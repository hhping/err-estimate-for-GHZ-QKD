`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JWHvWPV0ENh2SgFUaV+3I6r9JMl2KYBz7kYhygchSwjPzQVCmhjfvTSyYYZEH2E/
iRwUvfchhmWy9O9HBbHf838Nrl7WSogj+kQmG6nrNR4kRYu7B3ffQU4JL4PgVOj1
+vJJXZ9ZsaXrz4nCXxURVnLzUFRTwlW7FzTYZXXeixvdepN+DJq/EKflxzag9Afy
zJI5hfOLAbwXSf+vq2bmgLEurDbOR58qq04xA+FUvFVkMmpJlxAGYY6jh0X2qXh7
50MsOKUzrGofRfQydHnofurqxx76kZ4EZ5vdbEFzV9gWl5AFnnJSy2GxDhM6/fEa
swfWllvivzLX7n+ELWk8tdbcHh4V4qVE5WXuUvLDkDSrrRfC8cJsvoFQkL1niTzL
bZ3LtxxZ98GXqoHHSLmfA1/AgfEmYYEry+Z6PVqy6PWkbQQcUbZLXCy4pHr5fu5O
DaiIgMy89TfLH84KvO0IOTXpbqpGc8TJEZBZLuqAaaIvqKZYwLkhHZO0WSxH+fLz
a4NQc6ODGNSzD8jMDL4/2BgcEp7eGMZ/TiS8QZcvB5Z18bEGRWRqRpIcqoMU35we
Vks3whE+wB5lFDJnjnGXSNks/1VvnUbgtyIKcjAjC6aPBy2ZlxPz2lB50PXaqM6W
lTCUPs8BSlw13tOmndKXuiX36LDXiSrcYAo8GIcJRY907qRes9InI4KvfK2NQYfJ
zQZVWtDOuyU74wa79pqQjCNQFmGiyXqSPrldATpZFda1AuMcOANwCSjcI4p46Exz
t7qvXZ3tFJAYCWSGZcpemrr4vDIOJXc12TFMywDGzbf0bz4FcuLZWlTuWEs7JCmi
hN/zmSmNOJ/zM94Pb/JNCIyWBqSARo9ByaL+je2JdYkP++LHYSg20ddzmhzztrGG
xtolXp4g9MhOLF3PcoP368kW7OTAQtQcDV6A7el4Y1pBRi1Q0UXlRxbZFvxTMjoQ
NxAqXmfb4plKEXmWhbfWW/kw9aXWTI1bUokPAFidV0tzwnkSKrHN7PkLfdppX3EE
a/f52leYzyh/tLHCqlaZ5+Yo5t+FY/1KV2pXM7otx4XoNR9JhnrvAVK5DrnePA7B
5j05dGOJtg7Y6H9wuLFlsvC2w/MdI3HeNkDZ0rRyrW0Br0/5Z9Palo8tCQNZlGY9
yv1gs2aGARX0eK53eA4/5vMV2+5kY/vqWi5hlatbQWmachfmnIyoo2Ib04to2h22
CrWdpJ6Pe8Niu4s09aTQXhMineNbqZX5IkDaPNsgyrPMCRWFPWblL+vVON67cHzD
yLKBxmu/J7EPSzuNlOgmJ1U5VUHvBxE/Ao4jJ0SRJ+ojF0sIGi56s2BpYtnoTjJ7
pZSFwrgHZyrIxC+FhPKmsoHr1axDqMPhjMf4ONRg7A0jWXIrtl1sZFc8nRZ0Zamw
EXtrDXCw0OSNJSsyvqjBrLPl9mKtOc5bJlTDx7H++z/MMf9QnvEBlauY9McrjxX8
X+dST4IcIafruMIEji+zg+igPNrxEXHWVETbIjARB1PKgt2rkwjXe/82uwSXMPkx
20iqsWEum65r6dkGHtc5r+NB+wor6abf5bMs+68ZlBV+xlIiQPcjx3QCjHQhWMXs
mBvxtdgpbYgaMwuFWUeoIjVm2eYBNceZuzT00pLBkz7I0i2xTJuFAhZK48S9kF94
Vu6ch2P+W3WcP8y0UbWYy4piPFBOVrqmgQVDbk18vgonePXPP3jZDj1pTCG5WTby
Bfvd1TUBUCDNnQlE9cDKUrrXXRkgjTh7dfETbI66r0ret3IkhEMejOs4UD9xQWDQ
Fdn0FQQqG2MYH81Xi55gUvQ7tAvyMP1c/br8kECfo0l9TOG7uTdN61zyD2WBK8vC
TsDA+GHKkhy69hh5nnbe8bUTnj0nzxiX5EcRFMJiQJkXBQrpewRlJ4RUwfaFq+9Y
hB8BS8pWIBV0lrMmrv+SNaq1Zo1foKedaJdwp2UNbU10g2cQXbgMbjzUQEpTymfn
Bf2+i84x0MgLTWpnzy1f/+z/LoXt5RFm1RbsoYfuxGrfyEwGkVjlZJvtKB/+hsI1
Nxk7VZ3jyD8Fy1VfjOJ+IGr/Ef+Qcx+Ag1ozpUAkK4xpOt2msUvfCv8w65D4hy5N
jZ1am5/6caeXGAMmEzl1BASeH/ugTvdfh6ZRuOhx8NeT7MV0v7vEJ7r4zk7FDEoD
stfRy3DS10zOh3TtWeXt8veczEI0e94IsvcLFbqjgfCWSMzsqHhqtqdBva/FxJPK
58mTQK78bVZ7X5xjuKWzwtw7S1cz2ca1S2Q9Naq74NMnALWBAm2cFFsO0fETHN62
1SueG7SxYsZb368pstvpf3wpo1NgU7UZe5t0q+48yJspLnhKTrjqILoKW+YZfU1y
9o1Jxg3ueXODLle/kUhooE7cVJVnXoxw5upQhEuIIzpKG0QraLCKUm3yiWPd5Xwg
cw/RjxSbiEQ6wMgZRntgL3D0SGbYyakSAxS33lBJ+JMyDv0V/8JB8Rb8gWbAz2Jm
0InrMYaTKe7RX92+UruSKCoBDM65fxT4TkGLr8YZvPjb93hn/hIT17N5sXfo3fXh
hawjROdAzVOuFdZ+zsKUGkfToXrw53SR1nExu6STgEwnKrZkgKPr/qHk16yt4EuT
dx4iZkDj8/QjyMfi3oi4+fw1nwXnjq3gAkmuu8bJqMCdgCfYgg0rQvnr0BqcKO2H
JMMw19jduPQpY6DDarWecDQ6VUUSdwELO/lypcMN9gRxiHm7f+kN1erYU2jtehCj
ac5qEZ4kXthLAvKjTcwuNQLh8tEY15AhSl/iudd/SGPXb8USiWWLs+i2x51gKxNz
lOjQCCMsMK62fFY4x+v5gb3tZSZZkMC3rPbIQrthRzs4GbbbeJ+kmJ3s2RihgQ3W
hQZOvgqGFu/8vcWG3kppyHI9XZ6kbPZlISTrwx57ndUiCmQjgy6RvEu/urzKtBgp
PH0eI7P9XytIQ6Ph3nZFmwQk3taB/tCVKcJxzr50IFaAQSbSL3NCtSB37p3cLr6R
a8P+zYOpD335kJWfoybQhA734ncE2RT67fS19I13N3+Ho1XZrGRs2iau58W4muhB
725YgPY+vi4Ej6aYRPg068832qtfuxJ8wZmj9gHhBfqhqh6qDUzhNWtVJt9vQRec
EfP1KwKt3i7dDgwFcuOoAhjCRcV7CREAl15zoho0Z6zjXykAtmpSMywl/E+Xia8L
QybTbqCmLvaZXI4baL9SWZ6MFY2TSESduS5pdKYILOm3DDoooaRgFAH/y2OLkEXe
gizHtHqYHpuU/wR5FkHWxtB+rxRrc5hIesxhCUMsRTiHIzukP/lsuficnPKNmXBl
dxCyWRtzwnVYNBpfzGPEAtBmF6fsmZei1FMi6eRnklRo9CuedEkNOh+ZVEJydCqm
gx7NOWonZGVNNNfp3/ooXSN8sfnv8UKUYGjNFEvGp2Cbl0H8RmsdokdaGeZ1Ka/b
YVAqjTrHjh4NeGDszSgSUBQptmdpFPrH+NaSCfg9A6RQO22zY2CIgSZ7FTPlovpl
HZ8lRrqQamkduay8MqbPsbSFt12NxYxXAc2OmKclUDnnJ6kfWAHerQiMHi2cIpG+
3cghk7wGKQfSNxtpEGiO+0NPflIb0D2jAlUYeKl8sCA9NtsB2ZlnF1UVVgbXRkey
CMyWVVj2tz/PAdTjJ8VHQceNJnKuFOoy1DVEXJnQKkbpTwpD4JvB1ZaGJJRCK/jx
lyqhrYZASROAu6FTQuaqgb9IunfZ5WbOxEXDhmy+HEDwQAUv9v4r4HlPUcDYEPSa
A+8tTdiXVmcMael5D3kaPdeXGFPwRReuMhzFuRUU/DXp1VmuneFuleSTonofJLpx
0GVVHX7pFc0k2Kg2g9ZfIAyh3iiR0PoWJRUJkmAGz50wDpetbVp8HRQda4UM9dUH
vQgKxAlrCG7GEdO0FY8iwzZ10gF2LqGTGICX7KyBICkU1Xqq+qpJtqjdUiHsZYWs
FHUH/f14aPg8wCvMD7CMYHUDhyrP7JDQlVEktn/D+NXnlwERoPm3ocUREgApLcXz
xI/8afoc3/piCZ0HOZ5plq0isR4FT40LdSXS61//vGx63BdzAObF1hqxkEqqWr1X
wDNHYUMvoEgLGQdIRxszRGBzxIpAtiywGhnInyjLmlGsJgMmrxw95Cl19t9dZ3gH
t3RVPy0IZR9W0WU6M+yhEy+PSuBR+3BOxguPSRUcndq8uHLeXlwcWPJHvsCWsghZ
F37j1xzWkhtshrmfM4T64wxap6wi77ObiLzsLRusnszJxepCSlrHUYmglnIP87V4
2TCHFHSh2f7O2dXF5BY7y4XccFrRwPysTaicJns5du6SP92PrPOSMYUB9pVPBbj3
q0PFp106S+EbxtlEpjM8LGcpNV6MQdHFRnia0zt6404RKE1EvWjBX7UxMbJYUTNc
V8W4LxZzE57CTgGVIWfEYUbV873pzRvYJGn9D6CyIzAX0D/KX5xvcCeK91iNJW2w
CBtqn225vz19GK3mThaSqzRrzRV9vih3CBB3e0rjJDEVExCnO3kFiRc3bd4vuHo7
UENcmawHQQI1g7Db50wspti7tt3P0veSJ7XBg9Jwyydg5/JT38BYAKIYL2X/oKJ9
KK0u+mY2T+7iBDzSjlPMZm8f6QdqFro+2yTb9sWRdFt8Y6HAiaIFbZTJyzyEvjcZ
i4aRSHA9m6za+rlXXFKne7RwXJKKHtdjirUY5Q5pbB8IXRrUfYeKp/LBV3dEfQEY
itTeJ5ujDM8L9/wLnqDKSVNojCXP/cKf2Adm+w7M3aGyJo4tvSujvafuityylwl3
uJo5R3uOx04l5+Nv6kHFmIAGSyK74eRKffo7faro+i4buAaEvDoGRMnLJieX79NN
c5jDjtRf4OfaUKrecyaEmFUMCqVVNSD3hCl6jSg6+XZpplLXMcFryZnQkAoVAQn7
lQBGb/Y+sbALBEmcxbq2Fbmm3iHQGszWsjcAkJBJHJ+trKitmQZW1OnDiGX2huz4
6uJzNzJPgMfIJ7G0+MiDM4enDvkipmD/X0eAPH/eXK0aSXL6QGe3ha6eUcI9TwPq
dtfCztq56721cW3MTZ9xRQBfyWf4fndcMq3sAxy3ECiIAuPoe9iDQrRYJCm1ajek
Ba8LBaKwkFjHF2K2+r9gluTWt12CNMPSEzJy7J60dG9ThM4qLMQKZ/HQAvnUqPIN
5bEP1BXvbbiAxONTDc6BX9QMOEm7JVe7gqaoD5Zgc1Uu4dviTLvnMwpI4j5QSdrV
a3hUduRtioTEfk1/HLV1v88u1sngPmvfFF4crDKXUgodtEBi8uK9iPmvRD0NRR7p
rAC6UfKnpU2AIewagx26/rMKVHdFs/JhSebg9xen9i4bdQrrtx0OhgxwHfQo3RDc
GiNUMF6SfylARzOrCIklKSH2nUI9V7fM/4TU8Kn6qiDmjETQP65wGJHOJLAk1/IV
b59Hrv35vFrY4YkWA6v0BBoKPSQ2vV72YrgyBY4u6UPkormcYZ0EEWG9MMWrig05
wHgYFpy9iI0a9sgNqyaJgP2AHuX+vn1W/h1vEC2I0Bqwj1v0Ttkznb3t/bU8nc2p
SJlcTr4vXmIHTeSnxpPCWBcRsqB9rsbJc3vEEOyKdkVFA25sYajN8XELEsl2zLSx
MyQtLMqZdgVr+mMZtBsa7F1E2qEdh/6hevZIG6vWzhRGoteSqotU76C3akgoT0L2
+TNFKV2X/YRSs/KRJghd3lWfTX/wQMFNMkQlPT61YWtk6M5+vwfTzZg8I7gR/t7+
8uX5m9DoNUPD6I0ElxLaGCOzz993VpIbVfrfuvc/q5+1Q3J+C1I7KADP59BrvGjP
ROGyv6GtOJnVe2oSIrfhj+Da8aee/wCmD0+FuiOt3yjzPXoQiOBlOy+4Rziv3Adt
SZRDH3XQKAyfwUi5CVRoGXV0mip91xjTCTb2LIFTKUqGLM4oPCfzQ5L4w3Za/56f
DxwAkupsj5iwE9xmRFsEco5bdhmPYfn1v74n/5lZB544clmCWJbBGUjQN9FVNbNv
KvYfOWl78aCJ2VJ4g8d2uimy/g5I/SVgq9pB2dYRVbitRogKJHTl6bubxh86VBiF
QIhbdrusNs+zN5s8fwLtcZqsLAk5NPuUbo6XN/hJaSRM4Nzz0QSQuvGTU4uauA95
35lWJDFOYlCCJdntJMMHYka/aR+J8lJ57vtlyzOMwrCoy4bEAj8lgzuT0loGnlf4
+wXRYMvUeTRLW4U2dIvdYGwhqTLiRq/VMyR+bEpIsyX+F73VNP+ipox1jvdw/5PW
u4pUxQ3nSoCV1YWwqGppjmBw/NocztJx2RgUXZM8QCD21ZxSq2piQUnjGCgL/qCp
8ZaANqTO1FsSKgzUDiM1ZnLlclqyK6z79TXI7R94vMwpGWrGSPPw9ZtsAsnvzuRt
PwrF9NlWd5KckHw4DHko61dcVBjhj+Y2cMUuVIhL/GLKzsHO78N48veV3zze8sYU
8n/rwFi+fQgiMnNd661bBcwAIOgI3KsYD0bh14zPN2b7UXdQOH2EFlklA4rBZ0BQ
P44GXgMf82nBZ3m33neX8TY/vt1GwWWvQb3bxVzcHJCHR+kXQubFdXtTT/YrmYZQ
eQX+P3S1ehWkacX205pPs8IALudWvqPuzDsIk5y2cwsqnOSd3EDkhqjaVnx3/UPx
`protect END_PROTECTED
