`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ikFOBF0unDCw5cfJVtltIMvVZmcsNBQssMIVVeXT3I56Vjmv+rZ1+YZGkURlnybu
b/VX2tXS8Pyj/RjIkvOfmWGUD2L85lqApjuZdWmFTpRvxvQjZcX2UOSM8V8/chRT
z3yPHTYqNvOaDlH7GlODHVWdupIKbCjHlpr+yFBm4LaOnd3p2uN7113vmmPoloGi
gmz/Ae3ZAwuUKNLKGEfWbAN4QNSa2LU1wYN0/pn0lwRo+xPvVw33ZUOlfC4ckBkA
Xa1mpIJ7DaUd+OqdGXFcXQvFMMwyuHFszlYjoMaXb4+COGmXkxlPSQvqX3hPxetS
914aNiMMSNXr2hW4+TMxGUJdnyR8SGTQjg+eAuuW/FOFfDEIAhWgvSj+2kgTt9oM
YIPfchbYu6ZCMZaTnH6NqurgFQMA/ppkUu19EjCAJpSSk9xPXHM4YzOa0ODz6hd6
zIG1jNM7R1sXr5sIVRy1SFuNFRMwJGr+ddJ0ZdlE30ghqK3yDc5/o+xy62sRdxnu
pPFOIZqMDomVorCn99F0NbSnrUgIDWWC04VJmO/HwFoGOSaxICII8TClEApTyB5v
7B0dxWiCpAZGqqplufAmlFcxFNAlo4+Q862dOldnso/FGVI8bovHR6h4Hc5fUwr8
KJZj4S4tUzHEjfPtb3v9EIcIVEk7ThFHlfvjM+EbttQHkCxmfwwM9/OjOcnlYJeI
/hb0iolK426lpwJF35E9vE4F0s7gq5pIfMwtXIUNR6tzpiyo/KiKICif/X5Rv06i
MkSurIBEirIQyPm8/AkAR/WPjTmSl6wF1cAmYIsUOJy0kw95jFcLyCLdJrymDvsP
73WlOxrenvApMaRGhcXKLzvaL2QLry2qRCH8EduH2bunmwb1vokMVhRNyiFE2vV5
ZH5wi5VNd5ofFRSQ1K3IT9WJeN88YxeSf8QtPPkhwb+2F85lHLEXXOyHJ49xqZ2o
AGtxVNEb+tU7DBaNiHkRdSqzLYQ1S0Gccm3XLIY+pfh3KdjDLAttLpCOMPmBKPp9
BFsOOh5dZONeUSD2VzsnPGilqQG8h66FFy/gvzYfExGL2JQVoJ5S4r9lT2xBTYCK
/94Jrt8+abQ3d1m5BQj9mbltCZZ0K0aIeMZoa385+ZeahPDZrYob27oi0yDiL2Rp
H5CBhYB51aerNcRGv813b/66I/Qw8I5F5IDn6coj6j2iRe2LstsUit6KpltnERic
AQVNhiTv04xdJSvbVYgtWKBsowU1qxpW0MRFhk0A+c08+yqpZsFG/Dz7eW3WF00u
jntjsn/VdKV4lM0VaxIVfDsYTcyhVMwobGm0dPKiDD6c+ifFVWgkx66jHSiqKzZ8
`protect END_PROTECTED
