`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FWvXtI9mwno0dhwQbM6pQeTEP2UhjlmDsqQBgo2DYVuHhyWiHoIxtPJmI9UwXBxP
7Qnu85Ie6cg0yR5mgKkgtp7eMAx9IzSjyWXWjm+AJd9hHGFciZ/HQckRwE6zxmS5
iVFDjZzpPgV+rgr9QgEAGGqc9AbVzTskwWo1+zMxufdv7BEPzPfn2AVkAc5pukR9
TbMQ2JCjaHviU/T/jBOGFn28PclAfPfuthJ6KyLQ87C8asH+zZ6d2lE0c8lhSKFj
ezOOArx2P8UwqJRh2ZORtBnQxIp3YbSBlB0pJRgWS8jrw1VKP6MKnwWq5w9QWVtT
B3eeSPpA1E2L4BiL4xQPutVOgAAXLSMVfBhsFBbd99RDr9B7g0mT8Hn06HVQa+93
SC8xGhzM0cXRo6uFvpSRyZKw2p50NNFmNBfT6g4cJ0xk3RyJq+g0MT5KR8/SueR8
beJegaFX5lHwhLiiNZ1nMLbgXHKLAbI8NxPwSgXHuyfcuQbwpPpNJpBjIO42rNTL
Qaqe+zWy/rUOY5/tE9aDnD2pi8Xv8giYul1iyMfhsumq4nwyCWLvLz20mfSjCQDu
7PKfx6I01tIctamibI2RESupsqu3LjoT4vCTlXU+/5Tcv4lDs/hypaGwUSwwJ+Ru
+SwJi8eTX1qfVJEut0/QHiJq7jN57kxFwxU3HGVOLavSWMmLQFegdqCkqRt+7WDl
SMleLE9eh/10KUXAteRiKwsMqjlhU6zkOceadVuTkibbAeEnmGF0uB7DENjWRO2f
uvpBkaoSpLWQvlFdhqvSYuqXxmRkHG95jk39mIs8UXGLGREry0tdHzBs+cG9vxcI
6A9ncZSeq+nWq2hZrgwLPX73fxa8DxDDGDH8q8Cl7P1qbIiIvy8gsubuaQ4YELVS
fBpmn3peRQ3808w9p9Ws1NlJUVu/ZlZIIWDneKb3UniTO0FXZ7W1jOyh6j+hoGd4
7sY+cfmSACfWjUribI9QsAfDbFnWF2DkNDVn/stvNtrmxO5G/trH5abus7LbJ9bA
XuBRf0af5vtjOUUZ/v8yMLD2Z8Gh6PuWfajUANMDowAdKocv7cleNkkdrN7SCFii
`protect END_PROTECTED
