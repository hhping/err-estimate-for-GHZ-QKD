`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qe4d3OHHw6i13f+u3d1WAWAXR8dSssAcMMKZYY1ikX/oeaJPug462w5Z5QHUNLAu
PRgd1WxTTvmTeAMatViR8wJwTP3YFtOI5BJs72uzoKRulfkPAyretXPUa/bGrViS
mPI3TOlb0EU50wFC38G1r1/fXNvieb8n8JT2rigWp16vQQrNUYUSuPLfX66KY8wX
9aCUyxIDw0rp8k1JT7QtuEywoWjiVvE6lrw0vihEVboOmseStyFws+74Bi72vHL7
WoS5+CbkKtjFLm0VvkwRWp/dQuFx1gswySNelr7gjufQfeUekfdDV5i9XDRTan5q
cg+wSINhOfgFJsEac+TssekSttECNO7CkKsrpzAIan9YBJcxZ/jSOS3XVG21/YYf
bD38dLOnKL6f7WEc797duD8Usvgv/7TQ8j23GB5JI6LlHtibAZ24iccXXjohQ+b4
31t2vxvYw3vTN7ch5C3jMItkUaOFhmcDJ+27XbG+RmV/10TsLy5ubEAec4ITRT3o
1PtpPUT028MRluNHJfLyhp7tAcTkMOxecHXM/CDLk4sEY7Cw92w/8y6PytE5aip5
/RRbsQppZdfWk464RK8LGiQSS8LWCaDGBTQQRSpElYgkt2dgFO2Wg/ye6Jm0lYvB
ef2ACXrq7Yrcs71k6FOLEsVAqrtKclA4arUkBn5/Wtev+3wpSnuZEHGTJxBEsv2I
yheQhzHa6g0ScjZvEY+j8Q7JT9CQVS2rl6+W1TKm7c29aEi/Wjh1vZFknEMuialp
DDDbJP5tDbeGQIFvP3qkO43IDWZrdiYvIPGSFJNOumylZFg/eBrKWk60JJ1/76Ut
qiFNW32r2tLL+B7/vs57vq80wJx7D8ZqymOaQ4qjwTMGg0QAaU13vYUVXZal+VF1
gOS5wmN9hG/B13wEdZfl/wYFEG4YVELIKayUTgx07ZHrH40IkrL+n3gV/cHeu+v+
BqvPH2JJjt2b/C+APTjNUjZEYemlm4LJAAsLItmS9EUptiAGnolrO7RDHoJZMtT6
xzeGqDH/FXil9gH6AaR8UQUnYsIornhQ2FZj4gWEe+LKfwR770yWS0T2nMgnRlPj
Z4GV1RPpG+P6kteP2OlaTorOKK3eNgD9vuJToaeDNSQdznoeCf2IcBHRGbEYpWVX
uIqjGP1TuA65k2U1lAlQPer8/fMxkHwitLPKuZn1EbkPS+gJfdUZsrF9XBR9HhpC
IwhTR+Ko8ipZC/98BI3G81yu8vmyvYKtwetR+HpkVdewWzdkMrjZ8ZObq3AhZjyK
qiQafmZa8vM4KBarws+1o80YHv27snmU5Qyh9LIsxe1GTEm1vJr1o5jlZaxkOaR3
kRCGQofJDhgLG5vNvxawt4Icu4tg/PqxJl55mIq6qJFv3KyGHSYdlp4DjCGUQAiR
Rp79oHKHpcFRmrsa4DcZ61BBuNcscOOyUogO38EZoKCTWUVCBFGZ23HrIo/ibmVT
7gjMjNvBoiYfvsUa2inh9duAn1v8zfFxzFtiRre8FDc6GbQGEpDCraj+iTJHoM9h
Kayk7aKmPAZuo8F8wl6qcZLTCVF62ivIZd4GFaVRfZpMHQKV8aVgjX1bmohAti0L
ew636LxM1A3BG070JDgyH8lCQgmvDCTnkXqXaElvu5+7Dd1K6QmsQjnfuh4WPUtC
KxMSXFWBoh9M3WsQodFUFTW5UeGf3kmcVUkwS8Sxun1i9QOCbnUkYQsBrkayAmOz
1cx5Y9KH0YYfRaHZqeAiecArr/NC6O93qnkyswuHTPZvZ2daR83NyeWivrrIMFCu
dvfSQk3/tGbXuUeHA/QM+vxC30t3p6q32p5+AZnV93ySKP89NfgLz9rDwC3b6bTi
hYM9CHUY5P2CfceS5QAluAst51OPCcI7bBJu6nUeTwxG4yzVd3IFtQnAlk5q0ZxR
GQJ2mkk2z4suWSdrzCR57O0jGq5NoGiIwb3KfzaFZnXxMOB2zIG2BjMp9E7dwwpA
6fEPjdwdtf4f0Cw16LliVjsC8ghrccamQ+GYAgJBpEd/PgYpDMrNJDT9eu0nXJ1i
WwF1YXnkh9MkIXADj0csAyZXkxhsZhuDujlSpe34XBaiGJWonW+BaEUOpCsUQ07Q
rQhYRi2zPOwYVAv2HPHDgOtNoFzxB6tovxKEcT5oVub/3jjIrJN9ToSYkxFjOIhT
MpUjH+t+d8bdExup2ha0VoK+DMclWHL0NcglxPbtu1AGwX0/U9bz29IN4C4RMz4k
T2vkV2o26IS+0QzzcVTfZBkGjlfRcUSo1BU0ABgAymX2sAPIztdgjeHsIdYdD0h6
gtwMLouonOraKuxrcIms2skrHEMlP6+EF11qHrQXZ1wgR28yHWQiX5DKJ+yna3X4
h3KOQGYXVJaoVn8yRXySZzsjcXAtkyRbdXPlmm7qQqQFAHXPVL+NE8CnqLZD04UN
koicKzQ6Ntw/FIrDsal4pxNYmQkKbJh1HMKxACR6YGE=
`protect END_PROTECTED
