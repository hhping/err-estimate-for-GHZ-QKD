`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ss/nVdaxsESOs4wkz3HIsM8ZnA39SzohJ2nGbIl7rphekHYtdbbKreiUX6BPsuFp
dY0gW9MepfrvBvQQXyzubP1hRwdVY7lj8mshaqxbbSL6JgZ7RFDL3SiBGnQxOeP/
K71piKxDUy6BWL1963ISjNVeUlozcar6O3j8s8LSGReWWWgDkdV/i8HGAUwpb4Ty
CmTXNKqrEjq0ZPTegUeCzoizZ0t+Sw5+C1FRVzwKCvyRFAclbuqc/JGTelwazh2q
jhLX/ofOlxS8iBm23qsFG+tjvqNk4olf0GckZfDYEEW+ffNI6LTiyzqhwTmsAK0R
HMRtr34uVJy8zbhJ8QJUXLH6aV6jKaNMARE/kJ/VQm08Nzhry5OZk+jfE4oFRYZo
Jh3i24E1EaKXJI5Hs5ibQEV5uCj+QEmZWZ4vApVrJbmcGw8hYljUlHgj2mFuP+Oj
HCr9Rr0sgErVZ3/u8KOWqY9+0T9lt42b57zxuRRrDRgE8pl44eV1TL1zt7KzS1hR
cQJSY/HYQajGfxmD9SeCqi2hqlId9lopVBLq2bHSE2a76zTUQYDMvVNU3LhY8XiV
NIKKiHQTdyBhG+Gdrt0roKGxFv2uyZBkNYHZRpLkxQk8/6i2uOqplTtZYblbHati
1p3bM8eRZzw6JN29jwi0QIAyFtLkkN99uCfhUPbdrnuR6G9qBanFy4dlhJtytFT1
DXG0gb1OEntbwvmNM3JdG/xGsgQu40YiQPWY9C+28sM=
`protect END_PROTECTED
