`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wnk7FtBdZpxF1c+/S68AK5ZKp6wyQcFl2PjKqNn642OEBcNQpngnBaQqZS0GRsKh
CRpQGBCx1pJZua/ExPvNOCajgvbhh0fJ3VPwbXQd5Yp7UHenmsJhN9cu7gr+ScTQ
K0Jtm9WRCOtJTjgmClRZ6m6GJcBFZNbYN8M9BDLjA7qw8WiLGpy5693Q3Jzw6qG6
Nv9COCx0gf10lqcrz2RDC6fww6WHjTNzhm+k5b5WyInhvNWLCOEkHQtXIapinAXk
juP+pAZDFYWm9EnTVU76atlv1LPfntXxRRhiPRBMXMfNGX4sIkrjxiVvmGGpm2ea
Ckkv8eD5JdPlTDNDFLuU0Lk+i9NRGrZCAuI+SeNIwU5uc33gJ8QxBYKdVRoRprE0
EFG0KtTngUcq9XoAtWbnKXhNuDalnhqSkwrMiJ2yQMnI4L7isSlJ0r9GOc14ytAi
OXIs0JJgfx36xj5Dm4K3eH9mKdqoqt0dkOKEp3mI0kCB/9V8R46rEyDSwj0AHwnn
AGolui9wUWL+5oLi+cAzIQlRaZ8OXp6QoefJx2zwK/lOTyfWkVk2S0t0MwQPlhTl
3+KG3NXxYmQCRYk/t2zJzSR+Cx6gMPeUuFUwGLwGQqNrbmzUp4WanZm8kmuGd/Rl
QwfOjHJyIbutH/38FDBqdRGDr//xgSmTK/AhCLholpsiIOgtLKSLu0woqRzwkTuL
3B2Gjmtv9EdXeo8LQXvegik14Gc6SL1tDTlqTjIARiW2Yix0p5x98bpOUQcOZVfJ
b9bjCMtg77pJAjyfA9XWk7rOvXWyxxEozioqTqEc1gkslfnPmofeVnVTnjnzFkZF
pmTgwU6eV7WLGLo/+ycUuOv9u9r4LaGr+Pfli2uizfMIzTOdQXMgyVVCmlPsl265
hjWXxTQzbu9qgXyrdGp2mnggsf2r6RokkmTmDLwKfk6PJo+8ndm2z4jIBDmNhUf5
M84P/F4LDALU+Rnsc7KcM+WPWC4PuUJ6QHubjnNPWykbTQ5aW0LHnYS0mUwrQp2g
L1jd6eo7Vp4XE4rAbJOBN5TrPkIcKj+2cEIzXYPHz2wmPBMdnzpla2VprO76GhYF
EnSXV3H9fajIjBGK5ug9+orRDTVilg0YI34Bj1+T4xNhsKrsRK2YCYYuEBv7f7BB
NkxhFzlG7ZA8VruozcPtZm7PYnW2GsPQKD7tguc98ydwvDjNO1rxyoRRyPMUnMAw
U0aZPnH1CfYHYHEWZIwte5eBRFYpvks07sB/doRStsM/aCsG1kl5gcQqGtd+DLIO
k8fyCyf+75CMr7jCm92MQegbTRgLTSOsjLLE69Vidc6BkQSzPdhfzvWnCVrvGx8p
aqrRN3SGUqM3odCyvkrK/DkMtqmT6v1CujJWM+AUT1paFe/hi17BO0DQ//U1dw0I
VrCpY1xcPYohFeOqtNN6CAZ6EP7hJ9184dNoRfPvTCFJSlT77+AmkzmBNN0Lf1A4
huKOa/lJWZS8DGiM3wvSm7qGOyOJoJyl6pCCIOlSMir3lD/N/EZjOxosyCIj9tkR
5CWgbF8jpreOSjSKjNN0J77qYkT+jckAl01M1iM8RoAQkO49+yPyxbNzVumUElwd
A6FDoOEUPJCAteg/waVE4yTrd1kYPR2LrMkjXYhj1ccmrPGOKAYPTIrQCVS/F7MM
GUIQtLcN3GnavfNDCrFvNIdl00sNnHh38v1C1golXTYwCJpnUpeLRTA0buGP20ep
mAn2N48Dja+PVNXxbc9YaBFKwCR5ZvEVbjz6JjGr7VqmnNPiiYQT983LZaY0Dbmb
KbnluOJr5Z8ftjNRRrswJoibGPkh4WRQ1acn4YEiEvhSC0dt0nN8soIR7WlJ8sEp
OZc22ql/FNiLAewTDC952HBYhkzI6u9177vXmddEqIJzxHpy1z1TDYAmnF/I2IQG
vxOvk8Py9qkc7D8HH+nyDAaO9zAKXBQESxo3NsrIH5iA5hXfARIzFWbVVBLgmjyF
FxbgcXnGaZ5CWKQOhZAmpDwNtNYYKEwR8ijQYy70SaQkh7KuHKqtxquU/0TIqDu9
EPCCB/M9BCKKTs5oijyvL+7C9mHmC5jWd4pZgg4JAsNxibfDImw3/3h+b9ia7U4T
j1m+CQgr2t4kHiLm9xQbiGabrUrhpuIgK/ZJ/XvMlzwIfzzO6ckRUYTwtNkIKoU1
nuHOxSpRVdPOK78mm74hHhPle4uXpzCau6etQHXXyv7k1bkLz0i1DEjdNzCPHMlT
KhQOqTO7IWSaAvOeFhWJvPP71f7nj6vKWVVIPzQsa/XUnPTu0EiDt3bfjYhiJxwX
YeWp79eGS54DX5TDck0rrpRDnDhvKnyW/zgimYGtHbayaT8T/GbOc+hQI2mg2JUq
3ehxf3Yv0xkJJ1NuLt6i3aEgVf3l2F9vVdhKz1KselwWFm2yjH1vUhHhTNFxzwL6
qpIOywomms7nEcE2thp7AKtBp7GwrxRBFejeEsZNw8g9zbAXfmw9HFj4B2tIwRNC
NPkClWuvmHoP7J9XpMViNxrYThfySc+UT9C61I3C8XOWoNTBCm9bScKhTyTeUhY+
26PHXwHwUcY1fXk1B03j1LIS+fa3ZrNWoNq2LmLV5TzmR07R1XFOvegeOryotgkM
5FmlvwkW0bQdp9LMka/h7zQ2J2xEYjCKos6Omf2w4cT20dKSmAxFdl55ZHtTImv/
zoRa9NdNUV2UN22Yz03X+JwMV4nQ/eUnx2fqgy0Ew0BY2oWkxXNOWSwUlHjRGzAj
dmryS2xvwGZhmwrGrlRBqGvemgp4fIFuX3e6iGEGbZLnruH2wFU2126v3sc4UMV0
+qWTP03jBV7PvlHAzXLOJnMqXZ8wyhp91gcwbPT8Zd0=
`protect END_PROTECTED
