`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VvQu4B5i0qnG41CHYgj1H9ebV4b6ZSW/MscAYenQeD2MwURj3xWJrd8ladWQ8me
zbHL2etvdFCq3AGvNdJ/qRtw9CvxMK5+KwIQllUXNF0HPC9xmG16l2ViAGPgZCOb
xLRxXTy0hK81unQVdaDx/KlbNixqrqBBh2yye9AP7I6XuiIEIM0Q2L8r0eHfgZvF
WCRQ8M/M8lu50M++GcGFvWK1jb6m4h7OiDmRqwjJgddOwqPCAJGbu7KP7QTM07hI
ck+iOEaaJ6W+pOExp1NYRO2uGaq+6KRDX9D3+fNjz+uFUIPMJ6kXXYeGZtcxt9Hw
CVVE6cnWtPXxF0Xn3GVta+M8J7weuWtdouFqyBiEF8i41Z7wTfmNrhhznkFQ1lYp
P2WF1xls0BLKbFY57sJfdnyWw5A31M20eWZ1LzpAGgHxy5n/dvu3C5NiV2Udt87v
n623mnyaOXJ6xvezVChQXhjWL6WFrhjt1zdctJ3xPWiEobtbmmz+FfJzwkhp846F
fKSMOmz+Qhe5l3Qg+NfynUukIYzl+ExZqWh4A00K782We2LEgF6fTcCWPsYEgVcc
Pbm4Bkxfw30r6Hia1sqyjEYIBEbq5vJjp+FIQmOfKzrcCCWIgRZ/X9AQOSPwKm8h
a91PXDvYWO98R8lMRpGID56D16eKo5iZBvmmycn7fdlp3K8srZPrWUBMooKVpc2p
0aYChp+0L6jz5DXU7VvDK5kacVvBeURP687GQjsZZqc84WyHL5ArZZezVKCJjKC/
+4F7N6rBdEwoCt5o2v2kaOPo/A+UCUmTiZgWPhYTTFvsBIsIXq+lSCZooJx6Gbns
TZ/MuATFqh7OsCNP6rijkCcj7BXezEJzSp8zgt2b7UPeXBu+WI5NVCRmWTk+HyKF
pU9bI2EgyJaC2eiyjUzpou8yXhYdHSPfIPVjC4ehGRD5T2DypMcMQpMIgphqTY6W
fk/R4R1vwDKIhzRWueCsm72QVAlEFK7LMVd5jsAfZaii/OzosE5ulJ5xnT34ip3l
BpqFfCuYUrDib4TNHv6R516k8nnHFqggyQOSvvBxMLodpn5SEcmFfi/M6c0PBLP8
5sjfyZuZluc+Kw351Dv6LVhAS2tKAW0cpQqOuLLFGMDOP9lpsgkMXORmLcenaVIX
FUoMj3xyHPsiHertyjaZKLresdQhTR+0SOh/Izn9aWmtDtr/y/kEjXxbWpx3gmnd
KtkelGDH4cLYWvPy8YcJpjnhtlNjx6iSsQoURMsV0ighs8XKqgn+bpK0nOP3sgk6
UvwyL8/kvPkhkuihcxfOgISs9WeSZCcOGxFdvViIskHXAR/ak2nRSbjaChnt1mny
K2Wu+cLLvZ3r0MU3S3IMQRokNZOb3GEL85J3/3iOZHlRsKHkq5EnRtmwEllwIDrx
kSe2LklhZIcta2wQkymJbzlNtJjUvaXb5DGpFe6WWwalKtekVpIeM5iEh0NwgXLD
5A7sLnmyVKd7VQz9FzXEGovx+8AQTufJC7gDmnDUeO8EZBQmEPgJxY0by0CsIz3E
zTDm6z8f4IqJg5XWR1nNMg/7ACxWIgbNLvhPaGsp24C01wvZ28MYNrbUUSwH4uh6
KPQB3E0AmtFswtBNFRF2xldBrUrqwB6v+Dn52rGyJib74ivxAoguORXbpJtcSfml
pQPH54o+qFKcaPLsBebtYrjhUWcUVw5CIKLrJMorFGoLQeOubiqbK25Ao/8B5+IZ
u5yRJCJrjFxYauhh+xxDB+vI2WpewE8AKotvYZQTV5eN85PeotVv0al9xlCruHFV
LvbQ6446xGsgFrSERXZFl5rpO63pDWE+J+/HlOplo31HBS6zICJQfSVfPnGgLY6W
5bWcYgIwBGZFKG6Wuk2aayERu+eT1PosRXd+QLuH7avgER8xhDoPx4jv+dndnl73
6GN6r3bQYrLAKDXCw8fznymovyoRWDgf+25DU92LK9CHtpRICmUQbzXcgoP79Xx2
Dl/Af/+AjXpWpDUyipT5sNL9B2r91jf0JkXuF65usjgdUlpurJzGQH+ITi6KgBP7
FojhbVZzU97kAkir9dAiSqxfKj1AB7EC4sKLTH/heVZtFUSJDG7c8Zxjt4m1aNIc
IM0/K8Lo/325kfuGIB+fORviT59wTveuephVeMtZmRNE9AY7ZkMhufW8JIpsN02n
3Glh90MpXZCnNOO3pEYpnX3CXca6xXIBtHS1Q6fL8WBLqHhyTUID5q+qMpD+6S9e
Xnmy4ezCpgqdp1C75uC7wO4EXZx+vTstd5kkkWc84jp9zmlVAGF9cby3ZCd6PnBR
2wZk+2bzf5+vvbY4kfCw9xGYJOQfW6BDQvePI4svZRpVpTZA0xlFJhvnsChhyh9k
hWqWn2eDpBby/KJNiFEew6hZiirSYFgnrawd6GhgnHB06R8jMKUwqY10olCfGcre
d0p0l/at+GYtBD9BXb1S6mm+/brds8hr2zz8l1tqEH50kVHItha+/5opQNVQAORs
mjt2h4+L43BTj1sHE1UURSUZY7tx4eA9Pk6OqC0csSKJspZYNjfNZLuT5TCBzZWi
4DboNPeMPOfDPE9cygLaha2u3mbejHi0AG1q02bwhayzGHfR0nH+rSl9dtC8DbM3
Mf/ES5taKX34y7A3CTjiCABJ1k7puCFOtasXckN2x66RU8ab6ws5neqdkB4AumOC
PxeSdkbOOQnbZj7TajEzsuBPXuBorCxacXNTOzPWa6G9kQm8N42aShIualmjNGjK
M5G3frC88iAwkzVEcBS1/uoCUqXU6UdMNk8YhtrLkTnAwPWX+5k+hC2c8If0vWQJ
ODY4eCzf2hrWhwlJrIB0eI0HGL1Twy5fwQp5HsGqPrsq9AHUax8h7jPxffixfTRH
FG7CfJV/DenOtfUaKJuDuCNCb9PSMuDYQ4cnBj8jSgT/zaZSZquic5sFMPiqLwSB
m9s/QpMYhWtKh1x0yKZYCa4Bze22ujXq0n6BRV3fc/2yQ7F1SO3WzGVA+bpQZ5qg
BLUjexitv3Iwb4Ca7TGIKUedAQaghMjkPuyKAhy8jXXFmbCpERm4FmKnK1SXeZr9
bV4Lz+nmQwZVuRpg9MrgeyEGqZtWhfgcWy1vRLT8f6KEmgNwVWYLDPErsO/VILIZ
+DUPuKdnUu1397DWfHMsb9zrL4HeAJH77MgGD6n1YkpYMGDzUyWYQF92HKIVjCCa
8XVS0PXVmOBK5lG8K/zIbrtMCpNZNXjp1Qe6C9PfNPIWuoZaUzQ3/OIjn/9bq/pi
RJkQYMj8mOz51vrcRBMmq/5RKJmiJJ0WG2H28khyIAYqF6RuPPGxoRGzEh2tjAem
WdqxTrEqRtaZmIGfClccUv4vgqcu8V2nOfoGTWZUMs0rWYQIvOfCaLulNRnzibq5
Q5Qd8ESwpt8LUdeSTR2WPV0CekArESQsb8qJD/CORLtVbFe9ETqoCBnovBLaw+Zu
IvAx46aA2tYYEXAahbJyBR9aju8wJb9XzGgXlXht9FI4lTeYCMWhr7ziVD57tmlD
mc0tTic/JLY1JjSquhyGsXs33gnEZ0q7Jo3zXi1Opk/pD4SpZeWi6l009DNVVVzF
`protect END_PROTECTED
