`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3YJ3DjMqG1Y3KApEmpocjJR/ICH7xaXZFDp+npdnlRRiIV5UjURFIHEL5209NKkT
FuZzXMKzeJOWaqTF+0eUsv/AcfTJk3am+wENzq1YE4F61tvOtJEZ2DY71s466Pf9
M57zkFZ6jeKyxIKvktqXj2LGV6K/9kjrVNo6lbZu8y5oVRs7g5ukYgGpCO3fnnPp
GWEtXNEnN44jZy+hurt5mciVU0rSGjSWhuJQuilkV9Crm3HK7FmM0CPo/TKKKuJa
OmVKmsMvCKdZ8Jbrn04+JfdrSD/b6Gz84l79nzvr9UdIfVWUbVHlxvCMDZBulVwA
Lun45uOHYabYxR8OM7HRnMF2PdbAw9Q6nosAzt69QJG++i2wwVrqnIFt8+69XbgY
Hf+FrPRp7esQcnfQm//B110CmnQltMrhRY0bMT2zuAPsHBsuy0H2hj8Lq+sul9ue
lsFzXVpRfzo4GLg5V5AdIwGbBnB5NVzazXRaxqssCPhvEqeMxzBgmcFPkluXO5Sq
Zj62tL9QTtsFN5g4xYs6tqBSA0Kj8qt05fcVy5hVXLHwKrKDh9zV9DPnU99O+0oB
S2tFijqnTVh74fAbeDvVpCzKnfczgjEcmeC2Z9MI+rZCvx2iq7PSfgbGC/DEutgF
`protect END_PROTECTED
