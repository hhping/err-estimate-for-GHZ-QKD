`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVyaGqVVgDkP7mUuqVb3q+n+ChPnGoAnYdETyOimCM6O39ikqL0imnqodjjQL7FH
Xjwkow40CeyjNrbegjkApHiVuOUifLQlMlD7Lbb8fS1DJ6uIf9vgChWuiQUp3SbG
nBZjlpkuE48tub3PsTE51n/Pp40ZhVm8LHTo1SDqvBO44W7BixeNzsE4iNv+zm+F
QXgSIi16sqoXwkhd/rXXkoLQc+7ZygZk4WTGzy2sZ59/xVjfUj9fCqEYAdgqn9Gs
wH5zqC7vKOPrjvqIDYJeV9n+iM3Iq+Pe0NOh6E3UBb5epy4v1HxA2kYhrfhRS+c6
TUydiQtCuN3X/hUETIjBLmm70ZwSgTGXO8qbs0lNcwYw96AxExZEMOtdVwPd971f
2zY2+60A/KvImj7X8QqLdifQA0ca66djjbHGFvQ7Jng96bRgz6bbwgkEhNYekgID
iSqig+lnLa/gEWJid5qRXaIYS/u4xSzfir3sE622DprgwLjnrz0IRUV0k1pPMBow
cg878VXTiPN/Ng0y7f1HsSDTJMagyr0okLTgHZucv8/kB8TMbn94dcnx1AQ7aVYT
J3V2Juasv5OEECt2KyOJlJb6vtcHjDROwtycUm5N6Ny3fjBWRnb1gncSb07FSNWA
DrlwIlttMxNPZnSH4wUj7PxnsDrgOVyjDpTwOQrjMynaD7gUVXHfoxY7J/fhLdXa
cJxdFK2aXaZ/GnLo3dNEFBDTr0I8olDRYCQprsnGil3F6XnvgpXPmn/w/Pu0S2r4
OhWv0JfwEeOiXlvOkGwyYaINkVVwTNp7hbWWiUh6p6xXIeajtWB1B1PmBybi5f4k
+7NMIlD3MovD+jvXSzbn/yePiRYsm5iqXtmaHb0rxeLnF7IXRfRHL4FjI3W4ZTuj
dRoKscFbny1OSqsI+7bHd9xYrrFtjLwEKct7WlyMUtyeYeb4Aw9gI2x8LBgyo5HG
SOD7/NpM4J7vZ+bbkZw7jE8aPtiyRkgmdvWnyOWvZnbCcEQtvxh6v6obn+oQHeen
BKGnI/V3Na4GbnWXdS6YWWzkj2aDovF8foBKy8nRCk2Fxp8uQTYsC1gASHqkPKYE
WAyTZCZKVViRkS77ZvDJlovIj90ZiGBSVp08S2EvXOp9hj2s3wnXbxpgLojCMG2f
bL9q1+V8rLbNsbCLNIFB7zM1mgntHWZx/uearpBcx1m9FVea6NfNRAzY5iJvo14R
imbV8Gp5B6DMJaSUHAoMtNeus7MLLsI5ZhaQse2hyosZbdK8twWOFke8kxYPNgc7
IeMhJRzYT9B3E1gfON+rqvb5duT9paDXNZ3kuo/L2xYVxPZFpWjvqCS/znGiLLQT
i62PTf0mBOEE83aKHv6wCghSI+3ML231AB1rA8ohjPMpPsclDuQ27J7e/dU4tr0N
3WF0GcCpX6l/qjX2v/keq9hTaoUtYV47/Tttf62+2ETKJHsD9RxfuMwyrmXdNO+T
VjX2kztGTJJqGbg0aM+zP3taRH8+FQhHVnqpd684u7eHWInNkmdzrfdH3bnOk9aZ
kpPA5qBxIjpDlzpQ6IUgW9frGFErVkxmsECGkjGnjJayA1cJAJ7EmvVyX1fP+ipc
Q/4o5Jcaw6hl60lp/xTTmg==
`protect END_PROTECTED
