`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyiMSPb7SQ+Br2K3Dv8Aeiaat0aqCiwbVKfNX95LRleBanEd5n8fa0PMPx2Yu8MG
9cIy6jckQ5IlATccaGtIkA0mjYPfr5psYSg8y8xg3I/CuBHPWpmropar/ecn+L1H
/V6JbXgUirF4Ib+XB2Ui7NTKpHAO7QY/L4JPL87cVCng0lmXk77TUm66P70VQR/M
l5TZUBzpxDGV8lkomHsRYa8Jf9pdV9kn9SLFW2DpDa4OxkzuOwY4lEjUUp0Dcn/j
7r73ek4hn0KL15FHqrqnAlPI9RZnKehuFgN79fsv0uscZmJLvfLns/N7SqH87Frb
Cn3RKm+loUibXykNFmxTf5shSr8EygMydPXV5vyRFoaPVc2TjZcP9KTQVQZBEya2
IHcyQZHsSFUcqf3LFNByXnpYzaZpB2FmggALeYFnLDY/OIRcgje3GANqZWE41dir
L3nmZYEzG0zL7thnhIMUcYp0z+sL+e3lHaK4q5r0J9lMX7km1Tk4WMMpwnogfelF
H9oVkHv1ytCyOw6YRitTmHYyY1f5y+FDFoHW6Cfv0AAaQ7OHUKDOgn2NyufTRk0P
W6ftmKTJXNMNAvw34dQh/glru9nAMeUw7Ffvpx3mSa7sBei9bo+oY1SeAQ12OwaM
mT0F2pTO8osKUwtTYUePMbJloq/EuOLjDqVgOj4e2oGVw9qQjv4r5Lv9exBNjd0o
M8lW28CdBjDc46pCEsVtNCznfTfwG2a93o0QeKXUcAMUCaSil6cCVsdDGmxCzDE/
0aca5/be+CCQNy47I0TwhZ3NH3taKV611zv0sOJ3UXsHZP9h5idQSDCCxxS+jhx9
DahbW4HqjQOXxO7C/m1+fZnbSlnGaEuUX/9VX4rlWrLdMU5af+nTLjFhE9bt03/V
IHL70CIs2N3EKLTl0SWYiDWatqKZqkPD2s8pBg6hNSEd4ZzJQH6GeNuMBIDeO1B4
QOk+HXq13WnwdjzscYgilve3XWTSRyP776+X/13CFlxLe8wvhy0HPCd1o8rFINSo
rjR0e9Rc6rqlGwFIvc7T/iU5FGlhl2UPMCj9CoXs5br8q2tRysvtYjEZODd8ZGS8
PazHl7Bje2WxnzLQDKYfpdquAEMCX0LwPXiB4TBPoNstvjqVuxILEwDoM+YHq13J
tybjes0XWkVE7BZhdsGa4LxcuCRMnP5xal2Q2ZlhYadOAm4dMcv5yP8Jfkl63UL/
PaU3pMxW5mB/JMC0PxHGjsY6bDPvJ5CqZu3+0gi/Jzi0yK8DpnUQjldQ8hU0IRsL
gIeswUDQ9+O4YA/7HASEY7o9V0ZSxrKF8nlXHBBThBE=
`protect END_PROTECTED
