`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxHjnB7VQoFPwvZmMwzOPMbOQQryWZIZTESLNMXCNpOwVYV0kKwtjjHlH8FwEnxL
4b0hMFQZPSKbuixsx+X13P1CGTTY3YLTD+BF4tUIxd+3LOmeBhRIdbv8IBGOW10l
RpIEGHMIhdypMPQjGH9Fw65FQ0Zs1739OOY3tpw7bUKQcBdjfGbcQH2nQX01vZ1m
RIIIEmDt+ylC/so0C4PiPnDR4882MV3uuhXvBiGtJR+hRssbAJttTxQLvx6pgAcE
3gGcPXIUJXca7InEXI6RqwOylIjwi2tq+lVQ5gBS1YFt9k7N3NXvOCqeTIm7MYT/
Up/Ruri7KRBibEirwDMuhLgaw2W2VHbZhFQ9aQiuN07VcR97BUA3nB0uFaD+REQ4
r6dc6dRX7tBl6AzBNCzXDURMp/CFuqPqe8Zak495n/YWrTfC2Fkc4O33Vg3qzU9y
yFSzFpB69bDs4k3+JVZQhHWE59Cw/Jgi3QDWwU83eDQ9QZit2/lvDYG2umKVynP2
6Xp2pOqfZDH4v/r6xOYO8YFppNPx2Xvf90Azr8Vtetg0Lh1dtOrvteA+62w2S4so
fI8P4peAyinL8TUWxRqVU0+H07H15gQ/gboiAst8QFknTQeFqE0881oohBTwsdCe
DG8ByqWwO8R+aBFySaR9eyEgB68YLpj02R000Wgpm/MM8PIeCTELBqsawi8mPErv
0XimjGhSe7Q/9V6wtRXN9hP0a/Y6/pXweTiynpodJ/7CQZ4ec2pJ4FoeCfphI6qz
KmuxhzsYoqpIskgXmNfgswf5y1phQXri0brEdfybZmaJa0EVG81FOoGa4NALevF3
+LyrTWfwqMVygmZhNdO6pM/u8EoVeqYjIluzZzgTQaJTj5h4QIm5oddRDf8wsvrq
nh3CklP/RxEXkyweK1yK/lKd11Pb4+wcoUf0z20Mi3ZQaKedgzfurstjUgY7llvz
zRFmrD6nUJ/bDmWdJIzyVBukbSUeNYTP1sxRMxbnKG3xaU5VBvgzeyHQTWJj+TkU
/7faCL9whCJTpsaj8RPUeOLE3DDS63HHd5R7RtIxDPGs4qmoAXpoWQ7X0ZYlv6el
Fna4/Mjf8tVoqJ/tPwpzQzUPaiIDGudzA0Td8vTTxjbG3ZJlhTDNtCy5Tuval4Vp
Q29kemlV+eiq/gGXdvt52L9ltUvj4tFn8+kYHoQSZTM1gaeCsNh4NiMMu9izghqY
oW+8tfbd0XKE2i+WtnHnxyZMUdSguvpd6a+ezJa1YtQngvKOLJQOJxpCZAGVXaqm
0W2S1g2uSJcxkG/I8Mq/n6rFxCzxpSOje9rJOAnTfUYhuo/Hf4pploinTaHy0Fy3
fGWX+PK/eOCszmxE8FW7I74qJW3TciPy/Zzi2C8OZAlXN+arpKGJwJnGVM6nbrtU
fcw4HVp2ykkZgWJyuUuPztGLVTIrbLQ7QKBcB+6rKpFWntDi+tJCPRgGx/PbsOnO
udra5P3XbPF5gfT8rBYHYjlM62UB2RyALjmhZ7H4dE1va7wChBV5QScsqgNK2XnX
YO0i7flXSL7DBDRzRgiHC15J22Hv1CILucKFbM+X27YVt707lHq3wJuwSe2mL2ij
o5NFjK3KU4TLQpEhVe+wZ2s7hGKh/qfs2WnTzVaDK7LgHdHNQRJQGxh0kujKwNhP
JiWVo527t55j6WmpryEH5IyhsW/uLXRnYbp0t7rbzmOei5mcQ3+N5j+n5lEHmNI2
XovXurrJepBqYet9MiXY4sboH9lVS3/Axlt9nK6pVeaKg7C99guDmdloLvElEdWs
WW3M0fRKY67feO3rrQe6s6QrEXOWbBqyYVn+Vo59296SkaSHViZrGIOd4U4uHudS
M0715+p+bcwImRYJNVRt03wwzglR3CWFPq12iMFHCXGcBdh9RGTsDmO9rbPbVc1F
T7LLbnXptTFGCCEtghqnzCjKKJ7Qzr/R3Tvvua98SVpcglHddzwMRYcXfcC8BImX
iSOb6NcIAinU9Vj3loinXXbTCF/LlnaeM0OycRBsx8lIdvh493X3PurdXdIsOJCR
3yR+DFFwIZuGxslhwpvX3BL999jZCcnX7/9pByl9YdDnVcLTTigj3HSummYmPlHc
BCQvw79hEN6P6cgbE0xcmPgmXsS3HHR3YVrFfvjvrexofQIlG6JHZNeIMklJopvm
OHj8InoE8gckhQMa//5QoZUhINV8to4h3hMSb23n1JP7IflzDHc/rikGrlVtL3Qs
X4hUMHdqSVLZYPsdb5+Cu5KGxAyIDz3UIrHiKkieR4sqdv/xrSu6Fti71XFOKkxn
jocXSLK6K4oXLETZ/VaNwchV891q9pExg0v91IB19nABpxda5PD7zQURWIjn6XnA
F9NBvU6ZTW0S+KN4aOR8ngkJedYRJOqhYLmJH3pFLUtJ30LhVL4wEP+hDD08W83x
eVA6Yv04Yi8PpKS1ty53Jwckug7T2lsXjFnxyZensMIkD1mu0xaywSG37YdLjQjc
M4ANnAHWGMDAfNoV2PwSeO0E/ZIHRPGxb+YBcZ4QUyuMcCZe2XcXc4OhT5xkL3dr
2035A5is2ehF4L4vFufW+w0Cg526ajzTFL6kTGVzQWxL8JEQh3BNAUkkBY1AYf7l
48B7lcu58knQoKJld1Bi2tbRnje/0tcDzl9tck/wSQ6DzLmtRw2xM99Q/UDEqPhP
KixsRIHE4I9wHKepAGxiMp0BWk+F+qOXLflJFbSBVFM7ubjDR1+gPtNwVUCVyRwB
qE0VJhDpP8e19NVyUgWhlFTNmgo9t7O1SKXNTnZmDrWnulUKcU5RUK+q9aiOKA1Z
LyIK9eonAN7q/tUzsI5a+vyjgUQ+3vQv5rDs0s8ced/7ct+wtuPL+nmTieWEnD4g
q6v83rE5g+uuM8Ugdya/m8jDJZ3hibeDv99iz07u1LGJS8XYbFDExiKjUO17OZOC
ixGNLJmF7AbOtLEOsE56+8qkAuqKDjm3/YIZFeBRewlTxeQz438IWcAhPsvvLDNu
xXbwlaMW1B/SGXO2SQtUr0qoS+fmDOUqkzuFyyDllH0vN4n5toLtjuti5u/eo30z
a0kNdYGUzbc5nNrZRH7qNStB5M3G59IMdWgK8lRJyj0B64G2d+KIEAF8XpZY2rAN
7i097tbJCJZLQs1DecsB/8Iwn0VSb4VpAe4bJALJaC0APWpWd5obqjOamtdwYtNv
5SqNbVR3ybT6cFkDfURs2z8XPub/B5mGb0LQW0s78MRZV/CWs8f1DskqRtPyJARd
pwNNpMQVhQMFayCqu5WcSAbVxjFdusl0O+dZ0D3BCF9OFqH/xsoJECWbKGi54iZI
Qot4M55cP2FzHPOyu/ERyX3jnMkafzohmYHZ9EEIHT/1E61yVUv0vz6C45ECJmup
C4Tnw+iJ3FRYq5aswMxQFXdcaKBmT0TNYOJSLaI3JoRTjlv4Kj/hc76T/X92nVQr
L+qSkI3NN67QPvut3t/cljcROTh5QjauNy9cRhUdnJDkpWUoVnjz0o6g2SMBmEMn
d/IP1T/N4kYrkT5QS3D4aMelCXoU4CE33gTvm7yqjMMAtP1Jv/eFh8W/X9B+dqLR
UgaRVKsY1caTOCYvUAj29k+gD/gR4mYZLQy5t6LCS/B7fRBktnVbfUAgiHALyiTx
O/qQkFmnEqvUEsyxHV6I3Ic/rKObloU1zedyHj1FDRv67WppqcQiU7OLlOxn4ZUD
kLreS3eH1+zogYOnpUAiROiIy6Wv0FGwUwSD4SjRBu2SAs2S6ADJUyE6ZMUsufZy
K//+Ufxesx3iGNOLgIZZaZ1bGNjZzbMwynK5qmltk4+EiNjox49lfdS89PiniPba
CN9XfgVy0KksXFBECZjyhPSUcfvwQ9F2mL6yCmRN78zhDE20Iw7oWMQ/cj7nUcJF
mLrdz1+r9h0OfKUHNKpokwO/eXwV39Uu6fVzarKlwEm7NF2nfCehmA5a1LsoaCoD
i8nCx/j2p04djSopgobWmGnxvTxlK7whYKN6w6mkPqaSWn6McmeA/QcpQ9LeaXGA
kovtFZVT7CUDAidPLh9cp5Z+4R0VAZqP/Vw9tfKh6YfONkMSs4JagYk6qNcHGIt/
2ZSU0aSLkB1bwMzNMVsHyuoEgGJxlOFi+n/67aQEZ00YjgLEt+rztGi/ZGEXXfBk
o9WemvunySseiD0dMjQeS7m4W61aHdPdNn2BwXn0TOKlYP+1gUB2vAsTFfjX0p5G
NhqZyrYkx0UEReLXxIQup1YnFRL8BVjzUT4o6uwTfOheyAF6BIzmBhZxAVMc6ut/
5X95on7ylU/CbRdSBz26k33zaHFlA7paXUyhSXdlsOMq87/CCuRxV1yOE5NMBpV1
ZLw8bme3tE6q3qhqQUsygiekF+aXeB/ACK6f+sgKA+0iRh7YmI2fbaRYHYoBxoW0
vaZKNcWBcIw2yu01Fy7HVGFsCcKb7LZppT6obfiS7/Qv8pLkVf3q6K4SYRYuPtmh
zk8Io2+EYaMavjp4gT1a7Lkrpo65YhAsyG287cmE/8CpC09rVgiGjd8VgHedf1Lu
lkSaNawazH3LybDj2coyQYONzv/9srb7regAdo/NwZXrg1sHPJasabEjztllPbqI
vIVLwFYyO1A6VHUgOiAKVkV49cg8FWuqgIaiqTqgxb94dtfql4QDMF9nPh5FDuSp
siEcCctqA81xBQOpl+2ywvWMO3f4OEKgPw0Ehba+zYE7+F0IPNd+0bbmwthNtBCf
MpUJt/Fx6SceGFW9aZIkZFDzi/bsOU8HyOOYGkYt7z93gsKL349mKge4SGWoJ7rW
vn0yuKQ4iJhgmfwsEuhZdazx84M5pekbEz1pXNaGjg0bRwUJ1aALPuLkI8zl3ijV
DfNMszHV/2OlJiIVvWyp+4rsUxlhfkaFoQkQAFz/Cy9Xb7v7rYyxSYt2mU0/3La+
6yGPWB1sgi5Eg+pu2s/C9JCIohTQHpeIHEjTI04tbzESh7F52aCO51aedZf/TkOS
uUi0jBBguIquwYcuyXhNj72RDgHNvrnEy2HpVXyH1IpYkjymKs5PEAuq0kEy8d0M
4dVCpl2VqozOow+FdKRcaRegHvmj2D7HjCrj4GxIPw/8jbVk9m7qBFhjIuF5P7xE
74m5CuOv1SWXEaQWwM2+dLTMDnIQwkG8cB6yMKYkmchcm6tlmRtxGZFDK8vxL4nR
YqZtENWFydiy+R9JdRYX1WPCz5SyWAr+qLH5YaL55SD0Loe1g4WmeIplwOOyNuIN
RI+L7woVkb5QOpNzQEIQ8j84r4tqnlep2t9R2QLCMVI/yXYUtfqVj9iu2OjN6X+G
S7sILJfPMXexDNGZpnOUIDIr4cAN1y2vf90vDA6nhXAGuHS4JqcrRIbMueBpR3Yw
iKNs6grCFwmotBaPY8iWCh2f93Q9ZFQtTYX7CmT6cqolHdnSY/m+XBebQl2C8Ii2
sxYoBNMdJoGVvwcY2y7EzBlVFsSJaACmcu5tR5ZYFumhexmYfBk2ViRU7qMc9gYA
THz1mvsR2ATuT4bOrJiCz31Wblm0RroFMDhQIPNagR/43MHtAOm+fSY408f+Ksth
Atjba3Kzf/3WKTWnIDLfSCE5pO4Je8rWa1y3DwQVk1K218FAYYpTFKHzLQQhlnBd
kOr1DEowZC1+ln0184pWYYpnaiHGft/iWRBW+rSAWlHAjcJx/cN1DnYWDAJ+WVa5
47ZubDUoBeef5y8+ARLvn/sS9DgSHI3DYfdsWReOqjhuCRjlwCBYDBB4e1p56ELo
BLENPUL+/RwqM2dHcwxee6LyH6f0E3ad+te9aPVaOUiqrXrO/uzlKiZfM4HlfIur
DTb1hiYDBXgRU5kgJ07YsWpdU5jCpZ/4vK0sjnB5E0+6AADNddbihULRmPKSapON
FWy7oPoZMX/qSYIS3OXxmGruUyh2NKblaMnXWwTAmQPTbsugfiCMVb5+ebpFhEqN
QQDK5vSp7gDeCRoFzX5Y9mHaXFb926SxoKCmI1SKSjM=
`protect END_PROTECTED
