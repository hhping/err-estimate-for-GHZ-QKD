`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uZF/b2IAcLOnabHUwPr9/6PKQT2y7tH2bMNu/0wYyaw5EZRNBVWlFX9L65Brh39m
KuPdkR9eliaIwFgChB+1CnsGb8uNf4rzXM0o7eOkualPZ8jbCa5J44dEtyH84jzb
/N8XpekeHifUd5S1FUnDoRWYJSG/L9VtlkQ+dm5UrqYs8eUXXLL3KWB/ZLfwtqS2
4cClIUnZlnF3sxzzbr1Q0IoZ0jd6CNh2+MOj0A8bvj2RhOOTFWaTeRFAvTCKTJHl
IVy5kru7oFqAPSFfLxjB0zQBDmaqYvmdoAPj3xeC4vxFUEWZeJmQ+J2ex9cufR8S
hHgK2KRSVtD+0DxdeGCuO5HYp0uKKscynp0SlUaeoBW58lyCEzlArEfEmnW1DXHZ
OVaAZ1WKcXcf6fdJTIYSguV5BaMJrXAOkIXX0JD+SLemStd07ek75il5nm4l+l7L
JpTx+8aFyeQsfsvtsoKnoT8ilHrmiPqCPHOeDWWZdo3cMNsfs68iCyitn62F7jqN
0q1qeFpGiesNc9HWoQBdrdeB8nQay0p+v0GGhSevlD5Bcdf9B30P3Fe+ovt/GKru
u0zejHjIBe4T7BITVMvLrFOCk2LsziQzkRkDBphtKfCQJm5APX7wELfZ3lpir9tO
UwynoTz+olTQCh+NpXZWgUfEa+uA8kvC2fh2HGMaEfQotdTCpxR0WuYfvROIr6U3
VZv5KrTtMz8MasN8EtQab9n717zBLMRUUIQTlHo0sgj4wHequq9GwiqlJgb9J3K2
eLwS7GAx71JRci5fuyvdx/mCrElb/V13nMIeA/ecxZPglRLi5uqaFWivbpgCCO63
dHFGOM3d7BksNFSFN3Pjt+ss4+kgdumq0QTC3UMGk4QFbpXUoyFGbYUz/I3MlN86
zJxJ6Cf2ra2Zti7iBPao2OGWD9izxCK+dGJ/wTlVEH6IgqVOlH2q8mWNiHQw9k81
7W17sgM/XcU6jSH0P8JstommovGBNlU40PzRaCBa/9q07jBFLv/7joo3+tiqhVH1
xxj9n2tGsfB3F6UftvruixwuqA7BDsRhPQc2Frf6hsVcXeK7VZP1pStRfGot1qH1
`protect END_PROTECTED
