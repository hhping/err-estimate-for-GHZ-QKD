`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EEhYzwXUMOqoxc9PdSqtyk+uo8kttoQKWaMQ4Hy4V0HOu9+sXzhtucAFpvPPnp7q
DAodFZtnMrsKOo506dnK+i92Yz1/UbD8U0mu2Z9uJmhCuRIMw9m8BA3ODH4qx4t7
6mEkdg+16WYOYwBQ+QgLKGUMIxdx66F8icRd4mZEKPp8ZnxvKQ3GqxSSZFnPPAjZ
eLslFM7copLIEsqZqYc3K44/cBcPmi6Ffny8J0yjQNW3keyVnX7LRLv/sLJxKoll
4fMgQ+2/7l1d73lXK2k0UMW5XOR0+b40fSGRZFnlZonXWdFyqB7pJFS347+Qx8bf
l8CQ+UQy5a5XhfQ03nhC/CuwBq1NgX2AUySv+5p4vjDL6TwKtlKXt56Itg9Eox+J
7r7hdkHBYpJozQy22JSSsBZh4GF35lVNWti55lx5cYtEpHWpuUfiHBkfQlPUzxvO
+uweyeYhxng1xqx4sWAK62zT/t8skAsVra83zZ3ApGd/taemoRi5fOjMogbYEjcr
qpDD16LyBwkNQQJwG19OdhS33dwfRHxDKCpJlfVl1kbuoN/IN0oCU4WgEaCAgVxL
JjocEyXingfVOSf/YkhB5fvYkoGnRHqeG48zWVw9GOVgem2oVqfS7A8mpWrTIWR+
5ZWA1pZQQ4mVTET8IYRDe3sPrR/MRpaOtPKdE2w/TvcCoH7K49wJGuvNsFm1XF7U
2FV3urD7JDxSfLCOYJnif1Qs0PenmUgYJt0oPq1joWguj7iDQb+ukupQV8300Ckj
1qoHrMJ8mPd2QCP28Cnq5W902tr0i8PgnjBElZfVCRhtxlDvHZLbyODDIqwabDes
3UjYYnN6mao1Z+UpckXuL32neWmrGZTTcj125wYvsRps2qmxGV0mZj6xRY4hKZkg
1g9E8sscOCwm8fK+vWzF85OpmaYR7IzLm2u/WArniDc=
`protect END_PROTECTED
