`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zv3gyiST1RQxSY5TV3tuNfjEsOUZHlVewcP5CRhZUQKVOnGZaL5/mS0Bdmrkq+qU
6IzvJbUlwNWCDSN5sawl7lb4an8zsorH4lynAEaYEhhvSqPCsriXAo5G/CjyEvY3
yB8WWzgWUBtREhByxwx5moagGpIssQ4nCO6yptKrXG0l+vGxAA2OGp8VJ1OrUPAj
KMJ/01XRYwmVaSG0b0vYleDDoUywGE8a75n0fHLvV0ppmmr6yoYy91ZR3Y6ORiV/
sQu6AxmZ9kL+5LcRQ5nL5laLSI+yX/ma5TwSY2IU0eLD22tnj8r+mwO1+RerruPP
ChMnVLMGrL6aOvPr6QDf6550eysA/2cvZLAzOT+jfsJzy5WftlSuTf0YorAfIxFs
zreTnoxPFJI4wz6o2aUsZT4h7BgnqCGM6XGMgvY6sR741rv9gN1LxForfsxcdnb0
W3RX7JQM2RHOwUQNn3G5Hw==
`protect END_PROTECTED
