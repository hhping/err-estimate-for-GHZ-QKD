`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NW9O3/2cYLIA4g1FdHDi29oAxIHWOTbSK/C8N0j1pcb0l9hQW+/7+3t90DKafOi/
xILMMwPXGYV1ZgcHBBg8G5o+Hi9TsEk18xSxo63XNJwWV+VUpKk3RWC1dnL71X1N
LrpKsUnFbPz1yLWYOAouku2R0TG0T+vaLT2mfCVdST4NLP0yMEiOT3saX7AVATMe
xsjRgoGTaWVLa/UeK15ej54rfpN4VGDdl6C2RN2zZDfT7R07d1Ecy3FzVwFkJYrA
Gwy3KUipC8YQmh3MeOctGedcV2kq+njFVDy6o4qHmP7lKV120IQ7SBslURpvSyXN
PovgqpIfmrMucygtTbYi/vK/unxEn/H8H0uzmePm84xOM1iOZlTlbcJzGBzcmxGD
So5DItsJbcUHdzFSBfbh2osTgu/3JdwI8XuMvyG4vxH7Dm2ZFSP6QI1J7SvXvWGq
Z9bhzEBeBgkHNL6aVXsIBBMWR5fsF3eYmaJvWqnJA5e1gLreWId+c71oPM80HEiz
+9CHd8hTA3ImnmlGu7J3E7o7wy7zQ9S/d+YpWUGREjpNLhjMIPWaImk/I/3v6HEn
uyKXY5WlmYjsXvtZVuwkNkzMgV0t5FbhAfy3FgaUNR/5TCI14zwXXspJ8iL0yFg+
klOQN8ViGcot10GgFOOQsvhILVOcmCFRRki3CXXSPoQe9lr2AGyTyXx1SYG043v0
FlkMnmmLRdaOS2MebHGX8mFmX3uR50rucrUmauFjAfiiFa+VNS1EZQ7UrKmgzhVx
mLtQswiaiTDH0SGbyquCCurczsbzWboJcPTsbfQuMh3E20/DGXtw1Qi3wgMLsRd9
VmeN2AZ+V0H/jAPcUQPTREd+VjncYSJTzg4O7PHfgSgbyWWHKVvo2ODpUjJMf9Du
kO5Z5TFSJ0ngSyxmczs17cF++FIYUAGYiX6OD/8Vo2TDpl1Z+5keITu3LBI/6avF
cY14s9Ps6baBwcejZUlUePtI6Ui1dZ6Kb8kR+Fp3+xS+BbtfEkRjBsHKYBnV7T44
stxLSD5DfY5rEG/kb/GGZn1UhEQvhHJ0cRzouIdjIJ+2HnCGQNKzDBpRj0fC9nd/
ReD9rszkH2UeiKoSnyEF6sP6sIGImx3vdLfp6jYsPAGakDqTuJE4kDnSsf6FHi8p
7rIxMKHCJ4Ticz7h5HIhnOc0RUigX7nMxKyFqJS99bbxpJOXwpnslvMB3+GzFn3c
iYFZzfTj9TZnlWeiPA/Anyc0mABcW6LiM5eXQ2lttnMXakhO7Kh6KLpvMLtwD2K1
Q+NHF1KCjD9FKe23paMz75ORCGVpUty9jkn/Q4tEDMPqc+/VsSDD0q3NYTt5fzR/
BxfpZ5cJIvKQnIkF4mX7YJ69UQzuuPYBFlX5ws1e8bZ+7dfeO4jb3bKf72+QcPPI
iFF/h01AdWofe7haFp+XDTdCcAWiGP39v4eEEL2OEL8IQE2WjRhBLXgIwhyrLyMM
LcqjlUgbBBo7rMya4rE22a3OjKkq6PooAoiMTkiamACsp43jT9HNi93Va2SZosfG
nDejuB6JEnz+cZ1xJjewSsFOmqP79SQxYqzVgVEziYDOi1D0pwfqZT6GW1bFW6Ku
7uXxD08ReidRRHUGOXMHtjmifoiXrIu3auzQJAM7nRZng6ewf8CdPBDYMfqJzzyy
8ij4PagrvXbYv+9j5oOLPenD8dJ34ckPxgNXhiugo+/jDkj6FUpl3NLEEUdWkHpS
jZtWzzyFtztuV8WbczkjwyuWU+9bRpNsf6eKAV0mbBZ3bHVuajQANuiAZyd6+j+Y
I8Fv0U78pm31dKmxmf4Ua4YH0gAyld9oPbFNQCg1cD51qMpFwt2h8Xk3n3tczdeE
AslJlbp3P93GtB7BuNAsbCsJoZXwF6C1SPJYoQWoqHlWQffsT+4oMgNTLplxGAcB
QgpuBzXj8OKTtIPZseqOeNWvkY/ZIQ7MpvVJFIZHGwxjaC09zfBgb+2wdgszAAy/
wxVxVr6scapyT221QqFZpNIp+c/yz0g6Ay4RBnzw8tYLc/bOydgjfy4J+BVu+wEa
OqEX45zZkcdk0PUv4i7phwUvKV3aP5qARfsRZ+amt1pkgMAUV2rq00Gm46/+0lyF
cdt81/xrNC3coB19oFZ8qr/SzaOd1k4Cy8aId9itZM6SprOymPAYwLDASaz51nXQ
/fJxbuyqO84lSY9HPTke+WpAAJsj9qRlIAf2K49/+WTtSfzYP3odNoKgGTYuYiXS
mS6Fn6fTzUaYyr8FqMmKu4nUY4cmEckCjo8dRzx1DUvIuRbSPh6v0D96axT9M2UA
eb6Z5xnqFfS5g0kMBUgyYSj+94DhuNR25QupN63YN96rwRMT5oPun2kY9xo1QRAr
7D4SV22CWMXRvXf21fRG9T/FvMsOpVGqBO1WDwoxugbLIz7Y91K/QNluE6a60glq
N9cZOlKfqZlr2zRn7uVveiSe8laLUQMuIN2SR5BoB/zb9ZRJ+IIFJ9SdHSDM3hse
udNLlgmJg32Cd0IVlnLWIf7HLm3ECbVEYZvPxxLZbhVmXPkkZcP6cTfR87x7AgVc
SkhinHx+Rj3BKXzPEdyO3gvWipeyyOEjtDglZiFFjPWCLEddYqa3H2ZHCG9VzKKa
f48CVoWplGHeTRfoppp51bfKdbD90o95KAPqCOS7jr6/vNYfcG5xXoq6Sc/n7+0h
oxc7xUKwrea3ffVLIVmnsDGHSIGED49RI8Et1M4DINaOq48cW8wLNVP1cfbKAsIA
imwLYFhJS0mBJIeCH+W8I2nsFYCBg8JyVxIr2aHn4jouO5XmzoDShPvoh21Spk6j
QT81uHUh8Cv2vVioebXX58A0jh2MaxRYnzI1swkXOKqlit83LmwHd1D4uo9BPAO9
KPgJ2mdOaGSpKUQEPCngcjiXv3qeL/Ja/astdn8FlPu5snjPzABSLQXHoQ8zwrrS
cAjcmb/Y+hRi03YUCt+iAO316BFS0DAOGiJmUZ3/UICsqSckRsktT03wmrQ7aJXA
K7IEyXwDfr1Pp9CsPtwfPN1Q34ygb2ZSKZ+w5q8+Bs1nWcLwWB9bE96K/juUldAI
PSrVhGF7tcJLkkYVocyefEYOEkO6Qrj4xw3EkjqDytbuNV8UDIVnGNG54IiXzAZi
/+jcC+x+Sd3e00FFe9cLG/CrlnhDQD9akaYfVDnoSt24L8m6gIj5bmlnpo5hODjs
+hiwc+9qWG2epk81fhyWDICvemy/DsXJtpxXSFJilxj74qpv6Qu9pVxucB6vL7Me
I4zeCK6ehOk0hj2mgaI4CuNpIz4XD9sfFHvTKmzbbIHU44CdHG2NVLicRnJqNGmO
ocRTbE11qKc0Nyb7Jhp5NssPrlDrHBsCam0l4+mu6d17+WSUi5q1AtM/4UQPoNr6
BIP74wkjUuNFmjB5MY3K9OfXnWUGifP2L95vSmRz8KPce1Al5STMWFWgXXvFHM1p
+U1ClQ/8QAe3BQSy5y6kam5BRwViuZtFBJYQZL1FzVEO6iNjcTvX4bd4qZhU1f8j
yHvrCbTYZ/E+xh9AlXkJvN1SF+8VBtpvw11cosUIbwk47xluRpnO1SW7+opV3mDu
ormYTXmsnJNdh6VfKu2h3//DwLkfiy3FpZF4ime0sBYhBi5/+Rum6pX+joQV55m/
UXhGbFQG3nk8GmsaRbnd91jY6rsyxknvIdRdqv/yaYyeg4KaWYTtoMQ1+TYyfXnh
T9iMLrptLAL+lTSt0J/fkt54VByTf6Jfvq+ilIjoGzgRfq9A3mrLn2SvtC4mnvCp
E0gR1BJ2R+vjm2RfIwE5pj9zcyKYfqY/qfazlqx1TcR3rjYTa0OEeMYHGSyxSwV/
Ep5tFy/+I2+gTVsClIq4ITT5rt34Yt7wmQ6+j6dX6P0eoPxQtARbUgMtAil7C7us
syNfZdiNhUCJn13rANuZgomy80wbNL2C62VTqr4dWW526Hj2sGbYsCzWDpQMULsV
6D7TK0OOIfAjvnWTr/xwhGXuWWc6jPtVEu+XSy7+LMOZEG8qNS62VIGXqPHbtaLt
cvyf1TRvDfKYZNBheJg8j+t/QgOlrtBTHmbN5R4cnXnad34LY133EqozB/cRYeT6
e8pp/9VEtSCVBHLXyP+IHoiDN2zF7JPe7W/uqkonH8iFvTK1Qp/F16fD0clq3dQ9
qxI8kU5apnC7EW5INY7KOb52RZ+b8Dfv5fTYPsff7x/TN2Kfdykkb8ZGuMETPryT
zU6Ju0Xj6EblF4Nfbkr9WsAwLMwdAhLojHkj4+rR7+dUtt5IS5j89ISHGV6ApcH8
j0sl4SenlwDnLaKVYy0fEkWgdn83s7kPgMQ6wGjGaUiWzMJ4R/XYrOEp1fV3GuAH
TEkopJ/mCPag0uaMH1OsJfgBS9H6MavHGKcK0HZ/Qz5gRixOlCiYPpsxg+OaVUDu
SEkvU2wiCNiaWaFaWzuJfKJRKGB+iX+uRxQIkKDNc/K+0WcImH55DSvw83sj7xbR
9I/G6pLrEh5ID+4NV0ptAgY++r426t7SLlelsccopvBgRVYFYsvF0f7Qa55pg7vM
P+qOYNBrI+Vt2/yZZ7L495P02+jye0/+LlRLeGT09uQkFRkJtI7uMZ+0UYMFsOhj
38r4BIjaoYyF+sNBl61gcgFtuEhuXVq+8nrXLIFhqW4SsGPYBt7dCws+clC/ooVD
+Q71fyBapDh9rqTBa8EElCXCPRH5ldi3Hoq2u9R0t39f6CGumVdKxZZF1ZvPsGMA
tjtkPBczzoqNAnA1T9Za657N+GcJC/XbMv4C8hJ3ozVilGRcrWl6HHGQOFmuXa3N
ggMvqn9BvX9ZscU3NPFUwY0RZu3AYreLbw9ZIyuOnWiPSzEUwWKs5x8J0ZuySnRC
+4yoDsshDm+hkagjn5JYdyMbv9NyD4Nwjy6RE/fczWqduqYw8+Z1c+OV+wGkZ/FH
E5Qb767XhV+tckXWp8WttIs2XwMEW5EslfNoPUAPUiId4Gii2AYDiJX+cnFhPDhk
XuD3Gx7cIaEwhBRaK164hIO4qjBfV+Rq2n+oiNuXj8j8ozdJwJpT9eYC/M3OOkMe
kk7IyYXcB8LaxfWzzWmyyp5HXLUf35aVvLtrmVGqSSCuOySmODwnofodAudNmyjX
PoZFpiueJOJI0CSSTfhLp64/awSEc70OMDw3A1qG9OmFGzCB9x6G04jpNBRPxI09
YsvI16p9PkGNAzSh/VrZ3SjMsp60PDU0xj6+7QtZ/pEUBbKmUeFa+c/RLpynfbgB
LMuQ7eiLePucFIY5BXdIWsLW/VpYwMjZZwne2kYGfFxmu8GYFhck7NGZx7OMWYsm
DrKyPBkJnl/PDV1uzjlUFYs4jIjWRZrUK1WqZbiahKE9lZm+p8Vis75tEuyNQPdV
6S9M/FBySicimnBF9pg4ESj4sRUJeqBWv9iyOUR1NbRyal8r7J4eo+JKTOmLEv/j
8jzsoFhxbJRpY6bwh8oCHyO2kUz/nK1ONjy61MR4lLOTVCdHqMow29Z64yQWgWpV
QqsD879VRDl4qR9FN1ytJL5BRLrcLUwhhm4Swh/6drOpHXhyl+rXOKw/rhD/ezOk
JC6ifWfca+D/VeyYWPODhKARxp3bETd0HHaa0+Je6din2ZmCBK1dvk99OG+R8NDL
WV9I16pfrXMJGvcV9GLcG+fpJxDd7bew3KWKvNxtEu4uGLS2G7EynbRGSWUTovD4
c5JuySL66y3d3dBIjO0D2lq3w55HV1i+rTZkDql5/kvZFRrXNMTi6a1HAduHpLBb
78xZaO9IrPPZfahPjJywZHvEq0J8ls4s5FELWBUTqTmEKGPMJwBTEPjsOLxVqb3k
PVNIx0FxqM45GkEtBWnVJ1/e7Qyjo5Zw5XhU6FXjGX5bVKpqaT2MIs+FVrJ/mEHC
jmSnY7qws7bZnB1SRaJztKNss03PcsJXw80XEt7DyoBWL3MF1EWFihqraOkBPTNy
yM+nJp53On6yyCFcBQHvFfhpR9OzmSCEWqmMX3KfOlxX5gEN+OmCX+HXym4DrGoh
arTgO4X+VnV/kmwKavt9PD1LCCBwcvGyCWmOx58Lkh/mhOufiEECANXXTmFpMbiO
bZn0CVOiaXgQJDmx8bHVNsFRutLe95ZUSUxkFSQZQKVQH9cabrNwFHVAS/ImjP/W
sjU0uMDdCUYOtQuNdcJJosWR1bGo5FbQKXy1/kDHkxSGcWl9DT46Jx4HLWk0uZm6
uwLVSJJbOSqKNxq7+MH0ISaNA70NEb2ixbYwMFs+BbtLGHs/LVTPwuyLi0Vw4uUm
OwuTRCaMBqb0do9CnvhukhpHRv1pXvZqR109qNFwf8fg/fSFT4eTh/KjIHKJl+JS
0hVeWAmIKMfrkaWJs7eisOxRiYlxuh8BvZp5Gq3FxF6yKp4iCIauaB5NsfxFd/9y
8nLcatqrir5P6jUqom8/jZEC5LqOuCFMdkbv/ZqiG2xyCMtFxsXUCw/CIh/H12qg
B2REs1z0B5noOKaPBxcgw267+MnQRR1bEEULvAD/puzipwSkVCpBvksLbyE+8g0u
5VJq7Hx8GJBBvDGUuaAPoibgiX1h//yFX2bduPE0gaZIzF5O3W+x45tXNDKyB1ad
Pfe9U3+qRRm2uYd9NoMyVM9cuFzwQEGjbAB6U9ZoL82395pv1441+W0ser9g9P3H
9mZBerAn7S70KVhJ3rDDJSOcCCCpV81zolPT1QcfGKFoqz5cxIS+W5EItsFg8g7H
Sqyaf/b45FOYi1/WA9RBhB1tFmCu/NQOG2B5OOc4WHfGcwNNJUGaUsEHdmLJAvzK
uYhotAUUrkF9RBgGp3wyACka1ddxKsAN7hrxH1OqTOAh2LC1yalGysm2ZNbaW7cE
Q9HKAIt2OVeFscnSJfdVlBq5VhWO7+rg/D3T+6o+2HrI4lS7DxKT73mpKlfbmUXj
58mij+kohrhluDP35A4Nl6rJfafZmgzFxVErl6/ebv303u+uJ1THwjonPy/O5KE0
PzfyWKyzBYPiERMIoN8/SauKTvm4GHv4IdCFx3PFPB8a5d7d/76mSQHf+rRJFKBO
1Ha0dqRozNVGdOPPGAu4pJyGuuUb7J5VKTlRBrwG2Twk8mgAol8rLPqgOaISfK6/
+C1mheGXsd9AgNnf28ET7m86X4YVQ/81Xf955DQ1nTQi7Pgk3YjJmvn85tUd50nQ
qebZEru+z7FsQse/pA5dWyewp7Nit2JsQpmSD4tHSOJ+Z3Xn3+5MOYSN7vLLMKNh
cLfGTF7iKnwiR+Y5YJm2cC4Zzs1diOnKmKWbuY6iS19z7t9y+E/dmEjSwf3HRRci
720LIwFDYyQiZ4qS+S8JM93wff0gutWzc66ulXnhQHG76U89L1v6sFHIZ84R1ka7
FadRBKX0Vrq3ne9zLeHGfqme07CABZ1QK34Vgj/QTv8cDmR1blS11wsqSDltycEZ
SjMrfHAF3Gzy6UYpuUBIt+9ajR8ZqeOg7WpKCKuirF6GmJGGirNmZkeX1VEPkm//
Jwp+GC9Or7nuyp2/xmUlZJgF7/MIkVJ5pybm1ALXAlRV61EcwGimbrM3C1bej7Dr
U0ZGUnqIUjggnPUETJZLsHPW2d64XU3+oUEq+GJYzAqhgZeS6yHzDO00uDBGwhdk
PfsBeF3ZXP4BoR8qMU5PiO2cQ9geTpzMUU3FOZo7i4GflkCMQ2lb5L1D3ddV4Uvd
eVoXOyqBp7sNVHCZ4qV8DJ+Cxu5ftPUxzadzfiza044ZLh6xttPbvQryGLFv+0r1
G8wKAZ/rVHbHrgJZbdmFzFYcOoZQs32Cl5hvo53q06J/u5Bo4DiqieKNB85280g3
bNq2YTvJlQAg7EUqtQHGLlMULhqQbAItFLlYr+kRRNVshtJS97VzDy/YxJYkvZJK
Lsvz8TNQG5GJP9KnRCOOXAfZ6aagWqujF3G08xHLzmfcE9hdlK3qjrbvt8zl0c6d
whF6Ws83f5Id0oMAZlBmt2WF7558e4UNUCJkAoj++WtxJcIRDJTysz8GaiB/DsKs
pps5LCL6uYmOzkxENVfqfboQB7MEcyWILIva/H0G+puVCitV6sLOZSDu42WMt5C0
DW0ByAn7+gW6jkR09mJmtYKaMn6GT5AQdK90osgNDHTD+HXEeGiDfOhQigTXz25h
OliI8/ukylrg5ll0xnpN+hq2CdnejHkjDZwc3Y1pmgUcOU2bIDchWPD9N14cUVgE
xmJv/OW9BiVtVRPQNxwQqFBU7HxrWticYYRfzSNbuRTk0t/zrv7jqmT6EHmwVNer
VVhO4lsu0ISbQ4wCfZVV+kvPwpgiYarsQ8bHXdmHsGQ+vWRwObZ5lBQZ4Wl+NVtz
6lXHnnz4thfiRA59TTEJIIAdc50pjOkselQq2ZU0G6DvUS6oJ/0UX9xs0gmwCpl2
iDfdwlXdYdAzFXZvy+b7yqr1qS9fwFc+ORmCilAMxycdGbkTFmdY7uPZnzYJwKQD
qMxwbVVPFo+McaVsx2bNQr+WnP1Sw+GP7ggOcVXGvnrHEC5jrNEy30jSiOjD3PZI
xiEsTNtfa3xgWotAUwYb7pv5YBgdqo6kajnR8gpkYHnZqCSePsNnfE/isRLu7e+8
DI3WEH5fmoG0of2ai1mpEvmhgHVBGXVwq9WWVL3gSPAYrx9pKywN1OuFu5gkYSMf
Q3hi9AyyJtjXORndUG5B91eowMijUAZtuP20+5ZIv9dT3Alw1v1q6+dcJTbkwuBk
TWTOl+l/uxaZD8G1sN59uq18sdrJqQtBpuLPbNZNiYpLy0DhaPuQRgcM43Jc6qiA
1Pvf0Lwp/fySjhJjFY7FPvWXz3gUXR4ZjUvOvdWQ0k8yrASq3Av7pX20uhvZx5gS
QnHHIwE6bhKN0eLeZa5YrtcY350AxSvPW/sHWNLXWO+zsBFY9qvGruS/wYpCKHEj
R6zsmg9yNaSij7SLF97rfwkfodIM/WEJccF3FZxZnjT+nZCeyWWdGKaLTMt9OIql
w2NafKkvvUNiYQWZYe148T2D5uAGoCi7+ns3oTLd7yS9vmx0dB6sPt4IrkNDA6Z8
JEqgmS2v/wBmT1uoJ0cNNld3OkykbfqDXb3umZ9ekzdRwOQuYXvfqQejifcwK81+
izlwtAbAmHv3qGxeJlSjAHVH3iELrxRvT2Q27Fmo7XTsZvjfgvSibOGjK+ImHOCB
o0Q2sYQ4qkRDMckZLqn6OA==
`protect END_PROTECTED
