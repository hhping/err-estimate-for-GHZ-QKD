`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDK5UdIoBAiSTFU6HgBsutyov/YKgxVgEZv5KCVaqJwucAPJJf99r0GfsFDP7pK7
9deKyg8FVJCQki7LN5/SOaRbKF5ot3VOb4+pestsjvskeOTpY4gp6+o5exfb1Bue
wMatbofKu97jgBbvezmqRm/Q55UOzEeepDRGIIuN1Id5mC5uxOJgj5g2i9Ap5Wyi
KFPXcyxK3H6E9pRNRX1jiANoax+z/r5jj4RiXSZWnTyyRMk6W/kuyFWPHYFca0Vz
l3SzJqLle0vud637c0kfYHSGG2AQYwinWETDGA+Cg0pjK3l2a7zX/2lfWC51+9Kq
XCY4T0ZP74ReCYRpEu56O1f9rX8H3/RRWaJ8EsdgYdbTAncj6y88m9yZXh4zFYou
mZOS/+pK1xbvah0hEaA1aCLoUp/hUnedjish+D7bxb/XoFNh3zFvlePsuQ998Vzd
vhMWSbV7QpinFhS9neCfpvNTG6qf68wb/ZAB+dsqg3ocp778MCf0qd5t+VxB20er
RvrTGmstbMmu3XxgkRyJpfZtKGRrU+weCBQZPKe63ogezClM1GOh+/nHgnmG08dN
pdFEj5ej7Pe/xwNXh40asURWGzSd3vdZrVX7GhxoKrk1EcNLg+JE3cosZEnGSoaD
mI0OdaJ7h7nrd8C2c1ZgB5brePZePzfxeXOAX8gQez8rEPtSxyt3hpBIJ86Vnvvw
c/ABn38FRWq83pZkiiVHxebi7OYjo7xsCr+wU+BfHyDNhYu3kh+JIH9iYFL7479N
m+NjjDlXm1Jy7Dw1St+bclEcHkYJRVBOz22vHVTHZyw=
`protect END_PROTECTED
