`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wo0hfZJngJgyMLcBaJ3udsCVGagW+Yw01jNvYs6QiGaLZc5+UcuE3vBOI/PmCEj+
xcOLoBNYmRwyfyRqGUNkzDcaDQf9Uq4rXKqNFUEmn7fEp2g5e7m6nt5YWCz7i1dp
n3Gqwub20Z3lGJ+IInrMl5yFX72YvvaOR/KnHBygluiI+6MFpUaI0YqDQV/ah7TM
la3UdyGZ4LZVxzuzwd1vU/gUHobZt/6W82M8EQ075d3GWttjkKKbwbkJXmsMRLAm
X36RU5tNBSKNGTizwOzm1l+xFDLgOn9qaR/nsD/hjMXN3bFqCoWRcBpdflvkd9RG
H7hoxia0BH5dbkJcKge1a2+shl0pc3kWH7ObEWV3OERw4Co3KfURKS2WRcxXjcDK
ziF5EFNjuLJUyPP+nliQb+zD3B2xqMWyMY11D/qG3GJLrPKyLEcJQEBm/iJsqoiA
fNsgvLKH88zSrsHANTh3jiLvES1lZPNlREjSPyhzC/hu+gaODwi6m0KrOHYW5RbW
V2hEoklNCm86s0fdV3HkK854x6iDe6nMRAmQutywDR4G93n6Occql4ciZaJGVLY2
VSgkbeoh8/upUd+I/Ih3DFHLwNmDLXhOvP5CAUWWRwoCl4a5QmOFw3I9rHypRSlN
JFUvmmbc0HqrMkqXERdT8HNW9aznseln6Fy/UZ/batIGwnC0I5MjWg3LvotZ1Le+
fc3Bmf2i/9YCyUxUfRhEOVQU8qQ9zYV7Oz7mc2GGGHjR4OD2fULs8A3N4jmDBsYS
1xe6BZ9UgvIDJcRds1UrZWNBKRegUF4lom1r8PwE0vdmgeUXuxriqEwXu5jJTP0Y
DFKVvdmCN3XNfP5Mr6AURyZHVA/q63S3GXa5O2Sp2DzXvXk4xgbHDt3cifFgThIE
oXQpHISzMo6LW/jltg1EfuOEKbpzkEczFdWT01e7lQs3HRGjjH9sTX1SM7y2K9qu
WDdNY7q1lYxxtsSgrt+yTR+aVmdVEPE39DLamalh+6buFUKOLmZiYfGHlvN4rfSe
cZIcpxDtt2HoE8Eb2LC+mSIHUrSQqYQVIdlRRxuq5SJa9xUOhgvETycyI4b3AL9I
cuQ7bzmDIn5sIMyPVYkVwxE1ZBqDN+GWB6qKN4M3OHQFb5ew1TfLLxoRhin+JA/r
5LKauIh6NAqQnI5WwbZ2dViSd4qF/h5XWBKU3+KdEc//3qyAXqFFcmUoocHaMKjH
ATPC4bk2P/H5YjBnzYiwRktS2NPKHEf/I5zhOnN216Qiq5oBD2tQRmKmPEUB/dNt
W1qs5h4YQCGHcYUPzn+2r9pgcGnEEfOsKRg+rS0fspRpZcEao0cB4iPyzkE5NObH
YIOFG2iE/YC1oCfS+y0MA2QQcDGUlFUlYF2NgKHLqGQoXv9DRQmk1Od28ndhDgLU
vl/6Lmm09LmPdp5gOF61FooAiXJgqxqk+Wqof9J8IjTEHpHacQ6Ffk2qyHDydshy
TRhdsbA6OZHcf+8fPnPdikOvky/LpKnoz7pN1dlqgDXmmTRAOzI7Qw0S8pS1u6IY
d6vwpLOHmNYBbl9gBPaqvaFp1jZrq5cG6k0NxghQ0p+h/Hl+sQJXx6F87XvCWuPR
7BX+3ir39kcR5su7SMaPgizsVGauiAuSK8EmbL/zoVwz+vUfRImtviWfiw5NQ06v
aHomX3b0jEwroXqtoSuhAvx9rUXBEZJYD46mxzS6VCpB8VqeIo2l3t0kLhi7LXGd
j3uUUHJy2cn6GPeug9AYOqp/GHf5oM2O6CXV9QEZtez+c89aNHaO7KCszhgOS+AN
GFRVw1AgBpLzhJfyysOPeSUR/hE/2IBAu+V7gXCyzl5IuFs7KZOprnwg9MD+3KxJ
mIMZmIma5xoeTExUxRWqe60Ain6YRvqJCVDWGaFZKY/6CicXlv8rTpIxnmPcD1N8
gQfLGj4NfoboCvdrnrz8O0VsIpE4CuFpLV+S3AN0B4Hf/WODQGgKNIj+aNjsAx7P
/S6s9RjTrUmexq3af7IbK22ebr7rnI6Uc372K1TPKsRSVPqZdmCCgMpwNNT/Eg00
zyhUYNCpserYnGrlv40PpfupVzVqY8dKCIXHanmpM1ecYEv5mxfcNIJ+mcQCCE/e
3oR4ieWj5kRclPl3+W6tAw==
`protect END_PROTECTED
