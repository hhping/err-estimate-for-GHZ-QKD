`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIDRnyQ2rhaKITlOR2jQxrF0NQ1Q+ylU4v1dxm3udJzWW23TIxZh3sUkMeJobs3c
MZ6CKWOLj0+Rm7f3Fofps0qE8NuVH40hF5t937QHBIyFQfhQZmJXgd2bpejykz2p
C0JWqjdw1RlRPIze+KCjp9V1Y5kTOjfEIEjDDds+6cyxGs7QdOaYyM86ZusmRvPe
mID+mwcW6CvIBuogI5PP5yZpTqsx6dDFt22GwKCwj0eCpcptGkDAjxbg9Wlmmcyj
7t0pkpxw6dGyyoa1NeffQfsV4tzRo2oXu4TSzQS4P9Xb7fG0rpSDdfm0wEuUh+Zi
rrh4rA45TNsNfRBE8O9AFkDkcLUiVWlM+u8NeUnMsSNgX2Xbj0Ow7XTkfT7kyRZH
imvoyFZYM5ykMKYoq0QgQ9uff6jKnRv/0pHxt/CF65BS17pnbc7t/sHZh4ZQGRPb
yYtR4KPpS6zLhc+/nVR+K0VZiol2VyIkGOcpGiCl38IyaYww33f3yo4eL/nLPOEf
nnrItAyUlb3JpmoSX5evGuHXnEGGHQ2xKucOP/R19GbgT2uSxFyP9x/Z0Bis4Qrb
KofWHIWrXDZYZzNMJRpSh3XLnMUXGGZk0G+LmqSIm5POeN0glvt0/RmbAO1KQq2l
Hh4CUTJTKDH3IB4prUFoN6K/oWO/2Xwx5lCHPIW+x+4xwtdFEioFb+nkwKfM9FFR
xAWgsSaYBCOtqzpuMKS6a3NW9aevMxCUcW+9wyM5R9e0lamTUL05xB6VqGeavf69
A3LYEJbsYn6zyU3JrTo8J6ZO2Uo8BRLHvhaUbjGuDlWKZYSrKG5ZqpIe0xIhHw2G
odRk+EHFHk2c2iGUDuY8ng==
`protect END_PROTECTED
