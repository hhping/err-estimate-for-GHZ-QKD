`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPqZgNApqqke+uzRq5oPYMPFmUi13hgKVqjKBKZOaYy7i75SzMmlXQndJVKofWRR
QRSmJN195PHzE43JiggyQjIH2eKzfPP2xijo+nAfB4B686eFQkwdnXrnPaWHIhur
Y4S4OgM4TYJt6gYOuG7MwUG69RgYrfX8tMj80NXwbPyhgWwuTiGlj0PQphvO+5+w
hazUNzOV8WQVwIf+uzcqMJjgnKbteP/plD3cqnodO6qNU6T7Ff5ONphy5gZlat3i
wz3yr6qjivF2jHAQGuNyHSyM6P6jIigEbpS07k8oDlWXMChdvd//G/e5K9if1u3I
o/q2AfyE76YZ4wEpBv5EMGXkiqL/MOQHn6g/GEo2vycLQ12hLEqFqi+dxIjeAmoO
CdQ6VxA87I4uBrqEPsDCoRKC7Jb7tKBF4ckf5XvwS8rlZH38EE00KwrYjeD3KT67
VcN8pg3Fn4olQ+Lc243kyrWdg/UvvelAOTA6kPfBa+xWWLzkdvKvGVKJCoQnS0I1
+ybgWjBh2kvkjFMNR1l3jt5i2b5BfXAZV2vxk9qqoFg+20/LfKP85xhdiZQ8VHWo
4mAJD7IZ7nSQqyQ9kAfdI/1j4uzn+icwYY/UclszMXHcHMW2vCe3ZKwerm8LglZl
gwktF6YBIlEAxIoQbX6qYOsU0QD75BBNrDMUXAnIpLiFBVN2WWRQgjrlvHaTQAYK
`protect END_PROTECTED
