`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jMLJmIj8bY5tIKzNueSikIndtmaiPzqvVQxRu4c8FI3sa003OF15JFx11IfaK3j
ANg3XDTW5YH2pfNXb8F/tlPDVpwpjti0y56+izaWCzqZ/gQ3z7zm4l/d+a7hYQKO
uot52ikk72zfI6JoQ3cEZFbz0Y1e3OVbee+SW0RVzy4pfws/jW8m/0xKB18Z9R5y
kcGyD8DLr0O5i+QQe3iBEpRSfIh0GtlifJXNUdZvxNu0sV+/O9zpmMLJN3H+1709
AWWsVTFddcl+y8KX+TGxVku0h8NO/gZQn7pZX8jYdlBPAynhkDNG55LdGpDPGRkU
RqyADBRctsipSIWXHrrg8N1hYyiL7FJlWZtLqa3pCzkWm/AwugydAeJsMkg+cCWE
d7m5h288gwwbMhpmmNpxNsGOVsYWkW/MEmfEfIzVai7o0JyxJ6IMufOeVWdEgxpS
eUfxzQXuXIoopdNA6WnIBqUDbNenIkVpfddWn7mRa+cdZN5wcFrcFfs0OXmQICpX
YYPwp4iJlozmAYr4aE7t47oz2pm/qAgY05uqeHgc7KRoIkh4mWhybApmkRVGDH3i
3PHqDhyT5ESLXU5lydo+O3mV1UawK3NO31CiKRrWaWAn0IfWuTXnTn2GhGhbT0Pp
UEnDa7EB7JVs+0W+DCJivRDGPPSNGs/EvL2VvtqBt5pJhYR1YNrObRkD7VLtqyR5
QR68i7Gpc5QUy/7HfbBvLU+WWrr56XdKIhlTx/Aly7amN58PYfmi+sEtfICuNsh5
pqI+4cQa9BCKGhGta6JJQ2puaQSKmHGe6RBvyJxysm5q9Ao1O7Bpmm0Mv9Ym3ZJO
P61MU1Uwl3IpSpNM08Xc9vIbrbU29bJyh7+qCD9B34zJodm0ivt7KnPJ1mU1API6
uZmEa8ra96ips7frsvE/6AM3UfPAmbVqZ/hB0GohHfzxSsFYXc1D9BzknrnkApZL
lf4DWN7zsZrd1pIgaHL9a/9ECtOO6HNWEgxoSi3LnEjoilZMkReP6bhliezhF0Xi
3gvm3k2tW1b5ZU1L3VTr3VWYM0KwL5Q9yBe3Ud5hDC1iI0Xe24wPmA8wsue0vnue
2wId+WSryuHTNoxuNGeKP4TCIZo3npGOM6mO28mb5OvS50MxOC9lhseFQd/tDz3X
n0k1kE0nM38ppgoNM681MdogMWMWN0aQpQKc1bNVomNNx3Ofz9lhjYR2uhR1eCb4
fGofg5qolv0ZMHbuP0gEsbImOwnXr0/AR7dRDqe4X9VK/IqxzL953l2RzN6JdNz/
t3m8991i0GcBg+uWgocaHxWt9ghKgSAJGxO/lIUcaoQRrKwNrcmbd7uttAL9M8Et
5GRLX7zKAFJOTYABFUyA4wulRDfq6Ef3L7VC7gRfZYloIRwwU8WjKw2wVZeQPUjw
Hs9FqJkrfqfUMA5YZDHNt5b4IoVH5JmV2bXyqdBlxuaGm/+frU1DLqmtyIwUN1gz
2NnnY8Tt/vDYE/d5hznozhVp9kMsm6fgHs5dobOwRINL61s3reMPBHYNrVh3t4Xm
baqeup5Bch4mUNShYPyltjTgJHkYmc7kf1MOKkIN1HgNqtDmcc+xr5ls++hb4enE
/xNs5STHDtJIa1v9DHgzapuRup+ACnTqkr6tgiUB8qiQopSmzr2Pqz7ARJ1f4/LK
mv0yDLtprK3aRA47/JQYbQOcIGNkznxGchcNYo4h58Q+V4CY3BtW+q/kZwBLHnSu
n7+W8RYGQdHWna4hfz4UqbnYWTZ0dXJ87AomYgdaw/fWjcW3q2huza5zITJy6n9E
evyjh0IiOrelKEQXvqFyJl4LCO8L4ZMhyYkSx030mHd8N6mXtKsJ09VIMmfkuTfu
WD2Dfv2Assy6tMJGL/jikquZrA77B287HCsd19ETVvrdXmkFC2Wj5uwRFPSr7K/K
elENyJS7M7UtITtnxUu3DyLgI+mp89tCs6f980AKauBqQodVaxFtdULjA6DK+kmU
XiYUYs8C88yxutpeudUwwmx9gLuJ431kz7VjTW1gnsvvz73ZX/P/CfZXZrq9qEmo
HKgbUaBgwfxYvg3XbH9mu4oiQaNl92hmb3NzuWLz8CQVgqsNatbl3uirvhbmypyM
mk6E+FWKIycwDCFoX4Txf3ypNhfS298LlKnQfhYp/9sHLPQYNjyw3AFFO7joH96B
aOOHaWCcuXB82jv9f71fGoyvtVFBa0T5X9NLDf5KwOii7NJsw7Z+IRmvMcdKVdU6
iW1rfwESbCoqA/d/GryBE1wOY/hN3363bxZDPvEJr+D+fO0FTYGGla3YDHG8+CRk
LGCY6VuhAQB/dbeOzLPfA6EWiqlPVpJj1q5WEtyiLYb/obeO2u8Fv0X0qis/aJQb
7FBhUDMBDoNDjKKhrKni4XvpUP+F/HLwI60+oh4VI53z1g2ksCVHkwVnOBBmiB/z
+7URRBbbRRQqFwr0WaUXNimxw5dB8FfLVqJkK62Ly/FpCIwuI4kUBBbeya0SxnVM
jXVKU1IJYoSEsMRBBmr2sNxWZNrn5Az3IDr6JG8b8w5alVtebUzd6uXZ9GMTpMmO
wjSyKAcn7yKrAOdxvFDFRQSFVhQ7/4su0ovguG678PhtHm2zc/k+25Ff2xBg1oao
C4F9onaf9tAxxdcQ9vsxTQXBoWJbw7jaRYDB+y2T341bvwKFUouuDosmjzz6FJ05
3jNeBQ2NodfnSk9hqzcmL9X9FJBUU0BIi5qCInL1/GRLuPaf/HBVTiJTw/iNiOOe
UmzaZkiU+d+/BB0PzK1Z3ZCveiJSzjHekZ/RruOvvNmHmS+/Zv/RokWjZQ2tFrSk
2F6l8eLtjwlhgcyc7jJwxvaSmxK2mgy0YCbxnMgRYX7avlJ627UGUbMCYhxad+Bw
tqAzk/8JhoEoN4pmLb7NR4bDqzOSHandl5LPffDF3nbabu61s+BDJjk7nAu4Mi1Y
97Q5KXizVxz+l7yQIdnKiZfGSf+k5rAaxG1sMRo72z+6P5INfXX9t7wTyRPnFLD9
0as+qXwGask2SOSBI+g1Xf1il0Wgb59FcXAz4kEez5s9CBdnfhLBFYwKBtOTTI9t
zQqg9nFd/c7HFRKDXmVJVDwp1GPNe6ruEIutyQpB+TbW5yPvhCubbFibdKtwCOld
6fJ4mG62SGhGQ631YlVx8uKVrrCdeDcs0gRY0ypVLIBCeOds+M9m3d/ch19RFBUB
eZcuOKls/MPN0mXoKxyo4OHENQncUw7ZdhmhufBs1n8qo+bMKGCwMksgWGcsgxRF
OjAgUhzmywcHugioqD0TKGMzITCgsGyJeyJ5eEKrgWQxG0QmMsJXzUOoYnhv1ukK
wu7CEskeBx/6QmhU5wlH5qIalqvyln7AHLwAQMTNdnPYqLJV8SkP8VDotO3/QcHx
PCG+lo/aQFG3F7Zd60PSO6SkZoUqzLotJW0xi1+4uGkK3ad1ghmVoQknXpfaMn8M
3FywB2RmBO3A3LtaDyzIFgSSmgLAFri0+7GIJbcvX/8RBW/7AkCCwFDXkZVp7Wcu
TYN9nsiwAx3fWEdKyCiyDwoPtBdaXHHfr3ZNIh8ouyE788pptZOGahVPeQNYbAwc
3mQqaa1Fdvyvgjbbv8utGGS9XW24YTThhrueMMHgpxOLjBldoLjhF/3E9tOme8rB
3MH7gz8indrcY6tBCwmzVCc1bPw/5NGKh2CuRE17iTYSasZ5fybu0RQZ6ogNDZw3
V+aEFJt/fsZ4nt8QRnSvHB5ulKp096L4aXHMhNJVlKOeN1srIf4rvbTyHx5kEayn
LmxhNZX9B26jp3U5PHR6cl2URLSrZNEIwCdXzlCVwQYS2rkxoYID4SoOq42eVppM
c3IQ5oMTSaNr0O05abIlq3TyA2S6hGrqBIKBCnP3adjetOJ2CuYpho7/44CJrhD/
ADyQsNr2vInjJo0OdCjFD6yJgaLETTBUEGl+7mu/JSMtpNJBJmlDtOqwea++qQ8l
FAGR2Mny1gaUClY9H1juUphD1YJlAxnWflhbAbXcSap5i6SSxy4t6cyJA0+YLw8V
RlBloXylaMxw+AdKRWtUUvqhbr+4pLKDvhFqQ2noLcMGwE9zQd3eYbPbXeVVDVVX
upnmLvlieIgsXKovlthtfEKcurx/0uZRV5dVy56dIehta9j1sXyoxQyq9v+2lDHv
t1adApsLRzRWsImw1LK2GD4EypS0e2OLYi/Rn46vYYdTCBxE70EKKh4aJg1esmjN
pmB0hwfAfOYFh+mnjSFbXoxG/9UYGaD6E9mBmhhRLTBxsR+pAAenV53RmUKAuURd
TYtccCptIbjl+eCpgDQGGF74dmW0n6c5pGhiyKhVyAqqk+msiuKZVPgypcxAlemB
0xwHjsKYvOrJpmMf7U5NjZ8AJlk2oRTDicfyECNzkeY/kjfQ3YgEtuKhHcya7ICC
ptHvXzk6QknVa61VviMxuYpTZwXBzSDb7xWhP2xxuAuaL1BZF/YJeAzqctQhdSS5
t0jH27MQnYsKm0vPOvXapTAVetnMxS2ySlUF9UH96ZOkhzYbjXRq0ARZoL/DPMEJ
8Q/63zBHec/8Px4QJIS0WGFj0MG2dTOQM1oscx+2zw7gzRihwQ7lA2qf0XRJE/SL
16Unlybz6Tm6jI78KdfEx/rvgSJ8UORfbNJll3ynmCb1AYHDWxPPLwV48ZZQefy3
pIPJgeNkpPQLY2zTH9FcX2sEq2r/inDrpGXozmFmnuU8AhJP/n0d4Vl+O9m97NfB
HAt3ckMXlOjxj/Lu/Nw50B6OznQwQ78vHidlFsT/ZxrAh1s1dsGB0miVY3zZ54Rw
SglqxzG+2mx2O6nltX8d8HLEy40T5sOmiZGbrLXI0ptqY2Yq+WDm+KCYROLw1dsY
Ei/DQ7EeWB1xoKc9HTgSmfMWg8UY1FHrYo3MTc0BJWGfLRmBT2NU+SNP4SlQeqA1
U6du+d0DoFUo+aPxqpjf6NcFThP3GacRcLedODi2POR/MlEdfiCtPdHx0oL289ma
2Ni6aFFeUlJz0n/l/lxd6kQOoMIcriY66zVD/JwyGSWm7jh3dbFfKi+4x4Lw8TPb
kHdHdBij98BQYO82D0PrpgPfBRfnssG5etwIti9Go2UxhL6mdYvZ8JwwErj3hVBD
cRU5htJNU/bRZx6dVhlr6+K0FufeuCloZqJhjkKz8Q3jrMsRqu+Wc35jkZtQ/Ow0
MaOGSUAr9hSAZeIM5/V1EyMHXyWijDgL56BuukaI8Pd6+8OM5P1mC2g8tpZ0Zqov
6r7ugFIKEsT/AHHzQqCh0PQspPjwDQHwqDVwnYLCFMJzteCGir9hlSHeZeeWOA+M
pOR2rcLDz4Bz2TXpfA3DywmwgpROUBTs2H6vTBfuhoMEB99/pzV1+m16RH4hxg09
/WjPmpjkfu6RL7BMfpTMeNr4pk3m5bu+RRoGYSDiCQpED/nn473uhbScVNCEvdLw
qKF3lRgR8KXcgopQvdnveuK6qdFbL2139pmq0sY9bJKDLXtZVeFMm3L2z7Dcu8+f
Ip7RUzljuJbJYQ18JYZgG+syYyEmgeRxsEHmVFfGtRzck9QreUQlav+CXOyU9btg
/okgvTyg1rt/PORkKnuP1difjfgYYZLrqb/Zu2U3LG7a2SUzR+3lP1zXA+V/aSHF
h9U8gI675TCCAu8wpIc7MpKUkKVrTe+jUkRcroM0jnNwMsIHQ7RSsMZW5p3AhKeJ
NpBI1Cx+JOEQ34Q5r1byYW4QRta1d7gRu5MK3bzYulUETIVCtTeLrOpOWN0ItONm
5pEs2DaQ8DtHXbj4SF0Jw7EBsXSAhM/HhAJrA+/3EMFRlxLSUwcuYeyjLLZ7jHBu
jWVeETIlMUfXDUXfa3/aL6wtgLf/KuYskPV1+nkOxf9jMFBeu9+uRBYu0EiZAVHh
Im7Y7WnDpvNeep51OjlN9zk206mGN+eEG7YydFrtoIr0vplG/eHX2D97o4NKxv3Z
kP33dZ1h2Hgh/MZweTpcZN8QCA7FaSAFaYQdXKVCMId1O1glqOiGi3HOYrZVje+d
e5WKb8DRmiIYQ2tRUfldugsfEWoqkCq0nCvr5RPKU1drvzF8A8fsXVvFH9MLfpmC
x1QsCtvk2nrr1i87Riltv3xza9MUCHPrERLGxEJSfGQFEa5H82YBV3dIv1WWAtmf
OLSPUa1NUWrsK0rqLKP0vwN87k9E2DQ5UCXQ5+EHyvPvW4JMV4mcCBUi/S5VahlM
PaTxihWpH3XLGrr8jx/37ksEJdp3Lo/MIvsjnowr3UYq4QWcMrsQVuD3oIzkWMKX
gtjceG7MGcEF8HOE7tbgUY9yeSEhPgln7sXbYHuCMy2b3L2SJbgwbN37g4anBap/
fnpGeUKMkshhmQ6CFVJ4TsbdAuhG+IIlv8qCsDYfy4Jb5nA53+YjKVP/VMpEcMSE
CCWPeIL/NFJj1rm7n2bder88uaInQSwB1XnPKHUqay6p3e6KI2rroKk7KK2amOwT
IfqTawZ6B2NaYLTW1q9ImxTbVPxgFO3hJYZk+I3BsccjztDEo9B6fWvVexN/oJWD
p+9CzAO/290Qn7LvXjH1v7UIqzEzyGLlrRqKHmJSd0+DcXHE+hDoVhHaPLwyaNXK
vvax351JWGIX/z7dr6arlnQsU5BF4+69Jv1zUrEOz0SA9TA0gbT8pY8jnnLc2y3k
bA9D5YxCIe3EF8gEzn7jtysJBWxcnpzE5ZL6UmxPtEincPPo/KFjH3pEHK0lhudQ
9Gv+Claeip9zBAK/BtdN0L7B05NXGDjGRFi9KQxGCXZQ1cpG6KGsmKUPfj3BYLhl
+i+lF5CZdpD243EfvFWT+3mqXkl7r6tgYyruzaD+i33jk+5ZIMazwtyjkym3XB1a
jbD0f3JEOnihYl2cdruTLQExDHBqPnzcdKMNFBQALVakNQ84SWPxbx639E9vRNM/
JQu/I4/CCOWck3N5owY4o4nlqFtBuZUT7xAE+RHmDt9cMsOrH6hF3503yf/hpJaq
67IFNoKpZwm+k20FLosbiDwozTq1A8mI7RZyzAd2MRv+uGWCPCGP6x39xGnrHxLW
RqIGm9NWf9hmh2kEY2go6usZ+1/mI253fBIUGV5IK5EP43ceSr1ZakBjfUlZhZeq
nyL8f9ZvMVe27jYSZcQcU8M9g2ErSkYNuKxLiDrb08iRF5a4n4mHnUE6dMFSPg5W
auK3gd1Uok/owQpWSf97/NsVR3dctbKduu2oddzGfCVae/veWjoiB/FWHZEzPUAV
NmvckgTD6eokfsepY4TNEDxrUlPCUZSBaaAgqoJJ1ekNo4J59EDexnqWnIYr29mW
ujEVQeo7rRkq2AkDW/K4C8D8WVGx9NAz+KE+i+zuur4Jnkg1tcqrrb87GKJnM+2z
MDkdBQeDm3Hg6cpnHHHg6o5smV5+7l3lhaKd/3sHTkUWWbYHtbyOquLZqXvUq7UX
qA2xH2xz7U9Bi0zAxgH2VHcFvMz+DwP0gBGKWhB+Lf+GvF7TW6mAi2vx2mSZbHzU
6zdu9Q1Yqcd36fnQts8pGiT3nkne+S0H84aUoHtU9/D82FtBE6CZvWKGGTwrFmmf
FWOEwm7rwtCmMhMMhwxq5KWQhdh518H2DuxNB8RmEJHOqunNdUdyRUA5tN8Vb1T/
YHx7SzysjuI5ra69cOWTzhFruMEhP+t4kMLuVBJuVOZYNYNIvHcsXXIuYfOWKiVY
i/9p6DcwruFkP3PEN2KPL2I9pJEmHGtVML9GRw+BN7iQQv3NPaEvADb8rJ66euYV
9z1MoAlMi/dj9K0iF2tRs1q74Xzpbsm6Lp6lUwhQsfh5tDcN6HA/heaXV0m/R10w
RS5UB6KBvUQ7lWItlwzuNx4wnfxKtzKH1J3Nq7SmFL3YRJ6lhiVv2wuSet65Soak
tyWEpVJhs9bDJI8TO2ibL98uZa/cGCxkOc6013zMRainPzjGLxNLXzsdp/7/DoYo
WU1HP8EfmhWsVmxJWGDYdJlw1F3lF42uQTCvUpKChjK714+ZKXpFnWYk4/2ZI9Bm
YzfUp3WX9HPo9FL8UyT7PZnepBZ5n5xJwdnQBdnk+K7QldSCkppQ5Bd6iKirG/yq
ilbPdMUkgrp+/vD5nBbggxARf9vnmZu9+HZx7O8FaBwsZB9JVyOIdyVhLMiQWTPa
ny9uVPl6TjzhbLD/Vb3JLw7wmx2fx2vOPFHclcO5FhvdpnKZGtJRTnrX7i0SMqkI
fsjof2DRhA/qeuAsErpV9qEzqHg1XMc9Y4uVtWLOlgpiQ5OtnMKt3C9LIq4kO2ba
OxvqCJuq+h16hAW/U9HJ3Jm2YfqZiPGoUoZvtcmsGgcQ0fUgimwuv4slYmkdYiv8
T+FAPe3NN2Ua5nZGLYS29ZHTOt0A0Ym5IREgrCU/mHIfREl9tPiwfqrtyY3jv8nj
BJ6P4Y0WszW9yeAxDvWuS/gthaKaVyPWrNRb3is3mErulp3deuYwN9snluP7Jwof
yZ+xrFKEkdez1kkBklvGO9tt7ECQgdnm3f0YH2gVM4jKNq7lHoy5HCo7HIm47Yi5
Bxah228C0C0cMOHksDfeYvNQTTWCzblzYCFO+D/me2cVt2Qqr2GFXY1T2SwZNXwU
2pF6ME+3HGeaZw18x2tYYnc5emuZGm6L8YmpKDG604O/CmNkx0fXMJNMpZhKcdsG
UMNNGfN6oYvBzVxZpd7hzyyvsuq/a8wjp07AqsGCzdFsCkqvqvRm3krydbiWYTBn
gU/CN0mTEfj2Ras7MwdOwq+cOtgfCqaZ9juKNfhj10u66Qa7RPMisYT9uNz2Ib/U
ate9YBx7S6fAreC331nvP86/pBFyHfaZ6qONy/gb9cw1EWYRJsB1gerVqpJ8nx7i
TGe/NUrIxKhrxyD12ZPLrVHFu9oGCLGRE+UU96cYlDM+jB3CUqvWTf+zwMIZsoLB
wtBs6rGMN5WoHWijCIvM3zWv2fUr+ugS584nYEo1W6lxMnN7ZTbmhwmyuNAPoxbt
Ysg2YKht04KXCMwQVJg8MdaDkhK8a3U5R+Fp7FvhyEiopI5dVH3AXnJkW6b8vK6R
dWZu8th2n/me4aSqdLjl6+MOtwT49bG6bszdK4RQcXwGF4oNZqMAlhDSyPfUkZmu
bVnbwXTy4E8sqxiqtu8Yiy1TEw6HL41nyvzzuhpVhp8Ru+pqbDz6cSxUdZH+uzyg
+MkzvJwKZnPcxmMJvlzUOiPjmiWny/cNMhRsHL2paFAiiEX2sp9C9ISXwELdSkBw
bdZSlWiqLqfJpzM4nOx1gTy4gj0KXPVM0Ul2g+w0R4PaOla83zp+mp850PBmvAZk
0fvriAf00pNMbOUesuaxXYwzwfaj5qbd1QYCIG7em8YY8WAwGwmSSWkWoIWKMvLj
34cAipDeIwvWxnfuOMRYv6j/ToxCPmzGEGx4E1CS94Pc7CGBBOZNqXPJTyPosDUU
SGjwQkGYjDk9/hDyZvqPjcf+MWc+Hv8EzRTzfTBfeN2DHf9FyMVUfo1/n4BAf5iU
TBGpjO9QHsjsOoTBMk3tBot4AiOq+G5X2aB8xGQo3KYPChZj6PCjdoUh1YgKOGW+
tCRkis8GtjUfFGkyM6ZynBdEYC2ZY84U9tyvxJGiMmbRKw2DMtySjnqBN4IxRYn8
Daf7ULiExP3mCghmO0SjUet+GirhMARgKh1ksKyUUCPRRqePd9eS/8KzW8SrwSJG
LyJD6ebyq++v2tKS9XKeqJGjxP1MRwfsY4G+Jk/Zadje2HbVaZMsreg/hAMsA6BP
u0b5eur/jDr7dGbtYfvsSpn001kE2JKGYqwyS8C/IhHwqRLvYuVcjlQK7yJLqZdk
/pOktdc1H+Um3SWEaJ8mEMo/V69mk+WF9CgEzIjAhnzijeA4YFXI4kXbMnAy2G1m
lEXUtmf0x0zNtWSzyRyBaWChyGeaprHlkMYCmK0Ne6n6EZgeSphI6zu1ZPHu3ek2
2YrVNMsXoAa1lA6lLegsjLOuocPo1HMJo3BUk7Jo0J1IYsVD7JshlRwbNo8E9FZq
NNEHRLqdyJlerdCuY49HbaOauxu/Su3Z2jBWPn2Ed8bZGjudLDjNRfMEa7cLUpSu
JUMKlLMa+LeJicROFJuxhYua1GXLPfNNzRnOnbHC6UBT9okAvF6DEBrhEkI20M5M
hZhQIsKkcYgCHw7Py/1nRhIVR5YOKvU2v+JOywyzcUPC3+TghEHLD5q3fsj6+FYe
YLORRXZtRAfTD9vuQdXB820OZD+lBDWg4+s0Kk+c60Acod3FSU7OndNqkfQ9IPlF
AmIOg8CbutQofmhYfhawlw+iQwgjfGhvRaBGRTMfAcmJMCrpKgbV1ntS/0zIQdWZ
3TBrw93NE4v+HMwNxC1Kr4GyFAMCXNuaQD4B/gPouyqRNFg/HkP0lBMFqbfaTw2+
sR23Oxyr18tJFEiCX8aAf27BjDjQgrUF42R3IiOmXBCD5XWRAipx7n8BJm2jro5o
z7mCqpfjyUS4hZu6t92QMmImwmwhLhR05FDi8nB2nBP58AZR4H7CopvmVimBO645
EP1K7yixRpfZFXdQEDps0Vuc0lfC390pRpSTJlDokTtlydZPY5cY+A/0HFWULhSB
9Cg93G9wAjoPEHg3lPWz1t+2C5tyXx5plsbMwFxM4GmT6U77Crg5NgEqbbUUMU8G
mD58Hz2T9AzHWs5h0+/f4Zrfgun0MaO2Jky9lBM18/jHzUSKpjAG9tSc/bn2Rrey
qx8AQdiV6E0ClJd9ZUhEbTIwtSpqA9ptJEJ+f6TmnSlPfGYdM1tzWMj0LiklFYmf
AvcHSS/w3YGLfVV7UE0dv8jHBwFaWfoaaq7ma20Gx2hx05uINEIeblHJjTkNRjNY
qjHLB1XHNiIZf59nQ/DOSAPgpNqagCWD55nKsQlrhP6xHwZcoN0j6diMOGFMG/u5
7Ji6R8s6SL8vhtvSwJdC2dWPV13iiSKuPIbJe1kdL1GzTmqJP6/4K3HKcSmvCBiz
xCj59zxjgTJioEFyJbNoRYTFVepRcBj9t8aFYK4tmVqI3IbMAcXhRbMstEvbeGds
kIBkOCepf12pEMxABvMC4ZU5RfIigPeg4EcoX5CMmpNu1ZryMgxCeVu/gB1fBazN
pr20v7GyInfJpFq1yLV9ymr178DCVA2+NX0XqwGNx7PipZIyIK5CbHRB/oYESrZ4
mUNZguZPGfRoF+jyLhkQgsBS/W7QisoP5lA0J4rOF1MihBycvGHdZB/Z9ntElMsL
3O7vYWu20QUbiBfuHeADKUpZDf1Lo7XOjHBWDfDMOyIIBHw5CvO7JvQwkG0zRm6F
Olchst+g+gfkwDbgrENbPOSVW7lAOzW/lGvwcpOFFNAtH1druPI7QPuTsydsqwYb
rPY6yKz7/t7m12hVCR/6PfVoeVDszdUUwWgcMmux3noaIeOLPfZaZ233UyzTQ0Bo
wQGHm5lsevM32PJGuOrAzUORw04QenxxrkAUVtc/2PvHOPyxmZNxsDUtC8eYHSZa
U5XWvexuLKMF0M/f1Yd0GT5d1Gh34aaSA9hCMnWpBof4HL+kit/EHIC2v35cz2EZ
gA9u0g1nxy5BDG/i0ngMdBJicRsUCd1n4il3x9xfpUVqBHAqYyFE9YVLJWk57WlH
slGPxhfJOYYupxwPLTn3C0VXz15STQ/Iyna+lyl9TYZegEAtgSLAM7ZQKzSsJsV9
AeVaxVWH8DTgjoqyQctGsgfaqsOzgDOhGo/m1XXSrMjyoj1nF1DZDjvlLoGMkreR
NmAfxjQUqgWJ0zhrqE2Sby1GeKhT9UBApV9aysgcHJ3+/qUPqdE1Hl5W+YUknYHX
EnR1ksJTNl9hRiJbeJDHRUTGQmxLfQImRbmYAW+fzzqjX/cuiPoGgVwJTesFXFN6
uyDU57q4dgdYY9vhuSLzJh7X2h3FMCH7kZVgpjUtQlzHZaIl9PyDdZGqEAXKmF79
YMzXlOFyel5cjJPP11TWRQYrdfFlPE39mR4gjigSaRFAmmqjFsNrJbcXpadSMt18
G+zXufsIZvhjpudt1tOpd4k6TWTBXRNkjvBtUj3un4O8sFNclme8YZk49fQH+gbV
11uQW6ocYOstL+kHAnJ5FV4n78G1wDIBf60xl01cLemQTEmddVwB0094yWZBQRh5
qAKYTkz6MyZqIZnf7X/1f8pFaoBB4sVELb+yfZsIeBACB5eSw1ePCnwJrbKB8msX
RRM3/tpapip1gqnW9NEvViZw4jHNe98TETqbw2BSuL2iFHapYlyzFciuYIGgVSKX
Zlm9K12sNJUw2+WlJO3fCjBBxbsVH5644azoo6YFSwZzKGbqnSQymbixTFYFMcEm
9VcKENCscIoTNnMD66cYFeelp8PdJL/idxOk64MEVaKEixmQpGOs+8fEsGT+YCC8
P+0iuM3aHFGxF7qSqArqi+nwfdL3I3OKLJLwOEbRLef/iCADLIaMlOYyeU7sbHOY
b3QZhINEFz0iPkj9cq+Y8bQWx4RymBD/xHFIQELYs6sXjTIdCbqYkPo2hhxbiOxy
MgDpB68Oocgyixb1FDKJE5IzuzzlUu7kGCmGb856vAxQrWlZJPJ1bGiYEAodg5Z0
ZK6yaICDzwJV3BgFEeaxYE4ud8CoUyOkHwf0qTh1+IHJ4qH/MwXYT1qIXqP+4B9C
HCjsR8Y0D/bbt4bZrKQJWyHb/7RleP4VClS906h/HpkxKhkFu1iAkRzgKlwYPsHF
f+BdMsLaC5nAlNO7z6P66qrVr/cwwxgU6SOiY5qGLW/TiEM5VzBaX4U8eaGmZWov
8EeCKErMkNkLHODdMHSciLB6kINN4l87KAcyv8K5ePuCOzPWTP+gH2GNIVSfWvle
nJZPbG6fcOp7rOV2hiLiH2BEYxkQYXVZSBR9HbGDCvjbDSKU95qYPM22WegVQI1f
EnDaocu7Ehnw2cA1SGIf1jWCNWKOQrFFdauS3L3Q9etv1BXgoTjBUP8WEt5Np3gN
jfgBPuuYhfAkmVbJLStmG/hcl2t8Gr7ftXdyc685inJJ2q8NsGIc6l6P4+K/cvqd
6cF+dBklelRVSD5QZD3PwDYE4IOZ0HJybEBo62jvk6OPdlPoSyfsG47hKOW65Vbx
lL/pLEo+kk0MBPmxEdQTtWWkYLxk9l+qLb+qP8bAo6O2ck4NiDKI0Fxc1umvtYnT
soasIQjMSQAAx0rHFxH5PvuHUpbJASUehtjkpIYgWn/YPevRQ6H3m0L0Fvds99Tp
04WiQhLPh/6UIGo+F5TtloeXCSd/LuQU22vHUsLWmYN4LsNXxFHzEDjeTIk2OWCK
nLxOMJN++sxLBg7BpUMTBnezdrCkpKHhqvX899DXAsWSaocerciNXYyf7TDZRmq6
/XPQBYbJfEqhcDcwDehZbRrNuMuVF1ZUIRYeIqEWZWuZ09ekxxLK1yq0VUyXChBJ
aNwzxHhp32Tv6tJHwDRdeOyiR7m9FSWBhUycKxF5RqMudbgmPbxA+/aCOJQBZUOM
sDw9VrtVoAacjyhw5F67t/Fk6zgTQ0V6/D8GT2GYBOAbBim4Qz2XjMEfJJRpiSUx
XmFXeJqqp1TgOd/xqpZXzlvbKPQpee7YjAcmlEVxgziu0aCkJmERY6plBelKQKyF
gJU7ZdicPnCPrWbrRXHQvuT2CSaN/f2DkPC1lzbkuQ2S0ILbcTrM30Yiy6fdUG9V
N9jLCvlvfockWPxa32+8RrqxkTHxPIymncIoAH8ZRiwW7sA/GWxQ9VGG+vN1uWo4
r4Prp5DJ6J9PKy9NWYCbhCQQa7c47HModGqR8PvnTYBlOk+ZxVywHt0/OHLUF0QV
EyF0mXcBSefARd5utFpG69yhrcY2y5FlyJNMJOXW6twQ9fiRBhbUtKetMmocYEBH
E9VYpK3vWGm+mVr14odcjJD+WR4UtoM5JBzwL63H642rs4Doc7e7l8HzQcw5EUP2
MhV+DPcsrvvEeZH2W9ANky2v/jRkRacaf1uHqr68Q/LurO4RwTgemQS3YO92kn5n
IqZTwbchhUMRkty2SUid5yY8+PewIOX+9OCs94muQiinSWE7TAyk7klcBFzQ06oI
XHrEMrGKLoA+IZwsMj8XPgiIgQ4xC0FbTbsmYDMQ424bb9d5nQ7R04B4u57EvCnC
poP663e63iqwUl8CwxSZokJQ3gLvFPPeSGVumi3eZrUJbHQeHvdGb/sEHfSNObWc
1IcAyr6oiVWSx0pFNZTuoYYTUp6yAqJX5D34thx2as5ZSZRwWXGwQEs6PXgw+1fH
1mIalqei5an5vU/9VDQ8goOthdSglhjCdxyhVSAjFzPGwyRCXupcZkTnjR2Hqfu0
xNs34KmEAfEzNYzEbgvFjpXR2KdqCNGuVjIcDyIH7xugZzuB/1SV68EBK9FOFjgF
Se/xluv/r2obmJLpfDHkRIFln3nf73t66J+4z6CkIsmflDECfQgqzmsuO7f+AQuo
XmQDE2JFYIVamBtulFD5ahr6CY9YhmQsI6rI5cz3ivlWW7ZbNG/VIWodeJIMTesp
x04rIjPZ441Pg4mIE+a9NtCJ8XPF45iV1k2tfdE16qwHFC5SoAPdA4ZQo44JxWP4
Pb67S5m0cd2knOsf+RmxYnq3qyB5naIVrENkCv269vp7tt9gTGIigdlqNRPOYKTi
fVET9X+gzti4bzcwMaIdzDsN0VEh98eSdMOw6SnGA9ZsQi+JIlOeHkR1K9G5NFGp
P25JsIXejkPAex0QMoiXm7wlW/tV+DsccYg7Vnp3F+k72ZjGwjiCELuGdBWdrqON
z5cRjf2d5S589O+wdJIk8orirpsXKDSEzAjL7BeYzYDUcGH7COhzjyhrVNS66j9I
meJ6tmn2IVTMndyrSuqGuR0m4+q3IRANkDPo2+hj2TfhOYSA/eD0dxtkcW0mPcgv
2RnHrWvcMU8cz5/zBgXmeXFYduxccA4XWov+2KZknApom6TtLH0c90rVDeCRWK9s
ILt0FrXLYzzHITxKx3+4ePpOyvJJXS0DRAixXohFC7MmDxt5BAB6FXK/x5wbn2S8
WbNV+iyxskxrvIybVUwXHQTt8DoCbNQZCzaVhsvmidnKh+JVHsHuzqBHMft+wlDq
EUoDqzxiqB33IPuXJiCbYxIuNLkggFw6QNXfH4IgCfSEyRz40PmRKx91DVkOQfvI
rVtLV0BDOd6+jH7GBGx9yWJMdhOm4k0HorFqbIh48LgV6oAnHPDCkdJqpQJ5JEul
ML9ec/HEuxuSB+fvbXd0gCllFUslmbAjTtU/1J3ihAiR7yaFztbkf6GlxJalU+H0
K23lETFRHYXFsTDESQS5sEAGX8CMACdAYLqpoUX9qo28m42UYfIL0D1txnaTh/jg
62FBss8Zu7gOfeaZPuFB0+d+fGDPsLIi+21sj5rlxHThqdXXLEK9yknFr/pwrAzH
uSnUiNzptkFjPoGyFDrwJbo4PAEIONj2aDBByjeLqTprX1RLhq8NgaU2LPB4cQUg
IDbimRWPaZflW+fE9pPpcC8sf6j6iKGmC8+X94UL7gwUF1Y2XEnP4ca4XvNXT2Oa
bVT5dzu6LGStu6D9t0nFk5T9HkQ1U/7xA1yE3/ZXX5DJmImh+jygXlIJEKx+XQGe
z4zpWnJ2iki+quwxoII/9g2YDRV34H7DBZSguiQFTbI2yBU668QYjlhSDTN3o3Y4
Vuyy74K6tdg2HMr6ABdwhvb+NBsJHDWO44uz73ikdFhhoR6Lvk4/CoSfMztB4ZZO
MflSI8MlelFo/XK8pe1DBbT/XMGlGJqVt31Ux4C1Tvc2ZXPTQ7u8+tv5EMvCcARx
ghYfH6W88AmsfJNy/iDz3o4csfW5LA/oMjXXeZU/yCdFLM8XP1uYc20qIjeryeU0
3g5FtdUfdTrtcgNPGFO+YrhIKb1BqS34iB02OG7NwDhBhGIuHO04gorYdAeuSt8p
q0S8nZSkHwXCkS2AFUgFETCcQFhxjSLLZ1ZhCW381Fsd2TVNlji+Cgk38QCfoc6j
Y5l1QwqGz3bPzxO9e1KlF69lTZTq8dsAKAJ7kmpX23VqHxlXldaIlhjZVbHYpS+R
kR9VG+MSr1CIa8nNF2C7N7ArmJ/lFyn0s6N8wEysCDXeYj6CuTn/wIEQKhSLeahq
o+CUAK+yNmqoxRvOQcpvObwWsg6MUYKZr7uw4pF09KlqhCXw/nCTY+C01l2u7/wE
UcwP2u0D5XlmpYybYjKp1u0+tOou4JcTIjyIdImIOYV04ugj02P65kgPAKcgrZaH
LZYrae4EKjTJKCU9G+Eb4PAihCUwX+zZnkySD9WVGIUOWi8wHcWTRou3mlNCw+hW
zL1E7dSrlyM5bgU2fXj//hbxU4hOw9KNuyaYWC/xkFAnHGQR0/z+sOoVDwAIp2v/
20bsrDervEldZMPk3uBMgUUWkrA2Z8sAZoJct4WRc/6gsIK3jNViQFN4J9G/bS6t
y0cE9aKAJARcjUMojk7wodf4LHt+Lqj6QjjtNB657xobp0ah+pfQm9d8zbEb5YMU
ckB1QpK7f9c/wiEwSMP/k1p6zm8wWoSZmKEUDjDm77vExjri+mjf1bHfXSrKBYb8
UaTWTg23zjUE55F3ml4E6Aj5rf7XDOTXFDbvxth1Izh8fVyvUDrrAKegEp07DECB
SoZbQ1X+z6RNpYoNkk2wJPilrFPeLQ+2hwZodTwVQgITgfKUYRzU3d4v2y+1aMZP
aquRENLUgKrqDMgU24zR10iqG2S65xloZgtI9Vhw/nk7UvcJ16RrCWRSX2k1S56Z
rwoIQ4/SWqzb5gQ40of7ke8+/aCJheo4QblEknSePP//nA06z92sYbEcg6Doh8LY
EPLJAniYBHcxZ2su93W6N1oJqa2YPCnsJ3AZuborXORPdHvFFzNg4Hepzj/GBibk
MGcpMzMBDcvnp9+JjZzO4NN5Nq9DkCFjr/7hmkYCzOdd0AaWgxEW5yLdSv9Q219/
msnuBF8r5S9/x6VthAlLhFKkhNQEYeQu2uYOki0s2mACjRQT5ir1FPtWsU2OnUGJ
tYnulzqGqTSK9VsnYeZeGMAyZiQEmRPphfR2LBtaLeHg+c8JfdT8WgbSfHjhQ8bi
DIiXRaV/8DYG412PYLApRg1qDO2Qjf/j2OxC7LGLUWijYGk+ju9X+JYVCn4MV0pv
U+sqIK9NAVxe89M+ekScXCSv6f0tvmxa1L7NUKkCnR/WHNfgCu+XnXDqMSvLeJRl
ufSiiQCZa6h+XgyNS7+aL5CCQ1zYKBoq4dQhvAnb2Pl6uC7quATbZHeqCVcvmexU
YhiCnntIAw24HyNpb4iFlbTpra2X0kk1M32LVG40BEaXrFYydh6CaD/j6R4t/vBo
75dJ4hazIp5an/5c8OTHf8x6xo8Mv1VsxhBnDm7l+RgmMOEVbEmgElP46QR/4JNa
5cJa1nAj/FvMOmenFVxDH6rVcuFDwly4KLZbNDkBqshl0ZMNy16+nK/LuWtNj+pF
wT8KGujVlaT0N8DyDfo2kHD8j7t1JE2YTKZfjflT9WnTyJ+w2tgSBZqUl2niXoNF
B2AxYs8hHGzlKJ7ygR/kj/baHFXAutnLKUBR5YkxmfKQknUUHZs5nwRI/zfPOHMI
n0FI4QxIPEKOOMBAAI4DfmKWjZ4NTvTOroWxHppBPPIGVUhi6jSlpe7zfCtu/ldz
b8hZUWwXI4HIeg4u7BWPNcZi3LtHYWnGQJmo2oeLb2XZKNYsmbDc8pUqqqqYUt+a
IAYZlh0Zds0V236JLNBBmVDHhUOYbolEI8grYUSt7oMhLLpEe67h+HzKUz/jqv+Z
3M54e0NJTXUBw+jaH2t1k69s/DghDSd6rQ1QwKcS15qpzIxG83cPBmgrWvVcJHYd
bQrw+kEBKzyo8Z7P1qJ3cJHWYi95BIyHG6RE7drtA6Bkz/hi4jF6pNzgeeqEEyI5
oCv3wdtnR7ZcC8JuT1NVvEqXS2Ty0Ahpi5LqudLbF1qDgzOj6NbVRJJLQGXUyxQr
7Om7glca+djyFnWivUgd8t1GxXBjncIfs4uVrovc+AP1vSMjwZXHy0JSlivFoRfP
U2zsKLU0UUaNWqg1QFm9ksYrVIXQp37eRhF8CclsQUv/rzXvVe3Or6HDLYM7iTbI
2UuVlQscFtMueXkhHyhpQwBetMxxGYlM3m6An8e2ANjonyPTP9HevGlxJHMgapr+
NwxATBor8HQ3cFOjgUYI2LcH0fjQG57Azlvp6X7CcKmU+oKxhfts0FM/U526kAlE
5o3luvq5CdXmFegUhtj4iSKqq+j+MTdwNO6O+1+4qsS8CE3f6GWr+Nni8Wgb3/X4
nnUHjhcbLd7OZsON3FcGAgryx9XYCvcKn2R4N7absAm/Pd4OXq8naC3p3iZkVm8u
9Uvht+c0PWYXXBW0pk7mQ4fsdQqeq/rRzvnGHhk6sc9Qlrvr7XLOA5IzumJdFKRV
5Vqm4ZRtBNxrQpDRWFZX0cfdPrzeBInFc8j6QVYs/2jav/lyMRQ0HfLpIL3MUfh+
T8Y7qYHlPXJwxx7OZaSFUotm2GJFmND4xxzCt92guMuhr8N992DUZiLfm/jzzOrT
2SMGI/TL4MwbeE42VK9/jsa+qkwDsQeFrcH00dP9VeNO0KXYwlGS3QKOuNFAmHbU
xmGxfttVjjEZnnymnoLLiMIMF6R+PzjKURZy9A+J4vEMmW+BZXKLEHznL6JMXHye
PzbRFjVeN+GENzmD+m14fmHIpcSDpwpL1Yi18kiH4m13Ac8oKxGlJxC4CWVHWHNA
ft8/OHtPer8QW80a4XUcxUCqALMaiNzATM8EOnDz/INZNBFh4x2f56hE1xcFzwYz
+FPplj40AJ/qTz6iv9s6kRmPhTEaNoCWYwK3SIFR3V7OkO6qYaUQGsuV3jXL5HkN
sGDJ+bf9St28f+d4lFgXXs5mmulC0A6xVzqNKNNAdfkJBYaoig7sWIC960KhItVn
gH5SiBDgE7FqYMWmfU8Upu4fdwTo6+9f5FuZVJwPmzZZaBtuRS6x5vjhrQDrwFQl
KMLNoqaHf1/bLSmQOEEDplxUGk4xEQ5KD+oHh5oR94RNoLDf/M+g5lN989w9Q1cd
t7eRNP4A0Vn4kt7LVJfEsrCObYaQe1BMnkr1NHQZhYi+pqvGjRhJlnsPF4AYCpZ3
P/3NdDtAyH6av7haoMzu66/wAZY/b2K68PP+psVtos/A3MYdYTL290py5j7vi8/v
H/H7Cet7QGK/9Wckj7QU2uAbb2PXfWutMp/iDYaKpDA9FAyGWHH8DMrjNwRQnI5e
scz24o60toMmEhKrng/bl/Mqj/873OjIyqJ9JfBjWBkhMQ3TiKLVIxbl/sp9draR
To1Q4SizpjDLr0JfdJqzh5VuQBM0i5cS/eT/e6vF/1mmD3gkvthUEPg1CTK7HSyV
kALnLLatOcAKBjm9Qdc5VuXLhS4q1m4XUqeAUb/7MDLFVx+D9VfI/bqC5g33Yr0+
fFWmu2/d20nJsbdNNzFPF0gpv3fu2QIz2Wly4eeEk83rzp/WtzYbMdctar1YkThk
ytQZpGluU9zMGIQACtlZc4RwTehNG2vjWqNP9xGwa+Cvq1XDnDtWkqpOjp9I3pl9
hoUmNCXJ3ti5UB7FXVw646nN4GDPxZaDOCUhR28TX9HmfyvUJj0TLq0Zu245VvhD
ji4GeqK2UqQ0loUl/whV/6qCKK7g0YY8tkjwFF/8IDjKLwahiYxoEmysfGNZ+QXz
/ELTaK43YHpVu6qSKaa7H/MD/07fh3H7/yTUJKZg3FXkU6/ECDtt91oNon1SLO9T
eVlCBwx4Ao4LuHfGEjDsr6qzFuwjv4SNczyl7xbOIO+/KKZSwaDrvELWObqCzqCH
IKgkNRUVXg8pL83v+6whFDqMivDB6obNkvdNQFu42mCyiGA8o+rKqJolLeNuJ29O
Fzs/O/KxmNN2V8Oc4EdFhgWjR0fR7hdAgja7XLbrOkrQu2o7p3R7t3liX9+N0Wk6
hDgbORZg33OjSOXgDliTWG+vYpcmH0b66YsbZYXxicAt0buLTteA4blXewj93xMw
xmdIbJnGZulLCVIDGv8ITpXDzOtvPJGWftaB1tIAesH2jOtUXcCW9Cz49Dc2nEID
OnrEWAJOn5ZhzMG0gPW70Y+oFwZ/cMLMOc3ghTGliexnH+TvY5HdIomZ0jQWEUh9
fMtfPg8IFZ0aW5HniTmLflKzwXJ+1d4hKUxwXL1LEcKfLRRXl9PLPyQfkfYD2cL/
59LWiCyKiatN0bjY7H3U1XHhH9dksvU8mu8KAgmXRjIQhnKvjrALGCxR7MEwuYki
HhQTvTzkqxpaBUyZYUbGUU/Fce1RbhEPG3rUq5PqXbaIbV7waZM6k57cvsgp4u/u
Bs9NwPd0/CJ9A/X1xFpwJ4gAFzvgkPdpV4ldnrfciIszQIDCZZxi7bSUb7TveNlR
aR1HRT26d1HT1AvuyKEV2vDBq41T9/c+0SG4qC9ilioBqFoDE1jK+CHWs7YDYcCk
5ODeCnvL9QcQEMXsFW9788MKfnWFWhUKR1xpBxTvSynd69bYydpknqyVbU7OJzjN
viP5UuxxAb9l29p4VpipIWz4tZ8qOXGKwLacu3BzicppOHq/jTjIMvjp/5Wq5hS9
UGRg26TR7pQQC9iz7VFppBncWq0Simf/7hGNl+U3Fyz4AjBQJEoRQZyGg2LmK0YD
I5Q7BV6j6XkrXBBd9Lw0XbRX5U5D1EMdS6K6oRkE6LuzK77FdJdox78zQ64BrmeC
fSk4s3BHTpIabBKEliVklAJNN5p2uUdEWPEOQIAaxdeBn52P8WppY4+n79scumhL
/+rr9n0U1QrH3ZsaPUyXmGyfqX2MkdEf18uFrFjExVlhgYrcVjyPWS++HBgDIsuO
rsKXs67bNvttTl195YtsDpWbnu0yEhDNdliSwVxEAssZOSKPAIo/sc+R+g40mcvI
98lgXfH9UVdnw8yvFpUzNoWMbrwN8eNrkakKh4lTjibtyB1he+zmRc0SEOuQy9Un
yqxjm8KaCppL7KC8bhJ8RXKOh45exr4AjCnXQyGp4uIniwyPn3he2U3AuJa2zCrj
HNhCp8l1ds75F6Zi88yXNGudx9JU+2WlqkbhMNTRBaHWAt4NotnWo4NFjM2H4DCW
OPu0JgKMupbcCiOVIcIpsghcFus5S/DK0wLwvv0dywmhPPp9DW/WrSNP0Ow9miDc
YZ7V1LI9VLCKy8zNFHhvPQ6qnK1tl5tHb7YSqBuuOjaDLxlJ+9tRqnV3IRPVcz0d
Y4ioOL+SbIc2PbrXUAw4gU/jKqa8Bfzu9yZDQAVXJYw+y4Wc/Rv9PDNvFlimdlsJ
n7xBFhURk/CDIm9vGG4HtQVmfUBUkvCGESpZUkLmvr/8psw/ZcnRjAGus6mSuqwU
35xIA43wfr73m86hNK+l/YH1pw8d0KJutk34OfBYY5+mJDlL7Ny+U12gN1eyZzPv
hMoW5RgdZQ9OL2zVvmohmV0xbPaqYqG1kV0T0ne7pvbDx0ktsYmtEeaLs+WWk1tO
Il2QF43AMv+a/YU+hNgaDwxE8zD5CdJEMUG8rtLpxfBw5oyiJYOayHaaPc6jY3bb
KopcaO1HwFTjITExEgCfHfDH8RerkCK8T6tJRK7s+gyaZT43hzBEAd79HH6oxgmU
qGF/lnKJ6bs35uYbl20w4Dv7TiXI7Zsx4S+YVP9nYp0QZfY9q16a0yqXBl9PKCiz
MjntGNBH49p+yKZhwmQKMic3sl/I3DRkRm9PW9X3hffBHjWn9jyEUP6eJ+GiQAMs
2QefqVAx/kIbdxQwn9a2YFc+y418IZP1I2TGy4R9Gd/JmGxEw2syIdZitkXIs1hl
FVYA2DK5H7PuuAQZqmNb9eeqbsfw8Dy/OCp2kmYGcD9lfMUDHszOAiXs7SM6S319
nxuXWFfX9Q1ntZa+gQChgqulmZ+qqRLE1a0iqWtz1Pdp3OIZ4FcGrM+eayJvVNhe
1IkLIVShQINqXpcY3IeXIelM+QrtIyAuiyh90IRpbPUVE825pk5SOMpoekmuF17o
rsTJttZU3gy/H063lweg39oiWFeLc/Rg7RThomqaEm0KZ5uUdfEf4NiNKH8hLdEU
e1EoLBRDcRE1HIPDNRH6yWytSt2jT0BIiByzsC1S98vekblyJ5s4yvutPQc8NoIm
bUWXHiStZW/jzHI/aZXS+mr13sCIlFosUWmgA6qP36x76CMiAnIAyl149iO41TEm
dvrfMVE30byvF8BBTo1H6tsgldxlRP3VsIKnH+0KlrH1llSrHIliVhG8918VGCsH
uuNEKVT/R9kG6LE+eTWwAzG3TufeWOG56wclhkC+yKZTxO3YL02X8oHXwmyMDbdc
BYUsYSftoIx1CsQMXw5/a3u7qMXJEiivDcsNB9L2csLr5L4O2JFraVuNmcOA6j+a
BQpnxTbFuGFHHFBJybkhdJJvwLDzsYu2PXnLdEZIFMFjJFCmhv6MAip5ESVqWhuS
kycnarXgwaQQJxiDVtlnpVqmws7tO7QD1zIkW3ZJZt+IuPK8UK88rm+3GI8Sfkt2
SrGOk0BNGQYCc56ESKpMfTNsvzV5fJOv8zvLILMnoAauq68O4S6YcV67rEMUPnly
wM+Qxj2FvYTT8ChvkKeiulCnOukgNYPZuDjWnFwmRgBiHMpKyDNPj1EJseyrI3G/
QFvyEM8XtEon4oRW/VsPN+qw6ITcFNF06Fo1dputizlKeLMsPcTcxP1NS6RRcas6
NvXDji60HtPqEUlXrGQb1RWhB5chGS1iWRaT/9FQXv3HUMCfyYGBTHbpwzadD5TY
uT7A3yq5AgiMR5fsplOIoQzUed2FyKyFXB+HvGjyCCZWk6vvk3mfp6v5JVJIowhe
3JkhOb091nY3KWwXlW37HuR5SbgAw6cBaBz2ixjyBIrtYZL0KyLWm5XAdCZJ36wQ
rSyQ8np9EEsEj/Ehjryn3B5hu4TTuuV/vCdP1WMfoFURWMBHwikgeBip5cUAXFsy
HEYJVuWe+efOwnOXzNN2S+h4YIFV9A/Xf1dGuskl3QuCdMCzVHnZxNLwadwq9wFI
O4AV7XCtbanvqjnuBojqFatuMO3ABxHcNEQR6PI5Ngqk52SZn2b87KB6GrlQqtSa
cLb8/FCdUkfuGXqJ+VxX77Un77F3WhNTrZA1oCHCwrQBAj7SB3/7hfVkSBwknVJL
KheGi3DjNuSf/qPDvA90o6KQRcKi/cRap5lzwm+qN3UlsJNqnX6rUWzq2L6GAags
/gwE131UAsyD7dbhZ4dNpjhdPbJfss/1pqltYNLur0FNabVtuycZFxAU1BNNXsyT
QkWwtsZHmKl2i8p5e/Ox0hsd7DKynR+MD87B38HnAkLYNKHfngNNzSJinXZ7lhf4
YFRh84v1FNmY6x+sXnQJgKenhPbHUsjr1uJk/NhcYXFnndgap+V+uQOWhy8PUh3l
wbwehUcB7TqKsAtwJ+WLzizzsewaaAyLumn4PA3sQxMU5ZPXfW+hiVukGGQyQ9f8
tF9lP2RopaOCGwglHBmYNBQVDmgccvwF5zhrdywYIWhrzBNCaLMxnhk/jjVJnSFd
aELS+gz5ttpK6twHJ2S5zFn3WVF3PwxHXilYF+Lk0yChzviYQ8oH9m1ZweHw4kT2
v2k+PGuve7ZlYlm7LP4k+4oWqTYAo8gsBMYafRTOCaWWHqmFRPSZ3WEl7QJF4zZW
sDi3Ys6c1Y6WXOSldHFlazMW3kjLD0YOktKoL77shmzbRCVLGZfGMhds8R+xe8wH
8WNmktWhQAb2bEXaYR91EexA8YUgRIBKQ4GI2amFV+ydvdqH7RTRP5GxX0RHTpKR
754g1JFC6AcInexyN0RdyhbFYIYqCipjdFQSj1LkZK7XL/VGcYXr3rCaURs+4OPW
YYS4h1Fvux531RhsDJPKP2Ktds3lABTvqGdrQ/gZf6ql4KTzI+H0b+IAhmLcviLQ
I5NDctb2frMbWFkPbozZYX6doDjz3ObYszHZ93WaC6+ZuZL2sgI4YB7576u+KjtU
gHqwKPjYMWAlzNqGAghfjROtl43aM5w92ucOFZ7DtGIup+9VoTi6ZHi6ULSgP6Ut
FPbsdxVcih1GchkA7dMzeIFp5e41nMLnZra4dofK//Z4JLBExUTtfugO1+ljx9eK
PK6W5TzBMiTBi/ja+XqxwaN04TOcz2Ky5O6jYxpAD3Q5CBaC3e37EwQWwRqx4+Xr
Bi9aezkGWqbFHTZGShiOOpMaM0pZSfv1P+PZicI/+j//GGeIf6o6o+PahHs8+JOe
/UNaJ4ccuDbKiXwJQ2XDo611IfniPyQojy0dKuADFvDPRO8kcmaAER1YIH8HXXYU
9uR2CRrJIeBLUVBHEf5raG8Mn71ieOCtmGOlt8y3Kto+nJKsVnDuOoXjChtmEbr2
yKmuqIwkPDHhwMu417tLgHfRtyVUspuo9HV6y+I1eX1fLjM1yhBQK4KUyZDW7FkT
v07G9Zzum6GrnBkx9QM/O896Fb4rq0aHJXQ5f+hIj/b1q/cNSx6W/eWmSkbGoVhr
8Y1R1KsLI15fpaH3Fv5JR0to/m3PbqucGdMO7qm4i6pggSd4ambH8heR70q4atlT
hCfSpM67+CPE2IJ9IkMK4FQuedwijK5HRv4V691K8KIfZikDczhdNL4Pe0hc915q
C2LEWl3ai+sTUal0onNikRbYLB5AiKS+h5hEYastnRwiqzG9j7vvcoXlIZhL7OZn
1EU73vaJUPZsr3N/el8TcxsOrR+UYbjZs99UU86nJtETlsNAWcx4g2PRhVg6+9Lo
Sk50gVUoVz+Ng0S17U/6+qMre0CyRUrgDSDvK07y+NxPuU0g2J3DR3My1yW0fuLe
tqBwfzlVP2LfZUZzFijJH8mRoYM/T1oC2lhHtaxtlcEseR3+BX7cnwfwxJKe7QkJ
TuY4YdjJcaboDJsgcmTW5LI0orgfKH9AMmHqfve16trH0h3oB0qzJtNma6zUM6dw
cosA+IAGsXDcWi2XRQa8jZscnG/g4uGHwtePoMxIWdwNKqImvvaJi80qQAq6UO4Y
REfMv7PwnreEFn8knA4grFf+ixTFL+hmCcNLuc2gv/yHsRtBLHq9ZaCr9nJsY7Db
lhxDSUm/+kN1dNFUyDIAW2O+7PcWGjF7cJuKlhO3GkI4Bknr1QZnrTSk6e2MthOI
qQmm6FOnqgeAqPWTmPwalvgyjDhEEopr6EYzZaSBlIU21hYKaer0zS4HSBkm0+7T
t3HU9IfAJcazOlYkf0piMVK+l/fi3SJpiemQP1pRgvfMJO7bx9uaKAiW1Uh/eOW9
mcwrBMS1hzql5x3CU6YqUT/PSygSf73RKm9ax4d1j7pSmCST1Du8ISz+KBAjR7Wo
Ae8ySIuqx8OO/ahSRYsrsQTmWcYh4jtaSyY+DT5wGPaDHlF2wxd1QqQoW4mEutTD
+TBGe536aQ+kXgMaWXTDKMnTrEgAP1JxMbq+LakSZQV8+g11Qo/Edx/PZIV6mP8f
4nB9kRaKcl84YVCOv0iV88/qNPoxz/imj+X3u57hPO9niRzdHx608m2hKGSs98XO
eM4q+HaFe0X9YL7CUmAQHflg0+ADasLGb8a/BvtBMh+Sl+ad7PncNZQzhZsDYTqg
e3HZtH5nzowi1epPz3lahfQ7Yxpm44Rc2t5JXN9Gy3Caa/zEPsS1Wmxl8vZCRIqD
2lLK8JnJTf1QLXAFh95SKgHw1dYH3JtzOLux2qyjooSXwwgKFk5lfU35MncJHV/+
Xtdg8Zx90MvOvksghlU0raF+NGezpszqCHH6jXMXzAnileW16meW9Y8vZtD4TOR7
aBDrvUsLQ1MG3EO9Da0D/B++g6wvIZkMaBu1S79U90zAhwnIDvcbjK8/aeqn7sKJ
uqeSXQiTHZ7LQU/hqg0PyC5ghg3efPq6A7ZRkrjYvTDRkAyqePi9JAQZisfBBgAw
YcmQcJqdjU/rGTYI7xmB+1x7Q2pA3FruOfOjQg0FH+/JBY3fGkG8YtACGmk0dg+o
KHMcR8n4/xI0Cdd725oAV6ytHbYTPkfOCEEWr5DgzO3TtupmyUCP4Xs4f113nY0B
pc9OkIHk5DkK8Q2oYajqrtl4Ft/l7SAaV0aN0khbCDGMS+vfXA3HmiNEh4v4wWyO
ctzk5PiXAmfjxKSpY1dKmSN4+l2GVDXiMxQkY94HlK6AiINOWr5eE3Z+kCKk8ktP
nNvw0XLTskaG3fdOG21GDQZvt9ZynRHD38kUrBgkFJOOWrl+r5GhjIOO5i4R4vVI
MfIluEMjk4zDBDTMM+kXWDzE0g8FXoIcL2D+ejETDnRnZKOiHorucR24e/iUI5eF
l4jl0PuARJzysvcscCHw4sPiOln8hB6YXLwI+vrKPbIeBB0yXM+1e39EZXagX01f
iN98gEmWvWGJdrZBPJrxtfZuQRyebEWSxvOUnc1jxl3SCZ5HTo5ZyjyeBiV2JMTx
zqJ9Z+xGZQJrZWt2QA6X1i+ADWi9yz0/bW8SzZFxRCMwjt83pnHqlrN4y2mFXWxb
X3SNT9wKdVyr2xhAPPgJCm62JStt7CrkqvNwRydKPRo+HaX3UdRfgNPoOaBp9EPj
CfWS1TZrEWDenQllXc9sTiXvhHQGLS73vXEUyNNbwUy1t7SOB0X0egtntgRlYpjI
YawT3o6IJUuspqHi8iGtSDslmnkXQzClcgGraTio3MeF9R949xxgN5OLHLElczQ4
BpOIzQhEyTWhpDZH8Kn67sjPSlkWiGy5XAPUCWGOU9a/EDWyaQFVYiH0TiGiZmJO
0QjZKURxvetJepyLeu1W2Wiq//qqEt3Y1GlyO/DX7hASLIP4Vw38A6f788DcVjcX
2MxgVOqT6kYPHA2NySL9IQLydl7EESZo5ZNgA5TDAsSB8PwTn8818X4Jpo1dx0Gr
BDfY0j86k8JSu3iLH8gjK0lplyLk+WO1BlwsArmgw5LYlA3SMF+fGEJAhJTJkHG2
Hj0OmVZXZ4aAR2G93QhTzchgZ5hCL68c8EkQAK6gZU1pgGNkyg0A3r6F438AQMYc
WEjtIZdIn2TyOMit03AMTtkr2AXTJ0c3/ZLhdc/P2YIkE9xbhSgiUrIAPJ57dzyp
myl/1NbMWnNB1IpD/wFXwHmSlqS+XZzDMQbgDNasSfkszV+lBYOR2UbXzTxu9auM
Va9/YDzvoiPwCGjtrNHvbLn15uJf2FYoGhfQPp7IPt86JkjxIz6wX9U21mbZ6lEF
DSWMM7KJdPxFtOB6156Tt7rqfdRY0fQmRCtGFlyKNRRpvuOa44yRuachsE7FCsWu
SNYllifNbIdxK1HVql0EWnmI5HVpUXcZTdve5KkF2eA6Z2VLriB8dUBf9rnhjbN9
TexGRdIr9A5ifS+PCklEpJH4eB6GT6BTOsCeAWmujl0BKzwaFbbtTC+QjtJfRIB0
rYOBUY5WVVzwKRkbjhMvH3YSBs+zYg0ooz9GPNITS3U=
`protect END_PROTECTED
