`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZG3GLtmuEPQFnCEfsPgs3rXH9J0g/nNi/f2txs3nCXUhg5ZC3LtKMs7JMKDUzs2u
UI/sIq2vR1uOE/IzjUci0MAnS6TBGL6Dnz1WSYTdcrR/r7r1EQmwHln97QUuiJcZ
uMb5/UgmWWyk8TFf6gsNhhcl9xShNkPgtEGcu5cxDINmJZYT7Bpp0T+ob0NXgwiU
V09pWesMxI4j8QlWkIE026agsOdP8aSqe3GbCsFwqkmUy7pe2gcs7eC3em9oHYQc
H7WIA1LeO9xtLfcMJnFFi+fjj2H52kx4erEjhtNCuLh+RPmpRJ02XslgALG56a9w
CzMeDLXNm9u7lz5a0HA0pbY6SCvvuGdlck3deqi50ju+VVa2UEabHsGwhhXHTRKu
ToJeJwwaJPllNPc+WQjk7yO53yMod8zt2WzINuAqLuSGzbcRjNfcYuxClxjigJfR
L3hRkF2pYVyoTfYegSFeFtQ7jkBHONfm1Fs2+odUbkBKaZZ5yydnI9V3fWWpuUcT
aG9ZnD0AqyjRVSiSoL/Wmw==
`protect END_PROTECTED
