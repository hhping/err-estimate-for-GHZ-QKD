`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ir5Lz6o2eXLMLdzt3dxb+Lp489hW7J/L7yzwIG6TKfjZ7pBYWF7T7ovyoMtUPbhf
GVG6ipuDPyrq6bCH1Lw6JQVhqJ4zKIHFVrtWEOiCMVKPPuSGFwCY30pKa8MhZtLb
1lhdhEUxKcE9L+RSiQCBfN6OxjMn66QxdaOc6B4pDrFC5CEDgw7xDA+8+hO4ttBz
Nm9hkY5iJg4twZTkJauFA9wG55bRW0yWke1KufSWISa/goRzYOGKv6r7L9g/VOLH
ltSZ983XGzPY7O7cg0Bs+XPPrh/ONc25dldNwe1BjWx8S/KLlaWE2KHOsEcqnrUG
LddFX2XDuepB9raxWDBBLi9EMJcavAZC3yvUP5XhPsH8NQYYOZnGgs8kGdtTnOYC
hGyca81VEZt+4iU1rOn4MjkuFbCa1EaTzDHP9Hk20i5Izob5/i7jAPemn9pfBFwy
476HV1SttWQHIczoEcyoyh8Zk+Ra2Z4pyizQwVOJVqE3ndZEdjScA1xP40fkPRnL
2Xc6/51HRduYahVF3RxmyW+0jrwRVlF2H7wbl1jOlzG8i3LoB7vztK5FGzGFrdTZ
OGrOlPzLj+WmpkYe/0kT6KCmRjpHBXpZ0c8KYe9sfEg3ykzH/OTVB2DaCliRmM9n
xt9on7uS+MihQZRBovzScNYda20576yHKVOtG/19e6NBwymQJbvRE2eJ+QrDBS/t
L9sasPTMnnQhoOaXVYl1eZapSTRLaHJFG7KnFVck9fbA4WvuqAu6bVmIF3BFWw2H
FSIGyJD01xBYlhD6F6six7zEEBdwQjOf6J/avR25dQdMONacOw4I9TVa2ITlto4A
km5NTvO4wbuhtDuf5CXgElQnG9ylnjiidpn6HxF+ZFZ7QZpGtshfo4YlN+VTYKJ+
OhGBfMiRWfWHHsj1Waq9HNnt7ieBmbRapBRqtH4JrFtYN1W+el67flWEnXcXUPoR
oqFXJ53V62vfxkQcAkpgC/vHBLTGe0j7Aqd8N3tf5O7KOf5XuyRfmW1Lz4MEtcRz
F0JCh86h2xyN8zBSSfO7hrQO98sMvtt+rOfREqxHMNtn0lAXgAaaXEjcuKpdYpIf
GAXnKKIy6no4ERfw/8cn5/+yLvcM7GknL0tY9lKovKjbGVvLq5tZLTWsU410NzRe
k3A2+zrnwWNCuIZERD5W+ZuxZZVF5QseU9P2A4aK7uoiXLMGqqtMP9AvFqUM0/xQ
zBXxwJrVDueCmBG/SIMoP0lpQVAUI597rlhJ75AHoSuzAMIyWiLXQwhKCinMWwWe
Bt5QiR2uXIpTBuQIOY9uOf2pZXAvxV50IZDCHTrRbkdnGhV/44O3fbi871bE/IFI
kVs/cxPByvqJzyZtgisxbRi+oCOvV97Jpx0Ca/3ywl+8RABHH1p2q2LZgann7B/i
dMLPI3GSOU3lQ0jdfqRfCFVbyIMSKr3UPOSfqjAK5B+8Yk6Y+a8fiV1US+C3K2MX
AbrtNYI4fVXyXdXkwr7OP8kuOQSgVFfdZhH5TI4AI6IIZdSx+4xvr3fGIDBlEZvH
/xbnY/AczJ1pyg26jt8BpCQbjBi+E1Pq8ycTfgAu8+qKPT4Hp6i6KwA7oyGPyU9E
dFp6GB5GKvixs7UqjVqK2ZHmAB8oLMeeA2RcktUmNXNu+pNy7+8+eZGIjwXqlQA3
aDD4IDQA9a2rR7HBZmWpSuyprYiOvHiiCHLFlHwy0AfcUhSvYLoF/wG1FIaxLLb2
9nAbqwhaKOpHai/QLVQinCvAKSXgOw7SKIkvPg2XGsc59+/xCRkvz9H0QPOI1cGd
7/+HCg2q/oumhX+YV0x4QAVkkvR1eGYoNe59uWZEQigDtq4HK6GsYQsQdW9gW0qw
ZfSmy5DoQ6a5sUWS3MJ6vZqi+pXTz6NxJPFcbY3doh3POmIRf5MS8lwSsSdGTp4O
8UOxfGtuaM76f24XFmg8f/U/i/CSZLgSDRWON75aJvKTJM9Z+UEjyqM5qObwmTXp
9AYTMZvloaSY0dENUupSAlv5n+dpu/rIE3tQOHbPgaI3jbZ4MNj3YL9B3aHhVp1u
9OviSyYjHNli3upB0IHCpE40rM+H3zLHbvpXXO6uQKq0gX5CeObWg/z8CYQCs2Q1
ZeC1JiLYU5WD/JIliVlkxGl/iHWtxb630MQTqKQbANuxgm4DoltDx2ATST+/tbz9
3SGRz5S4+LdG/bgcyIFNJYZRUYm3ib+ZmRW4ag1cyjJ5yNQWABqGab7JNFeYjuED
DQs3UTdx/XzoavCumvjSwb2xwCzagx7xK+YPgn+RrLruuXFFERjVh6WI7ewL8202
AzLdHsNlzxoMNemCRLOO5XajImqF5iUCWF7JjhznojcMDYVBDMvRPsVJxVWQlX2u
XJQGJ3zYsGRYvo9FkNYjxviEzpAXkpSQ7BdH469CgJJyvVpycpQZSOHtGrDSz8D7
IEmcpSQ1ZFo3WpvrSdC+PuKUR0npZXJwiuhGQd9xVMkJIpSESxHdMOjarfbg7c3G
Z5V+taAeFL0Jn6evyae/prGMQTi5Tz7Mp2Xr8PGTsXEqbgCwiVa6eIVjGDedIFuS
HZJlHDetdI9K8/VtHE9IHHImYKWg1dR4Ix17KasiG3yWulb/Q7Ddh7AcEget2AjM
aMpkLvYC3RW3PH7X1VAmgD1cd5HcVoJ3IaWkZts+qoPfeqlEGLDHKgpVicF72KOi
rR4HWL7CiKTkeKRy7/0V2vFeo094s35HGbufW8W/zOWDBdM1GYu/tcQJ8Gx3J62p
/nmLq585k02Dp6iNOTpMLDonYe++Q2vUZRzTnxIZEkGmi9HUaDTjmFEQcE+jKqN+
IhdVrTMztywNwq002mjKI9Z61XckGNz9mW9wCui3wT2EOm5YTvI2zupEtW8FiqDO
B/ssofbABVAX4KB8AOvsM+3O4YbjwkIokAr6oCaZbhsG+2eEDiB+JTvx24oeSmV1
NmGUHJNp5ennGaaJinL7aJ/nGTAX9QhKXm10urUBtIysiPylkxk+2pV9Atg4c/FI
v9EdYv7hetamo2bqwaeaTiM9gsH9mxDC6iijwDhMzUV2q+4FV48nTw7bMWCX/1mp
SC4R1LUWpYCNriN2m14Nsbdy9pVBpVGD6JdVzwbeY2xfGWdVZ8tkXAtQcJO7XQwY
9XIT7zgF75Tv/CoVKoivuAOaAO7QTxVbdY1FQMs3frUFCUkJHX7Sr9bT8zvSlxrr
SiqIdKE0Wt9u6rxXHFst/MaPH7FsKZarFDLkuAWzCofr0XC5Qsc/9tZYWjV8cqxZ
zYzxvasE6g52FmCWNlMUYBHPRSH/VRiTrd1qOeqWHRtFGjjrfy/GxtFuzXrhHALR
39f+AGWJM5uA3IYTD+KSHsT2MYXX0dvhpy6E0czfLulxVGSO1zSRgRY5virQiSC5
cQa73s6X34iTdExmXR/MS1pT+FgSd8WN1sZXe2lfMnUqpMMPBS3LtTGtPLHkciAY
xlnmqccMRM3uaSKXfDxnJHMnXUlsN7hKVc9s1YBmX8RaoEQNFW3xVfOXh99TG8B0
8G32CintKrODCMZnRM102hakxWkqXA2oC2vsRVwfZng8lSurx5ItzoPrrniaXEr+
0V8c9MXFh7Ri0lhAnZ31DONCax9l8OVCyg21ofOvfqfWSEQTbqeByNWmzW50nah9
4zPU1jE+hGfpZe6H/m3XDqVhYJ3kDgVMM1ibkdDJizijhWnllrbVdzNr81Lg7oVE
tCSBAbCW3J+SL4i6Qi+JosqtZTBPmKGd/1HQubMYfP9DmzXJzc6FFJoYM2vvZru1
DABqAbrq6MGLi+0WAqOqCo9/AvalZ3oAjTX5q8oo6Aiq355a2cXf597L1jihdOQE
rFqCmUIjNzGyflXmGUw/ZMFK8tWQ2ZSRG59iE/JBhjLaoiOVk2gME76LxCDhtp5X
uv19n75il1bZ6JhC9tT0aAysA74ZNDxRup+EEGMdsirag/1naZvdZvK7w5cH4vva
/ORZqhQkFKrhlLxGs1+DgSfYlJvuo5Dc3PasL2Qk1ovYyY4ORJeb+gjfNmk6itHb
TIEMTGggU35s2NWfmUDno+EBgl0+E1FMU5ip+XLn7bV8LHLJG4jFqDppeqXNBXvL
Js5qgz04jGJdwrbrGG4v1Map0q8znyPNGhBlpWH3v2NsybUH3bEtEAtq7ZEEEATV
X6Gs7F86VHLuBaF3j7gi1iDtJaiKY8iD17nFmnA+ERBqvMW7gHJZTqLsh86L4eLj
p+sLYE6sA0i0z6by97D9TsTSaCoGwPVwNJ/YDM6+i8JOHm4pBGXbJJblYZn2yyIe
NscmvPG8xn4m+LnNy1OyDlYUHqA0QFKNIQUYEFkIIVnFpmA0ipKtt+42BlRgNzwD
VuaaNEtv43cWMoJ5XtgGT4sBUYsLbJU7BFNehflMewAYJHChPW9YplkH161imWFY
5SKJKEP65XXdr4os6qPoip/B8tPuadW7oqe3e1nZpkA9OTCWaMZGb0GN/rOvZS3W
nhKOBzMbmf8VlYRgqbvndxsc+3W4ZPknt/aKXox/HAPKrTkoipsF/bttlZ1AnPTU
ovMdin34qHBbd3jSBTlnIAHBkhmkU2P1DXfp2Aoa3nz5aUzr/RDGjPaclSCUjMas
fPF9NojR/rNeomateorwnZRt1+r32wDRKaIfTHWNQAClu8aTyJO7a5R9Xxyy4WiQ
xaFhHP8cbAX9t+oONyHhTJSVn5KyUY86YwYfdSmhPAdGV0y5uFh0yM0rb20N+NhT
zbaesFNPofSOyHeZQ9sNWcjOYLLqUW96HKgsDirtZ+2KGdnUYMQ7E3DAfvhelZAc
ygHYc9nRgk9Bp0uTRZEKF4N41+yfrysSOjCo3nE4yYNhPW7x4DQDaSCXdbkCISQx
uFp1bsaNwATQ0oD7YD8Xu4Kvm3t1sXmi/Vo5c1gEQXU29lCANiBym7OHDPUFfwvB
3g2nQmact9AZjuC/hlYMa0SVwAMkLL4xkwxf8rXj+nGaxvLecDFDEBiO+Rh6gmi/
/H2Jrk9BNfC9B0xS5SN80xTcQUrpi60GtYCjIGkeTTQ+hqeWb/+jMDGMsZuFvWNw
ZPDxCnUDq+26rSTv6vxav9mtjVvxOKnmhNp2r1KlxCJeitjnecdFxAfs74TEgT8O
M8FnZHIfsaIXkE0dD1mH+RtRMr24rPPG0iomlCh665FdjH+q9xBbUtOO9Dorr0/4
TeqSUrAodp9oyhQg4yWQ6X1NiAbKtjT2wQrEEfbSlb4+fzZ7mW8lnUOi6rzKCW52
bz3ebXomrqSNbhKTFmO7HlBhs9FbV5/oMxseP6kOc4U3+bqkW4I020H/Qoteb7lp
3O+l8slgz+/WvXz87rtxav0qluTKXcJIiHZpbqtUSpHuCh1LAM5uFJbI4bJw457R
ol+acafTrUhZp6p2QVXoFjpCb4cfmYhZNgli7djUxbJqxhzepQ/f5opcp4ZBSt6Y
QViUQah7Ru9CmIOOPYIA2vQ82ERs2ehzXxkEsG/QDTvB0ANcJcJcQ6UfqZjo4rFw
kcyyM+oP1eg+kFbmpRSCUEyjXsq4Z48ekaw8yg1VSt/G1Wfw7JfmoWfM0w91jiKa
JhqD4wLBbBVvYdPxxX8+SkKfgNRSNAoEYdoTAWJ0/wrw90mgSlkqx3ZAjjpwmX8B
24VhHyU6YfNYbtpvlneMQSw9i4No2MFJj9/pZBWRexVGeNsof/4zsVgZfF0C3U0/
5fwXeEITMedsH42sBlzoUxoBdlo4yxweD20KHvdFLofDhw88tMpquINAeSXoiDMV
wB1vJuiUn4RtIRtsafAkwM03FWpUrmWLa0dzH7O5CE/U1EiY+rGTU4X+YOu7x6Fj
aNoLOM5IGJgjyTHF7J7elsIY1FQDWfhsfruz7xJ4btEbhUgOSkzsmRYiEqvfrPqH
UXxjWbHhpBWj2WBa3ox0esvApuWTBx+CWq/ta0opQb0=
`protect END_PROTECTED
