`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjwWpgipl8JuGMOxP7BJnuibLtYj1wY59+CYIa00VaJk8skuz2DMic/SoZkvnHDm
JAyiyWGXzsWQ+HypVmd+apgLlhFrlWCVuB/IuEZdh1InI4U3ETacEnR9jiBYwgU5
j3HMmCr5h6H76pAjb6vA0H1puDUPKcWLCYG5gy3wwep0GPfAD2b5wEm4wbcr+X1x
yHxeytafhY/1Idqpalqc9HssKCWB3RC8dD9uek1JHrHY8BZP3GP+1F5ADGwtlw7d
`protect END_PROTECTED
