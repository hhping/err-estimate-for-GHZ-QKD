`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PmNFvPNfEEcI557ExKjdznHphGMpIbaBQqqi2FhJkjSDPP3zeBe6Z6LjNVBcUuu2
vHfzzH/4z1DquHpCdTtwQ7chYoo0A9flUKSoJlOfdsw5RZzVFtQ5rI2avQARDVgj
e5rz0nbqdaKBUpiW4iHxpkd+XPa1jgh/aWuT+u8uxkxUYc65oFbp5ffRlDOFBe+c
oUJXZlrjSQA56Sys5Vip/racXLFu3I2YhUFWXcq7jlRFsFtMVUDwqfLWJKxaNGrg
n83DJecoMOtpW0UVOCSzUhiQUoAyD6jAbPTxbyqdkFnEmctkBBtajUhqe/ggcjaj
ufDZT8DmMrOPOsmQs+WEvoFEB10hlVLfsvO9m2gq7p9c741WRW2x3qXla27aScb9
99MYboHfHu1NWsqhkfuaRucO3HFJbTIcnYE/+bgg/ldYiMT5t9sioWqipjMCFm3e
iYyKZfUapchCJMuxEAL4+bpQ8N/KFReZYGCWQQpmmruBmSTmEYCLh1UWQCrNRREE
g8YDCoox1xONUPI9J99jt3K7P5MN5qhEkskoXuzMOA50dcLkH/YmbFfRTgsfjdqZ
cerJkhVE3URQRlMI2Hj1x7sKkAAwr3g8jhQn+jtFSB8mlLSq0FYd18Sf+O1PFnD0
uJdMbom2KAS77B55l6xC3QoMw3rcnR5dw58npqOVWCgDJpVDrhBGMsynjKvRS69b
ddajtMakGcHVDQXfhalVvBuWFigP3yPJnyxbPDb6DIaEEq6nH4BOz/WGZv7NZeTj
nmZQ66qQfwekHSMvuiy8FZHqnOBNzN6DVUFZ2x1js0X87sUIBLCy6G4ELb8KJ33D
qVaNi1H9kqD0uL99MQS+WYlFxU1m//yG1M6OmtWJf+/divCIExwkOwqXMrD1zZ3j
2JdFyNvGyxlURCILxSI6Sub3W1bMAKtuRsBfMUeAAF0TG2Pldv+K5Cxhw1whC861
q0ucw3XbKiAfNf+fe9PIsBSH0To2Jj++0yzf2OzyS6ylKl/F6LHudaDNA0uPgle1
FwTZJ/eVUiPdiHBO70izRonO+PvPGtjNEvAfkaS3mAL+FzyMkODIhe/A5w8iagBN
XbyS+0zWQZ38ATvpWp6Rpx6vdZb/vWLtESz0GvRAE7U/31sKK+fu1uV7yP6JzXxP
Fo+eZAxkjMekcfDyuqtridYS7WGf2AFH+OaAMb7arKuIkm8p8pzfAtYqVbuqjo5e
8JvZps6+HvGWDrdadHQ89r6Iz7X5A3AFjQbG6WTvYYrykMoYYwCHJCbRreYOQuWj
vAtNF+7o9VXVmNG3wHIz3q2bSRbLnb45LVfzUOBxz1WVOcLbo7vL3Zc1Ubh05uhH
HgUFYW8Sekw6y0fck724oPEk7/UGsXYIj63aA6kohPT8TMNlXNLasYBuzKv4FaJJ
Yfh7ktbUCgOJm5KpSYOZwsJVouNqlilXbAhqHS07mNQqqChplfpR1Kb6EZnBd5mW
EA2b1qiBNZNYMNP3t9nAruFCp79qjdnSX/wqYQaM7um4kW7e9K+orc5mbGS3iP6W
n+XXKZEes+iImbNV1wc+LNikercIfSocN9uWhL/F/gqlPuaRMjsRVDEDgY8z84uV
81LYQayufdxuEgU2fx4q8ihrOpW5DHIvM3mu5RHg8DcvNeYGDKWD77zd+e2xwRzK
HxjCJBcZlC2Z8yNWdJwRaMC/LoQDKMva1PB7MjbGn1ZW2e/qIpiJiw/Tuthzeg0L
CjBod2aLBGG+kUIu48tCSLzdn/b+MbEmKtoSFO8zXzg7oDunW5AbF4BRtHHDeyBg
prJGL3Md2p2a13LbOssaO2LG7TDnCovjub1P/bkkNo/rhTJrBqGb8KX7qZoAs0CM
Wwh3Cgxz1Xpy1pk8qbMA6A==
`protect END_PROTECTED
