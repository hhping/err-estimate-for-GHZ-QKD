`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zc62FyjCmSHstbIKtUuhQ7r2NqFFCoJGDg01B3tEeWC4UvjqupjRwkpeInlh2VJq
GECcx1GgmLLQcyTl7S6D2cftRykTGwMjdSbeF9HaKkI3E1t+4LNSnCXC1vW1sUWA
sl/IgX2vjTPzHYHlzRMWy1Pd49wdAJlL1oILDKfVYGp3DJDbHWZzCQVHnZYpF0jM
5Z5Zx8L7Jh2/FbCCr+obaNHIxnIi+/iibnMQad6AEufzG6ZN2i9/n94KWaYIcQKR
SapDQVpY8vVqTkmBdtUyQ2Mr+9dk0iw8bMn6O/LCItBA8JIlHWVX5BKzlkuKgiKL
MGnMWSWCNiCbDpfRkAWI5Ws4Bchgg9ZF0OOBrZJLySk40G2wGxlCn7e11F1wP1gv
vz/wRIOLqgr7TwgTKOZNV+4Gc8cZmpHP9B6uBk2Hwgt/AqMlQdx+MjSV+COQOD/i
8kw+j7Bax8hbfzeP5CsW23/+9CvSHSRLxDKRl5UXSuA0vyALolHv5F6onMN1z4tM
wDt4lidpp5xjl5TJB0DakcYUqYACm93+OqmpoLeKkri8oaqEp/DpcrYeqegVC3p0
JOs+ogi/oGrxw0dif1OHH3FRkEBgF7GHN4fwwFDjobbGOgRpxY6vHEXK4OQlqutG
zWLwWknpLFRFiU8MkeSfroAlqmsELpYWyygOU1RhukXWa31ZDgr9caV01BdQy29u
s2Z0+gOSUchu3Ggmlb8LcnSfd53DbeEG2lmgGXQgFCw/WdUQC3AQOZqZmzl/Ao1b
fIrbI5ECDtEAFV1lW54CVDBUrjlb+5YImNXEnXhCMdQmOCSGrMPC+93LWzJ5dmHG
4T6yf4WfQg1nEoOu/vijKjaSo8f2+YwSrcvzs49Wkv3QTZreCIqzv+EyvUUkbB66
yZsMkQ7FEeBm/fbGgODr3qG1uHI5Zs0Tfm4W0wgd7M1fBqL03jWuiTuIw3Cc2XhI
wTfTMiGEsElA3C3qviU35i2IlzWBnHxr7VIeL6N2MkI=
`protect END_PROTECTED
