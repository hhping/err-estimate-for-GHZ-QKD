`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvLjCOkhKlLZ/QqNzNJY4Y575ZNPGoluchT9BbB6M+IJF2ULUvQ7ESIbrou8sW+G
QKRPxEaL71ELDRFCss6FIp08a0B1FHmRwvQJ3ihf35zW9WcHkmVFKASLArJx0YCQ
2WxjQzhGnJ1cVaF7bgg3nTLsJ1kFg9ASpaH6kr4lrl6ULDXCAu7ysv2nWOCUATbw
odYu1H2bRGqHHE8YTRy+EtI3psjNvKrciCPBA6dlIasgo0mgMauwTuw/SYj+B9Gc
d7CfcpBf+U4cyKPzpGUyXE39IxZMxjnMrXAMQYQPZRjPBfDLOd2nS8FjY+vgDrbx
90KQ26cdMqzXhuVkHMCnAsCnq8+aWhtUdmD2u6QL9OWMHMlbOXGBwBwI0zf8xM65
k8/U77pcL2ljy0ElzI/sApvPTSKpXekGPUlFfmZTE2fP/OSU49ocJWxNdzf8qIqS
OOiU+kuNahnEv9HgjMezoN8RG14TaRuLxOAqMa/CVfC4Fji3+0jcY4ohSA/o+ypt
FkIK75blMts0l4WXUZlYBUMFNSBbtEJhVgAJSC3HfE90z+HKPSizBajY48c8noJo
sOfT39oS58HdLkvdW+e1h4QnLujtIxUM4OR/Q/ckosy0LkFtzb/R85RZq8mjtl0U
EQQ2wUqL6WLy2gck/1HN7LJrGWIaWNecO/lyYFc/Bk5dSSDj5Pit6qqyB6Y2kJ9H
faILrkIBSZg7iVp/kUA9iDMRnD4LpxI/fAOBUaM9Fh6MmfPeD4vTbdbO8WNSUQH+
oUw2wsZvk/ohaPLkL0BNSja0kolZmlm+F0J/SZ6Dh1RWIAYsWZdVdF6/BdrSArEk
ZGCqtgG48YwloRgnIKrssg==
`protect END_PROTECTED
