`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SuUyZDJj3aDpZQmhCbGNwY/Rt6DQCyU7AwTrzRvE4aET0nqP+igKch1jK5/9U1UK
G3+hp2WfdTsuy2tpC6h+/QhyFXHTdNGvGDGSRHyjVvNtA+otYfXxWGpZ0wMaouKJ
O153Bp8k+p1H3qvHicSZdigrNe6CiEBri+vu8w+SbFK2Dp23De5hxda/e8XKGVlu
m+jIAxXQ8/IorqhvgxAeMDQpYA+wf0SdHOlj9X0PSbpqMJNMM4uEFe5l3MrrxRvx
RAss/BtnPXF9mujbPUfMgwBUQnrDlbZQLEOWib+RV6g=
`protect END_PROTECTED
