`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZsA4dpnIK1W7SezMwYDI8iYkmgSoWLNYReCh7uUekbn/Jy9dEgA9IiSJTxAZ0RK
VC5Xd9/N/IOefRKn/h0rjHi0jVa+MUPGda8zEHrhYBzTkbdU2vwY6JhwGtmNhLZm
0WtoNSgGXUMaPSjo+1DzVZ+gUFstwVsAkZTIwrC0tvLA2V/4Jtd107j++8Ag5Fmf
YFFgxPrfU/DBeGH99KeNJAWcmq2P+JM2tgKUd5ZTCKY4OMc4x9BJS+FxB2B+t3oS
TvH8vSMVmXoYh8yvSmqmTE6qac3lXmUvEZf6UO46hYMakYIe6+d0Nu9JmdDW5VNb
h+s1U31W63BKiJ+DaM23rn8qC8yiricodd04vzkhfMN0SCC/tEsS0jc96+SpD7Th
SE/Gb5NEiQYlwAmXGSi1pZha5gORXEttVACrudKXw8A4bSD2L1mHKAwOTJM/Apdp
unO96vLlKEInKtmlY+2QyDBRPu8fc1xIVXXZv0hWW66mfITPGIt1MUiJzJMV8aiA
rDmtZOb08MCh6QPxI6G7RgwDVBBHD8fYfxKsVyx9D8gxkFmc0g0RNiznVdAWhFpd
YlRJB4Hb6fOU2HWunYl/NV9AGUrZ86JebuuzDc0yg+lCndNgJp5MABYiZ4EaxMjP
1Xo1qM+QaeBfdEjCULQ+pnUpeq1vf3PVN9Ppgk3pAAo3z+WSFHq/U7ihWkn1eY6o
6zfn7AEPv/cv6E7J9XxRgCprc8aNte8Ol1R/+vU7ge4mB6pl/PNAVUmN/HTxrAIE
`protect END_PROTECTED
