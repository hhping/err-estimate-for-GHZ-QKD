`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzN6W4frvON2CV1oyBN2l95GRbl4TnCGNJ1mjEm4MLkzn0EmTAz8N4BZ7Gpk4sa1
bHVAikUjg/k80KAlHSTmJra+rmmr4KDvbqoDVnpgAiIX6wVVpYiDEnxjdVNKU6HA
H0A5axCLQ1HZOnOAYMc3NN3Oo7yjWXfM67GmAqjsMC0UewpSWDwcfkS4ac76OyC5
i0WEA1F/dRLCxbP7VYipDF8t6OZBw60qbg/dlkug6bOHYl+fChGCJboFug4nPUnZ
CBJRUfb1tnHPdbVPjg9NPDQy/WYuUgSLe0y7r8B9r2qVcHm097E0Oo+qPV0tq3kp
DV6Ru5lBvEoNnmXR1ukd6r921KGTDOgDodvGEa8H6s2buemHMSnwnKBqF5bAbEoP
Ebe4CRofkM6guCiCymDtIoflaFSf5XCN8pybtFLgIt+AyzVXw9DeOSCfgnyfe0BW
PobYhIgwK+5NkDgMeGjpIRVavbPAkow+FxLCEFmIVz22rR3z5i4Z/eOTSmxxBUC+
qhPsfshMgd5VWIpmpxgss3O3RDzB6+RH55ii/Y/9yMhR6X94o6Y2xuluU82cCeGi
2uf/6m+VfkEshtHDAa9xygAXXJgRXFwhi65VXJpdlAOOXoWD/OeWEWCnoWEb2uAF
xcLepepfxagYsGQjqBOPTz/fBVahcy5IzDFwqDJe3eQ=
`protect END_PROTECTED
