`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cw4qGHEMzOGJby5eijjPifp9MHicaP/rt5l50d+vwK9Q2NBRDprqamoNxUxc0qGG
06pXmT+Hv1LvcJB2f4w5wR2v3bE6GJh4CSj7PWpPNTIsT6IoBSAbvQtKOLv49sXq
Qb3UeT+Tsqu+WUH6Yq1IGMIAaHGlVD2S1XIOfvi8Y9kBL+KqIGebYpx8gNgtG8JK
QiTo1eC4MpiL3Xk4kyESgrVsydUKygIjUJFsAxgI5aBah/aLEUlqaKLraaBOn/zX
bZDZHB4X+AvHjibR7pJ/Bj7qQH6zgPGrClPxlPh6fTcbZuC2HWzzVxkEx6L6vT90
4nc00IkmDqTDHMDnVicKY9i5wGmSlcIFBxEkRFS0WNIXJOPieSjVQXVLmohSc83M
mWKqKwq6k4yk6R3vb8nnfVZtNRNKQ4uSQ2fTl1bl7FONNMSIB0S/vvJL1aoUg9M2
ZyV2wFLV5U6RSUIDJiUdM8KPy9DQAehtY9dOW3nI7Y2a3ddqtdcnky/FTw7PJpMS
i/meUhaw1pSTfNSlRssjusqMyIZ+LG+rFcD4VU2mP2uVlRteqk19m1t3tb/PL0g2
7JiaxyjCtB6/MXsYZ1YYD9GQVh+XupcW02RgHtWwg4xd6KcTJ+R2xCRPhjEBvhiV
SgF4cfUBMtZ70WaSYg2DWuKspGCPU3ofW6Zm6YDVtgfcoWjNlcgv6bUrHgdzGP2K
Dr8tiQ5zzmxfUT1anALSznFRhqUtS32DB49QhLXpktI=
`protect END_PROTECTED
