`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0j64yJbzjOO1CZJdeWUE7HN/oywZFZNvFMqMo8t0yWmxmy4+qEdgo7U+c6DDsrR
sQNCnYkENDofrATRo0V+JwvwYB/FITxjMrxelV1bYwXIqpaYRfSxpDpkEjVIOKYb
TwBmbLgsXWJuXx1nyzuWSPnEMW/ID7+ix+WbLRCIbtR5xqlwDeFWXJN4HFxe/Mfz
qkw1N2P5hbJshdvXVSMI7soyhbi8kh4M+CUJbQZOKbwVu+qYdKsj5x7qX8bOmfE7
wkwYFss3FXWx67VNC/kSuyGSjFekAZ8NrvuXmuG1NppLH3cvLeAAb6M9AyopTLap
0v3atL4u6BiVkO3+zsX+pDhx09ISsiYTXWkWid651BX/n196w1t8nqnphoqZfq1v
+KFtFX0PA1jN4xm0fY7sU1siAlcpasMa+b8JqJXiHgrrzoPDFswReV/omCzIrfoc
b1Dz6Z6k7u6NuSJsXdfOH+OUWEcNwweFo9D9f76r+EtNduEWIPMOgYHi8wDnTOy7
cvo6dk6AjK7QKFB+DldEGVlSI79zv6udg/lUN6ZI0es0BlNyqUAdAZDmjQdMi4aO
Vf+c9gvzyy4YSZfoWSGisviVuG9mh4QkXshi4xAYaFKEVCH+suEn0CHjtGtTZbiA
2uV3V3xOkFJx8ZrJSk7c8c/g1Qy+/6CbDne77WymjnP/IL7LKhjNZ8FAjtKn50A9
Z4F/FrrFYW64YvIRC8vwQ5iu581yy7i6e4/bCyT83X8GaexzZRyZDqgUmLE0sR1p
7JgPgUyfrY9neiOqxywaDrFbgMMoUlElHric4RVGoYhGl0/T5vbL5aQ3xLEGdZup
Ditr4PCcGIkWjV3a2kunCpTN+Uv17qQZsxmdbdpwX6byZY7WvLXJqINuyrMGU6xs
Xw7vWimn2tA3g3iBAfLgQToRXyrs7A9f/836IJTsMLFBMi7mSQoqvcMv9hu5gJzB
YLKTwVUQks2nYg4mv4Uu4Qqc2iuUsI0MU+Y5RT5M44SU62QP0Tc1ADk/WiiuCuT0
cps8JPo/bq0WI2MiX7KMrfJAvF11HD1FcS/E6aW7R9r9/WtCvmMeqo8nyD7wC20B
`protect END_PROTECTED
