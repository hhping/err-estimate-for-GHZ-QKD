`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXXk3io0aupL+WtR+WT4eH/MNrH6LErc2Z1nDnf39m168K4FAOVHP6gegdX3Xdue
wPhPKQCEW9iVAT9/rnajMHtxxpKYALX0Ez9JFJeUSfUeKi3teMv4/x7nS28R6lh+
dJkk88JmBR08tr+D8CAvnMhofM80FKssiQTyvw//KgXVxRX80nGr6FnOF4V+eJPx
mpe94mD1TXMGE3uFfFbNY5iT20hnfQJLiJfZBYu9J6+s7CWDoCXoLZq+LnvJhilb
Ot+mHf7QG2Foj5VZ1VIzN7X/w/a/eq3MRHJeWKVxO/zVLqcYKD2O0YazCnDguHrt
HiwT50Qg/47uveAkbHExH9XZRo2/OimrgPMmMkIqAXggXvWXDVOn2YP0zBm7SJ+c
QJyFfpHAMcaM5ZaE9y3tUPI9oiHEXcB+I2aXmUGHC31G2l0m7iC/SlS++EUkb4Hr
L0R8KxGL8BdLHeFLs00C1L9/RMM1QywaIQ1YBmp23NCkOCYgb9UiqP6e3/R0Nxg2
vmzDvjAE0zuN/Vai6Er4wZxZJn2/owYPwcXmYir8xF/aIIB0QUH7t+4/93O0rcSM
FtIo+0NzH3+hDTR79bFdnK5t4oAFP81TF6QmExvKzBnz86ty37rSY9N1fwvOQEIE
ipAEjnPogWW3vNUQgVFIy0euqaYwZo470g6U99qQfX/mPuX9akELxsgrNCjQpiVF
xwi2fX3polscGq1nt5XE2nYg/GKzuNqONt4fpNfhn7dHw6FXgFprCnsAHKowbLe3
cYDwOTzKGnlr4R94ZquuEEPAa8o5EjCSGKLMc46XexWxLrhe2WPfXO70AGumC8hl
OkyZ0WBrne5rwO4ZhuXTXQi0IGh0p4jz5XsCfkEM97pGW8OacAqpqPS1YA8QqEfV
3mQGR3UOOcRdlOTqxxuhM+hcG5G742kw/pybQgBi7wXmjpb46q3WDH5Of1RIPB7Z
MZmhgeJwGZxbdrS/zG2rkLqFsGEybV18PWZ641VI7NQDFsQk3LByVrhCJbUiomvl
FBtzml1Jf7nmPVRwbXFXYJ9MQEGN9dSiIQYZPfnpHd0sHjiRdVXK8ZWiwdTpS0jP
eFBYJaf8cahfTZB5oKHku18tcwbMyvqdzxdrV09ivilY5o/+QbFh8miQxEXHcc9i
g1NTeOR10+fhJV0FxiVCEPTy8VvDUeATHe9MZ6fl2qASuhqiLhlmNvWejrahzFiF
0fZPiCXO+HMTpRL8gghWez+QdRzLPCAOGRJET+ZOiMQi9ELQjIJ3NvUG1VD7aByg
N880WzRMyXPg/hs60AGwK4IpY+NwTkZYyo1oTh+emSGH3OSn++HUidhG/px01Wak
pD0WXQJnU0iBCtUsXnKiVjwUuj8uxN3ra2u+K2bGIeaBtB4RYUxk2VmCagWenlgJ
clVakFo2ydt45uk9FPYjictGGsD+RX/ETp3GsgCr45MGf+WrQYTfMJn1/9AgzvL1
8SjpD6Bqa3oyo5ZIuXSeKiLULyh5ry51Y7pEI4Hxc/23OYuN0lgjSz7xjZq01VaJ
/KAERiZd5PFbMc/UJ8jatq5ccrwSuu33nD4IMS4yE75uz5H9z/q41pFG4zGZ33VX
SMY7Kfe27GG9TW6Umu56/Q0Wb1TjsWt1kwjuICGRz/siBIbjAmarT7XvCPj0JVE9
A8Bxg0qcuBuysp6nyHhmPxflJd/AVWsxI0QBcURtOZ4wRLtA3utZ77HhKyH4F8RA
ydUUmKy8iETwk+hV77uzFBhsFWf+WE6n8pipHZVSB3hJ/GtvA0jjnwsfNtIMnPHS
ngsMSVmlcvBs1ATS00bHXw==
`protect END_PROTECTED
