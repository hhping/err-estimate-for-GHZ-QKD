`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PJsNOQ0y7DWWO49KuQ7d8ocXMtyCqiA+0JAyIvDZDh9L12F1efwIMZ7LwkVjgx/
GZeFb/wKcLcvlWsYRfk+N16clDyeJ0XjztKU1OluG7+CKUoMNalndZCy5U82tUok
z2Cqo3Hm967kCa/JYQiVHYaiLwIzd5haR9L6j9uDpOFJ5pEgZdoRay+Iy/B2/Ftd
7T8ia9CKKyEfxJvk8Yi89czqN1E4nHtzj3hRwwMbold7QnqZuXfx13UpkxaKDg5J
g2o4Hh4K5aZneIX562FVM8BHyTSmniYpusmCpnCFYsoh1aZ79r0p33roZlIiQ+aA
KvC5iCScWm6If+IG0Uzk0wxiZq5UrmvlgQmaRpPApBcH1GhkLphzmtQKRUYQDLOR
WYDvsxyAFJivx/pIkb74PtMy2ZF23DhY9RB7Gw+Nw1qaBbVC6ly/IlcCr9Z7AUmw
yD/Pr4Fnzh1vgc5EhYJGcONoC6y4D2MDMC4Ij6ezzRNm4xKTVtjMMD112YRN0l+U
2PqOT9iUBVL07/8UMYATY6QLLWUzAKfnX544868Ok8lhLnw9mT4lXrKVnPHO6B+X
3orTK3dEwe9xM5gQEhCdv8jHpwVugBqjeUm/h94Lg0zBKWVO5cMNV47JprnISXLP
DroW06DV7gMsCrQVTlIhcccOuWl9AxwOoYlbr9TzgzF1qfHI0y8vqwGVt3cPB+OF
y0fgUqx518Xsqif3PSt09RC+YU2iSjb0gqKPjXCAp05WIVS4/Mr8+v6yKNu9Q3c4
xn841PluxpTGnZV62PBeOzdEbjOEGkZ+/xFiEdWJ0/viKYwr69HjuCcie6Q32B2q
Kl6MSvOUTgY4VIV2pvJP9wzcCSaGjVNh5ETIzqLLYfOXAbJDz6eEyZDkpGtJiGUz
O6IuCTrY1C/nc4w2Ogx5p3Gv5OWp5H7a/1In3VI5HSz4+MWAGXxVTxwzqRMHaZvs
gmTjA4Gnf0V7XPAaVIR5IXxDEy+84JJS4y+HCWkpA4tjskNcujT0Aql3zviqEa4p
RhCDwRQpcFayrrRKhavIBKS1k2uOewiZQ1+bwrGoH1MBCPKlTz2cwTg0Wd7L0Mg+
6DCc+VslJbWgj0pAii9l7XHqgsy7Su3cE7j1oEpM4GCSsGFIBXuz3PF7Bfbo99vm
J/uEIr7Z3TjqqehnKNJDVgAxvdBBd8OKXjYNwzR3UhY/nnWXKWEjHXb3VpNxUXNG
ieg+Eb4hKZsk2tNjOgxsc5vgwc0+xq6qMQObkn0+cVUHeL35xR7cLV5WK+DLvxVL
WkmdW9v4at4z1qoPdn9p1X81RNo1cwFbCdBhCD5EqZ+BjBGOJpvNFHQY1gb7Ygf0
hsOoJNcieJut0iZUaS5y6vQeZzCr7hj8PvdC1KshgGQHGZuQAett+cA39HKKBeRg
bD5MV3Uf9ajpyUSL4KqfBCHZKhlxYqfuKJ5DtxupqLUvdqFxbENvdgdgmJUfL+aM
hYe4CmAqj4AWPtVKjbIPF/zLog6jkDXcoaU4mfGW6oZw3QaMN8an0UbqKyCNUJXr
TKpMS263PPXZEGazquTzw0UKULyKdjdQlbMbGYBlr+7edaE38A1Vpk8aQ4ZHrGuR
+9Mp/IQfl3f+rK3/W8Xpgl2MR6W6SgfWlpazuBzMsGiK0y57FrPTt8dOyXWt1RLB
92AxsNmjSinWcpLRjMou6n5mC0CgE2kujJYfcxjdlGPIiQKxwYbsCXf99+X9rxbG
w/Cq2sQHbx/h0UZ+lSNfBm81mADYdGJ8K4ecHsDLCIFWWJTrqBgZk8Ou6J0kP9w0
AljSCqamVW18mKZx4tsURTP8NXSdBuEq8I4TThIoq+b9DM27S0Z63jt/UgW4EEdQ
nRQRXhpi/tBIEUMoliuSvEJNihv9eNPpQMbsXYYNla0r9z9rpQxirinXQV3rkuke
mTZ0vIS0pbq1Oq5ZH6rl+7wWyY+Br6yCO73vyV/eB914YoclQFCCDp3BtNzt8kmP
loHRlArK04qrqTHeGliEL1Zjw0zEQAgd3ux9g/82n/5bLpZTrxrTBaKLZmX68NMo
FU9Lh2PDoiQwhaHFTObjaBYDkdjLhgx4UhnVpIH9aIA9/Rit+EJA3En9JAGSAiDr
DRzhrEme1l/vOhuO4DY/6snNzgqwu/AUQmZckpUQbpd050yfhRlQuqJKMM8ZGlm8
bmlbnXTtENMr5PnlNFGSG79haUiIc3isJ+L9NWycPQp0PASMSif6C1KNau6CbLw/
v9RW9CJzgZUfjNm0UXgUPlVTRaBkSup5U/jxjAwnb7bctDVPIymPdqdkWbuyi7OZ
7JfmEkhHA/JRPvAwSnQ4MBNIxvy5RIYAesv3fPetKnYt/mOVi8RxUtTDuHuMj3vv
wUmaC9HViYXW02n92yi8QQ==
`protect END_PROTECTED
