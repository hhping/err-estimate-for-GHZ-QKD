`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XW1e3J4xwcPl6s4U0mhIAIip8xe6TiNmubunIdtkSqJfzS89Orlae3obL9btgF0B
WIbXvn3HdjPHl4XASGauHC6wy4Brpl6652VRSi9hCaP4YomI+UBiuQvbLpdYE+0q
T1u3O/ITfUnigY5xt9e66x3ugyo4+cvLC2dcjs5g0MVblBmCDIofrEA5MG6bdd+f
b8octO/Kkpr964sjmHp1dOqkeR3rbuZthgjxccDPwZSLbsU1VoaMsa69EVWoDPHB
ETA4uMCo+k8F06eQ/tKbmVtbomOcvwGf26K0gT9ADvo7/XQflGyKRGqsQlfxwNUP
B+5sAFRHq63stVwYN+B8CBPC7ouVvIa/98alCwqHQYlf7GpunREQJTORn+YkVUfB
3XN+3Km1ipGR00zybuPlGw==
`protect END_PROTECTED
