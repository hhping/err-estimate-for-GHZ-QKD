`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFUbR4h0XoqZ6lqrsHmnlSQXEa6pbJKsP4XzAQeQZ3UkNFHOG2FpumDRNodXqNt1
aPgKLm1GJfz8uj/DiH6eXOlFhZ8jvM4za3lEwo4zb2OPd3zzmynVtdJ2bbMbnNxW
QXVOdwLevxDLp9FsSj8jAOXikRsk2dzwQjKXkoo/6e2R1U7JyfCYZbc+ADBYXSyQ
D08H5I/6FdA3WNCjC+470iOe9R22ZvgxNZedBOAKBgOMYPwzqSZPC2I20yWQ+paV
KDdVExoXnpgfkrCRI07pR6Rky//x4fJqfI/XI8Moq4pGx6fg/uScnQXvmahckqgp
94d/2C3ov68l8m7PnVc85D73hH1VmrlCiHc4HqXvZRexVohBQvABSSp2ig6GU68R
grPmwbThh2XqO7/9x+/1bqDHdnIjcUxnVWQlVntKQxEideGZS6+2101RaitmdRzG
9OgyywPyK+hTGzyVH9vhDgNjarFMmL1ERXyvk+eM0/hIY+HuujagnOmma3Q+3Wki
Dw3Fc+Zbt1Bqbvs0gcBcwYtIVOgHJluuY9gvzh3TrCDkaVLSZ8yB5J3wWvfczzmC
OknUR5ckEl/GGPuI8JzEBOzbnMkqfGMvKEM+oaO45Ojuj9M2/mm9Va/hSYEHPX5B
bTNL7crgUqQaJso6IpDDQS2OWKu/WhW5o7Cmxbqu4KZor3Wi79vK5imnG3R+/VV9
hP2q0v18XT/oqmLfdlFH65AycTKQOFwf3AOd4e+ipxbWJLpWSBx1INKi7YnihxUC
L/VBh9dtViv7ET+eWhtg7WLD4HTcKyhRv2X5NUcJRuO4ZKoA6jcKHWI1It0JznJN
RAXRPIOhkvltIpR2WWj2HMISINmRY80R7jaKLRpF+uzO0cfm6ZrDOM/7XWv7wwgj
j/5ZAM01un+WmpK8l1Jpeg4p08s9cSqNxxff5MkyVbumpuvNbMZwHMiCnDg+QFtV
Os1tNaOWv+AEa877vtoHnN+FxTJ/46G+cuJhrqtWrw3rBu5aeD0eK2UNhe1R9jIM
jdZwzXvtXzqG7VMqQlWdpdBorCdh+BiXP9x8p0tLvQauWfqt0KgfpACUuke47cbr
Pc59C7ELqJExD3pf21AoQhnUfjAXS94u+w7QQRwM30pw2zlYWCaKamAPm5Zl8ei+
kyBwAGY+IGBG9bHmZym0choy8nkv/bkF4TJNDKKrWCqO0HJEVpFOOCLp99pmXj9I
CPMJo2EFGiP4umb/asrc5OiK7rsdayi0LcpWUBr54+reB35qOE/nCfYqyRe2adeo
RLk1erpT72Ni1rlJ34IZ3PbL7ZjyuSfzGo4jEJZIw1eqf8gEy7O3fwp0s+8VmYMG
iec7ZR7kqmQXhjdD7Wq2CDkukb/V8rDtfAxKEPe/ERAeKA+UqdVhiLByukh1on5u
0epQYcM8m2SyTckmgLupeJYlt2m26RZQ4QjSlaA8mfrTQxvWkgzXN+gxxoR4lpao
Mq303nWglvmVRBNSE0DPWyrK0878QnF3sFWtVlwfYwROYdCGVTZzhW1XrN7AWcY7
oJg/u0jUYPL0RkT3lT4mtHQiiKMx5q0p4KH3taB4g1dg0n25tdtI4FaPuIxJnAag
9XdZonzG4e5a1DddqjPlf+mIAnqzpxzXlhOP2sCSRKcHDADaOlKxES2goecMUIqG
DK1YLeQknWV2BPRXtyjod+O7oh2kBBMJpl+OO1U1Wz7LCRbMNxWvhsujJ8b8hk8h
TMKxquZIvOsIcIDflIIoFzkqdCb1sCucPPzAKcuAMIrGE0i8ACtg+OcfruAtELTT
NJPio1Rm0VzqhDlm7YlyBoP36zHKVmx9hLMQKChXK3s3MZlybCzJN06Hr1Kbem4+
18bfgBp3Z7QpkuyRuxrE062jNIjh1+YSmZFhmH7w9Ik7YOH9qYg9oQNSgkrz2qH+
zm43TXeXBg0RlG5d+f4j+0GABGcw6lWm6fPkw1xeVBZP6HdykS8O7W8YRHGn2RUk
3VAvz1KdpMqJ655wWQyaHuA3dt8l12NlEHOe6AzKxwEJFxM0qBD4qaOWzN/AF7RZ
solknPcWpKFxqoGENWgSOScl1WrYnJaoT56QL20pzVV9HWgGBaKa/P5FObpzekgX
lXGXGw3VLyMStbKRaVtyakkhbaCrK1N9n8I1ePUXQH+Y3RgQOyAne4ex77LS87WE
iaPY/XiGhTe553WGbil69l85PXfml3eF0ifpk6+wU7moawBfmSadxadpqqgF3NRP
cZgdLpniGMKV3WF8RREsXCyeZCgrJ+ACbaIleaH/Aw7i267C+UVNoTdJhXX76V1K
06+yPFRxnxTrRfJ0qAJI99JuS3CEVmmeH7p3bBMSjFKunu4D9eK24hOWLP+Z0ljh
NNbFqNaMBig1lO3TWHlwiwpNWeVbl28Ml7p4/b9R/f3Y1bZYOcC8AkWW9hXnA1Dq
wbKsDjYQeb5vApNXl0cHIJAHXTkjsUoO7POWhO5Bo09fuThw5JmppatwW/qHq/Tn
MVDlqYEaH/rLaxcVZGCjzuzQ4hg4Qjjh3wtd3pnyFdNwsXA3RaIdghBFr6TXjquh
PhWnohLG5AwrPQFEqbR7q1/SZ8shC7Nwnf7KOfklvh11LbuvsBKBKamXTIb4rloN
Zp6oeTI4eIrwok/QScCE3hTNM9r6EtAZZ+r10hAeXjAA94Cozy26CcyyElzOd5+t
IydWRzeV0yg8RKUXC27ZgzTmYSK/WaU+GLnYIbdWQAtnbhBvlFK5rs9TBruOf9Gm
LIp3vUl6BHfayuqHyYAPZWXEsA9RrLHC1pIaFT9X3yVIYp6bO+pNPBNUVzF1dX4T
0wHLNe17oy1szAiJQgjmGESgY8ozV0xG0NAXPi81Dno8wp/6wQ6Zts5OrbYm6ljE
fW6luYu39WC2gx1o6lF4YspmDjvXZx/RWjstZXrOiVnTgJNBTsPnBrPv37N/a1Om
RoMm/UTTX5LT5KmaYT0dbzDcmA7V2pQhTm1r2NtP09nmZjSQ3pTVu5t19xARenw5
xI6GVSbmPU8W3OtOR6kxr/TPZpAxdoxmiQkei4eYM+66rpzH2UA+otJCZezdQ7XZ
07froDmJ3krwmft43E5FIT54oExJNdIjvpa30+B4mIu+q46PbmqmCQdD0Vp5nsEw
uW/NJryctFbGb4VNXnc9EJ3ihRTuMGt64de+yVIY+/F8vfMG+kKlHlm4i/vOKhf2
oEJuk105Ox/OQEoD6dse+YwSxbTlg6wZog4pBPsIlc4UQ80oW17oZCjp4jPQa0ti
ppnRbO9FIVU/B04I1HcLYP8CpBcyagI2tb7EXIvFbVJx0g0Zeeck6HcQJBqT5F8h
ZtF8eFfamy+d6WFAV40U41Px4PHU6LSy4+0k6frfC9xru9R89eJiZ0NOSyWS3CyH
3dKwrWV3uPgXEGOY0Wo0TCEqFDr5CVIPTyrTXcHZ72soZArE4MQGCPcHXADbI31G
3a6/cyr3YgsQ/oSCHEfSzfGinM8hmwMYxRGzCwpC/Eby3bF1rW9KGvl88OhkUAAW
gNZxHWRiSSBqbNSGysz0RAsGm4RzXuzjvF+my8RyY0AVZMQKTi7uMoBqkB01Kj1i
MaKz2fe7O5UqBfPSGjPeLGa/V/v5csJq2E0XIB9stM0pURw3Cgfso+l025wsZB5T
iZys/yXLKJYVGWPqPOZf6aASIwK22vy0ugsr6qbyOeWwRpOyfkVlsh+550jDtrU1
EBr7MnRmC3iy1Hb072DcEuEhYngsb7n0O5dnoEwBFBqc3SJD3kI0k2th1yru+51p
pDzX3VDUKPU0dZyptBP5/pi+qzzXayE32KxKkkBdhQpCKYtzhLuSPv3GRmC0CziH
ZaJKzkhNjk8u4vU+wEDP+gHfn3E2YmNVhfts3BQ6L5mT5xck/BygqxjdfbhxuYY+
k1Vo/xm9SlJH5cioAql+woJwDnaMkfg/fN+cM5GohLsYvw1Iw2rgZsrodTbbv8gz
7ZSA1/51u2WpiGMZmTI127/p8omsyhJ+Ay8lckhPkNtBrwFDxwNN7go3aB01Xkb7
L6OaAL+BeMszkN+t+RhQuush8+v4ZB4Uthutlp6QKfzeyFvafd/sdkrMYq1NjkAf
cmKW0sM2xydiERqYbLeAeHtbaFwXjwgXHSI1ZGc0r04kwkCKRhAz8onvC5U/5vGV
Ij1Nk+Ly2uvwae31pZXCfB0la8aZzK48Y3xRFCiAG7gQwU3qSbTOTk4FhhABP8OQ
yppn7UWcg6/lhMXGK87Llq8FfXqE/MZMEtg0ezBRql3vU9iiPMNHfg5Gm2Y5QuSj
ayURi5ZFp/xoB4f8t3bgffIxNC0GqO96aa8q6MP9HboYhWHX67y1zZ8wxcZRf82y
axYlBnlHh1JmLfGAhIDVCWqVO51mJvHT7deC7BBc0+kdvcFQ3KOhCy/ARyugE16j
1kYFAoVFc7AZHi+EakA2mKeOLMUgTvd3ygmMLOjNHkcL6ASeFuNYQWxFzbgWH2pk
O+SxnODZIXfbuThy9aUAG/YRVqq90hhKwQDz0GeL49YA0zQRf0nSEN9ReBKVV1Uz
fVlqevYcmyYaIGZzeF4QvBNjUCy50MBgKt6BJgs38VXOeVuhEbGZr9e+akNycgrJ
MKydPh4+OY6uMr0OxKLvb89Ai3MJJivmQ/rRUBn4pm8tNinXNPTPKKkEmhcGGjOe
bm3VqFgB9B9co7NTMkN34dCAwxoQpTUpgChz6be9UKTTsyV/Nto3eEdcLPl/V7MT
j8zObUMSgLOY9m7w0PxTrMv9ZxjhBOFD5wd/YHzC1RUg93/F+q4E1kK0mAptsoim
V33pScLm4yV4h7y/ltTB2ECofL9IW/Ac9cl3Hze+jHC5imyKHbvxHu3MQ7RKcLhS
Pl6FWihVDg0nY6PcnNdh5XO+2AHqNMZb2i7WZFhHuJ4Grc2NPSkGrm4vImMaOf6u
b4z35eSWJ+KPCPjpGC14Sbh8eN+iPOPhVxmkPoFhNP5KNcICt7IFXRibvbX+7wx4
3jyXtWE9kFEWYFYLukzTdJh+nIl9m0lemb1KYCSjC+QHKsHtMqB+Zu1+FNXn+zj0
pVE9WhKNUlZ9SYbBNkTkZrdNJ5w32SybU3EZplV0gUtwLCERFm7YPotGSlon0G+U
ZD7rK+7NwDDxltj7fHCK/nr6kjipL1KVauCPrtKcg1zEkwy4YdxW+PSrqYKp2F54
ZicWuwKz+u+ykxLPIEvJwEUhORhw/W8LtJrGrBb6hFvmUOVHQMxivGeg4oCGKbWf
kHFpUd8NgU1Q7pGEOnrcEWKKLEALP+gsyN4/595NBeeTvTFyCfoeKTBOtoUsm8c3
NuumHJIqzR681BDaoWa30htNYmGLIj1iwTNpBPtB9JvvCuwVfZfg5OLPVWwvQs7X
3NWUgCnfvdgSso17DQgQFk2g05M+RWVmiB/m35OaxNBRxePWEjSaGrHskvUxHgvi
LVReAtGlkZsjWUH7eFpuYWLTH39bS40O1yinYvLixOKF3rU4K6A/DAwxzG2CXvRs
gErY3gqkJwhKErhKXYWxibl7Ly/xf/JLKo03e1e0Pnwljc/UyJ+DeHI+8dlKRk/c
nMtQghO0RTb3a0X8YfqP9RTZ9vdKJ1SEXVIUCjPo87tFzpcMUn96MJdAijxikVWy
WUtoGe/imlfT6vDW2gVM/XGmK2Rp2+EBuy31t00A0g52cOYE+eZ7kY18y7Et/fCK
yfzyUuSXEr5PpMQLmbo4JYb0KRC0OLF07nFOhHmibmsVby8MxDRsLJwiOumIRP+8
joJA2LrMjxkQnqTLBS3X3rmHdFJEB2FvCF0elYNTyI6ZJiaH5X+8MsFaQ0PZnhKH
zMrRaxOas3uJwZ0nJrvMc0HliRIW7yKQz/SUAIgVRCu4cYEyiBYV0z7UxAgp+N5C
Qy5NtaiRSn7768SCJ7fYPqHPMMdbVjlO7kUAYHrUaS2MNeUtcZ2uoTBzjkqk45Ma
9uDDbAGyeEpju3gVRsCbWNqz+uePU7UHqhun7upSpGVpA6IgFvLpqMgZoGN0bNr+
qgNQ/5n1Cs0Oaf1QBbhlQ1YFv/e6gqMrzOHXnd08oZLp5OCNk1PNl8iMkY9ijoDk
AeG4eNnuGjXTVxT7P8ZC+BG7ly06a61y55JvpMQRLvoZwizvJahFM8nkw8p04X1o
Dlgi39we7cNZqQpA2uvZ/2Ns5K7oRqNnXxZK4lvmSYLKPwef+OuDGBb8tR46PUlH
yz6bx/OowjfhvIqzgatISq2Exh41TSJLNIWIaBQ/Ct9M3PBVSalHaxtHCoX5v8wr
/IqeF3U1znPMSKKUNXZVCgBZeKA0Fie+XX3LqtL8wpJLlQSNpve7PB+n91/1xIm6
XDEh9T8uRNR+Kty23cYfabWJVlBgmXYpazOKv2htOr1Rh2GXkRr91Y+3G0r4kj7D
ElCYOB34XZMVXGMYigiyAUc/bKy/LNSlYUKKqYWsSF30axruGfrZAl7q7tDhv9a4
I8W7KbCMH/mq/wwAySDZ4ussM7SjOjF+7mmWbaBXgyRP0ElMU8HQA9arOq/EEmmX
kQZdF/7lhVGSMzEBPAoCp27Pnu7CZIK1VE2nDv9CarH0fFB72KfkpgK+Impt9VV8
UVEL8tRTNW87viqTyALiiAP34d3Hizo4NyH57mDgH53tIcL3Y6gYrl1NvZwuONC/
m5zbxITazk41DKEMsVO+RnvX2uYA6r1mjUWSUtSkqNC1PWa8N4ceLyMm/90Zy+vD
Q7MmcUmtHogUNTu1RfPbAY4rE9Dz0SCseqGvjv4+A/DkLsvSGbyltOlEOKn+Sfm9
ArsLPOFq8M3nTr8Ec9KHHUKcGgUWKjcWl8IdB424h+3wZ4WVrmOLwZDVpPRDLkzC
ytRU8neAw52gOlCBt9Oj0NI/g1Ha5IbgoRzRLAOCUhKSIReH1QvrlVNlg6ylqQJY
dSPdWjlve3cd4a7yPkG7V2OXZgekYyIKIlWMVc4CENgJm36Z0wdXuurP0/nQ/KT6
n6PidhSBmI5rCr3MCuxNIYYMKZv300JMpnWlJentnrystXNQ22h4DKAiF65OzwAQ
xODr0KidvanEL73qEGX1dm5ZcYqyGGbR37tKRTn8OB4bWf5tKTSEFSKnHbrbCC3s
7IHQ7ZkST6EhNWdd8fqEMdDAs9hNmXcJ4K4hW4Qr86QnYbRcHLuqhDQ0l5wpGb41
+8dXOXQHlnX+NaOYoKnDc5zq88dm+a+bJTWmI8kWfsl1wUW44bPLDg0CpWM88BHr
laGjsAYgJSdfVtUAhQum8S0S4EjXv5NavbTSwmwVeuE9Q5ZPt4VhL7JA9IcRybvc
X1iyow8GySv1nN7t7GTw0f8I1nhatUH6h2JAMx02ZbGTjatbST51DXN7kF+KpX63
MaJdaWRRapjp7848aDG6wwr4VOTEaEwNDmb+ZIs8IcbygCE6bor1bKNKkVvjGop3
3A9Wa5hHCNTsCfbyTqzXIeuRCbvg2IgY8q73LNHXFwfil9vDj+LbfJo+5LGvMN5v
tNOrHhpQ+2dWktjvN+CI0VdudvffIfcpZm7XO0nOln95Gc7EQ3RWDh6JhdmiP+oK
P/HRc81YfGI1F8VJzZZ3M7K/eMUj6BE909pO7+tSU0Tg/pT6054dEunQqS+aYOEF
qflyL9R7qR5E6k7TCtbnH0baW9XNGmoDiBfZCjYWLAc++Bl246igktef/NFPQTP/
mOifTI267le5RAK3+HTfe2gnstk98xnjOFE5qZFDJSt4WxHuGrvCrikzG4WCK+f+
pxmDXr3L3sOfgEqPl99iSU68M2JIrql6cmm2HsX3rw+fUqB1rH96CZ47hxp5lcHP
Th/NkCFz/KgO3oaVje4ZtlDX8TUZxLvPe4Fny3cPKpyQ/b2YDQxe1NiGinouNIUf
5TvNyzhk0g1JUfsGcljxQ6B/M0GPKPUV3dtdi4E0YIqTrpsDhC4iC/nZFtMLE/qe
7H2+0SOeHewexlll/f0ty/ODfMCzxDNWuEpB2ged1gASpkQRAFRW2VJqCNjFZ62X
3ichrnpjJr+YhUL4kZsao/EkGW59jgatBKuMnrd5zyd9K2EDnohIbi1wcwcFXWlc
1MWxCDM6XpU+bWhfZTaiCo3+Hyh8Tz8e/ezKs8bjDUqHYPWbCuMQHV1UjCp32RmB
Bw36bW44HWGYtvNJ9G1jW5pBS+8XEsvhEwcxjd6yTRGB56HqLKfLNqnAZyZ7szsr
VoSN/gpEiNqlKRbq54G3jCKM0aQl51oFp0pE+O6RDiDTKbm8z5IcjCAaI8tb4qAb
4G2bmQVym2Px3Fz9dTjLDTPVinjBY+iVb/mCFdnBvz/E4wIljAscfI4LlpxpiT19
lh9yOeKrDT8iRwVUlcEtVUa+YDUNJXO0JRRDsfcXjezqK2ktmVUsB8AYlDYD5GoC
38sG74Y3APzIgoXY8NCazKXo6SLf5mvjVkivyJSkxWT13SDMTxi9ylFzJEpFKUCx
oj2D8TkVebmdiFgHANOVMBCJ0z8FP0+nJxpBY9SSLk8to/JK5N7jT1YcucCXr7lN
0Z/7SJjcJnN9tXXWZMnlS5U+TiFyFMP24W+uBmvjdcBq8uNF2WyZPilh6HXzHvAc
QRaO8buatyIzDbizjmYUqo95zt7SQESO8x+P88sQRWcOX1KgfxqEQDO59RotVBb4
7D7mCyWo4rDKV8wcFaJvZrp9m6h6849+Xa/HPHkRl2hjaPdoUAcDJt4VFHVYUb5d
Xe88D7aPrFyUppG1k6yR9f7TzWRhy2/WtUxc9MgVYYF4iB4Gd9PeSFqrM0yIaKT2
97m6GVZ/IVIoTklYsa9185qJqKrcYfkNfMY8qs/4+mckcMg/HXSjldz2CsaLz1X/
B4KgirIbNAkBb91hCDMIcDZ2yeh/hHrOpvEpthlNuppUNjYJOLftpyIGxOh5T93j
zoGkvHasG/ogTTNldktw8GzQJaiPC0TO302ynbqTPugUADMGApQnFn7sCrSwoKWi
Rx1pXJwP2KYS6APB+1Yw6vIbqrq25j88X56OoxQnp28IFFkDHzUO7goObgO+QT1Z
KyjeEA5svqB6kcwKiK4Da1aoHSf9jg5B8klVZucVijCZeNSC+VKskrEKLh8xeh9G
vKoHe0fv6R8kocJOgLL8gokUKZZS/49VHmQiXkug9xwjaVUq8XuxTOxIPqMD5l+g
ys0/+5GL/bClyJFYvwzO0bYX2WC257Tq4FJhxetmUHueFRZJC9yvKnL/33+FSX9Y
wZ9c6qnj+8p95K2aZA2UwTwdL8A7nHY7+CKZl6yyITw5boDCqKI25S9DOSl2UMKb
VO0icJPIQjCdZkfJnnHN+X9ZE4+ayr3oTTdEAtVAEUkdUpM3R1kZmtChRk4lLSlh
AwPpiiUR+EqYLgwE1ndp2aVEmt5teGpsWSMrdZ4ngZHBvUtgdzIQT2X0fwB0RjVt
LWe0yRaQU6H9upn8RhEhjGAOYcfE7OR1yIfl3AZKuGacd6C7K66UzwstfrWCZvJG
PS7EOdYWsA2qOio/eQ1iCQfCi9PhiZl/wNrdLjrp5CPr/0UpOzCNccQQ5lL+e06R
spWI/DHQJ8mFEljivUnbsiSi/+nTdSota6awSAlVRzO4CVZ39ugygSHj4aeAW+EY
dR3kORv/sRGXLuKakdsR9QGewDgkDruSfooOaY9vK4rxRAHjpO8Tes4u2QfHKQ5M
Ag62yV7NcM3AfyxeeXFXF0IOGUTon3vaTdb8SaA19oiumIzHJ62ZH3JJDdpQuYT/
24FtkPdQilt1KS/1fz+UtfFWy+Nfj15ru0Xn3++Zab4Y2MzluAIeXDWRVxLyF2/r
7YkRW8nwO8jiCNN2lVWezH20c0OsKCJ1BltuICGO6bYIba4M39W9LPThgrr0a2i7
84ZSwFv82XczUcgMt5L/Eq7jg5qk2a/KQ0dJQruYGnc9wUnwyhew4ABKOU7J+GmB
D95m50zHAFYr90alr4ctq4PM8qWyWA7T/JF046tRCrcLVRRGU3kiEaGpXXLNMzq2
KUk01fD3GbKfUNb6BMQEzkZgf+dxpj6tuV8gDGbSDlSquGd8zSpO1NJNfXm5Q7x8
APFZjp44QuPrIjFPYz6G9F4l2fiuKWqRt7n47jXv0oP5k4xhXB1ZhTthjv4NNYt5
y3fLHs40AfiYQzhvJYeY2Eah7BKoqIdpDz5iAl0sghTt8a/8KdakA5v2WJWViltE
TrpSMn4ispv1hRPMDl5M9ulIsxs3ENwBADYvV1yWStnhDDoj24DO/ZAWJYsp51IO
NuqwldL6PAkcdG1g6eLOkbIc0lYl3vgXC7QDjFkHoAiV/aR0RIkcfWqEMNZ1XcsI
ASCkyR7+iHX2JMD3PQB4FOvxEdEXuU0sEZPBOTR+lttlGNf7XqPQ2m+0683tQ5M5
z0nmwXaHsejxqJVQbrj4jVFZw9aCBCbmDB0ssiKq6szvnh24Sjio/u8B7OBuX48I
xJI9wZ3FblI2FXFH9ASAbnL2tfbkKSvPmFB0DE85BJ43vnuLABC3WVmwNY3BwVSn
`protect END_PROTECTED
