`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1m4uSA7RkC/uCYROEzBH+u4+WyxlfZvjDGHElxfkA5OLWBtP2EGOmJ6Zlu9LGLy
7lx4JS+f/etf0io/G0+nqhLCv++jgoiej6SACrwivNQjEbFVm6feEiXML3OzyJ/j
qLaUKWKYJczMvKJud1/EvgLpDJBtKTXQM0e0CnQvLs+n5yE91aNeBajPLEtfNHzD
Y6em+tp49e/cnuV+JP+6qcUW/AZgdnRyON89Qz/hRtv8zZOofFKi3Pf5f0PuAgGH
pp1+Ngyz16HID9j8hDploldvnTS5p3zsFOU6rGPIfZI5mmNUEZRc/Z5omayu4Mij
UVPxjSsU1kjmAbi3GsC4sjEqTeiKrHMeJEDfX7s25CoZqJUdepczKN53CSkTzt5P
UmHFbYryo0F+qrzTmlms5ddMMtmhGGR7oeK4IcG0CyxeVMZnsmevDXI0lZRe7GLY
oaI1vcFe5CSO90DIX4QKYnoAozwnJ1p2T4NrCnxOROTF/KUZX0HP7Qwridpf3IiR
pDbXLXDdQ1bbhXsaWUXzXFs+jgmyFD6hU+XmE6gBWDPWZp2iCHJWQq00UZhuvBmS
MjQ+hz65dCxEZJ7NE9Q7AKvdghjpiYaQw6GtzpGmqOBBnVwszpKsN64XYMS/zboa
98V8auI9QOLOcDpUpqg7epD65Fp4YMWclrCWiW/0gHjFUctrMRsMnatNM2aoRsyV
XYKqMF2m/FayfWNLCgoPdzMxQcearvJYXbJtwoxkM6Byr2/uFS6FyIGnAETRO4LB
7ZxrsRlwv3I288eSlBajYKSeMzN8WHLodbC1wxZOzk2FGKwIHv7iHzVIr4IjPG5+
Ls0f84F2BV1mmoPV10RUoawYDpgMW63YVxwZgJzvxm1luYHm65ViDxVffPT3DOmo
FsO2oZ4LIAzlE7atdCogFoUdTl5ylRoYHgyVlM9ka7vyVCEoGp+Rswm8AfoJVYQf
gogTKKbNNyVYBLAY2Jmkne7pruRkBPSTr2r3T49U4+/rm4d+WExnwqRe3GHlBeqA
NCHjVQAS0/Hp28pubEAKzZesLG4e8HDcqlQBgrypTAemeR/rgzHtSChrhZzbbt4H
bY0lIxf534nJaZ0SMU8T+Zif/96vHZXJYD/EltDZb1mjD4oYossWSR7OIAxz8FGy
JDyiohnkzirBUOYNdWc42rqe+rkzYCyzkQ4ipScJVUYZvqXVCZCrADPj5TzRQvAa
OO/gWaen6Hfzz6uQJrLqWLV2vCzSMwA76D79Yqc1n3rTQrLr9gvah7F0pO2O0/Bw
5sNuk6Yc7UijpbymvHqUkY+nsU70hE+uGm9x2KBMMIKV7Q1bliRtWIObGgj213mq
lVOUAe2NNTGfLe4AkYawOQJTwU0xkjF98I8fGWlRHIYX3LVz0ccv7SRAoGUKR6UO
JLsGQVXY/5HhQ4vgojF6ANKM3gQNZO7OZrmAycYL9lS+huxuKNgl61aJX4docLvx
vzkrdNyTqOjWdra1+MpAhdxyYkoXLVphicK878ToBn6wExfhsrPyk0fOSqmGcMmb
y3aEiAojx8J/msC1BamxDCzij5Tg+xa86ERl/Nd9RQxui9MOQtsz1fs4lVCsxEqt
7PlanTVGpqq3wzQalSV7RBYBzFJhI2zfxQ7hG4qFXpU9jUJh12DMehv//tPR4opq
YhZzEn+uJPhLwKBQsEM4vqPTyUvj3uO6S4FxLldYvXNjFRs9YGru44pFcoYCbR/f
yJ17CtYjLEPXOUgMvHdM/RQYTZuGPyF71eG1dch9Kew276loyXfjO3L+2GQ23BI9
ks3MNpNkpgZY6EEJE0MFiSj6n3bBVzX3C53lG1vPiUFBCQUvInVB50rzqBX4Aggh
b9c5IZGBkV4bpW15GBxjqUX2prpby/gJyer2EEJ9d7i54JBQkvR+c+lLxDETmtil
APWoHFJixnZjyNayxlkBBSw/Mi5lYP6IPcU+K6d16u+qOMsL0RDqiPGej+K7VlGt
pG9r/mnFHuXZai0a84D/+z1sSUFlIopj/5+kB7ab2mtciVQnJi7DXYZtnnGZ7xxn
AzN3AQbE+ALIp/KOeSC4DdBayKnxtVtfGN+0CHA+05T+XiLOeRhzWsSkxYqqPkli
II7vP/XprVw2rTzqOvEG9SaGH1ZxjafvRds9yg7ZsGD9IHItuouoF6g5uKo0IVwN
TM4dkaJSBcqu4VDQ0wrRZiq/tC0Q6/VkpFe2vZitvFSplnECx4vFjEbArJ8Es5SU
sX+jDPJPLZ4vmhgEIDQztsQzb4G7UT8IfDVpeB7K2TMneP3+zphqMiBEvZVFbpU2
1u/gE21UxFfUAdqR63iYhjKj+UHLVeZaHMhKYPE6RzK5RGxPJZq2Jcu6tGZ3P28a
avnAfAAFI2+hN1gwKoPtoc/QkfurbJbKdVmp8YZmTm4zc2tj9yGYMARi3mqcr3wX
6mgp7nmhtFvSSu5zgZ3TeVjLSfYl3izPel4OfAP2egqy66hGqD2sMtOBMIjvy5Si
iGO/xyBUv3rNXP4Ul2sp6LVsV04rs8siUYYIIGLdley95wM+mNMl4U/nHRGFJNFA
ikSfAQFsruc5A1uLTnWLNPfUZbSHgqLNS3A8bDZ4TYY0d+TiUs7mi6DP6yBS6L44
z4yjfDW7pdc0OFUGZi/O9nn7x5Tl9E1TUVxQYPFF+v+UP6xmTNWNhIlS4qY203dW
fo38H6Y3WYZhMcao5pwYLblu6KdirhReI+EULNIB2q8diKWPhG3TF0PgeDaqVbzo
sugaSNsQP4ET+vtWLRByub/10Eja4WTMqMggqhTxm/zE5U65CcNst3zx+wAHfJSB
ZGiajuCWzTJJXBabXQRAxPVz8mF8iGAKhnGW3nkr1h5ce1l7ws22ld2eQbaFf4MG
JHBRd6K9GEuOMk49TflEbv04q9MWANJE273JhfljGSpZf469eU1VBwktA+7fUda4
pJQMn9L7nlsnEk0QhkuSPsuR30QRdiVeTLJ5t1HPxLo2/7RmhnXC7E3TZuqACFTX
qat3uKI2zbgvkCGAmXEjM8pw0/aTis17lsHPzIpUu0LgwOODW/rsj2Z/gq82NmR1
t4f/AKIPWk3Vda12sg2L678d2vxdNF4aZJjC9tIJQvipPC9gi2LARs2M5OJoV2+J
IOTY5DHzdSFyPJaXSxo3PJ96oT03vvJ3eXrJv7iiYhHgiao5C76+xX1ZQ/hM6PYw
vGg4+tShouN8uhZihfKNj60hHDibnlQKWO29kQvoMt8b13tH4Xe9FcW4pezNY4K3
b+ZSXDU3vMxxYAWqaRn9YzduaWKBTVw92FuCTt4ueL7+TN4AU5Obrz7uq8jTwVfE
Z1jMTtheMDRbakwI+pCK5LzoeNNoh8+IOivyyu/aDp3vBp6Dr+EIKAt0V0vNJJ+J
+RQI2YMgnlpHf7ZtJ2uRSe121n2KkKz5Cx5z9OyIP11/H+/8FYGf1Wt0IObyZxbu
yODleuN5AFHV4PyNrtZ2iTLaCEoHgbf5mb0QPWbID2tlPr0AtvIQtV9dwkDVq/BB
8QtHr7CHngUCNJevap6zYx9j5I1VkA0NqijxKV/6b43gh1zh3NUbdUxsRnrawH5y
cXBOtQcXpRW7rqX+BF8ihfKEDyqdrV8CPs8QAxfrMQPwA3Lz63hQruOlhYDN3350
TRr254H+0WAz8Kjvry2hwGJje7ZZ95sP0LvJ5XWj0o2oZJjxliStt7doWeSY3duj
WjeE664bpetUI+dv4P56IbtomUElC0dSNwLRjw2Q7JyhMuIwFUa12XbfAJwmclTy
2j+rB8PCmL8hH+6SReRvhfEn23/45iosFu5AO0/58OLOPJiPP9msfHPh5FJDHRZo
OGFS6LS8Z5wZ1p3O9rs8BxKPcj4sC3bzH0x4gfJJ0UzhNMlRe7wIU07A1E13A06g
CWgTiTqlgEf+tQtMR8cOqjYTHrvlqSDZbIXL5LEe56U4CyRYAWuvB6bEC3KwCEOp
mq+Liuuw/dd8m3he9FoDKi32urBE50P0Sd/CVmFxFZ0BDJUH4fXuRK6EUSAe6uiZ
Sjw36yj9JMAN4e6tTixsACCmH84DrFrJMWtvU4p+MrLEPjWDHm3PMrRWvvMKVX03
IJ0bem224Vt09wpyRUeDlAK+IdzZcoLq8UYfa7DsCl8iioQUAN4Ljg5rRQehiMnO
kubJsWr/Zl2biOICmZNlRTjrvrnqidhw4goagihPmb0cK36ZxyCby27MpTfa6cvE
JO/akALzFbMFcS/j5hbX30cfkAnEmWXAwh/3AeEaSdGXOH6w7I4ZA5n4bJdaxvkZ
4zYl/rBZjU4IzdjsUeg1+gjKCjnQ2HsLhWwgHIM+1JnK+6oX8iz25elZNGLLGlsG
52BysWlIk9VwuRlIYExXmN4sFnNuBLT3WjqxD5Wlsgwk4WJDXpBaX59Q2/j7w2bp
GrsQKUoJl4kvNTNskJhsnY0QhJXCNnMlIXuD7fu87y7obVwLPBNV1G6se8w2jqaU
/BwLya0HCFocGZPLETCMm8MSpTcWWfXFL1qjA/FbuRDShmHD19zU1SrfkiuZr8Zx
R2m1+GROmWhdvZC+i8T+u9u9/729ReTC/YYT8f8IPzBneTtsBk13r6nlq2dUaV0Z
NB9BQtEYW3V2wIJ97J/rJAnKnwAW6y+5qXxy8pL57WIVS5UI8HHxT32MrpDVmx62
e0+w5tgMDD5F/a8vt7DoUH/QP5AJ5Qbt4rg0lGrhooMZYmCeIq40PZgXAkLNE4tm
oxRQRliGrP55S6zpN6NUi0oTZH8UM0tQBE0WoZQQ11CMt+s9UX5EdoZxoaw4P/xU
6eVZU2WwuUeD8hqLMog8pSATT81GGpFOV1enQtW/r4BAPrXg2qSSV6XoSd2M6C1R
xbQbrDW6vOvdvuIOO67ewEOMpUslfDiCCxkzF8yM/ZUpP3mHCcjiHHx86j6wZyeL
Ce0s7Vudgrik4QxIKocyJgynOaUfInNqM4/k923dHPF4eyQh7x0haRiTuIatJA8o
aAQ5HiMrLMrIRXY4GV73qg384aBPazvLnA3MdTsXk3PJ5lR8aA1TKLqsDAhQiMW4
ZptK18/rqP1cop4ijwBg8kG5IL50g4Gq5U0GVLj3Zd/toZOVd9PyB0tlEnMTqkgP
BHwFavxIPWdQvV8FMTkcxDrNxrykCUnL8oVCsqAqnxL6+6qRzIPQvGTYsfb7LDy+
Kju/PCelB/bEWIujxSbDDVB5+PfjKpNonyLz0sqMAgG00fRHek8cfrP2oNWRtCHo
dpUcYR3QrgcOBRXPiv4Ermm0x3jHGMzYtnwwCVouVQyVbzIVqLChuenxgK0c/+Js
fwnjELf8oLHez9uRrTD2C0ImB+UkPI+UXi9Y8+gCalbOwJi6NeltoDTBfn5/epRd
osAb97a984Yrbm3Booc5jbuhndbmyXfrJ4qMJzBgtJ4hMx2MugNY3Ixl+2Ld+wPB
ml51YJbGncHRtr4y/AMawqpxUK902hCS7lb95HT8JXvlJEpd+BkAb4yBNWUD8XU8
BBQs5TYzbtW50nB7ZgmDRLLLBs/anW8eHOwaqf/xdgOhp8Je/G6vaU/smWpoYnpS
g1AgS78Mo9P3xfVLHnM371JKQpgGougwU3mSVm6oZmCIvObrq+OizQeIwuFQg/wv
fIwlClCkEjpvn6vt86j+0x2iNu6swCNleCpX7wWAtFxadfTrWrkNqwwD/AN+hmEU
oeoft7UTxbDZkEDtSNk6qvD8GvrGPKFwckiUU2DaeWuGR7ezhmwj8ksCdWHFOWfx
RTKuFPLyW0kv9b58UKpTtMtw85MHENLdrKMTbp8b/M7jEAfnoZwR06lNMbzu0xvF
qM3I0JLoLhUOd9H7CraktFF1irfeKZkdwLT4dNXM1LZhk1/hQ/MAIINDEoW0FMXl
gmwPimjJdgZ9+twKmR8H+EDyfpfPFc7NDVeetfcV7iVgiHLlDU5PvGuor29gBb+i
M49dbj6jcTtZfR1p4r3QUfjl0x/BCZuaAncQgbevQt6zIMuDhOKC+9mhjitzR3uS
yuC54Lp2A5cBEft2F+cC4YrbYx1gbw1aC5cCYCSl3zX95e7MZ/EUWVcua+fx3hOD
zNtuqiCXykC9AeuAXwuQippVFqYYYwQ+Zc8x5gJmMOWIZ7geN82w0OlcDebu2OsF
AiEGW43YNIuiB+3dW7UR0JaNZT0UgmDV3VJQOoOMPPo8Nx+MZwrjWckWwmmvFflX
5FblIhwW6QzAJePGkqtYLezsBjSiFWaO0/MXPAWcY6WoYsbg95UjN7YP2QcOTjA9
oNJuYibgZtCpR65D1QuyOA6TpAf9XE6PI80RXGICWAW47Kxj9o0xc0O5R75x0YHd
q6/w/UPv2JZCVF6pUAHT3RL8hAvPx39ZRCWk1uKlLxdcyVW50QzANAYTBxk9fwIM
WK2Zrwqk4cAT/gD4NQ11E6hN6cYMu9ism2X+l0tSrScQHYaIKHwOkFFLZchtEH1h
tNWnv6dBOPiivpydRAj9Q+EJrLZRX7t2/BB3WupnMwJH0CgbFYbJM/gCYlk1suRm
dFxE+xxFshcBI6DjUQEqvtA9f4ZjRq5GW/6FAf68YKh12z6Da02K9gJw/mB/ltAn
cDOvwTh//5fUTlSjSrzsKyG3gYkG8XPdjY+oBhtMzjxUeiDNE0hlnm6QkA0bLpgW
N6Qu2wDHLqCmK/rWiAQzDl9+Qu91R5OkOeY+uTtaLIKPy4dLQghJCItqPh2+aURw
+8y7watcJMAnC9aOaZkg3WQ6yCPFvFfYWVOQ3h58yeWcgT4oY2apq2UdDm+Q8h6V
NoF43u3yAiDtmLa1+gSCv2n5rfTgmDx3tThlc0Oa9p94Obnc6QA7eW51Sxj5zLn3
pGsHVZtgwtRQUe0+ss9c3VY+6l3sWb6ChsMIx12it/xpwF7BAzMdfjRn5ZXCgK8x
DAAYWZqcUthUYEfKRov7t+u0+etv7BajJwJsmKwAsuOtMKH8YsJNggxbIDvG8WC7
lyZ5eKpAFdDqy6trrLRSAs2QZEUoedaMuT2nojalM/mLF7xHrR91ysCsWfU/NMMI
mKIYduh0WbxB2f7Uj8C8NN6tQlqq6bgnDHw00AtO+aQ=
`protect END_PROTECTED
