`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2sbOQYxZ3cVkQp5Tz4UNxl8eB1TWk7yIlNfOCLXVOHK2XdEwZxrcX0EwKCYIcUjK
fU+kSQymte0HeFuCnD/HI07F//9HYPn5/UqYNVOxHv8YqPr4MJR99KNA/jHg6CjB
60cjHJ8FCn+RWzJn3OO5S3HM18w0nSagVvkN+f9DW4E6yh5F0XsLhpEomfox+fot
TpvE5NQmb6ImrCTH6NQKBVEOkkjI+WCe5GV9pZ5xL77iPTJVA61iRYnhH3I/o3/P
LeColi/DJfZF+QuPxWUTNZUebvRmBdyeuQFcFko2zmc8AzI+P1Iyu/L23j5qmCGu
SmDwL3T0aUuAZyLNhzwtE4YBS008+ZUgBrBfAJ7yAUOLnc8qfPhfsAFEN+FvPJV7
QEg4+h2+gvKS6Qz6GyPi8dlBt6h0m6aGlgShLD9u37q1qMuVkQxlVFuJWnTESiye
rbk1wOVwYvGJOvgWL1mHJ3wZMEH1g/pfdHHEaou/UYLcCGIFhDVPmidM2Er3KXNi
709AIUPWRxB3TOtkpShkj0FLc3EJtGQzalB8E5j7hjfRdXf9+5JWbUMGz54XGDHr
e83XmseIPFpFoyQeAifPeZ6jlQl3uNbRcQEDVEG+56oVUJUgzmUDn2dfRuxdveYZ
YFKXR/tDeZZ+AC/FUX2fRZBHdc2Wv0ixEkk4yPcMs3uWOmb9Bmwex5jchnvrUjUq
tySFybTeMQ1q0hu+jTOmHaC/Jy9tS35SvstYilT5Cuo=
`protect END_PROTECTED
