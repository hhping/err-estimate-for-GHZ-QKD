library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pipe_gen1_2 is
    generic(
        enable_debug_info: string  := "true";
        elec_idle_delay_val: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        error_replace_pad: string  := "replace_edb";
        hip_mode        : string  := "dis_hip";
        ind_error_reporting: string  := "dis_ind_error_reporting";
        phystatus_delay_val: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        phystatus_rst_toggle: string  := "dis_phystatus_rst_toggle";
        pipe_byte_de_serializer_en: string  := "dont_care_bds";
        prot_mode       : string  := "pipe_g1";
        reconfig_settings: string  := "{}";
        rpre_emph_a_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_b_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_c_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_d_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rpre_emph_e_val : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rvod_sel_a_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rvod_sel_b_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rvod_sel_c_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rvod_sel_d_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rvod_sel_e_val  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        rx_pipe_enable  : string  := "dis_pipe_rx";
        rxdetect_bypass : string  := "dis_rxdetect_bypass";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        tx_pipe_enable  : string  := "dis_pipe_tx";
        txswing         : string  := "dis_txswing"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        pcie_switch     : in     vl_logic;
        pipe_rx_clk     : in     vl_logic;
        pipe_tx_clk     : in     vl_logic;
        power_state_transition_done: in     vl_logic;
        power_state_transition_done_ena: in     vl_logic;
        powerdown       : in     vl_logic_vector(1 downto 0);
        refclk_b        : in     vl_logic;
        refclk_b_reset  : in     vl_logic;
        rev_loopbk_pcs_gen3: in     vl_logic;
        revloopback     : in     vl_logic;
        rx_detect_valid : in     vl_logic;
        rx_found        : in     vl_logic;
        rx_pipe_reset   : in     vl_logic;
        rxd             : in     vl_logic_vector(63 downto 0);
        rxelectricalidle: in     vl_logic;
        rxelectricalidle_pcs_gen3: in     vl_logic;
        rxpolarity      : in     vl_logic;
        rxpolarity_pcs_gen3: in     vl_logic;
        sigdetni        : in     vl_logic;
        speed_change    : in     vl_logic;
        tx_elec_idle_comp: in     vl_logic;
        tx_pipe_reset   : in     vl_logic;
        txd_ch          : in     vl_logic_vector(43 downto 0);
        txdeemph        : in     vl_logic;
        txdetectrxloopback: in     vl_logic;
        txelecidle      : in     vl_logic;
        txmargin        : in     vl_logic_vector(2 downto 0);
        txswingport     : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        pld_8g_rxpolarity_pipe3_reg: out    vl_logic;
        current_coeff   : out    vl_logic_vector(17 downto 0);
        phystatus       : out    vl_logic;
        polarity_inversion_rx: out    vl_logic;
        rev_loopbk      : out    vl_logic;
        rxd_ch          : out    vl_logic_vector(63 downto 0);
        rxelecidle      : out    vl_logic;
        rxelectricalidle_out: out    vl_logic;
        rxstatus        : out    vl_logic_vector(2 downto 0);
        rxvalid         : out    vl_logic;
        tx_elec_idle_out: out    vl_logic;
        txd             : out    vl_logic_vector(43 downto 0);
        txdetectrx      : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of elec_idle_delay_val : constant is 1;
    attribute mti_svvh_generic_type of error_replace_pad : constant is 1;
    attribute mti_svvh_generic_type of hip_mode : constant is 1;
    attribute mti_svvh_generic_type of ind_error_reporting : constant is 1;
    attribute mti_svvh_generic_type of phystatus_delay_val : constant is 1;
    attribute mti_svvh_generic_type of phystatus_rst_toggle : constant is 1;
    attribute mti_svvh_generic_type of pipe_byte_de_serializer_en : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_a_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_b_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_c_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_d_val : constant is 1;
    attribute mti_svvh_generic_type of rpre_emph_e_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_a_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_b_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_c_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_d_val : constant is 1;
    attribute mti_svvh_generic_type of rvod_sel_e_val : constant is 1;
    attribute mti_svvh_generic_type of rx_pipe_enable : constant is 1;
    attribute mti_svvh_generic_type of rxdetect_bypass : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of tx_pipe_enable : constant is 1;
    attribute mti_svvh_generic_type of txswing : constant is 1;
end twentynm_hssi_pipe_gen1_2;
