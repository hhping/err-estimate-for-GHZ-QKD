`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfG8sPZpfbDPPwCC/Bld9frEiLa0x/Pivu3Uq9mrG66Un/BK9KlErR60g5zR34//
qcOoZSgiIjrqC37BK9Ye1J7SQ7Gfq+mxIURtBtQXFqRnbZZatAjPA5e6O1v69W5N
u7ii2UE1HH3JRJ+gon1MCypOqqmaf14CgUcPumi1JG78wqc3+NIHsVFDfRhc7Au2
/dI9JCqzFlKY/iNSzOzGJ7E5GEuV5TFKrPY819dnraqOKu4NeC2HE4oBpMIOikqf
iusTvHGrrAjB+Y9Ph0PxPg+IiYeX0LifoDX7OGw2FSkSufgtR0zAfrlZBuuXDyXR
1e5eASBZzbP16sHS4L4c4TIhGhM2+Kea9ap1Xyq6OqRpaiI0kPXqLSbECCKFhVNk
IMdkz77rMFnSo3s9tsQFHhaWDcefUIQznFejkFJb18KW7lOIKr3Zw0MC1cjXm9WI
dkbgR0Wp3G6uGBx/dNdk1TcdedwpYikMgv2Q7HYaiQMOvHTlPSdqekbptwursLMT
RiYSmGytmY8N57j0SKrxmlHYVcOlkl/BEf9mKTWSxgce4UHhslpm6HwhP7H7swsH
bdOa95VYeAbi66oZJS1zt77oH4HoDElZL4Dq3Uj/DKTMnuDjAOf6jrTwK3OaHpnH
`protect END_PROTECTED
