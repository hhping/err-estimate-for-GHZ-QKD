`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EY5GySiZjN9e66iwrL48TyDZ0o50AGSeqHFzWJyGbaK143j2GVT72dMX9vmb6lqN
7q7s7mpkCBX0mffjtTBasbh140X87ic5I5I2SFy9/XRUncdIqdkAOJZOyrsS5R5I
KhCk7cN+zJcT6lOSdgKnHiZ/hqRdeqoqi5YdbNetFkMfdHDLpxTZhmB0c1n0DeRC
mCTaxw0XzgN6uN7CSrSpoYmeWlQngTOCJdTgUPkltVSN/aq8zSuIc7M8YZ52ZdRh
GeWPsZ/VMcxARGbk9YcuAR5kICL8/kEiKmiSXTJdNrHx3+ntbVEvix7CTOwxXd2t
B3/XBOVSxdVHl9Y/XhGR9EoCUkRRlQd6tTgOgbr6jX8KmR2y8Pt1DIzzHCRtf9zT
k0qyopCGS57GIpLxuJ6kVB28TMTWL1/AAfCQNeR6qDcYQBIzcMjjfpun8n/4gCfg
8PFsmchOPaDbq4xB5ls+bnIot0llOJbmh+1f6C6tkYhqsKNchQ3jbRjF8kDjfuMi
rAD4pytjhTocWMR9k63nvCCmPKlar0IjoiA+BMz95fc=
`protect END_PROTECTED
