`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccM+ITVjKB8Ywchvcs4lFle4l+TcD4xfaDufspMKcn9lTYCcJobwkidl9R4GzD0J
kqrTdlYb8LaQ2FwE6TCvpNRXSNeqnuvR/s/HsbsVtHOJJvSh7jtcRWYrR1MVI6OV
ZnB4kPu6k6wa7X8yf/bPVnhwMrPgWQwy3Ql9Wgan6qs887dHUObsJR7vSV2vDles
xTwJn9M4068pSUmTUUlooap0wrdGDgEmpvkvdVyTq0AhCInr37lRGkjT0MECYcU5
gp9KCJKThwn1kL49vezv8sIBwzNpjbx/E+eK01kHrtl2LMM7B6mjuBCgWZTWc1yb
5IMpeG5TLlE5UfxC33iU2VUSwxu/8nOrUz2Wu+Tx3WyFGkBvccj8NZDgKQL1UFsB
`protect END_PROTECTED
