`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LleCfZviM7XM1swlRYu3oFoqp1Ef0rRUZUdDyGGgGHIB5YNes38x7B0YGXpBC8eo
stTp0pgs0r3qUgS/PX27RqkukNbOfrsMnOrcljAU5KPqp5ivgFnWc1x6+TReO/h9
O+jhSJJMohcAw5ozmgqrIUKJBN01Qlfj7cVterS2XgnNa30WV77eIL+shUv+53hZ
CdlciQ9zOtGPwipg96REl67anGhne6edj2O1HnkcW7bABFQjdmQ5hGdWxv4b4Ej0
5GSNPDJB3bJWAd5cHqkKFf2yD4XW4fq42bxl60NeC2nmDn7z6lRCZIA9ht8Usl0u
vxYKEP0a1gI2CY2A1ahKQ7b9RfMMapudulHwKk5n8mrPp01oEqcdBlCSpx1y7RR6
YPKCmLVV8aVAdgJQGdxmAk7r1sy+HkITZ6Ex66ZQsFT8OOEqPC/pAk6WQQDvfpC2
fsb9oviZYhCkYq35oZ/8vGJp3aghfkSEc1ZWQG+d4QjOxEmQK0+HoMYOSR9Y6LLf
nOhbrjrP0g+5pgo1R4PFD0wdfFP+jzoyY5AAd+BJ4ka1vC0BDQemoCNCVQsWK3I9
pbuXNA5ikcu2KZu9KMaJL1I6AagbXv1LX4jnCb+4350vb0hdeBfrwwyMBofSRkSC
STL0zEBjqiSrRi3op4ciU2QpPh+J31dv2ZvrF5GyTe8Qm7i3IoGWPYG8OG7H+P5a
Q4Zwq5/AgxdgZfM3GYCyX35PBbc9zqXR6VzPjucQx3XXP4FHQ7VaULlnWgPj54n7
SXBe5xZtUGNr1Hu0bJOO0nRU2HIsaw3dbj8W7HHWRQkzJ5tnOFhKSOj//kcZVB+R
0GECHfQ3ni7xXClf2TMFPvHteSTEOK85atrav5n36yqBlKwHIu6P5CLRGGgaXdWw
tB3TWC/kGJjzj+dyRBCcA02gEbUlXC3JXVCTI2kTBJrawdrzIQNdCOcRxc0Ux24+
Y6bd7CsIJIvonaZ7FS4HkWd1GwrhkT41oF7smi7/naXpKNu0zyYtPscwF/Gb3gtb
RvqK0nXgExUK4MIxXnxK2Sra9Z5ysJ3K53qf33p4ta4QAe+Xc7qOHfdHBFkfvD6a
osfdGzQjLn3MS8vtStV9eTkQkolnWKSUHbXSWF63Pg7AFOL5FYrF9KrKLNfzGpOK
gO3hE/C/cZ1tDlYPEuo+JDnEWt9Rge5gDVw7rAVumTM8PzRcgncOEhwhS3+1A+i7
LFL7XGLzLovUa4g96shj3sp1ZUL9F4YaunpiECek55GZmDtrDofkHDtPUAyxXBvr
fhAvNP//qfcJzb+vUahsSD5DdToyGCRs+UvwTBE45fHG/aZeOMlwnL6k2lJk1dH4
anW6VZzCrV0OXIIp3t7AhZBG0DfF1VlhcokfycKg+0AI9XnoHZljMww0qQE1KTvo
WvwtA7a59hExi8OnRAiP6dUco2GEX5llpdmrrzMzZMV52QvOeAr/jiuN4cuLqfNj
kO/WcHsGdvu+ORE9GrIW58FmvSAq5xWtQLb2d1qbSzUPBNGiJ8DgpZnPa0IgaD6b
1Z4P+aTVHCLxEk21tQ3yUctkPV+P9kIKaObYltYF1KRQ2eebw6d/Y6SYZAJSK28B
RewJtoD6u07hba65W3vb/Xz8MBIK/0NJEWPePzgPviQ7H9hWZmB4rmmsmq8Knbwi
a4iEIv7aGbByfT2k9wTAEBuuzMzlYrM1pySuAkQ+ax/zswXS5m+VMTqJWASxA+Wj
SV23ZG9Vdy2orBJaHvUKfVj9M3ewpcPfO3LNdtvtHSKLA7VU9iShvInBPjrrQUsI
InpLvSslVfExPVlI4vos0AMby70GbPpbFYtxARu3GyQcHM8PkR7Z1nkusWf/n2Ql
7nUPUUUKXaGCTVbT8qxj6fE9lUB3ZuEKe31PyfcVTvayHN3RMs0Ek7jKbEJJm/MX
jsd+eTIozpH9lLYJC8ll6/XTGwl8xU5BH0ExRN09b3OfTdZ1uUNZFHao2rl/3x1/
yTb3l5vkKSVbXuDm2hlje+RL4kwKEfGndk9Cz6TcFR5yjTwQGmhbSXO/RBdvt1LP
N0ZZjaWtg+P3wIZvQBtISLfEtP9jL98ENeRBfR6Udr2vRr/O8P+UwplQFJOO8Zsz
VX93473aCF3wYw/izVOmFaPW6OqnmfkDDugdp5bkW59X2sKnpnww0g7tGCtXanEp
FUX12pOH4QNNVAp5Ea0z4Pu+t9WyQlcrseoryECAzsZs1SlyG+nlJm1I/lNSg3w1
BUeFVMtv4BZQC4OY83wdYf6lNy20OVpJPquEsSOTyM2PM+Ml2j6nPo+LYtD1ClEB
d8HWSvoAQ2L5VWHs+oOIwiJuvy59nOZ7UJB2131RrZwiTktGQus7LGsi5eEZufgA
0TXUPT2VQXRaaepcuN6FSiCT8kAuJmYq9SS8t1z2TJfnbxah2dqtYsBrRyBC1I2J
rYp/C+seCM+WI0iUWkNXw+awcIAdw535dsNz1C5cGvAi4CflBHpH2keQY4NOILaL
snRBDB9yHJJn2U/yF1JBJskAMx4iR62tM/32XzY41zCEne4SbF4rkSEBnPdN44EO
YdTUZCOGFb4HgXWTJV8+qDtWWwkJyed/51tWLAImktPybi0+FH3dVdpcq9ElSLJW
eprZxlff5qp0OpGYq4nErg2HPAvQmdRd78S+YgfhkZTRBYirbVfnp8mTjnWZnpuC
nxauw94J4dk/Vw1+C3/aA4elOq7NSa1uMb5O5SJ8OgD6wWITLgrEbr62hL/UmXm1
AEZWKo1e4qjB/kp+vwsfd+nXuN5GmuFgw/wzsp9vOi6GAXqFpe/IX2XS5Rq32lhc
fA3YRyIi7XKsihJhTOYF5RKNR9Kilm5j8jvK994oIZL89hr/Y27oPS27S5+34/ua
Zov5I0v0mUjfudNaNHvwX0wKaMeE+OyMmJRS+29g0d5hB+Pzvg8ngo2vmyAFTCzs
xwVejC/GBKKGi3qPC2tWXtUwMLAb7v9FeMLstpQnHK32B7RBTzgCI5JOjTXP5Now
ufGoJSSbGUZLADhywdUwFQDW0XbzvBu+eEZQP5nWrU0P5ue5nETNi2SicVvP7fAa
aD3acN4933ztk4rO5rIAP2nxB885F9XJUflXAOe185H1OjtDq9zvudl9KH1lNbx7
ahwRgLP/5I+CtkrgI2j1O0yYAkJDQQkZVcFG2pq7a1AU4Gkl1El8xo7UwExhBIUH
ptzU93hQiesQityS3ICQzLT48w+jmKIK980pLubxD6rpZVlIToZfsNvkYdtVwpCj
Ojb3VBMvekqB0ZI53rAamMM6YXBFFJluEYHA2qBkY5SjML5dJfDMtfXEOa79jtzw
hG7cGS9ELQR24S8RHFvWu4Lf1gRobScFgsm80My/PGDv20yE4JTT3caMyP5xylLH
ETqymXTaeXW3lAAuUhGjh6yOavo7hYH1Ls8+jjjz7Kj+Bb81Grr8tGixCaz3nMiO
4O1LHbqvz/3RxNP2BtIiRnip7htPGaPhsc4926V17elj37eq/LbNtpFe7XUuJJWJ
0+DqcjGA1KBDlYvl6o1ezv5JGnrVE6AVCHsL/XzHOeOWgGZVb9hZeW0HWttcxmfx
wlkn9FI5WZe50G3nMhTIotyKW/XX+MOi8rmOIn2RZ/D1KT8ZEHHBrchUidJvTrkh
/6LRi78GMPb/8fTQveP3n5MDT8+TtIWSfzCMw3hD+DBRGUc1At8PDFsn+N1GQs3N
9GQq9033fxZtEBVump1B7R1WSZa7dJ/Odlt8CNknNql8fKT3mjdq9fgzDjLcwO7y
vZ6dl7kmF6Dv9+vyCbX0p2rNCO09J2Pu5GopIyvG+Sg0Sv3dcILj3gZhR0aVpj3a
KuTRFdCO+GmrbHlZ2gfy7J5iAPXoHQYSwwCdG60f2/ZHm2bPsutD5zgIRLuKU5z4
UFNIXfJdeAu32YmuBgoB4Tu6cVV7stGA1l4VsDUeP06pvaMotqyxQIxDgZ/HgczN
2kpTJwNowig4qz8iU+QwRQLvHcWRO0dPLUEIkYbE9KLguRzudVDyqPsZiJ5aLxDg
swaKMLGKt1BmMMYxOU89HJCV8RroNyTcN1fI4GvG1Um5zT2mOZ08MxBC01+y0JsX
ghBWZmqKDicqr8IR3Mw7fyS9FNH6JjCYBCs3LryIkt/6ffFpAgF49KN/MvR7vyZa
PJuwbWoMGMLnNoz5P9iGQ37NuAZE+6L+/E4YKhr/ajjr+cgJKQdQH0GDaSp624M/
I7IW5P+lN0VsfXupKsGGCGYPgtceIUTCeDpLOvB2Bp2cTK0iT26JCQnWCG+gfg5R
4JJnYv2NOxkwdFu8dblV2OxeIaFb3ozrwoZYTKub6RHr13kh6ePaUJzMGboyW7lY
cdIt8YvkirEZxDcskVvrsDTQcI+Rt3cuLd2ByYEUYVk8xj5O5e45NJEa1nLebH7v
NOULEiUZhY8+PLL/YyFE8BN9QOJFxdnYCLyzXX5vHBZoxX84sJdkZfpQHxa7y0q+
bGQKd7AnTI0qxcWi/3iOtFG3mQLYMVW+vRMjUbMgHGESITgBRydqmG1V6zFJCgu5
NUCF1ltPO364rpBHfTflVWOp00ytY/D/p3jwq/3QOGgkwJf06NKiuiRJLJpXCnZ1
Vw+aPycPCvj0VPwFCGsq1pWmn6PqdVdbL0128G6E/3J17gXkcvINUKwNGXTJws9k
BdDGchaTKEVsLDdRZwWAFFv+YdPspvF3vKBzuucBgeqvAkjarx4ImC9al95j9Jwz
k6APkBsmpx6lZD0eJ2nAcnPvN6rA7exMWA4zRsAjErpJjd1N07G7mrHwBgBhqBYq
V82h5slHcrzok4NqD7fu1tG6jFU8QlEc/mNDGL/Ar5yFb/LzLNsJTmcQ2Wf3dD1N
UdsgbpBI8KH0B764CnhUP6OCjE1YUdgRXUo/qXSY5wajA945pYi5wuYy5NHy0JJf
GPhxg54tEQjXEnvVZg7SdL3bzWsOv0o5LYUPyzuTGdLG6Qv0EuPC+s8I543HWijF
ISO5yjToN0UIN+VUJRiyYMCniq5Eqwa6KTddfjXaCQkBdGRVDO2U4frBf5YcXwLJ
7A0Z23QkWabro2TWXiBvJHnJ418HjYIuv2m+0LLM3SDgLbedulR24RIo+1VlgzDW
cio3Cd45lq/jKK6Uw9f43xcxgoQTPqu6diGKj7TqdvuQtrZm9tJeTGRk9RgY+gd9
njBjQfA0SiEvtN7U63I1ZZ7o/n6+cNnPWQdtCi/OGhoYBE8dkK1FNRWJkUYD6pwz
khYSbx7HZhs56wg+khYizNm0M+UBOyFKPBVAYumylpbV1PXkLqbJMY43QEBubMrK
EYFf0fUYun1ADNMCwL2YcKISlr+IGxjvT4Lq197LYxuY+CRmM8GfrQP57CKEohLr
kmevi1ydAsMmPrXNXjXQF2luJSguwUKpQB5Xyif2nltLMw6AgXE41nXpOeUJlD5G
OWUcaehSfre4QfGfuQOekG4JRkJ6aef8zVvxu5W/ME8XLl53rHDEj4MLOnDY2WzP
Lq3HtnMRFG6S/UflZ6Vhaav+SNAbbZeIxDgv3b6cRBJ3paiD0IkZ+eDaGZUjkG15
f2CimawJeYpcJ1b5KgMbk1OiRYjigc0lRAu88lpKoPkda2+Ne4IQrYjHuwj5XBB4
PQOaSRXUPzHQVzX+qdY6OY84uFIzG/o2lwIr33xlqqBWeqfvz6/N0JGZTvDni4c8
0c1qKJfg4olRodq3vwWhgVWlnw+64HZReWT02wnbs7T1ussEf/V722dAhoOFTr56
v43nLrLYZwrqL2MEamkS8r5/LZ1dklyYRreakeOtKEzkqRmw4IFFRpjSZ99zym95
xczm5Iv1iSLvm9J+TvDELbO1akugdCZAxutlehYkreyRuK84yayWxAKEe6uOcYD8
E81D4Qh5vJ6NdDZkWQiGBwE6VZEvs70VTi2BhIeo3e3+aNZHJhu7zgkoLJ09Dna5
3P8tKAuh7cgcGluKY7TEiLtmAn0fwPApX+tj4B4rFp+tbiqVw9eeFJ/Ki0sMCkIT
BhHWwFfCf5ztfDeCdM3BZ6uhN2NcoZUQuAtFV0ElHdiUmu8cPH33W62XVYFrZ2Pa
9DMUDfZxyvvGuO66WHbyZl+Ycuz5tIF+swcgx/Z4vpwnWiKu74eCGsk0XoKPxBlp
a03MHIsmoEspM1oJE/xgRUkHh3i5DKNh3zA7n3qBOlQ8xnlzklQlhx0QriLznizY
xhpnQf91xi4keR93FKSbPUxkKLDuQ4bAf1u9MoPkIyuLIfN64BSpxaQUwtyzxbCM
B9bp9766tOtuCX/egOdIwvVgifCYnBOa6i3TDc5xtocRn24+ausH1KdvjUs7+h6X
l0xqnqa3V9a5N/XoaCk/+v5MGHVgF1U2iynHtrqd0QmB0gCMbZ+hIXeppuTaDxvQ
iHYOY8EazlwlZNhvsxT+yeKtml/DtX4ldMCwG3wDT2w9JWmtP+ORLXIqCq+K24uH
qWq9e4ep1uB0Y48HBurjoD3dZ6iuTRpuMkTrkAQhDyT7POyPxmcN/xIn4tqrlgv2
zCQQipQJGfLuhHOXxcEbajggE+Gh6at9nfKzRSMazEWj91dEZpq5zp2IHSisXLXi
FCK5BsN5Qzyml4+p0UGK5jiX/fpug8mHwUKbp5ylWjCNU8OBfHQaML29D9jpj0q9
KakfiqcBwLvOSJzVEWfx+idMAK3G73rCKJOiK7E9BJuXsHaMUMt/0vb1G5KmAG1H
USMDDHdp1ypU8Ah5eTShrKMHeE3gQCyN9NPJkKq2zP3NTVU0v9IRqGbLP/p+sL7S
xv9zjEeVdXjZzn37umA9obP35+AKUJe8eODjgx64KYb1usOC9DjcHqE02afA98/g
NwDHg5a3y38WXxtPGgRsnMBaWQ/BL+88gpVd+bAuIzOOF2hz/Lz17h5cWbL+/lSC
EH+/3q3tqMexAqyCDQqGC5tOT6UzuD8oAn0m8Se/fnZE7L48cH9x5tOBBxc2a3z1
H6vsLQDeQvROq6OttVTYRkwINeNGejDQ5pIEcq1onzrRm1drjo+/OvmVJB4zMJZs
fOxGjd8Nn+s9fXlnoZt1ngigZolWkT8FTsj+MYEgsW/Rfoea05Urbm/55Qrl0uh0
as8iutWOZKLgR7XYEBY6HYaUuOvguD2uqY4lXsZ+iZQs3YbeiXyzkyo1HaIvnKtb
URlEzOreMEf7Phh7BapjT6KrIuhmHwN1uDgJxRxQAhuHLyGgq4tMA+/XzmbUbiyR
H6MXuI++ZCz4IOQhj4cQ88MP/6O0ajG8ug4WBqa6QnwOVPYmhnJh7qUrudk+tcyT
8naoRJI6UuNTbBQcNXbhUjJ2n/6Iier+9K59MapUpW+L4r3YLN0vwburKsd7vqjr
smX0t4YOisYkCWaKM7czk/0XIdhRnJgvXn062THLg6VaKrjB519HCKaJ2p56c3m+
c7rkGCsg1jSPwtGvxR41dbyxvkRbx/znJZnG4fp58hk6ExuV2i8/7ov5KPhI1W8P
F14Z0EU1e3qWgDeRyK4Bh+9Cf2ALZDMjfZqI4eOsnBgSX7JD+MzMqNa0rRy//I7Z
pQNHqZLNQAMGblvTQNd1/WRi4FbcxucR2UItBxnNmws7UNQtmk33lO5R4Y286t+M
O0x5EhL+1IJxh7eVTfkY1Pin4a8KdO0ITkrN4TtSO9iI4+WohJ3UCjVayZpi6xlD
8xZJd0RiviEwf5r37JWRdqlvRYyCdfKkdzTK35/ukiiwJrBcuNU5tatN5xj14KUl
eEEnqYYi53KhYMhaJTvVTqh2bhQGajjThzSAK0CVqM2dkVE1Ukv+Dg9BToaRpDBA
tnXxOQntzvCbv8H38Z9wO4azEJNhfDqnqlUL34J3rUXs6rd4/gdEVPYFrT8vW6M/
y9TM4C+XH+xPogPxTNTNEF/5szk9Ki9C1gX+KmuDonGjXA7HkIrMiPD9bwafAl8y
BKY8shuzRfNb+/HvxQmCM3SZSFppx1nHSnzADCsb1DtYUW695E5IQ1Dn5KFJYi9O
/JKGmqCu0UUWbTaAD/LQRQ9E/XiJtkulbuHU+XlBZ/bAuiIBSI5YwBqrZDETeRJ/
X2WpFBxGnwumWCDRE7KmPD6rHL2rAdhmiZymj050N9cMb4ujPRec/mfU+1R6CAG3
5Xbqh1NWcAL4YNInMy+h4M+LGu5c1iBTxWpsrOEvjMho68w1Q0dYb40qyAFhRwhw
vyq2XLGhcQdOAyzEOGZdwUhM02dNe72YrgQffL4M0a/ZJGV357Z+aMrETMUaEuCC
vztk/wOVoNQVynk5n8umGD8Aq3MoMCUo6speyLi0P5GewAEkVdIke7NlTQmVFSMy
c8oQ8SRi4QHG7CX/ismVNzKR4hSGYRJnQwSrqrFsMad8PjzxiZ0TfrZo8afbVi9I
88DiusGobB7Y8wL8sD1sq6KxRIv6cUByqTJyEIf6XCyOe1qM3grlDumAheHv+SzP
dedJTZLciK0H9DDvx9VV+1KDT0YOsxWIOVC+ehqJOtTKlRwODqqsx/sQPgwY7pAW
9+Gc//q9frgiP4uQyOmfm+F8p0SoQDKCw1ReJZUBKx6hHvHpxLG/NrYnMX8D13xW
WvhMRbekwQVU6nbsgEEa98s44Kmfnged7WkL0aZi2SEa3mz6rbJwW7Pq3+m68PMY
lTPQ+rG1UzFAwIfV8+23QXtoIkywfbKH9Mx/hlCCPKpR3x4lw2L58Gx8DXIHzTZB
8qrUKehFE+V6Ou3kk3ZoPj1rpQszCQB+eXKT2dsusgOmrRUqCDze/3qOetBa3K6c
R2DJL4Y+sNHeqkXNdTz9aohFmUg6dwo9cvJ+X+f95/zbYbwR0OcqAdElCNr1P77B
K/lcdeIW8DNbt3FJqIKkK1pCEMzonXlzOdYWuSQUypt2/awl6/wUFvRgvZK/Z1ik
YO8reCwpSmrx/kKn2mJWXKYUF3DuBB5FdUktGpb//Xen03EaKa4ZJ3Rwxt0wLOMF
ZiluCFFlbRGsZOhoSrrwilekq5l+BJWFAqiSt4PZi7sO/ia9U28UHYLuIC8PBjuD
Os5fmPuA0nZjaqKNsMLJITTpbVGr95kZPxHDQFLFe6MkJAJIe7WW1VE4WR4hE9ix
GuWe3PeH+sQXX9YY8AAUSlmdyEhM6/Exzk9c1d0riAsvQq5blttkSvWLZxlRBOt4
KJMb3H9buCzNWGPl9VuBmNgw41HUdo/K5g129YedeWLhPbOE+D98WaI/nxSKFYLB
TfWoZaxDvHbZePjWK3qwPXDGY4Woa+n7Avb5p/u5rRuzlB2KMiDV0jMznPiTfs3D
hZ5u1b1J5WUXjI8msfkmjt2aNti9LLpd2xAZY/K/XQftZpwh43OVTaaC8oV9ohHI
Wfk/McCnw8O/D9UKD66XCoWU6vpNs9mHBFYJBQujiaOEWqSLxmgVttgX//0Pq5pm
igYqKXeu8iEAOP+vHKwm7Zo/IWvc/J24cIxlvymA+GHxHW+Hc9Bw2e9rYg71S56A
8RmviPBoey+pU/4Bh8yEDQD/ObB8Rs5TW8pJZZoV+tnmNu0ttfCW69iO15AO9rT5
U4Po5JUyfaqtFk8V9dOo/jrszfZv25thIHkbGUtC61KDwzR0xBF7UNQTzKmzsLOF
3oponR+Kv5SktJU4luYaso/32d1zeT9s/emrqc5xw6m6cgwll8H2zuaVmlVZlgpR
eqhjuUuvYg0vs7QUpd12sw+4EQSnfP1LoipVNPXvRbUlS11OV0JDvsCGks+nvrIP
gPU0WSh5ZRs8eeCJhsdwsZ8ZfBn346SjQgIXYb458m73k4zYBGC6Ow+LLEQiat+S
lclOtnAUWTROcth2qsQ+DfPaQhYu6DokP5/X+p0xgMgj8VuP0/cnpyb5w482FQhh
8LpK4yS9i18IAB7a7IE/iNMMkbyn+E8Sj36qJu5MdSAjHZSFLC0p+ihzmKixGcpq
aT5L67/oQQVJaCI5GVYW6SdbJtDDBdusyk9eFFQKsJD41yGJ1lyX7j+XwOrX9Qp3
vrk4gIwFgZT1oBMQAyDwQo/4kE8w62ZDpJPGgyPvpOJjEYrLd+C4tiWAev0+GOdx
5ytm9dPPTs54pAhQV44gZ2rPJ1I9uIbg5lf7qftko9aAM/0iAMUoGnEGgxM1J5zH
N5xhl82r4JlTeGe0UNBWMESFfBnMc1y6VS3OO57zKtKkuCYEWRvh1attMC6D8EGA
Q/LJftQDG5VX9NPe0G+a19fGAuROOyC82PQa666Me3Ybm54qHv/EfY545Ls8O8h2
LlouLK9dlEkCYbyF2bYlTu7R3XC1RozDmbkE+iKzANJwnrMIS1QbtCOMUV9hNJCb
fiI51Kf6kmrApg7kasfbKAsDH52Tf2VLLOimrR5IhxJfdRhhxGyDp4fhqgnyXP5U
BMzug+84oRvw1GG4WccnZz8sNaD9ufLsVBN+odK59V82vUFpbst+7mB72ovRXhXk
6dLooNok3fbZ6QYg83gvgj1KDowasiMEYo5fynO/gjvewE0XzElb0qo/1xlE4Bab
nfyzxMCQ0P6lF7a4HGE/5bRYhDcpU8ORGV9xDR0h+KrwPTbBaxCVob/aFbZDhi7C
79+m+vqFVs7OSe4YxVWfdoBaWrm0zctKcWPgs4O2DJliZcL1uEQPXHd0nuxwqrD8
IIXqaZooXdk7/2YEuovsW3i5aI130dSHL9kYzw87gm4OpNii99TyYo+VWpMMCSFX
dCG1jlJ02D8TIe2RsAEqDWP8Tn10fQTCQk50txd/wdGL2I6e3vDEcySjJM4hTArr
IRUnh4aAXTyXqIEBooi/nfJbsm8qU+R/DLnUGSpqGnwQ4WEDpKXjD46BSkTeaTa9
n7pnSEvJGQoWAu8t0rlrguB4M8uDlqF27qFfGuOHvY6t4FHEydkVFMykQm3p4R5D
cjXOCNnm/Ngkjuv/FHg+3fAJpCWvKIx1/Fo4w8Kk4VpU0zCYZEKeM94zNLlJ/jiH
YY+h9O3tRfKyHihCkfnsht5Ma61gPQe2jebn2XV/cYgQZCyxwwhe56xl/uC4X5rc
hfYbrDmLdf2ORBOFfYVXGoy1FlUjhLaS+0z2BZ3UUSrGqJ3zvLOUKGiXwryfccJc
lIPbYbzYJ8Sf8mRRu0SmpqemzmOBFH/Gg4OcCwLR+TRXhtKSP0RI/x4HstX+csoa
+J2haeqldXMuxIXIZx4NyvYF8b7hk1y6JeV3EoVNs5WtJ+auWncOGQlgACSGHcT3
qm4eJZNRnhmqYN5FzQTZtmJnSirX25B6N3wLciuapc/jQ29KH148IW2U1JPY0Cq6
4e6sRZkyOHDp+bbStCELIJLEe+yn06e90ICCSZyrRgU8+LNrnmfWrPN5mFXI2YAJ
hCq/UR5Iq5OKrl2Q9TdNYBEPZQo3Pfp0nfHmyRMDAj5BTI8wHXksYT3GSi45nPmI
UtwpAWfGcAyfAa5bs1OJ2E/Rubujlm1ab7Yj8gPBjbKM23/F/YUo6IeqRg1b158q
2RGsmMZfZ+1PecOlH6x6fQlyKF2Q+f0au2Tc09HbDYUpGaZaAN+f8i9YfxAM4icl
xKAyO0Ii3cBrS/rl/GCSfEVV1DTQ4U3As928LDEkM+csnkcwxt2fNmTK+s2GdLPg
N+1YUCxD+dTLAKgBtGH3I1zi1RLUgnXg02xd0+1jzBECrnIKM/jqpUrtsB6ycGVu
eOBM0JPOiiXhmOsei3iPED8eoYlmDjaHPvSWCwFdycWzBgpKJQrLhGkaBU4HVVgK
v3IbRYGkdoHrZheycMO31py8pWQI0h32+i+CI7TWtxET3G5V8KISxWC+o/79bahF
hqcDRh9+7mvyLlbZ1sXRq0M0Re4sb/jFZ+E2SBHE5TvB7BcvksmxHIxyQSRWofuF
Uqzcdf6uNT4Pshv+/jAObkR7VfS7txq2flXmQ1puJow1AWN5ht5v5JzQa7Bu7yJF
xhranjBwEuf+63i1rIk3GDLerMbSgmdu8+kgZdxsGPCmARJorq2grGRRfwBZCdjC
3Ir+MdqZBTAiannpt863iIuotBpmQc0XTdMgHNplgGnSH6aDceHtDCvfRhlFo0e6
Wwp/JPq5nBttatN+bE0bSNrvlPddTNO2U2Zn3DDl/FGbZAuX13tKjoST2DAqsaRq
Nuy/aYtQqUHPWedfIx9OjidF312GNxqQR0njzoUoq+1Je5gqgV3OokbssmpVFQ7j
aVeP1tyxP2lUvypcTOOOA6woWUV3RIh4SWPrLcPfwK0TVUARqhCkOiHc8XBK83hL
Sca+Iz3ST1Ar1F5vh7OiSMlRpesov/e/0e2uaEuEj/uaa2KhC+NXcT+YnEV1W453
ihKjbmIa6/NNVKMAdG8gCZ7pNbbcbKj7IIdOm4Hs2Njz6bgtLBwcTcFq5z0IE8OU
s40x0BI9QvqYUqZD/ACbQeV0Dj4sdZxKxLzCMjsWiJc9RIn444wbN9o6M2EeRubZ
UU0fkqA1NKCZWpLekYHg8FNBDHLHWi1ZWaBd9c5cAaWOo5Odw8iRgz4Hr9eVIcPi
lagQYLnHL+AGSpG/tTMSir8Mi3MhEBAiF/idUqzQ3Ajv93K1xPjtWBbNdgynpVRk
9Mdif9PFcOpsIrBjgNpk2CQdolug1MFRK0KPHk5w6/kBOM4uK4OL2+1Bh/RTQ9dZ
MNGUPWHJRqwZG4xpwu06TtgVlxwdwIk8VYB3G4sHQSh2JulJgXj6I3BUiBqvPcDx
ceRjJjjhLqDBZMMOw0BerLhTOHaRdgFsIawa5L8+mtL6z+SwrGIMJNihh8TmmtDM
f7fU/2jiZXUmPFMHb3/qeA1azbdQEwT2IOprVNZnJ3p8Ueax6jyLbkOXpHuU/waU
8Vg0tZk1bfEXzBlHuHYQBQrBOoTTSjJ/suNQzQlp/eyJW1UKJ/dSvCJnnCQAKNbu
kpbTTqmDJbKJKu22LZb7SlN4Sh2SBXz6UlOTLMAdmKeBfzSjRelrO7IHj+7ni5ly
M2GCwF7XsUBBHJVBk9jkFYAtgyYtYNchUq8dVxekQnVGQjAdDH9JQS8vsRXGo9dd
eSSn88ialWl7dKyY/e1iUxeb6wWb6M4Z+R8DI7bBwlpnK0IX1ybmjkDM2Zp9/I34
iBISGwrFgBA747CbpGiOdUui9Th+su5h5qDbQE5rj9iOy1jPGLmO3Sd6ufecK7A8
g8d5tFl3j61QToh0r+SnU5thLSRGWI/FRPqRFprJ2rSkH6TlCVovXiUUGho2Xrvy
KeUeU9AONFky35L0/4PO1spFQEIVhEqA+JxZJl660OvGfjpIxcNK9kwU0+OBsVyo
NjzcOuGKxNLewhrtHul7Mim037ST3KpTe+1Mnf8nnqEqFEtJ8Qwr4qhAmYGJKpHm
9ccwuZr+duRLMlmohbGYuYVOpOFMzITC3quvmmOtRnYTn17PufNL7XMo9ZU2+RVV
afMYzyHqQKv4X7z0253SZ3wIwKfoCXUoDQspy1+mU9wxKzXKnPdY8bK3kWsYvPtO
yvFof01Q5oVpK7drqEnxJkk6hDlvro6J4PsoWHcVJmovJ7TqlMHEI8H4qVU3uxGs
whXRAU+0y6Z1NGi+sFDeTdvcPciAH+X/HcXIl+5xUGQa5LBYjZ62FLUcvsAiiugt
X9uKQ2Tj8rQvgUPLauwO6NNlSZD0oex+akPRsvYucnOk9zMdNGy7WbKJlf+vSZC8
I8yfzFUwZBXJgO/WBlPTpqo9rK/XJX6sJRaIwXR/vHtTo4qI4czP36IPOIemGV4p
uBWdMIEpMmoGjn6sBF5gqVH2pLLg/fPDKuJT8zG0twv1i+pOCw7NQHvkUMnvw8rl
pvtlKa/Ie/Mp8U9XHHyROCz/tb8hy0SiH3r0SPpXY9pkDFRvy7GNKgeiQReVQV52
a4jFuAjZLeCSePPM2oKfkVfCPmdPZcZCg9S6MHE6QAZZ5SqO16OPmoUR7MrXZVQ6
VJ7i9rKwQWwd7qEE6ctsrV6CPGL8Btg4ccTEwkXF3Jlq3TKBJTLvywLKZECwJmmg
hGNi1hRcEHgXO76MjA0zSj8HRnMMFoW9wgToBq1OGhFA385H8QI6KBDn1gQXRg+r
mLtyAiDP9lM3bJivkMmEngqk9v4caQ63oYhMCIEPU7/jG08aYFo6tWL16TX2m/cO
Q3lyNF4rhI8AoxycC7OQg+2fdCsfpJe58E3wGOCX2BJTH5YkLibyl8mru+jl6RoD
vCdSdVSK65KXw64BNuaW7ADf1JMVODsqoUQsjjee3JKSfQKjujuRSMKIBcr6tKAs
ZwDwYdNJo5hSz24IeNAILskO2+sZRqGJvyEkmL2su/QfqwEMmjCsdKkGkzfm+tmY
t9E2Bv6SUes3VF/7iG+6+OvXUWyL2Sk0bORagPMrS2ASK6qLwBi5b+PukhvzI+Ds
3zDesuQXU7UwN7LaapFz0rUvTklucvzGjddQLZ7n5vIUZ6QVwSMfXDHIdAZE3Rt9
IPaeO6e4gr4rwJbOHzLDheYy33uSgDMJG2okMWmNgDsxTLGlUeFE/CIemnJ47hMM
3EFj7zHdrKIAH+6sn8QCY3DxnC4I92MR6PB7JUwfnDy7HJx70YwW7v4F3MeSWNBr
T40ANPrCmiiQrRCdV8p7h5RZiMRLLicCKdUZE/c+PeTxyFTzseYCKRwyyxRbNaAY
t0bi9pqXFYE/25MDbaA8bN4dp3wNpeQix6QJ/hbHN1BUSWNMuaA8VQfX/vkgcyWl
1hzOa9OesxukzHpurcCQ9KVvOywrvbZHsljW5EmWKxPHiqSE70Fg9rA42o6dK9cb
qdo29GAR8c5ZxqpIZhQ7PjYPx+qrLB2G2vF8mJe30mzJ+xIOh6V0K/3Nul1YvrwU
DhFuz9OfYrNEvjjYxaDkzVqBVQ8rwl8LTQUSMLsYeMuLKvuPcO7fwUm4bXg7RxrK
X4V0skUaraz3kIieLISQP78zH2DJ46tkavgQjafDdsBhSKXfyJ0eJr8KGtfZlag6
zKTbzygQVQFCFEYNpOdzijMenD9GsoLYdgpgSSjHu8mTr4ahguwPAoQk1RRzi3RG
yFFZkdfoiwt/Dc4QKfjlhNz3LgcLLZ0JXt3pSjrINzYGjWnQ8ouP/8MpUhfwNon7
w6k+EbMEPmlgVBtMnLtdsiyYsePh1Sre8QR868wnrydkgebzVIoR9hwXi+B9ths9
7nKcnc08FFy0MX/kFb4CsCnhStcWBwIQiiM3xtkBAXDs80IVyOCc/ORhpr2pjfvq
sAqgm6ueGJQjeuZY+V12DNjd1FRWHf/QebCNqAeXXG7ozWRzf5nv+hLnHvqIin24
E6tKThXx+HNz0YFwo4Atos8URgWsl2Zf6oAHjbANothUSvBsWyAS8HRgu0uhcZ1B
33cKr0ASIbwY16GWYI4Gc9/wagtUfYdh7Uq8V+RiaBS1Kpof/Cum+nz05b6xn6Ww
6oxTsVGYw4KHtnx/GFAJgPB+iD9V7WxutA2NWZzDFT7ood0aoJu9Re+niOa5ztix
oDcQffhuTVvk2ES4pkhT3HZ2pxH3RWyGfw7yLJ5rZVY9Pc7snGNLQpJeacTKL++A
5UXKPDxGzujRBlYGo+/PoKx6dabbUACORfjulowcihSuHM8JLvddTuUC29NhtZBJ
Vm1zsAGKAbUoN5860tGU3f9uuo7XSZqz+/q4Ymz5XUWSUz/clR9EDdCe1gP1E9v+
NV/cMB4PuelcSZo/CGyv/sneLNDDx6NeGv3MvufKi+2WAUIxORTs2JP3SkkqdHlb
8Nb7pesABpvwda4+9FwUd2y/f5MB/pAVdT0GCcjVbztK5iptQxHwAMbn3t1bQv0w
1JLaxgqde3X8c0wb31usSmZvks1Rgrx6KV0nUK1NADLpbhs/hBINzvbquj4wQrh5
yfGHTAN4psoUoS8Hl9fkFjmq28tCdNV6fA35WHOQxDCg1hg2h8Ptk0h16TLBkPVn
1+bFQAPOxYDHHVMb8Wf5/Nzz3VV0qzdv8P1Uz8cp2znkU3A8VLnl6Vb00oI6aaVc
s4kehNeFomaibdb2W319ABNFhioR3MbH6/y+rraNcq9rxM6ZXZbhkfZPsF2L13oI
u7fvxYPrvoW4Q03ebCMP14tS9AsJORzgM5jjdbgS3JYVOyZ1Fwolm4kJpIPPKrjX
+INzJS0hZE1pgIuxwWrJOXKmggkS9yWMmc5GCgXOiGimVByir1I0jqJ0281JhQE/
fUuXTm5GHGRiROPQ0ppZvQDVQhIHQT5GHrz84FHEITTcc4LXSbUyBdVOvo+MEYDW
pHUL/8UkYxTiyZbfBDgkaRMlkBvW4ZWIKYXG7QDgDfZvKJryDDMCzaz6jZflM2YJ
Sjkq65PQNhdyueQSBp9YYpc/5rrVi0VG20qxdIe18etq9kzedRDGbc8sadcP7KIL
jWI2kfUO6xcw+LUdm7/KS/yxSzf3mqTM0TKkK+xp/XXJd85Yq41SHH5aYeWBk8WY
X1dp1J9NsTbVd2XjrtKgcnyTv7PjiSaNYaqVwunNs4a2brbZkJj9mhTmCcAd8gzz
PqEr9w6ipOufo6kbjxvSeRfAoZfXzXGzhJmI8hEoWJSZPvsvpEqZXsd2LxZSi2W6
BI6cnm0Zi/SG9d+QbBuZC5NCfv3HzHD5v4FH4I//6M3on335du2nyVoJNV5PPY2w
G7PveFk63nxVzi6Mrcgpxmv/uWk4MtmPl+xrE27/OEEfu8e/hFCMflET7RC+7PK8
I9IILPBL9l0fQvCkTfu8Uc4hcnTeXY036GRQfiqOavFEs1k3f6u4mm+phISMJmLi
FeGK5H+qoLLhrZuLnQE6mEGvyFlWq1DfUd2LiDT35eGKkn08D/bKVgCRsdURMOT+
7M1+JclGLqVNbTzxx0naOB0RJe757p1b1CSArkvV86eZYL4/O87IPgDUiCGstPWV
kR9nuFcMgAprqKfl0YhREeF5loyuZwAwKV8JnbmrPsx/dIfTTd5cxvODWp/Qjull
OZEyJDi0Do2xgJ9k3BuG1CZ1ZDMc5sdnKInHfVc6hYSo0d0eG5c0p1ZFZWZI9jg1
L/KxwR8QJ8NcVQYWhGCp9SKKtVra2SK20lve8ZW6/Daa6syRp34lj5kADenicf46
+6NTBdLNwzciCZ1ZnTwlA8hZCXiZAT6QanJM9lo0NNlAay0ywoHI4y5He/URsQk9
kQZKKnzyUd//UEuEBZ/7JvfVd1/XxR67jhHH8ce4kqYKj7G98AOKaloylU2X7NdG
i8EwcbuX+4HA70wGQVImWTjSD8a5/fnblLyFMopdFFdl7BwX4N41TEoXzFGN+WY5
NujLoDcjcapijZS48+lOJIzkRDB1RNvL2pNVlXgNnG760Ss184oY4un9uk/7t3tZ
ZnnCQIjZ62AowXG88vrut+Wl0NBcfvZW2Y+9TEMud+ylmylpmnPNUZRJes4PerZA
Yab5T5axaj7ReTKw5BagCBYA5yADhewzJVLyfb3zpUIgsehM1/nBMYGdR9kK/5Vv
tv9IDyATlr0kPi8n5SJEWlLJKnSwaABNN3gwGMJOaucZ+jHHgfJ2YeKihY13D5IR
i4qrakMl60MittExAOV+8DWdtOKVkN1EfWPVcMHfPv+Qki4tLsEE33YdrHV6h8ZO
ZOI/RpFicXs2mzpjm9b06RGc4uEOvwhMWb9SE6iKKA77e9P7ZorRKAAydsvXNMG2
CZ6hSrOHxTU6cZRv52DRo6Gd5PQJswUuG1zGUM95TomjZRykOX9vJJy+KaqLvYQO
1T+ufMNx0qyrC9D2nPqo1zt7bRKzWEGt1tqr2dM+1XZkL2/4UIUoJw7KlaIjX+FW
B5ZXcT8VTtO8LRaao0EYl3i4exIziUXuwrRUEqW7UPHycQmIfmqjVtXC6eF0YJ9q
ozZ7WE8dqpqO066mWHyl/u85cMN32Ob4nHP8E6b49bC/evFp+3mYkHurh3mXBUkN
BGEUeiN7nz4AKYqq53367YYguyBTfRWq+G/1xgsY04rczs8PIWRG3ekadxsqrHQl
wiF6Q44a7ESqwqH8GGdJqvrd5bCqlPBKl+BxcrLXAx5/LAqsulIyHdE9ylazHglz
3LtQ9+YaodRRmf0MCvnmy604SNLVpL6AAq3m+BprnU0UrtAO/xsiK97jmBeBueJQ
OOHLDKYlyW9YmU0LOZfzW7XBT3h3qeuTU4/6rRvVGfhWcD9xWwZsK8OxocI8PycO
cpmKjxTfI6dttwr4so3FQHI09ghnFlWPUmq6eiPxRWypDbCDFFfFA72ny2C8mOUK
kiDzxZ7UZaZTP9ZMsFnieoirtyB83KIyM5w544pHW55LJSquv1n1V1fzKuAfzvcR
mQ1NFKEYMmZHUPJvJSMmTgfHqFbBEcKtpnhcmjb4bHrQAO4l8heGreBGociwjnnR
b/7JHOFcLWMziaoY0kEtAIRyyS0Do/8jbNfDgJceNC9teTAWO7/Py3AlSQkzjAqj
wLooWLYOOtHktPeLCcGYwS3aTCssg12LN9LUf3hl7vPdeTbWrpZE0P0PAAvNpMT8
+RqZo/0FBy/rZ6Iyp1HapscZT/t4Ou/lwqPX0ZEu584m5zSurT8fmbArL6xvj/Ag
L2gsfYkFWkM9hmIQOSQo2rqrRKSYR/v3mO6doxwOHcbjG66U5PBva0F48VgPp9M9
AJHmnXNoufXCmD3vX/vlWrO/qdmuJcoFnT6y2U0ILltUUz14LfUNlMtt6SYgpZsf
3ml6iHprSehW6hzjQPAv7h1uRbqQdXozgXy3V1pV7RDyQxCxYKVKwVEJnPQQHbnf
siRWwI6wL0R79MPAqZfvRTVEsAN/TUF2GD0PJ053PyUwchJun9C8fktV6GSykG3F
uvHak3wuLd8QVWoOIRxZ6lSdID0gwVAUHziKoq767vt8IWTu8YjK34MArhsnWWiE
5aymiPQzOizeHhQwIJDzowS6XqpkLdRWPdm7bkpCSZYOW0D2P68paqL2vxLevoUf
T0nMAXbw3n1QS1Qa+JaSNK05qS4Hf7peh9nFE5XHCFnptcTJuH9259HU+HEJVhL4
uLsesMOBza2Xt7sKqeXqGK1oHBB8JHMMLY0j+MMZOvl6ww3B/Vn5YhVewK60ErBC
opGqiNyR7hXfBlt6Glx8bqhbv0n609Ed52o8n0uZ9NAs24pu5fxhb+es/Xg8nQ81
TqwTuNwQm+K4Z5Ei73V0FhiXUnAzOO2BGIFWf0cjWMHidgz0DtmBYsLZ62K6CouD
9xKAEyrvtX9Wnl5v6FwnzEKppSHbJOnQJYgO1WEPhq4AQDKFAhwYGMUHSOSqwSK9
DiXG3pUHdSUyJPuGexGaUAOBModOkDRqbZ7asCC+GXUph3QeoeIAYaO0XUksQd79
P7CS2CyZfrYO1Pr77NKrfMMVKEbDCXeaJ9Br34kK8GsmpgQ0rwJlgxPgZLxkdFn5
6WQEwrd/eoipofPjZQBNBTOm1mUrqUVogWm82lT3MkW08L9hOu6d0fFZN1N+FNfp
/Dhs7W/w9hEaBWbKoruWAFVX16JIoS1ocOMEoqkrtmJWTaIopjx452z42bNuUNFm
47dK5wGMlNTOZUn/rjiQLhziY2/1HzZ6y3WfrXNWUYtK0wxhUgzzSRDfw0894ejy
fVB0Y4G5y2JBgYzjjnVzI64CYhdGLQLqo+be8ecO6FlQyZZNmgPzQWfxKeqWliQt
0FJ9Trn8nXG9AJWWHm1PcEoS+pagh8+ifpeOeHA50rLZZmdp9ciGcsGFg6dwg10T
aqsKfdvJaPy7dJhZJg8/3NKjhVyZ1XOkHEh/SOXvHTAigU50/LhdNFgq484l04gD
HNxOjcDqUlycNksfGHspEK+I+D0R893NQLE0INnPGUPL5/huv+HtobIqWlDvTz30
CeOJLz+rFHB8602D07hamEPgdHPasM1tTg+mj5MHm2CMFWhOdSZYPj9LH/Ydybjj
9aor3sfFUegRn8hTLluOoAcFs9g43HVlwX8Mq6l0K1NiWThn4ZcO9BQATwAp4amU
Fb2PZXU65NnHjikAGl4+x7/PNl3tpuxNdJEuzQJhuKDPCkWGbLZKtkKbBWyufu3P
H3TUAk81fWvp1YivY03Qkj7ZEE2Xas92F49+JqbUIJyTWFgqh3oO/BfJlGukturR
9u9Tp0pxf1C8OJFGxGjzy+j4dltNzmI7pVM2f2v15cBTLv4J3FaeG4TlZHEasxuT
/nPMxmo3Jti0luoUVxK/9B16CwmI8ml6JlavqNYTmwREFJUaZ8SV/HtwTrPXbDwk
FqPdLSUIz1fTF7xHg4hN/kOMSq3PCJzIwl1T9rum0osmtdahT7vX5pmgbrp5CJDW
bq5Gt4+lQAY44uiPBKJDJ+5IHAOgD4bFE5N2gG5lW6FMcbGalBIY4pcsBX3kDsTA
0+Do1Zs+hDXadxy3A3wSxpVIj/lJVudxI2jo5RITwBUcJwyHe2hsZBlPOw/FB6yb
A3p7IG7JvbZEMShAyk462ouuO2UytOO5lpsW0mF92aBRdHAvDM0rWLssgTrjiTdt
GbY5nsIOCLL2dXagq9aEjjE64NtI+VGvuY7owUlYZcLtAh7lg+CJgIFHu4SNcvmc
T7bLWJFmcCRDHcLPX4AaR9t7xzSdJY3ybNpDtDflWc0rEHTFCvOdbv22ZgQpAIOq
+AycaFYYclsu8Y+eriX8Z/pB0eN3gFU3G4JNIz5A02OFh4963PDVbzj+tUJjNM4y
y3nhdAzf9hEBixOxl8hJXoODIygL2dKmjYr5jcWrEdqlp+eypjNQgt+7jK1fW1dL
jklnqyNgI6s/6go+4NHpW1dFfOxjEWUCAuNwh19OMfOpt1GT6wDncbMVa6Vt18p4
hV7auKdCHI91rrkQD8hgyfPv+X9AcSQNXeRtn+O2cVaE9pmg5nkqR7VmIM8fzot0
y6kZl1bs/al5poI/yifgAuINpQi2WmkAFjOj48IcdQNpVP1NoUgzKPBy8AahilYQ
GmJGRk9r72OOIoM/JhhJ0aHcTZeuyhdfE8PJR6gE8bRAGbduZWGTtGV7jgJaBZ1L
HLLEEnYUHGA6m2f5VApcFof6j9c1uruCVv96tRg22Fm7SIPsPLFDLN1H5V6PGjGB
VGfXtgxQjqC7rQRFaajNWBiSJP9AGUpKoUwIX3a4eDAobs8M9svepkqo0fiyR2di
Tsemfd1CRkfnpEgWqJp5wYO1gf2vlUYZuDVZuAESfLgEwzo0r03AlC9RDvaPF+OE
4j0Yv9HUpGaS0o8SQN6ezF7Jhj8yyJJXTegJcuBqXpRgg+K1Yln6dk+mrN9oGYUw
YyiIKZtV0cfKwTDxjLIvsMeGBAV89ATvHR6UBNJDcbSeAK2yaYRkVr7FIlSgxj9n
rr7iJtFyCZJWXbbJqJeOXpSfdm5WYsnNYdm6JagvhyZ6iT9rsZnXNORIZTlpMTYB
s2W1Z2tPnbZ1nbvUkgdaEL2TuFNII2ohFddv+ejDi6EfUW1DCIlT8EKpU4uR6Scu
xIWrl+5Mga+0+/gNVedKuQ79bGiWJL6bFLHvLagvA9K2nxgINhn8uJqS+vaumYmf
WpnWE/NGBhj0qVURK0fUc9zezU/eKGT8eTXCJcUKcfGqbPC/9O+7PA+lhDwSYIKq
gxPrEe56uhXIf8FmdLaF71+9aAGCWILYv/ue4WvVT5cMf3v9VxSfTOHDng+yqc37
iUr2Eh+paV8WTBiqcNFj0f3vos07UmdaX47k2e0ywgmjxOcJxdvadppS7C479YUj
WIjjZJIqVUOo+KbFHfm8LqjAA3qqQbHIocOPp8j5MnGSlPXlT0TBxbtCz4imegCK
2iZXE+Ij48WUktDzqPMJumeaH0kbntz0eTSsO1e+mOyS9y3NjI3sYx5il25TIlQA
yPa4t6IOYca8RhJxYWevXV5mdvvJ9nbNDHs2qWVdcjclZXYXotKam0tK3Ph1D91m
Jrm0GbjvhFT9tk9ckANikRVsxkA/X0YuXtYAa65Kwr7S9rfQlSfcEaqamFNhJK5q
Ni1SIAtUpS+//U7HkBlXdCVcaO7m42iaJ7HktWcQtdjONdoI3UqGZNNrVv44chNA
FANhILT1gLyZ1zQYtMADfgGvOVZRE3I/snA+1c3/B72cBUeMaokKodtAVqTP8Ci7
aGvkGU16/Ykr6pTPIiZc4LF9VXzk/wvdKmqo40KSKN6GVjSpNlLCmOGQ9iFlevO7
CbZqMuY671juKWyyHGE43sLEh7R2Q7kpewO1wCOd91FobSr7hiMlZ9C9Q5/LPBV6
YGwylKWKMUEP5xk06JW+ZDzK6wlDiSeMXfA9lk0AZX1hR15+Ym15OtZs5t9/JV66
Z/u6qu8ajCf48bU1e1YGuHxtFabNxvql9AjYICx2wBl55EcMcLhfg/lzDTiQy6XT
0UHGfDBDsYb3KYs5oUVAYkQYryBAzQVtySx+X9ZkZivTHaA5LmPCILLMuralpuQ8
Di8GLToTduJvLuGj9xQVSTCsR/krHnZhgXJsQv3Adtkl5Gc8jcznXQ7UYP17TsRY
wnG1irgdA9q9Fyd4DeV3UgiYh0oBblbYR+3EqIJmYKHHTxFOt5BDdQBhykYL3ioS
3P83UkCpZrqC6h7+rdT80+R8gpWSr8ir7ASoxILg6EjkUtGim0uoD/TakXajNOnp
VikIFaEwM0keQyEcjnPr3rWN5dYFLjkxPu6HejAppo1dgawQ5iosJimhbPRkNB2g
DDP6KlZhZC7pwgsFvOpTry6FngsKA/VvhQRWT/tgAFgrBHm98Rtu/UnJotU1qaEW
SnejYSyCFk09GluVZs1/E1AvpckyR1vct5jNnkuO2i63ixU64ULaYotOPIFCuSPg
JNs/4XY8A+QSbX/VgVYHAHiDJuS3vLnftcnrYO6goJ5tjNU0BkD18JU1H9MR5r6V
DHPahxNhcooWcd2uCnJTDez2JxBxU3fKs1BYf1dYyTygPDKgeiPpT9jHw1I5rOcB
Bs8zOHFYdpyBRQQTbcET+BxvNzmKJqDdggd7KS1hL2TEIxfjmKgubgNkTu7IVcP8
On4f8ousk/J48xaWM6jpCFXQNdq3JkCfB3ej5TDcIjRTNJgNhmopmAB2hFsJ11Zt
HLj1LSLNJBbqdojYMjwAFcoc/fubzWaz86PU4lbgImzN/wI8yZ3LQbb1d82QJuyM
RD5EXqyhRMQhlIjIiuhBvyQ/Bs9Xr7U/tpgCmhTQaKc2QpKbev2q+IO4RUrwFHws
k0kiaiHSRDdCYyikBgMgaMa5jQtf3XJ78nyRYpe1aphjcmqFEo9nTpzoxuJfEKxN
JrgWpAc0jSrTDRzJLH+vD4ggS5NmztACBKtT+CZAlOljUpLIiao6qZ1IL0g8RAjt
qn+i7nUJ52J7cqFSVV6RylDfcR2b/6AGjrdX1taLWSG0BM6iDENFms6A5WbMnyb1
j13quEOSR3wQAwStU0Lmz0QS1EC8tE0WotEZT1Oo+LhQTK/9b9DK+AmEPVxDfax9
CRWrGvO9FLrl1/dNAyDSJkjPhyHOFzMh7JuOr5zpPpO54VXIJawGjuN81sqDMOtr
jX04CYk47MXCIeBw4eMBxKiiAHXuIuCZ2x0oRAQOmE7sTZJFyHsP/oQL8ftYADbd
8A5B/y0WHZDs7+6vr2lYROWBqGaO3JfjQiT6KKeixIaqhVjaTtrZ5CHjwWbajm7u
dgnbwpiD8CBnEQSuX2XHVZhUE6sSmzWyg2R0lbRWlCGTFlU6XZmf5VLnfbgUp5oB
a4Nb1+3V+xE3HRzEkAN90bMvkUqsNfbNoofC0JjGr6tI3hbWiVYR0Uu2FxVS0SSg
dYHu8qDnnpchLKxMuKIW0zs1D4ku/TsmsA67q4XXzUXfYen2mM0iAO5bwyaCqC9E
OiXrQc/GQoaMgur6gsmygj0nhI8jXjzOUo/R80PBwkn5sANkWKhOs6206rDhodOU
e84IPSfw8WK5WZSMcXSU9VgJHkddqvLyONmW8DKPYr8zJ4pKiPP4Aqhf9kmCMoVK
O+tdK3HILufRIT1fy2Pix+3Owxrpq2jOmdx4BbcgfRQI6gmAiC6L2tJJQ3d/uW++
Od0U6XRmRJx3jvKB9b2U5rvQASyIN/AYTNohpUVyH+pPpoizYW2b4H1uE0JrENS0
iqMfXsN1JhrWZqNc96WcwoxYY3u596D5DdDTv7ekayGaDtmDwCO2AUWoRuO2l5MU
b66ZB+5w6ZinV20Plju+/snkdL754QPsmYXQKhVQmjvAecnu3lgzdhTnYCIlw0HV
+UM5rgB3iwBpnBoX5ZzQwPh8XO7iOajmojXD8WqP1CZJ3GXuMKEQkrmoAf9ri9rW
KOwd/dL6BtQ2S+OceVrlP1e4R+44BieL4Ggnb1rYIfwFtsGo9lIrLZL3MioXeI2n
FrfKn+5v4QvEvEjEXYx089JuZEE29skKQBjKOxg7fodm4mpFIHWJ8Hj4eU5nb5rv
V6jVDld6dusDUOk5yUekyH1xbU7iphEplHwmi2lUCCQhn9lnYWUAaEug/Fdk9IEQ
LDU1J0L0RjtbMljsu5YQgOpxxb5vOQd/vK7bf5HbDN08CXfEZMoHysU+m0RPcGpH
TGmP8ATf9UGu2btGfpwQk1YqCGhLcR4qX4JXedoemEFvyVF9oG6IwwM/Zpp15S3e
ySFemMvvw+Jv5yU9H4haBEu17V+rZMhA+I2b7qEFYJAZ99BQEPCUKghpQ3YU4r+G
hg49OUp/BAKaELV/mvawgRD94fHGxkza/9cUNbVUSh0jQsQ/ffHeE3pk6T1tTsMK
6ReFNRd3KuCq7vwmqofO435D+3y7YQp3yOvtwdjLFuEx2GeLSH9sCyIhthZdgVSZ
BZaq5d8+b6321q2L9AgCMvosjfR5AuQXkzRE7PGllLcISGsTrdv2f/ouzW3rgs/z
C+XEv0NIzXQ5DaMvqMdskcZl8+uKXlW3sRBvQS2pyyu/K0/OuiYtSdcHMQ9Sj+yF
qRkBAESUXAIGtmB05/eYuQ9kwgiM/xA2ZHLTwy/QrXLxY28P+OgY3A0+RnRtwTRJ
NT6uM2QywiZbhBWFSm5hcQNiOVhIBmt/WMG9+1Psc3KRhHacON7sSmMvTPb7Cy0Q
EQxW1/fDoQL2gXEuYvUn8NBfw5XAjLreFUr+gz+3OWTDAxhVXkS3EfjX5q4A/bwe
MWYIpVN+j1Feh9O9CAToDbuzWyg0/BTUjTNrmMqV3oOyZCN16oipMm8HC7717HCA
JpxJiOk/hzu2nKtANCTgTmLuIobh382LDFKwOQaYuIarXPr3ylstbATYG1fIB9TZ
2Kan8zWWgWuDgSMmXPE6gJvmcFnaEDa76XsCehJuX1zieXmmjKXYVWXnMZj0df8q
ngeopvSpiqwQ0WqHTBL15Ly3CxqsWPBTyOpaMO2S1EhkqL5xZW82kuTvyMUoriew
FNxQJVXH1Ea5rtb/EnAM+Ulbk9vSTt79ACvG7h+dv891fQIFgLq5hGSAJj0fNwGK
Bygi+DEKfVewwJYQ2OzMpi//wJEITiNKtwQdavu59UVaHiERtG0ncoeRtF20ty+i
Q7rfHqQ+F033MMwrI7AZ882m3+3eb15qaIf9H2UjxUpSUdlwImgleuDJHnl4rHeG
O438QFDDgcbVLCfD7YQhjjDQqh8faa58iwKfbCTYodVSxM/JGHcJOw3kWiZQYJ2b
K8FPcF3FOYXKoZ4UYV/kjdJOaOVi05nsCtTrGG6WPtcPLmmABdmdlhHhz4oPXSqU
goc22fF7Mew06U5gdFytdCw5Hlxcl7APqiJlcZjmlpN506rdzU+pzKJG7xF7kX9q
hhx5uJ+IFNTajk3KZ++rMOs6pj3YAFqGqnmIvc7p9iZFocb5zmxETpvSwBuniNBd
MAjC6gyojUfQreuOdAvwxBd9EeLfFBNIaOWBmuOEUfocIzIpAlghX5aGo/kzy1db
XucHdLX3BIuqyCu4YoSUrOZbVrjscJCApUbru05vdmQ2WFh/frljud1bM60EJyD6
eEk4jXukPQ33y6YYHcI20j9oljDmsk8uFWAXgM//AigIUBKWBlIZ6t1FwUAkpLWd
4yNBg/IL0dAthyjalN6vapqSXkRyzlQHRG44E/UdOJcdX7e/iO5kJHqqB96X7eFl
3vEjVou7ebSJBZ4L/Ra3WJA0pz/HREwkhQoJVYCK9jjTma6iiDroiAET3hitjlEP
+fc5bO71yyhdouN8rDK6lJLhgekztLkruL3Cy29jPuA2KvqLBZyKttV+2hllkKsV
41xZFqurPlrbm6BnaQowfLAIhwUD0x6mnPJYJl6mMkJ7EMm63BpKvoQjf2Ylf3sG
+z4mbPtxqQl7T80gnUW6z1iEPRTr1ACtCNahgm5vMGvD+Yrg4AogPvLoTbdgb7y0
7RcT94vZU4FbsSbTPCLQ9YlW7NMIqsMgdvxkoQdXF78wlwRH0eNyWN2nSOyghUBt
rUs3MFa6M4NM8Jins+w9/hP1Qm4a3QzpkvcPLZ/PD0wFYpEbbEOM8JWwFbQrN0a+
LPjTveVwzNwpliuRHpE11iDqEFcsZc++Y5Zi71SSAogqA4mMMDvPAQ8pzDvKlDE3
Iy+UUTs7V5T09cgx3+eB6+tMKPzcsi88Bsj8oGr1RTUgvUypxkr9neHtJ0xjTFvV
1AkewSP/ZBvA9AwKuCLsAIf4gpwYp7RiaiXd1JxaGh2NnVzul3aLxLhIf9u1mxd0
vWIKs/Ai7wZ10VAnz2OqG7mhG5rh5jypf/ITnelmy8U7seZW7Rp2MwxYvKKA8O6Y
ZMWorkIuJT4wj9aeIofL1DG8+jWYqcVcWqzBpiRTD5jw1Pu30fzgf2PXpwZz3+fO
lmIgw19kuFj7tEfvYB8qgBXIhbAPkj2Kdh2U9muFFiog6Lzo5z9HgiD8r2gNgnMh
u0w5+Nrg2Lw/8jOx40K2yHTFcf+m9iCgqC1SnhPSbUhiEzLhnnJ9r9S7y7c4xfqk
eumNNABROBi4NGQyctL5rsm1cA8REsZuFIoM1APYU5F6q2V7gl6PNV9vw7mvMaDp
F6t6g+RIFr5h5IaZeJhlpHMHbvwLmF+3nm1XjGPf8/dqidVdTGgRZgJhnZvDS+rV
3Fq2LRmWxfUpFJHDxFm7S3PmsWqNk4ELnz9O+mADwZ5RFfYsv64eP+jBUbwXaYEp
6X7Bqz7nU9oJeoEwOyGgi4yCncI33HEc1Wi/4bfZJLP5jXn5NNuE2eunaqDgufFw
aq4uBhrGyIHXP1aC31BcHJNTz+AvidgSRmGxpmqHdqrB+KJ2suS5/1Zrmn8hQl+P
TOsI1NvSENtJjs6b5ZX3sHV0FzKNc+yGagJc8V9V4Mhy5y3Qa3GjlekGNKKagbKK
iBUyT+W8E/gF0b6aOY5HDbii8N1htDZdJvGxXffu+4UC5ppU9GvwhqSaDYGc6Jq2
3YUcADXMVqXa2605fu2juJOxyWnc07f5V3NA4ldHboFqcYwEWHwI8NWCoQutgn/j
L4AQQ/8DetBNVYizFTZVFpkCReFfFxNPwA8YJzJslevGh7k9NKBHXTR7bL8aWCCq
74/VzqzZTqx2Sh7a1b8ohKfvdBXG4oOvm5HvGuZFJbCkz5Mkf+241pDwfuSJjaNa
LMz4pY/SW4muizyIO51nb6EOMqP6YTq+vqUeUcFz+IwCQXx5uEWPd4cdgTixr9iI
ie+Z5h8C2/6O2vCnorrtjwtCbN3VyTK6cc5H6yfQO7fUKTWsAMuJ4t8zYgjFVI+I
8KUFVnYcFsOTb1wxu4UNYBunVtj0VVrpL4BA1HDjcTpoA6VXczNoobLfwzX0kv+r
Cf4oXgXlIHMQacYzjy7kAP4M7Sri8Xd3Gd4W3F3qgYhlCDs8clo1OiAnlJXT5v+c
VHmJZWSPyMVFchdBem6rTeTbqrZuTYPyQzV99eSaRi5Plv7iJsSeiKDokdKVO6MT
w580Pfr4lEp1f5yfy6T7IIgauL2iQMZDYg956Kt5oQL3li4q2ELW0i4UMXw/oaQ7
1Rr4T1Kfgiy7mooH/6EvQw+Imr3qNKyuy33QKAoGtWSkSfdeqO96RfujAOAfxpvA
5Zluy3JSn5m3XYl3R8Zx8oqjv7D3S3j74TXUjGPgxfbZkQ0E9DJf9876ovHGRknx
Hb8TD21Af+gLtf3Q85EInv0/HfbjnZsFc5535Lkg0XNQHqWuvdPDKbfd4zeAonAl
yMdVHkVdvDbaxuxDtk898WnKduoMJyRO1P62zvAhymgy/r6bnld5rRB70QZ+FFYi
zc3R2iGgOCu4vcPcCnD76M/3+X57VfZdMHCFju6PYfpL8f+AWXqB1MS/ufxOgw+P
QO81ZHCmSOpqiH8ZrfkpbW8KVU43e/IbSDmKltLApfugm1aeRh+TFt85sNVNLMI9
vGl4VXC9x9o7Yv26q8QoSxmvdH+C7n0GkD+n3bbHUfFeu43oTlv292X1C+VX5ohh
3rPEE3SQwKCM9GtPmmFZRO4gDko8ehin3sk5U3WdZ2Kux7YZ22iTY2pkmYWi9ifm
fBSCUGQbiBWPVfVrZRMPx4M5IwWCULzqHlJG+m2QvFMColx0mg6m0lbp5e5YzigY
7O9CF06VlDIBkr1P6rOmCZTVfO0Q7UfEZ8u4p0fuwYIS+4Nxd39Us7D3WbxRAq0f
XdysP92E5ro9BeCghIAPvsyZp6QYONvsUWsY1JG75aRy1UYbNj53cLeSacbq2IPu
4OcQEetj0fZ5D1Ex+eJH87R1QUAORYsUvf/oTCpAstdLN46UO1T5AQ1GELzjPdj4
/EuOcY0rmql2wKKCvo7qttv2fHSCGql4NusB6FesZWhmogP4MeETCKPVzI7Ffwl0
4pwZIy671cIPLWoLg0Y9lzQIGt3gIXcD2XO7GWgGp9u+Zt38tzmx5MQNAvE+RqyN
eQ4Sl9q/u2b9SR4JibujJ+lrVVraeMDjkhejn4XYnw6XNInfi1JLfl4B4AoMA5Df
yW2cyOUTEVcAa6ATaqvYjnsKVaejG1Eu8gHUDLTGbeO/ghqQWrTXtok47bA+WRt1
u2GJ/2rF2tJxwqvYK7ywbtshu8APOExM6xgOKuRHgUQtRXwQR/czi1/A/n/W2crz
l4+kQvgpL56Wp4BUqU1xTzABp+olyOPpQbNaSHwxTFgFe7JtegXxOrnQ9nVNLNCL
xtmMdMp99bQRKyqfz+K0sNV0RVA0lNL1WNg78NiEj5gOXGo0a4J/Zcxulw2SYfHT
kCiFqmPIHPWuKbeNAAjmnkkk+7eSPiIDm08BwsLiChSEw3n1MC4L8SdUx09rL0y/
2oroMQH2X3LTG7zkViXdL9AHQhFJvvaTvRfmWhGWgEWZGSHFzDUFaga3yfQL52sM
WojqfbGsobEuCJwKSJIWJHxpXCIK1N/LmWvSk9N08YZhM5Xx2K5kBo5MONw1X9ks
HFjTaknbhJystJttBy0wgSfmLZBlpGRM+FT9m/CQbKlIW7cPcSWmtjE1KHhJNfc1
POCyNL58eRAGQ7K0NFS8ovAKh8EAdn/aQCT1O/KPETXSuG5mX2u6N9WA6uxzU1DY
goLr0JCH4h/8+uCZHZrd7ko/FSWw6XTUrM5+NOM4fU5ZDGeTFt1ZW0jt8jzfi+EU
4NsmwzR9EDTpmsyVCkczQ1RNC8NapO4WGdslVqtNosLhOpDyCJ7xj1wwTWYbIPUP
uTJ2CYnXKBKEEU+FawmGO8Isr+ZjTb4qAS41zqhyj3hOe6D//hryhOSeqC/WKd6s
/sT0SmraaMBbpyxhjOoyjtq782ekZVAYuUYkhNmNTI58TSm0Ree2SZGnWGJirSFM
CySDov4uBmEKtp0om/Zt5lafTIUCe5QhjDUTTHQGFLWUx2XtWrBVeH6yuBzalCiN
tTizTAqyhmHFcJexWoimKzodlXNBeljxpSp23i1VHm+oGL9xj9y/THj/P4cpbmOL
nTgxyaioFDIQ7RdWsGCpDRyddeaivEvLBSJOg4Yq2ln2pcOcQ5de28rdExvzg1nJ
RZWhm2uhr3Yg1pDbZ1phMX7Qmwclf7R9LSSG9voi79wHAaFoB3KQgQAGhcqc4Q0q
PAEMSctrkADNRVrAQLDGMbWL8zKsjbsshbE/fn895kR6Ier0f1OU44H3Kt9y6UsG
UcxkUJC9tcTppn5qNw8uP7Bl3Jy3dKCMgDQ45BIzsJJdUV8M08GrINNX5Fpr/YWy
mU9/76ABlEDBNHbZBJT130CnHirQN2aXEL4OefBShs+qGDJzRaUvvSRvAbNagOQJ
X0RPBwT/gBfa6IjuvoI+T+p2BG64TBctTmiO6sjCNoThcMN+Kq9ZYLUyHGsHkK+/
qdsTi9r1wPt8rnV/NqgWvKlldvu9ryBbfIMP05TiLKebEQ8jBThBkRyqu1XS/OWn
53M9o5y/ShSRACGAc3DTGhhkx7ahk7fcTngAJhX5RlAW/3CR2R2ZxGFqMD6739QO
Kf3o5cH9pJYX5RQxRzb80KZ9JJ8ulBr/M4jeZSdkCn4gLnkGgn9pxdCCUCQzWQLZ
TK+IxlIGRfdQY2ZxhuWPUT8zkOB3j4qclkKPa3lGkDQe/5GPqvU74F+IH6Cb/oh3
Y+ftlJjHuYP/Qn78dbWWzgPIgfBZLXZjZAp08Yek07kuDVIqhktdJBqHgIxXMW9A
yfas5+FWZqQLhFutfW//jaNCNvf5b+vto6AZNZJStkaMwm1RhTBxQijlA+DxXr7W
VT/QleL8XquEEjZZZ3kqyKBJx0X6RM4S+EndDNv0OEndQu/FPP2qhp6Aqu1tKnTc
K9Gny2trmMGbivcGr8X5VRNXlMekS5r3ezF5nLvJm41P2z7mFx8eEpYiN4PqhcrI
ObGZEMhgTzicZR4vW/Cr1J8PeyR8h4DliVQe/i3j9yPKEJGC5n9YVEUjk+dOWg7V
m7sSAcfN3zuxkqZkaIxIqmkFFlaaQGiPuhf9QPnPVp+j80byZuOgvne/yuO9+lGD
+hcGGj6rbTHpXpB3UaFpG7/KZYSdtGLz0V+u0m/0r26EsrsL/zRgL2/WQBOy4HUM
5tx22/uCyl5a8gKi4UbuSRMMmhPgK3Bn+ArXrMjlcApH69IoWDM+mRvJpBg0dWCD
uWgBUipiIIzwJDCzGIx+NnmLHr1sSA30DKfzqO4aARRD/BA+fAHItbAZGhYHjGaQ
LpW7njuKRzYUmyEmlo0xwAVHCKnda02gn8JXiVhDu+dGBl1Qal2onBshruSgObIZ
QK0IW+IijzZ+/+KJNjNHXsRmrGQztZLovH3o9FqIVSBgU9dnUSTH5qovNNq2jGiM
0KC7gzhhgAXvwmHhQl137G+PBAf7+wEmhp/bkN+jtWhIGnxM5F9Ukzg15RwoNkEH
GDl9Del8BbJVjPsE86xZj3D5npO15ZzRFksH/NSyNPJ2f1xdgBd9lfuTFUTxwHgu
6qsaDGgLPrkAMYjgRHLObmnxAfdGxe028mWL7jOZYHeKrJJ2lQTONWcS/plOGaJW
lPRHb+WPMK2LinIKmmJ6jtjP8K8m0UOBqPlO3o0bAJheIvXhq1HaOY+wdMwSXC7L
4oX3g0GtLDmDZ+gPN8TbGz6ZpvpNUjYxjezPsku34zOrVvrvst2mjRDfxDUqM0dP
fRQi5OhbXqlRj6UTcC5+JXpNoG53FU/ZWkbzS9sBThfZJFkggdrcCqFxG/Gw0pS9
zzqW6Un3oeqOaXaKHmLMThqVYLmc6aGrrtfs8mswWCfKIYTC6a3xxaQpBhjgsZEe
5/kDsOyzidd23VovGu0O/mRRScgSlIJAFK2B3OGvWjI/7Bw+68sZAE2GyKen3cm+
dNfrXx2ZLSjebIhBrRGNz8iadLK4L06FtOr3vb8wURzDRp/JTCmft1pQ37l2eExF
GTbEsEz/xYIcYooeFGlvwWVVucaGWLVrihqLAcH9ca4rMOMsJZKfyG7ZH/QsJlEv
cq7Bd6LsQnEzJ4GXm61cLkaHgYYAZL+I84ozE8aTZ07Rg7JzRpFxZhHNLp1vTy4R
HioLujrQDEtZGEw+oPX8tGK4JSZO+EL7wMRlYIm8C4eF5tieF8W+QZb5j7IXUHsJ
c7P2dLFou6+Idj6l6FQ1lQURfxA77OanWGeX1bBPhc4qhljnVMtKbrL3cR2UY4Fa
zk3qcYfPAhpZVjpbRCYusUqgqyYovC/BijXANBtyIHMRop5OuhnKjSjrKeQTUZLJ
m7Fic1ehmu59uyVOEHumqpLhgPoDxk2bIKDPr/UImxaIh7lwhD6e294IlOH4lQKn
tBsOCwe0EFX4JBYu5e/3cX84h16EQOCvAjGE/VrVErIV5SR4/8WsyMWbyv//+Oem
qnwmnX+DHPx9voX6ZosFnmL66378MeijGTYYl/+IiNOmFIz7ndcQgUnSKM1zCjQO
YkSTIg7KP+vmHH5cejhmKwTjkgu04c/O2i3W2bDzEc+CdsHAsnZGskl64BmZXMSj
Xn0S5WTkZcgCkHwULVPhIEmse1LFaiVBA2PNRmalOSmC+lCHbWXQ2bUa5ABbqqle
lVP+DUYZlobUjX0Aghu6Ed6fVFGSyHxXQPxThegt9ODm20+GcNg3QIW0CzqvHmx6
o1ek1qO3CtGxv+pL/bwoId5pX1eAcoolYulN1Co5mPu7TuS8V8cWHRaobGkwQShw
v2orEIx1LPE+i10gx4PW5XgYiM8PjOe+BMjwzMgLQhT4E1x8tFK7cg6RTrcg4VhW
TuyvLaLoOCqKh+nfzBVAAxTkzjMGlandzTCPKuIC7Egwkz1prYK3MGRsv21r5qBM
DSs/wEXuBOZEcYIaulvoAvToIUC6EqfvHlyQib3N/lmPFfaIkK1dPTdUU8KY4p4v
A7OPwN07sp41TmFlcLvBcCATd911j5BSbIFIXaxoOY2nnsmOyDWDjWnD/x7qSMgS
sQwlVJ2xdOeSSnieblyBICZzblDgCcE1DjNBw2Bgyn2f90T7NYUvc4MAqySaVyDj
9bzroP4ORq+RDARkK/HABiH7L+j0pUIRIMEiq6sS8vgx8+I+23V3f7vWuyN3ao0L
unxYniKFyMsIUE/4vIlTBmNS7AhcTEObmlmBLQJ0T58Gyyb+k0R4TMhnd4ynvOx/
tbIW68li9Dcqp2LAklk30UzRHMX6vhYNqkGQX/6ZuajUswpZ40BDuJk4ZvqokTSL
YaCsXGPNUtPCsujvNuL35L/X45xgJd34IVREWNSRieqiMRu1jjvTBF/zlEJMWOeg
HKNpuohr2Rxa7zanVsBd0ILm/A4DBfFIzRPelJI+MS+e4oNN0xGytTt5BCi50hia
ncF0pPZqx2Q0huxgrRYUsU+lm2xK3rDvbCc2WUpKRkR4J+AdhZRKzFb4pLS3mvmX
KeuNoZHQsZ+7H+xm46aTbPjDE2Y4+qCN81OxYaaw5cQT01zKUgjsz6bzSXTZ4fnt
zOhfJCu9T/4Vz5KQ/dIkY5q0pP3k07phouQAIhgefE+3ViI4U6lmG+dPh/+Wtpj0
IcJQVCXANy8q3XiLViD8ASfBjvYAzUqLpJ/YeBnXI6MtfZtkrwRXSCz+qAzZTaAw
y0tS6/LuqCDS1AJF88AvK/C0zSbbg7GIpOiXLIhodqJILU1FkNrbRVkCCYYEMalR
DOsfAIKJ4iySXwzLNyMeXw+0m0guPRzAjjS8LoK23OiTD/RMuoK4WnQmaAdqpx+K
UKxlXKOj31AJhFKPMdJnmcEO+Cex82gS5QQLGcvtyC0HqvauX1hSlpKtoKWmgRvr
H4aUKv2u7B0/6DLqIpQ+RAF1qz/MjDoRiEbOR0t6u8f1TKnr7PRezoaOE7ecT0hv
Qz8vtp/V1l4XTaEHW0cYoFZznMo/Olu7aZAB/1+NU5OGHPrmHsVsU5C35lYIDGpO
ufWIlfsZ8JYphWOGcrsS/98BVnIf1ViXHUUXxmGshSgvn4woRoyuq/k2upCiA9eh
plGrftXOyo65I6gGxCu3KCcSwKe+5kR0onZ6p4EiWqd9vET+5J7n6VOZylF57D5F
P/acEDg+k711VPlBs7hTeT0yzBgxG9sNZ+mYxX3t7y0VemGvkeD8mosZeG8z4RWi
i5KXiaT9lyiEg8TW3enNFvCwqbUUzsWr8i73dhs6OC/ba2RZnfROWDoaj0Wvekjy
T79UTo+tMa1623Flje0jfEIbgH3ZQRdRQASIJxH8LXNZMWteUds5odQZZXGJTpGY
iV+jdl5hZmhdc4FnKs7li7rBbvQu/dY79IY5O6ZP01+qmyDE/qArEPQPX8XyJSus
pU/lCUXKo1xgUw4ANK0XN50OAWdFUthnaaYvEeELRxcsQO8jCv1/ieKslTsSBmMH
KwvFmCG4r7L5JjLZN6Kptdio9dUtXfObwwguiC4khAL/p1EUWlC+tkBedD0C0RSV
ZZ9srUDfL0EpYHuO/UEdBy+LqAg7V96U7Dw5JYF06bjpNSxLz2+OIT+6GHFyiWQW
YGEWz3UKi6fx+2dLlKYjoW5ODqkS5Ow/gdP9lYxXPPhcGwU9XVdoNVbZgFKeh8rm
ScOuT9O91HAnPLHeXspLU1uYg6TIkfTwjcUG7oe6sbw7Q8lT8Zs/mBL+xxDP3Lr1
0RFg5ii7S4d9kti/2oFp0hV/m7ErLuwSaZzFAgvMSE8bzT+/cIEDs9fizrkcLFQR
Dr/kFr2qEQpaNXIEabzrEtzJmlc/myuPK4xvjos9x6hLUqEF6fuBKbDht2kDHed0
dXbOzbj4/C5IbJOJISQbpNzAoT6UMdB2AcRYA209gvDSd3xEFkqKzyPpt0TmTBkS
GoQVxuUvPCrifykWFuR8/aBSVKFmLT1zdPbz0e/V4rNNM3xFZ2pScu0O+h58GSL0
uGOxaHpxGktuwZsK7hx6GgwbXgaRBk58ExXZP2kvjaNEe3lsPnQLa0vHuXsrF7vE
rgN81WRJ1B1nAs1bIL9ndy+GnpGV5xpRi0cXPbpVrWIbWUlnNQ5QsAofEBPabGb9
dTrjEW3anumCoDPoI4bRRYYzgWlgGno7prbwjlfjPTvtn2UYeW4mpqbzyPSxvERk
l4WnUGQkBLN6CmCIhlrZCFp7aQUahGZQY+DXjMyjHeUGNj9ZcCnngtRnd35vrpMX
ozxa2MQAD7pdk6FyFY4nL22UgplwEm2rV+LHnQMBEol4O8UbXR6BKccQFj1N6Pqh
tBSFNvO9XiW/qBZ2KDQxwadDLE/YTAxwb81CIrQbRx27gMb/8yRPcFQnGqX2Co0m
Q1pJFl+IKmdTRVKHmx9IAvh6PSusxe8oCxsl3y+bBOLcWwlVyeyyG4NYOQv9OhIF
Cb6CvafOrTdzEHxcEaXQ5vxlAiKlTa0nzCzg1FMybJMGfY0yx6FZ9/JrHhN1IclS
Kpo/8zhErIxrpfGDCeXHbeAqgHGA9GjEMNiKPNGqfwBRvHOXA4RE8OMGeCGGNcQD
uc/q/LitNq3HdFWA7PIauO8QWtdnozfeSYf3jUl2OJDEnFLqEFKBiUgIPh2v+42Z
z+ckpkH6vzLIFutCQECgUrCBlfNhpqtpobLKoCujhAutjU0iIqJPcMGO+Nis+g6n
01eaCtLsGvc+Qp1kVbY/Ee2Dguf2XRB8yzChIQB0FK6gHdghhJWcRsN8vw3vXgUo
/Nk+L8cfpjIaM7KDkJ4bqqvJ6HwXnpsi1yvAtQ8SqAIvG1XvYMy7/+kVxBj0yBxN
3iVw2lWF+3vj9DYn+670T34b8wcySFz4PuuoNt7nfHQWhULP7cj733MlgIO6IwEH
0bmZFJdP43JMBO4SvYHQqPqGpRv8hoQnKAyZ81S78XDAouuyuSlBV07dMbYwFY1m
14dG6SP8tyzFc2v42IhOhlK+bVlILnEW7ehgrNPtyVcMraGWdlFPkHSTTSfcQK/6
ztMkmV3rotsg7ZiBmcOxAeHRrhlsSHvR+SFz072BwkpRvwE1L+UV7prDuc4CvBTt
9MjVO8eP1V8Hka1WnHQwSAT/1gliB1jazXbUb6ksTuCbBL34pM4y+vmqn0beMGR3
OhkQPUo+GrA6N3gu/pd8zoXbe8Id4wMBG/Rg53Hr0aE01sPcW+L/BeeMG3OF5bk3
Q3bbV5/XUDj7D3+WhukYwn4TwPo483jfpZlfOOwJXfjntthtGCx8TQ31oBPM7RFG
JofZc7/ErS7pJFM2CG8Lz08Vcp+LpziIrwBJv0dhp8rKEnKcbRgc6v7JnuV06E33
0SRyEjJcrxNAfnWCKJeqaLpqRWWKlaFOTqO6m9FJbNlOfF9m6sSUaE8Bhh9STMyQ
Y69uiCnwgRXKvpzV87Wcjlp6ssc2U16UjRwHrueh2cnmSRGKkjDcfnGMDDuFuc0C
sbQ5wOub6ZUFPSS9qV+YQwB7KRISQ23fBtYwyI8qPvwnfONoPYAdPr9oP8q8t8Vc
K5X317SGsICn4hKGbgGtUmPD0xE7/VOwMglfzo/7/JcbkKYNnX5I3p/9XfsT9cw/
V1KffVNxeX3UKCjsd8kedg8Sw+fgUkZVbXj8Vi7BgTn80OZMxUT6M9BZNWseIjYn
G7u66P70yjBrplD7+RPnkdL17wjpZDjrlS6YLXCmbyDhGmUlE7MgSw6sNU3J+TZB
VL8aEsxlNndppGuiZsZTiKapE1YYKdFqfYc1tDCg70teHkwwvC6wB0rpGcEsdVwp
+0c+5wSr75x64NY+cE6KBIn1UfdsA+fkwLzUEJNyxrD8GFJnoUZIiJGayXCRD1Gw
ucus4bl3wj7XVVz13ENIuTamqQC9CtpfI5sayFjc2he8vOBZD/AxdxW0h6jpGQOo
HfUEy/tZYnwoM0nIJr22n4cANpgt6Uc6LZMpmS9dEC8pAnz9qzUidlXFqtS2fttU
eHVs87KFGt0tN7AoS4M8AS8qEMSpsnEvtl4T5RtOkVHrW6nhAqxpbQNVapXPT1wd
C2Nt5XdA3E5YzyhCthdQDDvssfvIL2zi7oElR2LlC1jXujyzcSbsLZWRX2y7uZgM
Ms/oFULra6RkgeOK3dn58a8UuH/I+bDn315+ebYHSASJlTG8H5lH6cyLITTs/RcN
bh+WvP6feC3Do7S96wWPwP2HZcOtDtu8l0Nfe7QCQqC6WRpdyGwyNi3QtHmgrf5e
0aTHUp1gkGR5e8gnd7Z7ou9X8IbauocMemTuH/gNMPnxnvuqmNGSpMob4hVulW/Q
RElSeg8KbhFnXggG4mflm6R8ey/TCGtlGfu6308MuC4GVTCqS/2ceo5XqsnWdLqk
kwyf+JQkKB49K/Db6eUH/zdF7paMbObDOFji+aTZ5Gr6aWEzECWtTL0qXPjpxblp
5YY+7CyAIuQNIgciRu3Ovw7Ske8oYgC30bbqF23iS2GNP/ReHzJ+dI/Ia91VSbNz
buJdtCab5MIj8l1kESYk3Z51oVG30EYPqPgGx2/ovWrQZKNr+4HgM3nlL5yjSEk1
N8jS9YDBk8ProTNWQXPN7va8+RUgOcIcoEZk4uuFNn+Kdqb1VLQgFZzJR6MIvyKA
4+NYPN11EwYaYPv3sAzNcAtXLW1miAdXkVqE2C4bUXRCaS04ALZzKewrfnKgaAvh
rqP/EyuXyQNrpNmYRuz/Xor+eRbsFTBwSUjGHBnNwxXT34AE+zXQxn0bq9AUF0Rd
M5d/4XWdT0IarKFMMOw/IlLRHG3Sb8nymoykCa7R1L8zp4494YFlhb45f4Fh3JjK
r2aWRqYo6+K1oujpkFNzGe4xbV4uUzTYt22QL6pk4Z1PdsTyHPO2cECpbjhpE5Rn
zKXPhubwbe6EZmX4kzmvA8b0kfhxLdtrJqm/roZlj+JUp3Pg5P28Y2+aA+llDiSK
w22jS4JcdDqd/UiL623olaY3OPp4L3w615zHPvCAig4jDvSgz2iOWikFEGdF/C8g
St4bFGHkIoy5qDsxKeokvPs/PQ9elTW54Kmpr63yklCfmm+vlhaZKGvLQPMhySSW
v+nBEQg1qGsHyxugPfHhuqpuuXpWoHGI7+UU/MHRnKQ0535tG5Npg5LDu1iEA6IV
8kxuLw3qONaFMaiMzJg0w/h2fcQ3DwCuCJV3WOl97P0lUkEmPBg0p/NMygM1H3A9
nv/f/wg0q/aQLpgPqUjgvHKYU2MBnn5JioK0iuISVBAWp8ecbYMjpGREks3En4xv
9FAI0uEZLhCtNi8sRQderk7zrDy5MMGHuQsEYLBpvnC/7UFX7OOEhjELICtPoW8R
YcBHzBbMzbkv9F6VimqRgod+6L+4s4FEybyUB+7rVIsDngkSU5pK2FJ4ZDtERJUX
PtFJZH8l2EQCTXlcWqv7cXWcygshOQBu8HYTzOIJS8yO0SId934PyHCAsBzjPXv8
Y9Z+gbqkiYVAOisUrIFaHndlrc6PDEE93e7WM6dMYHg/3h/BG9SBRn+NKwPnZitV
fVcRWTZ/50ELa4imPDNGXMnSuO8Hv1H8GhLd+k871odt+Xppwlc30tyKRTniMzud
oy0UR+2cpS+ycYhArDcDNrRWznsDjI1i71Itdz/Nlleu+tSV8OW8vhtx1Ty1uaU6
DZQq/2ngm948nZOzrYJkwdkKFK+akeViJXEKOvnOlbQZoP/39ZxqDCC11jXDGvmg
UB/rU+1C9Kg7M5kQ2b145lEo/cDZMt1vAIWNjoOwwvCUCGcTpAFOe0+zOwGBLtny
YjZWu9uVzm/hIUJZ9prQ4cmVKqmq36U4mkQPGjh0wq4e9H01Kc7naJ8pqM9SZHli
YoVJC3jKyRCVH/qjuOyxrta0+B62RIXR5Yq8fEW8wFitVpmKgAPq93i1wD/MyRuu
T3/7zkEAw9Zo6EnajGZE3aDJS+FX2sltHFAIc3SxgE4a/VAk92UB3O1K3c2YncIQ
wFAT3TSPD6sjU4z4cHdYy+60JIxmjaj0VR1SuNSAR0fxph/aoyREB9oySpK+omir
th3Ge9PEU3ktcVqEWpaOoMb0vlyQ7uE3puUx6RAgsSBIy0Zp2JQpL7OqN9KTVX/x
frsqq6gmtZ1SE2HFd8PPLeNWlfMYxK3XMqkJRTQz7FeboaDCsnPNIes2zqUvTzKO
ctnn1/ehtRFHlOrrKz+llPzzT7iFdFIe1u6K/zeWoMqA5vl9tRHc4j1GEn/fMstZ
G2j9LouPPB5nJLW3kHF2YOucPD/7owbJFPkOcMOBVh87/SPwHT5R783GxG6XKSJP
wwFVGDInyP262EYbKQz7O5GAJPvQ4ta3QvmeaLTqpKRkmCBpmJUYx7+oGq9JvIyy
VTzZBrwl2cEUs3mrSXxKmMgkaBNAYkvxuuHN6pST2tZHewXeUjbGFtqyXhjLi4Nx
iC4qipgu8d7x7djxra3VFO7eMEh3VkViBsgNM1eigdaZl1VtpOcR1LD2NS1hSGk1
7N1MpQHsJypRu/mtTZVHJ2XSeIsO2reaUCSnHcBBYfRlEMIf/J1Sfhhu2sRACUKH
3qJuYwWs5qYJPopOy1rZj6FiybLNf/Xm+oZL26xQUVxmbonzF6/bYCyg4fvsTqWx
b9GqHL6VF5W//VcwIVWJPFRAsCO8N3pD0pA2Nd7KyKP/LdzqY7amdjyGpSh2SDOc
TJV64cdfNPC8xMZVRpn8/pzsGAgg+VPo1Icf74+DOQ7pRURBKAu0mCOpgZ0OjBBZ
98B0Gx1+N3QCkOiQ1w65OTxj5wE9+CasDaq835jQjs8ziwrxRUGhuCBAdsfXFyOz
1asL/xWo13bR7xM6HkMEA+rlz5DHqddDWwZx0ymMcMIksNgrCAktIh/FEC2czLFB
1Qf6yAdrRWa9O6YBuyYyhl00O8VRzGk5icgISDYJF3fF86uIB3hVTSHAoXEiMjIH
kB976iOEfkoZ7DEIjAZvRTrVK1y/C/gbJcla4wapUf0mvtDZgXIcl+6Mw9/rs34h
gDqJ1o2AoBqS/25HE3RodW5SvlD0KM+7fRKOLs9l3PFcEIY1HPdW4HW74QvJ4ill
TnXllVq9mY7W+cSfkYVU9slRGOowRRFRAi2xLD6NwWD5nQZC3tTPltn3WIdo0fGB
mjUwUHxlODvSPfL643/i9/aIHIs4hs8HxVY03YfZk3I60GWOPoywjTOcvF+2vk2C
vz8yAuRHSCWD8OJUZnvziAGu6qx9KFQbiCjYXUL2ymiaP/PmPqZVyTN0bziyJuFd
k1ClIV9SBnHD1ZE26iqsPSlPugJwOtVOADEt/0YVlX75zYRsOboAy/WmYHi4evpF
b7bUssWzAQL3Ea8br8Jr3dFeQA+Ug/pF9FFQGzuPiWhl9YyuVkGsKN5XPPHYdF6t
TsmpkMHCCcy0OngUPP9l8Trmx/0VK/FAz9R9ndg1qb4PVao0ddrWKMk/poMOrYP7
2qiQlkyiFFlbJTREROMIWz57yP78lnsVXYRNxaJJB0IyP/0fAXLewb4Y7HcdjYj2
iEc9RV3RzQxQSyIXfk3pyc3Doi9R9Pt+tK2MEsfSwlD9aEgqCmQGRvKylXFQt3Ln
byw1ce7y3P4XWc87WBTSdiqtnq3LMohOww60l8r+hpCkbAWaAhQsdKJABUurSf0f
MJ7JG5KC2u9nquioWyNdUORIQdb9crTMlQiCORTzT8uidfwwbUJUYgbmMI/mcyFT
158tI9Fw21qB2ptWOldD1tCDZGGlcPv8/GglPuJs9XoQWIprAuxfJoH2Lzx+XrHZ
rZM6tuOGnZicwuQi7zSCInKoujDe1gnSbPcmFywgLlvZV0llNGxCrcDTNGRPo3Zj
EUkS4UgIpTS3g8lee0MoyxqhQji6bWKDzACjxM4Yw/r+daIyzcpBtBsgaxtEjNbG
l3rdv7JapXnSBEbFZQLv4OWFNOKXAgewGs9R26NjQLqXBAaXu3xhxdlzWFzY2XSm
QbC7wFdFzD526PKh/2WPlU9A0ywGtkfCrhio7cZroJoykpUD1J5m6bo7SXpkWYat
v22DCK6yyQMEKsS3PFqOV0HK+gTX5G81rfMmgk4nJyHZrCmQ0lPAaGU5Uzfqfq/6
ZmukWFtzMrbJY40S3ADXVA1taKD4izrjcaFHR6er7chmADc+c2kPdUNUWUJzDQHV
b40eetU5+qL61N8rKoyDkHZikywMHlHZUwjHXSmgTArnZHjS42AyoD3svJ9J8GbL
DijMMx4DkujT1aLwNi0N6MrIB2hTvuSXo2qwVgRT2Gtpixwi8s3n071wku0jhSCA
qg/zHngfm++ay+Njvp+VK4AaZ63wKDwZYAEb239Sxp6kpmoOs4M+0fTnWQe17BhI
6c5n3275kUip+toZ8OCrdNHaKlWeLfw8mg+4QFH6SifwTaqibjoat8ZFxiSOXKUB
163QpcnI2e05oEdS6pABerrL2bAday69pHHVNY5JwCpuCNfiwP/ZxsE+sWwdNxgj
MpdoTjsCg6PiPN/Uhd4XiRcbFFjQJvgErI1MQuUzuLZFUin9gSuKJt6w60NhzE+M
jY41tIAviEPtBCCvLBkk9uhW78x62a+ritjdeAH2ucdlReSVLgd2ynvjjRdvdGt8
AQN4Y8gmwgdVt6PJgIpKth5tZH+6MHu36qzyYmFvWbP14N1KBin96NYzVUXpZLAF
jIWF4bR61SCm+krWXRYj2Y7uDYCsYdmqQ3A5vGPON5/oUfuAs9Xp4LdLtL2YLq08
9czUtKY2E1BFkNlvM3a9yUyyTv7FvRzlcJ7+eDRIi18KsgUcHwk0nt4cBQa+ozkk
Esbb/SgHuH4ja0CcNFu5HPdhRoTy6yXDzHf1Ypmzg40SKZcwB1JmNwEcrflnaidY
qorqKUaHIuQZxNl+Vj8EW00LBbDqhODBzl5rs6R5Y6d7uZxI5HcUmwPko8Zn88hv
zbh1UKbwlZc/lf9cAJejBj5nJxj41HY+W7A3poFVJQv1IqHwHSh7TNfKpS0f49MR
dBCvrdnTtde+ordW15mcth9vs4otCwTThHokoHflRxCWd/LAZu4BsiNori26NuKh
oAFzObc82GHlj4ZrnYuUGVWY0iiDO2cH/x8K+rufhyiSKal+d36yjthtiZIMdXd1
MDid8TEFKbjNz5BWW1UkX+SeZqYGHkloWgFkmckh1+FGn51DNQJt4pk5oaZOoD1I
JSS8ltvPoqQ4jqNWG2flmESiSu2Uk+bQCXVAeptqEWL8QCZ5cSuT0fVRpTfQuOMf
vdfbHQ6ATjLaK/cBBpFU/nNi5S4Jwz4zzhFNimlLMTXQnyHY4vYFWR6MOczfIJX2
q5HL+nL+bslVqUu9BShw58Di+Z8THDrU7ftPID+Su/tZ4Elus9CfimxCH6Yez719
BOm+RrqkuSLWMSx5hceMSevWhl97IZp6KJfI/K4dm2eKbKcfSja2LAT1OPO54dpM
vqYEqbUT8bgEYRJq/dt4P+QUO/nhiA1qc3LJkFa/FKOBp9uxnu4qRT8A1BIECLm/
mHHKhfs0ScIfID0u8UujuPGxoVh6cDipoMTVAfZ2Mgo6T7VAjqPKLOEpSEV3XRIn
q7APOqPPBMThWbnYupHEBdItnxt4nvRWRWKSzGf8Pdnmt8M5gvKy2V3FpdPIhkJj
Y8tsB8KO2ejoevsC3qIA11FiiJJx1rmw4TcLuG0qQoKa2yVGTcRIHB8+RJ0O4ST8
0PsM4TTz+Ud+3TVpyOkZBuBlqbJAhLp9gJqB+DZTaVPElK+/ZJAm81610e9Z06UT
bRei2xauPVvA9lZl5f5GxICa315Glj3O14BSi0gDcxYf7/+xfwO7XDydKhBa1c0m
ODkCwAckBYTU8S9YkGIHqVeqxfPOChUglLkVXlihpBrvIHKJELmn1yw50eco+jfi
uYm7wtLrgRyHQ7s5vjyZbInoW+bSX5IiIuNDQlS3byNPliIlCGo4oHwdUONpjrbH
n1Q0Mm7oxm2YVrXDX0zqIuTkeXr3cuCSexwYMsz2HwuLVNRmylRXRCYKj2PEodlg
RixPjiRQm9GWoeFlYQiN0S6tMi+zLbymtq61N+phUJ3OUjL+dBqKv15N6fsoiJzp
6Q18ilzOXZpbwm06nkHNfvyOtURH0kNkrt3gvsBzlwgDSj9HVwTkePWD0ryOy2CP
7sqnfLtL+gG4Bi8Lu0c+CUMCa3+9nfgZPby64FIvbiPKyczVFrb3dRfVXMi8X463
9ZdE+ZZq63H/KeCs3Y2fRZ4Tv4iB+7XETNgA/vb6dsPJzqhvxErqwAS0UAn/1cpY
Z7cbnAdtU6HbNXywNeMyImBovTE0o9lVb75KPOl7IrnvF8zdmH2mKbRUkrSE7yG+
1BQsjiZpm35VOXfVLOQCYKZHeBikyu7i9ZKkEYToL7NNJMEf9NWd/2OLxLujJPKK
i/r3SCmUPCVi8NATWcbLzvA8VAyIg6xlWqmtLm4OPcbdS7iWUudwCTCWifJ9qizS
tK0KNEjTYyswRfUD9S9nxEbHqlOjLTERCrMTxksYerVGExZM6sYd/odx8vUSpQhs
4U20NdiIeiqvNlSnJ4UFSNSs9uuUsEDN3mY79ZLRqeU512wcjOB+HKu7a9/Hz+mf
/ewPbceDOhEeFuQ9IQ5cP+VoX6qABGvClQXGaP0jsdXFMqRcT4UOujY9uF23ojIz
Mnq6g02zXdV3dXP8a94iyUJdliVyZcxjAbz23t7zVSA1FP+onZWBStaojvqUEwGp
gvFE2tiC9u9S3j8/qY+epMT3ywsLj9VYpaFXjBAFE6cLje67wbYKVAIfSzm5Orx7
ExQAVdlgafFzueCdJ0ia/l7OPadTF/wD7MsQxtv96u0uoCPeRD8+JmPzAtPK7GIC
X8iBSTzxs0EaMvoKfI7myYWf150cZnbyDvkN7Dgf5eV4/qIyjreE05q8hffDeooo
zkVp6kAEVum91GNmYCuTv3PVxBDeEgipjo8piv1YlSfA6EMADBfZ2PJvV+89r8Jq
07S9Ajsfar+MDwRW4vYVRLUml6UaNdhn8k79JDT5gUN5GHQ000NfbF48Huyhi9ax
ym+DWAchZIV1lRLone+QVDRPBQbDt6Py1FrrlRIvvvxMptAQy/gvLyJWVErd8BuQ
wQPJBOFleiDkzF4qPMfR2GPAl3tkIzXaoAOPNdqViyRtIQMDOKaBdeOIFt2KAaJb
Yf5Ka8NL9K+QUtgp/Ypnw3+SzKR2/1EmvneWnsKwh7TOltL+clvzj8Qz0DJrfvFd
vpdqziO/5QtImksEzqCvVZ7QjRJ+iwJ8Hf7Vsy1BSULsUCfx5cf/6vEZffcfLJCI
fLUKVf2jqr/ogL+j6Vo1q4dhxk8/ZUAZTZFdXCW6I/fejIWq8FVTpxhazNp/yAYQ
3p7m9HD6UKrI7FWF5YSwcAvuoWKqIPertbNAvip0Y10+ly09i0SpvgvmnqOdz5aY
+MHBbBWFEBqBplOd28Yqzc0tt5VLcA+kY9tyDUvRLW2Jxj/97q7rcGOyAPL3zAsW
oNCmA/UqcdvB9b/E+wgVRiFGUChDTKbUo9tbElSj1I+q/qi3aw33bXovblPcQEtN
WLdTuzvi6YZcYDgmRARLp4QO3bW6vEDJU4GYmotU1x9EAlsb24PSiuPrP3HBA7Ei
imW/2y24Nc2kQ/jmG2eu4Mdrj3NLx62vZXvJeIipbWhIsMRctM6MXQ/+SkMp3Xht
rVTFv4qF4NqLwci1wXq9VaB35ClhdwLH+hCW60aCRCo6gwzKo1HOJWU8kthhyZKl
G/ecqlIu5gJpt9WSdrzP+ovdgzFtZOdUfv6dxD5JEIzrUfqw7XuLaqfHBWjfW7B/
prZmd5Cb9/B7NUDWd+lGmZkdCq+9txXSKxKUNSzvNVOAIul41YwoLa47RD35wKGQ
2Rqz+Ol/HLV6Cfb06Z1CT/jYRTco3823LKjfvoFxDtvKOuVfx9E7HfWhcEn2R/9s
pQqY1vUJEBMtbRTOV4JdQpQO76QMGgFbqoWANRqomJiA9dl1CRud8aMAcNuMaxDK
ZL9Zy9QJ9TSTDyJzuTY/ZDdeDqG0JB1VgjwICfbmCQ2qE2nBCygS5kZj1ydCEsUJ
TedYHIs4OVNlOL33P6XMj5QhmNvPh37UOL8EWy8N0F2GSw4fnzzytOUL+9789DqU
eC6OllqnF7XfzW0RjBh7M0Xwi3AuA7veiHSaGdtB68v61DK9bjwL0/0xOpzKjgv9
3ANSdjKYR0hDkuOVpxpyJecyxrsrvb/qS/RUfFWTrOIP7V0KCwzI2FqusgDfvWu8
jvMCJfTCtgjtcoKq58lzD2/V9UHQTtmokNNi4kC6QgatKeT90xClVSfZtD96zVIR
8xrRwv+NlDZIiAD7G5isHvGFDMsQK2Yjj/d1y2PWmMgnYFv2z2ewWTeISjEDJIdg
RYHYQJT7b193qAg1Uw2MPsrxEzwPt42rIL1AGIK7pLmNh+lRkyNtZE7TrgLIoi9i
G7JmV4eiiriGKkyBJfXli2X79CfJxy/EQIIOJaUG0IQotCurzddvqeFpo6ZDRj12
TDOwBNCd9MKjQVWAm324qVfTMKexxBIxDHwsszWfFFj4A0xX3q3lBuS/rok9l1bo
Dv8zHO0WL0mFrgD5p/DMk3+LbO8DiAzYzH4GEKnXD+EdPpiGd7NX+Lf6S5mAByxo
VM/gcJ0oqdSzJO4hBKcl9PzyefpIPNX63C8a/qQzPlXCkyBJEoxPynPA1W49U5v7
UUhxYlWDfWC/vZf90dHhOFgIS7MX/TpM8HRASEk8WqFDtXz1ojbHR7odgQbb/Uta
aPzEnMpQY29WtO7FKetXcOFu56x0z+pvBpRpOaKGz5akkiFpoFjgvAzb1KlMPIGd
5gLJoSAcAO+cna5oG3MODdxVfOSHLQMIkfaY46bkw15r/jgRh3eGRiJpHsGAcpbk
WChhB4Eyjk838sz40AXb+1v2qBgXiijeCFk70hW2IqOJVJl9M7epVkzRlrzawdnU
0kCmwWKcFr4ePTB31qmRoh1c39pXKR0c9f9iRIj4Oyt7Z9qgBCK2o/Fuhz8smpCK
v1sOrWyGT9cCKhPQChHf7OJ2tNIBoPU3FYOv0kh9VtnB/+A6MyWkcW+93C/52TqO
ZmKqPmBcydp+oY31VMr5oMjqzRZ+6Hx7+PfkzTe66+WXS47Chb4L2QXDRzXCcD9k
fIMqcpCcwFCqV/tjF7+6sMseCHcX+fsQXGJ1Fw7JNs0NC68kPZRmv4tketQFvEXa
9Fsrpeh9YWEJJ6eQFLtRdCywDE6HoABMqPLh/AWHa/dsiFgjv8nc9KkvliHXfW32
OtSHSoPzNz66EOHxc5awNqR2Frh9K0bqOKJiD2+uiNp1pZ5woUtHO4TYBBugQGLi
vHEsinOOI4PxDlzL6AM62qQczjH/jf40iNN7OGCpz1w4ZcymrHd/tbE9r1BPvev0
i4CAYNcwzlXxYwkqqH+LO0rEJpkXTcesS8RAHZnExxjyFUJAg8Tf/kOVzE8VVlfM
T5d2Wx4YuZ8d8dsypK7X4ePfkX+LEC8JlPnupI2VcqsPFAf9EyauTX0SKyETo0CL
37LXTGg+h2/GiQFkS01J5IPohvaGFZSrJ5AGerwzIklPP5ZrC4p23brDUjQZ6gMP
umhIYo1Djav22iFMesTZeCdYSq5x/jgfqd0xgsNgL7miKD11ViHDCgLo7Hwjjk6H
zfxYWCuzq9PAzEV/3cWA0oaiiNV5JHsSNc1Ezizx94Tu3Zqm6nAASwe3vjoAwieo
2jFK4Mjn0EfBDUNrXydh55uI34jjByNaj/QuZbU7tglsoP0Uv4t8dONuHFACjrIY
NYNArLU0s6YyfZKMk7zl54UAy0loOMjfYAYI7ENlvwyue3o3gMhpboaBjElxruRi
LTKlFZi+KNf3TBAh58KrS81KWlb3DnHLOo+5hwdWBvtxoQcfAXdTOzqAMFipqlmi
Yh8rJp+TeqxDc+fEji4cStyk1o8YQxwoEfBK56aktHqHXQ9i7DDYK+MH+MEfsATH
2i6QC0UEgQ3gz18O07ktqR1/lk/NRfYq0OSAlUci7qcF2soMtTETBTx0755ic3cW
WFNZsgKz2L4vetjr/5D+u/P/2ULCKLekxHgLYAwf51DWrq24eA3QkczYe8fEXXCN
NKNLOHS6uP9RWpkHEFpne6/QmSvuuVlomrhBczmZ0iXNkF05F34S5BJ5wleAgT8q
iB0s8fBDIDwO9BKsPHicCGYgl+QYy3apAopFQ12Rag3+NO1/wZgdBP8KyQupyc30
Fudq3mUh+H02aZ6di9jFLG+bwPAyteoTWhwRlvylhZp7fSCCKLfqInyymhRQEEDZ
e5lhItjNs82dHpIV9CMrH22JUTJTMLiZXJEao3SAYLCbZPGGLjOeNr40uxjsBsYP
8aq20+NhtYYSJJJf185Ily0Dpq058IRAa8yomyt9OXJQ2PQYyjZXTNen89ACUtyH
vJf+pX2fOSC6rzwyW6bvD8xQCLBVNeiOVlXQtGyc4CiQxL24SyJtxnlYBzdYxE6Q
aBMkB5bncquxg2g262PYD4Z4tnn9AC3zdiMIfmWLlzgjE+QBjd+gyIAtjxxn/DJV
JUOjiosTCUsCz37J20lLsPd7QmgfwCL5Lyq1kE9FnsCZV1aLRR2wZM41IZeVwwQd
Dazig74T90HjnkEz8Wee4DgQH1k0nNhCNkmaZk123ETHSjRTqjJgOLs+t8b2gC73
vw70MVeZEdU+N0sqAC8W8yVatZLIWvho6IfOxy6WPQosaSiBXOeGO9T1sPA2sG08
JlwMLQvNRLsbhpISRWgXLwy0ukrXKZ4B24vwX8YVNhhVeo6WjsxibjEGrTflMqVg
Dk+wZ6j9kT0rhbH3gGnjUaDlSaYlXzcpwZQF4AtOeOWNXRIrhe3QU0faYWKfZWYt
ZY3Fw60BttryPYRjIGUZfQ683Ac0UTMs1YF5JAoN05ux+VU5IQvos5g/GwMvFa6r
5buJWTr6qiGOVbzlPSpYchCF8TC3jnAw2JymQ1frqEx6uR3giLbe1aEa+JtTdsQ2
WgTDERZtN1h4rNqGdpyWPpmGXAQ9CCt1Em3Gh2nPgdJKnBBKorBqHfIwCCTf4zuW
dC8fZ6Ex2WWDUnZdBv9FAExmGQV1bb/BLbKYPuYCL+/ngsXB7ZQSfHeWO6xcY0bl
XDW3MSMEPyoEIii9Hxolrltbti6Uz/kLCeNK6krLKBqoBgS7r8meSwfX7kqxA0iM
ebDzi6cNwCS04G4jkJOnxuiAHBBMCj/I850KqGtzxeAb0XWcezZ3mYMLRbwwIfiu
bb1CKgNDnRCF2hIuPJLyR0uuFFUPv0TtOhgPsAQqdb3DeuxkEWZDaN7d7eGNCeb2
tNiaPFMVLKeheoQdcfVJoyPfEcIWiziXoA/SoD4dQD3kBIUxSlxPYWiX1u1cdPdN
kA86N07RShtdtrTm+F+nKtLLBByEhyGw+fAPRYsLCKmCzCwF4csZ+wbcpQaZeqvH
2SaQbOB1pNahfoIxGDW4F7RtC+qHtHhv+wUACgPUFozZ49KK0xOxm8cUe0qNMB5e
JTL9PqVek3FDpmjSUCrFTPWWoQ5UxYEk5wD4A6dEYBGgKDBHL02SP42DZEuz67RV
rvphpU6dq9JmcRnEzLHnqYt1PFUI0fXnjCBnodF9YqJVAG3VWvtmfpWezgjoxvuO
9oL/u3JKuq7CKnNBvs9SiXmT8Rx19P/rgEmNkx7wqSjSa0cqvS6XGq9TC+3SMPrc
bphW0zToQ3mdO+JpU/e6+Sqglv93v7ANA71EWtA8MlO4GHCFAg5QzWphDNurU6Ny
sQck1vrWhhPUfeSgW4ow2IBm7fYgoACUmpKWgP8rHDIYx9Kb5vD9mDmKKRs/RZUB
dQzleIvY36qxwMhJoLmCBG5CpDguyZwG+fDcZMpqn+yytqujdA9fA8ne2U822ri0
ob4S0vAQ0yBedVTij5q+UpQ2D2gXeBJYy35eIR2CQwR4I+HH+aYskA0FCexSJPRQ
3by1jLcOv7LTGf4+DF3VnaIMf9+v+H9eHSF7FwxfoHvs+4m8x/qp7LnBAvmlaof9
BBGCVbu+hukEvn0YqGbvAPYLELr5j0n97shd85xoEeRrGfrL6ll3RM0OiNN1gzDU
P0cfK4RxloZVAVIXzQvgIUtJj7DS4HIKpww6q+KetbbpGNARSr8zxrvTED32ggQs
VGpZa7VGwVABe9pw6+oSYVtB9RR6C+fWengNluUUEtSAuYrJ2C3d5A28KJYw5esV
2dfvcpvhC0hUP4LOuX5qPR3FbskQkH+0StVQMcj8K6hl18gW/L5vp/dTNFct2r14
wZ/6uwtiEVNXHeJyCUvpRnIc1ZBwKSMSDPCh1m6dRO/BofnC65I3NOm1G6KiriL4
aS/2hCPF3bXWuBsVqIkxarIxDYh7/fTnq9kT7+SsNEhAL0bdzXb34igb51NolZ5X
Khw8prXr23bEsrCnSTAwEDlT5SYeQ8Qsnm3nneV/VfVmm0XdoYU57gKc+9O8GtfN
F/HESH1vCYPFQ+pFscn54SpbLy/9IP8RAqampcbWryp51FxVxdy/2AT8amY6/xP4
kdHUFfvMNnw4QIuJXqZLuXKgtBO9FM9d/b1/Wmx4+l9cmpb2TRFMRKa6yV5NWC8J
Uex7wii50sgrPfbejDqmVpmCf3TASDEAJQyMbLGZV2EcbP6odKljCHIUlTg+UExS
4Ewbv05KIuWd8W+qbxyeqqN6SRkr4ucL2zHPab+qecCHAALtU/XthJiR1pBAS5wU
r33lUZMchhakbuGE8OB4W2ja5kxJG5AgLomfymPLg6nck4o81V8cG6C6OVaDUnd7
3LASWsuZWAZ5NGMtdgGxLtD0ZCdbPAMgc+hfNW6cuwaCMv00G9jvPSZ/KEeNxHhQ
MEXxTb/6YDvYR17DmH869hAngn8CPHTZqKXVaBCF4HJxjl2Mqkc+eh00JZih7OaV
kywINF0Bx3DR/uTE1CmZWON2gV+7zA4WyOP53GrJ6e47DWYoVtMyCAYjgzn0rH+5
IIN9ge/seJECMuvc738z+DRUJF5315dpbGHn3FboIHI6ix1lcexM3Ze+CN3uJLLm
IR4jS1PT+bjC6jEzuWJUxI5tQUuqz/REfi5jCUxX/RrjZof3ZRDJ4QTpINcx4Syl
nkh3r2LM5akI0RuqOpA8KjNVPfcz2908MookN4B0QZjvUoXj7ccuk9CWdxMpb1DY
NmTVL1lJGw3qWMIc3lSIvASNxyyNGaSUy9qeoUk+rJrlVMZ4P91+nQ+KFd22aVSf
vrZfcbkl76GfBylx22Mw0hYjmMzXmerguHohB67GxKEpoZgRAxSnS5cV4VUZhuWc
1uR7PCiOv2+VyaM2dxQmGrOfczINopG0KgrQAt0s5KLivyMuqDlg51POnpyAWrT7
N502MtE1iF1pDkteSzcroV+nFf+TIylA4ygIJ94Gd5c0Eaqg+pCYb8BiWT6TZ+dt
IcpBbPgjZQuOefetba5x/3cOIoA/0YObNHNCSMNULYbLNORs3uig9Iy97Yo0BWfy
o3AzRuXx79XmQVj2PvvasKL6je91zkcbKqkkUkFMd+L3ogBgMuZ8ywEm89VNGhdC
cj+7pQZ0RIhZnYSFVmw7jH1RS2+tNFpKJAiTDs+NKAz4aOmDYlgKVGSGugHWFM0V
koZPDSeuEJnyRTEm5EIsRZMFdEZbkNtLthZa7BpH8atSbMBlbsVzwwmR0cgQypzE
uTYhrEH3487qrpoGQ+gVcxE0YmrSZbNmF2DSuL/kabOx4w9v6mwTrixMLlzkBf4C
aNF5tY+Q/T6gO5MUs1Xr1wnMx/2j8hqus1tkz+anemrJ7iGkhBi3v8/BbjHFekJa
8v0kyCgEN7+NiZFRJqFkLtcEJ6VMr1YTyiO8xTo8+F8HDfgJi/JTdHOSY7vRHY7l
jVzUgzodjZ2dxjYLicQk+0EluiA3cgB0ZE4ZzWHqtJfjOoaCyqKWk7oJQQgk7eIs
wyuIicKklh7L6vmmmoSiNS1hiY0PziqAhAEBBzCrJ1OlxyUYqedvvTi7pQ4UG9dr
UP8C9aduXCC07S4+Yf7d/Ftr4c4ddsl4el/zZbNeKzs+uomgae5WBKPKVZggxFaK
8AbFSOlrUm8jVRm0rQ4/kQ1vEquUaCOaGoF9ofJi50kllj+2rhoW726HjuOZaD3W
x0+Dge0q+M4M78KNBXrJUlpmhT07+VaqkPAg68brs1iANM8WRLS8NQjR0n/3CBF1
6dB2+ZHnRy+Qfzf6SBS++/cQCzT+PqNaiCjgoQ7vH+NMKBZvkQGcwWKC4dblHDfo
qVEugzjPyiIbXVJRLjFBejn432exxeZK5VDuNNtv+gbM89ri1V4iBMwvko8BRiZO
mb/TE3G0HVLY5H5DaRAor0dGV2DXQY7+8f1H67PJMPhG+D7ZGpeIMlyCMq6B8mun
QB2EL/s98z1K1DDSa5aryO4xTwekSz3M8kivvCwSQCNDUiQ+2CqnkKRHPo642m4Q
LeoLMnLRgUyKRPUGfDAyWLixi5HdUAZtqKDLC8BLVynBRNIi56irb0rIA1WLPUhg
/Xp8QKMCozCRaJuAtlVzDqCZCxNRHsVNghVI8xfoCHrLUQPWc/zrDxvRoZmpCWPT
1BHVOulyYY0nDknCpy+U2Hpjj/1P/FSta+xFxK5DOInm877TLSp4UUEndbEGBdYH
M3zIzke/TvlEoJFqAQu6gTZo/jOmufVV6ePgPEJ9aK6CDpVWuRW/zZX8IuTPey6A
e8YFSeIcKyVDme8KtPZAUMiemtrmVGAMG8A9xfYocj/RRfR5wY90Mlq0vVixNlAK
GI9KEja6wSJw8zMPbjuJgn0PGo2LQQxx0EqAZBq0ZkoWCRg6YWm5ApGI2U1dLwe0
iU38kTXkOABhM9ew3hny6fJFABi8+s0DfpMHioL8x6JvzjZE3e2X6ImdjDFxccC4
LiRjbWf9gmjUyR/5G59EXy9Y4h6SwLg0P1OaqrWDxABZMEsnp/dgRnYvc1L+JiUG
HfIeZfINj639AOZZ8YRntK2oXzvWFvWRAvuvMNWP9s36LZv/M0rshhIvYgYMWJ3X
i/ibzzdnkDW59/pZPcJlp2nUJZxKAu+66qGEUa4hI4t6dAid/UtC0ki5nto6KtVt
seBeguiM6EWd4NC98FbXu9RUTw34sp9g90Vhzji6XRkKguMtN/ORU/N6veg6s121
hBSECKc3Bi/Hscq+P7qz/3squvuKa/ac3/dhuf7hXh9Hav17Di6K8l9yO08fQpsD
0SYsJJEDnYyma/ebHpoM1sC6KeEcmbNLNJ3B1BGscXAAQmZ4VGXr3aUhgsPUMb1q
vez0q5S/YVL8Py2VGw4CSFD5TnThFl5GQ6jtbXVU+5BET0pfGTo5T34wYbRGqoaD
G8ThLIlSxwMKUtWuzlR6ka9SZoAci/PHRRzP45HV2FoYyTIPdwkvzmBDfKbKsG0C
XWtVwOgzAex+MoFWqy3Xk7ou4Rre9+f5pYKFkaX+JJHywGddLN1MO0w0X5YtP2G8
r5pSDeWl04Gx1n6XSTEmlwi//+6geWUzCB9tB0IO41E6llODg5ABZi9NfJLDZAqw
8vvUxw0qI3hQ6rgJIG8PVF+//aTy8RT0UMgyQqLFJJjtC+pHx+1OLnZtE3f0xEYd
pPx5nx68G6DUS5q4ccXpmxuk+LQ4q20v5KSqciRONrJ9KhyMiF3KoWIDEszV+HGX
q3DJOojhIZr5+AewNA+xuz2yrYGdGpFVrNDpSDU4Tya3sc1Q58EqqfMUys6m/qM9
7TeaenckjYxy89aVhnBZL+ekO8tgALxFpjzQ3Q4+pQMvZILGnKJld2varjVgBHqm
W8WRosQfDoHIk9hjmeOKaQjV38TiNtOegoG+mrrlPyYGFcYnblbsxPhTFEkNYqgj
5T2pudVumdxX5MXMEnxwFnG2zbL7R/FYPcCCWyDzzPvFr83Xui8fXSTzlp+BJD/j
yo9pc81cBZZwoC5WM3N7ktzBtgIlL/320o/qytA1erTgS8qmLpx96Ql/FLRHy0bS
HRLrNrh+gmxuQowqRvsGyuCkOWprvR1b2PX6NC2aXRrt9yFyVgRSzzVLbqTVGJcq
CqzpDvAUECkTOUUrwR0OndiQ9vAu4xjafK46e13g6k2IaLoW/GsMO+rUILfhikQd
MrgZ/RFyuYZXFxKaGZUYxFd8ETzoLYrYQ9jogZPILoYEMfUJfM6aZxIO2esMuD+T
j/ijtZ/eQH9jfwIgOd/44MXGhzR1kgiqFxAGEgcWXbnzWNUdBS6O0oIpk0lmMdtR
NaWy+T4BvXLVPCMMC7lBgrZQS00jEPCbuXH1kLTtE6gsasBuED6YTfvDBBNZTdG/
ChGu+CbpZmS2mynK8+PcYKbQiXcCzClhVdinEW9DebMyKIs3AJsHT9cb1B92J/id
PFUhewQ9i9cbbFLmw5ghnFwImA0jnpIGKLk8rvQNAjb2dvmfyhwJ2JdbV/EoF8CY
Rd4Z08poiM/CM5SFq/J4BLY/fyPiXhNqye9Nb0dbvkoCtb4ll6wovdsqqWcx89J+
n7MWiCyuzE793UpG79DEM/jVmELY7yFPLzK245DKHGvRMv88YJpZAj86OgeHq3AR
0SWZJ8HbjxBjLIPeV/zAgkRM3VDM12hlrlG5124XWZ6rtxio9aP98Js/2/qjjmGP
FJPqglJjekXRV5McTvNZhJS60wzDg3vYSZbmL2jEUf+N3PyI9iVBTURDVz5yseW1
pi8Pzpb5Kveo8u8lhhwe0SyYOaJpHOLG6bcK+qo9DPqqBvMo6vo0FibT/w57ZZzP
pYIS83fGs4izI/UxWt1ltgls5E6qzNTjlccSPO6J4wQ1Wi/kAdKdM6K81gt9JsI9
RK8bunFr5MnbUIs7kwZKUP9KQbLSFOk1WLV+E7Rhho1HIhcMhKsNg01H+gfy1RfP
IS8rOwqfV/us6N9O39tG5gOe8rL+P3T20+F4YUutB5jXJMBXVI0GixuzQB8WTfZO
DQxl6BosdQ93FAvNJH6m+ia092KEs4fn0Me5GKj0o95nH+U9T3t+iuadAlzRGkOW
pbUMqSRzu6bP2W4LASay+j3DAKMn4SE6zS+tvWsVDnhDLNjdoiPkOiJXl+XwtpYO
K8jEekp7F7uiaS/gD+4Lo7MPUUm0bodE1y2rXJ88gLip8prT/GTCv445F4mjH8gg
l2h/hADRvEc4EqjLSTtJ73Smf4Q5uYcc/pVYnxxSSk4B//ZjckFWaxyC0Zv4/LkX
dHW4g+7qbnte1151mMi8QZGRI34m6aLcdBAYW3TI7w0kSMXSWSP2drWJGdzUODIA
EdfzMr3rASe21IyFZnBYGc81HIWc13tkDpPBHSpuy5KefW1Ndm8nW/wudrpCM3di
ICfrlnm/nlgWEQGxmkKgM6Fl4uWIv1YKVqMRW2De1dOsr9+M3XIsEKDlIL6C+DpT
C2g5K6w3zujMhhouZhZFyGhr8KEWkjR7JN3FOJo7kq8olmXr8V2ROa2NbvOlM6Mg
uqcgpjHmlanUVjQJeHnclmCc6C/Zg4uK4LAQ3juLHENdEqOTTEFSOW2Ty5zdZcys
TQzLOt5Rusb+erO4gvEFSUKawdrL4Zs8r+mmMjNOYv+tYmhaCvEjCwHi7v1BrTeh
7fhCrxYO9fJRynWYiPtQmpI0dwKCsWwWB8FmfFK6DN+yesnsiVmxU1CtLaIxzxz4
dPLy8zLMaY6Jbn9b0WjzC/1/LudUsVduwipsJZ1c7jX4CzFMiLg+x0jalnuzAkvQ
Zj9EBYtRFe6Gl0D77qOi0z2zHgVG9KAU4m1zZX0V6h7U3fnBcneAFLH5WmShSGRl
E3WFBw7yk/RCcdC/52X/Q55nC7sndgOutrcS7drdbzPAugePvMJokpPnZyXyzpZx
dqswrSyWD46Ax3jh64FMTo5/Tl+FTicv5gcAZb2gdoA+WZt5TInvPSX79/dCshYw
j1a1XcDPrKJG+ek2XrjGnjlpgTpjcmA1GOPV001bneDvHVALb9ETQOtl2vJldHB9
E/cbd9WvE70FjZG5aY/i0b1Nn+rvJZmgmy/Gl39i59w4l43Aa0yL6UGpmDbom99b
D5gBD3ycb5HQl3lQXLPKFeuQ0bUpfVQP1Pj3YvaZDCCWPmM6RV9Unx6hxGn0YVwt
15x11/pGjSEAGT3pIQf04foZJPGgSnPSisv8Fnr2o7etz/mYb2WFiJIm42RB82Z0
W1Geo5e2d+eK8CWS2Z1Tou7XKp9fX6qQvfAazc5QWznbHYudVk2wJpLxLztgIzde
yNu2XhPUL7M98tSWruetZoSebQbUHkOc9C/VtCZR0iXv3R9l9eMmatELSEoT3iKb
NMgWR1TYnjV34yGDBQ7Ql1NhoWQ5y1BXS7bxS0KezeOMPiueN6Eo2kFOvGvAAXvI
W2Fqy0WEyVkuRm8qzTCkeOQQ2RQP0OWVAEMtI2T6olMe7xLVs5WALS4cmytcndnl
ujbPw8gEZ10GBd8gecFLGw3fWX+VcF/VQPDys4/bcqGrnDNAMWXUewBOhlFHJolf
GJG7mOJ4TPFKeQniwS9KzJjhpu0n4uYgl4rghI/wBDO+JQzZWZjFzoYdoDyAtCEN
V7kJVmbUZtraNNDjV0mtdaN9NVOYVTyn0Jvbvr2jd8KPheKWGdWSY4UpNm5ZQBzY
wvwF+E9toJ5UQgheG20T2pGAwge6mpaqGdLZLPN+T3atR7kWAYR95LZDha2Sz1Tg
Qx8W93G/OKdpDVOcfJpz0hC+yh5+BfbtuMbcApuw+UkkhLBTnIIy9ZkDTHqN35Ai
4C9aTXRCHO3xFgVfqe6cz8qa1lYuOdHobSsuVs3GkBu8kKCTaxuNcx0gKDXNlnyO
fmwnxchUqxsf6l5ZUbpSS+CwGDPnqz732CZSAckhMA0F/VJwCrAB/g+SkgbtL8X3
kg/cKtsTq4rLeAaAHPGDqq9KcqV0WtkQB6Zaaq8lvKpDW+dWGZRbPGCQAlykdVxf
6uzVLKDpq433C1s1TqLSfjePg5iL5ntNRHGRyK1HDnD2V5+myUi/77LKWJ1pBbqb
ujXiXtpkg6yYTEiO7bsavDkPQcVAc9gDYYFX3moTLfHwewN8kQ9t/QcrtSw3t6Zo
KfG8Rx/VQa892yoPK1AFNEu/5WU3nno9OI7XdxgfNW1J7oEI3dHs1osfW6pD4o0V
hDZLFWMfk/GLnOzkMt6DUFTg5wOaxuFD+fK46HS7Y0wIXWWJrQMseOXq/FWR9FJT
v9dYh30Aq6tTVismtIVVWH8pJPqEbiyzdsXr6gqKr8beS6VYY3gJwnswgUQQFxvM
/3SjDPLQR8PgLI1N/umxOx/w3pkkHxwSW4tETaiN47X53TT4SUIjLL5EM3xN/M4S
G2lGmVrcPgCb64JbRtcT//wwWs5ngZSmgZOa2NT9Zq+gme4l2WZjS44P0eZvOxtI
GzrClbkBfUVaHP+/cAnjMMyO0iZySSV8aUKyP9eK9tN77qW65ds74FZZiIF8PZx1
dLCocL+qUmXc38suGhCq72vDRw9Tzm6EPpwSqievbuJh+o4CyYZIgss3HbjBRj/a
hEjOqJ6X4VFdL6rt7Lw5TrvFUhuBpqI5CloFpCznomWY/UcZHcmXkDUV9vNuzPlt
HIV5ywK4jky5ho21/nx1cl/eQo6QoJq3TlThGFzdrVmqzjAIE3D6x5xz3mpKjEKz
op8Ugx5Rkm44BbU5BoEhB827updA+ACQFgaYpu6Qili+BZy4q2CMMYWgJzxcXzeU
IgrWAZXGGMlBiRdAey6tQuYgVXaV0XsnIWY9JEssl71FOOCktvTsYolV0BOz0Exc
Ts6Kxu/2tSprySaGGMwjC5h1xm1Mo21xK5c2ZNEMrdMyCRKdK/hTM3RLTdJBcXRl
IgB1XtKhAP0+vP+wK2E7STaU/N2xppn8w8tX+spIrMPIiZhhfv4qH4puUmlr7zZk
/bX3nkZQV15L+6cs/1IowV114AZoaYqH5JO3CPiU8KhlZJ0aymRgBxS1sncXXT5L
g3/ohqkN4RIBOfmlpeW3ZuAXRLgbFAxEf3dPGIMCF91BRikndgXEsIuIKar/biDa
85W3ezvchZ7PVzaK3ocVyMEvK7P13SB/Pr/bajjuX+pvzyKwLm5pdzAZnl3tMEDf
w8Z669fAOZICkmilS8Pw4Ixckk2snlLLzVD/tgYeL8KmFBETvl7oX+YH2FPzNAwx
Bef9fNYoRWU5Lu+n2f79zLsC8hwqNes64GnoT42zoPIDjiRZO/uP+kUzSq0pHIJE
LDeL8tI8PIZ75wnnjB+Z55sd1f/EGZvp4Y7IoF+hjroRv7CTjcrcC3VnVsB9Swba
86J7QfmPz1XGoK+Exbhg77MXXOyzmjLS0ktWWmK2f7a2mjNILc01eMKwXaP3oxbW
KCDjDflo+alEnrDXyVMH9+3Erv64ZB6p83eIn7kQ7qRBYppIqGNrpg2EmMWtRd8s
mw83tTPs4l/7vMqRPLvlEbwZLgZJIdvGsn2wlcnx+VwE7ClphnKXlJdUC8+bk1/p
GOFT3DujbnJ+DBcrF8PeR4se5/c18ZeuoQ8VMFtS+aFTQekSyXeYritjzxTJpmUb
vJLY9pjjSq79lAm+FnytPRuzrl0i9taF9iKFPzFyLaSI7o8akB9LAePRMOVLVskZ
zNuTHxdJW9DJRTKIvQZ+2WCy9RNzIj63iJhrOq3Xfry/tE5spE6/bGmG47F6Ukf4
/CAF47323gVBx70kzw498ccubN//dgN9KvKPOgxQHO230CDF0vtoP95D/ib76Lan
pYf2xS9rNU1ftVVPDlUNLQFTJNIq2pfdHH96AnoCye3eGF4aAY4cVgLFPG1wC/eb
J+G9ABcjq4GJwcRFOEjaWAKN14HPPIQAo3e3Z5ph+IIdlAGYD5W2AKuhhde8lwCU
`protect END_PROTECTED
