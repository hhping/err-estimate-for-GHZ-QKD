`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0SIfhEaE+SA5y6Ho2O8sUvPJ8uRopUxx73GTzWU1pCIetz1qsJTluxdrgVfKsul+
0N+6JdStTIEJ2ktZutNuZL8Z8k5JLyF+k5GmNSk7Z3ILYAr93jY1rze00+ap6yzS
3GUQZun81n232zmweLiNPtAer/v+Aa3rqLsfGfSo8pU9cPlnpWkYSESBOEKReGS+
QwXwUrFOEBaw+/2jZ2vm74EH00JqbnUc7Zrkx8/pt+WxGkCG289hbg72Ltc23DOr
tKV4M8atZJsUQ0UqH/RLp0doBBaUEN8e1rQEOfq1Qk7/HEPtGSfQzW18Iyw35SOD
Hi1BPwR8ghYdYE6oGFEdoBsJkYp5eYcccZso8g7XkNMLkP5OGhSmCcK5Ws2XIRp5
Bue30f69wWwWq+qTQfjzFSymai2B5yF8vkuKAQv+Mhe/I0sL/Kw6042cox5sZuvn
Kj9DYkUuHcfhR8wFRpdnS80QNZcdQTrh/WHuJHljoueMQtD5i2psD5YZ2AW8lEsy
PAqtUkR96JWsSoWkjQn5wu57EFxBj+Zc9thbvj/tTx1bb34esnn2yE7q6k8QPw84
zv4F2Pj8OuRYnhk3Z09P760eefADlUMVIGJvMHB5fTNJ0x2aHP0Go5vl+T7R3lK0
uWhjVmZEW6/8AmJr4Q1l1WirCopS22OdJwescbsGnhmrzXzBrGbJ8WFn3g7HD5PV
ItpQK0aKjQpXqBEh+BwW3g==
`protect END_PROTECTED
