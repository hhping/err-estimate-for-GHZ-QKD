`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkKHl9w7w1fzxS/0HMC622jTFk1tGUxpqBwAZZJb4SX/J4hz/SicUoX2YVzqK7DX
nJGDLNkpigVw/oxBbof6na3GD11/oIb7qftBB3nVAZuqJJsQ1eG3fK+oA6YS68oV
2kkVrxhimmJUlx6V7wwIpOE787Vwz3/bZSERK8IB8HmzcJXpZ0QIXRfi0M+L6SkV
u93XU5UKnuWMshH8Ahnej9G/xVlJHUCYQFsAUZAynlkUZC1GVj58T7fF4le1o724
YgNysHK3wEwN6n3/jwwiNqkM4Pmp1f9CtrXN1pM74xAx6qSQJndnUbgUfmF9hr2v
PJiIt4EWSZ/706EUFiDRIUXJzOOXx54Tf4oSQHcnHgdIM7NAC9YF1OeShM7U44JO
w7yK0oC3Ps9aCJ0HqdUq3qpsdSikBlRxkI1R3H9O9LAoW9urPK31mM1WNDhHrfE6
QN8rKOVoXzDsIL5EYe8uAes1FdRPKvuLNQgg4t3odcTZCXW+M+DCRQlafrIKAREk
NO2jISY4u1tYA2jsjidxgvKi8s2w9HLHIZUGzReme858bnRUMrRInKRX6xh7ngIB
KGqZEWkYwgFJKoiuOLnCsoRI7Ao6N5fjJ2wK/WUrnhlwdr0yFOY9OsbUqfVcgD9V
h2ViY3wpLvGODOV5Nbc5Cb1hW9Fz6v6mjaRXjVgQ6Ri1T6z8vQqK0frIzuyL1Xxp
0sfM7rRZVd8uiAcryMJNnVMG73jH3Ylo8e3U+vrDc90=
`protect END_PROTECTED
