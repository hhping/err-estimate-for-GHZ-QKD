`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uFWeibdYgZ4su8lRnvGRnxRyT8HxUyjz9qHOX//LUOu3ikgULn/i5o8GKRedXuQ
bPC2seh3Fo7T+xBpePj8szOSDvLqG/aIYL6r2JZ/fQOYLGTpUY5QgcmQXt+nKkIL
sUdR44mzymRUX6UiJUG12MRNINpIuvSU2ChZxdP58AoNgV2OqQZLlbGyXQdC8/Tx
veeTkn9RtM7JLSHTjIq3iXEdi/4YeC4UlfBLoSxkzwYDptHDfk0+v3368mImk54e
imAihPPrXJbmJBvchCGWQNDPBPQWU4MO9GAmu0QUUEd2qRrr1qImXVN9c7AxkXQE
I5ZIv/yRjGtJBVgYzQNSkfIN+Jz5+xwZkBSgNaCqvjR4KLn4VpfhPcQZQr63ZylJ
Rw7GFB7/JMUnbYVgNMMGyl+a8TnXm5mACfOg5nOtAfUF5IKP66gY+gxf8TsF3HBf
kNxGWHU1XBnp67LoZLnn/d3m0VaBXWDLmNl0kPPWnNXZBq7obBR59NgVFiVAZAdX
Erm2fWXVIwpLW/JGIProlGcB7sIBSdp1Otemos9onglflRIl7BKmUVEK2e+PXYMY
92ezCAlj+U/XIa2AnZDLx0VySRRN9c83y7a7d5Yv0ZVXh/PIAOxfGx9VzP73vAzG
mmcVLNqujDDX3ld3xgkL3C864mycx/y5A6lGokmPO6YqTCm2ULhdnH5UI7OruAT7
f2bIxGTCclTmrL7E7Jb325RiR62mhg0VIAyR7KQebCsDWQuhO6tj9LlmQRd87BH0
rvZTa/XL3gCAE+ACOl9an3AjC9yiL0TDx2uU89LNAq6UZrJHMMy1LAIAyLA/RV71
fFbPBLOhKoJJm11ePFEavm8BKHnkj3vLysw5vkyYgPhPtpPFynTcwcxi7sjCTFgW
yxwOq9fjIeQ4IX4hVZ8xGg==
`protect END_PROTECTED
