`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jm5cm6IXVM423a7tKVfv0BJJuPsIH15xmtSpk4arY9M+xkg+ztvFhTacVKpRXZ9X
zc3YpDGbrGCOy1LcpQtu06P6rmeUMhLqn+8Y5lNnL+xuMoQHKqc7Tw+4FGqDcXeW
NDfR6v7FZn0H6ZX0o85D2HSBSseDwXl80IfsnqJAEaoG8SWbJPEQTUmMYJ25icxm
C5VCAK1V5Ht4U5S3/OLKgWWWSRa/MFoFdWDVXfn1x0odRgn0Ug28RvcrUCNe7Rvi
6kdIsHo+C6zoBccohwHoNCO2Uvy37fXnrNzwtpOfSZDdobOx5evS5W2KMCCFdKrc
Xm98uhcMzn0yrtpnTkFiDaVDYyxJCZg9wgw8fj5FUf7XtjiWRM8cfhGfq/JhteM2
tI4Okazm7LkwFbPTuJXnAfjWccWAFCNCCnAZ9nTVJIHQbNQbCErd4enAynAljgk3
lRxDIDyvj6OMQrSLvsydZCKh0F6StI0vlPDzOpCrikPNzJPGZqC83YC6YGc6U5Ry
65MiU2NbOaRTX8o8Wib6CpMagYuz3I8RVzPIIwL/2w9BSdXsmtbZuubowClWyKlM
2cQLCrdPdFVdXfcm3CQB1gDBetQMXpqL7d0fIacHBSFK1OAkP7aYj/eZov9jsuDK
jf9UWprRj7CDY4QK+rsy9y154dm1TC5FvgSLNRJv2BonqjgxpnxKNaPXFAXOpJ+o
G2pHuTmGXvXNBSbhsP/z1eYVq2l8ISFmkQBvq8kl9oKREWFuv9Vp8NtQG9MA9KQv
dL2fLZhACGA914Mh6zfuwlAAtMxgjBXUcFWb9eWB7LI88PUGLGj62uOxmLKy3dzR
67Tq8+9R8TsYsnIIkT5xG6Rz4troXdg0wUv8ztFEUEwrRCacFdIwZSIZ/J3DETy+
PpIBBQueJfjWQ303wypqtnnYTfwoKLca3+KJbnIjFBRHP5Iydi37+mYBL2vBV8Ke
8dkPCV144GDXIKgW/aL0KC27YudfEvAnAE09WpDUFzaedC2UZNy74gwQ/egXXozu
W3oxw1N27Eq4LOG6zsXT1bptQq+pO88NRmxH9kcX2YoPu7ACgdV/gt99ADstw0Xf
E7b9/u1IM/ysFrkj8usVOY0razCC10vCpfg85VLfmBuScz1cFkQvqU99d5RSya6t
Fk05Jr8U74T+r/7ROcoroAHeApMo4DE7aLBb+UkFv6nFZyc3lGt53M+eEMt2bK/L
0nlCkgkRlv3YEjekKEhyQ+/NbC6dWocLgx09vnXxIh9ZJidegRKrsRFtYYNrD1TQ
NJaQwxp+qbqyyfTg4srziXVVD7NxY5rEp6tJ/RhG5kRW16PG0iEj4kUuggPc1ojm
P3Fb4qRN2agcJMM6O38VmNVYTPbGn4U5V2U3BtGgOCDpU0D5lbTXcFvEessMKcU6
nqIzHsyIchEX3aq/WpdFln2IS9tzRAcVjpVRXiYzeINbCGfRnX9URWswPbNI+3Nz
dV9N5E1eTbyYY5+13XPgh9RKwhpVyyOYg7pKsz+kCqcMRngMmbyAdUw8lsdr0HXL
oFQPpL+pKslhmJNe7tJhRw==
`protect END_PROTECTED
