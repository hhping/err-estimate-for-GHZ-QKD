`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xFPe+t8ygM0Nlnmcv8hSxj+wAPMfEfmUl55jjnt/ix8mvXuvI1f/MHlHyJW5iLhj
aqQKToGsInmauhZK8I6H6s9tCHg0bWhmbukb7Pqr3NGySgvWKXeFaxTt393KirM3
JRe9qdKRfJn24A5HdIPt2whbHERNxsFG9dceJgP5B/88fnHxGuSTIsFo3I6k12jo
LGNnXSXVXjtJSTCwc7IzoB6WE/ffOpIun1CSbYlrkoBsr1bCXwIQdDMyaF87KNql
bXi3UtgRp6yyLMVWG1xveMXUsJVrtneAMbPsXV0tYd5H7+kfYqdSZ1DuON7x6UAH
96qrzByNWb2/vRpYJLRxhgh8u5HNAsq7dJdbCsqDrvoyDBR8rLIlHgbyKMbCwSYy
vdj3SdwaYXWilQnDDGWLT1rRvuJ659e3B0f6GUDEMO3WusTgIji/n4F5OR4KQRFM
AXwZc3GhXUofcAEumx4elBJGJk6nRszf9epw7Mp3a8IPCyoh/FziXyN4biXYPsHp
sDkxyBAb0ztmCLPTZnuMnxyhTAx2EaZxHxo/Am8k2EX/fSpTPS3IQbCJc2wUgcvY
OCm/2d/pyFZx9EfEChMLiJstWoxRJ5JKk9xI4jlEFcqCe+Bb4Q6v0E6BJRZr7n+I
g9vQ6sorw8LCwT8UvPHuU9gtUiXISF+ZcgJVDlwN81w+F0IC7X0wvUB0GFmnCoN1
5VTJaAu1wgAx+SnYv/a8DoEAdo8AhiHyxtV3zpBq18eHsOkf8HEBOgPk0AvHW2jW
`protect END_PROTECTED
