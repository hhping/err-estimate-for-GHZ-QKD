`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lRWtV3CszB7e0/LwCMnfnsLC9frbb5c5a3OduKKbK+CDiUYJPrvC5LmamL5Pcqe
OezMLkqUFAVAybJkYiUzy5kGey1ag7R4A5DW6dqaTbjRh904ye1u02j16WNYSzQH
z5dyciuV1iLt78MZRMvGnminNUx7NH4K5hlTXQIHlLSE4HO9HxDjAtLKwLVy5Piw
On9WLYSkWROE8l9by+eC8aV6EXlU2aL3BrJGwmsAsF/EEzL4GAHABfp/cS9dSRRQ
AgNcRIVevR933ZqkMHJQ0q9FGby3F74QFSI2KHXKgTkLIlC+H9F80TZoom947Bz6
CJ4AZvWwIXzk0ZTzIBSBUCjnzMw85wZ0T+ACfSz+cywdCC7EraLca2QS6hkZYwam
i3Dd6Q+f5xdKLwvxYIssqxq1FdDLl7nb5nW3r4coU9iImewVxK6m+eCVhUzoL33B
mWOu6nSfPtLTLUx0Xf4g64N8DxZdVGSd6iwD6jdsDwy3dF7HKQuKh7sc3JkgsqTi
LgtTL3IApYog/0R8asEarFr1cYBxn8z7bmHloUCUAzsAKRRsUFxOr1hOolYLpg7K
OQSZ65Ff66QMqcko+WJ873BzbMYEo0bMs5eb9X+s4rfBbzfDAH8+ELoPUJ37edVm
64qfJKxfmOQbnPiAwr11fQDhclYoWgJTNRnqDQb0G+edddEOhE/L2NE7PXD0eDhX
P1o+BHcV4kEyohMVxjDm0N+0Za8/ke6MPY+2R0VNw9ricXz3MD6nu5V5tgww934s
tzsTOpXNkHcaAcXrYuO6LrtBRgH/WXDyhRuC7SDDrr4=
`protect END_PROTECTED
