`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18J+UWXBryKVmZfk9XTZXQ3UbHuZGGPNlSmIq7DAe3waycWK+rfZyREshV2LYYjF
CTDV1nGx9MRDl1qXIDddeQcdurfjFzhkF+6H0I1ELaytyzTg3/OtzO2Y2gUtw/bB
QI4NYddrW1yGDoKdSPYKvi0lIfrNJhKmTAwoaI/e7CZgFw/cEQ/L1uYOgqCBcaHO
HU75KN4UdVi86i+lk5JxQLzvlhxFtVYeCFJ2DGJgtA9NseV8tN4aJlm6H+CZAzWS
PtTU9Ay1nTImFe3hZtyJyWYJ/CeL6uDh1g06S5X5w7rJaFe+Scl/bq27rifu0dVa
2FRt5t1epTB/2XHsyHvAhLQxqQKC5p5+ZzQSdub2dolT1/z35LxX4bcIyl5sQjqd
hWUK47xqF7K30T+i67eAC4VKL+pW2HPXdGSVUpcggT9q9Xy9QHC73XfHB5YeLyb6
t7IwW8LwndpcZr9GtHsI5hWy8MvCiaPLeLaykxkuCOfHlOoT93lHMZc6FE8OED/n
NwMjzCAR0Q4h0EzK9WEuwCFiFSaIQ/ZD4lNiJLQn98ggmEfTJXv1j6MxB/TuY/eG
`protect END_PROTECTED
