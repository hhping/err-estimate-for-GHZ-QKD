`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+CQW9dcNaEguG6NgfEvujZ9EYCV0RtgnLywayE3tLRcpA+nO5moyW3dUbI7aX2I
6Uteo2PIOrY9D4hrgmTncxMuJrstl4vLQgnAu8ThlXhE1beE5JXWu0JdZw5NlhPj
oCvn2pOXaohoEm6PNcKmmCj1+DMt7E598w0kvn8Z9dwoeHWOW7UeH3KBftFNCKC3
gUwmKQVPfWILvVO7QSN5IHy4zcW3a2UMJRJH+vM3q8YCDzy+DdZ20B9WfPvnEoQm
EUlaHzzPk2YOYwvnQqHqgSVEhx0zarC2zLJgw1kij2mqa5tamRAK9GKk6+tuuybM
95QHDka3ns4vp8K4Lq5A+U3AWr3EHFSHfGHPxjnlI+pzjhyFlV7G2ceuXjEOaRMJ
BQuirQ6dAFPSME7kAZ9vUyIQrCx8ekTmRS9FliwZREOnQc3pfC2AV9VLR5xk0G4G
d0ndXAVixbOgjrdSwui8kQ+2Xy4EuopYjojgLAPGrocKWGO7Q4H3vnOclG67CIxf
wKpFdCeVXvQSYfFALKFDoBH389HXxfeQs1SDmDqX9c5XLsrQVsuzja6cmowPriww
J8r/XYIrG6k/WFSOV40t4co8f81jio89AoV2kJPFbDDtnoe5N3GfqbbP4BpTKLi+
Ds9aJPaWve0dDlfyDg3Ux7wgScbGEfDEOQxNpM43+Ws1mA702dH2KUSJs99fmoVN
890c35PJQ8NqAp2rKh+G5i101OGV2tk26rZCUmkmwZPigaIrbDKTdufWGliQzM3v
y+6A6DtRRpmykcSGTese5lqArR1N1gG6bzQUK3Yh5YH+tSSrCmOJuVVTrnX12+ok
A1b/LZ3Uw718I9ndD82qz+I1m213BlhaO5hPql1SoUvqqGKv+/V8v0UMP7b+Qfkl
MAnts5uc3/oeyqPigx3ItDoXJ3qXNcoHEap9a2s0TwwhSF8QFc+AyAIu70xnDEAQ
nbjqqHrmxJx3/VJffrsTNHNr+VpWBOQnzvSIUt5xN3Ex2jIx6IIRdfxCCZsGIBM+
irPxNnhFX1cF+ICpL2i632Rjf5k/+UGBwMm7MXIstQQ/nza9zhFavvltJXOqPuBk
lp/occ7PiyXarnWPxM29yDdPsfK2ktlfiy0ZNIIyfdv1LrBNtdYYMMgGNe0A+yDp
bu78UPNFkmJFXBtVe0GH6z2SqNOMMuFVoXhbajvmI29AtNjBaIy1WQLkHoyrVPq9
sKY8SeMoNJjwWYMEgNPv0GWA4byJp7uV5DWXhIl57PjJ7x2WnMP3P5PZ1TlbRRx7
9PdpQi9gGmjJ0WY1BAOh+/ma2UX8+wfoUGwuQ7vNtKYeqsG2z/a6i9XAwIzyZrru
IEamip8PKf/6P+G2c+CKBIv+LHjSXd7pmm7mzEpyoRKC0h8d8p1/u+fxl8dY5Rg+
vg6Ru0R3DieSoifJnz/IqqK6wGdnhEsA7tkUWiU47d3rdcKgRKYjngQoiCXP9n8h
xfDI4i+1HXvyd0aaIA3MVqRdfkcVhF2+L1oJevlBLdct8hLheCPpw3afkW/XSY1K
mWPfmnqy5UkTjtSy7FHj7wC0kAKwW9igl7xY1gawPdCrGW5lT/mxCtvsqx/TOK2U
HtiVFXpsNbhKAXQDlEjVbsADagtahqW6zxndknZuYFK/LJQVCmk8KEsLOLNHPTEz
PA9cKsLlVmafiuLUGRov/qF1JxTGHreYDKpJVq1H6oaGhr4QrgOBvQOV6w/rSnal
HbPhfcrm3P67D8gqqYfxDYCGKzSBbCfMnW6Xop1RaGkvbQ0cRX6kVKqpaU65R7n4
CGmwBQPuEg6Hh9H/KfLW1hhFYFW3b0bQh9g6/ROBKUeThZM30MHKyZnltDa2/xuN
HOO2j6tlLML0V6NQHukFoyDjMTc0htN8jQQDFO8snq+Bn4VKj6Yac0EC8gRS3mu1
vUau9gMnsulG6dTmpUnxdbW7lsUbPOZYMfPeP4sBZYaTFu9mbAehXfwWmRDHxYwR
zsBsXKSkMc/2YUPElAXc8wNc9LheUGeSfCBT5p1KwV9H4wbaagImanO/xL0ukg/8
XOezvqKFy47px6fFdp2iAgeue5Dn7pRzEIQU2HqHy+1uf4a5IQn58wthytDyRzxh
2MraEqUwwfn0RvHhD82kHFxGh+uNpnFL+Al5xyQEY02aVx+i6Jc/LLkQQqcxPsV+
StYXBZI6wm1pCuPe9RziIijDSF1OzkzzqYkHKYH8A73ZK+GGFz1pIDVwohTOClbC
2XOFRP3r8aPJ845PB4zh3roM6NobijagGmoVFMy4NhMjlkZKTvYgsWA3pOoxJgaw
lL79qEdt2dYgq6+xVGYu+XeWpUrkn4gjftELF5oJgAt0KMtLt/tz6idxrT/KZZ65
C8GiJY4Au83RwB5Sx4Tt+8Q3Po/pAZsg4P4VBEOjZDDulTz+gPaunBawwvxWvlQ+
IYho/C9ljG9bLJXEgUYTuFCPnKlhNZ0DZyBLuFrApaQz972EV0lRhNV9XXn1hsDV
oQxX5pUb0tLIsPUBwEAXYC7id9ve4Bmn7QdC9Vhllsq6kkCD2p8AMdrlMEpzs1qq
jEKEW5yh7vEZwVJnjfHMa50MXSRdteYZGG7kVYxuZ76SwDp8q3Ngz00zyHfA4gn1
93oVqrZQiRq+l6IjIPi4+9Gi8uiKwH6IBKbEvIRMf62W0H69d2ljKzppNhabI+zP
zRJkcK6uwrmVfGdGmcTcImNKPEsP2NujUvECoGe2sLQcrtHPMbYaTUKDon3CmTkJ
WcorMbXx0mSVFrv1+GFEESgeuZ+ElfcxCDFZ1sL+dmkHSMATYsZQBgyAfLTpzVyf
jrLWH70Foap1F7EdFXey4R8lwwYwMUfdXJl2jweeOOwtmOV9QmkPmhkKPO4AMYR6
EGy+nw8btIBVIubzRYVbC6JZI1f9cQvJfylLs6ibCWZezV6Ja/i/1XFseeA3KQzH
d+iJEFf1U1BrnVFiDtbN/5Bot42ACX9wdyV2cuxNPkZlQLwFq6ICjO3Pigj1oXOH
kXPdIzsTtu9vrYKqgku1UnwuGSVzo/FfaZ4xAJ1wOEzbWUetOZEv24fhcDQ5EBVR
yAQ4TspRnSjslcksl4Dq4q8bFWVTDZubbSfrP+lLhfjBe0ng99rSeesARl8l7fuI
OxK/sJC5BBPN+ajs+YEyijzpuNWplrR1LAjpcC3Q0HsZfMP7OPpd4KqpOLvNCTog
`protect END_PROTECTED
