`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZTJhiV4nnAvGOU4/9sOR0Jr4m6RuAdnSjoD1Q4JJQ9bCoNvivxVP4mlz9CuAcnq
0OouK+25VX/Hebn2dwJmfaGY1/o9AypbEJs0FQdg19dfKILabyofRCDksCuiXmM/
1bQnvQFGmAIJoUFvMcliD9SYhwMb/z8SjDwqdausblR9XgPNL5xCtgOYbhDgp8SX
dfQfLw9vFxvyyrzYCVzEb4zli1deApP3s1XLWs9vhFsb7FdL7CDRmvpvZK2rJ1Fh
MVrBbjo0zkg0AaMgMBsYe1GraHluHttIKDT16WWzTuBFrlmaq0qLF6IN3yME+HnW
u1UljixrT3thwRfXSvdBRc1zhhHtKLBxi/aIXGAsgyV0v443aV4iblqZuGd4DfAy
cLq26fT+VBNrrdzTXKiLE8Rr45fLZYdgqemZTz9Cph5kezTvf33CzqFSOaZztbwV
xNycA3b3pRZBgxQ2LL7HXtOQYGaawKJuEkU+sFyc/FfN3BmYSXcD/T3r3GO7tQbK
1UNDZoEDjCo/W7fuv57ncA==
`protect END_PROTECTED
