`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IV5uxMQzaoaiTOJJxDJK94w2ppKFBovFObMpd9Jn5GQ/H4BQqBSr9aTo/zK7vfR8
NkhnoI78xP8jqaQ4Bkkaa8wlQeCnW7NKyJLpE3RPCVG5+UXl76MDalSvzNFyDKIU
JbxsegygvUAhoRCewl2utbokIEzN2Cs6sCMIdIkBapdwP+lbWQcljbNh+e72XXfN
x2/Y+v7wqJMnM7UP0WLXPBbwvk5GCwOxxNfE7nGCC2okyZM9WJ1eY8Yzll5Fx72Z
X6Fo4/m9LH6pxIOZaGQjXQtbswzeOMMe9s/09xUn5ov5pzbxdqcajAZOlSxCbGoO
7PIb7Ce3SpNFEmc12LpFI85mUIHq3xaW2EjvhWn6xW4+Asm3oM4kMLm/6J1uyAqA
eFmLco7AExrrB1hwCmFAtOUgq4p0GVYDhuhvgZARREDJLbT722rT8MS2NzBD/1W8
CWJjhaaWUB+AL7pyswv/fdCngPTYfafLb459kgEc/+p3M8sI0ginxBa6pLJufr1V
Na+EwVPnbC/ek6rNZBYoIiB4CWi2DBzRaO9pMEOaJr51KkGB5kZR+wurksaaOf82
MPY38GnG/fyEU6iC0VL9I7LTM3BCnxGuMMqLWwvm5hEXVO/5t3bTvO53P5Ez+SEV
PVZuN1LprIAVeHO4E+gIfsA/CjAb5/ep68yOQgmulzgWDLGk8Po6YY+C3N8e7M7t
nj+d49Qn9Lo/qfsy8lNFluok2XFkbxe9VjOVV4Jgx41bHwfdeVy493C3CjjTgPjs
nnwvmVqjl0n4RWO1q6MQ4XXzrSbSQq1f6BK+oSfU79Ie0KO9MxJV8gVBUdWsKQUn
QhtbS5BweB2gfLQXnsIQ5emELGDGNCZOzkO6DlgnlBdZwGGOOILlEZax+F0UVzhb
+ZoLdZV3F3frsgsLr21h7TlOL46PnEQsDaGxfnRAsHdCh/lp1Ibc/3M4sJpG8U3j
ioo88PTVYkPDU1SiJSxbdKA1N1H/ColrmjaFeFkdLTTpw8BcWI56xuAQwCUNIGGU
lWyKhDixFJdn24QFyL/MPyMvTtZcjjww+4x0A1ROEalur1hcVy0bhF63SA1HsnjJ
o+Z4Ogyz06TO7m/sUMA30x9qLirmYDURqSDXxdW7XrA/s+xzgAd5zT7RBaR+Qque
G4S4BIpGGRaWRXXp5Pc0D3IKYBFWToUKzyRktbNet47e4wocQ9BXVA4Hsk9Whuss
1Y7emrnncU8kcHzkZG31MN0HQyW3Rw1Bs2iS+RdfTaCgPSxy+60sDqJgIHoHPGC5
SSj2gTpI/kr2JySEgmlpgAk1sRKUwk+TSNnC5Oun/ixlZBO+sVrFDUapFpBzhY+p
GxD7uvSRqliFOMj2bXo5QN90zuYqj17MdLMIbsfnuy8oSop3Dir68vQC7ZcCzve1
2PM5jUIwntL25ehjHVT3etyaVfoKhuLFR3+UOJLpwS543INin8deC+TCPiLU/0S+
13CNorrug32s6H8bl6+1nLfEmmrtpbr5myD501znYjhf1G+LYC6S2xyVrTMZixjr
bHpsA2PlDPDC9X4mXtmIFp3lrxTYOQvO/qB8eOfrQf42fNJnTSSoRjem4L0+mx9x
fqrdsVYrfg0fUHtOqnLrTmHciehGoctTrgwWK+9s/WhO/3rIUjkH47BHG0X0ZP5g
+ol98ANaFBFf7hilUwS3GKtcQ0mKTxmfIVGKAx5mfF/wfTDZUwE7f8Hn2EbW7++p
6FooWejJj6qNpila6EJduRgkRskFwxxb50vSh3KEBvJhIag4526H++DToN15hzjO
iuraq4R17JzRowkBO7XBwcis/POBpWAK7nyP7YlDhjB48tbbgYUXSudbJhPXBw/H
gsjtihiUZgLea6IL3KnJDJJSysw22ZEUlOuvORjMaoNx2xsFxijDl53keC5a6J6W
gsSBk83bKaTpQB5L2vYfVnwhxcyJqmhMwO2w+vOrd9W9jLFhSSimqpfqD42Y/qVJ
6YVj0DquvvCBv8YXVQPqYxO7xbqzynDUK0Be9h6169D7CMGRjZRiLpVGyEu8Rcnx
jvaoSH4kPVK/Yt97Cn07cFX1FIFKFWP186jsUUJTaoTPnUZADVtCaKgRxM32bTmS
TmDEOfinV7NgjKulerpwPeROdOFLT6+7S2DrGMo9o4cedXOKtN0kk8bVMZx+edva
Ti5LyUDrWNRqLvBG7SGC4yN5KDUGqTVH3V3j6ggrLiLTVfKXEXWqQXY6QMx7YQhr
Rn+dKRHY4NltOZ1nSdYC87Q+Bvw00sbD9NSWXJg31gwrfkvLwc4EB6qNl3LruENg
ijQ79saOrdDzySt1rGpwViOHiMGvLvaaEDzv5fldbKfEEvnRq4U4k8O0B/ZEELxX
rIKhWv080SbfvTs9cQJGfotjDJbwrhBvJNNxvSKkJQOgczhgmBtIegyDDTu3aEZK
BeCP/lkF3fddGsOSYSaYqGr9d69TsxSdGTzqi8fMW+ptQblGacAxWX/MfeMt2F6K
Skrw/R1QfOssjZkHV5bMg4PUwTX9ftSud4/AfX4+57/AqmPYrL/hwfolLAoGN3wj
NWshwDq/FoUj9EC6ML3DsTvKWK+j/G2FyAkBtPzBAoWO+ughs9kmbMhxiYFACBRN
+FfxLTMEaPuoU5b1enl2FBizCPOxD3xzDyPwo8uJsZSHjq80QTXQmAunP8AjLANm
v47RdK7ff9jrJHpX/wdJk31egLz78Qv/Dj3A18C7lSX573rtMcRSgrWHVU08J5zW
vETwXfxcnXxrkeCBefb/oL4ehPCYvTzGhXQ3q4S+4fqkCZyvb7JV5F8QTaiRLG8u
eu0ozcz2O8NlT2eEvLlkARc695HzkpvQvpPkNVH87g89zHEFYlX16Nd0VBP3P+Qb
L8XEoZp4B3iTlUFvueauGMtJuDW47Zs0jqR7plkyb+LwO/N7j0Ky9bMBromsLeqW
ebYRXfXdBh0ftaA+oWIAefGqch3FbaC7Ho53dm8gBbHRoz/rnhxKioopfW6IdgY3
F3F/d7mAJfp073IQSi4aAZ+4IH31NbzToCqvOeV90y7DUkGUL1kYZmfsEPTHBd1M
y5Jncdwo23dKo6/MzlexLH7ONTbxwg6yggfSGLW0BsOszMJ4h4MZ9q1SjufHOZBM
5W6egl6Hj7kdVm49MJ4ebUF396KBE+thh49vtYGa4Om0JQzRhrr/mBnczQ8qfZmm
AstYiIkxFF0lXYHPKKtrjU7U1upPn/AO5wLhMyBrJdGP/2pamimbh+egVi+1+AtX
vnN/0Jl0Xtj8aj+IevboYsy6CMu73NHJTuUemGR61gIgWYg09QAU7697SAARNw7f
/avfO+CoYxH39EM9PzNjFV1fJ7GTyaYTJFBAVm9u1fPDWYmAXDULOi74bNMugEXX
hdh+YZma2p8D4ifZ+eMs41ByYsgZm2Szq+sa91oYX6CglBYaPCGxRPK0y6RsZQbY
fsXazvUkpXwVOa0QloW1W+Aj+ebsuhMP4hwpSIc45TXfCSkjTyllRu42Lv+V92Sd
s68MjmNs9dobXM7NfCMwtv3xZiz8wqjSC9QSI1yWza/S2mLaWyajDqC5coBBG0xR
Ja+0T7j+IXnTDAm7FOzRLGdYXPShLS5gTzPM9dgCdlbJOVpkjuMZC9aSvYa65Lh4
AMc5k3lKwaOVRI6qg6X6Hj1dFK9V6Dj6L4Loy+Vt90Qx8KzVDh78qc/czvphso95
ZSfZONA48Yzz+/zCHRKbz9Izuh89dRj0nzaaRXec4lwxaBcDP8q0LWQ8aJJa2l3v
PGW6m8my/gw48r2SG0vhOb4EhxY7eNYAQkwgHYB8xVtut1EEoAF/zPEsW8NsGoqs
4Rc2hXl5/pYKEAlJw0wK9zCs60X+tWgF2U92EMbfI/QhuZ7ySe0o0Ee8PL6B0Wjw
nsDRsdqDH3pUWiXuDZdaOTFv8sS1vSlaUVd8Z+eZN1bNzKoythj+AWUAPVpnzw+7
pCqkG/VSvIElm91sk15RLJElc6e9KesTKqjIRW65WT4ZcpSBLD+Shds1bhLU1Tky
Ip8FFcq2Ha15l+ICLf9PcNNhvchODoQk91AAqethsg0jrTCFgXyNZoGkRuAXEC9H
PkqUBttYbF23seofN1/9b2kF3aOF2RhnkzbE52IiXdQ/V4nd5otfaDTjFm/L9QKw
AhGcfrkT+Ve/sKLpLKnAqHh/910DLnaJ2ADQijCdRqKUMfaST1xBGc/hmNObFwPY
mWRV1MJ2iBYUKSyTI29KurpYoouUZkkxXkBrBxJLcO7hzW8GlltXzEs7iyUJzylK
An8Hqjc+djp/mMKX0iPnZTV1Kz36FPUZtlIfPnJoRYfbQKc0LFLtaUHISDIdk1Xx
wcBtcYxqMrWV/4AIpF7yBHDJWFqRAfE2peAuyv7hNfNV3PAcGshsym2/HXEqYF7u
5miaaN3WKF/UHytTFGEfvxS31867gyK81BN8jj7Uq4//nE1wRG8ZyNevCjEsCebi
Pzk7X4wR0DvkCl1gM/OKBPypx8GdbOyLW3g91cZG/LXExexY5xADJ4faDFG5KxNW
Dympli1iteDyUKEBHiuqc6TOpvXJPKxa+hgUASwmu63TugSPk7O/nH9gnFWt3mvK
wSPuhk4kCmCsZ6B/rwwS+HA0UN1wVGJ1gcHjZAfdQ4WLp2cx1HEIRdIrQW8h0G0V
Ljig9vRIBeR5hKpsqYpe2v1Ff1ksNxhEr1Qbeyk7kCcR3Jtjn1cAbrYRjnIy3BaH
Gx2HOrXTqwNp0wKDdM4M2J0Gi49ZZm252W1vVIub6MK41nXSl0gu82sw7+eMHaUg
NA7jUcbp0ezqwq7ymvYxqCN3Zt9xIvecT5D/PViHUFWYoplKO3J/OvOHLBvRbL/a
V7JJ9om+Rk4wH/Z6JL2eClEcc20BL0Lpa4udAynlwBVGmC7BWpgS0mzigGK2EwN5
A7NuRvWuElWyEsYa57duE4bHSS53jnbfvcFpzVFcN99TTf3eTsJIzPDf0hkSWOaq
ozTBcvLCHBsNiig3p4id+IZVrRFe1aVrOMvmEDprelBCejf2qA+HlTli1OjYV5JL
abkpuqc5wOeFsm3qv18wfuNvfekpaspCBqOSG0mJ1IlrBCdXURj662GQ7NyAbBCv
sUheYC/qq1oQYpOfmcnmISjXV098/Y4F2SMmcEsiCFG+WUrEk0KEluookMCCUZCB
PM+HFdvyH5ujfzqVPsEyDLAZ//XT5c8SctCZLX+NCHraG8bHSdBTWh5oK86ux602
xvJFil09lK2z2lJKZ3xYu7b/xChPeCem2/SOgNg0MYMmKXb5LCUkj5y/ZJaBPx5s
nY/CQeZGMDstOghng+MgYuba9ukrs8//do8qLjgSTXYEnjp+tAlgD/hO5JSy61t0
F7q34Qu5AhWY450Nwm5d1bd36ghrU1GAWyr4OpvsHLAFpE7Pe2+Gw/J7waTRjIBj
f/2v4XJxThnzRJ+AvVMqXbgMp0B6+6GK+9vkaKdbc8j01RLxddTetfhwksM6hv8j
TZCaHEBYbiBVp2KJ/WKEFNe5A0+7ONuv3LwPrsqOlV1bI+CFK8+TY9yLYfBEWDNC
E8MqD4aLMozGijN23qfeXQWnJezB1LrKQ87+o2WzkUqBOAnU7QBCI+uq0NgMurcp
flYX5RKn+3IpEtQ3MiVGvUV9BXs7kJuyAQ0+YHfkfod0Jm6LEnsy5nxxkmVofKc+
3YRWFIr4a2NqwA2yfadn9iIhlp7qLKdQG6SAWRzDbG2r9K632cKaeTJ66ZlsBZ+e
1gtbY1VFsIkoY+ixjVwLbLFj6v4v3XKc0iYtaAqSBsUQvK82IA+lwyACl6BxvKmA
cH2ReU9PwYA6uxfZFoGaqVmbpo9a3YaN/z7+7bSKn77ue61cHf+52FPbZAibu0qh
x4rnZgyLlULflp6eagkrjtqDTTjR9n2uyWwlh6J/ka0Hvysw4x3M6F0UiMrtwO/o
9sogEaAOpl6YD6K4k0KQWNmTlo2MyXN+MyR+fpM9tinGmNJ7AXzVXuM7gTpEB5UJ
r99e37SBALa5nxVEr1DpoLLMpkhIlxzv+ja2FF3NXtV3Bz9sIX7SgZhobShdLmDx
FXNuwwMf54F/1UJIrMTBJR/CDPFDx6GE2kVvnFzM63B6AgUuzvNhDsls3y33+zow
Baxy1gN58EhOse9P1/CO/cBFnU0Nc3b5OAzegOiLJ+L99lSQkTuBCUWs4kmPhqsR
uvPkJIuKd71+z95nckq50E94Pk8K64wUWKsu9nVGDKC+Ax9mPVXJ6efMR4HDW/f3
6mC2Cdlxw3AGLZh+ngB4oUgyWkz3v1TcIV/XzCUGv3ek251nBWf6xPcI4ShAadn8
n72quAS3Io88waODXwdyPFnL/ZVDLmH9aBIGKYB5Xr9Pean4DgwI7Z1fY5Bo/tdC
3O6L44I/xRbARc+aRZyfoT2DU7AXxjINvNCl73qlD3FMAlnQCAk1vh7TUR2YyAr+
AjLJPdbPxcz2LEZehw+6XIQjhPGzIBbxxOGgwagOsrx8FhtQ9UJMEzZlheUWhjC+
XiTyD1+OFML+/0f77QVJ+16BL2zeBPTg78++OzxQEeNzCO6fj3OU2dxp1pNrl01C
hymSm8cyCgP2uAyDf9x+AgYyb8dhJQnbOQgDHv/aJW+UOjMvWzBz2v/iED91XqjU
yZ90KWaA2RF85NmhE2SuzIJyEIiHS7IkUC1EUOLa9CoAc3XcqApvIioQVOV/LFKV
1Fpi1HGtMIkncV7v3m55DVFW0jFpCYFmMviGNMEhPr6z7Ubo8nbUmziNeRP/kmcf
Zdm9xKvsrYCskW40EN3r2uYYXbCAAQpEqaHIlDoorWRbtDR/+wI95QL/TAc/gehI
2TEJgJvfwhrKNb6kPm6/qQnQ4KtUZu6bSt/BduzegQgbFfPh6ymZh/EHyilGFRTA
IT9cPUaprJl3F9JBD0wUSp8IgvUwNcj3PC9OMMjMWkh7jHy2p07URVDokuPZIEci
faKG8lpLN2hYXchZNlzdZptgTGgO6HD0EUUPFyl6gndHk5k5hmAHr3ZTHd6xbn3+
Sh7VDp66Up6XBmQsLH/nxCUc2HwxkuY3Nbf26G86C+1qX0rWWe18Z5K08Tgvzhk7
MsiYFiqyLpo0v2yS+7ID15Rb8nxA20prmOU/l1+Oiy/VGJ4HgamD7dJYqMditTOV
sohhvyEeR02R7KQfieKtYYahLwOzCs/w7LRvXSlH0YRiLoVJ3r9Z6xfGqsNAu4RC
XidAbit9Gl4WZCnDm3jgs34C9eOaOQf4881zBshKqH4NqODmgIclu4DpANDAa2AS
JmDujjpmZsS77CEIXGJJo8m6Ax3NzLpRrgSgCArLj7Ykwnx3YWZFh1u2Kmr6oP3v
nccdbR5Gm50g/M3ulUNwSjmkC/cJIM0FN79PPCkxh27lYHSnZ8N1TDTEhCCXpHgf
6CkNfTkKZdHnhyFjRLJ9cDN20/75/IBh29C8cBlYDIIpMGKOgRCajLUmdhbAXxb1
aJ0gG9EMr/ruMtXy5sIOAsw9MimE5G9DO6PbxZPu4bSxYbAGGmD4ybR/B3ARSJeG
PNy3Eqaxxs7PbevEBYmu9apq9s0OtGEnXZ10Deykl9jWRUjyMEiZCzhktdD0ZQvr
CzYnOvQqKhJJawGf3CKcgR8pRNXoDYLLUuA2Kw57V5wtliQRC+t/YYcbXsxrWMrn
tb51girTuId6o6nRk9uZ5HdOGghoJvnnYFeVb8eXBdjbaV7NCmkv+/8zUKMZxSps
yBbgq8Fgl/6EAOfkwBoDYatmZfatNuyDsUCxGs8zhQ+D5vkcHC+FnqOj3TMH2ETP
xJLFliH/r1w/Xq3QMOl7CN0gx7MTgaawexudXe4LoOEst83Brxs9EJzIyYg2phA9
2qX/1PamRVZf2NSNsvkt4vHdwepoQHSyarcuFaSflYL2924Vf6zouF0zUsKDaGNW
19czD6VnfDB1tY4J+KK8TWGL4X1z64l3dnsaPKWX/j2Z6E585HdxgVasrUfbTt51
xMEqlVyjKLx3Gp+DhOA3I9wO4MG0LkQn+l2P+NDvi/GzCPQfklDozDHHy2vtt7gg
4caAQ6Ub95ohXxWR8GZ5OwVuJy2a+Hp4I/Cnu2uvYiKIEAIUoVAC1iyNf3V2Pmgh
R55McO0hokhwj0ojRBHHh2fc/L02fK4RPtcB3Do0+ABhBkas2ojtZ+k7/d7qto+/
ev9bGB7sOrUI/Xr7mWyO32A/m0oip09I4JckEwWbSD0/45D2iJM+BHu1QUJwuU7n
3Iz4RzSRz59K4e403X95EAXNpJyAupXze39MNtTf+gyxEVv1HKyvJqWhUa/hXlSJ
P0gkGBv5FFnd2IXOCWcUxyby2tK0viLNo1cMZGIS1IywjhyV9eRIaP1mByXWRKSe
Fy7hsKdKGJZrskcQ8qowVkWmR2PxgsnlMKWnNLkc8SLjyl/zI4l6IS66a5tp5s8C
DnK6tcAejUR2ye6u5okTYAHOmumbRd5+rKh963J1MmPKwECgntvZzbEwzdCC+aoq
32lr45nIJGdNrdmMnoABabZvz661ZcFJoaGRRdixFnibvrKmga8wPp53wp7yNjqx
U9xQcFfbL5ZmXSUDCI24jXdcOoTXC5Qf0iftyYtKtdEqCvzlbLli+6FPOeqJVlL8
W6L7VPD4si4Vn2NTfi79xFROpQ2yl/z0TpKP+S7lD5RyfYNPq9Dl2MaI7avnLZ+q
MmPs2+uSIC220nMd2OqCB3i6mWU/Gg/yQGOjWlA+ttkSog7jDqxEw1CTtpXpzc1y
I0k3NkpcXJ6mF2hmB4JsC6R16+uwFZ2NAL8Z+wr1RvK0J//wFl6Ss6uK5wBtmBlS
7J7gs5QpN3bBgXt7VlZuzj3J+3gN7++H7E5pF+Pp4LKTcphi0fI6P0KSdEcCzqH3
KPCEFTgh3thqMAhvSVyFC852Nj8xnYqQzjesgv+jH6LM0Pt8U2hVD4vbP9DVBOvU
d1CDWyC+Z4SITiyOnkv1VbXT4z4vq8TDk9IeacbbRB0gtge5O/vj7xiKSSdLuifM
uER7ajTquxzN7RUD7XrIeym2wpI8PMTOGbn4qmyDrqIPmQnGVt2JPlmTG8teiQCz
O4ER7u8FIqBoF8G2sZ/c8qAuImuP80CKYV/kdLQ68pPdLGfASdesszdV/uAiBRZi
qjUt2yhzkiwX5HZ0PMw7gfAhmGXT3dJA27eHtczP8Vfy1+IjAzX0datQHU9Xvrzf
ckRsOeqvJ5sSBvNjyl8lHVqZ8yjfG4CWz+fODBUxlXNUWrk7Ybavf93i/5XaTqWY
ih+griiDz6MGRU9FblgBu5eMGPavAva9Edci8cPJpZuNCud6GKsvKyoUJOlcsp5b
iTG1GysgFWJ6C+o51MuuqR3BlfWulL8u45nLSsT1nOMllJi+TLlZKLP9N/FmzXeR
IB7m+lStc73roVP3L63CmItOWP5qwlLRzmkOwx0ujS4mv6MoXiKKnwCMeNrlm0vX
b6VNUJvh7+rY9Xs8Y4HA6uoEFJIhmOSr1UgW5Ycz8PlN5LLFGdTN0EHEj26erVbY
dVMyXhTtrI9pmYe/tttN0P6/0FKBnYn0G6w4rTenkGGfauBOyQ4mbGOwheYibxBI
bG0T8IaoNcjTc7H3rnJGGgcAWIDntrOOswjAvUhzawSY9gQX933YlOVViQyUr75l
bOG+7AfpH1xU3tQc4ysTSXxopLaEDb1rX20TO9TXHEOYOc95fnTrlDNz3JpIn1zJ
f2oBKXcB97yOey+nYluWcMMjYXfZ1vCyL2+tvM8zQDbngIrd0TR0SXqaq3FLihfN
rnCYEO1HWawPb/4cj+hXCpte/8UJOtbmVE6wZHCUtCVeWgEZY/VvLWtQU80lIjV3
hJhKTHkgDi7d4NjKTcbzaOo/lky1PeSeFEgNuFyLGJZnRLCnC0lQzen/RC6r6S3t
RJ86b/JZ3gfXI5+Ksx6QcVyZBVPSg51IN8Bjw4JpLErHHhKQEzDlooqtRAMxzD0n
qK1RhlzYgcxXN6IIdoreJuTM89mFO5TtmW64/Eo4Quqq+izEIe+wiGzCRK05L569
W8QdEndzuQEfeuDEfJvI9gtXwx3PYr2LSKObN81xL388UObGtUyNW3cLeK8ZzdBi
7amMNupAW5CmdbnYIB+W27p8rknGQ61t3wMczg2vDI01cqA36Yfc/zSTOkBNNxWv
KiedjzWb++QZIKMyN+TyvwGzdOb50eysgOaWltP8XBCs4Vuaonv5D3lsesvWglqD
ridrmEyngv+hpVJ2t98BlRvx3fMP7k0SYVUgU7B92iHIweF3t36OH1EbYwxQyTfQ
2MecX1FqSQW/7AB0tcyfx/C3sQjF3DRKJ0xpVT13ih1AgaSMBdi2lY0e5fLU1vJL
6BiaJDQibFNuF9dE1gM5aT8DQIBy/N0Ta4jYhg3xbFwfWlXxuyVDxBaTQBrKUlTl
LZymmHJjIjki3gdvDFu/fzURTSx2yFImbzS3VSysKztQqxoW7GYpR25Y5oy0Qq/i
yGVbGhtVjI8XIQWzSAr9WBkWDSJz9OAS6/GjTFtfifvF0ko97PRu5LCsA2iqNFwL
8uSY1WQmVlcgKxHF70Tzx3FrkHl0IC1Kg4MTkWuAYCJMNPdQxAmcRdMB3mk6ExOi
G+hAGVyLI4fkKGqcQRKK+3N6BRXSoSdGv6rtM9ZlRxtUVkIK68oqBBVYan/o1TK2
tRtdKhYNNOoNF8Uc1AmPPjew5BPMr1z9XrgFxdqiVQCE0OnrYbCqReOElwZH8rSW
92MBSEHP4Qk1YhJXno/ugmnjXmLkxlJB8n1yyoh/p5VnQBZLeJ+IchM0bqSdwfyV
tL9R11+vgvqVRkboAKyENucTBVWCw7wvyrf7FIq9/Cz6r49gqi/f4CLqc40J5UfA
2O4wupstW0zgyo/Zw1E/z2wIhMYbQTH2JuSFpoI3PjqQNkU5y/+YuO1sbF4wc77S
GkwPIG4/6FVOzlemICuv7aKTG6et6EUHaeGz/M+kM0SoqaGI3qihd4+B4l/uAN+O
g47isIgbuPke3J9ZoQHDWz+6jhmjCDcMynvMIMhfg6aHOeeTwt2XUhesZPgdBauv
Ep9TXniETIO0E9PAVq5D59jRw5LHXGEFGHfM6QGnPpHfNAw28vjfjInyIe80Y8dK
nc4qWCEgrfJVPnCGkjWZzh99o3thbmFYWZyIcvl9HTVB4iLN5lfahETzf2rldgW6
EFkFsR2MP9fHPQz/MGXKgDuTfIVafjpP41TTMaLDzVPS0h2FR452TvjQVF0IDwOG
2fWFHPUNO5ZaR0IBTTppojaFYZh7gSibYrlx+w6VklwIZz3ebRcv7Nm2QwKWPoo4
1FcIZfk5sN1j6j9R4DL6TiKZOd0F0DVIFx0qgjVcPDjBJewcepuTB9whWahfr01g
LJTq22IP/ZjsFsG1MBVh8jDhiUY2TkTuJ/nL7abFLrwofXKd9RCJpbOEFpLwq/dJ
IxHly6zZ+tJYzfS2ni2Y+Xd104HE1Lm8EHxqQTGMJh7s2cLTqfGZJJLeNUwCK1m9
jobZwGIgjftKC2IIz9XqfPB3p198B0UVmW+qrg1uXpKzJE6kJiaBWF6NHEDxNMqH
A+Tx1d/Z46Dw0YPe3Kl+MHshKfId21t5Ekb6zIUAttdoRbxTG36dYN4IAUXr+7ZN
zHoQJVS0PnOmaoI3S7qLBduSYvb6ktFe30Tp432mTaWoq3c5c/HxKfwotjGtMJ/t
enrGmryPVxs7cmAJ0U2NBiSVG4vHI2BKUsVE9NN11T+gUkQf2cO5InywEe4A2Sos
RQ7KrxJHTrRLOlo21FQkD2a9sZjrF7uRd6PBFRbTjhU+gT5gTnAsKWgL8Ld+bEFS
UJcpPEbl0vijqGV48ad+Uw7Axy3QCGwpEMuyC7CXmK2Ukl7yO0FWlCgdXON+v9Ec
M2iH4l5kHGRqePbxVEAqitv+lfGZy/+B4ALwJP3ZCks3q0vo317xg0yrc7jzqz2i
13AaHiTcn6H1/EDBhZWIRTejOsqH3bKBq6sy1s4ZBejM1KiS7qad/fkDH8e5WMko
ikylJCjh7L/GX2vWUxrME7NgwIygewwTwkmAEZxIvusp6bA6k1vqQ6aSq0BzVslB
rEr9gofnPtzlw81jxc1tazGJJ+ZrKvp6hUZ3nKaZagoxtNTLKPy27M6tzvRSVyZH
CyBcYnxEU3VcVgwacdcjSRUBKOESbFqXaG4Wv62mJdjzjoIMejctr5Lg5Cn5FgmP
mrAtWQX/Sdl/quCwygnaSi2oGyH5BKeiUKDpdvEr0u6IZli4gc7ks7DQpaSj8c7t
5Jrxtb/41zs3HsUMixn+VL2HmLsLKUsa5oOYhc0Vw4uWhssatHrWDdvwbQte27qz
/02nJmHmIqL+j7LmtEUDQNi1AvN727pdCuw3A+KUxo46i8xMbYsydO53fTFLw8Yf
n8CE/5KKtUG3UEIFhkti+mgoXtTtcC8rxszNnyeBq+EwTPfQxdNs/dzOe3cTJA8h
9R85j/IktHazZu3ptCEbSUv62xURajJx/YFi8fK9UGiC3Z1qJWqqFOIiQ8fWymuy
4Id/oP+MwSWSkWBUc9Rr2xb0KEzTTbOPcnuK3/Mw8Dt8mlNTUgGGGb35NvNs2muZ
+a031adl4HOHjPJyglddpVS47t14bESSig5tBNEe/8Vja4NA6v5kA6iGNg7V3BYc
YyIr2FM+GNSBSBNMf6+zr1UT/LG99maYFxNdlV9Q2Foh11CULdQRPEPUo5bHvseM
OSU64wp7eO1bK7CIw4si7u9zGrQSrl1v4Pl9fOJu3KGtOFmwLQ0t3OhsSGr/nrG/
4bikgTR/4syZrbIPdubMmeEYFG8CgltHnM3wiJXtGWuNB18wp6Horo8G2eW+fXlq
nU8hvrEnL1g9NLdEr45vtunMYF3/DO51YFpmezrFCVAB1EI8ndpj8nZx67CpQ/N7
nUb+c1KEjqUoZyfAEbYRzhV7auASqQIZMR+eu+6ddlcndsPff1olBv4+7yw2icio
I4Ayd5mXoEPFS2fkc88x0U0Dl7QJOd8ecgmhibUT0OEDrQY8qMGBvoyOmj6PKCs1
V8jD/TThUUKWc6vQ0tQLBQC3GFpvemaVgXpGUc6Vk1EVW9r2teeyDikr7OvJLuZ9
ayn5eoKnAUZES5Y7WhX3IAnzjuTpy6b/55wcbHvardeXQZEbN8pgoJzMRyN6AYKl
1tomfBeZvxzX+5qpNmN0i98caGdIL+ilEhym0uiru5MTNWG/Pqo6HzmDumVvfV1x
FUsYGILBCHm5kk1KhFFzkId35Af0CyrC5V3ZeowIwmfG1qA0VTNlLT+PISJK4IS7
ya7yfK7bxWZ6g+NzI+S8HsWP7wkUaFRjLYKe301Uo1ZN50NRtb+oTdCZ8hZpVi3X
DCgZWiD2eydC+TrSGEKQRTvD6kDORIImsKsQQ/0ActhOgwmAg4Hgsvee93s498CP
WIRstyulmX4Z21yVpn/olvTiq9lCU3m5LbeJ2o2MeDCwwg8pXwFG6aho9rX/7VYa
iv3B3EybiWbkraU7tVdZhYc+XPBp2u4XX7SEWI+iNzugXgaseeuVp/k+FMeGb2Fz
wctOU4RBBbgTKt9Cu/eq6N9jw+7INisiSB5PkK8aAOqAvjVYpOexnbC6j9m1Qkd4
UgC2HUOVRHF0deTUGAYeHz8vDmFNtLBmPNizPWXeB9FASv5sdxTyNOdsq3OTUDUj
`protect END_PROTECTED
