`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzuDqpKXj4Y508ckaLcotZdnjx5rUFyMpTiCoONIvxfCBwrL8JqJdCmWA2JlBBG1
DBpRlEZenRXK0GXbo+nOOx0kOkZU061l2nnPiTdJH01DAV1cSHIsup8aY4sT+mJ7
TQNeb30NsvySdkXeY5SZPjOBJvblzPan0WUnNps4spi5uvpACfevlGrU+zMbmQPC
UcyXcUeBUh6kYzP7OvWO4cxmSEDKJFeUY7ka4C5z7WwuqK0BHoC2ZUwtAJWGnN2/
+IZ9bpO3gJzGRdD+KzAMoV5+LRnVXDdn7TSoi3r8xtk=
`protect END_PROTECTED
