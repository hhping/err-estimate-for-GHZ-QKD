`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XyaZiJoAYNiWLOW1ScuFURd/5j5nM+ez5z0Q7VkRPyBV5+FtTFJp7PCZeddCRA1
MNgDe4+8zp7lCP+Jz2D2Nsp7STs+r3FEixbw2+BltpE6/poVOijE9Ju11UXG/yBa
GIjyzw62fnOgUWwsYkgwro4YRAyDKZgu0YOy4h9w3gR6jmD9SG31cukaP/vRHzGI
OJhw2hgUqwdSEHvfJC8zOJ0eoTVteEG3pq6UXdSuakMISMJ+iRQuW8fJUjMfllYf
zOPJIfP2xKtYNTuRYrzi/vovfhU2z/o351HLEFdIwyczfThpW9PXoyIk0H9VQkQt
kTMspnn6bzFytSy4XKM60rV6GRCPj8ybm7cb2sjTnwQ4CR+iDxLd3OVDqIGBLWOd
OPcAgJ30Ps3w9FgPrDu9CUKyyE0QXaE1Ub7vDGuzfbbJ0bDOOUCrByYF6xEY8tE1
8Y5KNzG5inqQaH+s7G2QD+bEqWwa+WxMnurxGVU9rrrfsm0p71D/f/DKYaYcI8pi
UeAiunLpK/f3gknxjlqTI7ZFdFJGbMdWB6uf35fJ+w4jtXHS86qiHLE5H2h1JpNF
J9QjuGJYE4S/kkcJ1evxSWLdAllQFZggjof5liVTJAcdhk9llxGvxqy6atdBTzOO
SNKRRX0qHyrRxDNLj/i3k6reFcS9rMuwDemph75eLP07lM8kM/a++YGFWLMAIs7W
fRApfDuKAyRiic9sqdTatYdu7KruM81IZyhgHfinZaVB9JI5nlBSNMlb47LIll4a
RyK6UDLHnOzlRhSG99o4i4TWU9HPohZrBNXKeswCDP/C5NFACImfUtrwL2+HyNK5
1EUCKSoP98L2q3RnrJzOuPW1kEPxP3qXY4KagzFbarSP5xx/FZLpZQbLtNMfcYYF
wg/A8CKNoSiVeJ/XztHqKXOAroi8MSTDgB6jGMyKtjBfmY5OChER/WgpfUT47Gyi
d8/EZx5vUGDRleA2T1x12oLm63XmRXXT8/KfE4fi4fljVbVH3KOMkCWOLYxwgWMw
U+PHbV+nAXSECl901MWYT3TIwv4/YZ2+chNu7Mwk8poDTAAlVToNWeVYZdB3qrSl
4zDw06M+LbruFr52bhXHrUmvnvnGwqHKoZvYCkTA50FAvyCRIgMduom8Dl86A6W1
LTbNQzdfmTCxC7MkMGH596Tix72WhIud37M6tYavRm/8xwlZl1CJ+guxGPkLjh6M
8iICm7yDni0eHEsXtxnm7Rct89gh/p5q4nJQZsYDgFj/QXydbjh4pSnc1YSwiZqn
hYOQx/MqWi76Hvf2IpYwHdw+KEprCHLcCCxNOsa/Lihd6ILRQg5bJn5C9VDVIe/Z
NbjkwgZlGW4IONawN31Q4A==
`protect END_PROTECTED
