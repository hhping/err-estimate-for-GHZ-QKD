`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jPX1yy1b7sfhlMuuw4NYHz7RAHCHOeCfPhGN6qPT2aCo4+jIvbfm2oxiPTJLOhoA
RK+eXvFkVTTukwiKFZASJgnc7tGpGGHFr95WsGe+sQ//2VGsi7y2Cstzalraa0uS
nNac5UMr7ujtRs3L1pYjBPKjInVEpf8TQABWfnYv8TGUIEb/gu8zeucHhuvM0vrE
LPRrGhd/NrUkXovbBN+wIGs8HQddIzKPDOQyf/nHnD6AM65SYdxIlRimLulc0Er/
ZELPnwrtWzSuS2bHjNAW6WDVBEyogpSllWOx+B45DJcBJuKR7LlHbqcmQzYEtufQ
1Cab4qIcVoT7dZCfC8epbQcIQY6vlN1KlRXcUklvXjA26aK+AcIAZe/rhOs8/Ma3
HDLt6mIOT8Eou9Y/2DN4OcHjl22zSj8jedYOAYOsyP7sALwC5Q3OEy3Ry0pTgHFG
vrips8dhAoi6iSsY20zNP64PlnZB/GvRPdzWm8U3PKEe6+xpTg9KtNLAFCAm4KhF
1oGL9TqmuVizbhT2jeyRi+zKhrBEZsbXpFHlH4bfDCirw1IrJvQJ5/gBwx4N0bi8
`protect END_PROTECTED
