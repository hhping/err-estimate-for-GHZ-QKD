`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1EepMwaytm2fjbjm69YncKh5U8hOvcT1AjBTs1vaB4SmqFLBxjoxIEuyJOsL3YGG
PAUgQgj/hfEu0yxhNxDHL0XQEOF2wkaUaHttfqT1KNcIRvQODq8uMIC5T/TrRfio
b75wgf8ASo5UXCVbSduJqGXsRkLc1xkQhIv5CQUY7GczAk58i6djzuLxGUE2jCNt
fPvXAdThwAAawWOtSCRrvUaDXEaaeewlF01v6x4+EdugkNhozJ8TRqDxsJYt5Kfm
TehEHt1AD2cRiZ7WEZziyhAVUr3N5yFlykjnyn1Mi3Ri/eMekaufrcBssV/HgLX/
51QAg1mxWvL5rjltsVCmpkKjxIUp47SDw6pyOAN9UAVoOqL7IkHz2vwParK3sx8j
Tu/DEELsTGxJ8jSzil9GUukVM/lMNMpKbWBr/Rg5k9dtIz7c8/MuNAlLETOK8/il
uPtdqrW4W3UIzXqY9e34ZiMx79A39Kuws1XB3HNKsGOtg0Kxcf7I9PN4zyPNuAbD
FpJOBEH9Rhk8ejXXkP6G7JjrqiqTlJywOwnmDZkUIQrQ8cYKGJsWREk7YzxfpkwH
eme6JPukYflNLVTqNiNv0v7XGltGHxezzCEG5J8AEO9GL2Owmagl+Jw2yNuspVsI
`protect END_PROTECTED
