`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjGEeUojbOJs13nWuk5s8o7IdniAwyZkaW7CcHBEE0OpNWe9PWTFQaiqfmiVeupv
8tfowDTyWgiMJKpvBa9YNp5a2aea+6QOLGfnCUnoK4949Y0AyxowhXEHSzi3ePzt
tUdeptpHbxg7KeZs4xsyTU+US0oPfOGXAwsHs5/DG7DyKSyzIoUOi/H12i5Vs+O0
yCCVteI9P3QalMF2goTEQ9fUyk68vpTaZMld6+0Y3sCQHRQ5ZIie7Jwh8D3e6283
EdXYaxDHmXbLNvg17WM3tJiF6Lf7TreOeRvmKgrLLcsKo2aevTw3Mea61+tE2X1P
c39L6pGfwqL3mDMcca/DG0/CoiZa3k3pF6DXSh2dYnxLx8zsz5aO4JdXtGbCZve2
aS0Dw5JEpgYZsI1u6HjRypHb1DZ/zfR0zcOubR/iFF0ZjnJ156zS2Fzw+Nz7e4vw
DSntpzr80tDWGZs34THi/LFVt99WtEKr0s4992Z2NSjriKwNde8TWJ/PSoT96adm
xhGXzk/GFZHaT+MUzypn01b22AtR5SMJg1x8hsk+Z7M/wx8SB2yaBPgY2iiLJ47b
xQXIHDpX9D2apCXvTScBecrTguiz4T3NRqH7KAqb3OsbMVYH5EOIQfUGqDKiEzOf
te521oSETDSUXs02eAwy2kucrir8gu/BpA9vrcsbOy4a2dGkjP5vIM7slpEz8wzp
Nb7scBRy6t2AhrCyLewXVQ==
`protect END_PROTECTED
