`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHWfss+oipUCq5FQWtUU0Y3tR8Bib1VfqAZkwbs4fhok1OCv2J+XgcyRXqmAjw2h
jHuIWm0njMji0votysa+cqoJC1X3vl7ElQd08CXT9dVuhNVHY3DY+4JsI/0a+Z05
x7uCTHLBlfHOw61V5D5muz0Cb7otKdDsm3w+odPAV5BrJRgXJyquHynTnUXdxLrk
LSwyMh11fF5jahXQCql9B0jUzVPzraEA48aS/aHmBTnpMKPbN3tPAbh9/zoNO5AL
jLyZkrJkMmnNzrX3SZusbQ+ae3B7qU4Wd225mH8k+lSzr3mvUzJD585e8rd0djvu
MnSW+HeegqDjuyHm44+fW9rbhxr1uRb+RnLQJg1C+VhLLx/U6FRDLl5/A/+Umptj
9PORxEw2HKYOojSxHRGlG8MTDriCiWcDW9mQ1pcwRevxcb6dLcp9E9jGgQ7qFg+K
wReGi3URchx39v7asofm/kNfeCxNipx1LPmSkNkxFalEl7GxgdzIo6t7Wq3oGERS
IzNB832ldhnl1xUf4jVKiXX4a5e9G7xcN2eZrsH4KZs=
`protect END_PROTECTED
