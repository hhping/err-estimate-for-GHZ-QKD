`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AhcJv9i54FcymwXTxn/d26YhNsejlx+Eaijv57Bp6KBD+LFu4NtgP7DfRfCoIlNR
8em8IaVrSoEjc7wYV1mcNJlEt6zh1U/jhZxWTnA8r2ohEO/fheJ2llZiwjHTtQjX
LTVavLiN8PuWN+Wo7yr4t3Y1EGlBh6hQG/AIqlfJuM9niXas72IXpJr1N7E+OU78
CVT3FD5n9ntcBNCMcM7qcMq2R9ZYwR5gd4VBmhxxDiWz9kNRnCN4dtthHftUhRx8
MCufMW3yL2DHUILxbe/vCGbyL59Nmt4ZR0ej6VKq6/NYLG1jE4/A2jUqnXVELPrW
c3YitfZvuy/lnXpxRSm6Ed4bSyrqUXVrLgZKwBQIuICMcgzBmq9GXILXL0CJc+BY
rrJsMAGZHYkmWEjV9b39Px2YYXEnP22zFmRxgKrVShWn6DbH0fzAoUOfNtALl9yt
l9OIsn6jKshB5D0193eFHfI/73t2EKuNC1Ddq4nOD44bhL+me6DGqMb7tlQrKDFc
VKqefuiuzQ8JDQIxRFHuU3ZqIpL+lO7zdm+SHANhu34JVUFemZCDkictf+8gtzOZ
nhJC95cYa+oK/WTnm+dv+eDxWTiCmffVROnrBT9KRRAM83fXH+lY6jl/QiXgFgyA
eu7jyzApd0xDfGQ9d904TdWMH3/gw0cj1UGqwBr9Z7K9LhHWfiXRlHqsKBImKdeK
pDnSbLplMW//6JdpXU7z5qCZ/zyTXrXWbmxl/pWZwPMZtTaYvjr7F2OwrocQHGHn
WV8Oeh9E1Ox/hMXcEu6KU0h2fRZqLW4ZofZrna7lF7bnVf3a7r6KIS+wOj5d8iG3
G8eWw0m/9rm0zKDAFxvvAX5B8vUDKYmZqYrlh04klxJGMCd3/QCzEbfF8RycLLDo
6SMPsZuym81qVL9eyyyln35w6zRjON/TEzkQ/dTyA4QrpGUPhmzGVJ9fT+TnY93H
SlBYtLEhKVXoFk2xlJ+rsHQkJTOmdNrJyccQLWzZuLoP40L6KIImQLAZPuhFJOT4
CN/HhCjfn+oDZQlGpc+rR/V5ZiY4nE85T9ZrXR2o7X0TwBoVk9F9sUb6l+QZuRb4
DnfPILt0MQp2om5WvHLy9lkLAkThG37kRdbom0MPQpPpF70qTwoQqEAgqwsz8dAA
2L6uF2UYgiHB7d18YE4Oqsn8lUupLpXOMb+e7g8zrMGKa9uyT9D74slMa0O3/wl8
pA2e+psOUPyGmlApXZeX5erlPJhxkj+i/z1yd/FSTEAQ1H7Vm685of2V1RjnpuRe
vhBYwK/735wgKnH/KPYM0bf2Tmt/iWPG2tUS6vMpNNYiokQgFsng59PblfQeNJjm
hJPx9szb1zw0VEUGgIlVX0a0gXSEm0PXbwK1e9xxAMmfwpaLSCOTCXfWVKHKIxjh
w7lKPYAXL7qvRd0AwOKCWTTeyrmMrVe2uXpvGe5N0yULKICFU6HtiyoLpV/bbFTq
pn3oIgZJAAyiSyRSryv+1VA4erlmWN6Aibdi+SgBeCBlFD+KCDZauFkNpSN0QH6a
8ZUzrfYY44JvIljwz/16TF5NdxVeMPDJv4Jd1Z2ujb0pxKNbmRS80VmSQfMpfepM
MxL8ybEhhjxmc20BDQaQ3FZnNJIfCtcfeEpF/v1/1mVA52F3lEcYUlM6L9sPhcUi
I99l0RG6sZUwJE93rX5iH1p5NoAXFQeJwRiOTyONtciQSdTA5dNRMlgoXkYoJQSM
6IlbnMqE+vF3Bi12iGyE2wHmDshYW0RIVEimlKI9XVEffBPqWiH6n5MG3ZYYh1LL
SU6SjyHwgTnRcPvaf36wpCUuBzlCbOX1DK4sK5Oga3PeL0mjLL2u33/33Zbbr/RP
l/wvjGIH8tEvbg35WwK4WzZ55sbvri33e5DxW6G9adTJEk3Gu7FAo/B8PUBSv95E
xikpsYUPpiQgjMAZy6K2jaArzXNhyc+KzDvvfsuaWp/Cl04/gn+OzeHSNRD/elUW
2a6FTNCZ691NxDmNrifPM1zjXDNfN0AIyS0oFmNpa9t7ydWFTnmBg0NV0bvN9Ql9
ru5v1vvjkJ2vpzwP+ReeZO/ET3/23pbMgghdg/hbdzgF33LqrSEib0iaX2d9Hm5W
LrHLbBzQhPg4Kz8HMvc2ZMANNjZU74myG3WwtFgS2JSxBpz7SrIr7FBOYPTL4Ud+
D5WhxGbvrLuk9xHhTS57ccXvOw51uPryCnRa4XL0poRmwt/puZXeRYUGGBu9A3LE
ZnjmoamgCFcmLl+FRHir2X2+R8zjf9ABCuYBcpcXS+MlLhgjpimGa33Z2DBgvrCh
yEPaKSdHS0bgVplxHPBVp4tZVQtrMPLOY+nIqDZjVzrzRxOGrGw1TJqmeavRXt7Q
M3luBNaYQHd4vxJYGflflQwYrqVqNLU+ptxeDO8MrzBaAqflKpKK+OKsYej0Kzgh
IbKZI5URsoBGykYeVUymD6dhFgnkMuqwAlG0S5o4Zxn/BCbhKdu3XS3hkYhp6ULH
D7qqr9mkkN1a33wp68saIoPh7sqNREtOj8MbwaDL7nm+dmBHP+8NZU01/xM1v2BW
u0IaNjzWFbUhpKKgPyBekE9L6pwkdrmc7Musd30XBAA6Gdk7F5pWEztOUNhzNq2P
MaoH8YzZyBRiJET4K8h5UqooCh88GKYh4JQ8pEyBlpLls6ASzGarpie0nFKhUb1n
D1JRDB4KlMBOFIEKhMlnhqEyy4F3PSFVi0bHVybGGbr5AMqe1kv8SI8BZboJ4OLi
WbdDyL1vGlY5KzZ9Pg8Ku+IUG9ss4XwEET0aa+3OG6fhNgleFLI8E9myFgG55UNe
xaVl3ZHd4d+ZwGjCmOhpJqPYWXPcWB026loLVvm655UA5YIdTwbGwrpNoe15h7rl
mVrAN3/Zmp+k72UXS4QGiAmugX/AOJvza0/r36mK+otQWpzFHevAAqjRVwWWBGhd
HzmMSJRxI2I9koxpXoonhK6bHP08myhRvZ/8qwSk68cXTjM32PWNwZMKoDjmoIpy
B9ZIPwvUUmpOIN383TRygjejoIoLX5itnEJSxIX8d3bXkpARZk7Cp389Km299Dhs
j6YVhKVM/HewbLWVK1LFMdZe69+xN6A8/LdSAntVFkjhbUSjNFtqpfgt9GX2l8/x
QnGjR1qohZu8vfQH77nyYdHGbxIQYet5otGhZiu2zrzezsYnd0uKD7vbDiq7htrI
k61NeaIwajBpZIdBkyXyfoReuFCH8NoMoc2RxCaHKLPKtmRIfsokCRng2p+e+Llx
w1+KY2FYqEUfkE3cYNXl1DAHBogg1dCAO8ZKWpl9DaQ1nRMonxHjPpzK7dYBRDrR
zOeGMDDgqBCy6S1FPVtylBm8PTg5gvQXcq0yBnmg7Za29nt3zd4EeDosN4ro2Lmf
O2Gk5M27vNVZON1AETr0fWaFyXU1IIOltFJml8T6jJWZoBMfbwE1aaOLbkN0Wg03
2Oxw8gD+xjarYOWDPIXDDO5EeH6F5+kk95YzsIF3qwMTPC0+rs6cwp8AsLw+uE9+
9zFZG36bAtmoE816HSTMimletWSELRwOCqZBp9mu8Jc=
`protect END_PROTECTED
