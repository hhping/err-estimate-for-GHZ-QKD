`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qwJNAPfenh8GKZXlP2LDWS8+6LHGsIkiYA2FivEgQii0fmrCZ03L28xWA0DDTpzQ
4J/U45oQg9YS5ZpB9FUwuJggscis6SLIleZN31jp/jM2ha9MJ0pfkl1GqiDP37VG
3oxEsT6yljbpvUcDOUNnbmBq/FqZGmt2w04eK+5tTzS7PldsV12sxSTfHYG1FnAN
xJwJhP1PkoYs1dBIMAw1DujzsgyWOUd4gH52dFEfywaWFze2HisECHas/1NEtj8M
80QN0jK5nOEXkRvL/cd1wiHEklklR5OrJ0ujWMlmxRI1Lk0aHh0bfsIT5Me5O59/
14iJzq3yiLsi3zHcdYdh7o0nrs3lTbbRdBWuUb930IO9URVBBw49So74vmythWvt
hhPCW9KYpGitdSCxQy7nc4ZFfKV1CEz307d+IVHsiAfyZSHi7JY8F5mrJIGs/nYE
8OK1n2qRMRgJzYiza8PjkKILAdRP3kOvGpTNTF6Lk8M2UoUeRKxDwJgvKV5wTLXR
ZFWyEelMsn4TRRrp7s4qwPheRbRbY6nPY7D2cyQ49fZlKRWlTwzbxXC3zFfpjKsE
yOQERhIgyhmwLQ8KwOm/7bgTN0boGuEze+2PYb4AIJv7pq+TrahPbRynmTkvXdH9
koU/LjF0wFiNiBCbeoihz2ZojO3tUCYk5LHxeh8QFCzSA4nPiREOAbYSjyyk0DF6
PoX5oWTZ09AIY8R+XKPLoJRplIYKSeOfLboYDxkaEPYuW1EhbccjRc7o4JV+bCBJ
a65dKs5lJHIC9xWLrs32Vmhehi1L+bG2n2lO/F2tNc0=
`protect END_PROTECTED
