`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfe5oaUutOAr7mQqZoVONoDNKVZT/hIP9qzrZgyFu03wAFB+4eMDWLjDCs21w8DU
rnWbPXn9LRl5IK2EKywxOD/kyBhiaZpWQeCt5To5MUMdjIV1gKp8YeB+ge4OCfQk
CMa6Q8b97jqBNzsa87D2w9is058bf1SPmJ2X+KSTOf7CIYdg5EEFhmrKCq4VONff
X9HWW+5fbpWdy+2VnzJURBgKSip1V6Yu8z5dXKh6NurUGQEndJUMpHF3iV3NbDzk
n9IEPBIMNuYhdKdGOsQlAij+bVM7UC7HzUpVAXVGSVjwy9DtImRxPnrs/EnNYdKo
j8e4CEymDAsv98s8/s2jTo58hHaWVL6Jb4eVu5GHWm6WvHR22gfm5Xv0YPEWmJbz
HBu+69gJGmZn1bM5wlZgcrCFKHl1e+970Z/ElEM7K1QMR/JbTw14ZK09XckrGVcZ
6PKRd3z1z5ndLIT6vL6vvL4pRXXaZBIj6vMOUcWyyOP4FqB8vvugMkW3bihu51lt
YUUkuQLjVPQKYpC2+ZHM6/fwD3Yc1QCrCU0Nl7CiwoQZr0nyyaBlsMccXuswrc4Y
G/qsXwE+ptU0JVeMkeVpUzXnrpyba4IuCWnyzXk38tJ5JYnrLSubk+XrnVahvXcF
3qs+pKq0H+nwmqP9jv2EJAFRsGaWdD46ZDxLr3T8VTs9+3CLzeevvPf9jEtWW4SY
4iwTPSKVNiCOCOAXMUjLfGLvOttwW9yXUGIveTWp/0IM5CTreo0jPmnYY940vVRJ
DDQYvq2x4yGas2WXDt1mwPDffTYpFKbsw0heKl1WT2xNoKXv0sv+B3f2XXBo4O45
2SKBriB7jEVfrPyejIUi2memBK7vx7tEg9turDdA7oSv/5Sa+fD6vPZ4mcuaAiJl
iff6YEZVtsfmNFLIqcFCu2AqHrZCg8c2ssFcaAG2QM+QPTr8C9q7NQFWMyYbqhXJ
g6RBq8h8QGWEIR8iXHtsc3WEHNBh/fj9WjA3TKflMprN4YXLfR/xxMf7vL3lxHWY
kINDrPILzs46H3/8Hy6vnSqlrYz9L5JpYJqJmlJlhNI=
`protect END_PROTECTED
