`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IJsCFXGpd2B/yUWlTO+4CsisZtoH6xNl+UcXlVwb6O09yn1OEW59jsg0GsSub1/
4YK8Bnn/juaq8i8X8UhHvR8bvpR+vPl9CigBFWrs08D2b6OulYIGb4TDzY9VjalQ
4BU52lb/HrFRF94u5+Icr46Mfx6Hr43ZJO0rireMPfjEVrriiR9VF+w0eiQ6yNl2
84kDBDLM4jyokucSUPQL2Jtmw4sI6JLUO+eIR86/CzzC8DoOtjsq9nSL6abaTzUR
Hcz23P0iCSGlGzGLgbda1HPCwbB13h/0AkECKjPb9zC5kYufXIiG4tseecZvMojV
u8wLYYFcltCPMG3Mhsw6/zaLvZo+ZqE0qJAI4m1Omh7pgwvkcirvVkOtz7aS5jj0
/WVigwo6OuWXcqndhPl2ETFnn9+cOyhspKFB6/Bx8/LxLOg6aRnoKO2gfp/CN6F0
nTrPb2MHV+DYfh8X1jPISmKHQQE8lTZBGe9226Crb8yH6p/x3mdhOMzcupgQ8Hxa
iYyROMFzqXo4NZfd/tSOMYoA9ZJSwqou0oUDTcStfyaV5OUemGpQRgGYNofEpkoY
Eg2mYx2ukrRy6ir4Hnt/SwcSEhcsDZ+k8yk+HNqx7zfQALBHcJeIvRbfKIi+A3go
+Q5wwazmhhk4J718siCuE3ctBGcAfLMPK6NW/NGhnHWs4il87J0j2WDu9UqOIfJU
Q38fVhfydPGSmjGjSXQkMGc+1tBQqIeE7NENB5/2TewMDcxQzEVDNJG+2W1oFnDN
a9kNx1oWXkQwn2i0Kfv3VqJFHq+pooE8SUP7DToWdAjwlZ4uS1GlShtG8aw+zAwx
Sh2v4+JCZ6dRCaitZapaTeXKG/nsMguQKR2ONFt3mjaPHG6JS/oGkVKLFEr8o+P+
Qflwrz2W4X89YXCPH4FYBqAkB1M2oShrjw1o+fibQZkarvOeuv3icCCEBZiISmnR
nPGq8n95Z1DlWfaDf2Z17JeqjunD9UyHpEt9UUp7R08V2azac1IUQcFEgICEW2BT
e/8a3+kH+PHrbnnlOIYEg0NQUTNYJ/Z+eaQ7zwgab+LXfPYcxlWyxHcQNG3+EahT
jarDl9bEvGtZ4ENDJMbCr684NWoavD7URNTMwp+rufJz3A65N7ZR4F8wBg9s1G+J
dUkgjFhSt/mN+VEcjGPuW/P9HUZMnQOON4/O2DHmau4=
`protect END_PROTECTED
