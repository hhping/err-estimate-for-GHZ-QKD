`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X62ELWh9wDvdbEuvGkGWbTN05xKiixkdEPE4iQVQATdJON9yxN8dZA+jOSc2BZfq
7Vhm9vKhOmEIGIxeUqQCURb8LT5rvPXvJ1nF2FY4pwSIljLSaRNHbIRUwcCLM6dH
D39E+p7hYrxG9SBBR4MggAp1byIzdUgIGqNe05U73qL66k8IVpGSy+dsR0MYsrOu
gQeMhV/p7p2zyzQEqLmVDoiSKWKb9W7Y1en8mc3m4AaYJzNaBEfKVMm7mzcoKsb+
VzgaQ0lOS9NsE5wpOS5pqXFbOm/eOsKyEH28IC6gANzBNWo3yR0fM1XZXc51NxRF
xEz49NmYo/bAhqeshVDsPxF4Bbqm2OrrSXqNeQJXeUMh/Lxb4RRdzOBwfARDVG9V
s3oBPjUKqPKW+EQgkSknJ6XipOwgnN+0nbheKQ8dm6Jxp4FIeBTa17bnrOESZxKI
TPsDnikg+/W1dlgYttzF/20GaHNC+ngA5itKfZShPksICCuFaDwPEHHkbPLAQd7o
SfWlKL+zzC2hku9IMr1lMxzslUwFDYwBqxITqxKWJQugKWNaBaNhqoPaTBTQSMM6
1KTRceVLWgsYepZK11IhDTRgZMrvJitCGCZ2tFT2cMmRBKQ0vr3Vb4q0H4rcinY6
XZxI/skRVL1DggGu9wi/sinZxFnU2M8ZY+AeDUiF4IzxIKXfwiGyl9KUqbDnDpyb
so7E0M7RHPOMTX2yzMCfH6piZQpzW+Fub0aYoL2XEqBZGx7dpdEZ5h7aHXwEnN2J
tpWEIAEIFG9QllYSFn+rHtem8tJe6Ned3+PPw7GzPoP/ZBTPB5CrxdjJ/W7PNgd3
0dMTBKwe3CL7gE+YFKNsHCS3lIkdcDVK/+lQfa/1mhs3JnUoH7Wa2AOS3VzZqVdt
pcfuNwBX/0rAsb1dXR1BAE0cwv3PBFK2d9OF3+JdsSA/mYH5XtE9aC+wwL+FaXKr
fWMkuFJkMyWQy7Pnud0K5XgsbVdQhPU+xyBs4Yik4AISms0CGoSRgFmQoqdVN5m8
`protect END_PROTECTED
