`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INek03CRDGh2mSbZwcKFIRfQeQpSAOKOOXINluzticIhP15pH7t/Eeh72H35ZDm6
m8qI6w+YAUT2TeaLTaAgUJijqmXExYT5LC+EzG8YJfsUAO69K0P5O4pSGiri9rU1
zM0SPMyVPzjdPIV7dBEXIsDwMN0EqTz0vJNk8jbs8HXCpX+90rNuFervugcsDSRL
S4RW/5dnCA1L+5JY4brCkAVI88dRvcfUHItEjHwe86AaykuJiNHjK4daldHuKMdC
NngEdu5eI+d8D29y/imjF6MJPtAMi74i4fKvEbBMR3nEGB4aGjKZeXa+eqwbHr4x
PsOSX0T3CbEHtbz+y9hCtFmc2leATq2cey1NwUX49xWP75W+XWVa6b2FpTSwgOFX
CQEKGuOFuc+eCZZpH+wRXLVg0n5mioz9+Lw6t3i+NgwsqNLucFtn3Ygo2J2ayFQG
6LTLHU/buDW7ejArI4HVY8z8gJJVw2ilPTnohMvE/PPuzvP2uML1MGgXsk3NirLK
qul0T9SEscB1pJughCR0OB5jzEt0fSiVq0sONsZLMVuzp/9y7RTPZfcqObtAYqqp
MSAzDOp8vryQDOdKJQSxoZmxe3lyA8Y7E27LgwhD3qpT2hU6/ue++KdEpmXIbxnW
vm7SBfztnQetmLvfLvFMj3P95RqTTGj5U7hm5MGVwElMaITz3pmJwzPLvlG15Q8o
MCf02MlUg0kPk/sjMVM40aP71AbnxjpOzilkRD1drQwO3UpEDfk6G8XbOEZZsmeh
eDNLnvLVXwrALumpF1Cuj8xG4J4VW3T+CrH4F8bK4Ime2B3EEspaeLrBK3jhDel7
TkhY+TWFU2QkpizSVhoIfn+F7UJst7a9xSv12Xh0We5STHC3grS0ShhozqYGpXgb
Bv0A2CPd/1vlNH2GV1jF1OZzdNIANLoXsyQCP5Fs1A/p59qsxcMrDpkcxqdJiDqN
751qL8QgWDKyMlLPssANMZyW6V6kSD8d6IInis2IlDs=
`protect END_PROTECTED
