`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3EzKZOj+yeOwE0QuNtGEdH+H/xFFmp7YPll7hTDGx+x1u/r4xXfviq7hcrfuXcL
50r5F3whW/l/4u15yH3TEz99QcLuCWoS5z1RJHZjd5qbyTAU2xs8Kuo4Sq0ifcUK
x3pZoGsF5p2XsO2JqOuZ3u4DPUqxm8ammDF7oLfRi84VC2XQDZb77cw/bNZ3OtEn
ibOd/M+7Ogo4tjpZ/f1vTQqB5DvCRetjrS/qiwAw5WWwjfTl14X3Iah0NMgw9MIY
7TDtmm6u5tQd+0G5bg5Q/axlgj3QVX/6/HUT61kufhzl6wdRKuFePkiJ6BsqUJhd
oMqwbtRf/PyFwj/NggcZ0ZP+moS3GrrQAw9HWDlEaRpoSyQSR9ku57bCq/qpS25k
nu+uOPHNHfwrQq3S0NI7APl2c4Ma19G6guP9PX5Yg2wfD5WGaYS8YdLxrY9R7ijD
I00hHMLn7MhRNr1qjk1swKfnmWDcVlfZScruLo5ce+pCkz6opobvOjbDf9c+coge
1qCbqdLXYqm6RFl8NCGFwcIKdWOyKqmWx9zvT6+SiNdo0DysFU+TPDJNCkNCpsJW
bQmj8x/iPfcl168t4Jx0yC6+c8RNkqCWVxfbgSOSE5vfxp0Vc4K5BHn4DdU0JqGx
DDPDxpLjKoqkkbragpujdyo3+mQECkEZ12cb5tPhnoU/04iXO7+29Ah5TU9MHIHI
VBO8r4AhQRsr0DOyqNUquw9n5bP26pggRga+BAoxPeZZNSEuLNr6RnNfJ3tduj0R
8jacU2vlJMPtTzYN8rnXP+vr6r4HxGsLEKIgqLxN0JPTt/vIjNzo6ZbeRFOVeRK3
n56Wj5gcOBZiMWS2/b7mrWZMBFM+XLUJPJAB/9my86JsWu2iHu/uJ/8O1TqNi5ar
u+Do9U13mCZ4ea/vuatLlypPd4wMe8ItOkpyP6xWMW/toznjH65jJgmdpvaKcMn2
h21u2FKu9uObKuYXKLiEoyQU5O702pyrrkBVCrPWVLaV1rVfcgNdgVIrNmfM2IR5
depfNwfpe1UhZWSoUOz440HVk+ZHLywkTUJ5vLOFkf2AzBsZJpyHwg0dypE1m3DE
B5VeuoDVMvlYkl2JMJc3c5vEL6xN/UvNELQc/9hoDMvPxa6Ra2a+8+POVhA0lePj
lpQwhMOoVfBbxxYjrNB3yNwidJizcD5VMQV4mOuOpfMD5Hk1DDm1ourTyRwTnXOD
47PqIKDRJLWGRg3Nh1qL6Q==
`protect END_PROTECTED
