`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qc/jkv3UV7a/pjwI/tGlJ3J5AlNfK4sgvlO8mVsFKdRSIjN3Nr/0QDivgONd5XMI
2ut+SB47hwN8/qnPCG1uAUe5knDrCJD/Z0Q1tTuEPAwHmNCOGhrMx00sZTisJHF9
zG+OyRWR9kyGtdDjDq4F2IO1+AjP6M+vMvtY6dH6QF4c8cR419ieSLBVyRctPxne
IfJiH7xtsDv6PyXkkFDWGrI0h0crCoLoYTHEl5FQcNnZa8OeXb7md+SfzZpPCDnW
yqaA3WTa+Fbsox5QOilpjqBMDsAGy2TkVow3JA8BvDznrSJYadMUEC5CaEAl46LB
T9iAi6F62AW1qw6AtPZNLOCOiBpQ16Xr+6eAR87J3PIhPEHXdfdw0X+kR2TbJy4w
4wbxLcCmo0qpc4w78SXUkmOsfHs+wI09mb5sut9LdLYh/H109sQIeT3y3gRgoLYo
Zx9prL5pzwHsBFRQl9OYY0yNgOq2zxmRK2zAuKxGb5Jfk1QsVAMdYlEqISr5YE6t
b9m67Q7C43pt33YK+KwxC9VuU5q7IS7TmDMJQOmwtShajONacuQzNJcNrjyDsh0a
5+LBONzAapoPo2XTOxMyWyFrS/dXyvLgsKFTBqq2HXDAujkioDkDp6nlWlVdXwXx
Z5piI9TpRTWU4pDMEbOu17WLpVfRTQ0mf2soTp7jKgamVMG/LtVciZqyj3Ky74Xq
CAO07xw6zPJ8y/iSlHCLNqycUJIC8rdkRtzObiHNPZ8sqH3OeQjm/hbWszTb/gag
EE3xrQ2hZKcyx6UoPZ2K8DAgMSj9T2xoSpIBEK/jL110TOy16xB+X7Cg5bbN6qML
HMB7gktuC18PGeN6LV+BzvXHAbzWRe7mKhRSjapyvBu0nNVvBEZTuNphUlP4uLKm
FO8ZjtrsmIRvXUaTq+NsNw==
`protect END_PROTECTED
