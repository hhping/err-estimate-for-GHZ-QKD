`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFM5oPjKr4afsPPJpkslOCh1M+iKUH5PIBVzv/o8QSj9goXX9TdwPQm7TbqoRs0y
K9/AvZ8ch+fWGDQOfJH/7qEprwa57Ud+39WNQb/nIBldOAN0rJ19D/3zjpND+Jhr
3ppcUqpOZpbTJkhfAUrO+qNfyy4/8Aq8NFx7W0EOY4sCucfPm7djZUfnv5o97F0l
HZXVRGJYYxawoeQzmU3TMYamu+/jgoeZcTyUqcIXVWMDE0SdvgyxxegUd6t47CGc
0KU3kHT5if58mJiyBPS6fQHRPy8JfcYqe5rkVN5yUs4xflrb02v0YHch4z+KDiuF
MOy2la9DkGMx9f4HHF9JnWN0wbHNaIjIHwVq4NuB7ee/gas5nBF9m4NQC4PY1Zwv
j8m43TT0go7v5NMvqKV1UkdFAO/u/k5msVc1qwPscPGyugNCg/iIWmcASHyBnON1
qtgsNwYKi7pFxkgUlsS8nPF2T6uYrvpwHmVKTdopGWs=
`protect END_PROTECTED
