`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlccboAc8CLcQ3aMrqHCpdIX27vlicvc5cw8FW1PefrRy/v3dM2/sG+0hs4QV7/G
s3mICgrN8mbOPEkyLzASbK1rwb1tvRRU37gAYdYpYdPZct2aMRi0Mxpsm7DsnU7g
0VUcz9pUI192XZW5ZQz2KOqSNiSZr3irYuIk+7gmhDlu/43bWdZyV3JsuOGjfCw+
trZMZruwOGMEwaJl+AIt3KWVCy4p53HFjU/KkzN2hczc5ClXWOScmy/UDJ9fiWCA
eoNhiAgfLdUlDTxPhL5ih2Nq1pL7HIKPFDtR8haVmb+FYvEdQUTdWtkNmc0Elz0e
tUClXKYaP+npdyhFJFk0lSIW2bKK4VOVE54iQwHbYInKao8w60WqUoQhjMB881c0
aba7bJD/bwGcU0PBjhzXj8V2LJnpNMg5gTCbN8jhf44VwtPPfD0vK30LatAXIZqe
XMLVLFG/SHBNz6zBXwlaKUh/a/qjAHZzPlBrIUI9oa1BSxDB1OKc0OXSCfkHx3JI
JbiCVYZUkeBMfWQs5eQoHT/6Dk/asMCWA7jTYGJg25Ty6ntrBlU65hpeztpZ6nDw
r3WKwhHSSdonnZaxW1FEmXivejQ656NtuWLSwWOlyL+tZc/rYK1Rnzkon0a19eQw
vxWBoR8R+C36B68ETqRHYMliPvPzQ1JUeTVluqchqbSRV4uf3qbfwOI4AjEH1PaY
Y3TGjr7SoJKdAb/z4bM6OT5V1zMCesOYBIEVo+nU9HNPGqQE+ZvJWhCmyJR6GL32
IN85vWKYI7Wn/Wl44hwFFqgjN4bcsNsuFqZgpguf53IViAMrl/H6evIAYt+bXGG9
`protect END_PROTECTED
