`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ikln+n6iazHYrO1yZF6jdotEpT/3qFiz/EnBQd1vlobtsBDgomKy6Qa2pApGqXgK
FUN7XsefXZKLPPqi4kYhPrSvBZxKuErKqRYrYkkRyykJ74ZWrqw4PJCsl29rj6BD
MyPrVQb0IIBPsuHwS5SlwB4ZrKJzi/IEsTHubYQqoY8NSAKemI6MFyxtJuf1tilt
wqvNlczQ641Jgv5MWob4Wt8zbsfLerTQi4TWCRijSht4Qfk0pBYIw+qdrdFRPFe3
0TINRoZ6koHTKF/KGmODTDuT+6wxjwBZfGj3ibxrSgDSyru87FjQ+hvhgWdTBg1M
INlsar0t+dVLinfwA/OvF+Nbyi308i362KOtlBU2rLvDFgHnhU3CWgMEmN54EzLE
00G9F7tAlgrd8L6ljx0w/5xbik8LWZ5CbLK/ghLAIJnj9bsyF+y0hqzKaCEgqECq
iXEsqtlBr2tG81l3y6rOmyzAZ/NJ6aTtJn8IfwOR9Duw0O1d914P11GhL9ok9OYX
5sYFzHyDhsPz5EQm8L6EDqg56/4Zt6qyso/IrNkhG8v+JPaTiRMDahn0Vtj1zDDl
BNRXe/cKGY5X69AJAgb5RSAXGvAuORNfJhxYgACSSU9nGihHsTpppYRfrMYNpT72
1zChYsVxtQ+Ty+l05o7NKex1V+Myr8Bp8EjVYfYngb8GIoHjSSs1Lz87QZ9nElQU
iWyl6CKZCGGZEuJ3ZQP4fzmO0jwhrnFnwVJg8KaHlNtgXeER9uanXg8gY/1qCy81
/5kWejnZR35dAwUC/bvc6jCJb6vPZTBvIY9A8rF7UV/FRj63q8xRkGB8pbedX/J2
Q0DMoHowRIzJvEeOyUz6/UeXPar61HibLzkX4mknDj+2sS4fdUQ92xu2lTi2Siu9
mpTBjTXHNFAjPv/sYHq8OJLwa3vwNZ7e6h6BGqdUzxp4XCdAKxCNYGpgsui7kamo
44iML49iyaKPiFV3MTi0ycWP7Z1omCQZBOu/HzndQyfg2RqikJq8JbG/Vf5kuBrV
tJL0J82Czdc/H12LCYnqKXXyqE+QI4yZZce4SBEVWt1tbc/1pNcbwpduxtqmH0B5
lDshj5FXNDsg6iRZZGdTlklogcJSZj0IAqVVttcGcmAayjBqqYfFQZAkGJsCYkjq
gPI7ULyZ6Eu1EYnRNFiyUwCU0eBZJI4l77ud9nd6//33KpGFgrmU0EKAgzUBf7ih
UjHFRGY/4hHqkYLAKJfeAyBunLv1DckKT1RXkEbfmlvvDEmJsl6mwgDyqapopkK0
4bOTSExSbSH75MXmR6+0977od8EUzpC5J4unmE2ynC3LFwKTX6EobVw3Lmjw1eAf
2EPJj+Mayf9J87MLflMYEd7OiWR8o6i/Ehg6ggfC9kc1M3SGqPrm0UGueCqzdbMq
1s8+CfzSShTI0MSrZLX62cwnB3K1fRk6LRXg2DFGTYzbhGh8tKPa9248RG150vmW
9tWFx+pTdzzPcBcKyO8x3Zj3o4LoLWaMVZ0BX2O9ZOXH3590cfi6OWXNAiCFJvX2
awoJSy01LebANFdNKRbQV1fUtJUtaSpjUlGdrGgs+roUV4BVAhhQrULmoMeRH0h9
aZGxdz4ULVIJbgXbOLF6VWoILjH3at+W7JRkUDtIppCsy1ARv/sklFaUqKWSTl+A
Q+Qcd4vxhyTA3mRqhu4JIjZbKCoKZyPqJYktbPN85uivyHc7PJ9816VieIpXer0D
vd89YFGv/ifeGofT+DSMzjloOX5m4uKcvgIZExFmk6DubxT6aw8fV5DUyd1Vr1MG
M2hDjDBVT2a7Tk6UnG7AH9NEWXJwU2F6JVlOOhmXQlyUQ38iFjv5T2EBTwiW5Xsw
XmEC7jmaa+K+5ob7FXpORBbbN2SfTvvLyUPuzn4RYVI1BfJS97PRQY9o4Pkzrs3M
JI6fHszudrFYhuAVGwDxT8HLM0YxJ1ONtOEOmAoHKaksd0IOjTcJCMOylB+UehsX
TCeY816GIgM1KWqM+m+8Tshvc0cwwDvfBKYXu6ItpFVFcKMH6o7wQ1JO2Lq0rXjg
BaUR3ep2eMXQI0P3uORftOSSpl555EVCu21aiy+jUGWLiPCuc8iKNLPLeVWEFZXg
rMpoVeFHllodbD6agj2Zwk1wpyjSIqKPcUwRm/lVlws6bfwxDV6plM+gMOfWRatq
85G2kCJ/FhJt81y8zGm/FphUOtgMFtMKJcxWtkfphyRWWnodw3EZllh65dIh1E2Q
UEL/5g+201kjmqO+3aJRJuhRJUjg1clEv03Ig/+Timeja5tZH9U6YWPMzYUlRCie
dcVX5gYF36p7gLMO8P6cd3w2RO8WZN74JRxl0Wig+Pr/zvfHmhf04yXZDzquLSmT
0gbnGLYVXms3hbwmAcO0STgmWKeoJzrihKeIl/Q6jfsBpmQDHD+R4FHAHxeAVDl7
GwGpcTBYUVtEWsbq0GuR15L3snmSyZq6QtFRXwBOXz7hJXlPec8+qH1Vai2GBgm6
H9ZPUcccWcii4Ousl0V8duPlLSapJgHUKro5mc5YPUDKGBFDSJB76gec+DOGl1pB
M+FNzVIuAIUTpPb/Mbpn12YUJB8Orn68eLSAYqCRfl6Mf5U7Bj/Goso+Nt+M9t2H
/dAg4VvXNaMCqMWz5h4S3DT3mpvcQa61ZoqmjU68tONSEcZ7s3ovk4McPuURBU+Z
o79ZWqFG0GX7HROW8Zd2gFWFmjfimU9ro3E5SoLFI9QRgU+BFYfwTebOdfKDBBZa
05JnehUQyIHlusf+3iZsvPohvMaErn9sC4qF5hvjjXSQMMsI2St7NQh+WO2Lvu35
cuDQjECZVfjw+UEB1oX6tiaaBwn5Q6lIDON2I7rwnyqQMU6YwFwSmRcqpfyy000k
Vxc4i5bWKOKkEcWUonF3YYz3yHuuclrZy8E7fVSPIUA=
`protect END_PROTECTED
