`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FC3ImsX12rDitiGYTPkIG5iTis+mjT6/Cprd4AGuhA3OPMGgTFZYOcQTtJ8OZpP
iR9/1pPxTbHRWa8+rxKuaC9KCzLGxDBcl6SVOZf0Wz9I6B6OtSwzk3lqqfFWhdK6
gbitGPsMBajDWN03tYY+KAOt+k/LIJqfRIcX0wj+1XBGyN2Q0rGyB43meOflgv+k
LwZCVxpkxA7IIL8z4/Og32o8zZT07CqWxS0NBcYUmrPz1aQ9/INJOwA9A5vxR3WY
DgGC8dF6+zCMysDhkeprSv6CyJMbr37U30dAkz1WbRrIEo9nf/jpbpa8E5qNhgGy
KD1Xyt3bueCuKFsMGafkswZ4bMIraWlfm7KrwZjanxMyDgkOZpeXq8rBsOhpdAB2
T84Mp/bjHTLJlMGfJRktF0Txw6eadQDB6VqhbwErEhpkintKcHE4KGvVqe7zSUj/
bR3gzT2Dx2qtrRVyPP4AUg0jwFe9P0kZ+2Vxlz/yWms+P82AVj7msK3J/Ln9bOz3
EoXKwN7LX1/25TB/Ryb2VrHLaaZmCJl81e9+0wqiB74mpkXRoCHsikRSOzRp9//q
2bKhTKY4iSpBIL8ZN5EJk5zhYyEt6hGfQtgjsuGgtUctn+f3vHHfdYzKerXdEOM0
yXxMAGMsIqJVUSnfbtUYsKhlEccmtob/4H09J7uJVZnYsD/TnEG6HktpKI85c20P
oebliCNBlJLeDO/t72nxnvfjcTCVcoD8G/Z52f6SD5LX0WZaWsdzOQzGGtt6rFSX
G43u+SP1g1SGnWLqrcjkd5q86Bib+O+wbxJ/RDflsF0yVGErqTdfRE7g5CTnK6ks
g5kMoXM2VXK9L5GG0QJH86n9uZggp4tiUDz3bNFePiIhVk/zVslmXC5pdzl4BDBj
GXWmW4QYSCf+SYAzQqUETo7KApT2ZbEWMObS8E/9fLpywwZf3CBrB9CqnaVfkWD+
S55wTkNwEKdLNlOVxV94wCJFapnMPahHQEmVhe1Z6GxRpCfHPXeGW6clDq8MDX8U
nOdIMZfy4sJOZZQvQ34TNOlcARdhrcITdiVazVYwJSkZdGaPfNgGJ8Im2VrDIjjb
34bVO0sDuP5xqOzbEcW4yM2TYT7xPYHZSOfjqb1a9uSjIw30LE0Yo1FXo3LQbJrO
Oo3IjZSnPRozwCXRAw/SZZhYqLcnGqpQPUiYJqbVb09b7sF5DzjasZAo5ddQifc1
VVtPgSzk+qvX0vlJnPNgWHAef0534s8wjKAlnrRBfFz7EdmxzTQ4Rcbyuv6hHcjz
59FpN/dWVoR4R5GUiLhYvj7YOFWilBtWf5NQFoy/RODVKhdtzNRisRHTtuSwzFQB
9EiLvzhWZSSz7tU1i/WOZlBRrguOHGLspnQzBbd5K37TLD1OZpCStHS46ecSPNCz
Und+hnoMD0N1YwZ016eBt1+dTQgxyKcBE2WrH2X/nUA=
`protect END_PROTECTED
