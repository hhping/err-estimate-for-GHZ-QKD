`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9MRSJkaflPZRXfmNaD1QRTsKLaZQQVqSZF+NfDfmnDChXD81TYR5O1v0Rk3FlHSU
rYCczOPnhvw+fMy5LHrS8YF7TVOvhdjH526P8HvuaW1ENk4YxYAtdMSHPlpl3yr4
41bc5lB8w6j8l7cqb7fQTzwhNH756PAUXk9idsavMvR9tLg8tXyZOCkvqXQjfqU+
32thHuXX4ut7wvDdPheBcO/EzWfsa88Ww1A5gVz0toEjDWHDgGCwjfMZRYWj+DBQ
7MQAXW6AqkvRqMkK0jQ9+r/kZ6gqcJMVE7inxGCb7DPcY6LIA6az8bc+wdTdCBkp
/4sux9c6wsqVwiQxyxlBt9ihUmKBcIVrXZ3dmnDcJDrDKT4PUsdF8+ms2KDzMmhs
MWx6KmIuGbNYYc80lAlcbgdsaQdNW+yEnX+4lXts2r0VxWQ2zwofE9Rt2c7zVrPw
fk+4/sl3O27vuZrjUHDQeqViLtwlpsDYKyeJIBSB3KsNZeMfFWtAIGOJdGrYEiC4
nVwB3ve40U0rZn4tCQE8cp8CyjTtz5Wd/MVWAzHHqJKE3KDCjRa3Y1Yv/5kY/YCN
qhnT9UjOfSBeXPwaogDwl7ygAcM3GwmljlQlI9L0FGgwvkpCe2BHYA8wk7kpuDuG
eO1bE/cQMd68Dyj+NNd5/s4wsoW0juq9pbbYajqTkre2P5xVnpn4ISoTPxj7YBQC
/Fo+GqBfPlRcW6rCSBjLeiqmatq7a17hY29nTPCSuybgIq4JphBytd6GEDyQR/RV
`protect END_PROTECTED
