`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXl6U1Zm4UaRvUfOXdJquobxX5Ish8PvHjFN9USexZNI5aHQYkJkeuwurg/rbjKM
HGbGuVajXOBxKHLzyQ6WSA9Kp5vDew8h7fsjg3SaLSO+hQu2o4/m5d8jl1cwK5ls
tp4B8QjehxSC3EPXWd7rQI2QzOwUZnz5oEdtlcva4wXyLKdZ3LjNjIRCUevfsRaY
Url74ezDuPdBzK+D/P+ORYPs1Pm/Djo3IDqfULIET7aCkujzJ0j79CfXFW2aVvro
bE3b0Nbh6E69tpzuI8iUeftpC8vF7Ec6j2GY37ErOXmraV3zuz4Zgmv5l1ayxotX
vMZSdRWIh/1g5iCenpEVzvyXyufvTd9l2tfwV3XyQ/22/TRxqvebU5kq9q+G6WeS
46rVfkWPOjfnHUqQn3xsYWXBrca3ucUH6su8qJuvl6eQw9v05PJPq+Xl0CBtgA54
kwyWLtch6+YuoPEUKJ+fGNmmOX3l/bJ7+Sf3cE9l6yNtGExuMY3BRmeXenKgG0As
UIA2vYfEnOoMsb5CWVqp2W6hko22doCAi02h9YzfmNZa1IBLEw3wijq/F6WAtRIi
i7owdijNPW527BxfkIz6SdcdIhmx5aRfZu5bQHvdIGTiRB4TdBtEVVo9uU1OSRHY
miKirZB6qkB7/cSDx2nOIIQJCObNPu/Be0/Y99vz5ZLgLZ6tmKpNXk0FIo8zGI9+
PQOBCLZEhFKRbosYH4eNNe+2RLo61FqGYCehxYrdnk5zKx8ud71u29s+szT8uyz8
yhIu0jo+cz10M9mU7bfDxbJrfP2oCRlr7570VglD8XSnnCFC6Yk5ykaP/sbgwn1w
34V7And8GUJ7qeTw4yd3pHj4aU2rBXxZceE1NLThKVNA/0IqR7Pv0NyBQvKDm0Rs
qvuXDJqZcx/xUyPOcGAf9jjOGYHWiVxyDn5ulqf3Maqu9SwNwFG2WYY7Z/QbzW1K
jH3K/NJJxQZwMO8PJinxMp+oqGzwWFQLm22JfkP1kk00yBlngV9JQeC232dNAwML
lbgMVtpFtLVwUMHgr+UAkxr3qMwowWmsvcz6LPqoEK5nt5WMige7zfNcLHtWQXfi
ozrGM5aSP0fs7AtGTvFEzI0XdrF/qarL07X8qdYiWTYFioLMl6fX0+tmDZE36IrK
c+5oVLANtsWvPLAJI/R8nn/uxplULX3jpEQ1zyEkDxvJB8M+advfown9tFJb6gHP
KI+8g8f8keQuv+R3bVz/6BinuZAqLAaNCIUx3ZWR0nxnnZRbMUxb28Ha5pqqha3l
Ly63MM19A9SOCTuwgmVQMSYD4mTNVVcgF7NUme3DtaeHfJ1xw0xO9iJ9Ym03Br5M
TSWw1aHQtaxokFNIAOq+lc7mRChwsFmDTBbLod7GmakS5kPldKIWhKQToD4bUc+5
c6VSin1GVXVXPoh0E5yBjxgoOocXuIJOXmbE91mJT19nW2JH3QWYGIWe2cC3pJjD
muzrHYaAz8OqGehrAdKfZTiLBJnyzwqF7+g8BmcNfT6xmgp4gyhwiS4Ntatd2wLZ
j55WNM6de2uBFCMw5yj4CvIIaCrpj4GXEt4Gbj3KeokKNKoD0acz6gbu5euO3mEy
dDsFQmkLapoydUu3KMwgXt07e7lBM0Oz750KzLropdfU9fGyyA5slwEPDEsbqHMl
3gh5es+IdkC79EnQLFRnOkaYC6HmTkk5WHPGNtL7QwVC4fqCtqb/hSmu0DR41w8u
TFmJw0Am1DxJdOgx61tT/N4BNaY3LP/QxgjbKlh+6QOKcKzQf6aaU5ANzP/iEqA7
sKeLLf1qr/PppPULoC8yfEFa8bzzW8HOljLwBwZ1bRgfFtw7ZjDNvYiM4poN7jea
SXbGsJnPy7MebXWHP9r2NxS3fnOiSEK5zHTVo30GvghBokct77eKH0ON7qy6+Fk3
8+kTs1y6msBOF5MChXkLa/kPbBeh36iSlT4U67esiOJeQ1dun2zWS+vhZzxmGQ/n
xjV35HJ3HRwtcMroHH0fk79GMVbKeMQbimU45Uw8w2Ha6QRSZwnkR7Nyi7iSbEkx
qLvbQ8ReNsye2NpDLWdA7XDvDyPQjSVYYEUKXJpjsTDTijyEjeER3/3kcVyJ8Tq+
PiiEn+3udY3fgfiWqt1D6grLsuR6BrqSuf7gYcMwRCnmUFc71wQRHuaRUsVD3BC7
XNxgvwdzfdgFGCm6pBvNuvZT7wLPVzFFeA7h1YLiXZ3DGNC3hsS5fNMRjt9mr9Gz
C3VhN1gQIYOGjCLlRdCPqIP6cv83fkyt3i1HwJaOLi/wvp2ft/xiwmLQ9OxJ/VrA
wpv+8s/AHwzzGbNcF8f14f8N77fiTW/08K3EpwmbdPFzMk4AuGDrMfTMBixgtSWS
s+MlqnA6/ntuwTB7IyiKtoP5Ea7r4z/RlKtdL9Zvh6mpM0hy4ToZ1eZjfeg0epLY
RursLQEPIqTxt+DJ+5eo1fZytTOoG3boFgFBeYNQLHQ5Zr8ZBKhj0cY2Hfdrmlrn
wffeTa1GADvfTFqnmLmFadOqbCiCONSpSYc+ayVsemU+GPm7zwDfo00viPYdxEwo
3K3aeDF55ASIASAj4SXVywq9cI/VAeW3IX5qbD3m/ervjOjag5GmmST1za9xMaI7
L24uMVAWK3zQxKHEG5Fv/ut2wtdz7VGeG+gmVRtVi0JhUQf9GqQrbjKNqr/LeJnT
4V0x+GXJSLy2hoZ0ZY/Kd9y5U38d+ykc17kV96lNU8acAl3hZn7elrgwuU+L7LRX
5NB5RGkIv+Ew4S6jyWUmLjG6weTYsJBKyxj/5IzrKVuKF9rh0w3B3V9r0Z8adyrz
ZUaVdc5Neh5t03+0zho5ZqpYrwfzypqtDaTJ5MoP6g8eb0NkMQYoptFT1vAxOYfs
n8FyvTEsW61OfwkAGtzkg43SiGmEcHjOVtnODEW4nMZFmL/XwmjWE8WbBbkKaz6r
bACVJgVv83H+OeOIjRdQ7LTdQhPSophBN3UxJzigIQszQx4vH+rNQAUkawqpFjmp
7Monya90dz1t/8vltcY2kzZQo9rFT+5iAP86GrZIdKYaqUHFqinSDv/EabsRPqjj
1JTkjp3vaq6w3pN5/2TBpR6hjXO3HDRjpCXy0k0uU+Dppe7VMtnJyRQPaUarhD4N
lsd0u04IBgRgWGXBoqyWlGESh74Wx3Gi+et2+aCKTe3XsjaVj9o5HsZICUeGVpnb
Lnnldgvv3l+JfqaapryD/EzWNY9O4RJtIaV/sMLcHqYPB6Jql8xkX72OTXmcCnAs
MfZihBtlPyEXdijwH5w6nW9pzCUkZATGxdzVQvofAWDJdiFOGs2/HsJsD+NUFHF1
GRROQ/5/wP0FNQKfEvl/03HHeUpucjAEQufz1Nzb2MBC7xxHidcfWPHGdCHNIe7t
ri6XX3SMvWx287QDvp6zAx7IyeKKyDsyeYdAf3VLbo6vk347Yaau1CNh+40tHcx3
I0yHGJAVf94k2oKenQm0EDUVurBvKFmsLmX6RKa8MhnZvGpO/EmwXCIpxMPRCcCk
7lLB5zdVFIF6evz0s38wXl8XrcG2u/ZMd0nw7iaI4WeRnILXj5ggsRpva6geplGx
xL4/vaT6OQ6Bvo+manO/+dkGyFlZXddggDtSv8nQPuWtObUEMmBDKjnUxhaqDs3F
0fhWyYTa+LSXUpRLXlIffYljT6Og7MUPIeiobRoMzBX6buGATo+W8s2PK83JkUJ4
IBn2dimDQzvhei8BJRJOmvUtzzmdu8ryef3/vtQ+NKf8oZepvvHn0xRoJDmZDLZI
sayPUIqkjS21zCMkf5T6Igob/Yw0Pcy9uiIOEcV9LtULN1YsYRi96tVlN5v86Krf
EreU/YkC2Nb1LjR3GMLw2XwUM2l5MiMaexd2iHY/nwCNCiC8Oot06PZfjpCbJDHr
MLvNwVBYY2GKQLUwzRIABoWk5R8nM/NpBrzvXbqSBnIAYiaJgO0rR5rnsFWGsT9r
D4pAXu7uyw70FwrRiIasOPwRv8OE6VON+lqapBEX6ql8O1GFlXOQk4nveePsfH4P
2BjqMm3UuWJ2GWwlUYAylbrfNiiabwcxdevRe7U6MyjhDnd5pXWiApmB6WiZAGrV
+123MTmzOK9XNw1fvVo78+MUxpiuurVulQc7oag5WNdp4QV5R1Qixae5IvEuLRgq
FZvI0WlkM9TIc19y5UldfBP5oWLoF7cUfQe85p6OJqOF4jBSzOV8i4v2y4325EHv
4ZuT8CXOa0+yoe/NiIwKAqG1JjUnpq7Vc2Y+1u2xDjOM/yxHwPgLWgIuzfm0kYK/
L6JMxZO9bsIxWDlXKwVvmeAgA5cUSrBHXx0UClfnbsyFgSfxFvw4UFxRvRuUJy6D
fyMOw2EzlUl0LQDEt6B9NVnoDS3CzqdaxzwrbdsqAnf5xf7YHT0HzE1JL1HqbDub
sQnSosmUgCsgSAJe0FttBcNPX0euN+hp17FOG1CLu+RKGtkw3PkTJHmy6y+mIivc
WYwyt9joEf+b3NxAGmD6aH+bm2z/y8ewRyMRlEzoG4hS8QblvR9MulwBPKF6F7Mq
bEPreohkMliVvFH/AP/+wVizetuu8Lv4BvmN/llTRNC/97QR/YD3+4nAiYnW1yCD
3imrdTcNkIcH/wgYkx3K0A9M06R3Q9HgXFFT824w4Gp2wC6j2UxWxYkaHyCCCJyP
d6mLrImg2/goRvjBQtpeMe2iyK3Y40iBo/tBRSwY4BEix73hyCVLte8TU51nYbog
mtpDjj3vOnA/t9MiGqWmJ72lieqAinWVzLPn7fyR/i9+aQ1Rf2vFllD4aAKJDn5e
AjV0ioiO1lfIHu6n0g2QzYeOjFb5BntL9blZU96hVnOgmHk3UdD7xxZRRBeC74iB
RSUgdstBLOos4FO8pr0hgLfU9aOMwz1xElvUYHG8zELM5Y/jnlVu9cktqV6SqkPH
MBmRJjGVjjK6gOG7OFq3DLAIHGRFzZsIK0+qCYHIktAgYMZ9HVSig1qdY2jv5u5F
vuSWwsO0dBr5DHiWLQgDmBkttvuRZICMW0TjyGtknMpDG7EozXzF553QOmTIfvxt
TkYUMbv5SY3yAVShV58U3d/dse7JobfRcvD9V7beIHpojomj+H3XDhKJFlUFdoc4
SzPcYCsiFOESyic8sH3J7ZSPHmzbzCFaq5UaIO4MKa8gOct8yoPNSQbzD6wpaC0/
eyWIgfbYhYZX/HDxuZ3Nbtf/arC+gS++8OkqlAmDtKIf/47xWzVQ7bSb2DcAJ1OR
CHAQIFLkhQ7TvwXX5HpQJTqNmPsgDfyE2Jq/22HXWpQsgEXcyHSHa5zbgQTYySWI
4mPUJyKNTeZA/1BG8j0uZxCz+i0KUchCYZZpnU4qYYzndGCfItJEKwpFdnEopwlq
EmyiNPIHnE1aCClX+L5wXioKPZ9VrCK8OPqXli4a2Dj6ABygB2623Q6cjSrCC8SD
/O8zJDhCvWljoU6WTSib1Vr0RjL2hkNAmNlW0gNugxc4SI1/JTfjkIYVJ3AvXc51
91xVKt4yPBpmml4lW+yxEg4+W+95u5e6ZGLaec0uV/eTRX4gdG5oH43tyRqMg5IM
yYT9OmCyry2l+Jr7UI7r3oeWmmTaKN6inbJH6Hhxck7MPjAHab7kPc0CuTjm0gPh
0I14cyfcdcIdbwY9naNvGbHzFpyPxNWi3M1okRMlvgm2a2O79TPsjx7bskTRUj0P
ZUiJkyeEKlBfX8bP4lLBBUr0eQ4oGO0KbwqcGJhWQV0bVRzHEwBLAZ9p6cidujhD
6u68+S/NOZsObpX2DwhMG5/FjYFpeeZzTIMmbDzUDMJglyb7dxeHK3a2foTXkADu
0BXs74U3EtjyFb7xkcRc8TT18gj/LuvdqrJe9oYFdX94hDvNscuyyA8SvPgpwDrj
AHUcKd/9BZBLGNNkgqUwL9NfRo3BJgkcanteh+Obf3D6NRHbK/EDwActFPfMwMP+
LWZcDMfV+aW6QCbJZxw00B2cyIIUD70A/E2lp8lpvzUeSoF6Rns6j9q1CQ/BfqXV
I/SKZIUTJGE37Z2zg+nC+dBuErn7MFiWWlALLAOquMAksdqN+LsHtkeJLt8yJPgz
0yH4JWQdlc2exXrNMAFnf11rMENOCbXOGcvA3lxKQbtFWr8R2P6xgjoeRdYiw8rV
GYsHxDWJVZRoZmNQLe039/QJEG2ILyUcxE6nvPdlEfaRyX9M179yiFZMdVwJEr8X
/XMNyvxUQaSZr8FTTexnKQlkOUgxsaFwqMP/ctxJNmJyPH36g8venmPI4SY13I2A
IFxeCl0tiQlpYkA7qvFiRAAuveeeO3lCA7ShP7K6zVULsyJyT4U/n4dXq3Uz/fGN
mhW6CvpM+0vQVNsOYKQNKiV3ZdE2nvaM3NKQocJzo/LY4M3JM62Zz9cRv8FuUd2/
83kb1lWDnDGHrEwnOq902QwBf6JRnmK2H09ywtN6qkj9vJ/iBl2232dQ5cL7S3bg
mnKBr2MGInI08HAqILk61gJTVyc9JE7aHpf9K2U6LauPRKAIjttMuvdLNUl5KU+M
7UPt7eS/s/TFYbGhgt/QHx0JdTqgaAb6GYl4rVU0Yj19TMqvrGbXYdj6k2cIMVAZ
wGIp1Z3i0cSajRpKLLjAkMTm5Yx3RRVmKKu2fBQwMPcMDk0YaB+Xw+a7Yrn1eAlV
8b6u3rVGGsHo2WZardnroUspTXC3p7Iuc+CVQFwii26csQxkGlciCr36G70Velb6
ppIGshxePXdqPXRqhgvNkGeKDtQStFQvrhP5PlgSwHgRWOVDyOh71ZXY6GbAaFx4
ezTyG4qU7H+Yl0Qn8SeU0yibTknc9rI01NuMr68dJgoWB67vppTh0rpDQc7WGZRI
fq9UDZOgVw+5VBhJhX8GX6xdg8XiItsVfYzzEN5C9T7XAsjzM/Onkpp5GgHGa8D7
3mHMLg+lGuhPBXSuqIC8YnguwFBP/tcIpI+LI1yBi/XmvkJUW4zTSnpFrbm2hJcB
gaJ2GTO3uynK9DSCkILPqoMsmmocBxBtYWoq23ygv9NTawHuTmm1u+JUxz06HxWc
HocQBOhJZKTGP9jZXX1p/WxirNJCQEkp2aZSXI6AbTq06hR8BZ1EYHfmH5Q4R2D+
ObW7ECTg4oPn7I/WgEEdorIZ96B+9Y2G0KOR5pGmB94ZU6QyOLdxXYOJSxxW9yod
uMF079AqqEs0uIf1jbbS7hCulLPBXUPNKhYlLrCQ+Zwq4TIw7eB7SVtVceLF1I2Q
uF0/sSBAR0V4j+dLkCBbw3eB5JhRrKdKN2SKWF04Nc0Dhf0Et8VDZnFXB2vNHKJm
uj0p5W9x/wPLuA8BjLW2yltnwCaC9meLLgIEIQu1Wr8LT3WSc6St59DO5aILt2vw
sDTMrHKOxr7VcNNpJhWlYTzXP4qbe/mcBnaiBRPMQ97LWo5foRKAc7kBZmhptvMl
D/BUbmcPcek0V9vpIKqDOB1ZQY/PxgyivIA2gCE9vJNhD4oOGRDj+UF3yUCH0psO
lm10uxxZ7iOsrNMUbpTTEvL8wGHQYX8szGwZeGQa+TeZ7s1dvqDwfaFuIqfkTIf5
yzs94S935okXJlq9NmTMWkqKBMxbMcpkCG2RIyz/GXBdZgzwwReMEHanSJpHnx3N
GqIHI9LvGG+wZXE8pGZNMGZRTEe7Rhe2WAkaA61iKXaO9FzgQOHSlLj3DC8xQWPp
ME/ZMacHyMdZdPvU39Jb7xGwwWDZtS3Pi1kqKGlk9GWCpowUgtC+89TWThmFvxJu
jyCNMKSqMmdHH9AyF/6smnEifWFCoSp5i2HkefvZEaIG09Llhb7uDBIwN/QSTg5g
zhG2Tk5tfpWIMIgCUxFSy5Q7dcAOTYh9VIh3RVTAFYq8Jcty6oCFj0+xhOq+V90F
mnWK3+tm0Cdz7sffv9rvQQyJth4eb8hLvv3/lq7IbMBORFJa0/3WFgZ4stXjzlee
i+EDxLX5KThh74NIQyb5rH/UgtcPNgmnT/2VSou7wjKJUJQbF1U2hL0Af803VLSw
j2cvYocBwxapY7ZVR0kZYE2i+8kk6tEhh1zwTPtQVwMJGZyj9nRs3Gl7/G1C/1qk
G9LDB2pBVSTsy9ior0s9p9C9rUuJ7m9GBZxKPSv+LlsNI9QlnU+ihslsUWXYIkUF
m32APzTK47/Vtsy+V3sVeELZT/M5+xO8jcRwb7DyCHL8gNTEmiKANM2YPUn9x9Wc
una5ecyE+qQPeZ4d1bkN+GMUg6QRzUQWR8HSc9KND3ys54LqrurD5FWiEg6amyP+
eTx3qDUg0+f7FvjFitJ/zKG3XLGZs1y610JeLxLY7vFxO3PKvLx1qsV61paLmQb4
PBG9HdBcnt6HGigwyjfQCrftHoWQ9wPfttibRuZaFJUw3KMgXUxaZXS9VGfB/8Zd
mumotzAXTYqzcTA/ab9ntUyyE/IHD1bWNt5gDehyU7Hsruh+oBbIxXh87QpZaeka
QH7nGjjAzXok10cs3PwSI17SSo4SPhAZE7myDqyQRpfyXbx2rnnRjp0Dda5m6q0M
3jSUMOChEQweG+dQeUcSrck3UOZIbDWChCIAPl4sDX/r+JLYS86a/06MP3oYE27G
3aKmyoGFXXywA0oiWJeA5vXJ6GHFpZJnZnJtVs1ObkWMsXSQSEznyXOnYf01EmQ2
Dd1C0vq9okuuB5tVH2MnayGVIzx1kLO6tctS780hZEqOM8onbNz0ZdUq1luBrSQ2
VPTelf53Pn1idB5rrH6339mvpvvskRALSp9G5ROGlx9K9yDstfXprzmzlPo2XD4J
c2RIm0848XnftV2Etk4N9aE9rHYtaDQPHPOdV4VWl9BiPQ/fetghy/Be79CwdDxv
ZdQDTfy2lNSRAYaJ/rv0uE11SjYVrYL2ktOgq1Iq/o7ioyCshqS13RSfOyqaVHSZ
G2fHOl74ARH5tD9svsMa17C/7QWOnAFL3XRpu+8QJfgkjstuCUdYFm1yRJqzuA0i
z3K3ot0So+Wp/+KhvG+CYM9iiPfPF/R9kWX08/cxgzK03w/E/Q2z7yhHS4ROxy5V
`protect END_PROTECTED
