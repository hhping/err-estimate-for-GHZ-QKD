`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKDOJTV4v1cTXBpQuOL4QejRNh/BaNHJbIIg5p/q0T5zzbAqrmtpKf/rYFWGtPJJ
99gIzxaeQ7/n43oI0KeMSJeusaexNt8VA/q8YTqZ7uu2FsL8cUD7eCcaE3KJIyOK
XxsL1Q4UsJUwdH1CfWSAqwHqNxtwhi5p83n1JD5ren9+znxLCDzYWf7gzRR0JJ+Z
DB6dMF+1TTEfbYaUYqF6izFDtfawapqlCNUgZJaDSgWRAcPb+YwddxBUSXcA8XM1
pYeyH77YzMYsc1LBRC7al8hBmsw61kUsQhHy7yG3ngFBeHGIfhZ75s2GoCvSQlvr
fKNhWN+xQZZiCjTrAkZTy9baopkuKg/zLMHGsft0JJxCJUk2ct1suN7IgcjY3ikQ
XmIOf9oTF6nqltwDajkR3w4PieVRrlVW21K5o+cnTPyZhYpgRewKYa+pyuHJ3zsO
JM7JxjNpzBC5LzE/eVssqg==
`protect END_PROTECTED
