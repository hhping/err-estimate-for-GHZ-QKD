`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efDzs5QtpflW9ISnNxQ9ZsCyM0jEuduaN2FrMJuhe4E6IR7YFIn9/X1Q5crqOIyq
eHhDBFI6rh6mx0bqNYxFdXqoXbKpiDuAGB+FjMmDP3B0eiy9uq0lvHXkPKrM1Evq
DRUPMisSvBHdkVLHdxsArsYuIhmOU3C7VHxikJcJdfp/kQz+yFZotV1hAf9K7Wx5
xJhu/urU3leidElifNUSJGpuHP7bGQWrF/4kcHvb42qIMLmV9nYwXgGPC+K5L527
OSR3TGBFv1wtwabjq2Cq29kuBFDuvewpVp3panmU4MhPfTiJ/BfQZ6X6aWeusMCu
vZ0j5j3MpzhIWFtb3xMhXdg4NVfqOnNVkxzE3hTORbrcD5B6djyePFxUggW7lCtY
bS1deNxGp5NCimr6UnGxhXQPiCOQ00wj9aZ8HlCrj9lVRX7Sw1lZP/s4soCZcD1U
K1crOozY/ozQiNE57Au3QeDXI1RgNv6asKCP3V/znRYbLIDuK+GxMJK7c+4ANwdq
3/Gc+ZirmqWUlMmxX1EcUrlydV1vbV7mVyy9CIbKY6MyBHt6z1yP73fPwfbV/LC0
YaDom5uIxmVhBpTh3yfkZUG5yiyBGlIwIibrDWW93lyc/tRNgO9Zz00XNaBk8935
gm6jjXp/LXbULsJad7e/x15rchNEnWtwXqsj4K1anQSXqdnXFQrpHvBcAwG69h0q
bFFzGn4+p0Hjy04VL9AjfMIskuLQRR/tBmoXFY1bQC8gHyTpGLIeFAQXXqLw2O0k
xVsaIIrVFDpXbdK8lb7A0UM/HtKxc2eWyK7fri1p3OTrI7zm37GX14uCMt/+L0ex
2KtoLf5zTImeNrxf+g8GpRttfnn9Sbqbpg1ha8Syed+j+m3YfRXqrzzJA6G4yRwN
PRb6oNobXD0/EJ1YIZYtvdgYZ07kd05GYsCZpiUHA1LRuYUe2H7/Cmgo3DE8anWU
eKaugQS12DOKOsRMWSUVimgRq+j4k/Op+vh/anBHN+0wt0Ny9MBdEVzdvao669ef
QDUCbEkHbVHYl8yDKAsCLtWU4ASVS8f19EjMLue/GzNj+9V3e20QMUrRcpRRcxrd
84AmZyxoMO8cEyhfgMty0YXrjo48OCiZSw4uMdcOWfn1ruB75uDesUrQEKyHt37I
rlIi2Cj4ZS6M/OxPvoASZUM/W4UB5i4aBGgvIb/H2WD96hEs3Mjk7TL9aSF0lsTC
nQqUCY1ZJP6PmrWPUSsKntXif1PlEirsJ41C5bmoo9zfIrQ5Jnks995SKg2bpbws
ONCRz8u+w5IncPmgl0nC9RuiMaLmjLynSUvzQUq0V6Xgx5w+2BwwQyq2Xhq9bDE3
ic7Ke9BffSpiU5IP/ObKXegmRajRiItK7jJ536L70atqS1tUcF3VHPBZ2UMCKjB1
skFiC5FT0YyyD/wYGfdyXJGsnPIWinq1iSAbjlb0AHg=
`protect END_PROTECTED
