`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OV88Ac7DmhBrDiEymhJaHwuZJFlFh3pQ0NbA3qFKzPO24fLOkclIDOYOXEMdu9aM
/6e/HzylLG3BFrR4lscg0pdNJF8hUyHNqf0rv10TmTckHum2Eu7PEIab2TmSJrrZ
wvB6xFrCbudwe9Punbc+oGczgKjTf/CtV88lAOuFDdYcGUr5CBkAv1l4PHqClv8L
xeFrg6XBt63faFDjNufNUFhqm7XJFYyHJQaun+UILqZKUMxA83tLSDGLzcFBvdwh
apNg1/mspal6oqwERtWrUNITpH8CiG1mwkmQc8fFOjvvGr/rP8MHCDY2UrSEImZ4
1ZnWE3faXtDYtP49CAo7Qv63Whx+Qt494wMezvs7xc6HqD7sE8Tq85/OAQYK7eTL
AHvkFagVl9O6snw3DXBSabHEGbqoXWsc09N8/i2a+tv3NuWmoOJD6WXQjW38zBjs
NhNAO4VrTAs9VU0QLrdavghpl8m6nF9FWYebCeIHwhcfo6MOzKBHEl12uMDkeVxj
2MwRlC+b5kVgj7humK3by2S2HQ9Cn3i+eQkte9dkzhXSyWKKTUaj6eQlwq4tE7xm
pKGBXBRClbzZGIgQMvVRjIXJMDl7e5t+ffyAuKfNIfAmlli6kQLR9ez200Kdn0GV
yoOKOHYn2n6wQwfFcsHolqzzCAsAe6UcTLiZhVe51hbJ901+dF+d90rE3YdJia8e
OXIa/9QW7wT8FufyPtYPo2xGeFGrldjmwn0tbWwexISDfqDa2mlAuVApB7FUAvSf
YWKI+6XGUTAGnyhEILB3NUBP0sXFzohphSMmCZFpaeuKA/DvnTfSy5Ct6XOHgXVW
rMQETfDu+STomGbZbm8iLhqUCvfxf/C3B1AwjEV4s6jCKSX5kIHxpzMVnp4RiPbq
7nMmkaDYLHWEbVCtzwwIgzQkncjIYlnYbDq9NnvdVendxhdIcAteAZJlrJ6+75t6
P8DOwcdLHwRC+X/Bcp5EuexCKt/2M8rAitKNj1V4cNsg3Q5RmvFOGrfctbx7P8UW
ajMp4aLt2rJJCI95VjV3HVFc4KHLUgCswfD/npc3il8wFCWjGjSPjQuY+6CptkTf
XP+snESMFjhNqBkC5IPe8ZuU0fc+cP3LLRnJbmm4W7kYlmMNhgUHQ273Kb/JWB9s
`protect END_PROTECTED
