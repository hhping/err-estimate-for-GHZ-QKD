`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ajKWAAEyf7Sz79r+lAQ8QmkPQhGnv1IhJzCeX5Ac3zui/NcjtJzwi74SMMPvVPGL
GDUpq1CDFJG4BXfU1XK3JJZTfqjoM1OXRI4Coktu6t7MxgI4wNv8w/Df3/2x9tsZ
WF/qrmd6BJEt0Blu6Gv4TctQFcSsROpeErgnjomOthlv3LKhquh8DG8ZlfG5ZAoW
p7RlRUACZdduvr9XqkzACVn7GdWBJwX66nQXuN3gbv/EfQLB/AmPSYuXrO8IY/Vb
7vTdl0++qHAK0M0i/JJysdliqC+pkFoVs76HW6T4P34KaitObZZqRuCzsWxQJzAF
K+SkfRU0jKZtYOTzql3mnLv8H/I/7Gj50bFqXhMTl8aUbmNF5YOvjuJD5zTcTw3F
AanH8Kwj89Uda7tyucwGvlQOomRNsOailwEJAGO6H5/yXOzbHe5Tlm//H0cXmzCG
XLNBvQrsjwnP9jMzDg/3x+hoNZvO8bHHoqHkYQbsvh2ycKWN2P7PCY0iAB6LptXh
eKZSY+6ukm+I89HPq//Gm90JdcZzTutlv7WMIBsklRHSX5Um/ZkRYlTPeijSv7GB
mZzPHx8oRdW9YQk/x6I1WOi7wmDxDQyBtcz06KTvsIfSYbwEfOhtEjhUMT+/eY0a
UoF6Huhafa7w7tcSyLPwwbXeGOWO6iyKOPSdVJa4fbABaZ0oNR35zidApaqgTWul
et3hdWqfIv3Rda74I+l+43uKCns/e1FDb2TVk/N5L+i/+6JX1QGrSuIDzTP4kfRF
tt/Pyh+NkKn54YQoxqIcjEfiyp/wPTFUDbm77HWFGInLubKi3hbEaUCbZW0xS31J
gLB+yL52MFh+fE2m/kmbksK9YLYP/vZTC33LtRoPz/To1KjiBSMQKCIdkBlIFdMA
UzSCsrwMYL7DIuVh20uFoBjiZ7B5hkY9iN5I0O881v7hE2hIOtFHnx6/I0CApj6/
Am3hkp5GiI5Fi870DBX3F8XVXWcAEn06cds/pWL7eShqSjkhK96ogNOA55QaHCUT
ZNIgW7omFLAGPFgfYyg4DFT6lp8QCGOOWukTAM5m1I6lTia3cFoFz/p30XnVow1w
/IQD2br6Cj5N5PA0XNqOWnj4e3PDfJaeqvi7HB/j0i67OK68ODyyXG+rmEtq4vFg
lH4CW1SdgXPrNvqEXbTm+g4mBuDq1JYOG85zt7wqY4awkSYx7t6HxV3hPznl4jlF
FJUPGyH7ZYrXPy5S3b4pNH2ybSTW4YJ3UiHUsZLe4FEAZ/IMLww2VnRAo2rpt2i9
ItbXLNkkU8Lww80ukl/QfXxjl7JlyI3hDYXAp3xBkePj7zCtf4g94c1DKlE6NMG2
aAd/4KkURkbcXFypyK3H+KryzLDPajyvjPw5Fk9Dlc2UhvQBhmgxUfXzRJssj30m
Bbzvcbvcb5Z0dP94WNu2+ETeQp1qaJ3MKDOwCootYo6IVb6JFmz+8OajyQ9eNAEq
9Hac2O/0GJjLOmfn9r51e7ja3uExXAtooYE2HVDtDbb+2AVdap6A2FYaLouuzC1J
1Y7r7/wFS9w1bCWOHSGNrNY/hvwUcBOSh1i3IY+lm9LhocbaGL+GUBPsG+giwLMa
9xK7QkWbn6UDwAiBL4bkAg9xdNaoxRT0xeAjhp/f+6MkqlfoGJVg07xYsG6Rn6Y9
Z+3rO6GPfyeFylccfRfegON6z5FEV14vDmbtOY84eEil1pB0gPSHzA4s6fyilFlk
q1eL/CRHCcgNHvUpCg0azhM5CSj7KRZ5/vmO3XRErEqrXpRVyiJC7PMtifpsO6yu
htxtZ6AftAbsn6VP+1ZyhawzP720o41NYxlYDWVuZwhuKW0Bk+ujvk6neJqrSydB
N8yLF0C0NOJjJd2fG6kXpwIyHb42U/q8KbqnDpCLS97jxrYxPgvQYtheOMo7dJ1F
A3hSYv78Ra0gg62SYuy7FRhTy0s87bThWq3Tez2P3wzIcwsn0rCZLmV8p33ZEznl
ZtoZqzMRMmSNlfG0F+ShBB6WvwVm3lxOswIsq0swiUYuiAsB1FeUZrLUgEm80OjR
ThEShrvknftIkvN2V+vW07Xnv/aprw/9v/4y2qdhCrr2clGyO/K/Z2LR2OyHIszU
k/yMMZBFihv73v9u5O1vLzV4AIQLxisZpIdXCzANFJ4sDbONa5YO2EO5V8mqtcFk
S04GjcGDhS7wAxBOt5cuX2FAH6VlpkXBXavG6KmXfVYilc48pHF4rGudMZlVT6zt
zU5J70phXtcJD18qgsLLUr+cjCkDQfJ/bYcrh8nSXd3QX2WYKRW9zKaBIXr6Gt1A
Cjhx5nX09RcYvnl9p3RmQSkNRHjKLklj3cIrYUAY2t1bFHGELv0hy+xzSIRaUCHD
4/oG9Yyh6SCdMKWG0MpoowbeHlTPWJT8cP+bKjtg/h/cVvnLI/yLpTiIW0opHPOt
8wfiyvGfXwnS7TAy8BbKLECUwEEHJFzpfllNtbMcbnNIY7/xc8m8ZPgmRbdd3gYF
+4T9DS2GTs4A1W/RjFRouJE8bAFdIiCJSyP86E95dZZNV4EKoOA/fZ5CLvmdXhyP
fMIgnlaKhZVlYPn8ZswlypycI+xhta0Zu60DEUXIUK/l7FlaSYl5HbmkKAlYnL+A
LDusc/CIdmSw1+XdN8v6Pa1vj/xOLtwf7wGSXLFrRL/2s5KKQ9heSAwwJ8twkhuP
Vlnwkd9Sp8fETI0qn0g9slPDwfjSt7cZgH9VrhPwwrMzA4Rp0xUtcQ6pZ9CSovH5
NswRbS5Va4ttCnVYDLaSVWLLHbRJJmyB1wHphU8kFVXmS8XMJewXmGPEhgzMI0oS
orYPp+jrZh4OTKEJIpDv8bKShMW1UQbTC2vhMgmgt588Fwdun+/cTiPYhf3TzVlz
wbEvqUani91bBXRjOkXS7VZG6TPvfLtzkjmdDy5p/YDvEHv5kss1r6YsHiFfU2vm
3XKbrjCJ++AaEsExaSn5l5IAAppsP6jKuWYlXXn8BAx6crGMY0CpILt//gp1OG8b
M3CJ4Q+lIMYs9Ex/wb570PO5QG4VVsEra9IHHghNBtET65Q+RL0UtuI04IzZg1ub
YCZQbUcA6v9XCVKwFxRCod0Zi2BoJ7U5OMnyUtZ/CuaE0YJ64OpenhVleNlSFoMg
A9zcXmprZEAiWzTmM9mr0ZVz90jwIjAc9OPYPmhK2hDF8PEkc9QipUrRa6ofPmZm
Ue/rx9fHJ2eqf+ldkUo/1H8lyNV8ogs+sYPYRuvZ8iazPax3HDVyjcbX1zhoShk7
W6dWFQvGj8UhKrKc36B9so+4E4Mf2tKV6B2v1FIQ4gJXqhNiRp3VuRiMxCcp6EWH
lOJ8inqk1qI6lLluLG5h9ugB4fis2S490t3cUFBHxGS85hbYI4qlch2e0pj0CHg/
a494+grQCKu0bhjZtyKqY/35SN916WkXAhRnP0q2bmf1AGgImbmlMVVYNOCDLQ+j
Q3eyHyw2UiiZHkD4fdHg1Kv8aZ3NMXcSZ73G8bQZfer0PzxJSYN8bhdskLlcl1m9
/ktaFOCojj0G+GSWipOs7tTFagTzmBri9L1+Mz0YlGVHi29hL+WS54LQU3GoHHG1
wyzR1SGt7W8/yuUaKGAvFWXYS0lbTWgX4K42q6PPHhhORy/Yg87NAv7z/yGgIJSr
WmZ6/Mbi7BxaCILjvw/cjCyihKpq19yDtlozpJtL04AD4yk8kj+l+3JbIWxLgfRz
lZDRHQju1OggVfds9+hqSjtqPau1LgQWbRGSdhDnmLfvSTH72NbvtmJx4ZVlsbHY
hvCYOHHqT2X6vA973qBBJsb2tSUwkZEjSqwV8WvjZ8EnB1GUUyydZ4gF7+T47D+M
IOubDfF8fhRvINBVAcFKrxWiNibVT+DwbxfuwankSoM4ouThZ6gymkIfVHitkbl3
8MDV8Z1Pwz0/kEH8rMTZI+N4hOOspzwajh4QJMktJQo6cMg6DWJifMR21MSnTOEV
VfnPQIfEoypH0OAdUZhVRL7PxfDE+z2gaKAA4QPTF+ciB40hYVBNw1W4pfdWr4Ul
e+4OKWqdVvSIW18Tc9201kyseVQk2sAfJOPHUIDMHPPaHB0GgYT8TSPPSoF6JX+2
8L0HGH6V8PkHZX0Pb+c4ouhhIeEMzXuUoWyj56r+BxPslm+THFQDkQRxfXxaDQDV
D1OOyELbxbsbvSLOfsWCm40Jc3QAFt3gn+trviIASM9Oz1moFGj6xxpM8zpjWRu9
3wWN/lYfw6gmDeVfT+K3+h0eVc20rjiPOigfNoJNW5GUhExMLmg+VjruAlAy/XB0
thcxkXI+444amVWJqB9Hyjtwa+NUxuNZ3aBC2prLh2tibmIbfBcmZf3i0aPlhrRy
1El/ktHp8aX7AkoBZQ/C3Lz4rhTisrjxXyEyJkT82lg0Ug8jvdCrc+HWA6m0ctWi
/y+S4/hZi/jUJxcGi7Q8oM1Ak2Fbsgb+zl04P0eYRH/qY4gbgA/4zZOLi//V1zcT
8MgmCq6ezjAzGvJt5e0osPZ9WpIlt8zplOBH+i9/Rg6n2Zsvliwo7RaxTHbwNd1S
RA01vLZ/lQ1A53EEjrRMj8L+LCtj1CoYrlvVeyJ6nDExQfoM0cWU7r+9rz8Q4t9R
opQ9s4DJZ0pekndK21m5s/n+YC9E/awEpjZ2RmOB7LiNyMjoIbf36/wfj5GEcIdb
zAPoFrYIhh12ctNeBSkfVpAVYrnu0aIe0+VKMsuaQ/dQIw7qDYG0JuCg5z6u22Jx
Nd85PpLXxeIbNv0oXwU11u3XpL0OfJ50MRPZctb80FVv3rFyZDUsb5doTWhrmZ10
gQ/3M49xw7Qf/HUjSbqNcV6tvUJXXa77wL5PZelSecnudjKp6amMmlzYvhLfedL2
4GdStUOQj97a8uWblv2FBzVbJMckbRzDPOwrj3Kyhn6EvVwNHkUqi3y5zu9j+8Ch
rkvfrzQnr2KURW7FNSU2sjeYhuYgGKw560I6avo7Ktd4YUundhHzqCH0djYMuCHa
r7u2exS3f14EBfah5Zg36SrnGiri8n9Hf+pTA9pAL+ms3GxOjHIb/x6Ia7tJnZIs
cwKkcNxZ/ApGlyBm5CNLBiRQfaplWiPm44DU3C5kqehTutH5Xef+vxEO57/rfX9h
/l6lpk6ymkxdJ0xZrExS8liaG6eGjmSON1JwR/Qy22TP8ndsQSSyAHKonV1xiukz
Bgu3tTwl5m8tJ0X5pA/ZpTN+okMHQL8rCwZp0XCJhjeJJDmz6C0atvY+1nc0HGyp
od0w/P98dZKp8BUm1gId/oQQfsbfT8zh2MOx+S34C5bi9AnovESMlyWdwk6Ybnnr
36GBaEkD+h9wRCV+Fi3fgq1PZ4og832Y8xP4S0BCA4PbapAVmFqI5qyFUQvSMhnF
ZSwrlGQbaRb27+XI+82KkGZZ+sx99kK+ffAeW3EIOLPuv/6neSKolo55VnAqJdq/
k5fxP717xXRabIPe8a+ZPjlVjmiaJ224/AoUPmFEu4F0uoIp33McEfRHmco0WK58
wojQ+sQci2jL+Ya/y7aCa36qaOHDn+p0ZjNZAqKQ4huSdacbPVFsYCCuKztmiMBV
2erJnkNKQt3OPU2smXKiJChmJ6Q8lt3Tka32xH0h5K2KJItV4LX+gRZCcllHV0Ge
vQ8Z39UEBZCfd0O+B2uhI7UIl8s71wYHbHULJC4Ren8jcOfkHMonuhZ3cbE2Tnek
S7jBnASgcDUrJMCX5jHxr0VYgAUCrizvWXbmsOf4gfkjd4wVgn1eK7lCru2wLOTq
wtGvq0ca1aRLn7Vo1PyIHgpOCLAl/1MayIRbno8iVgG9Z4kQsdMjq2vD9vGhGNFm
1Faut0YL8uvi/AjQ4PLyuV0n+xRk6lMK7kFxVdDKc23NQr2Uz4lXXynrETZGDn4i
ikh5RET7lxMB3yfZMu0h/lNU2yfXxp0vsNTQFGeQnaVsmxHh46qzUL3qfNx8XHsq
qbX0i9YnBXqSRT4elh3DliSPu4lPh+80YnNC3v7EfO/D3z33NyYAGoog8EvQEZ0g
atWscfqeStF3o9i8aXrLqw6yweB+0+pXIAOaHVPwSBuJ0gWY3w020hDi9ZQ37fb3
lqN3BJrOkmJhLVFaumMQMySS9wbtfUQNAUC1jGRT1/ybg21CbYNV+2W8zXIVlZlt
V9Xe+uFpqRgmL1VEFu9Doef6OMzCvWcr0UXPsFspFygphEGcWofq5vhlePhxG0Hn
QgXBcgtCnDssI3qAg9b0e5P/8KI1y1N053FUj7hf5ofaMMFLcO8WK63Den6jz9Ia
oVZrfo6K5jzzRtQ9SVcYj3eyl7sv0YHV+KidBUPobyGln9u0YPy4Mo3iA8xtUqMD
dOaWgzViK8nmEwp0THZiyr5dd3UsTXxq2mDXSo4x6GaoqQaNluPake/tDHx3PdFx
aueRcDDug0lHqkie3rDP73UQeygdjnVE9ZDorGq+saUI57Ork6CjEKzmW+P/ThVi
n2e4y5LNiT7CygRwfkxyfNoInXMp5XqIkK1tnzW1Npl5X6r7yrU+yViTsRIpZdv/
FPL2C2L/NcKDUVBCtOUa7cQFCJ0rUKlPzxQvG3P5KQX1YHnTaKxhM/ZEElOv8Z//
RFmEsf75iqm/W3ajVHEAC0WdsAsa8C5XoLg1Fh3/viQBo9/K80kO9TJTmzbvKv6V
vqxzkomzSqCyctwZXUepNl6Xfb0xWeblM+u0yo/FWemUQz31bekwOMQLUSlhvP8D
hCP6BEELTG46IFo7aaFRqzrGb2EdKeSnAykJpyzl0wmXT9aYO4ta8y7JuTvBgogk
Hgw8Q9wsd1REFOVjRD4dBHONG6LzqrCkRbRewXXkKDHLRm+tIq0mx0/ZzcivDIbT
jnpNMVQbU3GhwmRozZJopo2IQ5lMfH9/PN7oU157E60RzwPOU+OdQf9X9MH6CCw+
36nr2KTvLO7ykc2dwIvvBfgA1/yw5frV5Bq4ZU3Pr/QF1+M8qbHr4oj3Z5G6cEB4
rhcPiyOKR25GoInL1c8qJnzdNmHL6qDBCu87FB+135WFxDeUJQGMmx/iSkN2pGkp
lMOXYu6jRGSLWnjIBvWN6R33eK1i6apP8NogOX+tF6cSewAgY9ZeiN8WyzR1DdT0
cbn1LrFaPZEul7+k1n8I5wLllESIeVAApAKx3CRAcxPeaYkAILgIDpN0X+twu2FW
An5sG4TyJOvCEduQ5YwQi6b+QqmcfDeFwyJ0WDvAWw6AjBrai4u8YcMmc4lCX4uV
OgQS9cNjLiTiVFrnOswCjMG29j3KrfebkI6nPRItoruncSWyiHmuv3XuvgyqoOqG
c8T28e86Y0cDWojNSOjwV2/Ylpdd3bem9O9WTGRLwY8lOkSmAF3RLdzGkvXrbg1m
689kQJpM3v3UeG9F/BvOKu+OQWXxphz6C7szNpBlzUKjL1R6Q6yVM0LAvd8wwRuN
Qy4WkOhkOtgSXx+LJeprCOBEJ9nELIpg67LOHGleZ3LVu1Cei//UYXdh43qrClah
x7PMqbwIDOu4R//s9jQrOy59wXyapK5i2Pdl9Fnpg6WKw334kzb5uOgTvRRavD9B
FlTnV/wBVCWxMHmKKScQaM2iobg2r9aFhQbztmbY+3UVAmWnfGCS5vNuSeGSPgcC
JR6itVjBsN/J5AirqeCWPzMqv9V3VPOYEBYzls6tJYRguf7Pqyy63dLUY1EYWVDc
e5iF1HpzIu0WjP5PJPzbbcuMLhY6X3vk6/MLvTC1cvlw/3NVmeCX/L8I+ytzMNkB
RJgMqbB/PRKrZF4WNVikUmSNTcOMN2ghb1UaLcIj/+GTjfLTyIHqK3hdi/grGCdP
z4OqwYqZVHBhkXcveKv9cRyC5ChlkluEGYio0Irwj+oXbw4Ye3F40qy+Hgsi1jze
gdBeWHzQPPQhGTV6/j1uT7/S4iPE8rzVoE68f6e1Mjjk9F8LpVrR1dGIXQCWIuOG
84IeBgNlWjodnw1s4wdJGtzfWUi2B34ZNucFh2zoDrrZc8GZDhds06hnfI8LvucN
UqMqZXnZ157t91Tf1hosDhAAG+cBPjWCZcEzd3IarW9x9zT+FWZHAis9EOFdsPkL
jv57bPp5pWlswzVbh4VsHQj0iZhBl8gSlvpvjhgFWhOmxpxcNAXK7V0hCbo3gNQf
ShOLhPz4oVoF85BF/72unmWzSbDHTg4tZzzUAdpvizIpLdqc7tjdgSvFfn3PlDMw
/UNqOJwLtqgvBNeec9cYqgejqbAnNEoqWNqsF2O2z9LAY2nZkqjnVC3gZVxZQdDG
+jnpP1D5gbGz1Az80ntJwZsHWtr8fadofFaNTI3UtFc7w4057zR8Dk8BYVEuMC1D
5n8LTURjCHx8TXp5tuZz4C7cavonId+8pcCkflhq8YzwLu2XHA4JJ7zBsP9pBbCq
ekWLnJRL+ak6a1/z7GcVJQZmk6TiOkbqicstcAW/4Q/jBAfPq0QYoNipqeRZHhtW
ScOVc7mFt+LgcOzA/gPrt5u3jlu1fP25zGcJ9M7q+MINvtMSKxGj9cAgAkxTak1P
jooV5mE/WyjVJ0UlwqmtLOwhXSyubHs1o2znGvoAqc61Ru5nErPCovQnqQ3WvOsT
pej/w1nRGjSuaB3BlmVxczy3uMlyVW/vRTf4O2K7eNhcyh0hlr8uzqJeyunteGpo
PVPRQusVXJGMbJnu25G1AqvUdsscUZHNlnqRKMBj1ytsLlNTgElmLQqjQUHfjOdw
BENzk5Fo8L8Ne+dUPNR8IFD3h5tW+QNIFNRRdzdCP2JPjEsJlpc95ynxVgwwluc+
ieCM1+qmm6YIj903Sx/VxJ22FDgB9/xwryw9XDaEwQUwwtCkZAkP5XmNb8aue81z
jrclxvq4sj3n8BfvB8yPFHZ35qrQxBRurcz5rfsiOKR1iFKQPSZuZtpHrregEl9r
S3wP3sZfKdZQYE3uKtRtENwNJ1FsxzPsTRbj8UYuQyQ5pQ1xsZzfl103pXsO8pC3
MPYnB+OesRN2uGa61gvovi+hFZtjbbURZsOlQu3NuCkhYpD98iZQ+IAWn/dMhmss
adGjcucSBJO4TN9wuRuWAuzyf0Iom4D1OXn2p82rDTjkt7rdgT7wG0k4ufhjSO22
aFom34UsXNT8pN8QJ55Xx7ZmkZaiUk04L8MTB9dUy3Vc9XYt/JSxtui8bNCZemMo
s2S6Ua1S/l7nKUXVVFiuDKquRtkXrVFih1kjgezo7EcPxqkxc5U5OhZYOHCM3iyu
1Pb1JO/WR36SeEiK4NYPM+ORiD44TO77RtsJKILIw7CxiJ+36J6mcZpx1gyQBddQ
T20HwUa3uTFWIrv5LDNDjep2U0YNdROeX6dg69qYtcP3X0WuX59RbsTYp+URCo8y
va0yUClKnSSTXXypKRfO27pf+58HKUZsQ5XwaROHmycYs0QdlMqhm+tHPkfIbsVS
wJJ3LNLsKftAv5/Z9a8qvxXiE1xlLml+2UOMpULZt7Ik7LA5Jfy0Ytlxy2aKCzAv
y2QI8CrxYGe7rWE2i3riOfAKwf025tYZY56a1BuYLYoRk19cWuHvEtPYhYhxxFI5
7Tgno/Isj2TIpiry4vDFRJwkA44RnklJsbXKILarLuJsAN0fEa+YpScqtvrmwFV1
nDxT91UN2kEkp/Yvx44EIm53prg2vBdq5/rU2rz5yyEYaoVMrKPGwDo21oEbNT2M
dwYHvnQzsYU7ziegZWVa1x084CrZmwSfxKe5eJHfBIZ4SMYxJMizzIBp+bSRYfVS
PxaK9bHyC8hyu88WCwU357XpATEKwVBfsWTwMWsYJlu8XvOTA7mOY6cnrR4bsWgo
Pw+EW9dexc3KWus94p/zuFi65n6cDSw1IZVxxbw0NPa0N+pLWDBiFWjUzKtaa020
D7FOqqTui5Ee0ynUbe+QhC064NyfV1zArPkNniTQjR7ownN061Du8mNwuz3fZ2zg
ECWtwu+yHsXInUZFsDTniKJTUK5Jwo0W9BYhvr0I0PNaX2zHVMogxLfQuQM5RTzH
cMTuWCHGRd0g4dApS4m6LeXjx6kFnEKhkPQrWKvzffxJGVoRcVheoeqXK7YOc5qE
hKK7w15O9mDUJQkshboguW9WGAzu8ykrx9YwIIKFloJbLleu0OSU/gNEAf3JsKB8
QDTL59IhO4gxqehGiSFjcxJMlR09MTvE+cg+PF4S+DMcIa+Pj32lpJw295rDdZSG
5qYaKbMjDzwdOaVpxJTQMJnWc+NWtic/qhfWL+kVnWiE0Swiu9jVL8pwx9nfss9Q
VP29W4qnuvYxZaswOb6KCy5m8KLvgGKczxBqXGhJiPpYWGh5aw0jnTBpmheUINBI
qgBDJLdni3z03/6zcxcmXjNOhQk5x8V1eMyLgxifCNnEk2sqMLu4lT900mTdOtTJ
z1fDpyLJXteghKGsI6LFSINEHGCiZm42rjvUqChxf/mol/UJ7CbT3f9W4xDq/KsF
MPZcp96c1WalgzzneYr431S/9okY8Cdwq4dJeC/k+t0DfxY8Pdd3ZBiR/rgUsW+k
olDP6kHTiL+Z5+Zh40l4BIN2yup4oTxAyL3opBvOQ68CEAjac4k51d6y/zFWch0c
L7mWUyf46pZH0b/nI0ATgXyG3a+OBxKffddHLc4NOvFrQNCAPlC+6rIOszax34XC
ck5iLYBZ4WdmANSdTvGX6ndpfil+MuoTHjMpAd6BAnqjfoRB72OTL6tkl+/PCYw9
vHmRH0TkCareV/JGJ9VMSDh8sagPGOBqY4XTvD6FuiEo2IpdBobEG8Gd4e2x0cEW
S3apbEBmGTj2I6+ePw/EQdVPQlVTLGjetvCs67KaxG2V57lo+UH1g1vsCAVCkmMf
r6+bn7+iMFUoAW6zQbQjaYua7fM1MGc8ERPW5c4QfwRxOO/VZy8z6zGprc9t7Lca
dmzfozrzb6q0i8Xjs5sluLm2gXix+nj5MerO/aH3gRTk9oTEKAPBWuAHgzyRVQ7N
6B4TE6Vvec/DTlV9GimmQBoZz5q5n8Oum88Lmh8ZdVZ+dXttnm8Or0dYDCNpZkdM
v5HKE1m+CsP8hiaBy5muBD1s9GvJa2/tsl9oH5Ezp37M6r5Q849OTJ8U0P3caCmh
+S2p8LdJNARd2bJlZaGEaUuVYcwxExq6ZmNAdtTLRk4rOFYcz1v2NevxLmXApRlf
lifgGW6Q+OsWz496qU+jpVn97Fogh9hTOGigl867WkSd6LUzoSbPG8fw92Rl++fB
GVG7RfqZtbduRsmtb+5gSHl54A5aqPGnKjKBZIKI4/05CVKt1YtgjhBwTjv3BLj6
+X9Ro/Nsia+cOfCoMzP8i3/vTy9v9lBO1t1fOs7M1Cl83AOtzbc9+/i2oHLVCIH1
6Mx0BmlihUTbRg8c1SSH4zGxpoLA9Epep4W4FtMaxcFPxrnDKup4DZoVqgfMHRh1
MJMa6mYlGSeWGtlojyE1wE1CoR57UngisG4Y0P5J0npOCkPUPGIDfZrr7755SRsD
+pTqa3keAzvJC341liC1daBUQaBDdlSuityIvEjDm3nQLJ8nqH2fjXhwHGKL5BpV
oe6rz11tCI4TNTw+P9Mn4bejsoz/wYzziI2fWcrMpBWXQhAsHBdBYSOiAE9+oV+h
8qXsnPVRK4NuHG778qtiH7aiJNGT6AZoGozq49QvxByRUrmfixO9PwePMrDaRk3z
ZMR0r51y8Z0m/HL4cJWtY4OdPvUsXTiGyzEyiCvFEfTKZ8QVcYt5yB8c8cWsmvFl
YCWsYcv9Yn99qnep1GWNvMI+kKlndncm7f8dB7mz7fIRdVNtCViOSv+gr47FMW5i
98eVCMXvruIlwJXRrOKg4bPCGFl9t53cKHSmrRiVJFvf02znfWEy5lqv7FH59oiz
VzfDt9XxHdS6nPVFuUMwRWrlloqnQsJPk3AFI77aCJ7SwE1HJl1VgNhbTX0sALoT
/gSYdSkCv9wILfH/RkYKrWOlgQERNyl8k7NFNBupTaVYJ/kZlx3FLBm0gLBLY8rA
30wrz8VFwblhtEBw40VKqjfFUFp3ItTjwCZA2zUa3bO5XA05ylHCqG8Rh3iuI2wA
s5NPato/J8xdKU1/HX3CUwk5/eXL06/4LoH0n7TgNCxeLNiBdC501C9tcWwQV4Pu
w6i0hHv+WDvH7SbIQsX0nv0WozDRpMG6groNwJ262ELzTBK9LVQ/4mpH9+grQAEv
9FfbVVzV+H04PJeoX06OEzBAhv3m/BYuTIi5T2CSV+Oo2eTJGvUSFQutL5ghnypD
NMB+OS4MgtrIbefqaCOnRYJEMwm8uJQAU/TunafuM0WW4q3GGK8vys35F5dVVh9O
Vb3pl0iunnXN/JnBJ8qHDlaekSBdtAwVBc7wTqA8RcEed+oR7pgvLU8jR4iVX/SC
8vgwxBQo4KPCQICj9lb/t+dtofM3Gvdaz9C1gVVQ4BHGwhpg1OvxAOJ1wU7Ob8Tj
l2bWzqeoc79tqfkO/j8+YCZ579zb5Z4JQsjLpBjyaZb83/4DY6GB0Gk4kxtgdJ63
1Qwut0QN0fHcNe3X0OXWIhpuzfgj+e2CAETYq320bC+aAqCjnYP9miSmFpD7Llu6
s3zsyYN/WMSjc9Hb2/+ErBgWVT44n09hpPdB9V+gKe4J+LolSna+C1N9PVMJqrP1
7Qc1e0J9OEsbxTN08UVGVkp+rvGCTGFagGRMVarTuyeaE2Meq7DzB8cFSAlJjOVK
xLsESbZ9SgRiTAgJ0xcfXRksLj2SMgWoB9zcJgbQ7+fdawoHDSDWbozueBX3A8x+
qPu1MFIF5q/8EwJvaVc5lh3bzFRsQMjaTVo+G2jHb1H0UrMYpTzRYawzK9R+6M8B
81qkQmmwBt7RgNbpOa4+2mPoG3U4JXr6jdBfOkwCk/6+AFbIz8q0lgr2gwpSY4mp
yYPyrag6b4a0iQ0H131URyx+Zp3hGZn6IO0pjnaGmR9hCeapX8baSCG1+soJBfLv
1NwI5adjNLJcPhfhk0Tl8uiliDfMdqp5pzs8iWeMmdiZ/ZoZgZjCk+Wl9xi7mHaA
r8ypTuWBPVkO5g4aAUH6H+ipBtEfc/rcuqr/6IPzYiPoSPFw4rZSkYwDm6fht/qg
ef4tJiCkpdVC5EHStv7d8KVlxam6CutCc0606kGS0oXw603jvdxesVkChfBg+cGE
pZGOXni8hSjFZy0eKU6q5pWVSPPBmuxkQH+JucB/u6CIMml7fpg/HD/KnsEy1Na3
c2jZxy9PKQu9pJXjHhnZvXxaB4Sm/49vHBlyBdNWG3ntvq0u5mrFNrFoUYNAFXEk
5FgHzFC76ded5DSMZ7i1SsZJ+b/Cb03H5sHN4cH19XXKP4M6qTFux+3P9bs2mGi3
GuXWQQOqRGDeN/aEfKfO4dzorQjB7zf/WgdLJFo3/32oXWMXkd9HQKFnVW4OT4UW
oA0e1TDih+RlLNRQS8XKfn1JaMaL2v52fNu0o6LRFNzxQ0IBSvCpdvV5BUPoH3EZ
IGzuVhvWJrIGjzb3NCguxzoiHokpPbg+QLN+ghfADBp5BULL3scOV4bnjOsfzH01
Tt2ASI/pmfFMzFV489WYTbndiT0EltgjrGNZKEGgy2NntHONOsKgy5q0YSSxRIIp
TGoBGZfEji9bxILfCiHLHk9da8XyPurqkD/uD2yDOc3E/3zfSPzXz7Wuga1gppDo
6Bx6ZwEbjucoguhELykJD+y2cGB7YzNprZRhPUAXbOXylJ+GE4siC4SYDJUiU8sx
NeCCY/BfJvybbC5S9MPBGQ7TPbhJS70bsuvRcagTseuK6NkYK1z41tqr1CH8C8c+
ggdkNW64hWTv4acZ/IIO9IMl4CYG8uJCJz6QN4hSWq5aIe5VqK7lvdgcOuvfdhF3
YLpK5R/3AyafV2QxlmmQ8YTy1QhKi4Q8cCbgrvWPY4KxQ2DAKQiB9x67eI3aenuO
OHtX4Z2tYmDWdW1rvLwmqogOHFy04IVRCbI0DkbOznqX7wIlSSK03LomezkgAfTm
Ahs7v5ZwdcN+PouyECWQd4uAfvl28Wj+rShGW4VRaOHYd02LeY2gNodR8rk+vsAB
LAMrd09ZV74UGurdUvawynDAMTKlXTt0HgLxt1IU/5tsymAyFqkomjG21ChLJwX6
GG9isf/8MFRU6oEqkiimoRb8BJwHUef/Dturwa8hx9fPxG9bChCVQsIofl9SX8z0
xvQ3gPL1LPKcJvtKxznif6DIunwdZ4ckst0g1dSeK16Ku/+Xo7boOdIMayk28ksz
DZFE+w+QY+emyu4sGvJaK7rIL+LMge22mxWj6/h63CVrzRj6On+fI2TxyXn8a9wT
SDoh28Bc0FDL843ADj/BpWSw1HdSK46R5N67zNxzQ+rwbKBGkxq2ikWv4V0GjnuW
4Y7g1ufv03Gtd0VxCeNVyW3WK8S6TnekXVRS95AyS7kwsno+hoGlN4pVUEG4csVa
1qJr1wpnvo5MOMxVROn7AAQzSOhzBXF8YsKv+PQPKGHF94vvl0nuMetpjlHL/1S1
85+Ir8gnQAi6nIzjMCjsMwT1ui/YbXfxG8CeVFosHBSDVXfpK31xl4a2Shp7EIqD
5p/HJPujHrhj5WKM1FuBqcUaKtpkJU1eiuhMJP/NhDYzHDL+9BUTgvdOKmYcecrF
yKvPJ7jiWIU9D3sDarF9jnHInCKkbPc3rQ4y9tskarerql5WHQAtKdtobgHzDtcc
MK3IXz7CKjazeVsL3bpTF0aRzGYrMWKgLBU20AqfVxlCvNSGy0Pdf2DWBZQJxPtq
bF7h4n3uXtWkIYOH/tXrml9F89lYzTNjqJ1MHxqHGtXTwVofG47KEurw5fePB51e
8wDpaxLadpbrrEH0KnhWbcZGBG35awi5R1VUhhczCqYgMWxONonONWwVDh6jA0tL
jktvDrs/IDfzMNVFMijwYuuZyWx/bJKGhb2zrcXxULbyCr2uY+G2U2GKbDFe9m38
U3YZNpeeuzyQ29tNCsw5MYrIiqIGX1JBENPWbFWXSsqd/3RZDNFzOJHpdJ/mRJi8
mTU3y5CN6ZPnU3TNyjOqeh25Gl5G4CdCJ54c7RAnKb7Gzj9bVO8t0emQlwLNOWss
nsI+i7ymDYD424fQroeXPXhfgEsLP57Nc3Whoebnj6jCE2gM8dTmr1+gvoYr8oMK
WJ3lij1Q2+pgM8p6x4Uhf9Ubjd+USvarVIhqeLgySNBkAGPx8wGSAFWgA/wrDLCh
p7UJWv58FzchrM9Kk2syQPWa8Qf870eSoeZrzUXkCHf3qBDeZRc+L225Tc4EJY8+
yuDlJLA+7ko27AhgJEyM1GgD1tlBgmaAaZQpAHFvXOMa5ZugCXUqvJIPyrZHKftr
7EVco5ayy7edlVL+VZzXdXG7v8t7c45iST2dco/U1S12Tb618thGYLrjlFVjgtq0
Mv7oUX0vC4G7k4NvQEZEbiYWXE393waY5rL5DlsIVGCtUd0+GBXowP3Wr5ovL1FF
PUmWsdzrREsB4cruswD7YrustuqKOe4aJIidicF1dwK3l6VqVeSj9BiikGOckqrn
NKGmxMiHmQDiZju6CiwYKnHYaw/C39W/v6eNvbSctxSDXzwU6DGEC8Y2T3KDGBWD
YWx3Wu+DRvf2Ofd5MQ3XcmkP70FSZpxpVnX/H6g1Jht7ipiu0GQKcMrF/KwEta1W
2K2a7OaRcUVpGBSf8JkntCHz+ijmfBvPfeBviGR1ewwHWSUa2/MK9LRsIWNFoQ6K
uhvkfLjSYidL0j/dDYqWDq1UND3zy45xYzbBLjZK2Ex+2ir8Hal+3CdB4itcWhEj
Nqqlgc1YoshpU1jkZXPrfka1sAiG+uAVUhbQGI25XwMGHtnvz8/aYBjY30I5zp3n
YVyGAF2IJkU/Y8N6iS3Hd8mIqOkquaxxQnxazuS/UFaGQFbykfEqxZdcvgwBHTmQ
m0YC++0RP2bu7nQkRQVN89+eb8tTueZYPy3CI4L6FkvE6Vb4TsUyscxwj4CNVQdn
uo/9t7pfh5x4eBVXA1nlCL9zDgZDOe4DmZxeBKcUrA5bx7KwMldbtiBvHlwzyD4G
pDdHGkBfPYCtUZNuRxW2Rpf0pZvDVViVUHL3ghTRuJy45rmMWIhmfcQqQn1P9JLR
i/JsDtp6/LWzU4EzcecDAWBHtf1WsrWIHG70B8miXV1TuRMFZ2SEDwkqzU1A5R7G
KVeRkGEqCFRdIh7tb5wopbTU7xaJEHSwpwras4bqwEYLiHD3g0q/yZZD18u6dyOt
dV+OwXk7N55dLZzOJzlFLjdSV1RwmMnkvuoU2Rl2AxA18+AY6Epe/ewTTykbiSFl
BOZzf4xNKfP7tKMCIiCj6Cc+ZaaMEqNr55pBrNkt0nG9aCksD1O6cDf1jinwynGw
ivOudGRNvTLRFH/8F1g/2svkPTIvARD4bOAxcEqB5zTWTr7R/5vuvkMlj18HCpBB
BCmA1Uv+y6VGCi6Yk2uSjtwiq/+8PMj07KSK7NXFpMXVrWa9VsdRHRmcW+q5al7Q
KBuv6cf1dOulXiKvo9fuhlw0GwsL6wMO3hm66ELNYzNAUusNpoktwqJgKGBmwAYz
Utx9FcLpr3pJIsBYLRoigkMw/N70WvFVA+rGL8T2/65nwC6HEn1ybRWFlCd2b55d
1a2I5i43YojYDVmJMZGfLJ40oQyucM4lfqUJA7hqIHfWQR/5L/z0F1dr8+d8DreV
mWbtwf9Ua5FMqujKVp469eJDa4xMJFiHB2LZhgu/wS2m7211Le6u+/yKT3vHBlK3
h8i100N/D/O45oKB38NNB0XyWJlEYJ1f+Nxzu5Z0FnbrT38BXnY7pnLlxzQYV+OU
v6HX9O69ON4XioK1a+RpgHELA9lOc8s5cuBlCM7p7H7BsMTDWBgn1G4IJszLCWS5
nLKehCFlLETBnsL1HzxGGKY9M/zv/CoQBwb64SdvHie+rZ2hlOLQoIuCtHwwcLow
zOAelKeXylsJClsxUT1vGKzGn4Z5tVyZtKoxeJfnw903YWWVxiQuRjPYqqrUoUWT
/u8T/BmrfG3J0jE2iz6H/Vy9Tb4LklEMcp2S8CgNBNsF6iyY+vKSrc+iQ28VkMOB
VWTDNyu/NRJHLB+lUC7tYPxq4KYz68IZCjhGbDhZOqlBxWDogdazrUEN3j7NYsQk
mZmRe0J2clF1cAgpFeWiiSmIkfxzEQNyVctAUO51f+1ktZrJfW6Qzll0WLvsm3Ud
RSvFzSRGMM+UQ6IcTv/JNbfkpn8l3WsJTCSLdwNGPvGl97sbfJFPmr3YOZlUQflM
+PZ9pRCL1l3K4vbNGmXIHlCRGsPW8JFvuMvDn9dNTgrcpAI6fJ5GP6uZICU9LPI/
Z8M5nCAw1JMDF8tIQgv+hDNT1oUhVye3LemIyF41b0nMwvePQjLWzFRkFEeT0NW7
+Gg+aEKDD89HAJhb3GFjjWZGRIlTW4bkUB4iTCchTI2GARmSVmcGMr2OJdQPkoq4
05WZ9lTGpKDmh8v3yHYfSMT8a1ie2oUV0cHFbiCTpo8qsvwMX8FvFH8PtdrdVfj4
bvGnvqzS2v3ulKRD9fxkcTZa0bkj8Fwqid46O3ItwBcRp5GmVGSBybBckc/ALtwE
FJg6mT2Fys6gd7LkIa4qbHUBzgPUT1Z+I6yLLbR2PHlF2c92wfNUq9W5ktesrtK/
KIA1pyKH97oYPZyrENLbWXq4s2tdzKX9icMPrWawoixK0mFundBRsoWIfieWpraJ
9De/MRLglWCWmMK78P69S+wZQCep33QaVt8LRpv2vyrufxUUevrm2v4N31/wx1+k
DW4NTU0GDGEQcbvAmqDT+LQGxYzK13DS/0xP6KM7ognWtYURzZ1wzFUdeLFYemn7
Kj+k1Fk8SuyLUlNd6CLGd566T0hYodMQtppCLf7Sa3MkuQHudExykSm8kRJVz9df
noSTJsnAX3mAiCGsDyOc4lAUiw1VErC0fKt6QDnq4XVAPnScJR+ntEkWO/FJKBxR
+ShVBMh/WHX5X2aDhJtTY6mv8Ybk72ZFwfcQGqSh/4rqqVzQ4+iiQeN/xB2EjQNW
RBtqMOmp0YTbeRFVx1i1rIcrGPMg6rU848hydwBAe8nwvgVOjBEks9e2JTCh2CRv
Rsg9jKgwj8YbGxDrS2hu4GiczRuuf6Juxkjr2ioDB2TOXko17Gg1Uml7yJKQspk+
AYkQ4FuiVJKTv1dvRLTKC4HAcyW4mFQJR6Jnpwatw0Q1R8bCSSMIwkpZS5y7SUGO
NPeavv51CzXR7bR+AOId5nOIWDlzOvp5x+7MS0wr0PgWNB6+3qAYKaC8wzTUz6em
kq6AV/DkjYg3mrgmBVQ5NGKJTIdU+ijNR0oRC8C4W8Rz9AqmIK00/Nzf9ehKnZCS
ZhUjqiiYDG1I8q23Fwurkm9XswpIPvrZIsDiKcgxXG/gvvYajGyMH3Qj5Lrs8iUR
zYY6OGkbjvhG6F1z5ZtpR22yMl4OuHeSaYpAs4hMa9AJ/8j50EVi+YHh5s8fHODZ
cFsbHuruezWKqa3wfTQcnB/pT1PLRcvEOag/7O4ZWp54laXrrIcY3emRgV9zfNoL
fafCGzKfQpcuVqSrxmrT90Og1Y3RwkaO4sNXUEVQaXgwWauCIacrXLaGzhbGSAe3
03z4VEzalxGanG0lC6dDz7Qaz8SMDK7zJccczU7HqxtdaMmXSTfRPJk0PXLEELcC
TamHha7xb37Oyi4ZxUpuF9JCT2FX8nP/ZkEFffxtBdon/uWePW24CXdMHkEEntUF
PZfnbXfm4w94qvrnD/wTWhmXn3Q6ak7w0kxScpb+XvPww1v+vIaob3/SPg5r0Zcr
wLt1mNo1ObNyx3v6Ejl/ysQwKHLf9kp1sRsACKTJ8OhC/kIgpFFOcqIaY2hsdUSB
0JeNoNFSh9mDSGonVmfsKYxAvaE/Oglv0KpJ9FZd5KAEsljxza6pQggkYhHqcBno
APWXtqHKyl2JhyPfxS6tmerngoC2XODNNuSflS3bIBWu4OPZN0EFWLXEUlPOsZMU
go5CEMOBdUXQO+470h0zZPh3LF3gzsU2pjDHUS4DCRfGvCNwTr5gEG30Q0wfsHmC
HA7x/66fMTdhKylY2lBkPDIWkC/SfpOIAyQMztXVe3SBUKEYf/c8oI4P/DbMePyw
jn7s48+2SJNdkl+iOhsRv5oU9ED/7WdnQJT9gMbQyxqcMiZ2D6ixEVhey04fpsNn
FOUBXNMu8Gugu1Q3wcWPrcT28ZCGJT8Sbzyi8MmLgQPYfRlXyQrDl5Cs4ehnDzuX
3VwP0hwdb3XAsoR1iuNGHbVnYbniR1mwbFOMBIwvblTAnxfBl80911cVEG6Vy6jt
5H0y6X9hFbptx7z0bnNC+WvrXL4AYmXfFApKrrgLPXBNb/0axPOdZ83sm1RQRIQJ
ZMBPmVa6IbtQwbnCulhm1E9wQPnBD0Xz40+PQq1VuJnzw+Qy4IaB/9TRg+GTkQPY
ObpU7KYTgMNHZ8i1/VHVO6mdNOkOk1nBidTAZ9QVWbXQbkKRaC0xzCFGZXK80v9i
Ma7qxW5j7rS3tmm3TL8agjG6oVT/ZwsNHtQJJijC84NtBSJSD6IXELpkQybQ/pQJ
hN7DH2HCpT8bN/0LmLHRf1Nz5vbnw7ktoURTFtMm5Gkm54rmkc0OK0WwvJbbKR4V
iLWlQ7bR8gQ9K7SnoWXbtEAUFBsyXAoxHDhqa9tn87l9Ga+Ho7Tpg7kfMtWKFgHE
4Wutr4hnw6Cz7ZJGKYRcdd80gSJJGUeqMQaWIa91GkAOnboVNfMnYwPxN6CxryA6
JVcWhRPQTm2zRfy3M+oPhG1oyrNl1GuiCS0z9IKPdofYXwvBAia2tOPz6dAyMeC2
dUedgwD1eAL5zA/WDhwTGhPpAvtUBNVpMOa+BF/wIwG9+nm5Q7tsxXp//wq5rRi/
Egu5HKtFluG6GbV6Uf5br/NWCdPVA7D5AUd3qw/mNZpB6keNatk/dv+AaeAya0LM
kjjUFnYAxEA4GcDsXBMl75jgMWIEM5WVXnVcthEpuZ3dO6bsqlAVnKga+0q5yVP9
mIQ8jQbIYBXQHxRCa64hMxYD0qW0aZPHELxvbknumDprMyFNjuIbNpfWhY8iuEu6
wkN6lHzMoYJmKfXCeGraEhUOw4l9GdwBCFZ1jV2gfeh2OGzGx+9gnGX11gNy73cy
0l4fLf5foDXVfW6KWcWKf0KWXDMQNBHzd3Q7v8lBZeA/Ct9+Eyx/njBYbyKyvtky
r0auQX8SMddZTI39pYth3LKufm1i4btA6dsY7gYeQ/Tlwc+LZlwRgm+xZiZWMk35
Qp/uYf+dl7DCZiDgpx/d02wE99yl0eFKcsx2afB+S7mkZyj5oyVrm4k0pL1F4f7o
J9m/OuHbNtNJ16uYEri7ezR1OCZF7wNDT4KOnJ3n3eHiANrM9zUI7wPwzcWKivO9
t9c+ap9Vx8uvbTHAtQ/Qy18D22eWTf0gKH7jeby1BXDJbNzUfyK605/ey6pgtcm3
j4HhrdHiqMwXh4Uukz5TX3EfeXimkRXXANumZnrw7MyjnDGppnFAnIxbsqNnIRHw
9UyQxP05dcI0r+tkzvs4N3Lvf09QfYSUotWt6P/pdvW4Aly3L08twOHSLbVXROYt
InNpkyABNBfOnbgIj2k4nRQziSqb/dywpIIc4roerQqkkTJwp/e2EnLzmE4MJRfK
kJgODhfKS7brhOL1X1rN9VImw7Jy631KtnQ6cLAT2awcg3Qvw87oeczKDLlb7/6U
MqvGSLzDkksuHTvBWCVEgfx0UulTZYra2CzIXZrGV5W5yU0sQkNqO1QO1Woetttp
Ibt73yFsexPkZoLGMZKbcBULSlQUxS3L5c3vLGzDQr1CcA1HECmna9QSKebwImNk
gPrwF8P8TJjqLJLzjyQTySau7uJPryVLzylhfpMtk5hGyak3zD/+wCt9/7eucr2a
qbSb8XzdIBgUPWGRILezBMVw6rjkFl2L8LclgW+1wpPgyr32CsVZzCJ0rdFd4v1M
p9pbbPE19L/JWgG9JYlHZTFupMRdlFaaefwSnYfLmJex0V0DjV8/BETqc472j/yu
NEoEV6G05YZkt1jI7ebRnvL8M8puvPLC37Kx/gfDIGymdXQyhh7OY8009Zb+izyi
bURdDcfBFlbMQPRPF8J8v/QBKqHTg2z7Bu2s9KhyzEVQN9hNlDnipYtZYKXQu5y3
+9D0qGz5iiYRsjHSCHvx0UeMQ/s+ajlD5mFH2hXVjB9V+5ElRInRk3GNSonXqkgw
SRqc+0vH47454fggebsOHshBZZwLY4UWR+ZtY/TJc/k38a9uqH4A3DffgdSf+qCX
lz6CrizduLf8ra1Giqxjaku5Df7RP8oso1hSfCjiz0CfZtg3MIKYD3bo1cvbN2pu
cv6/cqFDffTXqRTTOJJ6bfe9RpWi2axnF2N2qASbAKcvJtcOnQWbOaFAoP9Aoyvj
yZfKDpxCVXWYtilQ9Byb/Z04PcotqRCgUdx32bUIBAxwbulsChCixqqiSWuslYHV
6BVMaqhmP1KvV7NOdT6uym3OrDZf35wtZC4NG00pJcDun0DshxqGBDFQNsM0eJ38
wp1BirR6JorANyOmWxkJr3Oxa/g1Ru5diV+0RsoLKO3xfNwpws2eJ9HsuUEoxugT
eJ3MUhH1CFd/GyiAutF0WJa/FHjuHFXWnC9t+y4592bHyfk8m+JOdSjscMq6Htac
HGQ3K+meft8s5kRHu3t3CqKgYUSK2vZXueJfQkCXUw8uNqgvxWoewQ05xOmPJl0k
0gFFKZ92PMtErJduiMnf6B+kd7tpNfHTnLfW949dwErZR0ETeyJLVhjvvQeS22B2
uy41OCOc+7bPwbSsGaF1wFZ7+rSJXaqju+QaBxIA4hI253z4KDjCzT3HiQ1CzlD3
2pZfUafV+hkeFT/13H3zOlvivdIli8xRpYawyhHmUqA7Si7PQxF3VBQ/+MR1gOQZ
NkkSRPGQf63ge0xGGZNwp4/AE/Fd+S7ZtsGzJu0wCzq/H2UBJN3tWokJLqn6aYq3
exnBXl78fPukFnc6xdf2mm6uSzTCV4wvJ8B7ek8WCzIc9U+2Fawhawt/FG1zna3N
cZDAPinQu+W5x5MGe2aUTaBOAkss+XknU+ZJVAxSBHNIcKbbDNscGHpa0do6AXbM
BNJCy+nbzCNVI0AKmgM0NxjZVQ4cCmIbqZPsV239Hf8m98jOdhi+nSuw57Ctc/Ai
IfmaHl2PnIeIDxbn7D+THcEFRxtAtGglA4G+1yWPjcwowWmF7iGr1OAnjvcw+ebP
iHLoAHfYP7d0IJVLhGSgJJCSZW6kt/vFI8xkck00NCaSvFnXPNJqkbbOXjLaonze
IJfoMyf0G7PnK/NKsIisNjRgjsOuAXd3hl8Q9g7YOyZWPOMdXpXnmxz9oFy7wUzn
ZFz3xovW2o5u7PbnhAw3AXC7AvPB/5J3StI4b7LqijXSvqnrNBc088S/awzCd1Mg
N5VapTa5ElxHYK5W9oG6R/o0bWIRyJR/nVVPqKZTcdEyPixz03ehGyPVqtQQGZdj
P3AUyzj5x8FP8f+QoBaRikskxWpKJ4KDh+QeB/iK7LdxWXikEi3/8kA2pzrMhWYk
WvMlAQzvwZvCvl/2qItrlOgwX4IlinXvAkMG+1Iim7ZOIJFpvxbNB/60ABNt007s
C2coEv16f9dktUJBOFwiAZscJD7576JefK1TIQjkItZCmx+/xP3a+m3gHSEoyl47
pB8xg9TDDs8oVHi/zmf+5t5PluFEmLUAJYWcw13oeLlMv6MUmZNMAjbLCqjUX0tx
bTV2hzUsskjM/dAr55OyEfvISXHZt6ZL8iW7o9pft1XrWEBLA4C3i/9LeaLwnOOW
YqaBDZik6p8lGyggaAMj2stejQYnWryRLw8NQ4FkLugDIBk9dXww7RzyEY94Yx6S
PqknjSwqrjVykQEf9UvO1u/UhsXiJqHlOMMxa9rcVq5LYFT4VxSOIyvWWrhge9FB
i3RGq8Vp2F/wYxqLo560IiOf1kHNakIRUqo8ZAB3DN4d6It48zcDG49/vyrLdtdB
p+zdRfnk7d+9dzyrT60p1ZRqpQNVtpR6vjB586oA+SqcGhV3gF+T+Ns9tK11C18O
pU9ye8PzsXjsJXKrI+J3u4LYoTvT6HAyr8wxxHcVJEEq5iQzishCQXps8d45p1wP
BkBq26D4LFSTBeSaAk3o5Ymy2AgTuBCnFhbhkPKWrUULmwkIG1qNW2WY4NAALSO+
rbdMFvycRnSY1RG//GFM8u1Jz69/zNC2jA9gaSqeva6l8seCoT1dpKbawsJPbzCP
JTCWc8mfO2jcRfPMGCrVFPOn8aHA9147Hk+f5VLml3C+I8fktPpM5AH2cj1x1VkI
10tqW/YER3bKeUr3BfXiY/hJED1jeBhNWEzdnISQfPEPtmemT6rBraZp2B5y9JnP
a0UYNHDHpUGVh6katDuc4/zmNBOSwn384W/KL14i22RQmRPiAmiCSrMf2qveRrNu
Twzx8jqEgyRlUdqmsOTQUP23CsIPNksjSCni8OGLUyKn2w9N7BXJD6W+2gMzINgM
j2mZE8p8/zvbIgLZPN1OYtV4km/ogQl681UC4HBNtsm/0+rV598ztT2+n68hu6z7
9nsfG71OFfaZNWLijvn7iRBsa8IrYRERHCglUQlNDW8BVlged/7n72iokX3v6Hzu
R/1QcwqdxvguFUmAGYOEW0aE859wnPiILR1IDGQ2XxWdRF4VNtvYxSQNAO4NxsvN
Wq35sz7X/wE5ZtZGFr8l1wUZZx/Zdv2mYewO+me0O96wLZUFRnNAYHzeZ52MdZ+I
8901NnDcOXUiXxLyxVPzeekIW6s+2tgW7X/A1f8rBGdF4guoWyzLWNyka8TqnSph
c9sufK0PC9KWt/9OZ2sTs9FnaLPl2S5r2Ob/IahmF6sr1MCWqldPM3ntSNmclOeS
MTy9jF9dLVcYxak2UcAy9MzTWK0kvikKDC3vRw0f131gXx5sdF5iBl002sBSDE4g
zc5sQ921Ipk3EQWz8TFR0D84nwwXIMmqNwtXvdK+7bS48mOhi9ZRrO76xoB+KcNa
/vwDGQcnjkv6SSVZz7en4hm3HPTHmqSZF2imzv8BjRu2sbk/HlYhRRsQPAXmvTLv
uepSMsVKtJVzGfWWn9eEdX6AF2VS2o7j4PupRkHAsSPJCbgMYi4i7eHB28WldBi4
2CU2sqkkj4G7V++mDV1Szq5H5TJNrex6OGhKspmfVvvrSOmG09DMVwVYFr+R9EZd
5w4X38PqnnRmSqgE0ajxz2mPj/XBp55Huk/kKG3URftWAZbY3uQlOwYPTYKeRvQu
byP1PQczeDbhhSeBIy7vfu3WvNffh8ekYlUZ9OrHsFyCuSVj+cJPHb0CwY5X7Rpx
/lPMHurTMbbrr1Q5T4Dh3nJF8QmrZXMOFDoaqf320dfnOBvjCoIKTS5O2NkaxZCC
1YnGeSlu3WfymsXwSGd5EFhpPccPO8zBggwX4bRJNXw92C+W/RWXkzWWZrdypYD+
HIDklROI9hXJok+wtLPIx8EGzGq4LV/TaOZxCAQe//Uygv8/rnKYoadUpC0/FM+k
wTvIos+CoT+O4409cGMHJvT6YxxPmgDX4nx8A5eVwvwcrPxL5BE9Fy4rm7P3E3im
LC1xpcsNr/A22tE0CJnKyBLHYaEkPLL4wpG1cMIJlFmS6l+ilZiH9GzG1O73liG1
e/Aalad+3pDicG1UCUpB36Dsm3upfZHfTIjDWPT7OmmAXrxHEfbjpGR7JXbS69Gm
G2GVNJUJlI4aLSar+oP8Jsl7Sz+zJ+fT32J7RMqQ6c/fHM7P/ExL+U2UypfrySz+
DaLgUXKJrODXJuWvrYUflyOcwRelwDwHADraBKJOsTk4++DPq1ldoX18arapuWP5
+XdeIIuQAuOeqscgxzXUddN09Kj8swXLqUJVLfxcRS5X0GwJ0AgDvDxXk2MVLsM9
YEVvUW5AqxB4zoklhd/6H3/10pv6B1LpsaOnSm95KGghActNqzFc3Obz5NGGOH+X
CEM1gFWWJfhDss2tqMxjIRs5hvpZu0UkcX4Qc/Kv2BYFSGQA0MZdw2L+b7X+uUlX
xqSR8tE9VipV8bOchZJEULvnK9VwMfwD1aNTbV5CGG35JA8uVT/Ep/zViuDnjygi
W5WKT0ebBOrysxuKLI2rCEqB4UcIulQ+hJUQRXNEaytZrrN5Qf7nGkZp5SZzQoh5
2cZeLJoDiEOZpMe86mWdspcI8PnMvHrF/ENoHKcVwze3th7X1GUQHPIBMclJHwHR
q43VJFy4kKpvV9hxVs7dvwUluuGarz+6z1YZ/na+kTDoKiSpUBVhqw4JSv57bWPX
/8tN8U7E1D7eC2IZHGJTBjcaqA1j0xC8vjCSGfHjVm6PFyraFiYxvJGdT0MVyYl6
6V1+PEQLeHv0S0s2e/vVKLcBGPKFrdhARspcZCfnjsfnVlerXHInjildG3lPILbX
WW3BKMGvod4XH20dLA43dw8e8Kzbax4ZIQepdqNlCazSgQABBkpXm/cC2RHZjhCf
WbTdKXWljrYiwIBK9WZGh64rNTh7l7JLUO5pgYmvm8clSd3KZ50x9z0l+A2giAuv
en3C5y6mzONICxZDGDVUvQELx01UnCfCVThbDdGo7Utadya/kzGzTYO5pmCwrJJ3
uz8tLCo1oFcHJp9MEDC4hbnD8+kSoID5M3m0jHp9JTk5PYnOBnNOKlp5oI2lDtLg
Yhivj8g7XuX65H5Rdv0N7NxbsPg+J2sAudf9UdWBmzFs8XzIWKGRI4QAPxaVDh8F
/CT6KZOpEwg1nP6RKp+0j+zvSZ9VW/mbPiMAvXMK5/8dVE/u6Uj8zoZDk6s5tsRS
KQ0j0X9WUaedcUdkUMrRI7OJtg2avoGL3X0qHQylYMOfOK2yN/im6y5rl49aoUKW
CtKn/yhOJ+CHAxLvo+7rswA6Bm8oYFRejMSObV6nW9SoqL3m53i1HFlOqP2EwutP
azkWtday0xwHzJ5fAqMPpiOquCa7D0Hr6cgaC78ztoVMDkCC+2VnL35eeqJINusU
qDTB2TJE/E+LPvwaU9+FCdcCyNSYh2Gg2AU1Qb2Fm0hKqY4NKNjhA/pRIKqKKbc0
KfMJkI95RsHrn31KXbL96FHEj51Q16YWc5qdr5YWanyUMoh9EenvQqV1Dj92ZVsj
4RqiJ2l2mUkAx+1u1VkeuuzDuG8okvknOzZ5gZAy8vS++5YlE4JWGMp+h2eckvs+
rpAa/foG+7Ur336K5rKwUrbFVMrbByT3c/4ZlcnlO5nw+UUOpVZ0jYxA00vMyevH
IJO3S0hsOPjBxM1p3eAE9ki3g9oFcvAzJTCcb99wrhHa8tHWB+qJC7Fe5KStaqxE
nt7Rhh+dSPLM+b4ntMelTfdOVhpHV5caPPRLOKjjXCDJ6w70cADlCPau9sJbNSLu
VkqXqRFvlAbGrpK220rqfoOYWgqiX2/4SShJ6SGa2cWur9gA49p8bjzrvi6c249x
jHZ0hp71YFb1syFEbIcV54yjM6vfHvvXV4NjG/OsCl4lmqcxrYcVauDb1WfSceeW
aGgICWNjW2asRkohtpTRMM6BrXFPtKfAsx2IKm/DSAar7geUk1qdONEVlMa/Uyhl
aGwaHBFXKOB5RoMDMrChsuhTsVeZzjXEh6F62jixWbZYgRUY0hliODkGUXA+/3mI
C/rBYBpIz8zr0qBZAOUbCFpa2KIK3tRzzDeSzoqAZQqiuw6c806M4RZthRV97MQn
Xy/cYSD2FhJkMhVHzOWE3OB6c51ze8AZbMDZ/5iN1kPwxLeIALv5FX0vTDIkIb68
3mmDqgqMGj+wLsW+/K6PU9a5NYUj+Xa44an/mtoIDPp2EHXQ81wK/z8YUxSZj5mE
gFTScx1BPOBMl+h9SoObOrgW1ubZD6z6/lzxIPHAMv7BJWzEJitXsegdeQ9hC9mQ
dXy9jznoyKqqcOrefwQp6CsnqJezDTCPlb/xYWKRErYXkO281UecvTC7WCLpIWIR
1QraOd4ssh4EuhZuGTm9ehiXJ9afr4+fzWooEZT7P7vmBZK9UMes33PAqQzfUYii
2F3nUjU6A5NLGrizZ0OAUXmHGXAZj/Y6p7Elb9hq9fri3y6CcZ3P8ZTWPImSsJSt
Q/rvYZKoLYlhDXKOgX4KEFmm2hrGv2U7Wi3KJqoq6T0GBmRjWYCKCNFmuv6e0VY3
Ii65Fvnj9CuEP1rZA3hYvOLRAoNuv6kaA21mohihyGjAuppxqiC10qPZZHa7Bc61
B5/B6MmxDEj8nm+Ioe39Rszsz40tdLh5NyK37cCjgXU=
`protect END_PROTECTED
