`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5PU1VYALAQp12Pldmrlx11uv98IJUQNrTtbQGJ7p47a2v9Q3qwd/h9atnq1Sbbm
sIvSBx1E5qytUzR2mdGrbTtqqxdnqiFRoiPmm3FIIZX6hf7yk/nBhCWWdmS/+Jz2
sbgPO3u/0VFMMm4vUYThahSkxVGWSvF35lfhbkXFS1ZguRUVbvLn9GZaHVN6/+s2
sj1/8hAeYS94IZL6TH6tSy40ITPiDxuUMTzYhcg9osUXIoRRug0yAIesjAhRf4oN
t61PETiulDkG/8jgpN+FyTjUGAZtJNEQN0/XWRFDFyU4V3TOuzhJxS4BplQKqvsD
ETRDzYOTMN7t+9ORNXAlUHtvbeoUJ+pC2InVrhqorEfFDgyC4qEPQyIz1lmdo/Ji
xNYK3B9bRkiK2n1x0iyadczMY5VV5Ml6isUiNC6osqBgyMmJs8eHUWqdL1MktWUt
0guTlpy9mHw9or+LUQMdFE7kTWnoztAmXsw33yv973nNnnOb+gEj4pCq1U9PS9cE
wHUM+saFZESE427ikO/9T/6/xJjcSmxBGOOBOdXyw57x1TTUi8eZSPs1q9V8vk1z
5IoK2DT8bwiYOWu+blsR3VU0MM6TC70oRAZeqJ6O1f+WITeUtsYIL2ndlqsXRhRj
Ki+LVIik7P/BlW5g6iNQrwllyqF2AYpE0D9T7IIaXiFhkDM3E154VCDnc0vkhjqq
G93oU7nieeifvmEBwvh2Cz57uBrR7Mp2MOLMR5cY5YeEcEw+mIYhX0X17yBl3jDK
bd+GGmVXSiyO/hQ3uC+GNFV4dNG04A+N9cka+9jJDt2R+FF3sa7KH3fC6EaLiR3T
cllA1VpACRF6HkISQvnhh5govxid26n2dQxLBVFO11wtAZEEj3ZYyofnUgCTV6h5
p9Rec+Wz9XZJXR3t7sq8WZo2wtKHXJIe5n0k6w131pAEetev4DNTetVOLgPO/+rY
nX58qxC2KJh7atU5qbX/fhb8fPzo0MkBDw3PMJppD5QPiBXuLT+C5ZGMvKJc+vCk
mW+XXaqLeFDSgEZdhYD95mNy4a6InW/tyLeJCTwJW0yWOh5dWXToC5qrdESMx6jL
EfZLDLKVQWCZdI4hkIr+cGgTYQUu5GCIY7LQgQA9t9tJeUV/xh034cF//d58YW3J
hm2rQYRlG6DIG87wJZkZDq86pBxAqylHkyoft8ex03Y5/tOyQHLmf0jGmZCssUUO
pIMTvL6RJM3PxjWwG04mldzVSe33hL8x+gxQqKZlFClZ4g3dXnQ6NUJ8ZjQVwVfj
d6tZkx16n+qBTN0O8/vDgpWKwr/vqkegJaWSWtHotJx2L7AwYk2gIThIdkMl/LYN
0B1GJM5wYIzStam9AMx0Xic7oluiAt5kdWXvXMkp3+FbYrnud0OoNKx+lxsnbh1U
li1Ht9nYrqUbfxc2Lk2sIrGhFAnH+Sb0vC2P/ZoGip+gAkW8x2DOE1Tpyp5hpynH
U4fqSYxrhmtxS/KiI5MQqSYBdEzhRKcxAlO0YMjtFfhBEgAy5Q3tj0WsnnUZpnv0
jLWt9hrn3K81y3KaMv4CEPJ4U/MXt7LMyvVzGTZltN3BgV5BXxv/9ymPlX+fl0Ur
f0M2PPcuAdRMp+2kVRKLN3CgrEk/15ut+uRrnBB2LT+D4jbqI1rowXKmZX4sC7Ll
2U7EYTAUsU3isv7z345TRmTvc6VA5dB5FI/lx/5ypVpF85Efaytc3Q+07nhFasjh
tyMPd8YlPx5PSbd5akUWUvznFn39wzSQIw18Zq7HHZbBpRWuCrj6pTdv+ohBrLJp
17lPFNQDH3cnVQAwdeTItbl6VQE3h4DPatvK0oc4kB4NxsA8zcMrqVnx191Nz/YV
jiXXaV81V9Tlo8stHKwh8bOaFnF6efthiMCUGCml//Gu5xFtL9Wt3WbyhptQJ1jr
rgEZqDjR4bZTeGbB5wHjVJNncwSNVHu4aWAthJ35J5ycdqjX1/r0+T0deF6uTddd
ZnaXuHpMdx9uC/DocJLNal9DK6PmGk4kHwc4b+qDhznewb43gkparoNR2JQ+NuaP
HtazqgfEskw4USBJGo+yazDtlAwdAEpuFWG1/nK12h9M3Mevjw5VMQtJhOxqc9VW
tazLphQtubEw/kC5HrWkDkKYonzzTMFsozTLBo9k98P+EAoeUogKzskIFsNkVoj3
plOiCzSESzcol7k40iE6guUgjB16DQ1CDfr/LhJaIcrrrVduGAl6ha6glRg1OvB+
Rk1gnlXnzdqLT8XeSOYAVYIPNIo0xPPftFjCloEtdpDJv5HO1YkgzMxq2HHbhBYh
HkTpti2Kq1NIwIEpgLGv3Oie1uqYJ/2vIbSTLk5V/veKcHXkjtYsUY613ikUNLzO
R2VCp54WY+55Q3ZYJusAt+ArseDaR5hOKGR1Uxa/d2e4Hw2OgHgz1AzRr5qNeNbp
1tdF50EHOaBm/48KcYSCKC4NKuehons1P22R/Z6Yg/RYs3viK0DkjKJb6eSg7bP9
tJrW+utR6CJIiWRVpIYMDtSeGIOW9Qc4yOK9ljN4DseXLndG8hlInlSORbGHs6N/
64QwR2pFGKB70a84mE42Axofcxx1klZGivsqVvo2po6/ccbFH9TwMBhWIGQzUvys
vE3ttamkZmQHj9+NdTcy8fzTAHemPS/jUDFtekWxOz/sNPEgZAUnrhUvtjmoHmFo
DGqKG/YrJHbS7O/4a3ADFqu/74c9XsJO8qFmjwvpv1WERZmvNA6VEqSpVxUsawJS
ueY9zkGfiD1xqOo9835z42p7qU+wIzUCZjrqc0iZr4pKtMjZpoptHFdVLtkpoPTb
afIaLLk9DB3qvs4geFubFD/3hyfRgBLEM9kuYHOOOQ7HeU/Gd61Oq1tSf+O+VIVM
/S8UNbN5G2MEPLEE+JgMI76VR0x0209vIcpyjaQ/H9XyqOeNh9Uuu/ZJ13i+boYT
0u3wLKtX7ZdOUEtbil1FTWO+9hwIjcnGJKK16yxLaGmFQuF3EvLbP+Ntw1RHzQvv
tLudLfchj45CLNv7Yg2t2ZvhLL5T3r+r8Vp5IA/3DmW+VDFfPsr3+V4vpL42ektT
3eLu4H63Hnzf5hxGAKAqFhuheBRtrmAG1ek6LeaelXbAiQhTCKXkkIAkoBVnzjVj
/Jr5kR29j6RwZy03VJpviLfP4QyGul1yq1r7Exnmt3s=
`protect END_PROTECTED
