`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGis5bMoaOe+ieuVqdtZQB2tLzDTYilcSWbBmpcFSQBJ4UsrP0iMnLxXGyrac92f
ooUr51S+0huR+wL7a0fTWPBSwzkmHSXgsHfZAgzf7kaavGmrDuOFw3zryt6OPK3I
NsKHBjf6SHMoT7H+4hwVdIwdq+KiOIGDUCOXX7qUmgfWKaqTlupZaST1/EFUKjOA
2XENh+CPPzi9Wo3uW6t8KaPmqnvdpCjXrJHUtDDFrwNIpyQDajnOLrizUtPGPRo1
liQiyNJ3rUTwxtLJOiRbDAmeMRfBJAbnOWU+cChnyffhsG2poxFiAKfwv6f5pgl5
7odrRw/Jsk+LEgDD7CvhNtGnCEvsOGptjoFF9v33CF7WJ5S6j0dk1vjVtXZJmZ+2
DF63NqpJECk3KIIpXTQNMQSrKGWNCpPXDugSLpQCoDgq4UOETMKK1Iz4sgWRaW0c
YyVMySEznO7HDy3H0q2QnTNGod8nU5n0IhbxSyaFCE2O4kYd1Xl0b+lo/wEeMQFj
IyaXsSD0mqsQITJYWvheUBsjIn64rS40KRjAeXUDhV3a0eQ6QOvxcEBz9bZuDsBa
Q1Md9ZGCTl6kZmXnpgRu7nDSiT6vqFl+FAc+n4K0ubwzhC1Nfzv2FBF5pHmwbYnw
hZ6vtdR/hGqoFn0RbkRLPhglNQq+KriMu+JNj8M1+y/SHpMV9kncmGFmRydjYg5z
q39ZdudMPnX/h3if05PL7lsAsCz3rL5EkzDjWYb1HuM+otHRqj0ebbmygnYSEgiF
BIQsyO6KRK0ua6rcq1OyqLEcAhOnQZJ8A7hGjWSM0xeyCrx8Azq6PU/GnRRQimGg
kq1cxpndGdRtcfa8KSSjgyc7Y0AGb344rCmHPITC8xrMgMdwKd5LpenyNL8gvnEW
DHkBc/0I3R9YengQa8vrFv5oiiPFciX7JCjiRF/vXJ5pTVXu0bHkFV3WG51byceb
TsUPydw9+JWxme0tb8ex079Tl8TjMhhg26uegES1cUF5idRS4EKH/J2gyypQVHIc
9w84RT3fLw5lSn8AzJn+oTqWsqTMQIWMdoQQK2vP8nnRgHOsPE5Cz6IPaRwjz6bd
6eICPMJgxZedVVoKyW0zMFh4oAxEuJwjN/uiyaOlPOXVdNlTc2yf3ErmaX5pc/m+
6UJ8NaGBfGaGg4Pw6Ri5mj80LgIXScwV1qisq2VHE9OTB6Tvd7E0YBSYNrf+XiSg
+FY38EXbbz+3GS+Y4bR7lT2U3CSrZbHSF3C3/MtvrryGGMGBlW2gexj3J+FhIkWC
dNulPuZRs6Mb5z1uZT/TB2ZTJillJXW3l6qqgLpUZ4kPeewRar26yQorxxey/a4s
o5PGLivpbWhSND6uDmpmMlDV4pLG7JIYbZ3k05oBiQp3UMKLlp4xO0r2cCh++j58
23L8x8SCOblXpMM6vSYnqjAcXDpwDYLC88fmtTENupDAqhq4bLjfEUtloBggGzB8
qT1SXdfguu5YSKESjWNAEL3rAplbwxauTRCIv13Uwq/ZGjM/13XGB1nGgEvEF3Qr
cFpXVfSbpJuGSOCwM0wBeaGGcQRGw4PGR0siwwXLFYyeULS0Oex6177IArfTFuSA
lJ2P5lyVWptqoBhGlrNQhpPlDek9uTfdX9DwDGidjVx9ezLG2f/bSpL2mqjjp5Sj
NV7ilrD1N+URtdidc5P+ETNn2PdEBOPbJaemu4lKFiWVrVF5Tz83HmSjHmiWEFAW
/4a7kqm9uoVE818wxMvOa9fyXtvSdNG94eHVD9e/QveieqdQ7Fgc+pCUHnv1RCS4
Cs+DZM/hFOwcvjyFbNSpwFdJ5+jIwUHbUE6lmlXzSLd93N/T9LJ1AG2Kgqehqt9G
6dmBO7Vsr5aSNOK/26R4gGebm0btmnzW+Ec1p5P59AyN6lz5scdQJyzTcf9nWEEI
PIkOD3r1PNp0GzFtQqk9UDws/ra8WwH/oDZ9vC+N6Nu2HvCsKE7YK7HcdbLfVTiI
aEkgtL/PEKAT/v82oa4H9qTaROq7jHa5gNEv2FjNiQ1LqiWBD8h54FLSqA1mUFjb
T8UP66pwni7g3MrYztFSuj2kN8lNW5K7Yq5hbAKYDOXdINLGRhtQ+l2QiilwOpoc
Maf1rAGNURq86S/XcoS+Bh/aoXL7yCC+B2KtIgSQOP809IZrF/Segv+EbEVxs4oM
0vfEyFIOyGzsjIcdSJIsvY7nut6q6JuY/8qaKvO6yC+mhUM+yGkLcJehhQunQ502
XDy7xH0eAYvLOWQO7QgsFFEXUxUq0JGpHYAvIaYKuhRKZRlialRMnE5z14cNb3Yz
zdEgEHBg/DYOzSCOGwGPA1E6s/EIwWT2ulrBgBDkajvANFnZK/TDhR5fTVXW1wBY
3DQMUxxuczV+tSkFxUjWDZ0UJDwgFzfH98ZB7/q6/H0hYD1tVe6n7RP/0rWWfrbD
1c9XhWGnMS2AE7LUzAu15AgqnfxfDgvTPGOqg2Tp5XWmnugJlcFp2IpewLHB8z9b
7a7KSVStT8IGBSFBC/bV/j2lOKf9uOppP6vPojvS/SHX+gLqwSbBEMyv+Bb/y9lx
aRXihMSJ5pQ6aMNHTUq0ZdHzG/m5WC7hzrPo/Si5fWnq/0aUha6LYdlaHMUTESc2
y3tRA9AwUOqS3SgnLbOKFYXSZMcAafwMA+6A1aD4XKCfEy84z1F4JPe5f/rig62Z
fya9572mar+bMMG5BAwUnL5Nb2b7it8r8Cn/C1LbB/Bq/hbYBUTKvx6PP7idJR6c
UFVwvyd1GE8cRmS/S2dtxr4faynOi/N+A+WJ0BkLlxSNG3qCXZg3IprONTMhs7SX
LXWTL5rdaa6C8loQtfYBIu5RS01em0mPlB3rICWR5y+jDjFcB37sjBnSrbv8gp7W
8kHlF0dvvI0pHbba0+HGvpOK3ZyLwDeWofF1ZqqFqmoa0f0MpWdPTvDMkirxOtmI
XtGPXKSvYp6eHoHfAtLRizV/cH14ynNFB5QXgsEgIHh5+1Kwelnqg/r3ggxdSMgR
1HbTy4yiq2Yj2e0HX9MGk4Gs40uDwBOb58y5wse3of+VY7qm+s9lyB5Sz3gxf5my
1EqPU6VMnFYYQUla2ktga5beZh9CuGiCi7ESqUA800znW/57OS84T6YOOxVJlCQB
Bq74mXGWgBa51BrrR5VrN0nmpk4OLWioSl3z3PUzKLR1jhsAweNYZj+3ZopfxPph
Gw8dUVCEXiOv7Z+vcn5kep5QSZT8jYSM3Dv1lM1l8BR3RF8YWxDqfmZ/KpqKu897
Reg+rU7T8hVJ/agRcis+y6CXxh9ENShBTidEUe5Qw8bliLAqvgLQr+G1uwRHDmVl
`protect END_PROTECTED
