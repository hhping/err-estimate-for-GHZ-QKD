`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X12l32J9a9x0xCXFBSp8AgklbprrzGwZiVoQdDFVUV+dnv1w9fyFnDqf3etipM3u
CFp+1QPf3USKr+aIsUSRo0b2aRHotSp9MjPm0n5cZj9IReUyOrgnwcQ1sZbCiz5b
vjskRxwVZQ2yvy04FxzPvuSva+XyD66AiN7lJN8ovSToqgPHdJtijK+BNQdQBbYT
pq2qJ+duvNcioFVr+SZshUePaFqghEsbmA+0UlNc6chKLyZ+zBvgyJxufxU8hrQp
PqQSuIfL0svDZrvPZROE31SpYg3CXlZDkfiflJXS8blB05W+jN7xdLntpuvVz7+M
lH6KET+Msmcw/xSaGsYLCSeW690O1WUzWzzkXm3oD3+65k1OLLtaR5mwh8XFCxQI
IzpAct/MAOqjfSzdaPdV8AjtF9HnIvGIQ8M1oR9RC2HAfun1XjEzuij7fcIC0FFS
kMGMaaX898VChKqkbcFhZKrV75bR8hR7EZfVY7vI69oXo76Pqi6QP7avC5VRqI6Q
n+id9Tr9ARNkwtYQUbK/eNHRhmpuGSFRTpNOVGtYAUkrSffE3lvg9rj7SpY/vbbi
jV3FDR6JY2PKFlkRQ6AGNFJdqVP/1FPl4x4U2MCefu0kQkKQ0QX9FdPFDz9B0yuC
2LEeWkNKNdT9E8VHC5pCXvihAB6vMGCTz/Utdh1sInXHISFPecCU1XnI6aBcmb5t
XT+CERodVLlDDMnKRYCVOM4Ru4QhoSWhCgJyg8Xhj2/d8t66BgmlpTri9nV7Y81J
iNLuMS1/vpj9WJP9qOK1mJ6IUQffmlYDlnrRFx7Ik85Psbvyr+ngund4uPrG9k3J
csn2l7zY0QVhiifQRyAyPvjw/De4SCnCf2uW1rWHVkTuZmAEHRuC+ZOJ6pl/iU5k
wnu5Ss+wV+tG3T5z8E9JrJ0RZhkwwdYiXISYOMRLEKPTtKIL8/UVgSnFWApR7wW+
1OnpIBJ3uNYIUfArfAPznIac8pmfO5sGjvzX3SN55Kb72PE2gSIPXxS7qM13nxY9
rFN5iGPfvmwNzqnO1G7GQeVNe99M5WU6IcQqnla3K7WLb3I6Y0dH6wmN2KwlY3YZ
gm54Dp+Fhe/t5myPfeQQUPxgKU5WE4OfozmveZszvwRTmX0X0M2pKhNAwHlHdqfB
iNLeSrcluMxOCvEV3Pf4vLDV+vtsUGLLilsZae+z5EXGFcmEliug2tSefqtUT/6V
uTmzu+DS3b6Kzp/M/SDm/ftuwsz8MGt9jlN9kEWtNR4IDVzCP00Na8yxyhePjfde
BsESyQXTem4wPuD5+hJ4t7WbYsO/8WdEEqW28gimq6+4iyOg5EI18fUZES76ih1P
bgOgO+G6rZsVgA7CcT18v1SjJUEiIbMez5tsyi6minUnyqBx6ZQSvtRxd6MTR2cw
RRkz9G8k6LL8VMG0qGv7+mWekvhBIs7PD79DkpnRd1nKSiag/NsZbo5DQWhMDejW
lp4vynOAjb0LQTmpVTygyelkybT+ny4sFO74CrzujNeg38EWiaFjDiVxoTDmT5QX
IuLgfPrbj3kIag5/SLuYcEF6CGCMhlcOv6tKh5tmWD02RWq3oSGmnJdF1kQKaF47
AOaKas9MxO76Hn1xT9pnAliaCAu4ioDcjVtMJ6m3ZqgbsAYeL++U/qWTt4o0x2L7
x1gzXOlbtytwRW7UnAXbMTm+U97izx6PJQjGCg+bcNC7NXN3SnET4MIhmtobP3Db
zSiVYyvQRzELPPl1gMQQMX2Nr5NAdOdnYD5GGbBcPBDwvydeBOsWrRvGHyEmbLzA
XQWTxkRyG7P5XJtWMVlu9CcMiZ/kPQlhryr/BtIKP9hFvGrKO18MMK5RVrHjd7dS
svN2emzjHfxm/Q1tveei6A==
`protect END_PROTECTED
