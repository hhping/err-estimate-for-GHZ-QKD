`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+bgsFgdqXxrUZFPWeFEPNL6+ymXyS7OABWzmqBUbeD6IDnSS+7CqBFBsngkIPvfd
jD31hIh1ppjewKGHeDwRUzF3q9lRTlNkR0lIlNp9smYlDE1EvgxKXz9rX/Ez6WRY
IYwdA4105CFQt3q4M/78LMdydFGxu+bGSMYyPVbCAiFcEkVV1JhpX+SiXlQ/dhJC
ob6Hf7MIHk1kM+QXUuwSwgBQPh3b7UFWE4hQTKcYzxmb8eCn88h5AlaI2dmliGB6
2l1ic8yhfB8kNVl/ZryaK6q3cRN/xV6hccqzgvr//4/TsyCmZgWOgxO37MgFIFJ9
fAnJ3fYpdr6jybSHbw1jt0gZzkbsl4hvLlJrGphTl4mNsKbZ0OYcSd6aOahc5LBZ
nUNSLm051Dv0YKBuTJaitYdzXXJBCSkg8Qf2PRkA6Y6ExqGfelEpqASKZUqI3mRD
hg/KtYg85lElykK0sHJ95o2ZaQdpVn4VwZD2o0UfG5xEWSr72uYgzPk1dmkuYyfZ
cOad2PfOaWrPc1Yeh2DCKZsGrO9+TOlwNwSYD8Av9I9S7LbMPNwsnLC5zDSxMaSf
Z994Wk3kldjiIE1M6QuFdJidpSxXOHnSQGatyE6DF0Dpt66zp3tCq/nkHvMgbGOO
rpsGy7JywgTdfEBAnCKgNkO6ZmALUnDSvB8oOvcn2XKM3GUxHd3uOPL6C/raV0Wx
IXKVcPZjPZZT0/RXCRtKpquJZggG/abuGdI9h0rM5a7mQ2KXRzxZJUjicFHygkmi
6QMtJcOnFA8/pKTsYVBSDIWAZLvz3TWNSC9lxwdW4FPmUparDawLvjtqTplWvdqG
pV293Fpju5okQ1V3Az/CDBMLxb5BPFB4sRb8eWExVqX1jlczn7nEAb/9qXcRnSE7
10Tb+62WQrLaFGau/NVSFZOMNeIgijEbrFYkEjKk5q/DkXMN2ym9ZH4iPEcEtdXX
QnaDylI+uee9cFNfEuFbzlypRfKnd1xGyEycy+vkTBIehc7y1T+vrduVVbx12E6v
CjLqsdujxAKijOtYhBO0isdmfmKLyKCfNT0re+hXd/8=
`protect END_PROTECTED
