`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gFXZ3H1ENiDKgRbgqL4HOHY2l+uI/Cze+yuihaH4TOIVwj+2QvPQ0A8t7mG2lNmU
NpNISwg2KZ8VVeXiQ0WA3BsfG6y47SROM1UqMLjDDV/3D/d1Q7M+mk1igJLwSV2i
5e+ncmB2IVpihLICD/E8SGOIOJYV1qSEN+ZjSUzM8e+Vqb5katIEj+wJx12n708J
yA5qdEV0NxFr/NLh5fQitNLdFd6wkznnNak5O8xqKG3+Z9Mt/MUIIuiD8U6QKgSn
EqBIUGAxvhC/cb1y3+eARRpkwpeQLJPRkgJjGKWO5xbt9pbzzlg/5pXzCKygpPga
ayhqvFSqqrs1bofaiswUWBRD23HObRCB+nqtbNFfHIyfwEEuUxFubde651/m1pBh
7WjXWCnPZfr4S+WYN1fIQGSn062ldsZxZQZfS/vEAIc=
`protect END_PROTECTED
