`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGtU6o4a3PU9dyFZRSSNlc2Tjhwvo6RakEVKASrHhT6rmO22DJRYeEUth9VG4L8j
fRLIYzfu9+UwBhMkxypzzzJGJflzXUTMWErl5TCYeyDpzeFY8NajOuAzqr8oCPqh
RDxtZurVauAVqP1rTTb6FzS91N0ItoL1fQWx90Za+hFxLykpTzIpbus0FT3hg7AE
tqV1CFwN4VZByUIO3bTt/iHm6mw0uypDe7yWtDXPjfrRnyte31qy0RvEsz0X4nqo
mmZUUXxWuogeqbAXCxnq1KYPc95SoToku9rATlWw8jnPXQUaUzvNa7sTMPFeSS8i
UEmLka/crIM9Jd82BXBwByDyPkoUpRQyLqhix818Mlx4spQapGhOUwUMbo+1I+3M
dzJnyLP/jbuogAFB0z+gXbWZEDKNOjQ5FpBsSI1rzZAIXOWWX5kewkG8fFTUcL//
/zFfDvRljV8ly5tgZcgdg468SOUae10GWbmMvFDbaErbh1w1twT4oeGsIjZkhg3N
HZMehn1FUmtcA14kE9IszAPqwSPqwjFphoz1XQexGbIi2CJIytgHgMabWIVdXTEU
IddKoP1TGeo9FPL6UxUcedvNVBNGwRbbyIOAwa+IBF02ZSHdEw4UICTCOtkdw44a
DwdHf/MlAgIqyc52wYydxo6T2GvINN2jGaXWQXyR9eFNmGpAgO8Pf+KiICRA+7yY
HJN7K33HWnFCmm9rZ0KQWeOKhcayM9wP3ZmBAc/7l0Z01ZJJU2xP6mZ5zSsjP8Nh
+JoPbOrpVfludARboYRx7qNJJ473nWDud30Q6CKGazGVEHD4Tt4cpO6Sg5G+cJ4E
ePlGTJIC4amgT/86mCGRdnu35mHyoVJ8ltUc9p/jJxSvBL7Yt8/QDtD25oq0/M0n
molyYk9NEvniaxbS+eNyxQIY2RZ/E4Q+zpYKDDZOVLG+eATdtTv0136YnylK2ch2
6htkl/TtCAOopFZivwMSrmYsifNS04R1EDV5tWy5XBkcsSheytj4dURM7oXGtIRc
c30eebkPgy0Iysneg/QutFKOmjvK59Kg9SyJ84LPteJKRANqdHkh2antBf3tbs30
V5JkJJH4IFxLW+gbkhn/3TbcvUxFrtkokOVu+ZVbFcaDFriiEWDg03h7naHmziqh
uopz9h0QwU6hj01aFws4JRBojZGUrwls3RiS+kEr79YLA3dX7U42xgqmfojDDBWR
O5J2ruPJVDHWbKWyXsFkBgQED2Qo2G2A4NOmeKGgh/ZyZeD8tDvRaLWwXbYhbixY
hihnUCrzZLzOpCPD6EbTVbVBHIc9BhXJ907yKJdWgCW0eicBogiFcKtdMkp+TuTI
LDT4b1c0P3jcmdkApw3appy0gswTQyPkY+KR6NqSd9xxFfurTvqi3NrEjV5rpbU9
Sg7R3mLOsm+1uRHJ77w6ETRaHnVn3LNPcNxqGYW1N83CmvRBuvnZ61Z1lYkVEU8F
MKOGqvLOieotla+ds0wIsY3K817/DGMj7Sd0J+T0hVbxTbDnI7tR8hheCIWX5LPd
gyUuzCAUEBsPvSrWum9O42mXXtpdCMTu8D5ndpfMQ9zW9E0b7abg51A6GpXFGENM
p09eNwZtJ1aEWoyjE5kx7qly8AhF/u5GmW34CT1JxLbNtiKX5l8k9vYvOTOxd/Pf
RE4migxd8I2dHtz0Af9TvmpLQwFknaSqfGcGCJ6QxU6nrUpIwYngev0/XJ4gw5yv
EKBTrs5yuC+rCXucTKsQmWmf8MdAra9uApK0V/Y+YCXG3K5k7hOFqqLruK3erGKX
ZdHcoy7EYf4EkikQ918Mad8qtwearuVTCTetpzB9b83R14J6IDECD46gfMkHuQAf
TccTvp9Lrt/cnfDB4nVt/dLuRk8bVaPRUdUFXM+/UanGtowUgcot5XMVrzpwD2CQ
skACwFyXqDLDH6Ec53a3zFSw6aslaz5iGtNnC3oIgOch4AH9Ijmr9AH6lt5StSCc
YpoVemWKShxzbH/USJtBSu9gwff+RsdJe3i9VCgfvLVmJu/8tnef8FLfq1f3jm6x
+sG2DVyDMRTPOD+JySvNCKWX0MYbCy7mJTSmLypn3oFLoyJFmuDwud8EQD78TR0G
04iGF/pWl41LtkmlD3NzvmY2lueHlbUFN0TjyE2fWt5Oj2w5Tgh+I/wNZ2XhTw+Z
BeGSKDz742MxyAReFt0KiJZVhqg5ewze9qlwJkRHPpqU2EdRalShny004a+eKjS0
GZ17pyDHJ4MV2Ucm3XwSbffhFg1jABKVqs59t6BNlyWsycRFnzdBFKvJ2eoNXQsg
to/vtqnZiJrgEEwQOo45T7zcGl0ssONjmpGs+PDKgcn1egKaz7cjHl6zHLkdP8Af
oDgAi68QYYqU41IEkF2/FBE42rGtoyB4MhtNjfj3rXIz1c7gw8SdwpxOUNAQX/Z9
5cQCEa0JJOzLE6hoc01gA4Yg/sz6odJT3d6Ts5MP3WdTiB/lFLj3m2CiRLjTI7dY
/mys5TCIuhH+KmXT8J6o4O0tPI53QYqWRNh/n/bF4akk4yqDLnQbg1AbsN0BS7KH
5kSX0ALucd/YZ9riMlF8hi7FKsu1sRN8oTdrPyuLqAeubTNkKJXYLoS/HkbJmnpi
JMnEWFMw5OvpbGWDwTGBg/D1dI/YxHLIWNz2kuAre9pY7BwKtYhwJjFV22W4gWyX
OnD2qACm7119Q8Ucy+dr7Wqyq08AWiimPlLi/KuKxZ6eE92ZO99BHWyMKC2VPRRm
84C9u12XenRghSPiDvoZfYxZDOpQiRUMMjJ8SJ//oGxZZN1ilqGKxYz6H+t+V+Xw
syfU+LsAjfVhb1argM1DSiQdAgQdzu4frhKJJyVGxtoYb3YQuobYATJBtx419W6U
/B7o54iERpcaVXQEPXZ0pQwLN4d7Xb22R28LFzcmfC+wY2htDpPC+cWECWBlSD34
TXgxZ/QnoB87PsZ0wFrN7lWtw9YsrXVQupWDSsxMqYhj/4XUe6lxkkySEHmShkRJ
mAWnx/OV37NGJDK9TXAfWRWVBNp9dFJTHZsh5yVQOpvnsqNSO0DH50ts0gmCB5Po
eZNQmodL/Lf3gn8ywAY6zBS8gEDRWsp/GxEysWqRc7salRs4lWdsyvtG6Y0ZYHjH
u7etTKP0bp5usEvDFd37NzzELz3vkJUkvnQcskZNRSWagUNsmPccU+RtlXPlqlQi
V1Tc+iU3nd43eiyH408wo8xatM2giGZDAqOdyRRQQZ+/JZjIDM0+cacAVdQhapRF
ZNlvO/bH7hif2HGiYc/76DF3Bb7ZCkXbDvq0dkeL2CHBU29hsirOxptqgcse7doK
9DgWgkMv3ajkuRDxLHlw+8nMd4qaPPSKHv/9rVkr8MswE0hmZYT1aw3YIgI++hNr
YPUTEQPXeKiBYNMigyPTuSjI7y5IlbYu1cbnF4IRzsg+CAzBBQ+a8azsBPN8pJA3
twhauQfvaELRfKlSlMxWyQRgy382vYIomHvAXM89Jik6hu5BJ6MhyrTeZSr8c7Bc
XPVrmtfcZWJE8VNOesnQDfeNuYjkz+jsPmbEeLx5gwT36T7tYL+76cX59153ZKpt
OYQCtDeuor89CzVJoJAfwErl0Q0zFy6XYRXMAxUI/JYW4FSoaC4oVzOCLM9YHp5D
Eh42RzZrdOJ/4Ox9pfFR0/qEKKU/V1Hx7aiy/5QXbi8uQOrVrBjVK1c943O7ya0y
ua/ATypXHezusvfFwEUrJX9iwZ/KxpxSRxyE3+8xvXhGnS3qYdtjEPdg23Des+PJ
xeYA9sQoOE8QElOVOG6SZzOdtrBJLjGliiJTTmL/bNjKFW9CWGl26xTmf9m8fRnS
sCBeGvc3N2EYfmyZV1KypXZvvBMoSqSwhbsjI2/87Z356C4NKS4Rl8VlL5NfCfxB
NAcmhhatZTOnPLr1rHtx6cVNrwNFvZ0boEHFLPgNzKO0/+RW/MdEXCF3WRpD4xdn
l1lP40UgFopJPwnxBbhU0NrU3cpRDi0LPw1Y2/qnWka1Q6BOMX9/1NPZ6B6pZ+eY
ynfAdrsieFOqRhSe3W7gWU41lwJ+ZKAuS1wZvC4aMAH9kh14aefhckKCzEaYyMaU
GHtcQSic4zY5nvK17n8SnHfQHjJdyEvjIlJcf7K6uTLaOmFajK8Y5K5L7ZdjNkSS
0OZACglXqn164Ml2D8ySfdR6g9iI8NNLFS90Y30aA93P/JXsZntkRrv5jnnz2ZPc
zuFkcAT2zM5fs0b7hN2ZFRT0IAp60MxUiO+OdB+WgfRXdfQb35/ymuqT0xQiajsO
uHMXE0xMDXmMCa84+D/JGkqigN5cMHxz1LCXP7d/pXPBei03vdodN/uv1T7FG2jt
pOO2/N527obgbYSYAoiGpUMRQL362n4yCYF9CpvmvhQQMR0OGZgRwoodh5EURFt/
/Mk+kTdXVFJfZA34tbNHeN0Ld7cuAw20ptySdYwH5LilHCdX713s0anIhpkhq6tv
6V4qhk75inJcSIE/3+izsmmWBMrRQMtPFSHp50ge2Kha1dxmAPBOWf3KdluNMHnV
IWGF43EzfbzRa0kN3MUihz85xtwDDG5dPxuv5h3IA8nPDc+eAQWxJ8AWjTXI62+/
XM64CKbD7LblwtaEtE+GGe5eNBetTCs08coXnu7mD0JBBBw/JvA5nq/rbMZ5EnvU
6ODYoQCr6t3YRt9eTrXkx9LIcGk7iCtMZj9oypmNMX488Bs8v0PMHzKYGeQKhCYu
iTUX7MeBTP9RJOTyChrXTbRQ8OqFftlcGtdZbwJVDhG6VWT5goBaTPcs9mXKGWbT
YMrO2xmyEKGG/W3yg3mQCWdaLlYlrHzro3k18TOKUOpoRDKZaMahjsWIg+dCoZpx
cDfmeMbebCwci6N4L208PKMrwMgIl1WQGmP9+pCrbdgp0dIbcbxxn/IMXhOR9CRF
x0OZ7i0bf6wpCK/kfNr4/QdZZZEj+i/Awa0HMKcsujHR80CZU29aCohx9QBdTsJP
Z+kxpXQTL4ZsbBVbgZgw+QuESFrRedFKyUFyDIwGqihV9XoD8LfVLaBXystkpu+k
ocUL/gvwZ+INHwkygPBpkZ88IKMSkUClOyRx1TzSbrf1xc7+vOXR/8wz6VFvfax+
948DKnIqBQMdgnj2dZxCTUXSUDIjEuEnk45CEbpcMcVXsJBHY3s1DR32K1xACPTI
6Ufe0ZxZn7bnW6ufsUD7HB3rUlZAJCSFssLSKul0h1uiRmfRpOe368HFoX2Rx3D4
A4cHumhTMcRxG+w7cs4Ci3ZF36CML5D0WVsYu62wzoWTP2498R5hzoLraEmneU4t
oaA/xV6rWDf8Tjbt4O7zL1Qgo+LoDsrbj5omxIVPawF7GKbsJkjBumuyQl2zs2NE
kA3Db2Rc45bT9QnirKfZsV2XYX55LZyngQdBGeNaIr3wpEk2eEw0LddU5w3jlJeQ
V6wO1YEoND/nFJ2gq0Lr1dhmDOzr0bD9/VjGkkpp3alvX1E/0bbVkFundmTAKIoC
tqS0a9vN1NPjDzdNJqL5wO16ECIudT/cMOLfT7Oz8ob5EkKcmNoKdw6sqOOLadLf
AuA+ZyElMGIjBNF8kvbL876F1rQgv68VeyF+jlqzjNRTS9+yTtPyzH/P1ZBxB61L
IAKJAi3XFl39P/APTR7XKkDAO/wUAIcwLqkSbHT0yRwiSiUgTWeHubw8i/TJ7OHF
FA8O7zF5wStgde6V/+OibKMB9Rbzj7PrBG2tKhzgG5ssCqMyLOIQdHfbKzHIkMnk
90ttXfl2ZnyURhw+D7YESCul59/HS6GxWalckuiWs3zEG3HkLDYAd8pWs1zhgmZb
QYrfwP8g7f3Duq+8Y04T3n9AchtO4vMVZCvNlCeP7l/Ir0VE+EMrGsoHd1xCj9VJ
hH/vBrDq8zqUWHwviDtxo/AIIbiuJM1yW545h0KHelhgjrpcvSsUdzZRNdItMsKk
DB1LCHvmX6WgMLHS4rIPQwY9Y3RtszkeidzgHETFtHd49c9AX8q+En9+89jwFX4l
XucwhvBpwBjhQg4MkmgyA/17Ex4HCotlHiYXJp7799UUtk7co3x4h2G+K4FJnTb0
8WVGZ0VueBVpEbSWCBLyeAH17yvOyvC3RPNU+r5p27aci03XPFxE/Z5NlZcyoUVT
OubMIqs794KdC3dBXypeSSs5ipOGv8zI3KOBYja+SwM0tlnoZc9yig96EKGsCrDj
N4gyIIaxZAxQ3c4hblyQeybw2JkZePnMhY0henGDiUgE4upyGE/nbtgpq4twHuKc
k29hW7HWDTJ/kE7dOAnouu3rzcbS88SiQHQZjM7G7ro6uukuQq/QDDuJsRaq0cc5
H8sy82+mLYJ36DaCI6PaTLODBUj+o5aYJsMZQT+KYrIeY7yY7/6omFwxgcv4MhXT
SKt3Ah/i3v46xB3uC2F+/pB41NfhDVPLRjvCu7cScmn74beiwBfHpTVkTlcFlbgW
BPQiuwRRLDRADEPVUIYIkz/Li6xfKifYma+YMaV/miV+yxUKkDKhz1qGyWe26KPW
0gOBEa4jI5XlN8C48H+xhH9WZ/jGBB5qMEHyxunZn6bte/8+/18KroUlW+RG3PUp
AHUu606GkWUf6HcGw1tmd/LvHtRa0jI0uMZJBDg+P4Gbd79ck8jkp3SUoiMjQXJX
TC797rIt30/93ubM5CeYg+/ifNNNJOfqp5K00DSQ0B44duOkM6/YTyuYhhnWujWi
kF4lefhM7/iK/e/4toqx4jV5328MffFvnjwAgNKNQXUmq76LQWn1+T3Pgz3f6+86
otUaoOyBvRUbUzAFcTmBUa38mxH4yqbOkwGKdIjDNwuNWrz6dY8UiLhWCuW2tRCj
3P7DQec/OxmXimWoN5Ei6P9vlv2fjg4OYThFlS7Gbu9pzFpK/LliKF9ErN1wB1td
3VLjVgxb0eIl9yHGOkd92UBKHpdodb84YhCpBpxHkvJX5fr3k47XouFfALUW1eMr
TAOwYmcF8wy80j6a9/HI4tWDhAXpgP3Os779l7rf9TRwb26zMYli6qSS5dqTRhYA
OAeUiDXHskOElocjbcqAh6faj79eTCWLNIXjZN3b1wHOVQAd1YpJvlg8yV4w99Bi
zt9KKQ4Fr/mK8RrgyqTjd5SVUH9WhxKakaH2LK8MVvR6dmAQrn4ZgNrjXKGEVNVp
xlm4dSWBqefnH6iKVPvee52mh+zlO9Np4M6T2aXps9Ujw1U1Zo7kutVsw/SoJ2MR
hc/OTbS45Fj6BhwBTU0VkBHlVxRT/FKQA1fFDudYGGNQoZfK+idnESvJwvk2VdrT
/Z9VmYFiXP0e5SEZo1Jw4Noxi9RHDY0RuioxB2w7hR4vEImjMRH9dH55iR3u9HGH
/vc+RV3LiXZHa5j3o9BVbLjFH4jND+olei1+4nPkSpgzIruVr8uLcINS8Rk+52/Z
ixm/8LWayd0UbmQ0iAxqIBbm4STUKddqwwmwDMBTa/DAVZSd8XPXpnTtXGlkiUHC
UYp8rhIJUCY557OhKytEQFVkAH4R5rmKdO/37KUeJSO6zusGU7j6fE1/wdNmpcOt
QLYFxof4k4XQ0zM4qPWxBiyT3uBqaHhg3rNlhCW0yLm2VAc+d+wlJAalLLaHo45R
k7pRMkBhQ68ziWn/06m3E0QoVHECvwqGRZdz0l2EAAGejWj2yV9dm/+tQApLgzY2
ANub2/0iHy9qBMJLRvfaOMEElDDTPa13amH15n6+6AK0xkON4D0vutkTiTw+firr
YIcIUoxayAzzcslsFG3CF3yZUqQ2MrebsVikmoOUvCcgkH09vBQTfJl8A2SPb32S
WdyGaky280poQ5JGE+R3zas6/3ek+CKAWCnrIrAXbsVWifRAcP2cRpufMi3n3Zy6
FfQ60m52x222PludZUcYLVi8Dk6w1ZBuQT8MgHQklu5X30TToCwQhqfVyic0se6n
T03BIM1wbZWeUfofyj4GvKChUuHhBuHkHm9fFyM1Gcx2ecmiRf4VlfHGGt2h4coY
e0CfONCFaqzs/xwNI8FtIwb+3s6sdngLrqpBr4X7lGp0yx83b5NtNqAYkUieXbUZ
aTTcGhfcGmcxTRwtq8SjJznS4zhkhUBSqaRXk4rK0xYL2e/M5uGb8vgxaJDm0YOF
OnksMEgGBzRo0fkw8toPzQKh6y73P7wND52Y1U5P1SgV3MdhIrUpJT5gCtQ7ii3C
OpUPll+SxgJlIzF7a9Wfr1y+iFmn+qc1k/Bh1UIoJlA7YuzB3C7Ic2TkeZkiKcS8
b/XvGZnFpLNaV/NreEUsIT9hgGBllSrnpGsGCOPJvNdgH6B60/e120vwZUQDMiiZ
8R/K3QVJwuREwSpCRHlq8S3pc0BBPsFxTLEVf3arfzfnzDdZbSaOHmqBQ61ut4ct
mmDWO7SxLrlmDL7r1kD3Syi3cvVgrcUDfl74oABrT9Lc/t6SMtK7KTIX+uiDbqMi
CXn4PDLvLyNtuN37X0BkQ+cW3WEkYFTbHjKI/FZc91RtsPBUXV1jp9ptPgFvDwWX
IneIO5D9YWhbppr5Oa7umd8PyXYgsWzIto3uZyEbYwIOzFcD0CVryG7IWSzPJpot
7e1toS3hPqmLFqT5V8EHr88YWfaJd/lqi7vnuWDmmrjNoWediVDo7MWxS9dZTz06
D8cRAkD/EEoNstmXi7Hi+Vaa08Txo94mUiCTSJyzdfNl9yIuxPsNTxntGSASydSZ
e9Xc6jdOvv8D21PP6RxYgJ1mcpAIzfpxYSjxur/+7ohJQA3VYonEHxUdXV1eKu4i
wW+bMBp0+HJ4WM5vBmX0cwVGLc0U/j5fpSo9UOOvk2vZOAn9XWQg0Kh7f+tGDHF2
Hbmm0KU1+sdFP9T0NaqzYE988RalTkFK8b5W7KSINkEp2o9nbfxXIjpb2pzI7Hz0
4lKV2X7Iz//pSbcz4jLH0vqILVgKEdxOjMxMIrwUxMJNaTDwk00BmkXaCFGb8NeO
x0jkh8xjQ/zlIb1AuuacVRYhzrbQoyN6vlVNztRdlgzzyuDuSz0W4UjJO04DLvLG
Itpcz1VCtBrrQ4lvF+jVbmLE43VVZjRWYP/+x60hUYmS6dLv44CaDESY+PVj4X6p
m9fPq8dtclj3UivY4rK/h/C4X3Ss3lDabfB/IvrQMXT5Ae6cFjhh6zl+zCjLFPKH
5DRuulgv/OtKzT1NUMyFR+bg4OTL8JKg8HgAY+bnVGKkNJqBRD1Ku/2939ipWOAa
eZ9+Tuu34tXCbPOXyDI7D6iz2q5WnFQKWN2WSuSMRBJ23IPPBQ2cp35FsvEhmhS3
/lZ+QVFrrz6nVj6MmZCD8n5/LSQIFJqVy9orAL5F50aAWkXfjJsjbS7On9s8Btnf
ootfT/v8OnHqHYH3SIOcZi8f6dDPLVVE0UN92/bqFf3o6NT1hNx8KEHilf3BnOmI
8D7enWZOq87/t6B/eOvXO9EmbqVuplHbP/V/C64OtbDm/7PAa5svM5e66kTvUXLF
qanFSbzSiZDz5Lq4rc+E4EyPrN6urF2IiZwrPidc7C99fV4pMfp0W0zH0qTG3xMD
SA0pjB1Z98KMEFRlQHoKFeM4eytrjZQHNJqyysDTROQqz/Icy0omSQbIQTCkZO7F
+4FVo0F0mhgWQyxX8g09sdw5VKoFD9mATRrBk89X3cTtdm+pUy4yUh7noh3ZFdNM
dv6cWTqAN7uQaiL+ujW/v1dWDxluqzu4pvSG1n9siQ83zQm19k08rJVB7Ks2ULWp
1U+7/WZv9sVbHPYuDvW/q4bor5OVOcMs0LGu5WJ84Txrvg+U9JJRGZWXiSyNRFXA
VsKgc05xCJwOjtw/RC8NjOKYVrNPvjsGK6scsrOFInilaiXnhymGY322fqWzI26n
K0OG3R1koZyYUMera5i8LYnQSc8k1e5/uJJKpMEVA86wTjmArWGEnPBddrdomFYk
Qhlf2N59vnxCfLkYsBraQrB+1YWWYKUbtaneGOUN+IAqdZeOaDBKs/x/c86H9Ys6
bacNalFAmNolcWSE61RzqGbZi7YqEHZvJxuLE4LaD9d89hbFsuet03PxltTcKBcc
U0NQAT69zOGElM65Pc5Fsyvbc4VRQQAUPipah2TYsY0qlhHaVD4kDPvvrJLys9Ks
3qlRlUlI7+NZDRxXEobUh7yQyRqAD1GREf/O4RvqbRDWd6Tgya/5Bhmx97dcyjO4
S3+N7P/Q936GOhOBfJFIBegkdkqBNLKRo0t3fVKzETcOdVseXDP+Gk1WyX7j7Nbu
u0UAOHoqAlcXk4fuAiGVp4FWlH15dSGrnWspJNWXYzVrccNnJ93zM1aHN9cPa7eb
mKlfO/90sc8HjuZTgnJ4fA451Ojk0MfZcjBoQ9UYcoadosfpH3gg4XIZAcU0jDRx
liHzyyf3Hh6vTHARd4j+4lEPoFiaEGldMZTZmY6ysjTlqi8GompYZ7GQaM4dyP2c
cDQ2DPwjEpshENG35lBTXUzFrG3zADs6VEtk6JhrY5xu34NiwyKAEYTrK13/oOQh
DeNpV+WLIJD+2fv7Y7sLUZee2HQcMan5fdsBA3HKyIWvyCGB4Pt1Ttpk0vGCaGBo
6D65XXoJ0YkNpGMKmOa7WMXxZh9NY4mjv1NClzBbGy/otbJZTZcd5/7WjWIREM0r
LvoH4vHhJ4SzQWf7UmJDS/W4e+upsVduDDbkKzs0Q7Y/6JOr51VW4vhoxgphKTUG
TB9p0+04VB0ktTDpwhEYTelF0CmFlSQ40HMZWaT5tw9fblpvHmem3Aa7wC3qfQtj
lVMaESM/VTO1dCP4N8BROgv6U6s9+W+1KZ5wuiztV2RRwgnkEn9EOSaxP4bvO5cn
l4n7BOJq6vUPVJNmHfmg7b+WnPW5DsmehzDLKCI6ZwzR8ooXGyKf664lTy1A+0kq
l1+cfDiFxuRIaceiTiHJQkZEL+pMSruPZ+C741LNu1XEDjTS6U5UadEJa88+20Jg
kANKtYu5prcfmAAtr0RhScJ+k7tACPEMNdXEwWPVYSte3N02Kgv6n9RLUkddfAMD
sKCa0L0iUTIuXli7cI/0T8JE4IEVetbgIyhcgj4Eav7G375YbR8ozRFsbNJsScO7
6Vs3QNYt/YdIF0UZ5sGhdD0vOD2tk2EAHcAroswgVptYq2XqPtBv4edTJIWWc9Gs
1pN/vKWfBxTlkFkLKy1gYL8fiUjObWXJeWc2l1IlXMg2siGYHdhGrveczTGjt5X5
ThMCGOI67uQdlFE5XQMjHFWW4dJzsO8PUKyR+rtLvyOaqNXSGiJX2MMonim49MLa
TNUZ95xECgAlj6I0TSGGnHOH1iL8CdcYeboFrN9C1PZYrgXaqZL9y4My8QOedl6+
K3bnOwTpaVKUPC8We2yYr3Ot1dFAP7GfLl33SM93h6dNuBegecUAlSHFt0V6lerS
vkTH5hJDso93z6iz6QRx8AtBNCMyJRYfH5op+K6jOZV5x1qopfSzVVY5Mf0cbROI
uVvrE58Pb4ucpu1kyCSXV4Kx9Zv1GecyYB/Cs/CG28gnIMCHFcz+hzqTA2a2ZHYA
Fnqh+jTacbvaP3HP9+TjimlYpRx3vmzoqVvy++lgVGasi/rAznrKRHcT89XPl6c3
NwlPEALxSKU4PeyMwCAMOd8nqXLYnVreNI7bA8kLkAOTr3fL6TUpOW7wWvipLqZi
JnEoB1vJh8d+ln3Th3d5ZXs3oDxW4xDzd17NrTP0c5fYgppCz058lKox6lnMXkhv
Vf9PgUzNdh+4klxr/Xf5aigR44Hv4Ubx5ZF+glr4EqezVCelwO7aY52aFB513TTG
RiUbfWFDK6nC6eUeLrdKIAH8SlGb6R0tVBRPckBa+R/7YMsPCYST4oWg68kY7UwE
7WZPfaJOyaeJWTWuYtD+HV1FRuzCVnt6v/c3w0nf6Ln8F1KRQAKcD6hr1eW7KnZW
PDFQckewYBsQnotF2u58RY7vFujv6z5KoRbd2hgFiqw/aR84b/BZmT//o1FNXDYn
P/0x1e7GYE8/cN7abzUg8HIy/IvKZwsEp0qcs1Fs6eLcTerrbz4H8nbJ/rJdusVu
YF00y7DV0gXvd9koLYBTuKZqfB27vsbLsuA06Y1QItc923hzka2oqvxxDBdUmXS7
g5glanYPjlWcwoprJghDouSu3GKxwEciIESYNe6Qfh2UPFo6kqqS12UtwHjZN+JL
FAEWdEXpXfAvXdYnsauqW5g6tZY0SKNeS5XIVtdiyiy/L6N2BzWxiXz2Iat9zZPO
EuZbeDxecZP9n+w/RxyqmqEBiCDq6S9fgJRa+zobxVC+XXAZGhumGBI7AwN5VmZ/
I2hgWzAYluR0zwUYD5xJZSGyeIMfU9lBhyK8Ki4sRGDGmhK9bWmHvQO0SSXd6t0v
SbPB3QQMHE/xqzN2me6fSR0qNCjvFTcXj+GLXzMO67qo41ZiSmomtZbYUdZpvxWU
jN5sUHjgwlKIOnVULUm5DiHCix+0HLeRM6/ajcIY87bFxAnv/kiEw+462WtHlJx4
EgLbEG02t8/S9BpADuPayaCVyCQTqgU3IkxfGQ04fBh+jSSBKiXkaGUaj8MCBW1j
HLdoMznwEbgjg2niv0Z020Cx9ngb273+IMNbmb/ngvAe3QfGZY2Jg/rqJzWMy0Wo
H4kmNeRC/A7Pi8XnyM2C6jE0e5K0wv0rxT/AshV9S0pI+Yw/QKfp3lblSKYnXF3y
uHr4pQKGS4v/TG438kMnwbLHj0RIm4wGGa6jT3/YONdPqIB5aV2DB5amyfDJ31Ir
sQdCBOaxHzi/MExfiYW4H6pVhDtc8a8QAB53/zj+6V+XzDyyO3QWSv798bhlr3I9
UaCj5Rye8hIIZnqMikKNT8J8GLrDMu43AjPDcqixpMN7TK/2qWfx6YfM3GKr3Fmv
iV+Aj9DsFa10PbguJid1Luu5aJhs949LjCaIl9ChA+GOJuadxaJ/AvZmYRW5lm5F
n7mV/TN406uesUWaVH7smu+PiVEVtEP3iSgY73aojGD/Cxaez0minXfbvAafefv0
RzEvyIRP21cEyRqb3KhceT4lME0QCO9bNirM8uUt8ghvea/obXUgFOnv/KVwPJ6K
480ueo/FCrggJfAcwjdP9Af06M9mQOvVWZrOyLpTs/IoM4Twsk776yIaaoTYF96A
C+kyY6yndjJRvQHQYVPaqS4wBxwX/1Azvgs+sqwa14G75nvJOH3/eKq0b8VaDeBe
624VOxi1rj9yVZ5cbDNIBD8Oz6BsdvQyT0bMACHDYvcncKEvbALIxdKATUhLF1z1
U33eEAjce099DA/keswDVnc6hRT4rr6DTNZqEakprbzW6oVEeE/HoKRcjktCef3o
eFtdcH+wsRogRZaWOQNNG5jVPi410THZvKtLqaK+N5xKljaJhVCNXzFi2np7ITUb
0vuwoCbeLLah9ydn6qTkK1tk4qxxVjnZuM7gaxEe6WqnxU+TCHiFcY0LCfpcPOuf
sIaVY42no4aTYSyejMQVVLklJD00eIIoTSAUoPbC4jF9weH9lMBfab9hlmulxnHH
ERFjWZKa22Sx78VBhkG3dy5UK6p8w+4WWhVnCjoiwLutQFoQTVNJ2/wduOUEESJL
FmnF5LJeJMEACqV2j2XQ0m3oml2/VF+zkAFSlS2HGrj1yQrWwBIIhHXZP38xeclF
zH0OUB5NZMLBb6Wina08N6w1vmPav3adIUB/sRzmSPhK5hT9JOzsjTPN/X5B7wKc
/kxAvef1osb/kUcDURENedB0LdMnb9eVsIXaqjeB4YyVr8aNWiWkd4UkMvtaMZ7u
dg+pKp7FbnZDR7WUwVrppnN2pSzQGu5GC8J23lMmi1RC+ZJ3047Ao6IYRXkgdNlH
8Jck3XPf3INmIKPEXLLBQqnm9DMLt7VP6AXOqHfCWUX9rXDgzoqW4mClKDRkdWPb
E7AWuWcdx2A50bWUv1DjLvGFhQRlREqtQR+m282JZPKOjejud/aECWQWVArWDT7/
eiNCJdPtWszluJ6YjEaPvrQJQYK0Jmujq86r+EmpuHBKLoyGfITibZl9BBK41Fff
7pxVLyQUOMO/OqglhCERXpxLqD2fL6V8AoAjKKSZyVutdlfYYcLgURb8E5GpAXgC
wMj1cHp8dysj+DbBOUpQetiwtUeWQq6USIpvBKT6nDdrtdz3bDfMlRkLky4W52V7
S2CcxuK+sBpm1sG5tJTLdn+3wS180GYNYZ6DKaAT4vgMwnE0xP8Yyn93t5eaymCT
QSiMGWPH+OYPxhHo1c94Vb5eTYelrF3a82yd63/fu097XZ0qswl3gyXQO2aPaTLT
HUO3PbgJXjEaU8K6OXSt2fYmC+5UGnVEzDSjRYhp3cTgh3z3T6xVwCB7q1MXihgz
pld7kbni6oDNSxg6AX1HAR6gvrBqrSlQnwqzYxVzA7ixg94bNMJK+Lq0ZW1RBAeW
/9F/ujNmoNOO5fl5NF6uJesFIwxLPRoo0AvQD8SWMYfzosP+1AHx/vbpvYbhuiWY
ce5sKqmoRWzCGRD/LjX6fdKNmaadcWwim3wpIKOGN0c+HhJp+Ff3VmNzSflOPEZB
IvuEBmJtsUQYSIbttvzhopuISE95q/n3IYnWg57B0TBOmXmVQhulO9MNiNRsa158
z7r6siDyEInA4fg5eUzf46REU9iK8LxjJD+G4mlDsnT7wZS+suRgsP860PRnov8a
d4S/5DsSA5Gn7JKVrOXR0FqB7BhnvHkUqiIHipdM+QquSbkgd2ofiRRaK4CBC9XC
IV+rgjdRAOjPplmeDQMAN4TkYIft9KC/1h8Cj+IfBzd6akLng/YIlvozZo5ecJhT
3sphDXW1e+36K7vYjYo7QgoYC2FOFFJoZsgL+2C5q2lzJu5xEWau5g5G//LjXjX3
i9PBtY4gGpHHFggFrDEeUgC6jk4GNA34wZAmzB5CDKqNVYcyanv5IfkzVxsaG9AM
n/G2EJevmfuXmecVFg5oFDaSm1wK781DPfPwC/khck5kGPuEAzE8x3ncKWm85eio
RjoQAI8HZfpK9kuiCx4TyrW8NRe7UEGMFNJTGoY7WTupr5eDsJ6C9kESu+LM2Iu8
E3A5bzhXQ5OHOI1i3XKmZPdruC2wE5Uz3qlw1KOIvlcJKtcGmhRwCgr0f+EsqPeR
wbJOOa981sVz8oBH9WN2VQYyA5AK9Luybv0m1eWebNtKR17XQamdRpTrGd6c23XF
KWhJCsIRLhh6rYOriC8lTvhAe4Dd1A5I5JXYOgEAK0M3U9y9Ax2OS4TNJzrz77NH
+2Kz09EIMkxu7iHPk5Exqr9WaJic8PBviPhjOtaYYkIue1w/txYoyKACO/IVkGpp
xLI2eYiU4JytAj0ZPBwGAXaFP8i/QUI2KwMBZV3QueSvd19zKwZ8ccjszI5WZ+Z9
yN/OGbb57gCT8hvhOJSrOcwScwT6ZbE2Jb/IBu3e5m24lTkWZHZKSXhLG0U6zeif
ari5MpdE6/Cjr3KhGewfEUsl2x8mm1kYZs1tzp97mhTJhQo0kj5H5iOk/5ZRxsIc
Gz0RzojyljVMCskFLFBIi3LiWxLk6vNa28VcV/Hb8DD8c4osxyU6l8nZ3KvDOqDS
MKvIl88NX4zs+5otDzJ+WKwqDn0tEhk01kyFEOqJf66b6sJXA6yAJ/egvN/508oz
jny7aiLNz/qh4A5bbdusX5FmkbB7X2VyZr2MZ23UglSZjSLT0sbQgSwDkZxdY3VS
f2jbXH/tyMLzaGnGy3fnw8rUSnVG5HRXsTiA4l/sIqBziKOI1Zl3V8aQRDsjRDER
AdxIm1Y9JVXOTfTi2dI5UoCBkrUD6MoHTYAn+R2XgeXdJXhGM2tnOlFXrJLCbZ+c
9517MrJXEz4r27Wh4+TipUnvTm2DuXKYXOI1txKU1KZjH429ucevRCxBWfxK3dje
0CUc8ABfIlQMEa64O3cuS8myazOhvH/433WZBYjSIrQsRLX/rWjWKtPmXrejV0zY
KK+LhuTAxdMPZGE/PAjOAJXTy68zMSseWqd2hPM3ICmaOvPAwgOyPDsno5kSOhTG
BvZa8KLu+Q6HlK9M0GpxhqZIPx8lpVHA8ZFEn2MU6+kZXdjITI5sEEw/tiBkRJ1G
ISFu16AdEukRy4wE18w9qVCnNd/S+XSdDjJi3LvhacOCv6NNvdLCabwX5IG9Q1a+
zcY4PGRdI2ZtEYqG5KULL8HNl/efZ1W0S1DjMqhwyETrVt5H2qN4Z3PJizzkp0s3
R78SeO7jf0PgokcAvGDIyrPp+F7iLlzJ+rUhdB0yvpHBwnD1eSUt1KNoftCjsuea
6ziu/LCTPS4wh2/ipfHMm/kjxSWzPHAeJ4HbTAlFw0+V2IRucz44PqFvwZZSNMqr
m4gRDuddGNiXL+2z2i7TJfEYpAVq9ekamHouDwjXDU38KnIC7pZsyxdy+k8xHAD9
BT2yrKfCCpC6wqKQyw/AvJSHkLISZ2sfXI1hk/W7YUvCV1jpd8NEGQe6krWvWKOR
fnw9axbSSrAMg84h0Fv0eaP/mZhV/1yN3eM04RGuTDjGBqU7T3jy6IHsngzv33Ez
txGXjAHJOnSHMcxMW6ITkfIDSFb0tGwPPP3LLKUXFOb5N+Xfrz08IeyhmWBlgjz1
tNaN9/JXyn3sRiDB2pdVqzWjnn4rB/hMen1sxhCsSb+CKcbwvyoxzFNhJWR4gUTX
J+6AprKX0WD74cuN4AIDAR/b6ETUGCTQF2nufgpYS8SM6+TSZf0YWl/keA18T1JS
daPyGBlc5HCyylz1IEXbuzDy7qXi/ZyLCOeMOVI64z4/7CvBcXbSc8PaP9AtEctf
7pdLxFS3CN0NMtSGuWwj77/tFlZTPQHc2FE4jVXu0JsjtbIg6orxzMt8iE7/CHH7
K/8X6AxdFTqV0BEWmoDRcggcJOKcsXelfTz/b8EuN9uj59XCYEa24aj6BUsQVMMI
hSml0vOn/pcHLNKs3j5vr9uN+QL7MgPlNttqO69ttoKLqrXpMi/243lwMJXaYXRF
sqW7Z3h+wV2Y8iPiL7nBMHtkDD30OyxjhCtVig94Vh17bKd0RQWj9Xdbu8egohn2
ia7b2E8AC0HrCvy8mLrHz7hQ2yXhNKwoYlPBpAkxQwowfiGKa4LJg78ZHpfpwHNW
2HqYezeFOP0/VjYTEeAjAqEJG+NDwoUK1dQD6W7fxgphxqTYytfe2aAPet4XZ9ii
4Gtzu3zrOeWxNt+Ud2E4mHGpgzmdHWZ0i2glWfK04h+oxKIspxUlSjgfoDQcd+3G
NElLgrUQ0qg5Z22Jy2VRZIvkDB7+JE0JO4KS15rWthy7Y30jfhGGDxmrNxqCDf+R
c+NsLTmYoRwKJgiA6zbaBsjXl80juFcoG7osYWE/4ymjnVD0WV9GBJv9uQvI2SCb
Dfv/DMlimKcpHX/l5Vs2Fo0Spclv0diOlAvaw7teVUZYuGidwoCI/R2rec48rJFa
hv1uregiXE99tsqZQ7IdMdXplpzYTHimq/A3qpFLWewV0KPEakIrkECO2L69KReB
QKCLzRmwYh6xoNlO1k2HZiy3+Wmsezh7GZAyDYr0apolJZZvptGGV9MHNG8u66Zn
hek+dqXMBA9RSY3Xy3siddHJKUW9IPD8ZIm0+vzFWhz8duo+V3QfMHgs5aF2LqUx
X/o3rLxlwAzoiq6Qhwlmg+cAB+MNQXAZ82MkM8ryXtcdqZeOb9l1h3LAq/1fje4U
kLwaqktowCba3W2VqBsp5fjXDinN4jshvgeR+gl204bcXw1n5YKl39g6OKuqC7EB
0c+eykVj5XYN73FTEEAtJmVoL7qi1FmXLDzJ5Rs6wxKoGKGIizQ502MpnLck9ux/
ZOJeKAYG1zRytVCD/+RCFWHYLt/S2febgJe8TjP2bv0K7yiNd3+VEvmUkUftp18D
p58Tvtbm0Ljyf7vyqEbq4f/8BAVD/4mQo0WcjjrA/GE3tVFNuKiSqPUA1TET6aWM
2+7McDAvprzO5vdXcfDrrYkyKFbOhKVLBEEXEd6Hj+LQZmopjKORumqziLWfAqz3
1aib2YSvy67RNRLcXY5HWCHQVlaVSPjDSuCEZSk2znbMguoizmsiuMp5mLPv2Zw8
RJlCHDiA68dQOrqC4iUGu1knb0t6sPkt/ihXlfrRDTQGCr0Rso8/gcmgSLJqITIP
6urtfzhU7PKskKGN7cPDte40061Xki9FjeTMBxHhE/euqlmciEwcdyfnEqXm5e1Y
K89pY4cf9DhwCLgYYdgIclthZtsAs/ujfpzB5ri5jDQTNXSvhU3NH6jQf19sg++b
ic2zHBCXHKzmnfeMXd8LAqvx31ycl/m3q36+7kSRYq+rUzkE2NJmUdaEJLQj4fEs
iLtFildpEBzK8F9i6p0Uehh3ubVBuwKB1gQjxfKV78WDLSTj/SLO7+dqYghjwYoR
kdgrKnelA/QxBMYAyGnQ3glvIwJr4UnCGH+oprXAgy+0lZuUaZTt5NB/MHI+6zLy
clM8qgBoEkWRUxlzC+7JZ8Fa1r1rAm9mgXYyuQ8wTxyIX7OQGJyfly8003h7ZotI
5PRP5aLQP9EuHtfSOoL/S+6wr7Q8eVFh9VHmoCofrpjZ+uoSfcojWcb0eG78bqRx
YKew5/HxQkA6ige5U1hCR10AXQ3B+fPfREC9Km3IvPnEUySdfXxpSQm4Lk+4+zAx
A0eJsNPFy+60HlrStxw1S80gJX1KsZQiNjTLaJoEaXaOWjWtLYUzBBVJ+n2s9sVd
1uyA2G15AiEzVT+1emN3hdEs/Vpjsyl+9Zk2IqBgWzAYasDyhfUIjXm+FTCTdq+b
jSpusPV/6LtIK7HCjZqW7/PVaJ5ZSLYvVbAMDOkYQECU2Gp9Qs9aPKOVQrjteKB0
9YOL02jUwPgEzaVUrPgxRoFdToLz7oFk9YVe6xZ+I0wnn01GBh5A8t+rOe7Fi3A/
HAFuoeqY7VCM3rjhIviCDt+UmuuM6DnTHuaNVIKqGg3lWxMyaTWYu4358Seu7tne
WNAg+oKL6no7xryhl2VGC6n9Ru33xe091ze59R5BK9nF60eDzIUz3dIQDPNv4r5l
5PLUhrlgEbrVx2UtC+rgFnRQLUyfNKQEr8w0rMYuJegYylRPLsV+D3WhVYTFKE6j
ZH47+W5dIB/WJ0lxZ9SnriG7CMp+fth2Amm8vcKWS5DNE35cL1RxccUDP7S2wlUT
oW5urY4bEsY5hg8nVQSAic0WyDZ2QmXWYkjZ28KcRslSnc/fO5/sIwdTeywMLGO9
ZKHNOB5pDGHGiyR1LK86mh6D4/WP/l45r66BPw4PlKTp+30gKM8iFuuZ//MfWJR/
l/m9lVUGYQ5y3w678smJI7bUlIcYwd01pOCV6Ll5neXRF6ih1TaVYCSSfwdatSsQ
BvujVWbeejVqa96xsGYw781UYwOXRyDB+rwRE5YFICjr5bVSNLJYX4Q1aVs5oQkZ
9/iBWbhHIxjQ35TwSK/LF52ThLwlZbhbmHNBdC/B2YIIq8ePECLlyCXPPYZSx3+7
uEDqEXlxKyszaSEm1LR2xFcXxVdcK8Q05/50+aI9e8d7TRhY/msXtjDhTOETBB0Y
5DYLP/jMSISNrfEqtHvZAD9MHu29JB3YJiCxyBU2J5R8Q7ldnkBvB/fbR9ipLrl+
IJmRSp+rvt9xM++JpsUJffQLePfFv4+0XL5Jp3duyR8bXFf+z2bE2nvSNO0D+VkA
o+uRDSkP47uLyEe0MKbZY3CgDcgf4ESlMzGFpzgnWvpxgHArg65glWfjgoiLzAgv
uA1Emn0g1/ggJr4jC73tTQVz3dkrUDmjKAMxBizVH/XurDR3xcbQhH5rWa1BcYzC
VGZDJLWIf/gV0MqPh2JOwUFM12Pclgd+0kwVnS2E6GcZsi6i207QKUAW/54NbxE4
zqQdBndLn/fY+TrqVM8alvfK+p/IjJUCQfCQmPT5omchd+FR0r1M6Lz5esDfkrgA
r80hQtXYJrdrysItNkv5EeBlNHz1zBM7FS67lrWUJ50klUlrXWF36OpfD/Esgi6z
FSJfz3aSQpNUT53QmPtamnqMWmidnQM2Lxty/tYso2B0/GLBr2nIMzp8GH34zqfj
2vntlz0ehXh8Wa7xunRxfeiEg/Y9nkd/jqa1PdORa5d9E5M+hIVqe2YLDaUxx1v5
wp1N8/MFm/gM/gmM23mEwy/NdyLbGS1y2WUL25WdNYMEFWUI19orDWKJc1zRIr7w
UF5WXAfFRyf5NSCTTYpmR42uzksavt1X1rrjU6+YRBpvqRCnrha2bZedMXomH8ct
zz2tjEXDHw7VdSN+DswnpCEkRYCtmxKc04iHcp9Fcg39dX1H0OOqC17jiCox6SHB
9Pchst1RgHgrGGNUYMRlF/JJTOVL4ujKWVB1IkayuO1qXWei81KKvyuXmREhVFon
p+/CnKs8MMLFnp9oLrWve+/NIRt3HiwtKNSE/vOEOP3mRPcf7/pevIuXJMG1rj1h
dRMGxof8pYIBJWm256Ajou3Gq7uQmBbgJz2nkLyPFQgf6o7WSpznh2eaLA0GEjQg
oB47jGLlbP9xkJdRtXwmYS5GVlwApVgGSsxUAvt40ZVlKiamblVTWBuY2XtnEnkT
ARBc1YDNsN2WbKnsAEDciCk29r6zq2NYLM0kzzS1SNxPl0RTtqcMKIfCk1ipsT+4
MIev6nQf5zANFhj18ivPlc/DJwNx+ynN94znXhMSaXpsWhgXLFGQcEoHbsVlIpgS
Gjfw/VfU2N9dRCeq9ut7HRCRb2LfmCBHO2LLE2BRlsgFTliHMzAi/kBu9U3DFHYc
ujeOZdZSxxjBQB2wITEFL4/TKBw+SZTUdhalnYVZBZVeREDxgbxxUIjWzU1xGuFl
EWIMKeS6RStdpzWisw/qty8PUkCcVkb8NHP9ZEU3BRxW1YrSNx6vRaBtLW3EpcJm
csfRNoDP7wTQ4FDMpRjvzYGqPHmyvV9RYDs5OovSZdfoze26avuwXe6ig7KtRdHI
FEYePVBEcG7WsX+5UlRS/5w6rNPG5Dgu78x1m2olTGdgKz5vPfAuKi7cQ+XcPQm/
fPBur8BAvC7SSBp91x32IzeW6MukmXdDbhf+fk+hXthFunzlLqieZZJ2pIcbiKch
lQKZpIxkpQdQfOJuiqD4XIpia2ozTUhTkli/QMPz4PxseM3fsQ5VtGiKBOU0u3VI
HguqXD0ZfrFeTv0IThviRe7Ffbxt2evEfa7kk7kLGa0cCfUUQOoZz3msYD8Gl7OC
lq+CdjIsPV8E9q/1MX6qxFcn1Dt+zmcJtcoaOv/jho0EXLjLZiQuvxCuqaW8RayI
ngu6YBk7qUS4AEjF8x4lWow/3sliertM0shrXo1M7eYy5LR/Hatgebbli0CBPBtk
J/WJFA6v0OfC1U1QHpOweCOQUCUvVZAPzmzucd+KH9McmXzaQuwqZfyH5OY2jGvg
j3l7WyUTiyiFQJ3kuGhxMMAtCoBNE1dnewenTzWr4bFuwf+AT7aToj408L8NOnEZ
tBq80hkc2MdMS+etRKPUkH6oYz24q0NVr5FUGwG9h/Is/5VhSwPugEbT/I+b90V1
gUvjdbPQIH7oRw4V4aOd38FDwJE0KesGyHp2RsotFPVAVaJTivD996PuaqADfHDZ
FIWe/R/kQ0cl5w50B4k1OXVc8uWY46dqn6kwnAoDBvTP4GUplQnk5Xvvg3lVxWXv
JlummIAeuAZI9qyqDvdfurOWNVyzELdzyImt0lB/6314ZDQNfeaoPr+kdaX7tyZN
yvkfZ6jZCfpwtRI+ZD1GfDT6aHjlNcRnjQJ4EdnQTZW5t8YrW9ATPOHUHw8Yscxi
5A2pwmAZAfw9xEHIGatPNxGIaRGprHEkqg+RW1+e7zI0G5Il+lbXzcQqOCoZYDNG
/Hq2KIt/ONZ3+1l2dyJRjnLvjxLgUr56NtXp0nrl1kw5PWnvgPOxYs/DaQb8C7fM
6QOv+FthmTrvWB1X2siHUCkDlRUVzJgIJa9uVwX/dRkyozwKJ95LPpxVAVYhekoO
9PwMortZOiCnt8q/iSLoctJ00QAyJgI7f2RO96+4ilNqMVokT2jUOCKgatc1wEDR
WQcTBZVfYeddpjleCS4TqIYYcnISkOMCvE0C3zQYOTHYrGinByQ8ZrBRHHnyuta9
FxxWrrgpWVuQrS7BJQUMfDvbf3/DGCPGJR9LBleBeSUPzSCeWFgDE8sN2gxWIuxb
Enbd7oG2RkuHNvPmBi9S99Fw7F5Y50RFX5NsqqdZldyNUlcnY86xviKMUJNSis/7
QuN/KlrJH/p5GV3bFgFKJD969Z8hwlHtTZtKDwTfMnJaw9X1YoFlzdSHHgIhvAs5
2SnNRStl9BwPvAsqEHIlGP07A9VLwOxrNGYzs5zAq2TQIrfjbSNau8ZZbKQFogBn
lbjaFMaVGtcib9bD4VmyOdKAOrddtIH4J8u8ElXhxtZTysNIfc2P+uJB/KaY+98M
4RjK+A42PcAVISpf4M9E6xYQH5wXCnbBqkVlgvgj/15biv3FhjOT9aWMBmGnqxry
XWbm4JvGT6/ddIWwHjAnFhYzs7sZkVRvBXaM32T+c6zGgzeUxssOt5hPNALEQnXn
EV+TEEZJ3R73VuG2mh6iGstX+ODmEfd5e50Us5dccMTHGqOpcK899DkA0veiX3Vc
aldivBapWTXYwVs8vikgf9UI8Ihu6ZzIxeCnZVrMo20l4sP1FMqbZ8krdE4yEBI+
k4XyNHXcHLpvi9Bkw1mLF9HVFyE3dhLzXDKfodx6Gy0pcQelyIt8MM8NYzkTLX2X
Qv6cEdT5mSYqkdjP8hI3MVBgWoC0sXMwqtnfXHGr3RLFjrOgaKhn7RNfVeRW0E9d
Hgp8e1xB0AgLuS+LG93WVIUVC+bsQx+gJIp4bST2IRqgh5l5dWBrk0NEhMUX+GQu
DtwnUlJQdf79EJFw7gGw2eBJ7XqmZ55+MB5QwWr3OZC8BCggxZS4e/S4mCM3Ksff
7IH+6tsL7b61v8rN50z+JcPaY9BXGyFjBvZ8Ze+2cDiz9nr3MIuv9vvJ2JKnRBAO
YTQu9+iEQ/LfeAVcet7byOkxQrD80oAgdwIc9kWDJeCReRwXBXtI239e4t3yDL2w
s3oUXPHgGG3SIbHcpaHyMfKWBDqBcrTxfBGVef6zm8r4Nic4oNs/oej1R4hIG44Q
FM0iVownUUwAFVYRgAhl/RW58amzqviUA4siMyAa5CxG3L6lLbxaYpE4HBfAu/qF
Ax7WFV/wHirexFYxH1KdQs9GZ8A5EkTZ402BLXZR+9mGcO8D7x/vHtPv+87e1UYr
hq1pwVHuh+4V6L+iIs/6qjjjSZ+PzXYzGbfzHpe70P6r8kM66BnIHEMt5LDLiTvO
BgyNSAXgM2Rwft6j94SJ0OTeBdVnFwlkD193X1zGu8681I/5tG+VZP4rTbgbMoAC
5I3BI26owBleEeAlFHREo03dPfDTkYm1EVBvpn+/bTUv3HTY+Eq9+R24MKm+di4x
tZbrjWrjX33b5H9+DdYFUwKgE1Yx4EuuUf7zOlkQaFEDxwM1xk+bQMNnM3G7kDk/
tzepNu+dRFNNhDWtE3mvAAL2/PNDRnHXuUfSTZCowtknmbHfRJFoikx57sOpLqeb
b/9+vl506Rhp41k5MUMou61nfeiCFZozy+G1W9k+V9TIvM3ZDD7hRbzFtDkP+L5a
0Kx1GjmGKlKUuPbvqSvCI2zx3oeis8RWXitXbwiA5Kh4qNSN8k3nHv9oIg5UBr2a
zTf07BG6jOomrCc4aVlN6tfHUeu0wnHilqdKy35O7Iesqwffs2JdH/KnhADIp3iL
z8h/IF9P/VM5lVOBuWdVh6rFGI6JnzFYiYNdamtlrEgW7jIddY7Bwy54qo94t+IZ
Jwm1ZjSIaaruz4mTFNVqKwwPrYwfDMipJWEGYik48sKEStxzxKiS2pxSVDO8TySx
VUHm9RzFKv7+txSQspnWV2mMoqjp6QWRlOmiOWURVtFa7uSfwFPk1pT5MxboEYBQ
pnci8RRmcySmGZNnEO0HBavr545Qhyigdt4Y2EuCRpX4gt3/lu2DsvqVpdGdH6g0
N/jxNmlxOOl/bFW0ZpS215hcTk7Ub7qSMt5a79oUn6/hC1Mq+PxHDimnZ/pS2/eU
DCbUMdHigZ0mryYPoKuILVOPf1Ucyt+6dWI37fPD2dHDmQAXhI2azaCDNOfS8pg6
Tr5Z/ES5YG6b04nlAIy1JKjcH/Sjh6f7eP3/X8SjE+YayM3TYImQ3HwBugZAWpp5
NcuwwU1Hh6PeXsKW5y8D5TO9QGe1k76Sun2dJ4tjHg69ykKaNC5EfCqaHwjCW4eV
P9W1QGZWc+044PzVsPBN7ZwXHT1v+h/tyoFluMqV6VZJo4YPyxPFc6n2zgXxyyaG
x+6Y5CHbJ2/pgV3w6bGHG11JIubf6zNtbX0oHJdngQ55oAEpkUyX2FLuYLC/2Yga
7AQ1k5Fux9b2183A/An/DM8Vma8MQfBpfuOU9BND4m6FpPIIXx4M/JQFvPKpNqrx
0tTyLkaOpuePxRJxWYWKYWXIImAEwEsEqt3GfGeZzClZUukHoRa9z61BxEScnWHj
J1LmUePNfGH8z27mbwQeF3nwS1XRz/Sr9CITH63GJVwTVcw/aQXJw2nPNNJZtFSW
X7/DYnK/vfjquwjivy81yDraGvn4GQdk0LUVXfA2pEVs169iuQqiPWqNfL1vC0gq
WRC5D9Q/qygpddISyOntzGfE6qJ8f8MWtZ7HDjiHjLQINfa0/FT1D0FvNWHxshXU
D/R8SH4Ke2dMYHLq4OA7I2rlFaW65T3DFootmho0LuHTp6fi1L2/UpgmNA0+MEZE
WwAp5Mm0xqqDm0IaoFwRiEPKvs2+qYYKAk4hUvorrG+eEDETwmhBDw5/udoqIFhA
SH+st7Wk/VqkXCBstK0Kw2atG+TUc3fGjAIzUUupEBYfxFBfJtbIvdBK3qktDEka
bEzHYpWjFmZM73kejlZLhoMXNM75T6CLSpzMRu2nJj9vOP8omM80DdnGl/scdMLA
Odl4UcqbVvOjYxInBjkQyW9cPeEFGtVJK6wCAVXZzdhpIIpJAgfXoBenp9QS5qvJ
wjHLFGx+gKYZvfpDzLYb6fiyvpYgnRYDSAMXmG4+Bkj9QuDdkm1U8kcum3wLBOys
TlN/hGjsYIYvy+RoE/BsQK+U1JuAQPOFS295X7EfHce/pNzvj9g8uMFQZb2c9CeA
33nkqRIOXt0jNHVe6OCZmxtYd5wuiKJWx7bYwulTzte5HOVFZz+seyTJ+U6FAyDh
tMrZxi3OR431Pj35acZ+XT6JQkCBNxnZ8t3Tz47qCOtufMq4paGzvAmMo4fxI8O9
wiApS5OtWuAxkLOtRFIJuYYPoBYychZHFmK7RrH78Ohjv+Tnc+yXJOVi/sroFrjM
WF/Q/eVlJ0pqGkHxfCSCPEEly8a0RVpLEiOlMryerW9vyhc7d0bMZZIKy0HEDIrR
WvIawfNiw2+j5PGx+Wp+ENuIkhau3vksMOLu8INtOofr9qNMV1GyOO1MEJeSl/Nf
0u8foctLwy/CImdQytUzpuSXSio711hS7gA9pAByrH9F/NJe3/N+Fo5o9ZQlGjUO
l662F04oJoFQdX5syqByqzl2Io2/oYfWsp2n9N4Va0nlFTkDEHgrEMgj5EJJquzA
AXk1rBT7J4EpRB3JIol7NIQDR8WJzYYeE2PjCRXF9dq1yaC3r21D1y2VGayVDdKm
Y/MIjNdx4a63H72AMxvIDU7JaE9+d0JoGRgPYozH8Pz/GFYI7xS0tInt49oGxI/k
e2lppzofcbu/Bn97p6M6YVyZqp5xZJvs3OM5hFn2xKsfCtENTLE4v8yeHA3NSZSn
dEZ2lM6BAc/bjwl5zdxuuRn//smgOxk2NXle1mtSd2eU3N1yLd679VZ1qy5l0qK7
E3qgyMODBl9Qh/f/27arS1JEOU76lgGjmkxVGfZ+NfmqBrhVQDpp//s7waZZOmL2
tbLsGMhpK6V5GxnVvmnzSOtjG5sABqLYUfA0CuI9gEA7cJKE1v3XOcs93lBiHnVu
fUdYmwkH2ZzmnNOTWCqgoXSpILeS0ZRBQ+8Mva/4xoqw8883CvBOvpoowAhMwkXO
MVDa845GrCzLxurEU0LLoFQEccQ4a9gMH5THb/w/nERp1MJBBc+JYH/nBg8SWrMM
6qkmMao0+6o8/5DX9ts1RezAdliuB1aJGnZharEmVXc/V0Z7xxlefM8a9x2I/0Q8
oZYe5ev/yX3CxeSn6s3DNWNzd/jOCsq58TdVKac/xSnfxRlTOHRvCkD2HJU1yCAu
aTkdUyn/oxcmBaQIED1GXg+9Hs+liQkDVGv/gjGkDZKx+oVgs6d2TJm0cuhFRlCk
EBRLBfAASDNn+zi4WGNDYLC1hYinZCdu1b6UB2CF0XW4nfLXnSeJv+1Y0wufviK3
VkplyRsfSX84EqazarWZXky6uVcURSBXQUYsGcT+vAotH8oKMt+p4WrW2lBgeQ5q
U923xq8PJP6cDe81YwTtsNFq45r+kiqNHt+y3kCvWQWE+UT2UBb+J3hPWFe66j/W
j9gzEhJ9Hn5egltsEtgBILzf64Il3xHSj2XvS3Te/NDEy7IhmVFRaoUvuOEqO75Q
0JmEMpNx2gYgfHMje4MNaAo5vlsS04NAzWBAu42MM9yacH+wTrxWVaXJCtf/8qXp
33eiSxLOC78kZ8EGyI8E4V5JQhRFTtzu7jnmWVBa7wc4NK0tY3lXxNTaPl7t4cvU
9c9XpHvOYCS94AfB3yhBI9IogPRX395Ud5kIvTpo3NRpGeO/Maxs5XxxK9Me0iZa
FlHdKETtJeto7UflPbRIO0GxmMinms8vOVe72L6oRa6aB9Gcn+SfSN60/fOFdmOL
qFslVr+JjpwnpsxsN9pzhAcHERFk14kvDom09sLQbSN6SAKUR+e7Ww+b/qTSGRTC
AcJPrmzv7D+oDfHLjDHBAhqtGEh1D47+/JjgTIlSBKwKNBgpRshQE3uNwGaR/+8z
CkmGh8xOfRC2uEYGmB5yKNkXG9dkeNV88/DTvHlCqsuM+/kvctT0prAjA3ehkJvT
jsXAm2q8BvbxqXcrVGcgJZQ/6TLNyF5pptFGW943L8qvfl2VLy8j2YATzVMebKAb
htxOwbiBMraxtOj+2a59QpnZPbR0eBK61MYlH+LemGmpvum+84X4ahe5rcJpj50P
8EnCp/7vMaif1u61m9pGSjycQjjhKZMkgYR2vy0QeOVfz0lJYDZFJ48IVtYsPToz
cf8QVWGromKuvmPB3eWjzU4y+avT3H3VD6tA9j70kejvi55RAkuv49DANEmUkRrQ
Jy4ZWNdjN9GuBkLFWMz5ukyk32eKleXEDgfZ8awnqHho7G6YHMowgD0qt4Jb8Qfm
45UgIlKouDKfadGrupIdsfT5ae4Y0dcrmeoJxcLCYqJOFifES0k5ASvEvp5oqhdK
4G5BQaEXHnDwk86aCilOAAbQJT84KnrNJ0+7IqaJ/cP4huc/8JyP63Bs3Hm8u8Z9
HS6ohIoyyFB4lJCNZBVbhf2JFyhjRW6X41kcvq3/lpqDdzrl6n0GZdxopDp9m61W
xw3lUUFy154/CtLePvoeoGCSAuhfD0pbAMmCB72XruxrQuGuQFgZuT6Bp5iQYZsv
jzXZWYGMsWRXPcljyJ1YIxmFcE2SvZMDOUJ5VBy6Im8H7jPhgeD/3VGIcn7YfqWt
jVPOo6/tRqNFwr/wZ8y0nBL4jYDb81LQslwsy/GFnvx8tiSWJIFKwr/NLSBhreeZ
ME9eeguHHyKBXmPt48FOPTmqkyta19buIgkZwkKofT48dWUyL/9sWfLSgIPehHDe
E4kzSwxdMvR6LdpnGrfscNipNXTPZa3u4/+RhgWX4B0YGMJOITc7oGuPSaadaFuq
VHwWLqOUyTICtaejox4cZWV+lVYyRQGhiWjC80YBb5vhDmBoqaW5Ui4WtBfa6hFL
ZReXqdE8epO1UxPt8kZn0gB1VqU+zFvWAac/xi1KIW2pzvqU7HooVVtlV49ngP67
DzkaPo6D+iYbh3vcK2UP525MbTe6p1A30LxuHskgQ0KnJIrhPuJixdY3t85OCjXv
M4E801WhBDaRfJoqGkfaZh7QDErPZYtFwvrG6j9zb8fYy5AbU48JLON9fY3uyDH8
X0ivG+pgWfrb/8ZKpvM+zxmQF9/kVhJAKcP8ZwuFIhGB3xbQCCDxZBOw9frp82Zc
bpAF/3zAHyT1yjgCNt2O86Bt4jtcOuvnEQm2DLDI3c84IjddmM4IZZHpLp1hiw3n
VGQTs09vB5ZSCfn0UdqFSLYnHzf9FvG/5FaiIlv4LFNMAkoiix5rSg5xensDVWR2
l/Qfry2aeRF3F+JT2qIRREzi8CsZ2J+HW7LurEhh/jyAwCRMu4Q7qKblcfzPeJQf
kb1VZ/H9h50uMEZaHyHKBIPwsqNBtZnphU2vsHT9jVay9+V/jGB31BnUIYYtG7gS
ISrF+kVaZDBsSHR35KfWquk210ao68g1YQckWX3AidF0DG0I5/vwDGHEmUPThiHi
Mnrl1x8mpZzfoz/x1dQ96VTQj4hPzHHzO5E5tAB+WfgJxeisxp29QcUUlEMBUAby
jGdDMcxDAc+NemCS1+Ty4j+VBL/1MhfRsDY1s9rCKwXpVqIFLni8wyNZ6KmEC0NL
6+p8QIfFpXR4fAtt3d/C6vpwfGjoEcNA+MW111IhRejVALYDPHQdXNcoPjS1+Oh0
kGgFA9ZwdqZJ4d5q58zkLiRDO52oNG384vsRC4mD58jlK/bZAew4PvIeZxdKGt4n
hrnEYAwpqRppBlCevF/GdW+3fmPRVspFzk2L2xbML/+BikVkkj5deSh+KW5Y0SBW
MIlW99XlxuS7tcAXOZxYEqxZdR5BYY57D5N6S1ldO5lS2rRiG6F/0rkPg50TwOFG
VoPXWC60LNtnwpTXUsU26LjXlngnd5zrNp3UAhq9GR4qVAOoo+qtKGBu5Ku3PdZ9
ZC2FqtV73xRgr65sjCGKH1FBepPlZZXJNY5TflE8lZw04yYzYC7pRCEg3y40nJcW
br8+ApW7Pehj7HWyQYo/A0yumwTe8GWg3Lhbm1ydWPLxRAp+V5vBTNAcS+NN2myA
Id74Ap/0cZPR4nzhecDp3xi1K7qgjAtcKTIssvBGs2t4Z7F9bXxd5kwD25cJ/yqa
Md6nleZEWLtgO44sI+zv/TR/drUoHptJhrFmf7fXk+AgJtZPwHBGKa8PiVV8FqBe
DV+f30Kzt8dJByXns/FPUokN47Bhhk2cKm0sYQVsyKl3gGa/MJtx7nF17TltKsOB
E/JLNT2zrWDmzECrScO81+hOwWnOastsw1+gMKdyPQk3yhpeThQ8XL6XgI1lrJu1
qHpRatQ8yKe+14TRA+SMQ6pbkUWL7nAtisJoYinDzlDsUXgE5DLtN48BS6zxaB7n
vkFPXj/ipVVNpO7IZofJ8Vq1X5cetMPYRre3or5XW06y/KinpLrNuBjY3otTM5Pv
+3ysM7kmE/qLVrYv0tWoC365dgZ+brmojeOCdU0zN7jE82DVWEhjk6w7kxnasg1M
8DglGASyzFPngXd9RlA7dsf9gJsfZQCmVRgj/1sfghjjpCJ8PpaDjtEy6xscuQx/
7rLvGvvy2tSQRLMM4ZTbBKKEkJ8VKMxf0DqL/HFu8Hhft3icfqW+LoPzGeT28Bcx
tNUT1opCPNya4q5Mr4TFtzTmTDocg+4SQR9yDzv2VE3239bQ4cTRyFYPXitswBvX
MojA4eFhrOSVQdIutK0PmuhisXbJRHsO7FdQZQQVGU5mkg0/jmigo2BMvLNZqFYD
dYVJD3ANaXR1qOU09paVmZCqP2YghS0FC7JtWwVWBvsg+znrEDisMEGjhzaVNwAQ
Nh9s4eOuUYvY/+pa4+pMTAYq0Sa9Dp4jxjPEv/+EFjzNNnQweL6pdEpnQHV6I/Cw
X7vw+LXDV7iC7pjfXUkkTUDb8nrxzz89nyAHMuEGAq49roD8Uqz9f7uUdoSn1LAp
y3O6UQ7sZjUhQ7UCoy/Cr4RaWHR8A6AkxwYL6x44Z7bKAUsYe/uZD1aZI3dy423X
SqzX8FJiovLhlPFFWmHATNNmvkOytC4YpCzxa5f3yCekls8W3QPUTB34TyLgmSzJ
LaLpbqIO0TmTDqWtP3nq78A6D4wFM1xQL9UM+E9l+ZOajURtm7AtaTRDoXgI0gsq
hczUHdTOaLBocf1lRybBjn/JE32SsXEJyX6XIlgCbFgHV+9sZZXpv0eRawB5+8E1
whIfhyl1TOxnA76DhXFktkdWbP40RQFbJNfB6ZGeA5QU+OrwFsao4y2v+4ptIgx4
nPN0IhEATjVoLxc3m8wV/UHSF7csYhAk2gIjfbCJyw+ZvEzNP/AbESn1NCwMYkG9
GoIDJQItcdqMLK56UkLE9EMiPxD4EJ7R4SFmkSRqn/v5A+cDRsZBPfVa784ku6kx
ZSGhT1p4rMZWUsKOtB1p1FYYJxVV7nPU5Sq6Gfknc/w7+GViD3sLDWJkRvyhynLa
tTn3kyl7wEil6y+lQGbYpDqlvc038gFz951LC82aIaAXn0lTEEup5VyLItrI+Jpt
wCXv2gwm2Vecnhggdq8D6OOkKkDri+RypmmsIluY/lL4a4P7xVdPJSdjq3yllByw
l94xR3LbBK+LfYSaGjpl2wu68MSpO5W1aloTD4HAPoM0KM5++GjF2UEBv5cJM3kE
XwLmuds2SL+/ohrI9vpI9nAoIqZWY2KoenpXV3QRrAO1hurQOBLMZfcv17A2GUGJ
3N+Hpozvj7PkoHg3z7qd05AIs5N8Bv19JA8N3WoNG9GaX7JbJ6Ith5H0OjAo01Cq
Imben8k0Ysw+4BcWoNEW+tbf2TfRWqP+4trFr7kMHQ3WKi6VCC9sDwI+z+44ndkP
XLYUVo9t9/rf5PkmrYRwyiaET42Eq9XLSVmJHt7+W1ACr9NBoCpuAWUm0N44p4xO
ecrB0RgG0uk03HoPBo7u/o5zvhLlsfceLVe+2Xh5VlQBK7bR8AhtsJojUYNyYjrv
U+H3Iu+aq+d1PAfVfXZBMaX5XK6gL0GrRtO94dXXhLMJ7dMeiS0IKlJr/Ho2vHPa
Ulxev+sOHIR4kgevJMNMpqRZ4OFuoK4ADRUAMjmYyQE/Ifor3d8hiWDddJU7Bv8A
ls4MFiS4yEWFRMbkhmp2RFe20gGxyysrTgREvlzDSgV3F2c6M6uXVygJXswxT/nD
ZGY3lVkrz0sGt2A19ea4ERfJbHPouE9t8+I4d/0ve3kKJ+mm4ufZEz/83WQzOjB/
jEvS0LxMdjrhtLa7dE3zAWSc0AqOL7KcZlFBKShowEknc1y72GmSqVeocMMuH8LS
n08ilGFqlv3Ma23IQzTb4jTX/FKnpyVtJC2BW6l4jfopLQ4eNbgOFUbN0Ewufpoi
HTvtsbl51xwWJqn0NjxKAySy8edIaMu/NtQJT18ek6IqsR8VC/YyouHOWfmrgM/K
ig1Wzc5hCRv3OyHfGxwt7FMm2UlpjuaJK7mIr3cuC2mt5q/Lclf3ojgrbZAbQm3H
qpXsa1c0I8yRxhevJo+ef9F1VN/XP1xy6Z2w8z8dQcElwDlRlBwYhdNOXBF0Oga3
3PHMCAw0MPYMjQNoKyHLUe7/MYewyHHYi5yhiz62qh3RSIUi//1IPAQR24VZHRz5
N45TGBlNzVe34g4lqRA7pOUnqMvj9v+H9gehOlNqCUZTnplwxY8S6JY9JI5vNI/J
RTsTbmE7Ei69j+DI+QJFZDa+35gXM1kGsXCOaxv5QHXQSkSeOuxqP03LQ+XXVRpa
McHTGaLWyx9PM86RtEADVrhyZUP64TwR6juCHAWwb9/BlCA2mxeHhPnODIi+GtGK
xt+ejS/JwhQ/YmHGqJBFFNC//n0Lj5NqISvdcIHVHIxqZD0Jcwr0fBu79NtCMMpA
C3RYfB9FlDb70lPpK3Dih1N66Ojh6jaL6pzHzzLJUo1zJVMrnocotFTQ6THUdZi0
EculrhVL6OHZxP1r2JgrWrguw00Wnd3b15q6815JMQra9umJ57T0OsgSQmUwx/G5
e2sdL0MVF2pxnvheWwpL4DiGxy9t9n8FdCHoiYh7X4nQlL/k3k+THWy/Wz7b/G5n
+4tGsBcxfNzzupkKvDa2Y5HLZYZEZA+HNUQSCxAb9onhlkr4QDgwBuE8OJ6XS/vg
3bH6MZh5+46S9aQF1Pye+QQYzKMbAfTqx/1K3dbFd2YY5ruc4r6w8vqnM+/dc7up
T/DcmOrHN6Vbw6bmNcL6Bjg4umannuGZou2exQfrNqz4xiOANGhyeknIv6/qHRKt
VyMQhISka6jRaxJPJWXEsaQEGw5jJO13oRice+fU+cEirZixK1DFeLSWhAK9xSOF
zGcuBrH7e1AGosgknQbk9tMvdShgZ2BOeznVkodsOJh+ZZRhFyl2OvXGy7z4WylT
K/Oo8vc/v0wJxcCdlyOrRcEoweuy0cuyD2kN6kWpa+XChKIXDnGPX1nBFxBKZw1x
ab7pyq3KOWNxWSMZcGbqiUJLpf3LZ27oQzQ0cRQdccu41LcYU8eudw5nFlVZEvuS
/WGp3Gb9o6pw6NwsmX4BDP2vMliBnw0ydgzCb3dlbg7ak19wCPA8HBCNs0JCRLrM
8JsqM/cFgKThZoqyXisasl/qJJ855M9suCMyBdTL4wG6KTevJaxHA5ZuTl+MOgGw
fHYIGKKFPneL4tg2AxBb7hwmn9cCK6B664Xwu1lYJyY0oJJMISgMcQHhva8qDVwV
bMDQyxl7W+nIVPDDuxb5fHVQX84YfzvA1qopZB6d1/b8+JcsNzNA2Zowt46Dxihp
lB4oDsjXGnjkbh9z+aZMNGseTBMVeUjWZjZPhrJedJcCP0MozlUa1m7tVGk52pgZ
IwSovkcaXtOIB1vPMVh+EBVpIoUNydHvGli3+w7qGnTmpj/8KICPhPxuffZy6UC9
wf4apaWntMqqzLG3o50/68V3vp1rQZ0ucysMCCUg8q6rcuX3uUc07HQBvWLQ1rit
456GW/7rLdI6iIdNkTF+7VpsFpedF7xGDfVnpEMPJyog7Z+pH1rSkOyJWYnafB8Y
+Un8iRz62I52P6bRVO4K51mkThSDhdDuf2vyoUtPsEWZaIfdvHHxCoM3of5mwGNV
4ZmRWmvNDLqqfebATHWwcUO3yzVVwB5+/WIZvl+ptCsNr79/fzcvO5OFnvAQ/TVP
7InZHC3meDQzFUkrup/YZEgvp54h7uDYC4NmHSYAi4tk0VqusI7hzfsrM5tHOQof
jKOeMyEem+AwdJJ2iUgEK0qqXQl/vrx4+/P4cU0nJpZ8NJ65GexhZkPTzqKtJtpm
/VZJWb5EV14UpSNhhKsrexch7TBosolg9TY+Gb6i/NbMpXNeEy4ksxMWim5/UK4F
RJ/kko7OB6PgVRJGsphSMLdZ1wRbt7MCe2I3uA40NZE2a4mDiftOeHD0qySRW8e0
UeHr5GJxwg25antZzwa3FPPExQnIPlLkzzEi2yDXqlPtlWmvKTnpUTL3XAkhR62t
Mhir04Rm0IGEintSOvB1evYrv0tqDm6bIQtJkndCJO+XUGoslJrmgS3GcjHKyU9f
aupPalTkJNLfcqXhVldzlrTWfB6oZUXBoTP8p0BbvOQ3x2ux0X1ThONndnhf2l1k
bPlOnZoOPVsDTv1Mt6rJBmknMPXzhfAHUSrcwjxDmI1rm/Bo2JvI2mdW0RmVr11r
KkVK2xawE7xiCHQ608mevT1rl4Cy1EpVmjY/vtFgMtl7conYtC68QRZsDMpyISgS
63np2hwIYaqVNOjI6jz4ixptSVs7M1omB/U7CDqZ+q2flTlAqH87ebYIxl9T43zZ
zX3JUe5qls4z8ze7x3Qh4K2f0OtH10QrAux2+y5+YESpA8fIUNbrEvH3bkB9R4Xg
Xuzptk/V3MCcQYrIzUO6F+HtYwFngEkwx4HjjHqHCPnMVz2gMSpRhhM/Hl4oxJsm
gTUG7dWfrv6HqOoUzGI6T5vxfYelcpaYJ7yPypPY1ahNu2r5mSsbqyVUlkJ+9Y7K
MxhNqf3yEwzHljN59RzsD9Q9d0KVsZHOdkN++ieVbs092mI8XLq0H1EVnGm9WBPY
wS7VtvZrBFK6Rrr5WE9ibmrul835lEblicju/zc6lDdmnTmcy7hdj5H5UYwMi/mM
g8FVQYmZQV9HoX/w75Wea3xswbNvfyC7XCG9zICBsOctauaHnUXpyq4rxnaR+YSP
Gm7rKfZDrlLkExSb0qy/YV/1afsk4P7eaVlNG+wirq3qBuDUsJlpihtCqOwXbllH
ThGj3g1Dy+MyXxJXowjdCgIWvEU/BM3GdAYHx4LYs4RUzlPObU9d0daETjB22Tvw
pgsUnvQze4lR6+IYbCul0iPBzgHOppEr22Nxw8EE7SnMTyWu7lVvJyHk5k9CFOUm
5gMYgsePEguRL+YbBzZVUBMywqWjMQkY8yYknYNRcX4g5Yq/8yT3I9bwyiv4MRSa
OGL+vXjgl48ayyXgA47f0fbDsqu1XwvIKffcfGyWhUN3qWM3rY3x/Sd8gU+xt9AL
Gp+DJhr8kIOEyXNz98Jc3crDFtaVQrXNwaAlaQD9skvMU2JyGhWE0/o/3XgdQNGU
7dnHCXQRGnBaxpdcL2qfFKB21OjxcqHelX/0tLMnT1LzXGdqsA05T3dCTh+L+diK
RJXWG1VObuW33roV0EynI+XtdDEP72D+5ZamMf767DMrlS+x/uFnr89lazzm8d/S
K3jzfb0FESQi9psrA80GxCwK0V0w31/BBt7vQCGOu80+CWjD2EwcLqRmmM3vaYLc
Mb+e41QBBEw7op5wiLET5lrYG99QZ/Jn8RQeRHcQsj87Y8a8AK7u2AIzp7bdPzH6
/su7XlO9FzoZOJPAOsbg2rA0Bp8KzluZBeM2Az6qVYjx7NRHmlJ4o+C5msusCA02
3gdp/8IccbctrNXKFxJRhZ4YlGWaOpcFPmT/pPU7q4OKE+ukD8gaGTiqGuaK3HBh
bGjMg0rb8oHcsj9Q6FVzmm8gm5VKB8OgmHP69y6jDnQ+IdZVapgNlIUCHDwbPuGc
Ztt5IBvxcKe79iOk4f7lcFaAFKuWjDTOFQSXWUJP0bUzyAKtPMHZufBpvIW5NqxY
xLSEHYjk/ZjHIN3mQoAtVQ9qct0e0S33OfA5heq3Nl39UlluXEC/WLkwpprqo5lt
XWRETp5Ce4wf6cV4xSm7mDlix/Tw4eU+Q19cw49539pdlRq+ze/5cPbM7Iwqj0RY
geo3+aKRe1BISX8z42C21bTSvdTnAjyBAGYQg888vwkDmQwL2RibV8Mvp6bceJ5k
n+52fFrtovc3F80HuqucY0q8mBuaxkiWoO23MZ0aaM8iwCok8qv9JxibOcx6FsvK
S9/fUQ/aubQaaZyCquSuYDhfkHYsVOfflQRsyfPMfb6KbQ8FJEI2zcJrN8ordHxk
SD7TZBLHMKrzBusvmZA5SJRS0d7gk8T9ZhcFWYW8Y4fWFm9053rB+9Q4ZE+EAtNr
/w9oIIbK9x0gmNWx1hjfj8npq2dVmWmB0HiqlY+4Hc1UyJ6o24hlpUhqGLkleDs8
wnlPA3RnN7yCd26+f0owBWyuWo56ecl2PHaSb6dcZDyzkq8uHDB8LmvhlN60ituo
Jmm5eyecF/1BbVDEwZtUCLTz9q8NJD9YvovK5ChnE2bIWwC3NABSrAUQvrl6cOgG
0LfoE7IAn2X1IwkKe0Rp4uakEHv40ntT4nmAtGbTxfcskOavJTDzP1013wZ38j+J
RHkZEyBzZFhefo26pyOvIPqR7QxA7sdPfZvjF8LUFXy2aVRtrPCxxOzQNlWXEc1v
koxWkiS0CrlrSOf0Qt6y6WZyuDsjTvyMGEu/iiqPoQf19tQmnMzt0DCl2eXHTptG
uyCPVSLBzOKDiJJ4MyPwvG6Tkl7ne4hjaiog5wRbIQXbjWaF0+MeuagTNVvsLXJO
NjsI1dX6lJTMjVPG/t3WZQ7V3iP1/I1HF0DnisVez1M1n2eWu748G5j6b9LznrHf
eu6/ZlbT6AJJkYvUhPatCk3ZnLwiDlEXSBaUJ8lU8CY2Yj2qwmCyA4MpMZQtDXAq
ff1GIUULxF9aTH9kwlJM1ahLK78tjgY8ixE4MgOt1p4EaK+b2ZCYqhol5D0zG6su
0TgSo9tnfc62J2Lq2QE5ghg9CGa5WPbmgn9NpXDwxpktzuXEh9GbxJFCtHW1YcXi
dYdgySWNrmeIiit/PZ93OD7gSaxI6fY/ZEwLYbwMrHA5idSClSSRf+h8tjWSJ/AP
R66sVNjnjVRHL4/RrakEDSaEDkpMdflTSjCnCMIcQ2jTcUAc0M08mHEa1gLAfpQN
dVdrlUSLZGri8a3g8b+p6/BijghcLqHdbS2tlOqfQfmQn2cNIzaEgqDIvvahs11P
kIxK8pIAyeKCilzACtd9WHrO/jUA2XK+P+sXMcVEF44Rl1GZUYWZVl4i3KlXDJT7
t74AQ1TD9hpV0JF7Nd32Lz6YrJF4JKJCVHjyi9eKRne8334Z7iG1Torjhzbl7pX7
APG0TyshOC0y6cXg6/znqVQdEK2DB1hoiZfejFuJAMaGe+X5rvzGN66m4EiWZeNO
hK7HUrcoX7y9/1gyqicSX5KE+HNr3GxwkTF3s3O9fcl0cDcP7NSQhLzFyYEWx1sx
7GNzJpxvCOY7C0NlNcFFen1aqidWSqTR3jiPZeBJysOC4Z/Dhnk6rgdEyb1yD4UH
BU8L27LzcHC/CfxssWBAGlbrIrLyjrsQa50jdezJodC8JGWK9YGkS9v8JQsjvNDj
ChYEPevaz5ph21pbY5vXtaKvdAJDkcOdLHpmWveHEJIz5PSgfAo7dGDNiMgt+kgY
6Lb4/Zrz72lNK0ZuszF+JSkpv+idgmZSP2G8+5Cns9LA2mUctno+NXWtposIbXO3
jEDFXOM2qisFXo36YkJqyaajZQDA3fPXv10YnSFt+/HpojH1QBMNzPHPvY9f/ReU
zmHpD2ELJU+MuZbjfwMNlPuckt7tAVoTTD2VIY9PO+s1EfBwWmKIB4/7RO4Un2Ov
KuyknPbVuii3KDj1m3jk6QtFi4NUeREbMKsnOvCanUiHtTNUYZjhNUNddKfZt3UK
LrdWyBV2Q2z1Vwf8opllSh08m+B+1+2bPnW2Xbti+Gmg/QXXPjQjOSSqcq8IW2/W
bkrfOF8uxFf5RBwWQHhRxz2nS6DOh8k2159e13v/dO82/QBQzU4x8JdV2jKSaSTo
mO3fKNhBIPzFvlr1INbrakbkNDGn1L4deZ4rXFtFYlAwRl9UKlp3OasDWt2lUgh3
ygATD1NCIOlJw3xbvlkUQUKK3M67e7rq0Byi6RPLYenpgBpat3VZz8XdNkLe96tJ
mt0h3zq0NFs3gTzTUtWrgwylGgr2/R1SbHH63xB/I10fD2VWSJnGWSZwSOn+1NI0
espIs42zdge8q2jYezOZm3ShWG0rrUVxV3ASrLgB9/BPo8c7O7pP8l/GI5XC25b+
eFJocVCe9nCslkZggv/scRGmySHN5kIZm0b70FE+B1eg2MdqPiipW5Wf1WjzIioQ
q2X2b54xul+wcK1RNI2INTe1t74VClSLhZGNRVSue/Kha6CmWi3gX+kin93mxylq
/JrCnGfXnTHvMlq8JP+p4kfuFubbj6ZuDAWoHh1zbmx5fkzveIIf2tNuSLJmSiWi
TUNHQNYNgy9I0GfPcAwWfNQ4BfOPxpSB01UVzY+sQN0WY8yfVVUSmSHJmHZuNbwQ
BQGJQcKD8Kl8xjLFLaeagkqXpbbEeZ2egmytjRrrVfgkY4oQMqVc032pC6QI+FW1
fnJ9ye5owDxsxQ3YT7gOJ6uAkAcdvdpGAJTzLBA4XRCBZKrjg0dMhAL8yqEKCq3H
W+lEYd6i8Q3cWHkns+vt6lLG4WSqEZyNFP1zjAZTsemMu5klLqk2uK1gnvrJfYkA
jTQvCh9JK7j0jiR2F5bOQo+41Ch3d2i9RwTmy1+nvsYothSfjSDd0tKKBvskr1Hs
1CpIfjUL0wKRTpTlTyGN/Gk6fA1GsSm0BWFK/HQxUlVZ4L+6NW2MNdnt5DyZhvL/
h0CdaMjJhNode6i0w0FSBByon1gEamI6YueguWn85QLa9DzDwCKbPP3uDDoMvDM9
YJyln4VThqSAglNpJJsYCmPj2yohYh2nqROAykItYL3jNHy+WeevKgl9rOEvZtVe
NhmomIdfNvrorLK5+z5bD5HKzgM8KDkA4lQm/ACa7DavnKbkMdxSl6FBl6KsNIFP
4ktEeetkMDY29hqyhQTUFkF27ooJdGpLq8L5Hijyg7XV3fk7G+7J/KpOzHY0bnln
DVxLG3pQ9pISBQe+ymb90McUjs+c7IDC/Z9dinDpDO5l2SOd6ggLmA6OhYlyfVxn
TKjQ8bMroUdhNNPIXT3Hqgk6e5T/si6myesXK6F1CG2thCJFBlXDgSzuK2FTALKd
P+4g7X5YGKjKxRKKhoWBDcDT83xwXgqbul3rq7DzSe0kMHOmCWHWfkZUpl/lo1jT
j97jJ2TjhraUzCN1gwBacRKd6YjtV/bQkqnYhP/8uZVtcLXPMrYgdGXwQnBB0g/e
0WpSdyaI7A3H8uTJYcj8f0TdCmk2Gx7FNKVRmqFUgNCuDTvzMnb9T3IMu7WpBuiS
AKtkWU1gnIR892Nk/nRx+0hbTtOTdqQj6IDzVJq/gl+X7BXDVR0cnvKuXq8BqBRU
wi6ZitOjQ01EiY/ej9MwkP04qmMqNmeJafi/k+c3mB6T4YafHQSz6CdoGcHZCXxN
NA+8yswCRWyDSaH0gjVUJHAwM4LJlh9Bgihceps74RIw/UucRvZge45Bj1UNJSat
+45dP83rHH7iatxOgLawIbhOtfEBZAbp3ZNmCp/m+SmGNhkj/BB6Dng0NcWbr48V
c2ACEE4IVol7ELHGKv+IXX74KRyDwBwmj+Mh/TsMo4coBh0VeJbmQYG6iZGgHXcY
PftkEpsPKPLRb0Gb3p9I8Tnz1D/dNQsuSIfTuMsAPZco1G/LGLhmLlFPBNIelwHi
lBI5XeqtobzK9qDV7ApltDtl9KEl2mDv05XDfGdFaek7wX+kOlMlOCpD5RsWqcH9
GqmG6Kb8NYawZQl1XHJnsC8ZryZVgvEF3D4bhIN3o8GET+u2l1cGXsYCVcwziSG2
UpLJGS+FQ7tCKE2QmkoBSRu6Y6vZ73l8puLFO8hSrrQuMDwi/tmT1H8Sl3KldwpT
5hWKp8Ud718Zlgg/ZEGoKux8ACqzBG5bNyWQphF1LVUlSigzv6+g8gbgtbuvsDim
Njeo5Eb5jypWSTl7dNo71stNp5u7x79M526Tvj/zob0h0Iq9AV8SedPVpxrIj9F+
MjvFkuLma5JkjWT+X0Tzbulpzoj317PHOa/ksaahxXvl8d4fhNl/TN0U/kSlU1mT
n9FX7cXU4x/TQ8KXwkY48r3Xtca1rjM5qJYmNYeDcIDxWmaeB23KdHW2Ry+EwZ4o
Z3wUiZefCz3PQCwv0mDKNs4WIRAyfwEKQ+r9cEwAH/gSA1PcGgPcCXQmI9KIoH5K
uyayxrUUabl88PYGZHrfzVeah1zzxDHJsefXZpMfNLiJltuaB+AZr6erVS1ajbJJ
4o7WuPCJQ+T0LbLh3z0mKAdLuqcJvPpGINdMnK+609quMVluYtCVX7zYLFENm9MF
MPns2h10djPP3iVOALgujWgcaqrLiBSK9jn9NT9tX1B9YnvkXuzZ4gpZWD1gaTs6
TCGbKvboi6xKQ6tL/QNm0gxXo8M2YUk/2C0ehQAglnC4rw9O7ZDNNwrrYiiPFXbM
b3sYcyP44zmROz8qRVEricbeinZ/5cnFwCO4A+Ka2TUv6n3MjZ6GgoMhKBEMUFpo
RZ3k5xc8TBV6/Ii1jo1pp8hGeXxj5DAn+vOc3Kgm4gyQudKVQDk8tIcm0wZNz26U
NB2uHjJvNr9EJoprmoqwCoPRtHPWcyakObFsCmIQpN3sS9th/a1+yhG8dQ8hFeW4
qrsmi3MsZ2A/lqRgxixOj+7maaud/rUmeMLnU43Lmb0pprRQprpfRF9hlhh7OmQV
kRpH22JgDu432TJAtnjT0Sl4pluXFSMGdW6vlxRbxnzX1g8Ac3nAB9Re6OUPrftp
sORDlQQQUMMQcDICMZYMCMmKwuGO5LhZHBPPKgCnBWi0SlJKvfpwJXS3t1m1fV+p
WhaN+HXga6TGICceaK8J23/MRvrUJu9Dswj19U03nAvwvDKNs0yYo9SrSWOKdH5V
D2vPBF21Xs3DEp+RhKXs23aWjy+I3z0kBNbkw2n5Ds+D+iDmiUZXcplQ6nqZfz5e
JGRU1TFKmxwW11gdkwQ5zrAxw1xfswAc4EoTUP6BE1+tcbpramec+qiviaRcEaKr
QYKBIiRuZA2qFIenSH59SOT0uI6W8jWmG9pNOefYwEjFKr//hOtz7sfEkCxyjlJz
iDX5q38vYef/u3eUzK2jCtXslkX5en4W3bbg3AYTPx9AFFwtrzXJ1SXbcjwiAI6K
UXoz6ELAP6qckISg39H8MyWhsfxIE8dfS8B3MdPDMmH3tVi7LsKGJHwEc+TGmbOR
CBpPQw/3VjB+SMrulAcWcJUyzNfuAKcHGCHCk5x7TJSkfnJknzUNlLfOTt+ACQf+
ikuEH6fZfMUGMukWcAZ98Xaa76f967WbLDWaCsojf/ajRptOpsNPHK8SonEFN1eq
OggpVeXlUEVXu1cXZR+CTA/HeJixb+VWKunPacZBb6l17gnRMAlydi0VL8diLvBd
zyoFApWgA+oE4WbvC5XbLAKCHqwMtDvbCAsSs/xmCLGPxJm0gC754+xVw+IxKkWo
MirBGDNHuLndaW5aal4+D5fWHErNxoevQvVrjsOU/E0HUhhEjPG9tJWjYxwbxNPC
OB580V2qq7CnakxbXkI0zYL5LiBxLsMmI7UDRwZJgYdI1OYJ6ohgKLHw02yKNNRz
hZ6Flcuh6xXjW27Y8aOtFwm51vu8/HxO3kz+mh/LPTpzt6uDMsJLBg9fgoE1GRQo
AP2mflVgfbDQFCLRQR+mo52TTLMD7s40wgksRaAJkflJuAktTX27quNrRInaLGRm
sy7k+8MDfhXLzZ70tdokPoUTmKy356QZA8tN6aK/AvhEMtCT3yEhpF2ujHMAFjmf
RIOjioaetEri4eePvgT4RtLcuvftaR0dkNYuQLPKBr+TMW0wvmaaZhsty7BJveCO
SvfeNg0PKs7rGEUYc7mUOCJLpVoD28WDGOL3MOxbNdXcSyuZ09/Vz5Y0IsAni6oS
BxIF23kxT9evY73Sc9X1oXenaXr+9mjZ2yK+83bzMq/8Bzzgi0SC3D36BgCDuOrE
tZoMxFJtLwPQ0el/75o8ZH1ZAOWjkd5UbGIC9Dqgrx/4ppUX8eryypgwS5jqbITm
zWNWn6LKjLLHjgqncvvNbSvt+SgZD26uk2z8PU7auyYKXUrD+s3pGqaD5aqoufKm
ub00mmlokcEUdjxUZvLociApgsgdAH/yv/X2tzAyQvpFcfAEy+JJ/C5MUMKT9118
RFQmVm4ZUvJEB5ekfwCO1tkarhC07XbsI44SKOTBbuverXUQDGcoQUXRfxg6uSzL
1YpmJmjMoz0LNxxirGXLujf1bB3AGKu74G5HILv7vaP3Nz66SlolurcOM2f19Ouf
D67D5TdnGbvrEGbWNoebiYaG4uL9gISX2jfpkl7h3qRw57V8T8aLhJ+Ct/l6kda1
ODrsF577p7SX91DnlHdzeJ13TxrhotaK3w7qQiziLO4WOr0RAclktqSfmGXJZepr
v0RQGDli3HcY0kT3uWRfae2IA7lylCWTKDtzpI/FvBWGALNkbmz1/qa7wlFRkYmG
fZ86f4Ot6sIlnXFPIKdCSFQ+8pDJnFeewr9a6u+okLVcOljATSojFPOjhJsNNS9z
JlC7opSArFPESOtr2zqyJTeHY+GlgJHNzp49be3JqLQuwiIgaQma/Y5yZcVamnQw
5UaEKiPNQQ7fE7qL/i8tK7975NkWjsBwNx+EuPyk8tb/FuuPhkob/D8MPvUel1ay
cAvRlfEF1+qlGckCui8OCJ0QAn6aHmjZzEUKKCu4d7SDkaH1/FJKiEtRIQnMm0NQ
C5WUzEwbJlldVNhqbxXMDhLTKlK96yJQC+Nm24y9Jd/gvJAqG3mXs7va5ZMegRdz
Oj9o12uvBdEOO1hkx+crgIRGKeABDHwFCos1zlzWuxBx9tOYBV8U6XMzCLF6n39k
A+amMxMMaFRB2ItnscYP4ole9vlTpLEfr6cx8ed3+sh8TAU9jFDrzj7Vj+LzXZMk
Xk07+ICT/eGp8ITq1oi0XN1rcNmN/YDHs9df6yFQ66X7WOgb0mO3jDMMKdqp+l6N
jST4A+PQRbJp4xM/EmLdd/kT6KBpN1pb11hBareDBqmMRD91g8LVe4jwN8nWXpFc
Xb3jg2MNPrR69nUhYtD+vvWypsE5aq5/ArDPpTwQKar093lvyxkGzzV10h0vWnkk
gFm0iXleWjFfbLKq3EgPE+PVjiAks7sdhTIzYF33y0EGBuY/Sx3QSpgytFHZBBK/
LfeKNrujpS4xqh0ilTbWy2PakUJZvGgBDJwT4rJ/m9ncafj/0ZYyI1oSQGZs5Q+9
5hqaCNse5wsqh6OJX3AQDxpvFB20DhVcuE9QsDymUvVMtgzfzQcdz+NWxVLnrTLJ
zeLgMe0GoFjTie4GuoScEN17ZUL8XaTol/9ZY6R1nGz5BIrDjWx0zGQwwNyPAYIf
HWE9xys+5/WiSMt5r+pr1l64qumECvHGgFYlUpr8eQRkiAZWutdpakyLETJ9dV4x
0fdK3dCByHTx6H+uaIjWmDC8Q73ZRwxL7PJWSQmpgU39oRT+ouhNhn76LGZGMul/
Ejt+e1ZPC6Fg6g/w3L2Zb8DCDANNY/imFJW03mE3RkOU+Vo6Z5uetR0RCZBMaTMY
yc+2NOeKxahvXDbb9Nl18sOCUqys509Oid20SOxVezVdZpmDe8kUp/+0fucpIxkX
P54lbxi7TLSlZTwyFi3CLLBgzjQFrpoZmrdh/ekwF4f7IJpEmXYMZ1ZdMGkhNeqH
WEYAIPc+j0fjVgvElfCzzjR/mHKKfhRC+cG0+zsftjKKSNBCQ2eh/dOztlM4X+BX
3hRPO/Yzsw25COZcCGW58Mqe3gnjxQECvJEZ57omA+dRXGve8RL6+7Ni3Fs1OHH+
WAd1sgYkiK3gQZ06VcWYvqobK1Qc1mMeRXpfa01jT/9IlJgTrP3C6+6R8wSEkwKP
0NRwm3fLv0U+22o3MijT57qKLGpDu1pvjIe+PoALOG3IVoTpIZCCDUJFfI4+WxBb
3C0w4Fojz8eIlzaWYKniM3WXuPP946+pM/rY9Lmm5MefIMrr7kIO2pbZ7psJcPTP
k3bv8fiqFYSNi/dsm+D5DiBRZAW3OfDtUfP9+v4zh1H1lIIjOg5xFkFheLJM7VpH
8Huqkpum08LnJ0ILnOkKYIYGONIDr3A4YM20OGGN157IAoieh+OWjqNoGWYDtnHQ
xaoPyxgvDAmY84CI0fHH7P/94PXsNrZWCXSx1slY0xswnDT0vSo15syLz+bUf3sn
UzXcBO6+obkZydA28ckMoIJxR2hJUpJ+4X1lu+RTvDjd5WmNyE7sMGjTWxlwtv5x
5h+TUNZ54hc4pQqKsyshHMT55KwDxABwG5ysBpJyTbJJdCBR+WH8Z1eqR5hBsthf
+cxhslhFlN/dOiIWwg705vSktG3e3hcIce4V1vnPWbYzoH7eEkyW6WWpaY5St4qa
SPgfirBPd3mVoiibLqdguNRAZrNr6eFiZnAy144i5btBFWFxeUTD2jYyjKNrigGw
HRFgKf6sjCD/4h0D+fyXKoHLfxKaqe2u68LDSvJ2kgC5MIMK0zkdvuUT188o8F8B
Nqy73/Mk96BT/z5wqNiw2MsZg7u/VFH6T8PyrnbbrAw4Kj5CtkIHqixYVdojO+RW
HIYCzCGCLMEtL71X4SNyb5bOMKPXlsnOaUgKoj4Bl7ziuY3qs8VfJwMKwWZkQzyy
jHf53n73qNLI48ZXgqd+TzmC9DCR3wGbRT73REtqYBUz9TT4bQ+qd29SJ74ea1cs
U5s0U/wWm5XcfGkRvIl/FGcwz8s7OTiLxMd/HEXUzL2jiYJSMws0odkP2JZY7m+D
NKcgk2wR4MmJbt3K47IcvBTy7euswuA20HBtco3HCv1kW0IFyiPYVfEhRePA9sca
f4iLWzp1268Y7QGLjZcqxtlabExjwT5v3Xv5T7Di/uHFP/qObLajlT2+WGiurWQS
RA0BIKlVzBwrs1QvyUt4aI1fMFNDAbV4Y92JGcCCmVwfMe5U8BjepVKjG/jgFyaF
s0UrejIRQUzd7hv+tEc70JACrDNapufykJF+EzzKPwU3nESwi7u1G0Dz5cvmQx63
cfwdb8/k4ugp4HhYoxkovAaw6rS86tmsEqu2EiUZv0MSjzID2bZ3l6T8/k917pVl
jGO9r3pp35LqnQQDfE6tJHUCR4rcUiNX25+/lUNTU+jp20hzHHtC6DR2TL53nQDE
DSeIDpGbNS4GJ90suw6FufKoKqPVMdJW5+pyro9OJfd4XbGoSk7ZB4JFgJHUKB9S
eSaTkUIpZR7+beKKLkhBFiwJ1BNzqLBQFUHWc4fTpogm0UMr7zpvpEij7SuyyRKW
5PThxhAw6p9rECDlILwRjgqQoQ/FcpfP8aqC6BLM6EakXja1wesXd7jcG6Dhu9N3
1tBpCBdhWs6F9NsICE23AjRYxR0Y7g43EpYoyFPkCuolY7C9Kztpx6ZTHMLc+6Xf
+qYnqLEPg7dK7cGOm9SXpMeWtChLMJIlMrg528HslChRH5RDestgTaljkK8Q5jcq
DWPi2kXTompL1Js0N83DbNky+6xEXVN5CIl6ptncGlbuSRN13u85mwnM+26jqvAR
lEO0hE54ke74KaH9KvyuIVKK5j8x/F89fOCz+V1ecpQ=
`protect END_PROTECTED
