`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3jHOqrp0GpnNJMy/v+qMlw+20rOYBlh2wkRqlxXatqSW7tRb5/tRw3d2VXZnVMG
Wir1z9O5RpgS/P4ZqjuDMRReP7n8U2YKM1Ptp7hmI3fuaZCddAiiZY0UaAZ9U/cm
gHFtQFboFwY1u1qEEKUwCpLhHohcauyz/buVSD0Gx2ITWCEn+vBduVntago4Snqw
t5/RC+Vzv5Er2N0RiOdLl7EGwZbr9bQPjIsF4wmD+ciUZxiQtkBrKqCnXCwyscxx
LFwYL0wUhrpIoK+o+OKLkLtvqxJUTqY/8+qXLZQaxxopyToZ5s9Ze/39Q1Di5vT3
fz3N6La5Adlk5MwYuHzEuFhNpXVwyeQswMflLHOyW8qfaxCk9IXt7TFPqcoKE31M
iCSNxzwndIeEd8lg6bseJPl2yhn2fRvdl7UsTUeipl/06WWlOR1IEc5bQ5T8MeYR
cdWArRcxXeLK/VieHHXMurj+jvr6VCNo+XoJDtixtmZbt0d3CnqCpL1bYxqmliwT
eQHhRBlqn0cnTIZ34swpWm0pTCg/QQz0po3JSZ48fyWaD7Tfp4N02+Uf8jLiOmwL
pGYPO/z5vkRvMIxVSI2bXM6gPAZPFwJAZgUkrPDhtoTf3+Imrm6+M+Stf8VAT3ji
e3LJFPs3ymwDK2dfTFM9+aWnSjhCersb06DuHXb5Y7z9V3CIMxIJC6MiCyk0ZBkd
IpBTBNzTGghczFpSXL3uOmBpFi8foX8C+tfKPWRziLK+iQcgR5tIsDpJ9jLYrDgx
5Kvnq1zSi9XrYgxxTX+ReahRwZkpEjiV72Shx6mpd7gdAiPE1El2w0F04cOZ5UyL
W0XA+WV2Sy30TDSbYw4atYWltyEpkofMA26G+UwMQn+mojAcB+KahkzdmHEIRvrp
qmcCPEe0jV0W4OnzvD4sInWRbql8jxzqQ2shBsK4Cnk/ear5q2LTSkdDJU0c1sFH
NtiXQf4PyXqYvD9w85FKfhuBtuReoBUg/j5K7b6wF3b1zeitJbfVufuDKJFyRnBr
OUFssjTicElcRz4DT+AuNljNMX17yFQ2WVNL4Tzfs4KvL3+/fnd0c3clHJiPxmfl
KBur7125NelPoXKO358JJTMt6s8c+izIfC1pohWLZhZ50xpbkrobbnvA3dLVzKsB
OT7fJRkBDi5T3H895t8M/uZrAU1Sy2G/JahB0LMjPwFrC4HPz114BqMos2PMpFfc
y/3WHitPhby0Q4npMX05zUs7ysp1W28uV30XAuQORFKwgU9zM3C5gOlNR8RIDAMC
jh8gEVJdBVJG7pVdKs88Z/kIHmzUi/05VMOskpzQNpoDejSAqPla7F9tHf7VAnP2
FWojZTDUmbKuPLKzci4nO9/ump0ff4rspG145CuHGhClFU4wuAbuHwxQf3AWVKTe
muybIo8xP8rdDUAY98HoQAg8mH0rh2v2NNo85gvuPqNwRjeZIT4lI8VRni2s7MxE
bpaR0CQdHBQpyzchkDbDS+duHTGSIK6fOLV6ogYuq1OZhUj9e7MNmc6Ta/BdeQXY
t91PFwqHxmdOfIOt7+hxaTauC9S10D/pwb/I1V+g5VRXYdDIbANnqNE6BFnYRdkI
BSL5Liz6cHu48P+1x8iBBVcDKeIRAJtw8tTjgqKXtQbbT+5IaqU69bIFjZnA2DcD
ZANKsI/fAoVYJ4wrw/qMq1UFZO3U/MvzjsqmcoyeTGA8TD4K0Mlf8p6Vy9dTSkZr
0GF3b7eWNZwIdIxnxJFlEs5ZPPiiuM2WBcP80De6MwjmhG1c/+MkUw8617aZ/qH7
H3zgsrLHJQfanU+0HJUCb1bFdxOHgCmzPKLqE4CXt8mkuyLNCzsnCmRvoATUgFIt
ovZct0B/EyShTGjgYZINorRhD0HAUo/mB+akNGQr+V+hJBgHPtmB3ccdEQWQqff2
OCw3PEdXB/BOFCVDArhzLp/pvEPLEwDJXADMSdiZEeq3VWtO4c5HvSJ9dEU7V6dG
/qArJiBma1PL5vn9oy0C3QBpXkm40Pq3W4vN/Eeb+R/uMzcTXtX9j/dGH7IO5sqK
YBB4rJIDTU0XroUvdonzehbdR86M0/oYbidI2ApOQ5BuGGtgvA0amFNbtaAU+5NF
YO1jPB/JHa7JrVSocoGz60n/Wxs3haeVQM63KqFiEhprjvfj1UCMVlzzkeqD+5vA
jgiy8/8J6Qw8Fvhj4lzQTdyqDLurevTvp8B1EQQLOpa583FT4dgqW87+oHh35arI
nGRJo8gpWwLZhTAigT02weYhPw+60O0+qN5tfqi7wF5zBKsCafegq9KRVcBizgtx
D7CDsDn87AYYKDBhwqirhKS39Z6exrjCCc1TOij0BBhqcn8Sldf6m/65RofHNPdK
syhZnpfeTvR+P8fK6LPXB3Tx+G5MUMSFWkOUe3MzKnsuFf4s7DY8SPm2iJ50nnqd
AHwUoQsjwq/SAezz6rRmaKP0i/IxqRZTVhJOLKVtA9aiVYEFP3vpsmA7kjL39gE9
3wAAUaxukRU1gPjge+zVWTdD9PlITRRc4VyJY8a4K/x/yGO7WE/oDZkjvDObnkVz
l+mr5bkAaFsvXcs99cIWXyX+EZaXIVv3FwOmAIvJiK6nS5vJfqRgFgX9Os6IL6Wm
Kcfb2/EIs2RUeJk93SYBKZ/RK47th4EjSiwWflkJJqLajCURJmxYMYM9bI8CAJUb
KILz2og1sh/j30aThiQKRSYKpC8W/UMtkIevZh4UUaKlKtMgbfL7/VMd6fBOThCz
wdCg0NljJry0d7ORli83/tnybZYASk7M/7h6qKyM7TVI1g5VCvtk6DfwrI4flnHt
ER2ULEeqsvnws54JlHBJlgXLl2KF2Ok4tZUxAIO4cmqxkOpY9DrzfmvNlBb8m6xd
cqwIS1VCQN7t7amAFpIfeud42njTRrweIeYbf/Fp7b7qjR1vVTiWa9YgGqO6G+Q6
DwoyDCek6qQufhNzA0HSQgFuKqUx8q7B/7h5b4pvoI6d7iqBM9SmU6Hm7XmKfb1O
7JDZembxVMaoVp/wbri+fZ9aoOFYuA/X8YKZsnJhAOzIQnbWiTlrNcW0GgfValhj
DcUXDAlHH74hzyB0y9qmACAN/u3q53845RHRh/+fzaI7oNMdGWCMp4xmCgYw4ipn
Iq3YIAV3lbCYYrz2syyrp4eqEF9X0bojA0F4XnGEdTVfKTFQu8Fj36tqqBGfWJKo
9W0tWFSbtc/neaflbrwqk2wtc0wwb3K0s0E/kod/vAJUkTniY1QMifLzTUF6QBXU
Xtyqc/haRjWgin/0S1XCJDBMJTFYPK1yTLAj1tDCoDwYe23UbNuQw8RDFr9OEQSV
G4p94lIi+xXE8DkRBdjlpOBUK8P3Ue1YVnGvbCCJwDPq17Y+/OyM39Drv3RUsN6Y
AsszTypIcVwfMzEmF4fbjXTkivq35gcsXLIbRNnODzAx3ug6NT+ac/woFVWRnOgM
KA3AycUO5FOab9Fs+92FhAq/z2g3duAyNatDaAjX1MvOTaIxI3w4wXeQOtn22WhC
k5PEMJDWvk7ctmiUvSf9wOcn+QNoiDxhhD+6KCl5MS8mjUaN3EuDtfDnMPINXEkF
PEmrzB+JkxqM8ayprx/stidYI/qMuZRMOofFrIQQtFMidvlm+M1+sGNo9STOFUyJ
juFlZK3nQvYb+39+k3wxoW+ZIMT3duuCsg8WIdUP5ZfuaEZSF+TYng8kai7R+JGo
QziNfFR77Bs+4ZBdHx13PhTvbCrhKHYkzsVdP9rLyBJlakRgDtVQviUnmE0mH1V7
K9NOIoF7jnPkTmpOIAcH75ZvmKC54P5sLizJ4r8M/v6H/ZG0APBPJwTWfDPnMOS0
lifiYvZVGTgzy4xCRaJ1ue+t3p6LheS27PxDVEG3mWvpmUfLYYDxX/U+yqQW6sYE
3zvIy8Vy/eIytQkikek/iBSOZwVdFNcbeRGC5ee4Wx58o6JG94VVHN9ALsnJ8DGi
kd4Hl5beypR8LqW8VO94XWg7tdaE9F2F/9lXeUvTadZcEeIyc7RxYVcDQqlszbh9
bxn8y5XaaYRWNqAGUZ9D9eLjuW3K334bpU+bxJmxraAByTVwwIOESMY7deRSGKTX
YQJx3qIPelG5jVyCWcwx1nLbj2CcJCrmeHy2u94dJEqS1YdObyd4iD6NyoWUv3QG
8PNIKT4Jp7MtJkjn5DP5HmMaoYE1JUWlYPG1CfdTh0eoF3AAD9rROg5kd3QY+76Y
msiU6pANzgw98DP9rxvc/g9pEbtoNSn+Jm2Zmj2lJyLzOIiI0dDGnslZ8s7AWOi/
QKUwg4omoYVCFQHjzN96KOtVleb46sUp8xcU+RRd3gEEkH6eHFXbRhieKPMjTKMB
B6g4SVhqwmZMfupJSMeyAxNEQnLfmRv0Va5fySzRNTIzCGAv9U0cbAMtQLXGhhJY
thE4UmD4lpucMQ/bn61Any+G4m3D2KEySQuC1hpVt3jgMHRGSm6NtHQhIIJTbGK0
+6YPAhU6N0YYTRZCmjNjzC7bdoJiZ3piQeVA3Q7f6DThiXWGsL4EpfigvNdPBGlB
c2X2C5+YKCNB91vzGZwteWfHFdMTuBDd/5LBHMAZbhpLDTC0Oo33OB1/qYvbR6Kb
eQbApHYHEGIy0H2LKe0fumHmWu7FFYyIi93pMZLazRG5KWMtWAH4TrOm5rW8Y//K
sGiinHkZ4pAOuy6o/MCkKv5FVoSq3wetb/wHTW3xII4HuYvC570F3o5VmamXufuh
IkRtwz4tJETDM/ig9EYmiOhJgp0P12OYus+KZHUIZk5GkLTP0Z8ZND5MxSWhgr/a
crjPmQjUxzHOKMagA0jgNSNyTS2MyGo2jgnyRAQ+g7QvIRu+W6kZH8W+FHmhpSQ7
bna13Vuti+o61UEHL95uDSXAROBkkRck2KteiT/oo4DfbbwSdeRnv1a50rosQzRS
5f24hg4p76hVEjPuBJUHOkS31u9GEAqgokZmR/YhU2hfQWmL/w6tTviB9FgI95eF
SaUq5rmHnFXhPYk5LJuPt0fPdMe/ZqKIKXWqT1I6NzfyDArLYuLKu3ATEdfPs/OW
bFtdump1WOhpoSBnAZylpnzmOzOGjZhEIYNqzclnRHYqs33DcL+8oL7lVVha/Z7P
SZnPqfULz5u+9sDH+TquNGvYVvr+7d684djLVwFPwQzV1Vp1fgPQ1QogMTn14igq
aBIjwsRbByE6rXEG+g1qlPO62Q9Y1KeQVGs/8GPV+tW8nqd1LMCnp7hGPHWUJRHD
3O2PaD/lbLODuzU6V0aGjTjKIJO5bBhuXjA1uCTsQNrFDonJ2X1X672jOp1n6Lrt
LhuOTEMuM7BfDWiTdfNly1YeYWad+xBufGEszDQDoaHUHJm4imdYO8ZK+a8Ntm0A
KxkBCS3lALHVbTUjQlldexaeUkKXuDApvfNhaPFuAQX9a/HfmF4xHiWMvEUlvg5O
MlRqfUiN6AKt1vQckfua9jA4FRJfYCFxhpNa/mF7g4W49rKzskCHxElRvfGAahWs
7ymSiXTNI+vfvZhT8NOdrbdTHUpVr2GbWrGXccSZVBrU++Fs/2M7QIEM/4m3Kh+j
WuwrPVsRe/6/cH/FXkvLFOFxjJvFGoIXwYFFB+lF7ka4cvsbaRelPVYrsxA3KWWo
qkyokbPCzRUdfC2uVQj1VDqVmQ1nIvYvYtnVJVFUdKJOMzJkaV2qw5KadeehwNYz
qIRN9ZzjYjz8WARbG8h5zfjaksPduyu6p4TIWnN3D3CK/6qW89VkO9iqlZa/7sCo
ZjrE18oezDOUQqikXCkFgWVzg1F3D3liRTAPeA1xaJz7aJGQDk7jlDGwcU5Me17e
zLWZw/YQ8Yl1pL6PAmCFIq1cD8w1W7104tAzygt795Hp024p5bHwR0+sDayBbyGp
iEaT4J+J2et6Jp866348oUSOL1DwmhY8LwVzJi+MbQYHlNSkA/pg+/nz/aAzQOpz
Xyhadf+hG3VI3FFu1Mk0XAPmTJPGpdkQ2YIZOYXFx1s8jCRQWvaI9AX9ruWmR5Om
ulr8HM5o1nFHT71Cf9iK5AANieG8HrfsPCt2ff/WFscoZeYsZuB9yyRZFc3x5kvd
R8KDqDAVjkQUpkDG7/4THqE5j1XGIimPcew9I3ktqLXv9ycyl9OBirL5idseBJRO
i4JMZ4JfLmlAZM248odFIX5G7oqzEp2EfeBuwYEy5XVBkIhkzvumwYcyR8TpWNAU
8G6/I+Ui455GxOMYNXGVa9bt98dVAsiJ7bMNStgQ3VUaR22lpBFGmHsrFDiEflsX
9xAkVb052JdK2z4rD+IuNDEYZdxCrb8loaNtAwZRMlPXeRCCdU2awTG19WWAe50Y
+6xxQI4PlyeUqLj94mmd2AQtjhD1ZRzeyvX/OoV3YyZuaea6OriT+VtYT/nxDgS6
gUwAPKaH2S9Dbltnwb9VP3DWTcZEOv1BGaqRC7msS9C5TwaRbXDBXGcKB3jZRjlJ
0pIva2Ypb4NuXRzH2x5uvF+EnXNZi8+1OIhseE60kF0eivNCaH9BXwH3/J8Xzmlh
1Nz3hbdllpwPUgcqpyqt7A/qlwPb+RnOys/Sj7Ip1ezg+IYiLUnVn1aN/K3nbmZi
Rm1kiBIgC/Aq3+LM0TURhStNYE5FWQ/KJjd5qYmvt26P9ekiEQ5KPnsz6YjTT6Tl
LNQ237GZXFJXJ2DNYYdGz5r+uesJ4MLCqjpBIhlCRj3Mhk6BVEd7M4Ppt3mxkrO6
SZ1p+kbqqNZGOsIW1uwNKKfOm8NslA4pfxJ1O0tNhwmrU2Sg31ovPWPYox4TGjL1
3RSHxt9GlhqqC2ev0Qq95HA0VWaHxxS/2EwtRD31/muXic83QVPvcQfpIfwSnnyb
/8gDyYCRdZ0I0vMd8DWy9m411QBLuhDTC2uovCx+2xJaq/vIk4oSwQDAZmNMiqS9
IDYagzOunKREHQ1ES/KmG49aeJNDt/5GDBNxSn8rXvoxPgqWDk58B0wcCvo/BRAT
h74ozTX8vx2IijeI3pRUDLVX/AgS+Ou382Cj0D2d8TqsEBfg45PnrTdBHA6Tzalm
lRdC+oBB8ZKYldIKrgWICDgGFMrGSHOMu74XAlJsub1Pl64HlV3QJH2yTyWLNwvx
eywOWcJLk1EgHvPhbp34gFcgi58OrCv/XTIfEbQKysn+NYOeg+HXFimzNc5nZRTD
Xn7c1ohqncCb/lL4p12u0JHrKzuOANeqAPxic4LkrdLQXXmdogtQAuaVSnnD3fWA
BuPtyVZJWH4SImBQhaQAJwu7H78IgB1ymKSKKp8FlpfOUnc+uPXvUxfDwY1pFeRB
L/8O5RO/zdn25JKTBLSJx7fo0nBUs0JfQ3WGvfh+EfXe5RuK1bTQuthyBhkuB9WI
7zIQXe2Rbei8h71m3f4NWSYA02k2RsdTAjsxg4osZBtEWY2zQqmbsRkBaCjrUMgd
5xOCkeJaq5l3TqXDHwOSIIKWzJkUG5K8GVYM15ggYiyWtbE+ENTbYvcBgH+UkNHJ
7WR0yJFwVTnsof1rcmh0dxIamflOcGhrkPtukEkGIvNMz1aok0QImwOpYdl0b1Qm
0//NoM4dw0foaGt1LYL5C4MdhxeOYnlSiSGs9UWLTLSD6ladbZM65rxRGR3jZv6F
y1cOax3R1pN7GKoNh2YnYKwQhy+JTNgzmQoymtGkIave7F+1b/Y9QbXNw//loJOB
T8A9yvw7dojq0RWzR2BWOfNLjUxCNNFDZJsCL32csHnCpkQJW11Fheq4eP8Yp/oo
X9KdyGsXPD+m+C53FMLl8BF7j6exSmcN+dn0k3zNRL3kUmdDGMs6UR9NiS+AX+PN
BV2JQdd72Z51i3BlMK6A9t6TFLUD+q3kfJZoQp4oYld/aMSddv6eCA3lbDcOjSof
4ud5fCr2/v1PWUyNze/05tgviqbVYF4lUGGU5v41Ytg2HyIKetItJFaEPVzn5+Gk
hdC13WedRISdr60A9C3poEyNzsUbJkfLPyoIRxvjRuGKU1YedVbAV3R6zBlcI6LQ
L5PwB5+uWcTTjGa9jHd/ONesGMzRbH5U6YEtSM9sYmdR1emkD0YfmRz4zOL5WUtM
pA6BMhdW4SzvZ2RGGj9aaaBXbjQos/F3O7vkzeuXiTh0+pzIlnDDq15vblIWfKyF
P6OI62A0jfVCLaGoJmGcGjdy2NpgRVKqZTuz2SQVHd4nzLa2niU1gGt3mSK5JP7h
rBJu43nvGhy4EJlxowdaCdW5MeqzPaU7snvofKM0SyxdXFMTtQNZcEoTbhseVJFP
rnOmEPxD9FKtLUNt35iSS8EBmE+QHPtE37JX7ZHNqxo2E8kapSesZw7ji1q8Od1M
SmLuAQBLCyLTjcw5Yx9G7tgnljW2i+EQ2fkf19ZzOaMC3Ph6G5HaqLX72At7lA3v
xWOT9oSIi+2/RlwfqWUvV2WV0xyJVSP1hNjDvZaURB+2soB9xjBTWw6FfLtIWYyE
DoZSf8ujW45mcPh3QSikSfLdWhM9AMtoRTI8d03uhykC5KEEgOLebfmNsNEM04fH
ujrm4ob7QhF7zx0ylIQ8I0FAgepf0mx3DNlpUcFD8XKaVeLXxTAWUuLAA9wEsv0X
BDevO0GWx4/Jgn63s+ObzRfceSPa92UnNKOIcUJrnCkgogbQUAolUgwwvqQcoQm/
kzWUurlw5qseIxbP0mPtygEqFXZiGxYgR36UPhreHTKJwHVXr4ZOlzDK+SD1xAUA
3AzAkr1Tgns+OMJS3w2jCt+RxbGqilDhIGpbZj3Ls6kY21U7AYXMNxdQOpqksOvt
qNKE36smDGC+zuMvuqX7ED2UMYVjmAVY6QBdN58SMfULQWDqgqTJsdFpUkULzkZZ
aur/TJpJHhoJKR4nvaLPsezXikuGQaWR2QcLQNzn4jfmTo0BedlK53hNXWeW+1AT
eTDDtMjZu/nlUeWy833qUvKwnZUXv8dkeUNhHpZLuyTFUz7odQD3XbZh9wLSPLmV
muPsCUb/DWtYxi1CY830c4XUT495QSAPjovmHYv4liTw/3g1PZUa7ks9MfGR4BOA
+3fdadmLeOv0fBsdMTP8+8+ceVBr/KOrKPybeGcUdflxig8FDogUw/sprlEZDKDp
bH2s5bHSZULN4YG1vbKzBXjha3fvUgOhli0kc5hzosPtsz1QRxq+2nOoVkw1LmVD
2dwX6ygawRtmxJVv3pB4rc6jXkNHk6VCHtU8cHBBGuHSgk8ps/BwOpCwaPta/7To
dNgZRWbbKQdA4a1Cfy4V/yych5D3AtsVaJ2tQcJ8Wd/hrV5bxml3RO1sI/Fse7Xa
9POY6uK9lpI/uTyRWLccyViCNiNRvZHTSZJAIXghaAyF28y2iGfiSAtdikmjmOjB
99Ynth7SPlvG9KHAgk4JEY/dHE2fMYq5+Kf84HjG6meSw8d1j+2r/+ua+3UNlQr+
uUms+3R5x6VD0ecunrd/iwGyLhBEKDe0noFFrWqghjBpajC4NXTmbFl1HmAVPsbV
D+PuB6ZDcB0p/NDV/us/d+eYzp+iR80IrydlHZ3qmXN98sYONmmbDpsSe3ctdswc
C1LTGgjHsE6LPBUHARBGHa0HVKKovnJjwejcuEFrN9RhG+k2bp+txd+RwwDqBzS6
q1dE1cYEoPwsxG+eYJquHu+NCbH7kLMfr/HaJBppGKPIQY3YKqhHsQx/3teM8wKb
3YMqDakoBvunW1QBksh/FcbDImZR5m4Z2bXyN4YO+PGLhH0FMwUw3W+Kj67h17J0
aoUlKPjke1rM+TjuwNaW8K3VtFNFkM/3w+DKufaEbJ2NbJZNmmuiVKxe6QF+A714
0X5wht/nY1KQKB9qD25Tdaz1mBe2MLfYgNceuAv/DDVOaL9AEEDhCJzck2Wns4/J
w61Lj39qF+5fR5lqGRxqTyHlkOg9PFPNNC9Z7AHV4qziQAYucjCMk84kLf0cOdXx
vRIhdTSX5PVYcO7C8k7yeyrkiKRy5xajaN4bsh37Kn+6NvzZv4eg4aaGLDfXtmqF
xDWDIWCVz7xkirlJPCZPLDoFVz7XAi8UUCgk6rZAdsxB1U3j6AV1HXW7zUfKrLME
IMmlQj2PIiJQCgP2tOjZRWoqvxk0Qn4vaHsioorT6GTsDyQwAVtIoUzneQhUeQuo
znTC5fxQ+cRZqwqokQNmfo8F9qvCQiWYV56DXR/qdRovDPP9LfAyddmdmVg6n/0u
HejadNwqZqnhUEY5BfDAdnfWpUbiSwhsifAb15goxYDQPjWf7h9fnXDLo0lNY/19
LfkbPZOjaF1BAhOn90YrvEtYoGGosFl3H3nxKL+an4qoEHK7eHhFfV5p+P5nWJDe
U9076wB3VLshZw4kQT04ooizP6wRskgLg6/gYY34gPHYNBthmsmaq0VxCl3WAnBu
3Mi5MSCPOCDUhiwHqvNEn+A5qIxRecVxbHp7Hf9RpOPw/L81LNP4OrXP3OJuWpR6
lomQF7KyN2g1+R7rJ1XCUPs+B31FjB/GIXmHI72zxFgqi/ufSeXdM0rqFl081/WA
7wfOGNp+qN8GgoYWJX0bOGu+RZwmYzFrkageNe+AkLkXtMWsJlT6Jm6X3MhZjwI3
HAyT0M/k6OisL76liRCY0Oof4GBMCalTjT/PdR25fTkgIjMRHCPlz/+jSSFUaiJO
RYXPEiu0A2XnJ+nxN4CRGFIsSkF2S1hmq2i5skYK2Vh08SphlibB4cLB+esmh1do
rfpRYBkbREFFafNlNdPrnrnAElMAF4ak7x5Aa26I+5USrcnccAeeo0CzKROSP2WQ
ezAgKJvsnzrwpqfV+t8Ao6BCJohK+64R/pFvKgYu7jrAM47fDynmbeSLzz++F0yR
fG6tOvvL8Hwn2oUjsgQA4pBZPHBRKewbK+T+KN0l5wG5vZRzRfyGh39ujXJBATUx
tOJI+EM6pqJJXJm+OaxjW/oLTqjK8kJ/pBzDCh7Hzaq93j5GMB3pgvYHw9Ot/MQy
FGDRZkidxKkcPLMKVYpHx8cTsI/LI/pFS5SSiq8TYzItBEaW6FrH8IdfnSKndG+b
Wot1k8JsR7acPpMKYSnojuBOPvSuf6R4IeIDZRcAr56aeZpsuiigGbrVFU+hy21S
/5RGB4mdXJmxKs/aIK4aK7JNtLxCU+/ubKij4oBsQBwDba2MmqdGRtlkb1EhBMbz
FSEDDxa5REMjsGRFIAKUb+614S3O8zbQS8Ms7lbZ04B22sa8fU9IzDkESYdxyDol
W4gyIcNhdJD2X03hqOomZp9TVZuzJuiEKE7w1wjYqzc434Cj1EEkqGeD0qIQaGsa
VXCsjUe2nDWKJCGysctIXqvQqAfbLhUkHdkJmiaB/zHn7620mp4vSG7flIBNclQp
m7/Th6+lve5MDwCuiUUZEnkoKGK1qt27t3eUlBiaSsqjaecH0/75eVJmI8kZVFgv
xEf94Gs7ExGIGti1Tk/DcCfsYDccSbQdJXx4as0St2m3X6ddnxjo9iIZn4V6EYKp
sr9j0Dpfhmj6asFIDsqH6RnOhMAsa1KCzhal1PjEPLMYK/szZBnDsM7gGIk6IyvZ
DRiV5BVvdojMW1y1pzRFkbxK5Fn0CUoq0+NtEFjm8r94/OZ9BvUqomc4RcmaSZc7
C4wQgZtkeuM9+i4ldLq++M2TdkxtJYp6qFxaR1qSzHNh7ETi3YIIqC/5LLo/iWkx
C8+PNzZqAGVZO4nymiEoxofJ0kS7F8UEM0bAYAcoEXdDDzGLwjm4l9WVo29NOlHJ
aiEc5qHEBuI7mQJTi5eHQR9cIWqGWMECIeec36pZpREjFHmzpuM7aL42ZjZGO9Q5
QlWtngXWsNclPU68MkA1DwmeSCwumRLmmmwMtt54p84WL+q2CoQicnz8x414snOc
8bSI0C4i5Yv454nlNeYubUDTCmzQfz3oxKsuJVFo5PZVZGWe+mWVdgRiVZIkMDkM
DDbawIsBpqpMZLVC01wajEgcTIumKLNT5Axaqoxb+b/uZlbFCVrJ0MfmRZgp2Fhe
hMiNIfqGmDuMlFQqxoC/lXB9cR4O5eXYFPZXjaKo0p8FPKQOXxjRAbkxYgs1pyBy
wXHHuToUYon0iVlHJRGbdMmWOrwxWHHzt+I7XBOmaKH6aV9NR8wFPlnqc3ii00+D
G+QL1Yhkx4QpRofbDIvoKBt+516+SiZY2zfa41tkfi/4i8bnZ6Cb4FhD9h4Bt00U
JaATGL7s5sjbKWSPhFBjXixLkZv5GhTq2iVaaQk9XL4141P7k6mAYlaB/AEuh010
Kow6Oqfko/CydkY/BWnVI/RVHlOnaagoU/dEOb5G4MWkpQOZaZStVBQmvj5yPxSi
/QyM3U3863vYUC1I5qa8tzLjgIUQu1uCABkToef7XuuJ3MK0nHgB5W/GKBagr3fW
EL3mwJgcvRFaq2KQdl9OeIPEI/G+FWu6wT61qbP7NM/KGSvHc7D/ns3ku+A5w7L+
GB6qrnctd17SRnJERhraHP7QlVrbbEtnaHZZLm1VRGrm6okk4MhoR7dvp6TetJo+
gojr8zrmG+y2XqOtIX6trI9NpS4a+nvt8tkyVdCvS+CDUeD6RKVYY0Z82Vxjfps3
WFoxgGxM2U9P86o1zqYFdh2lh4vtf3sSETnUCayYxOTHopPh0ugcCI+pd9XdC1r1
BBu4yvzWq119yhCx0y/gfIBjGCGB6hbLez3BsaRYeGc5z1brjqEesrHr0uBZm4nf
t1FUROCIMzjv4yRQrxmgmZooFapzgcw0ksWhlkUqtcwW9UBwThMIFP47Xz3nr0g4
jEnbAGhbi//ZuDLLPOnBqBzMMHBoS2GapzGjG1UgWaIzYyn+FIzAu/chQmvxwTYf
572iMZMJGtpYWSAUHjF4UVgSfh7eEu6xKYkBEOT70RdZJ1mWFHdc0EunU+0BTFyQ
t7w/3IpB/EzIraeEWKDUyhWHWKzDYNMwdHQZSv3h7Au380t8wgGjq0p0BkVlJj2c
c04DMntk64XjgRVwAHcNq8QtlBqjIhei972rhdkETFRGV5e/IUvg8mZnY8Id67cR
TlhIiTnozN2N/aUd2jBrHzH9v4KqaBU4zYncCWvp9A1YEmlCqnPLslPpwVVjT038
2NzpTsxFUITJfj5vsSr1wzspQFrIrVY82MsqlcleqPFi+XO9HxbBuwT+Aj+FExGR
jBzq4f/jTTypwRRUZ572gvOZAns4wJOp/ZdWQDhMCD+tsahGaKuWC6kt+jG8aYUS
DYmoQWfSX+Yds5fv4DHJ2jbizGIQj3e9hf9NwlkzP8jb0uyeLfdmsr0reJbDJtJG
JhHORCyRc5KoR59tKRC+NjoatLI923ZAVl6VK0HgYX44QI4qUYVLSuPIQ4JzFnyh
hoOoIwr5bPI1Dt7LGrorqiJqbVwYvXuvcUb/YSbh7SLRsfZ2RwgoGd/aQJljikxO
5LfEqKYewdiqBXR1ESp3rmqcy0mKz9e3pgDC9Nk+QsQvGoA3hB3S4zLUxA/vxkpG
A5YHhHJaw2gCE0eruV1QgtGdXvKqDxeZfkUUrG87wU2jlIEHlVCjYIOGx/wWQXcx
iU3vg4O0VCgk4PB2uoRLEdURqB1FHHR6iVs8g7sOrSvf8vmqkprMaC99sXqtFwUY
+lCOjLJcIUuSrWHclqaRGa879doM1KYMqa98mAnYoyYBJa8xdBL4YHhVtPV/WYWL
ckj53lrBwG/vu0jjOIG8nQ1x3Yz5nweKCYYjzSsk5+pS+hRkZpf0FGPrvE9qvNew
VCVw1ydSL3N2EDXHFtW9XrBhohaHagetghZivA2ufZ4toeJdbmP4RPBGV7OnlZ+I
qNiYzgZog7cv+67SZsPh1Dsz23H6hNJ9ovdBx9FezRBiPH113XcipQCBKINqQow+
cZbnM/Mm45WIN7FlvtmU5sBt3VOEkRs1iw3lYmLiLOOgYdkc6Gq4JqqIioyr6O3I
3VZWfkENCMwrC9fjifnViUumRiWnoOWGkfFb6oohUPniMlJbOXauj9i1xjroBkKB
FYvQj1ek9wR+tW4baMe55zUqTPBUSJnH83uTV4R6uL5UFyI/YbkKiDPAH0P9lYHC
pM24TV9plSlxXI+tUMF1DEDS7k2omjgXYbPiZQxcAOKCPxfHLWNU/c45zccx6Ysb
lJZ35T/Dp1/XoH8fV2+o4SV/L4qZKvMozwsEE8mCQVOcUeq8/nQ8RbvjiD9CTgTB
IcHcb59sAjVWOwm6NzVRn+dG1MK3lYxRmexWmtzhkgny5gJ605da816Ndo9IiZne
0Vg8wHtVe9FXB7UjGcJP50r3ETi+d1aed7Y4ngCb6L3G3Fy9GehjKoLxQv4fz/WI
hHK3kLvzPQ6sD/z4nEh3z/UQTvsNUdxAVfsVw2rCh2P+OGhbnj+whPPwcYci+kA+
IWSieB9g04OpyAF2zezQP1qeoYD2+ZaQ2EKMqXu1ZxyFrC7CAjv8deR0THegJfUK
ep55CAtvhP9w9FQqS2EJdQblrz5p7y3PE5ituish9aob9YRZBx20FT9PVO1YbKXB
rFhBTLfdbtpUhZ1rDJNXjdCBuf7sMbpR4J7JHIXW1zPvV2NzAioCZLoB7BzqnHlB
oOpQ8XC9QYHcqqwj7e1YFspHaBKrkAbqHAkafK4o50Hrm/aIs7YIk4/noDl0ATet
nR4iM7Ilzbxhtvf2n2PJXtp0U4fvryCx9CutwjmeHel0EtcggCsPl82is5MIALbn
Visoz2tt+cyPehpB7/eh0XFMbDJ0WGDR1vQVBY5WAMNzf59c/6N1YCz2lVQbGOwK
ZC/u91rnlW8qjGgMy3HYfELzs0TepNPPmK9MC3D8BYTVIYUJhZES8sHoRICIuEHr
G36QL84U7Rp6GqEXAWUAwTsqMNAWOuN50PhL+EwesKu+/ys643TXhzgUgfVG1NpE
Di/rpLTcvbpjrIZgsacNVD9BRuTDZOu0whP6USRXuK0ay50uttmf2Sn2E1/cmJwg
9DvzR/JMXSEM7Uiamyqjs4IRbe2JplxoO3oSBEkisXB8BCkRF5Wz1G8EaX9B2KCO
IrKmVcuT5D4sByuO2sWynPeSH8seKqlTTW+rsnqqMc7hpmJwJ4EhY1ucN2R+YNWW
FvKKA+sJLc6iA4b4L5LpD5AyZSVgZqObSSkpjYFlUTjAdYiFI/zIy8DQBsYNPtgI
AhtpC//D3UGLaZ8pK/wFNCn19VWpiOc24fbEH8iva17Hm+EEEPW0uvxIGgDoLNwg
Tbh7CX2Y2rrzl/VPlGUMZcgwVNi93kAbiZZC+DHSu+4XKtpjmvIYXDx3wbN383ax
RIV36eYF6yKOU2Wthlxdpyr9cz4HowOyjVJZv3vZdKIxk3ZlcixDVOZwkC4U8mW0
85woZ7rSDba30SKLQ1dTJMC7tz9rxB5vnRcW74SEgMBTpO48QCGkNipimYGRPUrx
2PJBcuHmN6gBtpxVnmXdrf6PytzB4XZBWmRzX8Td288ZLBrDc7so/0glEXV/qGRS
pxaZXKrVCGXnrfAOkNz3tiN9XhkBogEMQsjcULtvX10iJQxe5wEq2aeDq/cMwmJd
K3LeabNBrXXu02qFsmbPCpIcYGqFkOyY6y3EZlvnutkDjJMzO//k3fmSO9sub24p
i8T8qLs95Y3/S405LdwLRMjbJdQQ4m4o7GTUaEJCBHR5nMnPaDcJAqM032A/iZVQ
zzPsYvPJQgwlEYs6srm9IvWLoLXHjLHD8ZzV5WRtTHRRtCWzy5gzoYl4/DFdNw6X
6/m8ve4O9mTsKptKgl6niYxTMg/hUQShPHXrWdHFcGNe4V7Dggdr6uKAKBNDKmnW
mNFU+51oX/68R8Aw6DqP7RmA/uEf24hiJWV0meO3SU882D0DqWkUizXJEIEpxS6M
mb/WNauwRv20bYw91dZsuzseDXpRWawcG/+8ZfHRNOiDhIXtcs3JgZPVWt3Aum+Q
OXkYNvWR14oC800qxtflJqmtgfbtJyjbA6LGs5DaPSJXLe4eJyavWGpnxWdZkVOE
19MqG9HP1JNQmHWQ+w6A2x0vU8VxwdHjGnXnYUuM8i4jT+FZ/rxsKzG0kctA2Chi
7Wg64edIxHULCHTpyDTJHC6qZ+YiPI0GGnEAx+i/PZ/tV92c3xrX0T5CpKvNH55Z
GsSrO0aEBcHSPdZdKAtujJA213v74XdORDp49bCcI3wBPcwpoI4HIzGuSRoLJ3ZH
5OXSRMDO0mMfYl9q+9an9swdYG5cYAaDfxTIYXxTxhp1HiKp69JxWjf8A1p9OLFq
UCaEPXMXleVduXvqgHg+nae0V9KAE/X/e4VvAoKle9XLnwgiKC7BqChq+x5H4LQv
RK7AeIPWoja4PXkp7PwlxswjmDn1+U/IUPJka0fSKpWa2VhIzSjNmqaX1vWkCK78
dzNqJGvhwLc623Oy066CD1dr0aUxSES/R2ophO2iYT5RPODrmZ7SpIixpLuqMYHp
QI6N+oipNOuC2zP8SwBL1F1FxnfkX5W71EsqT10M5i+PopVoGgnrFLQnkz1Fmr3y
0UtW9AlvtR0yMkTf8EDEuvyOoX1U1n9Q1GM6k6Z1gXVKuejbqi/rm5kAmitxIweb
hYnt/1hGgY+Nawowh38EVkO0V9N3yp9ZNxmA+B/X6aZXiuQCtEkItaGw/Donrsev
bju3a/QeZhitvjkH8Piq/zK5v3FS5xQ2QsS9vo4pj0Gy1yUYmogA3T+lx3KmJ8qw
WL4UWPnJCCH++RSAZg62KdluqzQgLpQMDW6vvM5o875UxFOLK4Z6EFIunc+gLNvz
au37qzeYpeIGTaCxkMfWSP+SlIEArhjVycPo1tbrCSLkr2XA610qtjs/lNPudoiX
Jr44wIfTLyQftwPSqWipUZuefEc28OPBdK6AC90Koa4q3mK9mgO3ZSgrMGXijx4T
3jH6CFG8j6hDCrdlAghKFYleXn1Xt0mp4JV6bnLzIjZERdy44S5tiqyS7agSZ0Md
ym9utHW2tOdBOYXSJJFBXaYgSPK77Q3L77e8Ir3HeyBCSyr/QAtBNqr6u14sw0WQ
CYgJ62BYbkuSfOr1CzB3MewAt5iu+sdP2QRoYNluiZFksjq6dYV6KCBJCryhTPEO
RUAY2uFvLoyQBk+A4acYU1Al7LJHZjqZ2pTYyRtlcnBKo1mu8dvda4QRcZteYTSz
g8Tf11ILR/LkkdnggsbXapzmMTmQ+Jfz0jGyzmovtJLmOjfCfsh8hrsLaqd+83mm
ZE1HXzATVvgj4X2a9C2wFoAxWKH8yybXdcPWBaLxCi6N5XvaTB4MY/Qz2YGZcHFB
zyFzURveTa5M1/QbmPHjPI+ilCn00P34E2yhCHbpiB1b1RK8vci7oFmmpJMlYyvg
p2MDkjE8XBlKDBuOxGG1zgZqp80YkBJzuPcNmR4KVlYSogpREcDAj48+vAIl6Rqt
xcsBNkDD9kcSMc/ZCcfuJpNA+Awm8ZORh/BMkG/q02psBHa7MmoxHJjUsw3rmxTz
nH2haSdvAcQlusXbTZU6UDukARFW3rsyRQ6WmU//ZfDJ4HN6HvgsQeJRPkcjSByA
96DTs0ddU8nzr4DNbT0mrNdXIRQ+6NpXbH9XsavjBx46gIgcIx+BokoNec2Bj4vv
D+q3+6qOJCksngOyA22QqphzwJ8B+Ol5YyoqR6LYmPF8zgO/hy7PWN/eLDUGKDbR
4FjKkMN/8pQ5hRMB+oqTQy7Lx5/7x5zmv+0bLRBLhGi84Q/8onTWuxlC8gi5dfrJ
PllIbXAXTrYZQOj8Ne3OHRPgbOUa37hOikjCwuteMYSrfJfw3MVF6kzscRy8IEuc
EfXoKwpR6NqLHj7jfn1MyYurwpQOHP9EoiiWU3oKSYednZnPYITpDw4X7zzySXsz
9RR4PMuSfRxBxC2ehvlgT13C4lP73voBsZ/PmXzcg+LUNFIc3UB7K8JiWeA1Tw/C
OOyAVLpA825MIoFbS9J8SHgKbIejuLnOkQPMu0NKNtEtLsF5pxPbl92k3doHYuYv
OuDUYSSzZmTOkxakq6nv9r3DiiWOhCQ41XaEI9ZASyzgCTISvHMQd+UxTfW2JmQ5
l839ZpakRLwFsHivuyY274czl4U3MJxdHHNhgsizusjv5mcBmQokEeF9yxaWFp8L
WiZTrLPNKu+JCtec1BCVyxd24uXCDChUh430aJglT3nCHLt26RTMT43ZqT4t8tAh
tOS8+0AbWBTgrr7Dqb8NhEvNZXAFu/7xVbZ/sClmW0o/fYmbBjxkDayRD9Ix19Xj
mnm4Oxuyki1ZHRFsyr8/YQB7mpawIa2wV4+3YnVWzyE2eIMwFIVFtuqYS1Llpdbf
tgdxHpVdLeSqeOVZi29BM/VZ4OD2V25/hA2cpJ8txluWTcFPlq26hZVGYhf0YSXY
XARar1Y9VSrMDaGivcwc1kvDtZssljdde/IEf+JZFto3KKtBwk3DARUdLXUcnnuk
EW3jgFadrRBoIlW2xAmx+0z5w2PpWffChVaf1La2p/+hn7h/o1m04rSdFA7MN2Uf
bHvuPj7DpJJ1NfcYWRH0sYBkVBs5uJjdkw7t6iXPeL/JIAhTOKMxSyLvojh6JHYt
EB0mKxsQyrgTW+Sc5gb63dT+EYgYpGnBG6VI76RURi2QrQ6znJ0qJpZieThBDt7s
xBXpIgF5IRg9ghKOqZyGXQy6/H2yNvhUGjHrN5Yf0we0K18joazuo3VxeoOcFMBl
Faigaclrk1OuhxrCo1qZX6YaXhzJ45uSPfW5MP8cYMcjD2AglBZBjo2sl/jpZQrB
iCx76zIqIeKYr4+Q74qbZPctQEx0EX354qyxY/qpRpwmvwAjI1OIQVatUIMrRBiQ
0hpp2Dk9R7vg14QtJVuQQF6K9DZXHFA2H3IZWewF4e7k77U+ayoXF6F/27jm398N
p6+kXYcx49wwImjKChSxjEDHKqgOhj4ki8Cb7wZcixWDpxrY+VwO3xLanyImZ2hh
UCkT2lkXYFzHahplJXRlI3KvpKIFLU9gXnYA/NSdqhfBM719VbBf/rdjatzbZJbY
iIE9qyjqCISu9gH3bhLHFOvb/WuiCJYHKuSHP2WkV+vt5VAd+ow0wL1xUfgqMZcp
mIvMXOMAnrMxVfA8j4sa74Ibu13B9exINy408N8GMNH4Zk7DGVCzFHkq+XYaLLNF
hKRTH72NteQeDFOr8uOyFTkiJ3hRDOoeYyrGOrp0S4btZuDA12opX6r3zklMyDpF
Po08SsHmkqm14Lqu0tw7bao7e5Ll98S+M6Fw9MfHIeP+Lgj3WydWNJLefpgcVlN6
t7EIiPtHVmlsMXXcXu37yzwCBzIWgJ9S39Fm0cWKB2ahfM/bqeMhzaTs2B0DuKc1
h8215wPuh/VRcNUgVcgaDyLMKf2529wlkNUZrvayiHXlZo2yGHABpTBrLo7Ftzne
o0+REPLYwafH3nbprUqPgIgaDN3oQAac2Lxabqa+0q3AQsE9eJ6pw/4xIyMEM7HO
Dluh859DBtKVHoMHsD6ivv5xkJ33v1zuKmKVEGDc8Td2xo0BGFcmLBTrlmkQOsJd
DWgRGqcBzccnFO7mjylAhXN+5ktkHWfVMnrpCPkXNhxX9yE/bv48nBl1bFH0OjnA
2dTWsCLLM1BhxMKOVZDZ5saBDJdCrfwIYIjlkPOjaxVHGsA1EzmdLid76kErcFsI
qAM370EEtoxUMFBtZa+Ma0Wyr4iwn7dHYDPeYToawBiQVH0dc3QnxmWp9fJ8EbBK
X54uIQOpXTcKeLmqOviPG5TPtcvwKe4TmTg6yausXLnUj7r5QkHWpKH0YbZ1shGX
LRZ9VZ5SBpjE1/ZuVAu8MRHTGSRz40Ncwn/hj3i5XNdeSNJWUUSZQVIXhaVm7nP1
H8oLNlv7XGXGDfhakbr9dFpRazrt6YY+Z6LZCNdWxPYhwppDlJ3gumw2Nif3qP9m
/AN5m8X6fajsvVzUm+DVJE5VLCI141zqLLvKOSaqYFWPl9VtkJw9//dlw1sXSzQx
j5hNmN33KULo14CP98XOfgK8lVWwQjjixqKC8d3qObPMKmqK1hbULEsB/fH7t6jb
2Lk2A9iIIMA8wVSb/v/WMxQLkD1YPxRrco8hPsiTB6PeyUxBL515cH8eq71Gw2ct
S+JeOZ8wqq5pFfrHY+OxYWZWaD3lesdUBQVrV4/YuQv58xSAoIHoObz6JAL6lL+c
5kdfigZMiGnXjsCRHX4cX1E/atYjnOhjYmOikj+5FyAQ2VGGmvbPH3hhjozg47SF
hzCo9AmRLVbFx8h/8G+CmvWbP4NDuUVITkHLFBfhlLa60bPCQW+77CmnU8Xz3MtW
btxmCEzivpuBcS0CkTSZmdBL/7qxydWLlK4nfuPNZXcZzm6Bp5WICpoPrnW1I+Rx
nDxSYUZzZPLam77P9QiRFa75F0PDTuBtaGF3MpMUTWCzjRF6YQioYbJLJyO6eCYu
OLHPWWec1WQIPilps874gOoawnRNp970bu4Jje6lzQc74MFoRMhnZTpbnsg4xb9Q
YCk4xKb0YU5dmNIxSxtT/4iR/Nf/b7xsO40W/Voo4Op4ij4isgbLkw9haB7GffY9
lJKQXsE4eCMO5IVuhG5Cioqz6nFhwDvi8fAn/H2Br+dXmbCL2gyumaFJ/xHZT2Qn
Q7UKM+Afe+h37zvSDQq/Ylg0eXGDM28Cfqsy/8O2uq1jIA6j80y+qyZoebBFb8kV
77dipvucZHnbknwH/PMJWu2gW8mI/KpG6Qwce7dyqsSSybRxsw5G4LKhBpi8ps+R
ZiHlctRe9TMi7IJK0pEgYGl2i1fXsnTnkUaM3HWk/UZLxye3KhTspbOTDQzY5VEv
2k8WBh5rvZO8zpcJL8h0V4u7iLta90Cr0j5hDCe51V6tKJ3U7HdOUwn1AM3DSojB
/dZxCZHTq24jpiYCozu74LZXZTN11HsTeLQBj1nwR0q9X7Tnlbt7Qbr/aqVJSFd/
pxaOUBQn2zkraGUIe7V5oGIfk+zRHisYIEHVI82+JavWuM8u5ViEvI1zJ5puikvI
yEh74pKQIt7VKDsggnuuw1Rog4IReU6NgbAZHfhBnKpEUDEyGADqgbjXixBvwzEi
wheAi5uzb7UyH42wl4DiUnxjfO5xcRTHtupARLlpQpXLWSFrGhfvz77I6GuzKIJZ
pbEzLNgD6dKkPmgEfWQ5EmVkPLOOeBZOJwgYu7+TyGRki5q6AUYxIxPPfeXHSg2u
KoELfJvIMSz3fTaSimvweu8feub81GALJd5Te24c13Ke9j11OZTUsnyOHYm5KKUr
782WlaIhoy1y+WCfOUcPMBtyvLtt4P94JWHFKsoOyndEL89KA3WG00wEmjMAis1p
Q2BvJtR+UyDwIdR2Yqb/JFb38v440oR4ph/kTni5cXo4SfA7vcVsClBdarkq1J0W
AiCbHYjwHEFFzlstC/sIxESoA/5/IGXQGpOx1a6Rrq1NnQ0AS58Jh4EkzT3ciZ/0
+L+BBxeIbIS04G28PiwSS69+P1F3PTzdUXlkzzWZP1GdkSK3oapF4Wt25Xgff5qd
f9EmekDpKVFJHySw/6FQLCh0mtE10o/29oqsW8VkepZljOiih1qrmyopn78R8dKV
mG+fm1U7PlBizvdrr1duNiazDeLFpYzfuXL17/HrNE+RQi4trnLOqekEsN1SGEW0
SZNaTabFw5E9ss1lBtNbRuTW49bOc1/R80e6jMcgRY9+yBQQ9N+Zb1fGWBlqseiM
ua7g/+2juFoOJjfCQXwFuKGRT/M8+lexEXuCZChdlPmoOr+977b5R8+xOKFeuZHh
ZN98ugGvSp3FQWWdlBD9iBr8vUZOgRaydqNtz9rpiyPaJWdbFtJcAqWbthdc+wRA
THPqtv66h8TaUVp8//SoRt57FC69oPsGlUJEr9WCBwsIgNBD2L/w3uZ96f+FCkF+
qdKSCXzWX38zSSCta0eNkWbL+1RksaksnN7PnQC8Gg5sX4JB4lff8wtbdJdirY3t
Kq/BB2Q6Cd1IWQOV/sMDAqtJpPBd/X8uRmmA4n0QvyGMmfCeEwqoJAs4XcA+zB46
fsVhOI5S8rMg3YCRhsJEOnrvgpgT1593tAfUpMjiIpyC15Cwxn9PecFW3cD/XmPq
axgeoeuy8r92D7/noL3ee00yIoDc88pyCOrQApYwdEYXjUfVag1CflkzPsFjidyl
ptjHEORJ3HANu4CTkF88mCAZWIefKj/vsiUaxNbk+rkOvmQfxLZbGyvksm1jR9V2
PHZ7Y0gPoMdMg7Nre/6s0c6lOSszm1D+QSf2+XPrE3QcELAB0q2QkGuY37iOYz55
KQGar/awL5QrUrmJls825DJL/KOtFRJNtOZ5goQ6P25oT46mB9vdaEZemUD9W0g7
4rWnzd0/iosQnBBbJZL/a0BnJP9wjLZgDoZW4mDwacSttb5rwizUFYs5mJqE23lD
DiKJJBg5fq26DnylBgLATR6izrgCTOJWE1jGTzUyawdBhL3xWdASE7x0L5Nlr+o2
g6S1D3KmKWz2ZO/ANvsNXp0dPc/9QqZk3chOwq2ILlapsQtyTcxPXwiKWePWPOE6
bc1CkWYn/cyVrvaeNuKkBKIQ5fa4Cg+ptVDucWZ3b86A/luSzqZvvn9vB2uW8lX/
OntIoCPjj6i3ZWOSq97fYIYKsgHRFkQgLF9s5q3magh4xO+5B5/FHwGpuLvtoy9n
/wkDZwbC/W1F/ODG6MySQ4DszDaccbsPu8jHaaVwd93alpc7bCgzMvniRdEHpzDW
sARc6xsR3Eo//l5X4N7K50CDv/8+edZD7Ma3ZU9eMDeEG5PnDdFjvMExg7WFz6TP
mr7msiZbEc7ZYjTOe0k/YDTC2AhhL6T0RhZNhptQEpt5TAeAHfpmfQTnVF5a3bOk
ePKSp+MXJYlCnWPRbxd3HGxKEYo6j6dQ2w7lWZQKt7sU8BG/7FQdB0/eR2GCjWDx
Q1v05Sgguaxxn5ROxzFmr8n+ftLbPLwUp4iMXaFTUsESTYs/sE0UHC6Y87obMSTg
0zqFrkbyitpzvzL8ipCJ13lG3nkK993au4cOcvqS+J2OKyZmlkSivP+mNo9f56C8
SPlInqW0ey+kWPaWH12MHA1mZTPj1PTe1Q9GCR9Ws0YmTVa788x9OlLVfzaJvBDv
UWkCGCtMu48Yo7fT1ecKpFmxFDING/MuWMoOltUVWuv+Nmlihxfbaqa14McphXFc
eN28jYvl8cIIOhH+qifjQzczbqQtWTZnPX6xCY15XvGv6JL7kUyDCfGWmVs+RwqJ
Of+mmuDZfYx4GHFobSnw+ArWDd80Qh8eEoz9EV2bgmks6nuMWbuSXBvlfdW1pWAp
pUrN0AbeVSIfzjdoRj6HPJcZ1n7fU6en1Z5V+U0V+S9S9pjkCioqogIeDa46fUFQ
FFWxDwXIyyKxhsgek2FgoeZ/Y6mhZmQmfB2hz9tJ4GOG3SnhiGTvNJk6ZxIwScoh
Z1f27BrH9woG8rWOhF7FRkJNvTq4inhoqU9Anjfo7+jbGAsERKlF2m1Jr822ToSx
tm4IiDEQxuzE9GBnJMVkl70e1hTBFRDfDlbmt136aKCZCcjAM5d2wgiLMgSKVle7
/JEV+p4qfSYTiXdYaCIUCVlyHR9v6muoFYjFzCqcgqNYHTtVeHSf3UsrH6QVgoSd
ruK98CKCpEyN2c7Ugm8qJYiclERU2brVDm+u1EL287y784ru3uqBhRIx7WvXayUC
LrVEcaZNQgqSa6Z1wMKEXRyuDFK0hsDF0wSIyFfGbYJKxNVVi7PnxQPqOgb0jJji
0yD8z1M/1psy9Qf1vTFDgK43HbDvIEjZllx5/jGgEvMjQdh2Dv4UIt+mOV8Dz5f3
Dgs9Cf0depbZYQz1gbcAJ4nga/MnuQpN2Rry2Igg/eFcf+is5f7XKjxIpth5MnyD
EE17zgLeQBjBcQhtXoUH4wes52qQ0E1b48rRynBiZ6l3Rtr007oFiN7lmUA2lPlZ
4ynm2qUSitbfc5HcXoPGxeACDj2PrAVDwTgKf+TuNo+l3dvJcz4JN0iOQUelFsg9
Tbef92LBBZZvoNrHywASbOjCPVs7VX5AuyB04XM/vigNMs7wYZrXtWMn9PAYQC07
wF8WGdUKsjPAQ+daLw5ftHCsoZhD8Ucj48hhjFICOnR3LJLAL4Rm3sn/ucrLdxJ9
iC3X37Ys6F9MWfOUkoj7eBgFQ0b609Ikjk5DZgkiARmqK1GrbFOQiAP/PutTv5Uc
H+6+424OMTMeides2J6q6Zsc4cURZ7d0C1tN4xTJwjDKvcTa9Cj3ezI8sfYmtMxj
c4TMyhYJ37y7kNPbhQCDq+9OPs2T8A/7UuSs5tI6VuuWG7x3+WEmZESpYwcxRVt8
jC3FVQXGlXSYZoiWxHMIlTiuA5jB45GayZ9/ELy0RyYi0vKiij38cy9fSFUniOI9
QhH6LDVkVO68aAFlEwJvCesEscB6j9SGew0cvTso5GAvih5DSbdP9wWROL6dN94w
LpUMb4qYQ+AYwbBYLvetk7RKR1ganW/oeYce3ixA12gu6OMz5DI4UJdJFeV0ZtA3
OIvc0QlKIVX5MypVT0EejC7YTbqjlehSNMf6y67bUeP4ap6y1FF3QoEIFppUGdVn
i+ZF1M/XxE2KzPAuyjDv0LMWN+vQqzdE9MkpoehV/R7ORU+8Q1ZNWllJP82UfWSa
S7Q/HoYct+cGmIiy7UPEkQT3nMLKZHOCrTyDqsvFTWkKlpBHrErkbU/m7FMMxhRN
jKRmvJ57Hq230cXez4JhUen2mKyBtey4xlHWc1Hr3XTxKo+pxyhLsg2Sc/Vx1rp2
t/iOcSMjV27N27ZEyQIweM5HnSSLEqkzww5gsaX5duQ3DE7JnsjEHpiuAlaioA8N
b23Pl096EVZRX2gLUyjfaRMx/6RGyrSjhATv3IioaxADSl+GXT7PAwaJ+7eb9YK8
cpLe+Rg+7Qvo+Hd3Ttws2HyXjSYHtiYUvLFLsYYMThBteHRqP/ZoE0yG5WbA7iV7
TTUp1f0LBu4NPsrLL+hi9iWyDvS1+e2hVahTEUp4hLvyt01xelf4FGM0dGJjzfUJ
RJv6cZiZ3onKfpZ007iJM3kBdBw3XXiZtnOWdp0jUZOzAiGKROTNnGNMBIj65Ubt
Ms/P8ThHkLdLWSVSdJQYB9Hlcoo6IpLaSuGtV8qZLIMsuhHJ0wS3bAwMs67c68ov
pDj6hNy26SV4x6Cd2tqewVdv9cjkC9HqZldqed+hPsL5Ga94hlzdU79URK59o317
58rSwgr1o/rgXqNOZ4ikh+7mPycvP9qwlPGbEfu48QghpU2G1+ZVdVnXVOOo5scv
LMSNJiRRVa4BEyeWFW9NAIyQPNktZOCxr/aC6ZMcB1k7OZVVnR6x4b2FDLb6GSzR
kbGzn0R1LUYf280dgjx7JhMFyDCjxZmEs13O23dTz/EK5oZ+2GHhakYAJfDCnO/t
3g3g8w1QQS+zhiDgoBuavx06sURuG5QiC0cFM7imIO0HTPtaKE0vozAifHK7EN/n
7qx7Ir8v4RuziXOhIxL3gmFtfdFIAM3Shb9iWH81tu0erxIse7FYP2EklEUcg+y+
9lno3DxDQ6gpaYWQxYi7u8PuIJ6vrXVugTM+Rggz8kLVCwzfQkrBHhRYSD2HcGkX
ShpdPloMWR6vWITJo53IYeI6FMPq83lJvBGbl+6job+TUsv4mPSa+MO1oPRwJV0Y
8n0ljGO5VNOf0MrjhmE2c/kAo8TiKDqFKIpzykP7MnIE1IdWGy8eoh6cESecT9z8
Dwiswy0yk1voJaHB6cFypKZU+Y9SqNZOB1+Bds6vthWO5G2on9pyYaigXQJcLIh8
Z1S5pqyzko8+5ypWmhmG2+pR2KtNytxtfm8k5JVrDfFa0whP3omPd9seNsFeqCds
36amM6mBrKIxfxKlV9f7a0zpMyhMIdBAtpb1UaK1NrxP1SZ5O/5aJeaMPfFaxvFg
/jyLblV/VFkLEZPNw+d9hqFKeC4/mE7szHtKnIIndhf5naPwMcAQcNPzmyTtLgYc
48llozw97j9pqLKyjXLb76BMHNVVFo75cf5Ze55uFNuE1YjpeBgV7HTdBq0SPSBv
NQdNPHAgKyyoL4Y2KOhpkL29ynsiSRk+R2rIFB+2UCnsaWo8/h4KgQjFnWyyiIqZ
/SgWeQSRJ6e/NOVmdtn+ul+4giyymUKP46kz/4KEZU/cD5OXbNnFlCpEcx0W+Pnb
68MP0gkViYWG4TYmYc7uvyJLrOM66wEuQWiGhKMasYVO5wNvvJHW5qOH6kzoQkQH
tQOU5uLVtmAjTU0VO5o1C416yUbCNOv1TJ7012kibqHLm7zqBpOebQ+bhHpI/Su4
3nquPJiQz8FUMpixRWn5JE53rZoRU8j3xqmXXZ7So5BkxGXT7D15MuIxGyj10dQg
QEr8fxc+219wUNq0wjte0HId+iDrlBGOo6hBkx//H9ti0Xzgw+fswmJaod/K93Vc
eHOnZjHPRb3Y3OSEL7BEnjV+usAjrwrjQ9VJ9Bz3/CvleLMT803c7jdwUCZHk8n6
Q8y6++nTKeCq6llOkGCK+lb3YJ1vNTYVDezu8S/p2uU3Z2hmvYukdHGVZz+B1qDj
EHYE5PkDtDO9d6O3sh3+OJ37XtpuAvAWiODjmtlv1sATi1v5IzKY7Q4J/V+0hrp2
k+E34RmswUPIPJgRSakS2MuEcwwxD8S5a5J5tljbwKBSReKY8tBiQs4QgDbObxfo
j5jbh5ko5pRsSwVbWz8VtNi43pwv8QDlkVpTlLT/A4vrlFAaYSSStkz2BhBxyWSd
l20s/0BeyuG8cTJVlWySYdHwaq4vOnNDwGEKBFJfs3PtRdPf1ENSbUoSM5ZfHUNP
8qX2v0POzEvqkSRs3grWAqHxSwnWfLzUCmPmZ9MFz6QMykWyBlGxC7KgWxPbwdYi
br6/MBYLf76EwogK2HlNh/Ai2blL8/z45ZWIo4HDgk/o3XAJwvBrhGS5iwHSBwcp
0L67sgB1GZazDXq6nOjEg0bfEC00ufGQMmJwA18evDs/HZRqRTnIqqjf4Q4VCGhd
awkotozkdsdMGw0isJS1DZ5jUt+QQo+New2S7nQ57UBRXAaaUVI286cBDl5zox+O
5eXYfRoQP3/eCkkWQ4TJkyM/W1gCOlu5uBldwmpni3qgfeq3+3ZmavW5NGA+LEQ1
Hs4bvdCi9oE9OtPgCmul2Vj4M2oFCjrmmJlYGjdBuYrrAArdfTFFQhgcjfJnZQnI
VLaDbpPK9B6ll0EshrAcDjrEzRrJqivaKBcIXMgAvpu12WlvEIH03mciVsVuQxAA
ZXMkSYI5pHaEJxFiUSQ8hmxjMybSuvck/rkgksGPOSkm5wdo629tQ8cJowpSbHXr
BbHuLRWzki9qQda9dN73lIZ7T57lGsQUHb2NODr37jorGtqzB0kog61AhalMXRAx
5PcYzKWF4D3N2iLwSB8jjs10rq8ESVQv4BIV8Off46XjvOR03jf8qTrzftKkz7/3
ZrPNPGXnhbEd7EVJ1xAClh2jBF9dqQa/XKrwrhw4eFCP4i2NA4/ePTahDWA6bnEa
bwu3suDjW4XG6lUgkiL943nqkRcSq3VCdgg5lKnWZJ9GbzlN+XVWP06s+EEbQB33
N4DVB/RhVXaGCdrKY8di+cAXBmtNf32lD6zRPxAI3bOjNEV5/icOfm+P3R1iAW4c
dhJXFeNm0qHD7t9Y4vF8jGsdpqMzkaRtCb7KV1i2ZShto8VZL9ASZq2u/390MJZr
GUO50dgqrSDcPaGGxSj55C0nK5M+G38a1JeRmCw6nFbzpd5so7BGkwx2WQqP71F8
egSmty6gUZxjaXOjm12I6sej2qEtMb5+5+j5gx9r8VAiW7OK6l29uC2Dhc5NJOWM
s+ozwM2uePn7456+mKMgQTfUHKrRjarZEDFwXOyu7Qe9ssp2Y3B4v8jj3zj0dGDd
+qRQ3BslGhkjslDaefY1ETd2ijvI2GcL4AG23/CeT5ogNfRSQvpQU1Vai7eEROdS
a7ecdFRwm+0Yb2z8cabtBkMWliuzBwXj0b8kQbj8jvjIm/v0+VFpfrjI28+HOLAa
OxqYma0RHr0cr/eDePRRAOvo153Rn/GoQ0n9o52FDyAHPZSiKDNRx4NGpY3oljO6
f/R6FMvTG1J+k8Inqmps0QAPxUsi4hB04a1Ak+YV3pzBDWb75uE5tK+snTxxJy26
Icai+ED+ahbV0AHTNqAsBPo4lObahoKJlRuH/Zry8HZrJ/pgOHT1GYdzvsk53G+1
1ZYQqGMSXk+ZAT9bIE+FM7FIq/KCC0RcsSS5zI4AeH4/pM5flr8hSCmsI12YXDjN
UiveebTg5uw3UeKT48wefQYJL9VbyFPyvSZ8NgNP/87Id7hBxpAixDOuE59n9P3e
BbsZ1gzGErf7xaK95hsA7bUg/aqvy9Qyd60Zn35No0e2r1ScT/qPRR8LmNInn1s8
XHpSuBJeaLEiP9wdfVO+TBYbuPiPQkjkPafqIrT7L7PBQQRBIIaUos0C8rDuir7V
6fXL4eYY3kNejtT4TsA7QHXrLEOFuRXbFVU/hKUHxI4hPxg7jSn0Y15hfQQXRNn9
7FWVmVBUnIUZHLimNMcaablJrlw8OViLf3S/Vjxxu8WlOr4XYHwYd2pEECBD/W9I
c6m32EwhBnviiIjZOJlPyuNXYbT04O1VjK9AkxEZ+o6KriHwWoFXQIW08NbPQTKD
GhJtuky5JTVCx1T853y5XOKph0cq50pO7fYNHZ0yJzmV3ECMyqoU+o2zw2sCYVYd
akNOkmZUFNrnrFaNj+6SRAHvFv/JBBxQfZXpxlvxcM9JqCJZRePHTuZcFbP5+SIv
u1+58FhNB3yhDIChpemO99NAtQOnbmj6LT+hlFIAkzOp1GJPjonGQ3fe8m6Wpf6l
nnk8LGY+sdfJvG5uJ+c5S0UwDLH58Eqec2gN5q6PV1/1EZQXAq1lrNF3l80dDQ2g
TVV6ZevcXORBvfmy7yAtkbGwO6I//Xbr7mKclkjeSzogD+08gD4Ru/PfjYGoIweS
jauR04F+CnMSQnb8aXJYnHF1KgiZ5ojGlboWEFsmxv3Oi+VYH72dyeEWvgfSbqX7
l7CuuvDNXkp40suSob1s/o0TSt60yRPSCklsEPVkycTlrT6+gwsl7IkRlqlpcnIl
9vR14ZX/8F7YHfwNU3xcNbBUNYpCdn8I698jB0E+PaRa2wAW+bIN1NYj3A7pCxR7
+iV8y7zrYYPIEYigzpjIHaABMwp8q/j51mQk8VxK3G+mVqGAPVD53Ib30MFtTwml
vT/dLucQVVi6hN19iMxZiSLUEth0qE8vj5Jwi/1UX/TXKUbq3qtMS27t1xgYauTx
y6zV0HyQvoxb49Wh8fvG9KMzndF/yRpDjrUjei9WssRaqmxfMPX2FI+Okjcqtgkc
3jca/BLjG6g3Aw6yytwoZWSbv5BygwbgS0khhHO5hOZNnzNpu5l0HUopMTge9SVf
MW46DEsu0lVlkUHhw+6PAFNjra2ItDevyYLXSMXneekOhIi0mxYi5/JqhBaVz1DB
4NJAlnrq4Vjvc0ugqSL3ZyV+GvltFNgLDx8DU6YRPzU3GN+Qg3cPj7Gbkf+B38ev
Z4LElKVcpsVhMB3WINfbMdpriX6XbUz1/DKqI8bPC4VRBAmlF21npnYhMqJF7Tlm
+ZXOTvbs2EvQ2xmi16uhATQq52TSiRed1fHLd/YlXUmoWnTYYMUYIt5n0KAnDHU2
vys5YIlUql1FkSxhazjqVSJPqei+ij5ztnUivmLRFIWk+qv7UsLolryk8CCQv89q
bic/kPt3TZgzv8UGNMX5tfJRWDKv0HbOHV68L+Tqi3/CI0hPtgwHEK4LXCmlT1di
bJzpbM44+NtoZrLxLJWYsoPg8D0E9ZemOIupB2GO9lKjCqxBoygUJxzC2qRxwVlu
dronEigRe23HCw8aJ2RBgJcUpmPhwDA8xUaxDSz70rpUdOE/ySEITBDZKtoygqUe
xgUBz1a2zgUHkI5NfCgtmNeTmQ5r0tI1Tp8aDGAS2p4izI8XpC+tmE7xEp7Bk4sD
V1S5mpzm8xqT4xEOuTNHqbkPESyXvfLViOmmKLvNQZo4IeiBLD0XAMm+nsPZ/uSs
WYmUSbC+DzwiB5IY4UBkn1Vr8NjeET5cVm+m+aiTHpr0GDPerEBO8q7wXwcfPXmx
m5WMe/hr3u9iIgJdXWockAm5E8bkeMX/FDFHICG5E5gww6LyMbUU2Iu4z1tPFOOv
VTA+0rRYIGa9/PrxUSyWSaJf3v2VEXDKH8Oa4BxS7ZFR2UVXB0yUhKjpsBVT+aYT
ETWEx4wMeMa6xfPhP2krdmsq3I+TJhCGdntUSRnl/RFXH+Vmf1ySL3RhkFzJ8Spi
9QMrql9/20jUn0yCkddLRoW8V9cLiWaUK1vt7zgUcoVCIzGEkB11b+UVAKqnDoMk
Itj0qN3TxP+QaFqQzoW4LnX8qNm0XEQCc1Rk9J4UmJErvPZUuM94sUCUmjzqW7fp
Nb0X46iqyQuHqTqDxiGK+mCpMAofLx46hRsv/mPjFTwOsmLWhbem6hTN8TNP4eKt
LHgzrlnfBPYIU17vdU8sc4WhXTQsNLf2TgFg33Y77F15AZZqUYj8h2zZ73CiWBVi
xNPNPbXI/9/eAIKFlXKlX/ELVdIr89QaycMPJnnTZyKefB2+sGqFXYef4Z+WCmPI
+Yz+H57oHeStSY7v2Azbc1tki7ukQxWyCVADZGAIiqnuG5i+R2ftz3BKSDicCjZR
WTtCbqBgrj1g8mb0mMTiCdNsBk0aD3xysVyNFJV4N9XPU4F5Xb7mFkdkcT+h+xi1
Fqq0vzBdG4gZXSN7apnq/E+QhtG635qoyBqVSD/5s21NJcqfMWZQlFSO/DYAd5hg
5+KGbZOyoLCi2XpntSlRx8Msc8yjcatqiaCq2d8VpnjDjSIGQBxkE7Sr31perLOD
w6SLa/1ZApxr5/3w440NYd0YMpDArtAZCHdvUaL68nj1NEDexYj5zxxu3h8HOuAI
mSPZXUyW7eF70tH9bgm1qVxCeVw6D3mHeLIoacrKxQ7+ZEqzKiognNdPOptdgACi
RYE4CWgEpstZt3mMMxTjVaobko8gBNY1wcdiLpp19H3gkNaEehqbYFvhM1BZ0TDG
nP5PasnRNVckMuCg3pWR66WrCRgR1QlV7nhg1YK9LEGXEFoXr2xw93P1178nCV10
WYq3RIw+HU02wa1Rr7QjRi4dwTRjlZIp/Cmknnp+O2IKV1r5enaQ66DFFPAaeH4H
cs6OTPXkqK78wb9PGb0vbAhmMw9P4UA151r09IbGJ54XGL5uDTFep0cLGRO9OotH
WoY3OyYNyCmsuI/Qwfwd8ZhLGXSubEk72tn8gl6UUljU1UPTWrIE9LoPUrlgrYsA
xAtkakzLUm9GJUW+wIR1uQmuHpAzPszr8oimtTL6R+7JOPxTZpaKbUad0ekx0j3d
jP2jKOkBSAhH6q53f9HbWAZz/1+N7bZANhTJ10opljCDFZrgwLz0hXiE0Y51COK0
dfqcRKrpngOZeuT9KXC4SmeAv/sQpRQU+jDgdk/uzBXB5kd29KVqPkZJOWDV4cBt
IO1jXoHwsO9oIr5BW/RIDbuxmCMdmJ9WTkXiwLPK9WnLdHGVofesw510gejWXNY+
ILUtNFZRdh1qkegFBgOeiigBINk3t1DDobO0NNP9rATw27DFQvf4MRiolX0KMTZa
S1Jq0dXaahCtTihEIhbp9/0Jp3MDd05yIL332fXorVGAYuKz9U9KoEle68JnbOpQ
NvO3v7f1W5iIEiVtIEN/0LuBsDKbfNierPjKjuVnw9Few/dPVooLPmtLpeV7iaMe
gw0/wc96U69docLebmfEVetrhdSQp87pdzn6M+n4Z3EFSsjSzGiugenUy/VnhCMw
aWVIJGYqd1NWEbuBO1yzk690HffX6pTtnPG3y3Rr/AzOYPAeVGGyWDqi7UqvgcIX
pwUbjm7E/3baYpxHTpKtP3J5YCD8x2dH3eErvte3YfbHaS6Vy9QTPfBMRn5KCJ+9
aqdPoVoXbkMHSzmKl2/RfXR/kyoCro5MM3pLHqR12imOfMALZ4UFNC7plJ2vuiBz
KJuZsKGObe4cEQ9kGt84wrk7wwnEIWLuxvh6M5ZuMqHjoBzx/THZ0hcGGWIgj0A9
I5TIAMer86VKzn0aGgcG8qouwF5GZNQxrLl9qttCF3CafMm6+IoXlvpql4z893hk
aUGTES4/b8XaDkObSt+KrY1vNinl301WY+fersPO1AZvQ3abBJNCK17hStFdZxg0
a3gx8PiKZoQIdyQeYW33jbpE3rCQ6M5Cz/h1VfSAIPQy+DF30l+mq6URMCXHicEI
f9+rgIOAXcY+YDuNFDAhiaB9eSbv5dCGVs6/hxjlF8pj6HZfhgVqmvzqkUFvhsgb
Q5tQL9wwF+meAnhRggyWMVlBOyCKOwj/rL20BkaUELrzOOCcQ18Y3WRWXDnTuGEj
FwLyAhIcIzSGgjHlDekFLW+8mdIxlEJ4oTwwpAEW/QiJCXe2yJv4skJ3rfKICIVO
GSlgOqfEL2m48KA8xM9cJFnWCAJEvk+qfaqjV4Ho/ZZJSlOw66RagCZGq4HqYHkh
UrnJFMTX6yeYwnkaAhbDXkhGNiMl157MN+6RT25QHnEgcfG6me3N0OFoMmoBN+LG
qOV6mhaBu3A/zZVS8FZlLSARpi0zuF+PnkqCO6PdUW8955JmZDeyPH0oIj7Eqlok
gvW/HtV9UHMF6r58xo8hYpIMXrz/BkR5uXgsSZSMH8SX6/y/eAcEArX1mb3yYrPj
mC+fMZLFuyTfC727XEJnuze8/1ODk9gHdD19kaN1kXqA3mEUNglvb0O03i/7rFQD
itqLBGgP5Cd2ie0I05uSWaiSl7YJQjyk0zdLSMHZU7WQp700BfK7ns1rhs9NrFUG
rYOnIaOhojZu1WbyTHsKOmRx7fl1z/MbwlKoOqCV0bU4DUmEv5mZhWttvUtLP21g
ykjHn1kSYeUJhITCPDAc+YDXZfoxNhSed5xY7ziNXi6UTWliwgjQPHp2pUj5IdIt
nF0/P/FH8T3WSNdaeTUOItPsjo/7krW2tAsLJV1VvQDonoXhFLN4Btf8/rAjWaN3
xjSwr0J1ieLoVxLIkRMgb2RQ/SWbsqg4VjpducKHrYE/fcsYv5n78q0+6xjRsfjC
Gk2AhZm2vIudlzK5cDICqAEk1AFoFAXM/M3zWjc6BEgMMriRtGAQUB+thZZVgcob
jkUpIW8JK3a8088pfC5/CLXP5607LImDv82mi+12gEHcDpZuqJWeidl6uyudQS2/
6ubaw6lkKbZenDNllERBiZq8sPyAoOeo0077BxO2sOQHs8fUBWAAZ+u9iU+dksUZ
lNPpemPlk8HsaE/dHrORq5FLaNTXO0SsJgAUUnbjTlAxQ81GK/JW1vWs40P6GzqC
AvsflY5FtkuC7W2DL/X+bH3CeFOfa76uF9I5E1KNcAn0+moZ+JVUNbf4RCIOR5Wl
BlaZJ6cpSgAXpfFStwbK2X2MBTXiPpptzxcxhaiXgCTHFMosENbYiKIfuZkk65Tj
JR5hoFFht/pQaeZUQ9Cw3SXZLNt8WbQM4N9QAYhpXPxqVTrL6eU4t1nN+do/Ilmp
FWddFeSs6WXxcHvDN42OOlibro4lYHXLx+u0YuRrbsdNYBBgI53efgAIVrgI4p6o
5SMdX71RCptfH1ZZ++Ip4XJKWeirCUIxNjR5IJZzsjdCaLMrWaq0Y9VtDjjbPOLE
azcXU7otukFXsmx5eAe1Zlknn3B0eGwsHOrqJ4FcsqrFhh3KB9IKvTYJNQ6m2B10
jJM7tgUsOrGfs27YxyUoPoa9XY9kHaZJ7UTfh0FB7LSWi2ZTUFYdqZgJePyHLSxb
n6ti2/YeIkCfIYXJ6Q4PzspqhpxE8EuRnG5eIDn8/RqfEEfRhjfDKG+AsSBxbOhM
pKOndZPQLlvjFVLhxzbjvcl76oOCkIoWX7sCZD9gAgz2muv0O/k2l7sh+GXKDu/Q
XrHYJ/nOSDL8nIAFs31AWUsg7OsRbAJ2jSBRiXSrTuxjaSL2SYaHxa0zFgg2K3Z3
6EZyILbMD87Gbrfv1Gd8HO/WCWMjePJ1Jor59+LZKeAtxNzaWhqdd7Jq22EGJywF
wte+m1PCiktZMeU6mhkGPy76kMUoLJCAvr+5f0gb1T6jilhHLqvLV4Tl//08LMNh
bYcvvgizR7qFqvl/Yry5KZunRqOmz4bC0Ppy4C1fLKhS8jPapXbAtYi1Bo1k4QCo
WdCJs9enqhXnN3TyL5T2fE7qmUevJUNUtMh00tGEDvho8yJO1rR/0eeugX0nnYot
9ACFIOI5vCegI5apYjyC3bac8AQxkOIzJGucsnB1ucp/EhyuvXZO8f/36wYriGKB
Qg6XBC3tTmQpOVgl0PuPIhx8Ne8FNyUeVCQEFTsr9v4JSWaw3LLriAR3MQAbLIF4
mFK2LE/7sc+dhFcLjRNpnO6g7sDM6LiMFv4c7WyqyEhm4JxPpgKfHleBnMJxTGGl
Fab4cmtMcCDevc8pLmT1c/S6yrYN+rAMBOXFPm1uv1UukzDwjwSR8kdWYwFSv73Z
o2b0ZNug7hBEXLla2u+mvo2MjUI3gwgU2ujabUAwPDmQEW98yGGiiwu9aqog2Fmg
dzZHFDkoWha2fNnS+bvpYkD6jnb2EDwuRb8tAlO33taEaHxL61L6CzghDxianWpK
+mV5TCq1mgriayqjtDXTR60+mlk6SgEShgY1g/7GOvhAQ/bJi8sZG+nFfdqHv2RO
UjbNy/8VIFsiFFnpsgrAS9zZH263QKSlhryDhbyRvD9/pW/EzKgdeuIqRQdITvkZ
6ifM35v2u+Q/HTCV6J63CbRrlJ9l0wL7YaUCLJhJ3oSB+71hMWc6yhEBO95yElDw
D9uOeF9PhHxw691LoMo0+Qbn61aoZYzkTn+x9h4oGisRCWoJv5j/W4ocvp/c2YQZ
nUmxMR+efFKdgPiwAwaMUIhe1NDKsjocFEpCwTiJOxGlovzsX7xwX/O5TjF49nh4
t5rGLQfQDivxA5lVdF69CYroMqgMABb+eAZbl93l1xDKaiC4EwcGcfS/C2/Nog4w
eqlUOxsCvhpH51XsKUCGP+BT5GCdBoN+bj+eyMai4eTdDGUGipyXdyhOGB821gyA
+qgIvt8PlE1IBcqN0B6k2EZz79GlqUe9wxCbwCm1s3tidu1bR/ITyzH5HqDsmg00
+ppiOP/a8jJDImkWo3QJ4jKJv7ZnuaF1rRMT+ehQPqLzvzYs1BUmCfZqt7J1L8qE
fxjMvK1t7zxiQsmtpVTsK6D+C7Fm4kFWu05hypHD580XHlcqJR0YyqFuikO3pRpr
e4BrZ3X2VVuPFlHTLnpx2Tja3xXjlOuqJ+OcpdIKRV2VGWdA2RlAI1wbfNd3/psQ
bbKPOfM5IdR5AzYNsJ3ULw9vLnU5eEnnKpJyXN2aIIG6uZ+Fw6IeGJn0OCMjOUdu
OBMMC/qflV3V88KBPqp55S473ja2Yw/Rt9GBMFPPPjqFMTW+2eW5Lgn3md6ngfsF
76f+FHiXwnmvvgmIScPON7oNTecubAWcG9rBtD3tkSptGDBcDz8C82ySjdhQFrTD
uGFojYJhXA76+APTvzzxxx8XOQZyKm2zGtybBKiwuBARvFfp5UVgBSJhaRFUrz5J
LcjmB3DLlmd71ImCGJfutET9YMuY06reYf7Ktvgry5CCiZYZe1ypv7/ratIvjU84
hZF3+xnQJpRSiW8YNLwZtNzBT21TRzW6U3w/iZchkFXz/4kWUAIs7xdxeacacIUq
A+G0xg6JYnWKyV2Tr9qvZ+QRxI2AJ5wjPRSKzwcrBmcN/Wh3k3FDIdUJ3btB64K6
7xFkfbUHoZmB01D6IQCTzjxgaE6rCh6C7nU8oxFXXgsA4ty7JNDzTCAnKrxc2Wkz
aMgFDJaqZnebJb3ytORR7GCTfurbJTfb4QrM55YrwWoji9KGNzp0DhfldbyB2/ys
hye5QWYGt4MODtzV/Veez5tphGArDNo5nW3e79nnnnYZBpBTZzkqszE5OF7eMl4j
RLL5XWC1oEQbprA6P6EjIvZV+LDYQavrqFstoMTetzXqAEaO5i+jt+AN+IflnB4k
hi0iV52B/Q0sfbKDL/90Mob2mph1Ag3KXtZkODiwrpWVALr2FPSf1AR1oJ9PzmN7
RFpctOQrbQZIMQqrw4C3N96ihV3HguVOmlofSTB8SchaPwGuAIA49a/l3jK9b5K3
1340cSxDpdplqcf1Aod64h/DYyTxUZqpuTcmzh5jYFnQqKZOD6eBMBp+DH+B51CN
dmxz72yhNwmuNNck0za940Qc2lcdhY37mpI7FCwZSGY9GhL7GtR+qS8EnlIrXFyN
MW4vlmxIzz93wbz5WTGH39N0hN9Mh8MtlEaRTxldRxnJeQvab/Glge0fo2O/55gh
L7+TcPkZ2NxkbHyO+TMSuh+h2H9fb+EcLXYocyaXW+MTHvt+I4QUfqDbXMCS5wfu
Hx3nGgm25UqUgGYsMNx44kpQMc2atDdzHl0xRrYfjvqSBSsdPkULkGV20AKo6sU8
bCpbL5791uKKXmjPDworZ4Xn805Trcr+oGnip5xitVwOLclFlQ7epHh/VLnEY+w2
bKA1VxiszUQ9wTL3JO2mtPPVJzFmtdcifyEn+2EGWvAu307iKdlgZBBZe+dVUmGl
OZrCihf3/8NA6Xf2FcDTbPBXFOkDLMbQct3Ko1nRayt6CR+kDy2XiOB0CQHjVTIj
jj8AWr9LrR1l8D7KDChydhwPb6FmSP5HZXprZawKOCMD/OaBPmWfKE72XacU1fQ/
unmIVyge8EisuCua00GlLjBhseVzTcFNNx0lzMJP0orIjZWs0uu9M0SGt9Jpu+pl
X+5ViJYOpn0BdfdBkfNpBZW0Zyg0MF5YRRC/7AqxQvPE/0Cwuqt8JfIhIGPUnemL
+jFnuNk5SIh/EsUeoPiupu3ue4hdBWMDVA8BurxM2lRUEEHz+ZYn+BBvFMBf9VKF
aGFe1ytaNz+du2z/GJhUO3Xm9E5XoI41oXem4v1iPHvMcEEYw8e1dpXVZzuewaq4
p9mXcRxiXW6Gc8RGpyjKTxnjyuBm3y5xAuRhnbjJ4TDxM7fF28qBewPUGq+PZBnp
XREa5NIQe5fzGRSnHi6doF2xj2i1d+v7qH3XLgV7swAAbJDp5vCCFJO5nJEXw42o
n3p/GfvweXk1zmx+fy9JnFZf5IEG3m7woEadVOyI+lxDK5lNdrOeBTl+qdvHvj6V
avqvhTibJY8lvm5UXl9Yxzw71TJvaLRNKAcPiHqlTvExk/MQ9s4xiEy6HCPCbYYT
l4M/1xhLZbnPAPcN/8XYtF/U0VSEq56iINSxL+FtyC+ODIiKos+6rVmaU2VzMy5g
9PMWOUOm1NptoNtKum5+1dbyedkacgouC2fmPchaoZ/agFOT9zKnxB7FjATXBmfw
kpzTvY73n/Osmi11N/2FE86MpAvSFKus8TqeYkvdhgqb1uLwUanDc/dHQWOGeGnc
GeUpXR7HuaGR6b0Ei8uPzgsjiBibC82aOSP2qUqcMd+mnq/HCouMgxIbRDYSD8WP
KRFrIUokhCaMxTSXXGxQrno6LRjrYdvac59i6sSwPTqq/ZONcjwqD6ODXDtBDzg/
Vwo9S3Cr6JaZIKL5v2jDtV4mIylITQ2GOpj6rD/ux4RzdLo1CXVV/F56qXeb+GWl
UJ5WanPpcCFc/1jizx0V0QmuFrXPoZXkPpnCYZ1eRh6Qh3EQE39PH2BJjgw0GDJZ
yIRE4NMum8LMDVSefd5tsUo75gat5ZiViEWYV+FsnCSg477rWvH/boh4ZeXq4cm9
IHzc45I00TiumaSkQDnBgn6u++cRH+Aj2OEt7b6A8zygzw721nkwxuaRaUcG+v5K
JE2/RmQMh85BR1En/xaDJ1KvP0elsXH4r3O2bP8crlG/JeDMTnxB03WCsMnNJCTT
KtPPljTuXoGtQLBGyuc8EawYztc+Knd49XqL1j8gYtUBLUaHH/ecaaqajfiJeTmu
aShjXvfnYA2wKuk67DJPHtnF2nNWLJNMl492ZmooJxC7N3NQ48490nRVNcCf+XdG
rsW1S7PHdubmEJuFVhFZFP0XPDvnv2Uyzhdx2xyYxijIjYHApxcwnRxOBSHmkwKc
7QJf+WVIWJnk9bIy0IkSVqYMapzQ9uw51gSJx+54Gvah3RtvpJ7GLi/4oBfmUFJk
RBtHXwepajSyq5insDJbO32TYW/DDTZ33LGr97jz0C7ZSNdhvvXxM9X4U4nD+CqU
e0fXweDBGztPsN4tDoNngxMJKZr0Z0eTfT2VgBYEyzI/am21RQ7AS9gcwOnQVCo/
B4zeb1eJ/rzaYGkSjotjV+BeZafgwU2sWdl4ws2v+WljKROB6xw0e9/noofdL/1x
GwvWWHIkrAUe0wQhyEkPgFyQdFu0wnqVYPQUTmLEp0FXIpAEr5tmcNvvA11M/bUx
atRna9KugABP1TnVlPAEtvZ7cr7hyYV2qDu8pUowErr3crBCgNnMEJTclpmHahMp
fKzV5SMbLdnm3BQt82Lw/98A3hOlATe+Xk99F/ZvzghW5IDVGdJVi6rX2JZhA5+U
zsakwTZF3sMry+NHFUwzdSaaBXW5B5+Re14bSfuct7gO1CorCy2i9yceb13OoEZ/
MmMrk5TlBBvnCvHihzN9sNcKA9IUTz3wJnzkITY44Bj8aZAam29GaLej/27zGpqz
mHtdpLjq53nrI7loFpyEhyuVe4QaaAxstwnAqz2HsQ4Je4E32xPzaBuGnHW3M/wT
XJHeTKcPbWFHph+eAeX2cCEsaRGFwkPIGhU0vFAIMOGbWoyQWByPJXsTdh5A5h/K
WDTanwfqmFAx0COS86WMsjXBLwyg5k/afpZGEDGzbKf4GfymmR3sFZqfeJEt/GwK
ic26dsQov15nyY8OsEHZKrgsPOT7EMFpX3tj6FuJgmHF1nNndxmonEhGr/mQIg5+
Ki+enOdZK2XsQ2+4O4RoEXre3uqRsF/3x4sQrfM0JDVsTEaPDPMOAV6s/SGr7qda
h3NRQsOjRKzF5xglPRrwNcwZfyzg1sxTnn4yxc5ht1qtkEk8Aj36Dl0Fy1ymIBPW
oXICJhYjLWmenwOb+qKppjjq3bnq8A/v/uIPKMOs9OZZdszEfrzMIQpzTiw0Mj4j
P/nsRXVRBEtsjhtU2o9mf4kD4exo8gjAUmKw3HeqNlf3nFU2Z4XwrtgOZUkDHnTV
JvnqsLZmTbo9RP3AvDxlr1E3+Q8Mfm9ewUcV5oU4Hsotk+qBNZQLWcPCYNG9nHsi
FenSXBdRvit9dqJa3uCb4REDxjBqfvkcH5oIZqhsvxCvi0CnqM3lpaK/OyPdu96m
Wn3W0L0aFPQzbVIPhuDsovs7O75pLUpp79W6VXkkvCPzSiU7m/5mQfcgJvDrCMCj
GJ9w62TL2L2agDu/axiZhQctPsWuLxXVIfZnIoodPZ500gmhuZeP9saZhC8SFGmt
xmvdysgk/UhI3afAk/a0roUF7qaNwzQQHcI6/pBUOvWOwjqZt1B9VBx2IafIIp4t
hW5Wm3RBuemolGBMFGxYAJoj4puJ7BhfUgKxCUKnqaMKA9lZXviQboWfvg3IFhyB
w/SMAPCHfWLBLxwg4WtvSbue1FIG7WUwE1zf29L9oLAvha442Vrdop10oYJqr/Rv
Rj96Mm4VtQ9gAW4XYWxxoLaUF7DtdkUz5CRfzjsPNxfq38rGApYTA7MqVXbzWvFB
1P6zi8r6ylS+vohm7HVUNzHC9hRcMyTy3NEqm9C0lYxaw79TlgxJuaQuAt9sSt6B
gHqEyjaGq5V2p1q63xLsy1tvMECLb5N9eAm3JFSmBVfy9pHzctVdp8kpGtEKda4Q
0OjnFRoYSWCnDAZlHT0wVX+Ka5qKyQm4kAd3uwjU8akYh034jEYyvQAzmuL/WKNG
LtDmtWcAX/SQA97jZE2OcQqnemjByxTV9lzkZtgYUaY3XO65iID6unw8D0fmi2Hk
cerF17bL1bmBDmJ5jZM+UWCQlIU88KDXLV9WoLVj3if9hMmsjqcOPNoiqCCIBGq2
bEQ5MlIJaacp3EOJl5H1ugQRQSY4VavSVapwXisyQgx4wRlcCzZ1j4N2F4pZlGH9
yODex30isaoyjcVdklZlfipEUfgKIXS6scs4kOfSZiMKq0FjmSWG7Dt6hyAdUXCg
a3hcdWc2qxCnkSSeOdnDbeGHEHqGJiQM8mAktuPGzbZXmLYfMyJ8nUkgoydByQNw
0Rlgc5x+dVgCrWMBNg2wkic/7wKZnHbd+e7lIJ/tVEPV/OQwl2nCRzikjwZx2zwo
/RvTI9/25KIm5Q1H85kCc3O/A2fv1FcagPKJpUannw4NwXojLPr+oJWH4DE7L5Ml
dtRQlAvVpRz+PFgn73gk9+WowEHET1Bx8WpkxHYUzwbnbFuALHAIfQWoqNT4pbIw
rEp3m/DG8AVOgcgHMi1x6NK6kG438y+9mp7K3PiJkBitU79qMOB+xk5H5bHKb3pt
RBW4+AcEVZEfiHGBa0pCdt3aMEq5PApVH3h0977cpQR58F2KMsCAmfgJd0sXIuK0
iP00R1t4QZY4eYbXWhmzmnF+M+M7EJ1Lu4Kqujq2HmBsNWqQSoAkGudsPqhJvoFo
YIvvDJGsfnTl9lLL8kKO1bufzccIRDwmiiNcMTpB3v7+6Evbt3dtJM+qmPd7badV
th1mKFcGH0AbBz59T4vpbdyEX8gezYZM4oYdpahi2VTMhntd8z0uHWgoxNemPchi
JKHJNBouaY9+JYyFvFuIlkL/p/BSY8r4vbNzzkbS29mvKuyBBIqryhFDzMRGAgcU
anG9XbXKL3oE9YrFKtRa6PnTyAuA4N6z+wvnBbYHJvbkd6XXSpeDueTZFagUCvUm
DmqAJnuSuQXhDGV9k6oz9+cF4SkioTqWjXoAMf0RRPejZ2fxYstUzhwYpSv234Mh
ggkYJa3kDyde0L16Z55qz4EwrzkcEoYtBJZULVLtkEwh5PlNIQzLg3ao0vyulive
5AYW2srCsHD7n34NZ/fH3TVLLTW9r7HOSmpZYtVRUOY1CyX4xwULsuPMh3kYRYfS
dRLYYf44VYUKUKNTKVcnad2WqdGa/q/ZxgcCR2rjntBn26rkDXTSCrSrqmeTplUj
HYdQcGeJMRKqJWQ+YOTQVxFxrOg+JdjD3XbBhk33swGo31mhohTZWJ1k4HPu/NDU
he4+uuBPaQAH0Cx/VUe9uSOd5f0I4iBYaDBpxb8GXvt9m5zjCxjZORQF3fxxOGbH
i9EtE88Fv5dKxyfKDviJp4Qiwt/l6i6XyIqedAtmtgcQELMeD237Zso4ijDbh7NY
oLQRBGy4KYVHJd6PI9vNrFONjkOP8ksG2fGeBKQbNP4++sPUPqP9Z1Fl5xWuuFkA
zd0KjOyU+RTe1dpKWnLsrT4zpdO5tTTmSDEt5nVl8CgMV+XNdfGm9Ir9zQ2ows3f
NAZ712a/923ysRh5yv6gzxIvZs8ZhI90lPEKAr1cN715bAcJVg10m5SbcL43HMTM
vi8zAsTHBrEFroYK5u8yx8Ysli/UlFJ7Q7BiliZRr1a2KSYaqq7lCDRcu+Hpz3EZ
y6jp6luvFEWdA1boi/7h9bYnW581FSjmcogGLJA623W6OnMR6OTFVJZ5n7kK7ESe
4a1iJEYPLWK5IZJ8K3Z02IgWQ4lzviYvI4jjFM3wQ0qSLuTxW+sbaOooTZ5HtHsG
3w7D3oqyfZpFo4vmhEWUgkXM/MBGr0Bx9TuezZrwdb+U02sXz/PhqKdxbhJu+hLo
7bSn04umPN6401omBSCcQ1g2iNW1fI9MWN8irbD+DK4TKNS18QOWcuh5qHJYlu/O
eMgLnWxHM4OLJt5ZAF0Au2nkpUCczEBAaD1cUu8qLt7SUK6TV/J85muGuvefnpHd
WMAtLxmlRKJRi68DcCpt+E/PFk8ux5aBBINyJRo7IXPFqfAYABavGAM2dVPyxK7i
8h/HoZ0atTtwrkpO2OjAhGEJIFskyqS8hG4ug2NoUmFBZF85E15vA6WfPBPEFTDV
x+v6lb4RJHBcwwwGVlU2JuTxCJ5MyN8c0Nr1YvVLjvMNpx1sR7hfUsVUQnmdHZeH
zT8RYDb61BPSwHXMNTtGwU9xVAUMz64I6AJjB5aW2UTL8C6TH1xtD2Vg08AQhAId
uAsqtRp6Pt29CFN2JjRBcsBSOGNeYJ/750dbITUpWzUj2rrH2BWELm62YmPFqg3W
nDbJIs2WxK6tm1PvuzhGXmSK1Vwb72ZS/gTunX3PZkhBW9uZ5t2Im9Dsmzsi1TT9
hrMei5Hc4lGLIeVNNtiMiZKaczEft4x5AC1iCMIY2AIixt0juelIXHU49m727eMJ
JJWOAb/b++fUYef8Fan0OXWVbwNFT1QFB8+qFRqqbvHAMEvx7IPN/nuDTrBEy9TE
xp7x77sk85Icd2Zviu0z3rQx4AdClgRmKekbWdl/m2HJxHQH8FFUeBS+h2IrPO5i
s1OmgRQHnrOlxUxCpCtS7zMICBTuGqCw+Pl9ipVZlnRfJgd3ZdtAhBuYKIVsq5si
L4qLH+tu+lt/ykyimNw/DH/Jv4tC/CF4udWW2/3/cn7A6nWTf0+161PlmLOuldqt
QGtiectFct5L1y5ZAEzAN3azPzj8++0W43aGONqvu+pi4BDvfKVrOoBIj8LG3TAo
djE8bI+0pRgsiTYXelLlq3oGcKHEwvMvXHCkTvoYlzqlYFJ/XhD61ExI5r3xngtb
FPeCBbR3kScH1JkixZKiqfLYIVEvxLodqWYOOoOPa66ALi0M98o7EnbKzkvPneOd
ETmbW+s2fSJW21MIhFOSSytRb9Uu/RUbm1uUl5EB4GQyjmppEgrq32h4e+pbD/xK
50nT7UOJg56/Pvav4sqw9UhUvbbXccm9ZKYtp2jOzUtPWCy4+yAZQLT7EMdV+DMX
V6rNIUAEwzFcUpI/l7DaUvH3vul/44Aby5fJ9HSA0IYZX/bOUmMhiuNfVO5mLW5I
UU5dYxeKPTFhdOle9vf/VhljS9Gw1h6BZy9fnqbIelQj2l4EHGCyE8IiN6c8wcmk
CFUAk+JgB5LW+xbPDtnDe0vWCRNfill1b/WNgwZOH4YyURwyZAk3QcMnZ5Ygr6Zk
C0K9D8UD7BxcHiYqfBB1H7KRVBLamn15b+ZwNzWhZSlzMUhLqOo/rcAZ7KeXUaHD
rQZBEaUHLJ1KhueYXUXtvmaCnZQ6OiFy1c5rwFfhPb/94xO56QZshY4MJu4FRWWP
TYeytpOyoHQWIL2PpqlfARYAEH5VpPE1JOOxqy/e5Uvu53j6b0n7bRyNhaWgPYvY
lKA1AIwsr/J9bxVn8gKz6G6OIdgzM9daGvOlSQPDhx1QSQjxPu9Jq7sHETqRUt1y
cbRwkI3aaUdY+Vzmbct1HpESUxthyJ1P6u2jlHuQ/jhbaigGSG7Clupt3NszPAAx
pZt99rDY18xF2siaQXTPRjJUZ+hJST5s6U2O7SzNE0lqTuescRepyOQRYl3NLU0c
gvfOFjxiseDYxcei7mR2E5tL/S9HjmVJMKH/BcpOYGSbU7A4ali3CYA9ZrtHpKFu
LC7wo3ZIOsWonYQiuGFgkjwsY63UMmtHxGsiMl/ueC509QYfVEa5BOSo2yly6lq6
DL3Wojzbimh/2G5jSIlJaD4mHDWHDgyJNtgaxaY+DAL9Z5oGF5oSCB5OQW66dmaj
hpPplEAPPwyXdYxvFFopYS1uA0ofQvISUBHjnXDlR3EB+3Yd+h6sFqkbnJLjD+Cf
we0d8HRQ4Xt0Af4RGM5ZGZrWsqBcUcHQ1uFe0mM2e4Bn49k/upApBCwxheaX/kik
/bn0EgTgFxal7zoVv/rP21pHe1W19Zu4OJ9iyLtBBCW9fzZpk4Se6mjiP6bCVnm3
eE6Wt34ITUvALNQXenbdNQBYCeRfV2UYsbCBz9NlDOJoVlXE25aYQN3j8QrTYlfy
qGTBU39LxezZcD7A9dSrLQgDZA3wPgqn4SoetcQKCHULoYN6zv6nKDDNwQVe/gsN
1zRcG+iiYmn4Mwtazun7uCDxOoCXSnTp0TcuvqrT/By64ZipEBQvceDJstZJWkKP
TDxtLH+Q8Gje02BxV+sNZnA6adiaM2afLJ07CgToOeqHquLdFE4EKPBqwPDPyNA+
Q2nWmZD7dVmt+Uknv9vkohxXrzbRgvBW+5OQxxqqaYfBHk3YHueZ5Em5Spq3yZBh
AwojHHbBKJ3PBB5iX2cZtH/H3sLsyYTZCZ80CG4rVKOAoiiGuGvfbsaRV/cSD31O
QyqYxb2d2MZxB9bYkwKGIs0x/i15aq6oL6te+4h4TVOB4aj8vEYQR3fyWccMHN60
L4RL6czP6U+yovt343UOLiHjCG3gdglP9n57OSr8sAtraSAswhiZIa1X0n1/7jeF
aLo+dsRAQZRWzF7ewBHFjltFrOaIVA+VE3qyNUO+ku+F7/sfBKaHqANzzUUE+MOL
VK6oHlCiCCFlmHDQObRZVy6Cb8T2A14mR5CIebZmdRhun9pZnN/WF8Y4on0fiQNY
CEwBFWZIA2oXz70aD29749U46U4t0uca5GE0PVQnPyk8WlbtVvu0Q2AxcrpRhuKg
hPTJRYSBUQTsgYk75ehyG2rcIO7lwYg7ciVB6Pl0/7kEyYpGP3w8BiJwrir7XW8S
2S+2MIMH8WuQPWmv1N8z2LJmLQaYtKXkcrf+ZKufAuCl4fUGoORwBRRj3NzOOswI
m1ZgFWPG5dovIotiK6t7rABbAryxHbMEw+/twkjlsEE3Qz7Jnj7M3sRkL9yORK2p
ndsdZd4JjuYTe83cK/Zj8vGWGJJ0Yz3p31f61e+U9bfTCNztKpmhTyfWiabEyH5B
OrPowMJkz/EHmYgqdIZ1Y5EtLRxnPx8he0FEjFSG2rKZV0bUK5LUrwDvJdAFnbNU
+I0UcL7WERPk/D489xUp7X/pPy2eMzX8kFfZLI3Bpe5UhyCVgWe37B1YrhYkXpOv
WRHnBhqeugWg7hOJgQcQZVRJNns440co1Sz85vrbS1azjxvteDCWJQj2ZUuKn/CV
w5cg10pkUNp5TwcD8+pxQOo3ORayMspPQGNjRMFINmVGEdzwl5Osn8aS7dIOnb2K
6qPLDIGvZQizExhCU2d6jvw6qUZx+IP8UtDZtW5xNZUl1Roh0C8KM2FbxRshQiUh
E1UouHduvy7EqagBLtvz3KGIDdrHiVRffJ4fLXuUbyCGkrEkG20EsvaI9+3GQtkB
pc3nH8rFE5Tq9T6Qy7JSfyNPy5I0rYUP0dTqsYkPVNGYYL61Qw9XTKB1DZ4yJJjK
4ub8K0IZ8iWN5D7oaowXdStfqqYOJnI1m5pWZmNtjLro/24DQsV+VQnb+Ws+ABlN
latHRDv/zScVfKl9MLky1KXAcg3CJq0Bp3iEPh3V2zrtf/U6bvKrQ3V4oJDnbUE+
3GlDGrJnC1j8XQ3idfqKq9oKKxCsltPtHQ9DZR4/fUoh7oG0IE+8UA2jPGkO7+Wh
GUsUtECI1Om3asuyjveN2sPB/hGwRkqvsAjEddB2UIEqrm081tXpNaQ37DLPXwf0
FKlsOLu2LBcB6Ok0mJvoaxPpEJq91qWyrrgO4Bwk9vTdmETC3lFMJ7UKIwD0atMj
mQ7X00+tlIX4tHew2utbVl/6jk8DL4ks/W8LU83Hatz+l0SLck/uGp5wBEIHQPFH
Aib4HWqNAZpzrKT0ePpQPM9GLwJ9+nYTff0MUq2DjlMtxF61p2i/9K3M5JPy2kg7
sWrIvlCZkzHMYASKuOTVzMFNHOSzlyaB5AMbRckbY/9OZ0q6B4h+eWleMRPH2UGI
Lhn+upiFWWtqPaVewKnX8WkyRGNaXxgOg5X3BrD99SGUh0qsy0lNeJUW3rXTXdDq
gyYLcOztnkfBRV4SdSOWgS2+ri3mmTKx6VxSdXBxVS114qW1d5WKwyi/unxQCTI0
ofNX6FkKQGTHFJRzwg1s0/3590m9CJ6B2XBlQ5HUJ1w+d0lEUdiSLSEXc2cvajYv
ieqgxRL34GZ1JaRE0jaCUemj4DdveXbn8eukT+dpq36kUUWkkG5QOv4oowXnL0OE
/nhyShrK8PNpyiav0wyjORomY0A4p9VIOr7fZDJz2ZZHeL1rG75iypdGrbbGKAji
Zt/bFrUviXVlHtAjmgwekBhZVteXnEORUDmeGu8e94HCzcIMwUeB0y2apGiHHutX
yl4HZAL8xZxtJ7D8D0sR4yDo2+M8Ec7dPZ4zUDAcDYaKGTKjTHz/KW2JvG5VH8Fs
rrzcobbTU3Mv99gx8Rxa2yP+2gPeaWiLFTLC06CqVp8uPVO5u3ZOGJcqKb1Ecsir
r3fqtEm/ZQitJaMfLTTjuw+etQInHIfPc4Cdd51VMSg/gZHZeFC6HNvlXzN7XMTK
cQUXLGNEi5dmGAoGxM8DNrCioRZsqkOt0gI2OSL0QfjdexjfBy6xgXIeXxlFP87N
5vNghN+To/rL4A/M8nVUS5EIvvPgKsJ9Ef/xKBJy14Z8yEcDanL5m3tT650D1HAQ
FPLvQabOOUcZoDe0DmGe6E/i+lR9RPKNfd3ubpPBnwUwiwWQtqVaKrZGkz+eLWOe
PlAAXovtiV94EgB3tXdzZLBYK4r44krwNYZLBM9GDCgnLFd92PY5JOfIMQ8InJCf
mQRj+H+Wh8D9QKqWxLElYC51193mBod4sdqEtJlIZ/+f17T7WkacTX7sW90ilpbY
LeM5XIsqFv4z498KLjz6aHJ74Cdydx/k8pIAkVIvfTSSR4cUR7RwU2x+Vp6oqSmt
wKT266uAlwR8nDw0Er0fpkIZwEwIsBqvsvS1iGPhzmhPC1t2EhJzofoa41MttSDT
HOtiCLn0blrBBezdqw21DSPUQPXID82NdnwK6sQtF8N4sYtTApCO/TbPcc5ZLROv
/SVkohTt5FsVJq237rWDCH01YpTxHjnx5OsOj5Cv0X+edUAMz423x9E2iM4egFrl
p12AJMkGER0bX/sobzqzzlADBzSMBMna2CILms7xHdZwuP7nMjL6Pc8Y9+nSmUxM
UccUsAU9OxWWwSUJ8Q3R8qhe0rkjnVSodfBoDlXI5ykQrC8L2RCFM8ugJkuB4jiP
Ud1MkhwREvkj9gVLbTf4tW4TnVHjj4UdV0V4DADrk2m2KjmE4UPE+/rvNmMTVyfn
MRXso/TXynz0w/7JY1RD8xFvRv7Ayd5L2CaksquMpCswSv0bxIPd/KfZ+nf/ty1S
u+c1cI62z07frhJ3p3CTKcfaaEIDkLgTWRDsV9wWB5trGq8E/1cTL87OGM8QXYC/
IWAx7HuECV8Zvzrf7ocqZLEUkUvuSBVpjiIt/W+dLox/CoiHebIQPdFjOBW5308z
UrFTnM703xPzD0rvhnG1QH1COGq3XuaKQLInAxDoxdrkOhdqJW/6A2WPv0j5nX+4
rC9zqGmQLkjTJ1cPd38IBF2FWlsk+BZq+6VjDJkE9npj444EVfkGzo2M/oGQbwlS
LqHWTiTcEN+6O6cmLUP07e/y4rPtciH42OUUBloqPs3ZRiNF0TyVeyfuSmbGs0Mz
/NfkawweGqU7o8aUZl2stH56QpAiRL/stX9Sc+Y30ZOF99XpSpxaMFZKg78amHfA
LnL/z3jee6PCgkSlrksKNb+mt7EOtitNZpoDdXLRnXaQGJ/BD+t83EtwIgppxJY9
GmPDqEm54mAFDHZ1zP7WFdvIIFIXD1oDjSbRkT6ZAfIKy0bQHULjfHS3T/4GT7KK
saCJps8ql15s3gM7VsYl0tbQsrOfLUyxY9yahRVTlX3XHKYnzOD8U54gwW+nUF+M
BIbtdZy2RvPTwxdkj82tO9b9H8aZrTyeq6wjo/CK6dzHvFBL1BMW9BvX2uV63TWx
U1Fm28jDIIIxPdv2FQar8hdkIy/6BM4Xj08pLKDEq4Vm9miBua5WYmMMV5DOJwO+
nAPhL3E+cQs5vjXMXqJFSsSdKcnKnv/VJv5ADCli34fc1xYEOpsJTxU6XZ+yp2h5
qM3N8+U9bkwCLZ6pkqLflDOYDS72BBqpQDowkyUSc1ecvLC7LeqnoOaRI44sYoP/
E+yC4YaK1vhi2AnZZWG8/fEmdch2kdmGttbvkLV+4mbKjYFtNE2e8hlp9UXRjtZx
IXIjKOLq1aCeEnMFe6jg8Lyu4CTHzOtajUCVSSClFn1Svh0fxtHIMq1AsVMcG6aD
b9bdB/VSuxYq7MKJJsQDAulcC+V/Ywv52LjRwZAbdc/IFRRzeeQlUPbPs3f1j18n
NAdmpPJLR5gfhgDn9inemU3/d9w29A1YEZc/MeMUL8rVMbLU6dr0Dj7hF0IyzFoy
KrED7zaG5dXizTu89qEH0g5dgXTrHkW1qf5nsm2EI6NSbEh8ERj+yIDHNZNSa+eL
cLNGthEr3SbwerOEDksK0eaYUzUWsSThm3kPIvzP7//mPG6+bNYPqpPwdGNMwBz3
miGNCETRHlET0phnohuXqrxtr7jwXe1T9CRDnKPCjrwXd84lZrDi+BQ4hJXlKqAx
Q/bSfZeWg8c9qnmaV8aVGAXt5qpNT3ppuo+Cw5xhTJs/bEpGad4VkI1EGRLllt/1
TEJPDXCHt/2iEQL9KbHtfvsK3v5NXK9nk87w/z/1R7WyVFHz+aZaNTJGaCh1M9nU
YeBTZkQXQZRTBukRHmjpCdYHXlxtyK1TXMy3U2Xk2sTL2ekD1P2tLl3KByxLyc/N
nPBncrfFmxjDpaaNVBJTVFC9pKtPPqQosog9HLTVQiqZKaHhv/tUagqE+I6NrfIT
wSEAmTfvfFpdli7wwkRZPX8QjhJR9GfPfbG8y3JanftKKYd62iXTRrxUMGvx9cCD
OLkvJ0IVaLESR24T4tWufdKCSnWq3SdlOhVhpbOVKdnkU/QLLRmR+KDgeSNd4EeM
y7E3Dkrvm6gM+JpX6RRUM2IwZDNqL1/AbVT5wwEXEU2ATUqW5SGOBTJXFIpnux1u
/vyV4L8VMXUum6T0EZVY/V0KvjG9O6YKkUCSqRyejENqt4EP5ICn6EvK8+G+Q7ug
7nDAbS5mpvXN3KgNfbzLlPVFiH8iXSRcxmWclBf7JuJrpF1ZB1myhedOVtr8Db4/
SvmuL6NA2ZMUiSE0kCU+tByxLnEF3dvWIiCzncesPe6i1OeW/ntiXIYI1GLLqK73
S42v8pZBUWgQGS+2YJEs2G2IWdbK74A87WzyD39hMUO0lB128ywOfPMdCbGmS/wM
XLoUtzaHtFfBTXbeNtQs9a3/3tabBbt43nUUOo1hguM9nYAIL9yumabaz5lLzzoC
q66ahLFqfDC5yPbj486srCUiJiW7lFIlMu2TOPbdoH3FAz9OTTeq9AOfK93wz2Gv
FihUgKxfmSiCSrTwbPUFwzY2+mtfDcxVO3Hp6Hhu6a5oXNQfhhRhRs90zAAZ/xn1
x0V3SOCdkP6EIOmhod5UbajlREmsI8JPFPVVX7IX9H6bQWcjQRM1n0C/NCxzfxwe
Jk4WLBqumrC06+MpWW3PrkGIG/DQxssQAyiFePZ8otre7u3kRrVYSYsb0rG9KPwu
Tlph/KnCfBfjoX1BBEKa/YthHmjpB/iDgkEOt7lpRPdt8sd3kB4wh77CtC4/90cD
9hVVmPIHWelKz4RsNWV7VGn/X2gNmTCd2X9a3UNowHkZEoWXiB0LZGHyrpws3XFa
URXtp+0y2Is6mOeC3HuWGbCnF685npjZZMwwJqgN1dlVDII/lWt7Bi9HUhPp8WUr
gdK01MtYUFf9yvIOU+ical4g70rPNoBuqA+wa+oZUA9k4RYQISETLYQnCzsoU3RI
MfoFTpWess4sByP8exdidRiuOz1ryzdfbJigX5RYz2bqEAiaAv22Z8QhVzW89SHE
wLjD+L9xombI5rGsLl8b1VOTeCxnlGLXQovlLCkZMX9/ZDbkHdadhQnDX+hUcZxm
gPOu7UI+S6kEfEMaxKj+yPAX8XxfFYPdJ2hu9IEji9+WYepbBAJE1DNHYEf/HCEG
49QlR87bz0xYBz6OBV7E9gg6ytpI0DzaaIgfBl0XaUVVmWJGTj/1FYTo/NPcJFLI
fR7NQZkitFHQEWYj72kbHsrBteRyB+wQSgSwlGWEMj/9OaeYX+wIyEkjddLPCbvO
mMCn4VUGC9LR1t7N0szwWvJB251C0xT7np2bZimgCCc8SHkeoT/Gchcnp6WvKnYb
kZunYaa/ftZXZzl+gIuH4RmpsynkTlSggrIX5j0gYyj2S6QDIVOsJa9qpg3zNVHx
jLYgZP4VC6zX7cbYwT50BCd0hT8WifVbn52Iz7gqY1BryRwQkjkSeDMhPRi/UtzX
eWNzeyE3tN3YMmdVfRl8TLHpGrv1bHWZTr4wkJRq+dOkbslWqr2I1Hfo1ncLt9hQ
f+3IyK6P8mu8MI4tjlMv1WyCZSI88SW1vqg33PyHtoa2ZkY+8SfaQlkgho0lxhHj
U8HAmoS51Gj+9ILLylmpCS8NBYVjNTJf1zQrufPYwrhLFPhHGwXwdf75KE1whCGW
I1OSseB12W8WzYDfWetK++yq72s/UyXjW2qaVirof/zrup0dMGGxLGd1JTh9uoRW
ewPqBWcoMk1OHn3oa9lGyu7+O3tNHQ7tMvu1w4PDHHVJJ1pFakvx2BSZe6U7Ch0h
aGNYzdC/qb3xhY8FDwl+/b15r+2PKdALS63L92422SggMNjAP71V4aIyP7U2lR5z
Kt5ma/dSBeKVQvzX3KZS9MkXfai+7B0lCVpUqdTDLs0POgKCXZLrY9F9svWTZNHq
/A+qkzvig26yhdFnjYTffIkrVTG5y1SYSkHAmyXIX0ATXaeyD7pNRSprbjWe4Fne
qAfMA+WJZVSs2w/qn7YgD75lA+idYMgHC1dRiEToXgtgPRxwBH8CmbiG22ENjSry
bvO8GLyRSr9J2OfAFkHHZ+0utyETBZ/HKcpOGjeAwk4ZZviDqYuWaNuFOcmkeEkr
HN2wesN3MZGsiW8gpF4oFd1dvTpnkLwenLALawd3003nOxCO6O7ohY9TFD7RIJ6P
rirBN25maxBk6jhRukH5dxzYkhEwHfhHSQboLmyGwEfzbg8OV0LmBRMhx0Q23EOn
Sx1Wm2oOUGS5c32P7Be6y4OHOHkBCTovq6ZDuMWhs1YzXtISOMFOgtBFYNLCPX3f
9n9SdD20wVVcGT7WVCM9xpIuwVqRYAVyMFxHYHBayR6wv0pkkwsuwlnnaKrfV+RV
qStenTCkZneocZwg9ils6ieofwvQNUIvCrv/jm7abyJZwn7bNFNB5zKaSjd2g68u
XqjxEj0Xzeb5QeN5zw5YYt/uWgJuKCZ/6FxKcQFWV1wXFp83/pF/YHXsz1jkqrD0
Knwxk7C333wZFTU3RtFw1QgGS9/7qHGBm3KI7NAX/hcHJaWOihufUCfACAYCyZXn
6Oz8O2zGvsEkDgeCmE4QDlY8VvCepdMbCVd11555/ic3ywhGah2PRFkXzSr1n/It
KSHo9QOuu+9Xi/c38hwJr1PXZngfp3glixg1Oi9VzI+xXiML1HzgMS6uAOsQSt+K
txAEfhGuXVdha6MmkwMlGmqVJM14DKmdeiQlXryGrRYqUuAdDF0ZJuacCG37Q1OI
f5dgF+ojBofoTV/fiOonnzDdRZOELekIv5kYwKF8xCuBZXmKhR0DiNd/AntemRm3
W4KYqjdOicSj7rX/0xGS0SLFd4qX6HHEw04r7QP0jHS3UyUHQ0ammW218BeQhbNi
bvdylz3AHNBValCJq3egWeBbtffNhaLdUXA7YgndGZAhrTsxJ+jgWKVxMpCFeIP0
my5ARXlS91f8T55CPzPFhjevdbn7PUwG+PVQ3ndZ1tF5/RSmGIzjaXiC5wEbg9Pp
fD5CokULH+lV2O1Fl4bJoPQMpP5MOZeyTblmUEUpFyENIa34wY6rlOUa0xM7Ym0x
uys6UUIiu401WFXAw5VgFiYCh2tbw0FiGmJ7o7T0zCPgRZFVwFbJDcBOohgap0Sr
klFXM4NvcrGO4FhnyakDk/7UwfeWWFn/4g8H8rdyi68WoEVrtlxzG3cxiPTkEu0t
w3qtt6wuwQDTCI7KgB/DzcGA3wqvjvT4SvADP3OaiSGXJK2zWWsdEvPxh05UL97u
0Jgq/045SLwQty9Yemuj6HkgpEvechx+kkOLn8pHW8KALi/YkuYZ23ya/d6RaPag
zf+VxIiA1yPsi/EPDA9RtMxByIXwb6o31A89LI0sjMcp0piLm/54x9BCuh+7ZtCg
KEo8dQotuwqSLRhB2YLoOG+BzSWWXGJfvg8ji6925/b+jFs/oILgZ9vL5Yd/wiq3
TFybFrHfasYvW8fEd5+WyX1VR7+DXzGxjoxLSX0xuKkXzDocJJUtvCg/XWLQMB0D
XvwbdaIZm5KoFjL3znXUk6q9t+D68K3j1HzxOSJx/97aDUi8rZ97GzENdtOrA9ma
u/qoUvtKflUxMeIMocIYT+q7zCqwPWWVVSh15FXG3NbpDS7H/rjYd+CdgR64YURk
UIpXD3/oH733qBPs5/ZMm7707/KnUtkRKx2fbRAL8ASosFzeo3oOvZ5/exDyk9aT
ZE8b7o5vSZTMkfCaB223ckrtSdE+hWAU7bBOT+CeN9s053A2ai7UaxpYcDNNy/jT
NcZG8yaIEconbhM2juAtyhgfkl/oC4Zc6pXAANefjvJljvcgjJv50IzrZOT4qwD1
vrTgiUiwmmwC0FDwDHNYOShuIOlLVpn5OI6StF+uc97MxRAvb/FKYzARx7aBEbrv
H79pIr22+xYZuSTONfeIjt0wIrmJky4rTkYJwyG7Z7B2C2JVSLttqIANltoVds/s
bGNUpo7KPUV+XCiXGOxkjUjgSsBtQrr284mS/vvlVRyHJMiJeeCdku8z9AAmlmaL
5nDWzx76Ff+xeRLrs7RviF3Y22VIHH5noKiSs+CV7uA5yxn8uISQjR0fsYZX334W
6KSzvdYkWQfNi87sLugXqU271hxwXqTOOdptjkjXSNJHQVzfvmVOXDrWDnLPJ+3i
tQ9ygsSymOEeZ8VW+eHFP8PjWLbj2U2AHXf6RI9uQtPDG0QfCar8NsFxQgxHhS6M
MGYurT77dPLS1UUgFFSWeyQbBDjDqLQgTYIIUB0/s5841vmTksh9UpkRO6z7nqXY
dZczGMR+rO1eQr0S8BzsyHYvWquMUFSt8HVSIuKMoCJtuW7l/TH+qYp8UYPjDxHq
wmApX/jsgQ2H3KkD66T+cEoBvk4aqyBqzdGrZ83vOpF4p9+E3n5lOI6TjQrbgQ3C
3RfaSXLOn9fWtkT90YMotmK6LOv45+T/jKwejU7iNdOjQHrKrdQMIsWcbsmpvP5X
o/46vDJExYoeBFFqD7Dizbgb/PPg7a2ocxjaoTVztpJEFMxzWP1Uo0SExJMFx/J+
gwuSNgGlHLOnigX9Vwe0FlE4nviDKXCYzOcjv45I6JB3Dzla5VUxzHf48GFCnjLS
Ceau2ayrJmaxyx1pchV1/DB/Of5/pENgP4i0K8AomhRmUAfVQ2P1CJnFTwCKorTM
odu90YEFVjekZUpdc99uxP8H//vK4uCHRhGYNmfZH94AtWGi4au5HUKXySxVFsU+
H7+BtaQ5eZp0d6zcqnaLVxEWLpEamTJHqDsUXBj21ZzwrObC3J7XY4CSCpTQ9/6E
TM0n2Dukqe1yYi9FcM9WS8rZiTuueukgpclDtkh3LS0XVQzCfbz2XuzF4YdA8H5s
jz4hmNV6OKyGF/mwqSEhOVyO6zSJh5C9X+qWwwaEvFxXtcAMAF0bYvUA0R631RwE
7EnqqXUbfQa14leRc/mN+1RB+I8TtYQ13U3TjUWBCJH7473bdvRv0bgnNbZunjNY
gycDZyUwoRKpUHDYjeYkGQ8ha+68yQiAuKhXYbUVe/SbRdWCD+SZsK+CHOzhKa3u
whjXs8Z98X5IcDTXOP6oqXfRhW3BfD01rj3yz8QVlhujScCQ6hOoLj/1lQS1iRCI
xarNGXpxVLJ8mVOUG8uekHnwvg/g/UeZ9cLGAL8APWE6fA0nWsJTSpSOxOj6GA6X
6g3b4onpxNRYB4BvJrNPO6H4MmfNq8FFLxyOZPIEOCab+5O3KI0UkAYTqTqkvU24
c1dspLQPyZblzsTvk9TK5dvebLFWRHVnJPC3c2LaTOZ1DpS7AiwO0lWowYL4BtVQ
0j4zhmBNd22Dm1wiEvQz0tVaOGUhGV7AiCYZOHBH2/ySOtRSR+79Ry0Xx7jTEkGv
ZxBZfRT/KuCrKa1PU2bJ/9o+wqIjp34EMZLIqqDvfZB2hMUH57n0g/esOuBcX2E2
R3PH0nxa3MBc6W7IiBOZvqnvPCQzQ2/fzm5Vjf/fl4XKy6M/wY0eZqE6S2m0x/WX
HwswPYKn6T7ddNU6MeSln8j+M2/dywL//SEMwMa10iFtoe+1G9Y1ltF2XHy/VhT7
+vS9YPAkgmDjpR6uTtPOrMiHt+BMoetb6upo36d7esQJxA4uZp/jYXbMn5/ynp8P
R+nuoQxY9U2dggNkCyzJgMAU6n6dGbbS5dDTKq2vA6YtJEXw4MXjVHWwcZj9BgsQ
SmgIhTXxs7Z4o3OrZRSFo60Y945ghQVKbHxFkB4C//c7MSxekc1AiKVLqrdxa3zq
rmdAwNcs8B9jAJuMmClip+bwIGthlF0Gb3+02OvhHufD5pVD6dp33mmFcBZPa0Mn
XsHOMoMBIhBFp7ogLaZMI3E3iM4o3epXw/eSDnJeg8hZOksgIo5z0ZUTogr3SxLM
FLANsAryFA/TCCIGI+rQhdRaLXvFQvyUDIlhjQqD9beS22wJfFnO76Fcf4zB26d1
IVnN5qZh16EZSGJR6EfnPK3ZQ6sHxF7GipDlFcUf3oxDWbNpSqcpjBvzh6ZMaFTF
aYaN2KbnFs76lUqlBKAB13iv3OSNNoS9HInyjQU/wDRnaKz10G6TyAuMumSFik7q
cDN4mN0dRqWdpe2Hll8bYY0xcPuxcHIousrRAvSQWaiy4umvUZwcj1iI2OM7EhMQ
COccQNSvSS2v767++ho4+H+exiUz37VXJH8S5P8AdWDwgqMJEpdcJzKayrwpN5ML
CL/9F/7MdzHbjF3tLJb3GSY8rQISdLxkkIZk/utZ++74IgAgo5yTuiPA0qbcCKQN
wm+FfPF+yNpft3upUyGNlW+jD+QQ72F61O0BQzf9+3VDXrKgiJD2ysY1F+GF8z6v
wyb9Ec0wQvnoBUNaXmEobdt+rYir2E+Thm/e94dL8gw6zn8Ug/xVgIZjk34nsF3T
VPuz4q6RWY84MM5XbKbBo25zhLB8wDFarH2hutz2TUrliGhWfnmRSVaKMVM2ovJm
CeiScKbjnfo3W5ZxRFfR974Zq9T5+nfAlhVrh6P8WEDDuN/vKahG+fbgUYaNhXRl
umBTNFARc+DLit4/FqPJ8Q1xUXgsVNd1G2Qk1487U9Z/o/jpJX/fCQlHwMlivjQj
ersbSZ9xq9cGYzKO4p1R2Ts+oyT+XfHKMzSMmInPgOnb9WRxSaTX6k9QPhpvOHuw
2fg20T08Q9YXcJKhX/LDZd8diYwFed5or4j2IWQ9Jh6AlbU0tH0r4RY1oUNdHTUY
r1SGJZ+2lk36BsFUg+nOP3dzMGCoTNsG8w6t2Gq78XU3/c8FvjXr48cW5IygN8TF
W5bgzmv8kFCXdc1QkEsBOwmUEngTZJEQt2yq3gu+CNotwOVGQCo6JCIk39SkljuH
J7ty2jDia7bnzuv/9BKUnV4zCYyyCY3LEAq+iQR8ud7v32yKxrOtNj0Rrspzkcgv
f+QSnNbtZ+Ec/UrQn/b/xtex5wY2ceoa0cRNPOYURDEh/fTMSu0Vh/Ky+m4Wnr5L
/C+DeW6XM3GeFyPukgmm2cwfhjhiGBNk4kww7DbDzxSfUBueX7Abnsg3YShJTLQt
HFmG60qs1R4tMo/c1P01U3fwSDixa1d7xlzb4vEUdeuDtZH/r8qqxTEbPr8beonk
fBnmnrR24T+QL7uoeI0WMiXfxqeahMIeBIl5zMAnwKide+d2SKZwYHxR26ORoDQq
P0CddWZygto6/fIZTzQfQPXQcnvwAG3hQxgp1UaVlb3xgwHBCuRu/8gPO5x7090z
h1huuoRr4xIQagmqfeRkawifUz8D5P9bqcV98mCCkm+SbukLqvijyIuq09JSIcSi
fCHZV+bakObxg2emONSOvLijbeHR/DBPfFhr+QTeZB1kFWxcP4TM9rIrVyKHVdA+
p0vQHS/8lPpYhxQTOdVWlmxnuvv8IDpgY+JwQSKurV3rG+7Lg0rqBtCK8PRHkl8X
uRCTiX+GuWbj+i9yIstu2tZXEMUguS3Vgtm9vEFeql94sb+Pa2XiFus0m+kx0STA
lYFboE+Bjbd0P+IKjNAU2B0kY841q2htKVKYwefPM8MfzGOTwtToB+nbpFABBZz9
fTYyBOErAKpYDUK5NKohpvBFq34xwkY7Ef1d28MsTq/vZ8PtM2L3Cyci//sbKrYb
+fTbxRgCGr/H7neHydQrT+1gndPV9M281Fe4VhIBVQJ6SlXB5voMdE77pf5tAYBq
E97I498GZrBxmq+0R8FUIvym8PBNAnrgxR7S8fRd161qBb4HDKllGlpd7lAQVrNg
mv+1zSjFa4w0GAa+W+gYIotbZcyHVFyWlLn7p4YcrkyPfrpSMLmSj6ACgYeziK8c
e/c2UvEtJ4ZW100TpTdksDcRn0SubWkeFaFlBh1GD8zrTQGCjY3/XOAVbB9eGgxB
2qvymYl8E7Q+LjicvzTdqvOvu2cxc8OOaMi3tcnbTr6IZW5HCvGcL49oiVcI1h+4
qnbvQAwFhp1NJw9iZWk/xvCYBBJG/OPuPJsGkloT1rLm4kZerCXxli2mStcam3kY
hmbTCPQ0SKeEppSjzOL06B7atJGl+CnTcy/xlXQ42Znjw8UdlQv5oelsNjXTArqe
/4FuanfrxiXxAfaqebYfifkcV5TIxSk0IbyaelzinGVV8N5sFOyOUBfkqZhXRV6+
4sh3vZ69ELLzwIOAFw6KhrWz3JPG5YaYRcwMZzUON5yKzMoL2brACNYUrCBt30j4
VcOvvDaiIZ9evPC0zSqkcZiSE+5mZFF0ZnKZgVZ/blh8IakUgIGExGRWcMcWA+56
ue2K0D48vqOTPmsrehOrc2vRLghxDSEbe/lb40FJxQUZKQHxWWH4I1dbyzG7m1cu
g0MN62BnyQy2vLd+Z5DGO1FO4l5RnJsas9rOSL6JrTjeMGrG3RxwUodym7M9H/g3
Y1IwWQ7Iu/unxuR5lWScSANc8J02GaxJ/I0WaP2MGjH5tUHEqbSsFfRAWndMLeYm
M5WvrTg5reosDzDqazZ3pK/VEeV+4exSJa2NicTn3OeHnVh4ftCECJD8szX/LfUr
3eKehlbMV/Rt74zYl9Mu0QT68yt/f49or+aNZWbNWYiwnTJSzlfHg76sfKhb+9HS
PjZjf3oepdBS+9E48Q7w6rDXzg3yo6P6vJRz0ufBenkgz13avSEEAbA6bMacrd7O
DufGsNfQ+0iBlrqq3wSD+hoTj1yl/pohvTyP1IEQFECzsB9XK4LkXjmQgxLTEVHy
OQVCLv0Hy2htURm7su0BlOI5vFXWoerNvlTQ/WS1MQ3MDt88nCGSBP9gtixxJ9k8
DkS4so3WxZUppfuQMZG1ls5YgDxlm637dM0UwnxdsdAoCXPzzP52LBW7koqAtk8b
hS5rFOVxvH4VL+GCweZBN1B9RP5yZ+bP1wkPyJGFvrw4eAfKFDuX7rZl3rRrMbKC
qBvplyFMYe0YO+rvDEpbNpJZ0RUuyLQgaSRtr9W9nqDCwQhwsH6jhEntr68gsoJG
07i8umuwlZQ031f/kaWqpu9yjSog0cx6DUW3MBhLjSyRjxi1UclcPovrqJSZVD1c
z2za0kzZ9EZMTgEsubcu+PF0I6ibIcvS5WtUuqGOKJ7W1JCWW372xzfKOH5T3vEV
s6ckXMwfnJAvpHQkEir793ZofEuY+AEX9a2/10QP+S/CEr8duo+rUivqPwKUWgT6
pHoJdaEjD/i3rhLNzT4d2VakJjLozdtFBMP4L3O9OzpYe57yL9FyrJ8lyXZMRU6f
Fgqy/Z6NFcFGVfvZb32xL4y0UsQdRdBBLNlldvpZ1aY4gPqAVP9MJZJrsNy98UHA
P9q0cg7wFpqF6mJy8SrNxHtN1drkh85mY2e2yIXjRnvmLXhQbwlJAXZ/INxfgRYI
3+gQ5iMsaKYTihAqhrwR+LAj06WZ1vrWuPoPvU8bI39Ggy5+VU714GbMu9mWFQJu
SFoWGGFsaso9c4TDEwu9sNVaUo3bZnEldRubnglP/UTnxF1r5NxrWsLmaVR1owim
PstIhx1Gga9gNyf4w8oO7XxlTiePdmUHddRwCrgd8igRRPtmFlT6mAkhSlJVRx0I
eZwwniDRIBls60AJkJd0siKBGCaLH8kEs19jjVYbOslkaDi0ff8sBf9Oxt5xYcOD
QzGXtIz2G+lyIQKruJowO7oboovIJZMmQIBNtQqJAGD9SgmGspmSgL4y7dm1GUMC
DzAQ3clIg9RJwr9vLCCPDaka5jFMWAtcYGcVpgyl4redwfLV7R8u+SfDG6g19Foe
FFekX43DdxQqJ/EnkGITG1EwfTMppzhDwq/gDKuA7b2Yeo/Wez/Z20Xu15aewYTB
u0UgogURYvTtcVBeSOJOWnIAxyjZga6lUWHJlHs0Ji78ChmXsX9FgapJtVGRtA6F
x1Z1vaslOmzl+srTC+Lz5TNOnXtUFYcy46NEhVZgRzLEeiYBeOe5GJaZN4O5QaNP
1KGsfDYfSPr4hoEOf6W4fwuR1X48akxmkYPsWeYxi+bmPkfBh/2/rBmC7Lvy2lML
HflWrQQhnon9PyEhHOE46GBac0G9b075XzNlcj8PQsTsqYu/dlLZUOHtV4QVbAMI
BhLuXWXx1NZpp7OoweJFMo60AL/enlQEDU3NIju2agLVbbjj1PwENH8dChk0Mu+d
nkc3eFlzy2M+a3TTiE8oJpx+p4NUOvf0ObJoUtn//mf6HQLRV5vmp3tkyBTrwmco
Zqyy4CG8zRJvMqOlPPDOZJ0XbnmS7SRJwjmDrp6keDI4kGGBXlm/VFTLKfM+o2CR
kQkYAcpSLlMWviCf9rcXPdEXaXFRsGlKWC95BG/WUDj4QM9Xjhi4afl+S+xV6FrS
0pVfwhX4AOFd/vMXMKcv5etFcZfvaFRwQBWvG7DpvY9BJ7OgB7mtSi0pnZOtQKQJ
LbDeDqI7ZFj5DdNvLP1A60yEPHe11oBb4WrZ3px3F/VUDO+5wKExxfVp3PXJQ9go
qz2kzZtdczg7CVf/BQD0yG11aeGqYBZ6/VzB8Mr4vaAnyUMsm1wNyEgseZ/j+idY
BVb+/v6MI5fdP5/CeAPWRJqc4JB8cDP7cVKWMvs0OieDNAojGSIH65BpEeOnENa5
i5F828NRXUZy5WyPGpkdQJ1EK3Xve0BUbIynWX4P/UNgUKLApPfZDd0SYtWjfP7H
399JMXHuMmX0NFNOX9sLbIKtS99I1LsIXJuKWTMQ7YUoBLH8qfGgM2w+TOacP7jg
+TV8/UN4JwKHhMh1nVfOnhE519Ew1GcXEpke3NdpbcoTQdfYBpqV+6mANvbKDUIM
ofZ+EWhXAHQrt/IRVl/F+Q==
`protect END_PROTECTED
