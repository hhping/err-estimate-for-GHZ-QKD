`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wc6jJW1wYWVyGFNhwWScJT5I4GCvO9FLEHI7KZ/iEI9mzitIvbbCx2WyBqpQr2NM
ykjkFspuNu6xnUcxE3YvqklwZMa6ap1dH2ca2i93ELw96Bq/+ioWPajmQ5SF3/S5
fT97Y/gx3NDrAsCEVRw1rN3N9IGGKwak204RGL8cGKxKoSbYYXBXBaVliU1fnKlE
FWcM/Cbb+8LF4TBmFlmKhGLLwD4he//Y8iQiZx3fwKl0WWHLbhtGY4tkRVT4hiP0
sjM2wS1HuCC2aRGQ1LcCFWSmQ00iisZrI391UqF+T0LsUsYQyPXGruC2t2Px6WTs
g8C81SSc9wEXYompDiwQl7/r19EDFD5Io3ezqqKbNXmgjZ5PrGmo0cYEgqrUq2Op
yhjWJBOynW/BeObNa3kHnyRgkFwr4Baj11l4scYFYgIOwPuO1yorkRRXjWvCatX4
+CmGE3ElTluEF72iXiPeVVfWudXPNyULl/us5oIZ+k9rTJlRM3TBTndJZl2s2Xgq
xndeXqGk1xtHWHqqVwe5i108Smv4pqPIaysHPqohtlpWfuuMnE6JG4PU3smLUwet
39A2Rdwy04r0e/PcDVA4LXrdi8NHzkAxdMdjPztrBzOPk8bZIoLeIOf7mSbkmu1J
CXOiUio+Iu32tD9XBVuxpL1g9Qs1rXZkp6UOkkUPhVG90r56NBHOKnk5xx6XEzXv
OT0zgCiA0b6p2/e2vtM3LqfYOkT2XaDBE15Iz1EgeKF20vR2pesr4gE0k6AOUaQ4
3eBCpYaL5P+gitOSLopxQ2KH3RAmSGLGyw0k4rKBHSU=
`protect END_PROTECTED
