`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+hVcrMfyN62BdvLe8ogYJ5PwTEGfGymCmMjklALIIW/0ecGdY4qU0VW6iNjl+xf
dHniLUTxWCByRdlHTIj3AsrDEwJWINj8DZUFms7Slt/p2HOTyjf9PcZOxqXCEwfn
CVloICZry9Ner52O2yxS6Z7ues2CvipzkPZJubzhFAn/ISGacGCPlw8UKjE4fZuM
/5TUI5O2IazRYyBUTzqdnWCpxQGqpatZhDkgLZLt/RCB32wVorUnA8tG/N97aXZr
Z+w3KXTlj7pe7+C6aQUwXoKUzRybNu/c0X5dgCDP7eoAgDrH4Klz33s29JFNLjEi
UuGK1vK7uA8lO8jaYJjxJWsNmYGXXsZSCSdfKgjUwicitX15OQQoKQGt3CdPE/jk
Ohmm2lu8zQq9/hZ2Xzs1crOrYsbEEvLwX9F0Sy+HrvCIw0vlp+TIxMUevkmdkFUh
3VnO8uvrhCeHJvQspTAcsjnIZ0NxgB+j+52Bo5ySEYkjrfahd3SVWKDSL50bZB1j
Ou/3lBFSwJryYYRaVtbl+WZItgPibmDCCektT2HJW8ATCNGK+a0h2ZD+MBwYUbAb
tK7t+v19lrDgz6x9zOceSZac93fLCQHf4bwd11bHl/v2VRfNIBsiDTfSpvsFzcR6
loUX0eJvKvXa4BxXGx8/g4nEyeb+mLyFJfkhJ737blOH528HPYR2ngP80lPZGDmv
WOTK9OjbQf2mts+COoL7PV4D1A77f82FCl3n6CaO24g=
`protect END_PROTECTED
