`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qS+nq+Mo4q3wvWjES727J4/uM1cNbvYEHXgK1jcATdlDHLJ4VmXGEwFoxtEBH9dJ
T2rXKN1ugjgxwGJJLzCSIBr5ic3RfB6Fybp38PnUAHmOA2ftDDLecfEKeuUo1RsY
ijwR9lhBBwzjoY+GaXdVsEEttdRS+Ep/04sQil1PK0twkU+8VQ0cD4J3nCk/8bdm
GlRNLtwb3qSZca7CaSU009mcbHZkdubI7mOsHnDRr8aKBhbhB7eJPixkPx8kINdm
EDkEDLQFJCvsMN6Tf4NgpN3UqaoNsZRVdFAuz1v7XGvqZ5jCGHryxnmXhWcu/z77
WhYw9dtwr5zrFt4Cpk/XbXMluQQwp3PIaer+bjyJIoUHjOlRzbajRosUl+73TyVs
OXDJtSTk+L2jsx35toBce8K0yZiKYT51L932TuhvNd3ZtYnLnuGbvgXRnUYXrtXL
NmY8wRnWOVf2YHPAte33Zkz3hiO+rZgor4yrMqvB8RQei0+1CDBaHomD/OqPnUlz
b7SkNLucKO+j93tkuTAWlawvK+5LBEaB0p78dr4465TZPNxcgWWMxwKq40Go1I8H
ayIONjU30aVet9gIAIMAP3hvr/Ph9RY80dY2KS+5wsRh0HcN2gkv7n+qsrvrw+NO
3zNavfmqymVI8m6tWigxvxnNbSiWkyqPlqrrh5Bgi1s96e5nOWFNNvTf1AqAm2iJ
hNVSfvzkYM2T30l55vCahyoeuUioBPAPrZaB0Aq4ukvy5TX35g1dZZ7q4iKYjIEd
Z7ayCtzr3y5ebylOg+nIJzXmWIk7nRyFOg1/VzbB5wia6R+HpjHwrgHYVDuAZX8z
EQeJH6tYgq5BtfLc3ciu1vTIjhmm4PiGkmNgs8eSKUmw7hjcvgYHn8yJYK5qz5R9
`protect END_PROTECTED
