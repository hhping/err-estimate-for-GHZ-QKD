`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbrG+Ve1gyYgbknxQo+yGsj15O2dWviYi8oX04SHv9/WgbaHwGM9tNrTv5efN2xh
bfUsHENCEcPgDQdc2elURoqkVELYMje/3LsZaRCl7akjm9fpKq/WH3ION2XBMars
CG6BJXkE+4EfdZbdJUYWSeUCOccLJoMxnARu8pwNa3JmAr+iyjPPRTiwrV9cAvFa
LCAan/SPxwK/bzUhWduBpKcVA3gJVpHumMO6Huru9ON+ldvOTzKPXCfaIhkne6he
rO5A2Rq3iARWBRiYcLgOKbo3vEQc45/TAfBXT+BZ4avXS9b1lxn+DLl51xcVV5gQ
j9e9HuzfsJkZZjTxL/OAOiimVXciX2wAe6OyHdrHkowfg5buU3Af2OSjPA5aM66F
54wEE9QMSc0wnOa9UWOtTokPe+yqwrJzYHQS/S1tRVqrrN08qUa8mWTnwLwHSg7k
ZFhUqv34MDkIZc7AVIyDssR7+LIjkUhCY2HS6IG/UjmfOXQ1I9GXuFYDOR0wuf2T
8qgYslGfbNkIGd9jD+iw6BQArO4RO4D9HcMA0jRLIlseJ3mAYlJL0ij54/hfFfWl
TXoJPQ9OOLU6awZcXU5FzzXDmuDkPWOchLv8iZN0FlzbYcQnGnLrjGgyMzY8e5hc
N40cu3meM16SPyeESeYJj6Cou7/edmbHcbIP7sXKLHfpRHwR3JfXaH69zbgZrpKi
qjxg0RWJ9uXIK+FEQopjnp+XWGVQI2d9rQXMtqyIfwbsGF9Io2EvX3R5DUv2yNm3
H5szmQD24k5lxu5bIm0/POMbHegIvVXZ6fVGKA39nmOpKpYS5aBokIH634aJz94h
VNO1b9MOfNhgLKAcw9bWmKf76TkNtaXYFnnwxlycQyJ9QBH6vY/McjaqpKGBFNUR
jdA0zvooFOnjBfbm9tqiGswebg+3jy5mMbOcQstGRTjpQcvSlmA8WsZteA7fBhMK
MEMID0h65flg8BIyzA5rdUkprKeSXGI2Y9vaC9qdvKEsB3I4GhDDtQv0dKvHzSKQ
HiKetvKnFmYK7C/siOSey7P+wuP5Jr9gCun9v2Bk0eL6UuQek8UWGYyLjzPLvF8V
JG3dL3GjWp+czpX0ASPxMuVnupxtMao2a7Wu+2TOG/YZjXWynWScDt70n29q/CGU
Y00C/PRHWl9iwj6VXN6LgryonFXJOizwYChRRo30YIeb87A3jOFROxY6/HjFgI2b
nr4FucMUNGR1Fw3hlejlvjktocqfb6UbODzz04tvgZmUzKiFOJLAsn0qWuUs2nwC
ZJWxu7VZPdAn+S+jnvs376CW8wk/veccorLj5Rijh4lGvHRDepoKoxs3xqbmngUN
e4PuO0DgwPJqxhsvWQg+zUr2yTELx+zC6eIc5Z51/hQqDbW5KRIKLmJXF9JYaQgE
OwgF40g+CmroO59i/oLpZqll51H+sqry6Hlnt1i+eay3t1itE35cDY1+IKVSSr+v
lr/nSUq1/PrErXkPGLkh+NgFjUJi6wN3mlp9U2JFmwfnv83q2/DeJUKRr7TKemkt
loLZuDv9LcffpgbVRMsKjOjyMat72s0XG7Y+eSQlpdAlUxn3p/kOfLDA2Ztm9r0Q
V2aRRl1tM+iZe0fsuFucwE6AM0/eVw3dv57UbPun0EmdasNkQr6W8u9eyfBnaZAQ
Mgq8w2gUnTAlybk+KAyrjTmTGESlZVnRFISn1kkUFG0wNI/Rrni5DNb2SWebDbTd
xTeFQfyHmNrCjQvK9ONIvQpyQobYVBQt4yp0qijxPosvvBfdw8zgLVaTQAVx+kcm
hT9NGCfXZ4vOIEHTQAJLo2EwLELcrApRYk+5Jxm90FEvaj/59DU4g8ddEDqDwWzL
uGcDlEkAvhDU3qeck+942w==
`protect END_PROTECTED
