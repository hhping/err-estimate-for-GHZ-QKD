`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
862x5Kllki34DdEI8G93GQ7YdV98d6kPhmI72hS5Ld7Ebkiz/AA9wAP49oxUdHfJ
0ZOVSVM3uzNndGlTL5zeC4VLtcM6CXT8QMWuINxaoGNG4NYKNIW+245Xzb+RwP01
zsFw+pAjVC9kiMQxZU8m0lWjlbM8X+jFF00HQQb3Zdcx4LfZpwTY2PvD18NOeiIE
AdmjSRiGzfACPS/Q3y7387/gQrpFwu5hMBf76VKFfBD6p9bUNR7FtLBkuZioBQYy
hX7BZ7cfJHQrzh/1v3QvRzD0Ys57U9Z2uPxu/Wv8pB5NRY4HwiBVmkFkrPYTDdR8
2kDGg4iUVJDfSZaXkC7dr/RDzMiSacs7UQudr2HMIf5XtCgBgQUrynKKedT+iIYu
DCwBjSU2ayNoRO8RuvbS0xRoqh9OqcE7pD4IHsyOcRjciztrrJRuBwy+3YMRlY7B
k4oVlbAu8CrjK1m8iogtPfAOzjmKyfIntwFqsKQkIDMCF+Q/OKmHX9MUx+MimF0M
DoXOzQBIjM6UO9nRwH2vAW0eNeiTsAdXDXGC3CujHmbfSF1IZF4U0YT6alKUEgVm
ywWe1bwtEyOKHAWDrT+quRnvxZ+mdEYekyLPmw0Qk+bnFnRr7JKoNArZWw8m0aEy
v3FM14Lbddk0XffO2zNS+kljFZiRa0qNMbnq6SeW2Ga3/4onO/2VTJxfeMpbzE+S
9/z8yWSzPPZrvHTSC82JD097MUQs4A3i3ekH528cj8xQnLhXPrus45LHEsAtJoVz
u8jmV7xzA8Wsz7K3tSDEiWcf2IcUikuI8qeW3sqBJQ+bxXu8xxYpvcADw8mUEsEf
3Na/811KYj4x04/XYFh7IA==
`protect END_PROTECTED
