`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5J5tx5ABHsujzxn45b/6Xf43hHAmvQeTGWFyGMGkSbhUA5wuxS+JdCNHHLPN5JU3
NNJ8rTyYHUU32tKiiV6nwAlRduAMl/hD8OJOC25mrVJs6oK/T5fwoR9ZVzxZIA4r
NtOZgB2VJSJjhiTJmrMnPwivzm453qsCM8UVU1f4xPj2OSAVqnaeW1MsKrz/JBCf
a9HbbQIRgdga6hdxzUkcemVuIcUtZvyrXsT6YKqfNSJRYQcnQ9pCXeLVH3AcEFdq
3X3ocj3Qcq804VbJQG89ksQoC/0PMg3sLszMt1QMhOs=
`protect END_PROTECTED
