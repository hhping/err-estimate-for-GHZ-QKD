`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJNNBnUd6I4XQLtWgWVa4CdZ/xn3b/EmjR9gH5J5DmVHOkvORFaptN/qX+ZU6Alx
WoB+zajXBmLr5lpQk5X9noLDwHfcRSxjY4EZzwxAN7sP8UmkQqZsu3NOdg6PhgQs
52FamJdgJALL/WVDviNuoTl4q+GsUOnzDKfRv86bzWaCdYnWfNkSGEbGUjaEnCbe
hdfBvI5s3Y+YnNCnvxc7dh4evD+FY1dDHZCmStpFFxi7RIY+floUC37ok1xv9OS4
ukPbtbn3YHz5fXIHajFz4sR4dr4s+4udggU6jVncmsOlrbeIHxP+WNKE9bwozuHL
WNR7P7ul0FUaNFdgjWzvBcodqxUBmU0zB8CuHB6g2W5W52JRT+3L6Ogt4I4Ga24D
M0+9FHbo5kBiqoW/tw6zKYbcbRwk3izQt/cR9iJ4jC2ELcYjKbB/J963fccX3/JB
JosWbWCGJTOlPUgZF8u8UmvgVjCbdFoIFNQ0wU1Fi3qcN29yeq+asLQgawP1kEB9
PfnkZTN6m1T6l6yw9ffW7Y4YJtJYTl7b3jkss+MAqEdCHmoMUqy47p5FeMMBeoFE
AUE8A5wJ+IUORlmdQ3G9wFOye8XZCBDef/ugR+ocSSXwMoP2ENCeAJmnCTKng0XP
bEfApkuAKwc2DXErnQJuwrMq1OWr9Gcnm91b/Mjf1R7mNAaWPfL1VmN9H6t820sM
GHEwOLy2kz/opHU47XPDusOOnYEaatcJo7MP/Q8srdvoP7Ml/V583N012XapM2Zi
aHKOME5g24MSkZovseePwRhUwU54VNlh/xke1Qf/h7NdmJpOugmfGfZvoB0HzupP
4oAGlIB4MJIcQs7X5ap5yjREu24+sI+wHLll0trtXpLJPM4R1HDxCyp/oarRDJBp
kZJBJQ3G6YRD44SAeYcz/ybNtUTxBpZOgqtFaMn+8xB/lWi+KWVX8pEJmSkDV2fJ
OtwNpBANF6LyJADGr2bX++KxY1bikl3U9hLt4HcrJfA=
`protect END_PROTECTED
