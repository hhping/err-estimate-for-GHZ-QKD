`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfG3Schs7RJVbr1p36d2R3IE0QaZ2Atj6oKa+UfxNQHFoh9h4wWqpnaDuD7/E5r8
QrNaugk6uxt0KFFvoSOxaBAO9WL4Oh/SD8M69t/reX26h3yoPaQqlWdXBff0ktqa
Tn8OMIZKvst2e3FiuHUnDdEC3w0b5ETcChBkxwHdBxcsMw5mApRiOoUK99IxF/4+
P+gtw0xEU6zB3LtV/Z2PFN8roan1Ay31bKTGsSNxceNQzkHLdD3LamI15u1BDUVF
mJsH2Bx7Uuhd0NghSLaiwOg6Olcy8WxtYMD+q0XZfZm0L2yfyb3jixlFdNSNDjD4
Yqd60z8fufTIxsWPfwCr3w9xqkc9U/yKCGZ2SRtlzLfw17ABo468d5c6XlL6YrAr
jGNEIJEb53SWPa5e3t4/PSJ/ZtQuj16SqUivsd3s5iQ0sr09FuC0OhN+xTSNM/3j
lQaDB0Y7aXVLlLqwAqUrNdpPy1YdJALMpVmnw6/ywjrJ6JCkXvb9p6f+VANSh036
2kY0BIcY7aa/LJyEisFk1mxerosyCPrMt8biZ5uiM2cxIPrhrpJ5QUFT++3ojuld
bRQIrHoUnJdCQ93WJrIcTyKf6g/TPZvhtB4Ou99QL/RNhxviDyTijo3qb5ZreXtT
p+XFvSm/BugocATxMsp3xCjwMalhiCPeX3IPIn3OkjPJQlx+Ga86stABQjlJY3hc
U4W3bgxtZN/BkFcMhsv7tPwncPFm+rRUgHSIKGQ027KhcRbDqo4vLxg7JU8aB80A
Jw6Q9N/DFs+/6FWs/e3dB2UzuCxXWEWJKxDB41IBEgp8VX8vBoyn0axoGQZAKlA7
s1KPxB9SysnJgsxMS3k0+uRSvbMEvWIE2sIINHoTcNQB1hW4aLu1Gs/SdS5/8Ohi
ojDvpyYeGboMMBrk597g9KCA1sYyEEfR2W0l0m/GyOpLIVqsteKqTSP4NUO3rnN0
SU8Or3xc9qZNsIMiQOZoBxKAu4I2iw3xuqmhBpMfvP/sIWcuHeYuHCLxcyRxo9cA
hZjMLj32cuaqMw7wLnsoRcKwl/sJ81lF9NlV0WXJsn7oaeVNLYfIqfQXWHf/uMfE
mkul445CYLuC9ocN+xWURD5uLR3w77k1yufC7DeL0uRvLYwQgSDf1Zkc6AZ2tcf4
mQlr97Ck6BJjkwnE+oovz/tdSgHM30yiCvWKc/MX0yLUigumjiOx0NsuVadCCpmH
DPo3J5gLkIJoE0RPbEOBZLup9J2uEpQ9oW1Rgqbx10fm5p5n+Z7+n7vgIfa91DLG
f1l/k3cjSbQJBoAJUoPXij6yYPBnDJ39kr3FNUa+0go=
`protect END_PROTECTED
