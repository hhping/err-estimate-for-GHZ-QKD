`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xti/ooJvpkwcTIrospV4FoRDzfcto4s/ppY4s8nbaQt5f6Fra9Eyw1XdeFpGECph
IscxsbynTFlPOMnZ2XVl/37ORLc3r8oysvcmdv1tOeMqCrve8cZvq3qI6oliPlFz
Oq6ePpk+k2RlELsXcpHAVBqxKcy9qLNjkqKIMHAsekulQ/CFOhrRXrqDkwA3EXnj
PK/gc9+fHlIB0VxsA00H3+zPPuSC0WInGduzSdtRr62rRFcy1nksFyHk5mCZsWZR
NSCUHepZO3Cw+6gicHdx3ROjBYuh6nB3DRtgH6K1okBiNSaQpk7K42c9QUWRrZRt
6LAMI2cXxYUl3AowczpG4nXa0Fyu5dqxYMGl80f5u6JQNfi1E+jFY/Rkbk0sBzAe
KUi4vzlBsn30i8pksCXOMaB5CUWNuYWW7pSMLgd26mWrfCby1tbTwcRqOT9U5/Cy
aN9W9W9KSQRSIcbP/LTLs+LyEL0xoYBF0FsAYRru+wqvIha/UYLqzRd7bw77NqrY
xD1AxVX9PdI0PRzI4yKh4yd0LDD/O8XyXEfUeu0OSmO+TzK9QaHHtDsN4bT1pM1h
1//YIWCUuuE28Wc4YEaOyzDh34IVceeyTLM94KLAiNzZv3qHIQ2pcUXaF67CQ4jh
7sOl6aAseCJEgkguxzkjtBULzwwJI2yaPhZdKyQ6Ua+Twsab8uD8truBDdOEPCXz
LDaf4AHk7X9VWvDfYhCUgotYXte6bn07Of11n+53vzdeHu2BCDIwo3Itec4pMCOl
UuxFZIWIq/9pxsHPnEizNjZy06J4pEXyMe/YQEh9N1C4Rp3XPTYoLABxCVltIaZj
uC0FqsFHhP2hcx0R9V40LJ3smWZqNDLPYf+iu2wwrFbK66RMOBrkkRl2CTzlU8a3
hYHSkFEhZQEvJ+n6uzYqCvj6vwgFg5cmMOzoOECBVT0KxJnADun2Cdh74E+DGW1b
9m61eQUr6QZq0So/Vc72Rn1qF7XmPtWNaQK77WzkxF6bzmIS3hsu1QW3bJBdgRb3
U6l33ZHkyGakDpAWDIvfdkyo3pCrzoha4hZU7tQXJ2+N6vVy4ZH9cFp0I61Wq1PT
c9ZexiocICVuOTE3MKSiET4a/3P4q1zDRvQgg+s8oQGDNHPKd6I7BaUidQhuinBy
KpYyY2CTJ5SwNPkyib+1FNp/o2h6HZeDVmp90mneWpgAVTI6fFE7oSOT9pBwRkUJ
3c3s28O24aSY3VYv8dPCCdbkcmS1AgctzqTQA04bmRrN0a+JcC2S+JBpind2BuND
gb5GTeoIKo3J2/7r53Lz0GCh8dxSLyCzuNFOo7VjHJQHB84th0vVZDD+h6KrUQE4
acLqXDFOVJ068NJcHfUgEqW1OlQtkNokBvyLtDG+NbXckSMP5JDc74Hg7dAKjUjO
jTtvBNVUm3ZApUukjI1sHjyfpaRR2fG1xfp3L2VE1m2F6BRnIy8PPdzaV3XXxa5R
UcWx/sx9IACQACFKB5mn3uwQF3p928jGDQkrnE564XkaOnIQpzZklhy4xbySEwXJ
jlh8nMOAAEjv60RuqVzUuRFVGwH5rzDpzo83fH+cPTSbEND4iD7m2lTD5FNz/F6V
zsrDU1cGvqzYvVHzNd98Qb7b1i/z8eDvKJbhLu7rjFfEydHEBF1beX7eXbkv+6az
7TkZRoYmsT01Sfk3YediJKyKlk7U7e066NTVtlC1yH4dUcDQfyvJO2ICTrkEBalo
BRmNwFty5g6JZFRDvOa+o7jlQw8zqJTigKaHo9BpuwbPuV6Npt40BZt2ZbhKh/iQ
sQ6mVy2lHfcAjQmEBTEUeKgH+3b/c/tfbgVrrAfkMep0BPU9ivyn9+wIuOKxEIjI
VU1xHs6+/0zXSjvYdFOz2HpTbfELDhnep1DjZEiv+Prkl7JdvNInuVepi4BkCuYY
D3DgF7HNJ9EREmBt/k7YI7ilQ/0TpP8CEE1jGpMbsMI7U+kAMLp7ckW22PjfhvF2
/H42xjR7ByavV4pe3V7ULX0C86u6uP0JEfJLE5JXFOU2VYcVc3G7wKskyd8vqJZK
gFaEyfBfXYii3vDZj2Ox0Q==
`protect END_PROTECTED
