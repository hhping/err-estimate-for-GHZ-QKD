`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u4Mdv3whzoKFqXeoe/uB0a8nWBP4U5afXR0HHFTe9H7l/gnf0ZuA1QWkCIJs77yr
ES1VwfaZRxg7/2SV6KVxzGHfCWaj+ktNzMiwVAdZ0A/AmHx5dtLMQb3WC3djyzQ5
DHgHud0T6Yn4sKvw5yjKnwZkW1AvzhHji5KR4MjHdMZ+nv/nuNsSPk/a+KLz+u8c
7RVITqM7feCiNm7eK9J8rSP+WSD+vZ6O+p0z/v9GLHzGacNMYdBrJhuiMNuLagVn
zTtGfmUoAs1WOEkaDYtFC9DRewWFmEfcwcB3GX0B0SKx0RMSGcGTGiWYyHk4wvFX
W09IxdoTLkt7d3qOjimfEjeBd9DZPiBu0nDgpIbiyRoYp/9ddBn+1PM8xoXuSoP2
JfIamasJ5HIo6Rcfdp4PocdWPmWk0pUUTx7VZGsvi7JZu83N2B4CSnlv6LX9cHT3
Q5tRe4Eh6CL5GzSJ6WhAMA12mCDj5vtDGFdq7z4CqSjTOlPXhpuHDDvdLyxEeYWu
OMFgsQNFNT+CNnd44L9pK8+Qyzubr2LYi2dCYJTI4l33ExIjpGe39m+5vFOZuwcY
9LLZw1mMG4clsQjtBgQn/eAXmWahWvQzmHs7RzgPSQEWIKKpDR4IhXJo5aPqCzrQ
VvaS678LE6ooV7mU0AvA1T4uGNM3Ziq/tCQYo+Xo2oC+yobuaq0rMl8fyILYmQoM
iSvHf1osq9yd3kSKjMhTZvQc9ja2hqJ2ZRSFdCmjpxH0cuMinZ93si/Y+OKzZtSe
rAiiAlCwR0yiJVEaXIKRepTewWaXmQ7QFrzelTh9N2MGrkDdw1Xg0H5Gi7cCRjOx
eVCIxMRTQ1GMrcA0+KmoKZJBvq+EzzqfUCPL1To1A0Mh09wQZmZoTVFGSSGJJMR+
BhvyV65XiNjUMK7bzulUtcm5GrgD+yNMThcJs7cbop4qbLO5gXHDy25EVPJnfAhq
kOp3sNe5YUAeC83dKzO02gzm+HrHWTCt+W6cdn1b9T0cDgaLkmel4/lChP12yME4
s4rIhaok4TTEVJ+K3241w/IBMuf6RnlgkpWxcff23cB0pHiG35ZARR9VOkYCskAg
Dz/GrCduASyZP1bTsFQNQGjwXIQVT/t68kFDdZvKafMosPE2xSMYWNi0+Lp1GmSx
wsdQvwXhYdRYnzuwiDrnu5g/POccxC1ZhAB5nW0vC8o9c5Q7833aAr4j/dmmJ98P
k7lLQqe6r+++Y78ifDOM5MwNVPLcVyW4x9CjCjINDgAaIatPH5epdpB6AiGU4nHe
QzGQ1WjTDYIaam7Ddm+cezXmVlTCZeUtbgHlvJWvhUErFRyYz9YJcXxd/Cxr7opU
dk4fHa7/vwHpSA0kaqRkScQfxqdVDklv3vWTc6pLHhIFGV9VyIagbKHCFHFV20dX
5NPsWX+QabwxJ8U3ZNqAD/2136/WQ1OA06QzSJ/P9U8XiD+jE/SaqRtWYBzy5nk+
4Y64LaFrI2vyOOh7SMZp05MFI1ANARs9g59dYMcgGP4/rejN7+roOIahhntXTsG6
hwec/cjVFMHfV4joOfVQkX/TCeSBgJ+1o+MpL/AgMv/yUtLiwPdHoYTNX90rGbLv
5AjvHDsJ91Md0hHRDtRbJ4bkAszmON8BPl7wV+Igv8yG2WEz3xPJ1AUCUp6pmM/f
9TUb9YD4/gveUv45mlCnNpjf8CA79Hw1+bIOs6K4UpV+OeUYyaEKJ2UZ32Jk2sws
BlaQAwbO3PQ+kuz6PRjQqsoc5qkIxq6r8R2XlebAeL/u6MufVQ/NHwQMzT/G2BEw
gnpXUtzPcEvOTMMawhgwes9/eR2quCO85Jbb8nXypZlqh86S/w+I2ekPSylhp94k
obx5nJybOrDWDL3gpQ6pDxlaSg8Xy4be1C1kitPLrIjzWokhI4kSjI7qUdGisDOp
ztf5lMy6tTNFIlBEGvcVwdP2tW83h5+RRCUa0jiWn77mxstUNG34RagdAIQV4FZY
flsmhqggDHJ3JSdcR+g4LMSEjhP2nkzL1o/vywuHT7DC2SRbIdTZiidzpvYujq1t
KemxJCL54pw8OS4rDzJZ34dGrFnkFVrmBeA+WvvTpgp0OTn3Lvl/dok5gYuij/RH
vg5jroWcQb57+1e6YexhPJ920+7ljOft8s3faeC4BGCyjaPPZQZZO9xtB/7gNKNr
qIaBdrAp9sz2qGKJvA8RiIb82MYAVoKjUkC5IP8cXkGjFeJ7wlfVP093EWpjdpJg
JoFQyJPALFKhVgEYQ9NTpepKnQLgDJazey0ZSgidGXtT/9LiPlOHW/SqCm6nyeeo
DNmKWTZZM33Vrkp03otMmMYNhsVnTO/sDz0WhJxzrt1XoUkfQG7XMdEDmgDIHZfv
g4iEFkVMoGryowNjCMdlP6e31KNQsb/vhpQrfSLyO1HsDWM5uXhBr+xrayempQeu
CDnc0Bh9IkPTaZ+ekMitYZ831UGzdi0EVSIrmCamP1nGJDIKbJI6blecBKI9+pO3
jche1VTUCKLEk03DqyR/qoXTLJt4dBYyJXwG1s1Eky/MWcoThCj7xM2xb7Ho5T+I
P5BEKORmrGcrytgS7V4ObzcfVNifF391+aWme/mT4OA3ZqZCgwHKL4PnKEbWuV0T
ObpMx4NWSkHbTVPQFSRoV+EX4UTxSR9DSvjYwsjteTDHADq4YO1ORg4cSGVHtNyH
d8xIOUZViPPtMLZqqrsaT+GUVszVW7VAkFubRw7UDSZ3n+qcO2cZmEK2m2dhcBXS
5PI5YqqvFKKwAMPNWGRrhq3LQ0M7VwHH0JoQdS71FUdqZFecZjm7ZMvCAPkpKtJa
N+avaJcfnO1rIAHjceo17COCdfNcOffGOJFadpVcRBTZDkS3TXYdTSRD7HFmMZl5
eLeiZnCohwpXwU/F2MZ6Ae3QMHlOT6xPqFu0ZyxXf5MuskQGjihXEkU6+yqreRUJ
ZIkDCV9Hb9rf0h5eR7/ldy0Oz4UuVG4f4TSqcBU1B0DMHKmZrABaszUQrAU6mKs2
q2yaogmo9ryW+FlbB+CkyOinDXQnO/ID0N2ESZCoku4jUSTuqcmIs6mUFN/oUz+l
CDKmpAWYG6BrvuI31V3pWcuTvbn33a3/XFHdUc1nNjH9d2Ox8WdoKgTWUjCj/A4X
lilI08iSK828aXRCJqTAVFZl6fJZBBLfiquVIGeH0OMSYvlQatSpD/Td5b7pGrEp
qgs9VsmFn1oX3KT4AU7QDhVfEzKd7d6KHv2Lt6iK7veOODVj9gC4w3Oqbftk+HcM
M4evkebH7hftr2axxhPNgnLT81HzpkCXT3B7MeP1OuoDXh9HVm3VrkAz66kYkEo5
SMtX0PgDXOLbRL8kH+9/r8v7t1WqtDa1REFOwOBNy+Byuxe/l2QVKVtV9va9lTE9
Hmh+qVU5aR3/x10kdAnBOn90EoDevd6ywERmXBNGpAeLpYbtyxuoW2gdNnoStuNk
llU9t8MOZ1XO96/3tFeKhlL3XWZ2kb/wWM4sB7O0BW6re84cSwK8aHXhb2p5NJrg
KbN7AIKTuGXbjjYRL+LSrIdCpQVAeDNVghaz5B3b3CGP1ngkP96EjqWzI+Auzcrn
QX/S6Rk884oSd0pjkg1DVpogreoVSdcvXOEIryqBsufiDemRUl/sMmd3hAfhzdcM
0YQEhnxpHanLGPcSSiadpgdhnK1E6Fv+nykss0gT79v8ul4CdLYvzriI6ICpXiyf
vI1l9Zy1Z4Iq6ATo3KzWjCwjrRWxxvwLM2QZUoMOhMCzUo8VOBLpGE0+Z2dQhI1J
KdXyL4e5ECsYsJAMg3f4fmNZkJoxfNrlbjZV+a0+lZTF7uQifcd/HCgdL3ZqVxpH
WikwTIqOAOsL6xKgB+FR+3gKfRnImn5ly8fIY4nBUsS4bYTxlX4tbFCPP72JaaTc
cZ0yVfq/LDvuVaLaaXnhABuGeFLUYs/L/e4NL52xJDHPjD2yqQEBJkUtPs//Omxm
jPuTJ8heOqe4VgkQAKNC2zc5QyPZfPLWwpQ3VWlllM2v4zgFEkufUkZGM2Y9EOra
2V7qRPTVu8lSUD4XjZxL2VREU7W6y52y6pCYRh5fCyvec0psCr9HxSi6+PWgqd7u
iI0DMH9JpRCbEZjpbZ+lwT3EkyElxA/yPr9T+0RS2yEw0ja4zZ3jqXPGJgj1smD3
k2m9V7i7WwyEJikuPXtuRnGd/OKqupqCS4I+OrR/oEHiuD143UQl095OTa0+iMAl
Vvh1+Al1H+83vTu53nF0vWy098ZdH3cmfLKLD741+k7+blF9FUrmBfp+i4L1ZHlu
odMWFJ148AN/MHkCSQWUTq0W/3uJ0tTSU7sTXdBQ+k3rd6hkmrB2YNvwC/rSYXJ7
PV1Iyh38xPqwyacBB+LIo/JbB9KH36OLq98PnzyY3Jg=
`protect END_PROTECTED
