`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kjg/pelRLZ4EBxOC/PgVn4N4dT4xysOMsnb1TKwfb4Zt7BqR/+hLf0xblUHUo3C0
8WgKZo5LOujK1K4wpHIfX9yHMOmldiG0uAwFTzVoH08ypz9eucQ5nVPfKSUMAgia
sne2zPZ3TfiM7Bl4svnopoRBvo9PsPyKzz+PVfntHOT/cSVqdn/PYT8szZCGxNrz
UYlaZkSgBPWbqjNNOLeWWnuRn9ljnKt5gBrzYWEEI2IB3ZRSezaUr45vLcWDrRwG
RpqlRral0fGqxLqaskJo8PgR5R0wWJPGmF46tbGy6WqImLK81cwL2avbCoE/2Y0X
kMk32pFRGOma/OfNTsGlQskFq+9+nVBMT/GJ+TNJnghDur6kAmigrWH7R/+GyIiE
GmOd9pRWiR7Bk/YJBa1KgMKceoTwM+wESvIIt/JkFXnzsmW0F2BBW7wcwPki5yh+
C1pQ4BXNnMyCOm+pnRgj3+jiG2ljnuGqag5rT2FgYps=
`protect END_PROTECTED
