`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvJhqY+U6Qi17oqEplYQ0kB8VgIQ/U8Foin7OJGnr9aDMiqtD9lPpuT8E4XF8xf9
SEl5TrN5RVJ5kt6Pug1dAo77g7GI0YJVcKwboIU7CP9Q4nBZqBKb7AiBiHui0L0v
jp5EsAXQIPCysvF3aivgvgkB+xVR5wVZmwQHzAYDkkiXtlAH+1O7Xy5TUVAcXMxp
sVVD3uP9VulKIzWiYVCVMk1rlXtuOWFDlYSRRQ40fMNxFoTD9Fe58WTDJ+GL6u5j
41ICdigZDFElAFvdh/ShfoAkJaI/lR7eS+Vuttbr2EfgSvYgc5zsBfsul2j4i3e5
FXIdrWp8lhzoyzfLYFTgGjbJtUoVieDwfTnXXUqd6HkpCUQ+zD9z5cEaXr7J3xF2
jcKyD+c/2K7+o8P6hcp40mSapWPGrsKPxP1VnCx2D6g4tSsBKBCXxlwpXHI3aWHi
sYtzJcHvwAFbDCQll9wiZDhebZvAs7t58mo0BDvOoydkT2sHlPoy/kQcGV96L4SK
vEcuEdOkVWlcxFCmxbbWGF5DGqQRmKSZvnxJoo9rFfgkHCnFfg6OF1qWE1gYn9RQ
gZSsZ+MUAMENvI4qdSeKYNz/UL84wgqLM2re44/ZbLjLTSsHwVWjv1rEvaM3iSci
5/oyhEazc7cxl0enJUkju/0dDCRpePqbymfjrmO+wp2Zrq8IQxpTdOdbT2GTweu2
hkLYH931OUVpXSSdZNl/if4PlPjPOG6RGUnWNCNE5UBrliNMM6ldN1RsV5OVZ7Cy
YiYm56AVxklmQrGsGKIJoA3PuIu91tOxdp1DjLR+PPv/PwUDKrpKnClLsPnvP2U/
QCIoMoWhM6X0gKTHr8PDy26bLokd39HB5rhw8H/Qh1C5JiTAB11PpTX/sxjEdbOx
`protect END_PROTECTED
