`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgsbOPFCv6fd7mI/XmM0hjf5bKjSSJSs1dlyFXD4aIrzrxHTLHHe8Av9l7pQ5zZB
1HvUjer9TPF2lq/OjHWouNBM+kXuJr4t3uSh9zcEln81bAJoyW5ybNy+0F5U3vXM
UYJba8lwVfPadSie5sEua3wgBR+lcSiHH1ORyp54TEcxQ81LNP/7Hz29ahcMcdEu
FsBk7t6prfxr+jNebWHZc+L3gdJ6e5LMTvA7+ecWN1sAQHR3I7GBgCks3BqyRRWf
zXoujVYkaYjAUZ4Z+CeVlF3UY327mopM7OTyz8RoVOUHx19mTvRPyxYDEEo/Vsec
9bJM8SNduVb8HDNzRafG/TKvrgcsSxxCujogPmC/fJ/J73VvE8hWkM8Y2E8QS208
I4kd9VKGGX/tri8n/w93tNu8yBIrmmx5kvgaDsbkLs2KvYE+wBL6a355N5gkN6pk
GleBZ1l1UsLNrB3v6v5X48WXL94W8CIWVtmG75YDGT00BEL9Fkz2XktYY+invvm8
+eHdJ0uFNKVacsslWmNUtjHtX6f2Y75mOPGFy42ErHixxjhSaxHGXqFs5ouEU1H5
/3XMfcVD/TtNl3B+AJytMgOJlUoaAyIKwKphOT+do+9riYLnFzmT2yF7lzYLBkrH
mxG7bW+eVN8W/3SfeKis2kfG2Tfhv/vGTcEhtZgrfFwJUdoqFBTWq5BvPEMmamgv
B39H7uldt+SLJBe2ABvVog==
`protect END_PROTECTED
