`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIUZ8AU1uX20Ot8haUm8VfH6RE94vCKgWN2j/HXXhBL2ggUpIpEKQ1lim/kyrOps
vg6+I4EdPVTdJUZ9ruFJt07MeBmJyOloS3Cpu9WnLq0zzUB0ryUgZKL2s6IkO/H5
ZWqL141SPLfsdC84S2Zws2vEaIAd2dnfQp1SAYJQQ014M9JycvRcYi+SuI8Ax0Q8
Nbz96qv2M5KLSHEha9CkWp4UHGmDFwJihKXneJnWtNleJAMZtKWXj8E+TB2mthbG
QNpEH4eUcUftSek3UEEBGzZokDJ+lS4CKFHNzCXz+diEE7jE4o2XnbXzt9oTXPAr
SyHZw14Jm7fQ9KrLji3XPUaCgGsL9LZGDhMySlb0SzVk/QXyB8BJNmp16+2g2oVr
qHbCFSPOis6j+pCbrLLuzqmzaF3GSb+dCI+ZacFbIMSSCvX/7p6ErV3ni177cnUZ
XICmibt9gsNJAdzJ/e9ZLvy0HDdTiquSnJudZ4bA/Hwx8X79u4sGXqg/bL2CdWw6
40syRHXwPqGQLhV0JS2sbynqq8jGHmxNL9zcQDxBaG89LFumWCv1DfDzjiXqUP2w
OADrXorb3vxFTaKPZM4fJJ5RTLtOq+d3728BucDbnaubcia+f0RCF1cz0bvlHTy/
AMzS5xmptCiJ+HBnAT3tev6ejh2CpkEiEFB8mAytdDPPRANt5oUAznced+HnglAe
1UIvpRXlFc9WaqzRnyRWVsOHqEDdMX+rn93nabDOD6S4xNwSvDI0TdZRTRjRnvWi
lk5Nz22ShmQ0hi/tQ0xRaDl8/H3vQ/+RPAc+ZhHoKG1G+2f7sOIxOW1+uZxOByE0
g522FvFQNX5xXr7yfbXCp+gbsY9tQAAZAZyHYh3oXjL1ZwhUaMXAKREWMm2hFfyR
qCSCH+7OYStDz2XU+Zx2cvPib+Fbtto/CfH97uXH+J++L14KEXDHYpqQS8glbhKY
CihG1hVNfWS/ssJ1w99CP1iasja3WAFPFSyOVnNVFT9Bj+L5cVX62CKRwSWhAUWD
I7Mx4ht6LRDmkCOnZPwhzP+ClcTQXYLDOUOzaRqjH/Ruq3xLem8bfQF3h1iJspYF
N8w//4W0fknrUHk47qf+o1qWaZjQ9RsiG3l85N3VWvFb5IcVHsJEPTTB+F0MYLVK
KspxNx8Wu/43jGONEXpYQ7ADHKWbtKWafN4E/0os2KeG3psqBfRaaUkYsBiQzOTD
lT9IXAd6ahy6REt7mKAYNyPcwykFbEK/7QixzuQDs+X5EoxxwL6UvfCE8l/IcvyH
twDB1HuCMWXEhQwDQDhtpx+sqTpn23DQbSSzXwZLz0eqw+nxWhNbvJBvAP8W3aYF
pHogxDQnuVauM5sM/L+LuqXp0hQ6rgm6NxXbeamoz1WsNs2aaBikKwAsPzDtXsK2
0ITQN//mMJslM2EwLgrslumgpJTiquhQw/xt/bLZ+ooSdwR+a5Kow7xQUQNYsyuq
0sxSRe5uwpeMQRXK2aEntsJbsmUVn5/GyyNRGeXMVIOpwbCFiIrXa5LqS/wDlZxL
cr/qONyc04EurDkrS5ESI0j/m9U6mN1IUYgEu5UpfrehNomdLz8Bvq8VpHfVhODx
7GwMrRIDLJviNayQZxJ6o4pC9S1q0ytOnqRG93y34kYY2cbMQSWKRTnqA08ejDF/
IKkDcA5frXmlvpNf2SvVEscNi1QixGFRACiWcGtk4C8tOSPntl/bPwrQ4RXzS5GM
gUGmuxpxg4zd2tCEd9N3iNPqz0yKcQL92krVDv5VXMz6rQ6XNIu5PuteWpF3iT0H
GpO9nie5NYUjfJZna/wWdsKuS3S1NxCGDhjgbpGuChWlq3HxqJew58CLUMglhzm9
cbfQrzwiTX/tetVQ4JqYVmP2e2rdYk2vVQ/it4v8gpjMDiC8DPFF8IyNEdC9oTgw
uDkCMwGlSr1+lIMvKL97cT5qgNRqQgURuiEGLm3f7aJJ28DPDVabh9Tb8/qA1G0l
hIKw29qBZhMVsBdbb5wqdnlhKvTcTcu80ZAzIYPISpyQjGInbLGZBuhpWVG0lcIH
/IIMvP6QN3+Gu4PEmKEle2kpxT6w8Ol3GfWitHUauHTwwA/lw8JvmcFPzWnr4G3o
GDiKjv+hkXcLcmVkKcLCe95jRlZUAFKeaDWWSmouU9q+dvtYH/yuCBORXCl0Ww6/
DiSP2QPeyvyxjDZq8XiEtPgk/VINtSPjuTvSlD0GMnF6ELwWex9FarTSEzyTyr/0
0zcvMBy45y5e+VixEzUNujHVJIroDWHWYNOeROrBqDPCuszxLVvnsuXJUKB8+Wa5
S1ibSWV1mLlBJ1VfWxW4tFRPef2O0BmbqTxAE/uyIglDeLSo01AGiCzhNDMy0WGe
Paj4F9+QWIyzfwRypOKpozSyMUf7vvi57BwBLyvhvFYO0YOvBUEjIl3S5ogIWvde
DCrjyvA+VWRBuhH02yJINDz74jJNAA86/U2mOIW6W/xYsVIjAUdZD+WIrYzh7Bcz
w+erXz7rh5bjoovs6ZkLgt+7brruL/zzakiGBR4IOVIXKDvFzJiFy0lCItOu2PR1
Agor20fAI7B0f9ppU60GNE5xJnacnIIsVFscD74VyCKDpU1q+m74Fo8Wl7LfoGE0
PfH2m05LwdUe8ONXBYqX62ALqdOFHea1B9oaCBzZNSRlQmsp4eC37ke1WQqMRj8d
Z0YYqSse9YDjU10hVng82efpPV10SRJqXCh3TpY6YSCKZH4rvZiH1kZZ7pc0QrJ+
ZsUXiN3IhhYHHd6hdSFRsDhR73FaC8nG0V+Rbsj7+9Sg5Jm4ZvfwwnySYguur0JT
xIZeDq9tQv9uwK697gKb/gD0C5KClfgT/Ebaud3j0H8NkSbhMwipoyWNsXXzrqtq
ioYQwR1Fi893D7e6R4zWNaH/fDom5HOggsWkTNINLrSMlF9Jt5MpyvJfXJernGQQ
MhZooDsgdJ+AzRwJ+yCdhnSt+6rU6r3ybIH3LpvSSJnrMyz/Z4fEHjFvrf2DhWED
9rq1Yx4kfWof/Fgvr3JcHAKX3+L4Oq6YlsVy/eSXBoLmI+BruwT37s5azKXSEpJ+
qdwZTtvy5RfB+55C6COTuP7Flyl1KyZoy2QI6UGczcc1hAejjdD4IRn+BIGJnJgG
RHaGY/tjGFBfwS1HUQ4ArKtgsnhqo/6EMTNllTwZDLPlbxo3SlnSGFJyY/colU+7
JQzkp36rR0p35dmPJN4u6hTiylG2yQeT8Hmq8/2sQqRsvpmfTDahLlb4nEiHYg1F
DargfwP4i8DKPmOF1eaTzjnkGki3JtcvPnemZfixU/VeDeSUgU9SOgXr1AHhqcbm
CT+KDptn+kKiqTumekxagozN941MChX9tC/RelqgoH6MPtfAHMg2eWkeNvyUcOEZ
H4nw7ms6jS8bwFoK27H3Gd8N+5OQATMBRSubumdL/4/MyKbQ1RmqxO+gIvybcs1y
H6S6sI6c83s0jbCTXoH8TlDhQY+y8tCCepJFz6HlJBGTjgJ4c/o4TBQvPGIvaKYj
zggagXfOQ2AiqtdZPsuy+MpxbvEUuk9f54LZy5MhSEUzQEHrGQWgykwKzAkWcgHs
F+HH+xa7OUsPOcAOTDkKP4mJV6mES37aBq0WMlo91vh8lpAQY/7zARwh3aeFEmhF
Avun5TwUVzyYz4inntxHHE8pPvipXxxr2x8QkgfpGQxxdhwEmBZa6WjAVBz6slhr
Z7x/rRWLXFN0Put0IIXyd1+lUNrzgtaeyuLkn93C3K9L8WTq76pHd6ce3OqlLEjo
yMfrxk9Uiu9athzSKLmcoySR8xN8i7uF9Q/EnOlzFA/s515bMC6F16kZADVrvcbp
wFw+ozWe4A/Kd/eBFaccTwLhjNtMlxxFM/DK+h9+Bw6pLeH/UstlLxG9HVGrE/kq
VuhEClAYricqgumakXfkJ1YHO2r5d07d6hWBLe6cXsJOsel1wCdCSI9d1ew40sW9
4yEXx9FldhkfRm7FAB9llYYqKHbrQjbYm2szNyt8antlOJsBRpwnQ1J844f2KbBw
iVb4/bpIeqBofODMkf0E2xc944qD3jABzTATravULe0C2ijVnN8Dgf4HLspBqQEA
VXBslqoyAOW8T5+CexUqevsSOAbpBqsisdO+18vdPfh2pFIKOWRjhjrKizpcjkM1
y9QvUsMsrpIGepRIc9EhABeVJ9SBSuWIYGaTZib+Ol2N++pfF6E0t6V5vYSHTJsG
lx0J11qp02YVko7vdqQYIaHtIK3xD5qGw71vlom8bcGZ+6MRhw4fyB1bpmnE1VsH
zkNeBCqtkJmqOUGAC3GVvP/5/5x6jPZ+HNyNQbIGFDLOILl0y+bM8/8nn7j789PN
qlJrCEBzi0Yznnt0xGR4CVgRbPc4PadHACsPTnNY8X/QsvNQ6IqVBiNH8sos5Rke
ZP2X/x8xd5UByOyODi7DVANMPZZUjYi0GWNM8hWRY6qTFAEsC9EwedY9lp5+awHV
gL1CvO9Aybpig5eg+JXb7pUFEA+FZAdOxIxA8Ml9zan5YXAoCWx41RWQ8XvjtpyL
0iyHYJjZIUjYoY0RlHMPlvvYQiNWFskznJAtqq2O/e3vI0H+w0Ubo3mY0/x4cHKZ
UGj54AII8fPuPxiUZUkU8kQb/PJxbA9wLemfjY6dVZodjJ7W9Bbh7o+3knmKSjJI
2Mf7GX+bIVnb922jiQeTZEDUYt9aJRUxH6yjb2Qypuw+h4j0dZspNZtw/1NeB5bP
EAFVrE406ev2o/rGrThOtLvSxJDQfiVWPTX1UjyhKeUGy7RY3Pa+GcN2sRLLObaD
j1M/evOlAzp8O3n1aO9LvcNklDfeqhqC8yS34fVDPqDt6mzBR+d8eXYRCVs8RwLL
i0/bkytmaObMnFyoG7TNZTzSD/5zlclugGS/GsTfaQFHQ02CpMVdUGo22NO0dniP
riqLm56Qua8093UYosvEsdFlBIfDnv93lsivg37uODKih/YFxyyKfnt63yH5N/h9
TRfFRzQIHMfHkbZn6alVUqzdE3SWo3b9GnTNBNvo/hSMnrDDVewCWnNMdHUeZrnV
Pt+RrYVXAVdAFJBYSCqFCN0j1IHsjxeAdZi3a8jKUlQQqBTEEcYO/9ku2wfP9t8o
IjlBKjMprJ1gdOEe8m0es9O891mRT88lM5+nl/WxT4U=
`protect END_PROTECTED
