`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/W0tXYCTIAaqlxD9B7Q9oe981btg0teacdqI41JmHl9Ta0FsF9ymIH76hw2mP65
u3OkNn1eEY9xgOs6Cl1/pQE7xEQK7m0EuSPxcPD0nUDwq95CYhBHNS+Y+pcI2nvp
X2uLwNRe0YvWL7P3DeExZQg7+VqQ5ifrHDlkCeQLvcRWCDY7hw/FVh/NBx+4rOH8
60fC4d9U9T/peoRyEHVh+Po4rwPIM06XbARhGgcvc4VpNEdHsdX4EWo88OlEa0np
9RYoxSqgp28aUZYnmrGADAS4pD/BkNTCF3ivpfGbuR08f/F9bS72oLWMQ9Mx1cJ1
YVEoJZIA2+yKU939zs9NNELWKOrkipRWLjgGmS6xU6J+fODHMsR8Kn/RxYyzGKGm
99b8ekWjGNdBgbpAc75Z3jo4nqi5zacdx1FOi3wdXlcXuEmwuRXrg++nY89xJFDX
l4QzH33hMrU+hGWeCu4IJgNDTbgwudWHL+y5nE8ckH493nIMJvcGNHDMulcHY3Va
ti0cjWWbuEs32mKJ+g55/lysotk7YUJoMgxnccxbt1ZqR0R0xlNmnu5QasKgvJwA
bAeZbVdOyqCHy4LnShvqTT3t0gd0uR8VEBZl6M8O+osIeuX31DVh87aq/wEnYNG/
VVUEnIooH6VXwuV2Zp/NktvrhzY8yWPYM2uQDJv+YGDcoXDE+fJ+NkxoK6t/bsfF
6IzX2DoL3mDXT1lHY0B6uPBAKc3uQX9gYiCEhVhwqiHtTNcYSuSiVGkYgNu6RmnM
uTzIUZMp560ZHATQZ2gWU9gd4tGUefd1WRoJ/nTO/O0zLCwWR4M9EI+gfU4MeI0n
2URUTSY272Ftu5bFZQBAWPp09rsJy/pwJAu/TjQ3mflN1NXiuVaP98jO1CaWIUq+
Wmt79RftGieJrd1adMK2AMdV2m9z4xIuOrJkYQMC4V6M1T4u2pQ+bZHDqDWFYdcD
leXlCTCI5uNknCKmYlkx8esXaKgKoNo1xsSeTpCgeoVd+LwqY9p9L8pEbM6argR0
GoRHdC9kt0GbXByZivMaY28ZtBDbbfsFAcKOfcsoF/WzRSERGhnXGL1yg+keK+F3
Cgf0MltqpZWQzpkJuWlonLlM8gM81CmcaHyMfjcIPB4trOOETM77hvG4KOKViQVR
ItUqPwWg1+jRw3WNXhqPaJANmyOu70WFLexgm2IGUTW0/nT7QJdVS1ulk/Q/4pcs
gVF2JAutVv4AcpULksTG+K0t9uPZrCMyABP6qko53zJzWbuZrRFw2sYKdqXWiZvb
075/XF0rgx/4E8RsiazL18F50P0I2F3aqupv6CGCOrQ=
`protect END_PROTECTED
