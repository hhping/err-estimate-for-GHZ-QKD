`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e450SuVUFJ57IduApKILIynXYsEvYf80YzDeqpCoQ5YVZTJmwhdJaRKXItIcoSUT
epiPUf8goThPGKsEpKkmVgS841c/+Jq9NO7zdUJTXsKX2DlZwLXsH87YbUpwZ8oI
KKzRk96zBsZDg5BXzFt5O1e46uKgORMBGIrJCv+4quMDWNEouwQSC2bPsKfCt34o
TVfiW540UGUzpGNxupZDC4H6sv1Vu9o8Zm81DEizoJr6n++Vey+fXTNie3oqKult
qgjwwM7ivS6eLNCVLtd4uSkVtMQSU1VihVz8qLZjQQPHEgV+WTbmQhZ4AZrSKnR3
cLKdyc+VgDafeSHkPZUB0FGcpsh+YGIfIEY5262Ay0iT/IBqmlltA+0JTL18y8mz
oQqBkVLPTXFd5PPXyHb7yh1xcN01GSnlOQgQE4HpImuv38PzUnTxZuQ+s/TzhgZk
3SUoY/nmfJxzD3cl9B2L4TEK1UOuZWhX6n0shSOvZ3i+ByriJlshaxD15xpmKzMD
PMHyJ2TrF0Ym9ri3TMgpBU64rHXt3KRUMNYFYYFn9W4209Bow4RNZHKgTxQ63TeY
Ugw8kiz4pOpfeatFi0p7PqNQUGswXsCmfIuSVUiKN8xze/NKRkNyBXfOegmd6M64
RtbpElbp7c4WstQo3k+jil2wRJnlLe3odDHALFUR1oS451MUxT7L+nM0U5U3+yZA
0iO7zrIybf1SN+ldTwuxP9gyUNgiAdu3OhKVg6X+B9p2xe/JLtfIYPoEG1zcmboT
rt+K9l7JjRoRhM2lkh2gDB9W0O9lh63G2bpNxoEpOCqdQE+QQkFdCbZGwPy9mw4a
DkOwJfkP9XgA3nqdiH7dyPIVqrfWzDjJc/ZM1fdHWWpK0xUYWNB+Q4dk7JfLVJNk
xGDm3nFSSYcY+GIUflFrUm/Dr1smK41FirSeQqbGbGt1lS5QROARZ+HlulHd9pWJ
/ykFL0KHKw3TmtgLnKmLfg==
`protect END_PROTECTED
