`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owg5+n5E8kBiOPtdL7iqWNhc/9b1m9bOds1G2cguiZZXq+8ywDzEo22xiZ6lJHvf
zr0kBA1wJGtU2KZJxQeOmOhiAzC4hUdkZqsSS7Y2lbz1f5D8C2FB0no82kSVkezL
7zpX0aBLZWMiy97vvROpXXmI35toNer0HbUWXfGgBaJvdh1vMGm/gfYY55DCSRoS
/giyVHDl3R53o6h+rNts314akXpBfETbWzY9KngD7+NJhLkw+sswhVvbnhalXpAE
mIj6fBs0RDLYLmRMtkMdFPpUhNZitqINN2CHiZdQCRPk1K6ehhsN/FO8EZIuhF0w
H35hw7XgXDrymJT9o058xhYw0vrkcxBZAgbhWeEl+3PMwU1dBgdpLdUkJu6cbh/b
Z1XlbV5gzEVi5Sxl2UJynQitbhe6LhqzxBF5bR8xIapJ/Q9aoHohzW4g2v/mb50w
ICyc2Ai9YnAzKlUZss5Hbs0ekHZ1NcYwfZJeABnnGkycOOAMHlRg523Ol6tbP8rF
8tTh7zUnRuB3sjDZYlPKBYtGzUgL++HtaI0WfYQFro3NOqVz32eJWwAqbdTP8aw9
YudXcYRRIcguXUfsfTV1IcFso8cpvAqdz6gNIUZ59nFIlSkfnn/N9XOevd6Rpg7O
ou10lJdWygxb4B85fKuYqmcA3jqUmgTS1YxLcVsSMhTMZVIv+lcq6A7l7oVjbDvB
ZgY+Jp1sIAUZyJsI6RHBYhZNjcwjXOjYFgtPbd0l87Ub4jL16YEeacy3jlCi9+l5
hSVuzOoQIo+Am97HceiwLam1As3K/NWoCOq5RU2n6qUdF3T0au5V26FlY5Ns5bDA
jjhjAKgTTdfRHNm0Ukn9cHe3GgGrxTyHQlu6P8B7o5sTYkH2oOQw3ZQAgn/CDd9k
VNEnarNJNJBBFeB3Ssubwr9LhM+cK9pg+JpEqZzIfT2O40osVDWJC5mBqUp+yazC
c77NBUIRM6vMk57a2LkSE/X4rfhCEQCphc75AYJ7oHrv4UJD71iMFTz9sPfZj+Ju
0jW+ieTBhd9+l09jEPZYRsALTSvyacqnntQ1PBKjYxKRYfADo9tyO9UA7wVQKJAD
I1Zo36GhkZNnBTR3jz/FW+PMIGECVnEQEvaz+0LM8G+1HOpIPSbOUI7eLfuRpGl+
zMP1r6jC+PdUsvYaKFUORDiPfZPYG7lvevo1bOtcpgmQSOdhLqkGFTIHWLOabE8v
BTK0SOLkfOsHHNhVQyZwhShFpPvLRyxK87+HY0cXUTPlR70pHp+mHSDnIjm5rniz
8DB3F+4xoatSzYhFbIHbJyaxm3G3moUJd/VOv5pSIEhk5R6ecJxpCfply46UfuQP
rgO4oDY5uVvTWpBFXFwxrjKhpD+Vw1wxVb7pwNH86b0XeAg4c3njec+UQICXr2Or
tG9sOLj9OyWGYPjyuwaakPcgAYTsXPsVOf3EFJeaUZBlpOP7gwiPMMkqht+dNpuS
GmlBt6u1w+xiLW1PYW1uq6DusGn83b7pCpdFy1rHeYT11s7JkXzWsFuyhpCxNgsf
fgSj457Fh0iURl0hsFWn2nOtLeMVQpTFHsmdXb8Rjvd2KKsyYg4BLYy4yM9zfrcz
WTTOIoBv+T2F9Rxfk5yUmaTtYgf7XrCzEO0x0YBNVtSxW38HOyYRqc9y1r5EYlal
`protect END_PROTECTED
