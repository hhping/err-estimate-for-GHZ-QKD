`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZECXLzj7kGdYtJdl9paJaUFZnO3lC5PstUJTxZxXPVqEiNf5UZAK4oSCC9dqWSBP
HeIKOvcoV4MtKNKXBJE5v1xxd3i8v70NPQ/U3m4JnT93O6tJQz7Er+o6miJpq+tS
Ch2YvY65cE0gjlTYAzzgsDIwzc3G2Ih9soX95+8F4PM/B2QwnuST3bun4SB0qx2k
aJvzX/kpD+pFDT6ZqvGsu8Avgb9hi8HXejz3JsG3hfWe3Un3KfRpfIjiZzyP0sBy
t80fXOgNYYFMYweheQO3IJYoYrhS8U3ftCbahdMVpzay8RRIDDZwCzIX9heaXrL9
t8w7zInY3kBgZb0iYxrcB5y/5RUWBCk8lALA2o2w8J62uVn1LxI1tcvroMfOEtgb
jjY/QSxHwb2wQQ22GxqBYfR1wecbJPRrAfUo1rEjC1+0PmCzrGB58TikrFZ/+vbm
4QABbMwQf/Zl3wiaU72DS6obBa2JndX+9hykgpGVysWkfSu/1/v5D0Nt3P7+KX4m
RhSvb5NOCjb84hCSHuDqpPosXcS0wm4SoU5G71mfBpD/e3nPV8UTXy3bEeUg2/Pz
/iiEYwuSE5bg5KrMhny/5QAGNfaEcD3KULljgF88UYp0jgJGpYPHv+DmJnT0T4yo
6bFSTV7HpmXFJRRVyOkWvmbXJI0TO/9cEH4Nk55OsSYG7tWSvPaQKbS/KojzqL6S
SSMckrstIU4G+XYDZJsj074am13LpYGFjlZPUQ76UfapfU4TPkPznDV1Qzhb6dtY
5Htc621a2KASSPThH/T4GLLa6SBmrISjQ7iUB9ySebcVri7atE0mS664hNXHJu8D
sr4bHChKvYAimGS+EaiuCcfUCcHdWtLj5iArgo4+O4+MzuTiwaG2/JzeHctDS1PM
7ens/S7ZiS/+kKHB282l7DSSD+DXIC5FyHgaiyr0Xc6OiJBiySYfHC6nljd4b9eq
/DZ8/j5I0A/5cqXiNcbAumZnH1KQkvrWYFJGjLiBtTydmVAOtdWm403rXBRNraF7
dIZAbkDJSxSINrqX/Ki45qIKTawm7hhIXoRXUrXD1iBZygwbVVRPqeJJf7evpVgm
qxvKK8jkt8D8ZDH+t97CoclFalwdphctlxBLMVlmdy617Oa3Fl3ffFaXMTsRJufT
03kUF/mXbZ0nbBOlfrB13S5GRXjwoFgg5cfgDC60WMASSi1rikswMREe2B7wDm5b
4C4fBuWlg0liXdPQS31BW5uPk2DYJchQJRbSASb/axSR20nXyTjb62m7ZGtkqYOH
/YbBaOPYvAnywIUyRnYRNlRCdv2YorTdH6bdEpqIH3uxRwglZ14dlowfOSF+1C7F
kiZ3LkQ6n/XY/+/OOK8jpeyike+1KO0Nk7GvM/KsujPY3DZ9NPbzAWaxCmtpRluj
rvg9+WaV1qJ9FJgJhxbACt9SqaWHJB5wehWQhD7L8Y6Y76M2jTs8/V9ls+ObXD1n
iS7z8bN/FBraS9TuBSqQshTIhs7vox4LW9NPOhDRPPNd+ivE/1+8JwllY+jbdKR6
QnmsnhyS+/CDK7jCsLi8zVg7HlK5U3gg1tmOkqWn6IHmsLHMDCm7b3SpiWRQuX/q
IZ7QYGibdhNwdwG2yw1vHPgvDCaOZC6ivDGXtOcgOk7yzz27+BgymCwyTKzeewGT
opiN5f4SjEwZv73/zsqCXZQwuzSajwNv7r7wWZMnKDWnLBITFv3MFc+9K2u/uCoJ
IXYtI74MlPeCjOztpVm8AueDTvbgBOZoceVSCYnT4mpekmwy/m/pxajKPhe/yENC
+3MbAWET8wfBp8YQMTEwgylURyak5rIuEMdniQkQxv4=
`protect END_PROTECTED
