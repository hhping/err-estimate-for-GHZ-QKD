`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M85a0m77b1EQQTMUjEknD3kBw1OeOBwWdlxYLWfK5xc0j/DkmYN8cYeBSOtlcPvK
JIN/S4htp49hwt0H83j0nXM9eVnX55AYALzdHCv4Tp8ZXRpjlq3L5I4k5dFLCntD
phi2uaoznnwPbMUphXUbPZRdgPOTKGk4ew8QdIpM1mIrK6UhWgPSwbbNLwmb8QHX
0rrQ7fVQD4zQP+JmkTK5oHEWBsRbUaHy1of6d8s62wg=
`protect END_PROTECTED
