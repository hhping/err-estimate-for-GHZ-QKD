`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sghn/FxxN0B7ghRfzlw4I3/3xILBKykzy5DtUZbQpsymVyZ9TXNIzAabWXCt7vq+
V7QD6p7Rnm3Z4INSmsR0lPuFjpfUhTLhE8ysdPYgTo+Grn4hopd63qNq2TbnCz5c
mLjfEPAd3FoLRvYCiNUT7Xqf77Y12IzYOdPQ8srdd84P09fTc9Lan52BiiavYC5o
f4m45bYg3VAoJYppcy6EVn+n1MUoNRf0aR8dTNFXNMJCE8FlyvJH7rswgmi1FqY7
QCP+wIvqb7C681jtTk4/zjmkWlCCEGbEpURbpryDaouocdvuYkmO+rR1bFKzO6FC
tV/5yAMp6FbINZcIzq9oHiDCfcWKaTeQJTroRtih+TJ1+YTgmliFdUTvQsPqOcnz
txKW1tl3V22CPhfhxalF3tT+UkXj/u2/ppEq9nH8Ee0jpUlkDjw/gtaVwPuucQRg
JpH1QAC3T5hTW+Pmb+BvgzyjrYGDHTeO7pSKWonVIWQ3g65swOqN6YCSRWZfblQW
wmrVXgqUwjeGx4J7ocPt66/ALmAqkahol8hWtTZkm+eiQ1xq1QKbcaYz63eDxJOi
hfhoDqkOITTDOKACqTBdPYwVzUUBawTP5W8Y2IGh0Gw6yIPi1PeZCVJvKl5kWqVv
jDI83QH+3TwEWg43pMRkTrYOdVW8tnoiDNmrncuaer/1ErFqjf6FWnjYiY6ZJozS
EvpO23ykQFozTktYjdtnIXrU9Dm8kYKdgX/tZjE7A4KwVscwv9hWerZ+k/diup4y
w4bD0ybobHZa5PkrYfl74mZS0bsI+sFnnl/L83YJL+H3jYuKUftMOXMkO3tzx4lm
hGDEz+wDU1NF3UiE6JJ59ahfILsIHMAxIdULQ6tbpl3hp+Z3+8zM37ZGtf8CDOjO
`protect END_PROTECTED
