`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VWvBCOTt7awzlcv+KtiOTrphJ4MQPR/aLL5xW8c3WR0aSzaFQy/rZQOrUd9sMQw
jW8fZTKhoeYbszyAR1qdXy1KWmMFs2pVWU7Y8prUtnNWPlN/++S9q3/lPzwQRLFB
J0GjE2eY6a9zywEm+YFbcY+Fkl3Xzbqv2qTh/MQkSZJG1lfIyRRGTI1OMhURZytb
4muWX35a3fhj96nGuv5Unw9YHIBlEJ46+Sa+Fys+o0vPsWsJu1sZDNnciwq+YTgc
c238Xc0RnTnLmLdgSzFNDFiiWqL1sW2gFNiToQi02BzdPkwvGihu5EH7nPocMs2j
qPFUvMSD+Vu/fHx2Patn/FlFyvLxcOwT825uYbLN21pRgyVjlpeMWZsZTU5ZgcHQ
862KVgES1cFM10mPH1h+C+9pWog06ybvm1VwFy5hD2DA6Gb2+B6mwDVX5JzC0aGA
ErLgP/nCPJjc+V/mlkIBLtNOUtyl4BUFfpWq0M8Rr0hEDwMbG17yHunfu4QT7j8F
cOq0KMGSbA/+2iNV46zVfwGcLEDYYAhUSdZ1ruSLXV/81ezv+0+PAktRfVbj39Bl
hKQEnOnH1J3ipsxQXOatNO3PRLib4k4sBPyrOxdt2B3EBEKqHMZ5qT5uKOCBqssh
sNuUWvItWGQ/JQBzbvDqfyCP1BOvl+5cnPBZurRRnUo8XSma9LHLjvwWN6zhhqcu
eaNdRvbB1uQT9F4m6Y3NW4ii72lWI/4fL13x71mbcQ79mk0KfNjsOIjvZJGGKE5h
YyrXjUOpZeGN/rHX8h7ewFFqjx5bas6A0h9j7kxCUgVMgHff720OLh+YOyTP7+Z9
Ul5g2JX4X4FTsdGGyApXlPn0fCuYWR/VYBuQgWviptl5NaGYZ9JG/4wRAxnvth1I
WK9TkV/POChhwzYY5Og6k+XyowlUyun7fYphY8fSDDN2KLduL3LVNvPbFvrbqGKP
`protect END_PROTECTED
