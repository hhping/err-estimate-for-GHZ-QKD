`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tS6QnYogzwDVorhPx79z3b32t2A/nedLvCOnVt5onhyy9a2a2UH0TRGemtaKx5aD
OMaQ2NacqOJejuEGVWFuhOq/NbRQ87a5uxJ4vshnmb41cv7ubmTyu9ww/R0JVsfh
vAf58NH10GZQsQ52fJ0V/wlH7R4yoCyEoK5yhjmxa8Dwof+2YKbaOpOLZQDRG4n2
a0wgb1TylIH0X8PGDBMz5lV4n1fxMlXuT6mFeA0NouvR+VO3tC5hdl4OlqYNuGxx
TibOH9Ocm33QaAo0GMbR6dBUih5qo0yJdMHJ7weGLbDRZ7Uif14dj7zBDrXXVLaG
aqlwcpzpMeDK0FfYWo5mWkjFhqhNP7WAHfCjzN6VoVwusxcQ9VHhnP6iXULFfdLA
lwYHeO5dtU2eJAByASYEJITiu9+SQkLxJYBal8rJmp9fza0WQPGKROgb2G8DuS4y
FUTENeok5x0d4xDsf9vk7qtsMSTnEs75tuC9hEUif8+t2/mRMHMDkodLlJn6UFCR
A3Hz0cJx0DgghW2y0/qY7SPvSLiA9HtZuuk/RRgy7n6s18ZKKQPTv1fiX4EVuVND
6lVVj7uTTEZsKYQ/bj7aXeRtIPcWoxR5lTU4qjfLirdqbT437bTL9RcaOQ4LpJyH
vKV9u3/OHuun6vihEnpNh21EFMiPh/AjY2kU3/cocciwRjElNN/4x8efMaQXetrQ
msIYdspH8Vfw/f5y3D0kF4xg2SuXuLyXLtnSSJ9ifbpumhZjrTEcXeSkUmuEzgVP
M38y792RSHdua6wbe3BOJbl6mRtNyAhGSp/dpPtxXs2PpY1xu61ILxMXzECsvtsB
ensneWdMNyZuT4q7+xL8pwWAzblWuNf5FltCfGhyeo0ET3Zth6vrAg7wsLxw8XC9
x2p3mGor3KgGXIP1agC4wUv/BvOkdxNsgQEgY8CEArjBN7Rk8soelAhezGMgc0wN
AOZaybAEHtGjx6Whkf9Uh4PnJxApo33rNe2qqoWKUw6nV0CgxoKvmH+IxeVCiSUI
T3+MhPh0BONfgLxJrUtsmJG9bIcgtOW02jibPCPVvGWA7bk5yURfrCZ1Lz4d9pTh
yktCzNuV56i3vRh4+ctjOGUMXbEzWYHeIxfopfCxAplmEnQveeP+OXbpwiH1C6M8
ADD+bVA0RYzhF9ownGMJbgQNe2o3euB7cRwp5rW5T9F6sU2ECXfIigji2OErg6MT
vyaygkunXg5EIIaF/iXjlVOdqUopNsVB9UJGrFXtcCFOqoHER/GdzaLmo8l73eE5
SU4ANTSewigtxmtTE2dOW6Z9GF/6qt6Oa+VD2UafBco3w+CEs7JH2IkXmSlOFdpU
AWMIuauYil7YOIdkssEbmHW4s+2gK2wdBYU0VLxlz8GxmINPACXMQ4inxu2Fpe72
85R3mgGTO0wvPeNEnObbgsOBCsjQLJsSLF/Koz1ePjTmyt76zI4/oUO2raJMXTfk
eNiHj0mGjhyP/zCEp2qedObDagbTcu5jd0bs5OoKRBF2gIiJ87uHugJnj6jHqlGY
aV333e2hc3jmsMwrsDtABzUpzv2vOqJjEpvBITrqeW1O0AQaX7hHlAQaoyJgJa26
iSufS5pFBogN53S0icn+tU1ROhd0wndz/Gj9Ve69aQknWc4rb9gfSoGRnw5kLD6v
NJ/NWtH7NyGiWDeFg7W5QCDBLwApr96sixDBC3wIH/nkvH0oSTe/OzBeTslKLyzy
H1kJUTXYw3oWcxGlTfZTT/QJiokIbq85jDddYEu24CiJqzcgmZDqhGby6ic/3ByI
peOWqbzh4mGi/x42QsuidaLNeXr4M6Acu7wTGK/1nRQ16YbQLJQyi0Ip0nB0M24W
/av73cpUgfPI0MDr9jVPTHZk6gGZ1Z1vs7FeCgbFNMqjmky2Q5hNLNPoT5dnHnfd
Mfn8VULBjKUOw3htA32Lq0BgNMUc6nh9DdUyNCzHwDAgEx1lRVnL+rMMmFbwx1Vu
vv2Wr2KFmwhf2VV/BYmZLLZaGErGfGBfbUwfH/6SW/0bk5wH522XCF2fRfIMfMyU
KW9Pk06yvF2+4XWPSUcOOqnpW+T2fF0OaRp1lYmGqXt+alpyNlhIZKrp9nteqdOk
0zNkdgk61gb/UG6zEX4IFbsBQ0aG90U5mZxFsL50Z1Ostd/0JGbN6BBhFX2zBWB/
/d9aceyQR/zqag9Ky7MQ21WKVTM0lZC3UFAMrcbiL14g3sGCkKpLJGEVSvu/xtK5
lzoQHsyvhVZ1omHni3SFYbw5Lid4Hnh0goal+VBRSaRD0MGA5YVe9Q939KzNRLA0
vFCbZBrEB0/OaHgb318EpMKtonfc1+4oxElTq6eeXmKjj+xKrPgIp8eWpRR96PFv
5B1EcVeA1GR/2SsZDC71KAjV0sskZCtMhag/r6u6lcovjCOEcAW40GWbl8obJT6+
mEQ9k7ja9NkSQCYVu5bLSVCADFAu7lf4ibu9KzcbxKU10aTPZOHVwXztOWcfrW9i
`protect END_PROTECTED
