`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCe8594cq7boiYWEkToXSbzGUq4VokI1g/v+OuIoiGHjHabruu0BRe9NLWoUrgkL
WpWwDLy9IDiKEMW2Na5NIQCa1W90pk9Hnzu0TMafOudb5DK6kRBU+DmNJsbNl0zP
aVckZVpZ2G0X6x7IA+4vmGC6A9IrVx1LZVe+K+pk9TDVDKNEpyow013Ti9CSbgJS
fNrX1QmQXDuspoIXS6vvniU4NmATqrtDJaPfueBdQjd9UwJbNVU+s1PVCy8T+JB2
z5dJgBGkRSNZ9ELWTasEkAua72Kb26uywzpAIUud4HgU4ohdQAcs8vA+240mzcCb
2sGrGpc8SuMPr1J3J0cNQxzKUe8Z5M64AzrwsK33O4T0qXsYHVeO+rvQOQTlyvgs
VsRAlSssPO+GrG6X6W70xoATWNbh1OlfjSraQ9m1aFrUbhb+hvK+WFvEiPH7iRCv
MJa/SxB9K/ObLIeyEPwbSNPrWPPK4URFc/OorRKpQgOPIqrRI1bZjGC9CutYRRcY
pwzXOah8fyNEziunqZAKoZ9cblma87950rhd3dGcIq3UKWNG8H+z1xNsSGbB0XRr
bdmLEZm6rvWV9NE7EGZBvQ==
`protect END_PROTECTED
