`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkIfvqTxWsxce4KDnVms256ef5exY6zQxBn9mQNH93Yx/M8H2rfg32yPN7nOHtbM
56wrrAuvG34CeIJgaYe4Oe6vvsaaczB9yQt+jQl3pwaA25kfsWyYGWdmhz/VojoX
JO3wzbTEcciguDgfEm4OHs7BWIpvaRbPQEgMcMxokZaAvb5GiKjVJWKMUhJI78SS
8ZfyVFfpC+7rExf/+46KaGY+OLU9JsJDq9F4tPy4ZaVBvqG0gpYR5pfC8zm9KyfC
XR/nkluTN3BagnkJ0SRzKGYENnyMFcgpvgNXZKtzMdYfqOpds2sh1IlfvIZ3iGso
J+u9w8dqK9DKrFmFoBxg3jOwhnW1aUby3Cz/URZypaliz0GrBNrgQjzsnyZPEfCe
fjOuaKryl21MJwHkMZHew1gtCBGhpLN/H08hC67YFjP3dKMYnirOXN2Xexi7ZMxw
9uWtxZCpkwdnlhgRWVp5sISnwe3eIdKImkt4ksc+o4dOeGBs7nnsmlursBjkLmiM
pLjCRqLmQqTCqsHxq7qDjNYXlVDUQCR5yI/wiHyZ9/gZjA5nYwdRyAOq8iMPvCBY
BPdIQUFqkNkzSKulWny55/l86Cv0PvjNHg1Fp5Qt0wQvJNS2Dwc/0DRCCiO2rbKd
vKgT6tikfnBR9rwzbg8fO7iWnzNoaZ2NjgsebEeAWNJnCWIt8JsVAjTkUfqPi9Bc
/tGhVs8YoP7QKhoAZxTjkoX0siptLaUNE3aT0Ki3XsgJWCovGGBBbexrn2x+xtUv
QgDXIGgxPUHhnY95r6b4JfjW2onXYijksIojIa9tNcc7dBH/Y9VTRxLFJkPQxVH8
aRbqPzEujJXSpZPqcAeXPsas67bSYach3a5YINyKaxHmuOb9f42DFRbBWSnffM+c
3OU9ukmY8aI4j4WZiGrbMXBgVaDMm9Qp2sioloPLCToxmJ3hdzMu+KXEehIdJIEf
02lh5mqrAOkQzsuuR0qLBRCUYXvSBn2v2bWZhPIT9w88TeVQE0hu492Tdi5hcYKl
sehwrRsw9iAH1b49isdFGFqVYZamBYSOoG3DuL+NJxMPzjs3OfSArUvPs3j5Nvfl
MLv1rre4xX70gOsnGNrYhK3iL72dKjy5iBUKOVjnXrkPUF3CSilTJ7BY29ZQqIZ0
9S4X8PaS3ToiRr+WHT/ymGumptXuvEp4L9sNAlXw+5DL3EgnXpLwOhNl/e6P9MZJ
ykngrfYV/XIaBdmOgxf+Gqmw7o2FeKJxcC77w3xMtmBpre0PImY2LieS/V1UNSmi
ZmreInNrB+NyGfO0pbRNoD3Doye9iUyeEBcni2yTR+qyhnJaH+/sdWHQFzYzTleu
xBWIrs9H/xh7Y3Hqbz/vP+LHRSA72OEs07b3E56OOae0Ah6Nn2M3FfAj/FwC4/Sf
EwMkwSV2Yt5Zod1A5ll8ppRIPmBWQP2gNFqV77eF1J+fewbefCtXLT2shjnwmE+r
6ouvdIQYJZZs4o42vAeKMAF4lopwOOKHnAEDLhu4xt2wRUEhfY6gQlTPL7Wf0kB3
+A9c/fONQQDYNytGTyeUJAyymROOUj7aHDeZ0lQD90dpjjPud+FcrsyrWQUt1pTV
UZt8UiwhckHC73z/NUC7LNTJF0ZjJ9fX4gdYodh6s096HXiFHOuilrGAdZBIxZgw
PBmulkVhrXNQGJxHu2zq3Oqh9Ty2YFqDHQEs05kudxeQKRIHY/iOvHlp0XG6bqoi
HX7cyxttO4bOUYYKR8WAuKSvWJEvXACUuiVOIxL99M0PStETod/2S01W6ficVKsi
`protect END_PROTECTED
