`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3a8G3YZfuJjyc5J2roYGJ5oO3R8Pex2Mx+M76tmeEIr3QiV4DP36q3+nA2qMZeB
FAnO4w2xfZoU6nExk/Nl1DTYdIlIXV2rT3Ox7k9SWnlUGNmPllAHIT9y606Jp/gl
kr0lagq8cqDqsfCTMI+NNFPxUGq9NTt6bivmH5t3Q9Ya6soZf/5Nvc058cAr0DyS
shGoGaZC3fnIYina4lw+O9bqkQTC+EfYvyxiaNgiFAoGbewcy/duAy3ajK6jQ7EY
bBIrW95zYsSKKPJFch6ZZBzGOjYM0U8yyTrBI4GKG27KpGgfQyZ4OLUP7glEx7NF
IyyFci+xGl6qmPNg+DHanzf6bj/T+8RBkJ9lZRWDnofKuKRasJpbx9Ha528YmSJv
BhguW+4lZF3qh2FCu/aeMY2GgID71ACMBZFGcueKfhGqxPQtXzDjQw/ku/3jfuCS
239eNZ6aebxYeCcJZdPq6qtzPydyvpeaC5NL8WUrdx5/7Zz6I//S2H9e4ge60NaG
hOEE+cJSzszG5Y6+MDNUpSyXBQoZWVwtv+w4UuG1eD9TwZ98RqyRwXZVSJl9HXIx
TEqmsJJprMYKRu3DXj47jc13j7q3FVzD/i/GQpAxMiJXYqE7dc2Wn+j0oKI26POT
+WfyV2hc3qZI/B+v9QnPnbk0SdNS5F7pJlek5tLJpas713jhmweNOJEACSlk1Myp
ZB0gbz2MjGjKlotMBiwtUvoAbyLv1Fg5Ss/19P/CoSA=
`protect END_PROTECTED
