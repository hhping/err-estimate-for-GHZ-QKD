`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gt+OTcJjE+rtSrxakGVpsPE8xGoqjPNHrMjeMHBP3tNb1AKQYLsThgeJsp/JxHlA
UfXUCNd7wAt9oni4iDurQOHgp6YNWmy6W4P8XIQNG16uSwOyiquF6yIQBvoYYOUn
wvYivWZ6zwC9xQNus76a4g6hPsGwxrstbmE9xzmsmFClrIv1om6yfsGRxrPTNQ4D
74TVXvGTVEcs82jKPGBwGi2G+7ohXxZMhKNQ12L15nZFAuGoUZqJhO5i4ElOhx7D
sqrgUfKwo8Qk6BNNO4ii+2WdvUKQ4O/G4FfoXQJYQnzaD16gngibJojVg+UGWWKJ
rvfm7gwMkLEHmj3cFmnJgYGuibKnFQ2PIMs+w3Z5zg9VXh/okYV+GGvZK/sruC6t
YDtbvDggx0qBSdYWBBVsyQqNKa1Dvt2sQttUPnKTF4i5ytccXeJmria5fjWUUoSM
qwihQ9hyENaAQCVDWO3d3RRHDw9Pqj2HHKtRjeRRcYVqZ9o3BXMzaSSIixjSORuD
ZU1QF16kUYjY7Dn/fLYAl3XX18DmuyXOLQPzGvasljA+sVUA4UJfw4nuUcOvVn0R
4AyeNEoYrpmwgnY8ZV1Vnw7XtTUNLBr8mSol0tWuF0u7qTU+0DefywGy8yi/nhWW
R/8xqvOJXuVxCegddbc8/Hq0pnbLr7xtB8qcIR7Cg5yBGL1QxYFhwXTipbFcMXSE
9j3yMVLDVZXd2hHQx6ZDWvPzWMdnRSDF6hFM+jeuf58s4s9/x8oDjHNkSoL9+unj
85hdTClYDV27iW7kOFgNmeUkxwp9QYMV7U8tIvwpqOKREojivK/nSRm3fgPJuwb0
b/NUBmzc8DYSRQ42Q9M7mGp/IDbJaAYgrZF/CXFXttJHfY+FmghrPVplyMMVVlYU
NL0yehiDUAaAq53xWPS4IlOA8FJT4rCUxNo6IrlaLorkj5qDLsoo3INeQ8teWLqt
aPBqt6BDJSpjnoFZIkJmbcXERu07kNtFlGs4VJfrz/FVcWik7IaMTzJT1S5TqUyq
h/S1ATX/eSrS546DFPbufw==
`protect END_PROTECTED
