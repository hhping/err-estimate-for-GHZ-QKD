`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EEbdejLfnmaWzsek8ejcS/9GulsK5S8akN4dHEvlVYtGzUZCzxbF1huTSfCJCe4h
I0V8a51sG8kTbDP/PgQZjnm3GQIJkYqWenETMTYGNXbbKgo+HlqLmdoIPRLDreiV
uytBn6nAhBffO9KIF87IomUFcBqMvf2MMNKZ/mYhC4rH1CVnIxmVxFQ7VcEp22eS
6ssIdIFzKTVYWERq6/897495tTXO3wN1TYmeULWUWIY60YOk6H4mhVfCHeRqFOM6
8Ksx3zom6iHniTjolgydYS/R13mqsX0PKSROWfN+L8fKPO0ZXsHMW2F3fA0xyVJH
H2JoLL1xT9pGtgSxVxk4aPtL2DjrzL9OJso3b7TDBp1m/xCmQuVV0aQo9I25fHFY
19fkCvdVfj31xZYYG+7sXf0Rr+MIfvmFemZi7QVjkucm+bBa1b3lYX3ZaCVSmmvU
K/aw//HPv7aSr5Ecp84bAnZsymz1DWGxABhkItMFLkCpmcycZp5vs2/6rkp7pqIK
iN1n548SzhTp57v4Ul2rbfSdFMoXtMzbCA1jGlxn9pIBcLIUgez7MdQBed48TrO1
ihsKr+xGK04FSkesOmom+QH7zNT+0OUYDMeXwtWOLpgSNS/dsnKPur3i2qdUCMiR
qOdl6AkGpd9GAWAMzBNrC1ACgUEqY9Dwf9yQM884M3RvTtGXV6yxolimM3+A+Jc6
3r+I6VPQvRKvIxfW+kf+iWdO0A7fSnUNcSTWEFtvxa7iYlsWimULltsDZkc0hiaV
7cbJS2FGq4NaLHYkOOgE21SSxgitQD+bzGCdKNdHxxgYyIY81gCQh0qvTCpxxnvZ
X85fuyaTgiXXHKAE8DejhnzxM6NeXWyRCWpvDL+sKe9xxDu1TcHmcNs8v2S1hyZi
x1LeqJG07TGgWXWEXuR3yuyCFOhIxGGC5Q1Ei1G8ZSHl82skbby/srMS5vDGgx3t
nqhS5161xUSd3Qt9RbyqejrGQ+QAKcpcIrID/T8T0LqQMkU2BkiemtLGUgIct3fh
EmQzZ76qPebuCl5QbgizN9WiseWYp6c2lVeggjkcON2fjrDq71wHfVVtuz8fFBMO
w/DFzs8w5moM1BzfefaoYbuCnoTi+tKGVPJSi6ALr3ld26NP0gmIjS/vg4amPSZl
CpYxaXHIIUdenth4qE/l5x5YJPynprwLqIJWCZMp+08ZdJmZRru/CV3ECDMOA8UK
ihiMpIUAyW6rrE1uZ1NDktbin5jh4Pd6FPKbZ3xhJI0pDcQfVUbRRVIPvNpguOmb
H7ZGxTJHUGbmijbiwNsUTicga2xxmWQTkyvXhYS79JXtKTP8msk3pVBalmgiRJPd
IaRHgqnXuDt9YasN85BfXZU/+xRHkDGmmpQOvxf4X3JL5O4twEN/TkdLNSI/H4r0
o1nbUgWAebuJkZEHbKxySYbVsAW+moFbdvzOsDwKeKuw3f0e37cv+KMAkN/cI8xc
vZ/thRm240yN7kK9iRj+ca3Ch2yAMT50yCY47YKMZafHjTysHawgV1RRqN2RixZI
5jOnFxBCoeyFHigMfFeOI7SX4L4Ku3Ps94V58srmMJ3z0TwsuP3GjdISisads8U/
`protect END_PROTECTED
