`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wn5tI6029KQrefseEmRzp6XPLJ8KRD3qy0P38oCOzsmj343/tmdjtFRAIKheNivF
81xhl8QFsAXzhh6sdasloEbWnkIhIeUDKear44PDvDbX5+yzMU5HuU7eNu0k6KdX
vBv6ftGR7cMHwoWX9Dp5MGkByDrXlrimyF8M6svkA3yd22UZQRvIalhlfihHdh2F
FYp2+YgST1MZXLtZueGgFRDhnj/1onOtFBzghI1lnn/uHFrq/oG8JDbWN0nAKh3e
Gb9UKp7215ZlAXbbaSktd5+s1Aoa4hVz+28/c9O4651RRNxLTGdr8hZAdXFyU0Wa
EzPKHPJesC32OM9R4c0V2odDhmsJmY5Czmz4YdksWEkHSU7nCXD6WSPVlAS2DFPR
tM1BkWFspoQdcWDDVbZBCxfH6TtejACGnXUS0xGbVv1q/e4+aDg3GaHsmcMFv0OZ
8A/PLoCQZY0m2UlhiF/smeFqo7lWMB/ULcirTgjJ/HRe3vb5oZkLofvZYriolXKO
kF7YQ7ILHG/lmotSgbddWviTFS6xn+pnR6wZIBLCNRgoSNr/zTY8oXd44eahzuGl
aPTEJxl7feae0FUPq0teqhBRS6WxaeLmF3qZOsJGY5OO5ssd6q4AycDiwHeIZP3W
3jqUY6sKfzctsoz6Op3KDVdEQdCZ+bRrKB6WNisyF/dkw1KqKqGVzAMRaVWq1eoU
idKSnu7SJmNiiK8mktkXGZHgoKbBxz8GSf0fWRBy2qGekJ6soJ/rTvdKVqOC+z1+
zN+7jsi6dw6gG/qDYt7VkpDBtsZbyCtPvI2pSJz9gdq2z+iMnTR3LLT8Rv3qq9Zv
HOmE5tvPBvJEZW8UkDTNTHVUyAv1cxh2+GbMdMkz4j8znbIsA7ESarR4JWw6j2Q6
SvzyqhI/AWwZsJoQIihhuEdonX/IOFr1qjhOJSN0WWbo8/zq5guTlyTJlCnXRt3H
Eus6czhF0yY2UpO+YNAjbgEVe/2oyBq9JJgVKPSWczkyp6wvJ/ug322/0I9YJ+Pn
qKyYFlsWclAzvAtXmfOMJLX/YcNmdDmD1+2zJJSJ59M6Da4jce0WQwkFjBAUDFkr
HR+So+0ZX+R85C3MdSVBZnCTcJcWTGLctCFoqZ6thmqwnAJYxki2QDlBQfsxfww+
rVa/nvl7dc9hIb0C8EDuy0vYUqBDIpZUzBDAmMLobL8DkVSKyIVLEe2L4dqNz4fr
ztxAJoASV3aQyairNmUlmNbY56KmlxMtCNMcwDpJfRQi98FLLmjJ61qMSjXklOBy
7QmRSIFRZwT/wYb/wElgeaSjUK9GxEaFxOWInaD9e/9LbWZuTSQfGCvDFFpTwOQK
VzILQDG07pdhnGrUur/EyFWaeWsr7R2gG5hKUMqkwSy+1Q/c4rEhGPBuCHr9HcCH
v/d3iIXdRCehEUPpOmuXIAovN0wy09qhGQq2jf72xeDC9iB2/w0LSuZH65cm2FN2
VkW+F9NeHWsXUpfOkMftT+ZbWP2FLHJX2g9UyqW8EizGk1tevOJ7UZ49fQALSQdl
kfQOCYiHgJ4U1fJDxgYqhG/BcBwVCqdfaS6tW9eLirb52GaCaTlfOMA86crK+bvX
kpIytfTD/YoVqLVLcIK8Vk0OzJt0vbOBeQGqbLMO1IRR0TpyveXH2t2XNQEMHrc+
n+QAJ4j9YecFwUF9j0cqax7PDiPaSLWX6vsp9CGADZIkBehb/j+fk+O7T2axVxwh
59Jslb9Qp0qYmY+ylX6yPj0pjn6k16zKTDj9r1F44naanwF8GcRHLklfGxWeRbok
rQFkG1dG4pnOnpfL6gGNXlIbnypJOHEuqXNBGh6u2PzRatkMQc7SnxE3tWYwE4zl
lc4pkngJKdHpfJWKtXUS2B4/ocyvkksSgZAo4sDt8Mmv1lSR1LE4b0kjMBO9PaqD
1L8SP4s9B1HrTtkk3D1ZqJjZ0m2jtDZmW5cXI64iiXRbwJAdoAeHzxYtwJtW7225
3D7C50MXJxLBBNaHDsU1+1PKyNGIGQCKfIEY3i0AN2Tft5aQqeWLLAbwmi6Bqa+G
3hzvvK7yKK02cef+Z08TY2VlIhAn33eaKBETlg7ijJ7GWoyNNs+VBq7cBOX2+olq
lPCNPvFsr6Xj8DrOF4x7edVxwdOSY4LbTQta5gazCAKnyGLN8EBOGb5Q6QU+oG2F
WhcuPRucmu8gWcwtxL0BTnkgl7bu7/MUvgcwHyCFoCsayZ21WnL9lbsdb4iNqyT9
k/3to2sJNxyGS1IPWaLpnxqw+PM+u+0SraPlVTzt0bEIyZt8FoQtabEJbviPzwW7
VrrhMfWUmJcLxIASM+yj/TyCNOrpvfrl8R/mQdjoS3mV+fFCTKgVKxxZ+IwnQvax
SsPev7bAXiSZC5wHAZRn2TIk5BVyiwTtftDf1UoUwd4/oqvCrvbLqBX99sedvIm/
SI8MI2YvYrEfKdPI9rp3DfyVlk/293pGqDrljATMU1DA7gKLhvIZO3Fwpecddl5p
uNtpgxdW5q+p4q0wjMTGxhSQ+ZT3KcyvHuhzH0wuEfy6DHTOd9/meyRPYMtAUCif
lOzDaIeFY0AEVzYsVqyswOyuSO+r2SEzVJvIygqo/8+7dVwo4kzA3aRw8ihePzsk
lWRDk1B1lvearBb1+LYXM/aNQ0OzaH3Pfv3zHeAEyF8l8syWmTMh6S3tNz0n0gD/
F6WyXDQGSBkaecNVei3jyNQg6NQrmINYto+6yoCXYCqNGJaE6uGids/1u4TWRJJv
ZFGlPbPjL/wjShNCV29vIShmrdG62vlhG7aEjwoCxttcZ1D5OzehP67UOnOq4Ebh
qnsnxCEsyriqv5nVD4+k77ZGKJysdBgZp7ymfORuAhJjvDWT77SOVoViYvSMKWIE
w0l7at1j0TJ6OZNmgB6oKXsY7CjfNi9wiqSHXrUFLwvKCjHU0q7k9FANgctCTIb4
kZsCxskz07IeVVW/QMAKxQSEq4QqktlgpA6/tHP2dVKZUJ/y/qQsNgjcO/fAnHKZ
aTKqCPqwBHERa3UH1MzQiRq1r/pQG2GpfJVahrdyWpPVYoTwFcXlzZWDbWUGyoiV
V6DurG6rfACIHMj+9ZKOSXVoKBulvVuDtfIOW96khOeVjTRhTL/pIchXx2+6ha8B
0lj9yA7zxZmSUQ9trgI/QOLEUmCJ15VwGnDUdMQNpc96moZh3zmHt9KDQCOYXTrh
QdXxUGABteFWpkGA67KAbjTw/U2slzdmSYkVN4DyyCrCfKv/MWBVYrzOTH2iDCUr
WfWcsgDO/YyNMPAybuiorgxYAJMcUYfeoxNg4ZZ3J0Bz5kEmL/EPUZVoJ81aXdtF
Rlv7Yfxevi0zQW02HZEOGgZjR6tNrY2kZzkx0cq6Ih7NBjDPH65yCDDJE5AAVrGB
9OGTM0ft2HKi5YwQy+TtpHKP+Rj94BvaDElIf09VdIvs850UmMLmmanWXr5jkUPE
fgD2PbZAzg0udc0N7XZmyXUCm4JvHnRgglbEbQTJmTeeFS9jTOlHHoAWS+Ah8R6H
KdgoeBcW81V3gX12SIisOz1dqbZhN/VXCK8Bnk8XUWOzM+R3WVxVjefFFtzpCrpU
PZFLUv5lrPLkz9KLQz52ruIYFe3ThxLohN3ObT5Em6uDz7mGXm6MRBg4lWHLOLkn
fnFoxJrIS9sC93mk/jNE4U0vt9hQVm1WI/qJ1OX6LVc4DNi1RCwf08mQkH3uRz0l
FVdWbsoU8uMYsTME9GoitNXjrAJxXxW0PYTNsi6PUzEqRNi056SIuy33vPQ/RBDb
EVLM5urU8E8eEiH+AUJTeGRJjYY25RTGoRCnguigVWjwQ/ZtJukIvo4nYqY7qoFh
zsZXqwJ6zB6s+G8VY9WHp2hTrxFNZ9Y1X6Bec1HEf/gesOCR9IwBWszgep51jV7E
A6F92ASpWJjoVbYOj5rGg0KJcGF0UGV5YfrUAiku9ko4fwdpHmbp2GFSa7AvMwoE
Q6iUngpTO/rooRD5yGYUuQvLW88K0MPDGPIH+u0lxk5Hd8Cff1giQyMnTVtegO5Q
5XgQsNImJQWgPvwUweztWCQq9QqYE2hfpCUvO6vU2SW31LJhCfoZXvXRNFWdHK2+
vNOJKDV7cgOzVP2wHRp8m5vxY0OXj7fStuMSzV9rOoJOhlZXI6hanbqW//YEIkRH
U1QQlyOvrE/y8VOKf7dO2MbUUaCZCl9x761Vtp1clHq02Y9haqnsvcun52IJ+giM
v3bSvsyaTGm8kBqeyct0InAWOEMtlWs79+iYoddxYT2Ml9iaMk87d3xOORgWPkCH
X77K9gkhzrgKF2684RRIAIgTAhxjQJqvKwRqSY0TpQwRQhkNgxVGYuKg/v1FFbpM
XYrSp0MNf8fhM9RM3Z76Qz2317E92sLNAyGgGkIpIBeHAFcC5r1FhFGlaJE1eDKp
nv/kzMsvTEwUDRjLLNx5xeenwDECqX4UUMMctgYjUA5nd6ZkDPDq8MFDP4QbJ1Yt
BJTstxhD3SLrLjY2XQ0qUg3X45Jl4uhmi2E4V4xzbIvmTcQvPnT2ppyuNMFc0M47
MYKWE+hN0HLWFe3DClYPiFYDeSVA6VOhH+WyjbSfnfQ+iEKQjDjd+OwuiET2gX5L
Ypsg8xYdLnEcQ/KVM1PWRs920OcnRjjJJ5oC74w57C6liSTaPGC+544kECSe+OFM
jKOhbtN1yldAph3Ym1hdbnkqeajCfvtzFu0599TsjEfA/WeUZ68gb62YD/OkvDTE
gEPOaNtsjOQ3DXbL8roy7jyHNs/l3fB3iGsshdfPSfZHcCcN1qDutdJSVYZqD00u
LJ+ghzkrHFvzgra9uHmQcm0f5/e1MpnGX5/BZylcWYZmIC5BRu6inl7BDTl6YFXR
31FP9c02chSZtMXGSp+NmnQccBIrjtCMDsaF6MaZ2+yovq5t9z7o5l4+4vNezbk/
x4p98srijGMtxzH6LfHMtvA8n/mjn9Sdakf3tsV5GeyRXEvABg9azglD+lY2OExQ
MWAc3kw9GTqSSk/NbPWxl4Xk7rmH41zRPWnNcKKTKHqaBuw6OaiIUAjFuOuWguVo
w/1zY/fwezVJiXGzTPkwezYzGbcENdUzzLqdV75unNHnUAzYER6TEvlknVppZ9jK
0BnUrCcfvgIjHp2nouQPosLRjsyGphDG6pWQtK5kVdHwksGs5/HDr+0K41wE/Ist
UeBgcvaIkenJuoGwLXuZuyj5qCFRc9jMSyx9tL65L5KX5lzmYy5UW3w5merLqcNd
K17ex5n8euuzffseP32S8WBicK+B1j28AQD0tdSZNnUxU6f9E7PpkoUN0d4x0h7u
bJ0ZgxFH1loBBzgWjchD94armw5giAH3ir1aoAAQ9Rdnqy9NoSEcrfllu/Aj3EFO
Q9KEqUP0SJP9MLEKx8gjp3TykPNWCob2ZDoOaxsh1W0J3EWiAEg3BgZNzr3nXEXW
y+IyrMm7E0JIxspR3RmA10ipksf1lhdmqUJi3uI0QrxR8rT9XcZkK7uRkJ8TmEpQ
6OhAbz2znl4oxCUvgWRJ+nmwn+qtRzCT5HthjOb/Lo9QL3ZlH+cdDAbhVGaAO3ds
iyFcXMhbndt2331hh6gDOjB50OIW8fFc/DogTCTXNusOX0F57jWdEAR9W+pt7u8n
wo7AIK/cSdnUI3mjskI324nhcYDfZqZEXbnt6ZIBJN6mlfLNs+lALVs0KjVqVjIw
NrqTRn5p3i7cgrci5SQA9175sw7afvREzpZr4ZH0EBO77Vehxackx1dykSLLURoM
OY1MS1JjKJ2UaYda7Nat8BDHImg+mRb5GajTFRcuyD4GCvZEYGoj34csxUpzALhz
Ci+eF5w9HR+GaAyGEuxvhmDrzJRBrOQP0PZBn+k0zSj/wzfmdEz87ym+K8Qe1rZl
Ukzcj2c+kSVdgCBrFt8sugEQ0B4bpgWTrUZhDpx03bpgniRDeDH9Wp6c7v8D9Nkf
Aix3m87dyCHNZRwaen+OgSu/iIkNMJv8tffSCHwi5zvtcAamzx66jSIW26UAWlV3
NdqTvntIKaTSla4+YauPO4WLt2TY+u9g4uiw8knFEU8FIEhXKRZ4+fKnihoFdx54
Q7+J/a8eG7IR9kb1MQSrthYdAkKwLGkaLi4CJ+ZI6solDdIRHFxpyetapyDbClok
2Tu/8KrEFwPtdHfYXaGtXg4ryn2dWgvUMZMNdllbtx/yF7BUXZf1czsEly3Xj1fp
TGxvwYv2tLd4sZIZo9QsOdEDyhV6xnfzd+16aNZ89r1MvcD1L7eltAw4YiAbJ/CD
mo/ZeOYA2H3m+vNEIgsOllpVaoCbJT83oMRcziFtFbW397Vvrl+Zjtmin1u38siJ
Vs5TqyS4h2Cu9Z7CIbH6GhmYbeeEoX6mBgInuEevbpRF9NWjsn2jyFTRSJ7FB4dQ
dbAbQDliSI/33NjRryU23YZtApWeu4DzO3rEUYMAvcypZ2PIfgFmTleRRCL6Ead5
jlgI88SKozSiL21c3MsrQlpjrajiicxQ7tc49zPoWHFo1NkqywnwqbpT/rPnkIi2
K0MQWerrTJMa3Ssets0beqKa+Dc5RTmrK8/BL72hoow+xYOUiWm7cAyq1lTrR8sf
Km2WcE4PNoopDgBm6rQDXg9hQl2QPgEYbUcg2kT1k3I1GxLDkcB7oDPytI3UuIXm
E1/Miw6TupVDTDz4MwadfAjqzPZJ4cQhfGZbyDgw1rUeE7Cui0o1a1BAf1pPrKoE
fUKY6ZjNmrALVAX9/BtqXPEXZqU2niCf4oHdDTP4oXKRx1UOaAkWHcBxP2lkbsfq
Ru/uZLX47qc3QUofwEUPs2bOLrNr3h6aCZffA1vK98MwdSKazf+IyXVsMkiFV2ck
m5eCnFt40KfUFlpLufVBMgRwrta8G6FaASpRc4SEIDf9XOkaO4/eG8jia7wH1bZ+
XQCGzAT4PP6s/IrWE7fqHGzvvMjFCNNLR6mGuiJtTumExILlXGugv1swmaOzccAt
RJ7Z1I1ealMjMRhEHPqcS6XnIQtJlghU46Lqpx4ExComaeHOLIsLmYODnn3dAqY5
vQvp6Th5C0qLg7W81v66/TCszbdAQvKU3tSnqGbp1v4G4oeQl5zJN1dPYmgxU5wD
eoa2lZ1nsMGowULDW5tOt705CnifEb6M/AOsP4MbraDIxwiSqaqrVUBt0WYwZejm
6XaWWNnXKWrbQ7zjawfwVdEI2bgsnq8dKhrDLXdj9Ly+aPgk+KD0jOtDSroroBb/
M1++U95ZvldRoocFyTy+qNCUOvDKXr9Tm9gkGfvyWOXKPinG8F2zqrpk/4wb4AFU
gZHiiDx9AdgMNkVO3Fa2/GcHclPoTYcMaUZoWuC5e5uGnJwr/6VIeHlpPgPr6wyj
D/mlv77KaoH/VydEQIs9jTCSdjXunLNcY7H89OtB7QA/RdijkQql7vpvGc97254b
bS3DKNyAOBLONaRdkM6tmTtD3hLQJCooc2iFzEzaqSLufaUygfZxN3zgoNcevzSV
xgCTTsiKF9+gviD9U1NDnr/XUf985bsDVPwzVrxGpX6ffcaGmS8S0dqilXqBD2KY
bMxla/XzdQ5fxKbxiAGhIuY1J5B0z1/dPvA3wJmKK/S70H3fL6wzyiWhpTtNYYW9
lvmO1bL0VLfcj46Z9VNFKSysyAxteff1a4Cw5rFCYFk8VZq7HMKNq0Jm6RI2sQC0
jQSdzBJ8RX1u6xMrSwdRRDGZaMpnsNeXymCaOQxfkevg+BKfm51qtwcuppPcyIY4
nBMy73kI+yjMnj33h7mVeVD36gLnrlWi6FwCDrBaOjpbAECdR6soXsl22UsNZMdb
hN/3kOo3jKCbFYqbrwQFa10XCLwWGgVA5J6I2tDSAbJ8NJz7Q+gz791ILwnDC1ju
mC53GP+/sOEww8uE5Pl36KynGATa4ZNjsN0vLPg4moY/RGqWfWJwKKQ2V1AM+fPY
iJB4FtlVXTPCGqy6A+csaju1k5AB5A+yhkiPKOJeg8/eltIsSzLPSiowEeVJ8c7G
PsqwE5c2hnjPTS4w9/+3cpa658liSyW5kxVMdBQHs5w00SEc6Wii0ShioFPoY9RV
li8wRiLhxUYr8V2sioTNwswe7KiSIfTO1p1oaD4TpKZg2QAJMBFbXEOZuuCrHbG6
0l8ba7rm53CDzsncs+a2vH1a0YBhUmlsgFE8dyfOYIMXtqJF3L08yWnP1/RmzPX1
tz8m7g5ADiCBVesa624po8VBlNMvTGsgOXR1waK+VV8MhDkZ4v2sCqUIH5AWftDB
USoNz7xldKWrvymjsBCpP9ayPhIUraXo6VLcqgSocfyPTKvGvTfWymcWM8/i0Fs8
vQpIn0xEezWMZBzWLxml/9hbDqAC98LChwcuNW+6/2H7p57gMkHx558hLrKovLVV
Gha6bRR8X+RPmCHhxPlB7Do0wLiEiQL/QTVkX+euC8//GRZiPN0M39bEgFaSrFpR
ew1my+LBCoxByz/fKDvj7ZehBNst6TXqpuaqiQZ/AJrrMFKnFwWuqSjyMx3hxUmk
m6h5fKTmSxZRLeOrFdLKvlwxgfeoJ8M1C4gYQ8wnpnnmTw9uO5xkwzW3sqyVu8Mp
P0XHBmFmZOqIYUJbjhk+VDttDg7A2K86qKIhOyHK8mI+Pnz6KTh4CuDExj8oQGGI
d/sQsX29g5nORdJUmQk4BPHvG+lx0Im4Abj/VUshBagx4Ntvd79oWZVH/mlI4MPK
bIDUmcqnwoyc8Q2IxejlBnP4+H/ByiKnFSziM1j/GJXMRtg4CdBZbzk+ZfKZH2Df
RJREVI8b1Sc9ZmPkC+cJJqeDML3wstoBlIh7T986eKEAT5KI/IzP1x2fqC9j5WSH
iUJ5iUExev0k8UDZb+5x5/aHQGtYEQLlIQkaZ/eV3OHIEhnFwOLbSIVKktFzZ+ko
hkEcLQtw7lyi6bQ9QL4qNZ0qrd9jkMv0+k4AbIqikpo8JlMiZ/gyrcgnEN9dzOl2
MyvJfmPfv1zP/fMaUOXoGiiitrM8VC9dxD2xM668PLGzGRuzsIDArm6fDEHeg+us
A+FSvX7t/STwV6AAoPFi3OnnWFXouD15VDusRwvMbSD9IE/CYgUZUz4N1ON/a+Tr
rswBBSB+sP6T+Q32np+7RE94boDJUBxJ6QchOHETLEi4dNH3GGTUsDKhoWo+HCWP
kPGsPlSaeNET8oH0yuDtEo7yf/z+oFRIE3VRpGz1OieW8OjrYZebG385PYS73Svu
FvkPes2Y+ZHbQ1HV12bIdglnaOhupvcxPpFqL0ys3keFiqUpCdzeUNufBXS5Sx5+
Pe5Oq0kNZ+kAg5w0XZwVjA3loTbe5zw4qwpPfPIT7VB9atCWJFPgxnDwOGv4zinz
qznI/PrbssA+qPfiepYXRyKzP6NOSjJqOtXWcYEeeg/YwB7+2iDK1UM68HwRB1SW
7X3HluLjNTVeVmd+Ni/oXP6X5Gs+t9FU72W9L4z7QST8QiWig9ytUbxZnaQsGa/E
Pz807V01w85N42lw7PnOHDO9ocgnvktxSAg89pNadKBuyI+1MWIvKy9ISwPgjwAT
t/JWBckHmI726jrodGLYskDAyaJBYQfAF8bohs9YwgVZDAJjfZBZUKxR+Hp5Uw0b
T2Q+sHaA4+/ItIojZ4mMDZr3j7aAoF8VusU2YnhChwDMRWAjG6qGARNVF2iGQ5Fa
54RFfqLa4XtQ7/PScNcuakqpVq6EQOSlieO/l5HVIRKR1xIUevwG4hwjePvvYTZd
EvzespfwHt6MMVzwiiuxjlynciVwC85sfae4aqlhLADPkjjCip0iPGiRlpObiYUD
zichvzIAkilWfRd2oZV95gT3EF0t92KxNps3OCSe6grb6QIgVyhKxC2tLmX4EKRB
e4opI2ZdIZZklXQgQrlOXKayL1IST5ViiRSQQQHwdUfQNUeKXqmmlYRk1gXtO9JH
acAYQ0tL1fiHFVx9/rNCYQa4+CJ6d52lgUsVM9L/klNpc9NZxXlRz9RgEi5JEQ94
7xj9IKbDGzp0N+yYeHQZShbMUgF5PukstxxmLdlYSbjdX2TGnoX2hCOD1RTur+aC
/mmPBGHVvBZc6CnmkwvbJk4w8I1qZl7HKOI/1tFSOSAegIzcsI0dfXu40KpuYDnG
3qFZNk4rRMUrh9JCNsI6aH8inVKRhEfFmTE8XsjQKUVTI9zXxrMIUeGHc48bwI6K
x7eOgYT9gtDAxEdYdU6Xrx7r1nrHkto1fX2wTzpeu6lojRUy/2SDyO8BucYPaU+Z
9Hvn4seB4aXJliHy1hEkqQEQ2Joi3GhOGY4RxhwnCUxSMzka7P9xno5HLF2W3zUM
S3uu+S1PcsXXTq9MAQE+8vE5nmgOwPj1qwf+f6D808hhRKUYPI0PI+GBAa/BcArk
KnZ6vy/GKG4vYSXIR9V/f5q7C0DtXFmfim8CWT9gwUxPIaFR4J4R8W0SjSmfyI61
+8F4aFwf7M+L349VztRjVT4uOHFfpKTStAtRGjE4isjfSmOorVGetyNCgeUiEMth
xtUtY5tGw7/7hkHqDN0PIvSUNqWPlfESV2iIzCgnWRxPoAl/iYVSfiiUk9xV0kBu
z9HbeImOm6eAp7wFun3rdb5MXHbwB3EvRy97XT9PCB0fDM2/XfQufb+BTltQkONH
Jv19CtwUH7wrmmMP6/sMcb3RrZ+gxp3zwIcrBG2UDMEW9NbG+E13ASY8EYHdk2m3
xccPpM8yeAkkz+zwQWDChKswn9/beQQb/qFstamGGWsC3Pnoen8qN447QIzMwmZ/
ZMpNrH2eiLFkoNHi1GSN+K+TGJPHm07K6pmUNNH4TKd1DC/8HxMsHv5QUkYO0LaH
QWvJ8Va49Bs7qvUj/uFBBbayXmMLOEtS9R1hJKPEt4yaX7Xpz/f2U8/FdvOTPFXH
yZeXGXT1HhMFeXgE4miuN0MtG5ykIHMdK/qAGidx+gkz4nZLt730tnypO6OZ5Arh
q2aVJjfpL2pnZ4d43Tg8QGQ5/pZNNvXVebrjDtTw2E5NycweIF0uhYWXMy6KNjn0
4I6skrhOYnZr7vCmu/iguFBDe2SxFeSeCUwH33d/UGmkHFm+KWdPiMsQmNAgiBqW
F2Jk2jLDlvw40qQWU5PN2O+4xedSBI81pAUe59wb+zU0bQeu0iwvbc7il/7HBXlQ
2sw1gsTMval0wjrqlsanv9bFvpJmcOnWG+ZPCLk8osz6IaKfttnOKZMgSmRXNW21
EEw46KgFpAgnORvzgWcti5UiUPVhkQENcXKdfdbbjESU2hSDNkgepYofItATtFay
LEF6EEvE82y3Br5qN9DtUIfYUSON4j3CCjYzIsPtGPPqdb7AqMmudDAuuvKbAfGl
C5w+Al+WHASn6WnbHlqjwMzhGWYYo0QT3M7xls+lbZxTBV5qWFVO1Lg2opr+WiWc
ilK00jNUQMqYgOHSehRttlXybuantGzfAhZoakfBLfWaifjHL0dn1T94VBgg2f9J
Dqce2eV1DSNnH6puxeY6ZGOzls6n+YJirdvvuDz5jnkPtVLZexA9I2cWxfVi6OBv
NmeDCsrDeoV2+sXhpVqpzRUFyc/tLqsxTILueYTTc/0yAVdOilWSWcmvahvKnEaZ
FQrS4iNcL0WkT6TuNuC8+XIWmmNSR1fgaQGbwbnfm1fbrWbFfbCaq0B42xsFR3nY
kSmFbe4vStvwF54FkA+HbLHNGoWCBTbtD+mdWY1jHhcSmCz3LnlYEEP5IVR1ih5+
15+yAmwttIsaq1oIISfTpn57uxCnCyRmi/ZUD9ekRyMWxJyiw7uBkqsXfifLs5/0
mS18hJQ8O8veSmNMk6tYqyu/9M1AGy1Gt0eU7hFQaA8nnpcfApIlPtravaUlkXyX
+Fx9JuzLGjEMAon0nl3TJl9aGMeUxYpKgc0RgtQhiwEN1XRi7TUJ8z72LT2HAihg
mUJ6V9jsPgzCOx6QtDR2xNoOqfsC4hQNJmye57lSQdlvugW4YV+dn0Obg/Tmmd0H
oYXcomf0x2toWiL6KSDU6PO4/4WQNkD9kSJWSp0pZQnCwmB3pEMX7/Qn3NN04RJ/
jdyDDSZk4pydSsPYRhD1uRYGKEkCQC7sk7cha4JbsLvMh/dzwopwFTF1+p0hGiFX
tOakO8AWDOTvTZYJjozWPxcDFliDuR4x/WMt8SyEsF2YsdhScuvzAa2ROGcLNbGA
e5UFhEOJlBZ0tb8WYOwDWpaSyUUCNfsI0MC81dd7MCHfXk9NM2n0S/2TD3GiSDDn
Xaq/XT3HMt4pl8n2LDAlc4DcWFP2EqT1ArzdriS8WuUNJ2Vo0Sa1eCSvBtTAaAPo
4qqSrYPVneCbY/+9r/s8jmYvEw1m6td9A2BR2OZHIFXeQUBs9JVgf5AKqf7c+efE
BbBbSXWB30Va4Wu92utcs+hmT+oatF36LbezrF1fCTahjZ/LuICIz2x0l4Eqks9O
ezOHoYL97dz4RU37NmaRf4i3YwX25HPwkEDWvZwcvpBvDU8C1NdzZPyrd5iw2xuN
X0MxYr9xgg/TTMJaU5ZZ3+i56kZnI6OwA2BcI0Sl9JBbpPgMDCpCzZ56R0+PyCAF
PKxJEa2zIDcDSJMl0wulKpC5rQjqQnEeKJLT+N/vrl2w3m+voO+I9SqndThGHSPN
OysjVonyaOMXHhAR+orhMq0yQKMKTdISVr73XnHqmWkd4KTwLy85kQ2FpxHQb47b
BaJmx4kchd/w92Klb0yCaqW/yO1NWltRDlG74B3SNi/N4qtq6m4IfZf+7o4C4mM+
5nb+q5+KrA+YYuCy+79+3nuJe7X2lnPv35j7dcXmkxEAL2WBKkrOvxMQz8S/W6JH
aaN1KmA6fjCNk6UKkVpr5cCydvpTZYInRaF7sOWYi2sykT/ZoH/0FmSLzGZ3Qzt3
G5+J7tg9YBrOnX9WAwgqGCJzNVzKUQcRgfVUr9vt0vcvTMVMFd1oBBDel9Z00NWm
yYu+CJiiKbPX/HNOGOvh/TkE7dsNuPifPmJf8aOG50bbTmZZX722+1ENR9DgJUq2
EFoRSsy8ZN9YXhXJ4WzSpgvKSMnhYnwIZvm+afG6rvCFlSPPKcTT3t4qtjHVuihf
TgJqok4QLZjx1yRVHuN8ZgRymQmbsAQ5yTsCEN05nbUcPPcB0T/B1QpOOoSboQ74
H6gDAOXDkn1iJdwVxMq0LKkkEOuarJdVP+IwaqR0R/nmtKwXBcnHdRQVPr7mLfdb
aIdsx5xDi6d3ws8KBnuUIQ6ZzYWXKudYufvd7wqngPwaWq6Co/nHBCMgHzv3ddAx
hixpcdf0nGnqhqehqceAz4OclQ88Dv8iYtkhrGetup6QmmCPEcnL5tkUWeWwRDHC
gVSdJeVeQFdDFc/oZJjb+iZGkdqF/yiLDGN5BegO6zRNKTP8Q+RFPPdjLhzyz1Cv
3pWJdkHA3tvAuX0aw9kibmDo7rvDwoQZ56Zb0KRctUP0z7w4JuN6lISOs+kEXeYp
8KFeNBi8dcj+l4NSWg2f9TT95Bozf4hXYO9fSgYbOl09i/vjGrDQO6sXoSv3CyK9
jV2k9YdoqHGFRg0qb8cEOeyo2srmLLaxOkDnj0vYz3hlbGByM4f2lbGfIZX3Unsn
4EANRA6AkPwQQJhMQdkuVAZntzq1kVvVnSGcYOg4Kk6Hw45VoAINq1mZvwhTfdqT
WpD0V8WzfPORNzrZ1WKFxE+JY+nq2a7DnwRSpdsMzDaQy50XWdsTe+5+TK1hMTqb
zPy7JtQiIbmOlt8QmOWDWLZ0mfHM8N0Grec5OCKv7L6xjLYltnBsUG2qTHsRzIAF
REygeaXMlTj9SJXjqb9sJS7cG4fkTP2WojIxXQIgKllyLqMwsjOF02M9nc2JYUeD
nEp4YzMjweINf96jURl/ee2D7DkoK08fJ5bLJ2f5DxCN6Xeld0SHzeGEI+zJy8pc
PX1VhPJZeT41OKRi1UE4Zi8p2cJ8TA25Nht+3Lvn7/Vf7+zkMRXhB5yOZEB4eey1
/Kg1VWUelzFytnTeHrj2hQjxjSY8JbV7wTnp6e2nsGC/wuqIl3qxzncklDiMoJu/
HUNaFZlOlzbwTQz6Svd5iERkDUG62s1QlNangKc4eSBJKKpbysC5sgSeyOxZdX3p
oMYHGSigOmsj4ph65PxC3ZM663PLOjia8FIZITHgT1ydosrgGRhLPS5pVOfvPyl4
7lVvVYJk+ws6ZGnv0yESU5wbwx2AKJEZKQ4IAOIFZk77sN98kIYf8R7tmdfXw5kh
NPG5bkJ5dWP1Zhx/cdVe8YpeeW16cG8oW0e4l9OlkDvJqijNycIcTMMICJDhwm6+
lWIBGBKoY/v/08axMcxwcn4GcR1uBYZIzFRMQPMwi4ODkmrAGQZBLVG5tYDT5R+W
L7m9pg9Kv0tbOQG4wmTGthsCMm9qd4/E2zHQBHDim4XVYZ/2yGUN52/pw9VPsvMB
sY9Nu2wo27cxRWX2VBpoGIOm9dd2/5be9SPm5ZQx8XWtIyAA6Guy3ekw3msNPolj
E9e6YY3GijodY+9wHflB0r2mMIqvjMeOQ1w6S5rUKMXv6JdU6zD+mVGcdUsd0Bia
dQ5Q/n+H4VMV1UU8zCnHx0DNfakfbgwwu+Zqg4t9xeaJ63lgpYJSz5GWdbl8jXcf
XB1EEStyDP7A/oIZSa1K+6DI71qB3bqfscv3qcT8xZU6dLW+gdcy+JZrLRtz0E8p
Y832niyzipYhr4VxJ87QQ4L08ophYoOvy/Nw7GCCfW16NuNTvttcNs8nuAZKk/W3
3V+Otc5JNB6vnTx4qLMFBBU9xmDU7/uDrrNMp2+URMm2sn2VH1xMaQOO7BZHDER9
ZWvaEjXbV6yabSCgZMH394ABBO2wpSTvne97MCtIIkqhPkIWCO/zcpnN5RKJn30G
sdvtMwd8OHWSe50B+JznzvoO3rI6VnMhF85l0nOYjXiar7tt/n9KPxAeEjegULI6
pd7Pe3LKw+YizFtSwJnpDTilFOn+abO1bGevIaU+Z3bEal3VDX7JMOp9Be+FDnsf
PWuc7j+SzD7Eoyk6IioiXxRFlugP+7OZTkt5Bc1BGvcVt485q/zcX5PlHbZv6IUx
BcecR9mdtrIOw0mpzPgGRGVS+Cp8MQdl1Qr8x/r+Vyhgxlep9XPYXxzOu6ushf7T
Ydxu9F6SgwsQMIAQlSdGWibSizApRXtf0wOHGe/nu9VAWUxxfkCoOEsScGa/iJbQ
Mm7RRu1xNuexkLhg6KSbEEyxNtek5pqFE0COI385ltwmYR2GO82XPCXr2zPzluUv
jQnbf94hrj4C6OBWVzxn8b3UWgbeo8l8N/sTJOjVpMfw6o6O9WBrhtqZmshyb3qn
upqs43a9/331xLwtGMMqwxginSgmR0xqMokQeb8uYNEyE28Ij0lzcLmF4Z1BiYxf
jPWluOsbQGyOzd78rEuPjqwnOfRTGGBaEOFpiGc6cIrxPSoMhAGfyMlF4MZKnZaP
VeERfXpH2UbddDKHkI/NJTJFIPOskDRobpGpVQaGfCFIvg7oxhmuOeC8qZu9LCet
Rm/1iI46CwBJb1D/ITpYqLWYRKJyZ58oALmNSZYPegAJsPKBg3oFCtLKmcwS0TBH
Aqmdjp9qwteEoO6leROJx8S/wzu1E8CP8IragtIcPwL7Sy2tzr/iqCq0zXro8K9x
rMo2iXeuoedTK15oyaADmLmhjCuWp5rm15GnavE5zUtQMmKWMizqAk8lkXBbMEM0
xZc8QCKz/2auKkhCFSclHwzdb2J3XL7htRHGF3KF5V6Cd91jCCcVHzswrYo52Rhq
ooZqn/2SG5hMlX3vPfGaORHqSQVMHo6+qO9W32sjL8/3UO3affTkiQ6Rj8Mj7bCp
033I/frmlAt/64nU2mYSC/3QLxplpQAz9jkwfQc4drW5dPuc2YBaFrhG31mfQoPv
dk6D5agRgQJzxuOJFxT68gxGh855UAAP9UolUchhYHnsZMtvqZNraVtxXWt0xfms
Xz0hcqNRquKEsqvG8pOcdkT1vI3naP5IhwXchDk3sfF5nHCRjTLs5JEKm3E9gpPz
U2GfFH8xMzISVD8khhLAajqLdxN6yTy/i7SQsRgntj/08GIm143uu9kEh2fiZFOa
oCsRAQ28AimyA9yH3++JNOrlqwaRExMnQfFd9w9ikoEG8hvSOI9nodLSJQKE8wWF
tj7FCMyf1mwUdmNitchEd8H8TrOjInxGfCIzrOyq6tz1s+68dtug6feMtlWa3yts
FikKU3582w0yKXbJwSmwaUU8I1dyi7oEX2+sFxYC8YiozDyBsW9vS/vwqO8X5MFe
tGGeLFx/CEl8X8AW3fre6Uj43mfKdjjlfoQAm8mI+eqGvyJ2wdiJSjNbvZCoZuGj
4ky0fqVMQbi/NsKyohKrK6v5DhSmVTWZouOGANmk5wru8kiNYKv+Vd1CKCkTCd8l
phEHE9arECibFfiQKa6ZCJEyM++GnHoI6xQKH5LjmyPrsLJr3w3fmxCTSWcF1fPe
MnWse5cMP27VLp0P82twUtpZv/IJU9mP3AvEfPP7uwNaGEhTPa54myQTw7QYM0xP
hV3V+jW8jWQWNqzzrGI94r14p0yhdnSpUP2TinZdxJj31r2/gwH2arA16YApmSPk
8G4xr9H8xhvQF7c8p3Zu5MTn7Z3pQt2zmXYseDg0ZAb/hicp6zj11sYjlhH+9WFC
kiNBQNffwDEyy4R7ftPAoZ3Al6Ss71MZeyp6b/JMAZIECWUKqmUwcQyz3x3dcNm9
c3+TifBDTOH42JhP6ZO4UHySeBpylNSGQ9BvDquCH5NG95KzYbWeeSpwofZr062q
3dXLufd2ZA0vFU1FxdQtIfYJXPU26Np8ogfDy2NZ61Z1lBqyfCpmy4TklaCWrane
JIVOamSR3rMGIHkxMgyI8Yi0ZKcg3PLt5ZrYESHDXJ3eTnittcqLRLxlcVqcK3LL
kP5OttHHdvxh4hmm5IqdKBc5S1oXz2/AqDUwI/KNiFN1wt5Lu8vx44NfgAorXxC6
50yGlv04fPWYOTgeQ39UhJB4ZgiSK47qC0lUAKxEpOOhAPIx4JtwwMENN/xcG2E4
W2RNu04QEGHZ6ea9HR0ph6klHnX6T+Ef0qExCDZzSvNvPy1efm/sMRAIizEuO8ls
PRb1VTGhMx/UomodtGNhmTmBj2uugotoSQ3fsxww08yJ90aQ9J6O7/CgL1fI0fhN
2boLN0P9t6m1tb8fdkxu/hRLj9a4BFfBgDg5HaC8+I178AWcjIlXd26ZeBkI2S/T
SFrAZl04m5Ftwzi5uTs6vvMmYDd6qBYVbzSbbQ9NLQfmmIe2vYqft2VHbfEVsM5s
UfNIXd4B69kJvALd/Cu8Y6bCmVLu46MZA6HO69RTsYfwi5tH7mdTANUfUsS4VWO8
wFcBym698zaFhxjxEpvX65MTvvNpwv+zODKLFQk2zre9iqf4mj5tXr4chL7670fl
Ns9ZxWtLYbEyoFls5iJGU1SgYXoD07mZTD4Y5NFi0XoUbgGDBXS1saKpUJOXXoK2
K1GSYiiPScu1LqW7/F+rXvkmCMw6fZF3ztrWBsovCqzO0jLpOb4AzElTyt1BJ44H
amJkR91XOpj3dIy0EIGQrQ/Z0FhdEnnPUn+EYrWpr8FC5FC5CzryVpqycbw4L5cj
hcBVCTL/cmtwHTn+dp2cHVwDwzcdbdf/pSiCJA+pEn14lh1hC36Ngm/XPvOUSKkD
8iKuaNw8dtSF7Ludgc5jYci/Hd2xkeNk7UjLZ4e2tSnrOHXCg/bwMfoWY85Goujg
oemWNs32PaOVpuecfm0M0MwADQOXeHar/Z7mieLZD9Uvhs01c+XqHNEWnw8leyh0
ctvjozJ0GYEOxJyKokt1OtqU3lXZ9on2eAuB59zGF5xDLLLFz2ug8/YU+X8q8HNC
syzb/9p6qBTm7csjJ6JSb517nlkgHJYzPlFTBqAmIli0pnSjtyAcyQPPMG1Cs0C3
dXVDC4SmA8vDKlPQZIMfczf6Syb8yrzenkSY9Al+uUCFtKYJrJyD5vIXfk/UU7F2
Qjmg+K3bdlHpPpYKiB/ZVQ2MebGan+YFDG8SteRtGexNiCyDIPajaUhr48wHrquh
TngeZRuO0HHHKmYCBUMDm5Y52CmBCn1vuFiW266HQ1YVJx0qM7zb7M3mh0CewMJZ
9a1tc3pye8aClF2am6UsS4umR34WXNaLqsgQB96+99MAP1vDSrb6Ktytu8CpdBu6
V5YbWTnN7T/v597llxiPHeskZrNcPTFN+SGtwwbNzZBa8xmnDMjUYPt/k2JDTKPd
0jdb9JQ+r4tJg2K7TNxdvGkDsChqUHQmgL4193HMB9Lp9jYomgFqURW1m7u7MQuh
QJ7NAinFzRbOVwTaMhIsYCMd8dmj9bL8RWdytjXYoBEjDmUv3eahUzinvkRe1l9I
ATehMAGwQV/murWso756JNypr2cfdbOrn5QsdIYL6Pa7YShOh07E751VzDehpG2k
7k/i3mFOlpQWkfifxb3uRen5/Slj9P5HFcMnRzx6b5stl49PH19aoIsvZB8HFkok
jqbNcgTaDPlL2tNJ+wLgpJRtDk6MrkwkCPRrGoNIZayv7whGcqhDJ9WmWXZAJ0R+
ZF+wnsZyMB4wFRyWHKtkAczxMoPcFAfEzIyJohf71Ba9c8X9pe3XvzJzlJx/QfCC
OGuxk6cNdgRLVFEeKtveNxdOEmg79WfkbH0MA4eWLNY64rlGNWCLVV/veExdMWv3
7WCU+XBnjdqjvR/1aocR1vO8+phOcVspuC208yK9w/sVK+EDzfLAvCTCWI11hxNq
2MOA89u+S7EA++GmfYMa4I1pfy6+u28rPy+YvX99gniMZu4+/xmJbUIfSpRv5dsO
1MHTZZukMqDl4cN0UTX4M+ZDpoNQeMLMPAjfRjh8qQ/3k8nv4CtQBghQufeTwXxP
wLfqAt2HldGmTHGf0n9ot1pY+xlup2cUWqpPOZUSSlrqkBEnPwAsToKhYHf4lcnw
wg43mLjC6m7tnX8he40EuxRaMYNoCgG2h6zEXE+0eYhwjUtYzsMQTvQgaTLaVIzq
naHh/3fGVnRFY/CycYfY7tmxdRvk/tz3+41IlUS8HXaw748bU6zmQD31JeYlMPTc
9IyNI+roOCmRLHsUr0rKAHOzqnXAR1+Zn3OY9wYheE6Kt8tfQgWoHkPxkWmqZfyK
kHiZU3jcTvlKthzFdhpwk69+CMFVyP1HTrtfoC956sMRTtTPtJuzCgA8ggfkMMJA
Rwa2SFFz3jwEzxrEAb6yb1uOLcoA5Is351/pbHC1xdT5bli9p8BZhfbxZ4bCd4kT
BO/VIhEQwrfoOIkeFZ2cGg3TBfr54kJ/NLtirN4RzFV9ZaPO+1AayRW4bq4aTnOT
4ED+iX5ySAi7bEEMiTRdU1TTEjotoaginpEQosVfNuNTHWcvqKsltNvK2j/xEvan
pdfNfaNY8xL3/QC3tiFOOitAcHgUZHBDYBc0f6VSAcwgyZegpRxaQ/30oXjD+w21
fKqZ+Wxrj34uDvrLv3n243gdlYSroj6qmDecp5idd7Pj2kTFD19Jk2aYlvKwxGwA
jEjeKxe1u3o91Jq8oHOO5VigivUlNIeDGPCIOoLVWuWI+5V1MQP9n2q6iw1kdSoV
KP74oCPmdBY3JTP2FVuK3v3fDcbhGN41FDfiRnoXmzlzHchmkY0AIYKRP1KEJqcx
767q2FqxOmswS9UbyUpszg4vnRoFivufDldEn5bc50qvm2MY7CLYQc1TuAorcBFs
U/UIfcE0cag7SxRf2fGRMvImpnBiY5xRWER4MskjWVTl6P/iR0l/OnmOSHVecVkY
0pkL7ksSvsIHZLzA56PQ6YHRzkthjl3C0Isa7vPvbfkSMBwEvlbOo2dxHEHzSHo2
S4RA40cX1Tl8fHhbTErnFsx27zdWjB5j6bZ1Kz8ojwdiT9Or05z0pn4g7FLxn5od
5ZhHDRoA2DDLvHjcT03m/+YDwEwGG1FdnwY4gNGkbiy55kry/VGYSmiuTgEL2MBJ
Gmj6+rFAD/lFkw89if1rR1gpIPPt5ST1GknAC8NWSlrrBRWFL8k+qM5BBHkOoIoH
Xjy5OQ2OIANqpauoezTnvvqqu24C9AHHsEKAetGDq0ChdkV6TGfjYNNowNnBBO5w
HwqMB7IL2kNYtvQJWnKAO/zqq3EyZ97hZxet5CAfsb+Y6jtl5WsNnTwVvOYRAOxt
39LqKKjYMgWIupIgZBj6LWHWQ3aRqAoU50szhHlcO+KTlA7p6a0KGnzn6CcNQvqj
dbDV+nniGMmuqY+SgOPLmbMIN6IO+TajXoJzbPgZIrWvPo95hsYHxknfUSQSpw1L
0ecc74iC2vaSFb4Enj4en0hhPtK+0vONP3okkn1hhD6op3RREBwrGOZv8/wk+Ndb
fTKf7uB1sC8ugp227YZNlEIbE5SH6MO3V0OafQWkgWE3I3DEuoE7kmuMGsbWROih
h8S6cXr2ojzH0hDtaM8qh4t0u3TMoUH81tK5vTVt0LhBWflWaJYesZYYFGOM+Ysw
ArNGKlkhwE+gJ4PiQ7Hq2hhnO4LAqmvtNRk3iZ4Ia6AcpUBKQHrW88pUBIRYMzvF
Rtltq0HZnXo9JDBhsCmWWEJYESuIR6JCLv9SfiM4yzGJO5GewkMR/MVzZjdh1lsc
L4S9ebiq2fUQl8tP+JKBD3XfE3sKRf1CBYWTkfl7xEu65wdZON/cm0V3ctWpLkEC
NDqBZVl3tkbGgJlDYE7MYmeJdx4R2fjbd0dKKAfNqcRsLQzs/hkH62xVMrs5XYXl
9kh6z07t/qosvn5rRDF5uwDIdtN6rOqX6iI9RrTpEOCGeN4Y1lxRvXhUjwtP8VMR
1tSCldmw0/N9GEk81d0knueY31ERjrSEXYHVLTuIzkws61/zYaasOcyNBi6QlyNF
z0e6UdG4YMV1rz053IrL5hqkHp+G4+NDS09NMr+KYdswN385p5oCJGTa9CiNPNV+
+vW+eqBcgIVIJCK+857gfwyGqhX/XuCFo5g0mXXO0fZR1rZM7TEjqI5lc6+452pf
2bBClvPg593aBe4u+/GffOgNA15U2WZlKuwdCH6cfiyD1NdeYr57p9SKZPwnPL84
thsF+bDhGr7/n5RIG6QZSo+1N89GJvFr0xCEzwhkl3lfTA0a6UtDRjbIi76oT/0E
TGKyQTTBTVsXZsqQO9iCF08TgcXYJQPJKE5hjPYlThHBij2bI2nueUVNqqpbrpYq
ai+KmQbPbEczxxmnj1iyI+8Ot7zKSSKP60P+6BBwHEIPpL8hHHrlrFl+mN/muriG
EyCky68H7m/CzOQcRo0EtuGd9/9zMmx7JrmDB8rg1Fz7hhv0T+jliGvlHf8kM/iC
h032JnAEClJNwCtebCKt+AGgcKFruGQyu2173HcUfif5xj2/wDT+LV9HuLzdl8e6
qjrhGv7gEUejQmGqzzouRnrpXFre5bTT7mG6UovAEolovfNKu1FSxuhvh7o4rtFw
UYeTCVD9seHkyn1czssuiTMkABUvGmw5t9xzvUcy4sVf5tJ2ZdF3ZsoKKlZZ+Ghr
mgWtt2IdMTKHIEBtmDk2hwtB4FfJ+NLF7S7bpZHk2osnOlAt+UcaZHvUOHdeUIdR
Awb1OiiRUtupEkJzwFPjePPBb2s3rOyjkpo/c/5sBXsX0/nJBWw4vmWx/WUGYgaZ
fzUUZzF+Z77Rn8+JyZfmAbkJprPBQCG/nPOZIwxZ6JfpExxhpdc9N34Gf3IslhTz
51XW454tZ3sWkJWv8HLrr6avgkqiqMvSWT/JY9unCEUpJhp/ws2rfq5wm+AKQMg0
P1l2MpDI5evmnzypK3akMr/OFG6yTP7UEbFUzvhZDBNeoxPv76+9nKPzNZ1avMC9
iWantY9n9C5VXJmCIzhI6zW2hUHhZC5QVF84hbdPx7umcJUk4QSdTaQvF4bynCUs
Yg7fTFP37Gz6by+FsaCkZwpfIG0eTj5AXgyxRxh2L0fjdLGhw3BVKqFZtkLxawVu
o+yPWh9jxzAiwigdKT4cDlRAg1GO+7ii4IVb5DJd+k3jeGpEmzF4Nut0F8nlqru+
exSs3NAMmDzWxD7koqCYeVIgWW4K1nDQwyPCKFe+BdDC52cVq+Sxvb/1b30I1sY5
h/+InzEyKk/8fna1LD6vPu0sZpzPBeCZ55g2LpU+4ZdVWnBxsxzw8KDaCx70NYTW
r+5fRuFkTw7itOoj34APtEKwL6KVNTHOs+IlfqOkUcEPPNhRAP2C3QFb4Hc9vytp
8hCcs4euWXBBttUGWWPSx7gngSETbe9qAtCfjDTt1sFDcmb6wf7kUyLQXCv6w4/i
igZNyGoPFojiAp4OydYXCc+VVrk1H7ykKVeB4q6LYVDJoyXfRzAOsug8xKUEZM7i
9GUamOBA2vMliBBOSxcVVyenYK6rVoihEGT4Pn055xBp7HV967jHyFyUNP+g3cx/
71++WQ23TRFF1O432itN4cCwxQAQHyZDoBMCYdaRkGsMPzbH9fKdCAZLY5rCa//D
cbA03u1f08nMZ9N9FXzg79naIvQtQ+aFFyyGcXYZtac1A2Xbc93IEkADOmGLoiIu
8DXIwJhuB5SFxVhZPmiUz3aMPdK3k35Y1t04dL6yJiXKr4IqJxqhOFTLlTb3yp2T
DAf+eKtkESUx6avcab5fZCzBdAgenvCcPYcrOxaCXOP70Apy+pRtTVV1lsGWDoYk
h/C8SzJ85M3ONqZgS56Cox80oTBX9Th5R9TgonVpQ69acLhrAO8WbEjMsbz86uqt
kaqQCoztVSEZXmA9eeb6iKKvZ8qDyBHUr5mN8CbNyU1HobpSqQmFUCSOnVWjiaLs
CyWJjPriP8g/kXLJJC4bsr9M/pdV9XA6I/doAZpX6ZJ4md3CjkgNN/IoxrDtdA5k
VhlPD56IQaxR7eg7JNDfBB1qDjcakz4AfBf3B+Y2YsjvsCZ3gdS1ZVaI0gwYpf+1
4LRsJbNz0VHyqERylsNe9hnC2+MWdo+oagKeTZhha88BVfNcOZLsQtqtabe8FtY8
6bHvmthsAx4nbY3121PJFnwgPp+Tlwd4CyMkoHRUVe5A2vAwmWVHfJEmsUJjjpot
LZSKf/ZZV/HbFIRzbSfng1R5sXbfYQZRXD4sccabXc1Qa+xWOLJB/Z4nbHuLo62r
N+BoHroDoICbnk/gEaMO3c/owugUcLRN5mjug++3H+ao1GWNBD29u0Q0qPeNE5WS
NBi8C9ntFtTcegLu8t3s6vf3TT8sxMoEph6ivKo8N5Odg7tizJCEeeqW2SzbIIIr
xQsKG31DgKPR4crUUmwUCyeYcLKRUdfCu2RlaMuus/Xqr9RQ9oRUsPhe+LGXN5VG
LIA9pTTu0lItvDh+Myvvhqx0g6KLInsJmR0zw7iDUiQLdtDw24dijlPToHWcdRJr
mHewBlBOuAH31xBiFVxF1JL0mB2WcotPa7uOX4k7tkX6TyuLX+mq2NpReWW3Nno0
5Gt9/StY4opA1b+i7xsP1EUTip30ev4U539HgY3m7lMS0pceDb9HmsCU3jSmYnmS
LB24t6M++Lp28n3Hd8WvObIaEZwhGJIhZgfJfz+BZSbU639hh0tPu199n4C9ELvx
BZy4W+mXPBINy8DEvZ7kMg3vZZWq0+j9GAa/kpQ0z7+DMFZ9qJkJ955j2qMIIGfe
d9+6vFqJbKEsqJslHTO+2x/blXLOOVxuqJZFK2Fb8YO5G2CZd1lm+rE0Sv/8mJIW
uGVpTPJkUOeCOmLQE+Ok05+7T444+NR41mrvFKCFyiNYWB7EZLGwHzoAtfJeQFhG
bcx9dVINl9FCPHvEsJgOqTbHLWI7yVQDizY2+xBW/XcZZL0EGyr+Uo40p+ryBUJr
pmZZrmE1uJNhASlv0e+KTMvNj/SgG70x2dhcBI5fwZRC3sozALgSUru+6ZAX416y
WA1grGOJQlbHn7fCvsyLpHaznFNjY2m2PF49RzrE6sS3VXip1DcP3/IcfnX05x+S
kTuMt2AeQl5QyWEVlcZ1jxt+EFctExHBiWB6sQHOUmd5CjEW61QDMfHDwL5VTEsV
SZI+QrEYZ/rf6XgMd8jYbZ8GObBrwNITvNhtvEbHUIZ8iJYqm1lqGRG1pS2xWuRg
y3/XoDhjcGc2BCpn2RTv8Uf/wgQHZ1M7UaCj4Cuq+jmir/pYDrniJMg/dqeE9Yqo
3z0EmeOsci5/bUtPS4lfxX2+tYhKS2GdLBJlIYNXytqZqZlZ/+1V9Mqa15ZCai6j
KiZq9cVmfOi6LdN+uSJAgQh8oemRHxRpppTNS4sLxy9feU/yNPzu/2bsQeZH9YPO
eYyMeDsYrhPtntQjjB9JWP8Arxl6jVlTP4ulLTgEu03w8CHV/NvCEjD01Rtu76xc
J9itUiukFt2/1fwhWX69DYJECmT95omnF3Ng/cqxHAOTKDtj2EtTlZEM5lTIUKlZ
QeUma3mzX4OODqsCgMm6D/5OXJehZm1+UUDZ+ieqGChA8QoNyvBEbSo9nux1/qSs
WLFxOQ9xw7Tjw7VwLmVugQEl7IvxDTxVzsMAVoh1cLvIjYX4VtJi3TzBzAiPHJPa
gQxxcAbkXX6icNf0LEM5gt8vX3fUqZ4IR350x5k+OnNYcyEvLiar3pCjEWhJmjPA
02YCvgiT0K6ONkwUgzLmlYzTZCcLcpXt+S6jcPBYxUTFokVd25tXVUBVRzOJuyTu
gdaxsxMnUL464/ySPdfz9wFR/BFATedhUzUYUO8x8k2zdasMMSKBt+6BEQA63bQ5
5pXZxy+c6DTAzsTXxstf0VWyV82k1hX5p33xC5Igiyg1pxMVI5RuueGcrq2EklfF
LsC7JIBKTpRYIJgTgPYyTswlvPrL9aUi6jH49V/CIZJI4a+kvarIAGODYqntKYIZ
ockDS5wEVFoHqsVVs0GyANVwy2+9ZGslQeEH6PzSLf35+Gsm3w1q2yqkz7YfmuKa
IytGweJPZz7gKbBfqnn9P2hqYszCyJk/jbEIBgwmek8yl+R9wRZJR3gRiYffWFnO
Rxr5VONWDttg864fLrM6SsVQg6BvXRtjxZY5i6iJNCpy8RpORjzyCU5w5J6RGSaE
d2rJrXkVf/z/xUm3XgWUNJYVDVFQ6iT8VKf05b5lMOx7rbXWMMFYwsee3n0MzeHc
MHZFlrFUWf34Js4HfwqTu7zgX7pO+0Kaaa9ufntJlalNBFGI8WJtnUJWzTLBPOVC
PfdebzNA+0b1HGV2wF+9pJquW05X7HQ0Uzz5kYJu/HfQxQ9V2P/TlxKkgipk1Fz2
xKta2yXeBqfn72Dq3/HBym2LfkqBcOoLlk2nlSQooP+84DsaeW6ZBJMUDH6ulnoL
MCdSWAWwQv4ucJkDNtk1Ufi3xjBrgRTS/GuSFftPy8EMV4kxGr5I4oOGH9A27e8v
j/ATVI5V5AzJ5TlXSFso1q0yOFSGHrbIDkxyFoYacDlXLOlBo0nHF5zsbW6ydeRa
lTSXadTTSSmRhwyoCNgaA+hstTZTl+bMWVsxkz56ZWBssZTgP7oSqwYRbce5fP5t
ejVJNWgWm81p6mF9TcPs4V7MZl9wEW2VzzAiYCPlSPC6xJ3nv0NMomzUGx9cY7Fn
Pa0zIvkGaze66P+ZYPYJw9mNXc0mC0MTtZEJRW8wM2nDW4bLxSV5T+diddQYxUUJ
AO3pthpO55c1MuL3RQuEMwH2m7wrTWEuR2Znt3OVJw+fokKIylqxk4rvwqkZBy62
UfpiRyT2FAy5ESquWXa4U4WDabER9V5icXd/huCnXuRpTgSi4G35NMUC65lqeiQq
2QG61w+AKKmimCbW2+FsF/uG7O6miEKQvVQeNUwxczTE0RjtLDGhi8/Kn3Gk55e3
WF/UXEsWPoTUk3Ul4J+p12EOqM2G2fXc44nHoJaKh7TysS7rFFWL3FJTs8GqWZwA
cZ/vckh5TvnCJsMCMgeQx/KME1O6D5EQG/ZuikLYtHOV13af0OyNd8d2CQHPVGGF
NVGDp9A4/eoma80REwW/WuWD0JmeMD1mCnApk0opML6waAqE7lhwzWgR4W5zeKJX
pubQOeu7WHQwMG3fPxDozIUqy0evHH1ebbqe1Tgyh5LyfUfis46Nr3hzPNMQS82v
Hie1Op3/NjQ/bfXOEnp1E4rL3glXvryMKT0BgctVGrMPgl6gosx5zErp6Jf3SHGc
ZZ/bi8mRwBriRFB2Ua/ETAQue5HIy06+1XHuxnPzyaAPMHHqHbKZ/htmSj4ybM6i
KHIWfTrVVfrNUOttN8I/N3yLOTBVAGpvNS8yiiy2zm49RsFOGs1vsXmI0BhbOa/t
c1sEJRmbo0t71tS8CwascCi03GtE1MttjYHBqe1cZA4cbJ5e0FkGNPXjrd7yvjwT
C2PmtHfwsnzD4WT4CN3JCLZz5s565afW7r3/MltAuISM8s9nth3hDmubBPT2cxl9
nZadIoOTQQnh9TluM9PHz41LnCj+d/20P5tP/d+hCjG/23we1Uscaqni+TCzNdUH
5qLDHDOi17ObJNTx8HmIsT1E4Uc4YF7ndMA7RPXmPP2wPSIBprc72+0mvbSHidl4
IkQx3IQ1P+M7pEagP6KSPW7tp89UI0EJBuhohcBz0GYh6oYY8p8+MEf7Z/ZDPNVE
7+6tInGZOKpKcI5hm/COlD2m/XPTjYwnwgeF9aAQG8A5H4Ln/4LTS6zg23dtSV01
QdLIF7qIjKDVHiwqdfB1ziZOuedkOsFz232dlNl5izWEnNB4C/NSbwuRmAxhaFrv
r94WP2OR061HG6H6BaOM8yEYrOiQ037A5vLwX4rmcdlypmr86GSutpEomMRsZeJi
WSJXH8qrBLS7nkGRgp0OePiP6Gv6wwjjj8Oq8IA1wARlJ662tpbYSlnjpBrXf7k5
va2aktMpOaE0a9HTjVINm8LFxRbxyufYw7vOF8YeHi2K4OJwflFjkDMqY+Ni8Pzd
hh+3iQyUHequ3wMLLOag7w98IJCo2KJM7TOLG5DwCO1CP0tFqFm9T8ILY9bJNHyc
lYLGmbhqeyUKryV1Ox1UJGSCTqLaSfBAZHStDNq6uwhex+cjQLxW5CjSRizNQBWg
+gplqBNz1hoR6GZw32Vw9vXNCTWBvl/UrWAEHOfs+a1OC+fslpL9+srRPtKg50ro
lQwlrgj+CgZOZVQC05Bbs5NyjDqEdxZo84348GYjuyRERl4ZUPv0IGXUy0qAF6Vh
gEB5Lfw3hB7Dx7IZvpZTVUfVrPoVW0vkLH0p69ZvEkWZTI/7E/Jg8QZjBJ79ApJa
E25GctirOMSuPQuEYnGMC9uHzbbiR48O56LwGS+NcsL6aZIpFpyBqN8w+Iqher+T
OHrBzyqvibxSYNzlqhYKOR3t/YbVrt5HrLT+nMFgKuObNYenbBMxZb2VgZLvmT5u
ZFd8kqHL/NYINC3WM8j2moAgpQKFAcDxcYykDREuwRm9U4f7Dw9LhhkhOmTsVxMh
wiEZMT/rbcvgiC0APTf4pJ6xrio6g+3sW2lK3I8Qy7HwwunOthfuoX+fY4hjbUC7
sODO4xHt0gQFw9r3pQHcTVqRi8LcMseOxyWECg/uaBEPJV1fN/dWqbwagq1Ul9re
SNxGcFB40Bsfeuz4QDBPdlDBwsaQ76J6lHtQYOvTm68V/aszY3dKsQ7t49mL3MJK
DpsPOuydEPJ+FKDpBvZyW/avzNLIpDXDqrelw8LK5x6eKZq5bXgQVwUqLUPUoY9V
syvkPhlaQ5eXXiyJ6s5prj0AWM+FFuJaOsE7TV8qskERzqSRx65udco03EJT/fj4
PjXweKBxOHQV38tqfUU1dnBsxLn1e0qOjvwZCnjRXT2yZyfUa7hVCnyXvIZi6eqd
Q9dRgpSbaUbImzhXJgPrgBNiF8Gz36fENS3v6nztvVesvpcoiYD9PbUplN7o2QIR
bk/clsBAvWqk21MHLsxcP9brG2zMdmE9MKNNZVNTw3QP03qSPK+IkdT8y7Hc/b0n
iVIE/iKNcLhBl1j6J204Sr32CnOrBtrTKyXHOCJBuf8uuGsZlqiiPZCcbkaLPh6k
WKKI9ufFJXF8BvvNnnEIiNEJlXf2mdhvMydbHUkEq+ziwCAtQFaBeqo2Ix1ws9yJ
CYo1SZP6czI6eaIZsXtQzOCyYBB3WjJ2f44nwZ/l06MRfb/hR35EgAqrY1j+o5va
bSXMoYffMfGp7OwIxRpyhQx4S3y/EPtvUlG0jn2mb8H/AZabNRbY0F5HLHf7nQHq
Pr7dr/9NEYa/TlIfQBHek5PyDpK2iNHK+s2SBl8Cs/4lliW+kqb8NE2w3ATEoobE
QxwFaSUDAyWOV6+zKHjXjldKRCefBHkzW+ByNwhJWxIk8JpZWEXJOYUfG4npGYF6
CIyHVi/SiRo+ESgBlHCw8jjzWoo4RCOEtVHk2Xf5eFIoO3NwzgHv5Y3vCwzpahNe
lf8uHpVeebdOUAMekgL8zD8m0vJBeTqD97sdt3jIoXkTC2zXiyQugAtRovwxHTQb
bmY/v7g9aUzaZwg9TfwQi9I2J9Rq+W3z4zl/+Fgs6KTPoaLGWfmFD38NF4/dfGma
kw0l4OCtlSx1fPvTVFnu/Zfvrdy2jw9YYGY5J9CpnENMts5gbU1+GFMQoGt0mZXB
e7EuljO3jmbv4rn0mQyeXQa67wJw8rAPMBHFWxloBWoPwHp3eCmJkXf7Dcki00Rz
M5KA9M7g+RwxtTW/tD3Ze4O49oNfdNwGsZQv2mDduyChwX5J099//oq7i3q4vPK5
PlQC1ORMWwFF9705sOxLcFZTfMwpLabVuvqR7AzmOAMCdbbJiQPKcwsYsETO9m5D
tLEX06/+t+rjFqmO2+0jXR0Ga21QGMeGKVzqK4BhJtXPDvysUyeinSpHrgvIwf4H
pBy36GlYCHvkb7BY1wG/U5zzBmI+EmETgKNKVEUuWKVZz+ebAFYScGykADm/wG7j
uDR88i5nTfHwktgsuJccvTIOPdyE6th/EQ3bZy+2/CyE8sGUojgEPDwnotfSeFRU
yqdkBHDsNL9BJYKwimqQbNy8+tMkMLb7DDB9d+RMwNX+ydqRqn9+uyUrLOhru/5f
PSNdawpd8ML+jxeUOKyUJuGKGNc5ehhWBPH/JuU2742BBLa/iT+PTn0slwHgYHqT
nOIKAdxIjT1M8oFC6RA44Gx5d4nSC8e4UYfArPdAswI2nRbBIhbmB1W55y1v93iF
VgnRRJdubEUQX/MWSFA1AWCrXwTctOhYh/fnVcrd5PMr1ZFR/kaQmU2qok5IUDOp
QBxpDlGKB3AFKXkN32BAbgHt1dTAx0qym/qdx6hfR5rMVlCkK3ZYqpVTLeRfb9zn
7vUEQHZTFCh1VdKwpu5uhIClB5LiFjq5giQfNkGU3R61qbi1dFjw2pecmnzBLSWq
D/BDiO18eks1O9Rx/zRxqcD8aHm57GlccBqm7boyYJErdOq1YVu+CyjbFRdQvb2J
TYIkTKnEoFbf64tVTGihGk3DPSN3xsPWUp2WN/RLk8wGCyUTuhsaeZmmpJYtT/pc
KqVtJMEL6XyIoqVU9grwUQwRBPJwea3NbSPrHo4WO0Tr0gToic0DZpa7XBbFoxFQ
oPFisGUmYhsOpjWdKUQKibPYnEgEkoYWLYMIFnCRm9Q7idY2v9NypRYem4DTk0YB
JPbKceZdygdleK05k0CP1EwL0DpIgHGVYUf/CfjPtsDxTY5j/XcU2pGyVRmTw2lT
PfE9CgvOdbj7Q1Ixr4cTR9X4JgpE80p3Eegoehq0T0dfK/m2qbNmHT+EDD3ex7h7
D+Lu8NiUIXJpJzZoK41bSXXnLynEDNaWKdVRGC25FYQybelGTZpoEwQpxGoaAjLb
xDkoHotw7tfLn2EfjE6GnQMeoiElpm0pKl7VMylcmbCITmmZaCED1p36Fk+zQHgs
WYzcTqsVR0gXVKZdYJsu5KtbAgwMPtH1jJhb+WoPWws001wgxPg5RsKq+EOkvKn0
lfdMh5gQL57RWaAZ6/6fIHDNH06C1nTvaIb3yZuix326OTeWf4IIUfe51q4yM9zl
eqFGkaG7m43D60Aw3LI69IbqzM/WqsdSBEqpC84epgaOsKu2jPpdBDVGEjpniiVg
+nKRetbBpwFhPryOMNni8HTcHtrp/knna2lj0Vcxb9lusau6/2a9+O7FKW9QUwd2
JTTok29rgMs+Z92spSx/2YtWcsMECLJMLWa0ikmxEoh5OyQ7tfsD0UT+ytFWOp9S
t6DkoTTx2ZtGMqyzFTFazWkTyzjTlCXma7tMrkiqm/bW8F/M3ATwD3k4kofwAzRD
AvjrITjaXqVMvBGzpZZ7O/+vt8X8MwCbzSLdvYF+c3dtTCsrET177+3CVF0YPMz6
A2WJkA0+LbeRv/oMI0eB0Rg7n6dufpslYNKqq8R0PfR1kHoBYIE/SQH5xTV5k5GI
90BLmExVpcJ1dVqOIK/kUygpw8cC/6QFu2RDn/YnqyjdY3roWaY58rU1cVwECxKH
qatZNQ9SOkst7TmJzfzbfNuVJWR3CXfkbr8civk7T6+RFCKiM08POs5j0vvH5DEj
FtzE5wx+fUSY/o9CrH/wOsnJDga6W2Fek2VCF03wSEE8M2mRQocqTslZJemp8/dN
cn3EvOlYKCHfXq7wzUHFtVXP5aMFpKCSPogdFBE2FyqEPcl+L86dp4z5eWrZQa77
MUdaPHu1zarBf9VSSH1Y9W0AGYEqALEYJZVE1hC4b+PrdYA+KU/EzQ69qPGvIijk
v7oZYNiRc9NssmiFHyiPzA6SR5LgIv2qHyH78CrO7gidUsIY4wXoO4Fv55K6yOo0
+uSOTvxxhtgWbe1gfw0mmJEzl/h5jtDUlhs4zHbmWyne1ZomFxBQKP2aJrhfhf1W
Az/QOQB6aRBXbbpCYVrA6pvNPLL3hmwLuL1JonVfvraBI+317hat3W2dMzHVcKjO
4LJwdKTTUgjNrjnz1bZFkBchNpHjGKTNcMmnSEHCaWmTSCk46g317Hl85eCI088i
74fVGpOUbbs+6KgObYnVc1ripJWdey1Bc5YuyZ/a+WfG0HrKcDHoG0pbqeUT/IjM
fXllmpVG6EWLp+zGcws1CoTXSbK7l9wALou6uIc9l80bFVpHqDS956LNcYWpP08A
rh5QORGRjgY7R70ZGszN1NTTkFkIQE+7lIGB7XbIVjDHwKZ03nJy8TqtC7+epiq8
PWwXEBp8506m1D0mlj6HK0pQPoPVv55Skjr6K4i29cfTd/aol6OHVX53S7lhCZob
P7ZDVMoqgczhrASH9wanYnEoDaOyvUVk3EuN5ENxILZ1fqsMl8y3hCuHoZsliLLq
HiOq5ELifQclcmJP2XAYuZKC02TiGjmPfEwH1J55EToHVfnOiOcD8+0OQW+Y3hlj
Y1asQPdejKqh1PCl1Jiuxqra2oeGV4PzHdMxMNLyjqeGL2XT95xM0Uht0+J+C07x
6RVnpdWbJNFaJ2kfcb2fKwcXlOO2XC+flN8fwKaAPqdj/lutXNO7SY220GauSS+u
2+0HQiFusJC0hfFzbdqoEbWdrbnukWGc97Fl92HxmWVR5cehSXmdMl5SQ+QxFzRh
Ra938v2ZyFGTW+BuRod6/5jcijLu79ulo3isiykf2DEYF5t18MCoK+nGsjctZeHx
YVxHdWC1tRnEQgcOSXtgrr92MwWjjXpEtQ9AJO3v9SzVdYF1GGvgKTC44xq2+FPT
HtVkbuQbHrfKAkakxahOJIvQW702nb4W8b9jZHpua7LgyKzICCXuAClcO3xXxMrr
1zhS0CbJQp9zv4iIX2BoPny3C+/dfKQEdS0nds72BCs5qCBusbTQ524rUrWRKoIN
57FXKLhDGgS6/rw8JtFvX0DgoNQAOTBtlTf+ZC5CmXJIfGdvT6yZdd+fDs+zVkfa
6skGI76d4MLAAgbob3lBOTknphsYQVGAjx24hSgcpEDTaWSumjKQ4LvL47dSSw4I
6T4Jd4swlc73ZoFb7ilgLLkkuVZs+jrKvM2CT6d8RiKbdYSHIWVXFp8jDTAPPnvS
NO4cucnaMgNNRrgoW5L5PoByANPjuNCCPU2hM4Q+5hRH6/T+FgNw0QHQj2NHvSN1
r6ZGIUG6T5cETQBIybERWRklqmM1MD/D6lU9uGDULOmcPS0MN9tMmFLw42POz/YV
31g99aOkGd+m5ceXeebfm9IyQc8r7bMn/OSwrDyj6v2b8h37b2DV6zyzf1i+BIyM
/vfAdOUDRDMlf0M1tPewPW2KMQc9viItVdx4kAdWLhdGwX8rnPRFC5O996/dkm+4
ptCVn4gABLHmAuRQOc+0rfxoJncaGnLQuyGvcCppMMBt8zYRCAzH7UgDjXvQKp0t
bPmW5qSiGydrPlVUthFKzn6wBXONjuCWd4CprxDxuIuYgWBhaLwZIayWZYgxOkAu
cDZmbjITc8N2Tj/gN/rS1CkO9OeYRv8g6IWWVd/NEL7KvWMfiLDNkv0gVzQL4yme
bvoSMnJZYbJ4VvHBz8/IFg4mam4DTIrB09AcT2cB6S9tamFuCK0bfovmiXQ5KsPn
617mCKbPznotNU631/9BD03Aw735YyKI16ala8vLaC8/IvxHwRTl7VLfGeg95kQu
Uq1v0LcNCM0XMllz1aX+NRLQbfxvTEFmBho4kWWeuLMNf1+4VxFBwLO3gWEFiOYC
ACJI4OzA3IJrYwBEZVE/yRhbhu6FTfMyAJjNIgSTBkyH8kH1CdGfg5Y4SlXCOLUb
ydNAQ244Rvd971Wa70BYv2Ivj7rA0Iyz2yz/lQTZlSd1k4qRNlIPiBO2MxfXXzgv
/m7YtaHfjBpIFHgPXjxQDVwmeEofL7mGSIWY4D9L/zdKMlknI5MdxUe88IIxBrl7
Z2huoafHnr2vgKal8qvblgNMZ2G7D1g9P5Oica98/c9YxaF+xJCAtsbuqtfeldwy
pJlLQHrLjVcOQPmzQhDwhwdFisjel46fxsAkXs6/b6FCnVdeoWKnPYMtp20E48Yg
Fi6a4wmD0jinkoNh0OXsfsdSbceNbLGlanrS3FYfU1L/FdmQYiQqptKkRNIKUF/R
eDO4QcdAoDkEU7fzi1F86qPfzzT3lPYu9A/CLc5lSlFTB9QhX5x+Flt9Ezx2GQ0C
5zwNcE9E597LGiU8qUxZrU6LcWWRgn8AN4IvhEni0AiVas9COmDoKq9fgX4tlXse
KgCaKi+KWDklyxF9y5iYel2Xfm8YuKr14tm+EiHg6eJxpNjx3qnNHlL//zwb7tUw
xjKGxQzh9fG1j7OCLN/8Pa1HV26S01AdrI494mJQlspCkUj1sIV9uLQ6qQPD/RuD
BT9MJwmVIzm67cpO0EjhzLnY/2zW63QTIxIox3W41upaJzDBsr7xYrWVSDv7LuWb
QfXdn5puf3lzVOO86SiW/0vUbZEDNsapMeNkYvXl4ELL1IcUS7bzvwzq+Z5ibbUH
fAPWtg5CmC6CHyqbLsv/W+h5Rk5XvaGAFBeBBf+ToYvr5sQ/IHhWSeeOcIPaRIen
Y4rsFVCVOqqbaccZXXuE+WAXNhgWsY/9BdTzLEogVf54GXiJ0cpiBGIuwWb0DQso
b9E4Z5j8hOxcUU+nvjuMhhHCD6GZeMv2vnVSFj83KB5aft96PWFEuTvhk7SqN8if
sT4TigQIDN64YxTsIrtub2gtRhofxw7CdAMr3vFQkaEHQzCZrsOzJ/McsxVdAPHq
i4avk20FJFUc8kiWqDiqLkZP84bcdd2InstM4MEpv4iNJ0REg9HPVGpcLzSOpNl4
ar/qd33oN7Dxep4P2KZGLgXMx6zmlXcxFcTwmLyuvX62vt15EUHbToL+uvR6asd/
5/RMpJkw234bXWs1iPNv/yW/BVvJ+5zcQ2sSYTa3wTcgiZaeJhOhP2pgI0yI1R3P
DcDwCK7Q76HWmnzK8c8BZxZCgZ3ZPO6NdhUJqORR/VVgawH9f0kYDBnokgxPEp0N
26eQNJPvn+5Zybk4JCfeSz8UsmGIDDBg07vg2qpYU7N0bcW6AMbMW7vvsjthdFQu
yMV5HWJ2JoN1K35bONbN3yD0Gi3gV7+Lq/F38N3NMKW4qiRj0bF2Pd8tg1FRA7gU
Vb4MAIqu7hCJPEdjhPnSDhsae5pTIhirf5XzPY6NTFxCqfWWQvi2luCMB2Bs49aF
CEYU1oi6fwH82W9Hok2cp08DqJ3aL3Lvd2Nt1ePPf0uqDb64RnieFmQ0oHzSKeLz
XRB4EiSoWzQwM1sKKfyGoxL/bZT7eDHDiyQs3IyZdHMlTMAfTLiWdr5bZkVrPIjI
nrjT22Nc7EHwXPNLPw0NmYZ4BYUzlNQVcTzW0Cger0/Xv2ALA/F3Uk/6vf7rDxyW
aP3AWhlCJjg2H2fJTukPs8dDNRsuwxnMx2whHp3DszCkGsBQBo2nxpM+4bCfAoQG
4zyQsM5Uk9eoqLdDT8jXUdpGmbmzwfqMsVsPuwkfgJjnBDO3POF+FuwSROmXmqjE
42qWGKKnQ7JX9k92BmdCYzspuYU4+rbkmq4Wv29RIbgzPgs08/eUztNBky6NPmvo
t8/BrFTgZ6KZVye6sV/Gdt8ZUAxHc5qHQRQgrPa5q5LgcsZZbPcctCS2aiGzbstl
cVAGGRwuThOtfe/GYhyOq3vwT7vh933eBU4NYBX3rZP0hMqJWTPZo2LOpVWIOScO
0G0/azcxR+XCc5g+S5NpxsYKkBkKhLCptKNILeJC0FBXvO0JfzMy+hs7yKefF/qD
P/+7wq/JBzr5252X8VGynsTy2/gRksze+QThf1W/LGYABDL4LTXS5km17ZZnSIbz
rjyoMlF5jB0gbPSZYaMVNJ1HuOJwqyjHIuDOEAAgUru1VtoBAoHWF+/QnsA51PNO
QvaKqfIZuaLb2uptKFLkW95XhRz8Q0PHW3wL4BqefEQDsPX/J/3E5muTCZK4+VCx
XzLrasQ6jf5BpuD/WZr5xS0amiocbtNtVABGulKVf2fZLGeEBIP9ht6ioxy3dInN
yu82+gfG0zfKjtLpn9mbsE7ePOLKq0W3fLgyYx1yaqpF+bzfpcgUT36v8F2iW+ZV
RRw7HvpMdsONeMhUjEv6mphM0E7hrZkwCrQpYf+jYxaAQLAze8NRjGIARyzfivLY
z415NBKjmNv5q1GPGI8jJpG5dJdFbWjgjJZw5l9F6A3wR0d1Z6Iyml5+eVXeSY09
FBncq27zqlhbaw6vdAdXhIkyze2z90SJBW6PouUbpGAryyVaiQIgdLbliO+F/IKa
DQ/idgsKrKy5M3RXj9livR+Q9B0c6BDY7YF/xfif3sZ2BThg+0X0tCCIIlcIzF9i
vTmTHAfJR7qk/WjjFGgIzOckLyAABown48Ruv8DalpKYmCj3W+ravkQWQShlf3Bq
kMqzBM/pr4r+MLi4KnckfR/YBn4wk4j44hTGxgM0MMbDzcsp7piTZ05jZEPkbnIx
3HtqEJxedWEbBmRyEg28cIXJ3VFli8xfU0N481Y6L8cKwxZtjetCdrhUvPzWIj5a
z9x5zdsBi2pjXOl67xmxjMmSGAs3V8yAZfFM9FLnlWXppHLNLfVtIWzX2XNtduCu
v6O9wBoNCxECLmyAWSiHebxpltEKQoqlXkML4NPxocIvEHutpjAiYOF9vlrACR7L
p2PVw7M8SRwfofBUQzgVqYYvBjIyVMvthPSLyLWGA4jZRdxAESxv/v6X7WdNXO5M
+gepA4nE+PZt4aFX/wXm2UhfqUf0lS28SBejhpgOpTFwCBA7DfhQUlgy0AvsZwNI
g29WW2ueAKWWyDooWSdv3v0V64t9dVngfV0ANzo1xCcKXgqjfjwXkGGvc4WRahrj
IS1nbph/oO7nxhd23fjwT495okuDpl5A81ztoCVNTidqYct1yu8DE+z1sfbC+BQJ
BzqO6kqH+s/5C65v/99ks/704k/k4MjtNxUk+e0Xdh0Bag4sxYlPSmiRrIpMoyg7
wfRlQCR9qeL4BEYv5/q85YBZNT0zjUSoKsCFTcdDXUApqWgw85FIA9qc4+HkB1os
6FKRp7cFPE2oDwy5QKXwcREXzTzhxTK/BSGf+PqzzSdDnSd5eZGPRDPJMtACcv2w
h+Rr6LfXoF1NDfquZ6eHhM52lxpwxCOy3SqT5lZSpvHfMCDW8F89nsZD5jE3JSTm
mtCahcK3DA17hnFQ9TUW5d3HhVQAVNFH7jsy2GVCheoVr+C1sb+6TvdAnr+VUTLe
ETBH+gPpQoQRU+yaRQkNSvK6G3X88fzee6xXNxGpc0yasVVMAqSc2DysAPEwcllY
YiiUvmrTqNtB+WE9ZfiEOcBJAPTON6ZbU5EmI1EErtRvncD03Jb+qzZ0xfb0eqEB
a444hbQEL4X094YOtZ5/RtqM4hSwvpvy5UafDZsxnVzIRJKvDJHCq0F4sS7uAEim
KNp3HjKojL1aPd/K0Fnl3/ek6rJFiYyAGfPcIkKCShss+BSuARz95hudAYiRtxOK
tF4z+J8Lnrkcej0CX1VuTb1ScLonEqYWNDOnwTKRqxPwmCoQc1tyLt2R517dkzVF
yhh/i+M5y+Z0VGowycO51zWvLeLlaKx0QrE7UluWbuxUGHoLtX76zdGoFOEovWDi
gwnrqKF92rcX4gg83MV64rEKiM4jy4npUSnuDgQZaOXGXfge6mGq1ha+h5WmsZGH
WVkYrUzAebOT+5tGL2pzp7TfESgP/b+8GlSSDSnFdu1VKQbXgv7q9A8bNEbb2n1+
YdgnUL/1ZYgrhwHmQQQxsJ0A1xPUpe8QJDaE4g6+xldVBksZnKPHPb6snYbNFY3a
YeKDmKNmc2WVOAxOZrf3bKeTGbcJk5JXbJwdQW43u2Zi/1a06ubtr/1T3GbS9Hyv
0fR3lq7zqIGzt0eI5ii5wDDwGBl6okUwdJCaXIFCPH2yELwLc0oJ/4oYX03SviiY
hx1lLRDSTyW0SccW28wNfE0MdEJAyPGigPXN9rQwX2AhDQ9idcJqXI65aGc63+fA
ggibn4M2esSRxrMJnbZ8RwDCEx3hdwF1bFdwRkcog0bbizaanxUQnSj4eYF8oCay
iuzQ9d8UTWoFwzMeg0SIveUmvJ8Lsv4/Yr+20ZCkrrCkZTK9tja+WmY8TSgfjpMX
9+fGN5Yd9vGtoGEhhel9aUjsehbAyXZfIMjg7CijIAc12Gz37H4Tvqw5hy40ygpA
APdLNeQwmi5KSxHXDikPpNf04RjN2Z6UGa3JjS6FserNT4auc1CgROYMt8mxfi/P
3k9OSgM6cygT8O7eITSrer7bVHf0eJiBOiLQ72iFtuyd0f8mPeCAxvJu3AWmKpSu
l+lEoaZCp909mkWIRamybCDHGfLv1qnLlEGbDZVeIakSKp/iyCMHpNHAtkrRxykq
vcj8bAE0Mh1WHnk02MU60Bf/lE8uc9TBD1BWb9/h8ehmBuJsNePMrff8tBy4cyzW
HWOY1KcWirXWRJkQyjPC3GyEuohgpf+QpqcjBnC/gAHybn/TY3tIiOCU5Su7yI8e
T2Zfrm2oZF3ZzPvBdfAnR/jvpdzTkXUPzBfwjbe43eFm1Vyts1BD9U6RBt0doWGk
5t8zlIHwJM0OrPBpDQ5Us1KdC1gPrXsKIiyg4JTS00CQ6HQr6HeCl3ohviAyusBT
2qaF7r8VkiEJtcuvEwJtGZFdDISFRKNLyptcT4A0lxyOw2K/Vk2bKBc/FCiW9Xj+
o4rkMv0U3vrSOq0vs6ZVF93H+xQaVyI8+HE3hIZDGsNzGVCDpYUfdlSEGP6dOomK
UdYLVdVcL11/cSIshGL7L7FiGEtlTRtgdLKMXrNwA5k/sGIcTdPSd3Mns6c0bJ23
h+xQVoui9vdh0hUGwYvpaV130H++eB20cJJotLsQq7bWELE56kNIHRgRfLJjeVaW
mpoOeD9Ql5vqamqHL9AYCs5xGuoJk/t52ihffNzNx5V5FpQYlWlAlJEGmbLvgCMK
e/aOpPgVfz4m5QLmIb7IHmXX4ogKjHbSFKtTz41fyFjXTJ112qv8FULVERAaWIbX
MA+w1VdltXTdBHNK9nx8wGcNnoXjo1TMXF4HSn0AX4yTzn09WGwVDwW1CjayrhLZ
lofpr/JPJfUwk3WWrZuOOjrj6yjRfCTOc+/OdogPkU2s6LegQ2GGlmZNQIJ8N4m2
AjYvWCL+EOfiTkX1fBctxAcWq2uOJjvK+mMcwxajyJNIRKvGppsI4w/EXpGoDkNh
0P2gnbAZu8qhgXoxa0bvf9zi8kL36PaojLVp+6/JzFigfuwR1bUJ/dwqDhBFoUOx
NIiWohihlJ+sayPzWv1/EBZa9U9CvOiCv1UA/+JjjBHhzRi+3J6XV3cNmyuU+quF
KCiVTv4nh2Vbbz1QDdIe5/xaNndDF4XOzrkUN3m3V6nzQKmgLf7KCMdxu3Z6QSAy
qPPzwFWRStBJOCxuiQ53xyrp5bXEFhb6naXCwN3hs0kCpltKqnWbhNvMD8/kpcv1
SjW4Kd91DtqMJ5OBmWbHkmnamiBD1dnST9r5SjyMmItERMyREt6c2z/sF4a3PCss
F+fZPSjZhZUXkFJqnYhD5VBT7xgJ5w64erp34oT9VVeuGWSmxRRNiZwGJpmehOPx
5GQG11JToh8v1Ptgvaa57oB40LZ4uUwXRrovtNB7eEL2sUSekEw6E4Ynsojldskq
y/mKVF8oi6FGATv48fwwIN9CtaaoayRo19fI4eKWGcIadcH+QQMtEDpQfbAaXlnr
rKFg90buf79Lai0NXg0p8LVCGTiAkzD0iMYrs2Z9un8RvJ+Q07DsVSfLBCbk9ELE
BfSw+iEKFFZBAt43PbcFwRe2t5vo2kBn0evzjgfEiH4FeC+S/ABqPR13v5dZf6xR
sO8oz5oQwb4UeKAmHgeh0rRlxdkAe08FnBm3dk/dbm+TcCAGu7HkXeiWQ4CyZMuP
7jS0Si5hILZOi8q7mu7B3iXAI47TuaZyE7lEVmPRNTcQzhGhJinkvUuxHdebVxEw
Ig49buKC+H+/Y7asWn1GSHC90bZqKpQ91nOeBHSR9hjbDtM8WizGP/jJPsp4f4h0
EWyKzfJsGbytp4NOGaYMqFLQhuZbi629KemMLlKBb5iwzoXTlvLZ1hYSaqAXvhvM
rNgw2UHnXCq1XAbSJTGVdSbs2tV/Xec9HETlc1t7LFTAt/m/mvjxbuBleujbYwW/
LjGoTuKJaxc0w36zYBOBZK/VLce/fQe0SXgkGMSD7gPdKKUcHyU+ehQqB6E8HE4P
VXYhqaFE4Pb/wUfV5eY4srGPFyHBHfySy5oh/QPydPw4iQy1PI91bbEZEOIp8cV+
DGvq/WaXQY04CuzRLcIitpWBt+qIJlKTqRLkUqElzY654BLzUgxnNA3Krb1ilEG4
kQb5g05KIcCcm94cVruop1/zPg+xyqRXVDeGIhFbNwwwle/ZGY9026wG0H4GSxlT
uhheXBSgXkN2zlLa4T47K8UlQuibp16n0xN3q1HshpjtJTmts5xLuv8Ol3GEy0VY
Z56DS7NaPrfJAe8pjAvi4WFiWSc2TCT0zyzD+/5H+FvchwoLrYdENizG+W92x3Vm
H3E2nd1xMFfIgjgxIaJOhzprUetJ9H/ZAhOyaw7YKZ9ioReLoWFHgAvpNhdPZ9WC
8XIhpgfDjTp3yqJdWMW3keiaXIr7ikyKzbtUsMU2CFD3jfutncmDRAHwVA/wRYtS
0wr73sS5vrnogl4LMwV4JoCyoPgxhcGwqFpBc8azjCHIapFeMj9ek5tLEkDzPM0g
DYmUNS+a/zSuudGilx1z5OAl+2EDP3R4LZhzeFR30ev5iW7QGSHOkTmRQGfOjlYE
qt4EQPl6nqgPKx/GmNvXbK/w5tL1Rfu8S9vVASZIXrPRqh8Ez/NpyzQcmxomn+rJ
MxeJu99/32cGS+sZaVMVocy7ZST78/NDKGIvN1fOYWe8GpwjY6wDrxz2EEbW8ejB
YT+c7B3lQ5flizUK4gxJhTHqsWhBj4Nx9QDaAKSaWwO/LBS8svZRPF96M9q1VMxd
OXLY+mJoq70OoB6wxIcskKID9yHmxe70upt1sWgn06VkGYF+7kHKoWcjjrWwXSx6
GPOiebRT4m2729cY6gwwoG86rLG4vtMmdZ3HdqSgckg4KkpRjZ+8HkzKK1iVF7p7
J32UnzmAgjlLrMRIFYRdb/hZvotzyaM2KI0tPGNwuiukXOarlyRCJHWRV/eXcN4p
VQmiGMdkEzeNn4X5lpRJIHwbySmvJc4cNLhtsEhCO8U7xsYVkn9B/0Al9wtZmW7A
hofiCCvBOyPRh7JAgZzAY9rxVcFF/CVD4YS/bg0UfNJtT5YGBYk1GMwVId4TW+uz
cPMPcDEMo8OoT6oHc1+Bj5oHtRpsFrUVRZnVr8+1NVvNGvsZuv45jSG0eUnfQhdT
RYgajreygkxg6BSq4PPY0dQW47fhQfgF6AYcPJIZVUmggsDD3yAW0cGiuUkjFqy6
CLWmZHX05H6CzOrWysPsHT3VuwURuNylWndIk/qlaPfDkPlVuaqAkoilqWRuDoqv
t4ZTMDT2fEU2Y3aMi3Wp1hsbSNkdw4Sn+IeEqBJ+Prprrkq5IGce4WBSkQETMLXi
Tf2zUh4L9uR9e6a1Fy5hS2aiK2Mc3gpXi+Xo2Ogwfzy65F0A9d7gVAoCj1MKt1eF
APgwD6hEEiZ51B7EdAS5TN5wkUxWjywjAG3zINoDCo7yfsaJjARKbMOEQr/4/OfQ
WPBxJx1KtCO8saDdS+Mimnvos80/8Rqz6tC+1XspMCccQ/MWJJ4btNBFu6QT9aLE
Cxct68dQx+I4P5r7TvG2kzpzD+yjzM6qZmnDHUqnoT40N3RhOaC0eNGUbuLAHLD2
8uW4GEVGnWhgCP2Bix1FuEf1JeFbGR4hB88yQIa4w54JlRh9Jz3udMLS9Rokt5Ev
sXvs5zgBc3CaqBkfES7O4+bGijHMe2TCYqx+Yk7hHMpgU/9N0shFHTE6LI0HSMdY
9kcdbSaYy2bPmsUqruY5X7aBsbKDEkew3vAtZmv8qcSzAPJL5MbaLNvbHrLt2UPI
H0rgaplQxk+XfEOnQcEUQBYih8ab+QMR9JywPHyo+dU+RUDiDgk52+F4a/V+lKUQ
pzNMOaR84lcRMAe8GAb7l9TIVTeqJmj7h7JFEa7j49rYPgYbZ+jJaGthORqkYjh8
nJWS2jEzp65yQ33i2A9ZJ3jpAIlg9M/QKpiAvSaxf82b4n08bm9npxzlMoCRTapD
ERvEm3Vc+OU+bujF5yHkBf1k9ov2Fwao8z0x+EPt0IcbfugQz+HDaul6+GJC5T6J
W3C5TyZ8Fxc3/wiPYAT/fvfzEsmsTMhUsKtFUPCfYeCx6ymLEnfBF6E8CCGpwJ3Q
WVnUing6Jhu2d7W+UcPgX3saxK6L850OHrCM1Tjb2P57Bon4AugWIhvxCepB0SYY
Tb29njwNTR6oqotRh9gZGVWlINEyrtvVe5RODsP0vuSyLRQvFibYESZ4+4u68eld
UdUyjjTepLDCISE9g7K4u5NSNy3bZRw+TkcyFgGFmNPnAhv59xn5mte7OQ3uxH4y
BOBYfORB2jm3M3CuX7GKG7XoehaU3eOL7U1e6NCr71/VJnqdGZ7aYqPX2n6UrB66
RX728LiO3egVxoF7XR1HBBJdGd5YjenNnaa15tNlY1VsnTz7qJQxkVJ+0vun6OMJ
5NVH/8VaMzvdNzyq4FDt1hCiosvcCGEORUN5NpcxR3FoairivE04nmN8TfGCETOM
Xml6ddKxZKrMSO2gZ5zzOHXLPpQfXZn2qVnpc3rTvssVn5IuQMtlLShku/Z7uYEO
0RUmHIxoPca+uX/tcfYwO1s6b3zGa1ZlyeE9RSsjhAWSRysqvZd3jyYO7IuVbgbu
UHP/cRz0c2zGMhGKsk9O7UJ2+wvlimPkpetVos4v6ibAxgJB3m48m/lboqcimMQj
+04zYGyke4UJhZW0mxSkZCvsblfyjVpjRB+KgfR7LDTTs0j2xV6qSTJyuFccFpcK
WIbjC+zhu1UFkDgOvd8hOtAGHW3RKeG9ktq6ENDEDKV59A/4q9RFchq/qKKsmxM+
ah5ZVCDtIpxjZ55WLr1Iey03X/ATH5mX7MD/RE8u/FcMy0jwjnUXLf3AnrSgHKx1
wgK69hWYekZJzJvUeHFPW7meZV93HG0SeQjWWGzOUu1RdZbO6AcfyRaDyEZhPshQ
wp784zty7P6KghpyaqviZcr7HXFGuZQWWMZ57gLfZUEpcO+92qM9D0hBIGrr3KDg
rl2mLoLf8p/10f1sZ21F+AWTh2Y0RDaM0jJQlYSGkiEn09G1cHnRjvKOTqZfsE0W
11m15db7UXll47jcFnBbSpn77dcObb0rBTfgtEjoUKl2drXrHchtngFEtf/qIN9t
vgieMquE37AgFodzkEMqXwq1NeEn6gz7Hs8tKoe//MBIe9Muu6kzzGgYaWxawWtV
noMC2Z9ROJ2M4C368mCibDPuHLEHX5O+dkRw5tiwmrCnhwlunWuSEulhKgKh3RbG
Fb7afyG9PpOPjJszGHNKPFERmxvNevCx85lsONGjufozb+F0q9/9WXnbhknbKV8K
13kyreW2XAqsUly4uatCWN9bAYPf3ZEga/ObJVfhtoHP8wJ0Jb0A3cT2xXsNIG0m
dxa8FecmGagZyk9007JmCMSIpBgt6nmuEO4N5bf4PMi1WZvnaT+XjCBj9o59mLY1
HMjU6Me/xn3P4oIQBd7Y2WFlXburpMX2Xt5z9ZM97p2Rx/YqkqfsaXEkvhwn//N/
QDaBbJGQaQxQlbRqyrSN6kCbzY3PL5ZCwDhaUPJmEyERFO6ebE+DUGGPChu2RB4s
VHg3FS4s+tb/aO0BvOjNBASgDffNgEtMB4N2m1zCpJwQoScD9ARzuru9xAHH6T5A
mF1V7X9gTjF4VJgU9XFBCuyAEkR3zQ4/MO5cN3oVq3jDxBty6FQYsRoI1rqBZ8Ju
A4o5iMaI1fwR2hHZX1g8wCmOnsFUM75hixBk6KaQ/RquaAyU015wgxdFEO3LiHBC
C0b24V1oxMqntdKLvuA3QTmwH6vozqIuWt2i/1OLI22w67OUF3x8X92orKAcjWLx
MhBkKB/n/mSyqIXwrPvGxv5P3Hi2Y6qRx+/ciyJTD8Qb6S3SmgVr6Tbm3vu8OD5L
2GyZ8tirGhjP0y02hlNyBYyVYfIhZqcJuVW+w0j9PDbna5QyBaBNfmlC0SSK0T6Z
Mh1RMit13u42G1Atp8oCNzYLruksNt1mCqiCSdQ0quKHOoyjzkrXNDMkIB+b8fhk
OG1HE1y5lxD1zw9WgX9qWbSDqLfPQ/9Q0XJgyBHdElIuBgnCLEQAg7w7XdrOkBwU
7TgjykC1n+ETQYwK2U3BQy5cS/1mfzRyR5AHnYsUr0re/aPMpDHCo26wGfavy+fR
AwYs13MxMRdSzuVBOP+J6Ev8L8O4L/gCW8kerPBwcOybKkWGl1N99c5tnv+LcxJ3
8U3X2yqZQlmPXGuCeXpSuYIWHkqdHJSABxRpG8neormT08k5gHrgpuEZaEak+hl3
ZYvhQNXdlhXa10Snc86eCH4d6OiL7esUWP1VksMGmRlUruWWVVo8MGDuEu1+Ch24
/ZqbnCQs5FDxEa9JBJjTegBtoH+fxNSmEVvnQA33ehRZg1ZKKx6hErfMha13WDSd
YY8mQ+hxoOWLEpG7uJf+XAGyfQqm++WOuieXHKKkxtyZc0NzLzaYdfmZ+yr6XldW
3NXWbGRxHSzqJrZC2hFyueV1F/WgcnA/L0QWIVItvttlSywtSqfnaELrSbIBpImV
MgV2JrDj0zXwxCSP6MWcOTTGURuBRsXQl4i9h7dQFLj3zQmr3YZ92+qtoI/tG64G
Wo5ksFbrcxDLIzf2Ryxbyy/rTuNs1rbYRxMBEDIHcYDatG6ZULjEMecSr33USq4W
dGAFlMyA6KO++7kYddGnzhj8/syyFaXSQA21ENNulOpb/aBdLGOuXL68PlkMI18c
cktOJNXAKMzPrL0Q76yq0Qc9g7rrZtyJ52veGK/2KAiUhoSgzUQTZZr4tOSyiFNV
pwE8Z2pjgCeeABtYnC7gr/7TlZzdkrgMohZdp6iQRyKDu2yg2/kFw2NlHR81cAuP
xE0b9XTJCrJs4NcqFclABBpczixPnw4B/L2YBDao4ODlA3UGUMIEJb1LE8Iz00q9
AaPQzH5cp38fOVA/Sh9oe+SJ0OUXn6PDsuEUUue5KrxR6r28Lbe+Jp9tr5EE+Q99
IOKJJTcfeM9DW0fjKvIKN0PbtH6sgSXciUvgRn2brdvtNqRnBbAt40mhKUFlroWV
5+/JKdF2Lr6Fce59KhjXsi6DbtX4NkcWf2/cn9L1jcvMEa8DBnu/PJy70428ia9e
Jdsjvhgso0gymDtI65emHGdaWHjfeV102Vyq+S3voDERZ2NGlORs9kSnTLpKQRGA
yHwplCKkyohu8eTr7+ycOIL/4QYw/L/J9JP6uxwcCTH2+09wornWjo5euwWTUtFp
smHvBZiysT2kd0H+uFCl/Gi/30iNuzQoMNMUZHQj/EmtFl4XLgcXNNSPbJdr3W6C
1YfyBvvF3t3Uu07hsLGOSmeOfR5NcPDokD8y4I2IQPr8tQ0BITWWLaJCTQHyIY5J
6MHkqc47l1+1RRIz/USNpua+okALrbnw0+3y1Gzah7BNeJXZwqZMVcpzJMTULS4S
LMp9JYpBeOpPaaabfrD2f1GAXZkvYjA/CVUtHcaWgWR+cLzKC8DDuKzjyeszPGWO
YR1o4zBhvWgzA3q5dks5HyIwve2/F/JKgwFU97LAD/3S3sJg/bib70gio0iZ/nrb
sPU1XEhvojYYmTKZgj0KI5uhmjGla4R3u9n42g5V4XQ=
`protect END_PROTECTED
