`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I+sqtS3nTLCrOFfaWKQCF5yjM59Gx01Vl9LzyR/8H4dv7zth+GE8Tq+pQlroJV6q
fxNJl5vqBVTwo3wYohSuuSk+MOv+fK3w78BM0XqTrLitUG4DxY4Uom9Eo2Yv8Hkv
YX1ARd8o8tUzPhx9mNpodANHekdOY7Z/Nz/HpUxfHvcM0wscATrtOcbTR5pPOZjK
Slr27GMwU5iCXdW8DrVcAK/a0Kh0+ONd4P1S9ih8w95a3Slp0gpV7aOC+NN5oUFK
RjQpPKq+b/gD2LT1H6nrmkzAUf/nAJ846QZk7fbZXtIvedxrxU/qFX5Cj8uYvWRc
QYzVp+4JnfZN9oIu5de3EEYxLfqhzCTgYFfpbYKuJ9Vwwf/3SCXlRni1WJerdbLE
BkLnu2q9nQ284FwWJ+Y74EAm49YLALET/r4HogdyE7Rph9gb+VGOApudOt3HIw9f
olGotDrN1bwLBuPB5p1yigPkQplfjzWTWrq/CXbz+n9g7nZCaknRAXFpTK6u5n30
wkuV3B5FRPq2CdL9Fu0OqsoHG7UInnlGY3e9e1TPswEIGw7h8RwheHPLJPaRn36i
72SOJgNevb8fqox99xPT8SNmsRae3tLZIEIFp8Bjse/XXIk0pILMVXyy+zOCvpxB
iT/LqTcyRloh+Kb4bp94SX+gxP43dVGBx0/GG6FHb+YNg5Uil32eElypyPu9srZ7
VAnZITbiJ1WOYfyYRJGe20+Pce8RD8cId8GfW44CwJdhyxRGFEFW5JDym+fM6s10
NCYeJSDyYzwPX8CvKcU3P3CVg0BzUGqch+uyy/vq5fJ/i7JRHfdpOf2vjHkeT8GG
EA9gpMxcgBE72AXa+SqHzxxcPHRHFtteQzbMIFdur7hKd4F6HirpiQlldSrbRSt7
uk0oN3GAm0t37pmEHs3wBU0hGAm5WZfGC+CzUmNSxTAS1+chxbYPvuX0gw5+2DaN
R/VBmxj3ne1Kys5Zu8bdnIkjmZJTcT5CRQFO7QMuAKmwu7OohC2FJy0mlVh2Qcyh
yd6Xy4HOLEK9eMvz9OlF7GEDQs54yWLZPAGZcwAPRe7jknP6ZMgfi039qQIRuY+V
bGqlDtGOu4ngq9oBTU652+1DmFouOkV0SJi2IB7rDy6Ean/2m5GcbVabfAmjAsMd
lFAQQf3KPTavCtmOmk4z/i/eW7Civ5LR/ErSGSJVBDXHCNXM1C+lcqdzc36xtz/V
4mi992HOOJpfRqJ4rLzY5V5bvWpSD+JMemDOp9uibvH/Gw5KGmtWVC3FZcF+umRC
X2DsUQGt94shV/u6HsPm6w5EppLytrRP8onqk7RgGgcuATtOh4nP8oIalZiBTpB6
GeD0ZX26V4Hz2G/dDk76UnVVzmLjOSPpdcgGgMqEvYI8aXe/gEiCm6cl02z/64K/
gxda8oSxjciy29Hx8gBRkwmXiFuQW+quHUPJRBemE7cTa8cGCduYuDS+sH/f0coc
T4nCYRP4yHizN0LKKodOqcIn4Doe4oXpCAn6/ZXYwCHNOo5StJEONFWDpGpR2d2d
La8b2FZignW169CWdQ8h9hP09ildiic8Lfnmw9XkILd9CRk9fyFXpVndOEyTZTwN
RMJLmuU3g8usVyymI80iw8UWo2FMRwdwt8gOpcRwj4Jv/BeA8KlJ6M2CORaRyEKx
JYYNHOIVwjJuIEntmXBguror/gyUIrj2rBkKAa2ubXNX99lZr7XEp3lM0XTVxdYS
v5UH/MKUegdNzFUqw9Qew4u3a+kFJhlcKpNj9FnJcs0Glp/hZ8GJ4cc267p57TIj
Q/bHSOvlvgd1PD0Ttpxl6aQ5RudOvQKI99TAIsOtk07C/DdbIpbLstM7yUBh3SBv
qLJzo6HotPwH41+zlBefjWgz3rmw0Kg50Km2X4vKYcfM24ZUiPcRQMszjAWpHbhJ
H0jnu6ubyGbwgX9VpcNejlVQmMQ+5+m6wbl420FqmMT9yiC6/L+Z6N18j7JSD+bi
ChG9KR1bvPnFZr6pL5k8qRgStLUhd3CYIMg+D1s2yZJ8gLFKyl4ZdDcJq3zTC/ry
7kgPitS7Onfnb4Yf7ATZpQUOLPIJ3Sx4Ppcgs8tfQ+7st+ugeZa65ITXO7LoWBNU
wqfSNPUM71vZuT4TwBVUurM888OA+xvNoOJe1DgyardH4rRdwlZ4kaylXABg/KCO
LxGvYgYXkQN3qtVQp3fNLH+5DiIvNj0UHbegGgsmukl0bfieEazeWwa5AEoi9wBu
sSGJh9TJFQOXmQuO7Ne1jUQv+cfAJjNinEHVGU8H0GRdchtcObQhIPDzFK14ze5q
hL16+eqF0NBYMF5/ycoQzCxLSV6eHEm9zbU8/0WaGbTH58ivQigpYfNdXJ95QAK/
8RDez/mGWKwu6NGWq9HmXHACRzrcHnbT/Mgh2WDFu6kiDtrW7/mD03ai17x3vdhf
FF+iDrokgUcQq9KI/uaR4mRdzr4xB1PgNmo8+ovgD7YVc//1iEc8nJtY5zRJcg+f
/LzlryWJ7U/kmZMDpH6wZWn8dmzpKgpAjsx2FGBJW1nsy276vDk8dia5snIG6uts
nVPpoVwSAjyDAJ6bEenflLJvcJ92QmzKavn8LgFSEB6QusauKUNsABcDmVs5Y9nY
BQgeAlFHjukwrlG75VjlJZt5IQuQczIBy+8Sm9tp+1C8fDGmyq2zJ4/9mBheA7bX
voQLopuz0KirAnP6m0ABu8NEpJBwXnq1XPHxs9p4AauPHes9FXfa4WJH7xTPaOu9
tpx52K/XuIsdvQQ4y13eiKRrAEO8UTZuo9NHf2l/YcH8T72TTz+Ip2hNP4EHL561
Z0LZ+mi+OGo3YPDPGq1BJmCN50EneDzSwcL6LVOTHwjk9dHv3NJKiiP+Iv5KyvJT
KXI5ZALYa8oRZ8SCebk3FEnrIETeunO8vWlJ3yNCg0SDhBlLmMA6ZhyJqaW+kUBo
1Y3Wi4phhzweHYELMGnvRLWJUdT0jztvJxOQb9VtLxc5yKwPq1ZoFko5cURYku+2
OcB2n4TGlW7DB7J4CsDDwIlCtLnXM+r/E7ARvOGqZL7xQ+w5pecYBpw99DTGHle9
z/w/OCCezjg4LOXvbqtZ5w==
`protect END_PROTECTED
