`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFx/g1xWUC5W2CFobZquswrcDEJwFUYhdGQDeC+q8/5sDZCIU542AJeCkQUq6XFi
Gbf9OxtTYCek+Fd4lffgjZUsvM1L0ZUYDzV4SwaS+bG4GSk58AO6/bREQpNlvF+t
wRSzu4eEmGbLiwMGyR9Ct924ZYEvARmfwdksc/+PlF7ouRLofmm8GGQwO6QIxt+i
wZyk1PD0coyhOkY8DbX3nP0y7SbpVwMAmZr7zraF6m7qfuJ3ZEGwkj+tcOXust6K
fjwb/gQN2lz3RbHjD9oockrsz1/lXemBq4G+5i9JkMdfRiaQ3VsEsNKBo8AP6W4t
wPHzvsIAqO5MVq+W2NJfUl6jJa1b7K4rZABP012WVUpsTNygmAMHBJnJhsUIjY6M
KZA807jLTsCY4AizuCyF8nBS1YTtunoRpfRqOuxIwPdLQZx0GKFMTkoG3kAJhwvg
dflYvifPmJ7lQ7lGYGCMyoMvvSkoHaNPuNVoN7lHsjRrrI52oxTuj3qL7p+1A62E
RZhg+94a9WpcfuNBSj17jkIaKEXy295RuRsCQeaSh5FPqL1SlNc7OmdgeSp6qSU2
m6vpzLP6lpfO8w/5Pfd6Qmi5D1Q9wKpJNB7uVjnlrRHstitkNecH4ZIZ5yzAceJG
OE9ivuvdmkIhX7+xnbahtw==
`protect END_PROTECTED
