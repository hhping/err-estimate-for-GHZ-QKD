`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oD/FCsAUOFKBNecp3xDbbZAhhpW40+Z0QR+a9puvXJjGgJ7nEU1X/5Qab/FP4Kbb
JPa0twWrbrQ+yuXcVTJh0jKB8G004ZRDKLTKpI2TD3UrH5aaZwqzSxfxoIkMspLq
qUKEPqw7c7QzZDwyWPD03XK2d0fdSvJ2xcvimxKZJ/ssG26X53vTUqUmJ7K/X8ig
UMce2oDt91v3q0GYFaVxw7K+eApU+YEdY2TLPQ7w0GvCLI4gIWP4Qvqo7C50WfW6
UkUjYjOJd4MTTM4TBR/xv9ucZS5wni93czd1TkOJEDWo9t8+Eq4+mibqdbp0GJ/M
8ZNuAG476buPmG8btWKdXKf36pbGuigbPRgDYByEeBFZbWBAqrLxaQDGpOerZaFr
yVn1iFd6kvf9qi8FN5CQUx/xtsufKKF75ma1fDmU4vh6OWgimTbh8/G1GXTHXVR3
K+L6z2J01I+lP/zQg8dfwCA0tu2D/Zdgv9BhIXNMNkYlLyISYThWs+WpQG0SpPQh
moX7ZB/LVXg6ShZ0xOMEENTq1CuwBSQWOIMt+Ae4T7ktUN3O59xnvV32Vh1xvaOa
aSxaQPcChboj8fMnk6baB87zbBb6xmma3Dko/WviaLcDJrojj/S4KnvPgLg7vpcw
KhohUguU1hbQ5gL2MCrmicE1SVvZYLZ6BXGMpUlHc2+IlrT98n5IDex4+ZPb0D18
30PuJ+b/hhPEn8XGYrMnrUkexdMMKGgBWwmb+GoG/lmx/taTZ+obaTEmAT3FVIPD
qNh0YL68jGmSbRmOlVQA6AXHaiJwe6y6v7f3bLVjhWieWU1s9SRxd3imFXrW46w+
rH0tbaAlheiAAcvNO7nnneeQtPaKlyFMj/0PuWCsC9FmXGjN5+ZhiheaB9/goTE7
HVZK8paUPjUraaiKXyRtB7XYyXo17oXdC/anpNp5erFQlWeK2ElBApJoaNjcv53t
lZqwlaFa4xEfJXRqDKmYBxqcEpmDWIiOmbczOBcPISfRZMrwzySU0SJUPw3Dfyak
4ni8dmVlei7M0rBGiPe9P3QNopVZABzV1N2lfxQP/dUI9yCuOK6KaFLhR2HN74f0
c06/i+sGX7X93H3FxIZPl4HmRw0BFP9dQr+4CcDqJmPWxEU0KzXZq2TUt0BuPBIn
WEGGnS7Liu0g+kjdUVS46m3V5Y79687Dgj0ec9YPTSuuzfPoEdc96WN2qAeAEEeS
BSs9Hf7tIt8VGjNZq5dSpIrLf8F6xqhRbF0zi3n2DHw=
`protect END_PROTECTED
