`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKNTyqVwfGZVvV4Nyvn33z5/AR3SrMOeJHts/RXG9jlZzfjO/Hk9luoSUT4MSR3M
K5f2hKJ/0vVM83nBclxn4Vm8bSK3bHNZ0C/8Zn4irVDpeCPtvx9FSRjZg+ATn2ca
jDFTJlzcHxhp1e7xka6m3mJdqSrA4pqTlhy8xiIshjMJjPuATH2m3zTyWt+hnS79
PfplyQVTFfUsEspuymORkGz9tepaPS/aRvUqHpQQ6Xra1SdbHygIez0X/JJPNLuh
vEUFJgKXISDnSFdFGAyjHZJXGX7rFkxBwMLw7/k6WIPJZm23WEicfVTbVDKgH5Ui
mzHTXld9cdXC82yH0suUPliO8I/U/RjZ7CrEiBWzsjAMm04IR/3tZoqDam84hzW5
bz5it4BqhiTBlglrUXjG2NAOm1cwnioqsRpKhoJP4q5QHmcb1YeC8VFHkTuKMThO
5FyrLDFpRRtgK5A/4In1T0GnNBag8QXxiNAYHCisetqlsArFRA0PC84JKhKisXRK
PQ6eBhsSMvH9DlKC+bWWoigBiVcmZeUz0BMNKxMDYbQXIdEqCeuKYcooC5nu6s4l
97J7DgICNXSzomTIMOoAjrrwXhd6kfRexxlTwNUazRvEot0ehIxrQ5CLNC0xiwKk
+61bE0L222jjUrDc00hl1T7SWFuv1tJJJ9+u5BYJtyEc+JWUVHmDeOQgFODIvJKS
`protect END_PROTECTED
