`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gatqAkX7V2HWyxRDQP27b8BgHYdElxpzwK1f7gebeEBazL/WxIDCZT8QV8kJ/dnR
aur6MG7A+CnZfkwFtbz5dBU6sAOlRNL7BMgIVlRjTaQjtkZjgZ/ceFdZ1sKSMIeW
TxuW+J2ERz4lSDubu1p5cS+lBQsAVcXGqRLlgYwJrpt29IZ5UYzOOPoDQTI4s5/5
qdxrjd55nleg4v58Rt4doi8euI2BxZ8inHsKkuJY7hI/kcFpHc/AFJvBcLQRbftc
xy9Vg6QA6ThyeAVL7qNXqST1/SmPwfXLXWf7/fbtpApEctP7fxY7nBVS4+PvQGG2
Sf4HSfh/RuVIWd3FXxpdvPY44xTqlqQxamD4d6ZevalQ+Ks+m+b2fVdCxU+4TbpD
RsVxIpombJR9z6p7QDP1vaPRpEzGlF2HP+jGgCIv1PfFMW4SDLYNB8CG8CiuVcCD
hWVvBuJwmDp+njL2r+L+Npls9ikGdknyaclZgzCBiRHIPqhsauaxaONDdAO3sPJ0
V7NhPQ/TwUsI+vWSJ2N/Nd4I9VKL4vfalX9u64uAXiac6bYlgKN8C5rUDAvWyb5l
/LitFdtUgyxUjwnUBDOp6/scjBY2j0jYuXAGrw03l+gQToXOvKKffDK9ByKa8/zV
4PrebFUIKwS+wTaDIajHbBFzGDoy0oVGCKcAsLbQ1oTuLKgeppGUIqkJw+OWxYUP
GkFFzFaEN2G+HkoeJW7do5Q5h8OhRKKGe2C5KU55O2U2sPDzzWWioSlyMSS1M4YU
req+wXGFDllX+5DsKl8tViEMl+sEoAYAsNm5ueIpcSd5+rxLuELpTeDIvaZRFvD+
6Yas0/DJQ0rL8VaRSx/BttZiSybwjdravAQ+E2eyUmoxPGZprhJyRHTTZQTiFMW7
7B5h+vtSDGJNfB7ISCF6ych5i7w7/nBYDNWJ8vhzzH8hCH906qCIl72A2GGAId2T
74sJJHDmcEt2N9IrXORkFACiHJDd+x9lfRnGKZC3f4JOMy8ixHj26PW/zUwcVaES
z35rR8ISh9UiBt3zkUjhzMN2LZCdmDZUbqjKifqkTFeOSKJWSV8C6Cidxao5KGYe
qqW/puWaKtLHVJR6lPgyRKgfAwGYOSUT0d3QCfumAg7IDYVMjEpfp4NfiBt007E6
el1LSK3Zli1xqqBCwf1m+jV1P/4GcBJDxG6DRui0osc7ujE10f3NL947yt9D+++H
W/v6bHcQt262jV2J3Hx/uwsCpsL63zbHR2Sjn0zklbQ=
`protect END_PROTECTED
