`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AXcnwa707hBXYs/WsyJeTOtIy+K30g4Zv7BTDmyAtwsEKt02B7tIJt/0XXEQ/oeI
exIrTusgiCtCnhG8XbBwUtByyDlTM+3MmsgN+jNWAjfwp8UA3ROq+KZz0OlNIPQ2
QWooWccvy/7S+sQTEYO9GBbBICqBkLI65zgFx5vAQJuz8wiHFQcqUHH4UvXU7BTV
UvUr14Po4ZCjlvqbwNbRK4Wqr1vrfG0hVr5nka/9DcTvywbdlFc+qliNLzS7Nhry
7DrzVQ1ZdXxa5b6cnNSe6ho5XpKvFd92JQUb8LdvjewY+DWHdmp7IBjP/MQzz3Yc
JuTLCy9tkAXja7I84DVcm8W8ivHdkgVQXIMP1r1z5dyQfD+cBxtAdrTGJ8mVOEPM
VejBY4tRSBMv7euH7eWd7C2uKZYTFGnacBuBRpe8s8dP0VGNvi0PtKHKSR2qaNgL
bb97xe1LJNNWUETbk+GcwXo+nWzCEfVDagJUZNDWMHnfUOFp+BdKyq01Yhfi5jgf
BvwBcEYDFzdrMn/s8zs5EvPf2DtEYmxu+Lr8zXrfaLvUy/+nEVqjwMOBMz7OceS2
4kA5Sqnb1HgOH/F38vLFW9EK0lBSv8sX6aMbOKL3V9sNZ9Xqytq44nMIUccNL8hB
/IlayP0yYyPzzVCAV6SP16bDBj1NcAT9qMTR4l/zuX0XhB8KbyG37EjS4aYtP7mG
cCoBo69wshazx2qtdHQoFsnOggkA5H5oYKXOSJyo+euhatXjV1Ck3I6AjWoD8Gzv
+0vHnXF+taZd+ZHCBN8wAnwFOgm3EgJ5sUfLhFnbXTyfITk2JpFZBDG0M3chKr2X
I+d+LVxg5A0JcOBgWcH6hHfrFyd4yzJMeRvzDP5bNVG84sBxq0sMo0xbWWfS42M8
tuqnZ2vJ+7+Ff49CO4IJqBdj4+9Rhb43jp2rLUFocBrjYuC1hygqD/gx452SRVmt
l0DMPrDYWH0gPI1qLj4Kv/LB9PBsWGlUqFmLeWwJXiVbgpg9iDvDo3CQJk8GjP5J
GiKSQ+3PVHan1EkbWEk14PLZD89KcsXa+b3FcJkYZtrGnd5fFStbrnL6OW7AxbYX
2X/KMDfWfSJD4PrSLOSH6cz+zlH3FmluTWjlf5mWOft0h8BtTclVE2+Y/QsX3cNZ
tmkZCmQFHNHjmwmwomj4t+/tDnhVfRKe8MBej/qsC1YaGnaGhffcLz0al4CdqikU
FzTiGoBH0C68lRClpckOsg8qac79H92x+zcYJXE8j/9t00x7vGUrlN2BnyebGGgo
gK6V93s3/s6j/UY9puX4ENVAo9hTIWRqxb7NMlV9spR7mlee0+9ydvsrDh08lSE0
ayXrfG1+gG/0TX9b/U9aQJ+p6uSRNAmUoonq5vBt/p6xCgvihZcTxmeqXvmsoeQt
dY/MhXbXPG4xYxsqh7ZoC2n8N4iK/+eqqFLbxwe32ZAdw5IsO4JTgmg7BfiJUTrg
2Gbjpe+3f8jG31UvK51S2nh18dBWVcfIyryucj4POTiCoKE1+hOAfzRkbfAFvt99
l+tS2FCSePv85QEJw81CIHdiVYngprvgMSqSY+qlJeuPP+T60KJbXciAPU+wIU6+
oDZLtNc8ri3vWKKkKm/4+yGIeecm45GPzHSeQ+rG2n9lJF/96ccchXRpk1VV/wKL
nG0aJURG4vWZQmmNnQC4JSAS7/qCDGce3gRssIScHavVrB+QSlMGveKPiyHorBhu
7HkHcny2L0g/IQhUj/MFKuso8X8TFPi4oiN+5RRG2v5uWKeg7ubV7C9I1N0GBtZH
zre9hvBSqCALkCvdsqO5s61TarEIaHh/l178X9/seciHA5ppf+c1SZXfz9yuBCoz
1CPEzIhxxNL7g6CKUjFrR9vhhgHMV2RZufgoKmDld0j9+xr64qZq6x2BdoCWut5d
47fFZrbWLWibHY/l2QnZRxTBrH+pzO3FBYSXzVeAisOCbfPpdPzu4Dlz61p5UR6c
loYl8IpHrLJ1reMzj3tLTleGm8sZW0pCoUpf4+ujpnxBOI2jnFjaG7teQBtPjbj0
AidEGyIdSw+iWk9fDln87XkC6E7hBZOt+snCUqGJtG9rjECE5UeKd0xvLFC/oRiK
L3MunxvRM5eumOVLnCkR93zwHJnhQh5ns6jE2wEXOj+Xf5irEMbRS4yk3hA2q0yM
xJ7nobVTz0Yzc0vD2RQQtypnNJGM+eGCktwGUJq1dvd1V60OYS8/IXvC5F+LWE88
YzH19wYVZL1rXHKMPh8qSav6jYlbhFP12t8/XPbabvTiigk8kBPK/CNmJBpSeAdS
jSDRdnDisMqmAAQLtsuv/OKvsYAUBHGegYp0fs0zjdBaQni9TTGP8ODjiIwmplPg
GrzhS6hoydXa+qQoDeQaFodzh4to6dJ2gsnpcMxS5Q3ODpg847SsjLB4YA+Pf5Lf
lOVzdGcxEQvRsPuE5Fk669TX7Gp49lTxKTNDL8icyix3Sv592RUDY5cYN7NM9KC5
1Jr2/vCe3cRDP5Pte9/YAQi6k0iryzz543h3+iKwmgtIHuN/D0qWk934BhZrZqJQ
j7d0tLjtZwcbKKxpp3OCobr/Ox50NJMkghcvW96byHBagssGCULCOdR1S5FBymoT
Hv0PzQP3PVQmsGkoOIj2jWI8poFLAqyEesW5BzgmfKZ0Aj1+Siao19KgNss8Z8cI
fCPQQHKnrmmsAPf5jPlcTXunoQKwnUlA5iLe4aewIEYPuBuvXxqpekvUdagU0ylK
ZIbV7ecl/YMKxcS4KYw5ZzT6izGSlQQrljXx8lq4pigf9gPtIiJmLrSdrYCJALde
9ZJGeCT5nc135BuIzkmLsEnaZY5lTktUIa+/vQJ/5pl7tK4woROsoydxQU2y5QRO
hk1um6wn30N3gq3D2ZMbnF4CkInmZ5tfJ6gQQbtvp1EEH5z7Fi+vI3KznO7YrTeC
IBiddqkSoF5gL7cAcrmIldwUqtMJPUnD13tuwGvSTpSZji8plcbVdvxOi/AFR6EG
45M2LhpUyPQvrM5yStDY5NKBmWJhLOUqH1STOZRVYErr6WhEu6s76sPfvqgp60ez
ZEcgH100pUCf86q5Na0VIghq1xkJujHqp3Xa5/UnGNt1GhUj2a9As8OlTA9vb5c/
TQNw9r7WouCzniINCWMTK/Of46K7kmIoqQUCt08VAnITX5CtzR+y2EkQtDezozZ7
dKTRUzHL0F153YdbeWnVfhgfA9kC1dNuXMwAXCzVsd99yuVuTMYwEq82rvzEYuei
bCgRMi+ZktLjRoOFfPvy6JRIIJ0hY6eoDl8tPGb8TYOdAX8ie66R+9COWaiYoShs
5i7cHdihBwUtX4RhUdnXr8IQD+cAFMewujnkLO4C1OHKZkrHuf7kGzOsarZMEZfH
J5ujYVw/UzM2f8gbpsrWRozdsZyLr1cG3Z1jbGVNTgR1iNwNA1eZHKTtT5YdUklO
3kjH4SuP+xuYl9+I44MWSMUBagPUDZ1ZZfivAb9wl2siCpyH5rggvyPS/jQxtfOd
fLDscUOKrvi+kSl+Xe7sf77UtmtQyfddstI+X+jUbXhQWjGJF1YFKEVl3kmWugqp
k7zBChIEaJ+h/SfvCauP7QtJ0emRGwu5z+sTi3LIDXEmhjnuO+ynSMGyWkgD3cJo
X3CdQab9Kg5+b+S6IeBuAD9BVRPVmKFdvPLgqFgsBPDfc3J1eeQBSOyHTBnzzCOS
TgAJDvIXbCDe0o4SAdlvabROTR776uEKHcMGRB+t0YkO4cU2vJNQqm7hkpZsesgu
OTZ4YjiePl64izQykp0zse+5mJBkLSyA46T+aWfzBolqiUFdLRYtzOhjuhrqrNpT
iLHO4ErMg56qLx9/cTUr/e/+AAd6Mz4WUUAa5GEfo6Me+6Q3UfOCobpPhl2t1oLQ
LzJ+chyPiSs1fbRZbUmXl6Gc4HXImQqu33suH3UVx9NcLciZ0eD1NoolYfDeXpmS
qTLt9C1Uojp0tkASWixyi+jXqeBX0ktckYKqeOf1nYFPVDPDpTykSEScgp3PvbxU
CjPiU2Ev1DGtxbq+/fGk57nVuYb6AEoa0AgBp4DNheWJenXmysmjDu0V4SKghAZh
g/AZCmvNR0eRqdTJNL4cNmbtkxQIsO6l8lB8rGqopfDgafzzoyTZVbAaGJjyX8rP
Vu3mlwBVFj+MkjLSJ0HKCj1qN6qePzkpdUgAboeHDz6uEsmkBHkABhNkfB9yjvfp
umYmkL1nM/vkoQBDjJecijUlkrAIU9Hs+11BwNBIAa2kHeP8SErbO24rg4G4OL23
Re+ZkIIW/PXyFTvCqBvFw/ZunFg6C680og3tX5NW0Vz7XsBGwF6f+tQs+zcpPgWi
zP7Yd5wVAspdic+pG3k12ybLdQlN2O9bMi33qwijOjA2zRpFZoiHBlp8DolSIkoJ
17VP1URDJ1+8aWQD4cLa/SC2MdNG+FqfE+XsSaV2aDIHxhkA/2e4z9J4QwCZvvhJ
onzpMLgYtF4lQYCryTEKTvdqRM1uiBkWnF572D/lR5FK3XkBUOTiNaHm9LVjTqHM
haZMXE3glLcqgOTGJ9jDCxtCcTcomhsTjNlREnkhtO1NEtxJKh//g+VWXTvrM3I1
iX9eYZsDT6r3LnrttIxx2SDafng3X1ATlVkaSFM24yNCJXOzm7uCyYaTs7FV7yBt
0ZgSVlGSir4r6mYTkZn30k3dftDJFtmu4Q1rvY3tNJiLIUXVEu4fBV9nkL4Nm0Kw
Igs5N1zHJdOs5DpDqgy3cyXvU1csBkJv790ci1G8zrTJjprK3HB7MwDUhyWAh1N+
Tkjv9xRHrABCPAv2sD/KoEMUWXVdV1Po2iZ3hEzOa6k7rtQL5CjZjVk7FLTFkqzn
EG4lXaKJjgY1GWRyimi7EyR2/CYSZxN80F3HPloXUAnKHq0BpAeNDJDGOzL7pxTk
gDSw17BxltrnvaszDIHJbs2VoY5Yeb7F9oOSQLEolY0c3hEUMgOj66PBKzs+EYCK
xxD7lXDjzPzuCvVY3YvfrScWhkGqnULNmTTn3H5RUTVabyqYV8IYHeByIBs1dspb
Q8CqkGm/JL9WW0ibNu3VRlq5d07iKNlZ2V793ZIXufL9F2Ft9fvwW+e2lGeELBIP
5F8jQ0gz0gOxeWjwsfZ0QtV1Gwk2CraVzC1XpU/+HSfuS4awpzL8IUYE0cK5rV8I
m6csGszibIxprb15BKcoaLHUUQHZWyMFrcl9IeC2VCYBhuCxOWlpQeqkkgxbXCZB
gXW19PNtb6K8XzPDXMumhTdoNwLt6Vs6DVKYwVu+cRTqdbmCcBAbAaqbvatXgnwv
ddegfiU4YHPcPM6Qa+1leF9d8HbAu85kdXlUV5negnoGgHcItbCbomQOWV9wblN/
wKY+qSQE+c+WfK/EawK2BH7ShkKXuE9qBO4mqKRthsgMnld56zpTwHZaI4TTf7ma
YbuZXDKUnSk9S4JFdDbOlBEcDFM+8oOBxgFlN87GeIl9YpinEb/qmPGpuFYHNst5
CvOYYemOoZTNr5uAOaeYTwUunHquEetGOYvDtP0NuyyvzcqcTbi/fBigGFya8SxV
wSwp02i3iOxNAN+q3+7wNg13qGnoAWEE/rW8av6iG+vnrDwD6bysZ8tHUOSI+1jc
8r9Cx4GzhvCNJYB1sqqIF0Tj9bl2R5G2dK2Uws6WIqwIRdOEq6ekYM06pItr3wyJ
KQO1+T0TZDo2UO+5tbhXllO6gb1nGqQsoSiSwkvrf7JFevmKnp+y4h6OxiztCRD/
gGAOtIOkWdYFXlxQL4Qsc2srJwj9/qbZhO0ugaDCZoOu2XnUU0SqgoT8Q8t5TWd7
1AGPS6jsEchi/25SqWItH73repQMiezD8oJs9n+1aHa0w/TucqowM1SNsTP1bW2V
uA74PIAMMxhzbLq9afgkWISarZb9WM/znfo9gYC17RkzH3S6AIe4q+RmKw3TWt5y
d28e98kQI/FGfG2lYJsnQrFMJy3yZ4Wapw7ZqRmp3Z/Eklud5iaea5Tldtq5eICA
VGyiiZ76m1fM3gIh0LAmhpGVlrqaVaWjfYOfD86A2g732XslGTiFNJTwuEhdvLEz
kt1fdH+UvRhsOyJvyJTTD+R7t3hRhvFqv/jqNjguSRzHuLDoMIvyLAkbZjSVo0g8
v8Pn95LYl1PfpBje/YPLaJtB+MPshnIAqiZPCMgVjW7G0Dai449CSYHCHd2cmxCo
t54cpr1ovXCjJ4sXtbyBbSgRfj9dgNVvwNLOIaDpd9sIstWcJm2eLK82xywPDFRD
5LcyJ5h+OevaaUfmWRsrSiAgXvZ4lvC7QfRhCXp+I8+ELHbmKG+PcskXxcU511lB
jVuOJHIhMF66CRbeyGNaeCc48970EsEZOt45qH4ai+ykwlLn3i3yxjX4kr/5eRQN
j6aU8VOa96tsY3+rZwBYuZF7ECqM2g+DKpS89KnDSPa4brv8W8v/2KrJz7ud6ycd
va7q/oaktbj41Oqc6EDkvhCbVmNjjd+2WBxuiMPLrQBQNrOtpbR+6lZ2qOf5YY2A
J5/Su9LoS48HzfyNqr2xHJS0Bq7D/sX0uJCoaFq26qI/qVuoUuOee8LK6Y8NG6Iy
Py1tAhTSXpOYstaQhB6rlNwwpOmhcU2VtD+ibuzN9Yq+MPt1uPg29W575RWem8h/
7QmVvU1J0i715RiBwLwlyuK/KZY0mZ5sIPdNEGqzI0ypuuFnl3gtXInLN3fgzG9l
+i02VF4UM2ankuWwOWMSUGVsemPC3JwDC7s/kKso3IuTvjKjC5jVwjdRN27aMQ9r
yw9w1sz5gRR4kmn72pQeiWpdwG3RPdjXTS4bWyK2AZgKORg65Hjsm6QJ9PX/VRCw
eU3v+/uBRIbM6ZCfR25OMLrLGLRWHr8VFjndDfQDbApJxsnWfE1YiRFD6tT06pJk
QxiAMBWFvtRdSpgvm0C+4lxUyNCWo8r4sM4VvCYJ01kyky1FuRibjTPUqwTbrDaM
yd0zKPoXAVeIgQerclfuLqHhkgUntT8Qrd/HwpO92ux6u07zjQvRHjUaMHQmonLu
zrGJyc9wh8zkKtNkVrUs8GrvksHliAuLBurcOqda0VNJOOhuuGCbrxafJf/mg6kK
4gb6ZecakYXoBVIkMpgsVyXBFpw9qfk7IwDerVzYHSf1lU7RJkyrkZtyVO/jX7QN
Bus5mW9SgE1BPFbxxrXLOiE2iQZAMlosoSNg/6JlLef8v4tzct9RWuUhVOm2QBrE
yvAhpB3h+oasqLjt29RnpudRrvPNaq3hEdfWsoLEdEdH+uSxc/udS3zB0IDXRBAx
UiK1V7MGGy0ZK4PO6zxYUxOTO7ijGtBPptQlqy+Y82cNRyJFrbB3mxbMR4pUloej
vgI3M5mesMA4MCxHro8dHemrE43zJkWfmtDeHsv65UESBSnTGLST+gRAH8XtbqCO
CeUf05drxDm7y4iYBEdM4qaXHpJ1R3FvoNymQuJzFgif9+ekK3LwWjpgwWgkpzjU
NZv/u6bLXRTPdl/SL2tq6UQYu7/kEHVgOzVs8vqTCUW7OEAB86rQ5ifsVftHq60p
gr+Abs6cHtkJZsh5Vj1ADrOPQ5TFZ79H+xd8VQudaFMbSU43MJ6nmBNy8sEtQ4uJ
bX0hZo6k+Col0v64ZYPdv1m8nfyUnl375gRBj8q2wXUE9AW+sKJr//3Ze/Ipji+I
ix5AuwOwoWzVSCIopezgqwNN8SgYTFIuIUSvWBnrroYSMNsRX1e5aK+PhGnzjsfh
a2hblILghqsHCgWroFwJnLcs50l5iMNf5DCeyKVtrRPXye5mOHfMHorvn55V4VHp
hG1u7ZAzHCJWCTBEjguuYVl4Fgtd67xNdACMIf5Q12NIXD4CFxbkSC2AFOI0QxPy
0NkNVzacX2Ov0BryHDUj1BReRfbf5JK8iehdNw06x4w65NfP5rC/Sjn5V+FzkTan
mkn0gEHDWvAWKnxAETO63M9gtuTmGZh//UBkkV9eVKZEpa1Q+NdHE1fiTe3w29HL
ehm1rEJ8tOSz5dw4pQ0CtuNHWEfOeempEmOgfQMGBDkTUw5ERGeUJ9ip8epVr8Hx
OFW02nfzAR7RLgNdsOwVxr579BVJVAglytw4HATWrphgYFWBA+9erGhM20M0sEkD
+CauIEcWkSXjFj3/07jVa2jVhfWAB2VxIHV29hLlIENXdM/4zYnQhb8x2xTGdEor
OmTDDeMU1M+seeavNE0KvEGe53A7LjMi2DyOfIMEl+23Gt4Wkx9pINv6I4Zbwve6
zh7+/EC29kikP0j7SEWcequQI3ybEtY5q8xG9F85/REZnwl3JeUV6aUKaq/ABjlE
oER9sALZbGUoCiQ9e25T7emRiciflXc/WfnEM1zEcxnrI29Yh1ddsLz/RAxwjswD
9BI1XHyQmtta8LUHkNRgU4VDSb1mQWRgMeUkTGhx+0yjDwnv2rGnJMSZcLbLpNGy
qhNKyJLc1xlwaC6BqBzfywQjYurw0QCHyDHYftqOD2nf1l34gMzEVc9ymqBPrDKP
TiZVqNUdMK2out4ObzmA6BpaM0RjDtaFkI4aTLfsCLWF9CRh1nDtIBl6tiEm9Zcs
WeQ7PbCtsAdi/DlQZ0NT3XtF6qSVh5VXWB6lY93hziuQPOD2v+TWCwTe9g0HKNnC
DKw/gI9mu48IsAOLyaDvHoIKHUK2WdVCVbtNkRuXZpXi2v1fy2uunuARJeCPpta6
NLamAWU+ic6mNPic5PQa2TPwtIDMTVAlZTzvZqe9yyl+rnT89iQ/2Pou1bLyZIOh
uya0HlpkptSARokmVIwAcuYKSOEcNxX/hC1CW4+ab2pC9KGKoO+NtuqK8zK5YNOE
TFdHwOWzSuLBFdZcFrHNUQBjcXn/8YjCjS6pOA0s4s2J0nC1o+K4alrM3J2zrJQx
DgU0/RhE/ajOnHpUPsBJ0pljquMG53zdM0ul2QSynfqeAskuDmX2BE4Uj5ZcNmym
10+awqUzq0q9bPCvFTuClu6teLoIaANamg9Cb3QW58uXH4YGYoOkugkYw4sr+N7C
Vm7clfRe8FRDeJCIc6TbPM+hKwTviIS3zSbnVwe0tGAAtAI4WRGu5LTIo3wwQpuh
vSb/8S22oYn4QLYf8ko8IT4Q/zEVCRdSYLAW+xxRzdtxcQ42CYcqzeD4ByVT1S/Q
CD7QE8dBAa6bp5hkJA6KhoT9tVHyWns6Y6z4k7/uDtEJZZwG67Ziac+Iu27ELIhL
L5eXjyHhjTzRycpqrGQ8faxg1EE1326FCsZWE6GQvbePCnPBkK1U1+K2zf33ZrMz
7Hx44Yg5Z8VCdTu1tBRX9z2l5FFZk8uEGAzV+Mvcbp8LVEX74nK28aRckjPn1i5o
8s5/FbUk3wNongqkyo4l843gwiRd8n+S2s8e+DOpqyDA6CYDZJ1Rd5YuSpFNZ9cG
sl2XPrGYHxyGa5OQEZm/3rFNk5b3wq8yzpH6+GIMGG8P7JZxx5NQ9jQ5U6ZrGWfr
IbS5S5UuCQfF0c6UC3CFxYS4bCrF0bItRoqO7EnL5KWzrJ3yx9ZlMXRp6B8OZYBJ
P+ZBofcZdI4RspuJZqLdjVfvLmTei86G86zgYck4XGRUkNSQGLJKltRg4aCqQ3ay
Zdhc/PhXgxdhJcbWrWianI2LxksYzx9y/gIE/fi1wPF8gdJEoe3DIvxwkenCmqxh
ZeDZzLEd2D9Odfme+YR9OklP4KdbVvAX+KY2LuydMhUFrTa6t32/Yu1oHPliPyV7
WlHA1C8QU4pSSU4UpduwRhAQo0CUJf3qHmb0+Mc+VsseNNpX3PFjmQZN+dqEDumV
3e9gEtWVRZj/gixGreMTdrYMFcixPwsJltyvSeftl11kLJqPwIVnFGIlc8xt9gVP
ujVArqEXKgu0+7YzPFmIe2Ps7LSEg0u4jI8hBeRsjxFN1NxGju34heiXWnRl37fo
PSe2xasogQwf4lN6RcI5w1VgPdpHOqvMUhJWkl+XwItEGyUBtfT25fpChKxqT+h6
CGDBVB8hzpXKr3F5QWvL9QQLwHhcshNsQlf6EwVabZZQmR0lJwI+V4X7SVxdRVJz
F4iyb8mRmDdIq2Wu4iwxY0J8vSzCIegd/PrQnFaSyt64tOHCom4kR4mWOJji7gyc
AOa90RqQhex6kl6ZNkK+vO6ce4z840iHOhtN4k4lIBVN3/9+2QG7LsaM/pwGzqYy
bQOqPQ3E6NvJLAQodi2SBrUwl0C24I3292k6zB3UB4IwknQvcAmOVkr9sG8W03+s
JhdiWtFz/pc+soxC+Ow5Zrw5go+1yVruyV6IQk7pI5Y0rUkuVoY2py1VpC/sYKhs
1Mm/tDJTL6J7zTpJkJzboR6dqkxlXk4dtzQ8AWH343JPIyaS2h7Ci441Rw/RS4eP
R17TZMjGVL7ocLnRV5a0CKMN5wZhTsQNB1+vgoaFN7tqAGeiAVI3+0grJchbuypi
usDRwwFrApONMtTCqLXuB86lHdyBZu9WjsQ5Gkk6mQVOnOmliDBCeyZY5G7u1rZd
Fp1ZV56cpaDjoJ+f6WXz8R9gD2uYJD8vVuz/iIqdzvPqyVQ7G2kNBoYU6ZewQYfV
y/1nx1JAsnsk36g5SsEqur2hAMmSU5+MJJuwkTlTbk2ED3aHFubOkmsTqtRn1zeQ
FKbSFqmUygSdUi0armR7IbteyFZP9nTwfBBEfjKmTsPMfHEZ3gdK7ZUR+jo+/H2c
/swaxfF4+mUTxwabQDCCADAoiJKoePwGf3giPdDsviNmsZJG5mDPhq2CXONrpSD9
3fGgD6XxDLsrNb8J4dheHW/BIlL29tdqBb4LNjdJUjhmKJNXFrQipZ4CXNTHUjfB
UbKlAovOWAUKECbq58eof++5srlDnQEYRRyGkSOZfUtlUdcUYGgDosdq2hOanMnb
TeyudJwgFO6ZH64OAoUMcnMdVcEDFf0Xx7AIX4L22KSQqYZcml3YH22zu3kSWklb
a0zdjmpkB2WucLSYO4fuqJwh5C7LHS9S491RJFLqMHw9ZA3FBXp3NbT6ge82G32R
/pHNUnt3bxDvqBzSixi3NzVzLLqMViU3Z4eyIl3/9W1dO8cyVb2o8mb7DPRjqqPB
7sXYgSOezf58i9WItUSTx+tTR2zR2hnCy3d8RLi5fAV+eep3kwl7tQwEC5bU2N0N
2Alt/TnKLCVukPBWU6DIZE+62HbFkiGiE5SCcjsZYaTOWwnOX9UMSnO7cdLc0EEC
lE+cuFoLDZlBbfiaIr6HC9bcDkXvIFxJoF1Y+PA1z4EXFI0DjJ2x2CawY6eqpYXz
e/jO1rvsBZ4jkYiBWed8qNfWsuWREBRsc8YeGth0WH2O1dypcZ+e4l17CHGmGFox
wKygC8WbU/K7m70XPDkdzEeGsEyFe1yXHOptLnlTwxzncyjlBcL/aj/AKCRRk9pi
GFtRe/gOn+bnwqj19utLmlP2LHOMZOzEh8eIWyMUhYxFeFvtHNBe8UXWzwdmZFSk
hSXCschoinlPg2c1h0d7cNy2/cxPmAE2UBVNBBKNyuke0Koljy+X24dc9cPtMZfM
PekpQfST0BoK3s7qDcnXcsybW5FLxwgptV9lvZ2KKNYAl5kcDtiRn7+EJohYwqwP
FS+gx8Ib46Vdd6OWXExYJK4TfUeWRGFjLkVb+0E5j1/TmL+EwVwgwnSVNs4yJ8+Q
QJcEwodzl4O9Hfywj/iIv/emUrhhhb25EJqtSaf9JMlQi8OfUjMfsK5mmQYjinMd
EM/BQp3OEWo68bCyDlMlgmiJqe5Vrx3pYI9geEloydDnHkRwyeUJzqaAHAsXJcNk
UefJpSh35Ca3p7+WPXnaiHZqa56cbecu3gLOVdm/cCrA6sNQrU+FH+Isi/fy8jYf
aFCMv2Gut5vNp4XycotpPME7A2+vQEcBzmoqNyuzwj+ZB+dtFRKq9mhJdg0MXqX2
sGl+qbmvSTk0mn+SLbhDhnEbVzPDX6pg8IZ9kWwRiGzMu3UeOvzsWxHOA8gtwak3
AAGFL3NUbVn86sjFRNQzwOMVatYj8o5zrnWng8ETy4uzY2SsgY7VkPziFWS+wfDP
vj+0m+umSnvYaiIAr+MLREu33D2WF65nQTeL2ArZXCYUd327jd/U28Nul2NF1jon
v5e5AISQVOBhXv7mWXabIJYmHPK/3NPRCIDTrC5mvRMKFMoUq8cd6H/6HmhDqtkE
epXSlCca//bcEP5oFoDt0a9gjHeN3YQ66RAWeBBo/uh5bzW9+b5y79LJ+HPpQCFv
DLN8ASaK8WVmBZqMQV6nkEMQ6oAgDVKD8kDrW+uDza03iLPC7fGr2sFK8Y2VcTwh
6bNtUvpBT6Mj489xW/rsw/oaIvK0TE6692cDk6LGcOkkQp73uzgQwGmzwtSYKGU4
3VIAzGVncQybrxtxg4TjRManAe+2bRQq9rDka47vMF02tpRELfzvR/NJalyazFBh
qqK1yvxUqwQF8JrpqcW4q6XElhRGpIf6Zg1YdS7WZ4LUUvn0iZSaoa+qzujvwSxP
rU2AP6FtNldI524Jj8GRvOH+cVlkKALhp2WFUdYCfVgPUojX79S7PbsKDAqA5B5p
9klijf2fJZZDbH1PgsmbY7JBibCTCEDGw+rQlWqi2o/GKWNtnOn+p4OUXk7R1oHB
AtxN+kKJP+JfvGmWqTeHM5I0IzbnJYV9EN6Oods6zIZHW/J3NBcHgA+ULa6mK+BD
JV0s9hgL2r9UpemPwUqNuQcWvYgEmweGqY4/Qw3Jw5acQzrToCXZtXC7cS0eMi+k
Va9TUV6Zr2LD/6YcdV5BKZRK2NZO9Xl5nE4JBkxggCawaaCX6F9ipPrgZIL4CwaQ
y1AgEYE+T54S+eekJV9AiGR2x3ZgZFoPtWAKnIBJgykzgLQsCsjjYyzZGqYNjOkU
pHACz4wkN0I2N9gp8LWR8+0NlbK/sf+OG2lvB7JMh0BvTUXViOX+9VFCgeWCrytJ
UpOe5kHg2Ppci2qatfivJt1UEzf2id50N+h7QQ+lIagL9wmfs9390czBE1cROc2Z
nkOygD526XjlmBXL1OCPysvGixR05qyB/15AbcEE7eRrhYNo1Kqrm3Ju6DOlQXKt
TgldIyBVyulOWrh6vyl0VVpxEXFzRtQOq6MambRdagT5UXf8+uiVyIWQoj49LKL7
LC3ou02Yx/LsR7rlbXPnnQxqqQjMgARfsSc1Jj4/zrW5uh4O3+vwtSheWE8IcSrJ
GQcLXGDjwP4IeTOxyjrQCt+PBh1+1IhKcUNPoqxN4sWBrsFpvPRahfkQaHP8SgaF
C8VVxBEreGg2ibIFjP1xyiGEr82aLB9VJ3umBh/XiJyAf2TC3czEEb04O/3+/Zzr
XVeZnEnVlKqQvSOJ+/17o2KaU8F2YglERStKi2eRWKLKYqY765Hf3mf1IqbVbA6u
g5PERKWNc7bsWDH2cdS62bd4jjMmZWnAv4moU+zmoM0u/AoaaKhuNCZOq18hXHCc
RYu24AwKYqdT7NLlBWCSccN611FD0EBqeyIN3rpvYctoiy8/nsx5rAcCziOu8NNw
lyxDzZpirSEPyx9zTNAawzvB0A77OqJmd15ndgRx6NAw0e4NpZGQrTXi30udLkrk
cgSfnYwey7DagGr/uSfHOHPf4UULjjtnXAhjdMo0irR65d048ypGMQWKpc/KEZMV
stPJCAhnvg5OSSrzgSMP8gmJwccGGGoJJoyGw0GQZIeIdnj7i/Q3529v/eii5166
3udxKbz+hcS1jUUZzcTFL8P5vhqiROQaEngjJOH6wVk4wxN9aMpi6Fj+M6bKpQB7
lB21cnfmGya7KEaVqWMWVMNzX+ZSkQys/QBGWsQhcpY/Tq10Oj8sckWY7GAsIjzs
SnqqHtBciSzPnQeun+i07ClIAAEebChE4XVd1kYORgs6E+78y3MDOOPvxuTK47je
EoMAdz1dshYa2sLHeFPLsnlWMk/e66shQKtpa8nId3EEWZ7EFgy0wT6D5YXNhVUG
nBXgylbBiStMXFZLLH6W/Yx72MWjzumo+DOW7OQ0YwplK+947Dsu3bpnDnEe+d7v
gAxRR+hE5cXL0MyHubimwuGpSoCHiXTCR7xqzmJkffavUkxFZ2oyMDpXrnpICl7q
LYpE3ISdtGEiNpl/0ad2uEYFM/DGLh/Yhyl7Nlu/2GYxwcrDpsW+ZLCuwlnUjQ0r
/LM/KHNbtkY+CWeGFwNYUCBNbcsqnK5zdidqgRFsqy4BsOhJawdPTQtzewRoEy4k
67VoAEDtGoHPkAam+mR9EnHge/uQKXOxOiLBUwb5FuDZu3qTrtpnNaPSxAiZ4hbC
2a9wnlpCouPbUTTB/Mw6KcXKHRpPsNSmxi6mCH53gl5lvUa05YWKzIMxm/nfMWgl
6hxKBCbj7lSbRDL2L0AnJfqJcvzUu+X8la619btM5IsDyrky3TP0/L1TwZ/zy8U8
5d0So+OJ5DfejIrmF2c5HhoA24PSWT4df8YV65zm0b3U2WbTf8hpUXO+eHIwquem
u36mu4fkiIvzQ9dzp0OPgjwwc1ynE5YMIJQ9F9ASg/c242h68oWLy8grE0RO1r9h
UPa6iyt5oWlFMlneC9/QuDXSHyEvclZk0E/8pJRKX+BGPxhSmY7aKuMFANTnTlDH
jopY9eplpsxTMXs4Hx8xnix7Co8toACtvLnzEAT9jqqQUFZam6wOvKpVTnWTnHKE
5HsMcAYmv0S196tE/eMWledjlnGMK9zCJ6g3gH50iisMMBR0FltE7ZEh94S53f7H
YaNiVOQcjuq5qu+FZsZe0U57I1WdqhdO7M8bMD1AJqLZ6U26XT3jRd8xAcwOatGn
ghYYHgGcfOFCX7ZOKsEdUADqNQ1E+CNSXkOdL8M+fTXziUQYwOU8qhloyCSjBotk
lSwOBu/hGKo7tOaAN7gJfJupRB96IFFvpjaYg0XO9Dmhktm0Va7VmWIn1slnBm0O
4lpIn9eyoZKSr0BKbgW68tEWhDKzsvO/iMnBtd8FerwrSRP97ze7OuDcrgaPl7nO
Ihq5bNKfl7yvVKTntWhluVp4mftT7HKfqhThTQs3T6zeUOSDJDZCC9u6FEopJbdj
e6yRVmnzOKcEptNVSkNBOx1rv00nOG/IHKE+WUYinkUJI5VPIS5EKacQ8ELD2ucx
mwriuO2E9kbdcauSlgT6RMzJzRLO5iK2r7IHT1cHkGbVzlez0UCu/6ZLNVUPPmVP
jKI5c7MDI2o8f5XRrfrpn/xF04M0+6gD2SYVKcSmMf5UyShAbgZV5+MO3vEpg98H
GW0ZsPR/NVNbAd7HDg0hYVIaX6Tc0pE/+OJURHTn6LxY95jxbOJNkcNkFVPedR9B
HgEAlAJfjH71ID1LLMLHPhZA5sSLvCrV0KbdLtzBhvtwMsbcWQfQPvoECsx7NBsf
RmDzjsGt5dGB0CIIBdFAsC+t/MXCbJXcoWJMH4tORDYCzE5SeK0Ho9FoRdWyKtnU
eVSrNGa4HyUGLv0zilMHjSy1QgvJn49UtDPCaBwV06HeFDdbcDtvwH115AJQicl/
yD+PVlb/7zFmrfR3RyQ7UY6IB8po7S2uSLupvCj5k25dKh8XsjiuW7pzQI7nf6CL
CKMDlI1JlAviEKMOW1Uo97Ji44i+N4anNvzahlDBOKWXM7LdUImobXIUN9lb8m8e
etBOFxStneKhFrF/WXIECaeXLPfBYrySC5OqOX0VavR8HS8pcQKCPSHmi/M7p2gl
d6Zi7WTGQpZrf0wkQj/9/sbDdbb6IladlJr81KgxajyK73OceNPzobHQT0nhNmi9
9VDHrBgCvEQOcOrU4se1xfv1njuelcM1j5Qv+MswDAgLdj6Ndkn9JRghTv4zb1Hx
7zYYccYUbLSBxkdvOa9jt1zbl1CoRwFUsm8ecrDjBDPehF5RlkMUWZF+xkYU51SY
HCmVtmlMnawmVSQpS7Qq1CjPASUzmxz9O9nexJtO6TvosjUN2N0IN+kEjxjJBsxw
YVeJhfoyII7X5RUVid2M25QyrAk2pu1KNL4GVxiLLO4TrZ3Ym+C3QMWZ1nsKIrJ1
8u9yvs96ss77vswDXgR87n9ahI077EKaoiE5AGKUIl5151jrLgCQXARaF8bdKdIq
eo3BF0crx6C1bBna23Z3w6ItQGwtXwy0rUa2gCeKmD9UjrFpu10jKuduzdnNmV0k
dwvn+f3pu2IfPF6MsaK5HUVmHcgKM/6h4DBrdS8Vh24r+Ixg4aHEKZ4HqvKS2ogi
YsXv5/F/6uoEppmZW5/XW+U0DZfcHSmnzOkC//PXVrRb9wRppImDeQr/7dBtKhl7
2ahES4WrXQ8VZ9cyseFCjj318KUBFEW8lDdb1TCU5fr3/+GlrkB1GqwiNvEXJq4b
gT/BkKOeQfIiE2XuPPNja2KaFSPNRvSO1FSgD5R24Cn3voVY6elRDjNnPL6tnTfW
VxHqTA6zigDhlkUwX/T2xBMAON7jEXriwEEG0HBg9UQea7RY0eQsMWABOmmgOlUn
e2egmbNhnqi3Pye1NgfboHfZHCqdvWcMw8szOkHP/X1XqflMWABgH0IcvvWPVVkN
F+q7IzDkUMCx4VtmU9sE3k9p/wjiTTAESODNIqz3MIYJSsG+2uZUmG7PGRFl+lAH
LTyECbYpS4W7YIZMJFPrikqNudUxQsRpR3DZ8KzczA+W8uGK2lwdU2xcRv0BxzeY
/9OTjAS28GFjMwW3rvpbJyvqwlHXC00l2ONFNt/zaHuliA+qK7XmAohxxad/k8xq
0ErPIXWuICm0thNziXylrroMGBvJBFKxyo4bpn0pkzm+B+FS/R216AgVzRRcvla0
YPVFqT+o3kGWrKub2j0QPg+unlmHVPMXJTOwKQndJLQ79Dap3EAFZmVcpeApR+Ea
wZbu8dE1h1uysv6RqS6Hp98u090KTabRQyyj3e9670WkPRQI8U4v9P9oyD/XM+GU
OvFy4jXWFrTHWzZHsTjv476SVHyd4qrRCFliy8iZYAqE7jP0QB9gb47p45fyH2kp
2rxBlzc7g0yK8gedsUKKqoFdcFmeZsGIlcNReJNGwrmHZlWvvgfA+oT3KxYo7FjA
6e+blXF3ZAA5Z2X9DG/yilsVeK1GuXYIn+pdoucswNCVE+QReoYTT0Tzw3ct3JQE
f9IgjXqNz/IoysOgVtPeitPInG8mzGvMpGTAQDNtJxj2PvcdPZsazyXAWkf39Js8
9B1n/FhBcGz4I1PMpyLtpUd86r7+QDg1gML9G53j36ygsiVAlQ7m9AytdhWGWcaz
r0NpRPPyWUngz+9IRDKrgbNL/DgB+AWkE4YJvJ81i5TOwJZbCzu6MKklhN/mFWhg
Z7z7D5bZwqEZsxoBiNq/TWUGxmtdnYwuPuCsVq4gXde+dl0H7vE5mzHsnWju7W99
v5A4cfWZSselYy284srxqR2hW4SknaP1Tf5zcdEzB5EQw+nby75HEf3cSomg701l
HcAnl2u/6ga2zernO/pU5K7AczJD5iJCXOSclJIiPIxXJI2pwD13FIz1NyBIuyfo
FrClsaA5MQwXAJ/3RPanYQq5lOqjQ4OlkI+pqJiJMdJIy09Fe7eD3AoB2VrnNw8V
yLTsI3/Fdb8KdDRJbQNp9gurpEDbW0BHvXbdx4f4B/SbETElPOnT+DBOxn88RIw/
OQVdaGnaCtsuZmnUo3zbTcb7TQugq78ugjs+HmQgDgSKT8u0ZMjrQdllw3E59BdE
eNUqjXa0Qu4ZcTckitbid00d6sjS6XHJ6RjgrnQZ2MIwfFcfo4Y42bhjhDeIY5o7
j+ln6D+AizeMZAOb4Dv5rsTfIJMfGhW5wf3LG8NlBYRjsy9Rwi9G6D1R4XFcxsyE
ZsVNZsNYRQO81GIVNk52aMWxaxZvWtwQrMOr5mMLjtZYV36lvqfUU6GEAi9zBUNy
Yq+KA54n+oKq6rK7WQTVGdjWuHWDZ9N6ichAFNN5BbZyYOcECcaLRfUAyq7i4H+3
FRR1+Bzbh17dl9WKCpAEtrKOQfduvjAhjEWdcK9kL7B4Sv8TP69kdVKetsvD0do5
4P0v7yxcSdVoUCBny+p4zMJcKwVfYr3nZIP9ObGTjtnyvxHfWLlDE+Vgb4ZOQIFt
lhCQrBxZwwfo6AYnl622iyk00pKcHMfWaFTzXcwIWvBoVuE4lOD4pfW/AwRTB9Os
70KY+eSF/r6pHYcNbBtQP4+muLq3pYEdDBi2WK2G7x8fQ0MT69ktrhSz2IyD+/d3
r+t6GTTGDgToAWUTFvDDCgEGDoj9HetPsmjaDnedaQcgpEAnKYrwd5Ia0G/ubbmz
329ChkdDX5KRiRSnKvDB3aJDT/e+i+0h6YB1OFZooig07I0RTIrev27vWjbDHLFj
odV8kZkEBULW6D/2NAPApmSFCdZuCaiswEaTLpjPGYEUBYew9Fb6MQaB/f56zJg8
VsQ0izPtQd+/kINnqlJYsKxVyWE3aU9aszOq4F49ZMEGIU07nHnL6aFk5cxs5HRB
BjGr/J007CPnVN8Er7f7mrvDQ4PZKFML0ZzPkwTLW+Imunbfj3siEcCJAZgMcfkA
AuoJNf1IFnygtdVtxJhhXQC7RTzvggHavMcVSZNSWBqEILpTXEx7KVNynxfw3HDS
PZGQlkLPdt5xFawJ4ft30xJJC4cpp1z0Oc53oaueoh1UTDZGVP+WZbWsHJPyLzKk
mGyqIee7vQp1EapDaF9ADxAU2iYaMozcvDFbMGELndJ6/hbtzDI5t+DJGslEwcme
veJakMziSZT8YCAWnRGxTUbzAopMtAjxvkfyoXuSEBOLwrmA7z+4oN5KXSWuUe4v
k82aP0HA049Ub5HT1ZewlPnwbD2RHbNJJr9zGXEJqg9qqGmVdqbeE657NaKbcinw
8dnpDxp6f5n5xNQdWk2LKwW58zPzEvXWL1ekSy09j4kXLG9OenfaCmdvAYaAosF4
2pMNnCuVIUQDqnxRKgyHmWYgFFQpFbeeY3QGMlBnF++dSdqGv2GZgkPi294iU75M
2wrvqW8757hvzIDtSuA9+Zwd+FMYvYwBarh847Ch5VElOkU0ChMSDBs7n9iYVTn4
QHYFFf8B+C6a/fraq8gi2OxCR/R784jGlVW83WLGygwldgLbs3oyaJTTQx6zrdS9
qIAxONlLBwvB1vmpgp2/VU4JF61bppaIwSwip8asRFonDPfSeWRsH8zHwn6oqUcW
CjIDygRom9Opqg+IyNJAsnGl4fcA2y6KHLNfxmaPcccgMxeB4p/OjDvNk9vxYmv6
M/j4v8q5hnbXeCgup2zUyt6WgKUWlk7l7S1KtVv+oUNq+zC310qDsGE6DlLzdWH+
mnR2QRMyOz29JyGudqfKOf/Bf7fLkODQpMdHJ1uiXuUs/JDJ+VDoi0zkfZbfWtle
IAf4OGzmGct6odiLx64hAe+SCtWg2pyyEhrFK21zUlkYWLJ0dumv0hHeYD4gEMKA
HnHC5RT6GO/b9iWfSdH9BQ/sZt8sSgA/W0p3JVpwlEfeh5ENnrgpKo7RYaqVCKq0
ocC2REVBFHYdjqs/fk2qxMafk/3FiTdxc35zCoP633jT2Ih3JSnZiVKCYQpf31Yo
AWISPwtwvwlKD7IhwglSwvf9j+uJBTiqXpnFlooR4lZ+Xh1zNGmbIDUm9oUKRcBj
iCmy6ZWTo+LT/2QsXSStuXOgaGWbder/njXFjXKZWmk7gEshqVJ03XLHNHa5LywF
D2sv+B5P4qD02ebx4+/6/Uzr/yEN3IbNPFDWQJ7JiOHhfIEwRDkJTqjTTWbGiGKG
mwVgO0wwcb0/uB9tDu1JMVsnRD8q58Wg1I04eBJF8YUgwzja7XvXrZA8BiaJr3TR
qIYTsqzDLAZ4pN+415D/EOeiBeD9yQgj2LLDFrb9HtHgJsb4bDwXeROBNODpv5SB
EnsiYK/TkFmrzPOpBY6ngX9iabEHiMRkbNHqgH4GBHFgPNm1I8cntsFbvUQikhHY
g/Nm7wSl+PDgziNNRCAi5eA2weR0kMggRpKLRYWVjkyjz6AVL6Sp+HGH45yOChch
OpIpKcfKPOOZ86ey0A1f/85vYVuch9wv5DE69EiTbMQ/bR9ll2T4tq37EY9WT43W
xUclYoSZUWvveDTcL4WSwl90J5JeiLPT4cmn+py/8qzC47GdlgfRDDQHdGvfjm3b
9NjvL8eAtBXQYV0Qw7vU39Bl3F/zKiUrCcR8JHRXsWnm1a0mnZ/vQTXjrJjV0OR8
RySdBx0vpeddpHrmWdt5Yw13Iij6M0EJyo5dIgQP8fVuzy0zEErv6aANl3Gi5JGz
Zkz0lsaEIbrR0ooRwN1fp/4ougrbiDtiWgPV6kLby3ON4icGUGIBjRtPXyhxyAJW
sgm+fSfR17elJ8zZlejUEKtE4lX1JRL179fvl9PvOvQir3kmmzXGdojjZcON8RAa
V1YjTrhk7+VM6Wpv09/GSmD/4jBqsZMdNAORhwgwToE2z7idXfDl0GPT/P4WUC2+
AajwSVT8ycwEWHzqS0m63J0zH8ker0PZr6uFdeoBNQoxgg301Jk14/ly6CQtwf0T
y9PhhvKT1OHMTfdAa8y765ft2ZhLVZgnOKIJRhRLw8Zk0r4oVal7VU1C5N2aKDMZ
cSZtxXHaYm2ky4fHK5MbYDivaNpabXN6vFvIf5o+VJsH5RXlAo72ZqE6XXO2aZKc
aeos9wc0PN98/f+4foJLLGKFo2OzHyjUrg/Ot7KJE9al2x0DZtHOCsPAlr6Po2Oi
cP9XODEB9y6noYsNhCt9QvyqayxB/CJwCLjGW+Ug+VnBAfdQ4AwZ1Ygpomh5lZEg
WT1A+kyvBKSCWOFHpnLn+IA2Y+LCiAbpKupPG0uNNoAVHQAm8lyMhBy95F4JiN7F
85omOgR42Jw/cSxl69f/YDy5J0QYusNVlZanwoDGYp6RMl5LKYd+s7SAqYknMeSy
AGOt6bTf8fc8EHYpx3KfADESrVwUelUjV0CrfzlK9qy+0wNYFxLGYj8x2AsU++1f
cC8Qs5phvsVBv2NBL6t1vtc34mL2bX2/0sUZCOjMC4wVzzHtvJI5nHTTXeUInbK0
IARuxxT+4AXTRKkaXp/X/iXAoKpnoHVbwgYGOdPwxppv41dvvAN9ZuwpieTQBHGU
/hlcdaKquZkiDAWxnlOa1iWcGBZPusQP8W4VuekJir88qh9Bfy2gqZ6cwuUzkM1s
2o6PFGkclB0tP/leC6A5Qn3GTqhpxijeUsJC3l0K4JrOqXsRR/bLylY3xQXKLxCh
HZnaB2rrdbOsKsLGviLCVEZPr1nEulv5wP/ZyG3kR0sDqfVNljtkNT5Me7i/rfni
rafSbBo/3Dsl/RtlUxCyi15rF0fipXpWS0PahmjbGiYvmNxPggGeoFkAFCJG5p+B
XzwzWIIb2qIcBs031WWfzMhMCvQY1ZQ6yWTcXBacCaeZ03tADzgZ8LCZV2ZS4yuY
9lZaCsciHobtHmP4e8TV6cVVetfJAeFgCJkG/8QqCxSjN2dJBcjljrANxT15nFMM
f7uuEaoqZOdjdTfp0rLmVwZZg4nrGsoGEW/8h8ZUJaK7iZ7voS/OA91TAj8tpGkZ
GNj/cSFNsmm5KTMjuRgk/1UVPwgzR7+EcflkD7cYwWueBtmpxSJL1swoBvGU5Tqw
qJ6+NJ/mti/oiS19LJqlxNCo+Pel2RWbI8eqYVRLWE3eN6iCuVtjWfjfQ5LhDF6Y
qG1rcTGEPglMlf+BKgesPyeg6b38ZfpqLYaKLd4FsQYcdE3qpgS+YYtPlqyBqlc4
DFD1yjX4+UUl15YqXRaVwg3PkISN2VaPSRTod6YPUD02hLVbiIEw5TTT9CZxMtSe
CjUA0tkUvUEJcC6yZ/GK6jgW86b6vV93OswRCXVAYjfVWiQ+kNT4fsa7zrEKV4I8
W/r3O9hSb6698sVKD/jfwZhp7kxzsBqiuXEoCaYqKu9WG8RqMI2PpWWku9RR983s
wtS/3xac7vc/3gzdQZZ00t8nER8jOPyDb/fYzsqN0+jXjbYICDg4Eavr4i1kvljI
MbXNkMuc7RDds+YfxTTiQJVsMZnpgUNh+zi5zB1b/9cR6TrgHxm9iYXa2cE2cqfo
6kj6aziBN46V1ElIS4o9CeqyzHd63N4CEZDQ6mrGVCuFI8cMOoikJzpm0kFkayea
k0XKcSNm9CwUNSa06w2lMfY6t5PaOYP4PgwMrKdaOtsjvIqHnM3K2MQvqkFbrIWG
7WeaFDXFYjXDApk1GvqHc100Fp8EGRp9+udqf7G2Nk3LtR9QAzLqXTgsBIKaaPKq
jIXt+Rl3YfqHqakSBPJMsutwH+oGbZIl9dwOAkVI+8GcsqK6OnyxKhM4UAWLkWRb
eJrwX7+vxQ1EEcEtni0BkGhc2f0MNe56qwMDy9ql0Mglj0SQw7JtI7lync+8vkc0
9oS3qMKOtPCt2vASb/SFLDymyh3stpbwk+26LirDeSvOKrVFyfGRG/ECqxtymK/3
+EP7wLPPTk/+U6e6jHTesommK4lmLLtidy8bVdxutvsfXcCpztFLq/a0KWA6+ZRb
RPZGy/wrMpVcarxUlkHdtNgrZEluTeFI8rA7gt0I3k+w/8rAQDi6K6fq4PC3xc/V
aov95wYEfvzkIhmVoMQP1I819WbQszHSH/0Sd+C4Kaab63zNXF6pVy43dGpEAZN7
I9nvKihgAtKsFsx8Peciq3ItkRhrC2QB9Ix0UDARttjE/CwFP9ktqmVCcs81g7iq
JXwd3WznikQMy/HmHQlnt1eVnCOJIsi2sc4aL2MV4VNbs12tGe2b/nZg1cBOtxZa
s/L5GW950VH5qh19aATWyBj5c4h3HST8PC7153bPxca8w3yFonSwOsRNB1wbx3eC
EonLUlyakOSA8PwEXlyYB8GwkzBk0I8dotJArCk04kZiHR0yN+FT44OBKQJK2t2o
fjghGfIdvT//4z6TGszNn7sQcaBKlZa9YY6JszM9C87K2tY/VIblycJxiw0vnPtc
9fVMfRvboO4+MWm8Es4NxIgxZoq5+lMtdbcz1xZMrNfpasAJFvPwX1MuvBOJJa0W
neW0j8AGKodwi0OF0vIdEn9P0nf15Q+ddDqJxz50D9ei71xekyodyGHvBX2jeN5F
TCsRnxQeg2VbaovF93iZSsMcsJAPejJ8KHYpbwzCqHXpnflvCjtFCBHOAOB2e05m
TxXZxDJ02qbZfYQN8imlybQ7L9+AR2Ms7h0VyuqJVYV21FfX6wY6GBsDLnkFJdnb
k7I73w18nOm8wrE0syaPtzl7QEyMuML36S0+Zj7hyGhL5hzc2d0LTg3rEIJfjK35
UCr7vBeDwgffxk4LmQ6fRLpAKsSc85lHtlTaorcKSao3QhOi8WjtjcAFIyAc26pe
AHP4boRxyMcIEXn657TbZvhTsEdOzUB3hKAjBmlNPoeYUpZGZ9dLAtZFO8QYcocd
ylzBFjESwJW7gkmAyTu1QsYCSPMAc2S9bE1M1sKqYtO8SuubyBHZmw3M/5nqpOzm
h3hVadc9s+KdLgtRyWopPxrgN0wyVfD/4Bwsc+jueNkp+o/uBk6LXcdzcPyNkKeM
Q/gwUSvTzpcTEn+HFpN1zLTgnLD1Jl8FlhwJXn0RSLIderFCKCSuJ7Txma3UVEFr
hG6dWO1oqSIi/m56TRo7xRfrjOwZKQc79lA4icS2rOHDceHgc9AgXpYZJfhvaBux
7VyIPt5FGOr2C1dCUCuQg0FlXirNmnaceOyJlyO+3kVVJaSIYF7GhAOPJ82deaNx
K8rBNwNzN64IycN0GEt+CnKa/3s1QensDTL+4epDYyYKSJlRvVXJDyF0ktrO9fl5
AOfHA2jKgUJzqo1dBn8ovLc4DB6eO2LpHOWGRXCvJGKznyxcm03MgXn8fnSx0wnX
XHJMY1DF3jl7ueuoMpSxhO+2rrYXqSfgzQF9al9g/w/0Bog4tC3UDvgs87rm3EvM
TeZs5wog8mnWuJsh6yWJozlX67nAl2n7suX8r9XvWJgkMd+YGwTl7tJOVPS1W/TI
jMz7I5Z/pMfoR+B2YLEllL4pwIrxSUQxgmph1gBQMUaEMS4/ZcPu5dgTIFlAoRRf
4TbZllwRpgwUvtoeWQBknec6EWw+fDa47OS1pMe5Iv0nU7xBw76guaK+WVt8FSSj
4JJcPLQv4ERSwBx/wTuq7swxlj9/0Ej99KVptipNORrFY8jTr6J2EeDHPb7RUgOP
1Krb7wPKZk9Y0fv+UKKht9IpOMTMta2NZHX+xp2LiCrngUFoo1CY4tCKhnWFiLxq
BQw6JqP9Ie44dSXWZl4+WoAFcpwhu/M7SAL2jx/RLIEZhU2TtBfXk/5atfIRP8f0
Akyc7+QJE6CfdwLH4fAwX2VXcQXf1jknPypVeDJzhF+GFw9mWIVr5O420S7McEQ4
QR9U2C/oo37lK9tTKFhKIMAdPUFHba3zvkuEZ3ft0Ek59z0KQiLm0ESasf2gSqV0
yXaQ9DJSrvNL2SBDmvYgOVVJ2p5JFm9ugs0aLRdLaP8Y7M7qQlF253NHuTBO8llU
hetIylGi8XcBfjqxwI2hHKflSCAi47F/eyR4p3saIH2osC6IaWIZbOWlvTQrFkgP
t8rpvPHeyo9vOmJn5ihfDEvDKGJrJsSc29aTZO9sznSqDtSEUKfkWeeHCL2fwX4K
JYB+AbHFVNyJ9k9RMHvm7MwSC1mznSM+HZ5Rhyx9uPqgMfgbRAy9E5C3ZPMnF4CN
03c7P+HoFE3cMDBOl1/P4YKWNomEsXILkMyI9hNVASSmD/6tzpHRrUyp8HM13U6L
2tNtoC5Z9e9SubD09nkMxfrs/uMtBdc234Bhjoo3wPkRljjSeBGVPPNAJEM2Rq3x
6DA6xB0dqdtI+bd2x8XK0U1NcLBXr3w3+fTx5lFIw9ZpcdS1sfAR0PV7IkIQBg81
ouynMuQIMnukUSDNaPaUE3hcO/a3WU2hSTbtKws1u2WAUg1Ds3BnBw7U7PExOBwJ
Wv/R8XQvM1f5L7xe0V8XB0HqJDSDBfh+JnCf+aztgaD/OuSjAslAhMAyEI5zhHCE
nQXGA8tnqS4sxn21AN/CEhCk9mJL9aIsggqK85xWhD9u2Zf2dCrEeOn27KBs3o7s
2pDVMkhwP5L3fc1YT+XEajayin/ZSEUJrgRatZBmFCviKiCMNuxIWnkVhY5931N0
ejfl88IZNO5mpqLW7AIMiCN67rNXSMAbQEmXjzCxMdRDxK4ESZkyT9vwnwpPYjgg
mg8UyZRdxGi8Xk4WK8Nspwlqq0azEzeok34ue3El076ZZH4wcQPCdX6801zwz1yz
7nnwfZOsNh0TZuUlhB2d/cF/9gRVB5Q6aDDd/OOLqIFKqWV5yNtRbumTuRNtU+xS
ld8wOmAUTzehF+gW2zCCUXMYb1r5Qbw0ndQedP3JsIq0f1epUvTIcdkeowaE22C/
Ld+1vpfFeWZLFIJOWXgh0H6B+GOHWBnAj/brk3LxUkNqEHSGwaJaOmXqEi1slf+x
t8K7w29VVKAxyQaPbSlCobZhlzNxbC2UI5xg3Ptk1yBsW8/3/bfg7J6M/2oXSgkF
gV00CoNkIz1mv8Uet3wdDQV5FDLYb5bpowPy+Pd7qwelxnlY1MLukPfMINIDVvYf
FUrgOk5N43fWm2P1sIXbYOU+EJNaI98f3ntwTyN+LRyicK2PscqsOvOJCOBFCeVq
m+bS9neQOqhsFBKrSokwf2TTZ77tCcvlhwBQb1VKOAnU3/Q7DMVDZdH/NgchYNDU
EW9CajqaU3PW5RTNgPjRWHpmrGEZfl40VahoFPWqsz3MPEGm4WUBVyYiPkAV+dcK
cyA6pxTFg/HQknrJIDKQEyhZIhoTgo/vTcF1g0ZjOq+Ylvn9VsS1bDupez/gzXLg
RtiUtR83XIslKHfhfK+jZcgtOQ/2Szz9H3zjcyDWmhmealAidN38/JDgZy4+Fs25
2vhSxZdYJfLY0n8MPLwsK011VBq4WAIa0Fo8vLVVK9IJV/F67JAMwpys+WWPFb8t
kyPmfRpuHkZyip8SexstZ/znURZiYjQm3uQdGg2mqseSLz4rwhsK5r9Lu2QHxHCS
qfhe0OBfok6oL6dLr4+LZX4KZeZeWlSpuill2bim4uJBcWtoaa73WMOfuVZ24qnR
0peikCP7MPaouJuW4UbS10llilVPGi1vvnCKEZxbvgUtiAlO88czN7/fwaBTKRiT
skfI88i+h8OZur0jIU4nLwysqdV/oTVhHrpjK89U9b9mKm3jrh3yHtA3QyX5d3jA
BGRjtyhu6uXWiSdQeF3W0vlAsL8gqXURdUrTmXd/XZvrcCQX31bSHKR7yFVG419j
YXhnIiI2rJrHPKXwzGKLCEseQa1FdfL+10xT7euOEsHaadwI5MtYrGPuD/yk5MsT
k1dC6Pj97MuLWDoBh3WQlJV6IocdaI1XoCCw21IAktC0BWAQnh6wRsUwGSs9tbYt
ATjuss/Tsz2oTxbBrem7u10D/umTllZ5cpxYNcG5yGtQdyfs3Xc0GXCt3m1sFhqb
lAd9w8yMwMfJTyxP8/Y4MxU2uZPgMEkE2lgKn8CTGUynmxMGHGiE/Z3yfPHz3iV3
O5sxt76daGqw59trtdrk8t4d/2NT6kqE9p2j6l2BdWOBLV9dEWMt6Ye9bdJPxYWW
UjDqtx8vnIP3Ag0qquYId2JJ4Bj738s9Gd3pk8zPHvoQcru3zbzIlGSPTKQw5EqI
5P2PsAJqkKiu6GcrcCPOa7RL+KZb/8kSUDQtfFZSfBVAP45pI3N+mB+fhz9YPUcW
K0aeotmNUDFq4/rN5YuhsyFSudaV+kXElhT8dKohn0JaOrcZz+2wA15PQXdCTJfJ
2BFuODNXwautLGG9Y7jGJaxfB/TcCsIpA5IKhZMWeVrGfVcbtR8nR9PG7CvooFt5
dvUZNeyklehnyMLXv1y+X7PFsQbGJ1ydQWNhrRTGHeT4YINg4wGFhSW/a4jiK/l5
FKYNZrwkXxYkf4RQNitgiUxiVHY4nF+xtMtfFLdAg6VJw3T2aeLE40TaJ0O3am1m
vTRhy/z4NJtV/du3hrBBD1/Zoymze+W9ygsg2zjq92xFbytC2B3njQHUoUdK1wxz
gKvipO3WE3o7P5meYAYfTSnRIajcZpx3UnSlI7PWbx5FczI4IJMWkn0AsTeYtBew
MWNH1Sfvo2v3eptgz9g3M8it2xfFUKGMJEPfAB2TQSYhLrIiQK9bXVC5lmLKZ/Ow
p98zy4oIb68puSjq5xRFBftPW8Yf64Fny9VY5XEE9wOpFuaKpcJqNRRSCGVuA94k
cc/HaSarlrIn5ZEe618y7wdWFbOqn7XMNZmR83Xw9OiOT9L6hdaYAP95QtxS24DI
L8bqI81KpTHZ4xVcbi89AYZHgFYFOK8JR6mTs52Qj6fenWFd0RvANRL7oM0q6Lpl
ocsBlfUIThkDblmnl73uPl1+31nPya1BAS7WrcTButx++gZ7E0wKWu4bKsvNtGSu
1yrBg+KMoAWVUD1h/hSMGIbtoikebyYxd6G1pg7QzEtMIAc5vxAKm9S1sdNuB2su
qEbPXjKYzGDZcuZ+tD4XlFof92DapkDeGaO0rFA29kcpUHORF6vWQvhNz0pw0utD
wjj9b0XPP/vmUX4MxQeVAiHhoLzn+F63CaN9VnCyYNynjoWV8IhXNBq+JsWPzZOd
mo1yI0YjIuG/qN+2mWkCk8z3QqzJ/i+PXs7FD95koAqIn6LrRIGt3lWsRZe1buEn
hPDBZcdYgtuw8shWu3oWGXkXUc2KJJiGM6ibEZERVeMq9k+CKuo4dKuyivngGsSr
efHJB6/TyL/sWc3/aaYiDANpGolshR1cf4hVLYbVm8CN5KngboF8taGe4qA8S59C
JV73tXDmVGsrOfsWyGbc/+//DJtYK7G40cQz5ztijbNvTEAKjEfN+/h3PyEgXbUJ
mLkSdqcHru5SZ4r2v6JFhWR7DMD/IR4K4UdO0V3079BcHOnSpKszZQPEdpOMG9AH
BQaBObGBUiOYY6nQJ3ci3qdP56jkxaq9lZg3bmb0YtZH/1+r02TyiOH31eo8+ACe
ZUyFJ5ghLM4eTPHK2+T3DwwHroQH0w1Iajd67XVViWFtyUXuqDqhORyqmLj59MLw
zQc61yDcXpL052Qju+SJBtbqSYqz+4Zaefu/GY4iUseXsvGJY679jzILiQ03UM4C
/w3sgwWUqGCWUFZupGkzk7H5lBEGTkF9/DCqKaOqT3UW8wbHGY07f36zQ8M6bPtT
Dg68GgvDCS44LF54D/AsTlW0RdHZXY2YUuoGSyPfk735z72bhXW2lMR2LWqkCVt2
gjVqfCQWp4bzJhf8CsiTzzYbW6qqFMFS4uW0IITfSeFtRXonNkZnWyGMCz3TCIu8
3jVL3anGU/IVpei/y1JsA6bae/3qS703UY8wbQYiuYBFgs+6ouX6vs2z2XEW1Vmg
Qtp5E49E+AZE4ZP33ySz2r3SEL3k9g/5s75c96xNN6OEGupiitCTsdEukwps1C+f
DlCpxYzGh865wn0cT5ROmn0600zTMWIxcxn6CYhZnzexyLVsmfy310ZtAnACiVDM
tsmic71oQfGfKnq2fZp58Pem9yjo2E0TRRVCrZzyiA8bVo3ft10pIRC0RXl+id1S
O2Znr37RgvKvqweHM28k6PQznS3f+IFmPDcQPDfo2WRLhQz4UmSQOMmchZ1XxWT6
OXycTeEJxqTODXNlLan+csOnvBTdmobYfKCJP+/QMOpHxAbxR0fzjU6TVZrloDen
DbHab4l5FWzhXDJIVxFtQiReNEAu6uSIdlVO4LWCQCTl5YX0adf2eE5r4fJ07j9J
F2lEKZFw3UJbls5CpZ3hl0ybUXbetMXtf9YctCXeBYpNpGTzVuh9rqBA1MwNOsD2
VyZYzoiZgvwN6doigtAe5N0veoRMeeQTjxyaw9dgawOtAgyhxtVA2q+8C0CrzU/Q
Kf3ixOiSv5NZKO6EHMELtqrsF3mACbw7cMTEfEjruwqDqGkB1L5iQX8nLwL0Hyj3
RA0X/E9W0yIYp0VSETify09qFbTBpuce1yb1gtfPzCrAMsPraMlSPiG/DDKChip4
mSDvmGWYXjudGCsMa5Khs6j2UNbPWuVpEnTsgX0DjtCRnjLVmu+UN7ORSbumJzUK
mEeVm59VufaTkMoYn0TiRSgLKpdPcuKWh9ZbDIFa67g7X6hmXk7iKNAzDBiTL9jv
20TFUM/6u2DCQAQKQl+npx9mbOUom1JnDA8EIQfZBClNyusGVeB+cEbu2R1fRF7N
ssyvEzUDWH7vsDLtlltS90Nhsrw0KGbDTEqoGe4M8992QpctlENYlJuNBsHwXHRP
zUGHNANPajUXeBOtJmlEOj3NiJ4Wmi3eonQrsaYgk7RCrISgo8aY8qzGQRvw+UIc
P8BmNLEeIQq/tV12B9Ph8R/sKreB9hYIxT2KGyPmIe69m4feecLQK0n04h8x6Zeq
M4F/VYmM+kTYNVTrhIpczaej/YWrDHDmfDzIMwJsLyTFeWtXquRh9p8F8sX+6isL
TTX1ILblzxtc1/lnFqjiQZAOkjlwTyTUZB/zKa01B3LWXtagZXWYqihkfoMlr9JB
V8bzEJiVJD9vBMf99Y9W0Bv+oTZeD2026a/lSJpESgc5ppYtADKDne9pS47/K6Gz
WefV3epWfq9YiSIOZu1dCTP82CCl7EOkEn9o50KW1XIWbYDokYsFjIIcWHjfgtI2
V9271yokqS2SDWiOProTWaRGMdXnFs2Rb5oBzYtAnK92V8Ygeb+Tih2amt/HVz9k
fr5VPIRWXDeiZKvjyTwffvORsx6ji7w+yJMuif6XkrMzbh7ayf3aVHtsrtQ97Y7J
AtYolpWEFcNTvNRXmLWiKwqun12po1vHysuYs1G2zYv9PFBkJjlJ+oPFVMrd27zA
Xd5x/rtX7Xi7SyqHRSCIlE80oYbNNQF1R/5d1o2PT5RtMPH8+f6pz/KdxOycIqfc
m62MDWuvOJjpSGxObOCivDim6gJJMWqJFVebqe/6SxqxiqP+xGlMuyAIkbcH1dPa
WFQdr9UUeHCZDD1ug22rTwnEl1xdgDZwYZFIyPBhaavbCESh09MMGo/z8l5Xao1O
SCanYPVQ83j5JFDjD7nfTnN0MrKZ28Azwe9ml/ELtT4trqc5EUWH5e+1sXVxn0kW
XZcTY/onsg0NtolYF8F0BsSmb0q4GdAR/EwpXaElOuc+xvlHVJeMjvgVADYoTJqN
dVgouW4AQ/7OEx7c6YNnPuClcovCbRnVF0rfxY6Ft9uh8kGzeRQxGSxuCrgUOZJQ
RlVfrBelM3aJOGeMObNTxQQKOsOghr1kYxOq4BlXZ0UIfmrPgeD4SZ+HYminwOOA
t22OgqlD2RU3Bajf71fzLnPBFKPCg/hnF5deL4KsxdLeSkkYJwvEUfCNG464IL/b
aqsAs6hpwI7LT030NvB3ROoGbfFpr1945sCSrojjaJNkBarmHqnNok7NRvSnjuye
80gd+1ZB362nWboyUnkokuAnCZQ22wyeYq4e6AOLc0o6nle90+BNNv7aYsgtEJd3
zy/RnwTEaUA5+xdmc6HOMCRhXF+o0L6mqBvfn/a6C/rTq7kpihl9W05j7NYAI2cx
C1WCRQH/imzEO8pO8xChBi1PHwGVr2pY+n9OTqT9AN2y31MztzNDhRwuTHaE0n74
WfZF/SD1fz3D4uSnvp36HEoe20hFHxD5g2saBt+zZUk5zncp78iu/oqq8Sv3zbuC
ltiI5PKCJJxzgRxfZVkXKPkvLtqvVUoZf/096+dAWGaY1dRQDDJLL4dQzQDGdQIF
o5/p74xNC+zscPdQjtaIj14BRWCzdFtOYs6W4jofV5jO6DQMZ5PdbebKjZ4LMJZZ
2KTp4156aoLMgXOAeZbctnHoXPdX/PEyGK9K/lGa9ynGMhRUJIPGxW1yh3n+MtiU
t0mxQ0G5uVGPXtwHZ4wZOCfwbHmLFuLZwp8Hnn0kLcqIBheVwU3NTSjhGNjdgBvm
GZqWSWigt3wFhpwC0vGaWknVrY/PtMLLO0wUBnKB4dmg/XixCJ7/VXN1xPC3/h79
IYYpYvaphSN8ERU0zsPGiVCuUyVEdUGnrme0xAHW4ChIl05M6o2M907TnhvHGaxR
RYKTUoeFFtYfki15b3z2ZBbjItsLNKl8p7jkgCOI5ykNxu6hZyCzElM/bwzk/1PD
SlAj3BsXhuhyBMQq2woeuc60eVjxFPH7oZYMHcihhHEDk1LtqM9eJaqVkETOaYYH
DJNAaXStnHY2ecDWzZ0RCVNO6bUZT+iNJJXg/IqaHAk8/qEuO52OtvE5zdiAy6kZ
trvzXw83G6IlB9KQ/51dl1PGtLxZE6DaD8oPISNsRf+N7mc/zOQOZ3OPKZr0s81F
Of691qrZ7rQ6aR3dCmpl2Y0PDPzrZfy0DAMB8kwDwHdmW/MfVj0HKJK3juN/ofmq
za9/FYPVpPLJIquf8VrX73y57nc23UzD6sv8qyZuTYzHwH7GWSl2yb8UPWe5bLfg
J2tyh+mA3Z52LZskb3ciq2SmtbOhgl4IW3K2O+1fbg53xwnmun8LQtnECss71HBc
FT/4oymkzGQKgMG22uf+7flONcw8hbtkwv9Ot83bG9Qbc8v+MtbP9xHRdfTvh8cQ
SnyFHNmRST32uP8KbVQDfJ/g18l8oatbOuxZ0Z07AQj9BNqIFkY2HTytzJyJQ1WK
69inc9iisouDFU4NyW0c682dLGfV55CMYVCATXNsjgzIRWFwkyo2uepPq5Ff6bsj
fTrEs588vxlyU0qM0WvmCryOQgZuTCBDtXk+I5tLXe2RDtC4RAn9Qhlq7qwldMrj
ceBIJ3WtCHDj2fzi9/uNe0r2CDm5GC73jCN/9hblACtjHibhE9makM3Mz/SAbwRH
lNIGA600mRkphg5m7B6CPd8CC+Vo6oKHMsBYdFidR94zSw37Jgr9vm2Neyn3oUqJ
yHCOlgXBZKfvCEPsKByPEDrTGLuwrkyjSPVb551OmY/QAH4biotN3YAIk3ROJo/g
ejAgFQtnykiefffAlFxZbi0oEkpaKwLvHu3aUgNzDWsRJ9Ju9HO4YbxfTJc5lKfL
lno05ZK+KOsj7nQVG98/NFfhadlpWnfFUOhY05bXCIToHzsvjNnRdZNqFMwj8lrv
MKOh0Dym+9tvVTPvRaDqdIa107Y1SYxTNKeryIlFtu+7660U5xCkUBVtYaeGFvca
FVBMpY6yRWoH4yF4te7EghOMKvtUbr1n7bLHOpVtegeG44hiGOrbvy/1gAob1v4s
sLXKgwzpKJC7kgZq+8Bfpy9qyBDyLZdgB2KRdWgQu4jWXAhJ3DvDPUKoGMytf+7F
3U6VWBTVzreeA2u9tp1kCJR3v9uPBm1Ho8EmRGfl3PuzGwgzVi8ChId+84mP85nq
On5QcWRnJhYcOcZAct5kCrvD0rMxNvZqZNBzKZC7zToq9tugHNaaASYVL1OXp6NA
O14w1IhozZv/3YkJva6bpG4Vx6hxl0nBNdZpCKiKEweBRsYuZ5u7JalBWPV5XOaA
rZHqoDigJxR+P9uTghaoERqwVtH3kw5t04i9W5RM8wP+bps6C7NgJ2/e7v8PKnIN
bBdzmJWgvYD0zYKk1lhCto3UjsH5/chLzg8zzDT4A65m4c2I44VC5lzxfGOg6iju
gMp5do8Xp2a2W/MrxTQWs0vwaDegCeSl1I6f//RwTOXErueAzHodntFVkB4x8fp8
i3HakaQGtC7yPU+1q+hkXSm6YW3dlmKKnHlaRpDW5agcq4k+CAn2fFX+8iLugldG
oGzXwB3FMOQNetQeXcIBUA7muzU7t99IuAYaaZMye6iKR8V+KEW6wxkqGBpBRT3G
a32iQo/41a12qQAF7gfV25zxrb2w1dObfqMJuhHu6vhbtfQTvCYoVo4VFCUQWMxD
vLOeeLT+fmw1tFOeCzYCWyT8AX5XX+d/4JtBw5Q0Ci35pKP6HSnj942xvxmb2nGb
6OvHvsdVlSAuXMUeGDv4HbLqnjU9rBxvFYukeZcPaq9xsL/3YmKBfnMMQTE+rL/G
eOFR8KxDmmqIX3ZMOB2GviH85sB+INNKK6Vd6UeWpEgzCGV2NKjrqHjnYH2XYITo
PfBbNLpkVuiCpwnUMn/OAKrgMQIuuJ4YRHSfr1fGjQmbW+fGVzQb8mP/mt/HkPBp
o+xT58n2qlOdAqqcpCqn9zWNzexytT2XRx4i5BMsEr7EtqrKhyaoRb8nBOuEq7Rh
nbj3pyfC5pdLR8fKp1S66ZESR3M59REW9SM2hjRYt8Ub1VFTwYj98eVIrshEJqzH
3iwo149E5l4xTdtGRngBxRcy2a6kW1FakxkZobp+h6w+7Rrud/NzdIyRIa/zESaS
GWFOkkmv7ZVomm8rXKnJNGH74AWSiqPlCrRWBqw7jSSKD491FOm6PbE1qKGtRn69
kBOBodhsiY4E4hbjzvJrvbKdHXrVlt9d9DLhKNol0EfuZh5M+AMGAvAU5qh2WVM/
gSM72A/JqhEWI37w3AIgb/keMA3TMqtgqoxLlhrPb7BcqaMbt3D9+VpcfJtNlSe8
7yZ6lAHoO5NWkXMZ3U4icm/QY5xR6rb4uDVnF39QZ+ruYHGO1KWYJRtUqtig8vCO
3IQtoyioYdaBb71XqcKgCcsWS0gUPvPGNusO9qstGKMAdUACb5Wj1fpZ16qkHaVr
1YCSkzbwhL8uXVUQNK5VBvSIz5LpHUhMVG3jdSaKYjBeiLnUgxLABC1HxbCCq4NE
4w5KWLrfbpHbT0szPDPTWyUWBNtbgO1iqeqqDVpFEO1NqdJ3Pb6pV16YVVqtuxNX
Q1vS7u7B5XKLQQohVBSrPg+TQ8bYQ0ww5GB0ZaN9InIUMIcbig9Lt5LS0IvbZXSS
qaF7mrxez/B7iNuGTMsciWKn+IGGwxQ47mkSuX8knq2PpT8cpK6tw4xFIHZYRZaZ
64Vj1Gl2z4bamQyRwoID1BNcDBvn8ozTRWo5tdR6iPb3QdBpphWPV3EURg36CazA
LXbiEwEvMBGMtPZaOmC48GCeZmwgPxRraqV4dmanAjEpFCHZPFQeotci2bomt7+8
RLXuTNbX3dHc8BZedILhD5zoYi9AVBh+5c3c0oPC9gkXDIIVNuDY9///E1Ncv31g
shLgdSa7jdJVsHbARKlORnML04ptddSlvqFmDhpRpfTGsf0wPjmT6Xdh6AZFU3iP
tPP0St+Lv5PDrHMUxPTIeV2/dg5xLXws55XR+vNs7Pq1MIs9iRFTREt9SXTXPbDs
R0yRKczoHhUrf8z9fy/QUQ0vmRPwZh1ncVmjwT/LuEJFVdbSyBbYRDiKzDwTqoxH
4+c+e6vBQQY0bwxVWZ/iAKAZEYozSRlN8gEc4r5elbtrnmHjga/dKhncKvwN1qRU
f0sDlmISasaUOFv+GkWFCnBqhzKQurmDkf2azcQpf9JdWYBfVMngNAbq5XrLRMI2
9pGQr8VGVhVIDqS6JU+pugazX7oQvpkCRiY03btJqoNlERTWaSVXcOwbU6zdBwPy
OIb5UFkhLSMAlcjcTxw9oDV/FWNU+HQGnGGt6uJVigC2SyQdq8NyOhpCNVCNR5aI
tRRwRN9yUsiFQ+dtlCJleqlIlnElhpOknNBrZXG3h0TK/IUb2QuhNZf1IHTpNpqu
D9mq4/CGyK9EqdbGP41MV7lAS7wjr82EVp8eFCxgY2nZCIrkMyK4mlu6Wo40JJ6Z
uksSGlnLEF+HgLil/QZp2eDDUZgPxzNU8KaZh9bwJsREGE5JqnKFWn5e+ngtUny6
EBieQfA8ElSFJCexGAG57qP4Epa8lansgK9+TLQo5jah/V9uwyAkAGwBDWf8porR
r8KWDeI6D7ICBwinbcir5vZ2ICNxVP1E+4Hv4Bo7KH6oPbozvnHN2JDBDR2UyObN
slbY7V9ANr1CPmIOAMWZtNxgZcbaStFJNb8b9cpDaNJEJqtB3Znsk6zyDkssUI3g
RSMrV3ZKNAa1OlYPF9r4r3ueEb7tIpSSJnGdrIwaP0YC3uwCpFKHpy6bFYcnwORT
R+3Y6uWucFlbrmt2TvMEBlXpc8SxA2Wf58NWo47vWzUgCwgfczBA8EyShzvc0csR
V5+O65TSqzy1U0y7IrASTZ29mFE/3YDEpZ8PG0aovjIZvcuhK9z0ckPxXQa6bzzG
ZyLobj1u6HX7V4BecN/kqVZSWzfrSv/GUkbkvQ5bUiJHHXl66bfGb9B3JWsQV5nt
3557uQ020q0lWLpFR+QWOuw7t7gpfdaSKRGcnGSM2QadWSxNt9gZk15BNkhLiMpB
lyB2zR62Y2VPvVr667lss/A2LmIx3zYUuZGZ3GwphOZpFKv1ze9gja68r2n+gtNM
iQns6+E8NhPr4E8/dZsopX3QC+P7s0brffWalVqTaioTYjQNLS0//D+JS4AbAhOy
Sehg4sb9fuKVLabY9EsmZ2phUlx6Rc3YxtT7/VgCdCpSCXKbsZd+xoxlW6btL9xu
geYt+NdPmfqoQd7wsCvwEl8vOyWDiNaNLOGAQWRM0xy3tOppVyupZ7Nm/I5vHiaS
dobIxam9+5XhGDf0hFP3DSxd0vAhxgeAd7dQMlhp7VXET/5TzIfpOXhdhmQAHh/v
pj5u3nwHL/2xQ0aJPc/NqBGcKXUWzqUXdym5EDrZh+QRtoRX6YO8+yT9bbqTYkD5
w3CAcI2eWY46PBPRSR5P0j5BGEBHD6utpkOroEDK1N9erFCg++xTwlMuLq4AExY5
F+fWcDuV7pjWBEzwnPYqSKG5mUNMZtQ1xjub+rCc4+63TJc7KOfzoZuz4Z+mRhKH
VqYuIL+MFPtjFNq/MJIqvY14SE1l+toVeZ0f/HqLhLDBEWQnfMotaNiMib2rrIKM
oSnptP7N7AHSR5uMaU6EEod72hV/Q+57i+z/WstLo2t6wMsfFm+48PJJCfEpoDU/
dxQ3y6zFUy7I8QRLceQ9hE3rCCY+UKxXfLg8NSgUqOZGwIj+807FocT/Y1JAibvX
7mkqM5t4lZjK1LAFrhAvMU4xDAjYA8lnVMvfIvQD87DHNx6TsD53GvtnOh5czMBV
OUYC8YE76X4BnAaRFPoIbY1gkLkft/aN0dvSgGNa+oCMW3P9pm8DlJ6O48dazBL8
tthZuuC42qWJ+ezD96BdMzQDP0CcyG60RlwYyEDXTtp2IOYXaXZP202Jn0Xs5ORN
TEXI1MBhA8Dmy3H8fRsJxJjB0vpQn0BI7v9mUiSyl0Xi/YwOZyWCKlXoTHDUA+Gw
B0PAwmXvV8kHVhTdpqae5Nehr5exfXpvXlfs0iChkZ//VQsudbrUbXklTyt4ESyY
5iFWABclS7Z0dH8upHp3E6lpkVAxvne60uqN4epwIClBFCilGZsnPgKDIUPfeHI9
+mTk6DuVvGsPoOF28p7FjImjPb+Qqp4F9Q/LTXULm/2AoT8p5W11ehtcGWuDm2jG
WV2J/ezmi9pPqbvzSLlJaR0OZlFh2zKNqliKtu1h3wIc+QtEIrKL5tVvJjT5mMWD
oKi/4Q3MAoJSusH8WCnyuow1MwZqw1dFm2AcYcyHbgvwet7FEoRjr0LOsNjr0eN0
htG24iz97hBfULHDSLQ4uZnwDGV+Qk1sksAEAj6+8/lQ4gBdxv84lENjrBD+Tvaw
jDyMcHE0YA4lX9FIWwZgbArMQ09vChSzox1nTbSkFkaiByGz3V2lhUy6OKJq6ad+
ZYvM8yFHQHlXOgjfJhktSXtUifygiuQMEAXEJEWSAj3FgviDCk8SEn/Ts48JRTBG
I3RMkyiKYNtUIdMo5K7SPWuwXtzKaqr/3p9DMXcXmAXP4tgiBR4Ng6rZZAgmZo0+
50z6GPiIY+0msXw4HV6MpQd4IGdTLeh+v1jFmgLJIAghoarAsqtO4zLRIqhSdVI+
48wuurKnZVpy61jupMrNu4e0gzSJVV0r8YUsZxsGhooeaMd7wILAiHoyXGKizwO6
sDCbq1EKsiCPFtEFmnnuPiINcaF4VyqB2i81lddGxL5xn6F3F/Wot5XZh1Hh9zH4
HnIwpDCCiIadLKE+iqLUdXhbW85TQbc0CQu4BQUmrataQXvJ4m56Kh6gHvSQXVjs
TZmnK3I8b7Gw0XiV/adrAef/cI+zbipnA1A3lsRxlLkSuzfgotVyPNUkS/XvjvYj
OoGr83NDBI2e8W7gemswzrCSakyO/KuPstNx4dwi+ZT+sVP8eWU47pwLBjVOyK31
SbXoNtcYwkbxsfxAAjC5/uoyWNN4HjValXfJvw3GG4PzwMWzQmauz70VDRngGMV9
gzamgVaB/xOSeXPeSIPbGbxRqcQWxUwf8ZOTV+dlsbGR7XO7QeWxqIQJPBgv2lEr
bUG/4b3o+hIugU6+fpPm9E4WKypiIUv1JTWX5sBcJkloFpgryPGkYf8dmJT9tixc
sQ9Cnx9GaugJryJyQcEvokUIu4iXvmF6uCL6OSOA2AwvTUel4nciTSN/t4TT+D/T
+6NdcEi8nVuUIt4XjR4tshqcTbBlvMwewkoCoPCTLbeHf8H2lmqVMf+QXfQ6e5wG
dqmOSlFvO/XsAO8HPTtwGHViiQhusvc6PP0565ULAZ72RGAifOxsLp91WGqGgUmv
DeUXWG4MjOD1rfZT+vHcEFy582txI/DsSyELZAF2lD112W0SzBAL17ktQyQL0ZdK
N/cXkCjfwrm2FjfjIo+AoQv9DrltXFspg/Y90GpSgWgIeF9rhge3annJ71/qDqd4
PhomorPTZiQRbLiNKjcTWF7mpslHPxPHffDrjXzVRn37JuUjkCUZB7IOdV/H9dXX
0WeBpuZH0867WZr91JLQQKZWBqddW26wbRIO4iyUrYriibt1HaW+22PYW6Wg3g7o
eFNIYhxpqMW9RL9d26C3fYxo+J7Y35A3WcAziWYqvZP9eWglj1qxu0Gmq+WgwPGG
MN7M6PAvwBJebDzo00cPPD8hbnIXEPTVWr7Y8lcxom2rFSblGZPmPIAKGgbr/85Y
cAiNFkZmHrHa4VDQ69SKMIVOe/cg4XCvmOdp1btQbjuv6u1tfQXmp4NqyTWNuYnS
efCt20xlgOFFHsBO8g/9pYeQrp9Uo+O7EftShxpCosK+J2ZxNbS5zzGecelAvAFE
84i/eGdGIi0xz6jcWyK4HZADeugnUCz/hnKXHa0PRn/hBwAlhPVlU81VQUwHkZqT
WVnW2jvzkQlJIwceDFcjVZMcJLwxfAMfTxnbK/Cj94l1kExONKLlwF6Jhry6hzZa
A6ZIJwxFt86DU+DyL1/735LFdSE9QhG6WHwWoFBB81HRgJZPS5OTJ0gb5PKPMKag
5jmM34dqWVe7j2cxMWAW3vQ2CZIHma627PfnqTQ/BZ4M/zM3oNaRPg8WexBBGlYF
zB5Tgsrpg5lE8bMtvCD0ZMGJa82sx0OI+a+alaxWoQs7xLgO3oOieA1tv5HSgA8s
ZQl0udVxDIlsAS4Bl3AgK0sy8NhrS+JgO8zuzwSdyGZvdt7rkCK+ykl2gAMvJGul
sryh+QjrPV+hrRmvqd5kq76nd5HrpoBNbTx1/49SOu1/yS1xmXQ8Vek5HI8MZKXg
1oWR1ECUl2SNh30mgZp1zk9pcrrMiHw8FEl+f/lxfMIDodtKe3Xf21pdfDo9bpxm
Sy0LAQ1zD8HIOro2X9mTRjGEZbz2NlS6YM+8x0njVm9ydbZZYzOHAPec8CJ0rdH8
IRgBb76TBY6jx6nIxHyXFxYL+QjejFc9UbKX4yOdtGIeiN7OPlUwnx5iGfoERN9c
GAEKW+hguSej0qmf+ZYH+NoV1K4tXXsyNZWsQjPrSuEFRnosTcDeewKeFVztVb/V
d31vETTOgQfYhsS8B81UXaIf4HAfyi3+bT1JhzaCcl8S862gAM5LjzWkW3FMSbmb
1prJiW8q4dCLTE6m2qpqehdui1qVwKMITWflG/UhlnZqNE6seWKvUFg2AwaTuhHl
kTzAy64nz7ee0538mCTEYaCUbagdSB2oAU2Nc3lDTmYvOdCsJhG01b6aJEi4CipJ
fsl6DkIh812mBAh5lrh+emGA1iKIwHjjmwvvFFtoXNj2RID+G17OGPmiMD4Q8W8g
9DZe5sxGgsnhd+cPv28kLfxvX/1CQATgbQVVoYyDnHAKTIDD/DGDyU5aVwf1FLwD
GK1Io7EkHG4Ea4ffMO2toq8qCe/6l52fk/y4tIvYgrl40ftzaIGWcuX2G65ve/m1
i0gkPNn5FokT2MtNl1K9dhtFHDIhhjMFzhp05QwRjaNifRkWPtpP2wlyoIC2IIoS
zePYZQ5Vx9PgJw2fsxBR0XYumyXBvlrNLf39yFv8cL816lKNGWFZ67B2IBXYXmue
uy3ytL8OCvpSvzXVpNv9i5wJWESV3rJ6IFJgWzKzVcREVQOJ03siaUSQM5+fhw9g
SllKYalHfcu4y1XjcAmhreuROqRFCc3COZ+sX+nknHm0lr3VlJYdTaAniXJIxbcU
2D9nwUeSTP3uUCSgCtUiGZ27ma9bQAv105c8TN9dGlGMzOSZBiQlSVKZOw5+RydB
d70m5JGlr0uWdi0SKVjW7kiuLv4IG946fg9qHKEz8ktwP8+N855uLPttCz7SF0gB
+M6wH7IaGoLEvDz7tvW2HZgo9/VeSdXaPpC1uoUecIsvgm/cJT298+wqAGXTMG1A
6hXgbcbZNRnG89Oaw5YAWqCtKg2baRxiZZtXE1mUZ/aucr2MO3Q9wIoYH2qh0N/C
lsEOX0kg0+K6z4Kkcieu9JiZ52kr8IEBR5YavZdksolzKoQhiHjBxkRLIqsXAPV7
ih5JaIbmXrdstekn4iIyCCBXEMdq3LIkJJKC1G5wry/H61hnZouzEPBKakPwFF+4
k7tqByEVYl2rfHuvYnqH4YqOiFCZHiE0iOauVftuNlcTT1zJI3+5P9BsvwqnOnVp
6H2ILLw07wvsAiNTbVWpUTRdxp+Nk6DnvgcoM7DTWpdoqS7zU9IYf8PH8BCkEsP/
UFJLu7RY58RXmRHc6B2O5LFLCggDDZHvnsbEd1HPgkBV39Hp6bsyftORrorkYQf5
5fcLexBfAWbGDWOoL0ex0YCiVEtox6KmDqMUFcZF7adV9HY7XTmz2Dzi7c45Hf78
MCJHXp6tGMELIY9lQ6ENJQ65SNHsViTmEt+Mrreqvt4S28wT4sHgq2eQywgF8Nkj
M9KgQ7WTPPwTjP1v2x1GIxcrTvv+U9zKnSbHlqF0h1yNyIpC2BK71D0Lj+OHD7E6
sB5Di4LP4qv9gmViDxiCEMhGLhd8GAw/2Ock9Xa50uu8EkUNj0PDYsmZtcGXkOu9
/DZFiy1wWoOXy0+9wXV1RI8uopKk3Yhz9UASwhExpqWBTRLcPGCiReidTJx1CqxQ
wJp9ROiH2eeRsW4Kh2lhITODiUPYRqPjHurEf+lz4vOj/K9eR4MjuN6H2e8pcg/X
yqPJRNOno08e5zuLSsYFP0Wrkr9d3UUHoLakvl1DzIhGsZpakiSN58fSMvh1Yw4A
/caErA/Cz2YmB84KepO3MToWo13XUbGiv4ZqHJYbxqpZ8apc/r/nKY+Lam9jOgrd
/69bX9Deh6NcDXEHG54Z4f2v1rhr5JWC+5SvwcOXXUM0FmeYAGR1mOpwmDPPhYOw
Ert8rpYron7exl7+4M97ZuxjLFpmxsmUzoM41khmhUhz9ppwNAnIHEUGcw0/bRxE
zLwWo3c1959cDjgOIQkNH+e4prvZyyv/uGrcy4QMIeNF2Tih1N5i1io5dkae3RPT
/rr9rMcRDatSqqdIpa72wECHTMTLwMTzQDIy4XYVBOMKYJLwJyTuxslILie52skZ
80pI7cO+YFigxLalUCjdNB+Pr5n6dWXfU/PbKvzIv67mg+uhyIiWcMMt2d35M6fb
tywVBhk/e5+OH3gsTL6Cox6SB8RRE3ysAo5qTIm0IXgBv19l1krRqYgajhhDi86+
KYjZJYTYwvt+KtIiBfPQ1ficaAum57Dlt4h+2//nIaI6AzdzMsadojqIg13F2Ivm
OmhmTLP8R826Cb5g+wwxbUWJCHRg4tKrb/hRCkfSR569UdDQmw6FUNEE9WBA/keT
lgyFdPHGHPW+PgTCjZc5nAYsemaoXHPln4U0TvNw0g7VV3BY1xvz9ilGWn0AUaXq
OhiXAUfbG5KuzGG1G1e/HoztDe5HUrIyr0yxrCTqGsGc/6lqNC9zI8bt7ti/pxJk
lW8TZm/KI75rSWVcDK0Wjs9yYJK5a3OeB4tC7iaT7A2vjgBTuCazIWWCSpqb3VQe
MyIKOpc0dtOBF2I6B7lALWqRDu+mhlguZpVD1+SHo6DWhJgqKRwprQLSX+46t9wp
Kksi9EMPOxxmnQLjQ6jiLth0FSIEEwZLHfzj8U0fUJQP1U9oS7fHgLhNxnpKgXsi
XKOQQc+aFNkmGuyt2nopa8c77aeSOU6HdpEtuPnw+OOaC2h3Avqfyxze+4s1hnjA
Ck2XkxKzRQoLYJaRwRrGvM9wttybClJvZnnlN3lKPKOy0WZ6dsXsLqri0JCTrjyQ
zmLKkZdJm34sZgwNH7mYe+1fiuWkMJ84D0+SFGJ13EBV2Hj/uqdbJxtlXzmpgEmw
RU12hKARsOXeXcIaWOrBkMaUNKbLAYsNdUlc9TG/p5k7oJ68E3u7JfiBlZEKhZAP
4Gy05o9peTBTwHsfXX+8X8C2y9F9enWEJb1d7tpU+2pjfgTMJatZnHVyGlIZeIHH
mfzWyCNoybYT940tmb4Kyfs3fV6VdHS+tBprcNutfvfv/dsuc4FjjpIRWQe8MdLE
nCOTzE+rKxw+aigUcbLn3lEJPulTtNy9CIuv0AMebzJnh6S9dvTkGuX+pCTGhDhC
/CY36sdZpX50oxd3tR71+f2fojwJijqwccwKN6JJA368PmKiBxgXE/oqkET1uqkn
8kavDPr3DUqkTGVMjXLXqPkQrUiqNN1DAKwl9zos/HruUqtC84HKFlBti2VZR2i5
QXMaZCzgjPGIBdDR5sK7OnQp7m+R/fRfr0JhtY4KAeBM/G2HjINZvsPlqjD2kYUz
ERezMrhU4BVxOEpq3TSM11RQkmTWUXNaSroBdc477pBKEAqBkJVR3xXxgZDXWUpz
GYmJpGY2caXYf1TBbpblGHQ8eLl7+Ltg417+nGPvEEhhoxeJc8qi5TH29wNarI5L
KkJDWBdzRCtXcK7RtTxdydPczJvwDn3xvWy4pPlDCmDHt8cACYKh6t8BGmGKmFuP
zJPaF1tffXs59dJV38cE/cBCWxrUvWFXG9fgTF3R7ZdlcQRwKsbESbHSeLmwrwmO
0+IBrTy9mwKs+gx105Iz+t32bT2i6PKceqSM5Tjn9uBAAFpwMw/xQfRAINm/2CXz
WuIpasclYRoJD2aZBRlp6uJjlv/dPzhB3y2RHNwBu9Q6aW7XW0Kmnhyd7ifn9TCY
LThHWbhjBW8Il4HTz0Zry5xipMFK3zP9pB/ono1TWpC/uZ26ZlPT/Q7BgZ3+r6fK
YXLajpgEOYn5qp3bskP9gCJO+VBOZu7wNMF/JZgSFI7chukuKIQgDBA90NOcY8jH
pYD1w0p0VkGfSAlTK+nQ79HgKFt+bIKloguGEKQpVjgzSh8vbxOCzpeO1tSGkgBS
5Kj+XpmXfV5n1nfexeb8Eb7oYpSqJJgnu6Jc6l4e6Xa4DcrnNBqWcl0jd6FuoAEw
r4qUocHzN6EFId9kZPCzUAEm6Ww8if12pCFCtkSl0Y8qfcBUudRE4SnllbheTOdp
Sb6nFSPgnsvrONGi18yJ+jUhO42CJ5RZHvIURZ9hS8qaDk8+TILc+dycQh2R3XP/
tLdE/DJQVNiydqzXzuhEPGgaRXR5b9qgaYK1irWsKnTSZIzrRrp5+vEVV7yEee/m
/NPEFr76dDOtJpaEXUJo4ydWBM9g6K8bKEz0a0tMyD/IpHvQYFInLQS0MPJ2Yhxe
Zs1aiyrPPAPHcGPFj+rc2myeSAoOlsOYM2sSrRt4mAu9I53VZhuLZ6g3WR3zu8FX
rC48kUMCe2mECLnWH9l7xDMzZoBQkxD4n4dKMEdJ0GC0sorFdLAUKkI81JNVoiYe
mwKJTh436TROwbbNmIy0eu6qej9uCJ/xpV3uqaJh7hDpg2Cptyzmdiyljz84brU8
ZTMh4sdsBLE2t86TxsjhzmrVtGlt0A54+esHlPNTfqacKc5S6mkyarNISVwOzYbx
Pn/QJmBag3kzHJ8Rsn0USfNQ4kp+rbFZhSjj15DuYi9EprCk/kBFYONQUBdXUL84
yHLIP/ZCcEiyPmIALRPTK/WKq+AT4t1pk5we+E+0kTaAMuqpa4awSvyeacqBoO0v
VkD/aB6JR1epBTlkaMZfI0iHLJ/p2dU+nojbwUkHn0Ccg1HrYtam5yQ8aHpXwKyl
gYSeXx9RyYTcFLhMU1Xc8uahPnjrZw4kLK/34bJY8hcSM3xguYINrEZELw0ua5Nn
UHRIXzl6YPkFsGBt3zUD/DmwOImT4Vi8+nlKqJZz+sgdF0/US3Vhx1IOApteTUkW
Bd7b2FeLcI3b4UxToru4TE5tQRkR5uj26EmeOKAswixL+YqzvUD7rjfs9UB6JFdD
PN6p7Q9S1kfFo2yCSrBLKjWd3ybWIIDlx7rnFTODSDlGIB+0QdrGFxNXCr5ZptQh
LW9fJURGBqx5mRG07JJjXJIBRMHjoiW9mofMK16/HEweIM2f6YS1GjjtRW5t+HHe
rljFGK8iA2RZbh+MRdR5q+lSSEkAM4/+ixzWwo13y+/U3/LrmQkXuOeNvcowM2U1
95pzBiV86jZJghTwEqshGTEiHBMK+ol/yIi1MG99cyCoOYKOwLA6UXZPuZKSLtIC
OtXEwPB7r1BlKOyy+OyjEgVfoFgMAxt5KrzGKF+A6wFMBIIfQtOWD0RI0hdc3RW6
qDoR3dsRO2sLnX6Eb0jENoTweFOd66lWp2mo6rSrY+fAnwgxatcbS6Yz3Wpavzxf
FxVwhU7aLLUHc7+5BKry5F4LRriMcdhe4dUJihbe5xoWQJI/ziBulcWIQOeK5uEX
M8cR++GrXlKFZzvNhw8JLmPqNVfFh/g4LHqk9VrhgK0klIZfXgCD7gOdmiome8g8
qkNSygDXXmU9+7zxh8tMEfaNpt9x3GsJcVjrCbElHqWbPihPY8Yj89EQVMUUdtqz
TKti2i2gNmfK0pYQEKKcFd4wy2mh350kXHpzbYd/Oj8xdsEpjHICXGU3UTMTp352
vWbcDRQglKVTUY7hnFA9YFcuezO64Q/9s34IwwoTJ7/qGrCss1Z9WR0LbVNr4ONP
KT21C4FcpUGiUuG0W+VtWi6c1c35PwGITxJ30uYvD9HgrEP3AolE+YXCv6sxZ3Mb
Yq1VyMFWdVXv1DHRBwUpNJU+/8utt51a+OKbZgwLeV77+3KuD1qW1MPGNMVDkpB/
iA2O1ic7IzRo/j2U6tSIFHyh/C5kZjW31gjv92JGAIwAsrzMt0KDK1MGEHB1mx9T
0SYKBcX+3BO9/k1xFpjkUeMW+cVwKu9a3lzVSYl1te9IplKN4q80ZpnCCfyCAgiv
cHjzf/Hk5mALwTbDuT68SVbt1UX7FUG7oZiPhsR/kSOFA6ha8TZeHc+/OHwXOnpj
RXz1JAnl+Sqmwl1xvj+BEhKWbwauQR5VyjPoK8/CfREqM2a9MeL82s2uvsrBpRtR
1sWm7tHJOwI4w8Fb0I4nOAWeErfcIO93LWAbGy2T47/3A5QLEdEBibHxAO87uEW+
8wwS1VC12+B2uQ63WKBhgX4qA47+EwHdb6wbSVso5ok3HjIUJY+C68O4ZwjsXGsz
Dcl0QOdEAZXB7NbZhwWRnEUauETtwOzSRb5MaMXTjBFHHCtQX8JJeko64AnTGMU6
cFgopYZ/Z29k1kR3//+V2FNl28TpNBuKvmK3I/l8la/oyvfelwsZUgxjs+iiCXuE
sHEWtBP0FkidDvKUGbo8fOdHgNygsd/ajMxri5YoPIyPis27d89xK4wwglnha4Mu
fXIg3miVnFi/AxlOzl1TnItAVJBxA2Ultgdn/9MxYvISpBE8XQk9CP7SHiZlM5wd
6omcQsKo0rspu6SXPnEdLL5RyLEQazWJA5OVpl+BC5rYoZ8cA4fwHxtxpX9ynl5t
9w+oZUGV+u9u4u7DTf+OCMyzRHAUx2ogu8D78KY/ny8N69c6yqNGNDVRV63KI0Ev
J0wuls4Q6HmtT1UF6XDVwrk48Ku+gqISHVXrkuC+mNCC/bBGHFf/TZriCOlxorFh
3S90ErTOzgBj7B3IWy6u1kfLsOMTlQohZY7fx/pOmlaTBKFZPRvF3eqGxxzEm+ON
upMevyrQeVx/HJNHvGkw14sTkmrFn7iwOodv8Hz2ogYhDwf/PunM4lESJriWUdDj
rZ2skH5Pl0hZrs0dmvdatTVNv2umGPfdUfaqqpNoOwndVG1uBnV1gtbquLRSBCPy
Pk7gncs8cAQA3yRG4YoEaYOQW4tMYr5qpVxlnXxRMfh3NFRuWT1JY8BYyDkm1Rzh
Lh22QJxhbd1XVv5sbEm4f2DHJG37x7wu+Qvxekv1uM8PwAskQHSWVG4LgOmM0M56
JOeX4zU5IloV0usiJIVgxbH5//ZKiMHsJnTDpmp2CFLyT33mo9ws0CaUKPr+2y5w
c2vLRIyOPzWH9q/DAVvrIpC4ehNWxNNy0VZp9yrE7JFKbnC9jOcgdZZ6J1lzZcKO
L5gMcQaMLvvODbTQ/7yRDQJwUgskJW6vpMec5Qa0/uNQ1yKqL7xIEpZJLoItoHQ6
lUfB5nn4MftB5FRc3h5QbSiPb0AolCYi+Hqcrgw3B6AynerfGgrlWaTd060XPJZT
BdiJPpXJ9gSzuZPhEfP/N9qoVq1D/HxZnxhGQzaR50QkhzPKxrPkHX9Lcm34njbP
nzXWo2UyOjNQnjQv0vkZu8JhIPsQF8njEkjJcwig9qT0GUqrAkeIjJ4DHU3qGaYH
USgU/3xmBU91fyTXHZm3bzGcG41RvAXijZcmcX2WoxO0LmNK3B9Mqs7v1HvQ3+fA
PbkbDNKmI94Vdz++p5ZUCzsa/bcBzT2vCyzaZAni0xxqpDztW7rPkRZB+gACjnNi
SN2bBxz8rRXgC5mu/uSnIGGWt2vFllaRvqaEs1H5szA+dNWmDzBoRUQHDocI+3m8
cnpYUAXsVyJxCy/KlHuVxj0E419RBn2VgC3G0dFsN08ps9pEmpnzypJO0aawdh5w
rQOEePMcfLJ7L416kQH2byVrM6tBba1W9hawPUejyYb7qxl3IQItx2sgMFlTr4hC
Y+NGx6R7SKQMzIxoove6cyg3n+RVMg97ACiM9WlE0l0jIudjKoE4s2SLP2KpkYE7
BqcBoOPLHHURHG7l2/R/eqophXZsBuHSHj0Fl2iiiXBtnBXl4fe6PIQJvwPkK1og
sgy6m6SQAq3RXgOCPhiLC081ge80M5qEQCM4n5dz1MBd5adXNhIv0KRTofALiCSs
EmbiaFMS+ZzsPxf8JVP4NA8MDfGCFPIhMjwmCJcg2uuo935wtZUFtd66Kp8nb5oV
n7gdSNJoY/LqiATNT2HGw0RNK5UDDehRsQF1+J/YwGiQlZ59fCkt4XTuGgm34pZe
drySMelvi1TLdLfY2JSQMOqzO6QSWRA/pBfbXPrnWzSfdfn9Hmz0asBhnMrrZCjz
c3zIvPsNpZcsDSQ6AejyEH2LjWff3KzzEYyNy8i8R9YUAn539p3pvqpp3nJcxHqT
6h4anj2Xa0wqFJBU2sC3aKiIHxcJjPVf7BNLpQYKT5i/9+HECUbJpcdGStzU1198
fSZy9e2syECG8A4SP8MIqxrsvFH9QKpi7EYsrzH4j8ELcNMKc8i0eh6udQjaGTIQ
uOhjYvBADEhUuv9EQ/3CXbRhhpB7mEbOPnZf88vxtItJ+ZFlij14DIivVV0aabyC
EnhSCWeV+J/oiVBhr0s0IiM+iYRfJFSeBLMPHtOo9AutP7he/KJcG2TelhT43jb0
bvlFxmTq3SIf0oiOiiKe9XlATMbQ9bFFXxNywGInzkPMZe9sVqzTzX2ivESqZsWR
+Utc0AUgyHIfHj9Cp/x4OPLyxfTXK4ideBU+brHMR6OZ3UVbfaIOiP7tQ0uRe20X
r+p6d5QId4w3FK9rVrCtQnWhr05aqFbecC2uA5Iod4nEWxm3TwFiW//zlM8QGUtM
p6IzdoWqp9yyRd4J1QPA84RQXbVkfd7ywzFW+5B9spjUQE2ntGEkoX4Y90AwTOAg
wWVGPDu1Cmr9r7Lq1qiN4Ut90zprm4dFbqKuAWlN83kQIgX3LasYvER0h76fd6YC
2DpG2W3Nad32t+qhwf3u9hO3eW8vPSmWaTPmxvdT392AWspHIKyqJdLmzJgNofYi
ZPEiAxUU4FW8tzWA7KiH68IMpP9NsAbJgtJ91kQp3ojul8rBygiLxYtlPb8ewxyO
kvQFF7RRkO+fVb7XdwDzUPZvhiQqyfBHH/vk5LhPALPZkebM63EButWBewC2GsFx
gVfNvw6W6KeIpTKf5y0HISBJy8oxclM6xfJjNIQ10gchIjuHtI4xJdSeQ/UeQlww
syw4IWtA9Vz0nwmAxqkiBrqRaOOSfD9SPN7OtZVu6bx6bvy32xH4yQHeB4YlSBbH
wUU95GjJYVvJvHeQ8updWUkVJiGDlJkSATzOiC6yq5vEzcSwyfehoqXFACTdJwWc
GG+3HkcnYZkMdP7OBRzsc8W/hYY0DnBF+djUPxTtOB9qYdjwDPizjw42EqgaxCeX
MAcCywxs7YLCOrbFdWkzO1heoIVCFxCUXGMWYiklyrqSrUCktOAmL7xF8XrvoU7v
dBTLr3aKgCeRZ9Siu1Sdl3+YltsiuDgIT5QtX/pAc0YbAKq37GcJSldPab6/SAA4
30G6VgZCsRSMAdM1dEgR+Ekfxeb2QJyHggvHpuqaBJqty00qYY3jFf8tViNmMR9m
d2RQQ6ikt7wtrf1yNFBTueoO1zxl3Q+HKFN657gxIwaA80d1iIjPTINldbxtI7ol
XtYQR3Wr01XGuy0ddqIAp6HrZv5rSWtY+y1km0g69aVcv3AEEsxWSzWUqVr/33rQ
P/IPFeJiEEl+W036ndfYIQ+X2qd/+syk5ZcHbGOu0/JSLJPCrQfA3O8mSwpvuOH2
X/SiVW+0MSNnSIBk4dTnDi2w5tRhO5IR2SOvadUs2NiEYYGs/X/xbIJmkgFBuD41
gmJHqqSZCTUilVH9uZ7qhkL/6KQbS3IS6r+aJ/VUjZV7pAZo0gSeXKvZX5rBoHjI
9ar+WqmHn/VHvQlpx6Hi1WpQpfWZQNhNo64CPxS3s2ZbUf7Rt6CG8V+IKmgMeMwL
xdhgl3Ik+wazWdAQTYg5CvFkDtb5T+V90mtz7S0x/NVzFmwhCJ40rZcaXfA0jTmv
73vBmbXdS7Qtiqknc5f+T0yz1teh4AGqvf6pJZP5Opa1nj3l3dvR2QegeBvRmldK
MSwrQXKmfqyxWZ5LMjHkVsxgFJ4WtbUlpvASTc2/5KwWB7r2rIw2wl14W3GICzlW
+/Q2kdmVxVg8HXmd674gw6I1chHxbcbVHziUuSO+8Q/SyxWx4MWhGYu3gW5earZz
tYaezR3TAOuKl/S26Ef7pq4X06uCQo7baXn3Jx+hJKfs3BfrvBeHfdvu5Q/x3xm5
SgxSfFr8NsoqAbcSoIjMh5EZW50SFXSkr9IuPgT1ClkatFygIl5N3OQwID10LY6p
maZ/CsOnmK51k9WT8zpqkCELf3VCFc8M934ERS0cwGPkzQxDd7dha1rWkPPdgnSv
a8iE2B8EVqXxZewDfAn1zwamdWsImyW7i/w7X/wz1SKs0JoZL90pPaYbucyvNIs5
rrCCSPIXbOjn4qclan/vAO7j7C1I+bnyZ4XvSFrzYtR/jpfxWfu3JO2R0hdn541R
S+8FVxmw+ERrvQlpLLo8nePVMcr6bVo75nzhv8p6o12EDJYvXVnhm/A2AKP5Nq0Q
N72MQKAQ17PLx+hAuN+oH7Usb16F/Qb5BYpHJUKTbb9rD01JSC03nMO5SNATFGVN
hPZ0emoKPbqfTfst/RbRgP6G+477zKX+ntKJ7lxJ0wXUe+N7zPUm8Uw5b5k0q9vq
Sa7xbJqQyiGNxAMownrQWJsITfte6SnFYyET0Uksife6Ks2RMbvOr2VmAwUEXdEw
uJ1YdKNK/eFUKpcoCpUZyQqW2MJU+wQolBMZ7gY5yEAlxkOaCytnLM4mBSw7l6OD
RdgCrGA2ZxeyYLNEKbWgCWT0r9fy02IO0IoEsDAuWaky8tzNoA0n6IJyRV2mv0ng
krj1X7ZKGN4GgAOuhfqH0G1EeIwENP1OspLy1UcPMOPkkkd8DfEYcrcQI+a8Og4i
0NM5SCfkb5Pywjy603ZduANBH6MuFdlWnftfSwfbQqPnkhDTbDopAOIz2FcaLgOc
yEHMFTVCpjykQaJyqTdAPhvFat5NfNEGXytvFn8UMy68coXdXGUX6glny8fthznh
ndknM9CoArXSZkakU++NlCBNfEOR1dqbvJ6ayghTb1h4Jezp5j5zBm0hBxcvmHn3
7k4rW3SXjyHHO3mCKtC6lorWNw6pw/PU3fa90JhVheOsSd/6KbCgq7tNUjyfVp6I
1un634u5PILpzRfOzJkGOe0itX1kml6zlGbz7wzTpVLkw4yAp0MMdt+V9LAuqWl/
W8MErUJwsu2KkAYWF+U1FjH2nnWy5urdPvumH3h+XkEwjKq0OHUPTxhPU0zSWD8V
aI8LBEIpfFbCch5G9WhEUdIHa/WJTvXgOozPRAhlvfTF63ToNUrBV7tPDI0PZcv5
FBdzGve7VEM86hsV/QXaH87/RVhnqlxGutJ9IT+7W7EMcSEL86x9YkBhCW+DgmME
73my/iMRhyKUw2ZNSCBP/A5T0oGptLWT68di5kTxhBGK1z3svw8sjmQBOq/RwfHx
79OlXa/Bg3o/8xiDnbrJGRwbLvbEhxUq/r4a8HQa1XbBec2Q9VjurOXCxXHFI8uh
x9+iMDBjWHvQaHdx6R2pDBHzo5RFGJpVu57DpwjiV4NWB4Vv9R65aL9B8VN5J/KL
EilTTd840g+eELjefKA+VoG7whx4/s10YqWu3PSKWLcmnV352DcVl/cwiIo9bLJO
HMRFmhUnZ6ZNtwvaImJMNnaygee4lsdwa7sxEjeav+1detmoTfR7/dm3sPcxYBIp
0cZOtZpb0aI9kuEy0SEuXIZdbcPb4rdmA0a0LbSYD1xy7A/rggfUeB5GgZ+d/Tb9
A+SVTjXUygjSLt+P1GstPXwIkIwCG8IfU9AKIsHvAD19uJUR1YTymP6HZw4RSuJ7
nge3cOWlVHWVKv55vZEP5ZZVUernM61Bo2I4uK8Z83uirLoBd6V9/FJR31yFHZE5
9qm0B78c+8lXno8M3YsMt3Bkcc0FZXLSR+/ljPIm1mpCHo37OnZU6PcB17z5RwBw
4j/xgapys5KP8n9FP8+PIzJindQXFmV7+h0lnknLvpJNhbUpCKxOKDE6PaLOxa6J
renQBMKVmsC8lfdlc5Y6yXfE6MaGiPhaBZ8jrTxTfsSxy5JCBvqlBXnvvbqgVC+U
02CVSngNWu0mEE+m/GtYe25b3klJ21EVXqEw1QVCDDyQpZw1uAQGPG6tWihlopXO
NmUo+H4gFQoCllIeX7ZW1Ip2p5p5cTQosKHPnVw04ylIMC1A9wwOXoU9nKSBsQtK
SfYf9wjzeUizFzRxemKr5R1j/gtUpAd2VBkrDs7Dt0fxLuMVILAeHVDP7YbVwr99
ZSUw1ZK3S4xQwneoURrFNFzG75w7FKJ0jghytIR2o8I8RFDiIHHlYF8z8IrvkHBb
BbyZvP+sZVJ+88ZxEWgfQZe2CgzbG4HXj4opume9AiVrvKNBmxLJ4eezpHF/quN+
xHbGLFD2zS26AAjZ9I1uZKXXncUN6n5yPXfxj9Rh2Th4Bco2nbXtHwQ7ncg+h5U+
JoLRj6Kmq39fadGn/OfZaifej6LRsO8IpU41z7MFSK6U2qGKbm5L8jdMIS14RO9/
Z9eiELZnJXoA3rwi8rUT4HhejdTNMmwTcagePMQw6KXOX35lZdCyFYbSERPHw4Ed
SMHTTe6S0WHKQoMe4PWUUbp5JEYG59CHSe7e9/OhgUdx5TXIMLapjqFMY3ih3VTP
NzO7xcGtx86EUM4MDf8hqF3KfzFfDRf/A03fCzqeSFNyjFJ3xcYUwVqBK/XiAPLl
pqg1ALipoo0MO51JnyGMV0xpzpVPslMxrWIZFHNT5VDZCBJNodJF4Oy7qdblvzdO
Vdih8Kja/Pbt3Hk6LWOajaCKnIwz8wkxopy9qaXD6SSGNGlVPjCWWPvtDuvEYwZJ
dvlR0I7lcL+2NGemPeSudgcoDPAtLT9JR2f0St17JC34ViHWUp+nfYIiJTKu69+s
7YVB2PeOA4ZTo5bX1s6RMRRjfDgl5IQt/haK8fmOHLZA6HSvi7QWJ21PlBGip95S
M5mInm+Y6N4jZQ597+1dCkXiamvCVm1AsQVrOvAQccFUUl17ZUVLLXF4FG4gEOf1
FTCnLbkGs7gXLKncP6POwIEybITXWkXgwcvIjx4Qs6bkcnn7Uv7cWCPb4QVsJUrP
xbvjoq8ilFsyaZfWCXh8JhFQDj7ZqacuHOp2o8RUL/GRDQ/D/Fcaqah87/zSBJWw
OvKaDtEYkn/g1uhZNayyQzBtjSP7kuc4ckIbM0Z5RFaTbSu880TgiT/YpOr61Mkd
pUYyx5vNmAgPNZOmYXyyhy4H2rn6cwSVKj2zj8Sdc44dJs04GmD7/Rg8x+FAUEoG
RR90ODiKJsi+0a4h+tT8AEQ8rUU5ePGf65caug8d0A7MVIuHa33PUx2S9iJHd/JH
RozMbRp9Uekdu9ZBm96idiMSm5sRNokIGhKmPgMIoovWM/voOJaTM5/QINpSlzvI
WWQnaXHH45GynwMNUoH+ooxe1sc6zAf6KVWoqSYWH9elMKEW+ciTqunzNFd/kaXn
gRBUVn7p5K2gNWY0gvQ0Ifqr7zQx4YxpzyMzogvGcRvafdJlDBrJJbFYDwd3fx8i
cZtpn52/2bgcZXvg3AmWXumTDG7NSBnov+GhvM9gKASuhe2sjj52DxM9ObKjEVvJ
ITBzzHtzynXaFtNRM40ylmsek9zsW3vzzLDx7rv+cilM0GOT5EttfINUe3vtTcyd
8jq+RcbakACqzSPz99Ejh5BKm7cSeSRoS61N0vhG2K0eZi4ANItAxcYBKVG1RVdP
kCpGzKIp8NxZDJwA1XwQ2W8qBDBt2E1NAR2Q8Z1JjLRximBk6xyGzni9J3QE0cD1
vtbu1ZSmc8PQO1BBAu04zZlU9E/eHdvkC6GkmAEZNzx9fWyKj+mETGiEPEZ+sJf7
szfZYepJiVhdYr45HEMO9gbnoZITEBen8BBjfoV6jJuACBVAlGkhL7MU3+KKW8NW
TEIlbzUsxH/L4gULVxka7yHIG71DbjElIT20aZw1GeCmGC8GXL6zUlO2EgOr0az2
hiaCYDdNwZL6odUDQHvMlp0m5YcTNRAIgJ/J/BjHGoc6CfTa10KNyfSIJJC13BXX
mbXvYt2GGedENbBbonp1zmmIIT4SGedMeHNsNWS67OQ24hNIKzAwGxmbjNjolrvb
dCu2CaI34+8OdCWWtgVWQLVccwwtEpe0xxVcZVS+M+hITwUvCsLp0nhPhY1LDeDt
7KIHGs+ABrI8edNOqQv5pUCD2u9Mumv+H7xgIo18V/jBn5wmsHNNPwodGXe3YIDq
zJgb9upXd0xxtm3p86WWHbSbuAnkx+4T5TexxlX00z3Ag1m1H+BeQ4+4FAgzL5Bz
cxN25A2MAy9uYgDRxon25p+6MF/h08+u3yrU+tPtYZ+jXhkpwBWCnY3w8J2C1Q6j
GQWt6KSa+Wv+g4TL2Xh6ENkQ5S+NDutNJ+0c6tzgNHsKY1WYneEYalsWVXDIUEWP
VLT+K6769ktVWMHGfLEkeC+8wLEDgjFMKEhmiJtcXjEIsQzX3/5Fd7b6dGBy6CY3
wy/fH661bOGSRNQ4BdKsSDorSDe/uWFPvkEHzDZdh79+X6nChxMr6kW1TtAzsy0i
MBsg55EpPpSKgcjySAmzpP/ZLXKuzb2E2d/XMDMHE7n/JvTOE0oi/j6iIlmqF8X2
f6ysDce7GBthfs7dj+FHWAt+ZeHV3OwJ/g5SishX1CPfbAg/ek7KxtGagdgiCQ2i
UhWD7l/bxOJOp0VEpS4pjtjAvuHKAovbFaFR2DoToS1ID80T0aIV04whveFOx/Xf
tz85Uke0VKe3NtW7QLMzp0xRH+KKTuoXw0MYNZ+lafN/iarVfuL+/f5vyaM0rKig
BXlBLwSohL2S4J6nO2X3qUPx34Nn9b7MA/huiZZrhXR6VOdXhimGMvp/YkrC5onn
cDtkRcAtSMldS2lvJdOJw3LStrhXo3ujPf0wSRfq0YE8IjJ8HAqpHb/5RI2ygYJq
F8xFoJ/tyGtwY3VWTlNiXT0Vu0X/hjhxHO2CpNSPxMtoc4wgDyWE/EqkKLwHRrG/
/wRcGObP8DwzNU+HfgkMWPSRbh0COUsZH3dE0GRE2Qkq1OugrjvV63XpQ5EjolvB
T7pd4yc4HbmKqzP0ifTrd5L/ccj6+uuuXLiXNPNWh3xa48pHFVstsxNY27kMTp7N
nlrrsiDO/mJktb09QeMFIddu8bZyi2wSLo1aNNGrVP2ZX6go88guvD//6gUSBzvg
TZhB40k/vwZPKG7sQ4sVXXgcgrjEullPpq6aVQ9W1WxDrXlgY03bm8j+wbEyuA6f
2f0Zzr/z1DHrxQ7JQ/Z5LhCssqAZxReMbUOOgvLCW00sNYYzWhwOY2xEqbvXKBP6
0Vwf4duEvPq9rie1HojmRbUgM0uNcxXo144Q3S1u9224ufw+BtsyCxF+PEiQi3PZ
hmaTx5ETWUN5kvomCvSaN18gdwb/AZ9/jBZPDBCD9e1I4vwDgjhhU23CimNqd8l9
rLgHYFQ5PlTREo9Sju2dsUnyOIuOXpa4pG9pDp8mb0i8NIcb8Uu7G6xlBCje+kyN
ceyN18tgTwfBE2CunQAK7khqw3mkVDwbCCt5PbC41MDHublJDVBLJz0vootx83fQ
wzIQPr8gAlkl3LX4dGtlF39kpWG9N6MxI7kqmOaRAAUWt78RT5aAe1Uk2RtNubXw
WLba6Bdhbl9yqENjWxiDr90nDMlFO4bKBK8mJS+4DqjYceGsQ6hFcN+tQxkOI/8I
rRzNxxxP15b+5IaEMfY7djvwDMqLCKJQ1YjFA6koteke2vi5jJEfBg2BXy6hsosq
vqfh7Wbv/fmrIFRQctDB9OSEzMkbQDSyDotrD7cH1ygq8Z+BIw5hq5lnD/YPc/Iz
38qm9H+hYTmfG5msB4AsflpjuOtNTpNPTJuATSREKixWCFoQ2u9/vO4ziQQdCgP8
2k/1rPLC2Zfnqc6YMxllzxMldYSa3/D4WEsDRXfMWPJUgaK1nfhWYGTBtJsZl1C7
jelZ76rGpYuYnzz0H7OVpFo/Ji4zqZri/OLO7X/y7JM5UDOJY4lK41bRQdnul5FO
aDnGfu5Oh/MOh0luiKXNs/GOCI2YaiHgCFnBADQFG3mwIciIursKVG5B8PZnbAvA
9OzV84oYWoztyq2c3O57Vc8RD7bwyjcRhWgef6dGnGm+sMOFKJiBST6iFilCa2sQ
O2MpSe3oGbrsx3uxoIGRFhnkoDcEjC+X4mx4IzfzuCpQkJl1ElRdASK1kKNNIh/w
jyad1rDwkTe6/6v+efuzzqCE80mqsrQxDaRDU9XcJF6+4tBZfSwpgfcvgun+IntF
iaNjEbnV8P+hIvahI7T8FxPdI+JzwNULIwq9Dod/1cMM7OE3ffPokWHsvT5EABbd
eO7fJyY7TT2Wt8+U6E73DEzz/tSsNBwsyCyvhUMO+9oFqdaq/hV9rZSruNAJvPDp
sN4PiIq8+DijP9TxHKw29YguIL/LeWuJcrY8kOsAxl+CG2jJ3inc5T15jKn9fEbo
3Nwpqa4YN0G78STl7VBHXJhhT6x+CFJR7kwuGLL/s4Ly1RarKkVYKSWmaAu4wO3x
PxYBqfLzgSakvgPp6lKw5GL3SPqlPVvYqoaVECYyTYWUmA5sifV0KvjuBwACuITu
d22kAuUWuXPKHioDv7e33Eg+9C0PQW+7TuuyKUtvsAY3/nZvVEQUWELm1Jtg1tl0
5bf7IkVQh09XG3xIKxcAjVzXW8YSDpX4rL43sgy05OmvN1Ah7WkBtpKY22QvvUK2
5FHS84TdASEa5SZFVqD+Y5ukW/9IfTs9HwA77EYm+abZVTteb0ID5/4HDj8JqHoq
SyXP1rkdkt847EwkAMQ2lMwRW7SuAJccpnkqu7IygkWqxX94qamaWoMJ9vL/GswG
NeaVe7QCbePuLjq2Hj6Hdz8EELc/7oB+G5jkygP/TNGH74SeqYUpB+hcrXy5G5uX
+scEJvRsDQ5Iel6Qb0k0I9qvgbV3jJ7Q8rIfbm02aW82AqygwmKopZrQZgb3jfwL
0sICsByZbQ/6o09lPRWeljMHxQFCppWjmtOdrVoYxgxK80fTKSLG5jwUckF9sVFj
XpugleeqYMAzK+DlANig03Oy6Hy6NSKUqTWwqcrjwuNcSoAqfa3WlK0gGnKuiRZL
LBeTpARf4dRocFeA1th85C5qKHYT9CaKWZyrbNfViTqR7cssLDTbAmHXwcyUH0XB
umINsZVbwlSRFQcIj5XwHFP7Y8SQetgc1R8jxcxkxs/56vk8L91uoc3a89B+Q2Wo
KUfbujKvrRgkTdUgxR0WsetlkEIebz+QxNgWeygt95M5GRVEwxMfgDpFOAyVp+Gp
ir5pFuzVtkCGsuP6oGEt+SbnadMfgy1bdPVxpt1KMidupM2jsi3c5w9KpFhQNDjv
uYlzakM/PcrlDztruZm5dZ5WqkHyVnepNXUIMgiamGsaPoQXP24HhF5xtgclrANM
JxFZlgTN2gtk1yv2RoNDUVcrqW1I5tV4My9gbPK8A63Ee5o41tAmCfVGenWH11qm
fL+pyiolGNUVHBumjRFMos1+Ouoaa5TJq8DdeSxNqMaWjJafr8IUx0Z49NpZAsy/
RWW7Q2YE+uFWGuz6KJ0NZipzzDPm8kxtynpRtj6VCdjg1SPpoMzizG5/B2Fcea8K
7QrsEnRh4wKXaUe0L9G5i1vlPrU0QbkfpC+eeOwHLrytrNt3tbr+PErgJVodc69F
hcJ3uZRR31SJQz4roGntCZ2tGGRr7yoyW3aHE4fFr1Bq6SPDSrdetDrHDrtWibp8
bttpo9sutiBWFkS11nIc86p1Ssbt+hGtJvYKr6XimFJs01GPNp97WWrv3O0QNQ9a
Hr6WmvSUjmsh5dc+v4DbQiFK1icqiLm1XZbWsViRQyk3Chp42jXYLBXqEAHyUs+2
K3PLafiT/a34uA9ST+nm7mR7BmI1TcDDE15AgWjR52lvcFLDZ51AjzQVBLHjZRRq
w9x1/TkqUqF81ZRHV4CQjcb/7j/SLqA9FyHHGIrEVq2YgJ+3jy0mgr1/FrYYrjWx
Cgyuauzl8Ss5GMgmPukz7M2MlqxmrHDWmdDv5B6iMiLdus65Uc1F8xRizsq84kfL
BvO6zWwSjQNbV2z9ZNtq4P2/GUk0+Wfj5wkhbu+z6KBa6ESywsG2MpjBrZk+Qys9
608TzxPRBv3NkQ89Nis/CnD8TYtoqa7/ACpFmleiJbLmmvBy54Ssj0fGjC7rIpZs
UxiBywlSaKFYJalsjP2uJV5/VoBINeJ8qhV7u5ieJKqJt7DAMZQZKvZF/3M3IUq2
JeqIiQNG3XRgqsyGaPO3D/h6I+Xh/xcTDINUUNyylIDUlmd/s4YHiPOfq4riq7Fg
5G/XFmRXZK0rejUflQqkA/e+zX6qGoOdA8JqqvThYLMVO3cNs//BzUT/n+0JEUTF
TgibU59tEHpmWN5zivL5V/ebV8bu/J51Lv1AmvGkXOEw4hIWvNeOKVPRUZ3QSLs2
OxSRjECHX4ojbq6K9foYYlQzWT0XTQH6tpYjX2HGZOMfoTsJpwqhs3LKxKLjfngh
Jxi5hmWZp+orBTKpkiH72Q==
`protect END_PROTECTED
