`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VcLNUV6l1epRFlqBSUmNUXnl+QsfyFl/BPZyde4Xl7GjFzqA+C6+ColgNAOuJChI
qtkLZM5HuKmY7Rs0/yrqDbSrpDfhku0FCx9gpFXMZGWR5BuonTALtVmaG39GpBsV
Ld+gmJEK1Yd5uyNDpw8cC427G53orjr1C27F64z7oR9MXUBSt568FIAX2ddeLse4
yORqAGzWk7DXirbGDXqTWDk4GdBSYdsipj8g/59X8BM9Xq/HN78qw1bIgfJzz7/Z
Qgr4qIQyeGHWz/sH2QxU383k/FbYvM+pVSSvxkP+h3k6Xi22iqDN3ZE0gPEdnyRA
sOex3Id+KrIMK6oeSTxr9VcUngOVPA62ulZomCR+0f3Wro6loPit2YEGzVl5OSjb
xHujmkYJ1axMisqGznNkSRoDUq3yk2rNEqQ5J0D9yGEGC/2ZFpp2Q0B2DuF+Dlx+
uuf28waZnBgqu+PCjql2+AxX/3EIS6PkhQC71+vh9pS+799VmChbduw5hybD7bI9
67oLph2xgXtUNKkDoxONJersDB5CwZnM6GavCj9vwHbwU2GZ9/TAKk0VODmIO4I8
nK6XriTedkF8+yip9syYiQUW8tCH5E+yVD4SuWYc4bo1Db1MOrtstlsq5QoY9beP
VrTPJODZUzOUiou00eoVFXAhN9uUs8vofKOEZoUN8PLkPtIFkeZvvUQMhQScgX3l
QTFedHMtt/5Y1mErsA9Q7kuosAIGAOwva26agfaSOPMBs0cprpJ6cP7xs29yHHu2
wZHtD84B6rOf/uyoJ4ug6A9yCDZ9aJThPn6bdRuw3DB5s35yo9yvtVDKp1Wd82Bu
G08AldtcS3jJvGeJTQymdk28T+thLchtCnSjA8y4CKM42FM4J9BD+UulWLDMrRLL
OpLjPd3ra5oN/oF+dfqW6fZFrONOAKXiSF0bPpmHCJcWv1hRyqRhpfuwKmDeIRnO
Qa+1N7/zJNDYuFg0HKTzroku4Rk6M6FGPY6wwnhMksXsPDcVi+Ip6Naz7vLG5jXW
hqihyJnh7QV2UEKyxAVDC28hHW8scVH39h8KRLKVHIvNqO1D5ZzTmkwVZRRsKLWN
PMEufOFh8nIDovSra7b08EtVWHkcbU6zpJlOSMdC1u27gtr61cW9O4+ZowZJCqmV
vc8/RBgiArbNZfpH8IqoWfZODpfeSTqHj8iqpmJhXAPf+fZetgpXpx0M6031BSqy
i5qMHngnUnMEOSX7c/ARAR83LMhhbIKg0+jgdIs/Mf+e6nz2yXhmMsWS6lix0OGp
BuywyNrJBTtmbfy8sxbO6qbm4GjMkbOJpIwX9TwLI/rX+qKuTfKBn/URy2xTp/Lx
4rHMzJFhiyZVDe3YoCV1gVQwN9Lh7gpAyZNSHo3Ul9d7otnI3eZHgAT+gGan6uKZ
Q9j9UGKTO/9d7Ys90d86MAQXISjcPNOuarGk0WIXcqE7rwJVHTvzeP1b7yrlNtN0
zfRGczEeq4raG39YPl3jX7eloX9CulfzVmj37Ct1yWD5OOTBV7zKcPvQVxQ0sw55
`protect END_PROTECTED
