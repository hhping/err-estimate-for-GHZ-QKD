`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nWyagNwyXY9iEZ/mUyUxetzPr2Z264qNCAnpV1PmGu9wfYBv7BFAw6hd59cl7Vy
jROmDuunfprtorf6lXxvs+DVcJKSwYpHxYY8kki8EVp7kzB09LEsKz3uRQZF0kZO
lyzEPr/836auporsNd12borN8CSoMEWJH6ybyuHs33urxUqxl+2FMyeaRek9ojP1
DgpW4btO9lXgMOo/BWwlE7EbPPVa/WLILBhx7BhkQ/VNFDwtI5CT8Ak/QTWqFXma
/iTl2qmyBMcYojdJjMBENJaXoXaP8MBi4aTLkt80ZHpLBU3vNMSdAjLfjbwP//eC
OaSD5y4WxWG63+oKHcvQgUcfoT7lKfFnyfBItsb7tTg6eYpT4n4wq8ZN6G1CkP8z
rXUbwtfvUK8z1xusHKoPx/qoW6zd13pVPhfC74ZWjtPGlS3nhVx0JMzCBMDpxK5B
9We/NZp3jGTD/+FgB1Yg0PlQQUXPvaal/bjKsqiVGRKsA+4KM+0BPLZXvqKTQWY4
RWjaKCRS0HEvz1jiXJYyat0/8bSz87OOQOpe1t5+jFJA+AMDItPH0nchJgnXQakG
ngwIly95xcKaNTj+7t91TZJPKKGl8D6fmGsFNjcJRDhm4KtnBhfaroepntCIAenB
FmXk1o92d16Ds6JcMPDuPjqva/hUTdfWMScYwVoNAH/ZgvSn7HfPDT1gx8hODjbH
BW7bXGZLcPRfuK4qpGWBnBIFmmhn1RfMaCi7snLnw36SxRJu42+WADYPwx/LSJY9
oFZK5VRRNS2Y3xvBJo0PUUYp94jliDd3HuS4DxAWs9FnMq+IEv3Ga3aUSTteedPk
ACqAdHqVnEeE/xlUMxmj3Sukx6CI+Te8xqZ8zn0QyvhnbVlUYdpjjy4Hjkmo1/Hg
la5zPr5ruXxQNzJmfywbtMgzWDx8iT98XC0c53/YU5JiHcNEjGIBUAeN8jOL+lhU
pqF3JEOKcXGVQ622SQLH1nspoXyETy183BT2Bn6zZO1OIC0ZP5weP/0WyYB2CCLu
hQKXkDp2383DV1f2YJPysUyrQ2hvT5RphqyZ9nrxDWswiMYOAV7+MegIooRNs1Xz
I0zZXUfmhn/7WNDzKpuFr0iXFI/kX6SvAvckzulvt6GVhk21xZRrDhqdr8SW9q3w
Tmsp4Pf0yuJ99Sgaik66VtwHNtreF0S3tBmqPutOIkgijQy9r1htGcxVFcYsgz4I
Wod31pqWkxjv/2D9yyNKMFKHTAiVbM87RcUcydiEgaE=
`protect END_PROTECTED
