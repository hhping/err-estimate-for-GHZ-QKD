`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QhaccYuwpRqI6vEYJ1XIPhXiHVsBwYpvul5aXYXqTiaCfQBi0ubvFiWfMLxiNBI9
knMKpsPlt54d/HeYEejs+MIgUqb3+DBmBIe5Tm6fBqvMQBO5ZVzuo2ndbnUMRXRC
/pYI94XbfLQjvntm9O9Ioi/7UWI2Z9hyclrt6wxQmmrIxWhI2foECxxxt/WPOO0b
sfqnyqyDB8QZAfDbfj+UlrWQLpgVB0uVKZZq/2rqLN+7wfZlsXXas/VZ+r62AEQZ
7XDSN6HynjBj8GcU5Hb98rvq9FMpJ+ENF8EIYw+fZbNV7aOdbZBF/I+3sXD4XTof
lj4PVCLIdw/noCoKDE5TbHSN3dRV6zsf8J+K5xkcfy1Z9jK2A0uY1irG7vosclA6
517OlNNg5YK4P4cdQKOgArWtwr5JBMTCeC7AaOhhfNRapaVGkrXfycmtkcKs2U5c
RvD5gp5FhSnbW378haSHxLRWo1JOqJ2SMIMei0U2/kK8Ej5w7vNKR7TofTb3mIpV
U7Q/ly4iF1k13GvxSMRPx34oZrECaboyPKCdhpPrQdAlv0V/4+S9Rufo11TGD+KZ
+gmh5ka4R7Lj6Ek4opqdt7JhpB23V8RxudQvGFbFuVBrTO1BNZmO72sZ0bq6DQ7J
QzQXmBeZjI/s6KPjdbtiP3LtwM+rbJ9NbkyGmg4wBVk=
`protect END_PROTECTED
