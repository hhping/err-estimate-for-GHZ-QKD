`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgpiXJsGGKHHvFg0Qo4W/kaUd5+8ZUyWH+QUc4np6fN0oJY14YO188NCl/gvYf/K
T60Rj6ADiwimlbyDfKE3OQrpUhZR2KikQLfuIPx5A0/kKXcypR05/T/DbvA6RnkK
24aR1Ly6lLvAPCvPRqxdDfEI8hDg89yyzWCCGLMNHo4LYJeUGEFq5LyykDGxjv3E
culCMuFpvNNfhfFZ5YYHKXGWs28g+ObEMdNkPlwfKaKLXtfJXpZrTPXJwjn1nYc6
EC8q+ZFI/0Bh8bPNxfc0kyt9guMhNZSPW9mnmpSjsm5Mpmeb+J7/tkoMioGvIB2Q
NfllJxv9UNKluN2L7e32mr6wwTFnFacTqmruAF/e+XQK8xhWFpIp84lCusc1046I
ZLWO/PraEyaaS4CEApb87EsFBr6CMGj2d3jplQ+K/C4V/oT3ghu2Cx/MXm71BSoB
8H7hqwbpDwCuEJPtLRpUMgSoj+CugXkHtHyTUNMphaUB9vmkdE3Ng3L8iWBj0015
AtlySyT0B/7c0c4dZKW2GCs3Yzfuzn62rvLI+CGoxAS9iSWRgSp9gjMWPmcO8vPm
jSctPPzsXUewVIWjecEwlIcwgg2OW3kEmO8CpuW2cLoIPbIOkSt9914QLSHVQl4O
/AQS4ps65NrfJMT5HO1t67GWI1haOKf/x8sd007+jVachze78EgYqi70yxZXkAaa
n/B1zpg0qz6byttZOXk1nu2Y/UhnvRLeXLX+pWp++NlNc3sKdkHKcqjU85FROqJw
SmoVAgkEI42QlUjGtXVO0dgfFg0xcnqBUKlJnBwNuhHbz0YPKmkclhamXDty58Tb
dqU/jozpRQnEzeZS41BtX3esc3xuSq3IPqFnZVGl8uOpF1eMFeJVnVDXNiJReWYJ
+sXeHlXrZV9IP+k7kpdVq0s1H3jwyVQ/FfOLDX79jdvvILAyM+qtkLaTy27uAbLe
GeyYdRxtSDf+UI3Bb9kyeJSNLB+voujRoFpLNqx0Pw77dkOGGiORpfGCu2iAUyQy
98OrunVONDTN74K4s7wiKxsU478m7NiQQRmq/gGeGQ8pT5ENxyt6V0hFS0OPQVQq
MrvihfUli1b6iYTjwus6m3penkn27apVq/dUU9XIv9OWRTH37m9Qe5yPK8BtvZJ2
gskN3rsF3ltoXYLKmhTtR1BImcMoIEkwVy3csMINqpgjlu3/EaiSHqgTkuHTmyda
WJ9iDX8ECyyoGEJERUqfZzHabHHiniRYx0iotoxS14tTnhL6S7aHMDMc8+zihtrW
OmZOF3Wkw9nT/dTNUGHESg==
`protect END_PROTECTED
