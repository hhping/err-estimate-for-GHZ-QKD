`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdwIvB4WT+LAb/qS1Nh7hZUDo8KokgTSbid1Ww/uS9JDtDbG8HqgLmvA+zAKHw+n
d+dxvz92oQWznttaDIjZPOMIRG4rJyc0qvnD90oubOmPKg0ujltqPwEH3Hii9Mnb
kw8ekCV0Tki1x82mwxiA3Vx88t9h2StlXCxKSd+gdeJzOrYK04rUvNTZ+ZTDufsT
F7TaWmIC4p6C7du05i+1hdkvHGeAHUZW1pWiMaS4d/q8pTozoX5/fp7wQsiB4Lla
8s2DhhnU8USRcfEzCeNIUKJxk3RZOrOAY0WJI04Cw1C9R309Zc+OqQufSXD707Hz
schvLgaWMDD8RRuVA6NPUG6L/D3FgPLRCdOQSQGeSQvltU4uu9AnpKEAnnNV+iaq
QPDPSrZiSELONTc58a0f/HN++SRWlE8a5p/+w82NjZULR+3NG2+su3omaXyqGUAo
Amh4D1xik8LLzgEHfxS5W6HQ9tMwW9bXyaQFhiZvbuDjonCqyagZpY41F6xkp4n6
/a6bD+NAHBrPBReUHJtHSJ410x4WrMKYAU6Rwm0meeX518UMxbkWSkD25csB+Y3/
`protect END_PROTECTED
