`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7q1/KqBLYkQKZWHWBAFcreWZohXNHH7hvhvfel4/xGHJvyhRdiP2YIg6UIQW9PpU
v6VH+BTbyBaiy0quEM1mq5jX/ZqQy2X9Dt8SVVxeFIbo7kOpSwdMDF/pSF2mOOR4
VD6Ezl1Ml8B6V+DVoN4X6cBzlufRlfqnw6WBNfMVC8XJYk7hOf3nFGAF/+vgBpWt
cQAa6PAVrr7tdfsO2QsBObB/gHOpoKNo2la5NHtMZxiLE9FHCj7SZEMh0ASkaetn
FWZNCuDPAGEohGuoTlV6ZQD9SGu3gqF5Chal+aJZmy7ROhTCmJKmBPvIIwCcClIq
omLBvBMslJ5myBHJEdeQOG4E1nEU4C+rWe38slRf1I+vkhRLPkpmkt7WpUEpXRFH
iDqHDnzVexGjLUn47qq8K9nwMiMomcvbbqCiSsn3ihNk/onSk0brASefqGTa0bwZ
tPcTt7seiYrTOphZJlrnUa9Qo1SDIPlLjunH4VvwcaVqMeCcuMA/9HGhmKQZ/aak
Stw5LHgzXDAdf60QJbQ517CUyqE791sl+lqnJfoWvldNaksYpFzPa8+yOewQtPCt
ylsXg3HNsGwVC5XqM3z2dm3X5fcaf99v+i/P/cPl+Vr9vNDI1F+VagcNEVPKzRPf
pu8ixJEyUomcH86KZ6938w==
`protect END_PROTECTED
