`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWD5cpDUkLv6GUfO7/JLqPK1mbV3785u/+/AhXPt1ANo+MHaNNMQAAcIoSEKfUES
62RCuLFCeon0bSKBa0ssLovDcajPOrcI0OBtlVr1Ut5lsgGfdShO4FGuu/D+uzX1
PzYH7hUurcAxdB9G647Ke1fu4B7aJilC0sdg3YpPkr9fKW6dSz2WsQ83/kwNKZsY
L2QVOEq5ns8ViRvvOGevoAO4/j5N5BndUaac8e441HiJtmVUw/E3JiWig6327tMR
HwvdCV6N8FgFCGo1w2B0SPiOlbZIo6fl37gn2/78HmC8KVap4aMt3QCszhJYk5LV
T7QK3JYyUwLb3PI25IyiIqrtAyAqrOPwsbZqEAGuh77y2jfPXqcV9dYqcuj51u8Q
kNqaD5W0v9O9FB76qMAfOPc+7AfH2EMvDQ3JcxVYmkvZldvcJoaqO5A988vBsxrb
PYUokzEnGpezG1rHkh8afrt+FrL5zs9st70TKytiyxA5vy9520jtWwCtbcyuK1qm
4q47q6SZzMf7j+Hr6c33GagCbmNIXY2cjKyOm58qrxvVe0HpDuSn0s5S7oUi+5mA
A6fsYBUA+ONgvAKkbvnZI6+ASFHnnboSXfrUPlTJwrhx/axrYq9HtRaSyHSZWCHK
M5eYek9c1uZ6Az6rg9RwwBOqxAXnQanusNipFTCH7w3p6WE7L/TNNLHqA6CU0Bje
jB1cjS0Vqflrm9zNgOH+huvd3boMh2OROV/JbqWqfYp4Em8ca5xHe6+rA3k4KW7D
MEfPzQ+nflcFK8/DYl46i8l9nq2A4TTP9RRSINkGdst66PZXwdE/VtlSKTNdls11
Jq84EtcDrzg5UuJjD2voMbWxw0UnYG9xewI0tcXoMQ7yee3zEypG7gqPT3AEBaAo
RIVsRdzdgG5pinWm/BMBBcYVtegszYPpx3Mt+JE7abF0fSTxltT1Fzv/bDpYpmLm
IGEMndJZxxjgjmIaK+5CK0weG+zjZ/SAs4Rts3clEkKwfq6yCSdPNgaYEhS5KFh6
gRTmmkuTWC+op36aqN/kUh/7KHqJ9TzLjik8A2N7zGgIjMioriaq8TSbMor/cz/w
SOMRqTkAoRiRJVXtKVE7Iom8s3mH1H45byw6auldUTU2+Rv6FucN3NJyu3+9plOl
qpl2bHkmWOb+QcHukFvd3n9E++YaZcPfbVYv0YUN31+a5tMOF/r40PyXQjL0K0+M
MDGT8kuMSHqS1KpsTIi03lD/Vz7ENQ2s6ZYd/xLgGpevph84juUP4m21e2HqJ3mz
dpwflbwC6ngPyKxNbSywwfBqeIZsMU17j0LvkmvfXCOI7KdVewi45gg13+q4OJ6p
kflL+zgx3l8y4J5gVuwvU+HWOmuVPfQuuCNJV+HTEZSp28W14P4OCzotPYlEidgY
9xErSqyOgesQNyViyxDJafpP/rA7jLIQ4xXaVaysx+2XMgJfSh24T0J8LT4vds8z
6fO3UcAMdhILH6AJoKUNUUAjfAWJlda10EPnQOKIEyAsOKDnCc791KXucyLiGILA
RL0VOyK9PKP1xXWRRKzXKuF3waTMMF8WMyke6WxLgZGg79MTJHDfj/SsbTcyFqRy
64hUyFyT3iRZ/nBvaSKgg8TykLfPzeb8gAJDC5et6eFobyA+HWwH2UU0WxI7kST/
O1Ur8H8tPcNwohRR+yekl0rSYPsmX+tZFFEyJMfmYqems5//HwhOt0rLSsjKCdcZ
aDBAxiHtpFqIpVCJR9E6TFt1s1Q8qPSzRIjoMxjqgo7Hwtw8mzxgxkM8esbHMu0l
VCA0j1fxwkeCoh2Y60KLFid9w098AJ/Ad1crAn6FGpcsjSe0hYItcOQD2iOQNghD
9s7m/kRJxaG+Z85MJxx7hXjGwdTQcu5/uUqefwu0ingP22uANJStdguhuMqHFBUO
nDTn5K5dh3OwuyIzs3zZkgHDrYkyUNW6MLW4SohKNd99ElBnRr11mgncTt9J/t2W
CiaBqZ9dWUduO3rFdE+25dU3MWRv5aEruE72eSr4SBR1tRtOUYMYbDvNIshqsZYI
5fXzouAUuJ6BGYpzgBx6F4ceJGCh3VVrR+CzQHEgfg2fHOSUswy7UMIWVNqb8ysX
ly8Jg4CTBIXFFJB7tSoemZT0HAzDm3nLJhpwcl+8GoEta8ka3erTM8MFpOcrzuS/
9/b2bCci408vwNiBgNOss8ezPVPSH/hW5AqQxEpG4gMczPmlxnmb09ni+7MfSMQw
VO/Vw3Di/3ygFFUsr6aSoU2OJYXOLIrNPdN88i42Ezmsi/hhaCnLiklhexRHJ5on
VyK2d9Hew/sL9ZyBu2yusTQspDDzqJFhcSvv0pbUj9aPEceIwUD8yXovtaezLOy6
SJhw0QX8MQ8ccLEW3lvslg==
`protect END_PROTECTED
