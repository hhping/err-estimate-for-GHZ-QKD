`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HrpxDKrNViJ4z01CXCqlvOZxBLuYH4hkd6OvdHcxSGACoVXb8+DDBtF9sK7OxVAS
iTiaY38DGSKixFCXibubPMuTL/Hqm3E5/Z9E++FK0StCX0uz04CuUVCcl2MPFmQm
gA/tKM48B+uxuj6AG4U8HqEjgb89xE6fIjDOCzVI0UX89RR2H77x1QbIgVGDYpQA
2YR0y1MkWSg3CNH+yma42w3LKT7X+bcD78bWj+YIbrJ1OpWrondkFSfetLKGMqqr
imsST7Cje1xhSsyWrof+ig6k0nelk9NSAXcnEEvAxvRjZXhcjiOuNmRrIP69XUoC
IQZFthGATvheBRp30DTwfAKC7CXSHgeFm6ytSa3NioJw3kVMLw7vydp26pttBfM5
Xp9lFF6m9Kg6pKbAWcdUm6tWMIyv4cZK4CYuTGUUuijqNgOVfc4mxjNTauoFo6pO
XeEaF52L5YkUi2MJhpxHzsn38Kf6YV9PAAbovTYPvBzqhlv3AcBzLyp05rzmqPIy
s4NZ50P+IimyGLJmhzQLx/UJAtji9TMFoKGq/j/aKVtlutp0Y93w6JMkoljc7bun
f41U/RzknYS97ZO2SQMkrnxO8mPqjSljGNteSnvVly7fl+2PNIp2S1A9+mHxqOvw
eUWTU/1vRxTw3LqgfqsjrVPgAZQdhhuyqN2WTve5C0tUAoHRmCANNGgIvOO0dDS8
uzgeVh2XcU5FDVcKSPXANmIV4/+Fbi6qXO/jqN+n7KumUXRuIwwtkqTyY14Gw6dk
+nhGjbhvq+GmiBY3V7CO/+/BZwZ4duFBWIyF7CHsUOFfkfD/n5wTbzLcyalv07EW
3/dGhzHloS1Dp87gK/IqElOQhjlAA37iku9h7I98rpjGmAEI6xkKawERf4LpFVbw
nxsctnOma6dMzybnlPhELr2X9+edl/zefiQttGFJdBfxyiK8w0RbtxrHn6o432yH
CehnjplGLXOXz9Fe0LwsYpNfbySrB+GH8XGtiRHqcuHmyO7YRXC4q0kBPDqOS9Rz
evM7FiHOx0Jv2oTQ9UY+RD6VI6+pYidTpvjWm7mTW+24WZ5qedL/KpNyn9Wbp34j
KLHRmesxob5/Vx5lwtJ/vodGgHrqwBPEV3Lr4T+AA6WkHNOCrMNEBK+Y5/gATmGz
KAv3wLqgiGO1nWsFd0rO3/MiKlHUqUvjcmHNg2voNHNjoSGPG85OuqqVQP6uEL9f
Oh3JAACtxryJ9/9gbPgILOqpJwUduN87ueayZBfiW+S7cFrsmfNMHHoP/Ue1db1j
WgGgwqwFVycWNAs9C3E0WCOmHcA1p8zzS7zs0FKJIn5nhGsv8lLqOX93aUE1+2rC
vkw2PFiEvWF/HozJQ0phMtUA7Ne1YWkR7daJ9mawT9VarcXU5b99xlYSjqlyZuyn
j+7XEHV9Op73MNzXpzPvawMpo78Iwu84KpUfAYrcbbiE2M4DT21vy07Uqq7fN8ZX
RoFaFyX6a+STAgpeijExHlroyCLu6mVMo5GqFtEBGLhrChrM2LGEcFYStOzQasps
Kn334GTJtU66ewQnXRF+gvNPjwUIMnXaVhcR05BiJc4kfVWnXqxISTUwvEFYpmHh
FpeItGe53aw7dlPIFIojQdABMecZ8RDn2nSqfkbz2YXJiu9LJ12Y4bvp6HqkqpME
UkxWh+rjDELAgtcVZn52SIM9cdbgEI1FtLUkJud3azzY7IV2fRNF1lCDZFYPHwfs
GXr9ZTiYwjUWdm0+LUBH4V62kFMvv0FyOlSP93ZZu+oNm1jvc+r02aA4PjhaDkxE
f2DLMu6DhLvchXhNYhskSknqxDENby4d2GPvvPJGjzAVhc7pNx0TEIapfwQtQXee
rhITYC7yeqBwbEGm0aFAZrEHGvoBDG6omyjuesC5MkrkWWgp4CTCz0vY8VKuDhz8
fYy8aeKMBYabZ7us6O3yXCjJ20QMReoLY61TVQaXZf1PdqyjCcQ7XjbyN83P4Eq5
/wm6jwnqZZ5VLaa6cn87dgsa+K6X68qGPloBfiCVc+oYqR4nKfQqzW0j7fStZLLQ
7OfAWMpnfJNoXUNQHXA6PDnhw3x1wefSrsOevvrr6SPRlKo5GD/uF4AvH5RPcZtz
HFD6g7Vu+NVH0ecGJXR12LeANHNJ0wOos254Sxci0Ix7ShpLmMeh1avKvc1dmBkW
HVsQj+YixE4d7KaTcauVqDcCsXB/cLFD8Vjk9YMBJ5dyijacQf2MyMZxMbqHFCfy
mxk/SbPMqpTFTbqKQnjzHSBINTpCFSx1N8JMiecg+Y8HKa3+iNMPewPNn1/O84KA
FCmGXH+/WXkWBjSHXY4fh6MohhlyB+XP+kXAxtNfIbwphK6bGG9u/ukZ7TW0dDJQ
Rn62HahHlkYg+iJO7QhVgc0xaKL0OZWDsWvM1CasHpnb9OLLqsgo6jlx9Z3q3onq
9QmuKbBPGCF09AcepnT0sdLJCxWDdww/uv+YY6f4pYIaEjAVrD/MHQSmz8DEqN+a
ewZwfixRQp/HyBiEollTLngtuumDBnZVcYUI3cwBiW6CvCbAoeKVN/Pyfamide7z
xe9UsdvpJgdYzDCxZVikyK76cTNoTX1g1KIDXW3NzLyzfCYxILPUY5SH2x9XrAFT
0YFVTkH/OPWtGAD4LdnSF6L5xEqjXnmtfo33rS2ypxevIGZaVxKrq1G3G0caVkm/
731UaxxFM4s5jtX+UJQfarQRYA4S23zhGQt3/emyVOucaJb4HVz+2NFaq5e8fNKQ
6pbHKQaNcWL5N2xcxhiBZ57jLu0gGAbFJEPQHhxleRbeYjjPYMT7shaIKs3OI+t3
HLg1hY7OzYaxyN8/bwdbkNAEGsp3iTtQXHWPQTDZScs11E5UT7oTaVpZTLvd+ThU
y1p1wUeurH5uXFq7Ofm3JhZuM2TQAgzml9W8sJAqMt+SlyOVYOK+t+9ZhYDs7YV5
PcH32P3ofnBzCUorR6DCXmTlRcLd1fTEgron0tRokmaiVvVNf14Kl/UMHrDMto91
0j2ugC0dlMeZkMLLpZ3LKJups5lM5Z/gyYzODmSJpJWlBVGcg1nZYajQIzH9/8rC
78w+lwppR/D4UwdPlkpJM3Y7u5WcPUjaWzdJtyhZGMIucTa4aTKjiqzPLTRzTqGD
6Q6TOK1na9nUMPh8ZFAYHnbuigF8mINYbdreL+/B2Y/Gge4HyxUuyIuM1hM9njP1
7TEG4+EoEI4TlbACObI+98Fe44rP6YRseoypmqFQyghZurpJzsmcL4VIv8Sih7c7
2ooP/KwIzXcTELC9pCqYzjtAIKrzLHc98+QF7nDG06eikz2sC3Fy+8+ch3ajPgz8
8MTG5ltLil91hj1+/wOHzuWEpE8/nm0ZTZseFB5pHIHJqyzmU6MrvG+LwkDKRCCh
VzS0PeJUagX1jhnLejE/a3MGCXFYDAUe/H1O4uRexGqnc6CQogm0TyrJjgtQrx4h
v1ZpGff+8KIogMUSX9W8mC6YwzXw1Lv0e1JtmsuKtkJGQPbOPsZoYdhUv2K3tgVp
MjrPSRWFLSoSbbdEvisjRyekv82olCTYOM98zRYkVyW75gM0KYrSGQSLXndF7IzJ
InXXXs/gfTRS3jwzYxO9buQzChqJZxcfT7fDHs5ky3TkcLMAN0dkNM6qseyAhnnT
TubiXv6Xx7Wi0zLOl3JA0RjY/jBt75EWlFj2nMoUsYSYTJ3e+aA2UMOcEGDR1cJv
CTIiQGt26Jdx9LvJ2IaMUAiRpfv+Hivqkw2pDagziNyqgA8yg2Cjepity10dLhET
o+ovsBDi8QHQrcsRraWUs7ZT/Zobb2QUXkmONjmJ1nM7JaD5vKtx0XPk2oC7fJnd
2wJoK1sUNwCfdzcUjCeaPhlOds2HHxPVOnd/AFfWjTzIP86QzF7qNfld8au53KeS
26bM2/X4YCL3UNqpgsXGnDgp5xP6ig6rAPlaBv4QN+K9unvrNyFLWs7oHzc/phez
xikDlQUc4sd3nxIyVH+VHYD9gYqhLFf2uDchxwQwnAA/udKelB0kxedGZXdalP7g
zmLi66XxIYJj6xI8O9gF3/iZp9z9lP4xOtf8R5oz7w1BfNqvvMNWlDf+Yks+OBbd
lcos4TlOaKdpnMhbstpiZWjMOY5K9GUDEqRwsKKN9BPxZla6uB/IPlOL4bZCFWP7
s6n/kRTOZJmPg+KTCcOzlW6A2bS+4mD6D5ysBJJ1wXd6sbVrwYFw3+5j1RDTEn9K
ui2+9THtVbeQIqkdpQaxPEU6to9BCPXIvW5/bGIcZmOwL7XzRy2PL8Y1kGoHrNAH
GjyTQbXluBVHtiOz9ZqAacn+aNyxNgwNlps+4cl0aUbXAxM4VYc749vnJKwByFD0
Gv1/6J2mi1SGIlUKUSMO8DhhdyWmSS3cVwL4ggzgdvK2pJ8jBh28PFX3YyVvmis9
1ehoz0ya3WDBZpJvged7ZP2fUPPWbrqv2fz3jOX+NQnbgLMo/rL9XPiqFgRV4yn5
X0sXpXUilrX84TWYcveV16YV5gxvD+kKQ8FaxTAuLIWv8xTouKA0v0QEP3vYlPkc
yZfjs5xRM0jBG217qtcBYg2Jr2VtcVeZYM0ihlB1eclk20ozjjyg0/sYHDzKiz97
e9UkjXg1ZP+FFhJtEkqZgnEI84d2TDm3AvUEIZjHe+XsxW5lBwAMkJj9sqa6I+IL
FQ1chPbhitzFlF766tIzYiSeY9D90Cq8Zn3Ul7yWp1aA4dJV9frUUtnxbb0HJBDz
TZTshhb8+EJcCzlSa8ksUDKu0eeKp4fht+hrwjgoi0LU2s+yFeQj1wwqyMsErwdZ
xbqBr5/31Na1v28heTg3vAqTbMUPi861OOE15SVxLQYoCIFqfYvgRuhGLcW3DylG
YmNSOv6AJ5yGlJzhd7+n1dcVuVQtfMcPbVfcra4DZ8mVd6hq5l/CvhFCfxm++MQU
3mJdfD97EILb9zKTiwxTsEoyNEqfhIeKch+CkPe1eOTkkjDpkHFZ3Ie3XhuEBsyp
lYIUr+9Wu2ly+jkUxzw3l1jy8Z8jx0whiXv4zmUdIje3mwz6DbRaaj0mrVBtftYj
4Quahcb41715EY8oFpc9X+McYiIxAemPqFtyuzGWUtgQ9nw0Nlvy45CCEu+aUHZL
oR2IjP19bJeaJhXR63CMlFttGmFnGkyWfaeWVihvA0/Ci8Ab7LLohL6pWGlsZKhw
acPsuS2sFzYMDArp6DasUAaAf24/Bv6M2TFVoI+ojl2KRLQ4BYxbWZAasFJ3V8Fx
eb50RlDQbzHvPTf6lYFBR+6ponAZhPaJ7svXmJGp4qmGeICO4mxFrqHL78UHTT4R
HdLNB+AqZOJAPGEoW6FmiAMT7NswCCVHAw042BXDyruPgWp1xds6SrnXuYxBYmri
Oh/oRIm0zRqVAHR4SdAyLyUh275Dh9flIdqHZqSXOOa2Uni1noq2EAF6IcD4BefP
V9g+ScS5loRxLST1p1vwEscN69tVUfN3sv7xu3B5/qB/JPUA6FAs0h5GOo2M1zzs
HjbCcnZri8mB+1sNqTLBJDrJ94PHQDHw949M0k9nxJRFPWsF1KNUopKdoB4wo5F/
RrP0I6lCaz2MPtZHEBmGiJrPs95X85NYdJFnmn6y96n8i13IQS5zOyyBBVpRxGjY
yIs+QPvIQYgNYT7IDCUfLzJie8PTc1BXrI0CZbVDGtN3rsC9tM54qwU1Kd3emFWI
OeF20TaSCzuB16jBU4TnmTEmVN+cf9/MIeZWhTOunuxmn+oE8vBFst8T0/y6YnSb
Mt9Je9ruYESz8TYDmLbTq9hixNbDVwgzxeBk68O4QsKGc85eybF/WMOufKfG+UNp
j+SVH97ivmzKuNeA+JERLU5jiasAil9S26MI82aFb6nQ4xxb7RPOps/Bp05McpUz
aR3GW50IynYIqHAlxQLQiF6JfWLo5vXwKt7QSQPS4cAKhbIE6WvaDi3h9lof24Mj
G3lWFuZ3iHMxldEmjdGp2kPZj+VQWIeEd7BUVkc6VKtlkF4YrvtgwL0soRoWi2IY
/PD6qOPlGIIc5oqFyscuPevS/wmQkijvPprt/oF6oJ9bSLqmI4zwyFm+dzU+cG6z
BW99QX/JnlmF9I+H2iM0E6IaKZ1aZ23eaLD4/Az/h4C0Vmz8157ognOFR7pwnDHK
pmxrO8TtTjRL3a7Ug58gqbnV8Mj16bRfcNU8f826igvKcPYg7Zrxs18hgyYhlCET
ca0DO0CjM6a/WI9nZ4JTM9UxHiraOvGF71layQHwOcwLn00A/kpcC7km+59AXNFl
NRroUBGEaOVJmLARmAh+PwDOV4d0j9o27YJeF2mKPd0/0tBPs7Gt+0kpil2ToMNr
FSc6N/tv1aq/UKCeLLhcLTTJPwzuh3yIKP2wKAIpv6/R5qLgHfNNYvZ3YNb8QSPd
W3zx0p6FTgoCuHOGxrro8A9u860J85NHdI/XpvuefynLUIqolJZm77+1u/wIisZi
bqfx4pwKmn6oOT6cgP1bFaidNQlC0+grsVvt3WtjwM6+Cqjka43nBYik1flYzuLs
arAFvWc+bLbh/Z/gV2WJEesXQa+UbmrGx1BUzYoMohj7O6c2FsSBdETiVSDj+ZD+
rrSB3ttk8bLvcGxHrTnVGmdvaaWOQuhnxd6qfs9XP5poUcftqz4foLoFxTpSxmyl
67PuiDGMyxBadzYLrAEYlJy2KXVmP9Se3O0QOp4IZ7ETBemmMnscLN0gV21VdOYk
pMKLeq9B0H0VpHUWE8bJkEONB5Lb6egb6yUTe5jDQpQSXSV472OQ1oueIRRrt25H
0iJ2I9Qc6XR1EuSD8KI/bLohVmp/pkJ1HsQVtZEqAkNBzcb9WQgKv75GLesNtkP7
t9SmvyqS7z5ri5a+kuPJBim1VQHCKWZt30WgumHzTKSB4TWU46x0Nq8b8zRxi/ZN
1742ccXiuLbggJlMG8Ia9xPcd9+RBe0ilzxAwnyDPCOH1jJql/cZ4Juol56e2tke
2o21QDXSrkUW3OZ0lNRhF/T83ycqwaCGmK4uHgCK+p/02hnvoGA04cNSj5mK7wXo
+Dw9et9CSRjDxgtIXekXNfUEwJdHRm3RCJapibUE77MYmO7nfK1reS6y0OPYfLBY
Qktx3ibl7n0WQCSqStGvSxUyiRmrpOrPCr8g53fIkZEcA1njBTMDrkYq8e2JFzFB
sUTjG4d+isJVr7x8rSiG++IkvdR9ZA9+Va1yE7jcy0HjJU2MMTxV5qqQlNM2dCbq
cLCCcVVftiRVJf+mW534RIuL04l9FXteKh84C6RGCJRKv1tydPdhE0ImoonxfHbL
ZgG54iUXfi3eJL0Vd6+YSPEMCohoSrsEQMidRMR6u6o7hkXqJIht/QlPv7a9WUtp
Cap58Prefh36vSCTDXfZhLxNlXRKUbjzfZjvcAfrxi8DzSFS/p6BZ4esyegwYS0k
G9JYqpxYEqmFCtVKd9AEwlQlyjopbr52NPEED75OkNjZu3V2p3OBtagCfLPzeUvl
LrdCpMrJZo4J6QWBuWngcLI/jPtCjdEwqZ/UrhlzioKsOaUa/HNFuDJHzg1aWS/X
MpOGvVQ2i2HJzPmk9l3gIpVbcRkY/mfI0KFd3yiZduumufrcmECFuIzHfaTUr1PJ
qCOvZ9/3JDuweEzKhGENsv/ENV8e06daO4i6GC/tYL61/iVjGLNRo1Woo6s4K3mA
NVPWvmogFwUiAo0HMpU2lqoYbns3NVfvUAv6Ah3FR7CKdZMGRVEVZNDyFawusXFp
QpkrFVB3DRkBhrDjwjEcc8UXCzQdVyERFvlYUwuLzWZbjoB4iyE9D/+r2z0fSw4D
QMgbRbzsRDKX9FACnQA8u1/Q/9wu9onzCDP6kyfWWYThkt6R+miglNpwmjQQkVgK
mXMZ26pM7UP9HqOPcrpWMKwQu/LpTCgnbL8ZvD8w3aFynwMqBVmjOSaf7Eso97of
PI08+Cl//Ugi1yhv1mdgqYFXAgDoQDAOTUqowL9p2WqxFhOwfgM+wALx5eyx4dCT
O2Iy1UgdYkeTdnyzQlnI0r/lcmjjSVaxWtt2+FU19PchD6NH74wnMJJicw97+Sk3
tuuBRlazxVGTAV5MNkNz32lTHhQq2oKXqJw5SOFF+iEkMCxLWQF/D5lprxMOQjrd
na+4gDq78P1/E2ce4G3PsmfzJSE0tKTHGFjNcDvX51+3SHcBADSHHSBpmSygiMYI
GZyPSU2gnIDp4KzSvvtToUgwMf2lZFm5bJzBg/cmQzN83PuyBHBKHM9ryg1H2ikF
aTL6ic3Ehj/kJXGyTLn7Qielh/NkCmb/eHZ59B9qZSzVpr7BR4VQnQ/8PtNYero8
GNTI+qPvCXZSgXH/Wz063MRWgh9G0E5e/HbLFdUt3HIFCX9ona1FUKqJzXu3cHUu
0fd+BduAP4g3CgwtT4jLsCyaWCIuAb2yq7I18tiDkuuJ5wcByr641mUHvdESOY8U
IO9OSRatbM6V5ffYDEDQGzrJJ8lnR2h69F+FmBZe1AbnNzpHB+zM8NtY5dF7rRHy
Kq7YuhPjwoU1LTOUGl8N1Ow8VcISNIZhtsniRlLI8M2sjFPIhSoagZ0LQ01ZOfWq
Q/xab/dEbMttjs//T5Ou0D3PcZdHLv0H4YaKSxnZAKyr8mkM7FJELEe+HvhUUI2m
YvzA6Xzj7rhxAu0+C4ikRBwzH86VRQEcqvoDib91yv6evAY2wwUQgnEUJAvPKrEt
6nshZeJAafq11rUecq5+UrtgygMiYDofnF2jCA9TTJqzytK+1xwhfibCdLjvTsWn
sKw9SVXZvpODVwsJzWGDYMhuMFeQiv/jf5Zy4JRLWkBAD08+ACxa30cRKaMZkXJi
BSzyNkShsVgbFiWJLp+HcPykUV58/6npnV3MEqqWUf4sEtqzAWpk0ST2klakdMM+
TExfdcg+ZZm9tnBkxLcTGkkGQp9skxKv2pjgaKmVQntQ0gnQQ6Mq3F0Gmxj5Xy9r
1cxXeD/Lxc/PXpk2JP7dkYSahWmyT7jAzYkpgRDhT3D+6fWIgoE7sD0+JgXRrZcP
QzUfBqGnKVlz+gTNVs389xHUwMFg7k2p08qGdkVZzU5k6z5OBekm7mh0SVS0RA/V
aTS9jHHqj2QAffzBmeJ08t9J7vYZLOXa+iXripchSEAaJK27aw5ym6kXxqWFPMbl
BfwvOB9vkV+C7opEkfPTD8lrncf25RjGJfhPG+oILOeF4DyshfRp39xWtF3jkXnx
7G4t5j3wB4/uoiqjuuj5OZyz6tsKrqgLvDdekilNYpL8rzKzrStZoSJtcA9Kdial
hrYcK7Sddx74gtigDdBj72UCCWjpSKTn6gNSn1OAdhNQ2VgbY0rDiITOZteBeqlR
+ygVIWtpbva4znI3oKTAXI0hHfJd/JHJlWwSVhsbAeXMowy1U/j7WeUgfmDX85I4
tOIZAF0+AeS3+GPsZA/UgFO/eAe6THLn/P+u0g6/zwEQySQ7So+P9/JSDtX3F+UW
JkEeWPC3/nc1MedgOFrUkZK3qcdzOQKOcX8dwJHsmmvs1ghJPoHMLvEk0UMx0J7v
nLPYJ0fnM8pwxNhzdvOv3zPjVc8r3TfGvEvHBfqjtpXPPTGi2TzVKK9W3c1vv+sb
OmMdZDi1d2exWUWYCY+t5i2U+XgNPGLwOzLUeME90W7rgK0ZyjIU8JFAxmCBK5/x
MSRTXo6TsKsroFpxphXIM5/cY73xnlHFE7yDlHrolG2Sjw59+grQ/cCT40A8JFM+
Hfv8c5ChOxAMlsK1oObwW0BsJ4KsG70cWulHduFHSAetOHJI6mx7Re+FEpLS6AXI
0qUuuUOs+R5eFNaUeSs/OfKrhKxMaypgOQyrYw/qZp9hC9HU24Q9cO22usk7bzlK
Bga9fhyFK48Q0N/dCPHbo5i0aOW6GmvvvE+05gxMxM3qAmSkMuwxGtwq+ZQFcV29
0jUMcL/UmoM/0fyuvl87PfhJY+3FFSf/OM4UvSgjLMnLyed9ztMpLnVeRbfN8WPX
01XWWLHarUzHkGULMEy7e8Tsid869nPL5D++A5WHLMwHrTwxi5EOO+ojikkOZjOp
KBXtIMFjcexTz9FNhPALCgGoFjD4tVKctzkT+2UXva0Y2vzdU3myY4bqQ3mGHp8e
TgqB6o7p77Q5Fv4XfWXNLUV4y3IzOmu+/iA0gV8vB0YSH5Rg5u6rEV0UBJKHHe8l
4cuzXAMoEDOr8lOotOmuC0adkCCh8HIfZAxa7Dl+3g59gIokNrMCZL/xX+kHad3n
JP6ynpt+XvUJKTLQ9k+gMs78YeTb6eX1cnz8Sb1RRZ4VaxifBBX1cbBJ9/dTeww5
WEHdNl3NWEUFK9s8CUv6utF679GhpOxLUYENN/afdtgMA8zA9/KVkmpw2sgBpr70
FpI5Ot1loPascTYOCcagTHqi4EYbtL11ochHCMy8JMaq4wGVzxqZeUgVwoey1xK6
gmixS/dHJ5gV6ra0k2EHYYHokbh4IdsC40QkpdtH7QcCwNbkQOX7OCUHBaAaMVc8
wfYkiYLdPFNdvITk3MF+2EEY/qirbT+sCBzc3DIhULts72QtZ3osYPw2jQDvLoja
kd4otwPbXJLm26a9CVQ2u3U0pCOjUw9S0SwZYJ5Ro8zoRUg/8kGuNLZmHx2dpDXd
ilvzg/FRSNwmjZxiuzRrCkNudzClbOILHQziDJRvfyRro2swKgdAECYXozVIg49F
vAseLOvCX3iaQw5/JXN3akh5qxA4ns/+a5RHzmOI1vShFUvYAzjHSztYAt3sgaH2
luOyrIlexOmPraLu2I7dOXVR6blWppOewYr/JxMic2P2t8Aaj3nLzvJKjf/FTq+J
7qTBJHa/nRHFQPc9U8Kz9gaDPpWCytqS2oasroGDPngFxfZPpMSHoASe1Yhu1nG7
IfAzt1HzONti9o4kEvp4kOMV4YjPaSOm7Py46QcZSf/qSi223F2T3fIVJECdDn3b
5+8ZnyKElN3MU83rm6eLdOSuN5SpTtv0VM0e48TdY3YYPG9GquNYlYVoiTGO4DBk
2hEsKbmvaz9nMIEiEyr1vj+W/6xKn/Iz4WYpS9W+3XufF0Qm8ccGRCRAYgEYvrmD
GtAMNWLKV2i/IRwgcgiVA2/v8/tN88teMCoZftfMubDe2kfrs3l1VzUu+lOHOzj3
2FXX6CEpyyU5SlwAwISfAA6lMIqotMANPRCPJfvpFJbg+aRxBlEUtTSgBY5Yz5zA
+1seesuGAKde569uW8FDafpJdmdnOYgAJyQ3Sug5DXMrkxDFj+o1qBTARrJ34aQU
7ZM1KWlP8LD0ToCK9wLDKzWvIsSRucks3rqj8hcaT1+z6z4BMTsW2nO26VbB39Et
2PmCb0hquC80ysasJLtx1kmarDF+DmKbwn2WBH3Jqy4zMzNkHpF3QTs+RNSocytd
TvoY78dIjsZGl2z17OOEAvu0F9kqrWiaAOMEZKSkZ6j7dBBsD6gnDHJs8CER1zpg
PGcq+BG26c0oZUSixdS4TR720LA9BChtVA6W8g06jKQXABUPSz/TLVMG354ml1rq
H+//SQ6uLyB8iSSu9dTk+ikYnFODJctb6EZyA9ZBH1KkzxrQajr/kwzjFVOa7Cnm
H4osxrMWDfEW+5isPi+7T+oeJaDk1GuYm1A4jo604zsQ0/geq0t77eWcQViuWO6q
++hS0KMfoLh7EpSXLJ9sz89dZ38iBVx7TRp9KKqgvb74YP+9NTkUnyRbe0Kw32Tb
TSO9rmNcf07ZpNiL52FVBQMr3ogWeTt3AnwJM1/5GwSzdTO9ZYTdkfBqUP0PmCHu
wXZZ3RwAyCewALr0sJ+lUGDzTPO1klGzV8EoMbRxmN/V/SyAlZoNKPdGkJuO9cQY
LrqXeN+Ihg1kWNk03h6oNt1tcM2ny4dTJ1WUu+5iNdSPtqXGnUQB+UGUAAX18L4G
ae3Dy3Ra+7rk24uzN9WJzETZTDKe42nBOoz5gr82eEjuxuBM3r/k2HZ0pTjwR9Xp
vD89vFn/wyGLyDncfiAdIr+ngno+dHfr4ekWCZBAFT/RFdV+mRQ4Ey2UlU8tsLEz
gcyaS1uSrigT/4WG7ophBi8L0e/MrouyHZIia+oIqUQTq7a6xDESAeputeJh4seO
pEGEaKf/b/TTE2f+NIjgR/BKTpshWcIN2QBOFaXJNRZAzErvsDjPE+MhVeJsf5W+
S6Azuv4ZkII+Jp9TfJyOuDrSTQRfoZaFWneMoSpFZ1iYkfe2nswtkpiFo66DKKK/
KG9KWvEqKSz6rewEdKO1X393xBe8TOsLAxUtjVpijX16IM20Akevnkp5Wsx56nSW
oKgeEjSBQK8HwxoNacveXHZ9Ju9OjZnmU2CH+U+W9MkZmA0umVsuHxBucmYQiP3C
pmEODMa4aQvERjosoWctJR+6TgNhTXuAkHirl8QPj7EURDvANcoNpPSTsDgKL3ON
mXU9mPd+waloq3zMdX3eIUJlQB30WrmzkSNj7opwqmg+gOQ4X8TA9gamibWhor2P
lqPWT8i780+eJMAjRFDL5LHZ5EvGRi7TPmfkjPLY7qqY2HYuo9aBhSgt129dvyKg
+WZ4BxSZ5Vu67u2y4tdHizh3ityOk6dHJgVUlv96SxFLxDr1xr7fOZX46F8dWZ2X
rxjs2tnZMVScFVOSQRFuL4ltu6/xV032iU81ila7C8ObWa/HtAB3i3AD2qreRgVz
rMpNaE6uM76BKSBxAABUh0m9OGQTB42NnlH9sjHsYOrwSSyGfkGvfWla35MABN4R
4xTprxhxRzJ30LM3ySXGR/sVwuq3duRQCMqIBM6OvP9bVzjO49aE622CK1ptEJ4l
3b/0prRhQCXlQ/yXtgxfXbQRyctpN/Cd+AEQ5fEv/GpPjqudj4a2YO1vfcahyy7G
iZ5omgix8WT8jb2+vnrLRp1o7p+UkTPGWy4cDPlWgm9tiulm3p0LUkCEzTaHAtE8
Mv7nz6EBrN4RCUDOXbLb+jM13AhuWqdfhbzo3En+9Nk1G8XBbYKIclxWu6vKYQCX
82lSt+bcANunW8ajW63XF11B4lUQmHcA+BdVilCvlNytpmeHf72kTOXt3+GZ3FFL
ODRzCtq/ac1TbTd/jMZIiQSP0/sjJzNxd80BaIaMN62B2X+ECXVE2LpQhdRYiVoK
CbX/sF8S1Mr+YJzEE32NFyEuNgpU8HbLSOwpJ+XbqVPbDxyxO3T3ac074QqBUXtE
rd5BTrEs6gY2eR0vkapI2wVWf390QxSYBDqaBbmPNhgcLkT0UepiA6N+bz6dMSXE
INu+WUlicMehfobRDmJT7uszE+C/g9JbE6cYNDG/jDJRS8oVQsA2ute2X0gwuTOw
fPw0tfzrBO9b339nkqXFtg4+CqrE36Bmas2l9PakTJeesS2gHZWy+Fm7Q2R1T6lk
CKV3D7ODuAggtiNmK5Mw4AaS7YoUOwptlucybitbE93Vx25ZDi7bDonFGb32MjGK
qnq+w7FLb8aKPRhrwvGqHmyK51bdJS8WLuMfu36QxoCw8Q3P5dnwvNWatPg9euLU
cJTLzZx6nIz6DJkIc3cN9sm1ffCZ55f8kCTk0UAUnL7SL9uWH6MJjaa7bAFLujHg
1btBSo1anb4PYKxBZBmtYgg3AfJSdRHbRp4QVoPs2jDjSW4HnGb48gDIySyOkMDO
w63zooJcFcqYY9211vQxV6WMjbamcPMybW1DF1DRe2RA/fh/Z5kH4BydGNSbYyEj
j5juDVn25PuJeHyGG89Mb5NheS+yJOle7ZKQccXQVSYaTZKtrvbkb5ZSQToTwRW+
uylmrowIt8YwBLkDS3uAph+tAvrh/7MmNhzTgpkjpnXcM3EaBU90tlGErZlFzt9b
RN01SN4dS57OnPBizT6VsJ5G3/CocGtw4u7gA0SbGazaHgygvWE5dRlXnhdi0iqW
96pGPBed2jJiSydArD626kuVDufSCsmBmFjUFQpPuCAwqquPEylFoD+Y9dCQPEXY
iO7Otaolj6zHLK53u6vDrDr/hTp8EsxFOc4U+nHrUZo2WEFdLb6l+ysuxO7bsMMU
BdLTzpuxnOchEnLAcEdx8vU5lFTW8PATUEaccXGpRhqMEOvQjwJs3sab5k3jFiGY
ceJCL+hG60563hbCNB4089uwCdWDTBtT+dXwrwSzKOG+tix/GcFXg+o4ig7I88fx
SBZD3j0E3StZj88Sz7vEa6ipL96cBcDiGAQgl1TNs5hG+RWZBoe+nVC4l0rnYWLW
CyvtH1DaEl80a7At567szKhd3/Er7Pyl9uCOea41+vS2FfQ2ME/SyEM5mivddi7t
ks3mk7fXzSt7lkx8DcDBVOhMCehthA4CJnZmfjPE97YJH7rKumLL7y1RQ2u3c+Zn
4j3j6Mr7SDx/s2BXjHJFqDFbLy5WeJlUIY8SSAv9Xr0+HM5Ws183XxRSVC1gUQYC
uitbId2ShjOjJbRAJKEZ03Ny/UfNn3o2wdyS0H3gZavZQLGwhNLKj0bpZmKWmx+v
98cVpkAY+/4aFnh0O68M6UGs+dU3MNU9MA/MWtvPZAu6bI+0AMee5qkI7wNapIWI
BqmS+h9jmp7eQPohj903CuFPVaQrwR+LAnlRZT4kjLcTcFmRqQAfzQpNHXP3KptF
HBqN2P0h/0SrxqQH5PxW3u2B8cj1NgbPGpZBNH7h1cc/y0suf4Bv1qiezUSpUcNf
ZbBqBSR+VRcJGPjnd8emN9IQTym1GN+m5CA/nuGS+p0rQK6ekS9bS1ltRyKrrmtC
oMvWY4RWlKlhBS3NQpcHslbFMKCV8yapsH5rY2rPx5J38oFiRZAHVAptbaWdvalX
AITSbGcf1z+lRHIxjfYq1c/J2HW3JEvE/x3jMJo8X7kflvAdcYbOZA+6srKpJJNn
hHR59ydYTA10skl55TMAjVaz1r6RG8oTXvk+h0PPMPVbAIeq3Ldh1etldvA6Qh1h
0lbl3D0DPCjn5NC65w9i9FvgSQ1l7ylTxnsJSZI6qLmXLRS3LQpq7pj8SVBSaALQ
sM5nygCr7zM4V/agT5edU4Ga1xYHYe5CovU9GMjW8kGBA3cHxBnWh+giztWG/EzN
t5qjTYLE0o1H9/WgBDgJPTpZ4n2P1nMuZr42LNGKG5Zmq5kJxqnRwF+kd6wTP5ik
wxbYtHuVrzrEBrHIYT76mEpcTWb5UNRZc4RfaqhF506YjCX6jpiTNFw/GwH7pAR3
lJWk0sgW8ePiTtyYMPYYNAbWcMQ90ugK6chKO6cijwynqigXSCQZaB8FUZqV2UsR
b8x8TIqOmugb/Ka3x63whqUg1VIgLa1y1dpft5tQQE46nvsMXxvRpVg2zDeD8dvl
CWhbQCfhoPeJWITpVonSjC8YHT+PRMpTRceJ0NQN/2kkrnh0dPjHNJCky2sYJ5tz
oHZqPCbgl+SXuECCfzEJ/Bgt9i7Fcg8IqXAW30iIfPni0uH7YhHWHJHH9tLhMmCz
HXx+5z4oxPD+sBGJN6Uf4qyS9JSFwPRu+H3sNNAgRQBKpClYK4Zzv9tFcOeD3dEq
mo92NBjUHg67i46marVOAPW6cKs6Ild52DUejHDKXSdwjQ92HA6RW0BI2UITlAYR
UFFSKwGPjo3QN+5CJ8WStO2qhuNojLk1sEBjz4uHVGYppb6cgrTqzc/nSdP0RVlE
pl2ik1Tmxgu7GLu1BJ2ZjA2GTh30LLDL7Vy+VqcY+MNqa4Omxuaq7QMeC8DfEiyE
lCWhsw7t1/OsM7moA7dYUfBvyQrDUhxmpMovrMDZ8C/oWLYYPneMvB5NX9WFZSt7
Bc0JO80B2V4S+dmT0a0a36F5UpB8bAW2CXr/bwRJhyhIPn1Ej3LvIwNrKxIyKmUf
r/wV5lLgOUyhiYknYeVQuhc75Fhsgazi0YnJkud/YAPtI1wCNDbtXkMkth1sCy9E
6suglQUWuDaOi7c4Tt110wyCnIZsCYzimBUtOB0LDjwn7dUiEFLioOPyaLWfjRyV
ucWXfJNn/rOTkozJdKVRjVk6laTScicwYA3QIdAvfgTcbr7EQ0RV1uGG0YDWvcCi
Rrck58hCrTh3Bjk6LE9jmx8LkfGc30uo4i2eoEKbyMJIxT1i1cgV1bFdGNbyPvwf
HOFwrHHV2ggMs4/qeh4CevSy6bb1UiuTaZXticwktkd+1a/qE+oc0w00MlvZ2rvK
zsPVNi+9CeLwfmjPyF3GExJIqTxFRlyF3k6b2AYt2sd1p7a+3CzAEQmWW8KRNf4G
6NFu0jpczxdue277jbdRfCmLXt4Ydbc5yn1E69dOm5O6iIsz4oNirqZfNPG0WKkA
LrhfBIRN5pJ5YO+viM+pkQkjPSV7D6qw1/6RdmITYSdd9nzl7VZEer0giHLXwGe/
wgCt0nbJdRTDS8RiOo7rtd7SkRNIieQbFWA9tXUKCfOtYiFezyXiHtCIzmJM9R/D
Sjhywd351GLak9C0DBxvHGWFR0WcC0IJSp1TdS9J6MQ9AtPNbXSlrSSeOo6EDi1N
fQEXXIppIBpgo6MsokDo32v+i9Oa4tMP5tp6dVjk+ifbQ75SV69Btj2Nen+cpdZj
MLWD8dT7V1SNwtjkvkjiNcjMo+CWfgydC1tEnaGFovpngjJtZyNZb3UrQdgi7O6K
mLt8E3YLIZqfHhLga+7D1dKr3mwIDuoafADQHfutkMY8z9LEPNwqjSbFEuSLwGnt
ZB3AHUrir2d/H/qPlls87tXn06wI0IfppnyFGv6X+b0QUkhqSTgdHaqI1rjzi8ML
z+887R8zxlldiprN4w0hS2/04yOOS/6FqWduyrlnibuTaLLO9cQz5noBDNE8NXzL
tJEKHTRhGGZCOcOBUXvoyhwnihdDdeE5TDDDTHwacZytIMfdMZ+BhoPiB/vkNeHS
4ZGG8YA918DFgts26Gnm4TrncjvJu9TahAWuJfAIPivEy3n9C3KCft8vWId8xM1c
3DugYdu3SUoX/6cEEOzCvjgd2s+jD3HRYCW3Nm0AP0Oc7YVQziuu2+GixY7oiBf/
ty/zQO5yAxxh7KByXc9uZS4zTj1t8zkJU/ScKxCPwhC7Q/d2AEzz3GagNXLVWRcs
j6bZJd/mnGRZ807iNw8MRG/PkdDEnqMaFzo737L/8hCgCsXLdApuTS0XwwWizOWR
2AL1UsKdMRcqe1PkFUcHAO49b3lkYbwbgg0ySyVlXAggPzJZL84+oyulF/fC/BMZ
5lyhxfJbCSQWsMSAbiDJUuxabvZQyDJIQGOaASE0ZxxkSI4snC9E15bUK+98ovnG
u/88f0mC4clEMKbYM83LDezvl5KNOvPFMLxmsAHmHu91lt5npZx7uCw/vp94c/h6
Qc10d+FbVx5lpy3ezGRlkYgbVFxvOs/CF8linLwN2wgroFiTmHf9DT4Alqre8/xU
Hvrr9HdEIEpJTti2tOKPYoz8EqJ+j+jBIJZ/e/n+ZBl+M4GIZOIvI5lWKUnoUqZu
5u7nRpzUDpoRrQDwDQbIEElY7cawDih7HdA2dt8IkmoCrIVjwiz3JPCYIGTMd7sL
+pMwsCEeX3auTZPQndVDf5Z1mFfBqQtiN+cg6mgDoQHn2O05zIC8o/CDkSrOTBMq
E27X8YHj6DxsRCgUkkNi/cPHEXnJ2MGjv/Vu9qiXIW/tqr1NKuJ20FBzY0QrlGpp
5kc6qeIF8PIhdW9p8QLbbz1Ljn0eLZAV0G39c9Cp5KPzKcLOcvPhP+ju6jMx0vyZ
BW4v0ZBz2RTZAlqb0xhSTMgSZsMDkGeqsq2v/aWCwSx16Zvg6CQKgqV1FqTeR1vM
/iNv1jbs+5z24qzfdRGem1bvYsB1CX5zgs93LFqxJf3T2l/QqHFa/+dd1R/2Lf0I
Vo+GgWRKIDoQahm9bxSs9n4Y4x3iVOVGd4PW88ch0uw76uOxoaGHDvXHiITJ4E53
GaYDHjFA6TzFUukhfY9B7cDFXWAuhyqJLrB7nIOitb5C/4uBPOMEB8tljHGch+DX
b7BSVxqeh+Ukq68JF/bnwJij6dUbRhR1PXKXt/LJgQzIvjdXsJdYSNSp0qtaXrij
lsqvfsllnziP54K3teuEBC6cjclvnDNiauwmk9zqVcdAXXfpvwMq7OMhksVzTpDo
3m8RorcX0t9QLGZli7FLHEHMT6Ne+enS/MbtB5zQqVw8KufTR95Yuig9ctl7yMOt
5f8slinfUX2cT9wBq9S9ACTb44ESpfjZhwuO5JfY6grrRLNFzMkDMlKYdEYVkIFC
CdY0X/uwFpyTkYaO6z4UOdoDDOYRpktcTp/pStCdlw1z+X3cgddnpnEPhzVg+Rps
AUOzcHYWZHQ9VVjhC6nCaAaB3H9GlYGFtxr5sSygXPZsXjNZZCbqJLWa/ZrSqu2T
xCTFtewgNnSxjf1CdloCzkLlJDcVa0gFTdNan3CbDPs79pfRmqev3mVB/dm6j3A6
sG1yBN7zh+Lzz2tLC8uG3pL++1LGosHtSWKVYYCl23FKwqZygGzzMFQ54Al64hnC
BA14z2GlKJGBPmUZTHgWdh7lYJVKtrThwm4lNbX22IY8xrtMgdI+0lDHGGDaIa57
czW2fVyTuqJdmw37IAt962Mjwl2qMUxQs8UCp5R6Qtu2WuArgdZl0a18DW28A5hv
dPzfrW4MQlLiIwW/baUDb3Kh77LOvsOIet1oXGpHmaO24bIYu+0vIJck1aokSj3p
lkhsxYC4ioIBVkAWbxV3hbhXY4gIiOHjTXQHENccTaozXsw/5FaW0jJTCgAvg+lh
OQlTsygNimUcidrinEz64qPCQN+EjofgFGYLfN6ZuL6N2AYE3vMBBNQtPBhZx1Ub
Bd1nWUeD3j+3oD3TgY9/yoNXfKCCTpCcxi+O79PgUwd3u2Bx14hMBI/Cwx4pBF3s
J7vXtbB1dwQgmiV3sBpBsvENYCZlCtRgOFXcSyxuhopstI8EkLj1mAvB8iwOiWpQ
91z0SK7UUMhR3lydAJzp4G0dkB1g757gHnD3+zbKH0eBJ0ubujasnK77HFSHfTZE
H1mazVxq38zO7nl7Gk1fXk38l/ZgJHGKXuMkkwXKfNSfjGguGNSuQLLJ8iRjYHp9
M/9hEFddcYz9aLk3MZiPKf7oF17oO30XURdkTQhPqIVctzKoQkgISNOgvusCagzG
QxJu+NYZ4ckUXYXwHxykD7/lNdzq5M9E2S14YQgjwdfDiPLvGgFeI44OZBBYuMLI
4ddP65VNGl1fOJ94+DiaGlnqKCM0KilgZ55uuph17cBoSMuNKvrGHWT220+j1+3v
YS448LVBDEq4xxlP8Fl+7Hyq3mGYsJGQco8TPvEBetvMfJuhogId+z398l+CzNsS
nAErPP1D3u6e0J+uvpsM4HhwFI3B1sawgafQwYaFt3W23Khodpsv/8AFONI/fYo+
qbZ7zOZk6enjLBGlz7NoNA0xBxtKotknPLVN0iblvcuEQX0m5M1UzY2zgMrTTbQV
lUwZaYcDrXEQzatM7oUnCVa3OWAijhw5QESoTW5PRI3znMK5tp/kguoJeJc2QmRU
7IgEHPHj3z6vPtytzdv8BhgBjO3Pe/8AFm/64uwm2+eNvUoP2iRzd0Wf2IpEsf10
9bw306nhyGBC8Wx5YhOrRsN3p1PQ20m7QxCxxTBUB3aagT7YoskadJLZk1KuJwBd
MrLGwJVd+QfPInIUnQ3fQ6Zn6MozHb1DmTkFezV3r4uMNzKv+YrNqh1r2OjnnEHJ
IxoHlomGR25znLqpMkjFKJwJ6H2JwWSu/8gMjsjnDGRsJF4VkGnojckSxDpHu9ss
7jy+S0gP6EV6kfudpNnLagp7xHZgFs45FKPe/miAbCV41sl1zJvY12SQrKc8KHyO
I8KE1kVPYtyWWvRyxbeQ41NRRFzCQJXBDr88U1XR16BMy5Vqmpge6yM7Zm5FyyPb
Hvml5HN8czLItUpZCJ3IdMEyCKKDBBiQ4bUc+Qjnykl+jzUOpgMrHgar4phVRVgQ
4wKYU8C9xcaMotGI0nh9+7n4+MzH0VlDF3OyzwnDOIp3RUx1/0WqUHcUkg5EF6SO
t9snsmYOiwTiQZnlhUHtqb/00Leb5xae+Y9pYdzpIWYG7M4Sk+8ZMU2F9VsO0BEL
b6WCPyfndsMWCQdOxoJkDlvg3uhL35l6NjMXb4spwC9zsh4K1NjKkkZn9gAomSrr
cVUrZ7TLehLdBNkQC3G+G7xo2fqispiTWe6s9jAmo5lcMlA1eevZf7FAYckpfU95
lmeaIsfZ/2BVqzlxcVqabJD1VyhigRmD7hoGojebshnwbpaFPMFD7jkJePFNegpI
07acEys0SVXYZAHoAgdcFdWauEvY04392lSW5DsXqsLneY3qLV8pZEEsGTAoiTMK
2ktbc4j4CJCXSgmu8TCQFen68Hd9AW+bGRWqRvhu8CbdR0g9Fx2oK4mx4kh1SIhX
8MvMPq+0mA6robI/F+FiEE6Zx7Ph1S3N/ZqWjZyjahANUDmH1vWBCL5WpcaciNc1
cfUPgiCNwn7g8jqUs9NFJ/3YpxErZAZggXCeNdupfsA5z5FMOGsKM98+qeFpXEpr
aPXrUE86ZMk1UA2NpmN1mRj6T75LXqXqO0zkwR8et8RcUKBi7TBapFkotREKBxMD
pVttfbGSrIRouys4vm74/faQYgFu1dAZQs+kt/4mcxOjb1DzrBXhVoBkrwNg9uwP
KK3mPO38tO7Bzkrr9s2Poul16WDH/NxXOh+ov7WN3r30+hUPDj46TD05VGjjShqH
rjw94fc8816F6r+1E42PTnI0dBVVlD0Q78e15/+KlipR1l4jd6/hHSm2BhPR1QKy
LSxGiHnuaqdVDvtdRRUEsA6+qpEWYWhGjlB6cPsF9EbhUwHvlAKj3tA6jIcxBsoY
Kqg76fkuzhqAJPMTSvt7VQle7PTOXaExl2HBBJ/6pP281iRmXgLQBZhEH9+mbjz0
8koBCuHhs9KYgSF1cAHxcrtUKFK6zRDBnj5BWSp8lSaK7v107pCDwKKTvncYnEgO
a/Uj2Ixc1Z3h5EFUf+dnIj6Q9+dG3hjjZ7uSd2bqvHiSGsL9ngvrook69AwgwxuO
gpsjoRfDswLtbuzFD+ap6rHyS6PRsdPztx808s4yeCtY5Eg2yGvKk+mz4ixlppDN
rszaBNhQRutzt8iQUsp3MVqNSL+iXPR60/w4BkG3SA7hXht897RutAVWjn3j7wtM
fFQvwy+3ZQs8Ct0O6WaQ3PGF5yEi6l9d46OkAhpsFeTxD/bVRXDaynDYj5c5k2G3
fgYty0NQahrZGR3IC4vRuj55BnLa4ZOpmoXkxHBtny1pmJ8JBT9uHaf2DvWzQMS7
GsZq8zbhSuTK5ypjG9e9l0ia1Y7VmJtjvnQXUTMaeIiby/OL1veQFpRtqHramdVX
eBEJQHqriyJ5tsCMNlSDGNlS42NoizHsoswWj3nzJ5McKrz0hP+tGFXKoyler8wV
T7FCB5hKvSUUa3m/BaZ21ajKGF/ZMvG8ZDK8V8z7b7LqNsl5e5BNuvNDsZq52cVo
mt+R26J1pQHu8Z5o6D6aHjUFueY+KFRIpImSf7MHw8X81StkwprSXazDdYuqOEMk
g+CIsSImcA+y2R1qEuYrXLcoMyg35igFq1uOp5ahVL9GKaGOeU2RPdrCPwj3Gojv
SBBtzRka3L8YO1TjAusPqfq0lzqTM9Bn6dqMFWDhaSDtalFDdq3yhDiDY9AUeHmP
8mfKxGOFYTI0mLCAelwyenRQDltATbXdsLUcbUnpyBuIy6DKqj/FhnPA+v3+ftfx
mFfLA0tqN/gSOZM05ynFbg6in1CtNORNkfgMdijd8omym+hGsCP2AfulKj7Q1aXN
EXJTgnciePaEEV6lLORDeA0ZDF3k24w6l/kbWDON9YidJno8oG/89q7+qvV4wqBm
e6w/lXxMmleO/51LCMQqFHgT28oKMHEvIzqBffTbYRZUritkJYS8f5+I4Rhe8k/M
hmEg4y5MQodoFxT32XY9nnaaW4dBaKLYFWEx7v78GnPQDOeKd+AnjYBoQyl0u961
nZ0+gGZLM99fq82ENwIMQZiNe98T2iIqeqSKyTI4xdBH+YPpioZtT3kPflCtkp2j
P3WZtHEOJ0HhHAuvOE8bjvXKCLW3fZSKNO8lyP4AMj5yDPHi3vJg8z7c3eb0MPMs
nZNWNUkHZ7VO23VY5oQ0gmEM57r53q/85qIc8t3K7W7pnRoSY6Dz0rHLCjjw84C0
rwpURm4U2SPWSWz2gkypCYQQ4W0VNv60WFMXF3ZV1amZv/AWMDUfTeb8gItmYOby
5cfZ2ZiQ5/E5eOHHT4LPhvwhvqJiQHD/DzNXtqaycuoQ2YofW+cM75o6e6ZnsoYZ
AGIAE1Heze9nEFl080bExRd2MQkOMJ+oLmu6MGihHO1ID0nRnxjbCdu0PgX+LZht
JOeW9MiihSynspvx3C/r+XbquOSs2Y7EAaAM0PrpzYZHR0/idBJoFbzg6BFnvIXP
req2c5ofcx+oA9dig4fjVTLOcip/CWgYteXaHCjcuRbXfiqqe6eL/sLih/3hnh6l
vWgTtdho/OaLkFoYI4EyAyLqz4FpJvlVEtATM1FZwJLFzbMhg8E+boUwCnQ/Wz86
Kj/XuPuFBjOILCjB1JQ2RoeD7X0fZlRhyIbr8Ve97PG+4dl60dGZ/q45hOBmWvgv
yvKtT/wqqt4AJlO1xClzQXs2v5TlpPUtqeprD5G4AdCEjKoH6DiR3tZ5D59npcGJ
BTZWdg/G1wEIjqmAvF/ADB9zFOecW6kGp4YFTxldvmKvnbezGOasMM/4FEl0E+er
T/zXk0kMm0CLYmLE2NLWPYTvC0S9h4PSw2aCN+QXh40TNwGVCB1qAMxVsPcD6nPd
kXpD4yL9OWiWjCEfc4Y0ULrpFR1HM9esABNvt6jrM8MCF4WPEwy5k9S6r1oZAGKN
2GsrYWdD99yoBjGL7i0fgqUMz11lyghT8U/l+RljMtS8gfiCG/UmiVj72LqN6vmt
5JhSiDPKHOpzRqHWZKrY329PzP48VSkQnjGXTAUh4Q4z3vM4/3nmAs/eXGStPu/+
cLJqYsFRl2b0EgXbKnXohwTKLCRFIEkJBSOvvHjVkW+5Z06FTcRfw2NncGnytKeU
f/jPi7S4+reDQBor3ci1fXRwUTFNvp7W14rlh6FDIf70yrIfD41Ml3CV4TIN/ZlL
3/jZdU6s6E9Xe79CxFDwtWm6LR+q3ZgTTPItthJGSL+6a6lAcTcGMoYnKaUdiqnN
7qc8ZfTootWMwYNb9vWxPYzTzPJ1v1kOkdbS1s3ijyQpNjEeDKV1fA26LTdVeIjP
QLO1OWfK3X29s99HyHGtIWMfwQzLW5WGj5pcd3kroKunrol1gh27ksGWl1E9Q9S7
ixZ89oziRh1PQGB4jKyCizNzEN0DcNE5jCzH9ocbJ992u2cwT1HABJu/8ykSOogY
X34c/zuIhm8Z08pSTIRtj4137+BaDQEGGxsyQ55B3SDIQIyjPXCy28AbmWN1YyEi
1+jO/Iqzi5NrcBnCM/KsPkxd6RsWNJr/mT/FLLd6JG80ez3vbTFOThnZPLiqjGLb
jDsvTAytALZGjt+rCCUZiAV9QzwPpLOyDgvvcT0WA0MOgrm33QBiCqOQIYBYoWGt
f31I/n5Lj/LDkBu4T5eTXKZK43mK7bZMiL4SKcxnnDBv21rLWgK0lRX8YulOCokY
HNZYdb8ZdwQTJm6ipfGbuNg4M5jp6efDs/RXTircGJjuH4ai9y9Ptw2SiGRLzQBV
Vn48DXpS54j7TywKkDwpGlqmLkDL9byJmcbZVGcz39c2aoEnh9y/4b6tYVh5ZuSg
x6JreKLruWX7Ecvra/4lCPMPTdbpYPlMNYrqr7sOZNfZsrq+gRXrkDLbaqiyHu21
RZyB6pniD871ELoSkMjCWzlGAHHhLeosPr2VjA5PR7Z8YpFFAhZ1WTOjgr+C9AdP
myYQD0IvoAGmp3j9G1tE13JSD84MZA7pMvFaAp1WykAa3CEKNI5wHCM+77VRyMsN
Z0TQ1g5AI5XzrcUojSw6/R9k0h3IYLJPwBftA6oA7/JXG+wx9lsH8q6plB6lZEvB
j/9K2HgubptAz/Wz2k0UyhFllJb/NxuZ96koEKFrOGurLF05DnpEvd/+nlSh7TrL
uhTkD1aprmVuI6ybjZBnuJjAEMl9YGY6xHHDtn078FGhichtpR+RT2k2rPVRoaBD
wVs6ZmB5Gz35s05Yt3VDGFFX7TzebBtfLCDLjNEM+vouzcyhccEpp2w1af/VCMlg
kUu/0iZrgLglj+pQ68Fl4F42uc4K6cYInz20S7YbeSqeYStbddquyGqvvVu5+d48
STz6v4yn7NaQDUDvfdUaBYwxZj0JqOV4EATlO2joEyS9cQ4VY+oUoHXOA28yqwV+
8RRuyRcoSDoPt389XA3t1mHghKw4mKS5CSyyOFtxKVv5xZxqztOEsiVum5TU6/jQ
fjEtZdLEF0l5csrTiEQiPDYZMICMIncLz+qWmxET7S5lmSwRpTpoNuKzZccepags
x1cBNH+hJGdr2W5/tyMNsK2wiuyG3iUeXudgO1jsy69uLlHQv77PURBR5vOyde/w
WiXZzA9iNmwu1a3GzkSMmCxLJz5njLWmW143Hk07y9uJanaZYXwylICn8bsL2lay
kDg68RNEgfLrqXYDfCij3IYRmiQDfl5OWp3Zsrqiqd3uDaXcIBBCUvz7APCz9olq
NKW/Y36eJlUhRflWhNOt83bukDEMO6i/lb0k0RbyQb0rVBkU9ViQJux/dR5AtdpE
5hS4hMYTUnyrEvCIfu08pGZlUqw1TFNAP4Yjm3BIHrv5N+oUcG9rmToy6/MgNHB3
iZZoeOXbyfC6LS1paT3ok/gUWos5+mIkWlcteOpCY9yYRy+/c6gkzQ/l5QRNFuf9
mHqxbqfItaojx2l6tdL9/6khk35V0bYU5DKKkEmWojhKQ2C+72UblnG8kT6FvVM4
Uk4334BArR3ERIg3Crgi83pFLY4hV8oj7DOqark28ENU3RJ9Ph1USbYNa4VtwkLx
QyQGdZ4wUhLkSt6PLM3UPnBdOngz+ZY0j0ub2yneSO1wrMx63lg66Tz66TkfkvAR
Hh+ZVJpXhuM4BFkJ6hlalGMGsrtBs676rah5mFAzYN9NxmNXyBYl5V+8++7WMGif
yFchaoOeGCgi5gefTuPb7RpjVaPxNnKMwAVlVHtIC0fI9IKW6ilQy+5KVagYyHw8
1C0J2Q/BnicsbhB1gINjAcUpvKaovOSm7NJrUQO95asOj3ASkqclhcmql+TEu4FA
7n8FZbUOz49u7IhTOJwgjAQCvUFk/uJWbeWno171uhLbnN7ntHjVXwmoc+Y98i9N
aQXUIJIoYtiHLFneWb5sjkXCF6atYJjDIDmYmVrWhKzoZV1bwG4N9IynwUrn67eu
C4uIiyKiCNjeYWFIpszWz/dTLShFcrc7c/dlNHHNFEa8QuBTtjD5Mh2p5H3LbClW
HiYVPjuOhbEheKhvrwOxFnwDRFzWvLgVUvaze/O+7cj1huKJzKrXgvdfio3eoIcr
1dpLr4BuYaHZqJvaFAQqJNTLtHHHCtsPaqRA5Oi2v6K5mAsiAc95CKdgw4Ks+tCb
SvyoiHKbY2aTBgVdKLp/zEytHDFcyEqzCa14cwfcg3bscy9S56SNLhgMWzldoEVD
3fX8ds4ok2VoXDO3cio+MCZ69J+5O8aR6ESPqdT4ijsd4a/OV4n3ONa9rz6rH86U
AtL4H1iot08Wqnko0uqphmS9pe7Vwz4uDmzHc2rMqdP/33jGwnKAhu3Xqu7zKF93
ARIw+boFjKNcBTpMQ6R2SgJk8raRGEtr1MS/5bDpTn9cLWVw665OeiBgtQgqmq7u
bFau+MSSTWAbebfoAOEOpOpcLM2FQtb2lXvTmGOZgllHZIAGmjE5mLypfzCTeDww
QwzH5z+J84fZSix+wBqZ5TSQNSmyhkVOy585adjIcTkSemF16YrYe350WO8EGBYp
7icZB+EjSbm7ga6vDtreGlcbb8P+xjBYxUVRQb9nOgxbrxnrPZoD8U+SrLsg5IZ7
kd/kNQKIDD+E2b8xu4vT+Yy3XDN/nPXkeWXjC5Ibj9kRzdL8nM+H1h2Q3CXhokIW
puhrnhTXFthR81mmgqQnV4srKlI3x0q+8xAALgjUtnZlqNdBrCPi7+S32yNh8Cfa
z+x4syxd/G/4FGeoMMCXe0AiZOGVWwvcjNfROkZ2KqtYVPJdkZH24qDMU1dOKRx1
65bNajRxNoQWyib8NRp82OgaV8Mdnbu3/uF0op3KQVdKL/X8tH0xrYgBOoULivVP
fb/XJaRGhqMkjGVfp96lFGPJn1BsxgloVweis7v/VgWObn8j85dzpJmMjgVN+cWs
e0xvKculxvTOtgx9E0un29AMCT+Zt/xdt7oJ+Nz1taEJomYqtkxOsne31fCzQNIR
fJFW9kwt1oRYOCpmD7UacwzOW/v1cMasfTvGqPdX9X4CQSnX68MlT0og/ATdctWQ
khpqbSz/e8Y7jKKHT3gYBK62oxKvOP+AKMYpfvZQleaWoX/93MOJ/DF2DkHggC4g
Bzyf4DeIN3ck+WtTwnMjPbslnSbjwgSpqH81+M03EF3M/BJxIvcjkVmtdy6fV3f9
y2lLO7Uz5dblhWTUn4Qweylm2BFm0Rprypn96LPGNJC0DwYCa/G0MQMpSZfV1xRc
Bysw0Uv9lIaPtxDQyC1n8zx6ERc9FjJlUMH+72wIGf2q2wAY760Ja6/IbgP3K5Nj
1HrA5Ij4m4EeRoJl77dZ2UJSbYj96QFRZcVd5F9ZF5LAibZhdfvXqDWbg8AILWqz
I4mG6A/YAwvOOG+ObqUHh5PtzwUCh2/Se3Fn65ENgLqtWNnh9+o6x5iFgojRPnUy
IYWrKLItHgxX6SxUQQ02uMEY/SvK3Xu+Tci33wjt/RncPecFRMc6KAcl5rI9FCC8
PdKKu8jdwmNRpiaDqnkvd1LAMLDf2DTSCwOjIupNIIUmyG7DEkhjzhny88PjvkXj
/ADp/b2cJ3eqHpmk2UXg67LrOtyXx4v8IuHM53JHBrf3xHDlPfqYgKK9eelUDUVQ
zoYfV3KBhF4h4udQi+PfAOT2MvXzLUo8kXX4cTnI8a5xiss8TZ6ck2n9VbtjbKbK
Xouu5+0sTo6zMZe2JBLXqbo/csQKrMyxGfG1P2VbUeiHNopk2TSR5cYkJ0GaQoep
JhKNjFIRqFC7nTd6GlByJ0+e3r8vb9eBzmSjSaH686Svgbv/4u4uiKfofv5wNMCs
jZEoGVBM/LjYVFFgQgesOxgiR7/6dHwMRuUXnTEIJUBmPdC82C+yHcq4+GA5L/0q
2QiKkcs0XwF1bi+2me3o6MIL/FGvPzS1e63lGC9lPpmAN59spu3VOWmfONmjg0Mk
foBTgrpNvt7KGFefDtUw1up4iRcGmAwlVsvOIVh8PxeO/E8B+HscwQO47F1z+BZ6
EbZhko64DSDgem0O+55DoRrj/+agh6ch2F4N31HIyylltsDfJFkll3SjQVpI67gI
/RGwBffGprZWDIcSPzLO36vepKDquOOQTDVgX7uYKlxn/AiPCvAleGo1JN14k7fz
44k0uzbM5V8uCqhcInYeuPDqJnyZuYoEl5z+oc/fjeRwe3TD7tGAcrs2VZisrUOf
lF6pnP+Gnwx7FRTANUddjEsQRD4wRCB7Q0eRe2TxOXcHsNEOz/6jN6OzSPEaM3B1
GTxL2GV7RhPycOkTFQK3dBJ611Iub53VfrR3mVcMuQQYSSZ9yE4hRq8TGRuC05fL
JalJFifQnLaxwjyiRTE5oujttSKc2iQV0O8j4ZdqKr2VSz5q6lMa7/GFnHKSur3m
ar3HrAk7OKLh4TsxYTLd3VPiDEFzL7OPu7+FNLZOiNz8lnxEKaQ0EglmYibU5Eh3
kEkqX4o9zRBOXURuC2IEMn3fC5SzOVNAj443s1R4bRTjgBxsprVCCOnbfbMBL/AQ
blO7S9vZ4PswO2K2dbxI7WHbyFZFSIcQ3yGI76XVugdE/GiOMKprsOHiu0pSFB2x
3CtyGI8/nfYlQL29Q96JIeNmKoe8Nujw/0lvNLlAWdpiOZpmOLNBaQtptDg7mndF
UWE3bxD4l6s7GxSDvcmS70YsiV0Nx650LH5Rfg7GGPeSA4swvxa5ZvB2Cv81944W
nq0WX4/ONWGpdapA8CrVz4kDyeaQwsL772sseZSC65j1QvVXEqAzc5ZHCnB9U1ez
BbADa0J6Y+mWsj/nDZlV3PJb06l/a0be3SArE8b//APLwJpXHajTMHH+AOm+HmKe
0v18hGnsYFeMyupJY1P5Lod3S1ABD38jcWNqDLR9bD83vH4HYCq0duc3qBbXwnd1
H51Iya/VB+t7Q9Pj/yOKfOe9r4c/2YnpuCV+UWZy757pkoJiSF5MeNOL/foACJec
HBbKS0kBEytZVrlL6r/FHrDV4pqE0BTi658Qpd1lt1fdXQc3OzDBdTZSW2WHZC5H
Pwk/BJaqm/oWb+vB1Gb12Q5EF3vJDv0yQ9/DaqGuyqtkn0aNGaDMFVdAO4/51gEs
YmVHTAe309qHgoS6R3r5dML4Sz/Rak70fA36XBqtYw0a80MLLfHyy5wepPngFqfV
BeHmwfjsmG64Gx+V5xdqbNGTq6c8GkDuzCFVTjK6JDqFi1nmHehfo2qhr9r/vILS
q/T7JuDQpL6b3p54x02oSi53NwUO8wzBqevuscTYzdEMTWzfvWcf1voWsG+eZaLd
W/8uivXSRBPXfEAn4yAjs5R1wWjiXmL98LFkBXyTfKNnq61VeeJnPqabTmgHm94Z
8vKhtnxSk6rguc5+FGFWOwd25EfG2yqj2c/QZircFehE531ZAx8fZFyjaBeK2z5+
vlpHlxTz6wgCJV5vEjv4tEmdrLZPg16t8dxzuCLrW7ZSbZ5hg06Sav87wBAMDRtK
zPkt4fF2FlV3ABj+C4aujTp6zHYedv2uvr41pF2ppjkhuMvHeJZxzB4r0Y2wwF4v
TC6zLb1EmUZYM+p/chlAffS9ezgTc7ANGNnHtcOZDWMw0gN3llNFQHfWgt7Fh83Z
VD3INPc8fRG7k4M6PVR/UyBXktyRF2FvOf3wk4rvYiGh4uR/Fbho1dz9EUJ9yILy
HPoH52tCaU4PxA45R3pc9Iox5Fv9WXF59xDutlQNHOyKIEALyz4eBu9+XnPaauJ0
cx+DIi7U8VeUTQ6n8p5WqkBVI6kS+7zLuNB8DgYeCd1rBaVbogngM47OAjpQ4e9M
MigOQJu0UBnqJPmsl+5U7qn4yuC/a/QrT/o22lJhGCzGDieV0808aZK86kUuB18d
2LrUj+fFgNF+pLVDp7Bxak6DoLQax869llwvoh2nujOzf2aZF9N9EY+h5bClZbQE
nFjBJYVUtRtxbgokPUc2QqnSFZJbZhdD+ptPrLYMR7JGWbuA/Lk8ZaIV1Q3RQPP4
2LszLkogq1+920vMWN31fXdjhHas42Hc5blVunNEKZa/4LCGHx2iwvxF3UkOItBX
Qv7phMM/zkY69IotWt32FviWCp3pfCrFkMIwvv0cBa0I7qmUygv3HpgSOEKFpi5Y
5Vu901vWD8owXfIRWen6o9Yv1OGG6t75MjlP212FftNI1d2bFwOgxqApCfYbmrtU
z1+Woo68oZG7j3xfjPOednIWcUhZ7Mi3BjUVKR2e44GXLOp+RzJyeGqfvayVy9us
aAjkvYsWjrKyp02RKO/zaUZi1PxWzzGcX/vYh5zE1x5ViEYVc2SKdK6mupNMgtKr
uQBxAaWc90xUs8twYwTpR8uWW6SxIuTRRYTTgxbkSc4dSzC7ECGQRRQYaoCEdyxt
z3KUJ3VMbcDWwz3icCyWoZcy9T0Hrbp9RqPHED6yx8njlqiXncG+xMmiV8P8MhWq
kOD/5Pp15kyy8nBda1gtSAH67rB8Qa2gD1tg0NqUOKl3poq0smmZwRRjyahRjDfU
at7ui2kP0YPs5YUL0dcQxRaYYA/G1s3ydxPE2eZVy/vOEAt27bDK2QYYOC94fyF0
liQ54nwYlqmZXjvMfOi8MXM12F7yXG6reGJvc4HNP3Jsjj2edQTBUVJU/3+HtF5W
LT7hneFKnchRlbODFgbd8i+yWAGiZc70sSoVZSpY6F0+QBdmgQWnDs1gxSvPoYXJ
PqgFGpfCRw7nuMj8o0vTT/ZnfgwlXmFkZ9i56Rvun+mObVvN/n23DjfvFq0sLWRj
tsCRpkrgneneF442rf9/4HrwryiAxN0Pt4v9uK12stz4Z9L1zIo00kZ1sGYE1vI2
m1NZorjetfjCq3OxhdTMJZGnb8ZHg3pBmTQYJgf+J+3F9VDrTLLKvKOU3xcMy0fi
gWPXKwTKPamMZQW4GhnOdL9EheZd1fAJBBLs4XSGBwKukvyK/cx+0v3NCwuPog2x
pVi1cQAUtpnczdIZ3ZG8FYxzp73tCO77MM6sSoWk39LfcSivgxcLGuEjBJlM8wNL
mAYkHV7acPdf14uVhPFtblW8ed1eVHPkjRhk7chykIQDdv3NLr4s4zLCodVqKoH6
4dPlRdQn8HA1M/5KE773AeK7D+5/KRoHodaY93QMWuvAIXxSbQegxtNt0b/jS2LO
Eyg+JECM0EFKz4Z1iW+ewsLXVtbkRYNB4td+wMRsoGoDBOz8/6bBvyDkONM4vqAt
zJhidUFfYMBMTAAeYvl3Mx7o2h+R7ud3JIAQq4bvgt2oEr5wnoqnlurdTatDq+yQ
doRadGsqEFYQkh1dT14gc2Y+F2oq9FswIT72d99VocTQQ7o+WpewsNlp63XJLpFQ
p4Rim/NZ7v60YKQAilILsSMDplddtZ9uDwhn3aM8Diss/bsNHn26+7n8CbaL/JEy
h01O1OYfQzGDIlvA+ItQjw5GWJuaMKtKX8iUs3xzNRqGBU2+HllqvUJNVHsY5kcw
hU1jMAwsHtwcEfw6/0XAh6SOxDFqpTKbC+vUk5XE+5jIxdYwGuROHe1R8WxnHiHM
R7gZ/Kz/WLyOq4kgYxSCMpadZz5bHfiwVFck0fwx8cOfsTD33iLGOwZHMCpiWiXX
HDVPFdyikGPfuhSwDc/hZuKVuSLWI+qi+Xecm6Jn01N0sfAZgUWg7/1Hg/cu6dRP
9lL7uXxMEiBDEtqP5w09rvNjz1acaLZ6bWyBBpE7JOrXG2bceIZJXFaV1nGaHtVl
dtm5ZU4ODvhCKmoG5HWn2ScBsiR1mS/nXcY8EtFWgXI/TNhV0kd0WD6r/TGZ4F6B
SRe9rcVa4a6Uma+aCw3IQPeTSFrjcOZawaLY9a1saQOLfm9/4BTkrcCX0XdMnxIk
+J4ZONtpcboskR0uTe8kAYrRG9zDktnKM6Q4/riJzZYE6m3mqNWJAZz3oqOq4+sN
tBPOlKzt6rFf5VlQ67UqbNm8ww3nCRqgykJCVGEk3GFBR6RpP737SRSVxr1+YCsD
EMtA+ry8Gd6NPINv6wzsU6GqXSUfE+NAenL9d7Mp2u3dIdkydleAGUT4TEPgnAq6
kKRns4AqKdg3KuvW4127v6xziGx98chsXEcTFrMrAG8FK8uAoNbcM8D3P+TWgCss
NTJHSTY+TCPSTOwPMWlrxiZxWFFm9aUOjXGIuxElT+I7DfReDqHL4mF42hdh/RQL
AYvP9T2uMy2f4jhCM1jDPp76qDCandlvsCCJqbQeEsn1tspGeSbxGbOwCOSGpadk
Bjf5CXpy/qPUgGZbZrnGMHlOhADTIZWJNvX1RpFc2YVbB8ztJHUfGbZ+03Uqkowu
QK6lmCynypEq/kn0gnvheSDE6LjPr0tu6ZlS6ks6ROInW9Rxla1ReuoxDSQrxg83
wXRISvu8wU+ab9tgVEDqKeOMAjl76bpSsii77MFIGNWNo+ZTDY71y2qTHq2ufF27
4wQxfP3cam/PrBKcQGMVwEOKH28ELccTBAjjC4x/UzVpUmP8boVkhF9k9aDeYXWT
ynkg/G4LI0tVBEhTm3KbpYIXN8lm6xv0VTUmA4H+v1PKXVCfjFxoE6pqqA6Lr1Fq
bI0sNjwBSupMwEAXq37SHtbcNG90x0sqcunLl0bN1VkQqoxW24v4GKh4JYRXGKvj
eb0bwM5gNIV1hCtp4Mg0XLHM2uqvCelNqOzfqCgV7Zm2a9jlNdu6hFwuFKNcaLBH
wY3qM2fpS/Z1saMHUY3l29uaDVr6FRne+oxGxC4FV0hS3js7TVEAkMezV2vO0Ypa
pR9GH2tjmho3WXGixhiA3iVKMfsuG68KZ2RJzWjU+O0v4DKVejpVaE2ywY6DguD3
Hdj/ko2EhGilbUIX6QeFAMM7AtLb17XWXCN5HLpaSziBGOUK4yKoeH6/WsDnvktd
X0xRmuIgAYdq6AZXb9ZsTLHOyWfgRfgZdB3VCGv0AU434Sj14ZHGdIkXElT3iFLV
xyVy6yFvC+CZ1m2/ZQYqJxEMetZcAmPylB9PNnwNoQpNSyHj3RKAn922HXccTHIf
e9eCil+vGqnD8hg5p5+4v2wII2Ubsa2WzxoPobBIYaIlvkghG6mTBIcvBD8msvdE
NeTOXWH9Nl157Jtzdrap91E+Z+xgQZLXrBEnke2qRGYOs3im/y5r6HIOXh5pZGri
d8faWmYTqO2Xoo9unYO0U880GZKNkIVi0BPJExfxB86OV/mbGr0jBBz5+Y3/1WEw
gMvHujbhbIUgjNR2OnPqzFL/3Qt+UpzeX96uwzrdJoLokdpUJo3B2099E67Z3gr2
8wOHbYy3XqUrLOCXJmxKayTltf98C+shJZkz/3FCzwc6XxzNJz87tXCAxAaShgJv
c+G1QcZzHHpA0AH5MtpTCZmupYya4i4dG81BymQR+qFrkvJ96VVx4NCQLhqIgS/x
K+OKbSnh6/dAZiEAQYrbkbFsT5ZH3iAUQaF3VSmMtq+HcFLmznueBineBVx2BV+s
Y4+06S6He3UCoO/KhdH/jf7wBJbSDeGijVD/EY0XGpe+Vc2W6GYdCb62NsdDluGc
az7y1xG+zJ3/mwxvwnL32Hlx7OJ+iKHmqH/yU+0AqDlZjUdJ9mmHTBezhy2wWCxZ
d18JYoZ489tbndN1MLjU4GQjGcL9GHPu/xlDI6G7+9oAlv0iZgO0WXWC0kqjSpU/
dzQaoTSRcsFlyphRUEh7GWlsLTVPZSrP1HHx0IzENyaEkRWPEPFZwFhbg8A9KoOw
6sOd5u2rwB49xgfVpgGWwvOAQ6APR4PtO5BQmQsrSq0SzwZ4cHVd5MQg+mNLfzzK
7sK3bjo3I0yAm0A5Q+3i02UnCFtysGqq2W54TOZI+zrtIPyhlaFsI7RKS6pFYGCS
OknAhVE/dYEkb6WJP4HuUy9n/NJOUqgV622ROjUG23uhNbpDuKZs0WsheKTNFnJb
abqjpmIcfHJopGI/xrqvmhxPPFAEGwhTWk40CQtJCWj4Wa0emVCgnl+cwsB66RMH
Wa5fekUwXsEEB/elxl6Z5W57Bxxk8LbDOIhA4gh9T3xc18ew23W/FN/cTmMm3tjS
Yg0RWJQ6FAqDYgR0MH6fl5YnXNxzdfXVgRymwQHjMdSIWMPaQP10sbSiRuVsV+dj
tBPcVmPO2v4/hGkgtuc9uPIaDJR3HmOXi/3Iw8iJgtpU5ZZgqsob3R3oaMUyF33N
Ws9zjY+0T+MRwdHiqnZ5Bt2pjRprp9fZMjz8+fnWBx2WTqGpMmnLiv7NP1r3RA6v
mAZHNJm7bvxbvxoghLT2UegvyXG+dLdLkJ2S8+pyoLkGETQo8nX8RwNllcl+XILo
ES1oLA4gSn7VFzZ3kjiCYepdpmGbdkVNm3Rb9pcbZR2K+j/b5vvvwxq12rPVQFiq
RjrM8r28sFSAbKYucHDE7MP06xLQbXMaoMXSsFpBbBgcJSBzttS6iqEqwLTcBHZ4
kM7hQcOwqpgAqfO4Y1e5HNs4pnCa6OSXw4FDJs9qenI0b3AWit0/FG/14wXwG7uX
nqxmDWZkQ6xSCJz+DLWaQryhQzyZmz2Zja5fVYplnXD5bwk/3v5qm9pbsJOpFZou
3nfIvNLJRgVrd3ZMgWRWOBLE8nT+HAj4FXcDIN8VDIx642OhFESiXPUIGS6ef6b3
VpVcEZIrzhvHlqCU/bIMmvjE1NzCtHChZLQOQ8Ke4TMAr1a77oiLtpnyi495qmp9
Vr5wO2VVttaX1vsyEMk+EJVzffrzDGQ4P0L4eISpo3EducvMHg5JATHVmCrrwQuc
+8OBVSitRXkwktBHw07SGyjREQwEmtE5xNcan/r8Dn+D3ia4PJP1qz587etIBsY5
krj35nc6wlSWEQgqMw6l6XebzwhbA06TkJ1WXcPl3MK2eQmaphcTVwUS3BtBoPUh
4yH8rVfnjEHmUlnPsVtwsridZMYyr2jrahqNl9SIFFqmcwxGDSeUOVn/gdBSYgPD
+UNCZZaqjHFdMAXGGUGRn18Dp8Sw6WfZcu3C2/yNFQOnZY/vyaYF+fXFR3+75uEJ
7KOWtrf0fLTKTg/7iIRukk+rYmWbJUSi+onSglCcjlR53yyDW1deVvugYfjrk8bx
FYs0+GSiSGl9nSzoUCpa9ubZ6gvL5Xlw/8kYBSlevxmiW5clB+kASmNmjtVtUkcl
Ine245a3VRniwXjsMQnv3XCqhODS59A9RJU35ukeDcHx1XNi9MdUb+PyUAjxgHi5
Dqqlaa0dHpncC5+uwvH+bFcAdgJPqsR8+0bVw4ZRKxieihLAjTUZ+krNOBIqT8uL
1RtimGB0FHpxDF6G/sIhn2H5ZGC9+4PbvCaThKe8zCILUwDiK3loHDoy/brYsvWZ
OxlX+yyounaONqVdchqWby65LYjNnU5u/9hvK6TgyPahH3WqYiBVs0qUH75Hde7A
rzdqCB2fYCjzN6FINyOSfvVArqHRSMJU/SbEjqDDdLaBlVw3UfqmoNc/juSnkV1k
7/GAGlVdrAl0pkBPe8taErqlN3k3Dy9+8im69b/4USwxztnu1UCFFBGbAMWc0RaT
3TACYb1gjMElkKt1jZnyHqy3kSpqVM8XPsWWh1wvdKD2g9qPNFDdPCrq8BqjX/m0
iyYjnF2vVlKaUNKQaFET7oCh3VS8CRsCQfzLlOrrAf3KITzTop/grET1HaWfoDUL
n1JngSpyO9nHJcSEb02oJAwL7+B2KY611T7AppYXW3fLgBXrS+Dqqqs2wimcrrMn
KBs/HqugY4R2IfZig7jnq37Ujyn7vCELCaMZ883ZoXat8a6A1F5tzVrO3W2iqyyC
niSAI6GyCLj6020315d8CFLgEG3fJAq/W/cltAF68xsnEwTo/ECNCkqX9lX+o5m5
GNgGPmXi8rPYPP6Zf1bSwoDqNMMHOEISZQgJhxAN6tYfGDKm1VlKEW/W+1EUFCjW
CUjOkIq9EePrdJixWU/QnALQwRfkYkddJcwU+3wxhlNrtwK8+gowhqdf2mOYYCYv
nw/CX+7xw+i5jyqvaU0gL8gHuPSPmcnWpbYDef14unTMuCgQT2mKV2s8o9iG2Zt3
l2aFGn+B57+hiE9GQp9gSkfSiXEhk493XMpdWIAoygksZ23mbmu7s8ZhlECfq1BR
WcIzRYNWUX8y+GRt9ZZeRtOQN/78TaJvdEOeo1ERALrSD8k8DuBo+nFH8DXnfbw5
B21c4IE+1qnc2f67RGziRCBZ+oSnGqzzUL1L3nPCznZtNee+qu441qYGidZsogFJ
oWmcJpdUS+Zkp/JDhMBqyW/S1M0P2TDoFFdC8H5vkZy0DVCEKMkvatviuVCDh3Fw
rYtTpFLUOSja/soL4PfLWWKZojS5wnb96RdjQl4J34iMnDSlVeIKOE2BMBfBs1u+
wROyCimteOE72q1pGBjnhC7xvfV5b6RJrLZta+wXsCj8awv49ZdXESnv0fz/cZX3
vS4MI4BtZZrAy+WD6dBz6um4O4cy/+K43oHEGOkaIdcev+DfLnQUhXe3j0vCVS4R
qpwShlmALMXaWpO8HVi8kwlFOeY0EJQI84JBt22mijyrSQ5t5bnigy8hTo332bjz
3XM9ndzsvPUOYBDpR8bkyWXy1+S+GEu09co2h1Pe54Cqh1uziqjgNCRowCRabVwH
AtF3KH5Q3CoKsXYkXFEskUdyGZOZPn5C+YDtCUppi12Y3VTvTGtcGlYXZWujfSHQ
AYOfBNKPD5yecg0yB3uYjpfUwtvOYonGXnEx4fPbKC2olfpyGIIiUaNRwDVhYlnb
i5ukjSlplGff5IsdhpM2c/+saW3PLRXhngvPobrRb2IIYwp2ZF3FUfUxwF0HNxWD
TL8E3fNwIEh8ADkZkTiCgAh2UFWVt03N4hDkQsoS9GSxVRkfO4iAtsIIPaOmdptO
EayMxNnB2kS/f2aHAOdzfslcIEBr0jpTo3+L9Aj2gFifuFiYAlm+QM8QTrUR5vOv
Lb07ODDXL12i3TJ1YpxX5E6Ww9zEErbkbfrBnXc8HkmIFAsFcUYGTDt723qnj42N
HebYvlWYQOvydP1yQGt9bbDoF53WrC6eQOhXLii/+6wlirm5TzMJRTdoyyN354YM
GRNHefUi9gR2UYfN6PBa2meCMPL+blPau/NHVnIRhF/yCjTt6/xZt6AbGglvRM92
soWSYNYCfmk4OleK5hVJWn37C9UG5fYkFKnuR3nkY+j7cxcPOlLmAC+KS5Cpsn37
Z6ZnzSluRoNkA9MCJS1otfeffeg0AzGnPpSzT9TdvYSxawUOPgy7PDG4csj2/AFr
iViZU5UDQ1/muZ0NB2A32HXMcnHtpGz7t4JavBknNsy76VyCHM9tPpg9MOtJ1S5M
5C3Bf1m/r1bnj6OZIH9o748EXNz5zSC9eDdwNgaBJ4L7q+34V4ugv/Q2zJpQmSYh
8QQ86P/30sJ+6EzGCeidtojSOogyFUo8bL27TSgmy1jXuz1q+bRtF6lGz63plhYh
nnxOyJp7ZhvCe9dHjc8WVG3gikeo8Ejsvq8G8j93eNJhN7IN0OotNnIOG6kftYmP
92neeTaX3qaYVYSK0mF5StQkWp2PIgT7PJfCCmChT6X5chgErRVAenlFoGAmIGiQ
vowSG3pz3rSlfEM3Oi65lC2xtCztqKsArXrWmUPu6co5qO+JHW46gqzWEDRh6enJ
l6qW7p6XW7rvrXDWJhAUX+NYFOsCRzxyFuId+n410HHc1ml8g7oNWyAyc+i2Gm5b
3O8jB3P1mSiUdrfZ2N27FeubWZex6cdckd6CJ/CM9qf7nXlA0SocPZg49/g5efGp
kEJsXyo509GIuYa8njH03UZXr7DIGIdUjxWjzzMRyDXLeTI7+XmeV3IGyWJUtkOt
L3Hka7rWsDLF2CIZKp0j+QTHrnO0odojGFRG1so3LvhlXLbS7TW+ms4X72cV6l2t
dmHiGxuJmb+6FFdQNASHUWbuJvyNJ192DevHE1ZAmoyyfMvEYWfWpRZCdKtmtfJI
qd8suLgzGFLfuT22QtulD4Xa4kKHJcGf8APok7Rs3HhV81Emcmy5UIsE3wyypsm4
VcWL013dAE06SR486rSxAZ3XvNxsjS6zEEP74fyWrtB1GMjuirxCGooprcYDmoh1
1JhYCRyfTJR7PfUAW0Tbtj8y05D996cqq3tekyBQl1fFBYWvTHiXCly0tOVxpkkO
nyvdMTxPAUFsK96DvfRAyWbNrPm0e3uCCe2woixoYLcuc91swpn89ZdGSGTNrzqb
AbQyB5ceUwl4NRi+5skMEkCdCdxlw+BOc0ilY77IHxEO14SPtMUd3wEUGNyVqUno
vNPcGQbUeb1kPS+ct/anD0ygOR+Wlm+sboEij1D91Ny80o0ptKLoaJVyHRiamoTG
KcGztrRUftH1vFgp5gbjLTKmPT0GrbaxjAi91qbyyTFL1G51gvVLK59iauKT0cFs
30iG1vVH7l3U3XDqiPyzsY4/69QiKOLwWiS86N97WwSz2bSIe+dTLuQMAJjKutOk
gnnkI4r6y4i5Vf+EQ3nxUgtruVGAE4pNlx17vuU1aNtLJ8nsApL2k3BTd4rpsowj
moaZPU5q9IBtq52KqnXM+zBfvZByacPNrLYXZpwPPnX0oH2WnhZIt1F+Cdzgg9J6
NHQBGP7sWPTykV54qXZPezT3hl9q9HMVvdLal6MKkYmI6eC9kQI5JUV/HoAAMz/e
7IsIX9r8nt3fRXftj3HIhj0eJ7JRnaGTDWw3UWKCX/99ClCzBz/z7t9PiFwH1xKx
ZqCGNZ4lWW+EQz7qY3Cpu5NmyfBQAKENJUDwFFjIY+Gync2EtzhKRSQ4RgTJVtPu
AOROqlxrcXi2ZJcnSyfhJax5Ytz3/dSi93tKahFKcG2hoJA+lO4Ho/gv0ppBTn6Y
VVvK9ieVup+2upzfx7J08l8nP5dJO1fhWjlEKYq63q9JxjQbYtvNKGqFc8qQq8kf
DowRfFPiTjFbVcNaWGRf21hO9o4rXxHorrBbwNhSw/OX2MnGv/lZeYVXekGmcSy7
e6U07YSvypz8fxkChq1GNduLUZal0gPk7qjajKwAVztLvnLG+JISmEdtlzFHwini
sBTb6yQ3IMqIyJzFhmnJmOcApmbSYgtbjRt2EtrO50RKZLbN1uEMyEpLku/ag/8W
r41gOU4kDGLRYgFoFt9ZLPNWREf8bNWQha5poyQjTCQ6LBuWU1RlqWlLPFqobSjM
LD1UFxnr8mdndN5aEPst3/KTio7QXKyBBhJmvCQAjash5kYYFnemjtEAIEETdQ5D
xy5Mrxe6aIntIw+pgjqyHdO+ylwWXmQRT84uRyb/w4aZHXqsxvj7pr1WHJiUXYLO
8P/XFotBH2deO/B8aadhbDSKLns+NCQ88Kg7xvQSr8I8xVdQzEzxjfOOyrv/XfyW
TaYEi52Wd/mZ+6NMsSHFnJ/lSzgmrTFGThEruTlBqZFPyh+WRgf7FHT125+0elHD
WUsdQrR4df9xO3j0g2MumE7IUu9ATGylxTFhINrQIErPtNu2545NIeR+RVks8d/8
u91d5NYWqgaNkEiWXUEyYkMqD+wEcfxivhgmkc5VdHsDRWaqyF762TmJdFaI4jIc
S+yO6YOx1i/EbCls7Wl6IS7FdAloEkmN5Y2DtqVGuNqwWFbPhZUViy+y10Epowdr
raM+I17Kgo2Q9QZfNMSOqPMKdLMIaW9qRNqPDh716frSH+IT63j3YAqPyPfBzu2T
tVoRmRTQATtTLArW8A7Q/2CiN6ZQ6vKwQFCVQ1T2khxqxvjCBTsYZSGVWdyb8Pjl
L5QsZAcdcepGlegpCKsSR8WiUC90QodlPsmIBt8asICNjb/+oIR6pWcNm1gIGjug
tQm0poJROeMB8l+p2fMmhk2s0akCaiZwv0A7pwt7tcTrPi7bRGFx2jc9vRDS9c7p
TGfmZTpGht0A9gtUfuQUlZDmUdct4J8zp7/CwC1Y99PhkzGPzTlbKHhiW/hTGmDI
k5IB6WjrBRt+eiOo2boUHrPX2q7XQowFDCZmjuBrpl34uePDFOxyh73Mgy4Qhknz
/tQPlsMDK+pUIQpM/3BD+/ipKyQx79wyClX05wvMedeegZ4ZdLPBkTrooXNslquh
kUPM39L/tyBHbJbxUwUaNDGKqcYQBdnh1vn++quO1KqQzlYtK8hFoj03MgVTofkO
YqDLAAQVtHkAq9VD70ce3d3aFkXy1dzd8DMxiJTgyxVkj7kcaKcSZUa3svKG6msB
vrAM7dJdoYxSkUERLRBrsuRIeGfzyUOe57Sm6TAHj9cLv+xofZnkOzB2sHsDVMuG
LsscJY6aFL0exsyko0nalQOmQYYxeL1FhyAK3krdN1T6efbIQbeUvY1yYFVOBKtz
ED/u9zIatlVyDGodh9cdqFTP1xNzmgFWcxlfBut6r73M+QBcRZXzOXN0oJSsXjgV
FkRz8oryKkQU8AeNQzQTcvr+a6AQr8JF27qLR2kSCQTC9AiIwYBiJV4eY9LNwKRA
ZVdxjB/5ifGlZSwutb6C2ECutxDZri0zIpGl9uG1JE/X5kEuJHaEIJZovdQf/+RP
E6ufuIGcnwSAiJsQ0vP12Y1bZbO5VO/4Qxrf9K1Wz4I9uFtcdbORXqIPTAKbT1LC
ENIu2NfMnaFW0RbFrqMwR/rel/48t+5bDFjPwnSydWqJd1BeJEe8IkQYhBRClJxD
3BdlhRKeESyhFvDDbpJ2XTwWivs3gL3TRQgQd4MzdigrVzVQhx7Vt8CwltXpJd3u
WTAW7irdAo+qZyq2uZ17ycPaPl+r698kt0DvCe5XyLWIJLaBVvREt/kT6Dv//Wpg
3yHg2UQ9frONL0MrpgaspzaEHovLos4gTxLOqTA4d57GIMXJqx+/iH89w4eJXR/F
7x28vdE6WnxM+ehh64jXKoBSL2cjR6sFg/FbNX7pnAhw3mEBXQXebgN3hRZCKHup
JMsSgpMlfq3QQsUn0YAIVrP6SF6iE5ikLldajnOVcSAf6t/Ytrt2E/DS5piCydKN
XHxLY8qLo6YgrEP+Bq3AYPtRhzjdbbpNhyTFXE3zDnj1AJS2FeZ2RCEUcDJ7VQq+
QKyqicqrzgvBxa3u1AcRSsOJJ6Ya0p6aIHrQpbgIGOukJo7AP0DMXJJD3+WexUT3
qTQ8MrdvfEr5TlZG/K/usUbchWwOQ8p4pFclSkKhEh2/C4IOFW9nFOOxARs4qVCJ
KnrkoIHdyS6M5ZawtG4JlOz+HkKUSYWm6tdVvbTvMxv99KheI+VONirqkqnfcqJp
Dj2f7FmSPjbYw0yLCEr6pg3pOx6wxRXcioRSgB7ZgLhFXW4iJdrloQ7cJPW5EMZd
fHBKvOvhAbDhG9P6Qn3L5MTH2aYJlDS/RcsFbeETaK9avnykcPIc77dOr1Lt1nVe
Fvt2rGeDG7ogctFY+egvcT+S1vPASKHpewNq1wWXT0DINQ1YTxfbcJY2QFEoNuoO
nEtMuva0OkzE6bgWVyJtcMGDnDF4qLbNuXhvfvzwk3/cmqRFIh2TfVFfIkVNWkts
uqFfOeYOh/Jv0Juni9AQ9zDJBqGTl5102JlOU/Akvk7aGHN7JYHNWSvFR062JAcd
/n8dBOV43j72nmWjAH+iNkDqw+yswzzURBvaNwzMLecHjeo8iGcpZYSeORJme0V/
WNMPghfjVGrz9bHUo1gdwgkC5mTYgfpNaOReKGFrI2QvIETSri8mOCyz3++LAqyL
3Vuq83UQDUPfzpB8aWSLhd8KQnWOE+fVOSRgMzuBaziONhYGUuuCWOdt2od0Md7w
QJG84UbivSRchO1bJ6CbNiHmeXk98rwl8qz3J2LP8i0ZdMxdn/DNqj/nKRW2z7JR
QKMGtO506fwzN7URRMtVmaFpL5F24w/sXEKMDux67o9Kll/JKsDB6JjlAAEbr4i2
9hvVCVfUXemQ4rtysW6N/fSvuPl55RzxR6I50KIjDrcG5WyrOfKm3VSzQzQWjrZn
Q1Tuy+oQAMJRvhSauKiR+KGESd2dSxMJ2AH0QeN1MvSPwvzzNpjkmhkqoNGH+4+Y
BhN3t5KLZdAAtulzL3ZEO7PPvVlOzkw47ROKk1R9SwRAwS0LQIbwLAwN1BpGQ+/Y
B5FcEeSJirU3WiXYqVpbHWUegMv9slomqJSWswmhiwfPGzHa9mCDRBShVw9ed6wQ
uCGTNJiKK4uyfKH3v2J5WGKo3PCISE3swv5ffJPleEeoUFXbtnZisBY3XZH87OF6
hcML8JP6dytbNOuUf3qsuWn+jbn665nul0+MrhY9hb1l9m1awN8Nsgla2qY69xcc
m9BsFU3p6A1BOVDp9StUmpfvnRZX+eVr6xFSrSAi6MJcgIBZK3syd9hv4riG8WBL
GAUdBW55NDoLxFTjGEuzYktkiYpdzDAO+S+LR+1o1f2eM/40kCMY3B5v6Vz7WVWR
6x5z5CLqEVjq+nPQg2Svcbk2pJTX4i1s0ffhn4XiWSjuRSRWZJlXbEAYbCaqKacI
6DgMtK7htHsTozysfcfRmVh+oC0HPXFLnXo6ospBwaCDzDOROi+BY2n6ic26pbDr
hnJZE3I3WwNvMNKK0FpQZ/XaypHC03agO2jB4PtbGLXuIdAp4WUyCUj29fvu17kW
wEK5OIy162nRGxIVeTH6y6zlqSr1NMmzyE9vCbGc6ozgEl0YQDh8ASF3kPqsCq2z
WYv1yMN9NZrWgSpj27nhni2aHYi34glYfNaIzn+4lH+tThV8PhiCatFde+BdS9Nd
OVt4i60S5bZqTLrILAt1HNHo/t5O4dXoR2nafbEaLAZ92ZoBRAVK9w7i0uTjb5HI
Pzy/G4O7A2NUPgSixI/TZge3Uw7C/Gmmcx0hGv6LjA79HUF03dtQtXqIX7jv0Fek
t5l+P/6o59QSjSB16p+zOnaaULvNA75LuA5VXCqLjaRTBrVoxxZdavbnI69her0d
Y9sEh7HykNko7/Ah4AvR92kIFMr92JiXYGfeezQvPiAnR01OnzRDKmbW5+mKYhB/
AVivhtKFTBtoBLscjx4ENGunUKCCFsmxMoXmreZs6CnUECzeXoP0HsPQZnWs5LC2
DtkynQ03ovZM3MOCayCcHs8+RQcWUufODhAq+tl+E1VNDp+SyZhXGdX4YpDB5Jv4
uFWNDa0iMj3OaMLT9ZZhN4B/gG7KXmQRjRS9Abv16z+nBW0P2NxYlb+lk1cN4zZg
OBygI4fv6KWY8/lp+G/ter8kLGGUP2Fes/HMwWp8yOqS0BinW00YKh9Z67i8OhEr
XqCrm901B/DxMA2CBxCUPwBTBjr6zB0EVfSCmwgQd9jBdzU2wXTvP8NOOO0rc7s6
wRlaLJR6yGyATD7c0ktUeKS4/tonG7XQoOmFCADve/A/l5ExCh8uiJ2kBBngPJpP
IwZIykxej9fZDZZQsVL/aaKxFqRb5YbCIPCTJa68+bIC5RoVmlSpac1zmbIi7cjC
XAXLPrFi7gAm/O47rWhoK4BmlYWZQ6QpZUpmdEivDffXb4PuDJIDYnbSGDTod9AL
GTntJIqn9dqgSNMctlmwNM+EWZtFkt17WQ6KEUvPdcJnC5BUwJk5cDLPy0Z86aFi
kxuEKh2EIJW0Unngoo+UwCDz3GP3CU+1iul8wlzVE5M/kWZcTvpWNau+FXjbATh+
N/RHgkq6KbP6xIJAKIPu+DVX8crbP8WDys6ZxnI1rAelcT79uma7XkCIvbV13lFq
u2svvDyhSMB40WJf9G6KswtANJLZvQXLFWPwQ9mmn7eN3iwt25WJ0BdhnxNWVDJ9
qsxV3N0pDvxrxCinJSg+YjV5jG2h7zteYqhaHt+t08ZuL5G6ncdK1n2Rn0A0Wf1O
IkAgIoVBnaABdxBEVDkg416TFq3yiIoYJfBLJP2J1wIGvVoKHUxTfyM8yK+YjPsA
xhXfeIqhwwXmue3qStQOR7w4CNAAAE1c8RqOwVw0ZZpWcuTICMeuNH1lfTnFkDKn
6N/MbFFrqcJ1rW1DE7sfoX5hpNlsrkEoorbhHkwMe65OFsC8rFI/A8vO23A2WhCE
sjjVHWAs+CAs/BOqEF4nB5ZjdpBALLfFhJaQI4AyxTmkNZcIYjAo1jocYZubOxC/
Ko3reVB0Lv6Nvj4NmfhcwVB93OUqTp5whxaDrPZYJWC0xa98gWDCurf72D5PC5YF
xRkgH6/uzGQaIxIORZCD7boMxJxpSkPaJ104IHCnPNajfV6vB11XxRC41EgdcyQQ
A9wQtBexvf4DPDCGrb48apZ4bWY2T4JuNpFCrfu/o6hrW6G4XkXu6yK43FwRIV+S
AQaIeso9CxafdsS0mo24EqXyOWAZYgY0za7BXKqOALLu91mXxDSmiho2bcF8Dx0x
8Gtx+cswIGd05HP3KiidXXosh3WQ1DIR7/ZVG5DSFascKdmXVWnFbR2Bj6Xm73Xp
471qR1xDS/9YwQvjOd0S4J25NQ7Fk5tH1FL8flqcBCxL5FUThhYFqQIEGJFAvQI1
/UwWbd8ISF5wtXFbZ+WR64gfPFsrXp8DeFJc4Iyhest5PZei3bXheYmfFeZNwxXD
BDrwzKD/8mipr9I4Xi3tjGKiuLDOveFc2VJTbvGZ8fDM+SsOvzGVUvWuwLqulUDi
HSmWr83r5ch5815HZylxInZ5ZTRMLH0n1r0/XdTkpqDpC/VJTlp8ATMg7nFm3+8S
FSd+C4tk5rIZgeD6eR4Zbl00uIGpdZv0gLciTZtJ9WsK9eSP5q1tDSCzCp2KEab2
OXhYy8nXfqPhNbKIbCHIJakzUsaPXf3yBK5mX/BbthtkOy8vDjro0kgzGSGlqTck
y7ynzl4jeVfYZ45NFneMdlOugrA38vNaAGpe1XaRuam78bo2K8uJpJ1u+FoNFl32
8TVwbcCNTpARN/iasmedrs9CjTD7RST86wTVrma89r9N/O2+linRpgDXK8tQ3IRL
l7ZF71ZV7jC8Mr+3KYdIB3Q8U+0age8Jtu2yU5JDNbqtf8s9hRKYcirdoymFzkuD
yTE0SW0IQ5erpZBn3CT27H5jxk6RANmSw4CwskuX3xoknxcFi++9tG3YU59B5/nC
hYHvhuCFs7D09glYcKvoDxRnLtMfF9NAYR8Jyk/rMyzCBNlOMg8ZxCZPtXSV/qmg
D7EKROaLOhfGe4y9Llf0Orkc7oZ/d4VyzsBCF0l2CGm/w/y6fXf2Uq0i1XcCv09V
mkSNnCVdFBL707C99KHaVU+cHwRadNCWDVomi/uUwm2BpHcinKxhccCZ8fAjo2bt
JiviNfk6KNMY/ORLrIED2bldgwP47I1B1QDYczsZqzbqLNeSeDihvZsb9bOMZHMe
1vuieqV+iVlDuL5NHTEb5KoRCLpGmhszviaev6dwW+oj6VH2aqMBVJ76DUhihvd2
e4Oa75hlhjZbJhiniSnjBQZf7I5ninOmH0xrCBGUQVJzKDpNfBDzb0PY4b5PNAQP
je48h3uQMOwtSPNkdm6pi7vBD8VAPG86T3zVY9+1m4DrY7ZK+ym0K+6XLfEXwWfj
cEGGrWfFTxoWx7uIl8i9zIv6TYER8dmA9rVXJN0cLGNCyHmvV4i6z8fNx4g4e4Hg
XH2zHl52TMUyiUzdxp90Qyx8ISKKshvtLNvJbiBlyozHzDaDbTK8hTu+R4er65KB
UmKUf05iefqf+CsaSxEaqdIbEtZISU/ygVOvDl82iNcsZuO4Hr95U/tQkPlSjF4l
Z1rlTx2MA090cc/VUKWyh1bLuGWLTv2XzjCZhlvpN9UHHkj/FBDjI8FJEQYuWmLa
dFn9PTpZnNB8P7dRCvmV1EuabBnqz52gSG+1MGrBPfCDOT+e9sWq/wn7bDEMEpoR
XmbgdxgaIrdr2czMp2Z4raRT1up9ZwdelTsCCPS0Id3RVi9nCyaWXUTLvUXTVCkh
SnpMa7TwZHwrzut0G+Qfgg46MIxaFTlQCCNamYLBfwIK7ZIxTcdRivj9ZrZauWWK
xu3/eEUj+kM1ny529N2RGy+0GUxBg3ZbFguvnQRUuXTaHIhnE2U1jyDHN5XbIF+Q
sgePuarQ1LtM6xxL0tm3ZPRfcZbmzn1IN4TPaNYJviEUUGaye9gIp04sobnV4tUc
acbpCdjfM2oz21Ko758CCVrJESD/S4eHdeT8XbTGoDnMYRMWbrLEszOHB5oW4YJd
t2QZYa1UY44pNwV8b5c4MszyIns4AC+WMJaNBfSGPD080I3I4U9vqtYDXuJZsu+C
EqIX4l+72qSGzSm8Y7/CSTQ9gQ0Ltjq5EG7A1yaW25BDZyo/hrK2OOtZePj2AHIz
wT4SNhuwyfeVr+asH14mRKZPs0xQBdUoJLwGtfveyMAoHNHaZTcwxGee30Lf7+zR
wQAAzHtCVUgKyjSVGECOb6+WIVzWOC+h+6A8pgQHrN4ipIlUeCHGGDVjZ2Q0pnAl
GtUykvnAM+jNlH3k0E0kYp5bqposPzUVq5XAuY9zqI2y/O+yV5M2HUWw2gI3ReZA
yT1hNW4euJzUxUF0acWRkYRYABw0QuFyv6sv1my+jP91sc8zb5FOSYHi/XcwyPSO
zFLqYhV2masDaZvc61UfFcbJsDNZAjn+S6B+cJc3LeSG3t+OgPa8S1tJY6N/wNau
9g4lQaPURXkraMM0mjcybcs+xxaptaZxYNUxCHMJ0e2bvRu70mqbaglcXPlpivIr
TcZ5H7o+Tg1EjHbnn4H4rFSgPgH1HdeofU4aIavblECFj6mX6I0CzZOCmFj7Uc1w
KYylrfQfke9kMGwVdePpTuP7n4Vj1KmD5eKBgRaFJ1A32imKJUGYwVggjo5yQy8k
eGX8wSgoEdz24C4Qb2TfJa8vg+sr4NO3jVAXkkIELPqQ4qlpHgAWBaS6U7zltpB9
R9yDiINy72vl5BRidKxhbTj8dMxDOlslRkzhZNiDgaIA6FqjHfTovKu7wK69E5Gm
jUOgrxh8SEuYQV0KIAmhmEtUncGpYB3yGaLxFgPumOXLqgR5Rz7ZwnQDWtwGnHiH
IpndddfM4GmMyQHT52cR7mvRx2cG8b7Aqeb97ZZW1fIQ1Pks+alLtMlNwq48ihTU
+mIl3njrcnR/cCLXy0J961OsqwOwN5kx87t9a1vGEB5eWnsIt4HnoHUlV2Nvjlka
rkWhtpCoXZNF87o5muIppc4sCGdLEhcdocY5AeO3P+Xv1yuPasmWytDThOtv7Ar5
FwnSxs42dRnf9UmwNb3315MDVtVBLzGaVwqexMHiAS9OuzxK7OIHt5jvDtG/5Xp4
GjufmDs4lpSi8DysbxtRAnbLsUgkfz5E8SpiNIrZqiyHckfu4+JsxlU/uDERZ7Ym
TnRCPNy0yy8/PsGQutP67wihFgTHRU5dG7m1OULRnD6H5jg9yiWtKivRCvxpa22a
6NkQ3BszpZh3IYJZl8tnsV6CqQUMC+NpdoPQqT6BHpNB4YWJ5xBE59MiexMqEaiX
kW2wjgL15MTeVX8BH5aPCGNIAYndrpHB/qacj77Teh7N3/RJKFmQaldI+e8DmrTv
Xg3mR0ZKw0r28UE9Lqs5l+slhtmBkUSI6H3yICGrB+M2jeqBIrgFhCO+R384Rhys
iPYhW5N7W7gLkdj/zhU8pd4KtWRVJGgBw7lXaZQvTFiYDfNF9duuWWCxFeVsWoG4
APj91fikMlmC5gnAV4zV55m5wMt2YZ3dKP4DVw6mxV+DUJhPC7UVeJvVg6E5rojs
ieWWx+8E0Wz8yOvqpys3nzvIEe4QZQ85IRXu+opGaEKToBwowGlrUOZJpN4z1N0W
JaoZB85s3+UQgYTxPXLnk/s4WpQPgWY967EHMUOOVdiLOMSlNNkFjqMmKrp4kzU7
RqPaBoD/nZuf+1zYBw1ciRUumYl2w5gFVyjNzkn+FsBPeE27XwXo9ZDtLAZ3zi4F
8Wp5nEaLYnALFB0teunKeQYXZ65lxPPCoyvBD7tZdPXJmkou5ejv8GG1FoaIHO4S
9ZF9qCY26uTFn0V074rJhSfQB4laVH4m5Rru20tfeDpmOnRR2cTAJHF/MgAsOuec
Klrij5H/vmvLb92KfUoEPwsWKsQ+8LSWCFMaWHscri7wD2Vh32wGTEkeQoVtOWYV
yB75SDOeutk8+r18HTWMJSN2cFxNbZe0U9KQt0okRuDpsDLlxXH35rp0paCZ6Nuo
UF0XvifHJyM4+FGjZZKLuic8Hr+8bMuG7IiHGc6MIb/QHAAcpMvb7R3mPuVIbBUA
aZbUVzvg5R0WJGvaiugcMOVrSixgL52rtihTkSVmqI5xHleBPow6K0AoO3T4ezf1
emCtrFlVCmxzhDYCIopPc5c4M8FNp7x8x1pOCFE9h/tXppzjsjz2h5Fdl39UrT9A
RsZNrcV2tKf8I6WlUrmaXEEIfxH5uj+ynG3HuHmzC3kWzmglVYEEjKdg0aPpBBTX
+vB4If3pfDyWP+NgZCE+91s4BWfm7pQKKCzkBkyfear0Rc5+vMB1P19RCZiY0M8c
vj2xXuOWqW0W9BkCDwPD1Q4a0mYoTpmgzbBaFpkaWjTSwCxQoUYDAueGvHB7wvxf
CWJ+2hXDN3YjdC+LgRE3eS1NRAijzyNez1Py86KzZeXIksANDJWuR0XpV9vf2rlA
ehFNOnPd6So7ThMA04z7h8BpezG3a4RSjgWTWc27F7clIyv4JvYE+1ViNCyC5T0z
1J8a4waAFQnmxb/MQO6TyielbJCkn4lhfErM5+Cp/lEUEW4R1o3Lg7fg+YnU2HCD
4R2V+Y+KG+TwpFUuBoiUXEEgxVzInzzeWebP6hf1ZpT6+AffTtqtu8KSmm230zX6
bXdDx02qa3RJ/4MBubwGMQXar3btTkwYKuVqv0yFB55Nl+D411mddeDETFrfuEDe
AghS0IK9s5JQKGvgT417OiimseGHBasbIH+5CuDUmf+n8+9JaYH/TpIF+eFxzFIU
WKScQ29R9oV8nSkPGB/1unPJZecS2aXI8wmJsvohd60ECYfqNr6T2Yvu/8CL8zxS
weYmbmh0PDtgknuCAlstbagWRhQdxn2TEyCsrretgx9gHxInShL/jA71I6er0C4Z
vZaCQ063fKpZ4cdH8342FR5m+tcVig+ZgJ8huLij4rP4Da038e8XYFhy7q5huA8A
WMas5c01XhvzMXi7ILXtOzctTBMh+SIGZ8ErTw7E9oWXF8HCyt/7Z2ZIgQ6cKvGJ
q44eHtOXnP+r4ucw23q3RUwa1GfvJ+ryrMioqCy8Js/kB+2xPb45jvbB+WzxDPAL
6DY5ubxNNlxiLwvSKuWc903OXXVsHZL14XlOAPwHWMhueecUddPXaGQnGI/l7noz
n0yp9RbsHsepZADBtULfzsYChyuqbMc5mAKX47O07RkVn6Ham+f8Us/9sm9w7hLF
NkOfgHKbnb48xXtUpDbnEPogI4IrzK3DVQdsnClHPEX41DjUv5LwlKgrRq033Ayb
nd8XmrGhEfwHFXsWi3roEaKXCOpS38tqRtDz9juFVbGeQm3ulfohtwUWAaRDkLBX
3phipXbMr8GQsw4PxxVYmzPziWcaotjFZmGNF8f6SJtsFieKlZBi2PC5RkLQBQjl
m9VndwWsC7JCKmfxh+CFaMTcpYLRE32ukjx6CRoOgLK4HPKurKXkkC4z48rpeetm
C90cvH2+Z5wf3kMnQhX/osyTNDVNN7G7c42/6uiZCQcJDBriYlzQBhouLNJD0N4F
IhLqkT48lY/iVxcwVKc/HlKaa61wB9jSFC7mMkBgTzu2HhykEcFVpvX1qyyFnwTw
1/5hc0/8D6dekL++sJO/3sN/AdvbFy8yMMmVPo5FBjt1eVbxIoUIuSyy7UBS/Yi0
+T0DXXGikLlcZZn9DLiFi9rbH6eJd0aUnby3b67B8KXxhiztWgIBmDdoucEOous5
ylJUUQ7erhkj7JUPhHPNSkIqID9dQJhEOLN+9gs2TCSH2oWVsfOmAsWLfvcg7Ugb
71Qvwt+JLNxaOJl4eFO0/QQ9r8DEWWRHhtfQ7m3ddHnRE5PKyWP239Ola/Vp0I+p
Qy2ViMT6rt5bMSY776imP/H6r1BewTyWRk/avRSZGpPImgUXTwuoBQuYZ+NoT3Hb
3y9RuVb+cUJJ3WChLH//9mvxD5I9oX5TNsB4iLv2kzhEm8OwnOXXnxgqwMc/uxZN
Ld2Ttz7hApxmqc7dZrz88n6w7okpm96HTptXdHoVV/to1aPPQ4zhY0YjEzC9khT1
IRoqGOGgfVwHiZpPOc5c5D+F5V3alsnbUb/QFYWHbI5pICn7Fj0QzH9pIXk3MCb6
iG1sFotlsUlCAp8QrpnMCA+LmMfBdG/xeHnjSVy+Z4IktL5FlbkEajcPZfca/ZCq
qACGP/1hcwZjoZZ0wrQKmAnSCvWCICdm6+AOXvIKwN1G7kHOsoqkTHkiZ2JMDGR+
awVFof+seoZrH8f/8IGx3gYsILljR59N986rKiTAkrO5ix1nelO1nyw3pfyHOXi5
odNBiQ/AeFGITSzj/EPZzBS4t8xHVfk5ZOG/D/avHCzHZaVtCNQHJAA5EExUn5Uq
J3XJvlCZFA6bEbGuOOAKQNxJjATJ6Xd79O1jzizSHaqj6xtHpIJBR2vBDYnLrsJS
5i5ktqKaL8BEfgD4SV14Cxvhf6WXVfDI+/DtxHgSIUQwVo0Y05I2bqVQxQ79dIUs
ylw19LJ+/ROO1zfNEEiFCtMo0CWqnpJ2s4cySl4Yp293tc12mxc+x1UHy4ta8VE+
K/cHdAnbRtxWs9sd8To7oqbT7ksD7lx76YKPQSs55ulp6bftDUdsvvaDdK5hx76H
cJ5GZVSet+uRfOAIg2Lm7goqf2kXjYmuZuCWTgx5n5czXKlV3gaai2o3Ao5qYjC/
XcCAqt6SfZrHIQr2JllbD3l0i9N4QXN7PNHFxrYEOEuIuwCnzGcYcabDSjX8OVen
yi4mClahWt/m0e4bCJIGVD2kwpVeoEi8ElSHARD6JbW5DO3AJLKFbqa+5+/ZaH31
Povkuk2i3zFJoHw6WtWuF4N8dlZc3nsR1WSqhBQrjsaW+PpVBuwzYSFeIdSIuw7X
dZwyS2Lo0LXlWo9a7EKlKOJkkqbk8DQ/PQZQ4v7qsoTSp07pqUGSa6ISQ8YdNfZh
f69GgpCktiAftX8td6xSxmm6hUzHJozj/54ZUoPYdbkjCE0U6vHS25Ug1I4aHmCd
HX9CkgQT9F7yHtCE0yw18xr9v2VejpuTP2uK1AQTHe1y5CPQD7gHM+KmtCzlyvOt
IKfyj0/NjQkVNpyfskDDpORygJIkbv2gBm1sIsOx1QWhDY5binjDj9y560ug/LK1
9WATM9gBKDP6op16HhQGgBDZYxQtnVc822HFSGoQj05zdZ+h23Ym7v2/MR4MDMu+
U4XaZo/YjFxcd+VEqLaQYRgGuAh+iLs/FNkeT/Kf2s6Ynxc9+57fXpUdiax6THXW
bSD0JoZ6uvyjbJRmtAHAB8X89UwCfw1Ram6oi4RhINqXERrUiYWkXbGz5FH/4h5T
qyR+8OXGujoSyCX6vUUAQ4u1Ghr2WkI9rrfBuH299pWp+eAWprtWOeXxkvi9B5Xs
D7uir9sZliTDe7wkpsNsjq2ZwmpenLf5tD+6u1aFsnqEJ6o0hpgBb+yMAwLlQw9N
KwWy9LqXPf3xyYfQXSF27s8U02ar1ztn6McHurSzxwp5ePXkYMOIA++Wk53hehXl
Gihc/43zkJWLQc20rMBCSiA8AmgfVj9vpY+c8dJDcS3ZqDnGWz6LNPNxB7HoK1UE
3GiBvTOs4D50joTQnFzg3GzQQwj3yKqvyNOIALTu8ZKZqsNl+HR9UTys/+9tS85p
bKhNpLYIsBsnIdf+Zz/jHQlFNheexn/NEDYDLxh5Gbuf4HjQ37FrdmbxjHaqUYyv
IS5sLVy9cOBqPenazvc1ucVrXHaOt2DXMQBT57SJ0ifCVXnHYX8K3/NsprK1WhYQ
1fqlQAphaZOxmMdWNsGKdfbSVLWR1HfjwcFAQ+HOPC89L31GQg7vBToERTcJHerH
ag5nhaWQerPNQGbdq4QKAESs0ozXrfCA8rhYfVy8eBQYoXYOHOwZiFkchENZS39s
afuy6oovU5f4bwDQVYfdkvJVaMcEAphRW++7o804ZJAN4XkLs70jnuvH3/tBWUcr
eb3r+xR9bAjHSmjj5EWeAbQU2VGXQt/T+8/XMvVV3jbMi/+O4bihbRzdZ2PHzvzz
6KVxBR8lcU9c+15MJk6uEPdd8qZEujjWKnwbZjX++N5Q5ImjcEM0a7aLLOVVafbb
KLDdJUaK4OPFs4N9JynhPc/1YnjttC9m3/IXYdt6IZ9Qv4RNCF5WmdJ+ine+hf3K
TRi4tLKCmRRMx0rlz9O/YwZ/O8ymQr9m6mDi6lOxVz5HyhodN9YVzW5V8W6XRMCI
QQTYg0nfV2knCR6Z7+4CJHc/UIFuvf0sy7oZ9tlmVWWXpKOeaMkqJa+MFxe555le
KG2GF42vLN/CvK1KPS+f/yl5l6GJqC6Wq/PllZ0Ba/E/K6oLjR4y4KQ56uCZw3+a
uFt+Ih7jCGmQYXcw4UWAAvWsXZxGTupUvpwVVl1ZMndyFewnEzOzfL/yQa5eaFbY
YeVY6J6Ubw5T33epXD7YNr6tW8yrzl2XmSPDsK7bUAHt7NtFlBb5viSBlyj3jXwD
6chhRNhAsxCZVsNgvxsHBQZEm+cTFnWiahHFds/JPs3FyEbNo02nr5oru/vueDIM
ZSdCCDfVVYTyE50SnVwGQhFCpRJ3sYJwI3m++/PkrVyk/oj9oEOth4MT7n6VC5KL
BwGVmTcGRaqfvVgCPxFmzeTTRNCoHPFd0pJVJ4AmezHRB/wH9K5KMn6R/ll6Rjo4
hrO6iMIo4vjcTFJNcfoz8nNMXJBarLSO430BNnV4TP6HPEnpwAcaYxb7etn76D/0
HVNvzai0FBs2De+eBLt4nXh/BjFNnB0pYDx08XeJrZyW78KXzwqKKVARHS3pVg9l
ITjlxHI+tK0hbI3JiuDr/FkHg0hK/qJaee6EVpSzLkXBp8woqBKcd14pFbKguvsL
buk7FUDz58cLHi7hwSTEPAS5H/N4tVR7zRY4QwWCf9V8L+4GU44FnhD6peNDBe89
geh8k6H4VYRnUlTI2gxiC2GoWs5d/sRUBRZOX2W+ewxtJ38HGE0xtWAh9Vu+5T3i
4NwdQlWrcXSL1LN+0FRbnei1dfp2L/qan0N/RzkkoHB2/F3acqm71IbXu+Ax1NkC
OTDf2nQ78EdgQdx0CAHc4v1TBYpQNGcTS7V+IR8piOzlAwyFkjzlhFax4FBbtQyN
jRHqGzXKKPeYSUF78wi0sYcFkQNBBOi4bRiPRrDjp8qBD0Hq83ukHGEbCO+0hh9I
/tBdeirKBGQwLqn7uJ4M0q/Jh1ZHElVM0vLVmJ5JZ1HLfzXxhWwtdeQnVncjdNGm
53kyZZ5u2CIsErOVy0XCvst7Jy4pQN7f7w/y2k6J719FmyPydw+5+DUZDAiDrW8d
iDh4JBpx6D6dbqBYbjFM9PG2t0oq49sC90BYpZIwIbJgDuJRkiCdfaGodJZbzIog
JnSA9/aMNnnLgckslkfy4yotXyPenFQuSpJPCGyRJQWJ8hQ8pNz76u4M1/ALarug
meuAodDKMfbdZwZhK/DqVlY/QGFarz03TiabLKw4lUXraAKfeBgbCE4WDnHOXosf
BonVwzn8YunncYKI3EomcOPomSI5pJCpIwXMnQ61nYBGJHheO4befSeq30XYp9p7
Pf3y4rRXNgIMKL+wL8HV3N3V5v1QmEkUpW+BsHcHtPKGsR+aoPQmNAP7cOdT7XZP
SjMRXlbpIwcdk0QQrK1y/1t1ch+Mjjbsi05QnS99QvveTWHd4cuisW0k58nmisLN
DN2T/oFxt3O/9CLaAfydAFgZweLbARoBR6mGz2elDfJ7FrofQuaKuCeBpSoanr2k
hncbLaZIUTelERAMX3K5GEbSr1OVPyvIgaIytuAPTezT/VSy2y5jbozRfPFekPSj
rpltgiFPdSlKcZtSkXRq1/2nmGYMuBNzEYcB2Wx7xSSitt3roOD/vPpwzrIFwzrq
i+tFCHZBUUCpeqY2DdlPD5Avr9SJP6HA8cE2ZdKQ2pOnv6NuX1hOO5omj0n+Tlmm
ZIUXK0wkw2KCqsl65k/6OuJzSKd2qfxuKJBK5HWlHHghI9Yu64lX82NTRB06B++T
DAQ8MX5P36GKXrt/gFhzhEoeg01gQk+dQxIcM8wj5fyN6esDPHDulkkOyy8U07yS
AL+6TOhRCHVwoKbDn/uyp6XHfJnlUNzVhNmLEz/Zz1d5Dytn037ASMJUzw4jdzK/
9R/jCuk7HtvXzx6SDh530wu6qJW9oqotCgtqJy4S05Jj9PlejSYgIoyaLHwyK5gR
YFapAAdoaejqeUXFnLS4aV6KpcMjyz1KWyHmIQMHrzuoopoLuP5t7xx7Bi3iBfTY
9g03jX3FFUkXtkYUUxZJdY+ttjsIdIac7Xpdq5WWtPhUCXNsfk5TL8RX1aTsA8a6
EQ/gWaxzByEJDyDCF3211TJ41rKMq8JdYEmdnhgJcP3flJRPtaG3zHWM44F28LgV
u26cC74JlhM+KaqBadxE45lgYlnkSNP5K+djJhlbiwKn/h58FU0TH9+X1BGkczfC
0X8SfljnjCHG7Ize63AxwTMQUx+COdcrClnBI/Nf5XtXDUS3JKdujxruiDnyRADe
iLnXlUDmUPVCaP06UwJ34jZCdqjEdVdyIfkFpLW7ld9/ZK/ffitupvmHZqItF5mh
x36VvLtiYqXbwlUi/DCktXxRQJT0FVKwqj4WuQDoVt8xbGeuDVYWP6tf+L75K62r
ZZWfXSdx7Q0vRfJyGsGpGGiFJ2ev0ankm/A6MYLe9XKUps1J5Ktncq6n9Y8/pXjN
FkJPKxsyTvCYE3Gjd1pHajLkBN78rqsynQFmTe+jqiTBKv3xsicbafafhPIuXAVh
fzxghKSnvv+aIP6+YLMJxX7Ro2UlybSc8M8qezJmg+tf0bFoI61P/KIq2qRAp4te
CZH2HsJMOpyCdAolDRhpuJ3G0jyYM0DpBpw4JRxXiFYDQYFnY5QtpYTrX+BgM1XH
xkHM+JXuNbi068RsMxUvC6h/bmJcAC88El2aOeo8iI3phQIl5TMIP/RjtqZz53Jo
X7NlJsCIFDClzB7k2Yh5rRHx2JaOVLwqxRSZr99LIDKCCmXWRcgQZ36RQRYRDAqb
ZG6Y4Jpm3OzRllHr0dgJsGSz3uEEmDVQvjChxLR946MEwmCzf+ZbCedOwCNrAzkw
dTuJcr/d3IKrkfBHRqWHVlSGnI6ZHDcYCvtHZQ/AMwD9k7JB60VlKpBXtty4gUSv
futhJif+JOnhYmbOitPv/rT6F/gml1AoC35cGg/iVubZffChJppPIQIKE+pXPGiw
b8IRn0ozWMWgokYm+FYuKswPllut/5E5d0gNB6TuPPGX18cgNQdzo4EmEcwYmaS2
QlIxEA9NndbjY3pshKnJXLJriaTwJX6o4JyzrqlHfTDBFMZOvTAafhT+dc/CjnzL
i7THjhQO+dZciaLP446kpCpW0s+RcVEfg9/ZpUaCQCgVBqVD58k9RMCah9ndnb0I
Yiy4ys3FKcLCraAnwOH/lfo10EmKMvt7hv73K5ynvam8Y3Y5s/M91VrdeiEbBw6b
pSqPK+FWv50189k7EqkN9cIjf26OccpSf4eROUZsomaUyFOgEC8KUpHUSJNmNVpy
TVJWpS0GeC1RQhwv+86wIe1Z0hIXRAaWfOuDtp72AKPimT2+xpohDekbTCoRBVPk
eQShvDTXag56QgqJX9ueSjsFd9dXB1jxTRuyZ02YNtV3T4XHqO5bWTucdYwmOS1U
7M4EgDiSoqksIXy6MddgGqgoEpByK8Dwi8mUh0y3ozmFB0L/OPD/pUF4X4OS5OyA
isAok+ugLMaMVSUeMAM0/0gZwMObm9z6OU1qaNCF2qqOAqM3yCZQ+gqdWrcLMA0o
yL9mxmhErvuTSYMwLbBJ//2sfYkZ15VOB34bNGdRbkmctPS+3N/9E/2AH4e5aiqt
Y41YVquYK74T5ihMFRlrBvOuMHQEF1nxWjuilb+R2Txm6/4S+ESUNyJGlIFcywfj
VpKWzUMYW2l+8DIB/SUGIwhZuAAFJL9c6rsGToRVbf3iD3X6sGKXXArtuJroN5sM
NWdtcROyC8zVP3IU7v90j5afG6FQxqJ8eSVL6HibEnPmgkWJcBKFiEw75daBmyP2
aCNLcLAf/6ZuZk6T5soJ0duFB9zKcVJh589pC3LqzVOtsgoW36yvNM+zsp64Ntuh
sLzyJOK3TM89cDpoJfTsOp6JJ20mc/6xSRSFQK31n/wg48cbGpvxOK7BzoaGkqSi
RFGnUyPzVdoGI6Li5gHJbnC8Ybuz7a3j6bSiC/mU/vNun/vx9Q9/p9UMgISyYZW7
BdtH8kRncSqUtEAB2yDJl9E9UoHFUaQXOuMvO0Q4jBYMuoXTYnAk01XcSxJco+k3
IvzcoMDL7nkZp7VlukZwW2V+ghi3z5d30UML9csL/EKus43K2AUGeqTS73ehq4CS
Hacs0DWr4vdOXbtdgelN/ROneEQxGNPtpXBZnhwXRrsDmmUl817iYjM03av3VDVL
xLVcSsZwaWsUbo6M4tg0dqLb20gMxXN0YHVPIo2GcNOMfNjgMAtqE6xgJIJizRfY
utjBXaVKn55JRjA1ja1VXq1FCnbYW02edxQUKggD6g9TEveIaXdr9c4+YqDPn62z
WxQoc75brXLUdoi4+DrD1CvzB/9YqQbqz+PlR6kMr3uLzo+8IqR/gz6jt5XBLWho
1MQ7J+ykQYjFGaMw6RFCgkR1ds1ZFsQO772kG2C+i6JBgALKA8iMBTyOQu8j07RF
lKnS8QJJQF3Dx90nRZzIK1Q84GuCS+pdgCz4JG9nQlHLFG5SLWd4B4f9BymXYFgs
JX0mP7z3cR8aE7wbM5URqgM2GW9io8Vm0owux5+YiZKpqX7plC+LM6xTujN7mmqE
vypGOAw5MNp472fTnzg1eRD7NZybfw3dEACJAyxp9geEUvC98bFkD5C1V0MXyHxZ
/1+Rbjxq+SlAw6PPSg33COQ67EiL6coFcIxrGY0CEWh1+l47PubmNFu/Db4VbMuL
Lb377nNb0I5cckrWS+5nZMHwqCPNQukgCKmpvJW/DUzP293I6ZQnFbpPTlU6ShcD
UQoTCyhPVxvmB4G58pbje9fsIymuPdutqoj8s0VcSay+Mhc3vhS5sv9OT8zLByo2
oIi9jJGtTsoyG1WAZRm2dDvrkNq/hBjQxvqpkmRW30Dx3KK6zBzySB1IIBLqRbIH
kSxGZ4YK3FP1jXmSb+t6F886LHbf4zWE89L1hbYC0maDyt2niuHUEkH+Kv1AXkiP
Nm9mT08Dd7HBuxwWCxJW51o1faCOa5t2SRszOdPqB7YhUgNRqM8UR5xS+vUtOovZ
VYPT8HZkrbhBHC95boXbrGdhpMZeQgOldxFD3qFDjNl0KNhBmCt1vCpjfLrNOo/X
627dhBggp/YRtkGDWmjXIIWFYhvdg6OM3Z9svfx0EwWvgcgGvEHkh7uwAs7JGm2r
OiZ0N9PsFx7UxUyggFT1ZY6pUeH+FrvND65gdiIoKLnbiTs9I837T4BsOiWsl/0f
Ag7pocyeuL0mt571+qqpz+aRIAHORdqpOhxPCocpJirj3Nh7avK5fJJuHpl4ZN7Z
Z2V0Z7eaCdekKRYLyjytlxna+FTjTDeOS0M6t5S1IvYkhrtVKh9/Ezgh9Jq0fSMX
JOBx1ekII+amBFCr132urgg0HueYghRgQHeJhqg1CnSKax26u38YmJ+eK2TtYe3w
mZi+hn+eyvcDpy45Td2uBbdlS+UYqrdq7ou5vcpAfqN9CD8asDHoRI2SrB2QndVf
vXS6YFgqOIen1G1m8hKL+xMecB4tUlfh8QnJ8AOqE985evVT3YZebVlZ9faJu+Ni
96Eis6+gAjE/D5QixBNDib6ayM6mGGMel7yJp1EF4HX8+/83xJ0jfl83MRfGq9Kg
XKTzORaRPjKgwOPm92hfOwF5WL6OnPB4Hr66gdD0Zq7VGILEcgTcl+9kkmHmGLhm
OppQHVLPwM2/kWF9V1ihMb5xUgvLLYlc9JQFBleEFV4ZM1Rj2UiUBwhWiHrnrA68
LZtujPrAyvDr1wXjSuh9CBFrYp1TcAMLrbR9wRuT+SeDwy0AANWa9daT2nfnn2/a
D5lH1syQWN+YqYDUqz06OJ0+fKtwh7lR2ExN7J6GeSxUs8kSHfduCUYIsLQtRlZ9
20J3V/K6CAgLTkur37T4EX3u/gp3Y/S+47M7SpaLo9ZXBO28AN3q9G4gd9DqtfQp
eWRNhcITE0H51wu9bG9UVNR2Gv+ImIFpTCwY/vxaoqRmTX4P2Lm4k0N7kIbJUkFP
G5YfKQx3LWHPjCkdH6OS2HUS4QOgC4E/thpjaBi3QGEcEyQLAyvTrhMN9PltUJH7
8aGuuHQ0PM5zItKZz4JJHrzAy7wClsJpVCt11ImNp02ck5UBF51F2pmT+z3433ji
p2aRqQhPgAOjjjsrrqIVUHOYBwDcEiukQgA58xK1PnQ81rSAjxeQu2L8qcOXHW33
IY2Zpn6X/L1OcmwPY1mH4Utof5zgl5NkNuOHCAxIlsHql2Qi8S+GoSoxrUGScbcE
5Cs4d9fYziPbultGac4WQ5HobgOXBv8pJlXvW6SlAfHp5mtSNsG4fNWGsgm7xqSI
BAhswFs7UY8nUpAyNznMQidQgNBaF5webxel5Le3plcMXn+eMtNIvXzUOJ+IVcwW
3F1dwFydl5Duie8er91jK90RXYMbOiox/n8LDllDewekvNYzO35ClB++qReSHn6Z
6zfasMftV+oTn79f2j6o4lqtiZnt4DDuCQV4n+tTaF+2HjG39QHpQJVNhdi55O5M
YsEAn5T6fsAH+GGeK41Q2UqNj+2UzOCEUDzeFCqHBmQZ878ylB+kkyZtrlnw35OE
UH//XLhqs/FOaQac0R10+2SRArixdW3DLuk7CKdck7bPbyzyR5/0xmCf7ju9NaTv
3e9ZDXmiiMf8uHr0TQ+QXCAO5J42sgnfOI9c07+ndiXNUwZx4bpOw1xw+to76fFv
gsH6elrfgZXTOVkr+QnvK788ShwkTqxK9kvNbJ2dQv3VYSDK7vz39nqG6x4Z5wG7
g598L+emWCWpR+TJi5nfE/aG3DvKzQYom8eElmikXhMXQXnMJ1KUOe0cbcmB2PbV
ZIhKY5ygw3RxZVAdSrPE8dJTWqErrOnBk86NyS9uZc+xc0jonb1bQIj1jgS0bVPw
MaCznka34d9cRXy+adpDghK2+bz36hJYvHkO3oPqC4cpIAMaD5t9r0R6BblCwZFD
e9Q4YyfgaBzMpJUdFwjmcLyM/xQem5WRBBadj8Ajeyz8jqy91BICHitmVsrncNUD
svNHVRocnp2UuhzRrXC6uB4oZQLh7TbSIHbKKFh+h7mRoLb79xBHCN/6PqVlycCI
L3GTY49MwCiIujsNY/JlnT16V57bATvjAtahpuVOXsHg4T2G1k9oXgCd//1NLykW
0eUCj+jdxD8W4CHWWHYvCfnckAcDp/0Xu2r3ueXsiGR1LV4wm53m2++qhoRpIQG4
dAXB+xWvvD18ae+1EIa5DlzTV8h6AuuEPSxYYbU3yl58eB+kWGPWiHklIsQZZZEG
rmp6MPcpSVYAhurZ4d0b/bujqbyhUwpIyoUVI9Gk8bczmKIds2JYe5XAlsC8xpuz
1qWLoXV974S7VwwprBqcSb215X+hmw5V5J0BdDBz5FQ/H8U0T++uR/Tkvda6sU24
WGiwac+ClQTN8edDUXWJ4A7rkQwfS+KZuHaDvVGmdwH7rIBd1qakSpgy4NRCTbCU
L+D4w5rvr5lbDDCEAWwywvSmEFwdlufjlTTtUWtRzahkSt44p7eZAVcxcHXV/XVL
kjttz3evznfVDNEYAdU+Vsog/K6X62l/w9dQbmJ5sf/Dxhn1z/aW7rmrKYfEsY0A
QmsHh0bWoSgX4c/MlyIn0NUakKkOd//wczdtoGaYWfx+S0v2oWImj/r2ndz2RLrk
rXCSOUK85og4/AIhLPNMnCYZt6dX378VT1+7/lbgWJz4hLZi/eX2/6gtImlZeiS3
Pe5eqmAFchmOBllgx+P+cTkL2OBtSeMvIib80wrdixjSWmEeZVgWhAo0p3P+UJnz
DpH2AN8POpIJ4uinOr5zhBQsEQkMvpM5/i2AjOFkmBecnsCWmx87YqB13ZSVSGN/
t341akXjgSUcW5cTYjK3oUt32XbgbKjKV7Z50Xa0+1L8ZYw329ID6QT5difAq+Fw
5ku69Af8yDwYNfIqa8R6y7Am6tYzfwUsN5La/revWGceRHdnMBd7ITWOOXghmCN8
GxI7/2LEnqPQIZ+PDMt4pdo78ObIMHm5ILjl6olyc07eT10kSCXD5pqc6ZLwzXFy
x1v6NUbNO47gI2fYvKnYSTOKevKj14oFBrxuLmHz6z1v+ovGs6YkGo1sbbMzGYbt
YAkc0aUlzMoboixtMcuQERe6taMSTLZ6V59vC5FHp7Z4idRFyD/1KTJXch3rOnvl
sKefo+KH32se1KHsj6OIgu/iu/j2oHhxUqQrvno9BZGjyJD7rGgHI4Zr0ECN6O7r
UHFSEL5sSad/TWe4bOHahlw+bdc7AN9KhGsY4eyGGMayEZday0mDR43Xgxr5/osi
JbOVZOlRVPGkOp3yDOawsY7b14zj3hJLRdugT2ww/HY4vc+BLqHDhsSA/egRv8Ay
T6zYpaK6T7GL7/ABZs2cFCMsOjLt9Umoh2fpAWt68XPS4WYXF8U95VBrAQ3KrM6Z
XgTwmtJe7LcSItM0EbrP+9OEo53QySzf09HCvIeNYQRiQITQYz8kMltb+KR4i74r
ETgCVoHBLrkqrPgJTDYeOWgM3UpKPwVPzhoBSnAPC55UKSM0yxigr+hr5Uh5yExg
ac0hXGKR3f8rrR2Sz2QTNr5B0fRPtOB/TPzX6MS6Oppg09ynJOD7/5g+y2LvaU78
i1JxpM/7j8URJIpGpqcIruUNJWoAsVCilQzH9YVDsQOxVfH1D4taAB6c+qdkmrzY
nbno9OANKSABe6UGFl+tLKBxlEL+kn/iwlF/MzcrjC/VECuSypmJT8BZcGHik3yN
b9rBKHphMxqkYoc4Wl4n7vAOmq0pVWltsXHWJxVkGG+awK2k2Ff2cQaLwcr6aG4b
o9M6y97ZubY54iTfdsAWPG6Tr/mterYzGs6iNrdshUlydVHRUl9kTPfSKwl0tDc0
8/KREDxtwDNDsB+gX2PWkwJiDVI8y8JY2e5nnlrWoIRpNjcddjiKlis4yDhrTf8R
/ju0w1ty1UcnFgO9hR4cIAegDD+n8wrUJXMmMi86WrZIm3dyY5PltqogPHKtf7wE
JXJ6j7J0vN+4EatDVKPuuhLU9+OVxJi/ifQPk4w5M+aPVQUBuLFTQeEa/9ZaJRH9
6qnAeGKgyFogsXq7EV35alc3vMCDImXV0Iv0L1EH3DWz6Pd/KigVs34DBO8LhSLl
2VsnE7DZ3+b5yQqHCrOFFMr3nZ9nAJ2KiaHBQa7DFTKJ5kZZfGTYH8EK+rqzcJWe
//zG03qJGuWk7m+wppcmFEj/vT4rLjDFB0TPkVht4HzXeFe6A2iusQxiUuDMKKml
FItFeWlda7TNWtuP+qHrNIkb2KqPMo6Em3oE6QPrMZO1vipWhr3TncP7b6IhuSIo
RlrRmuM/rjtmxetLrstaAl6smP+QV4w1bel/QQ27WPhopfJyzbGaPK9RhQSPP7lz
3R1yF9JwFMhERJb44x+40qJCh0ejmE2NYJr2IPcsn42+cFG/qQYkaNJF/IONl1uU
9XG63wxGGUggSU5Gu4lxDSOjKhgD/NvxCiTTxf0rM4GXL4M/lKp5fR40sNMGjt5Z
N7z10XoQCpU17wov14BOvwR66a+594kWpBbmIDNSIa/oTVY+hDuQ/KenrMpDv0r2
DCxgQt0THoZJZP8X3edCG4qUnhvQ6FLZkn8qOTQalx0r14ZAd/3G6sYtMn4v0yYL
HQp7Z8qFBvuS9ghiaxjsN9eRTYknk1I4ywizK0YNK/b3yIYSwX3yHNzhrUABJ5LM
iqEMgcomVjP22aXjmxaF8n9/ZSt1gPP6q+b5tbim6mobHNWVealz3+kzYJ8a2ftl
zUVaaCbBGJgVE3Q2HErPuP5+FjGP1k+y8Jx68hoInrMcLPg/7RxzdTo/SjmO8p+F
5ah4kgjFKM8YWcrrKTKyo/XRMEby6mny+4A1KKTjj6a5R91gGY/FI7+fLkj3Vxt+
IygOvR/5xSB/8SJigTd6+esHvw0x07Br23/CmsSMftogf5GL9rpzwTvFp6UZfkra
mOBAxQhi1jflCYsdsFvYT8LnNYUg8MjQMUVtrrF95AK5XZJgjJui/Imb/6th1yCp
K1hdapz7PhHEm0LVG4okYgn01/UNkXsD+VijFLCIGOBeQ2Y5DtRcoqBkHoLbiVKV
7ps2GRjPuwCM8ut25SMtMe3MJIC01HLO6/9ewSp8ilBkdt9mvsAPZSRIw/rmOJ6x
A7rV9dtJgCZ7JQ81b/qqMrvtx//wvBjbbLdB0R3tof31iKF4J6If6XVJ9MjS5Wjd
AJtI28bpO1GZPhICEk9vpXRiCNcPw+IafYUY5KW8DZQG9UqAA1LMd/nq/JcAh4eX
G4XUu96z7zmJeACk00p1eHR2uDmY7BOW4hHZfusplRHHLRCWtrf/6CNurc5csp19
QtN3V/tEWqEGxdWPXjya4yJdJDFYi+6iSFo0OXV5N7ye27KT99kzU/6eQqI4KWTv
prhGQThi3USPKMjrVRxJX3w+hliFmKnN1Q99h6pqPF6hTNhiaO2Bh6RXyDhwmrt5
WwTdA0cb1qCpz+JYRUL5IKE+XmtN2lmT99xnGAs6Qel2TA/j/Q8lx6rn2lEkInZI
Cbhiscv4pNGA1gK4HwcFW69bfK8XuAzqV8CxKVcWjQ9+a6Fcq9mVzeN3HXJxDwT+
YuHplPRmy7cG+LImQfu13XHQBA215UvAD63RdA1Mq05fyJzOrl7JS+1cWTb8r/bV
vC1kMXSVQfm4pptjwzqtT3IUYV5u9tOe5AcwK5LpRN8TzW3E0K+NsyZ42K/T4K1n
3GnzhH80iGFykP1OEUyYNwfUth2jfW0fh3HJ9se6jOttoeWNm8CUu7zdGvOeVKHy
VogsrigWgqM3HhLVHRz5xcyt2hPq5AIpa1lcLsqzi1xeimysA/KikB08eRnI7hcZ
rjIUxMTRakrlqKl4fNFaFFSk5RFC8E6wMR0iMYNzH3f5CeR/ymotR+G7z7/6SLaT
Sd/Odga1jD8Yy5oRjdkpp345AbP6f5McghVfiQyQgkXThR1mpMmcIxq7aNElko0C
q5YxNSMcuc5vooMCZ/wOxLL8+TjjpPuDyFFPpP1KI+7R5WHHann8QGFUp/NtUWby
bh5XIlxjw0SpBb/QrB7534x3I0LRSBGC+CISq90tc34gfZhIM890MjSwiVLJRH0d
JnF8GXo4DOkMMZeBwFQ8kt/VAr+Z3qpZmaK5iFC2gu+K7oZpfwUG3PDB9x8fzpNs
MbavD6rJH4JW8xb2UsXtP5rDf2CSslLQtSEAn5kjOQrlyn9rlzrXeOJ5o+FNMoZ+
a9vHFk4hAT++SAGWQtO9qkS4UGqCqJDw3qO+Vl9oxc9jNiW9/VF34IsSNHNL+2W1
isalUUnxNoXi1TiYdxVxCbS01knomtY+K/7piBotEodaA86Lh4TnftstbCfRChik
sCUYVt9vkL1XRe4R3Ywq4UaLKpvWze9jkxKSLEc1WCezW7xPjztMGOaiHxIangWj
mWrzMh7UgTtX2T4vbni1j/seIKXrD9xkPuOZ6NF4v/vQ1N7vHUqsnrGPd+BT7rUt
zxrqj+bQB3MbJE4wmyDoK2jfkkbi035r7fF4CQORyWFA3HU4WSm6gP0JrEdbBNQD
CwBJv1lXK3suZF2pTt8qkJRLkm3k5aqXDspfH+O/K6G2df/QNek8q0If3vPFzYSl
o/9j4MS9dQ/f7LSFTQkyKWtWcRiV91wFGpYhdA/k7z4Gj/iqkSNcrj+qsKZZw/hs
PicMLtu8aUrapjDe4o8jDrlqqtc+kR8JO7zSroqnUr9eRdx+L4P2RhHnflq54Ndz
XnPuwpHGtKovATTIcNDXUtKXHqH30DH9PCXu4ZTMS9eyR5th6fz3qtMT/KbBpBaN
QTJ45jXBs9jGJBlEqGmUNIG4HuXqGCD97yR1QrfJUkMYJ9jUFtJMY+M0+TFH2icw
TAQSBPHpfhx1Ce/o9ekBpb5qPy9icAc44x2+UtyZoeZVHkGoikWdTToLP94qzTlZ
awLqjhsQagyHw7wQF8LM/8YjEOwMTa5YuvHdpIGICj5pIS+s0eVFkjzF4NncjzdO
yo5KsAeMrG5ZHEaS9SpW163Dt+6p0j6xtEB6BRlK8zgFaq0mlkNmDqDAgAeItvG+
6LRz5aVSkFlcRuvoHZjBxpI//Rap9O5ErE/1kjgnE/Ii+3o2jpfvFeyhqt31dLof
iTDcOHE+32UEeO011C1bmxlvPBWfoY+gH266E+ZfbCdDOchJxG2vzLwT9allWcFb
gDWuOy9EOFUUNBbZINNivu1jtDM4IEN+n6tg+98NlBKiaJRXu07Ta9idQrYFtHno
sDKbeCvQBLyyivLk+ZEV0OZ42LZJIYxDlA1K0Slrsh3UOXTMo2tWoVCFX3b3IJqQ
jlnGssL2gQ6/5qZ9mcY/JepseLeGJds8x622zzpJemyV1PSODrdqLYJq1BoilJrV
9iSulTe2a3B1/p/P70XbyVZToZ+Dm+6CAWU6LC0CfnkqiA1dwA4q6611DYrfEdox
jP2s2p4VaoCJstZWM0U4b1tT4fyXQ+QY3PJeDOAqbAH1mKAhUlwoY8qGFvgy6INI
ulK6Bj+9F+b6w4t8+6ZAGYcnHptvZ2B9r2fIQKab4Dz3cS7LmWjOkODOt8saCTln
ObyEkj5ZyBLO4yqu/eg5QqsdHpgbQtzrUZZgqyoCwvWZMYXE2wfyHPU9r5+GMT1U
4YRDF0jjDFsID9jP1hyhDPnRWktuw55skgPPWMqVgIgHdqiC+J745HrgmEI/eAL3
NGCohcru3+Fr+9K0pWlV1rMEyYjKq6FXgWLaH1MP6QpgabBNn0dCUvuyaksB6deq
lg8VC8Ydibg75SJpGJl6KXQYCKzKvY0Sn8mTG0NgGxQfCjjVaFLZvXyL46O+05Vb
83d6k7dry1SpNK90dZ20/3uX6/YAUL2+1/ydxc+SkYa77TYSrnnr52GihSCP7M3G
KHCrU3hGJZ+kd2H+NmmSLmwVKMIWxS/DMNj+jDnMCG2bZAFS6PkvqVvFOzQLf/TY
MzFF56zHcXxAAw6H/bz7lH1wcQYZ3d88Qr0kNTJ8pX09gvd9LmYFcXwRnIDeVt+6
lud3vdPra4CuuwVbKE+chBAorFzGtscZSP9l2r2j1qKuaiUbfp8LENeUjiY0GdgF
3mB4aioepDc9J9ctFbu8K9UlUElecqtCyOSc4HA12PBtVhv8OKLUemQiPMYQ4NWR
0QC492C7/LpTatO9bydG2+G78wMLO6bUBx292QUx4k4CB/mmqbzxlyFC2MO6+jSX
TFDxqsEyeGXRgQUxakg7kL+gF5gZNtxPYIUir+Qo4DRWfSrXHZWgzQldAwtm0Xhe
Kn6zV6ptgB7t+10cQE1P0e94NIqCNoD40xafmUJSUL/DsdleqktCDV2HiEsqOzSq
P5O/TLp6rRVZicOqhpo1UNqezi4573q09fymbyDFHdiN8sTUg0Y1jV6yn7T+BALl
TmZL9sZ+GAJkldX+Dhznl3FRSRBy0nCdx+SIzuY6XoSVBdhlkrnvuFjiatmX+cLm
zvXFskmVtWtmuXOMH0e+LApa5Fu6pctGDDGL9EOASeBKP6LNR6N9UFeOL/s8Gaxf
XHP8yfSKHr0NG76KAQn/WzQcMb3tkhvNjuSsRoYMGNVHiirOEHqZX/hg375GYJMv
6gJ2ni5TvqD1srcszLjOUBKRVdVPxU7JNOpoKOfLFdKdPSTvVM31RAhuE9nYlujJ
/0PrLNY8wYfDuBfTrtWLQPUNYwLmltPSVzZ0FVSNn8LlLtD2lK3GRUNvUaMCkFzu
NG1JRgk77wcxxBE5IgQDL0dQ73mh1qbB/oh8n5aEF0rfTwml6PAI980gtObI45ma
jhNXnBFfMI9UGrATQtAuCiWZa5sFdKb9+0lqKkJ1DvinCSk6NHyIg2MG9ZuHRarA
r6Vkk6ETzEUNzFrIEZoTdYqwKdRNqAX3y/Jd6RA9ZpqCZ8DvkzfLEPjZah7iuSZj
kXHRlOZ1z8zLaxEKaQ0mt5M6b+M2NwvM5O+IXsFX0bvywyfjzpG15zgGlEvlXdNs
F1hA5+dQl/yrZoGphs/h9qKTY57BlKiZYPCvIQ9ydTCz05T4Ygjw6MEBrwyvuaON
0QWoltDqqTOfpvwhwxjs5DZNZze8hGB/8G/6wrciJ+ga+Q7ZWwzblLIUL88zGKXk
KmeET/HeWLj8/wMdxfsV53YIhHLxz8O1ga5ciDkyj7QldUYXgKwRrCi3IR6Bquhg
k3UgQbHmhy510QKuB77QcRYHPZhQO7bcMavTieDOzbphuVgsXyzgTmsdKjffkAnE
0eogZqS21+DXdAFG/xkVWpUSJuJb9evLco2WCAsG99badXHhUoFfHaPBnm/9VVZV
kzj+QTX+ErY0FNqzWOzvt0sdLf28xG8ImLfQTp790YC1fajhOQgzvm44jFDZGLAs
pIXZnfbTU2j6ef/ct0ED+cfq5OduG/6u6lq7mhlHx0Ktg42fMTplEVZzMFsw2OvG
TFI+XLT4QL1fvT9gkvvfs6LG4iyeQAqHCvXEjuI2VqAv9Hw/LDCRMle8Ka8lPP3z
e4CPYSqVHK+jATUySgEXIWRqxpjbdD362xG/ia63aWSjmndbj5N6lySdUbASZZ3M
ThWL2fugdFYJiw7TRrnrDtKSBNMvPKzNB91gcVpPOoqxA6AxQiDqD1yPCILSjZs9
0NxnfbGiOWf8JPhXohUGJg0FrnIP1153Mt2Qb8OSfjvz5C4Y2I1mc9MiHU84h9cM
Fp7SLMsC/42nhNjnEXtblXIZU8qg3hgUE38fS24BC46Meg30ieiHTnFqbuWEsn+5
jGyoAwu8Zc+5wjsdcYlMg1ZJuglKVADAO+YvnG9dW5CtzjtG2iPk+Y1ERWqB0l3w
3tdy5grvFDMqOevZwLMF9vDVZQXzSIJvZd0N/YHbaE+khrGnmJ6ZqKPl0fcmP0Qq
oDjdmmcJT/47QM8Dvk3b42UedASM97/f+qcQ+iBxR6cQNr51Duh9hDUQAGy5CuUY
im3dQPKAVRGvFqNTQJfcERpIadFX6/0bRFIZSwIGBcr1YquoDxx2Av2e98W2bGCH
PSrkBZP3eQjh1HxSZZ20JS+KpYT0c81lchOUBdzfZnMOTM2OLM224ZowrFBWMoSL
h+OobNHlytLHzqYJaIn8mEJ+lWWJKp8AMLqa9s8hR8755uCFnA4JDknwM5crD/b0
W/gQdyCUMvd1cQTAGebZsbyvDkO3Ca5UrUJoBIeZEESNpxAg6WdfRZoDnoKg8Y7T
VMW2ypGGF7WRVxIuzJSHUHCBEbvC3RG+dHJMaRy6zdsyOuX+HfkoUeo4+U+eZItf
wYbJyuZod1r0ZniFDaARxAto0w+P/PuLq3GDQBYcdKNDjMwoXNRMqX9kun2EOIy0
lftrhkbqPrYe01fxGUABGiDUtjloL9Rlj97TO912HW59vhW875wXaSvwTOXQhNSV
TXWW0YmpMVGwFAFnoVHF9sK4n8vBLgu9Ab5Z6A0BBFKiOmlBrXUGun5N7sFoCdB5
ljbZSBsuu1ozcvc4ZA1kfLaebYWXXfe5D8dxOBySpv+z9FWq4L1tdRKg1TX+8HFu
v3Oemhsb0ajQDvzB/KdowsdJCeUItpEoUbkF3AumvtocQ52rdEREmxxyMo5MuM9P
zND746p02ldqdAu1LhnAtc3uO0uMF1F/lCXFHq6WpqQtn2gcwV9j7MIPyxqV/ODY
UMSkwvPTgxvWaF72/n84jlOOjMTEe4JUBMV35Il5C4Pa/l3r58bqA/jqyIpsmrAO
1I8YWzjvx4MGr9oST6zg3ADxt9sKm7Wn33JgMCiXsAECifLiZ5niE29s1VJjsFoO
0VzxaXmfozGPt0+SFD6e0N1Qy0tN+qTp0w+qtpmsmbm4RfS9+5rxCiqz5NxXv5BF
dOkV/Dusn7Rwa4/SwuLCcmFzAG1R+RcsraIjZdFlQGJBDM/0Ah/yudjyLvnleiXk
vTZfCZ9h4+aYyyA00qe8/vDc/Or0l4veIWUdUosVWiVFPq1a/EnFhGUgSApOve4c
YnU6y/jAExcksdVNoScCj+yKhZLBLK0RgkVa8TGlsNBBLMEZIClpOr2qpQO4EWIc
dUmhhjsG9uBr5/eL2PsOMnYuDZROdJpUKw95PQrQUszT4l4EUNHTMQXa0AZ4fLHh
EbT82qrQApp57xTTCHivNbw3OzjCrctCF2rP/iiXQnzhtT6AmGQh0sjV/9cVArUV
SXLj4tA55GwHXORN8EWdRpMR/ta0rOHca+hgtdzcuCzUx+zdUAkwE4C4Hwt/6WEi
vdka/BBdzYnD9SjfNOafc/ZoXluTw7xFhoVlB7uwzkC5DZ5Xf7+Qa6jT2B53Qkks
KVeuJ+TXY2ummYM4ukAe6Jeyxg3CyKNNhjqfIeLgvu7kDNdATmytUK4hRI+2OcnC
c0QGdXPRiAKroMVeaqts5+xASfWnJqPTogvUoq+AMJMwPtkr5OBAfz7r9AIh14d+
I1CdJHuRkkJH086+82H2zRiuiyXiQge2iJYiFfBgWDYU8c6NDwZ6kzfgvnfcSmOz
AbPSDub9SX3A3zo/KWGOdLaBxwECYA9zh2r0uBrvqUiE3tS1Iy1j1+mqpGH4n5+5
ta3qHOcR7jJPQ0yuBmPV19pN3MtJ3epkSUWqI8/6zD7nPXlMP5ZsQUroiygVXBLm
DoHPpE3FJPuOTkpgEloahkl+XEH1N2q5mbnCtXzyS2XqAjFCye7bzm8I64Y1ltLw
Z9zxLrcDQeoJePFXUjOldzIj/UjFBabE1T3nVm1pXwBSapVmV6KUdXolL4+GQSUg
xLxxJrKoVg4+3nvzE3ZL3ndATZC3+07UZCuMUS0S9uYTSXxn1GofEnSYXpWOwtx4
3ku19JlFXzQsAIB7h8AtDjeCVU80qh1JynakrgxjLD6mjbBTqD4SHuCQwGk+10vN
sHOIHmX7xfeCU572dcQ8plRPrsmZxdih9zI7iCDvHMcqeTmEYKdr8YtknmgsVeS/
aBH/mxz1X9BbQhnO6ipsZRwfd7Lc2VBRT5NFI0qiaCdeSeNmGx/IpsL6xntgbVXw
5d39HnGI4iwIJktgpoF5nAccu6zjmAJD/uzlZbF/8cXDdUr4Ib6y1cvgbA12rzhQ
haXS/9MwaYZOYEs8tRFBvUl4NWViucsZD0uRcrbM+chDiTY3pa4/HaClrA/JN0fy
4+OYK+sQjPm6fD4PNUcVG2wKPhLgwyVzNeDfFoTtLNa4o66jqjXBK/tc2JksJbaH
pUpqX4mZ8PgvPgq877mZ4mDp5tJ0IFwX6tjF9jhcx/eyDnqX4OirG6sGYD4LAV1j
bcaaUYst6+weiGzpkAWxoShjAxnD8KcEic77qPqw34KavlJkESqhv5pm5B+mfjJK
DXAXzd83bTFgWyzMyAY0fLlICNQr0H2McyXIZLQHhhB4CrcbrVgDj5hcjjEDP8ry
zWJReStjSwy1EaLXkHt71qt8X6ieD+X4SKcLNNnP7Xi5siPwbKVyWa4ErY569lot
SEozJjMhgdXrALvnUBaCALjTgJn7lsE23iyMaADvD5mmFVuz7dCTPdisgCc5YILp
zC3GtC7r+rtH+Vj1Ybg8ny1e1tMVA4LVN1FwYsk95kJ7UkYU4LU1Vt4jb9j5aqHq
fS/OD9OpautVDy0OrOm/8niudK65SVbHSC3418mdq+AW2gsVPZZZx2vR//FIqGFg
ThOriS2F0xwDq54K2xUIjsb1wZ2r1/gxEmigzLMFo8CpfNFae+/aRtTwH3HFNAEz
pWuHIT37OGrmRakfloSQ169I+ZsEyYcosZSbsPQdUGb8g8UxF69uvrkPlvPKMElF
WXwOC10M2GL9MYNh4qMVPlV6iK2VpTpMDtZGMtLlX4XiCZjQB2WlBnWhCxmEZAhV
ia76dzIfJcMqHt6tBR8+rdY02t7HduGrLwpa7oYUMrrtgZZxzbnBLkuIhPaF0O3o
PeNXUZX+7Cr+KIHVC8wcw3VFxowMWQwh2TXl6IfzdkY6AuA0OrYhKUJSQIPHxM+v
Psz+TGqGwSBm/hZrQFsNalVgOKyKSqNluZBRjJHZjvYYmEjlFFSX9IsUT8tmWujj
RUjStg/0IFrRAelVqTXssjJkQaEWQLwZRiSH0fdtIxneJ1bB+U2t8jwrZEvgjvPz
IVt96222jzb3WEV4kDefXJtK06/jIA62PPz/guZ5si1OkOB1wG94+DPjiQJ5mdi3
DqU848ISqeOjp2uACbdktuJYCToy5eIkXj4jpNI76FCNogETd+DIanz4ZpBfjb2v
QURfJOMRWV4gKRk8I9WHJqGFUfJMhY8v0cBjKt08Knu0ZiURgxbBo1n0hvV+XYwY
Lb3wFt99+jJ6HTap68EiUjhf3nbO2VNo5xDsAe6EoRgGktforMYpuJaC+7O3cPQH
QarerjA6O7L2QTiMPjGAhxjmgtGPeWlpaW+0s5PlMd9b+r+FF8bI7wUW9FTokDKV
yjBcXlLq2SLlNQXREubK3yaXengEp5Iw21UmhBISEOatUxFeE/ZBA+SSRVbiEj6+
cclHni4VrW2QKNEYL4/ooNhmXMvfrtiY8nn7k6aUZOWjO6MxiL8U+ZmSnEbN6QUU
hcNx1rcyWlOa63EhzqT6MsrfZLg9EqLImsRYqm/3u0lsLZzdukxmhH0EvkjR+50l
XsKLjudKzAK45zM6L6de8a27Q5BdiGaGjBdL3wyCMPkvuwuxWtA4swARyF9zC5w8
heHGV9Vc/bjLBfs7gBKZA4naAT5Gl6q2FbCcdM7AfDJbKdqJhacgBCWv+H8g/S/2
RPAfkUd347RaB6/luIc+HOvLpgX6fRlV2vb6PLqZ6wBzjy9kUCcFIINGkewWuCys
jGix8TfZREsmjtRCpbfCfSArIx1j4Z5Fy5+zVZ2A+SISwQg5lZBz4kV45Ifx/MJn
XzrKZ54wu5Igm5Z+PxcHH11w7dt18ImHRTcBjz2EFQfE/xrQ0BPLNqc8iCpB9CMZ
cgNce1PjI47RLh7EJayuV/LWzXP0f2tK53MCehEa0RTYJyEmc1DPfNVLQDGTDH0T
EpEcnZEjFPpenC1M3qTfcHyRt4zw8dxRCJ3VuXPr0ZZS8sNFcRhrEOafk1geIcUa
MmuOUNFr02sAOrqaP+VioxDuCQnSTxoTCHpoPYD3TJBSxdVmoKfiTrLVuwxKTEMc
lm7F21Ia8OD6MLD5+eg9NBNYbK4L0/ZFdxW2jfhGP1Z4bTqqZQYdOzwd0fILEgbH
60rm3gVzVbwk46QjiXUF7bcGBp1AjxLPavvgaaOidwksJvR8W39OJy+VE2ENIT9g
32KDdBTFqjJJDYN+cPtrUCIvFKadBA3zthOyCAs1nmbWL121sawQktMJQ8TtSFXn
2MnzX3/JL9rf9dbvRiwGAX1/yG4myRxOlLCYOx1vJbZ3KCI10tgr3ajSjUz0XbJ6
S3Zm1tY0sFvPBcWcDsUd9H9OwXjmXcr5h1V7pKKhRcEF7WEUPWNx5uHmeBdaDo1K
luBkq+Hj5Z1OH1QoOHMCzRdv7y8+4MYSwqoaRSGyc2LM1IEzsEywfCs+4xXSgsgj
bYdDi42MAfCLi86L5y8PtahCPOx6s1bcK6qqElMoqJzfxcN95meRYeRQvCMJrTdH
26FkXjL0qHC8RBXPy1FXNBngvz3gE3QLwUY8JGPiYen2aqQvXxBjx7V2+yCsrayw
eY2i6uMwRybtEn+UMc5iXCL/WuiQbYX04VlgpNNbTxQA5E9SyWqEeGxeUJ/1McwS
wMKseKHJnGjEDzVIN06OdsE93AZiT31wEG+QaYjkSWh3y6j7wzjISMeo5MsqopiN
/HnhFTbJ3hoRCfdXJVvX0lX9n5IXadbTYPdMvVzep1DlJcZj5vG6ZNHujCHD2iZu
xJdclRCZOq6S0BYh7zEMPzP8eFNYAUJ0yAYyhY9UTv2ZNq2TsE8AFxrRjS19/IEj
Apc4SHNKy8hdyTyC5n611JSbnkbvHFpek4QS5cwyBD+t/7KnSWB5cHLASm3+g1gr
7vG/AQl20bVUC7gLh9lL9rMHDhQB0AkIf0J5I2pLcKUL20rkRMHhFH0ZSyAx/9gg
IK+wiQJPVHK9QVfjHsHs+rc7VIEwzRsPuIDms51CyAMkvyrfZmzDOI/EzL30qtyQ
h5h4M2wFicslBViA8skE7MTywIpxX5LiDf78fj7JjuTUpqBoVqDrKAssp1FjKw4a
Vy7ST4rOzsrObYVC9UdKkJw5RMb4GQWoEO7heMUhux5Gf+XVrkF3SbklvLbv19E1
y2KNKXqLb5DDZiaCJrkPFkAcagcdQduvCLjZUwcYxUaSL7ddnVFJgeVXnBlqjIqI
4sbzmeWAz+S4w2K8FN2Z6nPM2Y6cpflRjIZHBr+EgROK30Qf3Emc4rISOgElQXb9
5aM19BRUx1flVOPOf6aKWOp68NedGHtGXW0HHYR281l8jp7kx5T4otdhp9wzcwU4
KXN4hqyTJDXeXEgklVlhatb5/JtTiQfm3v8SZn0+C0E2yQY0d4TzBYSyJKgU+WER
TH0b2L7/F5QjKIXJ2zlAuAkASoIfJSSmylqBuo0ZvARsY/tqmP5m5wdK/+ah31xS
filAnbCy66Mbaq22WwLkRAvh12Xu9Y0tcXFpganSYrkjZNemsxnuvjjdmgXT3gtZ
EyHKyw8g9j5wpLrLC/dHtfgC/zoWJ9qWRawq11EDssEb3E3grRF+sxJ/EYcsgf95
lLFiZbIXf0iBOb8EjiAzEnrJdty70QMIep2QX5E0sO2Doj556DyCDBrgqvsGAA5W
d/MxUUw4+c209iEJNaAXpNTqp6uwuG+KOXPZEMLuk1h8cPgIeqsTLceVNp0PgB1y
i4J08eao27Rv8eHaYknRfxBLECP4TjnUbmUU/Jvq/lIBB9WSH8Q/DvcUx63C6n/t
qa1eJWANiI3ZTQwQObxiac3PDLTrFmHzu073FWh1M4ndY2bmoPxiQvJvOLOuvp7h
rebZpQ/3dxGL7RsLAd7youQGXqE2ktxseClvhrKlLdoqOlhMdqTnX/DZyd7A/yxC
258BxTjUlRY2N7WWjILgss5c0KvC7aHesED5PL051PQYMZ9i436DFDeIN9CeyBu1
WSSMcB7dSiqif292w+UPhFOQUMIbgkpZzpehQ4ra7nUNcV/JA0u3ZFPrLOhOR2zB
/niI+Gia7qcmPj9zC9WbbWD4lKE60/WUbMWj/AS7/q2XiXUr6/OykMTEM9rhs70R
00XxWlzctDJ3Q27akiE6YJXfQyVXwVvV+OnCgl3U6PHVxJ/4n7OPlXtH4cvbz+dH
FjdxCnu5iAxbeb+aN7Oi7c4UtbBBdjQeJ3dAJRZuLUx/tUcYqu0Dq8l2woCioBSK
Zwn9GfWvdUG1b2SIznh5sc75Krk/kaR4G+FprrwVozCou/OeRsT9iq+hXZt2CG46
/1Ew2FtHBdrY7N7ayT//whcexatUKZcBJEEXdCj+hJ/GcVJnH6pH5WYlkmTlEbrD
cQXYqANhFO9WT1BAG+vGekqBBTUqqtlAbKa3ib7CuSNxz6rHr9eIY9lTW1bHdf8W
DT+TRNaqKG4wKgwN0PIXpHYv3orrDmFBng24Hh6mhpPYo90VO1Hjo252z2gHENoY
mTQGUZe1L+tr3TmG1vc/F9FpHZA5fqMlaM+ZsFKUc0oMTk8ahdh6pNWYywNYtncZ
N5bZv5QH+jrkO2UczHjOBpNk5KfuIGXFj7qZM8PLXLlFGlapP+iCGigjsJNQy/tP
iLM9HY0RZFCNyJUKO0paXL2lDIc9eJgFDXr1Q7HtE0G7g6iUXNFNIRTKiNUBuGRm
1LR+b2GeGlXzctFTXDD49/k4C4hCSWf57cZpXqmFUK6m/TF5BJ9Eg7RJCp66EU9A
htDmDOmVDgVU1fQFUiAL5nABbNzZktU5udDX/l6ejp4iIfwJTx2c6WvcflJIu4Yc
/xf/GJ/mxJUn5m1iF8ee2+39y3iY211Jq+PYBUnM+8ibo4ZAMEMl/Y7Kk0eJ340o
Ij3YgAdDwcGoNIfQjRLIrsihIHEdVBQ5hJBf2AcV7XWCJTQm1h334IADrkZYSw6E
ALaoIMAdZzrpR12vWbcAJkhH6GCL+nShxF7lxUAyFncxNQfL1P1KmuXK3kYsfMh8
GX6eRk1OEKN1JkwKeW8evNAIUmzuQpJxYTTr+ciD3XqrFAV9nPtFg+yuGdd3/qY5
xWqKYku8rN8PcOG4lVYuZD9ZMK6XQnlgZBjsMlpYSzcgMZ7HMl1B6G2Rz+fRrohF
oLzCG3rR8UFThz+zaSSkH5z2TJQtmyoU1UwFehSC1PwD+ncgCsCSi8mKpvPxPPYA
rUKnjoRHeAU5tM78N6/2ZuX92tp8BQ/3/cs7H6S1S47Kt3ypq6nsjK5pioCoPLkk
M/LxWRSPTH+jR8xZ1mBDy1vyVAR1p80HNfcaRatRlgzHWYvqgX93+Rd9N/ADFFkZ
CcLqm4wTGr7A0YC4rM4NBp8F/KxJ1En5QtpWbIaBBlw60yzzASxgRwcR17j7E4vy
Gmo1acHZjuGoq5Hvh7nOiRay3dH+vIwP4XYTfYNu+f7a5vsYuPMiVhACw5L5MFsz
slF/EnV5v71ODoaWn118l5fBhsr44Q3nAO6iStSm3Fhr53hK1EHP6zphkDZ/gbQK
UrkG+5XXkih1/URdr2EbgmoirhZ2yoHVOkZDpB4J/dSsgIVeX3WkiyQz3IuP4fKL
iXqTg3ZShnRjfjgNopa7Gf6jl1fPAhb4j9NrHSPnFFquXoB0PQoyjcmm5qgyxEg2
BiyylcUt1fF9Td8u9J5R4D4oIKZyQdZpsSp1SnJS87rUuXJ8d4mTxGf/fnYPkYQE
cEzBUtQlygMakSYig/s5uC2HAH2mUF+9imXG8aH/Sfe2RX63MzSwPB1Wk9YeLR3t
rVFGSwfpfGSHj0Z6Ay46HCQMg1hobJ+DypPJFXwNAo+c6RtzidodlvA9vFajGsuz
S7U7poCf60Lwednag1bos8XynU4oraiQQo4jIYqcB2vTfQwliTwaNZe9HKrPRVRG
M9E8ARURIWL2K1ZfprDPE+Ic1ap9EFv3nV0O9kfpRvSSovqAU1EkGL7bhwXdbSWK
y7l3/3AA7ZsN17SgnIYU8pA1fP/UfBWoeFBpKp6IGa0Mc+mmtrcq9jJjLlAI+N8j
TZTv82dkPEDWH2cRF4+crcjYF2hGmzZwilO7+ynycGdHaetyvM9Fr4XlT1sjI3ed
FMNtTGp/KL4Hih3Xpfc9N1Zz9oj/CcUnVft3X4D74jRHAKZnvVZ95DNO7Cx0tCeK
RjQewYNTzzAsT+/gs0FGtFfdgNrm5espPSd5qObvHNTRM6k/CIk8l0Pi++r192HU
VTqpnOCSpAKyNoxaIesphPXF1uMQy34P1UuAkjbY4bhsmNy+IMq16rz1RcZj9MCg
C3ZLHSdXwtydILB7i87gfSbGkjPQk8y4M/CV1OdRCs0aSGd2JrKAlSB1e3Bl2HLZ
PonU6jp48uzE8U6Bx7PK/wsOhcaJDWzEEIDsDabpn/z/rtH4S6KImUgD2xaS67Ir
A6kWA0jPMSB2uyrz2KVxxTcabmgZxz9h2AaHZKvlhJSSvyLuG7S7ZHculGApXW9r
BuzDN1yhG3pwBZCkpx5a301Yc7qvcBcaJWNux6kFch+PJhNjULD9VyhfZMUjA4iC
lplfN7yGxFfbTkFhEQIKFASZpC9wVcc3kJZPfpzmJSy/ahUPYrZ8r0aMx3ViP37f
/MNAYmgTmrw0jNo5u8vlt/wEQQMIXrCFRYp+WbiOWakcTy7XLxHfTIwLQt1FDHk9
U7DEwNc3oNjDxwbD5FRp9jctFwMMi4jKsH0ZaqlqHgJoJlAJTKX9JykGSL827hIV
UFD8c0YAYUlc7ze3EyRYNmtpmulyUVlw61F3QZJUeywSs+f3vxygrbRds8Gyqw9a
ewRIm3XkJ6HVOf/apWFsH3wErAliBPuDyx6+s3i9MSwZX9x0swmimU5MQxTRuTeF
nsYcofS9eeOcDEbgOxQ2cm8nUH6AmaYq49enwzAyQb6OpjuvVqjhwVItD4e791gI
2a67+gX9Vx2CYHFBwQgVdPEA0v9AaAl+UgWjW+2V8q5BeutPtjSQEvQUjFw/JDSx
XdEjNaqilIo/4a7/zJFsghwA/CP7ssO4YrlsZrKLQRJsfOl3LxBvdCHm9jcGGcRO
rBm+yXl93R57nunZXABCLsh2o1jtWqrGcP5fmRXqv48H5ZuG4r76oMgALKC6KpR5
AQ/rvCDL4TjOTPbVNkbbiUmvjRCzZMXhdXTcPdyvbhBxqG+DVF4y97amDLQgTzlD
j0soLd/v1BXXPQ0tGyJ7KsYtDMIjdnsO1nlA/aGgUOmomb7b2UbcROShfZs0Rblt
P6DUfYm5oG6KxdY2bYSbW5bWG47suuZ5MbuVlqHfpEjy1ZwJWubcVSrA60quTOjc
dAaeR2TfRIx3wop220zoC1l1ZTExB0e3aJCqLAdM0Al7YsEBJE67NQ9LG1p51rkv
cQu35gg9jT1r4orSfxtoQJFI6Cs4tmeOYy1RgRxObcE5hGSBWP1MXQB4g+TloIgB
jawejq4lpy+IB+KCrpe8pRwanC8CnfFgHbtFn66xOqQxk0dP+7e401wgscobmvq0
qeSY3AlGXAa6fhz77c5qREZtTmDYk23kNk6g9P1ALXhbip80GWn3HZSrvt58/frS
iBxMkfiFE2jsrTeT0KibN8Q1pb5PEAw9VbVrvXwSfL1uT3G3jifdyX84LGrdSKmc
jMS/BaU+Tm69OvHZu/NXawTn2kikc4bzL073wgLjBnelso9HIl35a4ilK0YndxfL
Wm/O/PEwK3oorsAxPypNIdw66pSbs1aOzEBipRC1iM+wEQnCz45GCWWKL4NKQU+H
ndi5YGcoDwd0Md4ZAnAYrvqVNvMstW+QuI0WLOBBtvQs5lTzBM/Ri/j8NscP5ODQ
08OZXEZAZ0AHHg6Ha1i5rfD5rtaveIIjfcadRKz1iwUs/hK3qsL6mWGdhNAVzONg
so/fkU3jMeTtyVJ6xR6AVss156Uz2zA5ESmZAgtpbg1CdycLhevoL/M0wHDuEyBk
tRQN49vNai6EXXRhpOIBvmhe/CjzS4KQ59B31zGsL0UdLb56Cr7r2w3dqCes4pPu
9CaDvwZT7kQlI3m083MykVsQmkoiHsG0HmYOKL8Ri4MSt1ns6g8bEHG3QUKLODq3
XwZ7IQcbocW+9X1VoUCF6kqiHqbRs2x9l+qTtBBQyfTl3jc7BNoifqryVFrVJTjS
dpjVDKd6tpjLQiOsWMtM48T1ehjNVRotayYJv+XKqgLMXERTXgfoGnFk/+huzqfp
oGWYeWdzkyQIRmAdSMMzrMd/J7AJ7vybagrcnz0myj/gCXXbAi0BjxD1StiofaGN
CotLe2jf/WDstSGqZ+DDXg1anpc6aFPiizAS1K/DsOnqvq+1GH4GzIN3qHiOn5j5
ffhDjrGP6ORlU99sPjD99FcCx94qiQEaQFT9lYhb8NER21AwoYGVuIvydjrJDddM
iC9ZV7oRFLDmmrVTwst9zPbQjO2Tu+YcJflb7h3ZAg0aCwjIKg3lwaG59gdZGhLR
ork3mZlZhCxaFmU0VdcwxlmktS7jrDGI+HRp+d5hWE2tWaAtqaH3s9PozUsaQ5pR
RMt5uvmk2LPePrBrbS0rpgGQLjfTo/La5cAT1hUATt+AZCWwIpBc1m9LrutJmDPw
sSlochKaiwW/jv1KejXX2XNXLNxRqZedAu5NALKnmvPmiMEiBsWEEpDyNdM5ji51
5MhjqJrjtVkV0jDNzx5zfAhzZU4IaRNC4OtGee6O0yXMmlKwW9wJzeRY17t4Djtd
uTwhVWopNJdVHQaCw6pYZ7kuZ8a9Up296KTcGbO6Bf4VjK4+d03V801MSWePngGC
pOIbgyKKVv7tsEBvsxHFPDDVpdmUbvyYSQ45Jfz52bNI62Cyh9Jrfzr9x2XBPppH
CwBH5p++JXpk8cxynCoCUGu5x9FEGkBYycTQke9HLKVczcqBRo/pD14UlIpYWAp1
P/nC/M+XgQeKE20n56rtAV4+qqzGjKduCdGuonwBIM8ohBEyUKsbK7obF2DSV+rf
k8EOc1tCIz4xEBfpz3dS13M8EoZdf7tMTKv8j0qCbRm0qWU6f9tpgRhtKEuFVrJR
9N1ZkMFbmDbK01Vi0CRxx1aeoabSqQCwm0m69o9ufOF5aPQQVsZK/1Jha/eaQE1W
SKD6SiHQnPngtlqrae4Zh1oJuiLhYhOPXBTFc0hMfukW1YbVOgxi4X95ahKHAq3Z
DCCyoS+R/FpM+PZ4Qw+HtEXVbkh6h7/ma4jaKjDdcvB3i+0Z5VxKPLgc5WJ80nRU
GnlkmY/0l5D+CNMBD8hL2ambv86mTByArAgTT3N18iF33r5hC4RPiFGF7F41h+9u
716nZtnxODzgQm3w2NlQeSkvoRKEnF9jpxMZ5PYFeE4rAGBCPyOIRJNx7g4oK3vJ
dasZm1pjgHkVJvKOE+HpokAXjlFqQZWg4W7Sn0IM4xdiPu9M054Rtxb1qiR0V6+o
KAjIxBu1CcpPr+2oYbpfZnEGRY/ofGAqkkKqajtOzu0Bt2Bj3g1uHJiA+fH1skQl
5xd5hriC9JKyn2Gq1zzsUf0NxlH9dxlQR28c9AgQ9Ag8gyfMnxetEbZulfIecPzr
b8g6jzXk4ZU3U3ICAWgB0nly9gzHG3mEF8FwaOsHg53R3Nud/IFZVQG3TZhyexfq
5HTS3WucrnFNWlbJXp3SqYtzl+970CE9jKEW2sLRfjJtyj8xI1doF4nmPi/j9PAX
0hkp4QbV4l5tOcoLm24Ci+3AlGE2XgEHtuLphAyhlx5OhnQSD5X1wX++NUUtM/nk
r9W1UIRA6q87EDaRNWxlOOqnB2uU/PS9/Ce8Mt1AdcQC8mOq8TPW4MIS0mZZQUm2
CWAkb92wiSpJHoP0sxudhWhwR7LE681QezvCTvBGVunC35aQhsne0CZC7usBBg4b
omtiEXLQUcKo9Y8FduQNnob1+blcoVm7I8MH3/D2/YdbVlhTavIuOQIu6i92y7Y5
JXocpTu2b9e6riK7wIIG5LcGuCGZNjPWjSq+8y9uaZf5gYkTKSglDiU+lue083dw
uYhLYqgPX5dtAU/fyla1fCSQZM4AXgZ14tggLsqZsK8AKkIYZhiCuQ/ksRcxEIUg
PEt7SP//CA8D3pS9rPTe87OjTLRuGCVw59a4fXuKI+fl5mr7mTrsz1utjbI8FciZ
a4SYd3h/YdJwktHl88I7CVRTUw5dqyuJlZtz03ZjxFhx5t56sbyYlmeDY7FPQbRd
E+JYwNWKwqLo/jrgpcGf7TcQJAiWhvAQnAUZMMIQ/FISp4eu2WxSJvDFpVc+JjBZ
8E/gamab2cH/8/SVY1M6o5tqoGCn6cjOL4QlGzbVtWAwzH5ZHPmb3RT57BqIOMa3
bPZ1dx3F+QrAPxxVfTtI964QdcV4BaQFkFNs/mWXNcb56Yg2j65OHd0jVBt5WQH/
BpHqbtjQtHdZZfo1OG7Bi4f1g11MASjI4pa/IK+FCEUlX4GHWnX+scEntbztAQwh
8BwP6UhlfVASW0uFrXocqvayny1DrCZXPlZA6BEIv+NqQp5rgKUQuwBXtfXcT8Bt
/KF0751hV7f7gkR2IsE3CJW0BP4QCrwOrMX5lLAjkIdby60+N/AgNMdn5eMcnMld
9b62KeO+dOLNaZKevv2v8Pr6P4j3W268iTK55w0s5pZOpcM4b3NKIEorGTR00lBA
hTkNJJ5LfU1TcrXQvAMUUCeujBsHijSSKSvxmCKlBErfq3Hhp4/tqndVCTf7QYQr
qYXiyDB1CPizvN+6/pjSOLDcI0ZmvrFOj8QvrbNBnmDKmE4bJQHUW+No65aw/Y7W
QbXXNfSHBlF7/InlEo3l0/HGedpq6O2/G1ucvKvqJI57S9KFCkYNYypfzg3l5FE2
8JGnKuiGLmugEHkILmibBPMY5WhiOxdiNHAsC05NFD+Q99kXQ8DdXGoEyBWqWXJi
G7bkHDTTt3sc8u2CMj9JJ8IG5R/OCQaueSS0KVcDXEXxiWUowZgBTEQrK9CO7FHr
ks6wlENjyDHUpNO2gB1ZFeetdWTgjwlOOXiRI3rmimRHCQMif5R5sW25n64IOo8G
dTeXEUE8TWTvRWL/15atqpe5gMx0KygAryeR1xH5RH1UBcZPgFv4E/y6z9l3ckxR
PcRE4pdMAWWziSvTkX708UBvgkp5mYoBJz2A+bMqluQXq8J4gFwH9SHbwXhrf6mL
u+HZ+OvZeq4eG6oQwQwj6O7T0Su+tUP9yS80j9CKUQF2l4bKiW2pU/RAy0dq3KL/
ERBHV6iB10WApEz5QUAt1nuS0Jj27Il+ziNqyaR4d6fueAaEfBZYytUZ57QFW4Y7
X2YRaqIsNaxYsDXB3Suz5zG7QD+QfSdviPuo5BTkG1rqMOJ4Km+PWRLG2yYeV5L5
domHMeJJBSFNGkYXvO1RTdQqaRbeUxVfXI8X9ArpANS8dMtNF7MPbQAA3UUopst3
oTIFOVxJ4zKrgvsBNqdNbp7FwflJcvyv8Wu4y6vdok4JDQiZQ7PR72hxx2nmGHP7
jzNS8I5n3j2kEJNSengxgyy6jbAlWSkQTSrh8TFtNzianOJcYbcJeRsp5jFwb47B
b6MJ5uiE0BHNVDdT3qcyM6FyDft3hcWrdte+bP8PzuTtbSVvXfYBl+re8jRnS5Ms
d9+QuA3fMH8SkTVybLdcOoJujaSlstl0ZNopoWKHfr2Y35DNRWKLhDfHrNJco4zx
2+jpAPEDeK1OfVgR1zffdyi33fsq++BUsSaFbJyw7dhSOjOAQs4VrC/TBMr0hAXA
OG0MqswOcsFg38uFixll/evEtnXEMA44pOBuZdojyz1I0oFxwJlqrufq1wl4R5dW
v+hg4bpuYXDuIq/wzKblddzjbAZ28dPCz3aDbkaPNWwKZ+OhFvHKsUZPJ7Ozpwlw
yWlX1CVi1pgj1Ej6o5/C3V/r6u0LwXEhAbai1F1rLFhx8Gcz8ILjKnwzsHjkXdmw
YA6LIA7mRUmY0ZVhOBKqxqzvN4jMy9DmvR1rXuPgS0wrRY4Png7yqRbyoY6TKcEV
KF530vLAV3Ns8IKcfL+KZhNlAqoN0zi4GPe37NqXoNGKS9EORA55bUGT3BMkCZip
Ne7JDyLNt1DQ3vl/AOeLlpZUXHj8qstzuYVjvMQUKw683BADi14mtZHwjaPElltF
B7yr9Hu4JF2NAkp2SrYBAlAVZvdI5orOkBZxNVR7BQT/8ymzv2KKs+xCozMLAntO
5PIKmucH/ffQifk6Rjd6BwzEnwdxx7o0JdXkaFDL081g7AH4bE8M/1ZHS+mWZsDv
vhuLe0lAaVgp2Ku3ZRH2Q6doaiUvffB0DSQG1/CrhD9BanOs2Ks+ymsQyNfMIklu
4nAVd8AYzk55KxkwIVtZPKhheJ7YK9n+m6Yu0q9FArWO7MwBLLJMYactGmf70PbD
xHnz3ZrONLLP+KPa+CRnOM3Wq5Jml6HFRaiPg5uM3MQ/rmRVUgn9a6E0sGwbMQ6r
Q6FfTweeFD1G3PhtK7TAML+pVD459vB14kE7inISlG0NGnECj2s0M3u5jcbgX5KQ
tzYf7zb2pJ3Vpb+QF6zRDIjgWSC8cW20rEAdXVeWDGG9iRwSEjKeas5dxW7k4DcN
SonMWkPZYZB/FJ6SfKm8FHIDtw7Kx9GnHD6Va7zvx9QM9aw/+eyt/ktjLCY1c6uI
VMF1CJYlPOuFYkH30NOkcffwOKtNMl1QDWQRy2f2nRDkRUeff0TE3nKm1c+Byeuu
tNNAwSoLFUycN3vLMP7CiNXrOziWHiwa1Rv9X54Xkkp5tPVmwk4KKKEt/CCPNOVY
mBWat3I+veolULd5AqBaHKnbF9FK6dcpmgXdVsLPQhXuXEbZWI5UDgUp9gGMwOeA
m0ENJQTAD0VgvdqR24O2BF0IJXvRDahQGXCgQpT+3+zZaNO8/gOok0Iovm1NooDe
p2Rj/E4ISlq8U5Y0DkYuEJv7eHK+BHwrSRVIqyx2tDUKUxguwurnLaLhrGwdZfcb
6I4vTj1ch3QtoopUJfZCyJCU41+O9rFwGXfzwj+QDUZ1QwZoS1U88M3/A/LPlZRN
faS4/Ex7RK+41QyjJ1BGESrWTozT9MdhOPgJPF5eWhtTsML7D1KHmnnYh/eTWTEk
UuW67b8SMSDnCvTiQJCKHEz/EvBQZuqVpjDOEJMKzAhSA02s4gYYXjcganGQLg0T
xgXd5RL+SP2dMVP3uvCIpKC4i4d2TLjkfZwPkPMjF+qQb19HNtNM7Oj5VOtWXa4X
8rtG6nXmGAUNrcBe7wSVk+wKvm/7OPx+LiXFX/XuUbyzNr34ALMRTVPbKrQjLRdF
WUOz+2WoNQDjbG4URVQgbcWDKaK9FKy3yatfKqhJvzxyJoK+hgb4jnmpOxs20HCs
Ytxff4vR5v6ZhO3FzrLRDX3GFrLJTAxaDFk9u0d4OQOU765r73d7RC20T7abuCKy
9V6QQoRE05wx3GeWKgXF0JDVRanbCXiot4kRqUcZH5VjJOlCwWQmP34OSJXhFYjr
7JUJH858b2kcFacQzp79N2kQ+m2yNfZofpGONlYzkqkOIwuyHs8kkXgTkoqIDzy3
IQf3ANCkDtzMv/oh9NNpNpDJYWvTUXRJx2RdI0rgMMgpc2wLbRGLWvwvHN/kLOUC
WzYbojDqQUe9DzpibMZragXr0St38FGID5z12KRL5wWcW0N2Y1SvJ6+Et7oWlsE9
T6jN9vxT/NVHjGkb+4W7JkM9BKrdc2fz06tF56ggk8OJECVDaXIVDwVunOnW/v7I
b4HStvCiiUmuX0IiBvYRnR9XZZbpAa6a2Y8SEBr75uApEmG6u9yEzRCZ9V6RUkWZ
QcWJgIuyNmXww84JUqF1vCzJ5V7iTo5oaGxMmcKyHmeBu5fQIwucn9F5pcqtqgYh
HUT+Q7BVFTuu2tiIfcY3PiFNkt5BAET9ZiRm8IQXz/YZ/7EOWfO/cA/SeF6mSxMi
TLssAj/TxvyQo1Bk1Un62rj/P4ysu+3PVK+ujSKeMVT2G1/2IIG10vKH7t5QaMJw
AE/q5PjuIXwhvVMvbK5/9K1bIh/G242OUx76i2V5Ot3NUQ6GcHylftjTwLnJOGcv
IQHumJjgqMz1dbzg4RDQCHDohmACEGlmOc+1Cjds09CaJLsZN9ZM3eThwmHYm8wN
ihqhwfOggK6ntarKvl7dH56k+ScTxWbuXTdz0lM9NrQTDUG3yeIJ52ogUFWntQdp
iaJzF7EM9bibKRhclQzPpVh6vgcBd7vL3CBd+EFq7DIBLceBeHb4XO718D2qNv05
q7DiMwvNCIVbi+l2LiybBj8iLgS7JhICbd+1sNXOsmFUZHct2PLvidtbJTJOp3OZ
Yx+xXwCoDbAA1GtDlF3XyMn+e/MfAtX3p+jsCg2b4AzJYDccDjMCCbvIIHqJwjkX
8/TOP3GVWCFyQ8q6xUwuOA47rhtZI76Y3eow5moZQWt0FJkUpimODbQ/twuBMc9G
8igNuJsGw5T6OIflhMKEydb6CGn98rYbz2noenHR61oIU18YdGO1v8RyuYhQwMZF
GbO3jYQ3zWxpE4pXLRaYJ2kMSJuMkaKpwRn10fdE5j2RGbLroQ01bBesKw0gF/fx
e6JhEj763RCtxdMUmoHx2ph63dtW1F1met8eo5bAS5WnABSjktofxxp2h2sAqN3F
LJV9BfeX8RL/DEYOVLhmtVKo83veeTAJLHCBZw7j1g6tgqef3GMpXWK1NO2JE9eT
aJQ4GdTdaU0b2B0xkCOHYFy2qYo4mdJvhI/uVOHnwGjDrf8A6zWokCZYzWI8NUIX
kLWWhROl0mv4V279dHSrgtrlomn21AqQNCk2Ye8WxuOCH+P7um5SduugjbEYU5e4
tbfM+OVviGMGlpsEgCtYQWcWi2S0jur3hUohyaTjbrhtzVncy5X2OADOCwOogLti
nm5wEacbs4ynulbh4ZyTUNjgpyO2duY3zwCBz43PPKc+MtBTelZcSQSxtw1hRR3B
yOki14koHpWBdFKO6xch1QCcTy5dQsx3o790wamRPrEgH41vH+Uev9cAak/D3EBG
+I0ppemoEixhW8vA1inhNSBAApLNvirMpzr97I0DUA9dH7c7H25o19VuIvugnKx/
zSLmQmS/5/N1bj5caC+FCuyJ0arrLSMBGClfl+YoKTJUbVGX+4zuSAWjv5uP6yIw
HzeiMagqdgX0/P2Rnj3NJnnLd40Tmhj0b8lEbDHSRkHlemStvK093d12PT0byUd1
9ONxMwxRj5klDzGchgVDXXGShScVghmVRPZ/jOLOKefWwo3fjQTd7M2lw4f8bqz+
ObtkGRlkros4q9X1l0vs/S/l9bdgQvoeDmQAyKAK3TnvXqNo5KiEbDi8zlE7rZGp
Dq2XPGvP0k7MCE/nIV3oNL/+yCJzpU0XHCEKhhlPQVtF7IKBnOGP6Q13sEI64D1K
NIwJprkRcNSBiLS6DjqaHSdYnARhxlzlbpSxy5PG8fJKlYOGFXGzF1pMW4Sem80B
80Q7WPMsdM0xThZDljzOEBuZQ5sHnkoGyzEOhpJN9ZpftaR1pjCM4EyJOFoGPlgP
fR9IwPVaWPXnxuuOakgmAvIS4lzxeBl6x4aChB1vZ7jB7W1PYa8xydSlB+geDQaX
wH8LsDts42T61tPlOg5djJLf+KqcqLb+KBQuEscMcVTE8ElLuf5AScQUkubsJXRx
M2FHuwxuvQVzf8/rR1MQMuYVRaM/PgYhRUE63kqDrtXlgS0pj1ORkogAk5yM/SSE
GQCZmlZChiel3kkVxEZcXgZ40nrhbr7epfMYKPoM2q65pQIjiYAUT5GdUpcqpY7V
rK8iGB+1E7OOg0CYnrwR0xq+ZandwLAd721OKSBySMWLXKIwJlJ36F65nh35SUQQ
JEKNiFn+C+u2ejRKUJxM/Oat+LAnZXSoRKnIXKh+KVyrOs1/hnw6tsmQ6OoWBOrC
8EWhzOVhMtZ4zmlfrQBFipQ7n237vsb+hM9hjefkqU8s1zZ5HMTazGl73EFBFX3R
tYHJW9ewSjzeQK6REVumZH3mr+ZLrw7jiyebM++UmJOtWuscHLuAJ0gBtF41V+jt
/xTO1GHvQHX5IVEYUy9LgKMYWe49l9/qp7G0z3ZbFTt5jug8OcTeTG/5Tcjcn3Fk
DNoi4ljr6N9o5QacZDGkJ2d/G4Z8oMycM2+v/Ql9fUqj1Z20h+95xn/g6WRIbN+L
FHbnDbBV7beBD9ayU4cy8O3E/IM5Az539+tcxu19fK+8VJvGavEXQaKEmPQaa8OF
mn4JUYD8TQQClBIvb2HVzLjV7ujkKw1mUxB1B7dRrCtF4dHnnbTiEU9+TaFcXRgK
DqironURxNQxB0y3iypHNB3/wi8jtlF049QJ4QIDSgVxBZkDHQCHkl9m2C6UW6W/
NZiu6klveQQprvk5mj35ttENIWeHZU6/C9FcL8/hNsqmkgQn+d0e+dkhqZK8NaDV
oN7Q0SLhPnX3qgRYlUnZ/YBJwKXci0Fj9jICMo3CnYxv79ubxuQSNh+OMMtydapM
lrogRbMTdPAVR8wMPRomhm+8WzmDcp6rtgTGz4XRd7YK2zLZThOgJrp7q4N5hbZB
MV4wKdKytRVlARhKAM8oHF+4Aa5InVUGdqPO3hYkTOp2U8qqDnI8Bieqt2LRL0Fv
zBbSL7BYwXHh+1CEUlC1nVUQMuB5jz4X2Ql4gyBk3kD9dj7YQSk/5XSNohstl9/c
xDquNufGpSys3MpGDjz1BQLAwxuImDDYz15QGA0frM+/ZoaG7+R0Gw5GOQPLOG7K
7FVw8Qn8MhlzfK6nxpPLJy/9EZ9dJRsXnyNQmMb/X8P5yGU2p9MRifpngISqNMoO
LB83lPTHH/zTRhspkbqvVa6oDHiHtbfXobETWepDkfSmlxTY6heBjm6u0sFMADjA
jocN4cdrqnDBG9cTpSn69hzaF/jWVx3c1jPvrFA/LAlr+Owe1gKfbgVv0SyPn/nW
zKfqm+XruQH0fM/NxKEPn4CZ21UFFeHJpTaiXMNx6Nzv/3Q2Ra2J+qOrVdM3h75r
swLlKatzD+cYRSxu5uXPXxDb4jNdIIeuu4Kv6jVggFgIp3qTvVBZz27+FzfMSlF1
qMTw0JRMVOqZ58a88SgWuZWmHZnuLzyoJTKyeOVzhrnGRzaVFKvlR3URoMOxCm+y
eSF1kHFpR4+fjcbvKIaav5U5/o3xF04Vy16xjqSO6sGhi7LasdA+Na1gVt0eFWsi
PzwgQbUQ5EpxfS2lIUs+lWWcAaARPZc9qDW5+IOBZ7vmrjd8cB081ckMjPwDRZpQ
7Jf/ZD32hJ8ur1xHApU+7ChIMtGdF/6eH/ee420maL2/eRkBaWmU4/8RX5UPLmAk
T51tzEz62si/ved7IlAwN9EWsas7M8JnjnXjoMq9s2lmBUnWKnz9zYw3FOm7lQhv
OZvAZ0qMbonr/EKFz7klMt0NQIHyPWDiRfMZoNk2ZjRmZErb1BTD8IMpUYa7dfqg
JkqAeOyIGSbbIYP7TRrcL7HiV92+1YmvvfLavrhpYXxHX+38kjngXyEfOpt78FYI
LVGmh4fs2vKeSaPQRnSTk9CR0S6oiPJJXgTW6wHkrm6sO0Vbo/ooScqVLMwtsVif
fCpXaDzgC2W7p+4+jyLpIT49JLkcudesFfaWuRKQPj2nKp1pKdkBXgOpHLx2e0fJ
UKjxc1DSpRrAsucoRrwEwcyOOLp05aM8++ipgJHozwt+YtPrv3lehCNkkLOy/q8z
ulrs74HoGfJsyW0VKEUXfneqmJpipmSt/pZLNNvBWRQHGGpMIxlAuKgJ5Pz6FeNH
4vDo6A8IZkQIhZjoHvHe6DtOH6c167gXd1V9fnG6bwwInLmSp5PGZR+CzL30MVOl
yu1LgqkgKc3nF3CZXlg5xEBK/YIzUgkA8AHOirmNTIZP2akpyMKbnUO29YFWf71G
YOoqzHuWaCdkw7Pvw55F2rsLrys021IRjV9EGER525yjTf3raDH7dHWV4G8MYlZX
qQCa6+N5v1vvGfDpG0Y/tttxHOYvZHlgYed5W/jq+P4+v2jCXLDGXdieh/FdtsTW
f468aXczGqIHMw+1T/NgQmX9RlaYRo9mH2F27qf/u2KwZO9+nizywEX5PvWJ1Vbq
9TgRPPxzMaKRbl8iP5Zz7aJW5bC1NfO1qVdf8pZbwWno7h2xfG20U2fLv57kZrc/
NquHYQGBIfwYnPLhD5np6DaGV7EQqqm49wOvgQ2fZLjZL/wBpbFUlAHk7fMyaEt1
YUgJ7qkELE3GVO2A+7865RPNOp06fEyCaSQBKLtgsN/ZWI8/TOaV/yFB2raHPKiq
3aP5VZnD7mfPqTgem9xzu2OOMnl4R5pTeuIFqrRZlhXySwpn/8JzBxOVZckRDT+5
dTpVVD04dsrwaVLThh5EY6EOlZAfaQyEMdSL0r6cQqMXoIsE0giy+C8Feni6Cc4W
20GC7i39XubxbaSbWQ1hWEHRegOm5mQeYzK3S9/ao32dvNFf6Ycnn8QcCe7Wrupb
6ajnfkq4vvn0VwVR3vgKHnRegGckW3awPrfw36KjqbHxYrzf4Q1CEweX4mLVdCP4
0OxIeQ5q1TYdeJE1ZPf97NakEmrbd2dQto51tAoZfVSXt/Pb5xlDDg+QCuFL6mD/
UXS5jkemvxWd3dmcDj/rW7Gg4aD7ZdHzlGD+MIIK19uBauq8VF4mGvndtCv4v8Vm
pT2Dy9nAT0ouoGooqLU+FzG5f5M7eQWifiZFOAL7ypFIrWwcT10DUyaLDMAhwFYZ
EraKN4GirXdWVw++D4Djv905/vnphS7QRaTndxetgQZtYSt67eTx1nfAtOpdb+qm
A3OyZsxTGsaOL2n1FxZPFuuUxouWapBHp1puo6y/2TNYzm1ywZu9uYT5CdhVn0Oy
ec7dWC64qA4Wx3hmRtS6cZDxyVnQ9CRHQftCgDygvw3/o5Dtarr3YWM4lAQ4PZM8
E9F5SymTznLeZw0qmwcKdvtvDBAY4ENdrdmUv1PDaTgosgS/r5vhaaucQ4UnCJQv
MQVtc2D4RRqxMX2E33M/Ujr2KM4IMxZnQRUS9WuiezvbMt077vfLXLC6FI5KUPT5
SGXlUT6gYV/t9SmYOcZNqYXtci3uQIOcDGeJzxseq9njmk/nONO/7hmORwe+dnJy
LtUYXyvVxqr3ibSAjjgtoE1nCWRS9JQFFrjxbQu/bPXoTU87V9Q28s4d9ryIp4l+
1J7aeeTwYHUfKvrA3+2x16VJo6DhrGoNQHA8xU1ulskQDvekbJlz/g5BtLQvFPKq
GvOy/ODjVZ0UaeI43RIQTQ+oNIfV3sntRWoPGf7K1LrwlXNjmkyEbvkUb/Va7ZQz
6ApJe49e6nLc0n18vBRUezrl2t4AN/JtTksqsdTDIGruiJMIFyvQC4cC+PT8nbw2
cRXXEMmIjlKIWAsiJwTlFhD0t+3dtpzJLQY3r0SvUnwQtQxI7b0bXUiNuYc/syr8
x5JP2Idr9NdUSWPgQFvLH3AGU2vdzpmjiGnOpV2gN55KQbKgriBccE3iwXVwi6SD
Gbe2eCSkxPtpQXW03KiQpHXtXwQUJVBZ/xgR9/Pvaeyp/FIYZlm4z9+oUBTDovUm
tAba8QzN1yXf2PANxmPuF0iXedYH5XgYAcX2eaOYqP/6J29jGEZIl2LmVUsUYf6Y
p0y/BCTKL1CX06kwG9Y74LI6zc1Z7nOhnPnjks6CG4+dpmVZfo5jQB4D1bSPPGot
oq+cbY/ZAkm+/vzITlmeQvIiyIlmLMNYpczdMps5cz3EtqjJMbN86TgZldKaPxve
WFzIn1CbI9Sp8epltuJRPKssb4xBX9pUMrTU29Ee3US+ypuOp1UpTA06r7metGhK
orAUaDDCaouCCs+QeERJn9zD3ymDy477lI8Z8PqX0XE9t06U/wifREteP7yg/63M
pLTS/Bxauv/rqus5cO1wuOV48WR8+jc1ExIqNAWSaLNCA9wi9QMH34JiehGAV2Vv
e1dr2YDHtlnPtWKFVPNlEiPj1scHe3PpwGYALfqJPds2Aigbe090qTKZC2zkf3Le
S0yimAUXA8AUxiHNaIC9/SBr5aWUrTtxeXyLo/xny19JOkt5V0Ff+SR6IclDYeUL
sGw83pNgCqXucZyQN7uEdYeX0my1XxjdadZOc3k+fA7Ks9Cpog+A723Vu+tLUcdf
a010BtLUbxvilJTW0bZsa/mvLq0DX6/FFFmPuttK4S4b6PbokpJt+LNk6kEOewv8
LmHMMEkoAopmQIdRlPHDvZ0VHuWYHIUt2My9b5QT/OKsGmTAW8i2MBj7BD8zSku5
8Rylt2caNI8E2R+Zbi8A/Dwanl/ZpjeLw+LQJ+AHLtMj+wZo4yGOiiup+IYku/SF
9yj6cDSP0P3dm9uJZeRiwk2ikcjRd95hcaCtj8apXd6/GXPZyBIZxhCa2unHSDrV
qwM8mET68NUaq6+MRoJR5hl8c08BwCtTPOeyu+tl2Nq/Q4afI7WD6uduoGecQaqd
wvK3DhxE+P/BFXE+pcRpoTi+xrwoxlH37NuRxeC2PI9twAKXc0TmSs0JwqcqKzyX
I/EK/PgcfD0PhswSba1BIcLAr1jaR7c45CceZ9Bls4fSBuTun6xauZRc4rxWTk5m
P2n/6Jt5ZNdsX8iGVFv8qgLSVAcy3oxs1sNezdG/R+tA8MxQR/y2vvdgeeNrqusE
NSrdAsMhJyrQfeZiqdcVT0aavd8rLIUXXSNd0GhtycvKmW1H+JlW6q47A/j7Tluq
MAgIQw9ORQ/9RlmP+yjGW9siaBJY1LRBdJxNiQtONwIXdquIJQXdaXHPb7E9BqsJ
97zD2UJNCxU3Du7k8mPB3/LVf6DrazhxF+l/J/CWfhfPbQ+ggNEUnefhOy0P8X7Z
LXXjj3k52EioiS95faaD8OJmDyzYVNZhvTQrZlJzaBQ/o5udsdtGSE7S6lpVfjwA
fEjlvciOEEZkTYJ4y1uDTYHZ+mJR0pDj7m8jVmATEPnbPAtZs4TQ3WJQ8qXTuYJo
WpZ2424bmL14XgqW8yBu4TaDtuhi9XPMler/r2Qobp+PnUHmzbCYfCnKAVxLxIqN
LEWno6kAYdN5kPBsiR2a8sAt+2RG4UYmrVdGjjsZdIVtj4NzNF2Y7ILzsWKbnQx3
uN4a1+31njH7o5tQYDMIvAu5uMQL2yYjex1NaOc7OhncfpDO1x+d5EUhvS1KfZW9
Axbuj2eYxMUS0JF/dozcpBF2JU3rZKTJ4gzCAVdPbQYObtjIbw42nux2MZlgm7Gq
IsrRwvrvuNWNNYlw1Xz6XqboPsmJdZo2RNZvAMWCkbPYePRkAIbyVLk8RYqMKsUH
uK1/plCMAGPhsxzD6UDJJ0+xD4gTGgc7YxWPxBml/gQHdA91Y+3rZ2nwKFyWtqmq
GjIXuwQjY46yah4kmII3G+P8llNTBIKHQIO2YQyRMQjIXFISR4+U/J5ONByZ634C
zcgPpynazsphw9WSNY2b7ZmgRSHI7B5E3uS/VpdcTPGiyMPFM+SMF23GEVmIi7Br
FphU173Da9VnrOMopZcoE+UAnRyBJ76g5yY58D6zK8WBdnDoW3XT6zJO10A482bZ
9249wclLGT6w7QKFTVhE7w2mc3fVpZTiVDGet5O6KSBKn6uM6bstDtZV1VZGydOE
K4vfBXdaYHIRljaCa7ec+cTOxRyJRVLlSNRpSj5Kp9vxuVPCu33q6Z/Ruiwx2UFw
a64TvwsnDQ9skni1sVGSt+ABTN2Cmx0Aey3zldLUvxg+KeY9Ll2t2A5brWoK8+GR
Ow/7s6qt2iYpvANAD8GRjg4uUbJ1nwlM5mUARnqNXJkQdc6IUM2PNey/VKSAQr19
KtlkQ6EuMr8f0ON1O49GijMssYIDXJrY6Teg6dIddo86BLjCwKkrvIqnLFZVzK7r
rOXbN7rptg9TgboBznHPU6d4Pe4xrMciTlCPIa6GkRIGQpVnSptIIW6z6Sy2ZVoz
W0Oih9L8GSfSd8JqwxSU28seDSLp77RoT90oGbhSN5q0LeYgOzxTlTm3hBFvjR5o
HdFGWH7O4YY80x7nq4DoJO4vdbrK9YicwIF4hjEGyGBdByG41+pFu+4A7+snH6JM
rOOt8tVuV3alm52x8rjpOOZYh5hLPVlKWVpja07S6sytF0tY1zAzcT4pjRhrOWAT
Hc4OXwIkFiTjEgP4EHLcW9TcYt8Et2S/A/keWcTzKaDsI0nWfQk5kQNM49776kuS
i3Ce0qck5j/0tBaksLUEg4rdJ1H3FP6+tt1vhN/nMLBE4G5Lr8AX/U+WOdydVE1h
kjem0EzjgOrweusxrXg2VoqHh2BQUZUVaFOyP9PXbiUccYhIyZDyancijD+6pcqq
NpgBtlwwPOAiRgAfsTKCgM1oZxSvJVFvQFbb+8XOPXhxZKd/IdisKe2OxmWnwkRQ
x4MJsRZoskBLuvKI3q1l/C1xlWw5D+QFUcy5t13/iadXCBhh9WkXDGmg0ICjPf+G
5TisnkPEnFcs2eXdVaQFLclThnJKBR7+umHlpuJAZ/o1ygZyt5GQXMesK1iiZAve
+GVGUcXfsrmMTVYgEWZfH1u1sQxeJsRAw31LBBPjqpogWPdeGT5XqPo0DFp+ukxt
+ukIH2p3XWIcmbfhoAVBgME5DWZzVm22Tw9suwReGAik81mtLEwiErVqlDIHUjL9
qA69oJ1U18MWD01wa+0r6AY53RwtR0FdZlIOgb96SQs81QaMsUeY+ObOcuBe1hmi
OiD5kxcvkhPulqEBqN5mEP55wQrza3Z/54sQ2ZNE+MTJDFkvf7F7Hp+Joc+UXGJt
IasJdiDMaywkTdArBcyLv/wXGV8Hxrjr4bGm2wvKjdclDy5o9L3blLLygx+YSIZE
OO3xs7/MkU6L5gOKWPFDk9Wex27u/3jwwF0L5FZCkljKT41gLx9utqdIeyX2JnVh
IH5pRd4YMB6t8pjII8PD0Y0U1Ma60crt+m/XugzDm2dSxFYX6iqzA472FV/KV5Lc
YczhEi4rz4/yWgKn8ESueRYzUGw8q7B9Z3EJa3k6du95bwQtEfY0t6hJkPp+7akv
Nt7E1fflOr2ry3BzhrYK6DOhTx/KclEhfakhurNKEluyfyZRLY7SwTD0j2reCR/z
wBKbwIgS8iSsh1RfVDiqKDaJALVoqfk7IW29YHXiE5ZYueJjEXVaZk72I+7s0pl9
7O5RXcVTyaq9Qeqr+EmhtNsgFllB3S2QQxZL1yh/yAXO3V9kh0+tvxvQOs2ROml5
4R8kvsb6tRCvdOROcig6j5h4lXYFIF0vPqZ8JXstsm0lU0Q9M9FSKsfdVk7ywMOS
ru+Sx3Tuq0F3VtqUHLca2PGu0ohH9Z32X2/Onu6Z5cf41h8C5ssHwugLiBYiMw36
J2gT07AWbsIA37WZ7xg57RhFtd/qfUaV9x7GliypvCJ6h5stl8+ifE6J0s3YA0B9
jzYRDjOdKqtoykQKIDJHAmPkRpbITxwQS361rSd/9JS+LF0jWRyWxDy0YL7fLbkS
Unqupq2pWDA3o5OkuIlI1pf2+SlrjUdGYOWcggjGqTCdVr0PPOk5su89BUivvPMq
Rn4W74wSPEcBU6guo7KG0COCbpcd4b095RUNqUOUG/kt61AFvPOWeuWE8fgztoUC
97eVBOO7lcAntr/qUWeH9tUocD50gMLxBbi6m/b7TYpKda8C0Zufj2n/amHk6Pd7
pwZc8jnmNKL7h9HBy9BxChzcs6T2ev8UhHaoRFznlWB0rKy5gSHNh+xBOQJRCLko
AQ/RFnjQUMeflUEjHf7KYs5nLNRGpwht2IB32ovWJod++orXIYngYI8wfDMQDjOD
otz3QU4AKKmVfaEvN/LRLm33UnOTwSWRoBy0aN82BG0paE3qGZzC7yJFOdDPIUZ9
GAPNSRDOuhSh3q1/9oRn9QPa6M1d6SIbNJnGOFE3QNaljLV8RQJbLWxWIseuxPIj
d9p+m3VoU6G77HdxSP3GsJAkv6E6sKWmJNj6y2biIICeoJNUz3UHTB3tPtiB3Lst
+hWVfrrNf+IZ+H+jwcbPaqCN8niqqVAVPAQ5XMbduVrAx63z6TCEYzhJZqayUhlp
a1wyXfxg1cLyeAfV2JCkdvkfyRQWjdlJlU3imq+oX4EJGdtPRHpbApZx2DMLTqXJ
gf43SPNk4tnX+tsnxgGiFl+DOoT0DA9/g4zE23mlOPzXrNW0byNJhF5UVpTzHM9v
pkhXeIPUuo3Ssmny+DR4qcWzwFjR4c3vOkxmR6Ya7jwV2JE6aoriONVUFeiY1feY
osVVh+kjyS3UpFu0R+fCk4yKw/DewVx441xj4g55U44lz8uTCnQmzlLEj+gGWegy
KdzzNO1nVZserOVcHHh2yrNl/SJAKqsBdkq4Edlp0I3wvjwCTXGwn/xwIpSfsh9k
wIKYzip1JQAEvHWpUMmbu6c2xuqRND2zWcD5JMJDOlBtClORb095G57Y8+YziA7V
khaKtbXfiNQUAsfeEvP0RNhi0d1OMVQEKkqM10bhU7BFm++Zyc3VLdGfnaNgdhg1
eg9lcp9hGyzFw24lPO6BoiASqPf8NaQDxRzIDdb9sRHZWghEhRU0Hm39POgr34Ol
dbNX4rLmnbm4LcPsRyIAu6qYumECl5rwZo2d45s/BgH6uDZqwxy3qYWkg8OuFojx
z4HfsdEVdn4o2cujJImUYrskW7V5t/5VU2mtXRKQfrT+Xo2s52ZhmaOa4NDJDDWB
0d+J0cItkEAJTujanNkZARg27Mkf2QjeRjYJgmdh53aDFiLu6vrsDfgQru7fS/nH
S2XMmohQ4nKBOqrOdbqwCaLf50jkSy3RNMjXYN4hgFY61tvIpwtYjWN4u7ObdxcB
W2jjN70scRuDpg7MP+88Aq9uyNsymPe/T0TmHwLbVmFrLfR4nD8kwjfG750mFq/R
zsDugwhitBtLUs5rW2Gvv9N6LX+42VyJWfLHYvMibNRQBAIco+lD/vf2yq3GBuH6
iF28kTk5Xy2qjoU+R+JLxIaYTkpebirSCMHAxmG2YeyyuLPa8GUA5Ol8xd8U8iRz
LuW9lYFMhki6evPTPwqNqo9beGdfnKqeFDE47NFxd5PITYHbTvOdVWKHG+uPIFi6
zDJ3v/npaP2o9jJTo3ZjmBhnyWVt0DOfhPn7T3SB7p0DpAouNGCaUNj+WKGJ0/ar
iRlt61pBCvNQU5WVYw+Xlp4XcyCaMdIyacL6X+TZDVy4IM/jr3EzYMrbc287/AnN
wNCsoyTVH4OBHlmsU2zdxcio9l1NRzTrJzXjaWDqg3SlBCLss4GgKrFUwqPsmIM8
3FXLN49UX/4Y/z4iP3iossgm9l/eDKjt60bmJYUaMXZ/d/41Hw34A0J2uCieqaHr
nzhgdkLM7HrfizmFb+NRNNtQ6JS1yuFkAJOi69hNZi+ihhDsOFW9CZBwcWsEEsgv
7G6sJzWkttyw+m9J0A8eHGG3qwdRO1CHVeTBwC2i3XtECEJY1nMtcAvLG0NFSTji
LfRr9R2ycMg9reFFyPlobkaGPpBioEvlzdpFIlq1hSkHhlak/UVIrGVACiZjinfm
Wvc0gwnkX+aDEBTk87uLiAR9DL3TXCFLVWBSM1u/4yIOLgrahQkFtlBOS5bOiuc0
IiU6e0eMe5wEUiCboql8rg8/clquXb11Zb43Sa2WkC9+ZSunhbB6D1zszCrrmvgP
O5cqLelXONxmyhZMUQ4wxdAPzdyFEbcMcqYGfVY8H0RiRMUn5yn5dY1iPAti2a/S
LTOXIIRJnRiktMW4YQ5aWe1YGN80cbJqYRkSdrinXbUleqJyfSls0dqY/QDuRXBz
vcuqw1xL2wQUidbwaM1bE4q4zlG5FYiTawekIZ8yZed2lhvuIcca7Ce1fBEReB5M
j6QPEeHeaJFERMaBxYvliId0tsrP/6x6diiKqGhHA/sLUk9bYfHwgsLOvTVNSmz3
Htd33zj/V+dExj6Wtmrq9NNFe7xEQUKcztO2CwEv6Y6RAa2tn+V4BV9Bi/Qc71Yl
tob+dlIlATQAf8CgCMWRhKR8ZkuLNnGFWFanuJBj8qNKT5LzRcf+U93EGNydx0v3
GsyktjwDMWH0Yx73h+NW2TRpaG0rDH3y+iIIR0I9ervv7wd8PgbUajZyWtgzaUIV
/InAES79Ybc37jl3hW5W31SXPdhdzLKc+hNdypP0imsiI5zZTx2M5rYVCkejrwG2
azIXw6WK2jBLLDIUVzfBzGgFMLONPxShxiE7jrI1FViWibys0t681oR2/Mjn87vj
gnc/lOinkuVYDd362Z4+FHvJJKULRdcJ30vEU52LeQBq41E5V3AE4dsdNG04ijeU
Lf/Ep8REPbs2RWttr52fk8Njm78fv1Ab/mzMIfZtGd/KOjjhLvB/4A1VnKH8UWBq
EUD6osZ/V1H+MD21dhf3t9MkuDs4RuPE56NML7ghIVN364LwPiuouqcylmlMybcP
Ha6ed2l9CEDFGeTDcvUy9798aF0itLezGQnDFo7p03ID0EacuivftdMePh1dPJHr
dMq7jQT1ziJ7u6lCYqvBqjNFr9nP1JQH1Ie5BaXFP67hlI6sx57FVqDdTrOPd9L4
T4lhrMaCTfxxj0Fbp9TgxTUB9YUuW5DJOWk+pjxZ111WF/BmFQ9ekJ3GPeMJ2YXj
h8RrTf+QgJGft+Ug/bgSHqdfeh3cr7mUmy1VjjIogLqA1g//Z6omMa7HtEpgwaTc
DaA5uH9k8mLZCVKrlG+RwYyTtsuOlzzY122atsEnqVEfiu0IeXlAsZqoKfH8vPvK
UDhKFWBKuQn/VazRTzzBVLx6HEC1W+adQ54pB5mtWVptYYnNuq8tvXwUdSRMrTZS
6e3VBXEUZ7NF6Av+QB0V6ITR9U3V7gQawBeAO/lmaShc/rXk2fVh2FrqjPvmoOWU
mjPgTfrE1ETMtjvMRSQNjFUcKuXb3psUNKdMX+2tKioy/pr+9Wpn3nt7Epxf9d8x
q4y4xfAc+PSPMLHOG6IwIvtvDzORgOkfcNuTCXj35H3updpyFHYisweIO1MTwSSK
zJeOjfeJWZyWbNYiYK8yCTUR2rU+qrOgAvRkJK1SU/kFEYM8ZKSN/q+rdcebr/ln
n0XLi9yeGz4LVyRT1lJgBIhxjfAu4BOzlwvObCswd8z9hboBfLaEu53Wz3wiensZ
1D7aAUvykPIay3K/NeqjwrXUXuePgdIRXK/THAFb+XLJLuYRI51LOmgZCrB1khl4
yXF0GJ1lCq8tQNdVU6oKgCR2c2FItXmcCxdeIDYbfzvX7a09ADgYBt+DQELzYTi5
hSczR7kettftLD1ZlGI85mZUiXcnXvao9EXAu1e6AfrtQuvd/Xcnqpg0ciAYHXNl
csOAALBWpbfHjz1LfFn+We/1+1/YKfOkZStT5I9kPbGbDCGXd0OVZFFQZGmzQ440
HEsaFr2aiEM0q3ovvwr7+s1cpset1l9gIqjm0UCLRG4jQFYvTMTGIsWxyDgJ/BnW
XR6IH7VYp4fe4LzHHcCz1IyQbKPa0/Kx3lH4jSQGWCb5Ag3I0EL4OUj9bScxF79C
Evwp0otcMeo5goZdBFzvHa1/jSP0GKEMlxQgF3khPfuvahp0LfZMyildbvOGtkXu
gYfCAQ/zEJS1Fe5QWp67mPXA5GSeTzfD0hQFWGgCcsVnrSHXHR4lFssPCUqm3lDy
RFbO4kToZH8P3ui/VJsVRSoRlhMltyDCPphpM9i/NF5knzhrVWIMR5uvSAdkuFGs
OXT/MfRw1w+CdWUd5dh2PZSJudZaWbl5Nf3rIrXT5M1PVmeKd0ZOiy+dAdbwJ9ED
VQ8Voo6IzpxCR9v5sn8YcatuTNbb2uvSZ0cgRbDYDqcHmjwglNNMIZkbFl2LKOXh
n6HSPSXqmvtMN3CQZ0wYCEQa/BkHDpYTovDcR5jx8I60JTF5oPPsbi8mWLH+OcSv
lVP1gEeQ6RmXqoMMtaYeCMUX5Ok+ehmvwJdg7oi4AkRiRudqeKh0Sn42rmdNxwyy
moAmPVcplAIG0oin2g69q0tES8kB2gw3XD3WP9/MR26oOOn448uJ1OLnhz4o/eZ0
+Z0W5QKMgwu5k9/LB1cepYH4cmzzEHT56td6HSUXnOSskLZ6mR92vs6clEQ0ywc5
bRGFyg8QkUelwbjhlg4Vs1OqSBdz/J9WYUCzMHfv//pAKwcTIbPea+AEnkmbhBlj
GT/E/6MwcjqdEH1MLvNnr25/PhZDBwHDIsnTSFUu34SG4W7vDzxl1nK2HrV4FoKP
n5NCEhPoO5C5MnwPFPh0iwl7FEdfx9Mxsqr0+p5aslrb22CejyqPHxZYfwzuKcjx
1mRw9EKUwttbRuz5rREy1FOpSAMrRmPmDEJ/c834EXfuKqU0JlETMi7FUuoo8i6R
9R6qg87vkFoxqeFgchE15DZLYs0vVZNeBnPEwldJaruVzrxA4i4Ji0+DNyqfGmeJ
jwrsKfn5ylYdM1enl8Lpcfn6mbFM+Kyv7Ag+DveRnR9rEI3JkJix9qWehfeYh6Wi
VQNbyYjKXpImNmwfSd9hABmjv0f7WxX2vu+0oBS/x1UXqrVZh4+pQKhA1e92vgCa
cbfSPWqS6KdhoLQFKHNmgJLGKJrh3UAva++vHkoM5beGPt7nJBZaeYKc54VH828R
AU5Y0cpnMu/PBVQfWG0uESz1G6SSg4rF//U/VJXuAS8Hpc/qQA9tVJ9+ls9OSXBO
c0ksZZuVXGkLt5V4yaTzyTt9L66ADrR14nLWlIWzNVFVk7ehBqCs6wJtGNsTz2lV
paDwt3B0xXag/AoZYWMojKKvVrtqdXPQ9RQrx32+sMGE44gRF3LE2SyKIMEmVk9Q
evgmQQXbaTWnCSOa6ZUYT8y908D8zZw5FlPSKcO64FMt0lWtKx+PpBBtwn6zxPjV
oYAyzor+mmucmGUR8+Zhd2EnVaCIG0ag1pJbLK5JxDqRqmqRdAygO++kTS8u7Mvw
UyA4gJr8hjAcqrTGFQeOIIGmnjHECxbHQZfJLN7ML6TlRNAYqhLReyPZYhAI8e5Z
uYbv4lvjEp4HP657fPfSxSPf4xcfT6MEQSgEHbTtV1ATVHKuP1d98rmLuQG4O+9L
0HaQywAB4LKOKcdtGKvBsw0FnQizadP60RlJ6tIPk41DjYvsZsS7pjWkUyq+t7ud
YTUSMoKTIgBcyPdVUczYutILU5ONpcVpgv/Nz4T6vHHugfDHGmOZnvKnJiiwx4rC
ibpd3SO7iDLoNmIFHwlEfzuFeIumWkyVzreKOOIyMmFv/WGu1CRa6eZ82/tiJAjt
UtKeZlv1W/u+HCeg284d7igW6ht87cJ9thagS9xKIB/ALSBPyLadOx4y2KHE2GM3
6LX65E2psZlQNSWmVZr6YbINVZtkV0fs/GYxsUKTi0Z0R1zM1XbeVG4cNEnJgxQt
z5ETXJB1W3EM96vz5CHR8vZ+jbshp1VynhPHWjXZ+vnBrWBMEIFq2PCJ6cDT7zp3
hYj4zEAumzIfB1mzulyHPViNj5FK8pncBas8MHXUySldWQApyckCXMFL2CcBRW/S
AwwZVA8J5btoYTx5Fx0gZJv5uf3FQ1dNiXiSxQdUlVZjrJ1MhGXf8bZNaEcNlB3V
zM7UT3ortSIeRaRGDVC1h8IiOsqrmiMwV5aC8N57ZXbWslehxoVIwlEDyIELMdzl
c9PPoy9AfcjxhqPvmF5ce3Hi1XSn11Cm1KqErXw33gV/PH7yLOcVrLW9qLkZuiIg
ceLLfu4zziATsNPVYrv2JMi/TtRzZLq9vAJ2sr8gxiRZdxN7hdqicCDKul3lYTex
05dWmAJYnJjHB2Y/mOmR76oboT6XisiI6Cce7vR4rdR2RGA5XMr9TEmKNOWnqrHr
a9cw2xRdr0HseM6Jz7Wk+xj5oL2JObbONA+aM/mr8LVqOu+bKhAieYO+jKWLr+5K
ZetoRcf0ZArXMx/U5iwjZG3dmK41amQaJg+EYk4jnNKm3vqJFc/rYNtLZX0CQpdX
fB43FdHnYhfCiebPj6vh1OzQ+7t/GIBMhA57Pv9KPCEO+NCi7FJwftkTIrGaWlNA
vvtLIQFeNffQMJCoqQcZULYow1feQlP3iGXK9Fab0UVQ0IAcEZmI2HXkg+gYKkWO
AAb/7SkzmQjqYzwvOHn99tBbKc0NUcCHY1WYcMthYBlF0wM/Tfq24RhradHrH9ok
0UXFBHcPCxt4/u1C3xVFXIofYt1YtkjKveipP497Vg0aZG0p3Es/tGSqwpIcVNbe
ZprIKBVsWLiYsE77OE0rg4ktG0EFDktwwgFYhnme2+ppkqnO3hqbCW+z2sZwDtUx
5FtfMQDOzEpjUT0n3sYf+gbRQeFYCvKwU0LAM7+rwlVVqG1+Do/Zzh/NCgRaeeHL
SvbMZUJpt7iu6lVNIIsxMbl4X8nXPIeysLV0GkAGsXL92pMxQWxtjxzJAwTjZzSf
sDl05v3s4j0vs6gWWZHrhQ4c+9sKgt5B6/70xiWpcT9bev6BP71MSpq7UVjToCb6
fN/TFgUswGz5D9A6f1N8kg7BCUtqbXjoNy9GL0U5TS4T9jGLPJYY1bUBxu08dWQS
uz7tI+jtb5aB0r1Hu7z4O7dhERZOxNQFWmmDo4bfpVHj50xR3AxCAi+JMj3S/lAA
ruaIOkRqnXGcnGgyxjJMpfdPxDzALHcovaQ6uEvAr2DCFwwPZwZDLNS/jWPvfhx9
VJnrwJHPrW3U4xlei2xmUkFMHIUfT4Tpx1i/ysdAe85fCILz+HLF1J7D8z7gX6Mk
42obHcx0ZKxbQTMVDQWM+1dQajtJBFfAmNfJRxuZnCvh9KsiVziP9/da0S/crPkF
6mLNZKyJ98CzZQHoa+J07qTDRMKjROy75ypdSeghPkW5kEW6wNm2/9uVAt970Oq/
ceF9D+kxZUYstpMPdU2llahlvLWHwurGhdPGQJhorM+9mxj3vpQBuLlNxlLsQklk
synqkORYYwNrVLehkrVbxl2o07s2pgzX5nm5IQvyT4DY1c7FDY8b3u+twKsjkenP
KLPtsF/FA0kW6xPtMl0bcAVh78P3Gk36mvq6QF7sTs6LDv6XXqW+ZrVDOJUEBzRn
yt6NlluG9h2+T0KPejtK/a/VfYe9rPCCjs7B16e6ZtHYUMG89q2JSgvuXfs/4o8T
NhgL5hWr48wsSJh1hZKcAo4bY2V+vJZ6KaiCqRGRg1hDDB7O7uOEuxBm/UbZABmQ
zhyAvSOo1cY6Irza7XolyG3Fbxi0by5TWi9JfG2ShIXuZ3Hh0OXHr3yFJFrxggEU
qbvjW8faMbp21eRWg2HF/Ji9YNs6vE4M1vzT0lDEzEiio7QWpw9FSWFVwajsz3yY
bTHnv5QtDRDuTKRS6uyrb9PkRYJ5H2SYM/QUXAjA8eFEt6uZKGrvxWPwNj4KUf70
/IiPxoaoqIiYXkQQL5CQS4RPwxJmolzybCPHW5fl391aCfRUJZPio2FeZS2RFud2
Km30rbfUsXwUbUf5Gb6dgUWTQDwXhTm3g4AYV/y/5Mx83igKveMC5LBbQoTXIzA7
sn+RMh2t9ER1RQJKdaemwbDlY4kFw3zZVyZNM1zG7kxYvKENMKsq+PLFAcXT0uQb
AZvGtN5GwQk2PRWUNrQW0BvWB/qBirJPtqjloW7HhiuSAINBu0Cju+1wzTELpIHM
9VcNS9/1K8cfmmsayv6Jq8uoGnQUUQsjnzGNSguFYFeSa+7YFxduxcpmlnjWP0eZ
NtN6uXlMrpeTGopXIN/lW1gtwYYoH4PzFepYt+sXeuWOKkgfARlbzJiM9jmBCeXv
bQvfRGWQPiea/3PJvhQi1z2qEOJXr20MQp0b2THnKW3BdKwehlqvu1swiVTG9Dap
GBnAnRi+SDfmn4Gc2uPu3ksNpjNWnWXFu33+qI9J1LMUnJXCDjsUi59tVuPFK9Ot
YhLlW5OohYqBCFlXsyeeaShEehSXlp+udQUXf1KeyTM0OmcRplqUB4qoRwERGmiw
E/DafEJpueLvPk3hBTf4+Jg/YbZx/g0iUF4E0f7zre5vJeoTCnyxfD6g2aEKwhhh
Y9n/FEyZOXCzeXNS5OtVv86C45DgXoWqRh3GlUNh/ui74GivvS8LffUGyWYX9dzg
RbWJymSc+/KUVsP0cRK6pzXcTLKD9WUs9v5kDTD4SLemzwriYI3aIbnaDtItv7uq
gs/lP6WtHM/PUbtarMiWUoIGmQX+7Zw3Dq1s6I1tne3PLB8ug0OekSUHwfaFY8IZ
an3KEhPjh/SUN2/a//AhliKDRGWTkXs8rYKJR5qwHHtdbM+TKWcUf1sGaQMN23eH
B+sJmEnXG9Ev9XmudoQdZz+hxxkKp1dghF2KvshFQhptlMpAanuaXru/jwNV8Qn3
r+w3t3wmVVKDZW1qBFGbFux9ilDWnEQaFPgjAPUik5i6nQOZhTIJKDm8T0/EoD5c
+kfcsAtheqARdD6D1AskK151F/grGQA1+/2Ju9p4k7EyhSsxno6QhWHJ7xOJzEai
XdHMicJTDBnRy1ATIZxY5THKpXxn7lY5B/ZiWbVFaNhaLCgLg6Jiz3FAFuIR6/Zi
5z0OKcuay39Sbq0+vp1gE1Xg+i/VjMvtZrql3MwVKfPH/HbH4Mx0BXXEtzWnZEN4
1ojGxeQxnIRGQclFUu3Y726ETPKFkyc3HHc3CgXHTyEZE0a6IID0iSVzwbTF8HK4
3b1kljyr9Te/TIAUNVHmQ1lXZpfcdkQUNDYeBRqH+J+XXHQjcq9Nd6e6PrgwBI9P
dJLfxxzlZk1sQpJBcZofE+dzzvzh/68AcgLPeskwdHT8Ub2zSAk+DY9sIFKRtr8m
loLqd6ZXZeCw0RA71757t4dFKgnP03yV1UddMC96xKs2wtbChtyMMqFMFlcg+/d3
Kh0iXhLuNAnsh+LSp1WuIT8Hw5WmAAJA4Bg9sQh5TqQfWklxO4QIbgR6rNsfVokT
e60lv7lqdAhshDtAawHaZ1mtPsVtciYXn17fiw4Pk1+jsrZIpXglLKSSLHb4f5gQ
0+GrDvhaBZ2mN2W53yi6Q/whbt1BjwUF0TvA3u5UjZTYuzcycSeGoGfmOhbPWQAf
oyohPiDVDO1lVifKL6RHxrcaD9U5GUl/VMtd/3bwAaV7rqf8ABPoIFltI/JGHqPG
LgIuf58ZKPMnssMqkGIRPkV26aO6JyfS5Sv4P2/o93bWADSunwUYtNHMNppNVUS9
QBGd613dxnUrolDSAWNCPzh4UnLr6LM6cdyl0mrwUUGvO0PfeEy1fi0qdtliSN9e
Ve1Ehp4+cxeWy5XvfPyQap1qVIkYSJz/rp/Yo3MBThxcx4L4ewXPiGtmu3eURk4k
YFVlhwmH+N1tw+4+OpV62m/mDWTa3BDDFukcHuryy4Qy5QwvxiIS/kqYE9QIDy1u
hOJfmPVXS3dxq0+egstUCwsw5htqfM81vYdWljUincmyfD3qTRlPgIFLfxyPukDd
l3iAK5ULzg1T8MQD2qQkEqwXafzd3CbdDVMqhhqK/qCCyMjDTebuLs18ExUGEYv9
zyBkzmF1Z2HZUzFtJKJQwGgVXI9fogBXb6DxqRGoX8YOjItbjJj6HN2ESLue7uF/
JLhZGPlAf/9r78tHw4F46VRg8N8tU/XbzgFi6ZpfSDW+mC+H8yqJ3YLW0TOJIxQq
kN/MtEYNfJIyB2nVCimtZd1LiWdMU1hYs2MkagKVBsqytWYnhS4kLFja4nSvC3bx
3vvdAIC/bie/7Cm0CizeMAQ4lPRpeo2UcfwDtO9Qn7XiZ9tPBVawIVuEE61bdGMC
rnCjlHT7bBBWIUs9RR00yXWeMZblV/eecCiQhUOfmXqO8IGEMlYM/y9LEHhLdUqw
uHzdWvO3hCp1+LNI1k8KDCGgNAPJrov0IhZ0hncbFX8oc+xLnGRsKj0N2+Sb4iQ1
6EBFgxs3G+bIa8zNhbijoK2oIDjWPgvhMU9pSHyG+dzKRNwc+j/DzZQHQ84WHQQY
zk/9tRQ/1ncu6lA+6xFLy37uxi0Xqyyc4KOqzP1k+gdk87gtgxKKSpi8fg4S5/h/
jZWsY208reqzdTFJruRwWSNOrBhCOj5+QUnOOCJLXunhHiyLvdiqnMyh+f63+wBo
ZQeYMfiPMN4Qw06rtWqMe2xBer4NaMe+M6FR2LgXlgC33J4a1IMfvzgOF4/gEuRU
2sgtJrH7FDodzRXfVECpTkEFR9nRDqYuXH9bm7QfjivYu9szmc2twAND0btyaZ7g
boP037guTjLoa29RHQMeh+sqAWUjpTlODsGLpJQAKqRxTZ51fFDjvcF2bLu5h15Q
53+lNVMAzG/IgZIZm35Lj+uxMtYplbMID1qkPeSUBj7WVTF0OHq84rAOjIWJ8EoP
nc5Df5pdOefR4TlTi8FmB0AdkF+K6Ds18trMZDCGoMsIAqsNCEW5jaxv3ibDqLgJ
PSUf3C/Z3EaHd4awOfs4/42I09HhFDUnzVFM1NoGX7vWkelROXBqtIqQkMA3zJPZ
euLQqKzhVRtIyPl5BpMU21nlcmhm+L0UksbeGYV+hWAYofD1ECkqGSs45tKZ+YBK
1/NJiVWwoLFmLXo8E/CzHc9MozXCyRrpWY3rH4yyiVNVzpJIha3CZZxAyaHRsct9
+PMdF3nqi+wtwNcjDg9CjK2l/62zZ6+aIegg1V8OZ7+THGXDN9d7ucuF0Wmo08JK
SQJb1onc7wwyh0Iv2Bv3+hsjqDSOZMiyZmQFu04p74VFyF3vhAe45pCz5HHEf5uu
6iBUb3220nRhxjg7qckf8RJcFvNhGQcVMoklKGwuMRKiZhBlQAWoYImKaGMp+fos
05qOwaccTccwyVvu01vjqXF39lqiGx5OFb29ldz4ilA14CoPOzVxGdl3xBgRrD8a
IWExwt/wTNCcILSpZ230d3t8dQxHkkjQDVc83FPNUL48BdalBNcCPyJwl9i4uyPl
2FpZmRggztRkBW/G+NzTnoiZvUtxcphhr9NqlMoiYrjki2Q5M9pz1RKhzFbZw4VN
sYBwic/6uoCHvxi0Y+hJJX1y7AUcF8IeB755A0J4ZLMkov8pcik/cOZ2AJ3nCOLU
9hZD+hD049PbzSc+bIQ8Kd7zsbfqr6XNAXhi5Nq4gOGNyNDweeJ55nBmqFZmHaaA
EKJHvhA4kIp3vKAIk/KWIFvAJdhHNN63HW0eFfs6cfWqBCatYVPfTIRX6F+4kRKO
F5xYSuOeTLfBEu1060DOhXXvZC+xeJT/xyV4wpgoSmLD+ZjKlatsE+xYNKzeroOx
R1j2o5SGsm4obt0y58qWfQQXtyTQbmjAXhazLk0MUUfioyKD1avjTdl1P8Kd1ITA
Q6grdqUGJds56ve3DjaLaIxsKfcd6Ur2fTW6uPX8SJlJTz+ksE9FV02SOHVDoHRl
rHCT8OQHYV3vgm5fT6Gf3Z0BiFhIdQlZE4wHGJscdVlWS46WmE7dIQbpCBhWv5Fd
Ke0phxEuQ2oiZ85UBkjhcl8sD9Htgb70Rcur8ciaPVe8RX9JC2vdaIDJSpvI/GZG
bawh8QAIRWuFhRUj3h+2U2Coht8lvOZQXvrW6NRT+mAuz5HwAbFBEPLnoNNhJ7sU
2z19WwVVcMqPUld9HHTp5arbo4R8ThPlTIkkWa0xesR4zgF/jmic5zVbeiFh58Md
p2hIF6+bx7qxZVRrwbXUbtrM3/XJe7e1iGUgmR7/apLYfzVnzfxzIFhO6GJIwpLa
4K2aGb/56XiGVVfYX2dFiMaEnKIRcOBvcp76nmkh0g7e28v1sN0PXAlou86VD0Mq
9iaSKgZHJP9gp1ZvESCg0isP4vWUrCEg/gy1RoFZOx9AcFfhdqBEVizlUPsOowhI
7YWCIht1rJ/zsZHnnRRFloOd2H8LVQDvyyLLrmGYRBkafSMazceoT+6uoVO/VNUz
7kZLdx4BP5XN9kYWklyY1QKCrSRzyhuBwfVGVlszKguRGNI9nA7IQZ2hbIVDBQ1M
ieoqPYaiGEgOIlJufv9JHJu4zrHHYnV1EDVUMmPjHQAblU1JTbf4qLLY74aKKjjd
rfAd4x5Qu6m7qTCFyFmoJWYTlYcxLFSfYMZlkx9yP/PRi93sCB9+TXcxlUxxp6GN
Bg1Vlxh+rpE8IAQIJd+Ih/6I1J3Tf/dPRB9XJGECC9iEKrFxpxpHTjNViMyKB66l
vTPA8uyl0SaNMzYABTLhVANaIoVVHwbMMlUmOGNvtMgM9QK+DLnNyc3Dw+hSPfmp
ZJAJcrNIiWbY9IA1ePsB1isvH8hM/k9WCAjs0FKA3tTSsEQ5RKFZjf9vY9MWwA+J
Tnga2d/xA4dGwIE7O4wrk1j44JaNtd/B1ycvOUa5ggCujiMsXn6yTf8Xyz4IcWl1
2rYQooHnfvRC2jD9V8k0yrhnCdJzfMyT97ts/e9QABnk75OZUl3u4TKmT8vX/82p
P4kXGtGlg6fc4GEiu1P/ro+Vae8cshATKNBTrrqwXaZ+I/KujPEOqlGJZsuViRWG
pJmWoeT4zMYK89QWz9eW+PVrkydepxVa9j/WL3yGwDi5HHYZ1r5EYW58ojRxwLq9
eNIR2uKiyGXxz6jJX8GXTpoQ6iBNYn8Is9V+8Sb51GEbqbYgM2rJPBr1+5K2i7JE
Vx4WL/AatPwIBHo1DAIy/bv1Zz2wSJCxoF7j464UhrVndqLnh2ZNarYBjb0FvMSU
ucVWlc/R5m/H50LmUO4HsEB5JQjyY9VPDbqrcomzeZFn36/67sg+iHMTXgb32XqD
A+ln5UzNsIIS6STHM7uOkDbmBBLuJtKVX4oh1hVhrsgGiK87+oUId+WHvj/Q8GSO
68/l3a2Vs0v8KUNKRFhlMnrNTb713DG5gJu0Y4ECz/MBgty/R/+CxpIXZVSpZVKz
jePlI5zK1ph+CXzW0fCCJR94QDpLTzivlXTdvV0Wt8aYCOReUxfBlePdlSzuFVD6
5OJs7ML86D+RcEuXfMBtHJB6Yw5PMYwwEHxpGn5lY6btVvkzCE50j4x1qYju0xb+
3W0a68GSra5ZVu+9e2hNU4efU0pt6CwfUUHeIbUpJEE140FSwiHXWEzup+ZbGwyJ
J3OP4wZSip0GuU2pMKajLGjV9tEvtcyMWq9lNaq0KUTUKD12nMRBDVL3ZOSgbWof
aoWgjZ1LnvS3hB1w8Zn03YEq/nsQjHkyRlIJN2/ASBSeN/RTYB/nwCTNqSxIIOIn
5RXS89qR9oxZcgD89xmMGHIrpVrbizfnqkMWCX4byfSb2/9Eap75hcQH4akdIjyA
ZazW6syiF8w1uF12P/WF74BD/Gd7r9rEn60No9EJICOCSBdcpc0NxRGEOovTwa2+
QjnZrZjhiNP8lYHL54H7KKG5dEU9v7Z/A6YBk8tUN4CPtmnNXnAazbmKceUqX67o
DEYvX9BoV/jSVY2z3grgufp3dT1cvl8deTKgnSLIsjnpuB/XO8bIVfHNcJJxAR5F
Te0K74U7zOfGj4/V+p4iu8EfPJ5pMYvxG3d9gKpXBcS5S61ufB7gwxWX5fxqqz4L
K42HUC/17LTv7odIJdp8MoAI++6VHNyhR2uCgviB/kWyCCM8l0bJpYJjm9Mw21Bv
DocLqFSt+3fQYAe0t/7PJ88OkHA0JGVCF4etrPnG8a+2nQjAf3egy43wy4/RMDUj
SeVFC5TnPHmFrVttEmN/Woq3sst2uhrd8UbR/BwzbDisCTKK6kDmCFNUaIymDy5m
qdVtMJaCtXmvteywO2ICnAwLFxp0GAjgCYHM9eXaTqJnv+7MiDMFw/kzIyXx/7yE
aoSWi9L7kolG14q+WPaKxjSyePf1483moY5lly2IIMp/ebKwqPFUSr4f4vX1Bbjx
l6rsLAgNH3ioCtrLvEM6+qNpUf8h7NJOrkVlPluncDScb3Hxv4uuTQ+9CDevDJXj
Vx+XWOmvJbOdP8I7/POiT/LlgJhUEePeukzo4Sae7Uc6jYRFdP2WRwdgoHgAkwNV
uRfJakP3FZvigU83LQMUNu04cu1jcXOK6Bu6ETQWWusdfguLgkmobM3NUwbKyEs4
0RvuOt/ocxcbdz3lb/747wftHOcK2C/84aT51jLmXKVn940cVCSpsEqCfsJnzzzp
7G7TBZf/5iNcZLpGRCQcEzwhh1sWbfwD+WmtJjflQ/mVw2kzEiuhDJOebtQhvk+2
GZHSJhxNuKZOaXqekgZDvjGOZfjf7yL8uoLnhkIAxKCJ911wTsTeP52pjGQCmg3k
LFIGbVpKPs/ETmGoKchQIibAXPbaBG1TqnUjZ/DqlkDgqGr6ceI+PsIkVuCnPdVR
ewWyJyTr6VlleAlu3P+S74g+Os9CiNS9YUi1BAtDMyPyvwGkegYFfzr4nv6ckA7j
PPcGqPElBmhM7UQhhBuIK3x2VyNlgk/JuiVOguoju/cNrY+Z9Vw2bOELhd+FBnAT
rMkfQ8XpOgtOly2zC9EK2jt1Uqs4UWzt6VfwOSz1ix8M6j5BZCKckM1DJINVTvmA
vIEr3HUFyhPBUz8hS1Z8XtmTWFMjRlrG813ekyKgJa+Z3AuZOEDRpvsEgo4pt/9i
wrFw9XVBgKRWDtm9PTzUipOpSBWc7+cOECWZb2dkAcyReJu7Gdz+MDUEkUTEiXXu
dnFytMw77+SDE5FawuCxkGBwKma7ffel5bjm7SFo+BgusLj1WFu802HkWREUnV0y
9bPZJZ9ym55lOVovzlsrjGcRY3vBBdQT11y6Moj0Kw/dQeYJmNcKBTIEADtIc5jG
dJXU0X9Id0Ua2fNnKeRruXhBv5hjAqKl1OhgFQopMCmi52u4gy57mxTWiV3qiFCU
xxPCrr0q6VLx4sYweUKDm75FTCp77i9mFxi7Zet7yw8SqAvAuABLihJScwHiFGBF
ku4vhEc6x+Vx/uw+jGRq9Dlhn7CCM/V0uEBHgAAaKPwQJPQU3c6syTbnDlESDPix
v31uf8LT+Q3LunUmrh0BPAmtTKiibS3yb0l+CSJXp8RqmhF81zZaN7u2w+1DoOPb
nepq7SdpqKluBrO8i5Z3Dbp5bzQ41V/SoiX5n/l69GLW0/4yOLB64iG23iUnqMcF
nNLGkQHVbIopz1Vmi+Dnfixkh2tYqb90Z5FZfzQwIX9Z2359cKzeKruMJ/efcfic
j7MX75pxcDjlDxy0d1WyElZdsakF0hf8xphu2PTCe0qctMz462o99Xq8XmIHgVfL
c6Jw+cYIvZDrF7y8LiDXPJbmxBHynwmpb7icnS8qFCGjScYc7unZVH7DmKXAgMyd
Yhr/6AJg4czySoAA5WqSs11LXKxjQ8gW2kxL5l7r/jxoJ9DQWAOHgdz5d3QxzN32
hLxeN6RgKkT57PfczaKuGH+9rJ55Ty2585IwXz43/KUFvUxVW0vbU2MWcn4HwjOM
iQ4T1VhVCd72KqRVUICflj0UAA1bRvOOK7QmCPlwJDuiV+/eQNWyCfiT921KygJJ
b4lo+/2ubNFyCQOfz5jqmB7AZ+jiI6PFUJpZiCYupaLoo/BDcUyijKKzFmWI5Dh2
sAmiLCbMvWqZgUIhViMPBk5dJ8CqXXV4OOT5W08ERT/afGVuucA5xSbT9FbWFtpx
xiBRgy4qv8OEF9ZFMROs+M1zfd62uAvJFyQAg1muxD8q/yED/6X4nu2hiHka74cr
6sLZkNRUUbcX43DYQfNV4tSKHZCyKn4t6roqLKENqlVmAPUs9bbsVUnD6k08vZRD
bgbZlvBky0vzhwmUM/BLhx6/JJn+msbC08RoeIjCmJzmjr7RlL9XzY1P0nUXvu+9
69HzIT0IU+iwAw7E3RSqjDCfVEAiYWRR7eIWGskl1/RJf5ZkQW3XVEB8/r9vw5tv
+EiHXRwZBe/sJHAtfYrN5GWlFxMgHG1DFOrA6v1nYT0m7E3h26FDOkWY5VFLsHWR
4GLSXiXfSNj4qQO8A72pJQGMnI0yrglI+g2O0EPQsUD9NIZ3/Q/sIqDjua9ccC3q
5IUgfjWSIUsd7wGzR5s/hb2pJBg9zrIi0BM2Ta8jUx+bE8Bei7RGnaDAFEIEduf1
ErOlPtyFs7Q9uaacNMsxL246MNUy3MlR9LgRMcJ8aWHZgn4tTxxdLLAdhMqupLdj
nsh5Nev+txJAayIAC4KQ8fJ9q+qWQ666EMqEh85w+TcJ8Qga42+V/5nYsmFp+bnE
KlCyFdqURK+x8adRlihRncfiB5QRTO4fKWdgVyXW/tHCPrOFDboCllC9zafas4k6
Y/i4cH9NhKb7xwlQxwsBnrx+OzKdw8G9Yuh0JCzF0nFx/gFolTuIcpdZD+ft+BjL
h11wgtJxKzj3MPTrM4z37YhAqhZQHVplp6LImEfY0RmRKnYF4NDTsWr/7CPWuURL
2BhbUWcGDsKeORjw4ZBKgcviBMfw7z4eUn/YITy5HKDa1yRlXkWZrh1uQd1p7DKW
KB60A+3i3WjjVk+foXX/pubAdavDu2WUywqdvyweMudkbpCq0nzmTtu1vPzlOSrU
zshh4igzl1trFYXnWby9sUUgdw0N9EiL0keLUSO2ySKdiy4mn8FKG+0RNzmfEANY
cW7YA/wnyHtoG5SQNN0Gw+22+Y3v2cFAfLMjI+ZcmFI0YrLL1SpCY/zu3x6ffplf
xRHnDK11kfvxnEKAJ4x8QHSUoS+W19jrQkdzyjQ0embsDlt9PtNetabzav79gCqb
PoJq65mlvjq3NGbISaOwYCif6Zn+8lRM8Yj5oDdjeOufLr7RUw9LQcPClIEMULgn
jg5/EysD18h9N1+n7sPi+qt1fxI5aaRhmD26A1hVnHWARATT6sjClQxcUNEyn5E1
8vy6G067XPRhjpXd9nP5Sc4PAymrSV6SbxHb2E2JohjXG+fX2MocmtLHQVE98PVG
SWafVateKRXzgETJFX2tdJ0cQOw2wptqMxgtCjE6v442lk8FrZ0OqUuCUD4vtwlo
6WChopxsyqhoLTzaRg2kyAkG7gJq7c5zomIWAbNzpMJtOIz+D9auP80o1GO0QcLJ
S7cey6izcS2+ovldyzOlBkJ9+XPqxP/xv7rclptNgVKkwhK/N4ZnVtVAzCLU2yRj
PfpK/vetmaIIGpjiY543x5UM6EXBIcGQlkf6emCMIS5RWB6yCSemPXyPrtGFTZP5
hLTFQ68yvPOw3suyRnsqDGzaGsUd2wTDms2i5PHnx8JoRQ1Aupe0KwbAeaI4FjdE
D8Ply97wUu48E0TdsmDh6zq4mGLm0fm3IAJ1sM/Kva7z9JmvPMfW70AcNZKyBpZ5
qj24WX77h3hBfSkn3VCWx0I/6RWfk4PHbEB6qQ+VzPTQjaFjj4wl8e9ZbheXyfhX
OEAV0y4TJqM4SxlzlWscas9xXiNfFL/OdKzvHG8JqiqlZH1isH8WS1WggjpX3gL9
UnxC7bgg/8i7ldLuG3UkLP4jwf5uuYZjSatsKXLjpJNbrTO3fFHcKN7vLjSB+hTo
sQ4fSqPEMohLwUnAOwOUhVg15iUuHirRua0Rp6OC13q8Wz+z6XWUJnmdnpzidDVo
QNvTa4Chw3CHFkqHa7BbWTVoTvH+7UKkRB/URqstu6hvAa2rKH4sODPDnPC8Albc
G2mU6oX67nWcrwtgpS6kfwp+/Uu5Fe8THHae4y4/v+KwV6aDoooQXZVeb1M1uo1O
KPH0A1nrpqKE9JzqwpA40TxWBIciMI8WR3cPhziz1qW3YZchCOESSL0cKUkUNlpP
C5GruYapp6wbBzwAWYrkSDLRfCc3Tx1DMAnR0jvDFVHPVR1EN8UJ9aelSRsR2FX7
lxcJ07dskGom/X/FcucWT1UNZBpgEhWz7ALAIO0JMIEf3EaL/31cWo7djxw9hAuv
Is0Chimr1xwCvr3OW2cumQ+UwW7DCFxAdkFcylrN1xcR0B6WaXgYodc0OJ48yOcU
uKU02CRHJxFgeA8aPzHe7D80WnyFWcjEGkDmCkL+LOsCOQqy5Pk/1RzsIo0aUTJn
pT5z4UcY3ES6FwmiJe4rCLUhxgisz1MGA9qKgd5mSlZOVQz8cGgPYgKdxDJ3vSQe
6Ha3SSRhzpoqkktDMUiACM61j4J+mGAsxERhcPsFSl1ARgAG7fV0Hp2wj4G51oyH
a/4Q/nLTZ+LYBMAiBaFtpCcu80ET4kBA6CW217BUHhrT4npj3rva5H6du7pXNU6r
qi1feL+tn5OvXaW7V6oUM3+eLZG1sI4eeOkjyzpOwwY+s9hK37kuPPiWoqqquSZn
j+GtSegbDIrUtHyONI+NYA7M9f5SnDNmpjryJmZIQ3YTVTjdvHVTDCTZRZtqZcIy
HtAL/LfyDyq3a0g0G6+6wpHVfngy8PXVH9XIibz5MkB1K0+RTQkoMu7S2qo1xnT2
fJHDG6WPZ7IAnuVtNU19+9ySE1BXleBmcuJzglaRxxZGqNRAD3J0yo2rD9Uz0mCQ
N3MU8FLc/Tjc45U8S7BeRWHJpH8ph41+kDcd++/qJiccn0nwLxfadeldlMJwNihc
M2jMUVKjPODu/Y9a6zmWh6eFqKnvVvnXo8GTMW8kDT7skwk2beA8wsEOeCrG3QFB
xHEgpopaAh/DMcGxbI3zlU9o2dTOs0u/XjWpP1LwetUWygOkbNQqZVKysznhfFmW
DfFMrrEEkiU7XHiwoFmq1SifOstJVjfszRW1q0K/yEeCApU+w5tG05M3XltUi96Z
A8Pol0DJeSesv1JnDN9Z5eP6yoXc0PqI5IbZvl7UbGDO2X+JvsL+2gjy+gJz2lwy
I9BPDT6fuVb/t5Y2AwPm+IfUuK03OsyAYwFx37w5Cud6j4AO7mIZ7tmxDM8QRWx/
v35sLlErtU2HB6qwCBioEdIpd1sN/EMd3uLYZR/cfMDjnrqYwIxS9Yyn+okQy+jh
4EDmfjH/1RHYv+v5sxJXJATM+LgsU4aSdGvmEg0gmSaIlPonKS+jBvm5e1ybtFkL
L59wH3ZwXP8diaUdMVWsfmPTNgzzW1ToZojJKMVveONj4kZ15ausK0tdgLcWQ2Vy
p9ltDUkdM+kZowMrClgvbiKijITgPHUHhX+zQ8gm9gyX6C+Kzs8ARKvv5rhFsRxb
NhY52XO2a6OZSEvKL8WuzBHm8q6KV5kxHNxEbLhJ/c3awoBXjs59vtAq/dF3KXWC
6GzSVLui4Eo5LLIXfuXGOeDcuptMaxCj8bwr8hrBVq67CFb922cgvG4dtD6kxdKD
mn6HWN3IeG4MrWb7ua+xu5NlbgW/aPk/UvGEevZ+9yk5CrmOISckXC7ikpM1AeEI
whA3GdWBxwEu/LcAamywMk1f7NVtygn7OQWGlhQL4RqsGZYw7BFTxec0r0gaUT0G
j9OV+WRnaj0joDlxGJD42EJvx+o39/Fdnh96+C6rD+Ms+YijYOc2n+CJeBLhX+Aa
sPlRqL2aCh8fMxtj9m4jWp7ZOS7ebb1/hh/vJh4uYHrPznap1mV/XC/fZNmGdNq8
exTFX0+1Dg2ft2O9oOk3Pc84LpGe5Wc9BrfCo7S/yMBT/lDD0WtApJN23RT/wWGo
GdReJsZGOD+MA0sYRUBvM156F9cTTtznp8Z9W8WfOnd82nvGZh6fA7SJTonKg5DV
9PhU+hkH5xRoO0iP7QGTZLYEi0Z8feEorSDw5ThtUscQmqNEqIYQije/0KR/UiZJ
TRAKckgSrIx1RVpK4my+k5B9Kf5P0ngbnG5oWvhEFs5wbqFbQEq8vijOYyYaiTXL
73JKwjaMHEwEItesKgO9mdqqQWXVxf7PdEUKz0/w2elTJrvMgUrBiUX+wwH2n/5G
VtctPrTX6Xz9UPQFw0m6XGHFk/5CvFi0RoiTrFlcvtVl7QqKcv3z74UFVOXRW7N3
hLTriLm2Dq/0uCmPcIL/gDjA7PWbs/i0tvn79FZFH7iNjsj0JMmhlGyk+tkPrETd
bjYGagktovWWAbuXknjUidFsp2U0u8osrDytIL1VEroiUtRPVhmQmdhX5dhecQgO
Wf9GnsSOqoLtmwHddGKLhefMzXBG/5pi3YJunUhHsFxxAPtywtXwgPJcTsqNDa39
34iTwj+QPQrmlFRYhYLqinK/n5lVhaKUML6WJROVBFwU2xvU2nQth1qYc+lN8jbV
ivtcsZXclibPsQEcIdSkwQb5X7nyHGHFgYScL5w6S1CcsAy7WQv8IDZAAtPb7d1U
pZxgr+yA9U8dJdzw/6XOsl4y4r2KV0FvD2Agyc3ZYoR0J9bYP5hKnfFtLw5RLIAS
2MurisKaPzDmp2qsYeeAR+WAywuZC7CrhmW85lw7NzvNqfdSzfa0qJWHlbg0LZqJ
/CaniFrDXprlmEfxM9PTygON/Bs86eRJXeIDc30y2J6nzrhbXW5re32tiBy3VXfX
ZthZudOr5uKRjhv4dPHQoW+JeSgvBIaQKJtKUTpvABICmeRV25GOxKGisQnvjd+Z
ZzwVxB1CtbG/36Ve0u1DdaPg1aq2tjLWI1cw0ZiytH8dJu5Q5HFLNuBDD/wZRcOd
0VRbWVhB1m+wB2znrrs1Fr6w4ECZkaaUIGeKSPjEXAnXlPf/2M53sQm7Sp15XbXT
qBt9vuGoLUegDuWV/gzk24hOp6kPVOSOVXPRuJogmdKNqcLs9HZmbwYCsWiL8RoN
cHyOzmPEHG40p5QqPMSp2vxKdsi4CqMt6FR87IZNJ7Xr2rxB1LqCQ3HsLpV5EJrk
ylRZHNZPxHkUMVfe4bf8jPJ+UAxgi3Oar+6kRDsAXJK90bbNubdi0/zysXzzHA2O
ugXzi7+YWnmbfAkwFpEAfjVIN33QD1wrB5Pv/2eVgC68QM0aIfMplLedfXcoHnpu
NkWpCLDYGXWNqhCQ56f6boqyB2NecB/ApleFcSY75cx53DYmhEWQi97VUFjnpS1F
xwPm4N47azal0mWmVRvJ2p/jJPLvszVXIUW39x8KKKIRZ1QNkBI092j7+x9LGzm2
ApQiuzIS7LBsCuRyN7T1KpwHVV3nk1L1V/PQpwzEMML0KfZ+Ng+wINB+nN/MKZr3
Oc8ca6uYyIMBnMx7u4e6bk/gVmqCm1VNSZR261P7+/SF1eSM5l1WbbTHaO5tshOR
hsUniheuiEfo+6VHozCjfN34IUzkV+RqctfKsIL+iOZgLyLgudTtGzKKuZz5KvtQ
dWnE4Iifa+fwD8uqMvhHuW1RmAxsSl3PL+aY85hGyXg2H6Upo6pBo4f7GNKT0fjn
RJFsNRtR/da/+ZRNRxstVOlUaNyIActqgILYKg++1tMyqEiJEGU/9Hnsx1q9ifeu
DrAhZXYxMPIEIEz0YfGwuCb93SQLLgOtkY8KtO+zLxPKYtf3lboRSK4MgRlRhbdX
2Iy75lSfOYwXs40of3s6rMpbOX8F5fnbIXpUKJbF0CSeBQX+oNfVK5os/apJOxNh
GaTewzARHuqmNi55awVx4aosKWwcbNwhBMzBp0Dm3eCnXoCoj0XcDyKxsV8wdc5h
IFYRC4afi9d9LoiGw9CYxQ9Dq/lTQ1koPcK9qcpxBxFaaowbopsw2pgezuPuJ9aI
rR11QEpq+WmTLn+/W66iGjoKu0jCJ7ts06mSTyEPJSsmB/RBRnO8GPywk3MBJBk8
+Z7cpHptxDiQ3yKZXQzrrM7JixQjoNVeICxD/qsTToLodIKLZOppBrMCjr8M1j+7
M54L9kfh+yFXwTkMy09xt+vj8ekzmDYGghePuBzWE/OXhdDIBJFaG5SCP/2C3q9O
kptN6RrM+QOTw6bIhoNvoMKxDunMwWnWhHukdOjPTUDMQBe0DzKoNifKh1XjRxNY
MxrgS1mSQG0IiaGTSSEhO4sgjHuOaO/nswTDQA2CKAi+NxyMh0inZ8oy43z5LLYN
FGpxApn+9cddCy7bkc8SLxe3oUXQBbpJOm8CHDJzXixj64Xwud3jCSorEkJaNvPP
uWSdFiPblFLlQVFMYp1rwwbMBLY6htNBVV8GOzHGNKhWUYRFg/f3ZT/9hiAQaFl4
M8hh91T/IwDOJGBMUV+EFrp+chHCpGOElLqzqnrYdDBsjoAxUWLsGjiO+DTmgUhq
hKCB503wPPfIyCG3vhPuqcI5cD39eARFvAka1shREhwoD0SAWk6s86FA44mNvoSR
XkYc5YJwlPg/GTi0tW7umeXqx2M0oqiOSdvLNqLOL1asYh+5Z9PFF63MGHEr3tjq
0EHlvpkEUwoidbq6rSPCqU7D/BKdc9ko6EKxiwLjVHeQxYY4NlN/Eth/TG2xKK5X
rC5MRdS9l0ZwzB9Teglk8KWEoX/s4fa3Z3+RH7fGknUa8kAWsThqztiTUCtDwP7i
oMWbCaLK9klpOCZHZ+gsJgB6uYFbrTyQ5P0qM6vK+To/8rLNnbUF016Lqx9soSNB
2rCt5viY5i8FABRQ6t7zdm1l3BE0KeM+tUaR/IPmS64THRSX+IIJRE+WWXUNVTl8
3NRvYc57uRTN0ggAEXFEC5uNeVUgcLw3YOV57+290Fvp9pTL/V8dqyVfbV98LKj9
cEjPogu8h7E2UCY7gUf494mTKGdB+jjIrh+yDi8Ah95zjAxkHhNAkuu/HxFgNeRs
vF02o9QbIoN/zPmu9b7h2TB/9rE/fvfSFndSLukKcNq0/6oTFGodPx49gG0HvPzD
5muUIqjbjcLiZNiv2pfQ9nkIM6GBIQKEjogpIvLrXcCukkCRbKQCFB7CWo4G9eBg
f6sqe1qd2jQB7w3OKXhbIqq6vosjNxWK+PrW7GGWmnef6oYSvTZLJVRUMbdzzD2M
/namp1QNCluVXSD/5E1Q5yX2nQ35qv56TEFBw7tVHAY+6/0rezlOsi/gTj8yXOqc
jx1xDFvAMej6tH8P7NaRASqOicBq3XpP6mPlBO5CbxqYoitrWYMXPWQJDLE4aASU
hheluEZ7XZdT0YwVph2grc9akmiPQ5dNIaUm7SLIH/kC+YDAX/rgPA46RAFrbLkj
KeuSfvVMr+FLDqNcOap2bbH0wfWrL++IvQUJPaEcvvBJ0o5dF5O/d9AeWdzARGGE
RfdbTvuvDA6IDiCvehvXELCyiBw78VYZDUijPEJBKqLitJVts/dWPA1zmLroYsaZ
t6BnT1o8Y+/bY7DYVOfGiJEmUKYDo1hr3CHt5QQDI5T7njzKhV2xbblk3UHn5VVN
0UoA+6nUJmOISjapBq6qNkPYnLaRFyF+GHuyr9rnuNwdxhSKQRWhvCYVurWQ6kB1
5sSMMFYxdCFGQiiMI0TgtQoIgzT2iHl0GptVVqm/Mzt3O1x87XclIxHNBh5/cIrd
/61uxjYxGJjC4WBRe14i5poeWYeeaPzu2HIT+KIFFR38SLhOVHDAIQaNrNy5re47
aF8+tgo6KMVf4/RR0Gz+aPK19llD4qjvOk7zR4qIKWGmCQrVU5MfV1e0xoQ0a8hM
823yFonuwPnoWqZeDWeG68QWd1H9fha8geakOGx+kJ6PybBnS0a8jymc6dfQB2zS
yFoZxwCWDZfmmY/a4XjBWAMLOxYhSy9FKt9jvTXUdQFh15LTZj6fObcwUl8kOaxt
TSmbN+b1JtxPGqP9LeS2oFDB/eiEMYG8wluvJHBqJ42HehtMRgANWEAzjxJirbYY
5hmBF/CaIvQOVPYHJTYe3AxWnXLaIk4ekElrJKGqeFOiXd/ZjbH0uqV8Hix2et/X
AvmQLnoGa4C5gTrPhBX6BmwABmdXxRFujltiz3wi+M2PoWEkHHxxf/6wWIQ5WwDT
9KNgmae28yMC/er4udmpOqeU0NROTRg5e7fb5KyAgCNTeQevbZBON0D88zDXNAV+
kb7atHSGc4ko/SvFXV59MeMdOIKBxDbQHMfiUg1J5jayvgpKbc2cjlsAIt+69FnD
L2xyZl28BsbEpwSp3k0PucKuvrOEVu8SOI4d/Hqzz2jhRroWQTs0/LCvQH1gTqOd
vyPRCEm3vH7wedtarUkYateadNKVSchgvzDaPn4lHuGJYqam3GWUUy40lEa9thHl
8YINrzok8hO0Aig2DUMNLvZTfVTO9Y+iR5KueMCEGOxk5M8jLe6249ISr/WDNJQk
J9RCw8uW+pYueJKRs+sx01VmBmbGTZdIwenve4NKzm9Zf+wnNNcDwl309C6RV5rs
N7oxMk/m/WD25b93QysiY7r5HGTZcFguuFdDIv3K+Rd6CMRgdfH1U3KOuP/EPxMD
CclyUEtjtvd3FxiOn3Z0HoqedRvB3A6rOoadi7t2yHlMZZ+jpHd7iGQYZtREhU3S
TG4kxUy0WMchQoYExef6BPo4sst1H+1JvH7LPa71tp4ZVP6FhPW1ZVx7v8p6hPje
2iJrKie6wvarcG3o9U+LXXtHv9dGanHY8ntzQyKk1gRmyZVRoGUHZC/ZQ0efQ4jd
GxOf4rBPfoLHV1WIWPAAOxjKGqABYojTVvNXmWd5e9wlsAXVknDCfhxMdJBvRRtS
Bh6Y1yBkPkU4QI99iliokIlAtJnkDJQP5HAIGw71GdAAFRojnHkCbz7GyQ+Ek1t2
mNR+k9Ts8gyao8GeSq02+67bSKlBIejFSdDCZ27l99gw1nA9LY832Xit9qKChvGu
z7lV/69ZOMAfl6FtCAm5WsNtpayotXfls8WlPVbvo3KYLjERDTbkPma6GKRVVvAn
zjYRr1iRx/ZxbBFtKbyjWUAZqF0WqDSCVBQs0AylaudaSA2h14a5oQZot2FKhbY6
rBAsXXqHu89ETTVYH0SSr9hfr44lvdbPBBReD+WCpmW97C8k18N2kDXbexdX8hgM
Y7ycNZj7R0AhUqZLqkfcj3NFEaR6UQ3aaEEanKjrohPwHh+YcweTauy411sQwn23
Yeba1+akA3/3vXvE4LOzJ9TvvuQ7R8Aa71m5T3elSTlkTGXc2yewFAGPVFey8zxA
RKWV/9dExFBLCri+0RlRmd+KLsD4kTja8BBwxneQHE1DvCOYRgkWtnQXJ56x4SnH
W7h0BiKpmxo1aVQqToagPjqafabmPcpkBzwbpEe5pqPwLMX9ikGNFsBhSOD2K0n0
6DNY499tJUxRICrYY02ZK2Z29C9/65JqTf+SLUo/JcyB4fbJ3ib/dGtr8EXgI9BR
oQjWHuslNdbWLnpH3w1gTtbHNX3aCYZenG9psEPcfmGHbcsqLqBwfVWQrhJn0keg
aJk3gcokeJs7tvE7ZLHJ3Uk6de8kzjg7BPTznGq6oXstJ4A6HhVxn8MY4XvmGJSW
5xm06Xsa6fF1zg+9EztlcO/SqvuTXjCgbH9dCEMHFpILC5AeReEaT0Rcb3tnlgiy
D504xZiJCYZyFpQat0mgEB3Fho3QlNODc2/3mu4ZoHJOr2+4AyNC/G+0kbfMhQwN
BngJBvd00CL55vcJ+yfK5pF2iWmbNWxQmBHESY0dzHZF6SbNXkQHvPyAfQlYmiE1
pJKmrqeiYIENsehlHJycEWw4Z1cS1CJjsm5wcfGcKM2CxDbcRgxd+oqnzf9WoS7E
WStETsPrOAFgExRwbWvBaFSdGzxrawm4sXOG7rWZEuACeRIlNbXU7gjRK3N3KXdd
v/f2aZ0UzbFC/0tIcTcUJR+qLybEsWEyVFHNFpTvGylKWGv+62BHsv55uQbvAjum
P9ZMMqfFhcrIpN99LMI9GaDx/9E4cPBMwuZo8cSJQRWuL2alC+ZZ0ZgdSuuKAoXI
iv03SgnXRTA2KCgQxBTSwWSIkMp5YgLmne3eWBrIotfaUUoBAmwXwCE/klKhmNIc
bcVeRYt0bbdkFCRfNAnUNOn4zQPPOAL9Jt7SRlxbnHtWq2KKXjX0beiZta5/BBmu
hnp0rLecNVt7YXBGaG1k54Lm4qwbRAcMmW0XrpyCukscZyH/FzgOPFNDDVilLtTv
ophcEH3L0FG992qBy5BqnCS8SYKb6UqmxhMyXU5cVU8P1c5kvw9xYQcHdVQT+4er
iiGPusjf/c33qGvHFzFTPyXB5Huo+92sc/62tsT/b69QY4AsM6XMaiN61tSgl8qq
AQRVkRwL5NjihG6r3sRHKSzfhCn/d2G8gBF1tsKVVc0iBOBLNtLZnP9X8Tv+ljYt
soK3oaDOIzry9iJPirjWYd0oUaeKlaCymbHzcokDAjkQHfaFcSgRSH+3UFwjsTuZ
GvAMpPNQfvFkaXF/m8jVRvMCoWKC7zgviC8q07DrFxmYapur5y0+i4/o8f7OOn4C
ixKnp02ZbTMyaT0zGiCRGhxYnjNZnhhGzhGnZIbYMuw/WRTbM/aGiS+RU0F3giO6
EDNMrwOvfui8JLHZNvH4cimy4b6OsRLzpgFzJsPWPDZfBNXd2XPW1Ct6CZ6YWUKf
jo3RtKspCVuiFPwPEBxgxb7WdcgCCCFiIjj15Wfgk1BjiP47L2fyTomMWfsdZ3Ec
vnBvWz5M+QqbKFdl7ujTE7KniPASyW58xxC9XfME6oyrAgLDfYIsqdbn/ACGysuq
//XwyX5dQJBB0znFhUWhxPxZyF/0quyA4Cw/TAg1ZF9DKY2/nnJ4z0IPyFPJmpbG
taXBIdIHiWDI/xpJHPR0JH02OKP6dySvSUUDbcUPugXDJVcQpEySW4Y4+fnX02cU
f5rWqqsc1pgXM3SGJj8JVxAGGqbrq0N+mz+9xH6jB4u83S40RQuuZ8PM4DFzAZis
Qnu3dhiCfEqFPjOvJVffJxo/62RXIZQLwPEcmMY1RSar/1UoypZnjnuPml9lcPf8
E8SS8NWHbEaM+W9eBY2MEzkuNQLNJYcB6lrUS5VRWDKGwCuTk3w7cnj+o07yvpaw
P5VET6iw+qoo16DVbH4rWm6YbJHe/KeNSLEnqtmqyc9g6isqssPlvmAcuXpVZ7eb
PXfEUAJLuyI4/5XPQukniwKKHR+jqe38eEJsJbeedx45DVr/v5n451A4e4w7AcqW
/W63WeqjIUOIvqdHTpf1AEhC6xl73ygvSfbTbdc/SMU2mwb2qZ7MKJe/zt9Mpl2E
rRZaZ3qalwEdr2ZCAg3yguynxufjowTtcRyc7eyRCHQCCc1+VCoGXgI3Ep8TTjib
FZRPrQ3kCHGiX6RLt/DwuozVyxlciKYe/Ajrlw3XAz5YEjVrVcEVeGdmEAPBKfwV
xSpeCs7ETG1joWP5TLcklS4rf5MAo2vWflP89xLs6B9yGUeNBOVSyyTFnIOk/UUx
GdJd2OLNWKIemV9dgwelaPcCI/pQVDfZqwBSkBjaXvp6zrfr/fPQqd9fgv5hh/pe
qVid6mhPzzbB6L/gNz4krAr+dTCxHC3MSTEDEeWA49/ZduH9j+qWiLyBmeRd/PKd
XxTE/LRBwUi5UotdIR0q7DnS2KvIYBRcLEQFSTAq1I3Aknqt81dRfNVC3pyx+d74
nnyNxATsRdOxsGnSSpbkswKNefdPYxUdx/9hxiiMQsT88bw8t98swVguE68rb+17
u/Sw9lgUtai1U0/95ews1mZ5Fn3rL//7iRahQ+RVZlu8Gpb/Fl3etl/DuWcMoaIt
sZNPosWdXuiyFnjZhdiGM4mhhR4s0yxLwJtKj+hgta7Z03WP/toZ3ci3oK5h1K76
QY/KR30agTVPq9ol1bcAiqSKXVr2f2/hBgqVigDPdDZSjZZHC30nEbzBrhXU3UK6
Sih7HGcqT6s62dFXRoyczK5sirrxs6/UqhimYisXwSwBJyNj/RDuJSo79NFocqRC
dQ3uZ9IYCccl7udHaE0eYsN4iKqgrUt8f86+f76ZLOerE1tBhn9Ojd5FlrHPg1cB
HS2uXiGViy1ZxQIgMjhvUQFXqdW8Z4KCvsCRQ+rfh394J3P76bPdQ2F7BQrPzL6i
iwbNJRR4LzwZAFZBeCZZ7ZuedZuV+1cEkJ61kBjCByS30FxEHhPOVoVTNWbGXCzD
tq9ph86a6MoZIa3fCe4g7ncHQBM7zv3fts7wbL4RNmzDvs4C2krCaABH3eoPTeYJ
9sRFya4GYNkYN0IVM8A8hAoY+Vl+MZc9HxpAIDaTeBO4NHI/y55EZZ6OEcY7itvq
J6LBIp52VEwsyZxjNXXBsiS3qrgPsHkpuiDzSQyvcaPZOvKvjL8tmuAJmy6y8Owv
kIOM2hlaYdo2bXo+hQPCCKh/NGRQEqH4V1OPFhMfayzZWc7Q25GA4Ed3EbsqTBOr
qOcDn0hmVl/YepGzk01X5vVC2xRQ3IzN9bAoLV59SzX9rp9lIp23HTwNzdPgWbUJ
rxda1HKOo3RN1ZHARH+dywYjAy/uR6/EFi4wfhKEJAc38H+Q6ISR/4Hpv0jAngFu
7fQU/v/TkquaKc62lXdCEGJr18h5zlzZdH2eN7IUmvf79nm58rmjieNpcZmAV7p0
+dQUwq5AbftqlagmhGy+WomQfUrhna/26e6KbzwLqpNc+SzVfSZt/wHsJ5wQTb7a
r+cdEmCLqFd0+JhNh4LWR1Yu7ApL2i1d4H+8VQUGSjxRm1wrKAYzla2LYvsiM+Iy
N+OG2+AaKScnkCQUFpAcwRNHQ/BUQT/1xd6eAUDTY9yctD4tZ4ve36QNE4MBIj+f
2O8XlG2qdHeLfQ5cm9SihyBjaBhaaVJJ9Tfzbf/qxfWTrTYOPUgM7Bax7869STrS
f8OConxHcnwHlDvIzn8RTAamYBYjiuxUmL8Nxnl/48aeCRU2Wd7XfK2+/8WY3pss
b4bv05YxshPV8UpywLSJQXzuZdcGYCXAGtJgqdCUHZjQor1/TQocEC81+jGt0S5l
VKMm7L20Hz47SxRSWOQuPp5qqduYCwwvheLziTgjctJLZvUT8mHrJ9zQrhViSxBg
iEQTSf91sIjGaDSUjbegXmTaIvVYZMCyVUkxOMkJR6O//Wg+Li+r0aITx3A7EvtI
bkDPqIllaBqNTLIqUt2TmYCAVQTcel4K/KUy7mmcO9HO0J2Tc2ObyelCqMOnPPgx
OnpZu9vXK0PZvNGSyGMSGRtpSIPg2dT9gLVqWO6rilmu7CbKE/AELP+hVwTVLuG6
XbwNbLsxAlwvoATvSgvcrFo9NwO6rTWlW4X+GZWleBj3KYL7pJ8rcc99pvV/PmQp
NCtPgU3QCrlX9MfpjHIeYtGrlrayELFqf5LrTENmwc11WmadEjOVlmvhFzpHG+n+
p0B9WdZiR2jgMYarW40GHlVlN2Xjt6HiWqKa/CTuoYdb78UsBS6+mxJbpm4FL8kb
3bynfSUiimM+8C/Chpv6n+o57W7ThZ3jHVRDhRVbwbAXoRyQZipg0rfcyiOc08U2
d9MQjI7DAeIcPs/sZ8YtjrJjDuzeLYsVE1ChcP76CmYdHw6alhK1syweAPgjMAMq
gXreuCvDsj3BeTOlPfs5lL2xth28tb8OPjUMz9LMBEHbzcUkhTW1eTmlhRN2cpj3
wwenJ7tx3WPYoWZgv0U/aDbt/0VlcGgd1XzXYcqwBeY0vZ7Epai6Zc3j/el6Xig8
3sDBm/soW7hWCzERykUT3R58pfZzAg33HuPw6sws5DjPJoSo3cb1HKNaK4Y0R5qC
mL9vMFvM3ozXZFk2FzpGgh14WX0M7bToz2W1hFah8jU97jIqHawVhJtB2vjGXxxo
nHutxJND1+dOC+Dy6bfe7BgP7WqdkpTp5+sXsEmdB08ybAUVhsLMN04Dx0Q0Cs+X
gDstvP26UWiNUaCZaE+qhe4Ds0ZflDkUMe0s+EakR0KOhbEIkNslQn4z96gqB1w6
7A8PL/0C3Kg1jA9rNJuvl7QfBi6RLnhnpB16TBB4yavGzwPvXFDMh+Aso6cnkoOy
2AXFUw7Gn1nupgtoxclX/Sd5+rBCNNie/A1JPZDhfwSlKOSOZ8sJockrAHRXZnys
JNvlmSAN1CM2lxS/yDC52yADWq9MuBlYAmXiLLhQZZkv9wJ0Wpchx96YsxZ7tP8K
N8MgRg6loDll4TEgUywY+XgEJd2mzYu4tIGPjwtJN26cJ4LSCYW81KNMxp+npodv
yJ1z147xym56covC29NxaJ7LDYxZB9UUK8nUKp9Q+ms4EnBojsp72Q1qD317en4b
MN3lCKteBfxTqtZSVdDf9nD2amW3v+vOZdSAZxfIW4VXHB9moSlAv7GITNz4WFLQ
o9oOjONT+qjW6KNNdJWd19nfwBBCN1B5100AQxQ8bJzS3LMcgZ14vz8AALEhRS68
JJQoVXFTGMhNbUSjyt4wPYNljrwaSoEXqa9ksQqcpuoh7QuKQf8+Bj1sOEPeXuLA
23fhN3ST/yh9oCheAOkYRKillkKAUFTaxf/4d8Ms8ogDGIzD+PlbJ7ZQby6kurp6
jusAQ9q2VdGbskLvSxLl9iMW8Yh9ubWoqPOEUrYAAs2UvhfRD/zDByK0tI9l0CK7
6QGtaDu3x6bEFIY6Td3xTxSvATmzRFYpvMkW8nJrUOGajiCpyaTjOUS73yBvKpiE
vy1LgEM4UNQMYwW/dmKFIROARQhrxEXHlSAY+bJaBEnFdtnmS5hlL1Qk9kfnetxI
1dXy735ttaZVDzqUEqylEA0uRrjx8FRpc4fKPP+/WC0NmxMoY+PYkn53CnyK3SIE
Tv8N4Tzqrq0/2OGawLVrMByEnaDWoFkx4F7RgSAbG01tPlUQ0zMwRyvP+MmeO34b
ulwEKMrum/Mw/780PnOd9kxnk8DSeEX3tfLCltmp7H6H6fS+C2dld/NKnwv3NIQ/
4U6AxLenJnvoNbkFgcXp3hoeK3EdNko6+pKVrAO8y7Y7LBndaJp3l7vsTcQRoTFm
g4xY1U0xYoq3Y8WNfSqPZlkPK+teMHDeWJXpSCHtTe4PjwilyZmA6oRdUo1l8i/k
2AchfBgdijmIOh0LDsFVqFB3kZPH/Sd6Ye2gBT3lmrmyDecankhzkkraG8qN/UWh
MdiotiGnCR9PKt8GTXZ5Y8hD6EJC6N5/x8NqAmVWcsXOy/XntxSrsGn/9fGnVmXn
CLqP1WFIB4yDOTK753pF0gmj85DLMa+QTInWN31XkYOK/ZIGb69rnA+VetXRShFh
wSBTL6tmeo5M23f7mG4q+cxKdl7OmZN6diJCroweqAuVvde5ybExEMq+U91B1oMw
Poamp8Qas+ofdnx6b2r8p1iZjQj84ujX963GiXVPbSbIq54qRzR717aVu6o+7GRl
/b2SyQMXL/XjU/4+E1KpDD5Z0dvHPC/oi7t3tp3Kwx/4ax03vm/y1ExH72uadi1T
m6F0RHgY22L6AfZtmlGqA+ubjELoaxfVrnpnpQwBykK7JXmPRdPLgtE81Lo0ZsxQ
1I1Aiy+x1zJ1qJDK8vtyZl4uGGXFLIUcUW3g39P8YaiwYvDz6EnkWEa0r+ASa2SZ
Ykn738vyP2KCTPEJzYP2EX1ga39ap5zaHv8Z4FVDWlM8AWWyqkaW+zYDdUWMtumz
IZGb7YGvpM8PuB93uoRhf1KZXgUVD8VA22oiSivtchoSG0xBB8coiHNTgCSUbggm
iJCrryR+tUzigmM1CFP+ZsyuwwuNfaXJjRA+gUT99o4RdDo75AOn2M3YmiJ7ZH4g
qFNawvw5LETNNUHuQSkb1DKTVeE0iXz9Q/cDPTgE/p2kcfpX9ckCLZ/xXRkFl3m0
cYJEfdycaWoHdDU2Jj2o6JblcfLCXXvDoE981HvoGr+OYX53Vg/vf2X8LRDYgxD3
prqeCmIZb6VMnkUYZsSEPkdAQYMtFK4YhWGsvJ6OqlsF+Q4ASMycjVrGpsK/qo7I
PWFWOKRfVJE9CV3k7aLPxvanxDiu98Q89Xg9MNOKZ/KauSmVdjbD5mA8hcsuzCO2
Ozv0xAThFKKG1cGIREy3laQZ9exqN7oKhTUG8a1zy/zpt/kXSr7UgMn+rtS+XEfR
Iy4vmuFNCKV3TJdpCTV3CHf0WCakf3+c0mCuDMrxaIFv/fVb82Y80U+Zsar7fpsG
X/dnIIcm9tyaUjPg9uhaGqKWpdfN6/FdfQugdy78YgeDgdblOxQatqgoYZcg6AVT
b7VvZTasJAufiHhLduDS7sftsS//yKomg6ucEo0blbyB4mzbKBfJfBzeSUf5uGCa
6JwTcxwYk8YcZOdEpJ7aMm+QD3ZPD5hf60sSnE//yh5pPlydP8fU0qPebV8e+RKy
+hIb/L4j6pXf6Vi5SYgfZXPuW1i8oH0hygwda/8pEJoUV0VrLhFfOBVYIb1bh+8f
on/3bef9rE6S9Jn0DwZQc/4teNJ/4YZb9o683YfNqSxk6uMYk7QI4AiD1HJH+GND
GdyB9RMxzjF5stVoYyeQMH2E2VEVDSJpVWY2j0bs51IxvpIMIpRKeIfZKFAHA+8f
8IsgcnUg1VaujH45qJhLTbPf8o+8vFAg9QdMSDKdZewfunDFBbm8c1pgC7RRoKRN
+5mp1VuhiNe8DvNnBpOl3qF2f81lAiUXGLJBzkqgF9S9n44OvOZiEsG93bachkr7
HhudnASyMaLlc52ZPPEmIbAUFB/T1IuvxpBeT6vsX0ZMouX9jREolZGe1YLMmIgg
2J423v9Uc+g5XS3jg7QwOrzELtubzsaKtW4QjoWtDJVRH0RhL7oOhAcdIrNKHHYZ
P+lezzvISyQOdL9gM9QsQ9tYA/+AP4okI+riTB49VaV6ZroJNPBXugOOVQg/c7r1
wBctXM5DCZdBU3gECgFS3e/UDm+GUVfkcZ2I3fVV7X9E7Hpwv6eghMQYmPboGVON
vObECKTuRccnxLsnULRDCqKk5BJQqRSHP2+HWxT+shMI2tQRY7Q6zDBw5l1LySSk
quqXwXS6fqxM43x+lKr7cua1IGIXh9QFUMIoAS7toVoybY81K+tliiItgTpkawX1
I5jB8XGgZ9XM1VflxTro6hldllJhJJkrOFgL/zHGHtykzQnWclHtKb6We2Qpkiea
mC6WH/F/TYCGaaP7Xyr1ZSG4Xev88KEA9t1HhEmvUyV7FgKKq8o7nDnrF0R+ndmY
kYrZlaeJrYdfLlzTXsBDBqX8u3TT1OBf/FeEMYW1KLVILWK3mFHyyNtstNmvL6s/
ICKxoq5VsURyJlTqd6P3LCsiAvp0YdwqS2Md/9j2AS6kPNyddkIOSX8NlwwVzknP
zEvkHr5UQI6aXdqvV2Wxvve3xZ5j43vPbkZip2f9uhzz1jxv6UXfWIETMsDQJ2Ew
IVk1f8g/67t2ZeFyuNgoR4DN0GA9DxweCTQSbJe4+YL0eWYIdKzmCAhog6gnPtsu
reXCofJdpyAj3BXfgda4fUjfkgDBgcnVgX/gdLbmA809GImrtkdQ4cnocJnT7617
QGMbGHum3WVYq4uJWgPSdr0HbtcyNH0Pm4ZC3/SbhcdM+NZg6YDkv8NsKO3vr+BJ
7dWdgJUCbA4Fj19tJEh3PUJGY2HTte8it/VvJOs9CyvMKgKRlaLOMccOus6MienH
LM1GXQRgI/SYPx+JCT7TvQFj/7hs6pxtVHpc0cejk4AnTPilB0A259N1qOxKTAmP
G2GcNog8A8ywo2bnDbCiznU0j+QVcSuNzs2RIRUfo4ZkGx6XFrf3GeBuqdfeEmTS
U9HKC8bOUxsKGuCTxuB/6+f2kZrtZqpvW53mLFYyfesbrJZcCQDTU6WOnhtDQ1dn
fwLNT/t5P6ER8/zTYSwAcsaKGhZJXuSrlNJ3Cb55nsa9g1DAI4ZSHHxW9tOV21qp
/t3Q2uc3RF/t427+ucwE20svjb9d9Y6eDs/z/hrLFP5ES57Ee8CxcnqKH3oRP1xS
onN6lIMZ7xsVPevCBek2i9ZVdU0bWx3i/kQF4wgyC22i2dk7X0syd0Aaa4vcY0Qo
QYGFfqOudO5kYDuysrS2Vs30j54NLtD6W47bfGbKMVgewEEFWYPzLmlGnT31E6ej
QSTh5sMMmllwUnu/BjMt5QfsQJSWROVC75IyfiXYl/L69xFTCuWw371z5p88vdp4
6tQJauZ3llpUAo02XuvTTBC52JmJjXUqtdCp5v/7l8oSfatVHzXVIrf+JFgkCSNN
0wvyK7C3Cl1K35ZPkIrCpnDX7logJN+LCCEERygcM3IIGR0Ut8CXPoApQLmd5ckp
byfLS/Ez1OGzSRxaGIKhEVzWi7+uH9IE1Ri45RYKIzaa4x2TyRAwE1I9oPvDaEHn
8Eh4w/KWChBnmnJhIR72NRTeYqSRwkD3SWo6vBynk/eCNtMQ+X41Z2NC6lrKFHlr
Ci3wycq7PjEY8I7uVGpGQv33UIq4jGs55XsEgv++yncYgHvDJaVJipol8VS45sBb
7yFWso07V8gSfuLPw7GR/tWA7k6hJwIxJQJ+Ui/wNmLCTTiPjCCY35bNSHmpuMVX
GYl/HT0nXYWtVqLxbegjEsfuZd0WMShMtF4PadJZxkovYS9NEfcTYuAVShbYzqXy
hNlP3V62EylVInb+lOD3nlRxJksJG9BHNL1GMtB0+raWtKXIgQI4mlgDBMIfTXF8
CREeQOdmWaRWYHEzVew9NrottZSNrlBpJ1laKE8A9W36VBugoNPrVizX1TY22Mou
/PN5IQCqkrOMS0ShM42/UPBwjiocuukI2K9L0npPnidATLogcjv9Zo+db32rVPY+
wXOVXyWM48UeOVZdpFOBPeetVYRQJsK9aPqytDQJeRaDVsqa3FrEI58i+hsSgiOL
LqIC5y5jytEMAvmci7Kxhj9HFVL8QhMvdRV1CYgIVUC6gmLBSqINsqc/e8P8vdG1
o84Ki4RrUhG1j40QcvbN0tJRX/XzFQHBAyZLtNIsb6802ogAExtoeHUqPI/H62h5
z9sIwWYf9JOA1+VBYYgqoWllF94PDYpJXW931svkIE70NWiehZb6NEXh4ySP5Pxl
Aa6/1n81SV2WBs3DUEBYmMpmVpU4eIpO8ycui/uH4uQVh5h/R1ZjalfMo3GAJ+J+
UPVCDcObLRgGFwZWDw1BAb6AxwTtNg+scIIKCJB5hWKAfMr7YE1Ow3X18Duli6Ey
AvhVn8CFvwQBPBM6uQshA6HFEmNN+hJGtsb0H0FLR9JJ23SATCXXC3SW9Od4Y2ho
EZuk7shOzhlc7GUSGVgovsq7ZyrVfbnfg2SWBzubN0IVXxS9bt1FCUXLcfugkW5n
j65J+0f0ukaXIvl/+JUY1+NAHFG0pzMPFq2jePahhFSJlNC4bfgLR3Qve0cPjqHA
7H+zohIjRl8zmRaEFEObOSIMx2Cb1ZdlBwOaZy4v1QeWvIDzyA1SndkDbC0rTdUN
383xTlZOxs7/HmKyD8uQESLlZngvCQ3/BwI+ntsrf+L3SCox7dO8zMT2BCKd67l/
1XFaonL1M5i0a9qWGYe5v6MLQy6KnWpe7D/Mv67cVTWM/Lwf+crezHTDeiYBwhvi
wfiauxJUHjC2zDFJNz8upai+lFTt8Yb8TmVDpR6VkPigLvO+mRgyy0P2sUKHc5Sl
NDI/nyN2feg3/T8koqkK+nmevIhSeoCilCybwQnOjenKPIezlersnsZMA3lUbfQS
p52ppgnCl8BMvSBAs9QxV/RCH1DK4Jcc39WiD0Bfq4xCgxtbbG+QhLEBezKLnL/L
PcAmqLZEd5JekyiGN5WG5gplP9+jQi8Eh974yDl2D9DRaRLGRU6mo3pzDCsgXxwy
zZVg+L5hwAKDc81yrGoIOkhgnGOF0/tSrcHMybCONtxdlZpoDYjii9EhqlLeY+FK
96zZU5xvQwO8cSFbsQ955xkacvb7iK4FxHjgAyHO0OoRUamZcACthSRf91H3DmC9
sjPaQspyMLtPG9FivWwVP216r8aDN0tujCx5/Qhn4EJK4ZibysoADBlytyiBh0+C
F/AdJMLtaWQJ16Q21xyYYxDgMS3WbZln1913IpRvurB49UcKQnSAuHAy4aM19aOp
vfBleOVqAmW/iXJ8UoWaaN/vafWooGckKl3pmFIrI+ZT+XfzDATYwqBqJlDFKgbT
1GfSQM0zP0b36njtvZ9Y3nbxWVB4lYs09cccm6/cdfbCRiToachiickPAGWkhsgj
xP+/n92U/tgeq672tsGcRYs5CRUMU7CFH3NiTIVMb/UfhzTObI57kJc35YijfRHb
lfCWUyBey2OHrSjjDCsEgb9Ng8b7meZjRL5vIuXDoS+LWWKqhwwTCocQsiPTjaMS
8t/YaPMAg+9/7pVEPZw9EfyVzodz/qbXMPTMWtttav104HALEr4vIWJy3CCyvw5R
FsPX4W8W/RVtp6+WMOWWEe+9tAORMi49zD9PG709QREZu0ueLXvSx3S8Va0iEMeF
mV+Mkr3G04Y+6hcnwvwOKfixev7r4wAFoHGHFh7B2306q6PraEfxoxcH8kE9sKq5
PlG0j9DKJbUFJo7JEyFMOVSUHZIis1ikAWlXoV6h54zR6jnPk9LUbYf5GFjuLVbJ
dtjtmUz5BTQpMzbhRMt3xDBfZL+pnItmxptgFDBGJUPVM1ls9ehufVJpoVjBV8DE
3Z+t4fWD5B4cq7cqtzlFstiVn4Wc4bd4Yhl1SwUd77WzjLyqtbk1iapzebT9GeXC
nxmFKnlK8QE0Uw+BSS0ocUvpAYeTRkr9iDIG4kgqsdwNr6fobo5m8rNYV8M0SKG1
qArtVn2Fjpb8TF4sitqWYc/1LgJBD6KI3zU07Ts0AJiC19yHAh3te3sJQuBXu7le
ONh6GKA9FWOdHGzjezpT7KTzKdR4tgnfyTHJoBzuP/OHyEPzRLrdXH3cUeS++2e5
nme77NgDC8JyIAespx09YnLXij80NnWJsoxQ2IjBIhQO4+d9fQKKS5TA830KOmTd
7cRaOl13LXTHCJOdHEjgbJXBvmZrKP4VJrldzu++InNWXcOwpNqUUHaoqXrVWOq0
14Atzilre2U3ksqRbX7BZdZ8ystAQpLqJG1cewN0psaxsYI1O2F3eI85t+7loOuV
mbp3G8xYlXxU9coLk2Qia+kSaVNaJ++F4yV6Gk46PUdis0/eFt0vN/r1YPV4dl3I
0T7NY58V3yiE1/Zgm/Pf0mEpHBNnTmqeOUdjbS5tIbey1ZnTHHrULh36u0iFV9jq
ZR8AYqQYpTZj5kZ3BzhE9vrKHEMw3+09fm7Ofg8/4aQpDIHjH4ar6GRaZm3+PNa4
EviZrrwvGefS6bYK48CumKtgKq2PCtnnAbv/Nx1gbihbWwyAg7BSJDkeOc4X4M9j
ndWh8FagjgUOe2wGyBNoadyvcXlEuD3eg208d2hcvU5nF6QpLOtBItG6+I/j5aQ7
pDuB923dqpw3EM8oHQKR4h0+9LGNC6rhVI9pMwSKfj+Sm4i/P5OoFML3o7anMy6d
RzZRJE0c+OyGgcprUTs5+o3Xugd554sY3aMNN+3ugKZeS1DP2qEtfmOiAB9aZ7n5
wV/3uuSodx6ERPGVMPYeo47CJNdyLAYy78Vykb98FsrM9oQ7g19av37k0psE2PHU
hKrbOZ08xXJspniync4QLs7ypfMTN9zn/fB0uqzmiz4vZMgs7RsVfiUnZGvFpjKa
dYOdrIn29XuSjqP7cB9OxYsv+iVG2yrUudMohsfpgLxqdnlS9oNpEeX1+hqGdcOL
EIfBYhFGkvxCGlD9eueVkCWekNxD6cYRTiHNYvyYXgs4w5oSOShstubPY9LnlWhX
nxPIaU3xQIE+lXdgEJM29ubTc838dog8lN3KyOUFi7Pq1QexjwwBEiUnogPaIHZu
2Y49VT7Oi5DGRQSSnNVMMSdpiZ/9ciSCKSdpwlqvtAP4u1J/et3SieTJ6aZd1CR9
+ISBEM2ECQT/egHEwUXjAjmMtIo/Lc8kKSBipMTO95xfzh0EbjSOzHirPYh0UmIc
z9dd8zXgZ4ZaKYJB/aM8okfgqjcPHmfdqtgwiqTeNkOAyZInYzceTtzGuBw4P7ZF
u0qWM8zAC4M8YlNh4twzyDdI5IbXTndhOZCSSocqZIMYbdByc5OmAGScSbB1bxgz
hjsvHOrli2GMKBY5uJeV+P+aaP/jw5GZVY9/zl+52pb1ZiigVtMPK65QxGhztiYK
P4L1PEteiW1VK4hZuXTlDO6J2tvKtsNSBJdLr/plw7XAZzlVxm9+aNzZ3bDouZ7s
JdgWaof3UOCLeA/VXtara0//KZ/HZ3ijqMhS+hodHblxclKi6MxPOk52gMJ8nENb
17R4ZunKgz7bIYUlvuFwcrsGXgV8r8H/g9dE1AXzxd7P26lzc/4yV/uwUIonQ0y7
F7cPOsOSwgGdFNjl4yFTnzWqB30w5JwLLbKKRKsYwM2M0isKgjKW/+ug53s+t8ft
p50W93iGP9TsLbOabAztpGaglkaWtbYkYWYaW8ZOSUJKCnzIer8Zgph4q80w5KkL
yVqi8PtIEleY18uZDsNCypQGiNvjZS1LNlwHsLfVBERr7RaCcSs0Ua3Pfto57nFY
wx93aOpAqeKanadAR311O+9HznH0+FyDretSJwXVlKzm5qNHWEwjj5RlrMFoW5kn
RNoZ8GoyKUeL5ljK7/xhsZ4nPGQ1tHfoR9DNv3OarhubLk4P7iQSmoQLmDkmUWrh
YD/MQF1Qp5maJ+HMxBPp7EYGAxftMjg9Y0lU6uwZ9tCg38+24Q5p5dZ/vA0Pfa7E
gyxKMqUC1k7CdKxjj5qzC7w5H2ogN8sfl/rxCjbLGWjhJ3RLkcOOKYy12IRRpec0
js8jcMTHlF2sBUr8LhQmfju/oIGi4X5mj8V+Cpvo0w60dHNe24G4EFn3rNzvzxVP
LH6goE22SXosCSUNFnUGswHz2LcCF5jTL3I3U6+sVRX4BPJwWeTuaZwrXli15cyz
iYzpHb3XTCAxXSG4u4bIVoHP0etXrrGE7lXSkb+JsYM+vinOaMI60fkE2LgBZkTt
NPcPHnyuIrPGtYvM22UnvbqLRSHUx+X/f9gnnm0uuFeRV8w11K3rSrkV9CtKb+Bi
s6c1eq5Aw8l1gDtn/Ofj3SGe7UYfDVRrNj6knC7cZAXFVhSX5s+8tEqsQtHPSPNV
ddJNhHtfVhm4TyzYMdNJDVeQp3jK8VfeYm8ec5kJ+0qRVfSxDTlrwZv4nKOA1yIL
H85ZG0Ek32u0vQX/nTnae2qQv9Aa0eAYWadHox62RqO9Ku0A1MHLvtIKke1Z+Izc
TXkUAywEzgT0w81fW8H66cY4RRtHbdMXkoiAU7YRsGgBQ/vQ836rMwMRuQXyoc5x
SxW1ELfyp621ElJOPEXL/Sx1ZuEgEpj/Vwc5H2CKFa69TsdGb+le8F83qDGrx/1z
9Po2O1dbXc2ozdA4PS/ny4ZeJE4fi3NR/ed1UsSe/ceeXOUXrU+XiAQrcGUYUM5O
UDRtr1TuJTXWyQNKNzqnjCQPaeuAAi1Shne3HZsJlLIafCnEz/dsrsEdawQUNB4c
44Fc8YJw3bmVzNd+61kzIMkzkm+pyFnW33562CRUZyGrttPdAX2xf8x8XeD1VUUx
hIJIgOlpWHztAx5cHq3YXTf34UZu5CqB2pdkGlrlmBHXQJxJU0c/68O+ZZti5fKN
GZly8PAbhpm4+PWC8QR9fOLBkFtUFqt8M/9bEf5RWsr0JxU19Ds6UCZ5CbauRR4Q
DzhTtaVBK4mAbI/Azer9Xp2lCBKUnX+I5qEqEFuMuYHVogdR8MX/Wf+vZsWRjgy9
09tQa4o4cTdYjrrh5UQ2wF12B2+arNOMt9SajiAfbirjIXLXxVF6te/PW0s7MYxe
qOe3ca6ZA8Htxq+DM7VdhcpP7P7dV4s8tV6ab61JSurjRSup/oTyusjfucF8S6kB
7etTUInVQEHpv5AuxO8/Xdi3mU6eDqFO4UxSA6I5cM7evjXgE4l/LBG+f5ve1CwT
lmLH0sEw37rZ1qCNuwG2+wpmSt2czgtipNe8JbW2v5xn7AjFKnUZxSwgPRNhyQa+
etUahDjW4/FtwRdm4Vn0dPs8ZQc70QeomgpKU7kF/y+pwgwrMA7/ItJtE7T78vw9
irYsT7beHJVouZ/nKl6XG+7Lik78bhYQxaIfQg3UIvourxpm0E70bLfembklolHY
l7Mj9kF0/O0Jon2OqdwZdf0RF2vzn98aeKAQWvI3BcL9SPy+ZMPaVO6EIXHFZOcN
9PO1KtS3uD73TBMN8uz29c5KsbP87OmOq2kOTr3fkwTC3pwsVqry0cmwFHz9sODE
DfCRO53DBXCzFr1azizQIYEa/M190AA/D+2nASPayTimEry3S4KssXgzOUcYBfno
EXGwpHZbHXNdlGsZD6JuXNYNES1B8VYvW4yyFtl8JnwKhG+1kmRVHFI/Iooi6j1p
Y8EYsaCcfkTnorR5KomZUatZ0MeJotrTBFq7rw3xz1RgKXaboMpd4+q3Y6wVjspu
rNHs/TrnGmSqhV907ZdpkxpqkDzxErveKw7mhOuu8RFKxHPFpJAAEwdANC6OXNRe
A26q8DZsadYM/N6JelZq2CVuBBSSzlPbshajL3jSLvr8n2t0cyDzG04zYVH/V/+o
lCnz1/IiPXnM8egVqlD88WwopQi0osWitoFkO55skFOnKV7jIfhw1IXt7AZpMyDc
o7MZlx9n6HFopLKZLBDHrDdbCcVbHEFVLJn3eBn1xBTMzKk8dD0w0A6s/vjk5Zcw
D3cByDixo260W24YcfYGdtcSomuOrmk0DvFQl2ofcsbnC30sb/zIAe3N17/e/PvX
+HrE2lfbp38OgfcRQ8Cpb0b1Z9ExIZkBML2ARh8xcWeg4xie2TilISqZW5GbE+Dq
HjdBp/vmosy9wdTGntY6t/Mvf7FGuZxeJhjAC9iV7tG/tynd2mdIGarXYomiZ0KX
NDjFIMhYTzJ6qzz6sLJYE/hxfeVrgILe0UTleAftGAP0hL074w1PaFZeSBWaN3Hb
BdsMjno3luWcUMfAVXFaCkEMVDaIZyYkSNdK0Zr3xwl5maad4JcTutIUAQlXAMah
LnhHRSa0yRHff7vrP+M52kFn82k4VeDPZ0+A61eSfGI7vKceT/g4upnQxqELlVAc
wAAuwyn9Y2tGesP/LrW7Q1FDnudnimW3fahzKembpYqi/T2isDpekYMDwKvj8z71
13h2Z5DyQ1FDjssryJVW+5r09Qv8R18ccSSXr+CVDxZnmGYyM2byYtfJ9pVlOLNU
i1kREe2PkrCkQt01/bXvz2E9zYUyZAwUH+C9OohY9isnfhbn40G/6yA7rmWwyi7e
4ahSfC2WfN+PsqUUaZXyks9XMmT4+g5DqlIwQCCkfao6OXg7AyX0uJHHOuB7csUd
X6mf3AsGhZwXLiw8FophU3ovEYcQkMxJrj6HK8fXKJg8TAfW5mraVSFZTMGSCZSw
2Yxnd0TK18bi9zGoSsPjIJmdHmV1XT0wrFhvtI5hNGlp9ur/pbA3Oa7NduGz4evC
h/ugmT8HUhheKNB4nu2539s8EhhO+0nKQqgiOVhJy7BifXOV7ij3a3Vs2I3y3nd8
lMQU3B6iBnB6rP0mX5S4d5hCpdARbV/AL/KE088DiWosGgmxChC6auM4WKjrMeQI
JZR6vLLxUHq1kpvEs5Y/WigV8JnDJjAaZ/bf67/v2yMYJ+wgfP5pMoYlfQKsYqav
loF5ax65LMYrpIOIgweHI0zVTVAXkOvn0qJnT1TzR5qztCzlrADgrPtXmDtawkI2
j3SzVgCgxVX05/7Th20+XzZLEE0fvL6hCBOZljxBTqRTyUiO8vWzsG/fcuHEoyGf
qvubNaGz0ANFquBwygON9b0ltS61Dz04mta3iZlIptPedzbtSdulredl4ZpM4w1d
P2MPtu6SWYuyEIA5SD24mIX97vANUUCbK+9HqQVc9SqQmdAskHflK0ywFT2zCd8c
2AsslSjWYCjgvHYuXOAL/KGCc/s3j/bR3drDsX62r81UwKLJcT1UHmG6KXLNECom
3quk/gav3Eitj1Z+Vt3iQBi3l6dMMFo/hlrkv5bCMPRnxEBmVTyFonbZh5mW7Oxm
GR6OuuXJzPHl2En73kzwKqj7gN20fB5/EXJ7ikRs63PzcPFXKkRVMwzkhQSItZhN
g+kz0LW7FOkIUYOIFa52+31S0o4pXP805ABx0G3EliTT2Qz+ttXAmMqHCllu9Si/
RmKRepv8V3cpUayxvtc2vTVtj4+G8Rht1njUf4P2XUngBoK4pTyoRFYolqSL5QTd
WO6Qk5MExVLkQE1w8Vxy9MOTyd9+KchPYzWs85PYz0c7waMinnKnJguwO2Pc6FCF
tHVArKa/qwWxWNJLdYzYcYm9XlBCUC/sBEmQRIMZhCeMBXunRO/ZbPe7O+wGTZrg
9vkAd0+a+667Kw/xbXEaJuPuSd9AuI4IFGonRfjCyUkgThhPibvOpkczVgoxyeS/
CNdaINuNmlJzTSShUPXrnOSdwJvmg9CK+rybRBme3l3IpJ709mT7IVJuOoMLoX1B
XB/2noVyvIURwZFJHLbPe4xjqsa4L1eRxO9QjuX8kVS4dVx/kYgaQqsTLDQy1QHl
MKNhTNlBN0GEvjiULus/zeZ/8Y5y6nGruCyLXJBIv0XDsvBFrdCx9S4a9/gJBd6P
HXszddyGVhSC2AOVTxQg/Hd/BpjDIqZtwDWjt0U8NWIOfCZuwcAoSsiJZK/0MkcQ
JBnHOURCn53+Fy3UeVm4ey0fnXWPmiRe1No9iAxY/0TGxQN8VhPr8xKi84A3buqt
76L8ujM95+Jf1jjlvNS8zQnCZh2vD1WNJPct6A0GQFt+ZPHuDaIz5YcfK2ANKXJ/
k4uazldK7zb2AYEioynLHq9Wh2tVvVWEttIUK3B+HHGlM0KNmY/699Zs82E3JLo0
7rWIKgYdxlzG4bjrGpuSLLPFKKpbKHRdc5reYQhbSMf9d2mhw1AFcTek8F7z7E7L
thMt8BTW1IO/+yFXNuxZOA/jlEvl3wD8QZrzgMiV+bQTk6Q3l+XAoc9yZ+d1w4w6
QpQxhXJDN/Q8uusUrdEOi8ds3wMrwk27XgAP20YY3TT4+GNN4yYgs8L5E10TkVDX
NKdWzV4UOyO5L8yWEJUVTB8qD2QItRZAquqhFy7JkD19dKSjLAXNz5GJBEa6KMIC
Jzow0YGYHUowaw1JYPNvoLMsSmbkezZ+dVIl5XOSJBixH3TFs1euMRIYrLpRhCTJ
nqOK4FpD7KOIO7q9OqwTyx/5COgJuMo/aGoYOVOCLo4bEEf/rlASNlPyGvj4Zs7r
3rz30fO/GDSEn7tMmV5hW5iC2hzNmHl7sKlhA6iXor9TdWF6UdWjepIf/hTD2Kh7
0U5ZFzKTr3XJQszSdCYbdtDLbqdA9Uss+tZMJaHX5NVfyh+D+uaO6AadR9kbn8aP
mHjb+pc+i1UlN4lrsZSDHkcwdQGAs0q+iFXbwKjhFMi9HZ+jw7Qm/KVUfcRfX3ZJ
SsOWBPwp5zXLrEslEDceYANcHjGa+vKTcF+eNjIrN6MKmo6A+b2UakG1LNZEyPkO
U55f+vh9JbnT3Yy8SZgbTPzngg8NqBSXMvIRrLKJ/huH0CgFflEPgYKzw7l2KXlN
JkeAFg8DVYxls5bjc8V6jJoXJVIsUxxuwAac3sFQ4il6XGfyt6FsVT7wpXUrcLn5
Rg09KllbPO/ySSEJpNHna/YZ6gEpdL0VCcCMBdWa9uyw7NaHMIZellVbFBbMFA1B
ezLZ0foBxChbSboJYaEaKog8tcwmUc2wrB1ZUbxCkiEUA+VJVr838hhZL/DUL3UX
wJIBO39E/JKSeRDtwrJSIpUqw3VaJS7UQa6Mb2ldGXTAplFmtXUTMBI2BFjrTJx4
jofjIAzhzNoXDrNIjt/GI43opfobkfx/bdWfmBVDwgz4G5sPniIerhF/+7vXCyBB
jVyld5bLiwkpZU3UJ93LEGYnJRvlIFnvFe7KhPpxSjpX/quNWMo/LSTX58ZM0/gF
A2CFoG85XcS3woFdwmq64wGN2TbWgKHZiGsxWu60ZiEj4tbJeqyP6QswdxXV5qq0
dosgDQ870HQ8gN8nUJr9dqraCSEXz51TaDxGZxZtuLhjavKgEYJxZl+LnwQGxtr5
iPRjYKB9/Wqy8TlfltL1kLLYfhWCK5EvZJtZtRHYVe/kZXJcGK5iZXeBOh2ORLSC
g91g65hHi/f1th31yb+ZtkW4kE4co2adi0iE5v5x/84cuFjsZlwR8zdkbeCTzLN9
TungYvpe6fVMMkjMULuQD9920eBW8GBBEKYNTkgxMmLvqyuXcIUZnA8Hcrr/EDjs
c3WtyRjup2VQgEdoqXUWZ4+vqOHKnXvxLYCKTo6LQ34hslJq7lildbrcmcnYgfn5
O4Yz85A7MQB44NcfIjC1h3Fsx8k3G2Vq1qo0Ve5xdP+7xCfT+pgZYBGgDXLxk4KN
9E+R+JXdu1j10OWMepxARlK/DiansCzOeZ9DmV/11pGGfTJxZmV9Z/iG6AdzLcPK
9qc/pH8rbsXKLX0sKH1YnY01/JpgVFIw9fcOhZn7iIVQd4c0/3zSBMpj2/Uh9kfF
YpJWx818q6MjjBJZlFSuudZhOBrMzSLL5zlbmwQ29vAe7g7LctKsn0jPGc7BzRSp
tyxbLOiT6iOBGuig0Vk1bp+V+xEBvCH1PeKO1fWCM2h92VDKury0itk7ugqx2ZbX
lhMYQljbrCTDa5CobW/awrrORBkr6reFiD1VgJDmCVU9Pss1qzhuCW6vWqTCaSZX
qkHVkHYzMshIoLp7oS4kfG7/raACXQVwUI/8vwUt3QNrc/2tfSJAbx1Z8pBPkUZA
L07cbtbr9CgkHXNUC7dONdNbpBdnD0ZBzT/YMAM3icgCvQqW0JsO88oztq+mZeqy
5ut5rIEGgGmGpq9WSnQcUfKf4JB0qBByqVZKegifRPgIuSQBl8E+agtP1Q2qzJOR
UqQETr2QFzP5XG53Fi10D1TUjdifi/XIobd4m0FZEk2i4dwWXpYS3MHbzj3XzuPI
XdbtH+BGHmlE1Pags4V0OLI3k2ZbnA7CBz70+Sl/DmRc6kxoG0bVAr7EYo+KubDb
rDjwirX+qMp7w7qJO1Aw0qQuo6pEN2FWnpPYqz11tLHCFmGH4NM7K5AAcLWB9jbr
4Nst/7y0Oqsk+s6tcXoB4ycbfn4DrtLC0koawAJJUF/ZRIcHPWUCXUYDHCutPTnZ
Ko8RgqA/DenVBifhb+MS8Qx+W5xdnvLMtlhhbJHS1KycZo/UUGBanhjX5BWC4VxB
+hzRVrh9BP3MiX9/TZrKkbb84BK85o0MCZ8vTEW/zjf+hEjpVwc9tidwv4mseE2r
kyQx6Jitzyj2j8m/uaPzMSUx18AXmN5PYvm2iYLWxgUVuV9LeYtaz6jvVU4kMD+4
3bu8AawV9bfxE+uVHE0feDNr0BZJJQ3CrCGSDSsxo6tWbIqov6QFTjY7/GGI3SvP
/fcfB96gLTzWfnZXjledAzdA615yF2f7nqGqv0cP8um+TsuxYsqdWh38uOWr721v
oxhiE79+TXZfd6cyDuao5zU95AWRIAXsWyoFAE6DMsF+1d5joFrLBlE6i4YvsQ3/
y5pJdga6PwgqZ2gF5Lsenracs8/LTnLDdyLYFZwbZsCxYZTDq+oKLTQVW9oiE6sh
ZofAs+r4ryuM6QqYWCux4wpaAlpLPxv8lSdPcW5Jg1RtrrnUJULc5s+Pa+UQJ8mc
lWSecQZxKjavtvhOSVetUTvju1g9nq95DC7DJZ0ziSZO8QSx1km1rgsAAHuY7SPp
GsJPBdJO43Nc1LyDwFSneP9t281pRDOCTFMGQ+tAZ+jqCZt5LNhoZYNiZNAcbfkc
y9aQ65c2aZ4unj57vFRi1y9vC3EASD8ASU/qNjA9ECPbvzugTOFQm8Va5BehQ8ED
UGlXGp8+Uti4s1kMtUUii+dHK1xOlU0m8xfJxEDerjX+zUxO08W8h+nT8FCJg5BU
HjGEoviczhN7GmWCCjUz3Q33X5Pf/NcXpPn17xt90Qrh4rudv9XVC4/mnHJGfHvx
ZMkHzQ7IxEr6vefgyKQ3gGG6vM5DFecHo53/EJI43Y04r+kFxB4PMfYB6UwZ2HNP
SKNsG5KEsp3WKnbYJGTtSgCGaPzO3cngk7fAu6sxKFxkDnULpasNj9L0ZVC0IL/q
sfe0EIw7zPHP7RuSiB1cqLMna2EeFD3MgbGqx2RKNo8chqIenFAaRUSeP50Ao2Ww
fFm3dG89ZAvJeYs1ASjlwC5qnxDeIIl7tDrjxEz10SlAfQp1fermAc5DXg4zdnGc
++IevAplG1hWmqhq0NOWJdGRv4ifpxzlXArQf75zkOC8mrAp4JaALRezM13HzIVC
wxWcQEBOBDha4BGz6mHv/Q7W0T66lnyK/UIX//xHh4s0R+2gJmfDQTR2otmN+ZCd
o1pfsZIyh26j5QrnA4fTQiDydVQy5AdwMbcdxQMoGr/fx4uf0V6xjMTywgNbOzhe
TCT9kKw5hJcKgktgJ6Qck4u5bZejam6lE0sW3Vu8jiEWX/t6SFgbKPjiGMehjFPK
R3z/4cn+T6q0MqbdKa+DIPw3QSrMBQXwa2H4dKs6gsBL91oIJgultMRx/5XTkyi9
yJg5doHH2U1f253HyrQLSp6s3KG3+Oc57FjRkvcPGPBqjs0+fbxbfU/U5ZtUeltt
+R3tyh6mO4Lw/BH540etYabBlaVeJhqJ8qVXgbfS4pxlQ4UhHecfgt7TaQLiMiwy
947441DUGk6c77CGDlgdIxD8ElAgwAJ0vE+6fp1j1+4h6hJb03aUZ8iIQuEv5m2d
b2CQF5HiO9xm/fos3VggqtAEVV/C12yyp47pgdJ7lagISPWpgBIlKQWexfvubgxb
e9KMMCcaRJjJ/PH5mKcRTVsyun3Gfdz+sxK1xATRp473OeA1BbTFp4k80YJPn3yE
SBov4lC0MRaW9OmjJk9zUG4iP4IBUR0krubG9lT5Cn+ATR+zne4d7mkP6QvYWEsD
gj/f+5ffkPrBphqGT4JHNSFalt8e56i/Ud1yE9fzQ+UFxegLAQUrqD8CROcXrV+H
xriVCx7jon2yX30fUuPZAbSjIyQ/EWP5H3WWN9qlzjkeAuH0jxZ613GFNF0J5YM1
+vU617d8HYIIQ1awAZ9iHAmbi6oPwdZkp1KCdyZGJBnugfwq62BnPiBjWhgFkgLL
A7EGZs6QjOJe7qY5tpLROdJmMggQrKlb8gBCjw4Bx/o1xC+Uj/tLce2iuNmWH8Va
QicATeSTj6IuV7at2BFMx21P8FezeWzl1tFwQl9P7D+cmzvQe03aBfiUVKlpoXVR
7u6uKlcDnfLAZfGqOUOvtAeTLQEekovGp7TECp+FWkzqcplAc6YU2t9zgUUjcKux
G6zvftEPyUHVbeEOHAa+TDRVQldVt2+WwObSYTwtLIlf20sKJXjgDd4zQNw2nEk+
2WNiD3sR6ROuk8JtazcJR6QsTET68QXo6xMypmgKq/KVXy66iLee7OSEwT2yhNZt
nKmcaUTkoTRWjXGURPMtB7xOLjL833xglUderD/yrkTPLVOW5oQZnFY2E72VQkaP
B9AIL7CYzQPJMFQiQgcQO2pr+rtnqQNNywAWBKoxTd5FIENK64DC7NuY+wg8a9mY
UVpkMlFmP9Y/GxCjpD4aZx/sxL+XwOAYPuaAiicHaPiVA5+VL4xmiA95Xx2I6VBG
gZ9vYRVccohSBT4wa+K+TxP9w/DHkSefH0x9M+wrnETEYD24U4o+PVHK0H7XF8nG
XknWSWry+EV23WbPjc/KHlxqWXvqyFn64l2xArxk+OC9/tPrQ7lPMRlhUv2Nsaal
u4w1JRBDBxIbDT5b8lJ32qYZF2yM/IxLc5iW5umoX5j1ViNHob67+gtCTHSZY4nk
BdCNI9G99c8dzQtu1oze5mNCGcpx9mldlaKS2Vb0n3MnMtAP0iXSrN7Hu3/krHA2
4K3lAH6YIJyDOkK/2x1shVx3Xj1ew2GjAj06Yb+vU2Sc68uLw9eQe3LTct5siMa6
pXut9SvqNNw5er+W5qHZqgC8+XWUw8gzIh+dIfQtQfvZqj52/FXaauWh8kv4CFeC
OvxAhsWxn318XIL1SMoCr6fDbDAmXlR5iYaER1KAi9illzNnMTYATKnUUKpnwJUk
d8MyksR29/Kj2Mkli95ZAa2b3y6UJ9/jE9oa9/ojxhR6f06+Kf3fCyjSsF+5A71R
1PojB/KFlAZ26xbUK2Bxym+vxhuVVQ7pMg5jtI47kRqeD82ZcYf526W4jZ53bUOm
PGgLcE7Lf2P38tMXjNIDdsukYgBkA0S4E+8x8bw8vZlpUOnhPjnfV8G1i0ouP+gG
/Earxe8SkKbJqmxuIUDMD1O7sQ8/qCkhoBvE1Gz/p3RpxvK24Mvw1YUozuwukHth
fT85t8CNtUt9UWvC+VS/Zz6/BzKpa+8Q7pXJLgSD4GFu+10TZ0x7qISau5p6RDks
a07UgpO0HsVoVbIeU9D+L1mA0yz7V0aNRNBMGou7P7bWtgM00s4oUYR/Jjy/5cTj
6SoYEQBX3rJ9qO9K/td4FuCLPDNLy3m3LXnvyvAkQqj4/Elubokv0spepdbtg8xF
o2y3KPWMj16S2c4goZLmZkvHiAETqoadHhjQhHOoXUOGnTj1uSQLktRYdxjuVH4c
Gz+v4O8FgayobD+LWxsZSJXuW3Ki3pWWj82EeB+b/A5neu3C52lqS0UTyEQk87US
9aBmsV351QLpLaDrFNKcdxWki3kANQ2CHUpoK8W+lYVVpcKwl1Cf972341Fr03fQ
CMuDmV1wu9gJdcCVV5oL/jsdevB76ocexp0fX3cyR1ar8RA3pwtdYMpL/+CiSVtu
QUlfOdsW51BG2VBS14PcQbAAnkBSfaiaprWyLj/9uIvij7dvuYA3YM/7J4HL1wkO
SWN5/vuvqso/1PriUGaSBmiTBaLD7rySl2tLETd2vdb+HsgMwCDQn8VcvM2jTyqv
xAPW2++gJXlIfTR9O5ugm5o+5KwvZX8frzvBH3EDCIF1/NNirFm9GqJV6Q26q0Jv
HskUskje8UhJ7w21uiZ+nrg7MEb9JOeVwDmOm/oZoVEmdk/NU+IcSdq8kRNI7hOC
mgE82laHmIqQGhV3PYjhONb1QNyxvpG5lMX5IGZj3taqLSgixuob8M+OtIL3PlEe
CXNgELUT4iF872aJL+NK/Eutnn9LFM0iiDk9+89Hf3tp+0RTMgvzzdxnPQFFoWmv
9jmaNcIfwDaVmJqNaDVxH/577K+pBeVXm5cBxzbADv/ktkW0MS7cWwV5zEuVImHC
iTXzkRhQyl6GLVPDqXv0RHM+4IyuxzbUzny8UTWyJbjK2WW+O28ciSXANO3O5EBV
+7jE2zCwxKHAr5PS7h/G+vLOxpIbJgQIqq8yCmTfh1+n0ku1teiZe6BkGm6qp3rT
x4zlREYUd1n8pbIWWsZLrCmzWybJGf19R45i4jfUU+ra1nAtA3ATfGolFBKT39b/
psmGVWW4nvKynHgFsazLcQFYtZ92qBDEkLdiKIVFmETObg8moEctIFDzXpM18PaS
YbEVfp8JZKZ0X64RpNCIPph6SsY0uPm1crooqUXkx5IdOURpglJPmmTrP2i8KVyn
Vp93bvHHDgQSLnOSSV3ua/Na58uoa5rS4qKWoZu8bQS8Ud2KDe+WNsoSlyVrbIpU
P4TQlBsbX+aVdWdEmwrK7CmUA/484PMzZ02akO9+5PKk2IBHNILbVmgkEsT309vt
qGhLZ/4+DdQ3TOBBKv6RXqDQa96l2rGleL7Wi0xa5k6CgD37ZRXz3XXWF02cqy1F
E5jwPBj26LFi9R/1I5CE1RMluLpKx7Sq9AvK1byKnLwcDrfyjNiiYhZ08LqkWjrv
qTmd+QUkqLqMhmsGV2+lC+JWx6oJ/Z0xEI81D0uLmZDE39ct4ojwIuYcc6BTvom3
12hazMpzMQgOj6OiRnd4PeI6aBiz87riuCSqOu/rXSCky6NVcmhUkkcozQK42bOE
+YzWdd2yP8dToXSvi8IW2jNWCJu9OQnr12izof7HG+qcLoDZnjw2nMTQyfm1DbA6
27ti/00woxrMXeqrljE6P7JedgqCyg72K7ebLyyE6WQOW2OCtjKHSl8IgKq/UxZ6
+NR3m5yEi+XwuAy8P2YtE8iJKobcDyVymp05LcmPDkuQGBiOfQXhlMzm1RLMtsK+
tS1imxye2hhWNe3winc/OT2D84MeC/UW6VZRf8ga8jZEtgTAJ4A5duMIo/BLqY7p
CwzfKMF5onYsH7PraxZtpF2HVTcIMNxO0xZB2e5NcBHpcPKXmHRplckm5tILtAZZ
anVvA9TRQ8gSp1KjE3E4X3aMM0rcPWV+g6TrzDzE7zvhxR18c2lRKvE1RD7Hn6f3
//fa//7W4oUN8CQf5srjtCh5lI6F4GqF1aUPleVu8Zi5dMvp7A2TSBlSKaE3iXYL
WPNEZflLXG9MTGU6cSLh0fdiJSLBkbYGrO5bp/gTalCDnAahjrkC5ww/liSCxtf3
+qZYVmq7sFGIYcrBKi1u/XUnoKKnYol9oO6jGTdF4Q3tDeKpPFgKaaLgyBY+lttZ
0/R6+ZriTRyZAecGwuD1vaFw+1ONJtR87PfllIAE2INDsoF6yQFmeM9OKNKrELFE
Hx9wXvQUbxnTY2+mr4YbXNhYVCdo5+3sbKstH9jWAxhC4Er0cLkNFPZGwX8Sw6fA
+5kW00YMPTrGpO9uTpVKvk4IakPG5bpRniURcjo3lgMna9pDmjq9lNEjM36/S/Mu
ZY9HNurgXT4ZTCZYOJDAmv6MYOqUiMz1aTih+oked/MJGf/t2gQUKbtxClyApg1U
Rs9k11UMyveEs0Eun80faZ7HmiE7/Ed04VpzNiHPXwtWzJ/4i+ig1rd5IZpT1uSQ
NxTFK4Fxsj4jzQYa6sX8PC2WxM7An5Q3t2F2n8ooZFcv0hR5dzVsr350BnEdlH8d
ZjcqlFRTGUmFy6kk4p2yU9PjN4XWBiZqoMIpdy9pjIIk9iyiiJ8NgMWpcxK9eVte
q9k2KRZUhnSZVr5EIpkwQ3jrV9SwrNt+j7OevFjYqp2etsTS/okVt49jmUmO9WXF
l5p70+olATtea1XR424DJUscWj1zOi1WYNcuV2VtmdDznROgNpKGOZxMuZtSlBej
le0aX3gu0B1CSVt9/90YjNHI0IBD/jubWx4yqi7R15YbWiFkzxz5ZUmWTh7w1Z6K
3/B6fectVhRDQc+C8ha7vlurlXx/Pmzca0H8dpBTwZUrUAYPq+bRf0UtctPZgGRw
o9pz8luApat9fq3aC5G3sidM2tofJNdmQvjhQwWL65X5n33mK38FFwZJluBOPR9C
hvt4doMsg0I3VsdjfuAIQmLQjXxkTaDWJ1nqRWTms+v2JFdB7VMbBG69vGvRP8+J
UPxHTPekP+6YyP1K/qJ6JfRHtMjG2O5Vg/4OxIqNU+U7FozQ0mn43QUvxiFNkMsF
8P0k2Q8lSg7u9v3vy6zOUluswsX8stUeAawEYN4UwbWa0sbJrH6XIGLiRZJaEM+Y
68JwcE9l12g6b+qc44Ko7FsiCl8SKwjGI3wlPSnCHprM7CASq96FSIUFY2oU2+lV
21TbkE60WZcwnrzUzv32E6d0CLni5R9KxgwDMyeGAJ7wTAcO/oBZeFm6LClzaEeh
YYLvvbrRzFoiiDCraEj6178b8MdQdKJbRvW7vPmD3U+fcZB9eszbbASj0BxYKfFX
jgnjBWjDLpAS9pvzTPg0yDMb+qDc8A4AwoQdLYagk6/nIsnSTFR0HiykniO5stCg
e6vPgpcSYISi5+XIw2m8BWpL/h7jh6A7r475Ie501IgLppOesRSeHYDwL8MgoPEy
pB73UKkK4Bf2dyHhN/nyBSDoKfMJfKYyQNZsAGQvbiV07Ky1R981vj0aPhzzpb92
ERNNDO+nIz285IyIEc7MxKM95PMVzRAj38EtD81n4q8jfYsghpVj+rAhw2pqyQ3M
ZHKy/6WoCc1LM6jp1Elt9MAOkcqc1n6eGrqk3muREbRV1Qj8vhjvvc9R0gl4beTn
vmSKVQJu4YGsihIobSJLF6FUYCRvxaOXyjeaZM5KkaV8Q63wvB3MqqiHM7p2cGSe
TBgUsmGSe+MLbyzihns4gi2WZc1H/Z0I0ksNPBEzhJ16tpQeJdqGwo59LrQlAtpY
2EgduMAh632Jn73WvKBdUE7qzAx7044LjJCJDc21mIElyPRAyYWH2MIRFkFlrM+E
KJJGNatKXf5RDt/CzLfvcScTO4kp0wVgeV14+tJdd4WDRSZG1Cd5X6ImtLdl2RM1
g6MdsUDeleKidZpf6fefc+4iIzqzTTR1FNsBgO96I9de1N8OJWu3vabVVxem7E9Q
Xx+fvAiUHRV9Fe1Q0chYBgoSdPffwlRwleCDnZAQybTTkpdWCZqjaL4o5MSP4M/Q
FNgWVvsbnSX8qKZMKC8nXAlrOSrNYmZTeHkfUopqC6k6zUV23OsnLvh3htr60whw
45+QJXI03Q2IL9C30SEqhxXBinHZw6PJrL9xCGR+EkwYnmFhUDCF2pyh/T2OfXoL
LINhcILXZecndItIHydp0CjttdLGi+xNz6qV04WsV2Di7s6bwiSdgNoyHOz6J++J
8CfNYMKISMQRHXqqVFRDjhPc8ilcUzXaUEWONHytXOV7OtKmjkasONn9qrB+roSv
pghHPFryIP5YeVV8eIWCNmdFs0mlDC0+pGDoB7iCiMuh7ikH6iikds5ilflj9CDd
m6GMs5Hsc2ZcMFk0Zr2uurfbimsy9pB3OjMY1zQo6tXE8/xdRMq73+kBWbi3FO6k
Bx5E3fqPSyA8++suVjSFilW9PO2cn2zb8SHw2J2aIUgDJb9TViN5cmhv5KVyn3Tk
2njDfsdpDAAAL30ALcF7g3xhfBHJKmw6XlNMBnUQ1tNWU5kDpLkHBtxO5dXXOzap
SEX+oE3qVhFPB7VlaUI/tfZulVIIXKnY3Px8xTHCyKogkztaXAHVrPGIAia1S+sg
DyK8STjocSyeFGcf4v0n1l1ts1eMrzAM9BRb6C1KaAGqDrqvzOpNpnJznwyFITF+
KdtrpPqUqPB5dbjVqdPUbb+Q7JBkLBVBUfKpsGMZH1E9u7uWz2XHLTPAnwFxXm96
yI3iUbBIBepW3K5Y7H1yUZ0q18Mr+mybHFEWDum3nqqHp6a3TC+idxWD7dx9YLuL
NTY/Iw/th3R/im51ArbSkBQrogaxIuyYVx5cpSCm/j9FpZ+9qSiYfmjV45DfyJlI
KubLOjJohasydpriG0jN4EqsC6ECnrXXAU02jmomqBy6q5h//NG1Lk+rz1oQTl/i
drRkPTaDj3ZLgQ9xUWs1ocKtVA/YP+l3/kldt0ZmIfWhyB7tBByf9NPItyI5nIk9
scLGyPg5au9y5CBkLU32MF6CMK1IDq/SfMQLC+LIIWu7S8IJwafWpYbEdh0tWrVQ
8H7eh6CBvCUoQ4XoLplI/BlngRgKdlO6Je67+37diKUPsI/7r7L+bs4CImuoQe1Y
9dhDk7s5JC6QKAeKPo2aCFIE893qPFj6ArRxZzRSIF0HaFlTANY9+AwiFhEAUA1u
PB90gED64pk/UAlIY0SckN/wymE46wczuYJj+jTDZWcee7d4/PbUhP7B4VNpNW3W
PlDyihh4SHVpJb4vIbWUHkL7t9pNgEP7bF2miLjzwYJD0Y2bb6sqPIw/LCZ5mFPV
BlFNJavViQ0a+r/1YrPUPcWe2wPqIXYkoS01/W/5kBhwxd8+8sD1RO85gvkS3bg4
TFPs9DQwUeCaAbCQKklvdidGwYbnWASrIuKC+ecpSYZDBy3iI0a1PoVMG9NACZze
PIGbEBE8pEwP8QyheE0apK6AfnwzL3WAJnCoMc3WQrGfxTCXkitay9KDL1eXWlZL
o0ciDnfGxPDT5oFAI+Ic68/fF0ZDSH1GCt6wHmneVWpj6EhZpEvypK2GIVhRXn3U
7/xAv9FVPEd9KMB2byF7i8WqNDt90wJ6WKcrZXkA3jF5IX2wIr+Hn540ynuzF229
QvJBbYzseBKbFO7vPdMBksDrZHFGdWaiL2plYpzVjuFgjitnr+xWky+uQQMbO3Zn
iIr5g6e+hkceKIVrJbzIKgURlbDV5hoD5yMWRi8Ddrm9E8mFGQd8WYK0BXi/GCOx
huQgsPRJRp5hwi+N/H9ZQP9/qvFWYHwRXO+ZSTrIb3um+nRLsTnkyDm5OBXTIbQX
/LOvAmllgXFRsnFYVeOX1dI+HJ+GOoZDFhNpfLMNzdAU0vZu4er8mNOUELWnEmsj
+evFGmNDo/dWTF5O6EFdHU8yfl3isodyAmFrLkKD6yplKXg6I/u1B6Z9cI/1Y0ch
BuhIDzpz3kZ62L9zNz9SSTvJz+QuVP8gaU1YAFRxqh5+01bz2vLLDXz4UBBYDcOA
xj6MXWvPx7u1B/dwBA3xxq8hwJ66UqOj8AD2Ed9pNtGLvORu99O98Q2Vmc8xXv0s
alIgvG3YVHe2cVY8tuiA8YE8/gLQNFkrVFnHoWy6eVRBx4AOhoxJTmp3+SBTjm6A
tBGLFV54WASTu9hMM3vKHzp0/gBedDvCZnoBo4t9GGr8UbksmD6rgMbQ2hafDg0J
P/OD5YirHvRUMdzENqBMMQexOyD+PdWUz+fqhXFK3CxO2nlvKAJdgz/8fLdPIEoS
ZPH1AF5X46JEPLJd8oc3McQHmn/Bo8uhvoiLsc8BPY0uEhk2pnjyx8fh4K0tdADD
pJbZNUGdC+I16Gr9oCsg/p5mbNdKku+t/Mi/m9K9d1/6mtaOSXWUYlFTkTDDnpdx
pteuJvgKBSKLwxgmgr+NDe5yMDidV/oOmo4LhTPAQs4XPjxw5A5SThaNRvBBcyKG
+8qqZB65kpdjOMG6gmc9WQZPCsqMgvCi9qZbg3ibwBnpOy9V8TUJqUioC+7V/1I6
V4bHEpMLwNhJUBFFpbHAsniiE+tz7jFe11yWtfwSAJthclIPh7BUzlM4eAzK25jq
tkBHar/qWwiGQFY236PUgm5c63B/3VXV2HaZJk1lqdrnGJjn4FSIIOOVwEdQOsNr
0e7UaCR1sVhnzYHDheNafqNvJj5rcAUkQg4k8nkuwBeWbDFCAEbr9rgNFJr1WX2l
KivOLfw7pmsr2D6ZGddZ61GgoEsaXCVVA+A36TmUbQP/cwHasZT7kkgAYtxi0Cf8
GF6g0paOFpYGUGBniiEi558eiSqHVEt40rAXGf7pHlDzIpm02cvT8H5fe6HSmmVa
YYhHsdPVrV5TIoEh+O0VQkxYZGnG4eOU4K2KZfKV2cV6Kd6ukRw/e5++uel3eE5t
p4gxmMHbjGFRRzoy1om/19/PJdfTnlTaRIMk4ORx3EB0JZWQIWAXSDR1vK0Wt5Tf
A4wvf0Qznzc6AwbsBVDJLB1aSfDK1zm6ifbw51peTk7rX9KEj24iyPAfBeASx7RN
7yO3fVSJ6uPo/gbXr+9EzTN6NLHb+gbgpOLKKyuB1uPLq3ET6V4jCyPDm+Q/tW+6
QQcgsjsK46+xmJUbMpy/ahL26v8IGp6/zz5bNVuG2spzvoV5UjBc+jfBvGh9/k0q
UALm8+IC30acenq+2COhPyuWi1nBKosBwiLlTybjKzBg5fDfvgtEaGZKvtdqq/8y
YGWsumvRYtw2KuqmO+IsvkQpmAFV0+Jx1dPZ8qi34Jqsg7UoCk6eNxTQ7Z1cE+My
6vlYZfHQ5dH4LXwgtrlWF0lZND5PFF6KjZqyv/1YFPQ2D6PyJJKWrcV77VRv5Wyg
4EAj3cicUO4ddH5Qg3ZxAR3P7vNp4ugV+6xa3ZaZIdnQ0wWmIG4bMmJauY2HD8jg
OZ6BvnvyVd0dG1OmfIX5r1TSSxh9HDmA7cdj3R3SR+8yDENcKjFt+3uUpMgZYUx/
Lh34mWLvK8YYAIDoMBSwrILOeXxX2sesI9AO9qwq9v6Z+aW1DNgTinHOiKD3+hFT
8mlaCPFJaG9ng8eb6G1lBfOQsPBM6Wj8UNn4YVs9IgmZ3TrvIFle15ctzh4R8J9T
nmVNf9Vn+yU0CDuSzS/lftE99KjB9dylx8HaiMTpVjP5A05pUB3ZSWiatYU4FD0E
tNG2b6UzWQ+OHU6vOdZsqJEY9eDwabgTKLgMYhINBGG6eyTD9fwdx761OvdCuYiV
CK53iOeNrZzxPA1EhL93EJWNnxy0N/CtmZx5GIg0dWHMeByvieyz7rDkcyi1oSNj
jeW958GRGy7P+FE/wnjjl3/0Z/bDZ3azRzOFnGCkmzGrwaeFj8D5a8/T+W/Is/3H
9oEhADNBq0qtDzDHXiYqSv+BzaUH9aDTiXsRvZSQrXhmUAWSvzwfGuAvbdM947VP
mNGO6Pfxup6FU3uBtjtTQ7pZb5xtg3UQ+K44HLM/tZjoaoRloeL2I28hXLKBHgl6
x+IfBVXeEvB+hbyQrDTBN90/MwrYRoEdcFGsrIqKqydDX+Kz8x5C7L3FhCmoxNcV
WHPrryGrAU3Bu8qtNO12Sbb63CQE/p7MjHL0pW1TjcGOpMSFw1FMVgWO3ICzOvKa
z+6eNgSuY7cPHCo/MCcNAE/AGcwfQwm6pccKtAj2ihhkeCwqZKII6dXUdVssi0s4
xvP6zeVSx1Rq7TnkAT08RNsTNh+MFwnAV/nVdSX/TcP7Y+wv75h1nOXOyel3fXWM
BKuSWSHo94cgMaphq145GEk+26vGTYx5vpVIPbQZn9LhUnKpIZv4nbaTv2WI5unx
W6m7k5cCL7CsMogFbRrRBnpA8r+9ZWatSq5xbAU8MiQ8Zb89wxcUx1nVpgZixm5d
fSCBUjAEfdC8iE4e3f6oJ3wS4bj9PmZdU+n4zC9QNCmx7UvRga435ng+4G+rC+4V
SPqAquzzr2F/IBL+XNNaTh7UQ2mixcT7rxHvqkKCJbHXPlXBYLE8EAfcd/Mrt/Mn
L6JK/izddwGisxUh5L1Jd3swJWiibLlDhr8U6XTbeolnkaORF6QgdLp2KINB/OnQ
7d51APpcq4sgUlk6Y68LpTlSxFp6cLgt2THBpBxK+CTS5ujQtpj+fOZWROjzi5n3
8ReiV7VQuWJAMBLUVH1LYk6cEPtUbXjdTrPSu+pv/+d3Whvc2Q3UGKakN35UoDNF
T8AOQ4vO99aOBQyU5g7Bm2clyTuaBKQ/epLFwPNfwTdYJIu8V8py9OSx42uuKx/k
ue5/iA/wEZ3GbvYxRfvL8X0aIv3oI5mImJF2gIPclxGd2mCnTf9VRcJEXIoCHwI+
24P5b1UKevNGvg9x2ba43Kv4nM8vNsavyjppP6voiKNNrVk/MmWtU78QFqM2gikE
E8hjXNgBcObVm83/enqEZFeBdnaCwW4Jdz9Qfn1M9HpfxEwT1eznJRKO/IaVLSJi
J7Fr+smIekApTlzifqf58ynUCUYyc0ZX9CastnDZjhD/sxL+4YRCjyFTzbInh6CQ
U84WmvKcj0i7r2Iyl+H0tbBydB0SksHdvB5jVIoI0FpiQCJ/yBc62mXCVurucxIZ
ohKIArIQtFRy2Pdp8isGaClS8/tSbULRbOSuAxerxfOUTId2OrEhFV/WtViNQGWl
JZkOroLHNhz+ttQmvf1QdYCJIcvUTa7swkSfr5zWB+YHxmtZj70aLm9Eb2hNWjQe
SnDLUyuyV+9ZfXGbtLYvtbiBAcrko04Qvd08eSgj7N443a/puQuPisynUhg9bxeo
C4yDJeW8JvBfFjYLnG7KDpgOvdObSM1NCwY4emz24HBmGaqfUhchZjPxVcMnCi14
i/4ZeYmHMJJ5qIJBSyCs1Z5zzz1yYZJaVP/Jplwv0BAwmw6NhKCZGf5ueKJoZyuS
+8IV4vInAgX4AgK6c5BpAARPH/7kKMcHAGPOyUJRYWcVHn/bOL0Kd6IdSzBHcB1K
UTGWdSuxc3avcrSKPN1x8LDomoknfkjeMevVXjuXJbGtOLj95NXtHjrmEErE+Fh8
ssoAJFyqUfEgMVdFXeSme9PfWCwNVEzOqjNyaVGPMD7U30J3gINdcm4Lu1mi5YuM
f9kVpjYoImIuZuZdub0j3dNOST3jwhsZob2/2udTYNOBbXy0qBQZ9Mx/swaqr+Ri
tHmnqFwljlFNFfxwYlFyte8VWPfOuQ8ljMlKEQmZ+VSyH+QsVEyvlAhHHldPTzZ5
v7GbNPQxV10MqOr2iEMmlut6Llp1q1lTlomUHhaowpa1k664Mj7BiLf1ie1rlPM6
zHaEep08vEKN6JOy40xk0aAmhpf2qV4OFYhwX1vyIzwHUWT+btsQzxPt6C8IFlkb
7RGZolVmWkxFvgJYFzwIfCmdESrjFupoEyeKShaZGeO7a5KsN58tO6AooQHagoAs
aE3+GhzaqCdNJC6igU+8rDUkk0be9GlhNRbcev4eBl8PZv8N3kgorNXGekkhcMzp
yvJunM+F6yQ7YehDzkcDhCFWIY4yLnZNlRf4og0XzgP5DFyzsLH7hG81LSE5Bp7Q
zSu3foeaR0FSRXEIemYJ9BaqgBZ0twHelcs+gy0Yz+od4CYZPDf5Gw2S5eNkRQd4
9U+ojAKnpuGzLA9TsACcTuhuQ359pD8sxXvYl02q9PlJo87rV4nRnRQGGet0JJnO
guiBy2eVPwMwRs6VyGAlbcmHDwS4Jdgo6cncL7g1NxaP4x8ISe9M90iVyNnDcS62
1dH73AGYI5JvP5WkQmSSmj7APND/Mf50TBXHOqpXLJimDlqPVnEkHIEyNeLT+7QW
cEsoTehwHlBG5WWVkqwsIfXqCPtMVZbdTMOYT9E5o4p0VOk3nwIx45Oszum4/rVL
iYgha0ggoHF0wZy2Cno00l7A9I7qvjnuvhWWNrUqrgdjca47eMCDVUsiNMdipMgs
Wvo4EF6GF5apihSZNft1yJNttEBBa/ZOXeidLEprmyBaikqOqlsmREI0Pwus56+m
xCi88h3UrsuvD2v290ogYh3g9Qpz/w16j5Xid6hqv6O44lpcAewNAUIPCtjnH5kz
wfLHbFl8tFDfDZQySEoWwFN/NTETNHYqW01B98yT8ewFPtz7eHZfdsmJSNIXE6tz
oYvKAcwJHR4e3fJMIoDFHCoRpYFdiWkbNyxnDOMpp84DdWLZ5sKicyw4YOGGCUUV
KNObMD+5aGeSZo/BJnNF3zNvh8K6j1evgGeQZR9fNLpjfNtPccNt+JvVJBoo0xBn
OeVnzWVjVSs8XKMqxlV4XU179izfPhgbrJcE93MTmInOUqNJsUUgxgQxs8QuuIXn
VKR/kXUGOtBPMoX9lzzb5figy2Bb+fInGEtGvsK9q5f1d6fguZ98FKrW/lJsS6ni
pS2+5EEdTez1q0jvn9JEkBF14BAo6JAyF7S91J+H7VxA5nWKjUSqkN8mczGgawiB
jTNkkFC7RcAgLTp4yutEybWWbBQcgABg+NN7AbH/N5u2zIyDm3B6M5dk+ExemNsO
HaY2liu+/pTG3HJ8nEoPGJv5QDFUma3tqa3oGSY9QVEmcdQ9aFbxLOxyGMzeTbLf
Kamw/EfxN1hN3FUuqopYx2alTb9ETupqhJrwl1g8xfNbuA4/dQFUQ4yUdHPKl7b3
FBf21YCQDckSMT5RnFuzMy+EC5mB+2zUH8RG/DK5vMbfmcr0bhf59JaWabw4Zo95
iLHDKr8JLNjxZejbrtYlOMRT6gHVas3h8A3xpcZ8yLB/mVY7jiKH80Ib4N4CIBuw
VSRvFf+NKnSrswDwsyuD4p+xE9HpKAa+5afRH395F5qvEjUlr3Ubn6S/E2XEgOMp
QBD2BkIdieaLY2bkTQ7pqwsr29jerhNGw+T7k8qFMCFJSN0GuT/P2YkHKrPIVT01
qsQCJ+SS4J55aWTzU4guPceh4M/ntAnJkJ1SbkafKWX/hJ1Tmkk0WOlhfg5MtLbr
XPfUA4eg7OTG4ej9mGio6vvKTXUOEXu3c0WHMTEpQLKmF5LIf38W51EHt/pYzpOy
3vark+8WBAZgRAnX5sb2XMhErrvf6DIeIrIenBNFpufYL6oQq5AA5Eu8kt8qI/hq
XK8Glcdiy8XeXzSHVhDWID7JwWbBsylEqowrPGhNox5PHOyhxsGX0gmvctZAflzw
hf0/i2o3dk/bSoy4qaUnYqXWZ7W+bSiVsjSpbBfDN6FuZkDqpcRvx6y03QlHqdSN
lPSWK/rN5jhjUPrT2vrq8NXbiID83+sDja9F7jWDMS50RzBnTzzb1/Rm+TDhO2PN
tL7q/uYTy24oUlKN7yHshsdZiiZyMX0dJzH5QFCCRtV1eKP2HbcKX86mnnb9oI2J
+pkQf1514bgXBVKZ/p9dbRE6PBwMZBOb44taPG9e2SVq9GiPAzbB7RStt4G/LURS
YVq8mFwe7bGBUJkfExHg0nc6Y8/BYuHWjo++9XqZYqSpkmfBM3uVrGlQ5/aDXf0x
HYScd8yQdozIZ80WucZnlkwVlwQkgDs27RhAeC25sUPumwIgdN5pRxKJ7XNWCVK7
zJtW2WHfbWH3wR1Y94bOLJsioLlJOF1qotepQCDbgBTBpEm7XbzUzt76uLD63Bfh
VMlRvOjOX/Ymc+RRhoLorx6TST4AjyfC5fBAazM+YaKY/keYyWH3gMzdF0gj2Fun
Xslx2o8MUw0pokbSbppAiJ1sNY+HmTRFgNo+cfswnM4cU+7NreocvXSm/FhrE7sb
d4swRGRZL9+ml2zgPXdMrua7kBOq7Nb4mWlw5WaeDPZHWXSLW/bKjHoQzlU5a6mS
nW+bXg5FAumVTzBv2lS/9k/ZEs+c/xMWWXKLtdKfFF5a7gWRtJpuDPpBkMboYK1c
aQLyPsHbKW/5df7nQuZYeuuxunCcTJPCtBsbGEdyHbRXla6RjwgPI2fZFmkimQQR
abqDd6ZpPP/mXCn02Kg6Bjmbbwsy6KZiV35iUd9k6Ekv3H1OyHclyDjKPU7ior5i
RpPk2kwCgya0QZAyPiAQE9KeeKquAaa6gKIQUybOUhIE6lEloBDrGP+QYl3Q+KwT
+8jqYLM75vSGvVG+frmL+iRD94btFj799LDP3E5riPhHaEe1NvUhZRuFVl2lJThT
2oXGAY7und7Gj9neVrEvrc8O9Cb5HC55Is9mxi61j46a0c1ISp4OIAa1Gbhd8tu7
/xEMuwIie+YKJraSsZIyFFVbH683uIm84XMZ1lJrwcWjgQ6WDPAEX5vBfDVNfs7d
OjMrc20lJLn9KZqV/GeSG6JyXV4N85SffmJXtmRWMLINqCpD6OLQWwgDZcYi/UQQ
rHhpcOpq6KEwj7D220S+6Dfe73c/1zvboWK9UCuwMbc9HwQgkJdWHFRXlSx0vwRC
/EknNZsy0+3bV54jmW5YeoJsR6DghkYrIbOzbWoTFaHSXk95F00Qy1T0eENUgoea
kiVsJUKxiKhlgDtAqvKlb+5JOh8+jOpjRACrQw19FlHoTilC/D72J++ry8iM0PiO
TUh1ojeUey3wiVwF/lWps7O0IFUztZId/B6iX+vrWCD9oOtbYNDuEvSxvqEmwpul
354uG+tIRCXzZvGTpA6nx08NGmA6c+9fAhxqlAUhWeVVgTcmBYK7XzQOmiPAhTnj
B3a/gJ2VCNgBpPmVeYoQ0QtPiQInXBQQqH2mTPIr3Xg7vdfAlUpRoO6ssjeKlusl
R6X8q+qc4sYDDBFYK8WRagT33ULSYTnSRntOv25LTipTqeUBbHqkGj5TFHmFpPQw
4pdVuslTTXC1lO7qG6Vk3PjWZAOPwhmfwHWeOC+I7Nc2TRBRh1rLI9L0Zoxk4kiB
+76tE5LfPbyEngrt1FwJKwYivI4Otvk1QNEyuOn36npqVzW9YOd88ZWrG8KsyGLh
T1CnGKjtJjG1suv2qgyxZta0dTvpIfYb9HN1dqyt2noba1BdcrvJW36L1ciC4/dA
nPCaBCTz7sxQtp8tlA02qjMAlYHMhIOwXq9EB9adZ71383ugghZVoh6q+R11oZ4R
39muAaLyeDqrUG3cUEqS5tbVnNg1poND/Q7Tk5KQO0JF/2ku3ao4s/16ZoTLnYyp
O9FDR0K5cni1JP6PjeSN121PG/9Um1xPPTYjVtuTdA7YNGLg36qzcBkJxItE17hI
1kI0iVwxbsopdiObMZ9hkvdPeqe4nECMKdn5H0a5fJE0GnZ3JhJASsayV574OjoB
t1/mbF96ZHvSCgNqfxIvHdUPObQZlfh6E7bNma4yurwk2r7IztVowz8MyK0VS1yy
MEWAgC5/fCPD7hAvYojmwk/X74ViVcKC4tzTYeMAko7TuZe1jhoHCN7rqTiZ5S1H
aLXw0vPceKMoKJQzFhZpBCJA5ptTKYEVl0QEeOamXPDitsergGAW8i4zYeRDATUa
7MWCaRyt6zHwZpua7ycHidvMy8xWED18VgP7lCzzixZoJpNbh00a/OCiswYxNwQ5
mAw2p5QP83v8Afm5BVPBli+7VsKMdJm5QOq0+zs6/w1/Y/EdmxPyVcA+3/j56eI1
T4BAc4MNb/sCGZCuv9UV9uM0MPAaV+UkJBFjWtQYCAirVxj6Zo357a3S9dw/lr1a
J/3AY53OV4R1QnDNLYEnJSq+TyxWQLV8c+6RdyJ5JEQedoZrBMGbFG+9RSu2Bmtz
arXpAz8RitAduxg7sgkGzeff3zx1FiDdYL/Rub0FOus5UtnPPADgn96TyaLcE9Fo
Kj4kUiquj5K/7in6AFBY/twDx/2KzLS9w32DSCoiKRC3HbxY34kZ0hdrSDL0Sytx
S/+oAdJ6x1D4v9CdK/XAJKjTi222+6tslDnyxSx026K2dQVxenh0/DPtCn17Ynjp
+qaQ0tRpEePB+NF4teGwcpK+Jt73zDpcF0Yar2Nz3gVb8HSVvIMv3aqdb8B94JDR
liXn4MhXvQDhxgy29FqWsVpv8Y+MWg/B38kzcFP/GdgNK83OX0SJI0phBCmiSdOM
lp3M47m3QWIFpeZL1omSoDnuO6Ol3uuxLNJVf5YKd9QXQDdzhR2NfHDdzwABuXen
2IOki82A+WbXc2zJiMOSPu08tU2DCjhs1A4wehPJJMVFb6OEjfHqjc6XUxKFYBGC
mDjtLixy6ApcGxsQTWaTurU/dQtPRs8MzOLOkKF2snUmN7zsNaw96TpoRbv3NWYw
NKLBXHQ4E6UhBOTP3RgWnBlcI1tiEhTKxoxMR9LOQjOpb+CxVuENbywV76IhhTFC
8GRhMvIc7A1vu4oO7TyzbI9kbv9DI8lX2cgyYjvgqoCUAYWmBUmDbyWIjfvQRHC4
ji5qyfJebYBMdO+Bmn64XWJ7INfAEM4vorfonTaqLh4y4IEKYJIv5brw40N1FE4H
a+QKjVWdizrDssSBExgVzgYr4tJAHXrZA7ZfoCdhgFGmMu0DeYmecExryY/0K7Z2
LHiNfUY6QfosAzTh/NmK8Q5BSXvXvMGBZLcJb2QdPq8zHKLV3B0jdS86cXFB1Xf/
B0Ko2u99DI6tzejMWJveqL1/K/Dx0gC4mL4wGb5CSs6yzT5MstpNd8bimAdHXsqK
Qp+oX784WRQH3rq67odbEag6Tr2vuKORq/Tv+KyxXLZS3AaLw8N7ncQaKr3n9a7+
ZEHrF1ShCkB8r9nacIR+wBTleHmSAhurLC08HM/E2kZIFkzzI9tai0oVX9SsfNPE
B9a3Q9Sg0LINN5pmYtZT53UHFmG6SyPVSPdK5g3V8wbyNy8zQ5DU4bUEg6lfPa6B
cJ9NVrJpVZ7zQiGXc6a4rSkkdcELfsl/uSUHgjJWanjIXHbL6mQZcs85svTtFRan
spbOhVFPC8mgB995AtFPV2Fcz93n/VDw8VRPjPz+46/19FfWgIX6svEzGJsEBA/T
DBPd8/eeS/8zeZPemOObo2FvK6AFCTviuRjriDNGr8GN6i6AprCP8b4k2vOiOVxy
wwdDEoTAGA6dpw7X1D7HVV7ldIf0jVxwgtduVHxN8uk7z2LhNj11yEH4jE6AwzJI
LT0Q0BF80D2WC2a+qfBDdoanX80enLK6cEU8E5PIofetx5deMShP76eh+BxMfDoD
h2CJtgcuagGoO8aGeDqXZ85A6WinpEO4i7l5Z78ToJDyMC93GMdDOVwszV9t1+e3
QnmeroHqpnVrzaP/76whvxmoJ6FLjVklu+dHg9naSRVeZ+UCDdiaCT176ZrLTPWe
m4vA2bXPt9LdhhThcVb0wvlTAwJl7F1N6TQJ2pzd66WmSheAz3rQi6QToUQCSM8s
sjmaXDTHxw9wO3ykVmq6rtfAmQv97NOycXJt11QJKq8ZfmXwgjFsns1z10UqzTkd
9tSLIHO8CHw1jsWckqD0f5KSLIWlLodGi25BL89pPdveBo3anwnYhfcdVcHLv68M
1tQ08eY/dNItPLxPSAMgyBvEMYtkHO1Ma4r2iM9cB8h/JcBP2IyLUl37miIvWuw3
KXvkuDF50hZ3hABl7SQ//sqeVOBskD2b793wZEh8ZgObPAEF6EXdcNf0c9SrIgem
O0FPBr1EwQ6ZE/iFp8WLagYkY+7jKw45CW0u9gp4tgF2JmDuu8wutS+htPMMFHOG
1l3dFVEiSIlqdZ8TBEWBrgBauvPh1sAePj/Um+ZdwUNv+1oQi4BMIm0T+H9SN3sf
kM7nnE0sByYYXkQQwLdBRXj8BgRN6ODXfvCYLJvTahfE2F2DrNZinsMGXCtUtvR0
wQSdz7I83RKxcJuv8MvBId22x3h90Iqs+T0KXuO3V7lT3UQAPqwLiMMN4oBFOSpJ
MwxHZJuDatbZ3erv4RqRBs9aIAh/5QqKTftVzqxJqHtuQFdUc3JHx2IOMT/KnCyf
sthtR6CcP5WuAcJ590wDvuhGtWF99cQNxay4IAZ51Vsz2fHZP783+gMU6MO9PCaU
6WWDFFnXZlgW2y7hXrKYYefG0nTLUEyBS3/+rsS9Amjru5P3JDXkETGO8PXBW546
ku95ZXO7YNGE65rF5nYNPjPD+udtB3nNgEKIC+09PVpUIX8PgtN65m1mhWHEx4hE
DGEPBpaLddDCpN1zbSwYRssNrhjY/macpiC7LDcgNCLDKFRkaYuz/HI8JhRGcx1d
fhJZJbpFB9shb8pRPQ4NLo4aZK+1QbiH0Ib2OLxtCLzoMcfCCvUoncpDwujinxYQ
v6cVmh7Bu2ezhZuO3QZHd79RT66gD00bsA0lVG3zOeTGhVss92+2ASATklRz+S00
+YCXc7yYpj5dVnG2hKi49Nyxrfvq3cC/tN/e4rRs1a4orksoFRRUC/sWkpj6g/PR
8NuvR3zYdhnFRAKzBRIdQtYnXG6cSdKX/bYPp9Q0ywtFVWueVb4kSqAKM5GUk4Uq
yKn2UkKjsTkyILqYRIFr6SF8eD7/Df6xg4IhGF+TwQ53Ji+0BZ3TqeLoKl+o8Vzc
/WzaxoF1HWRVeHh5A486CYK3bFS0bA8POJrkR51OH//ifz6B3F3No3qxb2JPrP4y
18XWQXgC6jsiO2Wv7+XIDBQsXdVIuu9xXYZ1W2nqU8sVBP3tet+g84TpHbFq4bLl
5qTyjAwaGntg360bGM5sTfufK6OG5jQOa6KY6kkyk1WsJRT7UYvQm56eolaJs9Vl
pAHm8fJd1fRaCD7T8JMEvre2C58jvWqGq7DiiAuM+a+Q1TAvVm40P1naeUdLylpP
tWRtA92sfZVUuluMCiUSINu+gk8wmaaaV4poB6Tx6O4/Jau6TfGZGGTc4qujo8fP
0ycygS9rNosf7sKCtdUh8N9gccNk695VPZRQNU3zsR4wMAiUSwM/rpB1MSupXcKe
/enTA49Ei4HxZX3bJSW5aewaZ5n/vRvnCLTbIP2LFUIz+jG7Z9OC7S9esxhIiCl4
wj/bJ1AnU++ncakxgGtygOaFNow+tmWG444m8FkuNd8X5HKWYL+LntH/KCjxRah4
GYRuhI0Ykhpppi9UE/dtE7jebUPq6QKIXrArlRgQw0pSBFUd/6u7mr3RdcJBA8Dz
ihDI7qvG9Er6umP99epSm7BxhFNK+jGGJpLPMZQNpRRJnnq1Nt3atw0eJq4NvPAL
n7zz8QYNX8buGHA6BEWBQ4yh/XPHF9a8D5YWuAChkpg7WqRJysnm538ykX2oxKs+
+gtHPpoDC6JMNtAvcbSFBU2arbBGcpDHu4wTYDpSFgGBuSEZzFNK9wCN8+U0TwoA
0WXr1dANVgPnlHbn6y7VcxpYbu/XfzxSBCwuQtNf6jc5CXpFzYqxsQRpJgq2RmZn
9JsRlMBozgrqnIEtTdCeiFwLVqVrGj+PhgnsXUn58hYaEp+3SkthrHCoUGhzQ+BA
p1FzQ4PX0lIIx53YroGv7DltzkfXEsC0OLUChq/6fPibeaTU5ecE7MjtofrUIpa5
tguoYQezjBI3KXIAh58Bbny3sySXdikICZMn+LBgwXMFyPOrJpCw69QoySMpJ70b
dwcAsSLhtPd5lvXd74Szh81CS7ENkdmaKlgwTehYkhdHzG9DO5zPfe3Lrg5WBwni
Biz1xeu0wKl92KDadxzoSs16Fgeh4BFTasXRZecyz+wtXf048efphyag2zggWZb2
zbtAVU33uLGT+L98Utplzg2Wf4nZuSsYA9HgIC4TrhdCgITA4Hc+sDDeUkL5XOCh
cEhwqeaYbnVIhjH3qA+LTHFBadOXoLXszKWZ/lOJ1zHcWNaIF8ZCNWeFrFOAazr3
79vrrEmxF4+VYRIDpO1TZ6tOd5Gf+55RVAe1ZLWPHzBPt5D34QKCzNxVaeEw0rJX
4w1SdsbWQ7ancdviUGFUsDLfAhs6TKML6yUD6mKo9edelKa3w7I3//fw9Io0DITU
qbobLOBCvajYrJaOdRK47ic2iIsdanPkQIEEcAaRr9nexPvlEqMpfvA9mRtH1Tbi
5FNE3+dhQBZVoaAX9VCgXhhVhPnrz0NIUUeRJ51XWSjpDptWeQiomM/fFx5heBXE
aGQ5jd+TgtKCz2Xrvo/IhJElNZNnUyYtmsZ4pZbcZw02+IswClfpIOLtHebsuLQ/
eJ9X8QJztutD/i2OsKiYpiXVnQvYMmwmVwnRNvr+plpPbca615LYAut8pOu60LRD
cYPTbR3nvxep50DsIOq0UxvKh09s0re+S1e2BseeWIEqqXz42TEC48xUK2xMkvuO
0lH3OL2EPSXEiREIFCv0bSzw7Z4WuVgiTBG0Tpob+RgPhSzdWvDVMYkZnHOVGz1/
3I9gQ903szhasvn+b1EghR+9sPQ3zEe/Cx6dcpcSa+eCQ77dClkJooX8SZYhlgel
6pcwCj9oRHW2WgUISBG/ehh4TDnupKjUHdODWeBast7iKuOekRfDMxGynPBzQiEd
bx6uRY9t0CIimn9LBaDTYaHsroCYgkHHltmzhnw1s7gn0r4B5ApalMkxO2kjair1
0Eu9Z8R4RPw+MYWQn+nvVQungm7BEPYU0LfbaiDic17Q0yatyH8APNlSKlZD0DbI
76ewiQx6nAS2t+H8/OnTwyXxNRdn5aVt+iMZJwdAZUToTd7SmARUCy4mmCYEMdd4
9YbnmRX7QgbehCt/epMRbma/Pgmo1F5tnblfx1JcWkW4KxMb7lHZ4BRHaYF4pLwJ
6BPOEBUmpc4PP1OUEfpnzVhq1Pcq4129yL9O/iEZZEtZrrerxkIj1m1C244gHjga
s7ifZZBB0KxciOa+qEY64qqudUQv9zVWQ5jiyd7v4Xz6ztoJd6kd5FxnyUhHbtZt
+MZGzAGhYkt1grMjjoLaVweugIEBowNLpgFpi5KLYlnB/nBYisvuQZHiJlWgOX6j
wCJoXbXB5lAt0Uwm+1jA3bSX0kgrrOp2ScgCdfF3YvCCLJgXvQxHE/0GoL2ZRio3
TqSv1dM5KAOoixGUCf8RpgzueKVMADm1cvUhBvtuYQ0X3cQaeCIxQzZSInjC+/Hx
RPSfc0gKUhicaqWYeSpIiDRug0jyedeLTnoBt1uYpyGrJHzD+8ZA+ATbpW3n8yhX
VUXivJFl8OEbYHCi8IV5GJPOtI+xgH+J1RexyuFl4iusKfKQD9VNBB2AiVIWMVYr
xMdO3OphP1gnApIlABwmlpz5MTNlNeQO83JBEdKck5jhik/BUxxOcu76ufO8b5PQ
x/ceWofFRJ8rLCkBHo1qMrHtx++uKGE9VoSgs/3e61GdjJBVZe4CeSnoVb5TWnl6
bzvTQFEHqmCzKJHGlHy/agdTAlVGgt+jbJwAWeUc0LqIkV0wRMoQhfAI/Cjo8Y3h
284jKcgqqU4H2iCrumxX/cMr+MmgUf5Li1z/YV5x5+sHME13ImCYECdxlpQhWUTt
79CpUc8n04eb0wU9JXIBNau4XE2RR5E+TKDWT3QIKy26nQDYkTyp2mYDafW/zWi2
hEGBdT0dFmp2dzhb5v+M2PQmAHO+SIX2ztv4FMhruMQMs1VZ7ZiuXhKd0A/qPzmq
BLCx0uaP9ihW6mKeyTEHmC+Km5+2i75n91pGJNrd+PqNKvgcllg5qtg8b1A3zTCB
JKHbJKYCSb0utaXVE3L4H43DLUAp8VKYRs12fVkNGKKOnAEdb9/PTfwlDEDQRyZt
uY3xePGTWMufR9RAZng6d2Lnx/Pp3EFANAf1ERx0uDDs0YQFBPa9ncxaC78ZzoRB
95aBeUej72B4o8Wjy3FFqBqVyBY810Y91HZuj/ojXUSoV9an1bu/0yw2gZb0Kaf3
DYkgVVDN0gW1SQeyCdpUc4B35SU5Zq1mSqNAs+HsZJxs8N37LzrPO58UbubBoLK9
596gNLMYbRjLrPJlMOWGkn8SGuHp+wyjCX1ahy5Ze+R/gDwJSk7bf7PJG9f5TVJ4
hwLO5SDQX2POwmKiVtu71IgOQMTC34349oBwjDC3ylfokN5tL0qNyKhyl8gtjjaR
tATLnI5KsHvp0TW3kJRJYZnajJdkJLDvSFh4R3sy8I/Hr7ReNQY+b1dIu5GxFlFK
EseeBDO+nXtVCC5TYqHbYbMsNWjvCqZUTLWgU3No7j6mzImn8/B4dieERPVw1XYJ
zX+9O24jRezIH1CZQRSQHxRj8UjiZqUrGogm2N93S+1DfsXHDHO6bLQS+oQd0BX3
JKe6nVT36zysv4vmK8jA5Wl1dPU8tMW361i8TfhlOflx+fPkwN+lqMcu7t+M4Mt6
8vyS5I67XDuzeyZLYr7PziKwCXeKMZHa6qE5xm8r9N1PU8hQHIlsVqZmMIUGt8Ay
IN4oeAej2gPNeriMlEUfBnj/Wx7YGwayIt7hhhkxuC8dB7OOWqm/1aliR+VxLOLJ
x2g/j6QaEp8DzhrkwIsEjkLqttiOrh3XbtDScgSlZW+N8i3Rh1YDFI6bFzR+sS+B
EwraKGDC7B/U1xR5cef/09SZYHpy+y8x09pWafPTvAcS++fzrjXFA2bHmi8UhA+T
i6OVyxgtfl8aXIGXXNr+9M770+fjQe/wT0QMaPT8mOVEzHqJX8/lR/vtvVmBXXbJ
whE5jRC2n3WrYBkTE0QjaB10f9huBakdUNFfWDRzYJ7Ph3bIsA/xMC6bHh43V6sP
fzSQnM8VRyATV6oLejF/F+uggbgUvj6Xt2Ma+WNk2IMCwVz8SrodmkWRAfhCFVHf
GrBHlm+AC1ip2YYMyHZDyxMpKo7urmRkL3xB+WCk+Tus8JdP0PtFhuuc0UeD5GgX
hJ3/XRcS0wm4RuUuoOBzf4mZUAGklLaHwJJGOktS2H9dlNz63FyJUxtajGXl6N0b
Ib4PuGVln8Y51tN2pjgMj5g6hqRWSiOVnqdqraMQT9c6VEztfU2WQNDxvte5J4wM
hBfMaFeC6vs6ROW7v9MEDFFmBSbCDCYj3v8H+5+Nk0d//ho+WLCIGLXe7mcRNPa9
HWh7p59Qy+dOKOe66FgcSLASc63qMnBcG8/QnZ2HzPNmfhP8NEF5Z1lZW1bXZL5F
IvHHlkuUH3oPzfDIczg8gN8nDCGVkFe/w8H3Rsr7+U8pM50mDKzfO564AqzrhZhn
w+OZs/68WdQiYeKjQ3RuBAtODWSJoqa6eiawTRI5X9a8gfOI1ePP57/7e4ddjRh0
WM/p3SKhUjcEcKcpqfA2I+vwGrRG/8zDfHe/NINmMpSg2K8PlfRbgrI96crdEhtV
xBnW5KG1t46zphd7K/vRT3GPtqvW9LjN8oYOQ279oWVasVcaVuQrUXi43SQZz9b9
D8qxamlgrJ9THgpGRwKxctOUPFZsBZs0hx48dqi2tLp6e1UeUCssb+R3rRymnjpc
5XQmFzmPXJBFePS8kkqpup5uplxPUg3LGTw2R60joq77SNrvpZGLTY+kkkmKe4qQ
8/O82xeqaiBxX3LJHGYJcfYW0vhoOU6A3UeGOpK6ZHfP0+a7J/T2bDajmM1NkJUj
kDiu2jeuNd8J6QwUyRTqapPsjJpiBUtz2sR8qNVGfHDlw24wMhFMZKPPofPP2kMT
Gz4GBvxKlML6Dnttx+Jhd3RyCPVYgSXVxts7OPUROw5hrkYk8bZCNg1e0VRXO4QJ
kkZldzxrvLnC9j7LvdfMKLulvdgbuv91TQSuKRlBp920phxL801JZrjYFZaBrlM+
/b1jpoPiB0rBBkBwLuwSXYMWD/j+iZehuQSNzaPxKNol03wX8+4ZDvyOxj8ICy3t
GP9VI+gJfvaaAP4hRj4zvQ45pV6DVclEgXbY2WlGhQuxJs6F6iZYYmkI/q/62xC1
yuTu3H9srUjCBRoQ6R7Avk6oe5JYcHqp3NdAE/MGzENTDXn9nIYIVvG7xEiyy81H
fhg81DEAR8ULhQAabPCmL4kjm5fkZR2qlvjisnALhcOThDsNLGDigDdfjCKMJcKJ
x2llWgWhRDTjHbN59T7Pb8waTWYBD36kMUuOMkqC02J6h8GypoU6/WAMYJOmdu6+
7mKD+is2vWI4oOiT/yn9RAmZCQJD7XOXhu/BLSTmMqWUqhtE9nFBR5uDInvDU0Tg
uL7DeJfW7kZgWEpj1t+POgDIELpVwBIL4suFXMVF/0ZELhcZMxtd5bVvtOF328e1
C2OiwNuzx3w9iJY16XfRA48UDMqD/Kvk/CNZtlXTL3EurSGpIromOiKZ/qiPWMA2
xnQzpcYGMyPnrS49HNOLlqWs54tX8vdpx51qeGJHBx8ANsf0D7FjHRdlpsW8colB
Ihv67C9N5x/fe2dfLfdRZVitmkMmNNOiRyoH3NOK8sAH1BIamA9hyYBEs8HZdQKr
riFwHya4nrXcmKifqHqifUnHBNWXfsT0RFqs+SQZ/LQJc3wNMNlmglyTUSxlTuLO
nRdhVqkfh+B8GkZ43xeGxaCfl8cmZCo+9igE8AszwYiBT11k9jf5hyl/WXZP8ZDx
Kt06Se+/ARGfvZuQu6RJmNIgMn1oIsfJZZ6Alawqy8Hi21ZCAu4Fg3wYDEKOJ0uu
YYOqKesSsB3z9GOHhO3YUvAqd6E06rHrVd9ChZ6eaJ2k3XBm8UYlqzzPBxm/t4gw
EVXcJ5rJVfmIBUoW9bYqY8nAa9ctx4u15hZdfcWScpUmIrVKuI6YE9RxzcEOZngs
/1PghGFn8PLOF/5RgkE0FNsa7kBE+pvlPJJ+WVO2Eh4LPMxShYMZfrU5EaJEjXwS
AXbPXel8FlvUOJIol+qqVzY+cst9qOjwtlA5JzoJgzqr9MtwKDpyTNoN9aMcOukQ
I8b9ZarB99IuSS2/cNwmx5KYQzP5JAcwU5FQSFfrlkJEFZXlN4AktYPiS0OPZcg6
alIlp2/ZgFljMBHQuSbkOXOJo/KXMzouqYcUrkyoSCfapW4L216LuQ4IQzkulN/z
s4zn4a4+FQ46CGct/yzhu2Qngk5ouFTTBku3Zk/7gyL24vapC70CDIGvxhE7VpRT
tQgnFj1yKuJynCJYj7h9VIw9NMk1uNNH/dvkVfB/gsQHgsncfFQik/SvbK5THDfp
WqSp3IlLHj1QKRYgMe/i7uC+it4+KIRoO27QzH/nugLdeH4EM+l/1DWENc6d9KVg
UVc4q72zO3t1/L6rLL7JP8yoMFXGkfRl/7MFHZbvVJYltAHByqM8SKPe8nyGBYn0
WEjqDYRFdFTW0BMdX21VEvzkErk0SixG6guz1RLhPROc5CuC4/Q0bRabomx2LMvu
dgaicdk7PgBOm5T4L6R+WFpBnQdk8vHo+FrUCKwY8VIIoSW+RX7TsDzbPSJJEEyn
lcmJfoLGbi3Yn3t7ld5J17KkhvEHGiu8enhx4pJix3rOuXOIceH4/NUu434ognR2
/dL74DRtVL4uRDIEYvvkmjEp+qg/mGKsmhX23y4/L8S6j9g3Tlg/cFEJksoSdnSn
JYwKB6zFBdpmhyeFdnYs1xYxiXozZFHJFXIUDJ7n68X1eBYjPEkjAfFDsEvn4AbK
tCa0MQ1tLJvfqYVV3w75lhn9aEak8uPEOaeBqlxi6SGDxR61U6J7QeGhcNok1M6C
9OrLXx0pOR1GWifp22b7op4hlAFTtklYK1THpnv4qz3kN3CmBobZESyV7Xx9z4TJ
CGBv4HY39E7lpr98MRiXRBmSBJB3yT5B6+/ju4dD7cvrtT90IlwIGsRoQ8p9pQBr
YOgtVNRbnkn61abwNpqukpdDwnyV0HYVXqsEqSbfUyPjB087GZLm1ToF9dv8z7lF
dG0GiLq4a57j5rIt4zrqcjzcHA6B5W9oBug7Z9qPVFB/cKjlAWyLnJc2hWu27vhe
bCL6dZf2lKBW0o8/xjqZcyNoPprJfk/u6oKkINWzy6NTxFp5ZSGE1r+1o3WKLJpA
uBN2mXfbbad09mbD11WHDPRLzt7Z9YaXfrGHA6JPCNw0CfY/ZPKZMnjvCiQ4v8Mx
54+yfsAfLpG1W2n6nW4peAffmZm/WPkTcgt1YZje4eZWfCCg3ESH1X882uUWSVEP
DJs41fmZeNNFcovMSE7Je9B+VTbG828aOY4/lCvVr8D/xbhbxJekeUJYG9V8kQFW
tEAd62diOAN+PkX4W85A/EDEdpOiQEF9shxyE8J1FCrzmYLQn6FYoUdKHrRpZZD0
sM/F6KkuzIrefd6toUZXzuVGKqNY5gyquVbCqN2zy/o0YkUAEP75AGnQ5EyPCHzb
Bqlwu8eX5ZOw/re5c4/MJ77XFYsQ1C5LUpVd4Qt6UzkXj8/5msH2Z2f+fTqeIhzv
+hurtmyyLJRTDNuWHu5Q/DMrfm66EtYn+W81xi4qI5V6EOA0maWARh7ZUw8C3pvs
RcQwccF/0smJ02JpXrkupv+04nhI/5K5vhNsg1//NxhWvN3pi0+uVwtsSdbVR9SH
ohmIDNR9spbGkys6Y9iO6Tm9NZPNW+NCO/SPrcNfBrMdEP4S+iNLrSVTeyePswox
M+6J3mNpiYmEbanOtu+MDzr/1KP2OQbQkIplNtIQ2LsusGcjPDpXEm8SR57rQTu+
skAArF9aQ8jTYi8rl/PBZRYfVGn11jwK1ld2BTzUrjJytEVl+cEhqJL/QvUCsFTi
9TeeNLaoKYz/2JLPapktIHoh+d9Z74pZdxoe7EVg7Xk4Qahg0KOV0APUCGgyLUex
LpDqKwhKPSY109VLWlKfx4AafSDN7xYi46i7ZD030WEEhHLjHwGlX6k5LIrqmh+y
ynYwTm7Pr6yNAyPhFaprsNE4kK1JL37mjA9Fo1ToRakgNzIz6HP7uv5HKE/2n9Zh
KcaJPWmvvOYA4qa+Tc8cIIRuFgYLDDY4Y7Xv8jMyzJZzkvWk+JTzyio9yUN++YRe
+JOLS2BKRM4xOT8YDohtnE3d1uPlLmo5xQI6ZSkzLTPUHaj9BPcBrIz5SEeEY8Dv
piEvM0NZVZZVzIZVLsq+qWRmAFLcgU/g/eYA3NRrD/aoJZqQ/nk0bEcIpcf5zabj
bSZ++MSScrg4dLceEDnlO/Yimhc5eCRvzAAHCPb9m9vYd4ibh6kpmp1RHEp+e8JW
iEAEr+YEoy+Um9F/fBvzWuxuk9QhgmgJxldlY6LyW7ACEq0cKYLz4hgV6t/EPVDE
e8RqZqkh5jWH1ifG29tNoo8FN5bJW6Zw9ivMWu5SyGyq3SbMWXIwCxeVkBFM9P5m
Ch0kwuXHHm1TvOxIy6IoSOwp4uvB8Br1U8TQeiqyfCm9xII67FgboaRhjyzsxIjn
YO7jA/k21eO4yTF/a8RrX0S9CsaM9cybIlTdV2uXhH72NTv3L5f/14eLZ1JgY/TT
mW+Pjp7ZwfhWuV3UODGjISUJ8a9PxO+HqQrggoZjWWAqIg54EVeunHaJSvb3c8G5
jeun2OYUr44GtCzvTq+52+50pBQYj9sSalpO3kcKPnsJ6+llrwatdcPvFWryl3Qg
+8z284BFTW3+8Pu3KOvHVy/st/DiTfEQJWe9sCkpYlQwQuhPzJUsK75KAbZfxm3U
rj7pOiRAUWqjVVl/VT63cbI7kt2FZRFP7z5zGmCnX54JJNCOGiK/g3HObuvm7+58
UFMuJQ6sAKeo0zV9fa7Q1Vf7T4uvSr8erolyFKMa+cYulksOH6cCUYh5mwOkBF2i
0QPIFi9NqEt2bl9Hz+FQl30DUeh1d6t/be6RmOxLvAVJLpXckR8FlPT8Qxve9eab
1h78FaqKPbEVswBgxC5oQtlGlODaX7YmD2RduGSSaMf2Mc8SrjiyuMheVQDo/Eqv
GZpQbnfqRyc1KaUzfT3imGrhb4UzxCthL/kVgfTNiUUnTzVPJ9wCEnsgx6VjC1KM
LX/a/t78PnCwTWw8xfwf1iY7JEjLZ+OSImHq6vJNJUCaXJXSqR/L/xU2XlRmNaPm
BzfGs7Cq2hi9VOKjtBvht2DRG5f4p5HDgJQHQ6XP79TOFly91SJ3rzf/A+MO8O/k
RrUN3NP+pS2J5S5cCYre9bjM7g3v5wblk/5UnIySWOWmkuy3lDFQSjr8Pr5dquiR
QudnDea5Hz1jnxyZUpypVV+HD3BLviPcgXW72Kv17k1rq0IaQTejVIdeTQZc+eHh
2ohsSwBhB0dTuTnTU0wtZjaXJGLDYucVHwqTATCuuBMb1BFZ0n/t38YA7e44JWrB
Kan3ef39fv9qIn7aktdsspK4QEF1+5rdhoYeoi6MEBcJ0vccJa78TUb0ZAmm9NOO
g3ouDx8SQpjOzCucKyVey7P84EGlYLV7cwaRFVOnxlp/Up9MwR5j44rJdrUdM865
YnGsAcyLrZs9q9HGNjvy/hBs5jq1xblfzcgerFeMDakjwIbrDoV+fiOBsoBVEneC
sRfucsXc3AtSm8EAcdYrbgjyPJmn5/Sr1/Ttj+g07j+W38119w4LKcfZZd+ZmAoc
rx5w2KNeg3GvkDQUKyICSnn++9RK/9ovM3sHNKwrNDEN/6tmR6Kd5W+w2tsevko4
4L6GS6+vPYHeJLBN1dTu2AHRr8oMnslxc3y7uGVzWfSOUdZCJ+b6BxnYarR2kk7C
gW1aLgdS51CSaHGdWsScJ+JrduA4q8Hegsdm3qSYSVZ5yjgVGXu0slYH2DQSs1/w
cqs6ui+m/K8+/f3Zd8eDmBuI6BU0hRRmNZKq7F8XBdkIVCVvKQk+Z75ZNCpvlYCp
u4hut3JH8nQdGjDfEZGMBEXG4PCOazQ3kDHnNS6XZkF7kQL2srYa+tJpZsMY/VLM
ZiccUIE1rfD9FwcTvGw5v3oY2V1+Euf02AHCUlVI6pJMRl7pvn/Tr1AEFUyCXQ+W
XWC1Nzg2fYhoAesTN/0+pFa0TAL5CqV8tg/w/qL08CfaL8v2iRG6Ec86g+9ip/BL
XBcrgp9wUUcwmZCsWTm9Q09YuSFIq4PfUUH1TFZlSvj3IZEmDpCxSqzcQDyXeF9m
tceGCGHPU0dJl2qbZ7zRoGU6GV1C0xSMeQW4lCTVQqeALeKoOfkp16Aa22RD8XtQ
1Zy0rB4Klc3aGxZeFDR6SSiSf6nm4LnKoOyBnsQEEQaN1XDygSY8LIoXPyhRUU3D
uYx/AQFOwqpGcZ5goaJM6WGudQV3vD73KmgGfRXVdz1MyvYUWzCKWdW9pQ6k7W78
80+lZ8xiaIYidndD6ffBkBJ4zY+u6u2pQ7D4Y3jeticsvks3ZPePfXuKCdMevB6t
VIB3sGYhJIHGygdFNeBf0jy/ED0n6d4TVfAqxsg8d6HLGHQEf+bbSLsHAnZ+IZQk
Ttj9TebJMistBzhc5aO2/GucFLAlT5XaSoxKFJpFkll7Qj7RDlQs9rr9uS5Z8Q/f
5jsSk9MP/apGZFxEMKb2JlBUjeCRfq7blJZCh8K/mknTGutB0iivRGUVbkhzuHWn
gLpHrOb7BSg7UsiZHcLtlGKDFfBwy5UlpxgkegrJ0WLtUyrKs4kNt6iLq9PAqwJi
lER/X/0g94zpD2LdA513lB/hlgjvTu81WeGKu1Xm099wEEHKSJEsvr2HzB8m+iAB
yNite2VAgZ/IwndFOhlJo4+Yy0c94Y08yazSS/NBl0Trl8gaKDhdX7LM9Y4jib77
k4umqcse46cSESMoQ9ofWV8nOCTO7tIkngid22gltp+arWWmwFgN6eLzE//gBe1W
gV+optYjuh00k+tXQdmvpREiEqrLwS4vB/n4d7KKJr/+PrluqjvupesRo13W4Bjx
p4yoHooqLcIk702NMmpyKuBJ6VP4Q26dYF6SFq42sGHU2Zsp6csNrt4ix1oNbFks
LpcJtfgFOExGlVL2krjhWVg8Xi9bfmyVwGIAOIoRKi5DuvhhURlqk54/pR99dTRw
3boXLEdf0Jecl9+N8rG1Ttapb5fLFde5SvKGgxeUkZr63iUw4mHv+BZGUkdC81Mf
jjHmKksMhBRGbdYZP6VMwDtSqAmgiiBX0ri1iEkSbrkVj1piPfH/yuHQALj1GZTT
6VYLYCpmQAwDH3gYGggZqoFit/AQUgqQqoa2bMF9OeRxqEhuSX8yvCJUbaPW/RG7
3xGvhd20DD+Xd86/eP58v1J73RSDeqyjMEsiawhAyMViZHlvQ1MQ8ckKxvMzyyBS
/e/F4FuGAIG5Aw+1F95DT9lUPbf3VY6KySkyrFmPpv1GcNMykLifroCkNTedoRPr
l28WWj2X0cMe3EFw911XhQND8955dQt/3UYXowwq3a84sh1FumNd6MMoxBiMcEN6
R2/AUeXKQOuNblf4CQHUh/zM445ajYA5IAqA5NHXugKjVpEQ42esp58uc3CElIoq
HZ3YuhTmmhDkEWlHJ4h26tMeuw9f4k1NIHZRckenYhuyOh8ree33VS8tgXT4FU5c
Yl9B9sGkY4xHX8GtH4gN+3HXC0Q83AqbgTQwj3llcl8P/BQAJ/im/G05OOZbeHYv
v/Eyj/zjQXNaJdAkC9Opv47n8mwtbU6xp814LD0ue3nBzssEyfWyj/gczD/h3Meq
t2luKi2hUmpGlVO150wHngt1PYHXP0TqJnfxXAKXQ6shnxJVufAgsowrYfJTOVn5
zsmvelaSr6jpEmFiFXQLcWS0ZJtbX9eVE1KN55/yk3OCr0mcPgGxR+qOIrTYyAM3
j0dHNPvGQOo7JZJApr1cxdG1vTPcls0eBlZ8wHY78h4e1G33PPrbfjoxK+RzLDAF
3RrBsPXJIAQadaB675IL3PrDeDJjbw/hetF/BzbU3dT3GEL9jTPL4/fKOi7W3PZY
geD1eyxM7mjumI5x2FZytSQPLU+arM2tXxV4a3RAkAJTpgZOr4BgY4fPsNbCDJQp
lVGqw13u1OoyXAyEbYyQUu19rfEnP3NYQa0RBJ8lbVpgeL49Ju35rWKEmWxxyOt0
jz4P4ld+tmPgVLISOW+P3+bMGwQsLxJCskWR7U/e1hCTxhfBaOR6Ki9beQKOcVbE
p3mfGOsBiD190axpucAaF8cZr1Kd8jTLOceYmCNJfakDORcbmBHMJ6MGZIMTN+bI
T/jlIioSwkhTT0Eh9GyVBeggP25DmPaZ+mrh+h6aMSMy0cRpc1OaTKjaPZRz1QPJ
N9qvipXm+RwzjwVWFX6Y9haF1v0mUMv1HOusPPhTPKU15Y1ybucXzlwNv+BtDCZS
GRin/Vrj5bEbTmAmehd9YikOVg08ZPGCW8HeDa7i5ayLuBhwqy+A46hopvx86j7Y
wesfQ7+S57VFLVWQfsydvZMGtM5XNYA7pveSmlxlqLiL+SJ9yia5p71Lu7a0ICKl
lavP2Ed+2x/HabygC4bY8IBQYFe8xU2Wqyhk9EJCBxQFH//cUZCXH/dHCHgwDWjG
/+KGa1lkhIB1UKs4k5TlVoEIDGt5v435Bf8bRVu2Sj81YTXOMODQR6HHALjYR/SH
RryUaC6Y6ygip3ilK4i/bgm9oQKOXxVsYS29jX2votSv/s0D8x2RHUOEomwAgFaD
ptJuGDw0fFqAcPcq8FE0I5zAjZpbK7aI+hqcokhBMT8VCGNVfvhGnhG9B5YAeL/F
lOFTyLTtBC7wicP+fmNmxxOQMzRvV2j7kmvyk3UjMM7yFxINx8wsj8PG7CouVBOr
YpL+YMI6oM0w+IOcOmr5twH16O1xdC1u0UGFu2f0U/I4h20BLuUMBkiRxF6NP4Xv
h+xooWmufpeQC9a0qhIHWmAvm2LVPcFvjZJcMaojOmZnK4qY5T50BTSc10R0PQzI
ApRUqFRDf/wMo/6+vIFVvRYUjXzPdgBoI0fuC8B+e55yNTWSAaQk1Zg0O5XGxRH9
cV9mh7XzM4NNnK/ELqsJykonGunxUHwefE39o51aIL5YvWKqxG3q+HrPgvwtqTgA
Z/z5ReTUYzUQ+Vrj83LJKcFyiTZ+r0I/FQoJDV2Uc80Qc3LfEQoKgS/QELAziMID
PglI9opQjBllIkfsUJVhC7J8Hqtkl/tLQjrOC9ctU9A387gKHiHIYRwYaHPa46zD
B1L/QfSg+g8EidGF77IBuemlRERiCFAfOAulbFv4nPYqGMu/JrHZCSjcdf9XR8OG
C1zXfRg848FfKqtkwQJ9sHOjkb+3gc4KnkSRZ2skgMB/jFrlFBH/DpfpOxi45TUu
ET0U53p15DbVzTdH4zbesl2gq8G3piFlKtNqgWtOIW+mY5Fy/E4IDoeYtCVWNxhc
3PMFaxMJB+Dd2uW2xyMAN+Ig0blweZ0o//saov1DcncSVlN4XkcFSOTeqilRGsqm
UBZEaKS9EnXmaQz8FvGaF7nWhL4KMWGH8gGJ1o1gC7YnV1LgJzJYXj0IKSo9CNGy
5bCOgo7SQUx+EbrOVTn1AQxp45u0ROQ+etVaXb3LVQ/oaM2nnx/gOo5/AVfJ9BTI
WByX9EuppSzcKWpjqHNJbDk1YgWAUwAGc49EfG/cEv+RrsMb0wL5brVyYGHBJqf4
oDJ0GbCMyoGO6cEVc9P44r1B1YGSfGo5OYbMjCJNLGkbto2EMZp4QUnxwy5sJoBy
33wj0t4PNjVvb5gKRSjEUrhp1hBTv6xaT/ebQpxyieLYzPjiKzo1iRXStiK/fCvU
SNdJwk17NK7FbMsNoYTwpss7scs38Ttmjg2oKAKZ3uLgsOFndwa9WIerRDXxqDrY
WWwc8qmIPYlVG7N3yEvP9lUT0FgCYzAg3mxdB/jUnUUA8aAyKM2aI/5WNhGRKbOM
IWB4sshUKh/OGmRvXjjlBpOHDCUAl2zC8gv4nn9XEkgfn9ZBkq/ArwppNTG+InPn
nJk7iFEHX1ULiKBbEkLJQfM8rCgr1GdEjSxzOdZgjaL3Am5F7a4P5GtuhfLws7yi
XGXiwM6+VUzYpwTB5Dom11FAP7noaIocq7KWUDBfyi04Q955wyrfM6uti6omspxo
TWZ2xGw1WcvZQm8NoBrLKjSpJ7b+rUwkeadB14XIsfIK2Qi1lDvqnAAjcimXOojf
LkCb/cq/qUW3adY9zrM/ICimGmpPNYw984s7/5igCKvtyhQnpG2v6cJZgpaYv9DY
UCYhHwye1ho5wG9GeqrH8/ah14xxJdWkwvrscwIC7XijpUIvf/ZlG4/TxyvQ/vdN
lLpBfgZEZQzm6HuLCJrsLAZoQe1GJ3NQaI0ELqxmvBJPEVzRf2LrELNcxC5xMsVX
dIEpgIx4kAbMkHkOdsC1pgnJYq5k2ghexDmXLMZcXroU2Y232OB7HPF0YrdTMjeb
cdwRU60BV4FzuG6ouDdKI7bpg2RgF6hMZ0r53w1DtRQADxiHIjdUUDNC+iXIkluK
INhAPiQbFxGKUzBmabnUh7PnokPtxgys4gxkZ4RR1JNOqcYAOAkgJec9AuqaW8MC
O4QteNLa9mCL7D1EuEadvkXiPQnVpAUKZzxj29PsCPn+AGmQgigP36WrA4EzwF1d
N2u48zy0INWVX0DnDUnY5F8RDsGsdLGjB34sfGZffYiuvwyon7zR4xpJVw5nkQmz
P7uuGg8rHi6uPq2mxk08Z8tHl66DNQ33ry9viUGh9M8sUy4iJSq3+ZkCjnnwiflq
5Y310SknsG7hzokQ1VPPCHSMEScdx80T72YL2Fk0lFKdITEqcS+OxZajt4ABJjRK
8qz3/DtQySPfhdJC39KEqnV6WwHK2I6//+VNYCaX0j4+0wBNFVRiMcUKGQZaEowl
2oyXPp6/7NnukxiY7JmSOA5N3YXhykhnFEUgsr8w7qdBQZOsyw+MMD4+rRwjWmMa
JfWhBnZi+88ecQqEiQbBTDfVAc38HHOTm4q9SpzK9d81f/UjQSx6bRBQOqXFVNDN
i8RjbxnNfrQMuS1ZfLQ/bSSGY4Mq+MhJZKK6rueuryOh9kXyPRUAwkaRYthGqqE/
f0Q7c/w4DTF+WZaYM8TVzSu2jfDhvfBLWQzW0TPHQ3yzbjWiOpnk2qx5f8F3fLgZ
IPKdCSbFIeAMVnUI3avjh9RHIqmrshab9ie8eUeku1Wi7WjQCu+M3EDhMQRSJHea
RAfv3uoKSJvfgqBE3tbmgHn2/iwZtNVEapuCWsgx86kTUHaTf7cSSf7Xama57RZd
JioxzrLf4voY6qASP0lY+jyfJrqDNFOJ+uKes3BVv7/64Fe7pKKeE6tfTiZXeIez
98j7wy6sH903i2GSdbGw2gueuyWOD2tM5+xpFZe3dQogFOrEtixDcaApu8F570IZ
8knzC/tzUm5u0MmjJbFQ5qerZY3LOrRcxFH/XOkv8RCFzCAFos0B32YpAMRIY1ed
PgS1wd6MCEva4a5mBkaNgk4D50kptqtZuPu7zBRWihplTIIVycGePiT29dcjtHI1
ySE92SHpNhrNzaTEdMglJ9nxjQmnpRc1PUENiX9Pxz2/bk0SnwpIAGLbaSv5XOzc
2AXA8lmZarF6U0IrwgMlAM4Ere2uFqGD1bFz39y0UMDI2Mz0xNHUXDQ1GQxBXIyz
hbs8SN3SC/YZFG6npbN3d2tKYj6EQBS3Kw8wHQlNUGOYL1JqAVyn6mHjxcSXk3Zq
zleCcJT6MOcL2OVZfyU5I4YRFWGSYKlqEbuYRJrspVWRgyoDgLhAWAtPuRbO+DAu
izYAH8y9PiRs/g1spCpvjycdr/6h/zFgdue5ZrI1cFYmy5Fjp+l4aqVbK2mrZm1e
zhkApDy+bE9u5hYSRMds+cCFfcjHw07EVrfa5LyMLS0MTQRza45z2sxjJF9thhZO
6iLTEJSuXbE5HLixAhPf8N+U3vIyK9W1yrR6JmydUwJIZ3zbqbEPHYQhDVvG4M+y
9xTJPgeoIPzn+kGbs3wr1OqaZf665h4VmcWobhFv1yOT8Ko9zPLC31LEKi8z9oaW
msV9ewIPGXgsg0LB8nob9pvMpoY1V95I5MVMx7z/1rjTG/rD0/euSQwVYQ0kDDvo
is7S+mGvoOWfELGypFxEKQvr7cXh+Pc9oFEok3pdDcHwU6oUOM7+gBQgqV0+lSSi
Gfw+5zXkQZ9LqGGBbPXS1GHKebEKS/nz3b9srHQorS/q6bYRUoNbngd7Dot0OG3i
PLtQDMzMlFUbQ/sghYRze6SSyfcQ3PqM6+GjybPoLFxry5RrqmekS/mvUykSKYbm
lFVGJ+QcjedpLP9URGIIjFSk+xkzt27CbwQsDFB0tnfmp7Cyss90MmynTrq1CGCt
7olAMxL/PygtyZlF2zG3ugpXEVCnFUV5uFkHgOVMCjm+PDCZpLqmy3DvxsBfp+zL
E4Kv7MVtaHlUUGi+bnH2+Wp2vflVGVAr4ir0gzneJM+EnvuPRm5MIO0RS0iN2Cyu
N8KdRxUgYYN1x6uKefDUI0iHjm9KG584/Nou2/n+juMJjgy8PXfn/Yn8l56647Mv
PkTtMxZ6qz619xcHKI3UkmqW2K+m+2FU1qAEYV/7GO4cNBwBWTHHBODBzdjP0QZO
rJIUxHY1mCBs64h4osg61FY7O1TehPgkEowT4K9g8T7etBszcVuF7wcniWnEpDzW
ZVilV9w0D9tFXknwr987tS5yThIESGfhH66vPXLTjQRRghYlleQWi8aZGQA4iiM4
zAyhi1DUpQogjn8HU91meorTNpkTnegrgwkuRO1WUmeYGe9h10FGJBLh7B1bnHsi
ygmA+Xbhryz87XzRK//hZtzBmaiFXRqHSC2NF2wJXm6XjYD5rA/bQ4ooAK21FIWX
1P5wCEKjNg6+ObQsYAj4MHx3U+RK7e8DvWbS0gR/CDN1lC1cb+ubtYKRtXtAIjKS
mczqN9uR/FJ1FoDvwhC1zHi9B6PWDsVl7lX3ZIsEHJXY2Jn7KLoD9LKMfwK7h9rb
elttdvsavoj6tMljuY2ecqy2cTTTjbjeur1cUIRGBGVh/0aFzBpEQep8qzlWSqOI
gRsseaNbEVaB5n2In1w/ZvEofymNi8J4olUZAKIyf9aQcW0rXQWq61ocwM7w0VQS
t/MWMsTI/XLOBSfg6FyEICJx4Dad0ediUKffsuY8r3jNsPgFZdIx836asnqcBC6B
a97AiqfxvsDVHxMOs9rz9aFXTCRJsk2TkmgZjMr/io6uANpaaJnMR7LAfVNzlNVq
jyMVMq2hHkaATH4sU6UbuY2z+kN/ynsvuCnZ9KCEdum+MUk7jdwKgqqBneg7d6dm
ooCb+A2RpC2f1w5g+mFEUnH3VGwbXdaNXImmPxKGzBGYQ3gS/PYQvkfoDT46MWRK
FirMapuO7fyK1ur0bIc9dj6O6pnIPmTmZSN3OPBnhQiL36zWCxi09qERlmRUns7F
ZXxktmxPjBsWovzi92kL4YEA7X2duSVDqV5vjseJsRveeiOtHzsJ8QAljKi9vAxV
U+eK4Q5ixi3Wyf9A/zI63pSYhddFKpaagw/Up/GUN5r8pkkCGz4HpFQq6n01oJPj
5+GJCyTfe9ENYCSc6NpdqpzXKe/5UEPiyRTnEnPJ563iayjhGCKySB7S/yp88Mrg
u6TTjhLvdNMbyFhDI0Mr8yXu8CWk9lntHh3Szjy1aay99qipX/iDtxj+c8qFKmXh
NnI8NfnWPqbJTfmr8aAyzTHxMYuGc8e5UmrEDAe3FzfLtJWid45KzSDvjsJP86qJ
9tK+x31N9em8f9uJNURvaSP842g/TFLr4yQypEYLxYNSSTpYr4/gXG7uW1oDU5mj
XaE9Yx4ydxYt0epsZW03Vhck0H+bIrOGXBdlne7qSXM/xWyihztqho0SjNizfvBI
PQOJO5aVy9feLbD1g/KmuT5u62W10HOrfUPycKNY0jzkAW7+sUGGzSj1NyIvcI/d
mTiRiKSgVwLU7dNsTuQC+iCLyUuQicOSrR+R0VlIhuAyySkomrWqoXibxwIC2v1E
ZLDE+JxIdLbQEtwWqCL/KH0lF25+JGB3C5z8Q7wvjMX/G8i+ptlNBZY2f/6MZ2RM
y0U7tzxIDRHdzc7yTgPKuL70+WkVdYfqSsBF10cTbb9u9Nbmgv4BJ7muFGCt+D50
kh1L2/xSgoTO0VsWqasQYf8L8lSERxI0ZF3Cu0s2tBks+OESONcHCp3o711I4lOk
dV4jqaIT9EZAG0MrX/1dv2r2xFOTHsQoBJZX6LT258F/hQ0tbhtoLLKnp2Z0ePF7
QEYYNy4qK4oeLf2KjSNMkIHbX+FGnaCYvfJT9EELAHBjT5WFsqwYx3S8eLoEfHvj
pNxN4TM+Zv0MryyWrZpHZ2xKkYNFZ3iJt0TmneEd9mf2cDnn6PYX8vlbtrGeY5Nn
VLuUyXj9eXoZLasZ8/lochs9knB77Ei0Nwdk0RaQrX4PwwZ6oin+VpthGhJA+vnW
keAkRAlEdNBsiYAycAISjr2HrD5USDxgNe5ClG56EpOaShqHZQA6nNvtilxsOWxe
d0gHwa1d1DBFT3L0NsGA+ALFoboyCq557K3+2UXZqLQwWe04HfE39NtL1lnDOc3D
p1hwFPv6UHX3SOwqa4tHbExu0D7yhEJ/M7xnzsrVjUCd/laUpgBBoQhWXxc5D+kd
FS6YrvuXBFHtsj60/dFv8PV7RdVx+gJ9sNlR6QdHf3xEXH3tfWtWRgQBZewyv4K8
o8tXkfRGI5qbOTdTHMHJXpwUb5/iqqL1cOO05k49zLZm4R/i8Tl//K0DeV1yOoUh
tSOBf43Y951+A53h5+GbVoNufsDHmPTBIFO26S26L+RSg45agd59eO5G4y35jI43
9tLoFw79hLXBiYv5tU5jstL+7P27Et5uc77HDsreK+3aiVtgxG2XVQN0kbIwKTlh
vgU1oKa0eopPg1xuTokfvLcfz920j4S8j2xBKJVAk4WyQOtSlsSzt9j0hLzKhNJH
sLy0PJjZgslk+vhenSNYe8WooBLegDqnHH+0CFPo9hrdCIc4pX8qza+WX/Yr3AXh
0p/YKGXs7MHRDISfrW5QmxZVGq7zKiEIA2ChlDzZzDCHDVC8COcqSgUxYgXIrkO+
IALjt4zKhO90loB5uRuCDNDX4Ashy8uF3WwCa8Qo+gSljoA8r0eU2FwL1xF8+3SR
DTfKvODa9w3gUhxfPnjknJDrCi0auQsOYPsmctR1+1Nm47sINRO4OOsokFGw7uCm
kYhvyMhQcRB/FGUONHFxnzhLXH7BSv/UjT0Mcplcc7atDz7GguCjlyoW2Z9RyDoZ
3PRUwqfHv+NTGNJqxj6h7jAyjPRq0EagzyauT4bmzxmZJh2nBjDpCAXIORmcjkrc
V7dUyFjzlPF7zFAxYFgwWauuFyapu2lJPMmDmhFJXzRufnkQtovUY9YfylCRJM3y
MIZcjL3X+iX1hw/mcd7wwbCYbuvaUdmUFo8sJO6wMUOHPG6Yy6MKUe9IV/S1MUWY
Jm+KYJ3hWAlbk6ofbCfLMR1GK4eMOuRMFeDmjs/yKIdPxI5lEcCOLNJSDJ+TObIn
UpwVZm2w3LX1kYAxp3rBwtmi6ldCvORh+BaHkBQztt+1IiY8R1hIhvEahc0FYgSh
HPwQovLuIf81WMhVak2T49/KB+j6sa+IvQUKxIhB8hA8dQ52Nj+VIZgrgR5FleBi
QhTwalftS/Sw+3hK9eicvLgBAigvIDoDZrrHxHvWJQxF9gROPajkNLirjpj4toJc
q+0kkCgfyRVsh/eXYilngwZcIz3ZnJzNNIyVrU0/ROo4QZNJ+rkL+ue4oFujP7Z7
CbLplH49/W2i8/27LCmh14WZekGWwdUsq0xMjbmjgNNbmsEFecrYMihL5IsXalAq
El6c6ofpH8tG4XNg54r5dksdVAKX8IykTL+btjPtKgQNHZMjlcGM9mOL58KoKshi
mkzTM5fiZu+tmaWCtqfsDSXOMSCcE7BeS3ykka9Q4NM5r5VaQ8k/U8AoONu2AdZ3
3f6u0/WW4JTmJkPCOUwWdkue7oQZ4pWvl/WqjZ1iOffsZCa/GRCuTNxgTkwgVG2C
DRP/W9FLIveFBET8GLNi/PqE5De29enFhlPm30DM7LDV3IfiHh59GDN1XkImyVI+
ENUnmmhOuv4lxPEmskLRK4AEy4XDcWCj663tB/uZ8/BzF/rXRBYdqDT0yVQ9HsuD
HHtnLQ3RKQerNGAXrwrtGHv0RFGKTMPmM3sukzAPnmIeYeir/dKVCTiHz2i4pxZr
4FJMAsQR1smp6yNgq7df+0g66LtDq+P2m2H3nfG3kbIuc/SqlC0WEtSOyiCxTrSy
ELnBSp4nbkkSUbiqqyVlMhrVbA+fxv8eMfyXV2FLvcaua4Udm9RRpSRejEkpca01
hdkg2tMGAfH818sihj5xB1uo52/mU8UPFsItbAIFUuwwEGE6WG2sOI2pkR29QPuq
LkwXN6WavKLpEwxDS0Th1/WOGCZUtOVscrbwN7rM/QG7zfuS+lwKb3WfupRyP/Ke
0iIXewQHSjf9rCgAdxudKKSm+o1ZA3o71qYHNzpsxlqGoYB002BQjV/9wldOBJly
y9TlJvoQ0azSJ50V2pb2z8fEuMovzBre0hf/CWn13K+iAz60EEmLSVdv8MymbHuk
pqsq4F2C6HorovCk3Y/F5Dtj8qFzDR5CWBdt8UYQcYIGR/l+xGCKpM6X+ukir7zb
wqkJm8qIb4FmasbcPrs3jckikdZv7wZn6zaxuLDSjDG/h3mCr36PWJevjz2upPiJ
/oJIy/mKuvqoAo8B+bR3Yo6JsKmEj/jULdfAgKuc+FF2Ce+6ZZDgg5aY2Cj9s+Rv
kGHfU0FTd/hZjTumC3Hmh6mDIQdSPps4+XyINO8m/Oy6S4r+hzJYFsExB3LPjIuJ
2bP6vy+ulyOuuljRwaEghLT6jaGA7YLMMvfdVFJME/Du4uVpNm6k04+hI5qJSdac
XrdNE2CQHitKc1pWSW52xsWCmR1cAXUcA1gnQmjkZB3bjZWxpbBnsOK5UTqlsCVC
3wGEzSxTxa1bH2XA30cSniyL+biUqEBTrwFL1ibtf1EVwxPLqxdZyAXcIs8lkNnq
IFFL6IxVuTzFdy/ToakzI0g/6KAI4WsNT6b0R4HwAHx/RnBCYNKOfFqPenIS3YtZ
DwXYRF/IErMUUT9gW4vuM4ZpMu0mlpz/w6dYxySFpnNbWvo9I5DJIfedf4sKISXC
jxdXexB1mXmtjbDYgdmwYq8aUHhFlHDy59A64DY5KYtss9eUmHC4HJLR5NvIdMHN
b0wljLLglyNnB7BCpeuU6z52i/oFz/IWt3U7ZNB/Lqe/huM3799MX3LmDcATsl2+
62/Dv/jkwJXLehepsQ3V3QdHMVyXKdrjT7lmczk1puY4AB6hfq/Tvjzbmk/QKU4r
wnSx0WvbjlDiVn3nLYEIbXAzWYsLe7ge23s2lC5GvDM65/mZ2iG/iGQTx+CKtgu3
GTJeruuV8ydNCtOrhOj0Y0DDd+im6YMFXz9tbUStxbPo0WU51Zr0rXp41lvZajNo
tGoBdlkmladGbs1ACohN4oeX03D6V1ucHuL42SRmohwIPyHR7k+S2/pSBAUIRq6B
gm+eui8QrqynsAC7eVXlYcAOKnEIbNEHNY9PCkJY+lCsurZ0qFMQvt8gqH/q779u
K8OB8fzcjmS4DDWPTkb0v6rYnOPsSdWX+pXS7T2mrTFlh0vLAFxYxtcEZNi/wyMP
EYdeBx/mfl7lgdZbo7E52MzIqhqHs/rRoHHNIPog0Ic0LcBo8XvTiNQzg+XLkymT
Vlp8IEANAphVPq4FAxCwmg0PnJ4elGctINORDI4uLMSRogHMdtHF9s4E+kK6+jed
YtH3sBujHCKO0COLaPonXF4PDCZWmsBPU0KefebKqnAnmYFp4EAXCkNwWR29F8vo
948grR9JJWALW1SjBnrFYA7NX9HQb7l66sg4yqiurzqEJLnR8yqh7dQQKgtBm+gm
/uWt5NG0JWXW0DrSW/mI4dzpv5raKdT4E498Q++PybPMJf63iJQFsso1RqM0cPId
HNxNJhURvv4c7bkhf2pinSFjPG3csIfsbMFd5wkUGhk82bvBFNm90x2W7sZ16LMI
D75yIcS3ycbOP0zCg7KaICB0lwoBbl42Xil56kg74gHVk+bjQo83+o83gl7qLgIC
7dQejM2KRP44/C2G+19cfi8lSvbDi9whn97pVmrwqUChDN32rM841hNjvMwz19BC
Hpee3ve7OTcpDyNyRzt4svMfDy/Inuofbbqv/eehNiGhBbg6FuUfMlEvlwuPzOM4
vLoWdB+sZ7qvBL+hDFuwRqJ68HivJSEwiHJYzeIBUJPcLbZ1nZ295Z2z6+/K4bZA
+R8T6HFVNxs4mb+tiBs11og/XalZ674PO8BpvShGd7LleiN25ZR42APh7a+458cv
Cbjcwlc0HuAUncqfKIc0mY4nG6AEhVUTtgiA2Mdsz7thWJs35y0zZiz254CBnaRk
Q8erBddYWo4SyDOIhf29bU8bklzdog2/T4NOboBaMwqdw5YSfTBKyScG7MhKlBTP
NcASgKO2warH8WzymBMlkI8xTMbt8dpWY1gH9TjhUllpshWwNz7Jnfz5DviLjCMd
vjsyox6WqRz7uZp8Baejw9IW79rftczyO7JuA6DJ6aRnoPWXW2a7gynwohfHPglj
yJXkE3auQ+izTLZdeLbXbJC4z+9PXjcG3MOZapyI6SfAgAiMXL61MuGwDmJcZF8O
7ASeOtTx8X9Qx9KGMOSO9Zs2mru6TvdfUpVAHP9PAU5PQXuGz/cbC1LCwQmgqkK9
HqKeFdWY3u3zt/wJyzYq6DaKtqiXGzNU3Z1o1Kt3e3KDkd5iuhVOAkZgs3oqytYB
ySBkaT9Ym8imGhTgOhpNNcoseijaOdJwx7imDwUE69VOpvKKagrYOrsFwiDfddk3
jqfIGMZLkmnE4tx7NOErdc8bONhS4Eh95e123IuuZ3XDCFrUMqEvhezW9y83Qi0J
CXXXrztZzflvqr3hmyPQC+zUyeDqAdKDjUeC4BOSA7jXqOVpQESlqUiU/LKymV9e
TiFOrAc+OcynnSsPoqMZ5BQgqmbA6+9q1YkezDkM4jIDnrpG6o5geBDvNwnmYbe5
eFmH/mBKnmysnDujPCjbPaGrNgtug/Djotl7QhI1VQ+ZBotHsic2QvJy7jdC5MjI
tRiSFJgs8lCpK+tirndjgKhLQKTQ3ZTE7Tu/9Cm9p19tgMiGQ3PUinJ0ZCaa0c4h
5HVd7RJOCVy5cNsuMg5qPL3J6+86bkDqblTIZ7p8bV4HoSs3aR2P5IDhP+C/R7r1
+kBUE4e+oVQ0L5sHA2ef3RmCS3VBfcutP1aaJHtkG5FiY0ErIYu8zSMtjYa//YP9
wb6iASqcj2YwZk3jdR/rYQS3mPiZiDAmvTlvTsgY+0TV6UW85E8MSx728SYqJcYk
sy9RqZam70fpq1lPyiUY6RuFbHSGYeqr/unSYtIXe5zoCnQCILNXsr8AGzVb9QqP
FoJpTAbjKHjqXIg423YMSv2qvRbqjw9F4jk6nJrU3xzVNlLV2b+alxGgXc7LkFIw
nVDLqVtwtOh8UuUmoLKNdfJzK0oH/9UuP9JZzrHkGjSCLrHeDN615YYo6ZZ5+ZjC
eocY3eWnFnSaY7kF/vx3wV+IXgMAaoDAmVj8hUgldRQwyVXYTrJYXkvZozQQK5LN
MIBMkhHfqiCp7HbIKpIbEwdIWKz5QhK2Eyl7dGFlzZ9KxPN45gUojbMx0pWTBVMb
K62Wjdbk0AT12qLiuHuXHj0TcTxtd2l6/M9mcGWSpAapiU6ubBdWMNfhOChYh0nm
MzuKdqHrVpoaSPMEej7FpezcIA0FWaqtIxdsw82MLpjbPES5u7CjnOUf/2pSg3dV
DM5zWdyE2VJtHVAb9vFidqS/wNWWXddarsYRa7To67e2omC7npQxEuHkCqbBLvOn
Pmlvdncz+NMKUiYbL5xJ1X3AUjLZkdEE/G0X8i90L4mwzzOd+q1yIm6InPJyrDbs
A/N6Ny6lXXIz1IwoL+NlcGJaTVFexeeuOBFuAbHFEsvIHvbRIJNj05EaS5Zqwnzc
L3OZYNZzZCkybEzwhtvS2CU8Y8IUEsn7C/HoQCZcKbyOJV1C6N3pIQtDJGI4p5O/
LdTC93vlibUq9AVVw+GoxnQo+wDBooN241MqfWiKZLQGVrzj2KM7+nIOJRcXJ7nW
uwWQHoRCfVrKyQ5TiNoBicsFEV4Cco3vjktn5daHMvgSQn2KOpTqWD8ytsE2/U2a
Hc2VZKSiYrbiVklVI9MYQ4dmQtvvVhnQeiCpprZTw5BdepqHwc68B/WXcdnFr7LF
Svpu5uOh3L+HT2cFyh4VqYnlRXVZq+FZReatZGgjRTXRYT0kF2qWMsn5Mv9d50kx
DMfLHYfF3smBYB4sTiJc87NXzaKPtt6eKLdZAjapiGle1Vh0P0CtYuA31QAcaiic
40zozfFvMVU+4jEetF1v+VnHvLuZP1pB76H45qoajJNCw9Z1saNsqzsGC2TOb4zn
81R/pIBmpeW+wVOxAcmo2jsmY8ni1nGRe5F38YQ3jFHLbxwPT0pUF/XoTwuRGdrJ
09PzQV3qpuPigw7te5LCyEj920OzAm5jsIJp6VEYXTZ4sUrOUIVyVinDn+SvTVMp
ZTvfIXBOBqdCzSxtfRyMPHq18kjGeTGPUosu2PKDILsvcBCJTilmzitVPFjSm7A6
LhDisA8EQk2Hc6vw1Fi/w2uprVLniyK15So530LRihzoSK2Qs4GWfW8dU6Q4aTYU
aQhcbFzvPbCk7prTfAM8OOJzapdfCLsQ0DBD87Hu5XD67a3v5Q5K3i9GPTgxqu7Y
uhgnjBn5n1qTBrT68LngjatpZLYBf6sMvLekVv4alLcTNkQh235PTGpbd2nthpah
u5+CvhEsqvylVGtgl90OHQLVUgygxwD7XzambiVD7u1tfIkJXgds6IX+NUnZERvz
e/mlXyvMhvbU2OSoqU5fhrWmfy9As9EdnJsOnviaVhjpqlF6H85B9Mc/oZNxN+S3
5ztB5cNhQakex5spkbMy+fcy2WeoWe8v7K+Es5e/oIf5Y9Yo+C8BDzfOl+yeNer3
68OJVqF0IMFtLcJfA6PGonqXXltS5Nv4SNZPcLs6fJnAKz4PFwLbYSo4obmc4KUM
oi66X6V6VNUQ4QKMm0fcLe8lsz/y8c9nKhLuq516xJk+4L2hpp2w/Wzsjxn8wT1z
m+KKtlIfbm4QlL+xiodyJAx7rf2W9G0K30zOenDNILj4Xfkj5nI0tm7pEpeKfq6R
V62z+i1i9k6lyzrYJ/mbZKpP6doT8h4Cwr7dLOmTJvojDYnkLXvwHseDbJccDpBv
iPxUtSQ9FMsyjfPaBqvtIh92z2+bv+z8T7TkjWmD9fsIpV+wsX5nxuzvJsuqJHWR
LEMXijAQGHczthTQMin6SGShXSLXjOg83+wB3FrS/Wp6PyXXzpZgew0OtalXvizB
zdWEEmYcQesdVuABKtlvc3tL4/kkH15Jpcz79BV9ENB0IiGjyBQSGqw4hdmNRf2g
5+DduRa6Q7lkMEJz2xFKvh6UKSgKwY5c+LPzlHU6xwXFAod4nQ8Y5DNNeJjs/2Ss
gd09Skfd4C7LlFkDVH8SebXOa++rdK5ThOBRilRtuk5ZYjgbeHSFv7fUuphOr9HL
69fUP0UVqtuZot5txrfPiJNQ4aeZuXrvbuaxel97l+eymqxmH26OfEmEhYlhRDLN
Y5YyBQH/hT/uiizIHpueLVq/wCjsf9t3DSM05UQCOyxE74eCji2YhWjr1CiKVdMT
66FnX92DJAwNTVd6qAbrFr4sXd0PdIf0JS/KRPBNuUH8Hr8rB4MT6dIcPsXikBWE
mT+9aT7Ox+2I45UYWLZ+YmSY1DaE5ovG/l+bxoUrBIMIIAVEPVUFooAbNnLJJQYO
M1hPVaSUImLvmpfRm63HCP8lXfTgG8mywWd4spXLWaPubOCbNkPJqnVQg463V5y5
vRtyor/uMmMHm48OJ9xIMXlUxTP/alQ1wQ7RHIYFYe1mqgArj6pKToOt4DyduuO9
eh2m4wvG3CdbL6dZQiQbgIHmdW6UPSPWTWooIinGgJ7op6VgpO6vzXyaqgnHypQ0
YpG62lFEMPgh1rbw2U0rJAYjdgZb2XsvG3RJHx5LfSQ53gFrANuQhaRJg24Z0aOJ
RLBTHdzkHMTJtdAoUYKh9eKnZBLCYaql/YjywiKgE1Pm1EoywJ5rz9gNF4sv3OEW
YsfjWWcIaMbOOXYpcirBin/fiklTTxJbrLSKt+JP0gtYVFTMdGa4LFa2pd1yWz4R
QRGgzoOSoMM0OiRWeck+ymmUJ3utxKQ99/SY8ef6nLkIqtYRW+anKjAdpiPP502a
hh28RydNauhTqv2mHL7zhAj+QoWa7S3e65MotDTPgeU/X53ZYfqqbBJt/c70rKYX
O40vE/GBlcgiss0T5bEyI+TeMWqj5R1Yx9u74k9SApxcdy+jE6LqOL5qbHntqujz
q3OOsge0BVxMP+4H8wyAP5rON6A2g3IQ/brE4i/wcR6Qk2QkPn5ZgyllEOK+q/+2
/QUKGhwpoaAmlXeTKP4RZKAOaPqj+EjCi2WuPfJWxkV6mlvI7jvCPhVItKC3ccoI
4GpIPllreNVyNLMIg/cGCkTfJi4IbEoKegjqen9xyq/1U0sTtd/UW79W9Vn0i4to
PWBtzifCxf+1PwTSu+5ocPWushrkUv+z2N0mPijgNwV2uT/Yrc7WKLaoapBlX+Ae
0Hn8TGM+DMCzE2ipuS/QVUwjHlV5VOAcBTegFIXdpiMTisFk9yduwcehk6YvinYT
i1s+G411Eu4m7MY+ebEcKFbJkX/uCJo3nytLQXun9jA6vGJ5SR0ow4uDpBE9cJba
vqmPdhEzQohZPSznl+ZNSNt+aKuX/jlN45TabZ3fSSZTsFb6TP+jfrnbdNvs0zmI
EY3vnltS2CBN4RXL/DxNXvL1Os9ByqSvokzcAbn3ctQDS5L+uXSg715ZcfIoOpW7
mxmklNKW6ltY0BaIgMJ4haVLkpYw1v5I+tgbb2OpOF+rsH5ui1Eqtt6KTno5MRvT
MXEtq1WwABvi5gyd98lA26tEeeQHrrQAUZfOOSe8pWTuOs5HspHjqeWNcZS4UMKT
fq3Mssk4C4NvOx+EWhaASP2aMu66uDn5/ruyIduVV95TTKK+FL3In6RL+fSIzNBz
Rq6teWZlkz8zvVA7V1hEEfdsCG+uN7EhKetK7fBtplH0pgeD/nKpJYUTShyuLydK
33tIg8moQ+1CDBNrMHLv3q7q1E0k/K1whtJnEHNx6vulE/LSXpyqsANj/kiguiTJ
G1U1nD3KsFO038j5wB3y7IxuDI54bnoCwGXSjWoNqfq4Cq+wEZ44fp58a4qOh74K
s+gLK9pYdSsz8jHCtmVWWeJqCOsC8SarkxC1CBkho9XTXLEf7uMRVDzArzcyI1CQ
bTtOqqw1SSa1JXbsk9VpLIP9bSy3RiLpqVNXivyIr0f+qBneA+nQY5lI3w/SHiYN
dgkzLQExde11C6VR3eVsD5EyDucumJfW/34nwXGV1XLZxupd+sKdhRCJqU/nlRZ7
59xJ2EKl8EOJvMms2hH+MEpbFzPq/qwslgQ3zf88+lV9OPfux2gFspxOdWnat9CY
IeNNCHUdN3kHgqnKnDRRvYsCsUwZNqYp+YU0QMWaUxWIAtbb8gLgMQsqb8yV9Ffd
KUibN3sjASC8sl0/tk01NTCXyIEdOlZSHUr2qklHLIvNdAPWjhEcamGil+gSUc+H
CMkuhz6fSTy2tPGuY/LfO1+24A1fb2Hu0+14p+CbjX2iwmtks/HdeU7IWghGQTVf
Ws6vdkl1wzJ39SrBy6R3d6JnfTsmp4AfOBurUBc5hUrspDOvWVYV2pPpL9mnEnd3
aNy0RHWC92CIuYCBYiwglF2xeAdbbZUUJXShaQ0xAYZdTZBkIMu4OBzT4hoYDCLQ
Zp/ek4t4/OlcC1tthrYon1VDDfgI5Pp+a5JKkjQJuzIAfH3dhsEI7PsDsZ1SuPN0
epPsJZA4lbzeDqAB63mZfP8cQYMqoojCNjmBb84USgeKngYM9sHegomXzv+4une8
lavpdKrtNJ8WTrgeNBTf/eiBSY98tJYzOvesmJ4h5BF9FcyjhlxViKz9LE0/BtfH
5T0IGjDE7nGFie2mImFk9Q/SKQHqiGhWg9+rMC82BLw52YXaQ0eytKvnQnU+DnJe
TtGXH7mpEKAhJeiUOkIi3uxz/jDB/9iqpoBSHIvF4vSee+JHa/zCMX5P8B8pYShV
b+s2Jx18qajr+EPEDpofXrgAAJ3he+9XCO6swX3g6N8vU3PDCYAJwJoehDdmJFV8
QqZ7ChoTpOqHAKVstYfAZMGefir7pGnlSfeU7oW/g1cyJuXO0e2vTYJR7yiLWCh4
gMR351jdiF0ZXIOw0QY6DQ7XUXnJYFz6U1H5hMBox0YyLIw4QAXSHuTyIBbjn/m4
F0ZHciqTIVAy8QrfDAx5fAszVdhBAH3Dd8y9QEWQJiagYpiNDR5cxgh/+GW3ImYM
f6iRNG3ktzRUH3hFD54FtnWgKZfSnsWoQwl1YaSHmFok4E1oVsTKRy3TupgRSvrM
lVT4FSrnfL8D84Wdpsh5LoKlFTAP5sN13GBNKkU3c+U4+APpl3W81fwST62V7nXv
wGGON3MQrBwwrbO8im0kS3n/1k7e6CL54OrBiBGE1V3P1VqrlaxCqTOeNbbhue8k
v1E7RRLXl5+xj3Vb5z9/+uFmcirmDh+kL1ypDv9daiWnXTzAmIa36f+Yqx+W8GAi
ZOto9MmWajHqJPfGEtyvR0611KEV1YYwX5O/wfgn1Gob76urZkqe63d3TfXJGzuj
ZJAEiNmrvqiZsjrlOyxPz07rHxrB7ZssEXhtmV8CTs5QHESISVnmy/nMGwsqWGdh
ifplXCAGh7/rmfQ0QTmN6+HfmomJHGHnjIz/3k2+dMxiKs8jH5WyPLzqly2Kzcxv
PO0clKhRTPF8/00G6DDpNRvyG9yP1O8/69a4UD1jDfbUp7Jd7sgpdS2ZQ+4hJQNi
iNTgx1V0bWl3CHO2/YxvsU19TRH8EBoryOqXlR+3dNPpmRswKCm9e5ZU6wh9i36L
YSUmdHMVzbgtUH5jFSJ8EOIqcvhZyfzbxCk3gLDdIDVEEfsQXJep/WMK+hi6Opb4
Mv5nwtBKhZdafrgotUU7+XpbHWR+7ywFuNpLj4CgcVCxz7fRvrsesVihscxnvXH5
wEptcMlMYSdI2S9YGtSlzkHVwh4w/LhnkMD+/Sox8k4N22AIEppSqxU3F7MaWqlA
b+InD4N6iQKz3BCkwWTWtdHYDXX4EBSOzOfsvjnP4FePEeq+vNL/rgsXdKyN+th0
8xbvwqgHHCj05kY8I4mrxDNzVeILr0mz5T2rwUeac/Ye6LdSAKpbQcpiHZYUHXkF
tTpjoqhsDZ30CGafpO1+dmCo9gzlbaEZ5n8yVmA02uVHUB5KDX5Q96KiWF+PcPPG
wgFMSxGPDf4ZftBDN4I06Lf0r0eEeiep3p6oh/or0nUVzKR1QkQ4NfGMV47iO0/h
E+H6qWWgDM6O0K2XfIFMOWrB7M8vDMs7xz05wKj62RyrQXS+lCMPMKTECad9Ktgd
BWFqYr4xq8Vpego6V1pS6R7lGJZZFSE2cqmHJaJnIYrRjo8lbU6wv4GIatrxHZEG
Q30rcsu1ysnvK9CA0BeNpOLH1DfKvQmbSoetvZQZ2wz1C4eqqChEXAAX+Wos48Z2
HC1InlKNYkIvoRizU8pc28bJOJ027JsxeHC3IfEo23ut9thYn1Kb5E9jIkLo7K9K
AR92B4rl6lpeXy0PS/DFeQb1Ya23ACVhdaP/6VsIBas7Jfmrn58BCPS2UCVtaJQH
2qbXLex4aYZCFKGx5nLg+kJofS/uEOC/fTOhuA8OWCPfnxA2sw0BwG86AjIcz48z
pmZFaCVwBF8s8gVDsRWVNuqL4uvW1M1QcQGcDW5LYnaQ2eKxVSPCwgQ/t1r83O6B
32r3rQTdrxVK7kSr/NMYDwtCL03zJ6GYfZqPbW8KbHwidpPaH6OQFhNkQSaTUUPL
StjPxTOZ9IhaYQHlNrPvgSOClLazXL50DgMeSqrj6M3IWQkO+tnceWZ0X3VyKSOz
U92NZpy74WHswf/aLdsuqxAfVLwVPhrNBRt436kK1oBdzl5w29XKDLQGjtMjWKBR
q98JbJyJO/Jch51gnGxNGKGDKLMV0vBOl0WU+31hQeVclIP/cuBm7k5TzqICnTqV
NHZvIQ3UpyduThC3OLxneRowZ3/xMLs5ouIhkjBqrm1vbw7+JwoTGOTZcfppCyyG
dyj5bBxFEwq5hnss6FYuQUMII8T0EXDvMtXwRDqROfQe2/KGatRvxSal2EbQVJL0
hg0hWYbtO1Qzy51bB2Z7mxStDeUjBoCHTPGvu9iwNZRo40zPFsS2vgFh9kvnbjef
zCsaZn3/Rk3M0dhgUp2dFuWnqbqL0guntEeAq1kH7+4w52UrL2gLrgH97osQc4Ms
lYFQe8/24LqoVoJFWo/UW4j92LQa56yQHtDNlbAkVBgrclqoFLeeisBsrM+EtDSo
Wy6ZvwJoIwlacimyd+Bmljgs8ALlonFKENaQ+jJ9OQB86MUg5cSSmseeHF2lneeB
q8q9dQ6lCN9/f6gsjIx2OzElxYgHIC+cXcmsK4Brll/xA3eptkScbZsXNJ8rmt/n
3eob0u7p/79DMDe9FyV4iZvL4Fstc0QZY719+RmfvFXJU/Dryy9Zm0M3LTPmrQSQ
/cKPjo+RcfYS+7bWFKvEeUNRFtpVHilO5CkBViFHvuTN+i5HPMuPJCK8JzO61oPy
emZwV9rXoUrw5BILDqn4c2bRcBuBZfuYu35f14MwFm7DprvnuHhNw85q9EVDFheu
5ge8x9+9OjcYtOVyFYs4/y9/D13vlcYeEIfSl+ZZwIP4kRh6+UNeUiv6IsT9zaOM
7BvjSHpjgVVEMMX/qjzZtgVNNZytaSR2OJnxYayUTGRcz7SMTQeK0TS6zjd2GwwU
KFGKUuN9QpGUAdd5B8hwajJQQrXltFnwFbQqwEZ1IJiApp4zN9tLBZ4twbbtJs9v
qOE3XABAoFl8ryFkSmg/6H/1llrKFkKgjljlCq/xS2+PL+LtV/oDJaghEOQIe5bB
RV0UANiBfvc4s4Ofy9YFbnoJJP4r9clvAahGHSAh9tLj4mrjQaRH3boIZyJYFs6A
GWr9fvOxOt1e+CfK5XwZbr9OHvNqjlZp01LmB/A+MGHL6l6nYjID/c3HNtg5HSfJ
JoHy4qKkTkGhAC3+OK1Qklf0LL1zG4p8SuE0/uuwe3S4N7OTs35216qPCS85iTUy
Kxe1xHAkc+vO4fEyystXVpmsX53bXPQlC0hIz7hQcPYeTLqen6dzD6cqcyvh0CfS
Irydy1ZSeBduISlN+D02gLocXOHqTnKBrBWDQBY7MquT4wT32NvDX2ONOG/JLiCM
IuSmxWdw2UqcusGW1n0Sc8HqdbA6fU1YaTTisx5AwJO+moqvoSqBkrI8Jg6a2k3e
F3MODo3i+GZZUHZsLsEVKGL2waJ3U8ZET8yQMFrj7D06seq6cRGvWQceebSrgtTN
DSSk1JTBiOaqKjZ7poxibhiljRfD5Ah/wDhge7AbGBkTv+fd7sWWqiH8V452bllg
FJCx8qSpdUUMevkElme12E4VdwPZ2qqKRRmUebGUXTpmsYmxOaYEBNBbnz4pPUYR
0RsvTfjj5cSfnLJOpPVqv+72OVOcT+zlPKetZhcA6LwE2bz0l5+NBKKK7A8bb8Ys
kJhfsxCrL9pdd2nE21oAcBGdOSdxcze0yRvupQR5a1FtPm16ayfmVuqR52jxb+ut
M0NHQmBGiyp4UnQDDLZ8yHmNEAtpnKmifpkqJNRiE3znLzWh4ZoU+7ALLcOUmxgk
WD60cCiGOEpUTpTmSQ4ZXUqwHi4g+sJllKWfQR8TeSDpeki7nIhJIHFI00eKnXMX
Ux3v+fzW54qy4/xW69oXz0Xphm8WevL/piaazG8kNckxTB2v9vf5/gWW2jPY3bsR
pia29bahDUudvs2Xz65q27s/nu6ge5RPHqSjkY1Uknk7TZWVzcd11hB2RdOokSSz
VNi5PKvpSmxt3FPlkX9VsZFzWtK5KUUZhAfqp2Fq+vTFnGhzbdhzfNq7wHJ2KFXf
Ky2TD8UA9RufemHFBzkvdWTgq8EZp+R3TG2E/jSD1OLOm1UUZnc1tctQAv+Jo2N6
cdxcUPIt9Hwdql8zy5Ehwz35X16RtcU4y2OpQ/j6lvOEhdON6FStg06d2SuAZAVe
hMU8XA5b933hw2qyvmBQKu/yic2NUZsHDN7rhu/bpVRFsu1EYLGa+ZDhSZ1gFdVY
mg9MjiFngMy7oEb97CersW2K2Mm47M4g/gux1a4Jhe6w3bRZifTvmGgGMo+XoRY1
MKmrlVPcCeSUKpsep/bHWAwmHUoHw+uxwSBB8wbAbFZOVJ8iuEPlldvB+a4mZ/4A
Bef9MNYxPp+lH1uCKL4AIq5GZMvJnvrGoGcMoUzdaWErGl5ykV9XGKaIxaesAgBR
sO+kyw584zs9yG/uNmweEdA0JWM/AxL8NwWp3h3xrI9g1lImO5Oo4ia2bwmPrbhc
o01IgQM37zTC4QHgdMk9uZsjEQwD0+jAJQz8MXACyRB4HQCOFXJaKcjGucqaWR6u
ENzD3EqVQkleP40GwqQ7qj0xxbxSzUiLmHU+vEwQ/xR0mugvxW1CpGWkPAswZbgW
1b4h75iFbHIsXTXsPFrAlCaASjSmkOVwMGP8UMxTNQJeHj2n6PWd7VMMbrT5VGoC
YQ7+QSL+BtdR7uZnHjfA7benC09WrAijlgrH9Edp2TuAGHDt1Xy1/oP2agkNAsYN
OxbXuksOuiFYuU/LgH7gkBtcUqMllwHJvlPVM1T4/veScqm5Ct4OhE+kOuZ+r4Vm
ssklh4Am+XXsmWwd2QYfzjKAn/eagOOMp9GHrDnzAkTiam7rg+kDC5fWW4K5MqRH
3CwsSHfGzJa/Tz5cFExK1+uJ1gfZx+nKdIOGh5txiSIRoEKH1+Cs9TYms4WwZDTf
UJI1qqaIaaIguOAxS+XXltA1B7EImGtfJ5evUvW/h323omIM64oH2H/WLWunODYy
Camr9/NsbHgNLqo4KdCPLQ1xB+4FsJPcW6PTAsqaThcq96kba27GdvhzUe2AC7dY
Qrd8is92cIquFazj5uYVlX8Jx7m3SwA4FkhKmPe5B/v8tDkPKF3RwgsALS29niYj
KFEbXBgg7EZHH1R6glsVTVitm6q8iXTtsTcq29CD9ZYIfQvtTUoyz76wzSWA/85e
P3weowTmV0sstE5axKbRdC/FMWqp+fgfBbCtKuPpPUS8/qAdc4n2NLLrVMgcWjbW
LI1jan1769kUbqOzgHkfSE/0PLV10Nnj4IIUV7V/qLoFNczSwLCtqXqsILKflmaA
ZvxvnpmkADuGYY6YsH2PHF/ZeMRDNxhiG7IS42VPrazdXbyQyB5nDBMGxejSj4WR
3VvIF3Ov7qWPcCCkudsuTNd9YuYBMZEOfvB6zESjg7V+40ydPv3avXVFMLm2H4dv
BoQV/jWTk5382IAR1cTbFPu1cI3VeTWUXpWqgoiQqmKx8GsZ9kwqVW0shdUh9550
Z0Kf7fEw8og1P80+7zuClIWGh7yY/IuHY8udqKAIQ56ZaXEF9XUQ3ajsCr/0Efdq
QfQPg7vlnpxHu3ZNCMK1rPWhySkT2a6FnJki9cVdA5MN7fKBBX2cAoPTbznVo5UZ
k9yv6QQbpKB0y+ImfdONaQliXBMmutp4EfugeMAP5jAbVxzY6w0W9jvzU0o6omma
i7Nf18P2gTaTnX0PlMqEsg3cwHUDw7CXjqOdCZBGuRJZdJnbuDN5nHlmfGtaGYkc
rZjwLqQSI+SmjaXrlL/zhUq89/PZ+D33T4MdEgrIPs1mrFbYjrGESn5d+PGz3+GZ
emNPLPbXygLguGeBRWV51ADibJqykSJc5t0nVMGUzStLv5PmeuPbC6LkrViK33Vj
hfSgVWxhK85f81F8etaBv8caywYXFbgF3ZR8ajDr7bfGmnkHyqbKVD/j/b5Hty3/
IYatTbjn467HU2EsUkqPYLjTw84jhgpyqQKSZfxUVE0LoGL5AKtaSb5Q1KMaSgb6
JQ52FI+Whwsm/uvVX48RR8IQiHCI3GmxiiJBfXs9vx5sPsDPyAyqt+5upau/T1Hk
UoayTI75zy0kCBB97+slQcjAEjYYbHKA/OKE0Y+l4lgebRrBHR2awO3iEfB5qnO5
RyjEjmAp9vtyg2/7mKXjNKhMuXGGK8uwVtdJYhkrj6lKqSl0ucaxiy2f9xYqt/OZ
gOaHZtZJV9xK9QMMIxrnN9TAEfVIUJFN4sY37pdI/USduZc4B7Z23b3RsBG/tnZ6
uMHYruUceosyN/guqif2yvOCmd2aRffKsJb74zoj43Gi/m9hl3T0HkzmExHOeKiY
V9JDPLGOoJKii1Uk81t5eU8jeJhQzixE2ODvsAUXjT97/aV72RAnYaLv/KjjUGq6
a1EQVLNbGhFIeNDDtPhPC92wHF+tSTdOizIx4Et3njnOQq/XAEko0tl9QcruEvKB
8IPxpqjY6L0QUmCw2nYZjnlI4etYKcJE3IqOkbtUYUfmympTCsL5bfNVYa1nv91y
9iBP294s8CcsqRtyeNe32Jxka0v8NlWJjzkN+Xh3pxhJYtagzmeE0dWv6wbdoJBn
G5M0RKtqGff1sE5m+gKon97b9IHCV1594ia/Oy/bh7HQwlZ65lI8wpmJjHL28LsT
ZFl+CYwrRSMoTtguhdsPGz3/6rxrljz5ka4yAMwUnOxLFX8fMx0TFfChwC8XCH3D
CYjL6O4xeDaw59iwYs2q6xxEOPwbNX/AfZJZiSnam3bv8y2H/s7O8A+BpHN8+wsE
PIDHxh8nsu/OTh+FXoT1W4nDP6Cty1NucCECrPMFYY6teQlOhKsxvgMJ9rWgeiUK
sJuLTaSUCj2NGYBxzTucNkqmuUGzrglTDk3SMfCUkSeuF9t206eAEvy09yaiIEEX
6xeLSKm2fC9voaDJOg+Svjwv70ZAF/9b/sfkihT/3O2fg9euLJqO66lv2NJUwvPZ
z2Atq2aRdPcnbOLuHBZoZbq9h+t7FeeFC9NfFVF/SDz9TFhtIavb3NyJAyoKcAjm
phF/kZFsH5KXe2Iz7x0SdLiv9VVNB8xLviTkV/g8U2L6ifxBSb1E1JSi0E8Xqghc
/cavMCNA6i2KxWr3ncO/JM5vA4/mR0J2yLTGJOZn1QifEjFRmA1YfFYFNKNm3XX2
8fL1YdH9di3jlnC6EGpFfWaCUTywUZiVFEQL/gAMfmhEWAm3R3844yK/FPccxW65
cEJgAJ/JIPVejjd2Q2FryPT1fRVaE62cg/DmsjU67WC3AEA1MwKH5ImuKW/rZvHc
BFSb/BopxbVBac8pvNUwPY7SCN1F/vwECMplq/nzv6LKL5cj5DAIpguzAKuDZLl6
gGKxcv5um2xPR29SktB6jGXn0DYxMVHqCGAqbmBUJHJj5emmK1vNzTOiaFX1lSAa
Z08KABK0ldI9TCdRis2M04ji2cH2qdNjPkDqey+ZoVmJbeUxTXHEznFIps+rmDOY
5bVH88H+WQm40cYPNynSJq2fsaBh5WsPuFNuTxg7xjdUf3oTPrhlkZ6TTijAp3zE
p93zx6lSPBY0ZGAamkhgBHKxbMzcdOL7d7RppG/ZjPNaVsEz8ur9yX8v4CXiB1TW
l+sQDvuEvlcsa5j+IT9sLE1ScLnDOaDYALcBYDm88rW9MGaNiI+I6I7p9eea+teh
1l29sMtnY/nhl9OL7PE0LXnCpMBQnbEbNHZwqZWXKPcUQegnhaugj5aFByQ+i+5a
cYggUSBuX49ZizLE8lPFpOU/If3fX02zW4nRPWkOxVc2+4SIsKKaw6GmbGU33QU2
eFNLz7JLG2kThiEjSPfQcoU6nzANA6gAzojh/M2te6oSg9VqQD0zhNp/eXNEGymZ
VuPwLPlra+P08ZCQoPgd70Efj5YDxg9/bymDm+4LQu/T+sPkse2dk+cgw7Zd7Z2R
y3c21IDO0QrkyGBih2QTTqIU5Oovjb8QpPTcJIcmR64avoqj3KLgB1t5lNnH6x3+
iT/oABCdtsD7orQ0YysHPKpY8PVJYnibl4Y8NRcQHZkiyXajx/0/szFqjuAnLWFv
S+z/nnRK7SdSHtT6ICB3Zd9SKvlJ2LLZW+9UPq3J850bSEjX45b0GJXfK8uDCPWt
RewFy9oNTTlsrYwtfBgTDtZ1SFMqU324icqclz431E4m9JshLp3gHpdNM3PNF+HF
iKWrApk4BFrJsRQnJ94DjqaN3RO1ZwcUwcBitAyIYfYvuvIEYUwX9np37sGy493+
A+kn0dRXg+8GvBiQUoeAUybb4A0klMi2lcFflrbltc9sumZid5B2suRDx/uVoE8w
4gVsq1CLujDhu8vFz49doqJhOBFc+tj6/hctNRv+/TU3b/j0MaVOSXqKvH/tsbBL
WBRJ0YBf0w2WAXqK/buGJPYW3mQi7LA19/oX5DonmLo1WKxS4ZlqZ2fXoQPTgVb9
P6eVSbcjSs1+FetKJiA8qrkAscnvqkMAzANwpB1XC4bwgwbkvJo6rwBC9LXPgz7W
xWPegQqtkN/HHqtOXY7UtJkN6yue/cFQb6LwulhTNtFIpfMhHYSjzOGJZ9r2uKQ5
5ZHYsA4m+hhw3/liXB+arIO6Bd1UPlL0Rd81SFfvVYDaPLbWiAEVdoROHm57Gqgs
s7OJuRgEEFCa1eGXVBdKrMG3mvMJP+p9r+Ex47Z+vIZjGMLNKUMiaKqHW6Vn8fSF
iKNotCDS5XnPx3Zd/cBDkEyItrLeYtPUtKvG8/7HSWwGsHB3bR0GZPD8+prhyN9L
Dy2BHA2aNFTgwV41uCCuT9MxJNnycMleCXlX49b9TAr97Cg/V1U7Hz/pQCzZdGgO
GUlK5doS3gZEYqI0CYOMNjWVikWK4VUTYv1U43r0lUIv5T3ksxkm9fuxj+y+E5qX
94i1HGj6lAti/hhGkN+qJQ3vB1okuaS0JUoQXq0f+wTYiuvgmKj4cRE5hLG1P/Rh
uNKpLlHqzePEJSAhh2EeKkcuUsQc4nYunAydCH1VmfU0SBHgS7NA4+vDfntO5FKC
p7H6kWZCgF+YocyUOORAJ/MKmyp0UN4kAtSaxi8cGvpNA1l7fjbu8JbEPghNuecZ
tr9lNTmraWua1bdcux5Ly7/XbnsgKCWgRtE3WERhWfOqVmGck6spaAXEjaW1Ui38
ZQiSxmwIVCWIBnBNPPiB66bIIJYQshWn2gFxMd5IEoVke4n8kF5vpxmDii5hcttn
owjwlWAvmlAQVthebt4eIM2cI2+l+FymXtuL+6U9W04uEya7Dy71PcqIYo/hD0H8
7LnTLs+1FFJF/Tmi2JmUaqYTsXQ/7wdkH9Un1blIzBbB4D5dz1LIbo12fomDRTb2
qBjpNOXZ+p1nGiuLvc1O5nsh+b5oH8Z2G7LjIFo7eDYHgy8PsFL6+eF4zAc1oHHd
ZQSPAulz2n+EnO7DAvZl3v0pV6sMPZjqMGFU1OfnTDH9uViDyuedQk8EqEUUYUfa
jmnW1lAtL1YiL41hrzdcLs2egHOknRzp4nka0k/WNU79O1rC6Uz5aTM5BWCdNiNd
cCG5Lm3b31xeiJw2PubhKRKI6g3HM/9DDtGMSazV4JklFhsSWVTCAg+22zUdEvPa
oPMw8NomsF07MOAdryPEI/Gv9Vo/W4UHzTTu6I9bdrX1hWSfvqjPdTwvmHc+q3JU
LZkpqJa13EmL1vOb9D2MqFxGDGBSLPf3PNciR2e3d4caSCBPtXdHYJCn2MoiZV+I
8OsmwuukAjQ/mZXSJ1/R3AZzHAk4Q7HglkCv0SiDm0XJ6nN8iqTvPfKsr4xB4ihh
Dz5m4r8pne0GwwcT80/MYWvtF9BXaC5GYLEfxRBz3jNvGSJAuBW7xDHlpOl3FwNT
xkRggfDUKq+wvMvop9oeadBwt1yFHTS11x6Ue1Q+aRn2iZeVjOZxD3IG7Yt7zB3D
fUB3zQLPsSl2RQvP5wyUb7k8B0SAr78zNkVLp0I2NPgBW4nyC/tqDKiDR6WMfpJW
q+HfdSWPS/+N2o+D3Q19auRxGoLSX10KSQrTOWg4pSzlg+p3BW4tx7b4HcEgYlZi
xvqLQlCkTcnlX/4aG5XBLm5j5ozsfbW+KEqCX85YWPotte/OWPwurr4VzeXXXhNO
YMRuSFHSqfXjXQYOHbLwqJ7/Izk9b7WrTGYIIN75kjG9NviZn2pYnblzfm8ocuY3
KzX/fxKDG3zI+DqBrcaoKSt3ZA5CgsoxeJidJqEpZ7BwsudL1tIHMdG4pwHYCt0Z
faOZMpXG1p/VNBWVQYwiSYAEvjH5Pd+6hQhqafw/mpWdQaC604mcT9+XmNXtKSdR
vNMN+2sNsH48t2ngg87M0YJbkrfxYYJLLQOw2OGZc/zKMlviozaYkR4yVWYQZGpG
lVd4/Ra+y0acXadqKuXzom0LLPp/Vm2QmQkLNYUi7/ILoJTwP0XdI1bTyhhRijiS
ZikG0vPm1Rs8uuOyRmpRyUkZtv7hAwXskoyioMH4O4QrSzxV7bPk8AA3X74fxYeR
AF62DP4SJkvPMT6JDi1RcMtJ64INUBa9sg5uPa7Q+diFRsnEUF8rZiLY/B4ZT7kQ
o7jSG8kJYLKlN+xJ7/H5uj/p21JYDdksGVU5Wo13x+qtxQHzwnIVgeU3RfWWI4ph
kec6OxzjA/skr7uEkqHJ96mwbcjCbs3Zr9Fkr1xs7Cr5sfllvpMWY2hRZPePNSBc
Qx7htYxVwwf14dNA0RfPYee4fG7pgRBT731PLAR7tIfHtm+Z9zdVfapOro/lujD7
pUh7ewO8cu4Wpfjzro9lFgPLxpC68SSj8D0/1mVTEqvdgi8VjOtGUG3aeFH/KLyg
GE9vzHGeYQ+c1SKGNITHkJtrVo+fDjSXbiL4AjDzBvNOsu1dZMncyYmgM9jccnDr
7dJi2Si7S6ylg1EqJb/ptwkKQIiUY4b/5jrSen6JKKIJ/RR2KEgOz7d3dnUd9lP5
xfZF0k3YaOjQT3lpsva8df62Un6sNbjBxoUqjYN8pXny6HeoLohg+dEM33/aSUgl
s2CR0+MoAZK91mUloHH474s7SMyyyvWEQpIUsC3PrcoCqyevXduK/ckR4xRc4o6g
B6DUZYeQpYQWE6DyXXrz7b+89fFLc8zboqiZjAeBTAkClExFzsuYxeTfuezSQeZn
mXvS7OXgZynL1KY/7FVqmxulfqvBYPnUAIvr1RoxunvzoZXPK3jlWG5dTv/8gm41
R4/LW0ByXU0KNYEb66jY56rlnyGb3CPyoLRRak9g6JoUP5byilvqYwovJdqW7pGg
9g94ukUswBKqTQvaLI0sOmkWaOEnzn9Q7uo3zmUcIr8Lj3wMY2cjeTJoFmqpcEWJ
1E4dHIDeAyk3RVNmaSKYwWnJ9GeTPi6Z6DK8yj9r82YYFsUAAGxH8vkMf4051KfG
YaJhMatddGZOwcSkKFO7IeKUZii+UdMKcBK7WjAiSvv903G+OcIXScoKaFF2dYWn
CTvo6wHzGSEtlHrtf4VoKeQbzH4/YRoiEW5uhpkKiSJttS3BUrPCaCd2e4Qp8qGz
/fRIRxYUq0afnSPHkhghtif/e+A0vvM/nvhJfC6zxO6CRQdO+HBfSzkOoIaCEspH
FsLfEO/2P9XvPFyHEkwSaw/wGcWhVCRYOkcFb+/3eLM3rSxhaTIwSBhA5OMz//D5
ynWXjcLq0C8RMMf/bgh/+4+4H9gFBxTV0HWmoahHhtzZBrS5AMWK9qmGSD0Y9KxD
uXuv1VrgUnSAfDr45xPcnrrmO/mo0Fjy7+vWRZUWwSGV2tQqAW8lwCJ1V5T7qWRC
PxN67tEiR9J+7Rjl7zTkAhtFtME/4W4rgDJ9nnt8Z9hbgKbIqt+MqrMLzN0iX/X4
iOnllfFX9EEfK+SnansfxbvtZtZHpU0g8/sFlRpn+GBq7xblpaL79QlA6lg8PGRd
oawpgvtY7lH9EZviKz3NOGpJkWXJ528x3EunBpaKKUnwiM+MpDaedpu6rj/mKjzd
RHSwljV2XSIvibHE5senK8k32Kxh0MkpZMu5R5j0K7zfi8SB7lVCifDa2h2GQdA3
4vJzMfXYp2WzSI1eX+aWxkkOh7dXDHcbU0g3msnTJSJX2ESkQS4At6NwRYlKA2nx
QjJp91+ai4QIgQn554mQPTIFVhhqvUHQDwVcPAi66TQ8d+hSJkdT+YTvj6kzW8B+
GL2lYA25ptjCCquKfrItK3rGxFpkMv1Mlt8biea9qkCh7+ahZOE6c1hq+6O7HslL
dNHwKvMsmCKYHm9Hi7r6ttJlBkEYJdGT5A6tHLyn7qnhdDrYnXeu4Ha6GR/89MTm
6dnNmrnWw723Nlaqbv1tEp/8n5iRAf5yjla38hKawsIgIuWrEhRRuPvF5rk2lwpI
iS0nItBcHtJp0Ds9aZ3AY3tWQuJ2TTl93vzIupRh3iFa0qZFLdG7vozpp9aty747
67gtDF6qqQi5NjVhpvF0dvrL20E2rVfghXgwTptgD7+Y7Z3JpYk5VdTKcukHxZ1J
aJLXHq/3p61yz4SuL9nQynFtg2jTWX4UvUIcj/DPVnMVtWKi4PdJ+i9Gl0U/laWr
dKyyEMaSl4X8Mf4wiBoTJO037EEklxq5FftkuUHprFXB5MWmKBTaLJHRCr/tfQG7
TPvyp6AT0NR4xyyTmkdRw5WEqSOFfgLOIyVpeWaks67qhU346b1pkGi/ZTXdkrgm
1DDurae45f06IO5vZLpnuGE+hTlO7LE+NiwUTS4KvbScbi6hUQOG/8PUvaZzn04z
p+yTpUAf5NvFP7Z3YHmJqea2AtwDNtM4MWc4tw8psG6C+9jQD5Ne8fetpXSjPE6g
Svy5JytsNQUXCBXwL4XBxF59IINNlU24ZTHrp91VuYSI7TiL91E5bsbL50GCQQ5i
3eElXY6zgXZpZqJUEg5SWnyDimdI/r8whybPiU7p++hz4Ke2NKsIm0ByN3ujpave
sqyC3Nj0uHBbc8cELhkgtUsr+3VTyUAw29noLB743P79eF/LxhMuUWPttunFbHoB
xNx6HI0z/O66P+ETLgmuhzEIbVtyVNeKjaXeOq70XGUxDVcmGDATaJ/b+Yp8x5hC
44POKaZOb7D9Or/MMvxMznITYUGN1MP1XKsEspgDcbZJl6ThEduUwKfHyT05qkAS
HVW3LHHkoCd3JrPZJyoy/sDlVH5/g4bOFyIfkDomJOz1zNZhwR6XBBO017yjTyC4
cR9i+3EIAElTdPl0sR0tC/gvTxnq2cyw+PL+grwYr3+ZlvxQDFj4Z6U70mPrel6A
Qyx1xkBJNGPpKcdmcKD0lYrm1UEj1PHI0TL6ZO1bpoWXl6CUmbxZbnLWmUT/EhD2
BdWCLladbNAmpDKLXOn7YZ1uHRhW+2HhDkzJPLriGrq+WBPoHowMK7REDo1VzquB
f2DohsZl6NeMOhwPnSUydGXhHdOfzH1c5WZWS6awuxyVU7frUszQBB9P5ynw9vQM
kEau3G3aWakjBr0WW3bSKAi3gTuFWLFlugqass+O/L6b95Kx4PQ4VkBznElQPx+F
dHQ+2laR8r6MuaWIRueldQANMgtTbqzGq4sdUvTJ2Q1SxGldbwHDvc0v3nPgUhuQ
5/v+7EcvC2vQ5n+d9Z0Yf1MAVhmqX7zl5PSOuYFJnd5gIguQpWpVDncJkHzRXhlH
xxZReuGEAWyDEVCTjKkZEvYImaYPFcZj4auGHCA8igc75R/I73TJxEgbvaB2eUhk
v8pSJSPQ0mIQz5TisFHKeYUzT5X2VtsbGodXrocD/nvDj8zy43aodyZEYiIndl0a
ZiZGLb/xDGeH8yyGDfQ2xRlpY+GzsS/wLkfAWfGfRj5SXrEx5xBC4R0WR5tbXZaz
TqqufEyqjLMy7+1Fo3oNe7TmAIPfKhFgVtIHF6Q0OTZYkY2/ZeKfl98xmzFex84n
Oz6BUcr1qWCZu7+pHipjeRJI3fu/lEozT+53s3VPYZ3Q8oWBTTBn1oxQ2ReZ9pPH
uedPrJVQxVtetewdxX4sINAknCBVnUCAFPOFdVIeRr6nvrGehyravyl0GKKd3hm9
Rqsjp1jAXz+798S3oXEItjFCY0ob/XJ+LFfYCvvdmdHcs7isBOcyXrnSSt2d2DUb
Xj2/eQ0h7dF98V6zwj8TzItTGz6mpC3eN8cDFKrEKmdik3fhxlPU9qZeXCauvXyi
7/ZVELCZhOm8EGLEii8rJARC1BZiw/D+jxgQKi6g14sKtX+GLiK8fGJlDLWYsedn
/cImGPV1AzIMOB3GgNAVLvZcRdZG4f4Asmyz5ToR4xsdDSZ9qjQPt/Tz61PBJs/i
PJayxcENX8YH5sTRQVFXRsHvWo2xTdKDQMXoK1023IYDzrvM/E+PCWP92obNiTk2
LfO6Q4cZrcqHufw1bx7oQfN6ecjOo4D0+8CYFbBjtRcwrzPzcz80dghJb9ncRP6r
U1IJUAmSNLOg8uiDE90cn6CkvJ7bWh69uPRgN+pS20zrdN9tN+6m0ro6MQldPyyu
k/dbJ6o78r6uDBZ7zMPuwq/IOtlpkddFi4EFBxqAaERvaQwBn17q0NT+S4D6Q51g
Gm7iui8aYFZjiauL/E8VqaF7UpSC1F0xWpG0ovp5aPog9Tv5wkicPg+9edevejro
QPnj7nlUNA08qDIh6uF8ogokueYrVFtOUvAKrbGAamcccfjOgWkWjhUQkqBu6YFU
LIRQ2lkwHaXLj8qDt0LMkCrR1MpJqCZyvXrjH3aDPCdgHhYgm8TSmPkuZbdQqO4l
3J4l7COmRg7BjZXdsoTiUBegD0J2fQ6BlMaqhd0q3pAcgFH3tN0jeuZHR94cu7oX
FeJbA73gnd6GYpjrwj/I8kT+geaFmee2Q9OIP8kwrvFu+aZ8hLtdJSTmUcX3uQwh
1poI9dnbcoqNHNiiGFlHEf4uo2wPy6+zbQ4LwJUDqSicNPaSj/xjEBZYWL9LUqdR
v+8AFTP8XfnZfaIyEOAYKTyzUjsA93vuU0GGZDNrUSmd5kmXWuJjJQwuHEQ6Ov5Y
orB3am5T9jONz7KA3UHeWMO7ql25WjfQhKmIctqkRVn4ME8okQfBb4/maCuIcXVa
z9cPONhd4jpwSfI/RHfhmztv6sjE2LVx6RK7kMBetTF/reWCLUpSK0bZPHbxmSVK
PVjLpvKZe99kmituIUl6vYKPma+2RAqj3G1ogmA/XXAqBnJ2RGJESGTa/scnH6Fr
13uQ/fFQ6Li33ujHEsN1Jaatcnb3jKqtjGd9pTBsfTdd9DLj08ko45Oms7qQqmS4
j0bVuJujoqeqzjczAR8uz1uzBtkYmIVF5ICNOJM5ds5/efmfsxUqWXGhqgDtSj3N
6nOxezwhc+ZKoAQD5OsnHDFlD/sQ2Hq88vhtqcevig48t0twEqe0nvLZA+SxiL0l
uw0v2N3/TRnnfSaTxRuQpAebdEWoa0kXvKoEgsxOTFXJuVG38J8aTsTJ+1yv8SCW
fPIhhEQ3GVZXVDmXC/il4jSdpdC4U/sqy1VBKYNmZwn3bVO8eAoGd0t7lgPZnGkx
/H8kc59FCNxmKdXvpI6p1p08qqCXjW4zFtDbPUkAfVLGJtLX/JN68VCZrfWpZwOM
HUmJ1aPoKYuc+Uh3nBiW4aXoj9a1313AL2wMQ1Aypj67AAz0g3S0R2MJaJJEQ9jC
zLE2H+aUgfrM7JjORqtpuiUKdPEdSbFQLSW6i8X4jvpJkLr6mAY7otuzVR2HvcJa
ePdcKp3OjNmTVxmU4Uu9LrY634RseOtJCG/jrw73fhuHI+7Y5IoA3xIeX6K98ZM5
daRAagSA2bMWN1RZJp/0HBbfJ2poni8IX0dW08We0y3lxkhS7bPK5mPoU+qx/9bG
r5kGXoMbd+CcXGXKkH5d29y+u9TyQijy1ShdNGN981jWOWGGmOVzWsH7NQy42MQU
rq0h6hYpnhMleTuror8Ov+TIzB1pRpkNdy7XVi5vuInZwNCgeoDQ4EHLfWMQdWdU
qiF5IvBoKgHXCZ4Ru7oZ4hxNx5cIMcOfuAp2VtloKv09ZOguCJxKxbS1Tg9cXHfj
O0Jv16m/HIODsR/g9hwVK1Gc06uu7291vDkzt2vEDAlSRXNzCvH47y1YAEpuMSbT
QRmuCSfhqHPHkMnqfL6D88ILkEkt5+3YlCnVil1cY55eg0IH+j3jGg771uiiMnsv
ll7Tpp5Y8a5BDw0xg7ujL7xrKjx5ukMNowiZy5UhryYAtGk+1sBVzm4M2Mt/QqTc
dfctJxRJgj1a9x56yCeSGI+COsDMPtlPpbMEhOrSJq8CAahTWJBnfVX5gv4B1b63
d1JtuN5mOi2POp0q06BHE28fZyr9H2H6CDVwnfiO6A2PlrbZRvje+ZxC5Xks9bVr
DsDYm58mzC05rzCDVkcz3gB1nuBNhN+0JfKYVWB3l0oHAYLmDtbrqTFPt/Bm/eb+
xDOQV9uE8o+PJb3lUF3pgAmeiKZXv4hwXR4aKhtBx2K7kRKQ0Lo4pCs/rHTFg3cy
OI51/fBtEuvJQKfCMueJy8Rl7TcNeLKUa3IXnvzEHW6cu+fihAkMvDpn2gmeSmsZ
+fOpUAe6AXEScACMQaCfNBYEg/yjsnN217HrGzrWmM3ppsGjwoVi9CENESJUotR1
GznQAl3Z61os6g4XrRF9rq/XDAwpMYgAdh4C4ZuR7qa3zBolRyU9PeUWyNzlIylT
fircScEPgLFLDlxR2ewOsFLtAdPZvGpArIbszPKijCv+qO2BcBgaiL3hEPyhPpE1
xI1JvN7ob9E3pKuzsvyUs+2CH1HRT99OFlxE6Ex7NzjnUqDw3S4Yriwof9o9X1+m
CbrSfec5MwFJKaq0JAGKYZJvolneNJ1BHe9LANTnAdadigSAze1yIXqP0ucsqqQK
ZZPZgEOSUB6/xQpd7CDWBtWvAQO8L6heKSsfQ/xWcc80h0d8PRdHh5x4Q96V22Ih
Un2Mg80Tw+kaGKiFfKGVeF1nnghwovcZsG/2GKW5W2U54qSXHNvyZNGxu54TvbeG
PrdfizdoLreljS1CkebrM7nQGN6vDUAnpJI9YF0KYSOyPao51Z4OFM1ZnaEAPOo7
cm+8Kli+61yxA6hl7X29W8xqv+4N6MDMnsMmePANMgDOLSPuGHWGR2o/E7MgD1G7
Dik/3oSvKoUxVACbJ3flmsg7/68KJOXzdsX7+fOUE0XWgjVVfoDE0caFh5mFItz2
qcps4seQXEJ6KIMt5vg3oCfEq8E8CJTbqNEh3KUf45P+nt0ABw/P7UKbAHwCAQi9
ubKH4xT8gdyzxAVwOm+EfltlYRTGcuV0TuL9rkoZY50KzT2eksvVeRtsWwAbBLR0
SfQmQY4xSzBzqlRfYFQmnmYHut0X17pwPrY7yOPKToUs0tniauNiVMWoY02vvMJf
4TFXfIqXZbPXekhwprob9Bs7AxoBWwBVY6nW9EMiIZBmi5fSB6uHKPBwgSrxdPFn
ZM4fYIa5YJ1g3VMPM1adECAhJicQX6WMmJSgxXNxutQgD6Ka9rg12yqFTd1pNu+O
e28PF2LfDQkF4gKNozNOwHgrnywnvvSN7EsuxqEuXffSeHWFIN2ImySuAwVpb+PO
ASj6RddTDoDmWPjA1Lj1a9pNJGVn8hpuBOTcBvutcRKVsi31GOAp1KZ9siXG5FRQ
9pX+fELkoDrEsbl9fX/oRggscCVE3vBvmqS5h3qMc0NNM1YBXXNm1FagOIzYG96p
rNe9F+Cj07d9tN6omZGYiEHO/9AvLhg5IJCWEoYKF5amXUvlPzqxHzm3WV6qq+e9
DR9AP+p4EEm/O7qveCtvkzd0KnoA5/aPt6GsOLktlyfcTddJgXHEPUymwsJnMyBA
s1OjX+g+gPcLCrdRJMLSIHskrHibEu5YnIGoJkaa1Uv6NvmqjriNiLA6xKeFcSxG
YOFxwxBZj3faG4bqMtZfQbLb9n7zItF8sXUQIPf+NXdeVD1I+Zxao5Ca5N+93xyD
aspwp9NW++aLNM/vRkCA1kPILOkAwcxL/VMKd/l7xeeOTo2w695ICHMk2Eosx9M3
zAqFnf7tNJ6eU0PDIu+9pDur8JrReag9pcnlK1d3KEMST1Q1GjqcwLCNMRiENkOU
OywtIrjPJEbL1bKzp8N1scqoFu9YgphBmOxrpYD08nNOw60jvfDZaIZd4cS2vHHe
Uu1miGmAjU8cdNRAr6UqxyLcspM5ldhHcTXOeV1zotFUsgs3djc9L3DGVOpMS8kN
bYv/H4vkoqKL7Jplw0b/Cx8Rs/fuLkt73NRO+HK5KF7SRWxgMS6FT1cwW63DjwZo
o0ZGslFNWWSc3wBP/BHP4n0nrOzUVNF8PXq86keAUjP5yAYcidcftnv+/fOqhRFY
PuTlffU9ZSeN/Hh0SyeqSPOZIrzZfuGzVJyzeeZyJghV/7Wn50WHhYFF0DQIhdF6
FqXalBJDSIHctAyepVaJqSIFOKFSVazIEx1HUUHnmsHsogMXE0MG34yoUFoMAHWv
JBZR0Yn4TdxKQrny2aowy8qfZp4Fz46bH5tSsyoU+iw8Iau2VWLbboaIHnlLt9aH
gwCa8FpQylabKIIOOKWSXxKy0ZWw5qkU6B5eb6OphcQ3RIJwSHihGQj0RKUzzCF5
U9h9A7bk6dOAD39Yc5sYuAb5VTrPE+loIE6sMl6Ig3W8CjI/fffUS10YofZGnVHV
7tje4utDhEsS3gDegRa5U40ZBbvrWdUrKio5QuwKTTE6z6xkibfxXFvgLtwfdGcU
mjsnNKeRRlGHD1TNpiNkg1LaU3I1rIUlD3RdBvGtAZvoTjr26tapI8wQ+FJhnyCd
YEGgQoZ0pyfJar6zh3ewDDK5dlgI6Kq9KzvCwfQO4PyGDdZxD4ltbh4D7DeDc8/M
Xc0InByOnRTUbb//8dcnwBvg/sGsEwq559z/8Ywy3l4ECjO10IeuqZvwhhJuB70e
sZ8tWzQFpFpD0N85TudfxLIihhMYxhFK+4vhxv0gzhBXoSQV4rCdg7P/TUNirGoL
vKWlQxzeh1muUKpkMhsqzLp2wxUcprcKfCJeACeIUeLIkQIVtpvOhCA/yUjrGETW
DoZxCc4g9ugCjd0jcJL/SQOZ3QvrlrLboFw6k8CTpTX+V6hfaWsebjo2UKJYIpbH
rbPZMcYrAx3sRTcj0EIBHprsQcKXZVbdfP2Imm3gTATmVyJRZnTCJbP2FApT+O4I
sq5ULyCAMMW7yus36WdefdXVFMTy5KKhfjyZWlgickMy14JhdO/fbq7xE+rEmSzY
LcZLQwmHEYMYWZwQ7FVrEQEZfrdBg+frH0xztSRDlsU8JTPWvhI0mTNu7QtikSU3
X4yPA36RaGJQVEgPMhh/p0ozDdWkRWag/tEM2O52CXjOfWgKpAQDCn/wg24xiu0p
P9QX+oh+mqFVYp5/MD+S944at1ZkZC5CuNt1ncbjelkI4qrxEGp1RAMCVZFC4qX3
XmIvNouG1h/AxGwpw7fAJOVJCOnqfw0mAV1J7IDBPaPFNUZj0Kx6SlhWxxY5HIj2
MUDeDlyugQpQJg7lZI3g65AB9i+uoqFB1l3RqmWXXKuqZ4KmU97KO9RFWY7sJDm2
E56bOu/WqlGzwM9PBxpPttiyZkya3nlhPSpURZPjI2GWOjuR/IKPrg4rghtkr/iY
uovBG5ciVNhZjLs3bTeUbFDyL3hhp/hdOpAV2zKT9oNXsBDhTQ852H/PUcM36Kf9
X59ow34WXgLSbJlLYZbU5PqzU8Hppc6RnT6Ly7cu2VBPtWeVFmYXdBAiD46NFOuv
YXQ9gwBFydvKDJybQminVB7TroRYi73o6nWcqcwSpN1GORdHL+cbNB8F7KPU2a9X
wap6tXw8MTmy+SAtmV9JApGMkG/kj1WH9C6yIX+BlAJkCTDdiXa2Qv+oDbtk1OMY
tU1YOgdHqJ1ShaJW8rVSjXCOXpssupaeGYCcPkcDjngVwJUnQnEOfPjHN/TfZkHm
ydpSlrs/kJ7XpZ1Y2sKo1MCdnpZl+P0FDONMGPxdbWBHAo5SEvHdBaWSZeUJovaJ
ad0G50Xq42sJWZw0Gh6WQveEIjUAxHDNgKWF4M5Sc60qPqn9c+36n0fWpKeeOXKB
o2f/Ie12LiS+NXbwM1y9RjwTnSJcCh3yA33y0oUyhOWcW7Al1idKCyEgkFDehaTZ
v6mn5RsNdXzXyGC9I6aiiD0xZLOx6QxKlqUQObdORBfTx51r7c4Xidom9ZmitAHM
m+4Nz5+Um12QeJZGHP3oGNWkOFcV7yjd5+QTXR71nnbOcFB/dRhM8zI3a+q7zoc6
y1gD00eZor2nHd/v1GLWQpS66i1ZbLS9c6FEFEZ5lRxAXMUx4K4983rfz0a5WQoy
Wm2xguz+T+avKXg6rY1SBdlp9Kh0uQCP9+JKQ2wgkYxvAt9MwQ9h4xBqv7DYlVAa
Vr6t8rAHiFY7v2+urtEYvArX8dHNDv8RbrIUCFk2NUuS32z8XvvL7Rsr2pPo3HSD
lzexfjy3W2JLo/6JENELUoy66ZPXjpqNGwTGvHxyTB2ZMqTN5asIDDhIL/B9CNnS
ziLKxQt7OIHLTG/AqoXwjJdPNYGr1UJ93ddlhgOiWUbcwqcWu30V83GajRPH7UYS
y2StEUjygwz0/uF19/Wt+rVMUEp48UOaiE1U2xZhOGwJqwSyqBHPuXgxj1OP/+h0
K2WwYufhS2Tdbk8m/qUzbQlbCtkBcmxdu4Akd3ezAPYXutIpXrk5u54Em5Ho/N6T
0i/YrcwC4zTyaSg4lM3QnvXIRudCJgHhqE15aAQ85Wbv3cMmVR9XWBCIaE+sQ8HG
gR4sGRON1Qwo/gpdSZMZYySii4u2o2xArj0lG1bXLvHuJcyAYANOEP2u98IHHgDd
k7YmRk5UhxLp4SzF+77OVPphrXuhR2oXCCCLl76+IdFpOOQobtHGIYgeXRPbpQIn
/EWxN+1MDdEKrlgI5CRveMoqvXM+KdvohCdEtvPNlzPWnERXsuoVwY9Fpg3nGmYO
HKtg89Q4Ie9IRfznYekqKr3fyyz2U6e9cUG7gEpvpkZG+wNgFfrCXUAOYtqdhoAN
/4Il1gWotxQyQR4bxn2jUYMui3hIz7dTk1pYwfpJuLjAktYe3nCyy3dcDm4ZStkf
RsUgawpLypSwHhbSXraAM8fuj/woMp9gESxDPrFqDniw8pInMy+Kc+hf+j+U347Q
gRFqL+FpFgh398Uk2uCpkc+h1nE5vIQkPyiI/p8Juy14F+MNvoBSpo1xYm4sVBs8
1TJNk2zpin9crPyCyQKyZT1akDAVkggWMNjOhKb4CCWnIKAkC3gkcLNrfI/j5t8F
p8DaZC5OZeVawqCs+EcVITX0YW2wCh8W5J8cWEK0G0NvLXNwHu9Zaw7zPX2Uh/sd
vAiTy7XiPO/Ubpm7+Tjtlq61HmyPCA4X8QGbA72w/y0E6n+HFH6vIGktJeobxGNh
oo0EAM3+msqMjHXe77OoJCymeR/gHcpPTbyodOY1k76g7oKa/knuRsPgLm548ivC
7nXYzJAS+eiduWF/EZkm5JDglfqIV3tCd2b4GSu7/A5YEVOjA0aEwa++SKCmgQnE
GLZoVPJ+dYAUvoDPXvinLCNrV3cJK0QQUu5tMXvT6Jm9wqFNUUMcv4DzUQM9bLZR
KvDNuZTqmTg+9GQrWTKpx8zRxAbCKKCZ55O/0whw/VAEmmC01EAF3+Db3jBtkugQ
cgvAbOkNLruB03gDAAHHFJoLcoNFLbxvVFmckWpq+eK7aWZoPEnygwsYxxb6Qym0
f9hi1nklWHngHMFL0p1lSFkGX9lzWlUMDCU+yt4AFTu5KVM6cYBCRnAX9/jAEEme
ppYiGtxqvKEitm69caTLM71SDoonY9vyk6Ow2Rqy+xGJA0Aq3qEaySoUfZPAXUpz
XvkfR6V6KMGyhbKco4jMxlkgvn++puDurkWtPythAom4v71NbUpVpHoXUUN8PKOZ
6KsJlZVqtIFSmYGfE4efR7QfJGeJookrTHUbhXmfr/hAceXOsXh9wB5pEk1FDiCK
xKs8Xe25rdi253HSj8SrWR987KYsXSvRwnoMOC3hpTMYkP/F97Np8sDDMRUZdj8j
XsbCUOWxWWgLeJEePIs6h6gS3KViNKMCLLRiVbPU6atbFW3p+qiY79pzNtTZhmm/
02JfRBezd9WLZ4YooDmqnwskTNzwgI3c0mKDrrPXG+laM9SSCtisMCmqzaw0sWjI
SDfgb2WEFtU5mgsJr+CQYb3x4PcrrKbqgdHEs7O9niLdV0UuhJye1pwdPuBEL/nI
Kkq8H8KcUmRsjfKlz6BM11KUgcbNilBOzctkToNUlhjuNrwpy2P2B5zUk3zJ05R5
P1Yqpk7gUvqjNSqKPI20reWUAXK7OjwL4cOc24b7Au9bMbpNg/gm0gDHKEsJcsoT
En+v9buZPC35I9s5oX3E25+F2VnLv/bVU75gbUexGcz14tBPioT5kMzL5Tmdfxf9
kKN3kITsrpIC/hmYbZfFbQqqeNhvYzPn8e32GIx0iz1HwwlDjPhtoEpjVOofKpmN
wAlpN4f5aOgA9cpspQ2YWwk+hkWoq4IEdj4LvqEdKXc6IipeWr8oEF6Lfe5twMK2
xsCiHqWFqy+muwVuMwC92akjYIALwh5/ZSvhIePbVvU7jcYImf+wSmcWsZJR+wqX
pelqZLM5LgqJMzIebeyvX+aSOpDYCrdvzmjB3U6orAM+WbvGJEXgBroCUSR153Jq
kJLhL8uaC9LJqk2rRD5K3p6u7uos7jaNWQNSd1uTUAMr7kbz24JTrw9Q9CPNfHKi
2G0jq3naF856UimldSUTsRfCK/1sefE4UUPjZuskUz7oprBJtsJXm9t2fN1DXLeJ
n52/tNmoX9RNH2yAtdT8cwy8WADZ2kQVgGde5AYNO5bSW3oLn13K3ubbl2WfC21j
okXdCAF3I8A6zHayKVI+QvsmwDU7AMyFdnL5rcqoXzHYsoI6CGTzt8+U0NoxQYT+
BOebrB5eNOsLOCScz3n+ivGbEGNEbo9WigqJmkhWiecyrCshqw/EKIiSgVtyUjUw
R/n5Y4c+dPic8fZXnunBzoQZOir60IV7Y673XPjDtaFnMLq71i6bNwzolZXHDwjo
Bt+GXlGtpfRve1X490veBeqjfXlB6d6kzGKvdcPBhR9N53QFrLNRqfhs7Rmy3wCL
uenCQv8ZHoP0JS0JVcgzgoj+TFUomd2hj9CQqzKq+VhquG06EeI5WVgNL2dJvnDk
/EmmmEmA/hhusku2vzYtukgu/TndkNMyyegYfalCjcMzE/TEPwMNl1t4U+auYw0u
gp8HjwiEqMExTIfHYIA08Fy/txg+6IAgaqS/sv9Nde77UcBYJriDx8jUIzYxjmAB
0sjVssy5OZQYtum/i/K1MmqiT3pgTD3Lqfh8AibFlDEjKxD4nMtKz0Q+25vOeKcA
gRektpp/OoPufmZVMcSg5gym4f2G1DVGMoGKFolKNJF1iSclGH4Q+yWJj+ERW/9a
dCBNPn5oGC/qjGJbrylowAjTyR2CLSGtbUFTI7SFznUfrlgkHlCx5wAgKNw12eoZ
834eUBMmqEo/lxaJt6o/z/EN/FwPCB3agFgs33E70XOvuywLT2h6mOkkjzJV1IYv
DDTagfXUikn5+totQuW7ghcbOVbZUd7TAvtxPT3zlVgtF8KjzcnQ/oknZKnicGWA
wajRm1B4HE6SuT584eIfcRVlEZdIklGR8/oNOdivEwI4GMQst9fv7D08HltZltBg
oxjXQ5Twfdg3SA0glJN5rq23FXal7YDEWgm0vHz1+m3sUaz1tg56ig8hUQEPL3at
7aYAZSzdV41f7f4VI3rc+WMR+KgMutail5rCyJ4ggUNCB3VLntb9BKdgoiJyTOSf
QtiNsDrsqxP8OMVUW/Kd2m96IH2iGGmdK9s+oUueq7XVRZTXjXICcS6KNhvo2Ps0
kscNfoxyigOQWJ4FZ0iq6sDKRx3CynZOKum6AIHV8sLc/2BYJThLCZiGjIxIa1Cm
zVG00ycJM6zS0sOmUHDFJa8CP5hfloDqpTFZvu3Qm4heg/Q58u+00UD63Wzv/EIr
Y5kt+nt16YoYZCW/aDH7VpyFWS13S1m5XwnsyYoisAn8HZ6a58kvaVmY/CO5SfyQ
aaalS7AsXYQXnEovaMbXiEfynkub6oSTo7x3E+LQraZGhDTk/9e+hhJqt6g9Fwnm
QEOC4HFK4m2RbZYNxw0Hm6EXz5Bms7Y7cmLUvkv1OATlW3yKSaQD8BBAhCwEVb8B
FK54NrbELrS4eQqgKEoo1j13sg2y3P5L3q1zwVUNVki+9AX0JslGovXX19XaDxC6
MKtB92luWnC5qsgfAe1Fy0Z3cJLioqT2201I9FTNZNPwJ/nM1KjASx3OAGw7wWXf
XjDHv4YtrFxv7mz5F162nXxgTSTqVXogqNNH2BXMgzV9LuMu4LqLQ2rMizi9Pni4
cPrRWYouBfUvXsCoG9q2ko3I5QCqT7+ElKLW0S63vIa6rW54JPCW5/OWH0Bu6xlW
ybR0WIa7iszxzalxCIf2FDK/6VWOxMdRXFl+vwq9L1AqMME6vCDe80FPQCtswOSc
VZdycGiafmpUBoNrzoLX1Fd3TCO4sekVJyVEmwaC/2lhCGAvtC4721TXumR0qOd1
ZiX/uQCssnzcEtdL0gqMCVc9bcgRfNFhzBewW6rOaIPkA8Lj0wOfUqToOpn/QCkt
tP0gWDRwsLZMkfOVG3/FyHW4B1DQeXfQbHyfByrdOjaZYCw6UtRqEyN/qd+ImriD
GXak3EuTvq4COZ0EeAg6v3S+1+d1I1RV7osq6MqkRdQ+dM0iud+YdE/a3W1CCMcK
AraH50v3lemCUnieXRgNglrVL9yUIqRIUNVsl1loriomGMaKH/CiXUgF2e7w3GfY
qIsnHDwUAT8a6weGebbW6ZBkhxcRZkRPNSubbDPaJrA78DTkDhhnrVGuOsOrpwtm
QG1DK8LRjRwzMg4eyyAgxPG+h814G2T5Gg5xU4aqWbjekHtomMvm0gwksbTxb49M
LVXGBespYNznhvJWncqX4eO92YZqCU+9vDN9jEXKe1KizfDSvKv4eOT3ywoyL6iB
8n7iN1kBS8te+TQtRZtWUbdtzBrvDk+k1smGIiSkx3PKV5jjixXrsPxAHlzKXvHF
r5ASPCe1mO1x3OJj7qVmyvR8ejKX4e9iucrFlYTTNw0FjN6fsHqgOkDy6aZNYynF
sAGPJI5KwNFdu27nTKMU8U2Nqt2IG+yvHXeAidTQF9BBPGQtfC03gVKOgTJOmQO3
yhsKL9rrBchW2FNloO+B8DzWhK9ksnK85I2Ebjuzqp6ircxvrQN/5s3ORFH7vp/s
sTdmxc4FBnN+lqVzkvAB0ByjBwvPkiHw3d/whjVg7cLaw0nEr6QZDOoytxmjAs2X
Z7F+k2GamJbyN6KnQTDGI3bT1aB7TpXX0AssQ0M8e2bGaZXP4Bj8ui38jP2G1/p9
Hyq6s42F+yeBEsy7iIhH5EiekTPUIVJAGDu7scDYCMcJ8tbqtNzExuBa2LloUoK1
1g7wUCKE0AkhH5G+P/qAuUuioKfhnCh38OwzMgVr2E6w2H3+0vWq8kVb6E+UDykA
4+82NGTcwhYZekeTIL6cclWZbnOTLss7WJi/gZuB0yX0zUGaKdOuVbO1CGHVSV8O
H+QZMy2XQYlWtqIkPqcGlVz7m/B2TCPVOE3sTaYKQBv162YW6YsP5lL7LahjndiE
AC+bdZTSWcWfmOznYXG/MN1jSuXBdckhK40rrBo+QRuuHLUD2+JQD9pqTavFzdBL
9PIKJ7fHNIGLJymEMAhR9bI8g73xz1jfCv3CHW8sLdyB8BndO1g9R6VP0BaeBPUo
OZuQWaY/rhKHYxYfQLGBicSswRSSQ4ADRXvFibbtH0lvvdfXAHZdkSWzwv3yS/ul
bl7K6Xb9h2NJBs2RpYzPOrTKrvOK2dA1wgNYfWzThWbOF2MBxh9B52WHNZt5Z5rF
4a5OTdMNQGL1xgiRX25dMCuUf7Z0LOMuI6BuWQfxbdau2tdQV03UjFJPULTuiTi/
5TyVWGu7kWidj7H+J7tSz8qRISAYbFoyYBjX5y1sYL4xChEkUgOtUm1D8ljOgfgh
droOmArvFG3FmW3I7NCDx0dq0gzcjR/mk2F6c6EJGe2VJoEpIbIEgkZgjd2tbUcW
o6fxaEdXXz+7h/FbOXnZSKYXy1lFn5cuWXidRNCIgqOuTXnwi7DkPiO6cWvXVOuB
UEaL3jDx+fQzGjucM50NSdw24PqpMyYgXMkzXnH2Pj+Qwrbz7HRK2kbG3SYJWSxk
F+I7jwT299uIPWtuC6HTPKjcM8+Hdg59SnZBvdbqB9gdlRuBONjN5Gfd5iqaW2Z+
4UvkILfA7JgZKmei/aQ+uCvq5okPXYAJhuiuBI/gDja4BQgjhrnIYE4/k1gWl6cI
5W3QuGZXlsMZg8eL+kAn5f4nn+hnf/w75TFuC0fSCjdC/ddGVADY5lXn9gMgVB3c
kpQqYrVe/hcQFZAWKK41zajMlxlUr0Plhpdz72DbU7pU5Kx7JG3zQp95H5zCSsY9
K0RvLO0msYrRQJKNAqrK6+I/7rvKO2/VRnaNbxk/uuuv0aXZW1vGhKFlubhvE+Vp
6Jk/I2mDnHe9sZPr8Twk6zXKXQlBWvU0qRj7E+S/Xs9IvxPKWfatU/Dqmeg/9Hr+
mGByMC2MmeRAI179wCiS6Py0fZC73NhU8XOfjMXZvV2YEpID3mzlDfjMChaTr0uz
2ifvLmhRipG+i6AVAaOLp9czdQ41r1pW3+oOej3w6NK22XY2GwV51yDg1lczOKUp
XkpShjNpw3T7AvnQqT9+Jriai6vsUYkG92eMzP2UQ4B6Vg39oPMwucKzyht76DUT
/J2qZaC5gqdQCuvDS85Ygj1zC7vQUouUnxBN9zgRTft0TQRyg19T/mOPMF1Oei3U
VWutSVsSI2n+mrKLu4HKOGWT6K0z4eDalX3BtDmOy3mu0prSuhu+LJRFrBsaoXCq
0Gh3uSljckuEA9cG8ANktjtpasleJgwSCYXRNur6w3Ax7EjiJiABzDOMVT10iI3R
rlxc3B6Ik8XC6jQFJ/mPhfB31/D7pFOFcIH47au6Yrf4NUB1/ThxzeTByjaashWn
VzgukDt0oTS/pWyUa4DAiNg9EcKl+jbEk5np4UsYjAzf3ON5K5xkS3PyAiQW7hL2
Z69u9q+K1MDrFNWl4w/cuF9etYRwQSe+3qaypKxnJsRhRrHPAuOW0j2Y8jrspOpP
LG0m6sBCysLagCmMA63hp57iJHPbLrrIxd1t/ud2HxMNsAVza8oMaNg1ofBaiq7E
DDlnVHSfdNyANUtHZ3uBY6Ddg2Dv+4u9CajuyeYDCd0l25rZp6Ib1b3fPNyXMlzc
jPqR5E71DEwe8U4ydwrPFilJ33DDk5Ks1waNTwsJr3p4T2erDP9DtuDOFKDyc45Y
ZfM8fLgLtKeOjgyBB6UwM/Pf2LJyCMNXkrtv40d2SOtnsSKvEyuwUQbfDeWkqNgt
xPSAA+xEJwX1wco7YotEBTwh5r7YgJHW0jBLzB7+pAfADjkNU/VLUliQVDkNkcFK
Ih4tqtgVdbpesvjR9NnFZaspL+1koPzsP4uYqlkW4F2chiC4KV3ToBhb1Kh96kK3
CKGr6lRVc9gUF/8iUVSGuPKN0W7Js+GHVjqFZvnHMN2FtI+P/6HV1GRsp3Lsv/Ch
RdgwvH8S+/iQn3hyXjYndyfvm/v716WEyWpX097oSj/bSDAmsO1cOpGgiDJ5mv7f
H6mrycPDJ5kHRw9V5BG3Epyw/vV8vLHbyzNrrPdZWALe4kV/ipHhQ1WzY7fE+IYn
Az0Za+4XeqkORuMem0nohDAbQbJWGrEmgZGu6LEmcHtd+oGQBvG/646yxTJ0BA2/
yANAFMzfBzfE6MTpuzOgMN0pAU6t/kVVATgmGJB4IGq8r/hJq3EeKvgCD4JXLlHt
/4O60WlZQ778p6rJz/z3gszbIEDjCkn5FIFDFmEsqNVb8ktJGjskfi+TUe8DmvDa
hYhvYuQGC4PyteQ7FEicxQjKwM96uKOdwe6KbDlEkfDp7fkarifkmgqci73Ne8hg
FPsN1jsDhWiaftvTXwBd2Y8H1q2sulBz8YZTg7F+ya3vaKJEA9PrlYba+FPat21m
4xUZ0MpPJLJc+UWLqSuQ5/cDu4YFFXccP3B+9THAF5XO4GSevl3lR9Z+w9r1QThx
RcnwAuwloe8U9oQ93Kjiv6+o1HyM2jvlKybFs0fhhK2pU2Vg/copkxmVSrxmETZi
xxDDfzO9bmUik/QhZsc/FR6pOXoQxFikkg0P5TiK5HMUdnK1X0IkQN0VlX3fRgkI
z+AVt/Fl9oSVDtUgmh0a3a9Xr+75cJpqg4CLojGkq5e8MjLd9S5mdBoc/rpDFeCs
jBPV+rjAderPYTiA32CbTc97l0HiwQixhdH4b1/96svkF8PL5o5tYY0dHYxFEscN
+m8mNMtN/BFgOWVjuAVRZVOeu1aoN15de3LsUx+EqdFwoKTSWUkWpTSBmI6Yzjnr
j2RtOvqROBMnt++xiEZVZt6G/evadUe2AtB2p/b3l6LSfP2baRiUWgOwc/VBrfTv
Xak/XRN22R1SKbG6CHrUHUdMW5fvqeQr3VA+/9mhOrdIQzCARHDkynNvctqmD+nB
7qZ3r6pfUacEwmGZRVJAxZj1D7Wi9JVZ6Zd1hHjVMcTrCuzrdUIsx2BOjIcN91Jp
PcV5WHDrmn46e1ungx9GkFNbmWYHminDDBAtZ3GjGWgMrjGPJgWuFAF7Bk+7cg+v
r7CW6hX7DYBZxzy9kP5/TUKV/w+meElvDwwC6uhsrv2cBpZOlQEcvbo6Udi9GyFO
2U/kxhdrIn4VHdRyLj20Hs235XDjTnJT4iARRX7dU1RycLuMsaAvoW1abiTumyNm
6Cn5Oaq6reX6x2ZzYWbKS9Z0ljw0bU9i7e1gwiXRJxgHRfA6qSrW/W/vsXe6QkGH
dJpQyK4e6y0ChPaM7kulvBzM4nupUUkeTUe8H2aanXGNBh5xbusJqFm/z17xcCnk
1JGmbkiCOwGlFC2mIMIquWy26uLhN7x7WUvI1zkHDKM26bdnbuLcf0Qfp4Wy6Tj5
4tLN0bqI/Z6hn+KCsoqlEy0+Ke8yvSy0UitGpUodF0//wKLBCo1yR1vDZmpkfaQF
6xnA3IIX0ZumY62rmdiqcZ6FbhzhXKHxZWaf/FEkLrnXe7oa/g/pvI6Dy1u12xqY
z2UfLDYTUX41+t89/IIoQQiUNoijrRZTTnxx0I8/Q8MbaZEjFxldrs3b5aiTO59L
rFhCx5Vqa3ZRJvcP91ZxYiHkgMAWn401fbwpeoMGUEwsM6RaztTw/HcJjl/Mzs3b
p6pJ7J9oDVe9kTVAFCzZxtK7vWyko28HPSol3jz5PS3VhYopCa2Ieo6/FfhF/9nS
qtOfbU4ZWU1C5vLJTk6AAVk7RvFLhgxcTLDyYevOZVF4mhT5hhC9WuyMR6zGJnd2
yHXnLJg6h4zGFshu8YuqQ/b2nMGY+F26V9KIyyiUjrYLuuObpGTjqTztbjo70Dxu
GRLkRyFEjicxtmtlLCcs1L20LicuWIOx1GWJvSp88AkswAiGbefr8ooT19+oq3Sh
nQKBSRSUM6vVr25YKCmu9TPV2eq+o7/djRJ1dC27e5dUIJHrwCoQsqSVgTmbrQ+L
lZgrFvj+wd4uRbpIYgbRz/ZGBe7Wr3sobdAW8/x42UwaE8gPHO1yihn5rmBds15w
Nr3KQy3GuEx87xQ87PyRZp09Oru44yLEJyWJzYyMmQTCzBvpaVdI3amF3wLHdQMB
X2eLO08f/fh2wZNlx8QYPzvo06v5CEyJm/9l84Ol+dJ9pPXONECrtrx+gCyMemtD
HLDkKpIat6FMn6YHMHHCKNeOt3Gg2NdAfWqZng1/7OZujUPXs4o6KmT5LI1YOCHD
/gM2BAyDe0jJEXC0A7OxnZ9zsHlRNsPu/BoXbQVnnDtceNVLk5zQUgE9RUX7kLXr
iF8CxYsOoa96p9ZEKUETp2JkIQTsT19MrH+QdVKRLTUnlHg9ElrgQ+2j2EJm87/m
DanhEUDgrUcJtfC07Kb+6dH88C+po1I0Ztqiaq7e53niHlq78EdtOIUL59BalQaE
CDvuXiVRn011A1wBWsWGk/rxdlPyoBM7VO4XLYeIRL5dDeoSMpt40QEoghfTkxMD
v/FGq4bYVZ90C7Smm8z2UIgwRlDL0OfolUnRH8fOk9ZPdJQN9oDt5V5LMruBS2cw
5cUAh/w7OWPdPrG59THscjegetW9SOpvGVwZTmMgaQ+ftw+g2qYyaoOVaXBqwaAg
tvi90x9xXO4DaYlL83EW4ujQUnWOeX10BtO3y2P9zfCT7U9hnR1dT+2n1QK0Ja2c
xXsFjpWRmWm+62UhjgbfxtUVeS/mm1XOrr9egRzsGsw9mTp4j0qHoY6Ypl3NENeA
jLd1c9TGcOeGr3x3ud63VMIfvi3pVvkoNbDDEKCI7zWrh5qgaY7sUI5CL/g4Yz2d
FE+R9SlOEKRUXaIRVC8FSvGF6unsQM2IbNh77ctDP0F/DOiIaeZrKSOV40s9ft6M
oKxNiDY+PwXyKSMG+L8kMpnlYBYCe4UHLnGQM1hqgcZ4O8TDS3UWyN2MVEm/ee2n
DOWiNDeaJFQX0stYvvJdXJeawCA5Eg2NWTbFc24oRmDHqGkTPAeQr5VciLv4h1Kq
mpSQOjV24fPg1FDIKirggNKi/UJWtKJl/S6dI0tvNA8eEqKvcmOUTRg+POrDDxCe
v5N6spPMT53bCZmS0BD3myMHvxmoE8SJIgFNOPfGR96McubkjUDtGLm+jh71dJk6
4HtficaNy8Mn3fT/3ifuJI/eyUG4omp460x0+oxQveOD1/rTpWpwzLIGwIuWadeG
uJJdA6qsfGz5L1Dax2y5A401KtOCCcB06TJcNIaOZWrF1zbQrGcqY8zmiwKz4nhm
PTGo/u6/cec6P/eYV5yjsx3jV63Vfv6l393L9jAENjuPLi+5o+L4Udy/X2ygrKxo
a+l/ekhkoKO+65tSefN2rqq9OOIf+s72DhVVgjX2bl3FKbPIf4d/OnztnHBcN6pS
nKrCu5Y9sXWx//2MRormDeaVh/3pOx83dZeEdpO9T3xm+t3jW2ShpZ7BFCBair0c
uxyAp00Ou3/AgLKYAYPuSqOMAulGf8tB6SaaDWF8mhz3RHWj0aNNcbcN6RCPWEsP
4Rk4jj87qjBrXTtcKr0osAVjLvCivYhIzz3xTrVBAEXtU/r3WzD/taBtXbLoRthO
BknKk6TEwJny4XOLQbRdY3FL/RLQd1/Ac+g7h6I81Vtfj4Qc+NUGhWr7Zif24+G4
F/5m8/FXW197quhX3P6hPqPct0Dm4bxCrd74kV0gPjS4UXEzt+Fj1rcUwoRYtDY7
saW6gesY/yGk6epSkxJT3uRKT84JiRV4D76yjAk6/g0x8XuibKV/ZBhAkGifP5zz
dwMRBLp5kub/uOmHDaxMTWbKuZisKeZLX/ZWU9i/R0sACd8CIgQ5dlZXDQsDUyKZ
Vru8wpk8KqmCZF3Q4ZMbQmdxvR+BW1HnzNDjeOrIMaMyWFVoeTTgEMWM103UlRBg
yb5/+6G9c7ayA58SoAiHCqBipFMS1sDD6S+8x2XiBGeoMccRp2dtRO9vJB7EwGA/
bOcxr/ueMtKQP2VTgdQnzPsSsAIhY3K67VYvKswGQnuyPhOskC4q0y1SQsjCjrGz
ouNW3rDQMt+lWHeQH2j9uD0RnDS2eZU9pxy/+DW9uq+TlULnYxMBdLMXKaOBtFRD
Um3C5HxsbTG5bGf9aFXFh8UyGxRRE5vLguXt1BVuPzj9IcCaNoPIstH4f72Exgoa
gYCi35/1Z3SyqHX+Bk+FenNIoYGA+u8ogH7NtihbUNqdYtHAlWj5JOHdY35SfpW5
zSjKbwstVeT9lWSuq/LYb307VvCSjz4tXJFWoiKYDg5zfkYjFqDW0QgV7J5BpCGQ
KOyWDvPAp7bXwDhKObquXK82+QciiE2VqsMkU4mRqVvqeJ2rhz4Z6wO5iOVA43qz
Biiqf/H/lckfk/E5c6fd/jN4s8SwCvdyXjUOmEMWRcbJNOSA3dhiTFGt0yWKiSDD
WDvT5IVmW/lUXBrG0GNHv2Grt2p2mFq7IenGjz5s4KQ/yS7eunLXoBxbocdYmSl8
Xz0QimibXRKlnjgkcoWF2bWqX/3B2jk2jk5KcJpiVjdP4/AW2HwdDpNwrsgS7Fi5
7mqar1vgmAaezPQG6gKkwCDjFH6lSIobOq9p5p1Bi9TE8ofoV5yEce3Ck2JWTX4W
N0EoEFVZIUuAHrkRsHJGXt3dD+Yzv8z/l6k6J2oWH0CF8bQ+tHAo5pNXKnKnq3Lf
jFdy76GbRB51CxoA8fWgV+aJftRwVnjtLT5tTIj1Q/sZ27VbQABLK1LUA0Xoqx+5
OZvdYBDLkHC5Vt/DX5Gv4novaX7618v3n/kArbWuj/dDd7WQ0oXS2hcKyNuD5N+/
+SRFdRd3twXzG7kLWy1G6sZ6pZNKUVNXwpn2u6SXYUSKgVzjKu0Db+RjU/mjIcG1
smhx2Z4AtETLpVW+X7zgK9sXAEFuQNahFbVZlGDlPGV22R3KuA4Zt72oFBfOfvt3
43jCRrmvnWE/SL0g1s4ksRWfBMAVNDw3pbxX44+hhRAS4P24fCr0FgCvBX7EyD3K
iTCc/alyvKX1+TKqffaYqBZSGBVPIfOf+sMou0GmOsn1G2K9OWlmmXJUa56sej/0
acq4sVBxb+1WWQCtBmMtmQ552vfE4xJp5mPdpP9IE3vrf7EMNqJZBxisBXdtwkB2
VZa/Jh/Wx81Ez8HDMJQ1zwiItWiKyOqGZsfRM9xzwMEkZA4y12Ryx3HEC1iNRqUp
v+N1MWvrXlP2SIfZEqZ2PPBFrVTGhj9KTLzkEb6AwB+B9j7r7vuPwofl/rDU4Gr2
JDrrWRZ1iBpywGDkd17h8ravKYxjxsD4xoxsr7pbLLJRbNFHCpZLxHkV07Y6UKe+
0MBoGfYKU07KgchlybptDMLgy7DQWlLkOP6cIHF7Pyv1zpu5tnYTZscmfj+L1QDR
hIMcH1KzOCjXlWLNvLZ2teU2RkrZ5nKqHDgptY7Lax0W8Rz1GoqN0lCl9sLnFvDF
C1jXOMzRWYLs2aa+GTmcXdxtWUIFAxfkHSBwZ4ppgSDdCXLLDs/8trt6fDpnrMCF
PBXm16sc1oCwZtrDhpROmGnW5vldAthIEEy82GBQ8JweJnGnA6//new0P5Viu8yK
7ySprdGrGjD8+WFVAaISt2oWShlT6cT7gFZ8iZODfWezU/YD2qFM7OTStyBJTKmR
srpTAU0CNr2Oa9rRJWMoTCGIe3+JHzh1gYFJLi80eh4GuvcYZ1URPZqpDa68QQYC
1gC/pYg3o7v+kYI9TKp4iKBkGAMZuHPOMJELTwIgSrB0gJ07Wd6TlVVhLBlzsah7
/NHJISwTp4UTysGwTGbdaOaQncJJfrR7qSRCplxvfdnTz7CJdfjzGcH9N2qhNENT
dfuOH4Tf+QkmiCdLOkamghFlE4Wt1uspK+j7OW8SjFB+cyx2/BPvXbX54efGiBvU
Rz0V+m1e+dC/sPvtDmfgK3Nf+y4pE6IlZiR61N1ArQqP9uPKdN3xHxRKfdIwvjEE
XTAu9Z5k5w5pJF7eysvGU6L9FYwJ1fU9zCUC+QwANstVRNMff/Apjkyu3rXfjGcD
A6PCtKPMYpHrRUbinrMycdWGPSKibFhyM/EOLKhVXpbGb0SpH4zN7gvySZkcElwX
v/K7h1QUl0VtaQwFfjmXYIZsDLTSW2UGXjrQ4JhU7/Kb6SSOeMJnUI3XPgY8Mb3i
nct4B3oYYqA5DeDe1KHQrCQ5hZjYBuzX0PI+h2669GBGKfplqua2mR2DC1tx5K3S
9yITwYl9oYrRlhdj5qmrN4eL+Al8SHFpIgAI//pabHEGE9B//i9Ska8peslq+epe
dPlzbYblfVMuDssXGGjvK08B1/qpSFlyTme+M1V/zMSZbksy7zj/B4U5cjSohP3f
gM7gFbKT/DS0iJazZOffNBM9+iJNfr/VtOwkkvAVSRXc6zonJIan+2nC/655z0KJ
XhNpAQV/TVZnfsLYnSKThFS9VjT9zDdS71haxVwcdlIRCOvNEGVAsF5pxdLjNxpw
mI43dVv3VmvHNXK9Ju8tIiW2Pehdkd58spz9YHPJ4NaXDPfDprsG4/jGp1QfINFX
c+k3Ob7r7PFjN6K1gAtFoc/i1O8A78TQlCLJGecMSA+hDHgQl+m7+goz40vDwSX/
hja/MiSO/OP/YQe/m03c+QYYtrOyd0eLaILsdDt8ApQyuC6tiv134E0msipc5Yob
TjTfWNzcrDCxOg5M6l3KkKUbXfvzRdw1l0u8enmAttbqk2JwT4hp6VAnBaZ3lGrg
g07o/AoZAdocPNLV01LH3RcMw7BE6lEXGIEBV2RzzLpE8kgvKELff3vl+Z+h3CjI
8hQsBr6SL4g69AvHfnQeZh8Q1fXEAbV2nuGWwmJJfQYsd3TIL7wKKJk3416fvPAE
nWiJCqVb0w8VNCmJL/WmwGbjYfyhlUSVZE9N9bm9fNFjgePL7XL2zSEMp+1ewU1+
zSv0jmAuuOVvEtOgiHKo5SYVfoab4RrTDXwdrzGTVFNGvT8N1MeWevvrirgXNX2S
n9MU0efPT6funNjGVCkirFKP7cYtTPiHKyrsjxUvOKyYrH5vqdxQ0Tcp6QXvMFI/
eTx3KtqUqAm9HwwnPCevdDhfGsXDjgYJKeHfwWaLLQ1NvkBzTYzi+1oBDKm7221x
7807dnajY8luo887tuagvyRQSXWvpBntHY5t5ORPtZNWeXj2RqGwT5xQ+9WAtLx0
sUDXJJv0hZIWX4rgqhjXNR+BbVSMWthP4+JJ5NxHtefbHTSXNXdcvyyxmvYpOdb/
oy3W1FMTVrsK9DpbJGgdXzRze/K7XEBif3e7RydvJekrdSf4ySu3IWWVlW5iS5Af
4RgEuhdv4Dvk6/haPiYaapivW5BT5BoFQtgdgGZwrhwBAt9pim4xiyFSQvkI1iWk
48G4uP9J1FF4q2a0ZvsCr/w62M46mo2N0QdVGbWrHY3xx4s5AxVOgdWDWSKIYjgk
QMhy19D9RQcE1tmb92Nrn2KcK2xamNSDawwsacRAcpfy3ZfqNdnELgIVj31vdqog
6CT+neMIrp+250tH8DGlQQa1RgfjOI7bgPDF3LjPMVLXDYRjpsqkcMZy0Ck9MZxF
oKXi0rSdspK0a9G28O+KJKairIHTjDEvHEC6MxcR+3P4dym/jE56/wLsaIBfN7cH
EiwbLUIlYWglA6oStxYyIWSvui9+uCyCZkW4p8lzqy/gtf7iH1Gq/Z4wxU53yZXw
ewK0A6RMbBX3tsC+2r08X7/6+zQT8QxFyyz9PoOiA39OUwb5PtHVLwwpP5cBjxeL
9XOGtkACk7bQhhtwmZb+C3wPvijkTOlPekNGsCbmj+xBfCssNbDAYLPYCFk9iE0P
3DQG7vNIGZl0GToJpeS4bq5t0fIk2x559UME3IoOTFLT9yArT2mCGvqAVvvK+5vS
KWlmQZhRlaRguWVN6d/xFMQGL2LH16kzX2UOFsF6m8dlj88XaaCsP6/ZPwgD2uHc
jNj/XzPx3wu1DHkpTOScc3VeYCPu1cmsBxmfp2oq7jLIeqjYP7nd1k67fm6eMm7y
RfX/PEFwvQgkwBrfvcBTLFgSrz6ocnTHcppgCQHYh/wmI/u31zA/qNkJ0NyI2fvI
LumnwJAHtiFG/sRbeAhN5B0b4SMSi8Jxz+VqbDeCQSRdeWovgN7PueExljhYv2gZ
Lrb+55Rh/bF7Z03f4wUdEY78NOOIrP5QgUxFza8ytT7rV1doae4txxGdhX8AZotm
9PIjyWAubr/lqYckJA7buk0xlQzkwpK7P7umvU9RlWJAnmCRU1ESfxWy6TFA+UsJ
cz+iAHwEqDmuACstoJe/gqxObjXAc78wfxw7/dXvduSjI6DnIWSuhxhBfI98McQX
Nn8IhiR5KMARkPF/ypSmSue5YpbyZ6pxIa28uq2F9XmCVbxmLugQ8/drTCa9hIH+
Y1V8DWlrUpJ9wF/Lar8RbhR8rl1vXGSerkm3b1IQVjErFJIaIDvDsipuwHHwr6Vs
hHsPcj6XVes5vM9XMTYWL5evIikcO5KjhD6XJ834ID3kGIzZmI3YlhaA43OOktoZ
4lqIwnzN7iRk6d1yPzh/WHbXsqhDhu7wueo1hEGA/FMTr4eix9QYVBQA8GuDurqW
hU/OXgkUEV63L3tJW1UZjaRa6wy98R/AvIa5eah7JZ/3YuABd8QUatL1AZ/3iMH7
Pur+/9F5ThPgJQl9SmK7Io8GpxvVgU3RfpgCIX6VjG7IeB6o+7NOznw7lRxU5bhn
kHHSn06ghMf6ZvjYWUz+yghUUApW1mlacOhfOkCGaMOulOmiBhFsB7+iPY/zoqLT
++vb8lPb1EQBNF+AJoxSsDvx4M4ch8ej8jPI/xDcQaZaZp49UgEKfboYI52d/AY3
m4RPwDgpyc9HuhNtmIhb0Uni835CoJfxalNM1JLcW956EWpYlzGDdtgjxicx3x96
HxD7C6CfTyGuxt6Cpvu3lyA4KVyXZkOfSwLBK53eqSI97BMvdvl0I4Q92wHtf3/Z
6Wl5fGIIwa/UZ9g2jrD4a5CcCqqN+Ae1dZEMomV1tA6z33dahGYsVlbibq4fb6mZ
DDME9jiZtu9nQAPHO5aenejG2QOdRtdTGyWHsW9gaxt5TU7bh8szBV4CkHTryQ6c
deNx0RfiZWU46uRU9YXlcRl0QII4bShpzjPeCfX0cvTGUw4vIITbE6x7q9tx0Pc1
9WUC4eTrW+weh9RI4gpYqfJ0A6neXPZ8DAVMfrO0SN9tUDaxl+wUY5nvbjZwR98T
uG+nYt/1P3nEZOZZEU1DYL4q4RsMWp8+aVHIZ8dfBeuKU4k7Aa8AC9BpxmgjneWg
qTvzOcR2UY/uJskP1TlSv29IZU0WDK2jAJOTWweBkiiPjrIsurHJRWyiEMZ0X8rN
G3EVraIAAcbIISb3tEivGGOShjSm8ag/H4b0FBQXC5/n6CtkjeUy3FUUIxz2VrJp
h+ZivZtypz6gC1GwBs4KIoa/q4/EI6Q6CyMAG6tdvjS0VwDQ+hO6a7IRhkbmVjW6
nltg9ggkpZvPnWdSsSVDrca5/Y5f8bmeCWyiPsun4wf3wTJLw/EUwiu09Hw5ve+1
lIVL54QQIovynlmC5YBWbcCj5P5aYQXK0xk5cVP9VYF2Yup/L+PgiEnfggS0/aMH
CGqF6C+pYd79XE7Idt5/wbBDwIgA/CrLFD8/KAELFH2G9rFbPwJzzMCXXZqRmbxj
bbPiWng6ake9rdJjOBDY8DaSL9Ub8aOpIcmIBPgEj3AUCzTlsS0gNou/CePkNfmF
E7Y+WU0uXlQoilxsrz3Y/xYDQcgJE/uguQJ+XhWRv+bOoC6qVzK+CpxkTCuVVPfi
ZBFTpQLZCQYQ4hwY0Aybr7IkwqqJFp6Z/Ok9Tgnzh0pug04lUpdQx3D8+ZtrKyQO
myoGwkgGA6cGWm5O7PlRbpbww0D/32ylh156R6ny+3qj2C7Ur+P8Q9DBeNa04/Z+
6Ek0QfaVSdP5rGxByPc2t4P9ILw/4UElwHqLhs8O8jPL/T3f2JaWUz37D0j7HaUA
B4TLpNkpSvKhrQ7SuvIfjZ/ttz6WqWsPS2O0bnX6yn6u5bOmJDSs7UMBL/bkSfs/
wocqtphA3h+zckOcircnPrC3sBlwmhiZLgL7mgmnS214ZqXLQQOH/tvrdkA8a6sk
ojX6Cy37N0E1KrhFtoszEC/rrawo4AQMRH49fkU3yl9qv6WcK/BKWBv8ZbTBnweE
e2lIW/CbtnKjJEtPl+NlwSVTKxe/ZEl5QwYIwc2F5nGSmgMOyfqr5w2pjVJQWZra
EJkmy9Q7gH4GJYDGsL8SMG+i8jK36BXsX9IaU5HqIBVdQsXBeH+n3jL4hiO9FLGz
TVohSTMoXFjo70mJe+OCoypzNAVJg/8WwMIUInraVH88dVVmGhKa1t6D83UmYc7j
BWZSO9+d2I0rzHRmNCoUIQoATiK2cEWxAHnZydivOXdfPggTgF9l3c8I4rkbiAl3
XWmb7qK7W8y+dmKxUPH4vpH+89wBLAAhZTzjDg+6yuLw6bMAXuEZUbd4M4M7ZqfY
phCVvzxchriNX9jSEBS4jBYDQKlRwLU9FOgDAc01EpMaSTaNl4k0Jb2hvmxq9ySR
a8T/tJBtd/v+pCK8f7CFKiXCWL15oi/1fTG6DU3RdWMKEE7VTw3EyMujZAMOhKro
qx6Pn5xfexNDXctsvHg7sZfLoCBEK0zObB7MOTmVZb6dWcl84aFVWhZf553YNWGa
TzOF/mbIoSmIYKoQBzaICLDlZIkCsOvGQWWpzQ4UG8AUqWLlx9lez8soDbtPuRYw
ggSLr0qUnBCK/ucJSn9QtNWPUH7ZOfeOFxjzz3+Go6K5L//at4dTGIheOu0Kbi3j
anixIP/nhCbBnjEBm9Z+TmbZXKet7ulJFJ/yDWw3+CdKIw70Rv1B3A+BtYniy9u+
/CPjD2zMzVz/Q80gri83WFTJ49nxnchW7IXNZ9ZbStaQ2yxtregTdSUsMN/Zn6Uf
DjeSLg8VTGiZOMcE1Ob74WiBsmQrg6ozRh8xQuzQ06XKe3HNTuWc56QEKpixKPzC
uM5oW7xjUxg4wHVO3JIf4FfgSJBcR2oX1XQRTiYhgcHiFfXg7o0ebvHwDJa8GS8W
0pqk/iLk94gRbSTgp4MEh9CF75x13HSprn0sVYxRuS9ZXugcml210BOb/lyufucY
l1Z5pQPWQCuDY3OjyMyg9v4MvuYrUHNt7/h2KElC1OKnHjz7U2/xe//DuAnC6YXv
LXB58Ylg5DXUv/Sl1biOMBjcsUPfVZKQQFuUPzJPfXHnabvLu5r63fTGKhvKJyfY
jIZycR2Ujb5Gf7LUwqgiA3LQc7BDB5Zoj27fFhaxr4CudHKrsYLXCubmsIvwi4sL
o3nsYV+Tzx+/GOopm+0I+fw+jcO7ddmzIaQlwXO+WCK5Ea0gP2qOQe4aaxzAsqIH
fZrQemi+3RYzzj7LbiuEEP2azvzWcPDOLXk+3Xg6u24ce+ibOKVkyUyEJH3yLbDo
7EcfL46K2EMARo+ZsuTOZ+56VK5suQidvMUDBiFGGwOuw78hXMj2FkZIQ2ccHhJm
8ShOvtVslLS4RXviE+X4B3F4oTPK2calVUo1bBuCeZRCTOzUmfYEJKZbdikE2tfo
rGXmk54mLz9TG5bXxjOcphFngekTMQURG0z+9zrGgSDBeVn8SPW+I75WL55mOrGU
7EdMDA3DKbG5KCqBqPFApOsBlPKWWSOrwmrLiU+9xhsmIsImPwmFGki9B0GSGpQm
ZtxIAHIcUX7jkVoD0OwLHsaW5pfAug7T78GKUFB3eikL3u8wo9aTa3nFDpmiXruD
90jz0P86rZtNUt7GzMMquEpnYHxfAJhccCMUIsBzu71RTfuHxGAsM2Htx/UKL/pN
BAWK0PIhFw8mglR1GwLHvIqHo6JJ1FqYIm4QDAbViLDnR2nbKvSGahjJxirWFwBM
1LmllUHahX5Gxfe4j62b8TYFTGqydI5lP4SUvaRccVotRUwtsYj1AKPO4Z7cDlYN
tniP15+EWrbVYVTDL0JvTa/Eo9QdNBi8j78o8hMFdpRvkAnvxO4r+5SC2Dbm4Myq
dJCHsv86ejoS9NhzuR19fZBU+7hM0NGj03cyonkumBU5AqzwsIKmmEAxsN3Todee
Uw9Euujcd+aBEsgStbcnk1LNyTna5rdGYI4qodJVK6oaGLzs15lL9wBUZTZwXi/z
5ZFbp0AMH9h+tfkFtVz+vyuLpiJnIvIBbtmicD3hURq7VbIpU5bP7TXMA61wWYgu
b+/uWL8zAtZe4KMOx+iRqIiIl2hUVUFw25UKa4eiy9SNQjtw1IkUX2S4qpmrrs/K
Zh4atdWnfmwmf/H5ZEMdWN16pcMRYLw6U0ORhnD9M9ff7UOZfvzHKS5sBLLN769M
vo9x2rromZh22CbWCUdYpVLVHjh2dQGcUIfY3Tl+kTukFf0CFZoTfxpHQd8pF+4I
0+BLJn0sKho9Q96cn134caV0kdvKw6IUSB5smgMEVaY5wTu0QjXzG1omwK24kvMb
Crb/gM4sWh8sfnO4Ca3ube6J96EMT1FIEvAyhf9r25fBeTM6AEy1Vxa3ewcNto4v
A9edT+dSzOoAowsJJYbdtMgCYmHLyGuwT0IhajI5GH/R4r+/EO951TVUmDzFKijI
JfmvqExfTIBXJZgEVZPCZ0FKodJ3VOcE/DU7ZKWOFiHRxcckusEvSOeEOezfzD9u
WT82uACWq2fhgBzZidFDQpUr7F5bDaCnv1lFZMvpyJi9/iYT4sEL0o0L2tE7l0x9
IVqkrJ4eRQfAR1iVNpDFKA7g2ZXCQpLyScDutx1jYub753LTBOua98zNcG7INRqa
g6DFmQdjVdOO6pM5SBq6Qb0ZIuE9qmZlF+nzEMFDWXgOHCL22O8qqTTaHf8T2Z1z
QiYfLBrsxO57+D2gz2guGz7dfZfOLb5Z39AhnTz70fGl9c05WfBFM+fnJaZs5mrh
IsKFaLLH0ABtblescEgkfXmPorHOUlh5smeeJ5r6EU3lgoiyH9TtJEwKb2tSr1Ge
7Z5tqsjiD8E/jum7wpW2mvf7gdp+Oaghh87ApRd6NvC988WM3nU+fPK6df7UTMws
8NSpbCMXZOQczXKM2VZhQQ5nLj9A62Jxt+2bCwxL+6Uwka7zlGSv2vr4fPRkeRsr
/jL/cyzv33uWyo0zUojsub5y9IbttZBNruZpojO9U72jct0pja/sQq9HIb5DnJnf
X8N0k73WrnLOEpvqNRM0s2G3s+aOw+sglqeegjD21AArPRdUovue5l8KIE/7Moxu
a5naCyIZe8SF9aBBX9jeQaxrNvqup71qGoH/xBjIQK5juOkgyIxM3h29648W2zi4
47tMXeRdLkWvyDZYJ1hqjwBFv1G8xR7grPC2lpo7iFKI4oMz7aXjNhuPiW3OuFOh
KzknnzRmyWlc+c9MfyQ+LC+F8evjOZ1JTPwi7PS5pwODVpG9BXXg8vCG4xlH2SvI
1WeoudNw7I5r8sU3SQk2oSn7KY/ckJ9sgramOihCe/itGV2PKbXCXVoXJvfNqYpt
VOk0YOHR7/uWftYdNFz95xr3LsyfxRkgqdnh8ZV6jK5ys+Gufu/LfPsBj9CuKPwU
boN1G/yU+YfojBu13qPXelomoVt56d82bkgtuEf0dtcLtF7jZiAuH6CZ2jGNJW62
KDriIASVlnFTaPxXxivMukz47YzweJ5/R8uG6dkua6zX/YBBfpfRK0fkVv9Oeqii
evOmNFDYLHELSCgR+S4teR/fwvlhskDHmaNcdS0qDWCOhqkFyAGBKExBkVPSyiHf
Fq3S9ohtCwm3Xep8DcTkSErq3CRHdQm+MI1bkRWLEGNXiuyiF7c9N57QgDckbIFD
5Jwzpzpq2YUOz6o4uBNHk0+WkEc217P/vhADffNUKA+8KkDd4vn3Y5WFL3awjbma
sq/VgXBqHqhoo15jjpZ5m3vDzsRY1csx+naPJgczhSble2KfQ1YnN5rZwFiEMcZh
2Ex15Z5wrK/pjNnIdE37luHIraoFmIGNGMjYZ88jbyb4pJWkCEZY3uIwoELexp5Q
AXoxolGGhv2QlGi/HzYk/oCIPGnVmNdsqNrXF0V9h4lum13xmhaF5j1dypZJbUMS
m4TgJQ5BEolnDvJKNiyTRQQsw4ucrViVq61RLmuhYBFVxIf5bqL1Xw2dSejzjQaK
/zbvJW3XPNCNaOs1O2PIHkO+XkeG6xf8L+bXvHwV43UeKjXQTp8pHw+iUPunZqq+
DrRVCWAgvinojJf9EDaWv9m4uet/Booxitpxpz9Wccaq4HYSX2cqZ2+ux1yIMzqe
t8E1bv6p/82YBTVQk6kdURuAG7/FRRwBWib1dmWqNIkEfkepypiPfbAEzImFK8Ac
YnPkFLpjjnjqxdVgksmB+uCMY8wGNYtzb5CUPDtThq9v1AMGcrmZtnbDO779O88s
1lnt3qy+U3pVuG1Qq/yQEkDZ7u1YweQcnUv3vgmGaRQJMllEebPQv1cUg6wbEqXf
DMvKtnp1T3asKSWrDUDBLzPdks+rBIkInyI6R62vB9yY8CEJTtkfuk8z+9MgokTz
4tlzVmQz99lZAeekwAPdXi82CSzAKCl0fY2zKRbcgRMkd+MpILUkf+7JnuD/wpDw
tpnrzVpRcUM8mZKLAVtPwnFURz/Y6k7NDI3Yxhk8A2x0VvOLrEfQgOosC0UgiZQP
xTty5fPK8DXqv5D8Zbob8qZtIottW8+UOzI3O5iviwZuHzLM+SK7Y9ZLR3J2xBTY
gzjUvz56/Zb/xWKR2RTvZJV7x60qKMlMJ65l+6qndYdMdZ0FlunKC1g5LhrEtgiC
WB+AibmJueDh3lEXGn/QiRIMPJjbCsENkkmmpNKucmxEINUx/5Vm+YpGhEWG4stp
DGJHAOTcl/Psq/qKE7b0f55ZhN3QdRVpmq6fnQGQ79Gp7GkSPsYUpMpzwoszH/Op
lwqPzc0HtpvSNvKErkJCsAwqz7KSrcMCewtOTr7Q/jOZqT4+p/Nrzd+1lGen/Dvc
plJ0ZghyqDqylOgrs72IVkSbH/irobLyZ0yd2xjXVrLjuCJW2q3usFZAmnY305sI
w2NMzdzulj6yhrPCf5VXfc63Rpjlk62hxZ3kn2CuM7uNwQ+EziunJBcqRhkPU2Eg
4UqVJBZyHoW/sdE6nh5Z12IlcYN/dFJTN4EV+/rqMbdFtOPY2kgpc1z9YcjIuQ19
mEQJwH1ycq3vKP/tOMZnqSN1IP1sLwGQxF6FDdKIef1h/bOyVzVd3mlmOjLY9ZWT
RVO13XO8lr2/vaC5GDTXM7EvAxYMyrq1kSUxg0+qpraFz5PANz7o17KSkjVtU3ai
RPsdGsyX05sJ87Mz0ha8rsheCM9/ha38QJK9Sfox1OEmRpq+iDyVT9q4FxpFDRW+
F5zisc/uogre8gF5xyHAgYuJMRoqYDriZZYuuEWFQVLkRdazoFJsgK4OIhjrkccY
0xCxKyM+Uxr2P2uMxcvFKWKtBHzN7dWsXUZOAra2CpfY1zShzvdyBj/5KvBBHvHx
8IfPPrm3lAH53EsbJD1UTobdlgfi3iUW0C2SKkHG23/5EdQV8+v/o6mTsRw5ylOO
lUoCUJV/05d1l+YSLaxSuB+a9ZGakAlN8V528eXjERn4MrTsRyJlJd0Lsj0zpZV0
WA9HrpDaK1q4Aw36AQRqSuQmI/be62DqPK8cl4/mfv8KrRRbnKP67pZPpLNU5Yyo
XsAx4Z0GCOe8W2YL3MGdI5zRFlV1Iy4n/fgO3M593trWTqkLd3ef7E7vGmHUTdxX
K/l/YyvVxqEleSlg5OPvnKhzHwE+a5VDJibE6wgaojidpHn63LhBTbouxq+6EVYu
on5SY0CZCMi2l5ZP3IDjVo+F2p3y+BYXrQId3ep3dSm/QYgmY5OPPOtiHMKaj9KJ
cVSnXkFyTvvedndhfiYLtzDa4SQ8jb6/IjKlh5fOhF3kWMG3AbI4JfzlEtYvpQHP
Z8nHAtAZ/lQPCnXPe6M1Lm0JnZvojRJU7M4koc0txxsIqqGHu17MLpnNnwLRq/X3
FEBCFa9y8ze/NDLOF7H0tYQKf7NFj7V7nrpDaKi5+1Ca9v6R7CqQcqag7pwI0v6b
ZYn6cPvr7Qs/2DlJ+fAogdKaRxovh9A7yXZydubDr+L2+8Mo9DnA7hP6xBvs76sn
eHnvNc6w1gEYB8c0hLfdYtr0PHbgVNKAPm5CZ/TLAEKdnJ0jtsiNcdmpShca+4ML
d5QVAmNsDS8rjX2NuTQRlneNfquEaSSat8iRU/tymZaYBwKNEc2OHy7rvxeQf8zF
uyvoplKG+GnSHnPE1WLN1UkdFMyEwWR46vxDyTYAEFLtpJzSNCbl+wTdaRxcr86e
lBgUmvFWWf60eONyR4faceei4Ixu8p/e5L7SYOEULJV4a5DliRHJcFFRCJzLfplT
Ao/IJurNJ31v+FzBWbA6+1NBuGJJHRbIPt//QctNMPSGx1OAG3kU7jeYNsEvkmYY
7lliiW6N3n0AcOovEf0KWqJaq2bxJEO5ILJVZPP8xaY8pqxJ9HekkOIsTbw55pgo
3lGLPqbG/ljJUccaAM1OM0iIWa0YsESmGUFj1DdJyVHjM1dHt58uNpli6vK6EQT+
AmgxGNHgwLfXkLW+zZIyutEJ0lBMquqqKu/+mXby2I+eI0dqT1vVHYQ1iMEDmiS+
ytxWqT5fEWkH5VMo6277WrmO0YtaB4stcJqunpCm3JatYkURdk975pWHI3QYD0Jo
nMv0dBcNAJgpc7s9rhunyth0saxiRTEp9q85aBuEkvacOucusLP9Cywafq+6+ebq
s2qe51wFxAVusdRgp4/I+WEsPEADTo0grihy9JsNj9GX4XISH1XmKssclpwVTJol
MEaGiHMsig+u5FEWCtKTv/jqUF8wWqSYxUTkswh6DkPsV31TU3GFs8p6hmP+pSQg
GPmoGjS3DJIwfLS9ki0/NFn/6JtzttDjNXlXVa+8H/QjekXIlvCN1Sx2o7vtOhLe
uZl7pQED0V9DryqFfoKEcmmgWpCwLXSOzdSz2CO9Yu+/jiXbV+ir6wvGrKzslr4z
1o469DgVYKViF4PZQ034LpAMCsZnoGvTS2FcPqYhbsImkVf2kPb+/WsDSpSGOl/f
YQHT382CiJelBJPBJnP/JLKRJFMQpwB5QwdHCd3dJYEEwhmi0YpbK8TR+hAmlUxk
/rHoQA2xm2qdiNMeR462SP6fucnG8sekGFsTp/cPXQbx4LCc6K+tJqDWR+8foalg
1ZN4IKs5dNzu3DZDeeCYdhexD0BCl3PV5LjFYFLOS19rq0XwQ+wRSTPCT98coT2i
Ooos/JuI6jpHxj9NE9wHHu6FDuClMdOP5FeMJy9pb11C4pes/8XMy1TSvckOsip6
A1lfsKegysCGUG/UZ6RBp1Rzg6sDRhE409jlvhbke131B9u4B9ut7Y3N/qptKjON
gGzY0qzWhGkaKmp4P7PoBvcRVInKPyIT+P47M3TIRhbJHANlUwkCNSFO+Ckmwm+V
6hB8y+8OjLy3bmodVOxoCLhhHlHPX1a/aihxlZtFIInjJ/BxMds8c9DCFFfJiJSC
gfG2vJME1z5kUi1J84MWutPaMy3oEp/wbQ36yad2hQXcJqm/YjfRsjq3p4/HDCB+
pI38We2rSXp62mMlUXYyNT+IeC6t3XibfPfNn8/GLLrhjV7MoKQKyumnSZalckL7
QB0I+L4KUiMijk58JEvKvRQROSE8gpoaJLg4Pi21rm5I90kocmZVak+pfHGGrT/j
pm1e75ZPpjEPG1VV92Jo2KU91iRSgLoMS5hDWX49Qr4aAgZn+2Z+qWrRrSNW+AJs
3QLqG/cXV/03tuyBXdBD5hiPpEUZXk4MM4U8dIdpYquUM7LgLLwqvT4Vgov/TwJl
FsrTD+YkUjqLOb0qbruxzlAGT6ervxDmHLeEisKXQ38yiWioSlq+YTNndrOXEmpo
ZdZnauaKYRjD4arOcKh580XYUS7ba4dOAi6NeEbrd4IjSmK/2sNHXGewMEW+2s4S
l+yy4bQ5Rx9wewoxnjQVUV30dgchh37D7jATBeoPQpAi+E2CH3GEpr9J4f04S9gE
hi51Rzyg2y0+hQeDeIcB3nD2JtOetKgo8Qxe+7/9ne8G2iP+fe4L6WsrVSkrQWuQ
Af4pPQ/7Vfiw2h+0mRl3vQ9KgS9jR9sadoPxT4a+Vcn6pv8/gritKRCAutmtbp42
vtYO0MDf/+FMo+PLp2Qpmrfg6MWAc0B0f/n0mgb59FINXHt/NLQaheuYd8Kbpn6J
tp3lktrnCdbt5X/BRnf/V2Js4Bg+Tu75eMyv29CR0GB4oSeXx+EI8t+8fFBxNUyB
d+4ZyT7z97cHGfBqlvLWqd/pPg0zduuJatsxMAaNnUp7fG/Y4d2d3wpg91CHrxc/
FTdFcu5+oUnRwX0l6qU1/HAageq1fQyf89VS72yHj8KXF0Hc3ox+p20/w0VOweag
kvLc17AQ5vbg4D3oPXtAJVRNcBQEtDDHOJmH0IFF+o8k+IMyqM1ExSZGMbea0ytY
RTh+K9kORHQiR3SGGnFjLrvFs8mnGUB7uvLGil8EavHiXcIU+NxiyqDJDDWleYL0
oM5y7bEbJ4vwiS0qLC8BnMZR20DeUM78YTbJebh4t1X2m4W+kHKpNECjOtjbVcH7
ttDcrEblnF17OeWvaBfwgn1GxdDG7V5wpeB9CE+QhLZRh5+Cs8+FJ9VnK2+USZ+n
iGYmAWrvuAXcPIdsFMfzEuvac2JdFSamzxE/xAgn3XQuyVKpoFWohIAiryPSrn55
Vv4D6Cg2VrxRXPJv3OnwkaJUcMW417lF4WDWWBd8yEWJZkXnf9IyhMEkf2ttFzmI
2oZhoRz7cJNVOyE+lC6W+s0AB81t8skqf35nVoZ4FNsz6v9D8PgNdjEvnnRa8Qhd
/44iPQOap7odnxWDqRNGdQbhsfm6+Skb9IMu7fqr/w/TkKA1veTRbUSRdKr1wUUY
cDXKN9hebhwY6F69bLvUKGyMYUNSRBIJkQvxwxe1VdDtW9dTpnjgt/treKftvtfz
yBUYiPlOavKDxL53zCLi/TI9+gE7oTalH+AXrDfWiGRjQOUAPSzQ6EGjbkyeiRWy
6I0n4SsqOZquHnOxGDEfHZA1byLW2LhLVl41aJZjrlccfcVRlvUZkW2qtwswVL59
pbEhvtbTYN8KtH0N+ropR/J9F/iTr2mVcIK5jcKQA1SDLWzHv4nPclSFRpm7uofc
7iCAKTJE0ULb2WqIP0hKjgSckiOw3sken8cPx87TVEnrSlPbmv9U227WBNT6hnEn
TxQF0M69jk8KnBinjm7hkYCP4Ce2lBkzOQ4dhfz2D3RamKuwiGZOz0gAjJZ227CL
Pc+TU4B5U52uqox5DNpXXX+gnMW0aeg3jQCSKaiyl8x2ZXqHvNbXUjMtCKunHfto
DahbO9/L6EFKvw7wzubLr+zt0ZSODxPXAuLkjZ0qvVpHPU9Lqaq37AAJUHfPhj5t
6pEoWrWYSRcMfkGKTZZraLiAPF3ZgSp4k8Cjv8gcYFiScoP/2Q7ayDipHHpidRzE
9rSXTCaGzgpGcyxZi0pESjNxtCMCVvGG9SXuVx99AW03DRV+C6xskBiNhYbppDQc
cW2KYx7TawihcBrWU3iwIx7cA3aevarAW3UO49BP3cf4Z2uVSkoPh4XeVe/k224U
i1GGWiSwdxYITD331o6F3JOr9ukatHTPOnsKQ3bWRNMRG8R5xV6yLs2/qeFlNcXd
DL33wytwY6je6XJfV6WmB/TYGd1NwB7oi4BhelT0bjvpauisJ9ksp1siVrzsSCi3
jzc4DddPGAVSNKxkD79qKOVqlnaPjAnRjzFq58KgZLUnVAR4DMOLr28O93pKJoiN
z/U9ohxYR7gMqrYPm0dEoqoNvDfmasDxKOXovtINhSghsc6CsJdyCZVKSS/rgT2Z
8xwZld/3xBafaQ+4CCaPorXnH7+eMJ5c8ug2noNJp6gEjLBjR9L0orI5QlnFc42M
sqk5qyMnE4oYmAiDvM9gRnGj1WLvwr4kQmlWbrZ5WsCTuqDDeFO61zZu9zK8Ae1A
kLVxHQFKAQzW47IsS3sWuo3HnzxJJ+t9RUSMsMHv5wYnuTSogIYC+j7dxXCGItpr
kHswoNhOtTpf0AbT8ayOk3dHi64/U5EPfm9kha86GDr6Y4xmQuJdwKmerXOxDTRd
wY9iKi6y6tXdHPyrLNDsDFF9nf+pwHQM7OsuxYQ+hUYisZxHnO+9hdpeLKN/LITe
7+piqIVwJntC2LuTl7HRH3SdcISYf2iPJNGMD9MntQmlFx3GoXpwP58wPwaRHVJ9
JVJdu7ng/iDXjnzLfLV3sKgrW9kdp3frwNp5hFd1SU2k98TCBsjOc7/ePHdmy0cF
+dMxR858PIi7A/ULb73Y9XgbySK2mGg6WLGr79eNYoJ6VpWMbtAJKzZ+3f6tVwEc
8IVqDJf/MYCVvNnD5lGGhmMttAY+A+pHq/pqLTYFB453YDUQwGwUF4ItxELJUSbS
BqxDW/mziHGRuyVx0eFYzorloLuchH04NbBbd6K3Zeimhpn+x+nMXAUnAEmd0Kh6
F0NqolFG6fvnee8sAJc8bzSGL4dzdpRmtx5AhLp+/6U1X/5EFf/sFsk3dZ32c3pe
Uvk0PXA7lY5KBNMmihsVYF0pBaooTsE8uo2n4/E+/umed1Ty5/F+p5yQ8r2ps13p
Hpz6y2s/79TRzGmAgBzpq5KdzdeKB6QWm5lfUDNOlZZET9KQLAhuoKLpOyAsWf6G
ShJoBoNT8o2tZOlrCCrH5UfEYvbQgLSsPbEzjirrTBQXw06yFrD+XO8ghAoumwMZ
tyLClvRAuFuIKUPXSGNXTXisUtlg0MYGhrK79Ke6z1qhx6x8qJFiL8C5Lhg5BaJl
c4vY8CXm9y6F67WSLUlWcl1rxc2jEImC2wF8WjcqHdngN6mGdFc9dJBuCsuVElt7
E/j+kDR+j7d+25zZBEV8UP6r1Frl1huOZMwGhvsYMvI1kn/CldjMh6u1V3YbLxtJ
VlCp8sM3JlVKJqHu6MeH2NSsg9AV5ilFX5o5f5V2ymp8vWjFh/cmbCNCqrxqScRj
SfLe9bA9U5ojR19JqM3BvKaqqH5dwhBAGRrHY+CS1QXAzBJks8Q3lBBDyVSziwX9
Hvi4VSMoY4QVqMIGiw6Aqn2sPBwZ7LNw7rzTNrPdkgbVjkjI4rvWcYWIv1VFQyZy
kSlo/Ao2SER7it93CbY6r2MiTmN7Mj12sIUR/sN8MWTA7aQ7dmr1ukk+YPdTNCeb
2K6vh3vmqWpC2+Pu0etQ0IlECxQtUmy0bi2aYNCNrBylXVYhnrWbfxcd6BxvqHEQ
p+ppqk2/RpQogMYaMHOxUcIHg6PLiwRt2an8uJc19wLsZETjp1BLty6H6Eh5fz33
N0Rx46E0ZDA1kv+GuCg5Sj6dQKfx7/oHxEYML9xM1jwadBNYEeB1+OQjGPoniCfz
Hn2CvC65dEd2Y7Mr/StYET/Nw+E1t8J5Zo9meRLhvtGv/lFSsZdCwtc6FRAn1zWS
qytAWiutQ4xI4QoRIiDyyN0iJYmWjCFGW8VqDyAWS5Hc7ubz822pEY4Z97Oti8ZG
aSieI5HIKWWYqkcqUHJYoANQ7KhJWuMMipGOKEIKd/QxqYAwfjI2OYP7iVE20fsH
8UycKQZIQjrUBZ+K7ompvNxCTeXb8ptMPSpIhULakJ6Eb0dfX4B2Gz/n1rSn9H3O
SuwaHAMNkgq9bVlYff6DeO+UWICQki+Ke0CzwEiaaXXgdJHq3TIKDcDJVorbUNYR
/FE9ALnMuY8aeQur9ya8EJanAJdu0QA/bBGeU06JFBPEyGQ1nd0ZKPnKGzsSo2Nj
4cGNv03HGMx5gwXKsMx5GnAt8nzEERnufoiJFCaAYKexFFDeUpPHvHGsdH0GSaRc
a5puurYRHhVQLov799WMkmq/ifCGAFBlbDBWU7IoZkL71a1I0Kz4zwcIp3sFeY8X
4Q/HwSJSmjvZMN0j0MEc3jDVLRYdzoUlwqjsaVxB2KAbYDVivitHE5HA9Oe+kC3D
TFy90Zb0EBWTZn3/CsnRl5UMzdeMrDdxYy3k4JcXq0XXcc8p7xcECQjdecGF4akQ
id3J/ApKEomgHipCgKBW1vlAmMEhepCSeccTz4RkxGt8OCeWvYrGoAdC449cuo8m
iEKETEycZMaVbbAN/VAj+p8mvWkegYTXp6nk7Z7oGTh/Slf9TwiDoGdJDeoXS8gI
c7rhY7jAhwH/aI/5RqvtfITJrFB/Qc7+y/1on0qxzuv2vm2AptLkwjV5s8gOymFy
fhx2SBYta8wvj9SLUVN1t4Z4J+ZDVFnCt4isgzAYfr/w9qT0u6BY6vyUJ7gK5Own
ewX8R2qVYbosV51LG1X2AxrC5ieND84KDBkIpJIueMqjvL3qIbNAdkUZBuoJvpky
nLaH1VjxzStyVnqh4DghLzXuQubZFRMVqpKi1UmRp1Bpz7OHrIY7CHQegkT5F0fY
J5adxlLfyiMfipo5y5c1X5HyY0QwoEfmf563H2GHdODhZoCkW3BUTh6x7p88qrca
rc73SvSjfEX1PKjuG26bglpeyEDaMiBXAzpU55a9cMkKyfbF2MzR1u2j3OmmVuLJ
nxS+GEXdYAe9O7LoMnSrHWDirpvUbGyVlDSXnnE7DqIeHOURe2yg++VnCtLBfg3s
gcuKHVw5Pt8CDMVx8N3ydGxbitL9c8H/flxEhVy1Xce6TCm6QRJ4I18B4LT5qa+q
BucNa0MUiSzFfCbSY2NZZIAKxEXU+nhouYdybcYKsRU9PYsNbMQPVQjtUfAvfemA
YU/EXi8mbOYn6Ku/QL61miDxzvOpoiam0FlOs18QByWIgiX5ip9sr/6tAOZo7s5c
uaABh/SM2NFkTXNBG4ukNj8l4xV3fuw0p4O8ZRZ4o7ZOuo/aNsyJPKzHqjkJ5Tmd
udJKc+euvTDDSdDkvYdqDQ/16pNXpDPidVnoT95XrZrAPC1U+8lKnv05SJla8cbr
SMroXE321XrdM0kkNLSvY5Ie8MGzI6TOsXyPzbv3kDF+5LUaxcuou8iBiENgLWYm
anFvK6yLqgyTy4+zZdmIu3+ZhBcrtEDKskez92+zmgw5u9SYM2Pg2gLUvThIluwF
eGgi0a982ts40ljwAbAs4NrPK1iHaSeWXWKmTXbABhxSM2POzqSQdg8pWD2rg5kx
jfoDT4qnyguyftCiQ8pWJGU6x4MK5bp5bbZ4jGtU9NOWDfQFWZW1Sy873rc6yDDn
dB/IsTIA75AQ+4rKmLN4bqgim8C41FzaroQSbCDun9ZMp29vbxkj8qZUel8E7GJo
QHb1JHxOoRLFwW5on2KXp2JlkU6OjS3MDT24EqbxhmRSQ+CiA08vcYMnrARWZlqG
H+/kYKdKE/Ysux8G6D0hE+Bpamt92F1Ep97XZGBjJPnXnN4yameqPdLzVbzEL2dt
p4/1snz+xhXcASilbbummTeP21OaFwtFwiY4UnJxgD3LzDiLQD7wnxg00GczwbXO
Mb7E8VlpknIaSOtj0aGxmavc3PcHzn5HvmdMfK0s0IBH7rdJQ1BckS4s0YaQLXhj
5k7P9g1059gT7KeNEl1RbQkRqlufbDqRVtaRRF4ABnyKCSuiwcvouJJgk1ellq1Y
7rG2FBnL/22NmoAjNg5lGDzZN/4y0N7QEFkmTjlF30rmhAMpTQZjhJO5clBdsiyC
ikALTTHi+5bT0IZjZJLyr6pe4aCce1E4bnklIdAlpZHdsA+jGlSCn8bakGiUdRZB
XH4mzHlXEtUJh7rT5n35isKlJoyJNLxkPrLEeNsxDu5tguYcTBMqf88ImjunId6Q
rvymGRwLuFamNg5gD5ZLXI4JTEXHKpBNkNbyhpwd3T3/g1l/uXpnDi0TQx67AH92
izuigN3kEK971mERkfwypqGXDfKmHTZnTAZ8ERvVo+z8aSwkp1zjET0MyMILUSmC
oc/rEZ4s86iXBh9U7Fv3Q9SvucFb2n1BkJL4R9RQzgD4ChZkE4cDk6lfAc4kV2tB
hZRpF84hNWHN1gGQ40PTJLd8XYrdzKeHSJ7febs0t4o8dS5PbHvp1lp2A5v/l6kP
cqNZKYf8eq5tlhLbB5H5SAsPO4ouD47ogXJt3a12Rd6Wel3+S7Kwnhlgwq9Ua5Gs
OrnO56fQNQDTW1IB/uoklA3t8G+Oyt4qq31ejYEy+tvA3olDwRnIEp81JQDoOV9h
Xon/0hrk3wehEi3LH9M8zKRGVF+15YYrPfCDPc/TwQ5bLhCaZz1YFPiz2ENHohge
eo3XnquisZ6VnVjp3Z10ifFFbTiIwYJ6cBbwI04oagBO2UPKHFAeKigZK9eDROVJ
I6fXYVxPJXK/iXvG5L+yv/Z5OHs+8cbjlDXltqZ/ihAE6HihNQ3u5LmPitJwUeTw
Cot3ZxwqVSL9Q6JeVNZkh4zGXOXjl2+GRIoBK/68knF3w52u2AWTN9Yx3fpCKuEF
BerRoLC68t+fAtyqOW9JWsrN076ilpzQhE0s7MXO3+4JcIi+lJw/Uxe6iBvWp8fy
/dz88fz64pRADvTUGyrPbgg/W4J6FLmB46mknMUnZ2UTUAhHejQPrwXQa7BE6Lvl
Dq2149my/TPwpHEIHNakdwqf1Qiib3bKPw7/6+0MiLfhX25e5HKRTJz+NwykjDSv
0dO0NMWni8o6r/U9d4kBOgLOHjIygnRfGj8tHRBCVV9Byzn/FNsGLt6ArTY11Lvj
aFPuynVWBUvcAlg5orUxXJwoP8d/7BAEkJnS4Zc0jLvi+YPzm1SLfe2D7eLdpZQy
4y4TJofSa9Jk5hXE23h8c8+H00Pw8vLR4HdIgDF23E2XKS4VFeYUzafFnrbgmOE9
pi6iO0XtaDtxA8N/8MbLd3LvciMTTkPcJThqy9u9EwS8hZhnC2zDckGgCJikn6B/
Bs2Vc7xSc4J8NPZdbA5Ou71lhV7veco112yYi5oRPGIiZpk3E4AponJtLONRLjZE
SFjypjUS93mI01FnVGwrhrWAxMR6VHSzh2P4p4ITDavTASiTEPH2MdNAx4ry/UfZ
DBKE0pKYpPDTC0gX9KvuidkjMDz5vvlfNxW5G94ruECNPcHdBQut+cejLVjilDPn
EKBqx+/tngQrtDz3G2KB7/NtQC01kRGY+AaHQhMTNZBcfWDwVvFgrosC1QfKvkYZ
sS/0Rt9nbEJAeW8oT72r7s+TQBgtQePdv+kH3N/4iq0P5fbb62xiXpBN/zMS+dJt
dxqO4+ECjB95QsEYlPEvZnCv7LhN1Oia+/sxYZ8dTA4kHywF20togd+k8dRZjmqU
3RJrcoJXtHOOUnej+10F/eSMn9RXAiY+olA7VICLNrg2Miw3JZ7E2+rp1sauLb7Q
TgitOW+NGdXRLjewAVexKiPGmSQdZpEVdb78xFW6/3Im2OcNUdOKjnwNToVUko+u
tMocusXO+yw1fvDw14kV8CD+jPzvPEFtTGYQarVvs38AaSV2U0VGiEeI2EGdcxJl
KPMae6mkB0JJuZBxuGUiqywfgUUQMIhEhfHRckdKnfEasHGB5UOe+kwjsng1H8hN
pMedkPKyXSKak4ZvVmKK4vlFLZ2dv9PKR6C9UgNuWOBW9AUaetXayS6CkUaUBkC4
lSqXlvI7mt5tX6EW3YZUu1m2PM/WI6xglHlOuOX5j1RcXtgw16D4/9/gB3Zn23cF
rAptrvbsHIRzt6pW0Y9EUxEf0dCQSA7rFvzJ/AFnBgmIFi/39hL0sS2iC3KI5aFe
ponG56G+JaBQWi34nIEm10F3lJfSXhmqu0kcXCrPe+IQhFfJpOG/XtTkFNcF7ygX
064Hosy5Z/8aUDYEDi+ur8Opfv8Afvg1KaH7lfkNYmtmYJ1UUbEDdOT2oMaFhTbv
jmC5eQjfTUn8DAGQc9rYS+SbiYdVctj7uCq21XP+w0hWjDAGpN5ZmxvzHkCjSSVU
GV34G1vABcrWKYVOHIGzebLTFT+npiqm+z04bYuiCG1NnhEbdP/kx+1BSyTDqghl
BAWjju8SQKro4Kvrj7YYNOr0wj6ZNpybsQfEO/8/SxbbAS0xI2pxJqv6MqVKx3Ez
yCB3THNOhn4UC1ZUyVchLDpftv9gCdGXInPN8lw6XnLhcEMrUHKyudkRR2RAJwx+
xlDItYTzYL+MOsW/VLgU+gdtR3jZ0m8aTtdXplujdiBQMYL1goG7LBIyuVxygTI3
UehIbfRBdAjm+MgHHezgf7mfUijDc5z6u8Xc1DUp/p8rEfZajzYF1EIRds16mFJa
fJQ0ayqn4j62gI1a1MtepQvyU+KH0d3O/sJT/U6gQHbyBn39bcM8H8+P7e1v0Ua6
pndGBxCWc5wsKYXbbq1jYVhIXObzfXv8sZjm2LpfyukYodvip7QZm2yReBVf9Gk+
czCpmfZpg8vbmYmPF+a+h0zJXtAqWlK1cGSWd8Mm3+wGpydlI5K6kupv+SkgKKx0
mFhnESKJOFmz6ofQelvpPFGAUgWlAXPcoS+8p8PDuf8r2A94/tknXVvwXUtGdI4S
0nuTVQDGGMoIsF3cKjyAedGyE5+aLC05OwHI9I+So/7lVliMPuIra8muBtbJNk/h
ch3D8Hjp4Q6WCkboe/UzXKmuk4guqMiAL6ofWg+LgnJGNuGoLFiPrwuO6YeDiV0c
bB/CeXaPf8gT1hSQAoTL5MohybgweM24CoUP0nlJvV+rd1M8FfuqmmXBioIn5IV1
sRG+x7OEAiHfufNTk+v8gOUUYAmzKiuQiOyGtuj3lVC+zoenvB6uub93TEwkVFft
W22IoZ0kuC/CnMDaUIP4zleK2eXMexsorP60bCt5Cgl/dnQOoOsp/pVXEMWTqms+
YJSpMtYDiZsqje7fM3Zmwxl/3Yib6IlgR9Z7CyZYBECxjJ25J3pScGMtZGZZzQEh
5+JmculF6CMX6PhdHijSF8cUZxv89GYReNypHA/PYnoU/Mo8uEg2sZo4piaeBO6T
5WrkdIMUYrp9SX/1xGeHcMDqqCfvAutlQhifKh8my9cpkrQN0yd0UQcX3xHIAELr
mQO49ZKtMXXtxz8x595e9Avwj/FbRnjxpjcOo8blsD31+ZgCWABO8KiiBhBFg6/k
ZGeVfY5vxdueZsVAu40D0ClXO2Xbs2Jyjv8UBMziR5zy/cQLg/2wKyWjKW5j9OsH
BUxibgbAgIXA1/UJ7wjKOlCkH0dN+XXqgRnBzzOK4bxAB2Y8sYc1/jwSTCKtJYi9
b8Euq6NRE58WTVa/QBdpIU5H5bNqoNnpwwf3oVJU0kETkCaQmputSj2lnL8Kfwrk
oTIIfrVaihqGJZWhnnA32xG4FoYxGtTfpCtfVDOAg9OBQyqa+zh4A5NbBVYbHvlu
uacZfeZfzBSZb5PR0DShOBHO18mi6bXg7PD1HFUiKAUnQyJErdZ5ISpfABTC1P2E
SfpGU8cIUQBteqZu61F9wtlqh/rKJWoSiJ02OQP60fIuTHRtajPp49L4e9U/VD02
EuENySR0ezgi7BYdXBhJ3FXFjRjUzIgm/M6SxmIYLtfyonc8AT45oTtnNyUw5CKi
t6Zs82xe1EFc0ukcvtTeyQVkH8q53ysBYVCQH9RIT+Ja5dgQrRmItH20xsKRSNAt
T3hGRkuM65LLblZOitnSpVITbgOFjRsxwgA5xNR27D02RforgLoBnv6YdpdXOccC
AQlFb6HMjA5DIjOR0OSKEM8INXDVjZexXhta1e1GcxruITx4H8xNIhNcmR1lrNuJ
lPEGRi3xgR2MWSHC4YP+2MEe71TzSW1FJGmQtW/7nC73e2Z8MQijPJwWNILfJgSj
+g/au7ztr87TX5J7vvEPtMZ9lOgsrEaMFqMO5AmFLF1u0z2c/mYHfevnRnRWBmJ3
hAYionAoK74UV4BKtCWgEuL57OW2uF8X4JgOFZ289MRF6meat1XBf3j76CdeBPdG
EvdFWMnVhHrH+uHo3K04hw1Ef5vpvAFEZ99/BAkddZu38vqxwDfwkO/T2VmWzAUc
98n+tJDubJ+Q383Ri8GsCxQ3wuX6hOyDP9DoFFPrr7P03UN4QAr/s5ARHBE9dLZU
+bqk9rPpoGQCoflDv6yHnEa1oshXmx5xnaZsHqel0KUh+yq/6NgVkWrrr6lTY9nJ
ynnADeS9NYH4JF3Nw0caA5XlgFezI4W5YTZDQPaQEnW1q0TbKqcVUz8nSlxhy2by
CSYu5UT0CDeM0s9GDsyLnhx0M7ocNQG8sMd+djFIK6AWLY5kBXjhO5bhemu5j9fg
5jzMveT4xH65+iZqMCvGFuo7sVtHwnpE2WhRXgxfQKGskXybNFagdgNdShFbRVzi
DNesR5HEEPvd63ZTu5BMOvE2TVN4ROlBGyWl7m+wedoEk4ZmrRohVTAtCT75aUEO
HCi2J4FHcO7OEWG8lusDSndZg3nNVEWD8HobQd4hGBN1nsw1Hgw9ZmrgMWGS3F5L
I/2MYEAvdFxunxLa7GLjCoygTcMZGWOv3D+fVPUmqdKCHVfxZti5GfUjYP/bit3f
aE5A4iNFNWPoKIRrx9FQB65vNKjHgpyxOdZbgqUH31/vQWGyj/60t6qBSWUvDp0/
tyThecbbXkXb6xOoUZq5a+mMSrmsqvlBphvVDQV2V/41Ty5iFBefVY4xSSQg2r8+
BKUoaXnT78EsS8ouyo8Mzcc3kuiPCLt0kMC39K72AnEW7Nx1vDsOAwfqk9QgQf9B
MG0HtlTOSi5NQ/U51fuaFK9NI+v+W7ijFi1ueRpShX50MRwDEE9wk3x9El/qp/Oj
rG+uOjgMmQOah7CEawcLkojmuwvJ/VpUUUTMGHW8mONqnIfzwgSKyzV3j4wMHihL
+0bpvgJF9Ss6zm87QozJkfgrcfdZr+fl3TViAZ5GvT/ERt5U1Tob7Iaqn4Asv60n
FEE2SqyJGtbw22gu2g9/3SZSMT4bmlZqMMXUxzTJ/hQ8kyrbNyPZ1NN7W0bcF+sE
X3jIKcQQtbIVXt6+vT9KrkzmHrpoQjT01/UT1OpejSZpNvFSeG9qilyxugOUiAGn
9vNCqDzF5qJER2tZWniZhV8XYO4Hlqm46IBarIytTd7SupFj6HHK34KbS5Y6dKS1
wZYT6BUHdiW/NXSuR2dD2E2l1dGI5am6Seb423GRiOungjvFtpY3P4p0DY6Bv6JR
C60mK/vwN/SzqzRFL56xM5foSOx432Duq4OJvjs1TxxPDvDTnAASf8uWliF/Oi58
0jLGEDs6TL6JOwp21cbSmp8bIsbf9rYGgl0Lao5/U+nIM0YEToIIBeA4nM90mEeg
aGHnyfJQyaJetj3aKDzeeiJxkFpW7nY+G5GSsLgsaVRdMvx94PoVcnEDWGFI3h1C
Y3wdnf8gjMZk0QLQVbQPSNTbGF2032aRVBH5y5C8qhw9Wib52hr/MY5lXl/mjZ2D
kJe81QiNMLPWj0I+7OzB5nA4o2st+LOwQGBOiks94SRvXktWbVtH+a+383xna0V3
KdiSPk9zQk1+cmSKG0vptuVV74+4fYOf/OJvWTe5ZKRpDdx4OLdbDEPCCYQ7JMkS
i+hxTtdvnfH5vOjG4M/3OzW3Ywhi639UjuJBky0Ohp9C/mupTFCquJBCzbFMBxUH
WzaY4lLqZFOuD1TS7/veDk0PYon0N4nkSfLgB9a5QU52yUax2ViPz0gn50Xp8+dO
4mTlwFtDTPg6Y7T/n8pD8VlzYU7IcmSVnY6r0msZaiukNwXMES+T9S49VxjwoCpF
blK//ql5I8XjYTZW5DZ/Yid2yVYuOIv80B8F/vU14ovel5aj9YQPaipSV+ltUW4V
TTvrtSlMghprJuBKVzC6PDVtqjWLHsMcIBZbxz9pamcbgRubQsTqo2ZLCUxdwzQP
jIxmhWcXKWUbJNAn+oB0nM6Z32Oiq5fzAhN+bGL+mQYlNIpRHtnKCGRgD5A0uPuq
0vVc/0kEkd9Qhqevx50qCu3+HQSTdmkeXXmRAPp767fkysLGzpaMFtMKCnvJbliA
nqCz/pPgxqghZlYTB399pIG4mLsUOwZrGR9CdTq4vAU7qpqcc2xdUtJcNg7u/DnA
MPtO1hTze9Yj1dKTVUh0JYmiJ2d9EAxU/uP0swv772lZEPZbnv3jahDKjFHZJyR7
16wYMv9f/zNrCkUj416JB7tBAuxKKq53SKsowY9OZcV0c8JXBjfONaS+ZSQjU4lI
0thvR3P6JwieQTVtnZyAQM7YsFaSf5WjkHYc70ToESXbfygebGezYoMIptBG3Vhy
5qdlf863tpu3Sbu4SMPIzc7GecQIY0PvaJ6sEFTUvWM8xs3cL2qAdKpzyyW7Rf67
/7opzYFxtmexilK5L0w/U/5yl9BIMmNZ2DoPiK6iKzqjEExWKXyqM2LqrMLCo26h
ucD/HOA0kK/yuGaNCQvauXVNNI9MPTRK9EZe4q0v6A9FfLHhATGcfPXFTfdjB0G5
FNzR8RJ/dTFwxBdhiXy1r3/anVaR6ZtOZ/arFTplLTCPQIrGHmw+RB/2m2ir7zAi
xPG7ZVwM+9ECbAK8FRmmHBBd/ubd/iGby9HKz4wpjsN9XYQxv0Qhbw4v1bMiaoIa
FIh5B6SucHL4vwAuLmUysxRurgs2+6t63PLsNhCJPYk0yDHEBEci+FzZUwOH+IHh
6W2briFZa1wBniSvtbbv0d0gednIdlo0QkbwgqU33+6G4WcmydWfa9jJKuNoivae
usg9PYn8InYFTsfG+v7pck6su4Td5bH1+kLSqF4p7VDNisI43H2ip54ekZuAM4+t
L7A7AC2WQUaI9quF874TRkdd8DQ0hrL3TjVqs6JKzobFnWI7jrR5W/aU2+cc8wNV
4nxgx/+bunVRkfCm3Tb8JscsI6QdfHb3xQ5pWbWx05YzXahjryRfHY+cwxBFYKNP
FexmcdjVtNBbItCXC2s9R1b3kX23DwX24qMfauzove+EffoqSOnFqu6rwdbD9U2X
macQihOokGrZprcOjLHFj7iSaFSqvjQGMyEUB10dca5+HG3zVifBg6kMrjbKMRZk
pt3QvAAIvrIUvv4kH+RthLKFrIL8ygprsTfH2ZKYHEOP1xWdWVtYQyLblr326RAm
HvLIjU2J545a4QRafb3w66cBakRqkNVX1+A0qP3qP0Y3Yb1q1DtthI2shG0PwRyG
CyC5u4m7trohCPMxlS9p9BHtz0vTmaC3EzCU96lmd5Kr/Wbjv/jY/T+oi9s550pu
biHpgTPgOiMPshHP6D5oAqFPNZT1H15O5xFRP7Uv7jOJZe0+GoUqgMWW9jnMLmuP
nz5v5DMScC7HXsLTg7+xIyuPyJcuYyQYYwoLVDc2u1T/Syk0/5yBPEx4C11kKI7C
Aep0LaPoAlbriiVIWs7doChpWpwKiLNCOv1VPZVjcmBKNFn5ZdU7c0vjS3MrVbDc
qukx8UqqoFvs5LXY0h+RZ3sQaVN2GrNfJFgxUoIkx3Gscqf9k1W1RVqYYrgMymRA
g4fn86CEn1xSsI+DsfO6EbnS+p8NWm8B/lb/K3G1aW1TOKfw3D/jIMmL7E1dwF/Z
lcb9cGqWTYzRgrpg8iZkEnjgYznvUNC0HQ8Lr4a6xOD1ZJNbkFFK+imLlzz1Flw/
q9xZ+NjTVmamzA9FrAFF0iAookLQRklCW7swpib/9laetz1Ce/czh5UjtWRq8+C4
hYoD3i9XZNfG088GWcCYJIkPY55NTgknIwrpvteyI3PxbZhlWG7/xIT5a7nK0l3T
jv6mXKXgHOz6McdZBZldl9tDMA/atXakB2Tv9Pz0eje36BQtxRakKNyon/x2viwi
XNCn73MyJPxuffHnsqNrX3c7RwmXpoNLj6rHTO1LTr7J3cZ9Q4tayy6a/4QpnNrq
HhUuzlMrAUGpekerziOwMVkjFJba7uyuaSGftxafbc6I3Al/0MDmwZTvVw8He1a+
/08jpxUxz7KBjS5YjSWNMwOIhyQG/6gVJLOGIv4sHkwsRlnUuQOhtMSTFmyq5aob
Tmyc9MJ2/6n2/HoZM75HxpBz8z1PVf7n8GQd7+X7+SCcpNBexn7fmi78V2vIupBq
HVVMYPcZ9NmzUNN+jChns1xCZjIhpDK/QLIjdH61sDYR984xZeoKoeSohnfMSFXb
PNqzYQBHJjVUzVIfweiQuWOFAX51wgmLPIcZDk/gm+s=
`protect END_PROTECTED
