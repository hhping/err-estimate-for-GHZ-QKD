`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvI2iEcZSGiFluLHPtp4e34xE9FpBktfhCxTmt+yh7ubPUxHEN5m1VwmaeWdGMss
8O5e540gltiOar3iqDXkE1MNJ9U37RSGEIrlgjoHMdslamYs4Vgb5hzmD82HnMca
XsDsVQi4PWzvCY9nHOQX8XOOTl+Fjhi3EwZcE7wH5Yel8GxONLuSu9u1JUCrHu0g
Q8CsM0YnAArEafqfxi0TmYRcSw1mvV0nqStKiu+1O5ShTgvuIzpKZdW7uPxw0Oz2
l4XhGnYqDjbVoMBEeqIuf6uzQvLrhXu903Sb4AlklZVDSbcXIJMHEBM7oXnUfzUI
HxU9V917/+xhwDIHPENMe7pq0xe3yWEbUfJzDofPNsl38Xz1zJdhf+ThcpSxikYk
CmUbN065LtUsG33qkbGEF9Y/My4Kv/v+Vvs1a0yAWZny9Csg0GWsexfq0724bSEj
qIxHPXc5AORCEHzjicAKUOWTMIvrFyrB3j8PRBbMPIGDTGqosIGH9qwYPvhVV8tu
2zSfk6/zRsvhudUD8O5PgxlfPxPLOaireSy4lgyudzo314LzOy2Qoq3nfDYinEg+
AyhaVbWZbnv5ZTv3UPADhatKqeuVnbQeFQxS3BhFcIpEs/j9S99redHWLwURGWeB
479RMJYJVk9H+UdLfWxTxneWdqORabS5q3sTYgrhQnF0iDDLM8qVQ3/m/DEMzsZx
WT5EDEvMfBtptI0l0H5dTzmMuipEHAYJso0syfoN1uAHbLcjG0BOzsc7IZTd11YH
Dwsv9dXUl1JCEpaTr3jaIRAAxnanF95zvHF+BMJ0dHwjvbsWqBhI8+vHZtifbM/h
bLjxcuiaNgT5x4nVCSC4c/HYUszWFm5RIAFFzWtjerZE0d4OuefWdTCFmRj18fKG
h2AbB7ZP+bVOkPGb7yBQdx7Zfb1YSaY4SiDqDA0vyZ/1sTI/cynwQsYutojI7dj5
sBYGLkgUKUjtMGyQjMOctg==
`protect END_PROTECTED
