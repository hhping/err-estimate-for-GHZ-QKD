`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1jjjRmKo7DRMTXmZO0sIW2e1glfUyHwfVe7V1UWj2Tz/LTAOvQ3pysn04UON3mw
LDcXYJLqBBVHN+T3Uos8APGqeIJUF4NzXAMuZDS4iwWQJlYfkxNVio86vMpQCkvT
nGtJK4/kovLEaOPUBEL1K05ylzOmIP8nwiOEUe6aR3Wu7VZp7jwmWDC/7jl7DGaZ
onsmIt6cNIq6HsvmJaHEQqj033jKzm9pCxqbYU7cBGMHNAfnzhXlUzcIAILG2h/m
3FpNEjtH1l3YpRogj8HXKqdD1jHuLzEe9HV0MOudHdDuONV6RnxkWZIr3sG+pgBj
dGD8fx8PshK4EndDT9lJyCANzzBgtnWEInJotYLotdE=
`protect END_PROTECTED
