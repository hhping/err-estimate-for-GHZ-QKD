`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CaqyFwZDRcBvHinLKzTCdctIzbnKDafmidtWMSaUqPlW1XoUnNu1eJCn/FiqMltC
UGioeZY/y+R5uKTtkbLKcpsFKyjg3uwpAue8KAHnXfbMwk80ZtJuh3ZQu2VEsxBB
ch78RFOYxTx+eYDBlr1JqWqn+n2iC45TLotGtM1mPeewbwrdtFLE6CCp/KlxHSUD
El2JqcoMMv9sKL21WkcotXTIlPJE9sQo7KWYUqXH6lkezMrpMPTeoWHKGutIhvqv
hDOB0/MAcEH9EvMxaJ7OYQvXqTGWvKJtV3zfVAUMcEluXMeT+7KoZG1d3q5C9E6e
WIB9iXBit05f7+NLReCoGxz62kI8/soLWpW+PcbL6tRhXnFd28U1WzDXMVuT8x6g
Y3Rq4RRAo8cCpyx1gx3xmqWXjJpj5H/w6qJJ2dLi+7S+v4MnDCk+YD0aFMTccmZl
Hir9tLUwXjEf++ZpOZ7sl1mGnqUKeIDzgJ3rGMRBc2lftGmlwkAP/VAvVeRhmQsg
1gSspvpmPbk/eX0SAqr5N9p4gFha+oIw6l1pd82u1XrFCQ7SEtZt8rJpZ4tCUi0r
k+Pp+djJHVK/oxA0gFxLj2xfHuTbIkmJwNoDAEqPfKw8Xl0xVMoOgEzofiKYooq7
EjsmwHefRvbHVhGuRgC1BNXigZO/K/WGzMloLfevUYrlK1rA96YDJNZRqJ5Xwnl2
ttwPftZN0bMnvkgCoiesWH0PGUG8d5nrTu3gsysNWn+36n1nRT6lKfeyMkD2P9/P
jozLeWUwYJNOLkEXnGUUJPNnrAUp/FSsMk2fNa5N98zmnvaMCTedkctxnASAJW4S
crR/XhE5gaEFxqxcFMsHdoVBxmQyKNEh63VckskR8Zjz5MfcPEPE0SBXqq3UwtAT
LpPnaI1+YfkLf2TauaG3ei5j9w3KRsHDh3nLe5Tam0BcjvFMmpGVm6pAOW1EzEx8
9/bX6Sn61ZvfGxFHABlroweB1aKlhsUq8UPg6tTGXnqspiXzjt01yk0UeC9NpgQx
I972QQlllycVS52j+FF0NHWIwv3rDNaE4ioO6btonVVY24prYAE7BaT4weK1MaGf
XmMTIrOj8RiGwbO958lHtMLHljrJxFad9iDUU5qHv2q+EOWJTHC0HDjVuTROKg4T
6yMzkWTxaloLnHd/Up3EHLaIbhyd2tr7mlwdAdFOXP4Gtfo0P0s9tXPE8Uq9dlXA
56naKLr6jcwREgtyvMloMSo3cwcUH/D1sFCTUdb2emeEg8ZN4lVAC6FVvcEgJa6h
LLXmU8rtQ8Zoq35lXwyGX1/yUGMr4NPRn8mKURGdb+Y0V+Jx85zYkf1XWVfwgBlw
jIPlgOSj5B1igXekqoC1oe1pwHsjEhzI1VxCgHy9ZrbKDCrLe5zD5hUhbXqx56EP
lDQwn5AY/c41gFSEE8mst8alRVpiqvc3Af++tFclz2THAXDy3q03ZJrETLGaINMq
zCsMmLaaMqBI5QdGCIFAAsU1WBIxii4rNQN19Xxxu9jMDD3rZX1LXjwID99T1f86
ltmU7xsDsz8zbmxM/53G8Kmr84TfuZBAdHNnpxYarBfG/9Np1jCD9EMfBGeTvxYM
EuxY5HMe446rJR+cHHwUKkiUTyba+yhXbEAJzPKKXvV/vb83WEfEwHKEs5FjmHdY
KQ64wbf8tzOpxq7soMJ2l0p4i4F3RRRJxfAB1goWsDhWgJ37mcXY0JaQcGXvA74l
Q9efXkMugiDBSv9NyalnCqhAPkT3h+CVw/TnrW/lE/T6hB532EF+XTme6Njo7cSb
wOCPtoYVvYsYbB6CRrOmpSFk0WpOefmhGmRc+sm+nsBhGEqxUfFLS0aXRSMnwRzt
bjVCGUo63mVr47WMrHVSld2KDO63PTEEUsU8mt5SpVrcZtcMjR5UO2BFwhzS4M4O
y43gHg1IXxFHfaU/ynJG8pvNfruCB30k6gMhyR24NGxpSsZqYegoGJVnsdfZcZhx
O4C1rCL11R4nCVwE0HCnMTVaJAZ3k5D9lCSPi0sC4upxhdVEL/Vj17xHbIwQvnZe
qkB9XUfw8Xj8ObTeibh+ymjoDv8xymtSCq8HC4g3iDeoHIvhGXlI6vvSPEhVxn3Q
BFY6t6DlbWsbkh4dOUh6ZvUbAm9i8otpIFvH4ih1g0yuQr7S2NGy8BUaJMto2ElL
a36Eh4V8g7oDh06tD9/r0R8pmpeavENSPG+JiMX8caL5jW48/wysSZZIjKYuFDD9
+YlC6amgciO0KVxwVXz9nBuTlxqYbGBj6AUvg64RYzcRZSaIvZb0Trl7u997DLc/
GEM477bw2A/1tdtObh4p9wYvqj3LhuySK7/cqw6GYlzSnynLq7mpVZHsZA5ohZij
IC3Lv3zZMPKt7WDmuhL3a/oWUSany9F9WRHM0Ug7kfA4Y7lGFvTB/ywX/hBznkwY
8pHBecYdkAIf4LvJ82rcVv5CypVZDxehzYvEZQw2qAVHeRBFIXUhIHk+M8Qfiwij
bF6lZP94H1NZwx9OZZtMxRhR3D6/ES2eedd3LA+2sJEi5jx2tpG4oFvmGwpzHhb1
PkeKjPKdUTbhH4Qgr1MEldINrtaTy2rN6A4pGz6bFW+E6UDtb62IhqZLlHs4oJFC
B0A1rE/eZux3Oa6b5GLoMmQ0RSDVocFslhpJSGBK8Gruu5BTCxUJWU8g8RKYwQMT
krEI2Ihh/xIvNhZ2WLumxuVPuuOiLCmseB8Baov4Pm6BZEdnKDyOiz6rMpkUwibb
LaQdJg3JtD638ZtClSCkNhlwCbLPy9vSnOXwy42aPpex1o6pSHlEsuSf7o75Cobg
989VJQNcU7tMnoGC7xcaJg82EMpBy1Mo3bCG5bBHFqVbB50xXJlNI7xl/dZQAYnX
W0hQUnNTp2TkjtYCHRUYuDT9XacHz9HBN44DzpRg8DjFiKaJmfwz5iEq+zGcX2dW
AKBfq/a1fiXny8XBj2YuO3BSsuV+QGhSk1aWqe5L50hgz14SD0B4SmpbYsNZ+GQE
HFWf4eS16mDOBAingr3GC48pB69oZl4nOmMYlZWRcjJIK+v9aDomvEnUV3xkiEyX
gvgibMQ7c4NAz5ZRw6A+kGf5jA592YQw9NqOKdasRFUXY9+BXfbhlHs9GkSl+98P
O0KHdAMcsafoAG/6SaGFLQy6kXo0siU8Zud0MclFPmcVxkJuAwSBeQRMjv4MBDMC
ZgC59mGST67O0zJ1dRxJuedGLBii5hWBzyTjFmXW2sTvSVG7EEVP5hq8GpUy9U0c
8rha9aHEpYPWNcChTjcqRgRLQc9YY9i2/Ryo7UWkTbaEh14RQrHknN13pPXkHcBX
Qfrr6IFI0ZK3IvoLNVS4rhL5AXwLXoL89bbnVOvPlFQkuY/cdjs+qgeIl9d5nXf1
2IFK8tflEYFdCXHY2Xmpf2/63qVQTGpyb7tDInw3fT/gWbUY/XSBg3Ys7B2Kj1to
JFgybAKVR7TwaPCTXw0REvyw00WC6kMbjNKEpyRZiMwVyq/wraAc0yOHE7mAwjBB
fcqamtixG0NEqv8OPaKXJqHxlSG/IM/YWV2oCiLkbRP5zcZdV/+2fughFn13Hqm+
E/B27pwAznQzy5DuDwDM9JpdtNXv59LxXhF892/jbeVqOi9bYDI7+/wBLAWCWm0q
pEPwXOmtSsHCS7Sqzl4ZS6UDc+l4onBQgv2CNSXvGxP30iu8ux4klCHHryuN+eSl
+nxg8AfTEDWaVXv0oAxqHUvvtf8XcV/8jNbeDyGREw1gnSrhXQ83iH1vZlu8/xGQ
9PxBxNT2FKh4qDDkmvsdLMhghHM+qW/4LmS6SQxd11N+s0mgDXZsNMM81rIDjpXa
oAysYjSJe3FsKV78mUVCxW4PeJXWirK0tXUMhwuAEPa3gNckpfArOgv4pYMbVrsa
RWFP83mjjAIo0OfblYnGz50Zrw0Kqgb9yH4KDXL5QTRvs6YU+b8l/TlQVkeu2lT4
FvRo8ls4Ybizz7WoMIZeoaRbqdQdHlQctUtCT+47mrbRCZM05+H+wkgDJLKSjqPy
mFwt7V8TfdjNJuHpEP6tA77NL8EUwwb3IbmB9x8v8KB//Cef7WICrZafC0dHAb8p
uHnx6F4VbkfdflZoUur8d+Bsg5kczIXDnEIcFa9Cz5SpghFgS/+7P71t8LTd5wHD
qsu5N6xkbmWPY8pKN6vWzLxOBbowRwSEi6IAqdb912qlYT2JUjWQf6kBPmn4XodG
BLZaWUsHLrU215n4DZ6HmiDcYEHHmS80xWgjcdLIjafXyoBMR5+RxtX8/fLXOnnD
sYwGq/n2Oqp2hJjZP499pEH8MQXgfBU0anzDr5+0ddsGkK/Jy0r0CutpaV7J/lEU
dkc/+WtZArnsXQl1zkv8585I0+dloOTFpnl96As1RWvLODoDlQM14T5TkvYfIPpN
nnuFzR/zyavUBznYP+gZ7vLW3bKt9l2W5Ot1SLeTCcsKyyX6gmczlZQHon/2oryX
Ad2iBsRBvjSZAb1yzMPSD4grdq95sHVLhOsuLdhT2F7rEF4yAmDUfvLtHSMxkONJ
lW8vmSTUCsvCsDG+1mhfVNQBOfxbp3FXyV4f99ZjZV1n5gAThThBv8dst21hTd/j
7rCQ8rHUeOJGkzKYHYvJi73iKL8uhW8A4Y636ILG2bqtGXHpD1h2FV4RQ+CMAL+u
TQqgthSaXNbTOTg6tncyWbmlJQzZpeZzIAIMG04McYA/JsW+Pg54eagRzPY14BUN
RpL5oQtbh344t8lUqUxTeylBj052TEIshV0ib43+58WkK+E+xIkdKuJTjI8Y/cqd
1Vw5lcQCt8DvIhzLxp4YB40l+1qJ8DKxowU30g9osg1UgqK8vkrC7HT1jedB9lsd
GetlrJL/ZbldV8U2I7BUaB15ZAfz7hzO4rn6QZgaJW60WaHZaLHwVm4wfTi5nAx5
CQS4jLkErbZYBvmFmopWUXcD+B+IIvXt6onL4FlhlKxBjR9spW916b9Yc6WIXhgi
+EueVeAI4tBBZwdeaIC7QylqxuHoSZBkrOzqZ0NRgE8lI5qG3x1KEwZrzXjWqLsq
HLyg+d7KceW7aORztlWAwy5NZnjvTjoFBxduuWKM/N+aRd3IqxcuPl+J0mUmABlK
NBmWeXhHwTYk1i5tHBTi0BkgA4NJCkXuGiE0b1DskqaFdm168wVy+JjVYlphFHw8
JtRe8RnXF3GZ1Lxk/drpjK/XrbBYaTTDknD2oLLG5fKotT/AUmkMkjuGAxVt0Zuk
VBFbD4pQ7TVTNXl7bjkcIzE4hkPb3lvNP0MZaHtTIAl60WniuyWMD+7It83yMRU9
ybivMM6cnC6FjapC+kzQTzmcWcyvIAZCHqPkuLmRhqOhWviD8mpiC46CmxpgXpSv
O0Rf/AmyiuaS0BQXtpDmNkPubg5kNnBft9Rt1j+/TqnCKCsghxJdhWydmR7Lbfc5
IpojOHh5vC+teAXmHjIYKt4ECgBunIiBtD6iNCAhtc1+OmY5mKJPaUOq52CpYRSR
+FL2p7+cYxIDJdKGJQuE/japt1cozfDrtDS6XLXqi+V/CbQTJriLLP3kHu4074Aq
Ewt1S5yfG1OtB++8R5yTdq/mHRlOQERPjfSqVVUmDMBEkHc1yJTKVqRQN/KyOIV0
kaR1lyQs9Ufb6K+JrYinA2nRmtmnvVrRxzxU+SSjODIlkR0uJmeMPgEp+cAsYvHy
i1cPeIwjm1AAqEkSz4nk3wXl7+d+sLB5hyQ1f0U2FcQKwTZDzHxg0/u07L0/zytj
arKlTbRAO/+S0/5kcU3LKbHxkHdHRmw6zAN8J0TFVHfDeyp7Us6lyuYZ/HVLX6Oz
bVoeAfD6QNorWk3JXxcc8CboKBFmhgtgVWi4prvvx4zxkmrYkM5Ahw42hUgpxsVL
M/h7s9o9dB2KHYtUlDHCdJJRXKxYYX4gucmpXNWPDED4A+cuwlfK7EN62xc0qjS6
FpH9j79GziZonsYO4ffrbXd+9R9D/DejxGENILVY76T3qdmryDRA8X+sHOODP0rM
oFtlsFF0GHaG6CnqI9J2oiaw5QXVnuEqXcdlKKk2Ow22qj2W2R1YB7/ymTeKSC/N
mI08NC/S5CXEbveHHelhu99w1YYpW50tq49wkFD0qAD+z15B4ubZnTUegmJSMqlL
OLlfhck5XiQljsIOwha6mXSfcHztWdL5Jk50V+TDjdNHqFAvTdrkr4QkWeiC8Vry
Yvx0uqM0no1O1k4XJDm3p6sphNNN457inGjtkRLzP0IgJik3QHv9+2AkJ+kFqQlj
z8PBT/UpBP1/UvRrO4+8Jq71yN83VYEp1A0n8DaP+bAmL5w3j8bEN6bf1uNyO86p
foBbfj0/JYda710PhO7YjtPvIU3Np+mlxvvCT2myoS9SPM05hnqAYMrWgRUPa0yg
ezT00VrIBxE6hvGxSrnnnIDtLFIDIH+1KHI19HAtxZY=
`protect END_PROTECTED
