`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2g0PiBFF91F2HXGNGxzsAP+TZk7pjUqJlj4lk9YxJ6nvdTGjIT+Y91BIx/bXDmv
X5QGlNYybEJY1e2B8moIZMrbkpsNFpb5fPB0Dm/7uaQv2MvUKeRVvFtDbTHnDMz0
hMwMjLiIyw3i862uvWqmgolSGdO639zHCP7g5S9P/dTlAphQ3MnDGBZ7rIw9gzhr
NpsK9b8sWKYLPqBMoPlrPoPfsWr5jNVqW621fBkVkNiAE9+IeYT7ZGCVXD5sL9s0
SxDiT9JYJJUu/XzqAWKawa/YJiGp5IvxJ3DRjLcNWtrhSrzACFHYCFWTZT5PvuJ/
Uecfg6fo+98IuOnOP3u8x8WvXqzWEjjhdo2zmhm1sn50udw8qU2uA2EJf3z7AH8C
TRWbVMGnQ1QiSdorW+6VyLapdPSM6moR23d0qEOrLMV3AEUnUkLljrX9e56O3o/Y
TW+7un526qnEnFIRxklAA5RGLA+xb4u3RNfw+ZCmLOWuZjqzKBFQQ+UYb6VL0Qxj
4eTPLXfn4bTVXrgx54GDQ4Bd4AC3aIkWm8Gx9fFMqjrmfDp5cfKM1YBoX1DJ45No
CxhZni8cFYvnJpJfZlaDE0gaoDore7w4pzGvyJKhm/8YQ/T4s8SfDkipcWLn6Zna
tIo5pLsuW+borlyJ4q6k3STm3KjvFgtt1sgZzP68oN2sIa3uRl88vpU/8blA/mfw
/CLkPCtIyQhfEU6Ep7bG+CCnKdN53zEgf4b4kXQf2h4APAcqjg8INSbjhWZBezjJ
GoVNcAl/qb6PHsi4HI2LhSGd8SFCUcr5suKjX2GRz8nXfWU70xNAUPlp7xO3NUsa
fXKT7Qb+Opxm1MRsZwrg5KLa/zt9jR/JFTI/CSMB+3UMWUqej2QYpiLGz8pkmspO
1y9hbxdl7IMMg8WyMNhXjceFwTkT+EGTvKTD5UxfHB8=
`protect END_PROTECTED
