`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0XJ9lmwsRq+jvEQ5LDmNEbtHPpm3RnescAx8zLWPRWm8Tg3H51UyhmJPDs24xGh
DRJd81pgzWrEG1Lmt4AwD+KWSN7uJ2p5khXKvKWEus3OLC0ReWerC4E7WV3A6+TD
uK4JUWGlE2mktW1XU2LjL+xgao69Eb8Pg5cJ0LmL64w9ennBbj8n/TDWoTmSGNLW
PaNb2Vbg6aC8NV31Veh3l3ew9xf8QynR0cJ8vK6bm7bbE3bDK/bc4SOhj26to7tf
gMVI0QoIf3/376O9eJF1gG+sB3ymfXJ53NK5dq8N4ep1SmmXeVHJ0wGxuA7quf9o
k/83FL8k3Z3jTU8a/D4CN0zNfaaTDA5X11qTz1eoPs2PX52VwrfxN6GKvjqOS/ip
ogzHl2BdNf1Px3iOy3OpRiXktQUZl8KqtJt8qZQGK6/bDUi4pwBg+W2ibkgRR7PJ
ydwzow0/KtG7+MBxIf+tciFVupPuLdc/RWRjLUz3o7f2dP1yfoMzSBZ+mFI0M/Hz
w0tiLenzVzCeNZBAls7xBgnlwSINyYyPWAn314hYZb4m1L8p6PEcm0+Je71i215+
c2m/nIj4rMA0PKi8z9xVg5y6h0oPKwx2Nz0f84UmQFj9EcIzzICbfj2Wi01uWCGQ
YsDscQVhe1jiLCqNgZmGzw==
`protect END_PROTECTED
