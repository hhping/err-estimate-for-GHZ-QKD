`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ZkkV91TaCrgZ7vxLwbxPEedrk+B7JV7aR35IeWq58AMnoKe+dH4UVdQibpZcTg4
YiNNnFAsVWbWHhcb/5nMIF0ldeQZybDVhrKlsMag19G3uFs7ajSgPe5Ctf4AIZgf
+XKJ60EfqEqEsUZfyv6R+hnFm9hY+mgnMtTfj9M0ma7EH7oPH2exLOePIcgTMVw/
yBDdbg4RLGiE7XoDOgYfV16sAoT2OlCpOCpORgzTEWz3xQJCIJOiTKfgEJHdLE9Q
rCnR9ONZ99eF/W4BVVkGcBo7YZk5DdRAVQ9U5wGv/kdVFIV+4vi5XzNkSMOV1jA8
y6+gvD8M/UEjXPHFTPOxauOZuVRdIr5d4a/tJL7exFwBOYbKsvKGGrnouNW0wYL0
REQw3/ajnSojj8X8042BUoM8VjupQGOPZqLS/lYN1N5e5yjuYESm51rDEpJWcoHt
sz0Zt8JpjpmBFHLkvk0hjbfIiC9mbriwCPeiR+/fwtmMuENyt9TIls4qmTy4R74P
647xWE78lZC5oyhgcPTeNeOMUr1p4ox4HC2S7WLFg866DGiD4b+2HGNiM0lwgapP
25XR2GWrDHDbQgUbzRVmHMNRbA+VbkyK8tLZXnxNj/kQnun8Wy6Hedf0O6e/sTZx
hTHy2ubFOKJrjqZ5+S6ci1fr2rrawaVoQoSA+6LPfkokP8JC/pucluXbbdWow93y
LNXgfSFKdiYvdeNjRFl5WtSS6Y6bZ/7cgRpLfxM/gf8QGVePl6aYW/7i1VFACcvj
4zVzSrO2ydFBHauXGGDvL5r5c8IdNaMJjyJyVikL9ONLYDllc38lb7WJF0c871kh
WbciRkotpD9VTOU7CoKy1+oIW73R0E4OYobhkOXwbfGZDC3SZ0Gu/5OUbdA4L4hm
u6Cg/yyOgxczYdVhBUR+DCp74ylhPbAyExkdpHQ/EEJZky2EN8rpQ8MYF0car987
5FTKpM4Df54qkOBCAvXHITa7SLUG5f1gI85VZzU7HJaSTI04Jf94ixaCCJS4H/sB
WKGQGh9ZkNH67n67yqBtWq1InGwiemtU2Baj7s45Ni57hBU4wT2Ox8aCB7bwtlVl
aaz+rAajryVwSoK/gKP/0CftiNC8v5y1oviWYC22OaIPDDK8w6OhALw475PVqZ9l
IS4bJPrqIkafxW96HcaHtSIyBPdPWvY4rGMKA/3QwrK70i26PN6fdQlSdNf0dNrc
iSu2FDudYbt38icuxi5Btnjl4kPEURHG6eXSOJHwpoSXV9aPIXVR4Z/mP6OPWgV+
iU/C8pPXKvePeDCVnbYe2UVkhLxFU2euPI9dTDawMYuvHSCe/r/vyCw8vHur1W6/
IUQJKP1UK6HJ2aRm11xJNCMHEkeZ9uHa8ZXYMZVeHbs6bQ5PNv1HOlsm9M5+ZGFb
gS8HeNW+1Si77YAaBf57JOSeYYZ9Uzkxo9v15Ybi8AB5ONUkkhknRaj5vcwavez3
1AoTJKivuVlP3qHLKUsMjQvUGr9fPB8DJSOVWcL1KH66iTJj3o0RrQIfXwTsy4T0
9WtevVTntlP6crrhEiQGUKufixD/tOAEpD4esmfR+W5WSjnBxjYyxYfPsDORccRo
UVOSwymUSjamICqyRhUxkzxNwBWrL9lTUHZn7Xs6Hv6xkZ3Pd3ydDRqLeLHj9D9B
0FPmrDlsx/M8r7mZy5uCXI0++/VUx0/TbN/+klTYcjegqZvr70cd1kzuya4JBcYi
26DiKYSUVYJdgr6Cyk58daje9o+nfdVCCWT+2YE3Em2sWpOmQ3GCJEgo0aT4PK+v
HHO9IIyCX8mmqCGlv5lh0NA3HUyb14zZtXG9hRzmaoUSokieapwJaP5Z8OvTLcew
3C1rDZ71tKt1ubfdzEbdNKIJA1SCyCe55T7g5CVzkViyZdgo3zJVF/YpRfxjthrH
FdetKHjjzXCi9HC/ndXBlQZBB+8LTXhqU2rOAtPRUUokDquOngh1Q+7G7qI/IUu8
Jz1uHweFzpvrap6Ceq5ihR45RfKKbBCXRWDKhxTSSBEAdX6go+/mrXFfxPLU64PL
E13tY9WCNqr9tSXKmIr7O+Ye0IlA84yo58D+u2hTLLPUna8Hvo/7dl+esGP4LAJB
a+8ry+40mMbds1DOar2NXKSP/wZqaH+GWIVu2h70uE25LQMlcwVubWo1CrNORmVq
ehrw9IjYs/+t4HlPW8SfAu6tMTwTYdqx6CO8d30MZwurkTBjzdPqQ/1ajWIljMRb
RufxAUPE72jxGIZrSD6kVPYVhzRHSwCvuArtvdnuWDMkDvywWwNBL2BxoKJQC9g1
Fu2HstOMcr9Zd54mxFikoB4Akgy+W7UId74medXDJQRlgkcHfHAIgE/37H07WyVk
S1CR9tlkm/PXvxz4I/lVCWL9tIbbLqNbSyZyepHhrcaGMLqKakxyXgsCLBJ8nP9e
4osS0UMBPphzkwFsEZprR0EdsdV0iog0rIvSCHqpSBqeE6PC0q38fs2Q2B2PJBqs
yEPgKPpo2FQwoKea2UhyA+9c8WrQQKAtSVuvJAe3ZBMDQEJMFoRPTmp0m7lFgh4m
oPOcXLId5drqGTzfMHY4dOj1y2N5ayaQOcCa6yXMyWT1bypUoxUxS0MryGvWYW9D
EgHtcCeNAM6O7689hFJeV3/npjcm0+Ic8lXVtjWwwE/3uqTzawQRGuibCLJ9OxpW
uyU7kkA7U29eM5MD4Y7gWlzfsDmY4PxDf/gKi6amCm8N7vukZkfo7IwHiv4n7/yy
3PP9c40+u5b1JsGEFGL/IhcS0LFbdy/IS5g8SdBQAo0zhsePXs+0QMAj7/i4viuO
65ZD16wSuMhJQeMDvEIbPAxECBj2Gv7ODD7E0ls+bQjZ78x1Fsk4FtPH0VNFqeTq
wOAb74bLpUWULTM4gm2ZWZ5Gs4YFCpFwWa3jvJIwn+rK8s8L0+4WlmvSktHSRHJK
aaEUPFA4GK5XiZrCI6DUi5OPr/cF5QLZ5UMDP6qub7gEW5lw8GtjXXwGtYa/ZsDZ
xXnaOQc1bz59ZNGmdP2k3npbjoNxjEwRJ+fR3aXCY5uZeo+EfJf+hOjQVu258BTr
tldeFMvAqdvkdRzqbJBAjWfkX4cuLV4YQy2D8kKIidmO2tv+xmd8zEaiEOxuRGek
Imxy/Xyme7W59rauvBoo+ZLxUGNtmwCOIyFCx4UnJMuuKA6PAClNWMZ2eD7qsLhP
jJYlFg80/f44z88iOvCXUc7NhjFsvmRQKdkGcgZvBhHmT4sUebEulOlEpG0bU/AY
OuJAM3/B5JsqPSMtt73cmaAzd8jaAqe3M7Yg+fbbyP2jkxzCA5A9+R8HoS6vLDkJ
oMBVz2Ra+Qx7ESZkLzGwk2mmckaFMeyGsv27BNIK5vWVgdKXd+QnRYjPWi4ZulaB
EhUfxeU8GAwaImz5ceZl2W+JUqgT8vpEyAi3LbWDDkFCWBuFyibyC++NPljuOkKf
fiD7AF8BDHNNM5AzhdWQaqfmjrJDvSrbglWAM9gWlDVokve/9sr0uIDxXA6mQ/Do
AibTM1p9XnqID3XwPs0zLYNCfi7GxS+uQjummhGG15/RqAA6Z7Om9RBnyapZ9ZYk
TdUtRg+npOJxn1ykElf5mLnUhcy1PEjjJsXGnxQD57Bv+22D5te2kdqnqnmESFIP
Uv1xxtvmbptqzN/6v83RUf4IVB/2szFKgYGzUIKWe7Y5d5jGuWDtUW+pcj53JgGZ
U/gY6h3ntbDs3M2jRB5kLTPvzQHf6ogWZv7U14gSpR/O425kV6oG+XxtHjiLNkA4
LnCANPgY3q5ts05CCCcnGfLIcoUBehRCvKNl07qR+/nqYLEVZjTvlUYl/qAEwuYs
Ol2+SVHsS89taLFvJlr6Fwcgki9wOglX0+JzU4Wmb8zwVKcoqSFIf2Jxvq6mhQVR
V6ghmQWXdVhwNRzJ0fwFfYt8bQo4SOzqiCfvGwa3MWqfXgV8yAGJ2K+E2WseK5mt
StKc2C3kkM7I+488poms6UxymECHqbTHV1CCZbUXyZjER1989bulmyVP5UW/bsxq
zPB7Wzk5axwG76zKd/0rPzFL+r7YepiystEaAyqobuKJuuLl4gjQK0rCBNRZvtAn
9UoBKwgc9Nqy+fVAdjwie2gg9rSFZ6WEqJ7PPySVC8/UrXfB0docnrFAJdu9oM56
GdT3XHcgDVjj+PhulB+RvbFTJzxKwSJXaQQrExQuDWNPZw1NBR8yV6UJ8lmooNoB
QCUKOayOF52BoRL8OnUtgNW9NdMWwfkcPaYAQ6suR3G74+G60XG7h8mlFbYlHtIP
DPCHcZK4rCm1z99ulSkccCZRdNkblIf0hrG7WzIub+04cEuRhXxS/++2chKJuORP
3SJ5pV6L+lsHkeMob06KtjNPNoYgnnCmyOvHnl1+yNr/DJIduE4D8reeM0JMMh+0
3xLGeqoj95vV8/xEGmvyiL+gVd8ZCvgWxcN37V3Xuw5Xkez1DQyI0uoP3CqgK5XH
SgxEMLwANAVrbjHfkgmuvpbnoFvT/MnluB9rnSeKZw9i+IKdnxvum3xs2hrDVo0H
xXi9qGzAf39WWaRD/XYotfkyGrGxk64eEXltuQH3fyVIpwYvw9M1RM0fPmpolIs5
PDg11qeGdlMw3Tr9bazhXjdHJbhpkTDv5kpnn3zbI1Mv+loUQ6+DQNCuhGjAZT2u
SbRL22QFWFANsuoHcb0UeS/WX0gD4x6oClrfKuBSQ9kEaS2JxPfK+DGXZ6hwgBdc
An3S19W+7wgm2kjT/kJURKxN+XH11X2Cdhcqvvc5YHG6KM0N5FwSG1XutFbHZyHb
aqHL1MTqQ0qb8hH9DSx7BYnUkoc0+TmzainxyErEUDQ99nKcYoMUKnoMuvZqxrdj
hwuHR05rnTE1vJrOcBmaGNJJ/njPBs4HVUqJedoy0CUSy5s/egUU4QEfxkY3vkd+
1hUNFX5TfTXuXks1dxoEY0SyZOjn5xQroHoHjKy3i5B5EqHSIoWEDdqb1N97ewyC
sW8zZMa2cCZP18V1gIbZKVBljklznXlnOn0xqFGhTiyXkLlha+HIVrDgisI6ftdS
PWalG57SX4vXea+O+77bKfORSzWE2FcQmHzX0qQ0slL0Ojiv0dh1IliZGId4H4+L
/GpGuqu9PblEIavT53KvdDCgPOYy5y2nWuoMuwbhg9rvvlCvTkc9T4YH4GVKssb/
CaPHyQYKiC+O5AcHd/wnB7so43WzUiUkRmLjC4vv4EdWZb3/RRERO67nvvQlZ9A9
hkOcy7aFR+SqeEutPVIcae48dm6zKiuJ4qKHRi1AEb9HGLHPwpKsV+zNf09iWtOd
1eJv+tVp9FSSdhZylJvBpYkDYWuWcxVjEbDC2JltwDJOKZ7Ar9JKyKtD7NMc3HbW
I6YqBCDekyphd/2r1jutnye2kziAgysU6sI24Bh+z9BgulHJlJpgbYPQ4/2kiKax
598r/JEzWpCgJGoIMUs2+0qO8xhvxljobe7iXdIdCwvif1N0ygQPEoxFH1qmFBb3
K+QKqKvk/sfAelrLyfEo1VKVIgXBmr97vKIvlz/EYbDmFMzJbG6WVL5szrg+pZkp
vRSgaszWpZ7RCHIZb2S6eu9nrh+59U21pski1+yX3AeDen1yg/DcNnfuPuFmKcN+
15eFXaLZjuruJ8c/zZKEUievQw8La8zTtVOdO3J3dzpkR0gWB4eoig5xSEUYz7MV
yl2gCmK2zyLShRFhVDLrZytA6sM9zjpAxxOTH4/7piI=
`protect END_PROTECTED
