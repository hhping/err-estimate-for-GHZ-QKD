`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gH4XTgvk9QauGCBGGTwrBmzdtnSWBwpgKCV3dnhA6Uxtj4JV0lh+dkLFaKPJyOWz
3splFDPRLxG74zCtkyV+brGAh+77gwB03R/1fcqLWMILJJFQIgFu//4rtTzncmoi
KaaEgLnzgX1oCyVykKg4AtRWZMDsXZB7vRiuQVit7rpV7xn4JIXCUiMfm0J8Mwkv
2veslMdoIxSJXiplmioTjso8K6tOoyz9ve6QjLlJH2dWIeFACtx8q0gEFG7ALxgN
c7SLSprKJRQ2LPQMrjuH7itzuN3MbA26ZJmzZNCtPfrWsZgVIYs1sveltj/Uim1m
A7+evTVxq69Vd/V5U/bHyYForUZaOBHfNVwQ5QPqBAxB7dwmPZ4bhpMBL27HQloY
FvTeklqSNpgN9/D2MwysM2F2vSRyVYxZbTPnD9ZM6TJDwTxG7U/oI2coKKrru0sN
btud49zbvFQd83CAgA84uOZzCboJWBM92SsbDuvinJX7s/H768uN/upYWVqNdV+s
nJ0TvjqADSkp/hffPt2AmFHi+u3HJA8pFmu0Mei2jOlMej/BjBSeZewyGTCp7MfG
TWsoXmmPpYgdEFuDre5SwGPQ12nw7KV5917aoRZOk8WND90+48thJkHRraCr2A/H
4PXKWPWMQa6f+H2Ix9PcvDv6lvICXDGRK4DagdCfvGYsfkjAVSY0myjzBYFvC07z
fxD06pg6fpigy5F0Y4zEiGpjRef4c1VnYX5CFBe+XaW+xEe9kLPGxC4ZfGqwRXU2
rueB0i7ToE9P0o9oagjFtBmwNvBCrxxE0DcgS2jebeGtwT54UdnPkKohdnPcanNm
I08IsHCfLfq/on8Ff3ipwXHzNgw8w4YR9DjAEPcCTPKrv5A5+/jB09zKxvNLotRT
8wXl4cyQHCklOO1ZrXbs3Ynp6TNChOnHeJ276eDNdmaj5oMehAGZxoWGE056my/j
j0DFpouT7x4cXd3s/+fZYFyt6QeqvAr3Hge6aYY2mhFU99b3jj7uTh2PhBZhT3ba
L7eIKDXHwGc3NkE714fdbCKWtA5ff1uZERHwm82w+ojNeCgZ3wGqB3cO27S1gxaq
OmTu7MRQjEVTRdZ0oFMGu1E1vxaIjzCLvBf5ff8gJqlsNRaUMWOtV6P/w6fCQFMO
21IlLvrX0h3m0R2ICtdV1K+oVjdSyFdk8SvefszELCObQVTRBTVbrXVW4PG3r+/n
OHYp69HucOm+iSrlSxKsws45CrMFsioAeRK0WxFKj5pxVXcTcFQQfdfRmyQ6kxR1
qMV1xmMt3NDLaY1S7UPzKt7XqhR6BeV826ee7Icj4FqMP1Q7cGlOLHC0BJUPOpO8
2zoJFy0EZn/n5V8KfQbm2JEe7D07asZjAbivrbDhGyfdtN30KDN9bkpHH8rZqmlD
8W0V52Ytp/jxhvyWiQ0L6dH8IxZ+3djXkG3M6Qt3/buqnHdq7I6zyR0/5RtDCaYr
w41quqgEK8+ZI2YSWsoov9XdyDwN+YlFjw8EU9KISwdrzHH9KI3NEqcjeJKB9wHY
v8Z4VKEefsuyCCdS9vxNs4M3fat3wXpJPk7x1B69C+wFXXnXuKvfJhicYxU4wDku
zzsq5sjw2r7wh0KSzoQNn0NOr/VN531OQNb0wPlaceHwk9hPPrZrWhh/nTlnFAk7
/QLfNrOocSCKFODTTatD1b9+h+2/8h6HGdLmtH4Pyw+1c+g61GOscTNhNqjzgEqo
9uvZHfI/1chkZ54KF1+Pijta1KjhhqMwD6tCdfOdDGGelvQYVZW4HjNBbo2Z+GGp
IuLpY1yL6kq2YW+bJ8Ja5+4RRpTwbhL0t8LehzINNQjsaZUlZUe8bsU/MKaTClC6
0Ztg15eYbtMXpLOfrYVEqNnfl8G8r5wxttao18KoDpMU07CL0pl4WJuHWecWWAi/
RhCDCkjBIwNrGQwvtJIO2BwwdljC6yQGYg4Gq5g5eXIFnYbLRQu4lvudT5Ytun4I
XlPo29ys29o+UBmZB5KlXI+IKvVo8D/GTPh14WoaJqToD0XOH42mglM/VToCIMx2
rTkIQ31BwJZE8P1qGlO7PLe1YvShsiAFN+teBDzufYl6VQNocJ0MB4W7YtG+9fAk
+ObjeyUU5LPsKbeDklNxFcVcRFBXmWPavWWEuS3aCu7JtIiqaK4WZosEX0WWoWOM
Kv72iPzFVKl61SzqEk0hyeGcIWGZC/2Bg04xR59mGgxqXS9cfxvbqoXY5SO2cPm1
++pWdUSABqgfJb+7NZUcXVIy8scIedZtTxo1dGjTWZDA5/FI0Uf1aKC3pYjt+Hj8
BH0kXZ9qbuWz+R9Y/WWe0Ug/v08CRrB9stp4VVBPQ00AnVDfhfebNLQiTvRIVGrN
t5+bkQWCDv5S3Y73LydtligT+KJSTuX+kzDBL5ixbq6yasv2BQhJwnYuxK4X3F/H
cj+AxJnEjeAZaNSYTvywaZrwxOqq05M6m2mgkhZP4SUx6lvyMJUi7JoxivxohNF7
kHRWhPzu1S5t7hosQbF4NWj9jRycuFTdrKC1muGck1FoKyV1nvX2tvEcifQhIKbL
`protect END_PROTECTED
