`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDqmG2QZWLJ92q3sW7sX9JUA50lJSMpNIcmi6fg5vN5s0CgeH8sgzYkPBSsuqFPS
n7JgsrfDVNSr2vGTFg7wT/EL8zXE0TPmuG58y5kmqSXhUGOIRrbp8i4NQYnh1GE8
vDM6Ka+Dv9e19yKLJ3oj71AlkOrSChfSIUDogYhRnSlRLSxWELzdo2XxIroQ44SY
1yQDD4DrWzMRQbWcwRoztCmfGEQ/XZFL5uenUuTXjVKZrsubuK36kMzhZG3vIDCv
JknLQIZ7XgNqtTJbTl3mDib5iDVj+tTzfLTzkHC8iEgZ78d5u5OnAHpyHTvI+CRF
VkN7VBqq4X7AYeOhvpKAnLA4/VMFRhvvj6S6clixZt5/u0kLYpSUsJFG+GpN5IPt
wfFXf9dxWsR8No6sWZjVgQnXT7RM0VrLEsFX3c+nijN7L95oEwqpwCx2TdxicFgM
Tamw0um+EF1QX6dDkqpJNxt88Y1nPR/A4SJXmY44JsMGj1YqgSHn8IjZjom1jhs1
+FMrARpNcoRnlXm7uSB6etR7LWKD5bIaO61nTWGDX1aeWeEC/2O9ScW0WvG27PXl
o6/59wZVag76Ji+Mh2cx16F3Zu5c1ztDl1jhGZeUpqELEyC0h+P4koVAjhWKOql5
ZzYX1VQmQGwG2hCJINxsUAQjEJ0OyOgnqTTpMF8eOIHGpzDdNYy+jsPyIO7oEsNe
dd2ta4uTyFnyDcfG9CkDlP+IsmamHE0vSM1YwUZbgPAnhZWdYdnDf3kEzkmJBcVL
8M0FAHX9ztJ+DvggMv5LE1OX0DWet2LCIM6Om1VN2DKNG2QXcom/F+1N0VR/foRh
aazc3+nwz28J4O4fi7N3c+BEmizo/DRwh707lsM32QYd+dxLGZSI4qeO2ycBgOLq
B9w/3s5l3mq6fnA0tbsRd+YiI2wdv9Whg4FOx+Qa92I0rSi02HfDQN4JSXMKTah+
0Ydb+gD2QxH5XSu0XiuHFPwTCfduCjedMeC5Mv/wTs8izpe9/UnHX5f9it/FWz8G
I8O47dWeF/pcizcOF4bq1/EPcaGEU0g+hDdsotJDXeI=
`protect END_PROTECTED
