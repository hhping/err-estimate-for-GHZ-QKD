`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmdbjyDBECDAZfsibBOL0NiZ6RwSDRizhgHge+YMsAtPFAEJQtQvkuqeAr3KGcPo
kGK67Udqhy5oY/eOY6v9umQx4TcsdZ9lEPbbNfcvIFRjq2RUOHcsqdi2WXOzw1mG
OLwzwUFBb5yryf9lpRQOg/Z9YbbVCx618TUyZ3r/5Nx7l9o0v2FrZ7H2Ha0kTXoB
jsj6jCEW9/N4uOx34B/J9lIH3c43ax73M5TzNngCSNZadvQkF5oe9DujcMKvPQbB
Ugk5rzB8SA+8ksCpXQ/+dHrbefrSgwAP69lMTf3zhdadUHjxSyUsJYLwDUCt5Wyg
9ibdou5FZCl26TTHcqoNGPg/NqwJw5UVBozU08qb+rnwVFCilB22meH1uhS2F375
+Vx7K4nwoF3UeQ9hMhszoJevCHK4G92FUBf0JsK+i7Mzskmqx9+J/HXFr8dd9d2f
R+Nd5gmKqXAnrjeiG7SaAzML0D2/j43wtG3T0GdeWbK+CzhsnJvNNQnu94fVsiW2
b0DWPRImkGJBYvBIZN6dHMefRtvARkm/0FsEENIenvhT7SiuYLHFtOGCyvXvJMhd
ucQoDmR3d05H0ljRw+bzIs1/kMHbcrFyppTZMO2xj4gh5sPWxuGlQY+MtD6yv41U
eZCq07FBtv6nbZaFNkERCapiTLzKGjcLTyMdgk6zedmH2q6fTymjz9Ueba927fUi
n64t07orT0PU474ZpQyvN4tPacqUztJujWN/71xgIODMTYVXCt1H/NG1iVC1N+7W
i3zqkiEgXSX6qT7pp45Boa34SKXvqBQ6PN+N7mCzOEq+KbooDSq6pcEtlhHk8EVE
knJQD4mEoQYyxeXvtkb1W/WLUrSfiFEWz+OIQzVka/IppkMXNzgwrGdabFuNfbWE
ZSiysv16ZOd5y9WfjUfzieEm83m7BY9eW7v295tSz5IFXOMszd1sHIeRyLXgt0uo
zn8q9+r2TcByr9vn9zqCapenoC0rZTM+soyITm7LIc7vFJkZq28cHxxkxEaW2fb/
yKLraw1LCLwVFfFEd4zAFa5ey1NNFZbxEYWwpqAJbupZDHRN/lhqRi2vlpNp9Ton
odUhud+MyxziVHuv5stV6tB5UGnwNJJDTzrLQz5Pb+SJ8OvIYPzbb6arr5gZQVVy
jHEUlq7YcobhFQYzCe3zniutkxgG9Yz4uyV+GZmvguBm732yqiBPPZobF/+x9bXD
rhrJFr/Xgd4cz5D9f4biwAMU2gd02HKMplJOJqU2Vl3WBobKlAnQqzaGx2WWz/sY
frl3eEJ89+ZUjcKDxqKOG4i9WwkVG6oYbiRldzMyhlgdPln8tNlqcSrhEe9Tyw3Z
YikTaM0h4VAn9lcnlj12Epi0z/+hqmIQEOcIhQofhDPLq5A1DYmPSVYZi7FPr3wX
g6cyboII5M8Lab2KaG09w4089vQZjLgr992suMX6SsL2xAkT1bIB1cHElju2L4Zo
giV4umH8RibDKK1EZJnJnJoJebr4nC4GxBc8ywIKBNNe0vVf9IsOgcUU3Iyy5LJF
hhJ2WCvOn0CCSHQ75HMFtYTaUZySLV8dp7iIjTTaTMUOCUjvf9yl59nEgkkfRaBU
xWp1C5wkxvz477msrjrECcVrDhZUdPmaWAp6UAdpWoSgQDKDj0X/G4DWSNg4mhNg
DE0yj3SDjihFG+pEIyJZrvAbA0kmdJ/qx0pFbi/i58xN6PUVWlFPnU7hKGd0C5m1
LWh3d4AsfapDPPlesZhitIyi8ORJPP0f7Bb4TbsYXDZH59Ws4FfBLVRVAFaJjEoQ
WgkmWFTSOFIrj/yfzWeq2QDLRRo6Jrn2xewIPLdAIB9+08k5ahCE651kKEfSn8zs
Otr0XAGIyEt9MRBsakFdWgqS24oi6J+3wCucuFMo/FRfKdwL1lW2U0/k1PDVKv4H
gskEfU+WzwyzA7cUxBuyJHjtuXuu5xRYKMMm2JyjiZjd/cQRdw3XBwn04knnimHA
vrnUqpX1q/l6IfsQ6iOJ9SGSKzcz1ev3HoifRtnUGxaeGt9gFhqm1oEj79x5ZCC2
l2mVDYtyL+s5q7u2WRoWg4NK7niMvNGJbi4MmZgdZ8BYynZRtZ2e8Mnrm9aATnQJ
KCRjsfdjGE47A8MsVG85Fq2+LITEHWzQAUXF964Pl9pFn6yMw2sQF/yRQrOuArPW
qTdJ+ZwRz+RXuvJB50yrwFZYxp37cvlvcIeP/X+69tmVadIM9ZgTHp/yvHXNyy7a
OXIDPpi4aOkrSDXCi2dXhllo1QSo4ojRhjS0YanJZRPtCd0UnkGsmLD8f0+Gdvto
PX1BQBwEsYnSWYFK462cPVhCcMRjE6EQofNPRWQk5zCkkben7a2F6DQdB2chtYGy
bHqGSbOrBcGrszIOM3mFIXovCye6HBGTYFYFoDvABXKA6uC7ghEvILv8wVvfqmqq
CG7QQ2bi/rSNuinCj4nENT6SPITt8gLQsqQsODdoltVz5HnKW/a/wlAXtr2SATMS
OdDByMkXByUc2A6To+mZqqsYa3+o14gfvl6EuUxmnjBpl5wZ6QR0lz0+xepneoB9
lFb/MFYrMCDushNP86dm3grHqSZPaXaUp28lCNdOBWxRX4o3LdAyGHrjKKTa8hQD
mmYhvMberlta04DGH7+MGRFq3uKPIvX3NazsR77ZdMQ22bj18WG3cNkCwLJjiOVT
5+4BViragTlBN8/Bz44ldFKASo3pGnBZqBxeKlSm9RtnjxyCn+brd/y9pFye+aGb
KoDbFWCytmIkdlrav7jxE43bN7OCQ+kR1fp6/J1FfYgbqs+41HxrL5toTIt4yFTJ
d3sxUhueCcndltEhENbo2PU2O+hhCzAYs4R9Wm0GMjO6V8tWRmZrfA3yKaJu34LO
joLm2GnTF5kBUoBfF6JXbT3EgR/5Qa9EyYJOe8vYfG5RBwFEtbNfz7pgCO1krSBm
Hm0Fp+EFU+IGudg6kaXfaH0rRcdiPBJ4a+/9lAHrt/4Knl9w1/i5b+CxCBGV0X+7
BV17KT+yB4c13KgWbZIJYIkQfisvlgRntXEIAe1+Nxcul/A9hB6MPCEUyzG6AMog
ZIhedUi3CoryZatrinUoFNI7fMsEhcxD89+qpopXHY2MZCM2DhsJ+UdZbDqZZD5V
H0p2jQqyAuE40QiqjVoW2UqK1FCnscv9Mf+XnHGkkbdTM6S+Clxvn/eJGY+9w1WX
pFFw1y8iHB1yCXWleVzXb8EgiRQDONAJAZ7dJbruwQAEqs4BNQmpqgWIPh0pkHBF
1FK3mCJsV5GVnUufOyvtvZL/AR9bmcfMnn6UokinBeK0ehTRjTSgJlGyYG4FJbWR
7bsAJvZumPCkdCuhQ71nn9YvTAsAVEk78uAp5qCZmDAqR4QY4irniHGpeI0UT1JA
exn2ko8PUdiznscvwhM5I738QzVXri2HI2HRlR4iwpDvba/FzvRtI00RNXOR3pAv
O5h/nt5HbNLLdqLdhqwrhpF+PV8nrPXsJqSDMJlzpMfh+GTRPdL9IJbHUjxUcsUp
hRHKHZ2ajEq0zrrAOcXWVUx2kYYFICF+vsBoRsMWETQ3tRT27rLQYayziQFZ7R0n
u+nVNKd/C98fuIxtC0ZX8/uCZ5xOPckoCS/HIhn22uOGipTD4rWuEKCPDhIXRvTK
TuoFKspEmsJ7Zhrp3zdc5z5nn3YrC5lHEv1dU0x9/CEFZL+g24Y/EbMwXpsVz6RS
RbNbxYDwFinRtIJ8mqgGBAGp4yaBf6mp2cCWnziBxSRzINEBdc06tY0sJdtP5JCf
hOjiQ6CD+tEdXJAYrhAfnpRcN/JF5tFFVk+/6GVfnN6MydtQ5WZi9FwadC0p0Wxy
SzbzLAGloQsvCvRCJzNyQManirLCgOQ7T9KRQH6PiDelk9fvSzpZuZaZOukYAYsx
Isu+ChFQkymELAdBQMu5lLGOkMrMMhfyB/C+SyvbbqnjwEiqWJVh7pksWYjiDUrF
NlELmviZ+GCTKRtWFJof+Gh7wj9J4Uja36gnnQyhN/Nnbkbmo9Qha5YebLLyoexG
MEhYxhMP9iQDzRTORwOgFtVw+udGM+LbNN5oFy8D20p2laq5EUg8MV8ve089+Rym
agEgm0gSgb2jP0f9eb8nR6C1f5z4Qinsmy1ONqvbu2CAyw2oGIw8WuQXsCw9pTg1
Ngd+U0Oh1T8NYsNdXUs3GJbqh5MZG+5I252cGGZG82Gksp/UUA1OzRaJkPKwLzfe
m/Acyn1J/R27of/p6akCmyuzc822TQ6e5nBtz/1ajbucAzaSUAv2bQFHFh1QsaJn
n4KPrzaj1mOojbiXGgjR3Up1T311HX2RXoIfSL97D+EyjHFZAtCbubTt4UwTYcNP
Lv3vv1kp9xAQ3QOtOF2MPJQf/dW6F5S291Lslohf7TWr/WjyPY9qMVSYEnvGFg0X
5LL3QUrNWsmE7zlSam7+bDXnRln7WzELGNMT589m1t6GTOeLR3p3iAwipENslG3F
Ih0vHjnYbKedC0wBoy0M778YucOAjPWRK6qRk/uvPfRPJkiYgaP4RZN9S+AdSN0r
RBObjq1kw7OhxbkSWH4Vv2QqiSUUkJqLPFBXoxObfD7+osIkMLjrFe4jmPP80kwA
I/08g4GzTdVJUpZLO9oy74eQahF2pK9jCey56CxaK6jqe2GQI8ZDk2prnp7H+7nl
UB4k8n3/unmJSyrftKwiEP1uC2H1ToCqCHTUUMDptM3HGpAKhkWrHhJ/GuCKt62b
fZ2o51Jx/+GAgSKG79SgYZICTIGKrv0KC8dydG91ZKtLlJm/YioeWYJ0aE6ICJZI
7+hx71LgibvvfjhMtUi0QBGTnsqSuCx36j3roG6J6yok19H9JZ5YitQp8cOLa1pn
TWm3D/KCraWEUJd+GA2U424G7aJuEI+oKwpW3AMjpc3DTCPclb97qywP/8erBoVP
Uhq55wvi6zUEOvY7Tgnv4s/UMspHBEEkF/guxnhHtcZj0lbBfVrRyn9tpCM+943n
XO23KvHS56/VnNbL9MVb80J5RqIRfiiEoLg0lxM6GBw1RtIkgq7UjfAWGJxXQLYb
827IpcP0Lv/AU0FeTqS11VjIfPiygshZneTP+mbFWz9pZsSiSzWuc+Vv6IMOaMlQ
WPvTgtaZJ37ogEJJw9TUBXU9AUGOEpjKDKkQXFHErNjC8ihida2HxyYncJ7FKXJl
f3bGXxr/MbZMPediyXXWzmqFQzkvAIdvfddEwaIG1eDj8gw9zg2CwsHwadZ5/87R
BM4W5IQTPyh//kB4UT96kCrzPH9YJ8EVkoVxdD8yUO1B5a038x+YClKWJfXhFERw
MRdX1scPSq+2fkcSBlbWdFrK6IXSm0pDlpBdBl/gOrZFrSxpn+cbrBH+RNzoByNy
zPaG6yn2yG0QqSB5G7Utuw4roVOb+XtLr0qq+TnVJOhscBOo2QorXvGYql1Derva
V7D8oTiaMXESZ+tci8gCfhmsNhWjQxWMSB+ezc4Qzm9UiC7/XjNapM5XxV2jEFVN
+lFt6j0e4nFKC2jvHcBlOFxNQ1GmIpPdl+YB4acGsNQTAAffMnf3JZx5EgixRL3l
toIDHBmMDvKrGFUIGb9M5yLlTs4sSed+pgZ5T1EGzBIXm1bGtpV+gYTeUD0Jnqbb
oRaFjiZFVXkU2v9sGCbFYCG+eEvTe0OwiR6vwfwqnT+Kxp27Ut68OoZc32SI+mc3
N3wkq80eokVaYHmRKtjbJM/V8xr6j5eN+bFJQQD3IG0wpkWhpi2YisNpT03LI6ht
A4pQX0Zswd0p+HZJMyLzF1aPWqAN4+n6gqC+GsDC8l65N67N10qqWAZZVGWD0CVo
lb/bkgs6O5Nb6oeZnjkCD6jCV3ltyUbyZydXoHq7e9Fs+/RhhaXA5zFkwpFkSr6E
VdWtSyFK7z8dmuTSxpiSPYKrbdxWsq5UXt7VbhxJUH82a7Ec25rQe/P/s6iePmN1
BanIiLqa9HkQ157MZqNfNKTeMcJHhGLtnr2+2xrlND26XXJSNc2UiPE7FBn9mxLq
qTONTpHE2kW4ZupE/bZ2Si0P/+9jlLi/qKexLuWQETGDlApwyR/54eQpYjrmheMU
LECCrZWvYsM2zcJW3VHW+6G0zTkP/ioZbIZGIJbbOMpjaA/X9bmL+xwFyz4dWW7n
zzwBwbgNpatuQ/b+QavHvQZ3zhflT/mdyQX2drwPFGC6bWF0Xpr7OLdWR55XuOmB
XxBAJhUF16af01o1jTmkqWbS8DCxvQd8yToIktnVp5qPbR+rIKUuSZsUz4xQjQJV
llDBNdGxsnbCixjmqShjd4iX/kl+elpepYb7bpPM1bdxk06Qr1GTK27TAzkcoSC7
u17AYoDR0qT5XoQZkeb1aQeJdYxp7a+jAdZLbN8DaIt8fCOhHjC7IL61zsTSudnb
U/bKKoaz9imGcwAS74QZX54lM/olwCw88Zz6omONPUAtfH5At4h79AQBlFtTLUIO
ZqdLBui7LTExzDLmcvrpg+dG4AGQXMKkV9awVu3ejOXFORKPKYacuS0Uzi34WUHp
MIuDnX+eMFzpZMIVZudJx8TKEHt4q7BqgUZKmcPrI/VVMRNt6BfLZNWiC8DSrD13
G2+m6T1TgnPChTMDKzZldkVfqTv9h9QfQSSijiUzyFgQFP/ZjJMQdOIHJVKNKwKb
8ho+TcSHsk9y4hdI/KFQmv5zrcraKJ3RYGltYPUic/3jBi9nBX55VJfIAHBt62IC
numaOqwGwA01AXF16hg9TipGgCKqXvQ8Qrc7MrjQ3OH1pCJFbrF1zFdZG+i2a2bB
q1fuo5oiRZhS9270+LW0EgcYo7p8Ys/elmdP9qMO5nrjrf2f8OViBlvx2HHx8wuI
ExGA/0R8LnpTk3IFO4GNZ/3FabhzW5NnDDDR/4kbwMyz5mMqJNxBawW6j2u9CvIJ
1nvBg0EbOV7Ed1y/QUkC/eXDf3Cb1AgpZFQwDKcLIisGYKNy3fgJ4pZQfRMVlU1P
QNnM2cAnItJi5/8FPHkqWuSxOMnaKzosgMpfD7Jqoii3EHosQwthM7TGw7Um09ok
b+Jw3Zma2G05+JcVgy/BI0srgwIyA0IQ/2ObNWdv1p41M1hC2IiBtwcUOWikkzOM
xELOARsAI7XkFq/qB2mIv5P3h3z2iAkLBKT/qzjtlGDr1h5St6ZuqmacUAQU8F/N
4trYPUvLmk9j6o33TF0l5HhlykGYVNhzgp/JGZD3JHPWT6Q+4oU23sgL3OBavk3e
dyJTdpcn8BLywObXHalpkElYBUWOhXd4P5YkY5nAlmJ9sRPmHcraGzzdfaS/t9yn
2mZb5TPk61TyyCGTR6UQoe7UcXtscBFAzTNibP4Md9AMU3y+a1HxXGMRpsKeRk27
NhASQUp5JErll7v9zSZ/q7G6OlgExBGUgCUDGumCfUBUU/yCT2Ab8GURU0AcWLlE
LHjQEcZOq5cGNCYxdcdb9U+kgjFPMIxLQGRV59saob19D5x9gi1Ai0GmuVcoQfI2
QCMjP1RjvO+8DH8Z+FzQrKXDC5cEJhMJA3wTjpkECM0wf0d5P+P89n72eIPp3XED
mtwaIXz5dkCcm4SQVQeaxUMnugORVY59UBfhWFOT1P8gUZnUzWhXAnYmAWFJHoO0
PfDBVyRJbiGarafJkXz4RZbCGS6Hagvkwi4PI5nySYFCTrTbl68iKn32dhsZJ3VR
/Ds+o/p86GmRQ4aWnAl6QrQoYx7xa4gJkvYS32b/hGvjo5kRwrxiqEJmEEO6rA85
NqnGXJfqKQJLIOgcwuBL76q2CCVUS4ZtcbRwtr50QgqzCJT4V3kJ494VCXH/kKm8
O9M43agTJp3Y1vnvYikygykT6HjC6PQEUoEK4nTV7ajmreeD4ctAF0q1icdWwUYT
ira/FDvl4S1i190U2fMrItaSTUOESKrrg8cbOHC5AU2kf6brmT1fVi6JsF4+RSmc
vIvidzOHNFOxa8fWqSN7p0RKClWSFAn7MBGupz5WDOS6jucHxjDR+8CLZJnUyens
YEjXb5g5bWgOORDLfz56gZItGIk4wmAc/QthceGqwGVakzntQh3sJhErf07e5bvr
utcvnNW1MS6tZPSRUf52jVLM/DTMy9Y7GUW195x2bjJL+8jQN0HfZfWCTJktHBe8
+rVCJ9nSHkmyQ9F4dnSt5Kj1iPYmRQS38fdygQe+nFsXINNEQkoezwH7mSKtrxu7
bhzw0X/I3KqEB/KXJ30kYyz8dJlQTlinUWb+1YjGLv/LHbVJsieNclzH2QoIZ1K2
U/PHlmH5tSs1a73Xfn6865B7MmcUZkWIpHJw1vl4+5bk20F6kc+/UoC9D3W61Ifp
l7mUZHPm3HvjgYgpJ3QdpUQEGs6rN4R7CQbk55KN2qULT75kJIGgORE1RBz5XXDM
Tb5h0CQyr1Z4BiLhKPWKHkqnsf5uhZINBGy/hYaMWDjVTAtPQngCm+pOD7dOcJ1B
3SWTuruM7UKgEAzugbPLAqjGBNgeJ6ixstIdymrfoJ+wXOTF4SotmUv+w62G1z55
je1+2Owf6vRCJbmCi+y2520vlVtiTeCImvZbELUR99cEGX03IzKnXVIY90NKwoCd
zq8IAfM6Fce/u4/pDvuZ5Mh63PH+FpMWUnZ2+HPn5PMGwPNKHRwobycyiIRPOp1S
bRqqb7z0qhuxq40W047/y3S+rFNY+g0BvU5lV0Q7f6IfCB40uPDCyp9SYg/fL0vQ
Xuajrkdncz4rCDY8khxbpd13IVThLFsF9q4TUWR9w/uOnMlsC8O6qg4PnTvbxkMf
f01460iT62QRxS5nTlcA/59SANouNfEP5yTZ7oHNNebUz1ubrH+7P9wnUQI4tFQ7
i361S1Qvbm3AJxRQIzFdmhEA0NSDpyUMm9Bp8k6BYlM5oIesV6B3SHAISR22gTQV
Jy3W+Nb46we0wNX3bxKBi81a9DgkGYgEede5YWzeuEZNV4y5f3V2rJ75Bg6ipD+S
DZMQwjS4kErQKPeqBi/cW+Vtk15/bV8ZP/rqUcpq8tkT9YFUq02QAzAY/Qpm5gEz
Gax4I1LBe2/bjlTN+rFyhe7cnvQ+NaO56GU4ulnua0roWPgvy+s9nB7tryWUcMKy
TINQOdmEQpcnLnaGrDV/qdVkd/Ncqi7btv/41iUyTaG9ightLQ4554t22ls6NyhK
ong8mUZ/D6UlEk4rZrzIIKznJbP5vlkpAwMKzSfUVrc3MwZhILDFhkSH8umn12so
EAkR2QEj56q8oEunM7eoNu9gNaw/fI+c62fHY4Iw4EKsEom3yCXz4tdLFeum4lk2
CGOMz8LQD/XKrjSRlpTvvLQlCWZWsKT1zTP2aXvLBAPlGE9YSlTlAVHnVPegRSLw
LD5PhtrJf+XXU6jZbbgJLwn+jePs4E4yR7kgnqvY4BmLngcOJ7g155WGBPxOyEMn
NkAgT0ZMFqu5Kxun4D/2PcULFTUnzMaDtW99XLvVIN7n0nKaFB3fr0+EejbQ2atH
Xjo13sdyBdKfzVc7N7AGmIQDKA8efwzcYCDvc/FoGg2HYEvBR8amc4PBwlPTMJIB
chgtrutwd++QgyEOJPpwmNs7OmvPS1shBYGpcOwOS5GRuuks7bdXVu5LI4X4Pf0o
X+rzd2iV4/kk4b3qahrhRoqOLV3epDxGOWXIKJuQkKvHCRfBlOaK5fM+MRTF6wD+
q7AK1Hmm0kTMntgNXekXA9dqrka1LIPwtXz4SQA5PtkA+tVcLccNERP0luvTr8+7
iRIx3DB2KKTV4kj0yOBFHP0lUJkf5ziYayx9HyPFKT61t1Em43hwbUKOSIrCwQ2O
dGoUd8s2EVyaLnJ4Li3zD1maZ9P6YUkzFDOhwl+Kg+XcAYLeIWtPpBsRh/pbfybo
6ltuJGPfLTxY9iI76NZnP4DDxeJH1CT6278Q9/MryMcgENBcE1/ungaR1hIDATMA
00tam8RRIIXcH5JCEaGOCdQNFPDeKPqdF/ybwwE4je+JSKfwXUxg7l7iIkIkb/js
DttnTz71c9HApQA0cUf99pW1wIQUzzjq46e76NQVYwnMeYb9GD4+kfyxZAEDtSxr
RIhlhCPdi0gwGGm7YW/SFxZUdYI6sP5+SwekrSxh0M18xcXqvTUt9L23dK2NnuVP
Qfz+UOH+VtULh9nkb/E0DyhTzmVfSizCrP0hu+zjG4UDTeAQjLijnOzgFuS+x9/e
qjuclOYT8DTHMFTy0u0pH+mOtn8xJ+2dl17LWaeCopS7tHPceTCm6IuQGH4SIqGE
Fbrl7JstnGewBJEUvo15JjBwl1iRQMFsA/syG+doc5DcrjgSnMXtAmHStUlkoGpR
t9ArBVIjYTBqEGfwRQ69nS5go4t8ptGLXz7DuN4urCFdIUw7vuWRgagapcH01dVk
zjZ2o5T3aPiyGDKsgIcDmAyis6t39uYvfwuBebw7Dz47VLcbm1yoc+YdXZ5DFWTL
tfafR7tn980aHjs1VofnykaQbR2GxHABLVaQNoo3vUArGmvfPAqHyrYUIRpA+gR1
5X0Bu72YDCuzoE63KSfhdL0oFZRndpVGA0r2K5EvjrbAjUKRDGE2S6R1Npqcm6iT
GUsxZYoCJ+W9G784CzQ8etNTPHxHLLZGXRFW0nx/4l8Lr/J3uQG7FUeztb1x4KH0
tyYAotyPlf7WYfxbdjo0N4bxgPkDxwSDz+oMjIO5Fq1LEflyL+8J1C5VtkykZCWV
PpmTA9llSFMOh07tclRoMw16lTlItRRHWotDzIIxpBUC2JTxAr/Td4sjiuMUnxO8
TwJTnjxFGlOjvI/HlzKYO0IjYR97Y8/0Ne+c6B3E/bUaLSv6WFMRIq5Xh/359TpI
0of6LBe9Wl2ohcDnPeWAtD6bAQsirlj13jF4GzkYVENqFTPSCLkPtd87IEevOcJq
VxAky4OD7laEFeRd4Yld8s3yfkQxFpzqdzVyeO9pz21UET/Ll6CBlA/5yvSOlAMc
HCUkIUJ4ThwHvRVIni5tw/HzBiNWRLC/0a4uC6DsOA121mQrDKIjJvpv/V5skXcZ
llzNNTRvL1S7pH3Jq6OC5xFcSuJUYAKEqsE4HTEZxsrYnND+5QisL15ISGrW4SBY
DCP1h5YtIpSXBs563CjEw6l4XK5PjBaelmakOuvoDT4tTqkLqgpi2dX2JRF2/f0n
ntz2uuExiK9amPhID49c0t7G8hzKY4mnNs2dT7qQRSmPYTnDUgcwJFDT4aN2ZWZ6
CSIp00xoAGWxidrn41bRcxsJ5riVhd9xBy/qld4aK7KcUDEHHulxVIC5GCjsagjx
WFHLVpco2oqcRC+3whBINgZB7y1tWXR6a6ZUPNJsmjgY4msNraxa5Jr6gNyL6HeP
pNvwO73FDASbOMg7PWotxagB57qD89IA7VUF359bBo+0+ZJx27pOTWtuEi/Uw9SI
8aRt1pK4avy13kZkEsmXt8hnNYMreZrVRjdXfk62nV3gRGPj3lnypxHIqS1QdNHD
Bz1OFzv836Iw3Npk7rGD+Ugcyigt/Q1KEobehyVyH9OZTytYDy+AosbT+iaYbhax
P8hJY3oJpwUcYPPUiADryjTLec4t5xPwIhszD4wL2acrGfKx+mJw9ppz3aQ33fDT
14kKZsA5BSMxsh6luL3M/WWK6DIELQz/DPMGuLp+V/XjRW6KWsj2b4A++H3xLp3v
NsfBHNqkZEX9XZUegqfpuNQjvphw8anXae2QiPbSw5eSCbIAoJWiUnFzKhivBUwF
Rkj2WmKzdlvZws9JY3igfPBdO6FErQCm3+zbPYvn9QiG/TEyIs/Bl2KgpfFXaqUF
unfnnhAyQWgDqIvlGwLbRQkWuqpSViVOkb8/ZX0zswRZYJGz6OMc8L7CsLKfuwmA
9kdTKE8HZRcfmLwpsYln0e9i5OMtkXs+MVyr6SUxun31wMiS4wkEL+RcdeOC/1zU
W34FGmY93G01E9iXccwpyueXx/DMkxnCF4sykETyUW2f/BqHbkKxgROMoTBoKhrg
JhZ1G8uIM0aTJgvG1H/SDBYoK1tcN1/wB+KmG5oZHcOJieSdLsmikmDwQ5pOH+Kh
bAUsKNYl2ZViqjDOqscDG2i1BfWEsO8JBJFfL20ZT1GI/fjA5wBP3fSHUWR4PuwU
3yycn4OxOrYD/iGorCsIRshLDTGWd08bj+kZwXaajlEweajNXkTK8qQ+zMYv/VWu
FzyG/TlelmDOhx+FL9XDbyaM6ZcZziK8ZDyVbd3Qa9hcaXX1iCIbNmovM3QEIyOX
wbGig8awrSOQx92DNrJmmHLwQGDFOSKhHJN54DK3EI4k0zavZDI+Gvi+64I+0JZD
e9xxVzBnn8aK2vc/axxd9rAhiReZ7kkh8WeNZ2/LV42w2SsXlGEJM7jAEF/Hx+n0
J8bJCRr6U9Hoae1iMT3ZJb911lnifn+BMKgvY9KBsAzUlEqR6q/d/iARLVzeiaL+
eFg0PRtKyXi7+IZ32LEwPLx1huA73m54tNX052qJVxepbfju5FKC+ClgeMG1WLAc
RbnDqFcje3hpVdhq3FMOg49oz74bHVU9FGlpraMACwhWmFcukjUrYOqX6yLaFT9t
kBcY2F0sVV9W3kLyFTj5TTa+33gJTPMVJ8Vol4WyAXTWDLbxNPhMvbrbDVdEqGMb
Lkv4oQdDlPB+qpx1cnl6diulgPrXuIuPYEwXZRloQtGVrwmhbA/rpZ38XJq6hTut
x7Tm3N3kUHqd7wbYVxqo2RkcCJsfAu9oEK8yP8k6Cz+lI9tvgQR3lAcFAPH0IaXD
9j+Oo7VZ0c50Az5l/m4zCDH3Fzs2GY+WVLDvL8AeXzrJ8FeqACTACd1r9fAIC+no
K9sdhf3zL7H5yvHMojyZr+FwpE4buwgXxrClzApj2k25sQRY9ck4P8IpMe7kwlVA
XiAQRHnAtk96Z/M8W5UkaIVrFqqtKzdCn/uzs15YZvVH+ZTi7TuOjWESQDAlx4qP
fwu4n6zklst6G90tbp6Hb214/tW5I7LNdoZ3yJSIOAqPcy8mz8s5OQgH4j/I/I42
f75NsWXwQx01w4yLmkyMdWiOq4K5xcFo78L3HOdn/8/M26wRfwS4SlIs1cbV9E+z
MMzN6m7aPpVJy9l+18iRZsS0PctPjTBiaH7kRAeujP5ik2x7C7RDpwLTNbf7Jrxb
tQu4jnbYN694BCWYrXBZOjaQHEY7ExJacrId/3MR/C+4aWfzx4c1orwMNf2A9BW4
W+YsyQi39d76ssTFRP34cXvc0F9l5nPNbHDuS/lM3Weexio9FvXQjGcthKyxmP8O
L4/Hvp55arSr3GpiQhpZW9Y2SM/t+AnFeGKL0DvnomwJHo8xIJpzVTSW/f2As1cV
O5Q7ql/tn9/+Pw59eDysbbK5roDhs0zVlOQU2LHz3ywRWbN1J2i05IUdGvRypVBw
HLLvzFi8JULDfdvrWeMwnf6hO8dUJU1I2atoGIfTz5xtYYRb6pFvtGeJ88jiVXXI
QueK7MgwScaDBno0uTJu1kzlbMCZh/xXDBjL8THAUhqUFtRhCb+da6odyq+AhMY9
pi0ohSpaxdyk27MxGmmMWw/yNgh80OoWJ0xgTh5gb03wBCETwg5pIgTFJRArVN6i
XbJ9TnY8MXS04HWWOnDMSFe9srfJKLR0R0HI+4jqOamXqGtqnKONSEkRvGc+ovDJ
ThA3ma4wDvXzIo4ytYnM7yU+mITp0+Gee1od62jqLxRKg84Sp1ztfTK080XLbuFs
m4deSEXSenbepw3iEgwYK27UAZdosVNHEK/KHU4bZ+ZP1PhIFtTgEDqu7sgS/w6B
c1SVn7MqaUvqvlcaTz4N+jOz52yPH03Db8XL2bs5mkVecBay+lWpMZ49pxS03vaj
XTORUsn8h42udKN4yT1ZT7FEkiVQFznIBfwV553EQoF80cBUPkUUvxlx96qAaS1Y
p1iF3nSbowrs/wR56dEpbJNx70o0qvIpf1b6Jw68g4YM+8AOFq3CXDES0Cemd+RK
U/VtPHHSUKazcyD68qU2gBjcbVBQpLVLuH11TrEYuD+ctbCbswkZrIAqGP54ESVG
TkukFT1tR8VAyrhvB7x0jCitM1/keRaYa7/+5xEy9WnJCl8MDKAbabhFPbaAuQwe
oKbxx3N6MDv8VnJGAJ6prQ==
`protect END_PROTECTED
