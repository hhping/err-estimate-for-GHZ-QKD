`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0axHe9d5Dsv8yJbKxJ/Ths/unInPicANRaL+WENO5VIJ91e1TP101GcSRFLRAIit
LOa7IhQInNyHXkWMePu8DgRX8XfbIEQUrlWUaxnZMcZBerJzC1T8eB2v48p8BaHF
gTpKxgIRn7H0zN+37nvw+hNcsXpJxPYkakrUAo8YI/woWV4VG0wHiETalFr9rFfr
kkIY37jIVNMup9hFWukTE5R0S/b+VYG4651c+oIbpZbFug6ULiGXBBvUWqxiN5ce
w9phdZa0HdkbJwSHNtzT0kBzCq+wx5OmezRSVBLKsipvNUKpFWQbQgYE58/BdP1s
hOtAzLcgG3v0yIF7aAwsCAaE1egWC0Ma/khqX6agV89LhYDwionvU0ZFLhQT89v4
dpJ4quhHRCRtWLTezLHnFEs39om/7YfjOS1RJgYpQP8Lre55A3l5DD0V8HKnw0jt
o0DegCZe0bR+us9o0FLH2lJp694vk8kxzxWYFDY5mSbExJ6MGbDyJUb/iZ5umCrR
YICnaX3Tgdip+pPGkI10rAWKouw7H2kU4/GpLIdA6zvlLi9I0FeAKJKbTCJ82qpd
cIxJ3M1fmcscG6dmUsqvD3GpIE6M+mE43UT9MLCquO5qx5TBE7bsR4XOgrkRazud
5M9gpsYxOHLsF2HyYPynWGx1hufMgJ2W3nDwa5JGzOuxlohvhPTSMdPPrp3rrdPr
VvdJ6WXK2xRF79nySHaYzrV9+oPGKTYkvVlAD2PMa8J4SGEZ1Ft6o6v9kL6eFvlM
5emPzqfX8tK7Y0tYJ+g0+gQbwEbwUUC5NF97VYq8oUlmARHuveqFVu/2n7kAgdxC
uu+YLiravDUZIE3SGeXohNEI1m0Fm6MVSpTuYUm4uYYd4FodqHdSYOcTR2/zAoQ4
Wd+O1QYBqNNulsj7qw2jpOIrvMgvoVzJ9oGxVHTL6V8t1B9fCTB8uU9XM/u5SJDX
EwCRVlF0uXJYcZbIQ/1MJ/lyTn5IUoyrlLXawXvMNe9TGKunQWbrtk2ouOq5NYxr
8uqhkkdBeqMBxcGIDC4rkeD/1nFbmuLqTKVI5uxz/VYAK1o1Nfzks2pd7uNIVGCn
eLKTnmF4DQdCe9gAYeadXwN9mdrISCpHiCCPKiuRlVKtZCCrnBzo4QO0JZ9hOr+b
1X6ZR9wcOeTrOO3oN0Vd7Z9i40WRuuXxjSi2NnxaEuBB/SoBNhL9779ROswty4ej
rhUAHMXqvj9r+7gpnSYH0SMl6OvfJE7o9mzsQwUkLKHPtyykrltJMMFYnSepz4Xi
gUko0lrB5iV3YavJptA66N1Y4RbAei4yU4NKwhZ4EI/KB7Ff/ZYAFGBe2kZdcrH4
AnMk3Eyq53GTvLj7hSAexMjdtG9iHGwnCMiIaTslM0d07rWZC1QKpW8+XF6sMZJW
mC1eiOyr3xw5QsjEggQg12E32s5eS764ll8QUeuIyM+qiZ/ypuj77bzASoTifThB
Y5QySPIG09cMgNrx4PzWejdqYqbwF9pNLvbsgrxR0AITQf+AFQ6R9YKwXRLdc9vC
yKox+eZm7eMUYhf2HTDoP2m5IrWtBMAF40sWXdW3R+Q=
`protect END_PROTECTED
