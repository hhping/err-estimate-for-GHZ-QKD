`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C03IT8Rz4Sg+i5gjN1TMBJ0TCmTPc6S6zB4GVargXUN9nvEHKF3+08A5VP5pIvDe
7nAHaK5FXVqESYTppgCT35/02pEGZDtWPk4iRge4rfaPEz3RKNmpOxHYFTzSPQW3
/383sFTmBj3f87VqpD/2gu8DIvJ9FPV6HI/TS0L5dDujIYy7zO3ppQXqY0D80aA1
pGvfc7U9QHgpwQoOJYGfr9nWLr69goaqFeN2PU0dTs0bO2RCMaYJZwN2bPhV8eNw
ZxIlvnzz5zXeZTSOkhNsQtV+AkT66/E+amqARLyf/cukk4/ZIoCuHgA93hrNOGdS
vMLDvizhei3MMSJAkCsBNtkyjQ+xQYE/EPUi238XIiHfeYDwflVL3b4+hxPk9zNS
gp7aLeGDe7pD4xGm+JufdF18aqDAFucrcS+fQg0x+RvOwiG/m9zhuLfkiWmD1AF6
cRG0DtsAQwcDlGPlsHppsakJaQ8XBZWz2u9EpnYrO0iNF0tHLQO9p7m+zcIEdu+O
dM9CpRCYsad5emgD7+PKTQ/u3vl4UyMauJcTp15M71W1JoMe36YBpIk1DgY2r2gP
JydwOJlhyd5cQu2JxgbeXHeN6pATd8luWsZOy6FpiNesAEdl8VIk4A8e0aJjZ/Ad
TnDJHzoKYgw3+tm3lXRcobvc21XjcB5gcF2cGkfDOkSlB6eEN0n5vbNIf/QUk+oO
mXlcKnHCeqHcbxY/5Ihu3G8I/NkR8qmdaF/YYuIO4LFL//v9WIRAIOj5KaAMGJYG
ZoNElqbzCBJN5osJwLSUQpBoU0O9V62aGJGusRjeF5bFxoX+vY/GumjRSy3EhD4V
pTKDZ/Gg8cp0kYd9dBywlcCU8fX/fUEolcmlLRABCQ2pn/uAAn210k0C0LnviMCY
`protect END_PROTECTED
