`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fLwiuFFiPhyK0/S8g2cIvoZSRcfELrOie+SyU1BX7RmJ140vJOGnc7xee4XFK/k
4w5IXpsHPLzRK7EikGX+LtmOzj/HmKKdYfqU3a7J3Uk4y8wNCic5mUXxmND+uUbC
AoPSK0nMjqUK0mrypQ3ZgsHaNR3Y/WHiKdmiKzNfGB4L0brpwEsQ3K3VlFRZsxFg
XviY/MMRL92PYmTMSVKKC9fNqiEhOeCCEIYFkOqtZOs28pajHN6PQzks9v/iM9dU
xqpZVe0OIcBW+MkKFFMigclgaI6fsDH2q18fuAIwGvENb6/RpTAT7vF5bf6JBx1a
Kzf8CBk8oQ/9NFv/NeLqtufRGBFVyJSLXhc8mp5hEB0sE6+CsBBFkdpjs/93ekMt
0YX9lkUXVdMjDgr+RJ+X2FlYFYdZjRVXaBaojAGH62BVtKGWDxoLN5LqQEeqCRZo
cRiXTMB8vSxQ8PfXy5ZIfzf8+zT6132RT+eV4tiRCXvqURsTdHUedDYNeyJCYPef
mRF+lWIFNIdkR02FaaCp4C8yIzs2/ihHIznkwinoi1BY7nJBbI8qhzU4rfg4qmaw
awgBLkAujRSHTv3Tbqjd4iFWn746fFnYX6Tjvsu2xm3OhDyS0pZIB4PXfH5RVoMv
446R1/r0djgLqhUA8LP6nxPKQdcWRe+JJHFJLu8CCNmxJVXYTmd4MMTR0as0j1+V
zdVEQAnPiTiiv0nRHiONO8Vw79X6wMKW1xY+oK9z6Owpb6T5G644toPliEan2epO
zRMLbbVC4Ikdr+lx3YqiZL4466D7H/ZkSPWsyCmOFLixrWCzGOdgRSR7JgcIerbM
dA0sWDy+7vpNDn+bau67rBRD6w9wdOEHEO6XRRz8VzIbMJzw2hsro0IqPcwgbT6o
E3ILk9+YfpJaCVh6iSzPZx1rcw98nia/0zVojqBmFldnDHFqL7UCEcEYiLiSdWYM
umUNxObh62z4nVFu8cfqcRD17G//D8QU40ylImHf7fOYEiNMVELd4T5gwfMr0sie
L2G/Di8qFTIPQgeJc+2pdtsQgL0DQ9YdbweQhu72ybrzkA0q0E/V0vW+PeHsPLw9
7eh/gRaccfWdZ0WRmbgTHDcq1JJOcW2CSng0gXtx5ZVPNl59RxCylxyQ5ViuxVU0
U7M9Q7f1Yi4c6nOsnhByb5J8ioTT1v30Gnw1lNGS7hPEM8vbOAUYX4Kau7J9tJlX
UjyaciqDFU1sksq+xdVnKxnQEkt6Ert9tKIHH1WkTrzZl3HCTnf0s7IHor3EtL9k
OoQZAZfljdNMxToMxPvi6f2UlfVA5UOCxZKy5a+aLi3uf+DlYuXj4s7LLKWPIw8z
ZwoL9EXWSC8Wf5nw6XDm+Sfmkmbgg9MFwosztDs8qtLBDYuQ4zscZo1uxX34GoGM
yNgauSwrfO8zzQHws3ilTEOQEPl/jGBStetrTC7bzqj18vvdLnaLWk/3nBZf9J5V
zr4Eh4k1RhRX7SczfPIBGcqpXJ7yKXt1PFUtkR6rU8QKDg/5cbCkFxTR1x/U/uOW
BhMWYvkDo0fo/gmU2BOFpP10a0eCVjqUIkk9WDVW2nGvnW+MS6K68DsXcVo/Cj+R
v929ZLc5Yn7vCPW7yGE26W98QirwpITO+fKs4fYHLubpSYEFXtNDsotMsNYs3HtZ
9HtyuOOP5hfTbPSKloq46AgZ+QyVvunO4AN9OfEEZ+8tOiD3tC6nl03C1sLKMGC0
r5yagjdaR+ERP3Xd86Mt8EhoYOIZAsQ39B0suVOs/Tw7QntygHkEwPewyk0yjis9
XAedHlIy8id7qfFf+m5gVCJBAridyRvaW1WubMLae2UE/oL4aCXSm6v0DMci/9A1
A3JsIEVmpl5/aH9yRaplMPCTl6U7Bv1DdUpAG9Yp2rFcLRvtH3bQwUXBuKAlzTa8
962hPXUERu0uael2ZS4C2/rD15WrsBD/983PlQxPsmZVg+w0f3SgZrQKeKKyVShR
r/4lRX/yFg6v8VUTlmFUwTgeQ5aDeRNsfHzx6gYJhJUpw39whLGqukMEAOj9JdZM
QsABvSWyNIwx/kfeCaPye7c8r0iXTbQBsmahqOI8R86RYkIZV3AlD9jzjLLkO0Hn
4OhBLAhLYE8S6UpYVCcZWYfr/TwIOoaS8U/mDeYDVCIg7vinuJjID6qCXkghk7e+
WVHOLnu4QspThKXRypCrTmudT4ioUFAykZu+hYSWf9InLcfvCIPfzRhgc2LftU+A
UNlhs6tISxW/bU6NeLR3FvF1jZdf4XwcI5mNliYq46fs7eQl1Z7AgTslS/dLGwmB
aGD5zu1jnZZ0bnZh25+I7d5FFBiXSFWa7/YEVLHOH9WJ0tm1qfclTFDA8k/aDkNn
L7iMxrpRSn8zntrcC6frQaPq3yAw6Xx07dok63wK50urXUUI/1ndB7roAaV7QiaX
6vSwNZViUlvg6B5RP1sOmF/UG0SDwdyuW/A+UQZx6NC3uMReQauTzloUU7FLnflg
TUHrZmd15do/u/3TUQxrYPdwZ4NtDEy4DPIxAErByG9sv0xlirk9e1eW2jJkstuv
Ui4zcF+Wd8TvACpyV9+V6PKaBpcKb8AqsB+lJdLiVSiBveUZRB+jdkXC0Ch0VkVD
kgqsREp+QqMxjq9QmIXzywa7F7Mccvsn/Ws/cl18MUxwPScdQYD0sJ3oIENZxbFd
9Zxzpcxep6JnwwtbduuhQPvJItbEH/XYFoNmFqz3H2alLCYoUHbZ4d3f5/1nA90F
DoL+Q5QVn6A3PSsVFdr9fSa2FyoNowFX8+8kLbQLtPya4qQM1hR0/uiWel5vVjb6
j+RV1KFOxH750b5gvsppe0TLI6N2PqMLYo3xLdOUspnCzSjHJGWnD7KPiYGkT49g
NuVaRMVg/0+7E3K+sh7K/qFm1ZZzSZnbtY8UopxBZwvpMxL5LO2PnIGSCZwHUtxA
xw9DoVOjXJ1NFAIFqwnwotXUyvlJTreNTxepHbtIQbi0i1IWlEbSFuOl5US1Zw7V
0B+zWU6Ok+3KYjaXWopM1NkDTvclRWfSYWBi0tWvaPcZkzM42P91sz4O+br1dQt/
a68IX+EXngkCDYyhQa2eBwuRTEodnZ3i3xqf2BoSB8k5rI7izVQriwlqoURaw0Om
oe3eEBPudooiovtCV3pEbzSdHFteOGg3ZBQlFgF1QDAmiIkUAvlftXlLrhPWrBB6
hATMJwXKYHpMNxjmzF//neO8+JxHPlvBjJfsZfbOhIgyVcq5P1OmFCBwEcoQ/GZB
JjALt8pI9S0Vk7iReUDJn8TNv8PUTdyOQmT1Ouzf/Q9OOzTfVHZq3cJFJ1LmKcvw
4VfZeD6b0i6nGUipUvQaT8eLY9K6zkLdW0M9E24izQq5WuROandsPbZCVOuJyE8H
ig8uZUd37eTy/khjnj6AJQmfel0NGs6Ny5ZXOioGG8ZpvxEG3csIKr9oRvUkmZD0
lOyBPrhFrbdVhj1N4VnjRWPBJD4iiPT1XYgQLZNAATPXf9udh1fC0+edU+U4wqLA
MoLjQCW8P/dRKAMngaeFdm7yzYkMM8+BO2pMvoajHwPZBAxnevDlQm3zXTHjJjh+
gTgG0t2R4FinHXuaCKAII5ac+a3E9ttzdnvaAwqfBnah9xpwI9rW3O2JhE7hHEYu
B5lN/W2cvC8ret6i/7+o/hinEJLWMztu/EW+rs4oxE+YRolL+Prd03RkFPB3EyFx
xrVkmHEg3qMdoWIwa61pSTrFUY48kLZuNL8SPSzrckNrgRXswF+eAmHNIICNfSxT
IzMMSgjz0USCuDU7HQWhcLmq4I0RGgyM/MYxLqTDg4HliRr3fNZmGfeiQeIyK+D4
1W6sOKvkoBzorw6ndA/ltOdG6xKf9FfPu2lFPi4zT9zggeWgP4wsLfml4wJVQ25Y
jPOO1Qw51KKt/F2DlrtBxYRiOeZgoqsB6PA2E9oex2xE0qCJbAT1lUKiG2N/nNUD
7bJ3SGYq7/+uhVaaH9vB1bsmpHHLkdl0+RiKhdb84SeE0d8ESetp20gIDPuvWHCH
fuqEQ8dHvkkWNq4s4MQSexXb2TWLfdenuq9IliAlWd0xg9uxmDq1uLcB8vZiA/hn
hdbwcXGD2yX6K26JKMt90nFVbVcWL4Aw0+rnN7AC9abR5vaVNiMgvqCcdjTyyoxR
IclARjRXAOHfsnrX8GLvQClShvTD9qyFdENrOFz/CN5FtTzRDXruRel6nOjUUatu
sJAWyz970rpWNCtRNXJZnXIJHvNqfsfngcZt/UZwkSvwb5RkQhXRka8YcdrKiW1/
PeixeEBzunhtv3gBi4DeEEXZN1XucbdXuzT5NvJLXAVX2LM/leUkQ853K1dne3XZ
ACCAXG5vRQrvq0lzoOqopRPnuL3gd8zwFycXyn+Je3Hyn3+Ts9Rw2MGuJPRfXUhI
yU+OOkvYpKgbUxhIjztDaTWykW+/OTbZAJIqBoR7mMfj+yhY3inytyCDgFED4Itk
ELdTfudpGUBiDHCh217R2W0ikvVZtCAaLTEGjGyXu9bVMVXR90RbCoZkxhEiiIgw
S9OQVi66jChHXDWgAin/zwHBKxjQaba4BUMFVuAf3tpVAa3aLWnKCX5qnsQJAWvn
/b6SjrDSXKVLkull+9qrQUhjf6JyjYb8O0gXwE8z2+aoUXx0aP7jScJHsWvBE4aP
9cwerlPq5D8hBMEQfuOx/amP/3HM2nmuvI5IxJe+tmrrZTPIiwtU1L9Ry0zrEgoT
QMLA8f812ajOAw8rFu/NuSM5QRGdqJHkd6uFQ9GEyGOr5hEFR9lSzqZ7nEAvUhlR
8vWZWqKFNWxF//x2oAsgbtpPy5pT30gMHXwvuBmXkgeN8+08rYPurn34Ju/8r75r
UwWgxJp+2veX/A879svk92VkBt6KzQG2yegE0GQ0JPWXqQT1m0PjcCNbYGzOnwFG
H5rp3FDcmmDkJfWGJn02bBp5VzDm58gWdEaoVqT6mLTEh7CW9O71PuQx9W8B0+ES
ePqzQm7Vht0zvImnVA5vW/cQzuGtzkZPhnHllAu//AbjMs3270L8RhkUq8idYsD5
t9LFPAu4lrU2fqO0bRS9qJDUhaJS75YdaZCOUBjkR4TqfvQ1dUH5hvl48uBq2foo
KrPm4beC3Z3CnMlTLM7dj0tyu0roW+mpOSXRuXWie8L4QJQxQ0sdXeR05+L1QGUC
WjxESufwmw1Mq4H9z0tNfdW3kSyEE4427PVdSiCQ1W1BmcmCBHnePKduuqcaDuHk
8YVgYpuF71MhltVZ+oWZV395mDFBDngqYGTwvq3pkjVIAyhDaJVqhOf6cX4KwFG/
aGPUtOdKSW378iBMPcfR6WJk8l1PMlWgodsIkcglKKUTc2b4ROTQuVFnur8fh/RL
fJamrzPt3JAiIZv075L8D1DQ8KbnB3Os7kBqWsjE27FgxO2ozQReoMSE2AYrAkD7
Kn6e4N8QUSzG41UzgBICYE/PGXhdiSbX/c6vWSkb7tItQQn9wfXmGbfbySwtiJzu
8g4+8ADyF7/IgQF8t+uFcbdRPoAe8bhB+sOT3cZCiGEmnA8r0DbsI1UmpJvXCIWh
VcYpzt5E+Cz0ZM7HLzPJUMkAM2czB2aAVTJzF180oUSVQQeYmoH2VdY7VaonUFG5
j6/YYMPKNQSkrXEEoFVznp/4J9e5fHvaxOzuyPlIbTKEQd9mxHDyN1pSidL1BA7Z
C/c95Fsc2dIDdjnDRnp+l/pplSz2bnc0dsZyzDydCRTRbtxLHiOtKLnCjhY2K8GL
pNrVUHCrQqSPti+HHEyz0qCmqKVgn7AOWUKPbW3BEZ3oY7NpM8npvA8Ye4guLcJi
I7Ev9KlmhRqRFOaCsO0Y7I90tEOrTm5xCqMu0d5cZblkK+dxGZ6+xl7ZVqdAmzE4
Ma3d6Bhfwxp7B8005igrRfswS7RMkk13bpfC79wDJe/XEb/eRjP0WOmBWIIUBTcl
4psAzG+GYLWNfbghtC4Fnb0VvQGjj1G1k5M0FhVPHXYH92FKBtcKio4yVTKLBYM2
nj5Y+e9KlYhGktzxY/BfZ3QMWPAqV/9abfaUmd9YLoakPebJ3/K+GzKhJfKqDcM9
xQVhL0mOS2yTM3TzXrBacq0zqn481KqFJmeHWTs3yMrPi/sSl+WAnZoDWVGP4qp+
YNp6hvTSDC0+OfGIeVipEcBiBf+t3rZFhYz96JlYKTHmG8YYh3nFMMI6SOQKcLzo
VCjivnmIvB+yhW1LXhTkXyJgPTxhsGcuaaKlG0A/b7B4wktHdc/+tCshqRNT3hwv
nT1XLje7SOV+j9gDYrJgmrnQYWfoBqecmWDo2VDmV5l9x2mhjqZvJmFv7cJQdQCj
GHnRR4D5SFNb/3u+SbXOOTyVTSNVANAUKDV81toRTEC9f+Mjlq1b0NYlw1Zfl3KX
sIo3v5HHjUEoxEc+P6tXAzN9kADAa3XuFIbIXGPmEfcDTJq78VEzEUdc9wQOB6br
nu9sE/P36epAXMTrQ5elEMKP6lumN9MuDR6fjnDMNDZTLaG5hhmu+3AP86Da/gTI
Fiy7pjSYYvmDG5Hy4ln+siTBsjaCaDmVcHK5rm8CwLeEcquDOeYdiInpDO9tlOqq
pSMHjfb4Vy+QNzUWEljJwiOCqr+NJB4wHZwyvU5SnvX7bWi7Jfc2kSwZNn5X6oeE
XXky2euU9ekKDdjq49b3TKQuWxI7Ziu9UIRq6tCK6w3r8yAUhiulSjId6NyanT/r
7YMPobD0X/+Z16kOEIZEgLttuaL+oWxKpd9wv44pOa5vtOhOjrIYCPTfekZWXZ2A
/Nx3gNyb6k0pN5WLfqevftESrKbcwUhb2jvp6rwndEfVHKPeRelk2yw33MV8J/pu
L/qTB9ZfNYmPbZQUaeEZA3qn97u0zjhC+ZX146G+gJfIyMRDVivoOR84hVeK1E3B
HtI+vgDKQ5WVcFE/mjNUY93TUnIyCldzlxXYVt/G4uc6bXhsofQtPXns/fn+43EI
+2NAwe0DglnqaDZ8SGwAv8iXM77Wj+Xu/CqWcYwTM+Y9t84uTTFYEnNgpxvIUwSh
6c+bmYNKDRmK94JC3pevYD33SQqBnqXJD/7aACTm1iK049CbNbuZm/RuZXSH2S63
Ws9oAhlyHgDtDl/ove0dLTNF2yTEt/LPNFITWek50phejFmhYY5+CH0CZRlhUf1U
EKiMCFs7EngO6Ro3bNJBOiIMkWgdVvZ/BMzl20iSftOSdk40yklWfeXbp1DAM+ag
L2CbrugWb2Vqtsi+LTOzPTRYuQ+roz7A987YdRVoUg79kjbnrZWro218BAy2LyDZ
jQG5wv2d4iLpZEf/eGz70GBympVYciIZL7+pkJNIaIvA1rIWOGmtXJB+7Iw4imBM
wS21nqxXghi5dWS63g96F5kjklRUGjNB3exCqqArTIEn+OH8N68qJU3jr0ue0MZv
n2TNPjdG6Ohj1VCaVvCEJaoDjtRp/bPO9jb6GLTiOKj1S7b0fmXpnQKp31pJjZpR
KNTzFZsI62/eq3uiLCBzZntIJYql42Q9Un8m5xkvdFu75iAWKumGmqMALWQUC24K
zf9cvQJsU2zAvl9OkLIj8yeXoS2gUCkd0vTKLgveVbs48DI2AM1Z0iQRee3dmf0E
TzNLvg9psVomGhc/i7KNzk2OCtanuxT5sBq8dDhUyNB1PXWyiqwo4QnmODKIVvgY
u1cxdN0Pi6r81PLRl6Ns4IsmOppzF+ZtqpoDta/BKDoCuRO3DKJD02JgFLh/JM0B
1/K4+CL5Bo8+1NDiQNvoaMqCQz54XOMkmoAeD9HoikVn/74XjYB4JjCFSfilxv14
jWsgkL9QmBp8xgKr+Jsz+SGjRRZDnSjHKQSys43S9Qr54o7vig5EYQnxILrrjDaq
rTS9/09YdLqVHJTQCfSyQNqz1x/h2awoDwZcLcerjCgXOD3iqoe9Sxhtrr4lsAop
/Q7DJ9qKKSMLoB0ciZSM9s6cVTS/QjYkE3CG82OzN/a70GlnYHkW+lbqRBCPcsWw
kY//W9wGHN3GzJLt/lvtTkoW0bztvE1Ws9DktTD9Yrjcv4HA+/yhFH6InlBtuIjW
EwMn6j7mpNqmukQFPrMWPt9s/jVuG9w4QKPjKJ8ivjApa6Tm6eVKcJ5vZmgd5ZGK
UucWLGDxZ5Hvu0RXUTkdodj8/t80SGl3jDtNSXKYjznSJrNmWk/JHjmqNiSRoo5k
hHjADvaXEJIc4GjdwakEZpqWfgsh6G6PhXhvY8eSMnQ9IJLqMfK3mQn2AwmeNd+G
mZhqRVdLWxf7eKlBitY8OALu7zCXYMdLF3HJ/qBEjEqf+wavRZVysHy5A6mSe7S9
8JYugRBSiy83Ca98Csxijnbrw90jTWrOsiENqwitBrhPTiClgYVtWWaa56c1M41t
FateTWIKMEKBa+3tjW9U8fU1rmJG9ftFfZY+JQNY1WaD3ThKLbQ1/5YzGNYV8D/j
6hdoAKvWZpwG/fHSlkLfrAZXFhUm/qZTPiTueD6rdqsUQeTimdLBc7BlurYAD4t/
Jb0BkMOjuv8v0T+dULMTX7dmP/OUavIb0j5F3lpCm41zK1oshLkB3KKXsxQ/Jszc
jMrQn1tJYfsSCmxjvUuue67YxPySYIzekGztTj87GMSZ7ffWgEDf+WDjqidp7HTX
la8h8hw3qisYXUjYglj2yGILBXVxim7CfGMI4TPVrTLVds9Vgy30K7DbmnPE9e1K
foStqa5v1UpRvnQd9FPT4Pk6Mb/q3vwTWn79pogiBUZOHVnlbxgyCwJVfiZa3c8Z
SUBH37lbutcsAic0Vryupn6HqyGQThaNeAqPE+DLYKMAvJhBHDD4LpbEgxShwd9g
BRQE9SMLnHaOl0UJrTdJCFMTNaAuJ7NkJn2IHvwBnEheo5OkFFOvjUcgV/dJNsfC
Dr3nnq6x/ST4clxrg1j3l4zoBJB+/GwIHeCLwJQ83U0Fr8z1Q8mdqJebLkCC1YFd
StNRd/bsxlqh+DWK+qauc6VvLiS/zwCryHfAlQEpymaTZUyedLwDvIV8Sb7GfeMG
sgiznvtgLwx/eih/YwuZMgiCwxnd0wA6rJIwMTAAP/bOfRttkqeSaXsB2+V3alC5
DYDFgxWjmJ7e4goeUvdVQdmQfkp9T2FWjFqYSeUuSL/H22RC8dtDbbV25rMK1RUD
LVKumrAxlBkP8IoBR0Rxdg==
`protect END_PROTECTED
