`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMH6plUwI89TmOLVrjIKWeOPfPUjxe4hVbIzQTLzNq/U+1bCQuXziu/adUmpULLK
m09Fv5L9WvRmOnSWtsuf5Y87K9oxdJ7RHmtJ8fFQtmA8TGlrrvcISGSyCaFH1oO7
m0LGBfvEfvtUxmE4aZe47OJK/N55Etbsc34+sAkTXpv+M1QtbzcL5r8dxUMb12hH
gwIxMflgGm/m3fNwFtaJtKC67L7OdWKj9XxXd7xfB156EKXztph4IA9i3lbAztA7
tB1lJRgWN68VHG24CWEflOHmuiAvRGevEpBqI8GcKJSfCB/iLJHtDPEd0USvwlgz
y2x37oVfBSUQ+sTscnZdehTos5J60pFstGGMkZEK844gMkF8iU0kJRRYWaatplpE
Ep85WWyYPffv78R6t89hY4cqgMyp3TFEU3/EpnrFa4R2bVRHGDpW6n1onQgDRlTT
UKbBtWPKtUoyS8p+BRpqtyZxsSQ+1jn5KA6Nh4tNPrmICHO1MQK5dkb0cY0wsxoG
XzWvmZQOUCG04hY3qBELC0Ep7JgDcmdzJthKnA5wSGO+bGYZUcbPjewVuCiaZZhQ
uVrwEQ04RHdkT2JsWhFubC9W+NxjMZtQ3unu82U0XgdR7uKkFMFSAaeAr7j4fDun
SlBQYGeVHQ8l9ThzXLhEgHKBV6k4LxpoHLADLN/V1GSLYGR2NzYOY5VFE22TRDmO
r2QQ/6IkR7GZgZrBC5Qkil8sT5y8uWEAT/91tdmPb1TQa/bS5FsSJxzChsZh3z4T
u+RFvgyRuHI+JLBJtKtpQtALsX++tgatslbrrfnX9ynx7tr4Dbha5rrgy8IheGRL
OkVzAgjY1xTxzeM8W/tWFX9278MjeoVNtjIz1kD9o9IDR5qwbADkHCaXZcr0IFcO
yibiowGioiWctKfFpTRySMWLAOYvj2wclcM7m9rkKvXAJD7TO7MO5tXuy49eTEvE
Whf/9gos2aIJ7Emf/clan8uNugZz4V7rnCze92pEMIMu+Xoq09I0PGlcufGIj5aF
3Ra27mehhDV8R8miIdgrN+/z06n5jUn3sWo1KKBqtxkrw6T9TSlhFhGGwCRBbJvc
fpKc7VjPEzUNF5udp0+vTflWFK6MyG07DYq+rLA0nLIkAmr0Mt8UPBhbG+LiGcqt
ggLojwDt4ifa/4VE0pvFOYAMz6a7VctJ+wb+3IiMvaBxvrghP9hIm0OBbGB/vumc
8Cz8r7wPHB0ybhqoxCTO9ST42Ywk/iNwsqOLYtzF+C0cEcgcUaKDFZP/i5L0jHqT
SsNPWcXrHRBvoKaNOGBO/gcYMx+SkgyhDEfsDpocySiP3KxCDXKfx2FeHe5oKL5w
7ynyQIYG5+LEy/NfKcgi4EZx1BgMc4dmC4fMCVd87eBPMn90fT2X5J4FhlFLGYXB
WJqxocqgA48tpRv7+2BJWWcQ5XOne1VIQD6Mk4/ZqgstgilxPvo8IN5fLkSA7Imh
Iexz9uUdA5YSSvKd58jz2lhsQbQ/zZmLll6nsK+mBUDnnr3D3gKiKgIlL2l92zzz
4AnkwT9bmm2A3qG7ooRkAxw1nz9DARQsye9RAdkSkxioaJHa72dSvKlZUAfRyABW
SYnhJlYWgaPTcYJOXe3f6YkMQVPhfediwF7XgaI6MfmEkeA3wwFqsbx+3xhutRn7
XmPeZ+QWuPgt5BoIdlg+SUn1ZKsHuBRVdXTjN9ZeYqkNkNIZScafcJfmVHW6/On6
CzpKSBEqcRQstx0drs5AMRWCqa54N28ulk2t6yipdBRP/k4xmYWskvpyiw4tv7LM
6tPaYg61FAPYjzCYSBVTsfu2iClYtenrGTMDQvIr0uUX96WMK4/LsVTzs5iXK70b
VUUaYOio7sI8ozmAvUeMas33Ulp2BA2hAQbkRnA/M0FV06lP8NhuXo+a25oaZTk8
aboudeFMbTBnia/16DkJqqO3DClalOsdMBJrORwhZZmCMU6yGIfkFYCpwnSjOMbG
UZmn9iQEcB+hYvomGKaRvk66Q/6s7kOIwPs+feJcfIRSxTi0IL3//hxNkSto1J3s
KY1w+nZPaMxn43Su/1yqwxTzmJ1GSP4tu8jJ7zpHZh4UYzJLrAaQBvWEZK3b7lfb
QMkuFDSEfLlVdwRa5q/FM2K9n0fcGeQKqQWPv9bQJXmQWv0Dph1QPpzFk98tFG/2
MAtc3gA2UylKRgLoDBsrXk3MY04js6F5bMH3/YbbH0xn9zS/xfdVwqIlKwFO5KRW
IPGKbWDH8UHM1/l7JrL4hS2R7cLfEWv/8TfyKYxlukCE4r9UMvqpx+YSqWsGxSkP
0hmNJiTN8hPPxWXX4IPsjJ8BGyMpThoSvJthgSMeXGccDq9pVdTCIc0r9jR/e8+D
/CgVWsYwCoQg3QFpbAV1X8XLTgqdrFXCS0XDB9PjsRrun+Acy3wswl6HubMJnYQS
rVmMcN3tkaweu7ozyD8onK3SCxwZlL8NJnJ4mpFqYhSAdSeDiCcySzbPfEZz+YWS
gq+tSXdbrYVM3BfBmcQ1UufYNG9LnGDFYk8cALZnseEs4Y6P/b8lQSKw/tFmCCsw
c9j/sxhpgD/siBmiXXb2FQPyKdsluaId+0AKLidAHzVhhDSFXBIxxR8Hw493g05t
tELLrkhGaG+at+ln8EE1ttzlxg4pMQ1vrCSYP/3LlAoecIywK+r5YWYQkZ8ej9VW
fIOO8fmVr2nqUarthQUk4e4M3Xi47QsBbMuvKLnwfIjANh1KQrvFznnwpCZl4yT6
2gsSdMPLzICsS5E9gAIQNHIyfBoeOFARwhQ/IyotFLVsILzybE4U7zM0RlnOhp+0
IS4PKJKNHFIScI5ULI13wt/9bDuVQtjFbN7TEM+++EMZd6n3SmOsEJ57gQ3/bc5c
KGFHFh+G1xs4a0zKL8JAagDu5OxJ7XGoG8fAOqASWUIAsiXoHkdp9/yflid2mOaw
G0nBqs9ZgLTOSwFGYfaX6sRMB6Gm06kc6NU9bESrEJ2YQat7gelZuAtndxLai5w8
xG9JV4OP5WJFfLVnlT45soQTOFl5yLi5TMiHfyHO4nn3G5ovnv73JpxrO33ZBs63
LqRG/UJic7NKNZeK2/TlllbaVKbDUFnTLFtMg64WoI/LWLqfudPT77bxVAjK5jPV
t4CJh39TgifkhvbcGECMW+uLfo7Nk5970L/6n5pT0slcpcgKSbwkAxVn8NEwGnOD
iBI0hzDbkCezBFi/oiiHr/lk479JljXxUDbxW82pch7Y4rwpmI+99goWW6IapW5c
18joxBTHFte1WC5BD1VMbJYkLzye12kxNeR2g7827dFfRQ7oS7/WcSU57/PsEkUZ
f6wg1TLgpeYGMvivgJEbrOzMmAt7+fUelIvhhkwPLUJVwJdCbXrzNNR4mvhA9QwP
8ZKIvJYpmRH0jpowEPc/UI28gZPa5wKYrs90q9qSxaIRJLj31JR8jesljx8NmwED
X9YFUqIn3+cE0jSjBaDoRJLKkv8peF924eJMDlxqHuJjq2lDiUGwQdeVVTqJynhv
pxjIupiroJPd2kFTVM3selaEGnPrZLqqAk+jNxiJw3X03tEZwIKnwC2SW8rwXTvg
PzzFYYaYv26aXb+4gagblVDl/uKZV4ajPxE7xkqRM6V0oE7Tqw9thbEuJbtc3x5X
+FNxI5WUAzJ72d9IlUELtFO/z8rZLL7muJEPLa/31EcWyNR8T68pWcLwLzjCVfOu
jl5sn0aDanIOhX6LBXkbbpvgNMeDP8ncMxbMcjjeGVkk0Cs1uPzxS7vXQ3xfrxbk
2Fet/fDOA1TjaELbE/evcwiprm6gz7jQFcJyZ5lf9m5Z+gZBy6k1fo9kszHLmz62
pmcTMPlv4Qx/duAPEMBugO3lUlSKV6e0P0Gx5EhcxXub67MNUgo9V3Y7/oi15j4Z
xkhCjdq6FBCXB9aPmehh8aLNBwFOz7fnsvgsChz9Y17Qg2GzeXUsLAJJ8QSyzvtf
eX+N7/2PP/EsukpHAmrgA+Ly3Ul7Y0wRuCg2KOblO+A66s0RqcBWMhWZYnRhF++f
w5fs33Drqtmcw+b74iyCxG0sMKp9zQylV/ubYIkBj7WiIyDItz1udLRzyNhAra58
JmaHKVPyHg8IksAMpl0uBTEoImmHhiyu+PYxyksXgJiNYnBAdWcsXqL9hje1L4Bz
55ftb6/L8QthejOLhL60dbGzDSH2x8qfjWkooMHz17eQCkyrDgzdY3bELeweopTW
2urQ2W5ZtqqkCxhk1AviqwsPuNon0qDJfpDHzTt3VPvGqvQ0SFcBcSuDPJ/U/I7W
ZOcHVToRbJav1ks40ogcVF72ajUF2QGMZVSJEXUPM09+zSjL66DPqan+GnylA1bR
qrBIcm4xgXQjYhsWarOpWjOyp2CMTol6gAqR/fRbsmFsA0+o/p7CNEEa9AfdCy3n
maKlSg2GChwdb2ZzcqnuYTuE25ZNYl+8sGmHEcHSK8WdT1RsbbgXg0ewW6KivSi9
PvLBw5BmgrNCre/ZDSsmF/o1L9KpS2f9WOTNiOpjpKJxhRFra2qUtLl5GzfST4jz
xD6Uy2oG1wLEEoJu9You/rNbOw+dbpcGioke1SF7J5smS/Kht2gzDo+VGij52efT
tgErw78FF22cVz3rjMCCPqoVLqixUnLNI/5mp5UyTBSVMleQhoIuiQ6B6iCKd0CC
uhCZuWW60QDQv7akDKxO6o+twTqqyaXwMFhXpCg8egX87yZIknGPOgdBbTtGpkkZ
shb769MN/BPRIWLCgKodvMGKNACjcvcVNXAfhL+hPBdNXnDO1iqGX96AQIg0Q+0B
ZymLHCg1ydvO+pvVnLm4WtkjI5jW2LboVSdY6VGOILEn8WopxbQs4p3jw8iJ4M1Y
uaV+lIyLrB7qSfn83PGjoro5wd7wiB534kQ0+cyiHy9zQTEn4sQEB64+bQ5IEYjD
ypOWzVQzk+h6WCm19o0hJqMifH+8QwCQdtRQx/4o6WTlgyNPA0w1Jdnpszx4iFvR
p/9BM7+HvEMg8BD50fjgdMLC0OET6qloBAqO6VDMiaDDcjvssNLiBQ73t3/pyPhQ
XPTxXgSL/5MCHjmaQ6S6DMkH1VwsVuUEAj8zRgtIbGjrAPu5VVsAjSwGBDdh6+oy
tHJS1cZZfOMD7Ivjqnb/zHt9/ZFGbfBE7zCkdALgyuStTT13ja0Nm9qE8w2cDTRh
AdT3SJBtBUHXFZmbrf0S81iFqiHRPfHX+KjheOFmBkqmkswSvqZ8VJKVRvWOFzDl
fWvPaEP3D6RTwpbxYD5RMVk5q+09ndUeXh+viYCWTsg/Zi7Yo8Ti7ZsIArkKTnhq
dav5kwzwDQKqHoCzKSojWulqtbA5XZb9zahCbXJW0BL78Wdvs22h764bsQjq0blD
jyOR7FhNEvtvkrOndUKgyF1/EmmnvnOKgmWyKQjKqfU3Cl/KN2a6Gsx2U7J+cj7v
NBNfNi6i3OLqOuyG3Lb8L9pfqc3nT47GAD2SX2MisadpTGxBZwx3kDwizuwY4OpM
+90gILNa3aLbFN8gBV4Xqcebvi8Z6nGmbjOIef49nc0bZJVHtNylDKiBsVs1dksh
YFsFF450zcyj7sy+cMPeR9qrajEIazg8ykrjCmxh/b1CODDL/VNdmGC00uTeKZvL
XZCsB9KPYyjEpJUD1w6XlWpuMJ4U6sD/6JuTJMFGRfJKsRTSyPuf/hB4N6YAoqes
ZCCIY9fkz/z3po8dTVl3ofICiQm5APJhSnhWP8whyKzfjL+QacaB+iVp9uEy4D/E
9llOE6KBHVAFlbvFg6C/mo7OPFM9a3ZExSSFX2hRmZ2ATEF4Wr2IZD0uxQtcFDSe
syzaXbN8ji0RzQhcDw/PwuROsh/H3CJeDV97E2snFRTTOzUTTWdww85LyqK+VajN
QizYD65Uspmojpfg1BRt/eDICdVwc9uFSkfVPE72ZqgiZ2k+4pMweXb0jD5ec8ED
LDmg4IjsPti2UGEDvwrxBmORn0NaIv82dJpTRmf4vsFTAiWFwjhCil2fKE4Y0BZh
u9gD9Cppr2Pi5TonM6QnqvvsBK2a+HMySkUBdWFaG1oQYrduEuBQBVdUiyInfBQG
e6mruDpeq36H7NY7pIoAuwAkyz8gXfVoOjq15ymgg/viPfDkIIPlbz4i9+rVZmAQ
19sZdYQG0PSd3sZEY12Jx63sXvr/E9MU2ulKQKlK3qqJLqs6rGJYyI2mrbvAvxvM
wcUPmMhMPY2ZMIeKykjXNlo0j0hLqBsgEAhm9QhuxBFAgeSs4nmTkvmtFKOQI+5/
jCVDCnD2ylG9QDB3X92q8pBiCaFHvsXksviXCO9yTUup5UwhZQVy05QXW6Ki08HM
xMnYIEuPKCtKmIhZppWuNfC7a9TAKws3bKyQ2bAz/089rEYVuAu6HYGGm2sHq7mG
P0wBAYz9ZJcalSmkMeu3ncC6GOFAGGlZmCPfycjrVoZ4J0ATWb9/pZf1Xy9MK94i
uu0giy98sVPo6tT2PgpF/tV1YWZBsr6V/HlElBEwpol6SWQOgvUkMcw5NrEakwTH
wfzFhvcqIGJ25u2dXTpa2zCW7GapFbpiggvH04ORISrTXIZi0krPtlZEoCjFEbUQ
g5+M1Ikao/xJT52yUMS4px/Bj62Cs0k8bWnlTAyjUPfa+y/cl6ejwyc07mpqdUpO
MI4lGXWohBaCvzT+dH/1Ye3ZOn/ANB6obsZyLJmAWbzGUOdExMjMjseUrJwq1OOl
vtmexljLJKXz4GfvZ6RUNeQC3TFxXrKOACa7dxvM2DFlq24Es4UHlolaAgPPaOE6
By9ez2Q3SACmZvIgOMtKNI/hpcck/+duVAZLDJCuFF3OnqC9hCv8maj+3nIx0kXY
H0FtusoFup6uYhkRZK5K/fvrdfyDDcK3CW/niodPcX2qlMdFq+arDrfeBrViYdlb
UVpA8DtKl1WN00YkHzqKqpRxI50QOF1AdOFUUDIO22dJ/QI8kmAV1b/4CWVZQOhg
kyuD2QfqPUTPcRsv6Ym1jUMHSr6MufWx3RfosMWWwAwIwTg4m+XfUaFTM/VpQqbh
h3WXX2OXC/ESoTJh0rQ3AhqClqsCNEZ7QluHcz3ffdGJxdKqhOLsCSei7IZvWUu2
gL02Dc/8nljLZNjAz/1f1UDHSaG6pkPrkexG9QMoDg9GyCdOChgH8/PoOe40uYt1
RrdTiw124dFdNeICmOWpZ4wTsu53yay00vwqP5YM2poKv5JSqoex0uNv+LqUOSGL
cpNSJSIF7MjyvdcYN47dbEM+Q5tixkZh7CFndHwDEHFhy3Af0YIvXaKW6LlCy7aD
P6t3nFGEaRRyNGaW0g86mL4nCNxL9c/t+ZDgWVtFGrNeuU3dd9lcEZUFNxIEKa/Z
GLBBEW7wKHgHXqlJHyIJZWqN+93JYPtSaeR7pHg2I/qY9wUAmvZn/3KZYeFB9QTa
Wa3hprdxHO+FddVzBbTs/bdDa9WXwQOrbnh5kYRKc31oBKJPAm3wXJ4bceTPNocs
4alB8ztPgWR2hy4i1hx3qGmg0KNAG/P/WV+VWHU6yXZm3QwjuugIj1w1Dvj82Ocg
cxT3Qi/mFbE2a0JJjuUGyY8lw3nljoUr74c/ZelNdP2tbHf7nVZBj5K3h06l0lJf
m8OoBfK3+5/dVG7rMGX4aD/ZEpc1vaMoNijI7rYk/vR9TBalVQ41Mt3OglNcN6kD
mzEAyD08bxJafNPn7rUro1U1+jH7QYxlCWcvwggIc10dMduMyjv44zPVsXAtg1iy
3n4LJvlBC36sloxAfYWHtoQZKKBeukz0w7t3AL8c2fQ/BGEHVQh1IOhoxEKqQrHU
0ZRlACmMH3itC4bDyaIHjXfcXxlS+VZ/MkmF3FRF+bAeOyRR6sncwUz9WbI0VuqB
4HGzO4YiOB86gXEmLogoTsNISsHIa79SY16+1DSvZG6ydkPkxGIfaqkhpIRhmu/2
z4kiREkWPmsJTuuNEjIoT6qGj+rthvzdGwVMmHOw1oN7LQ63aI/0uyP9OIDxkOW4
SpTRyDBFapdBwAjD2cN5tcoG3NhseAQvx3C72T0KDArtRbO7bcriqkCxXgL41hQL
bTkU5djrEA6zejeFxcvqlY8ek2FVsZLu3FQeTfq4ZclQa/caS2cE2xSCnwN+kT5L
jZ/7lWVcRYu950beaTuHlROxYg+PkivCb0iVYQUWgQ6+XhmJQf5g33ORQ71w75UJ
cwr+4JXnEIsSCv5cqsDSFcKPCbXzFAHv8pJB7qg49C726HUau0Ec06vuW8PqZ82x
wnoBZ0TSr7o+xyZeczcLGFnd8e3qyE5yO9l5k0XHRpGlqG2Dz0gQrqdLsxZtseGL
QgbzdlvQIbcr8tBaXhs7VkLMFYYejoKAmI6plcDUHGl5Fin6HikJr6UhCsPw0I0l
2ZVEJ9EMqgaEgrEUPqAMU88C5DLYoXY1HLWi8b0/Yt4sxB0eCTpQRQO3LuiqgBPc
AZijHilYDnufek/6E351fQETS65SITQtJvIavyf4qANuhLCEENdVgqU8z2MSpfcm
slsHKOAEJtWbLx5qzQ4ehaAn9YFDpvur1vJveAa6O1OY5RvZ0JkRECm/8orDj4Rp
FkFfRZHexxIs30iWAPdzxEm+g+vj0jlEIy/N+sWmO+HCx2zvIGRWkZ2dGpJUBIrF
i52m5D/hidXwf+DgIPrcMDiPrRAnA+cBqo4HHD8WA0hUKedPLy6Jtx9ODyAMS1GZ
edG2rncyVxRqUh8Pttbwa7TLYL1NRCa6wx4g1iXso7ltNGIdHofXUEiuAtXVmCC2
7/3dEPYAiecD7WZmEH6pOUfjkOgUf2SphVRrjshNPEYSdmhCAXfR+l8YzzDQ3gTi
p9Q53EC/nZ+uzDe9WHEiUZxMDojM0S9o7PGi9BXI7IZWtYbJhWiux5ojz/nuLvFR
fvRUU92DXLGR/3n1RU1fhZwc154hF1OzR8upnpr/waGgHQUmNnJs6twPeL0ITqEW
JxwMwCgX+gFp+gOnwuE/QodHVVgMdm2y6F+JAdmSHUIP9oW1tScwYhtIp0pQqC4p
5KF/ZY0YZ4mrQ45MpHASQFc4MSthQeE4HF4NRsqClexgC8zF8ozVuEUCVY7SRw3R
NyleZMcCQr2ZtGxl4tvhWPzerXwKfCtydjj9qYo1NDR9aHY+MPRU7j4UmcxJTVRX
/Gpy4YmEu12/sDDSXeCzDjyBx/Oniz7TfJb+gazrx/CHqaSJrJbJBt9jtUsl3mbD
J0T2LZE8ZCMr3to+ih7z7YKhf6vQGq02/Up6RV1D2PSAiQQ8j493HNaS84iXfB7V
SlmUeoswtrn+RHVZ4AA6dJEV+gqPEHa4fBe9ScvA4bD2FYUr7Vd9Rujb2/Wkp5KO
jxDaaK6HfvIMF+danO3dBApJvzaebelgT7lA7qB3N0xt3N4YO6zoE8Lil8h5vWCI
jQaB+gtnLswHDBSe6shhXeWuagvv+6GICeoKCtmMU11TeeEAVOafJGpUHrI2yTvU
CoQq9+9J7Ype1x14lO6ibmQIfx+mOjKsbMQVxJsIGHSILHUZmRHjFEAaQ8SkIG4Y
HsyatMVRBnEfRW0D3lVHQoFLyHjhrjnkJgDp0TQb5eqIoTFUBk1Sbj/c7PhB3QnP
wdt5++f437M3YfTowYS0sGm9v/omGRY5fcWHtWZNOp1RA31cPIy099xEzQtxKBUH
f9NuYRlDFJ74We2Bfd82IGwsXoQDAgC7eXRS1FImqXi4Ejsy0oSBKs/V6wZffPz3
OFP9+tYWQPATTSPOF7iw/6GiSTntIiu3FYG1Lu4X4VJYjpmxmAuCskXaFPNGqa5b
MbJBVTRd4vWlezE02nm6f/qP5q4isokAhAkskZjW1X1gHkO9618czMiQAmb8sKpY
bNoeJ0fhafgdOtY9oY8/MXTigxbwk2cxXpBtH3pxGdqNAFEM1OehKULARI4Srkyw
7Ocmxw5BNoE0NUl93i2j/MGHRxP8QsplFOQCCuNb84Eg3D55u9DdgsprZEQsP55f
iRUoKRBGIBG9kvNPzl/qaaP64qPqZGssA+sLEWIwk9/Jl4+kTZ1gzK1YClrg2+RH
sD62mULZj//kFypDLLJeRQZMAVYv9OTvh/dLShWvqIlxVMeOwLWVkb/Hu+MaYsiT
CLfLKZJSnPueDsmNIv3MJK9jf7admDovJ/zdKq/Js4Qzx2qIzrVolutC65fPGIp6
mEIz7+uDV91BFmeIAoG6K0WjkkhRirzlRhpjQL4+3xZAxUio3CBoXYVIFOSW0CZ2
ORPpc2ekkNY3k3lb21KZpE4kl7johO7QDFxs2+0ov0qvHb3YGMybBGmLv87aT2zs
D5aDGsnhZQgn1r/viaUj97GIwNFS0knj4WO1rQItxglQZchcFIA3LjOv+lGLlphO
ICF68KJyfqTP8Z/MJVTYrMK0W5xjF87cwXgFT+1317W/QL361lk2HMaLBUq8Y+Ci
deks+kmJVAlm7wD6UzNZ8K1Au4ZmjnvVI0jZRZZaMGBZMcgvY0dE5Fqe3NTU1GVx
bQ7BROaFTIRXLdDLNqWeHbW5BUjJM9HMHYQ1JYW9AeFKT27wLCTW5rsKF9DeKPjS
Yx3FyxkM18f5ofZs7oe6NQ==
`protect END_PROTECTED
