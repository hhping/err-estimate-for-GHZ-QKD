`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3uBUqTI4skKfv/b5DzjCtutj1S9ipXfDh/giVtbz5pPWe3pthW5TSUBLq2xOli8e
IfvBF8ZP6GAS032ZZ75f+bPEyAdYf88e4VNdNFyrJaaEzt9zGjLrCoiNagY7DE7y
KZFCyGjrdseiDPsMa/7jEpKd8FrW4ef9dEIEWglSOIyFsKNnHgOIlqLfzkJNuju4
bORSGCnCZ9fZjpcwhq9EVt6hySxhaMhm4Bog2QNt1U2zMjSxM2K+v+Z+60/QqZwM
n6ImDVBLDQw30k0It3kkmzdR653DdQa6oCuSHrzVrOZMXCy3qXso51V7V/E7ibIL
Tz+EMRoZ5LXZRRrH4lYO32gbu5sO9euolKZl2aZxfUw0bN85/vmeWdCuXCWPlUx5
J/glBISJBtwZKSqGbt7uhpAzgGjkeQeQXljIdBhhUlOECrdlIPvIZhCsu4JRVZ8r
Ldv3zOcsOu4VaGEA+wgk8K/M0Id++8Zl7GI+nFhyjvZXvSrpBakhNdQ5mlcDEQd3
oYgkxbFz7hIMn9CN1WcWQbpQAIhpv81ETiK6jiuJ3snsGTyE7AoXPm7huB3ODmnI
tuWmMJUXIzj2gEJj9IcE4C3+thpaenBt7Uv3B4u3FtMivzI6DTNq3JXubCwXuIuu
k5pinKgHAst83o+nCDrvPQEYbdvdfGNs0Ux3oQVIAXqPffBl3nH6o77VwmpXC4M4
rEs0cmT/iCl/jvOJoeZhqikMG3CijgvvLt2ivcZzvWdJbY9XXaqQvwXkY+U80FiG
xg8JAyJSfbq/M4uJcbFuvM0KpzZ80LOUDPrwvbSjEVxc1ZeZtWYEOjxb4oPbrZMX
GW8hcd1DaHT1oLU9TA3fN00Xrq1WjxZVEEv81rqoRWlIXPvq3WSMICFPpmTIk2k+
rjTMV0oJxH+CSULVdOR2omoaPge+gCotGd7vg0F+NmvkeN2FqUIGcReSkHF/n6D+
iYyQy44UvyBKuhPh0V7ICwwd0llII8/dGkR/SuGUKxSW5Rl9Z4Nq9gIDJGnY+bAO
UHMK/DjRHOC90g9NA/yej/SzXzvS0TRpOEnrtlCZwQUcCYQg8Rwm/CnCIBAo1pKf
uBhaFqjm/5jwD/ruPj3ApTdDduYMitl928CvahHlzXICq+nhLYGEoS4o7LIRBhom
Xfg54BQNUARtp284O7ucWNDPTad5dXAlSNtCd+3ZV+1oYayCgMmNh+yY4j51yUiP
dDGihZ1qoJYQcjGU2m58IdRa9hzt19cbbX6B1B1Tckw4PKViVCFYId57M9ywnUa4
SmXEmo0L1gPZ/woajQEVuwvzzRDWJ8M1EdHahFiwV1L68yCSMIiyxj4+19L9DGgT
vG3ynj8orBG+eT2b+UCCYLetUJ25P59fEHwoSzedPpAe7glkyAqeKhOrDNn7jC31
S11YOJdnOGaMqzNNQflbVcP+/29Rm60BNI1iSdqepi2VECNW9LDTs3wWcRS2UA7N
r6qufLYH8uxoX4U2J9Fyh+B44teH8VnU5xgVjux76ZiyOO6f8HEW0GB5pommEy//
3h4BvioC310pbQyUtKXy9NWxoN3pviXVgZCweaStcASkr5q1+0pwikzab49Yn/79
MCnKg3tfrROCrSpJEdWxnoem5vuqJ9K8wzAY29EUfMI4mqlGRZxRdbDHUij25RBR
uoG4jXl3S5BDNt/dihJjZdAWAN9T8/XowYTbFkp6Z3GSyS4Ci02SXSnILFB3uNVn
3iwerRQVn2lhfDNya4U2KbOUrirc2yoh8B2koyurD9wlxEsn7AY1PXW6pHsnITQq
ieaDfSfOAU21WaVAra59BMR9TlEEzPi4AOQTS+MZEK0oUFiBOwmjVHar20Pjb+iz
PquK+urp3iB41zvkWZCtrxQadJUnYOVkT5AAJNAv74Pt2cBBx2xMJILaasFpDuPr
JQlumcOjbqvxWyoz/vjQER59kuZXprAbvVFT5twi9gHUSgwvblhDlwMNwObwTfvm
EOQHOMiIVdBvKk2x1+ZmMZexJtn4R2BLyfm5v0CraCzdvzN18GlVmloOuLztVUeZ
uYpSxOKoicKS4pVbvfGiQ8LnJeYTB1E3I1jqO0mYXVg0CcYMuJTwHGK9pfJ4JSXE
HxwrUPWVfmLW7NL5hq3ODGtoebPZibxRcxSEp8ZonAFKWP8bQLOc1YbPO+1DGNpI
GLoTzJQ2l/SQsxyasIZTTy+fpSU+SihiCearULTfNsWJdOoAo6U/4KcLW7H9b22N
26wvIoaLTll9YV7XXGBR5w==
`protect END_PROTECTED
