`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgothmbvqHB3kH8zyX0G7OZTQhjKSSXh/AAX38vJHOByAM5la+3yDSYApQOYiB3p
qUBQyb5IEW+H00XST/OCNT3lKV7AgHNo9a/CesCZcoB2c6hwTUfoopNYVdchO5Fj
ukxxZAHNvVnCTE0afoGa5lClsPlBV0FnshnLC9ET/41Y3RMONahuMyErV/kwo1rv
8DxR+VcDMheVDysG17IQsF0LnRunG0gzefMw0Iy1Ic/f0oobYU/FGrCg7M7XLjQX
TTxKJr8/xyqoRIxqKypvxgSKIgBJBkr8zwkViwHXxSh+b5MYS1sACwRqQGqY0nNv
QQYkwxXV2QgMfHU+qwaZ+IJgugV+1PXTui8AUXK3yo6xbceDLRo6wmKUsmAB+Ts7
eETVa2exZZPxgBYhGqyIi/V6h3JzU3kTF26Vjsu8kxTN270UsBhlMbfo4pT7tdXO
PFsexoZ14C8axHk7p9IUiFZHcV6K62tqKxNo9c+sLC4+JN7J6BSWZb5H0kMCT4Nk
0wmMJuqvHT9Ovk7/Kp3PvVKkYjZdRojfq3P9s25HgzOnbgtk9zvS4twvQWa/2fIr
Bzn/M97KHitwNC30sGJCAo8D4IFB0ZG2wsKuk1FxOh5eAqDWQrmIEFRr2Pj63qdO
4o2fvOETLT+C2IhRu2w1giI8OhdYzL2zaMNlEeIzGIENS7N8aQs2+SpZt5kfTgYw
Oujzrd0I4xZWHLteNTL73KcACotKHAUO1QcHqef44O6vfc5t6eFBDbdj7RBtKlf6
GYjxL8iZ0cC2JUXjb/TwBcvbaESFlvfBHquiGn11GcbKTRPfHWgrVIQT8nc85/6x
s8dXa7pdgoGNS+lBy1KDpIhi3xkLk1LqQ0H5pMRNSSpo/VjjIe6z/N0+oMf1tKkJ
E2qJMun4L7ZVeQgbh7hpmkiTY3uJyU3ysJiKJyd0Q8H34NkOF7uIvMnzG2sOBANI
T7axzVJRiTsogEh0nsrcS4w4yW48DP9jXU3Eita2ucQOznvXlT21POYVoPx6NEc2
lk70DLU7/aT5dOzjoFDTFOU5T8v/mm3b5tnzKhL2thHlLjnu9MRUUW3ZIp0OFcrv
doP/TLIw5Qip18mi0lvtd1YVgFWr+pxNT0nEvVj2gVQvEIgFtrp7mXfgrPcoFk9x
7nW1iDviehD2ITqODkwdPcSu/r+N1svmSDl9u1Vm2pLQfTt+7e/pbOlRjOco+ViN
qKa+64FrxMn7kZRdlTxkRS/uMe2xK+2z6krN1RXzWD6zS6tmoZI0qMqjDMk5Q6XX
qQWjnIyHb6oPKbpa3fM5G0gpTvTAiLzgeo389RKX5M5LLmb6tt3Y0v/vFvme1lD5
RRbwychb3GLkK484MXe8zfxKVSGwa+37hnRt1W8txlC4owOgqTkbMqSDWzQSpEwN
2uJL0sS2GyeLkNVyL6KiiLSKuoLPdGg7zPi50e1Hmz4B1hnLbILdCRSRxtXZPNJf
jKXcmEwJ5FzQyZ7oQ6If3FYbYOD3KWMwPCI5IjzeJdYIeMvYlTU1kIBEX5HAW1so
qNTZzrHMSGM8MvBsFeePJiYuD1GGknNxKXvHuaKJZj1SHrfR+bFKC5x5ssqFhrqf
O8kVglFyVUK5SBFkc/psqiKq0Nxo/Ye4khtxqDaeWVpsmceOpoU/RAsLC9C3DYSU
YG94ZVl/eO1bWF23YUYsbIFtT3Gohtg2wfsPXh+WDcxRcJZYl59gDGn3tT+gTVj4
cO5fX3xeGTUO/b5QZYgsxMJKlDCMRetHSKUKDl8XdO//+GsTjU6pkAduQHEbpmbd
3lQfwIhB2GWIekTP1FcCJhtIGmwJN9W2Hhe/y/4ivXlQmzWr1e6SIW19udpw0Ck2
mzGguqqLpshnqWaI25AOzk6Kbjf+YR1ZJyXa/kYHEPzNF7Ui+b7IvO5R2pIS4jKJ
K9Y0rYvMtdNT3Nzxmo+QqliPF0TLl5AbaFcB1CvMHV5biCQermxkm086m3ZbiEDV
/s/9EZcf4bsVbDCW6dSpJMn5H7XzhreSFrcKS0+sQ/PWe4XXvtZye3O6j8b0dCZw
zzIHEu3mbJfB5FNwjwVlevjIerj7GholgqwPVWB6XZk0aVhnDA4eXgLNVEU+T/kp
QQYObHAJ0JGU4gMFdyfujV/am37QdtT99x3vVH+cOjjK2l8Kx8ZXO8veu1N5iAEm
UWDUbrixhJwcPuadA2ABc2cEJJaoRdZt2LMsnEmzifIqnvciUHwQSImNkhJSpi1J
JDqZXvvFtgddB+PDHIjrQQVbHVUibz4m1WOQ4CVGjWPHIH+2sxYikeGFCScBmXq8
erpK7HPnFI7Vvl7COox2A/+wUzTy46BgVeJnMhpTNsByIoQ/MyUjp1cTJfujhWo+
gqvn2scUlPbZ3dsAzPumv7+f+BOse19T5Ps6rJUzWbKCpb4ymmv9IWwrWBZFu43M
cAuIIsIvfCTdaMhZaR9r2/79roWq+XiW2fmvA1AKBkDbDICmE1S6yEQi2ugGu+wv
CZ08F/NIVoIw3ldvNe8NL+1v4LVhwlazGk/gE8gcT9DsgfX8g1kARTg7MjVKy6aN
bUj50V7miy1406JN9usPbs8qgj4hqgiJYOXqekGnbH2G5TCBpMO2EfXidqVgehVp
1qzeJ87EImg3lt4fZEdVQNyTOl2WSAGWzhwJlzgd17pNPgT0NJBKbax7Fwz+/RE1
K41RYr7wYXoRvj98crpI/mchxMH0UuLOrk7fe04lS6oMvjWucyDMcl7EOCywj9aK
q4Lajvw/0Q2ycAUAw1g2PSxXkf15YceyxMErp6URWbOt4MGU0Jc8a74t6qaYuLme
/Xn4n1F0uzNvvm/l2EFVWZLBFRciAfge6CkiCdi9h3NhotRZDE/JQc3Xtqw7iKqI
Ri0qf4l3ysIHdFcUvmGPJEEZB+N3Q0o4tr3I85Zo/AIAQ6qTqaNTQ+oe71gRwIb1
jb9NAMyxqQBZNvGTWNdd3ZGJnFvSBEl8qjJBMFsS1B7aKsgNFGxAkCu1VdKglSfn
DJhbgEP9SYEOENIxJPm5pAIie9ew16f6AgIajQDkrWq1Lfv+TzQ+tKqPcIzwuBIo
cRTO9cO9XkM2Aa3Cf8MIVeP0VMwoEAiEbXw4Gu1kp+g0V5WBZf0A40A6kBO+LwPI
ashWjmj5uD6VDIQpFoHbgvKWXL6WeFPR1eWcfkl+dkGJV4pymzMmEcZWvfpmJ6X1
GWWHwzEfbV4DGWenV5Yx4U6SgD5nEMCS9/IRRR+cvTfnwhRrUIjRZ5Gu0DziiLGn
E392GlRxpHmjuyO6bA+7lPd41wyC2rBCRBi4U0/m61b0Zw0Zn9smUj+JAd2JCclg
gEjvbK+83UOIhyoJf/lS4zHT8zVhDMVg9wVaWL43Ms8VHPLjY9pia5cdPUFo79q9
2JqNv935fqqzJe9nOmlkkE/Rxr733EqI1nzUp0An9+tTxVogKAhCXTuRrbLPnhx8
WJ80ZSnmfmzBaPxTdPAUFXMoF/J351z9VV88hgt/QyY6hIRNaFdAq+wEhWiAHIp8
fHLyUgonfg2M2qlQ0XAQqztYR1dReF1+UWjf0kisKaZJhbJQdfvfKkCMfHTeNfiG
aOUCv2P3lUn17ZFgR1rIbRbCNWVyBPSeTk/dR1Bb4sAtTKCVmlkxakk6xzST3snh
doFbD3ga0RLk9pYXNSmOzAZs91x5AP0YQqQbxeezpjyenedpD6kbSQHAHB3HwPZN
RhrHgyIryrkRvEG/bBJh8AXZkIQsP+YV8fw6XKqQ8c6USpivUsSSEsH/IPG6OQcT
R3et+DttVbSidzWYOqslrQbU4brbPTH+bDdkrd60ixR8F4Fe3KO7JRBtEcz62M34
b1/t94ka80TwBQHdFsNcYVb6fs9d4schb+M0TNpwAxCamxVNUyu4z3bezUtuR+/t
sCqRxOADsUQwUBzcuvGdKcvR9jpeBMh7sqL1z197yu/bNpj1kb+oORd+Pzfgtv3G
zSfQh0PPD0l5S5KUmULe4P7Ibm/mEuPjXG7HrMbGnul1RBZm7xQnwQ9Rm91rynmu
AHXENWxJAZT+nQKDRNSyslGGt1FTDkUUDfSqd1gE2h/opn72+p8+7XZn73BUcbKW
0iEMiJgJJz/gTAEE6fns1kqF7sf4fAbZo6PHPyHZRferQL8a/yqiBuzcyDDTR4WA
+eSW85zYjugM+puT06XXr336oTZiTX/bLRpxjMJVB0WAZ7nvyM1X1GtEGa6jo9CW
`protect END_PROTECTED
