`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOZUwEfi7DPdmgBbFgFbxnq7NMNf9T9U/3OL/VvpVEgyoKn9tz3PinLNR+32nzsB
h12jsnieYR3UaPrvGGZ60ziuPn4yNHiW/BDIJgKyJe+1eABmt0skdVUjxN1Ze6rq
2YPOXbZcFgCKqdRxkw8qdU2xJpEsEuxi7kZ5ArQKDWoA66wNEhh+yhS8fh0kZjz6
Z2LnTjk8yhFidHVASKJs/TZbbaIhNdnobuFdc2Kj73s7zKY/NIEPX4Z/KtOypHjp
Nm7PhWMLiRkp42wM/OKLY7bFcC271q75IQ4Tlo/edmJJ5dtnC2cVpfcmwGLOXchP
JEFk1tmryxU2kIecod2rhdvaCHlRd+DpJEd9J+dVsWj3aKzr7PgsQi3sAUzpHu2L
8RxEwosGpKKVMw+HRRhB1t6Oz0pLGutCXp5pbYFbcd3BAWYiaNSpI5xqsHl9b8dr
w3jHNg5dqBwgHAWbQyh1DuUsv+0CJvR41E3pkp9orCy41Sx40QtwREFLRJqWKyN9
qJIR1UGP+8Kd9CevToKo+Hr8Ej9PgXeCBnTBRnvyAdFDUW7eL8sYHywCgCeS3xrT
KeZcJN2aHwg+j/0Cp/5xfmaWIrgoV9IZQh5H+ToQjJcAwwlcs49O8LGUdazgqkJ+
jLJBitqxUgfYaRWDwqUjwYErdwhWh7QWj7Wdfnh3fAkFM5KMrZRwfa3VssHU4AGn
XWcendbdXPzqs2Ns7t6Ep0Vv3yCN+Zh7+I6Dft6rwhUsOauUZEnBDpwZQ2i3b8Bp
Fvb7x4ICq2GovDdtFYxC9zYTgbsjUDjwS2JHP4dhNopMHh46xuIz5PWAYuFj7shw
mS/zOSn6TE+RQv3cHg4ehfWIMIKlpxHUw9BQmvj+HisH5fybzBmQviXL1Zng5aWJ
OOWuzud2Mx9L1MTPcnRk8e7gKtt2QlNBK/oqOJ5spTWBsBrIMGOuEjdjOp/4FArN
0BTv8W0epdIgXjtQqUpuXwoRgI339nduraujmEfr5A2pZNX/ele4yb3kVL82nK2n
NDNdhXqSSn8Cs+CNVsUIZkCxuA8UNfp8VPG8Ogah3uX73UkWHnRjEP7YRmwini2w
SPKyXEvF+WeR80Www/qbYNwpbDf0r8PFwHT+M7/Sy90wrvI9mygXExfrNoStb/JV
ws4HhWBVDVR0Q4LzA3VZRM4m+meqlrKjK0IPcuehi1CBnd8FKdjZ1lEtfxZIItu6
Dk/aAeHHNuQ1pOSuJQIjct5rg9YpKKnk8qHE9dZ/H0wp2PteCZwDvSjEv/LsVsIM
VFSrpMxGE9thiCXCyZxth2TIQCDWrW07nGgESyfPoo2JV9FShmknJTNUreUnvEGx
i4fZ7pku7U79B4pWTXc7f+g7Q5z4wjfCG5PAo3ZRTv4JSx5gPWD6HB2jM3/uXiiI
Xvx0rNgIpLLw3UwpH2g6408/jfzc4LaYPRxwPr8z2zSO7Nxod3CYBHM4K8yA1zuF
M47yYVXKvvizdE5ziTunZcW2LR1NTue+UHf5nqhbo6I3/SVXDPvQafIBohrIO9OZ
iP6CGQFHVaDqhxPEZkSfpmt1j5oQrTHBMacdabj7GTNt4gPxHf2S4CsDe2n1sjSB
7qRnulKUjv38M3W6fipYPXiIpqdSJy+A0jFk0Cfa2HB4w5tmS2P6jt+NM9eVkH/x
SeHh9K8j/GZuukOXRTqaducu+jPfIJAa4VlFqqhTFnHJqgu0oCledNsNeAgO9Bwz
M5aRfKXtWIfi9NYVDAhodwFE0ktmvg7xZPX31w9q/DZCUG8aZWSUDLOrnSTUXtmB
BC9VzsQ3ZibRH975Q0xFMZtVS1YKOpQaiCPEm0KeIgFP+Yr61hcP6qMxLkvHZNjs
tJ6jjtEMRVodGnulRLFsDGaaSvaVLXZVVxhO0hEw4V9grWKdvbbRL3/53+PfvNHe
twR0ELbVnZ8Nq4B1lFWJlVRhBti6CNH0A/MLeXyM7EpUBQthGZb0njh+uZizRyXW
GqALNKmUxXMRQKdNodcblfBmCb/kppTqJPwH2Mk++ykYAQjso/0cjtW8IU+OTEJd
ikcg6zFQhj5odB6c2FFaX1cwJfgqJxDWAS5iIGU1HWHIaKexU/a3zeod1OykC1ps
Yuts0M8Sb3rBQUpdzV0DaUQtx3wGfyQrhSCprG+xZDR4jHrXf+wfur8cp6d+SMnv
Pw45vrYGPk+JyuBlXIAwLdeHNoDKDHbBBDh/Qt5AfBVSRP2/LueCui9mOYUtNPmb
J1XUiS2cjX1wtiuYZt7PU/oeh3xzZtJeN+KNxOxMtZMlnaZKVPKhSnf9i/OJI4dn
Fmf8PY1/G+FV6Lr9b9cWjxzELRE2XigtqedFhiU+fkgUmxUV5kmUKbwDVAb9yaMQ
25k4UTW5BIypvAGmrGZE5TJX53PzP9dhOrClPIeGRXKqfxCCHk1t7R473zluUMKG
6VqBjwGUnOsYCxL/QOHbT0anSUZcdM/A8f7PSfiRFbWNMean3v6jCKKCa/esMGo8
PbCsmedJAvTLDKZ2Vdk2tAMO52bD1ExBVCu4liJoYKBmzFi2a65bQiN7wd3DZfgV
Viar0swBgPF+aMzVOTjwRp1mN5AIZJEKfJq+8CEQ7jOdIjTO3MqgnB35W7eyi6FL
gGCT32bTGwXS/zP/L9iA3IrOojSblPsKDD4617Fsb7yD1J86c6GKFwLoEQNKWSbR
X5ZwwrlF8qu2tcDXuIaYI6X3tbsoXmfpMj5GZUj4qIZjs8sleMmayz4nlTEIvnSE
Dcn4vGW6P6FbzTdWKvCEW8llYKM+KR7806Eet3rtOOsmBgkthtYjKRrWDoVVWxTA
uyQZRSg4//Dy5knMXd8gHQNeC1LceNSVj8sq/F/UB08lhSSK13L4F5YUOYXyUv1Q
l1EYF79xb4ejKRnuc+DQmV/qlY5DEaoX2kYbMpiFT+ViuGzC8iCb0Qoh6/g29qwL
MxQpmF3Wj0FvPn/eidE8Rj1KHZ7W1VKsJK08FHGQiiirdkcXj+DnAENkpuGVRNM+
EvE0HS9Puj/1vevBg/xM2t6zNjQ82BLi4oPvTJ/Vz1aOc1H8ATVIDIi/32ImN6uJ
+wokeiAHy7KY1scps76/L5I3nW+dka5uy2F8yNE5hLCGxmSIXU8P804lqRIwvkQI
+W0PjnUXxLyfrecp+TLtdUZlnFLWQBnn9FiaBLqMnrh433GSk7vCtAxndQ4N3o3u
E5+DUUrsSIKhA7JQNpAc9Y22eNceD2y2hp6YVoZiw1zlkGrD+kmniUlzgCUbSQ+G
rVgOkI91Dihj1viNcv96IcvP1xzvzR4J12E1cglUUQMoQ2R74R5KL2z8RwzveFPH
gSPTvxaUfg41Poq5dvw20iflFBXBJg6tXpnp1cUILU9Bkw6Rk8ehplJRAQX5CNWQ
N1VdI24YzA/51jjxL+eztOJf3xO+smGBJAZ8HMTHA9jzjymzZnfXyF8La4cEmaA8
dhP48gUHOLYzzjABzgCh8MIhfy9Gs05+Fa6eWfBffnakdaEWkKplFjiFuVHxK6JE
Dq7sToAfoB8MYA4bUjg6sbryBGQ58OFiK9bedbWylrEezBcn6FfOV/kJE6sF4PB8
vgCcPdWPB0/piwSo1rHNuYGQHQig5sxSRnVNxgXHNx0+qJfuREn7AGixs4km/ttv
kUXPBNgG17uuvrMcg4QoK8S9Otk6E7g2+yp7t0OcZK+L2C0yBK5XlslYeqIwBtYw
4wb1LY5ybYuwMRDDORuiJ45RhyWp1Zio6E9L1UkpAn8QUaADP87f4vCnkIaOxAmd
5oPLUVOctXPGCzSxYum/SEvt+LtIzhqlWqJL39yN1RwYAtz7b+eSrvoi3pYm6+5A
T9jU2GXC6ArCmLwpmD6OnlkNYPLgDFpkZLNExYnscssbL65G5xkgoDXEjDqTEyez
l+Gb/1j+c0kW4jb9OBQWeVdHtL/QrpEcIUleC90V5HiV+lOQlfwU0rp44yTAvV45
pAbg7G4fV5E6JdiyaP2kQOP3RYSsb3FrJQV3aYwQRxTfe9mH3KB8VmrM1TGiYYPB
yJU3XfKm5qi1KsNp3RhYGTXzT2m8fTUoBiF+FxAcRJs7bQFMu8gPU+ls6T7TUUQi
maO+q2EvNZuKwKB3G/sthbP//BQPqkHn/jzeop2EmMHKXmRQrVUXR9Dg9ViPWOVn
3GtE/3ekGLITgCwqpK34HGM+vZZs5A5nSIJKRn0kM9DQVatQI/ho8sPYVxXrqVU8
wel+J1wPVTDDPo68aWO9TciJpD3LSXUjTbu6pMaqbt/O6YNOMUOA+OUZElod4B44
Zpmd2gsJjgUfay9KG9ko3rPHbr8hDb0sDgzNOJrfZqJS8ZhKBmoTDtqMa5W+W0fj
GYQaDQOzCgwW9imzL5Bap/CP8k9Gjtz/fh1UVOzlMQ9pW5+Ij3rOUnpF+REuqpOU
Kc8xeRG+0hwYNYigzPRE7Hv6Pg8Sn9Ab8KVREDWcWBOG7hA+fM+rGHVC+BLmm/Rj
1Io5s3N1o0XFpG17xIv1tOpOQdhYFRb1VyMP0zVuMAdeM7pAe8xirhWi/ZHokY8b
M/dT9atoJu1hrGGscBI4SvtkDm3LTcJPFTR6j5Fz6hRWf6tnu5dnUBXKfUYNfFI4
9KHA5Gt0Uqoz0anVqJ/0FStYTSczB115T1Bmcnczko/zkARK1PwbbwPEHcklMbmx
/PI58oIitXLBDO5f2bnf4AvFDCtEkJXEDO3sKm76TVSfbBOhih+yjbpIVDGhGDw3
YeWAz9iy8hM2lXYzU0igEbiav3Z+w0MkgS8lK2ELQw7eBl8i38Od2mU+Grx+M70C
vIov3Die0zxTpPgPjVgrFqloZkxQKu19Vu+nuSdFOZhM6v3pjhXVsJLdtlXJiJjy
N/zLouLYYSu2LqVOC/Hc8hd0NnZ8CGfk/qSX9U6EYulpEIU2cqSdwI968EfRnWba
/1QIP4fGrRo0wyBJFG0gcdNOCL/I4wBhMhvOTE7ljGAPXX1p05WEzal0NlwxhAOF
J3grgnriGHPusKE1aMORuElR6mfRdPQ6GDRy7oXMi0b/BHDoKVK75+JUMcvx92/s
Bhe/Nf4jddNPQkmjwrmwPilaJk3rttpkkEFckaZRfTkxFiDhRAHhK/DyDho5Ags5
dck69uiuoYvnioqzbzk7vCf1Yp5NMYEaAqmBPOtMk0HMtucl9AOW6cUeRettr++9
HEAo+ow9yKi1PRkGgbAvvhsH2qE2W0HrnUFOQs0RBGG61ZgxnP4uKnmdxBhpFy4y
3qso22bMQUWp37AJCkKJbP4scG4wu7BoEVh7COWk/WBk9KYl3sZT6wSo5mPTbU9B
JJWUWYDxnvJVeoBm3v9daHwYcjeXRyYh02u6jHLM4Jx2cS+9mjVoOg3PAbxgpF0J
DQJ0ldMKNw+RCpmekkTK1CQlKoMInoGkgo1aT/zNAeAw9oNPGAS/Qm/pnJ4uCold
Oy/UK7Yi622GJojhbZCd23u98tCEYkLFQH8YarLo+zAv34S/s6oGoZjv/jJ8sPfL
1IVzzZLUlxTJ4v/H7fiZ+46Gm40hpiXGZyJtt0YjkqCBQrGlnu3xEfNv+I9KDE78
/P4wpMyp1r756h2EPohzgVcPqfUaU8RZ7kMcDipV3DjyRUiNqQrus/wlyzYecotB
ixHgezP3iAtsUs8mj27ZTl7wNSS5rmPDDRTvGDc+660eUw2EIqRg3n88JJwSoz3A
0mrJdV1hBilRYDAsMLVBZFJWFFfpxC7fcm/4UZ5Ma0YmMYxrDU/HYHSsVSqGLO1M
slSdShMuN/WZr0iRzJLEg7d1J6VZVzUjQ3qzWpCLAvODcU5l8412azpMMP7QMgoM
jsvRFPENE6RlhuYTh/k/pBVBnWw4+CrtrDzE4BeE2wypQ1DdJaDZ+xajvUACMILR
0qwi52F+TRU5qRtF4vKrulttbf4vQEjXtLBpde1Gs+0owARdq8rvdh1L7jTdScS0
qoUuXEtdgiSGBB/5RxvbFM685ojH+yGAy3cNhlweKcSFb9OCO9ELJYD6z4ACptc6
+1iDJb5dPjeuebWw97URpLQVYzu2MdvF3PNpdFOe3EiLzuAh09pltobllmRLxZrM
es8yaZ9bn1jAXgILOiA9UbRxqKkUfvXLLAdV6kWcI2rA1/BpThzwQZML5EK0YuyF
Gp9eQECK0uxycp1C6itc8VifP13oSE2lSPYCDdBtCzfaoQI4jifbhJ8lDkfXEl3a
usFucDlBXsdBaM/oqdMaBmU8B5frYvYsJuU7nKFOsY0haIMcu+I+AOeiD+1BWEJd
6fCkYHhq5iZXfg0BB4/MD2T/1OKiLk3CKqwHOVE5H9ZOj5HeS/GYFcZOn+lSQ5U9
ZijCB6U74HOMD9y4zOMDhyPQX3ZWShT+Ez8d0IVDikk9673ERW2kMtX4XNQQNe/r
ilDiqjqylTgac+e0YhGVAmZHYtqnSV+VkDjo3rnK6TvqMTErtKloW4QbMvt7B/TS
kNOjUr9G3yTi/2CY656q50K9H5mJSg12bs5EIa+GwKXQMzg8WROmWmLuF1jTIjDV
zHILLNnI3bFvLClTHD3ZTurrsimKJT8Ryyv7W7i7fqGCL8lHikkwK8hWAj4Do3DI
/sRI6MrNvaV8+iZ5nAUjB7tMSZmKtj9U0K8qXDZbh2uM2lIxqhsdDK2AM8IF35f1
UlRH4gA8owy8p74bGJHZwQCB1qjgMDKjhKtLcMHsvq/MgdL/LpQxi+QPcfbKNvHA
HO0uwW+tzU1FeT5pXcJcZGt3ktUzjOshkHUlH4L1jZl3vIdR/hkjjFXWCLlIZCdJ
usR2yDpaBp2d3xERwajWHZQC/HzHql3jE+lKBJh0ULA1rmd8fliORC/D8mRZCWvl
8O9F41yoxQBS5parcdJXnzedylAAv8ETvHCspzJ6gsZ3jZa2DFV0Y1c/N3rFkAiA
vpc4F2pgDhOqmUGE9kwwkS2ovqQ/jKzUu4G4swH8sKZsFHU5qEhUMLKZtwlGO641
7EB420rioy9CWYlxQ4gXr4H+yJZgB3nlSXQsCQx5xu16UXE5Ov5k4hqzAjX5THAn
q0I5eBHn9fxeM8ED5HyGRxvj1OG1Z4lfyBL/rVO8SHiYBnOupZJoRn0aFuCTpuip
G+VeHM/qz9yo9X+R9wDld6iPgYmkdITmePhp8Kewgl2b3pPd4I/E5RxXf7Y/3nb8
nNwRGR+dK4unaXOt0W/dfTho48Ui1cD9KlvViCZR+SKiRdqXwjWbsXQkyiJ9Cgpt
2IqArFajVDgVJ3uyW+JWQ8WVDLM5apoFUAorvf6ImHOAL6y2mmNCGW1MJKmihfhr
T7NXp9R3BsO28VpGphBZak2XMCmZ2/+wn5FBzxwPQU8P6MRjBcERSv8QCNkIIL/1
zy/kVlprOYncDrVi5zfnH74JRL1r2Mm/BmUvL57ih8W9Og1HRHOTBfkHFMuCRh+N
pWsZkR8MBKif03Uz/oh/uROCc/raPxTA4eBeJyq1jqrYYjJXSOlDFfEyzqerFH7a
E4n8ZBSGjP5PhgsPnITNieE5w/LDNeDLL3zJ2ujpbT9Lq4sc7FCdTL1U7pTGcsfm
7WINgJZ98bf6r4g4OC3pQ9kctX4t/tKkci9su6uXykf92HVtSCsEJgtG1FdZcP3t
3Q1MEU6BvyG8nllW8d8V92/Jdw3adx6d1UBY5DgHwJJWoH2v3aGpzoUlnC7DKnLN
DWJZ/5t+ZG+G17SEF4aQKT+mtrbK8ul4Gho3IirbIGB5+VtZerpSXK9FQpmzWm4m
cOIVEBqWgpEsA2iELM4TAKRhNJnvaqxU6SRxiByxgCF0kYZwaRfEuCTjYN1BDu9l
NClj6sOorBvZfBZO2GaS3r9QdsUaRXvVD89SJMg+MkJvHY6smc6prpzDpyMVesj4
Qi59L3GgDijhgUBZJBitgvNz1/I+xVzG5+Wy9keXTEyJGA1hXp1eVzwz2ie+HWVY
b6yPPOHEQ7QcRSMqlr4wH6sOtq6wBiSgH+biP95CWSz3Is6HfwcoFOFaAOjp44nv
CSFQ186GEHRPHSRwXVJwLe4rzpBsAxab0Jb7iyiI94jEazD3rxyXraYlNUnnnvKn
FE2puYxLXnshg0+1HVXGnzXAETcPlexWe1x7e2FQLqrfFZDap6E1POPSJmtlas6+
K+DNzj+yUh8hGVkV5XzRfVcsjl4anT+U4CHTDDX+ZMp6D2x18gYGpaxj0dPxnRtl
N1NZ1UrYLSnTdONimqbXYV1pgxa1Jtd3+e/Za8xOudH9AH+skOrWj47Wsp36Pwrh
6q78v0T43PM8/9yr3PhUfbpi+3Hruz883VG8RTTlGkndrUnn0vX7DnWQdcqMUMqh
giR6fo5DDod1dbrlWyk5sbQgyFcaiUv29KeYRftsLkPtvKkr8jIOGIsLlgDAgLf4
erXZIU+oR+TpquMh96WS3IZDB8WGjh2r8ptMLW6CQFuoc8x1D0YuSSpSLjqhtTrz
7KFMpoTc5QHpnfEmbnUDSv7bBjN5Jve8L9v+diPlfYczaiz4gkbfcSXGuQDh0cmN
SkHevFn/H82U3sPaXdiX7HC11T4+0kU+D6uQhs2NF3K7X+SFncxn8tcyBWLwlfcr
oSQBpQ7VJWC4Oy7qqpurbEn5cVn7ix0CcpjkTtdhKK2BdeUmhiVQI436xKuz8kw7
qbt3HGb0RCXBFQjfaFRvaGEcOhjsWgkJlgOfXx7zV708r0XVpWcGTrafztOdEQsP
JciC31vgJxLm/f7i+riF0fmai9aKBGCKO5e7KqG0s5+VRJSjNceVJfOuu/R96t1a
aSzipS9yzkABnYXbAcqWj5KxmugHSIZWcrvZjfVvONtPjAn4qRgoznZcOoh+O/Ty
hNAX6NUWqNuy14mVDSXvEBjgVYangCwWNGovV+BkShBETbDSYYH0T+ZCTSp0RP8/
chiHkuvOD3X7YB0qQ6/AN94MvAkWSFPMdxse6P8eS6Yr650ieVP3Yg0GnaTB0R0a
YEpRreakmU4p5TVc66CZ2ZXKzQDizRfBKeHky5kHfVgbmdDeuvQmg7u65jlelV5A
yJw+0291y+0MBZ9MQxnhuS80ntiQPzvoUrCqtS+LXx0sDcio/DKh2TEQm8s9M+FP
8wI4tVK6RFDzoHnppV6FhrkuQ74B//ZdrO4jZGawFhLIOSfZjPirp3WwtBjTGzoz
7HHd2yUOlix803z1ijaZkHQzZoLdkBmXmKb+vYSoF+WcmtdSApquvUGuvdfluBOU
w25+5M7vrlyKChY2uo6EFNnLNKeqeu6at42X2WBjMzkXGM5SUYoDvpgJD9Ux9CaO
jWc0fA6fsTVeC1b3Bcg11ZmgY8p0c7pv3duR1ycZwt5tVjye0N4F68AB9W81s4dJ
DoHJUCfPOjycm1PPi/+OtnBYHTLj3JrVbwu/IxWag9OXV864mH8SDyRKEJfSNXKe
TBxXmtqLv/Spkvino0yO0taOQ2JZGjWgjTaRYLEgN4aWZx4Qvy5x+KOM99WzKx5o
YmPL0+9QqXqkc3HZIqEJH6FQcMhycZfS/SxMzA7ApKQRVU0jtfWdcbDoI84GeQov
fHqTDTsjlPw6KeR2a8vc/+RKHEU7aXmELxY61wvQZjfmMlW4eb3gKfXuLq8kqDUq
CbSzrZZckUABnZswskPKa0ocox5h/OIsh25g1knKMChak1vWuYE7/MpulqBZBpDf
nvXHc604R4NHxNWLdKesZ/xIHcrDF66As4RZiKtaa5fN4U4xrOjnl1Jbh+aJrM4N
5pYXdYtm/CtBmEICGzpq2eDWJULlx0dT/bQGi/JU9Kar0E1DJowHxmK3Vy5Acvdy
/WmhsOxul0X3wzaICjEr4M4+wffItpAETHKTpLkGfx+y1cbxWcNEN8mM17e/7QUB
QkGdXR1/3e/tkaZwY3+IM4tC6uu11qg4IYAt3EJnI3bl2frM+m66YirEknB8qCxJ
uVQcTnCjytIvRr7PPznBx51a+gC12B+w1ac1YM3wWJ6M4dTXwOiDKLooWOGkLLVn
jkPvtpqlFMBAt4LWmi9B/HQ/UZ3e50v71p8NRwyiZz/m5mm9JkP1Kq9p5YMdJ0XM
eHehWzSE/1wwcivAcFsw+3BBBagHGHvFP3CaAWk1qDL8Cjm9y6+L56sUsfx6L0Hv
jCPpeV3banRss7ZMj8PFINkl5Wd1vlsW1ZZjVpyj6UfVoz3DV2PKILEoB8Le3CmU
PdRoXON2frKUjZU0O+/82oz+pHFE9maocV/T2IlQTq8GQP0VDS1wiXKczk3QI9C8
uq8mz3ScxN6eIUmzHXd/nBsa5D1m+JNzkR5Q3SsGqRCABj0D2UW2kM+WIfOJyCfO
nWH/5FjAaTtwlw9OYmjHsLEVoOnnbYTm3H7m0Q561vZG/hYKeDHxd2gq/Q+8INIM
2n/guRSQB6U2BzLtdpK/PPPJwaRZV1VTXjYeGpDvtpRUe1NR8aacfgLdBhpvzBAB
JSo4KWJ48Oubt2Ogg+9Z6s+5OGYK61RauxJSbDduUsQrzA3ehtEysiscwyjb7AJu
uRHHw7eWypDa1rTtbbxjCyGf6djcMfAEsLLRg/71IKvwTEyFE49ic5Gd6Wah0Cxe
WygF9mPh3dKRnkwVNSCgcdJf2AgJQe05wb4Z87D34ZAPuFc0MvV133tXVRkLwSH/
LCfETauMHQ+GEmpAOQk5qqxVXybCgj04lwDpnEh7/TOosIMPFyqL7tgtlFKPUNpi
zynkvjiBRvzqvEW4wdRPHzJD7tsVmlKgZAgCpZKFLtXq/XTfFkX+Vd/LMx0icQai
rwV1EV4siJQq0xNuOLhGDJlV0F5Kg/6A6lTkOouyJhZ+e/XHL9+FXrDX2RXq4wf1
Ot3nqN5avIhcxFvLeAXJl04eqYHZm9vf6U7ExiR3d9KmUdiP9+FdK2IWperdaH+2
bfco3wIcPTjsOGVNfaCzU3oaAjLSsnWpqfG5RTIPIZMgLq1Zn6xtIgMjhuXwaR0T
ex+rbVRoLtoCv20Y+KQMewl89Ameo86aiNtzOvgFqGQ2Gv9GI6xu5Q45/VbwsqwA
S7z54Uv8H0/4G3UwNmYNuSIQethyftfIXEMrMJbRp385yRm5EnAa9N/dqUr0/0Ro
/pxd6YwkFk+2xs5bSn2Kb3y/FKszYKZoxBqidBKmyAHQGK2WlyxsNRIrHUIq2V32
F/JhsCLCWXIDOJgg3bHIN36VLX5cwMzSvRojO2oYcPdwIrDcYyz37YtnJ+AawwTY
Z641ReJuSGs1PEL0xr1E6O4XQOqf1ycYxnmFkjSvA8uh4Cot6Pb52ywwVfR3eAVB
ubZWCTbZkkBIpKoI41Zv4H7O9el0j00e0Pf+GgksWLuFAAwGxcgGZ2cGzuaD4wmH
+4llf6gBstcme8gxJCJWPpLv3b/6T4vNe4HR3090BL7v2l324V3wqTAntM0u8sCh
dwDgtLQ3EJQMQkQM9najVGoz8af95a06OmiMewxvYTttKtBKKQxpZrlTUIqQtXlX
jlgd1y4ICCFMcYaxqPYyf0kafaNTrUFg9qWnPfSj9dgFtbdO2vzJ2oNIrMgHzPY1
QkOQUTgwmR2Qr7cnSdbFS/yfubIitmzCifUKHAJLPRSg7Fd/DTXxpsEk+eF2EIck
p0jXb8+/dxvP3Mg/tiNe97rjbHuGV/uQY7Xxi1CZiaO5q5wI9dNQ6GA3fI1iplSk
T7iJU/b3OYhqY54Nq5CplN8nVrSdj3gLjCY5E2llcl24Ysz/424mYlRcsWb8NhiD
Le4wUqHPNrWkIYFzztfcr7+qF1VRpBO9sOyhBWNXkOFAlN/hn7LNA4NG5NwjcN7Q
K6CLIZCsuiyJXww4gn8gDp53DOKpYPGDHUW55IQ74SoWOtyCrAtrbNFFgPP2SujX
SVAUu7YsQSDLO8g3goa6nAF664UehsyxUBhAwAyseifRz2x2h0pqbF+c/aPDLSlB
KOxivfOImGbHr6wpNXmiyedjF3jjVtom2mdxONDPMVOCv/OeyBLUu1ZcmOJGnwmx
0FcXWwMBdRh9A2ielmJuw5VqLgiOdCWX6nJHGiPO5qHUXO1lgdqQ3CiuogLMi4aR
uGWwgZH3TQyhQWcrg/iV5nau9/ImVFAw7XMVmIn294xWr6pale+FKW3v0uF3F1I3
fysicvY4wm7lEcXWO7IVx4IOKBJx7BWuev8yJXPkyMCoJ5tvrMTcxmEr6xqC20x0
ASf4OLdlv23moyZyxFrAuGwLCOlO6irjcunAgWqJmU7XEc4T6S8db2TzwtW3FBvn
DwC/BNezi4jZyK5o+FWUIR91S2CYRKfIkDooYNasq8IDpLn8BianBSr62oodwZrM
IE5+bVFUSc19jRjv0umGT1yvll2NmTYXYGVas97rNDm/5g8p6QZxFL0SKlp7+Tn6
mbq5LL3R8ABbbR490xEIw4yT3DZbSNYQ0JgPp85RRHMr7d9BhtQZqPh3qpkrGaY8
DIGd5kAyUCN6pTu9yHn4jhAaU25QKJj4KrlBq65YeAR0SJkEMemz3uostrMXBpUo
5o4Er/JH5/AF41gd1Q4nNdAcFO5uaCXvAkjtcDIZZe/YhwX78hX/X+0J8qU2IdJ9
gkVZpz9R2N7QZR5GPcRvxngCXawN9JfRkviSCKW7iTLKtGK5akP7UL+H9ivd+rvS
YnCXO8m4hF+5Y2U4bieXVrqrLI59zRVRJiTeHryXbcBbC/kD5WjoewUcXhOsZnRR
zakmFIvW3CkKQ4vqkuY92htKs1iEMITaJlHRkFUo7FL1QoiiEObaOkKyaGSe73Io
6LysHgP67lZA0w0lLzxQrYX1nPjVbMKQlznWr1JkABrSzrjITcwBWtE4JHTBqO6Q
SAoyONYzsiQyXNOioP0enCrPuLTvnOjOltuz0zXh+x+FjcMOGGGnvMX5zKDDewsj
V0p9w6nCt2AnF0x2liDQOd8B8hodujecp/8K3y+BN8rKT7A34bz8Vvc9yrvaLj4G
/+Btu52hlHHUkiKLw/aIdBBWZkRDUDdchDBx5vWv2gFcNhqu2syjedgwnzi4hYdh
ygFdK4hHIa75ix1khtkwVLsIiKxKZdfrBSb07ZBIvkWSRTNz3G1lvUuNValutKWl
BHlZQ7FeTEtK+1g0RXl8yEk9WnR4d6vAfgl4YDRmyDbxcZ5VxyNniC0TbIuMoXR8
DJv8gvbZWD+wpn9+wMXvFRJUZxbVCLW8+q8VxD2tFIZ7/GZT8V0KoDH1UU3QtA4i
pooIwP6ESmB3/FfmKxQmeAbIITJ4c3zhgCETz7QWN+GQdwJg1nhEc9rjjv5qpESv
4rFTbYQw4mKl6nQqlWl944pyKOWQAFuKTgIqoGEBlUq7uGDumasjIQQqzrM4hW8R
/UsOFZ9NoKlD76w/CE9aKM5EgZFxsKmS06kHJqKr+sEPdrQAdyfcLOHpSp0hsybD
JEVZYjuCgD7UrY09KGwNnlAxbGxEEH7T4HmUbeVs4pM2WNSKx7fB2hz+Oxpa1lOS
skszEcbFiT4KPaFSv5oXcxuZgbAhAlp8FULD3EE/Hxv7axO+rOT28PkPxYW3ORd7
MLiepf+22Ps5Se84fEHyNct8tSxA7p3TLCCPq5rmdu0RI9cMKW85TF1Yi/FNgKIG
biK34Bpdr6h9NJSPTj7yfPu1HjEjEktLooePS/9CT6ODXD/2lZZq9SorbeiAhRJr
f8e7v00Z3rhSeWIpGici6jWhIPtbnnU0i1xdmiwMwtCmP6Shwm1KIiAKxFgtzBRq
IdbYDohpnQcVuEGm84SEQnACU7OGPdW8JI6T1cV+FEJhRr4ga4HyhJ1C+1KsBPtu
p4eo/35nv8ukcsBy7fGylUzb/UqY3pMK6f9CHwSDfOWQ2ISJ85cO7qei1tmnd4HS
`protect END_PROTECTED
