`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQPcNfqq/edqop29RgZxBu/Wj7/6OqbjinEUSutp0aGRDlX2Iwrz6zemLZ6K8rDZ
k9xphGkGIKB7XtPwyrJ6SGz0e0OfnaJ7omyGHxc2X4Rlo/io+qe34E2Zb/tg2yxA
1IIDq3I7IxE3xC6Fecx3S37Mcb16+hphgwOe5Z9aBqLAlPh+8n7L0gh3bgBX60zn
4ggKYMeebJm4yTu4oGazmsTOINq97Epue8e3iSVlcY2WOgqgxfzneAW5sppoBHpS
eFJynulePenij6sNENsa8Qg7FxptPZSsyLacrh1+ns77k8SnWttwLR6tt4wV6aWo
wXCTjuHpxGt4cZI5a7B/TY74YstSKI/p+H+XJnUIjDH7aidlwSQDnt2ZKldGiq1d
Tj2HVm1IwLHbMspEEE/1RkfHaa60aSgaPlje2/L8WOQQWz6DZ2nBwLkR6YFy4AMy
Fdyq1Tk+ZV5yx02x5bjLkokWjkpGSHtsAGVojyPt8Qcn6kw910DDIWthyzpUsVTU
KrLdUj3X2RjTJ00L0IbqAgDyhq7alGe4/g2aLFIVkYUYjADHFer5oj4unBOsM9ED
kmVV2jhlb/SsPyJkWDvlD0t8i9+4bd65I3ONIoYgXDfTidZEBxBeRpJF1N6H8UqA
iLuR4O75deFC/UJZx7O0W2uL93Rq6zDAC3b89EXtlsQVxbXcgEfXtmVDZVlp0CEC
8ORvyFCQ/XGPxxIYdeblYY1CHpBMsHxEtH8vJuhl9yv+7Kj450XtcgrTIm1rxl9u
F7EXPkaT6Ixm2QAKcxVh6hUgHcG7Yq85h+9J3jTLmvlEbDH452ChsIMFQxdyf9bW
JIHCJY7rO1ETSR8O9KNrYgfxr+YmnyqDZqZGjtyNDA9iiOfX4n8GfG6WjXIsa8V0
MHK6QqwYuMV41wnIsfuMZskorqDxK2I177d58NaT4JLdUuEcWfKE5+Z34Hf9O01Z
CNQR1aMABuahgtljc2JVj+nw4UIH0fhsAA0WLuo48v/cwE/XVevJk7k1Fzki3aZI
`protect END_PROTECTED
