`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9c7STdSnhmfZ5b8/+YtcsbenVoLT4h2hh+6k+NglD51nVTJRj7NlNdY/4PB9wOFa
kTrJeOZ5bQgZ3qaFsES6aMdJacPhIDLBYrY1ggxkiD3Rplh6Fm/PxiprYObCF25M
c9ccIR2eF7arGVhqAVOJDJpqhl98tOPTQ66Y20U+LmKS150VDApSJuBKYN8LQQii
GpiM8eng7ZgvHDekBLS3gHdPRJcGBkHCj76iEgpoB1wLj5iVX9GQjE94+JQ50uz/
VzNatArYKNbpmX/ShmhxfuD/UPcTPUF+kFrzUO1cyxtsv31NdgMi8nU0YFaRC2zQ
v+YF2LlWBK0/9TgzqP91mUr5dbBAFzULkk0VbzJStcaavZa/2Bkuz8uY1x//Sqgc
Iiuko4GoGDNR1nVWlXmoElCFQd51lP5Q4DnFeBI//qA/+cwsZtI/h/AHRQm5JVZn
ceYxCKDld9d08iFzgD8vVS+eTiSdWjWgcPgSMCPPtDin72O90Mu1pyAsX52D7Rb7
eUjNVwX/gQwBCPIMhOWao41qJkulNQda3uq+lP/TD6VRbFku3eKwSWxN8qbXPBGB
lbgjYTBI07WJS1hOzggmoMxaFQB2kBdiMtgZ6peawyYOF4e5y0QQYbZ/IsKu4461
IC+2ObdtVzu7SVdKY4l4x7805bw8BVTQp9SwyheNe+6cfkk1fDhwkKD7rVR5dKTW
WS39n2LJujwfyRnbP2r3sxIFdgxZ3Di70pFYSn/QibXjsxZJPwzj1r3OQdlxl0ye
r598HB/zEjIH0/zVzSTF+dtzA8Sn5oRi6ZFL7MyUOsZqvi/cq1ldtMdCvhM5Osjg
bYLrALFGvyGMz+ghOj1VDl75iPXdUJfpYvoqzgn394iw+BelWmyfzHpLRdiwkNIU
fmqo/zORvYdleA2vB03sCwoaa7jFdOP+a06bHG2nb2LwWpOoAKjZ38mK7jF66CTF
9W7afmsD3fThy52kG68bL3C/7UCk120owGIYG5kjVXDZkt1jtDWfyMDyBpHTCLar
efGATQNi+4HHJlv7Szf4xch1L1FGc6zZHkNwOtvP9Au2Xabl302hD4PuokzFsTyv
tt7ZM3yTzKQCRUnUYl7ljOXoI4t7OnJcLAT/jVwV+DCivN3YE9/jODYMIxsLs/DI
Bc0ya99Zx6FA9drCJjsC8fToL6y6C8WrTkumczB9SgTFeID2Tq7iH9+khdVsB7X5
RJGQ7PQ+8NXq0NZtNy68k3e0nK3qZgCzunr/M6TZGYkfUlvQBBuHikzI9TVLJww0
HVIih0HfPy9W+s6a/YNWvwUiBGGhEvWBOVobJXf/1gD2xTGneE3UUhZVhxp5uff0
E/SFDJ6sBZCsSXUFBfDkVZD+GJj/aWzc5SM2kGue6x9yOKP3zEyuoqO8EQ/OICYu
QN9K5yRvxhTz/pmkdbDlQxUbWd/+UZPPm54OZ2jTp5svkKzU6vv112neSSJZl0S+
t0zFm0+x264jVo1xmJpHEMgFeA3Etzr6jAHnouXnZZ/q3NCwe6m9W42HaY/4tpJw
NGRGx7E4k7ZqGvyql+AE7X2KbhfxL9U6WlD5S+ZLgn1P9WBTdtsc9FbdTEyuSuXW
mcU+/SG/34goQo1SwWuGnDHX3SxBf+ByL4jH0VG1KtKdks19JCvH7ul6YKNsrZdS
hHkoK0rKPjfQmSDRprEpWxCdILvNrvtBq8P4+BfOsenbTr9VxFwkTdv6mHDU/pKZ
86S7T1GseNg4HuxXmLObJUFS2U2T60iwAR+b0mQYR3isTVM0beevrimcF/ZGA0X3
KtnOxoP+FBq7MKJ1S0Y1YojenAackmZC3/07EDCjnDOPL8gFbHEHkdExWiZ/MT5o
xMbj7UnvzhB9vbAQ0u6A4Q0qyo7bH8pPbSlxdRXUIOq85DUWE4EFYahD9iem6NPq
zl2ndfd+pq56tlMna6ysXQwAxUpKfT+nu3MqHJ4RZWDvGjJIc9NZDiuhAi49K52l
+h6ReS4hi+EIoxrpkZqCA3f7foueSUK9cAyo+MxzHxF+zGvRI4qVWLJtbLaFn6CO
TIizRYDYiIOsP10YrJbtPEGFlMZlyUZSmxdcN8QnaLXpffKuAIc2oz2UFgrgjyW+
qnG6Se/4s2DFoo4fjKpTjbnZ/S+ojpLb2hl6PTTzdvP1VVHo9nn+tK2efmrzMiES
dKrbGAM4D77NJyrnEZvXVOSslMBbnnNImrTDdo7UcJtEc7pToKZ7g2mM+YFj5xor
lvlYXjVYJENf77ENRP9TQaLJfU0dafKAV0YTw/GZrjkq+hcztKKdkMEuASkrJEei
+8CT0uUmpABbxmKiEBbiftnml9aMRkVxwR4SgRz7uCPd44JoRkQLdzaeo/9XGQVo
UwEn3gvKTE8Xgw2cEIdOrtsVq9yxYHaM2NzYWHOHo1UjJ7MicJsnkU+Wzzmt9xNm
vT5QfR2JRJDB3l5bbhxGp32D81mWEHod2hlWx1AW5Ha3mJsnjrFCh7zgBf8hUR6q
loHpvNN6j/sesL0MtXmMLrS0uFrznzyVzMTHy19GRGZN63x58yRTyL1kYKHwu8JF
skB4EBoKS4qYOEUcHfkVN+5DiJ73J6+vO8MzFjGA28xrCB0juRjfWZRBYDquWDTn
ooLynUSqfCMb3OSr3cYt1Yb0wmItMEPInx2SuW/QvrTl3sbEaqt/fA2VLfnZtjz6
tvNMadgz3gBbnBahbLaXl14pby0QD7W8u8Fo7SsO4YICheNYec1MDSa3Ervqbaia
PY8udIoI0gMTZktH/iXus1ymu0U4UnLIZHYKZvMuZ5XPxzLM08XO8K5J2pxJ6XVZ
vLJhy70R6Uhj28W33YqF82ZsLELk4J/vwoegFfntu2MusbJaZ/XGAkzamcVA1C/f
83XNW2Y48/IvE2tQo+DTVJYcKFWRcVS5hi+1ooXQMMURQDEaCkQnYZj8vhh2qghK
KrZwpaZzpnUgsyhDxjJrvFYCRtRv9y523oKaKwMKVpDmaVcKWlrDqBdowuYZgRC4
evquvoMNlFF8LCTyzJC9wCOlv7z5VJMYEH5zlK+uaXOT7q0IJe8DzI9ATfgkJcAh
ZbcNlxhe2PeX3usAXI3qki8IcWnONMCOd8+tsh5s3SIaZs8zUlscIf5xlCFPXRUS
+Vg+Uh+IpRhXqhTeLoMDQI5ATSWstEBpFsqj4XIzoRSFXzO7sO6zreTGQXNeP8aM
l49Ma7AYHTrDEMiCUrTkZLGNCuAiGWrJr1sIh0V8cEUTMy+vwDLTsn8ZFbgvqooM
kp1G+3ZN3OiZX9WG7/EgjdzgRCeefY2kOdXgvN6kB7BEqN5DTKY94WqKwU8eGZsz
RTxs4buBSI1b4F2ge9fJeG7yl8ZuGvk3ahlKFojdig1WEOo66Sbp7dYyl14I4Cqi
QEmoA+cEoeiiNIboJbzdUM3X8NsNToCXAU3luwsSG13aCyTcOmugPVqDS1vD3E+S
ctf2zteeBEt5dBMcJEfdhsgpzF+d4wC9c7HwagzkujZ9mhXb83X1SZFkqZ6Wt0qM
lEVmHGoqpzGnNGDlBeGKsEen/dGhiHmtyHhdHxZoFfJlvcGkMP0u8glBQMOKj/AT
athW0b9I+nX0dVczfQ/NIEaXrTNemidgsligJYks6x9jiWxisQKwasTReqh2JY1y
DiGnQbTedAP1EqEucbM+ypzX6Rk8LmHKleObMYby+jFYuyKF17CydzS1XyU6D9Y4
KzqK0dTkeCgMKuhVxBAF1XJW/kUXIGK46bhmD/mXchvGVysbaUJhp4lHBC+x8CNn
RDFFaqsTVx+0qBPypdVNSxHI2ksqOIoJKXjtsUGKRbpiHAi+3OSm9YWWTmX/FjUC
`protect END_PROTECTED
