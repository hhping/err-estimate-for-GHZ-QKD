`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0pypS8wxZ5khBDeBM9hO0Vf1wjeQvZ+bC5MfKc+1oW24UxJ8IbfoBR1PH/GV4ni
IvybFHQRp8rSp3fx4wZXiBCYaKRc9UFS9SHAHLWtfQstPuMQfdoFqPudSbsh+5kB
E7xq+eRKMlqDLkcH//88eEjvp7+737u7cgufDR2ITWgCZ6mmGBQDbnI82BlvIaoj
WopGiLh2Osp9f/Stu4AITW+H+CKSJWyvuI0kMpczB+oAHXKJBT70AZQhY7IjBakE
BGIZxffM9xU4f8EHglKe7w7X5pcwLvW1XEds3coCit64vi1VQL67eLHhgamV9aIO
Od+hEFjfJSQcST7+AHl7jUlEuN9jfrJYao8YXGxtDehKeO+cHXDPhGOm+YyPMYiR
8EIChPTunvxeXw91DtbvkUSvrBmkIqoApdtninW64+7Isf04qphO+NMXrmJhZKzC
gFTjz2tiueqPI0xAixiitb6kUN3rgsxkR6YCnWUwhstDDfXB3rGbkmWCIqWnnqEK
CCEpqaOyTGdrsSYpXB+1vb0c4FQ+mQGNebftRzmhhiNnx3sJxdUdSACRlFnfJ41n
JYQm4X6Pm3A8vt0USOalvKADnMadONaEr3XJLeoZFVQd12kzD3ZUewQC9lszUEyw
oUKmWs6K0HJ5CBD/BWFZlLNw3d2CMs1S4b3ZrXe1ETbj5xqoz6Pn4nv7PAPrD5jB
n+wt3sz4e3xE8xkqDRV+2tdgRWpQyFK6ewXevFWBbeOJRuADFZ8ttMvNBFSkV6C3
nOchVVV6ps6jXQewx01ZPTddM2yP8/F/GSPPIzbcyD5ESd7GQzEB7l84MWPMZ0s1
`protect END_PROTECTED
