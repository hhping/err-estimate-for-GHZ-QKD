`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5YqIaJiV/5mB9c/cmph15S7zVGTNs0DXf8Ox4t+96WaGvixWQuI8GEHrvDBb4Qb
p0urUN6Uhw5fQWPdQXUU9BzJA2c4imbA6ncU3ybxJmb7jN+ja/BA+8NSjIVHazha
s+R0v4mRDh4ILTeEoSjqgFStcSsF4UXdERIBETFv+QLx/vBuZywV7eBvU2o/ZjeH
X7qoaAlH0UArqdm2ZX6TDFirnXV7the2PfwWujPYgLZ79hDYGJvpYwvqoAHMmwpo
bI2e3y4BHTWPoLkkN7hQh6eUKmQ1ZbWj6S8k4IYaXRB/yWKien56f+0Ckom7Y/3O
iAAOAr/4OegjIIzDvwE1e8PbKrPVSwRxR5AxxH0rgOo0Vfxg/ND1C6rT7duGyelB
h1Ze+zBe5APZvko0AUkHTX4SuBwEGmnq4D/4fLEQx94LzoMT888z1fcRqbNNLyLQ
ufmbi6jcSNeoMrw0lBPN64m/APfYL6FJex1zk9/qCmMpWLVIw90ogDRIDF4ZFk8y
54kja0kOg/4o3D/BEUlKit+QUGzmUgrD1EU0B6VLxHDgECPxbYeGlcOwAd90q8UC
Ycil08af90AIgscWU+T52ZnpLq055mA45Vr+quLOnXF62arpMBDNN4xmUoB7or/H
afh9xj7qKGZOOnR8o3mSwI7Y/fMqNgqh+7UiA4GBiRbXfLS+Zx/PPyWa85q2ZY4h
XPnLsiXOP4kkJ6+XU/hjLWhhQ3HORMH7pX++qnFzZAIHA9Ib0UEGZAU7Xd/gzMCL
WM+QEwxkSruSMTD/PXs2LM6+mkGvz16usuOVUNUUfpNUL7nqrQofNPRfajFT5NQR
UtxCzqnxQiXrL/bLA9MjOle2sAjl84pgHxIgX7S+D65w/nF7OVy2paYnI7KjU9JT
u5keAlvNhz9Acf3RYHQpO70h6XdFWPIKyTlAu1CCOIWjWlT+c0xxWubt/A6yZJgK
L289DBT584zS2Q8UqD54thXhjKmEeOfpfIrt8HSBN4NZmVoccMF523tZNRf+eQ0z
f/Dgm10Yj1D1/ZIjiGlsbxMzyyt4AKetfq4nJNsw1yscmyuCslbl1JPDL+VLL74q
wXA0K2W7CiuWe1dFqDAfRsLAMhOjbBvpM9+4BMpOhEFwhFMhBVA7o3gIpDRdVwrY
LsexgiWZAFmA5AZa/ZuGlu9XTnbiH6IQDuxww7w3T79vpdc+jePgKaFb0qTfspZU
1E/Pxy1ulytWVTzNqshygadcLxkx5QOk0rm7WlJPvu7Nl0pqcwR8KHY2TiEhwHFE
LLR9dMOu7OdmpSbFf6pe8zojUlcTajw5ac1WLjlKkRO1FPgWtOMrfV8Dl1LRkZ/7
ZPmuL1NxpR2T9wxDFmdYy43auceZYPVEmKrx7otJQn6SWBalmulVY6bw4x35DyA1
C08240VK9nsSGDHSVtpaj4xkyPghiVp2qTB6RQUwJLGHLFgo1fYL8S/w1s9cNUu4
WaI+np6XpBVVWn0XHTQOmFHmVCwpE1ydeyn1jWAPp7TSrOLiPpwEtplMM65hXCeH
eWR6iIk6ahX8pfivRagB+wE+dUAoJc5kGx7/4FzMTGJ+boHeahWmNxGh9AdebeoZ
jWoDvks4RAR1dci1MT02nbMyl/8e4u35sPxYWdgljvASYghM/0yF6+oK0Dj838ei
oEKUPiTM2XNOasgzcoLSABICu81iokuKe2JeQqExFYZmL9ogvtMk+vRg7r+VHbhO
Ye6eHNaye1Z78RYU75e30CrXLsWgcnIO6esXB84J9yonthaWxHvozRdVrf3TePS7
prZ9okro/V6v4M0KLjLEyvdw2LWcvnq1OPHEkL+KiaqCLk7eU6mrPNDYmM88dKq0
LFQpguyxbQwkbGa0TQIWYGP2gYVFWXFz4lsruLkmR+mQxY1FrXYM8RqQGaHR+/+/
Wp5XCe4Rl3KK8x688XZalnek1E8HWYeB4F4WLMDc+Nx59AaeVKQ+D38lvwllQtOX
G1l1WOz5xUaei9+nuAxCoySLlSWw84fkZy0moLw8B9bZp11fTk/5yNbfI2GzpnU1
pmpS6krqzlFIkch+3l0srcttX4jyPQIx8jAFtkYN6LH6LN60KFwnKjfwFpYuPVJR
Q37WZKrYWNDkr1Jqct6B678gp21xPcCZKKFxpGoVWQZiQSi09/3IJRibq3bW5UWt
lOwdBNEu8bY9MeHsfHr4TbdDT3M68psWxL1NLGFf/CObf6QMHm1udhr+rm78RGAz
VqmgBOxDM/OjgzEKO9l8ggTPNQ92hRwx78Nlh7I0LBYC8csygSQNuCDiFsoV8w8f
cUHRxXndQ5G3EW6T3vqYShsjKWFEticfDpWgHTmK3cCLoH6zm5qCj8Xb6TzkSf3s
FfMj14rWS34mmNEL3KPe7WqvAFhNH6JF7PNTaqw7qB4OTtBkTWLtcHjlQ/dEHWBw
f1YycbUzvo/UYStml9pc9o4cUwKK3Hi/Llmh8IOCJk90i/H3JEyryomazC2ARgm7
TgjTaw/KyYf/tU2l3jgHCo33ZRzLGKeCNjuRaKHcicV0xlniJsz8LBOctjkSqnR9
RdLzY1hIc3R3j9l6uc5Saa5QbajXNEWokHmbRwmkgq84RwE0bca8u1obBtAxQxKp
`protect END_PROTECTED
