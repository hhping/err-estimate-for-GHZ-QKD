`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9pVEyA8jY94J9QZz4+FWISq0+oM38VBI/PA/UqnKVK2QjzKfdkJ6gOe4JlTQxcs3
okwYAQjF0p+W/CPrxLUV8/e0uiEXS2lR/ERhiURHoBu0gMLFxtjuZ4FrMhycLdvE
3u2MI31QQysBp8GuxWZR+D3O/0E1ItJfnv4PECrQbwOfkJNDOS5GlbeoeDxn+qkF
cIxZ8GiJiXVaL+jYtMmS1nAzNWI4sLAy4u82f5JCuP6XbmYpWvAal2wVn4Z57i7m
rMIQP/V38MoF6rJZdtCBoSa/Ho1bwIn9PiEv1U3iDuBxVmoReNsg54i0DnMUKFRd
uH7pQY6JhRLg00alNBqgZ0y9iAuLfe0J0b948qSqyFjK1hCCBAon2NcQkv77lBJe
`protect END_PROTECTED
