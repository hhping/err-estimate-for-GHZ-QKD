`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2I487ei4zRdGAZRLoAFvjqe2wrIZA8nB0uXsHQJEs11+WC89+K3npT8ofWBnuRVk
jyz0B5pPw1sHbqa4ICShZBli0BoVkaZHzlUZF3nc3NXSsR2xpwsEqSaw+dGww5Rn
dvGXgtI/HR+Hkupcp3Trk6BC4raVpkG/7oroYyWmISPM12AG1AxLevb58w1uR0Hg
H2WQ8pz2E03qCDNvUwbr6b6URJdIPb+Ar2J4MDdAO3EAeDi3yFt1wjppHGINaEdz
r3kRE5pvLZA7crpZiSmxENfhbQhc6x0rzyCZ2I4E1fG7jsncT+YXxo91SWj6p8cH
dRpSfdKOEM3+Oq/OcdK2d0gcJ8Vnn7Zu+5ZMWND/UsbHucqro75VJguyXo7Wxr9x
cDh4KiuGCCEaNys+n6/AjFczQ/mLcBpst6D1b6nvFbTg36Se4kmDBCY/QuNfL7kA
HPqzB8ToMHn2j+mdDGRxRATLUoxue8HyBXIvdG0DhptHTG6lkKO67JRD2n9DLaF7
3RR9W+BEAj3lGaQRsFJCwMOxq9yIEodmJLdqtzzhk7Md2Vyo6pLvCDJgs62SZmz8
5AaYK4mc1EP5EEFL7o6QOBPujQ3TTt6mb68SN6BjDGc9CqaMEdQ/UgyACbkzjkT5
vaRxHgUA2hQH5TwSMR7yztJfFUDG4mCfg7zI+keHnwvlqGp4JBIxmpH9kPhtyXET
/rFb3FimN09WHtKKtVgrfzdlBfJdwGa38d1OfbCUd395ng5qNNVHy6seRDIwj+U4
7r7H6HH3YpIFxn2VUInGNYcRsDO/lS/ZGVyWqt83jhM60NxfY/ua5HX9snfH1mzZ
Q74Ec/pP+DHLkuTjccElmoFUvgTe6bj47GnOfEhzAJrp4COJ5An8butyYvjLpTf+
6P8ytOuhEz9BXbT4kqFhMI2J/HhiVDziF4y3g3XZTxzUnhmIqcySoIbyHdGvHn71
NuLPYxpygfz4p3W5Xt1HQ7muweni43Sppsw3Jf2Bm5Gj1BXJkey/g1cnNlb8MBQ7
T7xwbajvpU5Xxerejz1fW/zizhAYprcHhF3uM+HPQDLaz+e8rrCFxmY9e8hmY0St
z7IzHo8IzStxyLTmuNCaUDpub3bLY9iS5j+f3+Y56VJ6/igr76omC49pu9TR6xhD
SmUZUQMeXQGU9UQ+53btiDT0uQt/9Y965sYo/L0RJKh2qhjgtVOoOgOkDAj9ju5A
uoHDIj9ZOgWaNr1JBqb2ir9uVBSIgN0PFE09aYO4R5n/7ckw9t31J9K1gbZr/v4I
5lQdslggMczQ0B4gLOOeM5N/Ld4L9MwVX9IbyLY36GPccXjizW6weLSHm9Doxq2v
2vtKfBynz8HuJ5SyMcNv+UehHDSqlTat0U9tA4pZiApRSSXOkp7jLRWkCcK1Rn0V
ZdqQvRdiS3BbN0mwDWif1xjkfcrrq4iA0ax/wzxkMmlzvHyVHvEIloT2A1VX/mUu
H+DY09RzFgkoOQLPVNLNCpVWGDM+cCyf26/A7zMiom9IzXp0WtFjeeNJvQ+QnMOA
sJJ+Y+FdlTMFtPOrNvmUwmh4vDtVv4qmhMwo6ap8QkCUdu+qlpgfJsA1+U5GtkGf
Ar7wjG5QQW1Xw6UM7lgs2d3T8K2uUWBA9Y36IaHgGZCq/uYsWZuw9p3/LzA5gpZG
os3aElAohBrD7H71+jx15J+a7BdN3vMKa9ure9VVXREkhEdJakHStEe4QqOgnR2r
H0ot/3p7ZrxMEIjdAiak1IvXw7RQ7S67fbO4AVOrRM4VKCMy8vqA1D8rmcjs8onn
C663+cjoBewis7sCWvSvnt14dvYAHTq7P7UG9o9fDCjVQgDzvNME2tDRgU7jk4Ko
WNeJPmagbCpHMJK2Q5IO7dhprHx9bOAexqSb974G1RygfM/SwXfVFnnC8FUI1nY9
427Zbn/ZIn0pUiWdWg+LG03UdpVSHiY4ov1gShgsMVT2SyzHLLF8it5L2jxut2vv
JwxSkqabG0UEEONqT6QlB5viqienpuHMIp9Z1IQT9NZ6Pc1UnyhIzpzXZ6eTXSgE
ReolEy+ntiwKuEUIYLbtuDK6WWkqMB78M+0zSOvAw+2FKp6QSsoIilrrj/S1hT9k
DSpSEg9N6e6NIBd2abSdMZ7ATiGqjCFc6pvSTjzSgeO25Mq+jEvO8MPP601/4gtE
vxl/J6Kd32QEIJ+pLprP/hA95VzurViCICmCnvNWfRgMeTlKMi1E0N1OrdC/FXSR
O6LE+AOJ9mrm+MhHZWAlX7GM1irtqdDghKLiahKAaOdm2nHYUgvFJNOOAb6L8ZZc
mHRvf+03ZAaG1OokbDcB34l4kZtjxxzQCFwEk+mvZ78Ss4DdtT5dk/OiRmTAl4yE
PNUceol6SoGOHDx4oxzdIwLWWKwMAX2+6OcvtTSdbXCeBxYJWiwCLmuTr7Tp8jag
AOyZkRfzpjYSdf/+zaivyhokNiMiI7Ec37fur6xSm8kS5vPc8u8rGXHTHNzT0CZ9
nN9U+Ail09BEJzzDQaPlIZF4cZM5jAnZ/c2snoF38qq0KXjHX5A+e0js5rnIuuDZ
77Pft+CCvLfhmK1Y0NrT05IoI8StDYGXuxZG2CEYrCiG9LbMF79XXHc/bf5aA8Qg
ZINFL+K8FCHC1osyqOSMXRZi9LvVJ3cb6eIdIs4b/9Hkyy7/gVdRaQhbuMXF3MON
DWjXyx2Pk0RuLU/01KCflNjXUwo+hUjMBz0V83K8AupDpsUb32mDHowZWKIPD25Y
eukfB1I+nKb4O/GCpJLrTmtHvoqjA6rN5IhIQFzdQz7FZj1U7h8XutX1DVpoRZHD
0WAM/sQ1DOCuPxrpOhfZI2vDuSmCDTZhaneXAExMcvZBggTxkVOJPuGUqRsnbBIb
8AAfRcnMus9MolIkVvw6je5Us16Vv5WVoP7LZEiSB26fv/7KjYQuIlMGIt59tSre
6XpZ4Gv67by23GAdd9rPcYSLRBhcBgV8h60uOUeXDQuh1vN5RoJ5IXVw9UpspkZN
k9NVlj/SdaOTi5uQVG126HDNW7rNTIIKc+dIZVz8dp8QhompXKrxZxybGQLLudrF
alcJsmY/n3BnuunXS3fbyuSeU0p8GBuNcaIjRlfIwCgYXItB41OY2ijb7iwXSXiR
dU1z61Ud4mE7ZP5TGQnUVWHwXqtXoENWM2fAH2ti4ODdUNWBv9XrK6nJaZBfMWrI
+esFuG3TRDsFSruG2exXA93g7BkzgVeyQcEBAJypJBrLjT+SYJveR2/KClDi62Pj
oZCaDSXwKNtrK6tPE6UJC+2bNHyQwRY0RrFpTBuXLGdMmZQqIetlvE0Nk7dRGPy8
SmEx6z85Aso0QTZXUkGU5Qk0tHYMDahaWJhzfSshTptiI7X0322P0a1nIMtqyU0y
d5GfN3vmdqYioZ/2i8CkpRygaMVIn4gkYKWVE2ukcwZlZKVvKUYKLgBaNOVqem3R
VQDbR8Rt0iDWUvrJwFnKv/bn5JM8RkIZTYmzW2xGnWERc1Dq8tYt1dxy2yz40cz6
dWMoQoKAMFyY2uQhVsnZaEjQ31zSTURULueY9rsFUYcwwn+RHKE00qHh3LVVtEoY
9A9vpoWxwwAG/Z9GG10Nr7iTcRTLLTrbYtW0yvl9aHNPCYanxZE6n8GkKVgb8KgQ
62G+JmU0k1CzNaqplORAUlBGW4yR8mK8UyFB94VdaluELnolLTPPZ9p31wskVtuf
1XDdPOMCwVSz0GuzlBQ4eUdMgYuXEQ1R47K1FP4LB0F4Yq5pPPaJr8MARhZeYV6m
/tR8SWzA1w/tm46SuWNIclYhUGXq9v6PzJ8NF2xWrv69SDQbGPIA3eMg6zpqIiw+
xdGjaB5A9LY2tzsbFJfdAfVBMtP0bb0NnXOeYf3ZkZFhNmWCuCnf0H8g6phsRmpE
FBw5iZKD/BX6l9DmveTeGz8ZxhyV1lDOQ8Bf1tt38rIRfYneMwvFDUr9OPhxDPbS
jy484Sq5zATqkIKZVew2FnFwjh68sO/0ZNLqp7FUTadGHMz78VtW75Sv6KzmD5Ki
9BdoFnHlL8g9pQrowSX2P0rp+65ejFiiJR2cYKevksJ5gOrf/Gs/T0UMoGJe3aSw
2AcVYvuEGtV9eeE/qayj3p6hKrX6mFSt9K9dvW4CqOQJrNicGO+Y3HkWhQRy8h2p
Q4zw2DcVy1EfrbVMg6HLnTyiFKYAAs3c3qSLFVsjFRHNZ2EtvrRR72cQKS1Dmar7
r3Y8iqtzJLEZrwlSAdwbwvdS+xahNKEn86Tl1CaYXRqLujHgSvKKzUL2cM097GjV
YxU7rGkscdPu0yo0Lvd7s6dBhR+tuHzXHjBg59iirY//7xi4zX9WHitAuH+4h+/i
BiB5dOhfM9Lfq6VLRoUrZqGXIGGsKe94JiIGr7MQRfA0hrYT1l9jot3G3vltvu6e
R+ATevwCBDtyZMQygVvL1Lol28L7IAqGGK7la/rRQh5VT23kKd/WgmY7EwlXT9Jw
f/mKQiSZhTudxOjIxBZywBnz1F2XncyW4QGdCmKWDF3JhyjOId+/77YmmOMfdT6P
XhB2Vk80LAcXSgcowucGktz05nZXyryyguEAH4hQPoDDdOXpXNSUGC52vSCvkmXB
l/15J1gG8Dsa/IFcJykmqg+Swl7E4rY0ELJtvL5agxESzbX9OXKYPA4D+9DCIJ43
2NEk6zYJfYxwr2n4qUFkKdBs2KewsjVhkMIxH3LTxczLar1WLCujLbIJRkMvsuRR
vBflLsUnZbOvcRlPKzvvZJuy8a+mBGtF1UjIDGyYwbj2k6+WCNZ/+dnaQo/H6IPK
ag3E59+JJmqIRkUSYg/axFUPxAHnpZNInSpmzMfweEQfiXNKTUZ1WHo4JdUOtwyO
xhHA09GJp1zyYw7lb/O4AZNWLl9vM2d6xbP25xMVyH/I8GqLqIYleDYisqQ9aYIK
CN/qCUwKxycABQSX8eY1QQG+c9XQkDK4Gqn0Ogj51aT79Qm96M7EfhjVHmr17SJ5
pS9ngDnzJRdxkpfwVDcyjYityg+db6t2W5sjWZxErdDKaRD54xw+Vnv6hhU1xXw6
bYbfNx36GbM9jwmY/IMAkCfg8a7aGNwzC+xzKkg28m3c3FoPpHnQVTAAnfEsnxSR
XMjt6Xypu8JxOvonptta5/ZPyuZ5lbZK4yIBun2CKifQL9As/XJVg7hFh8gBTKNC
MGwaHOrBvnttSxHERjjrByVZrnNF0TQIbJWjy7s9DFUucd/N2YHZvxsFVjwTSYD9
Px9nY82xTi/cLHvxpUKwAzZsJI4Fuh9hozE1VKwnORzQd9umDZwiG5dcya4y2yX5
Og0HG/5RP70pQ7kpjbxOldHBrX7nBBDUzehB3kLxIbTWqEdOa+1k3N6jq9ySkBvA
+kaYOxB/6rlRXiUEGPhRMYHEYw2ndKGH1YrQ+AQu5KpQSHa9SbIBtstqHoa9zk/c
dbfnyuBgT26shlPDBArJ5jm8G2Ws6KiVB/i5zXaYlSZTC6PulN4fQAfplxBwHYPn
jFRti7falGIbIXjoJGgvZPE0GYGfxtIQvqwXA6IvCdQFEvAphUAhdiGRHXsBCJwQ
oIByzBBeHf8CE7tchCYbqwlWRz1FdzaXVzhkX6nAIFKImPm28TEOOLgXK23upXUR
d/clp2seR0mCPSrX6w9di27d530153cld748RyYi8YHik973IGLXR/69alDoa33k
o5cq0O55YtQZCsAEOLgSFxKrI6COJg8hBbuhrKSkRYFiSd90ZdiWJWMqASazgEQP
nVoZwRqoGhTygUPfKY0+dZC2ckOK5O34+oDD3HwhpKznqguuQ4aIXEJE4qIyQTCa
pgU7ve1AINvQje2Ouz9WgqOXp6lTJwyA4RtTWKKkTsMUrMqrVPfvJ3oxK7mFOORc
FZbTaRyFrCFkI8RWXKPRkgd/jM0C3now6jpH4raoaOJaIrItycgXNtryXv3db5Uc
hzOnmsInsWcamamnJvX4/J4V3v0fxs3XzEJ8+3pMNHh6+cxVLl9eIR4TM6Gv9Mx4
LoxVe8uob3U9H40esgh09uHIsYFS9irYkkIT5LArWDrloW03TrcKM0D/0E6cETyp
uBlubPiR72InNdGiuuxzAFd08WxsibuFbGt93f8FOwzRcsWUbGGvnwJ5bckzdXg6
zIjZD3XBbc4GpIxm9TxjLTO5oS6mq9/ALpVO/pPZkHZ5QxgEvCcALwM4nxs9QxOi
wJ7q5bcyuHGjUeFjbrPtZz15vz1I6dLGL/be9sjfeFkexqabRMrDmHZD78bJKNGe
Ci3XQqLk55iZZtcCnHdXWSF7PPBIyIC918QepTeh6hTQOlFv8Eb0Kol52JybNFpJ
CbYbx0duMhl5LgyTzwsA/5GHREGaTOUWsOf6g+KhEjhlNeA9+xyD9mCpUy9/XGGd
OKWOF32fLppPHWWTjWOugzpjB18fslTYv2xjE2AZfyu/d5KQKK1iPa5AYZPl9f0b
KsGTu4Oddhif2RxbY2OD/TQl49k2BB1SJAF5IjdKW4gGXkOxsdEzsZ2m5ABOjdim
pqjosvXeLa3OoWjpMiHCBe+HGl9yIiAWK5tQaKBjpDyAdWsjTBmvQiEu/Gm6Qbwp
O81M8NQwzpw/cDrKmKxAQfFa6ziCYVOk5KoIUrFx02KifNiJfzM2Kng7uMmTvOjK
Lbq0dH/mwVKRDwCM3yON0p1Eh/gpPchIJSmbGEix3bZoe9rJlLaxVXVj//2uarNb
Me54A/fxmdIWP3Cs51pWBU92pXh+Oi+IeJhcsmjuMtQ3t1M5xBVSqjcFZpmehisQ
EnRZ4FCm+BWs6BQs06cLZseabJod5vTwFRck2v3+tJlbRuYHDQtJkGXRWhcMCzsP
oGXIsctjF0BkwJ6zFg6EQTKvaDjCgEPP/rjMl2864YOjz0ZTV5nnVEHmk3FhAgD5
dsnQ0d8Q3JtqtSTVmI7qEdmW9fnzHvwrReDW1zRZuh0Aa5Z2JCbrl7CePmDcQ8C0
JSgX401+eg5INzSi0BhjhKEm6rsUC+6wAcHYkN+9RFKpVBBcWCFwy79vAQUsikkr
93IPqI0G9ms+EFxb5XzD/e8A8zEdGmSJ1j1QfYbwtXZC7mgfsA1Dp8DDcug6lJ9x
+hzm3QcNDbiyqoKSmh1kpG824p1f/IsJabuInEKHCbu2X+oqT8SLVkSaUbzGzwJ1
sbu+JxnHl0yytevXm7jgsrY653d1JKd+59+pAlFidn1VQLed6Apo8TSZOQvGTye7
OckN2PBtefvQK5WIaZdd/jJQtl4znJWJxPAO0ymClRKyOATE9hYTqPZqQbjsUy8X
xEEQ3agm4AGSgIss8Fm76fzcnHSLwGyegbLRhZu2JKKMG++630okYpRqgtwbgx9B
Vb1LXSl858N1CmFpFC2XGRoLE6sVdWQ2fPR4dBt+CIL9s0pK/5dYo5Atgcm+QzgV
WhKnJEgtON2dFYom57eQe3Iwl9mfkoo/ZFAPPVlOj0KTYIBQyygZ3VNSpiK/O6ib
lu7ap0/oBNWqfjS6PQpme8QmQ3yJ5oFTiceoExJZMunHtc8a43921NF2b1XIQWv9
L2+LoATVRnWUpcTapHZ8j7T2ZqNteT436cuOFo3G+y+lLFz16VpYdZs6thea+Eq5
Z/+YEuAADZg3a28OoXNY32PHrvakVSzkaZq8+Ky9OGyA4YzD5viXbt52QHR5q6ky
zeMh82Ww5Dx7raNpu3Ym5jUeBLd0Zn3TFCXSekl86awHQuT8bfLWKmpd+F+WMPUJ
76IR31VlV2pht6gNqVS6vSi6LyOstswrB5dmpU8W1Ocp0rJkaGVcu1LN4Qn7pivC
t5w/G6QbUy1xmfYnSPYkiXcEgah9MKqhEwdItkL3QTpJ7C+zg+TcpXHPTl2FT3RD
DuTicg4hSMMAe3cHPmHHdmIsUN0QxwrI76w0ShF6+gW6WJ9v9WDwafrs7rR5z1uC
nemVSMfISdRBAIf21yD5Y1zNVpYvKhDGMRsSOMsv5luwVLYrMSLKCpC615VWiKTT
+tAb5HXCDnbIS26yDoIwIaOya8/dkepqpirZgPaLbgi5yWDBTgcRWAW6oIMb9yhK
T9FBvIsCvBKm07lm+VBa+Fn+kifXG+FxTsLwDL+V+pdLkqiSIQyaxLakJUfGEIG6
q+y7Ct8neMpIbXJZ0GFlx5LkbEbhZ21kWIphaUWyKdwmZbUlnNmtlNWhhZDBWIPj
PgofIUGuvPnZD02a8nhZGXlG2aJvcE7d/4MKKfPN97UGSvP1qlgSdnBwuCvmYC5v
bqiAZ90zjfGzbqiBbXr7mARkHGXLWU9ZtheizDznbrg7Fy7Lpjo5Yu0RrJ/yZlNt
sCZO5KId11iT92v1FTRis0eLyG9KNGVChBcrkwtjhn3jIwRfL+j6P0Gpaw8gmJiv
0eO3xNL4l1ReTlIFzKEBZm0olik5104CDTEgklFoegBVoLv+IilTPd87OscQNtNy
zbVgFQ2Dj+lokgb0mnC9iW9vAXzkvjOStPdTKctF5CgOhzTg4Dcu+sTftAxIn1ss
cJcnGVDigvUJi8bqk90MrwyeEtKT0jlK6lrSM01EuYmD6i1ps1Kcx8dtQHn5jTRs
EUhGrWePA8yEOgZIKE/Hs4HZXog30WyKpQpZ1AVJzFZ8QtmaCI2Jn94udsWZF+FI
MWZ33/ASB4MGkzS7QMtIp7IDQiNHwB7jrPXBCBGCkltry9dKHaEhUjLq1A8o7pLw
9q9dDPyyjOchvtbGJx5hrnxOGPU8kxGuYGmEqVAGEUI/pUi7r8fUyVlrLKYghmkJ
dH0lAp4qi1pSy64yArIj0aN6okpBuhATvOjKpFy7yKFGuzjBPQL3nfwAOtGwVBae
blfoWilLw7UsgeuHi59SH8A3IRv5D364sUJARTujGkfCk9tjmWhW576mZEofjNix
FihjrqCRJRBwnHLTkHL4HcCuo5msUYA/leYuKyOvCSeRYEYgdy9CzdUNlA/yW60Q
59R+h0VxsXF6uFyOt78y9CAn8xiExN7vmiSVnJxnhIGrfnqWvUW5TsHXDj6E6e90
XOK3jEnnnMnw+WYUKbWkRsS3pn4yFolM7IP7fA0bESjBW7nlOrIJebBjh2+Y8lhO
TQxS23nHbyKvpUetQUB5qGM372P/MiWaqqx2KrtivnPrdqUNdGn6VzXS0VMw8SDP
oDjxtzWjrR17WOiK2qplU64AzGPJLTLw1G+HqzB8ROD8kd+KVYnCPTlDF2XT2QXs
hkL+IPDmqV1En1iSxD6x5b9R1b9KHqHhIs0advPXp/GL5DISMrIKhwES4j/V5APt
XS8XM44j17j9dSeqsy1YjS8ad8VX7wpv4qdKCZ/7lo/MuImKB2VOSqDpUnOSM3iZ
ykiCT4bAYZVgXkSImkUROwVrToFJOFHv+UZ+XejSut7jy2F/SmN61AJxWRyIIt9g
CT2joQddET+TWawIgJJXKHGt3WkjnqG3NxVfMVTzp6Yc5su/DeE6PjExTjRd4sXQ
1SkL0VfuiXo3BgdOTohlYogchjJFaYFzZ7nHVCUUemwr/CDV4o9IT27wQHCeCw8D
q0RJVqXpr8jDGVXf2x6KOdfmm9bgw9CFFxg5k+n1gM2iM0uNX/i+qjjnGtsquOtU
a1u+NGdCWawjWMYARpo9RJb+6mgkudmJvQqJ7NNu/DXktqw5XkO0240BBY2GOqbo
AG8qC5kFR3JcpHQ9nf3tqHppxpYLsKlg/lCJyv7rWgjBWwjCgkge9lsaFXeYxxMB
PhcHQT9Ajc8GNgs8GZWHN376IbmLDUEfUDuGDWQIm+QYDovu1JhDJBMt+Q2MCfIa
aiN9uLkE1pBjaqr+ORcnHz6jlKfFJVHOnMV5kFDygb1zwyMt7tjWEpyaHCtE1zST
EXzulPJ7WeAI/3L+L6uwg5vBzwhra/1UWRD+7EYmmS5PqEnRJmeIqsmtXY5VB0Rv
zxE6pf0rsYyqimZci4o1W9NUquF8NIvRJabJdtj4UHCqPFoOEhlQ4hvMvJiwR+7V
TiyJzJYSr7xgW/OjgLjvEDUNHi99JY+uXtCdGSqyMKseUACcyykwAB1DPMdIfWtT
y6adErC866FCfVn2NEyvP3chthROrHMclhaIe4bcbNx5NZYnmtRBHTJCOTKhpwXS
7srMphPjbqGC/ttxVSRRbuRcEWkJ1A9gMvD+okspwEAG81wn0+UDTLi8z+y8gru0
RGUgA1sPP3ctIkeZkY9vpZy5vHaoJ19lfMGdZprBrYsaVlJa4IvbPbc5ZKEs60++
LVvlmPPmcBg0eHnJQzcEots+P7/Iljr3Wu+otU8UvFxMYH9/hF5mpMf9NZpAhbtO
aEZZvEmEsjdzOQs+Iqh77yjiHaIvUMkeNrJjww5n6U9gq3BZsh+reYdNjJQoklwj
R2Qya/wemOB7NmmeJUQezaj9bN2RSH5LHACr7qk+E4FikMnTeuZyf8LK5/o8mVWc
gLti2PlNZslRWB5Le1FUbnvzQWgQlFzCgi4YGbVoB9PAU/c0Igea9HkzGOClkwXC
6LeapONqa5LGqnML+UKMDQyhHiPV3r/83n855kn8Y9r1OOaFFSL/up8etyjxYiAW
hCa5RNAk0ZEDVcCX8X/t+cKhM5u3vGf96/gAu9bMQ38RG7q1AbQnqdxG3uadsEmV
tF4Ik6ie5t+c45Fu6bDUH/ZMO6WilpBI4f2KjT3VNDvDBHoTwLDVZi+7duEPjjCw
UXObp6iJ5VDL0h43fcwI65BqbvryWWF7OoE53IsBvwun99bZBokVvVsaWMubdnWm
o5nr+2ji8fuq/3mjTavGkJJy90IF531zqmOGFPkXzZ8OSFtMN4GgvUuXK9HQ4Njc
SsvUq39Ba5OZVuBNkRLnkeO92WhZgFi0XLLIT0AZn2fg0zOIhc/kNj3CjI8IALhz
hOGTz7Sxhwc9v7O6HlRFXJH+OD8snIc8mmPAZ8vu2HqZteZMXWL7FEMN4zgdr9Xp
PbDQEVINkVNZIbIV1B2f+Y4TxBsGwsZhucz7mLLLHiGoR9DClSSFR0/9ZhZHwPe/
07qh20X1RR0mvcWgLuEUA2bLRQIf09hESA1WLjdghyUu8o3AHoNaFX3PW/Vw8T9w
do6FbUPp4GiIVjdFtON2O4p8x5j6B3c8mMI678YTTZ49Hxu5uVASot8qlvI+UFFi
Ys0/hRe55W+4pW9jMncSqiio6Y10yZ/zmIMiyioiIyVzstXpDqB1T5CKOZP8ygFp
pGGJGG06WGTHau99NHr+5Sx9E63122FWWi0VNsOXPUmBskXUig84jNoZOjpdtY2F
WhmxzRQv/+XHD4eA4teo+vZSvXu9ajSbz1NWHXT+VBJW6oz9PTji4kGn8PEO9TRq
qB3b25k2TeU3DsngY3WhjPQa9goUwqHKMOop13EmS+kCBT9dEYleMrdEcxmQ8aZG
tbvy6IyzfMyYOGMG9bdXU336Sxn37zJMw21nQUEQL+RAt51qitcVxmCVe5xPp/f1
juXLfMzi8CcN+u1abI1ATJM+Fd51zuAt5nDr1TAL8J1payBGmN5KxnZE3wCcWxyS
CUQv+/Bl4GntUhGTxD8rmpPijKaQ7iMkkE/LY1qUIJE3rLgJek1LUAOPSpYaJ6WG
d8NSZKsscpTbSyEKm+QO1EcnPFgBKzAkcq8JKNS8Ds6Cf6/Kvdxup6pbb/zOATgI
6ux8vT4H+uSNUcmTZYfCo4rpy6rUwGiLtDF9mz087EZF3czHUkufYsqpuXTNkhGS
5rMdBZRFB4Rm7O5CKpqe2dBFp6ni2Bypxt8MhKBnsRd2brTK1AsjEQwZlEDjC5nD
qiSQkUNaL2IC5WK60aBBjBekPxtH8gkC1jMQr9kXoBXjl1JChx4hkyeD60MeOBF6
2ajS9sz0dMBAZA737UYq82yVqvrICyfCMxp61bU4BeM+4tIUNdQFyqwpcJjsDdRd
343CW0p5L0kLkc0aTq5BZAfDXriN4BET9+g68/kP/RhbFdKTZmwHjjxgu4B7b7aW
ItclydD0S39Fz3rmYcvUBMEEOuvVtyufy09YYirRHzCrL5F1ZM2HGERBwb7qUiQh
bH7ISBOwk4WIja8AsGYT5WOZ/PgHQoSz5qgxPgElvV/E4HEAfgzEjKjKsAkHuXun
S5dQpKzokHdjtD7nrew27SBPIFuQ0Ldxkpfr4sYrWngx7nKz4oj4v9f/6v6L69ZE
fSAPy9/ncWXTZINSV7M7R1fgMyvDPpoY7eUSycXuKLLOIxPwWKhH4tH8CMRnEFUg
uQZArxkc2YXhGCMi9YnSWZvmJsVzUPvs880CB4AnL59nTwzimGKPTeJ0wm3QnqNv
JdoZIHeUbflf4N1S14Ke/Uw+sh4yKSTUdf9x6Vh9UzDzr4pYuhgiuwyFtEGb1dMp
ilPeoIppbwlnmTCjGcneAxKYZCAu5dAVwvDPPixXCbFX1kp0rf0l1zmNHOwpFd3z
pD8HkIjCZKDrPQP2w23VARIdx4DdSCC5evSMtWuPkNVwS1EbxOUwTgiq8PuVDlzE
O8i7Xm1k+ftARLXPS/ZG1wAwVvru/8aFsgLrjI3mJ+SaL9+tkYMzC6NJk7UV1Qrp
frfFOa1TjN/Hyzao6D/ilH868TnWgvjIpfcnn+MPMxTUrF4sfPkKjR25dGTsMWop
ZIrP3O57rtQ9AOn6YYf1EAWws9uNMrJ3RtKIODx0AXz9rca3pg00IAJmlem/e0tZ
cU3PYqkFKwB9xMOgLODWix4OvAVp5SFOWROkx3p2vb9qxOmlDpuFDPWJCS028EcJ
9FSvqcduOUhQJbQ2p1DdWyjjvayH+o1MvhaTuzzARIeWpsTqI5G/4X/Qo3ZjnDX6
b95eECbXJBjQJjKjQKX7X2/mWlBWQdG+3E9lv33Kuv6B8f1KbV/YBfWYQ8Axtuzu
Lr2xX14WVKucmGJ41PbJAq5vAKNdlt5Vz9WDuuQTbkqtLyJgPs4vhi5kIuOoKeEh
U0ASUMWiy33XNVUlRKT2fI4slZH74T6f8wqFQeWeKwyAZfPpU38LUq5CljYJ3zfj
wr58FEBXxIDlipX3UqU6ceeLm1eXokWO9/WioUWiYlOreHgONpoLskXwRMyqTfvg
trMBu0UjlPcuQFez5A3OKI9mGN5Pdo01WIazfNNeFaW06CBRJJljPcp2aQN4gxNG
SanvvydwsUsW71SnTtNqU2Sky8bojz9BReXb4GI8hkFwxfFHjO0oiNSD5dWbTrdr
0uNQhSGvIZ9YothM3i0+0jSxe2Dj+bCUD7MKWu44ILBDeHlCcyyqMRo0bYdrNQKM
ExR5o64ajF5TD7ZxN2pzluJA7J9TZzeHUKlvOLXJaYAFWfbQOS/cALFm6My4q6dB
3hxintUSxD4YSzOSmqPvClzlEx9+4uLg35hb5JmZd3GGbEmYZc3JJmRppI4pFB4d
woMh+qSCGoPJaJj9/DR5/10iArX87oiZuZ/JyaPYfqHSSLkPf/VW5P3QHXQWAWlV
IKen6CjZ0TmBgHZqMamh/hHCqPNmElqLTO4/JbdaIuuo+iLBdwTkZ3NESAwf0NI9
mxkhlSLdgjzIuF1Tx9OzKDEU+6ioYzy7yYMTSVtZyssLI4yWumu75cxQ/Z5zb8wp
adkyTRc7VcbnFy45k9cYLjX64rXk1ymlj+KPZui23ADPQgGVWgbnJ31XOvewyt9I
DVaucS3GqRAEAtghZRt7ech537a0ujm498OZS4k7Q1DTubnR8mN4wfiQ9fedFrqn
vd17g2oYKsSiR1+5Y4/6zmqhtWAwf2KgHuCsFUqxLKm2YBFWln1Zpz3qrhMYXPBu
T41kyf2IfHcnoUkAn6TCk/u4ttd6E065ctU8c5wVJJ60G6Rx4fmtBNwsg27yoRhx
vzX6vazwX83WDI7hldsueBI3io3uJfr+rR2M81SnAdicUc/NHs4+ekzC9f+qsJze
EVpBz3tIeZp9s373YPaEuvD9rncXK1MXMaX3IjL/Zm1YdtzRfp3xbgBn6jhraNep
FAojvVzwzx5sTi4DwpsiWkrun3fJzBGNLFcGu7+jMUiy1366Vnrx8IcjQQu+opSm
ZsoOX2YB5safTyUV21wNkDFdlZQbJeF2rqFt/qXT6NpDRIa5zGwxpXkWms1Vf/Zf
I6eJ5JUDYnrbiX6FlHmuaXJsHD3gboMxRhqUBpke7c08XS40vXRbGOBTVcQzUw4Q
XWLAHB43mbTtIPat7QmhfvPs40M6Hc8KI3o1sYfsSoVc+KtRKfbtAV9ZpOrTEoIA
+ssDFjjVHL++gkMSSXE68rjPtkCewkuobuIzeEhqafgI6bThAaDDRb7a6ZRigYUK
EXE4aYsZSHJVL66MeaMLQf77FCldWtMVvUxn7IQXYkPTauFYhU3eTAqmOZsf5uer
mNr168S+DyyzzCtFMeSEdjU4JyYm9isFh2ym8sqtcaJG5ljIZq/U3kbT36rVIxFM
F48QeT/v8WrzVcW6uT5WjCNdf7rFSX/kqyTWWeuaDf+5yVBRrSESNPPL/Vy3U4d8
+pxEDG2N13PV6SJoukJ8z0UQhm7dk621cgXzcM24Ca0J2MBFfbUTAXPBFgePy/tl
vIOQrMtQB6x/+5MC5EzjIHhMN00EYKvZs6g5Rw1pibhylEHtcykTpfRDA7Qd/XAd
jiXr/OSzSXpCInxkl20XGJ56p+axYm7oscmEkqKzqAh9ZznxPSBf/YM7Nape9RLp
lMJ04RXaCY4H5saGofdQPWyjA7BZAncgU5Mh5vFygwHUbjTz2JUIk8V94oNaE0d1
E5xYmOGpPQ3X6N/Q5baHLqyptHgdpI+VHbcFvQS2ymLO5gZAEfZ89mAVOY/iksQO
QpJ95/IeG4m4AK2D4wDjJRNbhCnh7wKaegHzEUcmWwHxyNR0KEd33KLZta9AOW6T
kImZaMEP/iTWLWz5h4RRK16qe7EqT1n9cojn2/4hvYK5ylU8rFtR3ejCV8pKBzOS
nSkNjLw5ts7n56rDYOqX1P59V1skWC9Or1v05iJhQR7pu9xTsoH1Q4eB/nR0lEah
4R080PfE+5WLKThlduhVqG8wv1h8Mzv7bIpuf61H1Cs6oyxahlkYPBa25Uj8C1ez
texILSuRgSSH6vNctw3fhx7VGqlO65O8DI21fMPqCDHVUa66S9LiwFGas4hqTWVC
YxZ8pmYRnlNIaE7GrRJ7tmug/CydqcJhY533ChJA6oYkzFB9uGKhIKx2FdrIiUK7
JI0Ychpe8yyls9C7Ay10GwN9wM7WIZFdikGAyG0cFict/pb0eZE/RftlJyXI3/Q2
hPArNSsSsm6Q9gc/7rO8VUPcKHMK6+YFx5rCMBxbwVH2yJQ+tQI770YgsUOT64A/
00NiyfuG0fkqMvoNDHGxQDSVHP9t3o4RhVbKZywjIzBhYb0olv7AZk26wz8wzVP2
bp2UjlFkwvCNq4VpdUb1Gcul9C4gG3ZTKJxATQNb/8PUQMd+nKbBbntqZlfYbszh
+UJr6NEUl72fU1/Mz6YPGNZtX15x+a6x2+Ca+FoV+6mu/AS3+1ulWMt/SFldCofH
8/DcDfXeOpoi6yQ+gguNRi3hsto9y01p2iKeGsaJBl9daIWNS+T/HwZxO9kenC8u
I60HYg7vkvI/8NJu25mKwDHgLi4uCeWuVbuHEMl3p0uWrb8ZSaOFMGaC4a4Adz/M
5PZ5jv9FsDMlC6Ns5URcZ9GaH9/6qzvl3yUhQ2Gwj7fj/wbdyKE4T9IXX9Zprpcx
caoy99tJO9WsqTPDEpZAUkdsZbAcO4JzbqysL2/4dwrCuX6Hi46Pt4t2ichIH8ma
wLgjPIfvdnDcsMc+7KWzLdRgN9wkEjn4Y/7XT58K8jKP1qKfr64x35bD9tgAUoF4
JTAoZGl6Ir6FYgGVlSaGWzHIuU6pIkraKk4DoLBUemLDVX3C41SkYIwOaiWin/2S
/nsoX3hxrCKvvTiA4GfDYm7q9T7csB0OSLsvkdOP+V4G2Rnd/XDTTeU+Kdp2qg9y
SaYjNC25lEPevaGZJTQ3AKzxE9PORr6RCOYdBFWMCazsv9zksmpMs+xWCLuBBKNQ
xNe3lCL936GYQDY6Wrb43hRTVdXGfYe8XOJldrcZE4MpsxRQEP7G8uW8t1AY+8jw
NFSLj5uzGbZ6GMtu1rDBiya2nguYgvUxC+LNYo8w40oQ5T46fQbMPRsfT6273jiC
vVkvuMimJg4GaWvb2XWDaXa5TPO1nrLSERqwjdYAhM92O55MbPcaLE3aCHWPmU6X
ASxM7DYP4ZuFFMDPPO4AURmWH7ImBbcTjDZ/P1HT5AmbbdwRWyyBw2qLCAlSYDTb
4WTgt2U+7f0ot9ohjJb9+n9gNY4+WL8mE0PjgT5m+cPm6NA57NWfVhQyko3WP0f8
oek6xCY1ef4TEbi33SGpJPAuSCUjBVSF9mTJZ53fqtxluJYA4XPyGlG70mIgzfIG
Iobv2+AJS6ZOBO5WoE6Nb8byIJ1h1StRj1BvPhhy31gXeXxn3qDYBobdkwZ61m6w
I75LTl7qYvcXPoY9luoh88uJAEqrGzIVxKBk+pvr1Yvk4RWvqDpbsKK9ETlBs2wD
s99ZzB1+RJ/9QyxgfDxqK9+u1mXvJIYWX5SoCGuKnI8Z5zmL65vighX1TAlU37Z+
OuL8407QMj7J8ennM86GTAy5ViTlpSWjnyshlrVrl6o5RxoGH4EWc1aAASZPEBF/
bbLXc9OOnmhUs0EEO/TvPBWXfPVhVXfZlqCcUPxcNQ/QEewb3FY4ZfadA7yHYV2W
fiC8ci+Z49LY3aulnoi+Hwpv96+FiyQSBM7JV5a+fENL2WAnOzgQNo9/4um1Ac5i
rNsOEdeS77Lx7OGNJuVWCE02D++tDEyvGNjq2kCKt+UEeNccprmEiepjxiYTDb22
/4Zd0jcycpd/YkV3EpfbcUm+e786A/f+1HQR+af+N4gDeIsftbPsPhjmyfBjQVsZ
F8rq7oVGUQyngoQZnrMt8Q7TIwGyK2fsmLUtCmEIykCbnisrjUrttQ8uvtyLzBpO
z0ay+sV9kQmpBnk1IjLimXOXLNUkjdFoF0+iRhHeLR+STLDBTo/WZ9QqqNibIeu8
EPc6Ddf5Un9NX6G/EQz/S/p32nEFb9xx+upboECLQXWqWqflYV0PzlsVlq28TIuz
jXu2obFy7uzKgChR1jZIqvjatyeGF3xxPB/+Og5YC3WMa5JmU9JZ2cKSaJjlZD3Y
FZZunoCSONRZOh0Nsbj1sUmhTATIyRQO4sBannBYER9ibybitG0SE2YerI7jlDt8
AD/r6K+ET2V39XWe/t8BEC3p1t+hf8HszVFLSHjw7CDzyzJmarC8zec8OK54WmC6
xSIXHHXb4rJbyI4GrHaB6xrqwo1P6/H++/Mbb/Y5NJV9z2NE0o8KOyQgm0aaiS9i
n0FpRIqCZur6ifKYPp1yn9vDhgGhwJe9laZPozBE/aHqJ00Y13g5wfnk/fNfHB2N
7ixgLjvqBl7jBB8Emb8QdqDvteAL+jn+eIpRFw1kKJyu7DHzZZj13xnMftMoGNGA
9yhUVQEAIO3iQCgpU+2OcEP4Pv1htFDZfJ1SGyQ3iQiErajIRIw4ZSSmFUJuBLow
3o+VEJ2xT9hV5xq2T/xizPi2vK/Go5vuYrfGpoVE/4Lg2A12xOU5ysOv+2ZkLAIY
4El+vYg66P0WG0KBnGZLr4s4a/cRUaonvBHUyYLn0KanPsrStNjfUHgLvX2IQnXy
BH1btNnKPcKF/ddWJpWvJucusidxxJ1I8UC1qJ2Dp+PQcycfVrndwcfL3isT1wjG
oqeqs2/VZp11Y4Ah4zy7e5fVtz/tvBSru60Fsxv6bl3UxnQK4naVL3BZqZ7IQH3h
GtXFZP72Bxu+7wLrF1uj9P5b5I6E4MT6ieg9QPj6p8bt7GDM9UaqyyvsmZMraRaC
en00ABVEni8pDySWvLfjAwvVPUCd30kMFcmaAaBYj04lqZpD8XibQcotzBrufrLv
VzmswEdpgMLnLg0KTcRjleTnv0mAkjRWx7yqtzva1RQ0yoQODBFLTZ3vEOqRa0i7
JTnzAxKe9d738PUi9OGkFgz0CWXSFEsP0zt72w1d7g/ETn26cXLk+oenyBW3ixZG
4iTd3HSXvhwSyTWepEa3EDAGIEcdxNx+DRLrD6e22J5/IgsoY8Vg1iDMGrYOOJXl
nJkJ6iAOpYfhWfqLZJ9LH7mjj+ySCs+yKBvHfjnldt+ekbiqjAO9eBYe4BHisn3h
Mt1OHaEVh3hvF6pnAuvgajc9hDJD70lhKAv5Fp1BIzSBE2e2k3jsKZorjaVxxxcp
Jg51AuSZzuZwZZf8OT3YgDTjeAfZUiRtzYLbPuSIAok7Oxk/JgC/VB9wWGbedEuP
FwGNY/vofYueJnimA7vUm7kclO9DNiqPkWNHTsMm1GItEcr5xP8E79jxZNWvFw/o
cxhFX2NOgIOYZ34OMfQMP9S+TH166l8voP/ceL/YLIB7MnKYaO57j4jhUQfCPiEO
adjI/0IEvXtv988qVoyD1W0bFvMRXtPDjYsJU/q+g6Ijm7oduB9y1/Fro8kcCy5x
ysP6gWCGu4xPkuNvX+gattdj/+D0ECgmqXXEW70akuT6K839E9eGVchVAE7YzCJV
+hD93G5tTYm3cOaeIs8OK052e1gEg0MODiq/CJ19NR+OuLh5xZO9bp0Pba/Dqpho
iTdTKrfd7Hp0yZRbQHqMmh+p7O0OQUclYsyJxg6HcpjdbD0QBzNPG8mhFxoR3JXx
A0Ex9GSnNaouO9MKCaE5VgecffiCrT4dmHOyxRfO8X9hgWtg/xzyC1My19Ejfnjh
3A5tEDPHmEJ4m7pv84pIUG/GVTr6BsE6+mloRy1MqD9iKgvFan/sb/hmwzrzBeAM
/Iy9AONhvLpIYENDMdwuRhGVRC/91py3vAoz51bEq4u5EbIq+//nVVqjnGG2kVML
f22RTYy9mq68g/jb7n2oqO34zefhK/OM8l9tf7Or7x4nIG50/HTWQPSAmr61aM12
ozvyvwWwbTq4wkKgPOWx9XcVYKy+Qc4HKyzQtGO//W07EEEmyL1aUgIqyiqw2Qth
jrDGBNqSPGiX4KtkL4gj4jKl7F2W5g4+FK0Zu1sFBKVOQL2Vu/KzzjyCx1yt3y46
jVkSxL0ts6beTLHpqPcsMUnV2QKDo2wIyRStxI8GfZNzAT+uECEkyIQBTCkqdnOe
dkE4kCAtudpot+K3a1PCPWQ1i6J+8+X7P/SYMO18kNiiEjFgDnXglaVZkaws2JH/
CFP5SMGU1KaURpBwdv4UckBEOwbv8NpNf2NhbXh2EkT/8XVsA7blMP6w4Ya2J2z1
IHVZ1J1Iji8/3fdeO+ShxQAsu39JQiDcxjyiZyy5nHorZ0nXPxSpvkh3U0TKAVvh
JpNjs9gM1HRpw1yCIoXuNBTg9vQ5elMv5s3iCwvGVQ4vWVanM64tAiCLcKdd+pZZ
S2PfKx28cN3/baFOFnVfoMHrcEbPFS0IO9tbai8Fey1vPxVwEmknzHKX8zKiTz/P
aUKJ3ZoPTfRGhoUxDiQK+7lyaDGqBis7QuLTpH+PFTVvcrjftpQSeQ1RUtOMBujI
0HyJzQsMlzMxInggUrZz5EBlZB2upk5sRTcxJ/uvgePK9kGwBXwhfdOBJ2DsU+r0
gNY6I4OiiSe75DFHbZEQq8GclbbZAYmHK2NyGt6MqyVI+KePvCzcs+TM3ds4y9Av
CH3aT50wOtl80X8WV/rY5DLEbFGE7GyaYiG1+YZm9mkjIQe5MyrQvao1OHrebOA4
vSPC7FLXHZGmK0e5HloE+WN9UUIjB7cOGW2iBb1kd3iUDddZuG7xFIMNN/IRkeX0
XXhshEW21FQSdJlIH+x2hfmk8Ux9fGocPXwTWKt1QYeGanufM4kxdyX7dfIOB14q
6gg6jdgi7Hx3IoLXLdr5OfDpeQWd29hl0BADD24m2vk9AJjsNg4ELsTgluwmfz02
Nl+6dx4OGEPajthWufwiEf9NkRLRSr+F8uSXi4y/bAWAlV/Mo2hyrS1taXSX82b/
Ai2CPISSRn7Tgsb04Ig1jhElzVyuXHcr7OlKtaramdtqT7yGCi6R1RzDj5nox7gJ
kCSAvs+C3qRS05rSdlLwkcl/oqtG3o1lElCMmYNrOpwKSkWABxsGHrFocFxVqSjr
IaBXA+41WpImF5dH34t7DQeuTz6VdLKuISAZ8ET22kEO4O9u4RiVYf8SFfqgw7v6
T6nI87zEenMKwXsyRP9L8DgQF+LoM6x5fbxuA5+5oUx3erPX68rQ9AyzyxTjK4fu
dxWIfxECPFBUPKEYahWLV8MT1nsarzmjupROHDQKPDNHncKMQXtMym2GYaQaFzyP
3JU01ARuk7gMOxjxTIM0X4m5UsUfq+nxKFcUbp4M0cr/9hsBaXX87cxKwZfDM03M
oFwwL0O+W6tE3uYjZ0j6nlCUf1OSqcjn1JKGp9nbHQhWCNMs1wFuccyuh5UDTjSF
XMUHVjGgVGcbbn5UNy9yOKNOIKAnXq73t31eMLml2+KKBBSs1vnp9ObzhHgokuKc
V7ODm7GDRAaeuM9oh/E5ihHl+n1UG9uB16hLp6iOCZ2rBiYi07FP44netJov5nMr
1/rJAQgwIsY08zluPtjyRGyrVHC46Ceajh558SbM9ALU4wWPvBtv41g5jaWQxhYV
J8LjL3nMw9VSImsRaBZ7G8Hu72mG/rqzB9tsRxLYKBBxmOBoeShHMAKijTnNg6f2
SxN87tq3KpIqtP2QogtLpGhoPqr4WEu/94O632fzPtOuuhRSnRt8srbsmpegWdul
s+7N85iyXxul8Jxe3A4fkn0Y6RY+sdMvBs37N9NQxfXOh9oZnVm3ZgPzCXq/uF8A
sDhVw0SYquYh2OcYIoCUSXWsP/9zGc1G2Y6pOWfMUSkfwBbEF++l+LQEWGf4pE/+
HF6RCb/dnqYP0wenEvvDB6A7mkuLMUJGaOrksutZaza0OfJJow5zMIEttFXFNjth
yk5WagBioxd2upW/SLuXZW+dDnc6gp1t8Ea0hUMHc3+GGKtKpCADJAK8FPpUhFXD
7jbOQQMYgEkFa4vtjfGS/3K+FCXZoJKgPZ/YkbLQJ4nJ+z2C3Ezq1t61h3W2++qN
Hs+u0VLMAOMmHBS4zI9nWvZD1csJ1+inCBL0dJzQ4sefzFbshB1uSx4yqAxmAPgS
s60cQAl1QZLdel7sGJteFY8PMx8jKu5jb9963wAlYgWRACJp4wPFDAdnurjUHNOe
sx3N0tFEt/8PSWInp38BysZJ18pwNXSlMDFSb/Qm3LCo2WI7yXlScBx80XRDOenQ
xOrZ2erRBxnxBTVQfKRywDuEbvQ5p/MC08cQe9UvExroHdJkDBFrZATiExbP1Zvm
NXtX4ahDncAhjFj7JAjMcurm7wPUQRhpaI9SMkjyXfVMcHtPBqAiKkzDABSdTeWg
nxtlUcQv1qt+Dw9JtXKr64+LMaaYnrPM6X/+Cwy8N1ICe8AturU0qB5ONeNKDpVd
7G8BjUNYS9k+vRoK6Ahd66hQKgLiGhB6XB9rP4NvSTeTygQHBXwkgdRX6iZGlqAD
EWcBJpiIyBNyg6qV8hcfN/2xutLURANh1JKlqw4HHIswFT6ELiTnYLEqVXzduCSU
mfFlfIMF9vC3GKl2YpMRI868nQSVjFkkp2n+wPP2X44tKrZMZh29qWC7QEmoNKf3
HNA1SdhKjEAqrCQkr4MT2iEwbtKTVzCr5gRhNOFyOmW9GfEhQnVHDFpLGnhavqT5
WAh2FzcK+gDk34me70w6CMHR92KV7oydiSJXm5gc0gFQvYc34u8pTGWee4cb0HtB
D23zqlGf+iPS37Ow48osIHzSSv854zE+1fUzD7dLhd1qhNiqftMjQS/R3Xirudqi
OSXuK4LMmYLBLA9pvRf7+3J9ZRo+C7m4iyGTuyTnymTm5VNpsdWrnLuWLC8sLzQI
9OkyhKWZ4MSEBVbrD6g7Y1OIVPm/VHAtt06z+h7QJHxVDarICj91B6VShWmEum+2
KToEqFx1IC8NMMdMT3G7WHSjTMOTm/mTa9XFUlmJaCJu3u6KyRvl1uTd/IcHGivn
0xQK+9hjuNQwVrvtN8WE9nozAXMY81BL9Moh4y3KWGBSmewk0EUY1F+qGiigbSBF
HoqLKvpqydPSkn3ZTHzdsVCDoabKgowwtM/Wz+3RczNSVT2ZYb+dtkNoYL2beKJd
/oHud0fszMbWmDrSuLylIJoSyxDYhBF6ppnrGAm3U16VAo5uxRyHQ/mvazWnCmja
S2h7HoBNNYAOo+xOoFew2OrgSyCmFI1KnlEBbQ9sPM9spaFZGGpd6vkT6T4QM4FT
fjwjqX7TaTAC9dMKjbTOcogAO8c8J0suSkmQci2V16CQg864fLWvgQN+HHQMYwQK
sKrEndIRF4AIAbAIDDUkg1EI4vaG1rhzLkpRJL57KgMOk8LkCoyhq9z6Cqv235rL
DVvHrWc4xAiwivW69u9Zfkexykyjuhxt9i9xHfNWDlC9qx/5P9WbkanScO45uuNe
MYOZWCNIJ/KfproqR3lufHGwn/06lfnqePud7bfUB25kEdJFzrI2oevG1Iqve7hS
6Vjh70KCPxnHmMl2rOXMDHbimg8OtAnZV9ts9b+IYdmrIW8UnyQHWKtZa2F4JRnI
oR7hgKeybwKwhre0QGHVo9wUZYthK2IIdchhUSh67saR9Dv9GYOE7gfWgoSzy1o+
XuDN8kXnvpTzZvjVLgWiDBqpK+mLBOozIAl4keW7f0DKEfxg0imB/sz0KYOP/OZG
LV1hd5yuMqYTCmMlCT+dd3Hawf5AdZQfb1ziICRawd0UxDHIP1SHQW8Stlk5oCFe
Dw3XdTMGs8QUqm632rZCLixo5KIVs8dn0xf0oAFuXf/gJK1FghcsSt9lGo75XQ58
RANXFd8JmsgB6lSi372DhYKYxZ9ihBAvsj8+99BBpnHPoA8KeWz9TzZo5rg1bo01
aoYNQvlKw8ankb1vTMCL8pvHousOlDt8LzEcq4IM4ecXo4QfyFsBtoVR4R6PTtON
KKHmjhrC0x7lp5v91Fm3dbogBYrDtSRiCappi8Ks06MmpHYyp9FtrOcfYsgpX00N
gUu45JfQlEiCaPNZil8YI7zvwE06g41p+9yXUzLasKBjBBBfOBPTsJQt7YrTxxSe
2k7fFl33o+vswPClUsKqhJyUv2XdR9BpR0Z4DoTM5kEe6DBXpFq05uSe1QNxSjzY
lWFiT2nGGlpp/0MV6xrNfBIyNRC76Om51GhkqjrZHHr5eetsIq3LuDSormBHWJ4R
anKPzaWa5GYE/H80dwYhStE8zkYRkbs0WkGA62o4OqQQkohQ0im572xgfrNsZ17x
0fdjjWkShw8F9KErlqNBg0v/KW19srDXHpA4+GgTBsv34nb39GpgDaiISMM6nQAH
zQBuI57uP/rp40FhV/Ft6ykCwkqrBnsZofTX7tQeV2X2Vtu4bejxJqQfz/Zv8sn5
LfWDWxxOcbDcX8Ar4WLMo3RV0kYjbzTMeDj97elhG1IDsT14oDUEOUZqP4q5atnF
6LQOm1TIRb8FqWM/Cj8wkZckL/PXf4bMcWa/rq0eduycwG0k5JQ/FeYcZINNIBP/
Q9+CI2U2fqJ2KEjG0uE2/Owevsz4KGYWN6m4sIWYpYLhFLbRJI8UGw0dmxI8BEaT
Ncb46eN62qAbPyrNbH61BR/va25Vs2quOOZYm0vZqIKQk2fjZwUyL3focql6be++
BklbJQ0nWR0z0KCCR4RoHofIqt/GYoaHNxYU++nfnfBDUKjUSFA06TaVX1UrwFx5
cEFHeyqI353y6z7KGXwyENbZajhbxA+wKH2y52IwPPXXYUpa5L21OUXJkEhUrZbA
+o1RIJaE7g4ybpifvZ/8NUphnquufl3vFlCnJctFy0efKT/TzfV214Z0/zJ9JvJH
MSR4ZOn9Hyi5L5BO7o5FuZGA4GeLfSeEz28W2pUSHjRrmYTsq4Kk5G+ttR/gT1/3
BuIvh46t0NFM0uXhWXmPG9S99DXMWE7Yz2dNoAskFFbeK6007gHGAGXiLNkwHTAF
BbgyYaIkdH3NjQi1inJZQjQ/ll9Hj5K9tFaHwxt7PUjq578JnPPSMOcWl1cHEPQl
z/dx0JVOtal899lfWfz1GAUfsxrZ5/Q64kf6ydHUJy6w8RxMh9DH9/sxXfyzX89/
SzylgVfp4aigSt7+wDQi2srNEPSF4BLhS7fWWjTcsw0fksFF1/CItKgS1m/yDYTr
iiHZ/KLPYj4yb3M2k/QVueOLzO0mKTFikjRhpJSkwCxy8qskchFuZge1NRiflQoK
aa59vSLwpYbXgUlgs4lpoBgGvb9JaBd5TNDGxiaiH1tIrItyF8z7q1521ItjJ1SI
K+sH5vl48TPi/rKqx0eB0BVhsWPhZnvk65leIkvPr2BSlhwR+8Xbw1e/HmdNGjjv
HuCxPKENeJrTKPOJb/GHW/ICSXXMdkVFfcnrSKNL0amGARD0pYRAW0F62HQse7Bq
OPmfhVOkYBPo+P7L5tOtzMkui/E+FGB/2uW2X8rEUDjHTf9nfAmwppI9wUV4IMQL
05treY2YyTaC2O/DablsVG/QrVf2SNY8lZS+5YZTLgpA/Yoain5BVdpHnJA9edqf
TXwAOxlbkmojyawIVPuapoOoKMGHbr2lTAg5tWJxpqb2kEZIZlxLstIx+iyCE7Dk
/GX/knygbqimxPNn6fmdpH/4vdexlGTsWVrtsvggaG71oNvcNqFABmY78hBAZWwi
CNqyDPKO/g4hzvebLcumzLQnSfunkw428EPvJEjbQCUyUcX+peNlM9CvqYXtHBRT
ig1jvRrmJvp6gYaNqykt/6sBAu2Vdo3HzWOqey3OOUksB/SvxlJ05TCJSb6IYTeg
pmVy0EgBhxZcFmv6z0UDYVBl1Rv9qlkEqGkPWumK5kelKj0RlWUvsK1oXb38BSQR
g2CzG7diZ6FkNnXyk3mtQbNikg4Zpn/kBXbygt/PNntGnrhRhVnOKs+djhioZsAD
KLkgWfvveRDG1kGriOBbg9pKPy5gXxvysbGOHrmRtiqyR3B6IMUmVrztd/uD3k1d
i1cez+tklqsZOgiH9z+GkMfcgxdcNPOQQ88h+doJ/2YYFTjDwxztlifWKr0Ikuke
cr/isFqNUInZwG9jObnAyB5ZSMoN2Xe24+KiQ+4eQh6c16i/qXf/PTythnB4yV+8
gLFaKH3GyIS04r09+gsYJWLUcdTrxcICDJmRIxYY1Z66C1F17MS+gKP9KbTzjEme
CfIw4aEgnRKG7TH/wDp+fdrfpPyfLCJbi9fR3rM8wqx79s+lXuGtJ2LLOw4+lI4g
pBhYn2Lx5/W77YZxQDl5sEsKN5qlCdenupcZDtvwQfc56UXFWJMYAv4SwG7POiPR
j/ZHDO554d4Fcm3GM+FuB/4AEq8RIq2tLVB/ckUv+dVDiTQonyKMVh3mKVUnEFsI
YGKTGlHDabLPLqJbxPFt4fmq9MHJtQ0GiZ9uSvw+ZZjMRZtJ8u7R3wleLNGlb/0u
Gg/urt9ES9f27kdsRYIqyz3ziKVWi18jp6e92cUuXSAbJMjq+LhGW9IqpriX3Z4f
uj3vrXBuMstkMQ/jPwGYP/mWqb+O8SQKE1o6unBGYbPQsiW56Agu8xLVFA48THNZ
i/hPVxb6PC7pKZhZ1Q3kDX9p9WQAY7xYJpDkpxdkj7RQJ+SnQk45l7nOddc9GhDo
yGV9/wRf1d2eHjED19uNztTpgPmUUj0k6y9HV6QhTgs37/mA1qmxBlIL00WKI5dO
yinedgqHLxQLMu2o4BfqIQDiLPBZfaL8ucZM4OwPiMsnsB9v1NdbtWYyrgRVtDwO
RgVZK9qoTWmPftzLeH/cDvX/Ti27JZe5gkNCnXNP3YzbGSftS6c7f2uLm0RyspZo
8uvuC1swWLIucTKUTorwYSrE2HmoeLNDObtvkRToqI/Dzqs1fWU8xJDIO0A3ivyM
nXSZaRdrzVOaQ4plRS65HEnuqyDIsndcb1wZiK7jKN+Im0RH3WdCIb/F8qBwSxXH
rnyprHveEuoDFHsyR6WPJSvNJi/gKQsVN25De8WRqyiW/L06clijOB4Klp21/8aK
/JKUGkxJesz5auqyEOYwdqJjkG6hvH+T4iRIormqbn+XIstuUrZgo2OrmwZ3T6Zv
vLKsbB+9zY8lf1/3KftyXfY8KtCPF39ngkbayY6SIG6XvNdcjwU2vJXE3LEkgO8v
3E6WJ23reFPaIijVUiYMVZr07QoL/aOqxwNVhhH3YjCG2V1JyuY4cpy547ta1gkX
E9MXtM5XcWDbUzgUC2Iav/AxhnhGW6NphfpB4KCF3yiagJYKhf85Y86B2K8OaRoN
l/u/j7juB5UcIQpZhwrwu+8JQqjGM8O4RcDk+nT8qoJa323WXr0pc8NR8W3PtKJ/
zi4hITakrEU1t1GrNTO4qqJNuos9OhX/R8JrXSa2fHKgWH2GePJPiOjG63veO8y0
0Lhnwl41NHRKl6KfZwLZdnDTf/yxaFyVLU1wxCnqNVRbOo6Y6Fl3R026Id+NXjxI
0AGBAoIpHJRtXMWW7W3SjToS9cFqcwTiSKlzO+XFM9SGaFyn+8RupAzd2g8tayNT
7YzKBcEOmJULC8R+zgaATo6XtLN7Q2wyAraA0exsou1CwUFAy1AahmFq0nx6rL+m
nU3AGfMtn/INQD79sy6NmZbRXxRw/ABrE3itiPv7KJLo4wejRgXj2T67G82ZGlER
V3d/IWU3Zr95/wxAV6fPUSi9v5G8WY4lVed3CyjuROnDnvDMyVVTU8Q5AGdbr+42
sZ70iHOituen9CUXWDoYblnuWouRQs3kJV0zvMmhfpbf816eZGZDMGatP/HpUVCh
h8qaWP7ejKY63NwsFx09XBGEmxOe6kI0n1p/er8gipecsHAeSx3ap7GJRIelEkDN
iHB2yn0KW31V4W3poz1jQPNsGW9z19HplTsnfDz2ZsyShav9KJI1bG3LsVrtOnPs
rW+2v5Y1l+Ptr7yvhPe2u8zjQi3BMyIKlbQXA9C5yApPzWO85vfU79viSh0zNHn9
nbfai8l008F9dqMz4ZcShl0pdFzpVyCciil0H1ZfuSxtmJhsEXfpLgX0QntzyEEc
ndFXD9H/eSHmqzmVpCV0orS0Pu7HcjOHpuqyo/1f2Jgm4qvUEf0eZt5fFVGCmjz8
oGdyiFhz1pVapBCtNzm0b2de/fu334ckurjCQ++5d4fNv9/noXH5ypnFSd7Z0SPI
y9abDuX3N6lddQnPxCHrGjt6KKXet9FfnxIN9xIsAa45ZlqOwhOnnbaTZd5rkLMO
Ul4PwrxVArLBzh15bO8BXzmMupCxN1YYSdAoRball4JanbmiDwr5U18Sdo5T81LR
gpHhnhhuNHgqbo0+2Usj/6xaAQyNPxAR/7BEtD2l48nsK3xjvcvdGjRB0QpO5cGb
L9t2OoUEYErpYG83Cj820sOj1ScERGE+eetHhbOtsBTCBQhqqjkvvvEUNQ9rIkF2
eF3S71ISAxOJbXRTLArYuDluLnDPSf0+5IXleL5CZb/XxWZodMBsFoDDKabKDV0s
hY4eTKsEqxFq7+emROLJ/QtsOADv+jOxCwPmXcmrk3L39qNyr1gG+nnDcPdE+5wI
Te80+XkyYt4AEJ+YMHEBxgiKBIdWJ/Px6IY/Pwbd1ZzN39t6MuzU/DbOLS9j9P9y
PyOUHki2ODeVNwetoBo0acyy+2hwNPM3y5xz2MgYUGma/ASOjSd02sQjuywUURvk
3nQ2ChiF+IKs7lSlxP0KCFvY4KYYRvQ6Thlz4gTXEzNh4eU1TbBtp1MP6NrHHhHB
va48YDJLO6GA+ruH+w0glNzinP0AVR7TwSIg6XCLpYY2Q+51TQupTOaXHOKFJ5e1
HfHa1sOkuatomjd52dTaD/d/HiKEteLlUM2UJ9FlTzn1KHgGbHn5LJGgOLwIPT7+
qAabbXPkwNB3xPmPfaVsaZv5bomAB+9UbsyiSI4gLmNDSMKg0YaBaISL+Yptoc6B
kNDogBbo9LpKHoOHiJu9/WAkbXVk5E7sfNMaYZp3/8C4Bs9T1kWuFU3w2ZPARDMf
RDqhAsDEVfm/gleSJzgm8xN3F8QCiAmIrZ4vlPbPaI9sh1bCcKJt2apiozeoKMXF
4UzU/5dnBG2SQAJiWp6hwrALCnm7lJr5mPq/e+g5hkL13+YFmMAPF7juuIx1dkte
ftbLZYV6OgXcLPvky/5Xou1pnjb6Sfns6bTnC25d9Pkp2cMQBfMV0T5l2jt4Ds4I
AqsMtKB4kv3vnGRLbWtIiJjouJxyfYUgg/iONxzJFR5fNaePm3rr7nDOMK+GEnd5
LsJHmFHTeoLonTeCZicjjf4obdOlqCUJR1anFLu4tnTWjRm0UUlFEKYyeKANW/oU
tduIkW6OdA3EokNrDOLjbq3EfL+fu5pXeNfSXQUwBc6bz0cS5zVNr0FLYNtCUbdn
MJoqVCmlRMcejMlxhoELbEl+ZK+XkX3sWSY9W66lh4uZEhCQ6Ezzut73fOz8uPnD
wr2fP+eB7euBPsg6m12aRnvxqoO7VFhrZf2OBrPXKD5vMXn84H7RgiY8dFm35J4a
Pj4uvO6fJeV/PmbgVP/9q4tP4eyct0jImT1W7OYDWd2TAA2X8LNWkqwjLD6DOSbr
B5+IA9WabmrJYu7ySqjXiiAwozXtrpd490TSVXuLyQAkTteV//+Y+Xvz/ojsq+62
VUWmIi6Hjq9ZLF070HT0h7m4WMOf66nh/gX6W5bXKQyJAkgDJlLWaDd/IvtB7eqB
H11ZUxgvCRmZK6u6xpLqSRTx7e9V15zJnEjUk9qQWbleV4/L5U0qmzh5rcyH9Q8n
lv48SKqZJLZntHiAjB5JxOhJtG29QX+4w9nKGdj6OPEgMQdZy0WIN3Teh3k2dpAI
Q5HJb/vLNU9yyo3slAiEJvlSugV0EBjuZAS3r2xtRaRjGb13zRhtbtX1YNTQjyue
pOkSKrjTCl8T5werFXJRt4914S2i/cwqr1J0niED9SuhUGbF56pOFUKV6I1X+oS2
9qpmBkRqRvLbUy5fyHW54OnYU7wCWgqlEsr3ovJSy8R968dmd4CR4O1+5euIb/Q9
pWKHPKj8hzEeXQVW6z4ywkNukoHBX72pjB4tKJQ3uRotQPlEwUFh4yms3bPLS3oV
JNVE2smAUYmgor8llLFxb8ISg5NA2nMLY0W0BAzL/gUEII0o4iwOF+TnMb2ojWZ+
d2sRqSGDItaWAWR1jENSGy4v2m3He0cWd1BZmqCq1T5o2Ksyd97MwJ2fRQD5btXc
AenhZPDTi+pfrtQjCKYYpmc0imcFk/bEerMinUuG2/sGUBFUlpGHWjpCBqACTTF9
QGSLkwmJqrRZJow3B86cQgpRXsfqzlf0TboyjWtoSg/fwe7VVn54EDnlGx2PJI+O
t5b9kPgJS/lXf6NBDcDu63K6XMOwwOPGZEBbf3lQfNNQTuWTZKStfxFixReiuZMY
XQoIQdvuDPsDD+R1E+EZ3cepcEinEyzCQc1SnqZ+SpK/IxdBWVdomgGeE3EiIPjc
O0p3+3SGplQRnRwNnYjQI5tn/5tskdUXsFBz+mAgA5kKpyWW6+nqp7HK7LTlr7Zg
aBtKZ8uKJSHdlVgutzr6k0ry+NqeqrPlW0hzT9jSLfZrnhX651SEVVaAIEAi5SBk
DPYNcAQh7QoQkpV/ddhof58HIZT44WrDna8M73MUqPg8q0ozvf6/PCKJ5ZUI/478
dwztGpxkVj6XOiprM8kJWa60k1ET7tSQhfloPIlkU0Ap+YpONUcp8AGEJs+XSOCK
1vCRsRbv588aynJL/v27zYfWc5/eontKDqTYaGj7KrcsI93NKvhSVgub654VusqW
TQaiGb7j5tNz/mS2s0904tpAMu/LyMuz+hU8AolZmnH6dFjvsovTGPLuQeyQ3rGj
R8VmewWARffqEFZ6VJdqdj0Pl2DRFzrL1xvRxaS6rQDjfoIg0kvMLCTTCrm2SdV2
IWX6CcgMSMpiy1PfAnfTvdMJi6Gb+CE6HH94Exyu9bT39QCmD+49UzRxKoBqUNP3
E69Ef6JXMysHbAnZLwSTB3LIvLe62F9PpFCtLGo9PPOAk71aB2UYQxD7w+CJq6NJ
BqYFP7nUpAkx7hOYpjxzT/jlF7L0EqptsiQ+SsqSBw0E8kWoPyZL/xKqU0lLLEdb
jJxH2xVoMP03X/xAwVsNPNmCcVetZW1SNjz921j+nZEgZTikyK5HmCt1JXs2zTUv
p4kQbY+bGC2bpDJalnDIhsIWPjrZY2ykg0wvISOlMkvARulyd4IwZ3QKHfki1PIy
jpHDf88KdLKlKiTippeSxv2zpGdBT1P1kvjE1/a7JDUXQ7oiwC1nxa1tISTsmB1x
Sgqz8EETCmPB1oqu/nMbx/IZNdFnWBJa8lhFaWj/ub9w7iuxiRbxuBO1OqkCMg7Z
u1bYIwWR8defjefSmJTVle4Ettp7KbkYnmwEC7ifLqJsyvqiJRrkT/Em9XkpjlsQ
knB9UQYdpNdtsmxFGF9TTJwa8P31ziPjqDQCYxpCkGIwc2YnTpOh5hL2z+ynX8WB
HaooUBEAJjh7Cf1cObWl1jcgCEDYcBreBFrZTq9McB4tncErAeiXIj6gdMRbwqAX
Jaz394mGyJZ1B7IGN3GGIxky2NVY68j2SXpfyVxsO/5lVbKjcYMSTZYcyihse+5L
2QLk8zvrULlhK5ELbRwmg0AMQHQMta1HpQaYG6F31PmZoDTDLYdRI6SpME0YNTFd
AmR+hNImGuLvFkFthdAzcKebzJN/ZgvRshff0IY40gcRAIFsAyKL035Gt78wnBM0
H8GdkUU+op4x81DHe3XDe2yC6qtNgTwZq+KETXGrgTsY6pWsrCXOH3kB1kZLeRqY
65XKX7+SdTgp/bpCSMIwAPTCLXT6t+khlPuHt0pXYOvlvVaAPehwQUPUkkN2T3/b
QaguY3hziCtK7V/kQcZpQ5bdHEKU/xtOVg0nDY15p42FhKE89RX+8u0J2QW3A+xN
xJahxvmKwiMSQ+oI2nHkCA+p4ouNlFTf1Ztkj46IqczcGbyr8jWatRblpA9xgj04
CZD3VSBB9Eh9JteLTUKLnAZBqiGSRezZpIlUKRICTS+8U1QIoDe/9T4IGPGS9m71
BympqwuKmbQ4Tldohrz/m0hU3XjXC/NJUOUkYAkqCKEjsSsiYcme5iNIpQvW3J71
a5nvZUihqDHNxOfUnl6p8DjEt7c3DLdX7Lg86vCe+bvoTStoQR5sGSmrwO/V1lDR
gdGCYSEi4+Hvyh3sIjFpGLxNtlGnaYbnmgq9VYoT93sjKeshE4sLGwvY0pSM5Azd
+VX3Q9OypM2pSva6ZwQmJXwjVGKxr1/ty7flrM+22QzDPda+XeUTDPkiaYyI3/ZK
ujY7kHU275J37zwTqu55dzuQEABTzBjfQdDaB6pgY/Uxp9Y0cS4teao4cDgxANHW
qLC4HSzbNQJHzir4YB3ZHEp2ehDyu9l3DBnSSsb8Bnma9zghc6RU/BWu6WnhyThu
5aacwvFxz/o2j2gTJM2hi6CtTQUCewjonpgaORp0FwTH2cU071tTYQHE5xT1Wl7n
/MGLvirZ9OPeoL/MEGwJcwiV97G35fH7tzbt4rRxQvEdX7NfUmlSuZLQWzs52/Hx
sX9uqSZe6vjpshL/FmbefpzIlFxZ55I833lyuZ0vteGwZXxSOaN5lQAOoNt7MNaZ
LoeO0kLzbx5bglf1GCKCqk0qcMqycd6im3wUcxqCjfptRlPQbvR1/cuOS36/CjCR
ur8967HyrC3s/eH+vPtEr5VUxCyYj8quqo6ntt1omi3v1RRo1ajGti0w8xNVKKL4
wKyJXtWoBxFMF4z90fBjRAX1bH//9IqoeO1dVzu/Ygc0qBSPgpkWwKPijtQ/Ofyv
HWWdkc8jBqhmpW+XDJwygYaI/xiM7GigbJMoR7wmYK5M0rq1VAX1A6zQcKrRW0QL
n8kC1tOPuaCq/y5IvtnmwRP47/nxOF+wGCmLMn6T7sjTrPribs03HfYmTkysrY/N
BdLEPMV7w2TvCEVu2iMYgeP9h7F2XyTtP2V6Rc3FYBZwp+x6ILb3YD4fqAEtunKy
yDewdkmPunZ/iOT0SIztCGUiT+4dhYl1g2oKZ+drq/VErAR+KxMMPlm4+AiClaw7
lnXWF8XGSo+1VZOcMon9L82m2eFPjT9n46lrpVp8NcgFXWu2Qix0yakN4trkgsV4
j/O2SaFkn+6k7ZFALp5JG7WW6+tdCp2O8EHjPkHRXyDih5kfaviY1IQ/oIVcZPdq
sdwNXEywm8Z9MOAgUVKbClROStIln0dy+UCPi6rqFV5bMFlGu1QiBOt8moFY32xp
EcqmsVqnqjDn4TT1vHc+216hi0A9CVb/zdTz6xkEUGSxI4/M/f0NNfm9QuXsTeWp
SnEbjgmyvDh3JOlkxMhUKQ0D2B3sjFx0719krYc1vhXs0nvr3s5g6Ru6ERG/PqMk
asLTUniQaJhP5z++GinkZ57eJ351Y9kdVaNEY8UDKqKFn6VUME6DtGup3ADmoC1Q
Q7GlnYBzwU0kug75lpGfRJsjStFzmgITXUlkvnu9siXk/964OxJNBfbDCwRIAL/F
bQ8qeaC2jbENhdExJI+ZOVCqCqGTBEpcurKV7ccNFwy7QuwuEmapXL2EdZAXMT63
2n8mue/ASgd3pqqNVJUsli15eXshEyFky8HJBmBRIOz+gwHMGJMUzk45ynshVvkZ
dgWGmIlJIJjaypQW96pl6JFwjlXyd64K3jxHhX4iY31QBVZJokCfuhKi3irgXhG3
U0dHcDqdJMgVqs2D0LjenNH3q0ZxlgSuy8xal2s31jtNtSXoUnimM7AgEG8lg0yQ
s19G2zBjOKa5dt6qE2pETftP1rlxIhGVW/DXzKX7azFM2vk3Jcde1ENeoHe9+8y3
xHWRLCh9cb0J4ZV5jQe5a2XA6sQRMKCo7MJSp7mJcNNLuEGNRf1yxgjbwgwxzd1K
Ajr2c+8CduM8iIOdnjcEeHhjdHfyxVGwLeRfKQ/eB6/7mJiKjCery5utr7N1YH2a
YH9pK5cVgiMkU9yibKrea2ssjrm/1PsupVupLsIBug4x7mIqsWGMvhN6PcxDXnLd
fA1cfUYIkcpcIYQwN0O08DL3t28aEzFVi3/0iUPSY05qjP47CYy6EbPjK76ux8MK
08xSWyOwyc8jFqA+E05YHGrQ6yPpAdqji4rK9y4LuTSPKMry3ATeRLldraWQ4bCh
RiOEzBum9x9eZRNV3K/q2S6qL9PeBhstbRlQXSHoI6ot98uVfqPwspr5zJ3pBcQ7
48VdULxbR37+MumdH14Pe5oFzFXvXilFgeMXVLgAAMdU6W4/6bXG/+EgB8Zj/jX+
BSU3D8n8rSJDP9yczCCn1MHmxEj748mjljVZDczGJTzln6D+ksnqfXmoUE5/Hs0I
dVg8FFSrr8a8bm8T8q6qGgy+lt3Upv8YHCjGxGujtVISPDy10kHO7wonicCALqXr
z/oLhAqh0ztGX9Uo+jTloalikQjRi41JadFNwAFer3jlQMtJzSYAfgqe+okYv+h3
PHHLKwNATz1ig80pEE56/WQr/cWKT0Cnb0xxxXQUbUakIwBC0wvgSqysp7Rz3dBh
sCU7X8v8p9xIhH08MsI++tvUtgjYy6aIQBbHN/ZHvLBC0jSoef1HrL74F4PUHgvt
bJPzCn68vFlK/05qlgrsIlFNOnb94KoY8uosgVtAkx/ZlK+TXx6lnSXGEKilp1/x
6J8LGQxbuyZ7+7HRTvHzjnR+aQvuCcipPbfJs8kGP4/vwxYDWSV4ad6jnJc4c4iy
Dpdtp7HGqL65W/Pfpffye+Kwh8PoIk63c3cl2kTihvnUHFXubQ2nEd3tFh0Cryl3
FE2z67L2y3/7lmGpQagFsNGbuqPbE8F/F4ii5561pCN0Bkbh/GlJa4hm/N10amHj
60RhJ9Vyk8/t9rp62LRaKhJFlhWmp+hKBc5uhNUAf47IIZDg7GoFxTwlz02Gzo8L
stvadc10brzj3QgevW0XoBHiz/WZ4BbTu2aH6LEdSfd8G1Sbt/iSWMrCKMEyMwhJ
STmkFhNRtun4rjMWB2U7HC4dmNfA/tpIFNf03SwQWK8NVcvkuIMY0/kICIOrnAVB
QbW+8yhUkPQrglEqOCrJXm5nWHp6jqmnczrReq8iXKH+Wc0MICa6L6yE8yIzD+cb
F2tdQzChq95aWAyfOFfSLWds2AV2I4oWKgOnX0amWnSE6Iw/bWUBdc/TPgIaskOx
lMkPyzXCdTx1JYEMgOWKZ/qu5DgsBsQU9lOC7jDeQQDi4+FaziJscBMPni4IkhFL
qTzgdu2329FzUDd4HdDSnxkAWyAUgP1XAXNAOIuVyI0EnTSd5JIrch5B1KLNcV4a
Ft0HcaSoeKuL8CFMFpO5rlJzuSUqkBjLiNXqUXcxFGVsV5NFXU4kOIT6WanrRtbW
pufz1Lm/3NCglcl+PYOXwGm7Jjuhd9ABjjJ77bh48Ie5SNM0UUPxPGIiV3ToDE4n
CQSX2wg/n5EYywOzJW4cjgUpphtARjxCiiN+rTrB0VowPpwnhnOB61AZIE+l+oHA
B1D2moVPFxG2VFQJIpdZ2F3DtTy2XMXI6/P5SBLdmO2LRlqjgyQtemI4m8vpej4+
vC2uG+jbUyWo/GnNZWvtvNlNu7FJxjJjIxbJ9oBvyziTV0iPwg24ixhI8Ro8EtJc
fv5yMfRuF1pINGUxhoFcPf8YWf42L1SdQ8uRrrQLKp6vZEVTH1ddGfGtdA16b/tJ
2fIjNoe6dWGErvLtrDTwEZRmM0gnfeS0eQ8iHEDUMoyqZbPLWXpc1/VtJQxxF3HV
n4rJ72v8x+BMG5cmFJkR8HRjJqHhrpBtJMNMqUzw3kzK+8NlTfFlxZwhQWrJSf+o
pP7WDmDzT4+n6J+NilCp5A3Y5EPr4+QV4/NdrFcuQG7Bn4hafY3fJC6h0KqNGh8o
1LuVouSvw9BmV3zNMSg2jJQsJGIM9GKhDUQ+c+Ediad7za7bIMeh0E3SO7UJ6ulc
GrtV3LMioBJtikoCanQSoljSK1tYhr5/43QT8ODgfRu2PRho/TysSEQnSVL4dBoF
TBFfl2NQdmLId9HJTmVycELTH/RhmRe+pIbqPShMPsPoXzbyuo/RwXk6QkhP/sEE
0b1aKBqX1Bl5IRmKQmC2ESRQYjFZOt1ZQ6Pm8TEq9PuYtMvG5KANW1eMJBqRBEsx
R/X4bh6x6J8jCBzR2VCmXfqIV2+TXezpmi8rv02dvt7AIsgZvnsMq3FxHqJr+zpq
3woSewVnaQUDBH5fdNz/xERAyzFRu8pR471l1ctgkl6Ti1HXqW7Mw8plmAH52Qb0
0BZdNGDvVU1V/sNbU/C+fzdpfNQGVYvClzXnB+E9XvAzQQAx1c4SPMzNGQUmEljE
r4Mh05xi3LdVjnZ5D2HV0lfduIetucUlY7aUIMDxjXeqrb6nqBqiaXDn1Kbb/4g5
48EDDPLWLSypOXZB+Apdf0xpy8zxMNXkr41j7HbSlTgi70TNQHwcKxppBeWYTQ34
viGLUwCEA4g38IkN/MI13z/ucewJeqKHfvoPJyioHwZath/5n4v8kE05jXLKMYGw
EzGQV9Lqm3Jyy8ZRC2AyUu3q/Bu1628zwjnDbYLq1zp0v0IRJbOk6afdQco9T8J1
7zUnXzdFMqkOfB9KHsF5oJ5mn+Dy3ciluteW95nKsCvExnVqFYtRE39hFEtmIu0t
YR9o9UJJA1b6Fld3+4UjYGSRVOTveuzeHPVBtRyBjWFIlGXl6cQvjbselq3QD1fQ
kCjixquqnvphMS+GN9ISoIjyGzFSoAiIM090TzC6+nlQvbGRluhreSxMB5ck86Mu
WCRiE4vsXl4wZY2fPTOVtdK+2xRTTVSPy1tGOZn9hBbnOvPXmJNJOPGEHdHnsmQi
yA3qke6wLOO4NViav49VAXmL3i81+GVYJY/CnshxzBEWX/Op8CEayHRHXRL7wjMi
2uyTAKdaJZNmyEbAXwZY+EeqNOZsOYu4WhEhUb8Ant06Qvodkn6YfxtvG/B3izFc
wasktqNbsTmWwBJFHL6bjGszyWq/RwgFC/Siz4y54ja2AswyW9c1NaniWt1cYaz/
HQsyVUrF37BeaCIWDdoqJWmPLNkPofISxVLgD5CRcOv5jbmg/oroGuZmwRaF+dDI
bTRS6CxrdAgkN2aoUXyBnLK8BNPp0Djc8bLs/TCnyhMspaTMm/ykRWLXp+OiHDU7
ZgLtMpvt6h2jbcqHHVcqlG1U2I6TaRin/bAJFf94I3frgjULH42HtfKNB7j38JLW
6Vjg0/G+q+6yW2BMGEQPclDuGLDjOKgsrsxHUnLXKhzjEYlJO5WEPQITjRm/ZOlR
A2xpcivMf9+6VbQ13rt5LwfYcUXT3jPrdZx9fV9M9VH4/i8BePUVn8pnNzSttrLO
G6+bHLLrnebWWefHdgXc1WXoZUl2UfNrTquslzBqq7CIuxcASOmlf7//fgbtB4sA
hknNkKfVEiUpI/WQy0se/t9FFfITy3g9M2+FWweQTiXRp+mbEMfINcS53x2M4agE
c72crRZ+/TMk9art9CMIYevGVoqk6494gaTPeY2UoFnzlGJIIxwojA8w9y9ZFyto
AQnkO57UUtF1/WgHcK+AQHGCBPDEc9kGbG+hBnkW+wMZ20FTKIsSPOyG3aKQ9aOI
XrtH5tY4O1t9T1YvOtLZ7gUrlpuw+051o3MbgJJ9aiMnj8Vdri0fiWMVcf5Hgbzm
VjvkPP1MZAOAYr8dOjC/j60LAXx94bChuXGViegqS/JKv3Q8lZzt7v5DlK1938J2
TwprzP3DH0Cfs4WSGBONjutkyfa2zjU1Izxir6bhFNUlQf30WS7eKLWzLnQF4JmG
xlvq5IUCiTfVm7U5Y/0xkkPC8RU1seOoTLs66ZHsN/jjgacEs+r3wcDY62e/g51Q
l0FwvyxESOx572drJVdAY85YfXdXxXlAnbDLgeAzohcGDkBGZEVk8yUYWDRc8EBz
D+uKkm84AXsLSlOD/HBiL7iUO3tI2xuS13eYi/yM0hVBqIhtgD4J3pidp+B0aV4J
AiZn7xuCuNqV7pfXfTjCPYLSdXQcKcSyOHcCfvcbnVmtJ0uRqTzMbpSWAG3yIvAu
neRgTxgadCbcG7y+DCfIMulH99VoV6nZKK3od7EBZi/GkVzsJEJtP8VljH1MxnOt
+HaevS57drgLWgDG9obSPaVNNysv1m3onGJ1B7nnyTSRJ9SaRmp6Znc1f19aCJSv
PBiTuDryXwGBlZ9O5n2WAQnPjymyeF4tWbJtbf9iLSd4NEDEbgPt4FMbWJw0f0sG
nv5RqYIx5ckJTN/ktKjqn23vxkVHY5oJKbiTS5I8FOGKD4bCC5wp5WT8Zw25TAte
8OD51K9ga4ytdPjMsqIalBa4YcrG3ZYJ3YapHVRrW4QKO/4gLJv9f2bGJXg55zMc
UHIKBir1+5hWSMFbPmYKg7FjcilzvhUcKBMeSrF6aXJ6zqnhtJuiArInKJhB+Rjt
7EbVY151HRC2mh/ueDvXGbsBWM5fYFGX4ZxKufCcq1DHqAd+SOetDq0eZ2h/nOc3
0fSZDpZWMJf0R0+KJEKkSGlbFIt5CvFLbqOSdFyoEOit7PoH2yhMCxNX+wgz+BQf
/h07WA0ePAnwexuQXeL1b38rm2QpcEDazvhLBpithnV1modCCQ6IPGHAD3s053hE
nAp/OLseJro43Mww4KHNF+G11/OOJnBjKPwY5JuNa2U68unmI+H1scKK/qKAccdI
l86fhCh7YE2TdHK0hRDwxBxmqNBR2A2bcQX19xkgRVXR3Q8X1zmkVSetC0dH6pS9
ICpBvzhNGLrLC1ccNuahsklfpEcukH7RtoT2gDJUJAlg4zo1mAKS2hqOcGHPw9zh
EXT5XIcSTVrWtMfYc6a7NyJTcuDyYttFUtuGKsJFxl2ua7FTL0tF/1LSeJOUS5aF
oMGiIU8JG+ctDee6lltZo092aBukY9bbbj+eSqcMoFcuMnC6faKxMtLqGcD3HG0J
ESfrp//P9REQVnyK4EF0l5QoIPYTqhRbMQkE2Be1/73bVavnBqB96OakSbUE9DkX
hhqwtDrx56IF/QuD7NmNTqxMfnzgzOClh6I5Z7OWOYdMxyWlZR2/PLlJYwrMm0my
CimR2Yzn2FuaRF92s+xAyVCgCeAYJRBuXPdSc/fL7u3y2gBL5uzPfaSQHdlrw4SV
bxuWkbeL9dJQUlQAlYLS4hPvdUt/acxuFII9aObIkVpo3ZR0qKLoN7eFtkVHjY/u
UBLDGFSFbv5cQ+Q56ggWvJ6BY+SPVKL92YWcRjesgZnZIIaI13UJCdCqqZczRLTQ
mfIt5+03S4ZyXntDDwvW3sMWqmhTVtkD7SRSrMjmj3MM8qYwqsuyOlE19RZpTa5l
xmMrwixMbXzvUgK1t3Pb5E3D3w5Wsz7kDIW/KW9IxHnOH0ymK4pmqX0dPJU/OOTj
FZmLUruzjZpzyBWlO1PT3HqdBl19zb5Zf1s2OtRx23aCwNR4lF9WykEv3RpqHXx1
LEXs2zKOdnz65Nz9RDx7/9w1CwGC/Gy0AMHxiQ+4izn6cc1Z3KL/zREBwB/7lQeq
KNKHA9ElzfqolXF6i7YwhoLH9n6amdtlDHU1XVR3ksNwyygePlTPde3yF2YJBnSj
SOGZ7Vc97RKp6+dt8vYZdpz8cAYuUU7hOo1P1Ye4Z9sR1ZIjSfgq7WbJ5cWkK9Pd
qbT+I3r60cdHbW1fBEYvvllQdRs6fwOcSbFHvgNPXgasN38ncQQWTVCdMr4v/xxU
RnN15pmvsfaptnI2dpnfVppZY9Ax+V1dUzvysV1ZPmTDIy7JuYbmgie4jfPBh/Fx
JYIEjhRAQcStUrEEihGa4aFd/cZfewZUHGjX3rJeNHAch3n7VJvgOcQ6IRgPdgSr
nXJmViPu7ZbqL8jWwv2VXmXp5vyFtmUpUvf5kOVM6e5PKUwxmrIjV64eyKInbqsx
jCFF0WFzy5/sZZg9H73s7xlFq0X9tfiwo1ZIlXGqeryA6UlWwfNnGBrRprz2jMw6
1UmiiSQGfzZRq/BqO/XrEp4G0LCd1Srb1hB6Ytk8GhnrELTEwjWHAB//XOgyBfBk
BOI5BoXWfcGESXeXlxOcZoE7jIUoFoSHzj5eDS0Lmgb82onKrRK7jhRDQBf2/cbA
6y1szDO+jMnIiOPvOQa+/Tweb7RF7z8csB2uNIojEvT/CkxbYiEGojJrtfiVgjpx
QzoHjuz5nW20M+vQXf1vH0PBPgcMafa8RkJQFJPkeKfqaANfF0m0RX89itI5ghuN
5rpGNfjaYaMMUIAUpDoKOYT40a7sj+z+VdjNIIFrAFhCr/3eXt8aefLcQB/a3h0B
/zGG/mgd+ZYv6cjGwUgPbtIVwRwmFH6p17uCBJgEwHEIkmuKUQ/6Zbi37LKh/5Ky
DCVzLl693SSr+7JAEggtrTywM0eq06px9litbjBvg9uf2ZvQs842cpoaGcLObPkt
+KNq23355fJKDVP1VD9VHt9VFsfU4pxaxjVLqqoOb9M9c2fcRsQavSSEkxcY0TJt
jTIi9S9JutLz96bFK8nJY/2kbuHpAPGJrtWSySwxUAJgUuwb1COjOKqD3epSf7Wa
O71duawDNBd8/wFViavXUfRaxqr9gbM/3+gG1PXczxsUP3y2u7oFHLjXMCvrY1hA
xvqQjT/jIGXktEp6+qyUyekkiqOMMuZV99Yx0nowg3b5f3AUzmgDfEuG4oaTgENi
3H54LoyNAJ3lQh+XuGwAVMoyig61jSMhj0FrGc5WbOjiIrR85oW2hGpGX4sLNfTW
PIiIkeD2pcEkfTmO6v3htk9UkyLnZ4hOpgUhUST4HXTZPERzm3g9K2DsOsbulvl8
30c4DZ1N5VAo3ToDOE8tgT3bjGnFq4Nnit4RthvSucrF9roO1kShb7sfY2yDluPn
sUmQUrt/mxzxOCPx+iwepvaU6Xyn9BGVXZqIf2aUQenadKNabtPj7QtB20rr2iC5
/YcP4D7Yk4J0GYSpdA0t5rnOKq6oNCuTUpZ/uA2oZL2g1fQ14EhI8VrsZyz4vMZH
Zw8bjgcMhO8nFIO/MdY9/mpKBXNiPpjAOeojcTs+Rtj3fSUpN3jSZqMvVFMOxiOV
EG15mmBdEI79+jFo9tC82hbvc6NyzrxPVmgBxY+ir7LZOQd8qlmaBm515jsR/z5u
mDaITJn/4OSfnsFlVbJm0yUEiLbvoZuSphTXt1K3SN8Iz8w5EdKWuDIQoq0JNYy+
pQiytGWMO6SFtbFH5PVn2ULSJvRlfbF39Us+hAEqRermEo0M3SgB4urq+rYi4HKM
adOcb/2zyEMv9JBUYXnP95O7afqpYzD5Qh/h1OW11Eou/IYmNRUOxX3hzUHYOm7s
qcseFshzyy/FEP6LiAWjaBP2TaoNe+AUOJkK3i5+LNYFPraltf0HJxJe4alXEOOL
MPVCFxT7+QUd0QpzISPHHddgH0Ey9yEt4I0NSHdf573aodBEPMo8zuzUNe1zht1a
XOxYC1IFgo7JPBJ8GKG78uBKL1D9VaKLWfqMQSxi36tuqK0U/3eqy0mDiyxr/wpr
fvuYohTTCk6EM47P4F1X1AatbI30D1LS+bSkOcJXHcAyGTK4jefVnGjlyEV3/wEe
aZnlNmcThU+RdJcwYAC0o+/4Ll/Nb258zAfh2lQIo1BqUsOTptyppQQChKaCZ+fC
dTNP8yLLtLkwZm35+aXHN+uSZM6kkUhfS9k3if4KqjD0hk5f3ALbemeOLP7ECfSE
1RQ5KvVZfRtlgy/eFZnaHCQFqBTqmvQs5ZtklNpUg4a2rKay0N1HmCVhACer4Mrb
dwxMeqwjeaFiY52zf5HljVvKZKnnpjsaqoxyKSbv6cu04G4RHKNSFc7eHJ0/GWrX
R/8GT1X79mbC8ApQpqyyzbGAGqAEbH2U2Grm7MNJwopILcsdNgIpxmVXb8kmsBgo
KKwZn8+x92k2BnXmA6IbQz4oSJyN9FZ3wBF1S3mSdmP9Ep89AMcogjq4+v2gbvja
3/rJEbuwA7N3QzrpG97//+T0S5ZAJecRHcG3D7H6eqFeVjaZzEZctt9G+mPsozA8
uZUPlHT2nHw1BisZ1W2bTBM13I0IIAREz9jXhRDworRisXgt80n2G8HdMjEuWdq3
OkE/HZctV+aihh/9V7hogIRkYxFYnYGJ9WbkxDXn2ek3kq34h6GVwwT2tP31rWcN
bBUYqFdyYW+p1VU6lpnPbJc54BxUBE94mNmG4c6gg6MaAtkhrZh+2AP1xh413i+l
S2kGqTw5i/+MCIW/BhBKCL4rz6vr4HtVwNGgi73xR3oeLEAn+IvjSKP4tttC3kAC
Emac3q6Q0Uaf3ytIFczB/nyGcuDMDkk2kOzjW3+RwQM1pD2b0ifAILhlHSjEho1g
UoWfn/pWb6ZNFV/EZaAKkNyfc8nZZ91Ceoaxyzb8Erl9dVsp7CXwvUVmiMyjcf0m
4falPgLxtDBxEmFrWJraS4z6TPtwqW5XfMXFmj41u2vJNXpEuWBMu/dPcgwnAahg
wZW3nFWXgtl0YkFA6sAuWK6PpFFCmgdXYXKv8efIZ5BoZcazOAWS1DFm+uWsVo/M
TJImqTLXtq31Xm9ZOd0ztGlrFeDAT/is3ptC6Oi6g/Za80/NJSCCgUHzwQF+yOhe
jdTIkwui75zcSJ2RFLaebEEeqQrSq/f8HRSQuXxIXEStQZb3ZKhW9/BtwubHblhv
5nY6FcW99RqYEhAeGFaKEPhNLsHuxC5EjUsENIk0HCXUxpEnjJQhZzMtHxheIMAV
9R+Gz4McDiZQ4kmuX87FnQ9atA56inYycmhWPSXEJ4lJNLd7bojWTOhDDDCWRhSP
bOFKfwEw4parpSlugs3dog75dfoWSG0jmREywanl1WEuNw5ibk+NC6aXtWyDBkiK
kniz5JtyvZdGnJft7Kl6R6TFcOlkdS5MFgBHeul0vCyzgssjtwKwI2RMjnV48yOG
Jb6HNuP4Clarc86ZyqA4aFTNke8YJzP/Dfd9An429uFGfqoZSRlewCw7fy05OGCu
j9PT0yUCMBoLt6tZhecJdhLvv6knUPn5YbxwCl/zkIMKC4EhtVbqHXfjUG8xQuRH
OfC+jtqf9uTQSnvm8UT2dxBPZDkemQg0nzPZhFRmAMoPHU/FZ01VD0/fAUMVbSo2
pvqB1AdSKMEQqmG00CbACU/3B0SGLLIgqW56mNvy4IQSE28i+TWNUrPey5jzibmd
LWSVt2Ecpl2EMNW4ayapSGsWomj20LtLdX83vOyOHfConrbDvydEJPbMpSreGt+W
tmcZaH4ScuK+/jQMSxUhgrRHj5DzTsbSdXxru0kVho/Qm7Pp3HWsk5h67ONDJlQp
kq4HwDstgBGlG2QCLJ/R+6/xgLxHb8VbYw4rZ3osf7ISSCvXvUjztCTH4nvfm+Iu
6BTLlcwJadnaNrb7MPnO1+VmMOq1SF3iHi6BnYi16nWVHXxmgHyf2MnlKRobXu8c
aRD+pxPuPlS8f3mHuT/py2K/Od9dan47st8gwaBphNnyzZsbveGWcGYG4fa9QRr6
4q9AdedBDjVEetnn9qb/1qstU2/++WwnANz90D17oHW+Yu3IR5KV9z2JdVP+KkdR
ITIb1Vc7HTEhEKjv/sGMoDsk0ASaQtAlWvZcCOYiD0nQX9p2M4c3i9ACzx0cHabD
DkHmjqYwjIvCVOcQHzlCTMvxg8HeQL94lVhpvYVwhJu/a+7hyXmvkdmQ963r/0q/
eZ2sf/EbAdNOP2zggpqpM7zZpvXTTXGYk2FlBSYynGcxWfWFVLsN3JMeFOgc/WGD
4b2oJrRFkIZsIb+K8jXplyh+hZ+mn5yPjuqHWbIkMpnTM/A9rLJbgpivTsqCcxxh
vTD/Hdh9oUI4OjFPZH9f/V424O4avAKcpU3EBaAbfF7soWtPuXAqFk7CGgcSOdMe
neLfMT5l/VvnNpvE6qY/4GE5sJ0wlWK2wp0nh5XLwkDBTjPv0+nnZcgxBLbsa6WU
dZ8Hi2SSjVOnWg39I9FEeBiXjfN1GB0Ya0wsmBUbw65vf4gP0/oM1F1d51OA1PL4
QmafdIYg/7+h/6knj8Cb4rI6bNNku2apP6dHR8yA6yUeBgwNAftnng0hYSA2oqS+
P8FyT8y0GgE09XZ+Bi6701kzFiLBQcGom3S8DD3PMhbRGKms8uLfZK8H2BDWXyqw
5VFwQGSUbYM8XqJcajWs7sTZer//PFIgLgmo3zc0YohClR6BVDh27iN4KxB5TPgY
OB50g4Gl8xGDQ7KGGEwNEK7ZfKhWlfBPzkP1rQEoMaREd7PaTEobiAfTn+vBzDcQ
HF8uINPuUG8IqYaK6po/1eGrQ/j8qEtKZcKO5Kqmq8WvK6oppVRSFxuLkjpBVvKY
KfotrQF2WVZunzVhXfwoaXYGeMg/KaMzlIeDvp4P4iFN72n9g83rdUJlcN4Y/zS4
6U+0z3b6psdVVHEL6tGVqVCAhrw3ymbpfdYMtIgaoEJYacYFRcHrSt46YEiQShxU
QiGAXaGbL37dvHwPcbSxWGBt7u8er/DRJbeHQcx4Fsfsgmyk/GgZSqbyQEqHkgAq
EiStTjbQQ8eGDPPCnb8+lK/KaoyQ5a95hJWq1otPvEGGtciP1Lto4b5SZ48WpldN
s9+S7CjGl4fBtwYQnZ6NN5Jfh6IAuVdZIHuJWtYI+Tp+d408047hL7V6z/UawKNz
lOaky6nHlZ1e/rYnFgPSr4rERhgPtZ60JpJXfXG/9B6apL00Adh49Eilm81GnPgD
mIGPxP3bnwuzYZ563VLDNt6plZ+xeQBJDpI6yhBIKZfKurfDp49l8pD0tMaFvZVQ
kWfyJ696Nnp0hIZSZhuGL1OWKgQwmXVnBSvHq7nQ4Hacj1c2MsHMNbZB41DOD/FZ
Bk5G71spsJiqF95op02pDNdRh0tVyuGh2O7MYuNEFjcJ4qOcbkJFEMS4O7kRi1on
BINswBVXXBV2goYd0dF2bdgeeQTIU8RebtVT/EbxHr51FT6r0lHKsiY7nR7b1zju
KPmCEXzjeWw2H6QVrZGZFkc3gkoKtpfOC0v3r3TQitqbqIWY1fl5m/oJ/nGJZKNP
vq7oVZ9DPiDK8I/f9vDteM2bLobw4ytgjREV8sTL+aWy3T2UUhmkFPcICz6iOkfa
PAXqKuHwS07jGOR8BPFLNRlTYasPXAeHDLmp/3xoWy+J9WtPZCXs4H3HdDLX6TNs
us8ed/cPPJq/F4rm9CxiDE6mcCDnsOkezu3LGVbixuZB3zbA+dSOBVzkhASiOPYW
9q1P3exlwLf2hdgZsUFEc3XP/rGz80JdqURnexov+CEPUe6xssI27ZLaYgZkUXyJ
RysrpZXfhxEplJxKIO7F5aCq+UO8ehpOhlgmJ4Uku/PdnInWDnxLuvO+xe3QOAQC
avnRvw24Cgv83pKw69mBrJp12mdbaMrK4AyR3si+v5M1EYfW0gKH7Bek7jJ9JH+w
KRoso8JriLseDNM3Qw54k/2PjDGcPClqncUUFlcUk8lLPNra7gtsqli3iEdRtPOv
ROwCSJ7Wcl24tqnox7jJh9Q+agYoKC2xrac7wpoI5g0yDukK3mzOLbVZaFWrpuqX
blEdRkHppIw7OBEJyOPwg41nxEZqg34pVnnmxFdVcjCskAG6H4YkoK/hKtDdeQbo
KUQNKBNSZXMGWS8+33Qc2YI8tDdPnKcbelB2GDwiYGRh/PpW5NLlLOqcuuVlUI7J
PiEA3Yyhv9qfz/3DLpqU7MkmmcrUx/QPsIwuZ1qUtA5dltvo4Zwt+kNdhG+KzMXY
uYsiPsOCsj+s9b+Fqb+JUiyXXnu5vu9xPo3HSBSIr9kvgnl7i5vWESHs5bCVTNmR
JYbvMcApmiBob31SowUZq5Iv/E1+6llALyX8shaf9uR8E+phkKZYEMnfotxN5t2e
PrBg50QxLHUT2IF7UJR+DVS4qfCFg552Z+m9wIdL21WF18CYHdMHEFXkN2kPCqoA
8hgph/cSdTlGyaag0wZErVk4HVA4OHbpO9NVr4CtvtkHn8YUvosF5W7esOR8Op1Y
bZXpxbXRh5IDcycdfzR4SWb5CSg9gMispXgQOw6gVh/iSwTgRfh/IV2AIci+I5GL
qOokbl9OP0dWf3DW9gnzZDXdLlpDG5ktq66p04vtUcJTRtvr/2O7+ebugKO0P1vn
xgTArMULxJWcYHDiY67Zv1RyS6jEQWI28y9O4dtH3flypF2yoozu2pzCvb5LqfKq
sxLis/wOhNZdO5j91geFkZxddv+TA1g/rYOeZlI2ILkvh/LpbwGXPePN2xBvuqGq
5FSSYXN1GZfkYy5NSAkRURcOvKUxf3HIWxIQj2H2jllqllY7LMfatupTdODUeGaF
CpYWjFPv/XSqQIZ1m2CsuwJTEpqFO8Q3u4NLhKk7o0ic0p6skLlptgP+nByKm0Ri
eAZ+4UvhTGIUicrAZkc7JkwyQb1U0leKUhDk8AvWL+FK56KFmzb+2bwczFky++fx
ZsYbPW4kvPZGkgKuajngaoqfu7AbD1NygRZ7w4D3W3wLXnvno//vO0jtV4KiUlZL
5JhZfVm/MhSGq6WmI91ksNwY0wjbwK2q+ZoGfbjTJd6G7AxxyVd1IFL5l6pzoPlc
i3qHiMhMd5kvYOmFB2P80DRZDz4ODW3hb31ibb22iMC8X3gd5htZ2Upq1b9CiMo/
k/b1xYuaSvo2KkLMKGXrLDCtDdDG1yjnJhbrJFcKQuaE0f1oNmanfoMiJFyfV5tG
nVzPbvUBGGvgMiDaGgGgFlzn0IXcO5rSaZ+nFEsxQvN/KF0guhzN1vZKAmfAdYH4
kbDuU4QEfIyxu6wU5+wbg4DXtnWx1Sgn3LckJeJnG7QEcMY88bUlo2JFfshK5aMc
EP5TO53o92ykR4YIaBnQ8zaiaWvbsFtf6ccz1qul2xgWmI3LsWnifyQYZ6+Ggl09
PF0wPpj/v8qkyqDifAr5qnCv6S+ylBxoskNv5yVb/EL6K2RFDwfxCWvyrV7urYnk
oTXvu0uJkrfjh9pKXTKcB0zfRxklqbPY2zu5xiP0+oL0IYI5EG0GBS3I8GG+DnHZ
zmH0gniYU1RiOjHFKXQ9ddwF/V4pvZEh6PH9t4owss8V0Oa+4ZGKPVT5CQFlQ74n
jNzsgQB2JiJgxpue4CjK6Pe3cb4oW3EP/eKGc9MTlmC7+MrJSPUoEpwPNCKEx5/S
044rUEtaA6ETQYfi3bcXhzjlefC080hn1kC7RZ5vPeezcsXLNRsYbjvMF44frRy4
lnuktJSZutKDl6z7/cq2wXWomcDK4uqM77A5PK0KEpz9Xp3KV0lMZE6ReM0npi4R
Ma/Mv+GXhNXFMqbLfAXvpyZIbiUHXSUK+NwprLJebBtV73W91V6Q/dGPJ1cKdfqs
LArSZbgN8eS3lRhe8G12FybrUUquCw78PydB0yhqTXSFewOMDzcjJIusbaf3j4DD
H6LXkeAU8CNSRzSNaSJf9WUQOGGrvL+g0ttW7TSR5nKGCGXtm8oa4LflIS2esehL
rVEa7bwDqXWSaowRHVVwpznwwoYOAxZQ2QzNesLmsE1FTloKj5HLAwV1pjNPCY6E
PJodRy6Fplb44qHkfGrutd9GDoLiTdS7MrhF8WMNnTd5YneBkhV9iNUZKz2d19+a
44LIbjCNT1cS6grX2jg8I/mgEteV1chzfh0sFv6FLu9CEypW+B6M8w1jRwSNb8L8
vYMp4iedtIhpXPNlQl7VXByISkmxQsJSmIrZUENKIwCrOEPpEd2rcJOa2sE3X9Ig
/3DbuAG28pc4ct9NaIlFrY/9irJv4AWuHfjNMXkVB7Lz2OVlAbzyomsRbB6q8R1o
5fHM8zGPcmiig79PKXMzb6FG8/9WfcxsfiK3jFb1j4mC+QWSGDj+pmOj36wg4aWr
0w1JACl01JC5MhPTLLhlA641NRCDE5LYCfECQcE/A8LaIEIVzaGsRomqXo6ONCBB
8w/bhCzEAiXThhcAGyb0EILz7g+zIfVqOVQsIzNMxUGNEwCadinuE6CIG2qlWtt7
E2FQ4Z+pjpvUz0DcO9dROWO1kQpIrbhW7rAiorZCN0Pd6qVu++Olkuf3Ar0j6IBx
Vj0E+Nva4xGRbrVVPrywbHJ3OhF7OosgcbR963xrWJJFjWn5UJoRdF8Kh6Ce+s/u
DhzvX/FZfXA589ah4FhjjaBi6w/5nFuGMJg1BvNwz3B1aIy8vhIRtcVNlKr7lTkS
MiIle7xVaok2Y7ELIcoyczltg9jE04sEcolXlgAA/XOdF8btfw3TOB3Yld8buTLg
yjrOh63p5OtqQOXX7G+QqLjSWatUxjG5Jpv28K34WGyIdyhAE4k5Pn89HbQiH99m
FmiFpzIXJZZfsdBaceLtQIrzt1M8y7L8RAoXtIyJcGGcUpKoCoJvmIHxp+tBFYc/
RJPJWCGak41JvLb14WVn/DoF+EUj/XMMqeOPgSXWoTa7EY2AI5YdxplaMLlkhEsS
hkWlfYMByhFV0jyawLOHF1ufMns/meqOi25Oj04RVB3GT1gJnqxQgxxIbqsyXcq0
2s6R7EYwcflKBQ4A5P+bCRqRETqjcbOR5f5EMPdyQPSw6QBsoFN+7uYZx957TS4A
ucOKBjV5lPMBmGy7BKlbE8d3uycJuxP4pN1ynQhjCq50fNhCCoFiqX+Nk84EF1Qp
MXiGuxm6/cnp0VC0MMoVtREuxMNxJ7P0ylKuhL5nHepxbNl+A2rZZNoFInkgK1V6
Z5XHbkwNGLdCeeRxLgyl6rCcjXMkaBV9eK8Rr+S1J/zoew5pBYNxRvBWqYnCXjv8
d8jrUcX/VGWV171JwLoHDpk+jq8m+4XgGoo3Y8NSMj87Fytaq4FdsO+bmRk1gbyJ
kQ5XFK8dZlf7bF+53Lr05rVsNH/pZuJTB734Zrbfv9YPqCmtgCIQ3dzXiKPTRaV9
4euKRT9QvuPkrT7CGcqMnBLnYnLg/EL7HpUWl56p+FPGzXDKidul8uedLvwHNmeb
jPa9sBaMGAlUPyPpw+6oWePind0nQZcuGdXCvIFIK6p1jLTs6ZLl6n5yA0Z5iKuP
IXKHDn9WTc9IFS5Qa5c2m7+B2Un/nGusLejsfmZojx33Keqm+usBmuf9FqIcvi5L
tiiJH6UYmFESXXfJ1fBvtHZuBRCIwSMNA0baRReuyynvbkkafDRtGcwz2qLsIs33
fA5HqTPOH60ERFnlQBcW7/llCM1u0MZR9DOwggJbEuQf2pksGywb9pFuZoYdKfLq
RavaNrke3FmL0YspE8IRfZxO5QWbjEQxQHRuxhLFzf40dxQbuomaBXiW2soSMJuR
oJoveOgM5nOtq3KdYO3JuUpNg20ZY9YRnFCFz4jdc6wHBrXfSYk9LCYdcfI5L49F
JM7jWqyVfNHHNyjZKM0do8U2mAgEuGhSnzxSnIPgMBy3qNs9fxmMiTm3MFqT9y/V
qZqRDk6q6zzHKFGac61U6dWAp5ypS9FtU8CBEfYqwDIF55EsTlv0XyJ7p6n5pGD0
gwiOoJnNXk4dwR25VrEtzWdkraqgc/tHK5QLAnOF71LWhAjm9r3wwGH7K7joT4Lu
xHCz3QAyFUoS87S8dgY944Sjc2/yd0zyhpi4NQEBTDS0LU4ao3ruLLbpt9qf3i9e
dIzXIcoWj+3MCMY5w83+nW2oQgUwZ+MPWaLKJ7bDCSC+AMz9fIaaDPOKqmY/BcPI
V8xigQyn/8fAMcSINwdav/3/pCVLR+lazuxglsVK5AI2wT+ZJsEtj+Hp+pQ+LIru
poOZXBHRgI8GGl25ucqVmd+SKVawmDhFOmI0GMTOe8Bld286RxDaX2zpd+iyCw3F
Lpt/p8Asx3MhbLvr/CBFVfezfCw/WNyArdRBlIyzqFDyusjkfLzd06EBwdFsvZCJ
0bXcr96e+OQsUIvetaiuOXkMCSVsOPzUwI8hVw5fl/+G6zZoWe/iRYi1dGT7HIgp
5an/ih486UV5iWhiegidrigRV8tshioDF43gy+62iR0fYT1km5gtARsb3k/okxxh
gPnkGq/MIqrPYdFsZRJGjAb6NyJvRHNjC7lcYPL2hYBM+29ErIGjfLPEV917KxIG
F27l+8pEsJqO4N5TAwke/+HKC4hzxGd6BGwjmdL8Pjas/F4j004Td+yPXM89/Hgt
KkM52mlRm0aa0HQKP1pOgVCiLqfg/O92a6sR5lgSB3TAoaGWqWq3y6jayHcCTFN+
WMNYBxQ4GTsO89WuVM9bTKO2X48VxJ0oQDl1887zDzyVMvIS+f7UBdNzTBUx/9ze
27dSS30T1wnPDOJDHKcAuMfcgxazU3xeov7305nuPqBu+miRxnMSBER8rO/dP5hd
VqTmdIJsiphtseB2z1o2pTKu+IZc0kTRQFuKU0dqWidF6fpigKuKwr+yCojqOIO7
lBW/gsjrgIujoiAxxDjOjWQnforBMDb77twNCgLCDXsXeaZBsyBz5mbt37FJLYFc
i7+ocinxJqd8fFPrJFDhtFAqXsyErGk3K2D2F9vsYeHjNmIkX5omzuWtfLbXMXnv
8TOToCAcXpylz+u4OJ8Wgb+GZPbsjosAFgrepL9Y93lygTaBBKdAxoFgB8HqxkDB
PCceCopH1TdWE0S2UEIlmJJom4v6ODLchfp/Ix0c51Gmt2KCFRiiiojSyLSysgc6
mzlXrYCfYXIgEnNN9Jx1h0HhpXPUoAiv3MVVETQC3ccTPm0Z+keSCfyuBdqTjnAl
0KOJckxTneTsUqdcnXFCkQ2MG1muFJKcvkgDfUUX8bniCuEyrCRNIY9y7V7DYIc3
fOKzmcVdj/jAMm7X8DzE7kqrLEmWefUoPImpDBZlLEv9JJp+ZtY59gqcv6H4CGgl
nSqQHv0Dqw8OMnKZ76iGZx4hjSbAIvR85tzgmDVk+UER04uFabnPOBDpNqCLAFvL
cH9vXV1Nr2rkRCdgvkA39lHIVvKBYNqXNsEKo3nvq4MCHIyTKvh7qaNLobXw1QRf
hJFhVUcSgxBrC/LGfQY3nF+Ir5tf5ueqjguJ73l3H5Bl5Bk8wNtD5IX+rg/7HlfK
Qv6jnpKTbQqugA73Vu0kw1YzM9WwwMAFgfYdjL41XXZWN6q21CHxExwfaMbHdhUS
KNOKmoVBGIS0yqf+UniRqbFW7ewCW7F7UQRA/ET7BCyVIF45GZKwHIckMHwtaKNA
kFVgewdry1b1n+aJWweSqk5TnmRMlRTppx50LJ1TGhK6w4OBE/pRaK9gWLH61+3K
1rwmTya2L2QCPUFN5iEtK8N4Eag75dDKkWwbvUkK9ysc9O/6mF0Q13qvzCDXqXBM
bATlB5iZ2hrZyxAxmvggT3UjjMr0QDhoBk8fD9gb2+Vo9jD7bQZW4xod8s/dlCNQ
ABtxchZu7a+Yin9eN4WNJ/qTmH7/Viaj+yvyAUCBmrTYKhzXPQIGfZpzAGQZPuee
ERccHQaWihQBj3NxkqFrsUQRhZFhci7fWl3/VHkbwweD+2CDM+0g/habdDDFdmZY
Di/d+Q33GZpTeSeTYESwmJRcWGTz/BoCvbnafJ4dUxcwMGGrQLmUrSO/BvG6pdjB
DikdUe919XuV6kkKya7UZlS7QQj1/1G33GvV5VGRyCs+xOT39d4c5GsmfEueypw+
2V55MzETNtwptdteeA1C8abhpmTrZjGZG3ysqZ/dm0Jue0KMK79dKmIupfhmZLpo
ymFQ1SKxcDI0un2LdIjcrXvPj8jR1hpZT3//S28GCldyjasSJjnoOIcfc08T6PF5
RjHIHkVVcya7+x0ZB/n+TTf+yfOpaW5MuAQj+nMujj+9zD07+W3tLs74MIludN+Z
gbxOC7eiPo6mOShJqeeJvnjaUCGxSVHeWt/G9pZStDQGJN65D7Zo6dKY6KEICXMT
o6afiGCdswmzWrB0cDQPzP5zbK1wRNECJbwn+M+sFW+4EHZ4Jcqs5QslcVsVT4NM
eXaTe3Se0gJPv2/YRUFjJRtQUKoMyvu3k8KSBm7GsgpuV2vQe/pmcPeJ1wco75aI
9g+97yHiJjINrY4UIqvQuitW57nhMngBcEukNT7RTfOha6LewWp+AH0YK/CIHwEm
JJ7UKKg++CsOtUZQqEb+01Z812ZCFRV6KgN93yHrNE4FVOL2gNcvu6uDt6FpfopE
tpS1sIPAB+e27uMJt+NgUsJrB74X9PN6/+s5NPhS9ZEUTOwr5KhY3fimBrH01mI0
QPBfSQbQpF703BaFWuNTet9XWnua858eZhPpeB++f67onweyXJcMTeUfvEHe9ubA
lLGy3V0pjB/+0MJOdg5ogSABuWjYXmjzd9oIKErRnWIMAiFb+jPvBYodeat7rLPo
nqcGrFBtXZbM1+N2yokcM6X4m7JmEEz5u1eD+Ezs4ZuuniB4VM+xyNS42zSNxq4Z
EKN6IR8a261B0kFE0Cr8d5Do+AonMwWJkx6EaN2hhPmcGVy2UGEerJTUC/9DYdpc
S9XDodN3xo14BxtfeMU5N8f1lrT3QhWwl27zII3Zclq9YEnso2vRb1wYtFulySGN
EFeSNZH74PzYgIffHcVw46bhrRNykhcdW17k6BHJpmvofBfzfvc9gHrpzTVJjeGd
di4I0i3fD5pId9NqhzsD1GKp5xnCNmCgLSy3UbVPGIXjM+nCoJyhxuUzjah2Nxqk
/n7osj3dtIaFoZ2tciAJsW72tHFerWsF4SV1M6xIMcCurME5IjTV8uX8GwnIFi8G
h61NSpzbrgubYK3dRZm+pG4HNcEI0EkPqJpRUx1m9wW1a7Ew+TjGt5F7teF9Y+hq
pwSa4q+GkXbmWZqhEpax1bHx3uWLNc3XgSxSDo3MsFliukKJGgYPMB3l9Pb+6+Ex
b9xkgRpr80mDmo6stxzZtm8cMU3Y/956DkOtc6ZV+l8Bhvd2mNWXlyZN25uNAKZe
mC8tcpZ4/mGEkZXmiCKR7NpLlSPvonU1/GmuSGb/y8G2vGDLaXI64/tnHQASNi6W
j1bZ47oj/bONJDHjaprJrzcDj3/eqONd4qCN/VAlpDLGLtsI5otWCzI9cdoura3s
Wb3Ec0veSZ95CU4v+ClXUSOZ/a8Tq1YuAipcEnPSWB2NrCUndMTrjzfKqRzuc7c1
lKK6dCuYbJ+SQ/kYj1PQW/jTWPeARXv9ui26tekD5TB/lrvaj5zcMRC9vnv9aCxW
c2l2HTdzqFKyPDO3HB0IzyZm3NZgSkIPgxniyvx5dqyIhjt0G1GfzCDqTYC3XrwW
jsApNYiveav/WZ3SlPxbDRhKZGyTa4hxEaL8gS+KEYxYuB6TlkVizE0f443uoKbs
97YEaDQp+Tni7Tgw/7lcbLTeqIdLvsIBGzU5eHqpQwL5lbS47DTJnVucTXSWrRIq
VbEN2OiwGKCDkhdeDDeAcQ1aNSK9aeiCejmSxkhKM4nZvTd8TH0qxogoQh/XfGjX
yG9U6uTeBpAie4xjqw0zxdj0Qp6kQqTxiRIlcBZsLBSZkvRKlZ2K0pH0cs2QXo+x
P0ziq4ayQ3BbW+MEah9Z867vILg7kVr3SK5j0kqTWL2gkjvwVBxUxsZCJjYnksn4
hSTMEn8CIjPBwE3ysA2QxEChetD4PUC+f5Jf/7MHoQyQrb2buPo7eDlOKqOA0OfZ
n/rU63p3e+HSUSDTqVKVY/aggMoCs5GrNtCoyW0aUPUIJAGiSbwA0JH14kcOUxD4
FcbAVYDcO2eS8eMUgdoiia5skcd0lzA16IKe8tpCekOoA0/Q7uK3znzCYOD7fRnC
ZuJTKVj7S+yH+a35ezwiZpnTwmkGIZID8DULIjZDkUXdGNdbOZJJXNWE6mrOCRLt
ll7k4Z94ko30cY4GeXwMg7FwzYt7YgDFbX59PHaGHyXQPXLXx9x10lcAOTXTgCpP
44h1GLiDyf6kijUwEB6siUs8/aI1fAYjYYYOxKvJxkZPBGKUnbkNsV+vldvhDFi9
yBBUmFQezsgwoc8x392BxS1N1c49DI7o/yrQJaLL0Rmal//+MfTVl4lxq9BPtRIo
CjlBjwKXAnWWBVEVcJ5cqW6NVfgircv/7TXBfWtN9t9iyrjC9bgk0K20qIxnrfZu
XRbi8OsIsGwV8BgY/enJxzNMZtMEX2o2MMeiH6cXqMbfAGUdNQlZ01wszralgrul
igK8p7QHfigP7Jma/BoITloAiHIZnThvZ7+Fc7E/k9TzYIJ/MVY57iVIW5LLLemo
g2VlGm2iPLdD8K85hZpWsF9yEKhksJR0UjQK6G4s1cz2QB/yER3EaU3cMrramn1v
/nJvOgHQ6T7hHOZrGvHptKyg8vRW6/GPcd4ZqxIk6uJJ2eGpvH0sBONW2QTTjeET
n6qaVZYmgx5KZV5oYHK2agnxtojEC6vMFhgnaWQ3/PHsn7rwOkZ53naZBVjJNJdJ
Zp/rmI9vG8XxHz4GGxyTIyq5ms9bkzCs3b8siDDpCNoForMoFpq9T5U8+FT3Au2Y
3oPnKs65KfGBRmNFiFTJCV8rD1MiPIfaMeVwImteS5m+XDeOzviHJvhyB+ZMHp6l
TNIaBAvkrmDRHNnto4iBwhME2D4PsOZj2mF046yfPsMoubF4NJs+HziY/u95K8rh
HJYq6P9w5yluLwrNJePzV05L31sJJQ6Mt4VcohpXzogH0z6yur6/oBZB7t+RiO8z
26q0dK5eUXvIJupF75ZOYuSeWx5nx+kaAeRT468AWPz9NKUKnNVY50Sd5KQBf6C8
C7Orz6kwHrZ1gzuaFaTEV99mL/lF9g23lvPRtz0IaC1vUKLEpZbB2JNBpSYZRph8
kXBGFwdZSmBUpM+80C7DAdsBnWdtwIAZs1ZZWOOboVEmtpqhIoIAdqZvfNVYy7z1
9YcP4HpqKGiljte6sW4B3kXyOBLOqRxAuqOgw65nqlWDYmHkxt9Db2buxCFLzvqj
lMK03HgitI2bFi6RuKChbQwS5FvjwUfP4UvsAv2h0Nn5G7YetDWGgxqiZR9Ns10O
OoHsNBFJAPFpfscPH+mKbEDBLpQzaG72sN6IIvE89EWY/AKjwCvogmBXmTRGiypq
mwmhW1Equj+Zk1Gqm0rM0owK6TxtnbHGoXocPMp/B5BCJhUiuRAExXqMQqkH+ssK
UFvnRbxojK2yGpSkevuz0lB4t+4hhMIl2x5CDSk51GyWtk7FKYkam6W3bzFXM2qv
Rbsj0+3kWrW93/1nfoV2dyyt4AnbKAb2RUu7X9SLH7R6turIcx6D+ewIUuDr6ROf
LBVfzTHBbDwcW0pGVwrsoFG0mrZhjMxO3/3+U9M8+L4UZJTu4t2dmkhvwcQzI4ka
rZEUCwg1FX+tIPLMvXMFlvd+kUgeqHmdKsSxuwUeV24jMOOoXl6RfBlKG1LJMrRV
G4/BtSN/lieoaNIFXRKL8AQKYo+MFQlnR+/BlA1yyU+HqulGxgd6QY5WeHi1wTHp
DLJP6rYsZPMYZjd2j/dKeLQcEMYJA9wH9saweZyXiZtB8H0GAHiX1WuvFuwdvI1k
k2Su+XA7h3RXHYxTMt3u4LC6WhKvf6EahK7o0oaKnCXQHu3wRcPZcYY75a1HVlJC
y++oikN46IjUCNfnO8VbOAankzpPeqzayjP6R2aWEzpBdREbNwnECSdhY5UrYR4e
/oACs2S7vL854RBebeQZDNqkVDm36WHUTjBFjvXUuhyb2RnIwsWpmfEv/iTYqA6r
OJgvtR/tsHHqWcY5Sp4AWBlfMHIewLSk0E84TPbIJHGx5QMRl5+LkVQF5qjQUwPC
JvPXUAOEQ5pDUrJvLtQOm7zFS3fAfWiA/ZMSQ0ZNqh4TCRK/WkVSns0kIm0cVuTX
CWc7xWJM7J6tb2DooIolHcdt+QEpMF+Xta9qL6jdiYCpO8V/8fMw3DC/dmuhu2E+
tSnLkivxoPbLQU76pSrcyBR+HDhtG4TjKvnRk+wCSvgGugFGWCfnJ+Gre3QyZ2r8
Dp3EzSCOThH1cVrNQF0uy83qNHcOfL25jX2svhFkBdRNtDgIr9VMxELgcMlpS1dE
g62qVKtBq7Qc77bX/DJ1MTAjMAqvE5N1UOU/JcVLJhEVOAevEGR2Aeu1mc17lxXm
Qz1g6RCM9Nu+/ODGkmXplM6V0f+VS/GXW8WIQkYMO/mlpCE2MLYXuhfGKbaK8sAQ
If11qsk1U2x3qqNmY0RajlmKO9ubE3pqYYp1jwmJwwfCBX5eJ6Xsl4QFX7ehsctB
GGgspKoIIO/pOrUz8MnFtkZaDDhPp/PoB5PkbxFHNCE0ii4w9khw+zko6V4Jvs0S
J6P6f97EX17t3HGvhwQTnHJRh/uDgiJFHHzH39fzseeLH90URnJGzHw0NrtVeu94
9Hn3J2KONx73NdeJNCUYfl4TadfU4gFs6AZCz7XuPErTYa3Zgpb0DbDOZBw/2I0c
e+P4h+FM+DN3XlnEXHgYZ4/yIvgCb8JeW9wmb7rHQLw5yD5fJfAbgvpQrx5CiQOC
KaoVzIefzrPJY05mEDJ9TVgM/zZiKk3E6abPrED530G5BfPqnaepTm00t3Dogj39
K5GCJpjs5rc4CxjdNDzprky2c98b/t66fWe+Y5m3q2uuX27/sDLU2mT0N7S7vzrD
OAM7mEGZLcSwuMNFfLu+O2RACQ9a4mrJPMiNlEGRM+PPauu61q2ZWsVO0LNsyQxt
XjXk/9y8xpj7PlfexRLXdtR6ggXhf2fS5BkOggmkydMHtu4NQHDrSevsTPofkCxz
Q7bGjtB5iWRKz/U4KP4L6LDBwMijawRCE+47HOUyTrMCcUGSLUXqiuzDs6XbNjsB
e97Hth5Oo2M1DpR6RV2NxYWo1GUs9HsuCMV2sakB66dN8z7Ukux+eQddFNdh0IwO
C3Mel6+W0rPVArB9ELl0S0uChM3K6N8/3n4iuDQuPPdc8Bnd15xIhpLoQGcfp2jS
CXJ2M5vIaIHi3bkg2blbPCnv9vLXAStfVqgxHksGA5AydEZkgCrOSMc4PhoOW2QL
miXLyVP92XF2GeqTJ2tDvYtli2M3vnjuuyHeh4XPr8mjjeoaKgb/LWyxP42SoYL9
MClL5p5nLO30J9+vOMfNJ6gxfaiI1N3BerwtV3fDji2oODpimQww7Fv7aJYP6r4W
LWbU7Su1ABrcEmYwNkDuk3h3UVzJB55Sa/y6F10qWn3JByDiOKlE0eHIFuXyPrMG
iWAzzW9yQAjX+tRZTWWfm7zd3BV5bDWG7mxskCH9COYaFLszb0PaSB0KKuiJd78c
nK6vGUr5TFgCXL+vmW0gQrj8POjIEVrIA0L6O2s1ImYxPZiMiM18Kik20hHEnRk5
eWmTk7NUSjntcjQ6EBlYGah8N5DUIHkRiU2nPznv9vc0PxMwC/dYuzbYPiNG1E0F
mE8FaJsNAp58ayAbgDRp78AJyAdasgP7LuQvqUjNkePezlQLMzuNw3iXT/tA/5dt
djr+p/MyxYzi9L5hYMs+mXkk7TxgXFbAwN0foSL4ZNbzqUZvM34/fOBuWVZuQqzX
WmF1DWuztj5jXyo4DPZ/1WF28cpL0IkdKoIuQxO8MON3IGOEIHio0QrZ8Z/P6LFm
WKtXeghZrZdeswGvKgHi7xzratpWuKADyFVbrv+p//KxKoKJEBw4lq4G1vBeQet/
btX6ICmD1FVh4oupyA67cwj51t/GZT2Uf/Cw9WYYvzClejhnzuF1yNsI/PGx5/iv
JkFNQWb5AxsuxqDF9gQ+Vrv96OrHbvGvktbibDHzgK2akRph7IrlMG710G4qb1rg
YuML6205kF9C7BFhGum2cRWxnJge5ILB13crBc/tvwPjVRMTdldJ0vrdb3m1Gf0E
3YIhAUT68eYKbIUc2DBrwN2YdAQIwZMMbVoiPNEUU9Nmg+BEUtsK6WGOi82pCVp+
RSwVb/tyCUbeapr2Pp3mEAny8laeDLZeKm+4CN4fsF+LlVwjgl8+l3vGk1HDdwcK
mJO9Jd5N40hEbcC4PR+848OhbSL0qFHUrfduoMaHKFPPyJE+jZGGpbrNgEMeBkzy
AVWh8l6FQfl6ajYI1+EbWrDE0S1b/pcI95AYXAe/rngqV+a1fZFwd8YNaGkfq5LL
wiq3PZr7JGeS1wCB0/4ucKs1z6O4coXItd3vj4sBxpTpprueMR+SXlMsgaVZ3Z1C
4KFI65bHnNjsTd3pwcX+Hyv2UjsTUD040k4zNLV/NuPE4BXJhGG/u4uBpJKzmDsP
EU995CUvF9V/SEVAB88qHDaENOKHi6CcdQp7nDpe3Nqmmw5H+2kNTlCsIaTWUCs0
2JSofVgV2ly8nOhu7Lub2Q2UpOdy55Wrbw5sQ/y4rPGi0l/hy1AX1eZhgGNftrJV
Z+WW6kX7UHesEaNmbXI2nbYb097wf3hxn37wREvLDDlSNE9mamOUENOMeab9jPCJ
x+/r7sjHKaKIQASraxUKgoJoL65b7ps3+0sHnkFrlxgbp22GbmQ1pSphqipt9vVk
f+3npaKzCSUHu7EDHWNz7RZqo4Wol8XTrnYRW+Mf3HTHKxbZ3dzF9SiadMubR6sf
`protect END_PROTECTED
