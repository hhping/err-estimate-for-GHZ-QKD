`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSEHPmsujSAZQt9Uvawcz8/rlSow/MfhyB0T7qTdqrFUkC7TfLcFXGrOjFoeHrYq
q0UT5fVdCBwzF1BoKfXeboIYIXgJzmIF8VYIAsq/jwislKwj9OF1X3y4b9+Ugx0A
AXYPD0uZCMQZKfpbClqUmuH+5AUyPMzJ988AVeWgjuVHt6grVYpEztr/qr4JleCx
HRgP14NBhhT+WLf1dKjaYhvpuxQl4+xIe0xwxq2piQa3cvmTBTnN5QpPPsM8CRcx
T6rnOMH3nyPxgxDd8sWorfg/KLeOoMDjvgKiURuAODeuyghZnuI1Z4KlnC8IISvy
lxD/sdqgUbWqwqON8qfIxaAsNQScSsTKSh8AzTltqofmoyym3BYkhfhvtUPfrWpF
jxkLGkB83MEg04Asa7Lp6MHMCbm+7YXtBCzGjKog7MxN1M4CzOviT2SV3MRQNzR2
0+FHu+25hWe/PXzOTujcSCQMmD/63QdGcJ5aFUudm+5BHfLkv7dEC8qcKtkbBMSd
WtDy3WAin90TwRO5/1RFSaf48kHAZIcO0nBKD3MGuDZE139TbMb/wMvCC7G6GKVA
144VbKsaO+56alxf9U5NsPc3rP4upEPlTjIOJOtSdbycrd+ztHWZkSZdZFmfKuW9
t+vbIOP6i2/DnNvmFvFf78Xwj04R3XEJ9c8I8nuS1a/4CKAZmr7qUGy12S5Cx/r7
YHcgys7fwm7NaNlizXlKpW0V35Nqbrd+JS2iHc70ooGB9j1JdsJzNpwXlnUPfyOP
a+QZ/Nfc+lGaY4toLzf76GLHZ8iqGQGeua2XSoNzc5B/t0dAf+6frwG4GmQOjVka
0hmPzNlvL8eKy2ffFmyXG49DMsnkax7CVYxBi+luTLh+NydDi+kEg7SK48LGgPDY
iuUePz6Uww8i4RopZyvD6Mb8ZEhZSWYZHJVGDaBt3XNhflLEpYGxRoXgRhFeovew
D1UPFhA/Kw3HXjMWOX/IJH9SQDHDAJ/uadY2P75RKMz/xBYfKgfrFhLDYUtayUbJ
qzQ2WIozAPm9lej97GsXVgUtR/EPtYF0LRjwTDqbsq899AjEqI3Q750KhBxkpwsA
F79aZESvq/H+IWgqPIjo80WnKwx6M7RsBcYn/um0HXRhNJVzNKvyDr+HgSjOpquK
fF4L6T7GmuL3VIbGvb2KKGnFFC6ZAWiqpIlEmURnVNw3YxWZIjQLKmHuOaLoqYUF
oknB0xCpEzgKA0zwjSMmCzed/cDXt23ATyRA0cvG/IKPQJiDQzjuqMhIUByDLjyG
1JR+vR/+HU/Nw/xrxdEwoik13iF/6X80SJSTyDmLzf53wXuCbwiRqZI117wZlxR/
7TNeF9j0QKZPVUdsb5aAchFur0w0UQuJKnAHC+w8XFgOSnabR3HwQWRDyDZZ4yku
7jz69D7gLBi6bfzZ/5kIyTLDyTDsg8rKcx89KttwpNPCledz6cErj+yGWfzuyH1C
DxvQEQjMUKPlz1JHxvVvN9nkf23pZjSWGtZruznenhBL5KrFV9XE57EwXEN/Dt0E
9nSYv8piHKgRlbB6K/CmeLilcpWa+mOOuGVBrWmm8+a4UYCOcMXxh+0g+l0lay69
s67b9wTSiCOSdwHgYi34XSpKb148ZFto2d9yUZXYpaTdbiLeIgYJR+rtzkKbPTtT
uQnj6eWwtsHpPquE2fppPOHCPx9R/v8VAumIU1ezkrh/tx1HCiIkEDuKMcVOyzCv
YbwfWILhx386mcm+lNMlE9xULeZ78Uh5UMRHxkzLDXtoGLQf1pInFQD+gwY7QC9V
fbZXmakR54YRnY9s15tF1CCfMXYoEzgfXTbCbrB1FTOTdKZhw+gMIguK2VSzwlmj
tfRca/2SvFWdOuzh/OQAicONBqC2VGUzqQipQv943z1OzNTnLRZ4WN2EJArfpNsp
JXbVWPkly2kds7QgsoIVEsJYUcIYJgC0ZTJZ/VRdDau+nsl00A+jHHeDq3SGtaV8
JigRd8gg1ITVccP4KA+PpkkyyCMV9IPg0WMwwI6d5D7leezGzvZ4qLlNjWB+gZXO
hiAj80CRpbX3DNpdWAfTMerWNd5/o5ae+YIjtmsmpF6+nrlTP1/LgKk/PuQjUvRv
go5HeWmKmIN/0XY4CEKtvLk2uWfs1Hp+JjSb/rhdbUZHuOev9+pAjna6pOab24d1
GfDsvXEQBgSi+p9D/HEHqBwOSKBlPHQJK6sTYvLZ8UkGGpsMBniughfIcBV4aSoV
8NuSqYd1YLybqP96M54yCg1qRf3lxGmGmKheJEKb2QRld6O3BB5Q5GQ2PLcYvINF
WyhGYTdHZNUvy5WLZvTXKY/ClYV9dZowPOrIrxo1rl604GnqIBB0BeqTL2EBgk2U
lWK+iNg7gWp0Qfmc8yp898ApfyGEvOag3xpvXt1z3mpmogh2FycRTlLe+7UoqELU
pBaHz/q4Bu4yYaz/jRXHv68KheATpS5TTJAO/f0g4gNpe3XCZw1vSp0wjIaMZJkL
Cw1IALiuq+3xmP/b0Nrh4KZpNBegDOzSrU/CPNXQAYI2D0YJCPUn+1sqlXXjULk+
4xJ0DJKUyVSfPSqnfBtdabOxdqMAvpl053IJv3os6aa7+pOJgbYn/+aJPdg8up6o
6pihFfSoccV6oCd2hSOBayc5Umf4N1GDUvsGXayGalkoY/eaqS+5ga+dyMZONXE+
8WfC+RaoyYHGwIS6KgqXcoSWhElTwYsxxMiYa3BMNBzM5XnnVvrxL7HRMt46+FO+
eEW3xVqeTJj1r2yXTZ9J0Mo+/C3dph3SOK0gnQG/THiikAmfTRSY6hNHozkSWpOz
V5O6RRrRsyan/ACQxlDsL5XyDWgARBcO8t/uVDyZe/VC2FyMnz6475iw0xTk377y
W8UlcZ3aiqz7o/iZ+2zt/sitAnwizqb+al27DWsMOlJpFlmfJcrx1M/KT4/Xtcr1
lSsKhMVw+eKdXCGUYTTIqZ630Sp8wtK/vd7pKK3VqMlq0+7IcCf+eqTbscpU2sTF
x17Zc6KlxBCggdDoBhKmPeom1JxvHOH7il4dmjXaf1rfRNzCRaMsf8GDIdN/Ho/h
4DZyQmYMzJloINRhwZ59Lf6NnGOzYc78ynx4z3zrEXCPZgCYZqONyZBTW6o9rXwK
YoHI3omJjwq7fTQdk5X14fbTHiN9bwrhJKUzOIFUMVNufTGLBVm/8BgE2LAuHTu3
s/9xdfRdxING3lDtRT6ncCxsd/E2DXxwL98kfuv/HI2T8ith6o63oJVLt/I1UZk2
+I+HDNN/Ab8sinxYqUqK8d7GhMQVfNDKSgK/iM+k8ggcjyY15cJBZeocw8HpY6sJ
/NsbMiheSbFW+UFfyzPo6aHD9490vs22ZZbdC7wlWm/p9mOrdK409z13St6e6Z1I
kYO1tjl3w5NLRPTxOnft5YFqvMu7JvaSzgJdx8NSFdMGotBWDGF0g0RUYFcoMFV7
gkak1+9N9t7wEXmcKviRk7frd48EndXHOK1v/a+KFAXPm0WBfzaGbvfepBQ1IwRZ
Psg9ux0HzKkjgL7uXCzwAVCeKi1GmMcOiKm8lkvgm7XmkgWYjhx8SjiPztG9+yrD
01hjWBfBLUxzFglJ7QtwsxQP6ACu7H3AKkjkIsqMtcisdpPYYtvgwRy+BbRvRrFA
64QuSKz02PAJc9+vyob+1G5P23eeqPodAevdd2oag7g+NFLKRdig7QUJzvCMkpBy
o3F5OA+f3N5Q4asT4NhhqYCx+9iaz//3PqiLbnsL2HT2BaW75RqGGG6WdeN/wkUZ
kiOCcVdLzGOEkCz7kzob4yX+puDkYps8HtyVfx9yzV1tGTIir9vRLppYOE9GVqPN
xo0PGBblG2IW1/ueqiCq2oYPMGcRWZlKWBdEoOUD0TsMhGP9HWWxMFobfZzc9lV5
RAvzw7bPzDqS5qTeINZIclWdNfcT6qSqt+578cWt834BO43mW7K0epXM9FSbCAm3
z1dG824IrioJr0Ez6nzavArT95PX1NFGYWZI3fMnZdBcUngRihHcX8/ooFstVqLq
2ht3pIEmSZwMN3vWkDID110+GJAqDhFoJyWHbYxFIXxdN4eErnRc6X4980vgABI6
B4/JJW6x4z54Cn0PwX9OOgp7qXpX3rNDKRhDaO8Di1VuAoX5jxLNv3CLny98QTn1
p0jaMUOld0nqcYU4bzU7FXhwTGZYC5SXymEoZ9KiMaOzhV6Cs+yM7vpPO2dhpda2
rYP5PRWa9kKI5isYAznZXWgAZb1M+OnFI+EYdM43GiBSsJ/AKjPJjT27Ln5PPr62
/MZ6qIrpuNxf/4jeL/QnJ518JsfH8AN572Tt9E+dGU8l7o/i+d+YoZaeEcPV3Ee4
kqo6/Uspb+ttFFln2jZe6aRSV514FqLgqGDC5cdnEUhU1QSl1JgrZTEduWcAcPpT
1o6g3DOQJqLVP3Z2DMGJKsAaGf3yUG3ujme5UIyMwgH8wuAOOSn29pJeAkpFjj3+
rdim+SjmDfkGAW6n8SRE50dDWfJi4v0nUGcOHuFdWa28N8Uw3sCwJdycjrIylONa
kbFvGWT9TGEfVm96S2x1EsgQH6WkBFpoj2P9iuDqxjjMkkLv5Zy9Aw39cQEdUZzn
b26PLdKoUbbEavMES/VDqcfR9RrZvOPHlHcSDwZJF8Na2n53vsh5iVhy7feeD+Fl
3WX2XWYv488maj56VcLrMMkUyFHz5oVf38fsp13ivhcVC/KOnaakiXep3BwUb2Uz
JUCwLK6rcW8tnbwyEpv0chFDeK42ftJgZvIpOdivUFB0kqJH+XvrVMu1UZGpKijR
CcHcPZIBtq9cyHcQITnFcjgdZ0QGb/p1TDJU3xkaFBi5LDzY9LXBbQVDL2B+Pxys
fu6yyjdLRhiO8Q4BYK4JHXcYsG44bqV99jrXsZsfAKNiRAzZs8bmmles855tHS1O
ay3dbUdh6KsiYTVguLPfKiuCBavMXkLFGCIgtjBBf8T46apzw+eZ9PhlEmRgxBtJ
NmvcSlQoqVusEh/mWrwOIuUgp4S98yF1AaxE4gz4fRum9QwaEOfCHiN2N8iHH5ek
cgas4RUcKXjXbB8Lygktt/+nJmp6Wb6dFb6HSLVt1ezqG30E5ZdGZnq/i24K+Zql
NdhOntRQdfOG6fbOdk2/bNvo7+8vNqLyagIFO8BWMzeymghHBiAIuailUoGGUwyr
avNw7nMJY/cwMIWDHiqzKMlWle1gOuL4CkdAPiTa05HjelBBgwTcc9HBeCpYcxj2
Fn3bpCZGvBaJZ7XqrSdA60SHoPaluh3Rdtc9AlRXRfz4UQxeVTIrKSi7qApRvPvV
cODY8UP0oihx/44mJkHgGpJV+DzzdYI7PFcYx+tHlVueL1lf1d+MVfvBeoQP1E2k
fWqktHFZNvyfxM8NPYIP8ispZSFDr7G5BelKoUdSwQsFr8GhloVBn1C8t1W88UKL
DMGBrfbk6zg+Ybn+9TgNNdPKcNOqX4i0kIdeahFl4l0MjZ8V7lZC8gvbKNTgDMZ9
fO06KX2rQveXDwjEnYwaEdW4OcO4Va+57ABZ7sZ7Vd0WIZ391AVuZPk5T+vAGG2k
rioQGE8VVR9LkZIdZEUSyEQeHrvBsHENFl9YLWvUCWhb4CD4BHqoE9dnsF4ESK8G
HxoaWsKzFzrTvMbsOFmhBLbG/VB5IVUJ381kEL5PkRBRllLL4eaWWEgYy+u7iXWG
n3348M9fqGoOhLSJV/jQdT03OE9/XzxuLzES3TPVZ8alQv1BPaKFeQs4P5boLpFg
Q7xmutIVqnsILHpX9pXDDXtkpExochCwgh3cM2GdlYIR2tPrNUWvQfQZY6AZ+/wR
/p8o+wcM0d8JmWmyakBLwvYHk83J0++yOVW3kkloWWhogJlQnaZDMdHCoUvosn8X
Ija2EvOQRaVCpg2E4u1Gxb68iNtU49V7awWTvGenzL7XwFDqP7mjzIxWx22DJ3fB
di5eWNfIU+XuYml4/668VUYZU1fxrz3kVHKiZPbL9NJ1RqbNfhcHz+dGNJQS3TYx
Nq568JfU55ZGm3yjyrhM0DbHLbMW8adQwH9hBbjgVAHV9i4ItlZaIp/+bfJOTeCh
MZ3lpWJIYNQIiwghIki7o+jwnZ3cgiUjk6oqgxrH2kK49MR1wq9oV/P06C2ReWJE
gdnEBWwu0IfBJ0a146Gk1eAaP0/Cocb4o/TKZwhfrvbOoMqGqleqjTJk/8+V92Kt
mjjnIDdpVJceywt7DOvrLFlnnwsfh6AKQCc35MegGwg5oIFU9Ind2xdUAAeNBDbT
stbm0Em/sKTxoAWqC2v26jqu5XtAYRh5XHmBpJ98elmAPSjZmnJo8vTXfnIgF4jv
qNzPbmwq/R7EVvkCrC1yAgW2mGORzhlGD1oHq5yiR06M1DWJOjcmru3xrNwqlUB7
ALcem/xlSborkEpNBR1i+p837BzaTxBdk5hBOLPcxkBKVLndbM51HsRzgpX1n11a
1eLRq7A7E7CIMlYFkFjoHO2sXwogqcAGAunz1BJ3MWe3oZj6j00vgA8l13K62rBo
uJGCADTfmIP3Un/G2yMekuf3KLPvLoqaesncnc4HLDw3NM+EXS4W6k8ra1IYN4oI
GrYSgsYWfjRbYr/sKBAlSv1pg3rG3Sd3DdQNhrhs1MywsS/Tb0xfeXYpKYEH96xe
9LYokiyKkzX929VKTDkNnshf8KgfYvPS0XojEoSHKXH/Ik6IZi/NPpziXdNDlHu8
2LY4p8KWNkaGYO7234D4ATdWP2brgV33CKe/M1jo0haPOUPYpObn0lik+YhpQ4P0
M+APPcTrRdr5J9ZY8qsyr1uXdBJGPMWyCtpZBahfgJxMaXhye+k5SmqUXb6Clweo
1/NPuLu6e+5bNM5MkBbCPVk5msb6ekcQbQVpSbhIdRCRPTZT4tmsEEn+23VSZD9+
WBKUM4xeIwNJpp7aQr5s02mYettC9JhKpa801G9Awie+8m+9fd2kkOS04BnxMkCJ
3iZENEYQA8oC587Mq9YPucNTrO4d5tbw/F3xw+PF6xPOheK/kT7WG5B6Tv8DWC+n
CwbcekpjwtbXX3AzAQSFKoDcASIlsqJpRoivaJh9Y9qvCG0o5dgkICRgllNa0GbR
ltlngUIBT2QU3AP9ofRo/roFgggnpCW/wICjFTCCZ0VAans+j/S06udL1LGcdi4L
aNTFHT/P5T6gzKtE9cYAwgOqBuzZizoF9nZWd5g1DtU0Jb1k9ZwYIYyzJgW6HM3m
FjtWyC9xTW3P8KEsoN8R4vMCbM2Fju0voYlElUI6ib4Xq+OdVxfd/BceV1tVJDHd
IRQmtGB///E8phh6v7CYtfLIlqpqbSJf43yn1uO9E5qV2LpVh8SmFipUIbs5Vkga
Sc9SPslhhbOiS8kw36oH07JB7lgUcypk6bgWa3amJ+f6Y4qMI37ZGzuIa+hUtWBs
LzaZo/9gshhcULvLV47fHNUmvv4cefB7HaHbep7gKSLQ3ksXghnkLxdWvfe3QH2u
akIgyjY5tedHisfcDvp5zcj6jvwpOiqoATZwRUDh+h2mOX4BOgjbl9bniCgs62N6
nMP6gMDzdfyNWf//HXm2XHHU5NF4mrQUOcAUmoUSeDS1RobCx9r2hTBjdr9CU8LN
oPYd3pwDTbhFvwo5fYaZ0OK7gyni/cJIvToLg+X8ReUjqD1pROGSuM+tbDccvPGr
VbD5hqzHy+8GDxUUcBMLeXqLUUsWgcknlHXvLduKPdMM5TRgM1+deJYPlzv8y7xV
pglMiR/dYGFllLpuZNu4niRGmK6RZN06W3mI1o4jW8gdK92OPbkabYwo4njO1xRi
3Xc3I9V34R+b7o1rWcR+7xf7rzx+XC7EhcqDbUFxBQZBAdvbNUTvBDcvSzMgrVNO
jqjkfwZX5syCZZj16uKjkESndCMfMGTIS0lh034F3BQzS9I2s0S+NkhDL1BZhnMl
YA39BbhdtshBaeEMGJ3IJCt8hKvEucIRx48TsAZwXzTZqdR4dEi/pA3xKZD3FH5+
bBaHbRY5fpJ520eqTiuhJI4EQIbMg6q21aJsI3lgpvFVLHQuV6F23ch0xmyJ/nyr
DCx+/2HaFNHfiVgk4xslDTyz6hLuGdkkGVPvhTe1doB8le3zGmOel5xSaqi+CN3k
pKsjKW+1drFAFrdMThQKYoUjbopdjGXBjgZbcNMSEOAytzua3xPV4W1Fo/zmRmo9
uCSZfcFWxZ8dxHxt5Bt5PRe5gE0D5kfM1BPkKIg64QGs2oUmeHc/FHDnT/0YB/F0
CCmabUo+nx7AnesZHRSg+3/79F7ALHSqxSpomExZ/Bt196+HbmnBwHls5BN33uOw
0mAy/P4p0nyGeXmXEwDUz54m3g3NjnCH8c1dlHzSJYnVatjIIuqqjSQeUgPk5WLf
Oto4UwKBnc1ci3yCmAoGqaSKdLeqYhWV3ubS7Ez2rH5WcBaYjGC49Gjhs5U/+oDf
iB+E3g20TB0M199Mn7CusmkfW5/yOa6xnkpmYaaFa+RBlOaBC8qWBCfMJV1+qAdk
tUkWTQFD2NrA3JMUfjtnQxH7ea6Dp0RxnKBJlIIh5Xv+K8EmwWarBtPsBjtaqY4Y
AdgkR3lnUfyuY54OXpJXpxlPBcmOMfevVRLUjwi89tj2M/gyPup7hYRWcX1Fulj6
W1zLRPZeFCi3LjI8usA9So110AZzEVPYDyYyQT3m5Cf94cAp+JyCd9FZ1pjeZ5Vn
zrmQuTbU/k+OfZw8DVDKZRhmTLg+Z/1KgEQRoMm/xJCNCrd7NIL3PG8v0hKnnZLc
RzSvhz2znM7EbIKDHNInYuWGp7PkIUAP2Qa5ioYKqy5pWn3hR2P1Wg46nUbq6Hou
vomUkgTfNzNZ2zEeTIcnxS3lx9Qh/tMwqbmpnYJrP3YIM0h5mDG6XnyUC25L7j20
m/Njm+r5BAMqZ0jVZH4qwSQq04Rr65wvi/BFpHlOjXKS5ldUITPiPVlnXql/61f4
6Jq2Pe7FBHHe/CCaYPX+c5rZBJ4rvTgxrurunqo1VzjsEGlh9j12fAuk/dXwtUsn
abkRFogdfE1xgTyIO0+VLbbSysHvLapatL+oXQNjppm0nE6VazHd6WfCiBM49Yck
VQrxdxCLC22LQIty8+iJS7UYJY/0CKZPZfEy80CSyuud+1ilzTg2Xo+k/gvTCtNe
Cw/HEKi/Ka4dHcuzG1smdZzbtvWamSnLopXcj+9bFxh/0FTmkB8zHrZJ2dTzyZJk
h/DfGF51S8WMQvyyx/AbSodMPCe2vawnKreIp/Hz+EWpyERztmUDdMMp+6IOrpKP
3zw7L/+5kFvGlETrN+U++EFBhgKMeTXvFbkeAoVRPJ8gt5NZqlXjMbcm/fNOSTcg
mArvbRFCCGZiS6ffz7bEHR3loPB6APdcnkQmie5/Hva8eSic6dm7kQ/WIz2YyqH/
Iu4YEmYg5rKuHqiq0xe15f7V5eBX8NHmFO8YLSohqiuARxQn1Vl69T7c4buPMEjx
A0rSwY72va3tsT/e/ftlfPtkwNRBXlKfGlREJZLDJ0PflLGVX2eTSQ99UOQbwODG
NUtpkVvr11Q3CXaDpqgc/qCQDhN4/hedjqDkAb+484oIwWrTjJmtUdwu+Mj0IVHn
y3KYvWZosPgyl3V8kCftzwPsoFx3EEyc4wUuR3O9N6m0uOMvB+OA6NSNd97eBxhl
QGgULRb2DZOJrpUDQ0gGlzO8IoCVsPSPHDRfNrosMw+nC+TdOyl2RAaW92H68b43
/KXA6QFubWgwk3P4lMTvcS0iiSgz0L7FF5ssaWC5r+ongI0akSzpX31zr3tuDSzY
9DfLLcPdBCeZbesGHag/x7vQaloZk/9UNa3XGmnkpg39i/DyaI2dh/aLNQMfa39C
DAT0k1kXaCt4IiAsIuJfNbdkjmSCZZ0ulG9e+Bgd6WSm73qdCSQQTr3szfeIRBk1
1EXAVTTtkFaiE2LCoDL3mmE6GW6pi14wDSy6NmjfCpqZAOE800u360bq9CgfKVry
P6uDzPDOVXWUav9vLhGA+Q75dgMisJl3Ea/Yml/7asbdLalhNksu6XrDm1ZwU8NC
QaExmYo7lOG0e5L5feino8vOgn6r5GygdqxYdEaYjyXI6E42nG5Lknl1+Tlww2S4
VAErk00fh3dD3o1nfbyM02fxYvGXHPLu2+xD9LaBb4Ke8cCiqz/3nPsfYBlKMYLJ
Ysgs6empWnNGBz7skCcJLpk/ejkRN9ZvtzlsmPTnzFhq1Ajp3QOANwHXDmARRqE8
O3NCrGDAvveFuDjP5/vq752SZHg9SktxUpKaZRj0PyKB3lub+9FdVCKhRFMmI6WN
DmdT3xO2CrprqNypDdoF0T7Uc9Jxct4l3wJVBqT0UEW/XsQdoRMZv6mhbQU+1ljm
sXUNYd0qrAUX3U+KnXNSkmWTe4wZQzqPJEpejUf/KbIKR5xyuAMfFte3yw/OqeOD
V7cgoPeCzCw8i48/q9ml5QRaK8U6GTqaaTK9ZWmui29G/mXjuvGH1cwO3KF5qAFZ
22KCtqFOQybfHrqtgkOD7Cer3jppfuyKrWL8rJOtWKibjnytowMvO1+b8L9aXorV
Np8WayLONYjyY/nkg4cofEtqWJTL5+y8Ssn+vTW/7epEe8rBfPj/vfL9ifLftlsq
Wv2WbodC4vhOcxqJZBBO+H27BR9aioZwwCUb6p9boIML19R+wjprYWQwdyvpAMaB
xUQScN/5fBYTXjKyq4YAUPnWUwwgZSS+JmSddnNbhuDjYHOoIZ6CaRKpNLM5pLOR
9Qlfv6cSxQkTWy2zQz8R6fiLqMDQiJTYuH5lkb0S3tHM2mHobNgPESlGsAWYXN7W
KJ8d9ZoOH82afhSl7Hdjn+nyqUo3a5gwrxqxEhr0kjSEt6CoRpcqL5wroxnkRJKv
PWN7kb8srDV1k85kd/DYtN0WkDvDyhDFHi9wQKpXUq34gmn5jYaAMuW7BgOU1oaP
WAo/6dU5CKJmBynMMOQnggxpuogKVqWjPOur1UvKlHh0BBOWJSG8i9cyqR3X0F5r
aOmOP07y/EXp0NmJn7L985qpMxjaDjOqPZVs6JWHtHKz1i/moo8MWpnc2z8DGRsI
6WHg5S17XITgldw1Am3ljHJmvfWPuJzhzccK0yOT4iwCgP/UNFOvXJtYhSRORBAc
FIWKujrv8Gs7kHswJTcvP54rekjWWXNm6T9YSpy7iBoubcPgXecVwPNTYKcpmyR7
h7hS1AxCT4Bm3vgvy7t4ZwZJoYuC9JJtxwdUARliamRUVEdU4xp6Qnc0u+UY3oNJ
Zj5wgXMCVqoJdA2TV30wHTMLV785lXk+cKRnsATN5Y7ksOH9KVG4ssyMtNLRCG7U
CIIWjUOsBNVtyqonAKvJPufJ2Opu4l/eLaN9D2VLfTyhV6wXZN2JeuGQ9YiQaJBz
sXYBZJj2AqS26SaqF1ej2E9zvTwUgCnGeeRUndqmM7Q0UqZKL27RjCYNBDBDDUGP
1USadlpLz3kFtrlurUwmsvPthEoJjKP+qxmBu9nG7KPupZBedpRjaXiVYiw87Ufx
wj+WLiaXcl8qqIH1OcUztX1f/WUKahQhUBNSI8fgChB9m/KSA6T93TsLTXX5vELs
Y93mbEEa+TMh7vu2kHUElymD+cf1UgUhll7mZI+O7Op/HgYWLxiEKSQfQw2G6yVo
H5PyUX0ogJALsm1FmfOzpFeRj05IlWWh3Cf0C/jkMLO0suZIZKc8X8VNiwoNFkyX
eRJYZwOEa0UzzK6U2FyttMVkoIo5yDxykg2pXNlEzLAkIFBofxhtMzwyU38Aeyxv
gevWUBZC1sIVck/9+nsH23f+0ZZoQNvtZWIBSToIReM7orkzFE5WArMb65bMscXq
cdY1+z4hnbD7bbVTxqngM3u+N0gAhP0ytevv7ipmAg0RBuiVFmqSxq52fVFaR3ij
DZtWV4LiMMrab5md9+f/Hn92Jfh9g4ZQp28QXA9O1VEjR+1XYtajYwzrPdV8TMsQ
+nZyaFxuuc8BMkxtu/8u+j6BqLv3aSffU7nNForDVIG/58IA0Wm9abADkSwfehks
I4EayAFYX8sAy/kdBXAzyM5cVpKD07UiDh8C7fG77IymoIp3ANtHSuo73ktoUJYP
B10ZCSmK0DCAfsl4rxsgNLNnXlbW13pD/PqXOdM+uw6XAp+VyNeDxp0OUYmVH30h
S8azInENCen8llBvLY5pUzxllKT5j884VwRoKbV3vCO3hamDFn8DHiLa5SM+oHxL
Xh7czfymtkcw1mjYxW+Kj+1cPouZ6UzV9TOBfw71Hsr5mCEmvtXA4BJhX689KHve
QS5AklyQDvWlVTOhxPCTMCR9Lx8p91kabNDLTuCgoI2q90rD+TrnHKDrELuZvg7V
SaNyMHZVcicH+mV2QLHVoXMShE/OSbf9lX+6dn3gLvPWT1aK7ZXJebe+rtwgDiJL
3PRDjbIQF4U9XERr39vdQLfIPoMm8F6nXg6tz2oeSZhq+m7rNOtUDf/EsPBVMMzu
62Rff6oNCB8aGRKCVCEAvpjlO0BRU3qOHfLjxkVjSDCrqLUIeg4Jis0ql4tPGS2J
NSd8iKRNJsaB3nx5a7ciQRs/ORfjJIKLpvl4fs/Dabf3hixFw4u784c8QsJnLaR8
U0Ydxbf9ENDDvQl2yTr4ow==
`protect END_PROTECTED
