`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrziUsqcWY2JnIAzFfH0ql3ouFJMhldWIUX3+/R0uAOVl0l5BfQzY33ehgmfxQGl
31ax0unFKugtxzrf4pURHRR/08V59ZPPuB4icu417281aDNzluuM0CYfJRgQSYhB
Hqz/8nbNY+pntiIace6qMHD9D8Jb2obknYLr04BH7VoOYWm1k00uOhDi9+CNVv6M
Hh1dLo2uZ+K85bjQ73jEdQ9vGP/1Ni1GoDQkSQy1yRlxcJLTaBnTtIq0gnuSe2P8
x6KlMZ9VBBb9TKptGB23LL+k5SebGhh+ocB6mpEzB2sbHAu4ZxjD7lEd62UY85pp
Bfp28qEcnthNKOfFnReRQxWZrSmo4/M+SvLHuNTNo6OxO+oq+q3uULa/m9b/30Ef
OOZGYpsZ193SPzrqn66ZrGR4EUCGlNkA5BN/mvFqSHxSDRXG5xVC7D1V6dsMeDCs
fZCCvB8lqwQSQqdr+x3W+A==
`protect END_PROTECTED
