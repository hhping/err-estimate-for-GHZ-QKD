`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bke6N9Z7SccfILIh7w1XcXts93qZ3p2s8TgNQOUJk0leT6bLRvSEKcmFh1KWO3sE
V3iKtS/APWuZjQ4bhExe7CS65mcUHG7Qx9qqGj3hDPvs+pmtK+lpRWU9yOwmh4Cu
BjIQN5jTvg0yuhMqNnPmEkQLUP00L+1BrRYWiDAeW0hsJjPQa/tCzkXC5IB17XHS
DOgYTTKHpLFgrDXNT5rcwSjVxqZjoUwZ+tm/+EaIC7JrVOnJFnuWGS4zCRCmvyb+
g0tCNOKKnwU+AkGgjYVkJyRv+ywLjoOTcsXmSQafXgm9suIbnhgWskSzA3ZmbvVh
eyyPzkhMr0bFnUww27/MT61Q+fxBKFhxSEWq6KkiiPUZpzXgGjwooyT0fYluEx56
XfUzA9PWs2xKezb11N2IvZDaWeG/dqLUNl3InxoOCustH4BP4TXW4708od3zkn/O
CvTWrBWEVFvJSv7VMZhmq94KrpcStB4FMrj3ywP68vAvyxyR4xOscKZsaJqCahQZ
qJCsO8NUPtVuqqUYJPrx8uvI7gO38s/QQf3DF9Lv1JOBGPS55EqSBr8voOPwn7V1
3cbw08ROP9z6oxy9mfS9rg68ciscvV9NcQ93pChw0RUGq6o2+jX/Riz1JZmcCktc
UQ4X1Hxxj56WwfVQNsy9ZrTNCNGSZyKi8FfYweEAQeyiUpN4iHRO2YnJHn+XfKcC
PVEM9/7lkZr9wmDnpM1TZDfbGksp9TcDVyGz1CZBAkqaHpFrfSD33EYZnRHTMx6h
ZOGBEYtSCLCRxaL3sOsFuStmj0nM7XB3ahPkcDgDWiMHUwdlq9gvywe0hUsY4FRi
PYnXI3utVmcgTomLeNXdrg==
`protect END_PROTECTED
