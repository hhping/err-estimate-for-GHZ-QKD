`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQ5joiloNfrNJPOakimzg0epXdRG4NkPoqm/n2FyLxEjhbanlO+PMaEl+tszD4i4
tgDYTlsJnr6iWZtc0KvtxucP6dZ8kDlVPOLDRl/TSvxNmaKK3WCvYUpbISTVnuKd
8LZsVagGuDxb+ojavLgj8+yRol/m4Ra5md5qudIHEMJviDKbkg8lLbbHnQS2jwrt
rCc5sM2lo6rEiuo2wew9gk7fgnq93rNSmkoD9WUt1nqR4NDDhbTqhmhs5hYOeKYs
GdUUm/ceGmm65xK0KiS9choT1pznPFjw7ALrthHHMf1rF1BLsyl0O0PMDOofe9m6
ThH4FvvAnyKzVqwzG/v8HyndgiRSApyU8X7xrJKaxVJS0L9womXwyCHyc3EP9GMx
iTfQruef7tGmsgi13wzqDcc3M0Bw95CbXZy5NqvvkxN9WPUteGBeBZ0PgU6NLgM9
XTHlObpvY+zmRWr4OL+yOSUC6R+bnrFUXFKgYnZ4Gb1FLpfw9cCT8TYHPdcZJZwc
vogWkAOoWJO6f6sT8j7vrNqufJ4HNkvVQRStqMQAITMLQ3oDblB8k3BkKpdPTP/0
B6r8jmzTpxt03p8UD0hm2NMnUxabWFvxmxpDuuumDA4EZQj+RzS08l5ThYjeEYQN
6+jVBPZJsRqPVzsS6BOg8Mzqp7WCeL7ZH9yHuU05m2OlbncMfRrWDtvz75AhJa2V
pkY979saZXx43lwXuH+oOmixHUeOkf+t0/ojTILkXIcfzxZYer/B83fsR/hQ7hO4
16QlNnnz12nRw1uToaO2hH6bdnZZJirB5DKYWEuMnOSpyK5sWdtpBYvlFErL0pLg
KgRcfQ3UnlO/1Px/Gezxsd0CxbXLtwwIvNhPqxrjfsyU1wTuT3HI7RyyeavtryTd
AwyD1+qLnahRFYL6YJpQPPTYifUSMqYyEpui4+UTa/9lRhS4Mnz2h+FiZ6mkhSmS
RyjOxUXO6rK4U1LktorYNx5HKJDPKmIiXQBHOxuCem1hIKv8Xzrjm32UT3BvGk1+
41CUXbQiJ+U3KPIv6BpMFB68KmqboitisSHSNYYk9n4H1tN58vlrF3E2xSGuSHbc
m+hN+WZldQZEWFZ6cSI9j38GBM6TaUMRmsxockVf0ttAfqhkzakY+5R+3xg7yzCJ
K70hDkKsYESC7Fmp4AU53/m+T4Gv9hvLwEQpsNBWQnTFRRKEsnsFR3cCiTC24fMy
OIO5FXfkvje5ufN1RDBhESY6rEZlVVr08zyYeDbDzY4uey+m0AS5JXSx3EfnTZYu
aXmB5rJ8d3W20TDmf8S9USlPRBmLGSdk72y82MT/9B8+8t4lvzOlQuwP39vTcMRA
`protect END_PROTECTED
