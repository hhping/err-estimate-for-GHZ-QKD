`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjapRyAlGUHVeXHcis31Dp13bv50iRrbXpy8bdKX1UJCdtNW39whwuDRHHXKJ52R
Xzp2UxgV7wLQLJKde0UXYvBGD7TETpqVH4DMQMMJawVMmWeyDkLxdHQnniU3i+vD
WD/+9pKiOaRvoWwunKJIYzy4NlxOhid3kykZwXbI96nwb1FiiDcsZpTPjeehAAfG
tf5VFs9ZfPGYh54OPuT7cZyT/pSs7FcvxXTfXO9eadd4HfvjvDxK7Q7K6/cdxPRW
qkhZ+7Fke3Uv3HesE8sUB2bWcUC7rZe1eqddGDq016Xs3u7MWmVum6A1PCNNX4BH
Xdnr2LGdupuwb+oDRFV83UPZyqnpCUxqUVxlFFpdUtXaMEPnlHW1rljY0iUvUpny
zKlbDROQs9epmC9VJnxoJghzXjW3KqtoIyDhARUMW6GwgdcXaKfZV7jzshs8S7W1
gPRap4G4510pbpJ5AstGNWw6BWXeQBOAMxOonnKr4/UXALlwn+5kP+eGVOyuSHQH
iQ/mLgts74qqiSRVlTf1CB1kgmSo5apNwmI+73il46UwFXQNo2NSITXdJx3cIsvj
q0LeBiycPzKB5hrnDQHi1ss4PlzBlDjevhupZmRLLOGR3edSvO88p1AjtaOxPhC3
P7V2SdaZAJSWPpjTVanKp0HU/S7C8htykV/9jCP4OthM74d/Dv3nbG5ilpQ32i+o
oBX7n8Mf/Mn28U199Q85EO5AeaDe3QV2k/2hbQXolIAONDku5pw631xDJqQeR5Hl
4lpptqmC0GprVu/6eBd07cqFINwv3RsMH2qxlM6ij909hXVLLP0Vqc9HJj3eajR6
Ejq9oirLZtljjMfQ+ezpPobA9OjYOz3MBnI1h+vlc0FQ91moLkCt3GTdsAeNVCQ1
Q/J9GI+TBiOCG8vCSBiLJZki/TOUHxSHhvshnAv+d+1Nt2KWCRb+BZXcsE1UbssP
kWgPeHGLhjr7VB5V9pnD+Okn4BtchtheI9GLv5DeY4c9MY6cl0vDCSAgwAYnumPf
hUyulcMSP/hVVy5iD50ZKWQDztWXyzpXnU6uu9Jt1U8rzQfmFUJO90eFnv81nLis
oxo/NT7qhSF/giUIZYB0zaFxNs20fCvF6nYdLRxhDtp5Yo4rygyFKDVpYr7nx3/j
`protect END_PROTECTED
