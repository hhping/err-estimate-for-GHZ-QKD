`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83QuAxe2Zu/n07dFuRg7dDlZjQLovIgYK+M0QZwQAL+OWYN7HjWi9vbzvDBreUSr
UWt+fKxXJJXxweNm1EsU6h50jY93n55cumcSHwEYfRQDy1I2mbn3rORCgEZ9yJQU
ktsWwl1885URa5vLGPUaTrykZw1F6pcYpEZ4ZKauv74Cq9NwYHK3oQcIiKHeW858
g+lqZmcc7v4Flp2WnbXLV0R7rD4viYGGxqTa2SEyvMqkqWQqdN9Obhgl8+q1Bdxh
9THo+4JMwLCzLBTXn1La1J7+x80RxXWL92lx7KLDy9gtsoO7KgN3ImXO7LEvxnBH
2/Mrz7d6rxmPTSfg91dUKWD0mW+/bICRRTf/s7N4kwneQvUyUkw8Csuchm6AJyRn
Td+JWWfpicXWdDVvfzlO9miZb2cSBNq6IMhQc3V3FiDHz5Uwva1Qc+/KO/ye1YYq
AO8mA63c7DoE+RUJ5QbrHK+Kar78Y6K5JNbEEiof4SjwtJIvlikbgrgaooGSntX1
imd8OotW8UNuxkgYHsn3Qr8mzm4IN4Vi1SuG04cmMfVOGOn8yFTbsePz0A83XEbU
+mD/+AbzYsYOEn+9zJ5RZdLa7nBpoxtKmXpy9Fd/JIXUkPMJpbZsm8SbD6980xCP
LdX34DrCGxt9Umni+fTCubcgXiihp9cl405VLiT6wJXuVqu1SS6D55HLket8KiTx
Pg9BjclwLCh1mLhy5QEkNHXESih5XenWIuG57AvTt9yWhKv9igTAzFYUE8c1QvKH
QQ/BjIKnS1Yjyri/dMSlId1oDCU+9nFKgVBJrqVdpZabWfGraxgwSf2fzvzudvTQ
0c8J48ZRQLgu7ZXnDn8u5wlSd2mi8b3603Lh5EwR9ugTVNNVbJrXQwx0uki1ECDg
66uaGKeQUNlZwjEH080F6Mz4owXxKgjoN+Wxo8PjGkLlYHxKY/yBPbX78Fs2kVps
fflfxjO8wkHAhOlND/r3+JhsBKjy0bJjclX4BQ6lzvU/ljQ0unsWdUBGl5aLB4Zt
M3JHZc03qAZPM5pZ4F11qbk9bQYv0dlQiaqrhS9fXHZ7luEy333uGiV3ViRGzho2
XOxVVHccsvWcn2uD53ig/VLb4WPwGEJ7E0Bxgeo8GUI8bGnOkFeO/2uvv6lf6OMj
euauCpFNhaUCGyV+6F+v1sKarcxGqBoAw0CHJMxb9ZfTxwjee+uGC0Ilm7J2sdeP
SooDR5c6WPqXFvkVQ5l//nFHperE7C3/aWS28JVclCeYUfi/gDxzGCIuWim6L8cG
bx7e93X5njLDIfjepHbR8RNLMCod+kFhW9FrYbXZxyEoiNm+1VLj0ba6ULiYrtXY
6Y1Bf810T2gGLwNSAt9FLkiygFdEHO1HmoAAtbEFQkfSK8FcLHU2UqGJowzr/FAd
y3IeaghxEZHgj8IFzsRhhKlYVFJxC40Ih6jAThHkT9NvfB0oMW1qyPav1HM3/uOQ
IxLMHSgPVJNSOLUCzmFB1LuuzaUrkFzvLeaWbvWVrjB2UHQP24V1Wt16mNx/Ks+I
sNtvb8kupMxQkCiQ2Gc3rGhcKGL2TmcT0/f3C1jvDiJRdTZWvO9TRqWFsyPF0kTv
zgBAFvUDPaR9D/tHqXViPI5XqhHQvjytVNo/Jie1MKda3qr3kiJwOmzFkdbb8VMi
wsSElRoLyTy0C0nRd2Jz9uSx9XXx9wuGVkdeX8V0f8mPKglnp1jTbBP27TLxdo7/
fBmrE0vEnossayUNbP33RazPrb76vVorFQV7N1oLU34=
`protect END_PROTECTED
