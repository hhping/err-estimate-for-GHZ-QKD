`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzUwTQmzaUiCH1cqslc2sufoj1wVxsUXyb/zmbkA4mlGQH3rSBbGsB7w2kmdmDN1
v32Th+tprb5ra1zCHCy0gOEF4aDbPLgmn/jfoGl0Te4z9CeDq87cizfDhXrsxqzH
MIfNw6qkjzChVGV1PKOjNru7/clWwdUUA+7wRWCYf6Na/7D0RSQwxS8fK7wx8mvF
Fnri0YCWlUrlySKDYKUzxa2Xzm/YC1AMJNXlLo37kM5n/ngzXFrfNvh/ZFklOCPN
Oph6S0PRyckVIlv+Dkef/U4wVhH58HMnEdN2eFCFQEfdLtN2JtrWs88ToaSOFvhY
vOOMClD022vj7kwX4ebWBiX7erSqT8DV2EJLVNH3kRXeI1puXOsLmM53awrGvthX
StqG/IFLX0jW12b4DZkp/OZYdfxUiJMv9mllkvqGgRIwfOO67rgl8DXMMhxOS9/V
nGGFesn3PsBP8i2dIFdSmAU1zsggRoVraEi05zc8EmuxVHfVYHzjR5RngCBoLtSt
fQyOe1PNfI3XPrepkkmC0J2o+mYywVbDeAJGB1wWWOLCcjK87Ed/DpQdak03P1AE
F9tA4wRypPUSgB9TtU9NxfcyCMZ53WFA5zMlYz1JbvCCTmJiu2PZGfcwBAjwBqrj
wJ18BzCm9bC1Bfj1tNeL1Ok1IAObt2YcI9RDhidjHeuVrXm3/ocgx/QlIXLiLXxo
piAg8yUQfFdPucAklLawxMmD4G2+ETD4Uz1sRthClUThrrAur/JeWAnCvCb7OdGg
LxeWCVvrjmcmo5385RvU1y8NJRF2aR1WByHenyuNHd6uNwqGy45fak39IFu3k30M
y3A6yDM/qRlDa0V12vuNOP1MHzdN4pHsrIa9icijU1Lk56bAz0PU4OOyG81ObrXN
U7vd+HX5a8oP1H3/+wUvLAi/k6EVZ8aNJGJy2Jr//oY=
`protect END_PROTECTED
