`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NALmM2pJvQMEwLH8tSDF7STC8UaJPGw6pOFpgeYiHscLIPgz+wFnQkiDGXn5HD31
UASF7o7L0yByOBCPQ5yHOE4RMyunXQrFKu9ipVJ2rrK0qGNVwa2E/oAwxyfxTwBq
mQtw1MYIRM4O22Xl20gAWSdeAk4JOitbFhUiqkFeF2Vooj5+HApTI1tuv1o+CskB
vKOQawhJdduMrjzDz9o1LutijSJ+uSLwlGf6uP7Rrh+yP2bHEH0Whceg3CrBFYlr
ddjs2jRRTTg2/K0RsVhW7kKAqRrWX9i4XVxpcLaYcOjsrBH57wAju8hZWxbUgTkT
mtFYZy+CNRJDCjMIjzlRM+KH2Y6Pe+b7yPzyCEaQyeGCJHtyz6uhcB6UbsKrRBfr
W1UGVYH4B2ZYzILoBmlE5AzK5KvI5/19dEsYxiDPsJ7viYVhc6Z3il/1qvcD+sHk
W4AZC617P4yRweum7vq6O4co5oxU+TEIRAJzfYrkokWFvxWGr4rLoRO7nYL3DWCp
cmnEOh6JbwDZlF8VQ3lvRrdfRsc3d/m3FSQT48OfTXUid2+qHVG1LMtrxeIbsEL+
plE/UZyNP1anNUCu9sgAHojtalbQyaqysXJqd1QV0OMLDofWttUgEj5FGTFgp/K8
lbpbLZyb5+irpPE83PfJ/A==
`protect END_PROTECTED
