`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1x2ZK0/ilwHp+ZX/TnuPoJUm6Hi+8Y+l2Wg8sTVctC0KK6FHVb54V3B1ep2Y0qz
X3jod0cZKHj0RyqCaF60LCI7mHU19r38tqw+3sidS699K/Czp2LV+O8/jrxQdujZ
uglY/xBr7cRHWn9glNLYZGyk/fz50+PxpUyxtP/VHf4B/kTTpy1xNtssl7Pf3cAt
4d2T2RGKmqiRaCOW4p1mgUo1ahruyA4ByCy5j/AKp21p9xHKxp+NUYjXR9xXhKFM
d1oatyIpdvZ6VZXA/BtnXmayMzxOo/rYn8IHIca+O1EdM3IOwuUUmSZHSP8LqWHq
lr/1e0L61a8HE9/DoUojXyCYI7na397VTdcwJOQVCNoVOGTblirbtWieBESsJdCa
iWeXhk1VXAIJgetduISoz3a6rhf6eqCEZBHwrxd1KdN42hK6tl9lyu33dvdQz7r6
A8A0x97Z5om8Ix70KCLmw1kHA0W76+gPvK/bsQYXYki1Sp7WZz+1WeF9G0cVd9e6
IRxIOb2Auc5mT3nqypLphvio7XGTwZiX8ZbVjnRsJYGWVB8bXLdKv3bklMqKEhqz
skSk/Yp99xsnd7wO5LoZEypjsZsPjsO4a8vIjz7wewf63Wh3/IS5gh0cbp29J8tc
HwVYNyh+q93yKUqjlTVsjarRIzDvMnG6sc6ybEtHEmBBKaCFL1GQXn3Hq7K6S1bf
W8kUJJCbSu3EqdxapHJFrFZDYKjwgXkOdnR/D06ikhUzAWjOJ2ij8mhnJa+0BvEU
fwMBr1K8/Lu0m+/hExgDOp2SZsFquGUbkgbt0ViNgFXz9LcbDzwar7NFnrcpsl60
WVHF5YHEZfy74f3ZbsCVdAOVXRxiDbrDCYYEe8C2j4BpzZinvQ95z9fyYVpGP2+k
cSfHVx2Q9icM0uLN9VSfcESswioUVHqI17eQaKhFwLeu30ySo/vKl8vDckdbTysC
bXdLRzhRP8kLqQeSgeZkXPyNSNC8D7A5Tvx9LX1yuiAM2aQm9aPcRiriSqcTJmtf
ZoyTfCyjY8UDZMFnf+6HZ7XozHwaYk+Ykxi1DKu+6hyScfE89WwasmmYavCR9T/w
7UmaauFMf2n8D9EveA0o4KXj+R0ojKTGJpP4nU4hX4HLmEp28kAGxMN3Zd2iGhS+
WOUx1Yaovf8aBl6YvAR15NW5s2YpCKRFaPpLGqMnWOSigX4AT2qpj2+vEEbcdgXU
cY5AqDRHOHs98PXOqajnK5xOxVcxuyZdOvqaiheaUaYILDo//b2usjBd5OfMTxO2
Z8Y7iNOO05MllfLc6fyCRPxkz5cp3LXbjSITCJ3jI2xzewyr6UQU6L6LIgBw1dtf
Bl+x6P4p7xN+gTuHZnfFwQ==
`protect END_PROTECTED
