`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQM2Fb4ikMO99iZBt8I8fiWvCyDQ3jpxzWUHUHcYLoSjw3nMqIpOWPlOUa8hdoGT
dw/keO8pb4XfsLSezHXMJc4EXbee11axybksEDZmtr0eqXzh/ddUYbemOrMwbx60
lNIbAqYOX3uVcaA8MSjAklEZTbhHWEtXNZ+wkE5wAqSgyFSE0FRpQVuU6mc0skIc
6X+8jCTDMeunQH22h/3uZF1C2D1pgG17rZLDExs4CRRZnMiZQPpmNqOo8reeXFCi
aJnpFpPgp9ufw8GaZJEo8RN591Y+Tj8yiIl/EXmvM2Y1mDOmiyUWW9r9mSvW9Gtg
D5rAkf1Je2miz4ZfwRoWC+eCZpfuhfF7+3pUCBj/KYCUs15PZNiC1E3iinKqysf+
asa7Cr9NNnJoU1cBaY3oj0ke5Mm9TdI0VPIZs6sqFEesVV9/p4sPlkvufxYnfJWM
s2NU+jPjLTc2hXJpcg7YjbonHjC+SPgu1PKXzCrSyujtlWLFQ5JaYl+dJt/Qsbpj
Fu5m0CCfdrCGBbUpazS1KIX6HRS9I1I8/C260U/eh7mjR+dUjArVgD9DjStfiptd
fcSYlkUOStWPkiwEtjvwvzLafUZErcdw3Cdr3Lh4QMXwqbK1URM1ou4+geN+xyTY
xfqtqllljW4skXUBBG00u1/wl37/TTucOa6gg+aUDB85+Qg7BQYFcngr2s5Ocv8D
FDw7mDNNN4+WTxMZSiM8bRDEtnoGDcAsypSjNzLCZQ25ylBwm5dlIR1GoPTRB3XG
81UV3GwndQKk7eC8fuRw5EhVqz1s6zPO8pwJ8hZSS+N3E7Ou++hJyc0kiWgZ7rks
PySmAEWwVwsEdMLe6RYKE3KIm/YcKJlVVqUJ6hBVVCSmJC9WzBg+7DDfByQf8nz/
ClzfgdcMYfK4NABjSjMF7zCe+Cc/5oaIae+40ufXx0ZXJi0XV7vUhrTA1GVnn6nb
iGkm5opdm8KGiP6s63b8AlCiDqjLK/OJFcWj73kTbYklZjAhHvLO39m8PaPhZoNN
Xht6608BV8Ct8cPyo7EqF+Aw/kG96Osl5Z7e+Yzymp6EYPwRMDN9PvFvTnzte6/1
jD9mYHItxtW2FjVvJ5BanFXR06E4hWeCkPD+sFuYRrst5lI6Fid2JhfpeE0IvSgu
qk1V4xQH4RnU3pYt4+SXtTcs7ToY+dMi0lJcy/uS7Kx+iR84x2HHFLgbhMpO+HsI
J1BkFtiSXqFCl6O2H/+c0sQLTScwJLAGa6mKPYhCRRHIhmwdH1SgL69v7lL7jq+0
ovru/AxiRmcwqoXmh76+XdS5etDvJeJpzhk8ZPaorLyXA9E7i2o0sZmwEFxG1x+z
8aCOMm8f7+R3s8Z4LD68MrXh93/KWytMXJ6GNhNmbeI74ml0W4zplBwJgBiRUe9+
n1OGXTm6cH34iE6VREYsG8mP03ZPNaE0BBR+de86G75M49YNemKaXRrlomBjosGa
0ilMM1gnMBdzsEkIKtSbHlQ0ZenQsFKo9NtoPNIk5cc5QArwcSOib1OuT+nwosjt
DyDWtCYYYLLbqm6f12idefxxjQERPnmbrmOcijYkwdTGJrlXumszPhGVaY6uN1Vw
IvKLlDHWgNlSCh4Io5kJQo5SOeMI0jF2XudyTS7iti/xR+9mdc3U5Vxjfm8NqADA
`protect END_PROTECTED
