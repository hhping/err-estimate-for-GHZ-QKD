`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JSPs4/xyBZfA9KmIDJjnECNRWn3dGkR/6czbqbZR1YdwDYALl9JBs5n+SwJQlfKv
vTOvVVMOeHDsOnYMccC7eoQ0rB655KPsTb+mBwK6dR5HET2HYL17VDP7q/RYktEN
DkwzOJRbA4GLxCz7JgG/0QZMWEcKF1H1zXfPKAYvtTVusY26IC2sWo47GIbYfeb8
rmVnVu4124D3X7nVCsXmhtKH8d3aFRythBBTsOwSVyGHmWfj0x6K9k6FhAAfoqgo
mvpzXn1/9BvchMHfNeqjWQrEKsVlsR/NlTSV5bGiPxAdjp+BjYZCcS5p/kZujUKH
YXnXg+C/sROPWQXQ96CeiA9UiVVYsoKWwusb3iyQCw9BM4MpFuCtGqD6NaZdqjoy
8v9YoEuk/xn9FUvaXSiVewlAha564jPzzMpYkayN9pj2zKP3J454WFrjyE7tyFE8
q3UZ3QSP4uLwbMUCruRKRPGA5gu+ngvEsZnBNbbVZuWI7Pywj26eHFwZBQ+Y+Zfv
xfYt8Qdxzmur8fbUdx/K6qquwLnM189N6gwVvGlmLYaJRnY/YDpdzzTqdQxQZCKX
CMIKFoXFuy2TtuK99TSldv+b5JaA8byLJQHLA4AMGbS63fgORhIwRq7TXxMG5HVN
Xck1mm6xMVf0DIpjm2F1qEqKcuI+1TvZg+kluS9dqb6UIesuFrQxV7zfwpjg7ZnI
agnAGZPvvQcGmWpLHjH+y2MD8d9ourES/JjiGcEaqdF78082JYk1Oma7oNgfg7kh
iQdPkmQzPXjCAaBKegdIz+5Q4omeYHaXb//OoVnEobpIMJmuBVTb9sGfLi16MJTz
7tZJnAjY1MQw1JL8MIhI3DUbGyZZ2dc4J7XmDLNg7drItZb1XS3wXbRtlDilzmgi
sFYP0saGeqE9V+22bCyR4G+2U2T5EzswT5itvkH5eUf8DU1rphww2RbLbaJkTASJ
iO03wh2ohiQow6zS4E1j1r4IoFoI1SCD1XQStz6MPIWAZ6m4RocU49dvijPLJyqk
`protect END_PROTECTED
