`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLMpEsYwJlO6i3710luZoWUHRDga6kxu21b7dWAc3IVprbYyeIzPKeDsQphqBGju
c3eOeh53GobQdoDG2qwthFQypG0a+gZEviJC51CNXbVzJKeq7vSe/5ndtGibbbjk
umD9hP9Imd1xK9x+3DvSAXaGhOFrcPXRNOv2f40Xs0vS39LFdZzsRwQSwzwCNNck
eN7ljrHfWYYwMt/XHu2LJSrnsrNFiyvZZmek3Gj6lxdTXWLLPk0Y+4jGiHXT79gO
InyeDf/0DoputupI2YpqpCVSP6/HN8ZrkilPidcm3Magk3G025TpxyHn5zr9b+aE
XwaRXL4wODjKEfoQ/33uQEo9DGbG8OdeT6hjD0fuWpBoJA3r/bHKLuCpEHOiEfDN
blnEnjL9cq/jPEkPdgFzqCzrLYb9+foBM457CniPfaQcHonTfgm1XsDAC9oKwPnI
6ERjnAAnOzfFjglRFv1PwQ61bqN/KPDBF0UeNbUMpq2UWyvWztpzbbec3tuPaDf4
hZNYi2oRHv3CAILbSbzYqqqXMc7xXeA4wVuYt2IGY6GEFzynde+O3QWAbMoyPcuB
xeMI7dI0Lhy2+tq0Fpb9sQiU+sfxoCWxl0BllGR4McMyhwQ98eSHo/7jUiablUlP
TRVqzWmfrB8c79hW6xzKoGRboobz0pXDFwWHdVE0VJtdI/9xX/GieVxBomciGw8e
RPT5LEqX4hh+e9VFoO3539iLBYFOazY4IYZO8nKjmuKxueZ44thFC+ZsUq4mvmPT
mnYDcZmnPsfwJwDYUsViPB4YZgn9r3xmsXmyM2nRY/38XJs6RZOnLWUmSAHyqCgP
fkRjRpLgXF9P6SZ+1LwVZXoprrVOInCnwnx1QY+nrZhZ75h25FFeg5XLuYZwG+O7
B0Hr/SaIV0e32na4Y3OTNnMZC8g7kn3vOLBRruJW9E/1BmtgNqa0by/A1NET9kX3
pE80CYcM33pyA8gYxx2Ysnfbt+leCnOSDZEWMMtfJd+QGl/Mrl2PFG1MzzeiqcGh
guecXH/AkImxLmc7GxdLyyNQspFaD3yW7la8vf2Atyxnqd8AZpUEEycnoHWIRNVR
koF68dS+U+6iK2ozvTQ6NuxsH2x0fYwIbaVDvy0OCBQDKIBsoqXIF1rjx+bbhdgI
jKGKv7y9ldXbPdpEbKxIyOACpLh+FQMM53X0DgiUCD3hB+UY3AGdSh5R+uzFtGsP
ECIEYBsjuEedOyFg5Wd9EUwFAJ0OfE0ksSfOPqouk0O/OKR/DPWxupACVUSMWGBT
dpmmxzfceROJapN1aghJcgIc3Hx2yzAiPj+rewyz28OPzdSYe38yvCEXt031CdQf
+v6TEf5rxZL/Xoj4Vf/Lx1HR+eRULiE0nzVSCwOX0239PdDvsBMmaL+QnPaAdCaE
6GupYVm1lYpDy7aFlJcPo7Yp9gUAgxT+dJy8hcQM03vKwyiyIoDru6zvRojDYVw7
tb6TIDrIzStbmaIIwcRNV0FChiVecYIkV5LBUAxtgwD1vk9gCAWXyWqpCol7/SyJ
cV0mT/vobaTeTAc1zWQ6OilLRJAHLIn3ftGQhHaV78fB/TBNdKWVWpWllUS6QK2O
p9ANG5bFKZ5HcuDdMfMT+YceFGoV+8JomRNIKRNR7r+w/s/5z78XHa8ZQzyBSwpp
Y0S+D+kuUIDKsqROVTjgktK3VcgvUwpji60jpXbYDLL3sucOOzmPxZgzUfxaU6dQ
nv6KLcTGcYTiKOpHIxzljM49nQZi/BFi8J8kZy1h/JFfJCNaowOsKSzbCV/3HJkx
J71hsPMMFV3pOs0V4mgwv+q3LIZLkHkWvPdyrqd86AlQlKT7QHscTr2b+n85eVy7
Y65k9VHGgy1+yH6fiIPbWjXQYWtcD1ZDdBqWDaikx+3667p1rndUftATkg0wDYGP
KRng5sinu3TmxnRAww8C3X9PWEnTMnNq2fx18/K/MH9siQoTDSuFbDGVXB2roC8a
f6GSPrnrTSB82mB3HHpq3RkGMCZfzoTwf6EzPdm0DdZ7I0MAlfzlK/l/kH7vTq1r
aQ/e63jvnWSiw9Pi4oU5EwUxcrVorT6SYQQTz4Ncj2it8s5KfhLG1xzZsCweuqC/
I8vaiAbcXKj421wyciyZOGvLzWweVhmjIQc15qBjuFlKUxNdcces/EtTHNXs7gE2
nq5p5tQmypKvoxU2b/uBLL7vH90Hwc+stGKS+KIKvJqLA7P2U3Nq2wDp0PFlUkbG
890m596mECYgkh0ACuDjNEG2z5QGK8Om5mXHXVCM5xvxt9nwAxmKS1Cy/Jik+Wwr
e5SP6h8lzDUhdvLR20HrZqqQqEW0OGFCExmpNKe2lDeBwdSyfp1Lp+vOfCf1kymJ
a5Nld3D5X0aTjnqJ51o5Ec97GG6jDPu6TxTmYYpo8XTyJP0CfsrweXZKtIZbrd9t
5Mh8MzKpHQixL6NLSpLeVzvXzedBcMb773xYP9fncu3KtKzJsM0FMpVStrbbblgA
MYa/BQKwRzEaN3KwScl1NRquS6arSgFTg0u5uroBrtO0tJIsGdNDNha5hS5wAhXD
XYWyZeDtnieE12Ipq/jtYwDE6cw+N5B+Vj8QCXZLW1p2enIAm+SssquI/RWgpfN/
FbUByg8qOLUzlBkEqtDICsjhlt4gMWi3CatIuTHGmHQ3Jwgl+w9VBPdQc2x+TxTr
dqeSrSY8DE1m+aa/8C6d/VcnrBnGTc7BpZZlXEZPpS2W8v6RuWYhspu/d/QHq/vs
xq5b9OGrQbDJu566HmJ767uWavTJcMV7dUKsXIc+O5fQrJxTr1XurJ2cRYR0f8v3
mcrj79BPRshlv0GD0gHHgMGCBQ0nzLlncQUHB04MwJ7xrNpvFED7G+m7V2L/F1Nf
fF2cqPf+Ico5xhOdFLxTUOU4+Z9+PwTua3oMHXaFv0BCEmzwZaN+dQ2YQNbxlBkD
NRw1b0qXvACODdlsm8dDYb49RA7Z7V0HV4XEand5qpVYoqmHCfoJQJ8cO2ERty07
+7h/Q4B8TRWWD+RPUMXP4Zdpd/ro0Ea6lPYptlj3tNDDKBjZa4Q4KUF6FqafAW4e
leLCAx7dub4Mz8ep7JhpofpFOfp4w/uwlphoAnYp/f0izQFu5X3cdiG8UzGzzRzt
uEbj7586MpfFdq/G0rQUWfw2LUGrpoMilZH7mpCzEd4fxD3tcbzZY6A5nmHlpg8z
9vTBpfW/ahHctYtd+ILAWvbBmO6QkzcAIu+TkKjdMdm91JaH6u5zsC1Xe9hfReic
/8gv6jEfhS1erPKKXW5pNeoB+oWOPpemNwBCpLIihwaKkRM5/3xV6wzuZb4LEE2v
Am/QjJaqGmaSPzCWQg3I5F9aQfxXthUdfT7rnrr3+XyuLR4BpmTvClkEnN2bRlCF
1jAOm2fNcgInfCNYu4TgF721jaXCk+JkZzkE6LzaL+rJdeBCy8tY5WC1Apn61365
X6Q7sfRYV/wGlw6/Y2fanHRW0VUCZa2XuNlBdgFTE+Q=
`protect END_PROTECTED
