`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUkqlwuqFClWCFHI/u8d9LoLwg6DuIZvNITrO+cWRjeEvV356LFKTQEE2mt2ibHV
LsvPxUmZgypyTgUZNcg2cOkuuv1ZlC/t1lbqkiPSqhb/zcvnpFi0NZdYk0PBDzz4
DqmP10NSmHP9FEJb3gjMAGJxLiw2Kv6PEy04cr9uf5ZFlBLqtHqw6S1noz1A5VEL
q86bA4Xw3AAtZ247vMc/MxB5ztS7kHG25WnCmhgl4X3ysE61zu9YUY8DwHxMABWX
tpWTN5jNKYt9iiA88XVoBwH5/41+VMQ1exRMBeXTkEFO94X0Ej3EW67oJjjbJIDv
qRXe00pce/63/WJxQ7DeLBsL+AdKHUg5XSi5z6dY5dhmRfAfWcFXdcqWxWk2PiFL
ns7UZugvI5r8wVUmP/L9rXqzjR2DApFLzw6GeCHtOo4RLY8mzEJM6LZMrPfBICAz
Kl40ppg/Be2E5S4OprdY4afcWuJBigyqvAzjugMtnTv448OQchQM+cdnlCMRP7HR
Rv1kXTe4DleFvN/zOf6Orlkd0EHhoMgz+QeHknzjHeJNb0NTdCYrXFiqDpuHhL0D
XGLoQBXuBXdUEWfVZnEI36xbmdQ/+f/b+h/8/d1NeYr4j6/Nw1bIOsx9NPoxxhTc
o2Zo3sRkJkMgLJkILbStiFjtH+wPfHZrIoT/OK6OFMtGpIxAqKaiOOaVYe2frE+N
rrQMsr03grPtNrmVlJgFaLNGILhn8+F6FhIuLQyjblWwhaCpRQSywJzarFJLX/st
o+UiUOHW/9t88q+kDwE6SQioYZqA8GU4/U2ZFA82SGBMkWelDtKntzP/W2b8V9+Y
M3i/bxWcwi87/9w+x0jOdcwd6/qtbQX6BiGtEN1lzfatyIs713TRZnXEc0imcjK7
oOS/U4uvNX/G20N43Jec9En93Jet9gQDLV/jDc8XBvI8gKb256Tnsf+L91qXRTMw
T1Y+Upga+dl4fzfAzoJ9XsxqW7dlGFlYSlJehoSiKSKbfjikljG6dj7jn5GunDHH
FkEH00UPqIWozb1q0z8bM78vKruTefEbzNVjn3Wn3/WdaimF9FpYEENPA28zhrB3
+fsjBxP8YM1PZDNTIjx1lgprFj34Ey80TPNmCRRss+BpqNNZz87kXhjPSpxro5+l
dtq0Mp/Nusqb42RFach96IU8JG2l1FfMOiZe8mn5Ea/2r5WmdLWYGLZ7rQLaaxP2
A9HiKAp7eRGLhvJ4NN8TswNJtRvjuzSNbZ1aSw/R7yjvQDk80R1WCqgmjNnpSPZR
R+ScUDcSFL8j3sGWwkDanwHENCMoZZMAOxq182Nngii3qii6xQH045JpmeRN0f0l
ykkRiXawUSnrxpsZGEKnbkXTpEIcHPvgyvzPKEjQOIsc8lK/5hNudOxDqWC8SRVZ
Sls377RLQOy81QlKLzfuAgtc37T4/lt8QdJBs2yR2dbKuxlpNU4IkUvTD6siNeQB
Rboxh5GO5VbaMkXhj36eGCI/fL/E+71LLysZ2P3JNrRNDbmgkuhfw6R0aTP3HBGq
+SEI+3mv0gGneSp8jxkIwFS6GlkWmkaIDS5DAOXaiqR6+xdReVK0VlgGqDnTaWZL
iuN6Ul5J9lGcdUCbKazQ40WMil0nTUTznE5odEgSIYRmk4vA/IN+NPk8/lxWYHST
DKSV/Ovl090fcPaE5sD9HrsCtCzcP/hvW5OqTswuJk1XV3BTFGK9plCFYFDjCE4h
QtY/kOa/2nSaF3VKQAPbcmtimThnVFxa651DwrH/x4Wg8wIHsELtC3VM6kqM6P5P
WjVtMe3Pv30jloxcTzS1SWpIsZcca3o4rRMr9k9xVsPNQcUE+tdLZ5tu0KFAZNgP
c42lKDeV5nZQIJj+j/CoQi+zbhLldabOtjfhdvvUyzhPUwpR+rtvYq9dp5QQug9w
XAcdesNAvhyCTayyxOnDEU/cntmnFg6Dca5Cc+YbI36OkCUMKAMsGBq7cQb2bPql
/ZUIv3t1FV/9cao9MJalfDEN6BRagXpN+KPo5Gyp8uuXdf0mnjPsc/xk0Xanb8bJ
WIy0GUjpVWAOFFx6+5UZ4WgJiqSs91F92y/Tk3+76IVVHvUNjRoqS8vdnXC05Btz
mkJSHO8LS8hkHX3cHgrMBnHJjpneCuFT83q+wcarHb0+sgViJKINV/vzgDMeNf9J
`protect END_PROTECTED
