`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMahe5/HzaoH+IDRYPPyCQcdkT8wQFO1n5eItwfKsUQxxLYc2WEsMD0pvpKXUR7O
H9WHXDw3ZRA635t4TyHSgdTaUgKfyt5dr4mfssEX8TohSViIweYreQnpIoCUFdd8
bPRHM6nbUYKZOBxSeu741n0VgAQaDqEaN5e7tZxMZ2HrtHFeJZfthZ5KDhdDp6IS
hhGWUApXaxeIVygxGAjbxNuQRP2/Bu78Bf9aGn3OaX+McPM3kDAetWx7pxS9KGUI
4MTCoISK9s2sdFZuGsRBoMQRIbiiRNweCpG1wyyzvVZSrG/3mlapSYDluOl59R7U
2O0nbXKW1FgS9LWjpBQuWGitACeM2m6kkQpVXXzoS5muVO9BMho+aAzsqMso+Q4X
rBLLy+mkqLE1mlh+aIaIihwa+VOrIUq+yOtKxZaG9ogbHZCB4/wX8W4ykJ0N+s5X
8L3uIh59mknwYNEEgm9jKDGqdMVH0JYH2XFheMsiVfi73Bi6mLIxtxyELU1gqv84
rwpyuauz7UAuVPk6YWqD0DRtzHUl8dG66W4BOLyfRukos/lkrcZw6ifqD7PDpnC+
`protect END_PROTECTED
