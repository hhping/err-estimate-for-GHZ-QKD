`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHe3Z0XTjiKLbT9hOFkUV92Gxj/C0rLmeirfW9k06E45AYadb8TnGPi/UA1rHNQR
47tO1W8y67n2qrCNQGWwpGjbkQ42/3iCiotvaLWoTnMziTbcGFoMq+ySkjRIm8po
I5hin/JQjaaVy/8ysCt2JaNaK3TRlST6JrDIG4xlJH/hS0Uqrk/9sGCuiFfav6G3
cql+NrsLQpO8CCT2ybNQLU9zhDfnAlmVEJFNN6VBbIhb1Y04Gyb/83NIdw6nky9c
TuRS1TkTBsu1uWwBqFb6NTIxFyVtC3e9wb9ZqRryEXc5Py0GW6pn7a/fFm3l2XCh
4udykH0xioDWxyJFasrfLvi7akbh7axxr69ha1yHSs55PXhYOgbph8hcBmWN+w1k
AvkH5FpcDnatkQnU1bmRumIBDCnvb3DbrsWG+rdw+tYYKAD5zrwqgftAqF8tafOq
I+F+g8iFavAok4aeTgIeAqV4PLkgWwk4tFTgWp/NF57o/lG3foXRSRmFvczvMTE1
ALK+zfmbdgRj0iJ+rBXCw/t3eNZJqCdrtFC+XMsZFsQg9NOOE2bk/WpdM8UgQZea
o3TFMos53tuUGpZIrKgoiuqnU0MJHtHqviQWLFPSZgxeFqZuWxctEDb6l2X/2Kbg
S5xNOz0k0EVL4DYYaWft6w6lou28ci29HG0xsBc1vG2v4zPNMbbqw6dUHv5Ray1N
378TBogRiCXdmt9LT0PDhu3u6XJtFSNrH00gU1kYgvfzm/9DydG0/nXjLG8k1cEk
CM+1N8wrtdATHlEb29I/66tYjy+92nAvaDqoUf6bF59kohzL7h4/fV7e4nB+/Rn6
INgJzz2D7jKoT9sPVF3JyTsrrcpTXhv0piwA4sWfenIkcOymoxlaZqZBK1NuJgSO
yE70tN4tXqfEwNsnjKJazuHUQEU9JhH+Ka2DTfjWCTH+IlZfu3E+PmZ/Kdzlm1bX
QOT92AKyDjxvA128JupviA2m1MjrarhhrOfhOcDAaIIzzSLthtgj2uuuppYKKChG
wwB0PhOZzCHA6ZyW2+HkvpzycRmkXGjeNUqYkhyrj0mDNQaLYBqqro8NIFoplPq9
u9IxEq7mpZslxR7JF4c8PJw0gTOuIis6cdJdaDn4OQN522LCedK0yF/YSkWQQaoj
WJ6cIpjlLZDz2Ilz3W4EjmY9eF50ZU2eN8LqfdnPRM9F18MnIr67VeERpz15mbGu
nB8ocAB0twrPdUb9m1u+vaNipxc1In/mTbFSLDln4jMAkrAS774QkQvzmLlm+3YG
uYDvdXDLIP041Zq61eWb48gH1j9GurMWaY/hzCe79ViUZb1HcprX/6+h7I6gIsbI
BvzCa/2mrzfWDdOsh1dli+ztev/DIUKeIWbXnMZHXTAGzVyB/HWPbnoDLP7Xd6L9
pa5btpgObL2tUlgF5FVWIsTD1w+7jqg9ydN1qsKkai3I942F6glCkkm+nfWLA00B
CtB7f5HRUPrawAM7ffZPtQ==
`protect END_PROTECTED
