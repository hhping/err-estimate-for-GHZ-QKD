`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqrE2hhlm2FqyArb7SvLJqBtRe5GBhewHGKQ48t50GvIDnPt05r5c4kQvH1XOJC1
Vk4gxOzRDM1zsB09FN2einEI7Alj1ge557vr+f02gboLMjmcdN7qE19LxYkceJSa
6UsIRhf+HCHBbCnKgZuL2ivHupc0oOluaN4+Wv9ElIA5kUqboEIvqSi6tjcZg0yu
Ge36EnASgDflPZrKImGae1C2lkxHHHpytioQTVeip95Z1nGCQKYcpTFD4EWKLI19
D21jP4NjGvVwZyrVk8OZkccya8PKtAp/+9iwCS6m4zY=
`protect END_PROTECTED
