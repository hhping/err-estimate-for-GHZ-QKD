`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
inBet9MTiIsBQT3PwYpWUqachE/cu2LS8oSGgQXx15D285SkY8J4IWZ70f0D/KaU
olohiB3ArN8dhI+SwMUM0XG2TrgRAboxqM5OiE9vMf8E0cR+k8YYZKnt5EEmZ2q2
BHx5Ag9tMZdLcwvhXq033Jdyls2CffZIwfuu0W4i+3j1v1TGXZ1b/lEqIQ4z4Umm
v9VqOfQ6czVWvjJ5dCCh2qx1Pmjf6EqVShHr5kY6ZmaFGVIWxziRykoZ7+gp2VWW
fZL5oCVIj+Qwico2TYNbpUBWQanDdtw5RRfk3llZLcFhN3qEKd4B61rerAd7xirb
bIWraOKjjwoyWksqoul5rmFOrYxPP/mFQOMfUe0T4gpWbXSx3RTKunfEgRe8mcpz
AD2bcNBhI6PdFkpt3J1sxvKPFScDzrPsGWFH0aEBxIHd4QztS6t7pjeUPG1Fj0cm
2kubk/w4qOlpop83kJuhe4KPGcD7jUKieZC+JPUbR09WvSZpjWYGVUBWZRDFatWv
ZV9Dd/o8ohW395A0OlMKEaPuxtnJwJtXz1Dx8fcpR8pgYdIZxrqfcayQfigRclSE
WIbEBQ23JzwOhMCfBqlWGsLTWEtEyS6fHZrshf1lJK1CZ6zDKdN8zEHWHRarSac7
Rt4c/9VTfm+/Xmnu7bl9LGjFYOa3H0da5ChNxcF4BaY=
`protect END_PROTECTED
