`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4380HN3yctrczeA0AMO4pnGSYKwVIf5Zl7hl3uf1z7um4oYy5WTuqC9Y4gsuI3y
Cjle0rLlDQ/Wk99xS8KILpRTVb1jJ/GTiiZ5ttxr9aFaXJXvcXmcjRntYv0aU8rx
XP6gTglCbCZ/yRh58aIdYoMJ9ytjx8dgP3CMru2aabUnfzTnjgDYm2FCVtz19cDN
JOVV9cNTgR/bRr+SUb/A3YFvG7hdR429dtjCTfiR1OQGl09wXv3W5++o+qRsYon0
n78RzhCTi47kZYcFIhcAjLS6cAUgS7XTNU6N2KB89PE58QUqR8VsUEZjfeLp1U+2
5Wj5mrLwhMlGWQskNFU01Fbn3KMyYymFY4mqTWoqN1yZqgKRT5vT7LUR+U8OnEzN
/++aHskwQ05dFle3jpDGIXm+WZCnd6+smL+5xPPV04TpnXIsEPQp7yM83HhlZpq/
Ih3kVH8e2eOyKFh2EvfqqzR+SWgHgHWpegeIGFBOsbqRyBMt7+D91O4a2qWzUm+S
f3tfr3ebT4vS8SqGkHeSsBtSguvFPQUmXJEJQsi9WBgBX4Xh24phAtEmlHko7RKB
T+b586+S7yASMkEVkUl7gfW8YUizMmUJTthCBS5txQIADOW6+Oti8qCZ4QMK6d/d
NGRzK1iEbWKNY5qPaXfng9ngmeTlmo6ldiS3cYSmoXbAnUUO+ADaNyyr0zXhIUXi
0ADxoWEQmgPntw64F/49Zg8e1HafultL/SdQviVaHe9rXlHL6sXYcXzgAvIf4Lx0
`protect END_PROTECTED
