`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+LfaiiO6UJDYEPfzMR7oCjfWYQIgGS+dGCL+CxBbQxHOnfAwSG6ax6ujooc6z2T
zfeBq7X8txoSzDtms1CKDaasfk7ZzLUXHnkWJiuJYjc6Hz8W/5yyUs9fBzaBDUvK
aqVmR7F3/4aXyCBKFxdxVq1VKzNlzr/WeS2KiGuWrCwgq0YrmtWcFh5QnWVh4A41
FxNQxQR1LUk0JAKMo+IcsIf+GfnDU3U5eUGS52Vsj/9Z+MY5r9JvwVGhinuOQqQb
xOPN2m6NUnCdgpVyNc6YKY2zhNWq0Thwn0QI/EpHW+bstwP4HCuab8WQFG3vr8bB
unrU6nNuKzgibdcsXjqxEl0qpyWENVsSl/IdtzX/saF5xCi0zK73q+jh7F4Y4OM6
xTsi4lvubvIxsosd8SD59A6RUqAcY5yEqwXnwKHbiTBiid3id1RMG4uI6OUW1aia
Rm3SLMzVs0CbhjnfMzVtsSYkdFGqA7CfMnzuBHs8bwYe0+gOzJlqbbenOknSRG6d
JalvMxngHHQx65vkD/MkN2n6RDSc/lC7qJUfhoLvgsZjVZSAliYYKTZltbn068mE
sCFu5pby5uioDSM5xN9EGFTQsL513HPvN0PCLx/PjMJQ1DPfuU5WRIk7QSCQgqst
OKyrtBjXkzfTZFN1Om6S6XL+PBuj6F+FPvMUMrAr/h7aFHEH614cdq2cOMIqKkfP
Q0MrSH+cokkrRtxGdmET5hPdpEXfsYncG4fRHj3pWLTqGCfuZvp6grTV8g2EGpnt
dCnicZGTzc7TIAch88s+vIkR0uxckqwYr7ip5S0FimnH+7cHqu1rc6eRuPz1TbNb
hyx5OIo1dgvt9KSJJ2pPepUBfNaqPEG74nAfqV2qDz8ywNoGR9IiPYsYUeMrDN8d
AR02/mY6OdEPTZXoz1oxR025Ul/l0iOAxWrBihe8bsBpLhaIVXWDD0io5fF5weNy
uyXm8Y6PyVFAgipFehfzKO/y3actyxq1f5kYf/QC9JTnTWs9+d7TZtx1NOS0wfp8
gxY9gI0iqxKE8xPPNPtJiKvt1XnQ99+APluiFjolfr1FRy2yYfPiCxvBdBT0VQJC
raIbHC58CuWIkahGI2JwCc2kNFaqkNJzphfXNjMFQSrGwK6N1qcA9n3+d+zHq26z
/5qRX9aLadbtgx+wqwuH9xRdtm/L5DkCmp0SuGr28/MrpYriSJSBUZ6/WG9DK98a
knpG9F2OhlStAct3rXGsbnCNzR+iGVG+4XlgetwbxyNYuOzTiEZqoLaRJYhUrsxv
AbGboPv8u8CV5rmMZX/rajnsPdUYM8OtozSlEo67MicOPpDtNGc3V7F3RaeffTbZ
0MM3EC1mcQL3sIpgs3Sk0M9jtZ0cPSS21/4ME67hoVLdXyCaS7vlxZAfipqgMvdW
b1zmnuicQKIrBllExinyJocyZdTaBh5SZiSeohQq0FH5CxcuHVio7VHbGx548m/W
bFkb5YJlrmqM2/Lh2uYMWqHCmZMkmtYeA4Z4HkLJE+lVo1RP4Y+OShTK0EYR+WJc
dky+SEg54gjdZrfYb+Ib9vv15MjhJaDRaTwMlvDZBerHTWeMX0bPiqvfKhBJE4Qk
jShqaOpUn0VUeKBYW41cDA==
`protect END_PROTECTED
