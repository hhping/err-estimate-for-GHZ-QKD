`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kU4U+/WaE4qkLua6mn4+qfRsNwA13e7vR7cElksZAa0YFhPQ36uodG/zLKCjRAo2
nNgxrPVQFCw0gNn4FqHIoVaLXprJ+PApF6w1Lxup8seWzws6RqiLTesgbddt5WOq
f4FZxy4K1jg+vcWsbCCkwq09OBdFgsG3g6gxGPnMnlwiXzk/Dty2mlD5ltmeA6VE
CFsWSN10d5quHycbr8+MzbSQMXdRpBsRLVn1SY2o/kvFsOQXRjg5ZaMxPCZzrCDZ
8/ymB8TXUwrcHVz0Q5U2FgAPdLwHtVqRk000KXlQMVou6EjsP+djLjQC8RrdDvJO
+4roGDInI2PQFHHxb+Xt7M6HK89heBPlcmP9KHmHtBUY/gRN+OqswEFWyR58hjUn
vucQvk2FflKpVFi98CTcMp2y9SKaIe34SWu8w6RWpcERhe0SoE/hV3ZlI9Z0jl52
YDtjuJEHoaSQqJ5VWXkUTCRt0zZ/xbkm1w/tSpTueWoDcYQGkzXLLa1FLQEUXn1+
5iWibHQFnD5EXQEvoAEdDxdy9LNgGnpVNUftlAKqJaeAO/wYKfJpvyXEFq40WmYF
1r5pcKEOvltws8S4zxCD89IeSqNMCwTHQth2+wgzOVS9JIR1llsSaws7X9DgUv/p
sI4OReIYL0o6HtYRJg0Tnz4SYAacRif2TMLeI6ZqMtULTuLHpjQZz2QPxwLt5Gpt
lg0MH6fuZEHVGRdb0ajOr3P+AjXgt4R7gNKW5iTt40fIqMrLagsEqlYednvZYaoA
7uMmyW9pSpw1kFwIZYhVWBOycVaJbrlrKSGU+9Adp/x577ogf/DVTN5xOKDYBqTT
IjkqziXw4yE3RqPNaiAJWTO5461qciZiZ3/0WHvC3urfewgmFG7Lu44M41/X2DK/
ulxYspcSTrirfOMXwxE0RZtRLzFTziK7wmI6wBPUOT086yjftyS6tjMznSZmpj/G
wuHm/0Vi5bkWMJN2oNCpp3tOmFOqbuhZW0J+aWSMAwxTw/kLF6Bpx2rFDHMEasEQ
bUsjkWwEToY2rEm/ryXUIv3wfkF+zUFyxx7myBiTflRjO8xHAaqzSGEIU2IhJXhK
CWOSBnP6Kd/IMJk40A9wfI9se5BclX7QtCVdPgqUqCTJC0gcaasFgxcdv5k14/77
GrBq9RpBFWAS6PAwPMNkDiDkmrfzgxB9XbjhC2vBAW7NeMOa0ckedxOS3hTV9TlP
QMc5EwnBnng8/aSmHQTiUibGA/+vvBu1DN15gZn8E9FtKIp+xFLuSiuqkXcldA9s
Qe/7fFE5eBTGSyiqiNtvODWX+yOxL0n+KdQXauuwXNH9OsI2KmNdDCBJo7QnvHsO
y3hiTlw9vdqkpxP5RqYm8p0lZZ18alBnM695Ws9bF5RGxMM/CvpZvxwosvwn7URf
zqcTXp0fKfUqTwM4WOBIGVpm5NBhbvuf5fmfnAhcfe02wV7Vijlokn/J7ApLCZdL
JAJNmxF7oEzMILyCkuWP/ZNDt85zGbsWlRirg+/JJYr5zduVqovtXXTdWARRsUQ3
oVR9tit6Fg+fmpgA4C5BwHG9SP8xGY50s4SnDJHf+pdSIyc4AfVp5cpqtn66gDha
a4kNA61CVspc0O6P24hYRKNDt9GMw1gA75OKU5OXQlTT1ZVMtMUN/v3+cg8Ame/i
pqWAu0zCSOuPSTmnvjebbs46B5/QDtBvkEbvy6d+NF5X8TK+2lAMYh+2yJgt+L/a
IbRiiUAtp0YCh5Iuio2FS/ST0r6jqv4TTDWIU+FqdsdtBtv8BacIQeJBUMK59qO4
mtoeebrfevynN3syHD3wTX6F4TWvM/K/7VahPDhAUam5JMc5hyqsunFB84V/jewq
1ZiGzmujcyghus6Qc2bU1rniYas+Mx/zm9EsqZ46zgqyZfin3ZlrWxhoS6tjEYN+
qJv+2v40us3+k8A6f8EPqrxlGp0jF2yVT5iecerhXLE8iZa4Vgkp5eQu42sQsG7n
7hpSMmpxElFQjTGr5My6leBgwVywyJySeRiei+id5dSUsd2IcC+qDAxjgfCEcD5U
txR26n9cfiHM3Gql1s3PuMPdf2gSezsV8ZB60fw3B47W0HVuLIcW/+ffSCgx5eTs
ajX33wPBoy1jaljjgnSD6ULu2M6sd0CGelk+H4UpLR/r3sbC2PLKpDdlcCvZdO4J
datWnSgDOPqfv8AKJ0UhdASdeCwey0BOWhQ3h0+hvlSbYMPapPZCpfq4RDzEYTTN
+arqkhCbY5T5m6QghBHCAUxMyEiop83mUTOp0c6U9v0mwXoec7I6AFnIwToIQeMe
74DGUEqtOCkAGZ7Tke2tBspqDqfrzoxan9U8dvZC4Wxtp91GwrA5vELpKR+oPuZE
G4wgf2iH8/R8LyjlZcNRTQzmBL9ORFyuF2S5RqG3F33ZCxtkAe24+ywwacxydfp+
bDj0XCjoYNPNxv75ioCCdqVqx6RJXo42MuhFtSa/3j9i+7tBpor3PfjjbHGyS8dM
JYOYwwxc7JF8YRdwK0WAC7xMe8XOIkKny8bk3jcsr4w8b7pScK9dhv9jtqsbtlwN
kPzxS/tQRfMj4wFkB9qzfecfHEUwQcBgfGwG6RiuhFmDQvKrCwj9vqWofXILgcRp
deSbnJv9m9RlUwDGwOjLWwsftD189xNo0KpZHd4JgYDt9A9bzJaSoMAGqV6RWtFM
Mu0CSsadiUKD/YR4HdKSy/jQH7e/ikNgitxf3Cwf7ivE3B9d9AojKGhJyO9aPl9a
H4+2KPAEBLd2gwzFhiVeDWokrpDGLYGf1pTbqLbbOd1fYtiH29AV7rLcfbSJk84p
UYEzL7gQKpdbZtKgyTrwO4XpmSqoo248OPEKhgp8f5aSpx1usTeMeg0SOm865X+t
O247CM1m31LBqpNHtb6KoR5UpC4hmStpxOCZEiY3/9QEh43Fky6XeLvK2MWXnFcr
M/bfTzQgcusFuvMBNQM76si6D0lbZrtoNUKuFEYYkm/KzL/VmjvxYsuTYy9PfBRS
8etzGGk/8irqloUBD/WATlryXFHKpLcX7I1hhzT4trqv2PGdJGknhBTj/D4ETcsB
/J8v+1aeCRC4jfIJJ4Zm2SEdWEPSmOAGyEIP74utT40f3L9iVEmOMyj2a2CArxCv
s0ixM1FlnOnfn3ooNTpmc+N2xu16SLHub75G/4aTivsFb+fdsvy9qvJqs+JX6XrE
PL02tR1b0VltPhqBYlfIHyeWu70CQrzp/8655qJw3oXySlx5aPXXA4zIvlL5oQMs
uSB+OFwvoyWvKCJuldXLkyrwAsPnt6JjWeCRPZ0T/LmQzenb8/XlyHdoCq4bJ0Ta
tRn5FAMnafFEofJpd2YSFjhj7DR393LM9D8pEbWSaBRKCpdfmvdFjwLyAbCSciqm
ieOLeh1Qn1W793ClXiXzzYs1n+jDSSarE+bKJasovtHlzlQsH4NJguxHAch4l+Pj
YJ93ELH+7Sk4b0MtknJoncwBjvcDDhLgPplRjV7MPUXsoluSN8WrJA6R0Yq3wErf
FZeLpXRimaMFnQtkCmg19f5Vw3VL+ngGja6K+RG0mGFD4Su8IkwywAgm1snQlMmV
MlMs1NE9jdDKRyNbw4zuV1AGtS92QNq007eAJUAYhm69wYjCvugIdwA7hTuRC7Oy
al+sqG1uaOGZWn4T7L22CbGBiEGnhKltcjPpdVCWlJuEunq64Znvsd4VFDcXWAAi
+Pqk7WNN9c42A52OXvZUiKn9bPFlw6mTS5dH2AYWd/ugtC8WVTmSVXK3HBgAlBaP
ohCo2/AVcquDOMXnpTHf3JGiYx+jMAPwad0mpdg1/SOUHGorIppJiO4nGWqybI4A
xeK8jKg1pEQ3P/ef6x6NVLzPPmTTUu8AC445sEhvUArkp33Kewcv0NCEd+oJs2Tk
hPvdyVmdogbbZWnMEa9gaJA/iYQooejyvlbf0Eg8/coRIaKPHwmU/T6SaKCh11Ge
TbQFniOH2alV8uHRg71/oRqqjwSYuglU8GCxkI/MZbRdjKFdOPTyHRdM31/fW1Ei
SdTEaRYZz0//xPa4xDP6dciYkpxETYZUR7sjefcTlJOOohkolO6Ph+NcwKLVUl3Z
AoVabJgmFTHFMz9zbHaeP+XmMa4tIgzHVnWmCStzfOFCYCrlohNznpKM8CMsojx+
fxKmn26ckbgOqH97CwOHTUcL8osJiukSubnGSpZvpRH9y7H2LKs4FwQJr7kZme9A
kq4pOUvyK61Wh51XlnpbY8bNmCcuEdIPM8tgXcN69lVDphm+4/ANKLPyMrRt9vkX
4lYODhwVaExT6wO95z7Nf3eCn8TT/KkTv66BFdAgua9XuJBoptmdISJgFqTMCAoa
ObrMCi3ZZ87IafdgycClWqLR26AOn7R6i0vDBn6kWpf+fFDkw3U9j5ik61xzxmDI
6etaoQije5JjRhP9PhXG6QGs4BNfKBXfFUAEdotn5QPfG0Z0vwtjiT6ghji/LkxM
PdS2069RBspNNIH1o7BpShZzyC8EJAL/hAWl5QotsqIDf9+E22DwZq7zlEXMtsF4
sq12fITxcKqozZC6a3zR9XC2AQ5b/+GEox0D/UnXFU3wctywoNM+S89JozEl2y0e
/nqjYod6p9vMEODby3Zk4slyYaqtUyLD/By2aOl6Izw=
`protect END_PROTECTED
