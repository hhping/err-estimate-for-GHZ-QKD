`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AoVhnvy8NYOxo00rJX6AWiuPP2vHMv5xouPMOrPnGMFVir0JnkaviCn2t3HquMjq
KvJ6qJmd1xhr+Q5ST2rTRQfU1AgEgY5LqXmF/thgbsm3znURbC19hLemSRTxo1In
xGHalSSBluVAlG9yVbXciilBR3e+TQrIrZDd6P11Ekt1hUw0g356pn1qLhfnhqtn
k/XvbFi30P4YD2wDMEVosxf28gQdu2npOSZiqzcnd9IxdxMSIbt+964sVt2LUaNO
5KuuAcikj6hlbDeSwDGEcQ0YCmayInAmejzJyac6GaVqv177d8+/oyrg0GK2HMzh
vtvihduyZo0gnWFwgHUA7nkzPTJBx4S2fygc+xgFPUVTehaH2TSQqev6omrEpOca
ZV/FBU6IOe6BXA1ri8E/otcbJm1NfD+EtCBT1TqPUidPUCXQOkuvGAh4Cp6pgNpi
jesN70K5y8jls/60wbuKC1Vc9xTOZkz2jUCI1iNfzuApSGvt4BQBi0BnikpXPkNw
6YYnUAmCx+nLj5FhuWRGnxYORmEQwEt0DqNrKuSrj/13XMw0wTgNqW9B2l9OpXbl
AAIxhQOJl+6yuUox/9nT5iH5tknWwwnPboAHDxD7pnvfGdwg/Ax395jpaAnjfyDN
i0zdh7on3PaCkRjor4rfxhLnO9MVpG9EmYdcgGqmR2KzZSIvCHsiTNHTbhonRera
auBQAP+QX0l6ueVzaW8V35H3O0NwsJXMMH4dVeI+vWCt0m2YehTC840qzFrUsTqD
GbN/MW/ZUXMZZNKivMlOglXbZE7PL6z6FQLMTQea3W62VIFirI45fPeChMnfFpAm
QhC9xa4c6+TPBjEJI9E2hXy1v9M9wsPC5+0OYXnEquFMK1Oxy7Xp433Ougomlxq5
yTQ6xigRkVTgpOmyWoxQha3FOSNRkepSsd6edw7sF2dexM6m3KvUGOjPKBxFV8gl
cqy2U/wcAMno62S6d8+j3wGPgakR92VHFLvdcC3Kkwdn/PnSqqNHd0xLCjdTJfD9
PC5XlO8MLq+vUZDKLzehsL6/PbKPFtaEDdDKFwTS8H9tAtNeDVum5w26z4RlnB5B
KumHBwfXSbjJJiDEq0xj3KAgo7Q33mFObFo7CiyKO4bLdgNbiJHYwMk11P4iuakZ
a6HBwQ046YkWLhP8xgc/RlpYs+di1IDc8pDFgz5AIldz3uA8cCL6GjI9aVETO8xQ
x2GFTizqh73S2Km1WTfRY2GJXPef4TMxHi2zLS5BfOOFWYmFX7uKqQbnknoNuVNf
cAFgNacA7ZLk7u9S44jb6b+TUKTsJ3BQV95t04nEf5k3BPuUHxCn0vwYd1u5FoHo
yVdajO1P01xSJ2ZyqgiWD4DFm/IGfeeqg67KIx1QcDCOYfIC8Bv6r8nCphzpUDkH
4Sd7EDd1hIBKjKnZUPu49Gasq0agPsJ2oXn5toTNX9FD/OIWlmMUsMeXLV4WP5nf
D/LH2FPfquEoCQJeAfIRVzVsxaquerQo6x4y7McNq0+n3EsyRlUMIb5n6sRn0EJ7
zyd11FQxU3R8YPFqviXAV44Akp6plpjia5ZYygnlLFOl5QMIzZgI8Z+kJnj9aj3j
NNN6ots5VdE4JTzpOiA20jfpV/vl6KsVbs7Wc+YVCIVBTZ4R9B/2APGngkPcJEIu
xO1pR1gnuFEW8TSLjCvP7IunOZ6Z4Vsi0ox63F52YcC8HEe8WzD8uNNjY/II7+0s
fCxTY9rJnMvsvGwIfVQAhGxD9B0tzTAgxuRmHscu/3SDtYFTA558kypgStUn5X9n
hydFJ1MNWyPtwg+DGNWTkfzkECu7aTM1+T+Kk5lWI3e9c3vy2h4ekczdCQwvbIMV
eSckNrCo02iz65JEhV9kmflQkwWTYXwlzSqF9YgYdyfhjLI+snaUh6hDiCvINJnv
cfVAt6HqXf5X5sjd5nRnlKRZdL1KxzaPK7UqRRt0LuSluYAfiL+3oib7M8jZ20UH
uT5QIOVwnl2HWU4WqDU24PyhV0UKp5k195AyxaGb6KO21LLNaO+Bu+HyA2P56FjL
mb35Ovr1VHDKfkZs0tGPpkiqpmG7nVkPDKlLkE9u0Ep0quTWpfoCpmNJJF0bleK+
hkG8f2BoECTYLfji1TEIqGyUFGiLsIK9nBN9b0xDUY9//lrl+/CXrQm4huGqV8Dc
/x2+/o/s6TeM78OvlFwsr1NbCnZjZ/7arfEQldez+W7cwcgKSUvL8uPgzI5yqUKz
4qwXhaLtKeCzDUqgIwaV3UuBmcPkEX0lIe+RxtQswPZaRCKOrZodmqSQbGgtGOoW
zDB/njisHjjAfARfSJuepqpZW9jxvYv4gBO23oOuz1HjpuNLYpXs0MhgHxm487Jj
p0P7obn+N3pMXe1MiKvXNIuNp+Q8+toSm5RUCHm9BM1mhdXZkXpBbgiiKUoD39T5
07ua2YOdlAaYujYBvHFoEzn/blPq5R9EBjeOZrWzjGGCEBuegcz8/H6MU9Oh95zr
jiZeqKG7Ss5344Hk0pAWz2msvgVrWbfQPIEYJUjiEEh0lch3Zd2D91FRyNyVVY9y
Pyr2A8tlV/aSz1GsN2TrKurBpuyG1v+O5YtlahDFZ/Lcu+6Do5b9b/LB8ai5Ettb
tiWIHHWoWKEzLIHO7H2ox+LV4QMOKtXTwdTuEyZCAyPtOSi1+W4Qx190MnPsCZPS
LSTKwhdjv+PHfwHqmjQ2sV3184xju3ba1ty0+G4Iwt4ZPkVg2AwHnev3Eh4+W6T+
2XB2a9lAAdhTyhk0ekXSC2HErg6IISp8z287pLDyIktuEw7N0HbnaSiRoYBQD/xo
rLiwJ9KMi43cDSEbBnB8sjWl220K0lpZP/7d0Ei9vKu2s8K9ZKle+dhjGplFLJoJ
mpQOPDRYSP106crhFTl9f+Ja1PJ7n9o1m8HDMyOu+c9AdbOoghp4/lTuDeW9YjE+
Kur3zck3ApVEphelqOR7pryYdAbyp8TruUlP4aepieEvcDjVuMrPf34opD86kURp
posgDMBMBxJjMbUqPBpvgap6/NXYIfNJP+jdJg732HwzIHGOCX2VnGYq+QNoH5nM
UueVeW2L4risS4LP3IprFzkt9m36swtmjcu+mbPfPjsuu7sUzUtatqbuLQ6OdkzC
I0XY+dJ3Ang53uWXzOqEwXPb4+zumkfn/JP1xWU0Pfb7nPMZB0rSBgc3rdTTmtTB
ntoyhwOVfX34HcWgwEId8mJoquxb17vXWyds8/N7EukWCcn4bCMvzAxa2h+a6LfO
hA+Cfhol7YYEudYMJ4LswhOIkCH3eyxZSn5S2VAKzLxijYmL1G8VfUlJjuf3JOob
3FYQU/vDwq9BZME5I6BBIZZmrmkDeUzG7q4HvcQ9H4t/iIXEiL67/Qqq0KwSfDdc
pYyypNh9kA2atXvT+V9sWbfrT3wN5N9NxP7pcU9MSfGHaV2yZPtnnT2L8GEGTrcT
Gp9rJOE13TnKXukIgG9BNvwKhobnrP/jWUyNx0VJKAKhRAhmSwqJE8B/1noZult5
fbgNP1taTn5NQ5dm4enLa5UfntI8WA3ki+9qTa0+PEPxqnvOQxeYCfvS4q/ZsX5m
bBLfbg7JwgsoOFJNi6XMI8okP3GqeNzyLqj7owaq1ieQ7CuKirm2U3Mq/h24DxV3
qu+a7g8evGTSq7hTA9dfvtnOIZjmeFJAzxI2Wd2k29Jqfzc6K3Wampz+OcfG0P94
lAv6uicc4D1pwEoFDU92a3Xi24plDNRNNjI/rp9hAhGHDvu/w3i9/5mqFo/pn9Td
VjwBwj19F8+Kg6G1MtmyfhPp4V1nisergOzhyGFUCGpIuBEfaJ1rVzatPilZ09/1
+ZoRl5KWFThpjFitJDIqjnUkaCWihfb0bYY5TxYgdQ0zMruk7Z7XMBCN2Ik/nA/t
Wyz7hPMvPxLc9COuKDZvWgWSVFSsGX4M51Nh2NMcBHbbUsNc9usj6zV60AB6Xilr
ITUHWDHtb2DSNNCGs+ftsQPDJf0GgA9OU8hn9dD0u1/ToY1nT6+psnTOCDMXQGsQ
db4vVbVsyJ8zNFsuQLbM+1/hPQJRY33B4dxGwVmlhlaiD4QnXXXCLNDzF9F9U8gW
LmZIO61dZC0+Sl+bAOO088izHeE/UU79/whS/vzeLycVlPOOPA7ptUWlLLeBxHev
8aR8F8KSkwxW9qQlRZU4PpEnkI/U/V5i9R7WeSL5mFpMuP1i7Nmu9w0Q4Y4PwuKf
V6CEC+7MmFPnQrjJ/8KhiSxoUCfw0ewJrswNSUuvUi01gmWVAQ/o2Q56bk+38bXk
JbqeRXmDMnm0QBGyAD4XzJeeXHQ75RTCL9PEsFU2Gm3tffJt9E0QItO9WDntZ41r
XiAmzgemEv79/URLEsibBikWZ5iqDb2q38H3IEoDtXFoXFHItThwbFrQGq18haSA
KbjXHMjJ9umwr3BdApgRYY1jPrpAjftj4wAf4aeH5EoEF4LErMinFd6w7VUMmMWW
Iea9LI1QcYBlRMCHHa7Z1P+eqd+NFk/qGbj+gbfirFPDL6gSTRnTCEoPnfQ5RSA+
Nms5eBr9MKfhOGeyq8p8XkRP0IWCN6y5n/fnU5TGgN5d2qrPVY23rTF1GGC+tb5F
kom6JVjPHdesIP5Yce1SiZWv/yqXXJRbFY7PMkm3mt3TlejlYF/0tUlI+YAaGOgu
QN6ghFuoa9qJLrkO+SkxKhnXXX8WCUA6HTHtpEqqssOtj7BcJW3AEmJkEiHJBu8d
A06EzWMcrZLq+XoGYvfFaUL+NWZkoSZI/0v7Z/+dZArsC4cW03dN1ORDVVu0vbf2
0AljSzmREgTP8szHouNpkid13YQwKgnAs2DU1qiWV11Z8nApbhlK71e2+iSiq+5i
nDe1RoviggAXWq68ta8TZ4JpRFzpW3ziO0XFhIkg4mZe6pMnqL4sdxvskkvn5Piy
5ZYWfSkEyI7KGZJjlIWuTOJioYFwS1OkZhWa5fTy0BNxayaStbCRr0kZtqu+vl1d
gaz4Lilstlj0pdK6xw6Q/3bmDdKBSEy4bWXcRXXZa1cnDVcbVsC5r5VEVzeowZSp
sPnrS7AVAm7izf5xv8N1Wa6DDeCHTyBjxR0aZCawYqWE7ANY0ndtRltXsYFq8m2m
jCvwOxbeEOCg2kSehxCA2cUeMBS1ukL83nhUU58lc4ZOxNo16k9U7tVeXORQnKhe
AX1Xxb+89Wmp+PEeV+As6f4sLOSDSj1xI3UnRWjJ/SGFX6GKRTEOm4RoPep/Z64Q
ks9L6SocccS6D5fn11N4dLLSTFLs6Y+wCr9rXDnB11YQYwrZobvukykJteNc/jBK
FPLFlw6g0O1hTMnLYd41bnyHVayBXOudduGvmLM6qkCL3a91P3Lmp8sRdc16KAkW
3HvK58ZXsuNtWrEdQnPQj1sJi6ADyLtVUa2H0l0MAM26f8mWgWryhBeFqiNS2Hkq
bYDFiReR8reJbCmhpZdIRCXqKnPHNacq7rJ4zOfn8F9Cr19jBZtacI6uf0AovcPO
AEkWAI/RYR02fIb/OejFDp/a6GT+ku+l5iwarbDaITge8mG3/cmeMOe6o/kHT+mD
lCeaVC/hBneVkmL+sc08BUEPsACL9tn5/6GutbVEp1huL9BrY2UADCnYvEWxYO/T
EgjxzppAv9xMS/6HI+lRnmyyds9ZUCnPN0sLr75RSW3OfIbHqj8Fdr0dBjtnKJww
3t2PxKucBk/A4WxtLvIsYZvMswQ6ygVhob2Jg1JANDJGOjrOqCkYiAgIKwR241ZI
ZDN6uSQI5YYkNAT3N8NGm3kRRdAwS7zXxQbWy7mmDuFHTB1Mzb0ax5JR+EKaYWuk
6QI5j1BD4mFdTe+jQPgsMb5iP6Lvv1hJTWB1ct/tvkKKaJW7OeFhlttQcrjSfIjI
HQLAiE+GCW/q8uxSd7yfZAs3IuixRc8/3xtqAm7dEVqUhHakDNweJFMhvJbR9FXr
KJC832PH1t0LI2Mvk4zf4jU8O0H1mguWBwKt6oJNJmUlasPQU0rFgOJ6274cH/Ai
sMiGp/ioMd6XoRISe/BzOWt4vf6efcRcmp+fbq54zEq030Sm4KNYldu51RfcC1cL
sTIDuEgCCVDCc/LA2OoXS+0rCj/bufgclIokYm+LzDpO3CwJTWBygfwWnO0B5rn6
h/iadmlqco9jps8U4z9sxWLGlYK1QpafzklQNBQ9W86gwPvFOckI5KMiv52tu+9O
ng/MTHGjPhcTZqIqGSyyTk0rqmWvm6Efh2xnJqbzoPdvf36GqGqgrSD/AHXuIB8T
LqruqW2KRz/fBdXH/G+byvV89OYYPkZHB1vEyo3aDdMF2UsuMebQC53UKVGftBK3
btAHFWG0YhG5duun4Fu7RfJ8tomPI86/xVQxbxY7IBI4IEMRiwU0I5GwFupE7yGM
2SWlVh1i67nVRaKWtS7wF9DvpjAANjdPEg3QdY4R5c7xVvXtu7RskPNoMjVMgfGe
rVjWxPrAsPtDFH7AHB/BoOZnhRIE+SiV0cyAiokapGAISZ0FqFslgp5HNENSIUHH
oTdJKs4v1OxbKgbASM8JA3kCJlHlvQQ73lobMh/sVC7kSHfRTlls9hB+RKR+t9P5
koPXi3s/EyPLKkwjX4jnYBWKH5u8lzkeeyrFCyF7FekuyxVwX0sHSayY4pfLXbdT
hU8mDUw5YHQ2vxCaXHAgFCarHgycuhK6j06OueVEMIfI1a77rXBfu7FWqr0GkFxu
aHTlp4sWWzT8GqhryAySJmXMQTUZogywdGAs4Ptb5uKK07LbVAl3qHb1TjHurA/t
UV8U38zfXckP7PUZMEUOO3bo7amnNGWLib7Qrj+A3+DaoeM0/f/ZouylyfD9FsQe
rKncYUL5kYlA+jPSIF/RKI1EDZPE/r5l2eNNWfqsFFDDL08qqxUxhQYnwJjBYWTR
oq3FNc39x4RtRoda8t5X8ySiUV+7UOtt4c6emoaHMZPL0Y/ufm0M1OgJ6BYmhWV6
vnqEuULJA1ROt8IoKTfeoIKkCxEQ63ZyEs1HVngkW7TM8H2EoErH/LAuFZzumN00
g88ws7kz1yyqHzhv1V3SKQ3zR5gry8hkk94vSbuuj9tVT6fL+By53sKf645rhB5/
VW0Yjq2Xdxdl0Dv9TqO83gM9Gtfo3WTXpJ+b2so1AHUxTySnw3jF88m7XEIXd5NB
Acoy5BvyFmfllP04i9qKwYbvj58q/ClS4DgcMJjhVMNPIfsssHxUZLrAMRiVmZnj
qrRxO+LGJh5+HRdyQvs6ZtsPbIydrKWo0IKoHxs++SBpEetfbtRRcoMZbx/0czi+
HtZNB+hPln4LCqZYWDNicwFgSzuiVXHHvmigBwfGF7ozPNT15C2dS3lzh14LqVWm
8UOqwUef2JT5cCnJ8m1dZ1+GEN5k3iugKFwt2GE5bU0LHnwAiUSLQDtfT2WBM02Z
2LU5syXgKBeXL5SXYP9umwMg5DFM0c91FHDoFgtx9PG0SzkkE5B2ID281dEPyjyl
vSwYFUGIZR+3qpucnhazFH+idYJYp5E9Ffnh4SrIEj/9Csg4S5jWUgSNTSW7bUiT
V7N9Imn1uQ6QkhF9Kp19XW5jb70nLsZiDTLxwHwUy8Zzv5ZHtRtNVg7td8jRDrnI
fCc9ZRp5SZG827D/+JB3JeTSqIh2umY7aZQKS08FCu7ZfwCHVNWisILSiU6PF9pR
ma0bu19nGWK8Aq4KruhZUHiK/qTP6joogOhATtbukZxYHM8OZUHSmdCMSrQ+ogP7
hX6VwDyheSnag2JOSTVFJ3QJwq3y3wSCA0EB6Aos7CvHyiRP1rHyLGNWg5dv65wH
EYRleYlIYf1E/Tira+3dbxe+9txJ+d6weuLIw4K3SKKvyVzeRIrrjWlKqt1G3jSq
f1imeIMO6IkMmpsNP7Z891swi64FJ56I9w3l6u/6jz2yu5mGMkm3XX9HlYnPOAYH
DK3Ph5LSdJcYx035KGUycrJ5SUEfJ/Jk4KpBWhtR8s03yE1ehURC2wI/TZUt15CD
tBlEx/BCK7hUgJ2eU3nnTXpohr7VUr+zwvBzX2Mm2Z+/Qr0i24zZYXlCByFHNzHf
4/gzwxjEBDM0624APHBlhE2LQzew1KbbseubI3HYjmPsw3jFcbbHINHz2E1QNK8q
queNoDEx4V3ombfQ307H74TFA/YQHlW7+yVrHaQTnaf4t6m1wVuVNhYOqRIfN98L
hJDAZGF9BfMWESQTGSk2MGlQvqOzywCSz+gnGQfdE4l3MyVjyOb1QUrv69DNt6Cc
ZYpQ1Yog4yV89CElfb7a1SOzlTqJZBNrrftEtfEUfpm7qkQLHunQpdq6CPOvVhKz
1EK0pAnrrrUNTyAUDbyyoxV27AefxZvh/gk+mcSF96bhxjdE8MlbYfNugLbIW2A1
ELEmISTdzfFbKjABr+VNx4zINpoM3+TM9csoASXbVd2AtoCMeRaU3OsLx25sEl/I
JznbsW4ABXaaFA0GQYgdWdTTKXp3nhOuWFy+W+/N8ncsNUgLKTgJELpxQ9BFicI8
Se17oLyIf6M0XaOoMvPWdme0OW9gRRMI2PldAFXVibqFMza5IJRYv7HpSA0WYNo6
APfbjy5z+qf527CJiel0GC/0617FABzzpGc8RWEXOdDosbcwcJ3wLXh8J9/HXuzu
K+GFNklANWihgQeLAB0mxtCowCqqx3fKCKFkKHMbTg9K0S2q2AIBIqVvl8PxPX+Y
3qosuOtsd9ZeVGxDEDlr5uHfoKliHvg9JmUKDPLwyDa5bplTqQn3wMqpmy7rGciz
GhNucRVJDLx/F7dBimSj/xfHd5b67Hd6IBJC4HYY7FZI/Jqw1InstGLyOqFFxauR
4+YE1c56jLt5eXK/V8fksOnzAS5SBsvWNrZiqe05Hg/kyiZoKsCwN/ZHfoEU51QN
yzNFICp0XvTiJRvfUBLtl8QflOGfYzf98hWZWDLznJKcKVlRrrIwI11ApgJaHz24
42VQEGQqf5Fz7+/Co2K0OGAjN4NUVnHnNIjtfcFGSy5KHeQx/IT81GwWbQ6Wgdpx
l3OU7BSwachB7SOqR+u1vVoE71OAn+tHzZQFk3x00LWV+CWOgZnlgWt70dAw0lZA
a2ST6S/FycaiNpJjwB32MKSp2WcXxORpvusJxBB3m4kyoHPwdMkaPCoRRadaWMLB
lrRNSy4Wt563qoMLsZpHBJcGxA4DGgG8m1AeyiHo8d+hfw9oC5XnYpKBNzbRyU2j
kHQNVdlx5WRyP8yqoC5/X0F4ZH5/TBR4/j5XlFFO06SpAhTyalZjEbIw7Hh5fRrf
3WgkXhp3fEWt7GxMvW9WZKIbaGL7WS70bImbgRQdlsyvfEfbI4RLUc4aqI4Zqjs2
RQLOyi9GrUYmVq5ZX9O40I9pQQq21o3dUI8wfuxtUrNHLKTK6Q2lyM29x+7Jnmyk
/KltOwGPSS3bLObM9si7Ft364iZfjNqO/5nmEZRgO6j0MlmFVFfzSIv5jTxPNu+O
zkqu9iCZm1yqRrtdRC6/JoOA7rHm9E2hA8y4xvBoD5fAFs5mXYH3jnUk4+AF5Hat
rwV+cw8YvS+oajpyhEW2p9WNn2HjdFvezR1axSurrsURlXr9hY3SmPpaVr6u18zY
uP2Yz8pzwIS5lFt0WnmxUAtH3rxhDr3TOs+WvMBCjhcw6GZk5/Jm+GusbhI1vEJf
tewWXkBp40Nn36eyqodnteCD+NH0ocJqtea5VqxgraNbZbzc40nW7ZI7LnG+sB/w
OqsmOOlR0P3RzICx8z5/FnjmQ1z2jZ56r9PyKDmluz1R+mxGsCCPj6sNNkQDSo44
UGLvU75M+JKtxCGgpXupvbZVOk3Wn5UWSdX7odwnvjQ7jDeRY3y1ssQyjTBEh52+
BW7PSYFBO0UICwUvRrJP4wDL6aAaEUxkzHIv028lwy71yQqGEcIMsDi8pz8P6I72
Vg3el/BybkuX+3C8+6ktquf5t9bxnf/LgzNcsMK5h4kAOcaHE+b8YaUicdMsWUPw
QvDcUYnmKswTXNXs4lEPdim0SrWMRxa5Y9nhOuPfIgiA+dZDOHuA58DBptxjgekC
kK3UoETATbYHUe+6oJM8SBYXdp+47xsO+wphjbSdsQhUJX4oKBHy8X7ISw3Nj+8N
bu7aqyW7+Te/oYLkQt+7wbGrNG1P9DnQ4XYDf75P++20sNMRDdqQBQxqgQWq6yll
2aL8P1S7gg773vwubkfzf+azCjpZTfSkC8z0haDWJ34SigWBF8jSlwXGbU7fv8Yj
Md/f/CPyzly6EYhJOYFC7ieOg9huPnx0t8cgmdc1LW2VKhy+3lkd2d2Px3B5fWDQ
+xGBbtZ25HjG9D6Ua1zRZV4VuzVztGdFsoevaNjbDwUUR7nWTQfPg2IreW6zFpq0
UkQ185YSEK99BhVCW49cfJVx16HfwaE7Lz6kSZFWlG4tAziHdalBNZg5VXisfSdb
KW3Rm7yyG+aJTZaeElYijO6BQgu9hoCQjlI8JW/0eh5URRUt8SS/+z0Ib4c0k16z
ht5NQ/xeHuLC9A9nMbKJM+6gYP7vu0FmY89KNW/jFxXk4dgkxHLhV+BRABLyO2uC
O9yywbe9/UAse3NWfIXcCxbY2Qr+yvLc35stgXD4bCrCC7yI7Vl8+EpSx8aakJ5A
UGBpAxldY1yuiaa4OuHqQbGL+mDJGx2ObrsMIVFAlSKZS9zHA/pcpuIrg0Eor/1p
kTxVLU5yjXrqe/OcoE5CH55uYKQMHR2bOn+yP4K27473j+6wrEhcdjFCJXiHksh0
IWCj9lysSj9+6aCVVOw8xpeJmW6NIZtpyRyzI1IA3Ar5bJ3kOumyfhgqnr+F77WO
c3MjIbPqopAmhsJ7liP/NXshwrZxlp5f+IUnYIiTKTrCx/W/JOMYwzRlglgrpL37
X7/RZl5wuZtLBVGGju+1NWYzEeaxLqZku4vvjNNH+6Wb0Vrij5uZpwX+XeGdjHQU
zezK7gkrrmsou39cuKTKjuen8ryUUD7j19NWpl/48yfA8rPwsAY7rd/TriSaKeuW
3mOCJqA2Z2HFL6+c7HIzm9v1L+9q4MSeW4xYeneKJxhPY5OWFK27wJigtRDhVst6
XOrX0pKARjupKHbfKFUIdJ9CxNHjeCiosmhAFyDsZkmNdgWQN/LzTrpTlERjvCdv
mxPLImN5mcRXpxNFIWJKnh65ZqxyFGA+Qo8/4SW1mh1TBufpXIybIM7lGa2bOPXi
JpVw+toiMSSIF43MDvwmVK5ae2R5bLA9TotFxEEL3nmAtTrOtGNWBY2+/Hp6CLh+
yyOeFC2jNg146MRk0i9MsqTei7UunGJvjscO1JBiAvbPZKV8jWop7GvWfDyOG/2w
Ji/HRUgvtoz33+lVstr/OIUmYBj6L+kMn4Hu46ICq2iAVmPbIZ5RmaZRCDGDQlSf
YWzcH9DQHvP2032jAERwPFLfJiwQj9YiVObYqvwg3Du44ZVKC7TX6eGEfFxd8XlT
vjOJYeBSlOyioYs/ILT9S/vv4tvWt0lopQUWFE7rASZjDoTHGxtFyEdnLlxcKDzG
19AG1oce/rv8Q/RXfDbtEaqtexid61wn8FuJhuSmlNuTdDJ4unYZTaKiV91oJ9kS
VOdzWn0wQpCRSARn+1BYCEByoF8TXxCCzrj2CtFa8Pph8186Z8Ndq/mObjFx7nKc
+GD9gdP1EofpD7ZZsimZbbfqmiu7hie6sbogzDBrl3oeRDesBDrs4MHnq2UqaCCa
EBNr464R706+cakosBwig735s17IPRUJZhyKyFkLeAvfMN6StsmIJgsUW0ZGSYaZ
t6ORV4jqNrhS/mNpp2awFvEj2Sn9DBUhUd6fBmIbI0rLT/NNt6ug/9C+LxVJOiRz
kUY5c1i59JpVoFfoa+MTVG6gZLOn3DNVc2Cxt+m33TkZx6+RfLDNFS+mqf1jmc3y
OfT+5rXGISBsR2d35pVU1nzliMPgs7ETlz+108B49TSu+VkW2mgXD1KQmEVLLExH
bAWQhhmSeZQMebN2TM4L3eiHliGn+lNJhjNM8x4NmzZ9vgF8uYWKly6O0ypKcb0o
/RFp0DYJAx0uKyKgn4wMIUR25gW02zX/Im7tIfnigMAW8M9U8QBiMWQz9ogDjcWW
Psde9MlADbALqdOfXBgWrS/GDkn76r2o7ktulULXpQmMiuSaFjZIr2oeaz9d7vil
ZtCUv1n0pskQgjTguzUTTN3+uUte7gMFhZfD6BTp9VRPJSELnEzX/1hRM9Rfy+6U
MFuwwJir9xS7tUr5CrcB/j9osMRN3PKJn/YyQ7tFpjuhWuDrwcpBFU6itL5QDdVI
swz7xc+Op08K2cAwXSwtZOyzY7aoX3PTwr57HguKZST3dF7oAw7MlH+RSl7kSU6K
eDKwpHJhkstwCmpntZNDoUvmREKIX0BIbPjq2xiPVRDMrVFBzOqiMZD88tQXO3GP
RZ/ByxICBTi+X+2SHLrUWk+9KF9RxmbMV1zuJe6kAKM4Wb03elR58mDWqtoQm9o1
7TtZ5B6h976q3Obhy2s9WepUS2LrKTBQkWmYaevoh9RZlrwkMTwIrmAVqonIVGmC
N8gXN2HB43NQQ3RpFrkC2pnJvjUAL6V8zNUwQNlQQyF1ttpQuSAaJHCCWoAsqtuv
40/cGNuuW0L9FU6tpkSbQTKHM9Uhdm74DFHvzsghxJQdxRYDPuIBK45PYgJpnZ7A
cg+ZeVvo6GyRmKUSE0iBtAzHLV5LmVm4Ey9BdLNiEcNsuhh7O8oiN9SL4NqTYLyZ
3NzbfRC3X2PFU94JudceU8V+DRwcd/7Sy41ZcZdVs7mXaNS2fLyPHSG8E8hwagRz
4bqAHyKMUbhTNbKCmA/pmQorxe+FmDBLiR4h+2WonHD/NmiRrJh6Z7XNiap7GQ3V
UdzE8aGkz2qwGyd0V7nmRrdKvP+4NsaeLCHODg+OTBRKM0mK0gpVLPJj3BIuT3fe
wAlhD+cp8YerWSianN5cm3U+J1bz6d7+MnMbX+Zng3awz5o1cxxonbFZi2VZopSO
c/h6C/NdGTkfKoN7ZfvUjJpFFwcJa59ds6wecxSn6bNyzXa8qoTa9VY0TNkOLauF
o/aDkxkAcqhY5X4h3CzQdlf9ofV8ZUET2qtZGVMBGtL2s8NX2ZvrQTETOn+xJmsP
Zs52GC8FEA6Hf9A8b2Qz8i1G5hfjMeB9IcY/SNJ+lfl39z9ZVLC9Vi19d3fKfLe8
0EsmbEXBAlrZfxlmpFackj4GzxHbrQHOT8gyqfM/QUltqTbFJh23kBy4llqDxjjU
FO61p2DsNsgU0GUVcvIOIqdf8eHLtQD/H8Jl5HR+2HJLAirIQXvf2zk2eHARZQqJ
s9anEiEoDj3ajJFSagEYtKUMaVMuxa5IrK5Jf0OUzuAQFnIVcA0E5wg4vSt9UoVU
LcJxlzvTlJkaQzQ5z3GvtkvNTah5nkjssMBUSnBv/+4s6g0SqDA1zsQjbcM2WKRJ
5XW88ZcVLD+QOq69ezES+snWi4EB28Nm+U+j5Iy0xSIn/G/2dZbmNSOagt/yWYv9
pbIuOmtqk+akIV6vzFl95VYAcJBvWuB0Lken2mtKaTPLOLN1enxIYvpuKFZNI835
qL/9pHjiJz0PCgZj2nrSFIryqGbCOJpDT+l15bgNtL5zSlKU2uu+4RjROwt/HZEG
G6X3KQxOT8LTX72RKh4oc2u6uk3pbgImjdV7WaQk6w/+FK4md0Zrfq1zMcWAGa9O
M5THTNl0snx2fi5OpLkUgimQGmdDgScStIdjODVrwH71GNdPPqkmo0Tq9NFSaKFF
WpR0C1WbQVQXRJZNViEuPZQ2T1z0TEUpSYW2AjxMyQJbEqOD2QDWXg+oukdJUxWU
oBbOCL/lN883QhrEMwCQGMUqmhQVrdrCI37nNju/XOV3dAJVMqPqYg4CzPxgOB5Z
UKH0H5G8f/mCOGG9d04JOvLWjUImYKCZJybyNBCgGfWWC/SVcNYU/AC0n+uGL920
dfVWFUBDpqO5Zkevf5QBPgY+7TgbgrEt8aikIx9Lz3J1BziswvWuMJhAhZWzY1CB
qI4u3yAZdhalTSwq17t+IvUVnUHWuPBBWdiHt9DjVvN3nsgvzWe+zDd+ptRuYY1J
a9MMtc8sqb12RDy214QRcbabGDyna/+g8/KoVNGx0zFkiLnokCk41g5xwPs63z3e
FOkfythnHWPc2jL9RCkQbHrNQ1fL3Ut087zcakEj4eqOvZeiZ2jxrjQxqpq6AMsC
BvHaPnMTZcLbVa3dACiKA5Len3FivQMpfHHWLBRSgO//+3yZnyGoxJ3pvf1MVtt+
nB6/BSh/yprjP+F+WWH8TM/HsGOxqDSEQy+VB7Mx1UA6E7nS+BG7DmWMIVLWVtpy
NU3LKskuQPCZvnUhk5jj7CoLUKmP20szXikmWOYDJx8iwtAptC/rTHsRflkpIMpF
jyFT3indqZ+B3UdmtAh8HRlwpsWGxSlWO/H8RghQZH7sJx2mW0augn7DE90VH2qF
lLud9rbBuf+gWYpdyryD80Co9jpQmu6BKnxqhbkpfk0fjzeXIGRMhBdn0mHMQmlQ
M5MuhUPivxzrRsCoLXkinEt6mtjlLXY+kQoQJIw7zmaN9njBeL+K26lUgTWZ3S77
RNKo31weLn+thSO7Jg3ouP1Rpu4rtvO8eVDygaJPPiQAxQt7ANMnBwvEEzn/g8/h
GZ5eE+DTT0Eup6w3tIxpyc7RZ0f1+974ifCUPLsp6nTJIbXNF7AMxTu01u9cnD8r
H/7PFC2iEya7n03pkBgmi7vbqw56gCeA+v/pKLPYCWdQVJvLx6jQ2BN5xhhwbOip
uFsbq1Nzn4wtISYFQGAtAV2bSgxcSQlS0LzDpMYFsgInSJ8LZR1SMXBgGSHTvhHu
sOu36y3+V+9g4U8btveoR83VpCaoCTfDE71oQCoYeYwZQFuLUjdBgjHLRm4dmKD+
zc0sRT2ava0e2KLJ1iakphpIU84ApGWEhYH0ddClrMJfRY29NFBzRvxk8vXVI/Ee
2xUvdgXQkY5sxNnoKA4FVLTnv6vNHvrI0SWVTlmIurOLaLQTEanXCkf8Ijt3cCgr
ZlR8XpB8nHoUS37Qy/aJ11uDRvuauRnMBAC8WbMu6J78XTHLvjsJEqgfMN8v0mBN
cgHHapgo3FVMC4sUD3eQpWMnfd9aeyaW9Km9jqtXWqSVirwbiYq67Odr3ES1oCN8
4USfaGT2eHs4VVZQhDI6MfyOeixmUBRkCWOku37F+N15Gh2G5N+ao1v1PoTbxl/D
t/EpC1ElSoHWWhG0Di55+nuFa7FGhAMePjufeSATX2aV3A80KMbb/dZBpFLWQWYR
nxTzbF84U/oPB+ziNubmrKpqqccQv8BoM3Gf5ru9HJxPDOaM2SrLHx0DI/+1wVmN
45t7M8TfJPISezl00mRGfzS/Ayzi3JS7NAQLesKoo4iF0CNAw229nG3Daf7JmGWR
l4qAS5kG1A5PLm/90rrF+Cc9rXzo6pYKdcmDwew7S8CibqP/HHnG72bRl0uUGStk
n3bqPavzqCDzcWCF7cmXhMc7VI0cwzUz34h9Fsiws2TNPtja14PGlAlupbTPUgvs
UUOfRIDpTz9Yjnfvn7g5x3n+CpHZ88qy2VhEVGhe/U2vxFJ007oEJ5Ah7eD+uM4E
clatNmf77vB/Ug9w3YjLKeC6csL9A4H3WMYWdV8a6yl2Uodb0D/ymk0VuqUPxrX9
yJYDvhqvLV4f6hjdivGcuSSZxOtQNx1TNvJVETK7/iJP2Afpdr+kK94AyYd+OgJQ
jYA9YDXUXLftvjrxhxERcnCXgJ9MgPEfZO1aWdGOryZMBBJzzXoUunpvMjsBdXo2
H2GmjiAfgW0Ddzdy5Zz6HZAvJ1JewF3Vsz9vEXtxkgYElieHP/upkarmoBARz4bU
vjGhntKqqn2WKOz6cRqqCuVMDo+p0+lyzg4fGri4aP/S6InXrAYH98RnmcpYfKKA
0nh3cOeUIpgKoLebuXCuWVZjSJEUgojGfHdcduQ2kiD0y5heJyckL2j217ZuxGgH
zNwmOUK+umNvcHCwIUokO0ZX4xHLzZH419SAle1QpUCCvVDq6gN3RaRRZrdn5v0C
Wq2rEjdBkT2Ybh5vvRYHT8RSiBf3chzH3P0wwnTwl4y3QzJOD4H4h0QktrwlUTwk
TP5QtuE67IdEHBNBSHMS/IvcBdkmFSmk8G4bPY3EOBuGKKl7/A06B1yOjEDjbTSq
wJHWsYVYWgplkykvwHr8W/xdF8DRrTo8zhfGNit+kcSwPhg+VsYa5cXOdybo+H07
3yA5yVYxv273x5tyqtK2uyTYU9qbGj36+dlpEmibwKpM5POUjsjDkdP/bdVKV6ne
N8De4eAjUeR9I/S5ZCLC4UbleAkeTkP0kfcqHYUrabjWV+5SgY9MOhSdiGjX7/S0
vg/qMCSkQ8bK5MnC1aXRtOh8uKYl0Cb05lZ0OBG4lrMbqpGso8V0ZuJDZ8XGXq0/
nKiSIaxQspNKbJ5HTKv6XSOthXdCP8rPS+OvtjKviAsBO56QKA/GKaEfiTekDR4c
8REnvh4AO/i504s8F5buUZUQzwwQokbx7vSUTQpjqOWQ9YpHTDogqhBmC0PMBAH+
BBIX5tw23hy3hTMmQ3rJAzoGNiqatbUWRpT0Eu6rSr/yn2PA+G1EucE3IOhyj38N
UnBceFoCBipeqef0XA5x22iUpikfMFU9NTlI4C+YAQqc+BG9phxvxcibIvISXn87
pIAxFXIFUFIRJRV7dgtYNXqR5AnBYoib76+kgKJ/BDxKN9I3AEmZIzLzAuH5CLPs
Yo+0GtQWbCjbNzbshHF7rinA7gDMyA6DYAP/rCR0GbT8XeTDSASg9qgLu/0Lkr74
bWYYAbdedx2J/0ELlRyG2acvJSC8KXmwsZa3Sgx5XCkpMBDNg4AAIyARG/tEEq56
75f+ggYWDD3EWsmUXb7R4+AK/8E+XwRf10s4z0w1Pdlhu1eA6/M93AsD57wuvDnO
Bon+VuHl6Ribvdd+mMlJH2W5VzrRj9mPDSTQHP8zdF5f2amBuH58oTlvqIVV1+q4
rigjvnNWR4Ybg+6uL7iqAh4Bl/TFqeJoCRYw/V5ojmljUYci35srlqs5nyo5jZWs
21HTj0xOeL3TStuJYhgRXctslNq8jrGtmhWfpzkZNy9MiTXHg91wyzL/0ph8TjtQ
pmvyjuZXXDZhIjf7l+V3bxmOT45jcSy9A3js/Ok72zlCC3GOb+AoeCZyfuY5QPcC
LbIcdVdnLLMT0PtOngfAXv08m1ZcAnYWrt+JFZqG/v3HW0pMRbvzNSY155UbE7i/
luZ9edO5C20wsXjRzxcCJfqc0++JHtlkGU3EdDyxtIb9LfOSHNTY3/R2ooiPsaNI
uOrh2NPHmwo7gco/qNoUELzjDtQWP6KwVb5RfZKnXGpdDYJttoz0T4Gwt6TAQU1T
I01rPwd4P41KpRQuK7NyQdg4hn8NBqXIJtxLWfY/s2xDj5SPRYnuW55uQ5GjyHkW
30Je+So0LmoPtpyu3fhlYnp/mrdKk2VXd4wc5hz46TRjt/M7mVnCLFtbexJTtJNX
7Bumyw8Ng+mD5Kkg6Ym2jWx23APn+2r1uCkCIcYVIH1grQoHFWou+xOBFjWOHEAj
jXTs26aiWtYiuD09cJNEpryGesuaD02urjuXKfH3A187usWNWFm7+Sz/nFsgcN22
pYgr9brbEYHHcfbza9G39tFEl6+CLtomv0GdMJ/DWaNJ05ZXDzcpbA73UGUY/j36
xrahcH6Qhl+O3MIfq636epCodhKFlFMKlJQAi6hs0g8fdddixfbcu7ydMENzbWWr
dbYYVrB8HuVnYcUoQZRxK0xCZ50CQIMnvld6ZDSlw5dFDOd0ma4RuaPY036LK7Ym
9zFIS8KJsDvrci7xRZdX4VggC6+xoVsfedeG0OxP3Dz9GUQuhqOazqNO+KjV1rG/
xFRRG1NNwX3NeB4SXVqNvrNKludIWTQhHRPUmbFwxbMkW33XHa7rKCHwsev7UTFe
JWjwLGGvOm6UDzxRZgtLtnPLT/z0PWOwz+pfM00iMV/PqmonuL0wOGSKxLbns7O2
4dpJzpIJJbC8Ip1iSeNkHC2wJFAyMh+lTWmOY5iAfgPeTeWh0wuR02nslrCkdQbe
1WlWnLYrPgXvqxD9KWykwJtOE5XjvD7zV5GqON2Pz+oIYepmf0ZktHTfXJITnFN+
OAlSSSQwRFEjLq8Bn9uDH5/FeRZjLiKo2LTP8lR3JyyYgSK1qOw/tOBLPEkTbK15
q71sW6DQDOZFGO5TX1iJUQVA4O40Wbi4YbfuWSm5JEb398AjHE+D+f7hAr2YNAaV
82/wcfJit8fSER55JX7Ie1fnFqxnpM9sj+G1+ORoz6cpHWhvQ11P8Bka7UNXP5FU
2E3tqFwg9RPfOHOW+XTBNguo3fpiJOR/6k/j0t1NNYd64WQ/m1CKI7hs3vNaH1dV
XHL0VgiH/vYuB2rzd7EzygMY2BSExgCYaBKcq0oIFuvJESixTLdyT6nWHlIZRLG1
Se4Cyyrv0uZ+GgePCLhvNzrMphVMXCYDpVHFd71M1DlVEPzqRGJohx8YJwgK6v45
uhBNzQSOdnUXtOTffnBomhKAJDD2IYOclwEOeFvYh8TIVm9QYa9ucZP4x7qHGhKe
C/nweFSVI+R1wg49FcMktTmJ+6VfgdKHhC4T2fEVHDpxSoaXcfJ35TPFXAVtq2WV
+M8bdll8i1KqIg7Fb4XB5N1jK7sM2o3QGSW2VsB3YLL/zQxAVQu1pFyvn0mQXNKs
2sPiwXNTSss5jvwcaGJkPs5JhqHcZi2iHIsnX40KxQRLU8qP0SAxG/yLDS18Z9Ad
3YVcYzW/n1541uzmjzg8VrWrx+9AI3Mmv0qZBReXT919w9nOSJeOYlLXhDfVhgcq
L8BIFJpYtXBM8hknXbcqeM+YZ9NGpnCjd0OxiRGHBkbhkRQlqdAvL2o+lhACRg1m
dfJPgN7VN4C6DuVV3vu+sS4YSpXAOW/2VUpgVJUU5NDEHmjCBOedIs4BsH2VsV1i
sBsXhfkGMFPKBEyEk64aYFfrE9F/t02NMCR3I2dVQLw5Kuc7M2lFmgMDBgRj3grK
QcZCWXUVhXn09ayna0tYAFof3gY/DFRxfZv7UmMi825jUnKfBf9qU+uDorhi8wPq
6ddNrZQZkhcD1JjUsiu5QiGDNra6RINRTsoe8M0gHClfqt9zcymxYvyPWiDzUzfj
9LeprHzivxtZ1PDb0roDSdpWDz/5nEDGGRDn+VJ/UYch20CNJyN57bsHfBOrCLGM
vD+/ETxKF4/1KeLKWsx0wJ2/QRB8nwnuBpPDq7jDDR3lQ7whaCgbt3Dx8LqYickZ
Ft2ISbNs4iWIPOMVbi3AiZe3eIbsRpQkweY5CGCCCf9IsOKc6Hmzl6ux4KhDZIK0
0mw5DXbXm8qVnzrq2+SqXuryS+aIVzuCNhvC1c9tJiWtEHT2UmFkh2DcAbVI8OCx
SOA5tqhVLNBbF8s6QL6fK0ED8SA5yCh+N2IdfbpKgj1w4uPPrFVxULgobUPY0H5s
A2J2uCUybm/S2XTby7Ox4EU3AcDsS0q+E9Cwg/JKYPituAMOXUdrD4bQPMsfGiVx
ERQrVSN0Bfx46tOnykNXqozu/N+uO6EPUtI0j0eZ++g7o6JLDRWFKyUlF19Q46Uu
MEcxqrjTYiaX4ppKgWZuZApgp+PQJLv4P7N1CDi8wglZSjZ01bmC9S4d0g59wrPs
LpqbnR/lISNig1GEwTJxlSQ6HEdEGA9kOmZg7NjA5/AMHu9oD07Nu9MSIfa/tkxL
axeMgUsWMgoMB0obNU/A9AjxGBEHxNr9qpxskHSo2zmDsd1IQ4JEni8ekmadoET3
stA0NuAEAYySfjhfFh0OHajv0uLA+EMfAxn4hIFAUvUWM0DA05L+76N1P62tTN+9
Cbnr6kITtZ5oNj90PA1VZCZNDgpqXb/CDSseeZwbtzHNSNLlkmBnSmnt6iw7TWo5
PdS5UEC4tTCDAdACXcOMtHJ0KijPiDLG8l41RDxKiKIwmxTzNOHTjUzZMCJb6AY1
3VlKNxqVhq1Uyth1v8wdjgjg+HzakMEsy+n97J2Vbz3i8KfeoXi6J4m1bU8BGKzN
HSLi/UkuxhdJbT7D4R52ErJVb266hJl5tQoI2NjMBzoZoQSzygCvK7mSwWxaTwyo
AvHvH+yU10FAd9KbatJrtsv6qMkDY0WfyDp3sL6rJW4AZuIDiPMtxvUkWQe6sBxw
lawAFi6TM3x8RRIls6qXGwDi/zMbjKNDcuI14J4F81jsqWWVsvQNYHdnC8Eck981
M2NveJLPL+SSR+5MEY/mtd8c6nn50JkNj48xHrhTGdYko+8fEGokCWLVm2R44YH9
TSL0n4Lb4Tus2aaPVkthq8/NJQuzFz1qbJe9KDOwDbGIA9xVy6nffhnCtugKLc48
PG55qVVsKwA7pOsmYL/EBlyla9jp9bmTXu8NyYi1LoISc/XiifGRlBHfY0TVZopl
iaRxwLqUzSfyRYf1+vxA51B6R71aNy+jZc5wab1QwtwR9L1Yrc7o+qswOwphVhfE
lEVjM8aInG3kjKfMFdRNVJ9Tc+z4pnO59o8h9/syRMkqOJjXx5+5VQ+wADCHbE7g
dJ9jgyrcCRkGWho+uELpYpARqLl+HthuKrrxmbQ8x7F8p+08c0U+QuqHDuO6Ghxz
YMxQHBo5aoDQdRwen7xInbw6Yq2Rw7Bm6Uf79zdRynouw9IphQgsc+nwJCoWZzGf
V9tHreaAAnJh7MmIVJteC2+WK/HUDdJtmB/RnPBSAdfewbU7fIkxYYXP+AtV90Vn
MCvZCe8kvLEdknpHrvWLeQCPtUA+Uq4I+ev5ltOoTI+Ji6CIVvqXd+R/EeHJswOj
Nc0tlcBx3O9rColA3H6Vo5RNWb6cdSkReEAWnSMsAVFr4PlTwkhjkmQVlgVAT4ip
DpVXzdt+sVkz3hjzqwhd8f4EzqIk24iNGVfxxhCuD30Bq9q5uWRwY7pDw9iGjScO
55JYqlz0kj0pmoILguqiJ3VRROirqr2No32d9bAl/2x5d0JqkcHLobugUyCMbHNT
r0CetLY1tSu1desAdJu+NCRt3cE823qklVw7hH93FeY+WJ5JfnCL/sh2rW/3VszD
FHONmuINw/SGHdQ764OrODBLl9UtnjSIsQOh7ai9l21iTiUXV+WEGYnOn7CqNqgp
2mwdUDmtGVGxrb3p8DD9n9KqGv8+5zuoY/7seQUZ3TxBxtzyVQ9VdgCS5YOikEOY
0MoVNMySMES1mJp84USyA7JNKwAq0F/wM6NqU9xwGdhUPVWS/x6dV1VLGgtVddVE
EpB4NiF7p2oV8HqfMKCnjd/CkF1sw3dtU0GC/2MsLV6XnukPxF/OjT0EewytuP9v
EuMnwnhQxUT3dFVuimt8+ila+mgRyusKwzzMi22LPKjeaujCB18cd32LuSwTJ2Xq
lbkbkoFmAH90io6PxjvmJge4/T0CeifpazOJNcpsQO6cqN3V8UnfqgNl3zM49no6
58FstxNX3B59Qf2zavSnLm/XnzG+gY+M5kXwcWaoN7MwZ+I1wCCI/2bItICN9Nio
YemOyb41rl8Axzrs+dASUQDXqysq/9SmiTXsRVaWUpN+wewjnfARy3V/k3OdBAdw
FLdi6RRMl+v+qWxPbAeNauYFx4Fo39AfhVCPcH37Rf2/Wq+Daw85IZjobHlQ5U9e
ridiGtdjTpHyNcPWavLQ1TolJPRh3lb07p+EvUkH9f0BtcMYwkLJlTF5QnLuEKLS
ozvNaLuBsBnm99zFoUVbTw75VkKK5vzIyeh019FrJsg0s/1cGteoJ38F7ZOYPQbW
aRGn6ZfGp4IXMiD/OIc+LFViUkdB6W/ZqHccPbzqqxGpf87/5DaKwqGwHPFWVDtE
jOvwFlQYohR5IAyUafn3X7WpEVRn5+CLy/uHb5XBmudg/vvG+8u5YYdBd+oKsYlM
MH/TPV0vcW/hfIDIvoe7FdVrDtKSmictBrMRhNklAe8C69HT5iZsUpF8JClmGpgi
Ocbj2uZNPNPBq0m8fLKrAIbbgA/MR7vim2Yzknb/d1WCMdjf8iaWTlilPBTSWEnn
/4w4ZEb6xx2FwhBAN0PwEGAlNgEspSEeBsCCrZXToCB+4Tpyy0SPcpN6R4bpNLmG
Fx661UXDmpV/EXkXweu9F9/EpQqvSq7WKkLfZnW7IKNxrxNWcOA0H6V3ZvCJAUmH
bVGbKxqqSi+ZQCyRILwG+zRg9kbIZ45qMU8kA2qyH2+M0jLbdVL3fYkdl6lws0Lu
9FIA00Dsax4H2RgJlHKF03trXfiiI5cg5t95ywka5EhKz+NZcxJ1sEPRGC5J3Ik5
8CU6qZwiLv9+no0r5TWP9ZJlw7bi6BBZxfUml+4f62lo8tMyWt2O3y6/fW4/jktX
FqYP0qNMHpN4uvoRuJXHwNtmxs6wJjib4/WqV+caSbISeloilbj3KXNcNx0wYF+c
C0VrXwZbNl+CTtybJfOmKLC73p4ZoTKtMoCSbSnpYonUUCsu7iH/6fiAnMtoRI9J
i+jNl338FK+Ws1ECnhSCqz8dP9W4ZHU40FwhRQeASW/OuKBCw8K4dd/pwY8FDDL+
R9UH+VG8qNEzT6v48O0CFf65MOd5MrZRs1ZtF3M/+AlAz6+Onhyxw8pfNu5tbjE0
rhUstFAOFgeTOO81ADBcqZClPkn57OuURaQNFZ0Tu+OxDTxWLRHpQ5jyPMiVWkNZ
ZXlFduVHEB5PbV7i43FlaPFwjYWfhEOg3FghLmtlOuX+Qb7nFD4Be5phVYCbyW9k
5dnqF1QPGzwktpca4l532okdCabMNXHOtqsmha/FIEZdfaN5jrAxqgKzHWt27M5o
e9xHBDc3rX9knJsxpW8XAIeanK26q7LU9Zut2Z8nH3QfgSBynsdoDp4fhg7Oi9dN
+Iud1Ew2/nAU1qhB4PNcMwPd2KQG8A/d+/AUqdvo5ju9/olgzveueLXpI4H/bbyh
vIV2cE6TsPPBnV6DCRqSsqrOLKOmCRXfhWccCnq5MMt7DgXa9Cyx/OAeicD/cDE6
p0t4EcJYjAkJn1JrY/JREyJa6OsnlcSv3lX7WfEQFN5xbQgIrFLTUPeH2uZwOItH
Es8Q2Om6a7WV3LzLmahxQ1UmC3FAatu17BP/qRrpmnBawFoVJatXId5vUKhnoMUF
zHCd1L9+J4Nw43nvt/y/HdxG+vTKSKXfCUSYLr2rWs33w2hepjgI4pGr+om3AxYb
dC3ywCzM/CQz87YWZ2uzj8gtcsX8GUq83SjzDTikm8tlZNjN/GB6x2ulf6m8cMyg
3WOCVPe0PON3oHyhkcs3UFr70ZFb4kdBiG5yitOFUUg7I+10n0f+pg74yxqtNwgq
MvnPNvdH95KNN8vHPifRfUhz+GXKRrkkwauhFley3KZ75wH0doW2SWi6nibw1LW4
foIovl8ty6wMfUBO/Ic1PcDIHh/qfS2QIR/Z5jUVlf/z/41lmhZ4ZcdiquXrHBI0
5DHiC3CI45UAohYkFwpl234brLYyr57TXlUzVNhZq//QqUNeyCsrrqPi6/ousm50
p6WD9x9U5J8IY671c4/OtMPWXZKfi5rH9TPAppAqHvmJMWI/IU5wlh9pVnINC0C3
sSosA2Y0yQb+62qtybxmlepuFpBQxR8TGosrbNKFrgg+jsKidJ+7+Lom22xTRNRf
uemaax5YSFxRc5LlEUkPdiZm3SNNDBtK1/JpkiVxddX3Vof/8iUqDyYz0m2fUQAH
vae7d7bmABD09Wk+6tZxB6XjNtawP8B77l/lze/cjJIo5zDeTCEZY+1Qc7R4TTM4
ipu9iJ6LnFC1sCrjnntxY8y1YimlBk9zHcUzaMlb1r4vgc+vZ/0ZsTHLEPbD2+dG
iQmfXY4BmC92DcUz0tiMRd0oo9C9Ixs39I3mgCdn1qprv1ynnGPctLyZmgLw+B79
RUs7DckM6zTIHmLiQLUiDVp0U3M78wsLertLud1RkFNSICitpIXU8VlkPq5tYbrx
KdoJiCAgTKs97wjsMmk6HwiZOs4gBbVQfJgeJ+LykBMFlp09zohUr1PR/A5+BnSo
o8WZ/LYauVdk0k9mu1SRgSWaY7xpUXVze3RLqe7nFnYC9e75OdgWAKH0tKpBmdCk
zoEHwNefI03HwWbAYEF2Y74gQVR2rVGz3XiZEHlr20q94K2qIScewdFdGKwlniOl
eiCtCYaYH2x1p8XQoMS6fMsLxtu1YPFGhXiiafYH/KPwVTYuVj15Icai0BJIECmY
KzYJXbHgJF4uBCErKPqVgmm/465tXfxk0bXpjtVvb7Au98JmdTkSxYNeMdG09R2M
cGPRae9S10+006AemV5oAXa9j1gnUwNPhYDJ6BvVC3YI6bYB0a+rsj5VSqDH1L16
p30Bu85mfLUk1mBr3aW05lAwPKpY8/tnFKIciK1qjYMDzibiYMd/DBXfD+RJvffj
bj19VmuXT8qemso6dsUu5m+F05o/dQ9uzhA0i5EnATf4Ng80/Vb5A3G+7N2TeWe8
VwLMulAWA9CvkeKgExTt7jUBG1yLvDExaApATzhkpwcgyBpwyMgK6MnWKdGBEk7y
wdjVgLJqfTh13Oksyxb5a0trWfarrinJFKLvp1E8TZD/Sm9jLQ3EsCcxssTySx65
9F9FcGAAu3WdIGn8WJMHdNie8BP6ospt+/yDk7EbacLBcC+tfaGgkmuthWYH6qvv
n0jrx0JU/tMLahu4szbYAi4yB1Xe8ZvD3dT9SSvo886q5oI6LhIjDt5rqfyr6pdS
4sGgb6aFr6SGkEfIt0cNK5D6lroRhoNJLS7/sYt759V3o5CP8C6egtJ/NJELgpwo
FPXOO+95wYrXGlMxYTXBb8OqCFOnG2863/4hR2tbyGIiw4duS9fPxx2YZOgqLnrP
rd8xOWFHNqNb3Q33Gg42B7YcwRSrbSWVcjKJttRGRlTJpYvkkbURlNOB4bf/vaP2
N+GPjZ4gtZe/0znR2SZC4H1ptOA7QujQdlKRykvA+q+PgfaCTRzVUKz7hLKqMJZT
Lg79+nsrFi+RRl1ltIyyVBoYYGeaecyAdu1vaSd52I11VxpNqb7V8KO+UOMHyrol
ocJKvgGJoLvxXRhBx2R0PM8ANajwtIKmRWMSFcyGjjPkb31V3s9PQLqwpQePz4X+
Sc5h9VHNsKxUReiD7xzjnQf0KQIeQLrNF6I7A5a+KE9SxekUwvCc65rBnKF9siTp
9C3Fx4jBQGonGYL2WhhkFQkJufq/CvC9zYks08DEII1idoe3EX+obMccnjneBv4j
JPn9SuxcZ8b7IWldglSrrEzD/aRN/A+55bwOj8GkNUcrjEKaB3SuNXEUw6lqBs7x
V/K+q8ZrB1zLAwSLeh2cZ/3LHBrBrqvGjtRhhEgdgO7h4R12STArpbqbpMJXuNux
pf9/Fa11Kf0uwMmGHbHTWDmik5BavHIPzLa2JA7kHvUHpbDqF4Mcah9hl2m2MmvN
Yaw8DyUqAeOBM/eaOEIAp7OEG7NM62uKzgB8qdQZrVHGBTTseILNFMOSSxMAQWK4
EjLz41ch3vofUt6XxrNzLvL6XCaKEackLyXy2NRHvv4MT7NqdE6mA7lMOmoR9wSy
nYb5vTUGNza8beHL6z+2NjgKvmqUW9Ww6sEJ4TxOOVK769i1J4sJ73QdQAbMz2UH
6HAquoXaoJptRUwgToKHq2UoD2vMrgr2TaYX76kkW0ux9zA1LIweJ5h5Ky8wn+4r
4Vzg0SBUsbHMRoPFtHNmagavx58Ks9FmZJJKq/abnieHQVw1aXCE3MS/gJN/XQkb
za+c+K9PHh4unt7G2MRH8qrE7aBTebxTOqsUW9814l9JmWwhqU7DshWZUQELpyHC
As9fm6UID68tvvfv7mQVX+RYDoW4wDFPoQPsIdjizmeAGNilTn7KlAs7m28egNMJ
HfqgsVDhjE1pLN+j9uNrlGSp08J+swjrJTr8QvGbBciy7lc/72bnrs66HDj0H3/1
CmU7pu0n5z1bwVKtlSaWJZW9JMypCgGAViPfU4DF5Cl6hibKxSDQicHRWZUE8LOj
j2C1JKQrdWjhPUdnIimsFLU0zlxI2bc+KgQSpKKwYcYnweJrgsfm+TZ50IRqI2ZN
UOiWr45szhHsns2DASiKLLGjUwXIO9vah0xB+fPR913Cxz+qZtbytc5go0KBLCNI
14gTU6D6fLXgPve9xdlcKKrhRfNqaeIthXFn7xQvDNmodICTrYomzVdI2LjWLLc9
HjOmngHdL8dHnqCcKuoheZTlceyG1sfVd1qOl7P/Tm9OhG+tT1+Ys27J5Dpuw16m
kWF2rYsP6W8X6YboNJ878Gn6FcmhatUzNB76YjF3W78BvRpBRcTNpzx3+D/JnRoS
KgfOFfXeIiT7yhq4l8OoO3b0hrbIHgohq2I1HyBo87iGFQ8Qp55aJELoE79Dbp13
5G2621tB1AGQDbs5fqa8RnUZYb1/aU2omkiPY9PYqnVUqWWB1I5rjcdntwOOFkF/
E7H4md8XE0P/IBUfUIGC43MnKwzjrRRYkXLPvouO4L1Z1O2EEnS1owaKqy4n4+EZ
ZsQtJGDp1glCOC9jT8mswjEeXIMR8dwYOpkm/KvGs9vPUR+p4/Q9hn74ZR+lHiX1
/UQIVAUZr9C6AkJOD2lcDk+2mXcjYVLJc3M4d/4alWMVX4vfR4uQiEaIiBVenfx1
s5MpaHEzqI+1gSuF6HVbPeEMwI/+ePymqWlWx5ullG01y/RgO+/p+qQQiSlVFC3Y
ALsIWFhXjjFh0xgHyh4nD23CBg19EmE0oa44+Qbo1znDaY0POj0rO3Uc57Pyi2m8
FWBNTqN/4aLABXtjRQw7hWGL9MiON7iU0nJhtbaf4hGyH7Ik/SrVrikAMl6tDR28
pr5zoeJ1ugtDgNj+rhoE8LbM0o02YCiub84YQYyVabujywMdcreUk1LixPtwmfCn
2UaRazuN7TlOunHzlp28Le9jNk1YWLyWqLv+akrFmJu8tgsU6yy2Q6ooXaEge9jP
JOADGnwDp+zfDB5jOrtMD0U7CepYx0OBMWhpz7UaxGTkZu7xdFUKnkdSwm0aP2tW
0fuFyimEJeGxngepLIw/PxI3VrpaPB/HvcQMj70+cIltUJsogqlbm3FSrlu8ArZJ
6VfdC8WyKg5ugN68IGq9hI4ycymGC5+vMLHks2LK0hNta/YYjPlNEjjAvcLWNRSz
HkQx3QBtwuN8pipdXB4Edd05sS69MF18K0WCCmbPPu59+8y3UyNp2U8dKz5ztrji
JzHL2MUqChJ31FOpqaN5+W84CgHsRDH5q8WthGQwM2xk3xpgxbbrGvhmJsm29bYP
RSlWGuhPlejywXxR3iFxX8cjiXTc5EATSOb0sJ6zmvS9+XXKUjWFG0KgnBMkEBNR
apAoWuFXO4wFf0MO4mAsYzCsYE7HBHNsr1XKNwkOBq4o94dsgGjjSvNOH8Is8Cx6
bKHvQ7qgmHkxN1d0G0YFIwyuxGsZhPXpj5P5bfj8x74u297w4C/LNWrYeaufgmW+
rkesBB7zjFPnVD16zN8i1uEWf2wDNKW8xnxLQ//4mOhfth/WD7JsuYyHm80DxPAr
i/7c+ThqwfSYjMt7ls/Y5kx2cpnJDS+PAyT89H8FlHPqwSPDoCJcwy70fUPs92we
Ugp51ScAuXfJ9lhiUABYKWa8flkaXmaGb6N7I6LdXzveY3ge7t8WK6mw8E6C8TUp
gF/B1tkoqIH8f75e585tpi7A9VJYUdTMZQqSN71twZnzggxSUx3mstIfip3tk47H
Ztxa60wv1Ko2MUnGTrWejDjWAZge7V9KZCrT7HIKIRBPeanKvrHSounYFcJRFCAW
4IZqAEB2PH+kIqmbdvxQF6Z7S4lZ0e4FUNPaZGHiM6wYAgyx3qe+Q9HV+oY9aC4m
scZPuKk5JbaTXSmReIHpL/50bmmREYS43sZcAw1xRINExnY/FjFkLvj+ANRINCmo
UtNonby2z6soSQo/eYgIOkBISJIg8zgv2vrmhzkRwJAdcwkMqOW8TtboxXP71H21
PH3LPkNvRs+XGEfa518ObJ58rbDUOWP7XZ04GZ+AizzbBZLyTvYqm0b9mdg4+9YN
TtlJretiZgPItP/KEmWXddpGl8zh06RKe/zCdt5DZs6v6lXwRsOkk7wffxFpbghW
TRx2QNG+cecAUQSqJFfdwPYYlJc3ZN2O4W5VJ8vMEOTCKxwUsFcNya9Z8+Of49PN
3yd1tVgmzqoIge66UNDrI2o0sRFxS3GvPHknBwDAEvLM99lq3PUgSzXmksVVyvor
93PwpuGnEsBMQLrF+mwp8mokqmcz2nolX8BI5gA+ldpdt6Ep0d5jbU16GZYdCcvF
EEzLI2E0NG9jlBjTIwkb55Kgx3w0+DuwbsW5v1QqW+LcS9mkpoWC0MBuPy77c8Hc
G/s+aH5+zVMmsYLaaNPPEmBPPwLWWkSPkjQJIEKAT7J4GhGkPFn6yde/sgJbv21Y
YrBNF/tZ7HcLKOAJM+qrpetnkECDk2MBxyHHwjoRXNUrCAT5G0WxNoOgLZ5y2KN2
1S00UC7rHjf4WsUmIeHrWMjfxQKzGISh4phzK1G3h9Szx7RaIPPLXy7Y65jbhTtm
bvfoZFDIFbEaWPO+68ZOfQWLP6j3038JkIjnyCN3mbZPd9FZS45zvnsldRf24w6v
OHCIgV13P1PTAobLGweyPUKCi4/JhqEhfVXH22dobnbLKx0bkFVrVvx22Mrql6Sd
2k63hr8w/NsQ28TXl52rUSEoa4mncJPDm8YDGkHUMRtp8WzUu4qC4iu8TjxkcRrm
1u7GR4X7U6dEhILjVi6tp2lQzU8paRE2ysEPjrsX49+r7KZ/SMSDvcI0pvNToTd9
4zhO/7vi7+l/Ft9AxUI6kNwax4lHvi2u5Wxg/4FmcxeP7Mc1k5tQyfAjZVjEOuPw
ssLjH6ipXIw/H+OzmBsKge2L0JFntyUHQsH37Z+qHc7hx/MquVOY9kMM1j212I1s
63HM91WWqKkY37NjGPNebhoLd6h8VLrKbm9NAfbj8foHZ3RpzKGmL3RdaIk6UZS2
uiQMqBb02XrNSiJA/6J51o0LYcSKHmIEyWSQdsYos+cGFulc1Qb/Zkhpi5Klv+KN
zXOFkcadUpdfvFeFDIW0dNCT5JGG91nEMHTNSDxlihDll5vySoZ0MiWGRn8it1Hp
Otx84shkSlF3NmMEUjC3FD1n+RVF94X9iMEnDS/zEbFgW7/3Vrkv1EvH6zNlc+LT
1WBIdz22By8WPjQ8BYOQGv5LejEXGVBb0RHb3UxLpg4HYifsck82J0jHqjQr7WXV
NyYG1cIlCY7RdWd7prR4TYEo7v0WBKN4y9gFey9UyE3KhK7BB/FhXsjkQDKFjfXT
f6sX0VmBIOkluibq/JPEVTwa9pRE7UBJuHVQkAJHwiJtVc5wAecD8AdnwnO43ice
PbETLnvHRsyooDFqiCuTGjAslqEzfrihxdCio3RCQ2CT3tFSDpRVNV0CIYHqCnFp
kpVhD5hIBW4YfO5yqRYFJ5PoT/TFSjIDoc86y8IfsYGoWJQdo07Ch6PU5RZ1pt7S
QjxJsuU5FI1uMOL+w1LThUul4rfaJqJvv7a61X8cSufHWsXw7lpnk6cDQcmPuPPq
Dq08W8oZwAv3dh2cebq3SswvhVxucLchzlB7tjHVxt5Ap55rQtrxZNllQziZD09x
cH8FODpYlxInIDmO3RvGaokK2M4VjKCY/0/ZN+5YJqJxZrOO6dJJOPyl5C4oUhZ8
Td7dqfYc9T53AzqjxhyyTAbCEHNPnvkVqnYqHFAzJ7ldxscYpAl1qWkxVH3CgmMo
LhgXzIIjrAT3DaMED/ZfNDFsUARFBbKGyQTa382zPFK6gek9NoqESVLJRtHVe1oW
sZzxQagqnuQ1FgIZ1DjKo0z4nVdni7Kj7VAHRCU2s1gdVZDeGKvqnnsv4Q4KPiHn
cfOaWLy7+RWhUp5JHRMtjNCqDEw3bJ5rIm7hw/JmvVegP3taWRk4sYP2V7c76qcJ
65xLFYfQ51/sFjTquAu1A08m2Shd+jp3q4qMpn4yaJye1RlHSI/Yc+9O0BVWNSlx
egzPHh5ygScBLafbkizRXK0pgp2wUwPSC6Fudbb+YzqbCDBIeDGYKwJm45eXzcrE
OdjPz/i3xDh79ekzdCVdaCoXA0w5cUX1pbNzSRTQziFKN5jgfvf5B0dQoKYfx+YE
bMTaI9HQuTpv6/BRhGQnA5cIciYV6/+LZ9StCZmXl88U4e1fcIF8Mbvjmx/yf1tZ
RBauN3PnPq0pzH1YhRTRj0x2ZWsBsHFGmkZKPSXFgU6Jz1FpyLAZL1z8kbAKDpiV
I1rQtomOtlkeb/NE/49QkcC2xAwLQTvaCQ8hY8fLmS0wn4oiwA9H+awZoFVe4PtJ
+jELj3EGldjhYdmGr7/iBgZUeqABQeQrWezDPp9HUgtYGh+OcfHNNqEjY7Ahcuh5
agYMb34hpfThnOpDcmgtwZ++geEZZw96C7Jq4icQO9pYcyvRuAHFj1yVAd/AOA4y
E5HfjvnLyM0dTHoP1/XKYlUrdOkrIz0terK7UNDRf9SJVryy3o0JcVpwHMRiTRvp
cwJ3R4816hvToLlf1fmAXJKZfYvWAYpeLczV4TCCckNV3tjHXDxtRqAYuEkO0gRA
w8OgksbYLTnd87tqUDXsBVNHRO/p0TiGlBU9RfVhuWdLqn2uECwhyNoIsNI40vuK
jwEVHY9Fwa2iaLJzbZtZJkBMiiELLmnDQTc1OTmK5pCsdObKuELSsD0PZn1wIKge
+VMOjD/Q+h5a2VRMpXdoNgJUVKOoiZKflQFTHBpUwtO+wa+lsYoLCsPsVRwz4vnP
TyTPvcyylpylSaRra8mmOfDPwMxrEsa2sHDwmar6FfJSAaoQw6ZF+HDXtA5GMpMg
po1X2KcmcG0C3IvN7jQMzpnWMHqX08ReOaV2IjvT8ZNBRg8K5p0bmjS3g2z26ybm
eDkFaXO8NcMM/vl9sCreP9lXyk2tjL9hhtK5Tru7mptlwUoKrsuPNX5upBbk9Z9q
2XVRsBD8v+msuBNb02cRcGOJ/fRPSMWewjeSll3NlndS6NP7y2rhMI6DzQIFFy5V
HWA8JvswIR3dYV49uWGCx1SQ+gZy5xclbXovdsGTqIq8vYCeg9lTiNPtmGu4FiLm
H3+EBw+83P43ijIEVV/V1/tQdiHSe8Tv+7GqJKX9Q3aciLLkP91EwbrH1DD3khIF
fqkPcNbfMuFBjhWslUQazAnBl1e1It25jqC1Y1GqleM5VAZZAxu4VnjT1GDSAJpF
VrjQ+7CyfkROirqFSFAPATQseBov9FDk3qzXzT7mBZTPPV5zIuFbXX457FvRRMX+
UGuCHoDLFRmdv3lbIN58LDtM0qtXU9c6wzUvDHK24GzHn9XqceHD11WlSdFFXKFi
wYs0qIkc/byIsF5UEiPpca6fYoKM1f4PGf7kCP+KBzghkAaENU8L4z+jlwqohlQs
dQ1zvi1oEo9/NQq1Vx8/nBRzKw8VraIjlSj3ch9TfY+6J13QjFTmPWJP2d0Tn1lY
1LvILVTLf6MBOMfI8xj8BhPpOtpX0CXDN80AqxV4YffM3axYwp6w5fRQgCyjyZ68
Hj/6CLCM5xaO140cV9JL/fPNS6GEZwhoAgF7yJsFLPaTIvoMAS4KMrXhRCP7MmY7
g8sAdEuYXxLlt6L8poO70929uswDGCfAkitOKk/enRB1M2j6wBCQxpUeVeVlSJ3C
St8xtMXoHyYRH9keRM5ChK4zZRNSSpHmi0cnLObQB/AKTK9idOSJ2KafFXfxYApz
n5AWjB0fg2DIsX8cj72ypoZU+nVoNgW5isdCpk8jK5ubh2sKCBQCn6aR5ZkYiUmW
g1E4Y6XaYnfeMqtwZ1cRetRZrfgc768BvVWedoU4WiW8U9t4gzMYmSKcn+MdHBBv
MPNxypEmOQaJJkdJhHtNR2ffFmI++LqjX2OHNUDT49+hsVqyRDMKOKXjciBlHMRH
kNuWMeUa7oxJ1dAArFa/CNTRXZmyD5nSFyeU9X/dt8Nwqvgq7gaefLL28TVtKY09
F4Ol7uijsxwS0CAuDk8/dzcViAH7MQ3QpLj2yhoB8vUp5KR6DIAEFrmSF4JnN96z
9epd8T627bIcEDpxHnDVRUFKqMboK9VHUbj64EYrDf7N9VXWTAhtgXV2dTpuici4
DwtoO8Nho1CkDErfOJGDmrz0nZkHvrl3TxzggYKknowAvBWyXq+I1p+i/LGO0SEN
GETDbCvIjQLmqCW1ssWq3rtIKJYslRCGtCsKbBPIV1fu/6X/XhC68CtJJaqQkxC8
NGDidKmSMgjaCVksHvixDM+3kfzrMbA8XR2RL3Vl9uxp3YBQbgjyj0aZISljvaI/
aZ7+hAR//gjwMz3adnp8eSYKpSjryYIZvHkRq5Sk1WH9i6g6LeAebCTfDuYAun0A
Z2upMZ5YCSFS9S0m7RNOlBRvqW8LvwclK5rZfLJrVA5Gqn7UcKypDNsrduRMzm8Z
OUA0NvSg4Bn9/A2foxEyJ9Yn9jHuEbyRWbq0Tet8N1i+WNEFMztwXTMxb7R77VAE
h7eSQOnSfuakP4yNJdi6PFYNE6Y++DWBJIYIrx1ZAvCd9UE5ubHejW6wCTErO8fU
r04n/GXTJQzKi4444mS0ziP+uSkb0zjXqju7vsjY0lkK3XePagrtgCpezjyexCjd
2oOwGMpsvV7u1/kEv47Fc8jaaDVL7lnW95t8RVBKeRHtqWvtZk7Hmu3nEsGB1Hqv
+hii46z80AOR2XnZf6DlY4aq/XEFTkuo200/qq6V56rr4PQAtyN2jhDapRayffcG
afdXcwFf6BrlNGsGprKdN3kT/PNu4Z3cSCiptEPBo1JNvEiY++WIiw4DfmncS4O+
zfdDREN1axSQxHlotidf2ndKBWQpQpTv7iMrecl7Gt0c3WA+gtnU/NBhsBz+XGF6
E0V1FbiuiQJ2MUunO+ramEPGGqcadOP9TZGmn35w0CcJqlxP1zYrfLjmWJ086iyd
BiCJgStmn/chhIbNBmk35ZWGaAyo5MXXBKaDFJhLpX82mRkqt6WeDnRWXGj6pASy
xTzu6YGc9MWtsmmJmigqrmiyGn/yNea1oAXBXDHu5ZgLORva8cudRzrr3ZP+yZdE
0ovnLvkNgYYbHjxFFY7xFFwqnjL6EFhCa0oVoMG5ed1vgY8VXU8+MAfnJ7RLuXJC
QZBnjKT+igoARNSSS3sLW2Y0XN1tkszU71awRdouaALjX/WNFRPQSckp7hQN4ZQB
Tk0soE5IVwA3gFoBrqovPkOCIN87SEqYw7OGV5WQMcI893amfDOa9etcfBPvQrEM
Q7IKVW2yi7EydvOV5SN6S50UHPdLEYCjtKJnrJCdVRCKVF+aiFLiERxTHiBy00f7
luLEQztFz5nPh3er1cdChjVcIPT6ZlhBAV3pDZHP83Lg72wjQbmOdg+HlU/Peikc
qHufXXyBdGLFrhkatLthScm2OFIFBsSHL6aLVrJTew045YR3I8DOFbidF9Nb50cC
R5NzDe2nACMJGC2moCiZsDbcY/hc6VN3qg6vgMZdW8aFZHivO7heeunBY2tdpNWF
Xhstvtveu0GZUNFRgeVCgXAx/21hdBDLdMLWUiphOGC6hR5aTuvtcPWiuVHHS9bd
mKmD+p3fzjeFZd4DqhsaS4zrms2w2I2uE373NDzyUu/ARwnjW+1WFJVIys6CUWSi
LSuLDu7ycmIeHNFJX+WyDdze9m2HOB/gJR19wqrA/2scpJlNpPCh9f6VryT6KyWf
+2DofVud+KEhFoFp3e/VnZ5R5iflKUE9lKIwRpzdyoGc5N24sKYiz6j0AvzoX1SH
vYZerpbJTXTg4DUdO6fbdgwENpMS6rMrRAG+LkhkyM7vE1x0j1iD9bfZHIRiWfYL
FKa0/k76PHuZ7EfpzHRJalMslvHSRmoBTGI+ZGUmXixYXxGHx77Uq/z4lNM47PRW
zRViWg0N6H6BsSg3DVTulc4m0ZUwrXnMDZVRkcg7UraD/HrnAjKG+GNo3zVcMUju
pZnr/l3J1LcAUluqQeVu1oj9Rs2WgxeEjovx2cZQW5XgGmWab0mWMZfOgUSZGrc7
7g1S0lBcCcqercm5l+fk/6Ujo1uiF2hsq4QyzzKlNPklgyYOrrLFLvl39OE2hctx
QaGE5OjjB0zWUaDSQyZU+HZweefJe8Us/SqcIrGhFFtPgTu0WxBO3HHvyrd5wxPB
ppJDk3Zvs38N/NQHWHwDIWcwK87BpqUaTP0o68EYJpzmdsGHBE8fhQLPt4t1SPTp
rsbK58tECILDG3yLT2ZikfeJIcXT497jfcMIU/1BSbyzj592w9Gbwih9q22nfcz2
vo22k//GE/oqgo3dOvzNJum1eDTDJs6z6JbvIyu0KfanRE6abiZ3gUj2it/BP1d7
Ztsmo/DobVSdytRi1KyTXedm2tnSDQ30QbGR7UL49HhnmXJCN8aOHFFDhW0D9gOc
7OOhpLPGkGxoBnVIfZcJGt0XXR8Lennaqoz8BoWbilJrQeMnyAxRRYNueFbxjYjR
ZZK0d9s0AX0y1QominK6kf3PADVokfVoEujDiav+XdUnwQa80HJX3NfnYEDIUj9V
+BQtfX49QQzc6yg8hofk3JcRRyFkV8UYUJI6PrK8MB+CbAQW5SUNiAcXeoVLEubI
omB58TcwprCpe+al2mb4HqinYmS5tL1XHFfphdNUpQtQOJIEW85mPgFiPfFbDwH0
+kWpxyIhOqdN4NaIFzs27jXAB9pr6fAGF4Wezf6BJrmJrjRumWW5ILql4CSnJSpj
0I5atJ2jkcV+U/V+M0RUY5lR0+JPWX72rYCIQpEEnzNeCFWTZJDWYtrqcobRvd9V
VaMtpkaJxlNO4Z4PAibCKhu60gI0XhJLoL17isoF1nFTSkubEw3of7RBuYnxqO82
I/EQ8B4La0L2ettT/8fPXWLGfUITN5Z0c75jQubEGY454Y+02m6M7L2ogZW1Pzxd
CyQ4wnn5jxDXRHZCAIvi1EwkpuNDBOJyYf5+2YkoM4nqVfmPMaq7zPZmr+w0XcF+
jaqcpVPhP6QWcJ+JRur+Cg/t4u7uICTCF6pPE0fO7wDBt75w7592rLVUsAEeQspk
UM/k9YwE/A4kUKSTHOPwp6L4iYIGEGKT7s0Vs6ySyEb+NFxHcJ8geocw8nEiQ+Eh
jHIFQq7j1W+EfC6T5DGCrAt0BuYikH9wBtcgLsQKQOynFcDn0a9ZHS1E3x0SP0SE
yChFa3lj3Y9QZG8wT2rBbyjSzbsxQ53HybVw278Llno1bV/hSJHtgz0M3v6dsoFy
1hvIGvBW5ZR5FqOQuRQdLq7dZBCyAY1u69ii74T+XmvCHr3r08aQe/k7ki1EACR/
tH628V45MYHqSX62bN8EoAtSK5ZA47sR3OTq/TP0orRZMomavrSWp6Mb4ADcL7W8
6DVVCohxMzxmNGNfWsNmhdQzCWr9SQSYzIeH9qMI9hMGft9UPjTviAEFHqRXTjmq
Q5NPAMnEwQLTVIE66WB4s6IAD8wGYeW1V3VHXVoLxjKZYMToqTj1rrQ9i/BQFPL0
6tPszy1wdOjKZEfSivVPTl4t1GSkFm4Hr4nrEni4HFaMU2hM4NriNY58HWxZEyJz
7IIKz4eHUHxAcoUi8ZeFxNZcrXyXO2q0NvP/zPkrH+rObYzNmKrC/DaOv7IKSAPe
Qh0o8cZ7z0ddF1Lt+6dY+HcmV94AfXBOl3+o8DKLiT4enlra6FNN1+5BE4XSrjM9
sELdEweBI3szQ2r2O6UAj4dhFFKfaOAaE41EdnB+kZwF2tHnR6CsPV+/V4+XcNe2
RJw0npsQHOKY6mx2yChFVDTtXiTQW85yq6pTfJ/jS//KYx21rzgNYIOM/mS46KL4
LknUs7Txk0TtoLVRyKZCL17G+LTenqdv5uLTtd41xYriHKBYUJVuv5SCdgwNF7Xi
Me3ZAKoW1K/gH+YxJRptFhfX5PNCpz+p9UmP7Uufn8tw13KxZi6AYwzXT+HlxPHm
/SFhHT8VlxA39TgK7ewPFJwx6h8zLBSn1vRRs55As0CbL8GS+cQ2G01FLK7wxlxY
U6b4Wr5UsqpxWDMYyQ2wizLttfw3SfUzdxjO+NTW0FPOsnm18UkjNUOOHb2l1TLO
/OF1Ap3PoV8+iBAcsiBzY2WgvYbKA05Xf6l9veYZWWAFFNdc8pc4e8urL0FmuZQf
C8gSxvmhzy/W2pYd3fPzxnRAxt02qc6X0vWSSHk21tIWocdwaog3Q+fzcga3F8y5
8KfJoXM8ITo0bDf1/275sHZjajocAd+b91yEUZikcUebiphZigNXzjRyWVStG/Zr
P6GTzbLGWUNToUH+ymkcevFJJnaU684IH2Mkk+nu7BwslzMjJUAj7QUXgN5AQ7Bj
wJ5btGBY3tq28paUZMgnBp02evFjvSRKcWi94esNC9nWg1iMmbddMoxLKUJzkC0c
mVtRbbbSbOYEpFoXlVUP/srKl2SHfjTaQw3Dm1CSC0IUTTTf03NqsJe964SluUh7
JMyyU5omJyebPa2NgAbIVdWvTHNGRtu4S3aS2kblLPgSXvCHSGrIz3xWmoonqAkE
9eDSiO4rAILArjqu4gUEJynPTnABSMPvshj+lefnenIUdF8IYzvKlnSvsSu4kx9u
H9EfGf/9mfA/JZkGcjwBhpX1oZ/LHHKCwV1SZbfxGra5m7mg1XdJYSeA03U+Jmlm
wxSCmBDN4tpwaST45K383kQaK/dWBzD274RhmydEfZ4eGl6appMQ9qkH7bQ8mtRk
Z3WapuYaaKp0ghN3QjG5NEB6rR4AX+XSdmHIlhm7PLw8AKwEmNva7HNd0uoHm477
s52AwKsq/Vv5v5kBr1oLUZt+orWrQeQDE1LDguoxaBW9OQHEV2BdtpmKGxaZ6/Er
h4j+FhzBsAv4gogZn1nL3/s34hWu/W1SLeZW8FX5qHOd47hh/oa0piJ8NKjkgDRa
+qExk7NLmJwxCluCqMjTJzJnBPlNpstmCIdCxKEdH1BOm0hDOIq3vpKFphYSyX5U
ikyvx23hbcnQEStdCXwVmwhvAPfw9v+vLsRxrLRv2R/305lgu94WoYwb4Si7Rh5s
9+dzG491I5V0dTyAdj6rQKZ9ijcI4C728DhSItVdAHuV8xiWoBxOXkBtKwyIK8vs
XSn3StsSzBDqLBTqWOjThJPH+5C/4NKttBQ/3WX4GH2/ofx6z7zqxNQWrm+tGUW/
iegQ2Kf+GxxTlctnprXmy5lbLkHTaASzNGoiZHfC0Lowci3hixvdfB7VF6trKRCC
FEob+8OTUPks32yIBEbi+iAMZNtFX4zDWY41+2uMYQkLisfze563HecfR/Uoo85/
vQtrL23aPltyvMtRVN1992jrxhoK5bI5TlwWgaUkS0DU3lrLnIs1W9wS9pgrWkyw
G2VzmQvwsvuIVDKyMtsE0VbW1TCzRV091Ob8GRfSNUqFZV7NmeO45mEiUpj1Chf1
isw2ndth2/kVbH8FFVn99gxUn1v/iR5SrvrsKExN49mnQ+zSEeClYwSfBjaMuNMR
h4B39gydEd9umADUrgHLEusELpnO7DM4VGi+APCJ740az9EA7JoLZvsfvwq1wgcf
3FJem00VPQXnGkU9lEhOOkLrsQ499Wh6WU3w62fWn/dA88+0guuJj2gL0woahhwl
0F2Ys5PJJnAcwEmHXun76uZFYg+YFnMyzSAvZKyD6mHbGFDNE8Sqcd64dXuc0cah
9Bb4nZGqUBuGiNNReSXf+9hq7uGvDjcHSFyoOxN0Ur2pozVtdjqsFbSB1PzJrrZn
tQoE6+TlYmupomzXlzNInxqQwQxRF6D/s5T394kcheCG9yRMoXudxp6Hhoq4OJIF
ppmMMbhsPjaottqYnJrvDaOxWXeUMxql4yBBPXtOkdlEcUhGf7ObFkRVuRMnTOPu
G4TA3aMGOjYhpq7DzDyn3EQJfzCgE3r6Y6TRkvgETJbS/sA1R2lLozKkVnDplj+A
AlkE12ereQkS3dqV4IRZTTOgG9DIt71+uPYMCdhQp8lWRlAsrZcyg1IwRcl/m7Ew
vaLVQn0hPWpLCBobruJwdYfDWiXeHG2hC5nIr4uo6VVuXww5gG1/xn63NrXzbaKS
nsYOTG78DheBjiJbNFq58q3sMdK0wUo2BaGm1K76in0FScIqNLCawA462hBC3/4/
aPClQqs8xM/5NNYEhlZeIAKQ/BVTrA9wMmGm+jMxLokicenVOZ4YJ8ne/J4mZ8be
iySJHWAFdJftkzVLrPBU10atBwXOp732AQ4fWvqxpQ2BAunNX+LvdRrustvj8fx0
IMlocStWOCEBZagp+ZvKQd8UOnEtpJ02/OshlBDHTLP0Pj6j/G5gRn2NVf4L8fIx
5jxSFeT3RXQ0b1ypc1vHzGOZ7MXvou0BPXVFHPk+7gM48epY5usW1YVhbM7a7QB4
NU5dczUFDwTlwZXhN1hJTbKtJ1h7EypPpY5DZyQmIYWnsYXZ8hS5PstcVoLJP2mr
KZHubz7CarwkFvhUJ/BmleU3udp1yRAf4Q44E/dHw+tySjT66Q65Ce47chFkGG6e
m9kaasLrFP+8oBg9AQ+Moqn2fhwGlVhRNUp0umuBQ55vbOZaIKqnc4qeVR0NQTgx
hnOY/I33BFJI6o8MIRPW+2RPgkgPLQZ/uXux6/Q1B8pdbi3vkTGRW6GpoQWojzHl
kwwbNYNZZjR9Q3p9MeUI4GNivs/2SnJvhMnXznV9j8jrugVUwnlsscpKKgXdKdDe
Qq6hox+9Cwq7RSdPkwH/CGX8LskC6iajQN2FdAbKURNpr9KlrplYrZLwxn7H52a0
cJnWe1rPkyuj0seG18AtFmkZLkHLaJPpY5qmxSJMchmahONTaPrep65RzXjVaiK5
y9nnDzG2+YY5p0Py2jyi8LOHdjpwXSBOuKsgL5czOrK+bnDy9+G6X7osCaOSvcIv
Co+/NSi3WK/njNCYuUDn3kTn05y64b3FK0SkNrIiRgX+nN42SG5SczOC42WqL6qf
CGOi1yqoti0+s589NeA2cfHHLklD1gKLPJcBG0U0tmda32OBNczaRi6BuWP0kByv
0dcvN76nkt8s8KUwWa8kQlJm7lVKBSMtFj/V9AF1t/kpDIMAokpmhFYVPk2Dhr+6
NB3SQfyBXZcvjM6e8wOLwHSKvMchbJjOJVh87GG2paw0ZbK4GNC0l9P7Lgt7O4td
syrXD/Q6qsw1po+EB42yMHqend1Id0S99sX8/PxhdJK06NGl6QlglEsahgG4iMBH
GZSs5kGoXsRETNQw+R8i/MdeqwjCY73z7zkCcT9PrcZnMvj32x5T3JBjH2hk2ItC
tx2gtIcKaryc0rzaK9a00LbnX1y9mGQV2ce2yatWwK4UeZf9OJHBkw8rwVK05uO6
J1aSXYhEH42vJODfjGyVwj8TAZIhk6nhCnLuZo6uhTY1rYSr1hapKBUrFghFwY74
Hv5NTHE+vBoxQUJaivwdBDVCNusJQKLS+wEpcJFhk2entwxTVdMTD5xjzWbyIlBN
INS2M7+Lotqxd3nRlquzjIEaif0ngj5KZxzCNxVH64I9w8jITEwFKA7WSmIlaLoG
h0csY2hVExsCk7w0ywnrmSQJ+pg3c6hzwibMZQGXFGlYAIms6dAwCY544tFtaZdq
qI6kG453ejchB6dNpDcbqRssFUyOo3N2llPVEfFFx/Echd4kDYe6jxnk2td66QiE
PhZ4ROlgMu3eOlmYkoej46sKAEnFSuXKgzBb56QW94kLKptBNVcW5buQUMyjlIfO
muCSXl3LLBqJsITJh7g94dfUXrYJuSVcs9khEykk6NqXpd4WhiqCBysPDYOZii4R
fkpgrFbyXkzfJo6v5FNAp+wdmfwZGly/0T2z/3jr+6xZtb5I5lUpWebA1VHzzYw2
a+bgL93kzZUbU9SJhAItlDGNoHGK0/tanHvABnbVrE38eQM3QfatJzVgq8CcuVlO
ePl4wzQjXukkK+YrdXWOdJCapLKS76wPuZ2k3VxFMmAGmRm0Q/74c3g9ZE863unv
GEbdUjM4bXpp3Z5Wj8tTmQA5uMv4BsAaJmiIRQ6xta+ZaFKCtSxJnLke53bUXv/h
5oIXjOjybdXSH1gdXrxwaFDAzcCg7JsAxdjULYjiw6hFEO8/0vr4lNj98GJD73Mn
Mx4HpLr1f/aKJGfc7bdzuLntPDJ/urKmW+9wUoN802kt5S0nt7Dc6IcsNxKvrYNo
hon9/dLZ5KW0mvMJgikk6I0bAlixWVUpq77Kpjn8/ZKHuelS6mtST1vWDQXwzXS/
GIgHg1H/6hf5d6ILF0obCS/RGUqkBcco8JbObWAfWj4/fJ+vUCR3Hi49PBM/Z8xb
l4J1TvnDkRYDguemxNpGxqwSgwlIZdLyDZh3pj/7q/KoqkXqyLDFvd+4ODTYXa2S
H36GFyYcwDHL221ZAzsx1Y/5nwjkifGYk+R8rrZyuQHQ8+4U8gZg5pfR/+DKoTXK
VafchArQRCNsfiNwd71OqFw3dGCi9mya45fyiPJZaTCINjZXRWA4LCMZplJg3AvA
dXbKgjb2CN4eM3wU3T8/u7+8kWNvPtjUq4CnY7oFhEBItrx/RdrAY2Zzi9shvEl9
EoHJzz1dUIcIrIEibxPkb9v0GgQcoSrIMxku4OvjY7Tw2jkG3octopgCgGRN/oNd
VhTM0Ep53zZMCF6Ys96PaAc4CqOSqLKFWC05Y9fPjV7BrcLAD9Mo9up0FcDaYPCh
JLcEsrMzcCF+AJ6eR75rq/2xVaI1295nFk5+0TMjxU3gfimHKI3zXt4FjMKVs1aM
ee3ShfTWirThfmSF2NdvncqXgocb3DdMIM8sOptUrssq00T2utwySTCajehXFl+b
XRLiNuzwvIOSjnaRlXXS1RLoK1u7Z1QDNQxOzq3uwYo4lWSHEWkTtHQ8hahHMaFP
DQrk9t6qnYeK3ID9eKrdmPAj1iUUkS1CAC3kCMmNCzb/SWZP3dEhjr6SSVwX7dBO
1qMIzph+siDfyj1a6ytpQ4kXG69t1k+dbZNtjW76GLjETRrphYkABThKtXtJAoqn
cNE54tx3l/7T2GZ8XtZLsKmDvQuzjAh01o6Vf7GHLkLSBfbMwjoAjmBgJMNtVFj3
VovdjBA7Rs/lcygXsIFDlAtkSnJqZs+RP5jn3T+lj1CnNpc4nOUJc9ogzFzbJgpX
Uh2xkKEKGiN5Rv7ZIpm+J+0Ra6nTtxJCWcF65VAbCTnTEJADpdPDGmMJ9THx8fzh
NcWVuQ6jVvAq1ch0MBVZ3OQryFCoLUG5/pZDJOBN6zTGpMk0/Xe53IuRQ4itwJbF
vS/3U1lfvc6C4pYYtRNCTYvFW7uldNqlb4GWuSQ+7/b3JH+siWintWdF4Rt8CBq0
tGe53hCDQ3FQlKRo36UlstE6pLa0SL+OO2Jnt3Ni6CK1NV3+KC8lngVezaDhQi0Y
zS5q63/BjkvMs/SOCiYzKfWYFMHj46DFiBgx3Bqvh+NhQGZ/pv46yw0xMbxKit9K
NTKof97GM1QWpOGeBPtiifMZgRqinP8fVVYxw5ZWgvkqFNdckXa1CkvkSa7rgD29
6zk1SVs3u0QqJLbFcCKCTogYEE6cedRPuwkQrl/7mug6pwJ8K1nUJIQfHhio9HbR
XyxAakfndqqn0OCBwWNJJBxKjN2ZiRONHpRM2S3zkTX4cXcXTGhn6sOH9xIfAaBf
OihjH+1bkIfeF42N9QHHDmPVjeVWIAySrlfZPkYVXZ9ul0Naac7aD2n6RYB8a6W5
OQtX7/OTRV5b/1w/2YbhnL5s1xqPNn3ulX+BKlT/zHdJFiw+VyoPz3wki0PU8TLl
+rR9WcHO+DeWY4Eo8tV654YMFTgo0eGojjRoUS8ZiUu7jPWSGXl/cxH1SL3sSZXq
w1rFIthgl4F+1QkdXmvn38Q3x5jSYSLLRtKWJxS+OqO1HiZ7f072JYYXpeH4gCjr
LIy/MzMy3ekADJSijq9h38qWblZXis8wWmlK81bJ7alDTmeXtfwQg4DJIq67Rokm
pAkwvVIX3KoU6/zDISe9zekSc9pb99fZM+v79BqKjhBihfJdY6jqzOYxTApy9Moc
b9x3ZE2DG8xd5NRJfPdsUHVfiS/uvnv2rHMfqGZz1Ix1Qh5WPj+5vS4yNMmMrIMF
lnEKv7zD5YZSSI6/b3JpK6LbVQErKyyxWdzYqXek25few6FEViVtEp97SgNGcmPl
xrxl/NiCREVIrrOdFYs4msjjiColH5e1xzTtyKw2ZeRvZIs1I6Mohy25pHI2wIDU
IdofXyxj4TUw4qt8QXfEmTrzwleQ/4hamjtBQ930xnviTRLWft9iTmhoMI3KVe2R
dlZnNFg/h1bNpRT9msO0EMw2niklOgQ8kA6bzozL22YfuDz93gsATRalodmqnSez
PMtSolgU7hhEXponZDTDerZu9j0Erc6YyT4xy/GgxGsOKFq3Z//aY0vxLtpRb6LV
eut1rFKSh89SGfuAdV+fiXOTIvjhwM1gP5j665gnTm5RwaiGBhL4MkjTPiEKz2Tp
vetaDuDDESeyPvWNBtsQNx+LqXsa5IWZ3wwbO+Wynqv8OL9TiP/fcd8Ctjh06C8b
Zh/i2C03kM54bv0xoa0gTm4heL83rDjV7buCwsuzRsEx/2bfTdMyk7DNU2WhaRfU
AISKAeUqXCZ9VKdvQrH4c/8g30uYr52KLgEl4Y0BguhH2WTVuZPL2UwYGNs431t6
fv6NuF117AQUa2paiQm47gzqD2BPvS243GzuzSnROalHpxf1UIiPV/QeYD5ux/a+
PUKeJFBfetWmN6xmjhNZELCY1xT+j/huF9oTBNjE3xcPdC8VAmy17lpVlniADTd0
3ouI24gSmBmAi75BU2B/37p1wvinJBb7TualJjjXJuwhVLYOvMcU+J93+xED5eHw
SuJLv9k5FklJL1YWr2/LadHa7XXL/KDdAe2X2XlkuIKlh4LHQ79d8F04cYY99eQB
Qio1HezuIs+B8zwH6VPvrdbjgaL3rqm0efCH43i6DxwmvpsC0kbRmpGzQa/EzPIH
q/njp3sLdDeBvafHr+XByTAFy+X4VhQSePifbG8l7IPlYMn+8D2Q5vbFUu0x1EtW
tyKBcl2lia6dwYbLuiXt6PWi6WdxwSpkKYKKpFMRIRX08CPEY3byzSOU0obwBlI9
AWkMxaDlZBMsSw+zzV5WsCIXByXPdzJBS+CE4qFt7wtsZSXU/Qz7H+9U4WW6P7LB
IHIU62fRdmFdGP6Uel30o7L1vhC/4rKzl2+RXz69FgUn+wLjHeUYjTNb9/WxHoXK
RKf0bIfcA0vl/sAO4I56YZpCjxse0Zr8YNL0jIhDXt/FUoj2KG1PuSluS3xj80qq
rfdFL/lFoG703zSPiBXcbDhTmYPABjS65Gf0brWC6k+A+EoxIVm6146krRfQ/i3n
0Y6WQBwYcsc0fArll65lLCBNH2RyQ2ffH/JO9jEjvuTtXUatm2Va9Xj4YV1RWjVt
cokI9BFG7hhfFQoMOghJDxZdQA6z0FmVY80oqAcWNyI2fCMX6byRo02gPg/f0Df8
JDmdpuCo7P5FA51NmyI9DgMC113ugLsWP+dIPdl+lIbti6atID8H0ABLtHcbBsyr
5nLMEC8DCkR1TyKcI5zl3ZcGvNIraAjfagGhYr9ZJfY2zgGhEpNQ4Vhu+K1bjiJx
nTNRe14k/3wZscvcBdjlPRLVrcBbyj1kH2YmzekI5+OxG9Cdh2rnEZHVkeIOB73G
LExKXenxVsVseVEJCaKK2KMLyr+ov+TT1psS5ZT2dnIDaO/Ghafj7izKJB/VmJOR
qWg4US0Vjkfi+cEnz+39IC/AOhn+rg8Q69GpH7g94EBOCXxOYiScMhkSCgOYsLVT
lHDOTcd19y611pFZFdm6y9bxGN0ABQz6soPVtCqRjTBrgbyXqdKNxK9pPKl9K1Or
36RTPGyYJCIvgjdMa4wCO5Iw5l1TW/0dPo7sAPxyIXW6HRrmd4BctNxbcbnFZKtM
oZZox0IutFOrRk9tHgY0oIMva2ih3cmbobquR1tjeeCmsw08Ix0RM4Muhtqd1Ofk
o8QUO7TEMsM2Mrj8lJL0f5pG1GjtrZydsYQGm6BRGnARXKNq1DvrZhSgqyEpuzlh
rNbDqM81TcgeaiV8QtyubE7hu4KOOKT5847DsXozsIjWxOPH1RDQFdpVORb2f8AI
Ji/phYhjmMoRiX0JHzQ2HlH3DB6tvv/dl3LMTpCW+/7Ocijq9ZvVQaMTDY3ejudu
8EoYwng1fS3CqEl/IGE7Yoksh0Im0iVbSaIiDxRqAcSvjwAbKZ4HsuCvy4lSluUO
4XjqNhjQmBjWHnrtK+beQT9T97QaEpAODg99op56O9CTRnKV31cfp3Pwq7viQaeO
1hvS1sHUKq3um1b5h8WxBJW4v+bM5qr3lyXcqoNw+PdWdyDRB959zWNZehm0qm14
JEMSp0oBvqWDB1NocK7cfSMFPzq0xxqGaPW0FsM741t1v803+Q6Rk0bzhgPVfRHN
12Zu9VXIJ6PC5p+7rqN6+y3waxcFP127zfTnTKr7qGw2n44PNU4O1JUG4YT2NSgx
RI7V73KR1BwuTJe+wuF0ZeBbduhxNJyQ0KKKJ118ARfUDfjK1DGsk79P3wsdDO8D
QSGm57Q+fLoqmhu9pIJNdphuuj7Vb5iHRTTpkr9muvSkG2RAeaah1hwh7CRwqUm9
UBmvb9/Y+yepLbugq5lDz69MqlaretEPbw/6u/4lCT2PQuTvXRDxEruUUn+njdwh
CFcGWsbsxcOJiObDWnOcHNk0DR4K2pEteINjxmydRAOgSa109PW9JW+K2hJs0bab
JWT64sjSV5MpLMJBgqOxWGN1ojHK66G8hgdVsX+Y2bg=
`protect END_PROTECTED
