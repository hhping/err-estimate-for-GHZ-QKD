`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pU8gwRCRkIpQSPQmcTNK8Hsp2LEXUBjJD1S7IXXOWYxuaWXwx12WiEbCFmHcLKS3
/RaWUQIfEUVNm6crlaRVQEoO6qXFxLBsCZSRj+0FWRuCr7fp1fK59CbL/zBxZFJj
ByHuGT9VzN6hNwxjC/iT7iz6bEr/7jhX/fnfynJ4kJ5m7Dc2MA8sv8qfX6uqXHOv
w4cdMu6Cky2k4O0hxnnSFz9h9TWLkmahO+uNIn/SkI2OhFrUPZJCJD6Xz27JEJPz
Becv7o2bvc5mlEj2SHXDlouzFUiqoK30CFG7uLbWCAT//bCMAkPQM8vro5/VKN+B
ylA+UeaITdk0qjKNAk7aeGEqUuWIEvqBNYr0GEylElMdkA1TDFLAiUpXSTVvitzc
yUXeZXmyS8vVxPer4EI69wD4bu6vbxh+Kcb7VD8GbWhf4ZxxOg3qzgugUi9TU8BH
eyiJlywabNpFe/b7ARuMlNbvmhb0ld9j5spbLs2hK2ouB+diyFQbNIRQEnDQq9Nq
+XCj3CGOsA+dEYNMr4RHaY6cEHWGu8LIaWW1dYZwaAflJVTJbwqGA/S8FB95fyeD
cqU4Pny0Fjz5wCNH4aPlxBODYyQT8qs1exl/o/Ogw0r5JhBiKeI4tcrBs2dfb17S
N9qQoXbvWl/zjUkHdtYWXwOMlpzjkKQAeQqpvaMM+z10mqVl3oprLhcgc+v3La1x
k72DI2Uu6+8d3rwEAh5Q2AWD9Od/RPBkCGQYPmi16Cl0SszAuRu4wWGon5gIObs8
l9RLyGLvCSdoQO2CymS+MMcixQGaSDWUFdddLd7aIv0FLsb64pJ1JymZP2FRziok
NzukiiraqZ9WDHY+6w4ctPOcZYkMYJNRfxXMzyGR1O/s3eUdxlNTzIwwyTqOnoD/
sfP2tE43lcfAaNoNMi8wJgFoh0YedEWdLyJxF5vk4yYhqTrQ7q2aRm3nzBe2abTw
6e+v9KfoYGskvjdA6eE1e5d9ib5vlFszHLiaZePoixlKGoM4T6CBMPImGQYFOAYv
uXi/0uJNkNp6XgBYp+HpcioqOZhEFsxGU1JxC8zVKGcLddxu/Y7hTEFUFzIZ7/0G
CDfgPz30vCrcImAxHGSTAPCdrdPI2pB/OQHiJDgAD3uvDJY5oypq/glTNxrrhbhf
Igh5P1WbMuzfp9rIBux5WVdtHF8g/onyIWLsWOFt0SgEjFOevibqJNb8I93/eyyt
CKvKgTE1TiVKNxbxzxVkNyVfqMH/2lDMWDtGb9zHANgWqii6/znNoi7bh/rS575Q
uOhCGgfJkAp33LtX1BfyISugP+7CGMIO6li4y1uXK5zQNyjQETfKAPRDh5yTxh9z
9WUV/13pxjdrXVcSuV6PmxLZokdmvJAGJrRQGz4T+2IcC64fEd71FaAKKl+PYbK4
bLdJgYKAA1G9O5BLbhhbr+2hQ+H+uhMVyThALbMk4tLFe10k5tBGQhycqxZNgJZF
I2djghXMTv96CyioImNftdxs7uJPt02W24lo23L72hw3s+w3URpqwfL6hKLZzz3i
D9VvsWXSu1HJ9kQSh7HQZ7swWb9Mc9GQIIGauIYvoSpmXy5Vl54yAgOFzrpUIMSO
l0kxx6iWS8x0ss5SKYDZFX5X0FalQ+SvP6CI/WJONugv1pDoqSpjxG6ug4P5v6hM
YBT/iVsxNgJYvnH8b6umvA1d9Ob4pjFNdlftHmfp5rA4Fxvej5QDJaiqQeF2Fpub
dYzsAQfB2wBP1cj//p1XiGjf5WQhIoHP/AYGU+5J9vdxY2GcBEuRKUFgQaldo7xX
ra0l/F1qfX+WyveTziWH3dUyGWaW7ET6DKQNcKeJLMAfFDk8BMdOxnEqnOjF9tnO
DuUY0IGjS/xuGIepmkiq0AWjIkjMZuNaSj9PUg+PVTz3Q22nOCLlB4DhdmI1GhEJ
0KcrqiLKWuH6haOWgrkHLChtMlDblvfDVzOBSc7cyTyClE4wKXBEl+5K4tR6p6bL
MbfltEr86zbNxTuTEYqd4A56SpceNnnGBbEkQX6yhWsibmSMM2KoRXFGC5UBmSrT
48ZEZO8CmokWkJanpS6js/oPQnNYoCxLMh6S6Y0lNt1xl32VclHJAj2hdAtt6+48
YeS4VoSVJAtDggsmRVECL8lT3b0IhOx6PpQbhU6z9FwNzX3FosAmPxZ8sXBKxKOU
SoM8Hz2W03iMdWuuwNPR4byIjkqjqkADwUStdguLmcHsrdpYZ9tx/4Ed44/QAcdc
orgOJ6I6/Tlslo3Ye3uqDnkI1ojTDfZQ6fF32sewG4lH+z1ffbR4izM99aPwDVs/
EZrBtO/nk3b6SMslmSeBXTpU83tHNrquAS8PcxHhd5k6VQy5HCP04BKzYk0/5pgI
jltO8n3oTsZpsQQyWHBIW3d+3W7GeRZwJLSJ0b5aq9VRCGuIMXA8XL5b+2KwMEq4
n/tCizrAYmes9pk6zUZ7ye0KG9lLuqT0fVy6jAv5QH8FlFMTgxwyC6gb7JfC6Ucv
dUSbtPnwlEs5Zp07LQyJC1sQ6mTBb6EoXadILS4PMVkJpBiqdOa47dQ2AfqqubFe
rZ8lQ7qEpcB/Ic3S7k4Lu1YArIhl/UoPdHI4beJQd80YwJLUHFXDWsXYgCP0lT3t
vBQfKT8/dZ6LtuCVWH5O6x7v4FZkL2LIznl7wJfmLt/U3zmRgWeA6RPVKhfxlFsl
BmhPIYOnUcMcT9fXNdA0WK5dPhHNdsVxVgmK8Q7gip80F6UgqhdodUlJdXh35Mkm
TedGllGB/S3Bjkz3H3jV2w5ucgxl+fEqcrII9OLvrs2//2y9FXJIHwmqSP5XPzbp
K0DkdtDHc0JXSOdadAjE++mjKdIhhJD6HIhV9ZDREywzzW5tECwx4C3ju5ILUaE6
YZuSD+C9padKjyQ5Les9OXqf8CTkj4ieve45ZbIbo2TynBOKtk4M5+H7BDDJWjro
aCnBtgDm3dybDuiOrPIPBkj8vmQmiBIytd8Pq/Hr6YYVNOJ8l1ZCAATTivS9/QmC
n/irj4EKOagQHd7FgZiQzPHk+ku5kvKXE0arEPO0aqstQZyagTZXpfnicLyXbhJ1
KzCjl+WTljLaBE2d0v/8vevDOqUrU6tyzoCvtVnWdZiQ3+pvqCkCuKDZyOPfkiid
wEEJZtd/1hEkzTTaDMj0tDVKx8BOa1lMO0Cdg6Pml2DB8g0D3usq/bpuP4TTGKgv
JVifK2xmpJ/+FLvtrl0DHnjfQz/cykARqj6gQLgecbhyn5GamHexWOIy+fswOoxw
YlU88JiC7fDuGvOvXYdw5mpMIBctTEYB6NHUbxB43Vjl7maYo8YNiXs+hgM4X1tC
F25IT5BdL9msBHs+TvHlB6YqUSDG+raJBSXmtRiUNbKkpr/PHHK3vjjQavBO3tOp
HKGKg7UWdMr7mrVaPuT2afVu+A5jH2LO1NWV4BTooS8CsxdDKU9ZWfMJcuNkGcgM
V64UY7EV1h7guzySuhDdOrQwGnci90PmEuCI2x8czCvjnTb391XkbaRxqUtv1teL
P5GUn3S9sxswlk/Ed3wkhK/7J0Gh2udK6JyPxylHLyOYNZYnYwE1JKZgZCa16V3J
w5+7fQ2xgc4Qo5j2x6zuB8FjLA9hD+J1wAoaOoMxAq80JR3uSyb4tCkzkD633jxL
d6T0ny5plLInFWGeljW0CnHO9wBItUEi/7ojYRDCg6543LFz6ii0skfT3VltMU+z
4mPjW8DBUZKgdQeWfXUdPhGP44S1BLCk6B2Jx5PxUVRgLd4+WxKThfMadB8oOXmX
jlBZoOnppUsC8Uf/qpHh1vJefekqpL/JBckf+GzLNa3fmMdyXogF0WzithiHM05m
+UZHqXmQ8WVO/vTESPI67csNCdin8Nl7orj2uMW3t6c/EtyXADY9Lrcntk9Wjj1/
Jcf9fBCOXWcPBjYDZh+95bG8oYTlMW1kEVuWKRZmpi+H9t3kLlIeF689TeuIo2x1
mjoO3fClUt5ygSlscKET6LvxWGhKBbqJsV2xfKpxZHauMv0Tp6204ueqVtfAhtRU
H0qmjwuKr/mwhcflOZ3L37vY9BVvD2PsKyQHCCDWUnhtl6CTjIRWwMHQXe43kge7
8n6mRNYsoZuNvXHSOiTMGDy9aMDX/XjW6ZVz7Rc8E3Xyi/3oOhr1cUeNTbFpgkYd
t5s5KWD4ntEGb/jRGgSqS3ss7O1cBgEblMXY0L/6blrhj7jrPcjsRr9HtEu6Ni2c
CY8jxkz2XsbDr8xSvZF7EfJpHNsC7guUHOJ98AduNpJjn8QgqUG8/4zGbvhNOIwk
CkHZoDaV/V1DaGQncn04MOFuzxcRZzNZ+wAIgk62gFbK+ZoYHxqXYBQDoF/Wb+Mk
bgOJyruZWUUil8+hbWAhCX/bft065UkdeceGgWwALmTYvZIB2syVa+r47I0g0xH5
V/W4llLiTsRiDbtmztuNrHZPKOiAr84dpJIHqm+M+NzaUE+5ASDKyvhJBBtx971q
jKRN49ZkfJtwAqZm48UsAEjXDYJKXY4tbVP2uocnrXIxyUFNunHX/CyTxbxiqepm
Fg88d0y8pVYNf1jvp2p6t0mQDyelGt93xMkaJ1hMes3Tqus2k/bj4KuPCDukVt8Z
yVIiG0voCKT78bIxcdcesqkrsa4E4tQtMqelbGvGiBRnCV+84m8HyzgzPuhiADEE
LfV1yBVgjfIh8DbSPDqZvivRgCsD3vWAzWAl1QaiWeRrW90IgjZsfM43LVCZeRDc
ayf+/37yFTN/K+qYlQtPzsn4jluXb8kvjZRblqObnbC5Dk4CIOXAw4yHJpTi5YK0
IHTQdKZ+abeoVPEjuqJZG62GU+zdEccw+8InhWG6W5ogl9ndDIljCvy34posOb0W
vDGXiXrFE1aahUlWZZZ86jWSb9ZLaZmQt8JZzPQUdB+ZW+yt+q/aXrD0dBgODfri
irY/Tml2ox8ChU8y/kYXcqZiCnYw5eyd/lmxtb0hcT4DEim+V/w9ctB7Lu6K11p+
rEeCnK8IxstbNjS91qZeQi0adMFDFThd34NHRA34OS5Ypn9gPDpqZP1lXC5zodn7
ehgh3dVk+RO2EV4/sEm76xzUOm3i7NZ9mGLeAP6yUnfAhVSuCn+7fpjBa+tO+X/c
G6BygunU5P+4xUfJEC+ssvVaGFJCKjARspVBMrNZjEqE3gYwhMLg4b7JJ+e4l3uc
0zXzgA3td9Yy4uImcru77+Yid9RSn73CLgVMQZRmr2s9aozlR8HvwXKj+Vy7t8P/
6jFzO+lzZmaT6oN5JLFUN/XjdNY4evbRtIHjYl21rg5P61KXO9vimxKlTgoOMZp1
ku050TVHZrt6/6kxd8YTs9LtjALMOqRBLIKJiLwUVHudg4OTCn98JiaO89fg78J6
BKwPzvQm9qOW5qfbh8xtcwGwnUC2nHeNZNTx01OfOa6nbgkeqrQ6oF3XDxkYOJde
nHzkJpO0ZXXGAtjDJUEPj9whu3gk6GvzyJbe6G+QyIgU+RjS9nCUYM3b9WueFpxE
PbmrJ2CljaVgz6fdGvhnR3TqC6xJKAifLvaGI6ch7wDbo3pVH+8Xf+gG1zKo9ApF
KJ8Kl+wkTNWnUlFDlIORzuCFUqMNYM48QMDhqVvL7vbHW0qotdCfjmAHTTvn7tpM
rjJoeh3ATyxAQHEPhfFGsskOnCZpf0SJf+CbGmtKxQ0RkjNERh4yQ/P+/oP3RSgd
8TD3TDy1/1Z/TlpiVP8cLh43IQZ9lppiyAZwrpBzUHjESOaqoCNFtxv3V0iAEzE6
sUeAUKhOj57+iFjYQGbeafi0tC0Y3O7sApMQKrs81P75ywNiUfmf/2E8MkI41LMm
vYYnMRu7nsGcpPcZzfiTWl7XS6CVr0cxZbsJRlKky0S7prsxvYPoTXE7pxKWj8JU
l2CFqKMKoPs7sosqd1cpB3wJN9fKvSxNDK0Qnn9wROOV0psy3SgL99aYzXy8cgQj
5fEFoe3yQLkkHyq6cEI/ja9BmiwPX6Y7NIi8JDHAVEExczHcBf1wCCTq4v3kqRXj
THnO4jJuUx2ylNzHWnnFSXe/7oS7dQ74J6ctYGfbY2aN+ZIXxlQ8SHJvl2GIwxIT
lkyqX9QrSEV42bjqarZO4YYRsWYQtUhQySgoyB593oQEqSuHrA7s6gEQMYDxbawD
V0TY9L9K6Vd/sTA18zliFSvGBbkFrZKvJtt7kSudFLLNFHjVKLRnznu0wsV4KjWm
9BYE/UvlRgzYY7dV63yRW5Sf2O+QdyB6Xa71KcGsXUnITH3Vc7ldUv4lbJ5xqh/u
ia7e2zHVtv/SJbh09CLwo7tkIqmwmED1xmq5i9bG5V3S1LUakT8671MifOM4wxtb
xpcZxtOP6vl6HVryyGRwSFlnowzrXeB/M4TaBrXJthtj89kZoH0PLiGmpmyZcyO3
7T/O1CEMuATiGVSl3PIX7guPAKhCqUTpRrzXQvTJW7o3DowOaXKK56qJHvpiiqOD
GKSCkPYc+/eWAJmTMWrlngTSD01lLQ4Gnfrb6QQO5uRFdVQ5k3aGywQgmcFZz83/
G7sXGVZSdjtHNQZ5Xk4BYJ6SZ3oCKv1Lwtvg3ifMj90V/piT4R2D9wYsPVkUQ1/g
vyuFAyilpHL/CcwPePFfL4wfsgCdKYWVsVoShDp+VL+BZQQbWzBGyqljdz3QjmnD
vwHFsaq903qb+Cg3NXrE4Rcem8tu/TAS6nu4merAxA5tgyc22lYhD/RUDFNb/e/6
5cbbU1k9I4CncnPxm5H5wz+MIQ6Y6m7SfJzUTahOHOyRxu1r+k23aMeJkqmdLln+
OG/sWUa3naE2/HalBtAYe1XPVYEGvRAUEjIHsFUjIqM8pPmQjzLAc3qrBEAf7WQ0
PgSfi0KyLDM6mhWs9W4v3lUcLeChkTXlaTwAC5hRL7gqN6ymJmw49w3HgkMXU+0t
Ksvc1OG/ptZ/500wNyWAQrQjXWFQ7zxOqXl3RHwC6td2wGLnn+ThShFPhbDeSjtw
jvuvbfjKqwlia+2Hx1fqXUgsN+pPHEKAb6seF38WAEys/skxYlcCGPg9b78LNjnR
PHrj2WM3oBVsIA/qR6Ej2LxjLSpFvbAzu8cUeAsZLF45qhyf4ytXYRmS3vdF2zuN
nZG/B2EsQQrdj3wqMmgv6VGYdYeod+Gunq/77SqYT8/xiuctsYV5mik1UJaXqEzz
1Le91VYMJQKv2gdZVjhjmFWIYN/SdYjFSufY1HZKhotfCWyKUUZsq1JiP13Tao8V
/oxRckwAwJNjESdakmbSNuHa7X4JRG49xk2gUad+wf2NzQwo4M6l4spVWkVaj7Uw
Z0tHNKmza0NoYjaYeXJRBo3dRVNswm/iGYt5NKzWGlH60T8nCnatlH1HlRDIJz/r
0D7oM6JKcZ9kbnF14RfnN3eOlx+IGV0hjeewJGIyNCa92LhiL/AJgrwNQwtLn6tH
meUrg/0QH/RSKxPzaiX9r5Mtiu+fQ8uXTcOsKOhnDD3p7OKSFsU42Uw3EdwtUdpP
LrkX1ix1UJuwp9x/UuIZvXLLRsMRalu4kZj1ddE3zG6xmmTt37M5QDXbD9dvExsQ
OLMXS2RJPTkld0TQljeaclR84w6m7RzyUxtzG1av2u/jToFLO0E2pI6egbw3jOvT
t5oP0zrZjJZJXKnXlL5eZLTvJPvx5gKb9zvCfCI6/5H5Y/qjayVxIX4oGObCfM5G
`protect END_PROTECTED
