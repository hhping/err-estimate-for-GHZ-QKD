`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdp0Lgfm0VAVAorQc9MyBW7W3gBoUneuqWY6vWXsXZ4ZqWz4SizFl9ql6rw8JcpG
jNI+yPqz4aJvrGgNnnqFoq0JV+sIaKLd6Ycl2g7CT91kI96ZRVAZkVrR86LXx9ID
kDvyEzSmQboODqcT+6a+4LoXSDvJrFzQxZBsQ2Bkjf/2JXAGMS6A7DNf+Rl6YywW
ibZJOIiSYNm4ros0o/Lx3NxfCaJvkf+2FRBBWHMuXhiLZpUdWN6eC75dLkOYxq8L
w/zIUr9KVqVYWAT6w2tyRflEITOMa4dobigaudtGqT82VUUdE8V11m5XzW/698hI
fg570+3ToQAMKIIb8oBhyEAcg/1Dl/8052Z5Yr82ZqgT47Bmm9cemUHkl49pa99s
lukiSo7VURwwJJM37YnPYn9kajuPOQcmlAVfLMtgpT6FeqGo+3E0m+qEaPB2FWdk
R3hnHo06roRMGZAkGsXKgIwqNZpqguncgccEWpRcj+iyPC2+/xFQFu0N4wj2oqTr
13i3a2rTBXit2CtX6GGT1hbzx+0utau2X4dogml9o6djoqpmZa13dMSQAxBpf+VS
WR8CwqOYNZqN7hgqAL7/A6rPkICqaoqEKGmOUD/UGEzH0vMz7ZKkXjNSer+2L+oT
J5uKj0GohiUai8fSqfi96OCwuY6t7ZeD8wH2OGFE+/UHXx4on+g9loHBqXM0g5QD
HOkWPMEpgU/w1iK8OIV1J5oDa4hfFyFhm6tlMLHAMCPjfPxlXOnuk2UL/zgBzdRl
H8sIpVOjwraozKWjxTbtojWIyij89hoM5CY+kLdfTKnoZbVsWo4jbM2EkwmB9DsX
`protect END_PROTECTED
