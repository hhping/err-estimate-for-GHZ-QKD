`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jn0kh0BamO/s6YdhE6z/Dae44UO7d8WwQx0KhBGXdU3yLbW6E77jrBXwMxx5C90u
LIJCrI3g3TLgOaBOdAO8jdZ9+VeRFQvqDx6BAK6yNgw86d8FYFwI4OqaIwezTYbs
O5Vn4tMePv79Kgu8mO4EzXvdTDbR9dxQAlLfL5VETk5Hp8LqsxFgM/SnChdhPchD
lQypaMS5Ha1Lzo0Tph5ffOkwb5SoMQwWqqFS1i1mLP0dMoQfQyk3p41+fvAuYxHs
B7yYjXc1TL77H2sm9F/ICe8O1wKtctK7BIZiXgkGs2bmtU7Sakk2zH7Rr+OW35a+
CVkHsfy+JtyFJu3Eq7bh/1MXQnOgMyfgjlYeskKLBf7UGEy0oofStwbkjg+44737
x7k3DtAFLAxl1nUQImdKVd6khTPEokWX86l95+0F0x0ONxV//eb2O9N0nlnRU/0Z
t8WH5ECYJ3Pp5tLRGdzjy2JWHzH5IsHFXoaFvInqYFyHYmqgIC1HUj3qnqbBtJa0
k3tPnWivKiaC0lL2bex9MWSH5pgAjHwto+Q/Xp/yFSy1k9OnvIyxNlMBBenirXlV
/p+kwbNZaOL/GNojL1QqhT0KFA3er1i344nIvbhO1ihpJKPeuvxaJZqgh6PAzI++
ml8S0donfCQWSwHYe6ES10az89L3zaHsjN4ynouOMBSr2Hdpxt9fVmcSW1BgRFEd
VrYX/i330bsBqOmUijAD3FzGAmcTpN8uD+YcSC48RxR6menAJpmnRpzBEXi26EIR
jWHzzJ5WFvOVEB/Lpulo4rfnu9ekxDmZgUCF5BBuCFwDt8nDtic01pZbt2pehuwp
XWPyh3Bx43WsUgBIwJNpar4dBg6P7sS7U+NUktdKn9nD2z+8xUpNd33ec4lOaN82
6Ceq3yymS9z6HQOTPzo3Mx7dD2aATB1g3iMEMn1Yk+1V65rOKZ1OHnhl9PuGISK4
Zw0qLXNeu9BZLb/LUyqb/yZtMmZAkh9DLCPORenO2W7gBvNLLt1tFp2NoFm+zEFT
98kUc3kFri5C06kxdCmedy/N5dOXfYn7p7ePhsEAZ6Kr47FVDYTSbFPNcAZEwaLm
IoHiQ7sRZuQep+t35IqKrCp6V4pSW3v/SKjYf3QqY367jb+nnwKVjXfXYTGu2sgZ
nKUWazdPusNnDs0iuh9vbCKtO5THg2IHKznaGTM9HtgsMmwg35wLdrsAelgHjl/t
OuvaD6Vb3LqeR+SgvGMdEc8DjAljLefD1Un1CW00YT+SUCu8YD/ci+dj3zXdUtjX
IVbNPGfJ9RZ/0NU4NiQvoM+ETZhX5REXev+hvaOeUkevi0fgveMHiblTsGO50vHW
crrX9QvmvJHPa/FTq7M7nAQfDDwWAt6kNsDCi7lp2OBUtyXmprZKKO4Bexvi7G+q
h1PdQt5NVkGS60/m0qWclbclpXjUGCT13Qtlvj7qmjTmi/BqtUFlvxNejXhja9kw
peJpWQziml3g9B5Hh6B4/A2lU4YsxgJPxJnlgDmpDtaMua/IPcUJn08KPKJ4b6Cb
HNasgdKoC08cWwJb+6dotcT5gJdsSI9kB8yjFzzYlcdW5E/nP55KpMKwRuYYotRI
pPh3MzZaERlX+yWuTck0I85+svg0coi5tyO/WXjsuUaq3z9LHlVQbpP98W4MAmqy
VDxeNBhm/fX4Lh5V6lh0bvFXJXWiKSGG+hG1cBc3ha9Mna3PbI3RD0SB4nEgMeb1
HvSnr6PCeMHW7ZSE0ZZt8Kay7EVg7TK2OnTgej1OJLs00Qqo6coJUZfqBwMo8nMp
h4I26iCKlwSoJdpLStO0sWGf3KusEc5HcWDk6J+zqS4iw1qUB56962yEikCXZKj0
v2ElsqjKbIauMBLTGB8pY61gL9L2L2zZAZEBzlLxlhk/ewfIrdfZchLxY4T5k0MT
vLFbL0IjA3P1mh7y72i4AYkA4yAsDHeEFSHww58zjomibhIwz8UMj+Laufa+gsMi
ypqpqpJwbTX1sExeygCPQ7gJsmn0hM30XbdOikx/dS6RHZlsZ1ND7HjTFEfhfioN
O1iUQP3juSRjCiocl3Cwo2FvI9rVDdDz2vmNplRhGHVWmALr15KzCntEMqx1oT6I
XP9qc4rV7a5kcZcFK7dRaAGy/JUZngbKgcKa7Wv/PTfP+BUYUzhAfjziJOfi8wmR
qydBl8btaEZQ+bcbWTpdSxgVDsHk5vaESXFoXCGf1is0XEWkLtTtlcj4cJuFSV69
uQKNZTuHdwA7cnkdYTRVjtvxQZxR1B2hjoCefYMqMOFrPdcJRU0VIR+h2LtnTGyj
+3RJK0dUZXqUEiiLT7Peuc38BSFOXqhggqGCxWD0/yXSjXygteYcc7xpLF4Dc5S0
L6NHBVi+FoZ2o9vlkIeSC+l6ofJC8qrEe9MkrcxD/IdsobatxVdfHcZZ9ozonzgb
cHiZeMuoUU7K1Ja17iMgdfs/7Vjithod3LVlS1wzO0qZqBKg3AqhVebz4bnlJtrK
lpuLE6zImVyBudDez8OZOF9H2OoS67zRq8xTdufsJUwYH1KRY42IKjtgPvakCLdN
xTBHQ8vjzXQdw7zB26VgRlTc88esZPrwZ6SxatSil/ihtDT1a1NJGFQdRBOrlSup
xbjEdVDuHtC23w4vi1w0ipcGqY7oXWdu4WJtFjgLYQU4ZnY0B2KdaVU/rqhHaSC+
ApUuCej5Cut20HPQa8dP4MB0/oE7LlDr38oGSwVrRLfMkelqMMcaYS4DvqJQJPkF
`protect END_PROTECTED
