`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jo/7JuZLixuSuU5TXlsDX8mwQwR7bcEcQ0hmv0yt+H/CwaqOQYQHJqZF43Qoxf7Z
Kyclj3Sw6TkvWGkdJ351nwr8AwU7JYsMneI1b/CQLxSlL0XGwbzvSADSzTYNFti2
3j8rsMuBF45fqmVaNLpSEjxVZPEXAEd6areWvE18bc7vuezqAztI5UHyZms3AqRO
Za35ruFwM25ojMoJWUVPC3LxLgx0lkNLjyamMjodnUfAs0QQwbu9q10JB5xb5Vea
I5QETEt3nGGdfGPK4vSdqy4I/bi5igLIoEIFmNzvHUOlW0SSPpJxCZNMqwa9ed9M
3a8GWmtoDQ9LlbrMHkdGfrhj83ra75B4szxkWlJCGzhej1dNOybtfwurDLwlBxmE
0GCfxczi4WLwOHX8pWAlgA87+vxXYaxwp4f/X5cZrwwpX/uyHUBP1nB25kfCvy26
+q/y9e7dHzsHe2VIXq/aVMYtkfmBeTsX5EL4tjheeVzPj6U/7mCBolmjAyogwzUM
5ENpeXJw7pcTba1xaEePSlMssGc0YNDaScADlpClN0z4o55nZYAa+yKBdKU+BSm2
jiN5VbkUVrvRt5OGf5O8MpCqQwYqX4oUaOd3iO9M0B/RFcUs71hi9ISxgx3ISW2f
hlcTbsMqR4GkKrAI8Az0isyI+eYz6T9+4lGsVW4d2XtM1izdLR1W4ZDz0MyW6g6k
gBrNlHeYMz6JdEwb3XI3E1k5A5YISwM29B77blBZgUHITDL478j6j+cFEGSuDhj+
gmf7Cqg7QaoclQdTGRGeIODYZRTLcwxMPTdJdYT/ngb+f25QhWE/nkwSDyxuj+1Y
F4DTeF5UA9OtyqBxtM1QCoiebXt4HWTrdkcpPdPGA7vuMDtEEq0obRJdGSsgW//V
4xqyDlc2OVjZH81lBF0qjsbVxhAkC4o88g0wgShjPnApQbcA66oVYRSy1Nu/hXzK
ah12WF8NmlB+UhYEWuSDJd1FM5eDF6adGGzkUzTkMT3wyzY7MqjRsXHo8PA523f4
mn45gFTZoivxnUUMZO45v5ZGIKNujgFuIdRewRxYVrMW+0q5yC2hyTJCjvdkxUTm
DYdMyLn/AqmmgWiJfE/6vfPcnXYFENTfgcfAKmzjjtw/cC4a0i7f1bEZZyAge3aW
sGvwtN0ptBmQciIyeSOcJ1lYqTQCXaz+LK3wm/qTNngSUsMB22yjZTdzpIn7gRXh
AEFMTh2doIpUHAh5c9i47iu5W5g02uBRw2EQctGP51oco9Ua9S8Wa7+7pRhgYP66
DpeSkDLX2uRVhiATKEIDVKShZFn5BkJjfubSoowLNX69u0/0tHjZaMCR7dczzPNV
tAz2KGiLy+rHCOXoUTyzgdXp2gF5EfdgVVvcO3F+rjku72osduXJlDzjkCcu8u4X
YU/PV+Cfs0EiCKDPEj6PYZ3/QnkXb90HsnnejoTuOHdxJlh2p7EHAtJfyhyHupy7
+8qvUGH4Ar5CS1exrnb5TflegaW1+adT4/DUHwIKXdbOSPgb9JQ0onVmaxCFqvOM
SLG32/kx9dlu9pspFW+9mdy5/wcZh+/H9llHAYYJ+auqFQac9kxgrgZ3bvlOYYr1
AlSMdu+lpBtnAUs5JHJawUQssMrQ91NigOXilPT/CjZhPebn4A+o392ZUyt19f3N
fE/b92Ip1ZWmOrx2ule/QtN5il2W7UVMtH9KRMhZh/bhEHjvATcTjT9ljlFjfhVi
BP4wXd8yi5eIOTh7CFle1Zn3Fy3V3WR/+C4nP8YzgKK8G7bG2VEslRgGPIZoaMd1
Ff08XK9+CUpIp7+6pfjVehc5zCP/1GLsaOkerQjXqqYDMs0erOutU4jOdTo0IL5b
bynQLg+W2sHIjqr8Ae7MS2TOLEL2awCbYNznubU5Y6Qllx9r5X8mfA6sCeaBZEVx
`protect END_PROTECTED
