`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xseRSrIMv6GWe5Ypj44KI/YHTErPqiJDOzVsHuL5j5xgJd2gbO576gBR2Y/pUOG3
t+0OobKheY2TlzwDFjXEewGRZMdCKNYiITnkepf3FDw5gQv1YnoyQvjOD/JJFAhV
3EvRTyVE5LyAAt/MLEnOt/1sEfkWlmM3FfQx5JZqueTADeUMPJ7ezw+iPryxGFUS
m8/iGdlOjAwr3Ze5EQg4GqDETeM1KtPLvzdIKhQQDUgwcHqFXHzuK49WkHTX85tW
fj4O+Bhdchz0osmDvSTvs3Dj5KEclMMo8eByCPgcpyoqxMJ01ZC98EfwzPFAQde0
ablt5ZBHUSWl1q50ohvTMVWzLO64CSKM+3FnuzpHmtZACW+FkNlkWJ9rO97JEqul
hU2XfFSemhosTWFzGPSbjw3Nyg9zIonzqyfmntu4XY/2mKKHwiwTQ12VrPJrMR5q
g1rEgnqMLz7cxeBV4M7dONrhirJxe9En96JhzccA25sgqAMqKKXCwUzyXvVC8bFW
38h5UCcCNRn568tgsE9hykBT+OFC3dZBoeQ9SzrUOTPCVm7+L2shqO2/zI2OJ9Ro
BY3XWsKXG7yfB6ziE8a9Znk8jToJe/POuJMVWxEtUiC8bHy0A28F48ZM7QqqikS1
sqt6A5XtR2a9wcYwBsjRDzIA3n/3mEcYg25LkKHdYwyiSzYOhWKTXyRGv4Gh2YyM
HuPN41xMsdMUxGgjm861hsFdu/3lEld/rXJY4BRvK0rARAQ1Hs6gUHbVSD+GjTFA
+uOod9VhvLuK4dfE6z9M3f0h9isFOuid3uHd58J9qztjmgtSegNB2H/joWUdYmxt
6mFMwzQoa43HTrgk6quKluJQTWPywN41qM5kbAsnzAmjTIEIXkStHwEep9x7IJtw
YyNPavwQZkMj9QWXI6cdYmSqqForeksJzXxaXeuXkatlj46G9dPWETPuCutI7kkU
9BJVX2abfMPhlV0imfkgZBofZp++g7kh2GWdBp1oAIHx7ugGz3KXA0HS135ccFUW
sgcRJLJ5DWQn0R06A8V6du5yImw3t2jysqiPxvtjZQ8=
`protect END_PROTECTED
