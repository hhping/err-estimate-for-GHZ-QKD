`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/bhnvVI2/8QrX8XT74V971EApsyKStaeZOYqBt0SCfI5aOjizgiAf5Zb0RsloJG
P+mwfy6/iQrjHkSpUkVrWrCINK5bwDgpWR3Tv5u+jdrlH0YXDz0sIbR0Wqj45rU0
cf8u/yGK8QKTYr/177G0ak1hXNvESLshAQSmXyHsvAYtYRdJdBi7GFLepdou68+L
3H33Y0nXCQWM7+A7MLciwi9x5HluUPlRcGnZbQhFSgNOlcFQZ6t0tLQ8dJYMwLTa
IHJkRJpUlYHSw0Zc3hR+yHrn/qzoNVR4xdkqN/I0Gp9Mz87wK2uiYvCadbDkq+r6
xZuVHZgl1UnVNt6Ji+4y//HegIQbeJkUwxUoI7el+JQ0pJzCMdNo4ZBVZJbSfRHy
BIlp6OH6DcotTG7958brfLzzaW253p2rb6/GOpFypqtj/VuAJ15LgaZz4MclNMN+
VBUcOTJ58C73475nBPzARsVRRJr4jHdNLOvCtdYOKmYpsjOYTVj8qsYhDz/f0LWU
Q5SRDC+dGVnvQwXwix4EiKTHZu6onTixEaA71JKknnleEjsqGgPT5fJsK2+o1NRi
bSe5MR43GmNozqLnlr4vntSjf45wNYG5cgvwEPXwF498CjA80ACivhOKPrv3t+Io
Sxc0vZ0+YPPVtKrctwhUDtAN/0y1ZCj08WVYngfrJK6EvC6GFsHelabIsoPfEZoC
wUiZWC7ZqvwwCv8IZtt26qygxMSAjaFGfgVrKlBOEY8fd47u+CWhzAUSygOo3zOj
WI5/3ELQDee28BAFnaAuVQ/qBlFqTN4ep318WRzkHeMzE9GPBToXSpjgUCiv1kvO
yrG2yoL6KxUDm/ss1R8jplKmh6JwY8TB841zTn3DjBV6O7xk3wTJ1lPplhWVAYKA
Isy2DMOf69ZVUc+UKmTYGgdtiacsjBUjlWe9yKrmSCLlo8HucPsWAH5Ys5HF8a0x
3GDh/YB6U9zF9ZnomxVG6FmgriNeCD0VEeRNSFTNK2XkS6h9F3LdZ7woZ3x2e3hJ
R/BYgaitZ9m70FS90PkA+Nw0O+ozuwou8J48lAahPvkADO42nh9t5P4/OcrU5z8J
57Dc88lorlxlaev7kGe2+faWMfTz1dJvSig5Uq5iacKey5dSEtEOz4LiJgKxNPC9
RzPIyiOJHDzQFyUyTLFcD5KtohYzRIL4cXonVqDO1oL0bXPOLlrxPKtadSDckhx6
6sP037U174kB5nTuFi+TiHdTnC8NUdlGCKM8zju5gDTzMaR9lmHNoFZ0cjWGE+iG
sYUV1bnc80wQYcel/4kqOANlTXz9JLCf0g0dK38GNl1Nwt7pKJ/t1I0CSB/mSzhA
qxQUrs0U1pIgGhEIn6hbKf8beHY/EQ8euPTnbYd3v2TaHyr8M/1XfH/mF0r4eRDg
u7W+BQKSBZyQAEyAGE96LFC+k5tVTD6mFbhJjp5Z4WbgZHjxxJ3aiosfOujfps2k
i+3Wn/0BzzfgI6djCBrRXJLaJ10h/uNECwbyk3fMzCAjllIvDRelbGeejGiZ0eYY
2c/GwZ7IhILpH2hA9YBEpPDCwbT32ZxdbmAYbgsniyuK8aV0ijfHEgvPp4JGC/QP
mPlC+ngTtl+nBm39GoI4yia/Xjo02DJ72OFpWWrHvXXnCANLQMZTdNT3R8qeUVfE
1Zgt+mgtqCD76GG9gUQGbCIaEuPAJ+HyNuLgE+mxRFsvsU1cMG2Pbh+1kz5oIO+K
BhgkTDT3tH/RldiYQT2v549wDnJXmVjRBs5+u7uEJk6BCKNAEoTxtE/3xIkSnN9s
o8oAqjUq+1ZcPprkjiFWcl3vcUKzdAzARxNNKrWeqbmWRYb6FqJrRSpI8tZNLHN5
C0RE6Ky7Kz07w6LrHBidVXUmgAwrRxp6p8gnnLwhJP9BK9jvm3BHDrYwYA5mXx3p
1cNiDLGUph36SPPaMn9Vwisoo7LPuGaFxAJY9nAb11s4jTU6tHh9DGrvdkQfXBuo
O7RzjcgsvHyQa6iDzP+hL0+IpjMOAcksth1eridZlClU7mL90nD8KxA9ovxD9mPN
xg7s4GMUcH7QeDVq0KczhIGD0erknkIDpR7tHIRfaoVstpwtyzRgVNQZ3jA52Wz9
iR5RFQJPrbKH4+PnAygkXmzsxVEKKvJa3jCONQp8G2pztIVaATH0CXnXEOqKuTjK
S0FYHKQ4P5ulXWVs6fy5QniWoBoAYnfTExBa9MLSgcDC7vf7vnmUlUBTbgbLSUj+
jd6yKihHPG7LOBK5ED33sNFR5EhYG+L0EMNzCDkmQ6dnI7Xx4JO7nhE62I1Il2LH
NEXMouo5FoHhdNrQhMDqrlKiFlmVDqO6scWmG9cdGFMrb8q5MqJSaFmWAfLTVWbc
UshDQU6Q1+lpNZ698ApAUrLn2cl1h6p3aAyZ/87KM4uIUDRBJ69jggibSz3ob/zG
pzwQ5NsuZnSJxqTEShkF+H9ZVnY9lYM7f0GH3+S8RyDd4+QXJ3NMDQ/ZefcXKBS6
3Muw/29SbTReJLdYYiVzgZugFTSZzrJMV1E/FCFvQvhc8g0lemQ0vlVbAJ0Rob/Z
zMFGORwirtqCrjl4X+edphDZx2P9lzWKL7i8244yzM00HcitRlu8B57t5Oi4ntkx
wgNQIclCKVxxYkR7pKhEPUTAi69pzBOjVO+YfN4L3YwDbymJcTok5V3L9i7UJezp
BZeKivAYswKp4xaARLEkVm06/Cp74gXbDPaIYLm8KGK9Bdv2lzrvx5fdcgO/PLPz
ZhV2THSRPCb3rbJkMYUsTxpdjDRCEkPO5IZubLhrJhGP3sq45XcKDcBH4D/FxK2u
ySS1GKGKb+80AH36YDoTabjdZtzem0IPNZH9NgOk5JM8UBhbvmFyC339/O/OTUe4
iMhGDNgVIZG8MpDt/J1+90m83llrfp4I4M4DJ8X8Kym7b/ntojqzCHDYcTgIjMes
P5lHXygwyDuGouibYnZQgCQnV4xkGkzvHT9qBG3cmzrdh6AIUn3yZibATZkztNq7
+cTB1p5er+9nWpkrJ91zP9JkJLtC3V3SL1leZ+4sTug7w70iLOgfaBZi2LVsUWwi
J1Fm9xJWeJHhdozocsMP+H+aBpeulw8GOiJ5r10Y5wKFGZlYPsPo2eixrOvA0JiS
qlRT8QcOnasEmfA92oTxe9rqZDmhrv5nd0swFnqro4TEtYyn2ys6UXAAqZAO9p1l
YEiiRMrdS7PFI/xswYbc0YwUnOgvqbP9Ac4tTJ/SuuNzG2XHxQiHSZ7aZ1GaxS3Z
dpPOMgVUTMqB24bitwdOEnGUprA/dwDt4D9+Cx6Lk8OMoRt+HldSlwXNuRZLf91D
KsWilofyNoIHpJRWXvMuzNWAP+fxqTjIG/31bjpFG3KwWOIPwlevh+LGmZckQTOL
q2i+/KaJSOk/zAKveY/SrKBEkjl6LL56gi4k7Ba77usAeAC1m7/cviujtzQrlMvu
vXz7nglR8TXn9qi3rjMlGSjvSCf5KpjZgI95P+vgtfETK9tsC+4qK49EbecoMj3N
cmsfoRu0aBMxSmuhkqDUzJSHdvI9m4gkamHR7hBQkXbwgxauEEdfAPWa+BKPRl+W
yliq8krB7cke5HT9GAaGB1AnppaYTHjFTeJnEH6kkic4Ql6v4SmR5Wlijsblsptm
xo4xvXPij2rrgmysnFWAFAi9O4JTP1qY0gvrCCtkpmyn1AGLL8XAIs54ZN7Kg+Fy
9SMqVunhFFLsbjOgEfMcG3NaKeGtnnnNMbhNzZdyLW4t9Bni11Q4ORsZU7nB5gAt
VKIFmcpL1FZYPhs94kTeznkbKNN+VgJ5Z88AnFeQ3Pyn2kpJDmQXZ3KvCd0zGwz2
8vrGI0e2w+qfUK2iRskZmwdGjm3rrFTk/7OQC2WSMIOCXPI8MfxCDdc1wcbYETA+
BYg+lzpQG6mQ0KxV8VCFwWzXo04hOV2ntosYP2BzxG+lykEHUmLrXa9gJVud5B93
uABm5OLqSoSlJTX5eYtl3P+7eE+EeQWtwQa36ddM+CqAyZp9CggJfH8AifHIPTUY
BUuz/hQH4OMLwCSjHCMCu8sN2uR4OguP8iCGQA+jCAbh4qZb7S/u6b/JGLqJk6HZ
LLuMmnPTw0oWokpghqy1qmmbGX5tsilFEHpd03PPbPU3+rD/ynMryfgRfz68cEDL
ZxG9dKhpTV6ZtCFT7VDrDcfTudbJmhCMKcKtKtFMIl72Qbig4X/f5lALjWO3rOfB
XXF+0kV6bhbHa1dJp1iJNV5A/CwVw6WcswBie59Oprp8Gfeqrx9OSukxeAxN/YmY
JX9NrNzjSzD1A08CgwjgNJNxn5QGerWLG6570upDGX9qMECwYLjgfJ/7+HqbGQIR
1TSAU5OD7rGr4j+yxDOIqblX8dQEUxu7aLuusNdEzwaBeDPM2fgyDOk5VMsQw6w/
mAbq/pGL6kbUkuqUcxarrSz0SwGWmy66NOlzoQO1pBmuQ1a0pITmbH27Tj0RcPs8
UrAWstnZqeBDoUH130i/52I9E/cIGdIVjGCokI/VczuuBOsZ1XpMzLIDSTDRIFJe
5OUuNL8wpMFqvQCxp1c/bbTAh4GYITSKhvm6RZQX3Qw3UMZet3vshGmAhmWSLE5h
sci8NKoQU0BAQnKaNxxQL/QG99TW5mga2hNPLIRIxWp5PBLzXjTFxuNtoAaauROi
3FHVociIPWO/Pi+ktkjHTNcqARWam5Wlhy2GNg96bjWu7fTH2epKp0hbWb4PHtEz
d+k/4rTnwxqVi7aL4SBdh/+0N4s6f4QSxo67uDS5Ca1WPcIMpoHpTiYyLs18y3RI
sRqJ6IGqrFbHy/1CMm2UPsXVvYpBwXSofb01nzLE+IQSCUuOzcHhSi4BAgJm4z0Q
qrz/p00vedFCiJnqiFhzxMD64/H6IgxgwhO0SV1irZ5RKzzAjXw1uUZ4ecK7QX/z
E2XI/43HuK2++eekPNUKQ6xp6GtIJ8bR2R8cmeseT31jpCRV2D6FcNbgAyZ2wkoU
20m1YMIR8OQVTQfIvegc5X5PXxyi1q4S0qIHPv3cIo7qd9aH9nI2pYhYkjsWwd+T
QX4wX4AqWULI0HOlch4Rq452b73pYUN35wYw4SaQWra9qhUoMrIRc/329RF+HhrC
K0kQPq8J/NKkOt9DIQkEpku0stGkn7nuDwRSPgEDKnK0jGZ9EKYycC9afBGTXnbI
HEPnWiZIdrYXmNdLlG8HsfwDlBpxZqAASnHw2/tpY+cnHg1U5K1KwlVCuk5hj2Jh
i0vtrejhAEwWPw6pVnnz2IW2y6q+mkDM/OK+83TOf4jE0OVYzzkRIBsSCr095lUs
EQWKW02Kb2U1wr+HJ7dcmPV9DNC2OwDFR49WsZoBJdXzzGrcw8dFqma2j+brxAAT
3iHrSJr99oif7+nDw5KG05ry2AdVqyAuVtIU1VFQ9SCkyVCOpImD4zYDOE+rUeXY
5EbTyh7d7cRgEc+IEj+xD342KXMBaYRSI2fkyShwiHgD5S3EC5y2oIX9lYUpmRBS
SYSq280BvaopPBCX56SLjxs3Y0hjOEyzw4C00DLhIo9amalXFI/KJxn5eqHJd6C3
Qx2u2yYjfpbqbxeOOW3ducrvG07KkgmCySRuMXK8S/ufpmiBg1qmDvINAG6/cYJ5
mHzdrqgtHT5W4Kbr2tn2/f8Smru0cWyPGFcYt7ycKNK2ORN90QidQfKQDTlpx11B
9Re1IYHdaf2a5iMDhTQRshYEQOTxrjSNxRS1Z+h0cNJwvgZUiBnIQNWLGneC1s+G
R95hzqoySjmx0x1i4dLfOydN5cB5VTISs/SABeBzizXSSLDBL+opEXZuzS9TiuXn
gznaxMZmukGBve6UXXZ7w95eMmvJwgvu8QuLmy5sTQOHd9oQdZTduwTGfzToztQn
/TvaI63nutyKEZvI8f2FtZFkT9y0FlpPKSNBetgFotI2scfLrIX3zqHT3XhO1P45
0RAX8kY1RcOxmqdLeJkszINwTfGNRnrMGHsz9TQQtjNwScoVZbERDDQT/tHUKhGb
tmRAc6lmBITXaoYTHUzv1qXf2AKX9zNLqEUHMMfi58UaXrz9XB6DRSilExorHQUs
wfpDaaR4ciiylWXJ5W4KArFfxK0KUxdzk0Em6yJyy7AHAfL5rM6x7tVfoqYes3zq
cnMoOZOMmoPn049JX0TAXxi2+JGlgklAZo6yKat5iHPICKS3r+pJWWS8wpWBEVZO
2T5fIygjxnZTNxMhkh0z/gUO1Xw5+laBtSIu0pd6FAIPaT2d9iraFtBkHe6L/hXX
KVSRRkww5AWAwLFK2ntt2D6wOCC70epoawsi6bD4kwnicL9lYvprlnps+Ab79T9z
j/iI+S6cb9uKIa2rZyDaBj/bKZH7pOxK3ysyveXLWCRCEyZKw8iWETcHWOO7h725
Eudd5kfOLVxLawzyczEgTloJjVfMnxy5gE9iS/xCuVzfu30KMXIpsdONHvXCwmrn
1TGY4KO2FffM4joyEYnrpQghQCiwkY7+InC7j5HNbAg8DGbIb5zQ9U4R7HwSWl6j
5rrOjNHIHyF44h6Fb2bnLkue21mLs2V4134VOBBBYpUucLHmsUNsuzVtIv4YJRIs
vDC5891z2SVPIsZeG5/iMZsXX3AITl5nwmQhTHRGZ581nXAGrMHBCB0v4yF7oJPp
onUbRXUdykB8hwWh+hzQBkHS2PREhKdHOTZfyKxqAsYoddI4Yuj3Upaknl//r/Fj
IH19iij7Datd/a8q2F7XTJ5itzJ5m/7fEUoq15htK+vI5B2V/0Ujf7wXPQX9ISlv
mck49SwkoeaozIOQz7l1J53VBw9oXEjeWILeYEF6aFlJ0YsWBhfENOC8oa3bYVF5
zvCqtkCp+bgsnreg2XRolneZUrBAY6ytkJMGdj7CX2rU9hRtzd+3cGRa0VnqSIgP
KfoFRTald2yk7aY5YRSy6CMf7AbJK/XVHFzgrDdEgZmdSihR2S/9LYu4qS+jL61n
zJp8Flungoi5/i89hZKSC1UM9NcTX9CrX8byp7RS09LJWvg9B2CHcciDoLzRKkla
M0Va0UAKNqhKjElTeXx87THqS8eh0xGwF1vZjZnardgr8ig1DoLVedPFb6Kji/Fr
EcJDnwJATyLJzYH/jQ7nAsgzd0LEd3BI8KQbFAaKOATEHPjL5hFhmcW/mJgkRgng
tIReCu2w/lAxHL/1OtHzu1bE0CdzsHksXUy3pIPj/MNtp7gnQBk9NaRgIvtRg3Yg
Q/VtoOUPl8n4gNBGQ4lQBnN+fOlM6awHAxW69/8Bm9LY8mGIplyATdzRfg+zhvBc
VZtLnJzaTgyN2wRAHlecWU4XCyviQTj0rdxih26pabzl01qiH+IHR4xLN5t0V5SI
RrebHyJvb6ug9wdRtSKZrn/pXF7xwbW9opToChpJG7i5eb0JgXVm/MDS4oFFDeKv
ZHzkGxxb52wJrd4Gu5WyrfsFtPfr8/kzLc7X539yDKz+6XxiWu1OD1gc2dzadXYs
SUQBgAf//PHIm1CXea7HdFqT32w94KORbgnzFMY7MO430QOqDKEsl2l1yt9ravgg
6jxzfEhn/UUsSvCSDXWOCiDpyY+Rk6+KALuH/OyG4MqHYiMYsL6Mglrh92IU2Vp7
AC4WxFuFTIXhz4SanvMN0mnWNv68y1AGBYJwJ4Pa0IvnLotmA1SuDk+ON4gG0H+H
VEt2vWkT6Di9XOipy+ztRpSFl2gBJHTfpljMoJ3O1BGzG12bSSsIeT7Ch5GpPWiT
/kvg7ZaRooar8+QOW5DjvRaxuzwhO6jXk0YZc0NK6oaHLUlQShrBoN/9DkItCVTA
u39dsvWwd4t/Bu5h6UJ+Bel2JM143l/ZQvdTlHfIzVxl+0i4kJyUWKj58P/f1nlR
d/Rh2kHXvPZMKwic0h2MgSp0G8E63Bb7H8w/Qj8CXySyEN/cKEALrVKJbFn8PyOx
uNU5pVoAcDjCJOZ4aGX4qQMRX3V4X8Uo/GOwxUTywZJRKYpta4WFLjuvtajRy1Vg
5FcE8387iOXrUuOq+BhgnPqjfbb+SKLaeMQR0QedyqduUmqi8vzY7LSfkf7f6Lyc
8PbR2e5sRW0vDkneBYsmSiEHjVClk5qciOgG3NXnqCbGqTX3+TY6DYwbREugkIAL
zwGwW+1ivObyP4LdF5DKhBd+SlhWAOaViUWth59J5f5fWwBvuQJPjhL/nCtOzj7V
XHCbxwsrl5pf5ZQbOPZFDI9aaHApwrfQEotcsIHvSAM+WrGF0+R3m0yq6gV1UXPk
EnDBj+imeikSD34hTCAZz82+FYRLyGRkaGo9q/PGFlXmEf7qX11b8ZU/VZFPRMx6
xPQSN+ICkpC3GMWi9mvYsOZHXgFzWgz1Z5HbUEWG0fO6rYKEhG1JCBfJwZT4OPwv
uyQzRdAJ5ZIvUYLRPACG30pVWGLp9Il5VzY1GjEnjBvgW2YB4Zmu5WQBzW0TkoU/
FqJIW1jSjsHpGVAJDPQnbgzQN4emyjXw6VwZVVxHJgnu8nRDIGdm8y+b5qoI2HVv
AsMOJleS/is18vqhWQrjDIOc/Vy1s5/oTOrAIKL9BYxHwD1V+oZKkX+s3W/VZp/K
WYuhiTwtfN/cwea+r58KltzP3hKCEQ+n8JWhzv8kYbdY6BgTw8Rf5YMpAOXzpK2R
6P8X8T4gZ03/fvEhvtK2fzc1TVLTDIIBRgXjhPlR0rHHNfYPBG5cjiWOJ/pnUNix
6XVmN9juQ+EHAInliBsIYUtof25Yznd+/xPNW0Rsx9kBwo6FoUb/RxQrlOLQNyhh
m5V6/cTIZDsfzlUQ74078kB2HmwCyQw8+BCV1vE3b8VAaWpth898n58T0Sa3+Kwr
Z9hwHG7NUWaeszc84+kWHxTL1nsIipRVtIJ92YOEdYoM1ZHHAysevbNWYv8EU18y
K/6xMzWrOdDrUWgDdI/wzi1qxlYqMuncxIxsPpKsnsGEu6d5R4EgHABqJfFcv6u+
0eO16QGSfKm/kMyFGDyGZQ26vjQ1UIWyyQIDGGQxYgaaCsX9lW6eRJOg/KIdxps7
N8mCXNfEPOkkMfgewHIKn2yn822Fnl/RU+VmBnKUlDREZ3NGCdzelXkcFRxGe8/j
F1J7LhrMjEBkRpHlLzHAh32P/yDpRx4v2T6MF78HRlhGBY+DVlFB4MKa7UsFmWly
E+Nouxm9w8hAHZ8I8yrdF8lV7rWngR50DNxaKdM+xuN8tT5E0c5xuiu5H5qvVV61
M2UGr2ZGZAcQzH0HLUtxL5+Kw2i3HOrIAm80fXFkgb/NuNjjpdDrKU8chsv3Degx
1dThRr45pA9KTciE+ntYRYeoelIkRY3iGH9WsSOSIVFMePRQMCQGiHhTLMade09q
/43LFwye54o+acpI1BzwYgndORd12j1djL7XDNh3ZxAhlP2pZb0QeJotwgG64AnP
xTyZYtMGkaDUnK/TMGsZ1WsHZLbJ6erhKPNwRdDOI54SKY5vnKEoqy449DNl8RCL
kn98wNMjOn48VgROWfbf9abLDIuB5rxVTyEU09nx6eTOQdYAuAPpg/DAB3yEYdL0
d2iXsScwNcu1H8djpSviEc327GwCiU1yqS7e72EDUwLbA6+fZLdx4/cMQj5hzq6X
pksGDvLNeQ1uX1h5Lnrx5kcNzKKHvfBnUErbMkqBZ2LUahMC2LsankTDSf+tIa7X
Edk0MnwSELiM9xn09XMhd03pnfYZCGE1CzIrC9MSnLWr27ewIWYll7id54mZYjXE
FTe6uYxodTZ3vXW9Mt4D/Ku7Z6I90ICAs+rzTLVOPHxPtyfgj8KF80hIDeQwwX65
x2P2KYiFAN48/ULv8fo7eiOWTf1yB4NsLTt/au3RAa1SFZTpdWRJTj0G5C6ablj0
c0TQ9/aFZ+lmYgLAtaYgY3tIrcVC72rctLFLbUiWM1qYPpQ0FQIlVVcybLZyeimf
R0oIwz3WpBPLdd4UlPxkdORsn+s6nR9nS7TGpvX6latnCXy+ca2E+b9PSs4pTnYG
K7/dZ0i16AAeSLtlW2+/FrO4ZDIA51+238RF8bi6n6Su7smiuRGTdPXrO8iqHwcL
q5sjZq/YXLHwkxL4gD6f+fwrcLeofX83m+pYsng/rUE0yE9Rv96787+CTvA3YAb+
60w+UPvPaglSaNl1tfATstZs71rgWxmbFSYTXuorFaasGCnlk/rW2JZQCdKUcCbw
QSjTIFovduBEexdEBbyy7am/6fuIS5nOh0dNZeELzyKOkocfu0XoMcr5K84e/XxF
X394NaeG6883M6Et2FtPNV5NayL9y99AWOPO36Pq8zRl7kfVB9FVPgnM+RLBGI+Y
sFGmusz3CtREoj/Dyqfu2xNISRXgt79T+855UXLgjzZbCOpVPpWhPwpjBmOr5QfN
waCw0TwZyQuLi7IeMVpTMQ9+G3JkQoRDLTZlS0VifEa7hjCIC2zbF23LiTxKv6xx
PZHbcAmeuX2E17BY3AnRFknkiGOp7dKCV3FMVmoeevui0s9IG/MuMNWUhpQvFNOL
L2sNsPENYdeFLTwOn7jNxUCHjGFRHgp4onKLjpHz46IPXzTdhj4m2VBjL45cYeW5
Hc7vYzWEOZRpFLQoRzVqgrFTrpoeRDpOFPS/aXMYWnPOeh/CAExMQEY+geBYsXV3
0NK5oMrZo7hld4os/+t5SZEaDbMzR6PtUEPu0UVFIp+nptJ1r31ApaIqxlIDFGLt
xUJVnpoRYqGxA2wJnFMEEofj614a9SLqE+2PoymjsY+jdATX5b5EtAp3+11IEV3h
npuDpWtUndGK9pbc6TnrhCZ8fQ9cKXSP1kWuLiJ/bEmjskltcmauQdzJuAc4hiud
qT8UHKOapqiLjnyqmlnoITCXgmaU+4Y9gHy6A9fpPdTdvrTmMVo42g1MGmLuOgZh
B2x0T4+eT2aBVwOTqgByJ/hMOuNYXgE6AYEUP9dyU+TsFxM/2SIAOoL7gY03dQ1C
jx6Y3FHwo9/tu5vX8jgR7utVZWxfTJUfzEbdpxxSwA/mGxIFBcNRfVjaaE1uGdCx
UVeG1AMPbnaL8KiGayJBjg8iDJ727+1R14E4BfY/v1Pr8OYQbJ6hs/mnq8tXnwzN
11dVWbe7dLHWiX+v61mV3pq9UhqXMSzwKtfvo39ZblgXXHN2xTNUDh9FBIbHSknN
YFwEeyEuJt1raR6Kuha3UTR8DXbYy5X9ZA3IGtvu6bqvWAWj3Mwz9tqb+M+ru1nm
Uj67nv8jIayfziOAjW+sY/zT78XD/UNVqC4+83GHsBMKNnNXtjwsE4hhR3DJi+d1
MdapiLBmkwraN9v1E9dohKWRBzaHUyAaVUKsuECPrSbvqG7sHP5xElY2JA2dXO4r
i4xJHvBZOkbIJkkOP6GGL6iWXmn6G9cyE+yVftuvY5DgNeSFYjhsu8SZqp97uGPV
vuczjIV0JaxxSCgrgXoj9oK6aHfu8mdZcFKrxryxkAATrAINcdJBBRqL/UrEUrAK
aKOzb8psyF4qYB6iYe1OG5R2sFo8u9hq6crVl7iOSOQo97Pj02xl9bSFTGoE0UmZ
vBzuzZvnkXqqzXSC01V/ghOOD6bTzEW2kza2HtfGJtNeob0ZuozIgQVDlu9J16T6
9+zyfZ87QeBb6aQq/mZ08jjcfQXSwVZMlS3sUfx996GFOg/NDD7Ovs3WBYAd3UGK
MgN83eXdq33oPYOzWqFnaW/YFuOO8VZ4IWmFnikeBIlGnvZ01OI+AEQBgOFF4YoY
CVi56OIck9P3IXd064QibvrPZ80R8sduLyBHhaf58B3zM3jxZrd5JAL1KFog0E8R
COqFURS6u7WZkVKzno6dnrCqyfdJ1XfT59BfFJQx886VK9UtpCKUrje+PlTSu3LG
w3WFieFrzI4Fz1p9PaSjUxLsffmCisUCWC7N9rV7FgtBKXZZqTdkotKqhldaItVe
whT+ZfUXSwEFNWkSuD/+eT6Hx0lbuLwdunnIA0K8zKzqora/akoOce+Tcf9Z5vF6
JjSwqFugb5TCWDqRzpsBNiBLsI/GsWNX0eaYUtAsHyQfXagL2n0hK8w+WwJ0rUJR
sDxS1EtdiR3wM/XTWVske8bbUFinfJJKSMRjz0b2zJggkmiL80OHy780sioLpSTP
ilCnlSEeN74wqhAbB17M5xwYKtiQh7owNnOySzoc0/GibinQiAGdGSwge1W3yVSe
6W1WtpFGa+Se8miyLBMNQE3T5w27yhxZkuqHi15M9Hp4KzWCEtC3yeG7hkeG8yIj
WLFpX8jdNycazhek6PuOD6ELkcOIwwPL2lqZ0fpcnpjFbeKzqLjC6fxpIQXmQ0HH
nYtJC/BKFIlaIp1A5DBs2DQ4D5+pkq3sPCJqgKEN1hG83YBwV7LcpW/2VC+/H8om
ThO4/QMsPiR7YUcxGMTaq6tRd29Z3Br1Fp3W0HdHH9nWl3fKmatpG7i7aE3m0m2q
68AQ64oza9whEEJvkFDOBpU6rz0zCrPypmtDlRIBA4jafKN54HraHQgjrgBuIf/W
GJkEi5B2d1no+4zPRIUMmwqMKFeeDAosw5EctZaKQv1wZdVNAH/Xo2/8pjH56PCR
p9qEQgffRuqc1Tzu5vtiTVf4PnEIu7agfqlfadJyDltFUSXgDsWOS5G8j0lmeLL2
3rqfL3JL/OOB9N0bnFQp5G/j/DceoJlYNr97t2pi22AhekLw5um/reBJ31GtZPMu
todQFfEFvsk8K+uEh6gcTvAC9OYMgRVLiA0rfuf32efChuBQemsoz444ZFjRjdR8
vycmcKnVPPuOPhz7UrbBqSiCYQjd+Kp6yO4Ii+J+yVnqtWiwogAC8rHhuPpUoJK3
fvdJf7iuAb3JD5kNLppSxjUTDIMbOvTWE3rGEzIDVqorWYwHZQ03pgbrAoaQoKX+
hq/KW+KwaPsNzmKADo7Qa8E+ySL37X2yEun2Z7sJJ9Zb7RBJL0QaT+kHyArly5ju
x6jfx87qCHemzLEQhBnzP9T0mZEtp1a8eeR8PqW5qfUzZU1ClbIygPFUFY6NzPAH
5Tyd50mXPwR7VWaMmFkgIZ1z0gHdRM/RstxAKWVrKhg55nA57GYoWD8ZMHk5tprc
L5LPNGo3RyIOy8YFAHg8MqYU9I92Tw5fWWqQc8unit96aKJwl1ZU/Itu8WmF1Qv7
owYFrOkDxw6gD+aT2F4az2dO+6ZBlN+HGBc5Dsz3jhh/+GXeSDfc/gjwJ5TDO2w4
KbhRaJZM23ihl2X+ApHBs3PfC95ZvrkdKj7CzebytyOn8+Fr920Dfsfl1hFmmyGN
s+ZJLqKIeiAR01jaR9Qq5Zko3pLILkU1kD44s50hRx/Ce/fEvFpUGL84vppBGQHo
f8RNxNdheLrhCQcF2tdYNT5JSekP2bV35HuTUddR/1Zn2sGwTVTdmMALbomYevl/
Cc21n1Dk3gQCOtgkHnVruPFylABD4zISo8LkegoJAWJeZl7KE+QUmBVI1qnZcfeX
Nc/nhXlOm+fZTn+3SyELeJyqbP2lbw5mQU7LsKXdV1+EvH+fKR6jaHhLyASLMw7Z
KvT3PXvFwiqD68mScwCrt3ZQqyGqNKfvaqVR+naXimuyzsBjpAQt3I2yyscy+cbO
ZwgTf3P1pAEwfyWiuJLtgbUfiR8TvsD72Ct+0yLAgDx9viiDbyVCgBp3L1+WTFjP
NGjGWDPB7yhKABjSbBcvqyy7wrAN/dBrR3OvAjwTjUKdf56T3CzbeNM3lk7ASUGr
B4hCReOMqJKiLiLFwjGt5h5Ty0x8kQWRC+6oMftBHfrYAyRjiAOjaGwR/vCeY+Gj
tx4d3wo1hTiZuT8XwiQgUSyFkaEm9KPDpfMqahxf7pOhe5s2XfcsL5ofnXp0mXTX
Da01AdhYM2EOFW3BrcHCbxLcrwClxfQSzwOG+mAhsdqBafXaPYAoRQ08sxHCBV4E
RGfPw/4B0BHdcxI4qRya/+eo05NimjuG/92zjj4L0p7+5p66+BGtJdeS2Y45y3C+
q0PnAJe2h96jKIYHGpYEZ8d4cOJ7LAkoH0MCYYuK2qna6qukpLi80q6zMxj6gq4Q
SEZTXGgfHQo/UCjyl7Bi7mPIG2D0D3b1dcpplsVtmy5hrChJJ1l5TRTLJ4Q5xHMn
sTh6Pdc+QG0R0h/wcBSxPYDCvWlRlgpAcjsAE4c8aB4SgC0PXl40DlPD1AaXavKD
sgAIeecdGR9ZaSZJmji+lC6wWQL6CGzfq2fyxnD1BqcSPnEotLWQqUTmhQLEkef9
qlJkNQxX29o9tapHbuZm61gFDYL9wPANZRBiCQWGnCQAtIDo6HSyumdL3px6nLqV
EB+LG5s2GL4nj4lrZLrXzmmRRlhk2j3Rzhz1wNtY21JF3H+aOsbO3lxLddVeGR/w
B5aUWfotmDN3xze+K+mHBR0hx9VauMJSnL40FXbd0QLjjUHR7vtE2befOY5TiJBh
2VRums1pa42+Y9JcgKwX6xjO4SDTzxFDhVbnq8dOQzOBOaXuRVqDXkjUfpZs9AgI
gKS7mOQ3D3Fe3hyzRplmWCgR634AdB2pLo5TDNtvO0C1a5v4gE1TWYgrUYqIDEqH
PKuUvZoHRY0eLgiYPP0FK5rStXs2jB8wQho/IIm0RDQ5z5n/ZYKWyHRFK4uRtvPX
VabX7iCMoZMaZ6GbDA9HXlpFqQjStKWFQCDKv1WyJx5Ro9kfoKikCj6Rp5HcOizL
OG9SQql+c1sdHY8rWNPVWfxGV5VxwEXnKX4QGJzrFnkNLmClgpNtYMc7vqUoNkSQ
AHyYGdIfE6JvcLgwaxDu3NfHC7VZTGtRlrdHX4seVS27Mz6BMUXAb697e28FmM2q
jkFRBujGT37QC+qqOyczLVoTxFDGZGWBpVogoaaRmgJwaby3MFyuLbL2s1dtq4pA
O21RNRDE9kKSf/9TQhcsiNpLdiAouNxczg9+M8vH7TflvnqhbpwXdmHvku0z9Aqy
wvnCaYLpkHX+u4SdoF0E0lmpe4nfxs4SN6tS6NfSaoL/GAwZprAJL6V6OkVNusD8
xndDBRN+hCZyv+87AAmNt4aJmRAaei7DHsig0EunjOYpGJh7TJEAYPbht2Y4XETi
TzEzPcyBVdh6abLnmYq8pqGPMyMcTl4qyOp5fxm+AOp8X/EcGEQ+IUioO7MdBFA5
gw418hjlxZ4cvQ6UjLe8EnPAdFxBP/zrAVy/2XB9MUatzdfEqqSacJr88lB/IDdW
a+1gIkLp44lj265oZTaZthoJ0/kfohqRh9+DafBUx4RCNsPZVDaj5oAxooErXUfB
gW5Eh22PUONpFtwKwoNWDSihK421zQhd6DJe9WTEOmDeJ94HZXSu8yCphG8h68LD
29C5Vh9o0+4pg2O4sC7ax2ETYh5gdsVn/kxjlkv0tz00NZ0PGPSAXIA8H0pdolr9
6SBV4iDYxjccVsFvRSagaOpj/2yWLlVil4RA0y4N+57ezsnDa3HC6/13m9q4p/l7
0xdCgEjhifWwuqFx89R54bVXy9GJyfeQKWilNkB0bTa5zNjD+ivmgxNLVnYyRGK7
v069UQSPjrFUSy3h6AYmZdqlZ++d31AmLmc28BvjWUx+ovSKT7c//CAE/dG6nri9
sab8qFZBYJlT1NvlsFBYWWKVz/65a3xl8lTq0gN9vq6cs5n+uWJtiecoJCUJz+9G
1Tx3qGMBjiiMzGLifC2icj2RxFuBbVI4BL+uQdckONfRIch56TB4d1KxEt26m7Dt
w9Mf4O5SX/OV3aTJfdv3T8TbBElmEOrq8CfTwx9UTC/GS3K1f0Jlw3xfN33IuFAO
AAM3D6ba/sPAjQIE7rfshhxe1LQGM277OJp1CvWF6jPdMMUfGXs1Hne6tk6OfW9S
7OKscDSrRH5Z4bw+Vy7n2+ptbpSY7Q7fqQnzObdtVvFTNIlxIFGpNVweWtKTOOGe
7bC6YwvwuCaL14GFIgQtsvcfY2FpZZMur1WpdTePIECnbJpnf+cuTaoFpszPpfhJ
56Z8qlC9Px56n6HvlX4SgzkrLMgO3EAElZ0VI8Cs/S8oZla+ToJGN9kXmzFSuHV7
RxfeU4ja6FepJJ2ri99jkrWSo+eVyb3a/GX6IMfbI5pRDVfGrA4uKAuH7JEj0uLj
CgiaxPif67FEJYbqD++VRAvoWPs+ToW1xrArnyQGZXDp4kR2lDfOLkAu8zq5AOT0
yBqOyNB/oaRDOKkCV1a10D05BhM1nRoyEJgxnxUwI8EhSWDoY9v0wQclwblbBlJA
xuhgGdeqSAJPKXJf/pAel+qxBNufRn3Og17MlxF56UwfPnFrElPX6uqm3j/Uv+e6
JP9ryiKbKrE3mFNQPotbRDDtKsRihcQVoB1LG9tn6qfIcQYhoH7XOWB7ONFVs7nZ
FiWc0QpK9tCWtzB8qHtJBlomNsFP5JN/zUrSnUFlDzPCNzK0znobH7po1311pd1M
ZQEMuBlChyI9/nokGC6YWYWjVExdFwDoi0rB2kXki0dE0g5coidAvCBroYy2CRjg
hr7WCdRf4JZ0goDLtLwq6s9339Yr+pY+1YFac+TwkdKDoSLTF38IeuplYsVYTLpo
56AYdu15CcDKF+ZJ66aZw0lLrPwQxvTwpqr3RRpjkdYIx/dJnTrN32SdMuG3wneU
0gFu8/XZ8keE85197fKGJ0hmPB805WeOdzyC+lPMre7Meh8nHdWMcyd7DUcDGjkJ
5c4VtxFbov4stRH8EAFqxKXKMYqowEbErD/Om4nqQkXwa94Vvyr89vFoHduiVG5Z
g/VSwjjpcPyFyhHWUl4jkURfuiJNBE0QZM9xcw8DEL7ze3A3gdpY1xbpx2iIUODd
dOirtzt0b+paiEhNjA0bmk/2GKQKG13BT5uzEbEpPZsj2Q3NXdS/Jc+tD3EbNmaK
l4v01vGNVXioYl/frbtOub/1ZMfyD0t0GvEcwf+3JWz3LSvmzWy7nM0YJ0cgn83K
6UhEloGjHg1E5P4JT+Iq0DIxjzlBNxbHfzffDHbe0ke8IYTtNAl1mzFRp9MtvYf3
8dTxFFV4chqlwYhH6fBXw+K7sZ20DzXlSBkFCAxliDtTEt+FTG6QW06cWR07XItc
e5IdeZecf57FsXCwSANkJGwwc/tF4Yaemv6o95YY+OwnbL+rIBNRsPkSwkCZCtcY
dOkIK858qp7yc6ZjB3ClYwZFETjaM+WHu0hjh8tdqQxazUAry6QGhT8KnKETWvVP
qRgGZ9UN+BSD8EfBxshHNuQ3710b8n5mzWESCtZKt3a6LIeOgI1Ea1SqU1MpV7lO
yJFIZRV0mV10rchk5TEZfVcy5zHEsHbzXPbMHXqqQ9AWx7u/WkFwTB2sL1jWkW+s
qyAD67QnV9BrSEw2+02LzS1tX3AZ0YUMJgx/AJ5wpFiyEHz506g1D60W4WGSD6Wq
3ElUjbC8+1AJ3CU84oBnaFRXisD/Ds+bwFXoCqtgrOjtz5sjw91zOSavxv9yByZv
rnd0MaXX9kqfA9cb76YIOuYTaVu4Su1iLEZR+fIxzKsh1bhQMS6wTqNLvsNnyRvf
2YnwbMdW9HfAcS93Sz77Ruic6IvjZZ7cceloPrOP1aMLEyD7y/tpwgUB4IrJX4HU
QLiyjpWN8wkbS1WHlN6QK0L8tyLAtroZ/CPMToDVEV80U1pAjiWdbCq7YqQeT/YA
uF7SGD3ln1EyX8hlyo2DiXkDVOrjbo9lrXBHauLi5IepeSmkzQfYOgiveBeKYOWj
S3Wmw0BNcZDz8Fo+8+iw+nwOp7D6x/nq3sXy+8U9ay9xxWA18emRQbo0RnQy/yet
37/LSgFTgQBOX+RBtnR2mfxDLXQWfWtYUlIcstnwGL94Id7FBz5EePob/f6NtPOV
hBPoI66ODYxC9cENp9EqsaEWX7xuFcydIXvsj3xpbnpqLykOmJmmNyGEpPYhaeuf
FMT+ZdVCrPYzW/8DfCVSkMF7rRY2+Ct8kvJPqiRqSrP6LkFK9CAiUReRiQJ7vy9Z
dF8iZ+Tn3sn67QegiP+d3HDBhzJIPCCLg4VQrStUSHqEqu0zVbDGnGFS62M3d+UI
QUW8e6D9gSUgmCgYyIgRg8p6qPsr8v+JNSTt6OMf89yK2MmwIDmDQa8uN3027maX
AC1z7hAh0dPlAPu7ccFuTY+y0PuI2szp5aP8AGX0D5FsH1DCui4DUgFtNkqCbrNO
lm+Wy0VpXuqxbxcdy9Gj7+tNF4juL7EesUwcnD+9uFUOamSX1y1WPMx6nWJe+wRr
xJ/BEnjBhAK+VoiHuEoP4fw5dCnlW+HZRRCUXs4XaA5MwF+IYEeIpM0dFFq5xT2m
jSSJE2LOQZ3kFxacV9RyQuQwe+DFfWkj23Rsn7jNYT8DWkiEoDwjhhEIUbkINrOD
VU+qilGKIafxfuvPIC42JBvs+Lkzw7syMQTXZZU2UD4xe0ceQL5kHcjAfDRW2xJd
apdwyLVMGcJNMCqgmRp3gjV3arjcr/CXqBeI4QTRZInwckmy6pn6uHzXzg9AfTix
WN1HOJN9ETsN44CexwuCkSF6mijPCY0mpLgUV0iyv7BWp+C0l83/hX3ZRkVs5T+l
FtZxSBgSYgxqTBgSWAd2fBEvQJywRQnq3nRjPeVUdtZWacD23NfDxFbBbMq7RKl6
OoHU8fEa6v6mCH8v2DPwy/NsuZpKWNQHIHLSGX2xrXL5fZI0hHkDdpT1RBItlOgh
H0ZOi+HTdY1Vs1NrVGRh7mJ2VDRc66dAH9Orfk6pq8muYZv8MnluEUW5ftVpL5d5
QzTfaTgkeRTY+Nij2/BGAncK4chPIOJAiDfHqGuHMM39OaNckgr/VrZw46TIyMmn
ecA0PiFeDsFDVMTRR1J2YQ+puQFVTb+AiU1TjC/vP9ed1J1lYpnxqeYKG3eX8vTn
jCZ255P3Yz/BWjEKNksF0Zdnh/4n87AGp2CWWpJdIpYUornx5gO6dBzVgZnl5Hga
kcmHAxZcXZCxKADJ4jNI+DeLwWK0ByOKpwB7kCRC6eHWW3yH0n+o+B+/nO3hPWMj
HZ2hlKywlTaToL0o1vxnJEDmsn+NNn9vtIJjc50EapLRM7NictVgE6jUiJ/4yY6k
o4pqTg3ierqp0ngB+lF5fSQWroPmabHotc/cOo37Iwnhc3gdi2+dKiebiGTx8bZx
Cd+QyMk8+G6zkV4Eze8XZQR58jp/HzqOzbFOlx4km6OPTNr/s6KyhNNpboCup/6I
IHo0vY1WJYbYab4N48HhqOwwYN08BRxrghgOjKXNEZ6e3OPIiVNjAzNslVV3g/Gn
SOPJ5ReMdQEHZVaTWh5+LPlsR2cSknfDZ+82TV/12tiF/CqRbjfoZe1zMum+fqb9
IfEHNS/Fx79s7wRiNLOAGq5ngq8jvJQLP+e+qPhnWCN6gar6wB6zNgs4qoZUEt55
AAzqAZDtE0NT0/CsomqbJLfgDmIyd9N3Y2XZyRHfrmgufUxmnlTHQXiVEIYiLnUj
T7mRryHRXGqF29mekmKwp2sRr3eR7kW0ZXj+lczlOatgGfgatjWZLwEkvk3wZipm
rdCJdUKqu/Brj4BBzhrzy5iiVl28aTC0OmPqX7TVvU+gIty+5Teqvb9bkZmUx8gh
mk2KhgSU1gmHQARlPkaRls5yKzMbfl9tUIG0uYfJ0K3h3S+ZXSII9aNxW4NQRzJ0
qJ6soT66WnY3YnSkPbqXA8ZK3JDbBgfVEZK2dQlcz7MA5+llFj3CVgfXjhZ6wq6B
zabyKJr0npDlkQZaEeDNWynfiO6nfZXBvAVBlABVtTg7F02oMiqOMcWNYCk1kAlg
dUWgyntN2U3O39KMl+gsmYZ/HmBLLUhb5DWgYKcfFGvF5imDB6o2zvBiq9h645RB
w8PakCdK7UbtMDMTazY4qJQFGfL+OaB1AVKIQGSrbAvqPbIax+z2qta/SYKId9ys
Vhe92eoBRm+mslFBmGu10ej3A6QNvJj3w+DsVPiu8pfFlo/ifz+M93OeR+tjQa4K
vuClJORxv41GJbSgAcqRoUlAqlghs5J+BecaNh5jH78v0TGef3OztxYb+aQiUXFf
RPkwKH55buVNr2fp17zVVpBiUQAiORztgFdOIpeulMeu/NaWiWqWrR2V2VZzKpSY
AuxJwlRRm1MW7E3ceCmNVmmx43UsBkQKDYYBu70Wkrrh0kAsICxbI2ysQazB8NMD
4ldbMqqqqdnnkXuLSReEIBFCgBKgjKFwyNGR8OpSbAQUzZ/n4SxwOYLhAxhGnCsa
22xSVMoTA7tQiWYMxDJnlfk68fv9bDGEoD36VV+meS/xwfn65dyeCENsYbZp9Nhv
X7CWeT6vmGP+GimKG0SkZGDrQ5YD9a4VJEP3kac+GBwRlXHtaS4CCwgVqL2KiN5l
AmSuom5lnXoHaQbLZuP+7A1MHFhYe99UChMp0gJqZ00qaSTmO6VFL3iCW2qSa4Wn
ELGIapQXP8HX+LgE/ZrJSvRLXdBQWkZIaWTBYJLtIZU/S8uvRtFfsE4OkdVOZAkc
3PFQLJQ2OJJ7/9NKg6cBrvu3r+xPh/nog4WSVajwav4QCKpKPU83YLXQYOaCNh8x
pSQ4NLP97C48QZ8cJfVVKtFro+t0I7KOhff6eVl0AbbdsfV5PUbysSA15WbJQlBw
He4yubTr2B47YXYYTJzwAjxK6ZlGKbPBkt3KMA7PCO4gtJSLernf5wsiZCAdS20I
YQceKP4P4hXBQ19XKDy2wTgnPJ/jnJ88xXYkIHl0XWxF6FiXAQgihiV/EiX5JAlf
PnUZOsBgaCQ3GxADjewys/dMte/HlX2n1VQj9XP8vkjs6ysmwzXYr3SXwo8tnfiY
Lg30y5cfEQUG8AUD3IYgaVDGgazRjf1lov/d5koGSFJBoaE4uJi9WDzc43tEko4u
ye4pvADD4IYLOQFBvaPu1+iyPhB55d9PTtykzv08en+LupgO7/kF1Whg9cUT4ilO
/XVOjwBZvcGAgjpHnonkqiIhg+h2A4T1fEJgfd8zrrbjczCsWLzpQBf4H9QbU0dr
qvS31V5Ub48+IQTtuXyY/clZBweryd/XZqDSTNm7LMdNhfPVQjwQVZ39mllJP2R+
evwXDJYmi0J392O4ZeVH10UwAR6O/UBvAowP16X1mmBWajcJzGFmwggbd5ek3Ag8
AfSR8N1xKfJljOKTNd8D9yewwT3BYl61hwo7+f0v91vUZjx7Ahz8GQe2C6czhsII
ADxXwt61Y1MGTpHWEkHAg8sF0CiGgxXV+e0jnHpP8KCM47LyE785BUOFGTk/MU2P
qFAfJD7zMifNW0d7nQhPAL9NKbg3rkywAxvJ/wo6+f1rDszD3bFHZJKPLME9TcFP
A5x+/lIRExwgE/u2q+TLWfbW+UeWDNCpQZQwpbnQgxVlVBDbL/UbFKuaVS7ZcXYh
mkUemEABewtWpS1zLVp9GnziOK6V9ohpuxly0my0J0vT7O9avsJuIZb33L3iGc4D
7olYTlTEa1wyQqk6M2aJK34n/NCW5fsrPgIJfytsOyyg4+9ZP/DTHnYvYFy1K+Fx
qhETkC2/WUZQPjYZ9DJrFPn5po6RMbr+PxJkzZqi/tdaDuqRwXo2EqAUyhTN/d4Y
GQt+I+k2uXxVJRhqDt+eALvjrg2Te0GFd+cA1Es23jHzgV3kRz0GOWntVPHj1sFP
AOJhKNiaahcAkvha2v+laVAdH/BblJYRVASjKyAFAlnidexWa1PG6UZruCCL6fL+
c8lfKYoGrU2pHRIGDdM7LBoUa8rEEtzZrtHb4is5FGSDIgszYnizjE1iPRQ1zq+o
rbrs8bRT+oX7nmN7JMwEEt14CQIX+4+QWkvog92IhQCZiuk83WzTUQHtvHIYv8X+
jKTnZwLZDuCm/Z5uu1fAOuy1cUUuyqRhbcnAd6+EDjs44jveEWLuw/RdOf43tFqo
P5ZGoYP4dEUdbAT37OamngvX0GUFJOHxkhGmol8QC4Rtu5QfDUiIuVO0wrJPw2lJ
qn0r35F/cepOVTgC9skL2tqA4eC8V7bHi2GcTrqqvy8hJULW7Rx6aCl/xTwe498I
0wkog6IElW1WEYs+ErGWFjqvy55oDuME94+AY0EVTQRAb8ivK9y5g3nH2QdWfzSf
2iebLshbEbvQqNLjRhiGTt171P68sMybOM9iun3mF22w/dkyqeo4b4oRuS0hQrd8
TyQ83DyK03BL5/k66nnXJco6NtSYv0GQp+XxuakqzsXuM8W/ou3AGC8toZ9oW3U8
NopgEJreLiOvlsH6y2DsRDS8//gYCqOG1FLUwyWWM7paq7l4bYUfb5t0K+N9ZfAV
QsF12J/1uRcb9oiniwrO8yPZWqUQT6ruNQ+4f3bvAO5zSLcedzq9VI2fB/Y7BVrQ
+bRqOX7hJDD9pdiWGySdzPYklAL28P2VrEizJdXdIo5zgisy7fOGyVUczr9vJ3xW
rFzKdAsZVZRYUAJCrAE/JSUY9Gc++qahJ6xIrZ72/dbZQTT/NxNaILP9jKPNMtcO
NjXugXEjEnnkfvn+eupsKOaVO4q3TFEcIZ/5GL72EcFPgeJm9NGlXkv6OSlrdUx5
NM4wteyJcux1Wcrm4azJ4Z5XXVs0CO6w4e0JO8P6offBleKj4vZWDNY13N1S5Hrx
rWBTdIRLbO+vduRmZNNYAO2eIEKi3+8PHCuR32rUZuqhNmecUomqPPBqEzrKbdUt
mzBET1Q3CulJNzKhgAiIQ1dY2FcTx/l1r09ByGTN61HSB+DCQ2XECaXdgIu8r9zH
MPVXJBFt2zxaqdJE4X0EspJLoyQg9zQSaxhPQNOOCWdW5Y5uSwTTk4SHXRT8wU9t
SqCE4thchhMoTQLzVH/UFxG3WNBFNFS0w4WRKoCI80b0MXwZhhFoIytVJ5hgwaA7
em1Q3+Il9UlMZD20hez2r9YAioFE2A8EsiU7PKSPFGRapLq/ZQUVhQ4MOjo2N7Jc
zaGpOJylGbYkJweFsXQZA8ydZ3hVpE6R8Oh37DABiqhzu+Jmyop0deP33dXbbvo9
q61E8ROka4AFV1mHxnrBc3gs3AMaHDNEv2eEB9V3EDZNyCJSeo3KxfAYdGWvoo2Z
JdlOegMpKoArxVwr0wmiBkhfRpPm/uY079ZGmpZNPWY3xbeeAo9gxUxJu5Edm9/N
1L1k56rQI7lK01Wf3dLK0djOSxWQV/Gp2RWVG0MWh+U0fr7MK4w3YXwTy/ygSrni
dbx8J3neBLGImbq50j+gOWsL46nSkt62/xTkwO7mchRuzkwT9k7V3Q1HNwf+XRUn
5rO0CAFZFfU3WWBBt7TUOJyC1LFIGg9G3Q/5gkRd7sYf7/euYrThFxU/gJrGhn+C
d21bUj4CmWyzANSiCtMUrgyeWHfnaXBjzcl2Oibiz5Wh1fuxT1QEWmTfEPsOilk2
ntk2hwQ2sKTw4xpOSwrfwgfEQSFlnuinxmXqflOthnWyupqmo9bRn7sIU3sF8bwo
5MF8wegD1ssweTVJVIXzPXcELkxRilPDDhYQWQaByQYBbyV12bjkhc9DXHTxSJkh
52NR/P8oxOc3ucvGcxwWGiyU+fHkp/2bBG4Ggkdm4z/GFA7TIjtkbg6cIE0w4dF9
uvOAPtVPDU7QbSEXSikuOSNVaxzb0UWBr2Qmw7ykv4gqyAW53Hm877EM6cUVHJiW
wMxwz0v3XyNww6koJwpIyfnK0H/kOliVyyf3IsGl5eRQYi5Bog0Sn+Z2AtAb6NGp
cCIzn3nZ4Xiz8hJSpB45ygajYbT14jO53pUuVnEcqd1gG8/8jKZRA6T1L3Y+wLQn
5omsTm7k9Bopy2ZhNCn6XXNr4UYbax3FhyQPGC914lSujtpTZk+fcBpH7mzwCSoF
K7969/UhA8RnUd6ytOC7dwMGVI6WA3h4G4LmsN+3tektfwPZBQ7azK93tY38ii9l
cESwih26z5Ql6FLUCBLxeE0MwIabdU4xOIX7JSLz57/TPDmfJPNj+d8A3GQnGRpi
rJPf5Ptk4zLbWhUymPVl+hDQFcHLfXE482ZCT5zpsoaGNoOG7as5SuFBBJucuwc3
1TYV1HID9ABrtm2t+AwvYymPL/ggIsZoqO544qR90qN11/sxYXBH+3ywoNy3x0P3
d/e4kOfb1sgmS6R4lWtEbPNI9uStqyTFs9SohDO06UBeKz640G4owcbh/5RbZ9VW
dv1505iphO4mEIj7Ux204tlXYXkzx4pdvHxstz3SYP563+nwReW3pX9GR4SW2yR8
cT640NIc3D4X8pJFqvpipId0rAT9eqDgaTwmPH8IPnhm1HIQtP0soy8kd2FVJ4T7
MBKUZnIwm6Vea9s8QWoSJfIqHcokWsuCpvFdAPAgwpT8N7elkcAPQ8IO2+6T7JW+
ZBLNcmrjSkR8+cDCWtU5+66uTKnZn5+cMTlvUKESphDxo8qZgSgVyATxxtDivnuc
24mYV+g89hbQuLQxo5EYymICogsm5dQhJ2dvo6S8LWqFi5rgC6CYUAVbIISJui3I
JlBxFMzK5tm2PBGic+m1df5vX1cpFFEOoq0wCIUw2qQit1/WZ8uWOG3lo0BkpSpZ
3twXrVLYMC0sQlla/fDoYHUQAUpLYTYYuJ4asoXFkZr8XmXMdLd56sDX/PVaN/bG
n1uZ5zuphXE0miN5v6ez8+Ao79SOt6Jhogy+TEKnpREsCPiIU+utKzBGZ77D7CwY
GkGF1Par6yNp2iFSMsodfM9qCputeqwskIDgJT+fT4kBcIYxwwD16vxQF2HxBpbw
tEBhkytkR8I8m9/sX0NxmQIpwGWaOASIzDbt0lrKYxySPvPmMwCRIE28+tldvI0/
KJLdQibjHdCxIMRiKZFjSl3plvz91HyHUK9cwwQor4r4gYQH+Hdum1U8YOfLJ0PA
RPRl0ROVfkG8XobsyHYE5ire9QJGma/FBzF9jTYpTDO7gVg6/Wkmc1LyKXublyxV
/m+aCAQPnZB6aQrZrdM35EbpJ+gIHkpyefG0H0npLaqyxDEuto9I8kywV2QZlykH
OK0s6/y39slMn6h1TiCifXhjOx1+ahyVvSAViEzbpsZojXM4CLMNTKilQTBEFXft
MDwjfMMcbm1bTaQ0bElyLeK+ABn5Wr8QYoyBzyCap5im9M/unpYBmFr8O3hDRtIX
4P/Ltz931v5vKDSi39v6PdSdAPvWWeHwjHxMW1QLDEtathcHkJpm1iSzY5gLT63H
eTxl6+6VSi/fOBwrXOvSWVG22MCB/q9ofAW5iFYqhZQs0I5nGn0TzsJ/Bk4Ah5fk
SmvtcHnRYCy4n5y3R5yezIF9be2R3Pw/RoTJEqCmD5/CrWCdEWymrw6VBTxg28TH
4M4ZMzg7qvnCAFTGVJvh2qjAuohtUdZKunBuR2G5TfnC3orjerbfNhCkdOb9Oufj
SmkxWW8HbHzqUu+2ZudN5YF88op+TPDi7mtGs0STmEJdtLzJyB5jXtLPwsk0eSV2
ABZkBgHQU2EcufCve0VuDHpm1y/LKd/zhPOspFigYDUGxratY8mD2Z/z9g8U1nsL
bBUS/TmOtw1qWh9PBN4pbugxNgt7rOo95ZJaBpmHn1HWQpq9fPtf8L/5Qwm0axgT
qWSEGOWWBk8yj+tnn21TmltJN88aeOnKYf8Sx4Hsn1xbwPQfylfcjoiOyZm7vuov
L/M1S0JuGJ2S8iOh7PY3ZBb+S2S7TNiS/Qw9u2Fvcmp/SqBF8cE6Pi5vkOd4gQMH
YeYar0RcyFdR07FvYvTg5AEzD8pa+DRFmHrEZpOsZ2oLJ+yQwJbC8xhto61dA29G
bsXhnDTIBQch0M+r/mKak5HR4h9prnueO9baofDUaXVA4rXZtNNbdWl+6y7k81xE
dZoHrhKhS0v2TAode3MDVpyiuv6B7NPCL6rMkCjOmpSnpmH3IDQfPi2dK7a6nf02
fRp/iDv4XSsyGrkiMTNGPDuOnm3cen1LuxxVzODVW5AZ6XScIi9eyUtEaqMMxl8H
cwPod3G+xBW7vI2efmV7SP4huGYoLR+kx5V4FAtboakXO+7AOppKrig933WQCUO/
qNrEyLJJtvLpN2bCyNfcWSW8VukdZwpVZoK2eqdkyzEnDouwzJ9cYJv1cLilevSE
xgtbhe/hOu+uJbY5fO3+eKgSLes1D7tF4+iHzOHh/t1bFE5rGbrKLIcPfBbRwErL
xOQ8YY67P123YsWwAJ3ldZ6XRVkEau6KiiVDR2TWxwSaV3Y4dBWZ2zLfFSx67aNU
rl50HiXRcyPa1yeQyEWJp5jnyCrZKBQOjmYxpuRrUUwE8fC7tMD6lOj0N+UPXfMP
xe08FNMj/ZBQ0Lk4Hm3I6yhPTTRo8bpwsYYINuVVgzBbw1KZV0GamZK1fNbskei/
9EeVU4/eaYsgoylgvuH5b/iSh2MdkFB3pYBBgLYtsMJH9tKLqNvM6OdCbxs6o/CF
8ANsgDAQb/Z12367qcJH5shUDnsjdr+HVLHNdIbqzvEiEQi/5qT4sQ7WjjmqkS2I
d5/btj2ZjabAwQY2PYWr4fjcSxvOnSis411jIFNVbPnjTo3jS4qN1qWfjcMRdmzC
N5KqFytbU00oJwAeC6zfP5QuQDMiQYYagbru+YCR4mhWxC4KdX441TwYP1xgGOxs
9eqoguoBjn0sHqQ1EJMjBR7ycYm9aEwH9AzwLjxI6QnoBgx6VGZjcHKkwslSsjrH
nyDiBX3u83Wkmm8z4VzYmdfQ1aSsys81ml1bwaky86dxTqb7UOPv5WnjeM7jQKQy
AT/+rWFK5ZjVBgEe4bOe6BrV3RbLxxR5UTnD3gVfjUlPSl16HdiaSAEuZxTrgTNu
vSmXyjUQEQlCae93UI5RrHsdAdKww7ry5hlbdqDQT5Lv+3jK3a/5at9mYOB3aPAL
9BUS0VrErJu4sElKsvYmSamrNa5r+jo8teooTGsm3pT0EunMLx+ZK1vVD60MREZj
LLx90wrBwcvEyQHtojec5xBwY5wokt04WC8iTSoRU+MhppLSfx+eaRbZJspHMv/+
5TzWnDfphKqxYvdP6ndOdxW0169RlAtIfclToB820LYXIZB1GTrrNa8C079W9RK+
xhBJtdqCS91YLuXolMpOu3R+HRPHMOq+szAY9PRZhI7CuA2vTXPSCMbou070QYhE
I0ik/1gl4mXz/G2ajGJRJAANAFXGOybefLAdS/VLTzJO2rWCUeGd3wo6s4JVwvkY
vXWK787MMA/Oczn6ZSvne7Nw6NBQtK0JLOjl7vFPtYkBZKYrajv67SzD4/W0JBy0
tGCztXgt8C82Rs50qLDjFZodzgN7C/Vb9RvgcZ9zEg7kPDYeM/W8LsOmHC7/R5lJ
zg80ZXpTOO8LXEIjsny9ZqYUfP1MSeM3MEpABt5tupAHcusYOTzKUeV+u5/zq9gL
LFQaawgRYmE1XLXO7ZTaU/I3vRB6mngoqjJn+02Q1YPMVZPpUppavww9e/nCySXP
fuOp56pGB49N8SEx9jWQe2zLfHRs0qLnvii25aoUCEh1TGOsLyYFbSlZuU4THI2q
c3FD79I92wwkdvf442Ouny6+QGLASgte7RH7v8uH6UuOKvwUewJutK7LCCkl9l3i
jKnb77B2E/aZSSzWyOZF7Ofx5sSKAU/N/nTxL8E4jUukKvkLtpAiW5DvrPizJm0y
7+pJ9dcRKeddZOp7HdxoPw0EsB2UoMgQg5/KJat/GbHNBCFnl+DG1/ZX7tRbb3t+
AmCmaVUjPwZqvtU9O1iM2O8NBYVXccbn/0VTYjW8/rSPXORUY5SSOJwAl3wrAQ4Z
RPn8FP4NwaMLDe1/1Of8OgeatK9LBWTY5vVI8WK65ue9dt8BGGVZYezRQ41FDhXR
s3/bsTYfGvUSM2X88YG8290Cdxz+VLRpjCmloBaa8gW7YAG/cyD7LQUjWruaQZSQ
YpzMkK6W78VyVDH54eK+yjRMTEACbu7lVmTB+EkLYpBykyvcAuNSpYuYEZRWCxFT
VzYsY/c5fTj9VrXCi1xQ1tzTZvGyXYKgMfofUvIRbPD2VCXHUaZfHfOe+K183Eaq
wIqBA0lVrkoAiqej5ftuCJBpJlGeB5r1vDUF/vGXksH7mKnE8F67K+mG1K9fsK4B
wP52yIYKgnjFCWbA6+4ixL5TKLuCvFFOSeL/ngbdAr7y8JxGoHnq5DIdDI6a/io8
9nIE/gEOpa37LtPDL7RqbnZbjqwvZUFDhdSoAjnHhNkyG0Wfb4LipxPRa3F6oRgZ
e2C15zwz/wS63oBJWlZNn06N0y0znEWcbKW1SYZTHSLbLx+NaMzLjY1gvW9RzIvI
moO8aBwQMNvOQirGv7bfL+2SscwqYZGSXzmix/3O5gNcBBYx57OpJtCYqWJnzt5b
5iN++C01AyQoLM4YnytRC5j9wu0b1KU7ogzLBLYpVmBoQOPu038Ul10gxOLYgthQ
f5VOxDVDsuPX1HRyB6ON+Fuo6Rw6qJFESTJINe1Vp4ARjYT9ZUYnee7U02A3nRcX
bprwIoKz0EPW+BQAdehWqNrM+VnWVRumBYWgxWCAxfrl9sFSYFWrsdE54igN153h
jz5UgJd9SvrslPmhwK32H0GjLdHKXErY/glMGQrbXHcQf8oHIzQv59Vc+R0ew5zz
007N0qVJb2sqajS5UUNTNG9cvbdiiNbisX1UgCjHjs0DDdu6ksHxGsfgVMAdjdij
2QKxW/v35SxMZ9J6gIEB5+mnAQXblkBsLFF6qLx11OM2gYTpF/tyHkCrmJ0v4Urr
GTxUNK623gALQbR8ChO6nM404caEo6feOjFuK00e93X77cFT4b7Cm5ovtjda99Dn
1VAGBYS8HuOnf1+XHjzHdl+Heuow6wajqq1vwbfTRFbQ1PBxLBQZRh8clkPi+Xbe
mk8eKkKXrkXADxqaQheJryJXV1XxvQrPbBpyBwpBxoo+h5OYlxAVXNdgTcIxG4ER
E8x4Whho7SK/3DhLPyJHm0mUxvZq8SAaODidR4qcQrS1TmkGztGU/Fsdg4nwuq2L
V0rAyZ5aAc0WT6hTC5Jx5MVygXOr4Je5W35vgAZKY3QrBfOKUMbbM/lptNaVxkT5
HETUthtpUPrgPZyfzVCoj3OlpqLdUlvy7TU9V1FC7/QtlIgC9T3nFKup5NOJ6FXj
yG3KTeE0/PqKPhwli55bUmxiFvIvjtfkIpiDoPzgh+OdGAtPch0l7XlQVX/MLiya
n/15O/z53Zxrx9xVz5yE8QhSkC4FttxF5I7dXrznq+dzINo1VUTamnmOy5Q/xeFZ
f8L5lb572VhvkfrArBoIywz0JVF2YxFLJPkTV5KskNpZZMte3ov6OF8TZLhWJnsq
UE3k2O2o5V1AYdjJx0XTRyUhnRT7WLS+NlQ1aEClAkVzr7KjQ554+Zf0mESRo2qN
PznG2Cz7T5YCSkcUzwUGcGaNt0YdtCWTQ5jjRUKAVOHbqob1Vrz/bog8lIE7dFpS
mjSV5OKV4hFUz27B0vi4uE/PqJf7MBtE52qrD8qs4g7Pw48OfHPGDp8pPkzDb894
7+gEZIogAwAFUuyTDgD2M2iquj9wisqrKP5pQo+xS91qbwc1Bso5M+qpz4bcOdMZ
4aWFkQH29oX8eEt6aFAG3oKeUoh5s8O6fJv7q3Jq9pGr4Ts1omw9RjmqFaxUMQgB
s+aMup1/PvKZiO81quG1R7JPnmIUQvEXFZ/0TzZA8HFiYSwTkEz2du6GJMSAXIO+
kqktEJc8epR5yelTAzW35PtogJMQkXd/edtbbmx+aAO95fOiP7f8BESU+2tekUPV
tbcuad0wF3ou+Oi0n0YkR3t97UKa5ktvPaB0GPFGjHAc0x9v507vRdfy9oDA6P7z
BsIIW2stJHxXsNdbTapDB7+EvIrGp5apQ2AorFPfst0CSRd9oSn2sBkmKf69YMJB
TUk7UTY1uhBAF1km7ofvkFZaCSF+QL+nnwuBNaHDiTWvpvxvF+7USFP642wSKp5I
zU7mY7Suj/hW7KdS/1jIwPL8T6UoV4KMbHfplsR9KuJPBimMFWas/ULB96SNzZjc
IvpsBWuO1K0zJV8Hrr5lvrJKb1ENWwOqWgqChGq8mx5GmI/Jb6lhLU4Lfk9S1w1u
adNVmWq1a5Z+/HPJeW3gsabm4Q39zoLgtA+hac0j4jL50jh90w9TYVLp98Ha8W3y
3W1Me48FaZKvVZk72B7dzxiCMP3YOSoS0ZkSxT22h1fdAMTQ0WCzSkaK/NMxFRUi
ucUQTA/13qaW1Hx6tgOdGOyr0XaGAzktXpc9J2MVaGjHr2R80TYimG/bHqUsQfgo
noW4zykONU5bau/wvMr784Nomb/P3nrp5NAmgLevT0yU9NMmmkdFtnI0zV3jLXQg
j/XzJCOvlU49Zso0fJj00ROcOQMkQwTiaBjuVmxojv0saPKx51/vJShoqDk0mKX+
2vyUhDOAoDBlwPlMp79cunKOeVAQsGJ+YOgme1/o5MY/ZMd4ksPnR/jXSvesMZZm
6JFR+pkawFV9+uhIe3hQ5+uCswwBVmIDNwcbsJL1W/dIXANYxFhF1PsVGGQ3iKjR
/lhC/MPrTbyRf5l9IWup07LKEjIlQih2g0yEpLj2XxCnTN442Ivi1Ho925oD4khJ
To0ihTAgVFNCeF3fpsYQRAdgo5g1YsKkotJknFlIDwJ3Uxpfj5byzwCY17P0OHAJ
eMdiJsUsNmJpBLEU+nWxdU2NYJe9WdPybJZoXivZmbbM6NCqr0eVbqiRA2YWu21T
P5AferCv9Ni5MC32sJBgjFnUnnWqp2uJhUIFWnL9KYV+vRukzpxEiHhvtaDCE+Qa
Zp1v1AXDDUCBLtunsfBqPsBBlTfbRNrvDWsbuK2D5N09zXj5wXxjZL1IiM5XpHMS
ys0kNRWCZJAqUijLgoZMpuPz5HU1Rccc25ayRLz/zAH5w6mqsCehvPsIQmsJXC01
q93of3Hw6Gifv8IsHObSzZWSjotd2XKhQH3bnAzylCsEJ1dQqpULkbHmcGhRdqfB
4d0xWwXlPxnvlkxh2ZdkT4teUR6nEBFD6fTq9hum/itrKlDC1VTLg4wcALZMRUm+
BerKiqOtM1CKq9s28v6SQnf7Tphzl1vLPruP3qiT6iMMck5cQ1OZVEBQwAr5VVrq
nLq+J3b/BH7MYBwdEpV/YBzIXI5TJPyWlkSHqJSWjbPqroopZSDx3XnFGjj5kOMe
R1lKSKiT+JiqcjOu73HgY/KAfEevbZwvJ83bEqVKVG4M+I6gDjmLZqRc4fv/qqUw
v3pMWU2X9OBqz8kwJTkYU05gcpu9DHJ5QAjcWxuOWIyQDPR2sUA90Sej0GJ46GhF
6DwK4hA0oL4hjNUzezKXqDa/D6chR6Ydt8SKheAjea5LXE/3PXxHERUNUOfgAZz6
M7yvGnf4t1IcDh+GGjHp0Rh28iqVAMiU0z8p2cjzdk6EUJwHtJiD26sZaSFSmPJ5
K/kaUdbIMzuJUGLLoyj4JlCw5qrUO/HyMX0eBOUiFxJ2Z2btCC0Hoee9nzTRFv4n
xGJGPX6oKoE0CUBCKF1XGn2xuxnMQaruQoGH4J77UddnjQFvUyQGihGIJy4aZaJq
UeY6bJIpnj/drlW/HajWHRVbqhNsx3g4jXW7z3eygA/k83X6ngpwi0iVyspN6M0U
SuGfkDYb13dRKPsSB9t6jLd46OV5W3Z/x+YEyxuHEx0d3t0vPkNr5H8V1p57R97z
mFYxc+aC9sA4jbZtWQLNC+CQ6xiMhC47ZUK4Tj06+PUP3JK/Lu0NOvQmwRYtw8sM
IzkUn3YbQd1WcFAPH1EiTSgecQ3C+TI6OEcXgwlxcQ/1Nxze2Va76piUSqHkc4/k
vW1PIS7uOO2GW3Nnxmkn0XbPdfKajbYpHciHhJmXaRQ4quInJGJw74fx7Mqcbvku
4OzSemMKm+8BkFHByLQZn62VD/L8DLeIllSWJ4+Ml9Cg52MMScFbpIjcO3tSysio
jNnvcO9qDb8OFK+cLR4Xj8vhwaIoM2pq25Gx5nKsONnE60pT0RSHhJX9J4zKnwdN
mx1VbWdmcyoP1GnPldpHl3ApS8sYNIaZZQ6gVHD+WDF9x17aarGDNA/RzLy6DWNm
p7fhlJxjDtZoPVe+n3vkilTbr5hLqnCC26TLTcbpyuTFtETd7w/pzAHU0y0ntpPH
cjnWLfpTXIXOJtZr/wyRJA4j7fcNUt8+mptZ+driupLVGqzMRTMNTybjh0yvb7w9
VMMDnqx0iaN0ZrtIUrORvd7Zcl5zk/zTDCgdWC+I2ulE4+P+3rTZq9FUZN5a+w89
/T4GR6m5EYMZTLvzep3rqjxVSWi3c2DKnSnakipkozijoPrn7OHKiuYUQMPKQeqX
63zTGMVISgO18ZspBwIU6KtJKtNLGNEzn5thiIemZhegQTGEB6t5KNMAvvHkvG2P
S8d0q14vEQ+kONhjV+YeSQlTWf+W2voDEQqNA28MEcmpcaCCordCg1qjFXekXpvI
cuHBQY887256FrzIYAx/0ZPUpxhhoydYSXGPcWF+i3q0PraLwgH/49yU4bPFAVFr
6lb3zR3txTfqNlgBp3mzrKKR+p6bccuy2udHKb50gK+2YNX56zpZE0w6dszp/uSl
MKKcDPK1qxrMLT4n1yv+82YkYEh4V1e/HHwfKX4yifylp7S5uC2Ei/9JMH3FJGFs
7kmfox50K1pKXg17sOpnnpVUSQsgHcuEZ+BNnfzdasmdAv8qF/I3Y722FsYAXwtM
NhBqDANqCH0ZYPmtUl3OnUeeJQpRwxvdGge9kRH/FL4A8AU48Ish2ovRpHO9TMkz
g//p4HHqwM05dMbsrFQkLmkXHAUKmr9w+qlgcl5IG0DH40VQ3YkAFzs/VDjWxTBc
vyOK37xDQgD+9478mOEKeW70JQIx/D/G/TtjQbU36KmjGHNazZc4+MFhnusCNOSY
c2cXynwh8B1AOfqIg/wOPiug8XMs7SODT7V4O9roJrSlOqI+DwUmpmJY+AcFenPT
0NTNN61uNto6Vn+ntbuu+mFZq4GrHiYSxS22zGWMJ37MukKnfKM5wnOA3Hv0ED/z
FcaG/t/LB7EG0X5aiomZUBjIOCL5Mqa/qiBRYnE8t+fE7eak13N3qMB2WPfjnFCO
9EDUWNxsJsLoT3Q9ZDWz4LwKzrrjE2NV/PqApQ9qHIXWnuERVMkQaesabik0QgYu
iYPm1KweyhSpm2/qiS0wd+r+MjtHhUf5EcX41i3Xqo+uq3jQUn0ChjOvPWbx2X4b
KMTUR/Q9SUSXXYTz0VpRMPCZNfNNUPL45fhUCJ854WWd2pgDFGJSwCmTrjx/wB5E
nCABrBHdPLToY6dnudEV5C8pNR7He3+MTI6mnVnX5PGzN6hJ+fWmxQPAiJ0g7JJ3
YiaN6+wVA05Lk7wRa8LigJvZ88n8oRUcLQ/c9KjNWi1wDFTrDwhQBderHsHZjQ//
uds7/YxmSx5HUn81FofN+iCjDD07GEvNN5IzBh8Ua5x4xuwxZtWZPkbwnSeaLhPV
MZdCqa4x36HcjbhRfniQ0WvNDbznl0F9euo6wghqugwIgOUoN0pDtKxvIU1ZqQNl
JxtQn/58QE6fnBy7XyJKPQ8XZWSvzXKkYUfJAadUS6Mar47qGf7I+69Mn5WfA1zO
AFzQgk30DqRGTBCE7Aot8AsrdRL98pZS9iV9WsWHS7u0yfIBSn3xIc5T7YldlQI9
pt67mQD6kDoqkGQ02Y5E7WCLBm8kDGDjNqo5QvCz5N5PnqyYghnexFpCaUaMPNdL
+PTMHwEkux9V0eqPVPFsXMHz/IHq1BoMtTI91Z3T+/ybU99FiTwa1ytTno3/my7J
S72NAawTn0CMbfPUkqPbxObFqO+4c5ExcWhS5zJPQ5tMgkHC1vkW8yDgdUDz+Ktj
zYkd7sUYz+M5KW9J6Fzrsa/jK/2nMh1j+Xa3htzUubL7EJiE4XHj0U5HuXXpxGI5
WqNHn9WF/bUyP9t3yrCNlKxKSVtcHCLVfl95C45CG4xt6T31pazzHVOYbMvotKcR
Utwm29xpqZPYpqsXIA5+jZj5esVEcum/wuMDCrkaeCCQKn8WN5bEHS0Wsq6vEKm2
qYt0a7WQp12cpw/qIMKDmYdrKi9psADvutlPgZTWuOn0K8qLRNBc7+hesaKP+y8g
HDQzOBEI1ds72dmzdlO+/wPa/Mk8+UAY3mWLM64yyOtsXHYwbGZJ9ua4nlqzGMSH
wNNBe/oBUX8heu9VeAH1yiIOM4Axa0+DoKxC2NlF1T1DY9fcaJnhRj0jOmLmePr2
w+VhQS9RFwKH3ZXYclgn23jE8sQWuyjScJAcne9U3y4+CaE5SSrGQ5JpuDNeJGn/
3wOL+9uCShACuA6PMTA7F0JcxM0RjbPvmfBZoBxvXp7I49nu/Ymlmb5oOPE3RnjB
6jIPAdIs0tMxuvWksmmzAjgguQe4g83GzNgC12sAMJ1o+6wEtqgZbx13ssbP5CS4
B8cbqsW5A+iDAFpd1ZTc0uQDOgxke/ae179guSRms/atQyXiQbo8fSHV7f6XIYII
kNLaEyDowO79UN5c98T5vpFtLZdyFeHoGyGo9B4QjpUS5jgdPd94/1SGrYsmCO4s
mvKgTFM+hWNBVgAa2Lr/kf9yoq21BeIOUpZxSDBKiWOZMSrjzoD8egGSLRoXtaQr
jhBPeTI19n3M0pYUAMaLbE5lU9tHzea/0qw1MHk4MBVY3uBK2tDPMrLJ5ESR21iE
FRjb/dkWjUwFVhkS27ZrCVarw3vXOkBsatub/mjJD8at//jhRovnq13UkI6wlasY
lZlJkdo37F4PISkar7RnArpR/v31gopgkvgm7m97SsK/lnguFFx4on3ZpJiikaG0
w461tqRTRDVdIOKBTlpONYs2ru/3c5rkPGAFkr9gRvkEUoNqfLD4JfWeLWB4yRhB
dLpWdEKEpT4nUOV8Bu/+HJ0ykT+fj/pcbTROFX+vmfyF46dQatwrjobKBxWv366C
UBnvn49LHScUlttj9s4Im4GzvqmL1FcKAGn83iSLwfauCJ0yXFReu4TJ9jLS71na
GTqKcr0f9PAvFKjiemGAW9Mqu594KDfcr3gsHKGorI96w97a1WnDXdoUSr3W/E+4
OSUyewtZDG3ExU1Pe+vn22hqYftMb370qszYZf/oMEOBQq99VPK4RpZDUAN0PQ+6
ZBeAf/ks9YR0Weik7FEmN1cfo27wg1dBSW5sDEImN8jnMaTpRT3lKKOzOPiuwMHK
IDcP3SGZhpRhIFtKFfHE04aWNP37QN6hrzJ/R6EciGKCYtBWlg2GATToERU6EUhb
5qLmCQPTUG9VgH9BvXaqDV+TY2oAcnYu1nDHT13jT89dcoxILVsavd0Mh44oYUgJ
oIcWNtSE8xhnUNGXEpzcU+Ac7NWqhDzYSO4OQnw4sCFngCOsf7q0mY+KwDkvXIQA
hw5FAmHC8XnuFqgX55sJdrYT8tmICMKAvPhZ2lr+n67T1plWc49TIZW4ZbvZ0pXT
8sPoDUGhoWuh0LTWz8XopWfp3YDgvwQF14+yUnns+jFLwGfFSISIFRAnXujGIXSp
c9xro2JsT5QXtE5xhoe7oHgm35p/hFAmkGgdxnoKJzsxyOACQ2rke1Fr+lGrtMiN
erdL16/seKOcOFognGilq3qgoL+HXmnK4iTzgrNcBzJqinW4BEyUbkAAI9KHKn+E
fEVShMCcewUGINqbgT8+w96PGu/AOKMSnHLS3TpzzfTctaYPDRun1o3Kl/V2xWsK
xAIma4aKriO4Av+rNfygGl4rGQXOTGnpzvZfn8AYP5DJ3AG5/B/+38KS2QZrNeme
ZnDe9Z4JLPbhDc9hOUKOSII/mzCil1D87SGxXpNMn6ZapUujDr3nEaGm7aD92g3A
EYHhvnNaANTKf06iwMkQBxg35zHEdwUZMN/EcNyhwd2ZsM8zpIbG+P8ufAdPjlE/
BFC+GFoVk9xt5kThQ6INX/uxNnCbS2xjx1rCQAK79WfcyUB5WyXG+3szABVEA1h3
VYHYrotNOiJ0B+LHzlZOP5hbbOGl9T6ZCxCi1HczOgG+TLDHcZpkmB4Q9AFRvtkm
2TtBCFf15CxuieVf7xSKT+Z3zHFnKxNcSFcASpdgzXUPfT2pO01uIgAvs2Ky3Oae
qI9aNu68inSx4Waox/YRJkDeA2/mCNd1zPjR69fV/sQ55HN1wsL2qkcIShx0CAwp
8XaJgDmXdeoh7AiHP9HBEvpRtEl4Doyr/vzOg0tz01xgA4WBkJeWjsfSpMFvTdv2
gG7nkw8kVuJcFq7CGsos4rkywoJQTyDofnweuaB2IDu8xse88P2OZlgzseaypmu0
WRWcAyifdIBSzl6brNFV8DxBTuXVwGhN2hxQmyvsbP2eLWXw9PWEqwcCh/hHRT+a
/HVC8InCdiW+LvOvAGArTQXNnACFsnI533Q+3DNROfDEuRhSroJoleMEhNmIpOiH
npWQrHB1I3u2lphh6mjbzeG2aKFMTcwyDevP5GLY/zPoit6yyfCNyDazemR4d5ON
Y4Qe+mjaye0ZFNa3YquqYoAOpcT7CjUd8bwmbfQlIeDXEMwA2KAIuQhydXMBxIPi
xwpYmyDVQJq72EBLR2FR273J7CdtqPyn2VKThSEefPfLBftT5T4zqt46zbkGKVEI
+n7Fmt7yx4iL0zoJZ6GCurh/DxMnyEHhh3aBuwbqERSOfdpYPU/KTavs+FdAujfN
KCKTOzaQkPp2wA8xc1Vqi56VUGw3sZw8T8M5tnSzgzYt8EbyEp5kssolIGyiHEJD
NTaUZn0nM7Y1nSaHXM8pTAB6+OO/8LUzQMXJ9T0WLojF/xiCx5/AxnQrTVeuxTDM
rSgQnYmW2BU2uMzi8JTlK0xR9LqPPLcmU9fOeXJthcoEtK1cZn+MeoY/AHPFWYpu
Mt98t3BZ9ZJWdqQfl+kTMokkLc3pYw0HWDkBcUwaEyl/yX+0y+TiSG6X6IQH8rDS
g0McqtPVo1G4UhQqo52fhIf3incxNMWQHp0PV9V8hWtl70FvhU2Ry/PVwy2cTfHj
/EvsvoyuaI8RhOHrOC/IYUQMtWnl1D7zyesjKRE2u5RTYodkPquE7mxtFhNiB6NK
UWOwlQHij8ycvWxI6VyjmdumP8dRfP0eHHm/R+6jbu/58lWTMHoAG2NfJ6T9ZAJl
0eiZASFRvtR8wrxVKnvITGqUU3CoIEWGQ9Bp6jzYTPf/jjxjnjRydrSIk72v5qqg
t5yP9aIqrzV3cX8WqfSRnHU9el0/zJuhBN0LSLGyMci8ap01Z1Joy+MkGJ42TiwH
hITwrVaKrq0zn3MTHP/AbqIqA26p356QFfHeps8Fs+YlhQTnhuc9M0reT7psPNla
k0UhgFl7bqwbXnjdLG0iR9mhACFuvZ61JSA8N8jYKaVQOhKxnx39XynfgU020iZW
uWOCVNdJNS+Zqij72mjQbkJY0sUoEt3dfZRjAVRu3kUdgQB+u1zbGE+SQBvrN3qX
Sv0Nd5q8zrJA3D08GJVceQ6R48UxSCHLcKmkqDoW+FYwyTA9zm4iEjCKLz+K1/T9
XUHQkVUQ1PUswGRh9zEp6f46bohfAZsMT+16qPvS9+aJ/nUTO8Budt/ZAD2aouRO
GWRWOyAzWgvGG8bupYXOu7o6DMTvnFDIzWvGA574G0Gp1gzdxcpUfER8qpxLdd+L
GqAPEfa4O5zdjPwn8dVtq6Cm/nRYTtC6tekmEF8VzYpXlsANhmwuWrYLYTgdWdQV
SAyBFpZhnJWpzRYV1kEe81zs3eiVNjIOGhwe5GGvuDvjmZORRorrXBYYKYu/QTLx
i7U3VooQ87ni2hOlkaSu3f4mapdpFqA+54LJ67vBmEjZzWuwmkYKQiAdpOigRfcG
eOmiq/tJfHrYvQhQ06dEZbvuEWDSzIVcPnBALrc3FzwSHVbM6pMmbPflFiYiBOF/
anh2HkzbAMz8at/zOgSHHxKSVqobR3iLWq0JFPRspeVUyYbfnKW4CGlNzBKVdQEQ
asoEM9+Wyz+oqu6FpYcwIfO7JkzQnpSeRbhPI/73hNMPQCPiTDzQ+zxxnsIcjDYd
YNV+3cZIARH45zryHktwEpk6Na2NVixiLIJky3VmukcLI/ROOFSL7TX8yF9aGFdW
hAtdd0PbeBAWjD4qya8rNFPPYqR1xE7gaJp4eSYCGPHNAKudeRU7mu7++yVlDBPx
ug4LgFec9eKy1TjHErM4ULJ9OmdER6fs4X5wBPkQFYW66NC9FFkfZCj6Er/xPZfx
RqqSbvrPsBf6iRw8sPGqQ9YbwNgPkS/I2X8yvdl/b3SKHxZ87xkohJPElTBbnHA2
7PXVN4uB9nW2wjutk3kbpW7gpEsdmtUm2BhVb0OpiXBLhjOEee+EGJtecVCeLQT3
l8jtkdxBl915zH8fe6mA7xD4fXNY6NQjmZjpnTKjYoUr6Gf2q34DV8uPr9dNeL3O
CcuBLrFskw4X0L/6p3vw4siGAElNwheZa1tapOG00iaU12EnU0/8y6Wple9ky1sv
vvpzk1fISwyXBaeyrxLDVvI+7BVcnx7TO24UEPO4a9Eed+kyOVGDQX/B7IQA1vxa
tw86FbRArMAdeQnOn3hL3w97hfv8r3fes189J2yOn3ibzuu0z13KjikeRJmoVkKG
qhzdLscua6fd/ganCND9p4z8E37T0agwpWWb46Cjm3R187I4lYhCRQ0jqkqhATWa
WXPPIy5HqBClQxT0E8dypHtoI1rz2QfVfbC9piVRh/Enl0iNTKXtZJUKKje1YW1i
V2AapnJXO/EQBSqRGNOXFdH77m2sunvcZG+JJ2uEcBGAhP9Z3OzFB2ygi5H105IZ
CjFWU1QvmOSZ9V77bmpVRN19ePFH3XSey4ZMtvAdNhzRSOQ4lkcA7+iqduZzUytu
wPBCdFvIt3Uvh9GO1YDE+kaT9w5w9qfCFh+psp7qAGxn9+pnKfy0cIcwK0BTLrKQ
lgTFGPFj77FyZStVcyZKT/WGPuo2Mrm7pF2tgGnI9LEqx0YUnd8J1D2IQTk5pKdz
VYm3GHLsCZyz8XS0rtr0Si9tjqZLMja+t9Q63DO2jWv+FTJRhyJzEjUG3rtx/NqI
4McKgAT66zoLy7aGACut6qFKNWFpUZn0J4y2a2N76W+JREOzptbTyTguWZCv02zB
mtQAQ1uwh1LPesQGtFeIU6VE4+uRmuBzRMwSJ3Wg+ZhwV2Gwq4+sjDI8U1+iuap4
/9ctoqrtMC9hEFP107o4hRWIwNZ8vNl3XbN8hhn6bDnz0EH5ll0aFCI2+tSkWcjb
7B1r5ldvx/kHAHBqS1ZtFasIeybAr0CZp4Wdo55osAMuorC86Q6frxaEdDavNbGk
s0quz6O9AddkT9IESojIvOqFeC81JGma8iwtNE9nQMzHvZ6pwqvbyuUTFELa00eT
C7ssEwJvRux3X4BiTxIXxZO+yl5KC89mCKMtTHIo1IbAcnBsQpZLsvoCLqUX7f2N
PvP2+7Fre7CkjzaQSSIj9dtAbp+PajqLlSqv3lLkCCz83xWhLqZUZsp35siPkjGT
1RLH16Bqy1arqMgtB1kRUYCYePbj+JLU2CfeuyC/WN5hE++icnCEgPIy0QX206i2
PtA84npImAOy4opgcTDhB76pq5ZpS/9hWKkvVKFdFxaDAI9MxMJs8AN7SRmE4Hq1
Wj63VofaNOy7klNlpTosOirghxX7EXFQ5ZZirLkVdX/3GSUylVMD1kxyDNgT51+C
AbybVrm1hgU+2LwCeF0qgiNWxbXeBH3Ty2BCWSaAreLunIKNkEWYXgs+FKJQAGiE
PtJKF99P9R6ONy4G6P3E87+T/j+NCYImG0ZpqL8CAz6rq0+2AScp/XANJk6kYw2f
IlxvfMN23l0L5GIvP+u/dLEo/Wo7lpkmQqDqpCyXEU/3+S3fKfgd/PAi0dcUmrZV
zln6tRqthl3zmq835c+hOu0CSxAJH7kU1j2HG9JNSrQM+0ur3fQmNFxdkNyApGNm
1VIJ4heUc3MwIlPHQsnm1UXL3gEB3Eptp6EpmVmmuqhiPqony8qMSXB96TjCm1nw
9cU9kOH5wvvZkl0A9M8/z4iyUvmR94IExZku3ZgyamaM30RgarxI1lhnblvEdAh9
yXqyKNl3wlk3TmnxnBOoSwlPg4J9i/32oB2gtf2NsfhhGKdftCpD6pK/dwYMrG9/
uRURDGPIlTtA1xZN/kGZejyPm8Rm34/EW4SxhC74aWcDaRl9k0zKk+wa3OmFgNmu
oyLBgBfbGm1TlgEBDLhKfLi2tRB58biX/d8ECV2kCtUtyw8RhRAmZ6YVQrBHpYZx
Gm+mq8ptHRD/5EB7MLWDkrvH8xqDl1y2XhknMr42059ca/55KNxf4UChZQUHGSFS
Jk2HjnPN8bxz2gbCb788ALtzDp6UWgNrYPM70d4iysL2qUKzRWnL1GmzFG7Pbnu2
o5WvFu4cDh1aXMSsLauk0LOnLNyp6Ak18p97ewa1vvXjl2ehCDCEMKBjEolednBG
rKC6zDGry+TtD+JTH6P1RGHhEAciuX2NiM0xR9miVTPfVA9mbCyUZB3CDKX6AU3X
XNQEe7pCVCQ3y1JXhHMd7T/hMI1rUPfu8zbccBrlIjvLxcIX6IDx8sKIxvfdzUwh
uic1bm3GWI6UNruQJx/0HlIUDADlllPPxVV5XK4obbRCwt1S1QBMCvvqiJetkaPQ
reVtNIdXY+v58SAvv2yg2C3drxmKpuzezZGUkIWA3dejxh9WiQ1waiwtTwSkSere
kT/Xg9dZ75b5AEOMgPqt4geFSdpCXRi1fIG2z1D88xqn3WgY9aO3R8g35ZCH02kY
dM7ej0+oDdpwD4ysmP0OPRf0LUKB739jnbfCGIL8ACOWbRQWLTxm8dMYdUm+tuzT
2yA2w3RDBASGQ9IYB+2w/oK1gO4a8S7BqnfkfOQF+BPM3E3A+RT+gNCIMiixYSQK
kOxBfnsxFVQjcZF4TEE8Oq81Jd/RxnMdkjC/lXHJHt8Kx1JDxJHDS/RARjs/am+c
JXZg8pDQGgoVEsSkdmo7MshaZtRBlHx7Ml7R7ebs6bQNsr9Nw2KU0NZ6sgtK9xIK
FGmpXanhJVhLL8/bNUUflKAqBkK7mrUo/NjercNJg8EjIk7klBquzoS91n//C/0L
zLwTexVyP+HCSyUeQmq+J6c2/lReeLhnjAoTJs8vQJLCxGvUJEbfTEAnC/H1dZgt
SheqcCg4laObS/2nO7ksdo+jP2ZwNlTZtsLxC/jBpgqGrcXaaGCm+RQGad6LgRLU
Hmiw5AW+zHmoxRHr81fvHwff8pZfQdWFjjzRvgLVkYdn7JfPJuxJ5W+Q9UgSsk51
x6P/AMG/y6wlcLuFetZRM8BBKsTqS31VPqvrUZgFAYOPI/HIpo8QtVnZfLgyTm3D
07sV40pPThUMmxu3cY7IkK9HH3Z6PSA+IbDBROogX+Kh7Y08VkJK6XC27gUd6c+/
QNqsxtXfmp2TUHjJXELQjLv7om5N2PhpbjMaCJwI2GUdVABtAdClEjpYNrbWEvJZ
Fz8T6quJHVSog8YqleEy3C/fMe7AwGVoMx/AdLD1ProfdwzjQnSSyWqcgySRz6xj
qzl1yK2V3DS8Xtni+er/RyWmr/YZ6OFd0t9oeQJY13rBPkLmMktkoe8b7h6dwpjW
rR746Db9tEY6zgEQ9O99FgiHazQqL+e5h/j7PRO5yfOWR+jep2Z0n+PusmjzLCP4
kcEbAH+HOY+LehKfr8BsNa3FiUVEYqMeqa3hZcMHEspQw5v5vwrxl8jsDP7AG40R
zUhE4XxFVtseYavrJtYE/dClXD8Okqw61RvjlEimSxeG1wGFbVB6grSe0fBi/QoK
JoRIopEbtC7ZX45u6oXbhjukF5dRlQm8Pk4ax99wNew4Z3PY2h3e79JFOAeH86Ov
KMmLkV1HkaCJJLqCo4j2t6UcQVqDXF9aSqL946wFNvoT+bSXrL7zonIuuFilW/Rw
k7P7U0u8Nw2qv0AyuzqT/8ApbrTZuT7sjf8mzp+HQW5nw5e0/BW/mBjSm5gd4ZmB
i2Jg335tgqCbNv4byRl/H4bAp7/hbzxBpDlUAy2y/WnwTfHyb8QpE/tOejgD/tlI
W78ERmCpMRRubZ5Y79tBTY/0Y+VbtNlv+YyacyW50LiIj9X02OfLu0qQDLfHq7s4
AtLeoq+2hPsAT2zOn45Pl3yijTzBFx5OiXpZzRKqHMCYiK7OiRy6HXCR073DK8oF
tuTTw0n239vQyffWgJyA6BENPwsQewLSpXEIntdY1u5GFKF8GMXyvJ9WfuHZoDMY
T+02vgBEwmuh+ADEsjqazvoZwGGXJmqwRMqW1SSptpIxcvx+SDe/lj6PBhVoQbNe
6WZwgzh+5+Eg61yL9RoBEwnf9nDBvwOPZe94GkZxM1/P7lGLnoI3TBg8h6IyII83
iMDpbd4GB8Kai8QZRGdXTqtv+btSUDL1JQEUk3iPS3hFBnS82w6mUTOHXamu0apb
Kz1H7hZege0jw6eihjC8fpItvNL0v+ea+Kvf86fCethCzbIEoDiN9cP+868EXLB9
uw5MUaoWHjHObFNW8qQzIHnHOsBRx/aln62HK5qlOUUkp3T3jvGxovUKiHT45XqS
ulWv+cfxIaYeLzWRmRTpuV4UP0toF5KGLGgUBa4TjW0RwvWqKMY0ItuJ0DxW0gRI
bEBVZ6vqPg8fL9fd2QKWx89a4FOf9NCOJVBUGNsOG1bhjFn+k2RpB7LefJF3sfag
U3Of7wYRYJCLoWYNDQ9GQV1lIKiMCFVwCZqGiJB0WlvA/nmGGGwwmpV4mPP+2dp8
iScJYWXEvhJAdTPo+PDQ8cVQ0hXx5eQEz7zxPsl8p7TTDc7B3kCEbnbetw9feg7B
Hcd3QJJKuxu2a7YfO/tT8hMVJYyeD8E7AzUQalX8Z35zmruq21Y/4/KV8qFOsV+w
Myuk5J4cLozURqb+9mKSRaZrMWsWUTMEyThXwBgJFMrtpgbZ4X0+JTNprq5QA4Kh
wQKJgGvNF42zbl0U8kPV5Vj6IOXi2euNRDee7bqjQ/FjwR/y697i9w+iMow2ymCL
P7GXxW5kZdcAVyyNc0gHcNA6mdgpifgW5CA13/4us3h3ZWlXjI1+FD7yDjqQbTvi
mQRpKIcXF38V62sxywWp9LtUYG9Cq9dpT7r7SWl54rjOUd2NADy4217Vl2q8c+BR
bqz3qm1KqdmCUhSh7LXrLI+hnqMmlG++AJvzoiYL1trYrC5xUe2tzYcR/8EB/sLl
EfbXEDcnezL0L1Uyn7zMOfjA+u2twyYAGT/mWLgX0edX65STedbozo7j4fgHYu9D
MoOoX44GwhfIparZ5zD74msBJuc815b3uDif8swfjyGoSKf3bDC7lzssSjCwsbwN
6SVNPgJgCKZX91g6FdbVKrTeuA9RmUWDbSvpo2jqLEM6zgJR4npnjrZKA/73tK5n
BPA5cjwzJDJzIIGJVDvpSxhCPbVRQmYzZUXy5Ob+GEPXC0UVq0oQJuJw/RBiKUdX
wumfu6Xd47uJfbqDS1kB774wxTLAbA6uACmvgF7RmGAsa4ikzPcfGQYPYffdfcvp
QwvFAI5eBT15TVvqjBTPxsvnO/Pt6XK3QGmjlUZcOcpdn6C+LmQpTPwTYiUbCJK0
iRBoNgulwK5iRcR+Q/ydcTSiFfJkBgl2vw45TXCUbfdJGumesSbcPJealeBM1zpA
vFIL16PEJUZbVVjNQCvkW6fWtXWXTuf79rjg9O1BWPya/2j4sRvTBohEV2T0VaTD
GIIEYI5adm7C+gvACQSl/BnnPgSNPAudUWHZ183A7/Es0vTB+TNJVy5Nm5E1dmO+
Yax0SielC6mTgn0bKtZBYpvyQxQooX7y9RdisvP59gDOeEsSycQn1mlW572yEiRV
jFDbXKENvKDRu0wu/MSX6mS6xrqYsgxTRAbj361nLzvlNjtm2mVLZUn2RFQTanSe
t+nuyBuNItbbhbxxqmsKfrjjA2IFCCSkmiDLz/S7I6XiMR543EfgRAqTxSWw1J0J
IRzzKyNrx1faXL/2FNtQCW60iIGnzOnv5fJsZFfUmcBXvO/BaD54SniMpxZE1xTA
sfS60LkKQnUOq+wYajUEVzu4+FYDa35bHtOS+RH8olZgsdeZNY5bPv5nwQf2IyS6
PcDTdljczTmRmubJ5A9p085CzCErWBpNoHo1Bjpf+Ah2gCKNPDiCgaK3R1sPWTex
N99u0MgWwjHqHIw0FJ2VipkZNlu+3oXSKhF6bbHAFprhsjleVXrz9RWyFhVXDdbr
mGXY/DIaXMPFV90j2lV0q9BuN0vfrIlbTyun2xs6evxyOChBCr8OPld8A4clkE4Y
NeKK4ofXH3QY70Uk1PPeoiuGoGxGxAGa/shXAgfWjCrvCqnKBs0vcr90C9ppNhO3
Xi4ppBVTnE9nd5fxdOb6HswHhJ1r4lzc6azRGZmOSJbWz1MARQxicdRVOiqfuPA5
H42JTX4a3psix9bnTCV0HUhsKbp2XX2mI1FAnaydtlBR/7atYNTBWIWwWRBSnv5b
hM7qs2yc+kThcH5BdwKD1s/lOZyEkrD4naJj+mMP+4STOUVOkcOy12l7SA2KiKVa
1tfNo++Qot2NQ2wyLgErBC7h7RTOGPGaNRWAu7ISwTjoouGbfe+fEIP5ZuMMxiyI
6cv4ev5BgfAhXjeKIm+bm5acKwek7socfcSA4XKFyuAmaJ4yoNJ+HWPy9d+xfuYJ
EPcLRC2Ei4iLwTomfjwEAUki8rqtY+XJxD4xdwPfGIaoOp3jUr3Lz5penE7sDW9E
NbHybiwoFcV8XSChMwp3Z6WYh0QE+1aayZ7/pvmFlBhEhhFg4Bv9v06ws1ufcTku
+JhHeXZ+Y4fhXHR/pf/R4orssDOTTv8EwZoA1VPK7drUx+VC9NO0vtLRMas0TFTk
3Y23NHFFmY15KQSagchyg5Tw+ENKNsFIwB6d2vRkmPqFZWK//T3iyV6wKVrMx/Ho
Wll0UrQYSE9xIAdAE2ZSB6X+F482wf+JQYFaTnDZcuoqAUj35XT40Pn97FN/UkcM
47zOpypvRMCGUgQFl9n2bMeXvdqV1iled80bNcipjZg5iN2aDxxVYPD44fAOjtLU
5/48+CeV5IWY7FJf7FCV764UpVgPiDTaehcTNSS3lKHFFrts3cSSaVgc8wA0iy6z
rjqdtafiQwCGnxV5BjTyreKivOMtf4h6/AhYTcltRYja562XYJ5N3VewIhc/daH/
tWwcgEIiPKOSFEIrmG8Xq289q0kFxI0A2RoVhC/NIIehHE44cvAzsTTZXDMvqymQ
ynp8xjNJ8oK4dNJzjVRKwdd9CsLrbl8PA0CshmEnMr6msjTjM/KkY/fSGFW2vzKw
Wo0ZoT2xHgaFc5xeobJxxkXRdKEfiVMD/dKKyd9qEJLHDrEZ9GiIhenuleWOFQ9a
Tll/FIZ02gUCvuqOQToRgJf1FAi9U9GGP7a4++4p6iK8quR67wumSWtmVsfD/obW
6kl/PMstMGn07bXtzqIWnaTMOrE+f2o4q3UkUpybPNG/aK+uW+b+DzQnHHPyv6mX
1t//hV/ZGYMH4bkO1Ut1TVekrI0BRcrjiUrxYMacSjjfacy6TAD9gN3ptQromx8K
22dM3Wqa9PW2KglcolXBE+81D80hh1b8VoMHpkSHnYXArMu7tAqJzeU8j4M8+Vke
uC2E5w6gIs1HW4UW/XKcKyUrktSdmAA5AE6Tr7pLBnYrlF6tKStrTto1HFX80Gir
KvDAqfCMBWKbaoih6u6/0I18hm0Ef9o4abSr2lRJ+hNee1JvlFB0Sytl8R+NpBCy
Ys+1IKS50xO4Etr3lCY5ufl+OdPT/IKg0p0qcYJATa8J1bZ5u2D4IEgu1kw1+w6d
niBcXacUsiGQETznmHanMFyrkM4X88njfJVc8uhfgJ4uxgCG+KEaMMJfGQqzGqCv
PO0E/qYfUaB0xB63Bk4f9dDFsN9+DUK+x+aj4aZaLnbUETuxvwEykreEMBBwjgT8
JOvnv+39JaAfqUDq6I5daCkVLWPt4umK6xl6fEYMEklOFrmdPbNHiqs6ApelpmxQ
GtOxMPL+5fsDylz5qzqI+lUiSRuVUXGMn+3Ir19oFkKrjnmbGcVD7yXf6ggGymgz
xYGjuK7Ur4UyYgiYZieicURiEMwJ3sD1g4MczdjbqtjA8QLOkeH2en8slIO7eWru
Q/gQcCT9fccFqQs1prgYSopOa6o11dehPasDPOjsBeMSHMUdJPcC/RZIHikA1fdp
WTAqO5ncbCw9CSi+Kz7RUv/psWtfgleEugQG6skNfXSQhQzfiTEsYfCnbdFDrle0
ZHVkTT15dE23I0jcIJIkp/nKR0M11VKl+tjW2qhuu8RlwjcAc3bXFPmKU5OolBRy
y928YHoC7+/htr/quKTj0S/bf+3WjxVefoNULxNfHrAavwdnzRkXxezpVwbjHBHC
w1dlHwTlwe7bsCuPvAVAXr+mu2bEapyDt/0uo7afCZvEvBV2QsDj7tGeDcEyuoFc
AN8mvAGsWxSwkWeZhSppjmXBGezH/bDeq0+9JsQ44qI36JUBnC1OIUkQtCpWA5jp
+AnB4sGNKtjOlJa5bLCS8+8cdm2KEDr5BAVcR6KdFKS460C0qHdtx1UzCDGBt4Af
ErRvhGM9uTogeGl6brXXFD5PSdHK9SMGEpNBOvTBbNvppV2A3AFDeZTuL61dd8B8
puSFOcmjPTOu7PMa/ANQkhWFTdg6EUjpQPLFBge98hebI9P6BPDEG1LYYXSptORH
k7g7m0APBnrtVlKw/5bjgDpNNf17lnqf6GJwLusqKwB7A6SVIvid7H3hp0aX80ez
XJjCPP1dQ6/E3mhvdIg/T4SXiE6UdLbJC+5l/i+4jS7FZ8O2vXEM810zQLw7Tain
WlHfF2p68D2av4MrZh8SRu3jzeT/KZUygMf0jdJ3bWVElFFmw4HCrZFnmDOPxCd3
iZWHP7Tb/eDHYWtZLKkR56d3gDNWoXQDb/GHe3TZBQ/+a5UbJ1RH8EHiRtjWA413
Y0wYnDR3r7eXbTFkW16DINzYnKys/corJ5O3sUPWjy6uSzAZB+VoAo3vwc32ef8E
yd1GcDOzVEzy8m1A4q9eMUNb5yIrjfvYmu4/ZnrAflEN+3dQzI+TU5YRK+9iun4I
Bjr4niT5+ykhh8ITHMk7SPtJEFaoKHs9SowdkN/nEp8hnNiYLP0tvVjIVN/kA8Ka
vqjP2muKRZyib1gKxTaJxLzFywbMKmozdeAE0TzYJxGo5CBmLBU3pVjYQIOz91u0
Vzn9nkpoM0aHr28cXgGzJ4xkSB7gzcQZxPDU2cL1YF7bGKOlDBnJFhYg1TdLUwGv
lpdUqrrsyXDOVQVKoiTKHl6iowcOL9Gi83ucKRWz3xCKNwG/UNV7PqbLmybiS3lQ
XQLSY8HrSpMOb9ciVMYmQ28cc95ISo3kZYFXsAidB9Sj/A5n8r09uF2WDUxCD/+Q
vfmWElUDlvoiit0o9ALFmgM6CEoE6a9xsS7LeXbM0RsN/Bgf3rPa6FI4Y2T/T9aP
WBWZlB0jHPQwxLhc0MH4MmeknosuXqSJuCT3l/rjJC5VwG7sjRWleM2X6fjPqxJa
tyyhycEr1eZH0drXjiwXvKzy9VBIJTO0Z1QONEaGZ2neFTOYAnIfAz04SV5DLVp7
r5mUnJgSSefWt4SX+6Epe5Talv8ILBYesxrgJZ3cFz5f4Irx/Grv3OabrFFWTu9Y
PDV2G2sdvfoEUxtouihnjOBjMDwHsvp1hmBiZjRiy6tsM7lQPO2yaTE5i6VkCcnH
1BuUm/SkCoZ/om8mxtKwYDtxTrAERshbcIGyMNFvhacZcU394SimDVe56hciZKOn
yqT1o73fZeFUZ8+gKxvpWrmMol/VrmCFiojBKCy3KTq2vLD19bxC9z56tZLLqfDu
BD0wSaOTrU5hEOQe7PnncLIYy7+jTZrs0CPMPBVhgwj+lbgp4H0Cs1219eSPGh3R
qJp2ursz0a2hVqu1Eh71mgsb0H1jW2SvqL16xw8diV0Bi/XcG5K6VqNFZ2x+nPR7
f/5OOWU11HrCQG8CnM7FR/lbZfAk1eE5tQuj0C+sASjDvf64htZu/XH27630Ivtg
4dyLM676cd4wtaED5ll0GFEwIVH1p4Gbr64vTT+ilCNIHHxw1PjmjZ9X1E7RGkia
wekybqDiHbxLqSKrVLBqGV1DoRAynyZMpbbwDmVCWmk9OeSlhQbxsud5ivJmGpaY
w+RbWPPYylySCzBTp8Fy0Qef0t2HGjUzRfGks6ADpeP+bgO5y6gXRiE/W6Qh/obJ
dcTNgxJOK+3zQ755Kl5PZm22uo1Lyw7AJ4D9q1I/wXQ8NikYvGGJzWS0GiaMtmIE
dU025RPR528nLYGNFIPkX6hyyf9Oofv7wt3Ont20SUVbkmyISaWesuJt7ahx0NJ7
IiMSUFdazs7jYdJikqUON7JrZqAqjlXAi7ZiHJ4esldUeRMm14Mi/Ut8AGfJF0PT
Cg7sf1k38oNPGjcDJ6ZPhaw77r59OkgPftaV+ZBczkx1lV10oyC3MLFSnYosUd3p
MYnvqai6U8XDeehDVyr0qj9qwaq44zsSsUuMbDb7v0oUFOoGeXLkdRV3ziIFLGLZ
q9LFE4R6sBgP7x0/7ci4DvwHbgaTW2sj8q6l6X26twDXROuVgS9VxZEKuZw86Olc
Ht/238z6DpgqFm1OOCWApyQ9LXu3k+zDCPJuZLHKv9hGdTrrDhuW4+KkE92jhNrw
iQFmFcroA7uSJSz/2w28s3jpWZu7eGiMfvgwQ0XC2yB3ai8WBXH4C2PwdX2jRGc9
G41Ge09I4cMDKlcpYTlB8G5ROntRP8tFLnaI5XZxX0Lt6Vi4eZ8auN8jlNvRl3gp
sbIroLtFc+HUnasJ2QcqZPe+p1vfVSnlCspGYjpSY5VD6ccrgD4/QgnVsmpjKlsF
x/QWQvOF4c3nEPgdsRJyVbuK2+KuYwnNQs48By1hFZ8CUN1gfIooD6G7BeP43vWE
xdvkLYNci+zi7oJtB/nBthDkCY2CSO7hSSsD9lSWGTxHDZfSOCfinkngOGrQlvaq
UOPBpbao4WBpgU3aPri9CHkhTsSxKXJzStZ0mseNHvPD1eJ2FlZKrHWt8ViNL57H
MF7XkevKQNXtQZSH75hA3LTLK/vchHfgl47exZ64ZHKzw2CoY9KyNslMz+Lel3k8
0LoSXLmHLWnsq7kMofYg1PRg1I2TMGeS3vsx4SsO3DUyrFGsZKvlk3YpiZdB4bsO
rgONI0GLDQEzoITsGOiZgIv2SHnDOhK6aECQgjAtytj2GjxnfPSXPXwwJOW9PITW
0ByAD3yMZx9YKyCb9rtQnjt53nbjNIxWk/GVhROOyrAe850fNr8PoxjRpHeyGwP/
/kqVzud5o4iRZi1L5CjSsUC4mrVmsFVgUvCnfRoqFkEJu5qheIWYkLgjaGO4N3US
sbGHUWrJlrRBZ5qYqjyxj4Vjf4BENp2BCbeP4jwLFfBXN9rAkscB3JM5ur0D2aK3
9LmDt5hUKjxdA64GjbvfvyeOSeDbGQeSISJ8woodfazUpRgpj40efiJD6ay23ioh
GZiVYNaBNpqm+WghWFOPt4PCvs2D8DJtqK+HfALoUqZUI06wWFXjPVYjVKt4tbRM
no78VQGx+OvbbfQZp5rVjmfpC0MIjBLMBfbYLahoz9GSZ9fYhIACvgIqvMSBx1h6
LogOAgiWgm664fowL3hq/Iobyt+Sn2plHx+dONyabZ8ctjgoqkDjo/smmFaH62qT
KXp6AT2t7VQHXV0S38Qr2BJxskEMts17Xzu4dzA6B4oaA1KRL/pdBtTeZrbj8w0H
DPhvhkxmbB3/oCCXqz6EHcks9IcYOvaYQjjsuzuEW//tSNpDajZPRTaoWYwPG5Li
nUUMe4JekgMgbWBYSq6hw4zWO0onMPl2vKCYBUbGfjFOikuqhFpZ7VJ+5dhT2z1a
Gl77cb+0+8MfLnaZYKSWXCPn1KnBXlzOKWzm9k23FxFlmNUJvckVX63REUSj8bra
d+UCQchptyiIEJsGOdbyRGJX1Tpc/PSzXc0XJogwFwBsb3aFN5f5eiB4o6N7yLcH
xJpdywES868CZ68XmExBxp264DdD0exK/okP32Bk78asO9ybaKWTLpchvFTRpEms
7LTzAinJdoHil0cd0CKCfgBRjfSSC3KgWUfbh2+PMdfyhpnAUIXQ4iKtJzb+622s
Mr/iAVNOFVeFmrPhZktLTMNOFWEvIuRlfjLJXTeX1h5Vr3QTjot0HW2fEqtZCnMK
EztsCMtC6JU/lLbaOacod27Q9RPN4lq8+7Hy5OwkEXuTY3G1W5L6ny1XUq9c0fPg
+n0gG6KpdwdMFQ5pf8Pr79JyRNJTHGRVZ1ipcYSsDxhABnju3GuBxNHvKsXTUXi2
JuSatXGZlH4OvpODYVGUGvLDlXbv10U40HXgYJgVEa9BlFfEsVN73M4KICKD69NZ
ix6+VcJRQKq7GtNcUlDJOyNEfyzzm3N3On/Q8nvxxTzJyTKl5iKhVbMEr2MhluNY
gzM/rWf85FoBEluFUmC6VRLtSmWbJYbiD485Lk4zvdOmyLCTyliTY42WL080+Q5N
xzPimy76kK88arOfu56uGx17/7xinsDgRnV/ouCc7Ys3QNA/8eVSST035qTI3Pvm
oJQ8q61uy+3l3l8cvUeAm3Q0aScMYFuGfGFMaHte7kdE1w2n2O17vQWYMLBrbgxf
zZJSDl+o97Nd54MzRVn2CxNqJRkl8HRBpyhSErjdPQxPVWkNso+zBF/zBUKMJFH8
VgfX3eCoxbHSQAcbF4tfztE3neM9J6dsEhYBPkrh0QdSVJjN/mKx3WUgHfP2xYpy
cYLEu0T8wyNbYUWEE32ogHiyhNCjEC49MQkFxpKZtH+S77zdayCzJS6Gmw/rjhQ5
2bIewf6Xts22C2N+o3dZQA9EiJ0vUCBui4Xy6JZOt5A0T266AoTxcaB2ikxutKUU
JetPciE3cgUA6jD5IJkl1QYbpDiX5pxA5SnBo8yvUFLV86HOubPcKeIkr/tB7J9b
Jnqszhy09LlUQ68Mu1Ae6rcyE//0ahKULjr1Q3AS7scV3bPHmrymlB49iiBWYBfU
kagNKLHO/4lx89LNU9BZGXCDFgXqAxHFi4JnmCAInYX/l3w+qvDFxbToCsP+fQu6
G6Gh+vU32kOPOrlbjtuwd8sddclUNh/H8tjNuTQuDQz5EqdrYoXRFYUqfC/xp1Hh
Nu/PVte3Ehc5OBqIDdHuuB4FGOVWvIcPErtQlkjxMBmVtONcKYVjJCf/u7I4aaym
4oxLwMw3rilTJqQsMhvCaG7F5hlbkbY79HaQVcR5e0lcR7o7i2EOpA4+jU+ZM5WT
bZRBAU0i4g0CEl8yq/equYyManv6LWlp41mlZKgzP8hrQatlzYTxpFZwNCvpuJlc
IBMsBkou5ZaJ0CHueJE8KdycVn/Fy5gjuc/FWWV5GwFmozE1VkYqOZ99kiE+kdwZ
6KlKvSPfeVPxAEdfEip1L98CJq9gUMTUFIlf5bJ66/xg7nCP/sD8lArcO/v9R8Uk
729tZ9k9B7o6QuDO5A4Kdf6F3lDb7O2snVxea2RavNzgyJvymnfF2cspX2aTw79t
xHl5RLIYdoPuGGcY+1YJxxEaoN7byKhmDyXmJYG0CML+2Gc2zAkScGos8x3YHQme
tgald0MKisMpkaomY+nIOqC1M3jLeHPmAR7bgVEA6Z6Gt7y2qg4RSLUVXqGB1A+y
ZXzg3xxaA5fOEbk6RtZgfeTLj2SGbu7xWtFUdq8by/u/vvmasXaWF8xWUhgesr7n
u2OIiUTUo/Cds/GlkeyyppiLsrMJDjn1UYOCx5w+nchkDxLhwN/V8JMWYR2Y6/Zw
Q+modtGAbC5qqm2xf1Hs2RRl48BFx6JAwax2qL2L7RkKccXrT+pOusSROIbyS2p0
L0nD3dajacg+qRqt5/H+YqrXZZR9c+z+xTSCLBuTBFP0bfxKBGdffJoMH5iVM1kD
b0IKZ1cmJQ4fnSBgSpINwydzXGpbmchMJTJ623Yw3nQNmz0Ee//Zf3euwdRXr0OV
rjCnGcB+1gdX8KhQ/CD2zr7N/FqMn0YxznjkG1MW4qe+qCyOSn74vJpAIBNRebKM
jAfIkQgiEJQijGsLvH1ERO8ntPK/TfHSbTdn9vJFO8jMzhTfKYZin01fMEVMpCiH
7PvT37ytuRBsKPvoybq0dVoCL1Ba1Qn5ytrExQ4eXLWgQ9S9ZawCx7SoIPuzOS1Q
AD+NwgacetyPJ3VrKuxdfaLQq3BnJFCnNVDmLUc1wrY3fSPEZxx6Qf16Rdi+x2Sd
eWAOOY3DSpYV+OFZNDR2Wn+TPokmH1SUP/0Idt0smW6iZzN6LQj88ZyKzHysfaaO
mOef/tcFRgtGFqQwU9heuRg/QCKcfyUqo4bV+XjjuUyN3QfsK7OyHwjR9g3sr4D+
lCduf7Zvlj1ceIUgVTERxRXaefjLpHftH1l41G++ZYbmrV9k2mH1kCSQBA6oZe2l
BO5mR3laU+zjFN5yiXzRjdA87C4SmQ9FK2VdCXkX+LT+uBum8D50gcwiigr7Qsk/
MHSaDlmCCnYLulF5RIOpLvl8LRzEaD25mRvynPsUIcJgOx5ETjnC715ATujAMuDU
YpVVSQi1J+I66tjwj5GOB5nNQGpM4y6Sq/TkD52uLZilCOyayi7FtJ39NdfNbfpk
z0TR4TUcXo+eoAeYqYVnhUejm9ouOYqhkOnQnYBNv0Ovy52Cn8+VQGeFMJH8g2P6
G9y8qMeXg0m3UEML7BSdRg95OOoEcrTlsgF7vUq/hhw=
`protect END_PROTECTED
