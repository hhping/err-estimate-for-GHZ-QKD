`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LaBNwyfe1BA28JJWPa8AG+NWDkc4nsDoUGn065NC2mST7Y2QTgKhA0+8uvlfoZ/G
8eyMIwI9ZUVZ6j/kyjoFG7cjWVvcQpYzJ/6p1kjGhHElRnjTRLUe4+Up2ssJT2ie
8zEOl5tCzQgXCzU+0NJt/GKH2+ju7zId7jXfNHDM8L0kl69CT7tKpMpmwm4rOmlx
6+UTlvOa1+aB6BlzFbsTEMrYMZVzhoz2y7nPH+lXtFFgtBRr0Zbb5OPYZxPAsW+p
37aKk/5teDfz+nOPNweReq4R5i4Lbl0XriQvaejTon8wpAzdO5M3rFZOoL+iVqht
EgG2AgU3yyylEnkf34KNPZqAzc4h2+q+q6gZcpOQKSBtDJe3l9fY8FCPThaS+cPQ
TnVDecXAJdsWk/HJD7bgO+sBtpJLOhlM2QGJE+qjJD0RJY9lWZH2Pm2iNprr08zu
r/GNwiSMlG2I7D+mGe+nkzNkK6A5Tnt3e8WtthoAdjRc6/L70NoGV6Z/XyCbyxMB
eN4NkM/R3yXNA+YXS6qjdSPLIvBvxhUTU8D4O26idzSoDRFVMOwnMStpQbj+fu0K
05XFK466CSrVyUkT5wXnoxO9X5MDjbiGAroy+cua/S0ISQJITCYOnONu6/YFPVR3
z3LIWghbANp+ffaFYimgbm8+TI3ZkwgEORmgqw4py3Ha9z2vpw0CKFO81YPek3gu
xxBuUHAnQMSFZ2vgtS4NkEOG4HZSRH4/HIQVFEtQN2Upazm6iZYDIueVKXQv4izc
`protect END_PROTECTED
