`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOT6Q+bTKEurSMTPG30mtPq20WrNDjSwEMzLLYooJPzm5Tce2wCbnDFRECktTwkg
pVx2IWgJT64wIm5cGyzkgKOf+/w8/X0rP38CCk9JWYtpMDmDKGicrnW0nyVOpjNk
p3EgbpwtQb6EQa7y/NubTUz5L6pRrrPF54+IX17DrW5NbkKaM6n7+8NbafL/h8Pg
SqOMNZz9FKhN0YUuDjJFs/xnmvyFR5kmf29NNX9JsWSRZlPmyouhNoKzxFiWsDje
Mh4P5jM3BaRkCN0svjMAib93G7xpxgdH+ajkhtRCmPNix5iigGllKVBTpmOl35WT
sZ0nDLhyPSj43woJtltbXDXZzz+j/Lqo3vGncEHgn4camjxhEdRqbOwEtVSwaiot
gcfFDY0sfUj5+YVgZWPnmisLW5ZfCLxW8h9Gg0s5gV8PaB1kOkkRhICApPD0wcRA
M0f4Nt1ItjSouaqL+GbBWceUfoi0Qa8MU7kFpfLhtTgzZ4XPDpNPqMHqwEcWE/1n
PUfkQUV3FfxGP6NdPJImJH+gYIjAa7MHqfI2MxWTHfsAfcvc4mxO5TkPK631M/wN
M5kaUODN14PhJhcojDBTh5WrecCUKHTc/SKgY4UrKBYfk9x1u0n3gUtMEc15PmC8
btTBNcnUZRHB97Xa3YSak/q4ogt1fx5CSbrTM+yIdDa7vEd+WbKiuwxYit0ZnT12
nythk0hyf1q6WMVNyqKcatoVdnBFduD4kHY3SlhmcFcC2ABOy2DO2nbbjCc6nsdK
N22waYvrrHsBwaupG9b2nQEtn+D61xuyeaym9ffYMkk=
`protect END_PROTECTED
