`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KUYyH2QpIAk8PSbyr81EQVUydoT/H7sY6gpYBhIoAKWPcCLmid9sCw+fJHvxxLMS
WXGjqS7DFTB/i8HiACujnEpcx5k3RVGZzdJUEizDXKQRwLRKQFq0oudq9u4kSmrd
GTG1XZo1rFHa4/sYN3PONtZk302dPMOgEl3ZmGpN3Qnd9u9BuXfIoAHObzIOp86+
L7MOQ9a6uGPdnDeF4VxnjSQIL7dyf/t/FI6w/fBLyAjG9hh0ceesaJSKaVMj8hQn
cLj9i4HGUixX1j9if505YO30klCfqO/D38JmeqAZe8AQjWGlV7KuQjx9VariPIjn
OOReOcOi0O1FfPCSHtjcENHD+6k5rLDSajf3M4MzvxtqxRhaIoPZBnkRv5MdCcny
fXsQbXt8/RAaqYteuIwJTZ+NIEm5IjwSJ/rGkrcO1hcmOR1oJAHhiOnIci1EMWb1
bvXozc39Z1Vry7nqyThN4T09/gzwVPcACtWX5nIMtYMLmvIecqoq65kUZ5NyYAM6
VLWcgXa+u5hYJSz5R+kzf06tkXSwzYqDbgWFZMo5vGlOfTBYnQgVT5UWFQVS1LaE
jCq87AzDo0QuWE7m6kN/pFnylSiHlVD6ZtwPQMNs4+zOnIl4njpo9p4fY6T3KCGK
9e7kTVpuIl4GQhtQkH4f5Fu1Q1I2SrI8cjnaBvOB/EwTmYzoNT5gzJ/PxWaFv6qi
C4CUvzIrkg900Gu3X/f1yeI9Gx2222WW20daw7hJc44HKU2PlJN59oTYpu8MBLOC
tOvvL+0FvvRe5lRRhhtCN/pP6WgOGpD3/zlGJ2ThD3apriuxROb31ctojLt2foJk
qFKIDIAHdEjKBAHpsgO3X30flOaOrT/Ku+ujnbSSJdEHMAJ5s/q86o7nM0fcoVRN
bBv7xBoo/pCAj0DjDpqyz5JJK6jFw+MgtFrEpWaUm3H+XpfJTYunc+3Nlvrj9YH8
g/+2vpMPZtuyUwKotHbCo74HPBc6HeVL/jBvm+SubDPWcfcxGOC+GrGXDkTjNLp3
sTCs3TewN8cTPqVstfAgCWtbFArasuaW+K0p5NfePfN+PvlxkfqF4VsajLG7EaQm
1tmraGKOZD+1fi52ELARbOKAOYP7aLfxd3t5scME1Snk6e4saKKBoRLGZHNwaSHc
gGrq8MVGfov8RVYi0VHEYzNkR6YFueBXhSGijDuKPxn0fEDJEMkFR06oXB6uqRjL
dz6B0b5szpBRd87ExFwbWG0OG2Iv173ql7qtD6JVncFE48Twp1NRb9q2bq8/lZHO
qIKb6UcLw7PNNObTCmCny6sn96lHx9goqYqtYla2w1DtOCssGhb7tgvMs4jKyvDd
9n95Wv0KS9lKpCyCzmpo8srV/jKpGjVI5ASTuZvnFCTQy/1FbQU/D+3fQesblRHK
1ruFjMH4Lb6l9lLSC3RQS+0NgrabmEU7XLpgrVbbg4h0hhXy+EYLZJGUMajd+6Uc
sWm7XFVXDM8waXrH3N9Yv8yAZJcqG7VSUeIANNa8WfafVInTwkhqkPRb5rs22x/T
eWJbQ6CZyQCFIIRk6s4KqwiUgpeOgFcNictPE1TJX/wIymf2Kij5TFJoIGej5v4t
hPGyGYlPxOO4P+agqyoJq38bewf26zeKJ8TA2T92xDNNnJNDxerk6cYcC05Y00Cy
gSfbz2nFu+uYJUzmJkeJL0ARvQdYWohCziLjoAptXhboRiirDRXwLPPDoxq5GKvq
DYyG8V24coBDDY3C09HQbXFlbWnl6mpS/5KY896CTvZ1EUrbJ06ZFuK9OIVhzZiS
KEOjfE17k6GVp2chYPPLG8MTjgSh2ZGvxXJjiQS7pwrTnjTxdVBWr/CmhS9UV1Li
ZYTYbJoHXEPgvacbXK6flAOsCJ6Vc72cnZHCAOlJDS3uYvb+Z84h5/XgNIcbksb9
Pi9Dl3FmYQ6v4ZCNIXy6hYgtpZN3+5aMUG2yxw2tVjXpYkMj3sV5+VkK0WKCUnCs
w+gNet7SlUC2F3sBVpsKdRLw/bM1dLz+vRX6OM7J07inh4BxD40p3DZ+wNfuF2Au
JIUzIR2RSdiUBB9bfdUkGEK5pX92keFwFcB4FUafJFAcc5LcdvGF8wSuzzhALjah
aaFAXdMPbBZDniNXoOa5xXbCXCyDSkRCE1DOcZMkuM0C0xrZ8x2mz4ABOYrVD4PD
qoBvm/V7Nf49J1C5bcay5/C9CoQSlPXASyLGfUi8Fp2PoKLf0KL7+Wfr8fZZ7dF+
7i7UIfI8zqJjtcSmvq0xw8hfPv61RM1+AI9wt1D3gKnpga+FryLiTXBVvGwDWIjw
fMp+blNsR5d8uKBsOemDkhucQ82KgrN3ZswWMlVbM621wIHYscEMIlmzn+NkI3uu
13TGmxfWv2i62k3RqmRnm4ZZTpWY2uHPgZy9zoKA7hNmqFsU9FEeSRrmuA4pWxRe
dnhuNNC2yQxHxUHyObehpHcHegaU6lvPs5xgLJGdDm29vfoAY/3LnAzx8huo7yW3
so9N62iGqL+nL8oArKsM1QHiTlOwl6IkF4qTKcheYNEe1q7g8uo+qSFVf7RJSrB+
spfm+9NDFLtNjVguNPeB1vaVixOnRt0/LQFhhHRh13BzqlSAlmpG/rK8cT3C8ByH
v16UXqPH4HAs7VVoTJXGpFVJ39NDYdxRy8VelO7bJ97sAW4r0Kx1w2OX3kpWS+Pw
Wdm782RPNCbPSrarTm56yQLaGHdy6w25FO3pR94vL6N60hxgclQSc9UmhdyO8tEA
/JAHPGT0ETwfs3N9zrU6Ah/nJYHfiXwgP604E4SxwiHQS38etgI9Xk/0GSpiz8+g
qStGHBKX4GAMDOKzEqbMMZUikoBHmECCVfj7aBItKlDDDyJbXe4x11Ygub1wlmU3
yTEGZiOk5gYaOQT9C+cbXmRSy+YMdUMmoF0KuQgmnrkfJEY+yibgRyQ4kbJXiUJe
HxLima6UrW1BWmysvYqaKhLm+emkQBk3eoUiRsGI0o56vk7TNr1n2L2qdLFGsEFl
Iv3NceevU4mWUnhH2XgBblwUNr2lo3tuS6y7RCQJvb+LJbT3YjLGZasWOgzPzsyd
BGKNyqKOgfeifAnSvHQnwBvyYbZlSfBRKQJfwBbN1jIlRXEjLEM0IKykN/8klm/a
Pfn9mTkQVIIsU3sqvSx1MednEZB6xSVpXiBKzkigswFNkjJey0kYwVRry8SS7jmU
`protect END_PROTECTED
