`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcSHgrpxKBFwKKDIUnIRf6Fn9+SayeCuPQ+VseUZo94cmGRjqSgdLf02zEytOiaH
C/2qOC7NBY5glkil7zon+BT4j3krTdbOiqJFy6JvSr5Hisj0xxMvKXhggoLyOKHN
iz2AZ148d1/NUFfx6C+LcVEwmZBohxrrjdw9jEIPdLnY7Z7tv9wOztEPnUPNfNte
xs5pwKVqscBUJQdRSmuEkpv9tv+iNPCxkEcVWTlO662unYEPaJ9h5FldLyc3oFZu
Ge9OkQSIz/UvJ2gwIOQF7qAQmNEr0jA/bgzor9G79LKrQsAgeOJkwZIWDLHWwT8e
ntq8KJk9S8YwYugpfkTwyRLCQVzrDb2NHWO58DFd2NEq7nhYKWRrlCjgJQrC//9o
V2ULtwRssfzhabCxzQKD6aUnYkShthAiOEqPftgYSvEhmQDFZbeVzo/HQt2OjvtF
QIBOjixP3sUxIZPdKKSRBNhBz7NdA2AEbi0vsC3j01CAnvrZbgZjwT1flrLXPu8N
FyKa9a0cM1FAtrgHmEDBwndj4t24vXvQcQVP0Gh5Y2FNxKaTcrXRse6bm0Gx7Q7/
FoXHxKDdlBAOsqNDhn5jmG9j5bJ0BSwFKwvlS/tiXdHyj2Hy54BB8USTNKGjnCBk
v0LBZ1ovfQiQlStlDv0cmf+p4oZ+h4YbB9tsqXR5ONsmeGtrJFAIIWJTPuGMh3DF
9zFZ38SSSmeMlWm4fxqIDXmsGOy/bXeIfJH/ykAFsM3NCoCtJw8tJkbh/bxCzdz4
ay+Xx4O5EajrlSFzZFsAY2nV6XXpyl44/hZO+ZrWOV+semYfpOt1p5riKrQhskxN
sFkW3mau3nidmwSb9oMDyhf0jpysxPAAKFDbROZn7ePrzNTS1rPxdv+pCkDYdAIt
yH4BLzpamzZjutquB0Qy8G6t2zKUutY2sEYg+vMRs2BRvud9pQ2UrYbkLfGjvU+4
nBDptvWROBwLMuX+89CAN3ss5Kv9BcmA98Wq4LVkftIdx36jBvXMiSyYGTS8zi9E
6lMiShpch9RN6b0VKu/tkWwgyOsBO5q4jFZzftUn8mAeThzn/UE6z6dZXSoKeFlg
jAHQNEhm43L70foGzJ/eGDD9gu00qN+/p/pkDtVTLJhloiQb7rI75WEqM/AGm+fk
TaIrYqE7fKpxvO2gx0uOgNzFQ9yIeoLRP2tGojg2eKd8J6LRozmlTVWbhpVlsqR/
NPoMkFcrUEuxmEdrmMp00K0EDAVtNvCeonQrWAWK3xpApDfXC7y6MNLu+/R1WUKF
bXkMC0LV/BgAYVdsqUCowXO/trH3phpos4kgz4W8i3Pr+nL2g8UvxM/LY7WAV/D7
ZsS+8ojNjV94gpdUT8bN24/qjg90lLgynHGxpEPBGcLajtD0CVVPTc4mmMVDRL+Q
dJ4lrfYLL5xcrUj2hK/CHb2DMtVPZ0Xz++y+IvFCl6Tw/Pk5Q1hH/z/cpqnlCyRt
tK+Gs9fezkpZrM8qnARuFypBPV0+V17mr9k+8x1zwPA=
`protect END_PROTECTED
