`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBt1JUQYCu/Ujj4B1rtvboL4EjWbaO8D2iMO8CVNFyC8vOH4eSZujSF8WPaSGnsv
LMfaUZlgmDAWmZXQgdUgmxLINIF/z7ERnS9FzM6VjOf/M8EkWQFTsA1XhEzB2mYT
xAerLlurnHpjWvRfTlOP7gi8EZgPXaHHOL93Rnen2j8QYO1preX6cLzCz3zMykoo
H5SeHr4FU9Mw5CKWgE+SyucT/3eORqxQEwfofDHQNLh++HkTT9hx9hwtM4J4MNOy
ve7MFlQ7KzXYfRIJFuc8y0/5Dm/vE985YFi7ceEl8j9skmHCX0VJOe8mL/gnx+Sx
x4ZITjorIi2Z3LEaJSlPwsVkGPpnn8nXU0m3rKgLHJGMqJT07UxUYT8d1sb5ANsy
ptPTmzGu+0Bdq1LXEqzX6fDFmQt5IVHIfHnaeqQQl6UFqnexNSPjcgICRTCcJKwv
QJkJLmitbLEZbyT4ZoTs2RfeWI9vQg5SpTnyUJjz5y5f9JiF8icZg7d0xrHPmfWR
IMbWH+XFPDT3OO72dphqsKbT7ITkG0KKHMJCfslzRJ5n/JglZbO73aDk5S1izZr3
sPJDgPHOYZE6JX2xqi8VeDC7t4MNACpdF6cKN9dlNSV853oeCK2jaVY6rNbtCDzb
9+tZF9ULmaePxCcS4KkLoa9g9cEOyzD20/PE9k4lVtZaV5n8D8Blei19lDXZcWGY
dFychLexK/ogi9AjZ9kxrex94+VW18+hvLol+Nx6JUM=
`protect END_PROTECTED
