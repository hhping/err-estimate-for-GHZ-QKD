`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hW+8cZXhUqfpYgLj3JtEeuMtzo8LoiQDu/JlmECy8oNpQJK70y806HvPwrLe2Pc8
jGbVpyiyhJl9uPSoy7LpyorwtAHjJy+qsQ7ZlQgJBuAcMyIBpUCsFFSc1PxUHvBB
v7HFdNF1IxzRU2VoOY/0+JaoK97R70SgJ3ztrH29fWGDmM83/A9Qu5TgtwMAUaGs
fhY/pAowpbKGfmQnkhb3NpnhOEZeW/i48TygPF1ZM140QeiHGmISam0T9ik4i0O6
J+nyGHpq+OOZaLTghnhT7PRLjrOPt6uq3R6gVah/k3AIJNso3Oyplop/WYvXDZCu
me3CN8l4hVm1n3hTkYbP+ShrkrPdTKAs5wSPXo49ppuGZsZ4YJ6txqZLNfKovMN8
6MJsxi3koebnQHkfTxgKclG+tBnvY59ieC4F+dc0qUjfzvvqFKYL/cp2yK6GZ2qA
+tjhy705QtxMuUk3uZgzgdgG1HQRHt55n9BpZR4kQ9ZMxtJtBg6bYa755bSR07Yl
4I+q5r+YzAgMpGe6iDrMOBEXGGcs9YXTqhGWTKvosAW7NMUTzs0wAnkackauYoTS
xsAoes+XWxNmMFarCr0CRDqb8gaiHTxmtpg51rgFuWx3f+ONhkmA9pgdmZtG7ebT
rQLPiHc1i1OTzDczzrDNY8R78t40oIIPdJKY/69MkCrsMtWMYm6smCrJjJHgWSNm
uxnf9moLjylyr0E76kGRQfMJ6UqD1oldDq+1TQnmKoK501VwGzsmS9SMaWzXOR4o
1ZfwNdUKRzjt/YSIH+S+ChhSPutpBAdiEb68AXBw7GVyhkuEYLSzkKdZ5W4jOzG2
2LVjTCJJG9CRUSk2yjSa/zdCJolf9HjN06dAzBtEMQvMjhja/qi1uc3HihmWcmxW
ZzGdfuFV0dTFI/eq2pXH2p3COZoqtRzz6xzQZ38lpImzkp+dyg/nE2EqLWzYl45Z
eiPbYVJO8DA98THcuEYobiJXEG25sSVBYFVAgzmBtiKyUFhNluqMsjJURxKMridG
ORUl+YdVvRocOZ/NhuiH0Z2vSUJ+4mgMc1Lb6r1S5gT7IkwTUFS/CYglSZI1iqur
Kga80COulSQVRpiDVmrtv9cbdBK7e542lo9eMlup0HKsFn8il3Y4qc5YRb+0YY8Q
vffECXXIWz0Liuwr90U15OpESMn8rFDelTwYYsz8fYz4uEIYGrXG1ID/tTrk8RkU
jo++1rJXUk3w1sMXFjb3oPvLeXxr4DaXnxK69cuLBni+2mIXOW3GNYKfkhUVOQfn
LOTlE0+hXsBwsp8CU0UA/KFqKZurjaLxaZQXBIFLpz7bFAc7j//KuYgt1q3m5WvL
8+43RjbLBaLSV3A6Dw7ux55y4P4b2p62YS+9EVesgQLl0Tt9nqbVtf/WaViUis6o
/rgzbiBZb2+wkRfK+Tu5od+QevnX/obJFUAgk3496nYqVyKw38ZbuhTmwr1URBsa
jJ9aRUiFwIqG5QbysRGiOX9r0JqKDTOm+FjQFWCgVyWrhefWFMlzYoeYeu5Md9uT
Rzv1HqR02j15L+A9ALkSekjhYBpFIODKq3x9euMZ4G7zYJQ0EYg1PyuU7EfXQJAs
oP/IqyM7nzecOvybczE5Z9voFQ/KkgdIapO0x0NHANxPI5seJZO7aWxK6NNP0GVA
N24ij00puXZAIyPUX7KNvdXApJMl26YLp252IZ6kDqJLr1YBY2SQxPpOOFI7V/M3
Dy+dmZhuO5O8fTcFXADhjo+xevS6EkByMHmJD6T7N8Fg7YB3w/ZJkgWF/c+VOjCd
7qDK1zlqj8Ey5LRTxq1N/bJAST/+uMRWZaB6wOGPkLE0r7LP4ltMLYM75dZ/613q
h8RkprntJb0uRcPR6YdmWZUDV1e4u2wv5Bmfjp8kJrM/qHD/9jgtfhK6RL+2+MuL
zAaxlhtTCYJZXXxMyJz1DlzZbSP3wCN1mMK8onMmCPrsR/3vLLs0WCGWILzpSIii
I7spMNyCvuZiC5ucQovaOE/74aFJJ11oTafyedTyrL5fUYkdxBRblnMqGDsqNMQS
EMMmT90JyBDPsq8WX0Aogh29etQaLwLgeOigZGDKKr6XXc7XaPsECkKJVmobEvG0
JlQ6kJ45Z0SG3lwCDnVMZ6Ri3lFUQLaoXO4v17Z7o995RbT+zyPrmA42KDhT0IS4
bNkApe12RLpCZ7byqJ30416B+3lZgriDE/pIrE3KBvpjUAilzyQD0ulUQlDH71RB
si9m1IsgZ2X6qmzz5qqH6M919XvcAsDt/bxDxvksaQG6ddIK2dVcswYARWwwklrc
l+KDc4zPFk4ACGkk9w95GO/8sYFfover6ayFvhUp4mSGPMpFFyeq0mWRNLD555tS
R1MJBCEwz273SndJKhyfnqOAT3g5V/TEIlXd3z4fUzDCnEvouhxWhGtwSJVfjC9N
F4u3Sr6vGrDRXmmjilgtHG5sd6+YJXRylzCIOA/5Q+riOGHpfanc/hhPoaiQ4DGI
pHFsSGnrracZfBLGX5fx3j98vhkuWTkfCoKlqNa8Wtb2AOJZkt2c0HoUaTKzVWO4
ktATkrcGmyxCjiF+pw39kqhs56N0k5tOuLfuQLJYqLTIWWbTiaD5Hsv0SIZPdzac
1p6BvIb2peKh4SNGFnceIpGbrm10XpzerflJUGOAbjpmbfXD4oHVmqJBcxQ5mpZ0
E0s2/ThjUYHYiQlUvz1oTX5YzotdqTAGHREfiVlpULK6/hUsoCBthsgkNWlycdAT
8TJWBAgQHLzbQ0ee7hvgRIouFcZ30oSGLxu+vIFxEvfGSqtie6Id7xa81symKpul
+ef5PaQw7SRcEUhqRsCn0G2x5l972HXA/jkSENrwiKVd3QHYO7yMTTWOnPGOYaq1
wDc32mKv2gVQMe/2Lv48AhrCkVKLfc8sFChD829gy1Va1zGpTA8DI1A453zRzSBp
9lxAJYKOXZxk0ee9nFcIPOJ9ud5eEAKIAcNlP910mM1zOfd5r/9QKqcENNrjuHQq
YPt9g7ztTCFysN6yk0pUnQZTxZBC0WgY8IR69PLQSbQyI5129LLmKPvxdZFjG0gv
qHwf8EuV9yeGH1rD6qNCnWpRz0fwHMqw4xANJ75izZIW1waj/gmWyVrtGIFgJkxp
6S2mNIm/XKbJQGFMFDLZXARc482Z7cKFj5p8goIq0c6SarYb9S+RRtuuk7KzmOx4
cW4d/IKpE1/85ozUJaE8tZfXtwJLnSTjYIwZFvpYaUK4UPPk0GGv3mCAcBP3uMJU
hTk6rD4gBPdfLLLZh7NqjLQidoI+/YEn34z3IkTc5lLEnnLXA3Q2QR2+RGJ+jxao
GBBwNio/Q9gyfJeV5nesMCHXlt3psBBEfhjN9PVqIf+m6LaBtFqq6urnAIn7gVIZ
DIRC3w3spYCShHgnAyqADQggsietpd2/2TlhwxeDafw10e81OJ6/KcZ0FBbW5O6R
qm8IiZjU8nOGFfp44aFELESZtg4rZLw+T3Urn0JC6F727kLq/iAL8qoHEdOmx071
iIU0DwvUNUhABxpGYBnL27eLFZ3xQI/sbsyAz3C5zmjzbwg4P2RDrjECoKQhAlWG
cD9IEPCplobIBDWIvAYGHvSdqH2AAKcr6YKkrq3EciZ+bZRZ5Sbg5BXhL3wa7S0C
inr+qlFD6wzy7JCeCK3dTxdm5kmyzbsDpNBOICRMsg9DAk6SuKQyOQY4ac28Xmh2
bqPxSbpFRQKWeqxfUsxVF8z4cYg9o/QZg+GPHnqklvGEsAPGNUAYXXEXngDLs+Oe
EEpJbWqoTNtKe4KBujsNTx8V9AF7k3KDYBcXPnX/s0sjXAfZ7c0RoMQ16OZFnifx
grMdVMG/ZNeYk6Jgp6mdHSY7jCpXUIbAYcRmTnbhdx7Z4SULQvnh8sv/erxdPLdp
0A/eRdgAh7OyWcJ5hAKv50YllectVmiTklQvsBGbAFkfzlOcS6xwgTTHhCRni6Ms
Vcfiyx2ItbiFH9eikYb2K0yL/fPU4fVhTDLCVd5IDC0AsbSB2ufnDmeqR88DucLb
NrtVdb4fR5qIv7pPWN2gduGjegM4gZNIp4NtdP7cWAEZc7BMZepJPF7PnNc9J+SM
J8FDiviCekC0qcggQFsRGV6z2gTc32bWf8gc5UlUVX7G1c/2f0wcBgksrKlLF7B7
QfEy12tz824LUgN1dpiqCdzic6KDjMg6JG8Zrxqa3d0J6UEbxPZClZIFTu8Jxs8i
hjisqvOz6cu1Xs+R5H8muKS89ThUVDgD3Cx3K5WH3aZ2e/tr0Xw07jOPx64rgXb3
A5v4780ZMYfB6JPuqx/CFVFWs2HBRZmBUgNEqZnBCjGj6+I9T9yyvHSu8MwgP/AW
FIxgsFhjv+U/Y0C1aDDbtf81e2xGAGLIsYIvpwfbTnEUkh4Q+23rHH/I4wm1Ejeq
RqIvmF+ABna4LlZn3uAM/q0gHRiByLyIZe9wTZBTKHpEWTuL09LOWunE9PUr63vP
T0SBextFnLqXODBgSienFprspfuF474J/5zp5zyBAux9nB7yvUCVErA00sBYquK9
iqlZtkM+f7uZn9cGI1/cClkYkZ3e5iwlYpb3tvWBchI8P4P6RWKvQnt7EgHjE9hg
6MVCAyv47U8JVlpgAiACxLTuRXYni7usWSgnObVATeS885lLGYPMVsrTydoNa6P+
yoJqGGHkgzUn1lhrRe59YJfLrAuieElgLlpPFggqvUJNjLRAUzrsSh/iq2LXt4U/
qzu/OMqRb0oCYgzsdFoUfL1jc3mJXQ3aIkWJjIBH0feT1DjghyPF7Zl5zgVSZXkK
6MtqClY5zeeeCV3dniwRRPed1RGqsnhX3yt8czLEwCe7O/LrKI6qj/moNrJyuDe0
4tZJfGAZj5Zxz0st3+HSoIN1TBJGousLzIASLCS48VbyXBAfcbKrt+D2dlvmo7T4
x1i1xKwMdJp5IpekYamVOqSOkiCKhRkOxGMSq87B7n5lJxSX7HYi9OSZhAQdButT
5pj+dn/63EWYlNWEPcQ96eib691pcjwsvqbAQf4yPh/GZEJlPOtVoLIj9KSh+pPv
pKWQLrjQhJaX5HT7gQCsNMkSo8COWL8m+ZbRSWFNGplG41wStgLSX8taMX1f1CpZ
jSq+bzdp4KKiYsuOxuVX3DNTyciglXbM05j8uQfj73wijOIkq8KTVS4QXjKIcqO9
o8T3qV56xEyuvAJhwMwFBiGzoANIJ/5g6RElI5kPbNuuN2Zc2MCOG7a10CBv6s1f
H9am3yFrSWa43KlqwAu3nEPzigl9ClZslxARLsWSKyGvaNt56HVJL8SoQlqGGxk7
Y/FAO4kyrHdGPqIbfhNQUH1EurOn5cbHP8Qska1kVQwc5NF1bORR7QmBqHnD9a8W
x5eDy/OjkcEg6mya8WHS6yKDrkUNtatcV0qCCUrqn9/XKCERb7j0C4a9kX1h8MKA
kaI1w194IpU0VF4fW2xjsQZ8QCw8BIvjv+2MmoAVYJ7C9HUypZZe2fwpuEtbk74w
Yiw8lOhUzmCxp8E+i1fcKEZMsT8m+Ks6QhPda4Qyfu4J8cAnJdHG6UQ2hvpsc2xV
VN6UquHKqK0SMlpn9X95+fDBGlDTPrSONdnjlB1ZmjAEcHuAW1lGkkYo5hx+yPOJ
mcKyk+ftcXWtItZb90+jOmCm8cliAHdf9jfflIrBEewZEh4l6OkVHNblnLk1NplK
+hlmZ1RCJ5vv1EeCmTSr02M4q+pMCF7fYoNAeH8bzOQQ4TUf2XHpQqw1W4WdY0vz
CQb83U4kagJhhMgJ8APn0CfEQAXuNRIvcoNML6oHYfNdcSzZvcAKmTs6Vo3U3mSe
+YFla6BE3bmvSdr/YNs85+t6GC0ctjye9xyYJvjWCGuxS6z03qgussjNq6szqPOR
C/9j0LPozRFIfH27Jlt6s/WhX8enHRRYx5T0nQoFjf7F1nFcEReT336YNVBMo3Gz
G1hODPxc4QmEowmeFmtguObopaUeiQsL3+FZCaBGZgr/podWvLVHPxPO9KX8fJDB
uI9geLFRrLLO0mmm6xQIYZvkElpieS9vMB/LJvLGsP6LjCbaRseCQNQMpiNkg/Cu
gsw3zMjTw+sPkwIlkr+KnxYNUox3g3MJ11v906qpVgE41+XxrsiastWWu5+g0o3w
2S1CVZWJw+QN8GWHPjXCVw+aBTrv62/PDuwu4pzr0OTPioUwnUcSsRxeOR4Ro71R
n+tX4sWH/3PGJ+mFg+IG7xM5+vJ2gpAHUJUbuUN/UektdmSGqcOVMe4sOXeGZFhq
M4rQmskhUtPRJzqqJCI0PLrkAGqOSXvf3+viYSOyjLMUdQg21NA9i7T2aRU8ETu0
ly7pPgcOup/12Lm89HY1z024269xpJdzilaGdO7JN7XXuM8+9YMmLxmlHt1wBbfi
2IKeOXEPi1ECaPkOFCCuukVZaSjmz1vv++k7pGsbE/ZaICUfHFaYlNod5c4Ufcgb
DLasoxZyrUDED9HjAUr885uFTlEdtKczBGZoxKjE5rzeJkFjJHGrbHaNOzuET6I+
Q2R9GnYfeVd6DwgsFmaoLDK/BvFtYCRiTeue+I7/Q9gFDJ3OvMuhbC9qhNvST0+k
ebI3XjwEu8lCRCdnJqSReu9sF9dyVmlZgAIWoIqWrKCkqU3ZV7p320KD37T3Bia+
r+EavVdpZFfrqv6NsbRl09LTr1Ny8Zu2HYjMJgVsdLIAQV12sV3zVR7pxFQbdzuE
GRUhwfwbhDLwznH69dScw9MlmXRln2ok7/uPpwbn2lgXS17cXZWW5GQQN9hlMW0k
lY2+xIsEbSavwd58IYlUfFa1r21QmFkeUaGl2Fsi4aX6/CRGyRHh/E2Px1BDGgBq
YBgFjkKW3ReOuyyqxpl2XNI1lm7ej7/WQek+2FMTA64N/Pv5vBlDei0shAZVAnA2
SJ1KV07GlH16q9nx2g6r0BCz1TZv9a4rU8+rPvs3xPCnoHGaJMITSeNbboIsAgII
0gs73eD3IWO3EeDzN+5EtNeGtnindISDQjsAJV7FMLqrFha7uY/ZUZ01shg5OUj6
xSarfP+1W1muPaEA1bM/OkTUSsG5dUCaLqaGaT0S+qnAs7TfVrPoIDrWUQ8KwKWn
A4Tpm0d+ni3W4WljLF7xVtg/sXEesd+t15zfFOJSWK6sUlkpqOOTqRf5IhP5QXvd
QVVM9NKLesNjuv+fjF7r84xp+kIGZDtjuhV7T3gR5+8k2cVexPEhDtiocRNjHax8
mlDKH/+ytWLXlP0jmvjrFFCrXQVnUkoMJn62urrZJ4eGZXS3iHK4HexxWMB2ugjP
0SUhXeVQRJG5qwKr4F3h5tHxPZc5NdRX78d/e9bycUIkcO5a7Jwxkv92Va5dVjCJ
mBd7RmmYg3HkSWx9f00c/8jxO+Xfn6upICbbM3da8tBUzBV/dVJkEluhYEn7xK1C
dzAdFT4GzFiOSLovkVX9vbyQX5Qu71ncIAicdfxWQmw+SX7fERS7oUCP7kUdu4pM
jPXJHb7I4x5l+29XGwyb5PX7RvHqmONfx/d71XjIC7bL13Yy9Z8udkVtDPxc5v+n
2aZitpSD0rSGbJ95J/RXcPsWydbcxkxXofPNURGiB88=
`protect END_PROTECTED
