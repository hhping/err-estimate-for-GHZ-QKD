`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PniWCWYWWJyUM+bBSIUm9hXLHZ9dz/lNAO7nHtn1H0Ct7eWZG/r4PEliamzjUa/7
AnMsT2r4mjgpUMrY07SibAfOJWwpoWTdWdb65sjOeXnOe/fohNRivLcKJtN/7FQb
F0M+qYw5DDZr5WRFESLy6EHNw1dQjVLIK7NTQatNwQXXqZQr9NDhQ1oXJ89yMM2F
49RpbX9U7QFGAr1NhBdcvnCS2GmFT/8HVxjNyZI0BqDEkAM7rSYgjSKIh10cjviB
oJaPE3lJaEs090EeN8jzMg==
`protect END_PROTECTED
