`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czvdb+2xccINrukA58oXGaOhopfeegmVnH5hCu30vD3QEoW0uwPa6Fn8tT9UyaRb
8z+lJoT4k58p6TFXvbce+eBsY24qa4drwkyPujDfxx5t3LjkjzomFxIRa1+naz8E
GUkdY9LNx2acScdjNzt4c5FWzO7T4p8V/Xus+cQlWJp5povAEc4vVg4RwLRZ/OpY
Enuk9mXWA5s8Vp7hKEXx4E7/3hUPeFW1f2stR8lYop47hTcOOCr0uQa28MZC59eG
LfXnqzeibsfidCpO+XWh7Izuia6jZwAn+kzTfALaA7Dff8U2S0Ew7x+Vt8MwC90G
M+LcnxKp3V2qItTRaGV7I1OVuISyibt85P2x3jL49+ZbubTcXVwp8Eew8YyLuBK3
RgOZBjRz+6GxQ5BMSRREd6rdTD8GDGQhbK3L246qjq+vAAtQ0nCY0jAM8vFMaxhm
oteL1BsKYQ9dzA2K5KCOyAlBxFhj2Xi8KyLLW68klRGOhbuzIySk7MBbaEayN2+j
wJQp61q8/I/oJNNq4kVJDI7cacn96QRndQXuvb/yEHtHupL0me7QUE1Voz9yzvWV
xHH1k+I9phl/ZbPUcOBsa+qNtGdnrh43qyQTizOkpm4wXU2t3svaLGHv3HU2tpJ8
pTsdGyJjYxLO26QlqHHdthcUFNpSPgQUb9qlvF427tKDacPcJrDzK7tq83YrjpFp
jxry2Kg0uvG4FCN8kUk49+5U3FtvwRPn8wFWKP+HjPtRN0CpqBXpdg6FJ+TKRFqn
lhSYNz9K9kDnz1KoVL2TRUcgIULwo65wmLIHkm8pW6GTaCRNdEqzULx8rjMDlIbF
PAf//tgH7sCowAovI2iiOYvOc95N4PouSP7bz+bIJNuR29xGwu/63hfO7aVWQskR
33v3Qyo76ZhS9avwFg+Z9zMQTWS85mTo8MlNDIdfSulcvakNlSSgQEAcPFUBywtO
NfxvaZ8oZW/aadH7BQJg2A==
`protect END_PROTECTED
