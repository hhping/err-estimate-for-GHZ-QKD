`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVClKnaOq+yiKsIJ8eoq89vherEz5hEDQ9DLWVTh/dgpPvjQgAU+yRQO9TLLTUwi
7kggmkgF22oBZVh6adbxTvOifN1TjHYLJxF2LBmvMLa11qCPjdta+cGd7BynWZG7
TkFCXWMS5jILoz1bEP+AxEUbL+DcBhbbr8QcPrqwXPqkEJlDZbEztQ1QV2IXf0l2
E7HO+/PnYecV3N+l3HHgQ2TetvbAoHY+C3v5EpVpJz1v/iVQs8oBEqP7iu7fg3n9
L8YMDrUVRv1MC1ygjEh9u2yfD6AKCxETztWmcgUiov50iiDDIKD67hWo9hvJ3gxd
tdT0A92Wkrt8Q6BT3PGWCzcTERzrL6uFg/P6+7TmUnBOfJ4sH1BeExnJcH+Ymrhs
VZ3Ny6EDlWzpPoLqtGqA0NejhyzjoNM0ukEBsaCMSJVex4VjlhQkxTPZLwsHC4Lz
8WaEfyJl3q92pXH1ZAfWid75nFwsJFyrpFmluyupNYlb3HlUTREeqLVWWmLoWNDf
F3AV0/XJPJCnYr3IJZ4W4S844qO74mT6vZDZm8qwVC6dFVfn1ELd7u+PaGQNmO6i
o7yHWkNf/SfgLuN0AU6tpyzApWXJ+nXNCJTwMUU1KOXqbV39WHdl8dLcEDZgnnRD
FuVnzdoPENQGTOTp7jwFhwM26OCyBuEsWmxvIwkA4K9pKad+4UswZcDjoT1ZruCv
lkasVSWuHoHw2eCVp9S5M8ScIXfNbRD9ohoaa7SpsEetpI3KdvtlB/CvfynvtlD9
AHFQZVUhq7ZxC0VSLn309UBr7T42wTy9hiF4u3hBulfYFJGeBeQF+3ffDY1V4dv0
GLzd6bNqVMDEDk5O6UGR8AWoughxVOOksPnjyE9kthxber9ZC1JnBoXVIpH6EuKc
sk+wBKBGYTX7ieV/q7QiNdA+VE+NLLF+a2IKLgW/kxFjboc6ztTXTXbRYCOgEARQ
qYYMlO9vLy+tLDl+mJXZByiB9EAJ6BTWgI5tGQLWizy2fpMYX0PxuBTTNETTX3Ul
xBPFIEdPeIvSktWzVKUV53Bk6nhxObPgUi6ifhYIbvApWlKG36kR2P2QIdOAoC0Z
7WwrW1lxcbUlr9rWuYcHzTnghn6QfwzTNGISuzgbf2FBqFX9vvKeZl7+UtJQ7TWK
T14S7wyufws1+tsSZLO3FanEHriU4T7b9ss8+5aXbmiBXb3WXovZYQipD1o1PVZX
WiXeMDZeDnNa8D2aGhUjuv8Vhno8ezqdds1JXM8EHJkIsJxNbJPy65UC8O0dYPbR
RYaNKoMl2MJlwvQhD7LFuYNAoI/5Aschvpk9Ca79kvcpAsqEnynUv5EMkLmz8gvA
im9RFwhu1kq3BRzBrQp7Cw==
`protect END_PROTECTED
