`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvaC9PlrKENdu9EaFycgg3SBSXFLVkxiFXIVvUzqRQ0LvuTP47kzRNMNIFKaICfT
1/DnAA38gz14asdBvp4AQCZSxvGs2950QvpmY+bYhm9vb6Hycr3pQCwQpuOiNRUW
evN3VRrvxN1Y+J3GnHDKzCu8Igibsh5w9vJkK/zuyXW51U1brCdxInQdl3dUlBgn
AtVplqNV1SgQeiIJtAnWTWUlqsDMNqmkESedLEsgjDi5/bon6GAE0Sle30wsftmU
Cz9957c9IDhfuGnX1NkBsOuINSjuUamxoualQiibtuxEu5PjCTnxnvpk41Wm1GLR
tEePbj4T9hohM9j10OHNE7llx4a84PA22MtlDglL67RL0dO94UVMNbcOwD+iJBAp
gy+xFuSFt1Km8nCZk7xVLUxkyug6ZyR5iJHP6Z0ZSm/1PMeiKwdaz8LvCLMhv24e
8D083PQHHx1tEjeEaJPyRocoilGsa6EJ8B99RVG6lkjHHoSgSDUREQEOmHqqSrOL
nOE0oV7rFIIVqK49CZU8fvCXVBbSJAT7vd9IflV1Fw/TmMjFwaWWZ+2vf5/EI28B
fHMighy22Oz8V5m8BMRaYgCDOd1i/b/TGmOF4GNRJB3iPxn1SfWtVogOvzmmVbNx
sQgrzCsb9/5qqeRbI4u4MHsDf4lmYt5E2OeBMIR/yJjjzNUaxaTsPdxiSNhfC3UU
W1kf+yfKw1fkePukfhF3Y3+T/miWWxCYAT91MNg3jxMhxD3kdCZWZ/NzzdfjxrFJ
zfo0EcAnGDlk6+/1p1400hkrJ/JfjqxXERldrTcM1V19IRMTUFoN4XdC/JUyL4b7
nxUo2ONGCm3PCW2wr1/hesF66RYwKk7duwrl+DCF2XgWOAPQkGqxyStxULfXhjil
SDLUUuyvDelWl85uDZVUw4biCRpq9c0YCUCJw/fuVoFRJpKBjSPyP82yg85jgMCD
qwONeQiihx06A9c2NW9t2eL5/Blza+CTxnAEvMYTGxinV+zBJT2GjxCNSqrFkIc5
b18stQYa1tD5eUdczsj00aXvsRdJhqM2WzCv5Cj77e7nE09SdadejQaAzOt77V59
2NCBYBbHT9AtoZFYhfnv19qLnRsKNKjCCgesCoQZ57EzwHTbQtXQXDUiOPWoNZEm
A1cffevl7CWLKiZx36KNINgXx74UZUInFsyke9xJ9TWUdrHYy8T20DVsVOK6v3aP
gg2oUXq5s+525sdTNElFj+3TiVtzRHNOhsI3e3kp8f9UhAohF5ydbsAnuuigLWhb
OCRCqgk8TezAbB4qmz52rAnFddRWJ5fTXTbKRGHHQ6DyQpMmGor2nalo/qSWeHWf
txaR/HtPh3OeHgCmqVXShZroDBcW1n6I6zoKeD1zNHTg2l8XxhfmIqQf0Gf3S8oQ
Al3NWiz7YYSrizAgSCixgk+Bd6d8wq0E2Z5wTnjYzw2NXWYbDwqKOZXq3zMTLno+
oCqyJrXhGBUPb5+we0MkIZ2+7LhAclq3invzaWImbkiXJdqNFCk8I5iANIJZjFW4
hhZmbIJCFePgCDtX7CT0Mbj2wCezMtQgENMpWoLBUJ4zZK0KysEbjx4zsoCwL/Ry
TJEAVD7Fty81FxdgxzQlGw9ZHGwnrzCwNzxXde+2bVSQYfxwejxpH1dqEX71V5Yy
Onf9eowAdUtNj8MCt3NKAWvHgPPQc7MlEHqMtpb3XLnIML3pLaxW4gYyG/L3+ItK
j/Gq+iV4upqWhOfBCPRLMC28h33HkEgsXVROYQ0fvfP2MHJYhH3ody+6tgRGuABC
tSGbuJxL3EfIDLeAs5k+7uZ5RJUfN6xl+wifY7hk+7XREHT1GjyKYxF/jjYQ0Vhu
Lb5BXHjDIzGrHEBZHnlTVA13YjenbTfHYLGZ1Bd7gQNXKq1TzNdG2xm/a38yrFJB
zdvOksvUT0l4joBlyIfxG5HbKsm+lQuWwtGD/7rvMGaY8NvvN3oHbxlYL8txTo/w
xokgup1m0c9QaYz7S9QjbbXK+dl4XN0Ex6fDuWXwiQglWlsn7PzImaLNmljpZN8A
sxRv+gfVUga6udRI25ykpZK/mpPrxs1CWaToJaa5XCYpm72s0uebj6DmqKQsmUSa
bQG8exgVBwVtq/dN7ewnjXnZWoSyqZXMCBlqABVC7NKotrZaci2W1OQT8m2QqRuf
GmrvVFPWHSVmL5H0wLpwCz+185dKay7UvUE+Kiznv9RPJUHsVRvrlQD28oflhSSV
/BuqKZ8yuWrIv7prb9eEHQ+lLllc5J1dbk/zb0kJIVTobstwW9yg1dMD/fMoxrNq
stjKHMhrj2gOrQdlqwTHlHh57+ffsx4iEgqFZuWmA7aGm1+AxxJBEENWCe1bFLIJ
4SX67CmtPGReh30RmO/HGfcDQbT6N6okmISD9u3y2THrSd36sOEU6zRE+Nga65v7
+PwAoNw6OhrFhGo6uE3R8+F7a/OhxybayEbpEUljSZ+GMsTb44vMkbOnXqqMaUu5
eDclyMZV4WoOYICqVkGOIApnagxemSLebHvUP0N3oy9dXDOsiACPIerSinS35FQV
8XIJUTHKp6PHb/NcR64RaKY/tOrpiaGK/Rdc8wveex3R5fdAcaL22mTS4O2WBFxn
ag6V30PYLXLzVZZzUBgIHjZpKvY0D3uVwJ0036zKVZZKj8f+NM1GlzSeQfVNYvQM
IrDAYXK9FjHXkOoHCaf2tkzo6etdy6T1OC/3YwVCjrxBrhLGqwPZIUuBmJYVN6TG
pGd9JJQwmCGbWfldRZ/EvTu/1jXuXPESNwFeBhC1pJqlgzRfv9oFbafcYBAKY8Rp
eAZKAOlJJRwKYB+ph5IFezBJlulPG2BbxgudafekQw4F8dW/1oXfaZow9MxrE8tf
mN39Amox2O1r25r9zgRTARi17DF7j1f8IUXZ/KkPg+MCtqAIXFm5F3OsHJYq53n3
fpqSi47w4bUZZFQldZvEiDg6xRuD7JiADUJPkWgdVjRXOSwDXlbnweoSbd8n/DAZ
bM6iIosY44NPcvQ5ltKg3L88pVhNAtDcG9mBEvNwyOdZ6sfWlHhGPNIn5utdjwpL
U6w7ru9mu21AeKJGMIKn+Zg7NhPzwkVtPLq+4XEOQ/8NohV84dqqt9eCPWB0fs6e
pDFQPPPMPVWzbW9K19c1vqnfBRmTDVsIWwLE9C5RDmyeM+XnpIlint/UuZkBJCkS
CWvukZwNeFzovUyaS6xWei0N30+2R9+mmkMa3m0dCSIYhBYOr60ZjBirPPxXeIEV
oOR5eALR7l0U5iarBNIXKNAAqSNEs3J0SJ5qP57Wb+UFWT3QqqGYYCCQHWj4D8PP
sfvpBrapRID0s5dM1lSluDATxovnxe2EOr/QL0SBshHtLjAb2lpA+PVnYpbg1xgq
/7YdJu5bE0WyJvaBpB4SdOC2rUNUvUZKqfhWVzBcD9thHLa5DHc1oSQzLIKsAwHr
AyhZdZEKm7aoYKHv5jIf0+zTkzpJcfSZnwCsfVhY906qzvs7aYAa84uZ8cTwWDt4
dB5J9Bp1wLbbKmYh1gKsEJbjtdaTSZASrX64HED66kfqpYo1gnnNq+y5aUcj+yeD
nhK/XtxK+MMh3I959Fr9RXUtFXt8sK1SH8ffRRdMyuwsPdIKNCplSktuwY0Rdqw8
EfdyiBkRnYGQl1kqnHrl/36w8OFbItO7TjfRpMBky+L8XYYH6e7x27GGU86pUivY
jKY9RCmSgNqwHCF4G0zxOspvYTalX4UNUZnvUSesyZTDOHwqCxtQGTKjxfc5OExS
UeRu2fgfFPxMQkuQd8v5QiwegJpj+z8/j88wdMA6yubNupJqmOH7bBYzYKF2gC7H
piA0L7/CT80AONJfC8dQYyyx3XMZqjnyQbE6JN79NaE2grs0qYl1ALAY6xONuPJx
mmJLHlOFyMi6xKv+7kqR7iX/1EDuutZyIiEpToiJ4/btuMWoGSzYjOV2BiO07Slu
kT8erKHXPymC1F8GQj50drO6260iIY7Ygw3GOCHKWCUdgwHX6IUFlGZLZLvZaByP
MvRV54PeMfC3JtQ11C9wNIsTLgWEX2IoaiGXlnvzIw7Z4s/m2KNE87+6qVRz6YrZ
2h1PIooYUSPCs0KklbiDxlmIcYCqLgziJjkVKPj2bulCglhxbFZXz+ihAguVfeNF
B7oUKaUSNoU7b0jPO28yMlQB2d9ikhewKb1nqiWuLnDT6uqUuFb/+JMN4KXBnEcg
yOS9Va919ASXK33SRwru7OCR1QSAm8GhBT1SlDMLWI1g6H2LqB7yv2/7PaAYa6/x
BtZ2vyfQHESE0lSNKswhY2Q2d5lOziJR+caNyGcpO/I0szOA55r81oWv4wOeUq8n
RbOs6yHWHB1ntujJyLQUkPCnJib01kow1OaMOVtIBdozGU6822aYedSTvXx635AH
iLcpgJFvZYKoTSHdIsLeunscLQbZYhO4IMfYBRiWa47wbDyye6Ok7ZUIRk2s/zR3
Pa+zSON//POedbLoCvjJJZhZ+DgB4Vi844QZwAOYGHX8OGET9H4wdnatJ6Zo09Wp
ZFBYsZxwX+PIXsnNR5n3pWLUfIu3UfBXSVOaNL/+RolRWagVl6FvsW7QQKdER3B4
HDvv1AG7ysUAjSHwvTd4vbD18E8iGbnKMmZwwhBFWwgFg/+LbgjOh6SVCT6oYazd
ENHSS9gPbBNSDrSW5u8Bcg==
`protect END_PROTECTED
