`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+gLVSHbcvNuOGOMcvl14z/KUB5uY7Eca+vEKilPIXQVCPSLWPudiwhL7w90qPi1
U8qzHH7F667k3+BP8EBY5Cvk95RF4LdyA1ukhGlSCuBxnA0tys10VBA0qaYGCPXZ
yuyWE80DdHM4idb4FRIwhVtxIwaxWJ84Vh/gEksNqhXyXd1eVnhOonDwWFywkNjW
zgPuIh7uG8uwIM5++S6THNVOLUufOfngj31TkJWprMpkn2CSKmjxyb3D6V7SUk0a
WyOE2qfp34wTtYqrA5Ah7wduV5a/RhJ2xeIw/jak4RbQdbB3GUdvwhSjdTUqszAf
NPhin2GVQOwofYNc0oA1U+TjX07Q4Ma8CzYo1/Zg9XrXCRwTjVupPu4zgDTBb/qh
lVDbrVuLaKsiBW0+Hgq1NJSEQcibpEoDxeotXxAWJk5WWWcLuk5eeZdpu0msrvB/
/ZKH6IenRUmqkbyizOUa/x5Ric3zIB+4byIjrSM2hpA1oWpAYbLE7xTLmki9RvxN
mw/O9Trfe3RP8z6E88ygfbzKauuw6AcwxZivOOqICB4sA5Uhu3fWu92uBe8xWXxe
K4OjfKZc4xUnWTPpys+zMzfReSu8NRzsSgbsGZIMK8dizNID/h+uiQonjPDOKcrE
YWVn6WhyM4u8oF9aToe5162WhbMBJun6qSTfDN0EzsncwBgUb/WVqnd3INR95HEs
NFD5cCXff/AlXh6DvbddpL3oOa3IVkOHu+bGXNM/BwrBWrSd69hMcAnzWh03/8v2
MNhiSC0MGiiW5DBft45ZWEA7ENlbt369a7hjAuWY6Vk=
`protect END_PROTECTED
