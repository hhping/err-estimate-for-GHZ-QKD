`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Es2Paft7XaTxaqUXczsidt9+3GxTk+74e2iMcst4/0+Ljbg54ghfpBGSpWv4eFO2
dqbJNg6v8OHV6N1fhzxAH/wR+w8rX4kxUDYAncpQQ31DO7XT1L1odKaVY2Q1ZZ3M
kFazAoOJkhwg9vZzO0rACGLhYSEOOufhHE6za/Eh2bbcAJ2DFHM7NWDEW2nNs4Bc
pVzR6MU7OD9pfLOWijTAOQGszunxSgYunpJbx8TX9hYJ2uTn8zIhMfTltcWIDyg1
TP4gGZIJXz03zYWo2OcMC182Eqfyh1iIvCAVACCXKYsID+1cHXT/WV3TcTrW5Sn7
ZZ+81c7IPRX0JfZs/M2etk8ZmOsJANTUdIGQaisMq/0h0ZuiCnzYP8IoEZG+wqUU
qnmwiDYzq/FFlhdasgYghBuoEWioHX14m0hJNN4yMa4n7osA/B6i3Tp4oNwp09rF
MH0//g0375SWgl/ldDbxew76QXM6C/NccPddgcD0unUs+SaKBIYnQNKOCZtlH5AP
r1tYWm19l8OVfh1IbVOVYSlU/MK26W425dKaIJ1aVggCIUkDrEfSsZHSHJ9GXMN3
kytWEdJb0ft1ZcMEaJ/KutmRXtvcHXXLARJDWTyRivglaNUwzN5nfoisjLwa+75e
2pMeQtv/BLJgHwU0ZT6PNPvfFz71rcHeHXaIxRPQCrAYBHPJDtlsHsvwjO9ERUNu
H+lmesK/xOuyhLqUmyov/8S0Jf8yyVe+EiroknyV10c=
`protect END_PROTECTED
