`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUwznkLFUJ6aAfhtqzOiix2FMnhbq+gnAUb409YPw2ijj3gW8rXakSwCkcpWIXjr
9aZq8XZFZd3J2xwo/2EqTV08wy9eSB7gxQAKHFqIKw/CLdfPLHaQ4tS0otqEbps9
kP5U2v1DwxAnT1DKYCryUtwoa/QMItSbtrELU6cQdBCsdkxVin/H6dsm9JMxrwMA
VkuqPppHc3VPBXHXB70d7MvFDhm6yAHZsFrecSTA3Cjg9c23C7bbabmxrL1lZaRy
GZ+nbbNOCOQ9ztjWo0eKK2px2SU+4s26h0Ru7EOEVoEK/WxlipjtwK/pXQNPEebG
H2Uj8SeLZ876qtaTcPAPi6w/ouY/mMkkpGPVA+2NyV32fKCNcPxWJfXnlUEqzelk
GYHVxB4yeqeF2aiNJeB4pQmkFycRw3MqL8n6aYM6+LUUnDmqLUAe1XBerESXnoiQ
zmdJbUadykLvND2BHaTXO/x3LE9BQMOCpRmud8OjDKvM9WoYH2HEXQpPUtJ32tJn
TC+jvqQFsQRfKy22di93IO/JydCRhVpAnJgROpZ082JWq5QCoQVT5hu5neMr4W55
9l7yNsI+480XCL5tNc/f4DByalVoHToG5h+PX71hhHcMbBFhSUyw8OnofuWkQ15h
Q8V2+ZKOYUgTWMf4Z9gH8boOsnKo09CVwF/WKrSvX35H2YWwC1vydzi20xd93RZG
ABQkiR+u9WBFk104JxKcN/iu5Xjehi8P5fnsDHDKF+B27cv/3tvS3FbNqTo+/coC
4QXSwets/j+wVVqwIu7HNg==
`protect END_PROTECTED
