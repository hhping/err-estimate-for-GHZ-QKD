`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pqRJ44hV3hM2ry3f4iUiOMpxWh5tjE2LoEL5qU5Pp+fnH418LamW/GfFIiH5cP5W
20b8olQ0VEzu/G14cmzZg62R5npOJZT0pcrAN7e0eMnoXTRRiaQ3phe6Nd06M8s/
Zmph9tHnaWDGl/wBfBKXIgD/ycX+LFyp+0Ls4SlExYzwR3OxkaUiistHaWBmKCaj
DZ3USsBj6D/P0S/wgkHVZFSvqpiQa+sx7EMs5mjm9EvMB3Y/UrNrb3C9xItkYuYg
CpuEqi27y4iGk2fYgXNs0lPj4eVurlPs/M8GV2zLc91N9XqszhTQk2Xea9RQy8/S
iAQotFEPz0s92SwelqL36ay6zrFqaSy22up2ePpbAYEKoUseLuJrwCD/GZg7Yohh
NHF5UMUd8UR1wLu4b6fkEzD0AwVre0sGDvL5/hAC5bWeY9fJ+jgXFwUG/jrco2yj
sv6nxokOJsHZC6Z8AZciO7mQFs20Ft2o11s7FPW5B0gxGBeEzRYodNpSKgvGQZJm
J0U2lo2BpRn4vn370Ok/PeWRB+fVOmnvN2hSBwms7JA6MdjH7W5pLph5mLKQAWqD
w8W/BlaNiJ3Kle0gvvUwoMBaTjuxY61rOD3Is4WUevSAFYUYIwSF0PDfFtxWk6sc
G7lPbClUyLmwSZAyv287W6GSlH6TVwC8D5Wq/DyjS1KBR6PJ4LHoFsQjlj5G9ujz
gcRYylbgU9QN/86loSxmu9fmTeDjJsfoBB7aA2WPLCy2H/gjRSPogiJKXjp16jLO
ZK4RngLAnJbZj6op5pMPMyw0cF630cp/NIhrxKC1YigvZrC3LhZGKZRd75XQ0qEb
jGFkpK0OjBXlLCYm4r815r91j4KHtrMEOGVjb2pViQp0ZC0PDF2nU1rmyQNXe1vN
bJ3lg+KGxTO2g0T8NCl3Y1OXd95Zqp4i0jYJEws9TR+X9fBDeMiZ7U+eIg7aNPdj
GOSUuFI7KS1EGmKRCYw/FHy1cBX2fzrh1XsdH2c9eSok4vWYN2WDqPOWSAl/8BPL
h55EXnkq4HZvn8Ng4ZPQyw==
`protect END_PROTECTED
