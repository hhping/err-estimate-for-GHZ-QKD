`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6/t7IHXNRBse78cnGH49dGboD5F7eeTp1v5DKg8RQBXjyX0rMZvcoKOOhjh/SZZ
ZGnM76rK1GLE74ii1rZLTlOiMKY4OL37KMiG6rA+I6k/V1L7jqKwk6jEAFJu/jqO
dAsecMbBSmbPRcKzuhEjl5KvlsHgz/rkfB51K6vn+DaYapQdedqnAbayi3/uq37y
z3v8uFiW2kwFHW/GIqNdhssX6jtN+CleL+utCQAqvECFj/L/a7DExcMXQGxNqDWi
xCoXXgKSsqR+cOm1LpJSn0T3L7zADh2ixbHYk3eykNDjnIqXBQFokSGy0I54bNgT
YRIX8SdTDJO65X30/Q6XhXmR1Cx9NthDJhKaJXU2UE8Yf/dhemGVAUW7i8T3sL8E
vcHMa4Z4XJlERZ8SQCr9ru58+/eMOw9yHt/RFWE3Jx1gSw/02AAspFpP1pM4m634
cP7L4J3l+wvrdjY3p/Iru/DZ4aDz+x3RF+l0CNMhJkATHPrDQAFDESusOYM91kQ+
+FTMLeZi69+IqG6tzwxuxuOV4RzDJew3nX68l7lLv3x5192raodYf9GzYNsSeWb6
/sVk33s1TxOIOULDTAMIV1/9zX61rK9X6sZ3Ax2y/Z6UmnPYLPF2PVqCfj6kR+4E
DE0EVcs+p1oIUn8F0OzvQsost14VBdCMpcLCtnZFl24z8dmE1XVjvpuA+2XEoT4J
BTFGanCwBSPHh1JEVfcOe9QmBAxivxTAszoNwEYLoF1CLelFefQGsVf3N6nQLfz3
WBAcrlGgSoqjX35J9OjyHAEHcePKBZS5LY5NnNaI7cEiwvMyEsg5Q0dvYdOFwdzy
vYzrIasyoqtgIRxRFNUIpde5G8jRpw8coJHJU2O/MJvpsAmm1rhbMWuSIWefpHut
PY0fDbkpQOlEpTVbOZDS6+BLbDgKDQP2EniaUPTXYdjmgED4pn3L+oAh+eCyJQzc
/abIrOzFqsiOwDwCZkQ/MiOqd6FizvjzC5mQSVjsLKC+k2NseK1F787rShMOMKlF
2+mTUMK8fxtE1Zog+Mq4niflMz3DJh2hOK1IwN4bA+r4fqqgJB6jJn1S1fFU2RLI
R8sKppv5MczgU9iPOa37TViHyACARQ8om3e7Yt3CHHuu5VioYJjBCSHFmrks5NRa
KyUUJNT4PFynbvnlqr2rS+758jZb5h44GJfKLtpWfpv4phDq7bh5Wo9kSFuHnFmI
J9NEhXb+ct24u35aShy7RdpWqCs2IO4q/6yjE0C/q3P6jcPbHMpgkpOZbivUFgHx
y/XBYQKz4NIcSgGBFxPkfoKtxWBgyjAjn6wXuNMUl+JIjhKKO5mQkfZIwi1KhAg6
9Rl5XEBd9VI/aSOvnQvKiUKj8b5SpjvwduQr/eEJKbGkw/DgDnnAUQ3NJqpoh4Qf
p895w0HCWDZLWgu4fmmRvgjPvU6LsU/0nnPNPcEVeIBL3FsnSR/uwRMizVeLWleH
/Jxw3VPWlw42YB17ScwUf9U2Apglhj5Fn+xD9bQZEA4O9ZmhbFBHlkbUiIUhdsJO
PiyT2akqN73idS3EE8bMEmi90zmHjveLX6lY+5NPJTT7dHkY/Xw0uxdelPKzUy0k
5ctmJV0hZAsgWiXrmMCok0qXC7jnxF9e51Zj9STfNvSgX7llYyqaaf18zXDhrqeG
JA9HLNKr+NvCTN54m+vuhGdiiji/4j3opLTGnBa7DpJX0nE52RylzlX8oPibuSSg
W5NDvtEr8EXCFZbSFVJ2eQFhIZ0R9FLTlf9fVADYCezLyZ23EpAEldREB4HBU+mQ
OQueDsyn86PXv9c62ikxq+hFWEW79na+PSBufU/AouhHfhJ2yuo0aZ3U5bN6v6wJ
Ph9xRznPPb8pA5JVv1+jrF7VzWZkKW+nPmGKauE2DiTsPY/OyuFxhRd1wsCoZzlI
o9ry7+HqU5BhcVflzHX3I7LWCh5ls5wz5rsPvGeWO6YV0MakCVNDHkSsAkCsU6ww
QDSKqIQHakuUatdkSktQANQzohXhiF1bgWtY5EIcznSS5t3+dlSk2FVjqJpwKm+7
MfXY7BYzh7/MxhqBTO+eJo7x5Q4aZujrfOQ3Tm6obPQ=
`protect END_PROTECTED
