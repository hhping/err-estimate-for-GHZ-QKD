`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67OYrGUdUwleuS8XdoToMDf353Z77V0hj4AUEYGiG+AIA1MxiRiIR0r57sH/x+Ur
tyUj96Nt3jxgMbGg6Lh4Fw0NrbtiirErWXKXlBkJkWcDSt4lOno/kOjuJ/O0LKZp
oZMpth/QCHpxmpXorV+ANPXbUTSO/EG67gbTPVVpj+UpAFX7JIq+0EOG2pLBznO2
/miwadpKIl8OY+9Udb34D8fVyFEz/7NSGalcCY1OuNqJTWC1O83gRwv7LOBA3i5k
h+nt58wX/4Z22fihBy1nG4Vr+uf+IucdgevojDnMy++TljHtpkIoSuMt/NAaWReb
dEZKPtxBNQDcZIfU8MlFUJrybcQsQQrwQfvDLCtkXO0okkanwCBtT/r/wNW5Vm9n
KnPpAKWAW/I3FX8kL+kiU3Hxg+rFpriNgADvSuFJ8hlyV5lgp2zurWcJWYGESINh
VNBSWm58w0ZIc3Bn7wgOiG3J1C6gebOj9xqpp/8mL0gEYDwhnhC/GYfotIritbIq
PmiFW6WO5Xgw4/gGGGoh+eGYfnB1ITwKOqQ+6dM41hdtLYSo629OdThibPnJDIBX
DuxPTaknJlI3H2VskyWpiG2iovrBOsv4SY7vwkN1SagbGhSPLOCe+kFHPtpXJVkl
9DtIhoMzAiEg7KzjzXW9434oJohzoh7Y2iYJ9ddT8HFBgVHBAMzMQiSRkf+lEE5s
6dM0AUqWo+Rtl7g6fX7begPurcbHbbC4Dh3g54Rj+pQMhHehsR/AVzOble+hkK0D
4gDX4eKfp5iKFZXsuZukUMCfs2itzFDcLfXAgh4ACfAjHDMEeB1GJfzLQhRdRO34
s5WR0ge621uTcopT8jWAeSa2UAnxZS0iHC7FduYF7nSgNQBA4Q5ZMNlD2u4WFYDL
VqfL1HUzzrHxUO6V36sK229hNnBnvlG5O/uKfBvbzFS4OSH+4wFSxIWcvaEmEMLT
DbkYd7a3wdhSMt3aybiQgAlHkz+X13XVdQHH5iy8lLqIhIOhM+A91UOBbKMQfqF0
VvNpu8vVr6y1ukzqa5/an4TQPudfRxI3YZbN12c0dYZvwA169CQ5SAxV+trtlQ8j
uv0MdU+o3bEXh3eZXkVd+TzvI81v3qS3WzJrX4qy1Nu064K+FLrHdFcdabqUbSEi
JTCdbCZDzdx7etmkwXJ9J0sRVanx2ofBOcvah4ATkPPRz05pfp1KGDfPUuLR5FmM
RKIUqZeF183lNtA+Vna93D7Gq6+5IoMlLIIOw66D+OHgzjDsnj/Z99pD5OX9dgOC
+RKQs3HhnXIv7/QtWapKbBNnO2tHYIXnPVq9sFHueW5hbLxvzcbAtsIp3CdKWfp+
/Ixrz87ryxi/N4vtg4pyfmhQSw4UDGygdbRIAERtMwAg4JJz/RuaXA5Wxh8g+49p
8W3EhXtjAwwEgYnb/0gaDrRPk2r02fQnMBLJ40lu5RTTb5oOybNE9Tc0p+54RfEa
wTBdxDoiYwuhHs8i8lcOJGO6YNfBvmUn9eoLpBjW2MwZxJ8gdvAq1ObIkUj3UR0H
ZPgKCvDAq6ZkerCm3x+X21C+ORpKh5q6yQ4d7BnVEYuKgFqPjE7Kwlwui8OIUq0K
jCc2ehwLFLNh3jdQnW867U5WF5QfVQaKFI1qSdci3Qkoj82JDy4XfLvEX5io5xw1
fpIGcmYuJH9kwVFB/VfIEtT4zBxyxNQc+Vd2SGD86JM//QpIy3+6+BXIJVu7RoJx
T8hG4W0PFo4l7DydPM8yOYeP1TOCBcve2xCB8Ntne1iCo3VayZ9gNylmL2YQrjAa
FrclJiEvPcosXmdYO0dXKKEyEJftJ1/AlmTSrhk76+yBZWXkDWv1VU7nbp+T/fUQ
7FjAaw5MyIXQNdhHIxV0uGZeEtyA0mgWwk+r8vH8YmQHTFzRzRoMVtw+gN5JZS16
w3/+EV8rN4NE2L6dML4dNW72zG542CoOrf4Fch9hP6gzTSsVnXgACMQhPyIqiAPG
ERll//vPGmKshv/9Y5qadHj7FLQWaxSSvx2jADwcHlIU+SGUUVedANVPlJNACEZ7
LocrMwiwbsGn7s6X9PdDwhbQ2vsHcLvrpEDWp5c3LQb1a5Z6yBMTACEJ6xGivMoX
EX+D4N9H1C33fa1MED9loPidQbMktopgkQFyFMBHISajIlcHYH5ZiS3eF5DAha4S
CMYs7jKYwSTivOsJN5FTIJqfDvm+godI9z3NEmNStZFwXmMnQ/hh4N17v3oorPKF
LYzP6ILasL4GPOtdEvsnpIVATw/yILWWnERWMGs8ch1+xHOLqNg8XfrN+0U3x2I8
1F8gOtoqKmBiJHPzAXvgpGPBJ25i94T+86j60F7oEsGa+FhtrFO/px6+4ozdPHz6
trihbXPx8YCj/3qThZL/kUmMmlN/08qcz4ki/Sa+psgLeTAAx6I+tiKC78kbwJJg
Oi4P8ifJduxsph62xIetlIRO0SxZP53tQUqpTQOTtd7aN6323noIqcGsd3pejcBq
XsQkfOsjbFCOpdpTLzY3daySZ2iEfYtZd5uk/QQXzMtKxZzZBMCt7lqd/zK/IFJ/
tHIbRhUlTAsfVtYO3TgAPi8AvDYEtrasxDnIJKz8HIfP9CdyvSp0zsuccMrnrxHc
u0yOXcBLZQqdujww+cVLlSR7ADP/7sctADOzRqR8+QoVMa+XrZnapNIookB6fIpS
3tF4KVMVSvgXRPZRJyHwVq1hxoth4lJ6q6NHGlwohQjZIzf6L/HrkhSGhbTXdNBT
W393eGDWD6bByYQgQOl8LA7SXDFQMcUuErT6fpcrQ33Hx1JucuY8jFsTJLPV7tvb
Mjc+kKmxvC2ciTOVFAgRHjhlaR5Y8YVULmogAZubXplOPkrnSES0g1e3ABqLK/e3
BSnoW1Z96c70ZFH3ud3Wl1VG0u/DKcBRTDCG5K/vTk2AubzghoPLkqogW2Rc5fWU
tK+738fqeqImR47FG4/ujtG1F86zD9qhs0iXh26LxaH7jmjDHknUIpZD6E2jRcqC
ZqLHmbAcpVPWlYppCKvl7gL807Asufw3prccP7yoyxdafL52zRF3b4+HaeX9dfHF
yG1oAyISpcchiIWbtGIk/QJ1b8wIUSQ26i3AkifAH1gTO1yyBTexOUAEsLV2E2hf
WYWsURVGCAKSHN8A0FYSE6r3CiZG/YcV56AgEvTkWseZtQppHBMYGiaz5K3U4fnu
AfXLkXkHtdjLn86OfwbDkic8/kXRaj9Ar1UQOmAPB438V9tOIFrvOP9itmX9UhDn
cLOVKDS6TiqjKBJFm0UVyqP+LlDWsQGH1Jsrzn46ovzmiU1XGyEFXDjE8GI7jwMO
+NAqi7zk2I2XWOeI6zkA5myV486r6b2xr2IgSSlmIy7EP6ojqkHU8m5dEJxuz97e
tlChjSw9BwwphymEIOvdDJQyaGuemJxzVJ4APGJszLoh6cx5ohq9NQ0aws+ZppAm
mD3E1mmd7DaZdIs9cK0bRUmZzdzzZKBPE+TwszDyPUV+KIziCsh3nkiJjDwh9d5n
0yYzRtP6Q0krm7RC84D+PBg3bnZUmqvGpeg6V4ticGgkY2eed4+EwLlkNSbuteFB
BxSe+SZ4CKch6ibCh0/zfwNdag6e97YZvFJsVCOVVINeDdjPbSAJ3Q50flW+Msxt
xf+wTZPQBLHsGdKUOlafVrFuaPHv/Bo62nb/IjrzB4JguINvS7eVF8MFkvE4hHzg
nuafaVeD11baAQwbMd072y2TNfdOKmZkkLic0YF+Ak+cY0S/dnUD2VR2GbhDFCet
qwq+pkEyTatK0jEA2F38WDs5PZrAGlw1ttgitrKMZXiN5LwSHZdMPqOUht6bm9/j
xgjKjRopRfTLjX6+eRCJKyhyeGiNSabhiQgru3eMxT5AcIVcwE9Q+OnYxjeeXAcs
bjArpyC80NcObBSZqeKsu7gOZU/Gsoppg8YInD1CuFUoEM6AisipaRdQBOhmUUpB
gBF6ZTaSjLPinumFqq5oBZLATYt8AiR2cRNHPHy/0S3FF+ncy8SESev+aup4w8X1
ZVJ7xDhZE9tTAEXBWoKEWPoXjFFQUCv52IhF4I5aNr+DQziiUn21hh8r6g0MMfAK
r4PHbo/SvITgYrccTHn7IT8uTe595ijo3mMFyWGjmJQ9YilJ83qMUtY0xR9VqH2E
NFOcow2yKnHrXrtSQQ52ndGN9GVyIISDVAFtDbg+UgaP3LcVqVfj5NB2dkHpwLZP
iTbhlZVdTNkRoDj7gvP92MepHRdDgL/FlGiDKp8zcNZpuDY0z2Uqet1eYKPMXA5Y
Q4PgVovvgRIk5YJCFLsH9dGfmJ4O7cHXuqvVs3g46NQHp0/dHchwFOCVJ9X60+kC
3COO11hopUAYcSMIfwMRJJTZKa4mNsYiBwyCI8Bgor++hR1smZMueRejyKKDIc5v
wMLcip9PIBcu3jQQ2B4su8eW4F2RY9R+0A67cr3HlMsU/Zurxs1fj8QZKbtfWjqa
dcI5vqu4u5be7OlvlophMxtGw0OdgmHTtf+Pu0VNgT0SW4Id7Y7uDUtZi05ER/7z
vRTN9wTlU08ddHDnS9KTwg3bPylJ4yMSCjKA4SBptA/D0XlehYB0Nf1Q+tkNwtp8
OfCMlCS6cQ5dcEmZ3P3uTlA79FAR431TVPI4OiiOgBpCDN4/QYGsR2ZL38vsn+vz
aV1t5PbTiFrQXO/j/JsG6x24K6UxWjibicyUczHqGhc56vt2Z4QSXAOH2l9MPNqb
vniQhja4/fxKxAIHaqDKNNQ1fAw4tf4Y7h1RcS8sWA2Pm8PfAX27pIPggyBK5suE
a0Mdb1Zo2wpkDFX30iKX1xLA7V7Dg+/UVhCzRjFTDOCJssgz0wNsML25KUXIpXH9
YvmGRvnckzRsxjWW2s9fnVBHKpm6lzZfCUwFHI+2Q+7mHe6sfBYhS51AMGrMG46J
op+tLuCBHxhKY5fZPa59x0DJVvTFBqq3PoG7a0PshfAGjQTSM4JsqkcaWiR8UOxV
bVt1gpuIPwM/hR6LBlr7LoIelPSu5uitkWDeS+O7uS6EjIf5ZsAuHP+CG+3litKj
tvXFL/S07fLDY3QkcrsWo0WDS/sZ+woEdvBM6a/ajrxjis3e3jW3MzssPbo04GCQ
5PewwIh+NY0hHRrHh4vNBNB4biHS1zAvovc028Y4jyK+gc1mrkPqExaLtXxmD9PH
RuRdolNuJ3O+spHrcUUji2CVZQf8shHzkIyPZr2a28ihC/O49Nch0Enee1uFR92u
qyyUMpk0oDcr58DqWnBGojM3/aZEkPree6dz2n2nQqCiP6vHeeUFyGbn1qI+PoJ1
zoUaZlBKYsYoNV+7QJjxL9Q5wgYCt4p67FScZaojIm3xLq1TcX66c/BxSqxjjEIa
yhGfvvD7WHgKDtJvW4LZEu+Kx/vZ3g2+iKTAWplVwJ43Fh2zIaZjy0oRVDhPFjMQ
BPcLJwUa0IZKdJ1Ktr3vMXa+G1h4HXpS2Dbbj7xJsvxUAcjWHAcLKm9AuNscdgZY
/cMki4FM3jAR5b1n3bEigePfNYTzVHWCTlt5aw8Vf7k/JenLaXOrSiYQ1WIYRyuP
DlzhaZnDDuDp/SxhZsdPjyuI7qzUhHtpD5ENaHA6T6MA4uRDYSQ+Qrm822Pb+0E+
68naSx4cQkFgUeDv3bWzu3yOQ3EMKdJVQSx4Kq1VdHQrMwfBMvp5z0coCeIWLpGs
sowI3VR8VZq9uNYJZGRZrdvcccCGSk2Oj2rvR5jZaiXhcly7naydd6QzYob8Ig6d
EQL0UznqbO1lDb5m26/3CkeSeNH0EpSYXO0ie1vvT6eS8OhUeggcrgWOA0LtWGBt
96qm2XQAWo6pV/DdD+ga8E6J8vLvlIaHZdX5/Py05z7klZ7Dzbd8YQKplwodKYhG
i3C/Jtf+VroAuuZB5khZATLDlA+dDsWhqFXoCmE93vnxgF2iRae05kqfI6qTNMrW
DQmGFkf1JtBExZ5sX/fQSPIsOGqPh96XFONuYli+mC+XEl1xYew+zViZfdQgNZpx
EZqawxO//xlXlyAHyPlTyNTFIAkIG70mGUnrWrvAUGsMEbgePVkO+RFogUHKc+XD
NeRMMDdcxfDQF09wGabtV7ZHvusGjmCn8+caAk/nmqXIDx4vf8EHBYmXnpXOPcs1
X80cDlDA96tHQzxLbfw2XcQhl5r3uN4dcSgm81UFi6w/nHHt1QzbwjUJYd9c0jcN
YvsFHCxV+7NQ29HxYXFL2H4iojONAl2w3oiqqxS+mVFp5efEvfk38lMljV9UAuO9
9Z9RBD12GPwVvhPuZFkZWHPOb+H2YKyFYQYyIvTnwrWdP63bGHcO0B3QyXSbvewD
kIVZ2eK1dAYFhXWk1PhTFUdEOBqUEj+6vVdEOLOWKpmhqP143q/XWGd8bcJwYMMw
9uuK69RfFu3W2jLVQBr3FC+Bh5cHoHWMd9jl5VWkW+kFy1FzAYOjQs7QZ8YqU0Jw
+j+MiypOXTjgbGnucb25SkXg9HCxV8CTktj4ZeTAKQRbRd16UUz2LztSBlaDVWum
nEf4jpZ8CLIBOcIaLyifbWy/QIxVR7cza8BEmV3XnsIFxXLvvfKDPkNLIm/UZz4D
mrzNU1M4YPi5/I3n5x8f05xCN8dYSfIJFOvSUzWhcrHveXpp7J0xwPtsb5mN8qTe
xF4lHYzUVBEhbztWGmxCqXuWa70HLnxgWbS8kCEgPSCyU2HPL1BQm1eP0DAYTDf2
JCugZnzYBKC/rdNhZ8XADldxzYy6ZHwrEAJBejGe1QQKPTC9WEylSB6Dn6BGuT0Y
WDIfpC9kSKvE2pVwhGkNRLgGBSiwDf9G06Dt7i9hR9kK/gihwQcxG1hOUnLXWnlt
OfCyc/ADsRzHTWt9A9YeA0kdNHJbIbNs8eH9qrfta2MOI5DGnvbKDPQjKYO9hpLR
SK72AU+hq52l57q5g47z3aNAi9AjLW1A1qgleIBDbgCtpeHNaHdeCC5wk4RoGyVr
B3OiLHAHAde8HPv0Q1PKAha1JrnybKotelFeYOrI4DLvwsmrRCOY7CtRiZCxeZJ4
LSKkg6kCDtYv2KSoKLjdn8bcGyF5kR6rPD0i6wruFTrUNE2ppkwNiq8egxOnmloX
7CuuEnLajxa8hX3HA0PAOdGZ3vVumJpw/yzpzIt6OtIvsu4uLrZpkm//HS8SsFtD
GFIqGT+mxJuscM97Nrnb8XzDI10wze64upkLV4hl+Mixzq0svk0iS1PLfKbDuj13
kqOGCHsz9uN+K92FqvanSdB/7wxdejn8bImS3Fs8y6l5It4yWBQleA58/TeCm1Dq
qoEKUURd+F1+lt4sgg3QlaAbw4hHhAf2O4pU0woKOc41PvgV0B1EREpQePhXO2gw
IcOXQiTNRYJjeuMd4amTgVzmMwAw6OH1M+T0cIMEt6RYGnTNvl5X76XjaD5mtgVB
afv96mZv373psnNwemQWEuBLX1ZhoB6MSX4Zo+W6DTKpSpY/ANFsd9yLi486uEMY
88P4vGlMt1s+WxQxIuNHq4mceTcXhANlRVov7pY+FAg69LBXdY5DYZw3oDdPGW3W
iW8D4fmE3v5MSln/bPAymAeneZmv0WOTPv7AimF7CClIVx579cvoqHseVjAvWNQm
pWCX9d0ljKQ0QundNysHN5xo6V3NzOe2nJyik5VXjLp4RyI53sdYr9cN0SbvbTwl
g5zbAN9Pvp5/SHz/1cxLvtGCBaljMtaBGs6KVWlRhKwX6tMhZuem+0GT6YxpwTVI
X09nbPCsFgxKyGR4bNqBV+Pu9kG98t2+yvugCykggBVNfMGaXj6eXM0GB6vGE1K3
mrxpId9o2unEV4rw53vZi9M3K6tIdLjZ8W1I/xjkC/EyNhWBMANDy57peAaj7aJS
Y6/sYqD/UyBbxBsH1rx0rGXugQRGLIuDFz+m3BRvBv2iqkhiZn/MEs7/xFDVBv8T
CenRgnXJRwUZugme7EBbCT5K60mWfXDjG0Xxq37vEcBdKQaHffZrv+YkNH/Lp9LP
CLs2BMYXuOkP92H+zQlVOWCOtLSL5X6jEqc+8FZfA0pYleBgf2fFloCGS6yjHWnq
mUIflaR6uKwhTh6kGROTRFONyLmqgucZxpvnqXQShwbroSSNx/aVA+1EuhcdOPm4
ibM9OAI1yHChejhaVE1Gi89JKwvpOKjrxzBD3Oi2rTF1ZmeCZb1V8x+9WeT4Fb6C
EiFf3tViK70GrpSo1gl8DAQyOFXf5bjpKCY3WqHUZJ/ex84L/dsnq4gAv+cxgvNm
1t++yT+lKMBnbFNKSAcSOAES0J4HR3TT8Benv9uT3E0yrQusVbl0i5LnRxl2k9hj
Dt4jJZGqEpJajguFoBVJaxKM0n3pmWEH3f783kdv8epvf/D096qmB2ypKHMqRPB6
vzxIN4dwGLiI/YQTopdhyCz9Ajgk2JFJCtfmiZVpMp4fKEQkU6+qz3db+sJmT81G
kg6mTru5FbN2IkZYBnN5S7PPxhZYCsitTZzD+xwML22StFqAC06OsB9tPgxpVEah
9dFcMGoyecenrWofEDTfDL7TnrH3etRtcII00NxvOGzYjOHt3i0k7YI5lEB+mPZM
LMigYHAxHEOM8ee1cDgpS4BbuKrTmj0ElkFl8tU4RHionsFGnZ4gQGNvBrFJzYRI
bSlckHGeh5ntPV9NXtVAQ2ZI6/Xz0i8zS0yHo64dzzCE78xJZC7MMGOQFaNQRB/9
K5MnMotx5a+pQBQbL7nXwC2mjv5bFeTncvHCclEqI+nmUY68cXZkCnCudiZXUwDg
GVGniZZYL2XYMYRV4UXk1cYrumqpPnG3CFj6jqLuFwT8Oum94Rkfe8pdYItYzun6
oG4bFQJA37dbKTrWFsnTa82dKd0Z/F/tG+VLcxk0DF4QDI1QIf1Il+9tT9XkVjca
Z3aRBAakPe4Vy39tMOo1Du9zjey+H6t598Hv9lF5yOtfiHhxYugNfT5YFjK6j6LK
DYKhOvnzIgmpyrUTmgzEeqWOG1PXq63S3+LviyowmHgp+7UBaigmiyom83qYihrG
OqScTeJx2VyUbuTFoZhfEd2Q1KvRdAG7/cwnRimPXy9uOD4p6ZacAm5W5I6xkCVN
zySIsbLATZxZ659RAo6j1TEwUr/nfZgNROOD7xctSObjDv7uWCcubTvQGl9YNH+y
fI4KWVgjRWEb4FJOCw+opJV7uxKMJY+YMWlJ/gHeRJ6XUX2ih+iut8SqGJWqwTty
GqwAiHDTWcWQaxzyUCYaeLW/AOuPzNbZV+SsU0AtOiugtVPMqHteMK6CAOF144F4
teuHe3lwHYAO4I0jIUiBeZhgi3bZ2NvzhAvb0Ub7YN+nQBMidqEsB1jfZAEFPtTd
keyjJxic0q2ltEtFrlO9x2Kdr3fT6L0mqpg+o2vz60leZGT5OCyr9mcBYNuXSsA+
u0g1vsnt9jCdHn/I3teEZwOJ4+ab3mWz+4GO+mfKTEXN9Zuii6oXlctaGOWAn3W3
goYSGR6Lp3+dttE6BGIY1WrRjxGrkjQMDgSNVyGHmOZSrgGtYqwVSCUdcoz3D+23
FYiDAF9u+JeSURuOMISIrmlXTH2ylUgi7KG6ipnZdGZus3z2d/SDX2JSOasp/GpI
W+Cagso5zdL0HNPMwsR2gd7pvbicRnZI1h8r72qUWLo/X/iSo2SW7Itn9gCDmyGK
VpjGtbwFUUH3guvYK+oM7ESVn5c0GVtB51peBgY5Fra5Bgv5emnjKcq8UODXnH8b
NjVqwwZ30xsCXkZQwVnaSNthRtjwmh3U4r1P2fNw12vVKyMB1rC3kOkCRTZ/8j+p
UbV59JsgUwVsCizDuLYbc5e226uLYerbkzhB/Asl63wNoQO4Xad4F+O+EJNW/MHS
v92lg7yrj8U0S2vN/QkQUE1zEbrAIQ+lwoggoliB1YtjmNKaTD/q8UEQHos9pfFE
L/XkZuWg8AGBUEFtdzr2odhYeiE3W1i/lDY4OFyRjQW4pCuEIZiScn75pjqu7jb0
wUPAzTZ9pzzhhqJM9nI/Qd46ZupL7Zzhd/se3la7FmhIHDsGaApITIPndVhgbuqw
hyIbxVs5o3dNqO7YSL/1WDrZckl1Ht02Bg/tMzSlEh0ZJDn5+cWRezcHnmnCznsS
BTmrfNfqI3tYSm1pQVhTfn1XolLcMy6nzgLaCIPmjqVmAeeJP7JLhawe41tyvLxY
qZ3axwaglI+LGU5vv6wgL8dbJ4JqOWqKJIRDNBkSK9XBrNv+gtk/Zs6MfOzlgt/T
DS6uWrmGR71fkcuQQeWCMJYGyTSM2R1b/DkqLTuxF08NJDjGaiezAX4PVgrcEIQN
ORrXndafqW5dsKdRrkLaH3qOahE3ZlLeefuQgfLhuyz9+fR41pMA5KqGJB3R+6oN
hYz0whHVJLL4QxPaDGt8LV0DkNE23NtozN4O46nYY6Us04ebEUJE+/HdHLPIAKPz
NR9a6yvLFppAoKTs5myAyPBy1a3DJNTs7+F1kqatmV0cdf+PGSsFGl1W/CGjbTZz
t5fsR2gcz9DOxxhob77UGXjteSLQkRe845nLUaaX+nap8woCTQKag4X8tgNfC/E+
K2wp34lO7yBUb3u0+BhBhP6w7CdoI32zuw9yl/5kbrPUvLwe9AINyRUDaD56RAIF
u/CJgcz1eR6T/ahznLTZN0kb5tzxdunfF1QIrn8GY61tKt5WJcnzY8QhQXNLbr8F
ViKZtAmWYS6/ygg4U+EjTlTwjh1G3XMmglIvJ+prgFKDTrUylY5psGuyIDMDCBqx
g+PD2Y+YmUaU2SqJKb3ABaP800Wjp+xgW1rJ3ebTh4+REONdP0EdTdOm8/iJ4RDm
DaxUX04vddrRgClpv2UeH9s6YJwJGRxa7ca0Nv44IrR7U1LfjHeXNvjxoSmSFqHg
3cRkqEcnK5RLMNxTaKnxjxrcuJhDdapd791ICR5ZwupucQARK7G8S5ilGppoNGl7
mc6dLB5ntKPsCEFaDkLVvBM4FnyANpyyAX8KYG56uXXtcg0me+2i+bpwuu9lbrYx
3ou1nJSWX5BIT/SVKDZ897ybL1nB0wlkQGr9QyPX8z4YCaUHpK9rOmOMRcjCAacp
kONt55CkOWcu3evThv5bdEwtmCvRQzkf85SHrp+OsB9kKx5Om2vdznI47dDl/KyE
cz8dPeWuvG8qmysB4G2UBRmrCjDT24pFHM5ZxlePrEmaqePGULhNOxlpZ09FPBrx
7LkRJMSFiMUtTDKYwr/BcCszGZ6rXR6LVwcY6fjPMP4ZnxWZ1IjNk4lSPsHQpBE8
C9ogtluiZSelsW+7C6itVnz7zlzD1OR8WahoLH1578b3mAF0rhX5Xe17xbxK87tw
yPahbMouxKQc4xHguP5AkWiM6i7e+UyC/PfzkgaVSQfkOogi9kPmIz19yPfi0XZy
j5e8ga9qaTt5/gSNMJ+76ss8HHR96/a3McbeyRo7Wlg6wrmSmxGEyzMZ6cBTv3cs
SD3WvijhL0mz1EmeRN/FVEfh3r7hsfOz+ZnYEchp5uR8IRDMF2iImr6KfTZmVNyw
B7vzQbE28ERaX7VJgAsJq9ldxUZYEyA0lfk5OXOsiIVKwkfDk7FHqCFBiIrHniZF
4lHwFAADPEGfH2ioWhUnZhaaj4KKTYU+2wjzQPxFZpwgaRSUPGz4YZl/aIvqXFoS
NRYR2g3TRyH9ehTkG+Sn4mvWc4UaarV5V4YquKpEJCtI/aumn7rePO5nHA7qpZhr
fZ5AYfX5eanYEiDLbOL7zMTPZDukiEnY8dYIWUbgx0uIgahkKhbklXcjJWpRS98g
hMjTVibva9VGY10RUABIuQpenjAzPbQYd/hXHC+M91uJvHOC8ghjnBJLQigUr+Ya
3MFh+mmu2fLkdCv0Ltsm7zdBOQYcMwSxZVDZD86uxaFkBYWsO4449rLYfjH7y1Pf
KBF/gi6LsTHt6rhGxelp66v9N12R6yd7vy9eifJ+fdOGQu/ErC2AMLeZLCzuXTej
9/oJ4oBxoHTz/brw/fPkv9mJde7QuFmCZxcPi498IYHEQyhcYpNUE/IZr3DLYKpP
ZNZVYMlowVGE5uUlUkye2DwAo9re84qSKr1RHGV+PszB8IFW/YMACVrlfn1GShF9
ROudeMPoH1wzXFD0kETmLcUH/vErwYyy0qy2ESMTYztYWyrx71DgYSbUCLB9zQc8
5uScR11qHZMdxQcyRV5Sfcq5TER9f1VFYORvspWuupbGGfWmqAV56WK5ZDe7/l7+
Mg1ax5d71ItyIbsRtlfEsZD6272QbLTVREp+J3t5ezQAs4IwDp7qlZpdiVZwTCB7
NCipE3PU4SnCy6LQIw/fFSTNazrjhu9id81gYY9c2rjEJPcLVZDKznlv+PAAXBmm
ib+8UnB6XgEYkoCHUxcT6y30WV7tdUmLxMkn5pedWA4QWEFEtwDK9KednQLmfAd2
XmMqPJFThQKYroHN4RG/AIrVVmWmgCPs5gG3aN8yxNtYRHPVe3Cmtld6uyVjTx5M
K/rkP9Hlu4P/wPXj1OoAIgX3NaYuL6r6htiw43RupsibHTVzG7pAlebVxHP3QGHl
XR5ZdmtjAsFEXtYPDPGdT/ScBI+FYGS66OxylbqoOhUAzqt+PnC6L7f/N54o1DYC
hX/nehPzHPAhFs9Gk8y0NjsotIM1cBIm4XWNOX8WZBKJqmbtZQbfXEixLp+exMpO
KEa6NZSAFZEAheb8+VMp3ze72PMwWPWt9cMNvOd6ph0rhiVV/myZrTOO6nl8bibK
3mOBZ8w8uuNhAPyIWlOCcQCfaskcNtaFDT35d+i6L5wiEuOb9TS1VkhHaajQW3vF
vHHC2oRFLUEjDYWM6XvCSk1v3qX6I/hOT9Ia3H1/g4Gl87Ur/O3MefWpTL235Qv9
y9MlR62IxS8SLzLRsqaTYF6DfuZjaeqekvkFYBUQFC+LUYehI3YmmFQ8AePOxfS5
rz2cWa5AZWm6E8IDtPSQWKPRjCltRMh20yOsqeW+BEF/ljTVTnak2fSiUn4SRVct
2bBeI4sjt5dUdot3xtDmHl7mSKqUNcri8Q7CdY9POBmKwTbZCYKHHZ+1OYFKaXKM
s6zwuhlARD2jsbKTTeOkfiRzpcDHK9dNtfIJ5fb39Sp6CrHfYnqhyoJhuxJDRHzl
iWxY3xpuHIF9QsRncpNRA10O60t8Eaf6zxOK7nmOpdzzQqKIsjSYd+B+higc+a4D
R0fOJb7p/q1OQNy092/9D/Km8PHnKYUwggN9qtdUe72ToGnhUSF7qWs3FrVR8LYO
q2uEb7hChP1d3YAh4wmU28igh4VofuPqakCOHGneIHykCZ4pHa23hVPtZFvtnCxh
0vLSApMVdz7+Im+3u41WUAQWYzyaEsBsRzu59od++JtoKAycuDVq04/5APciSwX9
j/vbbRMklEAuZ3Kx8hyJD7apETplHTqfGRKzyEKxV4X5po53tX0b0nvaz5m49WtK
dPS7BFt0xs77RdG1NNfpmQU9On4FBCaog8s60KNMNnqj9bJADFc+WOhvdR1AMA18
Zsw5gflkNatTOkMIvdU++HBCn5ZgOFB65TayS+UrE81BdVUQvBKNr1CPG7EC3oXf
LCyWd1vi02YtOxzxpOqCbchOsG0reDnTvM2xPia/X3nB339CtHMuDBCzkrTEd9bD
QG0hecl4Tyu1+nMZeV4Ns1Y/IFqH2PMkrBi5/U6jDwltgoYNI8tY/3HSOmT1v/vg
5/Z5B0o3eOscooNl76RjolxIaOlo0d+Q56paTtqEnlopThSoopuEy/kjbBcrWtkW
JklG1W5IR2i3Fy0vEI9aVpWBq604fkpUaWJYJG1r8k52iGQvGB9RS4VifkFkbz6n
XOS63Glkjh1aiuT4UeTxy0OaF/eUwbma3357gs3fiDaOp0FMZD6TU+Ghih6pRYm4
JqNHa9H6zjw9RjL5p++3cO6A3jybxg5fDkfWIYfEQLF0vTJMYEhVQ70EAmLaM/RG
8HRqeRZWOZc/SwhscA2ucW7LslZ9rsl4A4irN7tfKKLw+q7pUQh/KHlslAXGtglF
6KmqtUSQuDO7SMpYSyDIvlX4MOcU8fWS2Jivu1itzr2B1pY06TJLmSY3nj7Ifx7/
gQxtMorJ85Pf8J/VVi2a/Q0cWHHZ7owdZNz+JTfxp6iCZz7droYYvZb84KavVWx2
mnRiMqmHeKmAmpUjmrydbk87eHeOyU7xD1t0APcjLp30pGgoCdLPsj3XEk+O3M9o
/CExYpPY3MOGPfyDe/UDLYQQwMvqFpbJQMbayeYSB0d5TARzbyFL9smDmQdQPcd7
lZciDCGQxYINYda7hZfyIGqC3N7JQdD+qnYLL6nIJAS44TRGiiQ67ulUwuWMmJLK
wGKtP6P5Y/+p62ysnyMBYv4JJu9ESZ1JvsRKDUwp6Yo13JUvIWBSw8M+H4ttVZmG
7xMhM//ake43r64dh6jKTSwX7AxC0nw1n5n1qZR32Tz6TYzguboUxfRD9vlcn9GK
cM1X9r5aXustVRomBw7N9Pj9HZIKCPskdBXXRAhE4G9ce5RaldiLAcUA9QI/HwHp
tKAEMewaVskRQM/66d1X245Eu2mWO6KhbNR8210Cb+tOUYT2PWRWQRHpUTDkpWiv
+J6j31Y7ivIHD1MJd0dW3JXXzd1q5tvSTfzQ7dBa+Qn/IJyiIXRRQKtWI6cZFJkI
80rZDyHZrbPm9IGXeGtnRfLuyhkuh0pfTcqC5Yu96ZhbWlm0utI8havKAulyXqlL
3h6CyDKX5s0R3A0ECzTXeIR6Apq2YcUGt7rHw+edbpvbWRUZwH4vxPz6s6RNMgjI
06ocwLv2umYlUqfyiV2BY/Nmxw3bsAvG/Y8M+zDiIsv6a/NsxUhgZXcKewGiRE5e
tQN/3ZOyHpStceQIk8mzxp8u9xt3FuYWn/+9c6rDmeB3eygQG3MSA2N5xVnaFGML
CDGW7C2GDcGKjJiQOiMZtGhoj6uL8LDZtPAm5ttKuFFemPl8MtmArO/lxOz2+Fl/
YURUKqGd9bCrmWBC3lLO180rZuKyfq2dIqWe94+O3Ll79LJlqjsLNWh3062A/cbi
f7HKv8G+8zHZ/S4YPsAgEdzaMVvvnp5mRQQZUAX+TxZ8OlN18vZtYFVla0GhF/pM
ViyfmpTwuf+pR5lrt0u6KTSqgpHsdh14Q1jEaEOKM3FA+uLrwsn6Nchn4MoiwFrT
vqFK1YtUZuTNInXoJRkKBnFW3x0JZT3dALTvsjRhIMjupD7QKsg+J9SNDjPQxAg/
GF9+NZx1f+ICGUb9XjiwC4Zup5vGvBHrrTJoe7j+QjutvblX5OUoI6+5OKdOqcin
ny5r5ENrNpacfsSdsS1ozwmOF+tYfEf24T1fOfJh1jl1tKohfgQ/9SlcueKRFnSt
1bhbO7MSJmBiPSKpBnnr58Tb8K7HHgXWtYE3Sd03bqd6h/Y1flql7f9bJixc25RW
VCO47B9YkmxkNAdZloGbGOoalfOoAsK9H+bPnf+fbXC5E9JWmCo6sdjG82n0SQF+
sDMrzGVdS/8FFc+tETSmUIOInEXZUcwVgG69XMjC9eTKjebcXx3U3wyK002zAxBr
lDGBuGH7tifyQVYAsNXcpbF/s0Mf6k/jx9qOSHMJR6/8dJ3KOpLtzGB9o1qFk9+W
BeflVD2jv66J4EbaxkhvFYHN85+GdmLb3ZnZZi1w5LAJYQYSwLIvvKBqYys2M7fz
osjSFo4m5stQN9LcuVx+lZ3udjbWFJ8wiXxKJUQRYy1XOjWKnFDCIvn4ziKHOl2+
DsowygDwNfomtr+c5RfMV9Ari6fQGQS/iGEmyIX/a7uFIbrlc9hcV1GCwv5cYytB
RSUyGdLlPGIYFOIwUn86ZDqDQJx6G2YID2wFgF4theP97Yeu+w3ydy0usiiKL4PB
vj6JCqgZpI4lNUW2l8AFd1ZJC0FvAYAlzf/Cfa9LN2jGL56h6vbmgq+5ZZPmQpJ9
bGQERBwv3ae1XKXvGzcyjamXnPjQo5Czd4j0sFTwdP8wQLhFpaIr3bxSx9n8+95a
rcG+7lvj6P8la4S/Mjs0p8fyIWbHSy2sYdEDxiUysPPbziUAV4xpBZKIz5EujQZt
LmTU90wuQkO+F6FMmXolN2P1yG2QbUqhlx1sjFMa6iu1xHClLMu++fvuVPW3ZOuH
6PxPYlLeF2q2Ha1albtvTW3mgI19GF1oSc7QpYakfN3QojApeDrgUuSwp9rdmq+8
WQv6JGkR/KbbhSi7/z6rGsf8uM0iDn37HcJXLx6dmjEhMGbg6Meow5DFRWK3uKAW
0dg1Q8+jz82nL5QKfjPTmApW0pp6AUoD9J5FTlPqeaRHIG73+jIfs2z+vBqWFmhn
tZFlTDY9jz5Cp+qYQD21Ih1ilBhqc0r49nbZ8Pu9rFYKXJXYyDyNfFinFxBKM7Gq
qvOIuSV1BoyloDzsRETV6bChkXDzQY8OCa9fIPI1BjlRMEWSH57pucQEarV0bfWF
kcN7DJb9BHubxUriNvvMw7OtAc3fCl8JphPlZBakWAt7MUp679NSb9WD/o7kRP28
sQ/RoHxdg0u3mg4VtCLZTQgn/ZbTR0BUYbiUhLds85EpCM7ww5Z90T2FyXZXGBMq
UYnxe027qbCnf/canYd2wzkJrraUWYE3iDCAFJP/tqLmZkGCMSBLj5pJJyOrU+H+
80Z/H2eRNICuehVbkoLlfUIuvoftkBErrQwODF9k2v1BiCv/YbfqJeiOOKeMMyoq
1IeR7di6z6NdrrwDPkAQxj3VHWGGL1wwEgzv2B8JnpLVdVBpRtl55EV4F2VPEaKA
j0XjxXAjdpMJO4pJCpk0njoid0stA/Gh9kHgaz3djp5fc8rCEnZEEcqO2997jYom
2xA1/6CotKwXij6lpFNOlJBvfss5B+zn+lQCJu6GLOLX8j0ljBTo9XhzNMoZ/lL7
Is3Mjbb3OxcBqM+VASUTdtbTvn9eN2/aCOu9EpX9EY8kVoLJJ4TEz5lXQ70WJzYZ
vXTTRKUsWN3eadUi1jrklFxzavSvblgmYcoEvtE+YWj0l8dnkxKTkn9GKqjGlwXr
zf3hEDDlNyZQ3YNDZDxcyPQ34cgtU4w3IE3Jton3eSEo7wT0oz+a3m9H5An78mDJ
4NQo0dDD5t0cvD31aRia1rNG2ujksHWK4U42ZazZWct3uSANpSN51ExpzCYZuOYd
pkwZAsWp8lBSu6e19k1KYs3Zv27TtJHqaLgD2lQmvvrgL1glAcxPoPJEZ5J/UtE8
c0xfytD2H03yUY8rZyIfMktD+WPG3TGWgAkzWLJcguNgzlJw38dAGYXqWsgcTOvw
mJQ/ODXvaYRQ4Wt4PTjEyRd/0voKqBFVctCQN94VmzT88dHb20/La8hFaHO6Mf2m
tZN45Sq9AKV9uNve2jnMJsCUZVy1Ry9ETVILfwUAWTamFDzVnFqQecmj0I7/4BR7
wl1wIx+R76Me+eaBjhN8JRyR/MYdRv3i2SOYOEtrhK+Dz10xGDqHlMtZrwbiT3b4
z/yB30Siuhzp/+fyqEP91CPgxSzEdHWJ37le88FZKF2f8FkZEmJP/8s6j7svuMcG
5r3Rzgpj/55d50PjWdyZ0owGm66QqjUooX3DwqV7oFNyT2xDzCoe5T2mUmanyzAO
ZwiOAbpFxYaB3SJJ7kYOu6EJ5W0nlT4dLD6yUwtV1NybQjB6YWzYvF3dORXOnuuC
RNShgW/ESuUcNjhgAYFKo4t3SIFhRk+9vR1zOF7Ad7rE1ZuRy2CFhiewi76jmVPi
cuRXyyNXr2fzO9I2SIq3a52qjCI9WkIgb2VJ/39o3AP57vi1lmGeiXFOfF0MMq/M
aNvwyn/dP5OZ+iakyt77t/KJFnULl53Mp13mkJ7a/LbSjeY/M0jTPBf2Vzh43+Pg
A7Y6S7x247SeZ9LSSB97ZZ9IfjNNeh7Ad+UsjcEzsQ1/T3N3VVdBRUbiLh9vQduP
+BRya7YciRRk+UJKyT3ZGJJDxPaXnSIvEO3kth506UanytV9jaa8Mmq7CJWRrBV2
pMjIb977Fq6Fof9fNa7BvJ4jJFdrQxBP+ir8TCTakLkchBcVkRCy5zoiKSgvJf0t
qLqj1v0fkbYVjcDNx94gTzGA8qUpEy6pXWmMtgKGhE+9OA99QbtzI4hdtoZLVI9W
0AeZjPn12SP86eN3wpWdvniyE+NMCq0jOPTRa+eWOigwokmeWS49FhIZCju7aW1y
Ps+lZIgA9oTmhJPRMcGnKPEtBSSU35HEU6PIxgMhIHLvH2bO6LEaeHn58+aQnEOz
Mnf9ptmzCSvYEdmMAK6UucosKv43b58SCEiOxx/7Zj8SbrFnOMajkcuSw1UWFdPs
mZmdmgnMji6bf0vO4oGPCfaxNXf2vKi+w3aTeh1HVhNdoyzrDsX3WCzZj2Q0nNYb
oSoP70ejyIUqjieSyt1L6EndP3lndIFMMmJAfPAbJDFp5DtSav0ZvQRQ1zHbXngs
Ul8AsnTAbEagL7E8504pgL/wdulizVTaaRCBwJlEIwsV0AtQz9gg36PjqKpAj84Z
yzcR7eTxk5X4yen5blmS1Ezj8Bc6XpXFvsw+lZSI3yNyThRXGObNVhbRmI+PiRFT
A0Ig6voI2/dKYdJx926yy3Z7QPVT3YnCUbnrfEYzd5jVgUnifjLb/3Fw/8n9dZU1
Squ/qk52P9qBYGM2lq5grGLHs+TbD4Qom5t1zlivYhQly9KYbq4hSiBCGW8QwRnG
P/EORt3jXQv3zix+zwpWqOaiv+lZUt5SxyvcbUdeGhqi1G4ced5oCbYmZSnDwkek
LqXu6flsC6CJFxEfMrv+E6WyGzR0uQs9CV98lg0l38h3FaoZQKGkHrVGQ1DmBDhW
qu2v0uz/OGKKNdEs2b3N1E1yWLtMZZvCo3GnVkk4hweryYg7Kxw8v5FGblQ6CivQ
Sh/8nBiumG1ghAyJqIGgp1KtC78NgEA1V7+DKydqvVtu3Y3S+egTWcTRgtJQdUTw
pgjJlIVube2p/nwKEAtAR7k0EbGP/k50etEHEp0r1c79onlWcLQrwtVTXmOC0zVm
cIWW0nsOmZlUNEkeZ3MrSmFP46M1RjKJ+0xgMXvUztKiPfaFuxz/VbeVbj6JjVgf
Vn8A7G4FZVqEECORew8/bRBE5pbAN+3R8Nlx6avvjGmzXda43KbHK9ZB7tc+jzUh
4iX1j6gpERPlXBZ5SXCAic6MjnRplwz3JYuS/q5JEMrmZsqzKDF53GpGlh/v/pyo
pioWoIldSfOnNU8qFE7Ha8YBKtLVOcoqlG4Omnk6hrfGhyNXj7boCwv7eAkfI0sf
vtvM40aaIpjRddDzRYK3DnC9c3U7loCwSzbM2MLW8yUihr7H6GDA/7qqJXyV7Frw
C5PL85QzBUTdittvVNYCuf1kNWdO+aBXVWylFQjl09BnK5kJxknCEl0w1lH78FRz
DTSU9cLJQ9qr8segCzlah4lTxg/FkPHICc5taPijeptgUC2nxF+BqElpANHHMP04
oxNjpW1u+eA+1xLAsvZ78R1T2tkK2SRCsAI6+sWZohePyjx5P1Zq5KvgU7wITNfM
jPO0tzN1D6WqmFYTtVw/ZYffJhEria5RmeLzLEf3BDgOc6TzZx3ZDDgv55rUWkVn
8IOcjsNTKEJE6XUiq5ViWV5tDLGAzilQB7g5R2ZMmfwEe7cK12VsNjCT5SQOuYVc
1ANFUgzuRnuBqgb3iTmO4Pu/0MT/u1ZemioINxJxKh//R+b/LvHV4JfwZeM7s1md
6pR3KN9+OK/MiklDLlDbTAcbmT5rcruahB4cQLGaKXEzWh45Tyo5rJP8YiJWrnai
eS/FPV8iEuABa3LhQBDl/0xA1U10M/MuKL4tt3sqxYXTS2OUB4qTpmj2qaZkUeD0
68LY3ku97A1/T/Jf89w+/pHTqlzvq/WHdMtJsGwJg4VOCirdn1/Tt79TWoLE9yTC
L+vNgz9YTw6HuT0hrI6+RZ4gSfAyIRR/vWl7A3H/Murksln5PPo3IiRmsTO+kAbu
5bHG3RTbtJC7NNXY2wOG8FrQU0Pe+XieikYP7F1hYNTO4rs2ZoNjnM2XeZRv5RFB
ypTXIv2O3m5E1UtpuYDf+JrsJbWedZR9rjX0D5wfDQO2uc7/eYLxPCrPU2rYie9e
wX1UA0A2KLa28hdWI+lH4Ba8qGgaScvhYYo6lRr+4kq04+R0SqwAYLSrgp/v/xxH
j7JVULaF0bXVbLF4VzowEjYkgZrBxv41Rxjgi6cU2WbcLK6dxdEeSZvSStS7maX7
QY17FhZ7LleLMpc/WIcOV6AKBi7L9WXag8o6VKh6AnRcVthvVCDkEz0DSaPnPk1z
ZbgAvJzc+vRgctjdhoaxyWuRQwK471JenFrhXYQU1E74wVOpMhWhLKo2Tb0kJhHO
Ln0Sw+16My6/Uaga7CURXq6PJQq6UUsFVxyqx9rZ5vup0wwPafZMdB2ZAthgRdlF
iMk0lxSOdiz5bwFRQwrp5G6rklkPt512hc7xi6tHtQ33VTpII7B8t7+17lvZ3K0T
8+eSHM1vckdQmnG4KxmLN9x1MTENHgcB/ttgtsA+xZbmHZGm4NEfMo7rtnrhpKip
ktEytYgECqRXxsCSmeyo3s/Yb+7iHwfQFVsP5EyUNSpmH66d6aVNv28TxAquv8wG
Yk2NaJIXpzZqBs/o7XY1EPguvNJQtuBQqx/7xC23s3YcBBnAFoxVexiSmxqKzCm4
uZmxf30MGHddfxTuenn+1aq9NPPbVGdqQeO88utRCzuMab0+vQuIjU8ghqEZpEoE
HV5UJ/pk5vmensr95TNsku8Tjjgg2/9iYuqwiznJtHN3yG/GEMVdfYYON8FH8hqh
FAaWQVLgpe7MsKXdu6MH2mRNB5pRuBFfac5ukkMv9PhqPQb95AYFErgj3o8X7Zo1
BReh4L+Rax2BKR9UqQPFMDdzDuXG5RY87HK3UJKdhauIm6vyeRo1Co8trJlkAdHQ
BdFL0LJMjMqnA5CbZhTzyw6E2VWx/fhvLVRR7rTmcPKtjcgY/j9CbnxHhIEDojDN
UOGrCnPKdBvRZJ/d9pDHuWF2k7nCQb9e1AxPVfF4RzyC5HBz5b0SaXYfRNXooJm0
uv5vDi9IyzD86ABV3eF8W9LmAIpH2ccWTK2tSAoSukgiLr0PkAy2yNfjblmlCeK+
pyzTo0ChlemxDsg0f63FlvNQgWfEMYERvoRQBEPS3mUOtoOLFlzSS1+o3cAVw3uv
j0JAROsPIa2WoOlkUWalh1zxLbA4Kw3V+08ZTuNUCcTMfoehUrUZI/QpKSvfusCZ
mmmhotNQEZRF+YL5X039Wqj9o4qv39dcN6jGZ1I36W+hFJfFP2/lu/neDYO+Pk1N
uSbaAbOKe8N+F+9Pk03HpYAwlzCUV2DeIaPyz28cDNfwLvJOjVmaPJ4aOrJ1SxyZ
HkcJ7KvqVrm8KTAXMUk6ukMdtnT211LBI5Jstid5GqkYflUuT7m0pWCgTH9vFhzd
FFJaOR9twXoKfBkf5P2mRKL4xGMe5VZvcmpJ48x8rlzp2O1mwIXNu8RCku5kd+gl
IIi9t5/RE1QJNRA0QnbfpJm2/Jclzv+58cWsZ/i0VCUMKeUCy/nprIC9hjIRKJly
HEV1QU+PugigfQkAqpxUpOdgdJ+XmuTlrEyCb6o965PgoHcDf5aEZMgt15YoGv3v
1+sViiVA4/fxFS81ZEc7oCYR8mhfKtVtAFpAS4ziL5rY5sbPp79TEpTSBfijtoKc
4ARTbxQOEj8ImxtRU7rezVnRUF6R5toPec5oTloeVKpndO8U54YgThZjZW2a4OVW
K9UT6/uNNN9a8A/gxKdvkQ9yA1UDYP+o4MAFRpRjM7D9jscKDMNdHS3yJDkw/srn
RTHwkARt0tH/1NtFbGEGNVrvPfn6DsVjiKbpUnEbyFqstJIR86evq1HYJFHAoxa9
MRgnZ5x7NgKXzpQhWmUbjXs/ce5J0ertMA2HaHdklmLqWf41abyn6iN7PMUl5Zyf
ilXEuOdG+gifbQjdLDAf1o0buxBrV0eiep1OkcvdBeWZS4Zt0HWidpJ0fWKE/7/R
NUT+ZcdaHYiH/XwXmFLW3aSAcv5p6fqNWeaIhIs6XK6husMBqueBVEjNresHhKZo
UgTHQ6xYozk5kqUhKNkCiwruB9YZro2LtRZ3SsmuEva7E6eoKAzTVqOCKRsa7NKv
afNO9XCLAdTZkwoKEilLsq/oXX0WQ17U6njBODlVz4BC2DMyB5/AE4AyQaM0AXMw
0sawzQZSebPHot5Jry2hPIHDEI/XAQdFpWKNoBrbviug8tflrM+3ogKCa+9pueZV
FdNoHpIEo6d7XeDBXfCvIORTipCS2Oa0KmLdD7zLxDYKuRTFsFmvXK7fRhxPWFNf
pX1cmrehDHn3Gvmyc1Ur9x0A7uQE4QpBzOrP4yYxhuUclMY+G6QKShfXg/vfZPXr
i7C2sHdybLNcMi2BHXa7TO13t2OdLp856c4oGyefdaNEUVh0GVXzSq2mPcGaAon8
+Y26KI3YVaQrn1AJuNi8W1oiAwmDUeeLthX8D60+s46inJkXyYaTaaj+oX4G639u
0zRSuQ04OCwuQ1bgHjrfajy7bU6B54fiAUIXRhgLZJMrd63TLOdP8CkX0s+JWKsw
fso0LG0fV04HkdliFryDCAwiGvqG3Gl7aLu9kZ8m1fXKmGEjfy3HUrpN2DmlQWul
/M4jvqki1J/Aiw5h+zODnSdf6RerQC+wwYArKO8H/gFffvwWLlzUk9hCu/MV/f43
Em0cwgG1QLsYOCsIAdJIIXcuJ3WI+5CRfgmzP1g0s8rBsXFdJFm1sz1c2tLKS0SD
CJ1YWrh+DpIUOWrJCqzg1gJDg3pqBf/H/IQcADLiGb5CoxvJX8l5Lt6DedVnTEqa
Y+wEaM67szuMDja4O/MbsUwSdAqUcXMq2c8HOajuFYXmX4ekkASKeioN453lRKV4
CdT/Wu4v7vihdQp6g0YIiTc6umgVF/GMow7bcznt5Sc8I4yNsawrDNUgYBU6y+tC
lP5LkaSsFh29SF8SUJM1NErXbj9w8es6pr3PA0JwK572EG+HVWMuKND80bUos9ho
zNWK9fKpiKW8tBxhiiQ3OEmSdbeAb2XEcWTSeEZPtYcvo+jmKIQ1iXzIBQ/1GKqO
1/nPI88g7z7VAX0mRSpAZR7vzXGDQw3wVJE0Ioo/T/F057+Ov2LI6bCRnejfPwt1
DXYis7a3gqKtfcdArCXNx9sEZ3VAZp1quHLRQGAXDg81dFTSS2ldKWoTNC8eUFRI
8NAjvd1YSkxYSql6onHAgE8O8AOlVfY+MHIX5dr0fBRdS6DnC1Opfz4YWlFqF1kl
UM3NxaU7/ko4neSArjKjE94UihHzEK6jDSrC85igbQ/PasrRyvnrFNM+DuQh6hVo
oBf7PDoZ5WVUp0zwGbNYuMUpBPCLKzOSRd11ZqXx1QNB86sgjylOSwC45jxrXt2J
LUf61riaHTymokKdlHJUi0HJSHeL+FpwPythUqVkVnSXNvFrZHQAU1XcREyDVs2a
HRnaHnPJZJxnOlAv9e3Xbs/lRATtPJigg9NY1PFASP8prchcDGLOckNmjsSJ7tcx
nDslfA3Apjdf0utGx79ppI2uD+X0TDTrNI4/NW5eumrQdnaug55MP4+6DVsR2Kk/
S4r1Tfs8cR4W7Mpiu/lGUhxgJFOtsEKy5iSEyOBxOyuv80V19nVFBxI0JExzft6O
20K1VzMpLX5q68A/jEEA9g4u/xrlGaBnFoTZqOTkqUFZ2m731uzgGHOF9G7ud+oq
YJNhggUMeZ8uNLRisQlYGmfmA8rYHsT9tqlp97wmnSt80R2KyxrjylS3UnoyxrrV
tAIAdR3AQcIJvqTk46foBXJcngx48BMXiCbu+WFzccE6ge7WG0ML4dP+G3lqbZO9
Rh2wsio4hOF9i5fUGjEPk2s7VxVozjMDMegzUEyqO6TrEkh3t0vnHxKCiwbhF/Ca
bmqPqiRvL2HOVVftZTGPeD42C3TCRBDtMK+bdlErV8zReS+EtJawNcL7OvtNbneP
tFIPS67tO5nntrT8ObtuxOmIf5av5n6Pbjia1l8slzcRctLCyrAHHVICsAiKy6JW
yypXOQXw7PPIj/3U8vX0/QOJgUXEIyKMK4XMU1O+quZdGp1j6ftpDisY5kZM6A7O
79J/xsP7MlSZgSIFYiFqGZCq9JT38jYx9Zgpqi8DJtk8amNeWXFn6POFTHjImaNj
rka+S6bMJFQdc56VPLi5BDXqy2joHQgaH8ItpKDn5WRznFuVZubZRTw3n9x930tf
yaA6Ob/+wX4UMQau4NWomQlcjqQa2aW+6C0FKoULfkse01j2i3dlMxSwBlTYR7lL
Mq6PpgNzDmVdyctWjgQw/EYLPkKCt90sK3sI15QyNz/DNMamlHpvCMhpiq89ja3V
w9d0l7fXCzXU1N+JwDxCECVxR0/Ab5VkKH4o7HOChya0tPTLdNt464Mm1p8J/0qp
xLWNsVG3Unr+ZU9OsFOFc8SGut3vVODWjkJ6ckersNvqWgCmeLBl6BY2/Wof7HDW
WdRhNs4cTHjLU4xlyksc2W26jR4gFSl/n5XBCLvtegd+cpJi4mqKM8j5uWDUaKPp
iOK9F2FAMnSrKI7GJ+oKtHXzP3uXeVkarfrRKEHFMvB625Axmppts8fei4zvC4tg
6D9sqm9QRbT4T7X7dvs6DaH6hKlPPSYinr1w2wRbWRB5VnquwWklZrcUo43d1JWn
/WuW/cfAEDSQyF4hsrxgkEEB4LfYV6NpNPccq7OWy2lO2AKeHQPQ3jvJoB2692Iy
eEdXXlrBl50i3tNS3K8LCwXAEEPKLNcX5yX7uE8VsLeSN9xpXvzWdpY8gZ+gxN+A
vNvorxbQ3KOP2J1J0rJs8h9BguzBJbVywHcwaNgnZAw4wiyNPPn4admMtcnNsF2d
3c/neyOYoZbx8++uFagCHlXMxJwrX7T+UDeBemcmUabEthiGAAA7W7vAwiKEmjwZ
GJiKfnk167Qh18DRn8NC7wvt0G4X+9cb7MgkSvD1LLv458nsKD6wOusyf+5n/uya
qtKXKldFgv1D2YULTTu5OXTvNKb/q3EKy1dLSVqTbbje+Rd5Ef6XMfSjW8KgoCwY
0Uu2uU7tf5pMt+vY0rVzz/YSG1fIGdLAPaZ2jlQRRwBrmeQj3pPm3g7EaZ4B39FJ
dYHGQkK4WxXi2N1qRpf3MqP/UHPRSAV6QnbJhO3hIRI7WQ2UkFN94U+zsL4P9/Yv
aoRGAxOok/uDhHvFya2N2BAFKEFVCU8c0Csa9Q2bG4in2ZO//H7vETDMNxktE0zb
60MZ879qd//XeCiYp5QbeWct5Ah+sTkWtHXPT271E6+BUtfBqC0qB6LKIMgvm6o4
t9GDdjP2kjfg8NUK7zKJPjmwRUoWmRG2gzlhZ7hx440S5uGLuIep+vhG7QBOYZC5
r6cFvFAEJM94rz2szVvKwXunlJrLnrB7NRUI6JCtCMf5CVG2cc+LSbPcsFO4JlP5
mMDA6dJQYz4Q9QHPfhnt5LncRYKFip/XVSgISv59AQ9jFIb0AbSZcy/qT4jwU+Ch
LIYM7gpVzaqIko86nf2myHTzudUC+FgEjWu36LiiawkgZ2aqfHWgV/B4KcoBBbn7
Qd7xkWX4ePD3sBnWCYUdeU+x+sGPTFjQYhPXI6P0craitJQ9IzJ+UHwCy0/3i0a9
nBxtuGl0fZdhH3vjoBkEMinG4glrPJRaQoV04H9J4KsrIXfyxUQa1HpcMhar7lWG
aitNbzR5De8UZ7P7yk/d1kTZW7medxd5WFMotboiPudLzrO2YR46YGJeU1MK3XkT
RD8qDJukpzn0BpgQ+grVc39qR+/UNC/6Q1a90fGx1aXEpOZ+JEtCYGC29P/701Q2
4Hrks9Z3/jlbaLmmph1jxej8ZNUkaUWl/CO34TYDBw+edmX3X5K02Nvp/62PiBa5
Bq87NpQkQA/eAyjo71L8AEVJgn6xtZMFfg3fMmjzPavvV6EyMNZLZbLbwbcKbHW6
0XPGeaOiTkEWNvA1sDERua9RZfBSalkWYIDbklUC43FN0dIO+BV2VDHUbrscPbhS
q5EslY3YymT10nkDtEDI7/v+oLelIcjWYW9u4Juuqn4PxWizkabx1C2Y46lxXGcJ
7F/EmOdGpsQ48EPEzQ5I5mzy0qDCSMmBCsyclUbYonLa0vasx3dFJ3z1b03VZvS3
trxyG6IGse9nvpYwWgsbo/h+5wBaShKMLuHFNMN9vG6qJiyWYJs5jUScMnZz+TIw
WE5puTgDTWKdBmtQMxgocIPrhESxNpRwAJ2SxyGBCgOgJWJ1w9n5v511F4U/a/dS
sq544Ov7I6pPlUsOVK9ESU4urVRZuPpB28+m10m6TB132cQ75ABSb15Cv8m4WYek
GkcvWSUPz0IZyPkQuv6smYYwrVspwkRhOzzQBnfPgFjFtLVgOf6OE/sTEb/g9aTz
5nZLRTpS0IrodnRsiGxOBXP5DdT8ogINwoDBnnTfUijVhQmj6ZvK+g05EEZj5DNJ
oqkKAOYm3pZOlEx72hpCoKvDUn3R/Xyrf8JWEP072fHhqdPf4WWHBMcuDRx3bXwv
u9DoU5F7RrOQrj30qJD/NKut+sAFBaE5vwK5RcC3EkTIsXOyqBbCV7ZlQTqOhplJ
e/YG+tjCQCEV3s9nhc+tHRbLnyWKofaYcv7sRdO5D+yLBSTc/ZmRu408BFToLv3f
W3MVdQYTc5NiqvSMsWtl7Tf6EVC0wrf3B9AFTmrrFcts0DFJojHbfRk8wOgXebJG
VYU1BByMIgZzdqP/H/fqnlwUua9EgCxXAG51eqiaAVxdMZA7UAB7eqsHQJVuFLSG
pwxTEP/+d0uEPtgdy7Oy4dSS/wbwDBBm+tzV6MVHwajPugQOtN6zN3AMc3GgIEIg
2+641Utmms2g9shJGzLifSOzhErtZedP52N2ahFNq/LPsSq+dGASxT29MYplAQaV
XrJfeDiSmv7/nHKIqnLEMk8AluB2nsxi+E6oJybjFpBKGbd5i4XD4k7x05DIgdgZ
ORwusjqX31imTG6BK/T+m1HpaStuJardpfqvO1uuSdCzhxtCyIqrMuEDdH97TkRg
QyDOmy62KeLTAyAlAfrA1k9JwLZA59v93bqE3hAzN5C6Ydr1iEmfv3SKcAWYWjSk
KGpUuRTWdJAA4U/a4Rynkksz+mqZVdYDVl1H8iuKdyONSSKCchpIncnN7PvpIKnR
Nx1dudIZpoyRFY3VfbPoYzC3W44pbIluugg771t6raDmiHKC/yn7XDgQ7Z6hdxzW
oxP47OtkHGRZbPAQb1Fdbv8C7IJLBkbLPy3zrnHL87qMifNSyJ1f99m7/cv093cv
arezEfMAY/eAGTNum3377LG1R5xcxM/jTmQoxw74TO4rkNIg0r7bmycU4FOkOnuo
GSzT5DsNAX5UQW3CqzMBjgQP012ZpsyAX2zQwqD4CPYljMOwva00X9y5fSxD3HdP
zmqwU/rSPZMxRxf2hCYaYW29FU/v8Uin+4qIpTatSiKS0k6jpCCa8ZfzYwOVs9FB
CiXpxWQqprMsv/7KmXAdNv3yxWDb6VBC47d9XZlw8XydTsg9YcgMpAm6apvtKrSd
7BW3CNWDEINX7XJ7BAJs/TUDlf3a/5SmltjLayu35CCSfYUf/Zhv3T1UChryjBuo
2P1JqCjs6VDZ3PphFTlqe5on8uhHKIJPbR5P6p9WW7jq6rhL9Sby9tPe2x+z0Yk1
6QJyy+pWguGnyg+WywFfSHhL3wCFABdTxTzf90+OZ2TOL9eMHagDlu/9zbCpy+tV
ywZ/P2OKVPhPMbWR5XRvm8B3brENTE1zvQbr6j5dgWGWUKm8Ad3Qs+/8ue+OOxGf
LL1kj0kpZjCsiVvnkA+f2n3n1hnEugALkxH4yo9Ztztd/M5Cs4zmhMigeYhlXMvD
impUdQ6GRpqRzVOWhEXF54a39AfNILXmFgUOj7EKMj9L5vvkDqmA8f5ZLD/ZIf6e
FiM0+/prm8qI1oQZE0M47M9CWqYKM62PcPZYEmEu17RpHbmlS/oaUuffbYT5zsDM
lmls41NTGk2AK4cTDibnke7MIWzZV6czx9ESV7Wazmf++p/TgGLwXoLO/h21KDsK
l5OFOC7SQf4EPRdCk3+ReDxOGECV2jP3RzgsezTbn4xQlgqV4hwwJ9h0LAHuguFn
5a1rjgtpvspTO+5ncM3QDeFEfQ8HghX2XfaqhYBx2WQvkA5EmWPnHX7F4DBX8Iug
nG1g/uH0xsTBDAqz76U899XBqZ26FLKdJdl/w/whnd/pA1b9QXkVMr/YZFJrkov7
5/qx7pDks6xN6gHavaXnNhD6HFp819oVFAeVw15DOspRhbK1Wv0A3GcNb4jpFbNv
iIXA8dP0w8dZN2VsoQPnZ1QiJSC1YTOncor0deNcBM+b3S09k7pf0yrks02EQW8l
FotvH7sTzt8q/TMzhaIc7lt0gB1KsUsT8hjAboNntjvBd2mh/VLO98LcFxFMUer7
BVjLBcq/7n60/57i0If2+Mkz4jZjkADreyeM6aizVlVEKVWG12Lv92qDzhcHXnfN
eiK+Sn7CeYxwLAWXFt/NpOPChrYF1viPhRRMTfJIQKmVagfmT+Z9A+duyxAcphJe
39PDDVAfqknl8hNImcDmZb5hZ6IM7ykAzHN0iTu6YTeHSNuTbmhmABofLHn8StpU
qcN2XKqTlOw2xAtgZTwg1apGj6d47fjHUYpLTYAIQrReGWQSkAwkUL8oQzEtCqoW
OC4rVZkhCbcG1DKtk6suLst8veFWv2OCuKOn8rl6dvxUF0qXqwbhhwHK8z1QfaaT
jPYpkEuoIFJZvOAYqfwe/0poOl0spzfyqsfviQ63AZfkIvJtZxw9aL26c0vXCJKF
Tkf5+k0GCpNGbeHsPjPH7YkwKRcDcitzQi3j/MvKUZ6g8fWuxnZUl6ffR2XGdsFc
ozSDqhDxOeiMClXT/BdXW04XrutwmTAHgt+jVIBUP1TxQWvE+o8ig+/ZO7cytxd5
ff8XcyBV9fCB+aAg8F9OM2yvD8pQIA++iXoi3zh+1XekVfVFFEYfr8TfFeeOFFb9
rMxmLrDoCtUxF4vzr/RmlH9TyxiSa8AH0ePdoqlmF+qMwG0GrDpG7Do7fRIuIe68
ReFF4QMM/w+I1R1oyMNV6nzuRlf4V7fTt5Ug2KEZoRGH2FtAs12XQZLepctf48HF
F9EXGYaq/Yry5Tf3Mdcex+EMZ2O6PzXrF/aO75cgH+vT0LUMGGceO6Wzbq7mYXsG
RmTkZ+p29tJZ5ELH++bTk6yWxMjHWz5YapGlGak3LewWNk5mIoNWKxcA0ugSaeH4
GlVWrl9TKUdClOAz8UwW9LEcc6OHl5Cj37AI4ycjZbZbMBIE7y/VvOe6Cqj034+S
rvmKpEENc5LDNwwa3VuWtknd26216s0Bp6+788XGq7dlAb3y7+aT5AxE093atdXf
GXQ0zJ85PM4msm/XEcUHAXG/DTAX+IaaL9QG+BUjpwk5l/cQuYMgaNAsk+rovyy2
RuEHTK9JkCAAO6f/OYZTIIvZEuCecyyYCpSGT7hUsesmFVXOhkF9e8HJfgVfJOW0
c1XSrk6Ox042CvKshunLRhQCILmx68mi9lgb42QpVgPXGiPZrV533gQKbrkTXFqc
dGIwEIWwK+Q9hfV6adQfsdWhkKPWaK6n0g5Klq+LEW129EeX2e9Kxvi0drDV+ZyU
wTGLKL2C23v3/jLpI9FR/KQubrH2M0DhA3kmsoaNIndJQXEbdHY61PCjn3pL7JXn
3CABLXv0sXn28J/3XnUp1v1Vw/ovKBKSuoFQgMvUMsiuX5WIlx1XRvDl6mwLLZvc
10moF/ZtUFOrpYal7RQ8xhDbcH9yp8nlnRCGhZd7FfriIYz/AqIl44czHtB4ayAi
2yVBO3378bRbmMavWTnbVHD45uRnSffKGGH4+ogxA5Od6nAwo3MXcQaFFQQI6yQT
BPxOiV05J8q0eabawJc0NGpPBLIg6KDDmxLV6Yfxoxpy+T+epdMU1T5T2Q5YU1MQ
KOBVbGwhlzWAE0EzonqBtetv6LVKLFwUtcxQ0kTjeDMqBKoPnPaJP4Fl31+49hI+
+VAoNtfGJFxGkDnVABT1it2TbiuiTZThTAXAvtyuHyc4kd4mwC0abLwEr9CEMt34
JCcEGeJXjeUu7OtQ+0NigL+4qqF0rpFztqe1nn9GF02fe2lrom8qrbjhjV4yc00n
z9nDI0+ALR40S2yH7KLu7fsyRPVxEI4rUBpCb7ZznpjiPNcIlHHpcecLxdqlqJlb
LQ66B21CscnJteJbZwW9kWtwHOGFIEJuh0BervBiihtBBwKNIipr5l4zTCVfG9hW
nqgyccy/hplM9AVs9iXRk6Win8evONNYDQ9Qefuo+3Vb5dXD+CRxSGtkRQkT5DIY
BzD/pxeMbFjFu2iZOymrSL1M/Pi2F3qp3Y9H4cWnViKtyC+XV9amIBmEqEFsVtbS
HJ835TGKmelB6z69wWHaCjMJcnciC/kkCCzU1Z8pI8XlfdKHCDYjYNbwGHVhsLKu
PoqLhBnWL6YZKXCS7HmS0v+OgOVfM67BaahU9J3FejHmMVnEobmWAN7PqK/54yq7
GCp9S2uDyKeG+qBtVpthaXQe1UeurKG0hTpVOxDEYamBKzJEVux0OmReuPjVFSoa
Tk2mSji0gmlEHG6VUMgVenFQbwG4WHav6IdRdnRAoU4+mYwSvC6LQBax1aaFd5Yn
ran1Q/d7F8N9z8hQ0BS7TqrZ1TaxyeVyEttkz5bhs2e+wQcRaQefcG8vn/VQt7TS
Wi8k5oyzy1ljtVbMqTtxEtT8ozzk9LUucLAQUKwVuyXy/00sZ7PO1WJEASZCXzpC
g4zk0EZfhnP99jCKZIzyGIjXejouwmAl8WTMHxzerA6luLF3QtOOpus4XvADqMln
22gZElB9QlZjOsU1nxDfuJ/TG3vVIwnV4NUuEXnnEmrdd2aIlx+2FOnThBEGNKp6
mLibkaHa4jNw8zUHCeShSYJdLf5UxL8MiiqOZz7qFoShLwqVCvYvwk/C1Z4CCJYZ
5ZkhjSnhKdJWpyxnBHU4UPyWuF6A9p7bGKabtjf3swYK8wgmHQ8teAYhF7J4/fOI
cBamxmtSWQz93oPhs9y/d09Er0zjMWNGhb7Xwb/kneyLCpA7WeAMxHBvlgfb8yFM
51+wGSQ9+xuYgH8gtYA2Gq7lY1fllXMqa3dxE507xpfXDhheEiN8kqtEjQ9PWBi6
5115JV2SlRGQPYRwW5oERjATWqrS3caWzzZ4535csQV40Sh16hFmVQrM39gBlcp3
/hL9I3YbJOJ3LpnomlNY01zwEF55YVB4cnIxQTYVd4JCeuTmgDBtKcn9Xf1lN+ug
+9czwYIzd/6XxbpUousVccSkA6qyYxK2fXdcrzPi5Uiqnj7JbNrst4xCUCZtAU+i
L9/PoeKRLI7IP50yU7obCpZJZ2qJP97WKnzCm8T1ZHziQyISr75zveHPPjSxjzck
BcS6pWKtb/0GtGRwR0e10V0UA0Ae/iN20qkPA2o7SUwJ6Okou4+t+Hk9AfW8Uhwh
ftVw32JEWnPAnim7+ZURTevW6FjuVmGKH24N+eVCyxCL4+uP5FyibON6A/0CtLAw
RzgTEgFC4NPMaDMfs9ZrHqey5kiHWxR/dubOQGfxBZhFgnwVfDEdQoec/EOYW4SE
n2bXx7/W9TxWviTSiuxUWvQogEMsYUs/YXZEg0JAE17o4WfIOumt+1bqnt0Ef1tR
P6NqutdPRhSqYPY+Yf1Z1I4a1lS2ZXGavpvrq7XLEI3ZLZkNdf4au7CEYimYMQC1
9i4MXGgckgJRCHqvCNSsTLMHw27cUWt10HtrI44bD18T33vZwh4o4Kjr4Pp8FA0v
TGEtFpBEcLoSrvhdU6ey47clJyOtK70+ZenPhqFB5s7lbviaxuW0whyeJSRQEets
jMDjjr2JyGTbB75sa/En3+pHJ9CLlI/rkE62uLJL+YUKYy1WG+M1DpTGLLKnco/x
vbGt08IVSOPhxh0N1TSAgDKNwTl68unk2XfCv5XXpkPVvnNORMMB8ZBhamttkI40
IF0zCzX30USxO+d1I2Ti0AhKN863GnH6ZCqgnMKtJrrYdeRMwCqzw+bK1BdYEP8g
KrwbdZdqHto6Z8/hqlZzMEFK80Ds+SpDhOnaLXQhM6VZPdO0qDWYTirc5ERSaaul
3wndPduyIUbrxa3jrD+Xi6JWO7CNr48yY1a0d3ZemxzorPtVM5W5HupeLiFjNpoN
ND9djeT087+uNRTuklCy39cg+FWlEhDA5WPNsS+1v3ou2XXJx8ru7UDJHFSfTuZA
qDLV5RFbSMmFuZf1OODVkLcRwrjdIWcJ3FaoEJlAffQHXQc2Ed3GbE2bx4qFbo8x
CRIOgNExgCnFyL7qNg9t1OhaAuAMQMJ2Uw6b+wUY6Mb4mmYuiEv4dC+Y3PB/AumA
ogiMiEFqks6t/YJ9T2gRhqsMXWe4r+iLakmpwDc+nsL/7Qh+iM6H1BVJQssA9XN6
QW2clsdr0qClK19LF5+DAII52TztsemF8VCeXJJDxHZ8XP0v/5DvaWe0l3ZC4K2l
4gjrlqJ6dqYHFvEvSlZSYNBFOEbK0bjIciJfMJEJDthqLG8uC69jOmUMiA/xQapP
fC0SGqEXuxAaiDUe+KorCIoiU+hH/Htguk2MLutNTDjqOyXK21GW3jI10LhQQ9cG
jjLc3rmpYFbsb8610fPKzwQO9d5t5JE908FSML7Y+EfZrG5UULBX+guEXAKD4hqL
x6JAyD4NvfpI0kjgyHpq9HRDvVhGcgEz92jhSw0/aSaWFEuaAaODAxIa3yFWmzk1
2xfIIRekxQIGaaRFKcjmbRZi/dDGjhLbSURIFRax9/aUjUpGdkB+R1CWnU2bNFum
j/hW2V5WrMWWtLlcvAR4s5qTY0ye4/0Mb+K6Xq2XbOmOntC93c+11WFKiAmKy6Ov
B/lDtc0gbnkn0ntjemCu9qXOXup3V+uoTfPeS5iEyoLfSXCGrjtM9gqAMPBhcdUY
u7+1KVl4WhPQRDYXXtNJJ39leRFMDsq51Dp5iFHzHRO5eFUd9qQ+/fUgBmo+c8DG
pjStTMniYqDdk5XrCTany/6nR0SquVVrsFGRtbO0gCXn9l6MkoPCe0MNfEqgCLM1
GAfCsX7PWEd/jgjQ3mKbm+QFsLWJtxe4BIMEEt6/wDz5fAO4cYScN71rC7+xj5mE
CCmKWELQ0w0jSfSWzNx7Vw/Qktaj4X3wuElYQ4ZoYLMLY+BST4MjlSSliVMGGYya
tW+LbpRGrJr6H0PnTSl6eUhPoTScq1ECeQKN1TH0ZFHPlDQDoNhWxt88WomVPdIs
D8E0DVZFUOOJHOgZZPToCLMUhVkCzmUrVulqgivgCKMUrz8WrvzSDFy2vqqTV5vb
rF58PAuNPzIMsC0+QJEevyyzLVWAhFCNfThLEopu+bGuj+aK6GptWuGmOuu1jrYy
ROsfcWmtn6SJsl3loHJzuuZ7TEDqbO3MPtHxnG7Ba8wYIbFZk3CH5V4m4+uhQcPp
G8BrM8Dfyy9jFBT380j9qtkOMh4vUfiyu0Z7f9zTVTOkK1UrdUp6rT4XxEo3F3m8
rZxPYI1y+tiAOEyVZxGKiNH/Ju5tgBCz4uBzfrpwsZhNG7OkKXWKIGqF4ehhnmUM
zAHHokTCxzhRyTLQgql3ruhwj5JztFdpRNRTjOqruTnWerbTuofT44dq7YrS2m05
7/HO3p163VCfwxOUOKYipSJ7EfoGdbMzBnEcn/EE74RAAFHcqZJ95slEpH88oouj
HCGo6xzsGhPqcixg/Chr8z67Ash0ftNVfgYCLxzXBEQ9e1nQ3cEsY5KUh1vacvpa
dPfm4M832jpfDP8djAL8JDoaZ1KsAL4UWizjhtJ0Y1fgupuokuxbVrMlSqdjEM+i
cF5PmqlkY+JQwwxNEmZT6AWP+XenGiIRCItuBGHQIDbRMZkhETAR4hGycgnmB4K3
jSskqnsUBwwaiLEdGmtMBjSfYS2dubMubzZ77OHxdKx+1llFMFP7TfeJsOpAuKHm
uXz03F4pK9fVZfvQo240emLzwuEQNFEzOFwX304ziHh5Faj/zya8I9cTXvDdrt3H
vocj7ufN/JYjFe7nwRvGfDKftTjGc6qISpmh/3AyJfTeYiVhxN/2gfxA8w6tl4WJ
+UwgT7fOLZhO+NiwKdn3tBFUUkWvnz3zlE3NlIum661M76QeHCPUlA5TiDPQZnqs
V921bgJ/kcNPCEDe790wzPO7T+Agjp6HmVazibsmy8wzSL0X/Bl04MscKlbxYx1A
hN8QsNA0F6IYqDd/+Uh+u8dXfl5PoogBzSXTo2fMBDEvNrLOb02PNZQ3G6iIkem7
BwtW/14xR105PQhMrM+iKCyqtV5UsZ9xnYCr3jEAzrkQSuHmidmBmlKMt3dCp7iB
O7VA5wdQmzirYp914xFLii+x/2qNrfXsiE0+VHSDhD3vAxwRn5m/USJ/4Gx0/qW+
dCUG1gxArsqxsfnSKIax0IwcBv1VcSoOvaWP/bdUw65MxOjmKfdLlv/VS/RaUBsS
E7hzcBr9ABByp+OJa54jcEovKB8s9pF22su/RnAn2qtmlDolN+zeXNM56ob8bQLK
FDG9FhsWpP0gZ3+4yP72nN7r0D+7073FYPsWIsKZfwQkCO2b2oILxf8Yp4WG2N3t
WwgAnXxUbvHWFuySm6xdV9STepL5cwlGxvL1+11tq8XTxYPpYPKmVXBALt8fDof1
PnD8fcOIpQ2EElGj5rNbwoRBskGbmN6Riu3p0WlqaoBNATwIKZfYlOLebFojrdlN
RbVb991AybDGsXNuxmWukEh984NHV/t5Z1DDThbsLhpjEDh3UxLulQ38T/ew1kLG
ExyjederoP7ofQ+/DYgDMaFEllpV3u2heRhnIi9fDEOBKQDxGVYZMAK/2hZL1XJe
5f4VEUf/wd0qRXXXhkzHBnsE6/6X+JhFqdvDxroYC8J5FwR2qxNP7kU0n7Gzlle+
uoYI/OLfPv61n4enLURUctbeAReLmh6Hrx9Hh5xIy0fbVdt2pQ2azAZrhiM4VKRt
ZAR66hS2Grysbhj8qulygj8TXwAamlL3nj0Pu518cLOLWsNcOe87mX/8ds4Fr4VZ
G/n/UVHtbUuDxifpWIKojsXBQGLjCm45nYAKspBiSziRuKnpiTvGWK9HNkYivDvt
ou5hwyxqe8WlM8cm1I0PJRFuYn1wh0D+/6Ydg8j4GLEWMO1kIjuWTMAKfm29DXp8
s7Iqg3uE77KTHe/rtgx2zWgQF757BsGrVXmpNQl4Wyr5T862tqOL0J/zYX00Gylt
lx4Q8QikfZiQvoJwJsQyzYhrGbvXuNwx/FBMc07Oz1AtYzBCvdrKRQZpRWs/DHE9
4I1dNaMx5T7K6b6IBJj8kZNRywPoiT5o9DseTVf5hgn4Q7ALLnsC4oJucd1tmatY
DK4q45GSet/GDGxJTQBM/MSaBotai6TR5QekCR8o3HKbRPRAGFvSHcH2yWuHib6B
nVuwy8YA/G4GUh2ylxTWgkrDDsj0Ll0iE3RFroyEqd5IYeCpop5OoqHPghADwBBA
Bfq+qF4g/+B6TO0j5nqnTVfoICAH5Uvvid9cNh5WsNRMPykB8d0OmBqDcWQpQdUh
xjOHXKHsUAfg8Vx48oigLwlPrHBvr8U9b4yuKZ0IT61d0++KCvST6e+I840TfUxU
qELfmsMoBKX6rfWJwjkJKZzF90ZOBb8r2rT6x1MzWa4MyFL239vREWO8x5/LfH90
C6FEBhYqHOiTwbnEQAvxsbwk40SPL2eejw/XeKSGIJiTIh8d7SdVTGlLgimDJiQT
j2JHLCWJv1fyoLlsgldKkW4n29YY4bSb1Yv59unwffG1jLcCi7S4e07oXXSI4rFl
bQBpTGlKUL2NqaNUaFK3Q1TOsB7J8rxTn9Yyp3blZigIz5ZxZPJUQaDTVEnN1P/Z
WEs592xaTbGW7LsLZKLbtPzzPpS0Z3ODMksWRaoTOxsjS4hY1YmEeVam54EtLgQ5
iq5P2/K4gTa2v+tieg49HOMIwEu5SHkPNWlt9qa8k7Zxt/zjODvCKWUZBZ9o1XHr
BLAgg82+9UK73HZG7Vsxt2deH2OHGr5CAXTFVmifpsWgamWiUeumT+piCJ/psIL0
O6GfChifH2oiBOMrzLpSNIDecEM8ljnecqCxhBLPvimRzbbQyRoOYtnL6SEl3/9y
eu2cW6onTBBe6A4o88HlxyE2ljCS014RAfqUMxXKTojfU3HOvmk4+f22J9AGIJTq
Yc+BkrTV+HMXyG3YUuyVIyqMswlf2GEt+kViQP0NyrCbppbAPXRDJF06wHhh9KX6
xiLhgnqJEFw6Z+CU3isqRU6YfS8qBm8XXwLnCCHb84DMBIU6fxI3aP+DmQnWL+3I
jQ7j66GzjixMSzG9FIK2lYvBT3pGCGlweVFYIjJyDCZI+eNqSIF6pjdaORI77IAj
eAs30t0GZi7RhtebQGo30M8d+u00D2QWG0Cfs7cQvqlc6hx6acC183V2LaGxJeTa
aZ8JYCnm2S6nIZnLLxdxPnRrgzj2JNmncFNMVJrO4Afts8qicAmgtHnqZ84z2uQT
2YnK9y5zxpeAFYXjZm3NCYz6zzo+mCTw0RMbVymsc1t4CkPQd2hTHvLVxhZMk6NC
r5pQ2vsxVESbdpYTPfZaSlKKvPzvvA4aeUebCutM7dFikA99rc0n9k/8ckoHkSC9
J77+8lGHn7KZRSzIW+g9Ru6iUZjfbEyUwfejhGpnzS2JP6nWWvjl5zy/kOK8CAJv
RAV7FWmIrrHh9Ty3ScL8ZoR7mycMVMBmK607b9E4e8mzZ8GzYMh3bKb4uhrX1Te2
vFjr6YxeQmlnYDvaPEyDx75/7F/bXAGGRfPYzOJt1hLKYBi22yutC/STn1XMrwwc
QeLlNAijwRWfI+LmpZPBxcPXXw41XwJr6/1pnccWXsPqJBXM2395uTpXtA53tCLO
+bueRoeJEkZ6o4ekRB29IKrFtdYHb9Jb+vlI4aE91ScvX0b1KTncw1jeKix84KSw
7G0ICo40zLvAJZQ69FcP2Z7BmxUlc1ToMfmcpL2359vDekKNXdvYwYdZ5n8udAdo
HCYmSeVamCuMrIYCX8rTgvNVCDftac/dIuk3zQ+++xWm5QBeQGlHUpl53qqdX6Rr
tsoUOC4BtP1ZOvFyXxSj34ftr0IBUQstCf+SbkMoKI3uRnrYPO40ZhAF2ekXVvy2
55H+cXY7a/ZBp8OPXDcBOpM3dzH8A5qzTKVcFkWDI9ngYaRhw9/h6HFuwtWfXrbZ
e6mA7VjL3sj+P0FZeCFEXlyipWu78ine3BoqcG4Wqf9TkO6gAoujHV6A/m9mp6c5
0kvV/XxWVACVHsy1kBi7N88/08qUukU5ExWWDspEbfjvH2xRrprTCncKJDNATWGQ
K4a4fa8LzTs2HhKGIJNRfL7b9XVqzjbCqq673KVKnMPQrWzVAJWVXGe/2mDJYG/l
NGB1jXsnsKQ0kIxSaq9LIBLWLXt2TYJnF9EIbuqHniZgjZrAiBJTCWV/y0Y94kVn
UoaFmgluAjSFnulXSfkmu+lCUNUkkGEVayGRxhsKiY5S5lO+IgPxo3FXqQ/Z+V4W
sInc4vJayfkz2iAuYpDelc0KC+vTBdxOtSh9RTOk8XOzFz1dNOj266kzaVUP44Jq
5K7JMKERFnFWwzXBCll32XdzW8LSo9k2DBpaHn6aQvVj7aqfgPetBmOp7jjA4vKZ
RUj9SXrkRqwrg7nuoN9hDvjjfhPFP/GhjVJj9hsuOvNOP9DJ+YevGSHYfhJYt2g2
5ZFzjDDg1CsOIWtr8YpiNiFKCnT5eBz4dygur9GhE47iJeD6WvaL/bKvAb1ut/kd
u03NRZlwB1xT1VSN79Xutr8oTtcQ5Qc0vK0keGUB/2iAvHw1mzZM/cokGNDZVB4H
pu3gCQ5LqvthnZ5yi5Z/LB5/Ah64/W1Ewt0aEMZoiF2nZdCjaWKPRK25Zbep9wff
Z8vhE8wqhKmOoQONqE1MKwvdvvEJXD2k4wNKx6yEZYCvh3P+HXIjRHRhSU2bUWgl
IY4lN1om6YL/8zPCkA38FnPuzcVNp/F+/XJsYcvtWCJtdZbsJ5SAKfKfsV+hr+a0
pIwbw+7s7FwBAW9nVZ2cbfojMycHqdrSJ/eJedtcOBmHXjpfqn9b+CdV7d+pq/xg
3BQQV0GkHmEKb0upEHMIjvSX9aGJ6ooJytjxC8/Gy23U416oesFfkLndBIkJoF3d
XBm19pZjdVQL+CFEN0Hfh3KvGOC3MKJ8GohNvh5jJrslC4Hz3wnaoxeqDsABsfQt
mMk3i2CoOi49jZhdE94dfHdeHZWKgcvE4McL9oaXiPJlkI7iVWC3WUvl6FTc8jeK
mYEgVUd8q8e23o8AkIoDDEWfQxmbkRy+Cvq9yph4K+j+7aqaTg3pMd9Bee/vuSh3
J0Z74dy+JZiFRPsEQHAXT6BoOUh86uCd25QjAVZW0z9+IlfoVvohyOxuYRZG1nFh
X8ZrcXomE/ec4U72t71mg95RpS/wODl8tfE++OWqNW2jMn2b6Erz5bH/18JCcv4a
sMrOwu6gVi0T3mKV1W/ssTQGmMYcEJhlpOvRWyPersIc8BBVEyrZEIuSRCWXoKuG
x1XL3PbN7SHdkP6T1kda7gxd9CRUZMEzW5QPSmBKil7i235S6YnPYZPUCfeu8dOF
bXBtjKt2vdTH9HFytKs/CtyA9ohvMWwJDhk9WVKarznrfBPP9lQgoY5iTuOuMMOW
alNlQWGg2U/lbkhIO7ASejOFUtJToCy+v2c/n5KmIifTzAlD4DFehyjx/fp/APhE
loEVM8GhS9uaGqOKgj6F43uVXNsEtfvnUcRUg/lOv2Fj2BNCdDexGlrGm5e4rLTN
rylGmUFX09tsAdzcj0lI9VGxMQ7HPP4aW3B8+mlRM98ddFd85fH/u+VWRKA4W8Qx
IboP+xvgiTp9WT/FIinig0hLrTcHNzHr8pi7jFHRfEoIrPQJQ2V79C6kl2D/aIAv
9gs+QaYmOIXVU+zzJ6gzNLTFzZnJWqaTKuYDjksJod7dZEnwLtPMreqGI5rWa6XV
hR3fWqlTejFoj6mo/C9PddNq6jIdambMnNh0slWNcsT0j37Ly+ixE9aIUUUzEmGa
ZegIwnaVlKxUm4Meg7dJCXZXxPryEknk2NJsdIn7oRU0t0iK5mGpIb1QnRs35ZnP
BL6XIA45DxkX5CNVOm401kHKavN0kmi3yYRj/cB6ZzAzIWdcZnmg1Au0UHnV3MpZ
hGBfeii05bQSrwMrkp4rQY5P1t6mb5UDxvYVAr1pWrhNWI+K4cXNcolyvCFkgQ0W
UTtDxhCRIwrI/DUowlPU7i1pGHFYa3AkncVTwug0NHgWwsrGdLLD9lBl6tbOaj0G
z7G9HaUKXu11vXSuQxrGr6dzgzxbbUpXsHMB8CNGx+OohBh2jOaDUFANasvWcomC
FLeekIEWlawaPnQ383D5MUk9bwCEq+VWMVDj0l4KsCIBe0poLqgCo+3hJBxxwfDA
MjUeBB6+EB90PbxoYo2uIYNewPF00bsh+rNCvkcuqFTXsSVreE4DGaNgeaqoj/kH
9jXFyKFUJRjX4rBCwuwkP7bGjbIw2Lu91cyKvSQczypEKtstoNQviWXACcmAQqKq
nwIZ+HLIC7e11Df27pFnWBNiImvRKKCZDnHGWbhlm8Hdt5a9fpJQ/S6hbLcfGpXI
l6WZINUeMwVam1kwkvdkR2CIvBmyXnY60WwDRMDcAD2K9euqLuSXTZPGazV7hYzz
4cPxGpOT1ydf8ZH6TI7HHgf39VJut89TdF8AP/xbq7E3JJWJQCrpVbCvVdHDWqyK
HUWfMciiAo3/YKHln27vhhvFYiGY16hZc1bE+GDv44erbh8mmChGk5mbGjEyUAGE
Q+I7nEFFjo/3gIuLqLDfwLHgKs/1/HE9bdn4blwBTEQB/8FwYHovb6D3YgNrYyRf
OhH7bxp6Wp9L733p24+uJu6xW6LO9inyr9nrqxsKWDvDdZrJiOt7kFu4w+W8w3OG
NCnMvCpoJCsAS3nWhviZrN1t72Yy86XRrnSemTm4Z+q372aIwZmu8QXDqRcGSlh6
tBaDkcZOgvjkHxP5pFWJ2wWfDzDXuB5/Ln7KEF6Mc5/Dtn4dPTrRhLEyyaEgyyz9
4y6SIIYGq6vHjofl6dGBwFzTV929GRwaVaHPvfb/QrkawyjOuAf6eYsgA8zZg4w3
QHdfntBsIOdycVwiIbVkIRfeCNBFoo/ZzcMcirQVdqFLaFShIxyCaFS6ZviGlWq0
HD5qNJFAGGvhGTA7u2vmY1kWpggjGGfsp+ZOTTkTfAEe7I+zlsXOpB1d+jgYqaib
NLb2BjBbOJpVkmQxb8R2HCSk8TC4fB2gqxo9rUC3RK/MHYZ9w6vq2/e/mUJVW4Kx
066SLgk2/e33nRNZz4Bw/9cqzc8P+RhDXXVQBFkmGZszK/u1WwrWlSvck37MtCJp
RavajB5ZPqbjL0wzPxJ5bnw5LduYhS089EKSo5SiXlkP55QJbtjyq1fZf9SKwChg
irAqCn9qTZWgwOeSeU733UAnjWNVSQRZp3j98T3Azo2PO2Ky0/gqHmvFPqNdlrFd
pXjjkQyx4nbdF1orF8yZ1btEZZGr+jQQJ1u/EVgU0ekiry68xfoiTwJmMhxVZgDW
8TumUARNWNUNRuI4QK5bIwubZLkz70IeQR8dFQINpCgA+t0axUUcFrHVbvOFesos
HopGfn20MhlLz8Mlvs5nTgiRP13v3lyTaI31ZNUq2DhGGaA4o9sEpWNhbBrFaKfw
d/Oh0UtzLTpY+Le9A+Z/ImNL95020jSyOMU6Ms14U4rU8mgogJmuSKhzVo0TGDlG
rOqEcnhs7TgKoiUZ9o4IK8tA/F1pq+yqpJFovaGXUk4c+E5BpmzyXZufilCvnbje
Mm46DEx4QAKrWnl/WgCY2d73PiTkPTNL+T3FIFrgYst6yZrlOVHAZatxDF0cANnH
C1LYwrJOcd3+GO1+FScarJuWDXs7Q2UOFbQ/NxIpSYQ3kRfC6WP80W0LAms+8iLY
410k9DH2PJ/zP/cPOrQ1GVVkcn+LEh9S3oiGOkxEA78H5TDWLeVPEhLa94yG5mNk
1Y6ptn25hbOJWJ4fkILCAvA5vlmSEliyWaK1bwW8xMTZ/2MkXTlUWRmrcizCDvey
U6eQaD+3Otz6ZEa7ma24teSxyFIkRaq50ega+uZ4lmlr+qpP/IrDp4PE2UrmZgj2
8XM3KXojN9Ta/KSw/YY4YenLOyXXy6eCT0rv8wb7dezzCmgBS/ENyJcFJkTMoZR0
y+iH4leznTF2+C+xxa46Ik3neyWhGJQSPJFaelLwkZxFn9KHTGYxN2XpcR3hmZCO
q6Q8uYxsugQ9UHFTOZY72KNvC/CpGo+ueYI+QeBQAMs0IFHyU8h9B5wilLZwvPXd
iCs3ue3XzHVWoDc1dSXT//lHv6ur29oIEGTnTlGQpNiZJQHXvHfSh3r0dsS8C1UO
U5fmSJ+xFPx+jF6zeFw0rcIIFQR288inWe4D0fPINoHRXRlWjhbQ9XA6J1l3whOt
frjI70DPoOOLDgSdf5aEs+vYbA6VWjlBY71gXzGA7XeDBq6AhFfCUh7+Qbthboql
LeGeWFkDddGPrM9gA5FtNv8Um0Oc8vYpnaqAg1L8l/0heNq0gE/00Dhpa0k5P27t
ZkzAEYUpTjDBMd4PdxezBRqYFRysz/7ZpAgEPNTDcWYlxFLsM/Z1+N4K9COURlf1
kW2U1zDJs6kL1+oZ8IqmwalXTUp9lsr2roDom6LoYkkrNQRUJHW0UBFkLAfi6nEu
FOiMhYbNE3QjmLKtFsqnT+kdhtwtB/n4qaUYOc4RKCFo/favAhYnDzQC4txd6gYT
Oq6tsrPNz1BMd7FGpx4yhVU6jXP765BGgfmPKcUC0WkJk1ew54Ao/54mTE8dfevO
3W3QILlxEultUesdWba3MQ/BeYybZI8hYP+0Ncg207d5uLnyfh/xlx3Z5UUPCKLj
ka/cLDvcgVyfr30PyqAQHOXVa+rEk6+FjL/5qJkDvfrtpyZtk8mKBR5IacR7zSAV
VpXklWjz4McouFtKRylUJYd8lbXzM5Gp+c0liKNWv62PI9qM/iNPvKZ1fHVQISmX
nEMK8PnQ8VA3bvs/au0ELwWMhk4o9Q9S/hqidi4+MAKE/it96sAEJp899GdVG+Xh
n8YQTS9oo789ZEC1DfZt3r40zMkoUIsFiZ/WWC3g884BTO2jWMHlhm801GwEtiZg
RmPSWMpzbglZMk/yN5eZFUYELNH26hy2OXpu8LuZDeLuaDryvw7nqb2kr5Er+o7T
pClbYEfx5U5e6d5tbFuylhR/oUOLSbSpKJybaH5D9WfVYEQEjDm8MQHRUlOGL4Yb
zcQYW3XeEPkWPgLYJCf0DVM0JxgYXUhvbtZWAjY4FAW7gMEddF1aZbZ5zGUPRT04
52lD9zrzroWlQysIFAtSzyy2ChGadNJKRaepFqIcktoB/upIbNVUWkaG2EabpggA
r7pOZ7l4QnwtcFZZmwtgqs9cR0DIRoISeEQcY3rL5AS4l7i9ylbC+Z/l8A7QT3nx
RK7J0Ub5kNEune7MqMNxvc+XwAmELUcEm6SP2+tUINNubPG1UKtkY2u3Iwrg70Cm
Y2J2XrG0pPzxZFDYLKA9nKGoiJ+YHAyiliYj3BLqTbtV/rIxxLjLb7qYwI/sLKUg
Hwz3nagbw4C9d+IMSUmeTBUrGfsOmlbJWvYKGt4GEAwJLnYmIVeJ6i+N2exn8sF8
Mx00dhs426HWTwCTI/A2satpKLTuWbZBF0e6Gkevm2WomQ0MfEjZ6aG548pSV7UJ
auO2CfGdq64/rEX4oxmyiH3ArYGs8KXOf9ilLKx9P4OUb35GMewref4FAlMCn+fq
KtJ6CxtoR+o5p+vg50Es9F6Q7BheldrdaVpjQi2vu/EjTmGom56pzxIri/pTfpCt
afDGFhaa5t1B289dc53A1TeAu7bax0IJZ8DPjefWiKnFq9hCMD5FHjbS5BfVCrIA
GCPuZeRUqs6+Tq7E+7mTaaJdj6KKvrHAA3rXVQ5fu3Euy/OxGAxY+srVp7wGHide
4Jwfn+Dkq2sXzyPSptWzlz2uls8F8VMHAGk0N7XuWTqcX3zxV2c4agghhWyVdznf
yXWRMVDM9vC9uWTSkVF/D0n+Xp/gw+XwWaZd3JPyhhLeGvkOCwEtErdbIQUPaKf/
CYXLL8sk4Z2NAU8l0cgZFZj0L4rqQKXwx2595lksGgUHuakE0MkCuHZFYfj6ZCsd
3a63mkfX5Py7GzUHWhWB4jV+nXgp4n/dktfu4IaA7yYOGDjy8b/pbLZnNj9GSLIV
ibHNW/EDY2fzqpm+6fC0F0KR6fpBxGg05W83EnycKwNjMYq5H7bDTqGz9J/1mh9G
TqZYkIrPI05c0RATu6iUR/1Wc9EPfPGUgHe6k1fQShafyin/jRukXs8yIV7+/FKd
5yhk7XSC713FlTUJCl5gUh2YNb1MK9ZAJ+MEiycmpIMY1N+RlB1cQEp7O1SiW/Kf
eWAaxkC5BQdMyF2qLCl/LnayzWqmO18FGD1L2sPna/hsoN6Quykhl6GwEfKkhOSf
0uTppaecljsjJQXpTffXpz6vmcoT58W3IWSUIlPaNb2xHcTuk2jh8Ici71t3+1fY
n7UFrDIs2IiaEf1edJeFvK2+dbNt8K+rcc7vzJLCRTOiufpsDFhy/b6v85Ycs8/R
SglMU3kCbaQDmcgpe5H4aPXqC+qHtRSRXSHMxHUTpwpev3XYcTlLQxZZuQWmGFEM
wn1KcSAVsykQYqG2WL67GP1A9K5FUaZIKkc4lT0uVNg5fxbqA7lniCaKTigF0d2l
4wZ1xH86yrAvyGWkzxVOeWby9KXcYjmsHWn62ZQ56/Wqp7w4aRkjjis+j9z9O/l/
Ovlm4u088QVbqeL3mQPY5WfWANVKsGevVJ0FBXlYJp26SXgvTOgaH45sioMU3Mku
gEPB5cgivdHb1dGZShCCkvyCYLHfeol9LsjAXFFq77lOKqkuX5yGYSkiJqbV1ssU
/clsqcpGg3mBrD0Nrc0zX7vpiklGy1BJzTbfe27TuBNdhp2jSX/AKbxvGm9mI7vO
2PpRc/hjWh1Z7q2VJi+3t03KlNubUi+WnDWCu/iuUh9Xr0XmdONjSQve4b8zqbgb
wu+DOawCyhA9NZ0eU6jXBaXK9KSjbWVL4bbEffSVwAyOb67MC+sa4L9GQ8Xhoizh
YjoHsGDRTqUemiLFDM7gDF55kdn70kqf5Ickb0jmNHZ9EV6SjU2pDcTCVToeFBOO
RiHru/WqVAm/exuzKWTCHh3jqhSvGdHB6pLAdniDs4MQQJfY5Qw+f9NCFrTMs6mr
IbAHAK/y5eOns2cgT3dE324MyDkf5nQZiJzy3/J0UHw3PwNKHjtM9QUKJhIpiKMt
6SAf4ndrISJAPCCiudaqqJB6Sa5ALoYuOpZF0sym50oevlMq7FS0wgSp/4H+G8NU
M7g1tQpRVPddwmOHSpQLZqZM841+MAYy1aITP708BYiikZEifd9WAe8lYxrvZRp8
6+mNkS8etFMRIVyPEneJ7dLKYGrt3cxNXtCgtotZQw1UsX4haEOZxLKQBTA9Y63A
1VOjEwNvrGltANcgslqLlkrnWFHH38uTWjYl7MFyMQhjDRkjMcRvBjZNCg/coC+P
zWPJ4vW3Mj02otCBuWVQDar8MZ1wv0GnbFoR5MkDJMhZeYzeuSsFQfHKDSAf5lUZ
49sr5AL2eBFEsp841pBpqhNlZLZmrDKeRf96rfrTEvn6h4Wldr+3TMgVKNi9gBoW
ZeW7NAuUpNHk3nZBy+NB/ySvArKTEwgFRV4rLivM9WGUVd3yK/LeUwcQzMyR+R3Z
SgAAlTMR3mnjkC2x5BsFOWZVEzsaCfvmdnsd/MAYe4cl0b9MvZceb7Oh4r+qQM2p
mwzuXzWoDyrT+YBlaYhv10IFWekHQAnQe1kHWCq4I2HwXXb4dbUKGCoI1QEKfn2z
vs7tnlBB0EYOi5L47xgira8IAa4ufKZkTgQjQRAicUzt3zDDFLJG1CRnUnZsms4m
tgzJuYtATq1QeLnNrcoYizjMQPU3dPj21Kd514zsvxettSlYMbE+SU7Gy5b1nVDb
pyNSXnfROKoBklcWdDPlMhEPFtdJUfusubagZjY3Ke8W4oUie4guHXmNUFg1DaWn
`protect END_PROTECTED
