`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7lxj5JS4Fp5NcTUNp8cnCd+IcHKd6AKUFiF19zPWczV2HKFYNEFwhBRh9E0zZQT
4qZuxZmaqhN/pp+GcgKaldWzdDN4WDLPj/sKQJQUFbuzbf4bD4TfchwkDdjqQmFR
wdgR912Lhbn70CYT9g5i/GGaflQ6WYMbjEjLYBW8zwV+7lWO5G7DpTFgeSPODrL7
kDtHYRh2ozmbRfFIxqTeMA==
`protect END_PROTECTED
