`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryQCCVs43AeOveiJqvkSgNsuafoUwmxgYDNz2Yiw0t5ZggYSLGZ6uXo7PBXMA3jU
7vt96ud+g1rQJd8UOrjJti1UvYpb6Ww/Wv6uM2/2z1wQCOetR/Mo9f0l0iyEhVbz
0iuXXToNKAIED1vG1ElBhv1lXBeQ9x6APdRXBLZ5F6rXqxO0E3D91n1cgoWsOrIQ
4p8zctWnlK3/HOwfoDtDu5omZykzvpvXrs+SFETG2RoqdzZOskIurW7NlUVoRGY7
vemZ4yoz7H9HCsEh+xfxvirEObT/JR4v7Lkkn0bGxHU=
`protect END_PROTECTED
