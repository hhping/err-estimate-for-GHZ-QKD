`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPGrM/aQmyXU6pgilNHVtu7tJvQm0U+EZxpqVZZOPPSSdDxi5z3I9hqT/DkBoHzE
E3dOxUCC+AilZOwWbY4mS3RMtucbkMmTk270woFTTJ+78wwV8XI6J2bbvvRSYFh/
89WtPEN/FdcQQa8DQpzLDjrzqGN8fRh8ocMGwP2pesAtn9IBhL1coe4vyECq7E4j
FXlytbLZyi04mhKabhC0rkcOQ5wowyu9w2xIzLYB1/4qd+OVzpxCakXFh1iAPhKJ
tmvewdIPpuUxh/+WOCQcw6sumXWi0vwaUf2zz8X1lJC0XwTKNAWIwjHUjmTt+jQW
dOD+JYNtpcQO0HZjbtOAokrllntkDc9gkhVZZ/eeU7XXzULOP+ywxcwnPr+KHXf6
Bh9jxEZ6SwZHp5jjR6j7UnyhviNJscKPXRJrR1iWd1TDYE6w777bbb8LG4WPsJiV
SBi1/rRnHEh4PW/dhJtxpiTjDGC2T4QEQ+5rMetRAw6pt0edax2eRNAaxe/ba5ft
ypGw1aqyqDvyWEGcGBswGKYH2PIyZJxq4wOA9CVAW3BhROOrjvAy3byeMdj5I9pz
V4Kb7k962hb7ZmSYfLMwnBZ0nwG5oNcZyU0pSENVcA+7dh820RSG/xVAWLIWqVKh
jhv5vfzQRkAdZLROfhjGtGLNnwfbtXVYGNHZdiskOOw0bp6Hlk9g0/WzaMyFmcSA
ezrCmCGf4JQcBX0jGXABdqaw1RxnwQhRSNXKWbEcfzBvh5vgZkKsJ9wJI7HWsa/L
9UE4SFeB9c96a600wKP0lHUq1vMIm98cUhFbUCZmdjY6XMbiRohG967I+L2FDb7e
symztn1Qxf3bSrTuKpErsFtWwDtJWdpD0PMfEPQYlbjmS+sL+a7N2/czC8Cywlsj
b4fARIdJ6uUjFCs7uAF1oWq+9CJ+kchci4lJEE5VsXpZWMbgQTbq2Khe5itN970n
`protect END_PROTECTED
