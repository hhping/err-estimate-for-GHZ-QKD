`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFDIxH5rYC6F0MvzfcqR19LX9WtUHi+YnqDpWzOYpP0FbD5y4SMyu8VadairgTI3
Hox0Fz9zMkU68mPS7IJTHcLE5+OosdjwpGWQOIk6qOQi+14bgUFFzONz6CWTV0H5
yUQ/L+ywyaz9z55MtmVikiguUeE5oNzgKdbiIJaurLca8vDUIe+xIscscPeZK2Su
4p9rPGsiwV0gP4UZo/kjtJsKfJwe0MH8jSVhiOg0JLwi8Ri2+L1UcoYYTac2hVIP
r3nCMDZugDKy9RitgKlqXM5lutqiYGN5JYkcYcoOF+OYW4pVdcA15XlA8eWHBLKt
EeIy8gQiIKTrl2Id2dzV4zQLv96aaqzxQOrNwDrE8GOrR2qPxTyC+fp/EBoVXs1W
DYD6C6LFp8R0NeAKaUay8iFXUudxB7pB0GsknuzQfek+VWW5SVrKHMLcsIMcDxs2
waIH8KIcoajD0gl9f2RdQV1Z67Mb7tgz4QfchrW2atKBdBfc8M97Cx2dS6LsS6nf
nFhC2bCXMOMli670hxmjUpM1E6mmsHv301mz1voICfjIlrpgsULWkzdHVryja7qU
K6ZwdU/bWoxKpGQJvT4ecad4vgQfaBAxYsgSfGogSsybWMWFJzVpYDjYyAC2KT1D
jUu9acvfNsPOG2MxzGkj/R/wv2x+fUShAMXRoxVMdmO+FQ6fAQ30lhYyE781gR/s
AQmAJ1HCxqRk8TUQt2OzcXOTD35jTL8Pe6zIDFYNrb8NvRpYLEOjfuAz+wKGsnZj
kjPHF7vbaF2MDDVq9BVbb8HUa7Bq3f1GGviCqrB0muSKISgwOlzl13sJnZr6Yf4z
pQmNLxtU9vsSe4lK4onITA39lmEieKjFn9VqnQORMVDqpTYv2l/CvTIz3jwOLqh9
N7IDFH8EAliFvr5vosaImxbi6Fa6eIXgUu2LaPz3/GhNd8AK1ta59H4Ggl7dH16y
JXQdDKd0iTtA39ZV34j0UFL9WbnEHVmzKs5hiMwthP1kJuO9KMROjUPlwvZK/RbC
+mZjKdD5QX+DqwYjZUBFCFhwy4E8GkDDT9TuI7+8Vc0=
`protect END_PROTECTED
