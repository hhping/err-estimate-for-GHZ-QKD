`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2auBZsfjeqnuA8r3zNPsFIdAsfBuEvVrTSU3kMFuNfgQgVId1wXnGdFRV1GsrxV5
7RcgORRcnyca/2luCWwWV+fO8ozZwd0quRP5iGw4K4l+ys/v0iKYBZVGVmbZvcov
69tD4XznMDaGk/8ZDpUMZ2wcwOHyep9iIdpcOuKoXzl6SLxy85KhzIz2PVKOsWtF
QXxvRyfa7pNNCL6UKzaQHo+fSHfjM+wDaAx9bykV793eWNfUy7XjYSXvQqCfPDkl
2QoPUW2IDQATP1VJAdFYwSSly9hYyDxSYKAk020mgffVEpaYtfKe61eh/IqNn6ci
Wzq++2yuaao+ZvgnevdvFkVWI+se8g2yXK14FJPxlluqn/xq2vf/COrD8IoXXRuF
dZnPOduobETYzLpbVWmfnaKtH+1hBGoMAh4mRgW8q7hn8n6ccjDUlFufXiJ4ESDS
gu+vTg+mswBljLuzSomcmnhQYbD+X8dyZN8nlnWElTG3nhGbFXmSMWhYZhdESxO8
OAQp2DubC3Ot6RZgjkiTK54hIcf9tdLrw5zY+13SA/ld82buzrVKpO6gH7wGwM0I
TL4dtdD1v0POxNFL/C+UbknT41EoytioRSTJKgy3Qj/ret8Psl2hzeIPPN0a9J/V
4N1hr8eOQ6cOR1vFZVF4DK6ZBGK2LHlRZsX7m9RWypBrjnNWejJ+RAHMlD8ZIQBE
tJKC2/vsI4lW/kZWC11s6Anblhr0ziQCKGwf/HHFFaPyyTu2B6J5ncs45+PbVu95
KWWue7I2kLHFpYxS8FIHXlUGZ1NGSjgXsXnnWybLn2soyV3UEgxXvHc+fZEUK8VH
JWox5WtgoN4V73Rtta45GGHxgLCLtQEb79kFR7Ktt/kbfSAjRTqxv01rFEw5DLcG
TQZTUTzQJhuPtQcY4Zvx1qwMnn/A3zNsfP2rpIJ7aLn1OWprph8omjBmuMWHBzdX
9e23GE1LfOYF0aFNbNuFTnOsxwk2ruDyb9uItIqHW+a3LEakqwkatWoVTeq4Nq/P
KaG6hx4yujyxLqkhxrpXknJ1C+h3BshNkEuJWaqjb60vHJ0OXZ4IPL3jDfGczSr0
FPt6/2eJ/SREp1I7YH0RUTOMtwErVsRlVVYBbA8nfsFakFFzhXe4kxxdbaxKQ0xM
Yam7Ge13FEQhNwGAKg8BqeZkzzpOXADPlTxzT0Ncr8TeQzch+PqHURN/vlOmvUxg
Sg9rSrEJHtUt+867m2+ZFqePDCvHQdzysDRFykmdqladroOW7K3jlJJdFh9hr0vR
dDsGrokIeZ8gd1IK4VPYEhl/EENUOlHA+e6RwsFhUTe9COHkDG5BrCP+DXg2HAkf
ZDdr+/r74BWAgNGT0TwNLApW8/wLbR4A+8N7DvogWEUDuQTYFElZAjPVzECt/fqf
j1yK9lPQ0uDY5Gp9UM0W9RTJv8jY2SrneOMDJlWiNk5BA9kyc/U1ptj2ex1UHcjR
KqUZLbEd/s5cZdAUqBNesFeIPCMN/VPAI1hQDWfcLEiB3h7IPICKVe4iDYQi3SO1
zOIpfdKHEuiuXP9nv6Ku2yHjVK/I8VoLCNF89LGVJ1SZ5fuOXn2zK7bFg6u3AjtM
`protect END_PROTECTED
