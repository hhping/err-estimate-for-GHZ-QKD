`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+DAQmfcucmyaIR8oiCxf9kYMMXxHEc5HqE2FXUHvT00/lWOHoskgzDmALQvRf+3
b1ShVxoseJQWqI/Jc3GrGhQmPXHMABJO0o5Ccx28dcXB2K3JXnKvG47IpMHAMxUT
MmUpEJ7wofeXGa8bTy7vWM3RMBF+D5hgT+TghT91tR4ZYX7MznnBFY/LXT2FAWsD
6JtSzqIYswYl+9cPxV+juG3z5wDzhyk+GykQS853ZYKzQreFp+nQuXvRfnUNkk9I
PE2AC6PryszIgZfmRA6mIQrMka5z230bTV3GuW/VSzW0X7xG6t3Fk4HtPPqjWvpv
M0jCMUWq1HzvLzA+BduOwHwmimv64dCJlFLNVDUvC0S7vyvX7W3mHUsr2+kKg05G
qXioMc46IQeoJcFBV/9xnkQyEIhx9u4GPgAMYtvuPaZrW6PtgLjl+MMfCCpmESg1
YLkFHp8LUeJEHDgyoTXN/2xfDGSQeZ2hJ0YSEnXu3fRbkb+4bTm8eBCd8q/ef9jz
2uC8Fa6D3sdihAhYt/nHZI2s/w0KbgA+3Hv0gxd1aOO9v3VkEthkBtskWvpCjULr
EqBliA8ljh/2+uNs+XcOeg==
`protect END_PROTECTED
