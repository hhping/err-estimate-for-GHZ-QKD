`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1ugt30A66csk7SOkzhnpCAPxRDtyCqXEi9V14EmOmymdpGrLCE23ryJFsjwxRkM
vI8aYlltluyn6weGZ/yiA44aFBjF5WvhTiMjheQVd6s6u7BJ+0YIwrSG7Rrl+2cA
bhPhF7IOTE8GFoUqye5v0hhobNvFvkYQQd0AcF60b0W3pi1EWBzNgfieqVZC+o75
UNfRgGLBiLq5wq6aPVxmBBj8kD1jRX4qEdU3ntGWfW2XqKNEzZDtDuBvkPSUYNfY
91buu56V3NpifP3pW/RoYOz0L4r8VICW9yEx5NNmInBFH6Tv7fwWEvAF0ymvUx3b
6N2Pn4DNeUIIqu91bsB1x7yqIKrT7mZ0DGc9GsKWp11AFMz6cAu3OdIxWEezxSzl
1OcybiM9GN54H/mzLdP+rBdJolknlNfIO7HQ3EE/FkuyE8D310MPZlw3zlJA2VpE
ab9TMaljdUOB5Nta084SI1Rx4MCA3DSJeQgHR2kD+1YiGceuDY/RdyJRdKfLA9pu
XODPEAbeo0sjd2MiFGsP4zt4xMBTMooiMJ3+INUOsXjXtzBhQEHGNpfEk7Vl1hwa
CH3OghRaOlM8o5gF033orAFm2Hghk59kypHc6XbruT/eRCkRhqlPJneygJj2nP+J
zFA7KLFDY4/oV0VTPs5fur3pcFIYjQ12BeqAt/u9qKA5n0C8Gn18EH+dzhaAgFBk
/umh5TCnKu0/DgZbsbf9KjGpfZUY+FrHL9lDxwQOljjJzL9Z0GfSEFVxwQUEXJ4z
TBRh1PcBmqun2qMV+kBHjA7KjqDQOMlA04+y2YByOpW0hZ4lsmm0REhPGQkqeJPQ
DhoUQuebD7ZjU7pcl2+hA3n8Kjhi+6E8nKrIvwCZ7RVSnKIUHyzSAWwpGpML6k11
iIl0mkNKZ3Km291WznnJderJBr7pLSZIAlBtIevOCH1110qSzJ9xNdmy7a75Kcuy
0iM+ZoYvv6dSWymt6NtmUlN5TEa2P7Pxi+gu6XArcMFVAfiaty2PvgGYBzYh8YXb
E0KadTRM9oT+3XuD+5yFcxC643Cxa/iFliuy3VcFyOM3C7faHkK0w5nr68/QvogV
Gj7oHE6nIONs/Ov50T4O7BNit9fbkvBUpXoGfWgsVQMYM93VS8VJrNsZR/5mYRkJ
9hVwo43iqOpxMQ9wjj2tLCj8PTTkVeyR1Nlm0tJta36ygZg+4H7/gjEgOqN+2vm+
`protect END_PROTECTED
