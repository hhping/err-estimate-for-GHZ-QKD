`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JgBUUNG40UvIvuwYaiXcan7ew+z5kMojHM8lN9HDRFobyDvMBUdDxBnQK8veWIJ/
q/qsFV+6N5f4VIc9KIjIONN1F4rdL0P2LfuwFAqJxYz+uXxhuVtqPgt3NTg8Fijm
XmYHyv/V2+NzlFMaU/z1b6nN7UVl86RaoR8TbPEZ2G0pxkAgBztwTJEr7vFkxQ6z
OWR6rqZwZE6KS78xnlcRozV5ld8ywagV05CKadq0Yv3YH7ED9tsTDvyQ072SyO1U
Jvj9QNeW7zxul5RNgVF0nXBJGPtb1j1iuUpyOKMi0JF0Q7KEMg5GNZrSnPCKx5PP
oQImSfJOtBLPRF/Uee8DMJxkMI02MJYqnS1qj8V7jmFcJhr5pjCzUwSceOs4LJIB
6MfRYPFQIn/fK7c3wqmMYMws4AN92OAfW6a3mXZiY2EZpQKB8zt/fyTLxPhWM9es
9DQu9e0xeFcIk7kdznvTbFKMwRG0GsZdYePAZ1IycyrGVz7dCtKBeGS2vK0/Nm+8
EykYiF+ImNvOOyUNY5CCIi8X57USSmbdzcanBAV2M3Lczz1OceV2oTAjOV5ZiiPp
Hu424LUCrhZbntsltjLa/GTSQPSxMghXoVpPQvkRwyPsLU284MZmBdo0PQYmoo56
kYD7XbTWGJ9LcaK9f+8hJWyCzZQBS7F4i8q0mYmCwJIM980mHar8n4Kr1Sn9e81+
TZM3Rg0kuLYLP1fQ/zjH8TIJLM8w7He/kV8pNfD75C2/MNW8TYsP2WQOAa8bIkm0
lvfLSfDSdILoyzGaBZyaskyAlr0Sm0L197Ud9e/iN6mBe5pUbk2NWiDyjI7fBQha
Zdaqsa6ozzQKqh3OoSuS2BqHCWtcy11DBzKdKse5pSVtlxtMsFhado3QM0zlRR1k
AwhCsdg0bYzoivg6HHu3qm9P1eA0jMCNpU+dw/d4wafg/ZnLB6XYFG0h2Y+CKGsc
O1snMXr24uN+CQyyZLCIzI1yzGGrlUFay3e5hUqU5d+mr39WQmLsw7QreesvIPOA
HWBtvKToSmKhLA1pA/PF/uSkb5P8rlryTAyBLZ+o4oU1IklrsZOumNTWqPMCCwbx
Am71p9i5nNRzbb5WdQstrt13kNYl/NLAxPOrGDuSO8XdXnZkeNgMQ5rdAt0RwiHO
1dLNTVByf97pDLI15oIeI9cBPEXQAvfi6oZqosWhPc48mIuYJ68W2O86kBKjB+ST
M1z73iQBdVCq+8XTPPmm1DlUPB+SeZMvKhqluB8vcS3eUqAY6yi7IhCqWezLpdJt
N08MfzmIAgfoZYUzL3wTwm3udPYHJuImxpSxaqSI+IxqohdnynkZGoIRFq6jo3OS
Uq1XkD07AvSChGePpTVCmm2alVdrmohlV7XnRNd/rnUF+SxKk9+//l4vVS+Zef8C
duif2B5JbXXNinPIv5XHHnohCwLDFK6wHDEupLfP2BdGX4xrl32DA1EBQYzYUpUt
XagTO/jHTLqmbnM4R9T6cVf7enbD4DWU0U1KBBbbKhWfSxQ8Dd+lCYgSFvuyqJLz
hQiM4KXgkvA7QkUnalUAxj6ygmJN2u2MAO1iHxjiFRJgW0WlnGAlFjUnMIZ9DFJs
x+chIC4tjGJnAXRNhx0Dk0ADDyJdVzLxjKCWZDIxp+YAO9c6/SLjSDI28Nu6R9n2
6jWX7r5e0IOkF7Uubsie9IYQvAiSKomzV8ZHeP4AV64scVKxb5o50Pf1amqKg22B
58JUOajwmj+GkA7uoVPAr/DRZQPmxWdjnmSwT/Ax2d9SaoGmNzdgklZGglfsYqWH
wyhX1+cJQQ+LCzThzCBdU23lqfGPfW9CJt8v7HsA2G3dYhevTmk2Bw/8gpUON6XH
Ca9KyRQacGfoc5YG19ri5EPFS4KmGQpS1NTPJV5vHz3zi85cEig0T/bH7Z+5YuQg
LpHJaAy2DRtQw+1Vka8k70Mj6C94hcy5P3Sktl+XrrfuRmQaQjJkwn2Dqz75XvFL
wz6qPl/9/eMF1H5nMK4MSCllR84Kvg+yHx20d+Kj1jolACfUIyx0KEge1yHTa9LV
gyVx7QlXLpkNNE4YImiMfxkWrrbOtCfmN69JH/FtX7qmulNKdlzsY7fS8KMjhIu+
Vp/3J1ATFok0tl3ZCankphgQxLxZwDh48tjrHCM9jjIOLk3RJNETx2KQfr7p2MRD
LJfzt8kM3UVnCdbZ6e998zqudmsgA4IAc1TmjwNUNMzcddzUDyup6VX23ymCHkPf
NLf2+jPfwFW2BZg0aZXq/h5BhEIBfzgFR2e3YbjHfqZhjrMF2FjVdF5XKzNk717F
qHlUC+yLIl51Hw6cxZblbOF24+/eudtdDBg4F7u1+Ncw2kxIehtSLVylPmHW2lLz
OoiZFEIg6T502KGrlnX1jpnMwKoNUYhThRWRRrO9SC9CHTFmueXJNEbCWVMNFx8X
J6JL306Azb6ueHlV3ul84Xihjn5nKbX2qk70brUGynt23jolYZk/shiHqpsd0fl2
YxGnk3zvt7/DRKrJ+67NlTv1jUGZtYO2gNM3lRodE3zU055tx6j17dXlxLO0s5/w
msz4WyqvgokcTan4o65fqYbGkRIsp1Lv/22NR1+lPGK85dMo2K38bhD4bgvL3tTE
oYRHAyJrTIxoFBRhjFqYI5CXl2upu6t31gG2sEKbvgGsFyhBDFqcpDE9cxaIQ83k
y4VT9ZNOZ9GF095Uafiu7p7G4OV+0XzrVUmhRje6R79QwGb/pSkPQh5HGWC0gR1h
m+ZRuHHw8Bf9NEcwjwYkFnu3SkPm6g0PQLqhFm1kTCa1KdP//ZvWs7WxnMeHIp2N
0SnzwuZ79iz6H3KBkLz0y/TB1C7xHn5FkX3pDbX1riUCnxxR38oLS9smvG7ZSSQ/
NL/WQD49lTHRfYOgAmVfSQCTdETnmjRixXJ0K9DDjrdD3sF0M6QxVCdTGbo3HejH
i6pV0mN64ZXlDn/5raDfwJyIcGE8HAsuOz6l+MvPeyRduxf7SrWloRAwMdQYqgMI
7AuzlbdSu7bAwtWtWNd+7Hcl++HQunsdX3Z5BdR7ydj6m2SHZWa+8KXX+0smMBnX
SaZjNtdsnI8H7iq3XohDG8sY7jlaLDRfs1xktmQQrLpT9hcgX/WPE2Dr9Ybxx5hy
zlszVpHtxsiKu/kR8jpRLkyARvtcUEqQxIvJxsbDhP26PZxW7DpP2Buy6ApMSTBR
A2C84xBSKYg5nkVI2GoUqMAEso6mgBJ53AWqBtig1UFjmtyQdL1BZIFkL5SH+Zm/
aXZ854oP4r6Ccz3o13Lr7emLwqVuH1Pej6cw6kWXMiEfyn7yGfRvNxW7uKmzMh8Y
aEOEtYDLQMhsuI/p+ZiVXMX7gIBlKSiFu5q/xpt061vxEIElVBnmeTpNnij5Jpqi
O+9jtUw99WvsVWd4WpOI3qyMkim+qUBABdIXd/2WuC2/ODjRLo6EzTSFNnzWW7jK
Ggvm976+2PEy2hQIX+r8wdvF3PyI8Suk4fNkTgRQvfAe8/Ez+9mhHsBdmcwosoMm
2J/YkoBtFbwglIGDlHMx4eM5ziG46aW/8jfG0KcHkJz7pitMNSTScII9rbUc4MIb
4JyqmCNV9JV78eLqtfW+i3JIzAfzRvd+JML/ZXKtfrPHOeJwL0pW1udTFKGN5txO
Zg5nT/66b8eV6OKWaFvx5sJKzPkkYetJwEc3Fxa6mLdw3VEg9r4hyherWDXqAVpT
Lgj1VmVWFLnqjwMdctyQjZqmraakQw4NHBTiLn84R7a0/IVs0AplMQ5ka+2M+eBl
Q1Vt7Cdj9bFR5lxZeUC77Ls1yAFOT6e2Ml0vFzEsjcaPzwC49TpXYI2T5D7p5FEs
4BdvsrqaWMumptSndTFwQ7r5hU9R/v7jsNV7HjXF5uAHijGInbptUYfivd31tIYw
8w9nbHnbeJKJi+yxFs610oNoIa5Bu+/3DZySrRZ/geAOfqaO93DoqzqiKXckR/Y0
QK7yDE4bMysRjHavpV/FBFH+t3eZwuFZ4nc757Ll5yAVk9xt0uCrBCnNNrUfM5Bt
aIP12Onoo12WT8KyvYPUU0N7RTseCUxQiHiEI8kNOfWLtXjJ+s6Bvx6ImwMEe4C4
sAi0YeCTquqegoC7JlaMmJFUudcfWmx/kqVZcbHrh2KTGo8h5W8mQGDnRAVTFPuV
fb5A3RkudvaZ3YZOfWtMmtJdblUeyEYUqvPF2jTuNoJkqfZi7dODCKfJzV7GiD5j
zIGzX/zv6F3i4S8PE7U/TFqcXKKfbOwH9nLlYX9+8S0ijhwA0S2opBntIPCNL1Di
YDA3tyVqRxPRuNL2T9QjjMYWrDVAAZrx0106T3nxUao/9yuxs7xq/KqMbb2cGV2/
iMyytwpI5h+uG128sY2tj14kX8Fv2jVk15vGo7RzeMehYZ4Um6BeyOXwkujnpLbk
N9NP6RtGABLltDSQOnDQeY+abkBTHFzZoVTG826s062vY94rh6LI2DUZUSK5Ty8b
cHYHx23PP4gSspaYXaDJQR/CUiE0mcuG8sdBvxl6O4b4gAOBXtByI9uT8SPRd4T+
ix51diqxL7OOD4Qh6BkGYu7PgtQGA/ujSIwupoaHydWF15azCXsxBGQZcbLbXE3G
jpLnxxugFCiyRGXDQqa/kUVAgK1c1r02NYod5UBuI4oFRF9s7WAMXxeBC7dSgOBa
oNqrgZ7jiXenxLruyRytAce+zlG9rp2M8v0a0zzT0MwQ48gzuz3E6g/P85N7OkEc
qRLse1FSomDv1mJESszXW0zo4750vPOUSLYSKnqphnRi2AQp2xUX+FIet58Gst6s
mSFUp43vHWgkc+rRcw7WghBRLTB5v2zYl4u8owhN98hm4c6606pCU5ew+0Rht2e7
5YflhbwRq18cgP6FitYhZp6GmDgilkXDZ2PlF8h+/gBNrK/DlBoJvKjALo9mFaAy
rnMC+bmEpyq6WseiB1BAavdYWCgpj1Q0Fo7LFAQLpDsqmdx2i50KKY8v+1W3HqZJ
YxFvfADt5pBHDdjgCj5kE4okl+lnIK6Q76jJ4DFDLU/XmzbTT6gCV1s3nAq1XBEO
waARuzXO+SckXBTMhqyp73xCy+dKksOVkw49ej78GJ4mISIgWvhmjNgkoShrv9yG
Ba2MWfEFRODAfETw3ZkC3iMm7ulO6Xggi/nsWmWNrC3XVGmod4pmCO2oEsSZ2hoJ
iFJaAoMPTw4UoLmPydUmpgwJL4dU8C4H4KaGiLsRtLQBVhqtP8BCyfQrUz0UTQ+T
3JUu8pY8kS5Ut3AYKrLkqdQ4S9mJ2RCn1Y9KKaUOHFL72ZpaPOvei7BPDiZEGnn4
156VF/sYnUya+Msj63DOGf9br9NgMj8AHRtc0Y0RTVkokxKuV1q4nnH75ksyDp2w
l6fOQhstcJuZLbnK5Jk3r5oM/G4jj5XE86TDITBi/wQSfJxCsw8DJLpnvD5Wezhk
jQQHhTdT1IITY08/AhIf291H4WpA0RdTg29hYjVSqisvcYBi5Gszem0v0lcEBUX8
2ev/Vh4zSnLbSBAI3dk/lN0RjpY4I/R+RXKVIgCMcdnTjLD5qDjiWI/ezIiJ7UjO
WH7cXfwABufe9G8AkExsxvFq4+TyM4Rfabd+15m8fJj5CGKRfjuN0pRIFw5jEgwG
6QRi4avToSC9Ukz0O9E3QTiaCrOkOCfCcnLEoUNv6QckGfUXocFLkjKPnkMN053s
MLiV3P0nEY3WAAafvfhHM0Z5q9yVXW+gBgNZD3bojfHRGyyD1mc7fCPpVmC2lLep
2Xyuec7l1jC39TAMN4YtjVszOl34GbCi3KyTTqaXiJdgmnrvojXhhuj9ls0jKXoy
r4oOczQS49s3+ikPaqhoc7ZUY3X9+/A7RBOze/IHq29P43RrlzL9YTcaf7BlJ+mT
uGMEjlJ9shM2WcaN7gzERmf7/inkcx4F9J/Fdf4zuq3JSWPGuWk5lFZ6S7P5WSy/
YizZZEr0+GgMSySnmMekNQMj7gkj/3AoVdxtpTcNotaieXHVuxHFytmvOyXxbnNp
1WsZF+phHkbI9Xoz5rPOY4q90djogRIvlC95qHJxFPThvcYJBy9ptLh9+VCzmXPT
AuUfx2oFSJu5fldi8cMUkYge12qavoV0jsnqIsJ2mgx/minO+5qcIuHEvpCspAkZ
PrLZnJ48hFa7c2igNewmLG0OzGssEOknA5rtGnhj5MdsWd4fGJPGWejtLiab/YuZ
JKpVihYoUECPuK2iuJnSrZdmjrZ6ZybjfPN5d43IeQ9It9A3Y/iHUScvkyAQyxr5
IYc9N0+bu0JjirFmKuKRWO7V0BXtzl5XF1cqNOuG/BqQZwSmNhpBDwZObFFRDTNt
KLm2dJU+owAqBnK7w0SA/uAIvpOJn/wtmVhHQCUugCisof+lsZ41ld3MOPeqmZrx
Eq27aXAPeoBCqNL1o39+1rSmm9Ulhb6ZVHGjG81hDb9HL+3wjS0yQUB46WTSUtc4
3adfk8Tvrc9KgfplivuvJxiMpx/9eaWxVhwo2WwTsTt6wQr+vmw3tW4Ay9xVWgC8
etAzXEF800iZV5tUSAc+DqP3gySTIhzOiqumYvMTdL9PjqFV6DRHA5iK3EmDnXlg
d9oS7JO3/ofEFbzI3h/tlz0zLQnPCtKDpN/zk1eytvY5p14xt92Ze2qBzOso3u43
hTKC7brU5qu4FoCpbjyVThU7o3BoqtBfCzdiGzq7Rfk3jNvZojwszFUWTx4gbSmA
DleMQ3hmWGXUz/qMy9vja1DbE/5C2/vjT0yLbArQTs2JNftvMvFlKvTEZDfzcd3q
82KsUa5uej628z9xFfbo+HnMPgPReiLhZrkKTdgcVecrb1OTOFPDxv6kHtVdPROI
k8MDjMScT/V+hew43oQpO0IzFrLY1thvUR1RwEgLOmda7OaxxXnH734LT9Fh2ded
KGeCclu3IVnpEUweIrmejSKxyUGmNc+gOEzYk4wqrjdgr8IERLH2RKVfD9cujbfp
E2eg7Xdjn6X0yBrk7XT3nGy8XQayot3H3AKijRGfNVI9qhffLpPMrmn69jNFjNQj
4woWHweWFZzICgrGCctKKVqqX8T8yf9mV3GY+4r3Gmj7fspmapSUnhPGEYIneIJ9
Cm6eXU/StMPmHCaCc9SUF90759R1FUbzuglGW9JY3IE2Sc6dUHcOPQamami3ATio
1KPd4u5PzddA6C3MZzMqFXPm98YVLHkmRDGawo70GJjhG0/XBt3+GevYqvZluZ7y
zd4Fmj//f5Pj+fz4GQlEbhargUM3zW8JV8rdrI89XFypnxCOzkLNVd04WrZ2PHqF
2lNUGhhGddl03dd5DGifuZnItGaD34YWquSs0bOxrc5cK69hEttbFd5pwcbnu8fd
/sZgBZ78h78IOE2L/dM656ts6rm0Ut2WEp9D+mtWE6b2n4TkJ07yJ9WY7BamMfCu
Jm2vF3hNtAEUXXlLW2cAeoNiHiXDwf0/sj+ZCPTZmXgugiDKi1/7+enQla+H4cTK
dsmlrWprKf8vLT3mVydKZLfMwe6cfeEaWo3g2p5RH/68f3FHRkSRN4cIVqdgYtHI
mHAoEiRhWNPn4wLOeFfd98jZuqxPAFH49VOz5TZGaPy7+ac8vvOVP8FsLA/yzeg9
8zMF4GN9TeGyqlQHs7NVIxJstn0NesJP9Wgkcz4oerG4tJneEJ6bRtRTdyA0s7ln
9htn2eITOq72s03NpGrrdmN8ffjLcuKrqncey+GsonJBfHuxJSyzFaweZe1ruL4M
x9SlkrQsj85Fz7jJzM9JScZ6w4eiYUJiVEQcCbV3i8NfeD3SRu5H5F0kRuicCCDM
+eRlPqyUkJkMTu5gWAo4i1LF48uAuDcLuerTFIF9bEOnLoMKjWMYYkBtxvPwD6qW
SDFYAdNezd7YjpDIyNNp/kThyu6mqwCeAycx4XQmSY2/S3B6Gfd7T2vkbMDf6JQ4
ovK5sf8ArDytlO1gy7kh2GAHTxbptT1UiCuyn6HzmhNAEpGdJ0IZGUbUDCaA2851
6oam4F9TGvQTuHPEY4k45eUcod0EQpJFnd48IJrwV/mJ5MPh3/4Mn3pUKjZmGRYh
BYSFsCdDympZ+IUztQnvfwHrS0196VSfdt6t43p5DUKJJfKqj0+YSteACYe8Z2Iq
SP0SeGdnAOU4LYL/RZw3oNo9HsqjLpPCF4AribQJNoD3QI0TeGREiFGztlbm8y93
sDcVKu9Gcl4iM+5TxCCsTvirFGzCoo/2y+c6gxg996OqbU0SF+V22BiPX/2F25n7
HyNxMnK9aVhQnO0Rfp/PaAF6wfoXClN1tRKtTy5vHhYT9lvHyNwKDgnLYZHU1IO0
warP0sYtTYilyu4rbLBHGoBcyaFv7+MSRsj5RRo5pLzMkjs9cptgHOASlR01dJEZ
5I9bKnCdHeGNtu59dnoB0EFFcJSQPDyvMcfyHA0WD5b1zR3ghwbBTQoN0ILBFvaB
Va3/CL4wJVqtPdzFipuVL5ZdhE4sdi3jBgmp6W4gIe7ZgtBiRfgYJx67eXsV28lt
vs80c3dETC2Sb5y2Xmw8gJQtxTndKTv08B42QqgSwdxteJJD79P1p3DXkVMTFduc
gna0DRmig/EZZ9TkHScebQvkejXZTIsdMqaD/2ytEf8+nTtbZeYkOkmL+Yz+k5Gj
b629k1kYunDjrp5goxkjj7pOpQ6Rb9E26DkL7ACguyd+PEY+tKYN2RzbnWft/6Lj
rICKKZ3HCSA1MW984JDVFichULbNAKAiC+Rp3JB6rI6wW/3HJFeZ+MFbg61RVzw5
3JIehJ7982/h4o4OrM5Jm917029GKcy3ENeVmIpcRFrKSqsq8u0M11+gk3OCVYDf
6MsipHEfMbRh98AtICI93ouMo5uUXlk4N7KFldI9Pa6q6fxHxKeWSdTJqGKwDQsw
KwAYNge0Ce5UbBdZ29wR61aXbsOddAaQihWsN+9HDjw/j/5JrwtfPgj6aMjJxgGE
0kK/Wf6QKjdKhJazqAQ9XBcmRQrVsYSPPYxuQNMCoX3zwOiyNE0jkhGsKcyFQ6Bt
47hQjg5l6LVElafl1rcTVgbHoP001D8M3P3TOJgz40RPUViCCeN7Q4AtLVt6GH24
gx1ga+i+3Qede4fU1Tit5X5Heucxojx6PYPWj8IjiWDDnAv1m6GmhyisF6giiZeT
K7B2rMyCS47kIbzOwi6Hze8xjKjRQyxEuuP2oNOUa00sq/9bClQu8uguf2izn+Y5
sc1S/8058WlKOZYAvM1wrT1GY9Di2QTeVD94Sg7q7XJIFprdPyrm0eScIxcf43BP
NFhvqKJDch+W9FlTwywB7W9Uaus6SiiG2TrBS9t9Y4BrbWxSoVZEPgV2d0LyN+Ld
/oVo2qiJ8PnOS7XFYstwSITw/8vlVDr7B2UXTLgTLz3KKxnVvRiXNMeSxFL3cKDd
ibduKwYlxOnT/6AV/NJrVsNlBaW2y3dLCfFCkadrIpaLJ9TkC6UWlcQFI8v2gbrE
l1a4FQFdk18TDKOBHMe6/4TF7djBYxoFwubWjXzsTLPX7ByRk33w3Vk8Oj7H5Sy3
lstqd9ESM0rxz4gTt6n6KfPEc26JhoNiX4F8HKqFdaHIFU6paDretOkfq27gcmdM
ZkCyg9OXLRg2j0zwCwlLJQhVUn9C7yCbTSIzaX8gfiTr3ehbcA1CHh4xwUF4gtGx
CZq0p+Eu6/KtDSnD/88vrBzmw6lTdcHpqUod3aSicvL0yZl5o2FXd21FvnFdPKE2
+v2HQzYuh9ndGHFem2tpnJX3KBs/F1GpGgaYnhO5/yioNjETyH7d3cZep2T3/n6x
XfEjUExeu51JZcFEae3WX1pCaHlbRmOIRIl6LjPWzM225PeaC01Brr5h4R8LFuvj
v9/zAIxyKbh6brsRPBB/y+vVcLfsO8jiQTVam0jcATJn2Ks9mkho4gHqZ5/Fqy6w
SFAlDNkgxIdpVPicRaBS/QotbldtJpfmU3zR+ikO2r0fIlATxKQkt5JxrEO9j8TN
R5BCxPi0zY6YtHZhNppSn2HRisaeRFSHC7FaqO2eNr8oS1V7pNrBThifuophFw3t
2k117QL6+kyaYTDu1VWGZup64YIcjif1bCSAzayYRaqYpRRClhdKzRn/hbqJUWOu
ELem2M3fY4g/L9WxFUneKXSNSFtkUc2nPextj3ZE7dTnQN2QbjQPIG/CW5gSumgD
sQalN7Pe4T2222O1SPgP8azE/5XzJy8IYuSwG5elVDmmLXNv5kT8/IFa1vTV0y7d
1eUI+O4cGlqlJl8dCpqO+mzPKV1BEEsseOu9u2185DLFAxR84ZeEu2o6CZ8FD726
sFiRzefkIITYDOTfWXSv12EefbpbOvlLIgbM9xKwDID8cBlQAiWwoT7ciOiRZAeV
tZjcTO9G3Eg+cM5IRGua0t3NUH6PjLuGH6CeF61w01bJBeRgf0dDeHRdhdximiuX
LfpaGI2yuVnjfaRfuR3XX75uq59sr8CxWBGG50I34ETOESwHEwsZqVQyQV7Z0QdL
usmO50ijkyCcUTvDi+lYk0AT6q3e3MCEcVkKXikUp2XF8svTW+1THSomHJ+9avr+
S2vrNTsMnTo7aE8Rip2wqrhHkF/U89R+MA/gINlwsSjhlDeKBQ6WPArUf9DVFyB+
C++O8QJJgKVsv/RFMGuMVI4zZTIaQksmECzp4RdYkwFhkb3gnuO9ppdqK/TBqFks
aDOdQ8+PJk7eEqMky8bv2BboD3+/AO/Km81vUZsH0tO1uOJ0gm+AbRZlmVfe4CLh
G3U2Ymq1zY6wma20gmevjNP7gMYiNhRYDsCTLgqH4RHe3BGaRIKQz8wDQ49PnIYX
8L0Xdjp1A+PgvVzM5NAfeuUJuUz83DM55nYGSExuUEbPVbv0K8wl/3BPqZevcdtD
gKS3BSVZuxu4BsG0J169ewYEjXxn0G8wXtXsL/GdOr9lOe+lPgVaupkppLjTfgJd
I5ccvDflKEzG0ILDQTRTotFxmzGkx9qx0o1VvH3WGfPDdUAKzvqfewGTxQFPmUGW
sSR71XZOB0mXhmgYeeFv7tsjBETPcqRNeUIs75dEKPCZMHRoGx2l3YSIetSSWyWi
o5sbjVk4K/YLmGmzhF37DSxA8ajd+PgIZtHsLrK+7JaAlLpynFMqX3NfYPzmu2Yv
o3xdwYDCtluwWmamsvgpO3wXHUKR4LxSJmqE9TV/iikd9VGLBYFjbgX4tIa/IKE5
CQBqkTKzCoc4DNnMehmxt9oxhgysUuuYzuqf8J11eW8b2po5ecZlPWvs75fyZXXR
XkzbgZszcWwc+88sPejKbiD5ual1wuDNrkgChx6j1jxCsj7pH8SBJQzc+GR2ETUd
xEpmBSNqjVtmJQ4BwR6lNJmYM7lTQY4OzZx5k5ArPrxnxE6DlqBArOseklSjDl/I
G6fA59VTkX/bPFGSxbjrrELbGJn+OjtS3aKWqboF2MZKQ0p+bNYTfmU2tcuy/4NL
/br7U6ZD0zngeXZM3L8sb9e7FnDQZybamySOGQD84QDm6TtROWptft+Tzg0OAk1b
Ex3xkUMaZUZKszV3I58Qcso9QkShGlX1IrZVHU7fWy0cooALJMZiV2gKkXdvWtXE
RsDFlCINL7I19hMavw5R4wkVgTmNERmFTn24HyMN2o7miIUmaDQKQD+yQnqWMhSQ
4dFj4PIuMCfAUI3AG6V7O5Tjxf+x9N6+kzegI2rSTmBOW3XMxESt1z3BlutkP/fa
zKRjK1nfWUk+I/ZEZ0Bu/B/x97OLYwFk2tFvuoMhlxGUZVCyEwxjQ5MTE3PFVha0
StzzhSP4+5O2685VJEup2EHuw/MNGe0nkln7BLyTPNbzbeiK30F5/8qsvQokVVG1
N3R71Jgrg55PIUqFD0y75a254J1hMkK+bQgGn0NFyhX1OvfSnri3p3aoFX0r5uGG
yh7ThaiiivFz4XnylC+j2RG1LvaKJHo/QQNwtu9bsoGHtfLrhM6qSO3cw//hBs7E
VDtAH+drATSaWg7y1qgNpp1ke6TOQIsiB7Y/a+NYrO/sB3bcQmvMqv3pWsrWKqi8
1Q+C7OT1yaz5sFWWbaifvHuPHI9AVdaRsGGmL+KLcFFJP4ZabRIT0SKquTnBo/C9
izAHGRKBMM3wwf6dfDKZd4E6GnWW7gx+a1OG9xXTo/c6s6G5SZCn+BDz+3yX1kjh
RuFtMEy3HqAKWDX0lQUPwpKhXsY3O6qvr2tUjFG1GAIGPiSjY7KiuaTcH4bNcXxZ
ADwrzu53P6u30ACFsRK6jrYHxjrqqdfGHiS652LR5n2LTVBeVXJKrzxJSMs7G0fz
oNzmcXbeo0DS9xjKXq/vBJv/kPktAcH3dc5plzrgqxhRX5aVY4pToX5uw8/RIDqp
fiFyOa2TSrK+z4fyHVsfQdGgQsi0QTsMKn8DIiybbPKbfKIwDuCxoXWkAGByd7ZI
uFCj9T77jmVtC/eBw3xkJn6rqpBVPS1jQO4r8K62h/Gx/86K85BXHXknSL7xAgBE
9/7M1Yc9SySCm/vlQFMej8aO7RFIdq33U3a6ujgLqxeSs7PeNX8JzSaiBsIJpD3X
0qhmicm+xPjYtE19q1nhD+8LtKmJS1rxjRKjswlZFI8RijwG8993lF+rVbMPKHx2
k9304VLw6r2dEx9AM7mkdFjZ1O8gox9XpjbR+YgGKJ10XGLDYtvwLTBAXg0LSJLg
Yfqop8HxwqHqKvBxed+2WJQqeNUs2o8ItQHfSIVyRIxtl1s8479UsC/zAY3yYG1F
Cu6YIEU6uoGRkdoWnm/8FXQ2lxv2ETrDvX6FdJ0soL2WAYxMYA1bVDZZYU8lj7fz
w0q+31DhgattLgYYvl8OYJeEUysk+/PXgLlk3n6o2tUKmn3BzTditlbDV7BdVjVd
4WwX9rp5llBUWpbDxPC2+i5gQz1cpe2WoDgTIL+gZ8gLZ8qhEcTrr2KSVnbcBMRs
HjwjjEb4+bRSvL1i4iU8J+BrO0eCTjNuxRolKfdGUa2rrIjj4ZZjtlAiBQpUPvw0
xMMj5Qm3le8eZ5XqyxS05giR8VZGulCOeoWjDredF8QYvYrAAspsQMgMYAeoUPIh
5UBGZNqUddwSA0uU6MHvLuTgVOWZVpcTu2YZD2HLlsLCM+Tx01cThyadIKjrlFFK
Zms/ccX48I6vJNJAcB4POpdzHMmf4PPV4F1X6XJ1UzdGNgvQoY6uQwLFmKJABW4I
5y8eY4Z5fjqnMFxn41RQxA1RAUbhg9LrEd5nGU1IkqhM/+elQHf1OgGZDfIhcsV9
oBKZN2Cz+gPnpBwekQTmGTdbSQUSeyoQ6Fl6G4KVk7GFsthIH52WO3g2XlH6diqS
CjbPdX9YSR4PfHjgsS/8qIu4TW3r1DRoqWTCc9EAQEdx/R1oV2E9bZ3lwg+qTGiv
8gy3zDAPqfhFkp3BAGMc+bCqyH+XPOHS1ovpmtx9hfZQiDWhR0EnJnpt+x+4o2Oo
MX1817jPYo0XyfueI2+p3PoxqQyI2puKst3NVftx4y4SPdTtlkuoMnOUljdG6k9X
dS6k34JaAn0tO13hpJHiO0lbOm8RjDE2UN9037E1oDICv7Bibp1VX284CsP4NuGi
Q1dXSzvd4gdVS/skXItT7VNbM4cSTqqWCliswIn08eSUmUDHRXF+GC61iFMqmdB/
4f7sXEICQmoKU7ckSKxXKv6I8teNo2bvcucKuEdjonU/HMBQhH4FQqM8VInPTGq9
oFiUkj8xayYy5PWyhA0hWoG9vU4XASMUodNHMGOmr1ieYDUMyIQnCypPHhYcfC8o
xA0Tkv+EI3GaSJIZ174lptccJcKNtBoOSm7iCvnR9xbrNg2jssmLjx8rbP1W+LDP
5xC41p0OY7CIT/UhMvK+NZFD1naJ4RhPJO/TrlzgADzsSEsyomGiSzqkksuBacEj
gNkekNWaVXeUnJKkBCtZDAvtIliQL4AABcbwuU00zPGrHzyiw9SAcpRdaNzNVUPR
yAwA1sj/QJyArU0oSiH4U+/0tAEGo0MPIFWxBPlE1W+9snUWiG9NsFsOHLBOVa8u
tZTv5Ad/5D1wQcqe+O5j9Oq0yaboDHcdd8snDAu4efyECTPw+1k/QdtSkcf6Kt7h
/jL19Z9pZmCIXLnCgjduXBbFhrpSioL1Pm+t/n0hBklmOWGH+oU4JU0/VBzvgxSt
nPS4SoqWwGzrmAwpW3P+z2ZPtT8N1mB+pM8ApkWodZ5prhXv2NER7dNZ1AlVECug
PtauUYytbFcOp5AfVwd7iHeODOvaexV4L+s49DRRUbsIwiJLYIgrSjOH9YruoST1
OXu48sPAJrVfMU+n8tlDgKQRffth6pWJz4EZusCilfeXu5FaJBbBjAv//fD3U03m
55kOARevLHiLnImvZTihieppdatrEVs55CLhOhsFphMfNiRmxtwA2zNpx4UtZdGt
NKH/9l4XSzrH8nt5vmMt8FtnYy2IwihYarZSdrpa4XsDUb7qmSd6z2ACpzjGBh4N
UgRhBzT2GAkMaFkg+hVCMTUrh5XLH6onAXDHXMalXKq32re8Nc1Of1C2LGbCEhnW
pNLETDIjs3Qb/Jo2m4Ru1Dg78WS4blhBGVHrp911aY6NnKmin1tAe3XBVy4N/ymd
+08O7fTB7G+FyShXwoUw+gOW+bvfGvAMR3IEYfbCw0i2Tr70OGujSzB9+SjlpObV
VbWXm2W0R2ngEsRJeLvL1gI6RZAh4N52wT+8teuZ+rDuSNE5gfsLF+Vw1gupbLs5
ipLYab6iozDz7HkxbHS0Ybr/TjVhPN1pA5mMy/J66QHzMAZn41OZ/mXWm8B+fH43
OH3ayptXDIvVDfgTIaCc2QBnG091iA1xPZ9z1DzMNXPYKhAd9exxLqv9ayK7vYpC
oaXdG0z6IU830Rwklcu3MGIfXPeUFM7UlKu3SjtTDB+PvgHMZZuBaEBHBnz5yBFZ
bWbz77b4OZZ1jYhJRZTosdT10PErb71i2S7Yzmavm9ZIh8KrDvCLcCxte1tqAbUR
FIQMv9walMqRKhZI+7gYrUBVw9MjALpL2kb3bXAnPyJygrvXPEmwU4JvkMkrP1kG
ccz+G3IEX8rh0j2WdCJ33dNTiE2PVqus23F+Wbu/ljMTiAZMrTgC0knC9rtq3x9M
KdlJonVOxtUIwZOwyMgBH3zQL4TdfWmQ3proXTwF7qDSC96dDHUSI99ILDLzVjXz
avBf+BDQnS8/7i5Y/3aAtIkaxqJPOEUe7odY2xJaQ9hYE5z4NMU/eBCwyhBxAqTl
+s3TgKVx8bZeWklNNYhZavNl1dDHAQ5/fm883NVN094LO7WtygkVVu/h63vBElr7
GFaOcO/t09z0t+WYPOV/R+loPPNcQ6DffrEfRxQF4dTJu0x6lMBQSZjZx0DHQo4d
zmtHgCgioU/T89BS0or9ABBCVXdOweApPTg7/nXkTnaz58yW5q2LxpCu5v6qkBmq
eyaJ4z66zQDLUOJmR1jrhsjZK9nPtcd8ao4XfdM/rzF1+ySqy/i3f9rojcDCzwmI
u/WkLn/J5j+5Lh/x5R+PSNuY18HM4DZMjmSANvXo+XT4NLaYaMuWehWSTRt5oHwe
UVi/elXALEN8UxbrVFWIiqU0cEEGmxmQVLWB/vaL7wLIWWDHt06fxKb/vBYPGBeQ
xXiJ/fK+N3XA5IBBybn1Ih1gL3nHaqnwhDqSX5MSuYmbYVtIgGvTAmvkICsWc52f
slkXm00NEYcRLiYu/7X+B5WdyoSFdT9pWQ0UK5n4up1oDHyawHj4pSrcXSnvAd5q
YcJqhIUDG29K++OdYxUPBrC5h4QYQvkqaDuVY9u+FLftiTjaZTXPBA6cktUoNwfo
qPmgC5xFLGkqozbWGSSbBJXYqcHw5fo4ADBoJNHn5SyUZWCjTNe+gQbIvd+b2KiY
nQvfXCTP+SFXajqnNntEnHuEXDfkVP1lPNxxkMcIEUPIIxmpJkCUzy7Ga7dQNK8K
87OtmkF/aLPRsNPyLHRJJUmh2E319xrh6oVqJxabTOZDIFzXZr7milzTOrhodrgW
+HRYBJsoU3kwqyl4krZu4mIOJBCCdPJ9uBnAzp3s8qqpVhB243XlkNCtfxh/jGCF
EFbe6guw0A+whUx+M5vsNtXeNIi0q5PhfJZlWe4LJucxKoaAoTfXHvE5LqbgAWVE
5TEVfCuqjiqfQYpRXsILy7njwTyRvKZVh3ui5sgBR0evfej90SnQddXDwxVndmwJ
w+R0089HzlqC6yIaLlrm73k9uKLi7dlrlwEFW/x3sd8wukJr3z156uxVNH6kM6/S
FzgOUayuS9G7/rL3TBz83WNqpRbI0UZFgIp4W+j198WdkkPXZMFSe4IUv20DfjiD
TOH3XNiLmRS9NcRnY5bREKfDUuxylQZszurVHGSkKnRW1ICO/+W+XkPqC30U/dW8
2oUyc7nniijk3CiReiNt2iftspsof1aV6UkYswtT/nQIaOYhHZDgb4g3BsmgOr2y
fKL89ES0+0bMi4vXicRUiEJnMhSfa5tw1yF50IzR8NWChAnXjhKUwyhwPDDSQplA
ZuGxXw/Y+4xAB1579Uf9KKpCFpE+Y8eqEYgIKpj2xJEgs0ufQ55KFaueCi92mUn0
807Wpr6tp2IZVG3AT2dcuoqgrWmOI5WSXkx3MZxxcARMCmCN2Wiu5AK8QviUfMve
ekTFSTRvEBaq5ERvotkJZUgfYuF5u+Dj/8D1Xymm7oVdRJsq13Nsm1Ng5ddke2zk
Hhlcsa/pUBo+4EkQ6UdH9k7L+LcICnc1P+DuAhdRMiYGpsrBKCpAk7BTxACfSsST
SlB7+LySo1tzwSYvXJXRw+WYUuu/IvwvWQ2wPMYcbLA4goJbPwli4GFD/zEFZ3Ao
Sh8OO1CVjnW1u2gJWL+1dW/wg79/juWaVESgjRKewWrZoEM9u0iydZ4Ch8uVpnPg
RUbRTypkJmNoFqKJ/c/h1B8VhhOOaAbana9Wa2tQL/iyplQ9lUdmU2mbVu4wH43+
qVKba2e77r7Pjlamt/ZjWmZYTJStWbsRVygtf/AyEpNnFhLdPm79NcljKsBiOi4W
o83pUIi3Pgu20pCKlWNmp5NETlXr9pfeCieDM70YXSto3gwIDpaygUokh4E0DoiB
ldie6nDkX6sPk9LXM1Ky/xrp8+jyZRCBHJHKeEYDmYfr4m0DT4O2RJFg/3yTk5F8
azreMUW7BQmKv/etb7SHFUWhmFpRdddj/w7/cTzjCJpvQ1bWnKl9W2XbLNLKZH8u
AYvj0XbEUkpEvgbwasgJPnEt0glnH4zrWbD8xTnPSpdF5KGl3K0jZdCITrTHtPTA
K12O7XISKWc+dVeIlFnJ9ptd58ZrXCjNuz6sDGUBBHx2SNiNtNrFsGnNczqIsklK
REJQ3I5IwYR37krjNCNxSCDk0BUXRaOptzZQuaecjHeJtj9HqC4jy8JOR5MuiAw1
MTJPJuVSQZqtcrLMZVLiBrHm5FsYgY2yQglp4q7BDwgQrBrwA0szt1N3HVLdV4hz
JyY+dNEAlAQyA1E7dUZua0wacoCYGUWgdLWfYAArCUkMRzqgLvWOOrmpARzXk20l
VRlAOhmJgIH1wx208PuwoDZsiCfo1cUHbqXFOx6DkM5ZulL4nvia+VgM45jXmHzl
tZ1//JzuILB4cSSC4dEQYPFCqQeP297kOs3V15nHxowZQ23BmcGwwIaP1AEi/4jq
ewNXS0hd7urFGgPoMT/It3ecU8kn3qn97bCS7BjSegnSFtOjhm+3xdjIRaxuN3kS
LFNvx1GdD3nBorKy7Wd0nHVi7/Ci30Tz95NmKgiBgjsAa7R1rHDrCwEnHy/2fwZb
2dSzlohgnxMTyHwJCEzjiW6oSsN1xIy1IuMW/7A+4hO8FQ0u4BLiPzX3Hsy3tZVj
bcyfelGmIvXSme8Btzb5Dfu8EgEDqqawRMZ+qNvV8si+sLDyxfIcduX37Xopt6hb
5E6gKBkqhxoW+3lR8Bd4FhJyLqk0M2m+yDxekqucVBrsCH8oWpS2im0t61lV7CPP
5XsdcuAPyYjddbcXP+w6xb2y7tyVrQwr5BlTBKMKw0PuvJdLcDKScbuZw7fHCPin
L9Ux1VyPf75F6/xua/vPz1AQLIJK4kGEd6XHxRmihy04gQ+tBlQJsRHcwWmSp+A9
ql3Fw8uGXk07brp9vt35oVNiayofcc60sC7J797sreNnZHUxBauhh/jQ/ISLtOGd
5SAY6AuKUs9O+DsSfuzCoNOmpdw9gSks4POrVebgImRXAwANQpI03KDp5/0eUb+N
oQMYa7QkSD0khjmSS91sR0CiNOmo4fGekJaDc0r6E12IxRZD4KoqFGupDsuWf9Az
IPklUS3anD4wbxab3OrRZJdCRZMi+uyLHkGF2RkO94ZLimDAALRtpgT5oxwPxnja
RtNzYMNHG76PoheO5A1jbzshzF1dcqQckrBfU0KrRS3jfRn/pB60GLJmDSfOfCVR
dI11WhOClZvTx85SbkYVX45Uw10ABE6wMp0B26/igIRwbMqrvf2UvJAz3egyNKSs
F0srIavecyecLrJqa2Wf7NWDZ2jXd2svs5IwlWDni7b5WDBN24C9/LHKejbFBOUg
wmonBITE5ZYynLKT12zQAouECFDZRRaos4GcjkTRlxL/VhQ2TsWzbokhi4GJXMC+
tYe+WBb1jR0pBHaenVZ+kDwgws73Rm0hw8MFtx9qRuyuhuM96qia+/B04iXKDMs5
VNW5e+jg3OUE7Iy4V9BC9sdlUIORk55ga0aMKyDF6hA05XabirV14D9AJ+XFUTNR
5sZYaeTkIPjYSfBFh40ZpADFxvvXYCTog/ba//zvTAvS9/VBh3i7dRaacUoY3TdL
CQH86aQtCTC0E9RjuSsL6Oi83e65kw6etK3uVeA6ToYOtbwlcwDnaFgHnCn4NGHf
aiF9klhk5W68KSPI5rMjY8YIIN3PUHLdxpVuHSzvprHmVvdfOwbZfUiXOIy4NuqR
26lnTPJyb61b6QLVE1RZhO6sV4fzlOWgCG+XGnI7ajRBRBrnsguY3K6l4kpdkXpa
kStrVXtHMwDLp/0WaqOVWzenFJVlWh+ze2QnnUv45+R37KJSHNZ0YWt0gTeKqA73
xG6v8PZzEOoBErJYLMNz4+ZRPiurCZp6MxWg7hbF5IX3LCwoFwqrKdHmg9m12igX
980VI4YwlqOZRI2mS3jsUwrORNost2IYhVSz+jAKwIDuOz70FcIi+9sSrm0snKIK
IvoeJ3MXUjOilV7IZ7tdWhktE3qdpIUEoxw6ClpbdUr+JaiIipG/2wDCxq68wUUK
Li295AQceRi4o0y+lB1N5RPABbuScN45w5wjuYSf8b44YbrwmECrnCSz+1rFxSp/
Ot2C9XUlYm/SPW8VtOGdy/JsV0/gV/z4CvGlw6A3pyj3P3B72TjIDHuK15lFTINs
7/4QK9IuZbnvntv5TuZXVBG5RP3X8p5rw2GnPCVhz19LT+p8q6QFEqpGZdePSQTA
ykjvaS3G8qF8JENavR1bw6Pu4tnW/f5A25gWHpcDUMa60xj2bcnjK5okwUcREQR5
+UIQIGMWrup5s6GGlowsmPIdsxgomxq+HoIfE7rUmToEwUF4wrUk3RAc0Oj41ZEc
dvF0PMrzVzZb2ppDo1ZvwqENTY8TxEkJPZWSi0EfoXcC+FefDOaNl0V32Wx7akP2
YQFGUwKai17XHaYDO1hXv155VHknLuHzY5m/BwFgEZUuaD/IbapEIWoKlFiyWNxd
fxxSd9vOL5367B1XwaZbDxulDSnhPyNHTVbIEyu5ScbsrlytvBpamWSeNUw4DaMW
veuZ9jTvnFeOonjvbRrdrTvo788StmAXzD2dvYyOw4r5KOUnD2L+TwGg8/8VnLRw
23vWrpe4ba+iVBybGmhw2kZDeNrnd5TJGC7rZN9+XMnsGYtKxrXcLT9noQlZGpvU
/5t0dErG7UyK5UQuPc/ila6rKF8lExanf9MVo2sFDhbuGuucQ1X4xzTEvucAbSzE
fB/3cRxlw4Ww9rhL5JUwlgLxZnlsdIqB0RNBqP9w5phVS0Rr6txosHubGGatOxc/
OQwNXz18ajYo0fNut3hlf3/tbIWBP2/6K3xpDzKMZclugtmqs7mDzc0+qDRmsgQl
dBPVrrNtAO8SMvE5qWKIhlr62TTi8sloYKKEPsY3AbxQ18dJWPKIDiyAdNYSm1sa
465w1VWlKMD+3hNYS/02uXNkTd9nWckJZ3PYSLJg29RA50kmcJMM1VTuzVi+9cAx
ONwGMC0hvZfZG+TtxB7MxEtZdLkeZxQYeSGW4d3ChJMlWD9mP7jVXHS/qW/bUX3N
j+kBNCVYsNaqi14n50qAf0fKIK58BzR4fWOTj0oe9UfnBlz+cVQaIi+goEn/7D7U
GPo+VeNPaR3QClV7MA/ku0g231iXbX4RqmXKzffeQQIDz/NRQOFxFc61FrVMb60U
fPQBheZawM3nVBwHgs9ThAm1V3kukiDO8jbwJ2w1FjhbVOgnI9rwoIQjKqidoMAZ
RGOmoXA6DL5QrCzO/lsrFoHVLylrKE8133ftd8mp8W7qMTWFYeWYvQvNwcQIf4E6
LBR6iKR3eify78pwNLKPOQvBcZLojDshp3+DwN7hjIetEHwkJ37mot8sqIwoFQI/
WEn9eDkZG8VakH/2PIFO3U1JG6JduX5X6Bv+AgCVGVb7pERNvapU7WC3bbMc7ZVV
zqTMKQQEk42dsN9sW1w+SVGD+ixvJQKYfkXFdjJFIIXo0GdRN+jk+kqVI7S5d9Uj
UDy8RlXFr8C2dwQXxoU/BX5KkYwNjohwPGpNSn55Gcld8AVTQ8tJcNsRkHBwlieP
lKwYv/MtMhLFTWykcj1jJWQQueQrdm3Cd8Z5d9GzE1skIoGXRf1dbksm4BxNsjPl
s74lwtxRdlyCzhK4tb/oM3xCYPfZyRW5F0FodAgiX1j8dboAagpnLx8dY+KkD3nq
BBWTp8ijP5nzjPAxdr5ZZVh4t/mpehTQE82sGc7gWVyUTdf7AJBHSF4UbA6VEccC
DNOqVwpN5jqI/VOCwhwzFoz4Y6LD+pm0yQr/DbYydlaH99psZk1ajPG5knlNKIrj
C6i0ailPbUGphKQtbHAPSV4EwBV0glrg/k1+IczBuam1TjqH34nghPvPUAIqZkOT
uAqdNaOn32cBUL0wsGNDTf/UCZDUWaDM50oJsgdYvh+0GbsImog1vV0+u9gcBvtM
FkaUAI6IhMECTCxhvGFZqLrK737+u7cLjNLlBEdJUFm+2JAcVHtFbPYQmplha5ev
UnsaVufSwqJetoEhtAUPLYfzLay1F0j8+3e13GhIW0DmI+JsvEUuKeBLo0rRHf4X
+IwxFt8YmH+6NOLeFkwY9C1WgCadS+Lkswl3DlYAhcySHfHEsOrti8Q30YyoQ2ci
I/oALwnLBgFmMs1EO/ZMwAPX9T7lm+SLBnQecAV2Q6cc7gtkzgeGk3kmrQikHIL1
v8cas17IYR/Vdy/qJjvrDNeAp7RSuJ47fDkji+S0ZGglRF0ROEhxJ7tDO7Wr0syu
IFS3+76GP1cfyW8JSl3nxTORcaUS4NOe7gWfpcn50M2zpFBn8XCrEyeW7G3gcOss
dvSXB1XL3tHjWL8aImUh5HrpAfAkaL809ToaX+cLHXBhmR2d4INLdeY+nEAEkQVk
GU1pVrqnhtqswbtgk01nsNWkC11AXw0Ymdin6UVPdAq20es7DexyVnSbR06p8WJb
K15ArTd1HjlermR1MIrk5SJCU59rVWx6r5MzlLBgstbH2Zti6kf+DUcu9ZO2v+kK
hPsTsk7tnxrSfwUZ+N/SLQwmyeXmQjHQ49cHp5yGK2TA6MIVM8Bqs2t/u/v29De9
TzTkQKm9GEraKy17qzJhk3S/b1Ae06fBPoAv9A1ouFmGJvDIv9EoW9L6Pfrijbq9
0O1fmOGmP0wNso5lBjoAeHb/2iK0pS5CGxHQr0yUQMPABIv9IdpA5kWub72QghPy
ihxJNLqiwG9zQ1Xs8NEomFfs+qzAG/Y2Xf2buizBdv0YidPGq6fdCtT4TpcnbwvE
7XSJv3YwE0vA/ytPnPBLGmk0QlCXKrtEsDHbZQNBB0Ug4g+wqG2iPrN35TTZavci
4dhGpMWeS8p/6y3sgxAekMDfU8phLEIDTLQxRt3ttcZozVRv9z4iLk6vb7KA6rdv
XTixassMzj2M8mYHtXWUL2MzuJojO0OSRVNZi7ri8ribINaAPckme8nDU4L++mH0
c5EFHI/0VOg/qSgHrUlxQ8qv5IpIN6jCQ1mVaQHwZZfMBpszvB1dcH8HC4azR4eY
S4D3NBDnkl+zh5Lu2OTJVZ4sJvjhtShM7Ry9CvmDfJfLmF0YhzvkkRn3YcZrbaDy
LveKkj7HeHsPUhvX/yapAT0ULJC9BOTMwCy8Ip7VTbtqPHAApRbVb/1zFubmNutG
67VnoRIWLq1cTjtGJXuaheVxE0+PQWizKwlUdgNdr9Lg0Dmr+kx+tvThkAUzlMOB
Lq4b7aVDDaD9btdKu90v7BNpkxapXUPNZFyDwvGu+JCtcOE/GAghTrUO4Lir/5m1
cgmgAYoYv13uRSZFcmm0x/ZWdJkjHvVn9bpYBhYy6ItHNyuiztLzXobHRKqR5NlJ
pjboC4SNHkoZudbVILN2wBY7dK8nBiYd+R9taqL91cVgG9IpVLzbuE0OW2xd5tm0
0rDYOi3AuWt+aVNWUDhvzlQdO5Vfu1AsG4coklZ3N9EWgYdkDmzhLL1Cj0QRz+T3
dnHvN05Vj2FueNdGSpPGMZUoncRmBlnhmOSC2UZl3/m0Yn51JtceK72s9qjktoBo
prYhZy/Tq+b57+FeDzMMgrwJiMR9VKqLz9gH7NhB9iv6t9blp9YVvb8t14WIhHFo
10UrLCKkC9FxMyBIgfj7a83ZaXdshKRnna/mXpgli7UMuHdyeHqQhnHy3EXJ8MGH
wDmTZJd/4So6T0oNSf6H3pMApLWDNhxUbUpY8cWKyDptG6/ms8ja1CFWUxJmlZ1m
4rGMg/qOXdICUwjimHPnjniCjcCL8FG95GdqSQ4KnOQHxWSIFjjgiTzXP4TLTHro
LgrxjC/G0X7VKdYaqX2WEsLqVJTVkqZnuOk+TtU4EN2anaaN8qcj9CWlQuzBm5GG
htR3AaAQDqUkXhEGJl0O+YcO9xTFbRrOsWvlekB1Q/mbOHf0vifBfW9b6/FRS6fa
vE2ZpbW7uU2HCRg828O35cG4syMrNgxjZ1H/LVxc1XTWPG07x9pMegb6SpswgZNa
ykjbFaK4gxaNOfM0aMeICuYsGjr1GuZkX+ZOyfr3ULKrU0c5++B04cLHo3TD8Ck6
gMR6zkOxyXCBp9xaygV0z5omV1Jou0l5Xlq0ZRraDV72S5+9WmKsGdnYzSWLoW6Q
Tyugrvr0nQXt7H9EmPWQ6yGs6bMPTQG6xlFOLXLCErmBas5hm88iCBQ9t0QhV5NC
nCM2XcmLC+0NB6CuHOeH6Q787XiQQoKIyrylGldcuMv4i/3HTCxdX0gyX2qG0mr3
bxf7GzTSZqJtjXPWonjHclAs6C6UHEHUgZ4vTA2UCU4TuPP1hrh0IiyDiDqRZwnI
Tmu7U4CSwDzngRQ2wk3PZWb8U5WaiT2P0zdCJs7GLztoyDJuqFDDX+MI+E07BKKU
Hh3pHHdAK0Do8VLl936fMRiqHNBoO0HeXsvH+Ed3pmbscllX6NBC9Dq/VA51SiBj
1/FNUBeC85p5gqZTY99k/ZaAfuvjbPlr9Gk8tjR5HLJdkEow3kFvYTnEJuV+QXcu
vCL2wTEalYAPmMItB8gN6sbWaoR7HeIM9xRc1Puhc6485Mld1Cag084pjibo/Ggp
F3aHKuGYSuAIS9JO9l/war7OYGplaEI1ixuQTh90AX9CCBcyO8hFTJ2HCD6Fz1Xy
tsjiNzo0zaTbrIBFjV/YdjASlfSMaihOwAmq6DPKsupNT1HtE8FqfWfCFN7MSruO
QbCmaRXH2FMmEsSz4YZiFAFuhZiuVFVBmr0Y0hUPCWGmOBf4qdRNIoCelAdsr0B6
c2HmAIW99xtFL9XUm7W6vujJyE6pzjw2azHHeGFf9gul2lbbTi5ND4pPZDKjSiH5
d9Py5Q9u1hmzIXzM2bQ6GwhIhjjGQ/uODxFG/NTHIlBAikwe90zm70WRW121u5St
aoYTiYr1D9Bc59bW1Q0o9M8AIpb2pE7idnhwwLNNSSMyrtgjNPCpP/ct/qtS1+A5
RefLRp7M77zcB+ccb/O0aLkxOAjAzjZI8MwYSFPL3fnoVAp9AloOyo6TeN+s2oT7
KvBvLFOorN/nlZTJs+6pvyAGWquiGY1aU7vbUgQ96z09v6Lz4NqRVWjDTqcbxm6b
yhzCAn8Dv32+25QO6ouWCBTkuRWQ4T4967nWNVGNSSDxwhE3YHinkZr/ErAjfB+Y
NHVm7RP2mkVWlKZoCavS5kl2I9MmO3qWaxeLCLrJFNwP+nelGKeE1FFeiSkoXS4G
ws9fiNZzBmhe2y16okwu9ACLpE3k2n5TRNEfG4gZc40iV3noWDDHE76Xd0Wq6yA8
gFVJF9+ng2h5oZGi8i1ZHxnZxmew5bH9tjJNCM6F0ubG3e1q389QkMbbSEGG5U8y
qa5TuTLxq6zwNoMFSWwkwsaODvRad60ffLjzBoWtxmiyRqHA5SWWR1i487VAfP2u
FIMuiESVTD7ZMyWugIXZ8y16eGfW/cfK4uA8pDZ1yBp/kL/YRfMeihNIPm9+iIR8
G1AlWIWWsAxLrx/orPDBWMiaYORtoBuDX5gvhv0Ok1uJciDz+y9cz7MjCWeRiGCl
Sr/wl0hxEHhN/OZD+Cg1JodF51rdinF+QfF0T/96MC0pbDZuk7vfKCkS1X1kRHxo
1/ALOT5Er37TvPTMSbusaQ/QdX5cqbc72GKWUde+8MFgQLjAgf++kkquyGKNulu7
IEYfVXKgdokjsTh58N/ktr4VAQKd98f1ybveFVgBUWANmCSW51s573xZaiCt6Kxb
DvJiSfMiynHbgcALF/dqU8sDZnXcfZX37/xzwDoybrjQjpHyGViqOC6MEfcarMbX
QCiPyqtUtdAbS7AyEt1u3ST+uEZmZKMD68W7OnYs2LkkvbALWkYVHnuBGyuJqzYS
UqlXATSLwIF5j4WObue44aKi3vjzt0059QDCaPZIDI00S0M7urnXH309u9AieVHM
RhHu3UcBwzRkd5XGYaUNQTQqfBEBJgoAaZw1HASDBQgSP6Xx5osta/8TsNoAkvJ8
p5oWj8sX0qray7kWfeD0By9G8BklHbFZr7+vuZwRVACI33MtgmU/dwI3z4E6b/Y1
kOOsipVvH1hKAdwoMmQBPwZfI+U2C7AypftJNyQPaUq5NaqGRWVFViF0BmiLHpnV
ACSmdBN1cf8WphRhxLPD3OykrI68eAmTej+rsy++iMIPzZnEIl0fBA1tIKwHqipo
CRTaoSLXvGIS9MiJhLyluYHtCFXi1S/OLhjDkgxJzX1i7wRWjywoOTWntJzINB7/
OZAFZPV83VbevTXtkyUMMDt31Qk4S4NLWHMNOuQSQsP26kP6KjoSjGXfSsAy8LIP
J8WSjginvi6TZFx/M6+M/UQwnR3ccYidd351mhD9c8pWTUK2oDLrmhu+OWuN8mez
iJBaIlK97WnN7aPcmoGpOxmqQC87hHKonPBP/KXOgv+jd3Tsnoe4pcwPXs86JSSB
VP8P2AyVYH1wzFdoqNT/Q9IQ6NxpvUEA3QehYsqAIlQ5vvopjFo0MtvFLB7HgHsI
zwWYBh/XW/om90WGEpEZka38N6Zi5DwPeNrkuGrU88QfGa2AefmZoUDsY5IY3vln
Wdj8jYWFFnj/TW0CyWt6lVS8MBiEIZ9IszJlRbxydROGMdIR/zb8K2OVk0rZdreU
zeLmZaiJ3GfozWTkrSK5IqR+eTFjIiRL/dQARnrt/+tbPRY5Be+9X/b5bd0b+TIF
LT9X4p9OlR4s16blkgENRVq1Hpvtph4Yiv9wM63w++1x6x0+SAcPpIyYiH18fwwA
XUg32S8KsmtGiI34+dcTe1BwGP3LsQrWle3ab4u3+SxdKllh4YK0/TEM5WaiaLhy
N5EsboymAgTocmtunT1ZcQmqZU+fi7Jq+vj+IixLQm+VtbtZa7tqzmeogsrMC3Ps
vdvysizRIvZjKya7iQ/9bb7L6reuDbekkp3PcXx6m7ssf7Ns3MB2OfeMViwlp4ex
FHV25ameOgzqyUU5iKm4iiuqer6kkoWxRlnbPr7w0G5IUpOrGSrGHDQ4g/Tibuxn
RoczXYF0SZgjXaxdVbMHWtlRV6ZW8Co3BQbiXra4ONwV3eodvOpJG+JuCr+Lyy+1
HCTnDqFzKgdWJKyvfTRo9rKquSXYkYxKswermyl+EyCvc4KbgJofsSKMQp3RGazC
2h+QhSSHNIjJV+fqf869XA4E0e3wDHRe+vh1zv8dqP1HkrvZKLnTKQaVUZCCL5Wv
EBffjfQdekZVKRfZ+qutu4Wfbj28DTVbFDPzx59KnaMWNFeN57FwpmbqDrbfu9mK
JbvJHQWW3DeAdo2+AXNSmst92cSbpv3WkLfDQ4XKfAhSQj9QqTm8kaDLwA3pumDQ
XmiAHTsQ8ywPoiia7AkrSUN0+D1ng+jiDHg74Pq7i7xbHslBg48G1uAvscng4YJI
6QFe/eskTYN0ddJYne4vmFa51F/4/OjI2MXqij23EMAKF4jX39EGgTCs2Hf7+7Yf
bGNwce5mtm3ukYffhvXuSRhK8F285hqnnbY4FFjIPLOGWMgrVuSAqFpIIkeQBTTB
mAiPnrS6i6dgyn9HYtgc/IllWFpBaNipaBBO9hx7oHxXO6b8ALPKoW4lu9Epm08N
nzw+dVdTHfox0xYOlvlm1jnTOqmowRrAwu269BO4xaZMVWCPOXCqNCTDXwgIw5te
P+Jfni9OVzIYglJVzKs7cRm8IzdxuucA5It4SRSUT66Fiq5i2gJY0ZVgtP4eL+ZN
d6OHS9CyWiVxp5oVm7rgBJ7PjnJO4FJSD8yf4EhA7RenZ6zlO4FJg7z7nDELClhm
mMTR7XY24HC2mUH+tmYXhVVkOMu+SzHqOYU1WrUMIgQG/syvHrDbqsbnnLglZq+I
Ewg9jqf1UgHKWRIxj3OELDa7FMvwAW4MdOUDGjW3+DU76WceQ0VzhoZ1Eyky6c6A
jTUJwk+1AK+JtCbL1K1Tek84v/I+6y+lYDUgtmv2C8hPRTGfoKLCEbTL1r4kJuBo
o9gExXgHDeKElwtFIeWulkZsMyk953OEwnc1w9ITqrQRIQBTgMt3FwI9edWkIRsI
Bd1VhbqS7U0tabJrSgmWzEvLvxVPEhUbN9m09w3vY3vKzy2diJ515Oy5YIdgcdIW
qiI7XoEcH0r+GjVfCGO1L5AlRet/UgkKIr+o7aOCsHeRz5VZccqzw6KSeigaqgTh
pOPzTwLnKUKNcCIvcBRO6I5l18mOz5CLdSfg9S0Oc6vnWyQGV0wRD7YNGkSbPwuA
5vbYR1z9VQ7n5UNkwIZ+KtL4Y6u1TNCgMYzmJkRbqzqWGYQQ9hmSOICpo8XQiTia
2WnjG5OS7FS2aYO1ge8GdqJ5HRYdOjLaQ7jCyXMMEhCKqSr+olIEItsY/6qrDy6O
6ENMWYnt/0yX0tdAscZ4ddgrLLnmgDpT+ZwCz5ZE3E4W7U59QIBpuyFDfTjtSoY5
3KbGrr/Bcbd5LSmU9aXEa6cUmPcOWvgO1bfOWLWgDO07NYIK9J7MHdQ96ls98gtM
o2QOoweUoCn7vmLoji4Nc+KxTTkMUQx7KHwkX28I3ZmZPKCydOUFukwyDy2w0Z63
FLvJcFPWcpYCoebk8EWytcqfhpd6EfvnbFJJ4RBiutyxHkZaib9MFFSitgEFP5+r
yU4UwDRNYXsVth/J9Ytj/SD5ubB8YQ74xBScWgflLid9tdbEC0F2ue5FkydA4i6C
NRJIGnvHr4qRX4vPFYASS4dCvxPeptPBLkNgH6OsmAVIPREy6SHnXeyEl856Xprp
+EzzLoU7AxbBLrcZ9NXPIvjlc/ZUPxhorBZ4SflZy5bym4RJPdO9OOSgGun5ftD9
pGYVC4DqEhmxJEtbcpk3snFv6OFttFtJcZNipP59qWYfYj2Mi0j3AtJHFBrHnSZ5
XueKR8/LsRbK07WCAD8lnzfTogqWlX7dR71FyXBbXgc/gjb1t+N1jihxhAfUQFDE
QuCjL2K8ca6iwV51pR3JbvQ429TWhWmDWxZAZtqL39jjfRnhjomVkdVh9EJRzuN1
A/9eVTP6WfHK6ATg+Enzyk5FBEjsZZvQ1w0Ut7j5JsL8n9Dkn58dDcW87dgDzwDv
0MvqnTuV9JNNVswr5RXx8vX5O+CKuSetYqgxnaFUIS+3fDFr8aipvkIu0De0+O+/
PGkfEgDxyU7yoX/p+kUioSmNEYxoyL0qiIu88KLC71lem3k7giwFHZFdTyj0O3R8
wxp7JiL1FWXu2sSKb3LPX3HNs8tsQUEBRF1hHApkjARwBKXvjxz8CEqB3qf9Z7Uf
s/5X9m0WBnlxn0/FZLdKxW5XAKxPS1vyJX/mdHZosNBHkZnx7cInPLAoRWxSAFHf
FYp2kigXE7qzxYJGJd4S/lfo2AwRe44npvHgAVdS+Iwa+PVtU/YVk1Atcn/a517f
iEBOZrFXvXm8fNAml230rpBdZo5W4BEPKfA4HMEdBIQqYSyLMPOAuHKsO9/KLYjI
yGjqAkrXXE6Mu0XpMGKLT5UCznaFsklc2Du7WJjf43JO36w00UYEzO+XtIDeVi63
n1OycpmBL+NoVnLm10VLFU9+tzr4WolycEUhaz2d3zjhtYN399flcnOWKOehLh34
FCkRXh2R5ax2GJTowranVKxJHYdmIYg5IGat+55bC7a+tzkBGQEBdzO19Luq0GON
zXBsiAETvSsU48unDPYuVDdphqFUGq0yTdj6MmdJoVPRCrMnEdUTVmH0ybDex2PE
1zSboKuLiLgsHQy0Ln2OV6aAVNkfRcIBUAwvuonixheGJd5u+IEGgGQLU/W0VKvt
aJePZN9GicoAQ7neiIKCEnGXnLo+/ooCLqEiNShdxrJhszUl9InkClVJ6XkzAsGs
t8XjoiZeVqeEXEI9EenzsUouQIkSf4fQMq47WFMo0pQkrk2ikZzk2OAIPkN30az0
ckVbeXWP2ovw/ytgkQYUi1cc7XkWWP/VdIIugIoBzzZY4yYj6ClXqDXZgmjWFWpE
hPKHbl8BA4nUTyNkUN8HxzTU/a1wNz1ntICd2lSXx0BA3asFKs2IfKj9YTQeusVK
psvs8JvZlgmnppPMJmK8P2rlGfzzeWdZXZXdsdroliHfUglx565cQsELw1OLy8UC
McsgZYVj38doKf+yaWq4elueP9azH7PDo56+8UGtorlLe1mwcYxkcoA7s/5qnuB5
4YLPkZOBVzhgNgUyVs699C3fYUpXYIxfBbJw1+1It9mG5WXI69Wpmlt5aIaJWU9D
GIeEDR/sJob2BGG3FxaItUUpKkjZcUGJ6lUvGTBfle74b0JdvuaaoiGBevtky1pM
2UOrt+UpsP9262GCkQ6qZ6baHqifPUUOPcOY0EIT1ZAD9ZFqvtXKRHDcb26rfVE0
cfqZnUBK5RFMlNp/nsOaYecWLIde7lhDdKmndcTFS5Nyoxfrr4NUKlcqdOQ8RBLQ
hwA84ynDoVXVd7wq2Ws8+v9zZR1VVwQGFHg65NBa2fWqUnrlBUksMW8z9fWSSE6K
AxezFCd1xa8nkDqRIo/mI6vVM/+j91oTl5Ypu9WxcjNkhNHzli09+tgdZ5R489LN
37fr8e5b062FcSUBGkzwVJYOXybB8ecqhNa64pLFrR9rVv8ktiA3ogUF/SevfHLQ
emGrpK7+ZRU70+UfiCxaXTlHdKqgrSHtqIQXWnzF4IC/EVWRHyluhMxjFaeIfmBB
/TGKdtPdmMvt+yqWVPlI2Bn3k09cNU02FEQVlGnt44oRRuanLVn0IVp4uK//qtFW
JvwOg4Mt9XvRkseeJA/tSBKxg3noAX25wrGJBfmqguZeBYYreXq0XfqF6HKOh1k/
m4uId84zEtJZk+gmqoQ5ctMwoe6guLilIVE4XiUatR6SONEVO7p7o6t4BI9/KEb1
uIyYk703MfMC5qvhTctLdwMSnOaRuKGlfHRAYM7dbQlK5eZVvG6geD5XzdFtOApd
YxseF6G28DBdfGSv+53vguIXeacVo6NtKLXzmQgwBpDsLG2gK+LexnKTaNHA8VVz
eITOmZOVkojrs79wbd4a119czs+M2cckqpb55O3NhNDXIemF7r5/0s6a131pO2vp
YKXwlZiEkpA9duvCFGAZ6mFqG5eMr1tRqQtpmhyiBCU3clE+zjF+WXYY1AiqOtnL
uGlupu9Vja0lEiIUnix4GA00ddcmKFI+rzvEVM3FTFULyHFsnfhCO+2PRRgkzYrU
7bLCywMltWc/7FeI7cNX+AfCD1HJrleYUL3idZPhRrxCyVL3tNaDNMa/ZnTibOe8
ZMLl8mGvZk/uCwrNLvfWIoW/6IGuNcBGkHWsmGiFI1Kd0ylbJv1VVsFP39twwm5n
UW8UQz1xCPWjEWe+PiSaMNd/rFvwofQNwKcBLvD2QA6OLUpkkHPeVvCw1JPqL7br
dRQDEKsmaqQcZ5OOo/K4yC3leYVsFDlGNnsyLQXB31j4zOU2aFQ5aeGRml9r6PD1
tVj6KgVH6t9O4V3Mr8lYHT4sGouc1J01Xw6M3DmDQddUPoQxaNIv23vvz4V0NQ5f
2oxso41ffp63h6HbTkxrOay+jZ6KDgqPZS1GHsxV9HIgmXUx2+kOJCZ0TGx4xsoD
qIpv6SOiSkNf3j+ZunHFL5GhYY10xuxNiRtotvB2Rvp+3Q8VA47sWJvUVoAQpkVF
X9fY+NHrMjm7mBclyCDT2mY3NBWK/bhwJbNRxYzY4hEBaPbwHmmZyzfNIYduSppK
BpvSalND4Qa4Auq/PcCLlbSSc+GWzYWlSpziA4O8aWw9QFcV51gEPEWO4lkYzdqt
BVmpG0tHnT1EOAZJxriKabjo4+PmHfcqoWzJ2kUdywqL9JI0pZlewbbMQs7nNc29
gvDMFSwVTk2rhyEdQlFup8I91OST8sO6LkanlYR27WW88iEnFw5ZLI1myOxUCbFV
IiU4xXbncx1UGCmnhMKzUdIeMLEePWWTyDtPx2sawa6hX2zprzl/OrSVwdhB1fo4
f/v6Qbd6unzgxS7Wc6QoWZZDmSUnWR/kIjl6gZUrWVDdYpbz0GWJXIu51rSLMuY3
MSK6TWEzzFAFimrJY6fAC5YiBDQM9XgJuDaR42dEB7noBvEv9GFkZHQ8BMbw8khz
4QkxhwwAN5MTAzNhWeS4bX7J/u8sJQJ3R1LHiZD2/3BYqZ2qIwvVy1tcyZv4HJ9h
w1Y41WjUVOJeIPb6gu5sOQ9G6eJCtq8mYJWcVikvBqe6j2y9kfpROXvbyAJba3jB
+8tTkAy8tRHyH/1alrZIm7xO9Wsi3sMyPui9S0KzxaOhUVa+SDasSx32DZDhvnci
sbEMllFAJ6jtCSqcjicJT7IP7+lI1+lM+BkeqB3yklM6/zm6RcZGLajBmO4GfwpM
eiiQfKS8H/zSqXnPUZ2/hwMk3JXtT3Twx2Gzf3GqQLSH3BsZlvQZiE2i3DJR2Zxc
mi4hOmyUGi/Ho/6FevRbMIto0fqWn/qKbb+Vd80nW+DNxDeeNkgei0D0qBqGz60X
6W0ImbnGGFKoTVr2zhnTB5KiGjY6s+9cyVb1IyY9UoMeo47knkPYBhwCQcdwsLgN
LU4gq+RPH6PlHTlF8I6OgUEQI8K5Im698a/2OAFFeUX7+k4zlj/4DBzV+WJ7engZ
pVaqPVLqqRaPc7FHr9pyJegU5xgsIvNkDcjiCjsFQjGNr3Ef2BZWqWtf+ureUi2b
qjZhS39k455b+WF+Te5iXhHC7QbOk6hrzthnLfAwTFEBKcIBBvKnB3r3hPWplOpL
9yELRRcxkQvesGWqEO160TM0gxCKykQpiLOhGJQs2M2MRbBluC/ytcD2EyQgRWIQ
eVb4EZqOW4cQhITFUXSpct66vd6ometfYvbWZa30e06miCVg/h8UtnfpXZfnG2OY
/1srKeHUElkVdqgFI8afeP7PkdwH1HsvAoVV4lloctweywpujcKhF2b5zEahTiAq
wXDE8S6srmx976nLv3ouClM/jeKBd8xQt1WxA8a/k2m0FEhaTgOlYU4EBsTUPiVL
539UERRosW9Eti/qRyVU5x/hxCvfRtCPGv8OxMbm1dw+Mvd6Ie3y8eiLC2Bpw8sf
A6t/yLAp0q5vBzxhGyDORPsB64cYLTw5EDUSPA3x7vIAGX72MozaI6kJE/Qi/Vyu
N8IjgKvH9zZoO+rNOE9orcLWAQQI/R1IVdJa6+fY5z4TiP064QZ5XejxFVefkMcV
EbTt9Yzp5tte3Slp6joKTdBgta3E+5NQ3bsOCU2AJYCfKClSOp96deYfOrpbHysB
nKvfqNMqBdaBREeL+Bq7EeoVolTq8m9BTmAP0FyvfgMsKrebvpLTYhE/XThW0MRh
zAzqf1P5PDMeH60x+19nHRztnPFaJ3+S5lHGKSGoCi9+385xQwGdBAVA9neq1tbc
5piVsznQC7U+EKcdYsEgk5zvpdJFTE8LdKDD81+kGtr8TaxcoJn1AXH0AYBEr+kA
DLsoCDcSV24c7jMXX5JBoh12FbMKwFcU97vgeLnJ++JnnFq/I0gFo+VfR8EpjC5k
vKoW1ziyZIuUpTc/tdkI4cKwPZiJh4/Ln6aOQwzUDHBqUVRoRqpBY6ykGlEXnUQs
/j4rqy4MUz16J5xsiL0RTCiuVDn/+wNiCS1MIcYYmViJPiskzUAIki0RZPP40h3G
njdRN95vg2F8KNNbX61gCoOYgaezfWziDZvNH1cPxtVUZj+pP0XxwuK+biQdiEo8
29pz60CPMGOJQNyelX0Dkc6fVkx5uL5nenNXwSF7+boylGmSNxm6ufCkWqHTR1gj
77bC7oDYO7uTKP9MwwHjrpm1XaWYYx+Heqibngcpkx2OBdV870ShMAtN8Hf8Dsnm
47bA8Ie3wDiMn/vdNjlxYErDpdSR1ZIWJZW8y4DPX1aqSE7tLwmlhUWx7q5+JfKj
obuyNvJ7cVQPv2zMANEu+kF5a8MzeG1a4lMWZabk5kN5/jGCtxizE21hXzE8QEQG
twFA/0rBzCok/O6scQQLKvYs752dPd2tz1Lt1GnFogikEufssL3q/3i1D7Rspv58
lqKEhGMdW6+qamtegkSmuFXcbLhCHwNkGC2ymOW8njcAx8Xp6MXW7SwoZc2FJGaw
t4Snr+kJoInXY3WSoIIjkqAPNqwOI31G76U2hETVEYbk8LzcZ3qygttFwVO0Fr1j
S7kVXTGTWgaGjp6owwnCTY+sJZ3GLTQf4k3MlhkLqUzXQUjaImhVire5gsASjKSQ
NW0WHertvZN6Cuzl6cwxy7PZlxULK9fzAVyMXpDWlqRBvZOoujqgN55zFX+kYKSg
OKUXibBpF17xBHdULUeyz4zpqhjiyaESz6jjOuMkrJK41jE3py0kgbbaRSAFaNgX
sRcEVXsKukOVn2XjMRMZ3lLM/BaNmmj8uAjrsGFgxQBAN3jXjQzdwes7IyESIjID
TVmYJZoGswwaKd8e3dpDR/nYY3GkTuSWno+oVJhZW2P28s2QtwAGHfykHF1enRfV
qULcRovMpWmwbXh1MkfCEwEgrvrpGKWyd1xhMGma5yBlsksYmv/p3FFCUQY1Atzr
eHV0u/CK5i2slCHGM9lzLGYvnSasgjIMTBP+BGb7WGuXOXc8uIdUHIK/IupZ0AQB
jvkEzXC71uPK5aOuy6OeNcZp3tGN0aYyyl7GRdnzgugmFs6l0Iw/CY+6SVgvDCq1
mjVQyibUY3IcMg4gPnJTrlngEmOF4H/718lrs/a8j0T2JBNyAXPv3AeBiu/e7gpI
6pbNgikd1njEPMLiqj0HdrQFWji2T0pLVzFpQVIoNapLJ1jjQQgs8IIt9/w5jfl6
skUeaeNVv03aZzD2bcAxMei440K1V3qhOQm0HrPX8LxLfe67q3Mejy9BGPf2Tu8b
ptaPspCWstOW4/KWvcpvy8jReElGTBO2wB/vDyyFAX9OuyS2Y53oR81ml0zDFd7z
jidTFjKBNtQjtIdgybT4vOfAQ6KcMfOGhQqXsdOlxxDkyl/4P7sVBRhEXRri0tdf
VPeX+43ZN53uZ8qudyclzhva4fbg7STT58Ky2vtqLT69/QlLHKLCmmk2tj43P6u7
jFggiVb0ZJcnCAAFK1Fmj6DrizY/P9MqWJnea2qyoB8eGILJRtfOmUV+GmUKBdDN
JqKgLO12CWpEc44mcy2EZgDWOKOeYG5MMV58PZfDK4vM01/H5eOe4XaqMNPjvldC
YoNI56oj00he8Etvbl0YTWYwqOMOpGMmRoe1gDjW93kN02WJruOEaeVEeDxo3wdE
IwIZttF5mnDDoy/bVZHKA48dEFkhCip+FjNaxYQmNkyfHBdm8Ss1Wkp6seB+N83A
T2hlXQPDb7bxRsGey63ZLBp5Rn6udSGgW+sZevSyUfTHyuBxX2Fq2xfmSgquBSZ0
KF6jojKIv6nJjFoNjWskZzUNUkxungsPvz31Ma/xN+EJpnEwncjj6C3RuTdrLobr
HXt6PqxCoTHthM837Ri9+0rFxQcFZDhVhTmKnXCYuiejcf8iBPml/lDkjJ8pebpr
8NSW7PZ4/76Xiq5zXTc7jwrbdPO73FnaFbRzuy1A3eCAiZv8S4Rpw+vN6EAqhVqK
QwKUBAOzp8kqCfZoYHbW/UD86pcPu2hZ21mdZwB+DTmsF+6auUveMfRh59lYgs2Q
OD2UNsHkFdALVtmgicY1VXkN6SS+qSt+IAPExoDotrTz9Bur8hwEWACwOYPhBqPo
RGzJIODEEakxX+XIRVRFA9AoIJYuo291HUGbUTzupLwRMqtGW7ABwiKj5+3uR2+8
V6TD/S2RSLYKH+e58BZQfPJ1zKtZlqFoXdUO2ZWWpqn4bLAC/2g0oFfSjHeq4Rfs
28sI8lEuUgZyKvQTN1AK7Nv2FoLcYG7nmcNfq7Gtb5a4QlCd6aNV5rpkYriBMh0j
jwFBNZj+ITYeDGtVT6Mqp9aBhdrFE5hl8LHjNSwPMzQxi+9kAK6fhZm8EPX5WmBo
5iOYeVqe0upH+ixLA/o28XQN3JdsVWb/3xG41ZEKBi+/l9tl/X1ZK5Mi5n7FebNk
iF+uJOQdVGNQ1BhPJDw53OqCU3DnFWaRbXUDR5WmAHBxuTo4NPv0/T4i90Utx8c+
yQLU8zmE6QTg4SSTziqQE5hWmFhDUOQU6tIWxxv5tzqWUwHGV0lDmU6Q8m+feoMS
rc6mbsqDtHlGmzibBPcQttufrojsi8WJnhe0KgoJrMh2JDTG4XBD3Z5e3SzyirWl
PYTCfJMxR7YPjDGCUQw3D5y3l2n/fSLVSVuAWgw8FiePJVz1TY0SODyx6uyy6FMD
Grwd9h41X5kH8kniH+yty5mNONWhe9dNuywk3VfrKCAm/uaKEyR9L3yauH4BPMn+
AvrPXJ5iIQWuXtqdA44iJvwJAN8SZPHxI/mv2gLWm+yMFIKsfvv4mQSbRSbGsuEQ
t/Waah3RFzTiXLZqYHunwjX78Wp0M3MYtvDP7tISEz6hQJqlTq6RNqkmP+exh3H6
oivnGG4QtbyydTGjJV33Y0mbiDpE2rKu6Bm8Y78PzlWElbRfzn9pczd5tb9xSNFH
ii2hspHJEA4rmeVWehp62WWpnltWil+9SL+gBUcboxDdq7784tVbWiZOVTfGm5qL
2qO2caVsExdtFoze4nulFFQsgJXhezFdRUGGS/6me6GcuVKrNlqUfa4MUl2YUgpR
+ksCprzr4gf8KC1ym94KtA/xNP4XfQhqctpZQJZf2QdCDGKTCFkDGuXzYbQJVqnt
9mE4OZVA5o1aO8HKjN8IcHLmRMkbVCeLdL71Z5REN+vTy23VUUbG/0SCjjOoix12
C/14K4u/vvgAdSa0UaLQEpzn7T8miwjR4EFjwnM0v43sZBESoqhK2WSawRsp23M8
/IlBmFSKFe9GyI5kDqyAMhbJdIUDHZ0oREU/zQBQiFd38gcs6yRnH9hptJQ0SouK
OPX5fIK0uTtNjLwNxt38p9BBklYroqmeNg6yin5821dhIKiOunOfQVTiU/ri67pf
MBlbnzkYbfNiSrbhNVsczMi8mgeqL0oL4cUsPXMPFPV5LARIf6ZNyjsXymLF9qHV
4lKt2z2J98DJlKEaP5q65cqP08WPCBvfd9WFxydtcZGT4aBdJ01cQgQ9qqt3RSq9
xM9x8kpFmPnm59YLzV0/ulH/5jaN+kZ0/TZz5gQqWfOX/pLes9dXY8VcRbPdSU+J
5Qzn0BK0zhN3VfRtyO8H3kQ+MD4nJ88KWjMge7K+CfLJX6dQgvOLsGZwoZmhZqes
3H0o6N+EEUuJRfowBGrgWwd9vSZ4dQo26j/tRjJ9x2K8jNZOzXEpCucAYlBNohkL
npW0EVL6RX1fgXr7v2f1cXpbLGAkGnqKxb9i3JlkelGEsOJRXQY5VJR/f9bP5tg+
VYyteZ0pLbzv5EtELFkKOLvLV1GvG+QtjjoCYQCl3NbslSF0ZheaF+jGQafKIF5G
duDuGOe6EO9PyAXegaSPhM9WhF9ZQMOmhbE1fxAU0Bpr4D5QkBc/BAwWNQa44Ba0
AFhq5N8TxsguJRPlfPdikjMOAaYRw9a7qiaY1u2ZGxj+M8gMLFqY9gCkknpXJIC2
7/wB9ngspcpPGDoNIyThvNrgPI2izk6sAkZ86aNQvs9Wiq0D1s2AtHGFG3i/h18i
dxqcqsVXY9jpqGmQQbm8Zzsoy0ZjmHwzOYOywClPlDwddsDkVePUZHVqIh4LOy6U
TZ3XJqR0Se75X7N696Fkul4VbRWFsikiynLozBJcHgf5Orpd0jDMHHz90hkp47ZF
KRWn6lcsytxLKdD9SlleNYlnV88AumQwWvQ2WIjSDuv7NGNaSmP7+j1aOSqjY4ou
7BqWXSq3LkVSu8TlAsTuoDSKjYFuR0vtzahbnTkbWqvEpaqqqN1ZQDdMX+zrDFuU
jzjWJzjY0ttdvHB154cD9sd5m7UB9eLzYxsxbEQNi5dt60g56NSO5727t0dgcOM1
e7N0lgG8NMfXUkmVExIiYLNnzeqpcReeBW90DQd+qU2lTeZcy7gTnl/kwTW+rWfC
wD4YO79MOOi07n1JW66pv+qqXEtp00NUeH4r/5rjZq/s1dgEi5WTYpFQ/lsoKn+u
pkrG7S0MyUoPZ8yodcIb1CTyafEGxNgmD57goMNeyupKGYJkgnrQRQrkSK58tjhc
65Wyh8QyGaFycajUelPj0F1I94WgZPKZEDFoz+N3K6qGJcc09E8Y6HzGNb7qSAaZ
czhaeR4edPaY9KPjwpkL5BV/7QLuakmHXXO+PhoHnqNb7KIUlNgeNtfdWd+6WWay
1CtG0a+utZ/M3SI7LW3YC4ZI2yOyOxgrv3p6T7hOg6XTXGTdtSqVkWCyJUx2gcBc
ljRFG0HNIxb/kr/sqdcvDnXDHqP9YJWCDqTknn+ije4zv1iSiB9D/sBUksctYt5I
z2OVeKpmsEOTnxQqevHi+nUwzuh5tHDoQIj3hsx3/9dhxmNG6n7pln5UCCLNTgRx
17RXvD5dqRRYFE5d3l4rM7X2WWw8rRVox8hVHxef2kaNYrdCaIcDWq/hvNphgMTV
psnLlQmuzfyd969cU0tkEYLeM8vh/7PY0d2vUVnrw0InssCqEKKhie7WC5EbCC1c
ijvjWIv/ABQXLKgmTRRnE8I/8VjX30P2Xc82DUTsVyKYzp/zZ2DlEytt7t9Fs3ws
JnsgSwhpOo90xd4ZI5nOo1Gb7yih/1UsuAZAFR0Nh9IOvJB4K/S5bZx7C7Ag6G1C
61zfW+DXq285qo5jRWfBzr4IZlr/BoNGdEagqnEfuexOHpZSP3G0JuPW/sJc2GsV
4awFVbW01io+6XD68gOkD+xR2Q1VOKifwW5nS3XzkJLFaK+b/zcav32tWW5GmxK2
RusWOx4tW7Lr4QUuSKDuQXLrc0ywlZxHPJnMKPkqa6pLru9OfkWK2F5aRp3C8yUX
TFRUSbNAzFxQ/QQWCkdWek49Qs6p/qMm4SndyuAZz8HUqykp+WaYt2RiIjztaiUN
Hh0bnXYga+a6XUxQKbhRkaJ92LXImJidQwJoFBTKubt+us/l/y6TGIy+7Yccry5b
5Q6+CeyEkrelfjifzeLsZtVEAgg8TpzdARpE7Wj7lx+lj9gFsm8PEqaXtvvOmMvr
Dd5JYi9mc1bJTsih2N6zgwLLbgl015jkZpSARC+mJkzIKshXiLyg9GVPkWclrOL+
UCquYbaEowPr3jVT5qLf0MrHhBkJUUZcuc/5d/Jr5SR6CeAJVI8pECIlJWKmWPLp
pl2ZQ+yzIgC7JCBmYbEZZG0NhHV0Vu+umJwT3n6UqBffvZ7hSYSwv4qjyeGZGQ2X
OAw7AlsiJpkma7wxrSkiEPXvja66CvgaeXM571YgQ1vwfaqJItumJ6Tlcp8hndb4
hL/voh3M5keCabnbBQBVDp49OtdF9c2otrN2nBq28E1YFhgfG/cKWDF9wE1G8q3U
utWN2+oE3uMjAextV/V3770GdZ87yKf9tn60EUYkJ9atWBWp3fCbHoNnzm0ssiFB
P103dlFRPCatM/NZZY7jQ2Cx5t/NInqPPgpJr1zybwmIGbAX9n4i8oRkLwm1mf1d
5MVSMLAl+a6V/XA8Os0Pb2f/noZzXnfIs79Wfv8yIywecYxJ6be/r0b6+RXw74yK
S0i+zQ5hRqmpHjuk0mAY3iiRNmRKVju626VT13+R9TXobMCIR596ZP7GOKsghmOn
IC1/P1TdlJIzkA3uiuLe8ZW5YaEuv6oEMfUUzz8TEfNK0hg8LKmNDs0S/35F44mT
HJgSO0sNI2eWUmjdLiKdG56rtMJ3vSRelB3cPYIGYZDNkZHDTjpF6/80erCjdhhy
A17ZYZm/YWlVNNhkKvcmhuOO3ncI4TCGFEaAbJmjTs1MXZPAd7jbqHO9vmMFCQGQ
P4WMJZ1h2r/WK89j8/w0tCIpdQcnmzS/sAI6B25iPqDI+Li30wYcZqBb7bHcbYzR
0tqXbP4824tZseDsnlr07Mcly/v0qhk4G9UMsdCmvedBhe5PWbdJM7i1PqwAdyYI
Oaw9MnaujpG8vh+T1yu/+c6kweGBJw31537WWyHMVtjhtUBzfpUgewGVgRZ4kLf6
OtGoATmBZTgN3ZcjbPMn8eYvDCYwrQ4gih1Om1XZiIaPaDh3ef1iMl9bdAQkTKi0
XAoOvVSZ3fq6mE1Mk/fwZU3NGb8AXxlLU3BZvRUQkNM2theaw8HfpjdaKIidXWS9
pd7x1b3o2Z9t1qdNt/6uWZwC1oosIL99usPHv0g8Ny9H1OXAjgbe2GBzN+HpcF8X
9B8wL9Qy/NdEayvzF4V/QVZ5Amu88nIq+YpDRlB+BMcDY0Uq1YpOLKpQRf6B6KbY
8FJg6xHMH2vNZNxIYMFgLFCqAoXOTq4YuEVZHJ1JaMS0Vd8NGCt4HA7wEsWFdi1N
p+LejFyOOVq4EzHmXLLr7LBAOll+PLyPQFF7zU2/N4Z2Uljpm+GJ4azt49AhN+3l
IV1FHP0cqsLiVHjT69h4DHgm/OfJN2GvPEElWRise7APv+AQud1jsHMfGK5z1q/6
mecyLFFnaz14iydF7BLxu6VdJYCqk1z3l/MiFuL+i8j0QDBRF+CsM34nhEt8jCdZ
lt2W4IM6ST32MpQyhaZv3T8AFCF20JA2xvu/J6oIqizQV7y91/5hSNy/WKQb2nNe
3XsRR/LTvlmjnYCvOUBZdpu5xK7yzIQI7jJNtG3+B3eBs8HqOo2eqwqKutKlRhHd
FmuMcfo3dpcY3BD5J14wgWgsIVm93O4SiQoX58dYvU/aKrWxtZdywm1ZjAfTSSXs
cVMUkFnmZVgmjEVHO9+S2XXOk9yaR+bDOrIhla8XdF5TbBJnklcHlJ1rYDELx1VT
e3SoKWcWyKuBYv7qHf1Zp5TgQ5d0Y4eDNP1zp0tdp0geT45GlfwAySifqsNultuh
oFyPe22pTxqjucONrPIK+cXVgpw6HSjesr5QPEeqt9bLwM2fgPI14o7o3gXfH12u
felbrP3g/xssDqkPdoluw3bG/z+xqJH6SuCoylThhst0anOsa/Spnfcu/KGZakml
lcgf05M1tac+6PRWga3tyfupx14f1n3l2J8TsafE5mW3I7bXeSztbUuG2d2Hq3qz
MOO8ga+JKxG+FMwYNTBtprhxfrcyQJQGxYPiSxm2A9hpfUkRrbPFbcQUTCQHrxGy
1IJKIQDwxJC42jgNlbrwfPthAONQIoTPr6I5oDf1pUKhjtp5S47YpTtMOC5h22F5
EP74lh61eatLrcVfzajJK5CqqXZJFKn2n8QMdHyazjuCaR+etNJXq2rdQUcAtI0v
MDl81/IF6wKcUa2syLdBXWbom7UqABbOSbu4jDOK6p7tRzJ9OxxcXE2aOdGiQb6e
s8YHUtH35rwAyeGHnZDIxOIgyk6P5Ue5DD5nNJ1IOKn1hflkjJIImEVLfyQrZ3ph
aqsuU1OwdEPNpXDKYcLc/zLBP+U7nlMGYkG4A+UtP30bXw+5xdDolLK6ap4UtQp+
1X6YAAOAFOrIhOQKagvjhaDTHloF/qzEE5EXR10snqHO87b7RHbhE/vG4+eAdaVz
5p/yTz0YoZT5PcgYK0c/GBTRbLbTsImW3Cb0o5ARuUWginMdcpfGHWp9bO85A/xh
gUGya6Q5+EFyJLzrQFCYnhMOqtCZLI+smkzRICEKtem2FCmtag9cdi9M6007vDjS
0rY7icVAjI9VE998/wcwO2qYnpX6z4P5HweU6gk/6OZWzKw9EGtsSKj0agE+l0Rz
51dAJaJBcY7UzgQ4Qj4yl+erqFvLoDo7qzaoXBD44S3pq2bTrDFLqupF1ZBWO1um
U/7/V6rwC2JGTew7eA/xOpvnix71iYj3IqRr16XVT4C9FER/5k1zTU8pDk7DEdAX
XgD/D+MBp5KaCo4TvaCSThRAQ3Sijkz6zrG/4TVrLnX2ALjMw3G8DyDgQ5U3IVT9
KfNvHmaWgEo0xvP3yi4laKBOI/1GXV/9/FoMONMq9hJId8tVXFles3MeHPn5rCTO
EPYM5IO029BSNz8j2I8/FBDxxcRUrIf0AvRBxOvSlLmbioyWPyaKXesGEBGWbTjJ
N22dZpK4ORmr5evODVObGrRPR7Of5IOoGl3ouYRMjWy4ROF4RXMfzNU7Iim/sDCE
su3B6+9nCNg9xrvHqjf71kmEobbr5ZuGa5eNXTDFTnB4bxJ/ERnUWubWS8xnd75P
DFl8M/XJNl0OUtDFSoUu4I/EtGKFLsbkQmwJHIriN/I3xVf/LiLW2jpxNrgC9zGv
dft6DppZ4+53j2VCOXfCM+ADkBW/noCn5VPtJWGNCA0Frdu2J3Me+gl+u2ZESWQ9
P2vRKTHGu4F7kx62NOSLtkHyO02sHZ0ysAsXa0h1X2s6FxFfUBqXQKkaXIVefMjy
r21B2Vjs9Jfvt5NxOgsMvkpzxEAaqEOVMu6u112+/HsJ+lGJ3UkZwb658SaixK6E
EbKdaxEwxaKAwbb54kfHzn3ZW8MBV+5sfZg6xvfVlBxe6T/fpcsYyFL+cUglm8La
R8qW/iZUoQ6jXCsujqCAoHjIQkYFbok5ZWigT1NZUkphW8N4uzs3nPkveR7J1P+C
DP9ndVfF+L3Fdq//5WkcdNnnQAuy+6NMwIL0kXbDANP+gLcffobi4Nnhy7oNIXU5
My24roGE91JshIZT16yCubzKUNQFcMMqs6jojuQtSPXxqrO78qnxUIIpbC4KmWPx
h4C0s207UBGYQsECI6UoBb11vNla5xAj1yuSUZ0K9Qo3LxvIOAlwxH0AkWU/N0BZ
ZBC1S49vN98a741JS5Pa9rCcq4XoIDii6qaw39stZ7xK5fur/gLaRHIR0kBCEOMY
WxiFmNWgq7h9ODbAREEhWARTV67TvXX1og3hxwqbMUIP+3uaQLmo9Fa7nLxVoiDw
PpfwoEZFNhK8DaHxKc32wclq+VJvErN891LwKWKvTzm/ayyXs7/vgb5wxYpGXoeB
5QhGmnhgWY4dk/lYxZ8r80oZxHbt6vJe5+dhwjdAQk5qvRNyx1qai/WXsEIf3x1S
RLvc0XsqsglFiTyv+pc9q3Q+AYbFQWK6vRvfhzKFgRRJqCCYFKvrh7sLbhs94pdN
5l3xUj7JHA9HwglBhu286Mk5O2r95QsDS/YIDsI8iIC1WwNm7EXdAAJzSc9k94wr
uwyE3MZohxCRId1yi343QHUT2TaQMuKObEX4KWyibnSPzDBeEA+pwIoFPDqg8aiQ
KPF3SiX6R8wU9uXLPZ7UnNz9NaO1R7i2TmkZHPXnsfY+vZgbi2p8BAgjvBHcvtqg
mhSeeLmqmQwxGP5UoTvGyWOjak1eq0stGi09iKn9yydHDUEPGZIUfC5uuq08ALEa
M6CHJVm8xGaueaoEW6EEKlDLAmkxDufaayq+B/DH0noqzGQfOkobzEOdetxIQfu3
Ap2H6grDCQYQ7nZazx3g9UkuRB5PTvEgtrOg0CUZTEJxxLyHeMU9W9YGuUzaMgQb
RvIyF/EXkoZoUrYTjfSwY5oARE/45yXGKcBDtVIsltkWiZQbHCpxGm4jLkqO6yE1
T6j3pO26STX1fLaIPV4uwsV+9voU+rOnAi75rmrDjq0ZUAj8cGUQTjlHaFOUf+0K
+NYXfDFYO9bw52bO+xRZiUobFCEh/bTM+zEsivpZscyJoGb0Z0/mJpgX0KQH5h5W
BNpjNJNkllAarb747Qv/LReCBlI2FWaV/cyEqNOOGTvjFN/k/U49VoatOwm8dGF3
YVphMPIWM6MRWi7jePCHsWXZ5EiGxgVSRCv/VbrhKfEc+3ekoAh1udC5LnjX0o8+
d3t/4kBfT4DDekfgNvYiHzbtw0F15KxJlNCWNHcAIAq3I+sh1HWvRmpN+vpQVuc2
coc+51y3eesL0UG7x7atphDdQ1ZD4OC3KPIIJZ1O+AOpLWBu4vFaSpmqj2pDeQUV
w4y/MnFddsIt2dRp2a/Tej5gQQxcZ1w40i2lqGo50UAHpopKLYYnYuruiJm3Xdoa
3G4Mind6dVmlZPmQzALaN9vm1jgTbrS8k6Pt7udlncj2+A+hn3avC7Dlcwceo2Z9
qN7IhD5c5xxgjfmH3fwcc5Z/QkAt8iCT8Rt2UBHND6gOumCGGDrFnOUHGswtzcOW
6yVmappsTroxIyfmQDFkUcdJie1u9M33qPxfhfotgjfkyRwq8KKYHyEiJGfYwfTA
8AP7+oMdpT4VmqPfnAtIWFKpip9ull1me86NjaE2ejzf+Ww1kWSdc3bJn1jsnf2+
6BxTzMIv2ILvK8fBq2Ju5Rha4gKnotjmyP81xH5MX8FjZE6GqZF0aCW0CO81EpHB
98Zkth/nAWDeeEj7MZaikydDX2t7b+NayRQ646BFSQbzmuc5XItRnTNGZloy9UHZ
vM+y3jBB7RJK05DbmE1zWZmkSRF3lINDm6a+GNsUF+Aa7vALqsGMcHt5CQzHPH5h
X8p4HHSObKX3CdGjtIkAPvDf8DMB/3/VLU13+Gyy1oy1Y9VUr4Fq3sdzD1l7gr8j
0z9l7zot/GylRNag6MT5RGo8E22ImTWxT/xcDIrH0rlyXxvctlB+MycXNh3+gU7e
YiH59waxJZ0JqauyObCg6aDQJAMBD3t+Whefr3qOCmUQwUd5IzFpvWtVu93nEr+m
XCW8Lurm27lxZlvM60831Q9a4aX8oJyEIr/s2X/bgkMiv4q61fgJdJSL8ZMzr8hb
tvuQPBP+S7avkwPBTO3TGmkQrd44ZxOfMJv0G51NRnD0jC7+myueXDEPX3JNKNof
dcCB/45aDJIyDO8zC2NzJRay59fLTLUP+mzi9XCoyMFLQIIqBr9d9uMIjanEMn8V
hPPhirVjM9whNYmyeYtgQm0gC9WQRtD5eTE5Teexnw6Ykl7Ywefg5sF/j+T5JiDB
hOhQC9zYgMwB+yqBTa7njdcuoaRvrRGwoyfuKPSxFnZAIRwQGTe0y2J4zpJTI+L9
Ck4q0LaPSHwnGhW1k0IwlGFHGiTF22iOQyCOXOLx13PBGgnsXQBAOELkg87mNB3O
jpqjVVS53EOuq98sQXYC675cqhohlrtw2LhLa0Phru/fxdks2rSI2Pb/sMDuOcaj
u02FTN5amL7OsqZgSxWiMgMsKOj5eizPdm1d1ldY2Dox9iOE48X8qZmkeu/upbsk
0BDiRwJtIoyjlHH7b7ZI1Ls0A5Z+BwRm76/L9LrMUBgUrReAqVqhQIatBiLWcrzF
oL+Al0RYhqaiFhqQnu7knmyi2qRdtUQ84TkQePoQ6f/0Nvrcr0gZar820D04L7uK
Ifp9M0EVGcEhB2U4k0tpCoRyxUWybgt8qil691gq2sADVIIXboBBQkAuq7lseqGI
Ds4/X7uqCkeS8J5XtAjOmMPvbaZk/+9VSM+40BA/aDFpTCPktnwJ18gsQ3iTKkkC
lalJq+fVy3K80vwNOzazoPEfw3XUYKoGblWVpzd9Naa9qH0R5QOI/zg0HzUNfHTZ
Bd4Zmmi2LCX/DMJdas1z0B6YXUUhOI/D69GqA1lPlVckFt0i2aexPniRRgssSc43
S0MAHPAT/eLOlBN4KBS8lRLmflbi+Fb0UO36pRH+Gc/eJj9x2QBuFK18sHY1GLIh
5WVYQ+woNYVDmSdUtPPFf+y7t4SA1bvz3ascVtAfAtceIz/DRudTqZ2wqbwvC4kR
BWAMGLQTIhV3ouSkxpR4HLwhs4XYrByNL2ztpzUD2mvfUxXFnQkB2M1o+ajXQyAf
sUK2O4XJFbLKMMkzGKS7wt9laP/X+jaSZC8DPwf+7U58bjy1Aadw2L87yGs0wvPp
1kq/dSwd7KlIeWv9xB8sNbbJSWDNiOm615WAZfxdQldDnRJ74TO9TZGXmTKfAiTX
MKxPaoyemHcl/L8fr1GwYppQp24iTOkM9zV1j3Zf3+UjWlnTHxKls/IjacYmWh2r
g2bdPAqAW/NwKcl99PyTSB4A1G/1clS9GNtSlVQvwJOn+B7XWJAU2X4q+njfTfOl
Zsu3vdlBdMeTzPRAWEpFdnrYUQIKMdBbJyWM5a9e9vUzx8aToZREUTuBGGTnSwb6
AtDbd9JHZS2413MeM+XjTTk4/v8wl+qG9jJG6nrQbsNu/E7HtAJL050ME8OxD3oo
AoWDSWwMAZsv46/nrQr4PyJ5aBhz2bvxA5hOStiYUBZqareJiwigwItWmlb7RjeR
SEjC6KjlrPMt7UuJSD37W80cq1BNNUHEC6dkUpXCAcJ+PlbXNIDyOft2q9TfyMlq
CoVxqR1ugVnXgxqo7wbEljW/ChfVCm0tcfytGaGngrnOef/3yTi5jc+5Hr13BYBa
h/O8EbcgW7Nm3B65G1LmghAsgwWL1/i6Jdkpm+/JozWksrQaY/fDHbUQ9PO9PGUG
9LR+OjEDLlarkCprxZu95MDumT5yBQuo/BzeVBxacqreSFGl7rXetxoZBblPDeWR
ROp41mnBxxMnbS+97xJ+XftB8fVySBtTtXVWlB9VQx06Ii1MC1EwIDp6aBhZ5sAb
e6GdnNaSfwa2HNEbSBgJOr3Kon0fPG8HG5FIPpvGE8UPodAeV2gEuhIOOMfX9Nwe
oCugMFoQj2AMM/fxeVW5fMhYh5cGIuBMRYAc1ypG2FQqpAZI/NldcTJoh3PMpQxz
4TaxkFg2e6qBxPrS+6Zw381InW677/rVTYa8fGYEEEVvVTmTZJx1LTvZlRWIzOem
CoFBuJUU3pKGMtk6YnWh1uIcn5l0KBmAT5IhIM8HtWToJXemFQW5d/fMpiAGqXgQ
Ah0OLppESHFM1LhKK36m6yaf4YcSay/4TmJI72N42ze9BC7zCrbChHeoDeJWER9f
1hzmyEIOzPPyWkPP4rVELpZ/v11Utjlfj5ukLtX0RDPoTsgeqsuUurvSigpCBrEw
qWcDy/lGdq3pfOIIoR3zGuwSf80Owo5DPXXM7m+OSjb+aZGzfZaoL3mzWjZ3e+vY
rTYtKq22k62pEK9rsvVvqVlgInDISQntSU5mrO1UAkXo4pwA/zb7wbWdnSvHAvIf
tC1pxd8H6T2CSmjEDI49NYrRJYhNNI57v9OsMgy3EdfV/iaOu5Jezq/fowiqGmMI
o24XgmAqDmsF+G8Zmty/glacjDWIX3Al/CvpWBVm2Gg7JnWpemU90ubmM5aIO3Cy
92m0Xj6RgKmvxQAvQLUZXt8rdayicBBEVdDQ4kpvwlbZ9BxJWaTMbZSu8cbCYjYG
/X69Fi/R3mHq0gsUIecDliv8Fcc7nbHu6xZRfSd0VTIRPZzPc9DytTEbYIlh4IlF
yNZyPs0l4Kjq6RFSq15H6BQq/VvIRaoRJVHKqom0Cl6lD4jv6edZkzP4v5EwsDQJ
aehkwYoDZxt1+5kFePgsJxGpPtKcKwZHyi8RuchVI3E0JUjhqNy/j+7mgZMOgoyU
Ozm/aRxa5syPpkhkaA/PGnmpwUOdpIj9q6gTJOshT+J2mztgbOPts81L5SyYZ/rv
cWCoRRx+KIXiV4UAkTVv6IEyq6dd7Tzsl+yGWLvttZJpDKriHAMRG9gVMuGxOCr4
N1PyFtRoGp0k8eUZxGUsFhUFRdrLCDOdXmJbjkrLo7bhT6s33BzjdMxlHwdpKp6j
F2LcSo5zTcn4NR0fdsrbGVNcC0eH83CK74FPa+DtksHjMXLEZe/28K1AmmKyPTaS
OqbQTE7EsTEw6fKfcAjiizc2GdNcnWBYKwoAp/V2B33jc8KOWgyGJzhvrDxH+F9z
gt1AFEaPkLat384ebeR/tW8qe/jH1aYsZePMOcZA5p4KwZJWKSBwHJ8CKK7rLrRk
9GbmadMMfK56nq+qZprfxdwzjm/kzFLHFNXZ73pjOJBiM9djAYcfLYSF/n9AmLvk
lUmHPfz0QCMU9AtC/yLvXdnbMgk/BLakFEc/8f7ghUW4iwulgK+BTHSFUnwKvsY1
sU5QHeCrMagiVe1nI3jdDjvuJ+NPFX6kO9GleIMIG0dyQM9NI6XDuRI8iR6jLbOg
F693fHu/as/rQMhp75RAL9dJC7q2kc5eGFoWUJ8M4O8SyrCOeGmOV+cJ8Yhq0ODQ
qINcWNP3aySBK4WTwFJT+GBJOkv+aTnjE7Sr5UIo96p9BJ/uHbVdD3O4g0J4+pdt
lf+Lx4OH3a6UTmqw8wQWJEdB7tBTV5DtvDGuizba5KYFKh9NVST2OVaRgxb3jO8q
Qjzis89Q3TqhJdS4cJ9DXkZ0MGIL63N483uwwkuoVncV9ruP958WvvU5CLvTNEMp
A+pXVUHlKLM0aaAs+Vu/dFzsl0HImUDjNGviLFImEWcZsNbmbu9zQko67vhCY+43
MbEJIXCSy8XAIzmFhqCaPCBq0khl7lwiRrLouNP0a7ImrIMkTs85lEyjiT3oAngC
LoVRNSSwzkauLudgsv9zp4d+4KJw1bOPSdLWGZRpXFZzTGbhdXdiTg9VxcoFNXa7
35k9uiXrGWGjME3hwqcBBTb4MLkFZ/lr44qzOkRztVuiClJ7sI0Cmhr+g+WnJUxC
hQhSxCnbYCUjJoI6PbDAi3RYOflS7DcWvqo7RobmZaOCEA9lylCoQQkOxS1H1jUl
OYKzgAzuxzBtvmTt4orbSQaGQaA/qbuOby+KSb4N5r5DqMoYXSJZfC4WqtOB6NsL
p5+YDGUto/84REly9dCV6C+niy4PxF785MDSEhL1bVriscCMYvofHSGJ1Stzskm0
nb1YLLx1qCPV5ovh6v//NG28WF3VlwVuHEWVJSCzQPd5rwCHNSdj1GUwqGY+UfWe
CkRsXW/JN2fyBmqmT7+7k8gzexYy+6zp0xWSp8QAeBGr9YLBO3Z+HepyzlBBk0O7
ylpEkTzbdCD1TmiKs8cO4Jr6gjlFqUzRY/0Fd62zGe7A7N75PvYPQB1l1HSURLv5
f634awYpMb59NLnV5jI6b6hq3lCFqlKGijR/4s/oHiMIBc9Qqx3Dgo8Kz3Jo8+HH
sGjX0BN+mCVsu2EQxFnqp0U5HAgibYaG2tQ9FDJYqd5VKQLQjJtGN5vbi0uVhkU/
WOmRwUBezYmFJLpEWGHi8leKr4x2+a5dxDchZ6pdiV24Bnb3qId7DdA0OBRK6c54
i7HKygxxdlhVLwZo8k/ttiEWv65KMTvxSBB+FqcRqKmCpC5H4eu8KLqzJRc/9mMr
gUn4UKh9EzXnmbtoYzXd2LGqXzl2EDk2DKolwuSM/XEux16LxWeN4G7eVwZzEs5P
epH8sRnjNrIbsnUObbeyaRcD8Rv50j7YY8GNLxeUeVUl4f4NsC3i4OtXH98C72z7
RRegWPjHtV4owe5zYHSaJY2gBcJCzogKewr1S8YzEMeo4i8zS34uF2uHGB05WXum
Y/DeKC5BSXBcxKmTOy85oz2WtHZQJC3jd9nC0OU3VCdW9uLqvAOBeswAe/VZ6Xf/
f3Ssmu4YWHRBWkizlmIEQp6nsyfw6SLCwUoBZmiV9XeOk+cHg03s9gVmWGv6dcaP
EoxcYJWfEz0x4/oUzrOaSfJB17soKCGtqwVQh+xNuhp2J0NSwYy38bPDf7IGZSo8
mHParM7PQs77gexyC1KIxSjX2Uoc5ItjbeJ/669yjGJ9HH2LJYin1xBGVGNiDGuT
qJyLi10eugvv4rueKFtLo0IZXd1XzpVsCPUKVvWHV2dbSHdpd3t5nV9XTGOJ7nDV
UdlkvSCWkS2MP3ek7d/VW28txPizYcYOdijfMNPHF0UTyPr7G0i0t100iT1UONwn
4XTExgky744sF+99kg8X3DBBePQ/6YFDNCMpvlWRmJxOmALwEXp8sYaA9Bsgxn6V
tT7xjUBoMSW+pdLD32hMl52SEn4mMp/Jqna6EWcuHTQ22blXYadK4Pw08BpIf5r4
5cQ/anhBGD5vUNWneUPwuxYXdUQyYupxRa4iXaksO/LWtIA4BuwVu7DSNK1y/Qoi
vDOtZ+E8NkQChhalSwcFYAZe7Nvsk+Ed3C7vUrdyYicAQgizmXnjBAuUtSarhZry
fbZMM3ZzCr6AzvlKrRiGVW2TjcCXLrJQPXwyW/2LHhXJLmc7mlrlr1DLPqeRt+Oi
6FYkz8qNK0fMnaWozGIn99YtHjiDLtTkP+/UlEizkPDXv3b0YzwK2cQiDGWNKceK
rPtfmWhpRGgmlFVnzw7Ys6cZR+W3cidMM2iESHhhCIOxldrOg8kjKOmMhTA+ldlF
GLI05nysLo8p3WU3B3capkG8MESie9pEyoafxD3tfp1dZhbVWEtzV5EvGWmD34Jr
u6DCPU1qMYLtjwPRBOEwoOt65lHBJ15J/tiV3fKpcF7tNKx9JJCDK3CiVNuGVbEg
lOw4jLYmej7GnqPpcKZx+wjh3av6yqCUPiO2eUKaz9+oG/+W9bynWTDhX1ew8fEP
JVFwI3Nejv6gpHOZuUpv7zNBTYsgbY1LUvvE4ZLbziM+f+bHHa2x8owiCMcrR27E
ZGhkkLg1qrx1hTodjpgP7JXAMUVBo/U4dJkaBqXN2he5dxcUoQe/0oSacVRj4SUK
TMbTmMxngTbOBRhw1kSZ59XHO4tM9X+N1lxd5e4Nmi4qUODrSGnJQbMoEvN5X/69
2L0pkiTKa/ZaAKqrr4CVPWilY0IptUETGYWR6U1OYfq3GkGe2FQjHVyBjwbKAU8/
rCa/N/BhcbwXvPH/CBKFLBYqjabSdUge/5hQWQqjqFs/jiAAmnrlXqYCjfdE0JLO
P/m/KMs1xP6rv5yjZj7xS45p9Qw//7WFd5oOyF3nYdaB34PkdDV3rvwRCcTU7ySR
jxC0Oa8qawdmmnBeWn302zQL+sMfr1Yp6wCByGrJoCmMNKKH/ZTBHsYRtkYSKkH2
I1C5q8bHrTKum5BoqR9pIXf0JOtoz2Zjl8rgntxuRbLKaeT2S6XP/jOXc3vyWAc5
ZP6eChJzE8TjkLy6uX0i9bPOJNHQFk8mszKxBh2eVcNvQhrc7HcLfvesXJEpboRG
XCA1nuVAtqhKgpXTS3obECOFBkU8jUqydQs5rH1s/MRqMpCLLC/9i+UF0kje8ROn
xObbGdwzYYY8vdfQIYdBeGjrrNn4xAX1ltY/dqxJmfbv/B/jOZwDWamKvJf0I4IG
pikyo1v4XIRFnKg49/weo2juz0lBbuGRVIkcSHrRRZCTbsX+gKiJRrCLGai0Kabk
BlFxAkzFrjVI8ERxlUecc5w1VCcXzbEk33ZR1EZsMVp9quFZep33Bca16M2VhnWw
YRpnC2pvz+rzTWTlW+HCAkkmo0D0W8Sq7oZGz796szWjiNMqZ/HtPLgSLpy1XBoP
HugnstGUD7ZLrd0WutOMExEGAcPvcEjDLj8egUBn2XFOTn0bUXi71sYYIQi9Emni
8Mxr9USRUFluz1MKSxMYPdOB6a+wFiTLLXMbczkpeKqILLc0JWtqq22UqmMgxhnZ
dzB2z7r3kJQPPwMQbXAV0go+xXKrBCXQ7xB+RLyUGRnKvxkNr4LjhIoK2Jw3nAbj
JnhM4lzV1iFCmUEphQwZzjehjgCNRQdG0kErtgtRIHOwL9+9KaysdHxRUhYvTJs8
liHoCMxOdKCbkuTiwYXvG7elFYwmVwV6/QKhUccu1V264hzLIeWRQQ2a7ICZyuT+
16C+8OlZo4qpjeVj1G/w+KYtNCbQsYG8oANHmdgwrjumZrN8+7QUrubbrKHkoiFn
OX20adnVXc9p9CG9p5XeqTX4c3NP4x2MPEzL+Hwrs5mx+zeoF4xljay5UQlcNNyL
1ut1XefVB5Mn92PzuV2ayDSn9HKHA8LPPkzzRKW9j1lMkMVv6zSL3hwmQ1Jo8+1S
nyAQSZfsM6HdBSiK3Cba4KjOpJ7X8DJMRzEp9Gn7RmJaWxDacQbiV0mlJJVblxL8
0jQ+CSodbXMxIOVy3toqQ5GaQoKrBzIjvgJltfwXuWWVWoi/f7onn5tk9t5xd4FB
buro/D33GHqrk4RwNAt9fP4+3ZbYfQjnEDv/yH8MsdbKKEo1TU50mHsUwXsnoq0G
pggt7H0Ye6BTDRem1VS357d51SZqKrWt48JELA8eom2rHcR8ZTTvY/o9oZUQxHlQ
fOlCmnuguZKd5Nr+IaUJvKwncORV0JkWyFV94ym7pdeinwz8eKXFArZP1oXb3e7g
4L8BDuB55tyMShRNdwee+2QjBKrKvi0ShgqSTCucTwxCr5N/FDdQdCPrQZbFjgu4
lPFDMC2soyVQps7Lapcr4Sf08v0r5tmMjKLp54V/+O95pC5T67ja+ocrMM/kByyg
HHy/QXgbt1f0WpUYKhXruz5osoNoBtmEodQgCkQg5XVPUiLzfaR3+YUhJVprsrNE
3QeF0ieoMj/L6BEaC/6DSyoyEfVLMgMhWTolXCoE4onfZmPNBSThlqgqvzJJFU6m
7Tm3/HxcqXGacDFhxYM42pflMtpNVHsK5iH9OATlKUEzrIB9nSWBlCAFp5gLyzBc
CCi7lclarPbWHFUMDmrHc+13QS6sPlRTZpjaFyhtCGVXoWQ/XX0BpRf83aHurwt7
5JWB2nNF5KSGFa3kWPSd/J+mqtesK26Ksj6WM7+sJC0as7t9rl5CX6XYY/J3X1tl
Bk4iLHDoaYAcZ+bGz0ulO1nID+riWtDO5ca9B/TB+HheF9rocY2SnxEbe9yeHzTQ
717EIBvvC3YY/qnrvBw02YqEHHT7MbPmt6l8VKKELUnbyUcdtSahKX9TcDguqqy+
Yc69wR8snLYqYsZ6OtdNqEmnf5Miycv17ySZnLNmX2YZrRJ5+96m1l3dhW7ep90+
tGt7iMpY2WGC8l/Y3SY2clJxgoFjeWBP+7dGJOMvSic23ShM9u5lSV2euxhL3oVR
mwquoEMDI/FDdvvPKK+9b0GWF+Z6Bi3yvFcVEmoDZbkr8gQhIVg65LvAUURmH24Y
IWixyls6yOaLRLHvlS1Lhq2J6wEWeip7EMi7uiVv/+unlwGVIGfM1n5HMkkvgqfK
DiNkned/51pWiTclohRX1vYC3F4c17Z6eBUAKkQ2WfmDYNW0+JyN+N9p1i+12bRv
S/Olsny75y8zEIlxQAaOQ18TgQGDB8lHYY8oDCOrKmInOll6r84sQpu2JUVU+tf5
50sMccwQWJRSZ7jTJrh5zIH+POAajMmOyh6xuuYpEkGAGFlcGIuolcCMP7BrnTfK
+JanzUMBpoRcq0TCCtaVE5MfjU0GApvTaNCh/Ql3w09W1MtQ8cUwmEVlvALznuJ2
dhJeNIt/55G0lHdSs3JDhGTCVP+9oZunHsngXIQ3ZFfh+sskWlJpxCJeWd7MyZRJ
Grw6nMmi+Ofd8g2I1Rv4iQ6LHbg6EhlAfbTixljy8YceDD4jwdqxy2DFkRWGk2mB
7XY/wi2X5nDHiDiZUHdIEdv0Mm8L38i1Xq+HUas+EgPn5xjN4EjKXtD9gQM5f6kb
UNhabJMbNaB0b9bW/FESreg1FSrn2lT0GcTUI7/qK9Vt0fNxhHJwchw4vOmDxA0f
VvtGex4o5rMNNKzsP+vZMafRSLlxnupYpHFvkZW6asrdXJHbxkhEasfJn3QU+k/z
H43vYX1GYFn3uX9tBVcslqYEHtc32i+X5tZb+K36t2OicdslUbbNDOVu9cA04P7L
lwhb/AvddQlOzbnZXOQj6SxUMz0L94UCY8DBHRAUBWivSilfumupQeEhcMuAHjF0
M9DFbDG/iAD8Kw1u7yMTfU/CHoXuATUDFnzb3y9W8NBUrjwThn3PAYoqynLUrCJj
JWMR2aF8jXgnvgPScYNis6dQg3+Bh6u/3Un2S25jfs/VZssrRWWT1OdCMmMNVFDv
J7BNWwoc6Q2gXWo1PVetAc1eozX74uXUM5fsxcs8mJP0/Qcnt1MRWZAlc5K8dtKn
PGenCVXrpbnGyZcYJD1asfula6XU1xyWfRNseD7Lk4t84fLCKQ8LrM9b8ZgFXSc2
vMHmTN6/XFmB4IxyQfLsa/248n7hHZAVZhvM6RPVTCwMWO+BP9ZBDgcoiyqf6Kiq
renn3QKYSPMYnni2Am+nfdbEousyAVpVzk3NH8B9/c5/dzlzW+3hyjhxhaWyyASD
zuzxlePZB5mtTYZ5gTqM8n8J5HdDue6CvI2sAF4jwGYZhAfXVMFAsmFaUm0r9jt0
FbigB/u36ye389vp5RDQRrmbDu0mDEvYWWg+4YimdBPITFGLagv4000qjQYRhkrT
d6QKHfueGmSPq0Pvc20CX3m6OwN42Lq7meDa8VqwiZmxIKlhUhGrE1BbmDsjYCZv
GNx8qqoXt7iDBVVj+iwxzjS2ObQCx7yUXt1VmicVeywhwMJ5/w3TowPFzkDcxSSB
XQeHAYA0uuYtXAnoKTaxy0lnAQ9BhcRSBTD2HjlH11lu1/IjRUIApsqCwxT1bi2m
kmG5u03ALmzuKIdY1hPadSf2jevtmjc+0lwC/ieaEbXBKJs5cS8tgGxNRsNmQtoi
6JORhIYmhHjfpbTW4QmeycMhViemiDsAGiVaP2R8ohBl1IXYVlgVuQt1sGJdPNLf
N98kLEe23+LIlzawJLHdnQhyerYu+0dKVHXu6Y0wBx0bRfPpEtBT1g2emlbkdPts
MJmFE1xMX5yqIIMR10CD5itrs2qFx7H0bNGJzJxVKJ7BoWG7NIHSXxA6GXIIKEBW
alB4iNlYxlR2JOaa1dPJwOyymI7NG+l77xZJAw4ArQUS2IPbyAcpTR/TuHr3WWm+
Duut3WM1E+V8UqEJKDPxT6S2+bJu7StfyeLo19EF8bLw2vlOwfrtFt2OKDQRWKMN
RlqTfPQBvbov0XhBWEgnrPgcYxeSIAfPTKF5R6sBzCOdZD3ElCmYw3y4j+W+fd8R
TQeuv/5nQ/ki41NVlsyjrQ9OnX+kl96vAnmfMyGpWQXPyvmybXDleXUWrb7EiZ3s
subp92Vx0wY4wUXBHe0XBm4LIe/QLYQrV+IimpdLlWX8c4fnX8ZYugj2Xvz+N4Lm
CkTUqvfxp5vSYCfd49l9RvUIX4JqnlDDOeNkLLpUHuY1hNOXUX+89/RV/X305tSn
HjbJ3d1vyBxHFynV2PXoeQFGxz5NHzQ6f8z3BsnMh1/pIP4uWMVD2czxuxUMrzkY
EwPXm7t11QMazjC+Mxz7U9cz3os3N9HjVu0VAlJrxo+Y6yCBJ7noF4Reh0cbQT9N
cCrwbFjRF09XC0w7mb4eU2G6uh2NIbLUVdfZFbmXRj4II/bpfS8eL7+p0hBlHomm
avacxmT8tSoZLJ84pP3XpzJ15p602jkjlFIcdFAJhxRJwQeYwJmH6HGBy4SR2zvb
2sjpqs7UprqrCXu3WSymKAP8t7R+49GneeUavUmTT18x8ZYP0aVkPhhoeprua5Ll
H87CV1PGXAleY4I9717idISPdy/yNBTnpmDsw1zkyYfP1103E61Oneu8OfLXXsCL
VwpwP+pyif490ufwz6P4PDl378hRm5EUdF658VuDX7JiEgHFzs13uVqpDty1yt5v
dCHgpx4CJgVnQujpoTLnzmdQBJkh0DlM9Yb91CzlocuDth9y6EumpUbYBJDqBLmq
xzabI/xghvsT52WWQrqRdC715E/4Na8SVRhxehA259fvS+A3y4SX1g4Tb8CBwQV8
hLNzTCRgvuz9zg7tVT0uko/rJG6gVAtpMvkAMSm6iBvKUbuMlMNm5IPht1J+iNnx
Ms0nv+jZy8aYxn3sT39b4go1yosKqSRlSZWAwYQ7DiAM5z2NC3rDD6NxbSVA9AX6
I1Oue+SfR/9TivzY+D08vc6cbF3Rc09Q7EF8REAPuA34kL/yQZUIJCe+cKa8UoDk
tIQoEEG3Lr/83Tl1LYMhe6UEIIP/aCO1zrMeI5jRyApbEetD8GfihokTvkdSLQpg
7Ow0FFo03OZVAVhGlz+BBv4PqJ5eM5hRrGoJQwIGp9LVLzjUN2EricysCNWHTKyq
WX3ctrsAiJzjXSxgIW6fLJQZKmgoz5cVA44TFE2d/hxJDcEASzd05bzb/1W2wgNv
b+2u7v9HlFMEsvhxKMFRLavKJPmzQvjhmI+X7i+PxQVrFL3S66+OdonZghGbY/Go
3gL8qiNreTzzLFYCVjPFI1CyTo4hIWs/QvspdCgYMZeGBumAgR0AJVkyUfzxbriQ
2Qp5MBeVEYI5AovZ4y7q/qlN1fLPE3V5AzqWN6r1qQA79zyV3ku3tSzUNBq1J9eG
26p8gxcXJ/cBFC3Z1YXAFLu1TEQqcNA9KxXmXeQf7Z74LZ70MO1zepOuLLGZKd9P
abeT+tCR4VhXnPS4HRid51S8fvGpwoYIJJ3gtPWpvaMPB0IpaNWVoHFHf+6AAQwl
tM6FaoJH3oeF1vwo6Bm5QZIXg6+2aU4X1lTGAqW3opaW3USKfIh4OxDMI9okf3zu
jsssK9rQuvAzIouQE3reLByyAFLVF/8Sfw0r6piZGMBDw8Zte1mPyMuVyaeydM5u
oYNjhXDdNImMehwMdwC7B5/xIhkMdVJ/wmyPdJCFwHMVHNVrLb/1yx0dNR+cRJVO
K+A2C1Mbl1F+ttLqLNB5L7Vh+U1Mr0xQ58sQK0s4MJ8u/vQgMPKn2ME4v0EycMgc
0G91TLYVN3ykl1RrZYcpkpk7f63eWsyCE1NH1sEDLEJ7qaHw4VAyRFMEJBtFvkP4
x1BaerpoqGdBpCih0EIEsQ6i//9WTtFiEZK6JO3I+CDjn/iofz7Dv7y3BrZDfKYA
eE4kMYnVlrXt/o0YsDmjCtUhvRLmg1926Y4vTkc6V+7sy0ArwSkXcnWIHBJ4ieUV
h98MMZUH8mLTBjQfBGJihTKfUoyNoewCvA8xP2jLnsE2dkrj0nIMwBkpxc/pfjzU
Po+PSU4ih2c43vaZvdWwuHpsH7PUPmHjAfxIIM8r7c3Ublsp43Ag8CCvoSbUDaNN
4iKScidGrAWRSLQLKMeCawjGZiB6abnuVZMBJgW0TI3GZLVxL2C4Zpeiv4qTWJW9
ZCsvG254G/VAKHH3aYbbag2f7ppWairfvJuVCTjjljfmv9v4tPorgrUKN0zFAwAR
J+qA/XyGYAQKlMxtng861gikZHpnmlNy16ozJ9+f2tgl0ka1zTJveYurbZ3yMbxl
ytk+LlStsMNMP/29CVb8ymVvQYVaETtlEjj0Rwttpn1i6PzWqhG5xjsQ6WRZdGgm
XkTj8eFu8mcHmASl+3CCJlY4nXOO8or6imUeNubju/BlqsYsVxcHz3qeDCePO07Y
VuqVDyzyPJ767diSf8X5YDoFx5fIIoqK8gCnyz7lVTHc83QdOSZ8/n0CVGdn3BqP
r34Wi3SAuqg1ujx4hXn5442bmaoe33Y7Wk/6rCRZPia0c/Vc4Rla+fHKLVAd/a6E
PKN2LknS4xtvbd4ipaR4VJMT2ZM24kxFusyaohMDtNRmcPLcldb5t4CfZIYg7xU4
iWEJEX6bBZ5WdDbXNebBci6A/Hy8uvYVI1ZMSWljSm5MdZ6u1ATiGYWzlMAoqeVA
cl6tSchCxa9v9QPc3PRr3ueWJ9bhqOB/xH9O7AOAmbaO2dJq8UyiUYdTR85+9Bh8
jE8cE8uDmnKNSry2bnmS4yql5rciK44fPV83R5/TEvfl+JSyzEjE4kf7i9OGDvDd
Ez/H9Q/xuHWI33HNKaZyAtKaNrujXzI4KtaB30eULFnsI3FK7gQLCwxCvsWJpieM
T+xyOW4uoXdThc1Tv6kDNML16eI4RhhI1xTaYBb8+SCnRjN7A65nBDX8Oec2lbU9
hGnNWw8T+JuuojGh3FUculWoYSZabk/pMEhg8JrDt5bCyiMkMofa6KVI+ffN3yCj
Ck6Ch0a5AKoHBTsQUU/ckCfm/wDgw8sogahaJDMfUq74GZqp9cunC49X3zKR7zYF
ZIa7lEUb4SrHFvA9AbXiXxcTKuVuAj/dSkSSmduDri8/UHrg3WIsDR8jZ5upkhqH
cJ/GqyvoQgPFPY8hmkcR+x5rDGNYdl/JMJnFMpi8At0WllgtcWMpthlKFdeyvyCK
1abIE+9UoaeZMMrucaQHf4gjxIj+ykEaJOXhUGqojuBpeN6p3kp2/EyC7HZKjFSj
ZIespB4FDrHyZpFo3oE9RocDlYPD2A2MIqqR4gGsPa53dxEeyRoX0EbDQA9njSY0
Xr7sFvJ9l9vjU+Q258j9Gk6ueRvP2UuJhkGofNTo9p8w3GO3pbqCNP2RjHtVlGPL
03q3qfdDhdqhf3EHB2DInVx8zvyC1i/6hTPWAxdL2MHA5LeiatnMkY4Jz7mgHfHA
2+zOta86OmVzPqUmnzG+itFcE2mHUfwUVkcxIKhe9G31QcTAmjXoyXjPkwQhthzT
MN46CUZMxgJN5pXRYhyk3KYT42zMocYkq9lDmmw2TfeP9FXC9FEhcdpGvfp40ZlM
8wtPNR37DNSa27XQkhDrgoZZ+6NQAY4npCloYYuak8w5Ql9TykwJ63O80KWQjZwE
/rasYDXTVgkdmvD6tocTzl2WehUddCyh+lxy286K3hiGAfC4N/R4atFMG33bqZQy
RWGOGHNFDiaXI1PDyuYzaFFgY+YiyvpVXByUxEKeNpeaQeLrcGYpy0imSCx0R8qq
lV+Mnd3Ol3JRwXfaDbJSoalPSiQT/qLdJ4cMbOWDZueZBeqOohVDXc/UhGYGI72P
10QPrEk3EFAmlZadkeQtSFJq2Wd9b2M2JXTiDJ0WZ4gIWP8/6TYRSSUOGQ5RDju+
9ba3fu8ETLSqOmuypPejdgRaobH3D732hJLxk7pB4xFaK/hga8OpHJnLUCQEvteY
OJSSFVMD5twOMWKvwHsem1xY87Yg1tXGNqIaGox/isURE1QDOgEWkgH0tRbPh8xO
BUnOBxAVmzcHRraboIiDSpnsRbcZOk4pONQyTkPM23mUfth+JFnbUw5U+ffVjlXU
jj+18xSMV5u2/aFhx8Bw5DfmsejZ6ehD0RYXw90RRWEbgWNtMe+MFVChmWNH4y7D
AaA/BA0kdTD2evEk6aYoOBgAtHGYP7aULRXbe1WyVtwpKQ8VgPz+6CTIYKFLp16I
o6WJRJzOxr0SwanIERZ+est16JmlTmoC25OWPGdUl4goOq+DPdJ8xKNE6DUeCa0s
1V7uFSaU06VFDrqqPT0m3h9wACohW4YMUoLXsmPUZ18vXYHdm6mVsmzuCoevER+1
kx4bfjaN0OyLeF0xlsxPIVSlmuvqvgMvx4eRSlvcofY1HV5jJ4QVdy078jjbH7S7
XUKqtEAp8dEBUpahCamIL1AELUgf9Z8LSY60hpvjjHzgc7HWQM7ckL0ywDvzNR6y
vhM8Asfz9NMdpEUVRNikhPRtGkb9BWXXa/z+78ZuAQ8uX0EF6VNdcHUK4AXdn7pi
fh/3A838Vhk/HIGtRzhXOn3qzbDJDcP2r98Q44OhqPS9lAxu0m0ygYI2zVU6KzfC
1X5xijRCxIRvywmWQQBca6uxhI7InZ2s6Bv/viP1ETj4AiieZimeY+1ltUaaZqJ+
U98E8RHLXgy4PolyKzqB1LmoZUmNClF/Bwnk4EdJfrodcPrApM4pEFsD/92SrfsQ
PDKy+PmPyjroSlqmBlKyE5x8Lw+QKm0QZ0vzX/wPIgeHFGAJr0zxkT9jcWrzPhRv
mPzOjpzaNZ+PehTgZTxOzul29X8215f0LXfy6ZwYwWBYplqmyH4ZVZprx+ARcIOs
lLlJ31Mx02RIFZuvaf6cH6od89Bdcgx8EFTLbAPhOiU/FCJzRZ/hOQi+DGu4FTrv
4dOm0JRQQFnTs7L50rvhd+WpcSR0BWsRSFDLYlE4UB4B1Z29pEwm5Vrp23MD9y5F
TRLuK2EJei68rDScQHrnFtPpLUZ6tsokF6ZHZxDJPP/os4Xa8kma1JFmaHzK2/fd
cw5lUPDRebotKbfqjUa5ij0l4yDu15JKrMBTyHs1OF05n1YWtF9w0u/x3h7pPUSD
5v1G9EFUyELG4aH4UVF7ffQpPoPONIJ1xQo66vKoKdBPPJLHILn1l4qx7SkVBcR5
8RGcUOo8Ct+a0SGVs77R1ogz0kJakOLynvgDiosJQOMtQrdUsv8w3btt+bw8vCNd
/d2OAmGY588sXjYRWjUQ32qj+kSMNFY9dVzaJLrvXc+G/jzjCuhDTIfZFajAQBI5
rzblSPYSD8nwTQJnx+bo3w0oU0s7D9G9cb6zVQlO5STWI//FGA2JtXcZdtU/2Qey
qzBcJxrQ1uBd3WzWhmkzTwT55Gk7l8QMrV+1GY0ClAQTvdXWl/HOJCRoszhYLURw
3LvriQseL7vja80GnhK+plIz/JP8DSgCSsjTkCnF/ftLPsKa2T581I/yZeGbpOPd
wcxBpJKqfeCQ1Yxom7coPTrzqx3inW/WQ26gzqRpZLzMU58pC9XEXut2WvsiE/Kw
J2E/+3pHNkLDn/TiruxhQ/dQNwBYuL8ghuBU6KKsqm/TaDAc4UzxTEwoIFf2SPUJ
j3Whzc1lymAQCcCbn3oA0hl5BnMDj+ZViihCbNTSULh/9Q5uM0MjFX+VxcJFc/5W
1auVjSeIXXYngjx6rT5W/crtOzUm6KMZqbNkcqVsuVmSck1qlaKKxi8pqz/Czo/J
oYdAKIDvKJaNWZ2fgaLWPtObwSXup9IUV6OMQAUYSwcaK+uG5h6nUSND6quJ5LxA
qx3djnPkx299XcZH6f5zLbQ8X1eJx/dTjfFY8/n5S59SIeiFgoc6g80Q8GxElWeH
ln8hcGHKAySFyEHcaOu5uZcmLd6eNm+8cNxhoGJoVCv9A+J4Oe742p8QRsqlabuy
nPgVMebP5PIharxtMd6+akidNxkQrEKjMwC2gE1+GP6Min0bnJUt9RXlcLHY7rtQ
wGQxpE1zHziiBbaMLoJIOOuoYEwBSuewCKK1fGMUFY0q2kZ3RF22VBWMcq84dj8W
Gz6MIquhXsPXQyijQu6y6LxhqAEOk9JFsX2ViuYJ5SUOmkIrjs4qKfgv4q3Id4wJ
3hWI2Q3TmozrSq//l+tKwfBAoGxo74e8JJ5A4IJCAcjPpOFlLcesKMo1fbX4UNOi
zJL5zx5MAXRPVOq/TVqykyTb77bUjXyZ8EGm4fG/tkuQQB/n/00MjVxig3m7c5hF
wubI+DZLjx/rsD3VEvvDGfOWUM3NoueAp9lx2LxR5ciqNPedvKs3iszHRpc2egGj
BYColEQtw+e8ICAvrf6WmG1nTtScwDmW3alqk5OB+BDeF+XZlTNLYChUVPbzHO4P
KiEV1dr71L+XSbsY2D9EXBkc8V43Clolq4MlcwLZjJyiTlYTLDyLeNWKUwnTB34a
fWnGgf7tozMLhj584GrS855vUKmWJjAGEfBy7Rqj6CyGHEp8yOGac5IBtspalY9Q
1DyTkneZtnLNtJkbAdN0hhhYogBJoGxTh5hdOwxX1TgzN5qgUlZ2wSfWp05HFCqh
+IKOPFG3QObm03iU5SExJpNffWKB94gE+cINEzdn6VwEnZW3r69+87WDj/jYLDSD
JaKhVc5Q8r7tWiwSe+43eKDjI0EybAIryCMFZjuUI0ghxqMXjC0tL8UNqleETBuj
AOtGNZ75jkJh/CWG6skyLC7bDS4/oSQ2N8cLbCqmfO0W6NcemwjRHadPjv0BPiaH
qOdbhike4uKDKkM4JmPcExYNQhkCz/h/3+HdADwOdIR8iLuqZlWqYTAypcYolWFV
/03SnFGx8M8zk+24eNlgKkdQjHhVeRY42h15BMh9mkqEz8WP3l5ktYe6qrmwSopE
uMK+p58aHWeJII+IFzJq3Z/X3kbYCB9L208gVGnXAuwDbduRhkvXW35s3a7q47jn
9EBjRMq2puIsIq7dgmQHePEtQXHxMBxI2eD4JJpy45cfVMiEG25C9vNObSQsDV5J
UI+a9roW03KyUvZs4yGsctzang54wt7YeTTKgi9NT0ZZonj1ecTYjD9wMhgtcwPg
cHu+Zvy+ICf5Wq8MKuNt9empgiCzTaoJMBDO2cqd4Kgm5IJYmQEZ1Yb0OeETxWzt
8THbAAu3EMZQlVOQhiu9fFuzFebm4d8G94X6aJlRA04pW/MgJZqn/KoXYo2hu5DP
FShGP3V/+fOpH8gb9OHzzxbnmFcgQ/ETfGqX+sW7bZOKV3x2Cj808IpbjTaSnXK+
4LHsmkw3LsnSvZqHh+gGGScjYjK1tOVQoNVXIfyJowLIFusM//v0xLz430y2FU7Z
NiayZ3MfufYfUWggMvAc/bFchWjMmEjhBZWRoyXIH58kqU5R9kWGTdCk6BKLR72z
n9auBv9eRkRhWkurZkwC8pc9jIohFH2cAOXh4PwueHuUTAsdES4oHaL5qtNYgAwq
0UEOfEOOItG0DbpJVBVfdEd6HDxdG4W8t4AAMyLOctKZ+HodqzjYhu4mgYTgo6S7
dTeYe+50y01pt3t39v1Fun38wSMi1MzeJVJtl2KLQvda6FTStrdWJxta4CGcoNF8
0OokcypsZoOw3Cg7RP+o6hJhZA/pI+E6yVgQG6x8Q6tl5vManj1MmL6pSwBVXnFY
kSluc7Urbi3VfLE9ZnVrfWi1wY391OEhJgjLqjDBdsAcNVUrcllimNpT7QnypUKV
qMuj1yO5Mod0N1BXAEo1jCbyO0GCevjGCb7DmfEyGfqxNvbe+F94Wtz1lhFgDZy8
2M98ZTFQGJj+JABdjtit0dM90pC1/x7LVbOgYjxySUaXMCRdB2Z13FSAGYKYP6HL
snaH1zXK4vrR/zJUlZG03gIaiUczKaN/z8K8NoQFhK+vkzVyfEnYxB3/VeBt5frH
Umdgqo4BMQ/wSbFpIv2z++YKTKILD7G8J/E0snBgSkYjUXBN8WNbKeXVNOOzfQnB
WWNOj7xpSgbcEbik3XWYojj92vaTa3qRuKp9twWRl8lIcnpwV5Y2lLqFWVBiqjKN
A+asIk8hursYqLyy0WYQn4gUfLvI8Kklj+SSiZwrjNjevQS1xvXYgzxuPPUmHGvy
`protect END_PROTECTED
