`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
86TkGDb01Y1PGJacU5j+zg7lh3jhMttatjBcNCLPru+7RG8oAShjxdKgnp1N35+g
J1wKzwV2+ROdudi3eTyqTLrPi5lau71DfEhuQKzJAC89ye+Q5ocZhgGM26EqDtDk
Erycpm0ALzliHvzSzDbxqjraS2y7mOG9Bx9I5bti6pV4oAnnZ3cNFWgXPOSM3oNO
9P3pybFE28BwMA1wyi84p+o9NlwnPOv0vwhySA571+gsKhL19NviZ/YvFOq364Y3
MpGJ90Ie8ky1kyTKlAXfm3S5951yvwehLLpGxMPRd8QUfw6wCyjBXPcZk0MU1EOh
NxKT6B6dEm9fgie0amJMFt4gPRNyNrks9irJWtxf6jIzNTQavR+eT0zFtlAZ6SLn
YKg92zoD7MGjja7nKDmGfEnQH92vSQaqVq6CCGT+6AzEPhulryarwBqnn0V7Bmpg
4IqLfLjg/sh6cXmgJVD+h+guklurwAX0/e4wKh3OU0tL20ToyO1Jd6sEdPRzgRQv
y+7z07+1L44y1aREpuixJ/nqb6QIwulPoG+IuhywNel74GbEiG5w9nvBVA0jjKGO
HzsNaDOnHzIlg4pCK9lq8UsvMrtr9XyAi8MJZlxfYRByPigmj9rmnFCYubG7fewl
bt0IeQR1kSaW7PYES16cKthOsXd5vzG7KkurzXaORXDw5BGOZlO5f/pe/RAwN1zd
`protect END_PROTECTED
