`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qf5MJSsc9TlQyhLosmJeaZnhqQxmk8556iia+u52Zm/CICTuDAAuKQMgEVpK4gMp
rM2Vh3dzN8o/QlsS32VZSC3opN8YOFNGNjA/R5/WmzNLFP2Q1lGSs0HeBodHKGlt
VCzyyvikYolDNZxxh1O0J8ZurCE1bzXGETZIdTYI1iNrKP5plHsgNAP2KJ3ON7AA
qjLzDkafTK0KADwFjeAT5FWDAFQXbCvKGNro5gYrpDDf4q4wsMIRNj3n+cR4+lHQ
wvUJ5iTWvC0cxGof9eg1s8ePLGKeVnQMSw4vmJ6vNR3pBGAl1+poeT2ISjp89arj
Qgrj2x8qfMMqEyuhMT85BC1eQEtJHIaqWPzDeMAGs7qHGdJEb6tPJXH7p0Nol5RJ
swpPPkFqi2iQmOmUUqFJfN2zP+c/WbD6+ovl1+CsWKwMTBy2Re4ZLb7mR1qjQohQ
r/8KKGSceDSbU1WvNNP9s0OWzx5cH/LLiiIJCDLCBR2b+X+Zq772Nl14tLPA6dVY
RsWMWV9rcNz9+S6wHzJj0Av0CTZ+pTpsbUQsZTgQjvQ7O0DLzDdo72f9rqMmdegi
eHDch3/WwF/oraGgV9/kHXUGhmaxjFe1c3OEtTSK2hgbopvNq03GsQOspyiRSQiC
8JrtXi0pFnmPaHANpRpGyA==
`protect END_PROTECTED
