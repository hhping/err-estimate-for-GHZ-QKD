`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzWRgLwXTLTh6xTZWUUcaxLqO+g7KbgsA59fLoMV2nKPrmuRpzn/pv6MsKwqu+FR
eCaENptoRhpUWR9VdzAj7bqqiUldZydc2qMOH7Sb6Ng29PqNGU887d5H+QvjSUso
GNtwGpvxyrpkTNk98wnetWyYm7qS0Z1GFn++lrQ0DgsQMSiBrO0lpOSRoEWdM6tz
PlFg7OPw1IUnFeFcv/UYh5hVKFfgFTIqV34nUo9X5ydgak78dcu1/9Te4ecSmAOJ
7vtbFFxXQvDb4f3mh6Iy3CIMtodG8cNDb8Tvqu8Hm+C1nQinLziNBGGTYgz7PhG9
YWPdCZ3WKgRkBgifST0+qfz6SR5oRuAlhktNc9SA5U1Z/7cNz84GZzmvF5q70eTB
OULA7a4wttbWpVj1K8qkyxVctXxhj5DsC5f2o2Pda/EH8RdBesV8vFocn7VOMGAB
LcQRQKaO34NXBQ2v2q1E5yrjiQFop/5AmTX+AZUZQ8AwZrnSiM7Hv2Vvt0RRDJrm
o2Cee6Sv02mpUkTOiPcnCuPM+ovb1AtyHUq9Bb1LwRf0HtsR8YDcvsPlUsUHu36P
Hr8ituKPosoX+TAb/gMojeK0wqnOBPXKQhmfq9y50b7EUkrvNdg53e89keLcLDwj
L/W6n/eekokfiKvSMxfWgsDGT3EpHSodQjCX6mQYsz2QOAcVqew1FkMVhsLrkRlI
xAdER8s20ykXjFuuOPvZB4wjnTBojS+WgNDP/pFlirqKknz/vUuGIrAdNmqSXg61
HV4qw4sCuS1etltuQ1mjdU4fa/+g2Q2XwJLeQ8Lw9tZfrdMJTzsKjmR+Ns41K/G+
lOxTuKobXyZUS0JiOIyBjfF/Zcnbf+LFOgLiFm1gYWsKslqd1vnuSys4RJhL2xsA
vrKJ6vxC3s9xQGG2CSSeFPzGBlQ2s5O4P6UU7tRnghaR7AtOU1bfdhOMFTNSGyhv
odECoQ7qWuOlqfC0ClzxdX2aU/Ka2uUr2LpDx9xs7s/DkSkEis2PjxDqiCKtYuIK
g/gje5KHUsTE8+s9mqeRbj8eM6grsVd4A1lZa7ZzkK9ltG6WS9Ymevs9RBQ8Xvy6
EcZVecGCXopu24ZU23ZDeou1TXZYdiNBVP3b6B3XJhgRdEUZFAPmfx4nbkK86ZDq
`protect END_PROTECTED
