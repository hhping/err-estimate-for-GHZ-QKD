`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4qVi4aI8svJtE5uOZanbnJj4eqT7kddUrj8ZLvzZuj4X4lXtrYJCWeORXahIPTM
W6N4Ku8d+I2PUT+vh9ElRIjz+aFFuva43lmIJliTLsb/bclwId0WosmaDSIPZWrs
goornojLmwWCqq+1WViWZdIP4Tu0INR7gVhiz4PPqk1itw8KC50RoHzH2AsLnU3I
mFwjLPBZREszrqjW9zjtmK/VjPh69Yu2ytVGkjADgVKO6ynCB1bYilvrhtk93dpD
AMDKkTsXnoemHxqfXKdgDpVrykfTqmO21RUn524tAryxCoIq+jSCc5hxPoMJsUfX
4cEzdssbJSQFxUlQL+9YhZy3BMavki1JVnYIir4WAR5UIL+NLNP5lGrAo7VYU/ZQ
zvKS+GcYLmHyHa3RWPmX6ug16lvOjbJoAXZ/WZadU6L/Y+2P13xcFy+YBVN5fP48
oST0l5LsZ8VgpH5NEt/cokbRULIqNEOguguzAPZPuQpfmO3RsbF1kYszC6LXrueW
UcSK/Zqa6673XJiitETQU3Z/I7sutKTkmLl8MFppuM1+yKrfbN96y0ZzHEpFE4va
LTg5PZgLNCy/i/6WrUZChObPQWoHSu2xV3+WnvG35/G9WB0E07yqwJ3Psn500yE0
/weboE6TS0TxqvHHJyfHgaIRCFDnsU47Qvlz29ob01k=
`protect END_PROTECTED
