`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubezxB342wdmiXn9RcSKtLqglG8+j6jOuRSoVhDDtpHDrTbf5EFFaHuRcXXvs53Q
LJ3QQ82C69BgsS9GUCnBoDtZa3tXO32d0u6anzbvpgwDavWSQpI/xlmytLO6cw2u
wFtC2I33r3GqlHLK5HBq3x67n4iAQo3jHSMcDOuYVu3fcIwL+ShjFHEnx3XNlQbv
BW3jZhs004Ahzsen23wtHnAlPkBz8iwLrppJJc2AxiJ87zb4HkuOgSe2NWEatgSe
Dy/mY6ZxLTWhoG4aaSEl5GVe3x4dno/Qlu1+58yEokAiCmkkf3Rk3aW9wH4y5ACT
qKJ6lfPETNxxVHkvHYU6IvqpyDWgEEiiZqeeUsjvZAIf7aCpwhdyfXo2MDzR10jy
XYY2kqsdby0Bz0nWuk88BPZF0HnVH+yY9WaAogDDeY19DQhhYjYmNvZIA/LjC948
wK/dEXR7CFnYhkjEObc8RrDuWeI1IvGJO2k0bUXQJYAH1oma8XTP/brD++OM84CF
yjIBdvvz2fbwZX8U+fu+CzxWp9dywg6L4RDiIy4DWozkbutmo4oKV0398KZPbRaO
Vi/5VkI+X2j+eVL5QWL5FXwCp6HW1EStNnqB/M4o34YbZw6PpjLz1s8/xqi+kQh9
4ofub7NPu4g1hnZ2eMW07LxCdcYwg7qe21sOda6Iivkl3WS8rIiaEwWZ1hxY2Gf9
oYuIggGyfgzPkNlEqWe+P5pXyhGDmIxB/R6rwuX1RgJhyw2dtCvsQAGPh+USlGnZ
qvOKq7RJXSCcaSqPAgZ2Xxxnowu9etXwk1WT+AcxiJ4bVfOoSGA28wQCgVnZ5kPC
PLB+k4DG78XYPghV5P2lRH7jsAEuw0C4O7hfzhB4F1Mtlwj9VVmFS7r3JDFXM+f9
FoSwAWyc7ggtH5KHjndcVDKwkQiWVRiaQjY3DbJO8y5fxqgiPH21tPr1uLryodgw
ZcrUdR178DwgDhHqXaNcj3KPhBUWasYEdSo+sIqAI95/VgkVAk1UZT1QozJXMerU
VKJVAFhsKPFblcqmwnRbAiTzemtC3WHTFY7JhIrErskpcCCiKYkSN1thLFaiOf9O
+RzmmZ6OdLJLQbR5Rys6adgluIfBDjpD0oeJ76dePNCASdBg/9dXCpQhxxK16n49
5BJB1KX1xureKXvNV/3LNC4WfTeN7MphqM7MhqNFk+mY+HKfmNQ8JEo10RFBanMw
yto3nXRr2Tn6yOU4zIrrXSMqdb7SRtqmEwMODySurFSlC+ARKfJkF1KteZ/AWBUj
aFqozZSpQ+ULUZ4uKeZtgBmF8ER8Ws1jypuqcX58lhK3ug1Tu/BR6rmZxZWgR4RB
ecy2gj48uRKR2IQLfRVV7lED0E1AxKmpRXtlZJA71RsEOrJHuT+DsMPYaifPOfUn
2MYXs0PdtvFBYGFSZFEX/3Tn9pq6iGzooR7glBw9daNu6ywf82BXp8MhOvsFRfFw
+D0M5qQt/29pt6A3Qzu2m5jvFCgicjgga0QEOGaCSZM=
`protect END_PROTECTED
