`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+TFSEpmtju4MndQcDUF9m/NfW2jYZRMaXcrbdI326eYDYF31Eo7LRcs+ycmPn9Ct
hULLQeUMDtWBp1QZOaRJGr13r7PvVGWiRF/m8EHNM06t7iQz3X9jBcgNZdRCgdmy
vWH56USKCtcUOADrX+o/Dbf4n48R3Oj78OO7NNEvBtHCrR/QzkXWMN+Dh+h9I65/
hO4fSQ5/F4gqKSXPoISwK1ro42D6OQNK6dXZmVNSnd9/hXm+/n08K7VNsa29sTBn
IaD0Ikg144mNbw4tT5Z10K2jVoTtrvfiQbTCOJe7phOGP2tT2NRLWvS+9a20nbDt
WMwfukklrXmyH0SFh69bgC17W7FfRQKz30boDPs7536AlUOPP7huQPW7OQ8yLWwc
IadAGsAK6C083Y9JjYu6L5QYVvxCeAlxf3Le5hJqpQKPjmAL+noQtTQcDDaJCnJP
kr5jGdJGfxJLY83ipVqlgpvoMrDqhIu5t/DddexW1cZcpHuCoDQ0V1uyIte3mVOI
dVuiLVQN01DaWPh4RXqAn5raCi2u9KJgWqorPPNr6CZT2ySnMnpzjvixMqyklRzO
RT/3KUEstgwB2yNPcGvUMHLL+RappFd8QqeZIARMDTB7ydjCKK0A+USjPyNucAUb
yzlfu+5RawlDF6SaWo5lnFXm6mSS8nUw/rVPepXAQqOMA1ul4ACS3M2vNPF83HEk
RsOrHy/5/frhkCmk+9q5ZpZy7mwhBADfr+nBVfegt8bgy+bWJIZ5WWmngisSPClt
lrjaGQsklCmVxqkaPL/Kt9j9jzAaoURz4y/6e2iYoYWD6n1Y+dP0+6bovCNfeaMw
mpGFSH9qYMrX5uX2MP0ehluxnZuI3V6/i9pyV8JJWfNSFrc3kW5zNLXKCikvS/TT
1KRBWLYrlMvNyibKWxmeAmF61McJOpDGMbleW1V5wKEL0BDjMl72w9A9XO+iesfe
E+snoi0H2HZH1ycRMlYB++y/oarbvUqx58Hs7kcNi6U2nahqgOKTAqJVldzqXdU9
GM/8f3q1IoCAGmgyeOWITUS9G5976sc6okKbLvFPP3w8WJeqUvQ6ALJbxfTE2xwY
`protect END_PROTECTED
