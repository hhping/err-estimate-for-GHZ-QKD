`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RkTBxVemXIjfHxmbQse1bBc8RsknSJ/WJukiOtu0jU6ZlDLn4M+ah7h9DTbHGcrR
kEWMmaFTCTgF35dGi32sQ+CTbSfHrHJvKyrSgfJ9K5QiFJCwjMAK3ixsiK5W86mj
y4AIGC1kc5fHWzub1KVDqNFdiwR3RSMC80c1KzaxpFDLDKFjpVyBXLIGKEVnCmhE
aql1lm0xCsQJm5vAT8cEMRMYdwI77bM35LuukIbFt7I2C4cElc27fFXf5t0bNiz1
wUt7yk15c8L4NLY8509N1nF5zpQbQ89zdyJ/vb+cp+xsCzYDcUmIGmKHMYoKIDwr
9zfDmQHLSgxwuADO8JTjdTvIHH+SEAJS28jB7YfGNsQdVEbH8x8eg+mbD6eyHzmP
4kjyPDuA3rQe2JOQtA+mublsnuLHN5chxBhYpou0DN2SuCmedx2ELN4vjTrg1g2S
NvdjTTvfaTKQ9/bdJ4zlZKlHMLvvo5B6d4o9mfXnTlWyUGesX0eHN1tYdfihMRt8
+HTap1R6sncjq/DCMOP2aMAS/TkPBtnVwYM7XNYNGNBj9tD9YCB5quoFCC4XKhhE
lTvzhSjZK0ooyMEHG2H1rzgr0gWZGNeEW122oq4l7FRPzTVq8VoU01ajxzajc3j0
cyVF5IrvwR8KYd0LvreBccwGj6quxd1z+7vRorxtqXu9xYdejc00addquTUGHGkZ
3Db6j1EcViOCsENjuoPfbd2bJQ6nSo8d1nuUI7mqtcMD9itWdS8cTmZX8b9RguKt
ID/aS8QLHHM40zanPyRWl1qrP0ZQqXX/y4wgG/kdRjyDQHH351ZqAz996zKx+NfU
drB8KKJPUVJkvt3kLje0mng1O8tTo6rSrUoeF8J0Gk/EbpdjHqdsoOsb2uCB/QE4
qFSMmLtqWvrFPaNXEzY1AGEkhK4CrZBgZDXPozSOhs38XwKZ9mnVqUvfUrY0/mCc
YK+6HkGw1BalfZlYgODNBZRZhBQ62THrzleVJ2ky2tbzwdVcatEkzS78iH11elDL
9E1KhvtaHwu+9TXmgSKzz1rxeAyHZSyfGO58cmhI7C5YTBFMJUc2a5rp1veY5eFN
1SA6TYUSibeNyuzX7pYHDgJmuycwTrjP2X/I+JHRtbiRCF/ufAtgfDawZ9HqF4fh
9+fAfs2ugPl2VT7FWzlPC0ps++hjYZxGdTJMRfkUwSam7lGXtho/9CDc5gZsCIxJ
52ygRMLBit8Q/CwsqR3Ur1yXP57RkCObsaDTlgbNg863J7dD7Z4FOy+VuuoY0CgH
ClBCy9ME+CfLnPUkSlFJ7+Ro8BIhg4hQv9LYmAjiMmfZN0AhCwKLjzrQxCeWJ4I1
zjYOtG9KbaCsyW9t+iEbdc1n0yM7W+mhSSHysZgrUrbbNlWCL5KA2Kh9AO+m7/s/
mYgGHY732RQ27r5DBrFyMW7ZzpvQd2LZejyO5jmGEmIRfkLr4XnUDkmV2sRbmYUU
n74fh8cX46yfphq1VF1s5Zcrei0yUMvbcYv78XFuRo+AaHAm59jEO0lm09oYrTUe
FmOJ+JnygenTX1WvcI/CZq3DlMIi8uiY5+BUYeUJ1gxD/iNdLcBI8vc1+q+6JntT
a7RRClUC+VaFAuOnkanLLnAEnftLpqu0Z6sGaX9aG88VEsYdjRxx2r0FyG3XKsCb
zbVRgGq/2QKEJQ8MWDM3YuZasXYD2KCA1M3Q2LNmDVoKwNvBFuORBHC2r8b4P4kp
8/9bx9U6wn5e5LUzS28oBwZ9JevgR2ngtPrA6VEVi/BkMYSqmpA7+echhQseqVWj
`protect END_PROTECTED
