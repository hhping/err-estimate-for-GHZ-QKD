`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/48IXXWqkSQ07AJcvrLyYlAYoVlUYsn9Iysmos16mK1RPlvk1bSGN7sm6JmFG/qH
Cb8+lcUZKAApqcrwjUhWiwFJPd2mkk+dUd7GOeX08w0lhPFb1Xhbq2O4FbFbh9zS
v6z8lJ65+6ZB1riysJH4U5EwriJj16xBH7qhnnXkauTr2auNA7wJsk0ebGEIQYhF
aIilNmC5I0jFwR4MUBr/ZP3XuXtThxSbPMVgydZFVWb3Qf24COxSE3S8wRBjStu4
8/by4+seDETvMEyXc05UljTQDkKFDSt8/kkKMqgd5WkFHYn18TKLIo0KMsjuJwpo
+qfHRMH8fxfVz6yDONPlRisR6k364tSObGeKOJXegL7mJ0w1K3uHbaeWI5rMBhjM
dyJZYRCxOWKOgjTzJ3S25YN4ZzRCmUu6bysnE0Ai6PzRyX9a2vxL5hDwqJlzCXya
uliam/i57k3alNoaJ1evvSu8WGpPmguoo8k6VZ3K7EnO3pUavm9G0Gcj0H5z7uMv
Nq0cWY9UvTg0l5G8qsdwF50FbEzhpVhywoeMy+SKYJom0IE2/0x/+xDszbhU+B19
HB6hTGnAaO0sqq6lP58IzD2DiB6U4FskQGDeen8zQBv+ov1iqfRaZYQqbWygOWmQ
BjvZtbHxdr3qbejE9gPGN8YdmFyKlsYzWIUQSLsxvHl9NviUsp9xvM8vqrj/v68T
7D0oe8BIm7ZlE56GSBVt55FLDlB3p7A3Q2an5aB4CDhaT9LFyw3by1Yojgh7Q1A/
5n5Q1+VQUVf18AJaw/5G7pnVHGt7lwUFzLGRnyyasJYKhXced7qw3ysO3tL5LkxC
QRrdglxuqPFdirwyURAs8tfjoGMbR5XNvFj1MXW5TgkhhUQLFoF6ajRwW8zXpsaX
uWJ7d8CEAa6JVLMIhA5uakFmx+p6zdUMm5EIB1pCp51kSunMihE4ZM7kCZEnMWIa
ct1YSG9WQzLVIrZblRjXUxRkJsCKmP38D1vJJ1gnkZG/4lpXhBrV+ZFjkGRobs8T
`protect END_PROTECTED
