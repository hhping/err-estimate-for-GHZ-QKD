`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcrCcAGMAt7wCA3k2lngw50reZ74YS1kXi40VOZepc39b0537/vo9Q8ImD/BsJyY
h5z38ffaLr0JBeA/0dDbqfbHgJRh+QkXRuy/yp+znpbZScZ/8Onsur/3tciNSur1
8O0LcwMCOqy2VgAD5vlW0IJKRFNd00cgaYM+9z5kYpQcG7Ckc3J1zQxA9IEXAao+
yC+wZQ0Mko18bGGi16OkQt3YV/m7yT1J6MRVkBVcKadWOxsQ11SGd0VHwiPziLUr
TdEBnBmYjVhqBOuKKL2nhjWb4hjH5D8NQu9VaPvGEYYdfiRf2JSSHdDbQmvOqTKi
nrrmQJNCJmvhb+lh4LtLgKdxEvDZQ0uHQ702wmDnjcOYBZp1PbIwsM7/yrD4WOD4
aQruCvPPWIXZcNseLGIPgWCaoNDIo3/uCpQO6RDjD8QjYfAFPRTwc7ZYO738OpHW
q2A2gEevzBkdRYe8IMorxYNRDtiJZvV/Y6fm+dQRlMisdtWpghOFT81X3BQ8+Gdm
dlhpd07Z/Q9SOIhtejQZEZRbjL3nq0g4hlWykFSmLVnVF/rUjhaBYBtuXvI3jbrJ
Pf5+UJrEQ41Wz7XrXr+Dtl1AGOvSj12w0ew+jvxZlF2WTCfWy2N5zBqXP7dejweM
ZoDrUcF8LgEbsyNmnefpSNt8WZRYrL5pXHTrfiHwnOJA+2mFGwNhkhVtMtLTx7GY
VJJX/0aBocVeXEu+XENa6NzkN3kdr6+VZxcMF9fzDX8QS3lvuyspTeVcbja3pfg2
juxFxBCcnwsbGMODI8VjIaih/k/2bKs4v1UQff2ipninSEbiqGfeQB779YLs5baQ
5Bf1NsUKyTkutKP4g5O2NYuy5iYnws2g6xmFZaUhhAIL6BkieByn4a7ZYjD9ZxWs
tDa0kJ/wmJNfJ8TVgymL8Wo0LwOzOguGRdnBeheYYX76ijTOX6j+FKp85I32gnD4
BCIqvdPtIV68UTk7oN73J3ayTq/7bPzDH+jPPg6YFPNdzmMVtFz8+SlThlwb3tUy
wGP7/UgU4jnK5jcSe9THodEWZtmCi+BCR1vbdiDJOZhiw4AFxVg0r4URxD54ptwe
H2WKsYKt/f83MZRGdGacfLAyeAky48KD26X7TUkv8kLwhjRsG0dtlwmUWhqt9iYd
G9YIIPfWekWMWVbbgdGemGxHGJ/MazF3g38IyKDsDWJaTmZx/S0/KsalGZuLcRi6
+k4Rk4fh1YW9/oHjKf4KeRyPrr+XnDC/XOc4zdlE8Jnt2CK8WPJ9Enad4i6w3IjP
e6EZgP07GYh8rVzXTO/r1tXsThqn/9zZHfzolbf30QU/9kdUcecAFcKF0U3HuHUG
y7EH5ODl92ObBoAuQR3BXe07m/HeQtb3VzXrATD0JOSVqtg2sy09TLhNexlKOaOA
0zr7GSQg0CWCdEOgaeveLIzm4jxnR2Ncu7tqjF6cCweTLgHp/+ImNc95T6o9EWms
`protect END_PROTECTED
