`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SgPRyMS4fLNmvqYJR74VljrVGAuRr18xMYHIKIY6p5G/9Cp/vO5JuCVpekBAfaRJ
z8LmjnXdCgUrUvhriH+psWZmDCl1//xU9dg3ZKIMJmRoLvYqNeyJccr0WmOJU0r2
0RCEOjR96bEUjhsDkPCYjA3E2ZBcKid2+eJCu79wP27rTvhcGbewyvYWGsY3Mcmo
pvNlcFssas8IddzJPPLxld1IzAOXF0jVGHdV3ANp/14hC3OfFoJ1pVtz4IfjnTJi
q6hNFHEMhulqdpuAd9NnLsOwSKE1AMoEUhY5CXjeHFSdDH9UUlCi4Spml20GU57i
yLvjUylUKQk2d93nugx5bwgi3GDCQoplrCgvapcoJVq5RjQXSPTfugWOp8xZXMxQ
MRhKCDLCaDLzC3a97ywN6Fy9GChA3fKJHsbYWpS1yOG/NJehqBxzKyzXvZSl55z9
tLbSZGjiihTRzh9veuiD+FKHVr7bzUWJ15pSTFhcKa1Bu5tiOtmDpHnUnGWA/u4o
FOVFAAL01z55MYIC+IRUgm88aKM0vwYNwr8zuUaqImCwajMuQ+IZsKMo4bW31ABG
52Sv5eLWo71uuW0fh4Tlz+/4GKA7AwuxCDD5hv+sJ3o47DIOPAoXfAhcq23jkKjO
yC9LkNWS0i2i7iIqbkUS0SFTNn0cVhLZPEtBh9VNyYQ/QVkQLJHBwM7TQbmhRGcd
Dd4sCydWa0/3ED11zFM88Ce1rBi2MSQhLQE1SsVqkQmg5LZN/3OGXAy9+MmTguHW
cxBplf2UEJPycP4iPes+PQydl5ap21M7viwvVOKREd1cPWSEJe4TPdy1k9iWv9fW
A0XcNzLlxhllRcemUTEp8g==
`protect END_PROTECTED
