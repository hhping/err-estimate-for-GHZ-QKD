`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHJE3SDEOZpXX2CflD8ZznGKZp2mGUgOidwXilK/u6MDYjVbCPaC4MTI0OUoh0s6
KCi+YE+isiEiOP2wNOrvWsR/W8r5Lqckqf5+I1/796xUGpk8TwjoUJf5Lj+mmxlS
mjrBGbMyrKEBQ7rUsO3dc79TFehl/ifchqm/5WBkeO61SjfeXl3g5dzZYgXa3b/h
DBrxJrlsPIgMJ156rF2iFWlHEs04vMx57NC9ybak3kbzcq7u065wn02Quf5RwuKu
w70Wgm7pDUiOSkvKGyF9DzdFPtdCu3zuq/d1jxVElHjNMTUHKDgsbP42Srkhks/I
zxzUkOhnnVnUKYVJQIrer6tUCZms6YZ2qseVoKrJO2N3hOsK2pD9bXfKpBNtw2G4
2DGX7njqUDqM6zm3mjoi/D/CeO/16FF4t4NtcuyonfMCTKIA5ztZlyik1K4Knl32
+KQUr98eBmO4H0S4slaBKtXMmermsxDOZNPhFHtHhCL/hM7kJMfwWGtBpwwqVvfP
+8C9r681moVvsb5SFvZoig45AnAr4cauGVzAapV0gf3GcZuroz0nBV6WJqoJBzGv
R6MIG6ALAX70kRUhmJpiRg==
`protect END_PROTECTED
