`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Kck0q0SA+qxWtK3mEouMAobTNEF2YL4nWiEiLfiBCJkJhyNclwwEd2zXXNGWF7Q
KxQqJ4XLwvVWd/RsOwvURiWeYTIj8dAv/OF5ifAmg2uBTwAwhFS+EYpZ38Xm4J97
ro2V7UdAbuAuxwVTrHhty+Uu2nyoaNSjZ1Gm1j8De4hNOe1BoRAhk4/3HUECCvb6
5FwGqGUMontjMvwr0CRjpEcawj6WwmmEpxqMsCR9wDaAKZKySffAVhyc3nGmWSWV
Qt5D3lCNAdDI++KnKX4yiLlQdXjNG1pNyEXL0Cg9JelcGD5NFzH2uQ98HY3pF9gt
Qvyxqw7es+skXiH6BKGiFoq1SJ77UiJnHdpNxuDnLEgGFoD2ApzjdSWEzrRbJ+hO
HUUzGZz6iTEurCvzIdWUhsinzGrVJx22o2tmWaZYd2ZzbyFWNVFMkdos7CDEgUpP
Vrq+ikJcEMhX5MS0rrkvQ6QPGrrDDi3NRlwzAVy/e4VCJOTZwRRZyVGQVDGCpP+T
57PWzVuNzCf/MfPV58KH3PKefCDQHggtNo5GfXvDiMyElW48cmsyef+TeIiIKHsb
TxZPxltqlaM78/vPbZEv+k/Ed7djqDjXkrR+IIC+CQdCich3TNVqsvXL+7j8xx9s
D2sFLIQVffRKNsDdxbsYqaqGBA4s248ffgOGryuJ2no=
`protect END_PROTECTED
