`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeFIDOIzlECQ0fVLJYSyd/Eg53NiKP2dBemu/wMaosbfXrjA/fYr32+2HaoSayO7
s8LbiIio26XI2Iw8H5RV81pKcizAFlXNosMqnppHRrT1fajwAXqTL6XS1u9wGV88
ExZkISl7AwAlTwHCM6h7rzqPIeGdqOrRF/dyY2HXf2N6v9E7n8e552hSz1AUZKf5
ieZ7QJCMHnDg66MtbsX83sn7MrZkwpum6KXzg9+vjXkyonLA2e97zfCpUlaBrhD7
NiXkWHeCcR7xMXJhl+f20ySIy1cnv31JRT3UpkkyOS4nVbjcEK3MG6XdQfPh3Nst
cHp9AOIWJ5w4Kxp51RerwEkkQ26XWzCzJ1+JBXPk0wQbNAedI6r54er8Y2E05VBb
p0muoJpXyps8OuQxpLo3mSBffIrdEiDO5vIcyDRvn18iu0w9TQ6IcFu2xDDOd44s
bY0H/c2vRYZDfAqNhsrp+ygQOie5keMJQeTyS6tH/lNuSb4X8Ty+Et+HEE0YxwBK
DfnquyDVEYYxmjl6Gn2fnKjRl5p0SfZc7Olx8fOMcl0XIxkONwxUMzhM/Y1siUWY
+p52Si3gix+XmwxCsdU64HN1KnvJzCFqBa9p/tH3XyiEpIVXCFDF3G5dkhAy5sN8
6Gf0GTuP3Cb/ptVPTAIkJgmzQ9+HengprCRhGHBmcTbK39R2vp8yQVhW7/mypSO2
HN07YM5PpjubOytjSzPY5J9RDh7BH3NY8fvp1v3Oe+8xhQFxeoH11V5/SXnU0XPI
2m8PuwwpOrlYwnynvIsFr5dVfqds/nxhEgVSmbtHbeHt8qTM6VF68tSjOOwhtOGe
RDU1fAk/l9kAPE1GRpjU7qQ9K5S6D2mvpy8+lLWOazB4WQhOYl0g6uONcRnmnxrK
lum/HodgsFztuJNr3hO6dx0iyBCz76oTyxJQ53olu1Rc1T1QDv6QrthB3RDG1nU+
K9Y1e5qd4eBVV/i02FIA1oNjauskEft7CNijGAhBHvl7BvTKBJiMWnwym1mR/lRU
dGupJwvrR6TJ5KwzSPzkXPX81GiOtjVaBH70HpWIb6FHE7Jfp6Vh6HrXWkImM8kW
nyYjF0jyHzjzaVBPfCopRd5OUe/55xj3D8TfeyjQZQUiyR9Kt8EpzbjdKmDqsHPj
7JXMkMaWOyRGAEsHgOZGBIMyErRwRWwUp23cQRO2c/nA+UP9OkjBaZK3Bh7QFrYQ
cY8aH1SP2LFeJcSwjMSDz4JOPlV+x2DcJYRRxRIckuqBn1BFqWtM4Ysbg5i0D+AC
ParJ/iMsB25kSZSv2w8P1uhL5aCJTKvFnZvWnTc1gQXj7D0SlunuFfOmFAqjKa7r
Ww4fh3rHY4cRoBqGPuNKvW7JLrBETuAC6MlRt/nfImLDr3FLTi91QdMixATXRHer
fiank/5YMkjId15XM7e2P8M6dCSOx4y+umDfweTJvsYurV/6fE161ODRibz2MXGh
K0SgcC1eljZkshBtjjrNDQaiGwqc5PauFg00BYDGG3UU2a2yrEVsvfjebo27F7oH
ztMAVDe4AD3XciMi4zxHl1S0RhXkfAfJhzsYovVy74wV5T6VXUWlaQ34haDEgB07
MKyvUayP4F6fyfITvfLJta1RO86RB9iISKbh7pAvUULMidRUQcy3m8rnp+jJ9bks
WTJwBXIAhxO4fOyMUTnZRlkvVl8Mhldt8V6jML8fInAZIVgccLi2AIdqbpyeIMA/
TR64ORifaF59Ga5NVN22GmHG3uA47OSikPrdG40AVmmPOW2sYmRaQWWR5NBOeyu4
ZxBGJNrQcRkIG+Ednpk+x5CKfR06RvE9Sy8fK7A90HnUO7Z3CkAYqiwyaeYkUme2
Ubvjlr4tIHwja6dqDxrHwPYGaWeZSu5OIKwXp2Q/9ytQew/7YA5mEAnWGGXopmHF
pkr/aSgsTJ3yzAGYNDCrQC9P+JiHoFrPG9C15yO9d/k9FR+ySeGnAEEAS0BA1C3N
9x8BioU4LzDQVqvGqswsflwmXYu4XUuuCd1HAzBRdUm81ce9uc/X28cMad8A9UG8
cYKIuZ5wcYgPcpng4TpdtR/qrh8e22PIvMCvC9uU24EjKpts9Z16t+06suH16ske
A8Fgb55yScdvyIHLcvGfjd1eJWYTzedhc4yu6qDe9KwvkVXhEmRrBfPfjMneqtp2
naU1HW8Zxde7Usbd9NTwxvRMrCcUeNKFmthm2kEQnJnJPGg1KUUCn2y/6ZTEkvf+
1/goesWDmD2gJVk4Slw+X5EFBfkuM3qR5868cI9kfb9iikB6cHQcP0MEaFCENvpQ
n9kZvg/X4n6hPXcJYRQTnU/z4cHEMP/qOH6yhVETU0xDdygSpgC2nfnVKM/ohJHT
8qR/83EUh0emkRMNMyeC6+5vU3YViva6HpjZNfSauqS+hgCW8nUXtgaPXTsoyE4Q
3Tef+5kebtYwPuPjSzDXc/OJRQNWR0aZM8wLSi8IW67TcAdVnbJAGslhlrhc2BnN
RMb2qzI9jkW2Xfr0wt1Cns5KthtfMlYmzAq1PdJ35h8fBy462nqqqUxsNj2F1Frf
4bCqCzi28YYIyPaeQgrsqFkwa/NM53saH+H8EQUnS9sKZAPLBzQWa/Ml0OqH2BC2
+fJbqFPt6oRWwTo8YKHp5g==
`protect END_PROTECTED
