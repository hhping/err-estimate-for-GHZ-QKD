`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/etEhfttbF0xcob5e49Zx70x4ZusS66Edx84gdOBP8++n/F0pACmCCoUuW6JRnvW
vUzg2wa+G3scHVbYdzNaBXXRzXvux1VKvcl03zfhmkLVaR84Cvl+SsvB9So4Pn6k
znBZrgrX5A7dcSEm/+DllH3GnLeEFQUGcsLuhiwP09HOuZup92azgDixXVzT5I2M
NXPa9DkNHQmWFBddYdsI7LH/Oz73Na/Zs+ohUfhxzD4LtzQMdOVENRpKRAL4HZQz
FigWsJxRlyP8n1BONc/sZKU8uC8ajo2bNaw9lzokIbQ/XBo7D9JIUSRAtx+2uHlb
fsvplsd/NiHBQ8Fc0fN2muN4zHZ1lX7GAkbZbyBZZQ9dbJQ8Gm+e10SE4RVEH0l/
Stge0WMkbMYQkYh5xU1uu9v8vYmJ20eqko0KsS47PQq6R4PsUDyiTgbtVdq0P+iZ
/XYvwtKDmretI2HJTbkcdV3SHeJ8Q75b4xWcDF3BQHS3F2Rc9a39WUQ7zRcbwin0
0YFmJjcBiWE8a9vsXrrO+2gp6krdqUdYEFm38AvXd2r43vPKry+5sIHr7uoLjUee
d4QPnoNqfFWOoHpFlw8wN7rSBL5SWFTbsUuyMszO1xiW2zUOOR5HzA320fx14FmC
TL547XA1HYDg75Pq0v7VEgfXp2VPs0ATlbTob/OpzlJZ0Mg1LBIZ348RNQJwKAqF
Fut7+p+wzF6j0J5eBWNDYy+QXeL8M4ReVjYg2cbYID3HwL9nPmPBVWF8SJROaTno
ykMpY7EFB4sXf9dQkDNTMw==
`protect END_PROTECTED
