`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pZIxVPpPTpblMRJENQkUcB01cnbT+MkVM33ZP3pJUZr44BWa3n+P8H+F2HjVwCKW
w17BtksT41/hWcZJ8gMtJ1AJu6LSndzFIOyTKsqhVmqLkWBGoiWlWtN0YeXlLe9u
7YzmsSoW1b680CpaDzAQ7B+yHa+OKUrDmXyC15L9U0ZLgzGopD6Y6bGCfpiaGgGT
izQymKOEysk6TGykBoHaE2rDQVDPYn9W0YpXAJOCiXUFZdwFrgfBcXxcn4yj2RHd
Xhs8aOyuZjw3MhZ5OgSyjua+cihDWGoYfr5iLapnIuEzP5dpfrMTz92KikGZrpz1
mVTeiXZm17w9U6cRxDG5rthaj+xN968+sL22re0Np6LRkzs0WmAj9+JRRjGhlzy8
fN4UYgLAI76h6RKFj3SZ9VcNNMQnpoY1fmvHteiRCJoXajdpxt9aK25u7cF60m2A
LK2mVCR0fWXfFVq0X4YZivsITAY95LAMepYDwtdqWPKb2WiMXDNtWBN8FKAFJsAY
64NkqBZl5jgTY+glCxUGiH37C0ZlCoLymbvxjOddD7quyfoiCtYFtXml9++jeHB4
`protect END_PROTECTED
