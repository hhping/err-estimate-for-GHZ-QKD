`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkCui0rUE4857V4fXov3K7NKHKl/aH1chCJ6sZPbcbkGuTkYLTMiXQYLd5jwKJ9Z
c8aEdT1KapVu934iKxYXre+XbMmP8IlMiuDwhUoudOw44LtGtL8yOddm0/bwsDsj
jNp61devJhCUDQDlq34UfdbdE0RFu8VOPn5+m9mEcwhJhsa47IPohEruM3YrRWLh
6AVa8q2rFVIqOgpSnyk5LLmTjlnkqbkgdbBERv/snXiL+dfTnEhM+gWV3HQcaRhS
WtVx2/eLPOR1oNFL+4p2t4wflMQzDFttXYxNpFexugYVEa/vp22S86Ix4Urkak3g
uLy1TMl/Kh/k5PU229ppSJVJvETfq9cZ/gXW7Bu+aTKupHWxtSHtLjwNr4a3/nwR
hua4N0Iaqx/qomAXSDGtwM+j2yjPt/2ayoqm1QsK3Os0BbbHB/ytaRb//WXhb3Xw
QkZ+/CwHD0cC4AlZTQXs7kg6kT1dwgvmAnqbOqKuCNB2MvY1el5TjRTK3+AcSit0
5YetBegO8QtT7eH6ZK+0LQ0ju+hYuH4lhvdo0kEwjPccSU3tqIkWWG+CxTKg4TxI
8+It/otq9x/QptgT3NgsZPVE9uPc7EQV1FanbA7sG+Xw46VilyiV3TBqUO7OUo2B
OKRq0H+WW8YfabEU1QMorBhgKWW0bA/Vk+oZg97DZgsaVhR8w/cry+nQH24vIo//
yZ3GHR5eQafeQi05zAikVtUFH8eQIjv5YPnkZ7Wll4cgA0GHyGItigg/4sZM7nyT
2Pa8cDdB8i0RcNREMtN2TTpJwxqOOugctOQHQfok+6xdrPz0TJMccq7Wrtkh2pt1
HvtgKLeN7UC7HP7AS5OC7qBWuBIhF6Lg0pvgR7KxWzbFR+KJBxZ+l6oAw2EPgHii
v6dlcnx72BbqWyx+K1D5v1L1wOANt2Cn9Um4NaYTgA2EVHLFoS98aL0g8kZ9koQS
UvIztdD6P3v8ecFFC/2CsRwVcCEVPEHQCezvUF4leTgLK4SD337pP2MJVIZIW4Ug
PHsQGdW3qV3jjJ/29sjceFjRNWCFR1jyQEkbqGS37i9oKPR9QHw9x7YU56nNGT0Y
2ox4ID5fZOMmnkAQB5x7TVvVIuKGt3XF1wEwQYXDt5ezjT2svh9fciHm4AqqnEho
59OuWyRK4ok9GGtAX/lktQ==
`protect END_PROTECTED
