`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4vykDZsIfuZlNnGDDqbdPSIZme73ovcT6hoByHfIkq5gjConSbaPgBAX82LBXtm
ZhPgBnMhBVLNSamEK+l2QrKF2/8fOze87l7wjpE7X8vCwUY2XQ5kk3v5enSRGP7/
O4pAtApl4aEcSw8WWSlOY9EVbxaVVUIZ+0UXxUZ/7IArhdFZMiddv/2/RX0wKm94
K4WpHH55KoS1nG9KTutK8RSWF4Vt0r/KGzAZ1w7Ph5dmbHriqBzjQ5PQteaPJP9V
Au0DMFRyNeqHyUd0KplfJSQVrejiBnL46NqXY+n8Wr+Xsdjg2yRV5n9wlsCLBr+T
gbc8Zpf/pOyWInpJ1cZYNj1ZY5ozL/WJHXvqDrCl7zqs0k8NXIHAm3vvapv7xcLS
J4GJxuMiTiRUfPp3TGyxInDLjFvpl7SR9WaruiutgmxqyzAa3dlNH/KvyuEP2/Xu
lWU0Jusqg4par72DPFPTbSyQ1Wg9BHvNFDCp7czWC9IB+XN8KFqm9MMMOUJjIxGj
htl5iC9+FQG9G3uKbu7uJKKJbyAbvNUSm8TQq46tf1TAqQRykW9+zMqCM3Qr4H+x
Mts24UZ6hjNDIA6I/g5SfBmNT6AbYZOcbSfaigmv0Cc9StY25o8nKllPYKeRw2pT
8f7U3IhSwbe6bdwhcHQ1NvVYHF7O5v4ojBWWz1+Oxqrf+sEi0GI+JImOQ1Vb+Y+6
KGjgV0AWTMudVTMJgYrzKqg6pkwvlZhimkkmuS8KZDrfnVwEq8of6QVemsQCL/Nr
kUYcoCR89ol62vHEZVWqjW6ysIplk7LEhrk/kzNf7DgJWSzxDaiqVG2TYt56WEdT
EFiqHo49itRZ7dwd9LGjo/8UnPjIgb8IbTch0+f8BqJe+DMvnjC31ZB2F89Tu4dY
p7ZGqhO3kKY/VvHW8KhDNT6OURadYtwaCMP973OB5lO0q2a6Qa6aPbt9sRYdvBYq
/aOmYkoZGVxcfjm0d1zPB/3CeENw2C+rU8dIs+ZVXy8a6YlAnM7BHbx/mJapDkGN
sr0t6UgQw2WidZowikzvQKoObJLVaQrGWpmznrjtlSoO4dvbcGpRwjEBHrBt0uo2
0QFO/z+rPaN1HJTrsTmCasvGQfMdQ5kigfNpNOMljuHgGx7ie5AsQ5HLgvAfYs3J
eIkCJSfs/QZsKs03kW4AIRmROAMTiSL+JHtysTGa6sQ4cVp/bV7dmVNJ1SgHkRcA
vtP+JuygEHFVK22PFasip8xvd9WpmvxonaFUiQwWzAfQIF99mDYtlqSI5wCQZcdv
tXdeNCPUnfVULGA9YtoIII6Wb1QJ0s6zisMXN20dc+HauHbL1qsRozq5SitIlCz7
Id7P1xntrFmS22yHGZOhx9ZB8oBS3hub1a7FwB6kymePi1nep1TpWsg0rXzm1VlB
Bk8KyLfnHnAyaFV3jsDiUsvYXj/OX1UickT5ki6r73GhCPsGCPrOowq7/jRK7/aq
QgKSD7vEgN/VmkRGSomRCHTAqZr/J249MzafGqh85eTgI8By3R3ZF/xIvh4gzo7m
1SFK87WrPogYEp9HEehF468Kbt1sevGBcUKoe9/vH+CsHL2kmorf5IQZIsUfFACG
tvup6z/mCbS5JMScioesUgH/LGmVoufFMkqZZf0P2oxMoKRnWE1YqUOyA8mr6ias
WGlxaEeW8mMeosBTxPmqbaoGizQ5/XPXnPQlRYmqWVOnrbUmU60++zKTJw0vcZN6
bPV0Sg7L8b4h22TyKAbWr41uOjXTA9yzFQZkKrlbI+RiZWQ204ahRzWQ+FZqHXKq
5u2Km7I+UhfXL+jCLVlUjd+D+fUnmx0Z5lO8odwuESVMf3IXsfwvj1m4B7GLbNVF
RUiH3QfJTeg/LMvnRNNo5UyPS3UFgFnw0p+BY72BsEZx9w0MvZb3qnIdQ1/C1DMf
nHEnJ75hlrPbGNfjZ3ro6j/qoeNZl9mrycF9vOlxVbgxZ6Cpw3pyRvnIgZBtdBy3
YkeEIAxQ3/vvSCiD1ai8N1gPYlX5KlDy43qvjGIlcJtG3rQ0UlMpgB0ct/0D8E7l
rhONWeEBgMDqLMzIM05sM07n79yMRrdp9tissqJzN7HkqXp/JAM2y+uvxcg4ITub
ZfDN/+pNOMfoo2nRRJklQQ==
`protect END_PROTECTED
