`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZgZVwJUoAkeYEQqql+d3ZSE5oBhEAcKjC3VbmB960hOAYwsLbgL3wsUCxXmm9yu
8FmdKfSlRsdm6YGei/+HMYoAyqi9q452dLu4apPjbW4HU8JTBWwVu585IGXLnB7V
baPxC01OU6NdC5wXHN2M4VmNIloIlZf2qvpWXNfBJK+Nqvq5ExiJcsJN6lnRfmcW
XTwsyrCIkwlNdRpU8wCtw0NAqqHmqU4IcnTlIvr7J4IWohbBe5vsveoJPDYxnSVy
zqsEwjYFx/Wdyld2UtbOWm1wYLaf7o+jmOs5tWSQ7LeMK7AUPmYvbQCvkxcLIBqy
pRGuVrSKT4asXePF21+RkPnMVTAbU5e2KB1PaD1COFQ6ooBCB/CsIeWW6EXT9lsQ
/xfamhHjH9+8N9aGrch+MLI39wAPUf/pRbO24+Qv6fdCgj9l2hYF/OtszTjc7I/U
Zkg5yGNWYBI4Knmmly6k/sKsiOeeqkmv/UjeBM11ttZEeXOB5cfpDQzsKcxRVx+S
fxDxgBMk+FtomU89cKZRHYgAuH+KPO93T/cZweFeuqQfii3s5vIwWSU5nW+kSNjS
QIK3Kaug2b+b5Q14QenBfVRJKC6BCIyBq3nyZV13c3m4aMBul0+jQnbTiSOKWy1m
Q30kkXar0TuRmj7uFqXFsaGWPxWTa1CIwmgjV1o/5OdN1AJ1GKBZVfjT1dUvhw8D
Qh1Ppv8LV1BReKZg0limWUIypCskb7jnkmbPM3q7nYmUvM596vpwwmrVyg3UdS+4
FfKaPTaFWjNSUB/Co/epKwsWw4WNn6JIF6VGbTncszeURvUKBZkFSDg8Oc7Yqvy5
HBicnx0sVf205fzek+pz0lhZkxpbK2JCJTezj5hh/BtIRzfnqpM5j0bYRPi7Hg9I
MJTo1AJjHUCZ1Koa26p2G10jg/mVQrPjEUPUTmKZo+vKy3CpoF5+TReYefVKejzv
oN1IDySSEE8x4XnZdytTYedwa42h05FRUHZIMyzPaakz5L3GPG4j/QgjhzoZTs2I
47bypvv/cfJnB2YpsYnk3glTjG4CTXKKPL3lfShNhc3tWgS6zFCB54r+AO7P2+6I
QMPxbL6dn7ZPi0jPCDQ1FwR1Zld/jEsKr72UKGYBeoSS9+QbUQJiiiXRXthdSCgc
aVfCAxAWF67AVfxpRpYHz58SxdJa6s58O7iuTZ+/lMhrMjReImvYEQxE68lRfj58
hRMm1sMYPHrs9ih3GQ9zsJGia6TcCtqvQ9AhBUtCd98qqgG/apjfd2u1q9GHR9Tz
cxJ/1bOT0Rv28Lqup0Ww+hE2RcWT2kfFKl3gsXn+nSRGH82u4BO9kM2dyrZKfASj
evAzY7FYJIQrHZI3af0+W0z5Hsz5HJSdB9+zHMEvRM5gvG3j6AKQkJXvvP4kK6gu
OBfLq1So/G5ird86WLMFB/m39oEZEKB3edoHXBNX0lTh/G/VtE1CqDBFYFpcxUbU
S++tSbaskrfM8684jYCQWtFG7ojl3Wf6oetBqPgFhtjGXqKk9zcrQk2TO2Hx0MN3
DhrDOQkF2EJt6mk8Mn6JntV9umaoeE/BSppSKDlQ1Ay1oHlvYb8yihBsRG9Om4pD
09m7mNcslVCFp42JyHpGyFGixjaLCI/VCu8p6yVQeW8RmwbSsx9Z/svWpOMz9DrY
kmRNqmX78bowLRKzyqAKvHSjmpOsMb97EqUdYAXPn+PkMOr2uUNbS0Wph6JRdEQ/
NaH+RasntGxD9ahjlS5r8Rcfe3xgoA29qWT7EESjWDHj6jSv/CnX+PPZVR0ZiLAk
+Kz090wSma6lVfsf6VhBmCbpA8dh5JxOIo0khbOJzy8uit13gAliK5m6sVSSphnD
uVC5IK2AUUH78QZxcRAxx7vipRILD6+721vk5eF9xeFJVyVD2x30bpwAZkTwFTSQ
2VJZJciT/GG3trYBjrAf4XhgYgHdl/Kpi6EcCt1DCKFLkvyRhl1mTnbKrc319LsK
MRNupBzi+4m6/z8jPm31ZI14szypyoXd8j1vtI2KyGmYdkU21CG27UQHV7HzXPgP
m/4C5s2gjDETg0ThWp9xCht4nwNgKH49FH+oUq09J5+qKITYIBwLXSgphp4N/bfE
MxGgYYo2NOLeiF4uZy71XPq4p4w2Q6SH6YsD5kqhOhuTSzTtwcLAPBZF+Ra0PhTq
b1UfDUPgmlewGrnHxP605f1iXRoXbl1UoG6ZasuajX89X9v2Kb9TDLHxFGJ6JI04
2TCpXrUqlbUzrHWb6P0xihfJLPr0NxAFEsGOd14QvV9KfrzM1RXv5RmNABjZEka5
yw/zs9JzZ9XPtG+XlbCK18mGDR2F1kSMrRyeFvsHRyHXAISXcrgo2Yf3qIT4l5Xi
T+haqPd/zFBn82CBHGF8RA5ApYqRB7xVONAQjYu/HZCZV6iJGiTc55u1UHFLF4rP
raQcDcs9CBUkwCpdNnfZNkotjOfnkSLqEIer9FP5FOluiEm16WblmMLv1fJfrRFR
XHChiZwf1sJlv/+ca34lJB7sBhC010A8T+nagIVzRz5hOAyUxzZAHCIX7dC8bO4j
qQOU9fgfbLRpVdxty9hzuTjZQKyzix7b1txxfUk/F2ux/7TWZ17uIRuBmISkX6p9
yL1irgnw6u2vZW2Hwy4gbYq8nzKYU14V/uw393G2uLtS+VxEXMxrjrvWUeGow5d9
JGDiIWSIF5plKqzqU6JFuJlF/BqP8xNwpyKN8tKzvY5ODti+XszNh+yxtD5K0Njq
RH8MkWFv8A3Tr3RbrN6RDSdQ8+6Voqw+BTAqV0Kn2gjBIqLKol7vHm2/M5vYCIGX
Om4zp/vBrxeHgne6KHsxTzJbgSarne1Si81XZl6zPXBwtFhbwaDOhvpW2+gwrK3v
N5S08+cVwyGRHcIE0B4NviwbR9wPsw/zUPW5nvfRAfiwkj0xyNzMSVW04Os6bdJw
YdwvGWxf6mDPUSpvE0nAprmRfyaoN8+URm0Hx8rmxonCjDD6Bfyk8VNUGTR0v4ui
1yiZhYWyXufEVSAWH8p6IHXjWkJCRoY5MWg/uO/nLluqXKBgBaClTYxaeGn8lM/n
24ybVwSLLjvf0h7kqL+DsdahGriI6bCTCbQ7+/YhzrSp+99s2D0U+6uePaaJWBv1
9LJl63qFwRhBiMdw3EGWJvkMFWIi/mzjwPSpFR481+q/bO0xlTA6WZ1EfZbtPw5h
Zc5cbnqnv/Qel5KWeBVLtA==
`protect END_PROTECTED
