`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPPcAWQ/MVp5J67zsNZp0vRFY2AhbVmXta44zz2JYBiU+M67B/76Sj483RHsnE24
MdtcEi9jKBDRNvelH214cmUl3qOjzz8kpjo5nqBPEpRhw0Iu0oRueIQVoHPEuZoG
5seDggsMDt0JFkl2dGMIhJtt1QLgtk/gWPjN/khx/rzwYPdCG2bDF5QrFISD1xta
wfXiJwL6HK74RcfnDYLDUxvZMrigoPEovtmCEQ2t2+eDMoP9yhu05djp2KxFdMHP
OMQbxc2vhm0OnU0Un0J6uVryOQd2BZVbVGOqyjnfLkPdmtB81taha7IkyQf4Hx3+
S7QLFwEhNfQ03on1Yyq9G1I9lkMZh/DMcfFj6wAZwKn9Q905OdCIubjO+l1FXqqM
uwMT4BwPI4FkwCq/Y0k9gw==
`protect END_PROTECTED
