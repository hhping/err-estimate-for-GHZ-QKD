`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHNBEuyeSAbhtXS4AO6wHBsDP1gK8/tPL3D4bXZ7D4fQw960DjpXeJ2LWapVRLKY
y8UPAfApxJdLDLAZbkWIEsypGkuYmst6SaDaxEkc8UpNiCv/xAPgpkBIjmwo2Fme
7maY6CCgTU8GwH7HwQTcSaD8TcL5ytC4HWUdguc9x2i+fjdNUynXna0s1Bv3xHM+
aS6SyWTEravCdlFzh3I/6HIJGYahnXkRBAsPMzjxu9+Vq2W/Of7BH+s0vTlJjI1c
4Fy2h1OlvkbYTEIORcRxJGXGi9oxXOz2PBReBjD1aWNEw41OhRf29OUADEKkC4iI
oV7IuaZSHzIEQf6zCUKyREWcq7/147HZNhbHluv2rLnZTBteisqmbG7Wx4iWJYwN
83CWkSSKUjQV5ZyrwO5lTioU3yOpcfexPrP7DlvNv//2AO/bssk1tw3PjlP0ClRe
lAEL120n04FUd4UNAWIh1RHrINffZ1o2EWb4OZII3OELihzVqh7xmxlMGu4FClh8
hCMiqZSbqSomAyNsDPtTAad/YpshapM1FjeEOigNVOnOV3E4MM4i0fuB00BM7qNS
CQ5/FBTM6GJouMPb3HZCqxNkv9ob8txyYAIKdqsJk0K7wTymfWHZjMAmkNexhgQb
uaWKuxJeMp09TijMgrjBjM55E6DvlnVfm/Z120SL+qLOrRDJ3ySYoiAHy09REyFi
52SGF6Iul0MeARKDbBt+w6PREM8Zl+tlibC1yiB3J3ufpPEC3xvDgJjKbOfdl8Hy
uKTOcaCTtd7HE6FDV8/tdZ5srnfs2z66gdapfmCIaOQTpS4RPZ8UsXeOXuVmbRVF
t46qNNnhYMZmxCRsmYvpI4+Xs9ybAvkgcH0LM+OJFCu4GZtDcryAWFgtJ0wmPzMq
OKm0+2/Psz0rXEzA5lVJVx56KHUjOq9zuqlf2eqScOE1c4dvSiCc+nErzG8wd3X4
ddWixb2iq32HKimEHyOkF61c+ClJTHqMlQYaTYqXuwSfh48PXAO+TGnEycFNbq6s
PSVqHXdCRG57AKPWYAemAmZq4ncI2eML5AYjSkMwZHAQJRaAk5nscAOOtk7ryNXf
tTqLI/Hkq9PkMbrO0HBCjrWmTgj4lhMztd1cIC7Gjna4/MrisrLZ4UPlJdRj7IaL
gdRRjXwsLY3bd+6NDnTluGLwOR27Q5O2G4Uwiz2eTB043bP8WoazC7doOyQekVop
dYlpl6iZ8HnSdFautyl5Sgn57UR3sxF22hCNxOBLlR4Pjm1PrJkaepjY/FGzl8Zz
VVEORMBN2kL6z9Iww9Asa0AOBLPCpk8orqawSk7csHo66abmgaZI9YZu4nq7yycf
B9HyLG8TryNBnarR3q6sL69dWKocxaFDP6m1XI6o8wR08waiignZ5BNhKAXMuPMl
d9YrYzg5AMrhix4qIj8DLXJG9I6VCHcUfSAEkEWxxs6BxcINwsaT8HHNRon4UTDD
T8Van+V2VqKuw72Id0UWTHh0ZCuED9cHuJDDVCRDPi7ln4Jk6wzF1kAa+kkM9pDE
Lo2O91TrSE/MDBQFm47dLZokImbukjb9/zp36emefnPc4xXkNA7EnYXzzITJFw3G
4IxfnrLDoOeD5inT2HHASnORgdT8rZoYABrXnlprz0lVbq1YdRcVRU5esxQXsnfv
HwwJRVDWzS8JQEOXAlAXRE1yboIol7SslCrU9ymt1XCQspG1vj1qvUeeHqDn48jA
vbMC+Kw+UV5HuOjKS3Ffriq+W+gYDIPkeNSS7mI0SDLe/bAxqURwGWcPMgMJvT7e
Yu6Uqh7/O5T4TIrKfFhLroCgpoF94o6qdg2cB03JscC7C16Cesjut1451/j9oUlr
EKXjXw66Iuj5ftkD5TdW2OKpcSqrCA3/rtkGRhDTydNV4J1daEk/aFykTT83IOB2
ZPOCnpFOiH/gbkU+MoyA+cAgi7s0mkKBCeDwfZWglgFSAOzplzUziHcThN5oFtqN
8b0QbpoGMPfsNRdygOXSrrqp5onPmUK5W+WPN7kzNjmigxgEG/GzdFOr0EQHw4hq
ZvB1F+RvHDhxkU4KoJcCycDOMzUUUtW4NExJZ+IT5eAnnpCduqPVBSE5VARHBxMA
fgHYq60a4FGZuJUKtEKAavGFKvj2z1KGXqQd1RAyWUQLbO/6tHQwOpOncd9nZTD8
ifVvwbT0oWgbAwlzC4HvmTDu7KWEyJSF4l8j9hae/QgN7uS9xnoD0oLQii5Ali05
72e2AQqMdr+gRb++RAx9gRcq+XGnfNHxTxL8Aht7h8skT9CHuqXD2f9eU7ZVwquJ
kSCOUESQQLJw5f2Jho7q4MKqE538EyDQ/aJq2cBAwxwfo2wsYiyX/D/UBbiWrStD
R607B1G4mWOhCEuRvyZqrbSTz2g6kmTXvcorqKQT2r4pd4xORFILHdL1Rbz90WHy
T1uz0dYDRCYfYQKAAP2EbUu4BvVBT6r45CRsx/SM8AF6feg5zqtjGN76inBc7+pj
jyhUKdkFQLO6t6oQcDKoVWPOjqNhHC1VdPgWIMOoaywL76eo7doATQYd1T/mA5gV
Qem5xa3ziMQ/hkkol4qA09GtF6ZTjndZ1iDTHyOY6m95sQ7OKXQWvBtYBvu9rIKa
gvCmY0Mp+noSjK/+vUrBb2EDPGBr2YG0Wljwv+60FcDn2z5/QxPGQbcU0SHzFf6R
n/NYj4YRoiFLQlGruStV2CN/O0/Ec4uek0WIk6h9f9I2+HrbqnhkTv7qD9l60n9j
t0v7XtTIqFHn1o/Dp+0RFGNG+zOj2qRa67rBaKPj8cmAdkpPkpiY3DAHnNn5lYhZ
9Up4JDxeBwBNnd1YUveaDqy1J+t13qeE4UkzwtOQvcbRo+ifgk2lIhbcDGh7ZUg+
7JQIgXFIZAy6OzpW7PjbFJBNr30wg/mJ471gqLZJsZEtUjsfZxOyBUyIXJwHsyaa
LyvmjlODA1eDGSyWCjHZyUX6v7mVvvFwhqKRUvVfzc8TWm+bB+9tdqIvOFFeLhfj
lurvqvKAgK2xISprje41bmFoHpDokvqChM9xuq9JpENhUkHkrTtxt2AkX/IKwlBI
tKfeTPHGhGOnHr07Nhqb7pflmPJArIKokXXRcwX/Qsbge3q0aEcm7OAOuK1D+/SQ
nA7lZnccGupH9Ibo3efit+e537OnIUu0M2gYJEgFtcUFeYScBjAhcG/D1Qmtq+PN
+zLoKTv74yRVWW9EouyFmklS1dVVq/hJHkvigFP8MH66oF4IiehGZktUgU2AeCem
WCaMhOs40bdNKOyg9RJBYXHRGiRl3x/lr9s8JMlZn4nS43w50L8N6NeKkYnZzu3u
QUr/ASgzfAsniUZfSeLFazW4fh34rwDbZywssFuz3fB6VcUBQXbiuNpeaH4PKHj6
tICc7RBBXFhO1KFsR/h9W7OLBtGgwLaCqn+LQC7y1j+M8HDPqnxO2E+YcBhquUjx
aW2U51TsuHydNsCO/koWC+OwrTQQPY0pUn8OVMorwlhDHW80OGXI1h/FJtYJgYcB
Q8tx7n1226Gidsl8IG7ACvgI/151aeX4Kk/kTWG1Tqywkkfmw/blXkYRgplDGQuK
3PHLXKjtqSuFMadzuSrkaCvK3BVMmqnHhZL3KKB4tYJh6TJpUDlmRvhMMfaiIjTY
y8LTZR2P/vyoaZPP1Y2nOY40KBnbz694gzfvgUJjevxsrJt9cHmD++ARlrGl9KAx
OkZN/cZygqLv66aH+MNEv7zDpXF943lyWmjBnPEeewCWk6kUoApeZANHQRb/El/c
vq1RRj6USkXuOccpCf12gl/sZI/vePm8A0EKRJGI1tqZiVB7EF6mqnqGCf8xyFVM
Uh7aBHTSu5u1wG8agmAVybETbBjaUvHGWMOa2S3/bCUpUN7zaKuzmWqXRQevjWSp
A7qGPLYiRbchBXICbite8U2mfDiOKVmmYuyFtGPsPJQujtVKg56WALsbwOqtB5DF
eRVdF9TvNVjGTihJ/JLCRHe+vFOaPpuwEyX7/pC3FdUclK7PAFTy+n1wlGc5mT4n
a4biUbe56HAdkFn1a1Dkg45orSgkqQ3zJbkYNonbvDG/H8xt8o7t/Nn1ydf4HuRd
q59X+l6O8hU7xwWrUf23vzPM0HlFGLpleXJOx9EpuBSyoAIz962gNKIVUN4u/7s2
LSkRfJrwO1Ds3IgarExhRekZ9k39mzde0ndkNXk5+5A++1UtQJdFvUOa03RiDJnb
fSoXMU0e9VgxGKhq8yNmxwIY7LXOLM0sJuaPGGoLYYLTxNvmwolwP+WYrCTWlKI8
RnzrJTesVcuqmleE6OxRnOhXpfPIZ5KX7JaNyC5hdtd/7CFz3BPUTcvMan8Ckwcs
CBBucK7xsRmNawRqx53PZyICQ2yvyMcP8eUV1xYOGkS2Oq/UN9p626+alhfuOvjs
nHb05qEP6aEpiU++rSOdjbWDc70P2dL9VZD5gZkGzSOgeNfqpevcDQjG8Cd7WOG/
FFRbaUiwpeOmeQsEoW404YnrzHvIY6mZUMx/6bUm4UmGERcXBF+6txTEFm/fDIVO
921PbM5UE9cuiKOwX94lSKy4iHeqn7cxzqUboGRUEj4WP+xPFVJj9htPgTRmsDLk
OmiSYHWUVT+VT62I5g+DX+2JDAhcJlUSdTiQxKxUw04H+8gUqGFoQDMrnNtZ2m0e
u7MpTI1IQUJwQ91tD1pOiKAf0xAQpIHS7RI29dzmhB25ltVYVesKyVTlCySyjCeh
mR5rOw8h3kw+OthGMLpFCXP27M3YNIy2s9t6EWZxNpsytL75HjDXzQ3H8GsBuMm/
+08+D6H6dBAnrx10VnN13a1XBt/6t/q+6B6A3Z9zPiDet3FbikybxedhUQ4xjT5p
8J8m6Njv3MJIWZ6/mrMAfgWGUOvp3tq03hJwzJWnuvMY9QZ0gSYg6u6uGLzEVNjc
MAd+sx6akMQPrG1EWy9orAAjrxP2OmWyFOYkRM7QZ8Iy8yVLfgHs44tkJeQr0L8Z
/otS5kgNyil4O+m94wvA+Hv3q2n/BBsXeeuQDRcZdvZYX+A30J+OPkMmtS79Uqdo
cXUaLz5QNMC7G1kyqaWWkqOIk/uTXT0S/Wshg8XDAzxtE6wHe/Z/9zdWV4l7KJpR
GUJwZrAPE8CVf5gHuyi0c0kt+xRrGhJIxAzTfWiw7n4Rtw6z8R+0LQ0hLYqKp6rw
+6GEjp2dP5ooNKmRmHhUgWf0U5ezc8xXrjkOGNzf2oNB32F/Rb7uPM6YIo2Rhmw3
11qWAN1kqZGcINXTi0ISo1PJiXAizQtQ5yOr6UFXeaGCyAPRKO34sfK3FF/fKvmD
njKFi+W1xLMPa+2gRmqjZRQKMf7TjRMi78sT29VIm/+dlxASR++xSzx7JGbbE2R+
YyycjpefxplFlQmzRtM3p6Mw64fCISrcou0WLCXpPGQ0C9uOx4ifNrlibZaXvFcf
slMRy1FoLUDSbEdSs5Yt7VjySRVIsxXncwGI5nepfxTUUQUV1u6fn6cy3vp5pEsb
+Y4p6NzvvYidmdnjnMzEX9mWOE2wSmhBleQ5DK4GmWUVV6L28/Xi4JY3Z67c5TZu
G0OVQADcSrClEpvFt3qSStWldPBRjK6BdsnnoN3CR3Ix++wvby9GZxn0ymUxnnTC
mIN3olu9u6QGaIfcXWTGDauHNi9Sjvqqb4LKC1GXh2x+EsGZ/Y+MU22SICiu/L4N
P04Zni1Q+EAqWwXTC0lFrusovy+qXw5EYFsmMB3YNDYlUxtjcZzNpGBax8/1Jm+H
2IgEjt5x4Vvw7wA5fKE5ZM6TJqnJSfJtpYiCZ0WpJpdrq1XZMtSDSxcROka646sK
SqBCbfAO1R+iurtxGXYmsHYoLvGyYn0nH0GOV1ZdAgKLtCLNMxP1FXCpvPPBiuz+
9ZKbpavxGv1mxyplhtUnuqVDcVglgF6QkxB1MMBSotsFbDwCdBc3zkziPlh/5ZvG
nep0x6Ar79F/JEFjjFpVAtQ+YC8qbayDPyCBxhdMf1OImE6w2LHC4FYsw3+zkS0z
VeBobL13T8eImbWS0fLX5pbDHgnfK1CLs1goYiVxzA+QGpJYmZY5j8G9Iw2MFm8W
vFpq1fWZh7p+yvMiUvZG506la4MzyB3hgiRIlACi34nevOFSdL/UqK22K8w4kpg1
4yRvGKAo18w5Xwni6OPqwsf4N7IB/j5GNtJTHejueuu41w7JBy3IUf4iExlcYqxX
rx1nrcCNg5pGVY969/QcXTDHjCTn7TpgGDyF9vpG4ZLLRvbq+ZtLPz79fhVnc9Xd
ApdMzrAWpM179FlSBKTwQyGUEoSC/Mgkd+76wYSSlvN90d+sI46UE8ub/yps3SOL
KMPIoO+TIXSq4jKmU6HTmzcCcsMUI+xEERCXBQCOPGGXIyV5D3Wmn8H/37ugX7ay
YZzZYc83r6GsAUHfurvxLmftPe6iU/IB3ppUQp/XRhTSAUPYxvSPDyVnMFV4uKiq
YE4nBUOw8tPk3kuD1A6xYc2ohnlTQDqTNgcmhQhFIOMKvr9z3WdZKT9c932WWB4Q
I+Jne7H3CnDjkEl7ivg02sD7KDgybjd8cPE8b6VffBtsKbIgWUsQCwpLRQuZAd1y
o6loDiaeQN5jfIidyAt6JN4YEB3MvWQfZsIdI/6O0lMIYzuQUwI2omrBJKl7gL2C
+HHQBSE/pqaB6GLKype3/CqB5NxsuqsoeDjP2uLKjKsmIm1a73NIGlbbeGMKG0Wo
o6juVwrbehFMkPRmhcfY3tgZ1Cy0YX4JdszkkMRezceRMeqLaGC/aCNyS2gbegxH
zYiNfOlmv4lobEcgNEtgHQ6TpqFB0RXyMrskv+bVZeXb0rP5eEGaFjQG3jBE6Ynk
3bYKuSXIxFou0xlNbV5w9iP6PZflTFTuwzRLM0R4njA=
`protect END_PROTECTED
