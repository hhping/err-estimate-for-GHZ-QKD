`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdL52GqfoSdVX5tpUwQ0vCEYaY9AqSH36J+nCzsBj0Prj0Tgd02xIkpAP23PHrDV
6tZCRXez313ld1lYLxeEVGTj/swxWdgsl++an6aT0DJXEFHv0MIjtVU7LJDNejH0
mYV6RFDHrLbtpQ3SLhvkMGtqZGLko1EwuSSFijxz7yqRc/iOFgUz5ogD2qbHXcl9
VFT4R1ll/CbIHks0jJEEwZm2uK1Nbnbf78mdfH0Bd+r+vjMU837dV0hoIl9YzvV0
s8DIR3TPsIcdfPEkeKEPuFPlz69A5+aBiwwihewLA9pDk/SZZiLb6p6g/+1sfELV
CwpAS8EofyO7xPArj3LkexNWfAHNSC5DlBoXPn1pYubAJ6oFSGzjOL2VJHcn9aGi
R6rhtFttQeYpPlztsa2dPOBuQWUoo6I0C0mWHi+MYG92qYEd4O74stHTpZ/GTu+4
Re6ejk9wigT4CbG3DEXSV/0TGjxZD0q1GKab2Aym8DvyPtqi81EgYxRFoursWVEB
HdAnqGf7LTOVuZmyjM3ttMxamrktJ2Gf2dt2CHq0Mq6VGhDlKKjfKv14/TRANA05
FeUFOGAejcfL30E//thzjPBnrgMDQgZfRHKfPTSZz1Lu/mCHmdGvC003G+H7VCAA
rGYJx775P6Odc1UGvemjkMoD0xakAAfY6CRYHWdVe8oAgx4pM18++42abhMNaEfF
jWHwWOcQA7EAWG/AmMFtPoaA1nMwaDuhJRX9QunKeWA=
`protect END_PROTECTED
