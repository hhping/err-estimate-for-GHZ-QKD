`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8AOe2P7kzxFZUJErxa/LaVweqeSHMavZrWyv5PDzdOq+JbIu0fSudCKAOZw70Oo
4AxYjgDhwcl5XQEoEO53XyF+6CGgI0WX01GmAQDPCM6mK20oliXdebvsEYT345pd
YFrrdX7PBLOHrhrIuw+s4FdjCF/1H/5jbGuvsgAV6Mr8rKm0IHxt1QHseWhc3ze0
3qtttu3jfcDMv08ZY94KYBAHEEFLhEmMcUbnub+JHfu9+HE80EkAZ9aKcGq1nN3X
a8M0Yaxq5ntEu1QAJ3gVEpunEUWD37JEGJkagQcdpy+SsZaaTL2jA5Pmnnkz/5Tn
w1VfZj0cATz6tU7B6Nvbb+PJuYzWXVQzV1COYgzGrDE+uixYDOcd0sZ5ecBcWGlB
esqYoBLKqmecoY1HTGFaUdmNINIipRqUMyLCuVKVjrKexVOv5akYvjPCT/ecbcE6
R5pOhLiNXSiP08K5jWQEEOEaDgGT2HJ304Fr0ZYh/WjkAsSjDe0+VDWR5M9OwzRR
pw1QD2uslIiTz70gEs6WbqHu9fax8dykEon+es4BoJHbX0ODzRu1l5AYJTx8exL9
1MSpt+dIygFA8hb0QVyky4XNhv2F4HSnebqMkty7VBqFELKOfuDWHoZKWDtq/P6S
xmvhCwZX27JR89ne1snZCXKUNp7paR7vn8n/EzHcJiq9oyzbSFVxkOq83LhZdK5g
9ydgPsiV0jVIpjsiCN08yHilQ1v+8Fjdmfhb8htWHkPlXxYO0wMGjHaycl6XZpls
IwPAY+Wxz3/fbNs0LhSAHga4TNSvIt7oZJ4Y9HsIkFsWgRf1FkTq60WKhyfqaOy3
aHNhbdyki844zEsZn06jDeMzghCDhYPeld3ZeqNaxQwjR6dzEiYWsAVQTWQLjw1s
NUex823XDcyhPHeoLown7bOy0Nvf8rChtSYLKff9aK2suf4+sjMzRyMb4SgWE/QL
Grn4HQoe19PyhPZH/ryWErE6FrSWnvo4sU9CIu+MfiPA9H5HTX3e9DBZ4Fjpwy2Y
UKfdEzuuyQBngL3sVIMiyAxF2jACkm1aqZU0U6aKLHBMLtjna4ughn3uUyvxILA+
aXqTvRed5tbn5xuRvZfMEoLtCRaY2VcdRLGN5aeALkzqiDkXIjlowvE2L2mzaUVU
At2qLXxyxaNO0anzf5WNO8KevqH70k0CzLtCM8r9iDnVveWh4qWRci7OcDQ1sBRH
LwRoso90VlKbSH2lNyigvciUl8wYUD9LDMxGbycKDGMmcYnLvPXRJdN/8QE5pCSq
`protect END_PROTECTED
