`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhgYPbJMO8Xnh5Qfj51Im1V2JyU0cpQyka39O0HON5lH565J7hVxch/vcU2Y7kmz
gdo48eXeykbRIejWMOJIUeY14xen+mMgtP2LsqDAh9T0uojJNSEglbQZ9eg7WIv+
JJ0bRBISEJTbdqtRhMr/yA68un4bsN7WIAfFy7aU5yzM42onXEy1Q+vK2cjcyWj3
PO8UmuzmBa1TX5N/jMkKaBV/N9z1LkQHmTltfcQg3D6vORCmTbuB50b3s/qH+ZcI
QU8E2WkKyZS+IqvfQcU3WCKG6etskk6nVgOwHQ1WZEbF2UI2kTdnS7+mBHxZ3b7M
niUQmPLo7+4ba3tPKXNij0IohCx5sGxAXyughBQkPdRbMe+cQn40emsEGNlH5EGT
r5/iGou87Soq/3GU+WmnV1GodUdjowUU+QSjekG7Wb/NqPbM3b3r3H1CtYE6bmuh
SCitY7d3z+WCA0T9KP6ert92T2ackHP3F3gdR1d8jM+4HEaSONF7Rp2B5flcDdrM
MNj9tYw6HS6C8b2b+r1SEKCT8eyJOpRemun+plxS795D4R8lVRh2QA6cJtgU2OlD
Bz7uwZc1Nqhy5oxkLojJGhEA6/b7Vqlrtgdn8gg1WD2/EjWAh4WNgKTE+ohi78Ov
OehPxc9FEe1vw0PWVuHcE0edHXNsfZILDymAeJ/yLEuatRvv4tFalIGE0KkuNLY4
fyz+EkTZq8gBQ+klZcC7YqQAcp/WLToKs0IqH3Ve7OSE7UXlOx9tembaPUGWJnWF
rZeYTI1jW4QCcfVcaGgdEOIo9lsBWa9Pc7UoQiIcmFFlaod9fNqwm7CBJC1g6jUj
sMgarC3G7lOPPl72y1tlw1c2rMFJS/HjASCmGd9rrvy8bXVN+1WmXMRZ1ZdH+Q7B
LFF6nIL4l4/t+wm9OXyu8pUlqOA2w/J1Ymvoqkfr+6GKMXiEKcZEvqqR8oOVmsEn
U5tugyb/XFSluR/P7nue/s8CM9FRyX046WlBHBkq7F8RG4yo+xbPA0c1XD00HhSN
pPI3LBEGVQNJ1mDtvYwl/eiiuptS+3bgWmGhibd5o0fGKafdVBhDeGrr0D33dl34
WcKG3WG8bhMtKeUay9URiBEC/f+1unHQ/tx6G1CGVTYOZ0vJ9wnivJ0gXbwBiDkI
Mve/PQeZPtcGcuTwYK6kGyw4h5GIKG3aa8/1NdjJbo11SVznn7syIfBxE6stkUtr
nUFzuMJdIIltOD+Oab6LwWLWNV6QUmuhOORnRAGpj/iuknGV5wqbKeJQFaW/1blV
ajuAz+sFIdv8cWV6Pkry4tz8A9I3MT509BHiyypV4ALFhtWBNcNGH4R49Y/Yf1/m
KSocyyVuzS53KwI8UrfwogyroBmfYkN1G5FRQXLr+ENS2N2/yj0XI+XoGMnTUzHM
D3CNcw5yP715Uvm7XbLswSdUm0Yy4u0tj5l4R587m3R40TUPHm3QjePVnwHOrS/o
+rnGEhXeMj3tqRMkHLPuW+HRSlPew8GpgkMXsS99ZxB65zre8mbkgqq2km3K8cvU
x6/IZTREa8lu3z0tamR8Is1SlJKPA1x1LZY8TypNCqD0J5vj1oscSxvOZchTKQEm
+2e/w/i0yI2trWJLiR6ErzQs8BZpNtexabg7O2swh3EbIjRhCgrkGTiouiT6YoaB
i7mElB2kdyZM0w+1HjjGD8tWL1arM9/MMgbtvnfbarRl0s9mJfppdkrjpMxm8BaB
zH7gemoOLUVQ04rbs+xxPsxpNwxLgd+DK8KeF68QvNbNwKM1N6yh9BX6r7zAuAC8
2GKkeuEcNauqxG2VIz/3eQfE7zpOT+UPaeDZOEr8OIwgT6+Cdie7lWhHZ1Gop7ZZ
IWqCFFs2HAKnQpWxfFepTyznHnfyINkKgh/Vf9nmgdZ01a6net/3+PMskiq/EOFP
MUsVTScA469DwCXYqtl8FKipmbXyq5mEV5+U7ymjO9+k6baeuOogDpnX0fYBc17a
zFCRxEiEd37Hrbr0q00wVInaxex7xQOKKNXwtBjVen5wBSZTPH37J1IkTN2T40xX
IPpCRDbJYoTOOJ/KOGKVrD2PyG/RDILIOCsN1kPZe71m8LjAS45+CFw/YojqwbYB
L9Sdlb+o+ns7PqWT86KHtBex0tDz8hBY2Lq5AKQNpo9x976OAvWFYQFioasXte1R
4obzc0t/AH7nrFf71saz0buLf/Y3BwrACuEQtM0XfmiBa9xbm6yC2dgZ1Q6pjTkH
ehqSuLSA1GX1sBRwFVK4AhZC8V+19CA9Oasy36WMNMs=
`protect END_PROTECTED
