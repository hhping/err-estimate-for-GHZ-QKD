`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dy0BEKlhLaRmOTSrcY5KOrCeGVoFDRgKUBCW2R3a/I6uElkjmAspf2sNUeD54UMZ
z3oaxav62AGvw2KnwCXxm0BV6j69NiN52nufxbfQ15cjaSvUUVcPQ9NvapaxPl7D
nis4kFZlLIOXZw+VaBexjLf5xHn0pgvepwIV/Are+y8nSIRMc6ch/2jDiVIK8F+8
11ZA6dHcme2LkDD+WVRLWA2XyLGQgRt5Bt3Aw7skgtSlIYpp13tRdf4MnDgP6c2g
0WyATPWbmgdMqAPHMD2uqTZN3eqRdJvbntEHdwUvS5HOsxqE5eEjdHY1ERUtlP/9
DmUmnie9NavAi5LsFkAt84paKYDxQ7UyOP3snb5jXruRYAIp9C7AzSr30HMgA2nY
x+5Y7ZLXVvQM9/HaKF3Ch+E5Y+h+tBH7bqUJjm60lccCUCg2mzW/CPIaROUGV4Xh
6k/B4MNkfumr5IkjhgRz4waR4kjoEzSgn/mxKIz0LBPhgx2k7SAsozRr1kAPJ9/5
+Asjq5BtKOUICv5fnUXmeOCIlBPaKgLoF5NrfnEttX5Kc/w6okf+jtcJ+Jm0lzQu
`protect END_PROTECTED
