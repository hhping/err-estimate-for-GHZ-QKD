`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6uy7EtIdyzJlOUl6QlRi0AIqBaKM6G4cjgDOtvnqbtaTjpQhf/N4w/KbiWKX95Di
ByXhu+WVKUhjD6FHHJyaRnvbw59GuWNplbyY05NlPSCV0xo0xzUTIVnw7bwrICej
hv2kJy3NGr7hds36d/O9Tp4qJvs/dZMsgR9CsFZDasi9BA9R03W38apt/TI9fu2v
js07sxFT7k7iQMhZ5qFpzkxFuiwqkkvN3q4YOB8eW2NLbWvY3gUc3y3NGY2oDdLd
XoLeE9eQtyz3oT6x0FkPL4TMc3So440etjQi3eboNFWITX7qZvmb0vV9nxJnSaJm
Kq3wlDCoSCpJM7ErBMBuU1hsV3GAABwlWTOsgkVvvpEqz0KWK95imy2CwvLZP9LD
70UdwXVtoPzE9IeM21aGHe+Aj3G5UKzzGA4M/meo4p527xhNUS4SZnGJHqAM6o0o
gMKFiUkKl1YTygO9GAFrVamRlwiy5aaSD/Boy317LVDpXmT5NL0JgDnFt/jJisXF
yAd0F2IxjxvHebnJgipUjVzBK642PDTIvKWlQwW0ZGYr6fXNATNG85SAi03JkP5n
aFOgJUzl/STybY1txHS0ZQfz77wNmzudDw99CjMtwldpXIVik0ZP3rDXXYTA6FQg
ElwDY9XADUpnzqY4l/pU1PjUaSGIJlSpfpKo9YlxhAFnvxf0bh725SlE4Bntck2/
aNbhb107z3Tt3jw5zp20+16NFo6hbyh5BJrPtPldUhM+F40w+9unXeWhP3TBh4Qm
ZTv3kJdQdIl7k5/1QAAbbnKSJQWL1rIPXKlTNvawB/Im8rsrmm7UCGJiFOoKR9IL
2ajRCnvCjILKA48plNIaZYsX1ThHMoBlI6j2gyW9gRGHdyL465gw1t8xDjBo89UL
ZnjdGAJDJoq78nnVg7vyPbhFO1eJiWA79XtIH6YyLenkMrE/eACHJT1abIcISqL8
CJJTY4lwubxhTXS1hAijur488wcv2zqkCkkk2vmbGpMXrao6JQOfknQtargLcuV6
Qv3p1dwvNbss0ZpfccGnpE+uZbIQHg/S/j33MjQ9wuHv8aJtMKxY3CY4+mO68O0I
UQPBq0RgthPQ/x2OmF3h6CkbyCWxCkr++SKX02BhOjryEwJ+uooJc7gtC+OiSraM
11Kx3lJ4u/HQRUN0EpnCGUjTc3uAkXK2QI+eEJxa3/YcDBNBoPQQsn3Hx7YlD123
aRi0gDuKSsFMi/LwqoHPFIOFimYIav2WCp4GcrjF1bkiPjH82fPsvXUKIWQ660wy
guCO05W5R9eUX5YLZWPSoYhcHOYLVX40R1Y81IeWVLqdDsIey/Ddw5UDnbKzz0t8
/nZlp4GhfhuoUccFy4b6m8xoWY+j086b9fZ2riqND5diq6gmj8bCjNx18IjoCP8d
m03sw+MRCLR/7pA/FKM081VYKJEX6lvHws4fKA4Zh8Dxnv/zF9xIUtMihhONsWKI
Eez2DVS50C14gZmYE1WPvMW5Ko7kvnw7czqqusCk5gu/QcXpOV7LQdxGXiYWcbqH
agR1Y7i97xQ/tEIoX+ii7CcdjYtbQK9KqtNV3vHl0q4skjLY2OxfXJX5revxYQuu
5pGeaxdZKqk5HfZT6u4W3RVES3FUBkgjavwybkssQ4HrEV8n2kXbv4WUSIimJE53
hW3k4/cZst+R6rNb67/ML1RucV3/fSe0KfCziKmzro3tbTxvMN2Q/kX/2Mi53Ymr
xoFyeEC2HB8+BAdltLNHfZD2GeFiuM23wH1XfD0R3RUmJKfkOHLr6s7mYGPNwRuO
2U12kPqbJPi/ZILmfS6VcPeB4zEl8YOhBjkk/1ZlJVo8YkRHTtWaypFUJQ3pktdA
Q+TTL1QhvqVv26UMztNlipYyX8Hd0lNKnUHXGYtuPu3JD+h5udI7iu8B+GJlmhZs
uMx6eBPnOZhfKrQZPK38I1JjIwIR265yH7OBtiD82xa6w/0lM1CodbKSbxiorgA1
7ciXtN5fkgS+SduBgGRgfzMDCaA3u3KlGGHk0b4TpxArLBSmYtLHQImM+OKR3IoY
H4woxDy+8C/biXL+0a+8IgqZOx8zSRJYjP0sP/DPaFphcY34nialalMhytaKtHBQ
thne9N10ycxSV42AlB598WGG1SfEuyvNXJiUTYuSveRoj2izI3qNwsvMIRRi8mZS
cN9g83xtw1EXWd4VYqTQpXPS7Y7Tee7Ask0C3IeABMGoCT/O7TebPVmyiDIIyXju
iyyphP/nNek4GYgRuCojC2dSnfAh/SJ3hwrYpV831alK6JQYLBM9HuZCvd00uD6f
FUm2lODZsqJgtZU7mSXCvoRWuBrB+4MohYJiPFQH2HMkar4fcw91CZnZqklNqyGh
T0C++/mrdJqD27Fiw5y8y4tbI3dflU9s4jmGIh5a4grznhtqIlo4LXn13AY5pzcc
AWhM62FO8Fgzh0g/qhFGntiuRnCLgzYLwSyRLQTzL5ijKo+xp76Rj1AaHnw4EOFa
oAk9X/ThuSyAHNYVSfyPkUOBQTMzVzd/4iCARn5UjScY26sJrfEHxHFPKHa2FRRo
AAh4kEE5KDJoKaoj5K4SO7odXvOAildgiNjf+681OAV2g6XnVjKvrXaqKt13mq6+
96dgy+HR5f1kSL1558ZoLc1IV/ZRw2C8BJsk62hKK0MmFGsixPzWBn3wBg8i7JSs
5i1vw0OzPfI1wTB0/31M0HkBYCQA5vN6/RXFAm5udgwv3KHrAvC570ZwT/pmuUeC
9+qe0P73A27n4tBP8zXNZPFzRTUHt+fEiPfYa2rgu5GOv2OIf3uMEXg/wJRFv7we
7gKpf5vJZJfvdTVO81xOb3DCOKjGpTcF01zz9+5GLiQ4o0oAj/q5022RcmBGlJi6
xMY8LnBJY8vx3DLCGErdPhbxtasmtx3NXnBD6Phi9ZUSu1MBSFsWINg6Zz1RfJnh
RqwrCyDNaESoA00uh0V9RLNevDGBW7O/R5HJrQyPLxS0Xv1i378W3GoY9/U5Xrz7
pHCNHdUPlPItfM4dDjJP/HvPoNDNFh90B44WnTF4LtOHWvv1c6V3Po9ZnS9t8Fg1
kx3FSaCvf7tQgaD2ac2ra5HKppO4bSdI2x5jx+ghP/6ETM8GgttVE5Hzdqd9oFhx
DCCoXOPF1MbyVIoVzs7vtH1Dg+0AIikenx1i2Pzw8PNOfWJNApi11gbDh2Wp0EU5
xJHJSIpYdZqVjbFTi0YY9IlZWGgGep7Ayank1lXy+ASpM5pM/nKxXpw2AJ4/BXl3
u9LCfh0IGUDgeqV501xlt58ob6lHrk+7CDlKWZQeRT+m2CoqcX85nCMJ50r5VCXB
s/bvQRlb5wwyiDCwyhZmTTf2/FMK2lDE5wQlGcoY/G9+7dyY5RBnWTX+oyWMys+s
8ZRBn6dOZpDwGIjIMFB/sqU5R9YVK0gOkeRH8KiF7W2Ko/yeZ3mu3k41URlr5vzV
YG4Vk8cniQ0maPSJlqeGWiynJDWQ0h6SWdidNlEoHNqy93W7BahfW9u1utHtcn7B
iN9b5e13VJWDfkwJ+k0fjN6y9vo+ZOrNe10jaSz8n/QmSnbnCC/cxSGWU5ZowzPx
sT3hLHY7fQ6ruwNtstbtbeaG71JcmwXznDxiQ/OqUskltXxjcTP2cnX2XTJw1F+N
E7uyoAIHxxYRcuiMbFpuQ428FBU3iiOBI3RGRHGnv1SkYqQC3mEHHDVk+3u6k0p4
HWia16zDmEH52TJ/opJrwoxre2ho9rktnQRjlcPeYqQrfWy16mznMEDtpExLRR51
/hqjv4OnKyJNmjjmGICXkYIPXc58jWT2qPZVbvOZq/rF8i4rID6JklTlfCm9mcQt
IAY/AGuJP5a72erF/6bnPLgtf20on6yWAe3JcttEOGJ+Qu+vdvnfey2ijPDmiYeF
Ec/T1yUCU3G+citIvMkHjOfWtsT8CgNo9K1Q7jypH2w5Kdy+ZOvjeOE2lgVbJxwc
V1zMyZHRMZE+LSweEkt9z89QGj9xZDqchsGDikRQqsjE6FL/DvMrgvGtioAgQISM
HqYmGUJXjJj9IRA5mhFx0zkFZroLPt2dnlJKucy4nDgzPeTH/MeiboABI75W9iKo
Qm3iWQnTMiQA30DBaxnvVvUnnS0zN6lcmyv5muhMA75NcCJ2yPydEkSEdUZHcHQN
680264sJiRgZ3+sX3NbKvA+A7xe4UewsMTBRakyMpd63lYR03bBBtVVKhFa+RrpH
bip/evW4McmMI99E1ZBWEwHamkVezdp3Zmld8hIWJtQrwprCF32lDOsQXnsbEfUS
R56EYDIvM+l2fxKcCdwk7I5o8Q3Bt0Oh/2pV7k+5cN2cSHlTNXbMLBJPeZ6Pcgxp
hU+7dwlOlC5hBK5X5j8Eb6v41I49jSH0YGiuZdGVfdkmH9C1Vh16HEwod1YUr3If
hnEb33fPd/qB1YLZf1xf0W4Ol0AH+chyYecR/PY3v+R1GUrqm8nyNzKvu6iImI88
IHAQdSs9NzJ6lIHSde8hOZQn+B4odmJzLrBeECbdYtmQRjSb/lNngFWI3/QcOQzB
xbsfz1BE+RLoSOqNiy6ck5HOvM0gl6MlJSm3NaQrs8asvmHkun5KIK6eYiWf1Yug
5teWTHIvPTIaEBgmwAe8nwh/mVDpNvpBSPAf37LdQkhtArU9M5CUpC49v+/JDv2d
dHLs8Q+Gn9C0okEb1lEfbNWIcOtW2fGX5LW8lZuoUKaWkyv5xpmxiwl7rb9+1TtP
x5PbJUZZuU2GDbKo13FfLm1Y4BoiKuN8XHKJxl1ZT03ZDbQQo1Whk2GM5Aq8tw9w
1oc5+XYTk6RDdhQ8xIx3xm3qaufPN5eUyJN7+JoS/gMJLA9Lsf8RXm0K/BIJXpDk
afL1j13ZR47AElEO0DR8Ypii6MHaywPzfPi9LEjzIu8WCm3G5fy1P2aW5G1rAV0l
Igyp+15fRRB7mYrf2nEfN5ZdpqlJq9jKGudvnC+FVyHQI0xZac8d7TPL+TaSGqJU
s06Z1pktSya9+e8ry52xIdbqQjx8i9CuHq6SOevTB+y92ZbMOXndTTSutISRFYSW
z3KDaEA42cPXcSYySJZX8CiWAnVvDdRLRpOktqzVURZCJ8eULGo2AUIJAPRK+E2G
Rz5mpR5jSWVzeB31WoNRtmfQnfSZ/egzi6SQg61mcfqQPFFif4FIw0X0IQXIp034
5M0lcp5Zamc7GjxQPF9U3/kKj79YECwaA//5A5PfqhOXwcmcH7rKg3EkO3X1g/CS
rKRQun3W7kKNFufYodz0Ignc4AJhKrsSRPseY+9vskAsaLvgDDes7tVf2aLi3eGK
fCf1JSok0s0nqBTwuYff+6QBBI8I+02fM50z3oNfgkRgNVIIGopCF8z9v5oFlUkC
4e+/sXep5UFEeFeA6KUirWYWQwWVqBxBo8qGJ1ss6JibbXmmw3oxUhZyv7FjYaJ0
xZVDizOXmQa/qsfV4p2m84viDGbEvip78t+oXWESAxn3fS1AdwufSvK5oFWA85DO
bW31oCVR9aRgFOfShhqC4VhXq6F7utDkRhar6Rdw0Rr67vAlRTBQTCCMBhtqJfko
41QNEbm/P/Tc9q4vMOcfK48T9Evg0aVcd97DbmfYCysHPdnKquW914dA/tgYwvX1
rqSCAt6UJyFGbBSgujxiyvsYK0MXUZjTiA++JwCDdWtcfquoWxaDJobRT4LJ3Cgt
wkKfqaUdgaVgrJYW0DEJXk7FEjfVLc077BZPg3Ce2AH55NEGUdjl2Y9pojjgfZv+
SE2HlEEvtbDkK8mDHPaFNQVYld6KYwjh0mMUkSIWGmI91vVnGeCzRNtrshHlucqx
kKzLKty/o2sRP2TodIgqR4n/xTNF6Jf/esz8EiJnjdyMAzXYWQYdOxKfYMpgwsmD
2/PqPjSCZt1HzhlXbkwR5ltmj+8Gmvzsf4xQNb9Ylq6td0NntZ8uqK1HL8uLf8yU
cYyJHnOn8AxhTmYxD4TT3wXGWi0hNodh9i6gVy3qmHYqB/CvGF2EyNiJadxoi6Bh
HktUKezpnIFq5h9U34NT1RH5jTW00g6DrmGj3xeeF52ynRDIxKP5SouzMvlLLvue
e+m1YaA8g6tC3lFcbenPvBBtustzGHpZiw+JEqnzSuf/o9MjMCfaMVTpDdxrAND1
39KNUVaGXlAkFkiRyTuxETcH2YNrgxFYJMr5Kd7kk3GUuipQI66TKk7rt+ULfh9Q
1j8twjwT6X2IHTNk20r1quSbIqYvTZVxo0B0bsI64cWNhgChkv/gUT+Gy3FhwIFO
9BquIIUz6kSY+sJHm5Cp5ubun0uV1fS+WltxZXnZEO6WQKOL1G404A0ko7Mz1EeI
o2fyb1UcYy4z80B+kabHJkjBJo5MgUxiMVsF3FlifAd7Wv7Z6yVJwzutTN1tTYMo
so+YsQoqFfgSbwUudAgkjgGcHDl430vdail+yqHkRkGRiGUqFU3rF5j+B1mZ2p/Z
eB1H5vA3nxE9ieV6pPJsTXkS6nqfmnyd4CtkywboDqQymu9qQcegd7dvnixDvyeH
UOPr6XDz+FmuImPekUbGuXC6xVcI4FjKu5zm2Nc9LNpEM8ylZ8AWjpdsMbp5YwQr
tUE/AECih+MMTe3uQUAy4LuchwPwJ3qWY9Q0A6VNB/uhqUTsQrSnJpVvdPvpb9Vd
9xLI9Os3oElCL0u24YdF/Os+RpBKYwKs+Eq1A24JbhgQqRLxogDpGyOBXSLhPJIc
SXf4K661yug+mgx+3X6iSBXuCp6LelwtBXAv+/907o+ootY1EKb9NLipQ4umxGPU
tYuikZVHPbTE1N/OcdJUG7P7k8oO9tn/M7jO7K5IBxsgGJ4DN0cij9Ps9vEKeYaB
/7fGW65vIojfYheikzvJCNuWgh0m/bR82z5zAGVUFpJF8AzukuClkPB/VvnHrEHB
q6hMxIGAadI9Li9zvIeY7tTFrwONGGwA6gEy/umcOGUp3nMkmECT88HD2Xljg3go
wrGkY6+DxfmVkM5R42a61sT+smZ3hFOF41IXlpdVRpl//eA5QX7e0tL5aUuR2Cni
rQLojJD2XtdSKuuFmPcJQ/Z8TqNABmDrigbUP7oItTB8XGCmFqVt6B5z/l6HfuHG
5rlYe/xxBTPB/3jpYr10dt+pVweK/ag9WHptfwioN4Q5WySbja70IXS9TJfxqTTy
FmvlMBUX3vlF82wTNxaJ2piQBEz9kWQUTJU1SUxUL+6ak7PeqJ2nPxDNNiARAdkl
sjYfT/RyL8FzSIb/J/bQ/yPOloBqjdtq+c4PbNwJ8QGmuqmQsOkwd93A0EI1QAyx
pyGUo001u8soW9BL485Rs+H0dEwforQCX+UsAgK56m3siXAYq8gkCAyYrwxME+r7
2dAdjT9UZLDnwdDz8vOU+xpaIp3PHo3L0pWrhmTmC821cCjq9sSrDFqq3uwAOCNq
C23iaI7syk3yCmdlNosoTZ8YbziifjXms87IRBX9dMmpbVeE085MCUVdA3qvEUPy
G50zMkagLKA1N6DuXdGprGwHO31qqtqi7WeQXmDK77KewrGWrzdoxA2AM9Lg21W3
JSkmidMC04fuI4C5/yRsYV+I+Tn3pi7PYWejzyPGwJfkhlQHp2kONFIoEn6C5Wf0
wVV9L8SBku+YSwTMm8Qr1Xj1BT7kY5SCukKl+XlSflepQWAD5mfO6nh4y1bCVUzr
sxRhlwphgENkSZULWF0E5kAT9emYkVIjwwvSmd3BZGt1qI54B/rgH3fIQ0MeaHru
oGaD5ERuVgGnkixokyaRn8Nr+5D8Bwu0ikStxjVJHYWQ6RbV1OLOqhKgOkmeBzke
QDvNWCZCQpj1l6yFM1u6LIKzkmsrBLUA1nwEmh1jO5AYthAd1UuWW0j51oFGkN+b
rxxQuCWccYcYW34kNLHmOjmURlgWjSCR/tmKWYdNu0NljxJDuylg60DBWep7RzjN
v3WrdUqRRcfJ/8usjkmFRDxmpvZZayxzyfEBh5Yz7jWIJ23D4eDHK7SCwTxGi19v
ZuOlFi8gW12akhKNRdBWtRPdDs7fcOVfjKYnGq+H0bktrSpahAowtnNqDUhTNLHU
HTtL6cyJW51R5Jd+zJ8K3FSG58y22ZDGcroodNlX8vtsqC5w7ovrmh0jJ3/otFBN
csgnx1Bdp6vYG2oeMKXaK4bgG0zcly+I/EmuiTTnhM+rmRgaPOMXAT8MWF8Rd4tn
TU1lg2dW1jMfY73pGVqllHaZrTJyi9GoDG2nCwAPzO39odCkPEZUH3xXN1mnHlow
Q24EeCdcIXUz59Sf+wRizSpfzPtaNpKzsAXk8LhVBP6dq8ilN+i0u40jcUNT+Neh
78wAXl47zyqg5Q5dyKnxgUsDCYQufUzYkiuHal2DUDh80uZKPnOB526QIiPMiuot
wvV3hK9FM9BW6SZCFPIhgmCeROtKOw/1Ix0RwfbYMBEW2Whhz+ztjZWbklUK77t3
lwY3FXs8KoJ01KMY52499TdEkzYgIQLRlGUGob8VrDvtNxLu+RtKqjYZKx5C7MfN
FXuZGpiHkXrqkqqWgSYHqX2Q3jntZCVu687HL5hPFatqCtentPq5Tz2kbn7xwOqR
CnrCLG0L0LSXdjrgHgqi6KyB6oJRahjZ8iIZFPA40ir+imI9u0S5QjzpNTqmI/73
Va8lq2n+yi/czFcVPAsO3M01tIWAa/FS0QVSr5awTHVdWTLPZJfHPC7H/7ziVZ1e
eJFT9+IcwfkrEq6UluTK5kwRhvrmMQ/QE1Dc0/4h7DPIl41O//AYw7Gqwrk23MVA
ChwtKT7BGCtIUJx7QpUpzOfaGCI37bZFNWxc8t4lTszeeqy/fszCxudFUDhISAI1
NgEDUU0Q0eCv2mT0iLFTyFnRn4MRCFw0dJ7EZJuPwvHGeLsfjsDOextwfWh6Fsmh
ERmJJU8fhkL0G7sy3XDZHGAmOruaN+tIzQ1h4hx2jrddFWlTaO8Um81A/sqlJ7eM
Y1UyTK+nXWVQONyS+1Ck2JSIzgHUhZ/78pvNla5ea6hfKeaFyInCP1Zvz0VILdpz
yhVRyoTBYBM/ReEemFuuw4Ff2wYfuFDoBAb/spWWuTJb7UC6L4NeH0/WxPGmJfA3
BSUqq5Yt5trW3THFe6Uv2XMP0kZgnMp73HHGi+iL3eCmWxqfUMN3zj9S20Y6+ig2
aZcZnVA8l7kPINmvvotaqnAmJE/h7pFvIlMNZu8HJBPSJsRFvpvG/L13OSo2nfam
XPIz4GGxh8E3ybIpt65a+vrooVj6vD9y83gh3lNM1Cz+ZJNeW+e+8pV+Nv28YCH9
Qi2KlBdQTvZjB76Wxi5whHjZpcqPjLSvpn1B/TmhXsW6BXjRxRZpx3ziyUzYUkCD
fQJRcEZ6br4QUOHfhy4Er8ui/zk8RUHmBXouaPm34JOj6RfUMq7HNifZPIS9yEQG
jFSUxuZCEh5rrBJHLbNSHwJc/OWAMCnbEdzcjOVaTJFox84xR/DYNOGwm29X7WmV
0Equs7IZDiTIN26U+7z5OyJxcYIuJN2kOcHgG5S+PDcvc0V5V02Aeot8CHw/uerj
MbWj6YJY40yMuP0WmOmkFUdlUpEVZaczPnHW8/e+tOSlZ0jG6zVFNJ/Zmv5kqlCv
5njzeiUjlPyaFBOR5IRC4Q0Fj6uuZGaUhbAMZOrZrX8Y1nHLnDa1YaYe3/usTFuK
liFWBccYjDPgCWcLKsKTElszAu5Tg0GkbUAkLzUud/esYPF/vIyJh8+4NdPs58gF
f2xnOMz2irexcXYMb6jdHAUJv5tRBrm+E7X3+oD6D2Cp9mlJ5cTiGsncXU69Mv1+
uh8gtySyt9RNTbs64NYMwHJGLsgSjZ38UblmErTDZy8b4e9MtOFEZB7e7MP/upRl
b38B2H7v9otZK1lZWMFgRCZ/FsqZvyONS/sZzRAKC0qMyDeq8TzJ5xkMa03ej0Ws
5RR2D/hCOD4FXEJ5KQH4XqMuBhcWla7hI7uCX5XnRFH9h1WHes0zm7HXqbWqLPdL
MPHk79qy/oqmJM9rYyAWvUOtEKl0lkioT8Y8SfMrzwgr+JoHweJDhkjDSFQNx9F7
71wZd1BpfYqzTlWiiQrbJemjoXplQtZHWO9dSDBks7kV9JTYH5m7Pzfl9cO0ma5a
bnGZgAZ4s8ILm7MYKAt0XQnR/v40zw6B3FjkrEiyockBSTOemYs6n8HDfA7HE8ZM
BDYnCyCEEOWQrhKGU0vGcb1ACY9FU6+ZyFZ/WJKnev2AiouCwQHeT3/JEKQ16LqN
yyOcbpB2p+snwZKEqkCxokvJs1n/5sNBIOU0z0EVGb1manAbhXqmNPWVhOI2MyLq
VkyOl4624uZmswQYYL8t9Adsv/ckKMwFBwMj0jsdft4ZwXUc+w6tokvHnpTn8yEC
NbdcydzTiA2K/NVPEA0D5BFqlRYBKFyarpYIlysMgb7mW0L8ivFW2nLWFIAjS4TZ
Brv6l7f4FxMdjyRiX5O2CIDQbpZrjD5w5BawK/FmiBmlkPMPqo5F+e84QbeGct4P
n5x1lF651GxNh4mr/7aAAerGjSCDrJBycN/oXEM9KFzJREExXgT9ypow4KhS/lGD
HzDOi39gHmApdwNziRviyioXDtmGBYtuN3BJBD6g7FOtRd+hCCG+3Uo6/TkOEG3G
wmCT9rpYeEgCb6a58tfUpWedIjH6izGNorFqEAp1Ojdp/9g8/3UTSM7LuFgbUJMU
ibdp/GBTZ0GuAmdDrAboNneHyW1gP19+GgpB9h03l+8Js1F+wVPPmW4a2PDWkUC8
SGBxG456FyvkLIzmoAWsZ0keeZfexUypJIxiJmxaq0jxd1uDR+me+2oVwdlFaSGq
FejfYOnDwN0R5Bde/KQJUizVZui2lqC5SJw4/ou9IYvY2bzbERkYgRICw6bzzkoR
iNJTjxPvS/52gvdMNvL6F3uYENo2EMUSv+O3+WDbhFcngh7ud26aH41J2i6kbPIk
iVpJFgPRu1VRLxCv7rh2UKIMDLvnlSFk7NPBkpg0RClw4jo6A/UWvT9lTipt+iEj
EVa7tVpi3/4WNYaKyw8orbUeH6KdJxi6BjuuhGSonwTt71fChtRIP4wwO2Un8vhw
XJ/bLD2/m21ro6Du7QHTsqPIX5SqQFvGVHiKKcH+J1TQJqxLEmXc3ZiDkkLqtMcA
pRtqKCiCNEWa9caLm0I7Fcts2Q+ntI6MJrZ4AuT8ay6/hisZNSj9OtOF3j9cUzzq
uvH/djIJ74xj9ER3oyZpKMhQMpKs69Q4XOFsvv0bffM=
`protect END_PROTECTED
