`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9BjVJPFYoe0hIRgKdZoBN9AvagDBSGKyFxXbH+hdAYBAHvFJHk0E84uZCG9yXhB
uTsvh00WX3TUrcIxwsRXKXZhX0lln1EG4TIfsHVoyrL7sttSCoDltIbBeYWu+iNQ
TmBkNw1eJe3ZkyytcE3S8jd7TRuMY0dKgcPPWxaHFrFJcWIMrc55CUPmShPWyroo
V0l18J6MOYbQbIttOACSdw3sstEGpz19n1Y9V9godhcsoZWb5cdwSnRSHrcaUeo2
dhFivvercrFFnlp0Y5g7ukJQeAHsiFTe2FWyyCkfNV3IH7aT5ZkO/BPgD/St6+Z3
77yNQUK1Pqt5fmXVtsqa758kE27TlkPYj/9yDQ0BIhd7+Sla2RZ3gYzGqvcawaNv
4wlclhxhKXMAeKlIpyKcHnezpEdk8ixhXvdnvWNjHXf/cHuVaYjnxHR6qFIfzxhs
h7iR8Q6KNuDgUIEcauqa6JDpTG+8MkQSTGJW9HriapBUPbmqaAF/ZmQV/nx1e5HS
hzJVMwZ9/M28i+ZgwUyDqDOCnRLn7sVk9nb6KYfOeTgPqw0bgYsWXTyo3BzThHR6
NLP1WKMYVpKl15+fBzO+Gj2c8Z/wAcQrxgDw51xkSsw9LSbWDrPafZVHbTh3Ps0F
3Nt1HcQo++r44SOYc6EKDQbHM7bF7G2VDqYx7Wz/XIBlhMJBAABgZk2P0FqwyCnR
KoHpNmE0xyl1z1y1LkjqTrqM+5wEQvlOE82+xurKey995bDDQxcOV8ufjMFImxmQ
ErNEP6GX4S4SZtngYmzi1c1fJP9kt88JUX0hMMxAy982qGOpQ/Y3UX+W08jn8GRJ
nLnzdmMow9qjF5xc/K8niDm5tYX24w3lAZFLVWxNuFBzN8Kn+1fJfBP/G2KvDuJV
BwkCh45CpQWKxYUEtFalfjine4VExGkPFZyu1nI8PiOTulO0QodkQRe6YO04vAYH
IIVUIWODQkjPEvCiNtotj5tRkwB+EAyiDDRcKiU/x0uVkYkNwrVDFjzc4cqtZWSK
6K+1DYPoIgtC6YZ9O68pLxyRlNZRIFFWXRR49MtIj8DUgbkFYhidAf91mZnnhol+
q8zoou6VmsmkTwUPa9hy29WnW9wc2lZEbPOPXgqk0lHuCCmIxh9bNWX7TQraLbdr
Bw70rg7yCOPT7HpcE2Oxaw==
`protect END_PROTECTED
