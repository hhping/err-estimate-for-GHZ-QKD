`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QsOALMQ7KSSBL8NuvE87YSQAfb0XEZpOPWacs4dnsmNLxreXSIf/JqIk3NVT2+rn
EcoSD4MkjmET8wLeVDJVZx6Dy4+lePofDMPrwHO7/Qrrfc2BmaXwkuIiHqIVmjM8
el2ZRTBy1kY3QTdPBmhOXTkGXs2B4v4nVFrnR71MXTuXuo3pEcqzVy61LPnoIQoa
ubdZVY8391B3mQ8cJMOpPiszj1356yVtkvI4vpTfdcUMa96dQ54m/dw4slWzZoV6
qGtG6J/qcOroIDX/HHHjl8hkvw7N/vEWie7A65qjE/j6r311Z3igWgqhdcCT9U/5
7pJn5tboJ7dlshNMEzdNJiO9FeHsp5xl+V5BAebeCKP5QxyXviIY+ECYAS07kGtQ
RYtyAz9XEgtt18r9ReDkiGi1a1KYCSvL2GYmD48DSBEiM4l6/gMtT1mX9rMQp3Xg
OVnHiXDfimOAiyfSrVPNwqSIkDMgb8ljwnzpHoXlmqfZWhDPCJyTqQ7YXi8TiVk4
UxfEOgiTy81hvu83PKl4QSVOe128tWTTpwYjXAcA2NeQGy4ZdVRrmGOhHqy6ysok
gg2g4fqMMtinHE1tYjGXrpjWYdc8rjnmkb8zLDbG1L6y4k8+TGD6JSSomuqogTIU
KdhS0YV3kI6QrrnvANlpig==
`protect END_PROTECTED
