`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzzamWR5gKXHlP0Dw0sySEzuFvlIKjaYFy1X16Lt5CtWMvBIL3fadFQG+7JNmQDg
ok+raolOnc5cn/DD1VTKgaE/S+/mxmXqaKB8MVDBzWMq3iZ5jPI+PTwVB4Zi1Qbx
3LSXu1kvIkRAlV1gDaqAqlLlSHquGZn6XExSwTaDfLslTy1L62KbYIrgb/lKSLBh
PjMXZP2w8tLKG5MY098znWgrwpc5cRJoL/rXBSCUPAqD15zH4MeEmV3tJmUxVBm/
MJHyjC+aUzI0RQMJ0K6HJ1NZXw65OfESf7lvvCSKdYywhx8BZUHCHuXuXO1S6PRP
WP8lXtFMo+ayeM4Ro6RM1w7AC2rRJ0NwzBogU7Yrs1nzIO2CWSwgT33FXBDtQQ0F
JXvk+LuHSLuKJl+Yx3gL8ojV6XUAjNy5AQGTop6Tb9xwyjfOohYIFlsfevGewTzJ
I18Ml7afxw82aXPdPqdcgYqS34ibVQhEWaXYU5RTQMD+aM50JphUujsrpbv44o6t
oFAEXlUvuKxpkSccXBhopClZDImql5C4reRjFYbdcdmdgR29X8R8t2tUzrBtkwX/
SvxQJjfDQHudfQg+GxxU6A==
`protect END_PROTECTED
