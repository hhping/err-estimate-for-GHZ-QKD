`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFoWT3Y0DRZ5jcWip2w+gMF49s/Wm4kYnz1dR5gqW+R375gRzCj/5TkuypE3t0sh
o4QNwrfPXItaf2fOYmbIQDfbMrAkbEYjZcePHOUOATaIamqDzNc5VvlraULbfODb
D3uM8U3Gucsf0Qwr78km8ORYw+qZCN4WPyWkDg4X6n5qwIZ/yU7DTthEtNw2lsHN
6A1Rkmpv4IltzEJlrKxGgshfTPTNNCileUvPoFn6UlkxlbTi0lck4IbrLH1HzzoI
V3ae+1CByiMUXWq0uWm+fwcAV9FszcjuBxJq7oDgsGNp68fcqG/GeyHugapz3P7j
ao4f7QY0LNejBJ2ECzjI9cchRQv8jIV6p3mMudZQaSgr62Uabg1EazaC+68+oR/L
s8BzHDRUWtvza6J0kOZEg50T9LrUTsYswS1VZpKKJVHkfseN846uq7AdYQmfMHUM
m818WdfeN9slWiZI7mqG2iFKW1Awe2Dy8vD8AlekBStkH+qZp/hQM+cZoioVORaf
JUS6OUC1unb/yBJym62XQKQ/idNU2XvF6I4WzRoAzfz8UDc2jOeLg/qIOCxBmFQ4
Od5fIq6/wuNh81rMAyAHPWbth+i+QwK8ipV1nLqr/v0JOupP+lBril5p7IO8d57N
C0HAafRrTeMxa+KRVo4Nbh8oPtHZ7nMdG8QE2Fy+2y7Hkq3Eh726CAy169VW4aXx
vJCSM5MHKUtrDAizl94OAf/kBfNQtNm1BJZiPaivM9g=
`protect END_PROTECTED
