`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h868XXtLSeYjFVe+ab40uyMVh5LLRPaEUMsq7OjWKm7u7CTxlTF9XgpcOG+BZ7qp
Xxk2ko+QDC4KAV9szDsRUCY6RIJFgEQEm1D+rvnJkjauONgqaZi+Mv1JCpsrNLk7
z05pnpMjsa3XucL6n2TnqG/g2OJtWR48xKMzu/oC8b8me5Wu23KmMnxobRGDc25g
HgUcMhX/jCIGkXR2G6GmFvfgz9bdCK3W8JG3lrFlTbuU0QERTSRP+RUVvEF8Heyk
o8Yh5tmN9Sb0oREeOXoJVgrw5g4tZpakCmV0pSdunEk5lx8g4Ffbx0iFjhM5gdHZ
dKzXiY8QQBC8KHjZMyY6qfWtt7x4TbiDA5+J4DbqqRedqEy688F6gXuJHbvKaZmQ
OSuIw9cpbK4U+G+M4vudugi5gA7FEcE10UVpMLO+4eHQPahpWN+OnvVMMdvzrU/7
ddJmu5Wr0p74c/V9ky9eOm6Uf6jY3C5J2LzKZKv72ZIlRyhfedV8YSOoZNLRZZOa
x+UYvVIP1HJiFz8BblzZjIXLcsaj5482A7MGMsejvywlV9BZWaXEcs6vZFiapKM3
Uuu+9bBxpGBzjnNbt2jzI1Pf6MZj4nrNhZExUfRCCRf1QDnF2gXWsJhHVoOFUR2V
zOP/5UcrS3MOqjLCXhIHXZLRxrLFT2vzMqXK8jyS78oA3vOxUBaw5cjA3eUNWxj1
sQaI2rdSDfbXX308+XL6ubcl2WHYXB85/vRTLL0GOy21JposgvhcpPT3h7ObQuMf
pG8agtHeBFR0gbKbBPoZAYZu9SmRdJZqF5QazcX9zaz1W7NWORmuelYoPPbzVsPG
zO3306P/z3jK9f9+jwCMvsXw99im8GpQtDJOKQspYO6I1c5TuL6M2keyOZACmmeA
qtSl5lHJBmDm2fGhbg8DaQfgEwPcI/inU9hnjdmLV0hSswPinn2U+ihNMWAWwZ3E
mm9X8QL2WYjBnNd60wYnlKFl+2oNrazP/CQhhzp9xEiixRqoQmKj8b1KATBwFKB9
7oSutST14m29Skd4dH8Ky8EXRmeMkp4b+IfqWhlCqCLENKhWCaMQJlJkAzZyrUAW
om5rhBvy6D+yeNqeMLE2UUcOaQh/AENd9x+gevrbuH6FmUqTfMzCT8BANtfoJczY
RDBUIkXDgbkKhuPo+jGmDCiweXwq5t/73jGKbXG35iIroOM3gvarKAOpk0bhTZCQ
bbq88f7qjN/ur8Jpya4TnEVKdYpy2xORls98X0flexut8TMZ4PrkWO7VnKdhIJZE
mhBa/L8bnpPaLHI+A84nwlgpKvY5c0C4UpqDI1Tj1h6LS2DmrqlUPVr+ehJku4Kp
NHsrDySCbjPPCPEojgwcK3+K03npREmPLSUbz+iuNc5c8sVvxYtsr0RvnscYrbn7
tNgmbKFoqfcovTz/RKu+TAW4MY/5y2HC1M+aLw3FB5TI03edN+r8PK/A8oxSfjuH
QFmZd0pHAwoR15iIo7/fnnoqOcKCfyDCgbiJg49zJe6AViJUFuvqK1HkfLZzSybe
II2n8HkXbmqdZ2YfVAqOpB9r95D1P0Xjcbn8Ea7uWEHqv4TiYmQmkCsFD34uzrgL
no7mBA5NjEY0UrV+iCw+sjRso7x7raMb5Q4wTmWM6f0gYNuUTvAh99A+gPWllZFl
WDudUWf/Ra2CXK/lAdWBf0zSbgXpjP6CPiKABWe/tCtL9MPPbw57dEwI6Pn+VmV/
mFH4oGYFQ6bi2PhBLvrch72Ea36NzZUHIunqhCiRIruSoRh97Isv67lS2lh9IPcP
KLqKDZLq/PlO2I5yTAn4d628hGML9iOqQhVcOK84tHMYeO5QdToUxp9ZOpxNMPJ5
rMxUfKOO6GbOL6LIF9PnjtEbD8G79Nnznjq1GtfYBv17NCVsVcYG4oVH3ynR7Ehn
zLw4vAIvY/on1R7ycRmH4NekgPHrqurJSEjuq/6Pv6Vvgz1mMvXnc/MEMaC49xoN
`protect END_PROTECTED
