`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rsaKhjiTBxXxnXPNOnC9URGOOSz8fMEmQ/rk791TE5dkemY/avQ6gg7KSupu6FCA
g7zf2GwQcL+MdSN92XCpNJKR/pP6fCiPOB+Xz8tu40acobue5lLE7d1Rij2earM/
Hgm8VhwuDmD7y2e1a8lZqtOMcBRjLEJfVqocU7BlsVewlWVhtUGcqOF5ZhO/8xsR
kFlaFW5NLkDCkOmt2323Ybjl6PZPlLBN1FQBy9GI6WvGYwNGu27UY/aKGDBZzamY
8/3jdjTELhBPRYf1gG4MlE3jWhXC8LxF+qdKmMWcO6eycGqIuFco+dR4uzqH6epi
meaJONLmOPseCt6dPjJamAf+Udx7GJM7s0iU7HrpPgMisKiSMDt9cugKzgqwNiuj
aSdYduvyprc2v9jgVHqrK9+CCtnH1O298PN9wIStk64u609pHWUb7s90volvpqxH
JdUybvxlQ/2k+noCD01o1qZo3nc08lrDdzgCJzNs3vC6m9fFziGJAwPx4ApuUbXh
UC2BxU9ZK/Y46o9RzUX7jJs/egCoPzaj2iG5dNnGQMhOcVYnz2BW5jwbzFSY2VIo
mzCbYC67E5uVWS8NCt5uAoZMR4+f91e8tvfs0mlaVgPJ0m9P7fBQlDbyWACOBKBG
0eIhcgQgO4+jRvbfFLqtNmWhaJiqdUNah9xvs3AoNwrvj87C2Zfq2ZaXs6xIMJ3r
EbOpYrFeDbV1Sd9uZFcjIXxRRX0+F+g7xveK+L4/w4Q1Ki97cefU3h9ICBuquglP
ZmrYAIyEqmdUfGcJM0jZ9xmVXr9hePxdbsZlqPypYejnKFkmB3/yh6/J7h5LZrTj
cjmmVpdh0GNFpQq7v76rr+WOJ6TKN5lw2p9kV1xffshAgouVGKcCI3uvlGXLM902
vcaYX70H//y4Q+YZWEmyTKzAqkwv8IVlbJtGyNwJesG5zEfvZJsyT/mLCAv/2Npp
tUTOic/IyaQ1yE1jjXWWm0ZOEoxImEaUHK3HL5q8pw/j8zwDruZW+xr0tUIJg6Vu
EycTchUD8Su5juB/gJ1Qgiuj8GrSrQU8BhYR6ciEHyNvgxkxunwdPnRK/sYR02uW
nEO7qGgna8HP+/gr4wOoa9fW6dmWS4aN1LIvDnruVGaaKp0N1Nc/vo1AV+D8NqlZ
un2nVgofwdKwNXaSwaQK0gZZka6PpdDngBL8xOaJW2croiX0zrPQ/jTWEElgofyQ
OH7KPRMujdQExl+Mm8wDyY57slD1bnrYy3Hk9OY5zJOeY2/2TXrzhsJz1NlspSVp
R5fWxOr8DjyxEqg7vRzNdZjc884bONMM7UUxlCgAVK4ZDwXkEupOJYFhgweoK8jV
lBCg5PgD9Q62hFU+7y460JuLTvw0Q99naggNra6RcklUc/VlS3+TTmPK5WB0j0Pw
fVqB5oy5AP5eaEfQoGEJqPlY3PUpTauN7oJVY2RMkucZEnLa1c5lI01yO8xzVsMy
ZuzKX8CES8ztdPzopMcYmgXJar0vqja2g83G1RUPvbQciwEPd06/khaFGDj1cqQU
60Prw+TsTSN1pNJCZqZizu6NCsUMcQZvLanwDpEfuH6Gj78mNH1V30vpVbRF/C6Z
pfCoSiFp5NahaA2aSztap8T+ECMlttdjRf45drNNlnhdlDh8eUdhdS/EhagbYC70
wNdsq1BIG1qNtkFXl1plwP8GkUrlgl/iMSNZViw8D/DzliDl4NcZ4W64QzwWDp7G
pNqq3lH2CEjHr048L2YucG7WjqsZ6Ujud9uhmRMsVu4R88umkct77Wj0rX3JFmuC
hsRUgFmaiNEJuNV42xaEAVcx827vdg/vSEGplosvT7fvLMXQxjxHpgjEYWSvNjm9
BXK3NYTWjeqsSV7BLB3vpnf5nFBbcRBI30arPzdIfykxva1K76hHR7tCxBgDBTDl
KdozEPHp8SX4bgl3R7k4CuwBoW6rtAPxmT4W7XaXsnr5xacWXwUn2myPp/E7MCBp
xzN40bZ5Ums9uyPMuKwvDhxMkthlKUkv5zJXCeOgZC7TLnOCkTecxDfRqkJTVdxf
MJFLofND/c9gdV+xGLuMvzOGvz3oxBpbgMQjLeD2aAYLFzXBHgZITJQ8GYduMzIp
GWgvAy6ts3yv3Yw6949FFofI7pAQH4QfYcb2ZvT64DTJqdI77t0XwFyIhwqlWLR5
Ogkd+Rt0n3vP80ZHTFp7tFOoq0q/TeN8lmqQ7WDQsPV7fFxdAtHktgMhfcQTGYVF
AcuUTMzGd7TisZQe3KbVIoOFqMT4Mz7Ukmcv0KjztMZgw/VNyybl1bxq31M94GpK
`protect END_PROTECTED
