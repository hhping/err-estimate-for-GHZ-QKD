`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2GAtb0/gFQ5YEOuPxSfoqqsBGX5fCn3jxs5R+1St7HcOY10koadtr9iLY/NmLnGC
76r9iGRlzGMdFWhdDX5zGoAJK4pfnZlSPTqD2eJKyO72BKclKh5iwMf0p1gnmKSf
3XWJlkPML+AvHmZyaHLtQn5g42tkGnbmZVR3KtWzf1NlT27nLtZgoGkJqFtFYOL6
7++YD092jY0gcp0RM716R5Qht8MjJ6PV1JVGnTaMwhBQLp+Qhtdae3etEO/Z49om
VvzX69bBM0QJ4jg7bQ/cladgVSOMolrpzhRMIE8KAm5M18B5W8D/i0Z9ueUITIy7
l5JeodZ8q7gUV4UJwXE+Hf6qBDLq3fZ0l3KOund2pDkWLL/26ZmP8gXz8HPw0vW1
jINlfvaGN82vsinhwjdbYq55yg2g6PDBIuqjZsHaAyhvcPAS4k7inBRws/ZSstzl
ypJIZBCPY47ivXvWaCCYnLfZf6T1scyeLHeINKHJoPrk9gvt3fnet8dmKIT7u5n/
JiLQsQ/NvgV+kLqnNHwwRatxnu5d947pHsRE8EhJcLB9B0+oXmn4CL7l4gc1y3LF
iEFac4YirTEmL/sGeAJeuUwOOXllxrVFmrmElFvDbKYQu3B6N7/RtySXJRKp5dDC
zmefnhoKbXvCfKptywLKhHisNjsPN+7J9K4zzdLud+/tw0juO80lU0lvEAEEjmB4
eN4IaUqsh8iYAz131XUTQrjSXWg7v1ssHRGTLohOuKwSGhM5HXAQwydTj3MMJ/2H
CK1tCuzNwjZxTt39XCtT5ywT8tS11XmFY/CiRMaZJTFx0BtoANziDF9CmWwNyX7g
u6CicF44pQwjw4BATwvQs3tSLp3lhRIAxrb3t06YR/XcSVuOXXBajM11kyjZHNtI
LQ2JYmoHhjkE3Zc2ooWZ3p3FeD9765c+4WE1fcNwWz1p2Z4TL1S3EIT3eiFE/sM7
syst3SGx1fOjyzNExYqD2DpLlLFnUm8Bn5nAaHTXjRDsQQg8OCyXbuYlRxQA/KbX
6YMHUEjeqsM3eb9rygDc+LS4Hyz1BukWeODkX0BuN13gnbdIS+3u2Mz9Okqo+lvq
rehetUQV6vxXp4ISGl0tATXlQq8hnpdJRj65cd6xjZHD3fxWoINfkvkH9eA5E6D9
pEuO5i7NscgKxb24+gx5YHCkO7UPfz2L39mnOvd5TcQoG1kdmG15E5NFTAnK6zGE
woIzhnpibfl5lM8GVe8K2UTGUEsbcMZVwljNFSZb9W4+e4++a3SauxRnUQhrwseZ
B/YhVnawJXH8qHVVOzJzdnvHRmXuTaZ0DGZWvMZCkvu7Xj3fJ+GdoaB3weHQ4ork
`protect END_PROTECTED
