`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoXBFwM9F7T0QZZKiiJ+ScQixuiMr+qDNaaWyU/7JMhyhJx09aJRqGfXBug6OIZO
wUyUaSWbYi0DN54BX7+To34Xjps6GuyHvP+EmQX+eV8MupmysqCFRJ8H2rDiyNYG
NDuUbrolYgPVf3B6vQDzeYPEtGi2/qN1q54WIkom7vCSWgoPr/aA3/Ms1PmhTMPr
zv5P3BbR7MkUyyNjii526gScBTLG8pzqIKESjRnToPW5lOIEPwtobKSdRR1c7JgS
YoiqsnAh9wm+nnTQk85GiUv10Igyj9yOXIoUob14LjOgsjQ8sLl9OuY1SxEtqg+e
n/AE8Iqv09I4zugteWoZ/qi9la3TINSUxWKgAvGKZ0Nw5Y+nnagTU151IcIoyIrX
ELMMYzKWRm4sPftiayluE2eoSMzZ74WVL/1qFQXCmmCGK1iVyKeTTsuFlDBaNEm+
YF3lnAW5VmgEqTm04eFPdADp4tiAazbHefhu4nLqQk1qkT5/oaKGrtJGNrHDEsqX
ZIN0cSbjO/Mvucm6el+CART8goAgdKCvIn4zNe3Q1LbEcJzC688oPZ7DshpaNMTO
9kcpnDJxHCm/vDWGui+2F3sHCcUPs4ydN4G/eYTXzvFb6pzuer6bVZnRUDq95hao
EiNTiVYSlJy2cRipTLgC5wfeDz6qwqkL2SHJcDjj34Um/vhxkVsztGsR2VFw5A/p
yROPoiUsNXWODBNBapRGNYxSxgOlirVTCUaG5FIEmcnRO+M4KY35CtUrRwcCxB4T
rmKFqGW2e19F4r6OB5oF7eNOWUnQlkdJIn3ioHpquW8Jsp6adypNocLgYqypo5ss
L8N/IObCihsyHfnc47MtlopgzXnppr04i4Sb/6dG516YQeSVYHCkhuGRhUpZt0ul
b/ZHBOfk3g44BYJs9coaq6kC3A4+5t7Xmw6BO5AQVlz0rc44yFNSyt7pmlguoNNF
HjOeBsszWzl3OTEKXyB+O77k5XxIUUs2Udlg6rcRVKsbYse/MQm8jIRcHC3MqY5n
y82qck73aLIj6LAN8PY3Jit5awY7ol7Or7WqkCJ12V/wIxwcmGShRsQHMXXkAb0i
vUtUU5gyQtQ7ljSAfBkCyDg4BvP8sV4LbgRsL+xFA8bUQoo3JwjcO8vkHlAGGEWv
vwEge0FtKTWRVgNynugxkIXQXL3HY83VafHafH+gdzRqjGIEaShglj3FUH7sfEKw
DPss/nCzM59hduN/RJCyKOrxXkGa2SUOy8V66RV6HgG9DDvEPC6FjdcveDSJwYKv
7tFGzeo2D5WRs1gG276XbSXJcX5lQ+q+1fUC4TtHU79QjF2th7ULHY+88GyjjEsW
AJnAcuE3GgHmKM2MNUmM2qLSGvd2ZY03dllqwGoQfI2fKQ/nS4mTbEmN5sJe0Ht4
vvnxADtZWOS+IIG91MYPfA09PNrHBVUBE8R0zNFVTDd6nLDHHnh1GSOpk2f1CUmf
lQ4pWuBOZCRSwwH8M2Vh6g==
`protect END_PROTECTED
