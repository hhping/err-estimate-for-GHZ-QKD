`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rdG+GaODlpOufw+quaS73Y3dFH0iOgi2TtAjNMGlne84OoxEpmiqtdiIGcVYjNd0
57KnHaFUPGT2i5gxrjBMo5jmSE96tRQs4bm6fuAsMi1HUjvjXv8O9wRvLYAmOxd7
9btCIhbJ8Z0PlAj7cg9C2g5pLl5x1HUKcRIH8atmDLDkUjVEYdqukhtMOaocUiQM
odoasbSeJkarj9jHKWgzyvVacvx9WRAWNn6/4K8txv+FpLSiyy4MQn5GqOsnYwrx
sbaPNinq5uFl2pYb6kriYAClqY4TsnmqM1+rd+4y9oYylathj2kfc16JwCi6JkBl
QUDrgNeoZIcFWme8ddI5GPVJv3tVSd/h/dDSu+E/FzUGDHaIv/RNqluaZocJdxIX
KBHcfGsBuvuqj9kPvpbtAeSIBCIcQebqU4GeFAYY5qiMcBLg5MYqVqHtMcpql7tC
aty/oBEejwdZ+zuexe/4UlAoU2Pjv9USQEghabcVdiu1z6cm4oWtCy4C//VqzVhw
V2XQbx+ehjO6yeq5whiWGgCeKaO2fh/f4UZ+3cTI+5H5FdOF6dOzVQDGlkV9FhqK
2BnFaSwf3D9HfFK2HKyA4A==
`protect END_PROTECTED
