`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHSxQb179FwT4qhY7B3x/kS5dSvrNX41Y0HImygMrBs0+EQRTEZWqJHqjnR1VOao
Dsd3Jz1DI3VeMY0vP/vAHWQq7pG1N3KaN4uj90wi+LMCRIHiyClwNoia1jqZvh0k
xmRvxZYOKGGMGX5lv3WKlf4pTvtGGA6zYvXAlUCaO+Zvk7ZGuWG1+tNnrEJwUIt1
ttG/dQnK0cjvHItDhcHwsfU1vcPr0DqFNH3wpOJGH7bKU30SKRjpw/P8Qp0pm+DJ
Anxnzv57bEvnsL7seDlI0/xaaqyo58AG4lSb0oMpZxpDP/nYsfroV6C1eSeprk1T
1hLk/Bd4Opvh3NHqrP5AzkoeUBNaIYCmmsgiY6jF8idyevNg2jajAT8RNJUZ2OTk
k1eZ/FhXvzf/Adc+vhp/Qoa7EbL5fuq4Qw2ZaolRt8UFjSi7duxNUUx56Gi0otw6
ku/cffvTuP/kdNF9ugYHW56+dal7TG4nWlaVFbvW9Vqpit2So93ybEOw8gYjmJYE
YqhLZRKDbgsnmTbOYBNwWtYgKZpuRW6dyhxSFiYsVXTbN/SYJSHOJLCxvrU6LNBm
84ZiAwcdqpr9e4LwKN7C1I2sI38OcmidZo0y8xNE1hDQl4BoD3qje7IXtl6sk5go
Qqa+wYQGgXxb281Ux0lhjSmM9vLkcZrPIQLxNjsQXaQzngz6u5aWMLTD0cNSXc5Q
EhG7np2/pRacejkD+isz+NKQxJ7YpZn0hURKFc+Zhzxqgk6eTnLgle1XuTtH4n9I
orfUP/qD0K/p0+DkYkSmKmg6XAoBG/KfmmluSMd6C8lKWf9ZnI0OWaW6i3q2+74D
izF1dO4zlHwHZctuJiMMR4G++n2saOP6zm7TFQZmzv1F2njZgSE06vBmPc9xosi3
lnZpoEAjKgZdc6LblrtMvSdJRAD7zg5fhFZK48NrUw5ADpuKgykMbJ6vnUtgIn5D
VU/pA43nCvbBI/6ZYdC0SqHr8sMCZLvYIy6TRRInBr40SA1dTNE3Csnt4Vt8gpu6
fHpMfHj6Son2ijNSKze9LPjQtKVzzT3rcAMbM+cTAuKQlOe6b0bgn1bAW3MfdDRy
jJRrwBekh3VwA003PMslCEDb1LUNi4Mlt5rHp4hNm4IML9AF5qfszfthVpSYyzrM
raS/nq+//KyhbDXyoUTq8NjK+dpr9MYfYsYBbu53/dmkCTY9/eoL4hmjHY5AV0X1
vhmRdPt+VVtYF9X+cfB0DoI0NuJbKVXrl65Lv2iN1GkhVCaNIPrpjiJj+kzgBKT5
HLqtG0xURWYQuUql1A+a6m+aplnEDDpY78TnUpIL5CfxRKG0EdXqQHsaMHnFoGTu
t6o0bOGK8SLFQt4tbf1I17N4MgmGz42WtIqmPyGHUY0Ipr8pbKaAqQWcP7WJj1xR
AhlWICrrfaBaCuVhQPS9QJ/EoIs9u6ObA41ZLgxUkQCZwqi8VPZu0azWgsp7US+2
uZgoP9EFo7ixJfQdgc2vrkS95h9uWF9P6z+UH8iOTkKEjyGxRsJ4+cXi78G5d0uL
LxakQDNl2RrEp7HcxxZRDGncXhwk/s57G/Ifdju0Ix6UkfEfxroxkki+WR8v4a1x
vUcjfM2OubhfvOc7UMjH9axo1zcCkroScJeTLtWBpH5gUxEedNFxthsAzH2hT/qq
/4yxC7I+nYEEiAiuMfGLpRCOMHVrJy5bvt5KSwiWOXubV4V6wNDcLg4bOH13RlLI
ahjk19mPewnR8u2aIZcYPOF5CcamEeAH4cdHJd4f3u7YQK6QGZOAWVmEeLFUPLg2
jkPaB7hHTYscQy4rL2PHMOO0UrUqlr+PtYif1VC/pM/C37jYVtUc7DCnkSf9Ci0x
+f1vtBcU0NFytIBwbTXMo+qMp0ddZzu2KocDMKB9FnBOmlBUFlBNNaZhEdfDEQh2
+OfyVgTmvxmQo09JXEj7wrLCPt7YIMmjfc2Mk0FBCZFK0JF//eT1OE0tZGkVEgwS
pol8gyOeLTN4c7Mm8NvOOmIs6dvkVZW+QoA0Nug5zJGxWOxTCJ6hnCM0yg5dtHE0
DJ76/fU6Ef8j0hzgHokfA8S8kjBGU55u/YIGi/YcQHZl5i9pCwjkgl2Ev0Q6rWzF
UQlgscACSi588lO1RkIhdQRpDkKn3HqI4DZ82BluFf2HXSS4i4xrCo4hkpHG59zx
rWkFRrMRxhQJFR6d9MRBWPGaFzCjdXHnppWXTVZO3B5/aRNgu+v+MfHCu2VueBOc
MoGjnrpaskpXDuIdoLhFIwsbrckFGFNmfScP0Au8+rjtM9NaJSxTGikLPM+yvjFF
JCUR6qLspyq3woAe/2Ma/b34JV9P+uO8W1vMvlE48mHNiPuSw3f1AmSiHI48hUJ9
Y699L4anLSos0pafN7kSj2FeT+gZiiQTDO3c4ZGEN8wzHOZ5HrZV9tJq72JHIgbe
TLIMJwdwKr38hmrnAl3p1lVTeOkjNvdq7uWbV1veStsPk6S0+kTSLuwky6sVbSYa
fPommmvTyrh42h3tqzjLBvKXs3eVWS9wky61RZA9GWG0nOpzlU7D85mxLn4ZZb0r
WtgPs2fPaoijOTG792A3NQSjQxIK1DXjq1HcSf1UXI0yuxQOawtRdo2AdxsYn0Ir
ZcwnsapSb0X2DbfdMmdAQmlUBj9gxsKWl5dBruPVO66xHIlnDSozbfl4aIfp/1e7
kdHt3+klQkSKtiDNuCxcuR1Cf72LPK7oC0JPdeStHYKFLElrnXl390KDWhf7SM4S
nzJ9BtrwGn3AbgHVDr5CKsH9kd/cl37c7AqCacabaD4MfoEcI4fArYEZoy/vMu8t
/+jzkeJ+QkxBbFU4+jpHn8NHgBas5J5t3dd0AwpChZIVlsAwLt9sP4yQM06gxX82
wjkJnkZAenaH6eHbqN81wa0KTjTNyoKOHn03TqAqHgYkd80vScWAdcrKjwgz/Okj
exQFa7hkgX8h5YAkr8iIG3CM5OxDfS/Axyb6G1EVLV4cwbmfNubCqw/5qXxHiJOR
xEqE6noYuyPuSv6RdWNA/z7lYrdLGIx58Oq+ifttCh5K9S1iXthjvvefbe4bO74X
pgfiLwRXUEWMEzkuQa+qL/iFc422hqR3ibqzbduuF1XXOdcoP10vDLfgmMv6e+GZ
9l1nA8EcmeqfO7L+jue3aNndhUmWOjyZxdHOWOYMtzPGgpo8onNvKlR+EzV9tt1H
9pmx3oY3wk8hajX+m2+2Ow==
`protect END_PROTECTED
