`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGJHT5aMaR8ixRciH9csbqEesLXchbcmPCkW6Bjd5CJfpQMXU3Ptb36WKXsOgzv/
Cyw45kUhbdG7Y4b9Oaef/a6sqZdnS94Jf4zZUUJvAR0TCp5MqJK7pwLoMH4zDXS/
7FEhdZwzUfePHlcoRgQM/Z5klt2TpIXJpsUNX2PMEaRBnJpAO7sEkYP65akSjiNS
t6KR4y1nW8PH5U1ojbx1hNbcuDFRxrW2HvcQq9bzYVWYppBdhEBcZUMrc+ZRaCrd
L5QqXhGRLXZTMcoMKyshQzybcRM1wMF825FJM5lYOrZi3vgl+P0L24gYDXp0BzM/
/2KNYK3JZ97X3OWih5pr9L+k40y3sBAC/9r9F5WwFySA+eSzLBcMrQMk7H1WOEes
v+co7lX8mX6tbfvK50vK37OnflEQfkpFJIVB+BuuCCSbxIqdda7AUcGNPR1uD0aM
2k5Hq3JhmJ4owoHwrM7AmjuKpYZNTsCI1A8MtOrDfmkMhYxLAn/vt+Q7xoT+T8f7
iZiJ3+SoFPqixcRleNwFm599NWahj99shL56DLDpoA5omYtqcLvK9WCIjc+nWe8Q
5TQ/Qodlua/Scj7cacu7duBl3qPfrjOzqG+CMC5PNuZWZEw1mQH/6Em43cnToUwQ
LRMBZcrwIq9zZ/fBl1sP6346ViNPljCGOnZkqaj6uf2KRGfBejwqx+ua8WUcP0AF
rgcoSrGnu1Mbc5j9xxBDYoP1I1rkZFAJj1LJuDjjOeVLE4FNMzeGDIPKEVT+KPrw
32cQyf1JE5DoIiuXYTtS1MS1K5vtCL5bTSAj4l4ax9RBcvodNspXvvh8hTv3Vu2x
zAGlDyXTaYoZJNsi2zJGVH/q0zkMD4wKJi6hqAxT/wEUfalP4Tt/2Ngqajpglto3
cpby2vpFXHgjyeO7/DHHc+BYcaLf/97751cZb/QogjwoW1HAYX1QVIqICj1nuweh
HE9NpNCCTZbiLJKjsxNCmX4a8PXS8bW3JxgZukStKRAieqYlDO+9sGxZI/yxBLCe
BHZbbhZ1+PMQ+4y25BMbc24r0AoTEhd27M+A8MEzVbCCgDtae1AZlGT4W0YkANef
R3MKJvc75YaAFxHCWX4AHEOVnNu4Jh/yHeJJU1t5oQq18x7xh2cLLheuqbOwUbSA
vjZ/SWjKXCgVxbLGRu5cSRNKcdaVnU92Byfwm0rtbjYlPM7dCowaks0wrrNXRW6A
HFnhUAAhcNCTENTDH1aNB1Ogm4OIw+qWv9T+8gXHSsLDhCAjtdBg5dsTdgB57hXM
nJxyugGgFB6PWxnNXtXTYWf83IYgUZyLkfnfDDVFINFaIVgybxLk+QdFN2EQFeiW
V2sYq8a3w9JQJz+B4orTcg==
`protect END_PROTECTED
