`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Zk4Zvh30EQ9n4Lz2zmDThtfaDlwE91DzsX96jRPP5ITzmY++0WRDZ9BzkikF//w
zEhJRiZoxkzt9lmPYj7J7N/drTzCYoFGuQw/tB5skabjz1Zl/9iALLjznyCSlSmA
kcSUYLdNJqE/yHFbfZwSskBKbPVAxZS11vZ4Kx76r5lBJw+NBcvY/0WxRCu2FEwv
RTUE/z9UQeJE1xIz/6TZUL17pUdmZ/18+kzypJmObwZtCQQLhZY0WZYNfixYZCSi
Siv4n3tRAxGr+wunXZyNHr8P30E1wRMofG1nuYuerZ3gRsDRKSaC2jBGZm2Yo2KJ
nvqXHnlVftWrIdapezfhJk+CxaZ6EBM+VHFXejlBK4uf5zdzuETCbK3zMmDF4x7r
v2NT3RdNfaA7Uzdww2SEL0o1foWl/5SSkeiv/NWte9AKcLYadAWztdReZZzk0kIH
N/ZN29KFhw9npkXf+eCr4vdOVP+ImaRIQ3pe3Gn6+aosOR9d+diSBl29nYubZ6H8
XAkOMEi1OxCNJhqipUEPBBZVhyCuSnOr8w3+6rXovjGWO6nrNIAX0qIxk/k+2kmy
nziVMRmX4RoFg93vNXe1cM9hRpthtpztdx5pZlZOxFZXHOTxZSDXwxR6HAtpKCWY
E8PXGPnZi6gAUly9FnTT3uDnASrHNhEpuikLERzEyLqjCUbPv/5xhWMgWjEa71s1
MYzdTDgVAD96MCiXLTEhrA7WICIDmfbs1X5zmkoFlD/lddjLM2XWgD4F6/zssuSu
ps65wJ+zNh4YZvA7hH7RMTcxhiB5Sp9VehcuNTLoBiUfTtSvtSFHq42sFPg0gxW7
mi2uZ0lW1xbGpL2IfYAndPVXyxEMdRlfo/8NnanQ0ZlbH90nCNieae7GfxguQQq8
c+6fJlPqEJYFyoD9C5z4RtB7+IZakacb7MTr1U6uOb+Pgauie1oEc9ldsVf8ZTn8
lmljpYEO+mwey5goEaz0JhP5PsLzzGXMl//Qhm9bkE5yNNi/0tViTr8OaMhQg4xp
02fuR38Me9JQCgClc0529Ta5M9YyvCfxyFGnWXG1Hv6v4X6Z8EIN4UYrm9voosYY
SYcLxIHm8dEtBkRN1xB3YqlFyLAy/QFv/vyvDsRxE1Ft49x10CRu2HMY/l+/JWu6
uXRJd5CTEGVjpaKnX6PXm1Bey2KoFgHQWa2ENozCC+9rs3VGJGeGHrX2K624Vdpp
VasxqmQTXwf0B/kCHF2H7VLUes7RuqFgYVHFv3kTAV+Er2dTtUhxh18YbY2YAl4K
R4Wv++wTsu2EEPrXGAtbrcHWDcmUlCkOb4SnuMKtz2HW2boDEiGkKC2H2WRirf55
WVPFPUO4gxrk4JlWMNB+vg==
`protect END_PROTECTED
