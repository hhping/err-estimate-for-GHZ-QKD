`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htKxwZbLBuJPYxl4XAQEZfhn5ITDmh7XmI/lwbF25ysNotKgn6RGgCVGOxfV6ACT
bPzaTocSYBmInjfu+Axe69ji66y5YCQ7BIJuia2WC3qZspbffKHLDjbI7YfQboFi
Cqeg2duWBNh0aYPkYbvg2xP3Jmc4PIKjZV5LNQ/J/jYD5OqHRNFQfSSXEN8UF+6A
VxAvxJKy1a0WuxtOVkg6v7t68oWvyFH/AFvBAqD8zXAn6iFb7F+oxAqiLXPiWK5V
+Q0LWKasuodBMjqKAjK+4UfZy/rd7fOxlLVkoccjErO4S8nBsOU0hIS3ZMrPUrSY
YN2yYl2gC2PHbg+qjxKjGrTn3FAWRxM5wjY2bIFO5EisxCS6PkoAa3XRFqK6q17Q
cdTnoIVjSzLuJZN5Si4igwBMWV/kFC86iCl3J69Y3okAU6gDtT3R6Vfr8hE/tHuA
rNtxidpcc1nGz4+PKLwN1oLXZCmWXvjb3orVCTIhhnFnT9ZXtXfAIFoVJe8YJ2W/
WnkX6kRbPLQEEWur2FWbObV7bZ4K+3upHt/eDDATVyxRNwOlSe1JFSzLGXD1r9aR
qsTVDW3u5wjqEa4Amccmw0FsPbTal67wSTMPJ4EsguqWTBEmWSQREoHAVflKiKPb
MkpelbmxvFNrdv0KKIU8jEIGENOAAg/klkUbIeIemDhoEQgC5ZEvyfmvg1L91/AW
dU6IHtFuCXytAZff7lsOCNAP/631io/o8bOvPgXCwia8Wf+Qp/6tvzVjqZVBFJC+
LoBuFvGQGiKHZqZYA+Xo82PrzNWC44nf0xJubdbfsHKLGWi6PxJCWnNlDAFOu20b
wBmFkZU/aQVW4vhjOtk8pPjjHrASqRbG7R1Zd4+9S1Q0YmmjU24hJ3CfFMbGtcNc
/YvDs2TLXqzLgM9Oxqo+XX76EJ0R/Qi2if+p3EyjO0uJHyJ4FbbVWKtGcVTY22XI
F1FO/4WB9QBgfYWog1Ln6sP0Zso/1qSa637rPllFJa3KsdEbVaUCiuhplff0qB9y
l4gyKZSm2DYUsQAkOjxUYeQgfHhv4GHsP732oh49puOOFVWCPsekHu4u64whZUC/
0ba+aj3bBYfrikhUe89mEcUAp1ZVI1Dbmc8RzSZwWPrWxoDhR0pD8xhbGsJEVTaP
4Oh7STSkuJymIyBKpMRFL4gJQUAiYw63niwwHoxgplxFUQkteMhvb+SxJmXWNp4D
5xMg+ZgXXxqjDoxbC22it3WCgYWABSgjDb/StlkLVtcsLoBdM4h6KyIbKFbUJbsn
fpT3GbBaV3lLTr4bnNn5Fabkc6KEtCzRPg6V1jqvVBHvpHKizocP6sM6oPgrk5pA
g+V0mShvvWGGjy7EF+Lo4kKgUmximbRWe6yDBQjXf85Jx53jbBc2T7QetHvHweLa
P1SWxllq52qs3/JdX/Y3K3fT8njJkUMPEhsbsQthn934JMPKPLEGHHBwU0VrBSjG
fgkIu0W15DDAwMYQAQc58YTrfB8CzDjKAW3dSYQFP87+pZL3qdQVnTdMDqDwC+x+
w0I76NTQ4Pkt8NdVM9UQY9ch57f4qDsMzmq1F51xeonrhhuGvR7488rjmJC1vIa8
PdclbrPvqCtJQ5kWX0ENK2GwtUoAA0MQn2UWJuKrTCop02qN3dnwp9IalaQUlTfu
afkkmbaOpo+gaHMB0zl55BDk1c/H2UUHbYS2VP9RpAkTGWFnxu/uagS/mXTwc2mg
2YqbPJNOqAPC/FaMcxmB+Wh2YV7CATEVCpNCSFmNcJvjaCQyQzwhJj+GB3KFBj1G
Ua36vShx5FO0Spuz4jJm29eKddKBmXXGMzXBgsfzDfMYpiFNQUSIHz8jL10IQrXj
Ur/JHSKLCHysEVmjdotyC5UlZiwngkCdy6/ssW1chyMyNtCGKIxzgXG5IStC/hX3
rfho+7G24GInH0B+vhfhX0UMvvpMLpQPEklFHGEe8eZSfukaizGLjmSUlDfWDTLt
mZy20T8sdlIwVqxMZp+CCLKLVrRtR4sPeh1+rg7sbS/og5rPr3gNOY40/KqfL/3N
wVjHrh2NGVmlelHzQY6/0pQ1UrHmqy77bs5htJJFSz9nVqJo8OQYoOeDYC1v4Ko5
otNTZBcs6O/YqblVItCI+EPXkN9B+9qV8KMcsZZXaPPGuwJ/d9x2v6WOK3YHi1zl
tNJUoZZzxO5UJFBh/NhIwcm+L/zrzcc2LmRzykvPl9S/nDY2PWvgRFTbc9vOlqZb
ZhZH/KNO8lim2XHNJ7H1H5eGV7waZ8ywCnTlEwTY5KxfH3+mMUuY5tf0JkUMXaAY
8PFi0r+xCHrdwSouUG1AIcT0eNvsi7XEVxJMW/m0JR5uh6NiV/lh2ZDOq0NP+I8Y
TvLXFiIa573PKutk0/zyULCEFicL9xNDSeo3Z0Q7NLbDr2d5EeUmSi2Jde4B1uad
PiRY2NAEtamtXHVi8QAl2f5YphLwXwUZVrW6M6X8gLiLaq+96kM97xz3APCSZxL/
cNIaFJBvxKNJzt9O+U+gbstUy14//K3i6qErbZ9BUqlY5RdExwpJQwcp2h3JcI1X
lIcM3FchVbVnro3xY3NCIkAQELKU2pc22kbvi6/21CGb2bK//xX5z6EKcuOAvTxP
I8VaYqOn6MiuuMTVj3z1J+Pw5+05su8VMnSH0AilUybKi72UPKuT9ygH8S0JaNMO
YzQqe2s5klhqiWL1854GFDFc+y8dfav9jd/UtaaZrzL1Rr68qCOcYVmLHLNRkW1m
ynwXCwLeVMtIxRvIgLbKYNNpjCVGcfoUZtSLaKO1goGD1Bd4abK59wb/W/bQfsA3
ZQYpCw6ede3Fz7GnCsn2VtOc/f1yUpGUZbrVzHubPNYlLGYcH5gkUqaz2ImPzfuC
rog3ZSUb8XI4x6VFAX/TCsFzUetHKw/Eky7cEooFAPUYdVjdsUc18EFJS06HHev4
iar80/9e6N8CLTZrMblUmcnAQWg9jblHWtpcIZV+BR5i9EowlznsDIegrqkEnByt
uA7O0AY3zlY58abaTvqfNDbfRBqrO4YRp5tNyX52573ovKMA1mg24/rB11gApC8n
C//DtbrTT27UlbED9xepIXnmGYLKvmTmWyBOP/NlU3mDJvPnzaumEmu8Q6wWJv8K
c64WgcVa3/HSLqC7fVPbvsjFKgLM7+/w1GaUt59noU1vFcFevm7NMtdLcbPXSciD
VDOWVIpsRb+YJwUBBMup2Y9AnVLUBo8l3blkTGBUbaSN8YkCpt0upy5qGfB0QBLL
RuAX8jBDTXpHiogtfmRlPjy1fs9KQ8Lr/t8riNNVWz/g4656yiujGXJDrts7qvmY
4IeLITYhT0292T0NwWmaFE9MyVKABnWWPNVzCydmeFiVcGe2KpZYc2EgDHxOExe9
rOoX3KhHAZaiotr8+7o9oNBbrTLQ1GkhQ/IS4J3UxleiAiAWmLYKg3BqECUunA/d
RrYcvMP/pS6fTFanouMdeJqJsVT9d80YGbJASaLr/XN/oKd40gxBaj7JABT58Hmy
DQ/89O0IyXjUgeZYSIqNytbzXwcAtr+BoPYnX1PxryYNZ706wZHqyHwqmIaRHuxT
xP9ACUqxJkPW25LUb7y09FojGCHwn7KHqLWtMzxMDcf6mgniSFgKE+gQh5yTaYxt
AnC6VVb6VSsWlf3alnrS31vAhTQ95eh4u5UvZyVQ2UzE8gF9z/4Fb77ps+o0t0Q4
GPXSQJr05d8WIhPo0LnZd+C8RXClqQ8CFQlU44KsfRmRsu/LV+MOelBs/Q5Q5y4S
rWcGd+sRh2pYlL0jpEpSAsLtiCT8IPxq7KV0cbYmpkM5RCXgUsIQsRcYKjXg+6ix
`protect END_PROTECTED
