`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pT3JN74qG1dak4mUJ+WuqeIQ9f/O4FcxBuooIDES22jfJf6Rn4SPdx6uXXuMM5Xu
jB2MzGEPygm4Ewo8RQAWQch3P7EoR6jf1OFUX6A9sRfc0tJUvek7b4eZIM99A0eb
WDEhrJqNCrKjhNz11PxHczj9Bn0sL9BEEGQBW2gvu4ku8xYrafZ6r9tpAGIOepcr
Gd+JHldUmIT4JzGP0+9ak1sdUTLn4gwOXvOAk/xcvOl3qN4MQ8qKWT8r03BUhLxe
7cA2iYJ5G1fnPJGMCWiPq3bBz6rdXuHkHLPgQ/LFLsCRiQOkW+o8ancKNzBWKebV
0Y6WdYhsfHqBxNCnbzd6jVX7V3WvWf1zOm4tVF5AtsV0hMZGpV7qjfuxaPKD/ziX
A1rFuZMDvrW/ZA0f0dFwJdF7v0AnIFR9lr3raLBSKywxxyoJ8o4FRNoYhnj1YbrG
WXE5eZDOLt+n2OTQXUJQz7YVr92ZFTwBmjJ12IKJ5HBnKy/ih/FMRKwD0nqGQnJl
jNUlVxMIWjSHtXwmiQwhi8rpDkH7mluttle/Xx8+Tni3oxXvqvxRsilDNgSRHxRY
XEBpWESGtV5kQPGdiZkjwwPHPHQgi/BdCwkVEtQMQwTPOdLCTddagJMOwFTRLwag
C+aSF8uWxTDn9Is1rYXG3XIBCy4EnKHFHOo2X5QMZOneTBy9OSDkm6YrjJSg+yiO
0nVE02Yulj/rYlw/NLo2A4iWVqtMqlfhM9tKk7sECt1qGpIjMW+5kYXQJ0TAmyzi
QIokEvGUCE7x6++5guT6ucb26I0QtlMnVvx+dF2g6q2CcQIgMOkoQfxnw5erITUe
lF8WojltkSX+M7zWP1OE1j6CSZj8fv2h3lYzliETLjIRS7sXlp3J52alSXQ8GeHG
jZj2r4FB8ZDv6Vfw71az6sfbK0awy04riIIyIriJRUFvvxgfhhC4nO25hMfAKWsK
OLQgIKqtHPuvBPT7zaqFznzr0Vjk6nwFp6xw2k7RuRKdu9Cu8ysdbKqZwGA49DO8
aKFlptiANOZNfthQ22W5AA==
`protect END_PROTECTED
