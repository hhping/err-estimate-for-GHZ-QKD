`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YhHBUm19Gkv79NQ0gV1mhSXZExSKUCRwxLZCK5N+Sj3tZf8kbwlrfAmce76B4u3P
wFTJ8D+ulpOgqR4+qdTCOwk6UclWtrO7/l3RF3pa3sYtU9dTI9BM4lF/V9uHWb4c
9DFfE4bOA5EjZ7r1C9zVC9MfENTUUBJ07Fl9OfltxfS+jqMTbItyJQ6IV2hUHXLM
Qc8164ua70uiYfYrPdPllK25xWlkUUebXiY+p8IG5QBftZ5eCFzhbuu2Z4JBdvum
oNkRNPOTUxP9JDOjK0c+D03Kuqd9xkour42F+jKNwx+0Z9WuMiBvp73VYOChW8Z9
jVXJQNtHAJvqiLE6y/X8OBeqlfDV5BstJ+DanEcH8fRf8mVhHbWCSofhgjSRmHpj
rQUoxTpOR38TJ3ZXSl39aZLVXS8V5qky1CKRKHWU6oZptOafJ7MH7C2BhaZTePcO
b8pVS4gMUVTqfgz4r/GxHDx5v1UdUhGnhx/y+oef7tv0/dUU7DOrH9WsolPvXDWr
R7YBvOVXUBBe5vKjHucPryUszHEaaqwxOwawmzoqeQ0CE359wVZMqGYJVha0WqP/
gDtDyFe9309Qo0A39cEBeGAJuXqj/m1scpJePtsElbKelo8qMdPcjS2o43h3v7Br
We+f05aONSmH3WNOWxqJEYOeMUzqW0YfnMDZ4wV9iamuknBSUqONEbC4Eh7fCffn
Ojkby47Vm5P4vt6AtT6G2Mc/w4gjkKMDDhYgZt9MUSwXoitep1Ok/yuMzPEH4Gg8
wcrZc+4ist3MQuWrdEAcZZDHthPOWaUr8QqOnomtLEedOw/6RuEWASJ4a1zjmApR
UXYqyU7dLNd81hsxU/2jbw==
`protect END_PROTECTED
