`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cq3QQ3RQnbglZjzuERce+81fAZBuqhwXhbaKwgLyWKtxn03FFtigglqGJMl7thT8
lRv0MqRfKj7zqbAcx2EB8vBCHu2OKsMyFEb6dkk6R35aKUxQfMw9b4dj7AeDdBNT
oNyqM+pvadM+9eEzRhsYs1xXJvQcbMe4zUrWDRU2xMjV4lgGZ48QmZIP1tE6S9iU
FyMwWjL9KLi948zABN3Mc3LbPugb6rgk7A8Ed2ynNxE/SuJIBeWjEb0vt3NSd3Hx
ac2bhk4IKm2U64Dqmk8Sx2e5nCxJ9oILvYUMbm3sPdB9f7hKIA8+pKJZWV9NHOLt
4YX44QnJDuqG4Yh06icZy7iR1vUp8PdyQBqsKx8crMdWFHQB+RYRywDmwUXDWeqb
VUgrztafVpDjJ0tsDZO5NPCO1VgQXlD8/RbfufsA9+1so7cKYmN/nxAUezuqM6jI
PxTLXweG6vZ8hEtdtJNwZqnoRF2uTjuYinY7s6nDiJSR/iVRsBFhDyJbfG11h/Z7
LzssC978klYXNRr9SdPaouoNB++jIIYkIR2yAvU3L/ycW/xFIGU0Dc9rxewIxism
vmqiamDotf+N9lF4wJX/F+rlvjM1rP6aImisNucjMlpFElDRzD/yE2giB++o5P23
DJxLcV32l6gFwn5J5tL/SHcEyv1B17P4hAHBhlNiX7mcZD2EsNGHW1X2xJSfyEbl
tVmRP2n6PiFimqDmnA85B/Q6aR+VHUzMtGQQM+aBtWi/fvVKVTWn/WhVF35s8JtO
ZpCo7V1R76R3dlv/z5JYqnsKY42Uz5a8ixPUD5R+vDbbbGI3ChB1IzROX9B3YiWz
zyTqq77sCHy76z7g5oQe2u8CmB0L/oWdAnDWA5mkp8kw0NCkKPIXDFjq/+wdUquE
8o/vshbrJplb/B1hTrHovpkXkaCiqDsTWCcvddACVBziFyVMrw2nN0a6LaiXFgEt
kkTtCbtCtyMQw9Jttz+9ooFUJ3eiIANeHCB5jMka7cSOI3tgVLpe+jpIKJc0ej8n
ZHfnLD4phVlqt6EZUWhQcj4BQ2VL+2Vi3uCM6eanDubufkRQ7XpCvTEkqun4bEu0
RDDE7wuwPydgeBO+YhhpcVZxp439xgcb/9TeOPBmDOSsOZOwqayd7WHkPCVLXDLZ
8CGe9eR7WBqGMJo85y56uMSi2RR3vQld7PRlj5SaTQp/bx/o/vWUiJMPTE4e4Vuz
jC+4zOh2CTqrLdsKCO0T844joeJOwRSrHN4stlLKcItL7K+RkW3di0QhAnfk8c7M
cNiORPDw5WW+ls9mHpZxbwiNQpCUhAbZZjTtWOCzE9YuqgH495UJ7qagOR6en2Kh
mVxLPEf+Ui1B6Xt5DmK8n6CdMef1NjbSaJb034W/Sa/LgRQe48kIM9Ya/Mc/Kwba
ATVRvF6j+OTrNKIjywwuuJ6mPxvBq3Ed0tj8488FLh0SUs7AL5jCwu460vWyVvBB
47yXg5f7sjRh1Jbc9Z000q/CSI62a1g5sUMaCHqSW3t6lFMuKtbcM1Q1jRO/fpKs
p3af1S4iMT3YQlol5POCcGu60f1cmT5oyCsEbE8+nXLj4wSmdiUNDU5QS6gn03De
PjCSFJK8OAcnjqTyXkns4BEyWL+8moCyNTf7bUxgwW+kLQ8m11V+Qluc0riKoA07
mbUVC0EKGEbTrK9ElyAvxuLs9hFx9NO6Ywa/DaqrGEE6V20RgKdUOLZh2Tg8VOTh
rv8er1AhQdc9jxSCGj9dvA==
`protect END_PROTECTED
