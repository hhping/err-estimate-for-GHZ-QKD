`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+vHzl7x5Hc7E+MXXii8x7UqlfHta5y0zSkk6rG1z0smmBTmNj06IByIh+DrUCIQ
FCawqhBy85yExqH/8ofr5/0eiH0yXybDMrvlEASCPFFpXzc3D7MBLXiJxKmWQVCU
RLWQvZ/T4aM3Rq4Xl+7sFT2OWpHBSvj0SMumoYZcln+xAn/a16y5QLdcppOPPThw
1e12sgvO5XkaT9H5Xe8VzOWYifljH5YfQprZd+xBYLGzKs4wDrYSy+pBTZ6slAZ/
qtAPcLAKKhW9G+tkA0HisNuLNWsB2SjWLts7TAsu4nryE1Tzu/WDWvY+5j25DYrH
Uus7uijUaUiPl6yPHaN0uWnOl813AgofOUVD3NGVYm0shcwKegGXa+lIuzIU1jGp
m6YIkM7dO/81T6pyvyZvXcm9sAH+N+sOtEZuCGuZWs5Yz94VeNSNkPct3LU+gd7P
jUjCry1dll+CB9RWaDSuloW60upjU8GqI6KyMqIlXwPUrHdKiWAOJZJN4aVdOwIP
9eB2gn/19S5M02SgkWJpiifxGp/ncDK/Q1YXP0pg3qFlodHYdxTEO+Z/7rkP8jpt
N6cAF5HaJVp6ZX4ZX8FdnZDbZkiQPh3CcNnRSKhXBurRqPXhXJfTO8cBGrLTj62T
86r9F49hpWTE3dVNIOUmU+t3Gz1dbhWztqVVxUb2Cnu07jgMiNmTY4qtsa6B0VPm
ZpNrjMO0GmIJlMAhCjWyGSz1ULIuHhc/4wyZnc0GRThlD2QGuhdNa5hlJBTreMtW
QUnTirYfBKIGhgmrV324I23Md2nw5o78rynt4etMKdW4Fafv6elmTXAUsMSeIPDj
+p06N45D6dytoEL5V82MkqJw2pO8NFCrt5WuyuR9RHY+Vz0wvhi6F1mN7vPjjM4J
NxterDWmhlEjLDTh/DA9uh3iT2YCet38F0WMU/io9TObNC6PEIhd+7rt8LCLVrv3
5gLhwcRPuR1p9UlkGTRGVWG9aWi5/euwnkuVa4yC990uozLryb8J9/wKOydSNWuZ
Fo8h8P0jRwefJYg+jg5AA3PuRWHbN9odCFrDPuX/LWbg8Abw7931/Uz17uAl7kXS
w6x7LR3gF7upLdDFEjvopmTKdm3HRrvnyHGVhtB3Pz3oY4oz7xFucO2m2q0cNRP2
FUaD7OndUCijDayx+A0LSSq2dmKLCJQ+YUxvE2Q/qIpGyDP/KBLNEJ5a6fecK51S
JoZvkhiTQ88Di4wX7wiPsftzfeOxPk1legtLQ70Iv6LqqcPv7PU+2lkbr6p0cTSl
EwZsCeNBOfX8W1ZNCbyn3e1996dmPYmNgyFrDsn1oYWBb4Y6BJOvbOMzTekTnc9S
U/vMJx3kHptxlZiXJ2eiXCh+AlyYF9XVLEcXdp0Krdhw/SslV1rV/F1WxMCFZHuL
oB8pgy+8ljFzV4kQytJNtVoFrELh8puhL1fb7LZzjmIo3UKY2Q68vQBtkcHnOpJh
Ze/uMRnVG+J511vBhju79F8kYI5QHmqSPiwp1oPbDe3kKFhnhRIBTdzp8InNW8ka
+6X3ZWBhcBTYMoBn7zibQGpnxzExjDVQFk9V6GYF+IHbMrm5u6yEQ8d7QHMxUDjy
aus6QKnkOt3Kxf+XfiwMAAAjfikqXoYvB9CJOlUOgky2AU63vxb13NvM/Z6fAjAl
pMMj1SAqNlofcUi07sqAgCcHjGOJyFHP7RH4xQcEBQY8+MUUJGdh+M/vxRG4MS3+
hFCaXrIofugzvWy4pfoKwC8hM94lFyvQaMwi0/ZJkvvPVsMrAjP1V3+6WEoW27er
ahS0ERlF3Rd9hZCs8flvE7ovbwgzUnBUUsVsCniCR+aG3BcWZU3eiqx6eb5wH5sK
r0OcmYYzLOM2r+FcvTXC9KbLv6JKuSESFvX8jdWHV+Z42CU3X/+31wK/twu3gwio
uNPgxFbdqwSYb+jlASL/WbUf4fFX8Jm+6JXzxoTjGd+yt1dYHzzJ9sNir4cYRz+t
jkdv54+oyKJ6YrfE89rhtoEAe6pzrvQCPggOLEYU5dZCGD2z3EB1zqwlTcSNP8e4
bfxbmDuvBjJdNF8+F39ohwifzTOgSbGSC8YxgF5JqjofdYTRNQ81S1BYH+JB5u2q
l0Q7YorUc73xLcIQbTV1hUyh0mpe9ijoNJmCc2/tNF30l725wzYXsXStCihMT9N/
6JrfklaI4efjE6d4YtpgnDsyMEGdLV/vP1pxsmJKzeMBodzNMvwSsky+LilQRsmb
RkavN7/aJYF9Fw38lnxJija+A7ty51dnnHHqLiV3ukZGMsgJ4xONIk1Ivbs8c4OV
3FYq/SdUfTiwwg+6RJ5KDzRV3O+Yj7+FBIl587l000qp2B5EypTiUa7JBHyXeOW6
omhk7lTnsCjntNGSqZLwtYx0pYQNXewlbfbiVmD1RQb3ot4cJng7+bXr+sQJfMWb
4BmIGOK7nlLfMdmf70mNaPS+uUpCaokw4urRgirMqPcH+apsmwvCsrlaYPJjIvf1
lFyC2sMfENYo/T3Q3hhU5cEYEQOeeoXsroZtGvrGp6gyK4/EgO6KRrB+VkxU6Bd+
DCBygyM7V5b8ryRTEUwXKYkEJqeNCZTubqHeevPUBXeSz9cUeAUvT/BaZH8Ajn9R
aXjkSB6UWxr+NcNEfekvcn5y+qa7/Bkf/oTxySK7LSn3P/YBx5F9GU4gboa17Y8x
MY3rUMLA379aRrwYLeZis8+IbUng/eAAxivwYnSZI8ozDIPGkQOei4m+sZJluhfj
TNSR2cfSiazkjb2dd3p0/8zp0r1/ZY7GntnFMpTs8i5/v5SBhM6mWQ8nIok/iqBH
YWvQLRlYOD6SuMjmeNirmf8Ry2jsHlpUnRInPnDeeJsnfeCtKMEliss2w7tqeBKP
NoFJp6LI4yMXcKrTDSvWHSTGy39AMd3ffnHRXZ+5WClj+O0KoDnPIYO/PyVRN6AK
mR2eWhgxGwkQKJ3c7sPI25id//F/tlKwQ8eak+8jE0AhX0OVBOadOxA4OGN5y5lj
ePe8khBWVbjLP/pk4XW1w7R74bcxg4jj+VhHuUEpE33qJsTyaB62P7kgL/+ZqVBz
rftQIXrBFoHlkcONd6L2B89PI7WLGibHqQtl2EhiycPuXu7Es5Mn5m9bqDBbXCND
L+dJ3r4mulzsE45NVCy1/klsCio1DcdFtK+sAEJwb6l/EZJwJCSddFlKpeL9SVCP
EJ+8ikjlViGcexrl9dlmHTj9nx60RTW0hY5kumVN7zWNtUrScNuMOfq2R8AIPilj
KVuMVDnl5L50ySUKIDdQ5lwy8pjoMhxt+T4SXdayXxc=
`protect END_PROTECTED
