`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mysweCzzbp6wu1j6NEZ4n2On9dKPRHmO6K65O8RO3HCH6nGgjmd57+yKO3twMgnR
0dfJZ7XBccxUDnafbwSHVhZ4QBKnqa1hv0juElKXU0zUm3BIyLEDOiFsb6VMbCaz
hMiIr0LuCXp4bcvdK6cwIpM6gvHYAbGZnXavwAexxMSucx0ny1lw7B56vpky6Fpr
hicnUu/4bj4XzGffF/g+pYz2qFrRQeM4Js3cTqhCvnhhN59ppHDbKf3r0fn87xD2
RXeyE35DVxWFQBW3UJYFQradOBlqOqM7hCJu0C4SpDCOMOHogZa6oMmc3r77Cn2x
0Qn0Vr3RdiywDZ3jeIslDexybjldPPvR5pKIc9Yxu2p/30JsM+gz/z12mJBHJGb1
9KPhuB3+cKdMDRlSYE6CaOfHRhbO32JswZIqi6Una1da1DdkZVUha9FcXAwWs29H
uDjmiu2KJ4xVqdx5xouHBJV1OQGoq7fzYZ+NtxMWBzTXJ4DxcMxxS5eS4r3CVRYe
EW7Jv/iKBo1uJVGicINauM+qAGlX7zHXEZMElSsxZ27T1N8HLWaluQt7F1Ie7bCb
BcDBE2ouPvcSjPnu5MVwno5/IPpx3HaTkSMXHJYNAaTz0T0uImLk7iApa9mVH+hB
xPzeI3quX++tzXnWBqUvdwlB0u7Lmqp8F0UlkJzdfKG1Ss/FbVQm3ZJSMQKmHxKd
fxmzim+9soLYZdItTGXjbSWd4wAc/++JRtGZJh2/rx/4cyGDKn5FiMJ3zYOnF1wN
uUtyLm/R3k5+BlbOZq+oJgWEwTUMORFxCBPuC0KjrAVybQGxxhtjYV4u+IojEikK
UknRtTOE+NyCRGR73rKU0RN7FCGnc1LM2A5VTN0al5rSJSOrnUB8S9xQuvEedLKv
/j/7vrLAOPj3TeGSkXHFEemeXdqCRnMdYKBhLdkgEfIYSdBRKZbAA1/9bnuEzAId
Z84QJELmBvnq1Pixi8fwHq8H/VvTtXOzlBOXiUcBjZInw+qqxQxtMJc5pU6eRGpI
1J0AcIdnqvHucAUusv3yCIiXC+nVbJfoIJOhUHzIJfeWbagy5b7oIunRNB+3F00t
6t/e78a6OKenEKDIpCl6WzBBALGTHfnXGGPGZDymGI8mq0G2EM3GBN46L+aQk8ms
owrDG8Lz2auUGLlcgLKIAIe1Q6LaF4OMX2RIXQD6D6RQ+AbAchOk9q4sAomAgiGq
TkAixvsSXZK9zPfglfM/a/eGjPixuQvuXlPNl/VJRBZhmEvgbReyCal0wwCCjWkZ
xCzcB5Lrg7zSZpK64jEUUF8iahcYJr9eOdP+12XjtoiSMBk7Nr9TfA222H9x+eG4
bBcpnys9lbmAoQhfznMSpzoAv9J3IaOh9se6fGYhS49Y6LQLUpt9VR2TMW91bgM3
AUb+mFQTWxqOdXIeoq/z72HKL70z9gedGmOze5utvakrK9aK6gGfKF4EfL9RHcdy
TBzBf9GxYQW7bstYJK5pzulgAB0OPgKfhVDBQQ+1on7zIlCHFLeGOQpM7tBakf3v
ey6llWL5Vv8UiYXTuc/Dc26jF3pUCoOG5ETEcfYFCjy2rDzgXOSDu6pvo3DUPjzA
EdOEyjN1baXWr6dx/yhECAaOdGEM51f7S9HC+mWl6hdLw2ZCD+KXQd+U3nuWOgcK
WudDzRBbopo+LnicOOeccC2lEy/ItXjil21+2AJd19P+HJuQ0+KS+++J3qEU3d6R
5fWDafA4zSAVZIS09KD3MnvJ8fiiev6Hl4+5X9jkymycys9eheOUGnTzg4s+runK
83bc+3Hzvndc9PE2Kss9ebgms+ma/Dh0PM9SKPShzFDECFUG32UX9vIAWfznxs0P
wn5TywwappiGhS+NBb9EPhr34OnLzkI2VoYQc5GTfG64OnnQi6XKrnWnJNE4Ho1t
Ru7/hiAnkaec2cSHjN6ZSBSTf95XtbHIpjN+GvH9wXo=
`protect END_PROTECTED
