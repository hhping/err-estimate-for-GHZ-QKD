`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gD1K8+ZwLkQbivih1hb+C/xWcmXvtrQSrnXZKHTQjmmFZyyinpiTRGjWXNSwS/7G
byagO56PohdbtSx0jcS4WjAUHspF1N80i4sQ0QZcNKMZkEFoVSPKGWWFPcuarIms
gv0udGIQV0NIp9wEDetMzoOLP0hU3o7d46HaaBonDqVDo6OT8li0rFSGTOd5WRJG
lISaz6c+0zHZBjYqhX0xobUnOaBtUhD02J2nWMfo5QZcYrbLTZ0WdFulO4oNil2V
bv9UhOvz3aNemlMCFSI136eZ4bY9fxXfsMQz8tu0xT6EcbxjhFQdskF2vsO33nqF
EeOMNZbnNxTfOlcdIT5oI311rKknCstxNk9x/EIk+uypFkcL+P5MGbOByI7hmIaX
pNoDGk7E4VU76ZnW8ZnJ0ejg3vkXP+jU4KGA8+6KHkDONz50MwnIL5s76K0gnOnR
/J97D4HFrRVKEMJmBVwwm0QxXwueeftnF1+cHZe6sKpLsEdp91a2GF3vcsdEaSTh
wyQIUbefAdoGh68MZvqWTD2DH+J1Ki2IUMFSx95L++85Q1n1j4C3RYNk6YCZzS/Z
V1HAZBIE0ZVLLM6oNPfgtQoatz5ffvifIGyu3E+aFGUP5OStbCDGJ5mntU+xS4DT
xFnDe+PFD9xZAEh1UoFswzJX7VpsCCWmNJrBQ5desmEWe8o0KXUSGgYiTDLPAwY9
6kovLu3LPPQ11jyzuNKxt5g73bTUmDAY8jX4X/L+Rl+wuFOJ2vGHIo5UkRF3CMWS
HB1mzeZ1IjqlLrzaKicwox4jYhLg5NE234GSDI+6OarWCZ8OcxOOn4xJsPswFwC2
+gKa7olqVFX836F2UhrkC/5CklGetNc0lMFhp83pjUZAo5aEVlSeGNyh2hzZE6HV
YKmTn05phY5smxDrs2nz98bhVI1BgZIikW1PiaN96ps=
`protect END_PROTECTED
