`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WL5jN5/QUHfQMleEFq+1sdDGvI4e4G2pFKxN0hBdNKt49irXckX2ccL3i+SDzem2
+Iy/nxYBcN6v/YSKrdJKKZFsT2EGDeQngwbzzFAHEp+sfClsfYMKhntnvQ790Mvv
mSM718lIqlAP2PAXGsTcvWgEMV4nUEjjX/0SYwqGHUf1USakYEXR5/uBcuf+iDYn
QJRwgLNf2FLU/+MlZPDomv4rHh8G7xt1iFQyBtQHzYSktz6yJ/5j9YKDNSsapGnX
qqVLy+uFddPly3DTTpeU+xHHHlGsX4hObUB9+/IO8BFWiIYhiOrEaVdoweoCTeCZ
tGR7e9DJhk7b10LyVRByYEoXTw1MoDSH/VYLNd/Fp+AYfVaXZyhU+h+qzVWcK3ml
yGTCdEkWHqp+058sBX0VSOzvGDupFs1DmvlxxgaFYaaK3qaV3vzxxKc+O79fDMGH
L3NCdm0mertmwnGGssUyQvsvrx26KdQu8MUWjRsKr4K1woi1FIFMd4g9ouWenJMw
Wyj/PHBeTB3eYeIFu8O8yrmEQc9UcoRweXKSfw2eodiurp8G1ZfBP26m4uQYoyde
0LJT5VhLB/a02tFim544eYDGgzsRBCg/1QbxPtlOp3HxwOvvm0MB3HaSKWhrlMqJ
aEzFTSQ/hFGeAdD/eU/NjzjfeCbOYjD8sXsMSYgbJ/inf3KDJii6SUV/xygjuWEc
e6/xdCk/HP+K7+7D474RT3DMaTX0wyU/ceNhCPIO79mngc1iIUDaySvQCMqXmmTw
sVecKLo7LMnXuM1Uozollh2SlMsy6VHcVETCe3YjOiEBQlalmDxi/2i/y15UyHJz
hFCbtZ4CvEjKn6+6iLBrtogx1VcY4rIEwuvqGPOq0Jth4WP3Ff4hfwG4pWNn8Mjo
jKKaBOs2b9EaVIH1DzzRtiEujOqSCvlMIznJVheOHL4v95YCj+MtLWRs1PEHtMvk
uSs2fRqJeMV/+UzhDP5R2q+jH8uscF9BGy1sbWae7yljFrWwj4/WW9BA/Ga3jSqi
2Jn7k+PjFUHC0a387w8EeI72EJzDqjyEBL1lZKZxVlxWCgNClpmE7dqgzlyYYXYX
eKpFgx+G2e5DH6oQ+8p/qnQmJh7QhvEH2+aPBuOSL720WJvdIaBEdZimbWfcvm63
HbfOIhgA9xhuOU19suPQLnWtK/icX2dypug/+E1FbpMlUELX+0Ch3yMPeUUvH/4u
Hq9Rx1JxyXF4ZryqO/4zC7TbIKTMJyN+s1Ty1z3wUj384LBea8yWZMa8kIzZlGZD
Ip66URVv0u1gaOyI6HKisaqgzCYKW1u7kO02ztEpLuaQYkZdxfgN9xZHrm2/34RZ
+QCa8AOK1+AohIr//btLaMnWUwWJnCL3QW0ZW92CG0m7lMsIP14Q3ZJpPUf4+wgX
NNvNZqzIJqG+d3hiv7b5iznLXSW8XDc16O4tsVypCiK6Y/cfDl3sLjrviQJLigrN
lPb+1J34StFG5XnlbTKt/iFk3FqMqZ5czwbPeRAArnHLw2vViqSUbsGy794ntNJU
z5nejbEKYFkD4UpWHM2W7rPwvQZ7ohfy1KeuIhBk4YQ/Zh/X5dDnmbdHbFYIewUH
LtwQjr14eV3TcKb2L2zEC99MWANX9htLkr7eyUMdRYU/cjWVNS2w8pOek7mEB8F8
9SsTaTtjOO2/a2FZUuCgKrDqwxUvv4MwCyMhUBFZg90=
`protect END_PROTECTED
