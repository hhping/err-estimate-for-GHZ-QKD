`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADvtl5YL+QiTXPCNyLkRrXnVEWYmsOHKbejlsimjtLBlGcX0AseXpoUl1RFCeSuu
SCAQnz45ZALovwy6ESbpJJUsjin+FfA1dCwyf1WsgNYV89wqXbkpx1c3n3m/uZu3
BLwXUygyFtHUxvzcFm98w0aqcvcpe6DJvGg7GnQ/rHB5HkRkPbdDpPhxsq2IZfaL
sqPDjE661bwr+Bc1mIM6homiOexQ/qK5WZ6qqbUkggco/gkXJt6XnW/MadQw4Zbo
K4DrFlb91oqJih0FSHvYJbB183XJOswDSQrwGqxQarUwEVUJLdAQh1yGKDjHLMZP
geTcaGvrJdtnmb+PCy3IKsZnRdJyM4DU6RlI6GsIkLgGWpV3zfisV2MgThVXSFJM
rRDpmSjNEsmrFhq7EPLvfsS3YSulbwHV8bLdokTv+kbLGOY3BslL++k1MCtIZTXW
FTGYWmfbUeocPfulr74OcKthLXEDnVNL/UYBLMxACGYS7px2hfoW4oSImfpwfbf3
SEBpraOS2xYO0iTh+wR9cu8wJ4/RrcDVUK4Oea4iRUrccOMqa5EltzIvt8ZurJNW
NZJbhs32YRThiXhvHEClORMcunJPDG0QoW2bv2naguQAuymiG76OA+FQ/6sOCsIf
n3GiroyYR+HO+CvjxlKsZtngB0PsWxDFYod9RxuVpitkUi8vLt/4fzcdUwH7r6aI
Pbe6azlTu85+/wnG61DSlnt8yeKkTTqCpN5t/2iVKXDt7jKBp4FUDMWpOb3xS6o5
N3nszUpu1ctNjgAKjuMe+tJ/AwVUneKa5n82nD8kODX7QtqO8PXo26M1H/RThEb4
oRAm+VGUnCN1E0mxBaGxZE9veQaWZV+2e7kMlhA84Et3yDGe+ZI3eFKdw1nlsREJ
+Zu+UKs1vs0xHwv6mTQkxaBVubq2vK4KXl0DaO7QBNuFO3SKcp/DlKT+p7JZNydY
8Vo2TDSAbyEPdnw4+a6Qz7hPjiNt78ChlGgHbgXbYC56J02w9RJchEYD4vYDAcOO
OFM/biymzdc5lz2OA8OyzgDbSv097EcoyV96m+uxKXq61IYQtDV2y/y48Obd7lfY
XSDg/mcYCHsIgPX7GdJ3MAX0/GZ9Dj5vFdhhiIGrYu95ER+w3lbXtpRFlJ1dI30I
fnJHLZJqr9riHokd3jJb1mHFGBoE6rS2D9/ir8iAR1tHL1E95EGwH+2Ara8horDq
TF5y9l30+qzHBjjGVFqQlQtsIt6h1KtSrSJu9+htVNN9177KlDSFCeW+I0uCJqwu
ehJhbcTOBkuT0UikrEegO60rG5IkrLBXWO54bVPpjtfJ70qd64kmho/JRIOs2nJO
1ZvTGMaKWQsSEt6G3xNpmKUj/2pB60RL2MMLIwt1jxC35vuqnTXvTV/1+6khC7Ez
gY5UU2aG0dBUWv0T1gKYcJ8+kMZr7OCJ1+Sv6mGOXjoKMbqHwfCFmiwvW6EQXEx1
ec2KsEFMUZZG32qpV2n4KM4Qc3mdPjCJ6KcLTC1Sv8EGjfW3xdZq2vMzZMOJ/S6s
HsIw3wT1tNOf/7bBl4+n7t7UfUeAGhhSjGAyuxX96BPDLxCgZLn0OHILeOI5tUWG
A4EAad5Hlyn1TOBKClhB5yq9jH6UG4Dpds64+//ULgjUtAoBEmyxm29Mv8rj7nA7
p3fv4mqahdrUDrhePHa/XdNyaLKKOOr3vOKHJz0glaWWhExC/0Axsa1hS4+orJM7
SIzXbCH3ZEJfAPfxdVQKa8NjeiQrk/BkpseeQdEe96ep1iN+qRztSpH/gnN9GUf+
EYo9BbkmvQ6dWATrm6pzDwhlR1u/TyXdsSoSYyHPPWfsQFyCDmm7Ndw820ovy4jz
t/NXagxJPLbZVutG+S39PnMKP8KDwoe8VwW7OxPg8olcOGuD6rEtpig9mlWJ5z+J
qys5+hr2Dxu0+MQXrI/nGQ==
`protect END_PROTECTED
