`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gR6CegbYcErY+HhCkcymn2g+4ANySN3b9N9f+tkN93e1MzVQrORjlky9OIO2siTB
mdFRKd9iwWFt7SepHRf8w8FObzKG86FLr2ivSUB3pI7zh7j6kPQRpt/GGowvCRPp
EzHwSMLwZsZBJO0ySu9WDMgF95CG9aki1ZhOLHEEjPTlb9lwGe/VDydHDkt2/4YL
sE1hVcyWPypHrwN+viEQzR1ZkQIjxGLTUV0+cPa48SqZOrC27ejnSFfyWdfJS92O
jgGMPGY4MjCD9Qh/jOdv/DxZ9zJPxnN/esDpSQNNz8xenemJdbJpmksn85r3lCgm
/0NYECvEvnoCSAVlAOqH66FcTN1oiCvVQpkwRBzCNkOEYZdsHNoBsTR7AfmIoqpW
cjEJoJaIC6nArmAh3Ugc3uGslp4VRwWKmIq87npKoh/4gQDq9kbaUGldzX1F2UV9
SumJknf9ilKvGop2SkfPRx6KzE/aLis0ZGqLe7GGTEyC6STptd9hZa6vw9wPs8pJ
tY+3b9iWSwh2CV3v0+U8wm22Le/YHTooMAmLiw15Zk4XJ1Oi2homF427LsnPMeDv
ESzaCf6JQH+h5hVKn/vSiW4QdCxa8xW6nyOzCtYmSn4My8RFwlEZjNnSwtfNvYhy
jgH0xJ7OcosFAX1nPEBAR2LgGNolA3jeRoAG7ZlBpLhu3wgLixaXzwKSpppWkhZt
zwfNbU6dkSJBgR4tfsTA9ij6/+OQ0fB7LmVFud/R/rAgL0xJddmrWwcvZupAplUB
bjXujgVCXFjkBB2h9hi4j04PiIsmojMbPS2265LGd2JoiBoWFLFWAGXhD05NXwsc
zjt8q+MnH53W4x2M28ri9eErASC63zm4KfnEsrn1+1Iyvj64JNbQYrNC45CCP5d0
RGzyRdiu83KBeqkYswoSb/6ABfhuP/yVYy540k7e4U34yZUPvme4rjyiAPfczAVO
0OXrG+AxYJN0UyqAdwT/nN4irBnFxPo4+e4uBTTNcUasL9wnNGkgZOlaeyNfLiXV
aaUhDb5LWF00lhS8bxPw64EScmfN1Alsvs6hKxbKBhSaexoyfNlahCgGXrAzEMhO
j3t67KwEwbNkbucxKAadnt1EXJupaxIOwX/owrEAWk3VjarXbuOcJHd/YhNAooQZ
OsClhIgBN1ZS4kT+WOCu8PNHM2tN9PvzFmeajtqiKJ6GxgwW8Ko0JpqiCXuboTJS
TCD5hMZ335GzaS+EGN9dBeDPSVkDxCUhkaqJwWtC5kLyADJPMKxIrdpxnIkqB2rZ
Pa9iewKIOCxYRNSIpuPutjGUFHSpgZOWJ7pPhlW211st8PnwU7taN2kt1Ejoc3ry
WsW9goQpXHo4ytwrQZioBMbi8gIkdr5nTSLskHVrLytiMcxFGhnFGSJVhwC+MP8a
QThnJI8NPnTlVfRNS6XbbszD+DskWBSOzAeiiZcf/mwkeZyfv/UiFunShtiW3QsA
Y/iaeqAGGAvT4t/FZrLJi8LOakBk7iaL4GHZuiMexEby+9q9Ea+PyQvMfNT9PY3r
C7mOA10IX/dmT57JkW6z7g==
`protect END_PROTECTED
