`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvoNkOt88joaLtB1UyNfV/5mj0P3FwNC/B5/I6wgaEs6Tog7hCNBCX9T9yCzAOYm
b8H+MMktAm7bMW1jGdwD76X2MjwQa9HGfCYcryqcG7w1pKYXlGrspQrzeaeslWa+
R7vLiHZjnim5+rHqT5EiVOIhvvd7MezRv8qUrmA5yvuWkDByhgwifk96vNQAdS7K
5/Xg94lw0Hb4HFcOb66KdEZqgyyEN7HFWYwaKFPog2nuQK22reuPndLWoYKWf7mB
++nC+tT6TEIdXK+MFnBeJgNFVvnTrlKtxsfq/m+5AAIJLUYQQYXen4/GJSkSEJZN
JztJIR1Pcu+cpF5vjpP6entdRByphaKJrBgp6T/dS13/XRu3YmC59V8MxVrvO1nO
s9X7GLZj5XzXFfEJSnY8Dt5FC76Hxx7bkZVIwm90118q/ReN/qXGwilRj2rSq7sG
GKYWrw6fIpMykX8bW0hQYzPB0+ypmEwx9Cc6mYOptBSBsrQFfjGAkGUnUTavpT0A
zu+3290wk49yUUuYl09XI+7xId2JAUpWabl+a4g2bnI6e2oBNiRsBDJ7wINDLVAF
ui2ydrR1hFmbo63UtZJlwu4TugmUE1l85Q1MTtdsz3i5sgnYtD8psVXwJhRezeO3
xVUZEqvbR1otkXJghUR7hw==
`protect END_PROTECTED
