`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5Ro/5cKstfANerBffe+6fCyK6Xgof6CVV9BkIcBR3vuqDwLXNVKl0JfUtZJRMzA
McxBy6sAA3InStjGgPa5sbrmuKl+SWBlqbMmJEv5TCD00vzf0rv1e5uFOSiPOi+A
5IxpgKaGHvAEzjWwAKfevhMgC7JGvduIp3qn2JLkleVoQ/GjKRN9Ggbo1hKjY1F5
FaAjkgn7RttxYOxIcsNg8PRC9LbvgLDDxYriWqDETZPWrb54N6FRhGnMx+OT8JeA
TJbGMCQIXX9uY+r2H70LwmqSHjwMFDkvo3zqe6dANrFeuqwxw/WmuyS/7ZFlc6LC
pUMJUJh7dXyfp18JWqiPT3V1IfdfXID6KiVg2jCAVtVTa94HRBdRtOjZ046g7p2e
C0ZzQLzLScD6HqstFYMqQK0nGkDol8XLwn+v3T+csj8nv8yNarEY/up961Sffxuk
wrUmcxWpmrQqghvptiw1hvGfvB4pl4tBW3j3Eyu91ABgxZ01AgFNZLUuXcRCvloO
gPgy9YcN4ZlWZrkPdm4Q+5N/LzsfdkiAeu7wA0qQo7CrnFBdOH39f26Acs9HFkFz
vEvYknqspGDbT0An4hVARnrL2sOg1ppQDirQjPkHO6aTUsQSKKFwcIkxKpOpW4VW
h4OPn+1C+ZemAvg8cn4dNe1iqPV7Fo6/TdadzzfMWPUV77f0hLC6wVOn2h6dDgts
O7mKpgV/GPZ7nD40+TkKQu7hKv0LSp/83KcRZuWD0kxuRLmDNP+O2j3LlHUViKpe
yAYWz2Clm5eQAAB2+mwA5+uyqYpyyzWdmLKcJUJXEwkQ2t6UJTjSit5aQ858UU0/
5PRul5oHXEyYLCTeJaSq8Oatwen4oJA7DnjZzzxLC6uaCaerdYURDwNdz7cuYAHY
OJeVZLKYD+yH8+8SMUChEycwJdCgyCsEqVNGKj6WBDacAxawROS+fDzNsXoxfKrK
Yt/i8tpbsc4dkvtgUhlvcF3o7FimaP04jx5aNOB/u9p8cm8Yqvxsb7B7AQWNKbW6
SQQpQnRKb8A4xmv3kr/K3ApD0mPD+SV+Y1HlIsOW29cj+an8SjS6BzZjLh6PUML1
5MTww2/tV4NWJVz9OcGzNM/+UGVw3Xol1Hcz8uU2UdzwgVIv3ihY55a8yTX3Obuf
tD+C9vnepBl1k5ZiL4TcsyPuOo1aUYQQchgxmuBX9TxsFN/a/HDXjcLWA2eEGIp2
e8MfiOpzDNqKpZ07dhOHwQ1md0eB2mL7cBC214On/wQ=
`protect END_PROTECTED
