`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXe+rC+zSyjYLlMUK9LoikbXKW04IgdmcXRauv1Kzg2fpPHvPAOhUk3x1A0vD8IQ
Fv9ZdRPy+2rQEDqmYT7V0I8G55pnQs6NZp9f6cJnkcOHqrcQppBv2cvXdgIggLSW
WPUY7HK/timO8HjXOt2suZ1t3lbK3d9e3k+k90aZimgcFhY7Fey27Z3KrhuRDE1u
6Osibl8gaqXV7Q6b2cjpelNp4k18HMhSz0O4s+l+qWbIdg/qIvotd1ocjxNyaJ8f
6qleKTSRQTunjdh626IJ8uZnl664TJrwiZeXGd4GnUtPr9DRAOaH2ztC68MvPzJn
+5d/ajdfnQ8yFKe1XCIbUqgayF5oXcRqjVGP9XXbNvZDOJ8Pr3M6bHWwu0PyG9rZ
pUH/0mK3eFdMVt3E3QGgVYd2d7cmv9vq3AvYEaSrsTk=
`protect END_PROTECTED
