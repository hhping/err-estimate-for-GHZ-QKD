`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWD8L03UgOnuhrZbTEiOMqlwIFIiQKIhKVYPU5tK8rn+OdQJLx27Lgyi2pFbvJXk
Fy05TGD94yTaASKY0Opw+HqukR+fU+uxmXVs5NhL0N+U4kfu4yU7gsZPsyAj+ghr
8EiTAxzLe5Qvvxtx2BdgBs8+bXVgcP5essiLY8I3Da6AUfICfvA1l8qSfelE1D+Z
n7IK3UybDyimaLWqNb3HAWE8y/soG9zuDwAN/fL77m2Qc1IT1EtlQxoptdg3rUBZ
fLRTWM97aXcfGer0n+RzutgGrCbu0hOz7JeNad84ma5P268RQULTojKb0GpZ/kjw
cI4OOfICVNC0RgByG8ST5ylfdDKUXMNprJ8s2lylCg68aVkf8qm80+G/UfiUUSdd
CyT6JaRMgCWxxhNUwdXZrJqxbMBik8MXy8jP9GStMbmkDoirRzsMUw9FT7kY80Q3
u6lTRRYuxOU/CDWOnS2hrMNrYPm3ph7sBSKvVUqj2cKAc/IMnfQP3vOtknApL/06
XxW0EUXFX6wC3pE0lxBrEjG8G1nwVn1U3djZCEsOHlEDkt1uccdPsgVsk9G65jS1
bRlkfD2MU6ec6zBvGV470b5Qqbni/61TBKy76xAzaLNk+ZtVFgbcWMnbVNLSv14+
1WBD8gb98SJBvV1WsYU+pSKCZoNbUXi1Iv2VXjbJClvxASLH3uJMI30NbVlmUbHe
RRGjng15F1s8rZsqWnNj7MlQo2YL2PGm6ZinO2wA1hCFDtHC6Ch/opddgFb9eGSL
EetuLa/Kl6gJ7X5U8SxZatc++Kgyh6I38VcM2dEsDbbVWmWqMw8S9ESagMAMB8UR
sgBPUCgPm4cBcxTzYcYjKtRVAWKo2HDjQUOiiUM2ivZJI4/QqLUXCuS5N0rUTV9D
+z9jEAfN2bQXGevz6nya1Q==
`protect END_PROTECTED
