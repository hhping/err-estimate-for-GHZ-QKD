`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNNgYnFlJHbcd3JtLOSyQRJriMlWB7nMfiKqIwWR1SW4nGK0yR6zrpSnBr2ESIGl
jg5HtyxztCGhs/blBXj874umVmx27CnWL4qsAmr4kZSAL6YLXwY4pgoOwvq7jwP2
MON/eJ25aZhJUZgYIesVnH9yxlMX/wqQEq4PRp/J4cmHnY7YWkSQdm6UqcT1FLkx
S/i2ZTWqGdlP4PFWxxLQCNojXUl2HxqnKUpqbtj2OWsP4X9ZI+unZxVEbX11F+CT
kLnK+9nF1j7r59hiFzlRWjqeoC01vfJiSABb/LOkbz6tJCI4oXOE/7FVC+IZo5g7
jQyj6yLm8gShw0NVUaqYaEMISXXb9rPtpvnPF5ZBkgm91W82RbeZmrqaNaE4DRp8
5i7JtYBi1Bzzk/x7OyMqRUSwdjFUwil53mOdx1/9NeR3/boTp7S6UgEKg+PZH4Ip
5rxUkHtUJTVH+KwOtMYnBU/ysWo4BAjC9YLa7bzH24zCW284fs4NNqks6hQO+eSE
ymhF49jZezPej/Izd5iLZJWnpwpsXhOXBuGiyv7r91i2UBuOlZRCUPR+zdSFAkho
xcg07Shg4KOnSCh9eByooX2WcfWWn7nUkz1nWQTUvlYmW/rVr8rkOYSFcdWsgrSB
GuDpvADtLJlXDAGN5Umk55dR/0txcTrCedmhrP2p3k4miw0uDzIgTzZP6E3kTMcj
u7L0mU3UoPc1j+s0wiVYfAJh/Z6Te+vETo33QANKkdV11nOhbTtPR5IyuIXBThui
b/Y7mt6iWgmIM+wYL8aBorWMsZQJGDfzW1+ZdMmHcxmaA+XNcCvYojdiP6yFdhrQ
W/+feaCrELdPcooqeljNdsxVOFFayQLbex2qLGCOMzE=
`protect END_PROTECTED
