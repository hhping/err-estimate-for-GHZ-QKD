`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJsqP6NTlggyoyc169J3WiytXuJtlhNvFW7lMTELu4obyyV7NIigUGnhKj5MgtjR
X0jOqjb9/KtVIa+wn16+lpoFZuFlCHKjnSfiTGr8buOuh3jxhE5RKKC2U3WuuqvT
2XqszhM3wFVklYVsx1CW/48y5cVwh3Kp+b8/FSIh7Y8vsqCZO4GMiU6Mbu/jdqHv
+EK71F2ITg2cLla/GP/3XGLu5DsdVIWi+cvbjawJ9xz2j/cfsi3TG6wozt1eo3XI
/bbkhxm9Xxp9vPFjp75E4WD3sySUW0mkNGfWgxkR5gzllKb6KophhQyrAApGttr0
vatFcst7vpt1C6QnzEihQZgirFqMLegY6RtnJCtgQ/lImspQ9qDY2w+uGcr9Q3wu
9+2ZcoIH/0c3euAHIATZb09su+5AzbYrcfaWh156f0wYyBC7cmpg5kmHh5yCCL3y
sF4XiN5cjHVDKybHCJJsE7l0gBR6JOD/EMnjby56AcImNUG59d1NonsjnuV1w7oZ
ZJP1gQscbvsbtircntGMhU9wBHk7kiMjN6+tb69CQiheOrZcRkQFq+y3VUSigpjT
mwEm4qb5HTF6Ya5sFyfg2+xoIiklAprFvjHX/N5H18JxS2QckJK8K33DtbuW90FT
o1pRC/R8RPir+Cq75wivjN5p8fDp3zb21yEO8Jb00YFM0Ogcso5KO9MOj3uH32VS
8j3J6fXF3Fzqf8cEPk+pPH2nFYC3RcGrAt58Nd2pZF4PZQ7evOYphuktwu4ESirx
vTarXSFrhwShexgPNZyOyNIJnmttBAWeuK2kq7qvycOGKovg+0roIyQMtXyy7Y3+
2dG6egXhmPFf05TlSAx2lyQDPgicobKmylp93Ow4a9W3hWylo/tFUC0tSZg+gyPT
2ShfdcmRqp6+6N5/q3kJXDws/2AA8Dxi5DjbGC1BfA3Pd01qmH42K4vhvQlUWdXe
fGhrLuuYkaXl73MFo/bcS25vPeoiin8H9oLNknNNH++WWzcZRsCEQHh2ql48f4at
HYD6LFiDcBYeVeECrhUU0bqLUc/DDx1vGe+NkECB+EoDyu1Ghe2koz7owOsQsu+1
CeJM8ZjWmV0rgmeBPsuIal/Bd772+MdpQc19DlT2A+6JcVEbHm7aPRDQlNtVQOHy
qQZlZofMA7ev8ccC0Wn+a7TLUMDa9WFY/2Tdss15UDKGJO+NAFBfuzVVtiVPrakP
ESNxMjvDliD88AHs98lB6Y1BO52z/Xc9/soNY6qDmKT8A/94GaacbCUm0kKfgw7k
gpBEXymJci7DBC2IXFPhu1VqOy3HVsrLlEJ9tz/hSf3S6akB2VPWzLbVifXlDd+l
WitTzp+Fghlw6QhEv/n0ZLI+UyrFg50qvQPQ6LgnwzIxyWBPzcXc6/LNhO8P64S0
eAOk2+43Lyhxs4ELr8L2OJ2GMAwcspg7rYPHSo14MLWczX+fet2qgsZsajZsGGjt
8NtQpXMzdtR4u1cEYjpeVr6kA56Od0np+IdIC4FgDF6G9CXhZbxA1F4MaWwQO9jy
BimPaSCZXMTR+lXeC0FvG+k+xVYRJFp9ji539VRL2hvk3faAoGZQebHXSZ69uK9o
jFCzwgVCFOm3s1mjG8jGyPzR1D+/Vw4VW/u8IfPXV5LePvFEOz+lMIB7hzd149zd
mtVfJuiJ9PePeQa4Us22dH09ZBn2TNKacIIfA9VfFUj24QX6OVMmQMdeB/mfZKkj
fGzxSlmeN+OAdwoQIpjL6LznA6deG8pg1WYN6huZBcFMM5bCW68CmTdCVj0vbB7L
yafu6w+obFqiHO8pOOdXmPv0zSQn/fGYKP9GT/P9eUWmlEQfj9l6mQWC6X2SUu5o
diyUVTvkvGxov2Sq6F3MIvIgzTRYeGfYZE3zHcNqVCZX6zmEN+ryDy/5RGGfBIQ3
RU1lnnwe/SLNFw+ULC2Uvsi4vVH+kvpMoKa/3eHYuCqqGstwxjH5NAIjBl4EoWDR
2qM5wJBtFLdj1xC58Byyw3gLmb8tku/CRHb4xzoBmtZknnHZAqO13JYFYaXMl4gu
IAKxVGgUu8hJAg9R9FDO2BA7D41i7FiCJLVwbWfbhYxLO6dasuQik5g5YItz1kmR
zI6tnQ1t/sYTLCJmkabMr8Ms3b14JrYCXQ80O9QUjpwEhuYM75awp9AReGLaT8nx
qVTD5LQYWpZxVKDcQb9KKtjuE/qNMk3xC90WYuqHjNvG/icLggq9gDilDmj5FVrh
pp40NgiPAx33tbe3RyfG/v4GhcHXp0wUgHifWmWnWTsO0Zt8Cm0+uVrBhZq9H5iz
Vv73QjeuPG7rHz3cT+oDdHMAW0xnHi4MHIFCXp3v4wwsQhL69CGedskFW5qKLIeo
AVBjAOCkkOPDC4JFytCm4LCzjgtffqBmp6IXbOmx/jHwvQsdpMlNfb2qJanBqwvL
z7aZnoADyBBTyW5QrBCg1VkM0uv5iQJ86tHwEdFbz5+2vrKZ/yBZR3UEPSodCCVJ
DZsc0AUK8mWlOpwsERJGHRsXVDZSOzX239SZtMIpBVFgMYokUB3xLhIHEV7uCi2+
JvE8m598hqTyJcuVGmXhcg3Ejjtea/IaA+8+qi04Ybg46DuJSXNH7xTHm/rFYIRF
xIrHrqgGuXekydHWM0mBJuuZW6H4fyK42YzRrLVg7TBduLI0o3e290NC2FrgHMKp
rgNa6LVNj3sohvhkNDDXs06/mJ1iG64jRIbeWCNOIPaZO/jax+HoSwJ1w5qORHmR
rCsbcI7Ra2J9haWCfqWsJHQp2MCq/x6swPl4t7z6ItIUs+NoRtcXwkrj/Ep62q2G
DH4quCtD4r2C8uBe2jlb1IbKRREPzg5GmkAL8xQrRf9dIa/Z2LOTl7igAOwW+jU+
6iL2YxS6uYnTc/moGAKd/s4mhZ6t1eMeOO/8BbGfs6AxXq5rXFBrbh5Yda2fkEo3
Vgzs9xhqP2gQCoiyx88vwK0tonWR1EveMY9neo9WV5wp/UqICSsDDctDLi3ORBgv
U212WR0UhQgJRMOxCisEpA==
`protect END_PROTECTED
