`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fc5R4piR7hsF+QIagyNeRbCnaGEMA8JyO5tPH5zdE97eaom7NKC7vP9Tm9XvLu6g
Dd9PKgiasrKUilihlqJ9Z+b7VbrSAVxxfAVCLssf61b+tWRTC6/5QCs+7IGJ2VJm
YNs3ybT1zgJ9+UsvFKdfQQE7DFwUb30h0fcENeQ8c4u+NRp9xSkXpOpfYdGwQI0Q
SwdETPGU+3bXb/QehvMMTDvykMJlIBcJcRj7XePBfIeBSFRVM2SEkbj2SjV3kYGX
mYOdta0QGml4OQvWIDmyfV6mHuVGyCliFK4U3nrX8Gh1gQGL/dy73XDDxaBW3UVw
RhFPiMtRpVjjzvWa0dWkLspAjGwyEf8OUsInsg4oQ5vWBE3lpB+CAv1I0myv9UDd
kj0b5CfSVFZ5lnlszOfguuXpnSA0LMUO64B3Ys7333gFJ7e12mlbaEY43hBBrqXN
/AOol4wICnKEBk7ab1epAvE1jqoBwADemAi1FVZSqjsQ4fZDNiNuu6qcjh7P7xSz
o/qZMZlRDVPNLy7r+yzigq3eLBOsDlEC1w6X1V/ikLdXcnP3dDa2MFvhzbs5jfeT
UpvwbwSnIYB/ZeE4W8y5o+/quXqChSS0aDPWZtXaB3e0d9GMwubqdPaCvE6yvdq6
VPCn0gGTCPBkaw2hyNFe1RxxT+LMsA/PfuJ3WLCken016bOgt8NTOiksAnlFQi22
I7aSps+drEPYVpeVJLjXWw2iot5fvPHd78f7IaUo/8we8rmnNb6xX9S1SWZZXxwO
`protect END_PROTECTED
