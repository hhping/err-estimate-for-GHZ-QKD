`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JEPPMkmKjq+LOU2aTsD6z6fXmHAlzy5+NkPicUmpdZ5p2rHPOPjVDSI82wKMbZm0
sm0bMj2UeMCg6WQbM+37ZsbBqNtzwVcc8GPy+B+HQK5sxVdlyqDCux0LJ5KrmWfh
9Ylx+0B8o6IEWTh1wgtlCWX/mpjKQ3CuQBmoYgBYLPZ6ZywlFAk+HCy1+u0EiXha
2+kn1bfO/qI5aZgTTyAewTvigp1JoKYaZke8qbuEh2J83ODyZ5XvTTc9cufjD1Se
2gyT4mNSdTRv/w8K8tYP5an5AoxC5lp6FYmO+XqGNYOQOKUBG7cHOrGAPS8GjbXJ
bOQPJwIxHXqRbh1akHivC8TndxCQ3keRpyKehmI85N87tOK6NV4uZLw6q+HO7tSm
nWKd2PI1/KxXV2P+wFPpCDhKxYvlWsUmbvGqkBxdZaQIqoanzxTl/IOcOywan0po
VZiXgKO6ndVURk81hlaYEs/CV+gBwr/eVGfbkhleQIIEVodTqv5+LrCz+VtPk8mL
ku9yebAuvgX8OMJjOH3tPd3AvQIy71OJCPnScHcvhp5vG7uI1swwuAA5uJSiFVk9
OyKNRaHq92h6ul2EeI8peDdeEk2E7Aar9s1jKCVXAVcPXw8/hN4a+zZvlf9pP34w
nMCRK7npNOIGNI7rRPosfOfFKll6pRZY+vznx49snHocDjN8cAMNX8Vw58TCXP+O
p70Mu16JX7DMqmuZFn0r+EBdoyPCFmvBJRY/prfwMiJ7UQl8Ycgi3BOiu7w8clpy
xpx7G88FrUg6KQrAZCqylmbGzH9nP0S4SDWabtYDTHLnIIqI8KpjZb40WO6dyAqt
xesU2xRU32ubWdrNOLx9dV+LZVlzfWLhCbI7bJXfwfhzha+6b3UPgsTAi1rsNc2+
76sNP30XlckIOaI599zuDERKN6F+NvRGs9dFydjhBlaRHHcIZltms2Rs8GMcMwDY
55R8BmpJV43y4CC5RNg3gkUXk9HJvZTH4VLr/hB7vxY=
`protect END_PROTECTED
