`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sG49pdv/yNuHSTfV/127WnHb1IYptjTy9j/cRQvb55mcQal1UJsVNBv3fk3fxXJM
h7w2WpzoH9MVJyLUOQjuMj76Hbrteeo9AK09vSn87vTZXIvo9p5Enzpu1bHzlH3J
U+bwOwzIp7McPGQd45boY99B7TXayrUmmGwBTf982vvdaQ4riqEZcb6mG9wK5TZB
DdhAyQzX37WPINRpdew1GSjSN1f+sntYnupSt/Pd7gjuUDTWvv1kmEbeEyrlR3m8
eLHPA5YeTjFp8BsR4XSK5RuvUNsGkjwKdXtpxMBbP08r3/CJqqdadMu0GnWAvUYt
lbMyKTHozZgoLpevBepqoEGdZi9xunnlxw/Jsw6lbmC+kcC15z1BQFfc8Uf/MB4c
1Unb3Nemw/Ev7Sz+f8mDuGLo6A24WG6oS7em0S+wTZrVKJfeEUGoBNYWrbSjKwcN
tjp01wzolXdzK5vuuhb/zSuvSaTC3eYro0xE6RmNR0/YqgpUGYvB+KhuhrpF+Ihv
rm0EafQbLz/Ho/Oc6QSPCmFDxiTpS4acJiyfdrWYz3u4HoBFixN6nLjLf8lSQkt1
dZqlcGHmgNoZJPY6z0Vufqsb1EvlcgVA49pfUFHqUXHprdnrHSJ4Z1wqF+D3Jcyk
AgWCyipyk34IxnmPrqlgfqNmkgcbGMxnhl9xl8lVqPPt4kAIfiWqOlr0912ifin3
XoQ/Wv+9tizjL0TME8HJ6xYN029KDOJxPRzJ8YiS0KQk2hKRZpoYvBiiPOPCfiBX
AP0jT7AFRWGoeCCMsd7/fTSh6vKz+R/QXL1ArbdcIPXuWaJU4JEGDmy5t/nmZbQE
`protect END_PROTECTED
