`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/aTGlEvCN0MIyMGCfm82oVS+YmxC5867uufrUCUoMmcAWJOJQbPJnrKyd9F2I87
xlmF6T+R9GEVZKzD/qXaTSS4eWWcwfi0g/caZ7znJcYmxhVnhSJFC6OjsIrhnfJ/
DLd/Lf29+Stlvx2i7j2RGQnK/OF9xoM1cud5O+nwC7wcF2lZjphwGSpfw+ni3YIi
/70w/81JT91rhuLj9hfzGVDhPNHjpY1PHDeTH9Wrci1NzXeBwxH4bk38hWYkHjPi
SMC4Kr2ccvyaQyYIkb7Hh4lQcokQawG9UNk5lsZvUCVWz2LRJ8LxKHPuiFydJMBx
7od0SzFAo6T91HQZkkDTYylTYFJikavTmsN9ao/rcwq4KF2H5x3BMOm/AOmX7WQn
2Uc758MkDGHXvqdNq/WfGWCWxNlqy0DvHZIXMMAI8IL5l06EYsn9VDYk50w9+lvW
Se9sRKVzHzx/vknTjqMMRi1UBsUJjF9G4JQaCjIrWjNaXYOEwxC4Kl0b9lKZf0XC
LQqJK8I25p30R2Wadz6ODjVBS77LaRJcAs+ejQzKrz0wP7Nj5iZJoZ5vTmvsSdD8
WzQCBgeWmYdHtvJhoyu55uG9I+p5QLjSNRgwuUbdMSZVmHXfazgDG9h8/2uwjzde
L/ObkbN0kR5NK8FE4fPWRvY7GluLfXp14CEJFnWpeIwUZ/jV8P2Nt69Xn0MLSlfR
mMGu/iB7FbZU7zrt0joHGKzpap2xykKLjvrn1yonvpUdSVaPH0Z2nR+M8QSSthVX
gtdTeaodcYLs5BSSi+ZoOwlLTR9cm+VsiawgMr9tQhQOG2+1GHlQlwEnDGxyMGfY
iKB8AbQnt+aA+dfjlS97lbyjqk5ADoc/16Ca4cfqewF4SwvXXVj5JSsuWE1Q1WDG
xRLA4wXLxq5CceIVHmRgRxMSVwQ1yGPBHXh05yGVR22TckCcT2DMIC4zrHY9HfJM
CzOQkGvfN6pRmuhT8Gsf8cBZYdY38HT8BI2sdx7PwfyQCuOvaejn1dVtNQHk0PcU
d4KQ7gWnDk+sl9t8NCi4Z9Sa1ebmFDJQPxJWgRIufr8lZy4TdUkfoS70mNc/RjhX
MCESbHl3oEi1KcyiSM71z4owKggvpb6HJpIEFW5C1fJ9rgNF5SfoBG9XZHMPUDyc
IYbhhYThq+q8fZOtrMswP8ZV6515Ps1wO+jSAWkKY5EC8nsl1mE9BSmCal0LzlGY
7N+ykJWC+wBwwyZceK6x/RccZmxz/AJ1QjaJuHGBpIDqG0Mp78BkCnMd1P0tNuSf
+WuW3Q1IXsPB3pLkVfD9rJytL8eczD5UpC/8QMszHyvCq7ars5Xh33Irkxi6cYWA
3Zs7J/gxyoATMWsWDFit0W1vL/8PdHRNx1JAVfAAtzl4nFXCgIMw59lbSJwElYSx
og/lV2qSFZLHXRxSwAkfWBwVDH+qLPAcsIs8n6ZYf0c=
`protect END_PROTECTED
