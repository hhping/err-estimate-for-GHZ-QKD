`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcDkOtUZXI3dHft0flu2bjrZ5iNEzS7owSh+yxPp7qKvTWsaVS/u3iicCohrJo4l
1dSrnZA7nG7sWDcwWYicoaGR0Si2+ogNdJUwjMmUbMHv0djAIRP4G41tTXcZV9hZ
6DXTlNHfT7EI2uTC6bo6RUrB6dvgxjSYTPN3d2Omxz6cjpqleNGHNHPIL4o9mS52
jz2+AWsE0P8RMqdJzOtjbzoffLuxW1+7N405T+AStDboeETw3J1Wt0Mid0rt0mIa
mm42S/DeiH4+ncTBBDCr34Gnk6Upspf5D7CGYw19eYMNMBIVggIdkRbFegXz+GCz
Jyj1ZYGtuWzdF+yaMPL59nPy1Jnwq7zzrfkn30iTNzPCXyLQMZm0UKqGSEBRjJ7O
J3OVQPFdwvRkvbYL4bLQ/V3++pIu2hH5dwfJQYYJ51MlIu5AgsHB7JTnjOtxeZrG
LAP0oTSFLexejUu9t/gXFXMGRCieuxbXJttoUhGZzMyXGk7gKnt/2OfCDwATwKnh
8W/FrbFlKbq9EotJAkx7NgpG8JofLJ0hAFDWtRl2vf5pC0XL8St47SvX3+lHPUAc
xjSlpSD8YMTL+rBFXAMwaIi6TjPxxhvzgZ5nyCHRXeo9VIfuRwcWPFq4KNrRyuPi
Xg42cHKRVvyqStakdRuhIHfXVY3fnc7NRkmkapUlpRgk8/YOwf2JPzQGaAlWxUFA
5p1Zf3JtScOCHhb8CDbW/zu6vXhpHuvtKLQ5/iD7E6cKqN66e6pWVSA09QfiaiFF
ifYCl3EdREgyGXdKKpHHm9Z1GH8vN5jS3hSEdCGYjxfoDteFH9QWRehVCQiPCgNN
USPhTfh/u3cR+8YCAaQBEOfgqusIkhbp2M0Zc6e5FSbJn18JEN+5P8vXxA1OenEv
hPvqIy1e2KXr2YJnVrvFCbTBpaKXmCDCk0lO3HLAUmMVc8B1stRdcYYD0pUDRtPU
JNbzZmEbpLcnIniVI36nuxbKrcBKH2ry8DPnkhu9MaUiB5sc/7KfN2dFWZWnzDUU
XiTc1djmgrPcqojg+pbwXEYbf7g4/qsbFJIr3XvCK/oZWgJnbI8gD+3yIARfC8Pd
1O6RkApTBtDZwAabox9lH7l3zWwrlaZpxvliP6bVDZ9X8eZXpMi7E2IA8YCkiH/R
BYlgh8/FoBoXTcVTCLGOP8CckLmEkhCnlagBrc34xRFoaamp0jBe90MMFFN6c0S8
s2ThzlTM/fMlC6IJ7neGKt9zkHYfPOxLVfPJXtabu7w8rVdYpmYq0Qavb3qydpvB
S90slnOzji0b6ej5Lv/RGInKjZ/CB3H8BUCL68ylqFmbofD588ZPZZ30uahRoP+W
BZkuugtx1tIN49zg3bjoLUB50v8UkGIp9S0/o+Chvnem9XULyi5JxYVWRSibuEa5
HTpWfAtXK/7Fk1giYUZ2EMGgCsyRFoRCJ8mLDFYuJbheCVreRjpxrFe6KBKzR+GL
Wx3sbaRo8yXfgNp+5DefyQri/JJj5X0jtkfpn75KWEhBdC72GXwvgCNuvS0k8TYq
dHNQ1OcBVy3Y68g+TzWUlwy53QSTBy1c3OXPHSlCvsglhb+AZkCkZtNOj+/FrDR7
Y8fHPc4ASYWOAMtlALvZzEOlCVmxwDGICaIbgEd9GqgtGpktnl7UuFUgYlyFJPcT
k8qUWXWG8hZx6kcgRzZqFgFta2BAuGGfkm7H982wfB22UsAiIzdwG7qWL9z77nRm
lKvDwPQecsldOP/B/OHwzpOWREGUM4NcjO4YkC/pDN8YQhWBcIdoWc3N3F/8Bkxj
FY1kA7O0nIPSm2ZgvSsWr+E7EDphyZ2NCcnfrffRNLYLWZmDYJXo51S/Vlz/r/16
vbic6bLJpRajcd/Ocr3WHh5O72E5O+7nFAgi9vmKr93CTcnJAEpODUss1yjQlj23
EQFDbLmsYMjhYIcvddMDcNcfTujQBL3n6ILLF0F1ur0tGPjTCjvAnYusb4IAFwaT
HtkeIBeIkzN7C+CJsW/eX/ygeA5MTgS6tEnD1A2HvFdynCUbeSOY9NpmlJwpeUmn
wESucHrzxPw9T3uu9a+vDCBP82t8aBg5TMHwIIxN1BzVMPxbzhVkcHdNA06KMTzp
6meET/j5hjFnoNAB9GNi8C5mOdSHJGDi4jMj6gphBWxu8f5LP3fznu5U6scckqTb
6LDJ1p2pb0Kv6ACVccCaCblGHzHoHeQMqlMH/H/C6afWM8x0G4L8W9jdvKb6mtBY
Ctex+d06fWsntkQL9+3fMbQYWGsmL4NaoOTLW9SfIzdRbEkNjg24CbKrBpUGGgS7
ZFF1HoFyqCpCzpW7d3Jl2GFuKAFmSnxvmMLakI7spJm9r78jt/0p0uJT535LeIix
9OSIhBCxasasHQ3xh1ME4pRKrzotTL3atmd5Kq1i9ifUYF0KPx7OjHgwatM60Um0
CvwDC9vrneySVz5lI1rFTF0bI0bJ2OchZRn3W7soQnDIKqtav11HDSFf4qRVwl0Z
8DgyHntW18T/P9fISpn1YvNkpO/hOH200sPDbeiaEEyBtGaQ0cVh96ScfuLN2pQD
Bzr91NT89Q25DQr+DAvic40OZYes7CMpa3oeIayEyi2HnIGTR2U8pN7C8HK7yqcT
tFCgGEW/s1hNpPoDKUgA5INALkBZL+NyJ7hHA8g5c9cD9aAZnF4KZn3eGrxI6TuU
QcnBnfLo9LHhz1Azxw6D3sognAO3xH7x6c7QmjQ0HBzdAvfaK8W4bQh6tKiGQbVx
HCAPMPQemXP3JvaMihbLQiscFZxOPdXNJh8V5rgLCH06Grg52EwHx4kYiEja98ml
ViT0ycrPPXgOtTY8f12FgJkBXHSwodDdrgFSrr+xW3YQqsVwH0Mb532V3KS20IRx
j8YPyUKmiNVnCl7hT5ggw+8j/5AKaQCRQMiyb5C7I6KTUXGiyb9u5hj2AMzek5Yc
mMqoYMiEulPkUSigZAEdFDdMhDcRp5WOwHuvcEkW53PllCv5OlB/EFlyob6EL9zJ
ZjotbeFm5aNNpJwsntYi6Nc8iWrP+1tF9lw0IyT5WX7jmhTmyvQTrHY+uoMAQFHv
3OKWisosgO5/tXlq+cJqtcmR9KBWxrIC/QUUpJ9BuMcWUqZgLNGhVU5K/sPII0cM
Al/flfUR8H8kvTkIpJUXHmxC2jOGGFxAE7Lvqa1sE/UZCxv96VxSK/8f/8jDxRhI
k2DeRz9DUJdDRBCFDSSWxGzTiUeud0+W4mrY01yNxBRrcpjDl9RtLL9BpBrl7vaR
U4SycZMbzHShbGx8vmTW4y3c3P93sVIZm/xeY0X0bcl/yW9JCrp6Je0mQaTFCtQY
B4/4KJSKLINtUfL3SIHXmJ6syF4gX1Xo46KbSSKHW+ZVFIxN/SQ2Rl4cIsi5hnkP
8tP6ah4DZX7d3JG6aqeeUjCVjyrlE6qxw1aS1OaJuIEqod52Y1wf/adUNFE17Z3X
lGfDensHWXyTpCZ7Q/5AlWTAmNkPG4+bxyLy//1+WFtD1IbQWI7BKI1LrvDBc2o9
XBnwNvfTj30ABE1UJrt3CVGQ2oEnsOw3QajOVjijd4qRmdU5yEoMpSqndwFjMDf+
3mtg7E2YlpvBJSe/QB3rL43tQ0ZNaNMvOeeMup3P7ahXSJq0gnkQAdLi9KwAhgwK
hXURQwZ7FUHj4hcrnqTUeBLJT322BlWwkciB6bZw9NQS1hnjhwyHgvySdCnTvT/6
Pu1eZPohkqza1JjcWw4LEQsYgST+v8LTsmH+AyvOl5a2+3qOLkJ4xOFruCkWsSsw
573qI8fWVLmQzhw3n3q6NGcxKMxMrL3zOz28U1rb2pIASGNqr8Sg+1tT/0SG4GLL
f0fzzrrAH9Kh9o/1wHWzMwIBT0ymCDaJ1mHQCdTrJV59Wux6y2oT1gipyNlM/02c
XQcqviGi1qFkK8lc1xb2Ib6PNLtcE6aKNSLN/a3+tcOpaw+590bqWC3srMJdl8Xy
lvtbn2r8kHB/BHs0ocZ3mT/0rIzLXwOXx3ZNGHGh398woRMuJBlGAVlvlZqZq9vi
VO84/w3IQCSXyHfXSJBJS7IiBk8vgZHEby88ETkWuoXd3uKqo3lgdCqRLjxl7y4r
0SO6AAsQu5stZMKgDP8Q1YJvoTxingmu4WWCAw8Sz9StkOsYBg5kD/FsIxY0tidr
h/qV8rURp+tWNByUl0pp5/AKCbQ5vwwciI78tb7TF5d1hxyspMPiiqiKpPzDzn1T
f2gWq72iltdWfFnCjRTVmrvitEpaKEpbhGB2mP9z6g13ll1RvH+4fXSiIF596GF5
nL41XDe45u5P+GVIuzeo2J084nSqRBiReiRl+rOUxvz+agRe/cgSgAjtVtXIoREd
I1ZFQZTCVsjd9t+S/NWnpCGPNCX4xqnmo30alENBPE9m5327EvzHAnhAcsXcu71L
whxIyNENveM9N0aZ/9svoBzXpPLcDuNCF3Uxx6n0zUunnNYnb6l3jN2QDNCGJ4iV
wkVOlQm4//J0BuXeYo+MEiMrAc2epxBDDXIQmbQrjphfJ9LbdauxDU0NIo1twGpR
ONtZjNNM5vl5MescGFjTDDlJpzqlDm9PZKHeGb5rv5wobpX73b4J7Qm8Ag+S+zd9
pgp1rb0vRvtvagvx7e4gcXPouKmrmriW7SjtdUhyxygMKCau6jbH4UiA5aGOErI3
cXwo1npiAy5EzrHe14R5aQ1JwxFrveVdhyLi+bHjSesFnRm/gz1M5YrxmKTr9o2y
DwvzjOOq2Y/uAbmfGqY/zaRpsTisODvMaVD6z2WNimgTW6swzO5/5UYERMVegT5k
c6MaoPNfip6dhMQgNwyJR/+1+cTGnMlDuJDrGQnkVNF8g59SI4AfWXF5xUzHbivP
G99M3hCw1T0M+iX6UDdfIL7B5OVKf+oqimXVsKRFmSCJpjA1vV4GZ9ZOj4c022je
vRRM1+T3xOFPfbm7ZnN1FnGknEAZ3yJ5mkvkjvWY9KzXKXBexdToKFJI2kwnkQzk
uNGuvJ7vvglZdBNK9055oQQkQzHTjMGfZiVr4VdlzqcekVCExryP1cZj51Y9/PwX
BibDBIwCeBmWA8eol8A5JL2lrCbKyhADLQq6GDxhH/cf/63LHrRPCMjModZuNXsm
2rCYMe+nsIt6Ya1nn4ftfgRQ+4d7sLkV2wA43p0KbsD7ReGq3v4US7F/aRRR7chg
8H+7TE9euE/7iAtxQzdHr4w97HUJsXoXEpT6YKSv2HTScCle3HUbh3Yh3kAouBna
HArGUAzqmbE9npacUVmS6ziGbDdLY6yqofLlNlzS7HQh20JUlidTbq01wzSEOYyQ
8Mwnq2HkznVME7MLcVVBcMx+wlkBESt+F8edjOa2LCCl6XF6B093MWQsIVAMPEEK
xHk2ArZLHxlyXAbJ7dMmFgznUH55HWYiT4i0P78OQwIul3bcaD/wBUKI03D1T7iL
AvHiq3UiuXnWqKKCIS+GsvpcvMcWrN8ApkGneys6QBaQW59bWskGhMcAE5782wve
n4Ye0NFQXRaRLoNGv7LIjl/bTrsMAs8WNhFj+68sAy1o6QdqbRIXfQj4rln3pyh1
QsxyDOqswYeX0dV0FmdVfJfD36WCLqz8+SXnIYDU8TvRmteWgo0kMZDj2CJ5H+bL
x3WN+6XE/V8W8Bz4pROidfOwjswIKPzBe1GB6jRoL5pUlTUbTKATaLY9ZqeRTq2u
eldYD43uQnzBnWegt2HDrnnB8gfWca5QSWYPEZC/ZNuTl8ZEFgSrE3aX26dr/Y54
aiIBza2JaGXSKXpwYH20KKW9KL2Zor1iLYB68p3j66QwPP85uKTo8caZRXVlsVX5
r0l/ak8NBfJJnxKeAps41HsPr6t6UBB/b/K6AaXpCKggLdjn0z04SZK/zju8RAws
0tD+lGEzb5LIzCcp7l56vMt4PBMSLct8CbIYSKopElgdBDAAYNUOKnL4RHheEbjs
0Y2ieADtaEgsuSlAE3MlEuwvvMcIFSbOZTJWijLkXeigLfIrK12/tNs6MvIt0YcS
nFbzwZJ7Ch6tsjHeXxTYb2t9k4isFGwNrJ9U1PahyIMPGUNyOcYF7H4IBJVU61+G
ydO6xrtIR9THqSxqROmRYDjVtnc7prT1A8gv+54+bKBRWySooL58aomg8283IsSI
8OzFSYvMdYhhep9X85t2F5VoNo4Oyyw251B/pvogh+blRN96m+qRejMfIpOFR/Jj
m38B4ub1agN1QLZSNqwbyEkemcoi2kZBaM6m0LwJwTZg6LnRxCXN4kK7sDnb+MEE
gOMgsOSLkrv+yqfGfKaACO767fxkmz5WEvFw1P+BS3+Mg2sdLZvX6AiwjucAlspN
bgSOICgHL5ja1drp00vDWR/KYnCQdCAYnNUjGNa4QKrXjhQx7SWsI55j9yRyB3Fa
WKzWTdpjYT58arfo7xUOuslNdgrdXFBqDHuX291BeqC8Hno/u7L3tsJ/tHFubPW9
BM2rutFAEf4gcOyzX3FDjfodJHx6lAWcttKgLj33TQZgVrZDKfIb7NLA3Din+BTp
9xLTYm6JND5FpusMRWNrOZsbk7p+DslQzDWfiD1QiTUh3VWubrKVhwKY1sjMdH50
H6AWLsa9H/OxlzhJ74NtK+Pq6eroK+n3n6AvCLBrlxAGcz0cJ2eaP9YitD18f9eg
adQandjAuimEyeUYTZTmZkYW4S5FLrAmhuqY7+7xz+F2YSssyH2qT8UjM9HbhUc3
RN/jmu1XlQgNxjL88S2mux/qtVJpWGh6F2LkdHQTgulcVCVOGzrUcE8XZ4M+X3tw
j04QKiaNurXkMBFcDHw2iXNjMzqIJ5GS1kHLf4/XcnoqFxtSSYsXztE2z29Mrhea
ptcDB02pqXqw/mqhSio35qsgL848Q3M3oK75V5Odg23/WwaHYKH+bolaYUpqlVSj
L/0ghmohzhnkLyOcgSW94Txsjt4Ou4CHLyWsi47fHed/y1Q9b2SN8YTGOB2Kx+Zp
2tg/vugyiIGn+EyYnJWeBnL+mMhgq0IzybDYN9tAB3QOdgvtuUr9p87rzbKw8Ya4
qWkO9CmJDr7B9eEr6ghESDkLyOiAxGz0D/sQC3p/om/LD5n0ZbeO93vm8ki8GfSl
J18MUxIBt7j5A6NIrTvdpQNhJReMM0EqWXFXbkYRfZjfUozK7UEHLZktTd8fCE6s
00ZheER3mKgYuO2GH9Ci0oVbNkeihhOa+vcLWxuHFAr4JxcmxAi+oZN1X7GAt8IL
NxqUYk2XXpXatfFB6fSz6TAG86CrcrYmErOz4I05R9EHwSkEPLD+4J50Jg4TSw1t
vgH7FjhTUuOX115S59fbn+u9rfos1BcRjqi4N1AMM7iN32zWQHJtWZCiVF8TNMZ/
+BHbC6RVZL3nS8UuMX4ENTjTVkxuUp27xsiFqLNzLZnyL6zwdLeFIL9xDSl/EW+f
zADHfAU/1rEIDyZH6dyozZVZK+Zy7gnoXTMQJOprh6yHFvoiY7aywpLLtb7nQDTJ
aXd9vEZ6fEyaPSrcFtJqkG00uXjlvDxkwQDFSBnZ+c5mSZsY0+c1CZmYEtUyk4It
Ss4R7LcGabQX6dEZ03rafYr0yybeamqKgw5PxopSX0mcrKrVsrX87EDOi/KysKet
XAOnlzcebvVFgADXvA9vhc/HTFgxd9xxfrjkeSRPIEU6FdtRA3m8ltWC3B4KFHlR
nMQ0UyGgUmGNL9TdwJ9OyMIjeLqFdyzO34aczjn4luYQGB81aZEvuEBJROgTe20r
PhnbeIZ+piHeh9IPNPF5PR+kvTkukV1Ds66VDU+C/pyu4WqYCjvN7iNZbh2Vpgnc
ioI+GdezRGO+RDU3+1CJuLhAMTMPYwCTZNIrq0PHhjR7dTxLcvui04vS58di8MSZ
yUk5lKrXcPrZ03CHNvJRhnXjFg7JXY9l9vOESvFgie7obUkJdTp3WHypCf/qQ9Xg
K1CwptoCzb1dNOOBTsHD03EkjtQnbCzrxxvstumpOxBywMMEXEqLAj5o8e6EQEWA
3XEokiGNzqRM+fFGr5Yta5aQ0eglxr0U6LvcFjGXQIMFBrJN4iqdFQuFs+ZWtGkz
h6nU8rIrV4+HArzaZ1XYO5B9IwkKOw9WSSj3vOkMg9HNrWDbbrAbiT0jgzGDEdea
VmymU1BBnLs54K2tX5P4zZxIHeDlmM6ahoVj06Nn/ePOh6dnwg6yjDP29PQZUBGz
nlRfEZn6cAXx2sUq/q48H0rPa71PRg0tlx0XyTe9AaPBHi9OaMyuXczEVMc8OzB6
LsBBgBCuhhTAlIDuK8Wy1AC7gS7XSBjY5uXNhnUvLa7cS6WaGH4Vo0uxXCoZrmwR
`protect END_PROTECTED
