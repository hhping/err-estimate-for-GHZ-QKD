`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQCuwVXgjAhAA4YHi3SY6OvJHxctSH0sIUSczeh+Stz414XTzgdinH4dk5SmtHsg
7R3XC0tVjWFLcizCM3rH39SucYo5p6um3sbesEhEfybxv73D6vqi8G7i0fmwwlIt
KleEhqYZfhvNqkScYPJdbkSzhjsbf+pra9fDwo2UD5pe3TYey1QQoHxB9G+z4JPC
Y/4OXoIrza9bPyX9ZY7SXg8FwK8bDVhTnxSrmDNZRnEU1cOc04n7dFwb+IAv/2LG
jGUycnjR+iA5n5zhWWkbSlp6RdJGWl4tF0fbpZHqpFu4V+OKCv2Z3mc8Aw1BcT8e
DhkkWzO+0zayqW1uUM/puo0dVglv98PdRUP5M0+V87ELdswMvx1hXv4wiyz5diJf
F5dry6pznIbe+y4+YPnHv0GHi2jVU+0aBbQLTfuCvSg68e1RmStD4xIr2gvKm5hF
OTu7aMWk+6Qgo9j7SQLBYYAOYWJaQMpuBv8+W7hWd/caxQrO3Jv/sBu5CtuNo75X
Y8xZZ6XKyKW8yEXZpDDAMfgT2e+0bP0MPtGjXg26+jbzWhzq9Nuejn33y+JNhw9h
Ju/+S2sxLWVrjtcWMB+H/8tU7Pn1IVF3oKMl75TmEqTDSaVVjpUl6rvhFFGcROXo
XMxFb455CTxpijp/f1O0yf4Jl4jJJ6P5HnqQYiMWYunWGKvS+ZlFO+vSLSQf1WMN
tIex53nxXEN8PVrAdbcI5GSR1ZbJhHUyoqpnHb2VHB1grgGmaB3L5oRutRVJjZUO
+xfdkh3xVp7cse9HDSkyyy/xe4H+RbLKHbKbCuIxovTdyedXSdreLsipmGCind8t
tEa7eIUoij8MkcgpSEH2u0qyCFX1QCIDUqbodsBT1KUv6pcXzwjJQq/0M6sZrAkU
jlnkGcCLBYRLbhTktxDdkjQ22Cgggd8ZnRzp5AK+DkZFTec3K3aUlyFe0e2cqxCh
t0y2t+zQr+q+7mgcs1PqjXVZ1GMTwot3CNd5fx/uoPPceRCeMInxKizi/v+j7iig
NhAVrXNiCEDb99rPc6rdFcux/cz4rYVgLACTh9BXioo2he3wFAhrW1rtuqh4UOZ+
fngHunhcSmNgU9wcIy0hJOv+OLqyvHErUjs6IJI162Fyvof5JrSLEgNFHwGwzz4S
cVaKMLBv7+SvqXPWHWghQgirjqYuJmjh2NxOM//laCktQw1GQqakyqOZl6axSUaG
aXBYGfw6RmFCemV5ZFPQLj0/h1sY3NCFn/exOcbtUjLjx83dBN/I2xBnWzhHs+xr
WU2lK4yp9Nph+/ClRiNiaqk1cZhvjqvO30AHRzC2jcoK63tHGeqhd+Tt6T/3k9fL
89NWp8fyGOFKzSuLRR0X38fuUdb2IjXL6l27NGwgBntcNr14fBzeHKSsQpx0DOH/
ZiW/VegK/7c7v7SU9ym8XEU2ui2nUvulBorL+NrPoePnhMQWsBEFk9vyKGidASAs
1fqhvw6e0HgkL7EdeRXWfI8qkpwmtWqE+XZqqtMoiwxhHNOCeBOUN5wt37ew3luj
KCWjiPgpzvSd++E3iIyjWor7vaF2eq1tlHo6hgUL2zEDVeDPr81VXJwDI85kdCXM
bKU1kT/3GgjttZIzmbO3L7Kh94MhO1YjOG7jjvCfpCihDG74VVou32j/h/YyFdZE
HINwHF8QxinodgZkgXiCLe6pXkdweC1Z0TpyDbNCqu5c4/avtttG3VnWUUqAnntf
MIsvRdElNnWaM5zUY9lRm1D04quGor9J1ByJiY0MBHgLbd/N/jAqg+1mC5A+LVJp
yqo/SfFEjyLFaiNlMzu4Og47ZZ0G/wBeYkP5tmj5dn9wlAFLp5bMStj1He/63zBC
223aFng9yfIHJir7wfBxUX+86+BoZKqYzw+v3Ad6NLaBM0ElKiOwUaeGqg/F5uhr
MteqQb59Eop7392eTXvmJswO4kLnDpQgRZgC8kns0qfu7V679zHR3AvATScia78v
5E5C0oxTqJDU91ztlpcCAhehoBWE5MwdvQG23hURkJGCB3Pj4EXPZCvCUdYQFmgo
6Q7wf2E+8lHC+t4jfG8YrDUIGh2i2BVlTZPwXz+6zY5BTGMTD0qj0be6m7jfTZeg
wEC9FQuFaueBziYJjqiohA28N61iQusULbK/4UBbtAA=
`protect END_PROTECTED
