`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbVC3aLjFuLq3CSvwl+QTG5YaF5YQF4b5FHR8lFOI83CyvPDnZEZKmpDVHB0dfde
FWdZW7xBWR42ZMzqaPsrznOq0c+FUmLW+wk1Esky/CC/BJxPSHWOkcNJ1bweemKo
RrWfFYo3Hc4aOuNK2hbzJDYLrzpFgAnUP+KX1AF9P9G2j9ysPmmJr/crz4AnnTKK
PCcBZW8EAbTNn7883L6Zg6zFyn0s2IrHAJMtJs5L8XQ2BERzDHML78reJE7lO/d9
MG54925KDD+bWToNs13KL1Ok9oVhBXS3NClZcQLZ0lRiQLi+vnmTX82aU7rkaJ0Z
jqe8U0Ur7IYkrAI0lvhlqZZSRUDV/0fV6VgpfiYggt0cne4C8UIJCZQKhoUPK3Sb
eAxeNEqrGvLcpMpK37Do7gHFcHTi9qgP6Jz2SgshPPyKZZA+Md3TpLzQlTTdC4zq
B2G+Pbqn4bPOD84GseDOUfGv6v02EkdOByoVh4OQcleA2vkNZfsxJkr/FtrKhYGb
Mr6/S2+Y+RAdrwBbVnBx152W9PeoV/GlPYMgmiMvafSlNRHy0ZTwVHrN+KImgRGS
c2JtQi/KyyOW1Yxd/qvMYG0qqD/kCDKqZhs+SBtHLyQJIP9LaLfLlvBP2iKZ07Hd
+lOybDZSDBBKLdBDC0itvA==
`protect END_PROTECTED
