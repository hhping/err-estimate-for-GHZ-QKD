`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYSKh9Nnmg55+IcqMs0kHYexBXtSkzOWk0G5KxZZV1f6yDI7nWOeO+fk/HgZtcMQ
2+iADGHzyyzxr77MHjYLK/v4G4hovyG2a8oHwZm9HlrMNnkxqCfSI93xNAOKoRWP
GaSNobpNJddGV/WKwEtE1l2/JiVNNexnzI20tX3Z+taYrnIIHz56rtOrAqphA11v
eLs2OSsY6Eu7Heb6PrNur9hkvsl5U4JIY2P71Ruv/fMyctOIeceZYHEsCfW2ucAn
v+kUn8lh+9PdUjEVvlWt7BEVLNNrRSP46Bt6QJvaGHIXOyjp28EdMYyHJyF1zWwl
RDp5bCT2hGQTKK74wlJUE7p1p8FF/i5Qc+wDdRwwmhRzUA6HO9F9DflXdGko80SN
nDjaGXUWVfEBHXt+ooWYtR2APSxYNr2sGWw6wVi+EeG/Keqe90x+UZEfKogcicar
ArOw1bYwbosH9fyvfdX0K9v8VGZqvUrfR3Rr01O6SVohRrcURPmUeG/zbY462n72
3gibNrDj+Bqidh3NpoKk1c8Y6KAgmq5CoyT1p99PhhAhDl5+VyvzuUOvvybq9HPV
4S3qZ3OiWJ0eiaCUwO2G50xnL2Noz13ZcyZLzhAjbD0jvOSFH4uEZ4YSdyNz3Q3t
t5EbNMgnZDTKMeFNVESEYGBGCvx8V5F+A/XbxpgrBFUW03kjmN1SWR+oNRDsWVO0
iqmd3tzTgAWEaffhVKqbJFa9YVz3GI0fvTR0taG6n4nVh26Xyz37gTqXwR/8cxWi
Pv+oOgew7VclLgko5mZO0fpdJGZByrDRZz1JK6MXZvfsBYkPR/SAuu2ix2gb9juK
WOZ8dQ4zWg6k2Y6oGUZPF3MZGGOrWCUmRa+6yumZ/VrKgwNgxLasufjSF3+T9IeW
pHqB2/yH80CMjVwc85+jgzeSdC+MaFj4Eb2d8a1cAGoFQ0BWIT7KaAlqHOyD5QMI
4hzSUEgt38Dz4E5QpKii7RYDKrhj2kM7VAX5KqO90ENWhDr0+vF1tjrSPfldZaSa
DA2+sEu+bX9sVOcexoGQ2WItzqpRraCY9gQ449kLTFNwWw1+zTl32zJoY5xcoOQB
VLCGDoYckV9+w7bR6CduwyEpic1+GRoNqAb7gSbAOd2AyZdVaHz+IpMxEaBsJ1X9
sf8bZfUWMTdaPbH3CGPs1hooRhKF3mgq6DdV7RsVP77fe5HkVaI9UBINrEVylIBL
qHR5oh3NZegBaLo19COHmfbOVgTIxeVVDprYASypYm4yfkdJSz3rcrSORsuvwac9
iDgutMS2lBdxUyPyYCIVkT2qzm8VLgvwXOk0mBO8ko/Az8DABNRE1mYHyFOE5FKe
GxpWL5peC8I+PME35mENqKyIcRNMvxgYkwYAmZbO9FW2fNIcG0zCVn5PtwAnZAqv
mfXMHLLMsnr0eVGONwaUTsxS/b7ub7IlqfIR2u6rXgwRNdl+mFf69YsQMiEW9MKc
SpekzDR8QaYE21oJjBjc63mtG9IS2+ZjFaBVDEzUA3uPikLWgOJLe99NXQNeUjQg
YUyLKCddsptL++eJJXiazuLRNFdLiY5A7DIKvPNvkaGLW1SWJAgCzFO+xTEwqF7i
ZcinJ/Y25OsZoUF4NN058ngG9AU9pZ29lvWX5zEjFj9cEfIt2Gf/jmIyBXxv9RYq
83QxQEM/WinWouhDEK00r4W6eoidXXJBGTxVCpCrhRhaTGUP4CszqWkm8N9alOcZ
+JWMbbkQkC4uUHwXEd7hlH/nwbGiCOD8DvxWI2bPf/GdQB9QjsU5qn5wZ21ptW8h
PfgSRbpkkHwcSyxUrl3PK2sNgfvN4oage24oYHZrae4ITm/f1O4jmBPOFiZIpKOx
blD8ErzTvwmjBVvPLUXykRUYoXIInRllZ9ky77A9WfMIl2eSsWiEbIy5CKRS3Uls
9IRytZ6J24oIY2fz7hWrjCnKp/3QZNKePehEOxWS0B04Rnk4VZO1g/SHtpXAlKUT
KU79no3NGA2siXOfWY9QRuj/nYDzeKqdhbaQ8xrtO9xrDxOcRsjUcz/o2sfWkEj/
u9v6TqnO/oknkc7lvUJ2vK/9CX2thRtfHUSlgSGOlirLPt8KGCSvjcgAK4oZlvye
vBDHevxpohwqpyHupnAZVg/vy5lSmtpaepX9UhQPCRTT0pP6PF8yI/U6Cn3Xzw/+
MbO1IEEmb5PeWLIef5e2PJ1u/enNr9XF/kpJqtV9SWEsQDs824BCxwqqze2jZrEI
NqW5PxF/+PfC51/TL1IgxwTK+RPlvez10lNbCrm/Vfv7M1JMRE8U6CynBHPgw6QV
uBvL9VhQ0X3JzA8In+73XdfEOjnMO6+X7Kot35ywcgcjxqa6cyJeckGkFXNLlg1t
TjFweyLtY05rfqDFEFGrCG1QLcho26oKtyogAxP8nwvV3uwlQzg4Q43/xxkWFZbo
kaI+Jn7fMQXG+gCbu9hS96+KuY8JrWj5CuEvcDe7H5Ojst37VEfRBN7URlCZSpII
KTujvMLql5GC6TZhZXP0c7uMUXi68JVnJN2WuxXFbFp3keXtguF+Ermw0TksaOH2
jWtHhJNW5a2eav1BN9twA0+PyrBO7F7l7Zcfj9YU1ehbkHMCTjqNmMd+M0jVl6wd
JCPSE7RF6R9oTDpp6R3j/sb3Qcp5j42Osxw1pGq1PBYI38YWn7LttlPmariX2rZD
CWLXT5GrpmoK3pLV8lWXmeLyEr66tJuC3ocSLW+zHfyp5+q5LS7FBYolWA7EylxF
jMjGGkErauDGnlClHjzRSDj1lL1EpkhYgBhqUBiUWumALuLXvUMzdcPDcDt8Y9PB
cXACTnrsDqVRwVHFsAtfGIB/az0NjSKlYbLX1xPe1YzW9cAF6CiDrL2KyKvZL+D5
sVjayxdWMrzYO9nDKVpQ/nTMDb4gNiO33uG30ZUl92r6AxTNBkCVpMJb1u/T6j1h
e7mJ5t3M+7PjEj9gp4Myl3H6JWHIBaRnEw+sGyHU2SfEF5tWnWSA1z2nzcArXkhy
fFZi9N4mYUldXiBdRAC+n1tN57HE0mXq1ou/wbsAmnMjYnEuQlU7dXwxfmKZSppw
ITCE1CkA6vxzgjZbc8PWRKNeIClEmXAmaYtHB4Oa8xqtVjRbyxNsVyXEqO5kyPDZ
IlGP+NqyLDuu5wsbXXXYdA0Yj6yn8rlVTCgKLsVmFqQYp9F3JmUPpv/IOXVQOyCn
MiwtOFD+sgkRriFi2y5e/ZzR5RmveicfNX19gG/URCYxE1PErUDxElsl6lVMkNzO
e1M6YZ/T8cREA/IyifjXW7+8eq42SG5pU60RusMJ6JWsyy9GYVVPSYz0ZDz2CQIJ
RZoN7tOq/JxxX5VVKw0zMSVPusM3lz1AkMd5Hmffqsk0ijncWB1HHSD3hdJTDnHl
gXgVlVUELQfzJt9oIlgaPk6054wEMLLsQHv9yTDt4vXuzqt7k12e8A/Ta8wCK4yQ
xgVBoIszIvtbfq6epDQnnwKw20JNVUSU7+X6lKtKVSlIV/nmAc+oQ7/GlZRdS0jk
SXT3CEKZRDa346TD1k+RqOScrViHslfEsKryYeO5E+QZUnYW8hHaXqCx7ONS8S6v
MRt+wSSWuZ1B/XfNfayJ6YEggk/9pnHnLo8DxeibPGzmDOl1D87F1pwqxSoV3xeD
4XgmDD8MAP3///WXt9Omnqulh4fJ+pUzCQk561yO+D6BydQxn6WRxfxUC9F8gqEI
DrqvdK4yFW05lb/yrEs6hYyl7tF+GOA4PXtEnPEdBodImllY0wsK5BLrIGD2oUBI
BdHCglwUpyTbMaqSGJ0Yv4wpvVnvLrNjecucbknV5uSs3mDH8v48frj6GFTOPAc9
q6jHBSw29U8NqkI848OWi+wSnvW8rxANRxcH0YoC3t08RCVUI6HJU6IAraV2dB0X
y7lE0Je1sVn5cvuorNYbas2UxLwKKb0/0HqvpaquWygOiZNiSrjYN2sUGrDNEvXE
JojY1JEvVfCxsR27oBvzr2IK6EnFT/DjgzmiO4BZAEOXQmuQdkMaDhZRGkdccxG3
jT71pkD1mP44ylwOPOxO486YPO4MpMNHgsoTtO7fkLuLOH2H0h3RA1PYmNGJQkPp
mD2Pa3Fi6lTzir/ccPC284rISwqriIBjTbBjRsXg5YkBZQT1lpjIXmeZOjx2z2PV
ZrsX5QkPsGtYmngZpRKFN9L982eaZ6RfExy8hhNw9uSDhT+FKuNNghFjuOW6qAJZ
QZxuUXlvQJaFXb7NoPLaxsnZxi70LP3/HEG+St0HA+epmktlTNeME0MivGKuhcpE
Hk4PexkcgMLENpYUqHSg/RW5+Recwu4P2kEVw1FUMz6DzDBQ1kNYol2j3rTTwGHS
hIgD3T6dG2N0JEeYD0azrhTTVk/svfQl+NuPlOljBeDo6M9umfTsXlEn2rSKm73c
QRC9bF5jDTD3IlZ77ZGgI3LaiiOiz+Z+UPzYiGnH1zK0QYQBDheMtCgmcwoQjx9X
cha7hZbGSkwgXwio4cnc3rZ8XrzLxXhYKzqUOLZ3F5uU7rhbnmnP+Ny54MZ1krST
NlF64amKo6wfPg55QYjVMhAaYeOw3Twc8ePIKHib3OPcWnphUGsdu1BnKGFBYhKU
e6Y/nhVg2SfI5W2+g4SmQOWQfX6H3MdKbX6LNB/liaEPgRMHhN0qEuqdj8BTVidA
FC6A0dFCEUFfrJporoud5vc2PB0UQh0ED4bDOnNdvAAeT+nRXGTvsrTg9lnfbjni
asi8jFYnfumkOTr3DOUajH1hwB6AgAaTj1BYCKTbSO36ZlS2opmnEZfwJamD2qzV
l4csaS+4IzehrKkzMv5r8HkQC1Cur+Aw/tEh+P3x8STV3ywETmuTdYJxBfZZbgmI
9MvewJtSi/IE0ZivqtrVWmpu02J+krJPVRKyZW0+GZe+bbjHx6wOfJ6pMfbATxxf
l7lmR60Qe/FyYA5neWZjp70qHhz3wM+SC4IwyZjUKD4Jt5+OLtoMQVPZAiJ6rA9/
R6wePRauLRR3L5WLOgGHr3XxBGy/ErjCzmCTZwEV/lRc06y1D19XyHUDsj/PqGgZ
g1OsHux1BqgWmjZKDaGfGwmXSj7bAfRyO4mSIasSpugwFP+6h7oo0kg8Ioc67etn
f1PZ3XGyxYNSaJD6l0yoDMBb+8cr0Y+9tgwpUF90S2FcndQer69+4PmM97AwNOzK
rj1GcHqNmvINu1ZosGswxNBLprMab81fSqmDLZwRobjauFVyKsztlRT9gn/0HN+E
nrSsg2X2pue4kE9ZfKnYOhIdRUwfIqXPTWTnRxKjbR8mcuqkOGr0OcYvvg2t3rnr
0/x6/5emMYgke18BZlZKgylzd1BAZOBbNUaHzxNiWpykiQ4+bosGhAAYFAJd/6XK
lLuT+QnNO8fXaRvYfRU66pqsCsK82E4t6sYSFr00sJ7f+1tE17oDhqkkbzvBUX50
r5fYHWUcvicqRs4TFHoCaO/yfHCqhN4bZeMDYmQ63Ug6D7xOJ6Xt3r63GHgoO5EE
67ac9CwgB74g/ORq5hahTm8dAhEdvO2lnxfoefq/2h1+WhXwP4PDcGuBQCaGMRdF
htPPg0E3L8tWDr67Sy96EtPZLzYghotbsB0XW/ze0IoK9ydjdZGW8MqcQC5AkH1o
Yfxd/L21FA3ncWYICmeF4dgbwmFXyE8KKI60zOl8YeBdlwh0NZNzf2PfLdGlejl6
dTxnK9RUbzHM6iChxaHA3EHkHGEy05i92Co0636hvqTwPNklnpRMgE259NII5i2B
89oxJ4u0hhqIX/csKQ37gml9CNc1O7pSDCBjq5SGhHoGumHJBXvZlQjZJ862Ktln
4+L41BVgnmszQxNzVEjuPmCDN9kwQRKFwutwhIQCWSvjKSbPI2aMeKWjz4T1Tf+T
I4A3103QZ9igEO3XX2QjUkqvoUm5cpbHQQdvcdbRVCHOKc7sXTi2yeCKBiwW1XaG
wm3F/FlzSHVbv4zyb7oA/D4RFKLvOmKn1QfFaEnPXdLlun7G/cB0NFk1bOoM6CDj
JWoYD2wOeUIe3ewNkr4PONBfmOVJsNKcf2GWqr9UFDl2GJ3V4iB9jVRHJ+ExeYQT
xipb7Mvac6JZFFe+rO3ixBuU3Y7X4r0WcYJKclOrZjAfP1IO9sjomBumI1jFkwrQ
hu9qyDVAjybblQtUPE7VgF0q2Jc1fd1NNMx3hb6u3GOeqkM7vkfYDp/oXlJGcqCO
8VCKzhWYXZzyujTRce2qvc7NDr5W2Z7gSAxCbt5dq0sqdClemUMWlTQ9Ax7AsIxt
PTRQUcRAL71Np0358LYiVfusp7KNkX0Epr0GvqBYdE6bLfsZsDZfTr2LJ2N/mcAw
3XHJCMwAVtlw+u0pLW7/BIsnp+6P8TQXfA0AaFWRDyA3LQqvHmXgae6Hg/wPO2pN
Fs8BVRah4PRiEfZz5CqHTqiauirTNYjzj9tWWBQtLDCK0J+neyCYGhx9Gr9HEU5n
enk0z+gpT8eDgugKCZYlL7WsfANDnOM/7X7bzA3QDebzua6luyPe7XfFh9DbeYpX
nrhzK91+Symq/pA5eohqggQXOj9r8g0JNHi9iXPtzC3ay4TJVOmVtRuST/K7+MLR
AXzIbeREc4A37BWtoSsLsa4cuVIoW2HJ7I12LybW53nmhj4LtYoLKxqJhsCGnvEz
THKdhttNitYfNm+k8iFJc6amMJFOdOYsSjy1kJh4o7OKAN/8IMVvOFWmVBCcYlSz
oBrIlsS8hMpJ283CN2g3FGXlFM4U6uvTrX5+jZzyjEsHH4JwUtrD/P/nbFVHI23a
pFoBVBshSg6IyZTGJ7OUHROtMav2jGO19o5dcxsBdco6hS00rafqokROOrMncAIR
FjAoc1pV8hgrjc8NolRBwrrncdVjQCk3uctrrQGhMF7IB5XUMwxo4UL58LBaS702
95rmI+ztD/q2NRjAA7eDv42v5OllGbF07GKTBs/5ozCpKIbtNV5PAwuQWIyqRfrI
7TNc8Bp7T5c9B2ySJxp/87JYD3aW4IeRNhYBDTnN5fu07HUwua1m1JWrUCc1CEfx
OO6fpCsjdw1i7G+0knkv1lpE5yS+e0i8M+nuJUwUEFPzKndgZ2wngxV1UWn8aAMZ
a8ZDSB6VcBMpudkNYRnVVjuhEU6m1r7c0BefbOqrimJmsWA65TeiAIc98023X4JK
dGw/om1/TMrLlkB60x117qK5JvU30fq6GohNgJBWEwHW1yLlKXpt0QmppsRydOJ0
SZU2MZOF0v94jL3oi4Fb7YxqIShoPp9UHqMXb4KdZk5a2NcMoTP5Me0HKaOPF9xG
YVtkAu7LUJCDpVbltqIdIpjUSUAfIMoYxxxdPUX7IWTKIesbRpOFRiLGwv/RE9NL
QKMYZtd9PggEa2Mzv0w7MjdSNCf/D43BslbbosfBTtlkVLzo3w1WjkAvkbGOSft6
Im3vzuDjWqYBhc2LobK9piUlmLpAW30Sui80OwrhyET0/oRQLMbf2Kgz3B1GTLyS
BTERitSJeeTxlxRkXtUzr1OnL14mhT5fYhVGvmv1vm56eFMIMvsW9D1E9RyI+QL+
AxETAIAhCmL0g0mm2IUSo0h3rtf7iZVrYrPe1sbNtuOdT2UfoMbN5A6Gl7IwsUfj
3Hts2M3dXmwaEczFi/CwVLG9p8t82dnvlywd+fABxG2qlOYRE4AuK6Fx9gfLFJYS
m0PIYI+hu57x7lYybPXieOaMLzP4Oyqn/jFv7w5QkNl59PUo8rwsWhdTXqk/y25E
NfyiL1OsJLE/JAAh9RUrrOkB4/MW/PZImhQ4vjKRtgFwNuNWx0mOO5EyhUsYbEx+
0YpIaeEt8n+WxxCEmvNSbaB03lLUL0fOKg6ns2fYCflECUdqOkBqk6fVcG5pEGNc
AlEI8RCjpfp/kUeWrfGNVuAQSMynOpr3Idvw6nTFxJkO/x3ZWRTynVNxgj/25524
bzTgZpHfVDrq1KfUChS6+PeBUPmmGX3z/7SpT/Go2qa+KaZlM8jlqZdcSp7LtHQy
GJDWj9xb0azZnxoy3f6XkoEoaBQG7pi4PPiNqkrZY1HfXSjD4LWIRWOmgsy8uT9w
mxX3OzuwFJ6Za3OdnMMDr2srL8NrcD02MBq81x6Q55TRw1mN6nXRSACpM/iHp2SX
bChKTUhTitEFQytzdgKUOM5tAtE+NiX85AVjgMFR25RD9T8UksGC/7ro1dbFTshN
Pwt5B+G+wcECgORijZhi/IfdNB0VtzqFCiOka8foLCZm2gQvqXwLeyMqiYQwrT31
NPkpWoQ+cRsvPPXXlWuTW6NKJy5XC0W0lyt5I5kBOMQwWEdh7WaljbBLT6m25i1e
9EUVLOuaTqNlVy27DSCfn+icWgZTqOJzfGjvmKaJBVhW8TfswDzoy+skfq+v3ej3
4gr95SVyxPjinmS/qdqlJ+EzatKTMqQngTkt+dNycdC7kXD+FaJ06fN4GYjac9Ps
vwU0+/zk0mP9wL6TFbqnuf7DToUNc9vmbsb8K9mZs4pHm/oE8G4+qRDdml1Vm2Hc
ix5fsdhEvToRYAomVwTvM+EyX8HKpsV8sDfS/zg9clJoVJtn16EoGSz8a9IIDoQO
z6fKa8DxlTkCqE07jloSRrpKcKRGFRjMpHsWWU5qtzbz8ISvXoAAjGPT3dvdo1GR
RiF8cEASvndEbIdcmwYPBYQe/kUyUVh5ZgEj2vg1vF8+GVPKD04JXty51/Pp6Hqs
IRGCEG5+JiLXJBmpwbpd+Owm4vj6BHSvFdzSpQ54D1s7NJdgQNEPwJJX/hG1sYIU
vsC8YyVMA8pzzpqhuHXu3yVLD5rCWl6He18xHrw2EHl9DU6j87g1gb/6FGyxuCVI
pK033/Zk5tcvN2JkrQ/R/NrgJmVGKVh+DCjtDi5F23rci/s1abOOcRus/ayvHpSp
wd9aJFL56t8GPnPhOApUSBnvWzbsKp8QJsvjZHPoV8ucN8HjgH7BAs+OlZUMjB+W
WHjCoqBj3n7Jnp/zq5BSr0OlbrLtrBurrXCED5me31RJp6oGvdWWqXdNTdY9QWyr
CA5TGFJ/qvIfrPCAwPorIOYF173krU1y2CRSJEpF43F6+pAbSTmE0FfSxE5/dHHh
/9sb+RD8rdH74d1pANpkahWhYYrs9VT1HxwzmhI1WdbEvmq27SGYRRaAxn2gTZT6
KfrGzqSuPiy3kpTIIuBP+cxd3YN+sopRlO3sbESa1oYExnK4cX6wL6BfSqE4/9mN
GWod+rBl1CjneJ5JG1cVAEHftbqr98xWT7Oa+eNSm2cKklnDGcb9I2ZvDUp+S40U
Kej40McWmLGsKdvwkvaj5z8ASYMnv5m3AC8dWW3KGZ30GszwRplibRDxue47IQus
0Ybw9511zZR5iwJWQiBaB2PMnQORh4l7V2uCQJJ7VeWxrcNVh/2wHQFyZzjyVpbk
AZkz2Ao/kwXG9IC+XH5BCRTJQbr1BTuftkUVTwCIQKhqsmUKkHVW8cgpEbNGVrRf
aaQ5KV9O5477Ci0lmov4t/eswjFWALs6Ma2J76uR4Nn4zwiCs1k/OfcBNRM7NC3R
iEtWUPmfcxcwyXCSnC3c4WQD/mPzVQeP1xBF+suHxNlQjhGXnEKUeB/pPKXkWnu1
DZzoLSYPC27OvUz/coGP0WJBzy5F9IaPpf1fubUJBFbum+wpYPMjWTETUrU2dzix
C3cSI3aqDh9NW1SyEhYCWIuefY9S6KwQW7mJOjNvG4hXzHmjnREivnEMTF08YS2o
hYR/szXIiIFTx4RXA3c+j8FIOdcFRSma+G5NRp/y3aQP2sb3ITGBBOb26d1zR7Gz
ul6EfgXoEDJ4BI/AEW/RDakgG9W4ag4lqtqzC6661nitufHQRP3+Sh1f8Ky4+3qh
/V+mXUnjKLJ1w8cdlJ5u5zbj5HqnSon0aT/tN/xm41U/Bmocd83d5+5frq77sBi/
DfK80UaMvJVz7xF2nGkZK+71eVAXE6HjwIQTuq0PR52QFFoYrT7WVqMIEuFsG4iG
JphkqTtIxiCiqkeRDXoiQ6J1aelqKABmnkZW3kQ5tDNEnNN9ei2/PqIknaPhuNlG
PoS7hUYKrdOEMw3j49QEQyXGwXIDPvISffFAHeQ2HKssCO+7hD+ZudVMQevq17SB
GDlEdO5EacJmYFbuv9gnhfWVeUfvkQJco9Ha+RACvZsDwPwa/zAVAU2cDYTQYABY
LhZMHPuZLGfSX628XS13b8Ev3x70aKiH64mlMlkWmMyW+ecL7GVXcA3u93tJmPzM
pw2loeCKRw68P/OUwxbpnEPX2X4Hy8zne/v/QuUNR9uRjmdeFVCF2YwHvzvT7P/5
zx4QqFQs7E4rHL0ssvGVhZTpQcMwHM8rEXWaPqfLRSnIjzAFxbwRIblpGziSuGG8
cww2bCq/wglOPlTI7pf4R+fXL9uYzC6xRp43aZPOEwn3ZAKXvaWYI0lsY1oXhJ/1
jy7X3amjx2b/25kM6bK6PQQI1bFQ2tHosBGikILcP6FrHfliUk96gzc7MdrCsGAr
qa1eZOSKR7dwfWv7khHx8u5FalgWX0f69phyqpLvENDCIP38BElFNnWlpIggy706
5w7M2xO7vhvIiFH00ehzlUy00AeN4nmmbNp6Y6llPysX9J163y8MJ1TPEWukPGkq
UcHLU/4TegoP6ARLX2FYNRmGMErfYoEupq+XV+KI5xG1I+1EjjsX/gThNL5LOGc3
jKnUMPWQWQmQwEnSjWz8h5JDqdIIjA1hC8swe3agxINzEgAtDK07nAUfpNBP7rej
Jcu+wP5SgaclOIw+gvTyryOm/AeE0bfjhfnmE6Fmu/QGACfdzWj1C2V/iYELkBtS
ePT/luzCQ2rXIV5xpHfAinwlaoPpPPAGPXttekYWCk3bEaO/WLowka558bKKLgj+
rgAxiirq0FIg7CS52k3eACP0/w/IJrhPvzKLchewUTNxLKW2lALiJD1xoAr7DO9M
lU2vjp1uqXL/yTu+4YPsWObj6cGZF1zVs5amGVZUUINWcM4q+ziezRE0lI+b7oAZ
0mzHnrn3Mkmn/gHpv17ertYwGh6ZmMKy+KGAjY2ZylqDPK1y+Eof2BqS9VrrCY2V
rSwYsE0kxFsDLn7ivoBypZTlq6M5s3rvWiPhUbsv2AwlpKTQVoNqCHnff1GYyIe9
IgQD9x+AWlrCQxs3ffb27Wdh8HJ9j7r9a90TjQhVkuoFTFK34m9T+T4hKeSodPrj
7JO89WWLqPandf7jrph0OMEuiDhlEKvJ1wsey74HyaGhX9l/hAnFuWdi6Rx+IujU
i+Ng0mQZ4UBIJlisSiGZ6WkYwYoXpj+UqQ9cyF8N4UaKtZGrXSZxl+hgGaDlJsBG
Os3VT5w9gmnqu35LZT3vCoGOkWdzDdFEx88okK25FpQvIBsYxcnckK4Tzuak8H+5
cBqa2ZDZWtLkJqTpYo7vvTfuirXMcLk5xDeHncL8fmKMfaJRQ8kNP2xv5rJj1ycC
7pzengkLn1tiSTGjWVOpyovJzHtpS+ZEHQ/1JdI8UbHfaceuYVMDi5pYzt+CQENx
Yfzxa26YBmeg0556hxnDi3rr2o5RgczjYC5CCWcU2vo4sFMDLTXo9q2X5y5QL21R
XeDw00tqHbExfElsSaksTM/PF3+Q/G6nGc4cFf2Eqzr3QzASuc2j92ViqAe2pK1f
2+52PPm1AUc+afFfOsL8IPoCNFTgxA0ojsETqtgK2sViEkj/zqxnGpxuQ+qXdrTU
akSheMtjuk5Vu1KkzKKFs3nvM+ANFm/puznJ5CvouadmBo8cesuvovf7Ruqdkk6x
K1HwrCkNma/rt/oeJ3OKnG4qRWXWmWLvETevKWSuuDNPlt7IFed2VokNNo/1J6DU
xvDr1lY+9P/afHY/3k9ib0EwqO8+9Kcq1dWXj9yWTFxLMvag5CtbrBZ5iWK9jGKq
anA7CAChl0tezEoj+080l0k2qvzM35QHuzNMuqP+ERuR43LfowL2BaKNm9gRfyJc
XAMOc3Idj5WAgfNPyw+m3WvKSNppp89cnkMTDcQyygeR/KRjVfK7ZqyTUvITUf2Z
XDBFQ4LUe8ibsCsUf10D/ivn/8BuyQ23Vh70MtOsuoz6wfrkLOpY3gbmiV8kW3tX
TjlQ5U1NK8C5cFMZQNl1r1JOKM4rq4uBFMMn9z7/6hLjkQh7TgHj9MPPKtAs0wy4
VIk5zL4A2uhT6aqJVneYaNxUqDWT//kDksi1PSB/omTRVTmzrgmbKt0B3o9z3vNB
ABnqX1ZIrqYTPLVXaujiOupz/aBy2N94H3bYmfVLxLX+KIUcghRUG/5rFxyqWF/W
dlIzL0BZeaytrdx7I2Gs18SYnQNJQUBAfyJkcghlrjsQuDuKDa8ULNqJ8nmCyw7C
a7acJHkeqnn39zOUr1xUTux22HuR5Yy89+zsC/Fnq51aa6vnl0QencZ6p/wiGS1a
cXM2yaKv3pP9XTBFb8WD8DqFfUC/i5rOjDfyCrCPfmHxuDdASkTmfZ6Fyw4HaZLD
48SAOTeWpIieiGR8nfmsvXBUesbpNhQsO8UWjFS81+su4/OQnsvf0Df27L4dPhIV
X62LrjatTEjAIYKX3XugygeBLcwdxEcGgdq2SwyJDlEWOlj18MpiwrpxUT1IaDyv
KybQwoSt+AolKyme7Yqp88GT/xEMdWV46E2O/zMvUZ3GVtKznNEqcjsSOhNiSws+
EUvDCnDlcldOGNqdIwSlwbaB8/3cr4reze19DwkVvzhWQ0aQeoc2IVJEF3fS3qJ6
Ompb8e7KMWCn29k/J6CopUA38GMHvrUvNgI4vEvayHsCM5trGoFUitjwdO+IwNA0
we+Jqx2RVuUAheXSLLWhMz9ig+t5Vo35WxA0etl/XCZNO2nWuo3sBCCHQ830virj
KxrdrGbHo9eJBUGBwj50Fg8QI/H9TP4EBY3ATbOiQrfnxeAFYtZtglA+Tb/0+k6n
viD4aPa7fc9uXED3BozaXS/ZoUtZVX8UWHOiPRejQP2j0Qw9Ydftc6+d2D8gW7kU
eBLpfHCb1U1mfeh/3iTO/+P4Vh9BfKu5hGWvK74/msg7FbEaFdCyFo5cqPO+C+2+
I7Kf7polP0qyeR1ySQZSsBhAIeU+SlewIiasiD5shmpMhMdJ9oPgUsKOfofrRbHL
T7sPgOb1Ar+L1RgesWaj7uWgHaTU9zCc+RVr8IGWZVdL/Wb0N1/qPmROBo9E6uKU
4r5FjmWozh6G31NpnDLDyLhbSodSc7uwAWHZrPd23ayWToIAPjTQEcQMLMGhCC1R
G/P3FwW4b3aMZIGuLbuRyI+JhH3Ry9KkhrVQX3Bjbk7uOkeaTL1vb9PzpiF7LBNf
FkVWh9Ro7ecR54gWtDQkySGp318xXWNB50jvieQjIWscSU5VSzukg/p7k3i+SH+B
dMIcdzlCu2CqRP5qf5hIiXj4v5zJxfmF0xTwh45Zxcn0bVKgyCU+C8JWjZUpBaF8
kIaH/AUqwM9G1pCgslq9KVgrWg78JgbdKMTBXuQyAvFm6lbso2lyW5q27hlz926f
ljgsV4KkTksVQExIEiSYogA62qNUDzOIeBHG4LuMGzfH/ZpkE447DJxfvjYhARe9
g3rOH3VnVjP/WgVXl9lUBXd9vmjn2Vk7eRB/pWLB8DwvVeUdNYbRyFHr3ecCdoAM
cq7RXqXblZYY+ZQPTjcuk6+DhNujwj6gfnUc3XjdgbxRR6+8mZYi3cj/+eS+sb0+
zZppNp55j6c//kMrWCHhLoJ1uR/UxWDYQNLVTqs1BLrctPxulQcvkuMyT/8p1pW4
XxFwpVTqh3Hrx3ZlhCKk0GbpVhDYz2bqPwiPbD5NLWl+thi1m/hs2i5zLQM2UnbV
t1WhkeXgp/O37tQ/3fk3eC9tk1Uzv/QqeYg7yMjwtX9HKImMk0SYihovLT18LVqj
65md0bsMnIwfK46ocXMO75Z0AhsJ29nzhIZfPTDsar3PSakNMubmUBSoWkma6dzD
GaxwKib9kHhDwSrpgQWvhAX6YVgzmVLqKpR8Us9Azv8rDPbXN9n63jtTp7BzorAR
lyCyU2RHfZduWSMIJsedDH5tg6JgOgsCjshm1Hx5vrYUFLFoaW8vX/P2fdAamY6u
qVl1irTjlsySGxbq1mMGsUqc4J2tEkjYC6UwMAqTyqItQYhopJaSJ6BpCPp5QzCu
gvYJZ84oINVYDU//MQIaOc5rlgTpZ7udtbqiM++2xSM868YwmyKBBOaXszedSgb9
G2ntNwO/u15UfEnuQCThhtPtMRiABol+TzoiuRAOkeaExvz9SpKgErqAwg/dMLXi
HWi0B60MQKJkXt6cGZ9+zNYomja0riVVxvPo00Slq27djwNzj952HTAwcRid4Yoc
n7PqkeSweh5/Vs2V8Eecpu9LUL9GyGdKskZ3GFljYGgDULgzVxSxRW6ohugFKnS6
tF6Dkcxr7pIv12u6tQZQiNbhzSFDQMwZIFIQZXmJDlfxPx9hXj5kBnpppjRlYKik
ZcMJlUgEK1nn8epGNnB6lPZCFd9ll2ZaKZ1LHacvjjLXukNZul4gW5vJaXD79uIu
rtTq8Jzi2PdwAyHna5bz6z/0XaNomPb0ymcJkmU63KlJm1RsSxsFtfxWKCEp+g/r
lzDY8UmH4/sz0dkPTvikWmfDmvnTxMV+KziKh15PfpRqlZHbB4oHSMGo+43pn9hb
cMV2UXnOxgpNATVbVCI1kWXUl65daWi8QeQ+KPFW/5Sbpy1dQgF/BaaCKktqC5fg
sWesrDuo+lX7V0DJVccgEHYLR0u9EFz+9X4n/Q/5VKXx82OnamRUlblOo6SgrT0Z
g+q/9Kzmc+83f434q+uQIaOEV3hb+jDTQi+Pvsujc1qZLNYibWdhBK5b9mYww1y7
YoStQyoURWdyRRyikubD9tGTX8ePa+yOA4N72r53x6zsSceYIfhlQlvLmTscCFQe
UdiQe8WtS+r+ySSnIPXGspB1/q77zcAL+0lB1s3mMAmKpG3CxcKKMT8wTm4jUVNk
BLbMy8z4kBjPROE/ttLg1lqUUjnipNMa0tZMldyCjyC8Acj/GhV4BsmiYVHkKX3h
RmS6VebWMuTvVl67xKvTQr15Mq1Lj64kaCh6+ePC/8vBbSL9pXlUdV2Y1nyFCyzo
xX9p1f9E7r+8RrN4uQQ9qVa1YrYW8ZRnwHLhRKhDXB5kRPqSeNOvyP1hujT4TeDY
3wuzWxen3z2TpSWN5Tz9br+HNmelMkBRCvdiMmCOZ0alBQonJpzzruFbOxiA6hWj
UZITAgmhAOo/Sdy9a4d0oHL4FliwvADhe5XB6mYw9Gi3gVpFDcbDVHb4U+JEwqur
+jCPxUETGa1ixOJe9IzhqOUR5KtfFGY/xbY7RAwnqh1R4jBbnDlq5qWXLh0ba0y/
ZSfHSVmQBqk2/hDny/sHmzFVrToZPtlFJh0hJDsoBP5CVGYRgs+/4t+61dgaP33W
gZU2dlnXpl9f1r/pIIQcDwoMSL04tq924JDtbkrYu3SqZzeND6n0YwOlk+OZepTX
1oFQ/33tuSORP+hGD3YuoHmrYAeSLLlAzL3paasEJaGB+CRI6ao90IQ7qYWBr7nV
FSmn3Aa9uHtlEhnXLP86DUJeFflZXFWxcr7JLVi+GSJHE2trfhR4KmeIqnd3rFSQ
c8VBsjHYg9dymL27QuXjpKv2K1AJbs7fSMwDXe2TZ8Kr+oerFNV3Qb3eT6r0Urx2
xYpMO1UVsHtTonOosSHjcJ/+0dkEu7P7jq+qtO6nkoNhMP6i0SgOEaeF7VAwVz5s
HTKplFwgPgodT4iKBxbULWGUWr6k5GA8GxzvDP2c071l0d4pWOFf/oTy2Aj8tTxW
SYVftWP1HPYnsBMO6LHkP/LLHLnUv4VZG4fsWUtOlJVktTXRPA2n5wJCnG9Kgk17
MnhgRDL2124n6mbYr3qVpbg2pxiNQJkE8pBby4fFy7FbQ7pFSnF2hKPi1zTZnTvJ
bpj5E8Xe91Lgjq2SHcrrkl0gcAKaKQi3axM910MZsqOWsb4K83Qdjmd2x3AWCIrn
QLEZ0pTZAQF0jM/X9RG5KgQC1DJuhDa3lGebnqeHbIOiJjgC9+yOiTVwh+VIirJv
t1U1ESQ2UmPh0kt4VaUEygcBw8g6XbQGfgJnghHxphvQF9/V8OlUJr5Xw39CW5Lu
L6pMFfigXK6nTttH9NnTPPi7EVaA2V+OOvpb32eFwDnaCaTfRksPALyIemD8iz0R
pLhvJ/LO6HfhyS+YrzH/XsvpNTNDPabCgYooJLRv0AMqnxi+4T8Q4YrxyJCqf7Xc
sLdN8vBiBWceRSZ7Of+PvGQTTO0Yx82hZimhkqVlDw1mHokRDHCwMJLw9ogbKmKS
nD1HzcXV0LKo/LmcdfzVCXQWqbq1IKlCasWRqZ8mZvD7/SyAiT9GjKX1wFI2QPWF
8gVVmyjfL77Lab7xHjFcQawy9PjdRewghDwwzd0ne7ZMzEsgCdf8zyJXkaQ7a3rs
SoGpXpPaP/aT3F8+R4GhymtQe8eOUIiXCtGiApwYKo4khviHZ8YULDpdXcEkH8L2
h7tMdV0Pr+XWhYm5wzS5n7MuGAaNXTIBvd1C7wqA4NPbjMKsjG5yi0fXmcwfDNsh
6ZXn8BVHtvC/MV5UGiNxbFIP2HcXY5sXAqfCV6O+n4PoHVVO4cLJBeJwNVNFOiYx
wY7YPXVigtJlQLEeue2kkWW0dU9R7e/asXaPGnaKPEHhdSs4vrfPzGITvJji1FcW
wjZtW3uBTvNj4eDRN0WJYfwkLPoJ1Lj3uTcmuIxVLzOj7I7xP+eZgN2OzKAHAlwY
VIuScEek0oJgMXVsfqsnOdZ+VSh4BNMTAaGwFF4uv+Kun0iHOkBHBEqyfjmudDDK
MAlqOZUFZs5Yto69/3FOfjZ+VWzqYwLLQAZhWSigjkrKRGIpNRZbe5plW0GNYxpY
tVlg/edGFd79qWh7QOVlL+pt2qX5kCGyF08kJNUdKINEHu9no4Dh9f7ZRfFE8BcA
TB3c7+CNPTYgxMWS6ZQ3SHdPeW6aTAJDDY8YnK+BUV0O+f9W4rnW3az7vp6A3ZmV
JBqdb1vczYFIqc+JXNg5E9+DsvqLxhv65Zkqyi42Btf2YUv7UEJZzGlrSLPX+qi3
07Tp3erufLyj3Oa+CWzD241U7Y3bGXhE+KHqZSVgIWbIvU0ihzZWcw0mr1rUg2jk
ichHmr9sko2p/h4Toi9bgUartpP0+pdFsc8Av9O/l1NnlYEcB/NllFXcCLhQLYL1
9ttNQmZLTiEKF0NEu7wu1uL4WfjN9wo4eHIsDa44E9RYAlQ7IFECP/EG2XXVxNT0
+uMkvx19nCKj/e6ySQV823kBsGl0hh6dpyj4tf8RhJTuHU8SlTVR6KJvSQHaJeyK
TlZAKpDXtYmCA5dx+nL7en3QwL3I56B4G4fqY8zocVjPv7kF6YCDq6FeG4t+SFDQ
FBb3UW5rOofc5MtCBlnZ6DV7G5+xdFwGcqyWJXNk2S7G4+nkMk0AEwRutl/6+gi5
/qnVVulCA7q7E4fO4IpYeGNPqBU02ITb4mrxWgd9vpcd7JMcQDJ91nWec8GdN2AG
RbgxYPt3ai/8WtUGZR74JL6hGiant9Ee9W1wyUVCxQ63hVJek02D1mfDHP+iSTmp
0DScVgUb1nO7Ni2bQBClkiN7jx3QoYgYJfYcpASyXXzn0FX/pf+7VhoV1rGEjiI0
5uQoi5sV5RrhKeQ43pQZe205CZ0cn76MBPDXNXKN7aQ6ADHWdHSlQOqOpbJxot3L
Pjmk4JXxbUenwcnBRIirmYvxSB9BW6hlkh5bYC7wbajrnoKJ7VUNF79qF9ofEXgg
fB1pxqJKCavQybWLxnDoSbfqocit1BuWqlQ0YeR/h4pvYpl8GIEIGxYwVh3/JO4e
9/uGTMWeBBH7wTeG1Ih21rbyQfSTfxyDv38c9wGhKzOhQtlrNMtZm39zBbWEJdmb
i3DoICk7/XYAxrMJvHgXmkC9eJGqX6eQAtcYYVqKiEhRl0RiiYDiatCC+jAE0zNG
Ddt9uiMX6IDBC4wFG1yH3eGrnF/LX4N2S/Y/bA0SURN6Yy4h4XmgiU/TUna2YTHO
e97u0tXf5qeXn7Rkd9nGJEz+jvC+5EYdoZ6u7B2gKh1AaYm/LWSgA1j1naP7KOlp
36xUJGdGdRlPssLBRMFNbmbTvtyrrojqPOI1vQn8fLLpIY0XZyqtQxv9uYcHIfJa
dhCyLNXhtI7y+WpH9JoFl4rJ0RjN9wBNZsEGtv0u2g5gsg+YSKDDENQlq9GOj3IT
0/HMTGsL2vkQkEMRYrLjq5pIYTsGibafGY86RrIbMF9q+uPtPC66aMp551szzuCf
GgZVBDmphmCCBw14rX/huV3OGta+9DXtvISFZARU4FfomRCgrG2wUXs4qHuwaT2r
0jn3aC/kM4HJUGNSXCJadJg2XqhVfmyWi888L8ZYum7b/5qj0P9BJI4rViJopuwC
GE7kclJNP6Vo//lIgLRx7mqkXUHd/ArFUY8jWAT6ddtPzsli3UYu6YtXGjichu5n
RYaoYKBht1rUceOm8Pfoo+tN91wrE5zIhzY1wXV4AGeyNkgT2AkbkKKkYtOWvb+m
2fdZTqdQ0V4v1rpQU50kpZc1us/mYGWkZrOYyF2YZFzVAlXX3jsaWAo6Dk8NIHXV
TPaPvfU2weKSQEL2BpXcgKDRx3kz0KYrVHnWdcQQNSGlITAc2+XFtYnUlWXd4Hac
KOGa8c/ApL4JSWu6B+tIeNEeAI/TjdLZa29AePy0OgpJTjiJ5oFbP3stjn1shMAO
LWbfUsD/5aF9BUJzcBcwlqzTKtwiIsQEDUjUB/7Emc7/mw6gp9XxgidLowPX+IAo
0che83utTnfEBPUsY8wNDJmHT283K2XUL0bTbDWGA5GHIpDKjEEcX1sD3pcHe6Js
8Fuvy5+prIp7w5PfEyKmC5uxiIJyPGz0XRVzfGbQoPB1+h4EgwUoLkkijiG4sn9G
qTLZOSu/5CdMWzQe+iXm/59eY/BdeYUD9cIqv5jp/f88rFn3StOriWJHE0cCUf5F
8Tsea2XCJb6f2Gs9vnQta4OTrCKAyyfGGRCWKQXnPXZNMtDKg92JcTTDZnFc9dZ7
5wtp0d9LNeLHsX4tAvyegRciwp6JhhxlWeKcSXT0fJMuHCgIZ9lIDw2Ex4g4grHJ
VvAyC73BV3guaUKpgvRO6R8mIAtcW+HglB11/q6VUSUsvp/IoYeTRfOQLYw6f5IX
AVw5boNnAOh+FLugRCgYiIEE6SEReWQWXFhtXH9HgCj8ww5uDbuCkTSVOjWsI8xt
BXdjZadOMNRHrbvoiPu6ojeJKhwyFFhIZ+6DtMCQSipT120/KSXpGm16nzC25AEI
UJFH+DfpGW7TMA99Xp0KOC1ZwzbcM3zTm5SyFbneIZsvR1gJGdNQULh0Ud5fsDBX
R240v/sIm9LCaYX5CFh85r8Dhark7uyDwoEOSiEZCHi6YQSzL1E1xvpXsKINXsmo
E030lu1CJf4gD5w1WL+pXaDnFXqSE/Y689UF5VLdqPxcuG5CGT9lIodJd0IsiJtb
fIf3NJ4x/6Pg+e52GpYDlZEAMK8ptVbO9eHschSe8Yp+k8bdr7y3uNLnCkYOjGzb
XE3fsfDONsaRpZ3NyVIwC7rt58ttDPiAvoqMAf9BM7goJw91ewTk+C+eS/efYjHg
eb6loOfc547gyLF1hGlVnrTBJMOLkh93GS8rLGoc3ll4IyZO8e09Py4oneNwIuor
102UK0rVDR9CxOby1bpRnMlfUEEkS/0XvkLLQC4QTQxibIZyEsbTzTLGTRFBYDEN
qKD6eyXhnSgIp9XSQ6Wt93vwLSzrih+0Op6H/PHNda2BbRlQ3z2fdZhPWs3DW8yi
3ZR16fnGIkJ9YK8lI2IBeV5wnATb6psaFNXrWjSryCbNHA+CTBodR4sEg9a44eeH
mylD0vKPUyGKO5c+ZpkgRTI/X0LlkMNUhH60stYVRFS/yt6kxPWK00FR9u71WtkQ
G2Qwdy8xQaYLDU0huajnyjdcEdjg6cnla7rMp5024hO84kVVYRCez6zsN3zqe4rP
PeH4Z139In2pgHFXoxo8ATJ9KeyDrLrtZZQW566fp+i1TNtJaSM2LxBFm2klNf4m
XXdysm8WuTd5BG8R4Du94nF0U5Nx+uBSMXe7woyit7AT10xAtelcn5aSMWIUve5Q
U/2tn6OYhZYVQjb4dE4N9aVPQzQAAllREha+lVi7UFWueaZvWdCGmyWtoNUhLxCS
85/fIuxOKn1tEN9SfQyCn06RaS+WZ0A1o9GsUz4sgkNTEEiAdnz7qxzy2UyYQ9Pl
IEzIAo9YEciZDNc9put3u/AFbGAGeKQ06gRskNm2Vn7BxqyibcZGRfXwRCHqD8+w
vjoryWQbCK6G7u8DVAnX43aVW6zJWNw7H7ZB5048CZl01SohqfTqGcY6FkcIXsIj
fT7w3/3RB/X8tszJw3WzcPVurUuh1jx4OY2iTPT+DJco7RuBCEqQHOQmiKf90X1d
0JvnbBtgaf9aLVia5sMX2xnRgEPRoZriGujU5XI50d8spavMgfhSgXQUt5k8LN15
iEsyVARjs0tWuKEq8vKdmmswwy3vhjfPsk2VEI8K/hevl6QSJt9NIcsmAXb5spwu
IYjvlmBDs0uIqRmHEo44dZpunWyWyVhl8EtcHYb1xzvCXHHG2EbA8KCW8OHbcBh4
TApgrXtwhk+19/T2+tHWfrDBUMUAehegOpHZa1ciwmVbOtN8jBZMzNZSLg3AcSo3
EFpx8C+2METbO4VnV8R9h5lKGAbAjEr0D6OZ9jEXnSGlj6p2NrXBRpgfuIYM7J1N
dtu/WDErFcX9DYzA55UuGc29AuEbwyTa4gb4uxhhQnM/s2w+2iKPKKW86Rq49sZr
q0jYMKA1Xu6QJtRyRsYQ4h2cBeZTOu4Os3jf610BuxAW4OTZFOpiux8nW96YgzCb
DROb1nwLP9mC0F8M9CNqAvfwUx9+iuDe0UoxI9y79tXH8+uYB1bl1qzt3TwnbBNk
SkCeFEu5WLeNsb/FgfY6dDsPvP/z4IteGc5PAlz1YXQYNCjXvkrAi2I4bp56hMXi
gyE8kT4uD8NhSl1+HSGR7RM7TJJz0PgI185UNc5byvoulCqwY8ZOVgzx05GQ3Brc
sAzyON2Jj6vejMMD/2GAfJ8QyvwkmlkLaY9/+y5jttAU+6ymZ5rIsW+2//keTjCI
Mv+Aofe02igqC8XuivJX89zkuQKw+uRWZJFeiAmFeaPZmUlRFecK7QzaWMA0Zfhn
5QFeyF/Dmx/gdqogJrZw0L1k/MgGv/PTybLj212QsbyPFf8yeVETrSxtwfCornCY
n6mVozUGVaWNVBvoJmeWnq5DnE5em330ApI/WZ/EkCZvEshLTLMZwdhOA20OWlf0
6G94U3XTmHAd4UlYPXevJUTt68qdsfNjRsz1RKQizgVrSPuKDQh9H+HhGcvaGAG3
e22t6NqXSCmBNlUSkRBPbrruiepU9x9oF/cdPEz2fEB9EXyowXhDSK6BDIVXet/N
Uj82dAwAnYjYR+o0wBHe5A5W/dzlGz5Qn5EL/l8ElSr7xTs+Nk4TJqjFgQj3uL/n
dl+vhdpzwO0dj5AvbX8dDhMUWIwVqwRWZcnakjjl1qPvItLAeCi1honQnDq6IUmK
b9p1Oj1XQtvSi0liUnLfM178lBfU+a7e0O0hXTtuXQPCwC0ycLqTDyPmN3FPLOmP
Sze25TXHWqRPewvd3M2izCaLQ6IrZvPsdWbhgn1XfJUA/U6xmqIJRmZTmbj72wtX
zh8SmhOZHrWoKekZTvsOcEvNiqb1S6JRNliZPacUxuOt2sLtdjfvE9hhEThFeqxp
J3GXgvGsg7gyhtzN+maWbKPPkrfMAE8voyZn5aAHDURL0HIxQYWyuPQi19iXp/Tg
RcZlrrJZhtG8l5yUHlWjzyEicywd1hP9q1ZNihBQ1gsbNxrQIuaZ0SXznM9cy2iD
qFeUbBHStJRKajFK/IBkInDHobfkye8OYHwetKavJIeW0j3LGa90alF2jv6oJIhX
HZYJ2Ha8+M0tRS2YVc+Kot4+vbq3VIqJrK8peY6EjqDLOju4IYpGA+gtZiBSZsva
/L7lr8DdfZY1sA7m8OSgmlPHv+EmoKppDgOMJ33eQC1w7bOHxi+FLAQsN1XrU2DW
uIA7KMR9kfM7V4OCElZBpol36SlzAvIpdZRk+6/XoslgbdO8qiBNwm/3NiB4fY91
gpag4wwTTX6EmYtUjJEoo56+bVwcjQ9z38Me80GR6hSGPOqMzWYeZ7Ra+IbkDxQ/
OBHjhCFRC6LS3fxqbwdVYgnb/xwkNJx1YgfnqRUT2PgJDrb3uptgfvGgm5djueeV
Zu3YPHiQVDNj+qQW3GH3PC54HIfCDO+Oo9/+l8pPV87UOG7VUy31LaBvNV6zyeUJ
JMGxXUgOiFmIQYuAtsBPxTOrpr/Pa+BpgaHlrppThA+VnLx3f6WU3UCno9YlRP8S
zp93g33cZnsqR7CjxsqJpQja2VFhe2yjRUi4Kodkq/w/YnvyvmQ1egCw/SxqHHvR
AZMqbEpb9kCPVO6IkloV7mQlZ3qfY046gSEt4iy9Abl1dfshgwFuX4Ww+yMK6z2f
0G96u0fg4O3XD0gw1nT6EXogB874BS4cGHjv1Mz20hpUuFNCRITlvDQSmN1kvU+O
ud9TdQHamMoSINDYKokBa7UB30Uk6X6p9vzSAMXunLqNahWUO9FmSTOL+M0RHW9s
2nhccAk6p7UAh52z9W1KHeuEup04wgO3hYxjc6+Q1ZGWd8oD8gP7iplk7V5BIa8x
lZ6Zz/aLqhc0vjxRaTP8ucl9uHNZPfuDbn6uhCAeZGlE4s+OX/vXb3Zm6tULGy5Q
JVirJtH86riNA9KsNiKrU/tlNOQqyzYcX0Iu0fr5Y3DuAx2g2z2FRcfDOuvCcfIN
pTwCYKKQtTdS2d31egUV13ARKqhqUVIT3LKXkPXR1WQL3VztUw0ryOKaVUMdG6CT
tEbQWyZcP6GiXKS82zyuTiXZG/wiq551eJ2cFYb/Lq+Qwyu0sZeqXyeyD1g82MET
Fqy0haJJ6JsJlYvV5HMaPfwXXJW4X4iTL7T03YhLneSFbniYAf3cZBVDatJt6iwL
ZR2Itn+S1Tf4X6PaHUGiFBIHlT6RU5ULtBxw0FUJ43vORYT7c7matO1KwAmaC+hV
FoYEcCGZdFrqIXJC5K9Eh1GETdsUdfgDhmXyCWeiuO8O/V1dt2vBpYqHrES5T/+j
ZZU2gHGjOtYCdt2kSdd7yAUNvHmlhLElcfh0X5d8nfpmml1gQ+T5jd7MRuYJHSRB
s7dHPUmGWaG3dTC5LME39WWPuJB1WgEW3tz8ZPbFnGbSpMdUzPGXw5qTMSB5Fywy
Ui9utXnf3GK8ez2Evqmplma4GTicequ5S5K90X/FJZ7K+FcctL4/pmS3EhxRN3xZ
94LDdeuHmHAd0Het3/5mAy3r/ytxdRTT5nvHxb4QlVQlnmXH6UKs1dv9UONOGgWT
eY+gWiblRdEYpddSGMzI/CGbCcCiS0/zBIEik4PLrJpxwW/U94pwC1X9WesIAko+
FH6pL7PUnoDPNpOrFOh6D/HEUyQM+YkQzazZfORQj/zHv0ndOOYT1qUivA9xLMFN
KPDp8RfX6shwmGXn4xT+g6CNx7y0BDj1jX4I68FoeBVP9h8+SyP/3aeI2PEZh7rY
tUzRo7sPqsI/FaGy85NqXpmPzwIsAM9sPvJamV5GUQa39QRHgHFUzAnB9dO+fb5B
kmwusIn0PCHaZmc2KHeG4b+psIwI1dMW27yAZSS50WCydwvsFM72nJCprthesaqh
xEi2oKh6LoUxPZCuWWA9Qa72yHlEjQRIN+PHvnmHei+W89qG+69uptOaFjIm+whi
5t93y/2DylvHAc40iImSXkYLmQeSIcodtd3rnAMf1Ntfa5bWCNGiz84bLKBLALqr
386pvXuZVLtG8YcZPFe22mcLBK8UuCsc0o6plLE05LyjV89Ulg+6H59RGZP1JOEj
+011S2OCyjcdBNAAZHXGy0fW/CCNYZ0eiCVxmaciJ/5kdMFpE+h0EXZTMqqlroo+
BJhOs0lEe3lkYOYc7sDhnr1xMoPsNLh/xp4j/LIHugx5Zc29MvGale0hLAp2/CYr
t/2JHnqT+GMCfvcyNORtHEZ5VVySZYWJGUOB8gwP/ofJUKyMFYIitM0sgmnJ4ikT
WueNnAlat0gtnIZXkqHUogyLzlqf2TlWR7HWyHAqBxa4sZj6cOv9SUavZZk2yxF/
01e7kQfJum7qi7pjItuDSalq9W5RItdTcMLyljR6m0pB5zz32kuO+oCRcRDyOarZ
p0N2H8vxAU2JeJyb3CvWZdf+3I+MfQ2CWengRfj3FUmRUghXnkhfmO6C7vS1sNAj
LxlUFx/O4VSZrI3TlLaBDxd//L8JaWkwWUZxODrJlevhkbIES5t3Q0kehbLfSyvJ
0xDa53T+wTA3ie9zGOeQNX+KoiQSjLcPRZs/jkqSvkrw5EECF+k8aFT82R1ywJdm
EhzXHbvcMfb3M3y7ATzz1j7/3NjiKufk+o3TdMGQlC6f6G5eUcNvL7UFGIswrBar
7fZy0A8IKYcpk4ORxCAe62d/29G1/wakOXKVoHBbJpnoEX3cJlNfd37aNpKKnYQf
lmh9Fi8If/kOlh1vBwKmkXSwzaI2hrHQB3VbNubsrIukibGa3zwoXjfetw7rB7pm
+IxTgTqsNc2ezBLxHSnhsiqNUf2jr6lIm1TnJvBxOJbNcEdvr0A72t8+JwlEcLNc
82u1PHFJ8QTAWQOeJb9JDLV6sikrnIPLvsQLZfbRXGeclVaZipnoKjsWdPmQa5vj
g0h9uaNbppyaGRehc9RLEx5zm0I1SQh3vJbg6DElgrZyPbhqXhTMNHgaO+6LiQ0b
ravJ7EE7DmCubNJonHuq9G4W9vcs2/kBU4L15/j/1ClS69T+zEPvA1aJeeLYJVhi
I/HoT/GJH6+R6bcEPFZEkmz2HLYCzpHr3FP8K5Wp4vmhHUevpYwAc8CumZenikkA
iSiY0aAXjsanfX/cfypckyh8dwMcta1TVMxVV+qdgpp/aE+tJvm0ldBlLIPsaY1v
kZRNcnft12GbLTrkwcGLgAbJuMvFu6ajy18eU+zVQDBlf+xL1Lmrsr9FNU/OaBJ3
9maiYV9oJohx/VG+cFK8S3qGbf7yqrEgHuQi2eY3s0IdiKPAeFzW5LOaYWSN7WQc
SZDRKo3k+rk4eAe9OedtBjqDNbdHiVYtY6RV4/Rfl28y2wt4gOZ0+M5zSp2kxO2h
TCDURwlnCtXVUexd8kUGlN/6LQaYE8FFCUBz0qQYCLvXGYCVzFGlOjHA5uQvU/r0
PYqJrHDB2WNUM9d6izn5WBgyx4pBMhcokPZZUCzT+PbhkAh7dpMCwxY67l0Gw78r
pWtmFy73XCYO3WViYNjE+Tn23PnwNenbuTyF+95VQB1eVOTn57RFf7rcNFdsrATM
lc7oyYzVdu0D/1AyIaDjt/0yVa3HBhCI74hd3R8Iz4Lv1NN+Hr604sArvcciHR7a
kkJ/A8O6obwly9SSNqDwhOGxhe8zbRr2RPiHB2iWTsdwBjqt/Cps+d3QwISJ7XTF
feoltkms3qjyGYab2540B7S966gYY6MojOuUpVWh8iGlgcWEhiQ1SnW2gSo5RwZT
HAcIovCGWiuwd+TLMr6WITfxzIm6HBRrj51/1dAy5knerZ15gwTt9R3TPTJZ9i5Q
V1D/ZXU3BWLWoDBsN/g7Eun0U83kuSNjkb4gXn+GbUE8IUUt2smMRwZLDdkUPT0i
bfRkfezbbgmtHT8tO9s50MKL6KDFIJNZjAq6tfowbQ0qDBTZRXnc7WZX+nJATwHL
5jHWOehGp01XnJ28eXF8hOPuH3CCT01FONvCZw0E6zin7NuDtqBeyxCtq65hbUu7
+cYvPGYfyJ9g6kYVdYJomToTFXOQERXeHzglAY4OsUISfCCr05Ayhjc73/85TbZZ
3WnhApdkWBR0k3wpS/IAXgH9EMU/x6+6x1hsKV2J6UZrWXxRUyQ7YplwNV654UMS
u/b5UIZn3+YFKIEp/dAT2VKsHzPIqJIZejjQPsrlO6VJaIdVg+Mdq+Si0Ep8wELW
js0/tHoqLF+01WkPgJ1XN23dJR8o/vXEiGyqvWrk3VEGnqqj+iQdE7hGJ3eEGtzw
S3E8tndyeEn8i/rirgY89ikAt2gzv9z6HK0DWpu4M8v7klJrcvOPQwc7H9tSHBdq
4rHf+s7Yo2agCC5dE+YoaGLk0rxNeix2FmezE0iXgvSLIptOYmNqpl+QyFd4BHer
xjCQPr2yq+mvG+UF9H5Zz6qglRGU87YmTWcPR+ngeoro1BALEdJDhlapq7gDIKRc
PlY14MUan9mUwyfjHjQSQsQG7pBc4u1pE8DcrzlP6MsIASCRbOLlSnPUu76sSPAl
haq0EV+BJPSQiWYzqfIeRrTFFlwECXztdYTO+6xrC+sk+sU4LnNGVnlFS9o8W5c8
f4MZt8s64RQLkLFUjBPPveZ85+tXHkBGD2stq0Bu0imPZtIyo0cCD1CpFToVwieI
ag3JUYq3V0spKS/yUdiERIGjaXL8f0OZzn0zAUf+fIxBcvl5yRxF8rC1y6Z4pnML
fLEoShkUtIrj84TYPWoNnCb7Dhf87evIVQWOtZJyPKBkvNJ0koVFT56PkSMygl+V
53u4PPvugMfMPTryMCxYoPa4I2kM4cLPFfOh9MIMTve/ZvLhffvCgHDyyHZ+9cV7
cRGt8TFG0aa92rWku60p3nNF7TSLfWeNofVUs+DXvVV4FMYcDB1jSe9sMSH/Uvar
ILeAgA9cFAnBuRUmloN7P9hFXDDiaaGtJM+MmwtaHddsM/r36J5iu8Dwm+7mR0lX
5hq54vsgnLrvEN1jU6M2e1DS0QxAPqKv11gGkiBkheN6U2SYwlebsa2jHqTr8q+0
lv25zHyiIjP5orqwjZ9CuFVXq9J80JIAcbikzryLisiZQq2LL08U0Dd7vIsC3kAz
5GJ6wcDodwtEw/pnHUHV5Jo53QvUaHBasZdKhJoHhHbG1acn/KjCpOAhyKpkboZK
EprNlyQ9LUe/P1YPfLENqq2gRBA94pmj1N7AmF5CRNo1nOppd/lccIc9bfLDIuGB
8uNnYfYcxUx4oX7vlGJXuerITFojpNi/ZbUCXpWQNI9PR/Lm01gG93cFu3hRRDle
uK93ACqKWGCNWTvJZI97F3MVgm8AAEXgkwQs5IERtIZ60D61/IJKqzXmbOlHaeVU
/3ke4B0PlGsrqJ9UCXc1uovgY5IullNnZ0H3EbCBAY185L8FFURrRk7vTgjK+saL
oqsuWKgYUBS6fGKbGJmo3SCmZBcu+cE27aZfvXzUPQwuexEGDoQ9ZzPv87li6tw9
BGW4dtOcYd+9J4S92vuchhDHAN8VK8NladSXcBuUtq+rGWro4KDiTj9QxgRvnfil
w1oKQCnTBNBOqPkFws/n6A3eY+ZMRSn9sbGgctcWB2VVMq+gteO09HzMd5SHhaE1
Vs8IVdQcWOqUEev1jQc+WpxyWVKB1Ww30qP5905/F06kXy+uUH+8r2pCI14KRlJt
evqLaqDHp5ixyya3V8JKPloHPYl4ko6KrJwE2RWqOPclizkEm8w65l5wkuWiZt62
JGdQ0IBVhSUQNbW1ZqFI+MPZxx/9SEsMGfOn2JoiBxeFrMc8K3SqhdXu6Tiw55dC
rI5EV96DgzICqCxj75AYTNip/kMYR75sk3O686xYYBYpnjyf6cHoc2s65fKSFL6r
yVKkMnFJKH4E5UsW7H/hApRJk3C4HC9uy3bMJ5X5U1ip+g1Le/ZaU0okKugTNHBq
OR7KJYGdByLLIE6MaTeTcT+wPLkBRXZ95++RXact0nbEvrl2zzsSJ72rAkldLiWu
owG6O33vylpB2nHK+3NKpafUx2ZtdQTkjMD2TaLq3Q3PZqEBtype1zerzMBDrxRW
MzxCfdUfZVPEUEN8Pnl3NWOKsBOGHBK6VltlUlzr3N3+YrqrrVymzzl5Q9B1Nwzl
L/PWNC1PjjtUEZUY3P1gXpsOQASSTLoqCfWRtU8qFw+cDfDeHnDALkGkN+drVr9W
3NbpWSyKdPc3m4rxLJFiwo3N6hGpwmNc5mQxiPMErKoChixTIvWw3g+bEDCfJYfs
R9Rckv8imDcrLzeM7+VsDbTBpPKYHUpKAKKQ5mCc7VR188G44p8pYCRIHP75de+g
dwmi7ix7ADxdpFUe0zcbDW3ZUAA0g7G1TH9OUvJzUA1BQFPqIu89uT+j1Xjvo3i5
uHsJGb4VYsux4Ot/QqiZPGAGrTCXvP6o38PM3KpMgkXtveziDpgQS2cd6oBPS10J
WEA3hIqQ+ur8Uy32xy8vOW1z0kkUBerqEJf7gERNxIlLfUOB/gRP6YGjjbmmIFZ6
bITmnV7/hhGZoVBuyWuiuyqeY7rqJWnX5Nd3/k14g4kJF6SDLlWXdYvgkFNmCH54
Vb+X7kM54Jg5KqdqG8DT+RMqHVAv7figBmHMXbi/Us2tcHu0LD3gc8IJ+YqLAnzl
bcUifW7pVXAu8xXETAJGbwCXmzfu137F3Exn+9A64cHSnUI+fJ1jD1+BwGL+A6TB
AGPiICer4EvH4wWB+EjJv6PxvTlwJCeiOwTebnYV/9alxafMPaAbmo106z19NwvG
0Lg0TroN+FNx2TiWpDuy/9s+EjywKcMFdN7y5Nxt/wEVvI8IaHjAMuMQcBnasstH
GBtk8ofgge/x35+CHx9JBKLWK9VMmd5R23f7KGZxr7sHLXV0vATNMInzNxtqC5Sn
AOOsHOrI4vn2WM/gTP/GpB50TfgL4T8NXtQUIFjyuEp2zCFDkxoqtaqcMWWuif6d
glQ4w98YArbIVzdQTAefGjXtWy1Y/D9Wobn1rhERvIb8YU9MnDbv5PZNYYV5YXeT
pdO5cR9nsvf8GDSDJjdAZ8xaW53ZctTgdXy3lqtaLkDcYmh36STB2aKItOj+fvZC
GJ3yd6EwtgxzQOTLxJSsIV4mFQCMjF/BbNo3GgARyVOroZapQyr9MRIt3r3JP64X
M3ZDspSZCP4P/zy0hYSMOkvmWHyhvKKpwYiA9WNqlUrid5vLHKDrjXROUUTGwyZH
9uNKAgoYZ4xIeoh3/3Rwfi+7Y27r5a2HzYjnuexDwVEQ4a0+QYhQGTJJXC6sICWu
Id5C2D+aecDsQPW33yCy/XL+fHNa+PCZ8o8RSjLtMx/CuFfapB1vRKu/ymQhlKMF
k80wziJr6juIPhqbxnyZLfJmWIBINp3d+L5lfM7i+DvPlx8c1OZMbtiriDjStHxQ
rqnUwfUOrjizACT61ivm+EjRO2Vju/lmbwlNg4lI6YLYS1cB/MfNhEl13JbGiolA
S/K4JuJyj1a5G1QgGL8s/DkYrCsKaVsGRY/VZUoaE1R9EQkkeAn+w8sHCryMv0wD
HZSkqrpS3xMJvkRIKr6altkQNxmfZOYzvLToPg9RCaHIUaUDE1K9oKYlYJ6vcRXv
95n6Q7ybrBR50aAuBNasp3dRx9NyC1MPC1BgdnQxU0JPdTo534QIffdjomhqm7k1
X8lziYvtg9AkD0ZCYPQGUxfcmJq0l0EuR6QQvfp/0pqtxxLpm4vWtCapWc/rBW6v
3DFIVa2Z86ydEOctKwCjOi6shUCNMCyl97CgoQu1+VJeHsJqPkQEmvxW+5MyJ5vz
tOvS3LvvMS46MDTz1spTGH8CZdo7WWybqYehXZPgjyKSD1N6zY3M01d1HEfwXIZ2
YlR1YSlJoYPIyjjvQY6AezaxJ445FiWlF5YpU4NWvJLNrMWq5N4f+Vq+n36UXxWl
HVWXMkjPxNFQQWfaDL/toDXzChLBsDzPyV/jGXP/CWn7nd7uPzSZYDcvVtgo4e3+
pRsOKA7XVZcM3C7UJvi3kzQOdn3CPjWwlmmKO2i/w55D7Fzip67Q++mFVJK+hReA
DsgpSu+oM29lvhb+d2n/2aHm59gCJY+BrlnbhRtsIrAcFPPR8WeqpqXBGVap6s5m
LiG/AXnfKTQp3aNoWA84vt6Tn8tq8Is2o5Xv60Q+IhUK8qPSuITCrQA9Da0D5ql6
moO07qaSPTXZ3mTojayFDCx3uS5zsa7tWlVtpNKdHEsvrp7CAiyE2EyZ128lSEXT
RzOjpYqRLAR47B7IYwJL4ZxYlfG+C84BUa+fTrSKBxahP7DMKq+RscLuNLlfi0ug
ZkkmsFr3wVCp7w00nVmeG9y7v45IZflkarNa23E2ogfOTUjihwyuA/Yi8q/LoatE
QLPTbgKmBs+doZdSv6hh/U77iWQmZNEiiyh5b0DiHezRazdFI2TbnTKqXFLyPemC
iGd3zRHJyMibWXeNa72ylcBB96W05lBGCN5/pwYiI6b1Kj+K2kIeokZyg8RwZVw0
F8BGPKFGOe6vVe1oQQ5rcZ0l8dgg98Gqphvzj1T7+Yi4Mr0Zz1X7PAnlU4e/65PW
oUJ2UuaopkInieNsIYkdx46aWXxYe1doLAxLRPYcmaOzEm9rXvX4pwXAwZmpvhrD
8ICPX2ARAUoM/DIk4FL5LOKfI/iurskVQIT90OijsFzJfeSYvRqvuPgnUJ59DI2c
vybTr1aBnJBe2+K3aWT/IHKjap9fF0CV6RLeW5h3Q43gMfm1Ev0Ak1NTRP+TcQDo
zt0pPvzlEOP0JERCBb55T+NyXIxvso0EcQm0NVwzKSpb45UA3GqX73iKwghXTesQ
YXL8jJZRrlg5XwP6h8CiNVSSBigAr9C28oO4m1cDDJslVv64KcemG+ek3MNPcRs/
bQ92OmuQc3vdDpn1y7oSYrEMLgNwOOT8tvYg1rWvJdNz4VT3wzJwZ8XtWiheb/l6
yQZ/UBtv5OTuZZxvdA4lQnVbt4sQPTGqZq/QYMjjsgx0uBFkV3tSA+qpBaPi9c3F
yJZQ3kcWD2bDn8N2rX7gNUfhUtBmy3dLDrzIrM7ZvQQ9ulufe5VESCHHCPQ6Z6N3
SIuJtpWrlu86jVXfglMolF0Kv15/L8r6+jLPMSO7bKgsKJLFPf0hvy3XHsDxCQEu
p45TrI4329QP+kFox0FK+6vynxdPxFgXfbXU3J5Gw8TxCvJedE1qthIbK6LAFsbw
h0I4k1D9KnYsJxEQOx3eZ3CqVes0XOzz5HAcTFOh6lI2DhV9LqkQYHnOCDTNcNWu
YV54kJY8OVB7HzQWf7bbYINV10Jnm4aH+BdQsOItWPirKZ01MI1bhixHTrqaY4iJ
OEGey3Jz60lrXRSj6X1cY24qJT6/fCcyy2KYLVaG+NlZTbqnhSBqBhSPRR/vP+Uv
/koFGNvPOglXvJ5F3/nQgnOzGkHImwxMR1ZRElCZQzH4+Kge0D2Ccba1zLM+quhS
7XNn/En1jHF89hdmMcFjb4sg7hU9OQw1iGgM+7Q7GMRE7dJ82Y15wQerxwUIGpB4
Bj2EcsX4SgX5WF3ZYPKKXrtTNBOVmIey8ypEE/4NBy/FQH2cki7+QRhzFDCjbnPd
0ngKNO7PKyKXm6/kOkb9BK6Qb4/J3GQmFWPpaIAtIIViN+lARzKOfGxbR4wqETYN
Wy+YJNzFSUSh/Ev5RdvgOqUU3ZMEkb6wDRgdrjT2AEmm3D3mwMWW7hGeA7xHqe8p
l6HngMCz5+xc8e4apGgwlFaqk2h18RZfAJygn7fKwewqgy3qh1Zvd2bxDyFQZS4V
QXUmcwnZN2Mgm8ZsakddW5ahyGtx6p/JkzFI2Lzf4jJnSQJ+Z/geKYofx1jAan5p
kanMnbz5TD8hl8V8u2D3/GeEXBxlS5rasjbAYIBTK31Zsd8Ig4eTAl3K/3jK9WqF
07YzrWIcacDqMJ6Dn00FtCoGUkyP+p9mMNSvJtKtZKVaI+7TXaANwEuUjs+jon49
ejnhmsdlt5iLmiMKWq5eknycz2Iz1BSoOCISqsj/Of7wVFEVAah1Q+fDLZicS/qn
RdBzbPFEBlFjqFL5L7rtTs7stCzGH+fiyDwhQv+b5CHdlDizihZoPXVxXxvUSL+4
ln735LlMvYt+2g3N5vCOqqWRFPWkKOigqoUdhI6V5QPUa276JqWP2rsyuIKUnFMD
uCMIntkKP+Cv1m+KxwsmHG/EbZXEvLmJXCEHv1o2RCyoLVgY+musjx/p2yoY6/vb
vSzYzTfZuT8eoc+bVEB9LvgS1lcqMwnSoK0s6EMcj29HX8eWhaSscP4m8gkcpp56
Ey31zR5shpJXs+IbHpkQTn1v7N4paZhsuwPG4iWvNCYZrvG7cza1L9Xlu3Om0+EO
JeQVDGHRuTnD4uyd5hwrivivVDDefHkQu3yFzJ8KB6tb7YHOWKPBYjAzim04nI1+
ieyEzfuH8nyQdUjlyXQg/KFjXMmZSug4S7nTGc+hAuAk2+gC1uVh2yZdZH7A8oVA
Czs1dUOLU4vcCeU1a1FYfN9xZYr98gr+Xzk3oXn3BLovwwYcZ/nwnvt52EuHMdGW
2wAHPbuFa1KR15hegBkYfSgEGRzOg7g7W81zImfvYPVwS79tsSiPaZEfgrEYYQf+
xzKqpiWW43DkQBsguE2AGdvt//xggF3yNuY4V4nPLO+noggHuU7meDIgTCWjxw+l
xS2RC+XVIs4CapEjRRSc2nlcvkZtBgf/QLaSnq6SuLSbJRKHwMd4dfFtUGqKTSQb
XgqLy4o7wLJApOyYvEs0IN7omp/Wn9264gHlrIiYdPrTI9OgA7VaAouBvg/IE91X
E+SU6XM4oj5kQ7wh72QbkEG7pGd0dvfclA0mPKP1lx4r4JA250GEFsr5c+jWO2sO
ivBy3Fl1BXB1ftYduMoDYq21nOw78ZJODolaVjLarlR3UTAuKP/njRCobACy+jJi
5IGVNGTT1LaWyyWzkzxxRXT+SNrs6K2lIh+7ZGV1I13zC9y0W5uC8oIRlaD9CDQ6
Hf8+6JoXwdWhA6fGCCQlKASKphydXo291i7SyOruqnO35j39Xx3wjsIIepkb1rhb
YifBL2IW1g+julCItH1wJ9DR/P+Zi7Z6mnIuzMi5sw7/0I3KFFuWNeyWeQtb4S7g
9talcOyFlatlJeEvmqi/ps5vrGHoSfanhMYLRZRuYDR0AO6vOpNVz4WKXlBkGWQc
O4k9CW3LWPxrJTM+TPeG5TDsEzJuM5ruFxA779NhRWuxABO1iTMghFbBbFjzoWZG
LvzbCdS5YmEQxucpwgrEwIcafhQCJ6YSoG5H3Oz5iQyuODumncni2XbyHQhHyyuj
xKfK4Eh2NcB+O4Tbwr08cZWhfCd2BD3mtfCGEYCVyiIJmNShy+lVugN+YTdBmWeL
fQ2CzbF2nr2sLHtsS9NMYjYC0LquskovCdrPUZs7fq6P/xhA68ap+MhBBgXN3EFb
rBHWZXlwGKeP03PqIOHXBQLbz84b5Opld67IP5cyMILb8LSTUiqYgC4Fus4ARBk+
XCwwV35FPCFeH533OhpwI2gU8Nl6PGH5YUta11fq//VEzD9+8uvaLUgrT4H0o4Uh
skaxdLOqkXDGfRdef+pFWM65VtPodlqvXMu6qSI42cD3msBIlHasML2CfOo6XWxX
WxVP+yG1lMDO9qTLJ++P0AsLDOwb5YJv+Xry138mPCEbeJ6r6y6xyuoZCm6yNXmH
TfGqu3LEkTRq4C4Jk6Ai2tfDeFfDd+V/rpiheK+uLDvzF8ijwOl/BESw4vHYD8/x
gqipOQhzKM9seJlF82ot7kNpGcRrVd1ROAOnMWWWfpg6WlcVeyRPDoixSBcj6sv5
iuaqaVLi0Jfnnrh2GjWn+0K95F5E0KyfBPKBucTnwy9w2MHrI1CADhtIRoaiDjnu
M3qChY/689jIqSevNwK9G+9TdIaiesXJNCUyciwO+cN3RzhFP1ZHx6hehzURYiL/
pBhfN9MQDL3k1gSkEfzEyAAEEYfE89wJRh4B3IwrCDzQyEjC4Kz2jqG08hTY/qbu
/2sKzEHsS4kmCn1TvPFkW6lgwL+K0oTgggKJ/JVw4IpzwlylpNES/9vHE+/LQ9e8
IanEnWdc3J8flWha9nYduukCtWYN2Z0Vw0AsWI2ZZ0orBEnII++7zL6gCVl37Hip
zAFnwE2irg3Fgy+x2AoIWArmP10mrTg4ijs2wX8Tazx/g3Iws4FKsttbNEKu6rRF
f5k3V28xGIVUM724ibke3sqZ6gsnk6D36QdbZxVWSNqxzCtRultg+NR8CPPsMvub
DazN0b2fYvWnRjV7K5+x0VN6dgteBmXsYPsKSuffJOIoAHQuiDyoHWPKu1i1UTSt
lKZzmUTDwHRlWmMXl3WFFpSGxVCw/Mk8jXXYwtnr1EKmDuCP9JIQh/M9H14Dr9Xp
CZlk5Vw1ZuSBmsOV9qt1+SogVHpUGYwTZRD7P4oAixpC5mttqTJ8cGdK5nJUV/z7
S8QWHovyWNGzh8qGpAzb0wuLvTzEgjgSw8haOgSCRBjkrdTSht5rbVBH+cOONqzc
6p7EtgXT6n9U+Gp74thjYlHJgc0MYXp5Z1bLl7nUB4/ziJog5NlDtd8t1guSxZox
xLUSEvMV1KCwAv5HOJfmNUt7VOhYB+2yDwSkeYxVra9gNKFWJsS5b5cSMCMPPKIZ
TTtRC3LesHKIJSiwAv6k2xr0Kv6NNlg4uxd51c2frjDxDXawHOJNdcAufg+Z4Ggi
MoHN2WLqV9GcBYvQzCmbo5u77MvxshbrfTeGCBVnHVBRVvIWCZiWfQfQR2l6huYg
1oMImIV0zHcGJotXIM8XiuQwZsxwCa427is9aY5nvX8bBjVx5EtqWUYbHgv3lM+4
xlys7DA+R1wksF0vtdZC5LokKGmL/29/6QBOef2hDsMuarzzhOW1rohbQU9WS6GF
hr/V4rzziYzqnIdfJNrrAAl7FbkcZOSfTWFz9kAXhcwWaUlXuhfjNzgVZq4+0GPJ
LFh7wu4quaV2C7LD/I7IJNxlV1MIdceyUfSFdJhs8sda+3Seoixx3+HAgcu3g8rN
uBtiCQ1QOW0a9mkejrVdRj4sHPzW1Bj/5Q+59O+znJjuwHFyw56Am7H12MNv5fQu
yUqUvEWxF/EplBPG/dRaBBzihENt30zSqgd8kmjGGF/2AYQlq8ZUDJTxsOjPOrjB
ul32Ao7GNnMtSGfp+cIQp6t8J1wkv+nspnVC6TcMfKShe85rNmdh8fte2SLpghUp
u4wfGcdVkTPQUnA1J4MkM/IzMbe7738puX+LVIOhNce3xn3pz7bZMrpYB9xKrLTK
aF2/cgSdxBi/WGSjq88oXgCJiS5aeKhJj9SxFq7krAh0sP3NBe8r/fY3s6/WjM+N
U8pLs5FpfiqZlqZm1fGG11BGv2UbTnjGDXYlMhksxwUK32yw19fn+WPPDr0ZlrHg
RKpR5dYXiDQdv3z6+EVr6lad8IVXQVLlserOItMYgUriKnLzQwP5fgjDM/fcR+sT
oPLlnBOUTVQahgiYbL9jtZCIJUyjw12y4k/8krmIJ5VDG5vk6F1RZ4YhSFZhQIX4
5Q+O2V9iVpoqw5cVLsemN+N+O07agbV3GvQD2OasX4x15/K0Ee7S/oE7nYGA09Td
k034mqGa1yd3D3xn/X8oeQLbV+LlhNJ6BeKFAHmO/f8Wzk0+j/1s9vVkNxKGrrqU
XtzB6AXN7+Mp1kiQwfRWDKCxM+k1qQKKB3VafNp6y/EH2CGoSnGVrQO0PW7kWapC
o57WiJd3fli3rwNt9y2bFJ0OLyB0SSqQNSQ0zeLGy/zkVBfaVPK5M21fn2Wc0hE+
5nC7llJZvCOmkc6tVl31MZOBfSuvNmG8LWPpHqY+/wyyH1fnUIMs1qONhwnhyh1g
Z6edE9ML94Lw1dQzFjuPmFncS7vjGo0d1QwX2eTPZZMvPlELeODbnegDUy4FZ+mT
mLZBkNtwg79PMH3SvXprGowY71utyMkk9CXl4v5gstxwr1wGMqrPqiJUKVWT9Ec6
QWF6EyrjQfVeG4U9vLsiXEhV5u/x7EUZLfGxYGjyl6al4OdPJbkGTvgBFKypxXFO
mwbYskO3ma0VeTo6HqQ2W4lj4YEjO/B02T4sPcOzZvW+vmgOU1CjbmmC+Yzlma2o
Fy0a+hp0dbgLT2CVaAwhoSN/LppvHCQO9XNbWKzz7V4OvihY8P7BKF0wtZWVOpTf
Ea5AvWKiGTb8ExvikOfZbgVYqL51tudP8YtBayR53bB1iCApPBXDipDQmAvrJTb/
8eo/B9Jv/JBiNwUf4VNVUIeMZJlzSqebdNmlxXICIp2foGDTZwTPJoY9SvuTGB/2
VJfcfdFQb4DOSG+b/Pz3Q/hh4kXPwwTaN+P3g/7OuyR8vMCsUlTy0WzPw6qCyOCe
MgLK1pSHboWnnpO524VSSdBfXS7T3ZmVOcTeIOuy5lEl/4Set8hPQcThr2WtoSKg
8J4NG+wLwe4yECdwZoANBVtrucE4XvjFkiMnZagIJiqKoGuueatn/7kSkTE3/J8t
a8SmNko20OIbPm9tBv7kD7JdmeI9aaAC3FE01VG3fu0WBuqw7r/ds0UzIQkpjB5N
XE96xRw0HlZavJsTVlh+rq39T1pqRkL7Tw0vROQz2D8ClDxxwtbMRw4cUd7y2QL1
GlwgT6yxi7B8+EVIFUChQVY7AUVU3W+iHKTz6QMWeuLYHQ7BSzVF/Y55vDVJL8u4
7DjMiy4qrn3NpuFrOn1uK7ELa3zhXVNjUrRuCxGjjt09XBrTkuftrT5gX9N2QTtB
3bOSlId9ayyMr92XTCPTzxesZS0nrmqJkrUDxXPCFzd8Lwrc7J5/wYwVuAm+oVZa
N9LlDZe7sUyz0QsKJjT7SnvgfB5eUZE1293y8iOvFghcJTrepnrW9Z5O0u/yRHwa
awWuh+Xn0Epw1WAf2Kt8+X+Z+Ud5COfk/dFV6hsGdXnSg0rv/UA+xWYYsY02T+Gu
VC4tpwXkyoIE1chMN9EXcWJnGcxenzYFIWt0DNlmt6DA+2c4Hzu//EYovPlffIx9
StbVEeIh5bJrWL+//DRau64eHVWy4ohShRdFw9e3WXzmNnIkfZbuBnbTppQExctx
8vBRiemszFtFWfoEVw2DIGPOTjB14pbH3XCj0L3R6432oN/uq7r6DN9ehlAjKu50
G9rVIbQQdEcJTeeaIKJiYTyL6mj7y2CR4sXHNFsaL/nBzJIOdL8ortlutAW+b0u+
ivWbZcO81Dd0rHsUqlno3j6mKPYA7wOAt3A7i6Q5xIiSewq3DA5VKRwIjBrcevPA
jVyTaZiWDKVGlvDAu2K4MZ/dorKc7XUY4laj1ahowNODG2/WmvSRW/9tnAjF+dQf
JC1k5VvMzmHYGWCYf5H4vRYQDqkqVpHVPJ/GFoKyhQyRd2MnABjWWUy/CpGOTL7l
nVWz+zfvNNXFVpnVbJewhumIDxhKoo0BVZCXR+mTzHN2GL7E+8dWlRX7292jrKUY
SohwFN2RCENKKmrlDgPPUPjK1vzkf+x2mfbvK5ZyT6suyg3AG7rLes5xNG2THXaO
zNUuR4IcaRqYazAn8KIx7ZoT35kjbsd6GziEaG1Mya+yqCUrEQfuwM9Y/ewtubh5
sndJZPUOeIC8LFgsfvPAszaR0C0ziUB4rRRsj2B6cl5cO8IS2mVN7kQdbOTQPwcx
23ggwiGEXJgdyYkVyWYE/08SPLUk83lcayw4+SFgIKAHMNmHENPkX1z9pJnKa+/u
I4MFEdoAMLnbYxnUw+LDTtY8NZf3BdyVc10oUTEAOqGk9jtR9hDibpi9E9mfod38
wZKi9xtZSNtcGzd9EkrLWhNCeivg/zyArdlGZC7g6/VOLzIhKszAaUWH6V+s7qp6
zUEYhNlaV3cOTPgoVFkk/xfDVappcB04lOP4yCJpufvePK4EN7iDm2WPLJWOzVTW
JNybj7eN5wsLhJYzD259M9KvxgEQ+DhGugiXqXcmURR6gYd4RMuxnsTpOr6uFMD+
jeidTlKZGmmCfjA1CZis7a/VPzeZw5RXIUkRs9LGC4bUq0GKkLc5tRVc9nzJA8II
7KB6urLKzhLCtxFQszDhsHV9zsz5EpFWCCDRz3rsH1/aozJJVzqOh29Qc8UOVnFb
OwNM9NBVHEmQPhwWF5v6UjzG1UzC40bTB8zkuHQtjm2rhU+5/KzZym6mQCVkTf7Y
tgdbW6Al7Bflpkf8qSGycw7KwnKdJLasMTxo3JzGm2LqInZF5WJyCX2jjzl+8+Fg
BKdd4FHlLnyKuJXI07j+/lkg9Mjh+f5VJLh9uU8KasDQVQ+VSd8jpataE1JkF1Nt
6ayg3LKOqGhbitx7vw0gBwcL85hj2BslrEx7TllicG+dKeEKLoGRB9OotV45Noyw
r2IoGBlj9hSgk3zYyWlVBvpgE4nhXDybAL8M85v0tIehxYuZPG6EEjAWjSoYxeRS
GCFGFaghXabYgZoVWzNtQ1AWznxDwR/Zgg0bW1Pc/q7w5Huoo19XHGwSD6oAAcqQ
T0RmwR3VtJa0dt72B6iKhR+00KJI6ZUeQfKiAJAepRoVfzu+nZ7YfIFaXAzY9pwM
daq3O3lUIJVFJ1uamD1gGShbSod6jWNZRtTALi7l2xrnhZC9F6La7VsjFmiCiNSS
lUIcf+HDLZtZxTSdT77ck6AR3qBQyw2ewEexUtaBi16sWZf3ubTLVEKaHgI5LYbB
WEM2fAhgICSFgt8t3y/UwDK86wX4yoHj4l6ccYaxORX6yADbF/g9ryo44cWW1Yww
iriqXJJiUSEENdD+Zt7NclmMb5KLfoDYMai7KfvHNpkyhAvGmvHhrhIyGzLoJu1B
kxOc44EL2hDoDCwrON7Ypr+SKFqU4h9kEQwYGc4m3RzUw/XbhOw1q6llzOcwOH+f
/LmWWgzFTZ0ZdrpFzjLNCbUhkL/ARAUl5QtczfFOSBl2TxHsMbRr0Q3iKZCOg4OP
qvND1Ms4IfasqcvO+7GR3XyRmYlvkPTQMIAGZa6SC4/xgZ697ytTCHBOl8jBy0fv
5RQnsVojb7tN2Mnpr81l107FvT7IvrA8uElheT2KMx09urf6G/YKijmJZnmZZ403
2iHfwrYzjCL6DE3JMltzTwkvs62oCK20OSM6/dyatFiMU9SA774kGYKG6MHSvjRZ
/3alUP9pvNXNQch99Za1Rgs2ASd+zdwbFFQMzFq7mINC18dZhBLxMq8x3KzTy8Tm
r22nDu4vUzk1xzOzfTx5qM58J+cKuEbzGGL80ou8O1JhIdJ6DMU4Ng1T7Z80eo8D
LINOD0zmvbi6kx0rZaWUKIcQEYGd1SkYQ2TpbHwysp6XV4g0vDVWZbzDrP907OC8
7twVeg6WDRQ6f2zhlKP14yfr/XqhJvAGclvwhH2tQO8JBq3s9tce38mAIodCWLH3
MVTlvWOAnLMpZnKl4lTb2jbg1cajQYir9khiCt+uJxVlso3IZwWn+7ZFnujzjEd3
OG/UG7ICzfDvkEcKozkapTfYgV91i2M6q51I41CNpf2dc85lWQPmuIjr0GXAT45K
YMrGv5nN2uYHmvXUoEGBn5/pegPXSZR4m7ZmYoTB5weH9TnhEZTFDMJu55lwDMOI
ga+VgsmGjPjkgKcSKPGoG7bl/QgPz9Rs9x622j+7yyhVgrDt5eGlvq8Vin5rOkMY
Pl8/5CWIMG+46f2LOqYmYUPPD/p6RTb9d6BYGh7N9FrUXR9Mnn2SkxJvWgUGJBjY
LkcGTvshscyl8wwAMfmzpuNH+c7GY4ovNT7Uv+40nK/mvkYF6tuHDO9Rho55Wo9n
u8GsLwTdjRZqjiadK2BXPnj3vfdYhfbyUSFz5Vxl/uXN8VTwg8wiSEaV1rCZgiOw
/aR0JPd48YGEbj5Fm3KaOYPGSP+ax8IpDo+CMvWPvp0qf4qVykHK7dqmQ0VU3jud
XcsdGUR6efHbfygFz33mLNe0AL8iKL0J60aa+SKzc+8vtp/PK0RqHsyL4d0Xh5Jl
GLdq6DYU0AM5cvwnYYjCrYOP11hYPlcrQ6nfSIqOJSkdBhhaFMeXHUQaq6wr3Sqv
pS5mFqWf5uEO4viKhcpqCKo6u+xDBt70Axk9xKs1CXH+4N1KqKR8u5EiShkI85rQ
9Yc3GmE8Uhn6GTE5zcnubzVmiE/PW07SB+Hcaa8UyIvi+DX7MgJ2U+7/wGHK+4Em
9tYE7xOPo0xf2BSPW2dzLjpinFKc9RzXNOCejxpC602+/GEgYrXXB8vj4y7f2JhH
+YUmvLp5cy+tPC65xkVztvg29/hx9XPjeg0ZYyyRJ0nzGQe3XjIJunbqKko7fMsp
y+QxTXZvTv+TULWpnlmLoKiHNI1mBv6FhpVPhlQDJNH7TcwLvB8vubjlWJ/sPRsP
51Qiq6cs7ItemZF6wIy7Q0gqRGVXiLfLUZMnFfXsN1pMBV6BHtoc69Ml0zM1lUZP
+Tid+2RvmK3JJncHl/3QAEvsz0nQq3+tYeVUyzIhrNkg43RVYMgfA0hZ1+tVRYfW
jKgYJhyrjR6z5i+MEHPXyr9JViS6RZ+Tneb+rvfuUwd4Z+1fE4yhtRJC+vgHC8vk
1Z69MnDVoz2iDXkB6VZV+C8V5lNPLQnJpyNmh10pEEzkV17pp74eFzhTypJW+/R3
F9MSPQlIsK9KtfCJMe1uwEVREnJI23vi0I226LSgbFBRQ7/9kofaTDgfZh0ZZjWR
bUMORqhPFztacqslXOOICbhCNSMBHZVKCfCRb4gt+tR8Fb+jeeHZWnsH3Kn93f0o
2PJZZ+KmLotQYhHd63BoBHQlhg8AVAO7b61DFOGLTAy/Py4cN2qmCD2uN9tjzwPm
5lJWcDRHVLioplwmbCewWixkHG+51n0z5vgCdOSvkSLVtrkY65g0j25+kXPqLzhF
e4LXLdjKx8/jMV19reDIHRTVC3d5uc7QsxiQt74HQuI3ghQr3rTgN458CL3D7pu2
Kv86d8jNzM66jS765nAmYmfjTmP6lfmq5zPIuCMEu4l0rJYwTqd6SAUc6MHw/X+K
2k/CXy+0Bcl940q/CKpuGuoq/wWwoMIbtalRVysRvB7kvntAQ622uDDhzwInXvIL
XVb7bd8omJ3GsHdCbFAIBcqEf42RlKmNVlt7CRzWgOMS9fm1tAvmYVNgDkJr2tJ6
bRV9H1bYiqi8L7qs6iP1+fK5mHs3EORa2CMR2Et5UJau6BGw+Ev6ObBq98cr1xcU
gkg/r83ITBvSnw8336DwdnUvfpluh2c9guxyryrgnyfdP8onDSRhhCvDX429317a
pdZAIrcNeU0Ic/EB6Xp3jcUnD7KbTc5Zd3sDiSWyd/+R4JhvCfjs/rVr+LWJzwgW
K7s9au8qjAluS5aKDRddYOazWr/bCmNCSZYJ/Ic7xLnHE6itPjr6zI796ldaguCo
Mhr/jWJ8V9i81GBI+jNx9CgnGG/wrTs0dJFlslNxGIJeOfZCdvSyjhnnaaD4ucxo
QmYPEAHiWfYoSW4E0f5jY7qw23mVLhbu5tgT/m/NUmMJXS3LBRs7sa18ypoxPebA
j534+9ONPyP6fmShoPhVmkZrnPGh21yWVxb1l2O+FC6QNsXiSH/MO7zckJOKHV4D
w+5trW6BwIxMVl5dcGR3ruIILaBI9FLjro4x6Nhx+1jL+rl1mM7Dyi8KPIm+o9mQ
aCJoX+bR9Pq3+aeeEcwbkus2VInfLMM6aWVUVy7jpPqzssaaMrbrg5zWjqpbhL9W
6s7Jw5qncO4zvvWEIfg7EqW/IemoOK2A+FO0ll1Dc/ptRpOkdmjUFOAdIhsh2im3
pY9wKuquvLd0YirFgHojRbGMty/ViqUG4LGhRDiVyVCjLxfNJ7fv2JKxzRj1mCFf
RTxFQp5zSoVOZZyzsgllIDOKT9IKWAYAfCgDkqUzLsMQM2oTRCaEj0Pm68EKmZDB
YY5YQDcKUMAs3gCkG/eRtzH9SJ9KmRcTAlzcJDfw4RPMIA088iyRtd+1nLxAOlMN
Inr3dvcVjO+OX0GadLaa065CAW8eHD3yAD7McOCtfchlYLoi3xw1H9v7Tc8akPiT
GGcNUpVyyXD8Wqv/V1ByhAwK+1MD2W57mWKM0Jz6dHfCp1U3/pRVB7M35puxE5xg
u7Bu7lPsiSLatLHWtIs4PcwdMgTGZDxqrFqXJmlzKK7l4zSPIOyAVibmHUgWn4Yu
Gbgp2be0X2Eq/XyTRmwt5KGfu6QNpUJXfBC2RaN4H+IsCyaZdlRzZTPL9gsmmbXj
jLdvJ9m5KTgzg95x918f+LIwvoIpmMCVa1g4SLpZpbH/VZU4Q3/hPti4X9icq4F/
dVn7gu3qVDFnivwE/UUY+BxjxIhWsOmfY7nYlnlQnFJmvW7hRXL0YSpOZW/+uQV0
vXTu1tZhCbjWncbJHugzCC7dbAB9gps8pdb1iN0DOcjBcbuL3X4Nomi1apQEBmge
BEuEiwiVKwUDCUTjpk8o+jKPxIymfz/INXo2A6vALZU5x1pYjJfR4nRXtDox3rrX
/DgHu7sPm77pSj9nt+MBCKuXaFMkg9Q8yNySYHJOGCOXekxLJzd9RzOi+SUMtr56
r0toQI37Uwe9yEAZlWJPuqfNd5FVg5dl1iS3baTUg1ydPF/8duwhN7ngyxKUPtS0
BKuC7/c+eFjiRjpRi094TurUpnB31Upuj2OUaI1e/hBdqLPX7vuGT1CUcmgGIJfJ
oc01aPbztM/0dbzqzmKdQaDiubF2KzrtBvjqFuU06u1AA35wBnBiTzApTSQIrSDp
69xrPIkr+GfV0EzE7tfTaY1yt3v/9EuxZirZDPLkTDrofwIWeU6FUEZJkav//yp4
lyCniH3m/0qK51b7ORiQ0nExKmECJC+/5SqyLuxnSNBiteVFbgsXKZa8a9qmEcwj
ttahn2M5EQ2Re1PLRvW0eohwbgjmKTUBnMTsdZXx7FOXP3v6OXg/wxnjCG0aC/rA
yQGdgXE/haF+OdEvh5yWA7deFp0wy2JT2U0r38pVLQsBisNSYNDWgl0bJvGmqf/z
2tQZYV2/bUj/x3/DMFcXHyb2Z912XPlCa1STWJ/h8evOdLQaty+nM0kgPHet4loQ
YdsvvDw53HZCaTJED8YqLEqMFu4ziOlts9tYI7uJ07h5sx5s1qJNVg6fpQsHQT7w
Zo61hpBau98UcGOr9rtMxKLh0wBF/iA6Bt6mXs6hcurTdp15KMZkcLIZccQ5ZmSb
9T5mLNYyFj1DVneL1hQ+udKBzUjuHXON+eqZQzdW4PO6LgxZuwe95ugHTgQS8ESz
AkQaYJJHqLd0AbrnUassxRzxKmjQlqAE67HvAk6uYl6tBoTNOaerA78qkB9Qjviq
/+4/q+GhRCFOOAggMAAtAtpjSVoZQxD4puo1xTMSs+7Qy7+rNjRna88y4G2GKYRh
lTQPtj87KpNhbPXeDB8QppKVf33N3fxUw1A47SN/hOrIFG2XPcfmfs5IkqY/fFkK
XGp8ZtG5BA782Lo1hNAwN8G+Ob1shtMKmwuLrCxNTTWFqPnn9QD/sJJF+518+glb
7cQ4vBZOuAcr0dx13XEcNs2XnVH7QbNMtOhKViKjT6zsEE1l02TpF94Fqra893hy
WllshSd9EYuizuNLupkvckqYlHhgLyLQtzpQmKtjM5EdBf/nrxaOD3PXkLIFyrp/
+qGXmXo2fj+xg467lxA4hil/pQVAQ9gTD176jD3QAu6+BRmpug96v0Ft4GHjdEkR
zTG2rn7Bqc24aU7tzagb70ftCjniM7w8gA5t+xeASZyxaFWaAWqyVyACBvqWRzT6
NmdIJXmyGq/KKZBa4jRsAIXDLtgohyeMYb9udcS5Z5YP7D0eBiIBpnafXM91LLb5
n89XHphaMKKaTE1qX+rycpzEzl+9Eq9Bmu3fcmoZtZjhpa9/egy2++UW6xjBmxrs
VVTMNhelXS58P1Jz7usaeuTZzI1dzjry0CB9pOFikEvsloPADHCCNUfIi1QsHHmr
mACyYHjHYKZDnav2by2SvQ7FD6uW2FUfu4FXsTTnQ8ffhQ1iMqnH2kX87ZTwkuMv
wnz8WaFEEH9qDsVybPg/SMpuT55SHyploKRbiCQvFR3Jq7yeiQBcrhbFA+/kDFJm
YgOAEj9QvFwwN0TSBJmmdnhVwsJaoefiRtvNY0J/bJeSn0ua3fuRzk6NK1djYaxa
sEmawr62IGj/e493Gt8+ACYsmYYfZldFD0fwpHtNFpB40DvlI9vHflcIBEt8sKpl
5H4Z0rRUQPa53l4zW+sJTbKDENYoFf4PZo2OklXYAdRDm3yqR1vr9ehyVZ2JW8Tl
vH1G8h3M14ZWe3IXzm7PKo+5G+a5huXF7R1uf9tdgegYN1+w4WxYhG+giROX9Qe7
yL3nBhi5tiletjaGWkaF0vzEb7iCqQgTVG/CEek3lhQpGzf+rYFCMslKjlbUUE+t
0aQorruAVWFALwqNj9QkpfUX5iUaUzmTEBSGTZfESuYOFsDfNB82r0y5kmFopgPu
1Z7yW7cjTo34io6tMAv3QutI47UaDtKMbZxWCLxrUqRehotrqhWBa09F11mp1QqO
xQ86Y4NjBmwfb0HmbLjxA25TwwkkvPwpfoEiZyg/BBz3WcLJPok0GQtQkBrzJjkO
QYD+MVpAilh5hMoVnwvBDShrFJfkHi7d9tpna8GK+wcOicWvbw10xLo4P9JISGN9
2AdfMkBpEdDCG+kwFnQcxAWe36kOEYCx7O2//M9yMPyBZBFRyy5MsndxR1DOPUXw
BJnR2iWDOcwipS8uPsKvHfquttADv0RsMHtk1wcmpHmQaEP8ScFWMdiHj2LNrKaa
ORSJToKazjQrF2g/iZZxN2IcaoRmvL+ACUt9DE9KVhWYWTArvF73ad3jHq8MtYE9
ARrIvNx2R765lIrVXVYUO9o4dzC3Cpdgj+yAOEPvdiV/4Lqml+K1OaZapMUQ0SpQ
y71vJTTC//SSiG3YO8MojYbpaeZApB2RLZc6nBpsFtP6lMW8oIvyaURbzpbvHyeV
jx15QaICNwqvYfgmSiDyZwH8OVFZb5JVZdnS3PnFuZxZUblx1OlUrvhNdkKVRMFK
PaSr8CSOiBb2WUt5fEQ1qZwyN/Oc4h1na9e/lfwkQhmDrAWjGHvCz+IrxF+hv8yv
ohhXQocPYx1m/Os0Cxe7EhlQPkFulGyrzg8fkLw7CIHmwaAd2tXQ2+nqrjqAntsj
91DUGdPUk9Rzt31okxmkbfVuBy39ck89vXv+bVhi70NycM5iyZhZHPrt5zLl06AP
hLM+uif5UsSbJsjJEGbfZ+iA+p/WYJ7ujub42kIM5CUXD/nPincVOqd2PfVjLB70
wQZf/IVelKprmjBzVcSxi9G0VU4I3JjDaVmeS7ioshcId2X2BpybwEdeEK2XICcz
ROeqRuEm9rQzNqAf19jXxvbXWblQGZLtySCdwSdui7SpO/+kVoY05pLpxgevHZNj
VaAgkFRLjTJHwDMg9YEVAcPpxqm1TNcWDc6183T2n6ZaRqx21XDnPctUpmfcceh2
njGH/9FuXwKX18peYC8mSVxV5xFUjdWlK8Y5sZzB30Yzp7wuzb44fbjX4WapSx5J
4jkeKd33EFSVuXkdwgDN+O8EV/OAGwvuaw6/mmw16Iaw/6nmoW/dRCfCV+QY8dK2
wywVp1ym5Fj26EusQFPTjjyi2ZgVIeMvJ5x/UNpJCf68QmREWnEVnnPTutDZ41aP
gitfO0lgLAYVVRqyv1WaXCdKzHrejZNuXoQZ276kie3ICjKLq3F79XewhAxbDtDd
kHZk8hYRiLjtzL60kqC05NYdqMyk/MHH+PazMygW/G4bXkCnyeg2RLTB1vtKfjDy
YpLTSx5sWkR546yDXd2tfSLUjOblhI6Gfax0Io7VTeuiKe+AL5xgz2fKN1tR4weE
9FwF05c/u8sdx2S8OWb/qm4rKZ6MQlTe25Ex6CQxPeGPK/4pz9jCTK0fGR08yi9m
KQn8yJI3OMcfoGT2sNZR1b1AJso7oBTUpuCgTpW5qUdGYWlD9qgS6sxmNT0T4HcT
zAljstpC7tjCp6i+OmxNep54tSmtOAngIILed2wjv8IzXNUAK6IjZugNCEzbmL7D
KrjFHedyVO+1c1JSce3P+wFlP+WaWqNHMZIUx3UfyD1nU70OqrKcAymNxGht7Br0
kCMNrR+4pr19BNhBP/FNAZecJnxirtSGq0BrjCZz2Pi/3u3/Ubqm+3oNri/7rEH+
lDaUCi8rgOWeFUqI4JqoFbL258jrCJARKLZFz1Whlak99k37dGLSb08jVBUJjThg
cbTAJ5wGknzxlMKZiikXeTBFEWjPaywgy6+ae3sCERq5PmMWsw66p9sQ0evIIlC1
FhfYbUaZ+UHYr8tJrZo3V9sXlVfCz68sL9oIMR5qwz9ZtO4iqH+uKyX4XkQxJFlP
mnRTbjaPqT/CV03X0DGkMzLGq3vQGwu2NXVMYBC8flsgt2ROo1gIKSds+POC8tLS
WHZFs4DKM/2ckpk9tYqvxbk67w0B9/CV0OR6r2vvzGSQ0J6bsbhzSAhQOYQ/h5Hl
WpC1ZH4iAwqi0cDIRzqOT+WqeHu7jKORIr+c/OmZqwMZAiMka3uYey6M8YqHat5y
yr+NNxqLhJrZoaMXaZoCyk7OXQlYOx2/vfs7JuQSbIF3Vo1kV6nIphK5h8vS/nWb
bOn1qI3ZcTXtGDmC/6FQVxcG8HFNveiFeLcY9HU3WOXdfWHWUdTBCYHgsf+D4MDH
SWC+0EMmMorqUgK7XY/0XyN+/6uue+bzr1bzSiQtL5ozJWtPdchHfVxqo01F24pn
WOgmJWVlBtEO57VFc1LZPKHlYUx6xXqDlADBPTJHQIhwXFtIXmPWAa8icJzGORJD
MLDTshwvwjrPhjivk8UB7ZBeywy6vS7DAQ7VhCG3QPpGzMT1cheNvF8v7nsjiAkW
0dc82iAOb8KjjQuIyITVVoNI5bc6jlqYy8Csq1QurXm9zJ3/m++nf+0AUtNOp6+9
LBU25+jlzbSdWz5B5bwuogmr212YyWS7/U8uq0fS5F/DdDqgndAktoIx6acBjnNH
+FzxiOvFebZ7cWZt3hwtQC6ZNsDBEIQdFuxsndzYuXuj3ljUoloH08qo0CrHZ8KK
BgaRnBjdkmFLKUbpTha+QaWnP2bM9X0MuYMKqc7JWIpFMPxHknZ6cVwE8M2U8FbF
qoxmSOxH9qsITyxyUDzsSL3cSAjbjuFqV/Z4vSpj1NhX7cDzarM+bKUSrNxG7yN2
EMDo/v+skFwnqaWzZAzzVka4gQbNWDzfk4XHQlDEkpIL8yhtyW0ZpRFaI/iNr6vt
xs61grjj2YxdUfgvrTQ99PqiIkRaZ/WG4dW3B2Zq+t0mMt/w3BJXyqeJkrJPjgRD
QDPxgeddiyX6+iJKkv4hPu4JuAEYe4ssEFkPU+REjracjPJV8oPatVoGbzA417bw
9GtCSPMDvKqQDBXRopG/a/DxUAGdBsKaBQ6gpwaRfISbMlXhnSfxyGfBTkVwc/nT
gg+zDBq+UgBe/n9/lEY7qJpXsQKRLvM0Tye5vm70XZnNEerAYIqdNjqlS85aRiAJ
yzhAn1pkw9GTcWgcCmAFq22yrj1BkT7cPJRBjXD2ll/gqcD2emRgv2SN3REjBp01
U3qg3OFYqaIhhSI8eImwgL+qMk0vPjuYBTASIbAXfw8RCm7oQiUndYr2HF+90aVb
4iLys7LpWm18oJPiHmijbfNoNFAgWdzGgseNT0/yFroRAAHDHwSUs/g4PXP/sBpp
O34hGYvN6SOJME+fnL4C60DSo488+gnamAKC704IalH+ZZJeGNr1wrOfB2t6fKrb
aOoTW5X3cTj+Y/b0oknvng7skg8/pVUiIlhB41PYNiEVtbBS3pO0mXtkyXLfzaG6
YLQiBIoxLUvemVJB7VCDLQsq0CP0gm9w2C3HCfl13mwuBoNioqz6BtIQpdLGrow8
x5KV/ZDoyByybLKFLWo2+jtcfHs94RgpVUa6ruzWV82tbRLgB/yH2BvboKcCM381
hWBlrG5aPuIEJizmRbnJSFVJPdYE4H/0SPhU+P0YwpaZW6p9nBG34nyLAAiEekhZ
/j/VyAKk+b8u6h1nU/V/xfqlDDa2V7PQoDEdpP6pZWGkSMJVTdQghB+YOZf/wNBr
387Nfi9MW54xCdoQkrN3gZuM5Q+fdOjDqmWSscD/oabc4M7icZGZZ1E2jn4u2CzP
AgXnUls4htPzOjYiy5EiTPOYL8dk+FcLtqMDoxsnGTeOgqyG+VrJ31iyRhs09B7y
DfAgzu1JBisUEXvoOag/FDm2iTTS3eifJV/UAqgXBmBQDHzrbst9pYxMCFoK1Mpp
tP+SYoi4/gS4bCqGGuEEkGGbdhgV2OniItwebmZjnfO/OsXwUVtSBrcr0SPPoVXe
2b2NivXQL1Ve3dbQ+9TWU6SWyPAQQz2Hg+/kwhdlgWwqt64zjDI9mQP4W74uUXwR
CxfBvYl4uw3ppLVU6ANoZm0vzUsuqhWTw/BnlJgpbPgBcUie7BRPoECXIeGVQ4Z1
uroCGM9QKwTrZw2PLgn9B4VLTsNLhykx2oJDmxZ3pkQfDYISk2RB++fHS8hrwA3T
DLcwojfHkO2wF77lpbCeOpnNuFhh67EIkzix6Uxg98qSRiYIty/TY5g97e2+YAbu
Ixyp0QQ0kbXmYYJ7qHrpP1v5nHZ1wtdCCAapPD3c2w5bIZVyKe2aLaG64zrhxj5s
T3WtNNMfDOy+DkWXACWIuZyukdu2HOr4t5eUT0xFvaff0vJ8FIniSaNIgxngJfH9
6sxjxs0nxbEmNwRuHZ9dH+OqF+gDZe+XWRAqkb4qeugGyN4aMRV5HBB1yA6PKoyT
lSOTIW+48D4siMPnQvTOxx1dRBTiQcydPhvbN6XqVyeashO3MbQI9rADzdnihYRE
f9c3vUlcVF2iIQkOir82yqAR7roEREMh9yrLV3Dl1Y0k95sThev5vkse+60TPQa1
bmMhV2QhaUbuY6o2HOwd6rRuy/Zeplly3OCJxV+zdoCXsVWhbs7LzhKOyZGYq50E
xg8D289pUV4k/BkzSg9v2iWq5aeCx+cvj5eUwUZGNWXZvlsO/z4Oa6tk0GNtYynY
/ZAyYcZ8oFaymVMraQorVBiGEMWA4/COy+4o2BFyomuaR+u7ufoCFJ+6Qbzd9Fws
tiC3YBudi0Qmiu2XV2WHIfKbiLoYrZ2mXh1EUksvCpmGCFZufeyDB2ZvmVUSgDRK
z1thWMSqPta7AqzHZvN65WaWPTgJo8VkxCVPEtL+g3/utJnUIbzy1WppmnGQGw7A
t3NJmbV+2QrIGdsm7nnhGPB15b2ewQl89NrlIhyy1k++GOXeP//5icZjKIFbqYqe
fsjHZq3GvPE0+F6ZzvyH3U+kIdTBDXWf9MEaoB/BqB+cq+o4ppxZAKz+hOha1vxb
2hPY8HHrOZkD7ouVQwZ6vGC/DsBwZPLvmlTnVbyjzlTbaqhkGSVzBOJ3X/d2xyS9
Z13gEsQrW3nmQZJMz/LxIWZAmhEiTaKeO68vzVrGiK6fU1+w169MhSHyl4KPJ0Qq
znJQ8GEnWgb7HLL+h0HJgGfZyHBK6jRSiPGQgzDWLtQOciIEtZ2CEA+9bxQZApfI
botKZaDc+mlpKx8T5NiajHc5otTalM1491k7h6TiZICf9Qq1FTpvkM3ST8dTggo1
6hBJLQx2ovw3s8/D7doLuodHb66QXG//1MAJPQAtphf9tgG2Nx9ALQW44g1jgv9+
Udcuz//wFPa0J4r/oPxMXXHgLGwq0039zWHJvbw39oMLrWMpIiCy66RYKIdhGt6A
6RwzOYfFAz+H4+YeB02CLe09hK42ACw54voPtCjb3/Pd/UPXwt4xpdYPJWPVsJRC
qnQYEMk0C2DfvkiD6iA8lCgG2dxWNZfEnU/nQ+5IENkD6rd2nv/WN3y6t70/zdlp
N9QRd1VhckdIZ+kb5MmFN5nVJc08DEoqPd6BzLrVeQA3unpICrMIOnR8BtxGLish
MnQtoBYt8eumEdYkkgKLf/82mExjSBdzGPIaX/TB8afCWC3VvaPzrVNPnwY7zcqC
KY6L+ARecLi+v3bf0RX0tCbkzjIqnca+cPJytRJoWEdyexZb65jhQLTi2itFk7Ll
3hB0faucV5xRrdPqfiG/oem73fGJo397T/IqgJm8qYCKIOrP++iVrH1gs8xR0VnZ
cUS//4kSWpGEdlEBcsqM6VtSL5+D8DqeiBY1C/L0lSNRXEZOA3y57Z4CwnNJhdvj
A6y+zrPuizcm3dG921iHTBVto/bYS/Z/pG0sagF0aEfIraL1gOJwl2xzLMT4HLJ7
M00rOBkjyuLYvTxxawyAx8rcpt6p5OoX54tctCjxB36QY2noSS1JEhgpNjZ8X+9U
O/mjz4rc3EeVhvkWENAzBokV8kvZ7ShYLSlPCs74jSeLzRFvx5jFRJbK9hx4RKOG
cenmh/rdoeDuQFOB4vO033XLs60LfR8iT4nj8b2r3HuIb+Ct2nLGqgEHx4FDYYK5
Ib73gEzwvU6RAK+kh2WeijBYGOttoZyG3v4Z5VUlv/Nlz+DD3vleTBHFfNSRjimy
VbLTOhB7dhge5UMPLGQ+6kTp+v3NMoXSu2OxnTczZp7nV8FZ2tKytwCUnTFVe6Fk
k2qRlXafdKJogk72HvAZvyI2sU46wNH3woW0WyZuQwUApqYCPX7xSzDlR6Cvv5h5
5tA1ZVjUyPQyY3IgGiAVMDctiITaD29FeUq/on2rpBHnyR8DgB+UVC/zJAHw8Jkb
0V2t+X77F1vcj+EO8dj/imGlWHzM+8moZ7xwmKMV/JLwluMHkGnNjjGX4XK7Ycki
PwArHH8PJugdYwbMygJJShODM64dFNmpX0C5LmIBbLpD5uSBOjYuQlsn6Cb1xr8T
pNwGnSz2zlOQbSi5fhGN6cW+f+K/99FXw1lXsnkLhcw9YfhJmrtUPtZgVzKPOwZt
H0vf0PCpyZjseFmAumO50kuqqqmK2fECouidNN75aOxiYaLbmhHfqOx9/h4jn3YZ
XTemFAMnEyHg6XBtHnCAVaymDI1ePfBL7CQzXhwUoF45CE7gb5TON1cXyEuZ+f7d
JX4uf+d2z3+KCyZBDikY6M6sEps7esWQyNHci2spOs8VA+D6GFHTPFzgu4eDv27Y
NS8fMZ4LMOQ6/5GqSoIMCeI/ZwnOmM6MW8Q8TjNXZn0GbTuN56A1+UGov0I2iGDl
qmwPv8kU2QWnun5CHT6ou/YZ6E9b6hLEtIe2KAI72prBzVSaiW2MLbKhr7ppIYjN
O2tf+qBW2a+qV/xKoTiHM9GyA0WqMTxYbz6Al3sLRk7CtpQqtyKvpniSaQUoGhLg
qUgPH0xsLwHYphqBhaMGPPtlcJmf44mAOsxO+cftkCtbVICQHfsa2E7PYFu5Ms+s
IC5/YNb5B0a7KJ8Prz38dHunN7suBUGL9bDalG/GHpUy1IqTnvDCmLCMZDf6Jw4e
KkOKLyUapT+RV3O2ZvMXrql1xWQkKT6OsBE8E8BSrLGOm1NabtO2yIcjzLaZMD5U
GsthLxhYZC8NUFQTXPHh+ur2UESrxQ/yN7JoGB5SN9aQbdH15uGmypi+jKrvU4EA
RRAR/M9ONIE2u60ml8oE+yWxR2Cj+2RHHFb7bG6GeIJjYaKQM6vt2znRdOm+x2yN
GSHIWnhEAeXNrRfDKg3/tM1EbzTj4IoOr1gZ3hGQ7wWvMfPoJSiXS215ubhLlVo9
VFJMZjnAG6EiFkMvFvqJS8FRHbufsMiaz2+ts/n4KvMM9BvLGwMhYi+ENtTalcR7
K+Bp3Tr377zR9aw0srcSAsutvuGBy6LqOYuG4qMRJwZvlQpZaCMgX4Le+rDV0qp0
VNabB5M6+hT2kReWJ80K/ep+RRZU2h4eQC7zEX147uhGDz0YF13frkk1ZS89oEgC
ckzQXKHAz/e4uUaGDPOMLkg9BH25t7oSjHFX4kOO4DPjptuZKyZ1/6Mrc1SA2NgW
vcCo9Rfr5Mo3r8E5MHJLO8rjZe1MbtCps0gyO2nW17oOaRzgjSVX4kOr7CT+hlTt
rTtnPbNGlc20No+elg+wi2dxflvu/1a6iQJTQKObROeYW2FiBxrKXuNK6WiAfktJ
5GJqY3wMKKM4V7iUKsEDIyKEpk7t9PSkb23lOXnkF4MnBfU/EOMFZXmklytSZSO3
3w/wX4+F/Tlq4mNbq43ZDC2zqoQVxYSmA5UvwB84SbFGWiyrXG9JXU0Ygfu1QAp7
b+kxG4nC9Qq3KETFiqER6xE+yqSCirMCW56J6dyD2ye9TGs9TMGRiEgrBqlXYwOx
NaWLRFRm+6ktCjd0Ot4l3PfZCh+kQiYdKDWk2apJWbaqnRsIzWi9j/Y7rzIquaQE
hYiou8yx2xLscPS2HfNxYpNx/E+O8D0+XtRsrZCf6NS92u69ZdLnGAcv+rSCzbb7
IsgU3AI/BOw+BSsYzCHfsY6HjFA11R1raDQEh7IEjy06hSADiOVLl1A9ugscnXZ0
zPfXXIfkZ9D81s4SqfrI01v31aUAPMjxUrl4lGWpAEiIvZ1RmQ7ebXVcWi9QbNGa
CfApnT3VwFR/EhK5Ks7wXPfR75EERCZgPgfTdYTjZLpn5kGoHJ89+W8/bjkDLdyZ
z/QQKJ4w/oFbrPoh6SRUZRSMogKamjWyhYvJpveGO4iLE+2Aa1Uxfvb5n3wpcFMW
fBMaiiZQx2+ac0XAvGg1vCKVFDHv9djlxorij98sEWJZjCbRvu80fOnqhWUsbuLj
NCOG1kbv7gUejgO642LttKOyJ/KsmATHscBe02iWg74KbVlaOE+lhtnjD6rlCO5N
6Mt4U8il1M4GRSdH2Zv+WOPe/gNgWyr3QhI+icU5axNxMfgRyj1cXXuqNamluzcU
ODCCwwv4WRjYyTRo7ky8bihnuQF9DcnloxPUW71Urja55EB2VgY4Im/AcKhPVWaP
r0swjwUMjjpHUnBbKKLOtg3pCr1rgOoh3PH1/cbLCY/w05aB//lvPi0dofU/4yGM
lGd69Er7YrBsJtxqin8uCZ1eVPB6pwU1jdNBhh0wu52/gtOsH1ReQukBQnVKFiLJ
JOV9tWKZTQs3F+RzTj030yXFmU1T15AD5xiv0o8KUZ0zPE9FBHg0o0O/Ni6GSgai
fZNFNllwX/LO7EJvYkJ1Eju9LInsKeeFr3XEcrAD7ynCt5qzU0Wnr/FhQyHuI9Kn
GbuNoEq7PO/xsbgCFMEW4dPxcPzgQk/zzvqnIHam4omaqZR3cd/UUqL6f38qEba9
8iHi0sj3yrvEzyX6NEyQdr4w9sh8s8mtKyGfR4c+a0ZVETKdPU1R9FsJkFJu9nE8
XABZ/QCrZa1+kYo8xHt2q9Z28wRABwpXpayLUsAeKe4EJjutUS7GnQE1i89znaZu
DsB22O+FwDU/R1o4fHP6dg/wS+DymcEhQEwgxD1f9mHNn5bbuz6F7/2ly0FMVqQp
RCSkLI4AT6d1kol7S+hjldoB+HNZBG4N9HjZ7jjGBCLU2jNMMCkT+lWDO4HtROgT
U0bmcL4ruf9OoMf5zbECdXR+J5cF87xmYG3GtC1Nb/DdecLfR+jYnkRMtQczr5tk
YLotLu7tZYH00A/48bAmhY4RMHN9RjXzmm5sPvVlKP2chYsDkeAL1omru9pNEpP+
h8YMQhN9pCfuEiId8FEyZqu81POlxS++kn6HNKMpkcuj6txn6t9t2KNWysgUUmL1
RfcGsir9w0GKgcJFYeYihAXABHAZagHC37e9cvkl+rcTpN0Rr0vETzWkby27TPFJ
N1q1LdS9IwbKQjXGhqSGM+wcHHZBS856fnoIoahYGTFxPxIxBzkkrh6dUDiyJFr6
lFJ/lBRFU4I/xzynFgmpkDHy0j4JH9WComSEZQTVaAhM7u1etH5jdxlQXeQQLj2Q
xSF97NIt8bAgoGpMBgktarV3zg8yIKzxYN7VBNMKPGGgP38PFV9Oyvs4dxbKs499
V+NeTT6tRfKJveM4QcuhCftkxMcPf8o3PdzdkHRHPAU6bTKsJk2ZTQ1ku4g0N3lP
bCnvKIK9LNNi3fUfEWv3NFnYjIiO3wmyNma3+zP5tjcgTij0kpl2zW4YQPxwUXxH
VYEfsheymQDNAxROfzEeINp3FOmyKjVgpEX1NfC/fu6EnqVU8w4sQMOQL9H0kh/v
a0u974muFcmze8i3HGzUERWNFadKR5PWKNvE1H4q2VH5GFg2CNR3fLhMwuSfOPbO
ANJ6TP1zKJkJcaW7dWBVcLTs7busQfjgbvDt6sv6Bu2rK70yvsE/uYC5Z3MQz5iN
11FWK0c0lKWJPs3nlzm5gcZZjscQI17klmZKtqDLMVoMe7HzZY8hhWpPDk3CvhXF
tdmOhyy0atq0H753bfBBOwGWBDe8TazoqN60l/y2iIPHGL0YjcsXCurSKvgpeIcm
yjHz0dssOcgVmgfASiSw9q5U89pgv4UzyOGSDHD34J8PN8CFPvKRslMnsFOvlQJr
eVsRHk2ExFU2cr6v8vBrdcwz2js4SfXZ+5AHQj0kVwpg0v/JfWEfNe5zdbB6Hpll
HUh4MQJWaYTLZA0rkEyYXUT3R17w4JVmHpiwt2Z67orSZADMRHi4KEaXRwaXPTOc
6SOdaF5B+o5C/L1Xz4EWwpbCPvQf2gPhENBa492YW21x+5U/MOkhXjY9rsXdRryU
2f543UvSGWYjudy8aU2hwDpOR0vRPbfyXwGl+zSSLkZ8CjBfrYsrLK+OCKfnNOdj
pYshbmu0OOuMBIZGriouHFF8DrzhccHkaIgiH6EL+VxNTufMLHHWhPqPhP4urBYG
soS/2BF0sAIa0USgmHm0XTeab4JJtw8aUkdMKLJHLOXFX4ANgiWtJzDPaxEGTdxx
ChP+aSCWTx9HSTo7pvqajDJGn9pxxqPGhFqfl6+vXFcyZDp60pmiAAMFfSYGCqSI
NhFS7Nfjvvb4+SZWdphBQaGY7dQNMGTKC2ij5aRJPJBtaHvAueLLS6NmrjjT9Whv
WBau3+hD9gVY70dQ8G+0mPdkyw1mDXb0RP+y3VWK+7j60lO2pov9cghx2bvp3DbV
vDNxievQsdxz0fU7HbNzzQL+LV9oZaaca7+SyLH+bqLRAAl6fd80FukCwUVgPyZG
Abpgezz/Z+fq25F42nADiCto3qaJuNEFhagQ5J5fPZ+kUmA7umjHbBZVHRvPOQ6q
e7sQfi6Ac325BD32hjrpLiaEMlcn9WE0Uz2FkrfVw4tc0iVY2xvMCgeTNu+w9Yeg
NtPwz8hMMVzSO3MTkaHa8lIenHodIjsYmF3lOdCjdXrM2YKbRfptgNxDtpeSQLnH
6hg4w+B8Idem6ZKO1R73holdnIjf8f7I1UTHuFFZ/ykhOMan/TcrUxtTteuIDEFI
Q1FKES0uqd+9ftI5O1XdpmwK6QoOzIntzVGVvdjAQAoXRFeE31cZqY94sqtMpTQQ
MTR2zZhKnxWCCNAR9rO6dRgxKL6UHiIEPbI0JDJvUY4GDiSc9Jw+Y17HbuY6uDZZ
mznROYLVhYwNvsbiITxhZzCMecw8rycLYaaqyA1zQoua8wpQLfW1FSk+VtIesr6F
nXbjbj8c2NX1r6IuQ9sgbx/eqTPBskgUNRzXPjdzwV4BY6iSPjisoq8/d0q+ZLnN
MRPSe5yWEP0w5n9IOeTO1BAAGjzH/Am8T8sdlIZn2L7X87jdIavH1mkNJZPKyu0G
GwPoypXXj6th33cJ4BAW97Owr0zFGn9P2zOu0s+c37Q4y8Gba3O+9aBPXwYfuSrC
AGJbKTVUlvQE01h53JhI8Tl2ktACh6502PG28s5CpSRWxpHbNw7+Vw84UBe48qGM
IBCMjvq2cxnSINaiaBa/0w0uvc54W67impytEWbLqhz4r6Puhhu1Yr4HH7OlEORk
6oig6rlhHbt5yCRNy5oICpFN+6Xv8xHrbxDULGFJeYCZjYEqpe8FQTOwq5Fw07QF
0Z8zWnHxayBZHZzWbUaVChtOf0rP0Gn1deTkYTIXX8/+2u5zWGWaopm9vHvkEx7K
4XPAj6hZ7TBP3rGzEzY3YuhnfErFA/qSN9iodjgId5vkWUJZSiL5XRXDyt/SMyXK
gJ8QwRJ5AF9Th8ZldkIiApspMjPnsA9VXH7ATe3+0xeJtSbQHQ/UNYRPLMYezhuz
1gRWzP8vTGOHTt48Gm0+JTh3DCadj3n0zYUeJxzCutSPnZy8COX1WN3nCXIpOZwp
/AAerdNtCSsPWLFTywJh+zcV3lafVflWAnbeH9C3p/8H8GcOi8/fEHV3mh7nSUU6
aBFoOoPDHPI2MHEBNxn8EOlHSS0oCBzhDeKqNiRkdlh/XdX4GWWUXg8AJUsE1cdO
RhBqAzf3d9s92PkuDz8M/n5ln9675UGFWZvbg9KaWDI2xttv8zFNJ8qA3qW8waBb
kyHgKv5d421XNZN9EynKMI8vrk470NqYJHrsi+Dx+FQOICdVh8Viqu1hb5faFBv1
3C0PCXDnEKycPTbKSKKd0NScEWoyK/W/LQaywWcrYXxqUmbZ6QEkqCiDgkZ55jCw
CzTxEGnd09aJpShrkZGsmr5WXdNYpqSWDKerC9qPFP2LnKZxoyJpeALn/9tWYfa/
k4x0ZoeKJCk2+6+YdwdwmhnxJ6YmqstFFpl6CnKW8Rzl6cLFKqkVQTK8pIK3Iajo
Tr8Yr/MPCYOO1608IExvnp8e4gtUKC61qygBxLYhqyKMwUvhXrZg6aChXMSH1n5T
6pkCihBI+nXPqAxn4GWIYudBGsj/J23J9/pN7yF566aiRK2yB7mhCMjjRiRWi7OC
J6P7Lj6MhHzhLZATRZqrbZW0ggCwjeBT3jK3ROwFU84SqeW4MCH6AMWIvmxslqqv
1667BKutEli2K28GGW7MWug0eD5hkpIEC0Ml1TxgXrAKWrKjhjaIujZEtG3zVzOm
fZNgjeCDqVf3S2qFdVTr+Ro/qp2eiSfeFBdBI3SwKmigYvdiQP3CALjohDGWEPCR
0c3yzob6KuWfUV+iH/odb12XN9XlEghnUC6dzqV2aMiyHIXWxRg5x8H3098uY0nb
3duXhF8H4mx6FS+PANkFdAHEl+Cj7NfgrDkQbGZlnLrj0rmTpsOwXd8bz4gOsLB1
uFxFTWeE81bySOgLEnK4XZXn419SsKtn8KYiFaubJ1ZwkKQjxnu4Bqk0Kszdpb88
HozUJGykClF3+hcHAhD/04EXkpSoKXMwJAql9QuCh/GrTUCGBRgvJzn3yMu4zIgz
36/hu41kUUZSmH3rIOtV5ARJkyRL8J89niSjh04vHLcvSxKJ9Eoeik3a3k+nV7sk
BPDNgYXBc9WebehIv2XQBjfIBf+QaiQT/bd6Gf4lvAE0NRbLhOcGQGNvGyur608z
J5il0rT6ib4ZNe26b5nfMtKuQpTWX1Oz7a8/F0jknmoTLnGAk2ym6045m+DFiQ90
Z5tTU2Rz/hM2Rg/q9oG+Xx57uTpm7eKisLW4LuU5EsOr8s8Blp6dJYYLKWfmiuAj
mZr/Yh3ZhmcernAymIWlWPkegTXHTrxoUy2kTf4h0sYQs+VxFFaSE5ujNUMbC1Yp
PW8q8xinUpUXz8Mo6fhEW0g6ly7V2Z1LWCu/uCPIgp2hYaNTA3fuEEh5JinjwFSp
GIjRyl/O1rXNN7y6hYsziZIxwkCbE0oJoWQFxI1vDnuiiRhHpjLgeVAJkT9tmSK/
gnPEWu66EXEUpPxFH0jB1zc4MVhEem/JPwuEAHC8cBTvTE2bMfX2HwFNIt49oDGq
XNeKnDUHHvMNBCWdXxuetXE3Mi9FMQSzqNqq8PXqXcViTzM8eGL3qbUawxEuoEZ1
eBevzrhKg8syKSplJLrHPLPHm1fbuX+cdjcUSJMOt0bpZG3LLHpD4tfhVMZD+pSA
gIIJppRQsbdRVrADsqo6aUg2sLqNt5xE5oMHlXIgfLCtKuQ4RVY9S7qygWi+WaEj
GVIu0PM/vMVG7/Rw7Dg8XrMNTZKF+anaMqQbr3XcqSoK15VxmwAkatAtIbuyqE7U
EUJTvG8KCAFseALGdvmDMUyUoMaN4MGn/VkxZ1/4iBp3XhjEjrXN7cdJSzl2/li4
RJpx5gwkL3KP0Vn3Zsg+RkBi8wEeyOpKwOD3JSpR65celWub8b+Y/Ft1MILfXtSD
0lbJchQl46x9PS4QHE6a5KVoF2efP5ic9RWpNzV6RGrlOWfOQxDu4+jImztGt22H
wEWDg5oxk2CCD+1E+CHOZJeb7T8an6UkWekUNFkPEukzQHwK8Kk7R1kxP7nQBVH/
ra9ZyoZzUPjtg66/DA65pGmM7vacpI9P0N0Khb3vJSg++JFKERc5z+5VeFnf52qD
rK+L/xghhXhfz94tRlvAfbBv8o1lYZ+V8NU6UYwuPs/CdfpEimI2+/6ZOmW7C9hk
d3KCnF9Rmt5uywmCSB2IzOGc2wxDEYc8AnUvyxO6LWUyWtp9UlO6NpmAlfo/DiWl
KPHocOA5798/SGmmo/gAQw6hz4WEVNRaeExakwFVbAfBQ55G+agtmAxs1gCM56MY
Kas4lmMDthSTwA9FhN+UQ1mZdWsQySjY2McCIaJYvCrIXI+jvCtF6XUqKJgsLshT
rnIJHAiCKd9mywHKzTNF5xDX0Yy1ALPlmN4xsWYTS/o0ltUPyGFpDt1z7zIkhbi2
3h6VFavR7961ddwR/bezH3s3IE1DqgSTDvQGFuB/EgEdDyQs4kv/DQlYUtvzXgIE
RDlmnJd7G8FNNQfhv3HNXZT4DTJYyQe1bW+x0EzJXjr19RvZsD0ogEWLBirp7AiO
OcaSRpzQfLzqF6f8gstUftMoXiHBN6GPnHsKiX9VAZKinzaVe1ECJevdszbeP+1j
/yB8FfK9zhrWiLbtzuRmmIE6s9S8rB6ixdHjiXuF65eLq6qvBRyz95jdvxIX6Au0
SUcn8M8LBfypIkDUL5luIEM9fWz2fdT81PNx5kbpbSyLKiMY36f5AqPPY/kh0RFi
aOrkya8joh80V9BJJtdZYFmPAWVa1vFMbCIt6tycxtluM1HwymMfm0zxHWAro1tk
gMEatenVS9hkQ2d/oOYyMWPvFe5yDRqWKrqyIZwke5od/L/dvpRKiAPOpc8MOsEx
pe94pXmsufJ0o7llgUasBKIUI0f7ZuKr7bPXFHOtNy0Zyn99a2+MpTFBrbqr+/Bo
sim/mvKQHniIalLy6WZwG0Rf5sASVk5fWcufYowXAY+9GgYq6NTvZ1Glu5r2dwlO
S4H+bL8mtzirsa0LVaU1mIWl67CUT6iRvAjawsy61MomfdN7S9FaNIoxbcbybnA1
fz8T5jSZfKcxym+jcZlAtVeue6qYb/JCSPGF2hDKJgM7xMqfRz4pTAYbmfc81h/Q
tzLJqxzM2AmrciFPdXzUs+cP2AnRtwTvSSzl9LftV+N96cpcQK0iTvK9uUyNCdcD
HkmWK0P4vsm/H796UGOxKmB/qXSAZmqwPW0us/rXgF/CgWmR/4iXOT9P6ZvH5d8M
x9cgbqQoEa6gWMAIN3IdXRG3dzd/7YvxJLOOgMCoxHUztRSt9PZG/9jy5nFbki/i
TFbHBy688Lp9FgDsKZGhxKvexdulKIKlbcZg/QdwfCij0D1SZ4Nh6iytX5yPonHn
QhUWvb6cy0NEdomxIy/iCfzzyOuUM/fcwN+0165PT7f21JihQauPdIv/QMT4N04a
1s3+qdeoaNmk19rrkSALjPVI1Xamb8WJsgqvaQR0GOru5BPDFZjvZ/4HEbtS7iqL
owKTbs4yWLU5D6m/QBYAfr/Ped5g2N6Nz5Fyl5jkmZyOX55KXs4inNTW1wIca/Kj
5QgVWQuoo3f4BnQYAW0tDqH13o438am6n9XhB5Aorp8v/W7Criv7+PEsdTCV3ktT
zm+pX323MB/dAGVL93dX4bfdYvU5ZoRQUM90dwv660LyXpJ7FAEkvY7k2p0G42vF
NSY/a8WNTJvAKVvO4f0qsOsaICAhtezUQBCAS2Aunn8Quqxm3RifR818yN9rl3PI
O/62R18Gm4YCEA/jzZIXc6y45eewU5rZdYanHip8FFoyE7nFDysyASm+MLdYyi21
t1c92363VDVSwn5V2ilZgaqWFmHZl0SOoCBIo99fiGWB1WNuMeXD85V6Mii9R3xk
U/h0MG/BkZeubmQanOdoGomg7cXK+xYTU0N75kYiiTmYbqwz8YTPEMDuFDWl+D6R
Yv5nuZJSURx0moVIQtsdpxF3fZCgt1768k7cIDWo2KGUp8ILxiqA0rN67lBYpDLo
Yc6yWeHEOWR4/ess8QqjRqPgl1FTzJzfGcZTgOvlarStLyFOmnHAqyHVrZ6TdhYe
CLLaJ9N4tPXDrDmJ7JJ6oSDBoweNVEX8s7PtDD+B1FSKQgBCjDNpQGCH9fQEdxqh
WQZq4XENxavfrpxQHav9Mf26IFauZqvx3gkwqy41dtBMykSnwBALXbVss9kLZhkS
WjGVAqcINAPliQBDWw0H/fS3PbflDrass3W/ag2sntsXSDkAuYqTkeliivnlVdka
bCUxfntPV1IsW0SsDg+xdWyvDpebGzhC9Ls/r2Fg0sZIPuIjIrvpurkJ+q+tn8nO
gCWOwLHG89NbKXFgnUCqMo7eGtwxF24UYpC6f7RlKptd7rowHQYvojz8io/t8lw0
R7QTcUAgL00ssOb8BfoERLrf4c2CNC3cFSbgDB/9jMc8Dmdsa0YRPTtRZrMvEW0o
PJmdoyD0bJOF4GCSkQHyAeLWUjBrR43IrxTP/1ytPZDchsAYtUxvqSBufC5KILJo
VaorlfznUep1gcG4x9i/u3QqjhCj/Ur9862AENpHpQStRPOQ+zyp5SI3b3oXlHTy
FpD0VFmqcGX+gqjClFkVgCZhm1fC43mbzuv7KoE36Zbc0tOG1pPBDZoIRviEwp3t
rP2ArqV/738KSpOXD50VzD2cERO+sgmRno/YN8MgZmnQvnlcQSS3XV4cnzhsIrGd
OMIDInsjLxiFn0NR7ByB/QksXJtQLXfpOGFwqyh3C/jVl7z/F6D0fnKhbzbvPxVN
pNczXgt3mhcTT5WlW0etDboCdH95WrmjZqV/k6mvDKKrwCRSu84ZBNzMmM93Dj+m
87pznpGLG38S94etdlPxfKiSIgLRmE0n3kXu7nNyqHMJGDKVMBMSZJ7kNV8uabra
uSaeI/GwQJDPVNTiAL6fAHuUO8TH1tssGKaxaNmtA/W29rW1jpwrzrf33EfcvDQ5
pN67XjnnOmMUohZ6TagsrN5wM6KHxJaj5CwnGMKDpFOqgPodYTLJF/K5JtJVq5Xf
mqkevKCL9DTylti7O8PIpFfYQE+pVLRoUZPQmADQVq0rD3FPGUnmlJ5FOBzyd+mh
XMYXOY+3fLjwISrjoVQaZfEHFqu5U0VrNiWQaIDETXDoFM3yY1Bc1sBuq8Z/0wn8
FUfKpWcs9MvYHS5bNTQz51J+Oll6pK2yWMzsIveHmnZUzhBxTbn17EJb7jClPdJN
na6YceU455Agyp6+Zd+HD7kB3vn/OWlzMFMppJmKPxte3LP/FI/vVavGa6ji/nRU
9KOjhP94WGRQBe2k7AXenBFj4WQAuNL1+sUUYe+xXmCtLCN7XAH68ZVyPWAOl208
Mf1Mo5+FUtveZG5R5Qyhi7J/2OY7+KDPjiDX7dytmP3l5M6yKBd1Y5AqcrAk9ms8
zbJbE51bDZva0L++pebJmknjY9r+8Y1TlK5Qi7ShVUC9mBprYDRIUabvi2GYQKjW
giKpNF9WJsxuy7SDVSyUi9aK73jdkiaDW3D57Il0FPiIe0ZwYMv0Yz6cRL01akFU
Dh8SDXzLdyF+/z+fb1OSvzgEDOC6kmmG6jXJINscxEaiLfPmavuaXs6561W4BV/R
dLesr9IBf+zHInrQPNlOdbNhmeaaH2cKdfB95QDoE1sGimaP7EJlfJYVe28CqEkC
Hs62UTySUXCuyXIYDvSRcrig2Q7UZMWFHLGYx4QP2QYrooZifkh6DBOBLV2wOu1I
xsS67bumW6tNpYVffEiTSq0iHRXbeoSCllYrWfpxmfQecoRaLBB+6aVUaRxnvepD
oaVGAl587y6wsz9IxGg9VrGXrZHUkZEoUKSzj2m5IFdz5G4RwuS3w2upKNwh9sP4
ullt/+Lno5QmwvUqA2V83t0kep7ipm1PR861DqKBZiEo8bRQGCX1wROEWJzhRNGJ
HQlAWSbYbQ4iHQqun8l/j4Vs6Jbuxr8yaB5Redvol9cYS56lXaWzYf4BpL2BMEUh
isj36HpW44aJ6R2O2OBebm9CkJT1Axtelaw/bwQr9AQQCwURbghhxJbUZ+8atem2
FnNTIMFyNtJ/hzaZKvbAXl2I3o8tl0MV60vjJ9U/zJG596rEgs9TWSdTOWOCySHy
+4FFUnGmX/XB0AiGqJ/mRskU42SiSIL9tZvEzPkaChW58b+VtM6LUE1BCCgi3Fnt
hlFKWUwv0S7yG8rFxG+Y/OaKuHDC01J0tIhaGGuFnrDOwl5I9z8tvnk+dPkuFLuI
zI1aYqsNaBljQRnTcTHt6rcRWLVoE9y2JqxG8fttYwhoxCou+y51FDkWfL3WsXvO
C415wZoQGGNeSCIwIxUSdhvAHAGl9GEH8d7WnD7WYP1lvdtlhpnqNY7Engpn3Rkx
dCMoJRpOd3VsuX2DwLmrUtUb+VNuJxbyBKMUNevWTD+BOG6HWU2QNs4uA27v8jMF
5rHhp2rrvjijorQQ8LksA2HpJoVtCV8Nf6Zf7wMmM1DYZRYv/7l4HM84muGzbdZh
ETSsMKkSLsUtnjra0SIwkDYJwCiC6teOPhK7EIqTNIOVHQTjJudMIBOfWRNI727z
pxxqUIJc1wzFDOSJKrLV/cPgK8lIrFXLlZytzJnLLan+69sswAonG3iVdELElzbm
yNbWFhGXqrvsKKXd8ydnrJvxdk3SDU6GzO04CXLQDkVt9VDeENRZ9EyVkfvS3Reo
GwfxqBJd2vIBOVFcg2mw+b6O/5STpJRM4B68cwvR38g45ejTlZF4kemuJkwCTfCj
lTfuSgICH0/jH5kLfSb7ScjMw4LWiIG/JJw8CbLfDwPa8ayJrWGieRp5Ys2xcCWK
GJxIU3WBe89MJkjK+o9+WqpBZ6vUATf1yv1THSFky9u6zj0y8zMK/ZG55UfwdeFf
QdckEvIyGRHBII2x9Ir381s+liSwihlCAXJl2+spsKk87lCBDz2nqH1GiCTgu75W
keuzIZsnTHd85PU6RGyNofr+eEeLtR+rJIMRUTnZn6lusuvUEHDmS4Issf8HSK57
7aH+YNPRuoqsXZL+MDxkce7Cdf8oUajyWmq4XDCL680gVES9V0l6Vdh/VVp9BObN
qB0quIzzzRwtsBvzMuSQUNz+NG96ke6m3PjKvHI8NH/glm/hZPbDVtA8NjZxRYoK
9ZPZKnSBReVNYFzXP+5iZqEZOXjTxl/4oDecNSG744dXRxDzMeoLRwYPwH15aMY4
VkPWFh4fc60gS5XtSEFsuJOv3xpVDSwF5iBZRhmimde2u5qO10PurQpHcT1Y/eDO
zk3q+DYRw5EszeT3jPW/vklL5nDQrc8lFXIaD2ulsjoHihJ57wsqBE+hN+7zQCek
YUNFmmKuKNXBYTwFGs/kIvwzisCfdiKVk1655RCepQjAnbZHf5UKNDM61WAYQAZL
g9KHgbKIgjC3EO+5R2mcwYGD1X7Q+6tw3b97EjuGRA1iLJVlDORShR5K+5q0hCfi
FFnzuuYnLf1pbKcxVZsKdLL0daFRtwrWgG0T97Sq+FO544xQFF1m1A6X/F7rxrk5
44u5vn00265rbMOzdU8sV/66FanS9vCzn4cUQsKe8iKma2PZmCPEw/G1TX984Khc
8GfKE6Enp7QSEjotqssoStYoveudKtw3DouxAxjquPgolvpjNWcv9Qb3P+q6zqYK
NCIVYJbOdbHxiIJ7pu1eKPtqdXj/RmGglSzIZlg2BwaYtf/QRbUvFC/W+64g8dwx
U5qgPZtXmgwdrLlMDgOsQNvbQVA+wBJVZsdVSx110p0O1fec/ebTsVuThfp4U3wr
2P8G35nXxRHcsaDw6+6b3jOKf/nJAXDtVpkg3WbSqvt8XENmHOJ98Ejmx7CjLn6o
`protect END_PROTECTED
