`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRUt6KtBJZ9XgKOwYrw/ZOKhrnr0e15LDEf1Oa8wzRVqnP9fkuvWoag43jckrMkx
qbVUPfGZ9DbZvBPV3g5voJj7S9ZBOiyZCQW8qCzREVFUTJIH5gGg+J/8ZbeftoH/
6Yj9bhGT7m55SLSgKe8bFD6NJDVXB0cQg3tFQHzjOli9PJLZBTn08JBo7Nkj4Auc
06uLBi3mK9yrgwdTwo/N0cN8UTzuQh9BXvRwkPUB/lIhvuLPC3Kx/Q6vL7UkpA6O
S2hKjHZ3VKthjrSq/zrb/t0zFx3GUyTi55/UOYk9GXgy11wZ3GezjjYxeSz2SVcB
OxVSRytxAfWkdlouF9JgMA/g3EECMYu3M8exhVGjDfOH04jooqAo2EcICAk4p+51
B4tLIvnrFlgJpFGPwL8Tz/Y85rA3RikyN0Iwyz+w9t5DW/S79SBI7IIaPdvTlb44
DUbczwOEcqJgQkEyBzFGEqH519vqfcjTN1b6jOqsQF3grGFX6vycGGviwTuU9vij
S3XSEm7zhRlVvH+/2yeEd+c/Mawy8ErsYo0q8J5d+lysOi0MbnW2iuqIiTc7fArV
yX+15i7l84mWAF9wS/gMXEdauuv2JQlSPBgTjD+HTUXbyjETk38B3o3a/HIkHuTA
i0iegMMLs7FoKTDNMcEsh970u0rf8r6u/dtUCybame6jtHYLFko2b+AhKu9GmJ4Y
/UwD7Pfdxez1NW5cohhBXFAPNP9rmLPwPfhasl8v4U7HbllzLx9Q3Y0fQ3Zk/+OP
s3CsvDp7Y0YGRQUPbMJXaXY2k2kEumMkBKlK+TH/xDnvjwSTXuYwEUNIcyk3ypaN
3FVuq1FVglYFEdHFyaBR8IVn6hSwO78Wd88vuzCj614XogZ3lF0fLbpRDfnotn+Z
xgoqgp6+5kz2iLXSHmaejGhM/9H5SGdcDU3Nof/yIKs7wBqLTdXSNzww+bOASD9x
Z5Fh0IfyIcmIIk/RdhmJK4KaIcC0xoMEiTKllJ+7iXsrGWDsSks+dS6Yo9afc4kF
z07Yvx5+IpNaRsPBkVBvllRWFQ1XlRnFschlKknj73E13TXtqC2kaUR/e/iYl7dF
SR+G7A9ouPlkL2btbKub9iyYiRYARxfuEWD6lweiBLgqlT9+q5XSS03JfgCtT4rg
vWTErqyh7RSR4TTCgJ1GblAq9eXe4SpJn/vIj5jG05tw9Dvr410SnoIAxOepKN/+
/AIz34rZzFoOYJ15hjUUYNyrzLTIEVv1vkjGEV1u7OydzKNu9DIpwng1kuEzVwzR
/kB8SbpexIepLtcEzmFJJH3vnG1xyTKkDiLp73FX7CQgNCr2mwIGPwsby+udgeAo
LkMVPzyu00eDLUb0VQwESUKcqkUrAZ1h7s+H2nPDjKl1Y2+Fqu0Mem4XLvNJJOSl
1wb1M8GX0Y04p5EI0amt/jbdtogboVPli2fSH1qFtVj6nltz/b1rBO8a78RDGkm7
BWCPNFZEheG4U8xvVNepGCanvrDhmMTF9HUIB63Z9+gyKKXjjGUrH2YgSRWYh5kg
LeZvy7kqrus33pAHuyMlnRWxTPlAp05x1DLeUVHrbh248kuJGktBMmNvIod+plS9
wLmLoyTZMdsAcYJrgbl5D5gWpiDOVij/4xA3PS0NaXL6IxDzM4WXhOAE4KbliE4w
wLGUuECnVwTOFgtTupA/0BHnrMY8dJOVCA9wSnf7HOlJ1hMSJSMJM9c+43n9vipa
ud5aSTnCqU+wGsrArVW4WZPGn52lfGghbfKKBTTg70dF6g/7hJbbe9eL5PROvS6D
yzyQ+OOladsDR96oDu9dhMCcz64RdcuUASKmurcuVxYSc7Zma7XgP2LWHla1svdr
m4z1fyI+RMtrbqWRMXqo1+fELG+PzGdf4YZR3t6L5ce7FiLSCRgWKKMzKZ2N2Ekh
1Im3o1Ka8e4Sln7OzrN7ikw4du+e5J007VrpvpPTOmljLGvwi+k6wDvYS6L5mxH7
HMNX9kRbGPEKvAG3dw9KyZ/NLTmhxKWPbJC+P+661f/HxCFyn4GTtGC1Wup2zZ6u
Eutvzm8vmtKeo6B+GFuUvzvaXtkvFfmW6W9VzfdNKsfanRmsFCy7d44HQrwgjnZr
Yh5s5dFD0Th0/3BZG6eEbp07/vR5x2Wd4y5DAzQR550EB8y6OYLcL3BmWp71mPMQ
Xn7Z9en4TVUhEzzo52xbRARWtmixSr1h83S040uzBmL/sJNrx9ELFXwP+/7Dboui
eroImzUi3utEShQ1X9rLfDZETHAcL4hvlryHCvqSYXveskht+GKSA2B2UCOZ+jUu
yz6Fv26jcTYJsYeVKvOmMTwTUWSDaojvBpapSssXYIs850cINPun9+7QvL9pLAZ2
qY232XPAGWboZnzawvve0NFtgmNY+Hg4GVLT40A147oHaU3A4uy0mXl43u63G3ht
S0iZH/nmsOuw+djfT89o42KjJ75T8TjeVrPk1cy8JXd1aqfraFOxCYYNmsbatxkP
//a1tQnQFkWQDdYqmDoP/HSMgujpB5z4OnPZ6MBJCrhGLyrYHP8uHMemABhIFcaS
uVHxBkHmYKgl/276y0RxqSMxZRd8DrMRUcDp7/S9EcisFG5a0m7m8qOAFMIey9qy
OBSeSx9V+iN+/e9TyNduQOW5iDdnxAHeoZG1P1SB5cEZxmWzHAxiJih77663S8+V
ucaIQOu7fedULMlZkzDci1te6PkJvL+y7FakygJtgO9Y/XrWZ2KUhY8pQagUvKZM
XXrW3dNmn2LOLrUnWqBWswdLSBJkN2SdXSKcfJduCgfX7unxgwfFF/ih4yoOi3S7
WzpH0jCi+ZyJwfNhQnACoPE304ykdd2WjGwzfca1HNkgK747tbc0cwa/Z57BNAbE
PjhnuxUGUC6n8mXyUI8DS0mbW0YV8iGcafKATOSoQdQ78KMdBHokT1msD6lKxKiW
DrEXeCW1Yp8c7jN9shU2YjWO44i9Ogch5nkaGipfLZBUnrXsTUbkhjq3uC4TowJR
de4ZmIhc8eHtaOxVTqW5QsfIrZJ2X3tlCHiQsXfcl1nKLmOmbW+g1pokSvo631m/
mgfob0MtTiIONFlj3o1PsOvCrhBIVGhLI8439zek6yToWtvtbb09AV3ogOCkfHTN
UmNs9SmJMB2VJsNmjhdjsJMB+6QZ3r3mQU6olJtJrDFvRih81RiAFuk0zkzag6yY
GaGrF3eKIqoqn2Onw7PSNKIXA8Zm0RJU07fCNpdLwEdnKHaQJy9s90kOrbIPQybT
`protect END_PROTECTED
