`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4BPz60yIB5df0uq30Vfv0Hw4mAFDgrWuQgjfZbCOr1QOnJ+OCaTIVL72j3CwQKHd
p6qsWgEfU7bVVE78NXPx7kmYzjwpM4NJLhzU1pdpPbWs4bffKneAA7tqTOnOxq+D
kAxNeyL/Xqh0c8rbi8NRjZGI7R4rvKD7q0R3bmbRLjJuIExWsPyse7IDwyQNmoYw
JaArHNcq46qgwda0g0+zYbiA3Gls2GjgheZvH2fUuqVSKS4lOb4dkpiY7y6M31kr
v1XudpmMhuGrRypDklcKtHkeo/GDMaOdf5LkNacHjSrge0ZEi4vpK/A2IKmmGKZo
fc9TVUZCXK6E9JU6Snoflqlhn7oiOrDksS91ZS17GrMmfFIzrZXOV86ZrrxFTP4q
kKhz4pGfEfgY8QPE9cyxfLP4h0YxN8U0YVP88FA71SJltdJ99c9/i8PZx5L8WFhe
rbH7Kk16LDdD7tPGr713HoQi89PD5B4DKAsH0MDebILoA87piw/u6BHj5feLm6H9
J39OJGf1KC1yWdLyXin3mTHcOyPtiDbXUChwE7Wt7X2jdyDfPEsmOcvwlBfmjaGc
W18XGDz21j0IoI3a9+VdLBHRRsuuBbSUA6QV5ApGkEVsk72TZm8KLEtqjWjhgDet
XchVZzC4oEzpxUswUYKQwHWhE3/z5Ano9WfrPCigbuE=
`protect END_PROTECTED
