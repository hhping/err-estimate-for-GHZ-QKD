`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uT8Y8AKAirLAqQaHlfhzjhpauVmcu6yWYefAes1KEgug2bsFw12g2ONr5wU0MUWa
tV8nd3vhSOZ2zVwT3u5zxnMcuSvdJuFA5MU//a6Bota6ikah0i4VD1HneBJNlph0
7avlEh40xgG4Lov8lv1VVySomu0N6z4x4HD6010zuQCBP6rWruLaxKLAkfYuJjhu
/Lt5LMmqafKPqB+7f/ZdT0Dxzoh6Mn/xh1tU6SV5lYOmYykFXXPQPFhm38A52EJ4
+eDNdEtwQ0v1UPZo5lDOe3Zg0H7lqZt76psTgpiro+fCx22sx5eMht5sBuqQDRSC
ojJ157GEIcBhvpTZCYkMdzwjcp0KFBj3xmXsL/XigQ8dc5Hh+grG8FBq2lt0z7qF
Z3Ek0N3n5od1EeE9hEiUH24fRC5j4aKl3A+KWTdqBGdQfEpWNACVScBu+y1ETcN6
UQkroKDIa3y5xJOKt52ciTI1o4uCiMk31Lq3yV94MVIEbpVrcVoBZg7N9I3+GaI4
gpXFqpGs3Kuh1wo8X6EzUy4Ka8qOlGMF4TqvcYZSeCf4n1G+y5ydRjIafZi8BRsr
XijsdKSPnHrD1OCKvssjQRqNbocxbqLf+N9/gGvQhn6h4OTrhgz5mNoYU9UqK4Do
0yx2M/wAVioZe5ZOFIE8V9I12ZBlSCptZOb4Atvrsa+63YQbESqooZcwjkLvZf7n
38KxgXJX9VZtuScD5OZ2vXqPlzRR1w4GLinpBXvm29A59piiNpO+n7Nz7EX8uLGv
3Ivj1LEqijN76QjYezbAFiz6AKw9zx/GWpCiSTRwG/hnSCabMGtjejTwKF2T7zjv
iUM7hFuDVgsqsjd4PSuHIBwb97wTL9FGLrBd0Uv0OwfyM01/Zqdrtnytk4bOs5Pc
+Djduh1itX06FFv4bxgr93NDUXZwE53Jbv5k257Z1nKa+jSDCerLGRzsZU4kDq6n
sHbiHWnakNGct4fICbcXgTTq/D4YeSpsj4G3qd9IV+QlR0Uz7IqFXNYXLx90oBwx
wOFdtepWtgcjC5bCZ7Kb4CKLqLiBVnJPrDPxReo22F3PjGHR8QatFeD6cFlFi4yT
mXHUUiieuEKSlVwAnFNViqiM7os+YHrL0czXuaMPCYXnoISYkpgArek5LgcRwfxn
u+MqIu/ld5X0bkWo0Y2Kad6DOQKwTmlVGWpLVz8VV5lMkEMZ+RM+PCG1PSEK6Ggb
ZWN0YOXZdUy10d5Jfqm96SjkZRj8TSIxtTlgsoy9KjmpKIjLP7dJNAXmnIl3JXCH
tNHSuEeZ5opVN2KQUdPgIiJgJzRwh6HM/Gu8I6LU+HdMbTUw2iFW1JsOOQkaZsFj
UPM/cW4D00dIBkns5MNCEPzCdaeaVVXRCxrtxNf0nRQMrFOIYOpi90F0IP7ESeRv
hyu3IUzTk1HS1UWxNfKBjA==
`protect END_PROTECTED
