`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XX3Pjm02eIHG3mXkGI4wRbeY7Bx7ZAgQcKK0uU93xuEhbYFPRbcaCWuYZ4ZyaYpQ
n6jUKvtO6dOH8T4Nw8QQdh7/BlReoUkuRgrVVFjOUvITANbAjdQHJN96KwusDBvX
uUBp4oiCA7/xIpxQ/NdM8X5wt0LjdfUByybeAncv5e8V6Tt4NeKYeqv2sdW67A7G
Orc6XQWGfXyGuJchdnok8arnCRPLF4Hrv7uVXlms5GTTiW6EXhkPAu32TkgegIwd
eLXPaINKAZvdhnX6We2MBSRFvePaMMk03nsBhre/eWVfvgJDKhGuBAQKKRrhU9+O
t+xv/uCzjfZxRgRIGBZVPlP2DphU8rsCdlSgjWW4PuI3MY2Ts63CLEEKFgH9Kr++
TgpNURLmK3F/jtblVkSqBsP0Qw+cJP/DN1z/ULM7qg07oJWA1j5QofSyfqUGKr3M
fa27tkCkDswOd2RLKYg7A2o0aTfpFQ4E44psWwYTFaviBsW4sVngTJg+xPqEVZQS
dxYXHE3aXQsKrGRe/pIynYC74dqomE8wTWoCbGZbFxhaJtRQrP9uTAA4G1Dev/Qb
N+hK+R49KOXs9obJK7lANsrlGSaW+e9T3G3sEm/SLWuhJbQW3PlBk2zno0pEtnBg
bzUFfcAhbsjg1UIf84XIYJDGCIeY4gLn7UgNBx+4srkGqAdAaBhirQ5iUSXvFqxn
AGBdmuiHQFmF2ksju3d6p6pDQvg6maRbEtypQDPR/3KlwrthDlGMVTcOqtz8OCQ5
/afFRbSH2zKvsGoOIjo5HjtHaKHG850zilL3WLqVxn5XY0GTw0KqeMsetvFyUzda
Ehd380Y5nWa1ZNm8JFcElBQj9LAVqcm73jvVHRT8VJD9Wyje6cLmZROUatqcZ+RU
zQA5GeMrvOew68Aezzk+ZjZxZyCutxPj8SXy56VrJ7vEoA/jLUVgCDDEpwat1VJ9
0lQ8xy+h3TnULz4zYmW4/ICx7+qgZl3DDHTC7QUygcy8N8VuLRnJVi5GoUMHCuoN
Scr6h/E0oUbReMmOY2qirgC5av8bT0N5QJdcknaZMc+kEfT3hd55qj5pWOHh39lp
YSUdhtoZe94r5nmeMoysJcuDw2iEHfoHEERnO+hj8Ngoc2m/gbEOFrQqTyyhi2QG
gpI0tSB+ZehdwaVNkYcEPjG4pAsDBKKbY5DhSbLd2IF0FkvJmILiYMpcRcNB/t/s
GhyHo6pIBAVOape+9CcxOIpe6Dz3s16UMYVqi4KD/ejPsYav720BZz/QFXWgPcWI
g06ueN7fpQV4PzVX//h+eHHAj3uiPY8xqXePRCGjxhI2N8D/W4O8vvM7uGvP1qoY
Ks3lDOm5ZbFsEkILBPt/R8jRbIK/DjKtGljoCpnvQpMXP3OH9Jp34ll8lzhVvWRL
emIJD0aMhIoUpnxSpCNP5xQ4mnR59ODwcscP/ZjAPtTsXuJFbNmXJCuvCPIpvvEU
g9FUv2ulW33bwiQOn2HYM/IRjRPyvncMIypV5KNpZYboJfMMgqO4LREftzmD1Dph
kTs/wrU2BCJfzeA8ut9C+Siby6pEPnBBPB9FXA1hdV6xesuyh8DhTJ6zcwUW5fYK
m7cpDY9xCsvej7E/cjb4F39C2tL2wkJYprC3Sn8u96j6lIG0KJ8c/inbzLo+1RWC
v5aZe8/6cN5xdzl3eJ3Ynhwo1QDLHnK2St60WkOusZfonqZ1Lij/7q/se9EBJyzc
hNtNOgtcVqwpS8WLeLo+sTLcA2hTBinneuj8pgflOCFo2d96ryrqQXvXAGqmcECb
gH6hNXeqJ8DQsIqcnJpI2lNbh2KSmy/RigCB6C00fm5G87qixlP1v4Pqsk3m+8xn
OCOkNzzqhdsZ5V3X03XvCW7salBVWoGYgeWC5tL5qDl3lbYs29/kEHFU0Z0zcLhS
SdNyf5ztvYEFkzW2yt1kM9zkaDxv8DNniE9LWSXZElEmeEll8baZPDxuk4MT4qd2
GOlGg9Wal3sSdLA7pYKFQwtiXKdI7CesmvZrxEBSDN3YL4kA/2nPLPWQzT5Yl6LD
jUqx2pbah926h6ztJBFV4+FqHjSy6yrve3gq4vRfzO+40EhYd8TIhvbeeVm3hVwF
fiTfHKXsn1AZ6ixtmcM1EQon27OFBBwibfmJqh6Djoc0SsZFIhMzioKP9K1678xU
KGO1IzI94BmC02nbog/6MmkJ/RGpfTCQrl3VqCIfXt67JMbfV5P5gqQLfPM2zXHe
DQGwfHdzIbOobBSGDAHFzkm+Ri0nzmwFaJoz85U5wQwzGiWxYFmxEd7feGptpXFI
husyvK4LtDU/01fmm7we4+5Hq3y2wRiVoFEC485PJzkb3x7ew4T+3OIfuZLOFAbD
nhKqSIxlDn+WCHJCXcbEgUINC9GlYv8YtiQTyaNAYGdv5poaLj3e7v/5CJUEgY7g
8kXW5bmhbKHys1Hhl239h0Agujlz8ptkNToDEcB1DslA5rI1x55ohFnhqnzNNiaH
O/+ReMXqqL0UvPJzkc7MiMjxvmtXXDs1120pp/PzxGFlU5xzAwR0CxXYX0abUi2p
kt4LLjD5kXdGOCDIMa1RQ4VdigTWYE3Mo8yH5Z2E0c6ff/0rpqNhZj7HRhUwgZ1e
9AEBk4nUhYiCJUbXh0up59LaM+xtyDQlkyqZ6liD6ogdH8yq6tQGoHzhiXEkPmWK
K0RyFmLqdgmxw5YWrj+uv+EiiErkNjTIHCbWbhsC/Kyry80DHLJ8tp0tXaoOR1SQ
KW4SeucBZK5snQJtCknkcffMyqjGDA4PzdT2X67nsDnCVQ7NJtXtSuRDz4EIQYUL
cjrsCE1DeH8zLFKU2zUkW4ADTqTNKArnSoQcsOapIsWaxFdoTsTqmIkApsr04Loz
2Mi4xBKbOCUbPzgmGGBWDZfekZlw0C2VX82OZivIKDr0pCS0mmC4UImNsPh4EBKO
oncTtNzxTipMBG+25oDahxOoczABG5xSz/2l9wE6VVqo6Ezl4aSEeWwOGQFnOAgl
hpkhQhakfEqPlDM9iTfj9XOlLe8SHm70CJoHyFOJkSV4jxA7hySOGXxpM8j+8ECh
CM1TW7QlgHb/6rq316BE4CeApUzaUsUWekHUocQMjq30zvJbwIfHtuh61OYmo3P4
j6gPKbIHp96xH8FILXpi2XsdrPHsxdjmvrz7HdfUiKlt+U4NzauTyWwvuBFMskjm
6vDXlc37h4hkjKqbMDN30VIIlk2bjW+8pYV2cdabKlsj7KcAA1qTZ3r0b+HoT323
3/HwA/XiJo/o29GC1kSCR7mjXcY6fBSfQTtOsQvhPAAGoNQJEaeps6L6Q1y/RSPg
cylswSz7jl4q5xAvNHW6g1VB7ZHjIjif6wbsigxVNMjpDVOIJUoz6h6GTCQ3tqZI
KSRTSsKV9zq/U3V1rgFApw5+VcslM29eOYf09KiI/bUULFyNNDt5KRjSm+3R0flT
GYV+eCI0IhA+n0KiYj41eLs9JiLMP2AM8MqtSo5zVrxxlpm2Tv6wpzvHyKN2ryH/
GUld0tv2WDK8t+FE0ukM4/JE7kyKWRL1HHxfQVUR2ST2d9Ov+M2Y0w1MUjSOo8sU
kdWok6As030p6DRYJWsCPhHtbRZqStSV+3p5p6WDYBdU/jjjSaD/fp6aT2sb1JmG
EbKvSImrJfEFWQd460iegSjRMeGmd+nZnImk7q+e24d4Snr5g4qkBPIEJgL7un04
DlctWxV8cvUNrS5eTNA8ceTe3qfaGi49ddQeplUua4/hadUshufnrbrzDSoGjQUj
1hKxZu+D96kMvyuhE0zuMv87gp4aXKmjwwZmlURXy8MZK6ceyl3C1NLVNmo8ng56
fFbjLnVvMCcc2wEiN08FIcNtuPJ3UOLpQK4PyCAMdsPXNKTBjN8rmj8AJ0ewlWUT
+hcm/eI0wzprUsA1LdnEJfAylVbZ3wm+5T+y8/JLL007h0aG/76A+ZL22bxtRjUl
uAkc4hDiyWF6AraRha+aJRLdh09McD7WIYVpz9aQmjh6hkTTRgQN/qT0bYU0rt1I
12km+BMZRvX2gHwvJvjlnNtgAjPR7t+jcFx7o758+TUnShfF067qZlxq2Sq1HYbE
xNydlCNgdAvSQhpFl5Sp9RkGp2HeeU9T7EkI5Q2vtci/p94sf7HvRXApfXhQj6rN
EgAtmVzku3O9l8mEnB89ijTM0isdLe15flocUtrjDyZB//tWgQv28ezn9Wlui9uZ
DBHFor4VwHofOhcI/DfPsKXJ7Ft08zZZKv3qC8V+eL/N/0oAJQJl5p593EkEQnMV
ncVhumyPgrbqrt5r17MysPJ4Sl+vbX0HEiOD131OUFU0m0rjL4ifud/xCdLL6gF1
LXFX9Rmdm/hx7FzZrLua71uEG/0MqKtEoAEPERnqeTVMWTnB24b8eYJf9kIDcsRb
WlKzooQPCgILF5PODgxGiTBsHgOJXsPQRHmwswd/31B4wceBgM5WLDUk++dJVTg7
dGKMJ7REguNur+jPCN687yi3/sok7UsM8FikuN9dT5oclPqwC8nWD9755dKlg4tT
hvIu03LoRkFLs0mcpts0t7vM5cE1pvEg62MGUjHPIe2K0krIBci8dr9+nTVHh6F4
3AcKYwatDOsbOZBJeqsXEoVs2Qy68269AODd0K+OE8k=
`protect END_PROTECTED
