`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IVX8fKe1DDR0ny4V+gZqUKbA5Msz8x1rithtL2T5voEtVf/3jRuAQWkCNZCe+Jz6
9qZE/56maU7kkpKkvX7Q3yPGRPs3U4Sfy997jBd3KYVk5vCgY8LJBWyQCrALZ9eb
9tzn+a2scjkzErEYKlk08LtLOW/DMlP6cCzW9u4xFcyYVMFoStPVkmqqYr8RJ/j7
`protect END_PROTECTED
