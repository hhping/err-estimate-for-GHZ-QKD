`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LM2VQ+ItY73eV09BsqTVx6IGNedh3tppGdTh0GhBVkb2O1YCOGaLdgGFNK+mseIT
dr0Ibj2FT6vE0xvm3U6sgNg9pZP0pb+kQn5aM/eOmqRowKJp8t+W51WxmU55HaHq
YdyF6DRbnS0GdIpIrw3g5axKpZaxMpG5bmpz6ihtzqsOA+OD3OIj48AkHIQiR03s
8lRrbjxjBkqIF8kSFfvzUnKx7MbEATfrKcLxgnt8EGccP9nxVDs87Q0/TY9jP7Ob
QBP460Ew4w2uxiHQVlbRrA==
`protect END_PROTECTED
