`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BaqTApNWSBlVE/Ec3QZy6W36niaGqqNVWyQjKWNzZKP/u58fcbHHgqz/po6BfvXC
kultUeuBAyw2fl9iVKBxGxBxop4R9rjIq7xAviCHH+ODAshfGqLHBdAh3OUOFwO1
5XEMGZhrRYajRR0NCX4Sa3rOY6W5F4iPel9e1F2+W7WUBl4Vh3mFOPlOViqFANHT
wUhXzNsNy4jjyfBYsudtz/upKfkE4JvmoLHOHDlQk0oYmyqhFM51k4dYtTqbbB+N
NMZiyqgLlui66apFzcv1bF9YddMrqYslktI1khwvuivTc9wfS8moGZx6BxR+30LQ
Rm1sTLSs4/Jd6wenk8FgQ3HHzBnC5ZAyKO+147bm2/wkxpLxlIId9JA4Wi8Jf03W
y1rmzJwHk9HhAgdodIcV6Nv8mXUodOJei7WE+mA0Ipiuqm5y714vn7RIV40wnX5I
xX2JHm6zkGBZ/cAICBMsdEZdr+QnSPW/Xjm3ZaHPGpm9S7RgqfqAwPf+ojzKGjxq
jxdA5JAOHr0Rj4jWfTkp37CUpEsj8xmzQ+vZbKaBgdFiSswxIiRNGFH8v2TV/t4E
e/RLu1vdViC/Ia49fhCZprAdybQIvZbLQzdxE88ja93qYpRcC/x7WL0M6fBhGyxE
Y0DhRC0rHEr210wH6OQI0mxkX4ruI8Jwua21ZQieY7cjZCUFEJ09bgcYYzOLQyG+
kuco2uxI/qKLz48cyr0z4dho+KHa3rV6IPQg+WN+cHL3rE70LDx50i3t0YTNXC50
O5iTwHTR0Xtd78NYy7Iz1hFrbOCVLZ2004idLMSbAg+TIY8KNZ+4xjFe4PDPnMuh
rzVHB2vuRLUt68S6wIGUWCcKyDyZsbs1G5k4A8ATKU1Mh/DiHMM4qHk5H1wu0UNo
LyRWhs+toEyl2nzF3C0lnsNmBd4nQFJbpPGrQtD1BPsnNHGGvdAa09sut9JVNDqx
bd0iLZDkOnqq/WaqbfLlhnNvOIUnznUvaPlqG2x8ZRdLAh1Ede17WRMWwJFddnVV
IKB9v3u8TSTIIJWnFMkDhfMejgh1lW2JGy8qXQkBq63UHleRzNi9jBNAw3eAJGP8
ctVO+KaP+c8sw0FhWVPn65x1JNbKul1HGOVgq1zdXLLFzCMaIi69YLrNAsXP2DXk
UfmmPY+OEL0oC29RcjiPr9F/H3VK/+GF6gAQolWg+csdaZi83pu5DDf7qvUOU/Ut
9ldOwjEhVQFimgLzPxVD6WnYrJvazaYc6/zlZbMw2czYe4O9OgXVnWtfktiTZv01
OwdACl8eCRNpb7baSBAptROdF14olQ8/sXJCzcAchE6G2SyuKLUlTw5WH63j+I1D
uDKUcqSLGvxFcVzkSKUmV+1sFI6kEKwsB1uTag7bI4ZQNocqIsUSMDXO1WkN1GSJ
T2i8ichjvLc/IU5AETdXtyJSRKYlYswuEG3tS/gLr11MvTLco1ktghBviQmwzrtZ
HdLF9coNBKj/ymmnhLlaWliKfuBDEfccmSSczdBU8X3rzuATtviAfF1we/FIqzJs
blCaY0U1Ed5LcCO8NDoJIlmbYqAKgSewQrY4f47X+shjk4M+i7wXXQT1OXO5kaX9
tVEtVQFognWKRXqJ2/spzCjb5Drghl2pkt/GZdaY7qe2i5ICs/3ttgz2OvsZ+nii
9QWVeFxX+SRjIdhaMMTt7MDsMBwoJcQauNphmkEgW8kZsvhBd6bT4G1DTk2am+tH
eGpbh1zrXUhldez6rATVDMQoAJjKhg8ZH8BzuOIZByM44rVhAzQLrPjgFFh8VDr/
j/dQMz7Ikex6KRu3SyDOb+3TjZ2ngWhiRTWwDatcNrLf/JsPlHt64LDmkwqHh04D
/fjrCaIyYYeKhanTvLKRPTHvnqlEYU2Z+8v8pTXIOzqG1j0AIQeh6h0J4mr9mHjq
fkHEfLOkoz85a77piFb1CHnnMrig2ssOLDmSQDt57vbISLVFKOcEM3gNZTu4m15c
UQvKZcjiVciC2Xx7Wy6WfMLgQzOUXqA6wtWj2e2cTouYhQ1dbQGgeFFGdAo+L9J7
4Z/SIDID8IXNyWYSV80+1nP9ZUd+dKRxDhERXUvSFKA8WXTYD3B/BAZdSTmXGvHY
WM7G+ntUczaKpTNqQOSwoOCsx1hTmPW6I4LVZPup1Yxwa+qVpgz75Rl+OFZcdQ10
rMQdPrFr1pziGJq+Ijsf+F23aVo5cCk3FTMlg43x8GuuHDatnOWiye3cHwr2MUa6
Xko6AVYVOa/zTwrNpBWeBVK5hD+H+tnQCOuF5eAt+Jq1empfoOtAsy5q8J/msFS8
RWVdvtVwQEbiu8sqATCKX5Ww23thuLmROqGPXjQIaP9BcvfXnSCMuJ5z7lQdfokk
MGV7OU7YuoZV56jOrAG1DXLs6lDH10vOB4JSnedtd0FRdHSQ1fLd7NSHDDJS4WRL
su4LD3K+iT9zj0Ujs3j7L/xDHlx4cujcmHYt9ExCRJ12soqGLw0XMIKnrmYy5oq6
8JyXvKRDoNJEidMv+js1iF7J0mh6P8vgRUMzyjZiOZo6OtgqQIKyt4zne8LayWCe
HsuCFW/4AQpftmjcuO5kTyrFMoNU6p0DTTYTfmcaCZj2NQQCS6ktIDnrBbXltx5u
xjRkx1iSzMenGP0Sqa/VC2WZnNbEVoaSEGv7ZsEnYfeAi9rrMFuoODNc0Q21LPaU
05ISDLoJqYGvxXXnDqMdpS0ho7UXdylYLHLRglh6jv1u3B1pJLZJ3ZbUw5CVk0Uo
7o0EEQGxdK80RqTmAo7n2CgJkd1zh1EzxyRHYM72UUmiokgYo8WsDDRrsqcLJIXh
aqv84ljssRA4c2vVysBrZLI9R414Hd+BaNIlaQ/Fxp6qdW8NeZVM1ei9c+66Cej/
6lKRxlOudvenwTG0tu/YHxGMlhmv+stXvNd2jCmlcWz6zWizPOcecWZXl75xPRe0
6X+MPKVdSkORzWUq+tsD89G2EcMJ09NnuZERMWat6I4+unEYJ4t4M7MobqnKe8Jj
2uJhDmTcZkJU83g7X22MEI16IkN2Z9EF8RpkLh83hZnJ0CPXi6nVoAn2GKWdQqZ1
9HWjYufnK+O3etg1hIqQt2rLvr6RgYEt7OQ4qspmMigQtYXdxguEj9F5fmmCqU4p
5ucsLWjzmxYnh0fLwujdsjvJJt7p+WewbUODhhxYSIqjLBWfEOfc2zED0UbvaXYd
J7GczwnoQN/YBbtP+yTfH/LpgNqwzVjHR5nDT/Q1lO9hD2lN+MatebVPc/DE6UTp
cCsAmjUo31f5kX3e779SV5oKRai6wNxq1+M5xlNifM22b9tr05UCLH6COg6gJ4gF
KG+6U31nMEZxjcSHJCzoUGCZETXFO9p3+po+s9INkdnE4cps//A/vJFYSAT7eIqq
oRhj2n7hR8zIHlkBkkq+EHsevnnMhmJa0CK5vC9SYctBP9DK2xJg0/jmqthc1a3k
+qb9RGdmsTNTNuPrUoOl8meVt1lM61IliH4DsiGQWNd+z27bF5wGer/g8aVd+WSW
8t7y5/urMePLjlqpa9mAvi5GSSpx57Sa+QBZMiNMBkXyxL7kaDLhRi5W9KxuaJX1
JfIOxrw76U2QumgGzMoWjuG3Tfc/rI6KpOdrkcPdIt1lvTmluSciEWRyZ8NbZqBO
SK9c5uEPGENltAMtKZGo7odXOzvuszyEN11NhqftCB871/1UzYbRvFF3hgtR6A/b
1TneMW4zbEghL1RG1x0eOcBa+jSgohgwmRm6v0VdUoa/g9UkJqeiXgwQr6VE6e1y
dR6hEQymZACzr8HgN4roAjamjVIwDJIqJlpg0m+A0FzMzAcVB814c2ud2z/7PpHu
1I3dgDq+6CC70/3QQt8zszeRv5/YND50jAZu6vvfEpiH+ePlU3VBGbQ5AzYiDJz9
c98kqK36tjg50dwha7hxhBmhpc7TvboQt5AEVUldhz4f+7kMupMDe3UkRKAmFb4i
qn0jPb6nDY67wdtX75v1x9qndov2qA9b9gvZ/kQ7Q+liA8BI8AcP3oOD13966N2d
JEiyQJP7iIzo/uMS2dFlxmIi36dMy6NUadbY3YgRSlDb+aVHRM+7VJT+qo7NPxIB
w1GckjuImO3tIT64UHX7Q0e/HnbuEgdIjpMkSGOZoXidFtYKX7IVwJ2ZIYJJcqgf
PiYHGqZaqWMltfFGd+jyMWNCDmkcSQYanTodDnIrPQ2iaIJftimYres078PU2VI3
JjzwA1ikMs2H3LaYtV8zpyBe2lRi+enhSPj3+hXoCKF/YQx91Wu8mvXn1NYaQY2J
5jV60485EsPjxiCI2WgsFBBjmXFHwjIrqR1Uox+ghE7JW3EB7ISjNOhsutrUDfN9
OqZVmvjoOyIslRR5j9YMMzqcSN70bEWt3hBkGDI1NjWiqXBm8a9eESsm8JZobhhp
uynqcog4Ju/OhntYscRl/s6LWa+pQSOHXsaWP96mfH5noXVQv86ZBMBs7cYu3QHd
OByWyAblDEX8Sp7cY8wUMsJo0DiZb5ER2CQj1pnOUV6+0slemhsEaLXfQPyz1umd
zp/4qsMlkLzWYQlqV5OhTRHqn8okVGMNCjDYIUh42yn/xLcS0VbJy3JCsFEJHTco
h84xvVlKUFA5Gyi6i8GN31eCH2OZlbqerCBhxpxiqprTrQ5lDqOPZS81/kpKaT6s
XmSkTqS6U4mcdXo48ISIaX5FDT/FqGF5yCDASBRV2rCuiJ7bkNia+VXrbS8yb53Q
HVRsMalavWVVSHuOecM08uVQgwKLjxeEEGPUiIj4UMw55/vmCZKPaGxFloX9urrF
t7OTp5Aigex9Zbmw/ZnQBnPdsqEsJk9wRiQVwy+g4HDYzEecKAsar3BANmp7ZjfS
zr3QUmBTrijkSh9Eb9xgF7QrT+a5YXzj1EHV8LYDrNFtud9gKLMxz/T1KiY27ACp
/WYnnX2NjvYrtEu+L2KuXHrupqhwswSqHavQR4bltPwNrtLrczMbTT6y3ts9tzoA
z9+NHgsol7js8s04OQcRD9K7QW753l7eyjxTI/mgbKX6gjbxr+nNYX+yb0F9Z707
lOOlQQdtCmLIKzU9+JJD/TZOJ+zZjkBsRjSC97NBh0aT4G3ESBPqz/eTMxOmxduV
IqwIWfPJO8/7nCFOPCRVWsqHNkdt0doJHmMcSyJdneTtowhqhtteiRBXy+UtUnZv
2QIB+HrYveFNWrujwEOM6MVARQlgf0s2/Wvq8CCy6mWK7OaSGdfpqFScWE/z0LO6
SajS/4jkHn1O1ksxq05wfsHgQF1PqwBocnIfjfaT6dxkavcBDhQ25RQpUOmdXWHI
INpjeAeb6CnjXNNv3lms7WrDyRW5Id3NOQyxaHDWEr7dDhSNneWcjJGoI47gMLxT
gi9XtVSR76Vh8oVEF85W1aPYVd4IIxnoIp0hiAPWr/Pyx2BfdLeDzaVdf8KX/QrM
ZILO+Db+MrgLDA5T8u733VBkoxZhGjxE5jH5gjGpJ1JYra040hBd0JxKkF6dISdF
siwwf5pH05S3lXqwy+9ML2V5NICQ2CCGEpXxqv2W3dfrR2hUskdeOrrSFE+Rw2Ym
ThVr5X+OWUaN6XrNRxT/RGwvLKmffegh9g48EKOP7PTAE3TdhPGTuJDQZqoSSEBJ
qxPQJUHxWNkhipqYkHRc6MWywC42UQcqW2bJCl6jW9sC8PhePSIskORT/BFjRu+j
lILMEayysMacaLMaAsC9Ffad+Q7vCXymkOs5BOe7D6aCGBtFo1MaMDa9O2Wpr6d+
jF4HScMRTgBDQwEtk+6mzjb9iKLJ5EeG6L2y0jisR9bbSOvkar2xvO+3AwtfhdK+
xsVKIQVCCWinZXabyjfmq4+pprp46gmyBi6AlaI6fl1mGPHVYrECjqKnEfBqG0gy
IVfsd7XgqydS3+SEnoHxFsrzy9k0y8fxqGcIAJZhsUpUb0prNSwZdoq09o4Z5HiD
NxqCErArLbsWSvBiARXXLkDamKZXZT1Z6M++g4XMKKKRFFi0qBP4z1svyIlwN7Mc
vMMxY8LQ1dghLKLAeN+mTd6xLoDsqfAd3aM+l5r1rLyK2Oh7QW/UVJ3GESGV052Q
sBKb+AFDVVSPauK9rXIyICj1cSHSLLBke3sUIlHWZMriIbgE0P0gONot895y+38p
L2NVhjtIGPBejp63WqugKH74TL2Fpa679Wmrq6Xfni0JevuOuaAIKJZApUUNXzmd
6sj4lpdSIz+mVZ4UezF5ENemmAvrPCN1+qk1ns5Hf6o3+jeddHdc1SNxmuYdf/Nc
GbkJaUI2+Z1jmim/VbjuNA==
`protect END_PROTECTED
