`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mr9gP6+Lz4ZHbE8q/O88OZmLOV14qnSlkFpThtaSSGLaMWCF2yzfJeuhl8mFNElS
MOVJKMGx9Uuhj6b3qRwA6PSjcDeF/Y1h/vd9XNta6qpBDY0HfP7VTD+oB/T0LZcu
PNv7WrxMemdD/sqYiwCxl5ugqgwJkD39Kr0x2Nrk6jjwXSoE23IcZkOUkzz/vHoF
KFn8R8AOrZWpUBH6WGRUcyQsEBsEWrMEWH0YZy+J5gS15nf7O8bXtcV2B0bqWhFF
z4cqkhLrfebhiy8nbmu7a0s7azzYPj0V6N7kfCJuxeXzugLipZLKLEnRzmYNYWcD
jAKVPOnP/RTAnfXf8/QrfZl3AVzVuH1ytHplcV9oy1MR1M7Kz2B0tYEjTBVBG9Vs
dcC15vbzFfrZk9IL3XKUPKYM0/1yqDRNThxm8IZQxTe9EInwj1ZhQ6lIo3Q7Td8y
O2ai6snGgZz4x2QEgji04W9WbblA0Jmvso2i2zGXIJK0bNLAoQq4a0KsSTtRSr8e
F6wrnCQXhSF3renxC2397qtR0ggtao2CIsVmNIa31sc9pPmz7IUIUfeOIp0M2dsO
P2Nxy2Y0VdzgJ+IYgqS9Cqv6mM56VFRKwYnnkEOfr8y/JXiyeUH3k8x/Me4PUmw5
`protect END_PROTECTED
