`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2sa0PL0WSE/AbqrxNQspFM6k0p88RShI1/rfS2LQhNoo+RTbv1AmIAG0VNXgIqi
ZyCKQpOw32PgKpm+OVDrgzKImzy+YL07v+ByNbGiSdWTbQ28LGDFrhEnKBVfTHTJ
IdAbvMLN265XvmlEKpnPBqeUnigEKxk2+4HfeZHTagPDc8T7lCofSAEyo/h9eG+y
smSDjCRwgi5fVZcBkTx4ZdDoB384zX5o/fSxr4LsNZMXAfzcxO45Fx5pvqsl2ju8
myKLuE20lDHXoQa+6Q4/aJVp/39gMewTKsqbCpjkGOhi7+9C9wcmQQAsBES81lUz
YEHtsfQsNCQLZnbsNESUcPwLtxTk6yGNa76EFsgMM66eNtfJ5bo5lSI0BvnJP+n6
q+glz+8/Sjh751gs84iO+HhjSQrOeMq3CXqklJKLlA4C0SRCBSw8LqyQ/xvxxIqU
WhXSUwv/3E/NwJu7CEalMseCaQnKoiksYdHVALIShodR1ftcMAJH7bxR1AQGm4c6
iRuBntMacle4IAFpjmouYb/GrmLiWlBnua9PGeQ8vkA=
`protect END_PROTECTED
