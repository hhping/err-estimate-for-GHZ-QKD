`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rsACFts/h8iSd4zJEmzPVwsXEXc4T4mNTyDobjz5EwIC1JmwBxQ4Ljnn6uJYUzV
pctgnGAXXzf8Qx2hO12WrgSz3uoITVPNaQr6rQovkRHzW+d4bEjS8vPqDgo/LqIx
zAfnYJsBzYYwfXixwf7cy6HVOF3Ez/+XlCKaBpm6vqOYb9ENDIEm137JEpjLdZp1
EaQ+q3Zm1z5v6pfzutflUFel4G8poVTNT31shlIe6pYOzrak5VHVHi4d/pw4UhGf
ZYqQD/+hqSg06yatt8m5Zgc/jyINQUMLf0/Do+ViacJjniXT55Gs5ZI66btsGhE6
y/s5E69rVALwCVvSUMfnqjgdBRrNo8APxmk9urNAgA8zgQAcK4olRbl27Rs8qAfS
ZYOJmSRXCyBtAnQgWjFwMGRAQaN0WDzVYCVONWx4gUW5jk85yAO+V43EOL0vaWZT
+c4l/ZSGWge52chs9uwPh6yOKGKEYVHZfDEOrlAFctHwwG0iMXsafKzV/fAwSchJ
ZGpg/5P2j5cymaV+T2H5QLN5ok0D+itic2f+NVNuNhlj11fC3MvYKg5RshBZgxda
jCuBI1zC2nP+SleOwIGqQDwwoUblVoU1/muFk3VTHeufKwZxH2ufKwXSuNa091QU
3CtFSRZe5CT9Qla/yRdma0eYfjiHY5invAmr0QXNhXwX4QyYeLXMyxBEbzOTnWCO
CZW7u8YlV3SLcO7EvP8xsfVGINwlewtt02GDhxPQj1dzXKg9X64dAsmsb04wnQji
2myYbksfRopsTV0jXMB5aGDfhSlsLCah9zvFQOP5k75cf+65a259AEkRhHVNE4l0
qWNd+3S4UjQDnSrwxDD6lw==
`protect END_PROTECTED
