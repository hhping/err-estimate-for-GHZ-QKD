`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUfKkcNnLWw3i5jdurXlCX3ivWq4tYY9fzhvfn/PBNLcaShdt+g5pBFE70EveNBQ
ZFIILtQdKiFa9eipsTZjhVUCZ/2a6SVTvNYyXspCktO+ZZUxloHmJY6VnppPMX1g
Cks/09zfwtxouiaNvxtfsECwN59c4t+JXEyKNMs5YRlyID7ejmUByYfE3DHCbsIm
G1e5/ERH1mbYxX72wW0gt6UkgL7Jj9Aa8WPSlMaENiXHKPZMGc6knNe1IRCIT7bh
j9LnUrhbuP/pJ2yPvPq6Y0Jy79AEVXV7RhhHpv51Klx6jMm7cNLjxuio/NMOl51s
4ye8MTZZ8GqjRfvxdNYppZaIw/TXeP2NVPFe2e/arg+4ED31vuPAcrcn7NonnrlN
uns7F9UPpk4gqRZqd+TvhV5D8H9Gda+bAQ330qErlFt4WhlD80eJ7/XZ8X138vH6
V7nasLecF6U+Zq+A4CWc/ndlBg3KktkD+YQr+emI6o31asopysEHLOiBx7mP/rx0
oo4/yUUpGjcGw0esfZjKyg4FUvm4r0HVY8LXPZublMqFE5oXiVNU4PJczWRt35hJ
DF31Hfic4WGCafFRh7cPzoXqiRl742Q1A2rhcKWk3BbnTJBciHG5UKgHbJQCREqj
O/gPMaNVVEn26MgqiH+YxwYtkV0bryy3JUDFglbvg4yBWIKnvKC25n7mbpWuQUKg
JRWwyv4CxLZC+Y1T0vlJZb0dDNqMlhoSn5iNKk538mgNtjMfOjtKG21NrWBHc0El
n48I4HurDOF0rjDp6mipNt/NE5R2/QueNHp3IE0BViaZ/HiYOqou2uI0FGTlkp06
vTIjMfoStLCgWBroedYb/cR4K+Afnt1BwwEZyc3hkXDFNGp44RyyO6ud8Fq7bW28
QHhq8/jAtJ9EhVlmClqkSxborYXsEwARewRh2tmJoS+r6G5xN1Ln2FFbx2SQJ42J
iXQZFKVIX7KlO0z7KLC6/ZufLPaH12ikRzGXuux5KcVUzFUCYxF7ZangFFO44mrn
`protect END_PROTECTED
