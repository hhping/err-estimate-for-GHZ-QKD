`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bubs8NopVaILcgAZ9LU8uQvwFB3lqVr83bhGovIHb9gLC0y8kw/Nx/tcpB1YT6Ov
sLAxVpH0exR+2W2ytHoDDb8lvGS7sJcJWKfxW5fmXNZAwZqmRbSlPrw1K9KBq4k7
GxsS3cnZa9TvpgBG4uz+o/QbmNb5z5vXHXw44v3JvC8Gf92EPeT0PDDn4l77BgVD
K5trNza5ZRIKuyMBjgMThuCNDpzqSrSp6QidubjaCLeKL3hlWHVdMaYbzDrZNYvL
w+crTIEcqmXqGrWzwU/mTYC1lYaEPM9bjhMm4I7Dts7bJj4/qnkq51wgtK9HuQGR
iYefZ5SWpQRaehe2OL6e0iwAvYt6diAKuApc0P6HgwZ+2lULlaql8XbQeqGG62pJ
9s30xMIBzb9kKSqPF0lQvtoA7DAnRLTMSzXw5p55FQbx7txSZAM6MLmlmt3s3NOc
Y7x5mYtEYhrYhUcI7a/Lkcy9YnLwq3MO49tAZM4eb4Q=
`protect END_PROTECTED
