`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mI34GHaC+HrzbQ1Jzuy3/DY/n2p+uH5aV23b936OM8XvgRQ/aqiQCd8kVvvAaYej
TXtQpHszYTLh1MOeFVU0wy7e9e75ovExqL/qch92QStaMPRKe1t4LJ1qJ320Dqon
5KPH7MR9fZ7jElQbwjA63sshmfwyRxwaBMmDr94+Uv1oMAbUUQnbyrc/3FDV1j9m
sXZPkhVhCVET3N1T3i7BIWfRY5e+O37lfFjs0QFtmPKjwM1L3y7GRzjeySSMZO3y
7xz9x+OX6GAdwAxuftnVT6SNHokjE15l9dVJPv/KHn36oJCGvnA9MqTH/EhCj+3g
CmHOcraB6CiHpM6ql+F+pbbnbWyoX1ACYTLXgoK09X4roSmDqaA6uknt9NMeFgo7
Gfdc9cebrAmRg1o7k5V33/WlNwalwGUc2Duz7nU2G04v9nHcfyrqFM8dJsOqaJ3x
2+tE06oUHYQ6dyL4V7/R/gxJ4c1fyDAKZDpnw2WmVVAye6/e1gV3mwPcPw5YfAcJ
8EChdusLiMkbw8obfJi352Q38nZyb1lNu1TEckVPpz7EeXfSAiXyuWqONqFr65x4
SV/U1K3thDmWybkeKcTxpH9uYLK0chto4eOabBtjid1PS8BJq3GuJYeVN27iOW1j
/z0xoLl+y3TaPurwVZ4uD/cVtAM8njNQgMhNblGUFVBZylsUKsb1ZOeT+uOmU8D2
aTpJ1NhuihIpyURV6bN9hdMe1wIisuuXYwbRQ+WS1Ha6tbHk01uK6iabMuLrsUWi
395yi8c5vDS12v6AvMCNxT0Cmsu1MhG7xzqRNzL+LJRrKhDXS+15d8x2tqK0moks
Rpb5aTWV2yquLKt9zpUJJqMlhhvKb7UWA+v422uhCofvmrKOTLID+YEGWD/22iom
06TviTboIKuv91CTxTPNY/IXPJhVeaSWRbxSdh4CR/ENb7O2wQIo3wQRXRH6Pgsc
914Gxq33vxoZW90iVNG5mpEuyzQDTwuHD4mRUL5JT+jkcLSyBKb+7yapMyb5xlvb
gnR5yHxVDJZ2eEkCWBlg+l0l6iQmkOHkR6iKjxkI+PrMqbuxPnk78bFDbYM2R9i+
8llr+ssH7+o3+zW258GERLdE3oC6ItEfpcRcg6sZG67DqrvJ4+VJWz7pjfLrU+fh
Vf6AKPyYKFsPm/CwTMCKQFwGmYCOdut51ZFtBqAXkNo7rTIFeWtzpOu9HHE1UxFl
WKL3wpVqvbtrfNC9jhAjrJAZO1MTLwoNUAckQKytMCPnuCUmnkRz4Wkp95RLqjfX
XWzw7gvqUXbb2rNCpv4KpMYRiB54eEDIg0CiSY5uBt5jGsE5HzU6LtaCXDuPWkje
ILG1WcG2UPB0uws/tGMp99Zsxc+k9mc02bhQm0pRsMkYu06FMgV8istCsqDWCW/d
n4mRDDMGs1pcnooKxrtD9ffY3ccYhJQd6+IE5JhHogYVnoev/2Sce4ghvCq1ha1p
MK8ixmBuS9SRln70VLOdRiHthzyLq+BaFbRTiHAADBr1jxddJL+xe85vUy4dD+nX
wgfDIC4w3KlM4lBM5zjx9qv4Xwj8xCSxM7jicShAY9CFY2HMOrYvPOY78xzjqGEg
daAStT/nlZMgSq2s5q0SmCHjdbB/Q/sTDC06ZLKct2eqPwILYVAWrxUEOQDmJ3Ut
1S1QuA7BCJippUy+B3ElNTUiDVHz+2doFKug++ty189DNi2rpaVkEHLuOta1oqRu
B/Hmt/bzDpaLp91s4CofPipDrBEPSHov5NkqKTf7mW8F+VSZfPFPdqKkE4yiJn/C
uD3u8E+d65jf6HFlhY9jUAIgIBYgYfXXqpdOWYDxF72kdHXGf6Jtd2usF85dZVzQ
nItgqqlob2E7cZI54YUVVsIQNq8HxILVZFMrUDNquqxdxTQc8E8RYVNoy2QDN861
H7YBjkf/QFt9cNsSPou2DZeycVaFxRZIsmhNLVNs7QQ=
`protect END_PROTECTED
