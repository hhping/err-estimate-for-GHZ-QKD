`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8ksfo3ZdigA+8ts70JOEne1OLuJuupLr/KPrOJ1Jj7DnUa4XpbTr8/SALXVymK6
wy3Hz7QURw6vZ785NB4NOitKY/eP5a94ptFvAEc+nSVQWAKJsmO6V/JNv8gQWpjs
Mzx00O3J/Kgc7V4Zdyx92bQuFfKfOQ73tFbnilvf/r8KULSPjQyMtanTJROr+sfE
VTpVC8Yyfz8WrtnrzXQm4N6cBOv1NxXr6hEEi6REfdx9NRlN1hhndWRnsmZjj5eU
Ueyii6tmaZmGKlIOUwrFhXy+B9NeUSkuSZ0ERIzQ4DdexGT55r3sMYzmzyPcqVoH
+uTvOxvw2w+lZsFuJQ16Pqls/T7h9JFV0c0R0jT3Lm7RJOFYO0+eAEYC6QUu8SzL
MHyveWkWXM9dMGiBsxDKr482eQNxfEZRehxQymtik+fApV34TFQgD6kGrzwxH94l
sbhXOywN2+nM4pmU4dHwJUOHUP8vHxAFoGFwvPO4BZV6POUhDe8moxKsZ7/k4+EL
e9T8UWu40bh2MB1kzcI2vHeDvgYgYVMt2PWTHRDbkXpOVrcwxaaS3lKR0dupX7u2
5MXHpBdtnOxfaJERczjWlqihII1HuQgEFcDxquHd8x75wGozgCDo4cfXgeRwsMW/
qTHl6ihBwYd+++jJRRefy8U87LQ4MIQrsPrEaVzc05zsmCcc9lATPXaSh0Dw7sbu
03jd2Mhc8Up4dK5QdbZo4s0jEaipz0lu7dSVpcAUFdCWezqJMEckt3LbCUEqltfi
U9b2RbhjAytHjcY4ZWSMNecfxVGN9Nte2wwPByWdcn2AjEnRFmxYXBeAKHhXz9wN
DsS+LPHNECF3v4AZ2Y708tqkhMNtlG2IWqfD15GtgadKvQG4xnVCkMYjHpfEwmgv
TTO6hJQFs2Fn69+zA/r6KilwCtm1+NTFElGGnUBcLSr52TQnC0VyiWwB7kxGZkLP
/ISIJPj8KPIrxufnqhZOUA==
`protect END_PROTECTED
