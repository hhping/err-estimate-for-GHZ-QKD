`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7S+F4Bc2PK1OcRmz3egkNyHe+J/8SNnh+IaojtPah/gcTllN7evOGplNprrKsqUr
cur39yB1DeMuMF2+9lu6rWJwkqtUPCIffsZGSAz+8uYbm4OlhT+g39Ynz/+J+cdg
NsE1y6MpH/b8R74TeL5wt/FeXtDz8H1fNON+LEzpVX866nivJ49k7sNiciOCmQ9R
YjVklCBf1u5OOO6uLTcmyQHkvEuX1STx3mRl6yPw7CNbRVgHJ0ggri4qEHhM8u2O
bcYZZpWqZ2tp2Wldn3xycNLrjqkowPO2juIxT1iFvyI/SFxgDh7h0VlzxdPZ55z7
2UlM+khMZeeCTf84dH6zeTGdwkst4BmnrjAysVXBVqE73q6jb+pmtfpzse3dvA4q
G17P4WiW7OAFUMkZsoaD+PMBwXRiCOef+NWdt7Bb3uGIvUsYcLNBOe2r0grT/lWu
vJl2NjNdDVJHp7bW5ZfP192LFTTJIBsQD+JEetPNu6m9AGI3QapdfdG3AJH8tKzT
KsGAeHy3UstJJzLQ9SWku2n8rbnpj0nDg/hTloTqLhK0+2ZL5dSlD4yIXF/E5wJs
v7gRuj6NKIHLv+q70WvNsHeiVqIvLo/gKAV+pKAD2H6k1YdwwNW/KP6jd1YLPYAt
S7N4AXl4i90Y+sCYgy/yvwlFxoQElqo/i1noXkkym32Ji1lYi7qwNwU+eP6iL9gl
nx9RaZFan7jBWfMcQMz3AKBYGE1+lu+WWG9AyRjMLpNwrVmJi0fvO77flxSp0d5A
`protect END_PROTECTED
