`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AfBH66oSqSxSsq/HP6622wnWNmhhhtUqYAKNQKsT07VhfKei/VJktdVnYLDdgdsh
4MvzZJJ4xLFWzwwTf3OvCb1vgAmpYcs06qDh8K106rIZjud6kweE+k9gPi+8j0Kr
hTpHVT08K2+q5ljLLzwbWqASweMuXQKeD8ZDigTb9bqJObkycuCU4W9gqFqLVts5
ct/+S+yDgX11DWzcxBF8zIdsJifAJ411PWXks/SGKtOy83UnQTjG81YkOfTl/Jc2
DoBPJXwtmWGQJjvefJdYLtWGdtDtJcUvESjwg6/YqtIyPmciwHKzftbr5o4TS/HG
cjOYNxZL0Lh/xs/ZoH6bKFHZ9sojDKee81sMoSvSha/hJJHXSeYpQ20Ahjl7I0Ye
NCXenWvY5GhE8LHzVJIk4OtBu1JdD/MGs9LOyqpzpvPi9RWyMoaN4KRL1lC/Xnug
Ia3m0VFdSv4AJ4q6SZfE/5dymN/X5FAVlys3LfLmV5IYey/tinh3R2mCkuDFoEn/
NNwoQz7THYskVYHxM4IIaws7nBMnZbB7wT7pyF7dAgbUcGlKUD3z3sioVGdWhbZA
qCwXEpB/3Ml+OAgz7WSsxcSSOULlpLC2FWt7lyieuDq0230WAYsyVZaQgFH8MW9u
81u/DL7EfrYoEDAOlrgad7o76KRlXDf5lggjE5J19Uy2FaO6hxHcuZ2PBnqtbxTs
aFd49RDiKfg4Lq3sYc73i1csSmjq5GgARsyRinbqZHrI0WVwvTQPxIgIGWxTV8nW
KxdmxWvb/nA68UVBuRwn17U/eAizDOGux7ZkfhF/StlR3h8iK2yBrsyS+klNmKHb
TBQgi5FLZTEQg/EFLJpbQDqe1sJH2ySS4Qqxc4cB6aKUfWIzL644RCLvVwPLDVO1
NOmCfUOfGyzo1cbOcGx0dUNNQQPPZY0OtPPmngMftp+5rVenpDGQ2uhRzC3Wkpr4
Q8NTZ+u42aHAD1qM4F5S3zuU4f6BY+RuVGAIIIIK77Cp+TGHatEAhRpPpjDPmjOy
+nmJmH/DfRijO2sLlU3VKCsU0W6mAUi5OMadgdi5P8HGH2/uBhaxw7Z+gwl2PML8
Tbq/qEhVXcbSYkIAwZ0c1b5hHxcXAQUcIdN4irK9kun7M+GpgK72PkyV1DuToBB1
zh9oUdexFSn7L+LtmBcdD8slpdIROeeUCbkxcXmMbTd2NUy/wp1MyqY3ntg61YA8
crVGb5RIsh3Xp0VbHZHC0aD2uMNmEPFLK6IDp/RsXHVoTQ3FLIxUWuUpjWGuEWxa
1i352og18K4NcOn8xyrNc0aVIOHqfbVWampcRJIMcKfBllQQAxxzng94xgKxAOlw
U65g9K6NC5SfRKf/JRB37IT14FGBfs82ch1PTn9Q4dDumsFbXBNZJgZLb5fPnJxJ
Sf+AfGLpvhNe99w+ErdCTtjf9IM1tTGAnSTiVVoEa82KOQPlJ5FZAYqh8ob/UqlQ
YSAL/q0g9E5pUVoaXLqcFuvZitcI1vKMhPLJDaX612qKbe20ApufIyTp/1ATBiLF
HexRZDcFNkIndbV3KxbodUNU2X1ePBnpFfLXUJuSWk8FBrmmmDNsJ2uWTNJ7hgQF
Zt0BkydPbnNYwddWgcwv5A==
`protect END_PROTECTED
