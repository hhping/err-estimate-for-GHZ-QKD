`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0WATD252wWU8U3LCq9SMbvf5askDaOw/Chdqnpjw+2Vpwtc8xYPIFrVX0g1kYGa
701GkjGvjIVjAAukzOvkei6A86vjSpu5QjWU2sawfSjmYzRn3JJU2XhW+qaWB6DD
/RlZ7uQLZNGRffRV4pV9H5w50Bm9IixAQCwlJpxrmRPjdXB+pg7ySN6OPJDfsZQ6
LEpj8Q++yDYDdOnW9ZI4DHZh5t8umdblWNwSii9maJgaIz6PvtFv3yX/jiblW8vh
IryNaMAP9IYx2qCE5lk4DzZt+BY13JGrZK5lSAbEuWbid+dzo9WAnuUAB1lO8kBK
zEAbQDWopUWbn6YqUp3tMvg862w+XDKHHuaIgEWchAhI32ADnwy7AJ5jfv8VuqJy
MNRKBBPtPg2/X+XW65yjZds1SYlcQYa+C8YLywuexyksEsNKGYS6XKqnZ233QrMZ
`protect END_PROTECTED
