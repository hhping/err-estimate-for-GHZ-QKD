`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0qXiyogBoluGVa2jgkbJGJSerteyfkxpGHnGuP/eAUsDeHxwqFzv4l6OkV9ZBhQ
+T44FvLp7oEvLkpFYN2weIYpokhR+bbWH88HhnZ42CRjowC4RsPVktqkoTEuQmAq
ckN6qB06l+N9bVIg4z74M2pf07UNAkI/IAeRsX2445OWgdcuCIc2baGBXoWlLWi2
42dvR4E1vLhTqWydYk5OHRizvOIQzfJmd0EXcDT+PxeIliM//yjxVj0Q6pqpTQEk
WN1mOq6OpegcjKQw46xEB3xkP0x9OJ6NfjWNl2lBDE4h4qCRTigNa0cjKQZFhFTQ
nBxdHchub+HRtmQNgn0yDbgeKfFK7b6aZ3UX8HeWahnEv3olHGzYU0t3yKa5dnOt
t6lGaRpEkhd7FLLQVUfuH21hGLGGX6bMmyXd7EVcCZJuN+x8ARjEPvAJXpUmtxQW
X9JsB6d7+EX4kpXMT+IqTdDD1HJmEOAWizzUQ1NJ6I15GegNZPmjnSx+xYHwMHWj
x2BX9a0d5X1KB9fw1ZeVNTuFjn8OoPriG8ywhCn5WGkXQPQk88XrOGd/QpI1aB39
H/yd7PJU5JCSSK1x5cK1+M94/2d2dtZ0M+Y/0WHiWKwcKPOuRQgVsSN3tyUYrtSK
qWF6QoaEMXNb3QGvn+LFm7Uxh92a41Mamozjp+WK7q9deIOFabXpadJWPJuCr3Sr
oDgChIFCYZjpLL+jp5vdYxO5OB1OlJEMGw255gbhWAric8NB345TRkjLi54BShhF
+ZZfTBl+q9MX/jCVgdUyHTMortSWdIXDYeXT5OsGmF5wIDYIh8h50WiDD/edyfu8
/F+MrJus6+6xbntXEymomoXBTGvdQSV1+qkN0CG2crcXZvlnGT2HaqMXQQa25jeb
Z7WeQQEcKwaCzKXv+B8AyD+VcmQt4g+Pa3Cs0tBOf8FAMpXuM1MUymumtuCNRbWc
l2UurSPO/9r2PszMqOTSfPJjq5dfRQW3P65KxxkjMkye1rC6w23UjB9c3kR1qZ0w
i+gw8hRBA290knEiZvXpjSL3Kgk80qustMa8dEmB3drDYxJqk7nwbgDJvJThK5oH
8cPNTI7SlpPIWtaTIo+yu9Oc0DKffDbo9CUJJfLsbjAY2X5KdKzOG6ub3EweZ5RE
YHAQnACCnkVDihA/qWT11HHlAZSoE8Ycu0Cd5rvMvuOgltYZ7iOpa7646LfzFg77
Sj6ysoSnniFuzojO1Z3DoDpgZHnaOi+gzmHMyr7Bf2BDpma8GednETr8LVXSyoqV
mLSg9rgsvrGZXzXIkM/77SI2tmZD7enE6jsNwSo3+nk=
`protect END_PROTECTED
