`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csI60DACleW9ZFkvoLtUwACNjZfKSRPcE6qfx7NXiMCWxfWfnaHdHastEj9JWCZO
kCjx29cqmT4WHmWSudQI7MLvm3yfV08x48hRYZYtsG+Pi4MUzrA2oYX8VZq4M6cE
wCoeL2dv2Cpiz75jC1nR9kY9vRbeL4MFLpDHRKt2azrfP+6Jyg23iuaUEQLddi05
vuw1jUM71qbmLHRR+Joc11ScUqjrOXuZvj1iRyi0IdMswtAgZlhU9Dof0+g/WVUq
+NEb8E7D7R7SfN75MMY80rIeKxHAOoUI5NrpyVCRdLMam9wOy/wzX8awZ6319RBa
pepuB4R40E6HleLZlY823EWIon+X1f+epF7pKe08nVvwz0jqEW+aEBU6qcsQqwuc
8CLLTgxDUNeyg9VcO2mjxOKoKV2CWSd8F8sq4T1yjytetqOHHpf7FiQ1c1IlPOdH
8WPE855QkrmAoO7Fnih4A4QpkGb1EvBfT67Zb+sF85Qgm15+Q5eo1feXmRhfk2xW
4otqqGoUob82aQvH7ibVzc71f1bWroF09aKAd3tb0LjQiUg0hx+XGKLfhGS2j2oU
+iZOVNZKNaLuI9WwOhBrCpCjmckky8VJWtsuQjbv+WToCY3iMeoy8adsZKmWpfCW
SKRS5X1TSjxru2BGIuVo7jgvZrTXGqh4iaV/3gDKXwdylbPpzatCOmetW8rLQ/L/
L8GIR2sASgJJEcKS9hndmB95yu8gP9GPdgmulluZzmNzJAweYs9OGdN1atQEj14j
92RlCgDbRiSxV0d20XHKwLvTrL2UVbJEFa5XznEedHcPYSDGoGJV2nIjSKu/d8pg
r0XjXYUoDmM9hZpyzBrl3AL/h8Wmobr6kJ7ePK6rtKloGO3w25RPq3YKHv2MKPk6
do3ib+zOGRlvF3FVf+JKwpXIa/nSOqLJzasj4ETnvAnienHIFLJs/+BfbNGm0WUF
owjAZGqa5x5DnIFanW8QHNrLmU6rdkvGLDEtbnKtaP6T6QrtT1tVyG3v98oRV4fj
HvXTFXSzwsyElB1hBqUacAgGhX6fP+fSrz9i2iKbTbQE4cdYc4QY8M/g1VmEb4O8
ZCm5n4zG2JU7KurEIYoUJBhu+eh4Io4EBzvcL3aRS5wqpv6sfK30BoGYtuch6dpM
ypT2b91SIt5fgiMPeiZ+Z8DEEl3UnPrUsuLBBdO9VXon1/8F0ARwoYgSSNMs69oY
YAP6VRP6Zo3qeCSdLia9d0yxfa8ji3NDytKLHcrued9oBZ/ZzsMCJELFWSmP7Tnn
Y1jJdAK+s27e9/uwNCvUfkMoQYEMEiD3j+G9VMOwOIPIZKi0oygcs9NXV7vNWsiV
GZI9usq8eM+4Ryf9JxaZNlxduaOKmbst360MJYUCrrqYR3R3byE6Hq3W07+4nCKF
UpfGXVvpDPGgrWx6Jht5yUe0Xd5mDpu9UaTkEsqGztE=
`protect END_PROTECTED
