`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoCJh6M0Tjui9uRfyGq03meKRaYKoCyPRMlK4iC2Ulu8564uymr7YCKTl1DjHT4X
O5vucroEscdgFRyq5yGmbEYqqSl7oLtfoIL3oYx42JUj9BiEbLpfu7rIaeUdMMpt
ER3Ias9O0XxZwIvMazvY0mU1VldkF792WNjPAdqUilacK55oyl9dxfl8cWEvgvLh
/2WFkkwn6XcBFtjJAxzoKJgqzXG7V7l2KpWtnfgeLRelBZtJSVjp4Cz+Qg36jQr8
M7Xdf//PzmHCDawU3oNsSTcEBsLsmh5YPyAhE4YX0CoJ+wyCXRtw61GDKNpEc0/4
Za2fjXaywKEt8IJSJHHOQpnYLoQV+MCJqN92FE8cNLryxC3gsmiGA8mNQBMrwhuQ
`protect END_PROTECTED
