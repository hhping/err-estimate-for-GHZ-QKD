`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tyr3Sd5A26zi4zBz8ohz6Rnf7jPSIuh52y4eDtpIGxQ7V7Mo/R3eMMu+sl6qWJOb
DGqDIQkDdyAhGwsoM4hzRsG5Pd+Y1ziRcWNclXDsbHI1KryMDZJJp1soPG9BVHMN
KhiwiL68fD/NiajESAifzXu062TrkJPF2TyW5e5K3oK4olKCfYvvTnRiSTRRIXcN
5GOGqYYSbcy+vBfDPlCMLwOKjPWgVeLEKiJwPUsFrJpc/pg0N0Ef9Ahsa8iD/SWr
r1X5fpkqyMc7D0+MHYwnB5BE8dW23hcDKD6zBlHCr/C5/dLhwA48e+CGP9BlRqPi
lAnVx2gJ9xPqW3ovkXJLH5NOZzdh5qtaknz/GVJJlkq/EblaMz53/mBxGHZ9NtZz
hEqRVkfecpFfHazWD9CpvwDymoVDjA6ZIbBxj1e8GTvBaBGoAI/w22V4+IiY3z6O
bcoH9z7q/4V0me1Dp/zYoh9QwtSG3P7hr5E7vWI/l+VWVGbhHHvOPIeBM2fQylnH
zp3XQwTivJyRuyVPJgqTggiDvCZSHdon8QtIZYZQbcREDp6SZDNE0wHs8E3IIzYf
zYCScIX99jaCG/dTAZ8whQQ8LYf1Kp3n2jxfWD0DI25nd5Hr0HHQLrtqMaxeGUV2
dWi0Io5L0nHKMHLJLToGV8XtHf4HYIhvDDXdj/Wu1NmY3siHuWCM94HEzVia6Koh
k5G90gtRIUQ7bjosd06Gsl1GO8rC4byMfr9vvNCbPDGJaICEnrPEr6rPfNpJfyYv
baD5xUdHVv6aavpzuev2TwT9DJ4DfOn227SO6TQz7FS7ArQD2ZT9r5EdoSsjjjvc
IwlowEgXd07b4XXhLTKCdnlsj7DUjMntZL/hfoqU0oylQhXAJKTGYmoGD4FcGNF1
c/yidsYOCm2XvEGL7ioAKGJh8DqyoVkVxP6AkYiAMCWArR5HXsH0fGnrtWAOrZp2
ZKGK2tTm7tL7lIIQ/G1myyiI/b5rnTNVuwRmdDiCNDnTZZYk0A3nSoY1dMJ+xCcp
tONt1BcD0fuh7mPaVLvTeSKKkX1ZA+IQGsbHEgAWpBCcvUXg08n4Ulbh3I/a2s/5
xYxzj+vI64nUOdOHNt9mh+/c+Ere4kKBoiBSoAWZW+M9uLh0EwOI09c1zU4M9wX3
6TJB745P5pb19FrtTnbnQiXFikg6XUDgAUOpY7pm9jYi86ueUJjoXp4ZSMminmhn
bGN0BwKQS+O+o94+gOL9H8JwPIEiFHwIAF8H3/uqYkNjvoyNJ5at467i5GfChOES
N2SDZa8BhBu4pR+86WHigUey927a87zMprl6necGLmUBX5NOAlDqDufPQtLWIwHQ
P0sUdHRDLNpmPZoOOj93mZMYDZrDE8N63GYOllmMLJezb9dLX6kT6Vi3gwsBeVZy
vytSGOy3czxbwnxHeXOY6q4/Rn0gYIo+RKzA+pro/nnOtL/FpwcvE9ExVT5SAgv4
0QGG8GKG4cIihUOc548RrWkysKAIFqPYfHyoeLbK418=
`protect END_PROTECTED
