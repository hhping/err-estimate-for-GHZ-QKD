`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h6OUuYCGlP7Iz3UUtgvJFRTO9NiKqRzRYwqbUrJpju6eFiLU0I6k1W46UBlnx7+G
4K17ZcBIVhEp/8KIpEm8wDczB9sqV7QVrFaVJl4JFKqER0/GZp8fHGfoZeGF/6dN
UChLl4/rg5vhyBO8RqdJQrQqmS9Qs0IBnENp5vMVVMp1pLiTV49BLWiytKiD21SL
pL0F5INfCRVWqD9kMNpP6NZLyO/Sa1scEvhpgVPreVtw9J6u+4dgoqGanuu2jxtr
sGcPxgyZg/iRMF1sWBIq3q6QKecFgUaBZ0bzXWPVFe6+0ZZwK+ML74LN8A3LlLhN
0KYPshvkbczAYnYBd0yx1yot2FjMy9afvHaZe/KyVutB+1fI7eR4f3dmpejHOufO
M4PVgbnOppNs8H43HVEqt2gUmnl+xBfXRpG1HviEcGL7wi9N4q/CMogeOgN+vRfM
hVj5LJh29JHQeCX29Q5bdjRN6bnri8gwaK1WbRLVGWy+2tipOp4dlcBAib3/eyuH
pZHVa0R1bx5mWLnm7TmuRB+tMTgA4RubnBFuCk123zN9EOL3mzz5vsk0LwQVyXr2
JvuiFjApT5XLZIRfcdmTeBWRcyhwmHYE2KMgN8JNadCgSaQQhMFD4UKFlXahffgq
9f2LFpAuMYky9XtG7OgNfUFtDEvf095D/3BHX3bL/2KVqY9P09U/+djx3MqY5f2Q
cZ8nzbSZhjjPvpMAPNjCzFaXZf/XXvGp/a+jE511mo0O1sWNXAsy7Ev6cg2iwcgR
EH0Woha79ERnBESXY99bFt82GFVl/12GP2KG2vJEHlEqWFzyLDn6MpAJpLQ/gYmI
DjvbcF7MYYjQxK58fDeGXIN3czSWD0rg01DAFvufbSrOiODu/GUPsNBtrQt139YD
bxwAAtZnnwdNjKg8cX4NdMVdoXyCwWB5lNBtcfzTVDRxcl4qiRtdBvpyrQEe6C0k
3YTQUcCim2dPLcAzx7O/NmEec6DtM7ofji76ueG/UrxCN3NovRs2sG0wsFyM9+j+
ZpR2TohPRX550p70WPFM6pto15QMZwnJoajr2llbrijlZMxcawix6WFlIyiVXkfS
U/7sRIG0o3JhGNgqFmwKcJww0DJBa02qSVralAWZcNCLFZh1cB6vQ6DPVHAQ8p0t
+LUHM0m3PNAN9XiZGDf9NoAShG9ethXFQ4QdcsBtCntVaCX1LjIBIfLcwi71fjYO
gqzFq+OR7meVP0/bQHX+oYJurAomte3L8JMeuZI+D8HxgRV3tAhHdAOWPxCxZBh7
j9N2pHFg+kAHPwwjXlDnbeU+5kbVh7vqLxRY9yeJsLcKrZ7/gMDSg2hFlSD+mPjy
nhRIujCYzrnt+OMEOKbyC9/Dgyb30/YDuevx0pW81TPKRBzCM2yPLzBrWNNVZS37
+dKxdxyTgwJfA5QK703Sz/0R8qK0eKU2ViORg/W8/HFdMvKj1nSMr4NqfHBHWBDD
U6J0udSZMX0/xraRlInhkhnpMWALBY/mFdoE9xM6qSiICF/8rq65kCmR1sJ+PFu/
oOZM/dgdfJuc1FF/mN4vRBcr9sBLuVkhiOmyyqdm6/Ls/J9iu9yLGOg7BHHg/V/G
b15Xmw51B7VwjAKKwzuVti3fKTtFgoeeM/ql5jaSIoJABK9pJPPQHnfIKZ6CoAw9
IywwkfHYbcjvwhOT+aOVJ48Rirga9m+FRoz/taYRDDI9ljvRjx4tS3AzDsoWrnYD
Dc99qikRG06cartyaTN0OuWflE+KST/WWy756UB/fMZhLctjHFA9H6EvHgswtmlj
4nu4quzpsX6w7jiHN4gE3pcfgYNEwCUJbxZaSl0WCCwIbZOoUzUyg5eyVlP4ydYB
9WTQNSR9gufIjuM5kZmuxJE96Zr9lo10IHGjjITVjahXv+7KWn03m/ju2YddE8Lb
QAIT2C6jUYb4tTe9T9pzJh9af3e5FPqFJ3FPACzj2u9JbU7FZByZQds232WILGWT
h25mEZgX5MvupKLYCHvD9LBPprtVjp16fyPBFKCvbIAAIbt0lgrIz2VxSX8qx2pT
+gWKJJYv7LJ5aQbW7Nsg/VScJge3Re/6uDkGc/Tkzu+M2sjcfOPPO/yQ2ujxZm7o
XrYhpiLu4ylFL08vPFoG3NpU/H1W55y+FCGnubiOaQKlSdjy+FCULjKribqMcIlm
N0CgEZhrGV/8gnJzQYxbOsjDlDds6udOTtKrLuDuhL/IgsvNhDQyCkDL7mlAWwEg
sUs+q7/2KWZydaQmqsJ93u5Ml7GulnVqwPT+k9rYE4YAEqSmjW1n2/JB0XjC4qg0
LQoI6pos3Z9fW9UReU4tG0PE0Hf6Kns3dQjWMGupcsbzjYeWx7sEJpwnNAnZXe/U
jbh8YZdC8oEk4gY7Ii2eBNDDJ8pKERPTmH/jB5ziwPYBDphA1Xf0t1u3Dqe7bQPk
gkzNVXusnVPGBXold3TvSj1uwmFPyuCImhai7gCREzG40TfDY+CtDuMbdNzBVGMl
Ex22ENvfysCJOj+Btnlw7rSTiSjxS5ziw10qKKLojCe4mBIj5+ZjMY4aBnnQkqQ7
630EDoq5n1DwVaJk4Kyrwg+L9blWosXj7uUOdPAkywfoHUTg5jO3Ie/BGxHgB3Us
RAydn8LJVrhodfNtcIdTRy8e7xQXynyQBrLG7kiRR5FPoo4t1szkg25fMsahb1if
q0bHgbPP6uj37jzs7pNACFT2kdt2pSLqpleZqW+Q6ILBa6mg8pqkgh85fKAf0m/Z
1uDI/WYRkGhdo0hHNugRD3/AtxzqE1I4jrDd5wyi997VmasanT3EI0tkcrvJtfFb
HbJXNsqk9kWC+o7ggDJoZRjhanJgl3yO/wRoR6u8JPvFZKhEsYnBIPjAzVHDn1Bq
MmcGCF907Y2Yi1XSoF0dk4+yK+lRCF6iZ5PveNbqYAsnnTZ23jBI6jt1RgVQsg22
5SVggNwmUGMF2zM0yoCycH/zQ+3tolzCCSoyRbG2/WOfRxQ9MaedvpRl2+4fWU+C
msGfUAsix+9hcN+cpwKfucRHAw2mQ2aVIYZQcAnv4cdzF+0vWiUOot2u0TUH0iXL
WsBQIi6Ri4G248lhlFAR0w3U7RQVKraZ3H+wmxlriq0X8nm5hj5WIv4kOl2J+aOQ
rF0YP2kgyGQQN7dIwY4tnL4tQhOuYH7NiK+VGlL9kr8WgG0NQ2QLbMk6D6GcSJTw
01DVxcoXKgcgzKfRPLAs4v/nJ/2LrGJhAIMSp+LKOW7qlIxVfsiGIAAi7RuEHcDd
Ycy6te/MpEMZC/5FD0ZdZP+tmzFFsdP4cUPO4rviKRF0LJvExMy3GhKcJed6ensn
EZF58xOoWnpeFSTS8qRwyOv1HAlU/9nWjwkPril8w/WQ6zoYt+tUE8IwhYnwySHs
HmVyN5ONUKA65mPs58RwRZ3ygGo/+KMWHIo6jhcldEq6X+I5OEIAXR5ZGZGUm9y5
4LPgR2AkID91HNOFF3Oyjz+J5PZR8BwYBRjyS7dAik9HQI2W9H3+6RwQ+pmtOtDs
YYRoZPCNdXDKRte7H7lSLniVtLtJOKZkvO7S+JDwFzfdomz8TXkXesayi4ehgXF8
GGZkHmoZsla7AbmfShgFiQ0M8GM7AWJdk5uyaemcUVzFcpV52+Njm9Rm4dQcS5Nn
OZ+N3LzYFmme8qutTZiEEQUnJs4b82ViTymHcoceoWA6BOuhD+b10ECm/OQ1VDfW
54h7ruMyJZ/ZM25MqNQey433I/hQCQX3kd8e5/ODoHZE6V0bTjwwPqD9R+Pl1WEO
fuE07grhC/crzNCFTvilWIzI2pdhYAIyVUzB/F0S6ofz7WZdGeK/L2CWbbXUxhVn
ajk1mNSVfoTDpbGlKV8Ybg5izvEyGuh+RBNlEicR5wXy+fLBZ66BYpwo9oU4QPx5
/xdR93ccBzZXZfh3z8UJ98uAXfgKAMu7R5pcHiZdKHr2sn48AhYSxlgNUVpYa0XH
Biqeeo/NbGd+v89uCHR2gvNo9QLi0PbO/FSlC4bOfWKek0wEPyW92Z9/spOmVdkt
LnPiteofBqmHacihG72ivMZAan76oPgDtX/s57VLKBnfmbGNiW43PoBMhudm+pRn
feRtunnkPN1i3dVPRSdXzV/nRxseG3Qc5LoN5KWPhTqJXpXJoh8uA0j9AP6tpzIt
7NNodjvCgZduGGXWGFEM6khrYvB1gVqz0r7ORQwGeZaE/LkHBgzK0YZl0ExYdw5G
WgJ/WG5wse9f/Cb453sqXIDc6MrJl5fn9lk59cmpIxxISlQxe8byqlP6JqP+KV/C
W/GdU2SrNIuvfujkWDFv16ci2p1zE2m5N4R6GLfTDOBLcpDjKcDKLpKpszBRVOy/
C7vbrjMiVjNmUlsT7uUIvN42RU7aPujk5r1/etc4KZ0uA8h1gpPcSJIFFEgurRnr
8NROoMxrzsjo8iot6TNA4dUo1LxSmDLtEndKdFPg/u8cJem7GvoG2C4htPkuKil+
drTojWwWCC2hokITXIacO2CaRgCqf8Z++Jc7xPYLPwG8+R0iCd912ePdXKIACg9A
/1bjSiWcees7HafmuOZA7VIt2SBTi/lghScox22aAtMoVT7fiA6lBbi2kRR7sbYI
U5SvkiWp+J8XGNO0QUAMc1xhoVh856/JMtGJF1aJQh9LX33yggvWRWcWidwiqNa1
lzTnZRmCSRBtv5BugZv8mY0Xpbzb0pcgKVNOnKyT3HoD8qt+zp38jqGrIC1GPf/K
Zs/uspEszqzqdbA8NTQLqLSbImvsq9yWShS6+Q5jMLpcUE0xiIMxwY2sXIkYg38V
+fiOFbXaqfmbdloDnhiHKTxHLwlsyh/5Wa2Vj0NCBlkdl6SPMh+7wS1AE/Cq4vd3
fWt8hGfvFRbsFufWC+EuXQV4dQtHRsaKYz5KopoUFD+HSDW36lxgfWiQSxLLPyjh
VNa7YE+eSSaKqWxOWDfLVgoX+mZcg4UGQrJbKD90uNYn0N4jLvgG5XoKoiR1Yg22
2vKyNFvY+8JvWzwKgl5BPcAJCtmMZTv0BUAVa0wxCq7jh+l7uhQSvtHiGDDIuR9u
ggHlGN+gdQ1wcF+zZbqL/ZplEqMN9G8po/DxvuFcGzJMoXo4WTuK8MFeJ4E42mNn
IkhGzCcwtVLfvIy9X+vgwVU7YQVAhnbLeIeg46DMYNzBvlmiyvCJq5mg6YzkL4X/
4DflsyyyGMRgGXqfD97NeE7H1lLRD6yf45fhbdqTXJIWNCs1W2D8M3zBZ4W61DtM
vKRo7Qzd4nkVf51CkH4PpbS3BjqpHBHITl/JJwZhqSkTBL2WyKRjqQ9XPUuZ2zHT
JPzm3Fn4SCatpo4xmlzuSqqrNyZBPahhTNMOW9xATvyVrgPesH49Ne+soxRZCzrS
05OtZlWd4pI/gRJemmtW03kAyc6yIBFqPqw5ooHerva80xTJUlEeSl/qQ8aPrxYk
QUB95SX9oN6xbaH/VwTndo+AE2D+BJ0lhxAG2uZdXjGJedYotVdL70zalYs4ThvE
oM2hmuD7h/XlTb/x5HB/qneE9WiYI5WF2g6eYpFW5NjkgVuRppCKmSf2uvN1ZJVb
zW9xuyd+AS+1gkMZ9d/rldUnYHRRBks5t+NpyRXAb+ThcKlSsfBt8c7Pi01EFJfC
rZPZB9UdpB7+U+6a334ArU5DZAv2Ra8XD2dw0FiRGhS8FP9ULYtWZ5rOjmSd/eYh
6ZX3YasHip7WNoTGB55Nz2vxZPPwSvFq2qF9ILOe7gV+A2e8y/Y33dj6Er6Ib0E3
H8dyQWEnIomQu/3SEG3v5tImmtrApJ2q+XOa7/UbLamM+PYWITsZ6YL+HTt/Ktl1
faaeQEI8Mm9uGb637CXl+qgfZWtn6jyYhmtKG/GMKOyOfRDKR9hl5sD7r7F49n4H
3Ax8G1aOATsF6kW40dXWI/kBRcVDa/Hdu8QRQ3i+Usv7Ja3sPmYYxx6qaK1umIT7
Hh111v5lakvuE75IIygc9gjqImWTy+C82y0O3wKz+lg215KxFOpd/3GAS2CI345D
uzG04LW0XH83aj5bblyDUq5cvdBmk3PY4EN5y+0CjdZTjtKuJ1miQR6FXXcLizgE
hg3/KByZ/XKTsJNFShRjNg2TONaspfUjUT8QmUM32w4iW9ldX5KYzwJccQDQItIo
kWp73UaQlCMR7L+t2Qzx54Ba6kwlNgnS01Foho2mevMvcQUyy69r1ERml4baZVrg
2DKt5w3Y8EAqeOyOrsmpWwA9ZNhUBbOY8h0mEU2Z3uFjsreiOoxgTK4mCoh5CR5M
xEDdWS5IuNoJnGsXFYT1O3An5BcUwNthWccH6lk/dmGEIfI08cWsCE1ShZhgyuCN
7TOq8Tz15rAAjmpjxLigv9Du45TG+nY7rG3pjuXoolLWqZ0VA6zJ1IWjTIs9RPcx
56eSw/LkfAZYtIs1cM+ngMSey9xwI1YcLjSraiSatjKdsIgUoDJ7EfvE2D8o8sXZ
N3f8JBnOnX7vI4PFo5vBnIen28VEQCtpXFmxc6rTpCsGMUBRQ0FnA6gUlw/E4S3V
VJuGDrkj1U1rCofEz1McVZMLx8L1ADMch7Jhkd6FDPnnSmMcGnAE1CoIQmJ+aVBH
L8+3pfcaMuCJ6oUUZhQvsEs7hxx/uwIwm8UBJW/+VI8Uv889pjIDSjG6OYIGx/H2
V+eCyBsAp/qNG93SQopliP6A5m31fQLVtIIopfDPvRMUPGXqBsLwIot7MeeLD2J7
yHh5tp9ZOvI2zt8aD/U3BAd+78TK+T2ZKvZ2B/zbY/m77+cfJzos+1/oySuAIWBd
HxJtmVuE80tkiO2XzCHvQ6EOvF4u8BCvWKFn0Kr5WGh7PozOawIF9a+ls1Lcp6ue
CyuLYAX5ggvblZ6ifiW/MKBBsuKkQBOanyZzjmWwPUBZljlWOVXnJcnJe66Wg0bH
U2xPrXagsPF1aZeULQy9OvzbuWVEIExPq+/8KUddS9X8ujA4NGQZOKJYTfEWsvVQ
DRBMCMfre72PiLII+SXnHgZqn1z2gQRvNcwsF/gfmlAKiUbdJ2qqo0TAEMavFLYM
qmB0M3uATtflxMa1AuJGbAouth/GvECogfmZmVfl+lm16zTkIqEVEweKqrFoDFlW
YlAwCRVjw+zwyMHkonCkn8LRcLASGTKOp2QBUh2xj9E0x+wQfrNiOl6NohSoL410
ECyOWYV85sxy6kZK6AjS09vqWCH7hMN9pcNRvmi3f6HpJkpfgBmfbfvUv1B8MxlX
ZGeTldgw8bLvGJQ7F6mkJPqNicvwb5C3rQei3hDbBDn3BM87JGhVQnmDmz5vjxxb
OquILMKu0q8lq8Enpd9lvnE48aTSy8L6HhPsQCkSL7fMhkpL5jvUjS1BxrVwSrTb
QYkTgGRzC42peLDC499FDVxiYL/7l87hhfjTMbtyHZNr58GbX1HYCJM0GI+W/8GP
ArvFjZ9hd/k4ccTwrrYNkNbriBd2iImjLZG7DPXv6gleDPsT9hgBRTbQv7X9apFw
W1pLGYMg2LnXQE4B3uptk3tBBdxUXLaRyrN6Fmkbe4lp3ceQ9Bgwiz8a9D8hTz/k
cVhmSiJ7vciZUK6vAT3izfna3crgDcSi/ADnO5QhDsgtIDxWe2OdB1jf1l9lmemW
S9LvIpcUFFJaxY5UnyFkMfWEVc8vI9IMdaiJ8xgE070QFZDyZhqy7+VH89xh435R
KCyyJ2oarJ2LRxgMcQV+823L45TlZJGp+zSJOkkuSrQEXxGuCjmFcUw3PEMtHwyc
DiymLiw7v60mtBYxTaaejeu/kndTpqVeulmFCLRTy6c/qRaQQYS7jMxFAoAcSSyM
6Yjalrh+vaXXdftPbDFRiifyVhV2hkBHi6iqihgbEyHV10mU7NNdS5As++xQkeJR
DJ7kv9zekA9QMh+BojdgXVS/r3nai9vbIQ+dbzVxof6+3qYzkQXaU0wULxVFjbTR
s4x62i7+OtVt8JBK/d64rNFCkj8O+EAY1wzz/cOuNrKvMVV5DahV9EculgiSC0CL
mqUTg4/SGxSBbfKJ+7sdnB0QD8Ypnxnxon7+yavbN5p4ID3+WLb9UO6JObnNHYa8
vZLkweG/SS101k7YDOzxL3+IqJ3I8pckykEjdwT0UX8x8W/qD8taljBamW9/7KJ3
0RO9rzKgTbLOREFQJuGlGXHG7g4ho5ihYsDC9iN7mqEXGdixc1WKXY44ROfg9c28
hiYEEwAIKzfCQAebQ6MhXemG+U5++bTfDYajb8GttUJZXf02YbREpf6R93fwKOPo
3uKeqOawT9ZgqolG7Na5rEOe2vcVOnh/6uhRRVMq74M8iF0hVUwxYYfOAmkDhe6P
+EeXJ1BCv/ucvcTwbAHFhebb2PG/MsEpIK+w0LATnlD9ucVttXhHCevGUjHGr3sV
I3eEcb1MnOlPY4B0VMjw1kmMyh+3qOlxfUTnunMS1LN0UjESXbOVU9AIvtOj3q7v
3qZqpGEpQ3nQPIs6e+XMqJnBAYq4wApiqdGTEKK+5yQTqamgaRGbmlUnPFWETcRt
5xvPwA1m20r8pgm7Tv1akynkXewVWWb/GG/342tKXvaiLw4nKEjsIIGxVhIJDgOf
OoT0gcE1V1H1CCG24DlRYZBTRwzU/AQcgXb7nnCIXww5+X3Eu+c3igXtiDp4bg3i
c8WQ9nVeYm11DO5rOhjsNdz2OOCeY9eCBe2memZI1kObBrOzJiA7Ufqyg2AdLrEt
6N+kfFEea/kjeSax3Ci+uYcto6zbubR6E4UFMH7Fg+VdLYgDDLTljPl4qbfxFSlc
aLEc4qKYFQ8uQFP920kqme3QBC0fbRYmpxoWV620R5tMQuxiKpjUHjAmqyrFrCRz
gZ1bCo0fCbIjyWNRBTzkfYNp5e2JnQ9xF9+X5DS93G2khpXcnAB9jyCSTLXWAagG
iW3emxyP5LpczEl3oD4iDinZZ6m8A+sO3dyC20+ySDLJutbB6pK5iNdqZj+h9i7r
uFAW5vrlQZVM6rVR/GEtLexM1uLIpk/3D+rJXvDYd7MyNQZ2huwzDGyVxF80LFBB
JUQwJAzL53+cZn7a8rexCqkp42nsj5cfSqFc0uTJ63BeR0+pFz/SxO+3HB3CfaLV
tRjxf862JBed73TfyvCbJCUkNXI3YpiDP+b3E6jr5YGo1qEDQSeCjZj3abN3PCmr
uG+iIsKb/0Cf1a4m//dd0fekU2Xy7Fa0IJ4xYA1SX+aWfuVTbO+eaxhlg0EWoHnI
6f2rRmcvHd0xtE5ZBAu0x1Uabj2sqjfI8sRgct4u/3mI6szbneJa42n8awdgWHLC
S2LdMbqbLaB8YT/gtcoJoBbKMSfcxdv+I8Zh3sLSpPDO2Iatuax5m4o2gmaS7Rph
CGSbAB9rO/Uf7dPlpejcoLBd1f1MKzHZroYkIQ6IQfH8fEb6ammaoZpUNcdDzr0p
SiprXjw7MDBevJPT18bXtGdRukoEHD+Gzs6vM/uFccCVFwsSyPSbb3yuop1O7xmc
hO0QEKstVk8INQFCpAfcDmviL4VkAk4ahyL0gyd6OKjWYerpzD1UwwrX8C2qL7AH
vILbsp9xKT3YSBI0I9NL4z6TaAtszI8xRjm7AHLu7zZLoSI7X28G3ajQvwjecuzM
edI8L3ryR2HPcpJlBKuyvzwcdktTCCoJ+ohd1BNk8toohaucCVhebjBZVcgWA+JJ
MR6ArCNh7UBQ2GU7vAbGawT4VkKyxhypnlrfEjwnGshy4hiOD0+wgMEZVLZ5//MN
yTN4xdURpy8+P9fgJlgApoE6YvvTO3CUSnYRcUROPeEYyEf+00PJRIoLAqSW5sbj
Y5SNyolDEIGvk5Sx/K16e3dYLjrGQFFkp9jy/R+CbCcf8saSnHLYux+NoawhX3pi
3NRmf0sbxbAFhfrr6PBY0GI93/sRp86waYXecoqHuOGjUIruaY2OYjN261AOx7Yd
exrrQ3NLIo5+zxzZvkdkbUDFuPuikmHESf6Mpza0NWPdiRGPGBs4dlc0bTLIRfPN
hyE38SaT3Zklw8o5YMKsM1KudP/nQzcWAVunPI//wb6Qio+U2UOx7YAz5hK7ag6a
7UQd54Sanwi7KSYjR/pUy4Esv5de3j6JjWxA0xPX5zzZVU/D//F/aPeH9+r6oc4o
L9v0kXlV4Hp65LD07KBqmlyI49jKlUzCKfJl/TB+c8g5gRj81r91Gw7FojHiXTgA
5gHVSpoDY9ah46x/N5iI+uV9KFuK/YiP+2YuAYn/Y9KNdqPpQuQupkFG8Z8VTNYo
0fsHtoKSr+XHjdAbYvSx0E+0fKArf5ywlqh5nWdi1n2lmljQLt7KUFRKpQlU4BOX
NQuVKr4bQMwduEv7af8/RpZjOsQrqemC6Cbn5MoULoNMsSsPrxny7DOwY+9mVpGf
Xioqjb2HAsT6GbpFU1K+oRGx/qlExHz9YuyMPZRnKdjS0/crNGZSvu/D67Xd4gnw
8vPPzlV3//vorjvwwkDx+lixSj5f882wxEgQm1A2aPXnMdnZfv4vgqYD2znIrEcW
2buDz0Ehpu1mKfY0PTjmZL8qlR4yGhmWJmCzflAvAEExA6PIFspLHcWXMgH6/kfE
qO/ggLcXw4Mqj12n9ywYVS1UFv9HrTYo5poSrt+YFKC02uyQ2woZC+FSKa0ShnsR
6eabGqGY/S77Z4eRjMu0Avveb9G+qpjpS0RUESmPoe6EaqDhVXAWVtz0kT1Tv0AG
Dlw8g3Zcqe0c3hMT6Z0LPI8uQfQt0hgdfNppNRzIJ7hqmZsZ50+re8uNwjlv+rJ5
b2D7I6KF/eMs8gspnTngLreEVKUIw7lRoLRthdGSGmjol0vNcq1UzQfzsXX9wA9m
ZrOZNTKjpmu9Lt6pdiGtzCnjdA+rR8F/Jdxvw/dUugvOonQv1MicVpcOZDwS0ApJ
Xy9BH4Q4y1/hPwCaLPu5l2unQgI0cJz7gN8zTQHPoLVA8UG6/nwALBpEXtBV5bJs
Ex/jTwrJ1AWWG4S7bppuc2NiF6aKCqOvR/tu+1EneO5zCjpIkMEF/ihcl03ALL6f
NnM9czxHjnKiQcb7k2CxM05lziVecjcckM3qMstvWlLqYwGK0APk5C6c7jo82uTU
35mMGf174QRXEzCHTmIIM85duIOB52aOmz0yfgn59r+icN1YlXPFIhZSSwUIhPdq
vcMJv7EWBii2i7DEx+rekpz3AkG3owa1m/JtFffBXIo/5UxHszP/QOSvaHI2ZYUP
Jt7v65ofx6fGCG0RO137obrt28N+CQzPjEOzPPRkme52PIsSNCnRf7HE9c/ugKui
2LAmWcG7BZ/pFRCIaV8Dc6y2zfON08xgEXt2ofFtjnkoZqmsl33orRAKTCmGq6TD
lshutzsfmKj2Ygaq0hW9YJVO2IIJrLiusDMSRpA44B3KZ8iy6LTLPESOf2rER5oc
2TrBzxVmPRavwpyHdewedEo9tASiuSe06CWFhtE5q2nqCsJbf+RJUfnR/ncTnQyJ
M8x0jmKuL3xyo065H4xMy9Pw71Tf5GoQjmribiEZyEDmUjuEUETvIQNQKK4iDaHl
utMWD/8aa2nOZJQuu1X0n77Ggk7rPF/7Xa56/lRiKoV9OU3i0I47pc+Q2YVesDk2
`protect END_PROTECTED
