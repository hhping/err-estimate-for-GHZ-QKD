`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDq+/Wuf+9dFYVzOoV3KCs73i7jGYjQ4AOTBFBRILQJJDpH2pSKA/Gjsm5x6RIYT
Qb97nucMCNKfG3lKyqzroGQkwqBt1nlwiFlpaAjiRkOvK7zvWVEZyMpg5Ygdei7u
4+jbpbykEfQ/OSmTFegb/D6MRFWgPfFD5jDt89HjGIY1naBP2ovGtVcsqVuTu2iM
CnkzuB93xtjX8k5Qq/BFBda8QigU3l1qbYQAv2Q8z1QcGoz2IWdbI/BJKbuuvuli
bf4jKUxTBZnDvTLrrATQm0Bvn2x7rcHcBBQ6R2kCx/rGikYc1l+ughPuZc40daLF
wl2hQYRj/kO7QxgJg+Jg9qs+ZR/JW4pyul9F2Rd/135qVXNl/oe9jXH+VuejE4/z
IidDbFJOvTzAoInG9ObpvwJmEr19mlkBod6DSOvTsoCGg5zJU+R2u7dZPMhGyJfj
5c2RNViMF7cOL1DXfUHhvqT49/Bwf9ajiUBYfSImbAQ=
`protect END_PROTECTED
