`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q425KyEUwJRQBV6tn1MCFoXlGdF2eLCQ7hXNXoCRzeGRiFUl9SorJi8bZktwm/j/
4FMTxbJuUURjhMxn9Sc+VTrL8efkK4wbk7G0pHCoHMKy82JAADAdJNHPI6J7TMcQ
v1kcFA6XtmPZWooscyV8iJkuy9U24qhpFbIdCjdK1L/r56stixnOnYlxBiKti3Ze
IQJJgFRovYP+CI7KYoPO4VDN4ZKfxcQtt4hHTEspQBahPqpJL7XuOc1fILBm73gy
jdnM82Q4IeB1cu4GvEndoiN+4HROptV41+zqlfV12qCWCvpZzFoLkgYvwytDSnIE
GbjctCF5D21WrEXQwSfU7wCxrfbOowCHGLj3xUUKP23NHJQmY23/MEv8RN9LqDfw
eQYiiQD07nbKL4Mm4Ha9TABgCILFuDOVThInslJUwZ39hlGYBq05peZqdv9yPE9t
sBcKSfvw7wn/R8q1tMXCkLRUoxYPtei8aeJpgizwQKcIHLfHKVPWt0NtdaHC2uwV
7i4x9Z2+biGSF3w9CuOU9ZUhU1VFkZV/ZdzohEz2XRTlBkIs5i8SJk3NPsIglRzi
gc1QZgl2WTQbroH21ymdeBs4a0qEpsUoLI4tuEoXhbCFzA4FMQQOfYrstye40ULx
yRdhVvKFWpXAa2B1SV1GzH06G8kJCBdnQ0T0D90WFecf1hngPmEUO73xZkY6556b
xFDEQ3Eg0weXW9JhH4FBmjGLCfNQIHsLYIgMQM09aV5f9KWSTml+bsnE+eVpy1E6
J+hPDCB+GlFnySmzgJyb9DfBFzzX2ownyKNJT1vTrXZdEpeyGpKxf7v3jy+0VeQd
uBSIbHNGjk0wDcpiRxwiD7v9fn6bSUAcFU+130g1Kxtv5TdpZVfT7lqfXAVEschK
CWWrqtqooG8cbgZEprirzU+CfdJI1EwJgJ5B71JQTJq+0XDuXxdfWaOZ//NJZfPV
stRCjwQno5QPJ/o7Ld4EXeVOGv2Jxlw6IMWESSRdHJjRrw0uxxK5pkxlLCC/giOZ
mlF8+ODTKa3st7gl6ckEV/HHIgo2A00Q7SpMl6ywVzZVuf9Tk/nm6WqZKF96jHU8
ToMH7nCatHMJ+2n14WVks3//RQZRzaZ6dqs/saK2OeixSYuR/YJZLSgVF/Ga7KJ6
dVA1RsARBj+raGk50TKbDn1/HXU7xZqJKG0AhjeMDrfkn/dOQVPJoT/VeqvmZT/V
nMrZPfap5R0ZQilwKC3VEiKq3jCGfaY2t6BnixPP0jV5ueJ3S5KmmaT/lDVyVFnU
9BcWCT7EvhehoTeHV1YwBSFhbz6Xn31bn3VlAsg7ogc=
`protect END_PROTECTED
