`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aazhsINiO1OZeL3nxLUoP3Gu/mduDAtLWak30RU3Afzpa8C+iIAVSpK5KpMQQzKc
z6I5FHQF46PO8CEY+1mE/ZfCRk6d8lYWN5adEW2vGPAjslr2cj1TrsEjBxHrfpAg
Gtkw5nLW0C/cTqxZdMDkA8K9R+WZCz+NjmTvj8g/pCnaP/6SNUZmWVCIebn9fQ7w
6Y38GeuPRgIVjCP8QVDB+zXnSG9BMmD7sqjc8oYKBi+fsIPmUc5pTp2XMZqxa1OI
QWBLECmrycbcFJCqQnC9DVsUXciVm55HxlnPP1e/pPddgyDsDtmIsK9rDeKwIu6Y
YlHgsfUSIwHzCJrpuEjBLcCAXMn7ttunIVn7uiiebyZMNPZNqGO2XopJx9TlwJM5
EQSNGcEZqrylEY+B7QKugg==
`protect END_PROTECTED
