`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/HLKF5GuOeVduXrZ5V0pxeXXrisiQFpDpjyA3s3E6ugR/M+Gh0qwoz2AKfiPqeW
DJ0ygwpqgX2mp/YJWtclSS+cgil8rIFhUaGPhoT3ZAxl7YFWSD/nhiIJ5Cmu+Koe
jUtigayI5RwDpFQtO5m8XZaGXJ+voVohzt9aeF5mv2vJMJ9VzNcA02QJ1Effis+w
PM9zKUU2W/eS9uN3rCtpHzBZcXK3afWu2wEZLEtdTeeD4LT5XU5LJCfQPGdLXFAH
/s2NJKhpugHU8kn4q0wU2GzhkV6tFlhhNY6gaSQWWKgaSQXYEZozSp+O9YM4IZUT
qCm1rcUsSay1zEmClGTqmFHS0Ec5/8Xq6AaVn0mO6SkD3uIWJbPGcUwHKb0odfLH
naQonn+ChtiVsQRy+MI9vhTjjT5cs1ZL4fTiw5dUIeQ3lAPCk9zlwVf2sXXSrCqR
7HVIM5pvxRNrA3nNjxAzkSqc3e5nHUj5owBbSDFoZ/TeCTat4fpCxhFVtr47jNAU
4ZhmVTd0OL5ITICNidujUZ8T9Z3gVikiFudrdz5FQlWFjplzaoYbTrItEqWx5ifI
f8iiKu6YGuKWDBII4gPmcD75NvtKMxKxP1TRIqHr/woKGrIzeFXj4geIMzxz3VN2
hoEr72EP10sgNWn0/xYfx01TM8Z9KCNojqOZWmoFs4SqGZ4swrhksh6PjmitYTq1
qpwlmKwCMxIkO9tcgxqv1OR0iT9IhwjRdRgnyL7dnpjS2cAfhd5h7ZIEkKL1/OkJ
8pl1tIbGnzSfTGBjdHYn0VafByuIu8N+Fliya2PUnDXB5pU1C9F492rzE7cQCPeD
ub/vaeZs/e7gp3Dh7ZcAiE9cDI/6tqa3cnsorNa1WxvF+NAn8arkOzTmxTNB65Wp
3WQAsrHpmWQuoRqlLJgFPIIVgPbdjRe3OKkA3aWXQyVsiVlXcMYdmTolRmNPNMg9
J0V6oTi5OSZMo07K4nXbDXLnxQ/Rtmyykte67eQrxyX1xs5crBUq4X1+6CYx1sPF
zx9LSNip/lmnyZMxeTuf1dbEkFb2q53QuP3IX715ydg71TQERFAZFW6J+Fg/jNzb
WCeZ0XzfyZU+tFLKad5ABDhbimVseqPt/+tcDvjYKlt044T4XWUs5CjAbG1Vh6Zy
2g7PFq6nBJlX3nfgF0EcULAs9AsDy3og03+LClt0pCamtmwPCpfikfn/Yqmf/fb1
WkX8JoCX3XcWNknfM15Kw8oo7ZWftGT3uxOOSZysE5OBP85dNXQutIEday0ffmfh
0SdQXCAOXcf4cmVwezRynszScI523FNvG3XDnPS9Qr+Y167obEp7DZazJhw0RyOv
blobUwK7jPo8D6SGljZGkCUH8iOH3uTRKdAM4fQqjwQKaGdBJOLpkCw4qxfk580x
YX5dKFyxFBaoNzAykZSSmK4focMJAIKnskH+b0rMnmqJ7+KTq2WMGFAf9HeTAPzA
aoPg4tBrPe23XDWhkBZqpBEvqzYvtMguVNnaF0FgHoGc564E0Q5+LjCQLVS8wB3G
WOlNARMI11liD9RXW1kJW5V+hUgQzrR9SLegq+RJbCXYl7Pava7v2W2Kq3wGu/Kn
d5xJwXt0MkoEOBPoc9OHlXCdjILQYMGqe/k9FucAj/11obCRVpVgL/hcCuUZrBzk
hT17nyZ/Bv0f1yqadrEFdSv1Emu6peOBWJnUp9rC4E0ymqZsqUE2K017Y+KlexU7
bWsKxSFM2EOGnebJyW+5fciD8d7JzDpBw1LdRrZrLZrlymSF/hEaRhOcoN0rzfCS
6x/9IAylZJKAhjoHeM5qCf33w1vJ5MXN7e+40J1XbnmZkYYJtaBzpmKuioyzBhpz
U+ylaOIuNxnx85H7xOO1j9fBf9V6sIxaFLTsARqtXI2Jx3dASHwou5/sntKOGKbn
RMhZp3APZJtuWoPjMrQZg8SF3jOVWeAXZdX9FL/4grI+052V36mU+hfpUqNmQBNs
x19k7pZcQdxvsx9IIX9MjWHfYt+HAXhmTQzy+Waxgz5M2E2ttqnqG9M22awED32G
z/PxvanXQ91Vc96pkwHCXGUHHBgCV5zNVJDdHWnLGqXWOvCg5O6DuRolJ530cWD1
5hmKZpj28G7ZmCoaeVZ7Phe7SyAeiLmHcUqwVRp6znucxSAo2xngYFEKOMMFx2Rn
81j/VDMCD18XW5rVSB483OVLGQZNvfGU1+h3GcsNFdPqQ1/taO5ySw5xcrs2kB2f
Ov/r6UWsVq4ibn7AzRemij3NHyeGYcKH6KEclQnpUYr98tX+njuDKGoLDB95vjBC
s+OQ14U1Gsa4k2eX1gozot+GIdfegZRWYAdt44Uau7wlU8rPworEsilcLS4mo3cg
DDMzYmq0v5uCqdywl9gacTpsttj9teJ00woa+jC4NjGzMiXc0GdQsIG4vGPlH1BU
kjDELtZ8+UKL1VPlVsm1MX9nxPze+CTbfAXlpvJm3FCjdD9nV6R92dGIN89KkZiI
QGq/qN4H3uOovIWLXOZpDs/OFVQbwBGyG/O9fQo331P6ds6Nx/ck41AflCvBO9RB
dlEL4DvM3z7/yBlH3jBN98krr0Il+QmVzggr4XMKxhs/5G3+rswKCwI/bvmZkYb+
v59QSiunCHKjG0mL6iTsfDqU+6e0HwLk6hID1MJsiMGyxemnUNvgfEYr2I31EpS3
Fe2wf0RjsUkldrQcXuMzbMS5hBOQA97WqNJldAT7V2Mycf+geZboVh41AM3bOI4Z
XKcbBrdTBMuk6DoZXDbYYwEPHp5SBLIpAH4u6DcbLizd6TLroEySd8NkwnKgTtjq
FQymPFyMS91zAeiXefqFwy1nBXcjh+D33EBGEd+6UH0HxSG4/hbESC2B1Pv6OW2+
x629X2Stg6ftgRteqxNTyDjx9nmYf5lDS9h+g1d2zLMr0AdzAmqd1f1qaha6W9tg
5o/EmNSFtv4ehzm/R+EFJAxi5e0eNV4v9UW8LmSUJRNvyMNoDQ6+dEr4J+jA15y1
qL/7qCdvZMIhzJQo5hTsgklvINS/0I3fzGenV5Lrbt6hjZwVy5kpN63s9dkjQKcA
nBBBvnFeyRnRB47Vn+0to/wTGdK0rA9/9AtGEHvey0281IjzdrHWo36s+BPUkYs5
ZJpS9sublsbyMdwqW1/cnPVc5OR/Z0cdlp/OOscCQuj8H95nOvrE1UEh33NjCENq
+sl3J6BR5OzyGZxcVO4jsBH5Qwyo7WETionSys+1HAk0SckjiHHtYplZclyxNaLj
JqrllQR/FcP/YJ2v5beP32qJTOi/6efBE22ICo525c6VNKju4woLYSBvB47yjLLT
k7dcI+Z4+wLHvPo2IdMd4vGUX6QszFIvuCQdgudh078CbgjkVT5l9jZu7N36uX55
xa0GEIVUrHHyRwEiNAyIIFT3vb7jyEwD4oE48r9l9eeGmAmW95t+n8sAXNgDj/fs
nrd1NqHxS0ln0ZY1Jt8M8Bmh8DDxuP0nIGzPp2jMV9tO02eroU3UhNHsSq8jnbYz
9ml1t2rXvXFlEMqx+r1A7OHCo0ESqILnIf4Q62c6m8CV9rDRBBKMG0xdDThw7mQV
7iMOnLki5mEX8O8KSBTo8yAomeQAuvyOpfkgBHFBaL1vUKCRlw+ifsem2qiEsmu+
yFGaWQUM5WHd3DRx9ubKfVHeQsGpTW/q+TWGnW1PMqD7JD+RaWAfybIcmvxdhyty
uPtZsshGMa5hAwGwjwd4JoqMAEjDrtyz14KeVarQydTkaW6K6i0EZfMXoaFfGL0W
jw7oqFXAilRl+OQtHm6iex7tGmFxgFFSRu6O/UK8Tm34pJveXngRf/GKo5we+Gg+
GI16ioVXU69mSifKeD30XaUBey7B5p8yGPOzT0YX0YQZ//cDcwFrDhERBsqXE6he
/6xfLb7FPliDgHHEJYyc3JUit6A0jQXtVfN7Kmer1iFTxY51Ryc61v4sklf3noVL
9XprK02JghSluxFe3nF8Pxwbz7xWDJQ3v/lz4SLytwlwofGCqUlXwXpHmnJKy3mF
rLNRY/2Uon9eMdztR3aAYn6mmzxm1kjBoUYEJUyytM6EuUGLLwvpR2k51rIkMsFh
/ixKsIQArKamdPoxDp24EvG9xvvyiFTTTsVQYmqgwfw=
`protect END_PROTECTED
