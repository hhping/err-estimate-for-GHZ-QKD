`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
td7VYpXwNBsH2PMqNp0dRy//5l0pXI9lZPU5nmmfpkFr3fJAeRYxyBNepA7hZDN8
KDVDexWlW/eETxkYA+CLKQjGfPacciN9D3RsQhjuDzGHTA95cvSsge9zOgP0bldC
CbpDrQZh2A4timeIndm47jcsfdRxoz9WxxCcYFSpIVc=
`protect END_PROTECTED
