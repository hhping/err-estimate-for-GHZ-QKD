`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ckJWQ40WoiLQSU9Fz4wlAi8Bz+kvWNkEEUiSEXZ9qfStN/xbrHRIg8XB2f+si38T
BFvWe1O73Jyg+gKk1EpObToEwZrzRhqSz54RzwkKLcEqtrcO6V161Dxv5WJbKCqV
R3xsLdTbbMbnPdqjnU6rKINEEHEi7tw9CS2/cJOvxK7f/EJb+BwHnzfKnh/1NMVw
CPeMOstmb4/RzyjRGKNswwH/79ZoeLvNH56lB7IqUhjqafKOZWOUsTxJC4OAi925
r6m5SMqrqDsYxrqT1jjQzXc9SVn55zg7FQMdRNQeCCCheZ4DZnVnTEZ7VNiJj13g
lJ7jvQ3PFtdF1XGZsgVVwFq+RcnZyQ7e/6ZuN8I630GP0DO5pT5iSv3SvmR24OUt
eXKjq03KSgFRMffaIa7w8JU22xxiD+GDvxVFdhGW1j1ootrFx40Mv2nu/ty5s5aa
TsJ8usB98PD0OK7/go8Fp401VBsOz6FTxNbUnhXWTlQqOFaswbvRYtE4Jy7rpCOd
/DHKWosVHwZa0tXYHIAZQkiyt/9RJtDlEJkQyKA6wxB/dLlbyBwouTHVmteG8Czx
SiIrNp82FG22V9NoSt+Ab2+q+t1sHDwj3EMYr/B+ASZNI2r3ZWVHkBsg0CXcb6zM
hVHePKwps7cLLSGmiePn9pXlw16RZ4LpOJl2LFUcenyYaZVPI+d3WTUdFkArQFpt
+xU6C+juAbC7lLF6vWR/hyTxIWeYaPysTwz0VGZpliIiP47IqtZmh7Wlukox7s1/
wEEiphgdcq2Izqj6MGarG5gdrmzV1kH/QuHdRuHsZiBw6REiBgKILV/3rn9mOY4h
RhO05SL8h96bD2fYCoojw19eC4Ua7LBbPqa0yaCC93ldPpWN6TwlAQflhV1nm6AQ
Gnd8BcsElVmo8HyqcnRH0t71HlJb/bGtJCFv18L6vddyRhUn2DLI7lVVjPh2NFEG
sqzkwH75hpJS9B40tTmq2ArtjyaJiXQ1uZLj8AbRRBLNs/IC1ehWoDupAjLMCrz6
o/dB8OA0uyjm9yj18nwOTl+FuRD4b21lf25XpKwnQWpVmUnhYTA4WSFiZ/jU49XE
8D1TY4sbwSQT5td83K06dDRoa3Vq7QzN2KXizEsa494UxRQCZXpju6R5fSy9M+SY
Vj4Wj7njqAupMybuK1X6rqz+XTO/Jz8BJS9AhCk8XZPWHGkDihczyzBjPtWYlL2F
qNM8oaNpy3aDSYJHrDq6NKNLqbNnz2N2vBAzGKYOHyzZK+8O7a6mTveDzqj4cucM
Gr3L0easxZ0DCpmbon3rJRxLbWdIlLJqG2EYZstoqJVGwIs6KyjfdQ4iGi/CK3YX
wKdI04ahdrIxh3hL5BfB3nvdA16BMlz4nnz7fJve3ZS5XDDaXgPE4FoDQx4agesw
P4g56vFBipKHPytuxB9SXRmy4MQRfZaJw4vklLEpEgBKHFNWEf0mqbkszu1Re4zh
8Ur5tBj1UHpXlzQQ6TXyZwwIfXegqjCNaafvj72t8qEuM1wd7RJegoFTM5HeFAVc
ouadSDhsm3v737xWbMKcPrFbW4LE5anhypF4DmXpQxaszayudbWVJwrk9Kau/jjC
rsmXmXBFkySG7v0dWpUHmJbRSSoiSbcLVxPrgY44jwXZrlnnVu85aHaJUICzrMmM
/z4QCBZcgNA1iD3IosZ8jgVPQU30M0x8WTxoknQjHX77+DaRj86IQfPm5tkBCtgm
S4FjDSr06wm5A83bNebcRLsKRaTQLKAlERIdeW4YWeb3KMsx4A48kAnhIKbfhDM6
Yv6PtjTQLyh5SH7b/Hx/NJRDtaS3u7kTfurhs8lUILp2vVhCmrfS5bLWz32U9WwO
v7n3/p+XBsscRNoapa7arsxLXYbTryKeqeQ7h8RpvoZrCOwTttCbsjZYcog1i1Hw
PG1ZxhXv56p3ohj/TpB7MVcLuTlMoZV5mOaSOoRQzwiA7/14b5In4ZIoygZE7SP2
QhKJsXBbZwp7rfXipGKWV85fCjpsEnO2eJ4/QZGJVTtZsKnGRc6XSdRJ0qRrmfc7
JlynIX6AarzHTKFuVls7P7RH/8SmeO79NI1jf1o+bQThpqQ3UB+7iLxbh34cYO9v
uE/pZAtPj7Bq/dAteUoJi2tP67FwQMSV4lY+YMCDzimfON9+D1IeCyOsWX6Rt5d5
WuNJ1VYD3aDqpCvINJ83KWnpSX8SxAbzGvXr5eN5E0hDboRuJAa65J6K67jm/hos
7zaFVHvzeD0ayPh2XYw2BUF81tv/JkwrwAhoEP0MsJqbKwG+dGT8DDU3bQSO2yYo
TJKE76WvkS9rB9m/sY/EMfbrzIxweSikml5yQ/894ygr4cNRERkUIt5Pv2dFuT3l
L14T0b1vCQmSjWgCb9hxRPo6djbWZc3dgdHUHMd/9myr4RdWE5nqrIUPXyN+jNgI
1PmB1hgYT47MEPN1vNFWRx46mhJoE3JJ1Kt6v9oPLn68C+SHwcvlo1j3WfcKrU5o
DQRaRtt+Xvxy9dqd7dVHRBSZh1pVUr77udp3tUDFGlcDVNVLeN+Ufp8bdtAHSQnY
iyZ/tDbTl12dBppDBdTQq4tOxITyVFmn997oCrA2nriKauzg0ZCJNzgQ2goM9UXG
7F3FrdkUTLyiEtzKIAHRDcCpxBvnxhLJ2NMIRv9S6nZOGuMP8RbDp+/jMn02tAF1
abZZZLgL/XbfgDPZewwVx9SCCeOzOmd+Fm3cZ8Myqxk7xGZIeAmCcuWXXEFAUuhN
HpBhvYDQMz041rLk7w1/5jNgqNl+j8vig0K/rlalFF6+xNI7dWqEqNmgYQqVBkBZ
ufHFb2JfyQxeZPrr5btCJTNI7cU0nGvfwUzDssURXzNwqhNaQ7/IPaOF5OR6Epz6
t4qXXF0DQC5hFp1MxrPlCLmvAlh5f2ZCTzkIgJjJaqgK/Qv2mxAP96vs+LRuQf1j
Kcs2rZ12z75tSzaIbr7Sy0irI4rb5ZeMYhW8k3h9/IVgEY+oZWtadEkuMOQWHyUu
qgqDW1o1V2r8adE+DWrqUh3ut+8/EjQN3YoB77ko9P64MAVPiiNe3FEIyrMambiM
AI03DZJKLDU7mFJq0QS4vxUc9vcATKqfc7uNRS6O6yE1AxPLZlZ4QL1F2fUn93g8
EOeHvKO9RN8OODB+8rlsIB7eGr/EcOEt0DCLBEjC9oKo2eq52jlSq5ctUrO/GbJq
VRlx9+8p26xpcZKRKOY7Vw5lyckahOpKje+6AiK1MRGs88WgxV94OxiH6jfDRZc2
MOm+Apqp08SL8G8I7uMgjIfDjjyFWM2PAU0oAyOiB1Hect7HMzOp9P7Lcj4ElgNH
c8HmrIiiMGr84YEJEgio1XX+sOxoAiU9VORE75fKglFKoIX8N+lmsoukpv2yhv/C
Adead1ic0YG1nOVlehssLfXokDcL4o/SezjH5MKWWYGkj0MXkYo20sYqk94QSeu9
X2C9aOyK4mJAuY34bturAqJfgE8Jmch77An3kpXy7q/e8FQYMYp0L4ypGyzOlq/P
Ia6Gd1bbgXBAK58gJSLzdPOaWC2iJBfZVBlczL2RKSIwl2CyMn8LjAdpQVXJLQwe
O9u5O9U4fwpy39FksJjOkC03uC27lSBtO+whMInNbC4ZN7IMNHZn6ch5zu55Ecqd
dN0xYKAjrRGM6WkN+zLwwKSjf7ZW0dJj6lsLsegZhbW+PYOfPurbGov09ftLf/7i
/pjS8griAXRnIUxSAVICVM+ysDr20e7fk3ZREYoRm3K8p/ZTg+SeSlADVG4VSTvU
TQiEmA3dpI9MypnzCbzwo9ElrJnPRHYLCaNn/GMrcLEFEoYn/IZ9Vc+bDnezuU/j
95rz7p99p4F2g3WbNy5q3/FsHN+hpSnTgwvbR0H0okRU+6wfzB2uCx+Rf1PS+vzI
MxyVlNl+DtMUTDifA9U7gCFsU3zYjva5b1lv6VQTa/huci0iM7ifn8C+qZPNYunT
G1IDRoxw2MchizwByBvo02q09MeCmGAkmWtmqr2gP5UM1xtjF7x3KxuRzSpixZRS
VwT0mZYHdpFksI3kReAq34aWUHqwFKKdhbcWzBkVxaZ6LmGCS9ktzbRbu4+vF5R7
YIRz5EVO2+YJSOyZ3RsiilMkhkLC2uC/rLFoEixfGAwrXQOE7WBiVQ0GgfKozrpB
X44dwnfM0VvumDucYL14jrktSF8tsC6kAaQAt9A7XVFX/oy6JHmJywp8ePd3xU4B
/wUxhUrdn7By+F9BMZAZo1s0GeN++yHxJ3Cfi6Nz0oLXXHgOvcP/9d0vWJRP+LUr
5qp/S1qn+Zmx2HiCpyI0mvniVP8FGdXAX7XU4X5llQObDs5DboplPsHNRa2qxqtY
7oabGYdedz51Y3yeK7nPcV24vEdAc2BgyP+bgyOCjl+QNPgBUlSWGBIsvapEevxI
tVVhKkIKRxcHMGZXtlRZCHU7RgHJrOsTsx7pi50Wra+yr9dcb4OHaajn3vnLMSmt
um8dt3YR/4++opPndwy8AVuLCtJKXYMFRRgadbqxz1MuHKO/nwMjnVSOVbrZqpFY
XipJfCPXvawEyLeI0FG6tmfX/rjQ8pWtFcmNOwP+H4eglo/x6ihegSkxFRgTrhhT
lUHFdytQRhbMYE1FzU1chjuc4wHENGqbh7VImarwti1ghTCrb3dXfukOLaXBtNWX
ypkZz1SBLcgR3qTxhCkAMnyeoNWNiMMdGq0dwVCDQD3zoZrYIVhLoUYbOfCoL6xA
HUQ3pBficEDIXXSHY/ROc8O/oGlLYwErqbjWtxh7IB0o8Mn3SzA+G0hw2H2e0d8f
4uIrHcQ1Q/gO7XWTcRUFpUkRPmcORNSiKIukQZluJi1jcN7jjcNSvnwLmZV8ICls
asf+yiHlT7SNBaj5rpPP14zQaGhRV99JNZpoTOpNH7yhiiNwHrTtlKrLgBz6gsba
SggrBgmMjx+qHEwGCknUXr4IGcOoXRHvRe4jST+wafvPnRMau3UPT+JN67qBktZD
pPvp4vbvbNmyHJnxgmNnxpsIIMfyDbuSnviFY+ZmhTcNZ/qQQGIYTZCyyXqh+Qwf
nFw4Q7Qy++E5XexfnNYYGApQ9+0He/lYZ7Fi6cmNMi8w9kn6hlQ3l25EylPxHzDc
mA7w6J3t/A4C37P/2lnjN9IeRyfnp6gSdvY6F9vpEvZYi4Vtte+g3+bF/D9uQ9Lz
ctiuQ3web6LUuGzd1W47mNzjbFODduDfmWtO2mrZvFR6q2ovugvz7Thjo7zM4eFy
poywsbQ+9MnoGymwivZR4lka/zcR0DhI+qxs4NuDF5MdVkvmanmJFO67Mi580iW6
XQNmlmUlvvuLchY88q6KQhbybXZuUgclUBzzg8E+3zZyN35QfI8Ep0iT9+dWQAnG
LyTCQP35je68gnB4biRxNhhROxqOoFY2UMNy34sNonacHPkXjL/JgXofJ0lvtLew
fCHdUw80ePDwpYop4RvHtDQuqTs3eu/YcjN0R+QpOUsIRg4QEkAAyl8Q/80iPo+y
rhf0CRajjRq56lt+mLa7LS1BP3M/HhtecajqzlAN6VHdnadFumesf0sYN4pNOcut
J5/oQ5A+19mF3O3qe6aPXHuytw1StM9U08KMFBs2g/kVyVxk8owGC3PdWrRDadGh
SXdt/1aU9R8llTQF+qIW/N5kaDB9od/EItElSX9oStr6RdSeDuEWITMa4PIu0geQ
GuKK60cwlYgiScYaW7B9TnUydEemJfiT6DG+lVyVQzQ5GWKQYTCXFJGirVpiN/JB
Lg9mGaM4uGbbNzHY4teRf3hsPpXlI9J62+lcXup3f8um/Eb06+kKto9cbAPu8IGY
BeHnoXAi2dtRvG2z1XgzdHa4X48d4BipweKr0bimu34vtgcYVIBbKFB+J9c2QV2u
CK6Esfy7dfaBLa/Tvr1yIeftHIXQ5DFxvYoeiIYfM6Jxlq0Fv3EzZ6dV5zakZaBp
AMS1mYg8ZsvypXeGU6dUAFln6DRH1HQeawCozVJ8SiyGsmU0NX1gs8d541RUC947
ovLc1Pyn7PC1HZgvRPPXNbR4xZKAUDZuZCIsoOA1oug6rR+NFmYwQhJtbL4s3CDt
l4VSveNZzgMNNKPZ7iUmqpDDdL5EC/Af8sy8yrdmCrs/UE+D2JZyI+hup1oW36kG
a+GmICadd79rxAvCeXjrdvGVYNcG1+WkQylVyOA0Rn7CVLAUYstZAgMiQbn0+NY5
8apY7ZCuX41hRCYf5L7QlGNZc7HtLJ8stx/am+t4u8gHTZ3E6Y9mvKUWx9dUIpKs
aYD0grvErEpae8koqi/SZE6fb9IgoVUtfKeoIPiREttkv5yK/WUo7QZ4PT4rgI96
tjSrrncIqB9dAEn25/oRLC3Hlqi8ujcuZM+xx7YswilTTPEf0mceCI5kjC+c70jK
NAGQzNrCZXkwHc/pEhaAM5c3aBwvhusTnAjSGKLrEMFUCGPOWvm6M7qOPN3J7iLF
MBYnDQyqrhFD/cLPqJZQUlGvpZtkMMS/coz6drWgULQ1b0xcBw8aVP9P864TphAi
veyHiofQac3Do9qhbVd3phNrMp45IMuX57zhp1eGbmsII/cgbtZl7keQKBgbAEzS
kfyL4L5iHw8vKfCbhL5ZAD1oy2+NdleTV/G6iYFBshtQyVK7GUnpRKFHaglDBjdt
vVQnzyDG2V0YkeB9SRKA5ZPzGJXp+hfhDWUEtcJy+AyaM0t2WH/pyG+GRky0vJUE
Z/N8Y205Ss3h5/sYgyQzrQbaGb1pQFsayq/YgKnqpXvZv58XpfsbPdl88oJf0np+
XxWA0jmMHmHRGWSSsQiUFaTcPUnjCy/JsqiGiVjg2FtfVFgusQCnat8sXxjB8H+d
PuYHHK/FpWrA5eNIdQxUqOi1P6ZAd8OJlbp2f4JviVVs/MtAu+0TyfucnDa/S1io
CSTptDionqNOD5fxtD/A3UW9LL5iReh7DB8fqopKpIAC77npa98DpsqGFW0zXEyv
j2xxrjFo9wdYOr9ip7ayPsMEol/uwfXpY0OM8tIU84EmlF/HtsWV5KHauQniBdnE
yfUEzHeiFZ33tTGzXCdwjmQjrQGKc+mWBUKbpTiAiiS1oETcbm4/cJBLyzYbJ6RM
djvnFqh4opcuavaTV8sOsFI/9mTGbwirLRbaE/rIL5FV4BKAXt72r2b6cWm4+sz+
uVURN18VtIhl7c1cIVzyA4RjPRJPtta9u1GMgY0EI7wtmDjuwAo4I+4Q97xsJTO5
m0kbFFBLlp7FyZKiNSuzD6BY/ka2+IJNpBvzk70Ge6nFc3gWTwC7WKpWzPS5GN4y
pU3vWh0m1AJcgXL4BTmkV9dtcdlvLVRFwv78qIKUU1EyXcfAH7/dHl14u7Tc4Gh/
Xw9Tv+Ih9dipgVTBTAW+fwKj3LhSvkqjtqDkLg+7sPF/WT7ws1DqPAuPeq9EorSC
te27n8JizHW5YMTNuEeDJiutNM678WD7IGqgcIM9E7+0fVBX0fcB7UHUpmA3N4Nl
zPDCj4PSb/4EQlZdAGThz+ApCwekGbw4ukWS4a/yCaR61HIkBKzYigxtnLM6Vpkn
68fymG6i9yNTteaWT6vWcoEZm1nbW6HvZDl6j71ICO1hPTS3dgC4FNHa1120UQUh
gXIXq0pAxROKRuzrKQN/uguICrwIU/Y1AAD1SfGMq0EDStavBtv55ZJxsPhad5mJ
DsBX9wg9JFnREWWkZGVpfeke225mjDjLm0LQOPnyNeJ3LCVNjz7a0coUR89hRP85
fMRacrIF0ekV0r7ms4T/8IJLtwTJdvvh+SnLjU/9gwnvU0hA1oYBFl41FD4f07ZD
IQGn2s/oEm+K+F75UOiZxyxc5dGGXaNVbRVnxKtEnu2p5mZEN5za5+G73cq2X5LW
ReH2lYnl14FjW9AKeFh4y+iqWUt2uT4psZPPuiqJYThUIAoTSTvtBNi8KX3JoyxJ
3UVgAy1po25dsRjCdfGfaCUrOQ4RSlNTVHXZglFltzL4+eo12AZTLi2akAo0Mg+/
7m08l0x8hpW+Jo+BdWYddBrBy/sjPSAHbYP4c01i1q/u9FB1TODcdYeDF9q7lUfT
2s5k8THIf9YV/iX+inEt9gJiEJB/04ffOyg91v93GEsh3GoecsGcsG+ke6Isfw4a
MSZ5NZ5zTR9A+5DOjiaifp9ZqISY05Rm2Te26BzYUqTtFqLNcSGYhMe78hmXbo3W
rR7wyRLoKu4NNoSh/b1gbaOuj8fwNv0yIcqu6aVWe2d0CmrKv3L1CoD4kevkahVr
xpIkAnT/AYakO+TEMdNnUU39wTV/JjZxtMRNSHWLU0bf31ZTOtTQl1XtmNExyqaf
Mm7Df51I+/+ALvueyMyMMSopOSjK5ht0dyUjJWsIU8h+BKrmDnYD1ol3tAT+bzGc
+n2Ja1w1wNSHlAmnNajO43TlluyC/BOTOsyb9rFdaON/OeC3nrBgCa6zQ9qf5N/9
3OO/LcTlYj0XLUF1FvKf7M11kUSomaC1fXCPxNbr/OfTQ0Z2zF0TLsvplEGlJZpI
iai9nrm0NM+WFks9ElDUAFbHOeSf4okox5m3ICC1W/0f7wV/8VB1ULm4aF0ATKZe
EkfeXZFZJBpxMfn9g+NaAXye+rtIZif047SugOKhhcH8cLd/PuWktXjQGKwWDzd3
66Oi80fCxa0e/EUIgX2zho33DvkIOTDSZOmvcWLhuxkmo9taocPY4ocJPWMwj3Vn
RdzYDJGZ2rOcnEoZjUQaaFEcZlFe8QHdR/8EmFm6Ed2X1kjF/gbCTZiZws2RP3dx
wyeH3z20utzlTeL36d5ei/AzdtIx5JjBg43+0HNfAI7WmdycCv+jrbY7n+qeuZWE
Cr+5NP9auandVxHg7tvdqJOlAZmvwK6g+0+CiCIkE6JZFw066ZU+zQC1mTxGE4Vu
UjdYH8lu8CU307fwThhOzrfIx33LAsbP+Qk9rYuQukqZtk+yqPSlk2HU5r12y1OQ
aeGOXJQeZnl13xMdGhCNB/fYUn9NU4o6oaa1UjvY5FlT6KkadJhVyTSEFwh9GMPS
ve01hGVnQ5BLms/rPkRUUDg+7o0FPIi5mx6kMZf+uvtp+JpQnF5uIzdjAcwiQOGV
okso473KISKCLjEvwFoVcVtidEaEMSIGDltsBUGHvEEKxJxoLbM6GudTjdSUauNk
nRNM8Xsq4EqRHY3W6jEaNakHCUznjsPTF4dPdQpFSjt8IuJNuKg49kxALCjsufjy
QbZP4hjkpe76WdwXV/p01dvHvnUMmnXcnk86k1ox4A5CAE2X+oTwOYuKfbCIvT8O
nY/y2hMPhxh4RLpkQsj8RDjK2B+5fVfOJ1Qh43Xvqzi1DRGxmsGWxqNxDZ5gcOEe
xeZ7hzTtnbRFFyDHS7/6I/LT4HIsY6WxCjtHJal+qvfF9MPHM6/HibtFQMja6J/Z
P1AYyuoqApPt9br/aTP/hztRej7yNFllypkVeUajvH5vwDVa7zQKR1rfnGbPGmUz
1j7AxWa2UhmtGZaOXlJ8LOKn+++wl+23A2ykSTmMsDIUy0iWs+iGdGf9er+DAocj
br6JSHQjB7ZEG0vE78TtUeFVyQHMyG1mitIbz7Kf+/qNYHC48p//OtRXuzOzkXCp
71WHqttYAFOjArXSp/UihcOuA2Z5lJRuDVFm0zQQzliYDu2HoSb46kKMB7Sm2wWC
awnotEr6aJAAUbJOhELI1456CVnl22FFc7y5PY4pgv4HDdYI1wlK6gfBlM6pLCuM
ZEb0TwWx8o+1uOek1CIHtvjKwyE0vLgfs31YH4yXsTq/17uT3rtUoeUrZGHEJKP2
U/rd8m5qYoP2pD019HikNTUgbnJo6a3AktQLFbgiCdg3yHykVfAtYFwjP8mh/lBR
tLLnNX7JiruBOozlWiaBcYRYNkcrjdZj29dIwoQ4e6IXtoVKweXU1j+KjPEiQgGc
fAQgV+8DqdVzhXgT9YBJ1tsN/Xc9SBttEL7rYkPD01fzv+Vkx5qM9wqemE1Rs6WO
crhNgmy5V9NQjYN4EB89MpEXTzhQzMaP7CCAiHDgKA3Gq9H1iuHpPiJiF947N3ku
Q+WoMdUTYJtq13QC9EdOOAkxs8FDtEj1vY1y1OTu1NtzdIV/+htAw9WRSTDY4Br6
kkkW49/CeHv13nKnYswraVmLj13F9gU3IXUOU0jeOX28zWdsNgjj6WYoy+JeKsrb
2CGiCLLkUM1SI+3a0JQCs3ipqdLugsymGBZMD+rLrTyS3e/8/zK0Zv3S/LpsbSbS
OyNk/2et8x4ClzmydvqG2tZ2ElZFPA/OUWLViUO3rUWVRDmZ5DWsOD3zTPiyVyg+
VloYcDfD2U62V4wCsotbPLT+EEVOj/zFsVNgGuHmrtIOAeQhA1L+YhaWGxhFTz7r
nZwQQTcPVa9K41rDH378QBaREL/YAJxN4z+waCHQGsbI/+feWCJCUfClUWulY+B4
mtw/Kv06H0Fl554pGuKJUH3qryow7af/5SkEVl22erEgrMNiRUCEuyLVpcehEXKW
WX6pbe+wkGLKrpP8dj1uIWAmcD3i/eDdGGlzsvJv+19gY+7hPv+Im6Jlj1enyjsg
+BEa+tMlvw9gPhjvESg2uMCLa/HlSde2pQQ6YZMz4QPWUBRPV4+pJAZVtjtsXuqh
DQH5b5jtsl6j6sTfIcdm94OP4XMqw4ex8AcHAc1nqYRepIsOgFzzF66J8mPKAZDc
ziEn5TQ2D5ymwNHSlOCwHrfRLQu8+c9tP+B/mPDZLl+NPJIxj1uN9/3ZiuYHdwmb
1a90paqLEbIMWwT8MnIsD8wsHQvbOydDAmJQg1VOvzfSw+9ZOyfMvtbfXphLRT9h
7oM5rjID5QvJHMKBDqkBuxTtjLqqRL8TEtYjqxjfcPNdam6UmcIpbyRY2E4Qgjl6
7RGkNmPnP2hsBUZWUU9HVytdJGl9bQEI2/vM55zANvh9qSaDM75NUVK9LFcnzONN
69lVb6bDGDyqBsQiWxmvdcSwXPS8puBhPSPDpYe6dCTSewBTP5RkjmrxAVBZE6KJ
fUKJI44LqIEo5qm8jQ610Mr/f5MFeM9EzEBfIQzBagbowBd5I/dCvnQvygPNcLjw
kI17rnK3Z6Hd0bqWIk7RQXKTy2Se3NDi/oTR4omDS8u3I28gojQLpL/04EwU/RSd
gx4J8XdB8QQpx2Ef6HfHWfP5nAbma8vEbC8Xk2prfHTqmo9srFP9jeWvAYzaKOxJ
x8ay5usR8hTJB3KY08NVvWWktWeI/MnizyFK7QvL8sgiFSkrRFHYf2bwoMgA+m13
5z+2mj70k4MOM6T4oC9ttfwvF21wv2DLHR/ENxjhFpHgbXfh9VvL4DyB1Sl2jvkz
9sr2lLOXLEeD5yja3MT6RnSuIs59XDX57DXbrKjeRRUttoTAUbAShckKO0linQAF
pwNsMNlEclmAC9SDFDr9yfbCrY73ZPTuO9fPlLMSK6kzmb3+Co/ujyAogCAeqBiv
Du0/fX6XnU7f2Shyk8qNlXVzcQbFPjqlXoc7awEStJ0hzWq6xQL0U9ThSB7XNhBW
4MClmuFs1x4OYMNEKgyM51rigPgestvJSY9eZAXWlBbeMW9wvzHBHefJ4SfNKDyO
EgrDhPRxtrweG3RwginyqexQ5b3+PP1/Jr1sw7ig9n8r6fdRD1XH1zPwW57bttE4
c9YAVGpxPqsWADeSc5+WGMqEPfnAR+CIQ8i6H/tKWIoMc65AyxU7xWk2yimhgzrw
B5wqgvt9qtwXPiJMhw9dMacA9/j/hMJlB5QgeLxHKwGcENiBNJlPdHptmyzAY+/l
Yiwt7wPK8AF++oHH3lj6bKQYoiCkwTxk6YyQFqaqlF1+8wuu2aY58VWPkOyxTQZT
Mgq9cBse+P8SU4+glZM2MyP9c/bk/3cFFkQXD7CyJYG8Z5BH804e/g89CJkmLteP
+QdpIxCK+tDhE1+mopKpjJBhGG25PXLvKJJwDGxDzTj2ilO4eczu0uOUg6nT8Cz+
maSj7V4pkBRXJjxF54lrnzZyztylpwrWG2rpqRUKrTXcM4zc3yUHLRmzm9FkDpxs
dhyYz/22lI+yO014BDzhrp9dN4tzJTjPvKpm0YSD4916n9IejfGpFXY/L3ItvV8B
RzvZBWmfbDzn/z+Wn7sJ2NuYyk5lVX0wPTpHxRKBK94Nni8HLnkF3aPfY1wRFiJ/
oEpRoIVKMgAutBJ7PFYGRILmI1puMeQGs4Jsdv158SIkPapaDJKOglMGbJpBU/Hw
GL2KlcTsp/jZpNAfdE7Degl7Sp8x5gqqLigOSgIwGDvfSauDH49U7Kob8Z4M/Qlc
mhB9Mvn/uBF0r+wmJGMROkL+lWLzIyMpp76auimv34C6mAkdDQDyYvaThi45f1+m
7WXlSyjMV4mibKQgFrKvAVyThcxcTfolWIoeqy6cSdv2W+eXBVn2w24zDeB9Fw+F
8su4QLRfjsyI4O1R7PIP1wQUBkU3OXOb5ABcWu9F7eaxgX/bVG38RdD/y11LTs4I
klwntI9ehH0cUDcqhzr8nnaM7v7sP9YOCwMs0A1JYwhZrixQKGLXtdNrzDGLrQue
IG6dlFuWU6VfVVy7xv6cBRSULaiMHTzMNliw2pn1IuFe1bOCrmmIVaDhFcOoxCFB
bdbsiFWvnAFpIoGg9tRoCGxh3n67ErDNhytle5rWdM8KVB9h2VUbbKdq4jxWHhuY
Jch5A1Ex47TRf3S+NLXKcwoE/rnoqlB7lKKq6rRT0ZCimui12/tQIngY1O8SlgGK
rBJ752eRpIJuvfrtEowPlYlfk0436cxMtO+02QifjEke2FXWfrhnMv2FPTM2OWxy
Fou0l+y2vjxZ9TOAD+3A7DlhtrAO/TZq0Io7zlOY7wOWfeh+k1r6iicknYtIWjhI
A94E1hTvYwBDxo/f3VhHvzBP0d9ugqt4HFHdABEg4EgLgR7z+6l/cCbjvHd5/RVF
EeMsdck8Bymofea1/ernGm5jkUZvij9wQgsU7qH5cQJ3BhgQD1Z1wFT2+e5yMSAC
eqk6K8jEXguJnc6tUk3DF66jmt0gPMKHvb/LOLXSIxkiAXUvCDY18BVoQze5Pggu
GnlvwcuTIDewAbrJYAqlwag65iEJ5asHQyHnYn4cVItdH2Y5y3e2uPj2ahiq0M8C
9Aqpc5o35jxqwS1XczHjvLYTAWYlhIHY+k8nLZQ5GIp5pihWRUCkUw86ymYVLgxN
DCnGX5bXa/zfsJ/jP9eMWgg6/GbBk+mL78zk/tosJNhhHJkuUMpQM8oJJYW8QOy+
GJl9t7t5v0924hD15Zqmj3pTVMfNUYMbZqGSxofzEABwOh6yRyhYdgBwiY7xlhkz
mmDNKHBT2SKczMv6lmVdSI+SQ3LN0BMjY6AGCAKSU8yRrk+fhY67h307dz+UEDjG
A+wqVeiEr89GIVCEuJwS61d2zBncCe6iHFroFLsYLW4UAa9TEudN/yvVVVSq6Ye9
yb766b3bPz89+Y5EYzNdsLzcGTBp8xdY4XpyOkz0hrZKGteGMD2iuMR1gVpIzqrm
v+55RBOuixksrun/IMjzz+UMiRHiiZtX29IErKZ3iBpejkLSAoryQ2Wf8gev2y1J
l1CI/q/cGEC2IvH1yAdlHa5GmekZeuu29Usjh8qO2RUmJSo1YURigPnU/j3hztLE
F8hh17znD54HsPOMvFJ/mRaB/Lp+uGV1XGDrPOr7dHPfZxvZQUPzdpxb5C4McZBO
s4rkE6meMVii5WCDxze/QXkxrNj6+2dHlDCElqwAj36VX4ef1/NYzRVc8IT0co1t
Eiqks6LjqNCQI06y1UnoaWOmK3JPIEAr6zBxRpF/98xyRlwIe2NJfLZ/6pfyYrfh
MkY2rk/unfxAYN9czFBgGVBY1tDiAPIESIPWLdKl7YO/Faq7QPqBdv001ZOBOHKZ
zzziSjsvmoyI2BgxyJe0MqrQbB9NefkKB0/EQBaxCiNCVF+7FZ8HALqvAusMO+Ro
fd2FM7Z3Z+ApHM//VWsOtwN3JM3RIayNFlgGnS7XlcI0ZEyzjnx4eUFW4OT0nBsy
UJ5vD7tCYgw49MsGzuw7XmPfPlZagZSTsyFNlfvKKn2wJsqasGtttzbmo9CB37JW
wqKM0gmF6UIf6uAvjLK8QJc7Gk3pL0PfQ+25h7sACVsHpNhVe3s0y0O487hcoaOs
kBSVyOYIbCfjkePAd1Yd1frzAK9HN/wE8RXEcnH0iKGbkuvtbai7vESZIGEFTzoo
FU3aClsPZuOAk7G/HvhC5ApWOkHcqI+RwAP7dExC+I0SIJX/9VHIwY0+8jrsIVsX
JOrEXtAdxtkJ1Qt5ppl56DZyjgHXMcEMGAf3v0C+2Fepj7tnbHULFKd3h0BumiUL
tZUV/McnGtTPdeg53dL4foVEaVrdMSTgqXqObScuM6xu6jiqluJIGN5di8zu1gDe
TTgseNsq+EaTPvlGkenNu9ykvfbQAjRRUOtfmfQnWwbesHzfBExWNTRwKufmqgCu
B+xFhoJKENGOdamS1dIDpUYCqC6JQOtTaTcUmbpH3XcDbPhx9UI+jfzps0yaBzKj
cwFSV5aB06Ep+ofraTGQXRwWnWZmNHTM9x8m5Lqs492sS6YSF+QgAWM4ApBB7Jec
rv9gx8PqZb8C08B1buAFf0taneEwdyA8daPQO+eX1uBP9VzvgeUFskiHDydNqmV1
AG9RBuwjOZPWvE6Z962Y7ViAt7jjvdFacc8OKYvYCEse6M9G94VaPrWSk5HDipzH
XT+YlRtWcC53s8PaRekuD9pUypOgM+pb5LUHDtVtKl2wbWUUV6wIGA1m6i8X1NTc
S7r9/LRzW+IupsohPoYd+UlPHr3ZWg+u8gc8uvpBte/vYWtEZCUQ/lRZDP9pO9/V
Y0xTn22octFHU8bFMV6l7pU4kW0YTyEb/j2n170OqsvJBqDY3jEvcq5j4Cyr0ZPo
rlUDYhOW+7UKPW9+r8v4xMyAMXAzhS20ZNhN0ii5fbnu8wIWodzqZ7fnIYIO5FHZ
yhB/ld7uhaavhx8Ui3Q096DNIOn92I+fvg3RNtrwa/ei4fO1A4EYDuzG2W+PbBv/
+/tHuX+m6By/a5ep6iPwaSLZTn4xKfSckvbThrMwfikly89hLOSJLGaFmueqohC6
5g1grfUEMEekXuie+NuX4Zscl3rjuMJ9m5votKMKBjtrq+IW1suHr5T4l/2fT0Vn
vfJ28P3fHDQTknCoSpnOKgI5Kx7p5Oi9rB9EcUeDdgbQLNCOi9xtsnYjwTaawdgl
NTBBagGQaQGUOHIWwfDPQIVdKqz7J/mOm0ihE5FXgeL/B8dDlKZuKDODVLEectfq
ypQ3Jt0VJQHVMsXHiq9g2vXRh1l5lCvUUIal/Cj92ilAzXqVmzl0vnFceS9a8dZ5
dYvB9rBRv/sXuAag+W5jPp5tlqMwE0e/qSBLp6KoPHAs2Ns0MwHLfB2ukPPAIfuP
Eisq1HgoPU77sGopCgWUqA/WVLzvnV8n9K6il241iKXW/EJ9JwcatFBPaxtyvUgL
yR+CvLcnE4ERrSF++TdRw29bkflT2EAGIDFHV/e8v91RskkeuulpvY6NJ69GqTH0
iDzH5e9Vk/Mh2HNaBchLGxNUqiagNL6w/nCu7YMRREsXU6FqEyOp9PUBusElfVhT
FuoSTZiSZ9YDkI1eOc3viX8A5qcs/fgNYJLIODNyu9kfE/WZTDfIHwI8XsUkP6tj
N5hDGJSU5lHp8w3dWGhJrUBY15OOokz6LXv6AILjyaF2ioENQT0F3I8YCHMBFZ/6
IYRjfrXdgu+UoYDLXdCeyBSzzH/5c8h8bEDIM1OF8LAmQkYE0aypiR89a9rJFiHS
aMh5k9y3zC6MijWsUrLgO440nQwiDfk7VzykT5XJv6pJB0PSYe9rIVSiExPhAr5n
xYR1HFrEfJciFTUEB2on1n9fONkwQO9qDYBosIXf5GxNcjQout0zBDamKBOYEHM+
VmB1ZMQp0ql1fqMtBnJnVETuBZHmFTr80K20dkl+oaJS0SG9pD7vICNo8ZmQXBbN
zbMsfg+W8kju5pfl+FpgZU/5r9FmV/0gg0zBMgYklvfhGX7WdvsmkWdUe/04lpVL
QBJtk7zenQerxlTW/bsQ58F2Vbf6M7WcvuFj8tXjDhx4qoqiZHeARnwt48AMRqV7
7oH2Z9pvKHA7TcOq5AYx2TAyV8M5fHrZOl9G9/ZX3tzQ2A6O1QqLeD2JxPkXBAOS
ZexnYnxuJguZmddbOBi63yywEWtVRh8i4omXe77MQxUyFQA3U1aNQ+774h9I1DD+
XkwE2HdixHE+AoULhkbGSlMZRZqigZsmwOOQFt0P4DnYZHIB/Q08k3kJJkxoXi4C
M0QX5dJ6XOr3AUReXo3BiQXLQvA01qxt41F/JVQK8hGdKflumZPCApaN0jmiHBLf
rRFpfwlVE0lNRVoiS1yd72KFzNAUWQklTO3N+MmiVR1eNK5GzNi6KC8oPTi2PF5a
XylZKRvT2IjhpdFi297aqSEfaUI2csT4O1/5l0yyN9znn1Ps+ArlA59BcON3gZCk
uz4MXjWwqHCQddVSwWPAUXYO04Sj4T3kO0L3xu43Gs3QiPCKrLZ5netGo1ssztl/
6MGFjHZhR21pViJzudfGvEr6aQ7JmXVMuBcUK6k/wYbM4nT+2EiRcM7gUHoNS93z
5t0YCFH1UDwIgKTAyXn+lAzFhMEUWseUf5I+ud8mPP+7XNbnchi8vGp1Zli41JBE
Mbyz8A72Vjix2S1e+rU+nRRJdmR+uo53NdMmmtkv6CkrQ+V5cxw3qm5dbOHd4rOl
p7BEYt0IwN5O5UPwOOHsdeNmNfUrzVXZ92VISrj7+mCm5DzSWgQdA0dHwMmhGt5w
8JFCW+Qrn6MewxYcl8DqW62BrPor7tY2loP+0ywT24v2eTE2/pu07OQuMZxhSRhK
wzdLshCMzDmHJsRDq7VqSpxko2tPlmzxpTTAdtWgjowPgPKc10sIAYOfQdRT/f1T
OYASx1+7KjH6lOd2m27a5TWfhV6ofuvLf0c7EljAXnueYcEYtmOH/w2UqL03qx9n
SjKYTx29Yayl6HQLG14mFqxAY/g1UhEqKimDvWopnhseYPfkLd3TQ0f5cKv4xyp0
wHi28EJjMefKZx13qNbb+kNWjvOS34c4PhJ1xwqYh4pcMxlO+uOnmsRMKuEgKznW
nkyQGcTfF840rFspacGs6LN2QAGp2+5FRq1HvtKMIj4Y8wP3PzvrjLuSVsjHGj81
R5tGgg1UdjiOVxaugZYFR7D3ThoxaqJv/fTTzK6Ft+sTkRefnJZ00Y0KzlR/yGb0
TTZQTLRNu3FL+InmHiGikJl7fRXSLpDEmSm+4TBPczoHczBndF4iqdY5sAdX72t9
7piXBHRby4EQOJn+WVIlpmgj0gPZ2wSX0hqn/VXlpiy4000QY5tZx1ATPPd/aqWa
bom82kEAIgFezoS0rOG6tu7IC2tJi4C2A9T90KyXWFOWvVLQNnBrIl28wuPC0NUK
yLczKHFyv5mjXOB7TtO56U0XbdGB5+kUZe0Y5oYFNfcPEFa6G1hPk76A0D0bagAQ
NWUIb7qKl/nFOQJ9IpSrpOt/j1286vUisIrvYFMKkVr4Yp9O/X5rnaozxzT33vVF
c3fTpRLSsh5i8yRVaL7cwLacZtWglKCR/uvx7ef0f4qau3O+6mT46yefShmrwyXQ
OD9JGtKCBGKtIxHGCINr1XltmCneQqybiwUfALxDxwiWdYrt4gPWCTiqYSJvNrJG
YyybftkDhZEihTQ2oYjOfeAkZxorjziF7SZ/T/rjl7l0Vie/DIHlxss1gSMgkjvh
/gFSmzYq+91gVt2sDm9XkQuGOqek5bYw+ef1qSg6ADwVs3tweXqXuXVavWQHnj68
GHiSDyHcBHBCDfoMcYJWRy2qMaJcxyk0mjgLjlnn+DHAYwE0d9Njy7hjSGOLgyQR
b4/BKwNgsWS5RYgGXxi/pEDQdCiYWOzhJU9J1Bg0j/UDLLf0C2ZDcBfCLg1MXHQC
ZHs1VmOGJAkhdD04IE4Xb+ER466Q4y+eSvnWI4rZdLlogy39D2X7aFMDieFt9S/+
jhsDodBLmN5STOLMatLW+PrwIqeMgv9oSfkw4dJsUY9ZpvYYHA1J4UniT2Ly7dNv
xnqvoixJYYZI+rMXmuNTILB0aNQOgLbxOVHILvegKzlJBJoCCx3MHeaIwvWxnha1
sAQ1x2BZDzbiar37gMABPUVFMbsKkOQXklxNhlSCPCOpK9xNjZEagnn7UtUWLuIu
V9GzJ1xKipYQtBmVH26urZK54bvGDEPMliWtchQlrN29EDfHiYPkndVhGHE+XWUd
KQ5htC2fruKGzIX6GNEkBgTDbTv2aVjgPGe0A8HOUron1GIZYnPo/8jlumuLWgxW
86yQwWR227zKQA4vW0NkozWGa/8oQaoeiyj00yZA5w1VeanpYTlc4cl8rL6wICoz
AkoxuBh+K3dBmWoGfuD6wcL51daOmblBR6C74FeMTX/R/nTrj5R4fAPgdc4JTWZj
aGcsuSuzW7sLw05nTkfbJZQbeMmu9+ai67Af10sQGEvUn+BrxiwdoxzRZ5jhZObH
aBvgPcCTx1/rGNeCcmbc6nYfbxP+gBIilMaMS4ORAIh5QMQWEF6LDfxN3bMU6PbA
JHKkeqIlhvtfGxDwYE129wpKw6EqqoYsWAh3E3jRuk7faOIBqJRmRUgpLPHcakM0
Tfy59XMSMZgf/1X+kofdhS+mfNb0EGL8SUNayHgAjGHVVg0l/N+l+LCoLPfWQsP6
NHFUGoBVJoK2+y9hlPMuFctMNSqxpWnST/NU6NYq2ReA1K3LETcKxhznkF5xr9UK
cxaHV9B6m3d4YdpFlmGXB1PIU4iLCQSAGsL/bzcRjC8CghCXWLz3DwwhEGKFQkmu
3DTmkJN9iTphxIqQqmvvXDGivCgXXCamWBqmx0ACu087uiVtGT+CXkZdGevWnE+R
/6WaVGR+InsGXZUGLn3bQ1CXKOed94JzcGhc/k0nssQkBhGCM382vhc6UXcAHyDH
ED2DNQkdEYyJcx874OSIaBqoLIHNfzPy6dXELp9a+VR+QNYdKWNSjPHCn96SOznf
fKeUcsWGAbctPE1HLPmDD9RukQPxtL6g1YkJwMT2QyURnZFc0nvW/YKB6pZQc0CY
Wey+K0Fdqs1Co2rXabEHEv8S8eb3Xz2RT8AbQNSph/lxUrDjykrrvlk4JDUhlcd7
FCB8mLLEHztGGvYnk76M4JfHOt9NavJ6fRKS3tTkI8/r7HySgz1MGAczrDZGQhLj
h8XpNM/Zg8TSeXk409xqHne3vJRAlhqqkFKaql7qx1/yMORDh7tlZnPzstBsZBhj
KIkNlTkLjbd/07OM9PIyL57STwV2N4kiB/DxtTEfcihYq7bX4v2A3ucAWfItZC49
m7wECzlqPj1NPtgZ9fVg2EtygFy5o9Poya8bpklHpiJYdtwIrIJc1HShvTBfzemo
S6a3V4l1EN3OIlsV+RlfNYl5P9Vsu8jvp+ncVJiTDT66HKVJgWLHQscPcEYY3dId
yTSvfXHPOilbv//bSH/gRN25Mz/mEdKjqXO0AWQVZw/CkrKFtgjI6fszJvjYrEGZ
J6gSLVxbpe2Jo93tx0XWKICMUXPVwWj29pN61DH4Ivu/siMiZ0esBokrE324IH6u
qmklFq0ty7Vko9N5f28yK7KSZrsMfnpgYM9MNWPGuPMimxAyznDoouL1TFJSpIrc
XOz+0G3UnUjbirEWgbgjTHZBI92LY7kMPFnUO62rwvqjTf8AtYRK/vVsy8URgKZa
rGgCg1WmOqUxVMS9o/bjZA93mpiRJory+fmAFWuEZItHjLezMmdjsS5YPzV6eqAm
H0+k35vXjPAlgH2ypJl6fUEA0JZ9pV7ilTKZaRbSpAaBHInvYrOj6+VBYy2+ivIK
bI85CodoCdMUpwuz+8R4KWOcpqPnAxAkSuazUSIYPIgqXEWq4SHatAF+qhKpdW7o
seuWacNvfGwspuagsERh6SscQI6bkN3GushksFBbYtrnCKQYUTNfBXvPZ4oAfhqD
3E3MmQI0jjbARBnpqhqf1X41AZ6KhNzXadAmFj3i4XMkyWmsploJqv1fkliJgtpG
sRbpZ9jV71Drrwwf155YiHE/DEvefDR3bNZt0zM2DNQXjEziCsqxilreuJ7g3cqA
hmnDvym3rk2zzWgFPNwKgLntNxR4M2eyZ2vGTaqR8DWzPpyPWAMlSOJaeJg0Qkgp
HF5Q4gwvQwC7RO3rTOS+kl6YTxgudslJoPK57cXj9LRyDIVlD3bVE+9y5wukXX/w
TdySakPEMobG5ZfJHuLNkHWi6KF2XbDcXZoQUt1hBrXkxKDwXLHp3R29zoMQU/sK
ekyetrKeKf2rUA3X+l61Sp6SLZE/OIz5j39JFw620ch3aUlQ7u8hSiUcHPFKqC/M
vSxgMpH2FQDO1snV6m4bU3Lk0h07GvzlQHHcK1xICxzbY7cteccfunMCrD92KeGG
+cQWirOqGx+rlEWEoo21WM0jJryEOjMZYzcO1CaNID49NxALCyK8eGP9CJQLHi+I
1aPgCSr5To07MIhlAt4fJ+hjPYBqfhD/edQHPBzrgGrqo+8GAbzEG8yP9E/OeNsP
+DUqNDMSk+J/RYaJI4PQJAsfzPKAYDjVK/3u0Xyd/q+pkNtLb2OGfMnjy9pa62r+
ILnif1SYagMD0WNh3awYwF9EdvK2b56sC+DvmcE4qfxT0v6YErGsqPYmV+1IYM2B
p0DDozx1g4/jRYnWjp0iXp4L10VwODGaGXzLyWIIk1vkZct8f5ySOmNjMujz+U06
AnhV/XwdjRXpy/vbAQLO6mGgQv/NmQuRsXtG9nUwp3uTDdmpLFqrFPbmu8Mf73RC
8MFq7Blv2oLTjSFYN/vkyB7n8CG3hPPgavkXkhXsgSmMXpBPeHluKV8BU1AOyF7O
AuqPuGto5d/LWvv8lT3WtS0oyYCa2B4KYJbzkp6NnimJscccmW3GC6IKjZnVhBwI
DS9F4UJ/dtbn89ea8JJfU4ETbKKO3OEHOfWWh9bZwSjdd6FTeoet/WVWsg6fJAcq
nk/pBQX9nNdr5Q7i/cVI+pNUzsGTDTA8K+G/riItSMo/maeVdPwUN+Q8mXuyx+h3
wtNSuLHqpaFQbWaw+QqdA57Ix/ybxm8dmppnYkhBuIZLjcY1QqK5N4nzMNs0vUlh
XHndVq+Gz9nLqAsaqIAqFdNRmO+2w99odwrbNP2lfiPvQbqiLqNauwlcPiXTTbtg
QMOpzgPAuOBLKC7EISwNhGbCuH4CGa2om5XFo4dawm6FrTBh47VrgyNPPnrXvJGA
cHHWpPfigz95RzTsc1IvpXW+uoHENBfMhaE5RYBC32OiR6RNz58LaMxKE5w07TbK
vfy9dNqrO2Ed/moM/M/OiRtdkTDozrC/lZwCQ9en2T9beOB8gQFV/ORrJK0MJRPY
hOSeuZghYw6v6agiRUCX8sv3C7mj7QUp0glGDQSPHUHq8ud0YefoWiHVxxmgo4jL
ocrZcDG5ESHQwB1Z2aCCNmnu1eUy8ZFABxehyGK1ZxnOHyz4nh2JbO9lcwsDGTC2
f1yKXfuEKpEQ8e1N/2DyPd5cqhcP5WCU2VW1ky6kZdU/RvDPC/wYJba4/qfr1K2b
WQL1P1S63ZyOqvSg82UY4r9+X700SNR01zuOT3qEHE0esMP6ewMUXRYJs+MS+nk5
TUuL8YVSBJatpCTBGYO9eO2mJKdWldnJgHuV8qzgkKkQXw9S84V9iTGnCOI5wuIq
NxPYTyiJ1+UK6LFhjq5aRQkqAAp4POVpsL0mLtqqMewBydMqaAqggb6+DE3WgWkm
82jmwPIayKlwbe0/TmXZUfzvyz4bI/eeR+0NhI/Zm3jOPSTtiwIp+UpHpN+9JtHP
XPTD+Mx4Skjx61hYFU7fphU2AG5VM8BryznspbnB8MvbWAaTa81/3T2+XTu+AugJ
xNgGjpAjCJomZOLECOtM+JHvdSZQa79LzKItAcX3EDKWJpZp6Zzh04DTlgN/J6AJ
kUyqtPBSp1VbzPBibr+YKVfGqoQE81GWLUCx88sxieIrumEcol/h0F07WFGORucZ
VoPZfPtXIpP8WNAbZqruQCdlajymR7oL1mVEP5OwY8zV+XQwrnfzVHKwLeY58Lf8
9W5/iS7VMmt+utZZaxYN4jerB4quKDfLLTgpeSS39DgxpsET3Ldw+PplQHsFbrZo
znf8rHHbTPLbmj8bs/nrCPb1G6ftzBgYWphWY2OKlRaco9ql7pGHtD1x7uo6s/T0
Qa6r687IfPsrXgG0hK+MQ5+bzXaqUYm4v8NqgyjQV7HyuqjVzmD6kr8aAsbPbFP+
+rVLhR4pjBQcCQWBrXcTSplB14vlwYKjvGyWhdfDMuLlCTJAODrtg74nbkC9L7vu
1hYyUJVzbuVKqOxapGGC+WdH1w5+PgmVUmTm+CpazNDpIjxtIe0WRbF2kuzIqUez
Z92j/sKTh4YR1T5ByDJ+MHVzlqUwfN4rfaPTz9afGYzKjaFosX47Kp3p04w8vY/K
01VziB+xGlQCQIDSb2qngKIiC+NBR6evehqm0BOT2B3fSmMTsCVEEhkA6PN7xX8a
noHrd2t5rnThhIHbHyLDTNDG63tSKv+zCAvActcGmUf4ulP4xCVLO8/hMAY/x/dY
TCeq5U6SnMi/T267J0cUCo3SPGxDuxCCc1uCmYnJixIJdA7Qa3lLoTfH1YAhlh07
R+ViT0NxjlaVqrmce36Xbl2zpdVG2RQ15snMWBHlnIZxxAKYeXv9WzlPG0PuwMnz
MxBAFtYJQ78ZkQmskvcn3KOLx5/15TmcE4+5y5prcivEbJlgAOfoyUVV/yxN8iGB
zpV7JRTQB4smcCqVLHLNC2RsxkbXKDeQaIX6Olgi+3nl0Kr9KpQSn44i8121oxjS
wUlzOoMm+wvQ36uC0q8WvXxlndcXZrudC46TKvFfMfThZhVKxWmJcxFlkcMv/gqn
Bi/CUBHPaME34+MUTxov6bqXcE3kBjXJwlkkFKV+5O7ty0KWSklrkzBRdmw3YjV7
dhs3rtuqNT2fGiduIRIRwsdmYf+E5dXnQoOtUsd4bF6/ufL6Nh2iIYWFMZoq97RQ
1zJYrRCZrgWQrqO+Tkt1voglKizhRogBUYMYnTxO1c7dfkj0Dkth9kbkftG7I5Cm
qF6uK8xgtUDi7CI9FtEk7TDb9P7w2M/1GabSFe5Bo8tNbhIPXSCsjCWHQq5w46y6
2VaTNBQ6BZHScUqTugl4HOF4sudmPTIcLG5wJvAjOG0kIFg91TAqJBVcf6hdPlbj
TrTK1J0HF2WaZdt5YpE7smVJwd1dZdN7+7TyhC6IlW5HXtbzyJjXUxoAoNS0GziH
KqW4W+SaOnQ6i4c39d8mFfs+hz22Dtb4ZwWt9aOwbeIaNzfQ9zTX7cwUUqhKSIlq
mOix0f+Tu64kfEtHxqhS4sRpU5V7JOEOVCf0oB4VDYrs1L7vXov6DprCGEjq+Pzd
tnczEBao17Y9/ZtW5H8PexW0/faXc1F8TFBkPdmBW1mW/tsPrtS+vpD+/abbLRYs
bGU86lcLTO7GsZ/YOtlpWxLaA6K7lf5GysdHOIeLZ3JfjzrjYDYGesylro+JSrGG
VvV1jfmWmUbU2XZt3NduLKzRgrQWI1Cd0vbUeuLt6k8ovIA0rf9HcEStSenyeS6r
GmtnG8X5y6O/ZtlDlJz8mJf+3DM5uDUm9WihhURa+qojwWlbQz6Nqkyw+SHyr4zN
Q1UD3vD73tdAuzHwQyRkzuBT40deXad16jPDnbb72hBDf8b66TiiOxC6b2FOUreA
jElYO6nbNGWDN90ieYFVhoShI9b/ntnVt1elazTI2A20duUO1B2d7lZyCSBwifzp
wLqaR/pbtnXREqTk/Dp2GfdqcBeqbkzBw4Oko3sUooE4jkyMXtFMmGvS6vPInXXo
q82CFG5iGkWmMuHb6CjTKh4D+UH+rfxUMb/MenoaMIFPfLta4DjADSQclGA2Tsfa
X3KHu2Od45PFTLiMpmXRNgmnL3JQiUAVIV5EVOxtML+T+1hUYuEi8lTguaGZDK2V
HvMZ1qZA5DTxB5XYq882Af022WOWCr6A5yj7G0eBAfQfSY5gSSFv1XcvCNPc0AAH
wEIidhadoC26t7rFcNlcyodV6w/9Iruc7+wHnuaW/MFS4BSJH19QZfDuJqmdfY51
w60xQTQINaU1jL+qxLUuLKfw1+sIBJHmURej5pmtq/yODxQwlv5WaN+r9NPXQRDf
U4n8BK8jv1M8uhUNdZtKSWfVJh1ULWFP6PvemS+vm1aGEKQ/m2Trh41ZS0qL28Ys
PA8cqfAn7K/gSN7UopM1ET2/c1xxpEIgtw1GvV60kxDt2+VeUfIxNrzYudZZIraG
rL9R6Y7G3yBRFDGg+0B4lKCCfiihtEkHzmt2zq92TcPUzWPxD8pU0sebcFJIwhkv
HrtvoSynz5230DjdVrmFdqujzKO88VpZGInLrGJy5B0VVRNvQsE7asYqFIO7DAyO
E9pIpLOfBi/KSeWmFE0onJsLYOqzQX2KztcIDSE8v33MQpAmr59yzMzCri2RkVSw
AtOPlbPQ+vTBy0sDX1aLeu8vZG8QM65sj8C5uA79gkM2ithAC45VBQikW/N/ZOYZ
S4UE1Vn9j0cRyZ72ln/uvXr5L5+WZJhx9FENmdSnb6J5lcIm4DZajpJ4pDtKHecq
P3jiwMF4IWOzcy3X80U1OaTBL438tbM9Pw4hzLBd6Bx0ygFkFGQx21Ywxr+OMSIj
fG+oFUxck3eDoVUsHhargfu5rb4Ar6d3bXBM2f2fnyPsmccw2p33iXydiV8rIlNW
T325p5C1zxkb/tRXxu9jJR1GnzwTgPHQ/r4QpFI2EpHgWfdm0664jZnmIHH4QAV1
nXhQSpHiH3FQd3gslF08YZWtsNRYvgQInFisine7JVj50GKj2SrVqX0tUFl7KN7P
526A55r6TeenUm8LdOHrK3XlybkA1H/1LymqqWQl9PruM+P/vb3N4o/a++wCk551
95bGkipJ7zBktOgrphCksk7M3RqwRDqP4LWSYXYIE9M/SMixCBeeBpwdOrINmBAT
Q/w3AZfoaphjTC0zs4JzMd3W2c0ujtF4/MDxkTWOhdtTr8w8emnQDmVUjbFFzBGr
jYti3Rg1hc3Bm7kkRYubsK89d/5kYlz+SjeMNZCtKm9dwj+tc1P4197A2TsBOHey
iV9GgCfzcUWIfEIG9NqZrxSxFhp7dW+mMWTVzc9waoOuGbcYnBKiKYZEBOXezYQm
U2H9kGn+i3Txse8B7Wfq+wXjGjUlZ3xZJgtjO1xX6Zp5Tmfd4hiAaMY99dtGgCn9
4Tig7aiaY9VLNXPuDlz4Rpmmj7RqIegd8tH1jqSQMO29MB+WnaYRoRKdarV6yKRo
NgX3Md95mn638InuAG1maKQy3FuGcPKk/DweMHgNaebx9Q6mgCxAOprUKOKm1AWT
EFmKk5rCGNJqURfqvOAkwOruLJvbw7XWrCnVHp3ZOMuzXlsvQ7sa2ff7iQZyRZYd
hxIbvlanhR3hN12lYx+VUzGzujT/D8wCZbubwYbLRwBTHnJxhaImnk8QZDXErP0W
OsQB8HKExspIFwCL7d2sZnyFtjpjHtfqX+DMPVjhKKhvrUDlUgUPWfq69rxHJNCc
YsZ2a9qPDvwrc9XOm1YcPkZvRACgRslEfcssKan4X8X8O6PpdRTWSuYvTM5MD56u
aIp8WZ1no4vszEKDKC+NpbCvzKiEu5FUMJvUX819/tu4iO87rd0tESnAUbr0sknc
ZDFbD/TvnhVi4PaF3YMxaW9ZO+QxujTsF7V9ktvDpc65e8t1QAaBCIRxdBrfGpBk
ukRjbo0qKvA6ckzw9Bp+XiX36BUvjL1Nkbrqc7DiN44FaDgAlGhgXTDe0k3JtkPu
HyQoLIAPRngaQPUzpo3E64HA25eSvIxRO2j1RjEatODVyRUUu8hQ43u0Uko+g78g
XBkXdxNKeAeNF0rNxnlRAqhWBHoWcKl9o47UhJiB0JcrUfK1K4frPyWg8hH2H5xh
ljCow3QA8kj815UlU0b3krInrwH1Z04ictD1/vE9FzsehI8pZ5Dw84j3P+0E3eO9
RiEnm2YRoWk1UvGBZCizaGNYP4HLTKN6e2TRZq1AvhSvTG5oEVUSrVDsGp40TaON
rfs5fxQuXQRkfkB80Ow4HCkzaW1ksdiz/KbefRE6+dOTakUowpidurOFfohGtF9G
+CDlZWKkAu0cnfdZziOnNdAYfvq+qMamNq4IcmrJQzj9NvgoZIuwazBNs5QN3Bep
jeVB7iGp/b8kLElImSL+ccE8G9XmWbwFm1f0d9c2fbxq2HWLmOEK5VTsy7+FcXqD
soxzGX4EzdZf9TDKJzGiOcFc7mJlo6XIHNOOkaL6Es1nrNcRS3q5oJLmdUEWdvgi
YRtMzNmtawV/ECxl/koyeRPTrNuOfGihmizJSvjSfWmwX5+X8x0+D3hN31YR6htx
3T1PQNNO2uHjsz4pf85y9by/KwwU0Qd+ZWg6fvTB9NEtLw9Qv/qHIlhAKB2vf+nP
qpmmSoigiWZe3SuewEjSxcbheobYYMLVDRgrj3dz3I6RdP7kQYN/W+cv7XSkWhrt
j8EprR2GGxRmdSFA2s+H0kSNfpNUFYTxXWNmqkFDtVKLw30UgtCQa/o0VWpBMSR5
lD6gzQRnJFIMBq68ozVd/a8tm7FEw1lZjl1lbBfmAgpFbt3xByCPocLwjbxPpAT1
1PO1tGESWgHTJ5WhACXAIOTF3Box4dQck6tTUVPlEZMC8uc8FpiyaPx0oHIOP071
mmekKm3X0RErceeM1MLrlx09PWK5F0jweiL78yFnQ0UGQbTzgFVrog8lYK51OHN/
o2N/pWUSbNsIt5Fegtp4gmDqWosMh6b0g0rtGwHnmlAsC5y+Y+VZnt7oNQTCpInz
MgR5ZcFqNcwG5tZoRRjJ1tMNvz98fMUO5xyVF7qfMEivbAQBzVV/JP7+81EV8eZM
ZACxK1IW1WfZEpYu0owbJg/0gf/5JdcSpQIV8nlTv3D1Rg7ljdxw8H2JslDnUNBd
rU60WzowSK3knwhORU4cYCiUDCGXmVeqpwijfds3lcCwOGyNVjcKEn0jexKowSy4
WryWrN05N2AW9V3frSvenHX9I/oicvlSFD368xFDXFsNWC2OwAhJd4h8EgbMfFip
4RHwlDVvBcoi1bUYBL4G/0lsifZql3zOQH5Y4GGkHTuL4lybizcVMjndNzBiJuWO
fWPxMO6EfS54HBEYCnOri/utDI5lAL86wx5M8o5r/vQPQe6PAXJ3z0Y/abeQxATY
65rsUb1nUcamJBNT63sEfBNZOK9Rg3SsGqmUSyf0cKIMqR8ikCqZo6HXJSJLh7aA
cBoyU1oOn7gNSCK35KF1cMBEtzQWPurww9/gYApnQ0idrZ/89cYhN6nPOJCLkcnJ
tjYrVqs3ap56s/KlbFt9PcIqbRKDTOGdtGEDMARkW0Di3H65fOKf/Jr274/BgGsQ
TIdNPaAbUKrTMW/C17C7mB8etgLmjsi3Q8/FLYfoDalUwrpg9B7mSnVUHjh7uLlx
p4f8RegzhFBjouMKDecu85FSZ8L2LggvP5ZrM/NvmKvo7zXUJo+f/YyVWGw+Ecfn
9ZIQDo7MO+4g2RMhA+TX94bMBfPGHRnXTJx0W+19eRmKNCiliJ7sGwS6JZ3mKmNA
+rVVGTH/Nkbgjt40AGk7bmABCFsOKlZBcYXmXhqMf3oSTR5MJTDjrLA294VWMiV4
jrNBIROxIbM95zxHu/Q0E9SHrThyc0+CG6uZttZuB3alIgR0zTsfoMnuE4h9D5+r
uF1NpVkFbhxtmPET3ncVx+O3SCG5VhOzkdrk1BPW3iZ7dr2i25B6Qf7FM2eiQ+n9
/z7Mugdq3cgbfP/VIucaJunvHNYNj33C1smK/iOhVE0yASPAMN5rmJpe/z5GTHCw
2c22sYXAz3xzqDCHOc3HGbwhDQaO1ZSh0L1xxAZMHn0Pbwox7+g4D5lt0W/B+m2d
fwsAiKEpbrOhycNgD1gAC7rXk8Gn460U8mhOll0s7ypsE8+ZCp46zl4giG5bfGrl
BXNI+TBcvmRKghGLfi3HMLy+B4PRRr7wHPuO5ixMeK6MRpDvAQ/OQsZ/U1MNyd92
pPvXgljDTcqLG5ulVXG/2aLqW7J8NF8VOMzfFwROhg6vKtFRLe5cMHsxygjaKvFP
HPXfCGQUtgHJE7phqRO9bq5+SC6A94y+If87EOOiSd2R0VLpa1asjod91pkv8zyZ
g8ODH61eL7wnuafFN7LqyruvuUdTnjCLh83NR9wUA9YgeDAM5uaJLpp7bPkjxvwA
9x3yGsnftjPsvJoBRSLnZ/l9vIgMeTnO/a0y0Y7lgTlkS1dZIJcVwMzAuinrRHQj
aZuXAf7p37FlQ8PMIDh34XvVm+Jzf6+8uoW2qgmaZjgfhKSjuhjiyvDchF/WBOva
9dqGvQdqGqgAPZbkbaKx8qh7nDo4SEgiLJtYEsuXVr+cBHutpCvnDaoUjhNJqAT3
mbVNni8mjv4nwzouCZcOF09tA83G1qa6ZawrAGuhC3hdorOtlMGmPhKAi6+KxOb/
Jl2mLK+GYswiuNg76gTQam9zdv9Ufhp5mhjBPPzUtG9itbvBqttxVf4M0b6xgSvS
qBb11ad8lhgw2GLGmf3dtmh8uggBO44svaCnu7Sml0zEuHsfbRyFmdtJxf5XkV/g
tgYsYT8fZiP42+vzWnDupZ1cthgnmtqFSTryataA5W3cepZmd1p7IyKIr1wWXQuY
ggT5elAYnK1qI697MlP7OB+ctG9HmK2mnTawIBQ/2QtVkIB9Slof/Tygr1yoRO3f
clp2gU80pi5DwnMYoTwoh2k69dAGcu+140eV4Y5kBhmfeOPpuLaBLpvtet/XiBaZ
UwEBmbiLToxjke4ZwWKztO0uBQu1lhDpIW2PL8ympfe4hzrO1XjTS9nqXhvvOYM9
UpgYJh09U23q55bIKt8toC94mYn3vwTnY89W5wVfmzNdMaah7kA5WeEZSKUcJbIC
zY9kktVaQsnJ3h5oRlUV+eRZVB5DH0L6OV84ufo2xvqUYcJTHmZJKIpsXVUrrTLF
e1dSDBcWwm+Lv3uAf4FordPbLB/yS+/NFHN8Lr3aWKEHLU661jgMyt//DT0CjAoo
IOPp6Gp8x2UoIyd9FXj9D1lea8SQ6QKKR3jfmKyHlyqa7KFNJu3zImxcbx2tTkAr
4EthRJXPZzjRR9YzDYpTLT7unfX4knZFU8tccXVoOzmfPMCYK2WGfrl0CzGsGkpr
tU4DXvdZX0Qm7N689tZJsphfXdicno8+G67p/WnOO3RGLykyfb5U9p2/SccUrmYb
nppfdQyh6pc5+V16bbvLFa6h53QTr+qaof223sijSDRwBrZvLP3asOsL+zni98Xi
5tAfTiwyFST5My5cYz3IyUFaYQd2c71XeEH7NnJV2IZUeF/eb6OjTDlmH16kyuW1
0ii76c3Svh6jJJ0iysNR1nUPf2WEPWwKY9SNmcvpIobQTCY0PIh9LIxf6eNzhrsY
3vjJr/uR3GPviNqwAQJhco2HCGg99XbiyzezJrR1cEVESqM5Qsf/9tRUyqy9gpxt
LQKo+bPt20wOv8yC4LZEMS87/tdVe1z1P6EO6VkVQwyw9uArn2IEQ9zulOhNrrOk
5+WBKAhnjgqIXq1DTr+lccmCgaIustiouutXJl88W4gCPEnXpBey+BuQ96p2+f2W
713EMqMRnY/Ssu4WYyY4IdRi9XhQZtVVUiU4tc540YsRmA6EqRdkMZUlRZuNmZWI
4NsmfggPSkkquzYxcZR678QwgE+CR7LCScN/Q4SNBXVXXw511qI4H1o5v5IrJjSC
NclKACvNG6BLLQdk3D1mULTXfTqYH/GaNSoziUTMwKXPDJCrdaUPaCvu5o19e8Rw
jZ3h4q6ONP9DM486IC86Nn8OMiAdsHe/8frLUuwbSAPJBs0GpQDx6deoZ9yjSg1t
FcEl6wGQE7/vQln0FTC+Gc6eO3cM/hTPO1fQjGZDReJb6oJDcXONu9gAmsgsIWyr
E9LMG4Z5IkY0n5A56eNT5GlbefHCvvDcQt2M5R/Qn6iAO0LQiqKcfbbeE4CYDnu/
hJd0cqGYUKTowuginS9N3U8PReVIcRxH5Sqolm0DVl6ZiGMRkvkI4ZfcxU4RI+cE
FOxdOy5YvIfgfkN4x5PqAYpHJqUrPtPtGK4Y36SfioihCr+QKFPoi2Cn4RA9Q85q
0QrYuU4Ly+ExkPOm/TmuGg1NYqgcsfC3L+Iqnedyk8HBNlFL3k4bJ7+/WxWesuMr
kPrsUredfUo91TqISOBgouQ1Q2teRjPU8y4sNrci3ca1BC3sBUr1wja5G3a3iN43
UP37AeVBC6HGGYtcSxhg+gPJDbMnPErDXNVrSZB3Is3ZoWlFHy0PMR/Sz8ZZAx1/
SLhyiBP7o3yNFkqysnR1182DtSy9U1rpf8tL1UatJCA3VdFX7GAcGndNNpSTsBt0
PdC39fBHai3nNiPqMgGtXkhXsr144DRLVlLiSmW32lxGgj2mCHBlLWIyAxoHqDh6
OXJRMo/MfqwNgF8dfhijMyWXF3whnvyVAnVyVeiNg22p8+Lz+v4iyjVon9g0iom6
wgE9V/BpmLweeq4wRmrdAV4fLZt2/khre3zEYboMqLvR6jgbY3NVoBJI8lnzwc/a
JBpWsDaWp3EpT24Uj2+4WyHnKx3/jOkFVV847YHS+c4cPvDYI6oaUDctDwAp873b
UP+LpqbiAed+p3jEY5lAzGsp9UQH7J+oePqtXo2+eJ7HqiCi/yzp9T0Xap08MxGL
cp2r2sanyVKleNZ1bLi1xJyw7aT1jDL/LGKqVALV9imK0KuhRPRqW/8ZNGd7ZMre
YGklKK/FT4kZCa6VxACHQuZxU29YOSGqEviONuZtJmmezdEdSu1WCMau/acdZsYB
fDom3Yg51mfKMoB4Yud5okNdniXoFnuCj37i81y0/otbdOmUViMt5N7e6W/bwA8i
NbATe5GeIm93KP860Xnwbb5Oy1Q5oR4+0wpMVLUDQz+0zWEh3veyQhgxrOHw4F7c
/iezI8daACjkGUJMdWCq06O0QW6POzsKDzzWU7cZBn6dJmAso4HvGQhHIuoTBG/e
5vdfg2NS0dn9KY5Qj9nafOooN3m13MPP/LZ5liBMT8ZXFCQjafgC2I5RRHGp3d2T
UP0lmdFzH7pJ+h3NXWzaazZEQ1w9J/I1YQqQb1Vc6JfN9CaELZLITs7bRReatUw6
Ysw6nDccT4fP7pfUfeHxOiae/z5Qxa1ckSCnnXKEMKfFhVhIPo1v/gGyljhHPpdb
HFSSJ7vNY1BpXmbkDRhMXc88GbgwN6f6Dt3Ko+gsMHGjVOtY9iajGtJZjrZ9SEbu
B0tRLp9gfwOYEZI9UXTHwrpo6XX9xlPlWlChRqlo8wRHgf4wWNrCC+5EwmSOnfeD
44P/LwBqwDIf9NqIUXX0KMvZ9atbnJWUxAveUCVYzfpux8jGImnVDtSMvEsMyY2U
B0YY1eeq42s/cpJYNHIGYXq45dOocF51epOapqtT6W6Kletag9VgM1tqaDbd/yLx
YC3DKKdkEFwKBjrmxY2Ay2+NNpzwx+nawEuHhqlVgF0s6pCr4P0mMNlg/a5ndZJP
VUC//MQGM4E87ZSS9ujwA4Lu3cUQw26qmL4WkSiC0zZxwUdliNtvH/M5hFFwx4U3
hZAh4T3bEx0WatwhrtIeeEqVYzX+Uoi2vGRwMY29UAXDi9yovB41pEBRxHFfq2M0
uYWw37lAMwk0qOKgYGdIcIJUkTbkJc6tfHB2Oj5gQM1JUlqTSViZJJyQAh2Cbb1W
GgSwWEV/pajrCX6DXX+Hel85Pjuzq+Mh0i9TnwUq/P9mO2YGWWhEh1dFtMAMebEm
xgGzflacTw0yHrmeuOfDpv8oy3LRXIpOPuSRrUAfAIkUrotCy5lV19yVtT2akRvc
EuOSCTc5TWYXwNtanhhtMjx6K1Bxcp7Ep40JeI9Mocdc1iPZH8URa37QwAwIdGn0
X0BMRQ5+mm/gHQdVQQtX4CE+aB3AD6VRUhdwcoWiHg7D144R0jrSE9HZGGdxNOqB
13NwtZKtl4GBfOS0SuVnjlpNK5/JFKA7TQCkdA4r/rwYhqYATkFbGnQO962CCPCd
T2gH7A70NPNOicZmk7najckuO/gWToQ7/fbCrm5nC7q1BAQfKh/pG3YWNPgDIIdw
3FDiLp/Tp0Zuhvc7+JyYmFglmfLjklGggHobKjQn0el40BLBxPGZ1p81lMpdU7Tz
UjPFieiOj/IfAwE8Wz4iUk/aL9n96ISXidGp8TWX0y7UJEv1Vz+yol6ttV0IOpKG
l++N34jxQZ8XfDm4wnqFxZui5dq4QCwiYOY+ZI+ZZYt8nEAFxUEGJVxeWH0/j9ho
XeuBgLPwarqXHbItPMq85oVhLCT9xaBXDM/m+gOKUtHJgOj3AVd7IOfcU9NRt0NN
zQBk498Bhq45MdFnerSt72/O5hOFiryjP+6nMbuqU+nZoqRm6K9dcnF3WiGE+vhb
I/lyyiubD0xYWte9Z3rNOS1GEKlRY+uLUFbFvTJm66sPEFkf+vp2m0QsoYEkObXm
TqN7GFTn/F7kaLz4ZffAP5d2SQtzd+d/6nhVIKhz+YZERG/6ZJ5LTZLB3ihGi0f2
k9TjDKjedo3mbpdVPCvnGJ2qMUJu+7wMbeVIBinObLn+Iuw/wLcJBz44ulmEf3V8
3BIXghZX6SDOiCqr0JF4THD3zxkkDyxsB1S7XxZ39J3PPvsFPN0zxVGkL4ZwJjmg
/jBgJooxW9AVvGd/p97PHycuRyJ9P+lYShCdok8/mjv8NNFawfO9NSccU7VWTNfY
vHxaJ2Zwrb0SyTlhPwVfa5YwsVjpnckMrQCSIBqIwrDo/y5Nwh00Icl9/aRG2Ruw
BmlCNj+iJR+JL/RlCTFkyNeSnlcgrQU8ruRnX52lKjogY7+WC+Nd6ckxNoNd36Nu
qMB/rB1fTVPA/qSrbHTyCN7cg7raH6Jg52341R9Ll1NDxo7yC577r0sR6p5QocJW
abGVYqwNpbhW0XDHs5SWMihqjwz4em+ywh//48e4nNGUB38UkC7s1pzpC3pKRW14
H+mwgZJHd8jbJatcdW64fkLMfhhoOYXIiUCY7KjFP4BVSwAkIyxop3jPFirxGPpK
VxnWq0kQqAbp06re3EpPLcjkE7jDFLWaWs94hX2yGXVxTAU6eZsCg96r23nQ1D+Z
F+RmMIsGCVO0fGQ8HLun6SUCa+roSCqZgAxWMueWQ0YRcRGsfc7v1A+kAeN1gQWW
S7VepfAbBNR1S8Jg2+5rzslfZpW/+aSzQZeIu6dQkc7PFhmTqoyttoAapFMGiRKC
lIawQPeTW3R2gpdqSevBUno9MSI/FxGxnoN7iCgjaB09s3xeeMqULIr7CyN2mk2I
NYIvw0DIzBgyk9TfH/9lmHVpdlMEye7BMlcct0ISeo1M5a28ZcxVwQll6knDhAen
V60HdNeRCXOm+liD4AyfSoucR7eeDe+1tw+MrqbQpqUxKpLnbjCvWJUxFnZ/5d2h
JZWo9p+cV1q5P34B0oov59WUWfSzuopnMJJjeInJhClEQ+SvaY+4W5uFk8s5cIwH
/HyBCVNNAYXX7Z/4unpRLsC6vvv1/D7GV9PbgscvtiUqozusQfPooARvVLE3pKar
RO7nyrBmiRs3iv8Yg1PH9kYW+9R3UhkRpCyBcDdUpTu9dhY/CoKDi2T0sydyM5bq
LfYGeHPOMKCN8UKdcEeaAsKbQlOOoE7x/62oFrgfKDIiMzhrYRzPWFu+55Ln6IeH
gQr5YLGnugfGJvfRBEJyhCJ15gv7m5Zea1tD/gvWBRP4gY1hGrEGdL6OcGBTlqZ2
JH9gjcqG+DZssJZBTFR/q+7EDbzz7RWZTewMAsx0NJ0F9Q88fGaF4n8ei2FVLfGP
Yt/o2+apKRoA78BDziQDMcHgqgr6SzlL5q2LdouWZwqm+5hb5KEup29Anzt862Zz
8dlVb4MjELEQhkN5W5BiDEZs1wi5/yuFSK8xVv6MVjekPMUh7XdDddxDZT9WrXAF
BxropEWy2pNRoN3+iSMIqrRQa6HRPBuoGVB7T/JZbh8V1k6cLadwpKSZNtWIIK8K
guVf8ZWY0Z4t4TO5cjw73g/SFDR4Fa2BSQp4neO29zoY0SKep/9Cl2E6+NPjLtPb
Ec1Krf3hcA9UqqKjTsq08XJxLjewg2Y6scRjXBGGaRG+uGyl0d/Hsk8K1PksrkrZ
ZYFwJedc7XauzocTu2dXrW3EJddyU3jUIoEPVX9H9P6DFEpsFSzvebOh/EZaIN52
QUzUZLLp0snRrcfQQB7a4LBqcaA8twGWqAsmBsERospke58J6owK4gO2n9BCTTIl
kXcDHVAiLWL/rsJTSx5+6/Fy0FZcpTpqUjFcefBOlGnJoYmKXWZjfn1vtX+1uBwk
n/eViqM+evvxS2hOLVFTBHYmHtro5RafWug++Oen4STfXQ6ZQFZJJXkAr8WCZatK
RrS8+e00uAETRqesaFxDBMJXQ5iGhGtp//D4o3d+RWoDrTPb5kDaUfH1tLGceZqn
8z+UYIp1tEIJBPv3swXFnpAw7bXIgYtSk2lsEA6P1Heb26EkkvVBPL5apEHwZWLo
vFKuBalyp7d/FZR0LyLJ8lChQtx8FXK9qctGNds9OPxFakDBIAg4bkM4tZLb0E2b
Dv28Wb55T6TzUvJEgVfQqPzKduMnqcFAkus2yLmQBfti0P7I9w8iFXIhsKtm5Pxo
XgSRjpEmA4hMKl8EDQhcknI5ZVImA8JNopYLQPOQtixeBP2qnW6Owlu4zwSwl9+J
tMmbrK61ovdXksK7Cl6scyI/KisSsRoNBLhooL9sPrPirtMbAdp2SVj6aLFlBpWA
0Bpu6XdFTf5Lwx5uVWSb4eKTIYMbCPTdDss56w0dJKttU8SFG2g3DM4ZP3kVBqGe
/IazBCcBLmrfVHecThCNwrXvBz3pBMceILmne8F8LnwWClvE2LPj+wr6CY85CcQ+
Y8j1rCDl3TuBWSktgcEe1uBuA9xgk5kVzWcEPqcI+4zXk80LqlqVf3UAkuDrdykW
2omypLTlm2opSAroW87jgsbD9qr90hDf5xmdHOTaDOJUnNUBovI2ESv8EK3ss7bh
C48kxg6vf/jIeQVp9/PXUQOyGcmaKyIYX6LnEdxzfVCHVdX2Y2hroYpUfWgq2fQk
e4N93AvmGJb7UW4onbMvptH+ySmrvOBdS53mVXEv8yZG92rWXlZKcaXAbnFXAxBx
2d2J+LsIK8IyJxxkK8uNaOoZS0j8fEuvGe6dyVG5koS6dKDL3ZLqnSzVp5l3zHKZ
VtTjGwMdsueY6VnYqX4sZQdwW4u/rP458HW254GICJa7bvoB7rDBWmf9X36fzVXG
ytz2wAaF7yAzHFma8VT2cTRc+9ISGmANRK0KQxUii+nmsLCsYL6g7IEg9AQbFsuU
L4EcJGAWFa2GMxW+mvIYCaqaXBP84e3VCQ/J3viYJfyQP0S1sqLUEvQXs9fJ/l4R
pxbzggV5j1213FGQJ98PhYjwZdsJQdLiqHQEZiD3u7rhvVxRzdWb0AFh2PTnuKEP
ec4iZAFAGJ3ZcdDoFSlvE4CepzH00K+Qp/HKOYvyBMcX8/uOU2ZLOFNl81UEWUus
KcU84gl7VQxyHpmryvayDpwic/DnNdMN3NcYxv/x/DnpOyFgRtGtccLRVdP3wVml
uOSFu4t9ZqV9qkoRST+caHh2Z0JPebhi0fcwELUqyn9gYDXKpuAcRYY00KvcGDtE
D7ISGIZszqt7NaBdvJgZo6/dhjbYDePalM3kXkHjMQKCxV78XjL4kg8FCd5bhN2l
aQPOGMz/GLI/y6Z8EpAglsr3/6i0c5bv22P6u6TvqXC9l3ZU9sv/E7nyKspYHA3F
1GnvmS+SqgF4ZDkBirRT/VcMQs4fyLZXH0CAAbggE4MI9pHDLsCmR2F0y41Bjxwh
02mtG6nlZns4UXzuR3ZBHIyX/JiGHKeCbHMZnz4pJ/ndRVUIZ3ICmmHmjf8vyW/X
o2uMco9l++Gpflt0TvpzhMHNJablOKaOOWaZ5hdaUVix2VYY7ERxAU6tEGGF//mH
GQ6KGtTmggpzCtEBO55EMyGI9uG73ntY6kD31dUUm61zi5SDoeI6HN4BrRS0ec2Y
J6sEIjO3X30fuDDnXhWbfgr/2S3q7bshsUi4oSLe043vD0Xiylki4SY8M0rUPd/z
s7dOYXQ7hYno+jUzPLLCgX2vghxPlbku0UAIGK+wuDUziLY9pGEJJ1vsjdE6HGRZ
BJXA9xrHKnMYODhFNvPazXXeTvBtEmhn+944Ceb6qssxstSjveKHGaw0zEGMLDT2
KHbXeoAIk47c+sMuEhxHNyg9QR8aPb0+v5LgGNPPliXPDyKUuXrI69QmrYCeXgcl
9MLLsNcLCX6ruOCSPfYRTSyrcEqa4ev/66ezERL42h1vzL7i0m44XElAcGJ4td53
oj/1FgsDFYl2QrlNcX2XeOwoJNPIca2ODdvoIoW8a21PgQQPrNHwajoYouXu659J
KnsLA07YlQ1SfLoB0j1AvY9i8yVuIs/CloI2SlZsf6R9BAC8kKgZtwvrOzhNdyl4
dqBv5Kvb1WXp9pqHtxSv/XMOkX1b4DPaQqcLXGZD/MRpz725VQWz/K1jteNJmeGJ
0HTjqcxVGViDHs4z54FUXvWiwkRk+DeEke5s0ZAq4i/rwDKWwlt5lbHtzpSyblk7
+K4rZV+iSHyFX/WYqHIp1E4PWZjkuob3FQHBs3Pvx65P5Bv3gaXV2Mho2K+2TRc7
4JnGY+xRIfBjjsz7dPpLWAbot7476AihTNdmJ9AEr2Hrm6lSLdrC2vg9OhbtCZus
ihh0+kjlMBotApSWbVYtlpbRqU5rIGz6ZmZ8OzdKjihCC8MasTH5sUyf3RQAmL/6
SiBVT6X5iGsw+b7m6HwDvXL/RNkY9YLtkHumnCrP7uIQ4la7me7pp4KE18iMEK57
GY5dt7F0ot/1UBrAXlKI69IML8ocFuRRK+OQhB+IJSumrs7GocBWu7SSC1f4YFB7
2KfH4z3sheHrarjY9uy8VX3LgpOVQdNpNWpHyv4fPdvDlfz5F1V/q2SzA2FpxHuE
MMLmfMK1M3kBEtl35/DoOaAPcfyyTAmpNXBN4Ui3/78yPOtGQaTJ7uwSTTVKl4sP
6O2sUZ6umM5z9+y82+A+hkgAdbsiKazCWilKKVsIzPFNXwH0tDTbBwpCOwqVqXb7
KL32NfhbJ7NgomWAbL+01UnhZ8mfnAFiu0oUoQmsN5PUkU8Z4rI4kucqpoPms7FM
Fh9vWl6kBwX8FOHKc4HfGzBLt3hsgTVfRqr8yYV8c6nEMwRI92eSvvPnOOtGQQ55
SgSvwh1XT0AcF0EpP1WxBclt5qm8Ibw1Bm/A7j0tPZCpTj7OEqdVZg4wSmji9tY5
7KWroM/oZkoqHpCW04YHp3g+dc1QeC/8vpqlsx7ZZQ4naJtlQghzyvazRJeYPXZq
FzKYtn+vlOcs1lH0yo62bLdY6/r/75/jzW1FPTq3vrjF7pTbK5gIxiiQe9bGTW6g
Ipo5wGOL5TI+Gzt8m1OIxijXxfcRyqRVfUVyICwKmFtyiwbGle63tast8X36iCOB
8QnD+dVPNqaJHO4P9m11PKIGuVVgsY8kj09Gw9qMpCI9JtRbhsEKF8qfGiv0GUQO
7+VIurEhQjV70qXq15oRIQzaCTEGYImci96ztapnJAutABvfG1sNzgL4z4kPXaXv
O05WEm+u3IKBSnXByoZdVStH3k61PLwT9chUbHX+u6H2y2VIqJzDSx1pkbWYsMBU
VhI/IIUqJOsvXtO14hHAKUYV9WifJlLINzjnalNX/pxeXUlZjZfXpTCLmQJZd6Zc
D2wv44w0mOGXycRZ6o6IEl7k6GOV66iNv58eBeFCt0i6kNdwlvlwsKAacBeM9oij
ls4ZvYXh2wbTg+8T3IHqyiezOXaVG+VSScPAoIX/+oXEi5GHgg2M6Hvnr97R9Hvi
I0cQnql/MRwxVVrixdYGdgL+D8X4YMmCC/ochOgWV472qMewjKeOTfe1sYixnaGV
oOCmhAXgQhd5nAKjHLi65X2WnWgWOJQZYgJBWfv1lgahDRoRnFiVfhWsOzGbv/Ee
RkWO3a6JTuBgJz03xVghNuekZKxjNL+3EzSdh2APJSHoGB1C55dDfvccBiNg6WsB
utV+TZXtN85oiyG7Hda2DeCm3o8PG1FTxP7zcfQU+VJdEDl7udkYDCEV/zTV3pYd
OKhLJJhgX6L5a5ACIghapU3cQFxoqlxMS52VldpMGnXiAIUvrMikPbyPGUFpEQ94
AMldlW8ZBHcdBId5E+gOtabJq9+y4XFPAFxkGuz4DuCo4bNtFVZyrdjOwV9zz7BG
pjGagg9kT01cwUH1R7Kw52Ywo2oeM2S5N5Zc3gSJmmWzIX7LT44W+bYCDkNLbEWe
R7MtLLMykffw56YkDxAmLRWUlyVxjLUA808Ci7/nxv6abQ3nTC2UNU3Ny1fOwyB8
H5ZqJsevoyBP+FUxWJXfn6DIzFYI9bTBon7JjLziOhH3qe7hnLKeEG9Gq1XsDhyP
+MmCIo/5/QXMhdZFV+r7v83R+C9nYKw3MOO6TKsYLa3jUZUlsDFmVRS8RYvpOw3A
z/HOK92PTJeLYlT+aPOKstWruZXRzkXvNSqUEivW8wU3I7R28Ly7s1iLQ+uYEWx6
JsvBWz8uYB+T9jS2qKB++tSM4a+W0xJcLzaf9qYiTf3QDIzEJvHbdXuoVBAdR/Vq
C/Sqns4QjnCJhAfcca8ZRKVTfcjmRRLDHbCILF6xombyhw4huNkQI5zYsWBwJSEB
UHztbnoV9CLVIOziANG2ESaeU023J5ctJWc1NBWGwrkcbUxWnJS/1jtZW7hFYN35
spujN6n0pfZ1Kw0gbew1He3yBotxbzt2meXy2qBhIE4GpbbLOxzH2uaFsZ3iocFi
BPXCNA/pcncOB83qWHMXtggvwVGPDSfSn+KAz8DLwOP/T527rla/etIPlPq9vFAT
fHUjZnGgOcfPWAjb+l2r787e0OSGYLPsjllKeDLIJMxrzo7Mq6HUKfSCqzjmbNcr
yNrea5jqgz77aHmZVZ+Gg5fuMK76SucRmZVlQNOmGdbVrMnaBy0xhXAQoNHCFt23
vKkbd9c3g+M3f+B1eFcplaSjHVJNyjMoilxh3823uNSFNHamMNOjBUDqCmU0S20/
f/18dD17mwtHEGWB8dYmhG+0Qe3hPaf2bAHeve7nXVdgMfPioPJ5Fez4DFG3Yaru
tLq82y7HWFs2LWo2Q15IYSUcozKzaTWc76cPeLpMcSYutDx5aXzydNzSdzXF+dgn
ZQaAbvb20L7vPS+biocJqBTziRy1iZmtvauspXGPq1XTG8PlzBwwFo0LN0sjxofo
igKtWtO3R/Vp7Rrb0A0UajJ/QZkRUkJEixuzvonQLYT5YP+aLpftMnxGh39JotqT
6HgXtxwZZ4Z3DR19wATsDZ4TlneMOYgBk7Ny6sgqVVGfH5Bb7qCPHgIWQO2wm5sH
UR8uBoixetOuv5lNgUXPy7wz3LzUDo/WC0aeps6+rnkd5pyO853RNdrz8OcwemWh
alQRFWSL5cRCUM5n/kdSSbPKNtu0nRFuBbWVUhQrN6tXqoc+StqPFYRlBblnzuJ+
e8FCPro+TNNYuTDekVPeo8kIMKKasE5Dv3jsuZNf14NqBAdAbM2dr98NX5rg0HTB
PdBcVq7M3b6GkLx/DNL3p6Tp1BoJ1Cc3gtnNB6CG5KW5kA/F1qRTwtE3nT1NYEVk
HVN5iACYErel/IqpJicTDcC7dCdwd2NKYXMVEgwS4lrfKo6V7yVpexMw1h8NlIoW
XbK6Nc/Fd1tDoFKuH68SXJYSdfeQUXUuOWrs80RPYdKzK1kqZspSPVTDG/MBN4KY
lDASbndhJ7TBx+DilCutlra/ENkc1uwV5nWww4xyTGfuEqcMO0WEhB6gu80iMMII
PHOwij8zVbvghcELOk/akRPImI234JGoa9GDNz1F3yv13UqZ1JHQVR7IuoD0TrT6
Sjghc31ilPc9N51xqHm9ScXMJjCWrXQHfYtGKFSsov9yCSFXrMppSVWO/CpQ+RBI
RJ0LkyiEmOgiR255Jq+EuLPa8aVlsOSWl6HvoP80ZRh/BA7ND0iJcVstq/EoLZOg
3l16VuLBOUvVQf8Rplp/Glh6edm9sl/FERLhSy1YH0voj1jiMX1HVwP6bA1ZpAiL
2mShOYhwA2EGIlTEWUutIkIsRQNuIkXo74RmrIUKAeQy4v5Mh06yBowlN0YcJl30
BlOC2mb5FIbWOia4GQ7uOSd9yPH1CaXxyt8y4VxtnIaZVsG5kZjWOIhAHQaR4qNb
K50VPu8SRi3LhLHIhG5lJRJsEsfliuoJOOPf5aelONDemse6qYeZrn6+EgRi/MZI
usAA058o1OfgWOFLmIppCrPxZi4oX8UBtGTH6Ik5yw+ZDNrudLd+BnjYPPbN29vb
+S+CPGVs9Gv6chXQO77vdNzAZ9nvMLpsyuxzUDF5U6F2IAkqOBJOIr/925Mom5EJ
aV+rv3qSfV20dEWUG8xATvb/RyXgDL+7te+VNE5s+al2xCK/CToEUFuE1cF3MJoZ
pqK35m2vsW5cV1ptqUFeM4esZVEk05ksRWHAeSNFCrVZJVb/FeU2TM2+Ft1ZqNKV
zksxbogQIDzq/zuWPINrSsmBfdJuljstPaDt4o42VQXWO3m4flHgt2gC/dZTwowE
bRXhYjBqFJS0ueOW2sJy4tw+Z/wMZI5jo8g7QjYm3F1iKp35hgpH7Sn+VAV2Rw3c
gTBsgHiNpRRUXjOksTjWbaOH4K/12OzWkRpZy3FBP68xcuzwo7o/BFDQd7mpjLKX
Asfw1gC7S3Si6to4TkbxISpUkpMGcdwgV/xILYgLV+SiHK7pvW80yd1TsTuh9NO/
leYru0X+4Zk5YeMMOvlCTjGi1s8iuvWlAnEPqCuVRrPhnrhY1moFULkCUhjTzViO
ktc0d0jgL+giHBncHkEwSFWO3eUme37UXkwIHWPdDoPNt+8apsh9ntv+sNiBfezL
gDVH2bAcg65iZbDjnsNeUvoxgb07yvDrp0lL2fYPOSayBp33pbURkqVnW0tfPkwP
3sBX2Bo40/13EaA6CQ8K7Nm04T4JFCYrpvD4aPxAKCRtNwf8rqcN+JDGFgv/hPoA
/kRdEVvB9A04SRjm+jIaEBKNw8Q/yD8voxAiIoCMM9/qxnxVL5Yo9IVaXitwe54x
shmUuhnxoPIK+p9TgCTt0gOxXtMEvv+WILRyZ3VZCEFy7b90CVVpoYcJ3si/3D2h
MrEGkwiRUou1DadEhF2HbkEsldZew03s135livhmjrQgB3Mqf+6NOqcULXAE073a
nQ1zfgs1TjfmpF+vQAQ+Gc8DGNPasWtKDH1hu9OCLToOl4v+yYfLl7CG9dppxkFF
CelsMpD4scI24xwrT29OLbG43U+vpJ+cLCeBOwbL7XKKxW/RgR48nHQlbZ9pfXn+
Mbwlog/oRqIYlxNYDlKrwyWXw+tCB4SSFU/1vtxrpjg4W0rB8Y8PQ1kOujo0Wb/m
zUe97IaS1Q+jmCGC4JrpGSnNNlOxlVGMLTWWibC4iHJdrP/fDapOtBoJ0rVAJxpj
blsmYszQonownyVrzk+v8nqMRKxSnuTjR76UTATVPSQ+Cyk4cBO/dH1D1OSUPEHo
vuUU+B1macUmSwoacej+/B6ARMg48v2wQeKDeWeuYPZWg54L5eB5Hctc42Ux0/Wu
TGlYnzt0osfD74uQ6lWUtZ3/2S6Vt8IMgb2/Vy35udsJQg3rMFrQzvdekq9ddfmX
Nz+jWNZYplKQwq5xfqVClPbxgSC+0R4Rw6K7Iy2pg7zzbceAZQAm6zKkwC2PPaRl
XfQdSsI3jaEWnZNENSw8kVqh3mu0CfbaJiYaU4TuJQ5W+boa4W5V+UHkRrvjELNj
JZB464nyoeF7eQUseLS3oFq018aHcHMfjASwHVYB61D7jwd8XXyVpi6ShZjGyDjS
FSHrFN4hMU2L53ucdQtVgBC5Xy4kUaOJrX5dWMqMSbhl4wmjd1Fu7rAju+fntZRz
2dBRp46uCIV2AEIO2foUnXUMcOVdQLvzM8om60uyq4qglmf2OqhUepVp3z1TwTzo
7vQtnPz1DkWxlGdt5G8OrSr8bGpyvAsdsIAR1O+YUOLWU0b6V49vUA+i57Gk95ff
ldNjU8730mGoAJKzYSlw3PidLEu4GSyn0+K2SYFNEHGTnZrY7R/bynl3HqrOSvdn
6ERqoL3u9XdqQ9UGAtIjW44Ub5kG2FMeuyEpfJ+lJklh0GZbPyFrlPX+HcNd3T2T
K/ihjwKBglkT6khcZC4YkS56CO2SouL69Xx3iyV1xEZYkluKUHRA+8WBEz2VpuMQ
hHaCuOJ5hNDa7fznUbfud9DsoGW+NobWNwyxtV+DKGCt9Moj/vVc9EUmqdCObZF/
vju7XnfC6R9sFauSmsfkgAlGbGNFRPxVpc+wFykb5nbDha3peYPvg1fEn0JaB35E
MGB7pmP/Zoggxe9/UiM4ROfHvcRoRBxoS+Dj9zd3dDqJ/RPzUjz8htEMvr8vCvS+
iVUVU0mL+3kfjBLzN35Y0q1l4zTum7CliMHPo0lwvjgyDqB7T896jT1Zi3adxvcT
E3FlT154Th/+So6KzSMKKWmdBtp5H7QlccbLwXlEASxV11Vc4q4oeZ9pp0sC23rs
wtjs+OTHvydBjmRJQrj4eAF6Vsfpt/4XLyUpqLR38yt8O01XpahdnDk2naNkSmK/
gwSe1etaOdLFxU8T0WW0+5Z3qYyrSHti+6tFDBQytrHBgE1XDYz6KD0O1roqAlTs
cABo86xuGrvyZaRY4cXW629493LrKRRPM6HWl0BbehXCgRzYSow6pkvCu9ERmB3u
D4INSg9/ifhsBGwH0jFEMPatbfS1MTPhNNVUzSQMQnmroGLBFfh2K7ln5JXtwDpG
QlWtpxF+qzrauz/J8BjU+3BfuYN+nCF8sPr2v4KoCWBGEMN71b4NxrCGIGewKKKV
92oZVMaDPOEDNpEs+Z+U+x44bDy3elDzqAcM9r2LRvRLVfLD80fgz8y2Do7uyEK1
hl4JWnPZEouWfxANTCM4ADhd90E3SiVT+lb6b0PxMeQu0jwjY77SiIeApVgb9GKr
1EKOeVdPNsT1EqMS3xYJAfuVwGpAPIvWW5pnUYdCpHZUYE9Pqno9iUdHOmoac5Q8
l/1yHeBfZG0vSfCHS0ayFXXKbJDu3/WU+3bT+biEUzNz3vYoTbdecYHFyyplCwHJ
tZj8ZxCkHIWHCrown5SJb+Rc9PWFxncLPNKbHUEYr5rjT1+ssL1W1a2wAHrH/lxs
HsSiYlqEkmpxk7AM6EnPLDYrhjxr5q6a6sgbBQL2AaByuF6Obl7pw7hzvxqGdkAK
o/2frjnnLEYb6IeKLgRt8LfIjZPKFCoAWX6clgx+SLBtwylXhwqwNDk7FtNUOy6B
QdRN7xXpxNockDMDw6aLv/j7GitTDD5WC+CY5w/NgLFX8DLdKSEujV+48QUPZab0
y7+FyZj86sELElaWfWIK9DQ86Cq9ohoy4L0T80VrJynncBfqFeyJvxf5C9RRxLPi
xt988hUf0f8r8B6GE9didtgxTHMvHOOdIrj4UztW03WsOOMAqzLe2aJ30WcvaRpv
hlDUIXSnhAvYZ01JzCeEzP7N1BTpORjwXVlB8nNkY9+56a12p0eRgbUebnP5rj4j
hd8eBmsdKpTBfSoqx1GiQV2HDspMKwSxC2LVIqVngQY4O2vdeqg2F7uMQO1DBMSs
hnV360E5IWwfh88griIPaEuMJDFcTkHM3wi/wWwMCvkviNd+F4nQqxKCQDy8kPLB
F3ecz2gLt4FXBZ2hELRqFDS8lgujOFO23Gndm4xS4aur1tPANY63HX1bnUD+SzIh
179wwPGKo25KV7a3CCdVN8EOrIvEjdbTWQiAMw2XYZ8y1MqNMWgcr2ikgJPtaAsa
jcKBmo7WObZYKpwCso4IvuuSRSIfqXy7q0JO5WA5cnmNFdwC8a+rtcFjJMXiPtS9
rpyoqE0HsHvAQZ0IYsMYs3qFaZCApRdvuq+YQQds6Txv1FTJHj4WU1hCGn8Cf2mA
RsrElBcCkb9fgc3YZZpJIwvJdlwjokLgqRTgjbpxXQrYsQ4UcW/HbRh7AaJwW56K
Vak9eoehRI/KUBaBoN/m+ShYs/xnNFDsMC+Vqfa5jILOjR/J6S0P5OrjecLe4Axn
mY+t2M2rlaQWCmA+9kYM4F7KqsbtyfGI5C8RYI9EbG1tSlcYI2bd2jagDdVyJKZK
H0cAM8g5lcIeAepRsWtrzqdnn2y6q0MWOLCmOAN+D5930U4B68WYqO2D7SdKyO3w
gqFyJUJizurA0OPsqK10gWoSHqfaX8teJXAv2FSgI7tGVumRmgcSfEZ3m/jXukys
iAHP01fmAfF732NiiT02K6HV/3w3jTge363sQCzCDNNxHDCMy4dHOm6LlEomnGq4
i2FqeMOQ0KLz9dwE6bmh16kKr/xG+t5iV1dHeKmx8NT85sbRC/s1y2ZGXV4XsOC+
uciiW98JsMl68gtrKC66AVR+hYdIapoTXGXHYkoAd0RBZDf4RCyEtEK3/C8mqqAP
SaM87RBvU0XLrXgfQFNrKSue/kk7FwaqKP41x/vNasqv+nI5NJ1mcZcQiKlXq39H
LBo5L1yZaEjzP/sI3hEr0LR0PrP6t1FZ4iPW//nvjBMvoYn+Wz7gdLneIyHGys1f
KmE1nd5BNXzfALOGEpU5o/o5NOanZFciomKikpvEZRhuBqWl5LCo2EFjJs9x9WkA
mGK4wRJqIAFXwHuZV6J+wkjVVnZ70WM6Fyc0n7xkRjg9TNtfTbSHjklpGh+VU/Xa
I2gaH4rXWpQHqJ5XVcszVEjj7uifBjPeXDuN7ryeqkptpST3QF2z+GWFvxYU36AA
LzXr0pfYrM8CsBHofxW+FNDv8FfGxpiORi4nFFh+4cdc+IY2e1Iv5ll4+lid4a/e
f65Hx1Fd43334dxCku5lQ6KqoJn8Uy88na6X/6bkhqFT3F4EhImH8ptX8Ulk/dYL
MWIkERfhabsSlJNIwmcOWvhG1mC7WQQgk7RNrACww+Gp0G2Mlxp2bJ1UVEXM4/Vp
hHwiCsS0g08W8K8XgFQ2jmUM8sBxnkaub+gJoqIZz8G4TUNwKtdNzyjdx5XUYtMu
dS9qHTz5Ox+KnFx4gH7mmliFOtjMMbR8aQzwYY0klJOEeB/piwVhAZjnHEngLHzG
XjRMs4djHCF5W47T/ca1c4etXQg9oxNLzqVtV/fAXQnEnesAKMRiD5PGlMNOl0Bc
yBvvfsClqnRFleC0wWXI73B3tVXTHLrZ6ZdsyDkje2A17Zxryqv+kkifvL9gasZU
Z48dtB3rz72H+auajDwBpiCOcuL6j2zWay7L8x8pkxkeqPBxP7B7OXFEfHr27Mdn
rl0G1noP/Dj1u0dP9QcltVAoB0wdtgipJa1nJp4ji8zWDT521IHfLr83qKueaAKP
04juEHMSLbEcULwOWxO5n/fdmVtSFgnchUmPWxr5GTmcPq0iwbb5/oClNhzVdqbY
pKi6UghnHZ2Y0UmEhGDT/ajCVGj3qP4+rOqCNN8pr4TtOwN36ol0LSxYZJnhLQQ7
/3rnDXayvxsVqgbfyrtBd5pv1m+DQJlCo7HxTcqsChkb4dmPqT5FVpUGWx4rjYQP
IEPUyp1Zmc2qprSVMls7Mm0mlQKTUKb3Sa5Pva6xocuAe0ScVmKmWeJm0EU+sT+F
3yYB3GnmBNAlFwRQVYQYEnuinxbIWeO3hhXrOv8Am2myRrVtR0MOjm9+CLSYKQe5
CZkrlLKL0N8baivcooO/jyHG38LlumBkXyV+R6WPNC8HlPCn2ej/fgYb+nF0CwtZ
ZhRIBGVf3yZqRrce8aEs85MD9LtF/3bWUYH7o4eXHLuuDm7tvD/ZduLRvyG1rOEw
/3IiCrk2fGFcaK3Wg68etvDL5b12Qcy0vgohuAdIJiTuan7f04ulYuUDiwF2BQVB
kwGRuZ+NDeVJmpIHEWQPE1XnWkuuaSh+b01JvVyAW5jyJX+TNND6R6w+I1b0yYXi
M2Q6zNRCAajOMtpgjCC5JSjLPYEJGUye/+ZgCIZ34gFfkel+RvAqXOHh/rDd6vhQ
JucvAjekJd2EIdwOXk/zy1psvJv47WiqZJiIf5rMXHvFeSlIqijP/qt1XWysujGZ
VkNKYABiDElTOyyiOe9bxoVXtMAiL9rnRl9BQS+2r/ZNDvGYh56P+PRyiEeWb6SI
+ORm6pkm+FODuVURPOqHFUhPKca239Zw3ld25p5b6NPRzRmNKWwRxDGxfbAbdDaE
fFmST8bdHG6Bf5Dw+X+NpHPnNglgD/tGBC6yp3BpJWomz5pMoDoq7XIS37t66Mpf
+/utRo70ZTV8HHNscuo622OryNhuWLCD+JKg+HjNgnDstAjIgFhl+NITDvhQP2tp
0W9Uf0JM7KTmEdPsOCXOGEFpJcLiY4uiFE/BLH+w0cAOD1GxFLW8F8swisKZYobW
4s1Y66GBbvPqZfcZhtVX8D5Yg8PTv/dCAL0KGO17D+6SXOmIF0KZu1QebH3QfrKf
FdHXltYBVLpxiQoVXnSDcuW7vO7zUSQsS4j6fqYrlxukYUU9x+SKC65nv6E1dWjJ
nNQVccPIeYer9qsYoiy1iJopNP4w6NAsqAD4rpn/rHau0XqOTLAiMrk5bZQUpy5h
oAjjZFhvIX5oLAlGgUHf5dZ1EFDwjjtWCwSxd0mMMxR9KmWQ+PfDgOo2v3lPI78h
n+KN+1jom+Hi40S9YyWvWjoffAJUbcw1y/RBxjAbS7MhK0SNr0deY4xhAuY5lLR5
fINCCX9QDL1ur2vgFo3iKBEa7+E4KP7bX+fHdBbxaxuHxYfpgCUoMhNU1nQH/dDT
XzKMQdYsMuWVw+J2hwfiwwBV31NjR2HtkzgK3ywgcdT6mojTT8ogT3nPq9fwG/Hu
pU0eyyV4ZpW9bAw5P6YmqdNjeDrseFuNJkWVhzTHyKkT4v3hUJh/9HP7b5sxyvkA
NJ7Q/UeN6wmcVI8sCMp8nD7g9bJ66NGrvnuiIBNXteJJlyb2bSrSKO816PPbVv42
Hy8iflmSd0jBTxlsrKWjBPp7zSpM7XThQmb5Nh7p3Xx8ssIYctQ4LcL3EUXrLYUl
kWxoLkal1yh8FsEavseAzUv4sy8mzSS2MB8QblSzb1RYGdfuGF9o9Qkd8kni/7tm
O19x6OkvQ9NwBs9EzsNsJ3r58KOsN79Th1HLMIJ8A46MxZKwlqACZLCrVovZpCMn
y4WxYT8pfNkKnZQNpZBfY+3p+ew/NcGyT6nnb3j8XTRoKh6hThfB6Xv5blzRv3+h
DpNqv4f65mEmCFKZ82yCXmH252BjGAN1VgFrGkzoofcHH2jiKgtmLPgFrtTMgfdH
B7nHDul+JfASRy9YXjgFq3g1sYzRITOnhosI9F83HwjOIPEDq43tbazh+gv6Ts9U
EfRmZ/xRH/muLmhH17KmgB1mkTuvjJaNGqvdlh9V4dVHQV8hKAimLamaRa6cqEap
Lz13j9+XaHm9l3na0JkyANbcCKmYOXkP0CyEdwM3heuifONwJuprd+CxELhuDjXv
s+uHgjOIxQbxptKDX21ZpONBnY9MQzM/FdXCq4s3vbuA+usXBjonEpzGjpHAah2v
rfs7Wv3mbJDpPTPAs9hZ8CVjGoOEPb6QFsUrntz557RlgiMlaOAAbN2+iM6TyhTY
YmKZoJYhru9jAHfdLeA+x1E+cGo2OmF9+ccopf10gu4hZvC7Ig2FIP8EJnxVyQzI
kB7kzE2OQJbZrQstWGp1Or/OuL+5WDrElNOxjEr6uahGI8VAvplYvweSvnr8+yZq
21+c6Yc3vdn+cQVoNAAdpozoN39j527iwJOjB3bn99DeIGnTfyyzaZGEwPYdurPX
rzgKX0wBLk1Ax0gwRTeLemCs/01KqpGiboLy7uWhQwr0uFuiQ3pBZWkEm0kvlQw/
6Oj2LjmzB1C3kAFv/N72yRZOIgaqx1pZwf6BkVesZ0AY7JEAGUmkC+mTnhiFYQ2p
BDqrCbNPqmfcUGhbRh8MSmB4A1U/tctMiXenUKz9LJK7QbmTVNYGfQB5UbQizk7M
f7Fvy9fWun5AXs639BQaF08+1h7lgtRxF+ZdNdn4Wjd+9Ay6FGI5ah+8mOpQJfAm
Hh4MblhQXaURqiHLhOKs+LrXS8pKwN9qgRxA/HD8KDgx0XRBHwwEJ2MKtO3wXf3W
dc9irK2OQ8+hsZbqBdvao7wIBB0PqpBWsnRA4DX6iqFvsvuanOvetiV5D7mpoEZN
HASUb1cK4HCn+48ocgkp6UwWPwOCn/eN/nM7oBYznVh6gCfo2ma+vSa7lo29gAfu
4o6r6UtLrnCtxfCFYYTBsPFga/GN3yBW0WK8RDrFUv4XgtcvyFIV3M3NgQ8oTBRT
e9N2PYCFAt6tC7vPxuM7ZLTq4zVowHGpWGGvpUSpr7RhUjE79ocbSjdUz9ezZz+2
F7aA7pyRe+ZYGf/bv2E6n+mzPcCIAmwEMCo0b8wapDHnWMdmA66nNYC16P5ZgmfW
rRLkJNOxFuXrKO4JIPhehby84LbktH0FQlb6P6jrF85bahMB2dFakEyubmPwHYJK
0zxBHGhSsNwXiq6NsuV8m/uHwYjhuHfQ7Ios9zAmeA2n3eKJtPRsAClDWHL+Hu7z
kNgRcAIIyjX0zCvPZ5wxGadoI7gTtfiqENWqWRc3ngPc5cjMpvH5IDWIrJesao21
1Dog5nsUeKmU8pPtdwPd7NAl4VQ5ZpFr01Tm1AMm92x5UluJPRqG7olKHyOOb3OH
A/osXB8CfHCRLj2Uz9g4K1sGVUEmLuoUCteeqQZr6O8qtyE+DvXywdz2clvUYopa
3ABSLGLckF/zwLAhDhSG9rZSdSiNvIJSgyQhSeNThV/p0qHH0hWX/X9sB9d4BmP5
vEdCmnAiz73nFclF95e9217IU7EDOkEFKtwvUod/wVqimpSUltgGxr+/3MKcZrHw
oDHtWIng2XAwMUW3idAryzE4TPBWtWxcZ87RXNk/IS8WOpnv/X3GK+f7jNuEjtlq
Zsi9YXsvfGC0lxV5mi1s7t9hsYCu+4b3iBl1fS081DgB4yQocf4eLf1qJMlxXI+F
BQHPsMix7NUj8qMFAnifCOfR+qnb19Nt0k+rRVKweILl9FWasApcN9XAOEqB2va3
jWrgGvdWptqtUldZmuNISuNvdC2ki/E57v8tbZTKz3ZcWqllNOj3zLSrm4ucLpAv
7f6bSvtFe28xsmSRntQ8cmT7DhBP+0OPYqR4uG+verBOV5SeXkNSDporX7IDcX4D
ITO046aX9J5AZHMojIRryzYp+MSWWFuvRz15p3tDnmN0a8TTgb+rR6R7K3qn19RY
fSjLXYDDRi4hy4wDTDpK94O1tjD5Td8uJa4TSdFmbcTClsqPRS5CgntVBsSnu8aJ
QsNFXiNRCcvLv9869L5rhXCa8qaN6tIo5UmYecyZCidwAID/0pZiN6EviEVyG3ak
Un01NKsv3wf+v0gFs/72nO/PaSiSXOOfMWhyoOVmeXil5IbCEOcGV0uVgSS3IR+5
CmXZ+X1vo8Zk+3NkiCbMyxAa3OUcN2wj/hO/FSN3BJCuVPhZFcLErpChf06fV2qF
6vBYpAzH9w5Ph6xSucAre5Bq1T1IpSl8NDEz7k4ooaR5b0EUD7Ii/bZAKUVaCHL3
SQJdhN5rVr+01e26ToEJZ6takl5SX2p/MQ7Ay3Sjs99LUvYXkHsGyBV6R8R7U5XZ
wuluJ2ddOraEzL3eNoIZ82pIaB7G0DKIBys+rp1QF38x4uHmRp0fBqelAeNhXLI4
Ej6qUxJzWbqKRPaZpC/S0JiEG49NABOJeAi+2mwCR95ksKuTnXMUAtnaFeSyVQmk
/KysQNwfaw+MiWk716C5bELQgUwz42v3m18VTuzN9DqXkyof0Y6HmD8Hr5/DOFH2
GSf0hcYY7goYzTodnAHL1icvkTFAvsla1lEh4s9ZRvGpMrFJApM+VE8LR6XBSOMR
3UH+bYdTtddC+C5Fe6nTC59osUiew9D7xPoQdyWuLQCxeK7kdb18hVdZmAA+eBbw
B/QvOG9U/0EnW9V3DlQwQodpcSY+tXEL8c5l9HniY0p+Nejp6nkKYuV0ABPQIO8t
0OQ5Zcof6M1S7hgo9RdbnKXgDifd0pvrFMmZgbwIhBR5YvvslZkpXMo/17bzvh4f
i0dXmZPqM5orYvl4v6nk/pLgi6Fz4qGJz0/0PRjGSb73GqaiIBqJZtg4nfk6Aogn
/KIhg+72QLXv3nH3Wjo19erO31gNR04M+qiqLfIEC0aBaPwupyMlnyrXz7T9+qBK
eConYFOurYV+bS2zcCfI2eRa/etS6PJiuM77tul3pQdaLSVj3EGqyiUkgZyIdhwT
3tUtUqmKll/7v3wzOj0KTCFGevMABVTqo+Z1KAMhxU2GCQ1LjIklhJ/iwR76gNlp
AgqHY92PFOYyCTs11fbJ1wXZ2fBij6up3VKzrCKlB0VNgwNp7eW+NGn1gRmC7GM7
cRuUsXsC6ZBCFTeJ8rXkH9JRxBD1AebzAHbte2u4ZfZAmJsKjUaGwwDeOk/og9zu
mBjxWZTxHyZtyU7XV36Rd4SVRoz2sMA3AYVLVTaxWczriJAOiTLf6jKkxPkrio7O
D2xaDXAq/jl7b0w/A9lsYJzwkdIyQ+cuBT+SBYnOVcc4+s/2+LjwFBhU5+u+Cdyw
PNC4R0ZgWv92ij6nR5dc2CQ3Sa3m6+xrSTTOzV9kAadyO4xbkmAIwWiMpc9xkdyE
bcpjqRiLYgS0bzyuHZ8KA4vEUXaiLnxPHYJFkBTSag5rY+MvkGBla4wnEP0XMjXW
364Nv9GFeJdTVUywmF3u2D9XJLEUGod6Pul1YBVs8eCesunXBuSqYH3zGIO9tNUm
I3Y7Alee83qRh5qozWDVJq5REE2kqxRCHX7C95j2b+NLWosbHqCYLgRvn/BLgdtd
oVIc7BtYo89ICrw9BVCIrg0GjFYF6ySSmq/8ZTACvC2mrpj/f1NIjQPlEUvOUUJw
sLXaooDqRdq+SrtSYn2DMXvljFfCiLxw9yvNCAH+1bvWfEdwK1Mvy+pTMWdFFiaI
Bjzs0iU4z3TTekgwMCS2YTohf6z6I73GAiMZCLkx2TEhyDseLhzsNCfJTWoGSNDU
ALA4LMwDsZ78+bGaZoeCYJXaCwpoh5HljDj45wzzb7D1j4eQMXvxsXkV9RczUc8k
UMeHERKCB6Ev9/o+1iqXo19t5TPOZjzeRRXKpAyCrAzOnJBKjiHcZjjpU+yQqNLu
m5BmsSfNi4M0qZSO8d+RfQrs9izjnRJD7zaqvO+PfWirWjbLQG7QJ3eRPWM6gSkU
Bz0xH+rk+Mgo/nvQhJvg1uknj8oe1oPnQGur2RKrxJxmVrWOhG26fbQGrwXjd7te
ria11XlaRZtdThgaQ9sUuF0wutNgIT4uEH5/lyADVpQXqLlq73LWrvxXXPqY+xeT
FYcWN/QwP4N0ne3lCiH1KcQYHNRL3VfwGaITLzQMny0xg7vM4TdY9m4d72yGwsAK
W6XsIJRnhy4NP0FD81b+91hSkclViEkQD+yENkRThGw1ed8X2wsl0GRV/tfi2lKN
qiv2BrCjfZIcXWGJOKFoa2rpQYpfWAoEF2Q07nrNSMUSunM1zEXJMofx8pYwRdjW
KXaZZaLkmidhGlf8+BgBBDJbggexZuUdtnJhWJAuUwwtnQ/2BZUve9EKa41ykSMe
jR7hAEsuu0rd+4hgsgI2fPPnhaekl/JFBt8TREGJ66j+xxWoLV7Dz9hnRCyOi4Pv
eio3epYnSnYyp3D96lCwGprRac6mRpEMGImte4dec1PPHhP9j8xfbDzdFn0uuY9Y
jzCTrT5OdQa3tu3f+ArRgxFKsLijIR3Qx2PBcKX2F6B9s0rsD7MIwwffiyo6yjQK
l7ptT/JmTzmV2dfhbSauw/dCq4XT30Ssk++Is//+MPkfRjGYHuL6e2u/OapCizD9
eMmcZ1+aNaGElNTqh0gzk9CEAYG7OKe66+ROzh0/yNq1QiQIzlnYKBc6hbSNECb6
lXRTW24uGTvZTXYi9ke6sv5prSYOgFAK/XL5q+9mGs66aO+y36828oxly9COEu1I
lT1aBF+qxqg6Tub3/YX1Isr854+OHdWtE4RPQPmslgjxrcmQTaSVghxwjL4EnSlo
eHITLBfluaQGeqSZ7izTFqRtOpNld77BO1AUzizksBRllykXgw7hT/2Fff/Da7m9
XOoaOGa3IgWgm2uR1Odi8Nnozoi2LD6IvBedJPG2MsQelXsDXtoYJ/3behg1bbv7
3kdkAeWq9ttOZ91uaORQGvt4WXNVX/VWDAaeIjvBjOu+Dnl9WGfxSA4vVhI11TSu
JtNOd9sQ4cfL12To0aQ/+FhIXcXW7iYB7TaMU4BfFCsEd2PIZqMiU5KcwDxHF1VJ
sD0TpCYutISZpy4pKDQoVClgu7peM7Z4wYExyWHnvmaJkdKbHfIkH/VLf3+v7AmD
iRIQD24cnYAtnoz1zoPoD32M5gVSoSKNrKsoZYK0PUlbBhMKIWt5YHYm09QA2bzK
4Z3ydAh86CwfmX39tlXUqsZq9JCxeoT+2zeFyyh0HIk4iKRr8EAQqgzvlgMUlHjl
iP0jHhJFO/83fPN2349rNjstD6nYoEDDLnkY45i3ArKWAyD83kMbRZUmzzJ632k+
A5cpFsi0K8OMNhzMZzxoJ0JN0TC8O2gv/gnVqYRJWLZ9BPVYpo5uOtrF3bafi/MA
ucmVYAd4RWGWh2k3qY1XemvkEUHG/x12ebWtrIR6BY+i2qlUIfBNt5Cl7v8m4Fsn
Mfv9lYD9PNJHz61oDdAaghqRb38TrVBjm4L02oWPIAtI3o/qkGuXw7180uiIGcEX
cNi25AxMGqOQE3rpx5LowsoAbkWHNAv/wnHrSlCNxDDjitOc2X+Kdt0S6j0+mlV0
ENTsmfDNlaXPJ9IYZK+TL7hyzeBZp7TXPHVwne/KggwpJbj5WyLUbok4CXP8/wyH
n0uOKw/HPG6uHff5rxa35EYXCQXr1smBlrvDFo1SEWCkFBvP0t51+rZMNjfsiRLF
6dwnHWxL2qz+3G8UmLQIJxv/8OFQ4plyal9KNEanz+sQYJ+KPy+W2uaP8ug134RW
DtWtoiPKAgisT70YzLlMNr6qiIoWStPEZRmZEn3p0VBDy4Ixpf/nGuMQpXu7j9b0
hStm/lFy1XIEmo81D8GZXBqWaBY0hskR/HcopWHd3tWyTVoNui33m4Nq/dSxGHNG
RcEkwBK031bX2Dyf7+FbuS8TG/oQLz8N8cJQ2uk5Prrg01++Ty9DTeB6mqcTnMum
yYTKwk9elEXTy9xDdeBWL38EvV0UJWbXA5/LuSa0r5qpXLtyeVm9TsbiJcEEzknk
vFDljuro7YC0KUSrkXDC6q+6kJTMoEGRB0pL9R5EmvgE4UXqjx4c6/MugCtbO1r5
kSC0eB/t0ksRVVvoFSPxr4f+aOsBdY9IWUzXbBkQWteFGihW0/i3MQ2jV8wZZYWz
zoQPkWkXgL2shaOaOsB/t09CerIi4Kv1Q+aVYx+Iy0FB0oKO2p82N4VaFgonMgZG
Bd1j6iCX4OhbnFnBppS1zwzOXmll8rOkKOabfkllv8v/2nFjsIVT2CikB0vmzxUA
nDkRKXbuD2pW9B7pQDliyQ4tWDSVeF0Aqu84c/mQzvmxi1uyr7Dh4PwlPey+G8uy
Id8bj5vy5z8sSTQgwtB5NpoQ5/GCGo6pmqwTcJ2AqsL0mQATKrJ0nDpwbettDW61
sdRpuNDwirQLlezVIVbvuzVqdoEjONqoMgnWHLFcv8s/q/ZbIpN4fxc3tmThujHU
KTI0vKdszQQ+bfF3TxiXqLfq95/wDrL3IbU0I7yHcC8zOq8gnSFWjedk1zrXiqyy
Vz7TCkT/o6YNaO6DhZJHOuE4SVcoZKcHI3oFs2WumAn7YSFk6OHAHCZfmDyddzqd
M8H33N1ZUo4Sswbu+wld84Ywhc+79ky6PmZ9olJjhMdlv6PKjbpO1G9q5qlATZGN
HoItOS55cHrqSCELIqTKvJtSBGlCZJSZGsPVRrNbiJL0QuiDMRvRdGE3ADZG2Nok
71anGHksybA2VTlWYx5MWkRquRYhUq1cw1UqPRTf9/557F4hE4IrwKJYj3A8UFFv
VsAiKrTRJmXbSuin1AE7437S8u1U2aWvKN1DX2WDFkSrndzLn6eUCaG7+uxaXYG9
BSeARr2ru13UXSKXMbM4iBYgJYpf5TpZEnca3hHN4SMpV6TzGMVTNq3hD8CRhCsq
g0j6dTNYGI/olfnzJi53/5NMqHi9Wcrbabv4l0NDcOQwX6KjcE5TQ8ovoPhljQvP
PM7x7yQh5fdDMTXfWxTeoyu8zr/uvmANL9Vu5rwk2d3SRTiQJE76ThFi374elbff
iY6QMWkLzjYFVRoX4vPA6YTCBmZ/7Zpa6u64hJ2K3fofBQrxZNeMeWBNSic3YNZG
fxZFmrSoK8rGk+IkdXlvP2gWkNuSe+1ZkgO2rzpl82d+3ICMZA4zOdWDgO3NgBeQ
010oANqeFeFmSdcqmUSdHSgm1d0fFZguS8l5WSIXJ0nAJvYGEub1k7AP/k3ZdO2F
g3+hitN79KVKgcnxhOZ/qB3uKdc1JdWa+6lclVN24PTT+hAqPe4hoxCPXktjlVWO
CU06VbClCiR3qoTzZS9S8ob+Incoh0Xtyy2wzPdritSmsPoVrlwGoGaliwlTwAQI
jk4ZyV6uc1e+yGQlVhkqBWS4gTphSDrxv6Ca2p8o8sAMrqGXvKlDCFJ9HLExYDwh
fVZ1rLcdINfMsyaqAc6G9OyiV9vG0huDG/C5j83TSvwVDdku6v9rZd/AP5MWp6kV
1vDsYWzru0f+AF8oY1e89QJwPE+iV/6sJ+31rmDuX/uFTmo7cSIjnynkkHdoziuI
bH7LX1aRw1j/Y9TU2DVJosVsWQl3ud9DkF0XvYx2/Bp51b+64zWMaen5X2iXS7Jj
w9RbTPTu93Mt3ppaF/OdnMUHe5MmLUSlgEWA5ljODz57/SkdTT91ALigQ8IA+Ugg
UPzB8dlc8IsZSAvN1kgstsrE7lV23AalPF98+9yUR7MdBcz5TGY+pwUXv+usdRrC
OGaegw+L/R5SsgBxazFO7JTkCgVZE1uoQJsDS4Lgkh47BPYTQ9RL/y2XJBdU7pE1
7LzgT4HtkXNC1sq3vH5jMR9Q3r5Lveynbpzv7qVqp5OJyKOL2c8yFu7AG0vQFtqe
EXGO7pJmLL01WNxTtx5bCVEORgJpa2K/KXW8zbFxWHfQqfsLyvbBNYR0aBhODl9D
WtIfmCO0zbb92SsR55CxIoGxmGhk09xIetsl/qmuPm3JdycI3JDMfdfGKgJ8Jw+U
XnuMym1E392RPFnGV2ItzG5f4d9LULcSUcBXgXSqUy8Cfc9/F9c67QYgpG+UqFv9
NpMFuOLq+CI0iFn5KdpGTSfEnTniinLc0ipiWZSMkS0DdXeZUgmeKiPK5oUJsSgZ
NNxgZ19bJURUt84nERY187/egF5G6HU7r1fD0vFqlKCbMULmCJ613Xy59hB8uhZl
+3t+yHdGLHKAhI8C8nDjEhQO+0CMCgr0k+zc+ueHm0NsTr+/F0v6G2diUAkXPr/q
QqJlA39oZHo4uzAvNzpaNXUHFrL7hFOmJjetpQ729MPpt0+qjcULUVnd/d1x/HVe
JU8ErhdhsKw/mKGnmEOHUMjjHXDahpj11DyveuDrMnWU1cJyoeCYcCScQiVUeO1y
Qwq/r/BHx4bbrXXx9V+94YJ26YnkNE+3tyIcT4NM858JweeC5mwga/oPEFJKAqix
sE77oxTlg8fSEKRJYp+evb7TpodjzROqTNR9jlZM1rD0mUC/onpaMfRm8khNqEwR
3ddr5taeSmcC5VuGmfuUySswsm9NSGhusCBzXvp1SkLWbmpLYdoxg+Tc8dwIgaAj
M+Kl78m+0LaaNxknH1VdqhZNwv7SN1mjcYLCGrBNGC/n4mzn8Uj5zuWFTKySdXg5
mmO1R9LLZtheu9JU2O2fcCPSeZsvEO5YIjDFU+53WiI+oK3m/HaUwb846bLhIuh6
22KmoJyVAUkmfnO9Lmg0rjD2XmPhG8r2qQCcsw1VvxB+G3qwITXSq+ZJMtEc3wfw
jLsOh4gp+EWDJ/IC6w48x4M4dePZOqqTzCw0X/VqJVJMu37p+3/6/RjnJov1lJUT
TEc939FiZWE3gi+NHSgKbB9e1JQF8aFWeKSq2IaJuMv7ybtkUbVVCa5eMezOsaZ/
oFZ8UsAawHan/s/RCZ1yXUcj74002xoeIn+Lh4WxniT2aBgWlMkqMhjkC0vhLf0N
F4WdZOqRN/4dm1r/uO5I5OOE4XHvumvY/69TM9Ed6ENFmZINEY570VU44kaEd3uq
01X12daSGd16OagOjUVGYAdH6RokY3Lu5WvcMwLhj14m2YdEicFZrZhbK4kBGWyk
VvisCSEyYTeRIaTSqXT5HnuUT/2uOvrAlIZw1Am+eGhgfSPbqnvE0H90gXATAfts
g0eWeYLHzeRmVDiPuWpARS8sQ/ujafdrVnn5FYdphjSORhEaRzbOF7Qwv5v3PWLG
Xry8FQ69e2s/m2bTuvf80TYrvusy8WDFOzbs9YwZYEIOjptxV45sxYXiUgWJ2jOW
ZxD4K7HBAVhuWZ3upVgYHQiTQBPiFSly7NbjpRmXnL+Vzs4fJ+aOn3tVlvS83un9
tozlbZh4n5gvJdpcY6sro7vhsESiXr1mG3YHW87b+2QyiNJ3LUtWvbTcFlIncPrm
fnMKOrsyPcyuB6zlexHj2m6HCYFad/bKkAOnnWGZJ46nPOB61ZKq/UOs6a4evfxE
ZLLHHo8XywkabBplf+O4FgGZ0tEe+Q5bqOwfKc+R1xXoM2Fc7KpAuAMAGad9YhmS
NKt+BU+5/rYe71t+3lVbAvm059h0IuAQa+f4AfprY5gz3O4o1bJ6pazFxoKRoA+F
h2FE6ydmTYjf3BsocryMjxaQ2Ybwi3f0F6JU4kBgsVaZPIqa6UaS38+FSveQV5Sw
5joW3WsnmpGTV2aje1x5SFBsUrwCATNeTbRfLGGDVppnC+uRWHGzTpGRLVMhW/ew
p0vGdsFHN4xT9bhAmY9oy6P77K6kKfUezPsE6q41HsW5u+vfZTcAmqCFyUxbYrIX
AliUpc3Z0aditrQuDclh6H5pEDvF+EsgnSfFM67CqR+nc+FP8OejF7RvMkZJ4shl
kTsu2ula67uUHsTdzmV04WG0GAPajblL0mIjP9R4sN13t+KzsrY5Qhbwoe1tQW0p
WIRvz85RV+D9/CFs7Ar/JWouVXhAxmg7BTeBSmtWohRofoKj+9+OAgebfc59y6Ke
P5pvZ1P4Bqe9IqvrGqS9OBmj1rfTbNB69s6x82ukHIKIUTk8/Fn7IimpjsbYhs6I
+MRWJUhsep5Z+vjqPa8IfCrhJUBQjYl49IB6UZR097tYE+HFR6WSj3O8vH8vkARa
o6LP6brxKyeekS8DGXLO+wHtYADG/Mw7yoZVdL8fN07axssabb7jsmU2ZVeb8icB
VEuiZEnf34SzHLN/Orvk4c/8QGoT1jzU0GwwhVnzIKWKuaHeJfg0WkVjZa6q8G/a
MoZISNVl1VCL9DJEEM2BhE8PwWaO/GKtBsl5xfBsMBuipthWMcLvJmiuNO54r7Jg
smT7jzGsrEemw6yzrz86prt+eEyqiHJopJuQs5leaxOZlUpIw//Bq3Itg8g37tkY
23ADGd56VGIEuFr6oAvjAF6YUskBjy7VCQ94xQtrOS1Hydu5mcCKaZAG8MAEXtaV
cVTD5+2LP8gL0GRfYmvRgHxzok/FuGNj2V+7Vsb1NfY2NnaLsqh3loXX6mpmYln+
bJWegMhzv8ydCBlQJl13kuaxVzfH/UiBmnQaDNf0L3H835YI8qXJMKCjJhkRhsEH
RztTzj3GgarD4PAjMwtkVW9sa6ss0ZPxNJ3jl2qn5xxyzUAsTbFiAwTfgs3y57bH
6csYoNIaWa6Rhj6VRESWsrgsa74G8kXOG5umMgGFK9m0E3c3x7S/8mcsI7XgriEB
GvUsTPKwNtvW+eqhDii6jo9uMiSnbXVuoxjUxoFXcM505v7NdQJm72RyEM6eQu7K
Nr7gOJixgUOjCejC0PB34C0ImANVgDQrTCKir1YgbzQmUSLv/x3o6xCmpKky2mRn
QpCKNWfFI/muA0J2GigC3q04EtfzaNh2eXy9UheMVs8S9nAvxAY2QvtaPFcIZGgG
ZIlx7xbYe/fO0qezGZdldA1DizUWhqNgc5yzeMwhLsSr2FFDmJbQ7JBVb8K6gabG
hNZO2tMjBRNJBszleFwPzCuyRIrc8UD97J+19JEeQbY=
`protect END_PROTECTED
