`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yDsxEVrTn9ph3tDtt7+aO7Oe269QF2JeAYY1YP5wm5RpHLhOLbQYvR8kxRtdpjbX
9URWsMRp4B6CQXdCm5z/Y6/hJMoso0hSSSo8LO72f4iOvQYKeRmqvOCc1U6OLLqE
rdJWsHZ/BXkec6SuHJ4cN+v253T7JJZAcX9/xi1QKbqn24cNAykXc7Chk/rTpPvC
19Q58crix52dw1WM9gbo8EZya/h2eHYbJid1TjPK1cYqOPnKUqIjRIPMdMY6SIdT
2rpMY6aJ1FXnlyQ+AFTS3mBakQK+pqLR2QXlxhNeFjPMkONx/69/MEqK0dQBMnau
QjOkqIQZ6eATMLasLbJlQ3LVQXrWksjUrYxIJA48lsIUQbNGEjXKg3Y0MXE7GSxr
1GclQ/olrFXd2E7tbcGAml/Enn/DtGYcZaGVBqlyWxuvEu9DDBAVg7tAHOZiEBaE
9uv3weYjz1pZP0P2Wn8xJc6QrrorqT42ZQ8CZtwP9scMrNCyD8dshdccp4AFuQ4b
R+MXxYT0nfCXyivIa5eDvQfNyw3JAav2X85UMO1JIPs4q3PsUmbhTeBX0EuBSPrh
D3uAfM+HYRJJcm60EyrrmR6en7p/VL7Wk+Am1gan2suEa390dnnWif3oKNPOmGE9
SYNZMJxVBe1k6svMSiakPHn4TPINoe6ClbIcI62FhU1rn1H5Daf3j6Nwgo7SGJim
u8AESCE/ewXMXpGQJtfbtkt52MiDBSOOtkk9H5vck7cVMeNzhvuD9igOp/yYSzgy
GvlKj4SXVTmXnhRJ+WHYM9nWQV8GM5Yu1J+ROnb3fqXcN0sSO96jzi4VOAaaIIAV
3VHuv7fhmw6rwCLUBnRlU17aovQe3BCqNP++fhjSCT9h/ASksUMJLWzaQnWGPvtC
ISadS1drgEQW561CzOBOPWaOwiDDcm17QTCu4vnysZ4fzuhLQlXQo5OJGMHAVblb
XXIhL+ItBQaYz8o5kMa6Sil+JbmLuzF00y7Z7g8ir68yH63H1Ev/Me9+1689a1MW
jxPbN24tvCoSEbPWGO7l/tt0vvYmUNn71qbjJL6ha4I2YQzoHTd2GWHovMG/Ow55
mf6+b58hkJTDMTGl/bkEs3RjuExOalt5oG4wNumy1Ac2j8maBYouqkoIUWkm4SFk
`protect END_PROTECTED
