`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cve1a7W0q4cych6Jm2XXtjGm+L2hOLmk8rv6cwuWyeGRwXAslJJwAYnP9sfLiWqG
b2gaEgGo4Q3qC35yRJbARARTvkHKTlxcxcH86YBnTWauK6Ujcc+bCZnp5Pv6HbmQ
k7jcd9gfFC4hUAcdQAE5S1j9qGZjLhPUyChC9JsSUXsz1dHBRyFF1va2+qgl+IBV
bJXIDOaHTHuQlxB1f/lXzO1GmOw6861AV9JKS6cFRc+j6uTNZ478mw5qhxzCaHG9
rP/9Dv2WhBdPqyJKBShYV+7ozOjFYJ5bSQFWy7DblaF9E28XRXRuWigA/rW3EP0Q
7bqz8VMt73Q3AlwB3npL2r7CYIHU1VgNEWrg2oQ8RXtlPhsrn3eiGGmNueMSXuWf
Ad3DXpRCSEXSYI2wV6Yrb635FTvbh1c1KRI1AXU6akVxyMZiNTeBLkrM07iyMULm
ekD7ywxDiud+cKb2GCrDJdvm3oj1J51zHM++2UTZQhVDmEHWvdVg90RB+xaZqa7f
NS//g/jBPSlRa+YHCMc6OIR+kl1uWd0KjzYyBcwjcDFVqp47SmHfE3zi88MUaMNk
EhkPRq3NlQbBjNveKVhpIb0tHA8STeikivDdP0IYhs9bqksfYc8Rev73xTxvZsIZ
jNpeYUuT28fo0a2qWANPlF+o2raGG7wP8hzbnA3MlhUcT3bgAfAwQzhbxdQi3epP
TPqGfbjvB0ykhhle+n/BTdvbi7DpILBwfrbCjXkAnHc9ec95rHi9RAj1HEFfn87a
ycQhH5zMFfmIZR3mlbj+elq1WzctixmHAjyqO6jXuVMvJPBDahYMt7nxLpohVrQ4
3VTuby9d2I867J58Tc/+aWDiVcSgANBqAauU8uIJDEOQaoY5qgS2hSCpTpogMLIz
3ds79s4vM7IVA/ExLmG6F4YlXXCYS2CegTFMRUsniv9Rka7L3I2dwUtYaI+tF72n
t60aRS+2zn36aBnj2ELTBgQZwT0h5wcbF8u1QyaxS3bt4k6gi5p5eKDLDNKVteAr
Dz1f0nB6WtRqVgULNE7uCihBXu3CtIjZFSQ31w1qCMRgG58TENZxr/+2mID8D40T
pVp1uMpgKAAI0dSnRZTCtRCRELHgTT3GzJlzEGnTECs7Za8fKgKteBxbJBkOBGJc
AJOWo610nvZlShx2qs8EGjsEBs0R4AnH8jPc5vKxOtSTeGRTPyBjPjDMOo8MFEaO
0Y5Z6kbcdBZEoeBpVMHHYvM5uRaacr+E7s/3a38oJY4YaRXCAEew/yD5ox1Wem7C
lILXE/BK1v0Iw0bLBLhqmYm6XkqJSIQZJP97dg9ByR+GIrvVr5KJOzvIEjYjW5ql
UMtBGVMW82+8iAcvHuNsvjqseqG4Xx0z7S2hClKv/4tvkdTQJ0E/EivOwzZFmgQt
BTMfaskUYow8ruYjhKzxGOiP5HiOP8hRfqSkCbIE9z6Bogpj0fTFpuLDad+ptfOs
BwUzkAi0Jk5bjxSlhwCTTEbkfUwlw+jSaWOAuaW3yHD9nuAjuE9mo8aURKCPllt2
j/H1y9CmqUzcIjWD9MmiPSAydZTpk/VHwy6wW+pbdmbJS/swWpiEFqlaFuAr64PX
pFG0J5VKADpriMsYa0GseYlnDNGyOklsGINXpGChn/hcyEos9BkRp7iBOQsxkHSn
cs8KtqFO4FrGJ/8gYz3vtQ2UtKdoCBcXsXi72bHKJQqOCEDiFCnG/ZZl1gt2IF8h
3UznGCrYHJV9narJiPHg85RRRyjKbTzo4G2e9dzirCSLrC8JsvDC0r99srcB9R8w
M+agKulmcuAp+EZ+6lW6b/++TraH7xvMBJgBfnuuQ5GPFBiSTCOvhiKuvZEKqQmw
0Qrzbz+I0Tj6uHYCv9RhE2DkglogPivQxBBLmaulQdSQkHZ1MGvTeMf2YAFjp0J3
B+GUL2U31+sxNIrthefWnFv7HuveGOWKgYsH/+Ukw5ea8Brf+wvppw5LCA3E1BwP
/77Q9TDY1XFeKjRcnT1i1O7TeVswOKHqXyHr8llf1YnHdZaFquB8URUxC4y07bMF
PqCbDgnSObzOPf9EbwiOe3D0JWyCvyOQ0CZzis4I3OuhY8+4D3kaVYj60jxzI7ms
tLoHQH6Ro37frfGR9GoLgQ==
`protect END_PROTECTED
