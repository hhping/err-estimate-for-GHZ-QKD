`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/wGTJ7lnb5CFdrR41kgEBCj+NvnxkI7rN/AwrxV3PbF76HtJdXpW5fRDz4pjPUwP
/LigXctZf7K1hzpRbpdjkP7GwxrxV2yhfOe/8zJPTf+jWalnf1V621n0wsofi4fw
VXs60VmAtj6N7W78rkcsumdZ6iinTmAMtwvn5CCSFx9Pj87iZHfZfkgnCU1lShxo
LbPTObAAPCUQAHeWaePoLxmOMNo7b4rSh6svBX9UsPTQspWhEE0hdMEoGMbQt9Qi
mC1wnjRzVpIa4Jdh90xOg0zCvgp4FM9QL+MabSrqWA678qbbBWGjBO3K88kc7HSh
rsn8megS0bJ4TA0jWShNWTnOcTzsnfMnbotvo7fVU3DG6muS2mDchozv9ORGS/VY
fjlC/azyDrHDyrYFhiFG1jPqJP89EQh0wr41uPMdP/H51v2ZRxgKb+foLQvZvF95
RagUGxfD3bc1cATWlP+7/Q66DapAIlbQGHIGWByk8Yl778Z7d8hlnhEr800fXtwc
no+1BCZoKTzkjRC5mrLg+oK81RjtLUdpTTCD+WcfMjpF65ZU5P7VQecUwGOTOvmJ
tR81Oy+BJTxSPhvHB5iSUuff9p+c/GuTjyyi4SuiRVdIBmepRRSBlWGe+X2hpNSF
e1QowpHCWUtsEKfihEZ4YrAJtN7qQH3wAJrcEtZPfHS8oZjkIGmaeWlWx5zRq15p
D4ZMa3XQp5ukqA6/IpiDGpKoH2Az9+os5dvBIpnbLxj9Xwaxjb1GNCwgAEvxxb2k
bX0JmjSIWcWgzzgsx2DP3bsiFOITmKzhVSq+h2sFCX9eAkQ1rjS96hFdDZrQ9t4H
NFsBZWXEeN7vkSdoWT5rhAOuw2gGXQZaCz2ayOQLQamTL5gBo63z5/FxWIkPSEg4
ne+5TI4nK7Vu4yNeDeue/HfGFkUoFwiLAoVVhmWCf8w2Xp+8I88k+dUe2K8ySYcr
Awv1TXt8A9Ko1vcFRo3JkPX7euOdOVvW7o7HtNanoakoA16t0SeznBgXC+dgFhjr
ABCWxTwkE6wzm/Vm4DOmgjoDmuWu1ZGu78ZL1tHMeNDiFdHn+MARdYdmt7oHdxyF
7/1vlZbFQh2K92bI4rBz4RXuGKAlV6Bp9oPjK7b9UrMxuEk2+DMjULIle+nOJbMI
AZZBAMJXGaOvK91ftu56yBqqLYL2SJi5PgtCuHcYStyB/FojNLmaQQ9jdwms2JRM
5FAsOAIg6N0ZIvRkqgP1IiFOizpntO6kyRt+5nxNx7qSIxuJ1JWYqjYwwUDoelaY
jMhVYnoGaFvTcTPK3Hr+zJXZXJ+N4jQSQqXa32t70nbGjBtw/2aaLheh72OvBLKo
yqCBZLtTvl/SUyjmO/UiA0f6ETGlRt+Ro0cs7Lhov7a4J+Vm8AynSs81Woft4AWq
13hPsDvRIF5WKEQkoDWx08z/ooEO3co0NZlJkZd4oPXVX32EUkixhcG/2lprRmHL
2nk+WZMe4E+70jt/jqXE1INb6gwKNZZIgy59+YFFvafs9bKrpFhhoZo3iZxVBWJR
CWsoX4tgn9LlapR+iYRSr6Z/1Xf/5TFdMYF2PTmIL/n9+mQq/SLR10qVkJ1foTe4
sRfQ9Prs+lbRKb4RyVWCC6bcYigrNSbxLFkJV5WMcOwTntk8sRnem6cmVJi+3LUY
QD1UkTBPWl4/YHy3YLigDJaB/0KDNi7E+Di14C+wOqKONUcsypXxJOyyObCTcv/q
Cs7wxbYYT2wh7SVqvF79HgKyW8hEfd61ZqKYC9fwd/xnFE57qSOzrPfh8/uBunrM
HkwEF2CNXalgqkDgQaSaBvG11kW8LspNttTh+IKl9/YenoXMJZlue6MG9sFY0FcO
vvZoYBjlkCKeJlIQOP7yWRLuuudclV2PqQU2WKx18/Jm4wSPPZF1x32rpmsVwM2L
7rNTNaMItKuVrH5QpuA4/n+K5RjGbQCxFfl7vtQu2Gwk+3YpuSPLs23i5ZK3jSpk
/s5xK67yJrrG0CtTxk0gOosIqJ498ZJrH4QOxFtAJD7nKcBu/Ry/ikSlY9HbZI9D
lY1sCDimX6zUCadGeU6IS5BYDSzEVeP65z/182ANyDeCXmExsOQxpzro9ytHWVhS
aSvUsc+ddvd2YKUGYjutBQzts9d/kWq+oAzl7sJlVe8P0N7J4XE42+gmlYBwf4X2
eby7E+FfpUWFwe7RYz0Y3n3dAMG9OXHgNJ+CGycTP71BdcoSEccFw4pqEvS1wFnR
lbbmaSF+IP8MMnp2XhmUdDSlI2oyL5ptSN0eKrlPjnv6aZE0R/A5FGj2JD8OoE7x
D1g4QZrziBhZOOLHOvt4GH05xN5feKSoFelNhMYc23Ed4X/+7aAbtmwl1IB0OoNK
amtLRLiBPKfv4Av8zFROZ225xlgMGMIJ/0JZPJxKr0HhD/7LP++8t16FBaat/c9Z
TMnVh3WD+gEsKr69jt0rzaLLxO99AKDU0rFBIXntSlvjEeLT19sfOZZzFVxqY6BO
S/NFfSLe+9Bd5H1AwfsWzR8ir6HayphSa2FebIR8R9s6JtCbqBC6ETLWk/JaQq4T
+BHwanOOtrBhyaDF+ojRpRuww4+W39iionczTjK8u2lKbv/yqT3MZaRByAVVg6sf
AnIDwNfjEG7T7vtjfhgInCeoIerqipi+duDPJyNHcCKsDKJ4pjMXSu60SmIF8fW/
Ag5ngx3dvIIHiyNyF+d6PdcCU95SKEMFJzBhN9gFDRBrNV712lKjlNX81djS74HW
kRDhDCdq+N+pnR4ipMBjbk9/TTMrzRt1DwQnOhUqVQgAtcinAErukVTRKzg77b6g
HH4OIiU0xnQd8Lsp4tBBI9inXI3XKkVQH3VgOkcKYPgPB0oC+uOB4nbH2npcIBob
aeuBIQmy39LnwfHNYkEzVPlcglx3Sz2swwROx1eTZwj76amOR/WReEtpGpwxEDcw
C80w0wBmzpkHTdwVBxmUZtxbHG6fvFVJhCbLGp/lvifoRDL8Xl7ub/NrUGf/rxJm
nnbD/nH4eN9oZCG/WizTXRF0YMCPuz1ogIJ83rG1FgwWs3xEjzHrApgnkPAUDl4i
KjhGitWXjfvu2l9MrtYfCxO61xQoiALfoqLkytq4mOkWXTCQn3M+9jZhrh1plxMK
Vz5O1/rUxnx0Ugb6jELOcDaYrCTDMQBQIyVRo5HBekYaZFkjNXBv6iPzngdt9xta
yghY5LMRLSRO3X/RNn5Ozv1Cu5os7CeNGDKrZtFgEuFLu4iwoiaUBDFFXcBMmcGw
Fevq+aozsqRIdGvbUaPCTHPP0CM21S5XxgousSdw4Lql5Ysr9Ipu0uzruzyEhb2A
Bn8Mw/L2IQ8d+hvFtUyCWaEwmlY80rHO6eoH/yA3aqFUI0sqf5h4vJ5VjLGrPuB6
7LQeTLQQDtdm9e35d/catWhsYEqNS0NhuhBPplepHabeWZ2SynGcMID+ve2it0Di
L3vj61qCEJMGrSLs1YLImhlkg3nWjFMlGFk+TSPOAelgyQSSBBb9XlzoUBFmZef0
30JimMrf3If82JtV+NVaJilHE0puyxZ4PMGb6ldrFNLY+Wa9THfC5IMZofJ7wifg
9jN4tqG5ZE1nPK2snT2I7FTL85g2JHyQeDFz6NiaSn65WkQ5E0J4YRS5ANiau+ml
x0ZxN4piI52rG1j0+WZFRlLjywYjuOPB8Cnr+ylIDQNwwhXkLHlp4T7MPPFmijmW
bvbQt0ucrpwkex3XM4K2QLi1iHAG9ZXAbYyonTdwfnITfWmY/ddU2zTXeTKG2Unf
1VDoA7C4L+QM/xMlBG7imvDmcIK+Oao4iVpfOdP+rsUQMUoaGa92rhslJpDy23Ds
N/OUwgldo4mkbGHbNySxv8kR/qZyhR5CWQqs8fpQqJFQfFPrXW47T6GVal8w9INi
g6lB+43G9HVbD8XHVOBfFSxxJayaD495d6FeuUfwRhbO2J2FTtRBv9S7cpB9YP3G
k1IgBZYjRyg22tCxOeYNTKbi8RUUREBIFqhMzxX1bR1I9L8k6yqev5e/8exB1631
wsfNfPtSFU7uXEZr1yolr1kfmgkAWB6PBUSRMjv7n9ZQ9yTeGqqhvoDSPKmioyG5
EfAbK0Uw9FUeHeO5c1GB5YKEQrPoGbsgtZD8H3WALJDlG+7eMkIUHLMiaty18oD1
luvdxIKyFi6bNc9OSEoDGpImD4rAKxysSPys0zehlFc2a0PiXhWakzlqR8DuyOqG
TyDCDTg0MXKbOB0fUURohwREdD6cATlYUfXh9TOpWOVuTKGH7PYi4SupWSYPLbkh
pd74a0GFRbWsYe9JtiJNEef7n0utCTOSK7gcwq7eHRAL7jXn3AB59gav/hgUJBx0
IiBqCulpc/rm345zz/f8F+qkMBgZedqPnM8fDZKWa5Rg1d9eL78Ibt7G/IlIAmol
WOfOCa6jSKM+WS80YDBBbrgT3O0uc4Rt70f2aT3UUEuz1j0JgnPiaLd5ElA8z/fr
OQQsWcAs4AGUlcXHTixXwsQ0Uk3uTpG0KuzuBCJFiiklJs57dDg6s39yRb6S51U9
7cSjEVEWds6csyC4SHm6XA9KutFzi4qO2GkQrxDjm5AT+s2ikyQm3wkDf9dBY3bx
Qb6AfE2B26XeGKa6a/uqjVV0vbwFgGO9MI07+VwXgbOHNdiAau09sNIV4wES3Usc
JlLEETIe4w19NmLP1qhyQtH+P6Kf5imF2ASAVePvRwGSAGdUYYms077QfOkCfEVi
PpGnIYIVYjR0ucZF5Dkw7AhjtajVZRVnudjuU4eqSi+ZIbPJcIuj8Wyoycj7KnyZ
BMub/YNA5EuuWr+1/4Wuo2KFMkfn/bL51Ve/qaZrOYeclCxMvhnttGMvlxaXgqXs
6QTLM3aKtK6vAg/YqgYx30fAJxkZ9G5sQlE4ca1PH5XXiWoPgiAZKJ0Mrh1bVOXr
/QcfSgp0dFmJmZ/4IBHnf7zCnurMyLPlLVSiz+Xpp9fDTUhJ2hvk8SbZLQG/HIxB
hSmZP/umujEkMKmtcS9FYUTBUM1mt0KK3NxBh5lzHlYzWa34pKJSMjTt6k0IjWgq
SdpD0v1TOFtyYG7ZfOqa+H0+1Xf/dn5M120WkmXSKH3XPZ0NDSD+f+J6IaVZeQ4s
bAarJZwCwWAZRCn8Kc9lMon16c8oFuMkb0pr8uLgJ62JCr4JNiXy3rmHeX8uDbpd
KHlldi7RaEGgG1JEMn2SBc/j7iVjGPyDeRsG9ihh9cKqBCdX9z8hdwPDdQUNEdif
9YGtY0HJ/6q83QcpxYxOcwKyyhfHD5bWbvjus1GqhaYULje28V0TW8QjhaStrhRT
7ISiKabcqnDxdug4Etd3f8XsncVvOkXZnjDtHdVQBbeaz6CY/euNzmo2uLVQDvW9
AJ2sQ8+MH84Alro7dOawJneagzgG6LW8W/EaLh7cdpP434/TpNsDluzZJzptxzyI
xRjI40OPFCudqMKcBAEUaDs3OL+lGNYt1lSHWu8+ICU90yqGF7V38Av7OOzAaTTe
847c/5CxNj8Zi8MPRXPxJkYoFf4gTQwAkqv0moVx1F53dL7z9YC42Uct35BbzsqE
2nXHVALTS/ztiZgiSaveqk5CeKPcwoCUCwa9m0l+DamaiwkyACUTNOIU+w8q4lzm
ctma1tzfds+tq6G9d4RbslrNqPvbIMMJ5L9HNJiyJIYDRLsbH3jSLGcSUjflKxUN
F7U6ponHnUF58CZrLNpem5qGuwrh97n9S8odm/hXcj9mGvKzAJiW8TeKBC16xzS+
j52PyiFdmnxUXHNSd2zN0oGFNJV3/tm6kgqr+VPvV/Mj8VzB0pUI7apve3uPJzib
JcCNKq2gQ88lgsMAjKRkscHGQWM0jYHPaibCxJWAcI2Sq+0m1FJNnqbVD+D/0+Zp
j1q2LGj18EEm4c7MIZOB9GNqJf8iRwHcCHuuxfNosQHRUFi6O+JgzJ/WtbxuOcc8
9EU7RbtdrqKiM8k/i9OIm7zAUJ0IJcgjnGUJcme71OYnLt+RDK4bJnONTzslBFUU
phPepeObJrkL520/xsN5iXELYLCEKxnjfBmEusypyuXKCs5TEKjwQy+BESk+nZ7V
iHslr5jU7PuxrcxAN4RJ9KZNH/ruf20sCOMXHu2Iyhc41BoluD5yRWoKBDLr7heu
nsO6mOwsYxTcP18lV+pUO0x4pA29yDqR6sRA1D9w+3acwlCyOQ1z1wYWM+noc5gX
tTINw1LgzoPHECqhyo+jqxoxsnuNYDQH49FF8N57WdQqe6GPL4TN+39iZc15px0x
02FZKi69M4MDVncPuptcw92fTj85tQzvacwKtEP8iPoQ98ehhl2U6VbF5vtPi0XO
+4ynCknphHl/EDuQS8LDr0RLpUp4GLuLV9d3vfDYYOhKpWdZ48ABoWD/41NXgvGB
frgnO/A+ONtNy61aRR4qpMRW1SM0/PDB9ySbSqLgixF7eKcgNHdNPTisJIZO9GaM
pfgMD+U0BnwGEhKx/SmkV+9J7e2lgdcHHE4IqfuR/2U3Ql5btHKg8Y7RQLcmmKe9
1tjx3gRxYAEomx+1wCTcnQCY1yp/I+yOebV+RfNjGiUqEi4fdeIZ53Wlk4XBrNXN
FdtRkpNguOndUt5xphUUO3EO1Qbz38ZbdMCH3AUvA38xlX2wPZu9naT/GmndPlYj
BkNBQBWQBtkshMawwvKag7rX83xOSJJVIQAss1a+dXlm1BxOTkzF0umY8U0M8nGE
tz+AfTNvC3lIIVqOOgXEZYqANRGteSVz6PZUj9SSbGtKhlR/ziW9f0EWjc/vNHDY
WWLJ4/o6QubR4ipOFxVwvuu/ODFwYfpU3mspidUTiEhNlXNxbwpEHWA6RStrLckl
vNr1p1KaX9fD9rkwa1MICjQDHhhbXg2woLa+qemFuDcSEu0yF8FFam7F3Qq0/JlS
wSAvRnbLXzWRLUXtIVRCLKm52DwkJ4W94Tg++v+mkSwKPs+Hn+adJ9N0gEjmxvw8
M9MKyGeXc45G8CcNQQV/Kf7ExK183pHtpH0XJx7TUhHpmysjd7poCPmR08qZnU/p
GzdYwkHuk2l6pJYPMg/XmsDdm8ZGC5e438KfKKj5f48hrMY+em5E/7DWq4dbyrJj
dzL/Bv0+D9ROZIXFgxJL8VJrwZtu/JP7dx+clAct+tg456t/qKq/G+ALGglYz1JN
Nh7FB9stQieQd6yKJtCvwBJqNgpLYirDTAG3QpLxVPv5mXRMPDdQ+Q5bronsbu6+
Ym/GwdQJggwOnqAe0E3kS6WuNcEJaX8I6HFvGB5PlaXdHInkUzdSxG1wtOqpq8Jm
hIpzY70kosvXwSgEs9Zx1l4/ZbbK2nNhgMSA+NNvRPpLI0Zy3dg4jd+UTUDC+5nN
YuqxYJwmqRHAeq/F5SBfl8LDCzTyaq/L3cmT4GP3EC08XHbesOKuJSMFybUi4NsD
8KI+cSw2n2EfDhjVfXKaiXSgJURIGKbHo01ZZ5ysBcNWb+9IICWX6CoqQAxoziht
8arl4whMUe7F6yt/q/rjhAky6vQLWqUH2+KP0LGmasuFKZ9HUvDmEUITjFEhWSud
CPioOQ+hVuum2aDUVlUkmOI1aSu1fTeEV4MwS3FpLGoNgtd4j5Trp3fYKrYuzXMs
AFjG+D3A2EU2PX/AlfengMrUIOi2bznlp1MrUvnuqzhGDiDmlZa6IC617oDdKJVs
tuetLr/w8acS11zGb3VQrByMN09uc60wM99zRcFubpo4LnMraERL6zAlrOf54eTa
WDlnaXEN1H8wTNbnH5RAmj+asxOH1VHhr5wgSWAQvZn+sGVkJSpJNsGLF8VgM/Ia
+6+T0hYdFyegwGjICylMJZ8cpgKTQhUYbFIDiNvCyWKpo/OUhr+262LgG7VedzCI
LSEjNnMfU3bYhEpGHz2SBSjXr0YMMhVF30hLyW5YtKy7GP/BB3Nj0ieR5v8Fqq7y
8W75sbxTJIZtA9KhGpUjC88+1iBQqwRJzFFx+HNwfcanmDzFLfis7WVwxgFSkWDz
nSsU8gBb5cyVut/s6nsFNwBMM/Dv1Ww+x8oGWXv/rw5HG72Qz33vJwlq9a3DF4hV
h9ok9PuG79QiXmt6m5vfnBH/YABtBlxUQPEdW+z52yoL4eGPf4lp0OHT5eCLmybG
PoNQhNAPFaHqCSHKx1MWd0BiXIAzUD9Gc5Ku3I3dolN97GaA8Tq1XRVjrCJo4Mn7
NH8reyjFKeEdx0nHAgrOu3fMoYm+RXx93/fcexWNEDXaWA2ClRyIDsZHNlENZbwt
wVFHWJI3tnF6Xlar5cAKbhJMNqf/UfbYChqC/FcdLWyRns0TVPTHsJ3FGO2+FW3J
gSLmN11RU3C2BIMz08YpzmlFP9GazdYV6clfzvT9zTGgbf1dt7UFR2vN14q9wEU9
v7WIqnXhgpVbYHkRagh5oWBhaeGVFYCMxPg2wt+mY/I0aCJtFft5Sudk8up6N8D8
Hp7yqyQG66PhaB3fWJkpPqtHUoesIfaip6EUzHJNAdhkT0xfuJzjFza5OwXQHrET
4p/VywLx6efW834O40Uc40C1A7vVrrlgux2DaZmAmuskyaTjNY/1HpZorONZjfYV
EKWlWw/LNmdi886j3KmwtHKmyPCX4LAuSeixf8ngSYz6QH/qZxPoVchu2Aqx30uV
fFsf+WzCzZk7KRUtHLTqLHtQdRveJGJMtcd5pHx6g5eOdLV03HsNalBezsgR80vh
s0m+j/skKabA2YrqbwG2HSfTXTnEcKUo6i8ppfoVeJ0Dln8AvctghtFJD/M8tFB+
4LXC1jbL4v/zLw9ov81WZI37hMFcXmgJaeQ0XoOr6K74vgt7CEaavRsPcTH0G5un
4bjzU9l/DbnFMmvhKM8nu96ZcKHG4ZtMfdGPd5liPzY5TLqnWNZQbDEkG937BjvE
jBY2ct9ebC+PYNwbIJ3WoUIdEHa/OyingPhUn0r10pHo6Lr148w7S+0Ss4Yo2iyP
JVvyCueSULkMZRPVjSm7i2aQ9jK+ulNrNwFjd8p5fS90OrVYw+YSLP8nJbrS6xY6
jBz8ztnrd+WxhxzC1NPBH9CD5N1HIpCQIIVCwDWkkmyJ6T/hPZWVoNA2oFW5RhAu
oOqYFfDmivZnA/6wdLkuCO+fRfahcoIIjsZaY711GdzSFwV18Ew2Jj1IDN8QVDLP
AhveyqmC5Jn7CHiwBK/1QrhCgRbgadV54n2brdU9LGuoB8oumP7X7ikBoxppd9MW
IYm4nudGb7ZkBKCkG7W8LJun5h2kMoFq8swfYoVr2EUz2rjZTkkF46uu81sl6AFP
M6kAcXK+rVmXem2bCeyK/iJEoPOkkOEkpcy4jLbmVRtdpHop9VSyAkx5apox9MoR
jnOoWyt4HtG0Fs9WoH8dWyI6lHTfCyXlCyVcj7JzMhypl03aCMxwIjjRowR4lulV
rjDfLYV0FbuFvNJzHZz0uFFUUc5NRx3nzRe/w0AD0QaUoTpQYoH4aJ1OtTTlcWt4
1KtYHEz9nwAVSphLf8vQX5W/+pNXiz2k5+iIKZN+dpXQifTS6lVTqiP8IolZUL1J
oFEktuYjdDiHakKLNpgfeojD7dVEPpXyBBnGvK8hVfI2LBwik4oARM84noICZPf9
8esxQsnIiKlSQ11AxfjAV2ODwBAeZ90IdvHqzT9zYhF9omfmMwPjMsworaIpvlqw
/mrV2CbZttEcrzjZZZhKl1nNGcm6/9Yet7NUvVTi3Ldtiw1VHhAQevyaWnLW2s1C
y6fNnN0xkNqFzk0Eof6co5d+t0Tz9DO4mTwY+K1BRQm9msShmQYGAnDtXyXyLDmL
ne2a8nFnYohRBfVWLeQ7Qb80IhLN4koT1GBomLvHOOG9ixjHAJ5X2zoQwZYcjazo
UWkLIRNbadhZlI6J6rBYv6R7m83PhNBCWMUR6nPKZXwWKMDw6n1LhnC+RTH2cyup
FM5W8A5FiWm73rycia45VDOIrjBrzvYKpttLKepfRL0Wo8KJdMWdmYEHbwha44kK
+3/AB9H4WRTOr8qF8gvva9rplpdVnU1tNLIkgiDLSi6J9qCWqr1tERUqIxP3hbhX
LcC6Qs0P3vbwbDw2Iuan4T3Q0UfioL+BxDbZjCbdhj02T+mRjrEG454JfLpgx6cl
gfoPwjVOOJb7T29XOQyCE3+r3rZ9CxPBoynCOvJvksuQ0OR/Lb+5rdOvbTx+LzNS
XQFxiGeaLdVyO3JgqIbqpyVwCKtvN/g0WGj90OhqWBcmKWD3VH+2P1ECi4GL/epg
hAg1Ee8rBrZQp/TA+Lp+Xrw9GqBkQnaXaiwm4IBMTniFojU/VR9lw5JFNaG3mWPf
3XgtH4/qsuM5MstHbjbC85YbWfKxkpXUhEo42Pp4X2X9W757IN+hiucsAY2MkwjT
gTYJnQiNFeUA18auHayObYdMnKnMh41E8n1rcmINyE5Gh5I6avbW1W0lVMdcFHVT
IvAAg0D5+rUfkJy6GIqyzYm9HNhZVq2Aq2VGUu0b1evhFWzOawAbTGKvnAZHTv7P
VTrtVNTCQ+VBDg/OKX43aDZB+GPWVY0GKH/DTLirDaHlQSD6pMMi4amqQlA9f88h
jfmNFznTlFlZ7a1wE2SBXhLcey7HupWJnPcQ92bCJSfDNRMkVan9bddsgkJiDhqr
yx2XX4l3x6m6xtd8QgXWBSjuP6PwwSMwCwQmQ3EkHc8PCSYO8ohFvb8huzIcXo29
L+B+FMxnC/D07wufFb+T2KveKmGNoAQg+q8HWy6M3KGjHri85YphjzNC1AEyVCmw
vAmJJ6NlJR458Bl3gUQPreMeZv0ebeRrJ3ZKo1SPxJc=
`protect END_PROTECTED
