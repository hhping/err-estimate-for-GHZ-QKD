`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gixe/kBXTfl7cgO5+Ol8XQ0TU+6+Lc8j4B3FNYoW3N2pHrhu6GDqfI294i4zdlp3
wQrUFcDPqNJEwGZvxBBHEHxqWBGXuqd/+P7Gal0a73dAUPy1hYtC7YBk+vFBU9uJ
R0AKpc4ecDhupgFzwiN5FwlJE6aZHsT3V1/JqTLvOkvZ7XHp7deAuUi2GZwn5R8u
uquAtVeGaKQ1U9nIyEOHUNQ6b9f4F32cTPmsy0uCM2WfyEzGNrs4NT/ySBh+Pv1v
gqPFTlPCYwtvAhtU7dVPjxuE0gBueWOR7spe8sDzEpve+EFekNT1OkZOnh8fmRqS
hqof9muxukGqjCbvNouOvULJ5olguY+yybhHr/xQTr9PhItnLFHLrYnyIVnG4lmg
Q1UbhPqSgpIdJFVCeQJCLejl7YohFfqubWoYomtxtBXTMXxuvk9Qys5rRQojf0+R
lmRW40DSyVW4+UXq+pXsxbaYX7X7ti2RiLW2grB0UwX2iRDTCZts6ai3/jD1b7IF
GnReikAjvPlTzHhsJ28jUDeQU8C5rlkWthmVvR1Y9N/rn15zAkv9U33qnHBKZ7Po
NmNWmo3wGgZdrSXPJL49BTKPsiOgS5uRZBgQWkCfuXrfQZ3MjbnvSVMHz3PU0Eta
GKLOq/OBk/p95SU4laXFrmilfW9bPcIs7I17MsUQ+ndRp4eWkCjgqlI/HYJzI+iM
cGFXrG4Wvog6Hujm/8zo63dl+3bgiogl6lTEFZ2+7GJ79M0x5WBN3PaSXycGZ9lX
xz/wyUwrNeiCr2/U5cTnMybDd24HZFcudZFGRnQzK/ptWPkgGJ3IPhUjN8SEXQEQ
xvolIHCy1Bmi02FxqZ1I6niR1DkD/rQcAmtSya96IAos62t1/zOgQ+hAaScvhSDw
aH5rwOjQVPT7zL0I0s69DFBkpzXg1oZEh5p4NCTLy7/Hv+9gLd43eEgcJG14KTVJ
ApK/RGTmJpryEnYi05rg9ecl6viiHk8K/jML3gC0u5k+P2SgR+7wWL4NIUpC0JPv
r8Dt7t4B0uMEeR3CBmCo3vhX9GnaYEJu6yKw5FCGol2YJGIUayJOciw0gb5JcNBJ
U9s/lVok/jHL58lOVssvPGjQGGqgV3MZMAGzk6sM+ETk854Gq4cxYjyC0x/7LSsh
9wWBDKdpzEvsQ+i5p3ewakSYemCvvwyL06EDsiDuMAHAb7DySYmTDqt1DIaol4BH
J2Yemr4Hz+n9bFV7BzyvZYGUhT4OQjvr/RyQ/vp42QEN0yMO+mFuTTSggPQGoOMn
0skszDYm9YH/IsDc8MnMIS7CJfDJRuVUcZu4vB1wuBJu0EYBthvuYMf73JPonefP
AEBX2/AYqIUkKw04yI3QWqFjJ5hLe5gqnExGTRCl2QUoKguqK0wA0I6pVLbFhZOR
aasfSM4+F7Ghy8MjayYZw+G8ZvrGlaX9BnUGs8lyYv+Iux3g4m6m+qxOazlRbHR9
fJQF9/2dSXGcsk5ZOanDKeodFM2XLnuc8Ml6sOM3FBxiKbDo8+DqlYUS1INLnLk3
nDK/nsEvsjmNpmivPyEl5tXUQorBdDjmDIM4GgRlBhdzgxbUmjkzGoSs7F3b7V2P
4K85YTTHYrye1OWBtfFsCzFkMUHboCIzXVC8fAVU2mFv5miOR1UYto8tahMr25Di
qhD2/sc+sLwwciTUfLpS9jVNCYJTZdEAjiXK7zdoElsqu07ec6aYjurucsqo/Cjc
slugCcF0GqpxJwwp+D5xKOiuOm8iPDeSz49q/a/iB/6DPFANT1VWRqsbCzT/qasG
YLsy1NEq1bJq6tIDTBXUOT+1GFiUhZCGdFk2bIO+/CdWwX+OyNzILsaTlEzl2NFX
x6MZv0yoYabRNNK/hq8vk0k7ugLPqOhmAQhToGLvLAk/ezKIRzwrznaILaccvbRn
ZLlX1QI+x93VLqkJ4ZdZxtjfFDM9Y66bmepkpq6wuA59zyvKngBCGlTtMMlDkG0/
6+NQeFSr+z3U//y0bS7rfkNsaaYk3kH1Vh/aYVdcDxhT1xGvS0ZdmHEE4lSCopft
K2CmO2MQ6SfgliuHzjxV3zwy2oXT5NNtr+wFx2LcACYGnFp28fjgOjSE4AqC2I03
C4FaXVRbw8vI7PHp+on3CFN3HhJe3N7Qe4FdVmvImTeec10IXgpw3/412rVYnC6s
UpS5+kwSXiw1bXyEok7Lh3wwcFRf8YEnecAzvBUeqebYh2vvBWM8PioERvLTtoCD
ha7c2LUjNmSnOvJ24nbB7iTgsPBbFWElRU42AAqRJ2fohAQc/UB6Iiaw/jIQWO1k
0RzhJmheEur8VunZAonOe/7nBb2eKOmtZrdSSBHzj6tBsVAqfXNlaKDxDTS390sx
3yfsmLZ4y192MuSURe8YYhnUdYyxPTkBAhurCOaafFiVu8YwaEveeE/GNPYteD85
6rDvJFPWIBrSawNf9+SQ2rnuP83eF4cXS7LR0hNlgobogvnWdz154hAszI6M8PDf
7YBPxQoNZLXzX+9SPsaieiIhXgYxW/sFM8nWvElyy1VO0C1Fj0b5M5Jnk6L9GNZJ
AL4VVn47ONHhddHhwH+8F/wfVtUcsgWrnHgVuMjtjYfKsSAc9fIkyirapGfq6GsL
EtjRLlpyh7ypaf0IMzxyxxc4/RU+NEl9g/yxWxmXRjY9f4a9srmhol0is4tWGdcX
GAbc/EDmAZM2V+D8NKL7qyZND5rE9lKdtEngWO/Ff5py0N1y7Vr3BBDVwbPprYC7
7ISva/EH7onkYO3ALvxKcdm5THisQ/r0ddx+raN11W5WhPcGZApAJ/2sSB71eCPl
Soc0iH1eNDC/XcQbY4D+IEZ+c6nt4DFdi9o9Yo++ECdGYZIhCBrb/9GoS2RqnPxS
1vVy+TVKMhzs6ADAe3TdGBGZWulqBqKQ8KaOsZVXoYQTO0yWpDGXIP2U31kw4OIi
eUpzr942iB5nnaWQ4LbNgBSaPl7gav14f9rHmEDqdBN3Xtp62/gyShYXtOBk8bpA
80yPgDhxVKuQBogKl1a9Od8JE8tdfvZkJOb8b/dmO1ZvnNfY8A2+dD5WlAnbgzzI
vCsTGeNyYaiTOcCFlW3gNoEPJxx6TBYVQc2ifM1mjr8HxSL1z2J3uh6rkqTukoLT
Df1WiYDcUGCtIKYodcNTj54YgEHSejLUA75LE+NFIBgEkmnshhC1Pb0TNg0YgIvC
w9nDGKUusuWslMDUebxq3opU8VnEX40aGq5XGZ3/IK/GfKZnEXmlXfXWoE63jleO
akbyWyoXi1laIZXU9qzB2Y8k3ckK/PLzzPzS72i+zdR/5kKuvpoMcGie5kMiqHVz
OTWlR8wkN5tNGHaPP+LZ2f54Gn8JXyd+JRqFohiWfi2a4KT5gmTUtIH+e9SmcPLB
X/er3xeb4iVshYiKVRIzWaYGrKRJdSx7D+rMBZoN9RlO4/+VRWBdd0bYBWuMFdUj
RI8yaZ4n+EK93Ql2CSTpNv4GM7NPwR+CS71sz15t9CjUEr0jkCqN6fHATj24Y5a6
XhlA0pzLhL7Y1rPsc4sUnIlbRy0owcbuSUq9wi8YJO+yNGaCCSF7C/5BXwO+PUE0
VaK+8ym0BKDf637fxa/NTL5TwgtGhyPVCT8sdtqneHW5Ers9ZdrVv4YoQQZ/h6mN
8AGq7rCWoyce2ypAHla/z61EPb/HXvorrof9rj913dxWZwU0kIK634stdfJ4kZ/I
Hg1+EY3Kph1byOXYN4GF4ErNbKeLnkV/wk060HNCckt4aGQQXpkVyCeN/pWvgHQp
IzmUZrFRfkhOmyx7X3OMBtcHvhItTjCbT5hULkwWHddazbKc54Xpu6TZDeTscebE
ngsxJ5PgiSI6YFg5vBWySkjDbuqCGZS7qU3dZTRLNvGw5F24CaaiTojdPflP2uZX
PCbYUurT2zGFpgukvJQyUBXWSpH5q5escTFeCpiGfa/q/+h4qRN6Eh5WYFNex5ai
H7CSmOAdUlMxN1a0eAhytW/22W1L0Tx98/m8Vz+jxnTipqcB+pGn77jXTj8uRFRp
QNaI8cbBdsYOV/AgZ2Xd+B5i4h78JPJyJxK65VfEL1Ofea4WCeQROdyO9TUrzj4T
H/eY30KvoWJg1f6QJEWc0a72p8kF+BYPhJurLTmPWzI2DU/UIXOiss37znWN6/Sz
9l8KAaZkFm9mZ1RsYTUqJrcmlpRNXaPnIdClXgeDzlrCiTH2Z+iB1y7DN9zlzVyS
xlDxjg6lk1YWXkpnDUQ5SGCeRtolwtiRwDBWdyVHxuzbcy5kTyJlcMG7p0JupLtt
FzBGKV3AXSSKa9DlKi61PDP/GW2jL6eWlytfUnyc2YyhZH4bfa4FkAMPFvr71SIs
S0tX0kHEGqgqcH+Xz8j4Qb2lekuE/uToPdJ2+n/CFXeah7/aJYaQyAwUcYaz4q68
2O+EfHbNoNXkv0lNshLkOGo84HydhwfYf2UtcYrJHtFjGFKptd4e33y+j39bHNMf
+Q5AQZlgOzfRoMvzVQkL090exB5rFm7nlV4GdDr092UwHkDSZJqIg1m7EtshN7SD
TomRkU0lRoYXXq+UAnYXmcX91zXrs+5Y8l6DTBS5+jdHCFTGG5TTb9IXgLFQEfMG
/FO7zW/e1bklWrO3wU0DwmD65dSR93mImR5jut+gpHlm9lk1Weep2TaaJu7Lf4vR
EyA697zkceLyjDbfQYunQKUS6QAeRdLe6GgZ0iDY8skWfxhG5o60nxgtgTtqx5/J
nTR+teyKlssvQz45bSYdxloKG5dwUbybOK9y7xvEir/2A2chmNssGnGpBbuQnePR
QKwKb2FF2axy5nxGor1q1KQoL82Tk7FccLeJqGObThzd4PycZ3jT2F38nhSMJGiw
cFoST9CYWjqqK2BPP/32f44dun9x0nDJne9ZLy+BLras70+CZfhVrtJ/yIw9iEwj
V7mjQgJ78+CaJdhEz3ath7cDKKIf9h3Kn5RQeuNBh36g0EVEJAaKXnD9EK3yq55X
1ATMO/BXgA6Cd69XMAlTsQtmXTizjVQpdRjEP5Bv8s4SLID1rr/Ei/VuENas49oE
pLTlAWkrGyGydVOOZTb92o3mEaDczWDWE5OyxL7MQrCZ5uRMUdSn7lXxOQt1PmUk
eDimumqDwD22T53i1Qviy/wyCsj6omC6MiP8tG2+yAZrr9IujC+/rfe3N6O9G4mn
LWaojKt6If6bpd3VPFsjOswQqrpCfprJUL8aDS1D/sS+tR4VyZ922t0UTBfoLSe1
AmkfGhoNOYorOcz3j+7EF19DJyg3+Gij4Pj3K9Z56S2GPV3xc7IrM8NTsqK5bX42
1+qhCmPf2c+4/6tmKsn0nltaM02np8/dPjYe9xsVpKkGDcX/ViY3zt4BSKumF1qK
qMsCRTbwsFmgw8daXmxyZUK9pkQdklI5e/Rw8HxG67f9OkEl2vyUKK6pmhjkbw+p
Csjy79X1BC+jpiT8UBCmjv+y//EgAPefNcx2Nlt9PJ8BcTlA8QVT5B2veo5m4zSY
9w17+JLTir0RGGoQHG842ma6e8tQeL2mYG/hCRweB1n/TqhqPt7L4iKKD76RASx5
xW4Y/hZueawBfVrPT7Tz9fA/cyJKjEqasCKJXtpOGvACDxi7GMXbQtFl+81N2uJd
gqzVy6BxVNNQ1OLPPEB1plvoVK54T4icpOfWtS+44Ebg0RrK+Asr/6loBoB/bUaP
ZeSGU6SIXpfKonn8u7vENepLWUlnvufJZOvVubqPn+OpQGGJDiD0g4kQLZM/kdu5
1TnX4hpzI1/1I81MWYl5UHkkxdsTOQ6yXlw+bb0CJVfo/9uwKWikkPxtU7x1lY4G
dN0SvgWOEaZvwb6hPP+Ai2kV+Gna03e7eHT5HP5XOoh1OhWYlDUY7vXnAhc9EMqO
5GDZHRbl6Rs/RimbkgZGehy1CTMkw8+XNfi3Gz6dAAx8lSme/uwVm3swteWVo42D
/GoP0h/f38nDOlyFFxGDtu9L+b23sqUCviFwEluz8BY+TmYRn4Ubtn30CtmzawrP
scRwERpPRRwG6N5fFsKHETmYCFaFhpJbjBEjN5nSXzJNRLtxxTAZvAUNOL5/n9Wb
DCMyVHJGWpZmW2XUeTddz49rcKIT4KA6enx7F1LxRspQ+zt3R61rN8rJ7Cnrdbsf
bOQsBZmWPMmRF9n5zABwVEyETHjajfw1sT+FHuIztOqD+MMuYcsLSjviJDO0t7x9
qOTZIpBCM/dRBuPHJXPLnJANNCYRfVRtMbw+CRQkq5esVIJE9AgsyY6H3peaTzOK
9lMfSTpIPdW6OyxPeX+sJRnNnYXeJQTsBaXrqoQ6kDh7skDwvty7dfBHnDwjgQje
1bVVxchejWPF+p/fQ2C3sRppFSaOh/SflNLc9ahEEnCUPP63xNtEwnb6JbogJx2x
oLJFQq+He6oE91Vg/dPhTKY8irt2lfaCs/+c7DyDCoy6rzFCfT23VR9/0YWQpcgE
Cn4OiPBVB+fIAuPefNC/g7GkuzIssDwP3RAOArThvBL3jBjGbAdynZiaKSuwPHl0
6bitZC+3hdSSQl+P+tr9bFHmrsDVcv+Kenf2c9Kz6L+yFWpg4rY/CzYzdCtrHu4u
npUPMNsxw8CQmOstvdUuChv0CeoA6m5TrqNf4OAoCmlI0KoPHrER3n/IKKGlh29V
tQa8qGAew8NJpbvHaBfPfnC4T+Vsv4YI2jEeKA84NG3CjYvOtC+wxSVoF9RFaCDG
83LuLlVS0tMV/btIh0EMczkwvD3zM28htz6GbPeQmEQXjwwxjDsE1iYqbYdF+uOH
BhxPMBsANUwxBUa4e0iT7YulDP6AhUwymZEhU9w9XABnsXIn95uO53cgFdfOR2IY
QYiCrSE6uF9+9pUOgmNkKTro2cV4dMtdXc7gQGcDZVaht05WRvnjABluOu0VOPTe
rege/iE5a76tcJHjTHN2LHPO5O26hFpBI1ZZzpfIyeiFWGWhYI07LL3psjAHklP1
SGOinugINVcbHAThRcK5cwHwq9eS1JJVtWkPPqfbZq9K1TiQxFBDMLFTTiiofQ/N
bHpSDnd2s+GLWOwz1KJgAyJ6d1n2Kwu9PRM0Hc2Qg9GF+PSyv7Cn1TWEkv/vfLMT
vw14WaYBaAOrhI8dtBBh8DuoVbGSHv7b7ZMfu1kn/IXilsxCgXYabc+PjZiUwUtC
UcdChKlAfmdtNaJ6wia6zBpq9Examk3Y4xfNqmc8OUcmJ90nOrsBmgzDG8MkRszp
9Jyug6yNM+xQTODLYmndedLZw8ASyCdgfpU2ntY0vk4M4PtHx1VQj8TsGcBRWQdH
ueYq0JvkVXYe5Eqe0bPPcyG3O5u95hDXMJn7WSrHlQqZ9cS5vDUE5Qbw+S8FH/j3
hw689eAJOXfWnsRe2co7jfv+OgJ7+O65xof5vUtD6TQov8vCD3uPAoR9qEB+RAYY
NWcOObK5uaL3iRYV5X46Wkttlx63/MKUHg8Aj5BMOahCKIVf1eJzFQjyErAal1G7
/wITb/gt64+Vq7sswYCJ4MwiI/FzlAQ2dFYVpeo+iNQLupE/hVbVxLH+CvaaW4cF
dzw/nZLgDom/7kuFCNvkCuhQG6gr731XBqTSJc5JcLVGWvozhGZilfrFmeQf14JA
JEjFj9rwiSgtypjVp8rrpxuFnw3+zwouLG2OOpTuenqeRt7cDQ8N6D7danNiTDq1
ZiT5RO8KaqPrzNeoItXVDaPsrmLYzLqlhqSCKcZjWB2eoCtDxKtOIrwR+3nP39TU
PxkWxcwE5G92A9T7RNm+kMFzYyTDDP9OhTv7goTDaqIsdxKUKCnKJB9XXj1Cimyl
4GQanZhhYu3Jha2XHDbJqoM0+oOzF8fy1q4yoQy3KOECDCSchJGpIEMkReaza5C6
YkzqpMbIj8XarwW3L73zW2t+HwimHY7CxwlcCo63K6jarB1BpW5qH0ldyqEsRJUE
9D5iflHnmNeXzZY6i8brginnGlueHNSBt1+d0XlaKtJms3P4bKy3nTKbQlkYzGCz
AzG3b7dCYb4JJGgvRHmzA7+vUAW3wRLYrOjlcp+mrLAee9/IrP8uru9uXN+Klm63
AlTDfDoj5hP31F2NaqQKEDhuaJ0KOo8+tliw9qf+A1C2+o5lF0bRRhMc6WviP9r8
BxIUQYB1J9/h4O0WmR7lY4xtE4PH99gC705IEHH6w0iqckZat8IhBt8WsktAYMT5
Fcy84/Tj3PilEZ8DePne4TNlqB6D5Bqq1cBTspwOppUnYysChO9dQA++YN1boGux
Gse3zYjEFE0kKJ4tvpekEk/Pnj5xzUHR5yzl6eYL3Y03EFRtShOAe0Dx+59ZdXSy
V9KqndD3A32jkZeBREwx1hPkNwl9GbeUlFQxnzF3SObOJAOgnfsOOgVx9TgtBzn9
mov73AK9cq1OHaIitihz5bvvce6nzPVpThs2BJU2Zr1cYyWS1GFolpQukWtznqFw
iCsnpiSFblOA6ik3jfmQAzuGSaw6NuUi8g3LMToJAFKYWjmkjam19KnnQRmMdz4z
bfq0Sry9tK2594sOVGEPNSK7eNMD95KTu+nwBitpyEUvZ7eZtkLUKQK4M7AQovuw
VDkLG1jFEEW+ioeWVuCCq9bn75hr35qMWzaQMIh82biRJoOk8+5di+n//6vmaS1h
pKxDNIqzjWPfbiNthXPNSs5BE852MKwq8BHx91G8xRjgIa8HXNHOebRq1ztPIIFE
20wPG5Hfi9UMQGVLmUuW2PhRUzhWjyXSFOMHk7A22k1b30H3j6md7IfZek1H6ZTu
eFwcmZDBGeJ0KLO1xwUAzB2rfYlYSRVXjIqcbpRpg72derrzdHpbVublb+QAQ97/
8UnknSn+zjya2rUzMuO1OzdOGpb+PaSxGSu1FSHel0F7ihnR2hhlfSlvFwylqPeq
PrMCJ5aOQ+VB4MvxFuQxEgRTF/lyktjZrr77fT3SrAqE0NmiyaTIRb5GJ+7Cmidf
XGzxkDeGUKr4KwyZRt/sELg0AD3vG3PaBq3ywi0QmuWKNgpYstmpnoBMUrx+sime
sjEbi5WiRZODokgl9Ifr2sHrAe57j5iSYQRTx4knFTDuAz6qIb3M4F2D11rxRaXx
oOBHQjR0+KFyDjypPk3308Me4C7t13jt/Pbs6XNOeGhZoiRVrB0yYPX09R3fW6ft
a5fecXlN5zsIauC5kdgeK4xLap+fdltjzexznIx3x6YVOkw1X8A832B0zOiEyQIh
ZEWupdhPHssdE81NgoKfhvWVIlLymwUpwfxR4R9kbeuLfiyeEFPKMMuIeW3l4khg
uJ9V95NNb1Is/SGPqfNEmpimNMDWFZCLyuEonKvVjRwEm1rL+gm0DTtwWbYOA4D2
Gqu9RQh5ALk9W9a4qOj0Iq6zE3wJ6RZ6Q023iUHyuoQ1UemoEnD+XYU5omDWoQeL
AEZ7FLtD+AgTW7NPoXHMShMo33gJLPQq8Ojif9+7wPn9RtgoWU//hGzT4IDisDVC
x3LUyiUPTASSBnOXsRvxJPvzyHpuzg45U4QkXjuSNxgWC3BszeMXEwb6paNrsFUb
GwI9ick+vUnVvnZt3X4tn+5xNi64bZoe/RYmQPDzx8Q/PUyxwpYte+4TNV9boDLI
39NNQTajLlAYhQIMrZcr+UkVvvgfXGl8SjFQcIAziWdbs4XMPy1fbwzc3vXCRKVt
bhJJMIiCvOJrYVKBjD8GpWDZEmQrPSfa/D+ojchq3h32ZBaV3xq/j3LuRaC6diJO
1MFKNHntYH7nRxMvJGXRk4iN3jxTPAgVATmtc/Ro5BndO0xaKnqndjRc4P+N1qy4
3liwIHVf2juKceH0Y/O9Aik+1LuCQ2wK5GL9HcXnWdfEnuPrsAk1Nu6ij9wOBrko
jdbyTGPuoy9ukHGVGNZJR79w1bfs4iMjtJuGNSE0Kwa61EEyIUKSE7iwdZrB+3pb
fgTuITttPAXRzfGXcgA2rZXMNCsYNYd6QcesFKLv2ByYgIGYIbSzyovM6+zYS9gM
8IdzOXBRmeg6NkA3jUwBNoo1I/UH0R0fLvf5CfD+JqjNcLVU5JLu9EZpmKj8V+Vb
4fRi8n0UyjpVqAP6G0vUAdpliuSV25zRLv0W5iNJUQTR3NKP/5TC31GfhYLxdXlM
eSKqDN+xStUaarRs3jfV4Zgx4zyQnnGDE9IkFi6LGWrwOn4uAlHZaAKaugCrUpTx
HfauvszTP2swoPgTWZlxIRq6B0Ax8WVcnWPRnPg0V/H1LeGid4Iy75h4LDYfJH/3
y6mbTaU+WmCeOVpPZyHhHDPUu0AM7L+UROtPQoTbv3/gdsqluMHmKxtq8PqS4pqS
9OSFNd2URw7OYppOoIcSlj+c5nINuML0V6y2uRrInxAhZx3qmsUTX9EJQedy4vGM
+efjWPhg0dXJKBREcwhehsIBW30ozaSiVANQ8G1sDdWCyszanK7cKvDx1XX0oRKN
pNaPL0EfyPkKeZHXjJe24sA5tWVFKWBIROaE+yCpIJmbLnJJJwuFyWx6pR+OxO3M
t1iS/zVdyG4eW/Fkqs3hH1LVBUzoPPeRR8QeMyzk4cJdO4oMjEewr1F3SOMDu13x
QD9duNHnQX7CMm3ToNgKhLztQochFWECSpalUtss5au8tO/Pb1wBpoAaYh0KQ8Rw
Ht8RnKnJ/oi/KAV5AMTkp3W/ZH2LiRm7OTkbChpEiDnBmhiIHDqXTdf9FvG8aQ1g
nBVz4frM1ablOYB5LZAI4nTVTjvRJfPJ68pl6IRJJtjljPRcR6XVjozAE+eRCB2h
vKitW23qMLCd1QQVVBLLwQ7T7iAuzoCZmK833S3kENlgL382bgNLsvWcZQN8M6gT
jIRPjjhnJCtjaBcHWnAjCNJFoimR+28JM522x1+TihwOcurZsQMHgVK+pQVoW5G7
XkjXA8doTUgOYfVCgGlUrKCLpNUN6sOszcTiAY9f85f58z5c2v03q4IYxpgZl5yK
Tccq/AyrDgTAfN4D5vVNjXTHpUbQ3Cl/7R9ioG+5tHI5Mm7yKoqVziQY/hfj5SPE
p8xaGaH1I1o93ozSPM8a+W25UDhT7/zK9mQOMX8S+VItw47v4zszN/6aHf/0Ovbs
kFNTn6QT8ms0w73wPIHjOvNIhW8wJtjSYm0rA2+dcpuKixIF4DNtRV+g/QEkoIV3
A5KiEyhhRYcQGPRRMob8hu2JknvBgGjNhD6ODRtorn15pDfwdaq+ZzmbMaLD9fvq
FQSHX+gHG2JX+7XD6YTJsCbLH4e/E7cjXyqVYVINWPsm0GmVCU1hEvOptl2OLChN
7MJQPD1ipATKx4AFvRw2zM+NDit7J1iwSrBQwsfJcXuMy6D4tUfWgIAJwH/JpVkN
QsxBb3+tUVAu+VD3bTJKMS2ZZKrtFlsTyprzJDF6w95NM492jHNCVf7AiHL9LGN3
dtt43VTLDc1H8kAAziC81ETzicBeRsx+8LETEIFJUHVGuWBWx/CTWnoEXe7rzM1q
G7uZwuzJznpcklX+riYM80o5PSALFsskTWtRC9d9fKfqtNajmKxa1PcpPFMLMb9a
biYgyI7thdX1S41QFn6pJGhC2He7Ft+OIkEGzSHKCUPlpCVTsEMQtl4cN21vOLo+
VOAAVIT7mgJsI/eIsdBGutKSxjbhgyPXbp/SRULO2ZXPQNv4jAFoI405x1Hqjnlm
UaMgO8pk7zBjrL8HAREVw1GmACFqRneOT348dKFw630RJJAnwzqDLDLBMR0lwO4Z
fjhl8gRk3I0+eLSkhtO3jWT7tkeoZMGTBQgHJo0UAzzdX676JjrgmTjPGveAXuqB
tUXYvySrBGiBqPEsIX/6GQTBehtZTtN1dzFH+6MVwwdpCOkQttcRM9tjaaU9/xHM
fPODrTyC3VSBGCv/JWZ44jydyDtFZZzqOfkj5TD8gRPhJzw/R/ur/YWVIlnw6AWU
2RwMbtEW5qvj4NrCIb3xzYHu/iXgY600QFcHsgXL+uGPDgM838gphwiJWEji83ie
C5QzjlYOF9cG8M6kzUVAG+ZELw3c78ft8kQhwnOEhKHjF14NteaqrdIxVTaSIr6z
QMC6EeoRr5k5YjVzjnZluXPLAvYzHh8YNLe7zaKFetzLEpfZlI49Q6vsxITLwvZ2
k/pXqoe6GCOa2TEHbmwu+KuYD81kVueW809WNQKUqVDJAAsGtRdqzklhuoBnpka9
zFurLhucsgHW9KqY8jCvc/Xf/8hfgZQl+rbw15zVhTFiARGqQt3cD7C3cvGzXZFj
a2gL1FfTHRmfMSrTR1WhkUKj9B85AhEpPlGKKhdWpUJsWxvLTVd7VTC3f6LZlTWF
whNxU8ZqI3amvj3YSz+XNAdFoqmdWDU1bJyR+XVIkNBhLifu7iqjXCTi2+yLKPD3
+iSu7rAs/qvBgedWsaYooEAhLLG+oqendjk8cy8RrrlhYNdPe9r8iiR0LLxcFrcS
Cw2CPOlabPuSMyLPJHrfRjh1fJjT0bczAmqmQGaBD3UqsIFO4O44XX2JpuAEysty
G4zwqCuxlMMsEXYe0UWwwbLT2on7RB4tG3jxkKfQrGZDa74GZLxqHs7LyktVxspu
03OnayeV7qsobqV9HLS0cL/5LcNbgmAqqERREnl7Oft7/zEt0edf5obdPZdR8H6j
rbVke+JoAq9ZK9pPL+JDFlBD5f8FB72789ggKosQvX3sowQYCudTl9dGSry7aZ+1
4reyWz/W66pSXjUpCJ2qhM8r88pEAhDbJWB6GUD8lMg9mz9AUY6+aOVm1Xiksq/g
II2qVh4sI+tUKMTsph/NGUGlYI860QzeI+3mk+5AmiwJsqxR2kRs8gTPSGHf/rnS
P6SKWxWpft/p9vAcbD4KVIPtg6IS2FxJ5kqETZaYWocHS6WjUzuH/I2xFFXe3xda
IDryLpCUB4BEswBmY4+voW60O/TF4e17tW/8V3/UKKX8yuKKqf7C0oak1Y+LD9Sq
Ranh8MMpETU6Tl6w4qeonns1YeEddTe3dxqDvpS14b6GUbmQ1Sj7KlZRasJ9RgZs
WmlJApCUIMIzTop6TheY9Ocb9uRJITLDREFUTSblxCr+LzH1WSitYFb0lYduWKKM
LCKVmBBCuL1TQGwE+LhPzI1En+trdGSNNwFFcMCpJQ0w2sgIehVZBIEs000O8dvj
Z0sWFYk4xZgH0SVB8K+9xN0pE8VfOE6Ozn+k6w8gbSDQSwgIhXTftLrAxxz1ExV9
lFi5tdYu750L98qol6mH4HA9yJDqCOWIgTc8O9IYNtCkVnIQRTCEWFIo05x8YgNo
swYTVUzHBDmLPmAHnHDxYFCJZCl1nNXfsB8RVltdaFLZ/hW8Rs+5v3C0UI5GJd/H
JVmjhv16ag4BQA85+q8n29Sz/ljtSdWx+F1oS5aWxTgPUlxADGlBusN3dGkg3uZn
qKbHuadkeZGXGS5L8HvVlS8VRM9rY1LnPDhuEd7Yp9/hqi/gll3wjSm5TcpWRQie
n9Ry4yawLMRvwH0QJheB4FfjOcLwnSVRgwMROBy53SnmX19WgcAx2ofAKeE+yRgt
9S4fO12BMSPZsHYE5GrUZm5X1qg9wBtopRI49XSz1z8Wk3Z61l70vmxJSiM38esp
h4b7ym7/U1w19uSYtZ4dZoSUzoaZc2FzjaJ7/Zlzl90c78YsZoTkckeZ3ywR2CmW
H3mywJDIVQsNBli4dTHuEJAYc2fNA64RJhlGbQkeadlfrF3g6p82kczEYQUlza+4
12xG+ulD9trap1hNXymvPDLGZV8KHealZeJn5Dnzc9FGbeqZHPB+6HYtsBVPN81q
RjFCMQxRdCrTqV7fSjHlZhkUc3MylcAhCll5qqFDkdeFeg2xBRXw9L4XQsZLnPc9
TFTOD7jYsl+hqPjzXqdCIWE5dZ30C2m8YOclceHUVBs1gxLsNc/wqWH3o8IJOmvs
z0dY/mSLsFZQYXQfm60ZvJo29CGkULpD8pQeeFxxvdxTrLYkL9E2OW0qYb1e+9cJ
a2luMTjTLCzJN8pfRFUkqyB+2cPY0ldL1bR4WE+h4U5zvtVh2xyETifaITpRGxmv
6Lx0b0hrRFqTmdIB2hVgdStpPKz1ZYyBb9g5lM01l8f2Ba1oebWAZ+pApnamabCs
WXo5klP91vCCHl3vAerlYu5+EF3lZGY8f/3jxHeGVaDUfVmY9QB7n8147VkK1cLa
c35/1IRXQn6qS1zeE9W9oumVzVYbpFRamuaXWPkKh0hXcXo/K1xoSv5AyNOe2RQM
GaX/GApU5ne/tRZGGLjl6XwLRsmjE+DRJWeaNplugO91OH0QxKlelfAPp4rNtczP
KKl2DrqhjQqeZwPtcBTcFEkBtkCzoWaH31/0EAf9yVYuvetrsx2V2j+hcEoLIQl6
+f1MZR+4yeH0YFTARm5Xa3eg6EBCh9RJJ+XTruvvLer8sGsq7GTcNZYt+s4NpVrh
lyImLnMaYdKP7RVIhGC613riLYk8y+WVRGS38IEu8+jwSye0EcmjLtgi1faWSTzP
UZJa4sxI4bt1kOPlPOcp7N9UWsiF/ZZ6BO3nRgCIVEtvAU+8cZaJ+h3sEWjclSIC
uMyeNtM0etwgh6ZpjzMGxh4zQK0zcgg0D9rd1OFallfGMCWwPboEjwN2+CGgEh4P
HKkhF9JMhEhelooQsyc6drluAwepzRARmJyYkfM58Ds0GAMnhYIAIIn38IY4GmH4
cjc2fmLUShX4VlVuHNz/L1WixzQIVcQDKxbbHZ3LQI9lN8XOkly5H6z/5YQTyUJA
N1n+osHuyYvI7t+xZhTvNEibxpaVl0o3BogFzIJoIfDo0PkxF7e4daw0VC7IYuX1
EP/MajBKqG7RQPaWbh+F5aguCojFgcGbsLCZGXgahODPHqRzkfPiEBJoyU6uSx+h
1K3BqJ9zW0jros4Os6L1zpjsw3QfeIQf9KSFUA3BwG9GnrmlWfkKbN36Q0ReCMV/
SIfTCAcUX9JVq/JQyodbU6VoMPNDm+Jrm14pY2pd/+O/xMABap61qTZpwkOfyJwK
b/iAQathU8460Q/T7jofkpRKKVxwshtmItOD9FBqTS5UePIK/L+dF/MY8eRFGIqP
Mdlk1wXXfX0PDEpd1ZebmZ4qQBHeJumRNlnW/2YHeLFhBGpXmaQlSLVG3sGAQCCK
KFBpM1gzUD1gPAvU3xfYyxARaH2Kh5aBI8gRoPw9cO8vFC15OgzBebNeDCVzTagn
mvnBEsq0VBWtxDaEU0Z55z9sODXoUh26ms18V/mlXSg6s1Oiy6rPjiflK06SoI9U
m+eE9rC32hugYvUyg0KyuDE63S+jqQAfoyVX2ljJAQevm3PV5bGHxU2gomJiAgWI
oKAKIMRk6Cx0SPL70nDkTU3IDH0yMQaB0AZSxM/jg3hpNKrC8PPHknh5SsEFFbsL
ZVHLzKlSBFwYgb4HUyjq0sAooPeLJOJ1G6KvbZJnU5Qhg7JRedaK7oTB9fHKLsAy
PIlSsZvZxlJr2K2BAjdgNxPxHcPrXOX8uswFwIeDGEsU4RjGGaiGsCCbRv954UKG
4AiVQ0P8zFilJDA2wzMjPYaP7di4F2L6/QeJ7GvdATKX0UUk33F+XxZ/RILO4B5m
8DI52lqgwNH6pbIsjkXMjt7KUt1e8jkOL4+FdXStC4UciY9wOkonTM3VJQZ5Hrvh
lIoFvaHkPsy9Q5LQWK5uB9Sq7BU+yG67+LDeUD1Ks7jZVIeY3b3Gpfy+mvwT1qkO
ta0bMWM5cm4RMXsaD38QPQkNgkv5I1ARlA1gWiNXWc1kFwxLrvjfa8hmOPDncbxr
Np6B72W0MClqlIOIZwai4BUUlSdZE4Icjfr6vTZL8pP4TAvHn+MOW2PIi26cHAT5
3jBTzCw9wYXI+NbjWTKmOHsJs0988xyBfc8DycsG5TiO5VVX70mR0EFRGaKEEvF/
EQyxP7Nr/F3yKyWXNLPuzfeKRgDm+za0BOpCi0eMPPj2b0obb/X7TU0lZy5dbOqE
c5f88flg83YLDJr3gWbN8R6K399C8KP9K+0HlGBba/5OovTLVRW+Qysse6lsYZUa
3fdtGNKD0jMS5klA8IfFei8bADZ20Z/fk/7WJkHcX3H2CtgBlfOtFPTtGRekw+ou
wUZmAzYl7LcUueohefxfrm4Lwmzob1EpgH0ju8zYLEuwsIoBfG1Blk3Gypd64Q1D
TE2wgoVkDiloDQOHvta4tLFysW/ro9QKKMvHu2D+mc6EwlZ86O7C9CLz4NzEha2K
mk+fCkd4C9P6Vtb7UyIGTmsrzSV0MFIB6CYmSPv/oEKqZuu7RccL4iE0bL/VNnvh
TtntGgsa8YzcjRupG6mVm2n/OFUcMr3NFtVqqps9Twc=
`protect END_PROTECTED
