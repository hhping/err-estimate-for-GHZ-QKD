`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9n9CJ0ZVP1Hr88/dA5sDEor5FWeJbH4Z80egIulxpvnt7RjoEpuKeQTJGN5343S1
QiQfUZlwTnurnG+A3tGNrMXkhmB2J3gv2++12inMOK1YzzeE/yBDA3qlgCHj8RtU
mC7Wm/a2ToD4fjzRQXpoBex+WpgtnjKvKWgLL//D6cSHfmcO+oAHilz4GIa1Lr15
4ZVw574c5pgY613jvWfGka/u9pjN+9kF1WITUtWGsCLKPONbvax9SFDOiI9rOWqX
CJS9yG1FaBTGzT7eALaIE8S1+wzlhBEYzeckXnjtlyHK1HF/ggukakcaa2PVGBvf
PlAZxMenByxmxce0h+0SF7UdvbhWUgVU2ZyNXYwDinbMl+pYnsexC+vsQ9Oqkt41
sArI7uY382BaTeRQPR0pelWM3v46Y7PgtD1c9KSBhfsmpbTT86mAOEn76HmVZKS2
/gOZoJhB/nb14LqE/WCyW5DgxiTH+/trcJViRaDxhjxbD1K/v2kgACxMAWC4DQWZ
dTjVDmZytH9cn6XtzJEINvdLBVwltdPRvUDzXArlaTQHRJA1WQz3yrB70m3iuLk3
SoMr66skau5pnwwrmf3GCTQyAbpnLtOAHW8B9WuDsRd48a6DjRa+7+ml6rGjbu8Z
VjdeueAy1tjRRrn4ZyI0XVY72tmwmbm0g6A2zk3f+2SadY+QjwxYrhpYyJmxoLdF
Xwc5Jo7fAVDTDGnmc8URNVOmrWipFYMvl+O7WP1dWffOKk1mCO+KCdkaGiNsBR+A
e6r8ctxUhv7xxn3HmRUwcBnThg5/XnMdrq0aQqcO03Jx2wrEd1EWQI9wX5p54Kpc
yydHPuypigXSQTgOgAZCAlIPU3nsDG7XGusVgrfT6EWaU+kWbShblcK3IqEOuBNT
JPxyLzEXUw6kDoW1C2gvN56ujslTnhCI11TRdZMO/9Ee3GW82tGUyjLmQJX78MXx
rXhbOq3+SsRZzwcjHBmfJPcXnayWx9Q28e1PWvmyUNlHTzLNRakttoTJasavkbg/
Gp54Ri7ZALag7ur5iUXgg3eH3oGtFQQWEmb7TeX8SpHJ0kQ4hR4bCUJoKqPq0Wmg
xUvEdFmXv/st2VwVzS0WU2fG00Imp6P/YD11Ag5Ry0uQuxsZ8Td7RGCqELLOwUwg
TudVi5UiJF47X3EbOKYfEqtkyDvXtih83TPxwXkoPzNQD9OBHHNjnIP7GPHdJyXZ
tNLAUK5NVkhPwG8falds2xD9MV65Uwg5ujO8VzWl0Dje/+iy0tZcJA3eoZeoqdyD
TdYx3TtiabtuMgZBBBDoRbLD6BnuqskmCCh4GVLaEeY3poW3LDuxGn2TZ0CqM3OF
FX0sHnQNPIeNE4daGGVpXbFOfBfoVquHhZzlwrntUxspd89c2C9JyzksGlYZu9HV
kN6FgcP0ntVtX+ONMdaeak/nktXFZrkBdplaiNaZqcNV/Ze2+GJZrP4LwTybB0cj
JNdoAREVEQWn9B9KQ/03KC4fLZulwdEiwG3mME3ODhjAKPB6C3fhlMjNHqqE/RK1
3fHxmTpclTxkgbhmfskdUcru5sGzUnMXzKE6JNMpmSrPW6qgT3dkE2K1j6/7SHNk
Iv3jDSDnmCuOwwDrUkCsGxj7+vxRjHLBO5IhsU9FK32xR8GtUKPic1uLiES5fCBJ
a9ZLaop/kxeehGKYcBNYf2anqocZnAfCryUd9sAmU41P/nrckdlhfKkb0WaxjLcu
TmDul6N9lHgrbvsrJRMf2KyBvLH6cLuKfVfO55XfugaoFKrqrdIgkG1IwJg8ZHK3
v7QZ3MS1fTzCTWUCzD1mFVy5mZMPELPO8It7tdBRxqiGbCW/wX/JKckuYmx4xPpS
3E0ZZVBUQa6hs63MNlUgmlu02tC4+xrgs9+qonk2KzwuXhc3R892+3s4UEvQpP+l
3VlbFShK14FyiRkgLxnLD8eLstXNFnDA1aW0HYoZWkTXJ6un4ogC7YFEZr4AYVo0
savt5JBbYKlmbgtjWXtm9Gbm7gNzPRW3KfDmPGCW5b2ivJaxkNfGqdqPHfqxad0I
RPIiNHLfw+DayLgrkwE4uBuz6RgzuOBx7CWMaVtyBvrib93uvqM8k6xv6gXKv5A7
K3ud1DG63Puwbc1QP7mxzKTEDwx0lLzIOznjZrdpG7ugh5qQp4jXlLiFuHeeT9XZ
BKpDaJNry0M5zfiZ5DAHgI6DXVYO23dd4piGs9o1rjmWBE9+bN1ev9N1ZsiDYNBb
sZ2rF2yMCK9zYmuni1oFqfV8mwZJt4PtlJTwoQNZw80y7HNA7sWYaD/hENVVGKq1
vs+NS5rAKZATrDKDZVWQYDD6Jb6yjz7g89HiYEZBTUUgm7AH4QBbarj4yC5ytxf6
4pCuStS1RtypzZg6h4K6C0qmksAgtaX4m1pge+ApfDqdHFPPr1XEICFpxLg+5j+V
irpgiE6I3/blKBiLVg/F6PqhOCBMOTwY3u5i0UnlfK7uFzDhjNHq2rAcrpGvzSVb
wLpMm0pbn+8XYaGFvvi6kEGnzNRUzGh2eMD/zfaq3pkpirKyUOOWo5MtIGlQezna
EvLFq+bONIwq/pCOIDh51cfScVP6OJdAwcYSOwtZzrU+8Gshu4oIMdQFva44lcT2
csmPpuwxlF18ujmHwkEhJ1JIShzAOP/VPCvA8gGhZJX4Lv6x7/hbRgYfYDJLDqZc
UWaBBmv24qBWUekXZD5aykgqVAsClMiz+mXXVSRubaXtr5GUwPtyhYpoFy0qQDam
cU5ZHFeOEHNQmXaYNB5cWT07SXP/r4UJty2N0qv2CuJ5DwdKXwWbUcA97f8XEDDc
IksjRInPhsmE1SrQNIZ9jOMvWCs76F0dMIatE3NFq7m2t9eqpPwd7nnPbOjKojxS
lxBAIlZMAXpOfmrBlF6bngaN+eh2J/IFb2+HH9IWEn4rnhWTAe0P4mk79SmTq8r+
kZW4P/nDG0HJPDriqHBXqLIVP5sw97DWeCjtfXTisbJn7S3iDpJl0BLclPTKR+El
O/i0YZWBo8woRDZb/RSV61778SDkp60uuhj3NIEaeQvyPyUYr9wv8DZLw4zFS7IJ
34hHfhh7d4u+kj51pbWOKLRawbPW2QRsUif+CQI7gf4KorpDWweGxyTDKi5Puw7D
kQ3oMypQYP106nIkIiCXWYvS72WfxuKfv90m0KVv5cMUaZh2Nqkn6nvN4gaLgO7d
mVoebn+24Xg+7yCQqD4a0A==
`protect END_PROTECTED
