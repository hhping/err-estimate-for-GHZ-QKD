`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7VVj32UV0GjyVNDCva8c2q8r0grDeIi2Z0+M86n4urLiXNCu6727xmVmisF2kMxg
0x/9dGQolw/JzGe0Lso20Jhe2OwCrzraQR0i1Fq7GJJBp9UsO1iS4L8o0iESDT7Q
Ur/5oJQaZScxCjWroEYtq6ZukKBHAqn+AUwsIc/3YrPBzY4yjowM3v/K7N8Fgrub
d5jPil6lT7CdWV/j1IBhSZV6HNcVkHGr68LDFoABrggiuPlYMpgBYA34MN+eEklf
g7MazDjRslfJAI0h8BiRmJuLgsGgaT8indzYX/JLCdsAae2SXL9vxexyeA1cybg0
9bIzhmuCK25bflUsR7cRsq23ZBvJFRSShY/5GgPHUDkO2Kf4jJIe4oRmLTYNEbrv
oVcPTCtQmFEqnmH+gpyC/A639F2+ueDZnLZjnG6bvO3TDJRUYBeKqjn4VQseT+4e
KKjx/vD42B+k8X5hVc8H6SCcwc2+5B4JfLNI5tudQT5FTwp8Cok1X3q2YaBwYpxB
31A1nvoXFSNPPAiqnxbv4mM7ntmTHCvj48wM1Yblnf7D6lAaUYP9Vv1V6cRSrXhl
rrWSW5bP7eXum4kvfLR5F9E1+8XrlMrJnqS8ESUrwNXx+gLuVdpzAPIfoRU9G3pi
G0OzmC4cC3qHIXmZ/uX/xWiyfq9pOb6ZvdtiXuFDaf2ls0Q88N6NWqNmNxf+rj+g
X3/XT3IJCCtttcBVYgdhFTWeBzqBeJ9/EwnfEPf0xrRtbdtIhZ/1qUq6xC82rAYa
gdrL+rXyb9p2Df9Lu7bVYydummIhV8+DScJ332Ien/OB7IA7YaEuLKBvHEHd+G5N
cv1VbkUlE6J1SqPFMMmfwJeViW7wZwvB2iRCxMIwVFTNQ1+Gw0ERChFZ7atpXmd7
QEiYV9SacpIE+Qg2xOLdCxRUoNqBHhWRgd74CLpu3TCivtWXBvLlulEwtCCpWNLE
0ReY/ibgjauxTpOjn4VOWXUeC2++eE4A/51CkzuKr/d06SaOzsS/UIMqqfimW/2r
/JBKawuQm3hqrg79tsT4Fa/2PctptYDYJYYLOuHqWEY4yqu3Xwtn3+nRpCRzjDCC
B/cjFUCMmrJbrM4QMtmkfod9r8463TgUcrziDKpvzi088JyQ85+vZcpIOp4WV1AO
WJSGwc0Ja6npZtjGy0sPNKTphm24fG/yD++A9vSGgT1VmaEYh92iySWn3m67IVXE
Q3Kcb6BcIA+6zaKnKxLBa9nGj7TaGt/JPDH73vQVYUYXt0c5BcSrrn4WygzzHCja
Jg17rlUmmpXXA17DGEcZwLY+aitF4rqhH14fzWG/QQzV1I3OK7hK/VOpaA63M2c4
7ww+Ba46UIpwcgIXgAwdRC0NNQvHfW29iO2on+zUyPfHbllCyrEzCnPbwWcJzHN/
VV7oS0OVgB2POrIg0FVEYyZ3RAKZhprbonjYf5z0cnP6WEvBIlgVXj6z5FdzckqX
F4tfFTINw2Zga8kQxf+xqrBS+JZMDzuDYjYd2/kJCmlxWBFBEYgx6B+UzXxwgW7s
bZX23LMwjz1+M8EvZ8W9T1iyWAvTMesdClyPEJBB1y6N5S/2luJigxTw1ejD0x2H
WPUNP5XTQjTLJWkWZTUERArXZxQR/WXKLL+h2HUQGzsf4A2X2p1/5VzQeQKAoIts
V5pazNNEPDrjlxRoS44+uzuUMg9Bx3fwrqVIFDeyPfMECGn3+pDjVK6rpyB8DvO/
IwVMAQcveZW0W6qm0Mi8TAM0o8+NP2j8XXMbxsh2sA2EZxNSBRcSEptnK5xixsnh
mNv9ZBRyjSaQuL5Ket3LfvO5XBQPD0E02a9fWKNzXRxFFOwQ4Fld1a5w28ATbPvG
K9h2VypRu71ltxh5Zy75BUMhVVwi71JU2tsMByG5KpmnUv0hTwqyA/yJXffepbhI
p7iGvnLj9sZpY7ZsNGZ9qN1JYHCdCGXHN8dDkG2b4PNCafjfseGAPrql4Xl2oaW/
U++RRw/miResRGexi1CvK60osDdYDNHTaF8hPWA0/wxJzunceVaBzv90KMZO9X9N
RH3gsNxpKPDXtuhlovFdLKBXeh8hZ8UrrxHxAxCssF2eWdtkDeY7NYTncq0j1ItE
9w+PWPvoMpfav2e+b6C4q0zlEWBSWM8Tywoodc0kn5tVD6tPKMFizCl9ZsUBZoD0
dNr8bySd7jNmFzKTINTKKHldEMmTusAhpMg8zdmoTHzM5aQUH9YZ7Y18JHVwrwnF
/tgtXnIR4YEWQ+Cf8AAM4D1GmP38AqGyfzwqGErfEp9Iyf+0l1rq6rqpl6mc9cEu
+GqmVxJEU7W7NmOJUG6d+VRIExSUR9kWnt0RbHBKDHaQLr918cZ3Tm6ApN//L6yN
xMIurhMQ3bq4+YUbBbT6FsYmPNos44LDhI7FzdTuM+iFVhekgQasihdMnqlHlRN9
YxBAGO/KNcNdW8QZKbCh/BDBnS7KIiXguQ2MCIHP523K97xzk9ZeitVhrVeOYCz+
NvLxgiIiE2m0yo7GDUzegUZ7QLzzQJOp2RFwfOgs2GvVDT2ko1ppYrZNxzsh/Cvx
u5ZAseyhHczlSlzVAWhA9iQ8qBrc+/tMLIK6yrMDjmgtgarkr96xxkVqbtqWSUrq
CRz+hiNgVOoWsZFWrYH/KT0pRTynikqZeRm3QDX8oItMJadQcf1l+YhvbVc+Uznv
VlTShM0RopY32/VdF1Kp6UtSwFPc26W7q47Z6zWtAPfQmu2pKnJ6J/tGUg5YWrJ+
9deAdesleiyZktk/s17qb3HOpc6TRf9RfEXdMVEqZV56TSMMSlYL7gub/Q/tPij4
BjIhIccLQxofl+51M7M9xyrMSymurIrfmpI5IPshioW65WIwaVm+STAECQCd1L+9
rmcwQ937XWglrXknVNbHounBYl0/JwlcNCFOEKLvtsofE9UmWkGO8RVWyG4L5WHQ
uFXWckKtDrEZa2pbPjthhniqx6pPG4Oj7k7Kl7/wHlwvUk2DhPHy0tIIra3jqxG5
5ZQJXaEUWHjyIluJODOQAHlqZ11Fee+ygsL2kjcILjvUSAmjSqmbxYwbYCIyk/aC
hjJODYvHFGTvg72F1Eq1Xjv91zMD87aB2bCNZQaf7kxbVKt2lzEXC3Q9mYXY8vm4
mOPltjK83awV1KgwmqqMGj9uaqs/PuM8h1r+aHjgvVvOYz6fFyAQvRgIEp9BxBUv
PdAZ3gKfiUP3VVZEHzrZCZ+8t4/qdx1XC/lBBSJBGZtfYzSFX8nwar/lZcMsi1ll
qFpNzVrBuYLXy9oCMCcJEyEygN6Gn5EuYrjyWyF3y8nvfm5Wl+CnmX4q4zYLnFrP
6OnRz871LK7xYC48WlYLm5Dfw9FTczpHflob6KA9ifI4XxJCp99S6CkHorGITl8G
`protect END_PROTECTED
