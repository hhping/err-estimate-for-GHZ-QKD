`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJfkbNj5jD+yveqtX76Gh/uC5M5FYHgBT8JMgheOnu2SnhXRSIfhDr6yp2VQNtsg
R1263+0pS6r2l2X9ATx87fsegKEKwirAz+bMj3u8vEeXUFMt86Jd2xiLze6IqrRR
BMpJKpVNtZM/kVBi9kJ2ACZ/LN8wKOtP2MFTpUgmyHi+Bq67fapGhN0DT7zZNLDa
CYIhNurUrERPyqoXv6LzDBIDuInmML3XnpOpR4yX9HSpRtR7RiVnkbNSod7YZHsv
rK8Mya6QBx3jMwxAXEwxCW2HRqXHkpROmizyt8XC9WUwmrUJezY5ejohBfViDc4/
HRL0i+QU0xPz8Ewc3qBlsqFZT+HY+PRqzrJsm9WmrmhUZTM7mdcmuQrzUkBO+dvA
yZVeup8ptUaVHPTs/9ThNAT0vHoK2ragvvwp57/I9naXO7FYR8rTV4D3PT+v8AtU
KZu+4E2DZMK1cr9+Vyxo7Ml+5lzo0XE6RYPi90zalJzTZKX9FaPuj2k3SXhuu2qz
`protect END_PROTECTED
