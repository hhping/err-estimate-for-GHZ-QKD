`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
okVVzSKHjmWsD4FvOrflt2HDZFViEmIjF+2mLMP7q0XKY3nyTqJhkY14Ss0YCVur
IH1bhVLy/oW2LTRxm9vvCsqWmQwn0CeK2/x1MMSOzk7vi1zGI3p6ONXRO00481hz
ZScXAGzRsi4ZjGuipoKeayePF15j6Vj8hOm1zaHUpPQFOdFZY7m6quoTDDFT28Yc
XOi8O0Tv67XThCWegdNZcKlEiGgUmhzjYoQ/xFyuByV96yAEbdkIYQU6QfuD1L1Y
P8LODUzPi/2ZlPjiJSYXqOYfCO4uIMuugYMyCk+pAjXR9QP5abo3vQe01i2qJ++J
g/vt47dLV9Ifz7vQd2rsmwtx0K/TYx/1jvdlzhiGhRRDZfHjBb8aCZ576a0+GdrG
TdTHqzJRhaK/ZAEHXRhK5XUIJufgdUxySficLdc+hxoKBO/fSBozM1vOrUdg83F+
lpj8EXAGiw2t5FA2dZhW+cwGbAl/93nJeqg+Q5Fh+CIx7SfbDPYQVExn3f85ucMq
R/KblN36bDPTs3ObwRdDqACTf2VszsM33wHAizkclwOci9Qiidvc7waDTsFKNhoQ
liqT726vKK3ASmbBs9mhVg==
`protect END_PROTECTED
