`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sd8toIdwq5FIWQ0IuTAHD43XRNvyErIFodV39DtakYG17RLxK1lzCcJkKyRBaFn
Y0QmPR4etl/KqoqCGZ6Sjlt17zgshJjYSRUJ1RyRM0f4HgwW+b0CybRe42xm8V7H
nyXLGj5VOpKLutTt3bF+O258ZEtTcIGE00yp2nCGKfjK5VoRXnp4vgR/ZwvroYCA
/fhrbxGuB3VSY45OCChAkQ8vrDAV8NfF54h3hsW/o93DWTLYv6mqIjFGZTzCFVyD
rbXaQuYl2/+SAnuAtKci6abzmAHzN0cOf7qNYFzxHZ/rSvsyp8rOz5Tp7bBjqQ2a
f+hP7/muOZNGAf9pQSd3SCjTYhCPrsbIKTfEq13//IXbnWT5iOzj4WYM23FT1Wkw
y+kgbrmpl/VMxm06AVyPAfnjU9wjRNeiShrD2nyWJ+2nNH7gX7kothPuFwyiOtK5
L3dFYQaGU+6r5QqX6+QFhkBQxuZ2QC3g5DG93IwYTix8cxNCIZzvSL9mPSNxsR5T
Z2ebfMy7Q3BZdsYMUM/6VPisIbb9btNcMIa16j9Aq7P9VqqPXEsiVynE1nZN4i+f
JyDQw3m3lUrJa6wTwqN+fWEK8J3SqvR2h7tVfXc/PCOIsO/lAzA8GVwL9Utcu2jF
ESnvO1vFaxPv5sBK9Y6C35yiSSHp2Zx/4CaokBNKP002tGyAnpfjzJ46719hb3rh
ca4rsx54F1n7EwJRugUtJsoXIWmrp8TIlEx3wFToVBoYbrikL7bCepYRUSkXfmMJ
r/aLptYiq3nJvJRKPrJQnkzh9UPuFIdVaw3CsUqsp0gaLjvbdeMOw+lr7HrNB55q
zrMgzsBdoLZwfP0fNOusrw3UqVF359cqZLk3fAcrgarAnkn0yhE1quqrfRIQTOMD
hbDZuW1h3LAV8kV/Dkug1J1FnXRLoyFUgjA4pWE1l4VXT0LHED1BaeVGtrSsciTP
dGFgm00vHnOBw4lu6Ej2giUOOErpjsUhMLjnTvj90E5uKCHcLkMh+MYUEe0fQYQl
/p6LRqI2q26mbs4s+sLRUu0b2/1aWq5LOp4HCvo0oRiZxI8KQEOiU5EpQ2aHJOKG
o4aQjXr22cjUpqf5cMyJA5z0+zLcXgn5E/c06wI0StOqzBMppH3zvIH+GTTUtfVp
lGznHiLDEQO4ngSFvET1bwhgw/YHOk8pY0Gi14SyfiyYZ06DJyuPq01xkCCMUGDS
i3YI5o4qOtdZ8X8genNYU4YZfvcph57nDjwa9sPGEEeArnKIRZ3e3iY7eRDZkUZL
iPyzUl7cRbJTFoeWOdYU56yYe6UJF9UFMnL6v8046GoRPuYev/WQD9mrhMwfECXL
z/JgiNf6NjxrxXdIic9L2zyIuyTtTJkCqEOLe1nF4cWqAZ5WvuhZMk7ghu36eWPU
kFqi0Mxgvk8cc7/Si8DEG4nDfHWTtLRdYiNs6dqSjBTpwLIjCv81zn0I7Dl4Js8q
gEdAf/MuCpi8VD7TlBNsiyrSHAWmq0bCpempBVVh76x2vQsM4ybYB4jmqOnMpHbJ
4rGaI/fR9qeUbZho80ywXkQ9txPAHIMV2nnU1UCNeH8GWyzLLBE4Be0ZIE9FTooJ
q843YB7Yn1+SiAP/UfuEReXYJjr/xgcZLFAK9MYnXUyWfwvDOLRlWpRY1EaGo/k8
Rkt9fWKjKz8BuT7uyVbtfwN5bjikVX0Dif3XzxemCKqtC0E39jmdSnUrl461C5RD
tzFH2e+lFE4Su42RVKrxPxfx6681noMWjlKHtcTxchaojCK7P6+3t0Uiwdi8Rqyp
tiJjY5iS876qgL6GqfLlUu2IzoIizQuehkvJrVERV+ogTWlVvCaxJGuWXD0aJga+
iWbczFpJCppi5wG4cQxMMAajHDQVUDZiJY5JR4Fp6nUWCavBF49fWXFP2Xlz/ZOa
1Hda9wivdRLXxlHflcW3tY+BDdI3T/Tl4p0IqbICdD9QhEQBjD3KYyx8y3QWS50q
P00d27Ig/dDnmpUFJh06ud5dssJASJdKCtt+tv+GxFK+bFKqjWLs7RbuxXcZltR8
DjWzA4IfWKdrJAVz4HV/9+/YNeGMCEE+9ch44OivxuuOzcZ3VDIErQLsdATiNcJD
5/oYUi3uCkWP+KMlpn++FexHj3qmDhGVBkgQBVizls7W9FrO0N3t2i1jnzzbg11q
T2Mv4zxX1sRLnzIOzGA9aVFK7CewOTGmmprBrjTWX9dT/DUtm5xrl7Z1KSsagtaE
kLQj5ag48qnHqarWJqev008Xh0Rg++NA5oijIZAxhnNcC+3O0SHqVSx7Y/txBEdP
szginwF9fC8+gs3s6eI+Kek3gR1FvOxh3ENbgTlEhIM=
`protect END_PROTECTED
