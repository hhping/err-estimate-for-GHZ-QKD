`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjM96a5/OARCJa5Gr2e1Y8IOIFOHGAuXg6HmTPWXw8rmLBbLo9gx52OKCQsen9uG
eAURNhcohUhf1oUS2eNFUxvPSvmIoizek62JSPWupv0zozpsbJJUw7zLaDCIkj34
TzQEV84Q0HHf9Hyf+MpdwAjZifbffo3zE8IeVHPr0JbSLiQftwHb3KH73exPeg0Z
BjzPGho54rlagpk8duwnPWeb0BYsiAGY1eu7Ae1WCM+JAk71zCdbbKuoVgdvwd+t
1TGODMab2NSJb4TdwPPnoWLsUoiynjKV3Er12Pxe48Ja8MdyNYX05pTKyUkp9pTc
hbk6ooBACJWFc2OJqKrKVW6n0EwcH8G6RszU8mWYsFdkXubjrg6h1s8OyIBtSguO
b9QlyETi/wePiTSyor39S/VpMHbRgNbzc33ojfDjlUDM9G5wooNUQ7W49hKvobmC
n9dtp0wSdYOcptGo9Ql0RRAfDcNaADCu3mDTr42mhzRD1vfde+PywGWIigyClRC3
2Ky4720F/uz72LPRvf0sfkUJXaikwFRB/2B4a2rFKTKIRLAgWkQ5gAl2W5jBtbTg
TCcRuNs8zGzNF5lNxR44qtDIwvuMs+MjJwSsyXrE78tbgU73fSWL0brz0azFJv70
hQ+JF1GQO+U3jWcicbdqvU5g+0KDsTSYJ+4iFDPol+DeZloWrH9Q1oRpkqH0fktu
JAllrF5eYyjadkgGNID3TL1bn97DN1LeAEdAhfpl8qwU1Dl2JeL8AzwV1ImTKFHt
xIPVVb/qF0/JlaHsJigLXJqg3m3sQ88snwbaekYinf38zkQGL5YTOpxqkVPbMNPH
yW9lwg/6BerULjclexkMc4b74ZK3PLuPqQwhp3DiLzfruYIbRRkJYZY3eajojLyJ
1I++074yjsIclpb6hD/qVsZoqHMYYZK5n7qEsUERkLZdQySUC2HQ2wY3wLqPauk5
aZOhSD8x3CcrnP9LMBg5K0qDKA4C4Eh97OqhW12r77pRRW1fbgY5/Td+wMLxmLT3
9orYpOET05qRZRqmdZmwYK0YU1xmOTWaiKDpcicgQo4O7rHs/hYVreHt4vKK1bSJ
e/hi38OA0innhK9aBiycRTxMRMxceAsQcmqr/UaCkC68Sn3yjYnJBA7ghUfGdqbX
o3NWG9XdnLbVMaW2X2f1R1+DTCPU9Qd1fmutcylyTdWGbH/kQmxIUVMueI6FcZnJ
WXcKYx4t81syZewZEiGw7tJinS0Etj0tqYaSvWKPo8VvhAybrMCf+70T4KIzNppm
MASBbg3Wd49wTU2cJeUhboo9BcpFkQxMTcYCQNap6qTSx9RlTM5q4OuejQ8qha2k
r/NhhFWj1MnlJMmT2jeiLGrGcKYHduq2sWSLZ+NAFvrI9CSD7CRFVD1/B4bWmY6J
Ydb83NIp40lKoFg4+k24X8N1eAmLbXT0FoGS+k1pBjEIXotsdYZ8IZLMvIVOxspn
3CQF0f5gd4rmP4aSBVyQjQ==
`protect END_PROTECTED
