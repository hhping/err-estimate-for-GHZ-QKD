`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9YmcaHyw++I/FAQLpRxzhFhh5s5gk8+DlUUjUmEXcYKCsWrKbn1Nizp+8XKkwXw
rnEIpHh2tcuoS9eMXcabYvkFdm10fZil0tvQ1Gp0djK3cmqKvCWIGPVaf1PRhRaw
Irc5cOcYJ/1JzPRZYAYolbUBsZY5/Mer+23ew+vwW6ZAHGM3M2MpIq0KAO3RFzTf
oyvRWRAGkGdeQSligWt1JmYeIuMocItT2NcBfUwai3E58uHfLJZna6O53L/GemHx
0j2VOpqbhsrBVKVuNrmqhtYD+BayYGBFCjSZ0UUuK56YkAAL5lNuWn+el4r0cti8
UPVFzrJ5wPHAvvD0rZXxdM6sv6ooBu8ShW3eWl9DzsqQSCMoiKcNtQk3H7kE/dmx
JUwUVnYgq8zqDnWfv3NX/r3vJuagZsS6Z9yCtmyrtAoQOt3Zk7oB7j2/MbKj2a2+
LPgm7itAz7UY6ds1giEOjRMNyoExgNvC75l+jNVF+2Q67kEucu8gEUwyN0NypJyL
XuvEH2UbbF2JQ8M1nDglYI3nBkSq5rD3H+LncpLg5h1yf+xmMy5MOXz8AZH5w8vA
grOV5v7rhnhvFzJ04hlRYD9C58Xm9aVBPHV8HAKqymHJiv9gxBYOFIzR/fpq0rxI
`protect END_PROTECTED
