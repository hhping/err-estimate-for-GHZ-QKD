`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2HxYPSUOCAXwG/CC2UxsWDFYNesN+lT2IpvnUhyRep98TXNv1S/O4/z750LD3nX3
mSIs/z84rjVaPdVuv+nFF4lrxg9PbXn90f54NlUVw8pGA5naudoTLPA9nYu4Se2C
bv3rRgZuGxdJ2gMJVhJHJzFUZwpvYklsa1vIPcF0KkuZBfZuBgqDk+8F4CGa5PHT
WqTNpYjwZ7+b9k5DVmHjumAX5AJa77oA+1O6ILbOoq/N+L3ZGa5XOHhEYZOgEwRf
1dNxXcCjxwNifDJ3lrFYzpE/fPqRF4fNhZ4v2cApb05R7R6+v1B5u+kBObHWkeM+
VOnnslRZQ9AX07VMjrL/df3AzdpekkDs39eaDH0tbz9Y201Xg1Dl+SX28OC3uEIY
+34js+Lhj5r9053KBypiEtWPLHUM4SnGlDsUJjJiSuMda2s038w3TXxACht6O3NX
t0XWO87ZsHSwH16tYH0eBheuSfxzChCQCFy1NaT0bdgAG5LsFfZETvfeAd/aYxEB
Y7NS1w4umnFhm85hvSmfsM502Xj4TEU8ureIquXlu1ouF5WkSqV2/2ImlDjSTUY/
fdP8AaEnPBuihDHTZ2lXlAZL2TqZ/Ld4TNrJIVmcQLYlDEgnJjduAd+OLlgXTL9h
BHB9Prs49td6qTd9PVY39F28PgZcLdGrut8Kh4H9sko58oXjccLdmFpaBD7MTvhf
GsTrvJtLuFXBiD7W4TEMxu1fSaUr7WSLPMNJN4LVyjaRvXXJ1wud0Gw9B9Iqlmu5
FlLujLzfMjb/3AERpRybFsrX56JA7iROjFC2mWL8UEOpS7Ez2317ZBCf/sFIg1ML
KFcs4RAnaOhJs1z6DBq2dyHvSGXihSY+dZM9fzcXOzZ0AVI2/UyhZcqtCwgrBuTx
GXUVlyNrkp2foNVGK10JWmjEtY40gmDdimnU29zlI8fawaowhNf25pMTtgIG5k1p
hFK0prmZrcOJaxzEIAqnJA==
`protect END_PROTECTED
