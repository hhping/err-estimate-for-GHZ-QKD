`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0nZvVcEV4wo+tvWu2y0A7iiLcQK99PPtPXme22fp+gRJHO1pFmQLO4H5qrIsmfWH
qT4MBAL20KgakPT2SAnrNLH+Kv6OY6ggETe8PFzA+VjO3oxAQcTU9OAyke1RiRuz
LR8G8OmBqFASeszHZ3P1a3mqVrurAmdt9UeO/s+cFFkneaWC1mzeRBw3s1SjMv3Y
LT+UV+5YohIsx8BQRu6jesdkqnXYKoF7e4EMrW2s6RtKZUXLBnRM80svW9yqKT6k
VIWdwG8vF7q3uVDEOjdy1ArOLEJBOWIjMeiuIj82KndGl3L006zedyWhJAOpXjxr
SprZTQZSAXhnpklu4d/wM9ZwH4Tu7oZehYBa7j2gOcTKMHaSxj374CPL4q9w6HMd
9jK7R4vnsaiXF3XQ1okDS7Mza4WvZWnJEZas0ZSh8FTY+kZV4i14UJc+M+HMCJbg
QQriSaX7Fq5NM8h6MJA9e+1hwNI3AfBwT7Wmbb+YvVA+VJSWZNJ6CFX2y1CGIGiG
JTDIVKkiSRHMJtFntjZr/qca7gfG87/+iIdkmJKoyrP+zJXX8N7iTQD5PUVYy7Qe
ey4N4IGTAYf5vhHVs0FSblxeXvFHV0pShKltR0TqKNqCKngWbsKZps3/UwDaWD9K
WY+scGoCm+1aI4tFkWvoQNNnRuStL8rKPreTmwu/lCtSYcR1bkeBW/cVhmwO/m7v
G+BsM7TxD+RFaYaEjXTvQ3lmjFjwTm437zc3uV4cbSNqZCttNo4UiZXnStuelRAD
AvlTmIq2p8XZ7h+NDLIJuWRHgBlMoR6n/U2lXTghGI8l6ZqYDLreZ/uoZOT6sF4s
klNTRWUAq+7Z55hyOwl0HIlYC1IDXNpMU/2NJO6eivhydM5FvTx4dHfA1MIQlGz1
Hc6gjt+4+xUQowuRYf3B7dJIqlIJ9FDwnDmy8pzOssDxkdLl9ZwrG8jJnlv2VdzK
13rBdLWgE6TM3ZrOIKaQjhvclsldj6lv+wY1BxF6BzUV9uXbwzLoE6eCv8l45tNW
yuhBb1fFCU6err+W7wG1UtBi8fldRa/jOFZeY3BGjM6NhYKnOMlBUFjTTnYT19Vy
Cx6wht3LTLmnUKVXdVrcOSm57ZWeyOJkpeg7jkweJkgyK7VsRR4sIY++ZH+iES9j
`protect END_PROTECTED
