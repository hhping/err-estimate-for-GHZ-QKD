`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jl+hrVODzv2S3aRoxjjleaWn/9n45Szu2lI+mTWEyZwlpywGCPXdd/hwow++vzlH
kShMTfvkwy4B8KGa+L/PdP4s/zl4MARu3ObrtP0NTS+IgZK7ga2ay4mdFPB/FbCh
09mTeYv9bMS4r3mgRcYT/TYwoC1W9lCIbb6jVcplj0hjs5P96L83aR0dnb9kM4bK
mAwLpJA8I7GpJ5CfCvvGZ/Q9flvasq9DwiImIeJOuvXX0/gE0DJG1ZUJ6H4xrkn5
XHflABO+2/dzRveWV3k8fPDWp1IhmCxlNSWMx63m2d9gBzrLAOh7+S5YkAD7CixV
5iACPx0QPdI+oAXknjhwb6fwBX1Oe8sbQ2Wc8R6ehYSzKa6tZ3xuVm8nimRKoLcj
j9fNqxrjjISGHAkDawcb1GakMfzI29lh41w3mdvwfioYMuCTvdQIn4o+lgwfZV2B
nc2u/T9lrRtKM8ALgE0UaUtnK9xn/HhGyYRyucW969w7oT2ml/twToyiJCozf0KJ
bpmqv2AIeGxBikE1H0EDKQxnr6yOhfW8nkV4Mg9VdoCBquoPVWEwrUyOPm3Agca9
yVJSVqa/2s6zUJAxlZGg8V/oL1a18zflD/9wUYKV4AQFf+s0R2JfO5FQlc5qPoCb
xJt2uw5qmweLZUHnf4+Pm7VzF7IeZ/rrOMpmbJKKVUYdyBI6gi7W/AtZL2y2YvZn
eULFO6UekuuEQd01yR4J4s6DNptHfq48drh89nCrKWBjuhHvR5X47lyVRttIL9IG
lqRivo8VGUiWCbrpAota5LRq0kbwwNhv+cR/i853BvCuh2wcFb8dpnUN6pNhAgAD
QFj/66It9V4JwvNZ0P4vZuub7OoXWiIsHxhf2RO6oG+7oy0XkGkuDZMVnJhkNfPd
cHfdUtL5pyVtMqC7RFIt9zJ8lRybF7LNC7W/3V9lQtxngZTLgQ3O9xniCRmuYQ+3
lGqfQ+tUX+24iDD4m4MlIkGffljfKVKu4jR1s1npVWmxz4YLxtFyo9nsSKja4NRO
57YbMRHO2PopWXUK4SxBHV/+D4Ifl5ZFVKkjfp+h5+zklfposCDU7BR1i2Fb/Pu1
uZXcjlaXo2OBc/3a2n9jZvMkHyPtTPAmhjzV6/EK/kPk+GCwCG9KZvhcGmXEeTLm
0KbW5afUp1lgOtN7sTbrsLFuRvCPYmMjZIgAzmN0y+wo6aOpPqlWd1doYelgegtx
aBn+QJWRvO9aVBS6jNXbQVElZEZp3DSUTFTXP/+sIFE3aS5MqOPuWZGI9gG/R9Ii
Vxvej7WjPuE1spzqseDxIA+o7hgRcimmKJFXZznrzWOMYJ/Gii6jB1bHG3lZcSs6
ggp4zqTj0XWOcnOytnfJWWb15FUU8RxXZ7ErJCUuo8hB9Icjn+4QToirOMjPRGVx
i5a7ePhr5ChYr9nx4Exqzo1EgG1++fKLtpcsjLHRowwqLvsetRXV/Swp9HCe3QeU
emmbznG1dK7PcA5ICLloQpNdG5SqIk73J6cmdwXYTg0Gw+BRo4jrssstqKr7isXO
Wpbxrz2/8FwHk84KeC0MboM56HoSVs6TWOpf3h0p+R5PDelQu6WAFhWY0lNZY/HK
gkztEN8snznj7fW61JPeihvKqXgdQgdNAbl7xAyul1zzqK47MlMP4QaFIT/om3OH
93QWJ33qL6e4iHO3yzrjwuUlONU8db73qOwHYblzIBRnpYRQFvwODPCh9ukcGjyV
Ha6bx9pPG/tcLQ5MMF6klw/6phvm65grWLbCULoRteF1CLARu3yHkxs5/NjzAAao
pbF3MybOTOm/Hl9li5ZOiQ9em9ffVs/qGDoWDgSjBDv1B6lDZG4gM5HPeHzjZK8Q
2rHRpVAF4JeYiG+D/kXQ1WKcmEQjthUeKabn7dBG1g0UR5eotk6msKU7FS01qWJq
5z2kWh+xtOlTcnNiabvNhK4UIjx2bqhG6Ayg/OTuwf37v4iACE+EoYctuPMV5ihk
NfHUPTGSP2/jVDU+/63tV0pEz4O7J4qP9I81VqqSE4Ia6GA/Ts2FEYBHvFKe1t91
Kt66AGktztw4Z85LR3cwodDO/Vz37TCPH1cUou1NTdMZthm61b7+tgLJr/f9YP4m
pLzyHB5xVs65RvfsRLVh+8xdKhYEIN/Nb+7cGHyMZYa+Z3iHPihV9bbGx7PUrGy1
UZZb2Xa24XKZkQgmBYUz2MheRmYy8Wby3M1oj/qQKKN6Yt93khQePJQ+f7hLBME4
UkRvMkgZPb9PSB3bx+yvg2Launxp5gNZB9s0Wp2T2YYKn6YbL4lMjo7urPujR8Ms
UgA5wL44m4kZd0p+K4m49WLJQdBk8SaI08f+Mw4mTFf6naC/DJNA0J04DmJvcpe1
DvYuwycSo2wKgsplmiRbFKT1uFY/c6ayLn9Rek7oYcbrddzqXqcUnTmI5zvmDToc
3udogiSv+XhPgmMdvV3Yl8zZfIIXSHvmJvIfDMviXPb4O0PogTZhSvcuqCRVKazp
Qmms1ldqSEhsM3tYz24NiYiqWW0lOkzfQdDhx5A3T3bgPHDX+gYILjsBlgUJGH3N
vw+gmGUNnHAtLMFrmtmy88mhTu+GrwVR9XOQnCE67ZlX37kdcD0mU5+rBXWfSydZ
G1h3BlORHQU+pWKwf+D7N/t/18lgm+a4Rz+2jK01TPf4iKzrexCIi6MKphVWG3BC
GOJRO5+tqJWdSU13lGMSFQ3KEVa/k0RPwszXsOQHXrLm4EbAIgSfpa3IJYe4Fw6G
Wenc3tljiOW8++sGEwBkY59xwP+oNhsqfJYOg6e0nTdV7IhuxmoyIUSOxsoe52B+
9SwZheU7B1EwLpQi+E5VsOztdsSdRAHD14+GJHnJ7ymMyEDB9SOxvjEWkWLM0p1m
SjqcEDKoMw/Kui5L7CZzctUlbTK61/KOJkx+cDGSy3/fs9jl8RjSIOYRg/oi2bwQ
bdljiebYOZg1Hi/zgc2pquY6aguZMghZo81YufEqPH2mVIwuM9oaHh2g2pVKeEMO
WlmBDG0bohhOrnXZuUKo3oChwS5Jquskd+nW7ufY38KHtQKnsrhgf4pI7qWzgoZo
ov5iYqN++GODBdgGwnxpthLpt9HIuAaDJbeSL2TwfMPuupX6RcAyTwxlg9nmNfo3
Ff9QzgJUZL6Q7i47iPZIgous286XKWOidH/Camca0io+2sYY8bkVouW7sJcJ3c5F
H9gOvTdnO9DtlmIqCgoz7+ru+XPEt24/moC8ZRF2/xEVUiw5OMeu3WjlqLYfcvLl
b6x4JEmdi71kBcaVoP/OIm2F5+IIHFcFEgTk2pkukAa8EOPC6qIc4JHrdhUaCIJn
PDIBzrpCkGvloZb7ZV7tGSVOELoJ8JzCeN+TzhSrWOujxnbK/TNQi5YKjY0fXIA0
R4JR0Dszocgc2Is/oYiiXyNkHTPtGC4Yw6JzBIxQ+HHaBtwGmkSWtMEDJdSHhmGK
RkD4WSEdliy5ecoXPBDBnbTbn1cyDpfjB4l1lAhJ52lKUzBBO9ZB9BJ6KMk0iYsZ
Roi+I+N+losrP4HrC+OScB+RctI5xssVblww4jkuZywPJ4DySrqByZsKFv2LveyF
pOweOvcGyQJF+2UbC1pWKUHcYMRTqn6GLWQJRCc7TSo2fgpMnwZL3xUVi/zlBqWG
sA3OdTGWW13yU5mutttGm7LU5xGW5INrBUkcazSgjwZ6rK+H/i2In9ZU8DcZpgRM
VMit+9fhjCH9uvmpr01CRbIbek2u8Jiuhcv5NlWT9tbrdhoPxW2FK1udUcl4LI9V
UEh4IaSOuQRF/sxL5db0tbPCI2G4y5DNM1/3QWm8uK1IwCpRCIxVdItaaVo1fEGL
PSHf1c2B/EzADjeWRlNsrT4yt58T8uQq+W8thmHaQirZe1I28hEAuNTSWrQQNbbx
9GxqjAfIGNwaWLmxofMagG1ODv8ozzWa7S9VWGSmmCCVmI/Rg86SX+I2rUqiXC4u
53KpJoHpiPliQ60rv+heEi1ztkFXxrNHKMZjSNmXDe2B3rv6lLfSvskI2aagy840
cGvq9/r6K0z6fM43r6L1i1myPGKylZTNP9EXS3zDuKSvDimTE1gTbSb4ergY5yQF
E2kvQ1YR8Tsa4YevE15HVmUqs3JKQZKANvnfUPSiiDGd8IhbHgxq5whSLpM+fs97
j/NssMNjtV+M8A5c05dB0cpwK/FcUL5nywFKw2r9SyF5NVukGa2NESubkmccXzqa
+4q+eE//gW8uvcS9H8DESknKX0NZTjqyBsDzRmWel4uIlJTbTc0Lb2p7bOR99efk
YKF21cXrelfPD09QpdREWKth3YJLP7o0TDwkMzdlKcl264MzYzb/NuTYd2EITCOL
0ZL0WRWUkGRH/7GjHmt6FIVjg+jE7tnzGk8WSk05BMKzkLxKgvw+XJuWDMG2WDEg
8656oH2EAz8WE9bjHBubZPZLs5DylZKBTr6SzxJXlZq366XZtR4UFL3VV+7jnBws
f9TfuKbuJMsfutmu3vteFkUVCqu46mQxT3Yuwdt97ygFDgSKtOQd2EOLFLPmAyNW
Anav13uq8HaHdbe8CLL1uAmEB9tE9VYnPH0Fg1NWp8euZa08Vv8ZPwY+fVExyYjr
1acc3HkXQpPVw8vNyp2eZ98yKgdqIAa26oYA9BG+fJTE+lHwLGSlamTKJBeSmDSk
wysSvm1HHToAPPrHalGFjHkMDAzyxT8qaJtimXAaGFkDGEI0l1TZSAkKWFAx8/tG
WcBsHHh1fu1M7++MyiuhzLe3C+hG/I4lauYksFouXgdUERrmJolCfkIoE44tfxpG
JuGzS0Jxf/Rbvd5L5DbTandvxkEECrnoZ8yHWDP18V05HJqAqMyJKDwZsmWTVsUf
NtqTWxhMggnQfsd1JoECB03lQZaXQUuTwPwiXYeTSTE96gB96cWce4GhAj4iJLCo
y5LsrSktrv3kocM1os1hkO1jzU7qqtJPxy/gZYedxyOAV6GV4aBlzkaNe0wEsPn/
MzTbrkB7R3dSHZ2EsMKELJWscYZ9hhpCFSDiRXt5Iu9Y7ACl35Pw8oL0zYzC0RA+
z5LL4QpnzGndopCVLlHO+/RdarQpj97wmdSNFvH0PXi7Q2blDKcTMuazcDeqw9bh
aCEGrQUZSok/Y+yzQJsGst4+t1fJqbHVkxRI+zcluz6Ixbepyz/2n6rtKgSFAHHq
NC6oRbikTSpTENwmhD8mbygfWgzRqCT51UdmEGop1nAyneyTLsWkllBJDZ/rV/Ix
zlO7EEmoYR05V2ewvsej8O2AAkni8lbL4gUAb/Xbq615rck0jp60mDc7vs2o4Sgx
YX8WtM9sC0IhsjKojh55dSH5cvuvz4a3nqXc0JkfSxVyQG4dZvs4hAmd9FLty6u9
qM+F5z7iTnI0GTo+2ncWOv+FONkQedIkDyw1Wtph51pCw29itxG4VYxcwzUCTZQ7
z/NAixNLVZF58yVgHf2kitR5Ml/o1B/K/M3a1izg2I21o8sjR8pagUvU26a1ko79
Mq0gJ07xXsAGI6MyDIudOdIDjwO12ivAVzTLoU8nhJzHZk+DMF5FgCP0g5Ce2Avs
tUwgu18BVftpj3q3orfygA==
`protect END_PROTECTED
