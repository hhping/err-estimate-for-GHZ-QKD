`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrrkU75qLLo0sl+Iyiabp1GfOGAV5k3ZHpYuvNLJ2HD6NcTBxpTKGV1L5SVJKpXx
FTbowxlw05QCehLKzizl/cvpc18RbtKZ3ECQjrb9fvySsPW56VF/D4m6J0nED2M2
EfgewNmsA03fxydMjN95B6ELL3SCsDMF4p+sMzr4euvfUEKUJgNdDkKAoN7nncAd
HTlf9G1pZXhJl5qNGzM5PDZZJEYpH9Dmj/EhWCKKM+4POL8FKmp/lG+sQtKQhoJP
gPypws/Z7m5ygxh1WRkHMSWj/vxLccJIGINWfa3esCJXzEbyqruIbnrJN6Mhfq9g
V9+cZArBeFkGtpp8MqNmoNMHZdpJsabxryOxg410vXSY2R5K8thVY9+2lrrOL89w
+KjNz19aKNEvM4czfy1Kix4CWz/KOSwDuiccFqNeFSfpd7jDZs456vzdHxEw0QxS
IRMmOoe6aTyMGv+deKvcrzpbuANanFI9RfCrsWAsAfGzHt6iPVIDHWnqQ0HDK0+K
HAru/I3y81YRkWjR3CwSejV3bEYyDE9Sv1kwxj+1gfqQuYBta4Wu0zTzEbJa73qW
M666l8z+cZB/YNjF4vkx8cjo5W95yyPHFhOC+V3TYK/TstYmaivCS6A9Zh9qQ4B8
ShEe00ywHMMDZs8AVI/Pv9amTnNCVSpkuXAfDuvtHX130l8Fkwd78r8qJyMm9ta2
vb7JEZl3Z1Yrr0vU1JyeE43XHgKtqiUIn2zZhkzS9jxU/0HWQSqdjMbME8EAvcUm
ohXQj/R8VnTnaP7hofHwXV1nh+tc/O81pkkLBDftAqNdwfP2TEzOCHy6I75sOhzw
reWE7MztBCOfShlRhC2dACtpoAG6xEfLKTjzm3tIyy4DYiGv5FxqWcyG05eqSmNv
akWJ3C7ztQNaJKXCfvGasrMZf3IDKjhXso/MF6fG6uzPZ9QutUbd5NyG/SlkRejm
+vI7m5y1NXs+dLqZDczNWddWD928Gpb1aTyGreLHdf/2QXkRFtzJOqxp2rrI0Qza
GbVAx/SzOncFnAA/arFzSIuvyIc3rAJFUZ5w1AQascJntex5f9CXh9iju9QR7KuG
FJT6xcmQ6O0xuW756MT1nPdE+k7xKMEZZeb2VYCogOKcwrCTM8FnhFj56GvidSEs
dNNYAIL1Kb6/t0J6uhNlHJjp/yS9QdBgHjWyxbe9mH/gJkdnI0IFlnh4ct3yVYGy
tDj/5vm1w90TDGNfmP8jWYdXWU2yB46DAD4/dSTi7U1rzh6grvFc6UChI5KVDDgf
RHAGsde1rleuGgGlyCw68xDcLXINlNIYbkTWscXNwZM1bbB2sXXnUyAYwKxG9Aa/
T3AiUQO8c/y+BikP2BSevhn6605yxSgI3DXi/dy+Sd4xSjbYw15xl8TLszbeCgtj
NGxA8jK8RKjVI8+XpEabrr9UVioQ8X3EdfRlWBwWo+peQ3ySAQoookZqr8ooNo5m
fmQoSbSNJVpXqZBcxwZwrZ2Ybof/s2FDx2J03BYXawi3Rx8QUqiZjhc56PPyS6mZ
cROFiAwhbGp6kU3ox1LJwfkaYkKLlQ/7DTta3Rvz8FMSzROJgnnE5buelHA1vo4D
R/ldIwL4OYdKRcN516dQAY+SlHmN86yoVBhKRC67B0vSSRLXkrqLsm/PQwQJ3yhI
v5KMyA1gbUfDurhYw4N5/5eqfP0GYvTJSuR/FOXZQ8fBDC/jdT3D0px7ZoW3tjgQ
3PoKkB39qKq152kBQkO3o3vg94BwGTLfPNBFNjDCdghC44CXoGBODR15mnumXkqA
QhwWN3NAXbzkBlITKGKTnn+poS3qRfbi5/d1pAcaWvG3nCi2AI/8uoD169wnip69
RO1CrB6Bix6SJM/4J1C90z8xhSQtmnGyOPwhMdweLWOap8BqLdVKC5f6e30O39lp
KxDVCtSauBifbm8zTveMXjIcDs8lMQ4VoAOnD9jL8I8=
`protect END_PROTECTED
