`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFCORx4VXDg6uULJsKCLQkmvtuRbRnwhgyWd22ZZHiLEaAdLyaqEZCSgP5OVDfY0
dXsgsysAIoGLsX0VxuoPn31w2N2IPDcoE6BVmoChvuzr25fV6w0JQEOt9sZmhMVr
Uu3C1YM3x4mGpRgzVW5hngwpWnQ3xupuoFJi5hH7DtBjtNsQrtzs7Yav9PaAgx5W
e7oc3jHjCkJx4XRb4gMsqlpRCAYD9s3Df6cy7AB5kHSamJV/T9odYDHi+UcocUw8
7068FIO6JQ2VL+nWwvew8F7qUeXAdKWqI2trptARCg0aEsMZlac9vfQM7K6oBrgo
Z9Iq3uYP1ra8uFxVFnPI54J2tM47pjT1HsqqfLWMyYi09yDDjMMM0tFInhdP1vnD
gtuHVu851vIxY/re1rF3jVFAwr0heZXSvChWqoI7Nix8z/Wmya7bseNQ+k/e8HyM
t7/p25qOe8wuJfFYlYl/xYk6pVH1TJ/xkUHtiaC5cxJDayaUJPibDO6JOrlElJ0q
hc8ADM4dMzhMjPb7spHnWoq6tqD9RrktMU/JCdfgQyozlBp5o4hsmEBcUvMKnVnX
ohPNM2GFngJT5+GtQQwfsXLkxfBe5HYoNOnKCnXu0tAgUlP5il/cY+reZwAlyY6k
BRDTUSmEVm6ayYOoZlCLa8K0tko+uSLTtQH09KymcqMdlhjG7ULyu9TfxmrrHGBN
OAFakTel3lfYSfS2F/aL50mTHe4soXfluQXPhq1A8KQhcfoP6/fAdnFbtAJb1+GC
DoZfYHby8f3AsE30tezWYwEAFQ9qhhfKLdtntJk9FWRBYMBqy2D2/G0QDCxp/DEZ
ncgY2i2jZuleKuVfjTbqhjUZEreGLJ2lesonZ2HKElWxfPmx5cW995vCSa6JkZ+G
HhMosCl5+XS9eLMMNrp82LZdI3r5tW5jYt2X5GQmGxSCohy+8aLmYndRFz0Z06xR
49TFszaqDV0LVidFyO+KRNwMQcy2FA/szKq736FBs+7CH9jMmSr95INLwf18CI4S
ZA3RqLSEJIHkA4HDhjGRRMUC7tjIhZrTSHK/BjwPNWtouMc8Bvx/bc5ZITxP62b8
EeZVG0TqfSHwnwDUpA4/s8WKZE42zZc3X2EdGPV4wySNdEee3T+9Jb8GTbC35aw7
6HA0vBfZYnx95yVr8HFdI2RjeHremWqqtsSKd91KGmXBl+IdGvsQSs8Ysk2ba4C9
kIF+ODV1Z1DYnjsGYCCTcBkNUav7ERQ+c6bg/hZLQWHAbMfU6Kur6DE+oNFd7N8k
5ZbwLUFFbVMi2ufHs9eKlQ==
`protect END_PROTECTED
