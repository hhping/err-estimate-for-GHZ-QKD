`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+CCGlNpGARSCA+eBi12lHDq6X5Bd26H5eTPWM2SB+WvJ4AD7Nqsj/0TFzGXT/ky
kGpgNk5GrxPmPmnNKudSlYdkWN7/3kF22bm3vfIXcDLUjdsAbYbh5YuGNoDyZv4O
FMmdgmIWy/6Ew7O11XDqQ4Y507ulAcbdKbO7SisO4HcJAnzSepp/Q/eeapEYGkXg
pgYjGWk1ZUAM6pU2cQZ3rWmV3soIfz2MILhf/Jd1U49MxB6qVfx6piSA3YbMhuBx
p+nTh6Eth0lp5j6AFa7X5x2/U9Vyvf/IJ2+8I/jT3CToWtCt/nRZlZIbApuL7ByG
xYVcOEGoHyetemobxDZSk0CeEC4ubrsosBiMv9H25/SuAXcUY4EcJiw9Yl9Abnqh
HcpnWDKKYvpNYxpsH9yxPaIxhiqMB8vDUCHtY5qCZbbFBnbNESD9LH+rg7wporZX
SF6Xk+5mlSxlFdWEEb2QWcCkMLOjQRElGoxGyh7l2neuz3NdAVqJHyKs66/O6HTh
oMGEesIx4vlse5ATKSL1t7UoZdIqP+EqNONm5hQcAkMiIOVrnWPcHGbQWZHbXxr+
O8mL2RiFFHaht3eGBOu9FRnfKy2i87egAVfapNBgwix3AZCNM3umy+PO7TAERzyP
/ftMiixxio+BPDa4Y2E0Smiqkml8kD6QfienE4hFmqe0u0YK5IC8kSO92FcGhi8H
7Lnq1TDBm4NXgB7ifRr9b7wK3jchaYefMu5y69kDCI8cRK4FP0wvrKKPzlJquMU9
WGTTnXTQ6XWxK48kZiIfDMnY8rrKItWErBpL2bGhrl1w2bWKjWT653BBlgRFwo7o
lHfMPf3iIjIs2i54USXyW01lsjvxpHKNEo19VHqkxSKPZ/9RhuCeVb4b8qXj/sxX
Y5lLILlXWN3SwUjXufaUJnnNVwRc2AnFiZ3pP+w/U/iEyuvx+mdCuYPvEunP9ZNL
g55TPlc4u9QdhFe5kC8khqKUrVGj9HXomgT5AUgaJE8dyDqn7DHf1J6luzkWWWYv
r2MXpnOlUq26iu8VoMtjrdLcjkNb1/WARitQTnrFnhgjwuxdVT0YUrm283NLTNjb
p72ZY5zr2geKUP6gA6+pUF5vYNPfJylnwLeWZZwTC+VLARMUL9RXGTD+4VzvuIEl
08Yarp1CxqA2sVROmQWki1VrFj7fe1z/SH09s3tSRzqZVgERJPSVUsATnog7D+V3
Py/EI3HSxXB3oOAtipGtMEtatul8aC/h4eXeNxFyRdYJGTQwSoF3Ml8CVcLCF73V
OTRENwapME4DSiJXW2/QHyjSBMwHbj3bqNYmRm0i9rDhtyOhBOQuuuKbNPFYLzCq
vD4o5ovcEdQscIQDHGntHxaAaYJQieivqJZ+EDxxzhtlNUZYON1CfNSqpUh2dISv
zUg+zjSjqJHTEbMMNBvm/zUPFbToS+t9BTF7kunOEOUPSrA4aKRvPH3jbggDXMxh
23IA6AFNll6vZqHhtFIWgtfBSP0gq6KZ86xjv791QdUCaBLu003IGZ+fRWE1motE
mG/3gFk/hPgqAQTKcwT/Cn2YgsckQ2CGit54MAGin8v38ahKakTDdjzpLGaXRy7M
eKAE3SYsTBNQWTRykU21p9GF793W14O3eEq3F1CrQokozEeLss9JSe21qYXBZ336
tHQt5M4N/HFtqLX4cq8fVgByCqMHDQulFPfQj22gie2wA7i90m/Q1j7YE7tZ7Ugh
kKFi3EEGizgVXIu+s9rrH/GjybWeE5VssGaWG4rA5eaO9fTSno8JyMiMGh1kz5HB
j2XwdiUuxQCdwUQAQ5CV+LC95iN/hniyOmdEIOXImbIcsful9gqWfts5EvuVSJzw
q4Ggb/cIQewpm1Axs7mhj6jPO6EK72Qqj/XtAaySxkp7G+1TU5jCJ7QLduGyNVMU
csbLLa6ftZQywZfHcBOLVIE+pPaKuZ1s3jIj7MfGJ0MmXhb5r+ygDER7fgNaTHQD
Z5RnEhr2FZFvDNiluTmtnh9aQxsm+LWFz7LGC75tDo8Gw5iJAoOx/ByP45zIhwui
msJBZMLMJtBpeVX4UQrTfywSzIvyaJmd/X0BuHubDZuCD5mnqGwgyyv8FkRh6kAh
GkprmGcn1PtA6CA8tTJhYvG8XD/6IerjVeqxF3CmBVyziqUL93KQ5MjCDwOumsfI
KGUBxJQfX5RsgvlrzBJnCewFBwonnrWVn4E2opUPfR9HI2zy6ExXG8BU2X18Szt0
wrjXTboBeUOY2DDFvSzjKLGK9/CtiXi05EeTgGXgT9/uVWsdLaWgIb3tybmlp6AW
xsRuF4fDY4oBw12sccx+XHhiBkq9Wu0VI4Lp3a8b63LkMYQTW4QN2lxFjM3X08aY
I6LTzxw9prSDpUNaOumX99O94kxxhMDjm3vCnJ0F5z50SxpTASuUJJTcLz+yBNo9
Cybv+wzeRzbMczlp3H1kk7c5BtPYL1C6KOpAFrZT0sEXCsBUeVphICubeU+HZxPX
bo3AHK4DJQhd/qZSG+/GCA8duwtRqbgzrVF3bgoK0sgPAheBJxgH5lkHCYIRp8vZ
kizjUsOWSr2QusikhE/KfBlQ+LA/EXcuLVYCJCXHgQrlgMIp+/TXuXlxBndi3aPT
8qGq/NQaichnDoZz5Gy6/jn9gJkPORiX6JYq85aiNyQsGue9UgP2pHH9Ttvt+FvV
1hwI7RAIvzGPqMXGs5Nw3PxVBakkaWoaWWegW5P0OYjmDloa/7mhLGnwx3FbikjF
3kJ51BQpyHnnk0hFsSYZloyUKo7whKdFxhAFD5M3tVk0UQ0+7gjT22kGe8fAKQdl
DrAHVbe8bUgNxPAxlPEhxmzMZkkRvHke5K+EAJHcO03ylBgZSE59KeEqzwm6bXGg
HbI11WMB5cnXCAiZgVAEhQ1Ph5ujQLEQpR1ekN0w2gl0XZDHUFBiiNILJTTYazV/
URHMddwwCIhPXR6V8owF/7ZKjA+3Bigrcc0IWwq/H8eaoKE4rZIs6Gi/0bDcraNO
MxO2JoicN8P3LH1avpZMY/NeMSE1I7Q8l0kL/1X1ubSiQ9UPeTE3A4eWT3BDDQvR
yqHDGtvo4TNzerkIzctT9pLwA4qtFUqJ2qVBA42YPNnm1yJwotfXWS6Au22H9GIj
Sf/COm7+469QR6ORPp6cC+uHBVj/hQyH0KQTvgPGxaiR44xm7uZy8sfWDXB24k91
ImYeHxnCPoYihFRl0URqAIg3eztKVJK4jfK/b1G+N2XV5BnGorJo+P9WVxBk3ehO
SldWSbVa7ECnhe0Sd2Gn68YUuhkI6/AtAmxrdIQhV1mAzbVZ6B/GaphtAAD+IM4o
EOLWsxwMBt92e7iJuo7TV+l0WAUCTTuHJVyeOulsnzeZ8+nwn9omLmDynfEguuQJ
SGjgi2VOHbPuyOZ0MwXEE580Ba+oDpdlTmZLmv2yQJpIH3i4RDykBdw/aBgIXVvA
EQ99oGecW9hYB5ZHvL0PCBcdPmqZ6RzcYdCgNrTMya6xSqC0i2oqJaKTjppmcNmR
OVH+0+w+JdTzUZFBj1PrRj/bqv2MI3H8Y1Zi/m91e46HSzwBMF46sclU68jyzTc5
bLt4UREi/2wU47/8qHizOceUWMbWYRdiIvEksMeb1/2M+nLKiNixLXWpQX4MQXlN
4FdALjPOWHQh7obsD8rb1TScPXZazelg+tpWNOs9Yi44NFsHctyKTKOSbfvx/wl3
sTayGetjf8SxFeZvK7w6C+mFM/MEJDawGkHeEBBGIFQCbRskgUhyceMkzEQWi/3+
v+MA8zE80Zl4BqKSCKkowcZ9ZfbAnIvYHpr+5xQ6zc6N5lPfgdgvBmymaSGaVe/b
zeQXK6NIA/gxCSGGQMcZlsxBqMZ8USJkSxx93MrZ51vEwOtnk8Z7iooyuORtgFnS
liuZ9fcT1HgsclgkGFeLknG+dRHtGOpkIEyGrmztNgGj9xqXfMIxdbGOyUvl1zKn
hwnqA7DXUvmKe3+xAVJG2dJN9DMGmcVSPTCmCHX3gK5HHPkpPk+F8SkMVl+keXvu
uNcxvgKNHCLP+6+1Os6MEZk791XokFk/Kq77RrQTjomkAv+hc6U6WPcTMfYMFiSu
OVQyvaEu0KOSmoD6LXnfeSvFU6TYOrhwReexTkfIiPCQlETkzxgwekoSOEjnvpsE
z+BpWY5dqD5hQ1LeUq5BUoWED6Nh+E++5DBEYcMiEgJQEgRnSz4RTV8nTMdu1ODs
OAf2VlWHKMJfEU9FMCORe0x78l80RWcLp9qBH78rs7TMXlBUmRe5w9x3W2s3aH4S
ziKWWNBTVIdc2Ekn1KD7rnC3Fa35PhFrG9pjNlf7n3sud579izO3/0zccjZzB2vc
DE0amIt1/rrKWz6ASX/EYI//O2MtwWwUh9sQV+OfuBSdeN+22a34xJk0DsZgINM2
34h+jTD26rqIPtHews4lIIXiXzYdC6qb+TVyfPyvZvGoZokZmS2ItusnHZOBgFx9
u1aE6bRFcZtwqrgI74eE8ke3QNY/fwWbU7PajTvV4e8fcRHUfjoxfwZyCHtS0ej6
klFAilm1HmPpE6QivlYQXdBRgarJv5DY2sJe4ZQAr8H3i9Ih8GKK6xNPLTlZrBHL
+WygubDasdStmdDOvWOq9tmLESRArkQixjB85eGWb+dUb6jtBuGFwyE+HtzyvNOk
IGKKtq+RxVZ1ezbxKy1LVp5MltGAWf/f/LC/vgKz9YKmXAccc4HdFb2Kg/IPIwQo
14kJEwTIqxI8Vqoks98GctmJRw6Uz1OVcSW43TEq5Ra1UY8iWKj+BZ1JDyCxy8ZD
Lf2T6J8/6QsF0czDXYtidFOIVFfGQ8cj2qTGQ/G4JUzfQf3DJauPZ9AvcOB1FzWn
+s3XAr1hocaZ13IwnLMqRX8LpQcj/+sLwVDJ3B9e6Hdjh4DDSexoEcOGLPoLSKge
iM9wX6hntUJGTRSDtkA5jWLW25M8vUCof5Qv3zkQcvkRGgQ/FCWrvawXxY6wFYpt
rU8kR0aGgbwOuBXqpf3ltPoBoilJoeK/A6zTpL2ogvZvOpP9dICB9+/y9e4Aj4/f
Wbwj/Sy/DtsUgLol0sgP3ZI7PEm0ze5eKqnovfIxJLFowyWi4bv9WJ3FOef/0vuY
f1C/LPtz2bQNjqQGMaJRz/5uh4MW6xACBAzgWAJb8USvCYt12QXMHvzfKLM1gbO6
X/6ttors22bKkHtjbjEcOarMi3RchxhfpcFe6njRR3AZfXQwHnYlWa7erh5icNFd
5Z8O1HSGAcL9Iai3foFc+lwGrtv0kXir0ABy0WczFtTUgrn+bqypAbyL/w/4yLyn
t/4vlZ162ihZVxx1Maib/MYZMDFLH4p3vMSyTSRSORUNU7B2VTj/sJQ1+2d3QQNk
B2oiOnWbo1Hz27p3/sOpfyi6UbsEWF7A9c8rsJMzvblqw6Z52DKl9uICfdFkT+DQ
FiRue3wgWvrrliRRAB8HIYzOQ7xaQ8JgnEXPXJCkbpSeapqWccRRph6/mHL/H/fB
IEQWxpn2EmWmqHLivuUcLEQdGQ94QflMPd1ezJN6sFAicgaJ5vR88RyHVRdtdMSM
uRhLmPkZ5lkIxgO0HFAu2lPyr336QYXkaHW0aW0F4AQZbigM+L9ZRJTAFCwtJXwN
b9bX0kE9fwUp0SqwIPAZVej8nQrvQZkS0N/7k0kv5rJRNQT6woeSDKh3/5q0vVSJ
GW9hiqcJbvQ42hanezT4alUiWSLc91U3J3WkWIkV5coxr4Vqp6ReDWwKE3NCOxDO
DRM/deqKZOFeIeMQKgAcWCFmH0KLZCK6s9isjLBOcyopXyhDxKEXttBcB5P7toVY
D6hwFWflchFrUrQnRnM9Maqf7P23fXs6qepqMF1nNcZwxYNBKOLIli0cy0vg1Pg1
T6JPyFHQM0at0BFs1Fy4GTLILZQsyj6irBd2yFrQKLG7EAd2w0cMv3TnPgDQ1Ne0
bE11O7RWRSN57S0ALzZNxwGaauuyBUBCRmD2tixDfsvBa0Rzskfz16ftPOayz/LM
BvLtIyKkEiYyLOCahVPAuUc+N8/kXGQYWeDUhxTIVemlsxQy+zkpwy9p6+toB6Vs
c/t05Ls3y28wyA3Td6RuQ2k5H5cDss69xNmG8iKK6Ak6N4fPGD92/cXbQUeCVgGs
ge56zxPREzi+omjyoSfbUG4tGinMn1OTKJKwlO7gWpbTAmkI/PCXAgYupAujFmZe
H6bYLMcxhgkY+kFp5JZHuYwwenAcnPdn2f4t/2Keq3vN7fOSN7ENP1E/Navi6Csk
mxInhgE0RGdMVVP4rnKl16efywRO17bD+x7ZjjiwZ7okvk0Q0njc7RV+NkAn9nxf
qDYiRdl7nJC8+3w4rB1g7SABMfeAs0kK+hdSxUkFEQpHuQM9ViAvvGw/1owqMfF4
wTZd+n1kGc45m6xdTvxyvhZtltsfGkua2TwbhX2a2l6EdfKbUzzWab5L0MQEa8yt
uuOgHrUiwa9tE9LdG4b/kRIqjVNoPL6s7JIw5o/mHG4mz9VG3sscv6pnBCxuVFKQ
p/EEmGN+Ms+WXWurnb8y0ISwwrwpGD5EMIMviTSMYad9UU51Od4NmFCpJrw/9fan
qN7KYEeGTG8NhSx8XyBnYP6u6eILo1I5Mg8j8x7u1MlkAeb2QkmkqdgYFFcnS14g
KX2GqjqJR+tyaMPV16Ofzo2iYZ91TUWBsYdAd408cL3rgPQ0/7dDJ/1Y0D6KsaGi
ZodB+N+bM2E+0CJSRCka0uI7QPxf48eim2lU735dXw9nP+n7UAcwYShgQjzXCjfT
JcLKSayWA9GJ4TsasBdgpuSkYBYDPzj2xp2nfN4tKDkJzPk9nmQw8AM+GO4Mlz3r
HeTKvlrT6+aTHnySnaN2vCDprr16IbX6KHzj1QWmTfAqXijxwIQpsXF3FWfeisYw
GrD3qdDm2TY9vmGt/FTMRet1kUWH0BdWUF91mPg1QqnnM6qhKAwByRe4P8bSsBKX
OHM+Ph42wAuMR5ZiSr5463YUsSbiTyrnRzbbZpOmO3QOBjvjJbnuECDU4TjKohIM
Q6WBMpTTHIkDgMCB+XL4Yjo93tAtWHsyz0olmGfl41AD0KfmpAiBIO56ti6mAVKK
ZfhpDP8jjOgWAAaR1LePYlX13YzuZqj8XRe6vAayBSsZyAflI6crNpnR7fgszbaU
qKk4zmQUdavFcEIvouDp8NJNsWyqspS1wcLGZzxdDlLIUXGjJnb1cQa4CTYYSpp5
s6SN+b9pkMXefhPSulmWpyNxH1lczSCtPc2RbdcjnSZbFcQPGl5vJW/LZmZkzXaw
aynRDNxYskF8BrnZQjMm0c+/RZD4yO57huuQkysKosD7akiEeUwYr0IcqELma0nI
v3scV2+s65cyvouFQj+OYMTn/JugSZ2TD+DcH4zT0llt+Z5gJ7WZkZHv85D7c7s1
MVL8ZmRHCRs24NhTsLVCLlAjvrQPdoEyLsH+JjkRfzhNu5TEDQ/MBAdSbvk0ngL+
Zy8Uij0UmljD4qSUGqdfkMUhqpb6tNribkofdLAfb9bh0j9AIloyk5dGVwVy4N+h
HTtsTEw/kHT5xQyje1zC508NLrdboEEUpJT6U4ROhccG+nFYKqAhssC4DWDRtit3
u0g4KY+qlFAAo5H635ocTw==
`protect END_PROTECTED
