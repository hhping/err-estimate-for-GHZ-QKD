library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_rx_buf is
    generic(
        enable_debug_info: string  := "true";
        act_isource_disable: string  := "isrc_en";
        bodybias_enable : string  := "bodybias_en";
        bodybias_select : string  := "bodybias_sel1";
        bypass_eqz_stages_234: string  := "bypass_off";
        cdrclk_to_cgb   : string  := "cdrclk_2cgb_dis";
        cgm_bias_disable: string  := "cgmbias_en";
        datarate        : string  := "0 bps";
        diag_lp_en      : string  := "dlp_off";
        eq_bw_sel       : string  := "eq_bw_1";
        eq_dc_gain_trim : string  := "no_dc_gain";
        initial_settings: string  := "false";
        input_vcm_sel   : string  := "high_vcm";
        iostandard      : string  := "hssi_diffio";
        lfeq_enable     : string  := "non_lfeq_mode";
        lfeq_zero_control: string  := "lfeq_setting_2";
        link            : string  := "sr";
        link_rx         : string  := "sr";
        loopback_modes  : string  := "lpbk_disable";
        offset_cal_pd   : string  := "eqz1_en";
        offset_cancellation_coarse: string  := "coarse_setting_00";
        offset_cancellation_ctrl: string  := "volt_0mv";
        offset_cancellation_fine: string  := "fine_setting_00";
        offset_pd       : string  := "oc_en";
        one_stage_enable: string  := "non_s1_mode";
        optimal         : string  := "true";
        pdb_rx          : string  := "power_down_rx";
        pm_speed_grade  : string  := "e2";
        pm_tx_rx_cvp_mode: string  := "cvp_off";
        pm_tx_rx_pcie_gen: string  := "non_pcie";
        pm_tx_rx_pcie_gen_bitwidth: string  := "pcie_gen3_32b";
        pm_tx_rx_testmux_select: string  := "setting0";
        power_mode      : string  := "low_power";
        power_mode_rx   : string  := "low_power";
        power_rail_eht  : integer := 0;
        power_rail_er   : integer := 0;
        prot_mode       : string  := "basic_rx";
        qpi_enable      : string  := "non_qpi_mode";
        refclk_en       : string  := "enable";
        rx_atb_select   : string  := "atb_disable";
        rx_refclk_divider: string  := "bypass_divider";
        rx_sel_bias_source: string  := "bias_vcmdrv";
        rx_vga_oc_en    : string  := "vga_cal_off";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode";
        term_sel        : string  := "r_r1";
        term_tri_enable : string  := "disable_tri";
        vccela_supply_voltage: string  := "vccela_1p1v";
        vcm_current_add : string  := "vcm_current_default";
        vcm_sel         : string  := "vcm_setting_10";
        vga_bandwidth_select: string  := "vga_bw_1";
        xrx_path_analog_mode: string  := "user_custom";
        xrx_path_datarate: string  := "0 bps";
        xrx_path_datawidth: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        xrx_path_gt_enabled: string  := "disable";
        xrx_path_initial_settings: string  := "false";
        xrx_path_jtag_hys: string  := "hys_increase_disable";
        xrx_path_jtag_lp: string  := "lp_off";
        xrx_path_optimal: string  := "true";
        xrx_path_pma_rx_divclk_hz: integer := 0;
        xrx_path_prot_mode: string  := "unused";
        xrx_path_sup_mode: string  := "user_mode";
        xrx_path_uc_cal_enable: string  := "rx_cal_off";
        xrx_path_uc_cru_rstb: string  := "cdr_lf_reset_off";
        xrx_path_uc_pcie_sw: string  := "uc_pcie_gen1";
        xrx_path_uc_rx_rstb: string  := "rx_reset_on"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        clk_divrx       : in     vl_logic;
        lpbkn           : in     vl_logic;
        lpbkp           : in     vl_logic;
        rx_qpi_pulldn   : in     vl_logic;
        rx_rstn         : in     vl_logic;
        rx_sel_b50      : in     vl_logic_vector(5 downto 0);
        rxn             : in     vl_logic;
        rxp             : in     vl_logic;
        s_lpbk_b        : in     vl_logic;
        vcz             : in     vl_logic_vector(27 downto 0);
        vds_eqz_s1_set  : in     vl_logic_vector(14 downto 0);
        vds_lfeqz_czero : in     vl_logic_vector(1 downto 0);
        vds_lfeqz_fb_set: in     vl_logic_vector(6 downto 0);
        vds_vga_set     : in     vl_logic_vector(6 downto 0);
        vga_cm_bidir_in : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        inn             : out    vl_logic;
        inp             : out    vl_logic;
        outn            : out    vl_logic;
        outp            : out    vl_logic;
        pull_dn         : out    vl_logic;
        rdlpbkn         : out    vl_logic;
        rdlpbkp         : out    vl_logic;
        rx_refclk       : out    vl_logic;
        vga_cm_bidir_out: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of act_isource_disable : constant is 1;
    attribute mti_svvh_generic_type of bodybias_enable : constant is 1;
    attribute mti_svvh_generic_type of bodybias_select : constant is 1;
    attribute mti_svvh_generic_type of bypass_eqz_stages_234 : constant is 1;
    attribute mti_svvh_generic_type of cdrclk_to_cgb : constant is 1;
    attribute mti_svvh_generic_type of cgm_bias_disable : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of diag_lp_en : constant is 1;
    attribute mti_svvh_generic_type of eq_bw_sel : constant is 1;
    attribute mti_svvh_generic_type of eq_dc_gain_trim : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of input_vcm_sel : constant is 1;
    attribute mti_svvh_generic_type of iostandard : constant is 1;
    attribute mti_svvh_generic_type of lfeq_enable : constant is 1;
    attribute mti_svvh_generic_type of lfeq_zero_control : constant is 1;
    attribute mti_svvh_generic_type of link : constant is 1;
    attribute mti_svvh_generic_type of link_rx : constant is 1;
    attribute mti_svvh_generic_type of loopback_modes : constant is 1;
    attribute mti_svvh_generic_type of offset_cal_pd : constant is 1;
    attribute mti_svvh_generic_type of offset_cancellation_coarse : constant is 1;
    attribute mti_svvh_generic_type of offset_cancellation_ctrl : constant is 1;
    attribute mti_svvh_generic_type of offset_cancellation_fine : constant is 1;
    attribute mti_svvh_generic_type of offset_pd : constant is 1;
    attribute mti_svvh_generic_type of one_stage_enable : constant is 1;
    attribute mti_svvh_generic_type of optimal : constant is 1;
    attribute mti_svvh_generic_type of pdb_rx : constant is 1;
    attribute mti_svvh_generic_type of pm_speed_grade : constant is 1;
    attribute mti_svvh_generic_type of pm_tx_rx_cvp_mode : constant is 1;
    attribute mti_svvh_generic_type of pm_tx_rx_pcie_gen : constant is 1;
    attribute mti_svvh_generic_type of pm_tx_rx_pcie_gen_bitwidth : constant is 1;
    attribute mti_svvh_generic_type of pm_tx_rx_testmux_select : constant is 1;
    attribute mti_svvh_generic_type of power_mode : constant is 1;
    attribute mti_svvh_generic_type of power_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of power_rail_eht : constant is 1;
    attribute mti_svvh_generic_type of power_rail_er : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of qpi_enable : constant is 1;
    attribute mti_svvh_generic_type of refclk_en : constant is 1;
    attribute mti_svvh_generic_type of rx_atb_select : constant is 1;
    attribute mti_svvh_generic_type of rx_refclk_divider : constant is 1;
    attribute mti_svvh_generic_type of rx_sel_bias_source : constant is 1;
    attribute mti_svvh_generic_type of rx_vga_oc_en : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of term_sel : constant is 1;
    attribute mti_svvh_generic_type of term_tri_enable : constant is 1;
    attribute mti_svvh_generic_type of vccela_supply_voltage : constant is 1;
    attribute mti_svvh_generic_type of vcm_current_add : constant is 1;
    attribute mti_svvh_generic_type of vcm_sel : constant is 1;
    attribute mti_svvh_generic_type of vga_bandwidth_select : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_analog_mode : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_datarate : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_datawidth : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_gt_enabled : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_initial_settings : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_jtag_hys : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_jtag_lp : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_optimal : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_pma_rx_divclk_hz : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_prot_mode : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_uc_cal_enable : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_uc_cru_rstb : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_uc_pcie_sw : constant is 1;
    attribute mti_svvh_generic_type of xrx_path_uc_rx_rstb : constant is 1;
end twentynm_hssi_pma_rx_buf;
