`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JG6prAg+O5/5uPzc25n1WysgVwEowQNpP/5W6JX42znUI00VugdDNIb6NSfOjdRc
12XiibtbuBmj26y5zOKud/IeDDM6AuzazMIeTTUWnuJdDzUzi3g1orimoEE98XUu
RqRUXMIiAt8BUNbET/XeqqngKSLDG5Sw90cUtkjsgxEJKi0ETm0BncQHar08cm7X
9n5wA9usT2t+E58uiWaB6PL61oxZSk4WPS0v/4xGrh8LFAmuZy+Xak8yrZvMTwwk
ZnkVxZ8xPmSCl1L2WdKgmbGwCAkKZclgSP/yKfZr0u+tD4dXzVUVACE7wDlrDxV4
71LwugoaMW1WkuohYGAQFG9jVm18918y8t0rGlb7Gg2MAAdVjDJANg8dCAuBF3Bg
MIj63hT6gPEQ9q9dR9+X3kPnf6/IQI+HZ2oLBR1d1ZwVhp+qy1s0wfR0Ao0z+OoJ
5mNwyGrmtzx1vkpqBaHs7ndZXiBwQZR3lAggK1F3EiO1qGQtnGMLWg3TM1Dlt0gD
gZA1qjQkzj4HjuybT4rgQ5C3HRm9GPJWE6iIHTF1Hafi+zdDaFola7EIn1mVEN7a
3BL5gVHhtuS/F+p6VYSDdeE3fEYmatNDyXQ794M1PDGClKCa+1JsEJlcG/0/mADb
UGErbm4Vwi+UgXW+1KkJubVL1rw+1qYMM7cgCqrukJ5hLKosX8GHM7+aZqS8vw8i
CBG2y8vcKVnC8dAhs5m4HAZSGI345VgRqNdVdhiXrPo67G/HZQKTnFUDxIN/YceS
ZGDUTIifaja8DeMgFqoVNHcKdhG9a/Si5nv/D4tXmQc=
`protect END_PROTECTED
