`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r80zWNsusMyFBYBpdIP56EVjuy2udjg4V5OzBHFf/RPy8PVrz4iTX1hqLPt2uzKu
/6aKPtscIKjMjBDkGdPMUXTIngipl9JjxWpgRhkkdxmzcjuWf76zDW/rKaPiVWz/
hZcPNjTw4u3LAB7J4TMus48cbS8Cv36HhfILFBdegSdR5+waAbpjuyEiHO7bDvl7
LSGFSAntTYd5jlYU8vfeaX5W1VzO3YBFhy94m29vEXlG6tArtjxxl7pcET2zPOqi
a0yXJLIKbXOIJPd9hwoGu9BP31ADA1r1ays7AdNee793lLWMrnUPNbyqChRjHB4g
D3ONWDjSjbywE5ZrxJPtSd890EqzNrCdO0A+cG9FzG/NfPHC1P6M5CNgphZD0mz0
Lh4zg+6QUbyayAZG91LlVDr3IlDkwdR3fjC+gcMrEmbM2Ye3BzFN2GDYS+VO5iRz
YSdJjQMPpj8QJbLHM83VNCdP7CMoT+uCU9/127xJc+aXVt0zw0a8gt24SgFotUR+
lB0PF3xKFTtDNzvM//dI0NuL96NqT3L3PyuZRV8kzt0mM5Otam75pJ4anp7r2SxR
L3shg+DDGikxCnGBPhrlYNFzyuNIRp1iGkpuCUhNvA+vdKMsol944JLn8Nb8lT3y
`protect END_PROTECTED
