`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTFqsH0dnLi6gWvXQdYppcxhna/Zj2VcxYIcV9vbS0DvSr1L2mPRDGOXKPDAPVB+
KkJfxI62/xC7DJ3jqnUjy/XRxxjXb08M/ZglKqbwatoNfwkPu5T0ZFSU+QP3x2ou
yGFdqdpwvUIszP8QkzKRaU1fmpCL/hS1jR57bx7R5xUalN9RyW4xCCE1Bs8+5e5k
i7X3MmJ7PandWEPjBVjGrAdIAyfYdFLaILJXe7Uft5G3pmL+sxHi+zljyTmqdzb9
L5Hn8kB+MbRUykitRauDnJdDvCeAOFf1q8pdo/KRkcj/XtmMj5zkszpvDyVtKrGw
YIgpLyY2Lfm9xS8ISvMz6Fd7awtq8Qyf6PfKPb2dKGb0eAVpYqx0iROTPiUpjZwV
JIzK8KpdM3qL4jafsqzYgjOjLvQzD+RNsY3A7UWHj+n3Qpej/HyWr/I20WEv7xRK
yvMq58sJiq7firjFMWRz7qZfZXzo79BKVRMgITo/NdxhWKhI2DyDHCk1xzAhxt/i
kJ5bkaI8TMDspg6Z0Dp2mFFFNtzSXvTE17OMqr5o/se6un6FF7gYLGEmkxepCDps
IbnTvGtiYI5J9/oICwZFBSjFb/0Ox3djPCH12nBctwhwVy+0/YPXnotiYqtejUoJ
hetHKLPjtgMoEreZcldSXoa74nk5rxKeh9j67I4NcRT22aP0kDFENJf6JUmPeKkE
VhjKebj5Kk89x7U0HzJ/sPkTN1b6Owpc3KPIbgTfYbbJPktZpI6FYDsoWIJDng5Z
0Y+2wQQiBh3z7GYjtBM8P5VmbZHxP6cuIrlq21v9kw8/H6rJ8mr+fgAH0rhUwRFQ
`protect END_PROTECTED
