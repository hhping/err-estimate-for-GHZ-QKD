`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhQPmEZ/faU8nxJp+fizHtd3UQ29B9L9ceAupUvjDwA1PbDX8oWz7g5lWW/yFjdI
xWgaHVjAurROQY1mVMtKC7exhVueQXhBnmKWEytxdRUXbVC5VnkoXy+Yv9PizwTI
q4sPzLA58JsplTnvoUwbxnYfJpWLLSjpwOfOFSBdlY6Dse6rzbWgW7oi5oZZcToP
rXtr0OUqUHASJENZQKvxsZofxRtrIeAcpCkmZtiStiur8VwEiO2bR3F8XVFdLlFC
3yRPKdjYRWBCO76rpBQFw0Hdc8jsxppnTtYzUgKEK490vvasr5iVV43k3b71J1IH
LFf1BwGegOrJcuuQIQqpaITsfKzHyeeC8kOvQxqSgh5MJ+mTbA3NEOhXBK/ri7k1
qUp829pvIl14SfnRre8CXS857g4TnNHcekh1nrBM58a0Eb+ARwgpi2c7ffVqwMLy
GaMXdNBF0FVDjjKi4QfAmIXqUWbjgroYuKEfamLQHrKCcIJM2mzpJnm8cvYJSw80
CZra8NywqH7OAaB3MF+N/K6S06+uSnu0jGYTU+hL6RGynOcZOOMaIwb0fR26PSyH
QIjtll0dmZGpDxA3XechWL5g4KAvfIvwxlAxAMdlCaaDDhqEI7lEOzsxVs9ptRqw
2/F8HJ23g56jPIkzziZS7tmwumSi2BbSXq1fkpK7tjbABNlKPWf9uK6kRvUhO8bb
LfF5CzDfpKJ4UdzI2T1LJl7WZs/vhHovAiMWssNnaMuOldN7DnuSHGp7nvIRaToi
MHa/DM3MEb+W2S9koK438Q==
`protect END_PROTECTED
