`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6m7uugHrSSVRmx5fGc1RBHrvemEV6zf18OTx13/H3eON1qtMM9de+fg9fdaWEyG
NI5dilE/LU35wgqCFtTWzFqI34z8RpGgGbxZVWVqaz1F+4ruNRidmmjtlh+lZlww
FRsenDrvtCi3qxjXRGjM6fK2jlJ1jGSAWIPN5pNdIbRmnkrjbaUkSso9Pni6xXZG
Khb+BMbYESN149Y7mkaQHRhU5ftQ3wufAWmV2Ge9dV9IVjH8ubPfAA4jFdyMzK4Y
5M/wkjHpm/8PT+iVmkDZ1jNMtEdM05bT7xT/f1c458oO9XK5i6HhFPZbFxRpwSL9
k7LxCQCJ+rzQ5EoNQ88XcdtWDiIJCryRvPvlsUETC7Tro5DUqzEHAuYPLjYQlTmb
YKciBfrdVJ7WPESnp93qYRyqUD94GpzUWAqoDyGliL+HSE2IhHHBHcxewbgy3Zvl
kLZPZ0lNOT7u8L4C0Lf3aZFVyWp7iXFPK94voLYlxH3fClf5weRyg9NeaE04wqR3
wXUqIgseGxQhjcjDM5MSMgd8uFQm4hQ/qCiQ94a/xssGfVNUzR3tHU38EvUxly5/
/3uox6nQy2DNgSZkT3BWjMvZs803iPbeOXKjdcoJEV5uZFbYnUjcjohQ7QVLzLQP
bdpK6OVQmXt+yYdNeNZ9YDmsIOWGNZ8ArLV/VKIgh0rWof/m7KTZuxa1RNWoIlwp
yJhCPrXK5mhiyI6zaDJZBm2L7/iFa4MlzWj8kLH+cLDp5op1SK6NGZWSzilzvtXd
pKvoMcQGVC8pMeiV+gO9e5h5F9EXJqS632SC32WUg5RLYMboLx5NvBTjtLAxnI79
wAYFslisnDenNHSxLWtHvxKKatnJLnTrommyCd3jyjc=
`protect END_PROTECTED
