`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kl7HXH3PBN3+PASUocKPZGckxAURFLjTRHC6klrGNo43c4gnDhnMUz+m0hYAMxPg
jyvgSFoJFm5qwf88AnWa04r6unUmIRWEdPJJKz/FhxIVTXM6MxCxYATlvIfEvpmT
Z8fdQLimzQf5NGraA2Zwkb5XQqkwCoR14LghlVesaBg9xwTi1kONrhdZgLkQoQLE
oNAbknSMy492bD2cXCqCFJjNU+uWbyZZtg6/gh/1qGLOOtxTxKvPtXJ4jM/ui8nx
5BtO68M5+vL8f9hPI9lAMbkw/7Lx8a1BTca6xKud+7/i6K7Y0j6F8vPGk6Ytc+72
Yr58vFpgdx5lVRhDT4hqzLpGg+pGPiLigxckwIe8ogLMQlDSGdnN/C9zYjStiHDa
3e7gSRxneGdkz7KdGZ/yhYSbyKJ25gGSAN8PNwGO8vjBqusETfbVgl9xRE8CSOuz
p5H9PJAyupubOZ3LdOZoiu9s2bh302tL4zCnTnZCpOh2NiiUZp8lIRb3txQNXEqm
Crs6WbUB1D/kkAV7Q83vFy1UjfXAlad8/gjGLWikmh/vZSgpDAbCCpd5yhxvoqGc
M6DJ/+3ENCvNFZsxSOsN4mX2JqNXpYSQkPd6gko9OxZNB1pXIbvwUvrnJ3eP0Lek
BROcnFqqnEGAEjuwh+ZYwQ==
`protect END_PROTECTED
