`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFGhV+WC7ITSw+gg6I5sjzsCgxJGonnT5cFJsF5Hbh27JQV4IBJb/2jDR3XlbPUU
+5MYqHKvN3sB8Vucr2M6FeJxxe9vdACmTKHfcC6SBgmrsn/DgIDmEd5yU5WaCmGQ
nHKIxFeGh+radOBj/a104lbJA6vq3B8axslU3VWZyP+pSxWEoEPOVcvadTawIJMU
JDPPOlTbEobYVp0mI/Q3DuOR4MhKykkNZB+nSw80MHBd84KUY9++WJMAKlQ7PJA8
8DBdUMQJlxM81IMoDKty2qEphJTnZyCfglQEzykC56Khy+jpfHVSFmS9GrMBjQu5
ZT2yzt7+gFN2MVnzhFDszQVmHmeDw0I3zaS+alKvLSdm2oevj99FzFbjBPp/DG0K
/pRTwbbRyh16iRwCssGlZvV4FI+rq6R1PCbL0oz+adtZ9UxIDyLO7gfPeDvox6lY
kycDqvvbYZ+bJVHquqDuHaZDObCWinu+FpKfv3LlurSqvdCJwIMbJvJlHBaYVnoS
Cl8RYbzl+ElN8+Qm1KwFHuGskBvrqiYg9D5BM+h63pL6dnYI02+JnyDDGlTYTvGs
/N6yZdZl/2ntyO77WtlhNa0W2txiipM/7wKK9Qzz4wtxl6dvobRK8LvnRutdcm5b
ca/i6OfU0OXtJuWieB6+DZQLmt28y5fE5LF+FL0lIUUzbz/lO8rPQicZKdHvJ+dw
AJupopRDlUIiL2cdgv9RdOX/ywPbB8KjuYki6n0OwcujW7Lztu51uaU8o6cKnBbD
rrd1jals7PKzRHrIfqN6sVuJN5biEw4dplig1eri0T0pA4txzyqxAdZXJlrFvRke
5f1pq5Go3Vk5o6G7aNSrDUf0BqjjZZOpP3oAXw0tl25XbGnRr6oGpsXlHa1iGbyf
tSEYMa+hZke5Qju7vF/CJMt6gLPRlYdMiaMlDsBfo0xe88FovhIcZWSu4NLce4Xo
KjFcGSGQTNxri+siHNuV13BxuKNIIjOQ+J7xZRTKvX6LawbnyqVmurWKcr3cRxjN
ziICKLM4+HKsIGqWSkmqmejwFKy7a/15moG6tvvoOUmxAdRr1AVmtkA+fc1FzpOe
nKs/s+yYUeGUMiif/664V1EoVWLJGG8CaoDKVfhR4axEY1THu8mc6sq9W9WgIdPF
0R79xQsr/WYFsfbRoj2HAjC3kCFNS6nKVkOco2D8cnM=
`protect END_PROTECTED
