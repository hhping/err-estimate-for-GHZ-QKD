`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcEJ+uZc7ong4Nv+9HA0SCDzFEFQZRwBNwJoMRYp6B0uqMCPpMSCXfoDAhFbxXbj
UpwYpocLbGe8+h14IVhvN9keG9o0FaK4bYixI0y2d+pEDkhz0IQbG9kx6kG8hpKD
PpjNHN+GFPNFDMbtF72WNibHzdl84xSfJUbtHl2en2xk6zHcyZyd+vekor5vsGkr
wHXsQZmqZ9hqrvfvXKL/fOXLNhLNjjTBcgPtcfv7SszaKZoyi3lFw998UieqZD0v
z+1dgrjEqe7+cXGAKKDVGNySXvW/AnIv17TS0dXfxa9Gb5DcgCfr9GutPbksFtuy
/FG/fcrxBAop3FDigrXYmTTTtMTWOUNgX7gwCr9nQIdb1sBjxr2XB8gwq5QylyFr
K5mMZwkL87bVDnxdNAupYlCiBKQi9OXzY6X9PYszfWe92PsgUvzF4L1YESjJmFiy
ZsJiAdq50zK9j+znoYZHMqTF+RCbWKpKoDbF2RSUp3bKGbkICkuxpmVjzTmAX1KG
RYRuSkwIL/P7kT5X/yLglHsLbQpAhLY7ZSNBbZJWnkk=
`protect END_PROTECTED
