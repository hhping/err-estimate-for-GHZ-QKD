`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/FoCvAK34ldJevAFVzLro6rfELdE2994yuPmsSxGCm5p6G8Zeux7uNs/PAYibx3
n03X0PalIPGpIjkHdIZ7trpUS+WKRjuDewJiVvsA8jGv78Zd/6k+ChqSOLdYSAC/
gy048f0Q5OwUvNsiDQuolwL/4z8lqnVla+0Z8M1JA6dbzRAdKyqeDWxXFhBuyMAU
VR9DzsPK9guI2v0YSciCy08AZRJPmdPr211EsmvkSygvcj15iHwMsKMwDjLZhJB9
9BOipOcF0b0YlspbDReFCNUMFuac6bWqzGc2NsFJiQO/jsq+2hduIK94blAcnf9m
H0WrkSTpFokeejWNo9krnFUfM/YOco1v80JtgSDx9Qrvks7DtVYo01HOwAwBYGwR
C4bC0xkdgrk6EdMwFu/Z+uEIiKxnE+lwdgolmxM8EvB6Odeu2VWJ7boazIj6C7CJ
QHApddELsnV/fi6hY0i3E8pqWJlOtl/Cc0CpjDOedNQ=
`protect END_PROTECTED
