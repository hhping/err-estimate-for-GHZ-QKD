`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eugP72296+v3F6LOXFROrV4giK7L38WAdiGyxfBXmyNw4JNomNhoAvmhfy22Pby3
nu0/X7V/PO0IqR7MQu28FAe826m4NALLn0LlLfOWfLM/iKdc3JfbupkluoNKuGVm
VK3UPxedXIcIaLf/S1TMzPARLPxkQj7/Qw8smxtIG5azEy0ufbISmWyTEtVujrfd
ThjPRtFZ+ZT7RrubAKFmfIijlWpv5nX9uSEoDP0cQ+bXtdK6OfmDVPNdQcac1TBm
SpRA1YFTKXX7W0fCd3ppL5iG7t+tBmvtGkdglNclcXnB1wgDqrhg+dYlLcSli3tl
ryBYB5bnOF9PPwNntTYcEy9ofKi6ursCk34xjZXbGTSRweS9tdA2+0+VO2RzRkxW
zOUzHJbtG+PrmLYI28fAXHQxFqdMwG5v3GLSUhqbzCMuQKrZpPx6tD7sQyw3uLLx
EGr4csju/XRBjreW70ad0QhAGAi+4BqNq2GhemxRJD4EQsmVQYcR+8Mzu36sBQeI
7IGW+hvou+Qque/HWHIT6GRv7G14W72kd6kJozAki3j/HY+r83mKAPwDovZF/Kur
cEWfHOgP/UB6xtdCEmWpWrgwW5wVlcU2vwaBirTnmW+qCzqzTlNh6LlthsimoClZ
5146kzO9DGl7p1lNTUIotp4dq2NYfXisLq0NV8Xh144hBJYfWP2qQGXs5nULTPQj
ACGg247OUBxZN/ucRnqRjGlSJCZNsAJ/CQzvNaZ11WOszzjWYaYsgO8SW93YgW4E
v6sXYMtsMecZJqwDI1JH5w3swN5GfCyTiYRxwE+IKWLTeh/UnujcqNiFsSdFDE1i
Uj8S5k4+3XNc6Pyk+SJy4gCMLf5t64515slk7ZVHBT6hAAyOdfy9sN6ivrrkIzbw
FpHKN8joMbK1eK/Zg2uh8ckcqa3Tl7AedAiFgnl9q/jaeYLJUvODqaowrvnlejqb
Iykec8wuVbPzBtcDz1OPm1wDZC29Z7v6x74E0f0xWOk/4gi03v7Nap3+RAX+PvLP
UhbQ5GT3R/xjK/flJA0D+ZXkFRUKMknygSdrAQcB5uRch5eGFAz7bGTxBw7B4VFy
VNPRjpSh9kS5bkH34FH63gspJrFwSvdDpyiHP1jN1vs2epi5RhFMgTM44z3o/1Sl
8zSEbI19VZs5r+QkWO+TqaKVWCZQCNSJnt/aZr6hurVhO9AqRqKw6QgmJmwO6LmX
XDIQiWrlPouzEURDBsktUZtROZQ/d1kWVzIFuczv91BA7yqZ2x0dCjalWWTcFr4+
kqpVh3kDAoWcQ1FNy/lyhg==
`protect END_PROTECTED
