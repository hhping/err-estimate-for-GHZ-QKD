`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/cId7yeHkyNoreHNymGZ/jPNgNgqp5EPzLkafl7NbmBlcZdI559yBWbk+JNI7pi
dKnZfJEAVURw04EZBlJDNSkcPNpp/fcBcsI8UyAfxo1uoo1t8/ct66qHZOo57goT
Ke5m5V3DvadW2lfwGtqSkYC/x9zzyac2lY1VY2y2xyZMw77TzhD1OTPkYK39P+jv
YcCubaWw5Fp1vsQVx/vBn4IFeImDNE4IbfB6CbK5EvdwFe5N4ZPmYaB4EtgjwsIV
RjP/vjnLcw3p6tXtUzzqfpJJ8LdHAkEy/Gl64rv61VlIk3OHpimOSg6r+9D0hjR5
Xe5A9ud7QvZpW1Jp0hOfEWhJYrCJP+cO35829rb36neOOx0LbMMBQ/p5bUAEaWxK
kHTCjZilTPjF/o84v7wvg+D1EZe4zLRjW5GzyzeG3+z2UaymPbG++2GZcF2CodlV
LNPsUgGkYU6VHqitSox554qdMneL1+WElF/pFV40/5HMAHFfXvExH5lBk/mD+znT
gyvHjwo112U4AepeEXE8kr0SS/GD0JxEoeKV/hVXVd7Sp5tEBX2h/D7dNUN0HTvT
sI1pI5ExT0mf5rwmpVkDTw3ujKsOOEsNa9hmFH0gUqdV0/5e0r/PgsOJ+s0SqRKu
Jml+HEPlcOzvp0Il3BINHoMDBjR1UmoRy6vXQnL7znqdCHxqtEHOagZjbc8Fkaxl
iTSuTgObRQHo5zKaNaZqFQ==
`protect END_PROTECTED
