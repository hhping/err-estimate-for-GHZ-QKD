`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXu03R+5aW0EKEcYUzSdtu2KiNsTF9QTz+f3Zskl2YkD9VWlvtWg1juEkIuMnLtS
06XdKrMBqio5iArOXAok6D9dyVBme3a2rhYoaATGUxcSu3f0edy/Wyq42fHdXI9w
cyEoVqUFyuSYb2QVlg9G9hsBrnLfAJmrUQNPYllBVpcP131jiy2eoQ8+n4GlIBjO
Lib7oZbsTpNkdb5diWJ5SoZyGCZYdAVUrMRAYtReJq98e3s2l049xAMepiuoHyGA
6QRG1JdrdKM4PBcpIUZh4duL3qQAqBi2LRjcLORAgEt7a1P2HFHXeLU/ebiuwcdI
oFN9qu+JElSfh6lcTZYxgwaDopXyLo+YHBpl26S9iU05rm9lIkjuqjkwsuCccZXL
gkTPMCrBLh1vcsH1zya2cmAEd5LdRF8kgKnmRS4ptN1C85DKDyFdHABTSQtr2aty
Jp1vU60T5eIBDUDQq2S+WBgqKu8ZGvr7tHmfotPpuzUjhPAWEMzeLKWvRIpeodrj
NjlFmyKht9L7A0H+LqJ+AId/mLraI5JoCAVw8AhHaXHqxBHFi06llZta4rAVE2fg
63f3FrkPY5uqFL+GLyZ0krCf5Eupt5QAhb93dHpsdgmo43aOAeb4Uk6WAAkwp3ue
Irrfm8Oj0QtlI1ODo3RcjPi7Upp95C6SBCQmoUOAjHlQE8jgXXvfuDWiO7Eworr5
RCJTXkNu1TP44Jg3/uUx1+DNzkXHuqUZvq5NCM5iXcuVuDs4RKVu9hH8ijKp7x4O
9bYTpGqj0MlHEQrmwLNZrAQ3PVJEv/e0x0zH9DcRMyxdF6wNSH7F7+w6dvg6UfNu
dgqevfnvTXdeddaXFcWIFN5fS6MZfmyE37pzVsZisqE+ZNQ+HexPyX6TxazrPqTD
Gsusm5CHgA26Vi/avaG3hsfENu7tcrZ6EXH5LezmhEcf026o7ptJO2s4NZn/e2Se
t8WDXC6bvtMRW1MK/llWUwb5RfPmehCgVSuTlyaRXtg692fxC/IOMVegpIK708+B
PX4TQn51ux0FnMkiOP5u8MDqCEBEVTSVEaZuImNoPMxb2zvozpfUrCTOwrZT7W4W
/DnsNCpEFfmT+8ZOb4H1OK0RMzEDZk+b6nA26FKPdFbGSWcHMh1MjIZ/O9dDk2Le
w5PCZcpaHwTTUlyBLLBRpYBetBZyf3v+UpIPCaOhIIj1c4uKw0vYqxQUqLMNSOLC
hTCAoIHDmSEfeZ46LMiZYo8bKdXDZ6WmfX5Z8mtYrJyrnFQoKDv+Q4SzuMw4j8JD
nocOf9vSSw5Iru+l8Ccy98/pIHOkl4FOyGn5qzCpbC/6QJYk7iRfty1YUwntabwA
MY7FoIh431abUIpb9Ua61h3cZihM+83c6kLoQv9v4dnonLxMYFygjZFeqODi5E4k
Dtb6obSMAdPYSwfBmReunr67F9EFUPMnB9YAqZGyj32VTaX/K3zD4aiaimm6e+fu
lipEPeE6P7FSXeulaGzkBSf6FH9yiGvwzCNvUETqXMnWkPIaiKaM7ZGKMkEXLz7c
q6wIXQZUPT7/4XxvyVAwP6x5aurD6jv7G9Qzu9WpVIUa/3uBL/s2BsJlSZYyYbYs
8JXPcNe+gzd8JHCd6s4VBr6Hkv6HK+m2DeDN5a0pjjLsRuoXyx0QtrEeZltLKQ3H
/EooCSbQigSKlT1OyDYIhbMECC4xonE6YqlB/xyoCNVQUVXlv21ytwPwACiDvCMC
`protect END_PROTECTED
