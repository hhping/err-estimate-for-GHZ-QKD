`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVp6D5pPaC+ORAsCCuNThj/WAhH7QcI2L4ERivA6kDijUAxMhEAEZ4wWWpRowRcB
ew7HLtrM6JiWuqJPBXSFfOuSYUnw5K9dMU4Ny4hxU2+ssUUYYFIHtg7q9zG81SF6
7aK/hHRA4e6ZC9xzhPprM2YXbD3M+RWcodErZXXyGGoFfeiGzkN64B+vKRlui8NR
GAw6mLtOBKPT0CxvGBgeZaSg1xNPmds0PsXtSC1yStV9ace/2HUacFM1pKCjq/6m
H5yZkq0dkvJthWP5Qnk3YwARnpPIBLaTg9D2Va7KYQNxPIgayAQ3zZH7NvIYqs72
WUCarTCU9cIj2ojJ5iPgZrtXXxbRP7tq+Pfu3C6IrZpUSc+3Z9v8BaW5WHmHrSSL
3fjBIrDzuseDdhGwRaBydVKZJ/n2cWFmCfbHuCumjtpE2zpSc2feyUlTgWrntSKp
qLIbQX+C9fr1z7E2GeeByu1frjPccNRo0wl9WKL4SQEe1mPB/L0grHRVDdT4xVkq
wdsSrtYlKvy0Qv+oHbNRFj1WBi0bV6yO3Ot/giq+MKXMKDMO+lJeCtrPIXCLlFXI
hhNLBJ7Ap7FVNkZ4r2FIzsXVV01nfb8BRs4rS6I2OQNrHGW5VQgYPL2Z5tWBfeZp
MQZlbz9ZagRjwjsGmypTxc2dgBrCTdZvYRQRt4ji7K436m5NskB+vpdDW2hMnNZz
Sre4crZ8kelovH5bOpT4/PaHeIvP1DT6MbeqSYfDx/dCJPFm/jj2dORrD9LCmXMi
hzbOh+xT9Tg4VtOQTWEmm2aCYUwxzRQxgRqc7VuAx58KF0zBabrSEMpfUVIbOxgU
AnChMqzQVCeoQ2zkmBxheby5RIkzqVRek5UnXgqUI9DFCovjTG7g3G896+4jCKlv
ZXaxOvsyKCJ8nalkkn6qKXLAIve67ltGiXQaiDWZNl7rcJJSw1zMH7kJCY/KIDhF
KFuxZnRq+2fUHlO5iFTxuMLXA8UbNcBecAsJc9aRh6stLDUNZc7bO5oeYpAh6tzl
YXd4hT3/wMI1x2/y9yoR0dlIaafnPq9GG0xbILBUlG13DwB5lgZ+sqvlJSpQMI5/
KXe3lKFJD+dYBpxxFIb/jPuhG/6E6yrb85c3AYFru/F00ViSwAixaYURwlf2HV9d
Rrk32FlhtoGMqlj0smqBN9MVHqpY7/FnyWdZAnQS+XQWNjvGLUW8tGY9v0r4iu5q
xiRmz5tOho+9HFSzzGQdkWkcybrrW3IWuOpL3K1b2+qKv4PlnKO+63YcXNYg/M3N
YQDSNfXXxbsN9ig7uR/cwyNPxO/fj3QeQusOsq4KE50ZtSpqDpPyRxOdTIEn3l3r
sJM34s9GGlVcttVRet1hxe/wjz+BKrwf2txk7qbxrPUZG2mFMdZBh1vgqk//aQOd
A3Q7BCg9ykFyy9wV2Qi8MSikSa+kBCRT+64rUpiOZCXxOBIm09ujSjKesMPqaJgy
WiHtQeyKdccn2OxAv//Yh9iL8onna5s3x2L+tITm386GkSwm7fEZL//o7ZeimyTX
CRFIUK1ccYAYCaoPaXbjIiupjpXie6jhUbzpSTqUtBGmzL5w1temHYpQQ9ouaScJ
7mMrX0i9sw0QPCodTotARQ==
`protect END_PROTECTED
