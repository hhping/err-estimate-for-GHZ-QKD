`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ZCJHz+c4txyPAldUQ+DcFgFa9HRAHpDiuGIA449Blj20KT3yLFfChS2tW1H7IX/
OytoigOSPwEglfwu+HfxhceKVGAH3BRVXPekIpS2POmAfktUXMRkId9FUFxqkgdo
y3eagAgFrUeEuyAve+9H8vxbp1rV/uQmJTIVjLFpp5a/JAD7Zy7vR8tHorckLRGM
V+Gs/vtR47BHok8X1p8PnoeKpgr78U1NuNZjfIbXEnrG4MetKoFg2m+dVtmZPkYi
/7JLnTFv2FwLk2AJMfjN6aLuYaWH98IJtdHTouSzkOn+OvYmHAN9klOGBc/AFoek
DY+otepI5ZIZTZ9TXmQeer8axjt/ViyhpsEu12c9L+rwJUK813h18ar+yoeIr3DX
73Uhh+0IOCwg3W15TbZl4QR/4xtS84DSUdulRR80w66/wW4AnwH7FPqiJhahH8a+
cwzIDeqK4qxZEOb1Vag+AOIhXXMAaGr5NC/UbNnyB1lSujdU8czc4vPQ7frNdU8J
DfhR+0qyTpoCv1wHE1QQcyceB4r5nAU2MoyDAz4ZeZqY0rgyATGTBUZt/7IY0aN7
VKpANveWzrpRwNnGXgcGKXdbLpNth+WgKV8Alo4qszBAFO46qqFkSJdNkTUl6anV
DLrHDitVzqu0tK4eCUHrFdHSRrTVF20t/gae6NsUpT1BNveSUEjFyHtA8pRw+Eaw
RzEROmfbD5Td0vaBusT5bZR9BXaBqn+2SJMQYbwKFIPq4RJ0vCw38Aw+Jdo2SBGm
Kq0nommIREybCt8gGC2DqXiSp3ksYHwQbG5pZYXb/We5z9CRWuhTM0hqCIKhMDZA
Om01hTHAiU8lgFODecY6jlZinSv6cwgSTQhsIBkvGGYpFzdBbz50+4uTZ4COpKOM
cNSOyNxMsWbV/7aMtRrWiAOX26NQ94A095fmgDWSxpHWwEzeBK1aJFSuj3EvK1X+
e5og9khRXf1nRQ0F49CCVcmfRu5qf44cuki6KshQOXsq29ANCIi4rg+6eRqF4rJl
TSazVJRicXInyu+XRLVl3adKR4EkQA+ZV5hbJ+OUhWM9OYNVYBPVCrgpilNlvyom
9fLNHO8MKMHYA4m8Zj8Ds6KSAiInGZV5eROPc2omP3Yltdbw7z9c68GE+Y5RrQkO
UZ8YRlaeKaceg/pKdQLta1gpJ2yffqQgppwLwC/HUjjlgi49PM32XCx3STFdKrGB
lTC1uM1/804svW/zbIUi62vodACXkKMfpPIUj8wemJUwEWQAIxmzyf1MWGBD2/g1
dyA3HgKgf/WalucL5IM2W8V0aRxhvupCCLA4BpR5BUUBMP+AvDBBg8sqq237jPhB
Ne9A/DioXAB5+UzdifrVSjMTp994NNU2qKWWW2Y2I/iMN9pm/d2WJsuK6lc/IPRv
GDB9nuQNjJHti6FQFn2ePKbKQTm0NLza4POGQoVaPSCjqmnQRl/1LyO/ai/bh0qe
WJ+Y3QY0C97gW1Ymd/0ANta52RmiK3Jx6/BkRZ0vwast6IRVR+Vd2/oWO16qWDij
DF60Z7P6bdrwemLBsxgnJmtjDDW2fACXriIN+Et85zFDc1lkGzcWxIKAgLbOfixX
t1CaJnc3IGF4hVww4LhWS9UdPNW68/ZP0fgf2l8ewfZzHqwvD/QudOrMGVw+pKiX
GiZoBmNM32vWm59SfkzM1NceI+tfWm/osdic1JCB4RKYDGXzcc7MVK3B5MXK95QN
LGk0hcol+ipcprCpjx3E4uvD+zCwd3MZfoTwZag5L9n9J224sH2tXMyfwV4lVpOy
Bpo+izS3Dk7mq4plDvriRw7/dSK8jFUoKACoXA/RZk4HoiJ4EAYqS4lFEd1BRZgG
MJ01DwVnXwiXr8whDlNbGtvHiMIEfjjPPtGXdM5WbK3p/8l+CokRdB6djwlCC2aV
kpc/FecDuiHo1L6rdXCjFA==
`protect END_PROTECTED
