`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33mhUD2a1befpiapyU7zZNHOb2xkp1bROo0/hsm0DDIcwnWUkUjkRlT83MQ6AAjm
CL8oR/YUtkNFudc9hehcm8ZdxHM29M6pFOi1cyR4dqClFyhSbpgWule+b7R3Hn4C
we0g63G8U7eOxjMWk4NjzY5CF9JczEq31jfvIIx8n3ehAPNMqfXB6oO3J1t1hs5B
dw925J4HXKWIxEZNengOTSLuA4vvCLfaSHpkIrkgwae35Rjp+zrEdF6EkQXquOih
DGCMYoxWxzMJrNcWYIE/VV738WGxfOvqFYadqwdCiGKkbf2maJznsDRsLBsLfeUT
FfKB4tGY0jwffR9g3KQTHnEB+VM/cV/DA6tkAcymwjLa/vu4ngdVyf6tZSvwpSDV
QlW8NxWNYFTJcnH70PBF1nUvnsdTEEKQJ7CsofS6OrqecFxcafcgZeQWAPBl1y02
DiNcOgL8BJpd2oM5pIqYiplwVGQjHPwg+Uo5qMMU6sFd9Qx71ueVvqqAG+NlSEox
dQTI3SYTntIKnnhXEGMJdHbkpzDCVE5IqaTfXxvAVdgqubrTQF0mxcrx8rAMuRHC
TPwQBM5fyplTt1KmkELbACOiH6WQ44u+Qi1GgtGvSappwCdkuZeTFk3QXWVon8/g
UCF7kEySVKKogTLdqG/RpeS52b6EPHKFbB8J0+b8vSe3wB9Qh9galXmyOShAxmL5
VNpnBpIQmKb+RKMFP04QeCtcbmupSZJDa4HOjxI76fLDBo5BfmpszJBbH7t3YTP9
TiVPiNcD74jFYDZ8yMJXflf6AdFkJkF1EAJcm9kRRd3ST405+RH9DC3X9d7xLW9+
kXIw/Lihf0DZGB5XkFD17WhJdGacMiqhj4oSJSHXAUaLH92H8H2xph9iX2KZmAV+
`protect END_PROTECTED
