`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sQKGAMpgUK8/JN+o0TfuKJcfpWvw17XccnqPEzcv6MSz5QB+6+RAcXdl3mqe+zW
95xC+TV6PSr2lAjNaey7MKhgn2jAIZryjfoKbqlDRR0vpY33o9bt4RnRERvVgtv9
DiAUorL4WSNEwVraGjxhNzk9HiVtNn6nIZltcU4BAkb7QatcZ55N+hiIWuzL/AIV
qBT/OCvdj39cpRcxp+mPgHuQp1KAe7lWOoCbBq7Da2VVJDW8w8cWnlEWUsY8yMro
oVzq+rGAqPuTVCXZP9aL13/w77C7NsJr80HtVOnLmfuY4D/EQPmA5i79Glb0ENLs
j0qs1YuIQoHUjLhwPpKp094U1PANO/xjAuGMuTdIHj4R4HBTlrn3gC4Frsy6L6Xg
LDkZOfZyYMbl7985/XwmD+z2/9hqBVgjVqsSJ3TanmCrJOdw2yUsS8u4jMKtXEmW
aCqwVKriKoKIrVl45ZQdR+vmGdsF3+a4oVn9MGzFzsFiFj36LzrSG6MCY1UQP3qR
U2yj9elBz7rJCF4+X7bFKuNEpKCljywM1GwzXNiq0+FNi5nNXzR6VvDIiS5uw+SX
kiHJgpI9R//Nm26HnvTMw/Zd4ku3yGJeI/waJtreIgGGDf5caGq1JhLFS8AfuAjj
DLaNlaOiyX3JcYq+YqhYLUuxB7vt1OjicO8rSoHIYVTE4uTcae5Izy/gBAevPGZL
m1E5H8LRc5hd4pG02B6GxjF1EnNg+ruQdah/cVT+6tIwAwlkDu/AH86l2vk1+b+g
OnPvVKeyWlRMSIVJMRpapQ1vnkDuxIKNVUeuetZ5eSnIsN/v6XIeGkQYKu/rZU82
1cCfD3qJFIBoXQrSQOzOz8N/yLvBQU7ahFRlYJp8HN+zLL1sdmOQOItR2y9efgeT
RRgwx2dqkOiCiIw83y9DOe7UI+pgWm+rEV0YkCTftxoSUnhWRhSPfwa4WeQvyqZv
Tqz81IBT/1ChHVO1OEaWTWWb4riYPPReExFrKHAVYSBc6CoV3jADqjgw9tkHVs9D
xJDB3zNAgNULl5lTu8FoVTfNhmcmSiXuzXD49/XqcI2eEoYMNo7PaO3e6XkMNGOC
V6GVxvZnuayA+2bCu3rE/jn8tV1vOSHcglIbZFHQR1sckP/5eX+xyGpc9hxFpDFr
DvzUvNWKR2EYN1vnsdy+TCSRcQymE5sl3koj83Y3ZE24u9IyCZo+my1/KspTtz7K
HLn28WG8zTkxGkPEmCSaButu5RTXx/jYTKF/zzRF32g1nb0BtldPpAH5wopPRKS1
XvngVZ9PpOfQB/GkPLz/grsp7e9miurdNP02ljEsm6iOgsNZcg4r5iyO9MuKwAnH
ohFTPxSmqLWGYlGthg/PCQSvkZGaE5veS5Qa+GDsKC94n1QGGymdNmsH9fVfoPmt
e7nXVINbhZ/7lZrYN48ZG1HikN2HKXuL++6p6qhyYktdz27boXYoYDoPuCa3tjGJ
pbKnNHWAH4SDc/z45SS9uqKR6907eWP15RIxY2iCVy4mtAOLw+h6ArS2Om9DMtGC
SoZZns9BFjQIs9q7zeXcUwimOYVYnq8YwgDCF1O4Li1f7rTQWqEK4ZK60tl7DnDi
WWSR7bagtJpqby5GbeqwwMQE0vAOUz6iMWIn7zX3MmhiSTtyeWQxZtJyM+CmfIlw
hMwg66iGxfTfnO2soMen5OG0Ago0BnbPtEKAHHdTBkv4TniAskeJcxBcRE/wSqlJ
uiuzBQuhzJTAR9oF8x0Eu0GyMrKrItLPq80CEbPwEnqyq4ivsHl5IqRjKbkUS1Rr
v+NQYBpEv4cAt4ch7//BwM3Xj5XWi7JyyXFu7mNPDsLYLqYbmPc/BVOv7u7bcTIq
wyTzgss9VM4Q+TCi7iEqo/pwm7lZbRatnwuVtw5OC0m4K/PuUzPtfYFcCLfJgR0t
f9dVRZT7N1omoEuoSJ8rAB6kVVNUpKJWyE0LTiN/5+DNTEQgmMLpD7YYrbgh08bI
xEJkJMUV2zVRWSX6NL2PTuCGhURRC9+Jz1qkS4TaThe9qpzj8tEfKiK8SVegNbBz
zZP3qMByedNJCtVoMLnvmJ09ymnpiye8PDddFJt+nMFwx7OI9nOmi3OVyUUJjqAn
e0UfcW99g0Zzwfj/xeVoewd8mHIGm0dXOtUjvLeEa98IZSPl7RkbC5gxn4zOGv9c
dg78gg2TklLBp0wCdS2Diy6hvthHr6GiKxG94NJxz03qEAE4jo4aapFTCSDo9lqc
KszUyXFLbBq4czYjVFcYH3a3SC1VCgzkZLQBCf8o1dx5IVvxzmhrf9qofIW0ywP8
dqGhyI9iORoJDx35K5aXG5+PRRfPJpl7+NWh8DaQZ+mXTFbqdBxJtn06VNQ2Anis
+qamBRo9I0yv0PUh/RWFCxaCU2ynELXt9F8hNrv7XD0wzLJ+qg6dL2iAjw51E1c5
VoqGIXaSuk5eVCKnFDlD4RhUrZ8So/HZuUAd5eRrF6ABZmj5CDU72zyuwZtYY9Hn
t0akcEkyBiBbmGxHk4Yy3w42LGkC3I6KC4c8wuWujT7Tp3+9nNPMbHm1H3DeOZts
yYgz/VJBj2UGVI2sQPhioy2kaCfUHrLNq6NFsOxKvOgVCeVzsykn8GkSZcNCeKAP
KMhDYyQ3zTAkFitBcNfoos1iaAgLRn3qXndRvw+vLV2QMtvr5DAhfuwUJsQ8l7MD
VYkTJNFIrFlhNtUCyHm2QfEmI3pY8seT26ET+m05T/X1waK1XZ0tw5IkKrIhZ3bv
W1MZCtvvPSLMlkb90AmZJGufJgYegqvB/7hMOkXxcRITUeQB6cEo+7itV9CfWx9N
yyW94OsieghEZqHAhZ9At+1nD5GWdK7uGx15dwaKRoALQR51e90IkhDFaVhXTJcu
OPV15VGhKZSeq/BYobKdAijvK5Hk5ntXI3Rk4kVDKodTzvb3RgrH7NGOwcxYh1iq
/Sy5FgcX4T+ayO+HaHTafvg5jMUrprKrogtD9dKey6bVICACCkVZJaWyP0gGdk98
G/+c8piakUwaaT020c9jwOKuGh5Z7SzrQyV9oHxGLyGmsdFUBKl8lYIDlAYTTtaJ
Vwi7yshZAZjme9MevexCWPjmt+Cc+J2bv4EQg/h62hravwKXCkFYp69xoqpcT+6f
ePfl1zYRYCOz+30vuNuNMNKo5SQlWtoimgKAJLMyOm8=
`protect END_PROTECTED
