`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNiZaNzkFO+WMXKO2xeSRrSqbwSdhWK+4uTg2AWb1a888vCMhFZ7Jkve2hFyc1X9
+U5z+E2ISudhE3D/Ohvm0mnoYeuJ2PZg6GP75X6F6LcgDSl+TLqE+/CsSaoLuuUm
YSrhUsjzBE9rKowIQ4nTuLycFRVVYdkVZFyVbdjd/v2hypenqATebY2zcY0c8Bsz
n/XAJcnTZ0INmfD0yfoyLOrtIIJte8pflZ7CqCuOCsRGaqov05lseCbTnVtRlA3X
OFnH+m7zBTb+w4am8QtGSUi4ksAX0fHzLT4OD2ZWfyUhlob3HT9cWaS+7t0KjKRL
peZD890n5CKBrVFMP4UTIXfs35YlQIzt2izLyp63VzIVbhs1nH6X3V/+X5SsAGG5
fOY82q6nqKDwDmW81SikKH8vSZClNyb9OYhMZmFjgy7r4t0oSyvgumA+cLOzqVq6
7RN78K1cppXgzvo0cvpbJ6OL09fD0LacUsRbr4DKJ7UqY7fVNvqH/1aoZsg0hvj1
BSkIdCD/GBBL9SYmsy/+KcriwBJzEF8bXr+zOS+oVMxhyXtYJBjlfXTOsbEqxUoS
KAg80tJcZYvUqXjNi+W+Kp7jffKd/lGF+os9uY7mPeq98U+EFdKeitPohZQssotG
BNoCcw+eh+efgGMxDcqygTpoGvJalUkGmejf3uOEx2Sl3c44VfAM9shwpXuE7NTt
EiB66mRQCtgazVr1vtECGF2gIv15PXIsMfjg+IipJnBOcOJoSEU9N/wq/62z1vo1
BZN5QQXXNqN4wAxvKIRmW1G8yF6B/jq37K2lLer2usEkJtpBtdq9cNQo6FHHWdQB
6GCpQy9I8C5l8L1/hb/+AX069QPRt1PXkiKuBVyNhMY9r+83z9M/FnExWBPmq3nu
WKsNNoouufVSwmhyBnlQz1JkEduecbXRSblKTMc1/vOohbJYgj1cpvjwenqNaL3z
Dky68VABxtmnXZAZVdL+H6vVrYc3H+W0k6TxY2W2RUYeCfX9lmwshhebJn03/8E7
/KHJLkzEydyEk31SFDLk8efv/+1AfxWvzKjUekBaR8d2jEIimrrxFfoX3iHgvxRk
pQZDD11UP1lheRH+Ml2gD9WGdUtLXvbtxjyxuEbNly9M5uj5FiQYmeLvTrJ8zd8v
UVsmq71IVvQDGtb8NKthixwsXrWRIiHiSOQfyBH4cSIMZMf3DbxBGUB5d0FZUqF4
yEsVyc2wQnlKo8zAg66wNxyd8VU6Z7vlgmZNyBwl8NJpT6Ie2mbLLG7Wrx+FZDuo
FJlNo82BHL5lfHYXMvBPOMnqcmPHFOz7KY1C6RN6DV7NozhaVy9CkfbwvGZ/Mbc6
3id3sMxwcsb38JZUjmx4exK2TNxVVHbnXsIa2OhpAQD5ygpy1M707y7g0E9g2dgN
aFleVHks1sxKz/vEjdqA4aJrVTlBxI3xfV8Bb5wfFTarkG8/VaIAUvKa5IopVnXj
1K/K0++jdVd5ykp2QIlJgg1baxCfpQs/mtn1r7YCEKuYAuMBb3R6//IvC3WVQofX
2PEqipZNzxzhfcc8quHco1qrCFiE4Uvpj5C3inZ6ZJbWlYhDkM/ByS1EN6Zy1HSp
2cmlzAz2XpIh3HL9gZXoUuTKB10r7N5EYNtGatxf0MGcTjFGo2VxxWsS+RWt5pUd
vNuNXLKpUCtcF+ORByGTvnKuuJ0GVqzx6pVPXaqueBe4lBRXZZPrhgoDUXHNzwWi
hCnjQFckuov+WDuQL87B6KU1LFUdXirpx7JzBAFOmsxENJxMx1kNz2VtSygh+MUX
uPs6sr0ll18PkUewkgcR1SkdWfnIWsSoGunX5r8JfYWIPWAfazdYP2k3eVdDy1Ip
w2HIiVE9nF4mhZd2l6T0MHWj/7AbHAB2llsNNVOfitnP2eGaRI4+wb0ptGHomxH9
6hyJihrKkyxVAfcPbZBKg0Ki57IfS3K4Ul5bXjBXp66qV3ey2IXe83zadYjlTPJL
2buYOZ/WZSof1TNV4KR6Obub4F1dUJLf41LxSK3bt6g7XtNI4KUqEbBftLpeYje/
4++O8ORgkWIxDOWCkzWnaYToWOwI20Hant7ONWEmpGYqwBKrTIoxVAgEINXEWRYm
dmGk2DmNt8WqrR45llrdjjh9DX0XI42PyH/crQLLp3O/bWeLpZ/7AysxKS4MX5hQ
XdqjWR+qSYgT8MBQDRzTI3IgiqiD3qyLWNVW+as4YUe7rqNbj/mk/66II7LXbrlY
bSzi2bFITdO3J2SVxhR0pEM/qLq4Dom/usfSziRcV5/a3bvqCQWsahrHdPy3ZOSI
dotYZ8ltaOHfD7c563x+MYXHUecrPt6FuIaTMiz3zptVapRJ9YWZrJgrc81YRFJR
hwJc+TdVbI2xBjM1w7sfYXO2ttnmZyrAAOcuIMtSERSYlsH0jA+RVtetFKLaT2zk
ZwIQQoxDo5At9+uRqm7ONsekSYp4FjOFgAhyzLHzkrdWorom1MFYby/cG1zWSnkM
DvrHNe69ogl4wb6pWAZmonl8g8n6lgvz7wVrrsPocQEiGvuBydpOemD21s1Y9Ptw
gKUCNMFzCKyMEaNg7+wPHePQqzJlqYX3rWiHBETsA+pnk018qfGMDynQXQZM/WHj
EAUuA1+BMksftxiAUS3bIdd5sLTb1/+lVRvHEbWJ020=
`protect END_PROTECTED
