`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OByWZrxqdE2KRdX7MFTuDPKKDFLDisPr1ZWiNd8Ttu9hdSkeKlQ8TyeYu895k7cg
TmiDtXkHAGQGAFcX+rt1p1yTLkO3vs6emajQZ+h6tF4rGUHE5aOfPbUiVrzp4Jzk
tkLWLZ2XJceH1RPG4vXQJEEQYx8jW+30Rzv+12MVJD5lY/PU3muaec7Qkum4FM/b
Jap4Gk4Nr6DDXbduXRX+y5mBEFQhjAnZwrbrAFd8xapQKpmDNW4RlF0RIjkbii/q
TupWaC1D/04q+zfpsr9oUElIUAcrP0cg4m0nT9UYwYcEASPF/bIlrXb2PbFbCaLV
H4vdzLf1k9RqElOXsNxzSUCLOFh3SVwD5d3jOh+EhrUPsYecGpvD1UUJieiRiPA2
+GJ1IkdI+erO8wDARgGpanVs6AvujDAYPmijwXOUBaVmHIfgCT9E/LzlkIL4fUI7
YYbcJNRykf1GRy1b+4ecZvXmBhgjIZgEDYvcbuqO6DOETZv6B0arAMc9XyAc7Nfy
Gvt4YHA+gbAA51Ojaka3jmtZtsRMLLZMCPSZWJ3qmH6pUcSA5Wy8twrZNWXD88ZJ
8KIAV7AaLBA4SvfyPuN66lnvnKCLgEEYm2FqLuOF7cY+Vr7drN0N2pnHvOv4ty04
5ZUUwxVY1FabBdxt2UiRyNvVUaBoCtUd9XLakrGXwDI2g18BmA+HHF/Mm4mZUkaj
DnRB9FCH7c+LfRjqvRbVHJp44ToZd3fXf7BeSifu3zVWSJZv44nctPfHJiX4+tP5
v3fYJDZQuURF7Lgf4wXsOaSUla8A21BoJlpxO0InacYrtswFz+yUgecD5/HS1zdl
Tq8JXW3dp+nFsqZLHfv6eROfWWiKlQ89Vf3cQ7kT2608LP602G/k3DeMPa564ojp
H5hkDq7sRXAkk5fjPJawACMZ1UPExcMBuXgGv87Fl2UyGDZAdrwB1iYwtBNd6N3u
Ak/tKDJuDrBODIx3mOkyo8JiP4G/oZeBJDO8U5mP6zsw0XbckDctOYZWWsYVbsUY
hk5EIEtGw8ubZAeAO6uyAg==
`protect END_PROTECTED
