`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sz0YXuvYnHi83iEjwGTaoRP2h8p7amHp/s6RTTiyWLgIUcqxjHGEpzT3UHELR7Gu
5OYL0LJMNklL6sSIskv/AV7QIzKujY247rEKJaeDN6UBpO91sbDjIx5h+6RT9wwG
FP4N3wzigQXVX+lBDgubnkWpD2ufFQ38KzxE64how1Q3amFuNiMzfKuZN2/5Y86T
IdlcLU4GvweRSoD0su5OuqUvgHmigV4ojNmXdxzuXvvsrsqv8U2Z0Ur/BECAa9vT
KetoQ21GlRzUAbjWPhnqSTB0lMYvg2WqEB41DjEY+PLfshdNXS9pcPt/DA5n1hMe
VnjKV3vdDgJBBE176ehrCJs3IVb1cjfwIWh5YeAVQ4qpt8zSIWHetc+seVQ8q/lY
/tZpqt50Dbx0nzQM+tdPtEfOaEixKlClOmHenSi8EEGMO91LBdNuT23bGP+2wrjl
LU8USNByJ4ahP5/t+mNkNHetDBANTqXDsQMDzy+dgn1+L/a9pbaKbrgh0sPPzaqc
xg5LHmp9Kna0H7sWMiRiTMR/qE1mZg+KpDZ1nWjWNbyZKYApRvCMZCExp8WVj6/E
XgBgizsROanCRpkpvglKJmiiHa4W4cqmv1hhXzjXDUyjzsOvMhSAOh8l4HzWgmMJ
5fP/ym8JVWCIohuM5GMy8M8gbtR+xFwwT3sDeHyLcGn5+Q46TymgyDx6ST4caObS
Z52SSIWyosyeBMI46hEwTP9ugc8aarkM0JobEsjusGJL/Xp/yse+ZFiF0f6Bp7rB
Mo6UXpWppHrQb5FSgMdbI0otlUOlZVHN0yJj1H8qflfCLKi0T8CxKTKK+CJHwa9G
tAEGK1vRI+szoDy2RQwwAZuMrApXuyY4ISnBVYkfxMCg6BE5jR2sLL+r6IhgUHzk
mHMW92J4+Ak78dzKni7E83bHEH5IYFMPw68ARiB0qIZIBmzf6dlltlarQWNRqJWp
XN/i+2mSSvozYb/FD0Lj0M25yegzlj6GHTtuRhNSN91HsRBGIGr5MJhlm3f1v4no
CLrU4AAtDscbayjCoCJpjHqxubKYcfkgo2w5L/67EXA+hmWN62vlFLqTpfEu4UIR
lsp+wwDW2ABgav2pgn5C9c0SET9ThMtCrokzfOA9YUgwM1d368soUZciYWAjTBwC
LBoRkxWGDcoJlaBaiALOmh/fef5gMmDw5Gnqoo8AHU0=
`protect END_PROTECTED
