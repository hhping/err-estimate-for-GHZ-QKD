`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8LDR5NxUTd9UkxZ1X3gkRMG5lgtYEIsgIusssL8WUq9ciyLqvhP2Ur+cp374BdS
tHMyxQiKIu13Nja0n4ZDsbZGY4zvMyQT7yMhlUtUSmn+msvGtuXfn5kHWaw1KKsC
fyfNwk5QOnFCwqnNvFUaX0EiNJ+rmm2ep+qrMlb09WFvWpbKn718ywM9NnRnWfGf
InU0cTVNZFjJ60bAk70eKbh83pRB/kLWauwQRTgIya8Mqqj+NSyNW0V3lWIKXxDG
R/2c6VGlKlrU0+B3I8fuaW5YvrnDSyeT1XzeJ1K6f/+owbncjWHcFamPqrtBENKC
Icfdce71hm6/+/+YNRLK8G0MtQTc4DJY8b7UdpTosSZWCge3I+4i/DOMCTx3QgkS
lHxEACFTCRCHBXo9e7ac0cWV7fQ+hQ1sobsHac0mVqFjiqWrHg0D4x27RZ0IfNlt
IvwuI82r9s80va5QAWmb9w==
`protect END_PROTECTED
