`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4j+Q0Xx5RKgEGAIvULAINT1Yw+7/KpcvhLrA0cQBZQHUfXDbifb3XzTe2Ow9ELl4
qlazNxHXTXGe/mMGcXwvpa7+JP/yuvnKgXdZip4uP5806Th+YzknNfZRteL6rf6H
Y7JiHwyxGoxhmT4c9acM/sXj4MmbPaL4ewP6wa+rFLJekTKGeFDskKsumLtlYuZZ
hEZDIlE65ZRfAmD/KrTR+zsivbnOUI8g+NGLY7kpeDWvNTHNRRKUdiqilf8jDqO5
2mCvc5zc/LffKDL0Ng8p39HNY6lxIuy6/sDlvIXyIDtNmCVgehOfmJ2znQAl5oBu
vP/+lKNVuV0Zh9glBt+4jh7xnReAkCFlFLZYEJ6t1z2qyhX3JvniI7sfmYqZAfrR
b/kNlpt6PDJ4tLsJpwHJtQfukmPKhYKQAXYfY15taVGJVMdwTDwULA7IbiJcC/GS
oqDkBzeiRYOSndxK5r/dquAvu3AQbGhQwk7wMlat0V8c/52E2IFUXnAG/wbM1ouA
4OP4WZ250ECbpLoSFkaS27Ch/CV5/sb5kNqP3/Uoz7+6cf12faHO8Kexj8iB5mYz
gMt4967ZkB/5iJ0p32WHf2yI88Pf0+5ACD9RUGozx2Q7WA0IrCXoSIe1wGIopkin
w3SC2BXwEz7htfRtA7HL0sbRRi0Wm4/lhTZy+W+Cohph+HWnXx7w/kkhf/9hTh/8
TrsBiWlGLtdnUt7QKGyWKkdhfZMOuVL2VAYS7KAIpzYb+s7WOzhKfPrnr8PcDkqc
fSC1dSyULaR+dEyjIsZkSS8ejsLAEfX8a/tDpZ5QSTlptyLBDSHoTWGL0MkyL5FQ
TrVOzgbRBrULahEnbdY0ldLJL+k4KE26VZXn8/gRiXQXOvIuwuSmQZSApPbgUnN/
KJvxAqjFbe6877SKi4vBVl6Fnr6/MGz8sXKRuwveMWDpO34kOCTKSigHspa//RZj
tdAdTsMRyYKkBcTlqghBcyh3Hy39VtRAmTHJsltl09OTGo529ViQUjDItWYH4oc+
A+E0hK9AMFPGy7AwYySME6efCCfcU2PH8Q8uT9Hs9WOEWDIhPssuBnFqBtu9VPPY
TLWYKLcBFpQHvh7saakBb0oCst3ncaIb7AfjQnspRXVw2l6BsmdhBjcjzsGkEovq
2e5BuSxY9pfWrshsqRPLR+jiQM8c1C1hk778Ax8WIL5tAaQyFoemXZCHySlq+lpJ
wHfRxnN/TNXEBRf//wSpnQ==
`protect END_PROTECTED
