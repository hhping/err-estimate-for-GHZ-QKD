`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyBZvcf7AITuYxyypLplEwr9Ez+Wx47lxDPC2liJhLwAYORY0SQKKozZEyBMShOa
dR0WULkIODTksWQExbaTpx6lO61pz8gVuCaEyDVV6vwF4azJFfOKzrzxDKXDJdX4
l2NxxlHt3KCwXjZjKLPXOiAHNxOSMUBIjxTwGe4z7hcC8R+sCoP7YVqBlXjc2lrm
B0MJrKlYviu8v2pbgEGOl2b5HBW7kXuxYyrTuaWEsjib06FZPQXDwy01OPiSzSxQ
a/3TB4GISw4Fl6obAHzRhUnVX12A2xyoyQcZN4c9X40Fy9zSO1u3qnywxTqBH7L/
ZGyu0BpgCfq8NC/2SMJtwY8R3BXKsxlXfROO80WyUBEgBLFqMCC0GaIVV93S6lMI
5Dc5wZehF185lLC7dQN8mFFIGXGCoEKpBzAIWM0bi3biAY+wM6ez6BN9DS0jN6Gu
tGxF8+/e011LMy8B9qbwyIi5jrBRsprGOVnUbYTVW0VQFZ4o+44tMyyYhsBfjy0o
ZkHd4w6waqFK5UJvAJOKwUvAG7nLp8P2Jmorrs3h87s8rLHVXzQXGwMXmfuWirR3
djyzLjy4HWCXloRA/JNb9SLHUOES+NysGhcYnwqKrZNUL4FAucYfTIHG8NSfF7jL
xZIsqPyaehUqWKoO32VlGnEIcrN7mxyZ2AtWTCRFxykz2HqINk9ZsmjdniIrxnTj
mILk6Jienw2rCAOAy7yqgDMpDUF1gho7tEvYSOIWs8c5L5+bT0TppxNLH2fKxVoO
0jedVFWDby0FZiuwDRlHtsEaa5LjnVtdP305gRW0EfVEdnCZe50RXdOI4uOBAmfD
ytMwpQ42uShDfNzSe+WG6gVBsHMM76dwsSn/mdriYMfxRURqEcO/r9RXy+20+Ku7
IcjHtYxbE5FE+qKJvBtKCpoKVqTLhnQfPrRsvYdGvsGQZPvJQmW/hFRKX3Hba6j8
47lvabQ+QT1CU0Lj6oAMps3jOuiyfGJ8Dg66XoRiaAYMMAYZ4W4aP78lXF23HDdK
sLPoQBH3hRHjrlpkhxiY59lDy0shw3a8JoW1m6D7Mls1l8TUw2I4YLofMa3XQcIN
9K0eLh2C75gI0A0JAbtMNc6kW+NkmeAZk1XNFwaaLH2SXjm6aCpn2djnAFrgseHJ
awTbAk8ogCNNyyPv8LJimyOulE63FXKlBu3YzIDEVXJKBJGbBi38hgbotU0EN0VT
zYKoufu5V9QUhZcTwBM2JC2dZkf8cR4E9Eu1zJQpcV4+euSyRLHHTeaXE7V5bD8n
XG9bFxg6v5zP5XBcbeCrjFRLRwczsUe9WVd04wk0rNFh912WJQjeMPQmiWiQs79C
P0WzEPt+PLaianQTs8s/Js4eEZyrLbVxJE1i6z1XxX7aaWTmGKr/LC5XTLDQpcpZ
bhdFDExpCuF0S3/30A/bNymcjxVcGYc0du8wgXBst0qNFmfm/kYpI8Nl9IeyM2qT
E+Dyo5ajTXKpkzA98eAetRX+O7m1dqhGh1iGZlMMmM28GW1vFXqcGrl9mbHheKzr
gDQb8cXs3JRZI3bWRCN4enfy2eFGuQJ5LBZhMmAaEhM10RQHxgWhiz3ZFKnpKxqh
d43WwGNKq9KwLb6zLw7B6dSNpkxi/14LSYYKVH2/2qApu+W9V6chJdY5MQLvpn16
i3KnzAZnaQO1PvTAA07KvGN+0/X4ynqx9rzZsqDlzxssL4eJR/3RAQ0Eby0t5cdj
O/yF2g6ArN2qzsxFCPzb3oJbFZmioDbmQ+vHX9J0XZe0pH+V4XG/RRqnoOHZMX/u
Cj0G/DMeIRyrDBYLYn3xKgXzOIqF+agE2SFgUG8D2gaRZFRyqlNMP4DcwK9DGTOX
9qGgtVd54uJU3McLJTQtZFnRBqJNhTMlySVCUgSp9jcUi5GIOZ8oNHknEL/F5WCn
v8a1N6kFDG1kk6EpCae1tAkxGFWygSCaIaC1khDtIIg=
`protect END_PROTECTED
