`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7oqQdcwUuK1jk5mMQ9YrS/H2R4ECcI7rh1VNgEZ9Bq9AzMLvVuujvnadqmSGYoI
WUJMToFCVja20pD+QBZqmSWmDNaBAjbR1KRLd8/4Gpql7p4FdBvEa8zBa75EO1Bg
MDoOW7s581IX+BY01lEBrX4itR5Cpq2gJJh5gBFlDAKQknL0nIjMHjjxgJqha+g3
Bb8yatCVzQfc5UXflkbgbCcREmIHo6OpqLQKzqfngqDaZTdgESyOniAvp4ieeV+a
L+AzK6+cuckTjMxpm0JQ52+sNU0Ibb760w9eNnKkoHdw0iXyAudDZmBnvJc6YMMS
DUv87gzVPOWoqldWX/RRgmAfnlMsU3xBIhJrjHihOQvGtdgoFzM+c1SunAfMZAUv
hD9eoY9SJOAXFp8rDtL6HHpLjmd/OCQjTVGTtZANNrKj8pvL2SgKOQ8SJLcY0LTs
O8iUGLp8BWxid+ud4kIQ/DrT95L+N5KWQuThqPDyy99KyaEEzh2B7S4nhYJwq41R
pJ9+xnCvFteb/kECj9Kd4nAaiGGanibVTJgU9DCuz4/rhaVDCzAIo+75x1Rpt6kB
0tKUeTDfJ9V17SU2GMQZJLZZL0PPcEJ+6WAgOnpyxsLc/DQVuQ3pTYjjq6GUzZo7
0iU4MuysLvl31Nwwf3nMN8p+LWuT/SsqXTP8sTiYm7/LYhaDpwsF1jSTXT5U7iRc
wDFbeyExNk8dEHpS7flkDoBJjzAIk9BEUk/uCmSLZVWpQwU5XQKlJ0BIbpH/HNZD
q9knrJps2R3O2TTEmtMu3hca8wDhglSZRl1fVanl2sEFbubYFv5uUpFn0owW7vsC
7JglpO2w5s9oilJeUOehBVfDfEJ0Zj2MSy6hboh2G+eTcIubaIMYy7cnDZUpsPLT
2JBbB4q29nWuNdh8+VYYMG9DWOWzZia/Ut8zpKr5AyZ9OWjTu69z6Ezqo74a7oVW
sLsFY+BlaZIV7+j07LTfOTTTXM/dZBu5uw0cFcP+tOjplJEzu4iICMXhu6WmMvE7
ltS127Wfi9YkdPYdfZQbgTt0pa+zRnavfqO/5cDTNHJfNUq+YHfZB2k+tgFrVUuG
gUAadqsN8uZ6cHFbkrKzZw+lq/b1+7tOzWGa3HplUnxk7TUfhF56xj5tMRaDiAE+
K/k31CE0+y1dGOuD37t/YNccuef5rbfsOw9pTSQdbzg2Jgkt5F4dXBRChZKsEBj6
cEWTUUEmpLdfa1LLioZDdduGbN2g3bnpeIHFVOm8HAfNdm4C9dWWyJ3jArJUHR2m
Wj+hUNpho23QTfrtRoy3bD25uw3SYvtQeQq317pmQKZvFb+Sfw//W55d6Bw44JVX
KAIxd2LzL7mlScycImxQnr4zbpeo5RGFwFxBEgicgUZSi1YWocUeUfTu2JVGQt1N
+B6ytzYdHmFktdjCFjMO+x93msXLLkj9aHBuX3YlbA8iAiDkr5+BgzKIWb5Tp8Qn
Aq6qNu1x3dPK6aOmOXweAQA4DvEPfpUCzmtWljjLGRZOO0/LV132JS7ydjEQZgld
OvNPj1M0R7Qy54uBDgZ8XYqamOR1cKV6JUpXaAjRpi/Ae8f6/By3BE3FzOfM7LL9
OXDVtzTcleqZZ0NTBEuTq8NDYX1G1JfP0Isno3Ayjfo8MG7N2f7hYlWQpp8YAZfg
80Q9Tt3bvpfoz0f/ARj0eRCR1g8Jz/SqeEoVjkQt7KhOav4uNp0q1o9mas75IA43
qYCA3bBC8WjX/xcXfFgUKSCFU+Fo1GTK52GUj7U0HY3NE/qXqp3B4oYS8TVUdkTn
wBnGiNUwRJsudu860vdM2HfAHVzgyP9zjgXKE1+U/j1QrYuPvPIHRb454gYTu4T2
im2dowBT3eHtQVJcdXLr5Of/SrKrXDRlj8o3AffD+YrqcDSDMZGVC8iIm41dPHbn
S5wbncE4xE5YAfJCGS7G1g==
`protect END_PROTECTED
