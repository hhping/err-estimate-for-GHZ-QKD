`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LsM9j/SQW2EK4eNn11RPfMAppx/RkjVA3ye7zoMwFpRrrMJzHQJPil3xULHCS2Zu
vQ9Fn5YduoHjIcVfzhd+7n2fc9Q5hb2CnS2uc+9C9eyWGYPN00tHe4F0vF8wClO0
qJU384Kz8zZjqNirSEXeTCfLm0cAjL17Rbzx6WqeD9fbO7OF/BJ1oJFraAjJhf/T
KSZjypZvvRETSaFjymq2pgMZtd3CkGLjvtHfrdJL9xy+Jc1yM5JnSXigq26GQCZO
rA62QnctJar7El3TqMRhVL6rCBK3KPfbcYHrRcIGR9sWhJm12/QpRWdpTwgGYP0W
V72YaMojMFvSFrRKxAiMnklRHeOpcnzdmGwR81nA2NZZrHEzn877f9528zrFIqwh
BKSo5I/ybKUafYC3Soc7vxttNtOGjX9MJFvXzutDZ9bdH9diu6mOEdNiQQ1HdBJn
Gx1v+lEANXgnyAO6ot+fs8Syb8FnJ8PQC5A+DJXeRPGRvc5Aic6Lst8VLbjUfrdv
VacS8uoRoqQs8dz1aGdmJIYJd4Ds2nq49Qb8+h4qeG9fscxx9KKJS+XEvQIHFEbm
mVt5q4Lld74y87ziuKS/EVXq5daYrKuqZ99lNCfYK1baVK+O5IeN55OenwYBIZ0t
Rz2wLEEv48zR3PRIzcag3BBy0u0e+Hst7ec/teKvoIYUsVcsJONgfXg2q+pzHr/Q
IlHEqxFGd1vsYpAhOG53lGVcVhparPPJrilVyAWQWWZztYbtj7N2ihTex3lDsQ5M
xtqj92MIDigIGye+myFb3mQycqtc7f+dFwhv2taZJs5t6lwUEcw/8mEgYUX8BDJS
XcyEPiGa77KMM25LC/VuG2+oN0QL6TEW4IJF9gz97XhvG27xTpLSBeN4dN7JboxK
CEAc9kbPCbgCu/cJL+ngk0JLTfFwud7E2uUu+PAOHoqKlAusB8tCltJnIqHeZ4NU
W9oKW8BdVvwkLU87nuBX7ElnOYbMsaIOKwBNQ5iodLW0dPP8RGLsmKNueygQlYC+
e4DqP088BD6Svk/GrgmNIubqaTZv9nlBx35oPgkQwRCHTkRPnZIYiWeCf5HQeDZS
7GfjlEMa+9LuwuUL0tws2KIpIoDcr7DJi9mc79BbCr4xO2nEJykZ5SxAZnIBujyj
qZ0R3PEfrZ1NshZPLfKTI3KUxfTRreNZfo021YIFsIhJt0nLehxnanxnIYb6Aire
l34Yj0pQ9hP25hCPY1v/d5HYX7UOzLlsADegF1EKuZXGSIU4pMCDzwmxk+FaLKE+
K5k9K2jvPz6TG6Ab8iGTw5TrxGb2eimAuprIx+ggK/md8jGIcBg7SvLZRpR6PiG7
RRSOXiCP1V1IATA9D8cbMEmYpHHeIAV9J/9xOaYTmIiGg6wFSer57mipAnYJlIav
ueQV0vxbsEGad0STa5aiQulp51otPbXwOEYsh0W0gGg6jG8h/hbjceJh3bziV/nH
LVTfh+751ib0Qjo54bEX8g==
`protect END_PROTECTED
