`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xiy9JHa+t3GIrh2tqgDoghbr3ITB0Yp6RMcIx6GLb0gHvbO3WfL034KQNLOvAyCk
8Id+gp7l8GMd35p3IpzstFiLJ0xDdI4UAhj3kmxHJyKhWjLZJYTF/8cn48s8cRO1
3eguvOdLPWTZALUv6noMf2FsDesPN+WQ27/nI1UiIwZz8p7sI7aXfn3Ll3uV7eaQ
9L3sMduwTlknrhnn1n9chJRP7WHU75WKpaH8jYXAku6rM4hXBccUYTMBXisXZwMy
fmXqut/nJ5x71EXWVgzqodVlFQ4Z9LFhHb9XRJEZQ2AZ0Ko8a1OJGjAIHRYfJScl
Ytw1i1NA1Aji9hs00BZxgPnbHiOySPHBg5yFT/tdVcd2Gajngbs/IOkHcQLXtFgO
pKOH/dwvQXfVkd0TlLvkyEGh+JvrsDdq1/Kb3AoQcb8HhcniAij2N5RBGGsiVAsX
L36E5OcmG9NZHZVJQzowYD+7bGC91V7eGIYbATpsPG5OX8c/rI34SpmIVK5BGISO
eZPRFgeJJwzU9Mt8fjs66vxUEt/w1s7D/IrnRxTlJNjoMM6p2fgsoL2t1UbWikv2
F6ZfTrKxDlMlZMav72rJVJ6LOCLMN7uqr3WVeXYJ2y/ZHLGiVNpRuFW/kGJt8NX8
7EIW3GMn3sfkYo2ipRRx/rEGcs9/F2TW3PJsqyGP45s=
`protect END_PROTECTED
