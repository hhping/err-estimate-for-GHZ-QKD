`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMTkT4yr2qkFoxSuXauemueX360kBN/wyTliOToi0OUifQMH7jit115rj8op0NKM
lb+ddxd9f5i3fsd86pzvqi2y2t6eXeX8jbC2SXmzRifIxkgAEOy3kX7njxtgq/kz
hgsjZoLmLbOwzGvOtKqacAZ6PdBDlvHTq4S2qtqFmat269VgWlIzARUF0Pgj/YSs
ic1hsPo0YVpeZ+At+r/D6rGAHc5BiQmzgfmRfuxPsa3X1+jObNawoQ0IpXGV5vD+
+yF/2wnsv5fg+oXaG/pgt68ujkGFCOlR53yGwovur4H9E932dBVbwZyh+LCgskkG
9KBeBhjHo019XTLmmb5xYG3UwcbJ/fTmt5yTcl5gADx4xH97UqQxzHPhTwDnOzh4
iuuLBYGxDGaILJgNlubIVignLljJttXJo0GqdILh48mRH0fYeDugkEJaR/9dSMAE
GNqRPWJDeZz+imRpHtW4lKTrkntsa6+8Jtmup/OMxAfNblwAesDy4UqEW25rWbW4
9F8Uk7qvjeM38PJFDs0R3cSQ1CeT50yVyP+fN0tzWzGGRqvmk9Cm5sPeJ+NlWBPo
P2QXBagfRPGXXkpF/RGP4ZDtYKSEKsHCFM4wBfUJZt6Eti8F0U6AG3mwgPMLNUBA
JpmBu0N5YhCdtm9ZpMSj9lScQKhbP9LQhfkL69zLTMPkGECKkRLeLQkMbRIbb6kl
75ZB61DYzroiVZgFVmVIBSQ0fGvE2XYjTNeJfd5pDaGXUgOYIgBo875DiN0noh7V
7o7CvYj4rHB1GGsJRXf2UQZEx8A/AXeWT7cX1IJFrA6yYqGelG4dLfV1GJAi64DN
VEkuzfp9febMRkHkx0azNuhQSBmcetZFgZ4coYnj3FkHb0yln9p0i84neagBaFZi
BOTP0136XqSYz3LGwZEfWZGNjMWDEW+9Q8hyBuXVtU2DDj6Y/k+Z6esDOCjvkj1T
69oMM/bFV9c4anFgpPuxvXS7UD2PVYRqrry1NnzHEz+/fnyDS5lEUjPgTzNIfci+
tTiHoWc4LuvGNYwAvEVDXWL7QFLGf4gJ3g+ZyZsYP7gPHM2bPY23OOJSRSycqzUu
rH2jx0+YFK2Jrn/C7gFmiZTbMpjeXUyHF/WuidOkxAu2H6xoHKoxpKblyRPvOi/6
Loo5HRKAct+HOdApT2v31V5PQG3c9ciscDh8C5vwJHCxaWrrVuXmnsRHeaN9PUQJ
vvmuGvy0Vj3oh9FgqpaeSQtIHSv0pWN8mfBC0gwV0eLZhdjC92aR+FObuQ39/RU1
RP+iCaRB0itQyTIRq3gu67kRKd6Nu3yF1CCLHVOiEkMLp8GVGsAh9uP2WWl92Al8
jy8d6Wwr1x8qdMFn+V/NAZxcO65Ac0nHMjxsP5qrs2ltHmSMTGCa+/0YlFlsADrL
GSeo8/w17Wp8cHcHihNZ35T1cKvykQ9/KjniEqJC8RjCsXQYGBPBRysrvDjQ1ZsU
xQZ3NYp9rNDZbgNq6w1eHTrg3uuiM7Q0bc1lwiEyJWB207B0NEpTEe+arEHxhtyL
mdGocxqYLGebY0bMWOc2cfkomIMTLH0Yqfs65keYr4Aue86c7gWFT76XynP2Cjqr
SXVyLWvdM3bbVCywrFT2R5/kDK6KlamLzulJInTSI8vSAuj7y011oUXcaOjbJ4di
6t5ax5ghgOKr2PeKE31p4N9V9tvjrMCvh3MW17By+wAxA0BFN2H+C/s1I/jhHnxF
Q9Iumuq7JwRnmYO+nVn9jbEGOtjpHibFcX6iQyak1g21JPHH2IPapCcXRdgx3gcq
8F1rKxBqQ78xht2jJ8si38JXhkbcGzM/7qlR5l9ukYhuNkNsIyzzZSei6gUqH46R
H/SE/1ao1DlwrlgxXaMkxmnbN/MJ8j7i4Rxn9ysLQLv180OC3ZjB9uFNIBmfD2g9
3hymyVv9HywOP9dWUw4YQsfjLkxhP6tMB0Wix7cY1HmmFaLf20Fnsg2+7dcxvDm2
6V7XKSRrwalzPmRehRtKyS7qOnySGJtLTXuN/oPkaKjBtM1W5Ex9i3GpLvHwW3SV
uRXALj5wHy9ZALo2pUqas5c8TIqJxWB1AhrbOAG/r5U7Sh6suQ493klc7qU3F35g
73tnv7xhu17ndsnxLBwUSZSdwFp5liaP22GBZ93Ok/mmTWOl9k+D5y1t5FGKGXAK
C5ZjXheuzNuoS8rqTd5YitBDLCf01OLjMPkNjdoMba+cU+Jk9UGszRqP24Tf8v5w
8zIk6iGXd98h/YvJe9G7oAPVNesdihXRRBF341ozvSMeziH2wPciVHIC8aaBb04F
9nmQWBExgV4qECOHJY3I6NVj7NNMHpQnWI7ClkleP6c549xrnJzt4oj2Mh2bizZJ
XmNjaNk+7V/Z2+UtnfVqgDBQ+fZ6+SdBg//+zX3jcaotZgMuR7LBRJxUXMt+BIQK
dCNDupNMtuZybD/AEowW6awBP1CeOoG2MpfABy9WwSj+APq+OPvFt9UZrTumSXbM
ZQlgpnBc6G9DQMXNHkgN/DLoQK9KTUoFBeFlcAyBcEapDGH8l26cMYFK16kiFvjw
hc0NEd9DOFhEPQtrTXe6ocAg+qLCOo33WIAK8uW85A/bKqxbKYcyZtSvl6fiatFr
UgUocxOORTF0CLR+6Xdb+ia3N4K2xhAAi45ENj9LNR1rg2DMDWRaXW2u2/fLbZNT
dvFyMr4yZe2MldV9NnrOPc8YHd5X+W3NlQaMPag+G0a869X3w3+ZqQSGn3W4hx72
EG3XLc1eJXVF/64CEXVDJIhExii2hNzuJa94Kk+RtQezNSPQQ+/H8X1TOPYSFLCB
p+tyIKvlwcgQNrZfAyoVCTYhiosNrZOr409XJTRar3wXjENKCpcUA28//qLwGgmW
XULaPT24WHnTsr3hDPHu8+AtdsD/JT+xIp4kRiFQTrCQbfftCAKOvOHJCf71tCFv
BZQjvr5dr8hF4fnWA/PGxgWq8ZbwAA8XELtOKKOm9fhlUWC0D4VUZvK5/tJqnMc4
kZiriIJ+chLysR1I3BOklWcNkrhyAdLQs+iXG2jlUfKHUHRHMwIH3j/20/R9Kq7X
9bGrSv6Hiy376WrWRr4w6BVbZJTHOy+0D3IhfZXRz3MRnTH5GBXiPDhsnwCUvkJi
HhK+uE+lxhSs/xNx4IFlKZKkrKPHG3TVkkNAGFNH1bVcupbsKtHt8tGE19Jum8Lv
XEfZxG5/6wl4HrFwqr3bRs0LsrJVopby3IXINxAhV/rSSCkiEpJxqcmyXKVSclRa
rV8j2uk6afmj/laDBNcVjO24zE8tw4PoyBM4rYZot+gNKTtxxtkyTXCZoQvOK0jC
vtMx+S0dQvW/hv1KRE9wlxELZ1Ymrn3ogqlnC7y9CLRpBCWQASFo/Pmll/PK6XB4
IwF/RRFBDAi59+wch/0fh7i9HmBAVJ02LMdXR3WzkN/moKXUSicP5eKgWmZi9dhr
y17a/BvxzklF6mioN+M7ifwf8iQGWG1FL7RTGHflUh3mxbfZvVTAv9P4JLJ8jMNa
Cr47imeHWsXTAK3fbKjm81SjhFFrZx9csZ7vCsrnwexuAE6djb/QjqvlrP0GVKlZ
Bz9VT9/iJDoG3eOA0nPjKBH1HaKTmmFkEY5tEwtLumUPQbPnzZf4ov54QyqCL5mk
lRTLRKVTf79hDVV65a4gBJ4HWnZtb5JN6pLBnX7084YWG9eB05fTo7xgqxI1UY/c
PwGBz6pS57rEbO/oBgoDeCydihdixsggPF5KNBvePnoU5VSq69saxtOPX+4Sq+6L
+c5a7pDrNH1S6PlAlOW4y6d40zKqm+awmYWibeoGVPYx8EJFfi2QTBGR3HLaQnt7
+klPUOfI0nI/pbP8ErQEUN97L+Yi+2Mit+QNra/AvL49faTyBesT5R8a+ekxE9+g
Fvax02GHnOBT02EbgmrO9y2NY1EuKyLclxcsJvB/PzoEgmjCHdjh+uLJmyAhi23F
HZDa2mVx5EmOjZfF5+kgvbavt8Td8gI68oXgT9HeiZ3SraZpFNCvoh5UQ0jY3R/O
Rft44f5x7bTn5S7fplnl6BOhGzZbdr/A6ftP3+jr4q7+D80GlXH1HmWGZHxhONEZ
2b8A9h+O3eip3ieJdumIuPlC5K7ZCAQ3PfL8sJn0cWTMS4afLjaOS6o27JHqIs5U
Pf6V8QEcoiy4cKMNja/sp6RCoeIWw+A+0KYpXRA1mEBnDOTwZTP0HFUhQHFKXZ2q
qocmyMH+e+PF0y5qPD1ZjeYOTW+DY3clxJSWNJQwHIEqoeTKKYUCn5zpe/89fo5Y
Vj66AMceDWWuuEkseyLxcemfVu3E4jvxQlTrTsyrwPXmQtjlpJx+vGzpr4uZeKo5
OUkMJre/m7wV9Sk+zc8D8NPdmZ17+0Bk1nSlC9Xx81g0ZtU7dvPNdhYxQw4abFlp
x3vpBXOShpZTt54R4FUgyRh4ckwoXOX94bwE6krbV45Ah3dcvf4sA3tA3rBsYGMt
lXIlMnkn9MsqNv+JOOryKY3jrCOvPOTvuuR+Ys2kHD/z8+dQ41dxRxJSTWEcjID9
1nIfRPdYvcKUTcu7lnIgpj3Z8ukTqzTxDXQvrYCmb6Osqw46K8lxVOLuv0QSz/zx
qTwkUHtffxrxqCUfwhr+BP/DlsO/0sRlL4SEftpCtkBy4CnMPafxwZF3kWCpaxcO
W1THrt07J/qtYRwC6cEbNFr27bxbPWlOfB1oiMwTuSkeyxRiHhkogDa+Sl/nW/BB
X92KnjmCc+Y96j5fz1OARcPQ7YQOKDiAXl/Iu8rftn9CCFLqdK4uHtxmiolSv90s
QIS0/PhXisNaJFX7l2wq8ffUWz6UYrhIzwPX1eCJJYxea5qCPz+FZ4wtlRbiCpLl
jDiWqN6QWyxrglNquxpCq+bbU3cUN6xagAnbsNVa/GPhhgTRh5cqXtK3D/i5SVSO
K6zw4Z/FU+1sAZW1zL02x+0upaY1kjmmpDg0CEpGw7godvFjBYo9Ec3DcCkKnJsJ
WEL1yz1t9QhePbgqpI/7wEMeCeEO5mvVNzHnXRao4g+ccBS8CA0x5pALHRp1zi3g
/kWs7Vch5j1aSQvALxKYilYAjtvcPqaaubppTl++nVgnZLs6vfYdvbZyORN67R78
nahwvb63VEo3rzDjKWYZeGwR6pIQ/shrfFVQL2AKT8vrkaeenKgXpLQZ6fl3H8eS
8+pR6nsusMOVheYoUvwTpXOfunwVlP0onw1evDu6MPYTm63N5TA2ca3ZmDclXBap
uiJOIEEjOgLS0ndCtE8XY76E5YMfH0TIaUBh63PTqWoeIi6ECn81/XMaaOjfqaBZ
Szx4dI/dz9QyaF2lZBcKCMJEto1+I3NAVeQtdfMbj+zXq4oHMlDuEIFYKZ7lLwBt
+N0UNX4206uzpIHBbglSx1xw15P/VYvmieff/dDsLFANPb+f7ZWXY/gMCqJqMfAv
qzhwjpP5Gjl939y5uOIfaOzJcWVE8WDVgXYJZ1JAr09Lwnc4av46HPj9BgI/rBwN
n2FZWk4n9+PStAoY1tQx+63tTGwknUOqnTy2tcLn6IUxMNct58lPVW3QuIWI6zo/
fL+J3UjrNa2XI35Zzhou1r2xBycZ9558pSD+O1sQOFzZA29nec4Yxv6wj9IopFrF
UOcgYiuFT3HA6AH9Xlsyac/PXFd+KmD+yI8q7rV1xfQ7wmbob3cTq20ufRyejACd
fvnYaq9N+Z4zXyoGfJXXTNYEr4LpOEgR5L2a+22cf0TrXAyjPyymEnEcuZame+6Z
N2qyvB2WQz4Jgl7YUt5duSM5kk0qS5KJ7DBMAj5CoRhO1ref2SKc5ZdOJ9I6jOgA
WxkWNMknNcLFdf/NGhhCtJAD7QBXXm8WVEhvKyoO1xWIdGZAPtXlr4dnoRDz9cgY
fyFAXDLQOIZ15TwiG4Ocr1Da/gyYHX5G2Ab0GAvBEaMj6oA4tq7U5Zhn3q1TuXOS
Mr9isTwhMoUgLwMpzBoCN55MLpGXVNqXhdmLT0wo2dEhVoXPsnzgrIIxVfDDL73S
eJMSuD2OifKcU3mTi3+OVre70C/7VScy9TtacwgC48etAYNYRWdLvJYTsPLYZS8b
+aoPt2uSHFD4XatqlUEouxTM9ucv+JUfSd5HrYBeeM6PDLwE+630ZQR6PbYz/6Ba
BkLzF+s7evh+5ed50WX4BTS2nLVtxGlg+MDHfB+fXDq8MBqqe2e1EXTo8WQO1RUa
uuVHBJm/Su4g/L7ac8pKcdYElTUIfV967blm51fJwbX+pwkrQjUCcNTSTaCCEAbF
YiuLEnZlXJlc17RPujP3iRPtBXfbz/Oeul+lA7iq0+O2mNnix76awpmSIKb3t+Oj
WkJrFXboQgbGctV6XxHveMoz2p2/bSPhsyBwnh9f6fQCZc8conbHLvtPssTWtkXm
XFmnytTWmcko7R7nqDv1/nC3ukqJwPtY1AaeevePeF/vpJWWiAiUXWftQCuHZc1Y
HIAlImoaJ6OJVFuSjlJBUfnOgpzu0ZWGgLmsipZHI6/PI8rLJlX4wKiRcXIZeYU5
2+oUJLf54yW+cEJDi3HVgkhHxkHAMdHM8j0LHcKLb/9vb8rmLtGzKu5BZgcvOc0J
ShM55hhgscQgiy1yOH3t+twWtkPnst99c/rkSRcU92lR51EpvXGC2d0Oe9ZjL1QR
PskYBMeh5TOrlF4vudc4G8TU4SuC3DNuIWMgZ/5L2ApvX0YEFjxHABgPrOq5ZGT1
FRLZgBou+nB4NE6wlGYCCvW8z8yRfuTqgt1LAfrWyz1WGMEOYliFtEvjsInabbBI
hLnr07XYWRuRa7UeFx8sx/IlC8Fj/LgYv5nmbFTieAe3FC76etJjX9SODkcX68uY
OAu+EJPoyzFJaP4uAXCho63lg7OdMvqkEeHRUTAUxAoHJW6nqNixTB06lTHZ1x+t
XdPmH0Z4en10+fUL8I2aESDIKGI6PNHHwFJla95SjGPeWi42jA+59qe97HMiNdEJ
n9s2nKLmQWSgeCEAjjCb6IeqnijUIVysib41VFI8D2qBIzSL411Vlbah/i6eueYh
mOIpTT4T7Iip0xDQW7O32l45JsSU46DcBKmIkh7kLw48vZisMLNIEkG+o9vZMp7v
/+QVQbWlZ/9lyQ6DNL+uxEcnsuTqhD4G11a//i5XB5iBf8bscNrpTFhW8xKjyFNX
y2dx8PybzAaQ7aRjrr9XXEC1mRExl7JwxR6GAg5HWOHBXxh91KIMQ/zilKxydjkH
vc9TXGb79/+JYuSwLtUTTozagwU/PK40Bf4JmUsv1VA7kSMGg2rTvDY0cwKwD2TJ
Z++iZNnUigz61WkbQHILViwpyShlw4+DHj2zfDJ6tBuCYsBUUcmsgvJvViCO8D3j
dXel8nF+4GzpT+q1WoD3rerd5Cf/yPRvM2XzPLPq/VkV/9+lhMGTm1Y6GK7TIIe3
V7SjXbFJoTZmVddV8B0fPXhqXS+MbR+/WwpkWPRClRzr9JyHHuABu8ew2vFYwNwE
0VucRNHnfgeAGJYZwfBtsbvU1l+P3kY1QbekAaIirZRRFBE1iNGV/mzYRRWaZ1Vz
ooN5S061uEZVfxDuyRL/bpjL3/ItNaEslEpxUWGqXlSxqejE5YNcUH6OGr5jdtyW
sEjD16dF9DgdnSPBLTYAmq2NgFcSrwZnuKjAKDVbLlZwfQlIG5lAgiWlTJhbxBka
pYPaSrX24757gM/l+0IVPeQKZOJHRNNHt9nqQHtHIriudQynETkms/zuBc8jrXNQ
gQwbfHMzjoqLvWtkDnkAYZwAEd6qXO1HnnQoDR103+995KM4aaCFFNXDW+n+rQoH
2Cs46vhaAf0NRpCJa61vdrSp8WtxkV6S+wX5LmeJoV+XU5k/nRDWkVbjGWalzjDQ
66m/XyQtH6NIHW3GIOcdqdgMRvD/1nRoAo5fyZfl58pKto47bftQ0MZQ6H/z77fs
yWd5yv3iRv3T2htZP6RBR7WIOOx6Ocss7XYUugsGixpBwqCpqp58n19w+/eEjjZD
NpRCbbPwBeYNQcfzdF9rwTMlAhc2BSU9A4tLlIThFibfcFBYiqlZi7w3re5pcs3o
oqrKSeb7ddQ0IedqmtCOpfdUdDWz7IVo8admtSoI+Kv+1FAXqjn7JNlV2UdkFNEo
2n4nQH8iTrAg+Q48gIvVCQleixp6hC/yhnVAVnftBuFKDBzaV/+qkVPlip0RZyMn
XtWrYW/zT2+nKHDNhw1capzyfApYAZSecB2piPH/zNdyw6OPWQk8VyCAXBczH0Ie
qxM4ryMWms5Mhb+5/gdMLF8o4ro8KJVfLbgLTJ5XsKUoZU3NTZlECWKavdqJRWsG
iE2Y2BGFg/ZM3ua9lxRCMVx9v8EfveI8D5rFjxDbpElZTogBocLwzWkv0zCvyQMd
5N7m1gq9i/gqg3C0nFNh3l4j/MwDHPSOTePygeEfTaJa2aM2HfaefwO0J4Xn10Jv
yJx/LRhDjb5DbA03itCnsT9oU7lM4wyc9LESnsgHMbRX9aI+20puOhr6X3fngWN2
6TQ2f9KQlinHGee4drhVwot3KA+wAoxsL4axSlNdyeiv2Ft2xP3ldQOk029w/iEe
e5kuUwzQ1LpZXtGx/k4PO3zaeihp/bdSj7Vb9SwrLAh3l54vYdqARqzwwySQAirw
9lx9e3dSwjTZ9s/PeFwFET39UMjM8dFqJDByldGjciRh0TpbzCQjEao5dYw9K8mv
08zeYDuruoUl7b9ih1J1xjcrK64oDatLILxRO0tLW7Jj+XhkBD4IRRY6/+lU9mq+
BWFAlq7Adw2NoLYb1fv5zGnBe1BWLOX3RQOxLu7kp8x2vo2VGGP6qaepwfs9ROqX
ykQsTrksdTMd1bSGCWM73kty9Nb/uy621MIr9L65rx9EQgtLcdeIxHGqvBDDKSZc
kySJS1AkNwTMhbGQ77/md9LP5m9Zv9xtWTSY7Wpkn57dXx3/2vbIreU/+FVx6MSv
jXeS73JnMDqXABDTaZIjfCab+JREX0ssmd2KygLAqbf+S+jA5KbEs67xVAhawEvM
bKGPoAFKOXUFbByV+Hjt6S1xtIHSzXeJY3uc8tVs+U7XsoKqVluXXqEILa6DEMiz
ASqNk72eaj2cRFQbEjiIsHA32b5Bh3Yfq2iqVA42Imcibutg/mATdXf9zEtYef9O
55yUoTcIHtimLpeceoPBsmQe1Rc0KbtL/ThkFsqGoLDHAVueQ9WJANKvdpkwmgvd
0B5Zxb4O7dLJv8HD3Has3sE1f3y9WUHhjxI0TapHc6MlQoMiHXsEfYXfw+tczu7t
N6C+vpK2iE21wACg12SqLB/5weSeDthyRn1hmsP5lQXYmd7UbSOUD9aTqzXfUnj1
mCM9pCziRSO0Fg/eGktuz9mO/2hbjLC2TUlJdVUJsKZDgIMAXiZEZfDdlChtDYBr
fbMuXPzUUNBlO1feUaCLCdoXzOZTpsDfk7cz+i69KZYxdMbRdMVaHFU+SefSfIDH
7SKKNuoQxTo5NZXRGh6xna2OFGnWIXVYe6n02HB/KrgBVX6hdWpub2MtPs5+1RXr
GmVi800dQUbNawKqCy3YPZvNIYEe/gHNAmBSy4k++sX0eYseTsSlfXPs2ymYZfxd
cPl1MMjSMTxuNU4LBjSm/LZ2WmnNaCzcpn2wcRZABzlcqV31DWNWrl0JJAVWd1sY
ljdHAwqBjCwCu/rUD0bmiNjvVCd4prGLMq1Kk6wScUqwbMrDv7WmzL//EHh5eN7n
uhtPfz3n4z7yeNjd9KfLQCUMFY5RI8upeVVryfTz6Wqcl/kYJcF47fJmVEpJ00GQ
h0M4fPbC3XqQzzeMh+H7ucomMFx8A0klbr4vFLPgnGDlZH/pUEE8sFs/TJnHD6hl
P9hKZZDaC/Z8Gy8JpvdHSy/G3EOzHIZyPRvRRmhQQ6hu2bPgyx/YLbSVBwPjWV1g
ryVFAGLVb5tsNwdXDvetEm+lrBiktW2cSaiVoPcO5Kax7fGQILnkUNyd4Txvo8Fh
+EehvdvqhijfY4NBERs8z/2PVgCudmEKwqOvy9sN5yqgikqLcfOFK7UmaKDOBj/q
JkD5HKSS6S0G5YyUKclFOjEcoCNMH2gIAc328OKH3CN3dzSWNiFSCj2yANinMgGj
25W6Zg2nOQloVwwHjBvAmvsI5jhkQGFeK4mbldrCBnUqK66FV/7518+I2AfzztpH
dnIqXFD6aj1AKXnxSOKGRSq24hfDHo49Mq0NA+dWu7QmyfxvhAdAYZe+n9SXprBw
+X5+U5A6os63jQsywcbYvYjqQT0h41+ufBkqzxKc1XT7zhsqiDHy8x8NTsJn7ITL
mJ5/6f+DU1pmKjutJXQcKLkRFYoiA4elEq1dnFBmwl3b+XbhDTk0Ujw4oNlx96pY
NYhL01qLtkrqKkJ73RZyASH6n36VKGdN8O34nsJbKFd1OVaha7WNJ82JzNxn5AJ0
el6zAa8tt6kuufNgoWPz/j/DnqEpgbcDvcqQwAQwHibaME5UrRIDDZG8RZZ/JSB9
Qywp9XpHGVltyrxuFvXlP+w42Cw/Z/F+qnVR07kZH7t1Xxr39dNjpiHCxH4NizWq
kn1gYULbV62+DzJ5szNtJg==
`protect END_PROTECTED
