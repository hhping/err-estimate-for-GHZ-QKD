`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuhW9WULbcjBPCV7xlL454SQAOYxXYGiTB40Nd983SYNtSpgtZTpmmeTfH2LchpI
W+jN+j/ZO/d3PaUksUcEUOfeP7NTH3yHkDgCwlPlrEsLUsJyPNj7ZR0FO8VsERhp
ikrEpEou5qdDKA0vxzrVtAnXluwpMrKd9yYwtk4jsRjfmE+VVPYqQuMMv59ahZJD
86gC61UpD9a4XF5PeAT5fwah7XGHScKtt0KApa4Ij7gXAgKpO0eFGHte/x8M0Lj1
mpYglLTdx+cuPxgYf+PJhbouNIik1KHYRzQQolyyx1ROD0ME6I948mSakS/u5JSN
Df/eohJeEfxyXJwHdf+vZTuLhMOPJHrazo1PMEbRUwIOiMEVmAU9vcLGP+NBKGHE
HeOTP8hoFoggsOGa3gUd0nPLBWYU4aUUW6mo2d29Ko7nEeiHJPJy7N8Ic8SeowSH
RzBc37VTHZWH9V27csJAV3OjvQic/bl/sR6ObvsiqkONsP579qpXOE0nNplSr2o5
RGtqPET6MsJ5G1WtbEDjgWEogn/S7vdq5xpJ7bd/P+virxTM60TxSQD9yhtaujmQ
4QP+KJ0YNijVltWy2BKsY9cpj/r7/fr1DRvNqoSuZFu2muHZMyXFExSjPlkiQES4
eCDVo1UccKo5RgabclVV7F5sZ7f5QG+PuYJEtKat8uZO3riMxciEEj7e8/j1Sx09
JNvAszXH0IN0TSsbxa4yoCVI4kkbnbFQE/hOUgpJT/gew2Ndd2ocY2CA9+1RkLcr
bjKXyOGCtUTz3DCG9GeiXh6OpyYlca1fdVQ7CuTQqTJ93TRWI0Oq4yrOFKdM1D2L
3X18Oz33lUTltuqLMsyUj40mLCRxvi39WOtiWJLYtF8oVDl3OH5+PkqBDtyHu3eo
Sg/3S8cqBbcdnTRmivgJuYNHfjPgAKMUc49xUiGeN/B5gF4J5X7OoVr60LfNg44c
9vlX0b5Gjue6p4+kwsSJMeWsskUaXewHNaWSzG6mhs60ClFjBt1SxsIOzcrv1eDR
zznmn5ee1Ur/1lXE7hki2KZFoHf1qD26BFauHammAlET+MrkC+dLuH+qtj0mfkBN
6rgWgg+UT+Ge/l39DnX9ai77sd3A10/TOR3ZeTPe7aQriaBeez49mwhPAsczP/eH
dMwIm4g9ecUr44Z83puac8OhGfdUWgHbYr0Zd0ChGAkfc51eRJ0oAK9SRtLoC/ff
3SiogC4VPbrdoZhDYeTYRNataUt9Br5viwbLwWgvbTspUiIvv2BrTJCPSfNXb5WJ
LJ4OiluQ4y2bzUov9ZVYa1ruLpPkIdx7pgvK7Z1fwgoHbWGAOi3Xqc5b+C6counk
7VxEBqvUTI0czWcPKI+2KOM3CKpJi27sVtxUrXD1UejQpw7qSIjHOPW4YhveLrId
189cOXFg7L43uWVM6aN/uKmGR5MqBLphjFkjivLgfTo/hbiQGxVWEhoxZToeEGCD
G2XOhXRNJYgRGQVwmjjhZoAqsL4kD22tArxW1bydX1Enfaob8SFURlXTmOXUR2Iv
NzAkJMf4uHSTcb0yE+CQWWNQj2wxwtgP9DRjiUlcB+Em2uGi41TvK4xpL5tIBP9L
we7AbBGOcqBYIz8vpkx6t4kCVab/xtnTbN96UR10nTOoz+VSvS2WUfaARr3YIpD8
EAXpDspSyH+8LruC5dCbyZbAzMWAHRS3W+LM6WA4DM7CzuEE+eRAf/quEPtYsIZe
hVBtyJZ2AxnGAJDC4hqTKY6RGGfaY8Jj2G4c7NXIc+qeOQ1uL3jyj34t46DGzsox
9LxGo4fVRdHqJtzyyaYwgu3jfUuZu83Z7zCCHSbXcMBug3JMkNnya7S5UGcHgVje
/Eh6ialyydWrxSyGqsO4eKp27G8z4Lu+AmAX83YSNu325RjMe/+Gt/ENm52g7kpu
oLDirzXHFprgPFM1hVNTOSNhEx1FnPmzoDkB60g1nkNNnJaQgjeMmlnXzAI5iH5t
8JzpmZkzIvKMVftz+bjWK79GNC7iMptn3mTCsnNBKnbrYq2LWm8+Ym9fVmDCCm6+
Hz7HcodvquZ1fQ3KY9xE4cHb8nmeUOCwZe62giNa+uPT/uL1Gfy9UlJlJcS0F47D
ZKfoypnBo7CO73PZlSjTgt127JglGy87p5vIAhIy2/lX14PKpiU9QKfKUeXpit/R
O7sohvixLlujy8rRlBwbPW9+Zn60vhCGTUIOG4RCDmV/fAPj3KXiiTgJ91Igb+bM
uz9qe57vca8Hluqiku0GIOQVWrK5hnl7KuMoK5IJJDoFTxOkukEZ98hJ9dZffChY
elaNEQOt6FrJUvN9sD6MGq5AW0fLx0slDcjMHZ0FGLpNNjnDYse+gj6iQkHFAy7K
WgeL4Kiqcg0LBv+s1Lce4k/lqJRq0EJ1+r2xYXUKz6naBnTheAlHGPUhJKiq0aMF
wrDKrwNMWIb9ZEfgEt1uTDtlW28nY9Iwuh/WqVIZLZ/1s90tO98fz8lrV77Y6U9A
PpIMIPMgE90jh/NTcEQUCLBkthotd8umspq4wmDyj6obFOKU1NOu26PpIbIMihAD
yDBCEWPLwTUwULw2y5Z4/mrYaIdIbkv6JwxEEGvLAsTbMy7f3mcSaM4/DO5wErdz
pwVX4e/AjEcSNBIIjX0j594V7tMKh1Ur4udKhIlT3brguyl/jb7NOiSwz6g7QvlH
247teyuj36XGan0IPsn35oOUKfrfDF5TAg3vvlMwP3EgmtobsrxuhblC+/ZbhNia
Dw8f6v920fR5UujIFI5w3vKiKKVSgeQcjP4bFXw+0FXZMjCHqUEWwrYkvLHn0mlK
N99lAjFdhhsNkDbMKB0BzEeCR3edboYqP5AeIrYk2zzP/eYVELMMFGt3GUaIrJwJ
Dj5p+44m5WTlmkM9nuZWNlb9cacr2+MI/p9i2zW5m8s=
`protect END_PROTECTED
