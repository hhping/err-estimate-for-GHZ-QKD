`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLvLmXChYVSXbfDqs1H7SyE7LYgVCEr6tl8zkW7dJZOicUmmQU/xGxuEGg4xPFRn
4YtTvab99zLzj4ekBGw3xyumrdXeke7+MFjaFOiVtnvLOYmTPl/1X85IOlUoRcqp
KjeYy0sbJL9bcC4udXYLlqYzQgQ+3CfoZxQEKWc62JGTcw8cs885ZhSAhVObC9tn
SLLiAVLE5eUAh3491xzOudbMo8Rgiqms3MERgLcFi0+qOER1zhSbhnjNWIC9lkgz
dZ7LDpFNKTnJrP9e8zAAeYHnp7W9O+KTpTNgMMGyB8OJRP/ScdhBAjRehzrF1Qjq
e1I04vb75UA80HY9WVbZdUogKj90+rAGS85qG+PhZmMuUdd/Nj/h4SPhF7wWnB0v
jSj0vAQBMuoMNyCun21n1Cjodn9Lo88w4+Zysy9bfgs=
`protect END_PROTECTED
