`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RoQwCvO5K99wuHix0U9WWFgkxF1jzAbcyG5ESwH3fEAs7sAKcln8vXs8jZhtY4zb
+JPXR5BXpT8/CJmrTnoUMVdR7NQBfDX0444rQiNPWLEs9B+rV0Y59Htrd4OOmlgq
XKJAEDzrkFYG0+WPFmwviQSpYBtmw9kNttYzaQq57LeYs2/9Bj8xKBq8gyfuI4G/
m6R0FRzAH9YEP9RoW/U5l4jbgHiLIn/m9VbOTECSeR17pgndZ1Ce0MlPp7Fg7dlw
OXDXWjRlbdzFlsLWhFVyp4N3uF8krvTboTBQaLyEFg6UUH2IMLWNGJ44Qi2UICdT
KmzJuafG4RRZgLq0SikaFw/amQp/2lRpNX1enbLRjh9rcTkVNxWnPXtow+AXVM83
POV1DRbpQCXCtll6Z62ysWO9CnLFNzyQRMXaKUdYOynfpjiseYog16BvSTezL8V/
EG38Xb8XzXZ8DuQIaXXpnFE50HoEz1u2pirsn0QsAJC3WGnEJoACgexXUV1BRayc
+pruKbNhDfOcH+cUefzYCWwYaCQ2rAVKyhMImmFlEsyeQDheiRjFdi3++sjJfjng
yC7Q1aMQhNvtrBmuBCkJeP6D8ZsT9MZ4ODpZwPMnwI8ttpdLz6Zqxr11rdp+8B+m
GjIWILXsOLMDhWWo0WOYpQSoCNh5qRj5G1cV4ovHpBsBv5BWQXA+aEUZJhiGhvxm
q77OLvarF6l11pI+Bh4aTuHIaUAM5C2RgBE2D/ui0vvyrSgn2ueaoP1KLH1O1jWt
`protect END_PROTECTED
