`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsFKXwj0BkFi1azP00MH7yGCF54hPvT0Ynhq3yI/jNDH8Ed2tyTfcFMJWzaToB6A
QzQIk4UmM+Tp9eLOatH44E1pidsM12WqfO66iMm66PT24VP9VkgVS6sFOWl9WuYI
UVlIpvH4PufDnwBIzoABl7jO79QoXfTeQjahwqFKU22ePKc1wIsmcUk+lfOpiQwG
XBrPgH14yrsGV/E2r9RWrsAAFS1yazkWlxfkTGoHOAW+nr5a/zaxYz9PuQjpWWDw
vc2zNc1vdPnLqrupiuBIyQ0GLqe5rgI0N6ryF12x9sAQYUwChItix4SeNKTPwPDK
MlSKlTvM9P5+1IZE62cmbkvXbzIx8KprON9Z4TkJA+7IABHJDkkqxCgvVv51XF9J
N3d1FY21mELGwRpQCwMGjziq6IlHE3Bcw8CqbfH6zEKeqf/wlEq+8WXufPp4YQdD
+ogNcDoGxvJTHaXA41wx9EH8SsurLdAi0vti+a4qQW4NH+wJ80+JYK68h9NUyQnw
s7woVT0xEG4cfa/1lL4xzWw0AOb99FMr+q1U0DwFumtrgb6Dz3QI/8lU6MUGBpeW
4n9wCtp/2fyLViQd/+MlRKQFoeX3K+cTcW/4OFua1h9thC60NhloETV3pwoKc87Y
slvfwsY7zeWc9pXYUJkN7XLnldN6sn6DeQparMpYVunZe7n4zS22SAbLiP+yRVlL
Z3kmcLTrR+g1OXtqDM7lid6rPw95vcTGtULPT1Ba/4G3r8vMU9af3shNzXZAfyS3
4dyfVQjj6BJNwerkBFVKfyr6sj0fDYR8k7uhB3pfbXmPLY+y+5C/z/hYBZFjtS4O
xRlWaNIoo/OkWC40vqOfjo15wkIFdALhd5IHt0r/sXzzeMfMCf0Rj2ALKsClIyiD
MOP1gEFcVp2qVARedFBlrLtoWnc7XuDPmPdF9GSppTSDlZpj0xk6MMR2du/K4K4c
lNGnl/IczP/gacBTS/FrdOly2y2I1gGFh2u3fOK4O30dhh8BJ4p4SVfFAlLuZBRv
7jEM8dwTSQuljWxI9ZjWa+oSnsztz3qH4Obyg5jqy3ICAPwOCS0Q1yHUbY7TG21h
jKw4DCwl2WDYZFet+W7H6WAxmi0QDqpgJL0cvVOYZBWIQEq3Q4TQCBL1tEUAW8jd
XSqEfsiqb7Iefmb1zpI7oVhYwMK5FnXhiknktgfO18Hmhi3hTN2M1acEMXPm5chR
IrnHlYoVjzZd6VahrnQto1/DSU705Vs+Zd1F7xZdhgK3+YT3tb7Y+sW65cz4O0ax
B5IyCNidLb5z4/nn6/C6lqXy7CjW1Ab6xYc3xdiCCJDvp4lvsG9p01MmjA6P4SVF
wJOUH9+AjDGD1ufZ0ygVH5lCOa9SGQtaiOyvLjW6IzLvf8NqgiGysKo3qTuCLCoC
b7AF5dYx6AUtictx5fOntEb715mQurz5lvxkgpz6xXiOkSo4Ci5rdiNGECYQn4MJ
f622j4Zj8NM1k43VVwPJVQ==
`protect END_PROTECTED
