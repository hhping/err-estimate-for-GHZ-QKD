`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbspLoGe02Cnvnp1cVQwpH7Ww7upMvKj8AXAaRfHHI9aY4zxppTUHRce0lPrXQ01
BPz8BqMAnSr9JwczEs4myO9s73r2jW+QNXP/fIwI1rGHBX2IEyFOM+4qSH9GKAjQ
FrkKD+w07VU+RCZe/sE+1N0V58MiOA8JT4dqMlSo7sgyA9VPfH4VaZfyaaeOcCE0
EXG2awbTqjxwaF3pPb5AynCu21NQ4uq5Yh6VcE0JQ6Nj6Swqusx+usuHuJGw/Wzf
z/Qy6wiSOvbg5KP+9L7u8CMheJ0s2NjD4AHAYVl6rO7ZdtPRp7wcWywgHOKJLddF
CqNDk2QfEmDA8yrLZoB5+K+nDGdTjJu6Ikum2jAD1P6LJWr3pMiCyrX30nfinZa6
JicEUiss8biQd5h7vG91MfIuiLXVB/bhfODjbJM/C341m+aNUIn6D31y4m6Euj9Z
w/hty7Ngl11nxoe3d3PkmgVK7/6NVkN64YtdXTt3bXfL1NFahC3ut6xawNFrsHvu
YJ+mbl5GUsYeLsZTbA/UMg==
`protect END_PROTECTED
