`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88wxXv5uz9hr/iRSoUUiEP21dklmqHmtN40f0KLOkF1AI97NBTx/o/vnkXu5XD/h
LrrF90dkQoPitX2dq78JUwj8GM42oI1L4V5HYvnrZpp255x+CzKYWFlqQ0iZR2Ef
CeogtWltw3QpG4B7S36uxscVAC9isUOVsa/RVOP8qsYWRy/9xjckrG1lZa8eVS1k
sbVuR53RwfBVus6JPqg0lBhgWZPH4GRRzklNBNQ10b46WXA2c3t63t4UyhAmgYn6
DxJa/z5iZjmstzYE+A7RCeocybb5d9BCclsBWgqMpwFZGkTWC3A3noxk687MEvRY
zKLz0OE8yxzbRhsA4tEfvugXL5VpWXSkjYdB8saq3iVwPbFzi1fMM8QHFsFYZwiB
S7V0bKYkOYN2J/jbUVPh0S6aHhWYMejFGbhM9FiCRSSJiuVo8DoNsxols3g0GC/b
ptsBd6L91DSABLudxm1DDi9gIiwj5k06NKmtc41Q3Fn7DP0zEJglW19KLnb3eByP
vWaXhFd6MnSFMWSMy3f1D3wS4MS37DVC4gF2lgm8yuL7u2z5X0tfJni+YeEU+LJq
RG2vaYULUk5gMR9uHlIfoafFw14aqK7lpkwkxLJuWuG6cgW4VX1HZmjtH88W2vVO
uFFMkrdTSIoYxkgIQ9lUeLLv1WvYUV8xR66oHHSKUK0=
`protect END_PROTECTED
