`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHQJ7fiqH1JGAhdAVD5rLZPY4NEDcpJzVRSanNNhDS3Km1CCbVyTQtOB6bm55osz
xhQUAarA5zQocNw9okkyWpsfWczrBRHMKHUB4btPKGbsgiI4ZNMjMNagkiMk8rsq
BQKyyFmRWK7rsD+q8GCQ+72NIOuGIQVjWShxyWWRu2EknJfh85LnVwhEpWG/W879
iYaweqtmN9zuZWTObWrT5MQnSDhj4YAjqXMrPs7Zyd8K5lLKw8JhT2+oskwvUhUo
MyfVaQeeARAhXwCMWnm11oMF0G37DZELk+8QCMSYlZrIHYcIHn0mId6XBuVADW/F
64Kx56v5OAhhpBxikf9RXMASQBxZYM8CG+TvvHTGnOYauC6Rpr3vA4qwzpmj0Ana
yvJxcJrK4uHjOF9fEJBlVFGmWpIZhhDL9ebfiSu6MiWsqUXSDN2ecOBa9+6KksZo
/T1Avbz7uSNDxBqIhb+bPtXuBmb7SGhMmRwQsgn8WgPzgBsdT/TUtHpdpmpghPac
+9EpsfuvdsIgGi9Z7v8zhxuyYDb/WYO/xJhVXx6Ilhyi0We5GzCzeIcjAT70wVjU
Ha/pSKJLaCujzQ+IdFlIy69dXsLdMlPE8yyORNKu2h0fHk2b2ijq/tAOdWlutqpB
epQk6Ukzc36vlkFfrELkKW4ACgIsRTyjJiurI/CNNtfZ9SVkNBrCfWpeOhOpoJO8
EMC1H7p0ps5gghCi93zV9WEOvy+Hy/CFJW3JbhOk7fAdpvkX23TTFoNcKpfg207V
4WkxaTrf3cCGGCeBa4wtEGhE29qyBxBGpmH4wZUr6zxJ147zTbDUfwCUGwNFRk3m
Xqg62UGzT71LzcQWVMEA8B8CYL3IStTV3g/nMgzF8xkZkTO9TrppwPxiSZJV+Rov
JIqTIG3J9DqNxSU74qp0zb/Mf/mNhaER9Ur/DdJdd+enLH06VJA/cAsYE9+KovQ0
UDnDziTcbEqfggk+ZBgwzn2mhSDu5p7cw1ifNL7BVFsRkjGZ9ilPbDillijqxJac
v0JtM4EpOPcy7ZZWGnm8M2ctkf9Dsf8k0R/e4YHKEoeaKiUIlHbJLnlMLgRBYOMN
0y8LDIQId8n4YzIOrq4WCLskhTp05w0G6e1GVsT004D+SKb4Gi0+ltHQAzk5EQhl
RC16o+7S7uQE/Jx1jwx7U5KsL5LulBMMXA9egBeBdH7WblzM7Pb/sGsKvHOtWoyV
x7q0fiuxPv9wc8DsheKSgw4qQxOE4wd+oG2WXj/1jwVZFbYC3ycw4CV8g8ThmGPP
gHP3AyA+HLw19/02H2bboTOKTscnIlFvRH2WctKbkE/tStGCTIKUaDkXMscs6Un5
ppbSnw41cCx18MTAZwbAQ40C2b5FvtKXZQRq5kVA+j++S4zpYhxOeIdF2CbJOybE
5UEA7rnTL6eyF8mRUyOGtk5TjugUeNe8DFrALijdC4gndXr9eS3zwTYWrjVD3/7v
nkzczIWvkLAcL1TOpiUxs5nXBkxSWG/ZCAUNZoQ59CxBzwk4Wa/kZBBPOalW6KtJ
H3qxdjNuAlEP73jQAfqqui/fFAL8FqwnuS6imjnFg0GcGYAxsy5XvXPbJKlVhvog
akfg/U2gO5J+QBXsgZZAcTvPDEecbb/NpBGex0bCBnDfFxMFhqeotuhuF8GZ0/xn
5eTp1lQCxbbu3Ql9IRmXbjMTwTYNL1RpiLKWiGIgNv4=
`protect END_PROTECTED
