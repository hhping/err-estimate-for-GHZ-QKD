`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aypJ+SOcGHXz1eLzJOzdzKt28Vu/PEXfOjHZynWbOQcpsCWAGxlhwdDfs8H0uD98
AZ5gmf7+wg9c91JYr2C024kKMyCMJ5MT8AS45PqiMN6lmVrQp9/jEsUs0lqs4MxZ
HD9/TN9ve+TZ2dESZgaP1GhS3ssu5xD3jINSamoijnLfMnZBXI3rzxPF6kK6X110
lmqoGH8TTx1wc9ASPnVrnbKJ70r+3nuGX9aJnYzCcE4z4cX3Dgme64XDUMUN5gEJ
qsibcNLTO67B3I3n/9xDhLK6HeN34E5s/STE009JJlSu+GLR/9YCXnvvEXXjXlzf
pjcMELNEa7fMqM3A0Cb+UTSJ3Xt8jGO7Pue8Ig0OxsvrJk/T8dVccByRhwHm6HmI
NJ1Wkjt1RXEuHBHdr7dlLv6eoewbYMKXRT5AvAhZNhj7/TZBq9kJ+pOjTUFoHDQg
2Hm4coDvQsuqUz6msVMzsMtnKNL98Q+GQdJRhWEz3UOOqv58GD+X/Rm6gtIUwUr6
XvXLbCFXb2ATyaTxLiKHjKycksPHWCeB0xLvhJUEzr28vTCetIz0XKAnkyxZ/FJ2
HZ7nTb1A4eAw0mxNd/GIUKzvXBVQVGnMquW7+lht3f1OgbG33qD4WcJq6bed4NPG
vP1I6f9rYa5f0hSVynN1ZU+0pKxDU3TgN5nhlkDPNyf3r9X6dIphbFhXjFwuwpJc
vIOt2qnYObPK/3wT6S7ZZI8vgf7evXI6sD9RyELvh/7k3/DIo+XXmeQOOVoBhhyw
aInhearzWUTct6f6ZbrocQ==
`protect END_PROTECTED
