`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aF/wkCWexhNC9JsuWN4nafcJkTY4IyxqKWN8Mu2G26bo9DnBSO3RsXxoi9Rs4YGD
XYW77DIxNJWxGIHUFLzBkJ8ht6Vh+fvf3KJUf4NCllBIKzuKUMxlFFOZfVXuwhz+
df5KQhUTyF7cR+thhmRn6Yy5Yco2FWWaLm9nn6xtXyGsRmvt+0keux70lIe1KjFS
0EzyST9BU4WtkFKzFYuTkB1cJ38I0LmUAjakdtnejxWYZuu22tVoGNDhOIVNB6s9
Gq2Y/A7ZI/bpaxJ0yJY4OJg6Dp62Bb3Rli7o33lExj9YldwKMeplxcPOdPcUZHjW
4RebuQDLDvC8lnhFZHxvWAYNBSaRHWUR9mytAKTlXVDZEq7o7qknRUwEjt6PE7cQ
WsXMzYXo1z97Euon0p/EZPxqh6IwkJNEYC4GJXa6XoDPDSuRS9MYTFMTsnBybwgj
kZctvZKOFW/BUt1QJu8WBnPCoMTTZbJFa8OY3pmeU6nFHpVKpBlmLoEZw0lP59uc
Qgz6/E8atGXLkdrwHrgr/9krCQLoBPAahta9TKf8DcaTkBDO8D/NIsvxV1kVP+bS
b5znhKtSLAii/ka9CtsPeW/bXFxOGMfKBs4FQlIabJ2naiJzW8eepk/3I2C7p9fL
xvIbSqoFxr+WKPaicfCe57DM/D09sVOHOxbxZM4SKnjKDFgv264xzEF2Z8y/hcd5
/FCRxy2J3po8nky45lOYx9yrWqG32MX6s5XlSDOhguDMNbWyImHmaQUA6zFa3XwH
BPdpX3EewSl8t9UrpRGmi1Rr7zrV29iVUxmVQiTWFE7GigxoGj6rCPugCSTwog2N
MxJUQvmzxc+Mm+XI6aBx7DcNkB1vDnQfc9X2r9LwGRBiE2IrJY5ayhxu+vv3MPG/
OEyy9+GjLiyyX0MNh1Sn2muMlcfFmyqNwIgNOeYr+UxWO02owYQjarRx/acp2L3l
VoCcJj+ntpI+e0+ETxo+az+pqCv9A+WQ9IQsGzzFRY+RwtcnZMNsEmA5/sIf88jh
urh29bMOndTlOi6lpAOUcsEKHgB6G2BXkN3hwgkkM0qyCTvsdK2DFe/Rfg0mWjNf
k69f8RYF04BG3qe6PriDcg==
`protect END_PROTECTED
