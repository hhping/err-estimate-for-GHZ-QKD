`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsQli83htIvVSUa5YXRQdESbDr8sD44433m9rL2OdnDvtpkj4hcejectboNOn5XE
SKSeEWJN2jZve7A2IoeDuRAJ5C5n/JaBoMKx9lLpjjicrGy4GZ3pNcAW3HSjuoYX
k2Aqhj81WWHxqxUN4F+hOHrwU6pEnOfRjRMD+uy6h01ACS1szMMN8ZU675jhWu5q
f0Z7DsIp335J3C/S9eUUMHSAAnmVwpPJ4bBNotO/356bPvmL7UOIAV5ddpem8nBd
dBNuSx5NxDna5c8khpIXcCHS3AhP0H4SJ/Qditrk7v2sSyzE3nthdZh847IusWr7
LTIKdgB7dggvK0MYEE8IfgFjYnAOCsFynukO7tk2m5MDxuiYtz2nftlR1OTK0Tql
AXB+eFCEy9MJxMIDxqwK8Yo6MBo+tvCoF9eHGSyQvK+CHVYS8gDICy3GPp3S2C6v
4D0/aN30TfW1UKVXdHVfs/Qye4PTek6ASA8YkIn/CKkXG7V5rGQvUYpWDIo6Q22w
/1jDUKViCwUY+kQBTcK3ozb7QSffmNHHtmSBLJH82rfbZjuemOQrHh+nkoqApZ3J
r4ybld1Kp5eFfBoG2pRV6s7wAPgHsQGEQQykWvelDQFP7aE5CMKtNsgUZMh5vj/k
F9OYdPQdvT4tpZNRzyueN9taMevnRpH2kay7/OgvqKjYdEyrpronvQU68ockWjUT
XNRhUUehlvhATpU3mARXi3F+LWwjFGEvo3hOXq18tckatXKptLGEqe2N0Us3ca8/
QGJ04hvcBsN2hhl8qHRMctfz17gTYH4X5avPK4cbQ2tO6zRsx/1q67ACJRzOQc21
zbSAM5si0mEKapiR91jzks6+vglrCIuW1FFiGUkcLYdM4DkgcB+wk6Z61HaBvqSH
G2l70MwlU2nbOkhKOp4z4jX66FpGaV546TNaICvr7G/od8AmClSEB77DkWrIGDL9
BYxkFDxcxX7ceeND0U/T0NdTRGAlM4DNNsBPL4lj15TTSB/AF0dw1V/4ANGMjo32
MiNRiBY1BicmEL/EiQ7lLqyCoFIDqf9OvRBNnBnb/oP4kEWcfHk21OSKgcA7wFKq
FaoPjDP30kzp0t3Eo0TeCp02OeYectErTs7UBXqRcCDUhTyFRCPzGRF8PqRNAV7N
Gpte3Z0lMadqAJx/z7atGo4Ti/W/iaTjuqiDUxrZOIQd/s+VbGRyqyyqmJo50gMq
WdWrOZXnpx5J7/9GM/un38JIqtzMskQYYq6VmkPeLHC0xGDiuQyWtYtn2PXA7VrH
jcJbjEMEkuWEdW6XuAqqG8woEgRl5Wf6PlSldEOdE+PbSAhXZaMyAmDRtGTKm/gJ
Y6cccLFlEPGGhZTmHUliLca2ydD6GYydfGFZ7ykOzXD/VutDfJ84S3WxOxoNC6JR
d/svLtQiAhf1s33181Z9jAdhkvDn4jNcMaWf+MoFEC7/591j8J5Eklspp4viUkya
qGgfjieHjKAwmThN+UAZvK5qqyDThPUpSt+BrToWU8ifQc4UfB1hbZ88ahx7RPRP
POeKD3cbekDtPILjfzpPK+zSC12pwTA/fMlIsaMSP84IftAMxLC7SyOgi8RDo3jl
YFSqExAirnOFxEmXFt4cD4w1zwMi7imQUfJ7YkgynOTkYCAscQDAvgSNcOHhU7Gp
xbvAU7mRDdBCihlml1ZEzBjG9I2pn/TT3NqzU3Ckt6XBX0VNYAdU12lMx/JkyX7u
RmrMYtPVaHtSBY6LU0hJOLES2Xfur8bWvCDl7zKhqfg6+wIKCUNORe1LOXrhjrK0
rH5GgjF2kpAgErLSinbX2XPWLtjLE0CfN+xeJCapXlVRmul+NDPuJyVYj6iksW2p
DCxUo2XL3f+6u9uERHUZ/FYsqmHNDPgwqw7QjYhcNrKrQ3vAjthiaJbRksIQ9//L
04lRMtf/sR0nihpggEBQHNBMxK2aMABKKAMJwn0VunPwd5+AgAQ+woHmA7obAr70
84oj0JT52T9KUUcke0ZaUIT1jhaxKC1OkwsV9X3GmCH/WUKj+6MG//tgMd7Xka/g
lXr18T6eA7pY3+9V9cZzGSgdKjOjKr3fkgYg6vUquYgnkGrfj5xflAoN8SJqugda
OHhXCpA9Fifostqib32QJRNIjJffphPoyjliMsNz0qyoQanRLjdpT7LdZxKCIbBl
bSJV2GLLSGMmhAa96JT5FcrtXfTVqobPka1W2boOmEKRvN0nDN0VXR6xj+f/KErF
HyQ1lD7ppaKuXKs8F3DYiS+B2kbxGtsx2w32q4u0R2pluqj3cTQhsWH/wKZ0MalN
kJrrZpcx7Yne4XLpQIfRjGWBwJ38v+EWFUWKRwwOGbnbLXOiV7Pu+05bP84xSgG2
XKsaUcQQxTx4aI/BXIhOKcu2++oQdu2ep7V/2TfqIyOPMqLjNBrwU9q6s397l8GY
Ta+eJY7Wm1XccBrWAB8K+7NA6/2GPl1bOgo0YFPOVtdD2I3uWWBxRCj2EiCB2WHp
MIjGZj/sZOtEIKAxxW1QUi7cDoA8jRzSm76eVp5HJ1vT550QnL7RGELRWLfIKOMp
NZF+WrIMzB6nUiHfXs/ZfMRQTUIq0mPe/Ae/Hg1PLWuZ2JMktOao3T9QGtlKOOco
yYbXS24RSu7yQBTLP/EK0e3+aaIUPZAm+TR9RF0SGe6PSm/dVZpFoZnHGrA8n9pb
1sAZeDHEo6gTFJWLpwvDqYixkJ7gw71fqnAM2DWBxTxAR4WKo4euSX7sHrG4QRmc
qd/cWKu6yqvCdc8jn4v/+Y/CgThHGSZW+k7XRuVfRu482buEedpW7MpxugQtsxIE
qTXsBv5FKXeCYSxCWgUPvgO+KiLiiosUgBhwsYgbwjjWwXEqgH3rc6toSELynux6
A+Qv0Fw0xdD5wdilCOGuHspjlboqz1l4sQUn4gCzJBp5zXeS8CYFbXZ9WXzf3kuo
5gwB70UR63JtVCk8GM4qhjSiiToCzY5AZ6LhSAE/pN0mkGQl54eQDB3tRWguaEpU
AQ4Z6b9Jtq7S4Jrxk2fhHBFFZzg1nyvgk/dLJEQhIEDeG699WOpZRFGDaYNW8VNS
FmbhV/Dbel0r1ozwYMPcTFUGno49fsatw0urUIZKpPeOjLq2keb0zcZ4CkQ34mGL
HrisEsqTE7Fnh08zL8Yk2NX3ZgosyLXbh/jd1/U5FFckloTgvSUee/858pgbUj5s
4/N9J+GbxPT5V0vrrAYacfwnlaSkGB+GkDJ2nZAaLOT9hxbqb/tyz71xJ2uDYEqZ
dYWx/c6BBJbF8Q2Vt5UoFnSXN6ZhAhxE7Zzn/wyvxPC+RSVTlEi1vpB0xGQ/xbgT
X9XZnxpo3RtJjhINXGzUwo72V1yPsbF/Om+nszpkbM5x9BAzgM+wS12yWtAxAVhk
ekpwVjtXDBNINsoDq5ABDR4jQM/UVEQ2TbpZcpaVBnYojUjG032RMqlhGrblBAXg
bth6B8PUXHKdHTDdl3Swth9XFskU04J/8qlI4mBgpZg12ponodTCfDSokbdhdeKP
7Tk+shLTPR1/IdVuZAZ+LHNDx61uBz93XMsVQV8eVPNoQkIFh1a+1nxOmz0UUbPz
/YkyJIYvxt7Y5TKW/mihCCLC0RGXxTByunPvCvDMPKldJ4CJZYq2+dRJ0+rc8LGa
JQPlsn4eLYo5hWow0qzVzKatHh3vsU9yA7XUaMtDLg/EEhltg1y3SJPFwZILgXQr
zIOiVaoP/hyYg37mKRtiak78xQ+f3Eh0ZsSCRpyqkxkmB1zEbhskHIb03RS3kqLP
O2grzBrml0WRqF/dVswpE26CJNVKty9c/aHusNjKpxqHfD+XMU/K2poiXC19Q3rv
ne0vkQtEAKfypgHwxICw3hYWvldpflZO7uWsDfXvHltJErOhElSlGNCMwUd2ll/a
8nAlHYiqo4YTbMXAcnIC1qi/Ncnd5JTGI3mxLL9CZ7WIgzvCnhMVWINBbiPAcABb
GeO8PstQIYZeW/EdBRh0yoBYsahjCdUFb3Mx+iYXEInHrTWsKovgnnKRr8WyFf/v
sm5sJQGoSm2Fgb9Q2EQk5paxb9fc2nVB9dSi2ojUoU1frvigOHLh01iEQTwe4/HT
mUgsOoZi0YqhXi3kb1tSlsmAbJwFfjhsRIOPftEuWeKk+VxDwi9ix7xuCMQQULpL
zG1YlkxnF3x85mrT4PWyVkjc3LzzFyDO/nYBr38e7FF47k55R9F8QXSPMo4SV+eS
aWuv6uoGXcER5MyoW7PwNcgrbXg5RK86O5gZqrgg1tMAE2+wFiDUewp72PzH0NB1
LDhJ6W+eb8JDatj1nNP8lC2m6m9Csqj+e9rtvt2blmVS1q+l4lYoiSnREXsQUQV1
7i3UsJ7h8fGPG6EpoNZIDzlUBY3TnK3QOWDp7SCZqj8OLmMlCgQGbacG0hmMzLqn
or7Y4MXDT3XhSJGfjz2VVxAD2GfnyOQ+QOdrYQ9QZh9p4ZnAGY23i+MqF8+emznm
J0Z2cZqtfB8N0jnUzIg2ZnES35CBnjbVZUOqjGuv60qfIiIM2SzGwl2h63DuzgQV
ytb1AVZGXsAH7DzEd99wKslcUnyUsRBzDoKOeRDPT5YTcNBhSjgarX4aqjQCZxTh
tzuK4fE1/UX5f0fB2kUHiebMb4NXqceUIaXyr1Tj0c3E78p3C+xnFtGDrz9UsMJe
sGzvgv6740p5DyUoCz+vaDVzDhRgWFJ6iHTPav4kSHy/X4b815rcdgIBR8unxBuW
5KSrYm5xcKsPTAB+EB6gyTGMyC/xqZfYe2Llgl9tDb99FCIliFse4Xsh7TMu+iy4
ZHk+RQzlgLXGZTY0r7LXzSeD7BOCEMjm8BuCYuizOfCBv6LTts/RwakWgWQkVnXg
qDDgwiU9cSLf/ybUOvEJNXyXko3fRQzJaTDbIAqdtJpz5p/gIlloOf+GvtTTQ5rS
X/lI+5Lp4nTYYbI1IX0b8xhZ8iD6hwqFdmm6r6QYzqyuOtMFbQtS3mKGPCFh/t8M
2LcO+qiKl5ds9VzvytCr2mb37vjZPswYug6R+7xZKK6xEgTSQgM7LAflrRFqvXfu
4ta2XBlFL1jInYRumBKkxm/8DVz6fmJpreS6+oPDlj7LhuCn1e4JpbohN1frl6f9
l2bXMQfabpbSgNdHBnp8Y+s+N8RhhaFcKbKYb9I5x8V/ruW+0oWd/4rFo8RbTLCT
2WSvnfluv5Ojt8k35vTJ+Z6dkApBQij8hCmMTwntvmRG1pQLbBIGPeLnLFKz6zs2
SZWNhbwkGRUUtmR/ajRys1elgoy4UY1/zN+FmfqLF+wGhXrBtbUMZmDBfm/hhMUn
YvMW7w2kEB+Wx8kud5Px2YGH4xWcPlh9yWSemtKeYQSwRKWG78FzsUUblQAKTY6t
wkJWiAC0BfVJG+qSVCQ6IlSeMJVYJVSnVHVRoI7gc72nNmLzUlXQX14AxYeacVIr
ZGin9rPEAXRafUJLu0KZa3p8UhS/d/1g4zfawZKdmXmeM7jSpUaLc6PaGgd6ruvu
w9rBU2ifk7GxwRGT7+QVpkBthOXt2HZRcoSM6vSWJQi2vXVz55fEiouuLbTj39GP
B7TIX8jxU9tPy12oUXHgellwHskuARhYJ4VRHEZaRfF/lGHihQqU7y9cZlBZJezv
A4jwxJB5pDFwKWjNR2GGZQAuhnoS0KCBUOZB+Rz9olX1S27eySdKFjLF9anG1XLn
AZbP3iZp1dnTgK1cqzfowJy+sOLtMgnTFXxnUm3sgwn+rKSbG7lVwbsOcorrtJLf
prgaLsyvO+MyThdtHIJdf/lnC0i3If38NN6iNcximTYWxG56aKx6SKSqrT/otZTX
TDPtcvuFSKQxDkVrMWiZbMJuYW5Z7EWxzjmfaMKTH/C3nHJrnm6vh3GgkQnThZ1p
slzqASXvj0/Ng0prtCPMQEIrtixX+tiCl93G9+1fLNB+xngoxAajmU392ZX/Tqw6
3qcSEVub/dYDu8e9g6oUGEsLMgtMP+1UMzj5T/a/YGNBeSQoqLHJjxW2S4vVIk1R
U6rrYhMNtDeohKXEeGP0dhv2/sIUcnJMrO6aY8XrzFebxxUe3rL/P8tuDhjnX8h8
oVjx5gLfr5zOc6tWOKt243wAn79qQZzbDTH+vOKlHXn/5uveyz2bODTWJ552Od3H
+3WKSgUmnAT8StWpCC0q9yp04GYI7p2Zw3cdkf9emfWir0qa2GxE6V95HQK/JApD
Nx0obvLfMw5SCl3daISKjiftHfGVW4lC2/61icmzx4wg/jPwSzaJ8/t42h1GQ8M2
OtHkgdWr+nARf/9Z9PABMJlRNTyr5f0naaIJME7GO0TwLlCKvIi76oqxbzcsn6zJ
dy62YxBCmE92+vx7gAwAsCR2NqjtP2cs/j1Yw/LCGGu7P2vfA5xVsYHzEv8zwmCf
mXOHavRhCaROA9+LI5lGtMMP6Yc6R2G0KamAV3e27BNRqiPVlEhMWEkIIRBl521c
H+nOwoK7TeNTPq073uz42YfKFVDJBsePu0tROmYzZnD180Guv3zQHU1SF7YmNY4d
AzjxQ5zu0nhcmXB06F0DaZtZ5WSMdtBmYFIArQXD+VtU9Y/u+EhWgpMRUN4gFTEM
cjFqrjv9FdpYAXXPAyVKSLf9ptMAOg9qqGY6/+wXA4TVLDKs93TgQjkfLinlCaK8
t/hlf7/qF0W4PDd2/yLE4oVEPbs1n6fLiCjgWg/GWt/j7Saq8pvveubufiJKSgpK
CgG2PSjJ94swJ4fB29T2emI+GdW9gs0Hhh5NbxSPDnfgMQAiOBE5CuCQ3dM7QaF9
8E2L7frTe/1sorijV7LB3Qiv4ftTh2d214pneMb2Wa4t0VCIYyv9JPAmeRAJEylB
DD0fZE9He/5XHVVSysE6RteJo3bvZ5n/IJzgZvFtsMyLkDgCLDSm1dob/qiRA2+G
G0A/UnSc1xTPp0tiopefzrtwnHN8t+Bn8M0DOTbdWZT0FsxgePShcJAMA35sc/2T
iXRFTwtnYUMMArJgtwixofUeORr0clXtJuVnod8HBTN7YkOyQEDmU6nLxgA+kVqm
mAZTn4/r2Cvd1EI8J86varDPiwnZ92RExwW0mwpfNN26AfTOxaDgoS57LUK9MVOL
P4yh1bPrJyGnxAsMZ4DND87zJcy3YU5UG10IfLM0Tcw9CcQfxZTHgI/Wsjn+9aLo
h0dg5NVuajYwZzeswU/Jiw/mSw/W0hpHvZEUpiZKVqYLYlxgxw4UPEJ8QywnRvP/
sBHVUCuf9GP1slEd275yWBa05jZTMkjO2gcoLenJa4yAArIAmIdy1JPwX+vNyUvA
6R6b8mu5xatpl3EbiIIBcKtYjuCuUjwzq9CFOZ7a52oHF0ZW+27ixy9AQRFicLr8
Yj1ST5DGSc7K09X0NEoMC7Xl7YZz8C41mtfyu10k3pR3ptVYIORK3FMkPuOVBnSM
QBChR+OCadWpNkIVK0efahSMK4GnOVTdUo80LFAcX8IcdI12p9nsKYlt4M9VEtst
tcAlWRDFXiVpXGCBdWhP58YU/konc3M84GlKqmh04hMp3Vw0DMxOErTS2mQ0Oa1Y
wQcvozvaR5589TgkthbyIpaTARlEY0/GH3/YshMuJKiJsFZwfjn0yCn/siMx7sx/
M8m08sxWXk9YdG2IQudrdS96qkmz4OH4Gp2HwaflQwWAA3PD0HMPBAFP3HvPbzfj
AWntF8e/R6iTOvQiYOeB/BsrEmOozLWBpfWiIegYAEZ9DxbID18ODiqwTtMBusLc
4+14HGkpuh4X2SatZbPqJ3N1R/SIZIbL7lYECyT+c2g1mMP97TEBH87EJv807kvE
bA1oTIehfMjuRU/WfP+qPlr5RS5ciW6UdKjT74SXex/+pZqrl7UveVUGbeaBaG3Y
xHWCHPSj+n5Vfd62MF8Z9LMm99FFf8cAul6w+bm0CguwzJEHGAtyMPPWLCRJsAqH
DwO+7BQM/cfbLKCwUoQcCuEnBW9siO0MKk3mQioDehehT9f7PThwlz8aOqlvj48S
+pEtfO6ct/aH8+EhnJexG3ZHwue0jYxacACnJHFbN9bBuJ687cmPmElTZb1YxIif
Ua8gJ3Bl2m92ZEeGMkAPbZ1j2Ben2WfoOW4vFLajRMIvGVJSdbHc8j7Yxeej1fhV
mlF80ch2M79+cWCKLSnCKAhRPEMy6RDwK/R1EcQaEjoNvtYs0BTAspg3qmISbFxy
NZv4Boxx6dClWC0YRPiEnY5uW+/fQEsBfw57LUA0RpM=
`protect END_PROTECTED
