`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzRZ1YRx+Kk+7uZZHF86D9biYSR1ZT3l315P6Qq1JE9BeiZ4GFl92qsnRLvWBVbK
haXqgOBuIqcDoD1chma1Ela4ClEnJju6lfq7ib1kX1oXB0hOApknepSbuwI2ltyI
tqnbbr451mM78Wd4m3EH5g1i/PE/zkXfr8PO2I1e6ePtQRBVuPK1bublRY1+/lpW
ytHv66eCy5G+IQfBVl9lbZ+zhxyW5wDR537CT1OObg0ZVyaYwHbE99r8098gK7Qn
VKU8aZfm7Bna6EU7vCwsx4JPvzJyoAhnMJR0f47058k39tPm7MYRgDEDqaZ2NKch
KqVDQQvYKOV8jj+tyWVWSfofq/z6UGpFtN4A3nw9kK3N4PmBoN2ELtax7LbQcbFT
AiNumoLI4b5AdCAETy6xePfYcxH/JFMR3mcKMsj3JWOzN+y4jV5hdwx9MCdzuqI0
zASCkz3NRoESZUHLfpUg6sdt+faV1n6kBkstZ0M3LoyJGK3diyejnSnlZR4rkzH6
UfJrR7NRVKjbq2YSuizY3iA1BK9FBRGrGoWcwaUOHx2umUHasUke9uFcFuS8Jitc
Js6B0xf84lYggA5XcTgK602CNOwHpe1moDn6/S57eZ4DpanqfrbOTPOhtT+y7Hzj
Wdd348fJ0Cw22CbEuhQ9Bv9WOQW0+g6mJS4UpCHswbGX4+HY+L42XOxQiFOBczPQ
9fGcUhA58X2/VvWuPzQfWpBc2g0si8IkiutzsZ/UdtuG+UDuhY+eBDVfmiX9Xrej
ZpNJ4K3qlXPJQBea7qo++neSBujaGGs5fYAr5qJoG4FUmGwNYoN3hK65pSFqgBnP
qRK3m828xqDypUikBzvwnU+b+ytguchqOGZ6q1GofjaxSiQ8jltpAuBGCPXjO3Di
qlytYewJnztDHdOOPatARlcbrEd27HvDuavNWmymPKKPyAL3/rEIY4nVlwJjgzj/
m6v81v2vkpYkFGRfImKfdOCPtgglaSMr0mZRlY6U3l80D8L2RtzZEOSs2F3S8zpi
NmeE4tJJmKN2Zr75OquycnEanJjYsAuvRqQLDg7m3Lgm7Zf51MYwcaA2+lfANdbs
SwO0MyFISk98zKSXhpqTNVoKiWLDRqwFXZ3TXAHniFSkyjUyLS2ImfT8nA/68+R2
RPjSmY8N517aDu2UHkzr/Oj1/BYdqXn3TL7G41MPuxytiym4Ebqbm7mVQlObR5Im
fvcoOZb+HTO0U7/w2vhw4aUkGFc1F2hYQcAGkMABhZbMZD3xhQfXHsK+DcshDyoX
Y91mu21OGN6xru4BTGtaw/X7F4GvEtVLECZY2bEGWWPOhSDR0/R6TXq/E3++l5AN
0Bne2mjfqwdIMPRanohx3bx+BVxgA70sxq4wDzcmp8kAUnHIZ3wdscn+oSNE3WCq
xjW8AJ2Xq88tWzuag9OL2GWizOFzDSjSfqFcojq1luPzF6QHCU5j8k1VzRS0KwSS
+l3NR2sQhKQKLUWgM0bzI44SfJu22FuwQqgEC0ilx+NhFGX7BmI2c6AjzR7KKU5g
IwbrvHbWfPMeyEhK3ydB3fQ/otlLZUpL/aJGJujpSNqQB2dWH0iNroT6wxCEfjY6
Kq09OAjEU+yYHekAVYESlCXq6sXQAZuXtfHKu1fgOc9Cu1Ip5Tj6oruy38ICWYm4
yatRSpccqc4COdeajlWGFF/Ohg5mT9/ATaX4IbAm9S0Yi4nWCYDDQqXigdShL9ja
lcT/we7RGTm5klUv/dCzM8cSEwtADcrRjg3kiIwl0PYcdoVbZjL6Yfzz8ctPLChE
WW6Mip8H+svk5jaR5I4pp6Ef+eyacOxre/yZPzJUAlnDhoGRQxGaIAwMu7MOrNto
Rdpw0AUSqYyiRaL0NpJ105ZEj8+G10wLeSVVpEB7GR4l4ICaaDP8Q1eRNb6lcGIV
Ob3bGqMHfIiSCK7SVWEks9ivTCUyQhDrVI6q9md9N9b6YofmhB7wc4DFdzeVQUl6
FmBcJB2J9ZM0etYyy7Tz4sV70QUQtBGbT3m7vH6XGT57U5eJUS97nDUqJOT+Z2ID
YvK97F4UHK/cO4uwNMdRqb+aPgUurWxlxx5xcdceQCJoydXR8J+gQswTAr9xr+uZ
V2mK9sT9k13a4JBlJNsr5FKvergR4oE4B19nCAIHZkos02izLKxbNtrXuNoYgiGO
lVvjsBv4BOwo9XtJgjcqdj5HXJAgUuHhDfPglSalKmYr4LZR3DXhtgvmmf6ZSvc6
Dl19EDAZ5fvOyigWetD64wAofDhwnC89Jq2i0LHo+PWUFM5EA7NbIqnUl2erPBh0
Nw4k/OrWrhBGM+iJf3N5LfD1aKr566IofgagtzmaVhbQNr/LvmYN6WvGWtAKjm9B
hNejufePkLO3+yf83LIB0NW1G2iiLfkqmQ0/OXtiFQ0=
`protect END_PROTECTED
