`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d3CIza+pzTBSg6SFvZxbyzZ69PviwFWydGi2+9Xq+bmqj9Bu9oFCZpcoGvNELeRR
0LutiA5DfadLnEV7Ew1YonlRSM+/ONmWvDz92U+Fglhdh6F1z2gMVX/VUWDWTEtn
+YDf4QwbDXFloecN0ZBVC3TZem6qYxXzDU6mVK7voynZ1bKlJj3jrBUnSJRrnDt6
yP0RF9C0j3GP56OB8ZdytZGmvI3KjvXvzdlrwJfDWV2LGyvWV9V46NUnlpCKrHHj
OzTQCnLdY6OnEE382H4VkQeEZHwnHWVfHCBPpeKteTzkOZGLnNueMW3AC/BQn3jG
L1jO5vEC6EaYU9/bdnjjQAf6ARMPzG3Vd3VWK4TK/Ay7We8BoFD8vDndT+mwwQuV
1s7y7VvOA5A6llIQhZtSitT0Af+J7ya3bbxh4/8tlz4/ft0fZF6MNC++mmeSPtX8
MDUAv75qc8QhZE7tB2YSuPmiufAx6eOI9q2LoApZxwKeg8Dec+f1MCoQ+XVuh4+V
S0wPfSTkp6WvydFmFeLB/1v3Ws9VVMkSIqTyK4X0t6yeFzT11/qJKHUbRbNJ1noe
jbgFT0/5/rvqjvhR83TcGLpJKT0QquQ5dSIGJJSTLZu1WOijfqktxs1RLtBcEpke
zSOoBZjaIlFSDJx64bBfys8KlUlso3HA1O69g+oPKjaGbIR276hyxvyHHRanq1S5
wF0ADrTywZJbPAB2rioTLSQIU/dq+6dwzL0Dnjo0RXYBGvfVr0Qv/N1buf8Z0IOb
Abgvbi0zPqp1w559rMGzfcvjnqjJ5M30a6sSxpSe2Ut7XMzSx5MVZfYRBuaWIXc/
1E3QStNZCfVUc52quuyjDyzza2hRpWQlAGdqpqarmzDLfJkZjWANUisj8W1sfRar
iU5nT0bMkX1Pj8/d8Tvp/muTHiKTcHlKe5BDuJLFwcli9vO+SCZza7nJGgCDeGH0
Sy5cmV/scEnNdLOyr3+ZC5ofIZ+oUSCNoqvs1GWIoIlNuakHqw3V2cdJY22Rojd8
80+O7ruZ8cEryBeq7cVmcY2yi9vMKr/GwBpK5FYe1PVS+6R7FruMKj0Nh0dzY96G
PZB+7qWdXod59SLaD516Smr07uI/0oiJUDJjaQhH3Qm17A6xIg6J1N6SxlUzPjQx
JgLaouUYblAbrEoiTxgFaGS8IgWB4g0OjTKEFzrZc5iomilYiA8F0Mp9oBWNFZ0x
R0BEhwd6aSQ+LnWRUpaJkUWhej8lzhJvDRpf5OD3oj0WIPn9/W81TtBJlwKfqkjB
+rqJix1i+6cn1GJKJrK9DQFhqXX1C6+d7ifNJYG+y1z3mxsGTffHKPkromIvCdgZ
ajD0Xp2Rw/IjlbvM9N6WQ38FEYNib0rfL0yHN6J98oKg9XCCCKaHAUIO4TEZdjoa
g2pPEdRP6EnUGJf8KeVWGQdWuBndUO1WMV5FPIBtmeBcGu9+UIGlzmsn0zkbInFn
VzJ9mgTdNfCPztq6Ws7mvECs5aiY9HUg5lHaRITpak78uTuRwisCg6ZvDmdvcRra
`protect END_PROTECTED
