`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5ptuvx7lSegLG6yrRTEHhLRZksbnktixB6RG93Fl6FksOVBjPzZvgZCK7vMDgeh
bnofTQfUX6Ki2JdDb7F3qDiVS6paLw/YWuSGw61RPQ0aJyZFbGXfqniLxV3AbKDS
dgqFBQolwQAhnV9g2094vR6R9z3Bc/gK23B3YREzoeLWjaeXTI59nx+eIaDqBX0l
CUfv+kTy+JdsRnhqvJb9IPjxvyz1PZTrX9my/rVytJyZXonQ+BgVnH8Btaqe0Q99
CYXg/heoSPmPjCylXjjxfeIH169epvsQEaVfW/KaVt72ifh1CUSXtLriQiKr67eX
NppCUlSyIU0UfZkvWiccLBq2Io0TzI7ljdVAkmOG/V3CAqbDVPOcCGWTgpq2tcxg
cxc/kUpoJRTgrU29t+mHmc03SdH9QwQgQp2/BeWz827TfCguP71UkBtAyHxsK+AK
ejIrWv9MUeuG8Ybvd116PcGGYVe6VWy97rX6zPvgkOJ6BO7awYOaQhHM8gLwRfXw
M4XoiY3mR/RgeA/i1uCz1Nwch+nPX5APN9xWHw/uTUccPRLkMCSWx//oTT0qDF4V
2l/ALHoWda8Lv0W86hOqwuQ0VRTie5Cgw5rZ99MZB/+8KL1/9e0kWulauBgM2h+d
Lf2I3bTfgBxwh3VWNKY7Q8TRU2SrCrTrTlncR/7ZT/TdhDNBwz1yE3uH2Wm65PaQ
o4bt4zF7Jyr+vfNrb3NImGouyLkRMG8ynCehrst7Hx1OCFOw4myBTjvlXZU1mnkf
ayzukTkBVzk6Aw7v1NmGQqSXVrVP6SzjvCp5DL96/twQlgq8e7SGpeTkLa5MelTu
uYIQtafnQm9ysbT/1y+cCd/N30cd4iIyTGXBlGnFgnnsq00o694gacemUVaOL/tn
bgXgrSx+Bb7RbwxWvZVwjGynxM4NpOvoOXN3MqtNCUa8FMLNIiPPVH25uCc8tpAO
tRF9bSxRQpsx1WKJqfV5VdIZh+jS4uscq8eu2XjRaSJdBwnD1BLfyUndfYFMiP3C
1edKNO2TqhCcCTK1L3OWqc6QF+W7ajqksQE5Gq4G+Ki8KBGbXb6eUW6DUTvq5mxn
ncfXGpHG9rLIw0HzEJ5IaGkke0A/u0bIb2+MsFPKabo5qkyKOxhogznVxn0KSixh
SH8VJ3em9mRNTQeD9EF3k7vX0F4KCt0438oZj4LWDczYtAxA2SvpQptmVyoNppjJ
kXnkTWhAEslg/ZumxrtvQNGQqn7KSp9PwTh1Y7f7WFJjxN2HtYtGSEmGu3+g6zMw
v42+qnsLu28IM7Hp9u3NRzd9Q5b+aFwNtZc9IJI0//QoMYzfAqdXFXd+44GkI7X5
qcvD5+PDMjgVPRzHXUjr4wrzaxjo47NZzgc6LLj+2Ev6MOFzAK0qdAMOHjhkeyi1
hXt31MHBW1F61eFWPeA/D8kK0gx2ZEnYHhDrCtJGlvpNuKPAKah5TyFIW9kz3Brg
SrdqmU9zs+wlD+Rzm13gwC4e1OiVjnit4c+JCH3IKhoRyqvVJnMJeW3jeT4G+T7+
LGdK3UUcaJDYK+nKkE1TU0p/E3s22CWKclwoePxUTzZB/Z86hA63jKtm+qFqiQbb
IbhAu1m59F9GEyEBD6IwliLJSWC/LFqg02DsWMHqvwDJsPyPGEVFNW/Ia9Kch321
MDajFRB5pLS/M6TX3TbJKbploRU2ncTQOat2uMJBtSgyocHQ2HzsPseyFuWwwhMx
x1xoazXM5esGHEau1nkveq7dYbtoEckaPF4q3WJiol079g5uErxO+HzpfPBsP8N3
8q3J75iz5LlWP6F+6NJE7XGh2/048gSH/p1iQfqM4vwQDaZv4ia1aL8GGF2Po7UH
QQmahABkz5+o4gYqKpqOWMHd7GDO3VmlyqCCd7yGohQPNGRT1JavnbooIAiDVgJB
Mkv2jlcLFaiTalOcGn4El0LixcUGXOUNLa9R8pw5lTpTWwsSkek4+s3Ui3ZnZOrH
IzoUlL5XE0TJBwp5BMnfCGAWtBxgEMP4OX7wXV+vlmuTRwBYjC2BbH0lCiaSHckK
HbWbFcZWtCmxa2LDz+0eY4TI6rsZc0PfMirjZ32O5C7rsCkY6ww4T5x32UL5wVPd
cMauf7j2AnYlPVjtq8ca96aNwpIwigGv833s6VmqLP5qIPchFDXwnEDDbjzOr5/O
nRoGAAqNKUCyUFdIBgru3A==
`protect END_PROTECTED
