`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPIg+77rNPhCm2IkEY6nHA4V/8AS3IW0sZktXC0BgSxRM/cFbSHRRkJzaOHDyTZQ
HFU1wbdS5b2iep7Qc2z0cJiAHmAMKVPOCxpZ6SzfhiilyQW7kvnBt0vj6iIsBVOM
NP6pPoxBQOPvkDb82CJFkfdpIE9Y1s50cMrQ4sLCvcED0xdxtg9bRlutCkv2msL4
VBwv3IXyL3qVIJDgciXOczV6zvPYwhAiiOfMAiUNw2ArosOos4yAlqi0tu3tnA9Q
3ljJlcMmB5Q4ySmvk2CFzMgS9vWi0gGmCF+LkI5jkrzrbpbSGNbjfcBLvph2Eu3g
eiFjDxEFJ1RH/aFnKI0DSy2b0s/2hTc46SElOIA9GEX0BIKzDcGfzLJnADlr+svF
dcE702ycCqQKOp9TdHXj4UolSlTLdCHWjhhyWhci6oWPk6AB/5x+XJ0bdA43VTbw
9ADvvePnvRmes8LKKQe+wQUG7ZkhMTTIdGJIVezErnmA4VZwUy/OIecjFc8zW4Lh
rM0hmDFDwCmJ6OxR5mtPgWJUTxcbAHi2UWsGwlLq59Pb8bASJVxx1UfxfraVsY3u
TBD1D0ubyxnJzua7UzR7uhEC4yFEvM7JpAX4s40Ola+zEtGgCYhYXJL1d/83Nhx2
M4fszJcwyhiuuoszNzcvsnaXQWckuktvcVtDt98m28ZkwWhUg97Aia4lw9ElX1TU
H0eN2m++EQL/qwprm/M7zBJohAbTH1yLkGO3iD+Sn+kliEr2VSThCbFyGKh8hdrS
eiv0Cbb4hfOVA8UF1Dcx6EORgtkQzcKVQOix2MLi9BbvKrsA8OZoqTG/d1i20hnU
hnCk9vChdU4Jp3Y9KjQsZ22xTb0xVVwvxn1SZneo8cWXzE9O+VHdHQj7I+/ndsPD
JQ52UeX1zJyhXHmpBc/eE+jB3C9MKszAxaSLsTIim4ZEEVxY0V0VD/oxNWE6Dd8M
8rznwNQE/iBj5ooCPC7Uim+qKHcp4ybfoINe0fQyc8wUVFXlv9os2l+5tFUUWxPO
qKqjhCoDb5T4J41k3BhNxm5vWd9kWt3CwU3igRmXGVTZpxjtEaLCU1zaZND0pjyG
vwI6JtlQWKh+CoIMRkJ+7BoD56+4IaJH3CWEuQSGXfiV6VOKQ91dN3b7p7MBz2Ea
RMYh3o9R8j8j50Oml+48GdEkNozj97JNjDT72g2c/Ev3xocReN27pmzk4+b+y39t
cOlT+mzIV16gG7CFMUFJ44RKiyBXODgiMY9Hhzn89W1w/KQ9SuR/sc3eu1TEgiNv
Tdk6ghJ9bFP/IN0mxitmfANz3zkY7Zw0Ay93PU26ljtRHdk7FCQBbLwXl6LSZsWI
83axGN3ERc/rIeFnNj/EqBtPUOJDGhCJZqo+ElzxleO0J06bfRRx9tL6seCV1JPU
AmtfUmIM/8uehqtZghsJXy/UtXPbjfUCMppY3FYKSGpa/9hAdzSinWXO0xS2LnH2
cArzIrwCSqJkHmMFpvtzALC8Sqjl5xHhXlOGQ2GloKYqKWmG9bQUAnpPEVl1uhGV
0FyOtP4n/8RdPHGgm5pj9/apvVoTAqA6hbju/VbWtABKohUx7aja0RI4L8ie5eMF
cRbUO2N67v2bc/Ma7nyH0TsNXLAzvUqRY212jjHIRfWXfhDl70Bl7awuDzCVEWQV
0A0KpKbQoe1B6/jCEiSXhOTJY2KoyHc/UwA2r+FjvniHSX+DH0KeMYvm+SKOBZfd
EXf6MWfQfEOL92LyD3yJUPewvy/RSiETixa1BBg1hCsuZic5m21czz+jd9FcWDxn
76DbUb7kPm+iYlBkbtglo8qz1utWxOF/MaAxRgQ7MXoISGPyW84dQUPGMNvUCh9/
DULMcWmGhFBzRsb8Fm0fDtYDPSYh0j17XzxuioVLMJxHYPWowoNB5mgVQulpWBOD
wcXbOomEi/DwwhrovvwXBzscFBUnvl6SkQxzJaIFFz5f023UrsIWHSbBgpPPPlJO
LaKaIOtkZZxtQvdzQwQg27MBTwDvuLL4SwgmZNnH47KgYGEChFcKX4J4kRK6WZdA
/Ew3Ij+yhHvh28N75n14dTbApsZ4O3+GPouamiUQJ3CmugcOK/bauRpFpVH55a6a
ItX6yv+3nWStr6Tu3fUzgawaKjviMQIMgIGKp2U+Zk4UqMBDM4MXP5nYRPiiAZ6m
0CE9xMIaE96ZMHwa7Bi7iiQRWIdDwClIwDACFJ+GrAoLHMW8sO4IdruWPcDIOUjJ
va8xFswA5TLpQZzrzZjkN4JBuWf/u4D9crjwJfAxfLFfikHw1gDoE6CuI24dgOEC
yEtPkJTlXq+aTzWuOR7BI9bxexzPO2B00NF5XAXATgC5FDhRtJzMlOqeba4+8qAV
Xs+UTJfeBH5umdlGNRvJ5CiYjsJhbCeAGFo8Edr/yvewN4zMBuCmLh9uHeLuM4YP
WmaqQvF5fpz9ML88dEEjET2NMHm7yCDfcvRDTLOl5obsSS6bu6gsmccySpiN1DyB
c20OqfcRL/YNuYIpLWAVKnT0o5zTUiEHxcB4uIIUcU7/XL+zDtCzhBYCMUPUDXvM
i8/V8Ch2xBR2EZJwQFqjyBy4H1yNxP8kCY5J1jFbJHBbX7ngXG6aKx4R7qycWoN/
zWSGBrXqNRHWs6MB0R2LTvJYeLelZI5JRIgKuAWXhbT2a+724jw48l7YZBndH/0J
7icKDdGnWWs/jtvPaWNuWMf6lY+BikvESpD+KBaN1ngoZQd2ytJscEuk1l6oY87l
yT039rkG4KzaiyCb2InldwLYZJfHg0bs0cDSFJgUDwFqIWl3Ij8J66ej9TzK8rJ2
UxgTOnGjlCviZhLD/fOS/yC4qx2ODL0MMV0z0jvDldtTnbH6krurdivBq38rrXJm
b0Sfg1p3Qs+z8jVSGXYVBieeftTvdvgOUK8JIHKp1O0AWfPjW5h3TeOM+jX9sgDE
eYDAD8uEW171gaiHEqKWMTAesKc1fE4AFRL3TczRbqzP+2yauGV+7E1syeCQs/AP
d68nNthJ7lM0Hb1vpNgLyHcSRTwIrpzDmmeSQP6rLS4je8opVkeBW+QNs9a3EevZ
fR5UxM+fTW6FfDyoFg/o0vlL3/IO9aWGUYuHOj5Q8zzlQg8EejGoHt8u73DblfBP
kpdaf3lcRoTmWPBR78hadZLZFzFSXiNAuyisVEpECAvy8ZD6KMksKdpdQ9u3gR5r
RnIzf630vpiPKL6r/nZ2aSRQsfuuHjL1Io1puOA3i5oqmTg4Rku4QgiBaUIZkNyv
cKhemYGrYo+pMD8qQM0n4sl9sMEdfnwCgLMOHaEHwnZjQOFneCXBp/iXVWgvgvz6
gcEPTnOHTs7GwmvUOsig1/OV4ZBMkZerfF3Dxd5c4RdGf3tNpMqln8FTu8gfdSvd
GgFEfMNxHYqTcSAU53WGGfgn+BdVMG2iScyY4YMP8yS0NcBV2IW3yXJDn/IZk7qm
ZxRDi9afpNUlZ7RwGP6/y3eRiGmxjGrRTKydpfJDC8s4tV1VEdVi8zDN22joqKDG
f/vvCklfJ5zCXldaB2EQk6qFkHEqb8E8zxXDepy8ymo/ZMk24LwgemptSSNRj29U
/mP5eseIweqjNCBGndnSxa4bLVwrNMSn1zfCUTzs10aQUVo3tuIxJepIjEJGF01Y
wEORf/CBjd6lkTssoSi74WXzpL4juVlrP4jvhe6vZ/cWHGgLw9qIx7F/kWDMa5NX
+X0kGwkZU2vClNdz+hVre+E4Gbg9GLxqvCM8+ANoMCpC9FLXIuvvVjEj8JaBl/il
JA+GZiYsndO/Azs+X9r2oTf3cp38V4wipwW9xTqZKf4yGKn622ioVbWVSuRPrrQh
gp9joym0bNZ9hBzcaJKPbL27KN9vEGI9UdJJBlzJdPK9RX0Nj8m9Nd2ftzicbHSB
t/1S+A+yfN7tPVjzLuG9Gac8nKa2lUwpi9TNanKgkt2+GWsJnQJ4qloIZIHqD3uu
8+ZhPRsKXodSJauv4fSvZhauwoNBk5HNcP79Alpmnb2RzKukkpG4ikcDDwJNILPk
niyftQoKHZUQAuN9rGGfsK0dlQd7h6qEbJmuKNWlT5YwYZJF/dhSIgLBE/+5ucHb
KLXjmNPsJ7rUp+aMK/tyFUWRL6GyYvV+cBpTiRYDyEX5lIHwEK0fjdgnruYlMCEC
yHjDXGBeC+JDknF868Ygy4yL9KPBfz0RHb8SAr1CTvOzEjmnphQsBbbFeuzkFP5W
G2TDKjzg/f+e0PIAVC9xPoSwrMaiiEXX3UOngOjlUENGWwC1ADDGkgW+++KyGj+1
Y3CesKXnDQFN8J5VcsSAuOI9ssyMvwrFBVPVUSXiFLCK/jU1Q+aPnR1g2fQA7Ldq
NKBxpJzAWPf1CSFeEaOHusHCYaafhwVNI+UPZzS5l4i9vqDkT6MUpRj1s12mWd0F
YnjfhrUit3URKICUAg/iQ097vy4pDBRj0kkTUSEOBKamkcHpv3FD9aPA8zEoiKdO
yKyzsyWogvhlrWH/uet/3x69+UxthGLtP62M2ANGyfYJ48dwZR0pDIDwHaFa03Dx
eBSLhTqmibLG2/QA1Y1S00CioycmTsLWy5l3WKGDMxdyobySwAW3ekXg4FWhF/kK
xNyfsFhY70mc46clSa+1uvVGVoM+M84kCTa/BbvMkiGTstJaZ1XRUZ6PfdxP0wF5
ntV2x3BQts0M/m3P2IISfplp5+Zgp+rxPDpZZTSJFqd2BtryWMn0LuE6dKa/ETfu
LWNcHqJThmWIqi97ygnkG7kAu5PhaFgGjdgypJan9VqZwFn0OVzr0ACY4iztc+in
8VBwthD0ZGYi8khNlb7j3DmXPOz7EUHusz01xg0utBe/4vqR06LdaFwRLFrUzaNm
mczpIQwy8blyJGgJKiiO4XKxtjIG/K3mTVRh5eBoOX4+Sm1uRFhGfZVQdUT2gA/R
mqqESW7byc4AiSuqKbIplkhXfAc2ZL+KE23ylDJEkWDhdPP3NP7QxsLOxTKzn9z9
zh6j21S34vpzgZ7g9BjzSSThF1ZBamyouznkooAUri4RCpXXNmKFST7ZFhXjTtfc
1Aa7FhEF0YfDKUbMs+m0ZhRkpQYK+FOVSckRCogdJVRzOV9l9M8vdrnxAu4i/2Gf
YOSlL7cbFHLOOPQHkegH8PNihVJzjtLBKg624zIaI8P5gt7b5MWo+u0t3L3LmIV2
jXCNRXKWvWDok5NHxKiggM1P/ayqCBX6gprSLyBiZ9ZFdiTm1A/csLb6vcPueJmr
Ksb3Ge20ULHUqJ5aH/NePESmoMbeFgawLgKowNuCBHPpGZHRygKQYvM2kg6V+IwV
S4mrbLJ03ikcvto13PY8DYehHFxdENFkuTon7xUMPwY1UVT2+h3EvaqK8UEBnTfN
TcA0noz0ACTqAG7W3eig9ItCsrg1jTmmjalvN+gpS+rfhpZ/NxshYQDzJ9aZgNWi
FEd+lsss8exa+RjrFDUV/eD7K3TddRhdKIb6SS0NknX9hfbY7MSSjal9RP3ITZq+
qRjLo7gDNULInzwAvQCOe2gnP4d3jcTKl79bjeDxdvuKA45v658IktbeJ1wqV465
Cjb6oBtAY1S0Y1VaNsKCTK02iufDoyU585GwXZyHllq/VtR2jn3uz65RDLwohXWT
p4da6ZYv35Ht8wH4/feGSt1ImxGXJ2eLzvLKWEoDyfbaDqiUDa6QKuonR9CFSJbT
Ht+ntSPvB17kqc+qGEawBy4THA7DZDdEyG+j05PJxeU85kh+5MEIywu2ocA1Hgg2
VpfowL2uHsGcurpajzRwHgQy4sUI/+tALvZi8E9uwXCQ00OQpJ1mSRdNGx441GL5
ie+VjRK9KFYESpIJDyIkA92jDvpHaMDV/5ErLXmQqnxLFNye9BwcXM1hcbq3QK/e
OZjc7h8M2Jnf22okob/YHEgbVRol3iq1sT0Ec6IhYcmXuKsg2+AFUQ3Ia4fvyv02
/WajUUmYvCSZbik18R4fBnQ2EdWHCxqCfrJaD2B8QNd3Bf6xO3ubvU4crBp/CSta
nupslpcTSjndcj/OgRkaphk0x6lBXy/A7GRjAnQNeirTYOebALH90JYGfD3R9Xi1
tfxUTwtyY/KLMOchdIsWz5hX2JLMdaZVbs1zswKpmE9Lky+safDbLXMu5Kd2L77e
n0VS0jTrl7ZMdzOKJ6kiL3BtZvmyunpnLhEHD49y/P6uRNZnsNi7LYlL2Xg5I+8g
J6hRws9qlYl6c1/ZkuPRCWF73o5dcVP+rhttskkVepsLG1Wp9rBLfrDrkWtc8W5W
bccb0Smoa+TBaq5RXhtILwTIqDaNjJUUMXEq7ORHlu7ZbsjQnwhhB7R9WHeUu2cW
TG/8+uz7U6x/XLywSHhuIh7ocIKQ1kBrLggpEfJankbUiX2BYGK3q90KXQb3Hei2
BhCH2TOaC8FJuOggDY3+ExfD0t9Sc+d17LGAkPUuS5FErTZgYTqanCc/wdTcZQF8
J2hJgCPgWPp+Bana2IBUvcptLdMVk5wGFmljFYC8YEadPHzOpX5rfuZNcqXTPfZT
iYeSjXLB3Le2YJBjDjLvIK1533om98/V6w/5hlrsWaBdSImL3NS+Hdl7ZOpG8wJ3
cy8t82x1hLb0Hvw0ldnBf6DhZUgYfQU1S4g5kF4Nq7iB6dMvNqyx/0d8BvpTqOZF
2xmSVY1pxEnkTRk4vZkxczaoVv4u20CkJSYzAfa+F7Syzcc5DqhJZn0Se0Tc8giU
gEGxYlFVXn+Q/VqSO2xKm8CCxcKahACS7BTlsyoUXgVzUxPwUs0FhZFcmoe0wjOP
gZagcy+sjz1LIEki0Vb3AMoczfjdb9Vi6L7sbzyHAcZyRgWQbAj2qHfpGzmYaE/U
JssOXUzVvcmrxhBYJXOTl9CwQDgzRVJFAFKxPwsXB7dDfcPGP7S4IiMN+pU4SZXq
MdKhQrkqmgTd3iIdDjRvdcFr0FunpL2fLy+ppxGUvXNK2Z2L8bnyXNoZSaGhO2GG
L4nVLbvUrKrr79kVvvufkxbZBhRaxPIaGEX1mLAEl4Hh5Sg+QSCQ2Y6oEmkKlovn
C2gm+cntVdtGBQWcv69j2BxWE0NvbpdLYKHZhNynUtu1TQOri1AXczLmAvp4fgfX
idOPC6cOFkIQ0+X0CYd3V+stuG0xWnLDYEuYvYsWaaaRnH8INnJcRJZqGHvqKWOA
cblR/Ya3lXs+IV307fdvgUiu/I8QT6nFSe263gGiavN8mDFgGiqJnjCfyD5OnUB9
o462CkHhsCwqcITI2+aZDerfg8/OcXOk8yN/tTfDyCd7PMmvbzv+o7ERct5v8nBw
P3trccVYPZ/RnMwBDQBHRRCHjMVrNxSeHrPKdwbj4nxHLNWw9eoi86+FM+8L4Jbt
5UF1dvBTk2NV1jJPFlX+A9skO/p1K2HHLKx1fm7TfC7AbGqdK9MeWEmU761lCSG2
bkocLIRrwMRhw0BoNPm919OLK0Rj9LvEwCgPyz8JyI717tzJgYf47IBl3bHnrWwA
G3XUOcJTa6mnyM56ck4jrC0lbPupLXbTmvqakxeehtJB741xwnpVWSIY8w7LgTpC
BcQs/nAdSSAG9MESCFgNKEKogaosfpmLWMmwV44vYHQdsrIOHRapfwzv4rG6cHhk
YIbkE2M2/imFM8kimzpZX5AWhU3xnDeC+ChKHr1IA2AN8rMYfZTJj3mHiF4SbzAc
EaGDEj/Eu5+uEy5+i6T0rLN9tIsdjezZaJQHQXIjLIg4u/E0BxiIbNX+8KPBbXpu
d3P7BbgwKdsQCSe/QabI1w4xJeizQVNmUzNFjWbzIIQa1s2KGgSwDMfSVqk3FK44
99vGi0xSEAQHL2BfI7iOcPSltSLu7193k7QG0MmCaXmcLLOEpTyrzxDqiKJmtJil
Eg1VXRnzrp5h5Y2lSqoHiySY0r4X3QMCHrwA2qvfXCknkotInrQIajlFV9gA6x2k
SSZFYAncGBpKyySmNbspG97/rFKcvX2ZZq8GocGcCipMjnLhesOp1MfBV621PdHi
acxQ9kGcnQaOKLku5aCF+lrUdhCA4oDKOXAnb6ClhAdZTqTjhvC4aAADfcH25Wa6
wxD1AdScU724AkAb8HNsi5hnXm2kCe8rYpZzT+xT3eDDNoBhU/10Zla8bb6ktAKe
wT12nXHORfArV8umGtH2Kn4uT90vbv7w0GlpK9LTy+i3n0U8rwDWccjImnL35AZe
gIyLimiXUPHnVnVfQYTefh93BgyKcLdzk249DHOl0u3TSAgSJK2ixMO1/Q3JLvGO
kgSOhdtFAUt8u/YQeOEnaSjXluVLTpwDyuaHntHLcbegwstVzE209PKmX7Jnkyyo
TZdy5i/OoOb1y/B/cekCWGCAV2f9ywtssWCKxd8GN3CIs+zWnLJmpyF8ws7D2/3J
T78Jnmv1WMcfLdxPbibrVauSZOPbiLHIiTVdH8FUmHai7ryWBLHJWBiWAqe+mw38
J3gh9AQHexOCd8n5pkHIRFuOphGgV1Jp4o9W3nXm5Ugk8cw2xDAXKVO1kIkaAPdH
IgLSc+cY59AAXicHlTOBbA8tdAc/6AK4YXkIHha6jK69VmqHA2UYWj9ijbMCdbJp
sY4CLAUZIgukpOb9XD4dgyPjp28Vg7Z5C0OsvGmLWn9KyigJLQWx/tLz2ls7LeJU
cghrbZ0JQEtj8OBV1bFXLB+XdP4EozpgmFOsA6Y7413UzX7IhBv8BLAlKzddIHjP
Vj6K/zW516qvR8NLXeBMC+Umn1SH2IT7UuWiCe0CxWW87hTa1ETwcmOOfSK/Id8a
J0iOoAVq2Ki/SOPwrwurGyzwIwGkuLMcquL05g8aAh6pYYBL9/NOWww+2I2aLzIb
ZcyF/PgkYXPpYRjabxG8zpgnRIAB4Oh4B+aa0Eev/nvjks5i1Ng6pLEP9dWwlhLv
SVhb75xPcfKKhwWmaBi1CID5vnX3I0Akt+qYbHRdKO58bSndlh9by9wQMqhnABxd
ffrpX9R4RWUcgFXGth2Oi3ATQ5L+yLS4/zodJG7lQoQjGsoYVGNsYET7gIHWLUS1
PpalVcNAp1ZSRDjhXV1gK455cKdYhPOgtNEBu1fzZAlKv88TDoHCjgIoCaKAvlgn
cx6z1+GJXlNtK+NIG2YaYo2NR83Shi3SMt2THMfno4kb4vUM82unxqn+HotXryXE
S4Mc7r/nlp5mjNHBnUCRHaBCtyARQ1zpqY6QNuNV+7yQ6WMA5R0/qYCgUeVCh4fI
Ua4+f81gYAMcg/WpL+yvK91tUq3/qL/ivKVliVln6VrsRIPqUtSsbDZ1isP4nc1E
q/XzpLQnOk7eRFeJNXBoU+YaefCHm5en/AreijE1C7R8ibpLlcwJcnVWSxmaxfdj
fq2xOFWV8ssxpR8u2YjoVDbYtyDTYH/9AqNv+nOr2Q698Ftg5myp1e7lZUe9Gj7o
TwceXPG9vgjIEelDu2fPMKscjWarOUgjjuFUJ12t3H2kU5LMrGHCEVbIlrFqYncy
LA+5yMZWzXo/W0C4/QmMH1jUJGeRL6ndoo/kXNuK4jJG7oWdJIebVcijtY48vXwr
C55aXB18teMMylcMbGNMClrOfu6Vn9vx/GS/kLmByG2dbAVig5WR9+P5cl6DOcIH
fH76wXs6uSjhxdGpCfLsy3dUIyryAIxESkrITcao4cRjv4pzHUIqkJUOFrcFagSS
w6zIvSQY/hdgF+eQhrbz2pt/sx9q0VHvOPZADwDh1dMgMrmmVqlZR8VICnfbuL5r
Y5uP9sGWHrrDRz3OdAa50Yhf6yKz4+SENOufpDYPTdcIklgy5YXtnYLlZlnBUjbF
a7JyHIbzIQtk14hXyG6ZMZqkKS9QWN3NT0utjXCNueKTG4hL0Dr+Hz7iLFIJhNr/
yG2VqGVTXfevX1PVtWZsg+DberrzpQj4mEgFsSj8qTuWCyI0SgIG4KwlJq1tuPZK
vYGRsqxYX6Q2+7LYr6S6rn9qkTECn5CdidX+fMGEDNrbwxJ65ws3Cg5A6YcdxZx2
KB3wIj3SwLAOvT18TxqG/0KWIEGos427vfr8oM+v284NktE4VBbJ6uzWDqc2Li8r
cbRgNaB5CvZiEO5jyxEBali2+6G14CpUC6PzstxOPJoo08u8hP2fBHm3oFDfYiqQ
ISd8Cozq/mvzHfpYiRc9Cg+fUkk5DAERxcVvBONXR3aFV1bhIIbsVZugfON930Xg
nTTj59sspKjdt4TKV78MoWzAAhMgppb4jGGTIjENunlHhzym1e57KXDIPdxV9PWL
AB1d/bUoWOSil8nE38E3VoT7//8NLpa6t+bdDAwg16pJGRZ9OKHf9Hpxn3KmVxy6
yzoZ9JjElf6ECAwoc/GUbQMLho1gLjHbLegpMsC54LpJLUAYfk567qbAbM4+6R/y
jxyh29A9qeYygKDpcjFy6X85RcwZIF7b5SyRNnuMPcMc8hoTvjdxurhyZrouLUVf
XOSSYGtaeLv6X9YQZanto3STRAJi6Dbd8wCcwNnVYwfdxGjSa3XOlCIUq9psdayD
L9EXFSp6Epb+gP/Xz4YZ1lcfj/VWxBxN3jPAYzjv6lHlKugqZ0CB7qSMN+baCgww
RiUPr8UpZCBO6HjL7R3HF7+sN+hNS2Y6ONkK8wjgu9kMCKjDANaRIFwZ0pJGzFtb
RgapAADEYxOpni/2md9HZxmJo/yrY/KbRY7qK4XE50/0YlGjoLZaQ1v6Zc1z3up0
jSFvgx+foqfYmedM0ORTj9BJAPdKq/OqtY4j2HMaeed1A17BkT0KvNeGH6v3Q9t7
tAdmPVsP+0YzwZLB/j8n/5wT9FFfyZuO/mYuxlAyNBFaKvbG/Og6nIrmFfNE72es
2rlZYZeuTmZoZJklJytj1RcEkuiCqTScLl5JK3BCwVBeIZdLg5m89hnM8IlahEXP
JRJxPpNcQGHuHg89UWyNL9ijZzYscb6WFH+qICJeb8EukCSoZeEsJhvcgHuKo3CH
WEzCC0r/g2SSIefutu9wDOyynZrGX7j7B61OnotT10OUGGsq5bRwNz/j8lP9QyPQ
urWbLDuyek7DFCPh2bzQOLoQDAPTgHuLbmplQcjacjJ3rdYeKXvl/Saiw0+xhpxf
NUsEYboxZJ8+2UczKElYV1PxEBYQ9NhQ3MaHeB0vyHFa8fyiYCWAdlmb8Obbt3cq
i+u2JMrirz6kwsMhb0TPzNGoM1J8D0ItSmruU7JVFfTBELBdy5SR748Lp95gk8g4
xqleqZ2gi99UZ12AIUFeNNOyT7Nj7KcNo0nuS1ZMf5+TDRz7fBhrT0JiXOSbHGe2
Yy1RAtYPuzhWcIPiBKCxhkSuPhXCS3ahEwkrlv9g/kBZyCAfoR+xVlyxjnWA5WOL
VDsc8Y35D7rrDpCqHMrtlsxBNahmq8xBr/yjjIEBuR3s73/9koJucOO17DaZxxbJ
0h58Kr1XEyj4Sqqh3lhJdf7GPHX0E3fFYOHWDRetZvCPBI7jzGSwfxmXDfwsYK3h
ttXxvcsulWJdGUdJ/VrRwZdXIJzxGZ0Og58O6ly8DX43C0ZeDxyJIAOaNC8o9wtR
MmZ5f2gJUiXfamMAs7Bc7wKwAo62De0nnzyDgzwdG8ztuQeqb0S9yFxPCtQzNvgH
3cIBqgNLDXfYAweNDQBTqA86ATY3PjlGdR7PtGYFMbAoYtmoCqrNgeQQ2Tfk11RS
UGxHeb3doxMlJCZEVIkV4maIf3SSsxYYsgdJOZ5d3hH3cm8T4blL3QMUTBG0gQg2
vwYVUZIU7gje+nVf4Z1wJVVbhi+VKPaMweIB6dRZqAQdbL0Xtw3X0jh/JP0oDXxj
CcDsDGGHyXZK8OdG9C32mlN6EsZDEpKi5Xqa31ZUbxwpIBxoAMEub+KlFNt489/M
FP0Bt8ME0SHqtXie+gNCcU8EYI7PiAK8LcpV+zWZ+pgGDWd3AWDtyGaWn0KigCc4
+jM+6qWBLYHinsbvCMTxkVrJk4o2oWi9t5P6uBychvThJdXpNruOZR2ewlXGQk4/
imq/P1r/xS2HejtxJsXS2YokdkWSLcywcaiGXFob/qK9wh0nIkJXcg1vfuBsMJ3j
0dLV5sLaqAObToNVoZ7yqpNVit+inWqyfq6R2EWc0mgowPfCb6ptzVaDo7eM3FVx
5iHd3uz50DUwD1r8f2DJPG2X+7BQH1pMBfE7fzEdBdDYdglmizggc6ySxT0X8KBe
BUcrEDclC/omJ61zmjadLYU/Eel4TkwxCNIe93DmZzhmwC3RhxvI+bMSDP25pHZ2
P0M0L5I1h9zvb7H38G1owd61r3PjVS0uR25DrBa5BLGyiFsFRWZ6HjNtAe540OzC
icIqyplUFKgz4ElKH0mohRglYUtp79LJQL2ybENqKwuOzpG3dHtmbMObsuemq0Nb
MFCHFaRzo5MiUzDAEoVk2XZ752yHkhBfo+9mUD8Ky4LMfblXeO6tVnK488F04LbZ
msAgjUl9nsacWRO462utjbWhVACathXLkkK7umC2ABKYi3PJTRRdrBOM9UGbPODj
wypzj4SDFm0m0FFb1LMBRl7nUW4OIu6cziS6ew/40EsgMUfl9PluZqJBVJEeuXkE
f7St12Q1WRCLqDNXwDGk+AFtUwpqYeaW7fBfGDLHbsdAro/X2Y9q3mGIAPsXawfW
6QTJGpwJMMiMNh4Z1aqXNj7X9ryP1xFbpQCjn0UVAZVdp36Kt7QyZz0p1AqF4h4Z
5G2g5wrGE/nAul5+J1PNORQg+9OZZef1Uz5MaMqS2W4N53E7nI2zTqZAE2PTZTVj
autDNxZdpGccUAH0zK+szJrWNFb2asAlJNPeAxo8TqZHysRA+6kPaZO4I15bKUcd
LEaYGeLo04nNkl49SELHXBN/d7gjOXZ0caRyooi1qJV3M7la7Pj9Wlqw2l624Eih
j4FKIx1XyL6H1xyCj7tLdQGNg6zCm6RPm7cMnd+fdrbYEai/T1ce3IptqqGxXGkn
+1s2XrItRcEVy6AzSd7XWAOJ1jugr1ltv9Fyeryfuv5UAqCTO6REXtfKgDZ1mJ80
Q4VbcyO2KN6qwJ03HXxtsZaVHFkGMfGpCw937izSu2Qv/YH3gej4hnkk388de+AR
yT312PcNvKRD+gbYCRGzvgJ5fo2LLhFjWJu7PoJhaqc8YICJyzMnejx/zRLG7L7b
NvcNqiIeICBysCezA2Gr2u5tD3vccfhRV+pLQuTBfMf7MorZdtU4PpFbf4jGdLDD
7wYXK+cYjJ9RkXMe1qM8LGczrlus8JnME++1iFXpYZrO7Sq0ndbW7STyDII2kN4E
d7C4VE8g6eUjhs4sFVXPq2ytqUxWJnTdtMkTnHn66x6hw1xfBRz6Lbfdr0VozRHO
Oe3T2mFJfIyZx9IAB0/uGfwnPojHpN6AgFcKtN/vufVHU+skl5n0KEtA+ADbjqqu
BkkjwkBns7ZuBoK1XjB0HnOlrF/Up8j2NlxSKxr7Uzu6u42TqJ3Ywueu/L1q9o6E
W3HELYvgdJwiK81abqngZ1WVgITlG+Uav3HoWlcccVgddNB069nZrB8ZUmsnk5+p
8pPdzd/1wjim9uZaH1tT4aY7B7486revdip0aSHF7dDS6zEskZZ9jM0B8ra1Z6bX
VzTPXheXBTU4GjVdpEeMZeC9VvyMXG7C9K4uwoWNOF5hcx0ILxl7AIdd5Rd3hr4L
S2Gb3QgkQQAZnUKFCm6ecSJ0b5R7kpvVmQ3dJnPUA35OxzS0NYcn715MsSBHrv4A
FKngrkwWF0V57v/uvumuZdXtUqoOJNgJvhKEDhzSiNe8zzp3dUFvbxSJ4c8Stnyy
xyB2eKtANQtfKTPRLPKQjU8h0eehmlDPpR+wdVnK+muNInOla/VZQMb3GJcMQpyb
1aoQWejosHkbFdwR2uG63lyuUdhmfnyd4GPRu8oZ7DxFZ70UQteuguZcHZ+tbHG6
5YYpcU4w7yumDBiC0XF8FGoAxh8Hr99GRxBwEuHdhOHIYYy21sFF4sfG2X0x5Rdb
0KRB/c6lP9lBJOKGgb4ncNv7o8GykWfAXJ2020eMmfnw0NNpLmnjqSrn7nfTvh01
sTYSRAhgZR7pcIbW2TkF1+pejWTtmVISMnuZpw/uLOgG3xmVaVWaFv2QsywyTAOJ
cL8Y84jIyTz7Rcpn1SgrHApXTPljmDB7j4YPS5qwjKKwVuTA5sLbCcupGHAw/mGo
FeDGXuJ6pJl1HzugZtmQ4ziuukA8mw6pP2WcwuJSBYRddFJ1gE4GMavmQry+JHfk
0e+yRRMM07aZA3E7raBSWyoVgIP/mkDJF30METWRBQV5GSec/xNf6zYwvS+gZNoU
HyicS+I37F0bqJ5H+8dnXC8IfZbEyFC42oyVwx30U6cYJYIt4i8tV8z149eHc3f/
yRMlb330m+3KP/B8+4K5yGo5bMyQQ6ZB6IInJKqG7xbI2AhoJkJJA9PNphtVTjNk
9TuDExYA0U5zJYWX6YSwetaaPcDxCqh/wGP2v/dTLbWtZbE14GTc+kUZmY8nJcct
aayOrz0njP3xjYxkBJJf0aBudpb5eqwRjLRgf2XtqUfo46X/yp4vFx7yoqdGp6J4
z7ekNTVOtFHWXIlkhML+25/QuN/YCya27euUqo0AzPbNuqlG8l4KjtiwfxsXN/5C
ZAFAY9uoq/2RP7jj+ETni9WUnlM8twQt9zJjwibDtZZSJx8dKhgTdAD7Ih2IlAOj
so2wSpPnEGVd+1LPfBxidMwgjEOAbP4RfpxNco442emnc4+xJ3Ue6ldF64mggXqn
kw5AgaJnUinMPDa311D2Z2oQXk7HUVP2MXHcgzvuz9vQFcog+pZBF2L9a41Vf6aD
3kekO7wKGGpnDhabAIEvoJT0bVlbvCLERiLDvtTe2YGg3JrRPq4TfIhxVLbK9TKu
UoTOy+Fixk3fjGqrwRShw0HkebwTTCI4Mmju+b3aEqb5Vh/5MKKrq49WEow8h98p
6UDB6GuIBbNyHtyNjw60bDvu+UNgqfw/2HSgY+iXwILVe07BZwdUKmUaRPd372wd
G4YN8Qt8k25PTTvYTpL+9BuEU16O0dPxomi38hp07wmLyXhJcfA/hFhQLVF4pfPQ
2UPONeJaVHrHs5vqmmuHiYyaVrwR2kOIfejygRC5stiJY9qv1DdcCE4kks0VT9k3
FMR7bv70YD0FMNJN/YyQWlNK+44kkxLFTsDGRnZL8IsfQKvUB/R2I+LaSbwf69Ia
sdHde8JB8Xozw0b6x4QwgNfRO4SemGiFGvZEY8JaMKh5dEksUOUjElavdpg1cmWb
WvVaJUEiehw49qtSNBnwNt63bQWAj4JGue1mp9E7Ub10tdQhM8rLngeEUchM5eMg
/+LPhdtmLTc4+5VVGMsUs4XC7lZh5Qxraj9r0DHhbupNJtLEUjV6E4DSeN2YarWm
9KA3V7jX/qYCBozm4vBz6QFxvEOswjHX9v2LK915Aqk0CZjiunYG2FRptsKuxmr7
YQjKmVHruwEIh7Eo665Zig5pm5+X6RJGhZ0nEbWTQsgQvE1TBbYw6RanCvhWVQz1
xwL60EY3+dLCY2c9o8RdUcHq8MdJ8Eu6to4XgGCsS9+Pi6LL4he1nz0wv8IPywDG
+7sVn95ujM1IJ60frYPMEzsjm1qr2Y2nBT2U3OH1TEz0d/RG2eTHLqDGaKwLirav
ON/s+KXpbKo9u6o60h7M84WLfs+j6ktkXmrkXZelDNnI+iAlWptOOd0XZYwIAFg+
bIrnBPQmhPsu7suErcWieKSr0ibPt35L+QFFNNWsFVSOZozpJIK745JT66hSWlXa
aURnO6Hnu0UmEoSKPkcOaxNZUyuBI3NO+1M15iqC3aLry5xy+Hiaax1LfQYubvuf
YMLGL1npFQeVxrGIQP8fXL0WQv5LlWDN7T1rido+n9edRDnRq8cHt6g6eWPafYvl
CPY1o/cvyrBvLiNH+wzuvkiuAZwYNg0wPFfb1+kJbGLB1rij8wbwIWgOoI6Yoedm
BmBm1zOp8rxaiECndcpMUrre6DXYGO0AhShAbcaUecrzJ8WDCWSewW36wg4QGDlN
itEFRGWI/h/fNpNebMgl47Abazkpch652rZU3JVHy3Rk3XCgC2Tde2EWxYP/T7Nw
+iTGuqSPC81avITcdmpwKdDIFZen81ts2Da/P93Ve/nHj1woD29vcypRy7s8uG6v
5J+x0BxfeNprS68hvzk3XvRhnLnylhvAQiBeVNTm4AbX0MZ/D7ra0Wu8OaG2Jye9
fdmhsQNADHO00OLruV8bMw0VYsOPlutJYZvNqQCiGm9Blm9t5KK411ILLnnKN4f+
Zrtx3syYsiDOibSQhYQgB+916WSBP7KCVRJPtd/AbUJC9HegAUluiq4H1WZ4tvaF
UreF6N+ylEXYWo/eThJclhUZne5n1Yc90f7mwPTu0T9oBUZBEoo4HQOKTGwWOEBB
adnHciyVIQlWIZg6dPqFd7IyXab/JEldi6Qpy3k2E8M1doesTdDsCvPuOGi+BdLS
xi0syKWmWer4n+n3dclYee+nB5pbUGRLm7VazcOpV9ZGTPqPaSfUW5Uc/ikj1Xqu
j7fsLBS/1WaYzLsGwXAkEGvPXuar+6qd7rgW6nGiH3OHwpBwgEeNAt4dNB01OFNX
19PIOhYQpMD+RPZ6Otbt9KQyZXGTMyLxOV6YQgxABg3Ef+jITfr5IJl+7qFwvd5a
vHoCGUFmkAFe48EtBP/dJU0vjtqI3QmSh3c7MYM2X8GTQCW7I9QBFQ88uuzaIHvs
bpCY4ix5aippxa7nUJNp8I/uAZJ7rFqG7vUqdDgDXDIbnxAS+2/Sa5c6iUmn+uSG
H4d5GJBzfDIEFMHrKrp+7Ze9IYkDStKbUGQE6J32x1IvxpXQ2UV2rj+9qhWfNlJe
6l2sQ2NffoH4bsDjGgncLdKijLPaizXIsmCFtOgPgNQJxc9HKIaSbY2gKqAkm17n
XHDOQqb4rtVm0e0bjJDARntLKR2cYJO2KDvFoffu3s4nqgKo5LOAeZuCOMWp75PW
U/s1qzbv8GhYUriK3nw/xRLg7C1d4M2APnfhYIY124FkTCs8p94HLzNtt0limJPZ
ALNDWB/L2qsMxCub8Siy9cKJDK3eYOf9LBv7lxvA2zy5kcHdh4eRJbx9juEqddJY
RQaMHiF9CeUN1dbt7Q2dltHOSBwSIjWkgDG0TPq1qs0/8ADykAN+jL8OLE5eQlzN
4o/2cmMz0ulstDDzX/2EJv65t1E2jpl4m9oRpEsxLTVyB3vqYiNLC5sS48o167wz
v2/PVHQE8anwLzhencoRlA5ZNjNwb18UOprqlHAQ1zO3lYCcozFADuxHLta7h3ld
m9zY515Z0Cr5oddNFIsQy1ffnz83MTK5wSrg/cqkboIMM/P/mDVoFfRxvs24pof+
v9kVgXtZv6NVn0chiYexQdQsBgTkuOUaDitx1AusEFYJguOupGkOGx+UolGv3vq4
K5IfwXczLfu87tvgFe6QVcpgxAPqhP/mk1K33Q/bwtdNtqU8fMYldEm8bwmJabKG
/DbjTsIMAShv9MdFyUv3R+sSd/goi4UEX1FhG/Qq+o0z3j1kem0w0ce6VRqH4lu0
dwMVd7omws0Ql70Ng5l9ljDkhLhEazlKeuM4nelCAEBzd6guBAFQqtcdPu4GS3Na
5RLR3h1Pj7mfK0NT5JoQgdePjd2tUeTauwoZjUtbNM+fwVPVggDUedkKyTTiVK7L
hNfiDoxaf4WvaaQev1+Ph/BE7GZfUcM+JCa0h04dCJ+QAoKIEL3UGxEl42ipKSE+
/JW7e+Jb9CqWdqtmO77KaqJzmPiQ7nzKVhLqwFzjw9rtpUzRt4zRaH8hqfdz4Dlh
T08bBMUGCtiGa/tql4dJrqJkjMynwHlvgRxnXbCeUh0ORRKDrS5/jFk4BSY5Lfhb
PVM4OuKjz0JkDs5PQ3AkQ/KCI919GewVUDM14HBjmPN4lcmd+asrHPNby+vHvmCp
T0cvYbH5QQzLK12lx3CkdJOACwI6tHxBf+767R7AUmCDWT4E/+vXGjJxk2xvqvdk
rgmh5z2qhfA1WosEuOC81exTfBiUJigDqjxO0gjn9/4qgy9L/bFD4oFA+iUOnH9G
IL3XqQMdOAim33wI5B2rCgBzt6QnQTBEXsr6tndckyUXlUiH4ugcTh+9Ie+9zF3m
a5J+6gDAFL4fR9MFrG06jWzoIbVSKMFTleKOHH8dGuSXV/7/URP3KkhgLdszzcD6
2b+v2T4knu6vzq9tK+AzTS1sb8FNm6OrCd0icJO8RvHDJSB5rxHT5HicOigsjdS1
S9vlM+W9p4qwlhfXCTKOSORBlLiITyvhOHUOimeEgi+1hpcZc/i7Rj3ananitqNG
A3N1QxF+oYOzLkMST1w6Im5FYYug+vyu0IDWuh4riOYxMBroRb3+RYpnvnVJr3lI
u0gZ2y63tKbufH9TJc88qn0AFaFZrxWjJNpPDNXJnKLbkUKrDnGmOmOQEpPVTunE
Un4YR+ZK6jbBUGRWtmU+LH3mYhPJ0xinvE13aCSkjlrpaUSOGPsR7QgFeRYZqqrE
0nZG6nwIbCvGE70I8Hz8Hd44LqNnvpAlElYUiUZN3XxiQYEGTC4v7zRdbbU/bl0k
YhQ7zcSbi0sVQ4vP2Nkc5/1wrNq0QU3eBTzJ6TI2IHQWEteGGaUa7vttm4IdmEZo
XOEDkTaaxBxSBcR2ZzcOoiIJ2dqySbGsvePcWPmDmdzyP5jm14iyZE65tU/zXA3I
Sdh3bG1XH+kTHk40N7j9KzH79dMHyqccq22IXtC0yd5JXMEzj77pdDHhurgbH5d5
jNQJh7jDar6i45tJu6rM+/BjllOl15g4nvfBY/LgfmKnfHei3vYd3FGKITWqxkFu
Rc+oyzKh59zvLZqI7Eog++XLzpXtXiX7yIfj3tmzlkNPPfbRo3c7NG8Ply9shZik
JXKBAKozizkWQcpM3xh9a42FHkn5eSndTqbW4t3zoqzSsx5f/wkd4V2S4exy8+Li
NsQn+uomAK3lhiWOmVQ5o0vE8aW4pLikcA4GSEKQYlW3Ei/Ofj8iwMt5LtgUGPhk
ok9/u2dzJAeMGHsP42umnVFTzax+YORfcdenZ7LljOwWkGLqcUV5H6uc58bN983m
ZmLAoUlsXSBCGwEZOnH8YeTN9VX5cOaiKXDdZL4iGyJq8qAgqEJU1IBHkEenwYWu
gR0ivlZKTN5HY3hUl/TD5bnnzisV0p/N1KI7cNGWbj1a94hHo4+yKANJ7/hgLjqZ
fyDzNlZ97fc+2cxdACdwYPqGNPtnFZop2vVdxiHJiyDtWf3s8F2yEJrnlt7FsHC6
EEoDmoINiuZVEKQss3Ff7X0IgqzZiG0xLJxKqrFVWOhC90A0VIaRcMyAsQFKQe9E
PCrNknBJ0bjai20eje06bfZZ7vgTTMphwytxWWwUwxX2olT90fEfLWGUbx5gziJZ
TJtIddzhkc8VZOUl6IEIBLTNhgscYq1GYQuVPs9AMm/QOv3jVhtVmKycsAiTSkqK
TM8ZeKOA3QQgey+uL6xFLbs5Q4PghIIRc6ZQ6FmeLzQvSQ1DlHsDQdBTEawVBeFj
VK3Zh/BYtdDekF/j8tWT8+0oCQhWDMqF9v34mfyFxCj4qMOzUH6OrXw+2bvfNewI
bN9G9lmZVEiBm8h8KQuy3Ytpl55x+8OdMCMKRLN7buncdHsW0VZ75fyJMB13+69J
nc856rTP4KrCoCRJhC8pA+KTzK4WjXS6Tu+s/sBma6RMpqEOKAppxX8M4PIa9QEX
kRtkZF54y1DW7RpKaDtxa2IEhzIZafn+LFysPCs5PBj29Oe3wsuiT1kKpS4x9yhV
zHAKmRbO9TwHgLusFbEt78CM3klfM1p6RCJm4ZwmLlw0icBh4vrin5+A1uneOaKr
1w2Z2udmhj6FMRbuKjwigGJC16H2uFK7HSC7qnhGb+7zlhxn/u6r0ky3b8cE3Y6y
vEi31d/UquByxbGg6HRgX+DSSfVJXwXCn4Ogs54+EutmNgOcL3D3hg/qtoLq/SGV
WEoIZ8vCRNJ4kT1oHLcZqBc9hvIc0vYkh+qoqanQkuk4IwSMHOCYqMCV5fU8u+Ap
tWzB6wSNYByurWtx6aWYNnbRnN4brWM59SyK2lUPyJrjgxtF8rNZoxtQtvZvAkWI
7WyZ0oZrqG5m0So0r3bksLx6ozHWjLmp3KOsqIsPUbw5NItA3qu47skdSJIucu7f
tvA9NyjeWdhcADhzP47ggizsjm+WocnVhxe/YlwIdn1swCnWJNyet5gyevMkOzpj
uivD9f6fdMpv5z0TtvammYltTnro+uQBT02uALqFbF1llD39dpfvBvF+kXl425SM
nCobvl0oj7g7wI3tExRe6um8dEsa9vI7LJkhPLrpXrE07zrEPTq7Gi5g1o96l+am
9GR7Ih6uduDHGm3LSuwfRuf46dgR5dBp2bNFHbi8YZa4zOKpvMdksGc9JkJogOGn
NJbu3w0fC2CuH9tnMYuI0hnZSV+zKx2IlWBgMrElW8ILZNWn6ilgO0cLAlyvmTNA
QZpBs1iWXDi+QGwW9MYFkznHWkjdjs7Qb6eoRztCKUfOFG+ND9a6fY6jEqjHZeip
NW/jpj+pOexuRnvC6rboKZHYcUwg2DuTdwiS24OnHEGCowjr191LDXxah68VL5+/
wINgsJJ0EHBeNrgs8CnHtlDqhrpEC6qstyI5KtFjQznLi3RKmet6smIxBmJedL9J
3AUj6CaT0mS2c52IwdihOyucnVoWo/326sTLTvZ4puISIG5i0W+rW/hgF83OSJHv
eT5jyCNwOwOr6ZvUadsu1AJ+Fgf/td2PfRsGLwLiggAu+fQ5OJARbQO0EQy9WqzR
DZD37Jx0rFszu/+FDMsV3NxkcQkI43htnmzsQ64bXGznGaxl5tfSG+K6yvf+jYs9
mV61ALpuI6L+Q+89ZE8RRGwIa4+ByP689cv06d1uq+zdTYzaZ0eK2N8dTS8Kx/BC
3UNJ2LD7a7YVrH3aqihsA94eZuXUzvYiF1XJnIpdEwYinXwTDngI0jqXvHWyHW5Z
Y5R9cBO3YQ9//70coJq93L0e2yfS9Hdzbzzx0saqfZwdjgV2bX/0yyLL3YEzgnuA
ubMbldhlZler20XvTngqyWYwiO9shunSRuceQuak4YklLtSIVuMvtZVRq/FDmOsV
+Umn/2sahw4tvgkcH1MGgxsF6BzBYDtEciwWSOE7hUR1c9YEXe9CrIwZukS3pXrT
QrAbvo1I7aq0xjw0RxXslOTyHkyDpjYwp6syewLcEc/f+fk0s0IHMtXJMN9/nib3
Lak/mogt10mgSHa+WhBaunK2VbQE0gWIBrnGC6QiIPLInt1zal8KrmPCfsq3M5qC
M505fsRpajDxT6omBWiHWMViHYPosoadzzoD9pqOEPo3MZhi8OJuzp6DxlVJBbMq
C3YRYvjMGPv33vAzAYHza5AFqpnnlXOk/neoYhbGuLb6FNJFufMptLYfVGxw4Qxg
JZeWAeooUv3DAfSuXwqcLU1pojXk2ycGHwUlfMDSN7cCaQF1yc/rY3Mp7tkcWaJe
r2XhQ3LAX4XZvlVMCZGp8+pP0U/0fanj9ADng4cvduyk0g1LVLrulJcEkQ+1gE+7
LsWe17f1MM0BIhfgxtOiKHJA4r1YsHFuo/vVR6f4abc+/SH5Se3zcFypVE5N7JCD
RjNAkGYarPdHtJODbsLCFG3PtKmHxpOqkfgZ5ZWVgsOsQt0O0XlhEFHxDaR+1eWk
FVJ+nnBgI2I02i5NWUXlKrxT3VGAl9TVR0R+7IABoy1C5iwgzFA13fnKiOoBVcb5
oxheay+pGRhGmi2QqB4OwKbgTfKYHR0leBmLPHh8jJFYMs5sDkW3bmLHR66xoAIl
ghY9wJv5QupU5R9kqfNVYfKnpMAP5zN2HTlISR1BaZWGAI93QWHt5XNk1kQI+O+p
EJr7BXRW35sLR7ZjnGNxbozBGaAdsASjc3/9PPe36Ps0yps77tsYywaX7mfRe8h6
JJQ0Hw5qVsiJF4UPYNiCnwDYTUO2343tkQutvILc/R0w02jL90CXeOFO/+06QTey
/k4xkVa0F14PNE/rYBdr5ylF4VRdtcy34zdTyG8IejLORXixI85Sbkf1xWFd95dl
mbVyt9x9l2Z8bL0BThc3BQfVBjnbY9fnPzUJcWPU4emjWCovYkM/ZHC/IcIPH7Y7
fPr1W1WSCpBVP7vOQp3uh7M1b5o/SoXCOnftievOEdi2zjzbhwT/FTGfHJANgLyd
bMXRc4ryWMG5Iv3VohhV+SqP3THYWlJK3NxincmFzvCwx1XS5f6SM0YTDRgbdBmg
V2PS6FujPAHx9FfL04aQPiyrjgf0+A87xBiZkwGha+HrIhUVd6bvuMs3t+AU/bSb
s8xI3bWTtvDD1V3/saXe7FNHh32pS+GOU0GOwYCFzw8iFOPW/8msaMEKX6YmXoLu
fZzcbvtioGFYGAR2SLI/ocg47dKKI5OEE4i4+eFaQ/K11m6c3Uud0Y69po4qNImI
OccsdHvdxwsdUw/MGciT12WOZiavxr1PvXvE8+V3bwW2QS0okjZ+eIA1TVm0krAb
GzwQUwc8CVToMcZylohXsLfG4WazyJvfyqI2qISi8sc3M7T/mquBZHjl8YRqANQT
RyxWiDpbRsatGXK/eyBMI3d9jZgWifvBzdQfF/L9akAvVfImNZhZUk12gYcMzGim
uaV9PvAdBPZA6YcUxHaLwPgF8968rOClE/2jA0KSjnIU+TOAKSjwpuycKnTKRfgm
SSQI/3Ne7PTPVpTwBGQnFQRh/LIT4bBj2N8vDr8ov0xAUsUE9G/mxf5Mw/z31p8h
CUEoqZDfiX+QXT/735Bv7jARjiBvuQe+MzgI7Y81Y7qgkgm5X8i03AhhMcZyG5Ik
QItgW5VPixUt1SDAPqPADQinvrCmX6S0tq5ZrqxGrVJNk8jcaGPGKuDCknFAoyKB
XHUHz5ae0Bfh7QOsoap8YLSYeg+bHM9stt0srYBs83cPiJwXBWtY0K+2bqJpE+yu
IWPMRjfFF0w+lNEzOjqXDbG0vHm3hiqyh/nlVXH3Et3IDX/lQf5nEF8htYmBvL9a
d/Q1oE+5M8oTUwY4thn1A6pgmrxkr/DYOYxijjWWb3yGYaZMxQ3Cpsb+d1qVidO9
EkIaVtbp9xumnzRuT3Er32fE80eLswZPyi4yG3Qdr9sFGvgkjrjr8KiHpsS1tWya
Oif/OU9eHUlzxPCmXIF88zvs//QHUT8i3H2nm15XcVtMTPpaS8yX5Sky+mGbW895
TWV7qmcXVsgRGai4j9HMzcNPOcXoiXW9mDi+Pd5ANQpDK5IxlTVSg+hCZQg5Pr5W
W0HoZ2RSFiIouVCDQ9W2y0OHp2w23vJoPjFJx7RDcF3XG210csBfRAwltF53MXN4
mG33b7dX8dS9D0XKcsyxuulFT7ETKJH3SwTL2jkv2Cc2jR0hoiKwuNwrGflPS99+
5zULEYMX9A9FhNKH0pbUF48ObTWIPvdYavyv3yBy9omCv21eRoBmpsy0vI7EYmUU
Zs4zH4YMHrxS/PlVtVwqb/zn/Bq7rpGQQdC/yj0ITjuGFSsANA8QeiBvSpnXvObO
fh4evNwInnUd8L8Wo+f0AVIPKJsnnbYomBnm05a6sYrOWy+AKIQMw2R9Ge1sP4z7
ol8D2AignlFehgNrdyus0wYnzYis6VB/oXE0qydT40EY0uSA3cnGrZxCwEBtwvH6
BvNuTXrOALb1/wEKvxOctmEqO2nyrFbWZaNmT5Ka3kWMyjnQq56Zi1nnFuPXxF0R
7BQANXQO/qH5MikEEiBCzvkT/JAXkiO1dzu5ow4L9JVk2TiuiTQYuGPW5q0C1IjY
foAAh4HYNGFeOWF0KhTNJ/elTMLW/HEMj7N3xFbGAJiFj1i0wcR7SwyipqBEdHJ8
NT4qwy0u23UJZIJ9t9Z838XxLC0T18u/w1N9ul1oFNqzMoy7sWseNHUwZl9NNXnm
pUvWM+uvCxoqtD7xp9ageMC+VzMgo/Fu0Q8kwmDu1zDAXlKrSAE/lkTG7in9g3+D
rsbm3IPtSTh96oYmIdzTgf50lo3Pv4YVHUIYeOsPlMn3PBin3qhhTKLb/N70JSSd
YMWdonxGMF9+YqDzV6x8iNOjjrZeLnOevS6LNAXAmfvtLFZq7j/ix1qF95KdunO7
eNTiIoJba3XFXrgB2If2jzMEn8n+B5zAm5SkqfcD0eQUYKfsK/zH8RX62hUcYz5g
5GAb5WK3vzmnMrcZ5Spo15d/MaXzIF2Gfi0xpcSz4hp6mfCqoDD0zIPOCiYP0Ydk
/wUMJBMgKBfASLRjo0B0UE69Y0QSMl019rHNZ9Bk02/7zX+cSFcK7Ok86JANtNQC
79sE4tdJ68LFclrXnmkPn0U7gNOzR52L2gIPvs8q7KXjps0wKITUr4H/Z0B154Ys
phFNPAD4NaOz8auk3ye52sS6tSOxiWqh7j4z4X2eHbjC9eb5SrjUylCxNf+1qmpg
Vmy+qMTJBOSjGqYSPdt4YIaq2RdwKyKEF6LOKTJUDR9kQWFurDV4ZHok9pggFR3I
3/WD3FyY5mXqm4hg7eFNFxKKcmFKsPdLFqdgPJ9pS/T1WfEWE2lYudIL3ETcjari
f1vh9/B9ctZHB1T9Jfj8OZVXNQM8lphJJQqoE3sJ2X5qaWj3prTfk9q3PiuDxWjl
78MZuKQbjDqP2DDzOl/rIMT3QMkwl/pAks43bbKJAsmu8S8sJ0N4Q9cOzA+NDP4x
s17TY62spYCgbxFlP8xA+XWONXLCLwotU9em/sYbJN+B5gVlkkts+Br9mcAIPNHJ
8qindBeOVDQTvsPr7bjBW+ibZnBslaYbAAvUonSASorEBU69+eHoXJJi8K8xMzJy
k2qTJ2zmwNWCCUy00SJlEJtmogGIazlDvDZSrh5sK9w4yOyeWs811KhHqTKFzugA
U5XZqqJV76UxkPugamx8ikgOIJKwwH5pkHIsV03gUJbJcX6m5GZIUPclWtMJ8Vgl
uZi/yvdTspxloygb1EpzQs2bFM/iI2dK9eAWtXM3O4e8+zP19446M2zy6CsFGB0w
69WgYdsfmRYl7twzmgkBtsRF2s9p2q7rkY3kk3ZypN4U47WRLxpRUvMxYjJTewbr
DayimUSYU0Wk47R1AtYIoy+FLGM9boc5Z4JL5mUEknv8OZQZf+FR1xWNLgKW5GVw
+dCLdILmDIJ1Uywp89yZn/kcV91Cgx3ZjMNtbDH8yEiZ2ZSTgNQvaJveJmUF8ozb
u4hic5sUGQ9TM9+4cV53Kh/MAEKTyu07ZmFZm/Fgfy8aq4XLqXXxXEuhVto0vU1Z
yDvcTOM+lBbDxR3gyQsIwAbXiA51GnsjKPvpnAcV2a8kVtg8oYXFR7/cCPxCU41j
VOEKu1g1YtaevHtaqcKYDKLx84JxVGlIhCEw1Ydecp23IR64S9iBv1hD9HarrV9y
Qzdg1mkX8wk+Lt3oRIHbEyxKgr0OsIE6Q4zVyF5wwFfqNK7TSZt7RV9CLqQEmiOw
7GeO8U2sGqTlwYAeETy68FXc0mCpIigQUzmh1SsOTaG8NyCuJI9ZPJKPXxqvEXij
Onhb5Lur70gWbeW/CYK02HIYondq1SqOxEWZ36CLJIKKVQIti8zuEkkgtxbCwYRW
Wmyzg0N+WVUVR2953cqInJGVoJGbj2KYuJMrBI2f4iP3440EBdtZZL8rkpJW1XCm
ojXTBruoOyar/2aT/IJNQ31Odlg8MW0SScewDV3qecs+WgAv6ptjFobJRwyZCW2K
TAdSr+xuRmvMDVNaRw6KnqHE+QotQXV6krDBtnUPlEaDzwpTNHmNyK7G/yfTLais
CwGUVhztClgz4OqL5HPaRAIKCJa4NHwRvd2CenT47YSPIAm2bokd/JgOHAi3EDDE
/sABp234OjVwCIfcSm3AikYYGu6OubWk4mVZl0XUpNYpQ3RT9PXny9U2DVGqF42H
IF5IX2SNvYNtb7+6rvt6vkTQU/c7x9rDfLk4W9AgsOvDJATweLOKyyze8UnFQPjT
gTG8UDNVgypMXmaRhU7EYzRJgcG6zbhmvSWv2fnqEAyypYHgeaDWmMqNrHjId6+j
kyAoDAGzeAsEfU4/JLpYpwjHmTP6gFZYP4GDvBedFzUI05xPve3L1rgJI2Ktl+ws
u1drF/egWzMo+Z8QH60CjtzO4aXvgdaup413qMpvxzexTprT8ZETvYsO+oSGSvJB
FAMbVVWTWwlhBj+qjy88IfutJdj2dIihqrqeLwykWpRigZWMhvd62JvFU9YdVimT
xjXEvxFw1gRvLCPqk36HLugbhBqKjkw1tHD111QOP/fZgH9JzzXQFvjQ6ZZ/uoN3
gtfU6AIDkWakLOsxGfy98K4rGsodZEOoqNnwCC638MkTxlgwE+EHzGdcAKyQmJAE
y7CRR1W/1n97CLtJCyVdcXfz5AyE6fxtk1s6uEob6k2atmoprf8HQgkycmZuzNCi
VvlhbD9kaU5xPfaT29d+iE4sjmg/+qswiEZmqdcPbHbdxGAHtkAKdrvde23waUJ/
T4UiwkdnPes6GsKDHuFF9uu7F8OEIwWhh74DVhrb8piEldqPvjvJY4FkNXgnBP/Y
P8gcsY1kTpEqBmvc0nIGLZh1gLgFz/CnRdRWntjvJahuV3HI5IA4sXs4j9cA90KY
hXUQzv+KvLsdqMF2sDI8I+kBAhCBmmmqtoHZNveWehOC0sgPaOA+r2R6iBKOslS0
kixQ0VPzkJfS6NzRIS4zXcaqJHbrsPUpuRaRZFHRhshiDGrxEtcfEkhz7HZdw9+J
m59eag6Kxa8u6YX3YvbtqzQeL6TJE8XUS9kZzi660YBDfRpmRYqD7U8YOdav1QcG
F5koMQhz+FVSTECFfZTOIX0KnOtUe77DkrQZsCPafJVm7gXP7ikZk+8IUizswMpE
d+k6TE0F1c9wbdDAgxyQkYbG4fy/aAuRl6ay7e33+Zqy5QL4UrfA8mImOXWuBohd
n7UsSYzSE6/fmRrwbtVfhLN8uXCnsAvlK12VfaQcjiCSmvZIUh6x0ZMRipVf9/+a
NsqHlosO1yXxD3LZ2qpFV9usxbncaJyfIaCjKoSkD5j1tL0w6aB0eqijP1AjuYzW
5YA+faOfC23jJUbjP77kG80pbMzg3RC9CDRAp78Jl9N6F6mWlY1EWrZtXa22LwOF
rI0ZGKWwAiBTOUa67Xhl1wP0XRbwLFhhH6fECISKkJtX5jj6pc7y2SADwmceZTf0
tQ6XEy3XzJGyp/Dz8DnQius3A8rMCeWjAgS2MLVqgmBIUg706LI5i6H8slUcARHd
ZmDL2GDCgSlto4FiDMelrKFOPb8bsmKuJOa+jiJYfxJQXrbq7SJH2L0ecI7tu5TY
UTgQ9qVgSnqVyDkaQ8DcwXxtWNVUjYAA2YRJLIOVp5P41jh/jydl/m9zi6pZ16Ov
/ntLnoXkRR59owbYT9/Ung4CGRTR2NAApzRVXUGuvqYKjU0kzOvxiktVjCDh7oC2
+B/a8FH4qslFemRYhOxvvizs/c4BOLeQ9UsSwO1MwWIo0xotlkaDdc82D02L33Rg
UidcxnbFhi6VxD9DvVggo56AIb6xquu/+/iODFj+b9IFBJueqeuc9rKep9vIfSvZ
WfsNIvgWMhqCjt0tA+VLnjtJT9HTunR7sVK87UHkjXP2oZwwS+2fxOPObk8jnd9w
52rlTeUEa+5E6hFD7hIuiWDXFn/BT0wdFZ1ksW4M6Q4NhkAvULtWzH4i29Zr0vYn
dIL50N5voODUjIYSMTWyOyGeIjol0Zg07knz24smy3pK/ebWgPyaDbHLlkAZYUiA
Eg/j7KmwOcjr/YPwFjKqvCtWkpq0buz6C1e2k5LCV0ZG0TEHNC1gMNeXmPCPxjVg
zXTOBntImTaxPk4CA/zC5BorLjOcUjAVvCJZRXq8DKshu6WUgtggExwX2KSjIzmB
nGZQk8wrrvrvOkhZBaXpNtFAvhpSe/H2QT1qea0bmTeSWa8DhYbcbdZDfigFCDo+
BxpPJz5l3NJ6D5LNhgrgxbaYx/QsJIh+LLlQDFSzPvsu1TMdvOXBlitHgJqbMUBu
EYAKDmoCQBCvFCalgf7S6R2d1tuwvSm1qKS0UHzjGt8Nzgifa5S6ALc+YjHdNQ8b
XfB7CzkJCqMrVMh0WDgvJd8Jvmgkjkmsmj89mMNcMxy+54OnfLzIt2eFC+SZHTIX
y7W86pR06kumovdrix3Z6JDaaJQfsYEu/kmTbqN6oT8PggQtPV4EDg9a/ztc9lgo
djJPwlThFpOdNb4Ke1I19KgVmm5D1+TLlmLX1iQgFsGTFApML3OgrOqEbNnbm4Ko
nAkNNF7aB3RXnwi4hloV3R5VUTb0iThYCC9HX5iOOfxo9pwAJyp2PmpoecOOBc87
8FuyBLCvx0LPYLh5+jjfaPwjsL9AQhw1pK81rNjhMG2fnMPcNc8PqrASoa4y6NeH
Si1RRpZLtPH5+N7lm35XYukTHjAyGfVaOHHaGBa59lCmjSlpRhO7DffDPzcNaY2a
XmaXChntL9az62Rn8XTWIo3y6trTRTm/ySDRfLha0VtTZRbteApgNrUcQST0Swjc
phvVm2BbPqMlWA6yuyEDjDb08f+5oX/jDhadAa68ghaJzDjo0I3c3IdWVQX63iQD
5GySU+VtyoaUKySRqkJlbwnf8m6igME5F42UMyk+d5IpUVfI+n+d2PyPtm24MiTs
vLD8bHr4R94UasSR1sKrvkcAWJPBLe5WKcMm5CGifYMYA7325HT7IQIrECNLsqz7
QXwf0Wlb+kl6uisNyR2n06Qx7KqRQyLNWcPFXkA66mzCQ1ko30SwaVIw1vDfk730
W1tkUt6duigBo3w5c7pBUxTwe9qouB2dX1tIT9bAqJXYVztJmlRmFE5FyJsFhYRX
D5qsRPOExWiNsCEH0S3dcMSiMAa0elGRh0EQrjAlQ8mpbPuM0fpNjLvSbmZmHvJ8
DsfO0hhOz82wN5Ik3ECDzGE5TZt5gqV73y8WzLhryKMHdrjlylXjG6tvlZPRHRTW
Ba+lwECqq3DFwd3XCzpGi9uba6HEU2T8Tmiy15zHjBkBc0afRV3ZiZrPE0/ijclz
h4KhvAzWs7ERzv0K9+8Dvj6D7Wici2inh7FBpz3WUBIGGt033iZ2nJVV4BciePal
4rXhCtkXKW8WSYKZHIujoizrVrG7I5D5/gQoXHBnT0jKufNIZ3Fv2DqGbmZPvFeU
1im0tCFk7DNG1ylTQP4hiosybycMs89ARQgYN+TzzXn7fAi4ruCwfvu++VaSabot
dana+ouMkCebHGOR0oaQ9kf0WpGdllajT6Ty3jYUfsJ+8DuN7JB2b4snrRs7XZul
dz3RiTKrC7RGbjXjLWwWxfc+ZNTm89jb5Xgqfdd6I8nZbZLMwKJOKwYHMkmkP7L9
dZi5hgsfxcm44itjvPefH5354KaO6McfCF4o5ESOY1nd7CRQocCvjiebHDuNejxb
6nAtImG2vjgxAbxIoYiWlGSgwg8tnb2I/3qQY1j/b7imJJkC/lERS7llsigMEJ6d
cHQPS2F2//aiRXlLSKsOa+JnFQSxUBKtyeV3eBkRaiumZvHalVuCJY+Mxq4ncuac
sogfcj/GXtNfq7bJRgaUX1s7tmovpxdEUyEsEhxunE3w2TyyEecUG57pNUf7Cz81
BI14IPJgNl3vP+6HyLi/DGi42Oz6LOLhz80JTbiTpIVjZX/iL2xkW96NrAPvqzdB
FNZvSjSpdTKo6KYX+T77PP379DDkfB3jN5+4hNSStUqKJyE5khZYAUMX4laUWHhO
y9sA2mMIyC0JGFJdYTFbIwx5P8Je+8iz/U/M7HwKBWTQuUuSJecZvnzJ4KEWfzM8
yXjFtrBxhIzpMv4efI/+LIr0dry1SL36h1zwzqqucCRBbtEc9o3nJqBG6Zvn1eRq
YF2KHH0x0fu3s1d+GEXS+3WdEgTnhpiaP0jJ/0Q69bVPwCR4jLbFmEmGFrfVTq6H
arY89QNTrfcE3XG5WeBPbVO9RmojzscpEmPRCfW5243m0HlELlb28RhaLoRmVutK
m5Bm/qNkGTuYRF/mZR0OWov2jPSdwoERg9Vj4gb34uF4F7P2yfJAdYqCgEyQxxPX
IqGCOSvU8sIOPvSSuPWH/vs4BTK48CzoE/KgX3WLhZQ3pFymYh6/R+yp29P3V6a8
V35suTrqm3c675Ku1Nugy3I8mhg6Gs6zAX86+cYYRSnDOnuHKqhI516M2jVaNbUn
9nUsvwoRcnjY8X+Gti0xdACa3tS/nq8HGS1Hji8HfTeAAhWpnA7PB3Yvz/XvGccd
SaGEpDD3X4lsN0YEgTrodfVFNDv++BcrBpVe/PR8qSy7qESS0xU4M7o41gZplSIy
2/i5I4/9ducAG5XnALzdizmYPpuKBWcpAQ/7+DWFrIjHlunLP+tfVXNX0qD7nfPf
EbcIOuIB6OlP6XtVPRSF4dqtraisc+KuLoj33SUAivBNjz9PVqhuEB0yxHoNEogx
tl4p94MSCuMEMC7ucD3cLnQ2eiEbzUsDQvNE44wr4XZprQcRJNULbEe0dHurPT5v
B8siTHObAtFUhAW+crg1d+jCcJ0l8M6BQxTwmGlGtvhIuAgN2azCPOXqMsoKKb1f
YcPJfTidfQkmTOd1AThdX6Yy0q8BIMIqeq7w0GoTDLXDsR+h3s8eQJeE7+EpecyK
YKBYrNIPRHlhO9sKyP3GuMrI+iq56T24ZNYjodtL6eOqFxWPRCgTzw7Mg86w2nZx
wB2HvdCN12diMu64XKJIWSSM5kl7tKrZeyDaSmJEMYX88NdxB5ZAOjrimST24P1e
WWFRIK/8PV4UVPOzilT8jixMxitr0cSWWA2XQBgcq+bDaJm2rcH5ACNSrpmYGhnJ
HQtV7kRWknwqoWkEEjEqf80S4da4uQBzj+qpnpZrlI3atdgzMO+VIppvtBJ/uhM/
5Z3Y9tuak5HxxDwTVn6LI5s6e3xg3gPB12CbQlzNtfnNEqfV0wXrpBEyi/vfp97G
DbZOgDdalPZbc919xAJnzYzK669UPXuGfzbJ0JCZt1+YDzVS63X7IxRqYivDwZco
MpRWR5eJA3VNhGkiAAU6QxEd+n1wSCQ6CL15m95+1fN7HU6pEs9oGSwbLXwS7sjF
AePpy5YRBvzijSwRHnb5a/ZzIxA3/sokjTf3QsNA2Yo9NkAwsDVhoPeHUPYAhW7F
bIxD44vdw3ZcS+0aJRUPOTl1S+EFU/+8PxcKXH8TAN/mX7I1jZshZvUgsOxVADD2
TyMkb1VVs3NEKTq3rYR1nsUHp0pRjFDnnwNTkYXNo9tecyrAHlzY0jrjcuY6IZC0
26Gs3NqWgRP945YLjDqXgeAJGbO/7kjoM+VyhJLeXt/8yVMA1OQg1XwaQwQjbLS7
2GRZIK9F41dK2LQ42kJSnrb4nTRsLBdWmjGeMXbVkziw9+34Y19cPGR1c6ICqCzk
G15fHuU8/w5WBqb7uBlhkOys2Lv0vdVQCrDh/RnvA4VH8ER7y44FNn6Em4U+8Ju/
lAvzNb47qZTgkD27qjIlwXuj2L17bI6R1L4sNsRylYFg0dJ7N+xe1WU8/5q8RmRB
MDEHE4bIj9pb6uDwXrF7cFS6wjlKRIai/a1gqNAztOt50upysdW3kNqpLbQk7tD9
rAA/rAUF+u9rZyYuG8RjN8YY1qHkRJQRyl3fZexbHRhm97Mk7k6MlyWJiTihng2+
tFSUhfsaTMKcLQAvHx9COe0+uOCrdUt5ytHK00OaxR8TttZ1HMCPS2UveUR4uvzD
fekNiiHhlvoLtdaAxPyVauam7HkuoEe6LuxmSKnzct8VCFcVQF8Xjho39f0h5LxH
q5u/5bV40Lrw0PWrGoGYDP9+iNpsi1horN44/WvwhBEZTYKZoDRWKGe9dzBTEq76
efXGXCzUo+dPUsDY+hc3xCwPur4rKPlLNyvTkbCuU+sKRjPTQm8O3ezxkE0qGxLf
wxaMKTd4cyfnnGqdxuzG6QZ58O/8BmduvVlMzAbmApMMfI2RWYbaBlBXXAF2kLG/
n3wNjLCTpBJZB8F+h7Wtg00CRW7/o12OeW34EHizHhskf4lXMBr2K/m7mNSI8XNZ
6RYrAsYssyuBrLS9fXVi1zQ7ZvXT2CwpBSf8I2lGJzyoCZirL8Ds3OD1SQHfaFla
PFNcxKD+00QImez6zT3p02qHC88blHl2h1bQGylFCzu9Vk1GMQq8/Esg/3MlZG9U
YInHu+WHfwl7PRieTnNEbTNEsK/3fjdlnlfywnAXgfcTANL0KD+QloK8C3vEeeZE
0+rsG/JjXHRJPbGwGTh67NRLCoObmhJ6cvQJjVHPCXMRtmwLPacZnJTF+qDu2wLG
wfNOcvFaP1QOrquslJAGZs/o9s8CJNbAauPd6mA2g/FzDexd0VbtI1kW5PNMH5kQ
tKhliTMYLwdArWTQZjpqORp2YnNLiNMVybEzhbU8xKxvs546Nr2LdldCV6LB+oGk
VBWiqXF6uoAp7UT/IWJHMpwkBCgX5P4iGzMeJm7n3+mH01BAHutMHmHSXnFP+ZZf
A1LKB1gexT8KsqV4c12z4d7P6E3BSwahzO8wI7VqG2M7fwmzloj0eKafHYTpBs2u
suyEc8TYLCDVN14CY/oGHNb1DAxkXErRfhPF+ARTzjIlX80E+VrAAfD5wpu/9ItK
89Mszk+DW6zqj1wkY2nI6u3ny7RN7jVUz1HWarp9q74Qk3zl3hUYYQ3T1vD6lbgZ
+NvoMRPlKHvml04sQ03BUgEZgOvidDz0zQHcdzT57mOZQTw4SRaX3Egw7vVNyhTi
cMDNTZ129gqIpES9WEiFYNbIlVJH+8Lcmt9ptscwG0Tuvkn8XrlhC7reS8xvavEj
3Cz2axngCVDfNJimnw13FOH1KqpvvBLGeakxlcgNHSU4hIdNpGlXHsMGaYEEDbI9
sl4FftOgNop31oRzBeitvZihjuuGHC5maSArubcKa0y7us7dYdfHvTAXmq8heJqV
lKWd3Dw6khe9x0Gwq5iWONqCZ6rbLtEGlI/zC5RXcYbwm+zAwPBN6iKOYxRVaHLx
gaWh4dBXWpdewSwsGIvRiBGvrJNPFbnvT7/pkjnxyDpI3ZQB/Uhlqz39GyYIaoDh
UoceSm5dOqvEvi7L/Y2T4s2x9q527PSDZ3V/xDumYIc0cAgEniPRdY+4eMWXkTCR
4odXC6Hu6Fd3Ayg6pjsYckg6Pttljv2oZrIBjFdQ1yx8+B9q79hqU+5i8IVuANyr
UWw2+6DCrBuPe3pvIgtqbVEEJPNG+f1X8Ovo4ItLTrA5b+HNOcB3Nb/L0Iv+886O
/dXILaaKUrJd9cukOFxunfBWWEKVikxX1YmUyGCrcIGneHTozgikQN1d4Ew8Q7Wb
jYRRlVHYB/V9h0o6jWmWr6Ykp24P6N76k/049Lto8S4J5TeFYNFqzdkYPnCl2BE5
3fNGHNQtqm9QDvm8mZ6dFox4fAk9EVvAVB48cbxXLTNpp1WhQn7hkSpwhccu+gHq
t92ddoTQSbGLJh8xTz7yWXk66H0Yu+yME7MB33nT5jeRfwnoJ6TLtRMVmX88dMfP
ZQxya/B7rKrQr4SNgZzqCmfGt3i/2EM8+4S7+cdxWUfhF7cnUqKubD+ZB0opExVH
E4VNsQKAaz+Y4rg0FzhgJdJlvulqeg+rKQdRuf1pumSl6Q85mOSKC3p4lLlAEIPo
bGlho2rWFWnS5bRqiMrNI3O5ECVX8oD5pNMy8bJBg86Ee0Io7pQp3n5IxSVmM0UK
EmXPOyWpyAhOPo2YJmFgJD1nrKIQCf6QN/GVoD5s7voSrHlkJ25l+ItiQXAXgKfa
JYZbTm3aNKUplG3G/qOJAcGwhjEblu9HdZY/p31BQUjSQKZbSLMFzCO2BrW9dygN
laBTn1uLuHlesWRrh8LI1CcmqZpXP3b6Kq4LMKr61P8g4rgoztbRADzoPDPt+1HG
eOh7b6PGh40AkbWXwJs3eHQ7yQYUB4UoN8sQV3QM8eGzCtI9/xxQIlPHN+YSibYN
33tnqJxkaQ+ofRu5iq6qJ1CYpuE7aN4Y8IK/cbMx259omVjoi6dQfRh6LMnXeuHt
yB/tnkMU9TEk78gU+jyLLF6niJKJcP4dQFRbOGyTx7TSB+zDjTLpQKmAIAwDOTU+
aC3iwZSyuOn6SxSSQsfOLi/PSG/9IblpEnzwB73hfBUobbNCYICNjKIV5DJOlFoh
ZZ7keh43uJat558RF8w1m6TWa70DQ7eqP0szPgp0JGWSUsGvIPODu1bEBlZpyK6W
nWbXCwcOlokA+D+j4FOC7Gt1QRAI3PaFrl+bNIbPbION0kxvJ09YFs3C1h/4X9S0
aLfBxxD7sVQTvV281+vT4Yo7yVQddkSxKZMmHyDDhskIE7FVHlFhyYTGlg/HuLbL
w21TZAzz63YWckFbVY07+yUBwOB8pYUmZoGdjH++eRkyRsg9qE28Z+8oKgkncR91
9U+7zTDQXZSAi+xaDqjkeRxVUq0/fkBarW5z9DHhPW0aL6TyIYBS8RzBqKuiIOE9
1fN46cwkmieBbJ077cA5TeYUbmv+VVmjWUcVAVHQcPF9n/9PTWieQDFygXW4GMJD
XaPO++Z/WQFiCXu/nt5zbjBOTwBTA/2dPQLiYIbnQbnYp2Fxg65JiYq7n4uZ/0v8
KFiBEFy+57YbpEQg/GJSTMefjpgctXSDP9oZvXeCRIZv25r0NgYJVlkXSR+d37NL
ze4VH4kjKvwPQFWDToiri6snQsTgRnfrF05KpIEWYVXO2toIzvLuShD6+Fr7hMCA
zGwKPdp/eK/f7E9J2kFELHnCVsBgDc/ybvs6FBr4KNGUT1l7qHOwPfYwS9x5r8Qt
IqGXozSX7hlfISwe955YbWn8y/Lb4VOx3xGngbPaxSzWm4KhGzUCsj+XU9ODsrVr
aTt7i8kU1yVWfn96LSfXtTMncY1mdC4DMO6mB/I3vPljC8Bd00VJWOdxmHkn0Qpn
0R+V7RoeQ2BQik4DVR+2NLPdkrbLDbBx56pVpV1BtoQVXMcjfFC1jeS3fs8lirG1
9v5MRW5BDGv2ykuwUZ2bz5At9ZQ2KziG1vr+Z6I7DV/OOFOZ1w1HzP+MmEVNGvJs
qF9zzjfpGdeQnvtBd4dcXF+waG5TZz2ZsKtTjGgtahC2Cfhi6ge/8ZRvxJnhPwT9
3QHOTp+Lz2FQOhjBilM1V5iUm8PFWR8nbEnMil1o1WFL01DkyJyvFo/V26DGL3Zu
xAwHttRoNls9WInVbMaVkxy6jY+zi4MpPTlU0JUYMf013BqkHyQvSAjuKfPfxQHY
CbOxpj36yojXuZtR9EUXza3/35Sx0khLVW8uYy7BpU+1POmGZgZyNsqxvJoD6gUv
C0fQ6PxqI3Lpg9Mwsy7ygWX+iFYE+4Y2oQSv+xvPnjNcqpsqdKu26lx566KN8PqW
//lP4jNTRyze9ppLOR794DOqtZrP6x19W0WE5Nwt/UdEHZxCeb/KjlO52BcnkiAm
UTvar/yiMaRsDgL9cjsyhn0e79VXFzt3xeS8hkcBEvwGJ7HeFHejRkZLeeY41Wiz
1Opzni+xjdv3ZsrNC4hBzxZWNNb6URnLZN/+bviTNEaq40DStRk8+mIZFnM2oMjy
j+L+sNtUN0gdmTqyYEzQjitSV9cmP59wjY34Wtn9O33fhQqA2eX69xAmtbjiH2eN
gPpzL9ARcNczrjq/1PX4k3d/UbvwXwLRHj7WbN+TLqZPgrStGDqPK2mP34PM+sSc
vKeTuGPeQF/n/UKSmQlWneEnOZLQfDYhUJ7cnc7W6QhWBzArLQwIzeQBCPq6od53
ugq3bETOCD4a6yZAwVow0Gsr7I6p7NphqhWUYM9N2XMLYvEZEoBmyeEYeba/z9Dd
BvYuoGmM+v7FlUtFL5zjhPzbtXPfQ/yCnANj/w9Zqhw9I5I09T0njmxPuh/gOmGy
H2ovf7aX+ChIMvYymCKEIf5mn+o524ylY1tIGsGQFirWMpqZyD4qrQrk+FmgbA71
OCN2WHEZOy6RJud5eukQ/t1qJTwr8yMGngdHLE7doMsmjevmHzgDOnYMdVvXj3bi
EB97njwnaSE4geJLicw7xU907NMJ4e4b3ninK9mHaQ97S6bXwUarvip/MXIL1Ach
AVijcnAd3RdLGggWk3+BDXAoroe/VF6qQ5Bh0FuxJjr/OHNzjpXT+7894XQ1r65I
7yDo2hlbe85IYGsSX7mCBEJrLSHGGDlAHOuNGgjKclbBgdF9iBNXB5+B+BlrTS09
R64ZA1CUHmngABxBmCQRIG2m9McorVAmV0S1XjjDH0bL/7j/XaFmk9KygaJahMhr
u4rfwhT61SE8S7KIUBML1wYnsGstJh/jM9bF3vZVEAbqr/enro9RctQ+nDYMQtRR
/uJscNViEIocyc8taQVNpXzMkk8C+WValMY81x17qtsNt8AlxRYj6Fu7XWfdunbk
zgq7uVn3GPG77rJsAi32jeAwMUUvJnLtxjVNo0XZuhCgT9abH1OCpGwLCWNX+P2X
z4Su97xYuvIWQwdAPxyxRhFmcly3IvL7ZDkzamoWBamwWQ18GX75qte4QF8gr4Vk
zU8PHQLGSwcOmP57CJfOTxRBhJVqb/1GntFihe50UXuaVwhDyDElUSWxjegcZbvh
x8wF0tTtkBqkxHeBaxYcUkzT6rPfBb3FFBhMMNLm1qAVrBWCNQ+fK40NE2jq5zXI
UOC9Mx5GH8lF+djCfP0ETBm9gRz13UKBMcWwTjFDi1Fb14gdRFU/QnGD0uysihrS
GOyqFcjrBcL83SVpVE43YJOHjYH8In9op63S6wrVnimRs2L6sapD6Mm8CkDznl+L
2tBgivIfYVKn+3vfE8AduLWtSN69fuRZweCG4DySqGxXBdV0OgoI+lDpYuWR5x8X
PQTIXB7N82xsw68BVSYs6cR79eVM/5np7jcj0tj5zLNpBarBGFrPokAT44PCd22q
AziTGSlDMps6/HPA/UqTzF0uW4IYXyVhOUZYqSuJ3ahoZozSqeyvf6O9SANIuSZc
ddPndgTyw3K+2HIA48pxULiVtffjQYejpP+oVixNS1CnO9ZsGr2tnFyJp8aBmqpo
tEw8wvYBW7nlgRbdwj2qBpbjeclqEttZ7x23yhAgX+pn1TQqirCSrxOGRVWPYH71
GFN3JsKmTkccpItJM9mFfm6Glwq7hQ4ZNC0sPI8QclVV9yXytGlTlktM7jGyXk0w
8avVJcY3tsEfCpgRyQg6TOQ5smMbqg8K+E/7JvlTo/DsBq67adRZsA32OwqBYPe7
X2kMcbkQn7xdOseFBtOgR0i5eTtODFpaguVa/rUoKIIuy9zvZS09bDStpzKJMsMC
gUQFTGzj3l/xtKbE0lF+9SLKZ1HK4voCxN5+bmcLHh46SPR5nPb4TRrO4Aojfb0A
9WialvWcYqA4R1PKupKu+Bc1JhwK5qv+9r5aJwadU9y2xBSGL+nK1P7/KXnJxhtT
+PV7ubv8k5EaqDQ0vJ0qu+CZO5MBPLaaBEij1g7x7wbU6qzTnYvxksE7pzKrqKhD
VsazUh02qv52txpwQKexIpU83Txr2tTTSJHcxpspfsTymBK8ug1IMgRayEhs3vws
gJoZgN2uxUMfdm4TMzEdpqv3Spf67uLEqxj3sat2/JJzLiaPDAluFvmDv6NtMOKO
v4pWENhK3ddn3VYn8AnOobsCVh79C8B+AfgluVkp9qJqBlub+floSWMdxx/Jhs8X
GM1fzPuaJ2NWU40z/LvIsx2K2w/u7Vyu+Qc5qgk6HPnnCMf0QpyvSLC0i3hlQuVI
owlIZ8JII++w9gPUSxKwsoincj6uZqWE2S0aoHkXX7OgOp/EO/SFtujiPJES7g9d
W4w7pfa5QpP5jE56/P7Cvv+ZpikxwAxXJCCscNBHEBtONuXOna4humVVspSyGqX8
tDyAZYdrH5lZmcJ9VIThZxY6+Tuf5Z3N1HULNna7/TBKIF99H4ojcWJ11yJ7+1hi
BrtwNHzO9ZZ+qVl82dIPSJHWBUQQ1TobWsalfzmLksKUYxm04L/p5fQXK40IIB0w
V5YLXORTkKDPpd7UDxpC5ZWZQJs2t5M+2GctKbLHtpliuVTHQyhs7psoOFA8YrdU
aKNeZgSCaPuCRrjb3FFcMK5BW6cDj6ZZwcxEzD31tqfOHcgRymZIJpzXwG7ticWJ
oij7uwJrPkYUvDOfI2YyK0CevYb172S6+rbAne+WxJ/0v7AeP8kfoZ5l5x6xpb6O
4SzTOwwE4F/Sa09abxwte4nEOw70LWYuL/0b6RFvhcbMT1VD776r3muRtxCWodmM
MvZw5MKXviCehYGmgUDVkjx3lWBjrOEq4Bz3Qc0dZMjOxLL+hqF9wIHKn7NGRoU6
81jcIMmRHjpMJqxIm597TKdAcTqfmhQ1ZN/+R2t5ngAcZdfZuhlVQhFnNl5r2B1E
y6qf11EzOKkm/0fp0S8/J7+kYN2QSEbahmqm9p2Od62yp6Iwx47r7uywo/o34tC0
o/tUeJ4tSO1rLVYX5p3dKFLJPmzCDljWZlMA4vxo1neVQh0asgbDcmgv6uk2BTrI
jQ/SAzXlXOsdx8ycubDZxCOPNvrDPmC1oTuHtQSwV+F5qrqSBv9jtTnHntSMQlNI
gaypb4d5MDrrogROdz1kPYHEPWMA2dipIBLJs8T8MH+qrPp/JoQe8FeiA4VlIVFS
jv54rVGUT/x6lx+xAvYTUjdKYP4lbCiOb4XVfzQzvqXGBz5Z7/+gC3LQct3iwcvi
doRL4MZ9Kp+0fMukJUzcICZ2s6lG/z8lJXXzWJBHtZg8qotErAtPpN9F/ITmi1aB
9xymxtxHxDfOx/2rBKnGnXOc97+x+1ggN501csTvIcy4PXHVX53SA4HhS5DdFpcd
y1f/pwOOUpwds5YBYC58dIhr1Hs2T4U+roFDDbuDOaOqQXthOOsh3fRKBMx7A6Of
s1+fVc3M7pvR5d64DW5s2cAmK7YuuFBs5dyhC2Wsep7/JA2+L5e8YeKGrZLKN5N2
zdUIwHFtiXCc39GJiifDWgaxZvW6ob/Mzue7KXBofCPW+hQgRm7owchl2A3E4mIq
ipDuJwj65w2RKBHHMkqOmlunXet4lBGoTQR1cgqOJfXnC7ps3x/R4ltvDLqLuuN3
8d5vkMqJ8tuA0pz4i5KJxnlWH7ivAam2VHk16EQVUU9LD0MDy8/uEsfBY67u9QoR
73gmosELxJMA+tI+TMmztWRTjHD5TuhGRkZNwLKH2O1ydXwFxORzMMTYIaeqlgDU
luy1kiifx3Bwt1ip3A9n0XfB9QSAEga2yN6VZHYxRHpOOMe927ugIUTTxZGNt5M9
wDqN20Wf0IApCtn5HSTeUFc5dtfVAS7cm1wXXo2ZEOE96zet8tnaSl7+Xe5ETaj6
GqNLOXWgEU9xGoKCZLxAKkQpeBrG3dauBL8FJM7VlnIohdjNOOU86chg6u7MjEM8
9GnQwSVtlOaYDClWn2bAnCSuE2uf7Nv2b49aGBI/p0/1M4LlSKOAoGZVBzKGOX5I
DeZ5JkstAmmlmWclyPwNXUklTXxpG5O3Mf6Q1gNUt3LJ1hXktAneXbTrpP7fg3YC
yX7HnIEagoF5O6Pp+Gmrz9sxiSHEG5MobK23tNQyRE+hrDXsbUVpCRoMDAiQloA+
21y3b+fkQHrRYhEsPKBwQWWpbCGB0Yq24wpmP5f32m2KnBX3or+ENbQ5c36raSuT
/Qpg0UP5QIuSPcLYe+WPVLLWB67ArGe8mSLo1ela0KULksxq+l3lyOGfC3TjWgWp
jD9kHjXPwOEl2PQSJcvFwLzm9AbVXC2yL2VfirWT0UI0e410paK8HOkj0Iy11ROt
W4WwAW58VoGpTvprFU8Vl9mCl8XmmdXKCi14bzUCWbbxMhBlE0uXRLljX6oGmaSg
21BVJvc4kwVmxCP2dzKGS/yg4tzvrgJ8jhUuK4hCZXi62chvwGx03hKyg4B7qPVy
thaK+pnT2X9cbufKCVKWEHhn9CTHWPaHdVI0E6nSz7sCtw6/tZerASItZHu6xBtC
OE3fOoWJi8Yfs5MO6zsc2qoAoDZtl5tUDBjFvFNLH6YA24cBf+7HPdInnoDQqE90
Y30SY06UsEPh1dLUNFweLeUuOT41bxZZwDsWECROQwDHP6+XbQZUxie1JWv07hLt
4HMEDFahBhRPCpt2/hY7rjkxN7ZtmQURUIq/6OwBZGrWWmBSnq4SKLpd5F5L8u0q
wRMQHysduN6EF+LPQSxg+6SqovaMznn+3p2233j6yg4Jvp+zMev80x9Q/4DoGkya
Of0zT67fF0LZ55OWOS2yTJC/28MjFB+7+gynmgprbImTVVhqdvzjI0+L9V1xJpic
A/EnDsmQprUVoz+yv48DjM9yX8edRMwnUAXvwIckRfjAq9jd9+uprTPSWf5nXH4T
bZFP78Ofnx1nsGzYOv3peYE5wSQAh4q8+wO8EzVfP47qoYMGHhWPZqJNcOAyfs9V
1UIbyr3K4QLiDgoG3oi3T7+fjptxQHmu/gx1gfn5sW6vEmcEvoBY3J5qirwXUH8V
drqNtK3luQsRKTYLn0nnOn8hxn1bJTY6t+OWCK+nXuOSeFyqWyNKxCHybtb/tibC
S+LMwXv+KNqdGfrWqpdB+LUsLdX8R9mWAiIvz2k4NcbRgc3IGDCSi4DEhCuP5UDA
DoSsXagiHzW7kEHTi4RQc6GLAf8Rs8UzqKUGsnhGDxFdykpoDvD5vJ9KdhW8ThBG
ibWlVOaFUhOc0Qa+fNzZPymhhWeqTpUoQV2xeJfJDn1qKbk+OJrY7PCKoYtFaY+E
h87p8aWWlkFwIQ37xcs/rWfsggSYbEjBQgSsgZ4Lgnz7S+NAD5AMlkHUuSaqK+R0
van24a7kGFSeOhaw2DUCNgC10iN396zDi46iLwBWGB1C0+jXrCq2muJZBxNgbHHw
KjcZNDzcnhESCCyxQ+8Crooq17HYd5kpIuDcAy1IeuEhPRFxsa0i4qdjD60MSZVr
cNnv92JOLy0ZjWMHmGgy1ufiJPaBY+j6v9apoYrVHQ/c4hVOIjxG1OdKMwshJqCc
NJhMCxqXGrdgEzYdtVfe7gFONYynkBHTBnwdXRAJhaN3waJBiR0avk9cAQ4GMPov
l8kuiCGDSAEShjOKAXuzP8lMMy8zkNLXRV/898smnErvYTS5FfPVBnA+DmSqzBvB
tuXMvhbpciF+53O2fTOBXw9Szp1xXvw0zugyIjel9UpzaYi0pHQtJcvTelw2vKvM
Pbyi9fJ0sb9bWvLwljPQFXvkPyI9PEO3qhShkwIW+83uoDWyKS3UxQWFYPc6/89W
5iPJIlMoojB5BTKCJk++KbBtBSK5y+8LwaxyYfj4ria5ivRJWZCaiITD0C93A2Zl
DNohLNt4o5k1Ejys1VoeLkzyXisfjo9juKHUGtJBUsA+15jEZJAhf55Av+i2D+1Y
TrGTM1h8BUyME3tXgZfRqO+QbXPRmz990f4x7Y8XzsbsVSaaBLo5BQnWU6eBlLO5
ytjQTbvNf38UkVj4RY5QOQlgmycPVIThaJnZ6x4NLWXsVgvZckFJniaqo9QpaR4y
g/KUvS/3RQu5QOCHHEFe1u8LGHMXGyQR7n8OmqNPWoKmi2DfUo7Zu7ag5YDQWFQb
d1yykcWp1kXGshEqowhPbsqadD1mzwo4Ip/NzH9umRIgrK2DS6OvACdVkcet8ofl
erckZhZ4n/doScFPIACFy2uCP/h/yHX0+ytT4JlBs8OKJQzSeZffPwZSPErG7RZx
92p1Kcx9YKoWkmPNjsKeSfc3kfzjdGTfjuTFU/g3JMTbQuhp3OEeS8K78cBeca3h
iDigx5jdACN8jwsvoPGTEwDranQh7cGEooeZoDU4mSojeJ7ahJDZrauammrqodZc
kG2v0p8aPH9y2Qa7XxfGuen6HaLjiP0g4FlGOlA0B6aps5yrV9ZfhVPgxKO9nCiq
M2kfPwFp1YAHSlSjNGhIBSxm2FSO/9uRx0j3MDJm60o3Ko6j1nCw+aYlGi0qJyqu
99FgtvcYfsw703Fcia7MrlJFW+S0e2MnTybDXGilSvU4EG4bulcZvRrRIjMQFAsJ
TEcsp4l+j3hkwMLHo3iNCQ3JVJTyqDACTuCDamoHSWbMpQ38mi6Z1cSZTqrgIior
UrP5zPb0uVAEknMUug88FUr5i90hspDESk4fg3T+NQTAVS3k1a+7Nv45NjIMu/hV
22IHpjnSlhub9YWRXDkyd2xMXgsZKtoP+7BJmCA61PLRHw0TrMLMxa3yYUbnOsVf
1/w7Q/1Dw9cBxv+RXgLyT8FvnPAms8Hzx9HTopHJTGa2NwaC4xryXH1C9svKE2A3
rsxlmys88wJvouEKL2zehzeLnK+2rHsqIfEUZINJezy0UGe/7fN64leUzPhJXZju
/aP9ex6lAoXlPt7fkiBDnSSnap4u7qvGWyB/eOZO1i7DPI9e6dfMoKCHFflwBDzU
zKloMtApxQmwXWfmQyGjzQ/p3hdGq/ykZspBcpo/JR08hGYcvm4pBoDQ+si7ptas
WHC/b1JofaXQ29Kt1/3nQzdYTUeLZei8srR0pegU47n2PoG1VYbRhmxKcdK/Wne2
A6dJmA+bQ7mVkjdG5zsaGjXgi8YF63mpLBk/o2jOJyx7/GIbXArfl3gqnX5WZC1b
W/CPNOXVFUIgRTgzVnpjrZEoSQxZBkPPlzkRQNSHM3eufnr69rrus+YWt5R3kT2i
LMUpeiKt6nY710m1i4oLPccBIwyZC77L20GXV8e6RQ4oJeLQvpQcCelSqBgBNfSH
RPT05bxVRWtWyet4b+p3NPr5kv3gJRPHSPodZeWWEkjvkILHC+Ohp6vdcvP57cqY
/oSOPC81CDYgKzkydUmkvLgJ0gCGOI5EMf+tk5Eom0VhFJtgdJsrpVBTFOO4dGUr
Qi1RHY2L4FLnzAgniDMjMS+NCkYtguQ+tUCMDY+2Ant8oAvMzUIVElW546vdn8jf
Vpt6GsCpLQgweEr6sTm/VDsI0tF15ieyYaHd8HNDEziFtIVLWxWwc9X8Vo6DtNEy
F+/1wdk/CCYAmNOu90LjBr63KUu1ay9bahxpxzgGe+vLTn3pv7w3ugysqwnocyf7
NpeVNZ7UIdgFAGeoqyNDs0wqW9L1skzVsA7kuceU5WaWKDwnhp0urnyrjYVHjnet
I8h9jI+csUvVVY6UVMfcc2tgRVZyzPafywL2VbO8CKRoq71o2F2s48/8UYTR6V2q
z7CqpDxCI1zmyft0QitsXrhy+N42gucCyNjfue/pW/3VvEJPcTAE9MYFD7qmDGDi
oXNw1n4fFaawhZyHg04Jz7BkJzJZWpBY7Fu1lHX8Smop/PGoJCcYihFheemLlWZH
GCANdvDo4Dz6rrH3aNwhjKDrq20Z34n48NpHTUmoASQ92yUJqCJIHY3gU7+x1d/h
+Fn3ELaEwu9+U0idvk5gm0xaCBaPuZaSyEl6DRn/lDdbaemuu2pthBeFAT/g3+Og
K2WzH1nOkM8GjQCU3GmxTUYk92N0Wli7pfk5MxBKZeJwKhDcciElKmORdKIVIzsO
kRZ65C63rNB3YBxyqBlUGRvf1HcrzZ4h2kxpghWIQ6lf0dTgXNx89mOuR6GHenmc
lBHVJNd/8TOhLbCvPf72KAW2JrRI8qY1+nuszoEZRjf1liaZEBGdzvQGUNwD8ZF0
0zacXyTJe8lGy3UVYzVkFa2AFI4+qXbmowkPyptooIzG6us5yobxKnAuc/ay8efo
prvYr4GSmhUGj015QV4XF2VooYeyFnJEK/70BsKuWvfq8LJSIB5ZwWeROLRSk4Mg
0WPyplOkswqnhN03goEGhD5T3hg0aJOkor2A4cmnvG7oh98XE6nIfC/kBRm9whsk
5Psoq25LpFMtxOfhvDlSYNGk8U6jK7bhfthnMN5p2ohsXvI5Ietnlt1bEUsIFU2C
NspvDIeUXuCXgTf0Q8Um8bjo4eXjI3fzJzHP6nFhZ9+A+qtyZZcpR+4e8FsyWN5Y
iosC6vHgdif9Lufoo4TiOvO/xlzaxpDP3nBBP76S4gZxJvx2Mi9qGcosLBAy0PnN
aVRpQC097boMw2n7/mCW3rQqmojWVcoHrkjTS1ZXT6yCwlgMoV1uqtZ7/y9AaWYp
T1cmuNb/rucHyqKS0eVHot7zxiwupg8/O247OvczE71N3G6HvV3asEQwkEInFo5O
scnFKymWo9HkCDzXlMfTDKSxL1qHexbj/WXuvoyfxxoWdqOZpwQ4SqVh5868Bxle
lwJrgNblq6Cw98A83la0j2SCqwMMLQvv35otSL6ijNIjUnnuRnhgdT2s2VGxWLC8
KX1aUwKdf8fBG2sZ4ZQRMDb5SL5CvSs8+A8m8Lx6IOT9N6ZSarXxTHMlmqEhXDiX
p31t75pzAMYRldyYWCgWUy4IGlWPC4SIzmMqQBZJZsgriTiHtXAnU85S+8wz6sQ5
cdM8tDiJ7yS6zekItp19SX36sz2fBRHpuMUF5x6BQJ3YBhhVrEt/3ZWVVpfpVjl2
TRXnyszXIJqoub0GAm11YNqMWbBm6294ZvwlZVnIflR1MMiWoicgpfJIKz/fy9Nk
P4sOniXVJ7wAX9eWoHUHueYglFjUZPh5xush6FruZ6cXCTxPxkLTz+qrfHSl/tsP
ENtbRm6tsQNIKFTWwVIn2oeSGGpytFlgE1Pf/fF65AwzjXnCRZ0nUsRcPfsxXGY4
i6Iym566UB5LXEo8SY5M5KZv/A0AywLHEITrfjNZ4j2oyqYGKYVQ6eNHJxwbPJ+U
wFVvKGiaUQ3LsiHvbPA6Y4miArBs82x/56BO6RzeyWXC0u1HQdJuA9/oeJEjHvYy
z0w1ybqkgE+0MxhSqZde2s1GYX9uHw1tAoGSAmSDXJBOtEYKohIKjYFz+icg8a3r
pB5XEng7nA+1iqUr6Aj0R8JG0sHIpAclDejqqpwO64RpNwOPwjdT6QQ5cKCniMq5
n4CKbmbdLNFk/NcKF5t6NnnfKWuTt+b5tYooDDOLlZ4SnYG4SVqSAePaEIK9rqoN
47eOSvl0Yysks2Br3/2OfYaPaopWexHAA6k7SLvVGXpzwt1W40jAAl7W87SpNHDD
7OzHVDKxVz5Z/jmdMklJRos9Y0XfNNHKro7eo1hTh++/QMgfzn0t/hpOqz/sLy3X
OPTib1HY7tFFnhTcfN612Yv55XHasmT5SCW01EzWr3rcLu84/Ca2X4b1j0S5pyxV
gL1PdPYNEVkx/IEj6NnoeNKPDfA4jiTyT12eYjCoWkGQ6nOkLdqtS86eso3fs624
0EzCv7vM3A+sa+NXL9oyLe2cWgRgb640AVM9jWpDdxEcYr9WZiu9NqaTJx9t2a2F
Vw6G7y1LdadKlGZvAYYw8W2Rz3xpwqpZPbnTSPHlv8CoJ7+mXmGR7pQgZ0Ld6r7Q
Z8aHdzRvtd4agvrymuDz6JpzBQk2BS/NVVQqMkAu95Fcy/hCpJ8wPpJl/Hz4AmBI
x7BvFwt6KfIIMy1ftWu2zVUyj+0+7VSUqjqrUX1RV5FQ0NG2S+L9r/0jKQGST/s2
TzBZQZYj9WRKugR61Fw8lbCfToZDWFFJp62pUIelFq6P2wlPBC7gv6OrolxKLGw9
5ZupzdNMMRdTL+NQosypI4UAT3apY1210+KJinceIEdm1yC/j8Mi621MDD+ZvpOW
eRY5Z52+Mw7J7mTSDH/coXKdQHh7ktjsatFEIjCZmiKp5mY4NgjmvY/Joma1epA5
od/yLYo81qkTMkb4qyN7kjsZpXYxMoyB86lScMM85W9QTDMshTPer1YvtNxxsYrh
Qaru0xpUEOIV7Z4PptdXxyQmuORN5Strj7D067vxLkRvtS690fINgEc0SQGja1Uh
ebjmhb5xa8FEj4HqbORikDS1RyLcfYZU5Dn8ODDBk4GG2SkCjHDTya+qzScAUsJT
WGL3gpX+u2y7VxfAPiMXZ/WNAcBnKZUjAICg9Z1BAPEg22206Obf+BvnIkRImDhj
SbWWg6zW3eTYzKbow1DH4bYOStFLSlZka54d04A0dnSl2/RHHaf42o151Cp+iA87
nQiFTGcXMsEoh68/clr1llJFzXOsCJE3BWVTyJCzShJdMPMgIyKmYbM7c3VYHqZ4
nWTopNg6eV2hcUVkTBRaxKi7KASeP3NGmFkQgU/31iqowoeOW1S/dJR7B5DjxDVE
loqf1FLEfB1lsGBybtqYbsMkjdAXJuWjFB4iOO46zEvDl6lOx5vqVprxtzfLkPSr
vARtQF/LTWfDHwGkbLpISrIqAnyUNHn7HmY/NcoTPRAXCbWIBanrOTKE6PpoGoRo
wsJwB3Ba8EPEM/MddsU5wFPd/eNG+0zaGOdzU2FvznqkHDy+oUVP2NwVTq1Pz3O2
07PSVL1s6m8erZUytBpXpg9NUwODqKtUpGVIlNst2hpLBS66DE1EyFMlzfmy2Bnk
jSI4r+Kr17PzUg6Q8mjBbsDQi7kxt6eFYRAWb4RMKYvLLM5/XRcLcUSkLMAIRGzk
0dWpDU7/8bEBW8TlRc3LZxTQM6b6A1QLkah3RU1cqAm4a6um25rhJiXyBGQ/wT4k
wUanQps5ZqCxREjCo4JfTm9iSdNUXXfII23br9Ka+LkmSR6g4iZ77vlU+b99me64
sb3vC3OYJPqZfylEoq9yGF8oT50l5KWXY0RE32Bwk5TdHIVedfx6XqjDa8Ac5pms
GMJ27ptdzYDMEqLInJ1MlZNwledB7ghNL3LUK0/cV15mKHdPl3QLunWc7OM4e3di
UDYXy5L/RiHx1+aNinm/cfZSjh6dUgpbtQjDbOD8YDVFX5rL3OCusWBPJZbX+pnF
Y9hojG/6gxVYyfRgM6uF9bv1mGW6L8OM21EtxTkVilXTIvm5xlISqMx6fQer0c6R
E6yAGE6DElh99la5Vd0e5XIpliHnDWUMc3FznQqokT6hqOMwVcyNMGcrRHmsa06X
XKJV7g49Kv2YyCeQla711k0/53RHJA+o8KK4CPfOE+siRh5U8q7CsPWuvPM8R4MK
36uX9WeyxPk57Wa18jwSuU3tlcYABLYNrP31Le5J7Bx+EPzOo1/LMYep7YOEk6dM
YRqeyvYIfi9Y2Yu4OwCGKDEyN0kBsaRaXdxVj/D/qpKsIBmZ9l0M07QMdbxxnRBN
i4+FWAzyVlivXUbO2dYMf3WHUfGsqTLpG0yqcmVqA4c8SBgQqBHtOqHItWnp8to/
eZKm6a6LvzB2fei36xBX3f4UZne5HU48rvrUBkDgaCvr3ZvDAT7o4slBBaal3YZl
K0/6LTd+F6czErHmPdhnJeVMXqzE1VaExNWa6FqcJa4zRW8b5ZpuftKQEvsUva4b
BcbkSO/H0oWwfXNDaBiqBy1P/+bsDD1CcGYXTQg7G03DjpPu+w1QTdqk4GnCXbll
6W4TbJYGdBMrQy6sVaCX86Cf+FiI+j6/yYv3Gv9PO/h4M/6NwRiHqR7pnEwkDt1y
TPnhXr4+a9rcL8/9myczkA6SGmO6lWrBTvyyx6JGn5tzyJABKuSlk9EdC0nXHHzr
MED2eCqiF7VvN2k6HJvoNd/eNwzv2ZuaxDfKJGyUITQrMCxPVUKh7tR0dFm2c4Me
8RYRPJCpdYP+pLAeikZ28fcH89GkcmW2CMmnM5YBPrFas4tfNxLYrqRJjmccfbqk
aq1VaLF+zVauvSdaAO054/2W76pDA8JPuqdAYgLJFRt4MD9ylMUeDnqhkSd5egvi
dHVD6qFMQThT3S/W+oB+uY2o+8CeAYEMGgJ8sEbbjaiCCNhrFXoWk6L9b3Aw3Sik
+vQkq7ro1z+KaGXQp77C3GrakUkfRHBByPnl9pyQYD+ESS33ceW0rdCK4Xhc22hi
5v+bjlSt81RxokbSTHDuBtvHGfDEm4c7wVxmIYhEtX9RQGH+GnLJUWee74eiuqwL
nzfVmYWiFhDC25/gDMotQ8HYeYe/sYEEGiRuSs4aVDX8Cz6h+orb755wMltPFF9b
tdcMTFgd9ITTr6Vb0Ka1lRS3auxtea3wXvfxXZItjhBQFNR8K4742aM8YFBBxqqf
2MuWvwiYmmO/siZqtraE911y5DQ/WROZiKaTYJbNpdMZ9VkyBFhoWKmIcEjv07mW
wK83nIKlR8O6gVMEXAGzaMIxM0gOej+vCwkUTkse0YLItDGEp+UBP8TiPr0LT0Jr
SpJ6TGkPW7NaB31Od9yl41JH0B9UaIJJCi3d/xY7mWhw7wk/ExHNI41vVD8sn+H9
cOHHGFLRNFMJvQl1zCjq+W0BPYDOCwFB0WfU+vfVPfF/ICHJHPhzZ3HqYq0ZsaUs
5k7K7R/GqcomM1eBLb8JkdfVYCRwdGNVabxowa7IJ/MGoAXNWUS4Gvp0KeOjogK5
Vpb6cQKcu3DCZEVGGguWDDP5bgfIamRbQl337AQtJPVE18ea1f4Pj50GLuI+r+RO
92EUFw2uIeuUdbqhL7rQDHLt3b7WYpMTtoRnT12S5XJZFEbwQPXgHhAZp/7OB6/m
bEc1konF+yersNSyYPd9nDNpzpAL45oFArw6OimOy0SS//ErEtfXHgSOM8nbUTTJ
77QI1OUUrEKlHj2ox7eWL4/9AWUVSvLQ9VWoSuFzjWEMsA6mUQiT1OxxBga56sPY
dffIPIWVHplVavan0TpHpp7ShwJykVUz1S1dOYnlZN1xppBrUFcIXE/Zboi0P2uL
IJSg2jMn7VkVP1gQhv2Ulv59LJ7IPH7EiV8wr6rm0oRQ0wzMGihLQo/NF291h9mJ
GXT4YR/JB/RuFMq3S22fvc+5xTDngHMX81R0qzmbNvPvFHzffjDu51E0TQzFyqBx
YcqPKEqbLrmzBK78pQIwe2wA+l732OB7VMtv2m6bi6xSwv4l0SDzaVvrqDmokONP
DGM2cNjq/YVrp6505WGOjwlEXY2wDHJiAK6+qgBIVxgB+roAjnjku6c8d6SM3/5u
Dvw4YRm3ZbanqARg6PCedprv6kSMTOzSaVO1clm6Sx5NrbCqF5NuNxFaFewwopid
cMMmFSKJpJgA+ny0/UhhnWk07S4IUwHLmAv6C23xS6VtgT+a1l7Qgx163alHH+WY
MdbapbAHqFMDBKWyR4OVo2Ac1EL6wG0MMH9k0kiVCX+1UfPvuMddDAT/WbvubTV1
M70C4Xf1/QziyoomK4yMcR98d1JxFn2kQ1tc0xgw8sinAyvHw6Mpfvg+ogGXrcsk
9pcN8tyLTzT7P4p2kMY7PsRTpdQnG6NxpNYrp+VkhBMvwB9VoTSWL9sfnZaJgVA1
mkMX17RE/ECBBIsRywtILaMow2puMp43iuvKbCwKmZsY6ZPCcK3mLFuhZvkexaLT
P/DK4CLFsvT8WGMuYA43IAYdI2iIYwj6P2mC1buzs+uJKl0OnDQWkCrVk4QypvSU
kGB+C18YKFNfmZQkG7sRnerhK9JhGuOSNBYEkYdRwb1uK38UwZ+Oq9LE0Miy1BDN
GKkCzMYMq7cVyNo9gQG9+FE6nO95IWvXTESYgxrEpnCeYtJFAzVB1S8t7lKJDz/Z
fwcjGklyHwto/9h0nDYDszkecE8yDAsCUARfcwNsGBlkboa+2W5FXhgMaWdmLkTG
QBRAkCz6v983w1wArIB4T2qMhK2aVj5mWvQFISI9xDB161ZkuIvhUx5JaIpaVmBS
5IFIeZrIx9GOe3n8Nxnf57bvSvXuHv5aRQs3PbNAg3kN8tsoH0mptPGJwB1e1BtS
QDv+btk6i5+V0bor0nM2PCz7FzuciWbB9d12XTe8EVOq2J5f2jhePjC/PSkD+8yt
fcWO3vgHxDVZFR2KjH9+fa8PHFF69Nme4sg97719t4KGQedQYeDSQUQq2I4SzcOn
o3fi+F9RiXgCE510+/9p0WBOpD3LBgHTytllDVTJuVJHlgIUgn/SMvSJIYhEG4LL
pTfVBS77NScC1MhNvzJKpOmFVTCpY65M2AOEGaImIt1knQxCrZbF5LfiJX7za/8i
E0BBRJRc8ceW85mHwmVBjnDDkSWgmhiaGqW/xq2e/X014npjeEQmq9q6IQ0nSfea
xgjBtoxtm7KoP6xLkqbbBgMvxXFsNjdT3xiCVtp/Tl3ShmSNHZMVLDtPvoPcAdaL
yoYlbfgWnW25EmR0WY4GLWDKT1P4azenSy5QQ7Hpd+0mEbOrpb4t8KkpXD+NEtrX
ywOK5oxAmYCKQTsiMmRhZSAs9j2/XszOWIGDLkukaDJny223zQ4mhR7psUoCbgxC
P5XqtDi/95NercagG4rpLeLL6ooYiOMf3RehmWRjII4TjqOSdpC7B4UZ+T7sUs4h
TfMEWlhXTJngAc4J7KK/hNxtdCTw7ni6rFPZj9KUsiVT2bpwlZjhi/Kw5w6io+Vg
OOtoyIKKzFY2ir+vEBP4lEUv1E2vUhrWOVkSWLqqJn4K+Ji+pMM4S/w9BXltngG9
GSuM0z3Es5VyAofTd11HkhZXvfyLR/Il2+DX9qvsZo7kJAA8aN+Je7rq9j1nm7d/
U1IqqlS9sLjUgXxfQ2Z5NNlJHn+uuE1s6CYDIsmbLgIEqiOiNr+8DARJ2nwHfN0/
HpBnHFscM1MhOHH2o/2mRoiDDu2NErMOxkHghtFilfAhcOtlCvGXYK0o9sUDZVpL
tAug3vjBiQhWzf2BgtmddYM0kNkwi7T8KnjNO395oHzlklSvybeZztnsDU+tzp1a
bTrWWD7OAdcXnDA3NQcrhjOib7A3ca31H36rDeAJOa4Ls+xs8Hf+E/AFojuxrXSh
ejccI/MneIqLzQWz4x9uettnlR5sQJoYdalY4NbVy5GI1Me2dRXJbi9KZfKXpbD8
D/6bdSSRz4BtU8dR9vQm3ojj4fxQ/P2RSrIzfTirM6mOg+X/GYFOxRGZOBoZoxCq
/kePndBwhB6orGcpIMH33ETV4PL25aNv7wMf3KvDchylQGQPKJD04wowuNcpAj80
LA4WCNfgupG+YVkvGis2T4gDTtZLaS148RWEzlr93dHO91TqrJS4y5HD0K4jRja6
ldwpYmqSWwA4NG88PjuUnminQsa5O72U+J+Okzohfx5EUclBP9x1Oec7UHX8wM3N
uF8t6jSd1P6HmX3hsi2cgfP3ZE0KQxHSr8DsJIvj0e/JOwt+Q/wQotZNM4a03uTh
oftBLuJWScWUsoOmEiPqZk9LhIJQStMh5UyMroQ67oqOnHI6gOuFlP9jHgGD4l3u
z9535oKx/zla+p2ApxUexDW4eOSGWui7J6N0KL5+hS1dUCl4sIThzs3P5EJv1y02
2UfREtcP2PG1415szxo30OIvt1N7ULjjhv57EleKetuDDmUhywCNs9h0qtDi96IV
0mZ3QeiYzo+9mWHsg3R+UyAWXZnDpyxLPZli9W5Y9fAYhAeLREwd1r+XWlrw4fEw
bVFWXakmYd0/jbamOxcY4SbBh/4Z/F6j9chjPAoPcIH9AQOCRTnpUAAHAK9CGbmv
pSIvFyVR4GcKlz0MnrNNxPAFN9YWrUyWyq8oIST0Qw2UJLbVp3xKppKwMnYucCLg
FelfB5Gh0Q/Ti6jzz/fQJSbTw2gDqZeL3o4qqr5BLtkppiRRLaHoMn1qyvJuSYHR
UkxndZBrb4p1/bIm/bo0ECcr3jnx1K5Y81h8wztx7IrEifanoQWs8b7Xk53qDUvR
ZgrlsByCFLk6wOOVVjwYB/Ez37CvnXU+wIDdFYcVX+H7aehKMdq+DCgq50NLRWIi
we1MlhanZiOH+sbt538QUTc1Djd2Hj5Kra+WrgqZjJIqFObtgcdcP3v9So5jDH0r
ijpHIL5+CaLIMLM01THYL0XJ2JqWFRyo4+CBTTOwzJV4H9C/3q9Hhy3WEDQ78FhP
mjhhX4k7Hkg/st7Ngz4KMlvf5hA0uwwjRrOFUKtm8ksVJYVTAK1HXzcL9mzHXf/7
z9pmTKvVeoHQTqYV1I8ctkmrUe7hLwcfJx4m8VA/dMivdtyltHkvE0yaL3171LR2
94vXU9FGLD2mlLEnBqgaw0lal/nVSfqry2zDiS5Obf73FqCv7mxmB+xJ6yxmwlnb
RZbbkMsRafQgO0hWbci7BnVKpI0Oq4XChb+5VnKWDIl3o9ZoQv7NOD3LKYwdA6IP
TCHQekSF07KqVh23hvCdI2Ky3i3492mUVnBq1UCclra1h/urkaEvTM3c5CC63jRU
TXdu0L2KzEDqOLh+Cs9v/dll3MfoS5wxNhffLzg/ZZ9lZe/Z5ypXNuCC4sB7D0Pn
nOI7JzPDW3qVQdBQGDqG0omF7xIFfmxV5T+gP9rrwsVol9EXuHLiInkMr2E0mpuP
8ZfE1aGhoE6SfRMOTNHqUybbMvw8imjcWasxDv5zxrtL8pTHi2qV9mMAryXQUNSj
ZKaKD00Ieof3JqhZJBEweT5oclcua25LjNm2/LQJBAKs5JNTZoU+Mh8wCYp3uwMf
5MSKcsTZZwmHJydULHh0VHJrATFbQaR50WnvozWs+PtaA4IbVQVzfa6H2q3O/jz3
Z2ruAeIcOxbENMcDWFB/c+XM3XGu2R4Tw8/9wOuKE32Vd4gYunqHHAK6wKax5XBz
qcvCqXfLXLOKhzIDN8EXBKE7O+3DoVYtxAIFoj34ioeBFN+6tkEL5CJRlSgVO1RX
8G5pY6SiFwwSGsaJzTEWXoA/igOb8VfIpf+rK/m557XkAJfzTM8rBcHkty8D38ey
xGFnk5TbHNaAefAQ+7yJ8mUoVruP+nDiaWhIA49b9qw+e0RUalpavCKdaagZ9ZZE
xf4M7ESBhuWFGdkBxvubXrzGbNBtFXHLqeO4BVuMJXvaRbvG4CsV/8+yTJ+Gz3It
z/1Q9vdov9RRAog+SHSlOmUInM0dGB+1btnk1Da+Dh97dSbpbB+/wqo8ugLw/rjW
rVv2e/WFOeu/LZ8bbOf8rTkIxFnxYWazwijNAOsFMdntmIJaQtEaj+FR64rv16wT
BdAuhkMuILveqB4d7Fa5H0O51axIF6zp9D/wMP1YRpeDmyi2IZ53N+kSOiaAgbMn
HivLr1WnUp5tSv6S0sVOv7XIahDWPQQOWwTrT0pL7/pMqieC1HnkxUhC5a2NRJBJ
WwRkRC1YOAaKqI/d8YUk7YJNtn98Vuac1wUrIcm7ArgL+LiRCUeK6dDbXK/khnON
Cr5gMKdZDaLHgyCU45aO90GlpdXUBSrahap4khRvuuCwxFropDfmRz23RJLWgdQu
SkssORv85qEO1UsKNVJaqC+pgs6Rbo6rhKYHUTUEJ0/H434nAZBDl3VeniYbHWZ+
IyLYIaSVtW0o0TTPFEsmwhBsIcoeCh2xNi5rNAfd2rlJjBMJpPKZxfkVbuISJQCs
VwWZoOehnJr78GKX2x+jLJKl3NJWc7EKIFu3pCAormRWqwemiUZGstHnIQ2CNe8Z
niaYnr4u2duAWxmYArRzUoVHoCOaer/WTy+3JtT3s0xdkQzcgBnu+lEJGK9YF47F
9Nl0zyMmaaOMHdUNrqrL0jwhZIYn/xijygai7ThY2OJPhg4mowgBKM+k3sDMIHBY
XO5amC/PMxV2IK5aRJYWe8ijhMBHdFHZ32X/p73wr/aBDEqZ+aPhh1LY0oiqH9Sk
oG79cWFQZ/zYD/i2H72nAtKLlqTjDUznxEtRRYNesmnK76gcqwiR9AkVMaNC8fIT
kG9izqCtE3rlvjEY9WMR76l0TPpeAfqMrnpEC5fXDuUlKo79pQIDj4RuvuU2I7uP
xZTFtCfyvxLM/H+E44wLhXcAeGtJU8ZiApfLNPoQItsJa+OQM98wEmEIeX7UjYT9
1Iwy5QqXL25f7+J+g4b3Ih0HezFI75TYT1SDTWxdJ/8uk02H0qS5wTcp7P9YG4Xp
/Afr6BdM63AKSee5Z54+WKLgW1k/YWJE66Cd0H4LxWGRDTCkOLMKrztO0p/rc36L
YeWLmdV2n2A/o2FgJs02GkFfPoopXysxLJn9XMaCQ8Y+6xrBhsqWYVY0i4fLypaU
b0sQo1XPR4xfGHZ8T7ccLjpR6la80G6Kk51yRFQlsZMrXnPuvgwRv10NQPhwUAvR
ON/+h5utvAe8eQ0Hh7ECO5R4QqCIv1yLLGkDNChpKFHjgA5TWlHgWpzFsZSjzS2a
5h+WvVL/AWvQIVFjoZQHysVKnq+M6rM/GrsDmtbQ6xqAtzx0EcLMgilInC1DS6d+
0gB5dHyBCqPIT4YHxHtmqyP7Etu6+uHJ3C2J1TcAxy/aXlw89rYyOpIU4Be6+WIA
BKsneqjbNgza3BWk+B7Qaf9yMkia+nqOmHiEW6Erv2LEqwNmn7ivZDjOVxLZpeVl
Ezl1KWPUHO1oFLuY0mcn7adQWxObLYn7XvgtNvdei+MkA8VO15+JNgk7o0s27g4H
gqeQruFB/qKFk0MW2AgxELDeSfifavy4UEU/Fn9p4jsYdtS4n/D7Wb4NvVs8R6lA
BiUOCBR68MdVwT8Rze4l7PUxHw7dW/Mked5yCVzZi3vccznSPfL8HTAMdz6sn0ea
5D3ooJH3rUilXjuw6Urv///RLYlSZq83CT+5DScL2fOSF40V1pUg7odrKPeEUGNc
Jizw8/r5zwYDWueCa8Z1CUvoDDYPPhLNpa8bAhybX/Tw1P8d4B3SkOlvYOYL9BYi
ELU0rSWWp67HQCz/ZB1FsLi6AIOQaUfbntUiN849v9rBCkgnXnQpVo9ipVPecG0A
fRywwu5tm8TKuWiGMh6dTPnb+1A7t+GhbdaXTzuQgWtdazopr4cgAyHPmFCJbwkZ
rJgPk/INXeCMMxrBGSKgbh4zRDvTdeddRrcSN7w4J6hgfRHTUKqG8S6EPynu/F7p
is0KK1x6egaPWOTFGPpTgZt2GC4+/FHSAoZneNBne0V9Twa4p+EOR2C2KX2wH3Qn
JU+XnmwWDyqWPDnfjFrMKLOPpk4wYZWcI72tTaQNLiL/bYWVO1HDnnWe0Ft5AdG2
DYgsIkUxy1AlEhpSVNrrLFE8adABqvbDQ1aKX2kI6toXuEjx8OHs8Y4kI8Ki1Fy8
+9tMD7RpNrUqkUjdQbZU9vQjEwlYQs4WiBqJkLznqQILJQaFCPhHR6GqkfNB9i3o
M5iQvYnRGpaOzLC+d6j92e0pXtdpOhNi1OjemdZJ2B9lxIZZ7j301CF7ZRXnngj5
R4LKswnljFErx0H/Zgl6eHJkPDb9npX1kq78I4I+gfRYZ7QEqxpE+OgeO5UcR066
XpKwXDq2vDzb/UqDbKmL5wPU4Wuw4W8R5LCeIQudjRpUut93fZOa1L0eVbOdUltd
PR+38buAHIvFP/Depy4enUuZwM1md329OZK7OM/r4DJ1pvPW12pWRgUdyiSH7/S2
1NlC5i6Ni0Es/bYEkbSMCAwM3vV6HYnoSPxyW2RnazzaA9mVIDKoJwL3O/FPtmeA
XTCWCTTztG2zCzctUogEVcjoJziSl6+Yh0kAouZm80jmfCkpr5q+X2xzTJT0yFU9
TGPXzwe5R6YsGOYYrOrHM/DzCHL8KkDvwDgZb/PUsAlwyK9awAUj02+0aB6nMn4i
9NzgtCc9+m2TOFWlL7v9xSMiTatR1NwhhNO3UNAoPg2C2HLUh8KGTId/X8oABuyI
0lKFWapFmPHWwb7EvL6nzSokTaH4Tz0Yvi8BrIbevMvr/6GVcg9pboLsOz3wI9n+
ud9grwCv3BX/oofBubiAEeU87bribF/7dry5+yjlLMuZpT7aHSJXa8VKWfIKANmu
9GzpQcaUt1R37n+PXABINgjKBD/88Jwl7kbo4ce2rhFDWjhdyY9+q6Y8e9lKZb1D
rQqSIgylU2MviG3gXowSo6D/8G7jq+S3+ylbN92jo2IGG6VdyRaq+i0+U6KBdwb0
C+i8o890ydeK0TMf/w7lHjatrl0mGj/Z6V+rgwYmUvTArMK7KKf1tj5F/RRJVA+e
g028o1emBbUhBuOhNnCsLDMFCuQMyuUVko5+cky2Rt1N4UJWJL55/vNBjBQJ/bJZ
2nkjWkby58RY0S7olJfbqm06SB+ojFpSU+tfIkTZcHCrXBd+r/fuEySQC+h8SBmJ
G9qKP/0RPHiW7T5IhE425zGbn5ffJLZeLazIJNeYCVsR7B/y+FYPSdM4L73VTPKO
zNFPdtJjGWi7trNjuMEJcFSjilk5scYlfr+48eHioMp6KXZw/NsA1RAU6VX0+j7r
PkZD24HKCvOfDWj7EBbMXxZXuDx8Ye97/fs4wlwukf7H13eDAB+zkIHz+VqfW46Z
N5kdUW9MLEQREtikcHI319SLBpbSzpgKcMHeDpz5DklV6PYErBFXrU5f/SSrTv3O
4I2CRb01wTHHuA92mQkZtfPxUbdlK9OTCNNzWboYaYXqcvfVk/GLuWLQpeiveJ4A
iyRccY9VPleSwED6VYyt4Qrn7FKprS4Jw3491KYoFDs7VjB4p7zLuybeb11IhHdS
VbtoGIaSu0vssR8lfrbEJhXxnmtib6UaNLgkw0+v18nfYToJgQA0nvAqL+zJ+1PA
Wss+wuYj6b54vwbqPkZN3fBNuXcpglkNPNOzGmITPNisuaCS5TtaQz8OiDhNRz96
ad42M/4HwV4oyVc81y6yph0d/zKMT1LhLCZD9E28Fc9SrkGxtHaq3ZJyZeAtkG9s
O/p8UevNaxWPRR5RHB4eHCQIa0z5/HNFFEAQYxGQdx2EG/+0Lx+3B4/agn5XpYZP
a5LhUfpzaa/yO2BQId6J1LuORfqMtXh5FAoLc49Vw2OJ3VaRkJw+wM8vXlHp5G+8
y709WZSiYGdf+XRRybAR6epaZttP/nbp+Tx4AN6DnOxqu+OBNkFr00hAszdLJjza
DFRJgCo0fKWefb4wIwhqk4haSXrxJKwZ6grpx1IDy0rPPrz906rzcNc9DKOrkSDX
iWdzM82CddTOiaKIKoeQqDXxEjllJoALfYML/bFu/FfvckdKTu7RGmAihK9k85Yf
KbFT6QCJekpW89B8wJuRPFqghEv0BrI21hJnXuCBRsxKP5zoQBbmotILs8HRiGjV
098jwVkuvjOZORcMLy+6+NCgfF93wvOJ9G6+Y6uuU3LEkZh+iVgHpnlmPHkXI/6b
ZV6WuzyE9S/QoZdNBmub/66Du4sE1nQPxlYSf7aEdG4BLweeJmB3KCaup0RUqhfw
KOVvD6ZBFq9leHifQEar6mW5NUBPM9rQ/2pbaKVXtu7qWp+6ulHIqba2/uvs5CX9
J1j32dx+BmvPNUnvfbEg37tODSRb1Gx57eDkOffX7VHrZ8wpG61Ae5ag/N0nkOjD
HR0nC660hJs5lncqDskttL39bpXwKGeQ6b2zLVs/zvVlTTP/ThiDCB1Kj5w+Y+fE
vGMzFjZOayb32G2Rh9lS+htX2lRjNiuT48yPOXOo13wmPJxRLqiVKteQJ+WunoMr
EgQ8Dxl27yvtAfIyisQsaokmN9pdLdqQqC6yD464fBPODnlRTwoAMTYQY7DNwthG
YMBkweQqwhz5YtvdpSpRPIbFQ7qyim0S2G7kNHoA4zajo7rnCu1fWmADQz/L8uxj
L4mi+/s7LwdvN4ot7nx7z4UIKOtIfwenjPHlRgJKSey5K2Sii93ga+Tx7bWPVyGT
`protect END_PROTECTED
