`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoYdOl1mAXlGoyQuXGjcG3HgLYubjWPhEzYyvQjBKFW+YYzIU1IcE3WU6k52L6t8
6lUdw8kaKiuFcBeOnpgH0k6/9ZR6MBxyMiPtWQLNPxm0wta6LCCNKG046bu2UvXd
0iLzlifOPtVeRKcRWAmkhowwO5eWEIUWxKXflvG8UVtS1mixds68BZ6GSX+q5Y0W
9yfx0go7wMBH4XxsvZMX3tWFGonoYZzf6XrVJeer5HitztkQb9QpJPG7+g4Zao4Q
Rf4WZ+agZD6WVFeDznVRoTtEqlAjrUNXzzL+ZcHxKqR/W/f1QFTmckck1eijLDDa
OFzuQI1upW5T7hHA8HJ3Zy3BkDrHydT9z/QyI+uth4DEnvJFMWVcfld1U95vw3Ng
/nxhZGZcjoxOMmE25LgufI+a0ykXG/2bClYABh9nfmL1G+fgFH6nI9mkUF6bgW8D
MQsqyvrUh1L1JeZzNcurGTuj8l4GcMpjLqH6lIjmYRCkPKLixuk0oe/fc82zdEii
k/K4yVRp6hLE2YFQjelizEKJNrJlKlSeqbzawk79nLVl9I/p0RLlvlyUUk6ZWcKh
jgfCL+bQ8F025+gBsZUh2/BkXTYGMFIb7INs7UFtreeLAPhp2hOIr6kT+eATopdJ
puVA4LlXJ2UM/FrzMEAbrqCAU0RDOQrLxfjyPEsaNFjqlnAkf7DFjuIR5MVnkt27
QpaKkE3E2znh2OvSVHTYoJ+qEi0KUobc18eGbfbGBPs8yCFJlrL3fjekMLDzo2ky
FkDoSzCCPIPAHtHPM4FhcZEwP7LJmxIEhbJ/BvqQiH8/B9pEFb2FbkZgDFcni3dJ
n6blWNPjyM3w5lGPQbCK7B8hE4GXltoZKUKM4fS2niKEYLuvtXZnvW//y9JCIakY
WK1yjdpSOH+SiEWWvRIdBYkPLzWSGbdc5UplXA79KWU=
`protect END_PROTECTED
