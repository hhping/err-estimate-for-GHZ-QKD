`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1o0mIiDnSUvcOqMcFhud4fTV4lVmQVDWp869v5XbSe0M1uZw6MrGaaKI9RcSS0Y
IhqsYpfKcfFq7R1X+L6wsWmZNwcdpo11KDcCfzbsPr9Kf4wBlU5VlPXaKPcbASjJ
+Z8FF2Lve3hcrpe0UVlsyKLuEPf9KRcOGvn/zL57jAEnwGkQF5GVqyjrm+p8BLlx
3rCyo9KjjiFquDgfhA3I+BSrgeG4Tc9Pw86q/CMGyux0OQYCT3WLRTF0wHjbv9db
Brsx1Vx8d2r4oV9UXvGJGiMqh/n1JuBTcRtFKLIHAi9XxCt9Dexyz9DET/i4sAtX
CD/X+aCdav0klheKqFYrD71oMu95E71BLKRXgAihh7Pb7ujFLNmtzqhMI30wnPQg
D4R0hzG3cR8jhQ1g8xA8kj48SxTX52RP3U/F4QCRxBnlEkT5KCUt6Q+Be91iZaNE
RbkLpemGeHkjPQTGeOMhA6MdLsSNCEke++k0dxfS+IPReYLcJIaO4E3KxBY7Febh
lP1MJKd6m8NPlTL1FQUxm+WO++tNUgcE2q0PgRGnQbU9ADJYPq3pe6Ko78kUY3mB
l/r2Fr6fa0Ek20IzZhmFQAjpUs7KXLU5iutervIpTvzh+uBxtRp04aub85eL252D
+ZE8Cbp0/3LUjD4ZECRup1bRWrU42LMVIvxJaWN0h6FhwNW2SgYHtyBV+RO4QlWv
Wey5lTfv84tBfzSU0Hz19gKp60mkPNBkUK3BbfeyaD4VZ0DFpNFKbpaf8u2oiGXs
MJdhucIEvan9kaVuVaJEXBe2ITD7i4QHNeX3bkXi8VkUTpNErrMHZ17ERayQfd4E
Lu/Y42t7Kr4R4C1V3VkUVNu0xBbOYbCYVKWa5FPu5wB5f5lnf1ShuTVOpr4pnKKC
3HBHtrstFIgk6pIghF8kUsQr4Ep8tk9+PQa2zVomEhhRP+OmNJWJ2ltWKsU3k1it
DTq9UIZqj9k80mz8cqPHw9STjh47QbfFbDcCxmNOawA49JLUwec6iOX/JOCSQMqo
NJWlQAM2Lvy20dxJu3yIaDuVk3+77r/MIhEspcRh4jeXTG9g7C3+9OsdNAAQWLOG
AZb6OX8rB15oySEv3PV1PX/TgQAwsrq+X19kbyVrXw0fwy5rtto6SKiIyTKEZaRj
Sbb9x+2nT3Lbs27GOjfIDL30VaHe8GYR9TikPnzLN7iyKG0GHyQ3AScLX9jRwM7J
BNAFgcFwDiO9tDQaqic4m7Nms4/jqrfuc/no+HjL1L0C1TDSvTaqAq74/7Yhiw5H
bS8jkPuqMwbCCTWa5c5b40K9FKv+5AkUEN7T0VSntqXWw4bbaxAb5BD912TiCvIO
ziem5BAWntobee56dcUMxzPP0FD980Waby8qdJthfQGDQK2y7Fvh5e5PC7wzM7Q2
bL8WH18AxMt+zX/KX3kz/xwXRXE3oz1+Vy4QTT9mnXgnAR7EmjwDcoljcBe4Htdn
kfuZpNP84o3unTCrxgTzD9ra9VfQb3JHALhLNx846hoEO96f3gK098bKm05rJPcj
tRiagM/1Dl2+B7KSebd2YmkEiUjsydOaH5lAuduaRhfTBjb7LafQkk648WjmIsS3
Phq91d245DB9Cw5fG/FcxnGWwbPaHFgwY7WatVeBZNIwLyLViICnhwrSqMacQGPp
suPn36avmV7zpaOn9mOebyeOPY/FCjS0wUpv7S3LvkTxUsTOp5tqInYV+oeKLvZf
AmOg3+S10HJAyQUR2TWzgPCZrq5Q80WjZkPxUC1aJ+TdCNOSszUxxH6KHHFUd+EZ
XsxE9XsokoO6WA2b3GK1wbtES3VYoO+CQ+bzZbP+ef9YnbXKfv9OweQDcYgDETnQ
M4eeJFXPVvHaNSjhp4tiRIbMbcQ5B08aM0rzPaYARgJVBvzuj6cSniK7p/hSujUZ
I6uWNthqrenIFOHswN0k8jIVSbJOk8gLmWEfnoFdpshWZe21zVXIQ/fstSAKiebM
493AqtsfZpmVW0MV6TxWOOT23hF4mnFRmYT5nIhyGLeeyNZdbwtu8EjNURRoxduk
ucW6BrWOWz0levntpfpPCK/mS8m7e9h9WjK/YOynQtmctaUAg+k0TaEBvsW6xgPt
rvWt16q22AqnLOPLmBTrDWoGaRwc93HH6MAy/+hhDocgFVxnhjGwpMFrczV32F5i
3OGQIG5+TalGuBqWd6WjrumNdBBfGzIQKfYY2y1alEsV2CGeTJRWGqufLPdCRL3J
Uwi0+AmzuFszYsrXNTmz7wq49jEqQoGxtkldW4O5a8yak2ceeAMqmkCffEmsQtWz
MG9lczRwvnpqFQaSoFPKWwMorF/L0C7ydwAihQbNynkxT5GLZln9HDvwAt410B2P
0AachcIfEaR1gkQCbXDgseLE74yK4YoHDBh2B19Nf/dPKdCQRQwCj5meij016NA7
DE699/slu1/LKOVVX7j4to3ThLIkGW/iGvDtxUGhGdioUbIuIr/hFDr09Db34XbG
U/Qgih9gEz23l3JwLLxGhGTQyIyUBi6Et/DENNWe/NsEkhQR5mOMn25oFlqdIWaT
LxUsdtkwHjomosOJWWMFpgBprOb+xnCBgGcaKSyIp+VbsUmNQRzWqP4n77GeZkow
SZz5VbY/cJLJcTeYNXCI6uCzV92QpQwGh7yyWeci6ffwy6v+RxRyWEkXv+wGG7rV
YYS5jLoKf1v9pJxXQwf0RVXwBSVXJLTonbxQ/VQ86AF2Vc+aJyOUlHicfObaAjYp
ep90odahGYhxb0YwK47T4eQLcf943nJmg66/Fd+In2QzJZO9HnxWZneyo9IlG2NW
7yUjLGKFpW5I4WVnocl9aoF+QMc4GFL+DXbAJDtuxFoF6yeXntQQvaJu+DClA/0R
3Eg8a6vlTaBkFTCAjSlpXe/x/elAmd13bJye7gEu9JeHoW3wfICq4SivVYAKq2rJ
u3xo0pKIukGYiqXULIek0Tas3CRwXXIAKHQBbs/0sLcyjX4jnc1LKv+vpMni4Zi1
PU6QlY6Pd9/QSMby+YYnQlTH/D10PAmWqHLnQ+1h6FsI2upJWMD5TryyAuKgiwIK
wiXQXREjeFZ0kDWeqDcEId8PZo1k+StU4761P3S0bY8me49eVKt3+t1quBPSKLwr
AagUTBbNczTTkI7wSOGoiulrmCPf9wcw+aaKMbFOpQaQztp5nNi8tqE4EJ965Czj
6y82VJS/uCR41jueHpVwT57n7VUjHFu1qMx2FN+OeNhc3x+RrVhctKZnoP9bPNug
GDE4mcRvH6ti3edHmxvPM0E3G/E4sqfaffMVBzKfsBXl12q4jPTaEhHGzeSQBp1a
3XbuF+mYrdWpympkJ4APkju001RolNd09RrsiC8ixjWYDEGAecOnvpdsjhN65lTx
iQ+5A71X5nFdx7pBXz50i50hNAJbYta+UkRlO2mKtnKTSO9BHhDA42UJL8sHe/Wr
vqw2lgBrvtkvYR2IciRG1uaY2EXMS1VQqVxKI8/jjidi+Bro/TnasaKvUYYRicQt
H6uqG4EH+ViASvKRW4qlDUAPKxW2UbrcsYUMfBu5hQO6dzjCXZ1dxq64rrE5yknI
`protect END_PROTECTED
