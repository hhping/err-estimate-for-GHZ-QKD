`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lhn2EEzvWN2Lv3odcNPxMcYe39hvR7xR8mGeVYjWbzDKhovigu5W5j5utvSF1VLs
XEird+zuxOhmsioyuHTuNPyVk0pERdBIQLIiVyXl4er9YHu30BqMnlcw+H55m68J
6tfLT1CLE21AE5ai2XpwaBp2+IHt3Skp02llL/wlmGiJFLuz3EB8bI2zhH7Q6QWq
3/PT26m3sF0MWhdBuDYmItcqNvy2Ub48xbFAOf0PL4lMm6fqEzAtDV9u8ROTFhuB
lXykjQnXEftY0wVnSfY4Ftlisd8y3oWUggNIRorX48EvQzfBbHd3P4WckNo2++ER
7JcmAsMCXg+EwVHAXk4aOe5VxnmKucNHaw91ZdBl4BOrg62TQLcnSnsEtepmLWQP
5Hxaw3QjNPgysl2Cw2oAPd7OLDwA9p7zjMt0qhSg6g6oHpqgCB4MSAGY1kkJ4Hyo
0cQm/0BQgSeflCPasjIU1yshfu8uUK6SyXuF2rBRUy1Rqc4WY1SKyd/f6SkafmgB
774ov3jJzPdlNruhHI6OeaH425DzbsXFBH4QHTnlYtBlqWBrF5Odh1BrYP3/iPnT
epeYYEdSw0ficur19G4d/lD4z5mhTkqHaJjjPoQxxx6uZUesxmR89nRDrKakmIoI
4YII2CRZYNwULvxudqSJiZXv+jEfA6p2Ksk2SKWNxyR8A1SoQOt1V/MHwnG2rn+C
GNq6DoXq6XlWXivskKRp62Q3mkxvPkOGFKeLraoQAno7pZfI2c0p0AG/3C107WpR
XvGo44MyN5+QXccLnO6tuzUTEv1+jKXGUOdOb/bMwpEe52qgWIVQ4LnyeWmQF/oh
prJLA/2p6M/Obk+S4iHMTWhYsIXUmjjyfiClkQ7llVvSwvgAil7SjMXGHsDi5GY4
yMEfLCz4Rix/m9IUNAbK4PllCwgFvmSHZI1HhZf/1/yjAOX9T4N4DUphpO7Pfvbr
gFiyuxM3f1UmnZ0+N88zuotsexbgTHU1/YehgX1lt9FcDd8VBBVpXJbHv5Y1uUmN
xpORpXcTmujRXQXZ2vPoSFeqVSm+TQp0yR+av5c0ToaYXDDp3OhPhjOWcsi5UTTx
O96OJTO+QuwT4m82g/pR7xrlUZQq2i7f2wsJ2jzvDfVA3f/B+qEHCkCuFsXBJlPw
AEpuNhLSNlY13wmwOgNq9cJXjUCkqBf7qFxCRJUByarUsUsuNWYGt0IkYM9f4Gd/
W5vUH9BLqwGqoEvRDS0gcR0+a9J37L9gQ1+XFVsGQCg=
`protect END_PROTECTED
