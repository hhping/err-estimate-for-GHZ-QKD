`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ydk1CbBJ/viYnhucU5TEq7hWvaRcrWLHOH1BSxvcUPZxSyhf0a024uwAvg3yblYt
I/Kx7+rZ8yjG+DbU4Ju0WlU5OMCBUS1uY3hppzTaJHnEA+HwOO2nu6XdlbXXZ4cj
pE9Gk97nyWgOZj68Fmttvq24xL9cUHDBvn3Mq48FcAyryGkYmu0gmlXdnlr2ed0u
+94Y4E4NZJIqIX5ahCbitqLkb6B0D58JDJHu7MkWj0mnJTmMGwkE2RHzgtGqXGN1
jP62yLF0PB+4LmbRjP/5qfyLtrXtt8T0bgM8bDLpAtRPaZpfdECbVm3O2Auj4U7e
NFs5Kjo96X3xXY/zVNodynmkGzknBDpFAuHjvR6FYBmoeKPiQB+fu3BYGWdJ3S4+
YlTDhP6c8Mwc2/qVaArZuUG4S9SbDV5tMsflj86pxUaS37BtRDGnUWZNFv9AQjmh
XuUxzV8y2YwZLs6/RdAXveN1SAqcQw2Pyor71r8gkypaHI2oQCKLlXpY40oUCfVu
RCa6XhuLmvAMH+5xN6/IYgjDT15wEY+YydLDicjDU1agHooqDW2Qcg3YCajuWZZd
JjQMw51cclXKd353LsOdAsfQd9OmhL3yuThii7eqDJAfyU13KmAGPb5O2rng9AM4
rlQ8t6FtRTEjh5kAUo3l79EM0zCztQVG9nxGosi7IAer4+guSxNhCLswev6yql1X
EqdxOSXXDyy4evQXJAQ/MG8Qn5gVtY5jYnAnFqnIMPEl0i0ik3+epb1QRgqE8TZW
Rx1s0IMw2cCdNKyV0Sq5FfF9QtEC7l/MnTQDlxWQJ2fvTZl0z8uFavhzS04Vcg5g
E7HwQqoYXOuKZ68TedYIIP7ddjpt6c8p/m7q0lqUkLB+aJc4pBgML4MD7sQiqmrI
A+uj4FFqyO/QCSHw+hqry1Ba2DSQbWoDzxZCZkrIz+aOBss1ZWOCj4wwHvIMQmiT
Y3crB+3Q3b+rCuBrh+VXwaTN0PvGt5BhlliXrzbX1isBbiWk0g2WySGPrwAaGw83
PbD1A0lBMpkCEkhLVhxpmkZSF2rDiSn35XRrrYUFXmcK6m+aPewj1XbAJZm+X7Aj
fO6qFTDVcKNiGkQGgF1XK6cBIKF/WlaWSzA0OGuU70HZ/TgMjrcrccX/f/P+PyHy
Stu13iiJlsylgp4ka7w0fZiXYdVrK0QXhCGx4MiBTzlnN+wdphSW1raLLK6+ZPAQ
qumfFoEXscLfS2og6EeJFIuObs3MhkMJSCAXKDQMl2QoS5/Ocy2rx78c7ZyVcyV9
DIVSXyiZtcqeHORi84XrQoreAZrMQhqkW/pXVkBFpPotxHX/Rt475dYUQul0+23u
g4BkE6OdB/0kYTqrmCarUNErX4sBFWbGUc+MoAug1Sgl5jxaUaDHxjHqAGZP8gXv
eOY71C6E4rOZrLwdJDnVKp7a01kL3sQU2h+Y7GhgzpnyisIsJUZCJ0uf30EDYQzF
OCcHn1Km4yZ3xpIe4A2MEZ1aZVgptWKXmr6zVQBxO99zUqA8nTGICOl99w5FLYTg
3CoK3cUAKn9kGzRxSZNQv//KhuBqaN0F0gLpBdFs8Tal53+0M0hvLpahRGUgBlXl
`protect END_PROTECTED
