`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+k7B4JNfwIC0+A31Q6K685FtN+pvEi8VczMSY9abkAt+G1FgooJ1U38YuysuQjg
329XxJExzus6QOYTF/H1EzXIbpNUQmj7Z4iPeuOoVIC4NsOSX20AB56iClCbiwzP
f9WU61NyT2TCsXC+SgH3kmduDTurqQMiTzJ9JD1fGwb+T1LdYYIhgTYJ2aQ1fMya
bgypTNV05ljtH4mVoODKhzYOCVRcQdE8m6t6u8O4X7qtih1Z05q6AXX+m6JA5Mgk
7S5wbfb/vgGbVEFcd/kwQJGEsz1zFGzat9BB5hxV2zDXE3uJLYIPoN5Cr7GYM/Rt
F+BtjRPoqzZGo/2Ydsiswa4BM0D1y9oJFT43jkXiIpW/cxJxnGyrcBKDTvcVdCUh
j/JV4m1WDwXnqejxMPUnIf9JnQaoPiJAokFlfM+87qTk/YJ+HGOB3OQFN6pGRgox
le9NhgxhGN8VGX/90d+DU8AHANGRmBtoN5C7baXBM5GLXeRoSO5XBDtr9tebZyKu
6NnvgypgjtCmRQrruJfVvUFfTbj7hQ4doiE7bTMCceEp9FOG62kcyPCdb5BzdPBf
igeAp9soIDEo/a03z7rzKD0bEDAS2idjkxwz4K3RlKFpENiXqhVeTmLM0CXCdwFf
xIG5YxCVGGs4FM4yzdVTzQ==
`protect END_PROTECTED
