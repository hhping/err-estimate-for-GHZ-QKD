`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QDNojhjM/uIEWOLd7rOhjOb+1t00N5nKvbeR2RImMgSAGsx9w2pLvlfohqrW1TAE
fF64edBxYMuHYgspl8iJ5aEhHQQbq04CwSCDjwxhvE+6Fz2urawB2VZ1KDlWxpfr
joFc1OxBtBlw1nilzeuwH+JpuuVhCe2OE7y2MO3rGx6keacV924SwzkzPCYTVtSh
dyuaR4z3mo+bQII1oUw4/bUqJAFkPGgzdJxygZgrDVcQ27uZDvKRI3KnbBtj0Vu6
5tsM1YJvGJ/lICTn+/uE8xVHZ2pmJUu94ZyzYznMeWMzCpL8OXpEgOqkb4DT2sUG
YoALuyrO7BAX9aD3i8R/e6w3sBDpsgUfV3taV6q1sYlKEI4q53tIAsWXOzrXj421
6MC0YXNR/nCslentNuGJsE9U8M56HBLAA2KNIBzy/egfOlv9DH/w2cERPTQPvZMa
/5vs9WpqbMW1o8xs85FSVq+XCt7u1EHAbfkgc2jqpRneKEKzzbVQFUJ1el6Uh5V8
eY7AjJy43uZUC2cP/CS7glbTOCxI0fawlMd7na7WUVwx9zpGXNDNNsSZXBZ7KxJ6
EXLWkcHudDsoaBoHsZo9hL+1J6h0h1u2ZmNO1pGtSPnKVFB9IE7xSKiehH743RHo
`protect END_PROTECTED
