`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGZS9BwMj9Nxug0pWk2LXajEzzGKbNbAV3QHFWqPjB1BYPrL4hcGIsigdyDa6R2h
PXDWRvJIS7UdDHr/juzm4aIsTQXFTfozPY1jeec/swgxkDK77YivOxteZ+joJ4Hp
+VRpfhu+cwZNJzcv1eBQoTtgaYZ79EtGNLt0jhTbR6ccAAdGIECibTr0nmNQXnu8
nX8I5p1hHe2wpgDEujHvbvs3uTCZ9FpvHMaXt9oqjN0eP8lpNCVEd4j4pPus0G0L
vojQibqZQGxmRPqTp4THnIj8Bt2YGvOyg9ZDlmKd2XDrxMpYjlvK69krnwGReIwB
m3QXdLWep4nIrJtI+YukyMEb9EDubEw3c5lYnxUuuRvFu+RoGv4Oxyf31tL5Z3o8
3VS6jwfNqT0RmULml5TJhXju2YWXmlwFmHskQKLNWgKhI/RoE81DM/DZxN41Qord
7Tv1uzPPjUmSsSy2Z7oAAmXUttkUqb9raqZX3aeCoJl7jKS+9NzHQtcxe7vZtGIs
ybDSPsHkie3i1v/uqhVq3rR853uoMDRj4+f4mhU1gGiRPHSOdWAxh5f+yrc9j/ep
WmccohG3A2WzwESXhABJWjaVHJfi7eN52M77bh9xNSHHdaz1ul3WmP9NUpLf9j4d
+WFPzJtVYlhAjRmPI4HKBw==
`protect END_PROTECTED
