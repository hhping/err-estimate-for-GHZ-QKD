`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWt4TVfiUhR2AUq5/qU1wrRF4IWuziq+KNR3+QhCj2mPdLZsEFuWddHNImnlWHsI
wkHIXEZzZj11waHq14S10OHhOYhj6y8bqKFqN1XSzIZj65yCSxEvfTMFL0zsbFP0
FqgTlSoq0QlDPAOqXBlGH7x8/o+15yjWjJ70E1rd0FxAIxPA7zB+jW9I+JYFSTex
ZU4SJVbZ//HfsI/uh0rgak5uUjtlURcafK1d5osaesb8NUxEx1I+0VTZl+daP1M2
gT2L9ibKk0HTPsbo6XXY0fI2uamNnE5SBhyF5mtyVvlcyAgvOqx4QuzT+B3nWVnM
EEfaqx5NMgbWLlIU0PJVBuBmSj//fhj58OoYqPwILMXqb9QpUqo3iJTiSMPhG/Ba
pAHxIsjN+VesJlpu9Ix75Jz4xhGjmIR86Bt3fK9FEAxwwnSTLhpWerlV/J/FGbVS
LJnaMz+GADMGwwumECvYHILg73U9KcrRNbkl7MtbsbqUIA4WOb7xyRrH4ue3MiLH
+l0mXk1ZROcGKVEez76a/zs1vwEb8lCQJh8LgRDyEYZNeFofUJyyR4k5372SDdAU
ofcc5XZaYVN3BLzyvd9Id4qHf4oy8a0L/PSDmMdRzAa4fET/IGPF/j+8XcbA3hfi
NcY1G9DA6jkUY6kBkBHbxD3WjJXez5mHkPtyAbkfkuLc1UbjFVQ9z1pUKz1MGl8M
Q0jwMwH78w6YzmtNLO7NwdGaNU9bc8dBiPJcY7iq9ZTnTH214GnGBfTeTT+lhgSZ
PyUyXEPU5WtX4ze0KYGaI+/8cEiUL4fO4ro+gypUwJcAcuGlxAGnoDupCYC/GPd8
18ggLL+5dkARpPX94Wn4D1C9QD8XVIdIzpSaG/epY75n2PI0rCIZk3D5AyI6UeIB
6PaPOq/LQHjXZZTZ2hc0IvVZWDwGnrm6PD80x17RLz/9ZE7Y/80gjcqB15FGImfH
E2xX5lMVyltvXL3GWpZLIDChU0XelHx6TwQqc/e8p4RkQqxfv34p9Lt2jDeSNOV5
xh7oJ6SHj9Wz4pQNM8eF4Vm+LZfLxyKLAlLlHv5QyAIQb4WWNo5Fu7PD5hn1pA7q
jKVihRAHkZDJzdod5yyTDCqdFCxUy00wOJSIFF87Fvbpo79k7ja5CQqMpCbAWGFK
Mlh5jKcyWnoV4oF0opyqMzH1Uq0iAUJDaE3MPzgYpGo3YokMxsuMWXr+CU3VCBio
Is10M9oe16cZWiKsDCabOj3HMSCfJhqnzlKLmeMqakPevUKZiM/KQ9Y72GxeXSDe
+i98dGuHtrB2WHYEmDTGolAoPHM+jHO2kPw0/c8NrTqgcVg+lr6GCtKLEq0rSDuZ
7LUlgGOtHmbaUOgcDlMSqfn9QjkNjhgCgLKM+Rd0OCoL+ibVofsENe7TEe9zyIs/
VHGL6OYzEWbAA1wukJYexTZoqTvcul+dSN6HoCLhC4hSvEPIThKLB0yg2Q7Tybfg
zfhzuwvRyuPccxQPlTTNth3uBJ56hmEn/Tlik+exSSEewr7st/pXpuoXB/DK7gGr
zn+tXEIRcuVeFG92I5W3bVK58ICzflqP0tqJWsgqoNiURLDr8D+kM1yGjt1Pk/SM
EInKD7CbmWYJ+346xNEu3UVfDCcHuE7hfniUd/s8joRJBufUzskr0phiUPIRAPCH
o1P6CS4XxfBduhku49OgC1j7Q/4lve6CD/mDJFgw3Ee3LcwPE6TNHmaVrh2c9Eci
CPMDqD2+uj7WoXa3CEW5JHw8JebSp0xfb5Ya3rF2ZwAXLolcHRey33arK1ek4h1s
vyVld3btACB7BSlSIliPBSeEWUCuIAyPwdwD4BQyZu56x0ja8YNSjDCi4T+J94B6
5yiJHv9TsyzN5F/U5xWPNLw7SGW1aqYphob/VU1oLN5+f/qdBMxVkJ0z5olWHfnn
Psd/KjsG5fIaLcMU/VWrR6cfMC+WxFKdbrV38jf77Z/DelcyyBcO6RuSKgeGKWLA
a4fR3I2UaHTTZIIUjnA2g0V3pl1GYIdxfBdzNHOGA81AyndDBZ6Trq1xV91A6FGW
5ia7b3787jmhadvoo/VroeK60bqTWEPhoUDu74pVQ1Dh2xJMm9ZlcvGLiCa0kpGC
un2uwKVNwnCVKBVhra1Noi7rUxMIKTNX61+Vt1fH4kl4m4mul2I/ku/tzIQnbkoF
nxwLPSR07GF66GvaoSJoLln8k6v/GVXCYhm3PVc6BI+vjynoQxThPcOJUIKDhQ6n
PYaj7N9/Ru61Ht/sHUuW1aezr9GRoKR4JBnK9HzQRTwhXRiScCGSv/FJtrysX/+E
/FbLiR4aB6jHvUwMzexekfEMhJvGKAEP3y6cQSZ2sRCFVcZMWN19wY1AvBc/mrwd
c53N+hCZ1SBMuM98j2BAUEFQo286OqohqT2aTZW34dWBjhlaKIew0uppB9vS15YD
F0zBC1AJ+pjI3y8rsZV6yJlCXbH1wOIuA2HgLQ9V1jNdilEFUMGVpdeMOj/dsKzX
pLfqvGUrxebe8XMBZ5PTg02/h0K+TrnmL0VsdnqOSH2NAGP68A95/LQ9vliYtQTJ
wkc18Ye4hJPOapcf3dLEFqyQbbQ8g6B32BD+9qA7Bjvy1vU1EoakNgP7WI1GddcZ
xoXxumewDczbY39ZNTcq+Dqo8mAnWOYtXLmY50Ayi5ekXcVT+a2nyvHxa635yfEF
OdbLYb1Qbzf1kXt4sqquhru1O43ok+v7vFWjjKk6lfVu3pvUvSmdiTQao7GmwO0T
zCI+MCu2ekRks9Gv8MswTZnGGe4vqeAnEhv2NtJKlOPJ1X+Q8mjcz7duAFdydvUf
IfmTb1hSPwKQD6Scw7EupG2W0vtVEtlBuP/REpWY1Gp21JaVQjYPVnXa0NEZBckg
jSaIFpU2C73mRJ225JtIELlPDF2N9VWWlJGgYZTqsyIONBYUAjRiZQLM04SvXTda
PdIvyvnhvA9Py5cYSZAQpNTja5Unn+oy5n5RXF/qgu6a3PT6grhENNKRsgfWj5iG
/eHfvbCaQO6hxJ4VJKvTmEfDIp/RlFpQkhzjq3ktN5X840Hb58+uQNYzpc6GOMBw
gANM3Y0oKeptphrxJrKwlUXYaP4mocWA8PU6F9cGQrbA9jx7ctWSLzDtw7Yr+KPM
XOaTMTknwTS9ymyM/dRBWjJqOqXJgb46l2mhBxXELo/ie92o/TdTd1qgsu7G7U/f
rB9r+aO9/PnDngvZWvMo+CTPsZ7kk59i/A4t3OG991gRwBXTbHXEbzDOtmnz3J7l
7Ws7phfPU6svlMnyXVFnAeIGxeLDLqHfD14X63rbYW9K6Ue+jGMkxceY5HUSdDt8
2ETrD6q+CV1ktmwyWSdoFAHkgDoGo8ZVC3K3rNO55XPWRPmzCGh7oPZlueyoAj9b
myjzdFpKxTIiTwRXUSyGaD5jkv/iOU7qMa8zle483GEt6NepW/2DkwVvxv8KwAXq
Kb/FknhrbEpSJnWrfdQdyh3m253Ca3IDBftrcLVoSQgW6Zh9LzotykVe6y2g9abu
vziDPWxcjBhB1vBZKZeFgZ71p56I2xZMWIZbPMCMdUIkCPpkSDY2gejfQetUKvbe
ABLXCQs7654EhGvxpiNx3LIWNWoldF/JeIVicnO+8LTzNm/MsM5O+W8CIODsi+dZ
Ed8+A5P7i2YfM2ztGGNXIgTAujOTk+g6bAALs6Ux8H7iu3oQEWhyqRNUbwgvjJ7n
JmraakFse7dWyu7UooOvICS5PNrUo9ILlfbshTC/45BVHiHuxejtLuyYO2f/bcgq
JxvEi66UqgN6kDfhOAPri65tLFBbzYK7jhy2JD5LFyvZbMOUqeipjPVEX3zqm6uV
iHj31UgeCC2XrUXDY65QoQHzh0ndLEXeGUcH0H/seh+AD7Hb9slvIFX2DjOYU9PD
DmVjaWfG0RgSGIpDAYJBW9Q6vkNOrmpeIbpqXPMDxUIHbqcAv/quLQewkTFgj/Nb
eWw291ZmY7v5Wt0+35JtQh9twt6sJ/z0hP30gJdAZbJg6rd4owI+jgI955+MBnnH
O8kA4T0A6qJADF0Bo4yn0kgobDC438SKESRSqH7Nt8Sf24sbwYgTqKsIfs9qURQ8
JFyGAIeBv7kDHcGMyTjE1ZwDrBv2d1Or/5oyODQyDwYQWDKS43r/I9cXPeShq2Jy
bZWdOdeCgUQ+bfkWZWdL+hdFLsBcrS0L1uveatcK1qiACqtNjSogBf35vBpRQjZQ
WuLNftF34ktB0LOE8ougPKL7Ahxg503oyvIr31fo/J4GYoZ+/xUYFq8aTFnL3Ds8
6eTUfF6Iln1Cfeg878IO92iy9xJlkVGO1o+upkvRvn+BFPrv1cAPA2KVmXU7NAJU
jPI6vvSgYvmbb/luYA5wvh7+lO352QeLtpzqprB8YlxVzahJUM3E9Aje1Roxe1PC
CLhmZMNJ7tHtcv/dB99CzKpRap/ceTCW8mlS9tvhLQhx4Qg/IZ4kGoQ70sICcnq5
Bf+RD9G4IK1oXAHGRI1LbYSR7qDUvv7EuqW9OVia5697vlT8ktgWOOXg3K7D7Sjz
1xv09btT3BNIk3WPOjLpXSwcEqMb4Oq7E0eBVPWMhglAkpV2eLlyq8F/xFUgIEFQ
3E1RYGwYfkgO+aeC3cUoKyKhrQ5aYxRrsSuR2kRIsHwlpJV21RG5zIiJUry+yP8e
7OxV591atVY89GbOK8sEktCTrCkM2QrUYMHPkqmGjznEBgkzAoVxvgXCVv0eVFJk
p/IdNGma11JRPtarCQRvo1QMRobqh7YHXvKAVi1uUmp75GQbreG3o9l85n/OKYmA
B9KyvDKxmORSWPKaZH/0kD5RaqNTH3cHnTMoxvLs4FXZWmwJBINOJXiibIcMMChg
Nktg+E94JlVisqwNq9uehPwuKZAjqJ3h1H17FxCCq9uWvan7OSdE8gEcbnUG8W1a
h1Qg9MRpZHFMkoY4D/ZtJ9MqwzoVLhmCQe7AmiXkvqm599LeQjjiYZEBCJZEizfS
Vq7Nv+W6cJnYLLxRpnkIBnRhW7hEoCdkiOBPqrM/LvvDZNsZUvpEo4m/jIHGdwqL
5Z4hhDLyNSZFKbJhC1brMZ9oMiL1W6/KmWvk5mfUwBFu22st5zac8+fd369Dw/BF
xueDaQgaHuv5lZo9Gms8T5F2uMvfGScL7VtR5/bkfz9K3HiXTYY05Y9i0bKy3cv1
bRSuESbXlPIBOKzeLWvHz1zcSbKnArrp24FFtXFs/B67DXP2wkEK9WlaPWwx6PUx
di9YuRG5yrCphHr0D8885n078YYclRqXszor/iuCbZftoxpk/ILkDsj+IhQq1YXy
xsicu+Qf30P8lEIlufkUAEKaDco5GON6egZS+TG58eaNYA1ZklkCNUO/5oqiwHQ9
+F+YoyVjz6naUSZ9RvvWk5YEjCCQsG56K6Fvu/SQtMHpCHrNFZq75n9XP3Lu4faL
YsjVvo3yJ4XXSTjigGUUlkGH0cKUPmh9VTBs21VNLvHh+fLz3r7ixR64GPblnOGo
Vi672eqpDJcngVyL4E2S41hX8B1GV7tNUSNjnqnzCxshsv/1b0nW4v19ma6yF8lZ
6iXAXarc6JKFPbi3p6bPuOMraLYfbspMZz5C32CGXRB88tAF/U1YPcihZqPQfAnb
2FHHziFGAPuD0xd5uBLO+4ofmijPyCyFqUAVdpQvpym1TMjypwtIyE2RBsxWXYl1
C2pBcWlxT/Sq1XiHRL9v+CW0AbIQMG8xppoSVLfaAeGoxxAEZKlp5nvAYxsaQOR5
RayZ4WWfDZO7qRS3yUM+pvqvhipJefg0n8W86a8oDJFVF/DuOkxOjQFJJy9L5vUw
WWaPfJ7XA3r9xSWwXqfYDkZVnKHgYcB9DqwYTiK2BwvTa1gYBA3ANecKxtQrbmhX
ghWSWcN8VuDwZUj5RkqUH29hxREhIZYo3RZRRbetuhNCI0ejdF9eL7WxqXUqsV9S
kxoOp1GsWDN7eUj1hsIdLI9xagvtpeKwfFlVNtPyPo4NGpuPWktkKZcduBJ7gBK+
3pZulKG30gC0XDg9jePEXTpKkdwls2u6blnr+MwNy7IKPC9RqczkWVkcgOX5Fq4d
+g0aiArzRqWM0z1YW9yKDimO+q3gCoqXsUeAoep4ELFQlJJkAphKFxxHEjclBikd
`protect END_PROTECTED
