`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMIPtZpJtaiUrLLykl5foCFbIVxGFcOVMZ0yeYEVjKWS+fhp07TTJr1g49rBdQxz
U+en5e7FBbXxkflx6fkKvchNQzdHn3tWCchlFwmk/xOopud/AgtEyVgl1HOixW/C
K+0t4cEZB1410LTj42+vawL/ee50GML9dGtR6+la4joIrm6DHhSqVRHh2jWIqk1r
y19jJrIeAUssI2nZiyeoLjlMCNfTFsjFrf6AfDaaKBU6qd9dAQNw8URg5utiE9MQ
gP34DeHJVpi64EiPYfPRQBeQ8STbUE/+IrQGxsjsR87zosIGkpddtd2ibsi/SZfc
mmYPTCVdcyrHfs1DVd65F5BONo56ZDGLUA6s6PiR+MaFpmoLkVJKm1vsktBAzEfY
jhgKzqHeSy5NZZvmSNTfH1crSZnRxh4sETItbMK9nKromlerX3qrpam36hledw/V
Sh0itBqfPxdpKsfI9x7F/WiHXUWKc/cTmuHDMp3OPpNrT0wRRu+IaAv+nJHClz5k
DqZVRfla1laPLT5A08IhU1/nSkZDjBCy457zFtR8SPGwgn0BaFhL1cpebQ7RR4ql
S8xI+WNFka3X3ALYmYqPh115vKe4HfuahFn+VSin+Oo71VjRHK4tISmv1gRt5xqb
ioqnsrQv7cpMuG7dARUGSuSU/3K5flO4Gw+zipMeZdiHzW0J1zCcvfgvNF5uI/WD
tGUGvftVwVJxOY7q5YBqRGKv5Lg88w1sdoTzN285V5QxyUAjY+BM0mJJjsdklpto
DLbYxVQmtzuyGrZlEkanGdKb3scZ7d+uOUlu9N0Oh2qshsqhlFJg2py6EF0oP33A
vDlxgcxuPTxP5q1Iu3pAq4h8ub0NvVmIT2dnOuyDeiDT46tK0FiiZtvmTUysF+85
Nyw5NCEKzp9p8u/yc9JZgolNTzjpBb0UTgpo/gvJxKPL6WmmjACJy7TOhWktJ5Ov
sTapkjLOnMJPIEvXEIi5ocP7/sjtjzMjv5OCP2/Wcc/j13pSJJ/6DKhuqP/5rRcV
VLxmPjw6pbIa+LJpq6ReNn3iJDEmMBhHWFavkcq7PZgNI3Q+2ret9xRnEM1aFSc+
HWpKBAAX3LFG/fpHzwM0Gu5tjTPotnjmvxnQJXexYVAR3cmJgp7QQEZoyxP83yyW
Oo2H6gojLAACQzU+Vd22EDS0trvRGdQVqjLuDIU+szfaIfjedLJ2nyN2kNgc4ME1
xUJDTHtl67Rcl93wNqQK8MaWTLAnKjHvsSK60LRrQr3JETEEYL1wjHND2tNMDrl5
GyEInFfb/CD49XGEBbMjkhMLfjRlq+JiO6ON4D8FwbjZFcsBRPoRwZtX2O9wJMnf
ynU/BjIjEsy6Z9Y/CKJRp5bv7mH7Rrr2WgM2yhvdp8RHDTQNef9JCC2L+VGr1el8
qQaTdnZDBQ8WLFmsKVI/bwjmhx+lIaSbhCx/SUtCQGH3IOrJWrDRbRORpzFe/0pZ
ZSKCUg5G0jObdNKEYbB2Zx2u7GycHFWHI9YZVJTTSCP6C3zgxLaYTqZnppGb1OoO
5dJCKdHBei20NnkIk9L7xIURFOLPrPq0EjNTSPv/+Zo4a8FspUqLdJls26ATcRkl
wVg1TaHsnSB0uv/b2Y6DhG+CWm6PiO/FI2JWRJU7LVP/3LVSf1hgRAO3NGR6/Nlv
5C1+snOK0/ZOI2fEAEYjIF8ZrJvsnepQeqyBd26qb7wPfxalPuxQuHi+FqW7kgVp
epMfOTH2J2sm3NH9mg5/wHJ41uvoppph1FCgWjf3xw2JnzwRPM3SDHr+3gyF8sff
GR1E+jLtK2+vA3BThituyjlGLNS1YKlEqkEQGd6h89IfYTdGRMGqaSSocXIZaW5l
wL6/u20h72QuraEt2kz+8ZX8GnCJDxSW6xR5QiGqDGcc1a4G7JjzN4E1eKadUnpG
fYARnrqaUb8s8ENSCPBxN9qDVelv+7vru78e5g3SsBJtwOHsUG68zghdXOz6Abtw
W4YPDFoPfnTjg95NNeIumLHxwhxcEZNXHfYibPujTmAUp5seyvLgoAi0SA3PGZYl
aYskLt5EDxbW8+cvl+eFB4W4AqDtnsiDFLZo6ao9tld34fcsoOkaTY5rUh6k3o8p
n8qcxnvSwy8NRXVHb5P0lM72ajKvsYaJqlu/sJQwrDjN+ewBiES0RDXr5jPaq1K1
`protect END_PROTECTED
