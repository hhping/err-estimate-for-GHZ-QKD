`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qV7xCg9W0vDoV+OeZvec7BVeZuAXebwrN0PzRmly3lj+bntzRqUMaifR9AzEX0RM
U2m1Uj1DA8Iqg9FZ0jVGIW5/90bT/+wwufjzU1rP73D6lINHtvTlpNGvSxrAY8mN
3EK3qMnBx9JrbpnJXSuFFpozHlTnHr8MLfdKxGsCU4/rkz7aaPPrMRK/PVmOfxmf
Tp2DSMyxJ7T63+oFUpbkTlG5S5JxPWG99tle/3uKU5pGtBkYWbwduAEpbEiw8ciT
pqGKF6zD9MiVctKoWcnnSltSwJv8Jjm/dORe5zHpXQATMsZTPiwVUuBkkGt8XDvI
kTI+XumDr3mQU6jzcznLC9UEf5uRsAfBqQ+UJLZdMQKY8C6VWbkIA34vOJ+ea5rq
yw6aYlKBfGSFu2Q1NcGc+SGrn3nv5A8fyMqbVDwgVp59ZLSIeb7Ski5W/zV0dD1R
TodI8CJ4WC1i8WU4JKySyUTy6o2pe2Si+XmQ06Uf2gxYb+rFtpAFLuFLaO4KgjFi
Vdk8PGL+x4pWajMct3qCH78VPdaRmQClQf/6rSzQfncodMsjlFPUN/MDOqMnIxua
RWwTYcF8Q6C3+JMreSt2qJ3oiuyF7T3hB0PJK4ZjyDj0+W85TGPj69B5gGkH87Qo
/GWshL2p+NHg49kordjvQZx1VBWtTXPjwJrbjMf28G1ijmaHNq7cmkvnXJMdr0bH
3OQopyXmrF/eP1J3zKaP04Fg+fOAR8rhMZsXQulZ8s/c5zHwfUCCiOVevnKUJSAg
izJ1S/zdudldU73JVfQBVA==
`protect END_PROTECTED
