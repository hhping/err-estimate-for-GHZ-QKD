`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5b0WPiaYkobGeAys8X7FsLOeOwJPREftxCskInRjafR2gUQ1Cy/bYYnjCzBFc3zS
ZU0wXoitvi25rLI4q5akzxRLsqFQzGssTnLpjgFqoUxxN5Yvug8UsnYfK0NCRDsa
T9ZEUV2M9Vek6xsD3+zkyeX/3r9k2nxVHOB76/KedlxcShmxofv2o19xq0C5HAa0
RUNuzaoe5wQgRNdlx6HFKgPMIL1qPPzokWJ8/qVSDGZoahzK5dKd33qY5mOtDLHh
QzoPI9W6Nw89yJUCtCwIrR4uqj5KI0bOrOlOnk49w9gMn0sAAk6Ki7h7r/XQDA87
K/iiVimvoqpEPR9bMkZMLg8+Vhjhl8BIkOhumvE7aCDOdLpuIxxUh7//be+/kohI
OjN93tMnoKSoyZAD/NuZKR/PwgbySNMAvok55Zb4ICn7aC2yfDiPldU9pw+DfLcO
NyUaUvjFDIOSlh1kY7jSRqn3xtp39vKZ615tX7QXbVKqn8vKBWid43hdZ5DzN1CB
O8J23OZalVmrQXKOGHpbVf//y39Gu/SE70Hwv9aeI2myRpxfngVJS6RezNjsbIU2
eXQ+0BwQod7UabWfS6N5VCGefB+vJcoIuOEFUWcHjGWUBiBFPSCOCGP8TQB4kA7t
Qis6O4aJBkZ0LvoEdGJq4QzvpxgKrXnH+vGuzu69ATG97jSzFcw535hjjfuOCUAN
LwwZsO0RYzC4XTwTyGUjLNN8nx9Xj+kSESQbqDzk1g2U52JpMPntjjh61mIcYqbt
r9DOBTwN861YL+oW6rflkxIse9wPoyiIhuvkjebSMQMyFJWMN5CqD1olCxKyMRzN
cSewshiWXg8NuH82oR2WIVXrhGnJ2S6cVvHiY9ElQrkexsRCogx95w7nYqsYXbEa
MJ81UuocBriDeIDktncWod9pbCFYARGhlQ2aAfsXu02x6Ri7TCwSEiSfYV1gLK1E
l+8pLbtdbHALwmZD3J2Z/APmkKv0sqIw4dsQ4mTXc9wRy+tfHK/52ga7U1SfblsD
etMCShdNF0ZVSoruCqHWebP8GtdgpvqwuZ+uacTAC0dM0mRBB/Hzo1xOjKhITgAm
T0LRpgi5LS3HXVtDgv6SZpxqA1ZSAnhSBRss3ULsVhkCBkerT6VEONisBHrJJPS4
MIU94mFApD0xK8Zm+RiFoqxXcTvNop27zuyDy+dRnokrgmBc8Y3BjJW2dXdZxsHi
ckYGvJcZtIsaXJDmVa64jdLq8svfiALnyth4oZt0oNfXYCbMLHgcGprm5WuomD5E
QX17EI1MDemZ4rDMeg91SHt5oOe9BScolQHZ/+R7fV6ZEgWfNH3p/bCc/vku0h81
rYYo4w5FT75ce9aa2mDRsBS3P5cx++XJnXl42js7kC2ErCsinkkzcoLPYynrsW54
S8JJp/RQTfhrVdg3Qjc5ISUg3YbieMII1EgTpm9mdrvQPh2S0iwQtXRup7mfKdMQ
AVmFziKysKEy0MQMMtZR9BGwknLrvbmseqoudfR1NVnqkVlvSXKiS0eWvNwWLnHQ
O6Ch7pnYkuMPaR3vc/uxmzdaqywKviEJc4wH9r/Bsa3rMRLIK5HFD7oF/PSboo55
aJqhun3cBoCTnEzIHI3qqwY2zh+XNkJiY/GZbCSAPktrhsoloU7zYjzIXsgjmjVl
hTZ69rNivMN+livvoPfvJsb8e7O1qpY4g4aDmEvq8W5a4N61+IWeCYX5Smc1Gujf
6TPFGI/+5G/Am0OHVC/bX84Kx0hOz8D6YWarOms3s73OfUK/M47p0NchdX4h+rEj
Cra5EDizr+pO7kQ8pqBPBsoN3dmWWRbertLU63qSBxb4VuJh4YI4yqwEPh5tw6fS
seH6cP/VGqA4f4lqJaolmdlab9H/g2VLnX3Gz1ncCPqbI3YIf6IgI7J/oQejUkwQ
J41MhGTjKGP/XaZ6iWjly9zV+vE5t4sT+6Qg7V79C3FnuLqVgFdWdYE9dQIlZx1h
b3Be2CmueVDSTTWctXJkMS9iHwTEX0OFXb3GvcopuSxuNJlVx6+L3AK3K/FJhTJP
50J9OnH4Q/aPpb8jl99pNrS1IN3VEbf7Igf29E/FVQCyfYm9tEZbRVCKqXHTl+ZN
4C1qH42P9hbGMzaGcmICKky0PONfGGJp4lGKtn4xiwabY8bjdz/Zqbx+vL2KNgVP
EHOmcTWnjGnWcqyUK5dYh8ekyr6zxnj40peJMOSnngQ78GOsg7XTPQSRCnuRbRTX
BkTPHiAD2klT6rYvGQDmK8osGb+TViVMvREXa7fFkPGo4ALAJMYfiqaNSdx7NRGv
dK0f+CCyG12nMTN26MaJA8Dvu8k7D6rpfS47eo39ZRl+DjkR5oFVoBdGW9IGf1Ay
9jCFNCkgKAZKscFFFFhFwsuvJP/KlqUnWSGvnL7wzxFUcDKvjsM0BDU5y3ADbafs
kL+r1Q8jIoZcrQ6/4+HSA9s2aiu1ozV57ZVW3yEwQ4hjyYcdz3QoPTac18oC++s5
/wiOtaHW3hk6SsCzBrpukFux2iEMCdeHBnjKep3LdUN3XKhESNrta6e7iOWk6CTm
sHYUQKEiJVAuhzn1ln7Aw6kdyQeX9pzHFnQhwMxe1OKuCD2/YzIJWwKoNESog3Oe
ZOpA7lgBi2IojJ0bMqM/3VQqiuDKbdpulg8Ahh6uCiYCqrKkWUBDPaCFMG3NDx1u
RVf/u02ua1kt/j4pbZZRlqs09fezYaarW4EODyj/xoCAtOEJu8NcZGILGAPy5GYD
2OEBNOgJrc4+W5xjpfN25+u3Xe70kBuYJ/u/E3joVbi4hk7OnHjPjqjl/SUhUNOx
u1toqAEh+3a8voh7d7HGP/k2teG7bCsKY5w9dsm/CMEcBtxsVz7ob3pCWw/b+nbN
gDgW2kRAxuGPc9E4y7KfwWi6QzHMuN4QOiGrey015d4be7XLQsbUH/bmMOd8kSS+
8mSCJAs+Ar+NbnInHsnrLiEN3JVby0gf/iE+CtGid7uSsUIETceVa5WiOm0vLsBO
Lulwf29q/JAIdmNCGBCkpI0AJzzIcdSxDHgdrF2QYNed8l++p7Ci05YawDKa2Z4L
tN3mswNYCeqRkD8qHnYuKDzWU5iP8JWNKpjZXqv8i3fRUPCA75rHcUMeouHj8Ffy
HkrF+2YVrgzWAzhxUdP4ZkfPtOcQNsdVuitXV8/KKc4aU4nseXnQEmb6MvME5Uyc
JMazGhwV/YQ0dw38UE0D9RHSZPZn8375jOBGRH0vuSWU6Wnj7ej7Jsb598TtxUh4
FnyNHNPoRlJZXbyDWA8F7gi0aEpKDoxgaMNa976tytNF6uyaT9ak1Kwcs9F7YTd4
qeJjy1AGpE5Iawk4wdabcICw8xlNDsvRUs9WuWngu9XeZbuUJn2FgGSGF/WLaGMy
1uOf0sc5DbShjzT8pUV3iN7y0wX1cGfD/r0XJn2YnJynex2Q9nfRj7rSL1HECmGO
PjiDa2KCSGhEFB7BEnO5ihJ2Jmn0q1DVHKrTR+uJCdLW2N3kFoRA5AmUxerIHHQh
1f3+yrqdQOpoFTJ04bja5KEpa3DJjxCOsG/pNXwkJNmKGuTovcFTk9DF21bSN2QH
c+u0eeNQGDeVQya+KijzsXP6uC/kb0upR/kFRxqdDcPOGIRu141wVWk7wphRHKXD
z3nIJgMtnhianKMFshdpXQ8le75oY3fr5vLvtqhZdVsAMriMAmi7ifZWUKthYCy5
k9FyMUrwCdjmw+pDewM3njVaVhjSaTyKQ8zjnTS6FRj5MlNst/pvpe4XumEmxoDk
Wac5osa1UC1N7vf19YvMFVSpLvtOxxA0AesZbl4vxyp1n7k4GrYkrdbNNYhmYJVo
2TBobn+Xnnj1kCKZVhqHxvmoj9Iv2gNmWtMP7xbKlEflcjjJamusnDDjJOw4l5Nv
m+DV8klXzPfPxPLWJArRIDgeOaWsoE9etPa+r6pBeVXasxwdpG5+ivJ1svDpMTPl
VBiAcXTGvEhbicObmCFMS6oZ8jfi8ZjXSw/vesmwVE0p2rFw1GTErZnsvMQi6c2j
JunrTuOqZmUh2QgTphjUK7wtC8+ZpT5EYe7Lcnl8SwyiZCM3TXclaOW5uks3/sFw
1uUYJBSFBL0pHpK9vEng0amAk+drGY7oSNo1Cq086cd78ukN4Lta3yYBm05qmOVI
CpSuokv4qTMOf6K+hFFGAvI5EhsvRP7t4Cm6/lXEByjwKL5PC9ubdJhUbP3fApyO
Lei2GlobZGSoKUUPDpvJhfOm28hBQ4HD2ywdMMo5COu8a1QRV1ObvIjdkMIFjYL1
Q33NEfHdhPOmvQLSG8h2DiDkp/QOTf+uCtQF7gpdPx4s3rAsDJ6tHZ4brneF7yXQ
bIUHr9VCXtMP1AiY0mredxgxwwO2EEzqa9HTsSqDUBj5x1pHWRp/lrumC8u3UPmO
7RwSu2bMYNPJoRE+9ydfYiMJWL9sWpkIsSENolOMj9ieZSk3kCTkqlDCyKA/8x3F
rRU8KmGBgXdz/YPDiQh13SFfnQwylrkjPofhfP8gPXtRU6QZwid+zRyWi9y5GTtl
3ENcIhBG62R7KLth4Qh0Sjny9yjWmDFVrnnnrK/UkpJ0WBfwu3tMJ0EH3PBr+rq1
MAXOTYOcJ1jpfeZem7amSObofMIvIwZS2begQeyKvAWFxB1lOcR5qvnqQYeg4Q1a
TkNHmT4rFOdtzVji8hm29cqJLmb9eBriq/msk+44UGHBebpGhleFImickjO69DNo
zWi4X2+8bnb5VG/teEFbaXatyla/lZalVTQAPT0fZu3vvBvNDiu+WMuCQztwKS26
huRSRkE4Qmhqs5sU1WfFYtTZoKEZmYSHZikm6DtkDwx5NBUW1Tl90cAI0xvllk/a
Z1wCidlWr1a7fpcVkHn/SxtDmn78uWcnuAWP/uczO6xzAPK+d0G51hcasFhvi1LD
A2THb6N3IBSR5bQHkWQl+5R9ZtEP735NXIUX+TKkP1vaQcK9+/P+l0/rSLRDyIYb
IR1UEPtVnZOjKHlrN090lPaUrL3wyDoz94NP1/cbgTpOyl9N9K7VA4CLCCeijdbU
BgVTlaLVgRuUNPRvEpaBCvV4s8YdLVNHNP2sWUFfKjk8zCxxK0ZHV4ya/6m7wHpQ
rwSjg3P+LRI9O1hDA+JnBqFoNiRgZmgRo5mdNoWUFLOhZDTweV/ydqnVc4nToSID
HbfYhvhyZWAsWoG9aARneZM7skyAPANZGa3AOzCjkMPbvW2xnJpde9MRq5DdwtXc
cH9vX2DuoD5w2DpW052QX3eAA3BwkD+sP9PzVQsYK9+PR3g32FxTIW8USyuc6mr/
EnWDB+PXhsps9yX5WkaL1Zb6tSOQejmNk3QZ8b1El+MX31EdvQOM90HYJXHCgxRP
t8i33uFJjITCb2x39LQyDMlX1ZRstVI4nWTDuHVYAxNGb4MLuP4hDCAuWn7rLRj1
QYM51xCsFogiIgouEY/nfgXs0b4k8Zl/szqNYyTaD9uXJFQrGt3izEfu3Q5S2gEs
o7VFCd9MBUbFGm7ele0xxF02J/6i1ZO450TCv20fJOZdVlXvjCluKUpqedhFY4Aw
BYTpNQizoiId2qTpdR0ie0rgrN0P24deWU90dYoXsoKuA86C4KabKOgcrE/TP1TT
ybC/wUui7W6I8/ESDTMXqspskpYuXK91bzPJtE77gI5n8ShcjG2MFtaTb0gGPfq3
BhXA/yRsvkfOy21ZXYu07Afiu3aoXDx1gIHfQKfeoZk1YQbZMKWc7//qcC07gAIU
LBMJeu4qRZ4u4Jp0/X5SDFuD+iDuiVXO2Ec4nqra8PX4DoLpTsqydBW/Y5AECPVx
es/+hL6FTq1d+3cwVmEEZz+FfDYTFLltE8JaQlconIq38+WUY07+YGiwka1OiB76
AQUZtWNft2r1L60s7zyqkPUDT7c5NMsI+/4NzrSsa/fEQOz0MlfQdoJhRX27R+Z2
Q82u/4ixSh6vW3zjGngJdLkixBAa1NA1Uj7RISDe7eQmuHNQj2UkgcbFGCChpAj6
OZZEAIDUU63VWEdROOEVF0SJFWkaU3saiIgZcQLVB1Vv0vUi1qqN+RHwWAotrNc7
lePUSTptSfMS66khCBUWlW3QRO6DMuS3iRnukAzpEw8QQNG/4QcDP51Dl7HC/9y4
nMLeBbYBRDB0LkfP4KjzYX+HNM45uO4x+GAqK9sWImSTgVWX0HAxd0Tee/fgiCm7
+9Wttkn/mPkYZP9YywC9rECROlT6UVbWUR/KrHo4GXShowtBlJLYNBST4goBHp0W
n9qvoTP4lwjs60ufoiVAbY/WTMYUHmOadIBd5KsLr6liK2SNGel5cukk99+jp9tT
eDIdXQJvT2uz/Sul5oyTmbM3L8Y1k8Y5RxZCIPBggkBvZsjsIhxKsA462FWJq87Q
kDCgDbDVwqkuOrYLO3+AQtKbNFvg6aIYIZzhEQMdziVlo1pNMjW//oHULg2u9JPK
spva4+w12iKOodD3cTLhj+dJVRvc7SsGV/iW+6uvCzoCVvZ2EJ7YJbCcYv9pC5BO
fPgtMEfLqe57AgsWsGh1ClLj9zue78iQMrwioXXsY5eBubOr8upWBmOu1SvbDk+a
NOEaRKToFKq5bb5E4mj9skvVdiHmyRaZNlzJrMHuQombIFhupCbeOgQu2tK+gbd0
fvaWaBA2rHbTnA1iQLknhbi0dTkqwgWBYukyQmxklpQl+gwTn7MTKcaU6EsNKUcS
PpUi5NRD05LM39p+5mb4AmQhR8Xa3hus6CyOeeK9Z29GKFEOapR0qJvhiZHnv50b
ZQLw2xEKU4MFjatShzovaRFBqTYn/drrMDTfDq+5+ZSHbkQRW+19bRzI81KZgW6a
wLy4J2N5Qn7DRfz+5DdwxA+VrztrYtLrXe7tyarPfjN/6uL15FybCHtgXCj//u5Y
7LfWRAuMGVgom8C4XgoAORSLe7n8gdXk94wFy/aPcXTNwb/yELAjgA4z7VCifD66
PoocHw1jrKhJSQ5lmQOpxb7nxrEo5IBl3Am6PgU7FItMjrdT2U5f0lnGrNvk8Mh0
FtBmNcte7t6B2kcoKC9R23l49reIsFRiNRf/WL1HB1J2lWzzO0yE4Aqc9anUk7Dv
VYr9A9PagfCYt3F92b1CI8agQBsvU0TizKEmiAq8wz2f+tUXmiOYQrTpFkEGXkmn
6mBl1yY2n3oE05JwMYxvMEt0cC9xsLk8z2FVFo+7jErRjWBFnSW6TMUH8e/Fkwmv
TLxO6CPAdRm+oELUtJpjMIrVtrRqrlWonQZRE5XtW7Wi7/XY1WMDM+K8SQ5Pncb0
RI4MjAEohGntzY2GaUwMrxb/Vq+GEAYlsDwM3pOuAxayfRpZ0aggEv9eOPmXltzM
Q5Zlo+kUGEgN4tbI+wYbz6WoQ/DRq0yP5+FOCzboa+jCzUvLX7m1NOuUjqFL0pMX
x6SsB7SXdiH8TQ59hyX7WO/gSLVkflzRPd5/dS33toFS6g5lxlqzmOzKM1p96R9o
NdZ9SqpprxOOxBXMvaO541IK8DmfgCSHlVgRVvG+h0v4BAX/vBrU1bK9Z8GfS3NL
9WQBu7XIg7JVylm2gVlWLVCtpgGL/M28xEHalTS5VTMZNt3748BxiXqFC7xz6qhw
UVcEeqBZjFJu7mmi6gG+47Qpeqsq+L/VoFIXDOgPl1Hoo6Bqt9ceCKexPCu06+fk
IegOSHUBei9SYZresI2vHJplGBiQM5XZTWHdekY0M4T38Q0fMRa7l4InBYU2ic+X
Ks6ttK4Ghj/2RRyEFBkD75CW0DX0bDbzw3aHCHZkAdt/z9OmAOmsB1MNQSFRDFPh
uZLuGZD0miSa3+e2iX8v9fGYVpnEMXO+8qzAIJi3QyX1D3xYPMr75esBEhPboOcY
+Dt7UGqcIIQBX9ad+3zFG32oNbRurLmx333Smuo4OtyNJPlq/gNBJ0rddXfEveni
mUsd7sbAuzlyZGvZy6ylkRIPMYoUzLHi6KYhjM8C90aKzwObn8XBsifAoc1sqNmN
tVnh9iMq7g904Fmb/ejkvmKT4rkt5Wa7P1qWHAI331q/PupCDmXIb32s3tiD+7/M
IrE2IGHD/EXB4G/POHdGruuMX0YtQpNRTXWXIuGO/9AvtLN8FLTJXwUMFmxtUIba
JL8w3qS5AaO92PpJSWiv3DRFO3QHw95lS4+l9QUrJyU2Mzjz0jhTbqCbS3dVoLn1
U0pqLeNXT8TRm5CWpHZRupxqJIN8i0qv1HayMsfrPQd5ObcmK05/JxvKsa9G1rAY
l/tkkMoOAYbD6PkcAFmvddudkRM2t50rVyIeAdZHlByyKXWxIuE8JRVeamhr+dor
CYdeWOKjsMYP7uNQidj72kA8oDUTRPm7Y5RcInwzkOKoQnU61ihDykEmsz3lKBOA
HYMNGOhDQuK3H5QD5hvsRgVXD+YsIsKJETd4c8Z6hRs46VVYwlUs0T6jO4h72VLq
/tlLnfnxgi9zQzyY4zacD1Qb3wdFKVD1/LURMlpYr9/BUCArsNhnbSRsVSqeZoSy
O9AyaHC2OYkHwqce40DB+DAmvVIgvWQOVMrgr6tJJKTpewlSbd4ivck7BDwmJGLG
JbPCaxb0kPgSgmTHVy5o0i8o/gx3N/fEMUHNARIdgF8mF+hPk79pU4wRoh4GF5ds
023VhADDe79sqWKfddxn3l9V/asFMOTAJKz6U3lh9QEUcByNIAIf9guL7x2lk/Bh
mcwuZG8t0iRWTvcG9/6nO6Uc8cFfU26V6XN1D6hpv40FgmJPt054H1MNDHjE3Z3W
c1AbcG3KqrxCpekyRtkJD3YRhVzEVcXFOJAaAhxCTZBhxFO7TM0591jFYwfpatCS
66cEU7ByKPN4L1wLbP6mgTIiRBQURbN2cPysetgvMz6CMnm6EemaaHVHQfzOq/0Q
zGNFit/Wewi1SE8DbkD9lKZYVcgwLgpyO9G1/wS7H+IJ680PL7iMckusQkiFDzW5
zp7Qxm+zsOcsISD5Cp3FSlrDKaMcmjqIwJUASww/S7P4bcoq1hkU73F0khpMbATA
XZsYraLUCrvyJOdJqRizqxyRk/VtN6LUSwupo+zSuTstfzWIUJfmYojFmzjuvxdj
ruYZbn4kctuQCTHPEwm3s908dag9atO/5//R6Usd93+UrW2K1LVTeq4H+h4NeRGu
IxB20pZgEDh62egpCEvi6Q0zaE+9+aMRjPXe00VQjhwFQgNGY1PHlPYXhHjKu35w
/2JSfaudJeSBrvH63nFaqLT+4zotAWs400RH+V6yKM45W3ha5e/ak+G6Mxx+jbWA
tdRq4CKaPDFW6ppcC2RJLTdEhnV3QbI0EkJeaVEidp3prW5+5QVABTd5qgajsnDC
H9Tm87NgG6JlB/LhK3GblmmIg5z6DvDVzsDZziDLdccD+mN02pm/1e1iUfMcbbhe
6fA1vVt5Mn/B+7QRhpbVU41Iu/wWcI/CaHsswdW0PS/2j39mGAtA0OO6EYxKzpQF
1MP0ypB2G30nYOqpNELpSyW+tYMtpo/EOmKj9DezCWDYz89NCjdVMoo6hyVH6i1Q
RIW3Z2NI4or5k89OyBKNM2NvmSxdzT0aemk0qAArxDsghcD8ZmIFJ5Th3w40+xL0
08KNYDFzobkMco5Ni63sHMbA+0hzdV8zICdQcRe+RPtSL1v71QaE1mj1I5kd5uEG
BcpVPr84RY4buc1vazt+d+hIL6UVhfIaAz/xdC0pyOQAySKLb40TR75b46LwHCYd
C+T8Bgv9RAfS299Xubdrrsp24QzPlOSAK+m9rmCmY1UGHDQQ8VQN8q4ZDJ3T/ba8
VGpBnPZotJm2z3UNMWscgjihfdSCXJpfOhkBYIYOvvJmadMylOTv0iycv+5O8uro
Jdd5MiTxdgKCL2r9jlr3POmHrBLXC+Ne3ljOjFdGM4o8T2nQ9JQPkySuwHTE8eyu
LkCc7YH+mzOYALtruI1mOGhnM1+NwUDPwSYy5/o/6QH3V1DL9jYkofhyjz8xGm+n
33YVkqFQoJzr4k/5zcHJR0dnwvvvzOSXbX5oWpMfrvG4AK2isHPqASQImjAdjTzt
VR1iVM+3AJW9Wwncw3W2De4TR/Y8U6JakRUuvmSWmwUW7BrcsgmMGXmpBP/reTmG
yo9ooNqFfKB52UzpbEEvad9iHce98DKjRY4qDeeesz2yqIC2YRqoivLpF6yDw/E+
b8OiIOOYl5EzMhVHmnR0c6dhp0N5OHItLjZUKPvS/vKb4tZuep7OO8JYeRDgC4Uw
XNqg6MDoo3H1pKCubFjRI+/0tZM7rC0B9Az6W/jauvQI3D6+YCWBUb2idWzXHjPa
dq0VXFlbdkLtwPaYqa6sK3qSWofJtqL2dCaIt2Fr/3Ol3QLDAxJvC+pQ38kF7Y7x
5+A0ihAyauyE3nXupWbp3m17/xoKvYG16xtEUE8sQFSXp1yFGRZ9Q4/bzJw+7q49
W6L2pPgvs4uwSG/3OOStymkbCqsux55Y29Gg1+YFSR6r9oBlR/ljGZRtMGY6oPTH
RxnxVKobJejrFHXngfedAGwOi8RJa+EbFk45gYvSLXfHbs1rtMlmiiBURyPiDFti
tOaI/pdDCEQ/9KOF4POAGkiWOmP0wQkVEh0TyKu+GshUWCb+8x7Rcet0DnIwOtPL
I4VJykW7DQAbz7EkILr5m0CXnX9stQFfzfuq/M3WJXKdU3LAbua8fNxhErc7R+U3
XsQsMa6MFVED60LAmwAPfnqlpQClW+0Sh9XyMfjkYpjeGanHnewRX16LyWcsvTpt
7BUrCrp5QuoMtdyKTWw2nH4+ofEShAvDZqWe+zfM58kxOmmrQWprKWZiU8ueMAlL
0mxN/xVuiNgNQ0v3JxanFaaGySV9cX9Kzbmc96VfpTOThXjgZvgphgtpYrXmT4I0
4fVALHhByW9rrPi1gkxsKC4fmJyCLXOP/lI31ihhtj3i4xI0kiwbxXCfKLkrjoDn
ut2EyWacXbUWKiJnjHqbSc+gAx35pTUEiS6c6P2QBh5XKitAdYaP3U1F3WUMjjXQ
t/sLwvG/nQXETWqJ8PpgIaDHHuxgqRhSuyADGopwTHmrlUAcam9HQm1PyltQNiAp
4/veMYvYJ/dVAU4YURNrPqcyGMfaLUtM8tM8rg8Xw66uE9GN0T8KouDyKyAxPnrt
ihY7vzN7HQTqqRyOwppwMVmP5YL0XPzDkZfbETBcfyrhnOmaWQu7mgiZTsZMrrtL
R/HAOZhLK0LjXGVAwcFHRE7X5UYQeNBm9UC43mRNBd4YRv+UfS7D3bp0dmJeg+74
cjjgXlIH2o4uM0TN/udoOU7v8AZ91bAV3tw4GJAJF9Dxxc+eaLmdzrW6XsTYJoSj
qA790MqqYqMQo5C9JPySHkKRzEhYcr96il+pHHravJ9odDbR507N10kpD8NXbihQ
N8EoB5UR2vdjqNIKhQJwrW7mxs1emQ+iw2aCp0I4z81bWKcJ/UKeQR9ftPM3N2AM
fx/qJ7Khy8W8TMXs52xiWNdlYP1SKKUMgLEWpGHIBcVZmN4+lhalDqnzlODUPrNE
lxBLJb7YYGhz2+k6NnbxYtAWFW/gW7OmiwBSvkoCgfuXvSTCUcx0f/ORZZ+H2hRw
RzI1KfMopkX7mViuNcDKZ1Jr2LWklbEXEpEnXkNeBVGjts9gQs+Zr4z4xixEgMaw
7G+Sw55CL9PTtg8G479tISheLCAJvRmui7JWZYZYRG0/fhdRFqL6ayGIz4hf7G3U
CRJ8OHBXkAC4X59dfVXFKwCrq/JanoZV3UoYt6EIXdpVgd5azMoSJSgHnGe31mvO
OCjq2ceWvDY4l3PLlU1Vitm0TH9e7DDqkeDHZbMdTc4ni8enbqt7cL2ZvWOPEZ7y
xL7Ab5O2ULglEUS4Dgn0Ak5hfk6+EabuQMKFnEa4GEVZzaUogRWQp2g1Do3FMi42
X74xwpCBQcZEDI5yAD44wn2q1eXP0FoHZA+KuDqaUIRlpz8rgfliHBJEc3HsamNd
K8vBRCurA+6VCR6chKXncpGycM9Ts8Ry+Uh1PgGzqz/SjUEXnFHfN77H7uKGPRWJ
hksXgxDhPhFrWJ80BVcM1EshFyzuxite3Qwa9HreqN855zPtLhnSxWG7G58qaSmp
edQ8PgNDI5IL4A6REo5ciRs8sN8MvrkvelpDxiIDbid8zfaJaxYu138pumt6K/a1
XJW9SjLM3Wwq595emp/71fu4bsmMQ+VTOr6lhGJyElrUim8nF/S8VPy+N5QXQHqD
5c/eR+3JHe2Lswjzly9axZNmaPbmv5qmpdGhlf04JjfowZWqoK106fFIgId3HWD0
LDltZrG0U7mO/siBaRlzwQYYsHvMMZVFhTS1a+bnGWt0vzS5uzGuII98EZSU2x+i
15lqEhWnYnh5l5q44JHPt5E4ZjS2qxpBBk+CTepENXCuUAZB3jQFwjrw2jVQBPU5
5Bk5kh/gfkLAtP2sP5Hom0rjsivkgDUU76zQuQ3pW9+JyZCP7qXFSflhKkC53+Wx
sOCpc4tzEqkqWq57GAbg84r1GAbGq0oxYKhl4jHhKp8zYL3yWMAuPw/8rlKowLxA
evbhB2eKSwh0u25lqalBLAlkoCJxFsRqLqB2HrghPmWM0IQSQM1JtVspFT0fu+mo
BWOiL/sJdVbIhZuiF3Rbs28XIb7ECpLms1ccTYyLmJ6EaX2XSwUc4Gurg3fvlM5r
sln+wsbWWaUeOHe+4UCgE1jwZV03llnppMHx8OtXhf/gEXamCX5QlmzdkF0RSFqD
KSwCTCx5tYsP7NxvAeY+YIJem+oken6ICuF3o0Ts9nfPUfMFS9il+Fh/6Zqbgm8K
rrqnkMNbNDh9o2PCEbzS1JTKzA5Zn9o0kF23xTp7ERcU1FYEll2fiWViWRnQUXT7
fZNYYeW2mkXxkM2ItOSF6bo5PEdz4lNqJ0bm1SxV44lOx9Qh1YbLUIHRYqQyCx7s
+clSi50asZdfEz/IrfxSes+EL8fvHZWQplY6ELvj/SghFraJfeJfmIevDtg2r3fb
BLXMRA4r57a4GqrtfJZeVpTJy+lvTDzD0Z2AD0vITDQmxID6v7EBxqC9WmpX8FbV
bbQQMZf0SlvFwr/t1EKIsEk1FK+5FAcqcVD9Lk/KMGkhHQnn/ho1VPaGU7afVUov
E9wZFykjyqSj8TL2n0pmfPROK5ISJKMAIDy15Cd1aoqMhX16d8KRMa3HbtyaPoUa
RdhdV/6N6ZWOJfb8QIdS4QBsqvP3x4QlCr6e4Ngs0VXQU+0NEbJmWi1tpRCtu8uw
g+dPWps3ZRjy7HwTG9g9bS/yXZ03NMGWy+kD/ZXGB15tCeGP6sDPKWHX5YQV79wM
SjwPZnXXICnU+JIovoaZ5r75jHfzuAUgeFBciISAd/MSPVfkFVFUl2KDweejNyZg
3nFZfjY63dT4ZumD/wxEAv1eBtD7H+xdI6AiKfsCIHMLn52dHUW5E3uOVGjzda2U
gnQx+BSnLTKnWWEFz77ELj+xY38YHlqz4gguD0roB8pllwaNNiNjSpNSFWb6BHLF
C23rF145NZpcG/3GZSuwNPIaU0oshjp10HLPwsAqCzjfPk/98wwzh+d1FxRZWIAC
+k4voONcsxAi6YPxwz5kYh7I1EO5+TWuNaTtFzqg0lNNO+nAe8+TW2/+ePCPPWNh
hzv6dewMXoK24am2hi3Czj5iTibjkf/Udr6Q/rJcz+/fw/sPZ960Vx80o9dELMfQ
ppx6s4uhIdhxqDltihshbF8+UiKWFDKDULcxkkHAIy9PaYzUBo6nuUOtBci8fsUV
yZ52izRnEEpQ8+YPckRM6z+BJE3yalsCMrjitjlzRSw0H/P46KwWoOh/7BGCIP2c
rohKaLf2buymR48ruU1mtUPltVK1Gi6XziAgR7Nzjqw3Vz4CPMvVEtjDE5SRRykm
0oGNw8gZAQ+1koiRj6aJDMWoAGAUbS8uAPWsNev/YQHl0z3GOZ15OKG1q9vXEEA3
0RE5LFxpbCL/fmCc4gCRBkdywey2w0OnAnjA5HMtprIo7TC2ZubWuBuh2iWkRu6u
HJ5h2BJEFnvcn0cWKPlQsmBo3X/CMVAa0pWBTjYKcLWuKKCylvaGXNc2atqdALsY
w3WPzm9/ttNR7VZ1HXpAddZVXW6F84v228GYjl8ctwzoiTNio16wk2q+OZWEvH+Y
0BGqhT3oxMKrHoWNFWAF5uLDDEog+igEYo5bQy1e9CLC+XcNfdmlK6I54GjGKCWO
dUczJ4Ll0e4+QEHHxDYjjR4aHV5Jmwaq9hW2hcS3xR6Oe+TXsbr67w/9OvH1Cx0G
k6Ojh5A9/sJvkDLepjUw6PE9zD51hDDVCmV9BidwfqbjvBFEEwii9fhEFDN4mXGg
0zK4n4tG7Mk9xBKkLEVHW0g/lLax06yczkWV7fcawBYXhEAWueEaUllevTObRpOQ
b9oArNRZHoNG3JFKaOn6hHw38hFh74vgyOF/sO+s2ylRoPvKrcmgCnwM+g4jlxrL
Xw012X83I+juUqemWZIs68u9FMA7c1ps/BthObH0XlsUY/Mne3wPY64PwyxtdYts
RtzTHKNUETEdo9s8KEJ/pG4wQ40hF0j+iQ1U0QyduYecqG6svVIFEwPVNnMOlalE
gRa6Un5TbNc0gt9HAISOiU3w/ezYcqUofSmGxSDbhpWcO/3EESy55E32HwOkYCu7
EtVvzLwMN7BYcpxPfHd5hdT+6V33z5+w3oZZl8r8fiqDA5gAO+A/L1xeOiqDOtLn
hQ2/DHUPLOrGu7vPLlnwihDR593ExCpEHoaFKT6Q0oQr+LWBqjAyPfxonpw7NbD6
jfbrJi2bT4C+Tkpxiz57voAXlc40jIjxBOpP6VSWYFnwc5tqwvwphsHRPms6lN/F
TEvD5LWr1+rgr+py7LVfaLuix5OQYtL5CnCTGZbcKYfNmkdx5eLLi4LWj/6ROKHJ
4Sghts0xNw0Nr09506OL+nQvaKCMLCup6/gS3ky9x4CngH3oZoBIaK0BSwRcr57f
JLonKJs2N330EMrBz3jl/AgdjhHiGPcHUdr7MKiMrbPuLUAL9fw5Z5VuJBC0IVPU
ASBSqI/xEA0iVs+6qO0V/d3rXaLTW9c3feezf3MP/sl2VHcVYeFHATsDRlZBo3EC
mnsmNSN9B/6RtTPlo5AnjdnqGWyqMHqpXR5PPthPrbtioC9oEzuacJ4hFEa9D/1E
hyvNhg7i3bTYMiTso2ye/iMQNzEPCO2VjRJMCfdUb2XqvikgLb0weAJZN3rJBgMw
NrdDXBiDJ/EaopoXQXbStKXNnv2zAshIMeJmFSqoExq8ZtiRoqw08tpWINC0clS+
9AxpAS8/RzzlPyv7gwK72vHHg+9GuVZtrdgPGYaOewKnhu/x1DwEjMRh0xWIn0go
O6wTJyafp8MZ1ZKG/x+LjadDAkR9J3KI4iq8q6Uxg4AFn0+jVW7RSpVfjehvNJvz
37IvDPTfzSWcTGgZEMIEgwD+WAVHVbCGO4oTm5rAgYDQjL3Eq7FXgj7S1MBvIlEt
CVu3ZKExDa0OjMSUSVMiWPeA1q0sc5JVZmFzaTnvd5iHsDNQiTuHWKbg20hAyw1c
gmIR3gfBQXS3/eKPdZ8tPj3AR1lWLHboGvwcp8Xqi/dYIQ4g1VRzDArfyMZOrOk0
SoycUZg0Gkg6tXNeMT/2qMcDW+rvVOmh7TxdLQyjo1MWWMlxcSrLAWfHaoxP0VWo
IVDRSqdR+2VoEHnPBw644fg2fCE9msqSfxbY2xThkutwoW2CISI1v1R2ajbj9iF+
zAZ/M40KzNLV3NyqSJ4vOAD6wu2TvUbiU+U0/D/mWkeQFOMhuzYnq3Xl7VRYFN4F
Tpim4ZII2g5idHf6u7L0hog8qxrGsAWN/Pd6D1pxBcnYw9vD6e35UGwXWm/CFrTe
BeTG/fwPwKmAVV4lEn3libKYFToKDsjS+oJa9CFCZA7piFH8w9QXT70RyucSOhDe
cQJQcbMPH6UtWwwFbQ0jHO5h9cY+yQZNmfHqq8tkmYIGpKCG9KwJsAu6Ih2uLDUD
dciV61buXd/ZycylXDArwxiHjkZljF7UBgOvB/BLzQsz8omYyNqclYl5K/M+zT0W
EPq+yl89WyoAfSqt78HAbpUzZPYg+hl5wBT3hDKP9Swiace42kghHGE7Y5OAtwBn
VBvlY9A7g9QBi/bACnhhxbMY8fQRcTcWiu6Klqg0GeCX45XMg8W7RWcxVGFphCQr
6h8AZyk0gR3wDVw0dT3z/obO5Zvbek822/iTzvLmdv+4OBzdOYe4z0d1nCKS/wOH
7gHLc19y0B3HxtRHjb4ZmgI3xhU8xPUvN83EyBjtfq+/e8NbrmL6+2g9/gdTraYK
otFP7k750YahDt5TrNWxLJR77S1WfE5oleyipiAHWI2Tdt5VaV7jjN1ZL8cLuoxr
/VQp4J3DhpMtqPue7KgxtixMphgDqggx5sypB6v4s7u9XdQ4AoQ3vxoFFUXLGR/Z
Fs7TWnqHwnD3JlA2uVHQg0muOdrlOqqFYC0BE1RMyJIp2+vV5cb+WT2LcZAJLdBd
mIiBfSx+ovgagGlgSMqmHKxjVqNUx6jpQA5uW8jC5evhlvnvh9BBMWXS87MHotwc
icky8QYOT8rDTDzoLb2w/zOyEEi2sw9MiYyoXfC2eIhfQniCKe6IR8tSISwbsQKW
0r//6QsAyWWNJXcy9AX8F+UeX+ORZzc27OgiyP+X98pUSmKjGeUnTJDJvFCO6eBJ
F5x/e0LeyOhSXpw5JuQJ3mMKG15TsaLDt3z60j26iF5BFwpJo3xX21MU8NjY1dIQ
HBQKOijReN2osJgXs5kkiJHyvkhwNY5el7fRdTkbGKnr0ocXjDflALhJA6ayYKa5
r8MlcSuWMYkKt6VITesb58oR5AdPID8Txokk489Z8ULXms+t+DVFY7JQee+bYAWs
o3fOwIUiY2Y4G8tfoxvjv7vBV2L7+gjy7ggPjPAhKkgqeaGOtdfuYMFYvrUrXKPQ
hccqvZNYVZVy0IUVmvPqai455PGtsfZhScExgeCHioqbhOLeD05wjes0Xlmam3IC
pp2n89oo+hsqwX4fMVnUhNsyQN5pRp5XNTRjHg4G/f0cxOU3GT6OfKeTHjUAmXTA
O8yDadqHO5E7nD7IhAhGrMBAbiWXYTVhSKBS7eCN4wM8g1qiecewM89MIh5B2CPN
t7YM+IP3KiZ7m4HQ7wfXE3JuIWR06/l+xZT4hY20FfVeLR+uAEcukt0hYvDcM/av
Y3poXe3o26Zk076lNLV+Vh7L5p4lIXuC1Swbd9wJwp9m94pVg94KnBn3HInlzlMK
AK0Xeb3wL1iIFF83ZEs98XfzVKi8UM4FXtuGNjyM76QpZkEJ1cnmNs9RouH4C9Cl
bQZ0gFnMEkj0FGXcRO0x1/zcE9KYfb1+83tPWVNVg3ufajsgXTrlRRlpwoSttWgY
vXlWtudPNS00esZ820p8chNBxE0P/PJ1lDqJqAd5gEf2wtHyTj4N/Zv55GxRQXux
8c1fmHRG9dEW8ozO4fsHHOtqWcSQqV6LKn5G+08z30qsQbCmpmVA5dg4FjqHlxfp
4rt5TQwRd0HGE+9P8768XXTw9aB6EidGQXFcHw0lYQi4xiZgGkUOUfhyDz0D44uv
YzpKEJoFqaTJxdlaabBC2byS2TyPei33MytLcs/YDlyDoCuzVpqDplmPgWg9+cuF
dSu16On3LwkZskM24eAYxPV1ejxlLmTGyivVvJnuCNW9xY8Ipo7utGkfpxCQ4+QZ
K37AlXqWfOFeWJ5EHgdi+3/9Lao68sahf2QZ5GW4n6HsqDY4cSm6oIjsTXMzKQpF
L6YVqno6OHD7QFryM9tLvqZ4Kem3dXfhDf24oHtGW1BvMf4mRnKDwPumwl/fW5Zw
fwJcdk24GYk85btL4J2Vqt7NDBBkyC9FCF9ul6yY5nfHzWTJ6KJ5fUZzRMVuE71Q
IzN0ptbOsckos8OJqeRKOn8yAybTJ+2360PTgVpMJ3ysMXiovA4FWLr4CwjrfFjV
fKF3bTB96mthwpyiBqgpszzeGtqHEIitPlAt8f3xJCStk/NlZlOlY9ge47mfxSUN
+RUcoUHNkWS49IBekihv+Ax1ZV/9EJnRdPDwGnVJRa6FwDOOYoPvLOwV8bZNTz7Z
fdhA9a01nPETotXY3M1tMMyI5sfYhntXtv651S2lboUPf5asnip68/Ik/J963aAY
iGZnCLhwKSV6sKpa+/FiEZ5GE+WlGULT+l3XEokohqvkSCd+y+Ug0N/gAtYm849Q
KD719qqkveJkAYQ+TTTPkkJKXmzctMKaWWe+Z0RROCS6rkaDBymZh0w0c/qzYXrG
jFXCJFN8X58nHSSkqJh9NbcsTpc3Hb4zPov9t4nBR4R16WdGqzWig6kbfcBWYIdf
0eT+5FFr5PC57blQ9i1SOA3t01Im/17KWBhbwV44JkgIRh8tPpifrLuI6rAs3uXS
n90+gI+AWt2Dg101xhf0vHrjRGTfor/3b3Vo9kCSCfrAQHzJv3dkDIsJANKyzhCx
L+9/L4XObytLy5tyGSSHCV22wFUJxr/v3EHixfPphPC/YXEg2BlVvkCvQeA+51zq
mWzO4UW1FNbjyy6byBAgLUZZwp+ZApWyjQaI5xa6AHCC36524rcSMt+/DjjX5d+p
RTiV5klqiAe4yqnW2MdzQCWQ+TLbw3USFKzPXSAZFaf4k3yciqNzxSe+Ij0g2AUM
pJvAtUT4wwIoRWQyJgKxTKzYbWohhnFYZ6iWN2caYBoO0uBu64MO9Mijjg9yEfy/
hCXvIEl5BFk7DMqNlHGVCTihks2H9mbj9d49CJ9iliombQ8uajHjpdMT6b0gfLPl
l6V/VMSnYq2onMsK2vnt3WGOgcFMr869eNhQ/2oqSEfXbzRANisEs+jssF1xgs0m
vPccqTz3dDrbYE/+dzhgYYRQ1lAOHZxP9L9dopwSMoYFqlZTp7HDR/+XFIRV3a5z
atwRzl+NiaYctdXHHrmt4Mvd1kiUPbSn/sSkuSOYa9PGsP+sjCrPArbSgT058h15
txepDkuiTCdn5MGKJYaHkI3PCdm2XHRX5UBsQqqVA+LKU+KHw4PhO1tpqWnFhEFz
IMoKF4WpydSfC+QS+CuvIBxyFx8EeKiPc4BIEfn0d4gh1wyC9I0xS4nYKIJC+tmR
xu2SczNswDk/O8LPoeftxRl35iG6mMQyFwJmN/US881SvBXUYnrZEiTyT7MBczY1
Xv1tjPlpRMFWhsgZy+2pmxMVIVmroiQlfqjkEs/EZ59xNzlBjwjwYXeibgg7fN9N
ehybbYbUxTTsWro6TMZlc4jA33vN9VBALlW8a8/v34IIDDzdfSX0QHldxQC54br3
x7+VWIfaP8nPK+8Yz3UA54C9YQ6Dy5bUbQ9VKmAM+RRrZy6ewWjubyVmqPE3af0G
NrPFW90EZtlSRBLBeuhcdAOLCaLvDUCrk7mdrFeWvj91cfs9piiwqyjoJYTSQfJd
gpVxIfkP5GeNRaawnL4RhqZok4BUXdNbjjynAmJQWx3MWJOb3PlnTI2FIj2OjXoT
SaYaqzpCOC3Aib2Kdi/rzk3FxUTj9aZsqmkux3ug3kPyaM31DNMMlFRxISao5XBQ
LfLC0+hjmDki8+V8MUkzBX/vb6ZAXyG2Xc/tOfXUDwaQQmqxHWKXkoMK+wM+MIA6
pXMwgS0Km9Mcc3EttyHz41ySYyJstcT9dJ5QK6zuLDQKaqUcvaGvj1Xq0dhxLkG+
7rsjHXBxIj/B2RAu+H3iNXq5dBSm6F3xdCcHJbfMUyb0yTKFiozoZdgba3uLbzX6
VwtBRur8bUktqob+kqI09cb5eiG4L3/G/EPNArHmiB+st1302FHfRW2vZbFi5/lZ
PlKHNJkOhaJJmInl2/kjSY1cjq3zmrucJjKk/m4oHq7BGNeRpgyRnKEqbu6OAD+Y
kr2nyxg+uaJk41rd1XxNLTGlheLp8PVyVSKC1rtmKY479xrNAHvY2+kcvPhFXXj7
8RS4d8Dxz+bo8juKtuGu4eiwkluwqo77QQU+m2s6HnA4Dkw5E4TM8zyWNcaJjBYy
BJ1pMiS3U7PX2gIlsg7D/9cI7MiGVrOs/94ahW5nGDvTFL7VhJz3CfYpBBP3odKg
miqgUbgYODZxDspnBa+sEkX6WEPExvv0CTPdv/YCD+8Ipk8tVRDxWTtuz7op3WBJ
XfYuFLxzq0yvdh0JB+D1aMV/+/E28Y4Js6m+Hws4Nb5nTgZB6UJLweQn4QJdSbC0
WuhP1I98vvAEZtQO5I2FIVsbMkLhLn6j8/xq9gvpyEifwHfVoOghgpo/o8iwlO+c
vO9drY5cqnRDpuufI9QqqnSGPAZVvoy/PGrMqUrG3YESvcj+WgE8/J7z55v1s7Ov
YJVCrnRqxCnfBxUd/MyiIuAPfzD+DvXkSOpRvE1L5BDnB9akdEhpmrMQRPnCvBK3
MopafoKyxZpUtjM1Ght9aKUnKzvRxPbrW2WhArZJiEsqpd5wwEl97spNforJLgwr
mN8lucNUyjAoFbD3LqUSToSy/ld8n4bxXWPJY7dF/MG/qsiKMADG1HZ40mnoLQST
Q7T2EAoyTGXaO52JV2pY0OsWN3KXEe5MXWoa8989IpFk9fLxYjLMuj48ZZVPdWLW
g9U/xgEAxTqPY64BFAGpkj+XVjAJ/GO1c6pMpapU/Ae9ex5hlmxTt0X8AHi6K4zo
eO1TIycc8fFzaR6kRcyk8DIbDTypKu2bStBaujl01R6bVWIs1v5n6e18O5+7tHYq
28pKD6rmTz3i5d5Vtkm8sgokdbzfsUw0KgOOENks8TEu6nKq7RZeI5ocZZLmfKb3
gYcvDXL0Qpd/plIHPhDogA8URU6V7YmqKIpOIjZ6CepTQl188Li5/80M0ii+s2+l
lyCSFrix/x8BeSmeQ84TxfOnQwxvWcDQOoCl45y9LzbplRk6rf99USy/L5LWTtvS
nzpc+ffOPReDOlc19eTq5c5HlflYmHujC2MGfrcSvFGVBRKUBHA06uP3maoBJTXp
I94wO4z5Nmt3oxgoLe+eL6wg2dqieuTXJr0aZKBcrto7LmTv7u7Iyl3YCxvpPgSk
N58sleX5Fv9z0TjWdEMVQgawzhDi0YvB3JIFrExZKDfpq+2kNVjdMv2mvemhf+kE
BTa8QcRCq+2JmQe1zjoq0q1rZ+LfqDGzNwkjYirRpHIV00bFwqaRGTRdmUSnwKvC
hZvs27fWrgurEWpaBJMPBrtLQlTs9mD3rqLLCpARr0qwK2BT0SpKMf93dT86HI0D
kyUdSNrRSD+IPCszYVerieKWIVSRoVN8Jweaf7OEDN3qb6nn9uJz+1o6fkD+B5GP
3LdmY7gpag9oQtStLRjHEpXB4AfvdbdpgMJThPsSXX5TENlxX8fpqrrJJy3OenZx
cf38PyaXTe/IsxyYEz2KSX3jgDerNf9k8ApB5OmSOONFGuMx4HA5ocXlXFxfHqmN
ovuiyZqbtuu36+4i1jFdH0XLtw+BEwQiIS9mGvuK3WbmmRTo1CgYd7jqJorbD0SZ
mdJnw9k83BYIJWsmJeKX6colBj8z677XaKDeXKlgMxd6y1tANcTDiJTIuqh6rJFz
lrbdJbAyNFhYlmbVquzSMRlOCaO8pzTQuxGRuLaHqhKwMHBWPDj/Qi3UnNZ+KYgn
z/veUmqjglKlVLbbaHKb+gEhM2Ek2Prwb0UIcEFRDoqxW7LvuYpc9tKsAaU3+gzX
iPPoA7unOmTGwmLlUe20WvhlOYYZXIusdgVK50cRnbeWAFyBc/HvypL/ssZQ0uoM
fnpj8rqjXWC1Ca84Diy4kbTafLx3rmGbuuNqSQS9KXhlD7StHQcUen4U3blkF+hN
aVWupMgT28dxfgXvkmVUy2kLWzXlCl++CBLLY2NbiVVHRyC5yteXecgyPJW4AysI
0UHe5ySqyxCNFoLbjiZ9j8Kt/PgQfDZdA/QYCH8F74u7HhpiRaI8ZQ8HlZRr9Khr
EsrAjBo8UxFGN+/dcNbloiywYBgRZ8o50r6ewHOPbulY2ge0uBjLaH3ev5/FHHok
LyGO8VBowf8V1HUmdCYJXnRc0FTJv25yGTSyG1MjnQteFgRoohIXP3drtsk9VPh5
p9vsgoiGh4NukDjCUspp1yd6lQI7Uu1ZShQAMEOfKuq5bCmLh8qLfXilGmC3Snsi
PFcm5Rh+qDlyjH3PkjYx3aJOew83EZL+Urih3S+ULAP0VGjuItJH56+eWg0THJdW
ThYp49Huj6h4VSHmRhpuF8EDps65rYYMbK7hEGPNffv8dWSkUKtHisL2bsMVfmqv
ld7++LcLkqdV2e4jYQcXh47BuDDYOknZjDBBRoegYZr2IKHsG2s/XqaBWGHIctAs
V72tTNj4o7d6Ak/Axo4acQE8v9YDccYkzIdFjbA8zD8cQTF8yGb8AZ4tiGNpKLIk
6rDvQEATarNmSRo5+htbHVnDgT8DXsNhkPr6dooQXSgwN31TCvYCzQP/Z60a58uL
wfWB3PVZA0S4PgcEk7u6kwzaKtOCGEfp/NDTo0R/m8pa+Yp8zhHPoduTyw1fGLAn
8kq68NoUPEicfMbYpKLsUp4brmV664BD9UwREX7kgDwexlEqvQOpia0o8Mg6ajJq
y1Ij9LBT4OWsyS2SmAyF7iI5pMk6otp9qKW0d3vgNX9FjSZosP9g0VltRtr5GGgT
xxz8EBMijw59L1Zq79dtKbgRjWPqW6QGYAgnOPhcUXyIP+0RTTzOK6AuWcEUcuZt
AHa1QJy8fsIn0UAWIJsQYA==
`protect END_PROTECTED
