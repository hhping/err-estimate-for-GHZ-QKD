`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iVmJmgfvtup+cOxAPqO7rM81q7/Cv1Pmo5M91H+gBqy28h+sG42d4MhHISBGkXwN
r3yWIExU+MyaPJvgksPl6UPy9NdrTGsZOq7EPX+sRbuYAPQgBUelbsjwgrTmooV5
CIxkVWUdwEYKX+6UWvefNYfvRrp7f3ahXfTC6NTwJrPNdQHX/hmLBR+fgWbGo6Qk
u5LwJZL9HXE/YiuI/Dtm0vP5WlLR5PZFKFd0jjJYEh6lSeaw2WXk0ujXp0+Bhadf
bO7iXaRELHy806GuakExgpGkZAyAfmL/cYoGlddHIEvbQ23w6H/y7titb5bSGPg5
Sy7A05ec5Aw9QtKSoJBHLr/k6Yg2fa23Q3+jeZ28ucWQGeIcUAjB7K4HIxKu6YC5
l7FONGM9uwzJGduxUp+MbKVeMSIurJE8XGexzsaoeZ6Lt9NUou86248Io+llOPlc
rYDXvz8s7WE19PsA8Xea0I5/jP4Kj/OZd+VKtd2LcVRsRBuJH4eNNYeuOGuvgh0q
hOsdvVyzFc8wtuKSRJ1hGCdPJ7Z+H8OYQnh10Hxzor8UOg5kPK/k/hQOqCSf8pF/
BUKUW5kh757cZ07wpIlRxH+Z3QzEQSacceqcUnE+zoiel6YTTrCZozszrJYnW3q6
Fvn3CodY27qPViZl4l4fogMxkTZSI1cqG0Z5sn5PxpMgk0BDgcXR2ScrcE+gDVdN
b+qGzqk666GZJknITE8JMxO7GXyiHO8Tc2wDy/ex6qRIrezCgjfOVoBi8OGu82rM
T5LDebsrzoP8FePmTMyvOxsV8T9fvi8H6jfbFDPK+ACRDWOGaI9tM/IoygOuO/nl
21D+uIFZ92S2k60q+ObumwOxaz2KK75SLmM/UkOwO85v+2wJjl+tfqx+/MUUluIH
GK0imJP8t0aZtBSi2AW8Uu3Bp3/kXxspfjQkBkR8s0K1OSCGnbThpEVuPMb4YmI/
MXZcWxChKNc7GIQP90FrSxdZgcyb/eBL58T+be2m19cUefoea+RoNVbhAbyphzsR
tn0pOnR/OaRSWrq0uoUrlUTa0O2V9KjI66ErhToI/0FcWO2fhcTCVK+kkYPRUHW5
W3/IK3pfnjuUlScGMJSy9HGyV2TSlRv881YCp2q75hdLgGgm2jyx4MqtAfpwfMzz
g9bH/L1bCpFFeCFEAgM8nU3CfVWoJ8K9/18f7c6mkbYmUhS9+GwpwCEpQN6yu6pk
d5HW+7hQcM+MzKg1lemNDg==
`protect END_PROTECTED
