`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YprW8sNFCQ/0vm6fSUzlUOSS6DMqIY9aYg+Gx4dEMKtQdBJoDphbnJjaWB2JpROu
4Yrc2wUKysCJSGklE8ci1pd5/BFBNWrvO9ef0Bq+5Mw0eJe0acgwnsF9JcNHqvEM
sxO5kh4DnaeH/xvGyBAciTMCUPLG4Et+wYj8ye41G+cDGsIa53aC1081iBQcNWmC
JOyswyJczG/bk364+C5jDd/1bz0eC5Rpta+nqlTwNC4L3CSWqHXOUjzQieDC0WZy
XIc2SFO1DX10SoTN+iOBvqeEMQa/3N2AkebuawS4pxa2fi6sY2VHpNSPfILHwYv2
WuaI1n/x85IKciXDdLZBLfy38QxHWTTMdMme670itKxgP+myxC+Q2mkFTub0Pgkr
pSCsQbSy+MYuxKMboaFukERFKe8TYPy+/EYU/O1yA7WRkC0AIu7QGSOqptpXBqyh
U/LOK+ZFt5b/q4q2tO20cjWgcJ42yxjVBHc3FK26HGhEeqPk/Coo7sJHS3V7yHaC
xV7/+MmRrsL4zYPMfm4s07AS3MElu70WMtg2WhzDCWrPDfkeh6wbeLWbwDhIkYat
uO2Cvfe/ACtdTagaGoGlA/GzJz8rPKWeMORgLKF89OkXVR/fwFHJQrSAHFzMGEWP
4Sz1kSGrNYlzBXW5aEg8+89qo3X7pThbm7BKenryJTLSCj9xQBA3IxX3GiFu6Zbd
TPPg1B9pFAD6NEK/cOVVCYxApGsQl1RNXpKuvAlrzsD68zZwHfuHHNum/nPGvzpa
37lhtVWo+DNssb0sCGsUQeCNU2PJxEL8b0aYL5pY6HA2gwHhcwbuB/xbgWfOvEuA
EBuZ6J1O8col1HDbifB6Aw==
`protect END_PROTECTED
