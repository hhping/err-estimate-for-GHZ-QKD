`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVNOTUMhaAjfvi//ic9iSPEE1UsBvJVeYnCVRIXsfDLviTnw2eYWA23POkKGNW+8
lRxqTes0q4QP6LzxoanPS0PLfva8oLlRmQCZi5zONDnpVvjUHSr3vVhbgZJwK2Uw
138m6pE32fAGHWrv75u1+xFDWiiO5NLP8YlpY6ZP+BnuSLkg2FNxJIBT3UfAdyms
j0MBMO/k45YQs4fiyRj9Jhevlhr3yg2pk49hfuMkNWloT/xxKRuhys+RljFzBOzm
XyV2kzi7oIMQdLF52z5+wy2lQ902ZJSWpq+y75gM6Bh64ej5ZN2F+JZdXzw9/aN5
Z3+OXMFXjYF/OfQnYIOkOwqw+KEyT2aKPYaZztRLD+WiH3TYz2ebqQ7k7JOPAc2v
tuChlwp7uS0/B9i2PAyemVwwUv/fqKWi8lsGKyV1mXpS5K0iziN7rA2Xk3w7umbA
OhaqSWyYAeolmvaWqXLkpvOjSIRh5X5pSiUU3DhuOOip5uhGuLUqB1MYRV9VcfEn
tz2TyYRnrjVXUZkmw19j4mJbJyPUN3V0qcq9XyX709hHRgv9h1jNt0gBw4B1dDZs
UoLaJ4V5EuT+GNmINWW6r7QWDOu80E2yrI5GkQI9MfYtgb/7hSdMXDs+DuD7D0k6
qpFxaWWs/bMukzS8hKPZ/gkUaGA639MAx+gvP1Tiyf44WFuyq+sOjTSsxmAARLur
SS4NRgZWvGfXkcP1sV6LeqbRxeWc9U3rHGFEXVNC4UnIkZWN9annz+b90xfDN5b3
8FFzJ67pTX/OEFuLYVnpIVvZcr0XJPJRAiGxhcFt0HM=
`protect END_PROTECTED
