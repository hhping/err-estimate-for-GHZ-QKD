`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neENd3SoLTMMW1xOYlmkdbUK5a64iXYyz8OU3fEUuqvVGBARqp/0Izvgi2+oKyWE
zPylW3eCqAhQs8wtAStYfy2UhgAdN9ICHhtfO865/GJunoigdzvJmrV2Xguc69C/
XO40U3YgThc35nlcWem352uP6kFXN8cAZWfPaQONJp/i7h8uREeVjZkgp78se6gZ
JcQwkbtNq9p5DfVC2UjQLYms51tAWK3SYHiqOvAO9zBtArMHY0YG9OoDaHMSfUeW
gjtqliaSGW/H+OZQleMlJ62GwmXQ+cqAb87VJCAxAf7qRj3YNAwQVCiDcQEKC3xQ
o0mGKDB53OTUVosqNafIx48j/Jwu5MPIkFZe6s0whBJ+taId2nZGmXs+67IN3vNU
Ga1Cs3TCGO9IXdCGAFNx+JocDUxVyw5Bcq+YRIny2MndJp6feFOQryoUqatNf+9I
SbAgpO039o3/PUNYh5NKnv/OzcHmiqDzsAPPmo2nEBjMDhLzE+usOWKnb8IKNQUz
MMXps/ZcDv2yJj3aqb0Ybd1H78VzIGk/Tts1AMYYy/mH1gbJ4YHMDxAYVpO+k3CW
cH0ai1IdjYl0NOnFiLE1fLDESDy3731EV/29eKoZxVzxD0J9RupHi+oWlmqBTIvr
UwoiUqduDsSfbiRPAA1iRxHuXSiQsIqXrb91O7e548yKC1exxCsgfN0ByrNzrx2K
v7MRRQat98ucC+An7Gc8GJz36/Iw3a6b/YQMXiLLsFzP3mK1vIdESmoyT/P1jwZX
HPNsGC0R3vwCtTyg5xcl83U+Airmle1MuSdW5E57BUloVRUf2+xAp7vhl45GY0jM
kSlHypZV55/BdSvKR0f6ClEXxzzrn/fUVPaCWOUMvzE3jI0qlgVqMQzbjV1/XyM2
mOnfKNrpgzkSaKZmgEYEr1CXdje3xK/QPM/sCS8iQypmqdcLsfLICOeJgRqpr/Ij
zhizNym/IK2oSbJMW/r5+7QiGIVjbtB1PhJISaahrY4Bldfu/11xTajUbMTXRUog
IHa9JAk37h95zDwgq0Pp1AZGhm3yQGowl7NLHY4O2ufaOq3nLJgGWRHLFTjHZMU/
iMDc3DpgRfX7mRIcXDzcXo0dKGeM03ZCx0kiQ1va8qL0M1sOkoq9GmB/RvBpOvNg
n5uiNwpt3RUZ5laJ5uhvWysMhAlGUEFRhVAxVvENBqEaGRDqYanN+CZ9+0Z2+hfI
soPv4yayocnikROA404e0w5T9slIbsMov1sYIafzN63sW0KitFGgFFHfU+oxECV9
S0UUUOZ3NBcmUeBqkEZoZ0E2Nn95gQvB/69pXFQmO0J4U1HfoJc7OiDyre61UwlL
AEotviNa4NHB9Zu6tf5Yz4d0IzqtJl3AWwL5cjkJMusl2Cs/3Cc5jXBcZxVm902g
3OMbBa/bzTEMlxAa/OAWEp6W6iyAzeoJoBOssL+gX/4c8kJJ1sp2tNWlzBlMWvKT
dBRn8+uH+Ym0/w/A8HXNz2YalxOOJ+BbUQZ48I7Zf+JiITcvSAiU41rs4Qftk4hX
ScFsQpI35c3RtmUg3jH/T4rUNklczSLWc2OV9EY4JGc35J5KTOhkov3s5Dbx5AIF
Neo8mM2OKVvUgtwpmDcAl9ssda03X7b9NVxKXHpIqfhYRrnGXfmrnRNOsP7K2xom
k7/Tl5FKV+sJMLVk4KTUNJwXdDzEs9R6lPnavH5uyL6+5STmqUhDo/vSmUmB6cJc
4qg9gfG8ShGOfXWrPKG9F33SLlBtOAdrA3nh+m+B8DNhvmnSxEpu9KqzCHwHjzMs
SZpGDVXblQmjq2v14d2srFBxckwHWobOLlF4+F1OKsl7+qrUBp2ULl53+IiYz8+9
c/GmyQAKhnNbzjhhM+0wTdHiw6vaiz3i2ncTNRipG6DSkbOkH/AIRW2CfqQUZsGR
USVpX1ElhfA9V2upOi6e3gqWt6RAOMg7o77H5UXuqvEhP13v7STI0ZBY/kNaWlCN
EP8vNTra3FsB/v6ZkT+K7WU6CB0rWhvw/ag5SIiWDxG0meSZfPhIsK5zsKcvHJxn
szFS2tNSO6RZYYBJLAEd8ASUxhXbvqVyaeRSnrzy0yRcZIrOhcQLooGQSliikFdE
YID2CkhPIAUZYOlR4tcvCnT8tW4QlavrIXfkhIsyAxFuVgOgqfntDx6F9fm340ZX
Ex3Xi5QYTTmnQcbOtiJNWMCCZB1PWzPNDTWfAqkluEPh6EIcm72BUrG3xp6RjDOg
qcko4gxDGVMuPK0uATVaUqfr2wfthRaewgyqDFsH7wuIWZhVuGU5SBzvH8dqbfTF
RwAyqWjKO+szLLMgYL63px0niZ4v+3jbuYlbfbSZkK4ws6fvy6pYNVvBWMhpHBoh
Gd1vsHIEse4sv0ORlzdAb9w/9zxSbAFN+G4f55iNM5DTrWwWQf/x2AQJ7GcJmViU
awZnlW4/ShbSnSZ/xkxy+POcFC9WgUZXX7NQDuoyDoEt6KZFV6KGlZ/j4/Yjes8n
slYaSXc9aiNxXb0ivsEAPCnzcjSjzSPxMG0H+Qt54P2JFSGJUlsIOouZ9k2YqDCY
Hno+3+e75cpkXGBix8s+erIExMHiGGw5947mw91zsFZEHf9DUT8QLFJd3IOU3PUN
TW0AYa707qyxAldgOIRnEgRzX9/LJjyp+dNdjMwOnnKuhbLH0wBb7VCO4+Lmp9WL
epQ6NH7KygmMod6CoR/Hg867W09PHARNJeszjry77PkKvcFZEemabbGftPg+KPgv
kaQTysklPu/Y59ZTmt6fOQeOGHrLlklc50NeRuqOVH+/nElmFDdR2QiiDLI6s3/J
9LKzqmgRmtqEpXZWJph7kLpuQMk1RYDrh9kzLGGsCAdLeJOnQWRzNc6W1NlOLW6o
JrH2HskJrtl8FLkSfUPcL+Nju8BMfc2LNGLVi9Jb/nPnjAOK9pc7bqpSHV28YAlm
fod9HOm8XLolhMwPhBBbndSckm+w/PVzHzxMQHaPMhoQtRUsGRz/ZPwGXMIjlYcV
5+IdGFzxiNuVSVe+/7lJ9VyJfhlThhFAa9quopk1IoINowUWFM4/40XQ8BMHHsEi
99kBc9FtQfRoDZEv6H+iHxXrsFJyQWw1UrA2GNYSOSvxSf7qY86A8lnaJZHwd7KC
vAeNqj6rdRMFgz9EhOfQJoBOQflTeT3opccRf5wsMLxvyu8rnZsJlMQTB0W2ni8K
FZcDUgkHrLZmgrUaqAod0+R7UyIxr29VbJGb3Tq2zZMVZpO83gj19jngi3gLhwxu
QWilWh/KKpMzJTJK5TcXSqhbKizMtJ9O7lqTpvx0xTQW8CuJOCWBLVNdEJOxuk2J
kzCfygkxkzmP9moxUQD3GB2nXcg5OkwwGqdP3IQCUOZsdpN9I4p2Gx3o4Sn2+C5d
bP0zSQiMAAusCmwtBxxT0oYCQZNtUFdAe1RK7cUFDiZN+x4vjRKkdn0Qk9lYKjVq
r364M7AkgeERRAPljlSzLTLooTWmNxFOiYDTNFpFZdZNzt7OvOqRJ12tiS2i7gEm
ux+mEJMvnnB0iIXpdRk0GfBNf3kivHbt5Sv3PMwCXdZBF8PWG+m2b+u0H7M4ZATe
FOO2A+BoM5sNQldGhxKaBz3CdK5CBzqdPev+L3XE0TcbnSTKWsJAFjPWTEPd6yc3
m5LoiK1pPQML8dtKJN5nAPw+QPatq24vlKiDn2lGYHn9bhA1q3f7HmIj0LvYCrkP
OydxH4hHdGP3j3R1PBSG7yPOZc49fxNOhXevLZnT+G4W9J3fJY+N2eY1UFM6Iu8c
zQek/zgOp/2g44Vqr+YoDg22Ky/AfQFUOBPrCh4SBrtZ8kwQjr+/nK5cf0L0hGLD
a1zD59xPC+JY/3hlvVg3VnOgdF7R+p6p1UEk/u+iePt9eowjvi8ekuCacNdEJdWc
l8aCUR8XDPBsehzj4574x7/xW5hqwvBsHNzmgC670jUUA4b07k24puCigW7ghXaA
0Su1h8g2v1cvE+d5KJ7BXrA61/wrfWIlkMDeqCU6T4/iG2Nwq42wI4ecxadKIwea
4WJMy72wARUT4sO6JilJECAM56/UJftXJwKEm5M/IBZDIU7HMHfzh0oheDC0wNOI
AuKzrgF+rA0zeELg1sjsEamCXjyVKA+lWj70ujhlrc87s4THVqo1pasfmuBTgPRb
eE0xvMyEK3Q4gKXrrZ1EdYE+johLydm9uXY5FLHaWdg6h4quHIXKpa42+S7YERwF
wqoi9HE74GXXdAljfrEt39bauu+f58Hh0TB/kqohEvgKzpVye80Q2tREYnN66aLQ
5hCj5JQxJLft36M+5HukR7gd+ZxL6CJmIwyhqieEtE9HRe5IN3RMi0c9bPg+GacU
`protect END_PROTECTED
