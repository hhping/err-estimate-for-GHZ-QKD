`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0PRdz8gor2ZKWkJH+8ho162cw6+u72hERGDD0YcqB1yJbhsX06LIRUXL6eYZHB2a
r96O4GY5ti7wPk1mImljpaqKUQfcQqqlS52PZLR9xmRPOGEBLTsq7YMV7L4pcWck
k/gouG6Ab0pf54p1JkBii886NXvR6udqmhuX9PWymfwXL0vuBtrAR6KvUBr4iAHz
MXQuSS5yWs6I1Y2g2PjCu+O7rcCTE603YlMmRtXet6URCOMm58c2ntK7IpoIKkZ7
zzo1/oCZ2N5kPcTIiLu3iC7fN/3e6aSW5wVV/2U4Ckttsw++KJu+hnGvdXDxY1tQ
37BgCBGV5n1dKqQviJyGBBwYB+JPfcMj2lr40s+Ne5otGImxxIKCLqMHcbKy7dRh
WxcRPxfeM0+Ia9720LOJ/+g20xBC8Mdvk7wMHny/rss4kQO86R07RdBiNvKvzpR6
VbqHG/MY9+9oULrK/fFLKFLWfqz56EVkc/KvF5HV5pZRdez+zB+nOKxpu7xaC07X
RZybyYFtJ2+agvy2cTQv0+c1C9YJRw/SmpD36qI9IlyvDVlLrG3oHrPrXE/uKmBL
JypHmbV8T3In5xU0R5lsDpWHirhc7clV2yg6m15yuWOtD5BbwaLTvmJirWjQRKUd
3F80ti/ALQcFHSn/1ouRF572WrE1gOssE0zMQ7Kc2k23Ff1iQc4NMRfzqGxJk9DG
gu6EM4TJIvxTrU45/jtABN0bPBzkQF4HHzMYyu/TTa/YZA0AUDT9PiaNJmUiYX/f
i27Sc5Z/UWFF8OsUV0kHMgdfr1uHhSa91fqYb9/f0VQ8wGvDlkW2m5un8Hbe8HUa
4Im28S2GfjrDDAgIEaWtFIrFCbvIp+dfN6sVJs/c4ih7k44dCVsx2riCOvxZjfOU
U7eWR5UslS8D1NypwyALUmTtYUV+C6mpdgyraQdbH0dhoaHOSH2XRvngznmzikl5
x9QIv2zenacGtfQDgurWbQ18dqlZ28JzybPl0IPfclFD7ruhgA/lTSlFTqccMq/K
E1bOLt/S7Z8y3ItN9CwB3ABfo1DWp8egBe0iS5GR1KE/UdJ2K06ssE8oHMa3IPbg
6ES6NucfQals3OLjiwrZoLtHc70fTpahXGM18hVLn6jeEZjK7dkt37gVS71sGofx
2YwfI5T4CLVVd4fidsp9AQXEzrF19/3K7SnQNS1liV4=
`protect END_PROTECTED
