`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sksxvEsW59ZvygqnC8JNmEAxv1QzsVZbzctUesey9enQaZeZ6ra45YPm5TMgQrH2
D+CmewaPySt4lFuJToWCh/5O66oh4IO9yBrXNA1NP6SLmQA4xq1VUsMKkgqZl+94
AEZDCxOIGJrywONzcwgldnv0gX3FTVYswhXYi5rhqcaeLJ9oGdUVChQx3qX5tXHb
zJokuE070WQxlh3IssEOjzfZw1YaqB7jks5wGL5ri15tKHf3Sv8e8+XoOn2wiyL9
5EnC8Bc2nznkrARsDfi0L95ssZpPOmRrmmztP86NRdFrYKfvf609PptlDQmAj8JW
e0s+RLoqZj50vWk6zZik14sVNY9Chq/i7Kxur/MQ/YGHi3Grc3z1s3Pp/NxKwoQz
8x03j8bznG7fNi+WT2cuPeDWi3UqqetUZddAQfnB3l3kDu4BCIMQTfzNRp4TZ7hD
5aU5tRhBsddIFno26VNXO2sUAnpJiBdJa9z8No5vcmRleP1C1SW0yebVr5O6I0Wb
tqkdiPpjKy+wy9OmO8vvGge4VCurAWYrFAi7soLQxYhinCCImldK6TDjNCTiWx9b
96LlriNOwsD0/nEBkGc6stGzSXszHMMpVKFpSa/bmDbh/mQwvF/AEgwvjUH3earh
QxyzOI5p+oaE/1kb9Arddw==
`protect END_PROTECTED
