`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kT2VNQux6eY0BsFzeYgbIf8dazePdOGF89e20Zd+KcgJ814d0uTJ3gYCawwcdUI5
r5HsjNoA3SQrw+YNlLpm9vRP7NTxfB6IzYVvNabsNMzpQB9lx/p1jQaktOO7PVxt
T0xxJTeD3755m+lW3gAEaBN4pQcNVj3PWaNpinGZsFkGPqGlAKD91FSAG3LdDR+q
N/8vUB9b5GZ8Tv6YrmFQBaihNkdIY+SXEmrIClhXAEstjhVuwuRIi0sOXHcDizCJ
zmoe2KDgVjE6NNs1IcxAnohaWuuNaQuqv2uEbMuyWJBVWj66NMKpAyaUS4Y2Mdc5
48Jmx1CK3jkOuyQ5CKrZziJel+8RYs5xidsWcTitPYE5EReQm7eiRbt2eR6QscZW
LlcmLQaczCvEFJ+o4KSnFmJvE7gHt7MloOaAEzuYWBf6Pi5XpK96WqL5EUHu1kH2
2acF4wRRfMIWa1/mKZHkZPMfj/QYmaF5vNdZcVkWp+AMBPp3UKnmGy1YEJt633OF
022PmDjiHePbikRCuA0TEyn9bVjqWAdaeu0xJ9CHsqzAMUooQwQRrFTsdC6Cw2uO
c46Bq3l2qq8pZcekxsy2wg==
`protect END_PROTECTED
