`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3szCJ60z1AUAIkmgX9pZ/mjliZSp92lBzAFQr7anPvnLUogbN81crV5J57jYXPey
4X6tiMqRyVjIjIdtn/JbSCAyYctmXlimopVtc9zarNdlsRBW7deGgGPj7+JnKwmj
U6aPMcoJPV5+nMx0VUjMerVebehguM69lWdZ1NkqkAxTThxSe40CNYm0uYQWOcVA
WcY0FLw4wuf1xxbx3KQdVS+qDM++Zu1dpVRr31AdKzwWO15qsjVEjBUbpASCAFh8
5LkNKwzrn7XapdHQgVP4/aURqgTCnvka6NTXV5Cbs8SYjZHSU1sosp3nRTcq6+VF
ohYoBFx1GoPW8qmlsYlX1zXevd7vbHYnK/z6XStSmOhw6oa5w/n7n/4fl7m2hhuN
`protect END_PROTECTED
