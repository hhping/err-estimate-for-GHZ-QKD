`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ChCHt5bjjbC9RYiGWpg6DgouYVPayVl7gORkHJWdsffjMIOWAbSr1UILpEwMlRZY
iIuhJKKZwt4LnPMkC/KkJMdJbGXM3aSCHE0wETk/Qd6JfVLCRw9+GkxSRCFqPMOK
FUzqma77yWWZ/WoXgPB2itD96n8eCDOvZDeftStcLxdP5tTprLH1A8m8EU1ylIuc
KSgIDGNwSdur2FTlDxrD1Vld6x9OQi7jXFRzIfCJFjdFq4T76NBIwqdO81C65J/I
sdkTY2dxEM2AaQS+MQCg/ZD3qbFvc2q+ECy4vUxw+3NHOJxCIlX3Xlt/Bs6VIIAu
l52Y4aGUOavBEPRk1kCoCPIU/+kwq3sArLg94sCyz5uCS/zoKIOfYpyuvwN6pvzt
mg7JSBvvfHsgZCt24JcnOyh4Q9CZueqdBJp3hHP8hEMKj6bAEAOLi924/vaqUtrX
r7efC5niM1qCbPjz0wLBOdMN6ECF4wgUjYu/v5iTFa2W1qgoY1CZyPPTDzECO2xO
Ig40PkYe3rXG0bUFcndIj7oaqy8wXCwKhqg2kJmkV4078rVWka5hR4nZ65znBPLl
HO2Q6VGLSa2vZnspKLUqiU9UnPRY4dSx1qj/2OScsU5bOQQvEuGesaPKM3XH7LSb
ZLMj0/WCI5JtMYZxan/oDRSqG4vtWPLBgaJ40CORHZZ0db/MJXqo4GFl9S8i7ut3
FHmvUT54D3qiEF58RWwZZTmyjuiu7I9QNwEKHtvxs0eS2C9v+/qkSkkWv7wqYnrQ
kS2zmiyKS+sufgxYJFheNxTY/nGtgBoVIiT/yYitJqwRnYSdcTJpRouNeaIVn6l6
0AW+Ig7bPm9jQRa0Y5UPl3i0TUnZqpvnRYr4UW5yeFiljTpasGMFi2M7pLRgS8rI
OvMQGzjBKW3XCFIk/k4saVvpEO40nKtrtxSW8JLGJE0gEOErtNlTL75dUGO1JWPm
xzZmeXDIPi8rOZhvxO3JozSV1dBzX9PCqBNFXEHzP7Ezf1PQespCTUEoDRs0J3hi
UqqXC0QJCtUEOp4Dl4ygtnNpe/CRMAOChgjNFER5x2jWNMuR0eFxp9Sj5O4u2351
m+V+yHnK07Vzo+8Ct3Q9yTHEOjk2vAxGgmrGW8FY/37aKz72QwK6fDCZMMCaVO9z
8LoHRsCMVm2Gp+jyH+4U7XBOXhWRxGfUlRhLIbx6pH2JP44hSO/4Vnthcl6S5Bja
whSdLsAYpvWtG1mPDjOL7o38GQb4j2b59dRY1/DhjfdItwkO23mzId+vDyKGRvdN
+4FbeH/I++GvX0Fxiw6r7nWQtDQ/g7djLxEogmqrZTaeiwN43U4XZ+742x70OUyg
zbl6kchAP+K1tYIRyNW8E3gzl52Wce2zKcQHCVRs3OE+qFrNljAESm7gewPGOSxO
0+lel0RUQqcANXAAL2zgcQJ4NP04oh2rXujDVF24L1uf+2WVym+mMN2/VMtcL0RX
NXoFMZzfKJN0jQOXtT+ishNe8UuPf+UqH98NhNsjKDqRULdd/nxyRETBoaaOhg7N
I6e7+XNMN+bOYZ87lgflbjPmb8iYaytLkOLYM3v5Pr6HUqXCayae7pforSxNmgrx
cZAJdFWwmhW9teYiBNAd14S9QZxwTQCCUx3f8kSELuk9EaDPLcMz3f4HLMpmJ1ON
dJlUUzUO/G11o8OLuORmEmXbyWOxj0m/bfi2AbJQtuLdq2xN4+KF1XATu4RmTLYp
1ru1oNAvypmzhnd752s90wnOX6VJNptU0QbD3mdS5NTgfJfxqrafbdZe11t9j5GZ
3jalCF10J4ETJM8SSmYe9nQ++aiBXraSq+PdmOceWF3DVZdyetGqpHB3govuKkVq
IEKXnDmdY0j/nyTLSMcr57NvgM88cMc/YD2UaOUzvZ26DoznC77E7gdNB1t3M9c0
U2UwvLeWw5xu5gO0gQz8GAv+y6G43fulpPcxUmYni3PscItbE5mgadWk37DD0JfP
qNy6EfWYR/rtBTaJrDy4e+Z3dTcV3/DTMeyqb83+gwbEfQ0b/1J7Y5M10YVlKkeX
TrPNzrmDr13k9LsHfZkx5XyO6d7HGzULd51V5ESJ7L/8NX+ivAlADRIv5rU3A9kl
P909Aqv82rRsZGIP7xhnQ09Hrl2tofHZa9lgeJtgV80k2HcWmyHWvpL6YRiChKIy
c2hSZ6BgQq/DnCnPFD724C/Lj9TvSByQrQeasZX7HNioE3mjk7E9deN5qjxTWJcv
y9kqjtOfepia0ZaKCUUuborkYWkBgGMzumWLn+X0Fjx8Wmqm6eecwxBM1PuDqhVt
PKOKZj4vAVGlt1OrbQ4oYbUSgN97DFJ0uvJmpt3PhXHtFhxBXKe+Hq4eEMP4ehrK
sloigDbSYcH50/lH1CLSZ9sKjW9Gz2+bA0n0Jtz/ZLqqZbmNfgQFMESp9fI0HuBh
Zn/1NOglc54CUgLIYF9SB5BWistBM9g12bPD/zyrS+WkuCBHEwwdHpXiCcFuxdEW
QIHrinm9jmg5toegRilC2ETQfI+35pnBU6cwXCDUHcZx0xJnD/oPdVJGVuumZ+yN
HIZh/4KmfxF3QhxQpffqwjcSQDMH4DsL692iFrYncqwG9LN/J7EzNTsKM/q1EFsG
ge1qbpF3bWotBBETQWMafZ2I4vzrMJCM5A7an8uH/IYQcth4bFecVGPPSSmhAaGv
LpS7ukZZGaOCYSxj3MfQxBn4VbYXOfDHWVNehV77Cv7E84/6nDpl+q9aY4hSNhTV
S6XVNKwFaGSaJJHjxR9Js/X0QAcyp74JHIbiv9Y2UGml0NfJNhX48zMTkwizBnSE
cv9CE2G2KrPo+N845ALkdSCPoBn0rARMOnyXRh8dI8i/ygo5BzoY/uof5Lhq8M9K
X2nbeZ1hwI9WOKbVvz/NSlZhRnTF13hbwH2PbqMFKLVCvI/f2nLzgWOTyZJ+c3Nz
9YYrq04AdFWF3Es1bBNjcm0DwwlG+MHSobpfOrpj7YlnvNvd2ml/yyB6r8EK+gDR
+RQdoeVpr9upyS/ZpHSfcXMyFIvY4M9Qk5Hg135fMzdAYSQqqlSLYslbOQak+mpk
8qZys3tyU+GRvff0KlYTAop+5Hv6MJobC5d4MeY6QsTjFUjdDGTCZDAPx5p44bp2
BpLEzhM/j79dZmZAOsCLz1d8v9hb9J2nW+4TURw4YeSTf+18ftGXtCTn6wN5mxHP
PdYAj0rPjWfQjrQ+NWEJ5OIVEwJGzcJWcb7tGxEMxOFEnYpTUs7bE4YQCSFP/x5L
9gKoC2CKurpmniuMho573LwiaFFXryMLHSsUyXQkx2Tvk1PM/NCmuFYwm8uVxFta
FCI11pOYH7rRf2MjtDXEUJWl7SdcMVuPGpEi7pX1SOFYIUnDDUaG60CKoPoLL+IK
1d+iuS9fTnluE6qJbwt+qKc4zHmGBbLXKaWprId/38nqEmwNr2oVSXZWkpCsusEJ
dBulZKx6rnXdKoEp88g/pPIUo7I544MeoXhyCG4InbHfTB6bNIhFpiY13dMlkJhK
a+Kfhu9PiY3Vde81as74CBTzUTkugmHdJQtPFKsPleAY8mIIwCYkxXzpHhfRR180
WrtjlbTJP/sRzTxSXn3AsM8RLb82VAdnmc9D8tU4O6plJbrlxfXdm0x0Kg4Bg/UY
EXfzv1jQpuQBb7H24V5Rc5aD+LB6tX8AD4s+HnXNvNMkDb0+YgHW9rWqi28Z7T0+
6/M5hAh+EZj83EwfzogRml42lqFu526xHGd0FRYIRa6JTfcyZT3hcuiabRqCtngA
Bc22/3+akB9tAHow8MWL83gNebjdO+P4ps/gar/2rnaN7mPqhOKU2Tin/75D0XH3
O5E4qZaoZbYhxsdNdfdfhe5EBHgkV2hk7aN8h04qppH6+w/GQpKJJlF+n7SOSAb6
c7McDNZucBuSJ+R9gfr0HzqWPIlfdYA4QyZf2YdE8GElBqt0K2kF8zWcjmVWqnGe
CHqLYuvBG7IyDaBoqvigTXq7LqUwQCTd1zitsbqimNc59/7kS5hTvZ40GStp4ZsI
iubMxMYZuNaynDJ+IxfxZjM4ynh83odcDDSayXqOVrWF0lRDKT3kbr1Rh8yMB4oR
u4+Jzqh9E4Ah/1BSi3jmMbooxmXRxPIHIeMeOPDb7O3jktM05YSqt/yqGK9UK4Vd
XUpFpPZksQZmL7f/y5seh3UGoi0OxAqa9AMygLUCL3m6FF0sboG+uDxuYN1kMTn3
hubYGEoZAmFE0o7qqygYT8bhpAvL8EcPUmrGkwPC9jT0YbNBJNm55E8YlPUwDfAK
Ltt3nPe4TaplCFqflTMcjJTwQdactEH3AIXPimTDtr59BlGtglf8hHOAkOO+3iBH
wfAFtxXB/0cYcVGaOSaHStHw9cuimLTaAfLgsy/OYfqrGZH3xOiu5XKRdF5SnW1E
rxR7YG5L9iweCllpM6cjaNWhEbula9ppkVxzZdLTLy/6K/nc1BXvDsfmqzO6KECu
RBoaJks8EcwNoiNRsSLJUbnBM7A4RFxnH1hojK8Io0bi2o5OTSysUeNJ+g4U1I81
6GcNa2Xhi0giju9V8BCUo/kYwbsFEPu1xlNw4xsDDHuu6cuP1XI3n+IXJQIG/KEB
Nf6dJuwI367yIVYK9xA8AQ2nXzet2NspZ9YsFGKR0z9W/YT9Xk/U2xt9ebRHZKQF
ZCd+/czV9/DOKpAvoZjWHWqSUOAcYwwJWLXI6oCYqUYOrufeEDDdJdiTdG/DF4xP
PpuFGbm8swo2nkPeS98WOtaWG3j4dqbgHqUno6mJzDqM3ODJVBEkawT5HfrOx6GE
XQ+IS3wC1dHRYrpC27B1FRV43BG4N0yX4+ug7sPOi+t6lIDpR7k85mtP+bVxc6BG
o1uxVcEy9MbnEr7rOKek8pMKjDN80q+u8ghZwuHrV+1Mfxh1oOl37An9JkpaHWoB
5DcHqOpKbHavseA0eR8H1pN/wemmf0ZThi+EEUGFWLE1i6qRh/kUugv7BbmRFLjH
aXqrK+BZoaA8pzpQf+GhKdXptkfng7v5MsfGg4tjplzLc9OHVy2u10Y13c00YeOv
MUOaIxsG76QGKyRl34LGT/G8idcKUuBAoBAc0yWJlPf0GHoUQ3656KfICJd10FCo
4P3q7rZbz25o5ePMxd6oJtaF7hibYrybXURTly5H2YASVVD4kqME12QNLl1jvjNi
uR5gbPtpmX0ML5OQ5eVIpe7T6Ql+UbWckY4fzFwUjFjOevAu8qYVZdq5f0721AvN
Ed1qGA0a3hQPxAYLM4AelwB1LHAt2XmfmmvmSvQ7ef/sUsfC0Mw+w2nil4G8QeQ8
Zi5slzcqpYhQM6FmiE3oBvCS4BmcdhctC7tvuyKPOn1TUa3DzCt/OL6iKMPws9sC
NCsVtEZk1RJ644Sb+cdbCzm0iIew5Jr1JwjwpfgXSwG9oDIOP8/BoFte859aSsuq
3/4q7JFBJX4GpdDMMehHtmQGUHb+ci7MhZRMRVg3ZXpQB/vg8EkyiKGeNIJI2DBt
yljOkx0LLHGMQve2b3gDDIlMr3JS1ghO94Nqfn6WAllQsR0uKHm4UJwdK4umPPD8
i/wHuaRNaxigNDv85BMS7Ah8izj1JKYJuHpDOVca3tM1C9wlysDRyRbeVHMPNMaa
TJMnvdc45+plnOJxBmZDgUzDtZkWGlANpkyC/dNVozOW6yc3CGoBaA7qkO7ECOOM
nTZerRbL+HxBpRd7f3rUOu13umDIeHUe5GB0AyX95SegJQVzvQHdD2rZtXqH458G
kuF/yX+2fxelAaSpkGGs5pVpGYmbsUOt4Jr5shd2s3khBO91d6PD/tMz58ZOqWoL
FnQ1tDucfF2tEXYuVlDaZN+4VBrdB0K+SMyjLlfSjNcmLfNxbS2XqYOy3dcITDVq
QnSnemQTYsEuuRdzK6jr9apHdobsikwWXVJmQA4q37kpGK9oZC1/r5Hps92T5rRH
5ATUfZTxwDNQksh/STAxBHpFHx2DlvebHxAC9ZZnB5eGTr//NMk2llufq+h4tTNX
Ix9+V5/+RyC6AdFRL67qlFnCueJL/+8TViycf1QQAhKGqStEMEEHI6PVmHBwHkRe
A9xPcAWy02580bQNRTFKvd43xCX7GCro50EDEawhSOtjZY+ASYV7ij4fvbz7jpHp
0h6Fu+jcglbgiFEXyZrJazRxAEO0ZzN6LbNEIIWoyrHOr9wEHvWcZ5+5dQsskSFZ
aQ96piRbSuqlaid07rUIGeBG6XEi5xB/WqHO5s6pNDzLemGhsV+plnGM5Bpoga99
3lc+yrh0WpRaWMTlAjb4ZYCvFS51FCBcKMh+4E6psDppmsMdvFV2xLeK1anlvYzP
T5m+W1NXN+F5a0BJ8eWWfOtbiAV07mTdPv0GQ0ANGI655VGnqqP3dRNOCc40WsNw
Ev5CMw8Q1wrHEWQsSIIVyOz8CbieWZ+OSehlrnfw84SJUTSpiU0mKpJVohHvTT+r
YWoqtu0fS6j9pdoDhsu5OHDbW18lEIgWmPgJO0Dy9+vSHCLayqRzvMQ63oTxGbH4
5FDg0NKqyjkvUd3XD2fsw+83Bf9vh2JLdfv5duwzs6O0g+vy1Gm0nNs41KD4MiLr
F3GpDeMdKLh9TbxApahMkzrFRxPo/G3vhS+6GlVYYiJVxT2WSF3cPXXvBUqJTkmh
avYx1oibE8r8aH2J/04cuoD7mCYG+8eyMzhZunZJbUnovCCuCn/yF29efBQ0Kx5+
kjG/NOxs93n5v4aKkJYzxQYEgA41o66Pe4hVu7tePmdds0/XLG/gX6ghSLkJait8
WMHyF6zV/xaMyFB24H0w1EktGURL/diytf71qG3VR6eISkM9C3iQmc/6hMts56el
VWOH4R+NJh01WlQqdlBfEn0ISm8gwbZfOdoNHwMt7OpZpBJ9gdKcvBrVHWlk/cFM
2HUp+5V6eBw1pdBzXzr1fRDNWbQUgZrNhb/xGLgWr5xIdfRiggzkhzQ7xtjgcuf9
EoUvWXwsm7XQdBHkQ/zudHmf1xZc3hcfmzmQ5KsXRRHZPZ7G/Gu/gjzPalaXiAMp
IPuLTkHnwXp3AmJxHwdWsdOJ7myTVatAoU+ytvWYyc2wg/NSASKmjbrUYRrKovM4
`protect END_PROTECTED
