`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AbTZoPRKoAhaV2Fql6xoPp5/+HlHxJe+WKxg41YYnicvS2tiCZf55c0ixjjZBsgH
r4AWDDCytJKKIhbai3Aw7MdD6jqgTeATxm31YtM7INji4oFYNNM0v9O6cpYbscJe
xXqr9Fe8t+8i7HucCWriy0yJn+PwhHatCXQxFP3c1xhoaEojg/1jPhEg8VEYbRnh
NaNn/DstBtIFQ1RRrg30QeDwY83k5/j+Yf/KJZfRlPTCxNZnwRs5xDzFLVCVCATg
2rm3csse/9BKDeMhE+oo5ayvF4lccxfOeKVZjRgNnOqqXuUoS7Jmz7teFAJanhh/
3b+PSoRT7+C1eYUYcfWxociKaKl6WhBw6OTaV+ZmhDbBKMtx1IhORihYqgpmywJq
3rYdI7Wlg5sxVZwC79tjyYuPBwxoC3s8AJNX6i1iVJGA1PYW2ehU9w0c9p47PaDn
nQm6e2zWn2ehBpia4ByIbmVtTeREmk4+4QmRQoXTPJoisluXv3bg0SlGgIvChppN
sO/sJGuaqqZIg3cWlQRZpI/4HMvoS2Lg+Piih8Pt/eZ/AIjBhLwtEkmRCWTY8RUA
DjYMOqEaPQUQQM50WXhBcZwEqOeniDX1WdanZz5z3KwvfN+3wNSOZpjOVGiamVk/
vCSPosrxwPQIJX9VJ/cVLjhKrfzSfw+/+ED7V3JIRTQ9BCxtJil1Mm0RpNaEEC/R
5+AgNP8ueW8h+cLs1qU3VQL6k46PNvK+RQs+JyZxJ5XL7H+NV7kdCX9rs9ie9ox/
QncBUlolK1gat1fcLv7q/pX5B8xWXpWNd7i1CqXkaRo=
`protect END_PROTECTED
