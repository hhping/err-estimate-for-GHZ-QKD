`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MoVdsytrliFqg6BKGyuFLOpsSb1vdfupSZsR55V24CdmTnI17XNXLEEq7xWOz7U8
5HF3XBA9dD0FCzWfx5idoS+vucDgNVv8OUAnGM8CqzKo8jb6d9etkAKH2nrQwB+q
T1lAyRF67hGGkdek1i23IE2P4PfOzyLoi3UY44hquSUZxHaYyb4f5RX5L7AaE0Xv
o9Lj8ogmxKPxwrNXDYnZQtIJ0vOZybL57jGOLkrKPkt22yI3PoHneHdoZgddeilI
F1ar7f/jFxhKAqtyVX8lwF0Zxseooy7wZznggLO7z46jBSPiupsl36knqIyj/D7Z
E+K1F2fd4madhWa+Ue4eMA==
`protect END_PROTECTED
