`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jydq0ZGySEydfkLJw1zywW9GThJmA+xg/l3wRBD1iIJIbTYTuyAk6pczwALgn5Hq
4F7PRR4VV+J1OG64a4HO+/VET0D8Qsql3U6XARZ0N4x2iNprR9Qs1N2iMHEg1Scp
4vmuz5vMBbdQSbQemxau9MciAoc8MZS6wIZmmh7YkIAkRNwoXL66ixrpl83sxI27
DfwzYK81Bq0wLEs9JMvPQbAm6i4jV8OTTgEpR9BlY1WGoLHEZyKeR9zisisBN6fC
`protect END_PROTECTED
