`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4I+vEEp5ihW5rV8m7idbGo77aMxJOfXwigz8W7/mKuHQq3j9fKoE/nIeIT7FN2Le
IvY7Z9U2xlMJbbZKJqe6yK/wLSL/CzM5BXZ9RY5NWBIIgkxbiSownfH2nQjEA2Ae
6JPbBYAZwOoefh8O2HY8Y9NHgvoHZ6m3A9WzG8ZmJLXhOu4yJbfBCEGm9uMdvTp7
WbWTyP/ma0+Ra1zeTkpwOxxrB2SGc1IgoscgYujBvyADChaRCc2gTu5A4ML0A/X6
PYkIeUzZlhZOjBZPHY67LzmIpfO5Qju0H66SvmwgxhRWUyhgphKplJEkDbumYddM
nW2jMkCCtOl92pW7qOYBUmaajqwo68NndKtO9EJHzxDDud6yivHcYdgaQsw5R5fs
Z2bb0scefDoIwVDI6Uw0pntLZDWkHP3AFW11wjvjuqMsq9oMWeV755TKJZOkq6fN
Lmqc8HrmllOdg9GMc/vbZxje5311c97F8/WXM0CjnEw=
`protect END_PROTECTED
