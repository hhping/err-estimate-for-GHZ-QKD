`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pbl9SOR31s8e+n15iw1O/10fTzhrEFAIyvWr6DW9OO6wX0UOAsC+rFU0GAOhI+bz
ZDQswSHWcOhOcFX4vhAVgB9U4lLr4/eY+NM/h5wMb388o0yEka9G/dLOhepBBd7I
WieT6DygP3AnubQ2iiPnOhHj92UtI5FboXSYMiEkf0Wr+os5We75YuYYshRRPizj
E3J9gZpeiNQ9aEZNtlGDklJkTu599YQSgRkp2k7n+KdhpnUbVF4Ym9WpXIeYhCBc
EokHS3eicCbPHYUEAHCC7tIeLKcEEZe5NxOPCszc7w14T2sAbkvfyEuF0q6hyeGk
OooLOot6S0RkdzLJ4e6P8EjdF9Qeuhy6XfPzMZW8loWM9jMD6oBA3DKOHPmm2tqU
3DICJp7pKfTj4JRFtzTFfw5HpKt9xmztGMGgZEWaSif9LZsbtIilcF72gbXIKDtm
Ew/V2uFYuv0ytF1j7QyUvECmUrEYqeGBhKlzY3LvxBa1g1YNH4aBzYwr27CJ00vw
2BD9NBZ941R5wyRlOT88s+C5YIxUFheVB/lgew3g2hMJZHKilXKiYCl/LVuHZsgq
Zs/zHzrAGbmuD0CYDVey2suft7niqbnJ7xNFQGDHdNe2eIe1g9xD0yAxA1A6MfhI
ZnrlJ/3PWZ4Q4uNNJgxWle9uZcP+HFH3dXv60r46yDzeO5B8FPkURY4IQtqsI8lB
6YrZp2FyzSsmXWMMxjWi+UMLZOyuHkI7tRjcvalh8zRPz+l2c97jL9ohkSx0vn3E
J5MdyknPiq4Xp25xH83nBSa2aImtPTWZLvytYRVQ8KaJw6T3P7AjTqCbPuGhau2E
FXkP17Tqb+qpOiCGll4PXVyo0ZgGX0Gq535VVlYvqIavaEp5eOEbfrf4wCm1JPbo
A9OL3AIEjnYUeFOe3AECzZzEThveVXQDPc5E7DzzU6cs2Ff2aLvR9ypnUe03Fycf
Sm4c3YmvjDjYrFW1gY0GDAYTk2/WL0Tg7+tq2NERYW3n3Vgy8BHiPSPA1XsAOPAe
g/NCIroV9NXhRVShbofEvO7TW7OT7oycoTq/88GYmjKxO4ZzWE7v+pGMjRmxv8aK
Bvk5R9679jdNG3VZX/YPUpQZ7ax0trwStwMCuwVVK/kXuFq1WxzEZ7U5ThDbp820
S7m9k/EhTH9nrnr7E1ooE++PRMhDJw24NoAHs9jwoBEtngZHZsfTEAAeVqaCZzoF
R0+D91HF4KkzdtDHDP/oQ4Wq4HCmg86qDtOEuQT6ElGZhZD23wqHkOlk9e4l0F8g
ZZNkLz5xpZj/pBMarbaUcnKt2MO/o/F7NFL2q6mK3uegzrXOBOs7VOOok8yU8jc4
EFl4TJG7rz3EI4IcpURdD4MuwSWQU2xyy6GG+kmHNeSVM50lkGMfzyb+Yr9hUd/k
m3o+JuDgkAqj72Vi0vGfkwOjeF0id6C4BJz2TKSjQxqXzOw0q3vbNovDIJQBc6NZ
OFILLsWj0xUxkMXWNk1rZ50gI/xw3+A3S1ny4plrQlf/IO9rGNIS4C4y4pNp9sI3
UBjUcSjajoLqJ/GXI1fh8A==
`protect END_PROTECTED
