`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpxodpXkmtUmtYB3Gr3CkvJMN3MXiiE86RjEFiEiu9LodeJ1LE0CX0NGaE6wxk6p
Phd39f/TCsuIdigG0JPSTXxtqnmW1NflXGbK2OWasoTOwHp1kIaD2LX8/Gg3VQAx
tTwpn4+FK/FY4TtUfbtwgnPxLsC1A5k3y/nhwLef8z6lkBTuAQgJUKVKYljQGvuf
OjCiUpqe5OYviz9T83pLjouCQVCoV+a5z6LWAjt7VXy+H6WaUTyxepCKzmSixmqn
KUsZQUekkZ1vhbAIEqxJikCSXKSEzHIdGmeTRbSwp1K0YZb4eyAD6DNWa812jYV+
oNiMIQgelZuLQZREfjOVOZD47Zii26ccfFoa7v5SO/84aj4DtIa1zAdmaI0M3lXs
anB9+GWc7hE43Z/Bz98fdJsDvxkYEOjI0EAqddQ86sVvCSHNfwxtUlDyNSaIFJwg
eDvGz33J7adJhyq0Nlz+ip7OFlnOhr/4XxfBNaujEc3XJuW8H1JVRaNq//w5aYzv
WU8Swj+gs7rNAqvTf5qVLX2MkAz8RGYPqhHObTQXVE+JFtlPIHlXhottlC/LjZMG
3xRgWyCMfsFkRK2qgf6QWce2I87LaZmd5nKJb8mDEX91Vr5MhScKqiR70A/VKuEU
BKQD/syDEsmAIHBTzlzM6V4VlWLEfK1/sotKSJpQCMV53SM56+gxbN7Ft/VrLeZL
SHQab7Yw5g1gKUI0xR+P40OY+7nY53YMoIPq356Bo/aH8FgXatlbcnpq6aUjL8HG
gFOWshGfRqup0CZNhrLmWwuTbSzzU3jD8nL/M9aU5ojAhr5B2t94fKXGQ+vWU2mk
hIRGc6t7R+a80cmyKBLO+c2gErIryLulBudX+9Q/xoN76iDf8IQablKJnws4WjGh
CtjKskvDacUXwzcbLl20E63aIM7vWLjLc74YjiGDUNJ87N42ZpzoXnkGXEiAtWu3
Si7aYWhkKumIbw4B1LpFkT3PTKSg1/7XUELXHmx1YD3UmIIgAJzb1Ds0cw3+buzE
zw60LWrCzvJHCwcVPvK8dzaSBEieNLMYuNfaRFOh1/VsLXBg43URq42TxvywZTDW
ZvXCqB6d9RcBlRuNJ8WH1tGVbO6O3fFnbZGQt92WRnrqLymhoCintFCrcEbO5ZC+
yeVnobncyy3ghg4TMcARtw==
`protect END_PROTECTED
