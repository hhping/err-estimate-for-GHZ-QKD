`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9/MlNeyEkuVstu1dM3yBxwWlFWkBmXiEBMk/QHWylVpBThAvyWktclcdkLKP7LW
5Cav5n1N2jTQOsxvLKaLfAQOc8AW/OTqUaKBjzZuMaG0tho4g3pstByFm1xb1Dtq
I4s4ukASrtz9Li1Ye0N1V04mKoKU0hYmTdGSmGowqza01LWr8roP4gPILXK7BizV
nFpUymBl07qMzXj1G5iiZN2Qpg+9JYOTWaMvAZ+xs1O/AFT812BUNJfUztOLktPC
drSkvEJCIXLJB3P7bdDroIQFj117M6+rUsWYAF5SzYLYawV/r0IeCqW8i90nhqpq
PlUT7iSZ0/hZl3s1jV2X8tobekcs5NJEFq7fVLya1iDJV7u9TuZqAnJqPOZzFS5Y
0SsLlTnojVKG0YghlvO2M6XPApYIZul2UTd/a3S+Y9B+1y8EDPZ2cyS+DF0+r48K
aPX2iuvCqD7e2erjpj/pCaIH7XCMc3q2OtCrED8hGD0KDQCkmWxBERwwcqkyMn6/
ZAb75sAHQky9zURfzf9wh7CXpikoSSqw4OuZ5U45DWDyNyZxJ+oUQA2HrIAAersL
5UgWBgzKAvnxjj810iXn6V3/nSRX7bMMtjTcvFnyJ9W9y2yVRmIf7pIzdP2wNo4q
+0r7lX+UyvQI5EPtPZLilJ7l/NdQBUwlIpKgAd2Lncceht91ahk/a9W4G6F3zgU+
UIBLSlXV519ts8M1HrfTbu3628OKzZaT1RA92HudZD+SoDViRPaZwYi8Gf502EDz
pphLCwHrKiGuyaTl4pIJPcS/+FmraP3ClVrOe5lQAW+3hgKcQk4FdGuNNy03B0Bs
MT2aBvehJH8Iz3vontcC/gvujyecNOiJgkcAGdi65hUWzxyCS2OTTM7mHXtwwB7s
GemYTURrOEYJRCSBx/1pkwEXdC8SMH1dvbZzZ+eIJmg4ujQhKUaRR9W7KCYXgVNd
9B/YvjsahDqCUypRHmBqaVoFc1csWKjDRQ7DkFTkzOim5J/4ObMBhnklvr48zPi5
LcAWDrUoKjrzWLg7rsSQ4T27tYzods6n4zBkv+JGfyRqfJNbYwa0KD/rmNSCRG/J
dTWMDQ0aHJsW21QRr6S1uTBHz2WUpqV6OMD0mMC+5Gs6oGMPJym/w8crFlLK36gx
`protect END_PROTECTED
