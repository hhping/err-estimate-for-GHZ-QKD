library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_tx_pld_pcs_interface is
    generic(
        enable_debug_info: string  := "true";
        hd_10g_advanced_user_mode_tx: string  := "disable";
        hd_10g_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_10g_ctrl_plane_bonding_tx: string  := "individual_tx";
        hd_10g_fifo_mode_tx: string  := "fifo_tx";
        hd_10g_low_latency_en_tx: string  := "enable";
        hd_10g_lpbk_en  : string  := "disable";
        hd_10g_pma_dw_tx: string  := "pma_64b_tx";
        hd_10g_prot_mode_tx: string  := "disabled_prot_mode_tx";
        hd_10g_shared_fifo_width_tx: string  := "single_tx";
        hd_10g_sup_mode : string  := "user_mode";
        hd_8g_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_8g_ctrl_plane_bonding_tx: string  := "individual_tx";
        hd_8g_fifo_mode_tx: string  := "fifo_tx";
        hd_8g_hip_mode  : string  := "disable";
        hd_8g_lpbk_en   : string  := "disable";
        hd_8g_pma_dw_tx : string  := "pma_8b_tx";
        hd_8g_prot_mode_tx: string  := "disabled_prot_mode_tx";
        hd_8g_sup_mode  : string  := "user_mode";
        hd_chnl_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_chnl_ctrl_plane_bonding_tx: string  := "individual_tx";
        hd_chnl_frequency_rules_en: string  := "disable";
        hd_chnl_func_mode: string  := "disable";
        hd_chnl_hclk_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_hip_en  : string  := "disable";
        hd_chnl_hrdrstctl_en: string  := "disable";
        hd_chnl_low_latency_en_tx: string  := "disable";
        hd_chnl_lpbk_en : string  := "disable";
        hd_chnl_pcs_tx_ac_pwr_uw_per_mhz: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pcs_tx_pwr_scaling_clk: string  := "pma_tx_clk";
        hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pld_fifo_mode_tx: string  := "fifo_tx";
        hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pld_tx_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pld_uhsif_tx_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pma_dw_tx: string  := "pma_8b_tx";
        hd_chnl_pma_tx_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_prot_mode_tx: string  := "disabled_prot_mode_tx";
        hd_chnl_shared_fifo_width_tx: string  := "single_tx";
        hd_chnl_speed_grade: string  := "e2";
        hd_chnl_sup_mode: string  := "user_mode";
        hd_fifo_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_fifo_prot_mode_tx: string  := "teng_mode_tx";
        hd_fifo_shared_fifo_width_tx: string  := "single_tx";
        hd_fifo_sup_mode: string  := "user_mode";
        hd_g3_prot_mode : string  := "disabled_prot_mode";
        hd_g3_sup_mode  : string  := "user_mode";
        hd_krfec_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_krfec_low_latency_en_tx: string  := "disable";
        hd_krfec_lpbk_en: string  := "disable";
        hd_krfec_prot_mode_tx: string  := "disabled_prot_mode_tx";
        hd_krfec_sup_mode: string  := "user_mode";
        hd_pldif_hrdrstctl_en: string  := "disable";
        hd_pldif_prot_mode_tx: string  := "disabled_prot_mode_tx";
        hd_pldif_sup_mode: string  := "user_mode";
        hd_pmaif_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_pmaif_ctrl_plane_bonding: string  := "individual";
        hd_pmaif_lpbk_en: string  := "disable";
        hd_pmaif_pma_dw_tx: string  := "pma_8b_tx";
        hd_pmaif_prot_mode_tx: string  := "disabled_prot_mode_tx";
        hd_pmaif_sim_mode: string  := "disable";
        hd_pmaif_sup_mode: string  := "user_mode";
        pcs_tx_clk_out_sel: string  := "teng_clk_out";
        pcs_tx_clk_source: string  := "teng";
        pcs_tx_data_source: string  := "hip_disable";
        pcs_tx_delay1_clk_en: string  := "delay1_clk_disable";
        pcs_tx_delay1_clk_sel: string  := "pld_tx_clk";
        pcs_tx_delay1_ctrl: string  := "delay1_path0";
        pcs_tx_delay1_data_sel: string  := "one_ff_delay";
        pcs_tx_delay2_clk_en: string  := "delay2_clk_disable";
        pcs_tx_delay2_ctrl: string  := "delay2_path0";
        pcs_tx_output_sel: string  := "teng_output";
        reconfig_settings: string  := "{}";
        silicon_rev     : string  := "20nm5es"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        hip_tx_data     : in     vl_logic_vector(63 downto 0);
        int_pldif_10g_tx_burst_en_exe: in     vl_logic;
        int_pldif_10g_tx_clk_out: in     vl_logic;
        int_pldif_10g_tx_clk_out_pld_if: in     vl_logic;
        int_pldif_10g_tx_empty: in     vl_logic;
        int_pldif_10g_tx_fifo_num: in     vl_logic_vector(3 downto 0);
        int_pldif_10g_tx_frame: in     vl_logic;
        int_pldif_10g_tx_full: in     vl_logic;
        int_pldif_10g_tx_pempty: in     vl_logic;
        int_pldif_10g_tx_pfull: in     vl_logic;
        int_pldif_10g_tx_wordslip_exe: in     vl_logic;
        int_pldif_8g_empty_tx: in     vl_logic;
        int_pldif_8g_full_tx: in     vl_logic;
        int_pldif_8g_tx_clk_out: in     vl_logic;
        int_pldif_8g_tx_clk_out_pld_if: in     vl_logic;
        int_pldif_krfec_tx_alignment: in     vl_logic;
        int_pldif_krfec_tx_frame: in     vl_logic;
        int_pldif_pmaif_clkdiv_tx: in     vl_logic;
        int_pldif_pmaif_clkdiv_tx_user: in     vl_logic;
        int_pldif_pmaif_uhsif_tx_clk_out: in     vl_logic;
        pld_10g_krfec_tx_pld_rst_n: in     vl_logic;
        pld_10g_tx_bitslip: in     vl_logic_vector(6 downto 0);
        pld_10g_tx_burst_en: in     vl_logic;
        pld_10g_tx_data_valid: in     vl_logic;
        pld_10g_tx_diag_status: in     vl_logic_vector(1 downto 0);
        pld_10g_tx_wordslip: in     vl_logic;
        pld_8g_g3_tx_pld_rst_n: in     vl_logic;
        pld_8g_rddisable_tx: in     vl_logic;
        pld_8g_tx_boundary_sel: in     vl_logic_vector(4 downto 0);
        pld_8g_wrenable_tx: in     vl_logic;
        pld_partial_reconfig: in     vl_logic;
        pld_pma_txpma_rstb: in     vl_logic;
        pld_pmaif_tx_pld_rst_n: in     vl_logic;
        pld_polinv_tx   : in     vl_logic;
        pld_tx_clk      : in     vl_logic;
        pld_tx_control  : in     vl_logic_vector(17 downto 0);
        pld_tx_data     : in     vl_logic_vector(127 downto 0);
        pld_txelecidle  : in     vl_logic;
        pld_uhsif_tx_clk: in     vl_logic;
        scan_mode_n     : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        hip_clk_out_div_by_2_wire: out    vl_logic;
        hip_clk_out_wire: out    vl_logic;
        pld_10g_tx_burst_en_exe_10g_fastreg: out    vl_logic;
        pld_10g_tx_burst_en_exe_plddirect_reg: out    vl_logic;
        pld_10g_tx_data_valid_2ff_delay1_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_2ff_delay3_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_2ff_delay4_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_2ff_delay4_plddirect_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_2ff_delay6_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_2ff_delay6_plddirect_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_fastreg: out    vl_logic;
        pld_10g_tx_data_valid_plddirect_fastreg: out    vl_logic;
        pld_pcs_tx_clk_out_pma_wire: out    vl_logic;
        pld_pma_tx_clk_out_wire: out    vl_logic;
        pld_pmaif_tx_pld_rst_n_reg: out    vl_logic;
        pld_polinv_tx_10g_pcsdirect_reg: out    vl_logic;
        pld_polinv_tx_8g_reg: out    vl_logic;
        pld_polinv_tx_pat_reg: out    vl_logic;
        pld_tx_clk_fifo : out    vl_logic;
        pld_tx_control_fifo: out    vl_logic;
        pld_tx_control_hi_10g_reg: out    vl_logic;
        pld_tx_control_lo_10g_2ff_delay4_fastreg: out    vl_logic;
        pld_tx_control_lo_10g_2ff_delay6_fastreg: out    vl_logic;
        pld_tx_control_lo_10g_fastreg: out    vl_logic;
        pld_tx_control_lo_8g_2ff_delay4_fastreg: out    vl_logic;
        pld_tx_control_lo_8g_2ff_delay6_fastreg: out    vl_logic;
        pld_tx_control_lo_8g_fastreg: out    vl_logic;
        pld_tx_control_lo_plddirect_2ff_delay1_fastreg: out    vl_logic;
        pld_tx_control_lo_plddirect_2ff_delay3_fastreg: out    vl_logic;
        pld_tx_control_lo_plddirect_2ff_delay4_fastreg: out    vl_logic;
        pld_tx_control_lo_plddirect_2ff_delay6_fastreg: out    vl_logic;
        pld_tx_control_lo_plddirect_fastreg: out    vl_logic;
        pld_tx_control_lo_plddirect_reg: out    vl_logic;
        pld_tx_data_hi_reg: out    vl_logic;
        pld_tx_data_lo_10g_2ff_delay4_fastreg: out    vl_logic;
        pld_tx_data_lo_10g_2ff_delay6_fastreg: out    vl_logic;
        pld_tx_data_lo_10g_fastreg: out    vl_logic;
        pld_tx_data_lo_8g_2ff_delay4_fastreg: out    vl_logic;
        pld_tx_data_lo_8g_2ff_delay6_fastreg: out    vl_logic;
        pld_tx_data_lo_8g_fastreg: out    vl_logic;
        pld_tx_data_lo_plddirect_2ff_delay1_fastreg: out    vl_logic;
        pld_tx_data_lo_plddirect_2ff_delay3_fastreg: out    vl_logic;
        pld_tx_data_lo_plddirect_2ff_delay4_fastreg: out    vl_logic;
        pld_tx_data_lo_plddirect_2ff_delay6_fastreg: out    vl_logic;
        pld_tx_data_lo_plddirect_fastreg: out    vl_logic;
        pld_tx_data_lo_plddirect_reg: out    vl_logic;
        pld_uhsif_reg   : out    vl_logic;
        pma_tx_pma_clk_reg: out    vl_logic;
        hip_tx_clk      : out    vl_logic;
        int_pldif_10g_tx_bitslip: out    vl_logic_vector(6 downto 0);
        int_pldif_10g_tx_burst_en: out    vl_logic;
        int_pldif_10g_tx_control: out    vl_logic_vector(17 downto 0);
        int_pldif_10g_tx_control_reg: out    vl_logic_vector(8 downto 0);
        int_pldif_10g_tx_data: out    vl_logic_vector(127 downto 0);
        int_pldif_10g_tx_data_reg: out    vl_logic_vector(63 downto 0);
        int_pldif_10g_tx_data_valid: out    vl_logic;
        int_pldif_10g_tx_data_valid_reg: out    vl_logic;
        int_pldif_10g_tx_diag_status: out    vl_logic_vector(1 downto 0);
        int_pldif_10g_tx_pld_clk: out    vl_logic;
        int_pldif_10g_tx_pld_rst_n: out    vl_logic;
        int_pldif_10g_tx_wordslip: out    vl_logic;
        int_pldif_8g_pld_tx_clk: out    vl_logic;
        int_pldif_8g_powerdown: out    vl_logic_vector(1 downto 0);
        int_pldif_8g_rddisable_tx: out    vl_logic;
        int_pldif_8g_rev_loopbk: out    vl_logic;
        int_pldif_8g_tx_blk_start: out    vl_logic_vector(3 downto 0);
        int_pldif_8g_tx_boundary_sel: out    vl_logic_vector(4 downto 0);
        int_pldif_8g_tx_data_valid: out    vl_logic_vector(3 downto 0);
        int_pldif_8g_tx_sync_hdr: out    vl_logic_vector(1 downto 0);
        int_pldif_8g_txd: out    vl_logic_vector(43 downto 0);
        int_pldif_8g_txd_fast_reg: out    vl_logic_vector(43 downto 0);
        int_pldif_8g_txdeemph: out    vl_logic;
        int_pldif_8g_txdetectrxloopback: out    vl_logic;
        int_pldif_8g_txelecidle: out    vl_logic;
        int_pldif_8g_txmargin: out    vl_logic_vector(2 downto 0);
        int_pldif_8g_txswing: out    vl_logic;
        int_pldif_8g_txurstpcs_n: out    vl_logic;
        int_pldif_8g_wrenable_tx: out    vl_logic;
        int_pldif_pmaif_8g_txurstpcs_n: out    vl_logic;
        int_pldif_pmaif_polinv_tx: out    vl_logic;
        int_pldif_pmaif_tx_data: out    vl_logic_vector(63 downto 0);
        int_pldif_pmaif_tx_pld_clk: out    vl_logic;
        int_pldif_pmaif_tx_pld_rst_n: out    vl_logic;
        int_pldif_pmaif_txelecidle: out    vl_logic;
        int_pldif_pmaif_txpma_rstb: out    vl_logic;
        int_pldif_pmaif_uhsif_tx_clk: out    vl_logic;
        int_pldif_pmaif_uhsif_tx_data: out    vl_logic_vector(63 downto 0);
        pld_10g_krfec_tx_frame: out    vl_logic;
        pld_10g_tx_burst_en_exe: out    vl_logic;
        pld_10g_tx_empty: out    vl_logic;
        pld_10g_tx_fifo_num: out    vl_logic_vector(3 downto 0);
        pld_10g_tx_full : out    vl_logic;
        pld_10g_tx_pempty: out    vl_logic;
        pld_10g_tx_pfull: out    vl_logic;
        pld_10g_tx_wordslip_exe: out    vl_logic;
        pld_8g_empty_tx : out    vl_logic;
        pld_8g_full_tx  : out    vl_logic;
        pld_krfec_tx_alignment: out    vl_logic;
        pld_pcs_tx_clk_out: out    vl_logic;
        pld_pma_clkdiv_tx_user: out    vl_logic;
        pld_pma_tx_clk_out: out    vl_logic;
        pld_uhsif_tx_clk_out: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_advanced_user_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_ctrl_plane_bonding_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_fifo_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_low_latency_en_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_pma_dw_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_shared_fifo_width_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_ctrl_plane_bonding_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_fifo_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_hip_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_pma_dw_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_ctrl_plane_bonding_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_frequency_rules_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_func_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_hclk_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_hip_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_hrdrstctl_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_low_latency_en_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pcs_tx_ac_pwr_uw_per_mhz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pcs_tx_pwr_scaling_clk : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_fifo_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_tx_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_uhsif_tx_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pma_dw_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pma_tx_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_shared_fifo_width_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_speed_grade : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_shared_fifo_width_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_g3_prot_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_g3_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_low_latency_en_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pldif_hrdrstctl_en : constant is 1;
    attribute mti_svvh_generic_type of hd_pldif_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_pldif_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_ctrl_plane_bonding : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_pma_dw_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_prot_mode_tx : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_sim_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_clk_source : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_data_source : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_delay1_clk_en : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_delay1_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_delay1_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_delay1_data_sel : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_delay2_clk_en : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_delay2_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pcs_tx_output_sel : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end twentynm_hssi_tx_pld_pcs_interface;
