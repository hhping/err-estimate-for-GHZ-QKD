`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1oRtkMN+3MvxQ+Ba6KabuLb4fjcux5M5q3ZCM1+P4ZVt1W8jDFtCPcbdOM5sZzau
HOcoLam07YQjgX4B9TdKAGCgjwDhKACbBlSBAbgO02LFlmzLtTGPVSpmZ4ikNB9b
2ceshZMPAvSQpL5AC/Um6qXnxCS+1/CGRHrIM8kuQMkvWFFhZC1FBYCb8qyL3d9v
z7KRRdaT5m8uOitL5PCdY008Pp+Iz5jOS198jiusCdrRRrQR9z80ZVKKXjQFDikC
5l8vv4cVFjHu7yPlnUGmfzvssorALnkLTntwADxFXqQ9RYLZMotWYIazoM5KvdCF
z8kcUIWzGfv78kom/xfX17ivPAXCPofmg5x/E878EK3XSPAhLedBUNeaK7fOC3+B
nbzl1aB83lEYDvDHcDc9FvXpjL731BoenCMn9QAGM+uVinYFV3XyzFmzC+o4VsNa
etCSmpI3jW6b8YRg/7ikowTKZStjmblu4ZgxKGAMuovl2T3cZ9brEjAlz8Iqx+av
rFfzwND864DDYzDB7OnnB/BanG5DKb6UlEIHvuC9KCXaPJmEt7Xagds8WuYN7lno
oLbxLqR+z8L2QI4kPTazZz3RS1OW7YcIXlkWLqfmDqoyfX2weLJYzRE58EJw1H4O
BY6cBp5MSIRIFhXyNLgKMageW6Lx1DzLnrZGqCxcxTTGgCPnEtzFtcbUphAI/XyQ
25UGlvlyqcaeKRHdQCgeQcLjjp+TLMfFoJb1ImgVKIHizlCJcA3dViJWLD1+DUfE
`protect END_PROTECTED
