`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X09hdcNWSWEj60xSkd/7yXpRPovhdPzV5PSbvKeORDIe2/PNZOQ4G3nQHiUuCTPG
fWYGZpQWgI1xvlj1X0nMBQxfByZ14JM9duJVWRqKJ3H52OlC6VZfFUnJvyPdlkQu
CwOfx4iG3rKFQZ7HSq3TuKCtNIW+hVtN9Gkql9ns6T2AuMDUqkbNxUOlGtZD5aWs
yDcwsTdJV2UJgKl7zog33gkH8eVc4ljogIvE/BVBvD6VnWWefV2VSlfiyLyWEAya
A+2LMoD2KuG1pE9rUm3hSts+GNG1gUmf3dd4JOsQUtmByZo/vhX56x3aeAJuYkX8
MiNSdlfy8u9JiRkgS2bzNZuvq9+2jc9xycQnTedvcVr62oz3DyKt0KkXt83CnKBh
gQeHpH0U8LGWXCTFo+PuxJ61vDRs9VxpAUvACJ6LdRdAAfbBeS7oRq6D8YtTkyky
zIXlALm0F8ERCAkIO16eLoBoGDW1euJL/VlCc6PUubxI3olJLhhlJStchOdYbwLj
IpCSll5lq3CyT7n4FA4gltu7cFCHP9npXrZii/DtF/S9eGHx1AYvdWECie9PRJ33
xx2yNFptzKYEFmizZTMkdTzo1kIFeM2s/gOhSLVhdoX8cGMU8iI0G696rorjUaDQ
XqOBzdDcQBlpf+sMVM405J423wonPkhehIrBqJxCltpK+GzZhg1Wn+RTNpqQsike
zcBAnoURfQylwMtymoj4xvF7FB5+GM2kaR+w10k/fJiiRDrQVGqEfu8Fw06CJj4L
ewP5ggBD0MglU2NQkxTCWLmsNuzJZjJUHQMMj31cfcbAWOkP2WRGsKs3wAg9plka
gJHRUygVsR0rYcR1Tj08lnWGvaMJoomXlcVxLbQpeAdm9xFgGzT2ovX1uLkBfa8c
fUCjXQtNEMJt93WGq3UKISG0hPRqQJl1rI91sOLf04tmXE/JdO5vW9jDtOsDKIst
KcCu8lLjTYH9xg3PgbzWYn4sT8nllRA/Hy7GB+eBzEu19FKIFcOrfQSIQJRsHIx1
zpUy7e7zrc/Q66k5AijkJFVTvDRyol79ryol5EvQMr0nECvFuvl+oh+aa5NDt+TJ
UQCbTrstmtir91C8Ld35toYrSjNURXNTlitkRm/rmngR3rZ5JnkAu5NRGONkh9wu
f7+1ttA3Gmv6bmvRks1hAWkGE9rHHRwVqvRSRZWqH7ygPeldgpbWW+xlXQf6ik/P
+BtEbR9BAO7zZSscI0s5ldJ9TpCU6I1+0roxg+2iQn7IWvoI5qlKI39k287hneH2
6k7LqD/DN1uwHaHDRmD8v2951obX+hBuL8L3wlBGVo4WcBgYJZdhqxeUpzonlwak
dS/TldOgnJAZnkeO51EIxRmolrQwLLlBEWOL/fxZjSTbZyJ+LZYJvo2jG/HM95oN
7BOztK7+ds6JDGv2vhH0LdbhP4TKoqQkk6pBzM1AeK8pCzJUirMOtQPTz3r26zkQ
xnxxS+oPM9J/x5vW67wxpqBCOwvQPvJljM4LgWqTkPkSeB5jwep+Q1o1H2f0fB1c
h6kSKGcYFCFA3GrWT/jh+DyFn+KkC2GhWT0PrSyqSs34xkrKygHI5liWyvi2ThB0
dZMvtgKYvN20eYbEoM9MWwGoVx/JQtYOcEsiLZdTxQgwZTQX6fIaXIpPFiHdM+Nc
kyCsWINM7zjvBNaqe6jyMcOfH+Kgq+qLh4kyyL9Y2GOkyIj3HTfs5A2oHaPx7/rq
0v+70xxEv6dZe7LpzpTwgyp3n0yqKwgb99aVHhtnT3kS33KlOHrBIYJJZhCNQTz7
+1JGZOmirzgOhqT/avO6rtg+pqHh9u/Ft4UZkqNkZpeP9iTphMd0VDhG8Ib3cL4Z
KcKBlOSBTyP5kAhNd+lpVtHo1Qfjt5MvPr8Ln9xXbX7zvAKUMP+IL8zEYfbzz4PI
bsVxU4GweNrKEO0SJXl1FkyhvtiYmqdAsgJ1YMNcWT8MRDLWbG/+JXBCNc/S2Ai5
EiEkM+2R8SFdqjnO+9v6+0At3izUSxTcvWiIPFoWIJWRZ0fCeppr4EAozZF0wlBm
8nzIakBBzGXIo4NhOqv+obOBuIuEAjonSTjE1XRR2XDG+aKVlrhjIimdi/GzSsP5
UiCsOAwFp8QaUEWqhlALDKhjWYZvA0lh2PFvkpn8MNHEhpKnbqNyLGUVFIHVFmG2
fdjIyWwH6TtrE8Fs538/8gCK/Nq/2gYWkF9bE8JpZ0XIWd73NZ7ZpxraRUp+fUWm
LJRIVsDeTQ/sToCl/GKu2JWnFX+A8knUyf5eeIF6PRPAKtCzVGzP5Rgi6OSn3JaQ
jsEL7m+UTdQhltqFRhf+s6xx9tFfjceMBE4ri0Gpbr58gXCjMr49JvfZGLxGjzcg
O+k5HpkA1sD29WQquROLk5IGOx2Ksb3LDc1Eb3polUi/sRgnBZ/O1FgVQeXHWUpw
jFJqUxBBQiJC0LKmBeDBm0nPRSjXDpo0/xLt93NODKPgWMG8+GfvED0QnxC+f7k4
6Uh25hVnqKZYr5HhEacw0uq974Y74ornlF1kJ+x0NSAKokwIdc4IdvoJ+nHTNAGn
vWNkAqxDo2LdqhkI4EBNVNt3nRSfaCHwpBB2lmmgiO7mWRGSLAFIMi5GZ02nj4mn
IvMVe89qOCa/YNItWwMjP1HlJJBkzzxrtrNyJjFZqOfu10pl6dmkh1+nDbPDEYqM
S/XBz+vBv11hiPobku4Sf/rIYZgKDLMtHjfMpmD9WB+IpSF5BICptfjgVees+TwD
rdVGtUuI+2WoN2/5qEZB5DxPTXQuqkF8M8BJWNeo424d974coEolFEJW/wwC/86J
38smXp8t2h9Vr/rY1JVwc53QojL0dOivsuAu/00MfIdu9GJuDINX1bvC0ZS5FYlU
Qufff4kbyaOE9rKFTPoNkcma5kBwBlW5ob+xWmT2A1jR++rNscOzKpJOfecP9H6U
wl6ptAsxu0R/RV0fTJe1Ndo8tMaHfpWjL6g1+Xnw20NGLRDu9tVOUl98j/7ELqIp
y92d2ri8tnVNVOTH1qHEgUGsiCum2Q7IxFp3iXjO9YwnRbz+OCyoyJ5Pt/jV+uG3
77kWDKRAviIeaf+bcaMt1cF3h5qcigG5xUWHkurBeckmrKeoMqOBVHQc/5UgXLaj
iU8Vmkz3WsWk1gucYfhhev85vGurGQGOlcJFrWhModMcWlvQQdX1zB27FQeOq8bH
1LSkNrmfp5oIwqx7h9espqOvbdWHJ0G2IjGiocomsXQNFdE26SmXxwOvGm2t6+9j
eh1nbogg7Vk9aLT6pNweevTHRZhJVOMYOuWDRWlZY1XItt+NNx+AzgPql1cZ8Cc3
opGX8caJuoE324dD0wiRG+R2EwjgZX4/ntzI5jSh2Ls67dfiq84M01FYJadZK9l1
9LXIcsFg8YXAZZLBQ43NK+uuybLlF3/TlsW8lOVzE/6ecaqkgGoQFxmUHZ9Vm5Qi
MxPfcWGKHw8/MRbCEa5p30giJy2lsgXFSa99LqxvVdJ8VlKpWexLvb4KWz89JIli
GpXP7aLBwvFI39DqUgAsbBmWc/GA/mHbpCAgTJcWL0Gj+qzW/maJZrrF1jyIwHGM
DxU9KZnNkQf58F0QrC/Zvl5cwkvCC9V1MmcSRwPFdN/8tzHgFvpa3RD+WdEPlqvA
3Sklj3pckZK29rAdn//JRzUsxfMCV4n0vt2eEV7xLcYGKhL6HQ+3i6UsG661wXyt
cvNABFkaurQU/6CnrxSIa3m2sar6MphUD5RaXmK0byr/zd+MlCfC/l23V1I5ws92
mF0lFcm+nkslfSw6UNbS8GU1QeiyXFHwDeda0NVfZW9ptkCAM+loe2gxUcpu9DKL
obrolisIf9XdRnfzQgNtzNJUUlj4p79Bd4DGX1vO5pz47n6v7nO8Aoh9OLtdiDFS
B7h6vFHzJfAFGWNPoIZjAToaWYXwPQf4TVoWv8S+IxJDTAYeQZRqPB9YO5xb3z42
B7O3Xq5cRxrHHdc7CSRoJO365O2dUYLW6wEBwVfEN9k=
`protect END_PROTECTED
