`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URdXuf2JljYUXLrty+uZjWqw37OAqodGYj7qi3zaekTeq2hoIlaVNXvHRAuVaQhx
aBwAMXwnWDYcGIxb/lOm9+qWIfWmlj51lKxihi6/+yTr1kfVjgX2n5fFqwBjKfx4
BUJUrHySsraqLhkVRBAo10FX8oa4IhXybhvPV0Ivr7m0SfbZj9cdqHBqcOThHiZj
za+shw7RCuR4lC+QtlZ0bTEQzz7VAG1qBCWPD9DsRaWoIUgsr0ZU6tMWfGjrivrE
U1Uu1kWCGbrmd+ZnJ0k2edFhdLrcDVCOnI7nMeN8sxN4qoZN7f1gHVR0U659xDCK
0WFrfOvH0+0G37oREqIYEGuq4KX0pBI10MsDG1WLnwiX7WQr+iCBw66VI9AYIA14
FfgkM3goULQz2pN29eieBR0cSy4ELZZB1QA7iRdYCbqdaC4nD3EgVC1Kjb4vpow4
HWZxLiKEu1L8ipVJG5kzb6rimm/qGK7PVvsfsErDWw1aiqO0Z9vPxbyrgew8KRgU
KC1QsFpLSXjlebnbtZESpNVasPdExoP/Sda8oj50UC8qbmx0TLQxFqSHmBz2veec
y5qBKQ5tohYAJfpMSigdjswnL4Ky6vjSgY6+cAJH7R4eyuz+ppstKiV3DLuezKf2
Qak1aH5ZHzBvHWcrNZ7D0FZax843Q08bsalZ3qnTccGZAxS62vEacDnGFAmA95I3
xFug+aHP/0h/DuVhJ3jGW3VICC5lGBzS+I92hkHmEKFg0349TMYXjBBfDSQdLKTu
/7Mn8XjLHuXxcaUXTXVmxriff12OEf4Ml0t2kMkQeEfFzx8fsrW3DDvVjvrdIfx8
VMtZu03h3ND7/LjnRKWZ9lIe311jYCMTaBV59rfqHIXni6w5qQIMM4x7TmviRnan
V9+qA8EG+R2jZWzw0tT6Y8o9nJOp5ZXOYNx+Mv07pwXBhyJQUqPsfWmKkl7QXAJ2
J5+7DjBsvHJzAt+R753HX1N7s9BAcM7byXDFNU//AhkiKx7tokMaCG1UfOGToQDK
Fkf3ZK8KoJCRqbcHaJqQtXJpMieQ7Efr2OjRa3NYypGoYuZFyLYMKpkO7uyjcrU4
hcBbYu5xtBagenUL0QMM7oZFoYEn+RNBSUv71mOndTR7YC8Zm6VsklBwBxZhqwK5
VVjoaN0iHb0rUkq1B4K1y0kUWkd72BB32iNYj5li9lKWl9/n9kmQMzvf0+uXWR3T
GE0YimvN+X0qsym8yqU1+Kf8ruaTFLGSSsdDHfhcGs3efDF2uYbKjsM31IFwQAUu
T1jlMVJ+zTYxYL9b8qUpNZtvmfFbEd2wWNfrOOHu9uH6BU1rSd0sY5G5O8czV1sZ
4fH3TrAntPjWBOWmzxJh9zuYxrL07WN4tI9WBgKSD22qGspceIWV4W4Iy9Q5cgK7
fbW3GBViGm9586IG6F0jpca07HoZuQWYkeSiQBDuQ+wpbgFtm2j41DLnDLLj3XN2
0d/4kD3vvLw3TfQNiAbxtRotusUyNL2k2jnQ+28njpc7n0UaSi5xYPUxTscuIWXy
YKtJqHq6xAA5OhvgKs3EnPEqBdLToIzw4l+TuivQUtAzBFqK21zC5i0MZ9CV2Lk4
EcET4g+RJV8mrkKld2D6egMkXpAdhYWZ+6F5i2tzMbSno+U4GJzLZjLsgyDEMXFo
rsumCFGeG0m5xcmEgLg0dWO5uA7XJZFohbIpBgHGfVdFRMoESaFUMOTZrR1yvF1b
UbUMPZ6Egw90X5O2o/yxxd87Xlu0o4UmPMVM85LHvIu3vJrm5hUWa4X9qvy4eFxL
HXKVX5Lnb7Gw9L8ZO5tRUvGrirkXXKqVhFLVMQ6K408etk7PGI0a3PCQstnushju
HwNRYjCEtrSYwswEjYwnm7f4BGrx10XIxYy65p6v/5UaPlTMUhtEKpw1LDf69lXq
7Uny35Db8wZ1cYr6LRB78gyy2kLFSEe8Oe+sq9SUb8IzIJZ1cJtIO+VPHVpueF+T
mL4NHaCNY+quzPYgpqKm0srhIaQq9KsOX/qrVERNjbx4GH1d0JysdTFEU9lUtgMt
ytIaul76tLmq0iFMmJXCzH+aZ7tf7niGFyfmE/3aTfyHqXI94WFqpLVsE3t7IIHC
yHp2q9IioT0h9U4mdHzaUYDQUWm7JP+bTcvFqr+vMH1lra0d7LV6wNCqf3k30WSK
qoxdPYI+p6jr9wcm0Q5BQVQLxq2QOpFfetD4v1pMo4qD2fuv4mavackaUVOfjzAC
BmE552L85cjM3HH7Bej+y9bZZHxDn8wxRTR4cOBz1oe+yfvhokGb4Kkh9Hs9sADN
DQq0/81hwphU5CS7sIhDea0sSjd5wnvNjYfywMrzw0zLmi9ZQoYQoczRGQr6gZ12
I+lG4Y0y3aq8SXNOXUdnyPLk8/nWIgnvq+qD27nl+pYZzP1wWeg1reriajUIUkKT
0Y7O8ouwtI3B/t4zbexcAda4N8TiIOB35FP+V+5etJ4ZIGAY1Dp1jHXaaldgzTvY
N/y4YcK8Q1OvcGcVZh72SkrsEiDCCqKR2rV9gwEE8c0e/NyY87lnej7WbTTKYiV5
jq87XZXmdpufUMXcn/LMOV/qAweR4PeQrRvHEvhGbFLsk4AXzeGO/+WLg3Orbgc8
j2K+53GX70u+DVsHfH6z5Gji9I2cSAtWmchJqZAgZDMod0TyiZoORPFNJXrLxINH
SpmEA2PlfkKccNPvUJRVT3Kd24hF+AyXtAfbpEVPeoOi0TD5OIy+B/Qas4SsIaWg
/3p0GUTFAGMbFvKqH2f3wmEFXaqLatMmyKokr1idyN+5cgff+JGv4Nc7c2vSzI9l
rKiwp4Efa9XwKb83vkUFZ3esk6SPpnQjeH6jbcS2cVjT3musEdyWgSaxUCxtvzjG
Vmj8Ui/e5fPjma6bv6j690gR1TCR8B7uKAUOCJUkJ0BvzkTstsyFWVGA8tVEqyhw
2+9w8YOqdKQouzVYs7vx0CRWrQfv4VtPn3WgMhvqNwTwn9VmKbNHZP7vCs2ecIhl
eft7s4DXxcYUB0Y8ZfDgtmCHQT+KL4qmF6we2OyLTrlnfJ29+w0YaYN6MSeTWDyO
t+UIlOnPMWtriwi2IAMWFb7szpryppKDF3xZy7ByQGIMkGConDAywXnKTsXJJHuc
XsVQHpU3sa85lPPTQWasF+lq2QaraqaI9DLRZ4Ckem3Ng/cLoRVnCw6qL9y0ZNWX
zka5QXNN6y8lFiPMSL3XkArKx6uBYO3uHrgBq5JJKEdJI97hAslcnR9p/Or9XU+I
AnQeQL+dC3KUGQ5Ra5IU4j8il/3cyhpAy8M9CG3b7rNpPODip5cZFmsgVJ4+Au/j
U2HlD3nahovP4QtGjGBWCxNMY8NMq46+BvhedyGpo000vuNwaXEuICltVDGivscw
o57lTXFdR1Ztm1YKlQaeayBLizi4g4MmEyo9+RIC0NgWs2sQ4Aia853QRoQV8aqn
G9JlmMAbeD82A5WfeYqUIErY2WGYhS3aSrMh054z8f6iw4bXu7swuT7FbXLA5YnK
vE6FRJnvRAhj6We156cWflmVULwSWfPeNTETgsX8OpyJOiWZhudQBWZzOG5ywe8d
eHfmwJGnh10YnT0zPoe8CvN8+Dh402EDnrowaBlnJt2PqPb+SA3RrTqFcvRwQTQQ
liqKwjwCbE8JgsCNh3FbRTXfjmzVmf1WfPd8ePqmYcGyPMpCeTt5ZlMOZ2TavrjQ
3RDfqob5zxqyGAZ5DNDHnfU7k4yDmPKG4vUw3GKofdRSMuNdq8QBftTxZ24n/pc/
laK+1koZO81z3iQbj/UQOvyAetBrhN3MmGLWh5U6XR/EGv4kcEs1lQRxEjSO0VwX
LUZtC86W+TfnJGZrkEztnC7I23giX80Vh21IixOmMzuahuuEz/9C9mTAoF0exZPN
KiSO7UEroOAYduNtP8mzHZd4u+CyOqukjG6kot2rEnn70SJBme4IWfyAg9XPmnlL
`protect END_PROTECTED
