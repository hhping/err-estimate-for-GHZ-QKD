`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ko5uoutprbYDcxGnAav68TJBWd0AgdKQYidYWNbZYYT9WLr20DDcRNCxe/sYprRc
XTFIy3cBphk5kyv4AoRyPxpi0JM7vrWX7nGJ6dpbIgpQJtHGpQpTLFTPHs9WGYyH
uezyJUMpNTzFadlySwgOcEzjidXQtlHdyppR6kRQpx8/FyMdB8MSGkXprlC98Fw2
v2xfUEv1eS0Q0pzyVhDYgAhp+5Qi8O03jk8ym6DWIL7CecV+HrYYLZow+oGmCu1c
NMmoAjSnnpR3yH1uGYg6+LehlgNv1vqGYO7vJ66WkhCzjCHhC4pEDG1dYEK88BEU
PNWoZ8Gj5TWrLBO6G1s4+TK1KoYpHZhli0sjfKhehhJH7r/8Irz2mnhmv4yfKb2q
AiXjJ3vrpkzI8xNuaPxK3AL161tnMqttFyjMcJDrH1DfkbxW7gm4oI99ZIw90fNi
zmdUQNObRezhSihlrJsgLURXX0iWlruwZdurNNGe5Ln6qUU4q6uNnKepr7927aGA
LF+VXTD9arrjbSNjt8fuDgB2inp7y2lqECAinOTFBwsci0JFACoOgQTk4z2Wtoqu
mm+VOh/xlXKPmZR+5GsuE7jl4f76ZGPcTDiC6yoD8dUkMDZ2hj06wb02qO7cKakv
o421oTtIVN2cd39ufj0RiVIaWVOw2C/3JA2X69n+7VM1Mhea1wR1ul3mR4BiPkzk
wuht2kb/KgyitsOsS18oPVkjEicUswHALp5qsC0D8aY6JFLXrEAW3SYVgGp7ihMn
LbtLi5tncnfh+7s9yyr4S4ISRTdCz6kfvoR7Apevhqa+RT1ejANuJ9IWJgCWhePg
KWYt44utUf4ZBuKbN0c48UEFRbq1wTd+fH2+wIqHrO6ZtmCISZv/Ol5RtM3K1beu
wAcAiPzgDwg7Mm6YrDYlbxkQp7H+wy4xnQvRNCJetPvHsPGxUXASheRYNOLWy/IZ
qlHa72YezvFsWzujOIj869BYynPctoUJzv1VeuJnra0bOMJtsx2EqPTl7+LgR13b
oiqvMV5s0TWSBIHYaYkgNqWUurTMCt8V+OqsPkZd+KjVcJhQ9BBATKnkaTgCCroj
pa+7VN2+ok4/gPwtCJNJRw/ENF4Cmiumna/UdSSTHslwnT/k1nZNdZrrfuL56nVD
Dc26Gs6/zUiD4/QY5qG0igGiJqQJZivRzRSDBaY7SoU=
`protect END_PROTECTED
