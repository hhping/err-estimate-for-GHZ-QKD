`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDghp4c/3I06EZsbEIdfqHM9fzyavIv9jC91idAMrpsoOQI5TYCPL3l9po2y10k9
2BjL8nCfHGFCLOW/A2/S+dgcRIo+wI+XzHVe6AWxRskt3KMx6/QAvY3i8Rqo6ngu
1TrDnWGTt8q3mZx/WTrgjfo4nF/fI1p1WFpbzlDh4bspjJftmXstm4bGWbNO4CRN
mtLZqQ7h83e4eOSWNJXYrYwUZkjuXAA0yemGj43ldUOIXCfPtAx6sJjvVDjtZvFi
YzgygvS2Ko0IMz9lh1ylibnyMryOTb8dVCoLPLROXrGvXT27BHqKbgpaZsCctB+F
u0T2NyUTPrx1UDk0rQbSAeADTWVBp1cprnt3vw+Lv8xFUfp72t8UzBj15IBByl0/
4h5wGc0NZWa6FCM4tmXP6bwXlV+ka5gwwvQ6VMjzZ0yxNZaUzg0WYF3s7t2fCBfS
a6mEn5vcBri1CCv557/6gHdhqKwN5ydJMUnAzVmloT4YGedAjYqOxYJyzz/n+V28
HZe7Ci83tx6uxYo265TiiSlPMSfV6T0pyZwOVLcREPU51ELik1RD+E2q/GhdtO+3
1I0mPhV1kLt4DpysIBmahuDI+Ml6+MUMg6dqJ/ulJTsnR9B1FmoySZtb5+7HKNb6
LXnje7SlHJnMIrbgwwttrvbYQgZWRoFzuSaRgku5SSPfO0n8L1GTA4JBzVdvuzcj
afI+tnzQ5pCPNVU6+yjp3y1rWc5WWMYnj0yyGzQsMluhwyLZjNrJlOLAc5MGi0uV
pwJ83qSb2hLASO9mp8B7AiVGRqbwjjxBtwz64UXXyxLSiph8r4yxr7rm981YWtZ4
zINIVqukpBFjdHMaxi7PTA==
`protect END_PROTECTED
