`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftGDxBGf/EBiK8dNicrp+ViRtqMwlRywJSnUeyf/b2Y5EKqkcyeBEIMcODZ5z+GZ
xLfr7V+HcyihbfrqhWOZFh5IKKta/QfMUmvKkPqQTiW0Dhn9pDc8RurWbAAoCnVZ
pNzWO92z9em93CBNGbsUg647tSkBhMwtHU57fWNI6x7usCvQiSxh8K3UedxWRNJp
+/SUE0VWPYI8SorSwPTdnoq4vV/AOqdaGLtMXvotlDN+lFvhTGU7cuUasBrs+/sy
G/86o6BWQ9WtozE6e5jQLOv7SdgFS+LrVr0kNEHVl09+XkhjUraSQoIfYfxuJTLP
S7eg9LPNZNzkVZGWpSgnb++xkg6eFDcbEOG/i5qWFCM1cn7P/jfFsPgbyhhUrL53
Vr61DX1v7tJs22ASNuG52pftsD03gbgDGnYaOVYHL5GNuwt38jBVcYFGjLWz1qXu
ivCkpw/UBpBq1JS2zK13MBt5u0SDWn+wXS/rLKf2wkyRXp/WjGu5sXyxFPwmEffJ
sHSfpvJoffv58eT/iJCvqnx7Xx2kzxYE7JE/Bcvg7EjoHI7umYkfVM3HrI7CjWhv
QLT8pjRHai5cBQRKhjfqMzUQptI0/Ct7WoRO0w3eF1G09gPsJcuj/ouCtMu3X5/x
MZpy6eoKhzjDVHXJpiNb7yjotSSCasKH8nhZLoBuGQlok+u7atcZL1+oEPOHWKkg
ZOtB4AFKyM0iuD4sKiJf5U2/gp9m3UhSFRk+WmxmAzJxQsRAr6BSyGW7tMb0ZT+c
UM8lBmbzy/CDNJjKouFv7YEKgUI4zj9il+lHHiyimKggqzG6BxV1LNY82bvSWBe/
q17QJgOBcC4N+azhPftxdcquyvlUWgU7+5CwAb2ezGb/6WniVb/nyvhzIQXJ3VVM
I3eOMBGQvp4lBUHqedmXg8XiDJbNZ6c+5RA9jxUKkQxij4WvWz/BqAQkeiwyoEye
+svwNR3kKGDNdS76+bVCwpemRM3ZMGgT2awJlgtgObAeE4SrVitDwwhX/Mjp8tGP
W2354Me4l0hTk7734jRm7Q==
`protect END_PROTECTED
