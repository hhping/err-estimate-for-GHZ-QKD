`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6W2ppxvIzIu+Iq0S3+YB9O/v7KE2oWe87UrrVdAJElboBlYpQ57PwHel2HKoJJ0C
LpZG36FuGDM6r4xv5mupWyHTbdwwM+c6ebPIAFlmQA0crELC2YldStZd1O5EoLcc
+pr2q8SU3JnBC2X0d8W4rjf9yynmpleObyLNtG3XdpuH5AE4iDL1yLbqR4UirDU+
P9oVOHblHmAzNEJUVs2czrYS5LsQgd28Mv1dSb6l5gEMDnKudxmL0kwuYYU1p/03
CMwL1K4JKzpoFYe2nOn81D91jtLB1pn3gEqPXw/c7VBLdHVkdzvkrpthhy6XzUfd
Szptbub6fy0Vt6ziZix2Ilv2ygNSNbAAglUneCbAZCAGUOrPdREM1S9sIrBFFt4g
y3cXsBod2oCYuC5v7lbnDiX1g+X+1N9uF8TjnesfVHbCEaaUR2BskD83cBMuf8M0
XTbV8ijAWMJkMouXa9AUGEKu95WB2n2JKx9WxDytpbtBFLzTm/yG3uHzh58DvOL4
QmCS7sc+2pndvcxmcxZssMhAKZm1c3NRKYnqWJ9Cg+5uNPs/1Im3gEJkeCFN054T
8I9WmxSVtejYLee2doL3VD2uI47RorzQ7n64dKCwcAZJ/1t5FUo76E9yG3BD5oCd
`protect END_PROTECTED
