`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftPdd0BXO8C1ww/ugDPR3hiCgu0ekUWJtl+IHpny4WLL0jWAwyKN7pIkxBkCYyEl
pIrNQ40YpFyUAtKlyGbIxewfZ9vyiyPuXnzWR8XZm5DKhpbQleMhUD9Q0ypfEpqs
jSmIkpZ1J05PfL+n+8aBcupT4vEWEV3JLq62GGdDPSOBbmYRoDqek9r21M7WdiZV
ONMDOCjB4OTk3sEpfE4z2EBk5YxaKOCdb9dNkbSE6ZcJ8Owa8M3+3ee3j/g5m4JD
4f8Sk+shIaVBLXkyfvPLdI/Vaz1NnAs5OcN7swPUA6oHxOkRQDEgOSnVS7h0wT+L
3zhz4q0pGm/vEClNSq9Lc41kKaHez5cSbA2t7HAqja18DAylnKmNICM++Qtn1oYC
LAZPWaHw5NJa8Z569LgsRe/PjIOHOtTz1IOk79wCJ2ot9k+jlzLswGRUsJvQKSIj
sCUelGgUw8JAzxSs/PIRK6SZ9wAumwr3t3WlPBRfiUVAxPpKV6OeU2u2grjSF1NY
pJoMrA9m+PuwKJ6H62F64rBGVjcWhoM2NuufTdDYoNtCDPhqPeyig0o7rQtSzQMw
aJnoIlXFCVB2AkPL9at8kWcG8eG1neX/PfWlHa1tGR4MmOKrbems1fPPtFbzDZ8a
xmTPr7ZK+4otl0sCq1AELHxZDVaDUswOeFTO0JPBne5PCUcpmPz4UoLzZ1BVFldK
5+icAfc8tJcMyKQ9vBXrv6M9YZ/LKQwRbs1w92JP6SBB57xI9eiVxaNBo/fTEdGw
i25//thkQvtveX1o2cILytdSH+vDtzDqtPG1ee79ZeDjH4nMII4gDuD9K3NnuUPA
w1f6eC8OVxqworsUYTpuhyOMXWGOtLM3/2isZ9/JZ7amGY6y2x6qrzw6JjtO4AMt
M7JHUi1b/U7NGCNTbcfvV0iOaHtB78WEjDiFfRRgoOkWB/ait8ABTXovojydP9TN
Y55AzvEDf9fE+5eUDtrPm4iyYscCqurxgWnx7Teh7nsvL/27I/8XvwkkpKe4GnsW
TbaORj+7ouOFr9vfENVi+d9IQW8CqbRLCQUbzesWlHnfeeBJJcK8ekerbOwEMSdY
L0sQXV2yZLpTAoaayNHRB8CcNvsXhEt/+M795pAGARTl+mfsHGJRYRPYV0o+5xJR
`protect END_PROTECTED
