`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLjNKVTkaVMQ80wiIw8DnY+3WEi5bgVZyWFgYLTJ+BzeBpNWvJ9khKE5yu3+FF5W
yFFyGCb2NTxHD/OrVQZ48izrR94pOgwDohJPS3QAwowxd/2Oqrp2QPSZsp682vzl
hJYY8+a6iCR3ihTwkVTKZmZDitp6SU32EUVdxGtkSCFM1HrrGqWIuqjJt1Mt5JlB
UXsm0j2Yos5MWK8YVMIOW6MFSfZAsKiVFxHnA80r4FbJqzFn2uTQ91gzbRUo2sCk
AThhef0zrSveOu8VoolF/EwETW2OIJd/B3zvOAXn1Mm7U0f1xCxw6c81+5uDnwC2
FaiPooaozPddYyVn3IueyG+epCgFSXAlTX1u5ShTQ06RfrBYQ0nLWwqTq7/zATC8
`protect END_PROTECTED
