`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbs4mAV4Z5o/h5EQneU2gxaUDlfb06cGbN4CI9BGVuPDc+qaZRl6L0uxp6PDEuuR
XGoyPmgbPHYU8LocsoOwu/HmGJw1nG3FkBpXdHTr3YVsHa/z3yuCyIExzZkol9/C
8Z3AoYlgTp0nDhfLznq9bz0HK78mf0kz9e8jAh6xrNmX1Jxk5EKQnTe+0lNd5r7H
TYZvI4vSoJwg5u0auphHM2oLR1V2xpjU9cJmzH62TWgb2PerLAIiOK9P/bWir6Hr
7ETyGc8yD10siGisFxbuIQf6mXw0qe6cnp1xSEKnmtEJ896vvqrQknihFmreVV6S
8FNzsrDrMQTA4mBANDcuqPuPIOdzrU2H/Bk1vxKAZzDsU/wfDe542pg1jOXFURNW
ZmnqXcxoDvNhNrPR5h7F+VcXYkhNw32q9XOdYsG48zkIFntY6IkjtnZGYyOgu54p
R788xRpJB/XaOFFTVCGuT7HXKIoIOB2o0WF3Ss47bYKoTn+jAbBnsSfSw6afEklx
eUTx+KYGWOOjnsPxuULI2TXxOkTSpYIEuFwYVD3oWSx7mJLerj9SBQuAmZWwgklT
g6k5ddv1R/+x+PslIemCzAVsodBzXp0DoGHUN1ZWgKQauiV+s9VY++ww5b+kA7Sc
cExZ0EI3As+LC4RFuvf06srUjsTFJtsweONK2WmUwyRBZqbJzACxvEYosWxgE8EO
1ZfZkl1t+fUDi6WijH3dopov9XO2J2PavAnXRXrX9KTvqqHCnNGcIIpg94bRsp6H
vQ+sAVfmHKDr9rr3AXnwpwu49w0Pbgd1H2cE31NztAbS/OQl0QkzSQAPSokm2H7f
lwVeBWXFjfIhfVc4zTpYiIHKMKE2hoHE3/ncCY6C6QYBmkITzQcEpyF5OSh6ar7h
9fQGEW4ITQP7Xc6KFSoyzv6tYJKAnf3OLBkDaxOllJ3ACiIfABlljLOUo2VOfE6M
xxEg0k0AvzBhow0iDhF9VxKVFf5DnTntjuDduyljVWqChyuC0gDputGfHTfcnFt2
SFsWmC6NKTnLuq0j9+CfHFY0G5Mr7pAj/eHbgfnxJox2yZ9Ew7Ie8XaOJNg6uFES
DgSDI/u2/Vhu+DgQm7DlICumBv+wIajfLqg0wF7cYo9xUdeuE7YLeXyoWMC9J4de
gS7aEsM+XAvUNsQ6NKvjCzmCVyqke02VtYPsJVKodzsRet67ibw6YHFa7tn6WsiD
cAzEp0rhPTTS4gAa3WcWfFaZUXJeiG9qBYnRnqZnrRgP/0gyiMvkmDD8zb6xPngX
zpHHfy4VXGJxCpaXDtGFMdJZGmqcc359TEsNKQWbzkU=
`protect END_PROTECTED
