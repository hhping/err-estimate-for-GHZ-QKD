`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eEhugT5FNCbG9iChCdnBDcwTYV27fhbjiQw5Z51V5X9WJlLPlv5KJ4coTIxqUcwl
I2DFDthvnhwXZxJnJGBuYXmoFDJXo7L5oGwr7CQmdMoiSe+L2HtSHOv/etELLImp
LLxesE04bFd6RhUmMMXNwtBeNbjShuMLuNn5ZbaPq0UbiJd/X16S75by+aUUj4yJ
nwfiMvyonah9FaGIZ5yryeY3sg3ZraII0EaN/ZrP6TeefDa1zEgnZ2Xkw5wcMGa0
+5ApZMoZ15ji5aX7cPGyc1iznnD4YuENqs+Mx7vzzDjmNjBhBnJOtyphsHcEw1fq
CYRGqb5JeA624Joe/p832l8MK10GUtZvBkgQi5WuXemAjhAH4RLvnq0aHlYFo2R7
7yXa797r5/fp43hawu3ZAOgqNcNV8qFrZkngygIxtC25RU0hi93Bmx3CEQM4S67h
vdC4TwCWJ8re3aD98VjfMfH1rdzegpgIg221s5Zw4byMkGpSOoQ1eTK2tfHAfRQO
cplUa/Dk68FhrxTqtrsPfSYQgM/VnIIjgTzy36EnOlM/bDhLFzVihSg398aHh1vn
exZLqh13UMmAcPjd9KBBkY9esxicsDlZ7Txc+MLnGP74ku6jYa56fhCJ3/5To+CL
7MNsEGr4KRbdM/c/2kDU+BSx6h1hImIIZmAZwqcDJc4oB1aYDteF5MzMi9LwInRe
4bYz3FuUm9oW99UxxAF/P8dnqucY+/3n1X+l3tFGxHntM5L8Hi1bg7n+m91BwkHf
bh29LZN89xXGJU4RxSZ0m/IgwMiHgiSK5wQ9hQOiPxeK2Of7S/4TvIYyI+rKtR8U
uPP8ej1R9nvC+pqVioiEE+b/KZ2JACjaUnrMlDYDJyDbqeZ2LTBYh34oAm/L2o3S
lmrS5XFt1h7qsfiiYxdAQG4XKaS+KGgIV76PVjtluih4H6uXskAaGemJHQfrtPKE
cQlDZs2VaJ6mde9PllIWT1c4wleFrzj2RtVNfrnb9qk=
`protect END_PROTECTED
