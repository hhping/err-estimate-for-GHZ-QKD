`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zexg7I39Z99v+qcfd9VcbzaIWB6Hpe8NuvehL++A7SmYwI/V4xLgLnNITdX03ggL
Ro3M7NE/OQqBkKOLu0VwLKb43kJQcwpxzVXWSRV8Y1GKC1ijVeL9glbcWLau2Lmq
0Y8EK3BLWVRdg9jkomzJCavRxNnN5mJRTgarqAs0tKQ3erG20PM9108sfnw0qi4h
TO2mVV+3csIOcuC0c6TqVI03MhQYvx3sj2yZJhu67I7aFft5xMh+Pnbs3GZiHzhW
3svu4Si3KjndJPS5/bonSvuse3iINjAaJpR09BXCkmm3S/OFZxs2COvBN6M9w0Cd
RRSn8upAMT+FRH+mNF+nJe6N7CIHYMzhxcooctIBF2WqLiM2IwxzPeTMmP6IQ5ge
G67eGVIZqoW2oLQJt6xwKX97giwLuh1shk+aF0ws1Vio++n9REG1BgWcOQAXu6vg
iN7CBBxZzY08NmxJzy3WzbrL0gUwtdbLwfrAS5tIwtz6Km1xiVHMzaR/YOAPonxW
qMPj79lfjtmQG/4BVzd/x+9fYON1etE13C52j1ejP+PM9IN0MEy6iHZTI7qKIYwr
rlbWvIxUSqhC3eTB+eb+nG1mG7y0hhrcl8r9GMsFUpApbGwM3la+PolZOeaK+oFU
`protect END_PROTECTED
