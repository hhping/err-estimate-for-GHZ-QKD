`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ft3LDlX4g2Zi8xt7xQ5TU/PzQN12+/REMJXs6nxkouDAz00muSJ77s3hdgJO3Gd/
etLpgSmyfDkqT+FTFi7pNlk9i3IE69H8bzjYnrdRBFJJHvXMssZygKdueYBvPTk8
NAwce90/DtnrR0zeprvBDs6+Z/3hHb3UADsXkStHUGi1mkRc5NGH1C4bEw4o7Q0+
Qxx0WzNt8l42ODFENjVX3EttqpClDqYZer7wce9j+V5m1hnsqjK3EbiXsbMGn1qn
XhwYwSe0laLtqc9v7jR/uMoDMoqyU94Po1rZuLDfBV3R4IybIk4YSr51XtYaPZ27
G0m8dP0pVvAmxq1HMW5yvjoRAWe3xTziltlSqIry9EJ1Q6giQkJOqicWKHDchOD/
Tob/4LHJ4DTDOzepPW/MI99P5EEQxkIBk2j5pUhw4m+BV7fuIVSpgN7PCgVduvmY
MzuwpuGXRQvHkCMRrSiisXA0NFb6P3p5zvJaR0GZLChganXnGJXRRmIjZn0UBs9p
EohLDzMTEQ+/Zxt9LJbYuCXGYzW5aLnZ4s3/72Vh+MEADWRx8+OJ9hI8d3ObEeAJ
hG6oCMU6u9a5smJi5PqQ+XYywXaGpZsSX5zDU30sMpKmW8VTqaJnLXwuNIBZf8Yi
dSKkPVqNsxOi1Q/dYLKRGQoPMMBbrvB8DzBJg02aj4UM1ovKCzXoqWSE1sp1Fhx+
rmizfqqhKBGytM+lVJNAlvhrLgIIE+kueIcQ5vjwGAmrzx96IXUuYE8nQ6GVhEvM
ghU7OqqlVmGFJUUkca22xGuH9zEyjJZjvAX1ozhbTlc=
`protect END_PROTECTED
