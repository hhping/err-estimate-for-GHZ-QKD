`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mPizshUrKhYZzkQfeZFGjnOaAEGI2KojJTAKVRLlkkgQJmwbLIzmbo5lWUM41gz
DnYUUxjuXfnkwhH8PfSKiGmSHiIs643+m0BKFg4pd+NaJfVtz2looINJ55I5ebCC
qrYmg/QpfBWLTQupwfWL2x5agg9nGCx4CP0XXFjTPkz0KDiBsCNwyARyc6sDZwRi
3SgrcfdQiSqpUlzigphkWjUqL2fhsKxb6mTFkLl+ZccBDJWgDLlGQqrwul5wigyv
gqCJJGpUmuS6gCBTFxnSmY+66O2oPz63nHSfIkvV6qQ=
`protect END_PROTECTED
