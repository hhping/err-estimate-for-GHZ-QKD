`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GaEVailzPNB0K7Es9guSp+HPLU5g7hpjShXP91kGUBMx4zEqaBnxGCKeJiPJQEcP
Pvyi0KTS0qg1SuD/WLwKPKmBxvZdC1F6jU3XOroCemJKjsN1pwaJlWATuEYqhx2H
3f+g2EzPVL/5YQvZ/07ghRGTgeqDWcrSyEunQqcmA5saIxXnBAi24q6JkFjiQxz8
IewqXXbr8PrWlb/VrAnEXX5+9UI1mnHO4hiujtkFSAmDgCamm3Qcxisb0mEh+J19
sil9nME/uU8txYkfxa/4oomxI7khgS8RabuClTzosclTHreWrWQMTR2/Cu/NyzFK
NIbuWQHI0+fBtyxOkBSc9HVAkpsQhsfmgvNAtSkWRc13CONZhY6cBKw9fwDEYf0z
lqIAg3x9b4BRTDWQ4kseF5EsXVM0+rV6npezshgXe07uVSdriqgulNxLN2ih+6dD
+9w/FwjQSpgKEl5vSsr2DDDs5bpIygFzNZNwSRIvDCIqjfo+aLF+i06FRuw2i7Nm
TWj4goxhiH0Cld/LCB/TkEV1xUa1bU1RUIjGlMdTIqhVomqpml9ZMFARftOZDnJk
IjCNx7EtESqbvxDt+SVxaWIkSNP8Tfbn+0SLvtQrGhcTOT0Ec3wygN9ZKfPW9fUJ
Ww+HW/NSB7rXbqPIaLerkch6lOFQ4r4ZrR2YYvd+ggqp1ZMKvixHjA5Ld8LunFQt
SQU48SGtvrwzXYt/DkjbqFU/l8PgwjlntSAcOqGFQ9Yj/SLqQHhp7ffyhfw0fusg
vzPguncqSiMcduFcFZGoFU59RCC6gigeZA7ElaZyVfcOWZL4sEVoQsYuBRs8HwF/
INTUD+QNcRDqQ+IkN+a9D4JcGYNIj5QOPYaH0GmobhFtPFAnYrtSE4mCQ7N0fIDE
PXqPTm/kguPWO9nlllkdxonz4i3rp7kULUR03M4zk+NKozTiAxkZQ6tZ6joiuXtj
6QaXBECwlvsNgjJsX7DVORJ1EP8ee2gvIvKjfQjgvT0gLTD9FxJIpx+MBEck4V21
cSPgeTMu0L1nPg0M1SlLwffHMyddLT4n3P8nkj6FlZ1EcgEuXBWVHArdY8jskcZ+
rxKCTZVwEf09vohADbATzVXnFdjQWf+IPs/Hrs5FXo+wfACfxGu9Ug1tfGzdbKbg
qmxQyzy1jxdU72/bF0O1FAy6+4nOFdwC6WnKMYtRT48zRL5cezGPgCEKtdiD0jgH
f8gB94/enUd3FA4vTudNq0/Cv0PCUQQ9DlImEwwk/+I=
`protect END_PROTECTED
