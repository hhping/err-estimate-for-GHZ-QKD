`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvxbqbhOfdnMDZUMUau5mR9WY5CvQKpBGde2u/BJ3t9/JMd8oB16DjEqu8EvZfH9
/it5wjOpoJFvXeJa4SFtjVPUMXDQY+q1fHhaSkEX5ZNwZVj1p94WP9md8xTQ4BQ8
AIoJYmrQ0KLoXqnwNm/IxKKPvpurq+RVTq91g9ajUmRmpTtyFHcwAWi1ZjxPWTnO
xXkQC7H3OfM2RGtAHm1qW1A2y04LNpHI8xXEvxObaqDudWloLIFnrZ6h+MSg2g7H
oy6AUIJWKnUs2cVwo8WrR+S/jxIt/CXw6vlyKD+s9y7i87Vm5kl6quh9u8X52APk
bweMCLWYxTxbLaoBak2v+0MDkAp5Vk7ud2ZNZbKtc9HkfrPosVGTXVNLYn6G6xWW
QwpQDaZWmz3njHJLBgFycQxTnJpoAK9Q6snnwQ8zc6aiH1EWEkEPN1S6Ss3DDQq9
JPYIhxNsPHA7Z/VBwOEg5Ff6IYQC0kU2sAJikCBuuWNVGCFEA9BJJeq/0IVd7A7J
sd+ofS/2nfooABgD5il62EnKyFp2Obj/yIsSrlGvKbe5iNl+pMah1Bbzj3XHKbFV
YakaKlWRSJbyD+9mhKjQVv3fv2KVWJ0qMHKLxFAx10GfIU2As3/PP8k9z0qc1AK6
GiBvUf760HZb0W2WaYbMNM0iCr0/np9RzX127NatRDD/U25mAojgaEay5BGR7x2b
yA7Ep0w8bDHSnrfclH39UItgjJEF6fg05os4n0XyFMonWzdOrzXPEDtQixiBP44C
13RDlZ3tJXrFAi/u8j/XKOXsofPosFP1uoquPvvsc+P2N8RK+kwm/EHiiIxV9Whv
ojR8btx+vPFBrv4MBPB2QEvxEGLbCwVOYnx/6S7/4mCAC1pPrj03S3hpgDSClyYG
zdN1Wn7tERP8Z6OJTvbhL5Lw8X3XTujlqZXdcW1drGqUosNwVilf2mHKuKWXDV8C
BSgQgPcW9CPp3ErsR7kqZpCwlMvV4JECcdcVgI+/2LU4qUjX4tgkihjf19p8Ym/R
FJwtqCmbc0BYWXjILon9Hfi+deAgGVbHeC3s+UoBqG6C/picH2oXJt9wVQ3VqwMh
KgtvC9lCucSefRJyw9UT1P6iGCmsTIuLUhpZOHo96fx1JF8SlXgPigGHQqJzdoOI
+nft9zWeUCeLOp2opq8HB5Yp5S2WtGZvclB20xMJUK6lz4fIIcyW+Rw6FxqCUrfV
nOF2y1SdSt5sysmA1z+2LCp8NbVVRVVOvPB4yOS4PtahObtaMRkhe9Wta+O+MYeU
d7JhHIifKene6yNaPuE14vnkEzAbNLqURHh3Yd2RIpGXJVbMTU47Z5sSX7sdKuTO
Z9cm5zK6XIiQ/u4Y+KSYdU/Uvn/e5m5/b74OStObSwpsxISE0hoSY6nvTYBxgH26
vuocdEhixU4OcrZ9jaTyZgstgDhk5DVZaILqlrdZBjRLfwCRwV14diveUy3yeBEr
9Vbg4qlkRv9rbf5+wys3MtAEyaw0Q3L9vcLuT1p4TqO4atzsByxcDirGlrVbidXk
0wMr0Q1QqShKJFnP2/EqgiqCoiJoxTHj930zTsyFvx+4CAmJbSvHJePZwVnP5S8L
aIIo2eT+OD4PjKZcCIjnf7ZdMPNZ2TvGaGIMAU/Roud8e4udd7QMNEqB2qad/OAo
yzu3iwKl11fiqux/Nkw6KtUkXyNhAtmfUarYg2Ie8JWoH2yw8Ch6wni/v6G1dssi
r21d4IC519r6qa7v3k1DQiSCoWEl2y7L7ytiwUBzT7/qf48gDF3wMkTObXEToZi0
rjUCwR+EfiGTGBbDIYMR33RpXPY0vpvj40bBUXJ3+V8m7JJ3ia002IqLoXUUKyMf
L8Xb3cFflJFDsTGrHl6v03uVDjzINNoreW8qxmlVbkcAz+6VJJFwdGifO6TTEB/5
8TJ4/YbkX2HJuuqdkF33Fd+gbWqdoHvMRMMCVflqTzsLTTiFHwgNz4/8/ofI8ITr
4DXvlTKkqq+6u8MGuQaHuRh2HdD2i8D3yvO+Oxtg1IkmxeqRTHWYHE60KPWxjvrP
WBfQuTkuy22fQf8ulqz3gEKpI7H/9rwfwdnff2aQsWeDxt++DzdbAguDRQtw7Mzq
5QbNib/c9+nrLS5XPYke2gXgiHnrhEwVX5mcQLZqn2erDv//CZvtlsHBOMXV0y3V
oThJtcP3TJVb1CoxODj+JhW6sEhXtxYiJF9g5HoK5D8JDuPeX+QlckIHUSEDvgYN
9u0jF41CVjmeJjvobIxWG9tKsFDwoQiEFbfPrTh2EA32McGSFJkxqg6duTQkFtu2
zJJ9ogHba97UgZHxRnXMbael2IfU3t34OUMNbMyKJiLoTsrMgymWamA/A+goxxqV
6rxEyO4phyGrAPKs8awqIg/ek0qNYjjM/0/S5+zyK/evxLq+A5E0Yjey/B5Gx7q2
IPC9KDRNmzVBcOu0jZVZNB+qrd1cJTMLiWrOgGpWMJNezSHkpjzMsx+tCQm4qoiD
UBw/P9TQVtkiZg+ecd3F0/FoEN5PQbT9znuCntES5N2ZN7xcdvmYFxqlu+kAvCyY
ZswJsM3n1O544KEHo+JVx4Qy1Q3PLHIe2Y/BdyVktRkPd9B5R+o4iLYaO27urnPG
/cMFnFCoD3baMeUT5daav9U0+e0UAVU4nVF04PJGhdjdkd4jnk1AOgAUGXCdx5U0
i7Gu9pwTGuW+pRVxckKxb8kf5N5FXmKROMxEhS8VZVVxIepFVIW2RluEff1zWK3z
fB8ZlkWuvnnMksab6mUu8jspSscuvFOCf0ceHNhoedw0dlEZUMFw1lEf+YMA/ODk
+KVxrijODjBUwelUiqt1e0J1WOtgBe5tugjmLIUT0f5kJNOykDTNcQDk+H2ylPjv
Icplb/ThwBmpBdT3ObM7g+NZtW4+YI1jqI4QsFawFrq278Uo2uCeP6H4hF5gSeUp
32T4AWcob9lUhnp3lXnWOT3TbUJqpaB7COYHQj3909MhdVwj3H1kgN2VbTbF6JFw
CPvjvBCS5eVU9PavoDhxZ/gibfZDEr6wHmS7zrbe36CrhKf+Y8YOxhAyHJ2gpKO9
gC5L0AIs5Q0pd8X7V0z0m2cEMeTg2PBIe8ocv1oZ+uMBoA7XIrpAd1H3y+sSlijm
UTY6/2tbOAdm24TILNgMhZSr0au0Vh4nMt8mFrSoVWVZ3/6SiWdWZS6z+flqNmmF
qndzhC3ngBM8g686/z3Se6YXxBeUtKjK9P+vlzbK8KQcVKzRNioi6qwiOkPKzZwx
EFJdnWuHjXReb+Nx6vwtKHP8kHhyCyUD9A1YwMVzIo75bEqyiPVCufMAnjiU4+MX
kXQyIrAsF1uE9y8rTOEJweyBK4AN9fVjp/09mc6EEfNlYjFP3R7VT6sCAv4nECiH
+IUAVdmn+nHmgBDrsIObQv8Sqj9fFhyIPlmL0pduOMVMtMo12xppORKBBxpupLve
9mMZQFQQ0EL3+1X4rzYOFNpoYKVMBFYJL/oofRbhVJzJua5vOHw63HBAXVGAHhVJ
ZvZdcxT15qZjuGwyOOdTveyaZHKfHEtd8tQrojKSKmdJJiXFFSH1QCxTB4wUVZxO
SyxB681v0Vrh9V2QhIABEUvDqvF4C8eDsaoJaIyKFVK65NThCzUdlxPPd0qS2hOa
gdbq09bykZDZexX2L+adaHxXDxtNPin6uciESEAd3HVR0m61daYrxoJ9hOIKEYuS
x8kZaAjo1LfPgbax6PhTjaqp3GrBc+xc+/OQpmi9e41dqrHWARn7zHmh/boxKBp/
f7xmSHsygzEygHHY0WlCKD1YCVepuBFfMKSk/qPFrAzqu+aBASItJQ1ARUU8L59X
6wGidVvMMbV5HkN++OxP8raymOe4kVLQcXAUsP1XEZBk8jTrFLXe0lnqiSlnZJiS
q1lMHpfhvvOz6WzmP3HJOIWOECQ7ybG2vQVLpHJD2v4iS33p2XgC3RYXyZwYHKLD
3syivaEs23gEccMOZ1McmqYGqAchKiwdCHSSeE5DQNhj8mzZolXaLIkVI/iueyOi
V7nwqnWEt3/cX1ttAHN5YmuLy7jXx3e3WMogxqbjajkm3KAUEVCLD0RLleQpr03S
YS48e1O5aOFoUfzhsbRn7rlTeVGQieVM6APHhWkwQwNnEA6s6uWT2fYss2cWTM3V
eJusQ+1Miaf2T/3Mn1pfxvxUlwRUibFgv2S0jt/gmtdI0+Hfe/4eQRrPzzjew+nw
2jnJNYK3tvMBF8WT+VWXVD7APX0bXzosrNVXsPkOBS5/OW3tJpllAyoiC26iSsaq
/UkAua9u6TVkDrf46kBkcafGzic9wHgrJ+zl/95BEf7qkXc+uS51C7lxF4ZepNSG
DYKxUMCCuyAYLSrtCpfpMY2Kk0PY39sfK9m8n8JoDAgSJe2TF4QfHI5Z/ZRjZ7wD
RKzV+MmzSzZLpmfRhyXO9hiwP7WMgqcWedIILHqr4GayQxvrgTt9j7QktJ0BL5Xv
wp+st3Zjf+HQ/+7moepdWs5tO4MtvRkLWpuzo9p/Ne/ljga2c55J+2C14h625WtP
PcEj1SCu3FC4qLFhyOMeGzgEipcbo1caD1Tw0NsChiRH9FPikYAJDmlKG3vPdKli
zajirnLIF0YfGLLE/AJ80e35W94taKCN0b9wiOCtZgoXH9KdWS1LgB6hrbbWx70y
78j8cYl2IDxrt+rEh3rljATM6KP6ZSt/rQs1iwxeh2jWQoi1LuFTGR1RdZOLbIqQ
Ih3gD2xtnjpXkQYb8ZN/ADGF+Z5A8hJ0FnFLgOwCDfk84RVfmmgaj1WiEQhLJJ53
x0RPVvToaAuwquYvjx+pADtlL0RkviqhGboGsU1zJW/nUowRWDcsj51vgqGxKhKq
SYDOk/90o36mc+7BWeHL2bFEBCJudIJx2Mjd604rGknwNYtJx+w3Qw2GI71P3N12
VL9tzQL1JJWkKtuLgnxZLGZd59EVkyGhyDMwoBLNWFqBmfbhtJXuAiTO7QrH6u6V
eJy7Nn23C2RMIGmmEMPs8XuzpdSDeE72lpJQyuo4zZ+77E6qdSiUn0bCaPX9fHY7
s5LVuid5LIJscLLRrkYkr5N6csDLkir3LTQx9VyyuwhGsrwHrQkWp4rMN+2rmdzf
UGuPNixB3Vqn+m3idv54m/I2l17WKsk4UR5AwjCZyGaM25ZreNS8fMo2BcBgwpWX
z5x53hHqC3rWg2csBtk5qBVshRD27m1mS+0aOo2Jm9ELcu/U36lVFAcQk6k3nCvG
BmsrnhTiNCfZpeaO7GaHxx+q5RTV+/osQccGb0/3hD18ObemiTbFFmgNDktoTtcQ
1niVvVIAK4/CqYVmw8LUspzuvUiW7aPUSa1mcMREz3eNAaJsXZEAkkYtSmEdk7T5
/VDugA3boB+vOygQSn1P7T935VeNYnAHfLtGlX5yTJC2pf0ZdM8qKS5yI/kzS+hX
M79f7baqv0XK3onV7UBaNyikbusJ+6lFuP/KyrBRfmo=
`protect END_PROTECTED
