`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DsNnkQ42cAjjwI3H/Vky68bnFwuFuPl+RCaDdf42EAQV6i3kkx5UfYtp+gYonEQ1
u9gKqBN0FszOmjJdtvzXgjnkEztrz/C6Pgwm2AeNkEWIiuCMopqeOFUo7zhIudIL
t5JYuuNad7U+jsQooJWsh2Z1l5CktDU79sfi5i93GjZWwmPRnKyzNQrjvKl8PJkT
SFAGTnYn2sIDqRXhm9JUs5e2W8DVn+QpUHQKaQbBxNJdDrzk56sZ7C3oCqDXYGsg
a9qO4p+aOdoOSlmDHpbxNX7HN9D64CS+P9hNmLCzAg56tqjfp7kE7qvC5lfswVaz
YaPm0AASWEdOUDT3/5iSQwfVc6aLU5yw6aegrUFILa9Vab5BiVmbInhOETQkv3Gx
5quW80ntg3dgVqO9V81VdifvmW/ZkL28LILN+p9ohoQrcYlbwru1TWF5dGvREgoG
N2XjQlEM8S0/Xnw+DWcsmiS8/HaS+RSqKIIe24F5X//VOXuUR4Z0b/o0uERw5F/I
Rh7wWc1GET4cyWl0fq44NkszQCaWZyvrEEoozMnqQjPxNciyEcsYfp9pl+SzOWCa
Rr4bN9BtcwYB5yzypSp28SnuILsK6nyZvatAlwrDZARN0eyJ+G1abWlXIJ2M9ffu
hHd4DgrDGrbaHsEJ3YORo81yuKaYJM2h4JYw9tadqWEe5/FIghczg3g/OWhnWPG5
DocPa57MJ+IE1vamUeFWWcDchYUWIgujPGr5QELplgu4lLi7iYOf2ep8NDHFNiAF
0DnnUlftV19Ya0voBqOyGOpzyn/xtx4LF2b6AMamNAWh7ZkfkC737tqU7/4Vm4RO
QrYWOetiu2OS20zUJvKc0YCIERUSmC/YGGUvpHO0xoOL3yIjSEA1+4z9yciBao3P
9Zaqme5PDlqkh0zuZDLC1o7B0vedIgiJFNJy+2yz5IHBUAJCl3vfs3+WzRlnMcgM
uTlzv9NWzApVOObGIKb3cOViCi9VOwx8dz9aWCtiwZU+j7WWYapyKRD8B5Ockaqa
jmpP3126pfko23opVFbp9PvKL0RqQbH7Y7R5rOpqT7qkYMoWESLDLq/6+gZL3Une
NI5pU6DfIxkIVruIpHOhkY52/x9DlwpkNzP+RzufLhAngMLX3TK5Ro+f/ViP3XY9
zZZdAgTEkiGqrYI9Np3McCpkBXWtMZZ503OwkBUK7hu+HqIwHh8D2oheignwldku
V4aLg7tadOjUsCSyXcuYXP+rqTKwhzQlgTZayaRAo4DAAz6JLYA6WuywOr7kVHsE
I6bAQp7nxmI2sYP8bU01bSK1gnS/vOk5dVj9wzxcmq25rUJZVklfZA78a3clWcMJ
S0pYsQ+Ae2hQjxVwuUmjPH7wWAyWx/s8pmjGt11fJ78uKZyhh66knO8/yFFE35Ar
rHVYdp52uvvbpLmuhD9wiSY9URlKf2g9eGEIYfcEEVHTIYtVoeQeNqDlkOW8Dfrt
`protect END_PROTECTED
