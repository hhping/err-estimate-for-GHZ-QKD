`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TT99niITPdaGE2OZ8u883d/kWgrmzxFO6760T7jJGqEz6wrrl9kYm3bh/6b8WZvc
V6WwuNJLll2abu9gICYMZ7/WwBjLr+qQTYdl1DcMGmthPfT1NVwMcptJpZl8zBKo
gbI4i5eH+XCBAKLXhdu4RELNm0iZ6FlBA4V21bTWSDgiJMT9pLezXsKO3LwVFafJ
DDOvdF1Jh3cy65KVO+Dg3CL5E8hETZH2sLGs6ZSE4rngFuvtgokz+fQDP3C82gUD
yE8Vngu9QToZ6+tlTILx2RzLB30qFwyuU4xhSRt3dxiOYjZirKmgPMCEfY/Xe0cp
D8OTqDQ1u43YreUNPVH2m3BjDnxaF2OPKpEbGAn81sAIMCNUPJ5WGGh3m7kJNEuq
CAyx5Qn929zuwhP+G8We6FQOnRxE6eS9aYHG7t/UXTwJnRgHIJ0VZ0CTSn6FgQ0B
bp0BykiTu3OjI9bTh+t/lqAAeauGZ7q9i+l5W7GHHB5+PweZapOG1FYu86eoTAE4
1OpdklkjBq3BpRRBf4UJudq021TXdyEATnJObIewNYl8Na9spskDSGicNJ8Xeq1+
KG+5LoXtU0yLax2qXjLt2FkYAYEp4grFQ06YSrcIGPB+SB2cC1kF8WCQzmB7b1eF
`protect END_PROTECTED
