`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNGmK8DvHwo9j6QwiBt8pCYlMqBQdmT19mBHjY7HzUiUPZiQQHquv/1TnwUfqBM6
u+BELIn8O5rE7nobzvu+39J5WXB5UNXEKjMRbdqSgbI3yz1RwogeR1WC/VU/XaWc
4bqq3Wn40Rsv8yWWlgDmrHuVK2c+UZEMyI+G+TV6uOFf/YBEY9QRda29vAuYWOZL
rWbEUTQX/xI2rKz4PyLLpC5BudxF6b6gudm93woLNVBvRcZCjCeDSmnlvz3StS6+
t7GOijz42UP+Z3PG+awdAD3NsSLjLuldH/OoNa71mWEbv4p/+avSs7zzSuhieCYc
7uPHaCnmMkdyyETZG+FYfFllXFF2+fvp5qloIR6RGjb3a0Fi7rajFGIbygpjqvOY
EjkSI8cU1gpFlSTNYbyc9uAx1J3GxE6dqjxQqn77MnWyyYdffst1tUji5K9iz/aw
iuhk6amP3yKjDYT4Ykkb2Rt8zWyLuMTgTp1dSLyYufvwLBqJ7wMEmfULhR55DhVr
6Mn2ebQbEvfKOqzCswm3lA==
`protect END_PROTECTED
