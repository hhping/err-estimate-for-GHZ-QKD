`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1CMrEGQeECmDYhlucuyCE4NBBxJA2WzhYRrTT3vPR/nT2gq5j6h30FN9zA9SGXZ
Wk18im0lIoGCOSG+Q+cXwtvANFPI4vzkJdJoIMZn3eLCDqgif3pR7LBy84yZ8n9r
9QN4wzqUBgzrXyhLDuBFy9YyAYzw1LMY79bHH4Oem87JHRm8WRzbKa6fO8NLKldM
fhDkReX+OuCI+tQGT1nRawTcXOTPTjjewcHTTGbXQ2v3dwxAzKctT1PPxiRXouYi
UnPjwnUjSLyOVrU2FQR2QLrlC3ZHnlhwcIn7gPGD3hn+ri0sihUWCEQO/P5AcSO0
5NpiHLcmpYfedwAzZ4wVxmAZgWvo9h0MS2oH/03kSMjCz5tC4rVBuBiCBAOrz5gD
Ar0t/i+3WSuSXvBgiHc7M8l+PHIG0Sgl6JtY4Z7BIhVnexQMG3IHHsuAol89gTNM
irm0BeJi4mGnyzUoKCY6hg==
`protect END_PROTECTED
