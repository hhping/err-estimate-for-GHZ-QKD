`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+j5mrWWhMXjLDX5bFdAEgCqP1aSb2Y3rvZWIZqnLuH7Gu6cNK4zj020rJiMcPGkn
adMoT/jcwBVX3L1kWiew2aT1C0N45xSymtvC4JzF0QXMnXU8egSS3mO4M/lSbuPf
8evE3O+wVxsa5RvhhsrCXRG+UIv/V/OLh46bpDtNaMaBsL1FWvFuPQPKF84S3xNW
vKQ1//cg0Alj+BLAAvhsWTjBT8Hd3Wgj7Eqye7kYH5HAhU28Nwo8RnrS43LVOtYJ
xUmqPXH9t822x4oZzqs2KfBGilMucFXWBZI3XkxHNZoZBuqIdsLY4xY29Grimdi0
0GolCz8G39Lqrr5JK8EOigut9oXGa6MrkXF0orwzGxfEx+hyhvS6urD1q8O5SYk/
q0umoN4Enu90Z6UeFJnoKZiBvnXWTwmCT7YKUWtqe5pWXzrI1gE80Y7Vgx3ntuYw
Dv9UyoSaV7Rv50W0E9lruJOdCjLxKvmGbCdpKz4GmXUjdcFRn4RV/vPQ3Ji56qZw
lLEakTfP/j0k9f7ng4T9uLQ4n7WHMfYNMv/t1Zk7x1s46JXo2dyrNNpSR+3mBG4M
f4OQ5kQfEnbdCpgLkPZptj5GXjbsgPE4TBC4y3zceKcBSbn3TC7Actqy5XLwSZ8a
oGAu/IVljki24sfVmsLicRZADWy854o1XnfEU8A5r+OPVCx28Fpr6zegoNKGmvDR
ugPAN4m0gMUk8DWQ9cJq/yOQcOswviq+3vEE2X9CLN45qYGb3iC63+xxP7N0bI58
JuE1MnpVVSWiQO9DEJn8QuQS4cDC7siUJZ0/RkVmsJSQhlLsCnfDFmm5/0ciy/fs
mQLjyjfLf/s6T6q8Qnbsap3VHyAymsawoGk1OGq1NbtlLf2pKlK0cjcHMgaZk/Vn
bkg5O9nqcGR/Zl5GZEyZgT5MmAXgTrLf9YACzowAXt4oK1sJhMrHI0eXgupxbVnP
CkL9JOAscCrAyxMpAvHo2gOAWF+gsUamJEQClVQUHbA0FBkH+MyqwyF0hpZ+7nRS
Xm1WSlOXXZgEO/PjR5D8U8IVXvr9Bdkt4RCMrLlSz4Jj9AlhCNc8tzjBwJyFYQI1
+EqCbUCPargWbpntRt2gWKG76lheObszU/gBr4jCXHBTBEuqgx6Bu3cr33oGJFCC
Abjk0MhSPpNtGIZ8Rk1HQ7W6hqZWSvOsd1wLrDRAQgMPun5kFiTowY3xFT6Y6x+k
yt3kOPMolTqNxiFy5/Jk4R6mfCzhRnRM+5xtQxSK4As8HPQuKKfGQ8cvXetOCbgX
4PZZ7rpdrk/PLqh+8BiibkK3+uklgLnxXCtrWrUqOXlDy8pKY1It8rr14rA0rdZ7
KStT9xURUBkK4LUWPOo+SNmW+OST4UOXm9s4CIIxGooqigC7tExL1kmevlzstTSj
4sZiXIktg+NlxOfA/66wce5DWW7Vi7Qf1b+LOAF3My/eKO7U2Hy5IIf03m4HBouJ
WB2RHj/12CeP0O9ehZrjSMVk3o4SLfqee4ck2OtTdUHBGCJl7v7QGq6b4SH8EAnA
TThpV+huwNd/AhUn2N1/BtJWZHpjMUy3WeppU1eM0rbPO+poJ6DL7nPdY6ttCujF
pFgJ9njUoDNVPRUKleV1VdKJaHtSNh7/A+GvVWiOJlGX56tFFGZfXQjdZgkEJbxj
ad/GkGDqYmD0jBzYa1MVP/9Ja6hRirJWKKzT7WOBPaOiHZ82lVOEpNnqiiJ5Dpxw
DzFPxRGZb6EU/eJ8a3aYQgvZX5YIgN6Y/7y8H84z92l5nIb0/vzbJqgLwyyqAqui
3WjhYYP4smX18wS3ZUUNFWTFa8vqbt3uVjeVZhklo1lghFgJAxD9L1ohFigjmpou
gHL2+ZVZxU0eBKTZjdgBWD+m2Jk9Yoc/V5AGTTkiBk8X1iKLvEI/ptjOOexFpCc6
3UzbCIHlujvGKc1KEGPVI1sdOm4q+kncCfZELg0NiZLu3KAsXVIJVlq6//M6oLGz
LbWrCfxwqLa9kyysS53WhpU/5xrS/yt14OtLTVVlPP9nbUu8xpOjSv8W3twMVkq2
kuuwq2NU033r2HVYU5Iz14/6YllDq1rZ34BkO3pVWwwAdcc3qhULQPC6PxIfcEhj
Fas5lOyRsp0gNr0xWlblJlHzAeGgbIj9MD2Sk8FXnlSaPAileLGiVlyWQnAJ5tcO
DDU+qdHb9tfxITZIhqARtULVSAMeRQAfCfvEl2zXn/SZkZqCHy4XpN6v9hYDpjXG
r/1ZJCD6dGoiW8K8sxKwHdWSGUBO4RqCKkdgp+tnlWZBQ5oMgTxqM1vRwFTU/QCW
VVBtRu8nC9JNuaxDVzPfXhGqAn0QijQody4u18vIv6lTS3ekuJ0d2t1fJqdL74Ur
BzCAhUd+WULiwaPHMVQxkwCpZsHq71hzlLUUXkUEIVULEH54fhWqcDpueo8CjWHi
/dpyOXqYgM2j2s5yPRu8BnZNuN+oeVSeG1dQvABkg7mePeRWtyIginJQ4WsSHm6+
aqMfw7hMMp8w44F0z/Zne41s3Be1bAHsXjsCw1yD7jrXmxOPX6620p7nO8ooi7ZC
UIgmF/ez3owrDIJ2CHm3tRr5h04ZQOWDcQdDhQnSZ+Tm+69tbQqpCRfDt1dNu388
CpnhZXlxlucjBfS8nn4iBg==
`protect END_PROTECTED
