`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hT/oFhXBMCBXkklHqgF7YKTKw+pUfqv0awdIaCBIL0SOmkWsacGW092kf3OIzC4h
/Am7mYYWebaZxAzJDKVUsBfoTVwZBLU0LDcClWj2szzq1NWPksdP3b46UuYkZrAO
6psTTd1dFLjiejgM5dKtfXu8ygCtqDU3xBWmP2tfLbWW4pwDpWLw7K/yNUQDQLLc
uRUI09JLDfUo8bskEhG6MJMqZ+EcyuwfY5/n0lCbT+65XwTfxJz9yft+dFwO4uTk
kfRNpDiwlGQdkeUUzJVw3Hr3KU4f5vXrktgGyxQfJCOcaaoleK2XjL4Cfwc1lU0V
RVA0JXm48HHdhwtvbSfa1qusmg1BWal9BQ9UmEWg65v/YhLr7fSNWOgvWlp+MuE5
DalkS9fkHXK966Tv7cr8zrmywVdnJY6SYQnqEM8E4N44JrAYdWoI74WVfWJe8thu
uaX/qgZLjSlWq+06xmRxCzhfVdgXP2gAdSdrKE8IiJv2Tho+80p6qh+pRNOqXlWd
YC/Iafx1p4Z7OGTEAojPzJqx3nBE0m6ypes4KXQnL0AJcdy3+SE1TKwrqK+RdlJz
dPavK/Pxmsi+F0Zn6X80elwNodexKrwpNrvGxadb0Wx0nlAGUo8ltpIJWoPgojJF
XFMG52m2kLyNlWqEee0seBOLiH0GwXBfBRv4rB+vTjIuKaWzYtx/pFET5gL5xiY3
4nps+y+EQ0CS5ShRa4CUyppvnr/JH9h6Sr1Uo6i2TGTsqFGKp2MSqzDDbvTcODdv
vHUctXfr2AT29YDXIsPkwHKxUUD7/qxu52yDJwafRvQ75gIx3sbZ/Dg+Yx9emiQG
e1vK7v0ORgGjcW2744kB2nu12A5i7+xSDYpHeDxbGnsDfJg2d/oAkTbyNXLSmOqy
wCesGNDoNkwBUQBvWW6fgkxpSLCs4IUA2ir+3a/Ka3UdNXGhauKB14S1aTv3U0+S
qAk7no6wZ7IWnHontgSKxHnHFxY8mCM/hxUidzkICCcDD2ooOfGPl8FG5skKr+OX
ATsNZhUnX112GDMuwatBiVOaMiMk1t9lRGm5wBKoR+XXIH8uLADtRqOIRSu4bAre
S4LakZ9WTKCepx9r94K4DbO8OkXB3rXhAp5GnGRW7uBavv1rYFSlr6rGjdUUR4L2
x1n1dhtnIacONE4YtYuZ6PXTbjIEADAstom8kgAL5ELbUMtfTOtBxVs3h0w8DLOB
kh/7p5tUU7Yv9d+ZHqEhWx5Z9ERNO/USNNCG4Vw9zqtrze8B++3xKuqpF58PEeXo
yAKJvaEXIJ5M2TZtHeuGfHZquAJe7TT2FE4Jb1tnjcVXJeh+COIoGKTsTg0+bkX+
tQUB3UbkYjJxf63gzl2c80xz6ZDllEHlloTqgVac3Yc2WpD+NA6sTihX+Yvxrm0C
OgUmvWGqAPli7yPGU//6cEj+XmQLc7FYqM7kCQ9miY0hHf2WpNj1Vgtgls0eIiyA
UYy/KL8pp9P6J9Qhc75DzzXbz04NU7+DZPZctoY7uXfUWms8OLebK/R9mQZskpxb
vXW+BJ+OFV+DdXKKK4g5b8aqiQb4Sj/R8jSCpxQ0utb6FrPsVQwB1Wk5AJTsqlRG
XJgXinquNNqKyMiZAkt4wZ9Tn/0tcmdKuCILe4C2SNKEc05nENinNgDXmwTlMejS
QIvQv3e1zf+EwdzddPALvg==
`protect END_PROTECTED
