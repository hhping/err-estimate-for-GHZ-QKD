`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQYn7kZvrLEQ9QbiKN16hMLc7azhxkBcpvFSbWfL/4M+9+dXf3uac7Qd5zEfhdi5
DWhdBLDGQ0QH0YfphGdMKfGEzS++8ikBagjdi91naLBpF2agudvmGKdh9lVyifNX
ZFZV03DJ/WuybtLLMZxAiPEKepxSfzlWCY5f6R4PtSjmpCK0+2qlja6CMskHFpDg
Yqql+RNLm4PaJiLbDnM7WXJAcAOA0mKHsyot2JeTKU9/g40fTszBn4JMAMdTYmVm
yKmVG6wWCEfv6V8rXyghaf3n1gr+oJLPG3mpRUhZ2zYay8b5p5LsSXRIwsQCH6pJ
YcFwTNz5bxwojG/F5YED3MuzcBIU79W5oDd3LsnteT+TJJ4FBojqzWCIvVVFP9eP
jscxhFBF8y2j73RF3+THqNqHJ8IpG/EVYWAlEo/PMgxY1O3Qq9WwbsKTcfiXIeXk
hBhff6BByT4nEQoSV+y1bgOETAQNcgI1fdbEuAcou3c8qzOvufEeWnyIkWcq8CjS
OK9J+LCckL1oEv43V+fKbSavD1oMqWJhPbbxAYaVV+Mld/avpd4T6EIZOoHNfI80
INq6HCsAihPUUM/pbI17PvkyqMv6YWIQq2cyQVwRc+uSnQR9BtyR9YbsvwPwknAe
ID4stOR1BLTrbfdbFDtgI3rlsE5V175GLezKJXZQOdkzZVEkt7zByG7Mo62yJjZ4
y44AQM2Q6DMPk9HrnpmrLGu209W9BTA835mytoJ7WJx+S54ls+fX7AfAGoXkKxE4
7pD5ywERD8xy+se5/gf6iKl6i3YrfLOUxYifd3sUOUxZngSzaEcGab/qwuM7BIf/
AE/c1KfA/R3Y1uSU/lGpyAqraIvxSiZ7drJ94GfYvGBCG7JHZxUrEERRASTNGohr
gRJWTTQuLOCOz3fgNiKpYCHaN9oY5BQs4ZUuOlk2US3X9/F2FOAi7+koH9jWlKw5
nvftSiLcyLzEi1/ARWN4Dm+7oy4x1XHipofDkoWPnirAg/XV0f/xovRhZXFcabMg
u6KchSNIj07GrB8qSUmHKQ1BVdRrXoHt1Q0Qs4oe8IVxAkCqq9y0TNQNPXc7J+rE
`protect END_PROTECTED
