`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MwW7owAAgi/u5OD+gsnOuBNaBQUEQJLdPoIpQUyesAkHnnLhW9mIx8ZuDIeHnE4
Ut1AkE0EHHOI+dZHUP95CLXgKRLb8J/tQgfJYIKXkKnpVJMkKfWGDSQBGWz8iwFf
Ddf9H+U9816+sLQljvs4En5GD6nG1gaVrKSFh44fGkFb+M4+UR1HN5RC2zFYxabc
yEyESnZ6lJn98XcTceo8pViTTsqEzCnv+b/1NHojVHEqqQDhCVthld3DP3sSDva3
WxZzsi1zIo68EuZ/s8abrgkS6UQMwurz7h9Y37PP8W3XsfCH54FQKA9sQ4kSzYMi
8m3pFJmP7vdN8mDVQBiaoCApykbA+qa/Yirr3pxgJiCtxJ/lzGc5/IViiCSabFnZ
BKSSi6Z0GVKc4mPgTJf2s69Vyuehhi+278PeOb39A+8W22CcPwRujH8IwFINPZhJ
w22OHyMHtKt0p/riKVHa75Evcf2ZVDo0Ah11XiLNTR+pErxFT1p40P4QwYem9bY0
fIqEctUPGxg8DDLr/95+6RsCSdOQNJh2wGAcpQ9F8AafNjlD2bzk0b/cG0c2rVY2
nLwtXgZl7636GdRm6QyxU0WWkVdpSE2focmeCTNqJXxU8qw0Me96YKPgJ9IA3i/3
rA3G1yYkbCvOTSjvqvuC1mD2fjyTbHFklr25NmkoVU/xtQXlU1b/b4slIhxa+Qd5
o+ZQL+plU1K6xqDqil5QtklZj3nrEWy797Z8mpbHAg8DVaOlA0v85kTCUvBc9tlc
t03ZGFAYxciuxxhQy3Jc6+cqa/qNv196tIzW3/f7xiqW+v8xz6akduXGWSYxeD7T
qNHDOaJ1ovcCy10azZCtvKKtDcK6/cttrHa/wLJRNlFANaJ5w4c2H9dqZyzmxDUs
ZL7YtZ3aGXwp/N3sOHF6yyLYZk3Im9upg2CKuF0jG1JItusuRNxKzvsYc7la8hSU
IA6bGmgwqXUztvpoOXyMJzzzWI5v9lv9Sv0JgRY2M9OAvT9eRf/zqShazcnFaICx
tDnObPHMwEaj6WqUvxMBjSH8I4Pc40T00ETvB3aBqILxFAQiw/YNJT/QlzRRSp+b
E4rK8pZ6TX6Y3Aexm9loA4sY3XPSTfzKaGBCAVn//T8qoFBaA/qt+kGvw4B1O61x
dOgGDBcKqzK+KW4cybHNYj7V1a2v8hD9feTmIy8+qTx7odQDpNLo/rAGhWUm9t8A
CyuGDWqP4oY6iV6MJc2KDbrP01fXuG4d1O0vRWJBX3Y0SzZZsx8TbQaXnyQ7JQ++
aULwc5HAN4HlKwMvTkY3mP70xpu3g/3GIasptiPFvhrlF1Fd5KZl72IJY225yck7
MsJKq65ukWxuawHwlFCm5GWK0FtdzklHfMMOuD2UtdAsdKoV5n73U60Sqcy4Q5ii
/VdYumFyDNKbvUIYlMDQiTb1fGddtTQci9w34qBJC9Th7YVAKGsOMvVQLfKr1BEB
/7CYMAPShQpD2Dcc0lTiXDlmXCLW2z62my3gCvDdgo2sNJK7jr/iTl+t70byGzf3
yKStRP1kldjOdQcHkEywjFspQHEZkQ6qx5jtPQnLoTHMzRvNgk/hfts06jkqjf4u
zk7K8Y7crxDvYdJWHUlSHlUMmxT5uzFXnCXIxpNAHd2Ro1PMCtPIprCP9cUy9spj
p6l9E7LcuE038aaHOMp+/5lC3ALw4O5NWmvLKOrtUzksfY+putjXaqsh13OWfTK7
if2bugKGajsBx2PV+pBoiTlOxiz7SAUNZy3ovaaxmFeUcMi5P+FcVgVFG6Si2U5q
+RgJAEnSKwwPCmx/6jwBvn60Owx0gW7J635ByirZljbJOE8kFZXff8eUeBSK+Flr
lTyms+X4zlyIYjpLgr7696j1s1VO4++X34HDpxHCJ5/7pEk2nVf/W8wGGkh6qhfa
/bSdY+rerer2yBbLwl6dt3WFCmlRf+KTJExxzhtwoxNCfiLWc99cWkqOSmjDpJpn
4CmsChKqw3kkMioUtQ1xqxfbU1iR8kDcv6aUfRJ6eP4oJ0cjDO3EBjF2hi+w/a/G
yJYi+BbmbI8WDw7mljhvvIVcHlSvuczD54QW5OQ7kBPcQnx0IAwcBX+dJcSX/2vL
BAeY09emSQO4WpHwUcqpLGpzA7d6+3/EPP5si+C0Zc+2tCOBNXP92xyxEDy6BYGd
EcPOpmuK8BNaIsAIVgNFnh7/Voo+Dy5hir3G6uQMhVkQHIq6CUUC9+vIV/1s1o2p
ziR4L+uxON9STq5ZDmtuEBuS3dxc2pa9SSiErsYldb18jw4QzK8AB4tAiA05ly5b
RAZ1RuHDudfxKxRva6fUO4JsxZb32ePtl30gqAQt/QoIBwR8u/9lQ5/aK/4YAAjb
htLWbTt9yEtrzKjZQM+AgQcL8MQt+dd6JCj0x50cdHLSC8UInHCuyeWSbdgbebF0
biUw4IBLHUWAjCN5e2CdTwtrK3QWqjD0+Zb/zWnKIIRBc4bN3QPrwWRqft/NIbbH
sk1P3f0RK7SF+9MPjXmhBtLXxoJoV+b4c1/BSscmd6y4fMc7VoxQN9frwcqyJ9ZQ
IxymrzdpsjcG2AcaVcW3iRbnE+7bKfICx/LjV6vZ8CAOdmWdckFLWuDqSlHgEaWB
tsfnQ0RFT90hPSIYvTkdRASMDc38vYhdkEqBqryp/lXnulmlNEuf55HvR6HJ3C5q
3OestHrwdE0Aj0jO3MNmA/N7tSNxGpD+gxZJJD5fZM/DtoldrDMgNbNcts8HGLaZ
EhMIBgSySZeCJ6X+pvloPvWkLYe7387gegxgj3ltum0jjxjujvaG9/9ELD3l1JGo
DKk8LNz1FrZniH97ORYRfvZZMF6B5XZivbtjRNbDb8wvqb2kisUAhnDewLvibo2B
xNpwt3if3dAqkr2bCFJUzaMK7rLDm5usJ3pm5W0JbKDXtz4fo5gbmzAPsvmbffQL
N53P8Z4msJKfPL/09D/6bDjTd+/i4H8aT2Byw2XFyLKEkoqPL3+xH/sPIBxqYiPo
o4V7s5CzMPrm1siOQq35oxc9bTEDdjAvSgt9qmdb52ZDBu5qQMOMuxtPQvy0dwFw
w+tppBWar0pVfXj5PVC+BMBCOQkkG1qFM9WJ9RWZeumIYqPCKRgFRaxcERxaazvw
RnxfqL8ggCnb2oRYiKv7W2NrC/1M5krh6e+SLLbOy4Xxd0AUhpzfofKgAYpNHPQd
orlf6IdyWSuKlPhIADRUC7jWLA24M/0za9IGPnTPpY9BYw+N0sh4sbi+6+iK0n2v
e8ExUuR75TKz/5SgegR8s7WcohFWGgIF7Z6Ip6CNEEnrp1LbzLaSE7SFg3+BpIIA
kMIAyhAzLExReNatdIvJf7G1XtZLVx6aFCiL5BNcrSYx174R3W0vqdF5KJkA0Q+C
ysfcREgZKmZgOksU9X1kd1QxOyNkVRbRluUyOMOTwDC7AJ8RerOj6eX3OnO9oBtU
RkWAIiWYfaEAlg4BIbz8w8mlIXoFxX1Ws/UJ/9OUSp1Y4HROLALDsY9qGlEqCNEj
Nf7xd5lrmrIyzj9feaTc5ReSgJ8DbccUWmNtaUytzIwm2qeeXjts6xU75aH2imXe
DkBvjW5TC7YcIfnWn8Xc0PucfHq6tBn9+7LyKQ1LpVE1TIusCBto1d46TxQtqgGb
VZQIL7+fgQw68OyHXhxgXq//u2rNzm0F6+1bqEFjsZiQs/Evhob5VefOsGqelDVH
0yufD52nfZPJN5Y9fiQHWBaD3PKJFNS9Sv1lu7NI1pcaDz3oGoZTFPuZszurtisG
8FW9RtxXA2ODis2UnotNNrmblAmE1KxqEZBnCr3itcp/QCvoRohSsfzpUKlvMv5R
fwcUG9BUQOlg6PPH1C7WuqoQOkyPeV+qxh0bhmHWzxpFOPuS3SJloPDL8LWnGGrO
EyoOWO4NJfXJC0WiBmk2GpdZgGu1dvIPsT68Q4NH1J3Vqlm7ZBEBOe7kNx39fqXG
aCkRbPWvWjAr2xAPMFiaIckopmpTR4iH5zMq+hiUZu2idu6Hnkw0k4MrEQCTZGAK
Ryo9YQmc0POBXo5IFgNsr+lY6Vct2PbIBEIoAglhFc7jIXrcQeXX+G6yfKX6qP/N
f7oy9lHemthVpd9/6yhOksicY90IB20ES3ker1OwbAg+qm3/epj+tz0u+gSweX16
dGc1Bpf28VDh6Jp8lvdd1vmDLuZtHevGwCcRL+OJBcnzGZfhCyarZsAOt691Oxc3
Ob79Y/KZw8OswWZF4vWsRlCZCZiL75b5XtlPyBAw/XlhVkWHkwoS6mUxlBpkiLLF
G3ZaOzsXG1jQ4516d6ueRKcBEZ8WR/1lyoRzCbYSYYz8IcAWR4H8wDCcRJ1wTgJY
mDzCvq3sODMIRCD2HtUvxRzeauT2rUZusGjPy4iNpsgOOg34trPJIDR+o9JIcfel
Qsu+TKfY5GRMbC7x0oUhIljJOmAGZ3h7VKDGyHXDuwMfUkIGn+NYVEDUChPm1o23
6kyyH3OSP9prl6HEiZFa7Id9AvyJRzKaa6vh+AGjunz8gHlRhu+hvk27vqBFdILm
xs9mCVjqpoeOWcc0IZCMJlBiyhDt9pO7TmdmGLF/WDA+D4yZAhimH2f5NT0Bs+Cl
y6h4ugCYAzKovxfr1Hg9CP2oKTWFhwlrTXH6C73GqsZy2QZMr7BUrtoj/P7kGeXS
7VT8jzseaK8cBRkbAFBpLlIIp9ADsj5Xuf7SVxahtZzvfgkQe1ftX3nsAW1pzulD
25V6LWKQ9bZywMmci8ju1FUeZHYQnQhjztOf3lUtawLhHjCLnQNSe1RLGBtbkKRn
4Y2O77X3HpMNhUnz0p/s3G62mab2PCYqqADZxE6SLaZ1huu3mOzyffluJWbj4c+v
i0SsPgaOpWlsKvbY7K6WGUhLTjhGYAuSFopHRbgPmt98YvwL1r4tRG41mV8voCgD
m6zaRVRKTU9wc6qwJ2LWyFDjTrm26WvEqS6OeUsEMYMqk/+afr6SQphkB5Xqo4Mt
5I4Gk+lsPTG8akh5qCR0cCOS/97x4osNNFNn2QvrFdhsAXzK8cc6HbNsGhFiJIM7
qhic0B1HjV9mgSS24BlkUSfra6K6E/YRrW0IkSz4/oQtzKLOlxEBBRrAyiFgIZsM
SlQ6zQjH59NtBwaCqCEa3QIGaJoQ+rNmOE3tiMTUdsbmh1lgq+uaJZLcBM/PG6D8
RdnswBiYNRpdyNYf+zZ4CiWchMoPkN2PzVDZiMfXzlUv5rrwa57vKiCQesXS72w2
cnZMnE2d+fuj7BbT3cU7tlOMxCfVasemC/8XLD3HL0ZniYCuYABSYS6dDrRP81bY
LRZLnOPkCwBqXEzlBolg3N9ACu8bLXweM+UCWi2uMppKXde2WBj53D3RpFbvKvaX
m2PZR8O3dyeNpCH5RhoBvMx7BwiDaClak/LGLADaEQ07iPEFutSIjsDq+8O1nPDS
Zz18WlWycZSVJs6r+0U1R/ZpnyumndVWN0mJ7v3Kv4jbXPn95tCjRjS4OY/Qv/C3
Isbe2v5TDJ9A5qZEv87Ms/1oxJ2MdMUW+0cWAo/062kf/R90D1hMbHbCXTlViRxB
HBEMAwdxm7GSO2wPX8spii7Rwoy79juDudtMm9GYaaI5z8u8cWQks/RSCulJUfo1
iRK8YdosZYdZ5B1lEdmKRpMmWVUcpci1D+T4P+S39fdtBPdU0A+y2Yj99sOGjUQ7
7frGjq4+viNwmpa8TbOozH/R8Yzl6CkErJCmwLQlEVoH9rbGumdz94ZKKi4qC1v9
Bwczq6HY7QrPqzfUz/SnletY8b/jTjgU9FM+dbpTqrj1JES3L8TxcDdbefgdS/MM
9/2mfo4f+tgPDOnMTHmtJukmBofccPNExh5ujeh7x9bfGi30c1obWxroPEwA+HfG
hvp9wum7xjHgr3tk/YkbtNYPeFv7y53RJC4Sbiv4GLPem7DaNrxqbvArE5i2jYTr
fJFqxiMsISLsJqesRHbgmUFcHOp94XjX3uEKVrioFRInH6OpfY9lvN9GwnFLwEqw
PwlIq2JOLDeU6ViQKLxWuQJii9sv3ZwWc7q7EE4oattXoEt/m1NX1fubs2GKtQsz
lxn8VzOk0s4unQ/Sgg/f9FowSeJdUAh1sgu8bF8yVrdnLOuHHb3uAOeNqmFkpAYz
IFY64XIl7fc9JlkxmUDh26CxawRWt+q3tN0nhUbd+Pbey8JNyATvsIplIpQYaBOn
o/0LytHQqkEYcs4ReF3JW+vo8H1Nqtf8jhss/NzIf0NIkWvGikbY7bOOgDTAttA2
eKEKmxb5HOSLeAbyBgVIBR3jBDIhVO9eu9Vc6+RAuFlgbUlB1AlIDWcFs7QYKugt
pgXXaXUKZfmz6plIvl9FhQPsDLq6kUhQS2Px/iTGlaeq8baxm4epcDpETLfPdR6C
pK6rWeO/qon7n9L4bZcl2OIWh0UTjwej2WOKg68kI5dXlmDcNqC38sgwu7rF9r96
HxN8HlwaUoL+qLa06OSgZfPMjS4NGz5J5A6OZNRZmf9eRGB2JSiL7Q/Jy48TCbhO
z0fHcqxm6jNNvfrIyHSa7BwqbsVw2qNKncDuoDbW64QXXJnTJrUVle2JYoHeGq9S
APyqJZFtHHQ2hAaCvJsu7NIOoS1twg72P/ZdUHEqaGU6/ZqRXgwx8RQxIRuWPqcc
AUMFnrzEvX29lm5ekrsxIOhOYddAQ/9e29FAh07lRBh26PxvLyRE79/4Z05QwsE2
T0LtGVJn0M4Yy+DI6+z5d254uSYFjO+44hakNqX0TxNqjy0Hk17CMuPVptjklejv
q2TgM+nJwJrURl1b8NdIt3st2EdR8ugTLT+h7I8ui71hU9/GxhIX4Ti89VHEBkhd
2YB6ftpf4X6Vq6FJ+MS7rY44P41SKsJTSPgrvCPoCAy/SHIcR1o99aT2fz6veYs1
p98SS8u5Bm3W24TQgdn1UwuIK5BiUC3nfzNNQddb+U2DAlJnJR9/DgniMe8k8wDi
GcMPvyeOFksq7lGvLylI2tROdmgHQqfE/FWQDbSi89oUClf/QCnNzLHPmadO+zHQ
GTqwgDKK0ARtCvyJ6C3Lzsa7idy6VpSAAx18w/buULksUuo6Gjb7fqPqcbNxFVbp
noSFh2HInVbQCo9ZQi0PD5aaE2MfNitOZ2LR0AkZnRhvbmxZoF8/osH8dO5u25ky
vEE5I81fGKs24AHiy3dWWaeEcgD4xvqLuANJD1NQT3B+PuJXR6ST5iyToWNQuCI1
Kxd6MB8vd6jpoYXDROoVlhe8Z0Q05YNgvFFEyX5vKIBIgFd9skl1pLsETfahYKUL
GrYb+BMdmYPvkLN+3hIIFs+HhSr2C5M0wjQLl1cMiJOxHY8DXVoOiAuYdYumhBM/
6uIapVQLnOIwdMOBDeFW9IxF2+1AcnFrDWU4tgkwIxgtvXqX8u/A7jNAPxq/2MmI
xPqTiOxjRJtLvEU10mJLC9iUXiz/EVopvhRdbB9MwNrTMk4O72qVtsE/tQr8RzLJ
VgawJxwrKqrqVz/dhxGHZo77/EZMmD6KFQeI+PONCE2xa82ptaqoVC5Uw9Me8H3x
CJqyjSJVzoeRQYOXXCiur4w5TKHNWMNA3JiHT2WnmuX5zg4toekwi6cIYySZjsPR
JHJwjRUxU91cvHT7guvBn7z0E6yq6ADej+bVBPp+eM8bAu8BIbfA2Sj5hbQ5NvqU
T8zGNAVUXL00oFIxnMQwh7qoZgt4hQ8gpxtZ/qL+05SjW/SNgS19eFDCbcq2z2UR
HJXlHS3NaWngPJe+VrUl6zUT0QtAr/AnenhryNyNXqxOMXNiVvucOOE58froY0N6
ZYSwX2svE2uV4ZJaTW08ihxxPy2+u9VXnfZZnqeukrILs4D0p1RDOXxPe4eFrzyM
ywr7yMSCfWTbqZtitJR1V2fwoHbFDwe0J7nFSspXjbWJBNDYqti7q9lI9FaU8mf8
8RlsLjGc15nBjyUu+eowbCjcxRcEnNghILmDKJq5EjK5UukQ4BKAWwscu97HSGlb
hGFaFt0Tl8UdsHpJbHkBWoscQ2k3nFt1ufjlab5HfbNd4eOrLZ5vfOnNmUhc4EVG
8EEs8Yiy92FgihNP5WdxR2zZ2xQbPdYKKjjZ4qXlApmW7LQaPEWSyPagO4NE2JSy
ipk7g2fyib1zAQ1vus1qMzo4HvAYCMOsPEt2xWOLNCptTISY/ZrW9VYlElFzp3dy
OmRawwZ0eWr1/VFdgtQY0+E7LhAtVqjYQJ/j8huBzy1Z5hf/iGNWWc856GYAz9UA
15QkRUL503X976dFmZaAXYIvhHI8F2/Mm1w3usR8Y52mvHlIMR6a+YtxNRy1M8wP
AArQJ0pHf0MrMWLJmryeF8no90T5OqnM02N/F1RzqxeD5wbXzJGxYAIjTMMclni9
itZKxLIlD1npDR95hL235G/xRm529oMUdoOhHNsLbmm4Kq3grOXiAYiyqCmiXR5q
6Vf4uBYcASf7zwvJcfRQjNzVhHPQ9ziHCRgN7L8ZQHkoBpdkMHxZzbGxQ7ssu/dh
+/v74QEUT85y+XEDwSVKK3A8dAmF0HJpgZz7gbkgLolRni35p20aWNfZK5bmgPmP
Qw36h8QxmxQl0mX9fqDS9LHzMuh+OJyB1vPj3qJVuEa82BZwU551VtZOt9Eqshfa
95TU+Ja9kh0igikWahIYsn5Lm8jnjB5K/6IaNKwC58lVbv9gAnIwnT6SoNA6S3fW
mxHHRo++51BJq29PFHWyDwxlBPYOkhJl7xnghxo2IoxyEmOh9nGQh0WN2RbDNw1w
0+eu4H9gRqvKvZb8EsXzmDH/FE7sRnba3wYE7vTIGK0X7O5REpy6a9jcRRGXi69D
Yi1X8CLbYMu4M1NfNNrvi3gf6JNMssIJBMpzmStKhFh3/4XRF/S0Sl2d2MMLoz+u
PnqzY3KEW486Im2pnfws4NEBitoc9YVvTCq9M/Sjksgk1ZtkGJUgLwCfpeD1CVhR
qqrCy1PvmY5oxh8fORr/ENh6ZGxABuPM7Ihsp+5It/craLT7yGSXMIGFFJU+CjtH
6c6hp1x4IJH6BeGFY2d/4zSnAWqWjC1Pv8L1bt/z7v7Ox1b7j0QaIc7NH9pnTpve
HpANO7ucX3hhFTBFfYpNqcuNktqruCNDKcYclw1HFqF553yLcQL0pxPT1x1/TNw7
c5gxzkiREfQplZL9LWt2iOZWWTQiYZa3WKYAAbRK9Gn7So43BkgWgxS2fmhTeb2o
D84XwtxC9GtnlDpCXEk3P8H4hHbXyj8KRTFJKCTlvGH2lWYKJyiqRqu8hcc7FZJj
jCpirqSCxfDrkyIzLJhfgfI0TGv/RWAqBJzbaQQS8Ia46wokxd42mdpNGpWlAyTY
tUDu02w+O10YDBXbe9c/sFbRrLWKW4dnxtBlN9HbLOF94C3sXwWgM+cpsosrKR5B
cXWF8kU2mWwPqDSegehIxKu6HU5pTQqzcYQiLUyMHwBxlUhsNl6O0+Zcz84bMjbj
kzcv/oCnSmu5J+9AbMeOlYzH9GNVVcS6Kleuh8hHsEibnMAi+tDM0e4mupgQjKMF
/PJcYAzFbd33CjXWGtAls87iLtsrpxbXo5aNBo3mVVFtyotWC+8K8C2iSMf/24h+
Y6pgJgo29Y7S3o2gtrjEDWw36hiVUF4m3jJ3rhSDOMe9F/iqgVz+2Chz1XzqgDXu
cNgdcAEvNa8ky0V/+d9qdW13qZy6bkbdd5RK/bKbqF0jFIJfA6dT4Rq0/T174QEy
i1Xwf42X9Bd7yh9obLzzOYBUFusaHDYlbidGN4Ci2mHw/NWYB9bwMOhUTyyRtcwo
xjKRmTNqqXAxFJPOR/kFsfdl35P6yL80EdAuhkBwFF2lTvAQEE7ufh9s6bJ4DfIr
tmcV+nRKKmxKkqn1Tby2l72+6k9PPcVXLWQnvI0tDpbPVxmTbJpsreviK8Wdfjkp
KriA7FSmsTxVowqfZw5IFkgd4tkZbfOKT3SIM625BgRXKaIKYj+dVIc/5seJC3o6
BXe/Pw8dEOsHC9swtaik3bugo9crCw8aAI4ayI9evdfwElmPBzMImvJfClK1e9bt
9h18C+bB+bt3li70i+yduyRX247XELKv4+jEybJwTMniPo3o1mv16PaI/eY2SNoW
Ye9AmBkhLf2zN1lcezRjtXhSb/lkcQvBnGlJgT2ICpJEoD0z9ZUrKou2mVtmt5d2
8R3a0UMjsdJBJqp31hS3Dq3NkrP2us1MT2I2grN0SkmbRBoKX7YxQwRwZNJmDnrp
IVuYdsXX0rBxhrCyBtOlGxR5Ys6H3kULYZeO+2p3JZsBwMcszUJ0BXKaBJ73EwJb
xq0ZF0rrGb/YT/Gfdkrx4WgX56jkbDEnU3+/NfGR3+fFpJcp2RM7F8r2ldcje4jc
CrhyRmepbGZbrfNxBiTfPBDBqzg0W7MZDmqsr2jMLp6CB8387khhR2Vshm5aspVm
lnP4vtZFdDAzn2uFaaUQZDnafXotjDb02ZnNUWcb+5xqijlaqkW+2BcKgHbRr/RY
0R1qPAcpAqvvqVhjBWG5ZJoD26smKnCeXmw+H9NOCW8HPscqlhL4OUdxgHf64aep
1sgblsyO/6/GnO0ii+0JkHz5I0Scpq/XYd465bP7RiA8QerKmRvZpCMkZw6q46/M
YP5gxunsAlLMZHJ62HvNR04SvOiT8NwsMAXFkczZcy0zdW7nYDCP/88j7xBIhFqV
I0cbcip8nsCRm8ZIHeTTw8s+qw6RE/b47u2dQ/BNVjgtCjaS3NSSFWzi07zIclML
UsVzfajYOIkQqmEDnKDZxGe6JKuwwOfglBbyv+YyeYrRLdGCXpFm7gXbc3M09gZK
sJaBpXUo2VkFyi1EFjh0dMgcn5Wen10QIp8N7lgF6v7p79cptNN29iefno9fyKX/
QN621BNX+sIOYJH25jBj7upM/mwYL0aPQJ6eKcvMT0Ele7f09mIeNBC5pOGLTh1h
pmtoWNjFehlJS1oQLQVQOK9h7nKqBEcz3VSE65zeX0G3vElFS4y0xKJGS30Zzons
fxqyywq4aXTZsc0Gne8UjLzBJ/qJPHkbbEcHSxDCSrktN+aBk3LJCor51Othrarn
h0vjIGKDUphUwHwe3nsUD1mC+QN52Y6DIzlGdre/ZUAQM7BwsB8o44ntQSE8X/ZC
O7kguVb88Q5xcYxUd2Vvxmv0AlBYxgFb7HSfoIeoHhnTmf5SiF4W/NlEPxT/ASv2
`protect END_PROTECTED
