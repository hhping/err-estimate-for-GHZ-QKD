`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtvjgV7NNo5JEavE6o+Vmh/qo5G+WisWgSLIHVxcABDm4NLWy2fBFWR94J9h0w6C
9JUYhyXy95QJ9MeYqLjvwYocGsAdvxabP8zU5y3EnaAcPYTRSNJKE4eEMXjXnIsq
+dStRCf7wfJBFJmmwZKOD1Apglu87NICtzn60ZjSkjRf7nJecErboLm6UIPV3MJV
Hwx/S5my0AogtVXTyOaAb90ydue327N79LSpeLuUWkF1QNs78M0fPhErdxsJLf1g
hzlpji//clVZVrie2EO0Hj52SO6P9CldUmST+YuGywJq0FRR13F9XKpBGt7iuB+G
JeK5H4vUP/r+BxT2OCunR/GYPLcVRgsAy6zUx/Vt0237Rudw9nIJ4bm5S+C/sx/F
Sv6DQGF0kMxlTCdveJwOTSL6x/on8woMyNz0nEEoYolhlzLwCqn/PkC6nAx3u1vi
WyFf7lSW8Wo9w/wvqHFpmhz/IXK/0ArUFKb+xy9pM7A1ZAkOL8a8YGSie4oKsvfi
hP1hkgMpzwACp/qtYfBU8va/bvVqsl5HbomS9L5q34sleYTBYQLnOzLkZVg+c/wU
E+va3DDo3REs+vU3srINet9Rg8mZJZourv29e/Tb24Qwk6ndeREOkWTIiWisXq4j
kbaC5/jRrmAlUkODxx7ssw==
`protect END_PROTECTED
