`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r63wBX9ejAMjSi560C+vLt+DMPyUYc08YphVwArp4ynUwwtJhVG61B4UAoQt0YT/
mw81RXf7tMBnNA2kGBfaDa7gJL1sy4+5MkXQsU+Q1dMAsRt7tVbcRyWQpFOcdyPi
6KZJsI8rBM6pad6ncQMGf6aZQHGfo3WQ0jpDh4Mtc5vDwSfAW1Uhbtrx9Qt/MXni
duVIODf4ISV5kkksp4Kfl8BbciBcG5vr8nTyiG11B3gClHNwpp9Np14VGy4Mr0JO
oXq8XAV37mg0AbmYS/vL0Lo9tmYWTHB0s4+pWVoIQfelC4uBkddnk/6C9I98x6QM
KQjnAYHPxWj5w6vQ21X6VjQsXUJbyPAGZVGompownyTQzVma0eVRAvO+lqpdeusn
WPiJmUZoGAe+35r4wvCrSTwRYOESxQc7feWaW9cc3mgXpadM/x2v4MzkNeXFRJhI
lbBUnQFQUMHx7jpPzBSerioKg+iZE/TXwZGOa+sp7iC4wUtZZ0/6jM0WEtrSHhao
6meHWI+BQwOrJ0UYDgpdX6/C7XAR0Q7Rlt/0XaF0hZ1x+qJRDeWHlTi4TDq2hAs9
VGNQZ7tyRYFzynuxzvazzzoyDlM7RYLky/rYdfy+QS2evma3uy8RN2VuPhvEnyh+
A29MY2lreFbQqqwE0EDSZPV0jcaiuyuy0Drw69VvTjgwZ2iPuqsuVib8j0qNxKHh
jbIdU/GPb6CUGW03UEBbgKzTQt2eio70/+q9FVx1fShn3zmWD2ic5ICUOMTOx31N
qlN6ON0uYXNJVL9qXbpR3iOQzFosOESOVSZ+YuxXLbIYmZxlTcQi4NkatvUXIylr
x3hdKTufFuinYcRacT5nvBDfzWaB7Q7esayvi5cJWKlK8n9F0iHnvdlrF2UQ2d+E
8PLrK+EvVPzzqy4bBs9Ac2mAYckD/RT/P+pzkTlv6v8QkR8XCZ3R4ZK7Ie3yQ4DL
MI9axVsw7DXlccofqr5UthFjXj8+yV4HjHPGnlKQW+2YtOz1/ILQ48BYWHvPyazC
CiwDIBlCeTx2vHqWEtmVLfUqMGUxUnDd/476APsFxZaD6Zzo0oEJkZdkMj4+Nxbd
FFk787+6kGekmN4EHgTItVxqk0NBAFNJ5jufiYRE5m1+OyjtIOTCqb+IgYfTpSB7
k7pMYaKiR4Bd39aazTFIr6iSVsr6iaMPHUNigYNvNr6NxWCyvk1n53HgtbSndcVN
2yWacZIdI29M9ZBiTb0JU2/1x+L2+VQaa9x9KhvkzgJ1bvMzQD/4IlLuPNJ5T35i
O0JN+2Fg3VjXN+BOnWghVArgxHDoYtiwbJ60MJ3gbtAc5Hc1+rggEkL3JMv3Ni7o
KDkruB0jG/gGKrJRnUQVBbqyUifEP1FwcDzDK/+bYECDxn5q5fm2hlJT8x8hccb6
6vTN8akYYkM3v7HgW7CuG2k3WxusWOPr7vfyjg/Sg8emzHxnDSl0psJgsCdSAdxB
JXIWoTMwgdCdvbUtwdEnvhfMrTH85ofUQxGzU2RRJEbSpJjPcx4Za/x4G0AiwWki
uhxiPK3EJuMrRIFm2LyA7yBwud422Keoi7A442NDhnm4lIGlkAhPelJMD6SIXBlf
PrURz2kiBx/hKYdYP4AAxw655NYQ3rBN7LlsOhBUzbGBl1Id7TIRSdqvDZ5qXa/m
bNczAMSot58YeJdNfeqwAik9xncY8eFRYsgHRoFvzXU6Mj/iwAnC39K5yjUlrNji
zvZMCReqFCUnjy6Iw+oM3rIOx6xTWM3Q1V1ws7emE8IEfqRYUZ2Cg3+8QUJpb68W
kKOyFtzZjeOAIY9+VQsEmU11oigWTM+5tPu3EMvoocRzkoLaJSBHfsseUVZOElfh
XHCIukkKrUARFSqc2XrqBqpZMpJsJ4uvngNMY4hjP2xNUYhBAxH4oc+mZeoSseJk
Z5fs5qucvWcBXTOy+IZSd5c+ypV0LCRV6OH/+LLoXGHKqqpTZaDMa0oXHuFFFaDl
ACxFvohv47+lDhtnQT+tBvusp/DE5plQH1IjwY+O0P+XD96dzvMZ/yFLwWrIJl/y
uaRlXTsQeRGCZDEG7a44m+AkMDLz3UBZgAATobIVratOV+Kx/0jJ8B/3fZ2NNVaK
Cy07jJOqeJNgvaa7XZXl3uDq+9W1bCGHN/jLdH1toOtywqU5ZMe9X6w5MVKBILz8
eomhHWXQOowqcza5L+mQ2PvfqL9OxtdXk+m1oBWkQMMqd6plxfbxXMUkBqoUdBp7
FldlZol1ZMo2iHFGRlwURnSnzfwZNZ9A46LpTWZsLe5rdbvMF/VSI8vU5pE2mQom
Bvvg5rLU8ffaZW9NKlS540CqfwwMWxNSrJVebYGA2zhYSkg2eAsFpuybSI73tMsp
Wcmd3Gyfxnsbe9As64Sd4PpN4UOu6Hp33c4iQbT3V3tVCZcb/8ntas8swQeARtwY
Xg8BgWMggF392IjKoFLY4K9IQAKB18VgAN2uXsZ/I6tgvjy2GQAlRyW1IqnuDeAd
ZERJPwhZqKzFupv1XC4iGdt7dKiRhue6XA4zrfRvDwdECwxsllwiuH0yacjWLEdz
3/ppvP8vOsJf2E9ta/Oud04HXjMvcLKWUAVm3Tt172KD6RyAtlsoeyaiTc6ekYyn
QVWSL6/wEvflHBI0Or0W+nA/HscgYdakQnwWO6pE8OCMccrZcBCJx8R4jREZz8BA
7gbo1eLWwjxEYvkazq0w3XU6MLAKdiZa7RcJHG5XKpSKu6bcXBiWLVHehQm0sLCU
HKowWWx7MybHB3wbU+nkF+wVQyIXmd1r1HExvN+jjjhlq6nxiWjQwY/GoTuBi48A
EUl3IWeGnLSXGwnOr5vwq8tUv/ySrJ5bMFv0PCYUwDOBHTBd9iWF9IJ0elercZZp
+4BjC4k8Sd+hmDQ0tXI7W7N3s9af8MlSPYpShlxU253qhyYEeiGQh/buppfl7n+2
KeQ2Vzc0Yy2NlIDvd6uHlDFAytGIXk0eMwGuf0EFY2zmTGj9LXl/N0ohmR/JgjU+
5J1NCRQKfKSKPaPQ6I5Y04F6IeW30nDvj+UANGQSkROEslcaEc023NJRimxG8SDt
nb5ndplmCvw/4VeGLP6lIrLQ29PUZYLIIpid7UsmAKjegVdJDBa1KiiieVYkmgto
J/839fOr87/Y9lc7uOIxTNZI7QIrYjy708sBHDSRapx7hPXX6pmgeORrY4eGszhr
cnLGQiz6N4iy6ETobGkzD1rBEqa5Xvi26tyP8/ds8ngiAYGZY6yyc85M24V/1cAu
kVNq9r1WSSL7CGh/pWiM0jA/S8RrjSbep728VberagHjWNe6y+Bim2FSIOHCU4i8
477z9xZG0DgOSTNNVGfSiP6me5yADhWEm7BI0Tb9JKw=
`protect END_PROTECTED
