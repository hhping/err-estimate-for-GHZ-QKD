`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jy1cQdjYmJKHnhoFYQ5KZH/B2UkHYPiUlYXqRxZpGMi34Gkg4SU8SwqFslZPbY1C
TRip+q2m/EGnYaV+1ReFH+6iulyLEnz16d9mgKSgh24xP0TFV6qaOQsBwrofuIz7
VIySOt8fBXN3K8hyGFYhZWgYIyHrOwFkl4jjmT9uah9XNAVdEmkYHedkll/2TzHb
KSGQ5+uFsaovCoFV/fZ+RNA50bhcMjw3R9HKoCMZahutGk4iFTM373STpZydFfBP
wBjDbVzXORm5cnYjTLev4MA3ZRWFKzDOQlEgH7VtRZA0SffZto6E46n5XXAFgif/
yrifbCHMzVGCXudIcSW+PYGQWCeIC5fXtku6WeR2ETygZqnJhlm53/GRNLYUKx42
+ObV8FNCfvSw192cuW2ivmoHCTEdt1HjxGEmHFdGLjOpksrTkbyCRJLaUxTs1W/3
RwqAuMm8Dr24oWt/lp76Xjf4Cu0mJQpGfaEihEOTeUUF29qt4SPL1ayxxos/Nt2/
hHm+xCnzxlO7dpBl86ro/Fp4obGkKzHGVWVGMFr5+5n6Qa/t87h1obaA5YJpiOSO
zSo3j1HqEZGYe5YGmQpFI1JicHC6t/CH1bMcIiYQLZkZAOtpK3W6eKi85jKDi4Z4
Xrk+2x3VjSLr6zH1iREyW/KWi8vzj61DBt51NapuEmkRqDI8rWA2lUlFGm1K1V2P
ANVpbwpgGPeOCNXTIvDOchkzL7Jt6dw6QnOb1TSvaWfN/ijLRO4ynwMl6Ga02U1b
O5vn9+cADUrWp3A9ot4P0dFzLiykqoVvAYT/QZSJvYmTXjBnAl7yYb/1GPkYqC/7
LcCTg3LsbXOitb+A4Z7xSAVcXZnrWo5ETqlerAY8D1oRk5Vnga3c59WLAWFR+MQ9
3PDaEAjwaxNjbnefYeXwI2DuK2I9zkTIrRxVCCRbMd2bILkOG/xnpmAfKyl3ld+p
jsJ8XFsPv1fSDixCr/VxYLQj02x9I89U3J5FDOT80KC0h/Iz+B0l2Xwd9dESbu+q
EEm2XKIOYPORNwaXV2yh7Jwmh1C61kUH1Z7lUtOpleKb5u59CG69BpuuriSKtcum
gxTnIj1LxNJL2rrk6j+Nq1Uu29rBKnVPAaiiqOlDX/Xo58ksNcq9FVM5y6sWtZuP
ttFlHe3ahc30s7Nm5CZIW+6hAy5QBpFLhs9usWPmvWRnV96/v9mVGue09nVAsqHZ
Iao6Q1ay4N39tvCEDzBJgU00v/IwzkV1X6mqYT1ADuWWQ7RZuZTOYk4DabSDbFrs
kMs5XkCwW4KeyVjfTjkBdw==
`protect END_PROTECTED
