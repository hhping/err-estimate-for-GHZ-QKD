`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVyv6cjvuAd+mILmWvSN0uusXLZ0h3xchP9MmGX7F41VyrGwk27EdQvVXNRsq23F
UBWWZ2O4Ph6XApp3iOzDxajCdfVGtcNkXDGDOqS6I/ZB/EkPU5nJCoJJ6Qwd8pxW
rJEcYmZ0PuLZQgTFUPqd4GPPwLoSYdhYcqQo33C2RPaeurNIdjNqSkOeGkGE1kCv
Ti5ukDN4ug3SrwU93rtZQ5iyCrVzdKeVDq+AFa8PkFCf75HqAXv1Qi1ooGRuzaFW
pEl+3PjEPmpvZlKWrvoUgLMmKaHvQsK72ZcSIF5aJuyRQt9PJcQFgtCFajbHRWs+
UePfUZR8ReniweDujUZ3jTkBiGpKBP5myEuijkzq5cI79fbpFpHzqyX18fNivjgg
GbT/R4U2Wb9P867/R3BtToWdCP7UHEv3iMlPh6+ez3cGDrBXmLwfSuEwuRKKOgCi
kWx3D0zxJTOaZcQKJ6X/C1zSv59IynulPSldNTQFphVUZBI5g2xCiDv/hq5IFPDR
YIeHsxM1ApegHU8DiHGBHaGTXPnbVNoY66ZBYT5WlNboKGjnJzE5VQx586aYC6Xj
+2q4D4KOi3MBQRQ6T6DEY2XmbQs3xaoZIOPHyMRXHiZJOr7qKIXiGaAiBgAceeVM
k61M6vWKVIV4giWFY4ukLSY9V7mPJpOQ5HjE/Co2yyYTCXYjtxFQIfYRg16oUWC/
qO0DOC3HgZCpvKK7kA+SGw==
`protect END_PROTECTED
