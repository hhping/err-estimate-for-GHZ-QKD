`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8byEf8ilETMQxvtWpikUdN7nrALDDFrWGseCe60gYcBqE16X9kY1WetJFNktbhvI
rp8h6Wetpg45UkOt+1IooLWkcWQQ+2geLmyY/AAkt+SKNqDaiffWW0aTZslIUiz2
ah55FqwmXOZPQ7XnMt4HpleEaKs00tiTvbekcN9sTM++eWuV3PVoYPc/iuB/LR38
NGfbVv24o0pyFJm5w2o9WMkud4N6O+8KBsv0WgBBOCTj4OaVvDdsR7xswrHaqpx/
mpo34YfZsue9xdbKa5vBnzqcIC7lPJHJ2rQOhQEA0ElSvZBf9xMrlNMP1cao5sJL
eTWVYwAkGZ4/E2yQJRlcW+YECDzmi5roJQJ0sBjjDmV8zPmqKRuqsvxvwKVPZwgS
9avN3+gj8+w15xqTFqnqRh0tQ8dJ3LSXvEFUj5Y41C/WsuxlsBtvwC+rBX6u0DM3
9DlESPvswolwPIAfM/HNAa7CfOcx/39fddPbnusZuMyae5zkT4pe12qI9mLmgrsO
klYgGqLkFu9XaWG9BNXYhAZk/0fyG9vZQmJuBSABqmev1fYyEyOWDUkeCYmFNYIj
obcZg+vlQdcSj9Nkeal6BnRLpruIfRXufnHW8MLd/XS2EySQb3NdMXJVJLqATxP8
FPuKjpeWb8Io8cmD8voRvUeMNn/i9V23opIX1RuB7mPEPukLOdFHRq85MNpD5YMH
yRccBSbSFB7pXYMqUxircmPGuAS1s4Um3w76e1N1360+kxnNshNNlnRx+ftNfIk5
1rvDLloTpi+JgwhkajrddZEVkx3lHxU7ed2q/uMVpyIyVM6dOV3hHjK6jCW1fAk+
kHNN1jnRBWJLUVWs40OZ4TeIFG1lI0YzMjCMErXrM4fcoHwuS9X9MpHcoaZr1Oie
Ufp7D8m32RP8tvcGprHg9K39PS+bmRvmpSLqWmAahWHK/hg/s4CxC10GtNi8Jb3I
6nRrDFCeIjYQZ34CuRpvQ0x+0eC8RCbtBQ/XihXhHtlYSimqbHfvYQspeG/zxcbt
/tOiUjXpMFWH8bLipPqpvsRmC8eZOO+YUIhC7/TdLc/E0mSxTHdgBWitDDb5REKq
x2X1nvBFYNrxKF9G3WVbl3FXqibKu7flJC4KuleXpv3rpIRla7Wu0aePd0APShVS
JSBOjGNYWfFF3NTkWYGB/eS+0PFipaY0xWL3YO64bJoVyUTCo3zqYqBmZFFjRan9
VuPb32Tgm0KZm3ZRXa3BQlahSE0ZGPW9mCub32rR0SwsNIO3+Xt13z2+lDEnCwlc
NFUhO3cndRpqypXX4noPZ7rdwwBae0q/BrF4cU3hJMapbiaX5R8J1l6VWN3EBX2W
9uJsG/cCq1DNMuERPjRmPcc5Xyq5d7QN3qwVpMyzYbpogM/NWaEaKRJ/pSYgb3/J
IsXAYsNM9lJFj+3UUlkhRnNXCx6zBfPq5PBUkbE/p+74lV1vyzUKdlljZWN1doNW
FRVhNshodhflLMm6Yjo2edof/p8lUovEWE63RrGr4Io/ZQfwuFypVh/+ukxu56jO
QvLMfKvfoED4WzEVGXP07f86LvCMVn3/OJvS0BMj5TMEpL4hkjlNEehuDsx0nK4s
nJgFwmNyfnZSM+7tSJXlTK31GJgR1Rn2ekzyDUPs4eGhMU9lWe7GGgnbaQyYTIVK
qTtweaELsh9Hu8F/e0ieBGa3votj+FkL5xdfxbBwnJdnQNnw0BOo58/aQpDSCUSA
xnrSf3hdztsYSs5un+MNFhlFhcjilbxGQvyFlM7KgBBWGWsp7cjkOMPBMvojPyi/
hq75vHGHwzYBypFJyG+Lh7YiXEcTErlF9Mljo9G8CDcQUphZ37sfPGqBus63iE3H
ITmUx5l8wOTE+w4DkWUFxA8n7aDVG+hIEeiQFonQGobCYhbXebHhuTvDeVMuCRv9
8Om0BD/U0T58l4zePaiw8napkqUPk7GPXqLofI6rlU2yvykRyda97jLTBZPYhPbg
kKFfR71PwfGAt6r8ca+Di/8Y7IeY3IaJ5cDQBCIiqPd0yQ1CEuM21MKdE19Pmal+
1Ed9Wlou6qRVKPLgxEexmBLAskMAG9sIghQw6iU0TtjlbfJqgYeEj/JJyE6bO+k4
2JbAo2kNDhR6oyfsivjqm1OLnpl6d70iP6/AyM3l3P8CwLagpmonKKUfEiLgGZcU
hK+W9p0M026m5DzBxGWxKDMXcBJ0xH565DOLaUn9rNqeGgvsHoqxClnJe/Q3ImDX
AT/7szxRY+Lp30g+WUSleS4IbU82rAx1CsGbq8FFIiT9EF5MWy/ZwMBP1oiPjIcp
pOUIN+DhfcLjbzvIEwwqQ/XyWcTszX93wZ/7kr+fxHj/GHcCkY386DiQlRo0KVo4
BSb2F36nRq/eDBw/73Cr4JDdCvp+V8tiEGbS30UWWLZBrCe339BQP9q9wm2vhapn
YNRtlsdaPSigwpwNBvPlzt280L1LPQlMfzDNODj2Lf9Z4rlifrmyW8btiiy2ife5
tRTsBOb0mmP9IEd06WiRo5fBnX9lxrctIBjq7X7OfdRvIf5o4EceRbfLuSp9XdzY
Cnc5nzGeJKgSK7SkWwspxOxd8z1aeryCB/d+qQH+5Uqj0d/bqsj5Tl94Z5q0jxM4
6jXT/F8tjrK4Ffn6FlPQAp6CFH4ynLCGg7D/7ZqiEaw8v/C1WV1XH/+BH0+kUR9+
fhHnxoH1q+/MHKOuBEDaDuVuXzZ/Ff+ySiWht6sFXRWFBykBwAOVNuNyN12vG67/
tfyxXnSCSduvWSdxKHIKw1wFh9SPEOsRPbUT2rGgnkLc8ebvwufvqV9w5trZ/5Ik
QtIxo0W/LjExSKEe9C5fc9/w9Jh//jz5Aqao2A+txfH9Xijy38ZbMBHgoV++x/DD
7ONqTS53wNrYRIBEGJM/fK8CvWJ0dPVaNNupLlnuWaxYQlDKwL82T9uJQN+qm36T
32HuFZ+3IwWdUwOW5iRQ5g==
`protect END_PROTECTED
