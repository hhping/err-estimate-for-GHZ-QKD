`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7Cj+wX7cWZDsAk/K2BPe8L3TEKByZuW811x3MyG3oiBWbynjhPsltjjxEjt8zkE
52dB0kavbjouMViOf4uCqteawUkGVh3EwL7VdqmfcnIECukKol4Ex995OPpfcNKY
3X3uoGj3uPtVco9uut0dUHwyhYZls4RWQe0792+3BYCZr5i5NiA4/MeIRRJ3UmI5
q/f/Ba0zrMCqaMez4c3XNRd6KaL0NS/QdQEW2tMgS0cQi27d/oQ39Onr+aAZYrLm
fKjnCpcBuccLFIXGn4ExyEcZBpXSHn0VyrjvEi+Lm6Ag9+rqSTLhwJSlFMMqP4vN
NkD5UaUSSIAoeKNBvjOYgB/nhTa2j2r0Iw1tFlGvPqDznCiKqohTRbt+mfwFNonH
7oUXrx9ICyp4a2wUPpq7F9ubyjRrshaXrNdFUh3JxyX0adSq21SEySLfZSS0pUOF
TxxXXhbNGU7fkcTIlTUtbcca2XYADkA1X4ciYpOLLWUTtAZboNjj2zqwLLqvJPEV
L104FBk+J1Xo1C5WSceigZVnzmBLrz5j9OX5TBGFiMeIGA32oCebhD5mqkWoKEm5
HN0jj579zbV3aDmJDlQHjQ==
`protect END_PROTECTED
