`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/nTtm4zEX9oOEtZtDE6YyNtI5vy1tt0tZgzNNVxqc/cQrUEAlJtQ2oqkEvd0UU1
m0ZhYq2sHY9Tl4rJtN6Ui6r32NpnPbvX4he6u55rG28qsMoSlw0gC7KRSvYYOkXW
9ZGa8ATNlwfEXxww/bUInzVHLuef+kef+yGu0wdgY1RJnv3zhkU/JteAfXwTJC1H
YcXiz9k+lF1oJgdhgRM9QR5WTRiHNNLIS7E/G+3u9O3RNFJbvIF9yU443RMXtY8A
3RufbOaUEMTznXYMtwENeaEFeFeUhGzyreHSVZHNJ37kNnZlhYA2lKfpWahdvlfx
8suo8HVdG5/byIg6TBaZ5KuehCxVCQQNsTh23o7WTPqDYP7wMXB3RmKQyi7bfD0A
xlaCvv4Lh0/Dxsowlapihm6z5qFRcUeZQE3eAOtE9PwmcGNSxhubBEZc6hdk/CNq
xwD43X7O24M176rS41QvVK2DLWtvjlhxf3liM7KjRUDziqpB5WZ3fQtaq/bW4j4/
`protect END_PROTECTED
