`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+A86vXdZq5AlZuKcshawLcGCnyS3OvAQczYmlrUaMlltAylIDK0yxAAsqlgj6+2
V2MZpdMT7bGoQ7dBp8EICLWTMqWn7XvSaUbVwZ0wme6446vSCPVBePubAOjl9E8v
rn8G1pA5MAsdSwuphr77iX8H3ZKhJkEzKArFMlzaYIBUGSQGsAGDm6IjHPw9BlPj
At3tlHAWJbsxmRUatbrgPP9rPtFXtd9TUwmUAvnqOg3Lvo3+bJ+X/jNrSqlqfYM7
mC17fm2owTom+SCKKj3P3iyNYAvtvfmOKD9NRcngA2gwOzjY1FTZ7AFV8Shvey4m
KfungjkEVQSmzA85rLFcQcxbntsiBC09xm+9i1TJSEYS0d26oBpMVaIJxRRxA0Qp
FQKnvrNG5idUOdfCbsgBSQ==
`protect END_PROTECTED
