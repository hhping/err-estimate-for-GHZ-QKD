`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPdKdH5ZZWNn9hg7fvjX+OUmekznJOe3HncqIVq+pgyYpLMwXl1ydkJ1leoCE7cd
0Mtb93Rc94hYGrZUhx/IkDmrZdpt9vU9GnWPyR9owL+MTqaQw/MR92GxijUrbiLA
SUBOsukMBWohcVeFay1mGlNTI1i2FJVgRFT5TYR4ant5eBg6OJJLPqNJWQOFXQZp
EEVmrUcuQPqYkWILvAnk0zbyLgS7b7CYAnECuLmeRKyPSbwQO4DYUpX/tH+gemJv
S6wcEnBfIcpQPMupHkkMoXOKKgB0ML0Zi4s/nOiQYhE8/GW5pZqq2gE9+iT9vETb
NoQu+DUPIGikM74HDM+4miOC3lwza3euU4Wrign8gRjNb9nr8Mu7zyqKYp+FJAUa
3SbxKlf8RSlBBfdO458259Sbm2JccjccDp59TsEvA3i8RhrfgaBRtWkfxyPYEmQX
+MXuNoZcPULIMAbcm3BFTOpqiuOi3EWizCPvx1FLqvXIeYZ79zNvgZAFrtAGfR9k
3Vd9EU9uw+PuYFZt7ZawUg35rWtQMeqK7XWm3MJTOz6mqG+CTZ2+BhR4y3UU1cli
1wvz5K6QIlGpGr5VNyMNbnXiUJjLxiABapamshH4qqg+r5voj1TFfM7ZtT4rT6zy
DT9nhzVLeVVSy4bnj93qnXdBmtHmjJT3t6oirFoA0i9Oh2XnHyI7/kDrkLytxHOn
IzZIOdFYvrkcGgJNMr5yVSZ8fA+wYNr0juDVwFjy9wtnqdpIddyNXolMDjzUAaQv
i318IHuec+4rjH7D2ET9Qiv/mZyPmLkziBCJDAiHHlVIl2gDt3/l4LsuclSRjGmw
UsBf0LuMTJaav5zM0/MHWm/sM6RtkCpc1PddcjfqfINNbU1O7vmOgN1ZCqSXe08a
CfotNabF/NzJPHG1nsiSjthZMWvgOjm/Ox8kWwSuEIGVlpxd2HmiJARZgemYzLtD
O9JuBMOdvyEpdIN/8R2kyRcYHJfR3ZQq/fwuThC6DuVCClobOsb3NiH/KcERhWC/
ztPT2DNVnyEJoSHiORISezrpo0Qivlq0tQLD77yCLZr4pvmOhPGLCw9oVS4F3+ZT
YXLwI6ah1QnuNhaLC9+2tp0YQlGwr1bHoHdIVj+Ma918UprDvfNrcNNZSWbn2u7b
6cGM5ICBM6uuuUCsToZ9wGwPtmWh6D8xPMaG24ExJMqH0zLP2S0f+iVTx6AetcEh
gtyy3TLhn7Xe8Y0S+EVi9dsuBodezB3siSc2Yhbs/vL6v4Dr08KUeqgEGwSyFBRI
Fb5KNTFt6NAZIzc7H4RDdygnjIaTJc5KLncfNV+PdH/ynXGcPanKrFeza6uNtqkI
`protect END_PROTECTED
