`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2wSmLpLr9A48MR5TQSNn1EQEyChv6uaMpDmPV32x70B/07r7qmPDRVYyg8i5YD3R
1beL5bHLKO/99IBookXqUOosmnC2wTP3EvWoDoC8HzUHDO3tevSqU2J3fLe/3k5U
Cs/8i6hfn0btsRSHsN0lAFBOBSiM+18wu8maHbdsdDJvU+fF3pXO8pfn6U90eRuE
P0OSOdlgatPSSnxE8y3yPHIf6tjZlb41B8DLriqcihQvnqrUCKfE4odPSEgbvaTx
HRDYeROSLwxEoil8kxCzN+mdIiWKxujwSu4CONiVCSL72ZXQBogMrzFfyVEKjxi1
eV1kGLU/kDWYvAJcFw3PTioamufbgSPY+LW1vc2hfoK+xu43KC6A48kaeAitaKOJ
zmrf0pZRdWFbzQelh5FMjGGRD0SHazrcTM5dqRSpDQDhebCLH4Kh2BEbv0XtA4Rg
kMLbLvLWlnSYAq2QKx6rHLvXBgQjGQZBrtrW2buBkWdewChFmPntkptBMZ6HILhE
Y9bAA++da3PnKODES+yPkDYBpHV3A3E1/YaM8ofmktRTu1qEEuOeDmeAoJK+ULwP
dxIuL7dP2q6myuDo7Eh84HnBy+uMaAGgXv4nKJh3qmmbb6TH5ynPcA+CxAI2ipxi
yTFFFRmK4GNjvObbNESp8jV14BF2YuYMjvg0kEHtwVsAC1xKHYXLGLICuD/QJ/zO
KmO9QwU68YkiD7z1cAqgFldhYckvXP/QVFo8W/74qG2qOsf8mOZK7rgHH1Qp3aYE
dyFRAgRko08erF2XeNWuylrJ8QqOZEYdLekcTmISgFiGOUk24ElKMwlY4JpYzdKz
AZvgwkhbFqcRAf8S66qFbSf3QfJT2e+rrGKr+101qqGGMJaIM4aQrSV+w+SX2r3U
grCsjxs7cwykBclUgMBsDR5DS90Ok3ee3QtliC7YKAqPSYmNI8JfLMmgxzDy3+yP
pQ0vR5jf0ZrrqiaorFpxlo3WaXhpeeZXn/WzQ4RKjWFnABcU9gxOAEGoh1eXjDle
QWCkvJu4MX9DOqLyVJjxSufmVva5a8HIOdgYQYuKBYPlEH0Wu1pVGw8WTJUXmwzp
nTlfHAJu/B1CAeuOrDFvv6OgEIdADq5PQXElO500VY0u39aYgr5W8QDeoEv0KxYS
hfN3OYutCkolr5O78HcKs+uk5PT8+XZVhlDOidHMbCAdEBZyFe53Ynz+AfQBsXTi
7ZrCIgEKv2TM8ysPg2St2EwaITENpSMrCywoe2VRmJ8kY9q0lvLaiejpbrwGmByQ
3BDupnYvUfwow/8imoLZthZPNHfZI78awPi0C1AynvK1qlcrnkMDHk9wCNv9hs2O
j5R8+HK8Ay+fkqTGk9VDNArfP85RZqCx8kAN9BRvUDeoiMpAK0wdEKFXClgEWXW6
IpeKp95DhEo6xAWoC17jg2qfPL2CDBx7qfpHUp9AiElcQlChDpI9TCMH9ML7iC2K
4PfRNAevENmYdqCfoe4GbDZ0eGy+grISeZg+VqtlmOg2td5VPqnrH3r7FkloGIp1
wCwcXbxm2rIw3umPSu5G4Ke7rElSppZmdWsrLi9yT4JzN+ipouqEo/16E2tbUHu4
hdjvfA0GEzJ7JlGuK5RWsiqZoCHVBe12MSC7Yw/46uYPAw2BPlOjBXQiDuclA9LT
AFA4cji1dHI8nO1/rfVaeZExTRDEcoZHNt6gbttLYFa/uDBXThxh1tSuW/SqPVL+
9jhKa2fVqcoDqXS56XL0nfQfH88BrEQmxpS6hxmWWLEWodp/OkeDHaT0lwrayw9x
3nIO848RQ9MSGRFpRUEZJzj0CdNgS+/ubLuA9stOHGlJyScfBs7XaJc0gk4r9S+d
ylWF+7B0xBeCete8Ok8m5yCduPB5OpbWKubJgpv9EmbyvoupJo2HXZBlJUNIDguB
vf0bYt5vKa6ID1HdwduuAPWrhXOwDUIHhwPd8x9MXs4x+X13r71m5kvgfkM18CDT
0B5EcNDHQOXEeGl5UMmkP2qdKZLCMkB6p6NRgRusgXDJOoqdAUg2DrCvF80ZGqOM
TRSTIIzn4fXbkNLAOiWF5i0iEiohmg87YPBLpGpSeDk5mJx8TVGZ6sFH+p0fLvNo
JuUbVdrgAE/thrBfkGLNklUoP6NCRgsoWgq36Yx+teWo0hkokMcspIPxIzAdKsUN
sp228JtIcyOgqK4TzOet29l2t6eDr9kwqkEk+Fs3UAKIjlbCqZf3p7oE0WA6j71s
yE2zpNQpksKRowa4y0Zp93AkzSaPgvRovfpcOwZ7oXfSvnHPUQuKN1paPJrf9vbS
kgDom58W8PQ84F0Yj6jb5xrTfoyzQCUp9rEam7YjZTxFKY0fVc5xvWRMtcciL4PX
+2OnBh/oVZz/Zitk9dqU6UwCfh+PdYbzsC2WDedhy5FGg5id+3wU1iU/2AKeYV1s
i7QMLvTRy1TMMmcpYcMW96VcXMsc4ApqAf3JZnscUXfe0DIofE7hMSSCvuerNn3U
QLsj3KHu6M6e8AXDGNRHkWTMqfqikbsgz92m9u57nd7gFbNrCGot50m3ANBnel/B
vkzwtHyY5sdownDdj45NuiWitTgHoFnRBWz07FG8JyieeZkElMCe/ZGVsRygGzEv
fYe/sQunhLgHGhDISreB7P7P3WPvEgQh1Tu/LWDAO2OycZiZohOjsS0Ld2PW3pKm
Psnt/N9az5h//SfAKq6jsP+7HYQDhjAaRst5JtbIIgu4x3mjwMfPA5s8hqjrhYNR
4KnWccShGsUlLNMwl6Uygvuv2npqOa1fN64mQvM7IUIoWIxuNOzxWEhs1VzgLQKg
TE8YByPDwTXZVvbh5Dow7x97lc515eQEOP3XEmmsSx/xQyDk/bLZMI++VS/8Nu5G
NDn7JcgNBOTRgc5WaHGcqVr2GYO96j6jxsi5fRqAb4lVFX3Qhwp5yxu3W953bbe0
2u8A+KGwtCl4tE9rR4GqQdxy6G5P+804wZV5dJNIlLpTsUoKqAB5TJ2D3PGJ1Yk/
41zlHqdViUsT/ZvDgx6mnvuRz7xFn0uncouWDttPKoMSQNymhz3vgnaGRtr7gs/f
glRxpKuREuDfSW9OKm6bJ545OXLCo+08imvRGbm32fkBG3h9596Wd+4HaL8nYk0n
XwS7Bm87AndUN0j9/Mw1sSobr+ufxUbDE8A1D318xvb4zt9ggVidrMLadhV+AeHL
tI6CZlT0GJsbAIZPtzJOfIBsM4NpjOKqysCllGCM80k3zNVW9BO6qHhQ0zbLkIko
EhgWVhAfEJKwfmlGWW43NQsXOEra3slm9gj2LPoNMfOQxpnD0cE3w7QrDrjC6bnL
Rt02XKCWQyIvOUmti8ZQyIBIOl0Xi2f8RyonOvRAXR/ztuAG9rlGL7CvaoLubxxx
/26Zs8kCXKecMsyinUYskFDApn/yhzgBQYxql0t4p4vSVPuBxHiQfKEsotb76qZG
lX5gWDoR5M0iaPGKtE09h09ipJUw+Tx43IbnaLOJUf1IVAJ6g9N3glfqHder0iIf
281C4Vmv5ftkVp+8FdSFSLYbgf3+ihLo6t6YAg774NTos0aablqUgmYppKNoTrYM
RRxM+7ve3foLUPgik9jSslOmbFfcM8Exk+2BUXPwxDiYz/5oq55YIOwO8K+UM0Uc
XaSfmsNlrez9kDWsAGAXvuuq8cPlzDjwMmgh2QUtEL+D5duWhk0pXPTRLVkklzeS
RcGAC1r4hLcihYwUrF04fjgLo+z0RDOcNjNf9ZGV/JduZgy6oa8XF7tMrQZGZvEx
8FnfpN+LBL0LlhMF41eH1ltilMg4C2G1kjurjAff3uUB+QwAEQ2PpaULR8ljkuDC
wvPvpqxc7Dxu/JYZ4DbmlIw0hOiD9jQrVBUEL4zYD+RYLUSBRSstgO4N2PgNUs9U
QyyvXxUUJ8adAHG28l2tsZuopMgVRF4ecBhqdhS+4b5o/EBPKq6rQHDFod/mhLj+
P4QvOEJH6bwjvkQOF1v0Fvtt/6351Ma+Uu5LPGQDHmiIyfRP/eumZuq6y0iZzbmW
EWxF1DzPcKaBwGkL8PovVitvS+Fn8W+D3gm6ePIqmiEfqD08ITxEwi2Ry1oIzGwE
8NzmSxiIS2Fuc41ngmracSuWx27oGR4eBSPG6G/6Bdlci7cNjTpDTFqg2bHLptNW
UPzlHNbvprl8jP4eNITkY8uCtGKdNbVzMOjZsvOufzB7xvbqZGqgl8zWWILWDzmh
Hs/6yo3EpYoSLOnhUA5mRF9aMju1dTMiNgzt2QNoQV7yBZb/g643VAOSRNzMfHLr
T79RdbV25rgggITQaVHa6hfW05hvWJ6WhxV0U6yaTbv43pify2VbjH2AkTQ1mJ4E
Wsv+xA2WmjyTrYpcfkDbDJCR5FwtcglSnkjRiL3P2v0Dea2/9PLNGfLI7y+Y3L0M
PZ07umUwUHMc1gvacMS61YtV/c7r25X6pZCyQdxpapqKUWHcpPMVvIXoIN2WMGSw
Yav61gFue96gDZN9sx2cfERESFmCgsH5SKrJ9qsgnHUf0TyB60WpZL5lLp0+t96X
i/XTPgC8BhQnKnNtVHvnsa627WhXjFCDWQpDhLO2wsTyufORFU7jS7nWTo6htafY
KVVGtVlC/wyhkXVnQS5R2e8tLgiVgPbd5FhDpAHScAJgD30W5+8F6UtdZRxAD7+H
4zrsjyMnclwboy6EchPbo7QFNg2f/V+8o1qRJZ4iex5nloDZHeflWTE+cFDelCRA
OX5Ic53s1mgnTcKfJHq3/XIyj7IyGE0u/cbgul6J3MBAYxtR9fbqG1PsqdeG20Yn
/dKoQOn4jpHq5wFvOFI91+AZ38cr4eePkDcT5FxPqWARMGv3ZqO2xbFQUaOKZ/ok
+fM50HAFYpBIQMb2y/s5g2EmC46H5e86UjtNGY7DiGJ8KxHD1DWFQb+nEv+5x+M+
Duf5eujvQgjTSpg8xpSk2WSbVOCD45ujZ5DAXqbLP6Sk3EaNzOyxLMUrk12hIZh4
9pB8KxnBjlQNBQNjYb2mEBSNhkFjPR9Be8HMfWdSMw+ao4SEipEEzKRxnoRxlSG2
lDcq6TazR5j/4RmAWDL272en9ok4Tf04V/23DOF2/451Nzh21BF8QXRlbwoJ0oCg
Ih5CB6IoYhi6q1arcnk7ZsxmNZ1d/RZjIsotpWsmPwcSHQHFB2TnJ7U9eFUD05M/
jp7UwlFph99jVcJySrik3zqOxdHe6r/1FNcNl7vTlHIbKTLie0nPZKHCxEyGbdJx
4pgArViEYn2SGv+CO4KB76LXBFFMAldCn6vQQBQo1Dc5pCWYLoMjnNFkrxMNK6VX
FK/2AE5pRDATiRaPmHeQGw/xLfybfVwtYCZO48+RW6zPOv42lfkfwIE2DrflLEFv
Qvnwwo54HSL8jN0JrKRKJ5f9RgseV3IZurHhx6nF5a/H3lo5aBLtrBskqs3RH0GK
7RK82cxLMFiexwaAAl7dre+yrr2GWGz+wyFqmDWq99uUVmV+X8AlA6Pw1fttLKaa
8kJdYynrHv+kK2AiRvOEa++g2EXzCAzxwMcRtj29SCafU92SJTsZ40CrW0fY0VYg
vwWwecZebg2k4EaO8DMPSIED7LvNY9vkRQ9IvrrPM3BEKsD1VJEgu04vLXkF0xly
ngRfk3lsPeUi74HZaQ2JPeZOvKDNfJjbNM3+BullmKvaSmO44HcqMUAI7UKonk92
dU/xx8f8JVPq1xe14ZZTyI8y+rbQX3k9lsGXShI2OHPoHnD/5z+LQBWlFYtlNhbZ
MSrtnMiNP5zZRsFVYnS0o4RjPNDLBGShGz7Qx8U4ne34EAFo+7h/QPH/FyINBSzX
XWLKysGhlf9bObB4l6A0HgmY/spsw4x5VKj5Srrxgr4zfvUl8tN3T/yPjhr4IdnB
IDVTO9vUrBR4jmbo+Yr3acq3EtokKUdLRf7ZSeaxp2tniJmV8Uk4xY2SYVCvucBS
8MkcsS2q9w5JDJHc53D7EFFq5gdnmgDNUUrn/iPRE06yAF5RoiP2DB6SMEmhSmWb
iGGwbOUdMH7BZ0QVnlFsz4yb1moBXEO15GPqY4WLtApvRlLJftDviQ32qNbKzeYU
j8ZQ78MqbG5v0WC9SIgiAPs6RogPYTiBB60WWnbISOJpFpC26OtiHMJJfZPfWugc
Bhhe8+VmDkW2zvTEtm5RYZIebcpgwPjJ/lSRDYY3R0YW68PiVETKNJRQwh8tkdov
e/ZLQH9NbtNN7plWCiMJUR+1O7eOOXASEhHZLObeZx5tEkecoqu7vlm3JscEIaEx
CkcGqLzHOnea2qte1R50il1vBcrnHZxrsw543cTJt5eNrRFOTwQePf8GPxDxoFFT
rrwasuo4+iqDV/VA6SMuCmz3NFvEEn4G3JUCCbPQUvc5zvbVjDGjC8Q7X9P+rabO
te9/33t6Gr0znIlLjNsv/UgbEr2Rk+/IU/+K8FKQ4eEwpAAVXGZhEPd9CK16M0iU
Mtyrfo3bP7/Uw93DNsSKOPK9u1QuolvD6VURk54Wb+DiCpg5I+YC/zJA1cTALWWV
4Rh+ejPuZK7m1LUwFRxgfnyD31EV4j4M1hdYGuTeIfOYwec+DB5eHn1zSZ7Y2deG
FbPCLB32J3EQpe8SWXqMpkwWlgeklt5NfRizk4Kc3gDyxtrZ2VMMnOVeUWvTb+7S
ZdlPPs5Fw09mkcEKpKe/Ev1CG853fmqeZCJ6X6kB6kxPvdijx1yKT0/3roAjZfuM
kNaViW1tfHUSclHTXAVTC7gH8u9kQkxj5mvM+GpuklnWFBGtRVa4nH9JaAuRThjx
8zDNuog59/qlg+u0YuuXL2PP33oaCxzVlnV17ynfE1IdVK+ueDM9p6aheQMAAw9n
IxD+GecUgEoWdjQYt//cCgr3/6f9tdlVuMYpZuBLfJdEY82BnnaHi8QlGsftm5Ve
65TQcfk4okHdvjdTGp5oOxKctiR14ITuM6TLFIUlqv8gxaosN8Mu3tG9qynzbdsM
mCC+cZR9bv2KYeahHujlJHeKekEuYJcNChQu5uNvv+ewlkhvlJ3SfZrLHcnF1b4K
beN5/oHo1Ld/JVkuAMExsagwkH6eerXaCy0+P8majLnMrANyWNRkSYmmNgI8Xv/6
MOjYMyEtpe7xyQmJYFqO0qCkKic0+MF35XY4LWiEYcVc3IKf4mlnHbrRb7ojXOrp
YQ6CmXfcify/ihBZJ5eWYJqtz1HKGCRVvYejjrAnl2pQcOuB+9eEqyiSQcXdGcGO
gBPrV+Mty4kZe7B7EYEV1MkB8uEDXo5Pm3V0aj/qKNsGu+nR5yA1fYjoxl2DLN0z
vRoPVw+HQ/FyJJdL63dx5gAjMfcKeQxw8fqxMXusMBf0IJxa/GGy8+k9a+tLeYl+
njcylP7i3zT9fBkO1VgMedY4ohYzRb1oDFkZ9SRB8NZvmHCg91h5BrzZdks8HRU8
HIgtiRRaFPRPiTZ/hDfWybn58DnQEiqwuyRBzBctLbhmOPjfZVYIK4fuxc1q9Cqw
p29dvc+h+1J0N1T8EJeyrPy/rjuoqgxUB/Er3CP0o1D+YHOcgSGPKzeF/KtfFCh/
RuwWcqksuN0pAiyuqUZ6nUJzR3r8jnw6LgBFqxjjydwCrkbIvOyk2N3zG9PQt+5s
TWgmAEk03pwRAQ9/dI2lzfbsiBr/79RbxGxIFdkbOQzI+udA1+Q+l2GmsyRFklph
aIPA/8LRqeIA75kpy9n9r/QSE26wzOYClB6N4be5I3kCVmWOkATcdfEcic8ayU2q
m+9HyhS5iYy9xXHwQxWEnzUbyRL/L+2xYEXcg/uQLbj+5Nl87d3ahcu5cQOkJuL0
fdS8JCnBKT/IaXPCcgOY8yITzIpuCUAYLuPJk6/8ux6BR+IxZGTOlT6wQKD7djUP
nVxpeSa5X1W9CdzugNJ8AlO9X1f8mABvipRnJ4O80KdcW5hH7epz47Oat3Q116E4
7lryQtyokTZ9c8NqEohHFXFY72Ec4wkATqXpbJsq0Yubc1izG+IqHhethNeFZulf
7LGEwV0+HIqpHjYZXKgPS0dpedia50SAdnxq/XO4QqI699K1o0q62m6ho8+rGniV
gAsfQnXDCw4EN27xdPI2b8Fld+grQeo1bRUZtJ9n/mG+beafPtlbbMOQGF2z5eXn
bjZ7F+whcOp64sKnvmB1KLacjjNeRFfm85qVJdNi1u6C3KKAVLCxi+QNR09Aggd8
qo7QMS52xLaZV2ym9l8pUVhyb5lF0ct8w3q0EkygszmeRU5AHpz0WjHuqVjNJY2E
PS7gmleAYZvWTDZnsKRDLGyEyCcWEtCUcb8dXOJttn4ST0ubJk5xas+AIZirhteq
VpQin+fBAGosx/rwxiuBokGVhFVhY8toilChnrIZvzQ4BOz/OhGcY/LN0NYB9t16
0g6yI7mGOA+KVLIGD4WQ6+u/8kw7hL0e377asrbND5fNnaFrpVjyUXl04hguKUrC
NlcJfSpf+dAKB+5/3GEoEYbpCovSxnDcGfPNHt/zuw/R2shjo2kjecd9Isz0K66Y
chwdzE95lPvSSMAq64teVti09L9pjyWO2+/dV7M+Ff7DJJpYEJoqOB+840pyq+y+
XcmjJZlr/caBMev6GjpcAmG/6fzU6gEZAq97LSJIyQZUo4Zv+GkC25YNdT8X8bsm
wUdkHmFTU+ul13CQcul7jDCAyvxTgyqDdHFUU1Ts1hm39d9ISHhQaZ5FfKUg0qOz
Z7ljb5Dv2HgSIhcvpHxhXvB8V1t8StILLWrS+vSsG4SbQ8r+EYVN6KQhllUHj6Cp
SnT9TxjEH91HoKfhvhHXMYhiihPqfKPmCmLZ66DIzp8W1dL3cgDKTDGxrSMKtl2E
7d9jx2WBdH4MzrNC7bC1D0/01QXrt4jHmZJEwg4Gx3Vb7zlYn++0D3+jI9AEoOk0
bq5FytMz9vPnqZruzql8Zhk+WIqAQkbT3QAQ4BrcMFryT4Su+y0s9KLF5KCDwxR4
jcnwcv7iXQaYi4eziWbE22SPXLZL5eNuC3sLte2JnTIKAVfhNwpWZNXPeL4Lx/J4
7Q24n9YNwHHfpill2s4iNsmc3o/q5/CtkUwpMempIxf7gsZFJgtknH5F4gBffLIj
M1xuA4W7cg/dtAfsMyEInhKy/RYukAKcje8Sn8hATc0AeNJ+w84PlL97q7R2QrT2
u3SdCDcvKnXuheoN+4nghMD/fOgUlT0ZfH9jy43Pf4VLHkShfQQi/BK1DXT6QnUK
N08bss83qASWrVvoH4H9ZMJr/rny3y1ohBqz678tuWsuej8ZaJpjLZlPpz9KstKq
h2vUJGR3o5UIK88vvrmqBSfxAewF/1UPYtpgn0sWpeJNwNnDBxI6gsBJgaC+2QkJ
oO4HKk6k5XHPUE0iXa4+rh4qdzRSmTpY5xZHdzPZyI30CCr572yOpQ/PZe6fcCA8
Msm2SdVgIORDsSoN7fFj+fJszww9ZvOryMUK7qm3QMMMYwwDVSWIWaHc5vVVvGEl
wFPP5QFAypDamZBo0wqQuL29ZRlUf6BRZQKtcHbTe70jNz2G4qOPAdddqEaerKr2
fhzsFBOJD6mDH5yZ+PeWYnxN4L5c5s8jtoBYodJSSTjSSmb4rRGKM9Hv2JZ1CW3M
bSX9JJmZsQuzkbKV5avzjZJeoW8zmNWnMKkPatETrt2dVrafEPWYG8fu2XWAOYfX
zYS8B+ngyVlR5cReIRLQwZh8EAtgLn5j6m5/OjKHcGkIH/+V6Kv5E3rCR/FsPi5m
kB7/ov1b7NtOe4YvPcACSUz3Hr1v2FOU0sznAGf3aAAWh6Jb5D1IBzC3VZ457Seq
GO5NvxIpdFw0Oel8l3uU6rUt/46JpBl39L9fW77Fl/Co+EZsNn8yQps+hTXo0fUE
XwAEa8laDSu3nfKY6bPYnMTcbXAJKI9SF1shSfNfBoD72D3Ft+jMdcpR452hgYrI
/PKtaT7M8gItrDCoAa7O+cI5e1uaiQxnvLbkzdCpgo1rA5WLU1Qfi+b+E80RBCZY
vvCZ9n8ZsRrMfrOK+knEUp7MNbc7DPVvhuh6XRnWyF81JjWXRARVh6P7xBBoHDls
M/BpQ7d0ihyGjw5qKTCqurB6in49AXfFuYEcN8GEHuqPRbbtv6lu5WfmpxuJMiQv
df4vB2ejUz793vmRpWTPqF2574kjw1b3txoFM4PAEu7Cl5pfDZD5lbDisSq7IOrY
5CEhyJjBIvEj59ZJdWF1Aws+aKRr31L0AbiTbtLm0VOFbTcSMZxEiZO0IQ9NYyUw
Ho0cSttZnRgDaBaJxpzwfPVg0gWMC+7MihEjfEx+3EGauclJS1JaOyiPQ3ZY0SZ4
YMrMDreReRWv1Z0YYZLFDfKNPIyhpwF9Q330Y5nLvGwS00/jOC30mXH+xo3zirM5
+eMrfPN0LXhdCLpdXk/4hVBUwuFRlTLNb6Aw9ZxFcTftsV/vrbuHd/tdllN0gwsn
s3h7G1sYLlI6lJfJUzZE0xttGMuxjCJi5usQLn+N2HUva9M1BX4wPfkU9ZrOg581
ZQS5OQWAl8RZuwP4xd1LxNBQcDnhRHkFDJOmA2ViO/9i+CBnY/Ye1tBC/8Ps/AG2
p62EUikrfHRq/ma5aPi1TGIIGZmx7fsfsVrYDudHm5AUNINV6tJmaK0EsajCknXi
y9A5gju6prdJVeKSZlkpuHWK7yQyUCTYpWUwlSLrMc5wdmWSeB2SlZM7P0JYX8TL
OMG0d3Cu8IeukbknAIh67S5E63zCV+VOezT8rgZOfDAnuKJEF31ECSIw+RplVSmV
k6ew5oiQ6MSyhbzNHt63RQrI/Jva+iALEy6pEgaUTrsSwSlDLkyXY0CHsh+BzTCH
COK+4z59kxOmJD3h0ySo08Z3weuXhI4UNAt6ax2yDU0HiWqKww5jBR4bIwGirQSC
S9B6d0rJXWM9t0I9atXu93Ba2tzAijhHUNiLcmiwaHXuKg2vESn3EXE22bPrnan6
l2u4Ff8X9FSo0tMI6DRez7FClFI3is3s01XOnROE9rd92gDvOwoLyfjM4di4gdEc
MEbzRrLJ0jEkmbCQtM3MWNhh/YnmzComjTBwQV67T38/lhvzxCkOmCliIaZmfrsn
HGRif+x80cSbAs2Yv4g0/r1uWgux7ysFtyUqXaYJlkFC+jxRcxueIeOdBHWj07Bq
EP3bw4LRKgCLnQZbpLBeXbQDQNuAjPSGwgh7Jqh03S0s20xhYXkIZF8H4o0mOpqH
OvnpTAJDlnVvBJQeoSSvEVEuoVxnW+ZICfnhSusxtER+jL9shwGcftHCj+v4/sEu
9J8O/u45te94lp18DvvBzexBJOLlBoSAWMsQz3DXTABFiQ149QwscIdu4JmhUa8q
walbdUDULEjxM9YZv/98upzIN8ZdFq2DSCKqI4kABNhR11XxxO5W+SD0uaV9h7tt
jjnV6XV7zK9RCsyVzQaPiki6yCf4E6jMzEFV4VISFOXlYi2I+YGZ8BU72wiPEK6b
gT5kCEjwjOM9Euw+KPchqxVp+WEo5JapOuP3NsmmjkRDevsfVGvwpYEgC9z1oBfr
7VrN0r6mucIbXzWb/zB6EiEkNaWQZtxKHBIwgOfJgw5OCLNODfSVyT/0KGE9cUPS
aUs0nyInoRNt3bQDFF2WXm8WU6fy+ix7xyiJTPhGJFwPR5tEW0JvMZgIys78dD0b
g4jTaEmrvzoxE5sLO6Ce8tmMmNqkjBFp4UQw11tmleCYSi6Zn5QFE1Onh176j+Sf
stzn7nXqw3J1Rjx+vuY3DuT+PYE47pKIW+tlMshjERoVZ0cOXzRVNy5q3yymEr9F
1wnF7gzUuY5SHQpAcS1rP4u5/cSJM0yI22dwoSoHmwum2cRGOTeFehT4Nh5w94zV
rdgJRPcubfRGsf87nVpVegxcTQQPwwFcJWGm+UOZFOoEgoKmowN9kgl2JfY0m1pT
4In07uGbCHmy8IZQjIH4Zn3T2QT7pc6hNMxRWKhbqid3vm+EhL5O/KklCVHP8Tao
UJhB6pklSXpUNieTkbi/F4tNmKq4GOpu3dv4vQW5f05Edsm1YVDjZ4HgfiTBdXAE
otp/UVAr9x/4/4rUMLAFWTCf1m+ufREO9pSrWM5bLR8fXO9uR5ckpMhBFtlWEhuM
ftYaUlSi9pPy1ittZsHPiLjsgBBUc8Fo9HJpfXQOrkG3O74wNrzP8XBVO5iPLzv8
hrVmfvOb7qPwOAfX3b8K0FWrYSfAP55eiauvj+ISD4t/yZQMowKJ+ncjzUCZ7Y2q
lvZdWrjSrmxBzDjdVg6CRYy1M1YaKYyU2eHBXpWX7S/A+LS38XvFNIOsSsS7Uqna
TsZKrUhfYkdlXnGXriGZm7CT/ABz/tajB3wkC7cfY69XocmFA1WfaqgZtRUYUxeg
cLHTMOKPbV83tN/FUIwr2VGI+hgezVN77yJxmeBg/toLLPwin+myCkRzkOepLhU4
ztspR8l80fiYhKvSQhrFhNmDJMhdxfyIiw9ca1r5X7/QifPSZoRZ35H72RbdZZRt
w3ifAKditaJS0N5KDFs3r0DKaI4nPq5KHsoBPK+M3wbg2dNR6jSpe4Br3uzT5jcl
8r8TetXyrfpEJFrjz1MCG7tR+MlHN8lmt4NQoSWjSos5+BWdSp6YMkigJiv13K8B
cjU6+ioy1Va8ByRwE26/QuhWoMM9042oKBnBKrKACdcFoLAyDzLtLI7gxlK40Lvh
gK/AnWVGvsNurOYpfWE01Sm0BZRW3XB0uwoavWp09+jEEcpc3eOzA6qDryDhsYIP
FMxXDvm81NQonHGJ6gZS9wfJtRV+SyPOQekZ9fA1JEW6/Fo6Jpnu0sZiMMp0B37V
zrxkNIVFuB1aI6m534W/KUTCk4il7LxMIV53PSVDSLsLffiJs0eALlHsRdbTiJpj
a09ipYzcgOv1jJKdziuOmKZ3E//4kyVA2Yo70mQW1jXycWeoxLSN+L60Hdv8SYRg
06QlLLURIApbx5Wta7/cJtu4dylSht37F+a5A116hK/mUanswtGCXW36oWOsvC+2
PuryVQBS4upQN3Bu658tTmpiVnaSdJvv3OKnc6O11RvZQBIDU/nsL3eaYMyiAvat
LlPXgXgOg+O3YsIG9sceAI2BT4pUC/nghaiNfVZMnMV87j01acilyF4r7L5yttVl
2pe9q2StVrE17I8HIJZmfyahxA8WN5CSVs9iOM9dYHBDVGi1bNRKmnkjMm36ubKz
7TVL/AaOBk99ZT8EfXBnw/Ejobanuk9ZDHnjjVZoraacGpgPAoG1GeUJY37VUiMW
cW75kFZ7XDGDzooXzURJAz6sLnLYJ9+T3ij4titCpjlfzlMlcl8tup7NYXatyACh
sq/W9987XV87xbf3kcZRD8XX5PkI3v6676A82n+WrxXvPjuBQv1+AsBuP/d+h/QY
XMRN9GvB8cvl1cGpVFq9MVxuFQHn+5GTpXWwdxVGHEeHGRRJ4b1an9kKTxtbRIIJ
QDEscvkOHURDus8nIqRPPokq5hRYdX72aErU0crqqNAe6uWD8fo5YXScPpCGHl2+
ZSznZobMu0gGt/ePE2SNwyodMleUt6rzeEndV0yP5F+GHqd7CId4yzTiSq3sQ8kQ
wtiy5pLSzPaI5GFPVggFjYrFv6mWb2s9HVfV7NSZevo+9MEGjCacsFYlX7qnJOwN
WJKoyA5cDapzrfDVoVE1BDmeKNKZIsRCYylwm7vfCw5xY0QjHED5DMh1uSakZetk
gHbDIr4BivLzc2i1XpMguZxVS5sVBJUbwVtjB16bfR7LWohaB17EYoKofpWlMeR+
9/Amkh9p2GH0LKlFYJmhtFafe9jzTL5lTuv9LxNkgcIa7BObvvLE54PnlUY1cbh/
pxV/qfgojDhRu1QxwMVkQYsvy5tIq5s2pLXBnL/IY6F3GqtzE4pfn5H+HqSnm32z
0pJ5mcNLPmWGE8ho9fv5+2j6k6jvsWMlC4yBWxMQUivrG83BD9o/B510Mq4ouh5f
Luu13XmaDHwR2ULQamcSXADDU3AHJxOjVfIX+EoB4oeZ4Eu8OZfPQUMd10fkay1V
ydPc+nOuV3swj+wfAPDSa2TD1gEMFVUlknBEMupGZ2YmjIZkGUspW8wBtIdYHfTI
KG2XqQFpAUhUcqeHXvCy/wiZy10aZW66qZpw4rFiaPweD4ruRHWnBihDu+jyuvTc
XVGbU7pv3KO428zrnRWDeV2mmvpOuvTkHwVo4QOvkZYRIiYE2PgZq3Us4SUbkjLk
Zr03ZH5myYUaglmeyoc33mvwiE9InmzJoGRJoZBViwGmsXvpzDT598PDQrfWw/r1
87PJshZCA7v4y7XnTjwREkQap9eJ7V+H0we548qQpyBzos6kYoB6VdVmGcTDsilK
5Ihd/CtXNe6O1iOZ5pWWw/xz/WcMcIpeztcYS7/06XF27NYxdZlJcSt+POQraK5b
FUUZKfi6zRsMxzggNEnIE2ANU3Z4XNcN9Od1QoZTCOhqTg7Xg/KmUSNBZw0e/+kS
3CctuzR8qXJ12fdTMdLhd2LAESCP5BZC74pva8oD+am7noBgxl5C3xWUL96mah7q
g/Bw3kqVdVhaZXDy17SO8uz2k9TcE95YwOC9ZII7Wl99vLwzxbuEoGLppxPu4+wg
+yuh0VadA8/lkR8QIw5JOHP4Ug9i++GmuAkzwKpaxH+Xwp4E2QIKjTN7orhnKog+
6vMjeelpZjf1NVm8ut5WyYvS0NpsicEjWCiWDjwDenEjkFhao88WW1y4W86aXENW
Ui29fzw/KZNfqas2+SzEoYsqgTZgngE6f++ogiUAZtwOSk2AwK3FkANSmfNqkoPO
n5V7H3JuYnK3EYNncumeZad+u/MxiY7ZGAeq9k+F1wScSGCiTFyqj1TuwY4s2O0o
fTMgfm7vTKnU5WoOpIAMDJBaaGI8kqC+wvp8AYecKLoveSg9tXdwvEE1IQzeoo/4
xvyO/InjrSUM3eigsSbP+5qpPQ+93fqASGjgpujkw1MiftQK11NP/z3ERj7z6hty
SV+dJd9qDRfXDOhByn3FhmMlWsVDk7uSf40uFXM/W3Ak8IZi6k2hQZiM5iutBIJ7
65vl2N26CbzTV1bVwiJA6IsGxORSZ/MDIFu72a7fCXsI3usM3RrZBbZCRM7+h3JM
uackBsc/bgW72j4gQ0d/4ZNKCp2p62rZ5fHjzPUowTDI/g5HRiDBAyo0anxlWhhq
nw0kAygkFBFCgNHkjOBm32JlGKVmUQKGzIujyCVP4lkbb9WGP8amv6r6OHUPYmF6
/TKm9GeM4KKIcb58N+h0JhlYPyGljFqf1PauIGb2KwfgQ8eWusKjsKLZdtKNGzM4
ejIUglzBzDB6/fqJqsZ5G5/mOQLmj+yNvn1VT88r5f8bjX/1oMgx/NzjYGW51wZc
fj/edU/sIVeaxFfXcCVVOqNF4StqHY/2IP28QYtcS1Bgd63Gx5rOea+YUythEEPw
Ddolfwx/eqxODlgyhWDVrMC4ohPGGDhwVaG7i5t7KgISq7qrKYbIqL1+AxWAoQTM
mfbVjmvHvSEoV4VXlsoWNcMe4d75WN2ONtz50jXFkmAjE3nLphoJh2fbt1RZE9S1
wibM6IfvdqxudJq/lcn/ly/b4n+BqxoDhm7eBQYMbuEPCunh1KNAWVulHsRDjCcy
fCYrBp/RaIrzEqqOXWEcKp7X8BrVpmVH7j9/9Y8b2jefy2edU9eLKF4Yk9e5+uy3
eYnxkc/8ZRjqDGJDNtQbJJCLpwCu40U2DtFnXhb/0OOBoF4U50CDGogPQYVbLXoG
iYoEmq1LCisk+V7rgkqSZ+NRB4yaGsXta1nx/iqhDze4p3Cu4wevmF1Dt4Wr5Ll3
KZaLu9Sh6CGhfPLqvwWWs3YJ/ZCRdcnHOeTTcCMyZqbDmL5c6Hbis0RcUqC7/PNI
EsrZDiy+xAZRnr/hUgkKniCeAWzQqz1o09FEdEk2fCSJyTVpGt5CNJlnTIioSjE7
LrBoArWLKSJuY8Xss34nanSIpQB26PBc3Vv012WL0zoRiDJ58Z36Iz4xnrT2/YIX
S36hF/sSYxqX+0kr6neGws4rVX7UWItC3zHJZ+bAEJNK6+1gvkomhZvk5RIiEu70
SEErcbLRq1sUeuUS7zwDerZvLt/VYBGk28gElSYNW+2UV+hn7AOcgDZK2Pp5f1Eg
vhZrSKKx/OEqri0N45UlPA20YZQ8WSU5Sd0iEjjt9ojCjgl7/+6v5hd9q/1ITo1a
n6Qsc3dZn1xYv8er/E8fY3Fz/ugtsJtGl22Uy7RHSDe0Bsb09AqsqesQxnUgzovr
pT9785QNVUy9Ee4aae3DdQIoqWrhqj8Y0kmY4ki6vzm31oWVvYkXGSYIrkIFRNH/
DgwYzi/bis6KN0PQM2WqwDntN+/7pwTciQaxm9ShIO8HSDUoaj9yLXWdQdhkCoRX
/IS0sedNG9U2zVHgye5LwOZnaMeeK3yWTjkxMMK7hqGCPlzd24RdpZ0WYO1N9ktH
HhWA7xOyuuzOFQHwfLw+hmmjf/VAKM8AywfyJopS0y9ce5leHVgDD+uppyk7Sruy
F2D8WoRIpIoyGZA0v/QdfofI2cnLOjhxZTafJ4sAcMbzP3w/sIPr4qCMrspMSbWQ
XhA3cFLIESTmP4/6Pyp/LrcXmziCaI81cUPmIB4VW7yRqVxBLNCFgH5QEh/41zBT
H2NM4u+DsnvvDfchXBLm3IL0i6nsZ4o2tD5T2IZK5+/hydl+iPJlZsHeH6vTgtP4
lK2AssaZsZouxBKVWsT/7VMCGDsIhbG34uuB2uXfi1Rooy/6eW7nAkkVadcRoRrT
T4iOJQa8r2dHR3WjHfNWXXcfWLH5rT4mLZOrOTrBp/SKyAyg5zFiA1Ebh+SPT4Wi
L7l80CkbKnW5trI7nd93ZaE5gbx1aphpRVh4uBZZH/rNt/e8+oJav6KCe9iF2bRm
gyYIN97GhBr7JZfXq4v8gs3s3xLIl4GSa/tWVvg55wTXAUbiF1OoNcdP40fVxfrb
jZT1SqqPsUFq1SSQOY4myqzIsLn1q3Q6F1gqJON75VpRQxl/qLDdpJOaRdi5CsRy
05Tgi/5ER8HVdfnZ0Q3PTRrYwK2xBSKwMW5ft9kvn2wupbbyhzDcvGlcvDixixOQ
SUTbWSBh4ASv834Tfm4rSnf+TSaoQ3VN5WOXacNT39wgXQdpNDCXavthS1Mer5N6
jJiX/8GwwWQD3ygi1gFbvKnb40VY2BElp1UeeoDgNSQZNYbyi986Jeu8C4Op1I6Z
vz5GQxuui/b+t3g+VmwkbByMXuUb6x4APmgX/54vlUkPelDzCV/RE79QC6Vbug45
7tnvjPKk/9BjvF2yNjlwDdsedrnc+OE8SGl9gyuyeUZm3UaQn1EqnzqLNtrDmrhs
ZsnAIqyYQuqm1cl8BqbNspTy5Ibhn0FZf9tHPI1/0oRiqXAJ7owwXK8zntCDCudl
ywyUd7VM35gnzp78H2aZuYRCZkYtfsPy0rCTR6uYI04aIauDukAnTFHZO8AHzq3/
oC49m7YPOX3rssv7CGk5wOmPo7UJJo5k2iNC7OKX6H+5Dx/cvzKdOG7Zl5hVa/6/
6tW8efNGeH7MfpvOmy5r96iNGyV8f3TM7b8qIITjXZSV82bvMKgyQPuolf03aYMW
vIGv0CQ3Zkb3XtO1Os/NI6iKeuBqsuUfQYSxSVXZ7YF94MBXIGyikQQQGSm1lhrh
yW22bGkLHCiHpuscZARu6j94KN1BshlCqjl7IgTIy/PZ5VDoCA+CqAWkpFTVHw0r
Cu+H+e0ZGFIvWN1pnF6YT+XVtTdyJ5Zf2T48qPCqxdT7PkAbegKxqqtlUixA4JnE
lh0nBrlx2MNty1ftAEoOAQDkgF4akLk2ChErLjhg3H0S7O18toybGhqbzuhNnaXk
KqcnGBwLwxeIKO83XUQ9U+YhHQAmL9CpkkV9YObsrDe9X7c9KrH8PSMM1TGaaRar
4GzA0sfm+bSsIJjzmeLTo40qnyytJkJSEGoRmza8HHenxPaUKp3FX2ewhdpqUjA3
hzpvinwnabCP0giUiQGMOPs8WPNfpxrGTqh/FVcyrdMcv/Vnt0BM15IQAyDr4jEg
utPkyV6q16R7fwG5FQj92fVcr6GN2Av0G7b4fE/Af+t0gm3IOVtNMaOfpVxzVZZM
vzaNgiZXMC7XTtYbUBThkmi1JwsGVSZqscSerOF78dHV4eTKeWDtQO0sy9kg6HzG
gaHJTaZ7nZDGcimHrMeRYETzL1VAR4JiTE1vInE/I62C1niybbKWRH/r0aHYANtN
wUxXh2st8/n7nyqALWgk3dUzgkTHmK5RyqCe4mDTUhl+3L5sJgT5X3lmY2Lw4pSu
CL+7UVkkZT3FmxDs7jt6epEbcuTyCaxr8ED6tkC+R3y6TYcB4r2m0ZOIouhKcUP6
0fi/OVwe48QFAjowcQLbPzLj0Q6wWoiO0rtSUziB+QT4Ju5KBZaHRy1QkZata7nr
ZNSLs9tjTcaiJwCxMhqxYfhG/iyjKahf2brp6HziHGk/DBHBFUdV+s4iUfNKoq+p
DvPhgp7cWORHujmJF/Id9cRSIh+R0bC+FKI4YQjxw3BbExsJk3SlFKJ3DImliMMa
CQW5p+AJ6qw9uWoDGylsIzL0OvDREVxJet8ohQDiWq5+TqJHdxbXesg1ah76vTOD
n/8bWUDMzwHRLe6mIF61Wh4t0cs38CvqQ+SGBa3YL0UW0kMi/QXSp7+cJCFaL/Ky
Cy2j61jujO15SI9TO2uLeG7V5f0/c1KtzsADK3XiqaeH+Uo4E+WYF9DcY+d6EKdN
ZRfuqlu3JeT0In5f0+CngyA4JiDF0HxOjSvW2YvPi4Fiziu7sUT1iH7dHW3n+vdW
dyeh9oBSaxcpPmRg67H8esW649eVd4mhY2fq4Bra19pxE6xxmOaixucNEqB9bnM5
q+r9hDLXREDnO2piGdsNcXhdVpbaxT/aiHevC4CG5kZFfQtWEHCYOt+5clsYonad
S9PLcP2KnzvMOtvoOV7pPkrcEop1k+zYpWU8rGgJm9uBNzzFI3Lz4FlNeVcPfxSx
4vPtWgizIHxePDQBhfdd/1O6QfUHh5rVRDCU8suvkjpto8NY/uerJ5xeJWTZ1LK9
tyGU9U6tjtbQxIwUQGDFkOP3eDq5wxj9TLMNnFswA0EEBM0uUhJyaaOVu7UFK/Pe
HCWqfg8moAW+UMH8CmJk2f5UZXLTDcnBJe8kWTeMoY3VOx96u+CBvagtK8n3yWhc
FUvK/iwdtWMZx5TXrOjNIo7alANJQnVYvDQY4b+gl+kl6/MLPSMQ8nefwx3c78zx
D45HGXeHz2eVn9Jq2IhZEjD/9RgXLxYMxlEpBozOSm0kXBYzz7te6T+36Cc/Dd3z
fSUiM9DckqokeSWWD1QnGnH/UujhzKM84LpVf6Qlg9ZWD/uvxMpKdPtiHpebUcuw
cO82DIdYbnAeXonN6gagIeZPLBQnL4VVAA8tmUMBL3K89AqWfYNtv11ViR51jW2e
AeFE9AfZDWkKWp0ZGTSkVDELoiZL0FzPGbVTJi+3choZpIrPdY7/xKFhT1f95ABo
hlZ3rQc4mYLDhWlZAlhn2x7dVlGVysa6lRRudNHq2tuRyDiJV6MQzGOARl3B6EDN
UlRp8EoviI7iw/M0b3gEVFJMb8rNGPucKHkAV+wG+rXgY1mAoo3+4yPMTtjP2onb
BQlre/za06nOKsssqaEgrdjbufF5FGEXElQAwX7outAN8lYEEQuRRjZAnqWiU2UQ
7xnJ4jv0M8VcHcU12/tu+ez4YHaWxRsNUWIJfaL6KKHCNYc9ST5HVnQmiB0EXiUP
O/mnW8Xrerb3qxg7IGdID1BaZd3zzeU0kAsyOaUkOYrvLHt8HVGTQf7ZiBm+Us7Q
M1yEzJhdsvi+ZqMMYnw1WIRa1mHinkgaCtv8D2jFsx8tNLoHugCPLhYVFhiwFrSK
meNQXFjkm8PpmdClXJxw1pOmrMpPMNx2THOdL85jGW2agLLOJaUSV7+ZnUahXPgx
tsmLwdBiunacgI36p8in2PA7h7TCYomOkR9yYZIBmgVrgXOMVmpfkmR65Qxkp46v
UnsTtRz9nKJPrG/q5suVtPWhkvyecHtP4cAl0ND+akHQtrpOlOfW2nDkmswqEKI5
C7H3BR/j3PF1MJOJV5og9bbDDFEllajqOIGf4SLhNayQU1nbmYw4ukxd0PPrkK6/
esDXmkYTsoHek4APRb6jWkLisD7+vEvfVG5mvNUsYpkHEm3WuK6h74dMJbJ28ivQ
DvXftm746dWMq5OJZ5aUoWJPdXGyAuy9xSaYDXFddHyId+MA5qi80omeiGsjDWBr
iSe8yQhdUkTexYfoL9nxgYUuYqqif1NqGj1EVAlSRh91T4GMThelJBW3InNRjBX2
DG7PFVT4o8Rh2DteLo1PzTKDG9G7AbGSLwFGjjyraskU+1pjGpqrjnGepAoqMJ6f
iqv8WJUfy6PpU0dw4sJxG010ufpjqPS1bm0d/gCNncR30ket+PIHGFV4b6TyFgHA
O4pRkJygoRi3jMsllZwK3402zWyb++BQv8dfviEXrE0ssqKglgeg1rC3seD3BjMC
FgTrV2WSwMGD4LVk2eDS8KJ0qH5qhS9KxtazdWk9C6GYWro+IdhlnlCSphFgWb/o
x1htBsgsZuhHw41Zg+bh4sRupqqYnhcRfcOIzEBzY+/KNEs7jT4qHYA6Qp6+dJ8E
7dDqyUDNGuRj7T79aghOz822p7Yous0xUFqcq1LGaqR1CvnZxLbjqUxxThQnt7Mk
/+VaWLt+RxSlLS4QbihQCKHbJOab2LdDHlvPzggHvEp7d5X96sBemvDZAHfrdPS1
rYUsi4YHzz5F4N5vrgPBixKak+SF7E1UIGuUGPoOWzf0PnU2x8Ak6jr58kFhdtH2
J1RuxLTsJGthGab+sbCOrWfcOS42QqQV2Sh8BH3vIUwFyKyjwfBUDt8Gwl7zEQIb
zjLaNIEAsh/RiJ71dotbdvxD1ddxHqhVek1tpTkHoQe86/my5Wku4FTfC+/GXJwS
3FPddTsreXRLcOgpXJfm0jdFvQyfnqKV1mlojhH09Oe9D90eHEWtb0YdGcytKNge
uZQGylUA9OwpWK6dZ5KeNywlY3X+3Kb06WktgniZSJ+yeBEtfPeH4/ia/qu94SGn
QFZTSzW5ol2EbsJoY1S/L9bw6IxL8gZMkjTlBbN4jkzJoyfKBvtx2BvpCNef0gdq
3grA/uaRSa4DKmgVekZLkTpmZUSnRViPuORt/EzE+moJvGO9V1hS1PS44CwYZ7u+
vHLRdiwmUb6YHgH73UnLieUCkxyyL5mpJVLf0eOmEfLnWOBvz0DgflhK6jDZfSrX
Lt62Ap/3gKnojah5qgm5Oy6FUCIe4WY1DQrVvaJ8IBiOZFttu7DYylVMIcnUNYq1
ANieZ1tS8/5FaBzMIBM99piPdYKTNvgArn1q3+fBfqvvoZoTKDhrklbAMVmpecan
NrzCApOksTNWAu4N9fX3rwAi6rYUmcQePX4I5VkiJ3NhCGthvGIFqgXWdEZQEqL4
k2Y15xcUTAuKQwUFBdyYFH42VZLFYbmtA1T2y8mmhUvOEK9YsUKp4IMdG82fGVfC
oXYqyM1ltkzy8G7tH5rzi+qvr5J76TQxVM1FhChLCochuql/1GTJHh9WsqgilsE2
fpub/CCyxF1uXLKjRaa/9GiQDmCeDwqjrIi5S8KoFYg5VsSFeSEG+7Cm5HeqqtpO
hkJMTo2iHWPvvddwXNv6TP9mUoF2GGZoNOINtl4aaCm95SVV+A3HKlEsqVb0/PZp
DMAOSjErL97VSGDi0j/h/icvRRJ/7F84IfpFL90WZ93r2qvTDud0vY2NqWe1kbPp
Db6/XXUQq0hJpZei/x5GeiUMNvkAWOK8lp6PtOpr2c0F9AG2qxXAVFNqlepnZ+sx
dCb7BFoEgPEzqV9tqdhZ/96VXKw5Z1+MW9S88YN8SN3C8tUL3T4rwSLc4IKx2PdV
0c3uPth2en0JQhY/SJkFpL3OHIqKXqdADqs1GhoI8/QyAVzLs7qi6wuktnYB4Axn
zP0ZgI9JUWGiHRcDTpjyesaZoQsyn2uJq1Hh0wHWJUjcO+01I1xztSBTTkmyveTE
c4HQbYVo5h72UPA+7AJ7+lfmnQWEgYKJAVRvyFMP+cswz5rHqB91hmncXkpgxGL4
ik3VjobtM7cwjQBbRpva2g3QTYzvq1cU5oTID7y5gFMK7QqbPzNsbcQzAlqRHfZ9
ClJ355W5tmqlPxfEM+g9OalF0bnsDnSFEfiwqN713tVGeioFJTH6zMp4ekcckC1l
iPedy/CXYjPRcmLF8v81IlOiCJIXnElWVfw/vNqdkgCIjtOpmkiZ250LYlmi5CQp
VV/r/sKuiv7Z8zaB/ETXCi3mPY4JwqFU/NNUKQ1YHlq+G5laa31jYsDXAcxKHOZT
yniEeqV+sZEtlWWO5r+8ipUkLXxMEQuu3u3gFYYaGFPmoIaEiJOXJzqXx0Ch2bES
m1eAZmJ4HFNIMlgNWwNAUEq4EmwH8nZMIYStmiYCAcycYpsiDr/UMc/ESzv3Ifnm
R30UpKYbnHBEW1FStsE/wJvsq2hOVOAFC2hSSmaw9J0okz026RA43IuKVJGD0c83
RSP9md9o1FTToDOD8LPZrY6zBiVtXLjcVJJ58ZiPLUU59gheJgdWtQLK4tJqHmU3
ihHZPb3BqRIrSuZ5XfPw/S4Jnq13a8Xtjf5uJn1/PyoL3vypmGgTb4di48WlvC7R
BjZzcAigu/A5OYZIQla2+ppGF96ae1PUm7Rw1ZEJJ9IHsVaspGUA5LENk2gX4B6K
qYw2c3xl0UCZP5kH+7C1ch1/BOGZGfGC9t0EToAzO5mSbvn5dSxKwTogodlKGGAa
BIMFQUblGCgpp+PWprm/9iaiazL4sWRDB9mPX63DG2DdinqTupmdkk5SdSMT6MrR
05bzeRYK0hIM012meeBLwa3Rt3hu/8kbRgV6HO8i0ZrNARXbzrKriImmTbU43rbi
KWARVuzX9g9XivwP03y29pxM/vLjndAauhBPLX3cdUjZvvanIE4Yf0/9fD76qubW
GXwTSBhWrwx3ukHFYBBJ9B+oP+n5PsUjHJuuTJKyGgxhlsvKBBN0fjfNdcrh8ZbS
eqG7G0c0LOnZFXvzZIeq8G6tWrhyh1bOp8jPish52LoSO3mmmP28ji15BqPmh3wg
EkAoA68bezj6AtEUOVHKz4trxBRuMI89CA2z/sAmRbBPCa3/xTROEu6kUR9Bq2o2
Z1nzYRz7LqQDp8uIBuQfcmJjuEFipXLTs7s7DELLSRRlm8nTYE4S+DKQxadxwae8
yZFQzh5pNJbWMl6JcX076ArSO1PtHHdqE8HI8jKmegz1WNpdjor3Txs9HDVrZqMR
Dmo7iOaRNxUrvJKA4shkjODf0BfLAqGmLRjj7zl6jWZVpDp2k9YNuJ5xbk3x7xhs
LeYSueoAMxjnoIZxWZ+3Jtd+uJyORFksnUOhoP0vBJOhac6KxzHWkmekTb66LbFd
XiOjNFiAYHyXCmARle0MkEF/k04dcx4HmFdhSg23VectMOZXUOSMsY4NQHqnAQn9
yw133BCcsM/bkYgJt21Jz9wrd0HWXD0D7mu2N3qQyxsrS4ewVGeVHO9noR2RDc1C
u3Y1gWYi5H+3WnSJdGKGd0rCEYvHr8epiMNneIoFbr7yDg5bBFl+Yx/At+gNiake
5ddIV+JxQpp2IyLAHmN7wO3C4L5V1lURWPK1TaTPfsCDMtw7Wr+t87JKiPACtBpr
q7yTq/zL1Y72ck4hLGcI4pGV+FUUWOejOxYAiSQ7vu1zeDms6OW/Gqy7k141q/Wj
phLvyUaVJuTC62Rt2o7192WhhcoJ5ZU4bl647YgsbOk0ipfPZFq6PpzaygH1Nx5O
M7rzL6LefGoq8jaB6Etnsd2dfEK/ISu4V1NLKk4e42EcnMvhv5lTLtAwPhZ5h9fm
8QVAKVw+yreirwS5KcjkuM4Zqthx8jNUOc09xioi92neYq9REAf22tzYVfdnEOoo
JDAgY0L3nU6Z9QdhBD0lNJ6CPadqjpeAmxoec7b/g1WiwoZ5Ahh+LwBmGtvcXBW+
GX7YK6MYLUSKk0uRLsMl3AJMYfRQxiNNoIVdSs4dML0Fpbn//4B689aZ8/mrKobL
fEo+/z/kA1CnCjBxKYdTV3m0b/WO2e5HpSWeX3bfg6bg+fnSPvowNajakRYST++O
ACxw5BjhCJRPvcgCCIwir6TkbDDO1fbKhp6Kb77VfBtddm19qKTgLbQ1RRhGhdGm
/6dfk3g6NTK5wPwku5eQNyPQKr6uXzEYQtcp03T+Jz7M1o+hVudhEh3k9DIYNkfE
IR9puY6I6rrapa8T7KZH2NZ+WgqbKB4f1qg6OrVQ43rY6WijKO38dtIcw4KAwjLH
PDq/BPG2wgaIXsWycuYNQB/0GzZi/nGlglb/zET4uTNmH0gZNRY7jZB7BooOxw9A
KzLdSYsDK4BE/NMsf+31l8pWHCaVmvvkWQ40IeOb9/zq6rAGWRwqLbbKjK1ezudT
uu4MTPqm0Z6QsVdFEYN9qUiw+P4aQ+lNbTcKcIr7eQ+8SqlM9BRcADfGmuHiJmDI
ZK8+122k6zSIqDLhv1xe7/HxvEhzwva58W9hV9LecIySlCkDsU0EEE0NJqMq+pVa
bYmr51PufEA+h91TX9Cb8d7JHgjw7G3EiOsszniEYcH6g4l2I20D5e6dt3Bxeqtp
MhhGK7FdPbaJ/ki8nyrOqp04mkAAix4g//Fg+dfkB7DRckYJyYiRuNIaUKv6eOdH
xis0Ka38UjSTvYFCYl+Md/HHlGkxsiBNYg9CoHNr0G01iMB8ioEtSeIa9cpT37cg
dI24lPNFosOD/B23lUHp7SHJ4vgTrV9JycunUBc2gFHoJhb23kvkZNV1hBpGLuZl
4HVlmeEOQbO0uVxALKWIPu1E4h79oaNQoLnEPUvsPWaGYORYdtOjRRBsh3iuUU7h
8O9qN3BIUwK6eLAZqqnaeE9dDruEJucnmWDAUSMd4e9X4sdiGC1eP9/9oxhdk2ut
qDtJlw3H3/6113w1F8Yw01JbqwN3uy0iC/QY3BmQc704o6NaYIHlnp5nZ4RQ6TWa
PqZGppP8NbSq52cogKsqNxKqt53uWoOxujZz8e0mQq169boPIoGPQ3x5pXNPKKqY
n4ECwkzJ+5GXNgM2I3kWUgpk3nOhZ5l6cPNYKKRU25U+47XObJlUTN+Cy2c0keuw
fbkrzD/GrN7Zpu+0Qc5D1vAga0xFdF21B5HHoZa4vQhRBJ64QNCRhRDASzNHbb+e
eyZtsRRR1IBQZkIhPYRddDRSa+qBEHvA+TyhYspkMY6HRtiLGcIy2IUW9fIQq9wG
vH6YZyrdQk28xFTicnyySbrvkhNjOBK7KHwdK6u62ZZiwsEwlWi20ye5cnwDHWBJ
OhunMdtaQw+xGU+fidyNQZhpJm1C7hFRxY/zuJobkQeOwXWt9noRxyxpmiApKct1
a46mgTeSOMDTh7RyGbSQHgwI2CpuMDxD5Dys4OssZctNl10hpLrC984FNevLqDdV
Iu0spL0fDaihlNGKbrmyKephu3yI4VnrCY+mauzDokJEN1QctQTHi3aaf9jj7ocn
2Fxmk62FD5TV5acQgQXbEDWW9rlgCSJHdfBUUD8xLEhKy71rztIs39d+DPl5Lae9
KBS3/QkGsd0JloaJidz8WQKB2C+0pktfjznkhlj8I8rhx/EnGT1j4l1b9nQpqGSf
VkuLOvWUTqXg618wu8ddwVqGrQZIqADnEpwMkE/DpoqIXz4+9ES3BJJGX+TBmuRa
vDIolkkkmxq760Jb3xW2TGAI6PWgtRxHjojhFmM3NfLXs2+iLY5rp/4wKLneQepJ
FMcTWw89zLoTIhqUuDZyRosrQerMgw27to1ruX8axfYP+xWr7t15a0kID0KjP5/i
lWARQmnkttcnM7rXeM12y6DTMR0geJHPi5VZY1l4ehI8BF6PVUiALIecDMD6nQ2K
0SeJFQ0X/sj7PZBfZ9CJkoxR/OhO8QIaBuhfep7QdYS8ygoyGhw5yaIzS4JpGfpb
faf1mWWaAfeuGHdZduCAQtT6oK9818M7EZRBh/3a8s+U/H57SiHVjjxYpXP2XU9+
HitjJKMZftgyocwRvIlO/GdkzZ+UHTnd7elsddMYdg63Dm7zsaccjxUduRIZ7ovq
uAl6WLqtJlkKuQqZ6d4bnI1twqqK0Ff+y/XZAbP5QIkQS8SxJGzeKDDMWrn3iBRT
fliaWKDHwx0gGPKN10r06piMy+d6yHlHh4385gUGkHenrYZLqr+70mCNHf2ul/66
yM2oUaODqlv67OX1Bf/rJudcEwxkISMWjRZ7ZVqRxLnfSSl2PH6ZBU8qyZoWoo0w
tLo8pl7tB5EXlWzHzpEaPf703GZ3IW8yKxpKJKa/WRQZ1NeLxerDxr5fSIuOEfjs
VB6gTcTXL5cIM1vNXYfgPHyfPVla8K0GO6GJJIhtrnazMocK/weNVxTlBL2DpaUG
LES/JGrIorpAYEBmAAOkiJ4elzO02tvkrta2wQ2f1X+oWpJIQCqKhLOpQ0JDD9kU
CScpqXCxQdyYfJeEF9F0wsex8XImXjB7v7K50HKyatObptbpne1X0aDtY5jgo37X
PH1RPlttPj23HHs+/mlI/1L2dxcG7fyluCQNyK3YsWIzSzjshl8BPtkLzBFO8/L9
tdmsoA/RNXvVAyPlQcgZ/jMq8dOJkY/vb3kp6xh5yK9ytw/JBXQbSl/ccEpoRWT8
/9y6JjjZp6nchGAYh1irr0btby3oj8Gf+MkdT6Grcv3FzQxBxiz2IzIWA/EmU0nd
mHnnBuOAx/sTn7ALwh+J8JWMHcxG1iMEiCpFWbo8qeJVe/A4Atj4T9ZiRsRUVtcN
N7GuljAD7qTclP8pPwzaj+n5njOfWYy8hfhTPmaCGKkyKdJ8UhSoO7CJ2fBSWp89
h/GTVCL5gdK9KxExkmHLX2CtlCERR29OKBSuvYTZHlxspt7S00qRKCpM3yJdkmRe
zvW3LLm6tq4Dvjzsxfr2JThxyNWMPTbmaa600+ZXRdkGSCu0Izlw4A5ctoAOhTsU
47HysTRE5H6UIZps+zGsDhRnJmjADzW4Zo1zOltQS4E3GxtNdiSjlSfhYylqi4nz
6QnbEfJKGhJ9R2hpPreZW0JynPZ2WRcsY2gKv6V2qa8sD2bzylA03Nl1OIDi65GC
U7itZNCt2cCkxVi1M8j/Xgvb820l5ul1vwraNwfrsqmPoOubSEnZ4oBow0sl7hFA
WkaWNnQUJQFcv3os1OHFJY/7XHJhizSeAGHtpbncXjhTqNh6yZ+s6c1YDDF2HlVn
M5tvGzrTVLAyd00FZ+FzBRFmdrUZKwc9m7oHeQJXQrcsX/x+ZCUpf4SBqDIRG5GD
rakgGqXO5b9GWpYBxSwnDL7A+PbVqWYAqzu4lrrKwHJiVwZgte/bpwVMHGDiR0R8
mCjC7b0JmHvznBm6qKIX3VoPn2ruM9OZeuIHfg4oND1PZLdIsJrGxcr+gymYgsCB
K1Ay1qKhOW9oGYqLAFtFvlcfNGXJWarX5/KIeSePRY6ljKSfbKRYY4h8OOp4Hc5u
OWC8zgvNa90Pk59lkMnFrGsHmAPCTQgYVe4WliDQ7Pb7HEpNxYR/0ANtr7a/NaWt
UG3bpu1UM68Xhe/fqPDfDN7UWfUjEx8qlOtuFhLGj16hr18VrvfZjWVXKYLrYOZb
ahB6jZml7hOPrdEAkDczuhaWRVacVIKNyCRMlGUv2Bz4Hk1uI0ZHDE4e7AvnY3kN
uSo/LGij/1v0su+W1woCUUjXcOJq7ouKqcG+a1XlLOP8fJv6+EydSZsRfCSjyAMr
ucc+XHVSm7itq6Q9Xw/4TCRP7NRGGdWQdbVmNy8TfgAyp4NE6nrDyN2ovRD6lxD0
uUnv96mER9DjD0QQ+Df27RfdpETuPuC6DhtMdgnmJvRdcDXyx6+JQ/aONMoRrngz
2kU2q2NIYAFyslv7435G+rE4y1Phd+I6W+/ucCF4tS9lywSiMf2B5DWbRy2JRALv
9nTInNHG1XaHgRfid2/bJFzQTOitoFtaC0D8l1o+Y9B/OHIk9xVN1DWOF6hQvg5i
iZo9joFsqER3I6PI+VT4oaRbdDRzsFF3WxLhF7rbe45tr93y2HnuksE1WNMU21Y9
lZacADdXrvpS2ofF/5X70khhlIvFejR4R+0dIAo1V/PhpmN5QJPesVq/1MlI4mg0
DKP8Ld4FAAPQAAfAACwalOcAJxFPMVMHCol8BCj4b3coQDS6W+iDhSyBb3JGhRTy
N+1GS1XMFcgO/bbI9mLm/6c6zDcUgr9j5K/jM9tFV0Ybp8XLOxpUtUsR48jvCiwK
/oMy/nkjGlrGp1QlcoCo7iDwoajmv3JVwKL3eWZioV18VA/djYt4pq9ElXE8nxVa
N+f17RNAIMKlSn33jDOGSKAYi3ik9ulzHYIkuwvSFi0i1wExImI35yYR+LQANqNC
dRZah8/4MkuJOPR2irShzNqjYbO2v1C/tZWtCRZe7qpNIuFdTCMlRnVi9Z0S3Wbz
h9XcGOK/ufk7+b04enLI5MIUeJJrWc5W9h9hHQLA/lRFsHAnTzjW4P3AJz8oyuU/
4suBQG6xytQ8kHtlDgTKqh9Lg5JhAzlPdp8DJkcMbde+QNYuZLIZ7B6nTe/ZvYeb
pGg2ZDYHdFTNnwDTJ2BhLqWsPKT0SZKGEfMK9q1yE3nJuT4CF/2v/7dOXKg5a21d
ffuObHZYwY8OB8jd815qMYNxFZzrnMcqNu07xPdAzIFctYGd5fgVlIpcmhCbKnNv
wkFe7PzpVW95l/MlapGneJ4B914D6tbwG1s7cHAdfzZZ+sZGRVU/D2a22a4QtezB
W0fQIluVIMEYwKcHvi0fuOE9jFpOV9y+vdcJvR+cgLNoMxETLUr3KysAijPAXWmV
NFT6kTUdrSQOxzJAuycYNw+v1e4T/d9ll5tGcp2XONvrPHXe8X6/6tj1+S99N3Ik
zDhiVIJCmfBtI6Hr8cbeBvjAPJ5Ys5HxBxHEYGOgvz+WWqlnBSl0sG8bGfxbYArI
RGsAtBUIcgy40s4EkfnmraXbE8vU6CX67+xgU9WFiacRqYE8Nla20yD0Suhqp9oj
hl2qjjSXk6ki9ht6huns4jfr/BjNaFXgsli6a2X9PPkZQRX4qorB6uZcrc4gzz63
LIBf8tSnocZQDyQ7Ek5IiUZWsT6DxUc+Zl5HqZAHp6o9Q4ltiq0ssOHpjWhFvGhT
z1+cqO+cBJ3NS5O9O48u8IKK4igh3HsU7qMy1u8eD6p1YcTroduxUsBOGCDIEBb+
XKjVtXzaBQUMRm+Yk7VEtmTp0B4Bf7YBtOlEIpveyM2OB9WmTz1qOHlr/sMM+U72
CTygnlvnpZr/CkJkIwMoVX7QjHeA7fT9zgcQBOnHi6f/GAJ0La3aVwRuvvoIDBLi
ECbz3h/QrUDwTcFms/o64bAnp6KKII604KxP67eBqZ8Z7ENdGNEK3q8duZlTfHab
xZGz6N316d08T3Fz4Qxr5zrwvOqJn91c+IyBOru/SLUiRzeBWl7DXzohLtm0JKfU
rijDbh7ZxT5CvFc5XMPBhwWzt7d1Y6dhnVNYz3gdobKa+1oRngtkdWZiY1TtZgHO
ntJzCc24kY/Zi+AJGRHsuH2ASPCmT/IsmNmniH1T1/zCEVE7kcpDkyAIt04JEfn+
IM3DvGOvwr2KBEzTWopviRTZdOmcnhS9MdwSlOIOL5JGAyhlUClXugB/mIOHJKOv
b+ok6dLnoIP320e2CMmybyFAxYcDhPdeM2TOVvbGxg3bJEFHWfyfX3zomds3F5vC
ujzxCEbUMtoZcj5r8/1V1Xp7wIMsFi9uFjS08S6+zX0/wvoZxi7RWHKVJuEnxhe+
oPM4mekey3jkSyxU4oBg5jUrHo4MTKu1diwkqvpqFtOxhx7G2gFrvJbi+uJVk0lp
wb9i493hJIyf5QONrUlqdA1NvscFJyEp3qlctA+AHSts+CSaRxnJimTbdpdIehk/
cFWgn8vcv8zPaqRzZ3r3S0Kb/HlpU/RtLOgTF37wIVbn0koN0FPGpJTWIjxio8tG
hdk7RNQAOeye6o1p4ex8IC2aZOrh+jXmfO9g2GCh5FK2/ype+PUtaQcYKPucK6DW
qzMIy5kb/dXLpeK7ZkeWxDzsKoYshssVI+aIB/EyQPIIgLZhUuHU0lRDYphjOaH1
x0g515WOZq2dWUizhyhwhZ38kM6Fmwtj0cBeAxJiaIPhAbBGNu1RMsWKmOSi2uVM
4cXFPkneoSkwh64pQ9RzSKsodCabJN3TQtEKtpOaIuSMHGgeskU1Shr4ZL0a+GK1
qtGqJZUARigoIo7iw5hKjzSEU3sOV9zbBNjC0jS+LY4zAzjWYkaIuWmj66U9VB8Z
xJw+8ebggur0LzBaeAsz5AVpcWVanXGDWnpjgzJNPhVZCp3mVNAoF/NSYvhXq+qT
aS8V5Q87WqNm46MkolTYqi9xi3FTKVEpD3EfCjKfzzqbW1UN5qg/fBf6K6kez72U
2M1O+yISTjE02ahmPqd075Wif7zwRFjSIuCLV7PValGSOqRbbnO6j618pOVhOZbw
piJfFSTzlhbtNc1QuSOUa00CAIqjDr9NgBMSLYSw7WDlrw11c4h1BmnPUT9USXom
KomS96UYu/nApjRADok7/qmp+jKzvx7dpWz3vToAmn9GS5to4ngHgWukr7Syonuw
Ch/VL2i78zqaMIZ8uozb8NzsSNrWNgloHV233DGsOWA7aUBHZAHT3ti88jx+b2zo
+h+i9NXrn2+R1KR3TLRq2t2Vao0BhnNPJObdEyVDAwf1JQLSMGOTEIpVaaBaKKCn
1uDtZpoqz/qT63MdZj23f3xZRZ2+sQk+re+I6I6nxj9e1+hv5A7CJD7EKuP7t/Hh
TibVJ43goVATqu6G41skuLfqHL6QU3D0hcCuYh7zhLX/4vitbcCJn3vGGfvXHBWp
sbB6iRym9WAClngQL5vRU7kH06xr3Y4/ICoVqN27l7Nq+Ti0brEcHa449lQB1hYI
B+lnnuEZXbTMCGL2XDa9wWwuN318MCf3UBKl5jAdBJUXmRCO7aoW70fy3+cUCM/Z
+M4R21Zz2WAH6ClEe7lBaE0s33mzBAoPNyjbCNmXNx6iGI/tSpomCczWbf4iTD0H
wDCMaQ12HnbtN8juVxbGV7qqivCEaCGlN3Ip+8feS9EZ0xvhJZim5nCFiTcVWstv
AzaqPhdrXSXBLxBeig9pVk2I1XECjE6H6T2J4K0urfo8mLUWvCr9ecJnmGfUfLHQ
D8DanRca9MNqUKIcStsN+lExVAyO8iU/RRI81ryf1F1fmthgFY5q4M+Yk5YbtvfH
/mwogRPlJO/OZ6j6ErvL2DKOqqoZJRz98n1avLgL2f7P2y+QI3dQzh9Wfaz5mnER
j+Z3JbWavXyyd9ugYKiOeN74BfbQCYj6/qCsjmT/8yJS+wF4bNC7CH4I8GEXNwgE
XsjVHmKu60Ax+S112snPOFGZ8rdhQ2bnpii3Di6eyi88Hb+WsPWaXETzjjnJxgtK
/+Oud/LtGuL357nvqyBHvTw9fpJzkmFRKBCHJrxA5T7TsbttfsPkdSXEagSQrrWq
IMszUvy0KSGxS7FHyXX8TBKPk+E1w035f9gR6COxAxnDUo9poUSnSxJviJKJHzGW
VXbMCG0aL8c/pu6YPmRf1/EGsH3QJZ5ciwQYheyk8BlRdpg/feSA8wa606GY1JAT
pOEOZr2J1ue4yJZquEzIG5NwqXE8gO7Aikl1Jn0nxsYbEJbUO8L0n97l2kNZTizN
8gZ6xRncJbMWTWD+xCOt3eUoPHKF/QXBCHL+NLEeNwTvfihJVUJSXL1ol4eCA7kI
FsF+gIKyGCHXI9x5kEtKntyz+Z22BS73GhmAKFLPLwN18U4UU5P+wKD3mjq44cjw
fg5wMO8sIkZx/K1REgClUBaelLBfkuPIxn15QBh/CFJJYq3frnOe6/2WkWYyuSY8
QfqrEdOaE+yuYD/q9ezutTossdoOlMGOAsvRip4zIUSl6KE94rAjyGXJvV2DiNf2
0RpDELadEiacqt685sNSJgRDyL/ARcZt2FfAqE3y1DgSqYBGc+6hs9MRWB19Nx2Z
Jtsn811a5m0wqQARdA2hG8M7CdkVP6Bfb1jhHTzqPzicUUrn24D/GN2IYpO4zKHp
aZhSGi68wqEzu5raN2lSwjsd7As1JFOfbCkYp/lbUQmHolsaG8pd5pzFwKcNJxsR
WY0DQLrwllqfuO7NPMTbDJZR9KEeRa0LBqTGn8gAxK35V65AaFxcRbWTUE2GOhBO
o20fM6W5WAtDn2GqsRoizOl0lieKrSmop2EIT4x4hXsgnmyo9ss+u9829B++szre
s7Ixz18bwL4xhjXyVlNpVUpMpoibATcfxP8c5yEpwfyuAkrlfG1DIZWgkfmIzA0n
EiFRTCNtgTEjB61qkd5Z8KT6YQl1SlO7NdGT1dgOpsLHxmqXlL3sFAwLvFiGEr7B
+/djFn8fxq33QjBUKMwWzYzXgiAcOeUyrfEuATWqstnLBvmC0jeev9Rkd7pOVhpT
GfATjzVnaj8V9MLCG/gR6GQSoXV1LMfIfWmcFcM+d8XpJ4lLkm0gX2veLVim9x82
w4BiNLxmHZ6Wz5tH1bT9NihmHzM4kRPWkavuf9oNEwg7ytUXUdd2mJL9zmW03qwR
amvoMsJLXPouognvWd+FNtYJDAx9eBvWoLu3ssZp75sGfHGj2Ogwy/msBe1tO4ug
Sn3Zewiv2UFqDroa++b3DGnM0por4uYCefR8dIbSOMlGrkAY91tAKOnIKNuBVkLJ
vVcDQ0t8bYY8SJa5woZlEFXSzcmbKDH6rZWqzJjTj3prwj1bWtuQqFHd5RkX0Gyn
5YQaRTNH0uLh+FQ23MZkffojRigDYqLR94ZGfmJqTTfEpnpSq4WkhtTgx0K/CmdP
92zX7aunt55rtXtxE787j336uuA5+vDxV6dHCr3k5A/ADCEpvxAojzMEyDjUMVJI
XRTT6dRdtGehDD5enAloIY7PGx9DmvNlc/jzEZhA9XiiNuNV4FIzsN4ntLD9z1H3
Wv+8wi+mtwXpTRpMRHnJ9HPN4ubz7ggPwsfa7kAd5Z59mXRPHdgBC4d1LhmQ42Yb
qhGP7zAJyCOTsHXfh3GsfcplW7SDDXuAKsm7q5kxp3DCgfsmI7+izQi1WZvGO+y/
+Qeb1hhMZvBpx8Y5GFfh2W3eLNDysSXrBU3sRPgNiL3OrnzqNcXZ9q/SQ2StSTuX
kHQHYrXV4w7yxpsN0kfoYJVFnfWHaL5ufIQ6rNvFPM+4IzWWDiKW3MiG3EYi8F/q
Isc3H+Ktxoyv/mhPTUHgN3wua4oT5rUOTDUG4YAGQxGi9Npcd5Sq/FQWo0TKyBS7
UABMqsF3v6wMCBdX3iIxlp9HIvlTl/TQUFS0JRcLpA4HQpxpy9oFbVFZ2dAde2Eq
SVKS4mFKYvTJ8T5FWfTHahAmkrExIY41ZXsFYFkar8VVfgGcaCzqxnpM3xc4WO4Q
Un1yU/01uKNINjjvybAI+RQU3SQtLupOZPEQsCvdwCeQJWdqzw9nwkIi5kKvAVlz
hnDnITIoGsJnRdkbMdGqwb1amUVCxjYI2JgfW9Nru1d3qrK2+Vx9jAZhEmUxFpgY
dGPMfEQVVxTVEHNu1Nuofhy8Y26YberSHqi1F4/D0zMrmab7oQY5LZl6OJdhje+a
rA1cT4PzevY2jS+t1tCuLSdCLYrpLdFmlHE+vF6pc/IJfvJx0YDfkDWcLt+SXP16
tGLOXs48kpU+UMxSbd3anzGacVGSS1QLmPGgzG1rbkTelJOB0eLQRQRo7766Szbv
DUSRtluUUtVPuTntJ7Sy1fk8lfwzQK5J6aXlwbisyPbBUGfKKA3z+GEBQM76toyE
SzMAUHGCFeOU/TibNznn4X2Wjae9dqCrBBfVn6bO+yneBzNTK4npKhdlVHwLflxQ
XAERufY0S7gD4IfMQANsmOgq1rOxUFxp4eqX768u/K33zH6Cow67q+6hHu4sBaLR
TaGg9+iY2yJDwTQGRtrkyaIMnu8gWh0mckJz7JFz/HkBW8y6QY6xl1E7Vk1iSRvu
Ddd20coA9XcknDF+YX69k1gYuDCersxaolOAG8rtcbTTfXwUzRr5C1VGfLVljTXz
0goXciffqh+uSnpl3kvOSnI5O/oNn3YYTAvsmlWBiCaE0KaZZbky0pgAL5WD2NiG
XugJBdoDIbfyViAXxuNf6AGqHtcBiMyGrJ4MdYwY/0713k/OUJmPhq4gf4EV+z+V
bcrHsotJoSAhL9/sC+S/8MCAd72KPeAnQb23txjOIPeMeAcW3OHU+UF84CofL66Y
xEZo4OfFiK3+jKDSzAP7G+FRdSIA3lnDKeSwxVj0RQgeQ+3RCBQv83kgQlOtig8S
0vCWSOowsxrBwQFkk72ESPSjep4zyOCLjUaR+HHwqlf1LrGL0Po3sFdtnU7OU4r4
2vSS6NIM5WLPsTFAAY/eSfJcNJU5yHEJtdgCu9wDgjnXsyUciiphSfnccu+MIXm5
HPLErSKwJmdFO1iZOL6uZ862g+siMMxIUr3rYd11CS5zH+ND0zyvXkd7efg0IEos
u2SfywsYL2iPGjAi/HBQB4kZFMRO30+cbjwQD7RgjsLD+vD+DPaQKNI7qlhP9v8I
Hv9XtN8pj6tUrFpD7DHnnPFSD3rUy2odWkn3BCpvPNN2bYotFmjWd33QwKHcirTZ
3z11pkocVjZNUhDakHo/csJIPBmoCDvKhIpkJjqU59nA91G/xodr0NGnfj4fXH4I
bDZBq7066YOztpp1j2AkPDpx3Ahz99aLK6y9s9Qu9tCo/qVCYpI3b+odGTrKn6DX
CFkrjwqFCKpGFUB8cRvxa1yIzv0AjNTWS3nwY9sbMEsb/SC8BrLBnHEiRTvd+ezw
BAuCWfE6diXhKMkZyDmZvaBulxH7+rJjhXFx/trAJCO/sNljWNih7U9vecRyc+tk
6RiTVbD7VoHpLJXttdNwVPbj3sKoO2nEEUXzVWHN8mOaPHU8qY8t5O10xRBiNO0q
w8nWpRTw90yOSxB12AKA3i7uHd8vAgVugtMWQK+U8zrBRjIqxq8L2hISnDxYNf6s
6m6wJS01ibF8Pc83HPCxv6qlrOkYjHyx6v+/0Hz4BTnpxDa8BOgM58LxiDxJWm64
UDWj9eN3nqr+vbvQnbPkm2Dgx/mAzpLP6nBmyvlbRA9OSSBQxNUlx6xJX3Md8LKI
Hs+1+O7qXzdWP7JXtG0xOVHM6X2iMavNmOZZBy+xsyYHh3LoEWKBlPkGgz5xqDQX
iDO6x0KGaWG4F/0YGe91QYW+JBnPm5HRL9LNxTR0P68HzCsGhNVp0NEOF8P6Tlro
qvl4LVZm16x5tQmF7Cr8+fOrKK8+LqtRs3eq/Hi3DRbE5lXqgtiIF+AWBcQ9DcXP
Ss6N1Is1MVCqUpzpwXY5yp7uNjiJ7WiZvM4Di+pyUVHE1wUcJMIPS0Ys7UynzM27
ILlw2bTSxsnoUwIL/fR8+Gdulcye2ZFx+aDzrOl8Nl35pflVwlsNcnUM3gwPxd2C
I0SYZlNX+//kKSMCJFJZM4vTlGpCDqirEQC7Iaht6QTfw72VQPftyun/+qvOHfbb
7plUCKmIuT3wm2KBcuFLhAJjwLDpXf8fsL84817uhJzKyy0uFb6C1VRfD/rV4L3H
kiBCAQ6zF6oddCB9hbSiYs17VIKua3XVmeqxRVqrBr9V2cfeym3ce2zdoRujDeAB
uQGP+q/UY1pNwSktF0ZsF4S1tSm59Z4pJwqD+l1Mq/8Z/B+i3yUWxtfgr3GrfYdb
LqoMaIN7VcNMrG8Z3ldIeiQwhZM5hD+NxvTufXKGjaAFAkqwlrBubpBURad9/q09
TP/cUbjvMkJCtAm5wGdRgqQQjdIFuGHsMRG/qYi3NfF79dkerUZkoRC9ymJl1qtu
SknvF+O0mzTh3p/U8CBXmqEahYIuauKFmTlBkAD8hPGIDkeIxkxpXBP5JPOclVtv
3qA0eDViFxxRvM8sPD+kflJIFhO4dGxSsnw6bpnuUhCj73I+QN8eziIVB11w49ge
9fIotanXDxOhUEHePWyUKQmdSv7BJKd/eikpLknRPoD84TU267sF9BPHtwaOWjZT
Fep1653cP/ahBbeLO5RXv+AIouMooDPosgd29Pd1l0eRA1JPL/GKkOygmgKRGqWa
YjYVWN1zgsw0XRoUbEOh5vEsjXLddXl7CxEE3bwLrVCMKiNSH9h9dOKjoU3h2TxE
R5SCB46Tn0zmFPzSsCH1sZYMpSB3Kzf+LSf0fhX7znmJPFwVihbVSKBxMjlJztvH
uuPv5XWJ3NwyA1lbFHkOgWaLp0Fc6lfgBQSW18OvbOIdaoxgpp72AP6shXFieffH
O+3UR/JeZsnsz7jJ1llEFluoW69UWrWmtdYmUNq0qUD9pjInEPojE851GZmL7DM9
jcPLyi3vQikd4siyT64lJIypr9zgHlw2L/6AU9+lOAgAUjzLozAE5muTfgI8yLXT
Di+VtumMsLUDNCf2v+8CoFW2gFljv4TJPzHAo9sjtPzPtEw6zsXPXOYrG6caUsv+
jZzlvusGFlTYb1u8LKs8MLWh82Ujvv1cptz4EjFj4G9gNlNCGUKZA802sM9tF5VK
H83cL8AuYGv8yFOYnNzBCJrzqay308TS0KDZJ4bZY6JbuoMHu75VEawlqMv8ZxIo
/hAVCMZC6jpo7Ee0mMWqarvEM0xwEpoEB/0zxymKBQkF+QY6KGrYDTuY+v5jNej+
vjhewJH0IX7hGcrUIHA8TRolteKnT5ll1NEhBUNAs5uomEad+DqaesQ/h0J+erK8
TdJs3nq0ugSGngGHuYPIC/BhkdYB8VnJYsreMhj/Af6YOt51Fc5ABYPxSaN3U7KT
FblomSfZclrh2BnAO4FDs4kppWnoj9wvfaOfcHq+ILDZ4yDQMS/PmT37WDJ+Fuly
56hD0NngR51Jl7+pIeCxBb2BWXCEKaADFK1feQr4lP7qUCnBZNsZl8OVLCdl22Ev
GtIenOgG+QluliKCy/FvMga9jraP77QgPMf10YcydonkT/x3a7IIaS8onEx0CUPU
FwyHKFdnUyo3BNu8DcbHIbDEncU33ynJRu5xhJakBAW8QKXXSNykM8iTfZNcy7xt
JykMxONDCdJmpsUXpPHGnP4tlHhlIh6qXtkCC1SII+1kfEBmfGrijyMUWuAQLsG9
ugiAwhfB5gQnQ0XaLaSCoR1rUmdgkbXRjNiGBF8FPKfQLXrhvOUre5/qiK+XLV8z
txLgnMXHxHybSfhf51cjubDUzMe7/2G1zJ27rkMIJgUktaeaIgAGjGjHB3OIwd+q
UOYP9K6lLvAQaFccplRJtzzq4gJAa3hyeDXLjmAxwcd2pjH1yV+bev/EZ8tA72T6
Z4vOeNiQAcTCShJ9FFibJqQJsRw3+9LtBiYBWjFD8g1fwNXDRp6vj4/yjx96MCFI
Kq5AxznMx/2c6CvGEvAztuKnrJZH0jkKKzhLSVr7RTQMwYcc7ee7qn9Nuwk/1Oif
NsJxFJN7I8UuMVCppD78Xl35Wm5NPC2BzrvoTXheQbnSdyKleyLLr6ls5mCHjS7p
XGdOCXyGgBoNysmMsDZx1v729l3k7b9G/Ie3ZV1MKF8OByqC+nWwjtE4tCMUMxbY
U91xpid9D+s9MWcLce0EFc10vWKBRycef6SQVVXEKlo/dckMr5LtpQz4l2x775o7
Guef87jiIbub88habi6wQ5SuWPOZYqGubA/RFRYkT2CVdqjMOAV/WzuogqtWfZr6
LzSquMemd/seXldkIuB/reoqC3+xTa10ZoiiLNp8/3KqCyYBPAe+352xCxVUP+Zj
ZXP58mlKKWdTb1lBn1Xry5o5E/m95emxqSx6E5Q3gL0S0UvXTpeQxrqJ0gdk13nr
2ZtkeHnvJLhRsdyXoIGBskSFph82BZ1+tO4EjZ94Enf1npzNL3A56vFmtKn6mch2
+WTA/xbRj1buiFZaZxK15MSidDfGqca+UXk922+zu/VvCS20ARtGZu9SE+rtw22D
Aul3XleNgyjXxM9kF8Z6ZJlo/yic6paQcOvR8+1rxJDO0Rxr9X5KTDCEJXcKco5g
bLjQvwEGth3n9yPc5TvurGAhb5YxhCPjAXVTLHb4MCh3gEZpwBOJF3lEi3oHXd0U
LtaP680yVGXDjz8gV5cBVF4wLV2lRusGn33c/gbfrBoHenM0XDEJ8qRmrkiMC21S
Xpw4IAQ9Z1bLZB3hL41TpianOSWRF3ZLyzZUGt5WIGX3ptukVd0j1XylQRZf5WME
z9Kulb23o6h9bJVhjfd60+13iv4X6iO+U+TSeLi1C2j+6zdz5dlkYSIWU6aJWII0
tpukxa/Zfq2UMBijnP2IcNyF3tihIZ1nfcBltK+JcEKPef2ecyzsuClge4S9zQBC
R8cx8Q/Ac/ZoqKi774vYOeuXHF4S6fIZ52ER0i9ffK5mZkf+LW1L0a6Ppw5ip2nO
OFwTl9VFaLcyZaRE9aUAGHNgTEl+rsdTc0wSmggAa9MAlh/cRq6F4I5RitLNfTx6
G3O7lQCWUYqqhSeYpZbWovEprolB5ArBttyj+8sI5+luVlYwljCKRc7X/Po3J6iY
h9nPZhrf3779HGT2LF1AckdGIE5HqXZhs1ffAtyC1lPP3Yet+1eymgHp9bqbRYHo
aHqJORAQD/8EJDXkw1aDlT30TmJiGsAG2OwZrwhrH9uAZ/v+e7HdBBu5QcP03Ijm
fpiyzO5znpoh7k4BXW9uxdEFcxw3So2/W3WboSR5Md0f8acY2khP1A7qXk7bgxrl
wEorF+r6rx46hjrHp3rzP1ozd1vF0vC0alu0dO0V7t9twzaWiR89DavQt8xqPkXK
yM68pZYFUHja0a2j81MGMk/DVeG5FF3vw3gw1Zh7N8SJkaaG4jO7IruWbnX6YKdj
3Bi7kPH9sVk7IB97XLqGiSrn90tenNbA88GNdvR2GzcxGMtM4NaCy0sTYcnjOFt2
VFG2bZv4S9ICZUnUpu6uahwv+IENYCiEYkRhPXx77eFzKWpgDuZx3UUiRjMPy+qn
njBDzZilaCJq0MQo2rXq5SQAKLoQhzedD0pY9PEvZDtPBdAUjsjNcc34leWtctG3
XEYJVorA3cFOCEFFDtyjhfEh2G19sm/PYmhc/ejUNRF6qkp8UJRGNah+EjWTPZIc
dJwtpeQEccasdy+mYszRii/ckDxIJmb8q4WWDv6zuAbdVDybS3tG5w5gZGFkgVtZ
/bBG77SOh92JjLmtSjHjYLjwDX08Vpw5JROtAZxr96UPLjYyO4fDUQ8unjJX2F58
M9jJJPN2820bVq2b4JTrMSMLn6jemy1VUAs5KyHQxG/d3IfIMQnghpx1lN4zjmLc
yo7+0vlWRgTRPYX+QeN4D4aNA3RIqwJzFqNRd+b3YFFJjPIc5YbIWUhz07ZZ46D9
7PbA1Q5Sm4l2nmjByCLULi57XQSDfpKdoXjmoLG7EIszA7c2OVx8p0n2vy1jBa/4
rPyZykvt3pd+UcV4qzh2cYnL6BNnAVmPoRLM2n0j7Ee9n8O7pJWb/FVs9/zh6qxT
XiOzSCjvJ4k5WrWhFJCStINq5Nck+tqN/Sac+OhpKj1zNmrgVNo44ayTy4+IwCNM
nC3qIdlEGVX/jIEma9cJxnMMe0tVOpkeqm+1TV7VmG5+rEPjVoC6jE8KwS9gsXXp
H8QpDDs5MetkM5UjTFQ8OSksO2MSIOrMfZ0cs4dO6/edpnVFoY9Et1WmO8gqBi+D
VxddqiwtAbetrrdPCnqLGPWeiClcQe4uSjCQhm7pFRZx79Ad2x6ZhQ8izpvoGO6Z
YkXT6BbrCC1+LKv0d6QuuagODFCR6QGwYv6A4BUZH/0rqueIk7AME0W8PFSjg2FM
TGCOIfpK7wy1dWQ4MmngNFte9hL8R0yPj5j7kyvSFWnFjtiaUHAbeUHZZ5R08xu+
1JNmOZWrpcZrPs3nKn1UiJ3Gn6id61sD/6eD5Wo80CuOlbBmyqPmeC1ntuGuW9AQ
CcXNEzPJyB1UNnWUU9kGKQoHZH7NTs/32oqJc8w+8KyEi8+dIWxsi23VTjB4CCW7
PuOu5AFNs8BJk+4jT/2lw7+/S4yfBbXo9W8IcPXPfmfRAJM/pM2AJ3udHaQllskz
DkgYS/wuJq3GAPlJyc7ICTejJ8mYeSN9SIN9dgS+QUqbd3iAi/U9VfEuu4HRs7fq
pHV+MOTVhCj3vD4Ga1jW5ObYueyhvEGE1Nw7UMISMaD1P4tFkp3otQzZdUPlQkcG
g9kMo4xRh5vaeWnDldDs9h/kcQQuz0FzC0xu30OVoaQ/TW9PFNadt1foDFXu6Vse
CxNNkfPRI0PIcgEyOu62aywHRXVGdHlFD+bE0dytZy2eg3nYvDaaIrmLL+/DcVBg
g7khUnb8c2qQQuFVCbmvp0LKqW8CjqCfhbZ8KXEkywiUjr43SpW3Ds6RH2VB7afL
HBllALPSnJ+eqwpWYWO9VRavt41x12rq2DSfaLztPlHlJwcTHthtmqYVdDRQPZaE
f8e5tsP0utBw/HpqPqtNE9HXcLioUbMG2ycOHa2w45F0jOWbNu2mAwIWnbt60NlS
PoaCe9yuGx9NcW7cZ+fHg+xSEYE83uzENTANuKdbReBhJw7TIWebwZJTCDQuwfUN
aH4nRv98W9jMUh6zj5cZSXG2wO87QflklNdQhpqr5zd9yk7awCKMcAMtKoqtt7ii
WMGC0HpU1qw3oZJ9h6Gh+8Bj6kncc0uUsV+l2zKzNYvkDypG3p7iO97a/rTaST7S
QP8CvsWHc3XoLI46vWXJEh3joXKr/h7Jw+B7H0+IsLNSTD0MLde4q/On6HPxVAQy
cig5W95QhetEwk8AXbBmrM9cHcC02XdysSSEwHjEOPrEiwEqrv+XyWhJzY5c0gnh
EMUvHCHaqEg0Ww7c3wn6q7lA6ISjY2FR4TpIEod5hzsGzq+XAzgVYGsBrlQ8MKkd
ctfzWNvIj3VmWlx3FhuTrrTCTtl8r+DSSa59UXDRebXt/DY4+P58z4nyS3CdX+EL
B45Sr4W3w1CeND9BJ+eZwlkeYQaNaYA62v7ryPdznKiEzO7QRFS6VZcNiX0HjI+C
XWM1qgkYMybVLMVfCDd4RhypTAWeoPEjr5pQKDfaD2t7t7swnInjVUKzzxv7QCcr
EGQwO3M/GREx8zxI0LbcGN3TIMy0gta8pa7nUqjcJZY8G9fTiLyK6MF1zh48kuQF
0ZNViyWmYPCn3hr0BaUDyfXYkULwo/2C+jMTWs7E81TK8Oaj1dpvLghzU5wIjSle
uiFABSDG7KcEJgSAJgonR/hy0KL8CJLFVlmsMJr/5vyt+1UBgHwVttIZg85cPObq
i9n19emf6wD8ORoG06Sr7dVZszwa6xMhMNRahbs1xpO0mfi2VwhP2xoefiWdpz6H
bTwdo5kVH+cTWianU9+zdauacP/FLt0KB2mYywQyL9l2lJXuJAlPhZGVc8BvM9Vk
6o51Qcjyyvu8THcnRenTKQTw80Flft/8U7dMyoxZsdkbgQyNqUtsEYXfE61NGLsg
3bHEbdtuGqeqWxyQOyVP2+qAwxhEuSuRMJTmdKIukA8XTl6myQRs8A5++YfZxBwz
rynqBQnTvPGddy13QFyX4E+9/s9Ut3T7/OoDgBYXOaUp6B6cRCDW6XfCxQz34j6I
k1m8ACfl7PwGRVSmIkJrdZY2ypCby7WgV9YclBBid94tWgNw3XDcz5HRp8Sx1Y2W
PW3/q1YqX31I3qfdRxcr+qEctSs5QxttcEc93jKtR1y7ZfKxw/qiumUcufueQpAJ
Bb6MZkuF6V9KHvxI5k3qaSEJc1WsTjh8miXVO7Bmghvr+i0q9mFANq98J9ogDndi
dJMzuGkKMJFLVRKRYspDeV6Vzl02dRVIAQpbEs/AL/PwGnRpowQ2z1py//ze/VvQ
oSYTYkntHrYkWFmJ+ERLOGgOPt63W4m6mSFtHG4BCl/fidqBy+t8O1IkEIIlFYUe
7rmEc2gVO0GCbRiOxTtWre4FtOsA0mjNJdffCz4AL23IXCaougpuF7aeb4R49d6x
HSkJ5MCj/xChTZMEV347ob3UQ2EvZYUuFq8reV82zQF4L5h8VCm6VMvSNOhP8h9E
gHLD83MngGk9TKsQuJZLClg3FfPNA/udZblyADwIyXH0u6d0VoUQ6CqSvJPDYhVH
IZ/D/rtlVwSIPBTb1EkQWo9+1MP5js3hk3u+Tra4Lzq8NtVXvA5mL3nHi90Ds+Ie
wY2dKilhAk6Z+eeqW9yQabvk9ES16Wp0ZYvnBIfhd12H9QzGAvx74gDJFKSSJsFG
qmDNdPSUxtyQWz+dTjPvZHGPxIEiZfryWzqEPpfh1m9Qk9mQRGrXZ5R051DhLk2L
jfwLAvF17KNDs1VRO9Rx+HFtlBS03r/bypBt/M1fTReoJm9oRye5iKUdOAcoUmUg
/4rgqsVAI1LB1pDZia1p8tg6mZtNiC7zOgvtQ2+1DSdCJa57n+Ny/ciRlmwErs5y
wJbctmDEtPx09sWgrkYCBDnAzgAIOnPf2LRkq6dQg6uVgO2NC2aSNG8qESCXJ4wj
8RdpyZgenZOZYGYJzFTYI2sKObG7Rr7xUdUEQbdL9aa3WCcIp7AGVCVWyYBm59lG
n+XcPEdQtmimH9ovrzGKwj+yjLo2b6KTSC2hpnO65JBcfFYWkwzbW969IQhtmAmZ
kKGZUtWd8nWOX/6xYh3TfqHxGYz4mHajHSbxxlWhOCY8uCVdJqPbf7fqai2Zo9H4
v36mojFruN+rq0MJZJTD9iWT/f/7XBj0sN/G+8LzQ4R4TTcfDJhUIceKiIi0DlOX
/ZjxDLTTY/czPEEka6viRRWMUwx5Xm2i0QgP5/vc4vndCi3HS0QSkUE+3B0UQpxs
byY9h+Qq8I4Dsx7g2xJUjB7gi29TgeRSCm5otr+7Zuv/EI7ehXHDoq1/wnRzJ63u
Ih24NwkoOiLPEXazqDqPVj9NJqw+cFrzgNVqS5juEHSfGfLNGeqsJOKxaI9wJ2XQ
JrLSpZb4ykG58wT7tfAochPW/SnHlcF0fjpczuJcE5ZCI3+NJoRqr66IL4xAePoG
cvBoClMhsVUXUN+TvErlXC9zWqSsB2ClZK8JYOLUeKLNCDQzKRv3l3HT1h7ucFCm
pW8fe/wjRdBzq7XZTIItDXNMEMAO5kKiXn+vEyHzUifFfKzVvHNmyACJJ2Wg8DMv
agCrJTOCVhq8jZU+CqHWQrCbDJNq5Xf3q2rHORf7SdW+MTTgveLVFo/l254V3FVY
Xi8u0wA+C2it+twRXyo7yj/xA8oixycKeen/zypNseE5+eURDE42YLHx6/zbEMbt
GEXGfwazH/muuftoKaCusGNGiYNGStvBEogpKKx9f8XivGyO7f37fkH1GxA+aH98
KXWMC+sTYxLsCADcfhz3IVzJX1CCQT9Hx1rRNzMWoGIfaVN3Z+rrcftHQqLt3v1U
haSMq3Mc43DMXpGNxX4NZMt4j6o7VWDTuvSH8EwM9tGfYKvM6f9/jLwrA5Tw9Lyu
fzSpRVmpIHNNQQnJ9IOqSrZbd+HoRWdZ7FsRDpj3U7V5BGNM8DisZ4BQQN1BRCLK
ZpY8ohqef9jq31KqMbIRgS5tbDqjJYfSxUQoY109juVFNc4VjzpJwSc+C2cFnhLI
HY0iPWBeWgv4yo8CDE2G57NnY5cbc7PC1rMEcZBc1a4NK91wCVAlGZDgD8OP7NBw
tifwrF0haCumQ+RuQrUqRQeHmM9tQXlJIokb2r/VERG5jM5gryHCqHXS76SObSWk
SHisM++vLmhJoolxNreNtbPSqNsQjurVxwwTqv7YPIEM4VZNVhEbcVIRUcRFHPAv
Vh5kLKSCI1FdshWZqca1jFXlkxmVUzR0sTPvBkWIp0Qb/AsxeXzWvWA6kK9zcVIT
BEu+UagUurGQsPz6Sw0bfVOe601/VHpNh4nV70XDVn9/4mGdByp15Ft7//I5EsNq
rh5gAANNnd0wXi2jUijRxHz85mfDiVGhOlHYBiNQcw1C+IWdBtyPMA+PNP5ymFWA
abfCW3V7lWPzuZuYPHGSMpt7SBRcR/+qJDgaWoNwMaVmgB8B6QYQo7Lcvo6kLnw/
4aR0IAl4+mazLJ8jLhLNgeOyx9/OdrDBTFt9nUIjAtqbJM48ZiKEMNejgj4AFraq
THZje4VIdZ9MpJwsnzSgPcQQzFiPUVxjMcwAPw5nuP8dGxvHu8Laft5ZlJ355Ze7
xCJ1Mwmc37Pq+vixGCPKX9nrfjX4e+rTYpaLyCSGc64vyHF820oLYjU0a60bWc78
iBJLyC0krXMO7bAbqu/PnTkn1WFSTnPwlBhVXwwlf425J81A4mpAu6aKYvvCPZaj
4NFuUFWMST/80aruWcUETzFQqDCF+IhdWOtWVSsCrrhtAgH7KMFpCDGXhtBjSHdf
BongNF8aPZEfNz/Qf+IKEyn8Wgo9W08wav7PLLd+v2sIkNahLtTTM8oh0BxlBn4O
j7F0GxYqjr8sdCsR7wfNuw9Uhh6dNDyQ5T//mWEEAWRB9ah/n7f1rzvODfsQIovf
mGVpVGo4hAZOMPwiFMX+qSdMbt5Z14q89on4bLhOLTtMHX4AUykExnEJ+jReiU70
heulQaYxzSttbXn7wnABObrO+zX2PuMkYUygx+krM2ks+nIpnbxhZH3/5k6Tv/NU
r1lj8bEnsB0F3D1+PWvZMphhdHRA0byyiAYsarBqnEsrTqR4ukQPdVsIigTMhO9u
2yXGuCgEN4LnXfNz5zYTKLmxvNWBmQyfbJDCwoPE9ToXOw8va02AOnfI3FWm7Dv+
J+R6aEkTKAViOq/FPX8kNOpqgHQouRnyZKQSGaWIC9aCNxscrULrgBHnbnJFzb8B
yvXFirleaVuPphuiGltvXW9U6Y4c/utVCEjR7sNfjCGhQFK5AcPSbCxTrf6a41gm
L0lMyzCCcCmexj2jDuyiCnfsmBVZcXvavFuGkl4D3KZK8D+fUTavJK8kKNgGNYFP
mIa4dsF+qVO7NQ8RLSPmDqTAZ3+oM0DVMi4N4l+u57V11WzfYBxV6Qjmzd62tv7c
u12vaPuWL3BJ61EsiTpAURwevhzamlgeaeXGv34UvQb87stm2QBvACpTpqAFSp4i
iXnUpLYPiwk8qQs1fy5BcRz9wxLvIhzjr8CYNFDCmmOpk3FJbvWCgKcYoWmEa90S
phZ4LSTpqNxGNLVTiKVPMyRc4wovVvN36mDC4Zgu64BaddjJy9wNVmFCpEJMKvjv
n2gtBLRdbzUHhz1cJ67kXykNL4uLe6mP301jSclFztItpyg+zdDhisvYijsDmzvd
JwMmK26nwVqbQmWuPOa/Bmdu0xcCSd0IGnNxz3e0qyJ1NMfchoKZj6JERbgN5ufX
F60o98oXqdOT6BgRbkpw5WPmtgtY7kw1uLsqmVPDvGx0LzArwZ606aCDi7/CiIbI
kUJhJke8tTUVE5KbofRmjMmsS0RFBgFwkfyuvzTCDCYV07oCb1MrXx8pNm+Mysgm
0xiHgcvOBU2R+8IStsbVCUz4mGrDyZThWS81YoFgHsJsSzxEqJCRUy7u5CdIuZSO
bnzYiVOuCk+WQUoF93egeP9tOR1GNcvUsiFCvUbstH/P84DGeLD8yircf/PzyKb4
eKqHhL97OxTNj+rhi4pWAgvnIth2M6ka5LUU5N8AS0ahpFdq09+iYJZJscN80Xov
NLDjf+IA8dqNvqy7WIrp3sNcJmCdtt2l/ZNinIErtdCCjsS35yJ5XH28QqZVHAjb
kEpf2aqc6WdDio442/qEXl4UXNhCmvX6Rq3xHMkdGme1fv3ueFejPrZJ9U3Ln0JC
2qkXUrf8rTHF8x7FBjZQp/skt9Y1M5agjjfm6H2VFRo9E0mLcrm9r2e83CJ/Wbyd
+Fz13fsaJgMHR6YnmOSq67mImvjBeCEyXJQ27V4ofbihMXEViNyqfgrfoTr+XtP5
k8Evw6UJWAAPhu8iQCcu/WDTCY4c9EqsleDeq71nIq0BOEHEo7cjaSndS/yi7fXn
N2zeTjqBTY0Wv4AweV6phN4G9ddvOH9gH/fYBbxDubp2mQIq5wYI6T9GMu4oLP79
dpcKhQu574GAqKakPoIrp3G/0rDLhsIc5fSw77/3FX6+aQRes1MmqIL8RgZkpSNv
BRcIOmgWldkcTVO0ytLM3bCXQzqFbR1zV3CHA84cj82Dyzo4qqDGQwUGSiOmreA8
E2dX6Ns22jDzM77meUvuGWBZdCv6LBDoMWlMgRaH3I+gatjnZ51IAHKHVmSX+PiO
B+QoyOxTeYo8SnWDSnPV8RjeNw/cmKM36Qw4KbfliBTAKOJm9alp7r9xmmU6U8Bj
BEPAe/SawPDCzN2COuFAIPFaKZbl3Y3zBH2aW9X4K8WVBe9ttljeW9NDaK7v52kE
jlBtu9FaSReT3d1N4kBzpNqI80jSQszF/DMTAs86vSTsAF1QpIahRiPgMqiXCcYz
6sF29jq88E0cezBgqjl7oXrPgxrndY57qXr7aJBsxQr6Uw5pL44FQGSueXSlDzsQ
gsX+so7qGVFpvZhABkphQY1k/sWxKHk7XXat8RyAbUqKSqvikDNL5ahQe9mQeejF
o8a8/2XrqJuZE0bb3KB+OmrV2FuCIfKP8/VZxuD98nHGZywHZriwWgrmN/+9dkoJ
DN9oQkj631dJecwz9B0ZeEufiFYFQ17IPEOD0sCtQKeXagF9F7xTvhhcBxt9OKri
GejlVuqyCDL5mgMRLyr3iZgtrcIeWccm2DreaBrmUGOZmln/twEb+vy52bIQw2u2
JtrV3GPM1WBpXCXP03sWUqg4qzkvZYI17GESrb50Jy8Ue2W2Qld6v1mLVf0kkqef
eKdkhPzv77inECXwJrGI1G2RAbXN/qPb0RcYrqSgapVxY1OPOQbm/uUXdIUJmUwe
e0Cw8PIgw9mdSK+pLFB5AaJ1ArgyjSpl3bQbshcSRPqXLV10+izU7rDMy4F6Imr1
3MU7XB3Q72fj1ozAFgSPNQCpTWTQeocSqre32qRYYiAPrGWzRXqv4EA7stH/OIaO
tzthKB05WpFj4gBWuGy/+vfu7KDe2dnvSC5eYbFS3qS0UOtTGcyVRPzmxei0hPRu
xN+8CHR/XsuwoIg1vwyN1S5WUFqOLcCyvrPkfXdMZzVCMQZK2IM4zzlBTMwEK0lB
0wxwU0VADUXqqOJVHU7y8A6AOShu0IyEU86CDQr/brTMiLJxOxyqAJKV2DqHhsoP
bJIJ8gP+P8cBee6FbXYsHkwNpX9CA/j4gojSoi6OSbYjAi5pyODP9wtPEKBbyfBS
PXieq62jJqO5EEBOWfc9Rn/82YPopISU6tOma4o7Zd5Wt3PSh12vtkvlWz21M5ig
xB47e2R0V9tv34NlKttkv5l2v+Azs2A033LQ600fa5B+xIoxIqAqYUeBkkrv9wyk
axL6zDN7m6+FXVwXEt/x4IBg8iSMPNBBJA7RP/gQiIhfzIuv1dwB38+r3ZwRhMfQ
EBvDIWRhCkWkPAddjWnFTn+YVFR9SffOSR/yjK5OBcoComcqQd2LGppNw3vXRW23
1yEHoOugWDDC81u2VfCu8RPenzZO2KgDyuwynSYpi7ndX1iWe+WZXjAiV+0I3+8i
rLwGXIRYfNet8QN+Jdr6nGVsc8RWVopiqgbysLH9IVr7GJyTc5ROJGk51ArctIH/
SaYyJ8SuSb2wcl1D+m3gbedFxO9r/EGpXIpgRIARbT5uYOcKtgPwbC+HIjov1qJQ
KYssKtgLrnhWOmfa+z9SjajSijTojzdgWYinKxQhL1CgV/mVhsvSJ/9mIkSi5lY7
ACxmKAx/Zf4kxUZjVCbJm6VBgqiq3YnuLTWvIwAGHv/+FGd2q5NCfJ1kLx8pONiH
9rKRemgMHSuxw/XlmLkXQOdUr7hCallK4DL650SxpANrf2+e5ljnN7Aqw88i/+UT
d3e5xpHnhOR+c6ZHScSrz4oLVZZLl9XA/pINk0wpA4bowRe57MlwURuj0WQtE19l
NMaN5gNKko0kTGag8qLJ7Kq9Gque7OPCNZwxYvLX65jsEO6ifDER9VQfVkalEnDg
KZB8wEtkPjY2DEIaAjyR0XdCcXO2FiMGmd9wnUbU44UdDLGmtp6TJHT4Zg0lnLsT
oDD5U5Hwrj2IC4yHdhHeilp9ls+Utw0bw+xKpU6BDkkJvzwmP44vLUXEzHdA7EdS
aTv4BnU/nwxFeyofoeclnXlQllyxGOLa4XRgG7zcyCAJwZuYM9H6rNnRN/OSihiU
ZnqMqQCdWA/vQg6axET4GFduY0DBouhcv4kwd272h+9q6whcugNgGbixIQvTvIax
uUdpsxBDUefDJGNpANHVbQlhxardbS7BNJqSbLLkwRqWO9v+uEJimS4f4vfNS9lL
jpmmP1BvUtQPYS3Y1XMINLQJP9OBBeV9DmFQ5VbGxrlM7XgGWm6/SuHVHThgdENU
OSkkwxz7kVQJtAMKYEQI51/LsVZTNiNOqgdIWzm1Afs5+9t9Wbm5Qm7Lta/W+rrh
IBXdz24Tezrt+zTNyoVNoKy1mg3o77NrWURPU/ZcFsApzhWpTFsllohrycQQy2ax
98DxTU62d2B8fIiR5pUNq/iA5QjWh8m3rxJi3IL0A9QiPXWGRDWX8KjiHRQK9eYn
qrJDhmQ5cKEmFIZqwKd3S0l0CcQ2CinBodhBIc2812SqxsIID0AV3QaMIUOlVqw+
lQ38Ra4KLLSad9Ixr2yR1iXEuESS52ylU1ilalKqRKqZancB8sAHUaJEsTbukRLc
V7TbOzfky2r1tzDetSLvaVEfPgjjEUzrgCB0/FAsIY2R7kYtZylFzAWT4/ZI3yvh
KDNNR/jypPbe0Wu/V5r2/UdyUeMGU4luuKIrzck+oavObIWi9zP1sH7MgEjT1mXZ
PBpYh5VCsM6HL4g3CppzZko0fFE8ZuHsSaR/ns0/005i2JAo7sm9dimen1tgOTbX
OmAxOd3EBZ49Tm36UVABqh/lNZ/1ujDqEbU9QrydFf07DJcCDEUnE8nJGZd9t3ir
QLHyHDADWltbv8267kdt0tBqJdPBJxKI08Of10A2nqZavFVKBFqNIqeN8DCUkYBL
6xsdtcVQtKveK01O54ONu1AwC/OpGQ0PSRRmdDkTPjnhsNqPXGK1xV/V9A+jFDAp
q6UclZawsSuyaLEg1MUXQubTji3ysjISjGRFJzuGl9sDqNFbXper0UBrkPjngBQO
q8OmEKLs73/kcEuMtDwpCoUwsVpMJZaKuixAb5q5behHCzSW1NsvPb/xy6ssb5o1
vjA9428CDFOv56R/6YM/34xweWMFjdmvA9VGVtR48i91CGbaa6xI0RgHLiqLpdic
5Ut+SMtf0hmtmmKSxZJE8rGugM41pAUegByPTr+cFVF33w9QY/bygYLgTxajBLLK
w4Wo9H8bLJxnyGjy7iSzE16t+sVbmfHxsMz0VU8fXr1bI03o3DFxqQ73lcYQSN1z
Rm/CYEr0E+hHv5rCHpiVCCwsWwTcVK+hne+fwdY5Qhx8biC6J6J+sN2OV6qjyQbf
tPSTzwehHQ/qMRPy16rTeGa0+EyL81TVWiiOaFRiSMvnE9pSdxpJqmEgG40FSs8b
hnwgI67cuFOiS79p7Tm8oz87CQ4bZ2pIXILGhH0XginCpWFph1rEDZjvqXqjntGX
9gfEgLLB05CYKj5Ptk+exDx1d5QR9vHuMoglKBo+tO+2b9VXUR3TKlWunvh1HtvC
qCxJGYU7tKfQjkLVKoVY28cGczNsq2XomPxonmPsJHJih/Ck2J3aumy6DW4BywHo
J3RFn3U8M76Y9zluTugBx7OTI3do53sAt+1c5cq7aixTiF8PwatQ8o8xCeb9uL8h
BFQwNRmr3a4iqBRAOAsw5mZY1lKq15t2ewNGJUFHu/vzJXMHC+tSI1NQeL768/lW
25yroJKcZLKf9aE3yo/aSDjyajSdGkf5sNyUCITPwR3U9I468w7ToEd18tYue3X9
1/J2PhBaegoIQSEGCEU4lno3QZxO61JT4fuoUlsdBtEO/I8/7OkJkZSlfq3wBxhi
hg15vl2v06YLt7pFSX9lFOYAlyE+wTiF8WOVt2oUzzjSeOl6mTR12YzphHf6Puw5
T8tpXKj3IsuZnPdiUEyeNg0qYRUc/dPWOpt1hjpAEpSIg9crjBGhhJkpbmOM0F7N
PgM1J39+1NpIdRWs1/r9W0qWU3JufwJg0WySSDx++Fv6cdl/OLrU/12QNWz1pbhM
K7oRcbUCP+4SotNHvPOSZKzQo+iBGaAfawmUqfdqhK4w2M6kt3yRujVGcHYGaTXx
lW2ONQkJZliUlEXYqapP4C84uoQa8CrgNlaHc4lU2std0XmwsLu7v7RO8+IUUvUk
bJTD+SvlmT2nnMjjbYqJfWhxggQr+vvQNbjgNSx3zR6rrLUFsNhEh11p6sd0MvB1
FR4JSJapoeBAqgZK98KT05g1ladtUbySLdoQzdM067C/yEJftiTEqjPh2OKidaxw
Yeg5TyQ4klUyE/UkYEcI6isDamaG81mSiyOhU5tM/UrC3oS6racx6Fgr+dG0Mxm3
OOD6f5Ps90dYKP7piLXIp5lBHfQNp0BxIenFThjc/br0GaysmsT+/A225EIUd4pn
rWiXx2pBPoSH1RBZHozJyTgmuqflC6msYmsO3Ejt49cT8r6EwjZShU9qBDW91N//
5Jul5+K2YL+dcPx19O2xkQ2+2TCJ2oZEksFGYiPFOl51pxPNIFPT9iJzvtzvi7Qm
B1wWhBEijNz9NHBODwctUqK5O8k6XHT2qDepEO5SsuFf/ySrUyD2OwCnpPpTs2X1
NX/EqFA2bGhmgEiQx2iJBO55DLHyDhJYAbJRhprjqLtsqsJza5fZ82gaXSnyoVgV
SQ3rS38SkyAJe7rkUnpDszO8TNoVs4J8NjqnW2mIuaFmxc89S44BPCUFS9pgSHP+
FYql8q8wmxW8BCIDRloftQek6g6gJvSdURf0Rlio6WRs55Lsh/Gknh0Q4ryCwCWp
TwuStrUFH7uYNShcvrSHRxL4c7di76/agKcxJJX22zzq5CAHZLsPnmOUVCVWehuT
U1mssC4os6WejL2A/LZ0xdygHLqzT8oJtX32q1JkSAeqxt9Od2FXufQdIjewYUT/
g3cQlDnsA+ErYRBpGXez2/TJJyOwkHBq8Jsw0rqsfqEWP1SSTbWGhOblbVYAKhIq
xBaxSvQgsvP19qo0kGf6S04GxHdwXDZHZUB1CmNCYPcRXoa0GUOEoNlOgIdyVNTL
RVOKYcSeptSAuoL73HSFzVfH23O2iwvPAKfd0yeubCFQxNi4sajJ7YF1cJGJ0Jlu
K6MvM4trSQ4rdjMK+ySdd6Z1J8781QkRmCv1ewxhMRc0mXGHop4NBP77JogDOpop
8uIBDQ0+8zTOZNDlA4NNOIITKxveKorbsOD5s4YUC6pRjojT1J98IrTKknlSe0x5
Vcm4VdiUlRkr+CwZYv1j786St4ZEXFgXlhoaDUKhyh9U5/CXhdkTo/JG3N2UWSyX
Y+2FGXaTvRBZAPxyn84i32oF6AWHtFiSjmcRM1BRCUcGLsJj1BZWNuC3ELBHxuxn
iyjmBYbM9zG5uoepIdjNeN0Z2nolTLCN6OAZIHAJWTJgv9ExPnwWmGWKV0VKFmAV
/q33QAYqYthaG7sI8o4vo+JEX2I0KD0/HLU29aCVCWidnFPl4utLxQuQENMq6OC3
eOaFypc29HLGsDFG/Xtl5+C9WDCCRQ2frygHddGIT9iI4Qkd5HfW8E3jIjxwSD3M
kuxInQIzfbYoY6CIDcRexxT4uS4vVFGxVUzFstBDf+qTrhCNWpRM6GpNqyxOuFQN
unDoQqTWYnJYbbz1In+uDW7ohxu++EGh97hCdD3kBfT+fpsZow7jf+H00XdjkTTZ
s8k56/xbQEsTo+UmILwAvnCDTd9tilnGP5eS20QOFAkEkFljuVV7q2g3LjRjdXsC
0oQ0Fnx3gGPlHdiFVWGv2oOWdAb1sGmO1fu6VIMmGx5NVKEcYaKVrWFQ1Zqk+meT
BBkF7uwnoQMJaJBiVEb+f7Vq9l3bwpxHqs1xKB77ZzrnSkjN08tF+OLicNFT5ljp
o9sGRICwYfKcp6MwFEkgtitmOGozXEDunFoRXn9J6qZ0HR22KnkU3srXf/tjLm7j
NVSIunpov9Mxc9gUSld2kpEK1OhRQzF7iz0cc04JoMKDiSVVBit5Mt2GS5NhYRz3
mk8IYGzLDqLdd0RP/6Tmt3b2+xpyqA38ghIkP8yP2zzL5aGlHTwSx0MvriBijPPy
6RnwHbla+gtKnC0AXmN5r9/335xmdM0JpsNbMmanb9qtmDsxHsbIsFlwV/KJkUdn
si13uPNLSkXnPeTMafvytpEl3wDWOyrk/QycXPVvrWqbOSKsn8kR92f+OSvAHYj/
u2bC31SBJVZMfKArwHPNE+0c5ch36TQDo56KdZ7d6B99bro+NRGlN/scBAsFNiCD
PqFo1me8Vwv2ekiv6eVtGYWIoHywYXjTp+c6PzSYSF53Ajyh3WPoqgFoooCn8l2q
Kb7JG9Y1FemANdGXdfGu+72YiMv030r26crB9j91APwL67iFvmm8OdKMHL8F0hVL
cWeqxeYDaQfwRKg9U+a4Rrn73Ca3CHo8I7WwFoFWE9izfvpSkKhuLhhSkL2LNbtH
tThtSKZvqxMlmSnNGPOISN2HMPZZ9TZ4nrz49E9VMDHFs9aTRGXWIqaLpab1C7uY
lS2SxUH8/O5p4YXjXlaShshp7XuG1zCUk7r7MJ51PngaGpVD5ts9r5ucF/jCsqSM
T9mID93zvDDPciu4736APg1ZRSxRjVArgtAR7xoHFmMZTuC+1G1WyUt7yGx8uxvv
4vBejyydF6Rto+HvFd+ViJfRAKqYqpm76POSWaJLPpEw2Mnm1MWOBLLuazW5Vjsq
dn0uuqL9QiBYHWNmUroOsUlzC96jZyco0JtYxr2nvuTc2sMje52TUwzwEo/lmboz
tqVZtUus69Trv8Jrz8d+1AazcaFEmpbMYHAwmsFjYbeHiCRoPwQbe258INogKjvl
n5nx+B1FHvaLTz8mgzBvAnAk/bIsMndfKLfHG4fXGZwhUUKiKOdp+aV3z/pZ0kQ9
mf8blQnYLv6YFtMR22INPSPeNrFMfMURyTPPlMyLnh/oaOYVgwQuuG9TNvEOqEob
I/IBjw5bVTxDyaThO/kTvhv+ao9n6PTUBcoa9OMisJjFWslvhJYypXMkX+v9C7C2
rJw8wttZaXbVZ4DfovIZ0L2llspaZu9s9SbYmcMbqXXxuahmerrNKCUXaE7gisas
N5nEEbyiziYhmU72cFebZ2jsVawSts2SAYSPZFE0wQHnsIJ+bZi1LHlLxTd9FkgW
S6llTcVj56vZoXylyxit52+qf97/aoLyomxyMh9bpXda3Ues/gi/1MxIaK+ByuXu
8ZXGOuFdDc75ovFYTuqKZQO6Xrx/pow1mvtcEW3ZiIx7PTMDEOBxCUkW8eHFm83d
aTuTuqqLTuGbguojijuhpO+PgW07wJhwbwnjrYtPBCcGt/FImrR1v+9sPiS5O5Vo
z7h2Qt0fnZ1JKJtvQPIGfyvz30N6dtfH7SXpb4KMKm8T4Gl773L7se18BqPS5JwM
30r5/mRthTTF45ODcWyjRcsIV3v5uqdSKRu0jU4nLiXp1kZ+Jyzebda7XCTUgeqk
COytehezhj/63lc5m3YO4jNCL8H19IRakgke69ZcLsnVLCRhkT2wqC/k4dwJglOR
qGcKXSGsgJ0zEztE4zH/fN54CUCqm0LkHOwIAyUDfwTO62G7znu8CaQ68L2cPZ47
H0t3StqZnD/URF7r4OtnpWVbbOfpqRWCWQF12iHWmGap1pFrgN5R72Pc8HiEm0Mo
i2vLtrhS7GXSjzdO7yYQ9fuLN+gDl+oDGeLTx3SDoprYdccSKZTdIF0tjvpF+Ic2
dUYO0V5+Uuh57TOOnthnTRNJACTT8MFCCMMMt5tm9WZgEiku/U4alqLNvhPCN6MR
xqY0lT6H/ZEJvDD5ZSn7RrI39P50/h7RUVfz66fMQj14/oMjKGgoYf+FwolSenb3
02ZCSVrt9prZMXaARR1m8ZOZJS2xRYkD94K3xNGW/Gue/KxbKh+mJXUyfjypC3QB
8M7Ch6Eb4PxB5SXq7lYAbefob4uTPNLx7uzqnpAMKnPyA/3eFn30IUkIV6wdke55
iImq7zslr/5rrODCNLt5qvW1yA7/VA36qwpUIt0Hxqw3EL513ziBxPGImRFdzkcS
bcDp9e0yeJYoRnssaeqZ/B7v2TTnVfi+3A0/TD+Ho89Luszfx/LNP+T5JwmI73vO
W36ArAtOWKihmKQOH9yuHVhUj8sthK6o2CX5+aB+l/stIILh5iUJX58YBJfTq3q1
CC3pFQ+kLSssGKMsZ0foGbENyRfZ/MfAc9LRWgP1IbkHeUnoboH1tfeqOvVXLkNV
jN+hDdXV3dB8DC4qMeB6Y/JIkUuwwW2DupBQLR6jgeWJC/gE9Su+8lBebxrZPDbC
mFUy2t8i7uxTNLbnyZv977OmmD302WYL4gH8chmEXHXOMKmXprGADg7QQnSFPIg4
XLb80rFtB3H4zM20Fd6ak+CGieYsdHV2akXqEZBH1b+Rxe8FqmDYRVZHltOebdn4
9nnbn6FUBWjPoMRoIC2Qum7eQXAIkFk3oAVvu5oEh+v+Yb9Oo2yFmTXCZnSJniaN
fs8euDqu5iO5pN/e9JMFJAwxoAz8P0aeO0JgIkHO8SLr0BFocymuFqN2ck9jiTNL
WBl4lmCmRsr+Aa/kNJfBK9KEUls6/OxqzNJxQfyG6XOLJUkOg7cUTIS3qlP4JYrx
9UIg4ax+s75IP6TdDV5Cw4ud4UNPftm1LcktfPmz7oqWcFf4jS/tUT7QRKB6Ge6x
bNEKO3cLfX8F3SqKivu0vpi/HrpXdTzk535YPcB+Gfqf0cyROfQRIM85/5+9EEUo
fyEJbYJyME370cb6uURzAtqcvZLNtON5IfOYS0Upcp27FjUm7Bg8TXXfwA0CHXpN
nEyg3MNkgOTfIeoPc9KbrMoPKvQxVegdB5Nyu70KUezUBIqmoOX01+oVnLP1Lh3N
OsHXaGgnftd++X2N1JrYTnweQuLSh9Qc1f3eivKp3lPrBSdzHSj/a0ThmEkqMeyU
lhNz1Wm4wQioiUWWO727h+GiAMOYonvFZ5NboWL+hRH0OMsBi6TsEZyaaM9+LxxR
L913WyI0vyLNafZx92+O/5K2son7nuaYhBicDmLBmXs7iEh3cOvDaUxlqz1Zdb/p
F1xXurVCGqTzTa8WssX/IwPad7qE1/4E23qDQYWvxHK1RUFZ6PCWjz76I9DHvq6P
7EFSOmsOyC8mEe7pyGSqMDYICAkOVyQCjTGZVT7QxfSljf+mh+1rRxBQQVHQ7MZT
oJqlz89MHqChnbtRTKmEQvkk6d1XNDIWNgrRVlzFVnGluVAczeY2N9dtUKpEp03H
zAhixiMeYnMGLoiE5ymM9NH/CJKPzfVDNRib4VBMiM4qzGrMPFGyMYCgh8mH3E7t
G3ZzhpmYk/QroyVCCmaU/8NWw7FszZ+vv5Up5zNZJQ6S23ML6lwqGRH8scOoxMlm
Lpj60HSXYQqecU13U86gcc1p0iamCVaeR63A4kpBy5MuRT5+d3bEqNm21Fm6klre
Ghlyk6XaOBzFlL8bfXFEhQ/HMcYrTgV8p/s62J5M4mHlKfr3mXFukkSCTxmu8Ehn
LZ+DBG/dUoGT2fHNx673/b05tN8omx8yWG8IOUR3TfcYrxNU+YGxybN6S/0h/YZF
2bLV7zJf0uC7lHxV3s755gW8EYkXj03SThG/E0KfqZVw+XEz8UVfa4TFYv0/EdgJ
rj2GmiWqOfgN9oTRCN69e8Pfq+W7bfPRw0v9zjP28dZXeKM6yFJtmsyWSrqtlEVZ
bdO623QXGstXyXaytmk1wWrq6U4RKfeXKi6WAEZYHGEaAEXRl8EbR91XzsbM6EtJ
8wN3SJEG4n3w3Xxg3H1Hm467ZTK25X9pcNnWfCG7xRDL9BMWv/pBFQPbSQ8gb5Ib
7kJ5JvZ19WHooJcP03xmLJzeDwDUWMKBC6loynHiLNT5HeqglDGlTMuhX5LNmiDl
mYm+49s9qvVksRDl0Z2gS3vEcZ3WPySAXo1TXfkYaXdKj7dzVVeaSs4cznmmMn68
85qgN4rBqFH6yjI5m9WEziNDbv72oSUhlwZh/fJjDlytkrsv5EuKDybRXDw0ljQT
aDsT5qO87s1GD4dAt5Eqv44jzFzsdO2mjzaryz35KpeXsnnF6wM8qWm9jBWj9uPV
8hw8O5YuX0EwcLajhYLTUqzaVtsBvNTxWDv9NFZMx0cnBRYgZu3czMpaqMAdOhWu
ZHC7uRrIZQ8WenPlQ0k3S/lLext42+RLpH60lJjwKp1v2HMaztfBgPR+aragfYVQ
p7JHFOVCh8caFq93Dlp2aD7lSUoYn0lwpOLMOTYUnwXvcefmkfURIMtWJc5kBLoG
rRg6rsm+ieLz5OVPRJ9kkh6nhISpPhsTdd42RmoDMhqXs0xaJVyRkHAOh3RTvSt0
zvYpHAKgjZgdeyXOVuySYuf1n+hIIf5uFJN4APQR2VxgrayQj+X5GqhA919XYGx7
mjCj5Rv8dOCwSyXkZW5slCYCR8sJCff3KA+TZ6bYVLXKD5v7iRx/7oiJLD1HOXqq
0JrUap7p0qOHpZFNYpCXMNetLjRiUNrQNHwaojp9NF651WDoqO1v4vk/Y27VUek6
2oKcvHFWRfTMaNp44kYaIHmZOu/SJgqz00xlvjvxZE5QziebAjcbvCS8wyu4mhe3
vN2P6Fy/QkeTXs/NJUWlUafllSJN/NFpNNx3ie1j0kmemB2oGhzgvr1ZZTimjh08
yusNsyIe+2XxFIWtDsx7AbniLFj2NcUPRiPzb8c3rPUfzRCYvI1CWpIYfwG2Q6NA
c8kPxV+ki042g573Tmgb74iz56iaDOY5ccAYQmiUr9hk6WjMyLJKfQooqYVDfy6F
H91/LE6r4fWaVXS4WDhmcl0WreGK2qfvf3pwAIhO6kwr7uJyaEPWEP+dsQJN6en7
wP69p/EMvN2HAHTmsUoFxHeVH5ntiYCtxJMmljmJdkGnWgBKZvJsdHcdF8odqiuT
F4cLWR0aXiTtwdgZc1ptdXclejsrnRo9roSCu1MVQA0WdIzswjuNiiw+GwkOw/UP
bJ8XYU73QnGZ9yymxn5TeLB3y1rGPSoKDNYO4SS/iTRRQ4jubfrAzxgVXSg9GiwQ
wM3xpUmJB/DcVSKp3FctL3rlXF8wSs/MzU83CAq5dusMP/TmPUgKrm8GQfM69VM9
ca+sW8EY6wx2PmYQX5Yu1vPMcqb824wKjPBp+BIM+LcNUOrtSTzyVWdwrZRS5Biq
7AfhiM5pHKEWYYw5q6Imky/TZ3yqFGdsEKBWGL3yQhA0I5Wmuz+W55Y0omXCRvI7
7xzml4E0xBKpeznB22EDFWguQIYg/w+Apu56ECeQspiVLWup2ruvaXC8wWofOmfQ
4l2PLagW5h07R9Oha8dqGNxmxJF1p12+tGKkPAXProxzy5iy1+Y6UVSmvNw76BzG
8RyEBD0WcovQWXmHLytatY2kA1ar0T8h9AmeHB1Kh30ROdvvfATBEFPGMmMcyR+/
Nl9FuxmKdI6QJYeaudfM1PrjQAMXI9WMoMXLAON66UQDPsQ6ZRuYUXyxjhLSUj6z
5XkZOMBeKzJbqSbmOiljXj6elbRXgtIvr/N+iGAsj01rrYVfDAhYBmi8Ze2z4CsJ
mGsCDDkQjgcXXQxYG4JafGbfyjKbpEku6yygqDebRSnad3ee1M3vhifLfQKCF9PB
nLI1ye7+Guv/m6aXEg2d/UexTcnE+pkvXavTzg92GDyM5rTHTjaWKuBlptS/yDfN
pQbfIVnzQky19I/jsfeIjoyjUDijJfjVnGwC0shheaVtaq5UMFnzztBnfjeMbFl5
TCvKJb6RwVvvJ7U4jfTTK+tHfA7jVaCLd5eaxOS0UYfPhqivP0sAz86vmzTC1Bh0
6zEiXIBN52xBsXn5LBJZ7GYhuCn8/EXv8adq8Fy3dLPyhVZOgpKvQQXAbxjlxKG+
glhm0hcFi8MJUmYOkAgMqIPUmyDPOF7nVJKOLQ6zB+fuDlhvSMwolLewPDj+WyAc
Ojvvro0i8XFiI1oNRkWOukd1FNfuFs9hGcNQxWp2oeMS7fM51ajuxxTkI8akP58E
2H6TLO2nuIQvM6K9+NxyoNpNLGSk2t6HY2iZwVaNn9h9KOCylM9S4FkLxQDa6EDF
aOJYYQ2XsNoToW5JsGJUzfIMk3NXE19dSOoMfXQtpfAzZt1iHxbR+LKJhkEoYGXX
aPm7q/xQw5Um+1+yVHJY+JprSB5+phvMvedeoghfJZhjOh3Janfzn+OWqhAXinGB
Jv02b6nXfaGZhOc8kf1uv6UodLEo/BOTp9q7/aI78HN5P2ecQGUlkelD64r2WSMt
z8E3fc2uY5no2MueqUntmoRBNXyjObjUIqONTQtktLB/H4Neh6FjjvfqMoq/EqA+
eQJ2xW1s6XX48Lx0mJCdCK4vn4JEOPK55eC5qjkhbw5wwFuM7umsZ7KX+EdrVGCt
KrLdAuk2XPb56akgEqy4nE7BwYWQl2TsF9DjAE0hgoeuJ6NuMiACz1G9dGD5Jmsz
7mPN2Q7YQTT9YuwNBU/2l6faEZCIRb74o/L2ryZM8BmL93W61NBlU90lms1dnihO
zEQvpCzm5N8Zd52A/Nr9KKlTCX6JPSvMzqh7PlxZQ6mtxF8+RnS5n63f13BghrVY
565bdRuBTKxD4FoERT2lGb0dYMruW64hm/eHzvTZqtROH0qtKbKEneCANOKDLC/A
dlk+nutiIqEJS8fgwULGQMKapGkYeB1NtG3f2hAd38V11y1zVMS5L3jOa/X9TcU9
14wjvbhcErd5Rw6qvV5v44521zdaOfyS862j6VaICroMf/Xq6hMgGuQBH7LVMWOJ
XdiNH7mE+jHKhBc0YY4W4j1RK1H8xdfdjXvCeKVxofPkw6Y9PSrvLXx0I5LcUdXM
T/5AKlC+QO2+4k6VzzjqFQjtiM10RQtmSM1LXxB/nnOMZLEfM7fmmbgqdYVNh4Hk
mamQNKEvO4MYxDNXJ+5bfJUJcBTPFrtXb5l69PFvF30BHAfRRanYPjDc2ZU0ogTb
JA6RdXlOyeJBUpl67qB0xg6xGg9xlgMzKmWIdtskrzagR+UcXzKYYFhXr40Lh5bx
V8o1OCk19BOt1WA2WSF+kOcI5j67ziIzpd/ULNazZaREkD5u6P8N8I9w44c1seWn
vTDfC3+6348Q78OYTIz3mPFQmUvGeHdQyaJx5QtcYX0Vgyedszp6alzfc+KjZhAb
+9BQ4JI0FPtqnLBffgHXByCtrC+XsMRp/L/oas2j3Gs/TjRz7MR+yVSfBuafNHYm
SMuVDaP3Lba2hFoc9AHJruzNfQuBxfEIq4P8VnU+th3qrz8YxaNOKGUhmYHgS2pe
czpWvrJObykFtx+lt2d8s1zK4sPeVJZWgR1iVYfOwrx+0Ngzs3lPYE8AC+7hZORw
icKqYQ6LehjERKd446MzRS3Ty5e9nDBowekB/99FZDHXl+rBsaEcMV4zPsXY8P2T
p1aUP8KoGnOlWJ9bLj/NC0S2MnULg2PjLf1AoxM6h9EaHGfGyrpeuUIJB8CKskbU
TwxPX+FIyxKZgHcZ+zb/+sFUByW4WyoncjswTMSJIvGL4bQCFoxbNI9yqO0lgceG
BWNHRreb+ulIKZVTEU78Jqy5JR8/i/YEJnZNc2AjtagXCZmz+6bUOlKpFQI1AGlu
Xgk6gLp0hyiDtTmjg2O+knyICT46iXykkBIqHNREnwCFzyu/q4vhBDn/Ff1EsMG9
wFtaxw3czq67DdAu3VA/sN1lJhubeHzhskYYPJo1saJMfnHU+MDzIEhJCpRE9pJ2
V33dQddjKxhZPiY7Z8jyREp0PFnzbPpm5PCSkY5z/gnBDryimWlNkZMS3M1zlVbZ
7HCoKM6ffZ88BGS9VEArJd5y3xwJW4OCXxlKybJgRd3R/WYzv7IZLkvJoq5In9A5
L91JC3ufb0V9kaWCuB41CBBG1YpF8MO0Eqiw0w8N2otT8GGAobaUCIQpVwPtqRG3
7JZ6DLCxw/e+kNd6+En0+1rBVAk8IGZXTqpLPtb5X3D8Qa4aPul1YvnPRv6W/z/7
/ZiMO5qmRbQKO6NzKKEHIGMYQOw0NNU46goM2QF7ShArkFChLv2RNRaezYR7ipT5
IKWb0w4hfI7L0NRYxOv2kae4Sq2BEPDwIlOrn4e3u7U9ZPRJ9TLLtofJSN1qFpof
d5a3/VXL9avCFHuZPBFcxtBq+W68wRKwpDs6e9pG0CxcfhKpVrvjrk+R3SU/8br3
jaSRBPHhJa+7ftBl/mN3joSG/9y++SJsSwQYbKIqjQ8ancxuIRFLJTZRc6+uxbfV
9Le1y7SjLJVOFZLMIAPn2u///9ohN9pHtiBmDe1hLWWFHiBKSe7R51n1P++MeUhO
5MeOOgpJrvfQ/1/f/ECWqpXYsEm14IzTAWrYlyuXwX7ir9zLQUPWGfcgzbQOe4Yt
Svt8BoQtb/XKTYXvP1fwqw5ua035bowxoNuyiWyR+hB5PSBNcpOeOYJTr10dBIm7
tpNO8sYp+AL4BHu2hCkGePF1nWz+RMdeymrDfNSXObBPxHJu+2ubRl+89W9E8Oku
gwAMZUp5iJQDfRnnQxlWILenhrkqaCp9YqhLnZ0iG/oagxbzrhno2diTGGP0YK52
HRYt1ceUgYRfgn7wI6YRKuOqZvlL1dUeCapXprzaGD6SSOGc31gLsrGKCkCNE25z
FUVD4aapfxw0V9CwbICwWfDNfFr/iz+0vmRAQmzWWWTopsyPWM9pjkSm6kjmdt0w
JN/Hj6vs6WnW/c4OYBiQBVnVMNEKCdbGLCgcWSfcELR6YXX0YeaaMkRzrKYD6Mpq
lK+aYjQlzWgUpcaSm401x9tRojNt20UWH3NIBBOcUq6pSlIn1WNaheUUYrHG+Ken
MiCYk4IDJuFVbpgr3bu6lxyIJiMaOTTVLwlJASQ1eI9UdErKQx1E9z7EskQLKg7b
GT0q7a4anQu4aYaJfVBTxQn0UnhFfmW/qFJeMdgXrvzNPumsG02wMfIza/RIuHjR
244dFtHYOk8QMUWSuYj/vScJCJPed8OV26YWP4D5Oo4EfW3gtdfkp2gU8Cqcwaam
dj/OewDjYSw3L+teKdKQmusjVn8/Vee8QSscBmi3pV5/Ogb9DCKIkgV+3Vc538WY
wwl1JqQHbbYhYeo3tsA+hkTNm/e8Mh9tXDp+w4cV5DLYrbs1+Hk1cIDoDEidakxQ
KNhAAlkxL3OfmcMiwNEutSaX1ilMpiROoy0DOIpE3El22lbGREMUO/T6c7qejbmo
PVivHI0FrzCeb2E511v+pshmUhS9jBl49D7nijASPj4QxO5uhoeabAf8TYXUtRK7
D47tmjzwJgl4boM5K/Cx1pT/VrbObCouxMKfUp8i1/tGz/dm/OTMTvbDj0uXkQSA
mwJQ0weS7Y6XPQUfwlU/4ATN89Y5R0fkS1d7i75NerG4zRTqIsdz2NmNNXDlNZT/
z1oPL93jtoGj3UkagRTIslJa0yVKvI8kxThHD+OG+WJyLEOsaLwxpjULmP1swWll
EoIyUrzXr1bRuq7+s/FS9UnvGH6fE79Uc4oTD0L1k16PTKqdh61AovFwd8lGz59A
+JQtqRYxPWyM7Za2gC5HWyA+vepjj0oUng6tCuILWfki1t62aGrHuwL5YOHXmenD
H87LlGb4NzbQHpR6Fb28aqbocphEn2PuhbvIymxwxyAjC0YDqOa/AavqZx54Smri
3VQjNocK+nx9Lk2Ob5PpcUAom+5l84pTx8VghUQ6GvbAQgUTKvvdmFFtBf/hYZBV
h636qTsDslSP2U/5y8S+gWhzWan6BMeBUwJY+uQM5fpENbwddgw1KzZYRWzXYtB7
BE5hG1U1VZtGnAVEITjUXRttNh7stOwLy1Z+8r1M1ZMoM4cSc37ZcED1MJ31Of8r
k3iaKbCt0Lg/8daCODgcY/siY1/+VCy9pbSBcDBqyGhUxRY3W8vrGE2RX09Vv3Bo
6LthmcXNkpsmjmavK788r/Yk25Cx+YJQ1Fq/XBXDumGKTbvmcnftCfGWtyqz60DI
ELAvvicVcS6rCIuRAzDLV09r9hOxFlfmTEGvaFMIkyc0FszOqNi3FCGFCKT0mmHb
yWHnRnPH+2PTkE/5kx4KBsV7SYC+bimZmORMWLfBT6DLgNexZT6gILbpg6Jl6n7c
Ivk7X6k73IuVbBDfZXOvOvh+Vw+fBqDgNKN7ITVGTc/MkpO7iv/lcnrpd33Lj270
51+pFYvrgxNg1GDiAvoklXUi1R9CnGSmjYSwMuVJp1XwQBoFsI3e+CJV7hvMdJal
zr/1fmo5gf+VdU+RTY2l4LzQJ0Jx2ZflcqR2NkbNAn0H5djNC8KpGHeYa6jqxnWb
uC96n91rKJ0D7Us0bPMswjiilud9r6dzcqbVEvsjT0g5Eo+Fj1WeTFgNZUBwS71x
WQlKUl9jWn02M0hPYChrVqBQKYxGVqgh0xDdrZog55m455QsxYp87lpL8u5dL6+a
SjUmnT5YOsIddwtGVeogMzCiwGjY6RhuQBwLBzl9yDMuWSUL47igJoiPoG0B6lhO
zrtGJVns8qDkTVbljR6cYqzArZDbXcGMi8E3Eo06LBNw/smzMcymT6GNpYDLfN4k
jJOoWyXBXcArF6NxytBvTfZeIjm5/q9OcZ9Em5RBZPHugX44+wWXPEjy2APxRRkK
n8Q8ZMUdkIw4MVGt3JcDXRmMsNMo9VlN2Ae4T3KGpENHouavcrGx3Eul9MC8v+NX
yGr5M5f2tpq6XPcKK8lk/vpxbVqkL5HjjSUTJb+sgimoK7kCs5ZBHctP7m/wNks8
0y3N9GgtYL2ibx63yYXfWi9lfmgufUohlOqS/0niMPyT+cO5Jfju3ctjR+g7gdXd
3akEh/rayL9wlqzl8rtqZC3cywQI/sVp9Y2A6WD4Nm8IAWnDglL4I4hnQHoPncoA
ZaLhGZN334Cr6aCqyG6iJLNTtgHEvN0CUiokZZSL6YfsGVjxc1wQ3kqutPN+7TOb
uewexFpIENQjh/p5ItUawob99LJCOqHV0Q4drYjUyqY60uCxHBF5/e2awmeleFMf
Y91kvWQoD5Vzbnhf6gCqryx6ahVziijv1NshJ8pYa+3sMTawMgdaqjm6cwCAOroR
jeh9rDBxThV7rEZkl4vHMncVmxGUDu7+JqgIAS2O6AxEeSZ+G3IsV5mHljSKoIlh
hD9eN7ZSdewTSuKNF6Akju5/6IaXc1485CREjNfHF/0bYz9IZ3S3y1iAW8hnGzPF
GXWooXx1chGXX5AWdutOo8kwr6FGN6rG5eKocQBsrhf4RvImYQXu4/s8tfbUeEaW
EiD5vmwvi3e0YsRP0tzS2lLBnM411MZGVgSSu8ty+j+H41kTanexpdzbBJpiesaY
YbVLDhLYOj3Cp8eMwvC9PIVe59Yhf43e3NhMW6m/+MdH+qRh9H9aV9wjwBU0urox
WF07G84PaNW00BFohxhwqyo1KxlBPPIgKV3dqUonUPWqwB/Rw83Y7z9WchT/9Cpn
lrA3XkEihGW4WgGvfSatVNwqGD+JniUJIMjibyYbYXCbLHsqmRywmulskojwk9/0
zFO/EJ8ON0xVgHCMcpMGqgZuyBwF1dOSzGrgXzQRMA9PCnETdQ8WV1OAUN57NrvX
TB2pcG2pkPe9RT3R/kujcJznhHUAtHP9Nm8e3RsckfXP0MRqVFRMhWjTOUVAMxG+
`protect END_PROTECTED
