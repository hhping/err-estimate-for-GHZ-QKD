`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgQskkqAKTINnSjQKN16R2fQsiEVJkIeaZGDWEVCT29arUcB3jZ1Tp3vCxo9q2BI
Ulg8FFTe0yr08bmwXddZdxIKm1ERziGBvflgepusOuUexYqAoKSaRscKOUu0tLg5
cqGHRiCg/nE6Foneoay1X63dOyMFdnt+fjdOvvqNAUNkjVOgT4U5qDRTqV2gXMVx
qI5BBGV5ZrrrtICc1/K7mVVL3+T9xDugfy/XoLd4h7L1dGZ7p8XC59NjOyc8SasC
nEqXfVA1V55OpZSp7BiofxsXtE2FU2k6AdCUmIuRFWRORzTZr7lgFH+w76BPNv0u
JAxMFCDOBBmw53sMYdvn2/HoMfpDpcs7QVVfSKLER7YOtKbXqit1wqqGadWR34fY
98qZLtAa+TIJJlGpDYmLjOBSBq5PRfBrasEBwERnUfZKXSg48Ed8Op6oqrYhWn3W
ntA5Z3k4IlvKZZKAF1gytHFJCKOA+eddMNYyuBYSDinqPP2T6lpDBMd+ebxIvHK/
s5CLgn+8MWE2gSdMtlovHjo/uwKw11vuHijZ1/b1eHieAOZZvU5KabSZljr8wIma
DaGnK+DGX5XHb2LSQmCDDEkHiWCBxEbesc3RrX/K5h/NMuOIhTSFH74mss+UY7rE
dSsqAbmGjflsfnpK7cQTDSvC9jhDNtxVhrJVwMQfFOA=
`protect END_PROTECTED
