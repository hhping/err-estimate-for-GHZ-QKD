`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2I6FlX/DM6QL1DQqiByEsAWyafuf1vvO8d6REllsIqQTZkeGP4tya3B18K7luXZ
zEE7u5eQ4++abox8n6bs+AL77ni8xDYX/fbZzB92wuheSA5ILtAdK7iJP/T8PRpn
fSwjWl9q8mVYPIz+uApNnZaqtQmWOw1LQuJss6hsPdQdI8bq/UYJAwZNW1wVFqvq
QuFOWcnpdxRzEazxgxyg5+0eiqt8EP7Hj83tU0Wy8HFCwBQcfl642YqhvDOcjzs/
RNfX7CayIJOKC+kjM5RJdsrCK5MpyiGvP5Hlr5b+5/O9sSLMLJsxUSwCud96oF9A
R3Tw3qBVlGcaZ8vuuaPlNvop09OeFSYEiPNZyYNxCpjmwm6qlBl7sSHtDFD0Tj5l
kDUgfHrYMcFRSDSbkT7//sWbIW5Ir4mzhnO4QiGAeUbxfTSWb+vkufBO2mi9531B
kuUZiiDvU1aNCaVbOEN9C5i5PZrq0eVS+iuDuJBOhr3B96ppNxyrF5KDsInDYzeh
YUDm/zTIzMt/znxMZmiABZbkvCYXwrwQgcR0yk5KmJSas3oFBmYf+RPuujpmk7+8
q8Uw0Pqb6Bvg5AaD9JtfOzaK0T6uYbIKSgptrRIvcTFAOG1/VrWzdGydvkQqqE9t
YFedkqVWy7l2q+b0igpE2AAGwdFS9cww2yCNAS89EmRyilOJcqe16YQkY8zlWbqe
zV3R2HO1gAzVnVeAvyX9KQ+eDLxPyTjDZkZnIA1TPUJCt7UEkgWLd/pGbaVo6D9x
kQsKDqtjloc0ZN50Fc7RKI0eTLoXVKkEO6rzXveA9yGuRspsHZxUJUjSxwyZ3e+z
IAVB5anNCPbB6vv3BAZaJKxtcXzyf2KqNu0Gm+XX1ctzFLvFWk8oBsJojUbgIUMG
PL5xcq1ouzYieW44sNNVY75G6fUYcwOmK7KnkQG1ZUgvg7wx3a+/VSVNciQnDxQ9
By/Y4/kJz4XogQxFt1mxF0uF2ca92B53o6ruCy8uz/t4Fr5thLYag0xEAMUCoCzx
xMnAQKSA/4sL+MhYDj87MQkjXtIFH2as+PnVhk/CYdcs7ikv5oPYG6/6REQIBRk9
DSy1cTtVuzwMYrqnJob2TgmksFHZelc9kIrUzc7O955+hOSe0Xgg5IyUt5a6495v
43STMkaNXIJfP/M6Cc0zNvsRfcxczFVM7Iuk9zXfDC/wXyk5G/4tBdCfrYwT1X08
/32LczhO56HtqAPf3GVL79bm/BNPsYv3TMx0voKVaMqN/kYG3K20iGSYx4Begu/d
gyTahgtiTzgpJVM7jc/3NQK+px1RLMAubB/OHbfROWy9jvMRJv8R6ZTuXoG8aqaI
5Wwh4T/mOIPl8Eo3jxLzE7bzlBeeSF6nFczqsxwYopN8FACWtVddfuuhHJfFyEMo
2UMmSreROnEcohVgiuwYA86ytTcsluAm3/6Fy2QxvvYzVyEcPhS6shViat8AZaZB
HJRC61jIT4kgEa3G3HI8w2ftO2hQHxrMeAT40XdM00W/aMc8C93s6prpzRTR9pz6
+bizqKMFX0eAI13NiA0lm81JplTIyhQOS/ZvOSbWSnJwao+zXvHxZ0Uz24a0ihJL
/hdy8IVWnKqzXi3MFS8ZGB7k9h2Z7sRHsl2nh0OEoxAWZr/X2vbkcRz77Vu3FUI6
WUqlHAtr30rghKDL93curS08gQp1R21GkKIBd8KS1A2+lJImPMQEs7bNAaOTuHyn
0ZG/fTN7OS46OYOqdz2YFBVplNuO9FMw8uISbwP4e92dPfa+bQyARYUjiJGpziQk
xe8qQCqUDPSmNXXXzvUBi3lKsZfsY+v3Mx1PAaO5JNMXDNl6/6Jv8LbwvtEex8dN
a0j1WsHB1Mt8IBuY093io8VOUXI1kbngiZaWbzDrNH8i+6SrdWnRkk6uFD3UDNdy
JMHdiiTvfB51rVpLkJw7PgcXcAfiABzMcA7kNKlrAQnFHl/ZII9isqAlryOxtUQZ
+kWVgXqFriCIl86+XE8ZaCMiyYW9RMUrRkqQr/xjugslTz6/VfqrpEonq3OodMXx
iyWE3CVykUn74rZOe4co5u3mpYiDRaQq6Xacjyk6aMf0BansEe2KuuurLCle3MRY
zUHhgzPkbTlWNg/yi6vjFSYyOZf4p/3ZhHrRSzc6ymfuKn4DvlD8DuTfehNtlHUT
m9wiA8cedyMg3dC+HJcVEKaNDDSIj/ivPDf9uYtFuFxYOgfIxdEFXUJp4JM3sn20
t5AY2esWKSm0hq4s2rJSUstsSSMm/7n/FRemkqUOlG+uBN14j+atzMekoyoMOmxK
5BwJag+ShzEMfoJ7VTLFv5ODoz/sG22vwuQVCD5qZqb+9hXIrYK1Rv6WOr8guDrc
dbnRkelqmsQY2nNZI0yvM9MsBk2NQqMX329fxHglLmdOh6465HtZ4Pml+EgsLaos
kZMOAarFQDP9z3EzfkJQ4GWTah9KejGZs5o2ZQhfE5MgVs7B9sbJWfnslEtWhS7v
00EHe8XdKzl+MVH3HwKLsBIZgbSp/0jfDyW69NYxUEJiy26xBLrBj8yyMt3eObi0
l1V7WJJj5cSCurUZHoX4tHvlfiB5sjOIk9f8xBGqN708Z45N4YDW1WO0lY2hL7Hm
IPDk/iNAD0iga405QuTiIY7wnC5nzQuCD0SHJ1A8wQNyGQjMkHCOsE27kva0ax3j
RRAWOOC95g7ZCuNgXnEgZDS8lYIqRzGXIHBWhKcxEDlM8Amv0eTnZBgls/q4SHVt
7yr29YCsvQYxG/qs+RGrEE6M/i9UlcriTe36YJy7EkUr8mAaCgupEKOww9qThnY0
YW2BZcK9FaWtTSgKWr8nIZLGbIUqut/zz+WOBjeWDE6RtrGDOwdV3X27ehW08bmM
+yjcdOW5nKTtdgaFa0DlOJGHSF/6PFOv/IfnWGhu5lfJkHhSmc+icdHxiFikP/UB
G92cbMA7cb+xrAkKJPXW+6o5KY/aoyduy2M2ECAn3gnqdWAOd/MhVEfga4k8QF87
i8ZGw7cUctmTOCnUGbjevBaMfNH8E/ZTI+NM3kEni7lj+IP5I/u/wHot/+J092Lb
DKSqtXm7IvYYez5kD+h/BQAky00/SHmC8VS0qNcdIkWHsdOW4KidSluwmVyh/PbC
qVSzefQqzxpVA0Vynb72iijKpKJCKNviWwx3cEj8MYH2wQ2d6kUQDiMAZ2NWe4KB
Vmz6nLo36+UvujLAM/RVVPZQO/SwlQ4s5ae0kgVi/M07ZovmXQrPNgdJHtDGEsnH
XI7GGPuP6ouDSWglqlwTPauUHgMrTpTBDpIk+Uze9dQRwbxlIPrzHrFRWOXO6aT+
M1/A8f4+GwPW4kY9KaDU+b42eVFgJZHF0lBCwLz5HJa84n+lVwLP1Bavk+KO46OQ
om8x73KD83AaWl9Y2gzouxAxtcaps1XadQQ64EEakjG2oyThu5dHUrj6qFwZcyU3
MFaJtavlyKfh+bDdqtfaQLudzMKc7Xq0dwizvPqkgInL9/We5aXXr+bJ5g+3OO/O
36W/uUCIoru2YAE47d3Rny18pDsmUAkBzTPSJBGNHTaTxvcNaBNNJNaQREfRNvqk
x0n8pbEUgd6mvmF27Etheqi42q62YaJ3UiT9T+G9nxXek75+SXQaYIPkPWmgYKhy
Xd6/ZKMrVU+KhRuWw5xi0P5CETv8eS2oE/yl5GdlTYXcyWPe9SsmetBgvtI+SyEG
V/BY03mc3lU2E81XPBsI+b5bj74hrur90+FNqNMDNjCOCSzVXHQ4E+6wANPO1ZGU
+rPhQydyI6Jb99oIDe+G2MGHXv8YRxVXB3MwyEjSB+g2j1JCcYNs1VKPI9IN7OD/
SDn1ZzofgMTBP+vuDpLphzwzAfkKQsJSi5KjYQ7FTh0YHV1aWyUt51u/bs0lEaMs
SYsfGEfwuTXPFqaXaPzC7UMgx4PBblSqQNcwFBKbwBIhO7ADxpnrY1f5cOX9xeV6
bpxrUJkeB3R/CzBEC/+CJAedhDXISmW/BXqcNNLqwILm1CeI0dk17LOalgDOZvP1
KaC5lQK9UZcNYDW9Fm6Dhp0cMHoDZT0j9kJvUtZlF68RLEgGDDFkYb6RWE4ldMDn
Z2fxFtNModc1N4kruIanNHZ8/duL2u0KDy5LL3sftbaPY/ukzMJE+hexKyNDgHQV
LEYdMmNH68pL5BQJ9t/d+1RjHyHVTz9YhC+qn5GHXUA7UGpoR/i+lHqWKuFj6xFM
epwrce2+0lfKgELxi36W0lujvoIM3bjt7mMTRAy5PitVG5lF+It1qkHxseTvU6FG
0t9HH79o/KgA6ZPfFVShncvRu0ETAALSUgmrthubWr2d+xqlRHRxiwc9mUQXdhuq
Ui/S9nhfgPNydibVVD/8Ck+zV2cBuYxwP7IJLpvd2T7pPMijpBSgdUfukE9n+L0n
Xmm+qXnmHBUjAQvXz3DSQIC5U4xpWHh2zN/sK/yS+Vsj0OXx1Hs0gU2famDWwYcC
m7uQZvXg4E/v3eoCNpuWaD7bMxM0UoICjpzPYV7ZMftkNPzjmjkrR8cBfi0n4AZ3
o5f3A95KKZ9xzifThXTbNCvQkQaCIXt9hyNoaboyxkCGdMP8Y381dSaNw3iyMv+w
1Ye+j5NIAVHP9nqaMd4j4qyE7R6QMJzDN0bgDBfdOpumBkMWsRpwW8HOCwMP3qTY
0IcdQOzhw97e3giNVgkhRHLslrYH8yTZQA44xgfr7LynFI0xbveDDwn3+NtoHSFa
2nlKcJPitggVONijvFn1sfVbODWoRp6/WwSSYocQpVSKB6z1eGkFRU6v6Tlmj0hp
ve5cksnygtlKqPWa86MWEw==
`protect END_PROTECTED
