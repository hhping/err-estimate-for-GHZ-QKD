`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4o7MSw0k+5/cfkqbrYahGUMAHfftu98GHAdUFQLL327fEfY1mQuE0SiJrldduCd1
DKzFOEv88sqQ7qB2YrzP6LL28hBxcfabPI5QglgNgb0jT/qIi2Q/dEbKyB5qEPhi
d4g62/yexUdfNVh+wPnR9Wub/s2o8UoDh3wMV7cWviZqkPH4WsatVm3QsO9mfz4Z
aP/rNGNdLyzbLT8AwmfOA7u/Vqc+QErdoV5lED9m9ElvvwOlEteUSiSmEK5FSU8C
SItfMdh33qBxq25NMY7tX+AZILfiiZvnwwqSbuS1lcCMa2aj13kr0Rf/HsXfNsHw
kU/FKdM75E7jt0rPBMpy5lgB3sbBzad3bSB2phztX62rEIHyZvSV+geKWOJ+Ww+W
DizmiNXt8xxX3PPv+0i+5OO6fDUasnj4P3hoTgK2W6pGZlJjujoNBY+vOmwrIW7C
jA6LRRMGRX3wkUlwEiMhfnY3gNoj9o0gSJrPI090Umg1TLDDYytTkOq7KxYfX0Ar
gXYMHOillJN+X2BdtZpIybIu9iTHH8ZAnvIPtjPesIQ+14ElsgXVM3LCSqi8WU0s
P8TvvU8T0LiVQr41WWL7wmKaFrvvm82NW5izvlyOqmGwflH5X5dbhIH2vEjpJZWM
/rQ4Y+tZOHY+ikNu1tzAYhcXjrsl8xIgKnRvGoI1ZybtQVUqmAp0P+M234tHrBsY
lIlFn52MwR6EkCwiLOgjWIE8DyFDTp6HnxzW5gqtpgfzqYgMHILlRubwcHbFTuLb
CuBvUsEc+ZGMBNavpHOqafIud6DiBJ6iwhqn24S+BGCi791hP77wnc+9JHKvkgNP
Vscc2IuiHxfkacw5WvF3Vt6N2ZCFjELUBd/V37550cCu3t4AOJHqsUKli1XsUTNQ
kRwLa+cfUkrq7mNtejkE610TAErBY/zp5nceRFtM4cdC1Sci8DqTaVpXVQjGKEda
zNvowYrp1H8xb4pr7CPoV9bseH8kFhtbGDXu9k+j7SeB5AfAmxRbvGwLKt744O6J
1GkmGEBMo3epvYRqDMC6jfMXXsEcyORWBWfZrPeHtrN7lWMKwPZoSBQJRr4JmAgu
Cq1yUfv54DvU7l0DGMfdnY7tMWKxp3Ne7mxFa135z7VSDk9y0U9GWWlau9DTr1Uj
`protect END_PROTECTED
