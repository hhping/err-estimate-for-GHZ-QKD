`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kUyG4cCXVkFWiFsWbem2OFg2hMe3UXB6mdt96FH+7lHS7u72JwIjRCJlWDKT6dG6
wNGiiJyylW4gpsrs8CCUGDaiQTVa6VbCG2EcGuA7yKcrfp7opEMZRPC63SOLPvIB
N8DcbM4mgb5a8A8iGTz3EsjgSWaLNGUjn7UhnQTRfgM9VchygqlV+pWT8ZGk8w+3
g7FElXiBoIbY5bKEHHA+4KL/esHX4hRATm706OksxUT2Ffk0T8av78vjaIC5mKI4
SMaW7SCYdGOEZE9pOWxPAeB+24/nMvBzpPifqHcR2MViJ8G7pirjoDty3BddEuPS
iZdulYpbZC3G5iY5inDau70iXG56Ot7UIbHuGYrtHq8odwRGwNBQwYTe7lkS8EGG
Sun90MJoy81zEn59prkq90ZL4jNLXLxQVTRfzpw9Y/tEJPME1XsXhhFmOMzLLVd5
wAwA6VPu3MnnT+Y3k0KUyJe6P1OxB7iba8PVGg+wFnPOdfn6j+S9fB+egXLC2gV6
xGNiLW5KOdbilhBJ89XDqFzWzZRDrJZBW3/ISmRbHmKS6jlkMcV+0rCQu+adJkMi
uimykgcfwxH6d2lLZeZ5FMyw2SUbZlTB/Q+RrlhkQUksv7ydaOO8mojhCs+4rFLA
BTsL8+4iDSi4MMWISjCCL4QsT3RfvzzXcmvGlhh+GLYuczjSzmTHU9Kp9i40HCqx
jZsLMjuYQQ1KQeTRrTYB7UuzUBjruJTh7/ULFsTvtuArr9y86+z/e6wqBSRcNM1b
i2zrnrr8SqFOtVTzItwn9J6YAS7yk643nQ8qu2XZYiVFcn3SQY+NQWldkqT9cWQb
X0TobgAOp+IS6mBkfbdtHDGBG32tFlxd7vktcJ0KtNQyKcUmeYMgNMRnSwOD7bQd
7jJyUdiP0w1TDMcXs84ZI3Vf9Ci9gMu37bCzo19VkVw=
`protect END_PROTECTED
