`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7VaORvEJYbZJH0Qox0ZqRLagQFwqN19Z/UgGUiO0E8M3fdcmzDUsFl5gOKf3cwb
UNyiIrS8jBob2Ws0sOhp164jA04LGcduIyLzI/PtNODALNHKOSyEk9WiUjR2jGRr
aSWnt14gx1G39RFV5lp3Y60gFAWsWvo6TxCK9CIB1thMvKULlorKnooDB2096s6I
9oUs5TdfLhuIIzu8VPeRr0N23nZnMyhHmRm5r87zP73P+dhukfSimTWGqg/BVRDf
+qzGDv0R/+MENUZqZVZgOYUa9T/5EPoL0yXa9OD/tFdcQZnKdbR7TImVaQBltNB8
MtppV8LmwjQaLmTXuAdNUWyb/Hs1px58HAKE8yf9m0cHxefBvmi8qe3emQZK7GWE
0cTRq//TYCrbr6t5sfH/Xmk5yNoH+oLmvKnuxflxb1Q0KShlY8DhTzEKqxg7GjS/
EFIjO7kmTVV64cifJ8mXgmMn/lJqMmq4Az4qU+dYVN/vkdyWsG9E68mncL47lM7k
Jcp4+gsW1gSjbHxntQOgMeXsAQP6oWcQezblrJLN3aNJm+rDvsKrL6ttFhZrFSdX
OSp2D+8YhLq/dpT2lTsUVtwY7lnRoPXXkCa4H8+1KTzczhfBeyzEolnhbzdmWXKT
K003U4c76q3vUc2q3RRmgnDalL/hDDCY81EsKSaIbAroi/Jxh8fMRF0j/IRfyRos
rDV0BGlx7RDplJd967lPTw2grs7uwb3k4rViZOV5kfjT5DncRXRlcAsJhtLhp1VE
hc/JM0y/5pKC8VqejM05b3XPmpbcWcY+SkAEGU9tI/bDSrbUFj0n1K0+Z12F4JXY
849hjzvNXS84KJMl/osi5rGWStWE1tTxtg3Ht4knMIOJp7jxs30t1co+hDGBr4XF
61fpZK66z1LU/lehtSDq0fPx7KWC1SfKRybTbXlbsg2VgC9oY1O3934CXGLv04Zm
y0U2ASOJqpIIQSy1LaJRuhSq4u4oc1P+ccGIfo+yqQLwFA00Xs9vFM8qqg1w3oKN
m+a5fyYcmxkevG6+pz6vYp5+MnCFzQ9359I6NG2+R/pUkiONbW7lx806G/skptJW
5cIlzXPx/Yc+46LiZAsIeUSiAMFWbKLsNRMqt3bI6iYEeQ0xi043Q7Iv0v4RdUv9
0ZR8qGM0CviKXOhFZp5h8ufZ5UdxoLEcwBwwIuSDUeO/SFhLqC3AFtDCHhDQ+S2m
IdQEL43LeIFbqNNp2PpOWg5Eh71zUpstjcT4nbk2zK5Qe7yt5P9TRzu4SeDIlO7/
BZXKdgLbKyGhUemBt+HahwDPs+3skO3dSW5onJ9NYshbq3/szQKhBlQ65ZpOumsp
VQkA2zT0n5vEi/CRrNKBSWyBZywdy9ZDAl/qMOWKWQP4qZy7vfeiJ4usSP+Ac/s+
UFIyDPBc9laH+xpwCjToQuZlY5UQ6ji6/NmZrLwpZnTNrNdBaBn/wa7JppSOalRn
MFFjqjTMfBF9UE1uqF/irbpu9VJkaq3jtDnaeEAXrEpHqhoj6RMXYT1LqBFBKxav
9XGxh8fwLx5zTkBR0jkn7cAU3D6YHkuNelOj/G6aTr+h6CnI0GnKeKv0SRJDMm9E
VqxWQcHMqgkBIUqWcTdd7cGS0THDRddJ7eGtNTfE5/DBMcIh0vXY/IbZSvqIeAAC
aEcydGVdIasz72qHT7zwXLnfIeiFuE0JX0khH5f6qfh3va9PtevULbYszvCpPuET
lMaBhlOR9En2081S9te3N+pn+dNykc0NFXALqIVeZpsEAgws0//KkPZZzyqn7S6y
Ej3nLIOna6jfXeGBpOGM/P5D1g58iDxj0trgMgHW6lY+Ven2AD5Kw9KdGM3eANXW
FVqEqMsK1LyBrnd4/gge49Do807y7SIRtVLVmBwLMyzqv0/EsPHHRa8uUQbF2o3e
dXoymgtan3FaUWarOLZpG0bP+PBoLAD6p53swCg5uvgLX7CBnd9GMhIqI1s4/IWC
ywQO6HqKFXpN2306svzjcjX1Ku4W31VXLGnkfC+lUd3ekAIpBwGA3wafsMMxUzOH
IdpckS1DFIf1/xaoAKDMswt6rFoKnOuPG4x9FK0VUFU=
`protect END_PROTECTED
