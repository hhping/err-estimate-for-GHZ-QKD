`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFVAUk96UVH7wTCCpUlXFOs9N+xeANkgtLt5ido0ApRI44CC9z7te/Kjr2JKIGJ6
p/OAktH/pJIS5sFnTdukTV08SkRhN7zUtLmVXv3MSYn40JvposH3GNwNs25/ppFS
XeGmjdyJ2QNtqT7m4KcBOvnFidg9Vu9FGbXQT1fdja2FJxAbbygldeeUxLXxPP/s
CSF8tt+xjKoHpsqyJolF7EAtZc+cOXsupeNvC9wcTLzF91wumVLXBMSOmKlSNiLU
8QikDC5pJd/9xN4Wi6/TpbGhNNmdfvfZ3mgMyuRqNB0awOxHs1avr5iT5aGBlRBk
pqvdp4owf4HmO/JJQbaoCZA7GpzomMJbs3ioorJlubwPBrrttLDzN0q4QKntftC3
iyslTDs7NN5xQCn+mMxOSh+7rjJrMWgup2Dp4r1VNjbsGwAXO9ccIkeqshi2ulGY
SujAX0/g58D8DSbsZxBD6h5/8tpTAI5pR9l/lxzRinrBaG+lBY5EF9FRyvsKzsnr
TyhIpqnMq98ZoAOg7AswKRtp9qKLEDpB4st3XAOcdzKSBJfDn5xs9q7fzgfaCjd2
`protect END_PROTECTED
