`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ardtxA0TlUrJ5QtDcVkCJTAyfvLnzk890ekjx1d9euWjynRGEHY3mmI8dHiYT8KJ
8742+LrKcocOWz68YdqdVWv6KNmP92+/G7+n0hcVtYV4nFmvbvl0gSq6PgMwN4UM
QqHNi39Qp3/C8Y36ZWgp3UJnGiS8X305Br/BzNeLVFCv53GYMTlAKEMbCiHu93Lj
tnW4um3WWHiaxnmZNIgkF8vbz5rGWW0oNZbn4X75wpy9wzzli71r+0ZybMPoTxdg
kLrkwlB9/z9+DBU5v6YrXl20+2J4BEy36V72LhU807Jzd2tOGNkk95pdbTRTID5G
53hjmqiZFOt6soLrtOvQhb6Ph5t0vnsJk74/H8NaZXJwUQcTzd3Jm/Gexf5QMYfx
cvxOs5scZJRzCwfA9F+NjSQEsp6qpn9bYjb+D8DXi2WmeE3VoAQ21HpUoUKnqwEI
ay7yw7LK8Pu20SJ8Ouotq7DwBz6QMJBAQdgAnJ0pIeysNUkKhW9y4nDGfa8gj056
XZvM6z5UbatLBSg4cvNGupd6NI61HHVUwp/ukljCzvFQjjUMQb56vZihSPAk6alY
11M1JoKkgr2WXTCsz/OCyv8w4eKgqiMCFp4kztZET2uJHUquhBZ/B1hu7t6GupIj
UwTReC/rB5iuVhVYCXFvtklGb8S5VcxTBh3f+e8dfwGUC+qbbqnOf9fQcdw14s65
pscoiCnJRE0el83/4mjVIREwz9079YWfBcCPyI2LUAk9T2XEsl/d3igoVbtaGU9z
3rW/mjmhUa8UMfqmGQTg8//ZtMP2h//UPBTR6SPBy3QnDJw5PgweePwboo5lfI4v
FIDkODZlt6wXIyR+UdSNIWIwIBwchkDBSEhRmujVgRpRRbufkg8/nOdKtFqjipi/
YaflKkiJpwCHcBAftP3tdOqHQc6fl3Cb+WpSPUlpm9rPUwrJpuNRStnsuEHFX8Jl
wPzFxrKMlVM8Li1SRONXQJ95BRLzTvn45YlmAV3EtD4GfZgwcXfdMc4GNowfDA6I
hbqG8X6dsCATDE7X5ahZRhOd5udxBtduAL7Tzd0dwxzLAlTsHcSigK1lEXv+Lp7H
gOn/I33K4m4cKNep++7TxKamYrzCRUBsbTy2deMAchfQaf9Zuw/g6pUdFGl5CBeu
rN3EtZeOnhbum/yGA9/c7sNBqFeinE3ndrfna805PiEYF2bYFUYb4jWlEFMGo5dl
8x3wRpLcscK7qlHCCg6+fpM8y4VT/bVL/il63BUVawSdD3xVKut23Ig05FZOeVPW
K1EaXMI06ozgmF+IXoQmtI1ht1Gx2Lt76kTSFu9P4tDwYJadI6PJkR0hd6/I9XEE
Rv758ENoZqiKpg5ndq7hcnm3a1jt948tE2Xbb0bTST/p5GYMpO2aLw+SgUBCjo2r
BhdFJe/wT5TSwcN4GoLmJwMUbY2gx1gmWavRMBedoei5c6tocWEt4XKpE802aZef
mn0uIxhwZkRid8Pf1ozplaoIu8FvYirRb45sg4HuKqpyPUIjvYmQlCXdbkWiwwLW
7YFMSTpeAYUghJkoFUf4G0WnW2KizLxGIjvlrJgJBjL9rePp4Vei8kcQAXyCxfOt
dhhNaKf3f0Od5RoSMQzPPh54N5V3w/5WbqspyzRiv6kPpqDFvW7CImrzDi3QeCOt
i9UmD/WL8NQbD9NIKzYlEVkqJ9bY9O0lBZPnQOaZ67atHOB9EvcZRiIIidjmOq3t
cEclRWL3N3NP4pzMEvMVwzIcJk5P+nDurIFdIIM6q+HkF00+Rk4asfztEl+lXaMQ
OLjJTAfeil64gHK8vuXAr72ggv81YhfuHe8L9UTjh8GfxpX7mWzPVPoALaaF6uZf
qGV8FLi/hpxLJBSByvfVpFUkLCh7JWcgL21M+R2nMM0EHgNvlmSoMiSJbJHbFHkw
+FHgCDLiptlgn+yWikpazL3uGQ39i7go9hsuSPwPsCr3UbiWj/TXsvB8VtvE/FBH
kn8kjxdpJm3uBbPrKD6lA3Ar8KvljTvFQ1AefFBodNVq97ese2x6SA9RysfxyglT
BZYxtPN2OndSlPgTnhZjKs7UesEfmg9Pu1pW+xEK4fR/d1zxbtvq2FOwgs4giniw
iuV7jOOzZ/JCzw9iSabrxJXKpn//r1QaRIQmrE5Yq7Jipx/1nHiZodEKPaxPjKLo
O8OdPnbJGs6zitA/I7auM9RX1FBqbrWB54su8w/CUDdsvRDRFyWML8HBzN1xgOeV
WFvWx175aVlGLmQ4vmQFxLhkflkTSpIchDQXjTqUM76iQZt+HuP47X1HeZCNKEA9
oi/TRuMEu+WUBTaTS2BH+Q==
`protect END_PROTECTED
