`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ttn5jLWpAocFunJZnPKahuxNmamsaC7QK89fVCcAHhM9Kn4pszvI3iu/kWTERFJc
Wkxxac4prgAWT0a2Qg0JxbLKCfYsKzEBVq7fUnmnowAGl94ML+lL/B1RRSr44+1C
ytp9XeTgSeU/zB1hZo3S8qMin4ber5zkIYf3cYwxIDkEKx+Ibqf1ACGSIrlhFLF6
a7NOk/gjIROF4bYkdS1L10NVtgXgPtmdp6jCmmE8rP9HKcBpJLWtvql/i/YZaxMh
nPsV38SkRlwAmMVzlHsRpFBTZwnjj0cVQ53bthcpG9xzu4qezAnl8vxw3o3eSTXS
FxvGAmOrh/tm//2bb39Ok+iRBHYGUydKWTJRllp9f7lELCHy1aUMrywUpFmya/Ab
J/H1cqcq/K7ZqVQxVevJiDPjBvcVWkmuROCjGyWuxa4=
`protect END_PROTECTED
