`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pi1HKmAZ3XB6JkudANTVb5sQKYxpWpO2nsJo0knJJwHRjZaw+SZBgZLCLpDx/g2y
9Nh9MKF8iHHWdhQFOQ57safbg8tiSPdM1s9HYaR/9toRTvRI25gNRUGTi91YbfQP
uqKjqlXtTMKU9FGBL6EuP7rGzGNunMPuGsdpQ4btdlm+7mu4PpOzdMgojxCXg3i8
VOv5HRkeEGqzSH2LMJNa6j2Vs+rvjzecE741cGsskX1cA+xiPTLg29u/AHD+uGSe
D9353tvAA/GvG3pIJiwDrcJz+3Cm494lxk+EY9SpDHRyGJ+0wQvYrOWKJTxiEpBM
D9fq1zkDIqc/a3oeUkAcKqFB9hS10qUlpPNQmemh2ctf2hwXYvYa4xFCAlpiSgNL
1lJ/skPdLPc/82y2mmQ4pwuT0apq2tnkrAzDqOCNIE57jGK2uEuC+VvOkoLtl5+k
O9swvzmDlqhmVTJgDJ0/gaxKlxNT2UwFiZduUsS+GlcQFsnO6aJ8mXGiW6CsOGeb
q0ESxW0tsqYkNKRObVR68tHkuiR7k0yFnEL4clSde73eJKH3Qt4TJinMJUCPtLSQ
Ew5bcfZlHLAqcUZ+rx9ngn7PQT4IgHnIjgiyyTuE1YI+5C006RE9COGUnDyKxRkI
zm156aSY2uz0qCVBu1fgufvTWCWOEnzAMh8noPfezEmdLDCZYq8wfG3pj4liOg5f
/nZcXL20H4Bx2zzubJxtG4Kbptl2gYzRRnmIii9rTpnz9T+2iiyymTx86Tz037Ro
ndwXMBsf4qHGGPW7YxV23eT8FSf8m0taGVvp26G25TTeY7SDXddMQLpCOzXkpiws
HhAyRLCpyAFECH84yQGfafvjnZ1fZ6uQWuOCMNfjfYjXgo9yHLnl20a/qESci0Se
ok+b403YqplOjvl6ef+gdgz6VeCfwjhdbg+1k0j6SsEZkP5nB4G+sBdccWOOtW+d
ucsKDW0I/E9Ky2m7D1IhiHrxTPtiIobO/v5VEemQwMun3Fnbfx1T9c6ZMerkYK+b
BqA9IpEuS6erW25GqbqOmYrOy99jJwrGKVKv1jBjR2/OG+dLkRN2tzh96En2Yuey
Z4jcti9nRhC2f2TYwIaPjmLY0PQohQY2RpijdjZtWeDm9msXoLGT6PfAXdgQEby6
vpeTN2VhKaPT1xSUvV7jVb91Ec9LE8o777OO6rAeC2kANqN+QTrPPHnnt93GVzHI
OdCS7H+uJxaQn08qYZF7pQFpXJ0xWmTT5rf2vJqAJtJcBAWS1YbRZ2c+XuiFAQxc
w56824vQsfQF3qh4/3bFP4uS9zhmgnLJMW4QbDvST8kkcoJikJUNUxliFKPwbPwj
ExAfURqdL9K+Ai9vGGmx39Qn3qtsRW9f/XrqooB/bSua4YZuNptyoxGj0mTTzlF1
CAiG7uj43/ijNFnRbDYGHj+3cnd4luUvc84WzTZyHpmmPAbV/q6LypMo/N4JPtyJ
8obScqORlGykSzZyn0BFnjV/uL/u72SG5aL1P68NonD++KlhzaC2xS8VCaeOwlJ3
55thAmDPoFbj0tyxJz6gGpErryLUzGK1G/Y3GC/HaAdhbUojD8lzXfAJXUETfHYX
oONcpJRnEqswAZUf1cGnjz9ogXVGNzPK+2BG+ympC9hEU3h7hVa8cBnnl4lW69Wx
ZLLy3Fw33AfTbrtI4D/37tIL6IgRuKwGXRTY/+MJT3xPyVm8ZB6kuvDcZp+tW0bo
8b3DhVEcPdOYVLhwSiWZa6v7+g8M+SQPrJog/QOKP9c6Vob/KKbwlnprmqJ41s9t
QTU88Q7UBa36cpDxCKWotxc7Gt2Ry3ZJogrDbCs4obFe0PybVL1axtBXpqBN3DT3
EbQWEZ33hHkDHuKtnGpSijriHpFegIyZNfL4/I+Wdorc0Z22tZTH0ZB18PFGkdvI
IGvRN4QAmIKAeGkuoWsx5b0/16y0sADzLyLibxuZHiD7zbgob6IgvcusEEhOsXbD
1btJ8Q3SERoytcx+VdlWKcvKKnf9Atq7MuUBvlaDVicrBDoSpzHbgwzbR+5Honqw
E7PTXHGCIDVtCIPzufDtRgeIxJkcC+9IbU8srIjtYl+umF/N0bqF+CxQs03jeBuo
WdGlVFCBFRBeBrHpm+lLVN+Xu/XL/LI4eVFaYxzByxE3da2S7qIQXQy8DM8SjEWJ
n5BCGGGWElwgCUX4Tvb1LWuzOLjZXk2jw5xEokP8I6edKpI/PSwj7Yx3HTl7ixBA
Gc33ZuMhlMxKY1OBrPbqXna13k1KzWrnV7i/dhha3CKI/W7aOM8fRhkZi99nGS38
DEphSVfAeuNHtnf9UKqNt8cbmNbPT9c+A5OeaRNVgvdFj3Wx7u20eFSrGB74mmSw
jVCyl3pgo64Ku1J5prMfZbuOyXeK3tL3b4TC02wv0/U6+eGW97ftOzkz76OxM8By
g/MGgEGNriVqAEWI1pfhk5BkVYB+2ZsPR2NkQGWJzjkDXz3Hb847SDmQvHllN8Gy
bQ5KTJJIn++sViXQYj2w6MoqTgF/mBnIBLXsRklBsfjEK7K52J4Yf7lrucbaxwIT
VYnBwP0JIHw8nHod8uGnwhLmVZ5PJAdjFQ36pnfG8V2qdByL79I3g+nzW+xJJ6XR
77AkgzkZ5uenB2NcxKFF/XjXSWtD3QHgugm1TT9qvyq1jYDFLqRpcUzyp+ozzzo8
EkSU42WyE3Kaiv8u9EvBoH6xXWBFO9wsE6mr/QVfl3HaWhzks3hJO6zdanAWqsII
jv75uLtV9g3x1RLoxdqWnRMV99bp5P9D9N8VB1wSEoeUQb5ERydRr0Pjm9g1D5qt
hrMwf6En8FCKoLQKbs0gQ2aVIIBWDC/Dil1cVC4IQYwhOcBrniG1AFy9jBYdB9mV
SnExol2vHIzLof2TvT1Jkux1tJUuAtjfdbexaxr7Tx4IbWnN88TY7czzVuRujwxe
gsC6wRpjhmaWZc19XJzzsrzK+hOK/v+kfr32MQvxiTFBMri3LdfxgvoQimrpykcM
`protect END_PROTECTED
