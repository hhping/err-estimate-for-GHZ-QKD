`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZwwGS2K66GfLYHcNPi11PQu1KcqNCgrWHuXZrMVT9IvqNYfRBBVg3gtj+SvAbKO
UsP7b2Ix5A70c44ipifDdUTNIfCBZR2ZFqi8l3dX945Qsm6cNOALA9yOFFRtXAGW
qn66sDxrmaC7bG6a7rT2oejLqKqXvVxb1F/BB5OhkeuYHT18v3mZZpKJmrwsqWQ0
wPtO41tIxvzoJtsacKk8CrxQtbq2mtHVOpT/NqyjcZ5SF4f8vZccbYIqZRj0lbJO
9+Sr+OEwunGfNiv0Njbhv9WU08m4mpDMj9ABKTwBYea1Qqmty2Qxi+p6P3rE+RZv
yN2l5c8eC5DqsW8OfyFBLCmEkcf9NGnKo22Ubl6zbsOjawMoZ3u3/Ljm32Mg1XJF
fUdpxzOuEoLLHxI8bIBa8cHhp7HyVZT4sup8pLzL4warmSIz6+xKRhkImJ2CZ0rw
wRMWvpXjcCPdzfqN48RXFijvyJpE+B2MuXauH+A2gWk0vCZId5Dx2kWVfou4fVRA
qI3RDv9W5AEcsvypWldUQ1tEWeo2QBREIxhWhGxlE36JvruJo4mlZCSffRkrNmZ3
mXc/8VIoJzyHV/lkMYlCFOHwfvmZXQxSOlne2bvwRqxEA57UP3e1tetXYdvg7uSf
p/HxOVrV6smoO9dmi+HMnlSdm/f1pK5Vuy0JtTRvxcs8jIWAxsQiPf/sx6RdErTj
upxIAgfc/5bGioafTB2QUznktPpQcxHx9yjCNgNWPF3tKV9YIQMItaGf2uCHyCru
tRcNqgfVMnm/T2Z8vYBX068ysx8JpkAkXE8lpKlGnQo6wPY9U/wEkihnSiNqk1KX
+vHtKvI3Mk7jxWIpTtUlp4RTVZDz/cj5QVQd1d5UUp8vJfgnz0EMHDwyIxxpolOC
1dAifKtPKZwPKwFKdVz6NuTgCyUCZrMfyTWAWfSqJNHjiEXgRgWfZXcEPucb5n+Y
bxCgnLEKCgy/WA5kWz0K80h0g+CfUs/FwM6qJr1OtXFOw+reJH0Q2b43LTiuoCp8
qNSeYjVjx6U83MTtIVsLN2MN3lmVK5nzVXcwCuGv8XDJILZ24DaNMn6QZlCAMd0z
Cho3TNI9PsNoQc5aX/pDJCIFlI3AaCUbg0/ZxM5rJ96fUN4uwWBHsT7I7s5XjbE1
tJt2iVZWDh/D78P1j0M/4aL2N2d+tTFVUpiOBWLCwi23/gyzyYQ3j8l/Qkxt3dtk
4m91Xf+PcRwobDbPKoDccpxSfZIVTHcQyhhIoiCBBrpL3/b120cbe/hLgLul0RgN
j//ou1VliTttdXi7kqe9QJxQEjiTU6WSyCQUM3u8fcqBUNBQ9B8EkC1GP0kBYBP7
VltDPl4xA3RtTXmz9R8agyTQtkDTFWUSbPKbS/jRPZcz85BrnA4Nu98zx4/y5cJN
Dl1FOlmYlySTKUtEy7vIUgZ7vc0N18hyJcw9K9dP/Vp/nYRntlc/9Sf1GJWZsG8p
pS7wNMq+H7FGny09CkXFfyB7FLyEBEJeWLxCiCQJFXigFMad74DoKlMbJ+nDiIWU
lmMHQrobFrQ/CZy6c9Bi1BdElrF+qfgZNFOUh0wZ8myxucuwxqSywECceaYcuUH1
3qSjkQZe+Gc47M0ZYloDCq+yNBMg0tHu/LBOw/KQma3rnJRwaDUFE77ly02bW1A2
y4g1K+dPDOEk5feSFMBn5Iw/VJ0UMfmrpKaPGOpBx/atbV8t9ryIXYb6ttuVj0p4
tzIOCFztMfnmIVocXgYK8ofHmwMv1Wq5hSnULovyUDC4hsw6I18JHMNdkidi51Od
/SshJcESipGxbpK+j4IpZMSeJKMY7so8u/1/0S3noGwA+r/ZYZ8V9N7G5JiWNHnL
UNolSNN9W3L5SSh9lWNUNSLiTIvm1lZnzDEmiB1pO0dEdZ/u4i4EcVpNHixJ4FPi
mNk+CpS20IwUMeAxdq6uYYI+dwf9pVfcWFAO57uya1d8AAAs5UiGngt8ToXSI7vT
zgo26Q/cPjGGe4G1rfbDd8Y0IMZyoA0LgxJunJ+bT7n/gz3K8Tsds7XcU4LkPiTC
J4RFAFhWfkVLU39R9g9h5wPPSe7gvrJrBiMoklCTv8I=
`protect END_PROTECTED
