`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iok4kDiKBOwkmTgHgCfVjWGmi3DsJ64UT+h/Sk2idpFQ0Cy8dWikBIvfiGcTfIhC
bKHiACum5+7tmdCQi8gTsvadY7LJBx0+J7GPN4FaOt+/RBbszL7S3IO/5dCyPnVL
NB7HUmPLjwZP3cpintq33bnA0oYvelezigpGWKqVde/ftZfvQW+8W5uWgJ+ztiE5
v8bunMQdzoLMU5XglByQv0POPKN8vDzb0lvog16ZnKbH4/Wyt53CDTDDpEfk18px
KqHPe+52f87YsFX+CsszTxLV26IwC/8jw9yl3mJ6biqTZl8frM3+Oa5o+TI7xPys
APNQlmhsjR1UJABhI7gru/KnJP9mz9JF4oQBBMGMzcTpVH9ZFn5FEMVsPIevouPB
7EGWc28w3q+y8tW9YYrw311C98ObRLC4EIt8xrp2PN7SG1YCtOSdbai1+tJPemYE
RTeWOV0uBpomrW/IPAdmF3xDFAtoHs1mvhGCYYiUlR2aMEN3DGxcHPtjkIg1dnXI
YlMjk6/A5Sb5Yo7Y196UA4zUzylW9HzBdoUWFG2RdQUnf+L7a2XHUUBO5qxgCvpF
+jzRAZhgsnXRPwOVrRmdbUVIokU4t4qbLu62y6pLf/BII6EmE4V/vXBzuZ5aSpYv
`protect END_PROTECTED
