`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt2+ytJNEYREM8CIWQZK+JQH12dh8wMpCd8iSAG0mopSHlppW4Abx0rGxbwvVixH
SYtgdNOb+bS0AGI72Jhmpkb9bJY+V8qHn6EhQCWe0G+4OLqBz+isjtgghpwWWQ+q
0QmBt5dtdmwTWV/y3Yr1uGfdu0tVSwCyXA4EAJ/FZVf7xjRqfq755XtqycbRK2bl
g9oFhezGPpyuNGZzwThA9QZvk3Nb9/zOCktPzOHHBuebmKRBNAgQgdWp58vZsbfJ
KaHgTW8I9/IEUcJHWn1aaIt3Xtb/SetN1U4RtiA8VKJTPuGhSryGibnZ6RVSS3bR
tWHoZzQ8tKEV01XurHWulnxqeLiMgu0vwc2TFMG+FawVnF8Fl7NBT8LOReNdGgWO
3vaHAsD1fhNl8AlQHw7OKetabxa3DQ+mN9tII7qyht6kwPJl2XccHkC+fG2bYc8Y
6QSwArDJLB+do0HTXKHnkxnlzCaCYtrAw27u9P4zsJfMVOT0nhTuT7G5K9iwtk6O
IL7qW+SlhlOHeXcpTKx6EV9qcTo5PWSdjdfXUq0UqdD9dtJFzEZrl4twhsPYEJgg
jnqOatJgKegkyubB/dXNQjJEh2YRczDTd99vLc973krP2OSRstKtwM8rHPIFfkc5
cnOIvfqxKIlx34fgYLnntG9NCMQVZRGCxpJ0+1FR6dI+TjglSfFbIo1ZIob70sc/
yaejmyskHR1g1rjLmA4WzS1DVDGeTA1HF4v70yuwuI31T9mkHr+ngbRGKinOJw4p
5Cb5oM4a13RvU+FKUq5JwTBBlCfujM7yFaYCQlIBzV5aOcwaPfJwuf29Kod0sJ3w
rDBZKD+szAEQ1aVL9eHucjGdjtud/y1zDqk10Lq3EGpxu8UScIeeEJqcZsiUeoMX
TEsFET8nUPmm1a8/wT/hOUGLkX+K+9eVo0XS6El1Ar5yiaUMfFGFwzCIPg7M4vgU
Abi/Lpyj0/i1ZuQ3M+SVj8zBTQRassb8+9DJ391AdPn+BgJ8cqUjP5AykWm7hCEr
`protect END_PROTECTED
