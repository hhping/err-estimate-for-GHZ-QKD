`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lMoMr7V4Z01llUV26f+z49aB9r12zyNvo+3Ou77P4m+3Jzr3GXpCmxcvYiZBhec
YGlZ69quE+59pacQEDAAJf9VMDwaIFkDE5GCxxi2fVYOfX2Iq9s5hnYZoNCx85dq
PWspZB9ahvvyN8QkztsI2rWdP/fE0Z7mYYVm/hYBfW4oBIi18Np8Yqd6dqo3r8l+
e4k9V1S4cxj4tRnmI34O868EyGsWbTIiW3zpxQJhESJTdx8aOzMOvXp25MvsCJ0X
4JdTWVgpqOjo4L2XoaO69w9JUPytJtegqoTRdsmgV8NT5fNOwz3WPqHEsY6BGwhF
XukSFn/AricmfshLtpxVzqcXARe8UjKPTx9JSkjandfFmHcsm1jqT8QlmoG1MyFz
KNMNmqa+28cYrcQaCB36UBEZOHItfpkbFij+l4YjAiK3OKIR22cUdwbhm8QZL11H
yxbL7a9B4zbR3PWmOk5PEQ3CvQnfoz0jloOFOfEmEG55IxxqF1shfpwNBCO9tR5f
KsT/8UqLns6kQgVptfgZEFsoSGag5x+eTr7L5Sn1SAuVjllZB2ftOCswA8bdd7v4
r+K8u4VCn3XNmJqGEq+2brlXYi1jZGhiOk0QZJYwzOg7CR82Eozsw5bLSYLQbwOn
lbyyqrsCLC2eBXU5aReuCefz/DqzOUMRbuxxCt+0UdXPkTnW5mjmcVtPbZCTvrk2
Bt40i/70jzJYb16cAsR87mEPi6NNybGut/mIU226jzSJtiMK819oNso1YT3yyPCR
WtuwhQZp7AO+z460IceFZ7v/KY8eCyw0D69z1qs2NN2s99DxD8KO4kedMQY96YWr
Pw+5NpszwNnrIJrkSgLAD0KLqzpAWFY+GcsH5m4WUf8BFtS9R24N4Me0DQLtSMX5
NY8mAH+O4ZhrbynSHQEwEcLPxB8mO9Cth0DsofRU7jYFSfAqgI6MYFa9O02Y/8OR
qvG4pF/BPGLwt9IOIQ0iKiqCl+stPa+ZcoSZCAJ3r9g+b03goxvOnvuW3GpOCe2u
MWWCSzEloQmnGMvSOByFfq1FeQky/QK+Jn67nV60Jp8IMIwkwaliP5HBqA6NuEaU
NVDac9vzcNEFDTUmK1PSeIwpjUIF+qyy/FdLQz/2p6Nhj1AkK/Qoffu44xwRPSW8
n2ViYvIvKST0kWTVxnsAtJ417wVO/UXJXwZwv1BAfxx0KA2KuVO4Ukc8OCXKZtAH
p2C3zGYeoVjxnklO80kBsDKOLOY5DYNT/L09FnpkyQg=
`protect END_PROTECTED
