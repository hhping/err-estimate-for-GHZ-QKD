`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kU8MwreAuGDQg3qyxU2bz5c9jnpxwEcsIymEgYqbrIz3pa+aXIxUXvFyC1eUj6B6
c1it8WGRMXBm/9JPtW+iQMBhZJZ9+0mEhjQ+n5CULwn4Ff62a+cx9Ubgv1+XWDBN
HUeRw5VvwwMGrbp+guWDye5oy/mstWMojSXOQf4wBu/Agu2P1fX9Tnrhh+CLD8ZR
yBVpkmD+IGA6cpFLqtVh03t4rzew9bavKYf50wa56jYgVFGCphQzYwlpHWE+17yK
qANcPB3HeOfivJZLSsigMuYiXZ1bo3Z+wXexdgsez6Lg2FjuZGBjWVnHF7JXzDND
PgZcp7ecUWGpYcgBQy3g5Drqp5Gpiw1RfBW+FR5ULEXl/dL1pMrsaVl+qz0pf2vr
03vyFI7ihp3q53GiAClgELMYQNr+LvxJdFwA10blKY7ngQIIttknnLpj6XAvuFy7
QzIeN5WxQk4WdquK+Who8XEGlJaQV0SK58rFgbxlyUK6tCshQb3SqKJRU61bW40/
+U/IqjtDR+NLTFyYS+SXCOHvxaqHf4E/pQ38XFonUKjLSnxr4brquIUE57C1V6Lj
sec24s9g0UkxdtiCOO5nIg24OMqBEzlDHEPNkOz73CrkMfwfMPmfq4FSNmoC/Sg0
mZGq37KuJtyD4fo/ynSkT8RRJQw9E74E7zwKGmiJO0Bpwd3H+2ehyg3y/Kgjy005
ZyRCRqjIXnGSEdO5UqbBkPWpSTnKP51T9hofPwtDRpwFecyvulvDYluv/VGy91af
rjfvER4xLgBuk6uXdvX7xH7/RTHiSpbgZSjOEv/9UYripLYnTLRGJnJca8zrx4EX
uxH5A07fTeeaMmyO+N6dey7+UgE2RT34vnUC/qxHS9wfllcZ8UPMM5NMwfgl6Z7+
E8JKRS7DskHVGwKugF26vXCwPik/FNDiSjOKrr9CklYbfItwMJ9NArrE+U0OY7KH
MrdzuW5EabqsWcMx1jJ9aKhkOTciM2/IcYvaN4CXnH9iV23h1AsPbh0nTe/d7Hn/
JwgcDgSf7/+i8EEzHhwalbz0xMHgjht8iNgFjqJoR6nDiIKNGlRqifuUOT+2WV/p
L4Uigr27CNE5bfPsXCl8OXi/tL2r+B5NeXO3PTwOuQbrQXBzIEo1mRXq5AtJA1hp
S1z2N++Xv9/J2FLegHAvbMFtpnFpzuexZFq/QWD7exB3kV4lnXPTyi1vASSzZrbF
C/o2rBLS3Q1n+OBp9NnW6DbZHtoKHeYyuhC/Z7oI/KJeAUQ/9EOJUAUq2E2baSHP
P2dKqcki3Tmn6N3Hn2gY4SfWVokkck4f8AJ3U/2hTJ3WSrMKwB12aGvjvdnUhG3l
ksrDAF2An1d7h52jc23kxxUmGahY7rx5byNEofhj88ecQPd3Xx9W9S+Zg6yr0/k5
3njLQaFd0AEUHUWDBdb02XWQ5Ip+Mck59VdGI82YzxBsXdSTub68Cc7DAON41V2D
SF1pZwrhdr3Iwf9qdWQ+JT79XAtFum79FvWT+AnH23HchUKd2d97wcVHgRoIut0p
JI4LhtIYcugWcT6yF3Swop3L097fnp+Sguv9Hxa8rejNz/Xo4Gzn8MBeJPKX6dmG
NWBwY6uwCqDNOzyiXs1SNscIZFOuv0rsa69b5IonQ4l3TbS1FKaAf11DCMDo5JxP
IT94pukZemKjt2WOnMmLimSfy2tXRADUZzYK6R54eH+0feYlSF5CARGqZPfGd1bJ
nzzTW7ZZ2mnMBsvYOunJEgPIW+txVE2/PgT6hLoYtBm/Hsw6iB7IunJsulU1FL5A
qf74Ieu1n9fXvhLQonKesQ4gzXumGxtLF7bqHytGJ+wuGPpj7OWwHt779jSUs2si
KX2cOaJDrVf5sb6ui5L1JZgT4FTVy19UAT+P00mXzx1qmd/sucFZjcAxz5RAul5V
N6UqZn60+jS8MHCM43pJXxkimXsufvbUifLg0Moo3hVtd1FhvxGHmJjwJTXpXYRL
NP5fU8rACHQP2JmrkhRBxK2FvtqhvIiEZfglEpxWXfe9qjZa3ci7cVLB1wNu1aIw
FhI84hJmBwrwsxQ+yoTI+97B//lmSONqNA34KibGUgFJYNFPgck0Pjh+H5uzwcH6
YcxWM+djVkYLs0SQ1l2NoKrT4N5Ks3GhsgXNiaHZK/TCwHLL4OwQ/yGCs1+wtMYf
Urq0q729CA6b6ZbzatAHq22DndcTzQ9qQd7aq8ZWuIJdpiTBnJIyRyx7d0ouCf2b
QsxS4EQqEqiddOa5KhRn587T09UH+L0Mw/7Ax3Xjf4FwDDdtorsStptp5RLRaJMG
7RpvinpZ8LvHiCGqgi8MYUoK2NB8Tou5FwwO/uCw0jDn/Ncq7BMfuGAyJuvwIVp+
tHffArsIBQ3RH2mVLqavcX4t/VKFQDcxeGhGBV/4uROguLG1IW1uWzvrMVpBHQp8
z0nWIXDe6KeUhjnLpuw7jwc+CGSm9cBZ9HICFq5StfBcmqpX7FBq61MOols4SRjP
8WvqjSePsZpMJBwCLLMlzlfccjZPzhLQjY4Qy9JWBCIEUlkTOCvdHWCMCI3HJMf9
A1DIhvAznG8DvxdXp/aFPCV9ohUtjVIqb1ZA/ufqVVErdGgPnF+a0h1pDTSLJvt/
qX6I8dSIJP8OBPWx3k80EkZIi8uUph+xALQf80uYcJSInkPZ0/iKT9ti3VSDybsS
iBikM4dk6R0nbbyYKsXYIOsLH3d0rt0IOmOOT+EngwsdwRqZGXbpgclpyw/uvRkN
FuLDneDYknDZlXyqY3syeJ4VmvMgXZhg1Qsv3I2yu+YIO87VMWCnMbYE4JBZp9Qp
too+FMVsT5tu/R3uYFDoTd4qgnp9SFPxNGKZdUh0z6yieyoqyc+PB2AmvIXCxONu
P3h8PM/Q+C5+cdLyho3UDFokoBwhtWtCSWVKN8ODncQf/3VRGgg2die+NXmcQEse
FymcvJD4yw9Xex0ps/wzJPlrNri9gmOOzVbPWaNFe//+k0nJ4JicJ0Ir8CUtGwXH
HNc+m8z2t7TnYk7saCvNxiyRfB1fV1nBJPhOxrFlKIyCa9jUxQ6t02eqExUTWcWl
Hzast0jg1LQMKPH9an9GQbyTYBMoWDfBfcs9ydTSRGy07iYrC8ldQvN5iAr9TTsg
7VAAbRR5eOBM8nOGV4tBRKdll6p4+whJVPiiL7dccMYPkbyrT6aGkpmAyv3yvheF
`protect END_PROTECTED
