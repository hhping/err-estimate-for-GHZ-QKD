`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDfFKc4lhtwadfn56FnPYf/q7gxvBA+MV83Odw0FKjomRsF39EyT5YmKDm2WOWse
g9QDIgOE5u8nLf/Upfntxxjr2QHQT3ZH5WkPN+fn8SadDjWMcFM5cUiuHNV0VrtD
RVGUxrYHSJRRiZvSubEPATjUZNqd4sljgw2AOOC9451TW7sClN5L9hIYgEC+bfvB
PAcc49a8TfZI+y5/SBcgQhLg2tuT3/D8BkMGlg+334GTZKLAgI6qHtsvjSt3n8sF
zIVrbRk+0i3v4UFSRzJh5WYYiAdV346KwsH2Pp3LXEVAFCSwnYRukmh73NkgqFUG
G/iF1PjgxeJrA7wnrkRGnLEI2DSbrGj75g5H93EzVhGaSJZDISP/H0DNFCj/skT+
I5E0wsojjS1+U/pxHtg9dYU/3WO1CgJg3V08z4T/6/0gEKlzJbsP6vBodHDLohtt
AgV4gAfNYMiy4oLEe4NZXzBzJPZYq3wfrOdHFJdIxBuf+0nBo8+pt/omBjPOesPU
6hAyHwEtaao9hV8pXVidoLOI0jtQEO5NDtpcmLy+fyS+Md/P5zNyzB70VdwG/t98
ku2Et6SOB0OH05hnaoW5KT0wDlX9mH9disxDEE1edZHCEn4JdheGJvFopjqQ4Ilu
3NmUOSRXn5KgWUkD9sVWMc4AeI6BTnYWejPibORr7AL2h5anweHXABTGo4s+ThV8
0MAn7I8DR2X3IvZmCWUn4OERSe2OmX1d02W/2wLYi1nP84YaacK2Pom19SQ+Y1ky
/dnCIQjawJeGSMZJVwHlVdYxWxFbNGlfD/902yTQqJS/bjQa79f2EJlggVIu+A4V
`protect END_PROTECTED
