`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4z6bwclEoNMpF4TnkgGXl8rvvyHeC6HDa1I+ssIpaCuOHhPnxYK8M/m/yA7/k//E
ATm35qO9HR0y/Utto2vNyW2VpTB0IEN7P4NzqpizCM/1DhuBquNHNyX/Zy+cMgL+
w+yDWEFZH0wJE96NDokuNf3snRpaIF4BY56zuLkXiCm65ehR08J8qfbsRQiolNDK
DBMDwnmrQyNdeA85zTFOj2fS1c2ui1h97O2FmccgaQy7yC4WrXFz1sMgwjjZywfR
nBUNa4CqOgtHNQu2jTI8CQSZ3GH3FfrPVWW6rPTxz4O/vJtx9KpHmwrY6dsCyHcQ
fFhnt5j+NQvtGqAJCxAjpJ1oG86fFby+kxT9yKTtTRW3t80S0QzUDyv2EWfqPnUc
5Zrqnc3dwzdaK2Mw+Cjz/8ZHaDeSnIXAt5fjp5fZA+wMNeJZRFNeOAwEXDxbbTgj
RMaQIin1Goazknl0IKu40RLIO0Jfttaboy9D63A9cMm3DC6Ezoqw3Si11e65Lb1y
`protect END_PROTECTED
