`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlmovnzYOu251ULn1kKBd4zK2kslO53RF0P5eMpm9gzUsSZQPpdpCq1DcW/HeRTJ
tDUjtkI8ACAk5RwfcQ2SyeJOE3SF8wH+4l7SkpNJa9sT+22LKDEaWgKXYHXhP3KG
5MaWWSu4F0K/8983NC5P+xO06nabBoGqERPCeeVi7JMs+vU0Vp3SQK30TAs2V3Mi
WJrmHTZu/EX1QeFLjGlzBL90eSEx3xQ6IEzaP9zy6D+EstL9+ineq1HKjXkemRTx
mFwDuujZ2bCeJ5qIcZVZvbkgXFSpQy8tw7LUx1eAHZRj3YK6xjiNQQBK56dBXfYi
pqSMh5igv/XnyYr4BMU1Qqy++fM9ZoXMK5KMX94Rh/ac/BJxPLa4dpcDqrbH9st8
pVntC4A111m2HWgiGZE6Bn/OvtBXClSqVznyKCpSy8x7L4MtVQKK0BKVGSDTohpc
G6RlZhE6/AdLuMALqnGjph1jpUeonTqE1JbNlTKPrZyJxFKQM/RSaHdEdIdDgGu2
5On2dcLWWZ1uu8q6morYzRvfT7VEXj9l2LcOf7vWYVrm0a/ePNICV/WOhjP2F+S5
M+on7a1MMKPDZW3dU+iFuPxpg0FRwNhIF59xHFteIaokZwX4phxri7r/tex3uyOp
1QI+RGnVCPvtuoUl91yEX2LgBIi22IqPbMlardO1iHOrFBoT+xV+FrWNJhBFfK7T
syeEdbHjZ/t4cGkimDfMcQBuA3ey9LmIEaxA/hNziaq3k4MB1Fez0Ir2doU2G6yk
19l8ZYS4xaRNczRSjYmmgcndH0KQpd4xwJY5azQPvi+NAOs/gTz37hdvvlg0Skui
Tr2rIYowitiJ9GpyWIcz4flaVyq/gVOvLgds7Zm+Tdlu1flW+EGzocgugZAkuGYS
W5CZHPXdtYu4OAW4rmYoeALCx4ylmrm/hMol0stqd5AWPiGMNJ+Mb7r8ajfpHrsQ
+Il3TucHAdwza9IOhMT0DUJcnkYH3dfV80CoszomzAbCFrR1JSknL7G8tuF0TYFw
xvVMvosRzaIvewAY7dBD4xsu3A93APL7iESZ5n8LkRBnMZw2Bh/g7esdj7MOPRQA
D/3463s1kHY5o80VL8/aw0SgmSXm0Rtzc6+MjTQHghg7hPMdYT4iSnfLz38JjWF2
8MlAMrr/FJZg4CCXnGE2BjTVvCyWdVC3WGFNxzQ1RcCBh1ChnIPRJSFTBlKds4+l
oc+GnHlBzEjURepj7HVIX7LCEagRHQiJmyU8CUCHhZaEjdN/IxAlmSLvpdoLzPEd
nEFrUMwhUvgP+AGAujWzcDUnyLVJRTsrJ+Qddcg85enlxtQKU5VRIBYkbMJvDyY1
vn05FOzIWW4Zmxv4HvMgnQ9FnX/k5ew1uPUWCstNpghfhKPpsjE3/RDR/eBy7foo
z75dBmSoZyoqK2p8M18FpbayfnDikeeYcNGvSBtdDC7mPNCOpW7Yuco3xmwsMshh
`protect END_PROTECTED
