`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6b56yMWQ5H5wqW/+LVAkZRod4+x7m166MXl7LbJekxddEtvdoGrlCOpU5mwdZwr
2Yw5mDHtL0RE5BhCM5kKK+i27ZaksaSUvTirPs/EvAODMl+bzH362lqWEVqrhQob
UocSWjxej8pLDbdQOZxwo3YnkUe/UCN2COss7Yz9EtSsaQrdEbe7UXWE0COpxHZp
51Ctyk0H5wM4lYePS9OkYQ2yA0RV5n0mOmfQtboRn2De3ZuyCTBdmlT7OhsqZ3IF
n1frut7WkNOGhJRrqn8b0ubXQ9uAxrU1/AWBnpG8oxSoa7njr1UDOtuG97YSXLXu
UgqGSevIsaDJSsroRX6Ep1p5sSk8RDJ+ahQ+mNCSqEzKumtqe1AqFyXX6EYU7R9A
m443HnaJMztD3rUKHc7e89DVcdOqZuHGgIBh124iKRLbjj9aGvdCu+mGZeLpsHml
ETx0BHwdAgiAp2AZvncPC3xW614T1aSV0c/LkCGAltwvvmFSo+aH2rTG6C0le4pp
swEmeEQbcGqQ2HoFed2LeW3KtLktVsTwQ9wLhwc68yKjVyz+NLe6F5zsJDzOcgr2
AFzQtgZBq7HSZ+Ej62V8qQ==
`protect END_PROTECTED
