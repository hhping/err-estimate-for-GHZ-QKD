`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gm89e7oJyvRwVUNL9KRwH1YCWu+Yx6QBApn85GVjl+w+LHr2oJ6Bl2LIgeVJm3ha
wxisJ9dl7fc2nMYIIcBbkGoaX1aGTrCruYBTPoqoHeStortMCS5dPXs0yXjIc/xs
liodvgL7pmL0SVPwVugZLN4Vbr3ct02NQ+YaJXe2i0IwznII8lsDCkw/oO4ryx1F
jA5OkazzeBEDEa5zcEq8v9LLM6XUEOMFUvZME85GJRrcGd3rY2/aWG6p4Ae9/O1Q
t3knfBSGJJGy4AOZhv+2W8beofPl3cARJOfhz6j+DQ6hbXUdZ09Xvf2shRLB6TCc
GZ/Q44w1RsKdwUhCtg92wZW/fFT4KEceg0XiPPOvkOARSmTjuNH3EXBOmST1GvMd
c+9hDlcK/M58CeJx4Mf+6y1N1CVH3GAa3CnpEH+2erwO7LB/snG4PS9K0BE/3atV
`protect END_PROTECTED
