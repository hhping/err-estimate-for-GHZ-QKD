`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIX7MaC9irefi25CDDeu76I64ZTp90B+NyvrgcBBXZa+Rwx/N7iA5Vmfjmi6nO26
VmgIKx6InQAoiocJXMTaHJTXCl+bQffabsPUZ2iGDMF9fSGtNSeB1vgW4rLkgRYn
XXV6s+hmlX6A46xhWb39vVNznC+xtXfhdrczizihSCz22Su8xNkewimG5DNI1d7c
tqnkC1uAUyb6Q0J2WmWzlsk7UIMbIKPlBbvi5htNyuhnzvA7fir7Gjy8XdsQoKAs
YHEdaeoK0pQnhmIGh2PMYueoplLixHrsLnLdZzDp/VIHANfRS6wq0AaBTa3ST3rz
YXlmN7kIjFisoZBshe+msO8zkXdxU8Pd785ME7svjIkoIHgeAjEARMpbfJTh02DL
ZYHBBXjoLnVNBLXPg61fMA==
`protect END_PROTECTED
