`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vh/j3pmHBtHog2ClLhtnfySXL5jYLs5DYPKHErQLA9IL9ao/2xFhV4cpvjuWR2GI
LKb4EokigFg2dk8wSYUq7tzfzvp+wqWTfjuqCjr3lxNppAAJLN/13LKX+ROMlMJV
3KutDLFsTvrEBS9zq7i5m09G/9tXMf+rFjEKbRXFqEj06HsjcKg7/6EGdcweGPm2
+k8LOE0l7S9Y/q621fF4C8sc7TVV4wwwQJlCxDP8uR03sqQ7D2q7mhfaZ9UFSNix
wQo/zdnyXo7yZ8EVpYkGNip/vQLrz9H7NcDurQ6kHNMoyMCjjDIPCO2Jp+Z6xQFX
DOL3eaTHWqxwNoUMqNfQbmS3MMkNs3KQJBl/7OdOq8tblO0OURsjQAD1rXsIzK3a
iWW/NIBgJVUnbE9xYQ5ldKwWyszkaGS4wJQrfFuv4YkNuSsyv4yeUzEtO0XTVwnn
`protect END_PROTECTED
