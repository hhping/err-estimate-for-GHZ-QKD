`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azfAOpGvkdXaz+AIJusNWMWqf9voI0hfuqU/SdjhmwsgzJCMrF/DRYYGvjyJIC22
Ppl0ir8OEnsYCJuuagkaG9GON6s5shT0bKKTGJ+6OdPrai8G/JpgntnZH60lORFa
1F9GPWyltxLPUDrnBdXfOSMW54Q8BrL1ZFq9nVIQEFEGycm3D32ReHbXmTvep+Nx
GDeA2YUstLYJnQiA25RXFFhcRebUNeyNHb3XK3qtwPf0oHW9XPDvhdaRwPu8dj8d
4sP/2Kkm2lrvX3putbh7PKt39WGDpPcRW+cVg1C2StRcKLhYLNmmpZS5WMx3Qx3C
XZYakfrGoW3F4HcLVPeGvsICuMCjMNyy+9OupH1OmgR0GZ5RKqDTfIgladp36dsh
N5EK5bVw3X2Tw85vUYaywVyErqbrK0oMrmWvxD5ywgFX1sysCwPLZGnqqNgHZWbk
j8IwUxke3GnUsU+FWagSQdj7VE3ERc63rWwqXTpNm+2aD9BYJC6mX/QlCidBNEiQ
4r6FGvBvIWMQ0o4LsvVVFPj26BuVxtQLfeLxmlV7KGaCtzyMtHo7CccGZH7B/DTI
pixOjPEFnCKR4vSWWKueSnaRrfxqYTSD+9cMtJN2FLDkLx5hbs2azioAVyYr9fT9
3/YRBY8EmQlu96uWU17n4Xh+s8mYVeVk/+cI3N95aXAJ3s/vDBdxL/XyFhySwiwo
ifNsYH1B8id6EYi8cOXz8kT/udth1Iiw2tBbSPjRBVzby+njlp9wC+BJhi7i4+eT
fCXBqZEl5BLPfq/5bw4CkiLZGg5u5ZmjYL15bGz7z7WaZHpJEIP49sKvkB4vPhhu
s45Edk//8Sxg2MBdWQgGmYW9it35N0mdFnS0NWymfOEPcptny2Q5vWG9cc+DJq7I
OuK3yeJk0V5FGep1sl89V06s8FCPtSR4rVcJIvoalWeiJcDkMM5ha9Td3qJ7Iw8Z
ZWmEsZED6doamgQSYppySvgBnG92P+ZhtbMTdBsDved/a846CvoTvALZNsoDLODz
gxs5gZj+RjY4wDFNXNQ9GAR7Qr45bBCE1IUkrPt18EcXDD8tzohnWMjdym+wqw/4
4WgzhNllexgvmfw2Mg/6N6b9/ZTKoyMSYFQXVnsRYp5KQcQfOBOXPNNTYvj3kaO6
7z5Q3ETsAfgpayoDEYFHVLB+RD3OZEspl4EocNxGbQZFB23hIhEPxqdjRE/I8HTM
ePaLJNWzGm71rNwrCNX6cTMhuafpeQV95pwEU37GQTcMTpz+moKy1kR83Vy/F9Ih
L10HRV5H2l8PY3uP/K+SLcKEpWhD7lI5ACRDnZM2Zd+m8VoMS2bjc0N7ocpeHvFL
tDq80GCdbC47sv+0oqWjGBMcDSCQV2VxLh4oV07fNR9L0AQXSPb94rQVXEPt1Dn9
8gqQdRWgbGVzRr1mcYnisK59C2TmE9K1x/li7/bYyABMsR3QG6obQY6FkSa1vpUO
S1CBj2RMWpGduBCsdEB694ahr4pC40Lk3GK8SIJigplvNALAEwaOFSR0FLI2G2WA
UaPOO6E/Xutfxx4Yohejcu3JGEnoa83NiXAdiGMxJH3sNHNaMj2R1HmEHiQrvzht
4EZeIqOXnIzDxSPdoVKYZB/t/TFlP6bl+Cmu2fjvMzD7wRhp0ANM1guBrPucXbGT
f7mIq5Geae9L8LX2upL1WSO6ZG9gPe6oPe54F3irkUFyA9tNLLCTRy5cEXpsCvG1
kYqC0DF5bIp72aHmH3t8lt1EE5c6wsTyuOw7rTwCpxtF7hvmkGAHiJvtmMDO4/Uj
xfI6p937aPx97U+7DfKybetpoCK+tIEFYDLALkotXSX86GV5aXozmQTz82jGwUC/
6nOUcUTQUYmHwPlAva2DfFazSj2zg7Umzm4U5dPuwliTXRgTr+uR20DflNLdTl8L
v62V1t43+0szOOp4frCTeEhHVXWYQX+KtyOPdiHuGU2crwnS/hk9EFfsymfNbT2s
En8jAR3XFn4VoE70pezHV5OYJVvepGEHOh4waw6syFj9huy8Yo+f2t3FuKek2mHc
pm5zkC+XDs2VyKeWv/N0h0t9klnAV7yyTRZNoFNPf1yqoTA0l7j0QdSlrXD5KAhz
+ax6ePjd9vNhYkONR+96nH3mBOnh3omk44osIlglGOS1oEcjQAQcagY8/80xujWn
Oav5rPv3oeFjVGdJB99ZqN88grBPG+TSQma0xMei68TbgY9c6U6qaNBVI4t+5/OJ
utMlOFx5elaRdKwUe3IiCNZNb1iPNSrBoddLKElM4MejUCS8g2TYrXCN99+S1JjA
21KQR0ybAc3V/ZW+nMuF8ujiBBKImd2WWkDZhNkAsG8ideeEwa6or305I631SD87
wxGPXzrbS4OmaPCoKIpec8v80edwQYwXAnTLgw7iqSXzcHRmoGHLjsX07CO9tjsX
XrUSAPVj904V81AeubzUFGKO4kTdywCT0qCb9rR0fbx/VfttvefrbnQQF6/3W3z9
2MRFzFRVE3Stm5PPuQX5sEBWwX1gusAa76b7EAkYpQFAKqWvzXalpQ/nWSjwtozG
UhLZfeJRPJPtj2V9YAdZnDuiycyH9v5g91mzQdoxRFlq9B92i1vJ1CCmNsl3HYod
GKfoHACIz/CXJmHenZGWaA==
`protect END_PROTECTED
