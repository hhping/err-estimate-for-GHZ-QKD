`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kRHCOyFxTeqqy3nMQs+wbgXUm2R+oR2CByfCLKxm8an7z3PNIwUJ2iHYFFaXYF0I
xZxlBOTU5wPd2kiNUyTsF1GIkggGbcfVtAOFAX+vB1SVYnNC22XCs4kPbMTTa8WZ
uvGQBQQyGqGPkhKiPJ+OFg1doH/jPlPlIXqQeLmTKykWwEWCXpTf0hjjesqhZiCD
ht2dYvd+ndNvT34qOXqFUDlzpUfBA8sRGpS4R3nzTOyJjSOv0lE/oPUpERpa76V/
aRL6dsuYJGLuoU4KIDCT69K4VQsiLe/IWETy792UJt5gCz6HDP73GwGi4NM71js+
6065EP3x1mdAW6tNxd0byp1KrxvVqMspCM16vULPTOOrt+foABSK3xLAvwjpjv0C
5E/lcGNL2LInQGejLBIIFg86g1X7JXJskes8D7IceofosC2hBM8mXkKlrdUrIuCK
L+9bNRmYrSLL667nbKwMqdRdeKGy+XWliomV4EH4DldnsHcqXEr6vqhcEcazSRIs
zZW1CiNlLkTcz+n2MPptevGDvdHfswPEP1uzU/eDPDtHkefR2wScNE78NZXqJhNV
QQYxz6Jrsx/O9zCwnIpIfMVnLF4jM8S5xr51Qalt8gwRrR4sUhrydC/3mfyGViVf
8gohSTiqQiZsNsbV5lzUxjyg4Qq3PduFdmnZb7t6zDtB36xl2v7GVDQmfLX5W5OM
JHHgJPo57MowG37zmafHOUzBqskEAXcNufMo+qt4uuZJtA+brtgleS8qK0fewqoZ
pcVJT6SFtkWWbrhZ6FsD5rnEpjzd3oF8tIHDX3EOik13p3fWQ/Z7AwQUVTITbrnc
PF2GaQwGAhEqE3/IdSQWV0VO1HmyRFBQSyuZlsJMqIfQagfVi9NnjGmLS4D/V7nl
awlfLHan9yQdGEsh/CZEc3AVjzerPiu2tMgZjuZGtvlE0cwpsuJnJMNliL3JkpRk
JI27Gv6ik6ZUzgL623S1iJHyaVVVv8ZorMfsO24m0JdtuGxWLvE7Li9R+Wgfljc0
U/848zKi+Ys3GuIXJL8QSKLSPNIx+rWHiFKn7g2sj8x/S8VKuIeGYksa1wa3UJr6
NXmZOTa4yVkZsQqkFaxmXTgeNwMlEl7impjwXQHnOSqfmQvXs7l9JVauTM05ySrv
LQXLC28rSnNdvGL42dp9aloXPz3BlJJN4vJ16XMsYGrfq1AgMjivHKv2+6MlthRS
tcQUET3fjC+tV80R8KOW3qpftTjzrJVfGHNvjWwlCyofpyFJ+pJCmvtMOBh94SfP
rivxV1uk9ugbr9A8cT9x9ecNsWpNbr5YqYmLgg1M+B/e65Dt3l72Z0gtZ9RFbfCk
5wQezgjm71W+/Pyatow58uEjmWkNx6NzWQJX670OPG9tFWgN5OIyPLJF6o41FQay
iN3MmJV1hFHvDJG56xGCrPkHjwovZiBE71u87FtyxcWL1/o0wN84PA45e7FZ+5Hc
19U0QdUEF2FP+ATEqKowh/ZD4lBAU4gAE8PaWz1QSc7dRD+g679Ppp8Jxxct5zAC
titXSzr4Rz3QFcKf12LDrlR4w8NNAgYUV9T5TifXkI98Ctar92u3v34uB/lAFTk6
KfpFRGbtgX2gPPFT/dL1p32CMwVzZ+xfKW9KJWS9CSOgAmduhFXPF4XEdyf6ztMI
CvNVL6fJ5BYDx2e8TB9y9pN1kqFgYWcuVtULI2rzdJQ=
`protect END_PROTECTED
