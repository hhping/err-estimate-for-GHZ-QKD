`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1z+FmcM4e7yw9hpdPGQ7GASEzKARqJwbw/b38lC3Qqd9K4D2dw/auGzWIOZmmnkE
mL29bCkF2Uju1nGBO4JbqtcrPsM+fRe+aPu3rxQvMCgE1hqoCB+/1KuEzOJFd2tr
4ri0uPGCAX1qdy/xU8j+4oLGcbNaWlW88+ETfP3w2BJMys98m4Xg/BsFZR4g0TOq
NxKhxkZTBAvVF0t/zQw7qKpI9gPCKDVLgbL7muNovfIhbWuJJS4K0cRrMRIQZW1q
19krlQhYKUjPerF/mwZDLqQuj+0sUBDi6aOaVFRZXxcPcGJV5USpZkUiqKmYbcko
ZyUPRYC5wTjeQ8T61k4hBB1glXb9sh4rRNe7UwTZNFbuSAIEorsafrZRfUVW0GcM
Sky8zNyj8hYER69vaJFS/DT7ULviC5zx4RdNAOib/UnZZWRc5okbv378MkQ2nxsH
nhVvehfTdtk5bZpbWfb2Zna5RlHYWqc/3YcJAdq2+33lnKYABPI8u/p1xyOW17n0
VAbm+XruRE/k7bzgRLQ2EcQ65uyOTAitus/WKAiVqpNf1J9nNcD1cY4WkAxW8cbh
RxyosF9LkcHupSU6px27CZ0qMI9rtTK+7k4gkXzeHL7JXujOP/tbTs0cm6C4xyYF
ltdMQPwNBZsUijUujI6eSZ1nGPi/pe4WoZLJkEpV/UlES6XNlYazegvqUFYsxiZK
Dmgpun7oEvAbpys3EbTD2xF/8ADRvqqXcZ3x7qYQc8ZQXqi10dDaPucDhJpSHq0J
DzNgP0ekduDzH/eadTC8ugyNdz2bUUlEIeuPv/TO6vkRFy+Igbu1IfNImSXG5V2u
4R6DURHCEr2OO1VH4mfquaY339ZxltoOW4GK0ejkJfmww6fVI9KmTFLFI9QzGkW0
8n8c/46ohbAIlv6L4QBrgwJaak4toXS5HPj8CJ4AWBg9s584ZjxVLNWV3lTeOMvD
nw5EKCDzvQvtISch1lEWg/vDMuVde05LNbvueppYpHldI//C8F4GNE0c0x/GvCsf
jwUr2iQH5ETOAttC8FwXccfaWlDw+EFrD+kMlPwiEnQhgJkRMYwq64UOLtoALdF8
11TdfA2EGXjZLSzv0V0GNInt2P31zLhMyYHR5p1hgf3MkGaeDKlUhZOlktSzbzHq
24SpEWEOzIGLEHHjiJw7lGylvYeTkFBU8Z1+4+HCf8vrONbGhLVVGJCfXYrc07kl
V9NmFQhS5v8dj5uS+YBofMjNWu1AKRVL38BExKq05vA=
`protect END_PROTECTED
