`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjFSu16oEsQMQnjo6God2bymZdc6mnqv/9jM626Z6TePeNvjfSpd49j/qxFHP93r
tlThZRKYy4YIXSQPNKft/wQwHuaCt79l7PfEiZ3qD8uCF5VV+7QIo2TCCZp9d58c
TuWGLtfuBYK7Dw3n71RYKlGAyW2UV4NMJXjwK5R5kT+um0ta5snoXUkR9ugM1Hpc
0uFwbJby7wWChO5rkVs4JG+5pmb8d9rAxut4pQNFAaaeKU1TdvYsRp2yp0gaH43e
jtCTOuzXaV3+ygS4SIpXTqMyiQ9cXv5drFT3fagGj3aR6ejaQ/ZZ6cvb2Ll8V5xa
Q1KuioZm6cRRoHkt3knKRYa54wpx/BINQHFIyLs1XtYJM/1odewGoAi5T5na1Wep
ta8EIJVq+yyWjjoCrQWM0s5+wBTLGfARHHSSDET0XWgFD/qxUpPnvBYOL2PqhNWj
yDzT30CpzQVU5VwjCbfCEYbHXQ2riHux+JTqVgDTcn0pODu65uHYqzU/Ggqx+gcq
yLmqB9qlw9EGDsjZgNxKTjjhioWUzwJ+tRpfVaizdCH2UOcmWfzUVRkjA11n+yuk
YZgneWGJ3ZUAB6TJTXvLSkHQ9xeivcA9bJCS5APPbeQVErEnklnmdjkfUrgCrImz
mjJXMFnRlRR1AbZTpHMFOHkDBIhFIBW8L9IjBsWJ5TVMIHjVRe3+im5tiSWnqaAl
XzBUOBIxJxjGdt+1b0NI31HYwRogRUiw8Ar20L+fUnpzlbf1YqzZkbVHzoRu/xDY
iS/x/8U2Yv/b5kzlj9z2G+y8+0gja7e65K5kIXG4BT3s/mCB/bwUNiVG+CJy0qmt
lR/0sFZ2yIngYnoZMiPK5FhQ+TMADeKB9+RZpko5cb9klh3n+k3R+zY1/dCeNcx1
hZz8byDrPa0YpxYJx1YlTghTmeorytA2xxKtuV6wUzu5f+EzWCzNmK245U0LYJun
sXFXMVLbZnAzwzTUDQ0GQHyie8fZivuZzOJFdDisQctournpcRjeCRU9Tq2U2oPQ
4Vi8k+Pfyi0+SeLrjF7zg6OD7GlzGk1frlLAVnQ86zK43eo7FptPBFwhgvfu8omW
sDWuW9AJqHLC33imxeyZ7wO259RFQXNcIvBhD6/oHRMAXw7aPsyLbd+wWwSK7I4U
Az8RujStpfbVRQJRMLldnKYkSFa3XpsX/pqLuI97zI+aYuRIWb7IGxnMTlnC9dUt
omDtqcD+J1yUdh0VhK26wvMX71x3pyqszZ/SKkYSjMeJZFV4hpVtn/qOdRBUVAyp
9zY54SJbZsao/KjnB3F+MpB17F72TUHD+Cj2gmicsIoptBYHHABPy72VurMCWJRC
2quxC4rELPMxutLAEySmVLSibQbLMmVPLgqj4c3tXssGqbMI4wXnhelGJ7rFCNPQ
ioIZxqvDTNKc+biIjxWXQC/BP/zfAxFgW1zFbUJz+2tEvPH066vmeGrJqqnKOYJ/
B1hesrW5/tHujmcODNq/dgCZWeCtjNtLGEr0aXwpqUlU4s5Z4Zbu6hAHRlAylENv
mCWJ8gX+tBukUxOrRqwyUMS1/ChNplR7FrDgUz9qEoYij1g+vwFYM0Vg2Wk/ruaB
mp4KYDhm2KGPYYa52pr3ceKaHSf+vkPdfWTHEH8JeefUZD2tBGvQYcOjSQ47TVSW
uaijk6UyXuxR7tO0rg/CIXkmpf6hd9dafh4CPfRdAPcn4SG5zbjhf6lSHk8oq98O
UTMDnUNVONF/+JxLKpO0U21S/cTzfXrWvu1d3UpwRecdYugTmhvlWTzuiQ2IsqBB
ASyJMV3OQfD92fH/b2aA9M6kBHkFfvaFP7rCAs7sO1b0jTzjMdDNRoh/skrFgEyA
bLZE7mwWVRFG5gAY/WwZrpcN5ymqU3LISIzUyCjSC7LW1scy5Tran9IG+Yy9IPQv
WkgkNFc+u9saOdi9yTvhE/H0O+G7xkjpvHFlrZTH7NVGHWd8mYHu/WTEQBvwOTlu
1H18moVdgv/vMxPmairHSZvqfSaLrxfKnu9ANGe51Wb61z1vNQf7aNUnM9NouUNQ
Lt48w1mhnMwuF9GPgIjE5lbNsP7KB+hahr6D3pWDz9F+3lEZsmp9Swf9lvW9z73j
2JtwoQ9zKVx3dEFJkGoTzkUthb4pF56Be+epdTXuIzxzU76sOng6r8qUCSgC2dSe
ehvHcU7fUZJLxyr3VnerVpSbc7bznBsmyNvgfWb1gJuYqekr+zJ2GY/lWPejBJFJ
r9a1lnv5XaIA7VGZdzWSEnNoIRHPJH+UvCvOf9Jdvhttw1IbN3Fboxaf+oyM84fh
SNKnwisRZRG0gthVd7y07xx49E5nxQygUWaqTYqAwHn2pY+R8WGevIAoC2QHxGyM
rkzXiK/OeFUFUUmv+SljYyLeJdlGM5HXm+LNL3iinGxHoqX65ny+8BLuCdGBonKe
Ih1wELKkcL3j/jn+IVcOIeo3s1O27axr1KRHMgBP0zxAp0GKgFNXMlYaX8vexY2i
3VZJV7yyG0GOtDqaFhDufnWh1mBOQoppRuPWsvcH7c3Pi9XsVyFz0EdclVusFntF
hL+gimQ8aGTiaNekPPB/nrdwj51t8zfKxh2HdxVvf/5k5eK4e0HJKOso/JKG17Zl
iD0wAUNHPq9YkeND2FTyoEpCe//euUdtTgRa3l4ilk0gZo+lVQ19XXvp77Tkg6TS
b/RNMUjuIWKmbcE8FuhJMFeUqmTOK+Bt9GPEY8ToPJ4E3HlCylo6tTDO6eURRV+I
yu/hd8wgffhn7Vp2zc1FbLBdDBVABdTLn7ZxX9NMetKs759PpApPjumP8lUF7Ppc
W7lvZgKoM2YLyeG1uWeQ45sLeUcD9W+3iXnQQr7rwiSqFSSMdNOTAgI7ud3D9hVq
9+vV9uFGkppZg/Mt9tALCIuKrKwsgis7qY7ubLYclCpe4v4bF9F6tVxVClZ/DahD
VoTYoeXJAA5gaK7eF1WzeQuhkxvnvOMB07UX1HU4ey7zYlSw2c1HO5E/Ag+ejtla
jdHIMiRnwCDMxgatnjxmOmy9OFAKwB3RJGGVLoBlGLWRifxq5g52TFtQpfpd5Q7v
egITMiVRHF2OuxF4L3AuRPEMUUgSSCBIbBRIdIRczOeK9F8k+V0J6olRJkh83NK7
8PIGuyBhosG45xhrbiCkK/F6SwEhO0rFVsSnv22VBsv4HkGEcDKxZQBtpj176xky
inyk8Uxe06qSF+O5Jl9szfDNGu/2JQzyOFyr8vDTZ+HqDoJ7ApMfriADo/Xo0X64
GrMXIT2HjaQqHii6pTtJco34ct46j/8qMjUEFORD/9QuU4SDxC+qoCCGkk/+qFXq
oM3M1XCvS4OyFoWmH1g7phuNqRZqOaw44aqXhUUCvbeRMpv0W9Q8pjmRPUzwritm
NZu/IB2B9hzwzGzzc2FkzrFKvZyiYh/yjmPZsNwOsULiueJ16AEZg7WfM3ksx2aT
ggZ2E1I00lQQ7P7BQpV+i8iZKArlVhUC+68MRUa4718jlXICfkbzXs+93pm7oe45
np1rjLtouBQF01u51VHroQoJbrrAUhmATaY3ZuUP6w9ESVIY0hzHmrQDZ5iH9blU
hDTXq2xKTx7cXb7LZF8YNdBMQR6ramMaQRDHNSEB/bFZabyYBOOBruEb0+Y3+0os
arwXAAnyhljDbD+GRJJ8HR3upB6AohjdlVZhj4ZoaRMFS2A9Jb3SWB8R9/5E+bfd
e75egyn2CMfKvffy9BbbDBPnXySfI9bN5ZhKuToD+FnTVU0WPs1w6SDBYggFv0wS
Pcxua3FHWTUBuwuzHluoxQ==
`protect END_PROTECTED
