`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rkg1vRAhoZV2d35CWrSpeefF6S5IJ8REAPBPVmDmk2aasxAv3wsvnoY7W5qRMij+
cvxcPpAKp3qQIhM1AvPr0DXmEeiIrCKBQiK6MwZQd02LZk/GPBcgxmmm985C3ewD
4PZzkTwEkrvkbvSjjhirwhBJMI5ur7ZQT8NgkxOv8i13kZ4wNTz3d5oKrxRn9Y62
h4kukalbwCSX4vCqMakRKvZ28RITo3nKreHRFP0GGvz0CPpiOmwePoN1p4s8DUiy
7YY0djDfFG1/6OQo+zxA+2MOZ3E2bOZ2W2ebi6k5m3ZdJh9991NIoYyyHaKZM5LP
RAiGTAB85ZxzG1YST/qvrz2M7GpSV4LbBbAQaePkFFin/k9azbBbFqbU0LSptALZ
s7tT46SRH3gFqeCHboLRbmAVALQFgt+WO0LARKjw8yiJa3t6HmwlPwQJVhO3/hVy
Vu0wjxWlPsfKOQ3REL2lYrjJsItbO+0eBtK1dyvpMJlAWg4VQtbI244Nd95Q6ieH
PB/zq8BOPt+ba9TvLEz+PkkEwyof4j3ieqYdxm8zl1rdGmeF/TMmG43ivEO8GqYR
Gd9enuA6RgcKbhmIINIGcWLen1pfJ5d46bMGxVhjem2XkwOTqk9g1RTxXo9Nvld5
Z62mEYU3iv07TpI0ye2wnNnC+e/9/t1IGxJSw6DGvoVDVby5DgLBSKGwu6X8+hsc
uNAdZ+lrxYviKifD4rW14fg6r4kC6uKr+eCi1cgvEifeid41P/52Mz1H8Fs9pr+i
`protect END_PROTECTED
