`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
co1af4DHpdT4MMsjZLsM2n9mMpNLnte2CsXJS18Y2/myg/0CpH8Ayl6Npl/9K9uO
NdsW0gVTIaQUhAubEahL5dszZjefGiApiIXgLxyn+8pypPhBBQQ2DgxdkgYpjE6g
yp3dcHXAJE7+psxr+nyKA8U8jLQKL1wOMRMvOkpHgvlFjurtEpwYIZ7sFQ7R90wa
TVXnkF6i5v//8iJ6tgzb8qy2y4A6fPSLPXpgweIN1N3ZndOCCQ3YKwt8/YaZFOwp
pr73W8eXoqLg3GvPQM5FfG7N3C7M8EgcTFXNjbrgmGqD1PlvhhVZVJEK1qrZ8L3w
uqm70CuvMdPhRHNluI3xbuVVZzFw7Wk1ZAfZcB07TVkJQDZMwa6FYUae9lwIUTx9
6i/VHp2GsoXkwvutEo7Okz/mdAZAgI+iFC5c0qo5SupOVBPfetBVXagQj0GwwrMB
pa4rToC8NYiekzKuqveUlMghBALEcpqoBjXyTwaGT0Ik8a/deoWIG0RtnURfcoYg
ZKvx9cNhUpguis2G1klloGAHv0TbvNJL/eU1ZtogPfjlb+UcP7vCtsngwCXcMLNR
rRrOCpoYrS8zBsqHcJ6Ajg==
`protect END_PROTECTED
