`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S9ztZfTIUWVlr1+Q3bnv51e9RKFWTFuXBqFR5XexqZ+1OuMqgk88jWsYfhG23Bxw
BrEVSkLphllRCRDhJiB5KN7CRXuOR1WMuG6JOA6CZvUGI9ttFgRUmWMq3TSx2XmA
eHetR4sGVer8O4v848xP5uRsK4BmqOsIkN437E1PMiLC88DN3xRav5VfRaGAsyGJ
HWEJuknb1+qqJBrxTnbcrCJB3udnQI9UmGZOmbbKerpGc9KEHFB59vKt23upwexp
YLX1YNDbabvvGWTP1YtQi5C9yXGr7qiuECXQQ7OFEyOEkuqolc8qte8nVY1u4eOg
UjxT+kApSaVJ2pvL+gkoe5zkwuEQsVqQGTuPWTKp8ezlBAbUYc/7PF7h0vv9effy
1ADwXiqFtWq+En1y9JJgm/1vGPbWRBHtQBsUhvOpRreep2r4oNOHsZLiZ8XKFIJz
dFMTcw67uYYAejdFIXI6WOoKxoYl2FiWAFUHPuRgo1q7zKc032FIN/uecKZprQPS
EsA/n5trtPnJFt7UEwU9JujFGjtehIsLzcT3y/H1zNFrPo3Y3DJpQOYffolkc4DE
aZZklzSmlpZAn8JVBFugsyfbwjUKwr5sI68g0tzPXW1cvTdXUlLxFu7SRWfo4KXg
RffEma6HmTs0vUnSTHJkzE0AfKYBtAtw57o4WISZ+xYHQm7XfpDLSV8vB+hsfxao
KECfamm1aaaYtV9tXRI8juXunlr100GxT7qHFmYtohfJK0dzg4qRM5kGOTe0NB7i
1+Mwgnk74R+qSEPkRES9YdFAfqY/GJFzqhb1JQ2LX6+QlnGvWVVR9CqBn4QGhojn
CYLw4rH33MgsKhcUI/5kgJBbI9dfhUWNvJfM+qcjUn8irxBUZTN3uO52VXjHF+eU
`protect END_PROTECTED
