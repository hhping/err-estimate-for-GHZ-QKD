`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3ugIoh1UL63nE0IJkZUOsQG6XR1dbXuI5wyoS0pzucMRmI+WokGYImEVpheM94B
ZxTFZaP5N1wUn6WE9HRCBOir70Z0wpPyIVHtSvs7M/7IWQ+PGKCq0zQBjvyMbOFE
VDpOAZq3dBYZtXnrlNOYmTMdMJKI+dA3gIo2LVWsVmJ+NHBjevlP5Jn7PYzq836v
/UXqopn9ePnSvozBemwxwyxZTRms5/fyDYHSP9AzsCfiuLLyEowH6FSFtQ7Hl3Ms
oWIJqOvSflbLXLcw06+sRLggj5jkNij2M1Jmyrzhqa8QUKnHMWtABgomONNt/w3K
qN+bTpADMd4B2zscpjonnKznAyFIt4OJEU3wlNEmO8gqnMTTAZ2SgcAZ7Z7VZxGO
82KdAYcGlOQd4XfzHmJBXR0933WoJJyyb1QheCOxn7EF+DgS5K8KeH/xr74Pi38B
Y0DjT7CVagRWTe6KD4i24ik2z/5Pjp54N0WkipaTgEA3lz9svx7fXbKT8Dp4tH9i
BLMHouDsl1fkVZ5k9HOlFImb+6JJuyAQehsBfA5u2bIyJyp+JRF40YKojunIrZDq
mSCASKDt8GT/uRFJqiypPq3ExadfT9H3ajZg8P0h0GjtgJbE2GCETQEG2qyRHix4
ey6vhUxZ2BHCe2KVHxaLGp3YBZIOqUSlNUi1PFPhUDxbdBoW+yEN6VAZ/D3G3qsB
9pK66lBP16QnzOGeUpBJ1No42hEQv28BFByM9Yzks63BHpuVA1MdPFdjoCTRrp4t
MtSVJ+lJv8xTkCUL6/sEhYtX6HynW8HOBuaheJkoaEl9s5PHf69GboRnR3nOzUQ9
Mrukyny3g3nB0KeFV4XFMs6PXuZkfsF7oGU5MyUmmi8W5V1iEe3P+dn5DioCT2Qj
byk8Uz32GD9J9IbIT9V7Z67PJx+nUoSAiyOfM9rJjXKkXuNQBnZgOzxBTHgp4LvB
upCW+1RkHuTJd2aOi++DUgWwXrQwQqX2pKGTAYqmIO8Mddpn7Lwp5WQNLNWOe/Kz
yOdsI+mLupsRGQKOpzggef4ZNsra5pvvq58w4LSLSPjd0FnTwlm4akDzJh5dO2q1
8b7GgDyCFd1dEmlDY8j2cqclPwM6yTGrrXek0rhq62PNpjxgD4Aro5XsL5g9SebM
pYb8e9JNU5nDbNWItJqsFDUOPIhXrph1oT3t9Le13SEyNvxkZ8j/qpBygTMZYkOk
v483YI+80o80qdCvL87YVp+1ufTJIm8Mult5SN6+Lah/UBmOuCtmpsWBen2gghV7
hoI/M+pCUaBJe6boxF6cwxT1H4k3OrVvKTxYOwToM61aQNb2+AkWLIAuKWWQ7d2z
CO4Uv78upobR3BfuuI0FFa5asWvQByVJnlEiF98MfdjZPJecE6/ciRIn1xp6W6p4
TeC9VOwcEBMPvz57I2IjRK3549bE4F4Cyt6Za5S0qy7PHkS4v2slDh0F0C7CVCxd
m4rSXHuIDxtyTdaS3IQg6ZqOruLoHyd/V1FBr0mTIfR9OMUXPqfSzt890bJ+NPRP
A8dLww0UfEKtuLI2edc5jXSCL1G3ppnkNYcizJciEan5rYQFN8XnjD4miHl70gHs
OchX2txGSgA8b6geIJbhxTCjQX0/iRL2rxLFHXSq/t44j5ou4mYZ5HJdpaOgYvyb
4hBBH43HZr3klutOMnF952C0+bzVlmzd7QWJeYhjK5hJMU6K1/7QSLLhBtxwHxhU
WY6pYFhW4TjUXf9AtdVenHDeZc946HA9BMALe+acdL5X0B5+M/+4x400HZ8bjJND
ZiykijJ2bwiEkL5LtfYPkImFBxm/bVAWVI1AfC/ihNlM9F5ZZay/F0Sudq8LxstJ
OZGzM2qCIWWdTxan/rHkySEQ/p/mySJTxubgAjZocPhjFXPI6oN40bkRuHP6+Hpu
se2XnwGkndBpQwzR+a/Cf3mzVoSa2l6MFNusgFvsC8nR1J2o5W/+sA3UJnz/xKnk
3looft127+tgGVpZhz9RgigzHM5jHQ3vJPKTltsU0EvUE8QR7bDkuN1rD20r50PY
XE9C5kFj6f859TqsvG/SgAk29gfYhlC/ZkTYwVUFK0ZA7dOmgQnoW9QrU4qrk2IJ
CAISBHGnpAtwb3+LMUoIqOeecJInBIsTFhTOFS+l50JyQkkwFgNiniqswyQOv4id
PD7v+nMEhJ3tKaEFcQqpvX+8YZ6jVog9EFAXnCUj1EZTY8vSooO8Z4mnuDIVCsRm
swSYNmZx6czr+5Zxe/WEx1n9iC8U8hnupNMIN5pvft/jxG/JM8zAmpRO8gA4BK5x
lCDCMPIaXx57xZFuhCUWS7LcSjEaCxFcYx3hBrG7lxaZzyqkKpfvEUxG0NZIOYaY
0lI4ehplGIjhHCmHPHm0usWvOtb5YPPXUTdiSvrZXqocbtrNL0TttcDG+QL8x4Ww
LLzGrmo+2h8JAS6J8mj1XC4PUUUrabL+ewc6P0TVe5Q5zcaHs0bE580TR55a07D2
L5/C/zTCYaZLHSYj3hLJS83c2sLKVineZDT26VARpTUSC/nS9ny9QJi/uAu0dZ6B
tUkerZh0ia/TNCZbGB8TtSMXBBj6rDr4AVU2u3YSLgHCbrX62jILTGmIIguEnhUq
4rzjExZ4Ih/oX6LviVDHQbjwGrpE5PzzIJD5zi4sOHifj4OwCpcmASbO02TRihER
eFl0urF6WL3qpmyumbOOKRP0t7CrK1vm1r9T0E1urOfMyCbJQMuN1ijfImBUateg
k4+56hYAXWQujqh+DfiUDqtOgO0OGJKVBd9dAvpTPaNI6xu4MbuUyA63pfMbyUey
coA1X4/ielxxVtcfDHShWYLAKrfTRILtWcnqVm1xT2mDGFRaTuBDx6jzN+a3U7dZ
W9QjO8dWaAXTNaGWzDfO605ErhhyLjnu5WwHTfA9T3pkYIUUl7A7dmJFD3sDjIse
c4Sn5nwDGkYAwBTiGmlmki9WUfX65G5tsV8vyUxPxqnbQ3gEMqOd+IKpMd8UGjpD
hb9ikpPd4vodKlfPn7OivJKZ3DZIzna++ZpidV8AqELWdLYF5Dgk3mtg/FNmQ1Qs
zuPbrV1Alx4epmHiRfluUMgQhQofR5gsQBg4XcfIilU+AKq0sV1m61zuNBKdiO+a
SqnwfrmUfJb2O2+kQVu8OO6dqmmbxWOqVFXd3N6zobtL/DkjNA1JOay8eh2bLWrS
pdClsaOcKZFZHL1XBoiFi/eSiMsKVVVta/nEHBK4EFWBzFSyTcHZunWfXSBix+kI
`protect END_PROTECTED
