`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5YA2ASZd3HrmLkRJTg5nOpkKkNm8kl7mGSgABKVhsPDLhKpnmorG5f0mSlwv4Pjs
pMATNcTtfTmuiw4FzBLvuWnWtUgT/lgr1fq8lJLcEj4CIiiBrPtb4v/vJgEu7mdg
smEIjnvdX6Sx+eEjY0k+P3HV3TfclfKoEreDIUzXXFLD7JviAuKqJmkRALytT5bx
nKK8U8DR1L9Vo03nrBln6d6nNSecALaoFH8qQAGdg+xxy+s3XDMazjczfSEo5cDj
086AzIsF8ZiPQf2GijiKpwNbE2IW+4EHD+xebkMWx+DNTMJtrGuvsHaZZDXJcvtE
se8Za7VqJlj9EiwKBAzxPbmfyNzS1QsSUYeI7162bQIZ03suIdP5KryvVVmWk5nB
BooNFtPSa4rlRBjP80xFslHb2t6y584HfzKgT0/ktFOXjr/PRQDU/+RR+KYpJFIx
eA//ev03gLl2r3oGwWH4e+j5PldtKjTL+Cf5jRU0rvsS8Qul8eD1W7jtfgWvJlDz
`protect END_PROTECTED
