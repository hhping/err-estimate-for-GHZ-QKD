`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxGviNMIwux91PLVYIMwAOxg7yPMr86wYHK27QElk4JxeuPLEwlnEMRrN8KpekvJ
ERzDC1Z7bvS6LjGVRcvO8sXi/SbKjl+57VV0ZABz0mvFJap7UuXqW0tuI8LnttsS
DSUHGhm3WWFe/HPLJnxSnIw8tcXJ6pVDkIFe9ECuqV/st1H3B8nT+3ZdChkXOyit
qBJuEaJFSdLyfADo+YJPGEjXdr/ciIKYhJaIm5foeAiPwNDAYjfxP3MNYe8HWw9c
CUgfgH1IRBp7nApKcPuN4PCnrbl8UamiTXQ5ATkLc2yHSS90lScjVS/OD8CvVM58
MlKZb3+CFm2xLof7h50JOkEyOTKmeyvYbEsRohS4sml8JGO0wjxG04pFY9SiwJcp
Ky/A5ikBN/LJ8/7Ua2cmbMU+xNXOouiANgCY3+SzYrxXDDkjIDVkltTt1OyYNutD
+zKok/B5Y3gIfLVhTNLW1dO/GX7px0i/B7fxDEXHDkzEKIkmnkKCyIm9SUnVifjs
qEdibFkdy89OKsqaOJJb0kVFfPS0oCN78q/Wr/86N3MPT3GZ2uzQQ9nLMiWbKME1
FH1bYnk6EAXjhjLzpbcAu4gxvAxCjRMuBWDiX7j+UKsSLZEkmqmCZl/aJ244D1I/
jIqglt8K6WcNaGQWrPY14C6VijROzn0dtCh/GfZ21ZnBsVID7353ADa+p8RBC8WZ
fOaxc2myKO+InZ08hUO7QUvddQWuhtnoptVZV0d7uuzmfjcfj3AhtS8LsFDMgEP+
pkgS7oR+d8ae/K9imFLVx1Peh4qiaEccUutM09rqYwjzOgZOtNLeTEOkahGW2mQi
pvGObe1cd1vND0wNDI4At8od5xPnWXSZ1Jp85tgLfZiH0+HZciGcSpLu9v4nPxEg
oe99MuvfrooOArfo4xGHMILjmuXEEJPfQtdEmYivBxox7xOhC/y7sYFUmqpALlNu
SwcsoGkpGwlEKvUTwaothbBpSoYNjF+XC/X2m/0jImCFoAFilngs0k4Lfoj8/MP3
jcTWayfKhA9/uRyJQREy7jnn7KALD32PreC0c0mzc1yS98NNsMvpJHc4+XeqAOpe
0fmCQyyHIu3NiZGFy4c98ShhxdeDKQqNR0aKco7bJnwWDTcvd/F8K4Gm4LtXLEMZ
dph/lSo9volTpvikfnN7zGWLOl00sSwQPSn99Oq0qIFsNbVVKsn4/wFWHz2kANGH
n5xvjBYDH2nxPkGUKaWH3yXUmUYojeX8Ntfh+EN0VopkgfdsO+K1V0sq/IsWV/du
OOjgdHKiRff2iUh4wnYJKYHKxNNNs/AxjXls3h3f/fhaLtdKewcu5cxYU9DRjdva
OGCUQlPSAQTEXlByKi0deVD8wfH1WBM8lsWpOTwdkLp1hIJ4jL7p7actAZKnxoH6
L7CHVs2PMDad4s6esD9qXrrqekcKqopwwTUxWJuqH89UXKeofdnPWi1I7FhKZWIm
jeKEjeIqfMRnv3V/MSSeC3J9N7H99mDkUF25O646ydk96Ui516cPHiITAQ6ECCuR
2frBTWlr1F3WBqURq/x8uMzX5K8xVqkF7Hj6bAkiUgUu0PW5kRlh8Se+uFnuIDBT
RS4KiPGM4x7E79m7ILK1JtQkn4nlDGOquktRq+KT7sBzeMfvfwvB0lAXtDqcnOth
mTmqE6cBKIxoh0adn+YEaWihvq9DtcSp8S7230dn37PbvN3lNh3B6PMlaCrrlRMM
Tw6QwrA324PQPeXOFJfg8vWa3bKq23Bc0sizcRktD6KFeNLmhLlMD91VCGxmfgl0
iUm8V1ZIxUpCGTwb9RvZe+aqSN0iBszYR3ouEOZaNbrGUbiCdYqXcXdvQkh883RR
w6+mvkmuO9G3YUMSaWXhjwi3YApiS64CEDRJYhg/QcYBgPgM4TqU5tkMML+9Z0iN
dcTgiJniNRpPkCTFyqN3EbrAyoYFk4OFXh2vKGSMVfNlbjwM4ny1X5ImRcYS32vD
nDVQL6usGPQf+Sq0U6J8+hyPj1i9WMtiRpJ4tslp6FFO2tvbFwp30LYmkzEiJIe/
6mZMH/iWBczdQVnPpQqfJQNXzPBW6GEb2TpsDqb2NER/40/01PCaMHd+gkYtAW6Q
8Rc2YL4q14Gi5ZfZKSbMH87omZC2loCSadxOIv7PFYBRmSovnbBqdWc2v6/usgTR
7zdViWAQzXHg976ETX8y7HjjwW3TcCoRicAfxC5W7KjuNctlQkIyG9CbsIWkAgcL
g9euPlMwGkgCxVBNKwQO3rlJ1sBhJCmSuGMz0dEHo5gx0zyLBldN3ASUwJCUtG/g
Q2/fGqFF9i9WMtTbcVYb3deJJNAI3FASekNCKDC1n3B2g4F213FEci3L6bW9947W
16AMicurI0xSKt044scIB3CFopjB1ROK7Wvo6kuasaBdN2BNR646eeXbVlBE+yuZ
Bj5xTysMv0NoGiHlkbYiDYglcqozRvSUUFMjPXI4e/vwozhfEHbI9BvnZKRemYAf
XQSQZgpsWbR9uR82trDZw/HGIP0Jq0AffRwzomQJ+RUmPfxgWb4Ku1MdsKLVKDeC
pDhy9Jo+iagfE/iCIIM9GXkMO+qmAvGLaoIlOq2V2l3NyQsHXSakrK1nKtDd6uzX
xDb4+TqYK1kjcINDhUhDRx3Nk3uNUvZ/+LIMZSg4wJ4SMTS49QK5syMfV/LlOpw3
hjZ1GLOwrn6f1+evJTEgEPKq0s1gR3AFP9FcVxHkqU6mPH3PSlXsQURMIzrNSaMT
KXl+64SMv4wrgDuBp/TJnJQ6VxI3AbDSm2nJf6dxY/4H0a2ZA00qtzNkcCRag3G/
mCfddGZ/kNnaoqopiy5dfVtAhpUvJKVEBWkuHk5dFCVaYYgOikhZhLJF5b7bVF64
04GCYNRY9uCxNDmkKGPhjJONbIDBa32lyUUZweUxNunK5e98p99zRGpbGsmhjUaD
EITybdu57VkJQoEiAVsccdsnJMGqwrIb753A5I/ve8y7WaFhMjaoiDXgdPKTVVRi
iZYFAUrFYCtAUnSibfsNS9Kkoliub6n9MYeug2+g3WoHzODSkBvGB4J3IvcoSEON
1mGWyE9qjSGggutDRc7ldmWHUqEbyjtmO2WLehaR9maON+7zPCLT/tjyimKiuTIl
+cKq2DKYFtTgM/REyIQDyfyAQHruxt+pHsi1shD9WdVAkWVPqxAkkhn3mYeex8VL
Todh6HWTGH8p2uj5jRYq7fGc1VDVYNKddKobapXQZK8xcb0f2s7OPLEpuwDRIr3D
JjxmOdZMuLO0YqGhNavGW7vmUNI3u7jaSi2pDBYsuq06ErDEgf7rspVS0AYhSFeT
pfeSuD+9eX7VrFGQnYSQxTPlO5UeF48Fz3HjjHtFe+I3XLHrf3N1N26JO5dYHrG8
ms8KbVdlgMbcdOKhg8NJOaPqSd3i6FfOoOvE0+x4okkbImJozRM+6kIwAviNC8CT
KgJzggL8atEYIRZBQVlCP0YCk9QUUHrG9fchU4fBuRXcco9I8WczYB1PazzBX89n
FlMLNJlmCmjIB/QFrnO6hLNnGU7skh3270SWG07dukBkY2Qd1DC+h5RS43NrMv1Z
2qpG9Jbts+vQQVbejPwqnQ8mjquwhF2Gn9STZjcSELmqdNaVq8LarIcd/6bO0Jhw
PuTGJJdKC8IRrS7oz5881GFl1/2V72gQT7L+/v9H9ZLk1Hz0j0FR40n+YNeH0p9k
GqNJMIQ5rhf67Kw4iD3TNG+sj+T46E9ELt3BjqFU1/ukTOBCKfvRAU2C06IoxcRy
+EoCDQDjrdIdT83B6/R01E8vBb0IMyFjhms0GyyBmUYJVV6NcSwxvHjgDoULVrGQ
u07wvpEkaL/xii4Nv64mW9EcLNCH4lWzrft/bGeRjnEbSYjgZ6ldJ2JaMSo0GYg4
/V3fkKTwMFE1MogjrXxMK1GhfFqCZ1jofF/XkiRAPlYcAujgl9k97u/XZEzUq92y
dxpf7CUEp+kJ9ohuZaT+gndb9cBu+awNvlF6tTm/iEyCcr0QwDswNM1hrcHpW3+p
COfY9uSeQeDqgKEvjzYFyBR0GbyRFU+Ap6TPZoQlyjgoouJE/25nTfQt9+OBKPIQ
YpS29xE7StyHgrlhZvf9z2F6pzvbQ4u1xhY1PZKcz9quP1+Xk7a69AtciYrm5/no
0AectBRO4UKzQY0oqka9dOGQwOg2Bfo0kwDfsUI4BBZYuPnHIHKhDNIKoKGukjzy
RYudPPi2ufrrxJspKv9eZZX6VgxOP6bOraYRDLNFRi3gN6OPjA/VYzrPL6hoS14P
/ESariDJ29UIcNfwDynokYdNr2X03fPv04a2sg0VWKQYuC1rJ2u4t+inqqn5eqDZ
buAvPMloGDK2s8vCKsqz1JPbixeHFnHL/jA+/uBLsS03gqIBfYoirkPUJuQynn3F
oZgKzuUFzVUclnFGcGiTp619ow/EKYbuh5UBmyKbYibkvThCXBtqNR8BftJqqr0+
sgmeairTE6D/iBCWP91K2zgoyL0z2SBJMHQveyeiXJGSEdFmtwddx08KHZfseZ5x
cZhDXcchumae1BqJwqcVB+7/FA0hWSXF0LIucP69AuZMaNycgrYwHxNtFsQ4/F1b
uJrPWMnk1NJ7qG8upQ742axSnKGCQ+cxm09kSM/3EhGMZJuDeDVQhsmGLfebYe8w
kpXdOusem37Ntm5NJpaw7uCJrClWJ34J8O1m2fJRLOYEUODrxf/+tBb94iAR4g1y
QaABHMiaoodThjFgUVecqgu04eWBBXBu9VPdgzxZoXsbUplznEsxnQuWxN0sDlQ7
FhvsBMnsuvESYoSvGUGOR7rvDF6sI+xjRRcvsqu59U8hdh8IQsWZEDCHQ2+DNSNN
+S6IKF91FigwH/j8ndXkpHHetjOuI60TsfrIktZsf8RTDLinMAH9SnYSx2MxNv6I
jd4tHL5L/raT/kRE0LI87xzllK9qWdpcKaxi0/lfLgFtGQHQ2EDITn0FBSojs+Kc
itY5S+cf9SZjqZcfunW5dyceI26jMcOexNACqykeCf2IZmHGORHwkwkt9oxyjj+m
T9jiY/Xzk4hnDpE8GYvb8AFSJNBKouAksBakM5d0JTmVdPFh03cSrjZrMjb6ABdd
AI3uAZi7NdbpCYQ14DuH9o0bNnePRdUpjabHHEyvjfDEwhtJdKbJHL2AfNdwXHKR
TvPwAFeJRLyOqStWgmQc28aJe/cXK7+rBIkAmLSsL4cWRCBpvgqtpHnPKxlfxmxh
Yt6R/gAXH/YqnbymTVa5KM+ccptfsnIPPfnG5jjOVbkdAEyxp4cq4QhIyX8nM8t0
P6mpRiu1lN0+dxkh8j/0VIAZHRXI97VEvlHr313kBAPcqkFqUKvfsyq5bzS+90yN
ieZIAw0q+ZAvDTgyV/9fSonhCdX5CZt8cLEvjY7yNCjjRpVtRONqkcH3TpzXfCcq
vxvpBr0wmt4eZQl0ONCR7/m+S/+Si4Cx/JV9oAOH/EPHtxhQg517/OZ/8XSC4JzH
eU88sNW8z1x0uD4ISy/2GUCCPe4YD2LOkZ0DT9a7wFTkvVmn6Iu6kMM85OXVNbTv
WUX46jkpFq1TBCaGRckfbtqhl1EeZONi5hH12oSwoSH4Xa1bHi+abugb2ahML3VP
FQ6LYyBFEl+HXvDjF0Waz7qM3cvKZvx1f5ElFsGjP2GPQ4sZEyqbgThaiIFpkHm7
3yw2JGzC2b53zBT/uzmPRuVG4k9Z5VuD9m4dg4PlW0qO3Y0Uh18dxQ0t9r+7N99S
Ss1iO7FsWwXBisSrSzZUP94LEglRgN0hKEioQECaFsxfbfHxPR2Z51DTJUnH+3DE
YQxbqZIfjrRBQ/BFlhxrPGLCXmwiYy8TwEgNTNV9tXpiZQVVncouyNx1jenk3S0M
INxU/ViKT0zQU6hhsnk7oA8aYZWn603kqbipyvTDrstIsemyMBWV6VZH00D2pTgo
pyw0e4LRlgQVM67VymBpXUJOz8dN0byOV/JWgmbyXvedgjO/PT0GX5yqn7L8Mmvf
lTVnO1DxArXUl+s5+bKFXy4MI5T2BAs52RfIxVlVpeHWWUGwL3JfMY5a/Gi8Bg+Z
ZDVLi0aqT8uDzCGW71GC/uyfmjTN28pzF6Tl5hdZFgHzFBdOSoscdGzBiXTKZBP2
xWTiGrsm87hlzwbbtaHoUXTKRILC4vj/SkoXOnlaQUGpo8hgGvEhDmqVAA/WqJo4
yE/OxQCTZPiK/vV+QrUOUZUZtxq0w+UCTbDaU6sVjI6LLEHkWegvLBCEFt1v7pvP
zyJRbrVVCj2EFyKQhBqrGSDvU9V2NJ6Mrk9zUCaqfhBgBoWA67HP63/IKGugYQfB
A12IlYmtdxyK7ZYVusSerELo8GxQ5ZKR4qqs2Q39Ul8uWwKAYvladB1+aiJd7ou4
ARsEcwnPQn0LKHIqUUjHY4xgvYm2B++UHayEByvZ7U8I85BFHjLsebVrN9W6cqF+
sttdXiihsviHMcCONlmph8ux4vjtEqy0rMHi39plzJeHTDFozf1U0kwPd8pf0Elj
ZxV5AMAAMXUIcMdQueZsNZnu8E+Nsgc4nL7vr2YtMtiEYhdxPuab1KaJ0vUFTsvH
RDeXe8+NGJo2Be/cpMHMd7Zhmf+Ms9aQLYFF4KODXr6jJi2ygJs5I3ZJib6WFp/v
8Gzf2JFsxiynvzYmj8lWIMMs1y8BPcDZE1qRfotX4PwgyNEBkLmMfUG1mWjdGGPM
rixc+QlyBC17vzfx2uZkZJ5pLRitkIuiQXx/MH0Nt00OWmii4IPISZwKrYq4PFQ5
AjwV8GsMS8ywEzd70zb9wpWA4Wm+IbSrACfagF+1sU8=
`protect END_PROTECTED
