`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GfwZeYQR90N0+vibHXGHwDQ1xdLtpJtoOKjyhR/uDqNrAwL+R3bK0MnKpW9+UWny
NnuPBRXuriHCI9EhCtvlxg1pVIprZtsqYFiK9Woh0xz8himESi9CsCsg/F7aYY8L
2mf/6Ido7AZeQbvxiEWuRNiEm5zpJboTmC6gdnEZbeGtpRc3jf0Gj+0XzKcRgsCy
JU+CxL4e52vNVpOoQBiGWFksJhQ7XEnvt97PkXGchY2J4qPzkGibGj7j5Kz+INAo
dYnd6Pl7InX0T/3WjxfAvtQ/F7lD0S+NWQpagYnymOVZe41Q35eY1bGz1wVaIUFt
mPeF3WIQhHfDBhtNlKC/MDA5PqzNbVQAi4I2RWS+2Wq507g49ijr5JbwPckUdGDS
XDWm9hkkNxPF9AtWZvn8s2Okg27cPOrBWq8Jnboww86h4bq/Y8q/lWoyG8h6fOcR
Muu4glbmpf2+WVETnIoKCtROWw6weSyN5tjpr/hfqU+WYwCCM6axClhX8WCo1o25
rNxuUjBaTQpKW0PhUZpQ9GiXNs46s9uO557Q5Us80g1Hj/UstNMuOsa50TytrsNB
i2z+hyV9nbaqpi5FPiep4MZ8N0CVOdX4kmnGtTgTtQ0ZcDIl4yASnAIQp2U/v3Ea
EwaHbycQIYpdyIH5LPKA7HHePxK5fWyZ07w1LHmksEeG7kIz0tjDzQV8Zrw36l8x
+R11BbtDaHDOS+SFc+cbKNQSOuJTTWLrp4qBHrTtp9jlyZNP2twJpFuBX2BirbT+
M50roOFJCixovgGoC4s6VDl6dZ2iPj3atibqmaq6QKtnK5ZO7guQFhpa+Drf2dgZ
XyE012IlQlye5Jce2X23RZrG26q5hDcDobcMPrSpkBcW8EiTJ8FbA8dAMgjGVPIL
3Hov/Dgk2z68sZ6dcCRQSBEZbY0uZwJVDU1g1+G8amiyvk73JjLNOu8wouO1ji6+
xHAj1OOLLRh0KwGsruB/IqN5PVPMvRkaeAc49bJCEDHwsfPC+A/IblqacpmIFZbe
/ikSWauZ3BnaIouDCvzpi2BCwsXTD26P66LXtS+qb0Fq9fd2Y0f7hPq4I8LjYBgR
geJBsYxBxkGtUdIdtqu+spPrVjZzXyd0dN1cndWAj6qpvmEC/5xKhS+5ghskbfZr
bS0usHaFlqhh7v2Mq83W8+EZxvtpLx545uupPT4ATnQ1d6LfrAJ7h/nAzepdqWc8
kDRvzAAzbp7coiSIxmmCcbpkUCq/uUIFGRGGo1bWVSvqc+zIUI7m2MQuG3lhBuwJ
azYmrA/SciurLqFYlMTTcB67n9c+yKKmh3uJWnszOXmCO4ZNc4YXKmG5iiyi3znU
O2BlP3oaFvHATzffOBo3VNXBaBRVzKwJZbiNgi9njiLsTuvFT7AIVCLz/Y6nHQkh
sfT9HyZKfVI+BW8NjA4rbIfNOwkUszz9MHbGLlpxPUy2wkEzbhLmse/0eArxZSKS
fb47tROg7nVB1Lexa3jx5wTqMMlWH31/rKr3VuNQU+pCRID1AdtC3yadOzKqEPop
spTOto+gMTKmNGnEGystz4qcpolYIhYXk2oFjyFneSSrMSF5t31SQtlykVn1JwFr
fN0eyp8XcOxQ4h7p57ua6ptGqUrg5VB28MpvIh6Qbj9qaZOYozDSFG44qsx8vaor
mBcONr4rT7AzELeh5hTmZLJcd4hDiOeA7Q5sZ/EpAU2TvthZscgem0MpPAC9ayjB
zG3bhjC2/6jVz68cnRhqtHwi+GwO4g3tnCTz0NvSkfODJn8OGIn6JdEdXIy2OO19
//6gZ8tNtyOpLORhcn1w+dK+zctGyIJ/lO0p5WhXJf2FWdYL6q19++I4UV8sfo8Q
rvePswWWZcLzm3F86mFi300/PXpcNal5Pwmw+q78T9uis6DK0S8/OMHYem9/j2vy
TYFpWzJTyhG7PByTef7E3g==
`protect END_PROTECTED
