`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvaYVnaybj8T6wXyVvpNHmVbOP3onFtTD6WwHxPY+2OViURapAyBj8P+l6AuL/CL
iGlpF+2OxC7e6C92SLRnDAdzZUB+vhMKJaA3ttMifP00znJMQELgAe72fXCsMNtm
lJAb3smsmpF4cwbyisiPrwLTuyrAysCAXpPyH34pOuHVaBSQptP4PHqlswkHzaJF
SS/l4TuIYbTOeU4g5TmACQmnbUxoK4sxpceI34oKVu1+IHmOsmbf/S03Tq26qULH
Y089P5f2WgHnH7we09AbhoyjcVFvvi5C6YZVPgs/e63lv/cj/hARKWOiqMGUqJU3
b6X0tsyATDeJTchixN0wV8R2LUavzGqZip83s0Q9rufps//kllYv2NUIJf5vXysU
sI7bfOvBxQgWumPY5LvCN1IpxQdz8/tRGbjh2rEWL0BauoV0vqsuL8/kk0ZwOQ+5
G7Xsbw/oknWegJlpBKyXHdTG+ei+WP+Qfl98JDKZJlrrZiM855Va/KMwNNp8MsSV
0A2YxirYbirXuakSWo163aLU9+0c72VwnkFXgg9vu+5JAirTd30CKBKEsxyknMWU
BHDixEJ15NaWZvvoBnd+HZNvU41R679ipWnfuCNLMoHmRUIi7p4Muwl9OCYFej1T
Srt6k39cx+S+9TUzpaWJLPQSR6NpLOMsZ8VmNN/Ela0aHmde+pfmbLS5qXsBHxEy
kXlmw8Yi8s48szFROIld1mATEPqLdHBH2Oh5rNjHQvoXMthH5rKzM5MwrwOeNPGv
7t+Zh6h5a3k9UKmhKKp5j32NC21Dg8vqTb6sWc5rzRPVbUz53gloj6ydq/lIrlsJ
V4gZKbU7l+BPdswfPHDEm3lw3f/BV0DfEZsvL4c66MjjDPAe7GjuxUUnScVPiUg/
KlyqNYyy9T00U0A+u6f89f3jWsNhBuu77k5iNPaNMAjVMYNVTkrgWmTR8QZEah67
tbcrs4Wml0y/Wax3XaxbhAWHuULopoKihXqpPIwv5E9cah0bAJuJfZCXJjyh75Nq
6k/BjOpMCOrNrVDK9pMHHVGGXWxvQ2Kj5IRJ2mRsWzYgzWi5jJhHoG7y8h/cOotF
br7dlWo0Ci++PTPsjEXkW0dbmk5LHaF/68nb3eTrB86NYKmDbi95U/icIAoy+DzC
Pq1PnAkAAJ4GXwbWhUDVfgjUqrQHwOr28t5+4xYpItttpo+5myPjIn86QIgHQf/q
imU2m+IZ8CfgGeRXeuhi2mt9cDutEbLg67IbQbCeM/peaQ0rSVx24EI1wdC+gOKN
SkkfT7hVUBS3vv3Dc45rMMQdd6Ogf2wZY5eTOIsURcg1mcON9+PuSuOcWoBQ/URs
`protect END_PROTECTED
