`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t8T6SXlvoUuoVC/nqqJL0QSH/uh6pbEefvB8JzAlaJXAyJgcgLt1dGFI2RdNUY3c
0BRFeJgvAueO2JuvSOvnSNBsIgIXPziq6e/O3YgoLb64HBAado6/h71gjbr/XruS
EUMh8TEIqJTa7v46W9XC2AUR6K875Fhy25HKYXRCMuAtrqmkEwux0RnZJj5kjZ1y
keaRTs2gAcdOBK2jl6j8DppkaUN2g/W7MQFjNArN5U4kxTMsqM7dxrMjiUphUCFQ
78hXS9OZ8/k6PrWdW4Ea4M50y4dPoXlnWtwQEmyDHC5cuxz38ZIkKvW8hMwKRKS+
D10ecltFehD6axEw09jNwzkSbaeH34YDSAAJj69yD12TwtEl/185siMm+SxDnkOO
eyyhw0dM+AdqxcOOn1q52zURLvY6NpD3X6wqm3HjOEv20YP+bHEX+9kvYkwtL+8A
yiHl7WONpmrVP5OshGwXKSBljcmtIGZHtFt5GTeLaVCCXoAWsmvvXz/Jb94Mvab+
BttjjSFiNthcIuS8Xg0zqY+d5OST1Hh5ziyQYuG779Bxq5pbdTu96Pq5X5fCj83M
MLNd6uV2wCANJxpGwBJcmE240LdQvIAiUnAi3MYVGRbJaeK7A4TtGWLIO/TWIomW
eNfsMI+Kz3yvFK9sVCdvRkJ5tfRmT16WIQPIO4JV2lTct1d8QSu5vfHexq1geWWL
aSsMVEw39flqWMagn6kPGtGC1CKPq6KrRQSYsO/xJewcyT9iU2BP4bk2FUdHYyxP
huLobXVXyP6otfVXLKHxAAQUVNyWn/U2ruZf2A1RxN9Z6spuwBuGpk/hlSN2KS6T
g8SzWAD86oyjHpMOqYFhi0RBNclOkX3c9yqGIVVttu5NoU5eGtIPrGcX7tmF8zKl
CL8ZdcTriHjbaPnRhidwWSgAZZwFVGyspuI7qGcO9It1J5L2ElVKfoaB5ZwzkhFG
IctYGjWZlzpuwjEQMfqJc2i3pRadYeRdc4NSlkC2TTe7fA96/3o7Qw6peo8/MhCO
kOwY7JR6S2NuJbUptp9jgsuadp7xPAsErMhkHyRC29Mh38TzrNj/yMCFQkHVmqO0
UThgPac2+/67eHedcI5MVpYVEXBfJGVu7eW7HSJ8GqCH9E19SlTEvgnS7EzRsEmp
IOFaVug2TMQXo94guY/TutsFDSrgJ3mktty8A0AQ23g+vFIZN3e5ouAfy62hOU0S
Wj79NR3KoEZ6Ol/8LOQvcOkRf+YLt+RecAbg4NunfJsHrbS4ZYqAJuBZigcwmaOw
8OwteuHq+TIpP1ZU4REFWpPtQh7q4QJiLDM5mTqbuuUKCA7TgKysnO5EYpAyWMNn
TxJM3xzt+3V545nPfou/kMcIENuSDw4vQ10iZqPBkJPCU9H0HgvLoXneiDjbcAm8
Tsai6Vd7szNKZcfe6N9htZnLdpBmGW1eKde03Iz0zl7PGxWVZxnrnA0LnEmk/Wyc
hN9fYfz1YXy7P/tmRFjQ1msGOC/84eBzIgg4509V0BWs/FycTS+EXeZub7PRQX6Z
A/kmKpQZtag6fknEYg/hVTkoPtRdurf9yD3d5juY1dU6QDadQPJjz1gT2Ha5sgou
DOCWirNmC3QplcsrRD5O/MRBQ+NbpYEVV6x9+92IoDEus2cNWs8SXWk7Jpp9Shqt
ubrs/Yw8Lv89Kjtfmp+ApvEcmXjuRQNAli2CerjqDfhFhhZG0DF6p4Dd3yx95xb8
ad2gs0YmDxOyxvlJ8FdUGyGa2jWwiCH5Tie/QgG9nobMspEWFhK+0WLKdk9HrXu1
daTU4+k//gby4aFW29XPRh05eST9wzjLrwYFaHZ/Fu7jSwhv1Zjf4BOx5a9modYF
0m7sz7hRxop19/l+jVMDBt+BJfgLxgVlSQIyRVu6+bOlHdcGBn8XZmPN6wCo7Q9E
X/NYbEPNuBb/bQfArWON+HCUwXSlORI/BQTSO4eUbbvqItWH5+ZXHGXTS1Vr+dWe
ouWHEk1fQhjnYDtDA2VB2jZxO88HPe2kmEVM4UiWcu2HR3xChJzCJLUWkhPvFjw3
3JGtT/6/+cdgcW5wraNV186OREQC87QCyxcF8nZ4C25dpGmSdQuQA6W+xstStY9h
hOX+jom8yP4C7BzmpSieWMFqRsI90512FFFHnpGtXhf9b17lAst3c1chKOZ3WmSL
kAFIaRyNiD/P/R1pi1yPtEdHiV80ivJT1gmhow1EuQoAcxQxET8GNbMrRFKyplWW
iHZcgFUXkeDX708Kh5+aARsy2qZFucdl8O6em8h2yIPRCewhze6og8sS3MUctj5H
lA8VqsM8IPg55FTyWN1R5VE+k650TRPqyl3fKM6GHcaVKFzsXQKTFzv8P0Oi4Nib
YIfgO7BkQQ8K1bAnAeynQnNa9/wErfqUWLvGn2c/07BBE8hfS4Wee0K1nRrpr60k
TaKmC72Ae0ZbeV90JsVaLRRuR9z0SFKRrBpDq/j3g/XMPH6N/xPNUL52kMCzdcq4
4FUVFEUhqSoV7UdhEsxGJMhxZnVngGSyS7REAMqdGRgeOeRGq0f5I5PL5qfKmLzI
NwPKCP3Cho3hn97KLcku7jnfqbEQnJtRzSGS/8kuK9NG0fgQIXQs5K7iJumIDnFh
SRvJErHz3gowOZ64xci8x9ABE7JBmbKH6nyrSTk7OjwgY/GieaIyAjEBVHXysvxQ
iUKADXK6X0LW5rpKjCDrvxEHvU8nsp/aKOVhbd/8t0rzRvVzKKRv7vfpdujPrGEI
s4h+5uGrkYm+PS6EDQJi+DPrvzL1oeQEHhqItvdcIP4MbK2ThDDSW0RnFn1WBOAv
ns0189LiSQoueZIq6Mi2pI6gHzqsO10pt8zIHema2gf8YKj4aaS7/Y3Al0Zg/e8J
5HXWHem5npdHILq16Xa7lg==
`protect END_PROTECTED
