`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQDWkBmk9i5Ldf5A2JBJGiOybaawirCXc6SbHGlwmm7ibTFkPK5ZaaCYigCLWpkI
m5CokM8gxE5qUNEfXjB0vGZqWGyAdHbjFFckLTKobuEyl9I+kUAdDfi4+UBcYmyQ
Ps5RJ1d36krTVFjEYKTRtwhEmVFCQ/QDLdiqrY1CS4M28H1a7NpWLJtjodcm6Lqo
CkaXHZN6pAzxB/n1UdqCc/iKBKbR0XYwUPqpG/pIPuQx5Dm22aybdLv8pYEY4rbM
TulAK3P8zG809r+dsDmHQ5gfqe5OJFUJbhaW/1x1tg+mmwt8QXODcAb/GdUbCL5t
m0+M2woudlLdKexXcYJ0PxpZ9l2UIbtWpMQfk5qYU33k9NJ+euBdiGraN+7aBii5
sm5sZAVxN18j01cKYYKVIbF3ajtB5XcMFkCLrVgDUN6nTiYE7pDvUcrsgZMPAtfI
ka61qW/xjeRNnUx7zLxorNyOfm5IDWo9F3cS7xcX+sk2RKIqmlei6MpHaP4L+6as
+SH7M17LdoABZI55EjOEvGxYqoljPL6ABWogk09KlVWf3zyF7wUlUwL+4Bameaf6
f7z33KHxB6G328a5wrdUQRU03Bnyu8DLaCYAWkh0TdK4eGpT2s3uwMncQNvJKcqc
UmmGdAXfRX+iriAPo5km7p1llGzKc5FLzhCPy/+46+Gcsc5NCCm6WYw3exjE2BSM
NIkeOA90YVnJB3+6pLmKCbnCUH84AC0wM7P5sMqumfjG97G0XtGProoXAypmTP7/
OKCHjfLibXt/+5uiAbMuhi0sGbsjLKv3b063B5VJKijI+JuOg0urqvE/AWnvKT6y
XkgGI7G8r04BooRzto+32hVfBBchcI+fFUbv1gAX7GqYCTvsqFSrSmTMDOMmzJfk
DjfX48NpuIG8QnPUQ1s2iVzvVBiyRYFSg0gqM1+zDIvrMM0gZJpe1D8CaKVD9CFN
kSHcV03jXJY0pglJ/cAmDiqzO71JFqcnTNI4TsiJFwX0RiOiwL8aYxJZLhD+9jn9
y5n0378RLT/W2wzpiupxZfms6XUG3cX+4Qcj7Cq2QChqoSGjy/rohjkg/vKJ8KqQ
bm3VF0dPSE8NYWHBQ358Sl9xmmtXE/SGGYR4CfO0XqzvI3sxTh0UeLUIUbiWbAd4
bqnFIWHkwqDy4avfq+dnK/iLUkRwiI+k/swfZACE+Qc964S2a/T7vBML+3FE5VhW
jlHvZJaB/0UH9/otBmQJK3ZiGvSOgnVgwr8U7mDIssKPR6OGTtKcopcsVM9XfbqM
/mbMAWqs8XwYkP1Oi1kgqZ06Si4ZqlVhSjFJCSpugUsO9m9CpGNfBSatzjcbvV1h
Nb9Zhwj7/zcXk/mIJLf+pLVijJNPXN0mFR63hh3cmg7WM/Ai1B+BwZP1PxG/mOrV
1rBfxEfqkZecY83qzbdvmoQ6xq529C6Fu/PphQ+rxf8cUI6OLXg9XoAIg4bfO6yI
3I0rL7wJbnzRMiRE1KmIi7evr09x2LVXU4o+8/7+O/u41Ycw4vPgw0GaExeTCFxJ
0sPFk3A/NMYsDaqBQuAt3rbEkpTCX/LmxOBGA7Xzt2zl51Ngn43SkYPLKwtPANf3
2FxaeyWRzMeWNZRyYow9PgcHNq+dh3MS9sZuSCiWe5upkPR+oS0GN8I93WqBsZJm
E9LaZNCMhW+H67eBlOQYmDtqNbcfHkB3FabPsaHP+GNc9mIAawgA8uiql2cwmtoI
GvhUOAa3dFLrm2QtRy59dLq579n8/NUoKm5blr/1jTftxHgKsgHX2y0UjJxZy6ku
iMVGqH45mQnFpuWQGRRDyGHM71IO2rF8mZ+6e2c/tKgF7Nv2pR9WmlxNmXz7ajRb
HcXD5Ta8+ew4XMPhJjULYRdodwvWzG6sEwYe20/eZFWsdYyrdgnWuh9Bcv42SPvE
CqqmKrT8aZgsiukmhVnsKRoUQLkSn0YnLF99ZTc5UIGKv/9RwYrnj91SWRdEhUtN
yv5d9mzu8+AYcwYURNAzfDqoMMTe74LnlVSSbdugyWBaHxMXGWtPewowq/H1XcoN
/Sn/XHRHaNuVVoz8NvHa5VZHHNjebcF0BeJpBIfJ97H9V5nU/Ji//x81Kq5CpnKZ
6SOykgF/hUx2mwjb5gDtBkNxwZEW9DhHL1P75p4TF/3LvP+mZw8dl0zHGuqtk7CR
HCLo6BlAwNWqRjCYcP3Aq0Hzg+RwBhjdz7p0QWK9CwLbAllRttb0tivGJ+S9TL9h
yloo4MGDCA2dBObvtsyAzrbxrDR2ivHTH5pNzVFgJ+nSaVIw1Nv2vcEdGIESuEXS
8/hvqENErTPNK6EGJR0uUIhejEd+ZGm+Tzg1uvgAzasUykACCfxU+JhHJIVETNlU
+8WAUqQis5lpHw0M6g8UX/I3LaQ10Wu6Q5JzcnXUFfIQPdHi00cZFzPchm8i7slx
RDcPLmaEBzxOHXaFKG5h6f/pxTh0LZZkmtr2KJ/TYUgNqyeZNnme58Aiw1jxQXbf
5nkgFZ9V7K96LImwV6L0Q1ndnpbIXOw94O7IC2P5nNgaxw2LjRIw7WULvB0rCxnA
AG3CRW0eTj7yc4Bx7uTVmAI8BDyI5vxaOZIO7YSsUQvk0tpuFBh9tieYEw12n6ZO
H5NmJaOtKORjlrE20p285i8wsWoYrcxpFq3lNsvFDLYn8717TfbJVZFmyLZTJcMw
gdJ43V8mN9Cmj2zrwsZLk76VRHd9OGxv9M0IFx99bfhsV8sYZVT6osIew+KqUgLT
LQ38f8efqMowSn32cN0YkuQCET+aGwKav5lKhoo4+UB7lWAJ6cOh3Pa8usFpUjep
3FBUIXmJOxn0Gb6jYVMFSB5cQYDcR5+1I9Q8RpPKMvq+dwnNzou5D9Qyz7BNwnLK
GemAKBzfw56mKnjrkRWVkuNH5jsdxeA6WXY4hRTq/GkPIRyS9vhw599UvqXxXggT
gm09RhiOEne8p3PK4lg2MAaNJi26R9JGFsYkI0d4Owg=
`protect END_PROTECTED
