`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sffsvPyoO2DH40m46/h0Y1aggTLSdUcMQfyGNIeMlXdIkuENzrTCBoBMmdpIq056
nkXUgNZ+AjkJFp4UwM3LjvVDfPoW79zNKmO/Zg7hrlpF1L1l0uvfpLw9w3cmAE+Y
Q3eIFIAs+kPdB/vXHw5q0jLdRFqk3OeOqSaOZAMolmPHCr3LyP63OxfhH5hJXXvA
ZKEu8m6QTh5yHOTUmduo896fIaKRUnDVJtVAl9wFrgk5XaCErDEycrP9GRMfuBaF
NCer6gfj5lhTq9PFuiPmKJqvhmsdX5Wgqe2TE3NT//guwWkXF4Mii7xyZKtV/pvY
ksWwYgba4/Lxfov28VfpzFZB0bVLuDcm3kryA0T/R2tso69p9186qlbrp0RZLFYt
+R6Ovn7cRReEI3fIDDguEnYJYrfPqEdEdMhMRuDv0V5n/mtbx/ScV/SSoBgLmh7Y
0u4mbjzg+wEfg/Ix6bsfANwUNoDNs6gU9vakowI501j8z844BkGkw5HZ3p1pBJ07
wNuvC8MLRO5aRGqB/Z2dxO6UcdryziGdI7V0YNI/bFK6HEgPDGxUEQfhB5X9QyPj
ZyWIJXk+nuh5cKyxX05gdsPrCFee7E6ikS2KRjfJPaZBzlTmzTipRR0rkjix7oOF
MUp0dqN6govCbOaAiVNnmKh5y1qRE99P4QEUcSC/TtZ1/ZiZpBEt8apUwutFRc1w
z1eeQk6MhYQqezta0GhNOrhuIG+QY319iH84VCnuSP1V7RRJttIO+9JzCggQbGwj
Mu4oqxKJ+YJO17rm8WgWAWLqkjUCz0UU0P3A0CJsjOnLyUHrskycK549sI4hrKTd
a5aIoooDR1lfnw37N8MRI6Q/IWeS4Pwayyxh8IF2PD9tju8lQuTZzSdP33qPokkA
c78g618zwohtOCKZ7V3qOcarkUDk03nNk+sZ4K3hg38/XgQIl8TAsnP0yFguyZgK
RWq+Dz1RjjxgEvqtQB3is9z/p0PSpcsgOSHaxY/+A8VikMJLLQnQ3GZZv1C1ODSv
iLhGdw7Xo9GbQps12caTnBRaNNxBYJCNxrHrSEQT1VZ0kVVluVUCaaZxzfm3XsY+
Cr1/zuS/8MPOZQL9ttHv80WjEnGiTxwFQDvOF5QmwikE37+JLMXbrd63AoIrS3mR
BM1myd9ADKSXhV2u20Hx1IsIhmGVZyuGVJC3M8SS3af0uNEOMURCAwKOEkKPiYR6
Ka9FN1pJQY1UznYiqGjJqkdKEO4ZNfv4WmhiVnG4V4TFVp6dkY/I5SS59xL98UWh
FabZ62Ql5qJ+fgrw1gzt/K93TKjXSepaHb40M0Qnei+QJXxdxVaEt4hvXXaXYwzI
VQpRtOdY8lZXngwC0bt62vgKOElNgNxDXbwlHdjXLJeWbgEVP29czOIBwHwt1vxT
pkuGZhiwPJH9BCvPEbEu5WZwEVY3LyUcFWDsSYgta/Nq9e8MCGaIaJZYOP54ZsgS
nvwU2hUd0o4D90t/DTcZk6FL+kt8dIjs6+BdvSmyT/WqzwkXvpSYQBcGGNAgKQml
sHnLUuoh2dQV+V66QSBgw0S4nhAJmCyuZZr+JGOcVdgXz6M3YXGVvNQSlHnFH8Zd
3E2XhHaN0FY3o251M8kvcnJurhbPVPFOGDwo6C53sEmjX1QjfH7/Up4tnYRfsFOV
Lh+9i9cyFGboHJGB82+m7jKp825y0t/c5plODZTDMVrVy7B4ouRSlshMSk4nOCqk
0dBbwT2/JFpp7HlaE+4gTWFjfu0Rd4ATJf0dLfh+WyQs2cWfNEjVvLc1eHEtFFsZ
EfyRpuL0J11/hap2qJTmlmAGv9l6SDr/acGQDJrKpsvdIqz6dcFi3XuqX5zHw02/
rgg79Yefitm+E2PHiSNNpatvG1O2aPNHXjhmX6nRXVlWsEQBFuQ+6og/5Ndf3I6C
OnW2CLsa/IEcjDwm1F36d2Y8GWdy4fXOTeCfWyTyTeZtHLaGCfZXj3mn9a80yPpH
6Uql0LCF2hm7sCu6GDG3Q6c6IbWSu/VCMKMkBrJ86iVOKHlzWjI2r0H2grtlzkqr
UrBmFZOp8t4qiKW4nnzmsxf/qcsdckb1/J4mufHK5NhvhS7zXU8+7C0t9lHDKNMD
rbHn0Ys3PKkPV1gBuGeCNckJwqscFuo/vVxNSycwF57PBnx4+9BEJ3q+eJYc/9gb
PGEqdSUZQl1A46VA8NCe33Lhc80wfSS4CsDmKEO2koPfy3mqlPDZKQuO+9vAhq+E
`protect END_PROTECTED
