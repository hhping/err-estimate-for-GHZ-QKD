`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BkRsxXvAeR/io4O5wGE+HhZ7wIPALnjv0kkpMFez35gdaGwEsrZJIpD1b0u3bxr
pk5tRX6UIuDIY8b4J3gd4QTSE1+5obpfizJ7FY+pOYSg14M1EUM+pFfLypQJxO5D
07FhlZw/00N3dlP84G9MxBcp5lWIz7gqqbJQEp6JjQWp09qRPrahMf2fjxE35Hqz
cGXcGvP3S3vEjw8+sw/3fFXV9tzPTCIQ1VWrMwWK+DAOuBIMuxnweEgNoWtiEV0p
u7JSvnGqDPEIk9cNe61Q+iQrsRXGOqF+i7SMz8hbmlo+/MOBKvu4hJlTdnfPfXix
6mhcCS2IcKIq9aazGUR6sFNLAsN7EEiEP1WgqQYxgkEDRilrngcg1uuLwlaB/JOt
WvD17eNwf7K6eTz2BExmBnZga7cmM3FOc9FxRs73fQsDoSmrJ4XG794vpOTRdAcC
fCGju5WR3AG1ifZEiNtOuDe+ASfuOookL7HrofivBfiZ36vgCnScf+2aaIw/Cabl
b3ab1Vow6N0ShutiNE384fQIj20XZ+iSFcE63ZzrT1ZLrigryOvn7abflRRSZWQ7
ugCTq++2IAIfxdhnHDukbfiuuUcRpuLR774ieTl6HGk+t+xPUE4vtgI7/i34z+PU
mRGmTL+qYXO1kBnml5MBqKG/1YqaN23sp9lgzle1/fVByFRz4dMCCb7BY8ahy7Ln
4vTnwOva2JLaZPDSLuXl9yDCpReFjTGD7EPkXDJcP0126oFQ3cAsadloKIntqdhM
1HuS/KwyVzbexNOxc2PdJEGSumEn27/omosVn85mwvat/Rk3DhG5vCBDK8eaWZKe
zO3L/hn1mibZZmDzvv2AgKiFmqQWsZJQ9ZAWpiDEnxeyjzdVXkmFiwXY53PaOxnq
6H3v+U9Xw/YoTbOG0jFHD4tM3+Yl1AF2FzBqa15OUpSrueGVPJM0HfDQKykemavS
dbCNOgTs0xv7uucbkNPPbXRY38vH/CaMYffrNCCY9F4Uxy7flRrzXnEAAAtnWLmj
UhXP8It7dRdj2ltAsGbsiSTfvClFKS3uMkO7rwn3/Gsr+VQt4PZ7+vbDak6EVj3p
IcMnG/7/ExPLDzvsiFGFCYLuuhE0FN/cxYO+gKtWm1WZb6CYCpOJUcg00s/9tRTL
7MzWRHOyISkgriGZzyzFKBlRAYEaqMQZChvovCjgfREyFdQA3NG/fWOfTBNXZ+Ji
fpI8d/a/GCErhSv5GGq6zlxCFcbTZeHBg7kT3fzsIONXJjBlKhR/J29xgVeHEze+
tckLomSAxczh+69aep/8uvALC2gq7xuuLDGQzMj04h1pEPEJGSLkgomWNhg4e9wC
P58Mb7grgEjiegkLwLa/Pwu8Y1aZgezPLvKPCQ8F0R3Ubt/V3IHL4OUothUUkwsS
pGLJchU+T/NUHoQhJzlfoTbFeEDiIKz7znoaARU8e7E=
`protect END_PROTECTED
