`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nSEmSvmC/ng3cvs7HtKmGDhLMjYNUo89HDg9RRaiJpOvSGWM8L3o1ApJmMc57By
fF+PDZI62QZ2RSkKCFllcIssLJMYhnJ1VljycTqXIB3jeUFlhXNS/NEJUTTTpjpp
MFG0ZpcpaChWVfsU06d03rG5pJSfIErW2QXbF+5xoLPlnaK3jfsq1bqX7mbwCrlF
jl+RUMXDP43cIAod2TvwPNvDiyRhGYsbud52KauldcxLKCd0xfwEUOJTTt8j37Jv
g8x+lmaRZ676oC74KNYqICwJIBeRiZFFh0aZ60za0dItL689ju+eIX8rmuO8lmkh
swt83CG3kd9TRbmDsDvNC1UM1DaGyTiYAXc/EmtlK9NzizKFT14xWWSpCwg2vdcb
RQC/G6fx8De5c1Ubc0csD8UT0EBiUVxnOTRgG0eLNjjT19lhex83euAIP51C64o6
C3NJCs6qnwtysDxnBAL2JG9ZOd9xK6HLCdlAjbeb/rCWT+HK+sW1LDwCGwKSOclO
tZQgNmNTu6HGcl/vI9lzSiC0+e8yCtwkjf4n6PWxGaVYlzI2BcHgm28esBElwy3H
lrZK4gqIo4Dta/CHJXuarT9UB46rG2Wh1sgSAaQPnmKqu0/okPXfJF6hbSGqDm/2
MaMI40oXCqf8s9BPoscnd1yZEo05KMa/g82x9tsSPKpRpP28DuaRNnNRT1ZrE5S5
iPT6JC0pXayeZfM0tyyK7aKaVuyl88vIKdalGIwL+ys4R3be6ynIOr941IGw8tmW
qWmQizdQ5oU9mUUDGhvUbuUUOVhzDIrTZMq5ICXhByto/ish5Fa2e/mhK2W3+S/A
XsfTzLim3F6W+Ji8okE0b5s8R3JEcmwEggw81akS6rxb63rYOB7QQhWsUCMjzbcP
mKA6g2SFL0k5ZQijkYSlO1RW3yxPNva54c3KWB+EUmQpZmbqG7mdrnmA8kgTdo9S
RJndBym0zuRjwVUeJnFY7VIvsUxd61A1egkO0Qw+PDViNS84uARXsTjquc3yWR5s
dwcbNmxJ+L1fekOYCPTimq6h+4EiE9hrkzzn2sxr7OdrLofQF6na2Ypbjsjq3Bs0
GQutbff5gMepAfznOfyySM1Vx3hlo95yskGwOys4X9dNVj2dEHE0fsldHAknUtRn
iNIwoKYaDuygZbAJvlsK/DgeqH4SVkjXYrhWSE4mo0bSXHOjvT7tjwnuDEIZOSOt
rzXZ55GCeX7b0WUQXuBdDga5qWhdtUCTjbYHZ7lN3BV7TAME7DSqQks/wIwa+/v7
nnji1ZqCLjS7tbH1huQjYLudvHpjsMJISnO4eFGIgcImcm56FNxWGK+yEwmOhoNw
1svjJQqBuDdjPjnio0v87PNR0Sbfl1HGfqKseRnngNggn5ZxI7qfPb1Pd3yme0r7
OJV9WxQLDAHNJEFumOPCbUoOUDAp1REUzxvuhSWgk+xKOZbx5YWSnNO1K+13TY2Y
Z7sNHBr3Wzt0MjQ0JO3vOMYp7KftmeCXCRQFjoKRktP9abm7NahUDjFQI+WhUGBk
j+5Td47UJ9XM3btz0gyfhDXHPUQvEzCF2pFeYc8zl3VhecHYwnkK/xvQExdJS/MN
IZXkJqqcof14QeeF6lXp4+589RJtfeGtkmIigfY1j0TgbKuxH3m3o+Umuqr1C58S
0SAonExxfF/jpEFYnGvo+D4pfleHizoT+oiEldN45k5mJP8xSN4DgyuN+noJpLMJ
mwe9LdXy1xb8zl+/uz3w1rOgQoqLTjNCBBAzsMFuYa6Wg+1b35bDG96X/zmvsjmy
+uGw9nH+YXCntz7vYh7LRLPcFWLPAaCdAuhWAFPeJWWQ8wVaykcAI1dN0+qkFDKR
Qq81VdYdunHeLZvNf4bJYA/coSb3p4JXDzZUjOs07XKVEsf7vf5E2Ydf7XcGpvnh
Edrpy9FOkLrcTqhBfKujosFtrCTh+TSt6d0ROPbdQEpeC2cnJ4mlvXGLLD/j7DqL
vTjBPS6/AZtXWo3qM/NvlkAc78vqwvpbJMc/1TcNlqthTT3RWh2Ic9B+N0WzgMRI
afqYtsRyIOApTEVj2S16qJtI5vVoigaGl3QcwIOHNlH6tFZMgL8lvudMvZwSzbWq
7yMKyd9DxF3nuxQ2CGld/zVlVkZ2YmXUj++rkufguivcJz9Ll0WpLFLH5w18lXKk
xVhpKW7BsW/U17KnI2zpSvma4LS4UEg8p0WY4oxUmt7IT2vb54alNGRFuapffSFu
gKe0n20LMLHIZFkQ1SzNDCihJDFzxNLh7c3k6kSpe8BViScuoXVCLn0uIdvR8ufJ
PMl6wmFrFbzMhVIWGMahdMbNfpRB+CsuvGRVaDiMQmozQYCvKtnzWPdPlxb4t/zR
VUjlOO/mlhlrO46EHIFHb0Gx20I65MBmVC9af70nG7tSQr+nOU33UczefW4Xji7z
RT/mQEGFa/ygmTgqmKpVumHCh89qW8k9RHJee+W8IGDc0khSsP2jPXZC32QW0nxW
/qxzLR/p9g1UuvexrSixj5TYhfvZJYUOH/KAZcn4adHJAtZaEfmUu2fANsQKJ3FE
2oQMZdihMZyZbI/H4bokbWgACiIUpTo3/7VY8i7vepwuPAwFVTp7eWi4+8+KWb9v
yW6fiBS2uvvwtqUkffK/A/6rC1aKuf+A6Ydn4LXr74If0Sel2WbE/aOPEsNdvzvV
8FpUxu3RvSbCivDw7nvMv8lvs1BJg7PSmCrS0k4LNftL2JHCmQqOtmy8VagROXPP
AJ8Wu0RwPfwCaTeg5b2sS7rs3vZ+w9bxMwnXihtbXorP9W6Z8lKj6Zwa9LRm6qs0
IfaBdQscfk1Z9Vn2//w27gLOnOciuMRgF7VOJZgA9OfD/bXoeEwvtYHRfRnRwVgt
sWQJYgm9QrxQ3dhu9DsNiXF05Ljl3MArWdShyFPlLd2z3BV8dVCJHnLqzRZI1sht
38URRs66foWlpdyDo86ORQo9emJ8pNA9PPhCr7jKNwVoKDBkAZgUAwXKJATNRs3P
13AONfaEER2WtLsnSZObRq4XuHmgs5vPhcCDnp17soSabKmhsYAjn5jEf4PTVBEN
vW381/mVTbgN8SxZSTYBhuyS8G4IwL/Q+RsPLaaVx9VVEY4KxeYm30PESM7zYDZG
0kk48ZmiwgIzDVGZgnk3AL/7aKvG9J0EFwyFZImNKf5Zr8wlSsJxbbv0ybGkBvxo
BlUYnRQxGJYUk4pzCMTLQuUrWiyy9EIi+rFOuJ1kOqwx1oHMoz4TLfqDoSbv/o+D
4K72cM4aAN2b+s107+I3QZa5ZLuU8i7wx0A1ipiw18ZxTHDAB++vQVYoeXRkPYcZ
AuY9cI7YVhpzoinBF6pFypQl/jbuPrqf7nFJKD7BOKh2+SO1SABRCTrKH/mqThw5
R0Ey1AbQMt0XSL81+ou5LbmDP9sGeV3ZrNkaYNdygVlO9gmRraI2Qz+iMp0/ihZe
TUm469KQ6XGE0Nx7Qc8Q9rOe0el5ZLYlGSfYetdXitYHX/ys+kJRt4AoGBDQW2KE
yXqASJ4KWmulJSNlhGPRqQJqlFCn+XPhUTqZg5b3E/akDWqvhjC3Jr9ax7dqK9y6
plW3xz08o+4jCZcNmGP+nAgTvVWYDLjEmEIAxJBzhHEQLsAOYBASwmJOtWFCnzOn
gxeNp+vLlfUx7w4pcTXsuR6c8S0pGIOpY1ZQaQzuJeda6F+TsPmRo+DGtosdkpzq
G6bSy/TORg/NTvZ/AhNCYWQ1b7XC3C8dRz/HFEOGLZnjKM4ga7qU7qSmvu+i3Ffl
II8FOiXfZvMjIaDhB8aTjg5YDatpRAAdotqK3uF+mweEBYHrhXJNm93cfJ+wRgIs
Z/KxA4TY5REv8eGP9n+VwzXGS6gl/gaoyfBNqbvpi6xT/OQS+hA06/ucf4mJXmxW
Z/n3O6WfRnGgxiSw1zLJ7jcphbhoCu3ih4sxoJn7gennKymO9eiEEhat8qQUweTQ
jey2980RrPW5rWXiVfYaSmOkzlnRO7SAhjlp3lPWwqhh4wSS9ll0fij/+iLt2XWv
bvrJAH+SNJUAOYxOOSnev2fHULcqDjoeo9bfXwG7mwEAz3qyCD+9VfQ53aZaJy6q
9L4AcMoWrKt0gtfpz2JIa2TJ8hrsyAjJ1LYeoZBOuPiWd40Af4NRG52ZR9qEITHY
4IAI+HDH6OBCbGHWPZrE153NYpeVj3gNZnQiq36G3JJyj1JMKn99W32ll2utrx/L
VSVTaPMofupvMqaA3GmE1veFf7aTDE+vPWPqg57Wk1vrdDEo+dFvmRVRanWR+z9r
gv0cQv39XBcNTPrG/cwgcOmeUNAz0WEGHfAfATj/RvKPjF43HQvbfs1OFUwsJvMx
c9G7E50P/Lo6sMWoVTldBIPsLvsIfLOmOxdwhgCjoLXVST/C2favBC73alUWF8+v
9+0/NKswlrWAILIld5Vlmgs0JsVXfzs93YJ5NiVvLhm1NluO9IpenMBISDnUEbul
+waHnnG7x/9jzOXKySZTnKRsSrMRR+7mQYbam7NT4uwxt1hft88HC+zpZVNu5z5u
8REZGGsIuJPUfmC/Ft3smGrHqJqWYawBf+ANhmiOfh6bqXFFv5VxOaBz0oR7eKn5
V8nkiJ0FITArHFWk7PFe8Lq/YIoIqRm5IgwEc4aTTQ0Ivwwhezcw8Z7+jkK1oPuZ
gKQyrR5/KGgjx17fZAKUjw2S+gOoq4dkED+UYJSWLlnWe1DCSJ+AQpg65dfRGr8E
vxc8ML15tXu96K3AZpVRC3Qpc6cerLLje9XPl4Hp/MoplbYt66+iIlYUAmfVpnAo
PDgYpKZ2ziZyUscPveYRhnbyfnvNA4oelqxPb50YcSTQ2qWwbRBV6kuGWs6IJgj1
i9xm4rj0KqlRNp9OgbR2bSWKE5lKq2mfdC87iLDcFL7Zf+qEuupyC9zai+HoHd52
TExGn695ntyJBjfcyMBhT25c/oAFzTA7Ouq+fqWcrl7cvbL9ViWb7TT+oZYMYQvq
fdzhhlOucmi9+BMTssN3Mqv9kukUG0p9gWtzvoyNkAQY56OQJC7DJfcgG17COoo2
LK/PjPdLyeX/OUvY55DP/3irTSpZQ4JlSZveex3kWMNTFQpyqxBgAkWuwfThnu3L
bOGp7JbJ6QeVuNWu4yFjrG5lTYdKEzifMpC9jhctl7cgVprAe1B/hI7ZjXyBjnrK
FPjG7cJSlJ4cUs7O7c4aGzbqs7MogZUM6Ci7jV+4LAYm6dZsUvAgrHy+X6JaSZe0
w6/wu5ad05CY25XdgUANQUp/B/7ZL3AlHUJuAyBJ0r+c1UsWIZi2WL9ffg1KsYu4
4ZfnfTfzDGVrgo9qQfp+mnf/53zAugbbdXzGfA5ohtztqvdPKktnN+fBjYCkeNh2
thPp8fjZQUIgL9A4UOOcvhgJpOtY4DwZiBxUDi1CM1qAehmir/DEdpv27ROE3SN+
KxTIosS2B1GJ2PJgBdqkRe3eowjiFfiKMP2t0JiXkkIJgxoAMZ7ZKtcrBGm2xlD+
4KioDv6YV8ETKLQ48S9doOUYNBa/rXj3Dl4MTByUSJqkzHGviSOYCdrOIzI8biCz
mzbXVZTBOXsRHBRP0Obsq0oNa8Jy5n6948oH9udbB6uqJtUJHr5NPjU2FAYFWuY+
43GEMTtS8YstgRrW0nh1rcj5sblwTDe93ESz98sGWh14jtRY4LFehwi3Fa0+dpyG
tZOFCQuI1Yj1WfBEl5gMQ2SXY4l3rcOq1YT25eu9p/07r2J4xDbTJQVLdLZaSMWr
GzO/Ix/jzPPsHBvdKjt2y+tq+InklT5/pAvWJtiyFsVo7pz4RUjWGSRbJES/g/oT
Jl7U6ED3hcDLJx2qKAnMRqcrACrGo+b/qPNzSP07j7MnpYH5/SkZX11oxAgR+L44
PXnp0xZMRnYg7K5ADZmbjb9m3UPRt3IhT8rr+7Adse11688TbQMCswa25rEb5QDj
idW2wdvGjDdbL37ZF1NDqFt8Gpbx0nKrhj33NV01P89ea55hv8+WUnORJjelP3DQ
MHRFGF3h1ROkt1ScGCyYqGIxIyAxs3dEpFxTsiLvin1G1cINFbDNJjLjjDkIhp0k
6N+kRKE/m67NZSXC/zxRh7/n9utSrFywNFWhuVzb4ZrI4B/HSyYqpzIau7TB9MlV
WBL/L22Bs/UyoQ9Y/93OwKMx96aNBxpqgD3I8A0kRxNLPymeWr06RbGJ/b6v/NF3
8cSQyCfCuZQaEPSQu/+yQhijNm4MKXYSvMN4LMfF009AcK/kDkSQyyHpHjSU/z10
8wsvDReVsXC65yFdoN414gc/9unX5YxGJjRIcAFM6eshlHsh74n+k+3Uq/S8xmNe
gXgGUk1oAsloO/imIbViCoKgD/ksqw4zjtKGyF6PK0ceIbdysyF4G+weqzzNATV2
zEufl7htUVIp2xWH86zIDtvcy9wXEuDywMsoe1ZLRVsR/kWmWjynYwN3c2FGFVFM
CcwZWeHEoKTToSR8sjdZ5L8cMFRutrUueOl6iI37bpYGqgnNFYlUT5AMH6p38AUO
V2XHnlU9loFxhP+bXAb7w3sGPwODPNHWEUvyUPCSOcyxkhWGkEkBx5UNtCpEVjvh
iYUQia7V2JetntpUEyi42IxSOu2tpx/qkIoZwhJ3r2o9j9/PHucHDdwIyg3kwmBn
3Ud4Rq41LW3+uQMsrepKt7smkh3EFvzvXFtvtfTjlNtwpEgmAmmbKbSE1hal6v/L
Jnob5+ZqxYDDxEmBymUwY64uYbX/zCxW1SCqMxHgUE4J6A0bMA7eDQUOJh+cwji9
7+ClyFxeLiVKHs6gdwP+7GapQ+dKuebRo8Mbiy32dbBbK4F8v2T0UbpDvenqnLPz
F28NRFfofU4SxmpLr2FAZNoWry02vou0kzm0Jpkg/PwfhV+P0LDBLRoY8QOxdvX3
mhC8oICSs4ttQuMMXTwrJFCMgJcSckKV6HXytQwlVtx0ycQKLaK14CAGuOI5/z/i
AO4/0CH0fFym1mLhaQHs0ka6mrAn98ejxmFcJqsGTK1zrz6yi4LZWzZh5UCK+fDX
hCzgP9tOa2CBmmav6nSC/StXbe54T4GzNyGRoo1DvVc+Dszt1Qlr+XhvyCHXjXgv
UtNayLbg1QvXbKZS9OE2DjgDC1wgNkzzmN4DybP1hGzDIIjVzD8ODiJKrtXZ+8Je
bqFZmCgc7ybLek/hv/ctpOf+0uEpuphjwBikQDsV98I=
`protect END_PROTECTED
