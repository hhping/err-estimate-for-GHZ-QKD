`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v6Dcm28fRCbrFV0MNVzdghFPze3FQ0utFdj9wVHNK8OYFQx1YjvlNgpfcFqsqZsk
EQgDP1P+ri2W78ss5sAT6tPXmNC5kMWkubTCfYgoZ58DasvC9e6lGfGj+ukoE+fP
p0O0yE8M3RiFuPYMXylmSCJB5hu4y7PRg0sKhF7QfpJtJQw1CcrQz9NTMiHg4M9w
7NovpmvdIMJIIjTE7nWqBSBhDoQtpv0YCAj7QBjyt8EyL+0YGf6ifIedJClHFHGV
NZKDHZtYlulwGlZKZ8SvIHwbEfkkD5JGC580WD7zFnC2jOA5oCf6DSjlqR0U8KOd
Sysfn/lPfVRzywZGeWnN6vXcBsNg+eTFR7baX7z0nAuJ4UlMgG6oro6aR24MymHw
IiAhrrJcosIc0KLiFWyfpX/lYDW+kKkJ6sMc7C8BlAjw/I37thXeDgiCgM58JG8g
a7N6e903QfjqW0IKFHq79DRb/hK4f5MCPzgLNRxMIfScfBoQpYQPw1eA0jnPsVaH
8eWn7bFcXGmSaEmN8XOWcd1PWsqaCgAzCPGgDOkSfOb74dSc36PvF8Kq3EDLmuh0
y7wkx5P7LiHrXXTJ/uwoWcxEgQGKtf3YhtfwSTk4Lp6Nz65ktOFsdREMOLTbqSZr
T1qqlFmd5KWerpQpk3A0z4YN74uQK/aV2tupseXkvXuOhVmgcC0t0mkkFDsIb8Gg
k8kt+rwjHvU3g8ozCjiIarK7fo3nvUeJ5qIGgzf6Bjf11pEU7+dKqRZ/s7ZPPB3H
IR3/Op0q6FNFw3ViWESAsKm5W1p+ukEYM7pwPKjlljv0x2nRqIdofY7VRYvzDltq
wNQnEdh9UVQAMfuJwsOuNLI96VeZc5miVjClfkB697joMPwEz96hRAtuYZ45gIuB
hp7Yv8iMT4HEJnmBDor1x96UlQ8jHu+7vVrCxaX4foCp8qIoaZJiWpoBJ+XB0wku
igHV5sKkiTV16McQM0GI0u90N/iSegznk0hYGibBhLL7zOY3ceoyerEoQaCW1ElU
PzvelMvNix17ACUt9AfCI/FDDsqTgfmoGjMp8aw+fnbCjNfPwVLCwz58L0WG9+J0
5mKQ3gbaRJCSfJ2F+MPbKw5QLWrWvAwjxLkvlNKdsOy9z2DBHvapBBhn+QHOhSOl
RpQ3Cy1OptE4gb4Nb2VlW8JYL8CTDNWqpyB9+C7AeNcvJWtquf+G4EPbkmmQ7K3z
QfqW7G1QQ693yjrUJ4txn1tYA09QqDDzQx7CYvqQE4dEMk2PFPidzG/WOKQpkf/D
HopQy8bCyE0Izj48bfv7BFgvERmyAHJaMy/tFwFqJc8KUu2AZ6wktvs7dfGyYVjK
50edx9QvIKBtfK1JBG0JrifBvEYapF83+gQwhSHF8MKSiTD+6b6PLUsFSeKK8aZH
fPNTCSnVgjzsYjoDqNoMB6HbscQntBOoE9sHuF8uIPaZfg/PEVIjLw4jMU4PacTB
HTTArl+U0pI1TeHSn7nmkoe64+pMD7M/LQI6rKzmNOQ5WwSl3X9dWYJSIzrElleQ
uX+UyZjjNeTw/yjZtIg9SILyf5RRju2HnWv2QCB/XovcqxhHAuPNNKRs1HTrHOuW
Ja7Agyr7wkCoqwaDeqQOpL0Vv7hjosyD3rhawIG9IFZqxLoqKa7o0XS3zhtNd/3+
gBafN5uEXGvWgzgixMMlR79NQ6YnRbDQiYaQC7OeSrtvHCNmg7/k6agNyUO7iasn
LShDBEyJ6lQbWEBV7hv/JtPydLJ7HDLKCBslsre8/9dR33asMsPQCrD1QVI19Crh
TdDAfbYF7AkmPUJMt3/UpBF/4KM/2egz7ivvK+AaXNn4+KvNBc/d+UISf6zgj/7O
+YLbz6S7k9FdDF6YmPED/B1qwz0YGEHUwVJ0fd4LUiKtCwddQETQ6KVawIOcymSr
ov7f9QUHFvRJ/R536V6Bo0/QepURVHpqMtEsS62Ym2ol4YOeIoQBBFRUTgouHwV5
MDp1leQwDXUKgBajLICBrxG5+eMIkJAATgZAnr1yaEWk4evXYNDHShDxrG3tfvm7
/50Z6ykLI2odXc6xGpGS8Y5XO9Ao/MVNc5g2AaUiQwTcKP9a5+/qAfyxqnnkVVBE
JCSQEswKAYjYkwfR7CV/CjRSOh+YuWSD7yq+HfMkmNLMTmIcABz7R62Jotq572i2
tSQCWXSBTdU59jLBgA2XsYwp+Hb5cS2wxutyELEVDeU0JM++P9TkIX/In/kuESHI
OhCgxjy6oIicd+HWiCHXZ840fQqc2JpZVgX4jIy41zxLLfwHstSB2s/n5fptbjQU
Sg48S9I9uI6O/d6s+J3HaPBZyCHi/S6tm01f+ozNNDFZCN9FKfnVGDAX1DU7bmus
HwZ/pZXjk8VV5e6yRRf3xqYbdcDgc/4BG23OLVZhEDl4sXq+PHFk6nQu8JRuympd
zDy2q1Yu1fohUj9gsHbRWzu6tv/hUCmcWMxsaS23x4GTExhBOjWU1rJuiw154enc
doEOiVmHTQWkpqiUJZ+8aeTAQNdHn2vA4gYL9RnpzoV82gWPY4kPVPuM1V+SoYw3
7Z0MMjeNIfdq7kL9zJG9Ip6+4iIu8Q0QfI+GQJFQAZTVckV4WugU6h/EhPAtLP3E
bhz58mDuDZaLROEhbgtahnxKhQUKNns4XKeH96To2RQSXJd2k6ggnPTs3/PqdDuS
4SaFrCQibnKia18aRYrMquBuIQozdTrH3J9BR8RALUJtVb/dC4JXZYMl3XBKEm/o
slWZ+2yacQti/OxydL9IjPIiFqG11a99GU0hhNTw3/j6iAQt7H24FspKjkUv8p1w
mjClTtFXwAUmhx+m69mpa9DvQKRGt+WxOHnd9tvN4FMFAQiCvVNZP6Ecd2080DH8
k6J25SjBsFatP6PEqnfgL1aA0mAZlg14jDqH8PvMdCXjFNEmq7tXGl2gb0UosMqU
qstGZxjfELpYDOpcBbIub7lyTMTJsd7RVaGa63f7V+f1sA3zRIl/Dv2w16KteoVW
n+G3z9XyMmRrdgcb09D8msn2dBthkGOg+q3VJQyOUe5n+ywgUAjP/9jKgbUDfDVT
QVYeUet1caoRWXcccM66GJ6RvcI5hleyH4efzKtjuXgUgsWOw8Ggi3dm8eG7kQ74
FvDkhHaLNqkXHXYWOuaoi3VxqJ4WrCaktOF4KBGsycngOyFOWaVyxKyBjV28c/Yk
yCtQLr24zg5DgKC2B3Rov4HlncjJldfJ9g4VFBO/QdH/yZ+Nse3UkDTjW4Mg6uH6
mNgQVq0wRFhGA8q9ccxZeHB5fpVQb+RlDcKvO+UMtCkzg3EGvUvUpQ4R6+zgq5OH
YcSZSpTxQKrjiAHW+keaidFsP4ac5kyGcpDLZ1Ljyq7wGhyc8uRLR/GEMfeBR3xF
+yqfOvkfQtP+Xsklvn78Z8gjHdMV9m+aiz5bVEushEQQIrM+dcHHwnEvZFE98jDe
8HWjWyovhk9DTWpFPx+EckrHBFyCM3BYpOjJU+e0DKcbIw554x3hkoHbouVulIlj
7QnJOEa5moiR1lGDWzzoTo/UqSF7eEtD5dOcdaodLw+u4BX4Wr/8mKC24HpKcHI6
xBc03XOTQyqm2yJ3b+E1u0CUrUB3cXYGLvl7rhiegoC8rK+lDtq5/ku08fPKhGi1
AJpaVvTW2ACFqC7Odl+CfOwXFnsQQ9acwAGF1DjA1tgcA1ZbhtfFhUYFZaV95PZo
JdFChzFneZOFZ+Nxuhixb9dIw3bsaZmCFvhnQnBHC3Dp2kk2+cGJbwOH5ZWHl6qQ
CpRm0Kw/OVWJjMjBklp0oIlxYb4pQOikNMngC+iEljwpRKZtg1CFiWpt/UnhyHAe
46DQAnkOO2EcnvwLhBwV9yhvhPhHJ6A7MxDN4ONtIzy5q/aDnqmf/Nra7uvl2lqC
zX0/uAVvExf8CAWJtlrO7z3Awf8DOO6durnwHoe9ddSNkZ4hVmpk59cj/m6HJSzu
BXdvESeV35s/aa/47INbOXw0BUvskVF+8PVsoH1/VElJaMBcg+h3rowR3qIJLaDs
Wt+yYh9APtBLp5oB2zqKv+kTqJ2KMS/HAK8jeVOsNIEjYPcFVtZzdvGnHI0KF5C5
C6YNEriykEUNpckQbiIkXFN0tbr6GWJFqw5vaZTak0Vs86dyzfRDS7r+ZpgZnk6F
8cK2QO7W0r+cJ6TZ/eaxri1UghYaBPMbqG48+p0+SsM0Y8HGN5Ef9R2D4LJNwRXs
`protect END_PROTECTED
