`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hO5bnda65MPL+IE1YginfNF3ZhHsEkKEWWr08m6p4ok4d9MQXFLZ5r1PQy3XQLh0
wns4YCzBJOTRHUvMxWLw6lsZPZwn4NiLS2qaz3a7K+9+wlquCzpxIkryg/SNKTEf
hCfBTV3tQO7MYJgHaN2vhNPHaPQAD0QLJtNQlLfx82SzT2LQPyv4d+KUSI4FX8Qb
fuJ2mj5W+GlnDikx0Apn5scR182Yxi7f453mo7gcBcrBLiaIuHfuosIk8VZl6T7M
dbobxiBDWM2UXu8qXulukDRHojaUFDojcHjE60Qzq7Nj2CcTd0SAKSNedCDU0YHh
DvcapnFkv9LrM5ODLbXFlVDrLjbZCsxP1qtKXD6IryD6zptxRepX5WVnIOFfA+UF
a0wC8GJGVpv2xQZyMqTyYs5CfXVHZ6fg7baJh4Trf+yUnowPFDJEsmTdeu/WC2Fd
EIK79y4CV4D5Uy0q/71e0EIcJKqL/ghDHxY5Xz5Ob2I=
`protect END_PROTECTED
