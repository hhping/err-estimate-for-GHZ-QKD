`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HEjztk+yzs2c2z5vMY0R4n0C4ixsq22md4E2jKz95OlmlrCBwzUayIucm02AUVx
zFnuqdYFF5HFpS279A6qXFhMePJfhnX2VQrlqW46n3++zrckKDuXlu+9UlDSo1Wp
ViLSAJPQ6cyfLw+aXdYRwJF7+rhTk+3Nc5XF1TZmClG8d6loanqwRg9Z1cmWx479
j+vVc2JsQ7zbDM4rZ+63f1leqVoYAaUFznm6oCMYHvLjYH+tmRDu2D+nqGeheXLS
uajGDp1/+vJQ+fPnIy5WlgmREmnx4H0NklJtVFtW7pn1kMKtGrDK2JjBrb8cvwyF
ww/UtZYoGgeqI1AzyceLVrEQPtt9RUfXZbLMKmSeEnY2eSsnVukOMO151Ungavln
/mUKgZ/sb9th/B3L+YrnHvZDmDCA8Iwpta5S/NqQWwlsBNUkdZnHlR+9hpk1NiPM
ox5QgqTyUobJfn66c6TMxw==
`protect END_PROTECTED
