`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxTf2vIzxUfZcqEBCnPkZz9bfbC/6e2HvzDfqoY//FC62f9ya8ifMhQHon1Aokqe
a5QIKwkEmOnum2g+xZN7pg5/b6vFiKMAipB3BXoIjNEP6XwjTe93k5H17mvUV+iK
op6f7kQDc+UARIk0yWxbrfSwdPfKEh5ySKL16Y7G4rdLqPb9pMHGXLEAlrnpqLn0
/QZ0B85+kI13EwBvAqtQ3IginXZT7PA09EFYQ9qS4Jo/euxRoCWENLeqnUg6o40E
WuRVRfnJFs6FqLmd4CaPs9cPZvI1vQO7/jQKvy0ascuH+6IcoKcieqRqSuYMDvoa
jgT6lwDSZ636NsuhNrzRUoJsT4mghEldcgSS83ICn6zBzh6drgFl/NO1v+uypxBX
5pO3WLPZSsx8oP1Tvqo9Y8zNmf+0scBYyw45ghMFu3vu8eH1pS+a3l0zl2wwuUFM
n4oAKQiFWPtOcquSoYdHYtHpxWzu4Xt9PvHEwqvN9WzqA1siYmtzM+hGO7HwAi2n
dYwpQd8tfTHZz5z4snNUNa2gpP8HuBfwrGCkDiM6pb+u3HzhBLcwM+EgeWJ/HNpe
Bqwk5xh6D7y+s4/XxYIOCKgHJ21EvPoOrfHmMcfzOYkifXvva8OpsFIkTSX6kjju
DdPll0Wg8hAt5UCNzTHmzdlzHekCXsknvCl4DQup418a2c/025mQb3YDTv/7SDUh
ZUI9sLPJXvnLTqRGwT0gLR8pxLhRqQ8xovW/T4DeTtLm5+EiFa1jtZI7grFGLp1k
/cPBIT7pzjv1ByAMUSSbF04Hx6Uql827TCDvfgI/0rXturWdV7i15focc7HReK5i
r69AiysAWU5ZbRK3aYB1m1jm8cXggX3RtYdlPegDHz1hA6tyIVQ/kvBjH9uCV4MT
3ufaNbQGS2+Al7+dosMtBaIEyILEbLzhmkj2E+/q8B3prToAZj9Da8juidH08Zpo
XHhDYOC8sDvjjXCrLlC/dzUScICuj1fzBaSg5LYFCrbEa/TKLDlwwV9SACktklxk
MYvKCShcQoYyl8WEnQGxpZArTQs0iE4FDzvoYghq59IASpd0SzLC1lgLzr4DjWQ7
xYoP42HUQk/8oRy/rPERQ8QVI8+HMEG/Jddxl7mjWtRIk5eMBXh+WAPzQJmFWmah
jZsxf0qSSAheZcJgINUtMBb2X1YhxU8Jrz5BDgEpcrBcXu+hp7M8L3vSUWHpycqt
0J/e0qjfpWEnsHnqfw4fOXqbwsgHMaDwiwsFBhPcDB4HjmYqDshE18yP3xuuH1gU
Y8zCvYMYj5xpqL1mNxFyRaosE8lMZfbRpcWoRI47wFcEV+Xda0vDYl09xW9O9cbW
tghHOtHmBOoTz8DlFtifGEu+Xp1dcJpb8aNzl2Yx9N6D5Ehq9l1mpLskttgPYrpH
HbHahNkeTet5jAIRZmiFsGo+eR0ffw7Evypoi9ZEfWUYHFH09waI2epa1IhoLZWL
5YIr5qhH7TfRbmqi9EpoWKyjlTYUjFL65yHd/rGPe224Kt531Ad/oSXRl8S58NBH
OYUrW6O80bYw92bfuShqJGO6P/t148+Di8NX1xGnVZav8rnwYfw9rrAM8bog3YkW
ym3RVaoiQuaFZt8wFkkKby2kLYCewVY+PVIwhBiefXoII8FFQ0oZL2UyWpzcEhGR
ikBKFCArezhghE2NnRUfDqC3fqAAKPqE1lDF4vjOd8IujIpWap9nqeeGNelvYxfn
VGKnmRf1VmOpfHWHRJeS0AmG3iSVewLXFaAYXoOeW80=
`protect END_PROTECTED
