`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1g+ZKbRxNuL19rtEBMTki6GIkWON+u9Ajn9N5QTMe+/h6J9V6SSIlNF/uomM5lo
kOvOxMcuWTTjKHrVgEvmRlLHyPudLP5nckMM3QGKgZojrZsbDVUK1V1T7/7omNTz
H+J7sv7f/rmMU244GQFg0ZmdXow5pw2PWm1/EWR+FSOziRATjynQXvqhEHffonB6
UVTWMWlDmdLyEjuJQRaw144bMBhvXXBk/Fusw/llL/So2RgLzwM1oh/Ca9hNvcpA
H0klnG5WRn58YmTCkCJ9/IdrZ1UAb9XnLlbTRi9gMEFmpJ3NZab/wf9xw0V2ehJe
vSeXEi5OIeUOULZND9eh6WXprEx8v+G8Lwul1Kj6cL56se4g9+u9z8HXj6i6OpW5
exKpbNKTMcD2zotomReB7pdWYrBrw3HucRhOE+uLmoPf7LZi6SeC2T6hqpaYFnyU
MzoXDPvcfmVTZrR4LuDU6c0go8fUSONafYG/EC7muB2Ye59IrBtOf9trkSeXPuP2
94XtLU588L0SHJbUA8iyGrc7nQk+aiGqBl4q7ahhXGoSo7GTmpeJuFZGX9xNOl5b
2ss+uLpvIWQoMMZ1skrX4bXzVeES6T+ZclRVPnX/bevGqiWTwHH+kpcgDHgI3LkY
GRGMXA7oYdk+yZAE4O8U43Eh3cU8XFFCOPNFkbVZV5dAAkUahAYu1YzcSSkZ//F3
SibuOIvF7qe5B66I7kbUHQDFg+jVPmeIi/wgEJZeqLjr7UmbZcDBGPsDtAVeFqIo
p7UWIS9gOAx/X1hRKY2tCscDKXdrXhXQAEcKoS4ULmpBo1NacBnSKvxce5cbBSKh
pqH0CWaZXR18SN1EqiKfak+BbeaMMWWELYkpK9V//Ub69XvWkM8wlL4ydu36fv/M
bxCTB8HByQpiRUMllrEdqQAY/hc+plI1ga0qD24t5/Or9T78bS+sMeeXa7e9z3+G
Xc18FYr7RSfJZ0tnq8AiztGXunAKQu2uLYMhEeO6v9L23KhWhtpbcUa4pjqIJ/2c
`protect END_PROTECTED
