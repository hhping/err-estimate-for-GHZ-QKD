`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ke6Tao0SNB1M7w+99NkduS/v5B8NW/y0UPw4Vgkvj/uk0FQZGAdJefYu2A1aZyS/
hdtn3ckoRFbQ15wZLII1PUXxFJgkKk85hKDS2TJuMEv57uqn+jO5c98fjdZ/YaOT
kKRuXgesxlGYWgdciuICy9n1wwvafLg5F6c+LgPGBuv8CN1DobXAUmrMXqennieE
C1lP+W5l1cYOcnm+OgMmuoQPoySeK6+Lg6ovRnSWQWIpjZYx1+i+ZSbYC0Fyl6m6
ZWTrx0Xay7+3G3pJ1lb9zJafjzC63LfnYIbjIJDnNLi0gnycHGSVGcf/ShTl6GV4
Kjfe5WrHXVtzzkjcVvR0QicLdwOnWSA3L/vEN7AlhY5rlpJOx717rlzBIr8qKagX
wTWCSzCkBEZweXSTJ0DZ2JbRAie4rQaXAs1OszT7AYBmhQGhY2gBL/54FlNd2Lr6
vjZM9KVgX5wofEiDkyOwGk/zSf1T2N68uC5J+IZDSLBoiCru2DTcJvIg4BMAWbcU
j7gnAPyDouTpScNUr2tkoH5u8+85oqBwHOOdvSOwM8xp+Ug1FGWb334OxdZ0kYrx
mnOekcESuYUPw3GLThhVlC/cL1VP5xJFN8ERhKxFoYJSjeWs6538RciIQbIr+IxU
tdqDSdVhRyI4riMY7yRnrFTXWQrf3rGYazQrCpN8WahBDpyBEUR5dVzmS7tY3sDg
Lo6yMo+y87BpAlDrSaBedlZrf5dd0/KWi98ZqEki50WT0pgyFru5Byk+4IDqYdFS
nkbCLn+y3FjWjBxpflTXRMEXaVgLsNjeB6eDzOv1BwUYa42D3cpwhu8W+mbzyPyQ
Ti/oDsZaycrAYFrI7f49S34z33I2VCJeTVvqLGSsfLbQPXNNLh80qEVD6Ayd412A
hyQOznXWOXcwsRzxBuhFu5b2Ljzp6Rh552TuXqxLKBEk808Z7r9wnehzZevKknLm
mrFqzO7BAOz2yLWp7T894UEmr8aRfLWYkO7hYT7lbB5kJ40xKeiKAQluqLm5LaEi
Gz4mB8Qiz7Om3e6r+SVOP46q5P4WniFzbKEjCQ4vq2slqQhOx07skHkq3CncQaKU
+1jQyH4+sk7xfZSTa+QZO0BJlDVJlF6zm0Cv8Wl8ISy+01PnbFyL2UQHFdsOOnGu
3MahkXmle7gHTY0muapxSwhFgbvnTejFnYw9j8eb4qygtbicUgh0Lo79NEaOSqqk
c/XtQT8R7zEqHnVAGKm4Hfi+Vhxnabb/NnLG21Wyr7LfNWJIZZYFZoUm+QtS0lqE
83x0sq4Bc/6ZiIkZsBQ4a2ee4VoSq87Em5HL5OoRBOS7jBr0lrzqeih0lSsX6ekA
/J3gINHFtzpH/SZxNHmgZzveTz0l/bIVnPsTGYT3U4859+9Bkx6Zxzem8IBkonBl
u0NW9QOnuYEkSifwcue+qkQAPVQ2oQA5O2R+RSgpSKzrAQnlU41nW5b49L7b7XEu
VUZDOoZ7pTWwJ6Vo5NVxShg4Y/WJEvctkegGrinw2dY1Gad2nDHXUWdGL1Mo0QOE
I4H6AeNn7ChP+gUJHGJ6BQApD/aD9YnUpLNMhAkHRPPUZJAlF8DI02/6hm+UjOXv
/DOxbtDUBEgKVSIIekT/nETOtVpvOxKkzcyp/rvuw7+GI87+zayeKzGVIAd6s/DI
1FED9grFaCGbUqRspCkqWBvy3cy56EpZ8VSLNES/P+nwdq73jh07HzRGmNTpbSCV
l3liWjyDwexwD5Xe7syoaUQ2HI35YMzc1sFuV79ReXM79KY1YhQ5I74TmJWdmTbB
n7y8aCLg5KmepA6FKlgUlkJwUL6s3+fIrBd1A0jvz+uPwiCKNaFWKd4Nmc23y1f6
sJ3wjFulAqKHl5+y4BABjGgn4eqjG2AEL+QOvMA5T5xvjy4AttdjY5fJwR6EgRAS
Qr9lE1K5oP3dBCd35VW/JV8OctKytZQgBO/3ZFTJcd8nWt5TDVJ6RjyoewwuCSvV
xm6xmwvuNFn6b00dfS2/YVPk5ZJtEyFO3YStQmc0KXhDUwJhJ79COM9UJeKW+pza
U1cFnWhQnKLh6aeZXgQQA68BcZi7PGdHSdWody3hFwoedP2d5dJeRDnKq7sp6AAJ
lxuh7MstmnTdXvDgE/1wrHTHaZxlZ8RJm1LuIpWVp2zNbrZk9+8MSxmaz3zlAqcW
Jcy46iLcT0nLhf7d04oSpi2pEfrZUjxEUHK6NHdg7CbUGFTzngUZK7SVZTxeJJfY
2TW7mbf7yi2im7vp8s4e52qKaIRO46ix0FHkiDK3cMMRIHWns6V5KMZEp2KD+DT3
h9J4rTInTEh06/+e+Yiqoft+BgxOhPHuKLuPHUPWOxeGVcruG9RYUeQZlCCQy2s6
YsoQp2MqpFSERfoCH4tJgP/NUIUb40TcKw5sYVAf/XKeyROtferTwCVSTCooGKlE
eYvmWJgiR4taO4csV/6vuEnSwdXXU0KlLnSECCQsIzr7kN3jLqIZmcDrddgJioJE
cbBX3HRenwaPO828pAHVJyFcnb7D1rwpDkzRayiAeGtqFFUTvtZX3spl6ubk2lB8
+odH5YZn11WLRmZREgGcj2oDnVTlNucioo07tH/EPjdT/F1lMEPU1hQp83sQjOPH
h6aitp9koeBgeEtB1UZ3R76/44QWz9m8+YI2nz3jKCPcx+euyUG34jg4a9eXjnyF
eeHf1uTlNC9ev+NL434h+wF/Y/I7QHSWEfsd8HZNV4gxF4wOGZjpg970Vw6xsW2n
ZejiYGir/caEjYxvzRgZpLaR/+33YBqeWDvaDitynQCy+1HoMjVh2soTIMAsi9jU
+Aj9CdGyvjKcEzVRseu22pa4lxDlmFTH7UgVZ2+aA3zAz0YlUPDhuF6qzz5Nrh6j
VS/v16n9O8LKlfn0MUYNYFCFUgLw5sMKmHA+0TmDgRirettO+/s16a0jpZjejylQ
o5gpbwHtZGY2z0cAgTMkSXOxlTLMs7jqGYNSpAxPv5zC3B87I5x/yBG3fNL9O0dZ
cnNjQzzsOAlflMhY3X9tBOonz33vHXebKG5hCADVHrXfcLwlCXMwCIBmQ6THXvcO
ZtpVFT4ELY5kcpB+bHaUupUo9rUTIL6Xuj8wus/8rrZ2dmcrVjA03g0emMu8HxbP
ydNOf5nn4jF2h+fPOFiEN6WD70qt5VMxDBOg3NENQ2rYGOaDw05RbE+LBlhNz1AR
GXx7LOBd9l5xnXzK6Z6CkfAwnSqMCZbUK/pn4vIzMAKIo5hD0RVSIppb/QaotWGj
wrGEDmY0g4c6Iyg+x1yj+9JfLspDkTISw85eetkIs1eF11PXqkOUfmwWhFANArmK
2a6fHio9jftCkH1TvBilErzzKtmz9hz9USmqHhOYSAC35ATt7AEo1uHoYHLT+yY5
frqRZ01Gg4h38SI/QlwtW1c9/Y30Lb07VWVZkUjsyFlS5bazTx1dUDA68cbbQFaZ
qQKdNOicOtoFwNSFP0o/Tw90b9CkZo5tSL+66Bj8YxtyoCeYPX3Z4aOgzThDYSHc
cCPM+3w5iBkbhS6QZCvvj6nlLFR7Qvxj1zty9UgPdb4QhDiThkS57V8DXd0YEgFI
+ZJRKqwonNdGuZh/eTuozNUvkuhB5Bsa2iEMq7Nrhwi2kPa/CAp256Zcc6Gc02Lm
ZVO4Vvu1es28O0T1elEIDx3lbVWcuQt14zG+U9b4gTygaIYRgOb5NE0aAFS8KDym
MsiFRV2ftmJSgyZNd/EGVGd8cllR7hYqfwtR71orOsfRFnflF9kDEfXU1T+URPrb
gd/HWyi0WlvXip1z2SaearKLAN/Qd2CngGu8GkDgvHyspL5vE/GExckpMDDHWu2E
FLEkfPkJT0xMYQetaaM3goCXOI3+uUnBeLRCHTTf61qN6Gszp0HbZqAohiL6oxqm
XY2osb33P7AZdnuVBtIdOA2TZ/iHoEuaNOhujAHgVMrQclY1jxPVSyxhJD2toynb
oKBJ1RNnmJxlFz8vpk3wYXUAQn49q4a2xOBQill/n7ryDjvAgeUg+lMqNhFPqonV
SO5VvVYmGG2SWZZr7K1QgzXq8RXYs3STYMoxHhANVSMmGctNrXsZBYA6wjoNhT8N
4gn42MOwnvMVytWcMA0C1sS7PmYylWBGvx1QnI2jNauSyQIbByxBeDexpTLrmITA
JIKs+w2bWg6+d9Vx3bRBM3nvdy8uKV+eenC6LRJiYtf0k38mA7kcZ/R8ijNM+/dy
r6VyIW/oSaTTEP+ugywMvc1R3Dw1BASsimEo9VN20CaUGEnkZcOtr4Jm05sRbPiH
hjm2UjCKlnijdW5gJhLuJbI1E56XmKzxIsTcN6VWjhEnVEoF3nWH5p37BenFYaOj
rsVJN/M1gWLqidVMOytqnISKXxD0Grb0sqwzoi5tQt6Mou9QTx0fuFJILJrWqCTP
IUndzSxzxxVl+JQMrNSsP8n7RlDSrY0oate3QjYWxwoYliCFNN+ptMeHxaZowDl1
gkG7lL7y1jlpriuIziAb3clXU0MRyuOLT4+jZs+6w1qtcuyyWL2TA5V+JWHZixbP
I2Z45uN7x1plUJSHNkWFfeDhXVfK0+GnSRGuhuPCs1ty1DqeMPBI578RMTtFuMGJ
SBqEhBzU8uRSHfL88KUIAsIiQmuU2dXM9Ce1WmC1AoIhG8/IToDqSsrbbMrlnl2N
NvC5bLYkf87/aSK9NNiVx1FiefToWOsImZFCMTQfmwIAB3gCtNctIpHjD2zAQdvF
Je1fvdtCpoeNO3YkpmkIHKOq6VtwSJS5UQxiCkgHao92RbhJtVyIxhkgNqaPUtxC
vTpBFZaZOunMfYHExj+eZbh6bWj9tmskLqg7uGUTCtZ6zUQXyrgQIWUXfl2RW2Jt
ojl8cWvwVCqwWRqZVqEEtJ43scbmVXOiKynXoAdS7AjGS+0e/zu0nkajxjlNfy1Q
TR1nl8LPJWi+7nBNZb9+FAuQjHJtV+Fs2KAuRuqM+KXHhNoXpQppSYQLWu0d3Rgw
tZhzrdWZEtjGRJCG4WrYeX/GrmDFra0JsngnYmpbiwZw02YuqgBlF5VywodFJ5WM
SAUgdDVWhTlFzAQ9BLq4hti3o1MBz43kKrVFS3G0OEiHCbyoTBA5DwhWoBUJqXHb
/VpYG5V4mvsyXuSIWgQY4eIuZw453yR5WYOe+rJ0qqg/LBqnzfCa0pxExlCP1uEw
40SZFVNQ3YNxI/pdgC4RI5sk+HaKAwEkrBijlDkBB7YBDll9mDh/1U8cGRTys5/W
91U11ub1PDcMwFeYh628lLvjIZvDgnxZNxOY6wboPrq4D1pdCAXqeAfSHvwMP9tn
YwbPS1FH19HgCBdvH5nDBk2iC9NOi3WWR6d6zwmbUob+2GgdaNVwEbPBLEF6MsoC
QPJMfN+gZpjN6nf6KrusNi0wwie18r7wUBIeQRST3sScE8SKsF9OMn8KUAOb0+IC
nufvEIGb25y6OsAys+wwxXTSA/O9/QGb7iVJSu/+6IhJWYGLhw11uqFBCScLzBY9
HKunR3KtF4xWmxtmEXpO0SOwAudVzVIEvLTYVEYSqpUVBECkV2M+rIpSDcaa1/6I
IXc2mtaMw68jsfCFQdmLBpL4RBcwQBS0zg1NJqsYUuyj8XNAgwsXN87+ex8STQAw
WZyMbGl/ap2kr3gCfFbiC85tzRaDwG4JEZfdiKoA3fM8RVl6rdlRf6UkMLFhZPkd
wEB3JWENl8ukJgnlrrjnNQon4lQSPg6q2LU1N00szIooTrW7PKRER9VQhXjWrAny
SM2w+ikD1K+eESi8Y0BepFnLJsq+lqH4qfbzE3nj49LZ97265+gN5eTj+KPHxg3f
zZPHpLJ0KquvUSEZ8BM4pZUnuuP0PAsP8sFK9uS29LpU0wDmUtBHNc1hCs2xaI1+
ltvU05yjexwJ0Ar6sGFJInUy5c0mT91rs8pgV+rfE75Jn4blHV3+e1f3uvvxSuHT
+i12YXQLgjnx/x3lTnytmgN0bvmSmYybw4Orf914AZGP7xGnwkG4y+dZDSUH4ucl
kxZ15lOibuHNLfqIZElsmpLZ6n+kYtlM33fNh6FyPuKeEE/NP5amIoaIOkyoJ0rP
J+uT5i4jD7Fy0ftmHg5oATg5YWN7rxAf7dF+TlQWEoneWf9xN4Ea+QEz3UOK4m30
Bh23k1Pgjt4XHnrrHLUzNoU/CruVZYPf2EydkBlo4xbk9WOT3mnZ+9elPIDd591y
XAFTMJ+nlL8F9V1gC8VFzTz08pvdmXsrTDiRRGpSRurCddDu/ITn79Z/dVVKvNKa
cjD72/DPjEww5KIbijaGU67yl8t4P8ga4nsfAy/d4XzZSrgo50Ohy9mDqS3fBK9J
klQLp5N+UkfWuArbPjXKE0qWTb2KuVJpvLk8B5VQesj8l0WySNHftiw/ugRQ/BtJ
HWLTnYGaXb09kumTojvfASWpQy9TU8vCGeSMhL1hI/ftUcFq6WLIc+8n5CN8D087
FmUrVbipqmemqf+wwKeqfD+zvO/NuY8X5fBvs2kqrwqEt/fyrHvBRTEVM5cd/JI5
n8eIGGepgv0/wzrF4KIaItALBo3STQXzADSAN0XtjyAA5WAIzIK/H1o+TDNRHZr5
qW7KiItDC1Xam1V5v28NGo0BI4775JKbE5aWmp2dBuYQQ/g4OGVZ3j1+sKeZqn06
WdcS131TvEY6aXTybywEbkBGAKvxTEPDldcw32LP1WL9UMQho6iFDtdAKFq+25y7
V9oJWl4M7bmbRud59LlJ1QqVjBbE3QNAkL6Aywa2YBYYD/qNRMfA2ZGVcQ6nx4N1
QbXMAiqExYCbDc5mN/VkV4k8TMtxDXq0YscgfjkdBIzHyW0vq7dnh4kgHxQMtL2U
DkzEA7DFCI4O36cTkM8PclEADFtyVqssL+hmXBE8tg6xNOuasx23DNixEUEM8Ouq
HK2ENMwfYyVuCXcH8roxewMLIWAiEeZ8xN7/NMXwAdjSTIYv0UnT1PMvNTiHQJUI
UUn/NK3qjKllg/3w+O2jcaueo6zs4tQ0OivzgBop7emW9WBcdnRjUMLpPoh3ht8F
cfA+UZLA64vJj7vW+CexirjRKRpj1AdJj1OTGp7qb3AtNOG+EYCrbbITy/xpMSXR
zmvVCQi7gztsM0FBujaNFbp+41LIw3MJs7OmDZfQ3vh3f87LUaGaNdL0C15SFPGT
Zogvir2bIPZDFZ0BJ/SDlEXGa881nJSIvXgClGXR5pY/2srtla47hOap4xrDn4y2
sHXIJnz6LSKiXEUtUCObOLT4SbWx3N37kKM5e7ivh1U8RiJq/WHVGzy9rTcvXp5O
RzeJ0qo1xacyvo9E+5Sm7t3THjD9GSsyxNJZlWTcFVwcBMxFSrjhcEG8sGwCpRvc
qPFZtiF8/ZQQDODKaVK/houzGM1Xia+eGLeBOotmXIU2vYEV4PicxrbTEXBShbOD
9gjcHhYnmzfRIY6fJYdkGFcI+idwAcQxGYBmyFlSAFC3QJ9oRmWDPRQsQGPNQnfO
9OiDl4SPk/Bwuko5MQdYb/eb/s9HRo7uFZe2NIrRyYJWxsDJrAHe6kbmTB9bZ4Qc
4RLjIHPuHzTZc21LD5LyxtDdvisjMoT8h2JOP4wFCz9pRvXnJovrawB83TjxTE2C
j72ccl1jT7aVa5SOT66liFmVEXDlI5bZ0zkD6Hz3BQKBNCdTZBxiOmxjVFp2evB4
M3tu9GbwoIdkrbgryDsf0ChJ+hWOo3ttIRAQi7hdKHmrH/UOuz/L0WEcnlJ19whK
grenIIZhN1WYPKeZdY46UMw7B1b8+lifyIQZA9/I8A6cTPRKG9vtA6O1TDBJ96Lp
bK0noDNS0k73KffEXdY2u86Kg1cXZleeK0mlMNGcEc6T3S00Y0Bf1XH+Kuuz5cSO
QQT6OtQbixdwCyeZjupXUNgMIgHtwj+Ut/6hKaEJp3/RcMZoBE0FsEdcR+gTgr18
CX0XiWimSyRQHWkxynKWmYfpJEt1fBsbsowD+IOWr5V8rDJ+m6F96WIuZiRBdBRH
yghq7e1FvqMFPPyp7gdhB7PXV3gmwZgrqW6PGDe+Mr/dCdyflaPymEgITQ1HB5zE
eS0YwjRxu8ifz1fiB5Rj0xdOnaJ8HDwJNY2UO6gg3jL/OngrAcb6JwBHFV3rnNxE
gOvX1jY6uyi8q7sfS7/SS3iFiH2nRQfZXpO6t1+L4E9OvqFoZY8ZK2CBTOITnExY
67Qa2qqP10g2ZonBZ+FveRAi1Dc9HATYzW+cW0qChRXrz9sms0yEsvWPg8ayVXF/
pBLjeC/lFwVWpVUDMhBA0QtCDWt+9aYncNR7TO9ToawcfKXKSCT/RWLYY1x4NVzp
1OBxNP0aarEg96o/d5sB1GZqEb71XVBHcbkZOME2iR6T8z8WbjJ/yLeXR0n65rmo
pzNnK7zyThh1mQDZ9JPzlpm5EvveuOT1QuGm1zsZL8r4EDrsbux454KagggnYTRC
pC3rDVKLAUBvHlXqsSEdr21dBHoK57GLiDm2UsbbCnisZi3sTEj8d9/KrGkFh8Ng
vur8lM4JUNuuq9v4S9o90lRNZhiTx1ikVeblJgVcALk=
`protect END_PROTECTED
