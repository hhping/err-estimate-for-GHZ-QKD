`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KlKjVyTWRyNTX5B79phAl/sbmqGvn4KrPkA8XtJTdf2G5MrCuxfqniRGY3uHtgZF
1gUOUhmnkHwdwa2Nj+vM7gEOst3jD++bgHCPWWjczSWVajopwh+eNyu8zyOjuNRh
YOGZPde/3jOx2AEuIv0L9qjAxh49v6drDlBWz2XTKRxWz2PsNmVRx5ekvQNqWb8k
Bentcm8CtxNwS+w0EGhZFD2XwrSH+j/2yhhwtifHiCCwCIRCUaKlRmkcq/EiKmw8
t0cqDqvTPZycMNhpdV/npkx7tCsmF0jvnbPzsLUN0MYJuczbw/VDZGkU8ZHJLs6k
luQfQMyqFTcSP43aRWUlEnvLgbuVrbWtRRiJf5lEwz0EiHjKlTmbHqVkrqkbEoIr
sa8GOctHUBCDP46v0jmpee5Dufw0ptxuEynrIPVCjVCARWElW3+6ZnKQ1Wtr6xIE
5yOWjMKEUDQ9g0DMXrvw72AHuAFlj0XhBY/pFcXmqnCeCGI+y7cir/oYpACjyMWV
8a0jgqFaKISxawd4lWQVcSGAB1TyJyMq8FARj3ROq9DvsoRixaoHPXyo3Fo1Wb7Y
ejprA2dJqiv7AJh4NJ2BjeLLYY3kveX2aXLfKca8DMJG4Mt3PYpvhW/qgIHoJevk
GfKeh2IpUUXEgUOedxk7i9o38YG0w9j+itk2pTGLY28=
`protect END_PROTECTED
