`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuVqoeJkowlNew2MlqzzQaCzOsebr4Fk7gidLRtq/3QqWFwbUUCml+UQtT3BAdJT
RUCiemjUrd5QJ0fsehDBmkJblWRRX7l58Us/+sM1pTYSM9OtQMD7WMDKBlJTlRrA
srzllpmWJ7PbyPd36hNhGCvNcgwdnWsXqbeuvANhB8g1tfH87bqgnpRPL1uT8YuP
NxoSCyc+A+9XBZE5lnq/xombyCeeu3YxkXR8r81mVqv1TfSSiGBPyubt1pRvP67w
JJOLRunvzuG9z3I9JGAWQrbv5xKpQQJKz7WAJNq77Ckrdymo8JqB7PrUYVnxTF4p
g3iFc+LENbsSCctxeN47g7HGivDDccGK9o2LUtCYe9WDn0oRBPmQNQcbxF94gZvL
B1GpPQTnFqASZ90JQT/dxN/EgjT18k5tz6mUEG55bdsYyYgHxsBkvDUX9wXg83u+
XCn8DI3XSILzXADmX6a33vOQ7CY6q05Jq7tZEsVq5F3ULLmmSZ7tS8Z20pHnF0k+
slR3vYE9N6/URQSGN2kMYkDAvRuV6TzC7RoeMXYlk96zqPFPvsA5RfnhKBNE7IW0
Al6xoZk62KAS9olGrNbVrUqz7VAbjC076km0MrJlsxoohueSTlYsBN6qNOrjEK2N
10kNzeO21pVnCdOOTa3tUoTUOUra7+anCelr+mYleTgjAO3BH4/YivbcEgTgWqTI
VVK6B4GpYLiqQGa4sCjlHoFURXApoGPMVSrhzxBNUCWazTHZ7M0GIWERSMKJERl1
a3a6hlB9n+4Ts3yYRXVAVWbKA/rc27Ho7D/GbFDSPBvboZ0aXKOVHALahARvOJa6
SVqv37KQK2WgraKOVH2SI4MgUQwfbwVGgiG2WYu2lFuDgQz7QS/K0FMXdogTjfwv
qCJXX2LdoWLvQ55mAWJMprOnxkl24Tf92pBv3Yax2SvSYRTG8u1HJm0kuZHqm9lz
4BR/1rHSgdPcN6pHacQfW92prHY1e8fIpnblKt/jE8xE1QvA4ki82pig2F+iEnS/
ot3zGCwXOIVNE9hM0vngMIPt5gOx2MSEVVbFiwEs7VGsnv7ZIIuCDLuo9r95d+as
WbkC4BHNV25KCk+8UHf8kHhIXeI8K9h3uaHaa2JZ+Xa/HNWaSrsYuCOU7IbPLVNA
z+p7ZUouQbzpETH/OTFttl6SKujJccKTcroHtjV9u+UEbRrjV975K8ZnGJ0WziYy
uN6B6UZMd7lVGj8NK8UQXblaKnEvsTnB1a/umawXA2wgwI0pgOAA6A4dorjj2ap9
sIYHznTXbWJiktTa8brdgAeMKIqEzD8ZBxI9vd4SQ59klsaxXAuxfenIiA8Q9X9U
WN96QrDcdTrPcOHSaFa0GXjDb1GqxGfAsSvqRKSkK4lqwmZVrkNrvKI/pOVuwAJM
tY8YAr0RLjtjQuy7zTp/8ZtSJgseFvdohU7qd3p/6KkTxH8l7CxkKyYl+86D+6ZF
0EvKeG/TACH/V9CXH197KbTH/BibUGVLlDZiz+qYwjTpqCXy/vKv/OahBqyLOIEV
+kLiQn4HaQGltrXRJPjJQZftWznwWo6HWQLyWNFRKjxNpFoECYDRZDrcV7N9MmBI
AhZkFnzeZZqM+SXIajZuf/jlPXKm+EJERHg9v7zwh+0WyoS2azY0LwfSAWyksfn5
`protect END_PROTECTED
