`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11E6Ms7G4y8jLvpHzQ/P92ItwAT8YyHucWx49u9F3UHeBTC5SYgr96DtyAXKzcYh
kXf0vp5qihj+4lYgW+DAsrU75Dq/FiaZZ08RgolG45ZidvD+tcH2V+joTy+2mb/b
h6dfPs2i8Pc284cG05Yk8JD5XBw3atKV9Q4QrytFL126OEq4wIGlIu/JRdKRYByt
k/WIBuz9C8CiCswnGUl88y6Ln2md3NF3ZmTNJfCP2ZU4p2BsKVfqFUXzez8ufwmu
Fm8tHK4A2J/ghYyELsEE4F4gGKk72xK2d3Uv1b9bbJVhJ4onrSMMDiCHBQoTosdO
BAbWEUOYQ1v0a4WLrA/IcfnM6QE/W95Z3iESkyUl02ED/+7VisV2WgY6pM6KWzFs
cLlsszVfw9VR/Kmogv2eIA==
`protect END_PROTECTED
