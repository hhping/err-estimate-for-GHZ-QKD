`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMwggc2exFpwcdto0E9V//eBHzHXarCgACHo4f7MMrJez8oLF5K6JeFmcKwwFBLI
JgSWxh3wKmFY2c4pNaQTeIfK9MI/fieK6aOaGg7/xlQVBdClTjSw3qvAOymK9ucj
uXOSVFxb5X/a7RakyIY9tdRHJ2ZbCOi9lXFgajHZ+D+HhxHYQv09GRUgwIuz/TWK
8EMI4eHOqI4dU6w/AeVUVIXdXlhtb6hyy+sc38qWCdpSN0n6zSD9lTxApc5+Sff3
U39Tq7iPjZFJz6KMOo+RZP/SxNAcvNYwjhhDTlSBz+bWwkebj856+OHK+CIM/UTZ
4DIE32TBtIcfZGgMvDbR+NAm46lkvd2e/co6uAyxubRRFgvCUvKII5mmiXXKVWKA
F2qNyQN3+LvG6ostpWITpzqT8wSSjC/6b3/HmV3y+2bxT1iyVpS1zmhZ0YCeD515
vro7S6FJ9XB1caBPI4cemfdhC7lp4KW/KjPWiIBsIig77EJuTBw+28LJ+NiROUm8
4z3d0UPuFB/0ZiBDIJnTOrOMm7ATm2YJZLWalWlTYzOTMpaAHbFHIgVjeg39Tw2A
NPC0kqBxHfCZPHyJRXkS1j/ffQFtxtJ2u5bC8JxuWNuZnzTQFfg5roJ/lJILwW1e
yOx2c+jR0d1ZU7GoVuaLjQ==
`protect END_PROTECTED
