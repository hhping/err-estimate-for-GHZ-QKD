`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+el/dwDuQ/KYc3yMThVVK7fB3HFgkyTztt+t3t2rm6jcLq9qXcVyPQ+ijHTJX8Q
8/OlVxHeCQQD/wt6hcrh1WcaWaK+mhFvEQRCpTwU6RhLBq+81OoluRQzztxJNK9Y
da07CR8AxDx2BFfcL5aj38Z3xeQps3WTDnfvGeu23agGAvW5BGjicgBqRwrUpA/G
A8AqavuRpQ4byxcoRCPf3rBqKf0QP27acynqImWWb3dVhxUA2RyRuskrWUSIVAoX
6LaJje6UAg6rFEp0gxTL9eRwzUzqh3E4vbAfhnjxJzE1eY7fWJ7FNhL+x35/ui/b
kwzrCJH/FRX3zJInKKMPaB1aPy5xdNNMnjXb2BwdE0INbgrokU7q7oPazjMnBnsQ
fYfimaJqOxFwLLwBVKDsknBZUWjkc8sIbKhkEj+k3wh3riZTDa+21fAot/r9ZCRs
TaFqjukmi86ZoiPmL/6Oi0BjWvttL/QOrLAe2Cc1GUNS7PTCVV0fUbGqbfwKu0hG
NdM38i+jdz49UEmnHY3pdXBXgXdw5pgidhsyCTXjckD8UPukakFgs4Gsefc7/3mF
7zSjDiG3uMgJxlHBQiduAX16rvvjFnmc/DbpeFaOOCQJpVUCVwcrd5cFR8S2ADVr
QzanZ+Q9LhVUZxYlwrSfXytC853NGTyVMRnFOHf03m+flWHLhlQXI492SlW5D3Uw
i64cMxGtrMTBuK59WGGTLXiiFUr1BjCx/kRPiDzIOOewrzL1tGKkZU7igJvqdPv3
ITk1/jEcHNBTjH9vNZWaXEF2QBZ4GoLiBn22uuxy2/1oAl6P+dEmCmSaPco7FanA
woC5amKEwpRLQEfbs32Do2XAnrFy1EKy9TS1fhn13zxEXyDhve8Zu8AukpC+yqKN
tJMoPvf8TUjHIw7rZwcBJ60l0mT07ifeBHojMeb5hDzk9WDPtqbWeFlWAuCj/KcZ
2naVnPK6AB1AEYe/jtVmExgnKLQRGy5cxCuat6ePfPOnR5pgumiwo+Pt0TvgflSE
D9go2KD4qFZUdojCtdxs6HvUKdcF1VJ3fayP+ShaBw/VF9VwkqTEVkxJ2Gl+Uqvy
L8bHVkT3ghw9D4IggLPNuY2J1qxRh9ksJSS+sbGhysB7cR7mojci1+RdLBsaV1FC
nNGP+PBaPKg4eyfBNmxLyhJWeICbvnj+ktyistscSkoJI43H8hyGAACHghg7GPYm
olP/CqseHNfhQfpR9eO8qaBltGajPoNMwHsXWP5PRyeU260ZMlp/QQHk9T0DwsK+
8kJfEWnhGtPOs5/tW3+25Nn/5Hzws4wa7VRFcZsFGQ5oSmu6TgYkY5cvUQPcSXTW
zhb5wJ3K9GdJxeureF74TedPx8GfsSFbyFMQqrVTvL70fEvHHMqOsTIWRA8vEWVv
v0u9gd22A8BbpMg/05H+F4+SACCqkuFgoPGgP+VP1LQ2EJZGrFniQnOwq1ftKzSu
i0did6WtemYCy+KuMbI581CJiqMlGC5LZD4YCXf9zOg=
`protect END_PROTECTED
