`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKdVWCS1LaVKQwUsMiMS4B38TkuI67UAV2Ae6AV6W//VpmZ9RPUeR6c3bQ3jtcga
PeoOxckDcYtgJ2Ratzl4adCC1Xud+4PkBI3ShNYAM7FQuSXJGnX9bUF1eMPh0Gwt
cWJHoDTIcHnRLgatcOEeSXscyzhtdUMBb+mLvYgr4idxZ23ZWuW/kKJb88cCCjgI
Sst5v/3UWNz5aS0XBMJ0WBQNQ6d1BpuGNj0PNmJr6+i/8V2EiD3R95dWJG2R9z8X
yk8zYMBNa2ecfOl+YWCicdGNYTLsKHLzz7cSnPrp3EQ2dVTK6OePrDiISofQKP3f
IuIno5tAz6Odo3czfggNKnUKawS0O1GOS4tHlK/2teR89q32ywYGVhzmjKGShkk/
IlARg4P9cjTvVeZr7flIEduP/2k3zaQcLSqxJQ8OXXI3Y+VVBRDMJGdD9WS44QEw
rR5/DXuUaTPU+10Nm3pSyCRGG3g0OnkGWKq4yA9B/PYa19oUfgsDMSRosFylC/4e
SOeVVv24doVOBLidtTz3pZZo43I5KweyFJqreoCp/WAbHCGqX+b8XSekIwziMKP4
CYuiDiEpVlVgqECG1zls6EO6YpoxvXiU+jh2oudz9W1ZSegNOyv/Y3Bgg9kncaMH
36AhvvBvUZq+vEmeyLI8+H741ynbwRysh2jOdIFf1Y/bHdHaRUz1P4I1dLfVBYro
KpqBPavDgoeU7FugFARGYp398zrwre/2Hw4DmNIf4oWni3pgczJDJv5R0BuSiN/t
9SF3X86rYfNtv0JlJO25iaNOJOUUR1+n19xTxW2bHRzCOM4U2xqFP+5ibwnkEyUG
f4qNAvFg8qthZHALy1DfmoKjiJxo+/5QBOR0uJ1UkslQDlrd7plGX+0Y8QCTDOqr
F+gw95ZroskNimREVYuBeDEfxry7xy2OSYjYTcnOJVtLnwBosiRgO2kQq/71NmJ4
TdNakiQYQOhL3qvGEKjIJW8llgTspksbqhAkHil/P5Tot9CeUeIqs9uC0c+WcBtO
VSrJqBy5JkCqJtyJc94mm9JzOdss5Jv2xgfl/mR/jCApDWQlSIFALhSExLJTsP+i
zck+h8L3nw8zA1dcZXwk6O96hLqrPejSfF1OsOJDSvUazzeB56mJCFCDie7CYtWc
h14R95Vz8ILp46ndY7KGBNpjy57CLaYAdUomKFuNznBeQwlSg8fTRB2RWmpRMDrQ
g1tD27sE2FPQJWlLwR62LNHiQGuhGGpDD9zu3GM9OW97uQyU/wZ5gbDjnkuEiepJ
`protect END_PROTECTED
