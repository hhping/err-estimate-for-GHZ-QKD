`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qbx+Dhkp7Byf5j5hQV3lIwo88aL0jtf0/m+5jcjqKCZ6v5qHhXTYJU5zr7HMp0Ur
Egv1/1Mp1Pqd6boNzuxW12PP9LHQR08plnxSw0A9ygSRAnV99PEC4iMU7st6i5GA
xKPmGMDOW4RodA9sf5WhjxOeNCIKcqREKZlpPg/i1IpLX59yvw3xpPfVSqxAf9GK
PRuqEHgnuws1HlFAbHzyvdn45c1R43vZ0kl9AH5sHl7ez1cO8tIB7tMcLPoI0PoK
M54MiScCWlBAXQwgj57428oCOFHLAvx24flGIFrFDzVvRiq9D6wE3wdC7HkdXf8L
4H0iT+xqukIeHWN9Paa7sSqFbKKXq6J7voCiEiUbrcj2LFIoDcS/a7qo2SIYSdgm
e4wGVc91XdBlP5/k+T0JBQ8ZExusOHw88ecXGPVDhbQE9byP06zXrTj74KUEV5gm
oeuee9fX5nBNpeGYohDq8tqcrxA+4Eh6m4Vtu3sFTbo8ap/ReCJwIqi8PE2CAsfe
uf/iT8wKzNyGjVE/pAoK+YJOrMZq0OrL75z+oxLd2/rSiYDRRNjP1wA5ZwBU8GXc
reaa0eekkbE9H6fE3trq30zCZ7SZl7MkIg26qfmwXA2vtWeUq6ahzOC/ezO23tsB
kWw2FXYRSZmopQVkCT++vxHDRDbrAx1O7sDXtmaEBn9gpB7Uexym9nJHPfpeQjGJ
2Wk8tipYV7YjMOjeUEjYsSumnSmjBJjcCauwy/8QlTSi29AXRDPboKgeYgQ1sJFW
YPaZgfz9EUolnEw+OBJo1WRY60fXBuALQgL3LNyxNeeJ2askHBbInZMVcR2s6aOS
9GgVKB7a2Ui6n6Sfz9dnrWYjzfreinTxKTnwUVYh5muYEymRbCxA2+eqlwbgkHu4
p7rOhEOOr6RZcmpVjqIynGnfOowGmVNX/ue8n4I5Q8EwMmWSFDyung2sL45lSWjr
zHS6oXrl2c8QZ4ig+r1z1ECWC3mi51CI2xtdA/k+UkqegmnZvctvLgDk8ZRIosdl
3c/j5HQyo00OsuJsdkugRvS8tw1NyynTmWQCbhrjLd0Mcm2RQPsPPNj7ts9O8ue9
IsdRxlu6C8CN8g+tTznhKb+Xhvdj8NyYbVR1hk0QLAHh+KuBUoLIlfrahPcUlURt
H6AZX2AYpgKuX8LcKcbmARNG/uhbLFJ8y6ojVo437/QNNx7JWU4Ls3cCcxR1IA4A
qDEQKG191kj9yLjDTvA9tvXqPxIQeatM9nr9ME1FlSa41OpFdl08END1wea24fO+
kWbDnG7mAMJqAf/ipEDvm48vRMQuskXXiT+84pbf7HvPASkPmbxpE/BENq3SWR7j
AWmWbu7/r8v4onOUKtQFvnOioCaX6awVJbvATfV5xNSyGhXyGuDAe+txLwrMAOaZ
JQJcfoPx0yAG0m8v+cWmPpTGBGXL0MeEJTV7W3AWkhNKLygZCubM6uVYC12K65aM
DcqkjU9dq8szjllR+BCDlo++9+8e+am/Y2gFBiiDrkTX5Pcoxq2kg/PdUB3WUF/e
DsOGBQYH7JUe1XAKlVPSHxv46AvEhucKXBlrH9TnH4tnYi1xDlub05bSdMWdfeIc
RyrViaQKD5euWcn4rrZur4OcIYmcenzaB2Yj7WI9g9EQfHn71KpPrfvDv8S2o9Ic
B4D8+vXcQO7Qg8m4cx0ZkH8beOP8YzMWNmBPKk3gcTRbIKLMUHFDNFR+D1OtXssq
mFpccvYn47zoN+8QEYaQ6kgiGX1EjK71Fz6/m8Pa7B5N0grxLHm94ENDw+pQS+Wu
QSgDB0w7Retr3aAKhp0/s4+At1EsBzZDof4T4Ht2PrIvsdjrtRVcyhS+hgckVzGV
hjqrur+lI/UKct9UeWuBq6DbhnOEBLUtug3/1Zlmtqrf8zteL45ZK3WvkPDSivfK
IS2gI7JK1FfHVPmTDTP6vGS/lU7evwlZ8kuAgmkLsZoBvhWJVhnYdMEtH/R6Nlha
crRPnBw63TcoTcPDYFhe8P6a35WVyqivJFkSzLLSVAmtU8iCVJ9FyzilLPacTEqy
2c+ME9aOJS7JUX7j6zigyNTYneOmEXWxGYTzPiIMMIrAOdil7f4xGJr8xFNGa/Bu
QX5lp4BiovZMvTNt72BH2JNAgssFhyCAaL12Ioz8TPmvRLQ87/+uzoIqtvEJVTML
niBd3X7Mqf1YSpXYQelRRc1hl7MqFL7XqxPtRsneBnXYOglRuRmpTuzgsG1b7bIj
uHJFrClXzG9AinBRr36zMSII38+CLqtwuiIYp0DcxkXa7EuRdHV4Nj7TLmUfdj7r
ved3GSsjBpxkVlY21hkejb+e3F9yszIIL2QoGWj7t7ZrH10S/Q7iw64PFj2TnUax
w/V7STWAqr+6yj19mi9zw6LnYDMQtckA6satDkGD3/S8O2TcOun7lGAV6s5sWWeI
ZIKIlwvj08fjHY6Q8N2yUOcTIxmC9KTwdVYFG+8LFNfokoUCRgsT/xwCPcuyXwOK
sKMkZkydsVTZ4VKxUa5LQtgr9KbyvUVXxWsMelN9x1MWuqTMHTA0avTw2pqezrJh
1v4Mjpws/HwjVWaXxOFemBc6rrdOX/4YkLOoXoJHW0nkguvTd8msHDmz01mXXDLb
UmxKy7pBLxDRPA9euGQ2x3D3fM92HC3eqxE1pP4QJb7Bsw77Ov5B5RvyVRELSJtu
z3E0JAFxW4OK0n/fTT/igUpQhz+mJJ72sCJv601uf0CYCGGgGBUOKBQBY+ZzaxrX
uITdpeomEHRGBhXgHoPaG8yeJ4wxhQ6x6y37x4ZuKKtz3rmkm3ISrDBJLuzhjYmO
ERSIRvIyD2SAsmNy/ZfDFPVDTcySvP8UT76pTpXMDLrhgKPu+NB8nSseGv3FE/LV
ub1epzZ9JQseaxHRBbh2C0qtIDoNccnXH3mca7RxJPjsrkAkpCuJ4KvKUpTVff5O
98fasLJvtMPYtUZX6zbHx5/a4evIHQX2no88CiVbFQiDrwfZLiQLV86ZLGkblfQ4
a4WtkgHZXlIGzyTGE21BW9xwV4uRWnLMdnNOwqth7GAm3PqAINrBzXH0liU+tajL
PRYq1aGaebcNtReBCY+c3sKREm4+qHq/la4tMZNqsUkgjjGskzTxfmrmlmHv6Sab
4M98cw0EjbHupwComxEvs9mcGeRGAvxPc+fmTfQkJz0csEguEqmI9h4H/T6lwz6c
1dtS24y07JJ2qcaPPvyqIwRKo8E74TPEvdb6ibVj9m35OXljwoS6T/9uNsF3prJy
noUoRby6Da03w+axhlwXWBmKDJffhvUmcM3F0X6J7CTVV3oxYdHqAjOODl73kaxw
DisYunEj8w5RBeI0kIlH2Ag+ZPuXm6FfkoI65+/aKMvz4uD3fgxX0vogHNjtmPP1
scSriSL6lwyV1qW/X1c1NC5Iexc21vFSUCy75l4ZJzZODimHU8hFrKs+XUf5qA57
hXSD09ba30PTDollJ2+BO4aO7LiQzlEcfc90VCS3xbefCZrakp8fWpJpwQY4Z1Sr
5EM/U6BrT2/GuwJv1OrG7BHyBmMMcPsjwTaTK+XSZHgKEzYpPDpSh08x4B8dY+sp
1dZsb3bSEZb8BQwoCKdHHM6mbeDzAIRd5RbbCKbU1aGgBOMX7+3K3Et23bApLql6
HNP9gZce8Ca8s7fnIPIR4SVOIGoNTQnL4i5q/oFILl2lnrzZDAw+tD+gYFc45e90
kY+8OVCTCjIvmxIyXOyf5njGY8kASXGoqZCvltRRiBmbb/cosNp7B+rQ/ZpwoJEA
z1VV0HqOrPC9q5+W8hBjCtWTbHsyQLeiRnGV9y2X89+y5WDOhM1nYH7/3m2Mwegv
n2UOCl2jL93XaHTkJKfJZGoXFhO4k4QJWQJMAaUgVSJ+ns05nDk3dEp0ZPVtgPe/
RlUP8EARSDZEkFVnkxWsy95QdjhqKTi2UpULqS+/DiD3GhygYHqaof4HYpAywtRN
T7V2XLTRF0gi0HAmK+AQyGbOmNX3tsWdg6c+GgGI6o8aFZ+cvW/qFnrEbTptFxHI
Uzd0u/4DJ8xt+aDOoMEE1hCS3e80ZQYz+8LFI1M6+DPHY95FkLUGTOx3DDGZ/xjg
QKBGyhOLzG4oE4UCLxlHMudk/6ocmJEJ/t0Ibd37cjGGHptqtakL3wACH/zAkfmJ
RD6RHYcnyjWCjK3TOT9xSQ7ieVQPRZpkc3Qa68673gQEETEvfiGzPQ+SWNvMQ4py
rr1eEEEimpwVvrHEliWq51KcuUUr+q1Krhj0Fh5o8uaLOu3XYfxzwPvWv9RP7wZx
kmLzopz2uV42o77nZMHsmg8V9l1s5xOKO+Pue4xkSNEHTZAiwlSIvcMjdCH2wxlc
9Mt/bnPFFHmJjgs014d2fE8CB5HkS2mznDDZJvaSI5HqHDsg8j1ITLgLeBESHhGj
/YI+A/82RhvZhSzVlIfwVEl38usQ/WmTr4tebUiljghs0wEdO+knZgePN4D+eFL5
VCBHNpz2rp/kkY4uMnxGO8wNufvJeUsxH/zPHOr3l0xRqX9l6vmnYXhUsUJXwwAy
ZVcZ5c36rOzjFrlVCyWmd/u6tJmSlC3BAUeSMgLTe3VWFF7mCfbmX2GYUUThfr5n
0UPJyvGy7/fkUbYWYcbExBnxpis5YwRwmIZzR9vrGGSfOSx8dMchTMgB66ne+uj8
5GjoVxY/I13NkiODUfpeBiPQOSmfWwIUkK5RHGBkNuVvil+at21+KpdTaG6JRoqe
320iR+FxQt0Kl1bCMzh6SgPfHrjei5KmWJN4L7xs/J+Hd5N4os2ugIsrOmd00jOS
Ft0jrIhnXn1euQvEXu8EXFDt+3tIS5UbsDZYsWwedeJ6dmQ8kd8sJu6ol3KmAXf3
svW1ASX4GTmM9dK4jrx4e74P8u/Xmz5dt9RqJgsh2jTqfVrOMulCmzZoeGNvdPbI
axjQvj6alA5uBNXsmrMImzY5YVanlVjA2Yb7PItEUn5L7P9dNUelArerJRJyYQj1
8Kkde5KVaIeQx3DWz0Y48OEqYj8FNHuwzyTmpCb+JYxSPSbKP4uYj95Te/G1Yw5p
tuXrryx5KberjrXxM62T7bCcw90jYdWa93XqRasgQubcPYkBWuHdF61uR8JGtzM8
A7H2dKOR7VMWtFfKwos3yD7NBNc1Joe9F2j1S19/4alxslLWWxcQKTWc8Bvujicx
zfXOpYaNSZJI19BUKdxxhAImi/ueQO/HKgjEMvljWa32rusbAeE2gzmnvLJ8Gf+7
NUvp+iM1w/RTCJDt5dc/H0jcZqR7rsPqCZO05Dq1KRO4DxfyGHXGhdRsjGhwdOAZ
YowPhF5UfJNiftsuDSOh4CqZHgq+1r5rpKL+WAvrBgCeVM5FAlyTo20LZg9zeEjt
JtB3tQi1TDTL4DejWPh8zlrJnoXKxMauYde+v/pQvWnAsTmPeEt00m35pRYbAsMo
P/l+KyDaDkq43PcUUcHNYgBOxfr2VUfqWBtCN4t1YF7Ra5V+QswTsjujaybrdSBF
78v/DN6x4Hq5746sy7VoM4NKnlff0eycsgHtuOcb2iPTXGIH9KCQZ0afDEz7uCuu
5NnjgzlTvEZ3ZymWJBilAJwhng437lTjD+5t/G6iPmt4sbMmXGvXngYNt7GUlI6S
hD24fxiVSbbOEbPpYbewKUEcE4Z/qL1aGp4CsGgurSytW3wOF4eNjvYeBe1zADI7
NTXGoQrAY/4Df4DBAoJoY26JP+zE4IBfnPVv3yK3iBnsNOnCd7vGYLLl/d43YKnv
misXhkc5Y2JXVanhCxnDuiU+sAASM2RT4ZwsClUf9Fp6XlCYOVk8FxJAlIFbko+8
k9qYVzGcb5weWneFAOOek1hiT4aUj/Wm2renrgw+09XuuqulIR2aZK2Rj2czp5jh
O810nNF1swXH/wTpScSyhnEkVMLI7R9rI0wWpaxbsV7gWeX4yxbqEIyBdPAojkEv
QGmpq4HPQPtKoz2kntvrefjobhzWV8lkPOTX9MzuDBhPJgvNFFuXvoMLw5kCXnj8
y9SpVS0eZQ8MtGQkhN14UfhrBgyc7C1d9E/FZQGvwxX9rFhcDLn+sZbPIzlu9uBW
AXquxSb5ketKsVrI6hZxXw==
`protect END_PROTECTED
