`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2AvQywGYMYrhdX1m2vovMEvYr7PL+wi79rDmldK+LNYR3fne2tuidkkePzGn92S4
gs3cI1viuI3NJsH+SIk8QBR6hxLb7S0dWmxzo/mKT5qlZS7ToKs9wwFXip3vFcQW
OJFVJ1qAAq/uwDQrvggvvvwQEG2RKt0Y7VYQk2Wz9ZSC9mguitX0geY/nC+h+G28
bYx1xKadXYuT5SvWfHSHBIbjZ3eehtJnQ+Foi23xgKvRC3U5ECdFWaQgIk0LQALf
sJfeV4Om4PiorprllGWXBZrmt7sILTSAMSTuq7uQYTxo00jya/d0lt3W6KPj4X5w
nHUllUjnxh8CwY7RfqLIuNl1FDqKD7RMPYGDm2k5y+y9AJTLq8HWRnqpDtGAF1JI
0VePzlbhAucoitx/THUpFFNl6bIM1K6nWOWu3WaxB+XhO5n/rR4qtq6dFw4ovW4v
gFWfJ8CnKRqZlKAJyiTEjSSBiiMkY6yKCxLvC2x0YoWtQ8m+6WjH7+6MogFjHEos
jLO/izYM/jrY/j5Zr2K4iI0N4j3eFT3hmwL6+OosY4DBJv20wxI5FIDNeJfQqfJO
KUNxmQfxBmX/82dAeezs0oyBiRuxC7eMmbOsWRAAfWclOY9fTw7T9KvePPHsGOP2
2wfafE4kBMoY8x65uR/x944MW9YR7Zvh9QIasD0dQyJPe7rPB7zHWaQqUulTrlbb
w4NSh+K5Pkou2vRT+dvDlPgQK3sgTK0kEO0S5RyUMACrAvP5Jhnqr1xxKiemM62p
RLXYNIJkxHV+ZjuFAa8sSFRPcB8eeZWDEVnDqP2/rDoAVZj8yl0fCpPdyxNKTn1w
43KcuAm/nGPCD4m1TVrfUYgYM+lo2DWT1wNDrpiTIsJXYXC4rh4oefkn7ZWoBEVS
k2bbWxbBsOWSzUJ9X4d/S3bVVOEVb5oYHddS5XcTWzloiPO2rQnqDlUX01VDMjF2
qG9hfQd6kD25EZlxBaQqIlZHYkSJSuWdWL/dKVRLgZyZag4iGFdEUMgJjkOaBasl
pqtJOXiBqs3Sd/t8crXrn5VJn7N9G5oVPVa73YKb21bnjgWfmA3hNMe8zmE/CVAv
JWcbpPqxjFS607T4axiJcFg+Q9GZ1YORKHZHKkNtVukbg4sUjGl0H0DZyRoKXDBY
m+f4ygcdY5JBWSE5tBqOKZumAiqUeEHJ00s7Qql6f8BwEe7zy/kBg4G8LdfWTRtL
qX4B5bDj9WkQGhWHLjstK78wmvDj3EH+sL81sr0rBAhdvvJrNJZCGqTG5lHoKIGv
d/72xwQSLKNcViuSr2jKepQCrLrvrlJY0YLkxqOo0Pej6XiEym+c2GFN48KKr9sy
hdVyjn6VyUAhggPDdGEKLqMOREPSMsANYSdL0Qu9vIWFJmPMAnSiygw4kJH0tqO9
nHPovwJCSXtMeljePA8ub/N+6kOuqFBiqe1Bw1nBljy94Me+2B1pYKp0/pdXSvku
5kGgUX0FahV9BKD/ZdIQO0Rr1u+j80o5ixDonmBby/jDDmcp073HsV3GmGmxH1+U
G9SjYKUikCPse7IKfDCgyieFbtuhWQthxvG7kNC3vwu/X8jCrv+azvkvOQYa9tws
ySG1EY8mLxzyMCkfKqMDaY0zpPYzpH4ose4q3H3vnNJ8+8OT9kQdhRALO8T8npC3
+CwY+UE7WxI62BwZcbs9FiVKCbW6lJn6lZza7550Q8oSEBQRfG7FkZ8WL7pGJ8pB
oR2CVkFCHSmJuxXWIWXfJtxFNlkQUaE7/dhZH6WJaR/5tWPX2pUPtPQFEbgVtEIv
peGmnI9ay7JLLWYutGlE3PS8KKU/6L+zBQHkpwNpFUcxVUoiPdtJ3GjfTipxw0SS
A43mP8DDEOgcDL+OKCk7UuVlibk9aKBJzuRgAbmGt0yaR+p+s95yKnDhJa4ROVj9
fKhaLfZF3z3SibbnHe2nHVSZYgPwCHj/UMdJSlLiurivc/HCC/0XIiTCIPe0tSv2
GDK0wjurYMs3OzkUUgRxz1l2Q6mY/v+B8astCcBmo25eeytCcJEBWCxAkVaAq7ko
pA2o2jEUMRorEAk7hEdVKfSDq6B5p5G8+b6FSKZd2HzDJ1wzREUVtikcR2QPvrI+
UFRqu1g2mVHpUYw7lJYyftl+MA4rOxuJd+zRD/feWfcJh4z7WJCJ40NGqyzvKPxx
vWcKtR4qI+F/f36Zna7iG9WaPCZtXtGTaJWRLmuKssuaIKHvrqN9MVNRWWnrRqnN
vcrY5CGWt8fYXbIzS+lqhO4EIQ4z2FFTBzMT8TcxbbzQ72eaiksG1aWq1LRSfuMg
oIZzgcktBR6tfCV0JlOeHs3/U6vSNv1qefIdC3xHto31g9nZbzC4p5/E1CTIj2Px
KivNuIC0j0Ysl21OL5isYvqHSLa5NDICw92ZepOZ5TCA6Y+zqDcUmYO1ImEnkiqi
53SP01D3i+i3d92wT77/QmexlkOBng12AuwGqiAnPoM2dZeUG26nUOA5js6aDEVy
6nvVe8+nuNfmagRg691aFGedhIx3+zFQ/M08oBojEJTZ6LwlSWpTDoosCUw2gNcG
sbWGl6aBysARJyCvnC/JkJGUBW0BmME0QEzzbtVF9kCaKpHvZKF9+0R74IM7/g0X
T4ufn73ui+DqYrfJZBYof7FgicjD3CJkyHtrn2QQe1KWPQcaJV3ZdNDNslpoO7z1
B2abEeKa3n5Lw8BT2oxHgJve10/oQq9Q4EDZPiMayTSucY976RHoyGbQC3QaEZvT
MziKjeJ/EeKCz7yDmjYDfsSOromRffXBfvmUEJPJLzFO1oxo4j1sHfY0lKk9Lv3H
rMjiiI3TT8DY7QLrc3udz+MguMzNgHPjVQY81KPaWb61AMPr0wFLxbuUIaUIJZ8D
vdo+sPY0d/1lIcF5ZAjsNsyorIsBMhkab5+aaXJAscBO3qxfz08CPqa1rRTfcx0J
0Pvpy5mtrdvQGpJrsc2kWPAVpFVWBWyZe/LxsH9EQQa/7S6t3Y2l49rFNE9HPqR4
IrMd6w72dPWXzIwxWEdCmHnHmbbhx3a2FAWaTEU042OERicpWHYpwlMtjXVPoId7
dtYKWF46ygfLotB5sDzuEKNsaK573Ns7cUF5tuPsn1XRhMnVUGMJTRZdeKj88GoC
pju0XL5jUNqZ5SPHUJf4Og16jxa9DzKrRiyXt77wSL2FI/VX/iTdo6yZGJJVDFHh
2eY81Quc80x91K/swD5IohFtaEPxR0ZYlfl1VejIIUi+Y9iRGgNhbHfcjKNuRalH
4Kif/oRvvBPL4tQkT0QEaj0AMOKMBXaJ6/xj+0YT0OuNZCAPoJ/Dww541bllgmJH
bkMoltstv/9iro82CpuvAu6G+wnE5iZFOJUDTjHaztfU0ZQyqIM4HwbPCiIDcnmq
V/inojMYJhLftQxPGMkdXnY0JM/fCAYS5/0ckOqeoBfyEVHJ3EP7OJ/i5Bv/zM57
JFmY5wYWVAEixsC+ZyKdpN58HxSVqZTiSowaMnexhcH9H14aDTMDczsBTNw+52U+
/CAsHctPu6Usoq70WAPB1ix0L5KGwqgt6kRZ3LQ2VV1fzzjfO7hFA1FzAQ1ablaj
nCtZSe8JVOs9Wtmg5OW5j2UfqYLmFYiRu1+hoc0mtHvLrJThB5bID81r3i+JDD9V
xcAvYaj8U8g0NOM2F2eDCplsiGS7ncsCCMDHhbGcIm7vW4HhKUVHgJU7GqZP7p9e
U24xMl8JAr9o140eymp8iixOhMDj/6E+U0ihKI0NgskO87Pz9Pz9+zOYgpAMlWRw
F2FwxA1ux051mcERlzXlTash5NpDKf6r5z+aGvHyGBD7FIz3vzn57Brm5O0Tij4h
shBbHjmQI2Zjhdj9MZqeWaoS3FTJ/ThtO4boKmW/14gZo6GOvRY9YpnX93sBnsTo
NNDH/9bUulNfkvAPOyDXo5FMxuA+Rl3ySFqvS6c8y4SabnrwGhaY+5SyNVmnm6im
9GPmcN9ZZa6m34n52h5CYFDuzOyMBhAG/3SwLdnnwUB8Z6R4aud8MZ/ek7M3Wsfe
vFCTuLD8BWtUnTsQHzNDzZPPzrKRJWswo35fkdfcKV+DRmLG2BzHFOVY/MuR57uD
IwzC1WHx2qSfdt/bTXv3UaWAOCL7XPCVxYkfLGoUjHZKlxnuuaw/db/yMEu4NIaE
UVuL+Zf+NK3uO1XbsoHKXagKVDOreW/9+tDLo3ORwalcDRwHJ4KcqchUeMauo0Pd
e/1LSnaIv39AXx/APTqPWSLT/fIkxlae0jgaDTuvfUmeXuulg1usBSeCBvVfzLot
mLfSWaoeBWW+tkgvF8+YpCtMsDDj7U/WeI8dFxpb2uCZg2GIJJCYQ+jWzzM3lbuH
HZ4Ws0GeyMscQawBinjfrpihKVs0qdK527kqMSOAayW7nnUXDyUXzqx7rGkxq/n4
bHH4oSQ6+I2V8l6cc/R75e+5VT1e5su6U7bKMrXGN61M7HSHCRW2yQNR9b7zqIeD
lMVNqssPOKLiAMz6zHIR/sBrXo3QDVLFQdSgw4yj37kvxroZVOrYEe9ZokW0x1Xl
BrCgn0iC1Ly0lvC12PmrxcxYNsQyaEUxxyv0r+hb+XoESeZbF9dhVLQsKdBV7T9O
yj1KlaNQL7a37D4A/sj+lDi5rpPu5K4Z285UPOVTyOCaO8mJ49rL49fgcZj5Hx5c
KhY03hcy8Pd/83V7LQY8sIUKl2SBUI32sTVOeiv1t1pRj+RI13C8y0RYM5C585PK
OnaUnPvJio1hTNrpiPsn+m8ZYXghsubxlG5hYsCfoP7ivZdXxfFRkRe49ciVgGEU
TtsS+XFas4G232lp6MUrFY/mfp9wNdNb5/SvrTkbUJhiRiN27q19GX6Ju+Dy26pg
Mx7n38L8B5iXrVkM+DCK7O119AxblyuzgWsF+bEJ/Uiqhq/TLPZaRKVBfK6hM4W9
J48OUO4GuUg6SNRNO1SOVmaSwj0IXxUbp3Vo/d8/QxjdsN4taal7a43SRkdoqlm2
a7znKlBVmiSSXgAkj8uuHVCIlkKw2enirdFW5IjN49tj9QJeEDsnoo7c2Ssu5xOF
ipGrYUrUmQQNq4HZ8HxiO+8dZwNC77XsEH7nNhSd/Xg9nAyY1MdxgTVku6yzhh8m
oUYF6kCRh+30sYn4s9YUut5esCYD42dzna6XjrLYE4+H7kixpOn8Lar35xivxiBT
MK3jH85A91dbpqZmJZVwYuCUNoaseIL70rb39iO7tnOxMj7jAtnb5DYeGgwqFq01
y7QhTduRwoZG546/POFQKUACdi8KFvWi6Iz/J+MPlhHgQ4sT65GHY72/cQk55eq/
bGAipEwT3HpAygDSLu6GlHrIRohAKQaHvoosj/oSyZSIuqyO0qq3/u2yqU11Ux5G
txDuaLpldoQpTo8gtW8Oz87fD1+noPKJLR0PlYHG+Sh32dWc/Wqtp+VeCMcuLGX8
JUR6yyrMbde1ZeQJBYH76uumgho+XPoYoemHk+rAmPqW/wUfxq+o4PlKVgox3b/e
8Fp3oVg7sKw7Jv49Gybdt9JxIEmACYMYVEP+0sge7ZQ1/2uT2Oi3tA3Xnhgcho7W
KsyKpk1MjQfeVk9PZRHVNrICoNkT255q5xoT8pgFfpnjEcTqsC/9TCzjsY4aTCi+
ZBLgLr/wqe6ST3L9hpVEqX+OhRYl/ZhLTuFjK8fGbiIxSnWzSxF8Myg5SGJ+c0BL
aqWCNhBXxgKcpaChfDWt9YIU5YjEa36phokKln5YZTpp+9aPMqiKX3Tv9iTnhTtR
dThxhgEwZu2NWN0W3T8yQOdlmpW1N10SS+MuOU4EGbHqmYxqdGoJwrLxKXNza0AY
+k/nO14P6UFPF51mcUsuleFhl6ocLmmFk8jIIJ605mURn5Z7fjGzlteJXP4qE7cX
GB7/XIdfQcQHAFq/UMXX30dWunXPic516c4GyplrVe49MxjmAE6ddRljoTWlJKX5
OwOlq7OFQfsBAo67AClaVPkmanamQo+GgDXjjX0sbV7X4zOcg40Zifro86AINIDP
4+BNg3Ss+9ylZ5rk5ZKUboexyL+QA2/aODVU6osh4t39p+eVo3L3cCFAwTqXToGy
RBFmtNOUeli3cw08JyUGEBcNtmkArFwr+K7AL1bDxwXMc+g4k6aJIbP4NyEOcdpB
1x9wiJjol1QsiTLXII3FwlM/6bDVAikPj4iqRmS1TSZ/sEjUSj99iTAc58Se+gsr
m8phw58oJevi96TmkABVa+VIBlqg9dvvwqBGQCjdl707Rte9ie3BGP8H2rnYozAX
Kr0gQjjVhTZHnw09OTc9CePjefGngArB1xXKymlnCK9esVLVeDvzpxtAyGXe3TR0
Z0lBNsdJspNbFJdTysObaHHF2x8mY5EycX6pMd5xsHAnLqA97irdjmgbG+oAA0Ui
rLLsjtrdWN0zXez3tjxM/CfxrTXE07imSYvIJ7vPEjra+KynlZnHSPymfAFuT1tq
mIzEioGEegM7XwjMpRwGrolXtqbl/vJTH+8u6nJRgM+Tsapy9PfSPRbTdGUgT57s
a4NX+Rr1my/d+EDqAQMJ4wI4tonN/XlM34Ne1ve6Nr3KtpEI0j3oLh4D4taqjV63
dLbLXV644QPZCkVEgp+ds5dBJLYihzinTpxduV+fj/gF1YTcPCEYizmdfx/fo3LB
5sptCeJKv87rTohvxSnvmCMK+JIvq1+oKCBkzIF8iF6UhTGFHTI+T692Gxxs1DGQ
gPNrDsqs6uyMPWORqGRUGqJ5KudOVyoxDC5QVK9yvoZIeiD4cvHGyt1yCmVw4/En
MlvQVZN0gAliDBQtEmw76EKwm6Gvp5iXNJDDop/zEsiwVwI9tIaXW7jNGcDEUqsM
s6XPjZAPZ/YQjtt81NoC7yq1jDqBZdbw0K+Dh+kSD9HUWfapxY/Ha+dL7wGQPApB
NZCSuljjSDg/g+eIPx/A9Oy4OVcxoYGcf2lxjJkbrm99RcXPyWcafT1gFH3UQ6qN
KdihbxiDJzvllj+uMS2fxwW/yms1fBAP4dnQujNlJtSQMaBLBKcZOf711EAKkVOE
bXHlK2oBVp/u6g6b8Ydir9/jiucmWm6zoIjgTsTTCoJbD64VO6ih7/iCaB7Yk/em
7v8OgVJ6ZzkdWJNgid4LzkbgvR7U1+aenl/RwfuI11J0kAeSaktI+pZv5TjdkJu7
BwROVJmSXVR3k81dH92q8TnHjIn9tptg81M4KGuGwcsAQd8saLBI9WicYrlpnHvb
67Yh8bbGHBSymgMXc572rCbGg1J4FE9uqUHh4xO2DeWYwXmRxI7hcK5zg45UmxrL
N4L/21Z2WKI8WurYgDEYGForYTy5G86a4KwZwoWkc6jCbJiOWMVZnw+tuPMxbikW
pVfpLsVfG4QWkCuXBEaWMZyRIBSYrdDmU+DZBG09yj/InTdK3J5KanUWjJhGvF4a
VcQRxmsKzXJYjeRT24CbIGKZotsM8USvkZ5gJPwcDOLPTtKTMkJHzTgNRoCTeJFi
m0DCNQLgrd23+y93Iv2g88y1uC8n4MvMIvhdgzdT1Po0N9fqeLyD3Zztdp8a3zZ+
lvKMY3OTCYKhIye6/2c9AjD42m45eyAquC0iQMW0NOVSjq1eeoM/NgPshbBfYQ8b
ll9kKtPvrC9LDswbpm84RAYPXEagtSRiAXnpdOpXrfYe6BVx832+D3lL5y5G9rUN
jQaci1w83FHmTu8ZVYq21RtxoWjLlzvCldtUJqdLpkcyaAapbHqs4OgSkDQKYWF9
BLlZ4ABDKDSNizSsBmBH1R2W7rscSLrO/NjKROdkklM4TaROUfhGRW4+dsiHUqM+
QGPsu5/WruPpeP5CjqnA1YxtbAQ7gftCQO0C1sGgvFZnXJrvEOKJi5XuW9mt8jNw
lbxZ2/SZ7DhlwQLhS7AlyOyISLuUFLR3bltBFvDnIwWwsfKGFXmldgAWm/nDQvMu
ZC8FCPWSMzZgQFvjxXta8eAjyo0F4tCbh3bMU4DiYkXvIrvHZ4YM8H9MFwolIM+3
jc21m5/uIeucUO/tRAad5/wkUF3sQRHOPq2I/5jnipUL2WbLSv1CX3cc6UsU1JnC
biEXIYM3MSqkqZCBykT3553F33SbLHW0IPK0IxBubSY9EHZRBM1xT/hKtwXH//fd
R/iiqc0ODJlh518kfJHAaoeDfYD6xcwgmfo1T+33AErQFdku7ux7MNFjmUXWkN85
NqQnBEqXpTYrm5APt+BO87M6FNP12W1bu/CW5dk7R+dfb/KwKKVGZfGaqw2HP1E5
Pm1t2JTbkSlM7OTovzRXLK6UEiXAiVR68LFErU0LBvPv1U5tblXHa5xWcY9nqbex
0xEmQK1b4RYneGeXyBLnMBrmqiZFGEK8UwUrE6LbaJ61KgqAZeXJNl4io27rcXwY
jTWSEiroRzTpHr6L9BTDlJbKmmNYPKNrbsN8zvwGuf1hOAG4RkoRxbQwX0y14s5S
hr7vne3+ua8LxsiWYpzEMLe7YmbSe6EdOL+Wu1HZssNL4KQTarEnCG4YW159LNoS
JoqPnKNlqSzBusGY+dKQ4cB5kWBAbBT//9SDMIYa2oAatXTmB9M1Ygf7mcqzdDNC
l/yJKdNmiRsUwxylWKNHHEZogwKJ1gcG4txl71Uf/S2Q3Hi5qugEqim7oUL3jIx/
JXiGJ2Ax3Cm2uoHCx29SlPKv0FDl/HEJ5rP1C1/3I2ZFivSsTyTDV2ww6+egJftr
w4IjADO8CGfWiMAhyo11UeTuXO/CUPKQZ9lJJtZigufZVWcPfXpEN9HgZP2bO+FK
9xm2KFb/0j/3V7OVNIel1kn79bSfwnbUtu6LzsUBDkKiWQIXWXWzEe8hPC7n5ttI
maM6/3njyETRwptF/HbqHaqFO0DzNLEan5iAWcQa/TVTlDaJ1Yr9lvixMbmp/Pai
6X3zHewDpBdiLUuFlX0LNiQu60qxDTpSy1VyhROsTqvzMQ54pe7aaQpYukCnpg3Z
FqvR6WcuuNEp6k6EplcH0I11kZgOTPb9tcnMpBsuH1kiitopnOoMFty0W73H82Oe
xddPPV8PrBkt4AHzdpUEeDBaNpOph5R2mFHLMR8rEaAP/Y9jRTIpJgZF0rfMHN79
7kvz6GjK7dQebKVIxxDFxYOaZh/7+eC5bBHvZWTr59XxGA1wNauOi29z5v1SnPCa
jyM/UbpJEU6V/Fgig6SWUAc1+BrgX7y9jCbuzbSijQmw2YU2M4Hh37d+Ce/KV0zn
nv75lD5bGwOKpfMWj7sYOL2ljd1rKDpOYXyHrUrytRpk2KoELoX/J0d9fuqPyUTp
oWpLR256QgpeDm63uCZ8EAqynaRP7IRqTgZ+bT4DntjtuYHefNRL40J5kMJK6W7O
07tfb15eS64NFanAygGKYZKYscc6+k8jaw1qKzKUd/gHJ19o2JT8s6zX/wo399O+
rsP0bxCgmlNCjcaPkJUwtO8dabjf3qN5SbdzWMxO6DbIh+4C8xk/wHrZTuulGlsF
nII6mFKewaG4goHW5sbAdWyWj1lOwK885cm3pOawsG0RPE3DHGfRP3q8wVeUdRYD
oPjYgoyNWXA36GrPVe2tYp3Kv/rCf+7Tv2nrwdnOz/pEBP+5lfzYGHB57W/Mm9Q2
fTs5/SQFgi4wpcLIzm6rtIanYd/Krf2YJXaq3hjVNVeZVd8VijB4yja/wtzE0P0P
GWYxz1yGEwhkDmoUFfF1LcNQfIQPl3Pg7OEbEQ2582kQj9B3UOeDscvWkBZH8VaF
4CwDakoH7rrATkvul688b4ndS4rASFx8C63rtL5YN23YlLqCU5SlIfqEM9RLMHXv
g0ssTmuxdYF3raHEknxjOz+uNCf/p4z8U6Pd34VVZgHUUi9GPLKw1fm3m59L4GT2
stAfeZYnQQLeyJM7903fBTcv7YbD/m4psz5ug3Fvs+K0o0CLsLr7KsmHDbQBAb2t
Wc1+Bzc/6tar9mrvjW2oB5kLrWUwN7VuHpSgsY8Ni2tpkSx4VScdcLAubDeuJPQP
r+LakVpCQ4Sqd/3IrUA/rGjrANPCfy5EA6U0ZU9Ubu58UbCXPhZU5cozxYf44Ezh
IHNzr5RMsHr2rMosiHP9xMOCFBSRsRjSYmvHMNyUia+eXxYLUX3L0JwOPQbszoIm
vq2/9vJFmAJnQ7xdHXECkBN45IdAPeFl6lISwJPxHH40tymo8MoeUL7CIXs2w3yF
EgmJGlbvOsR/TzBgGEt/XEJQrmYgKoDXPWsvnBBmjMoKH9riZ+hUOELTfS8Tg9it
S66dJsEtCRcQzRvsozIsVvUuwFHR9V8g8qWAf9EVhB+bC82FQqHAMAjUWMterx8A
up4rzqmdHinkNRMF/nAccx976XIrkxmc3uaEmoVAHl/nfR8jyH2AtNsSw577D2ff
1kUjUgWwqHuCT276rZSvNPMyIpO6wxtkIHn2Gzn37MEpfbxQ3O4bF5WK41VqlaH0
lpmsrnAgKpPSa+juuh2OfpmpkXvw+485CJjNeHTMhjOz8/G/OspDmnpsRFzL/0Hd
j/3ICyE2CW3DcJzXBkK0Z4YfjHGReNMu1cQFvr4tLNyChc7cKYyvP7P0DdJH7/wY
CqR3zBgxvSdJyGI06mXN8Fq4rGUeFdvCBG46Nmi2cKT6L/be4KDfR9RLCGNRhU3x
0IYJ9nklNqjE0ziqy8GPJb+X110jMAYZD075nBM4smbHfxmTN4EECtp6VLMgF1QB
8NOJ7QavcStpoNLWwGQ0z7ZIs9v7G3lQuMxpFk3imnvR8KJX/RwozjkU2PvOybuC
EoOMVKZfqcVPMseoPtU8Fot8FTpUNM7uctHNxDZI3U4ZnOclKG5fFUoobUYG6oyU
CeyBjYoK9YsFgTPUJCJyi91/+xD21PVlHN6eKLM9IV2Vi9YRG/UtmR7p6iMkHlUI
qI8WIsCKxoh6ARyzBh5vx1bMhGvoU4Us0ztNjPVMpLk0pinLcr+CmMruVMS2rBYu
bYVR8l5i4dsk1SC95FslTmvnabAQkwx+YTcZ95MUOlQ8cy52UCBrfEy5FAMFadvy
grZjabcoSro5MK2mVrE38h/m/6Wsb9v+BStQKn9v6cMqQ3fEzE7D+fnXANH108Wc
Bj8Jzk2aBgb7kqicqiRTTDaYWjjUZf0Tpx4JE0IHAKyxmOp/JMjhgoDvOCYXmtEm
xr+5CdG4dmHVBUWlsn8jIrCK/6JQeYfMq2RlGQt8Erg7LUz6dOOTRE1FH1eJia69
q5zEDvyjSJy4gnAbJFSY1xRDL3s+vyxikJ/QnYAuTZTuL6aNHx9Ey4ex2lKSqU2H
8ukoZiViDY5rAcDb1spnJQRUYVkTOjrdB/rxqKVY9XFdMHb0JidUz9T3cRjXBfJD
rs95UiU5gPa5OJgTpSymSKiBaoNB2aHmAoAlXHDASdXrILDCvJOsFKadavhVYOxR
KeKJCMEh93ddTQfkbsn08zGfav8heiFahpIPqZYd8hMyWXSoRndvaKbEiZXS0jVb
K6IipFmrgPtKrYnvwNp98Yx4yDLst1iQ3EH9sNT61TUmTLI6aEJgAcg8tSzuYh+J
44yXP3n6mV6SynXcrQ3ZPnpxxLY+QzNieILLgkF7GEqlDGUsGAx7DYfE6i2gdFR+
S0+vlVGvufhneEqk+q7DV/t48mCBi3RenJXgwAf7NhMx3jynJGNC16FlX+sJlqYu
lIEQkMCtGfJJRPik7D3t6CsaBxv0x+Qc8w/HpLzKIPNqE7qPztnc4skB5h8MjTML
5+wUJvbIsni/4qIevZQLuZSpv1tp5ZjjjlLCGorrgeAZ6+Y4+jTfESN5ug6QzV8C
Irce+wfIUkYRmuQ0mFLJ63kZwrFqb+JXj9PD2EYk9caIBEKB7GXY02QQ2Mt1pI1k
mOp0l+n0mXv+ckRHFe0JBNDkmiV9ObTMCBmXWJNO/dsnWHFLzGwD38kDtd4gHfH/
oVbHTz80dJbZrTgJY/kbs1hmmRhuep0LVSuwt+2rgASUD3kCv5PALlB94zwsexqj
QhdBfatR54EKvB4WmIv2fWmBoPnleJxcfUgMadGOucipiTsZURVMwPh9tJGSE/dh
ps7/u5NSReW8+RQhsBGaslFywo8KZ1ivdwJ1APVIP2/uyp1qaKvzmj/LVxCy6PtS
WRinAr6VqAL8U5pyWILnR5zbuQDylsYW/sXprB0FcsOu7wYyIp3QpNxG8d/oeTSi
ymT9daQ9anTf6U8SPXnOaJXsXt3TmO2KlVieLz1AztacUD6suXpjxm62oQNq0PIY
REteUU/xotxX5H113Z7zFL9GBNgPyKSum0k2Qq+Eh/1DQ0Bz6vh563/pj7GOURGH
k2MTDTEDrUb/ceEVkI62Ag5KPSBC6u1q2IAtlNfwJOdqKQbj0ZoeWIcb40IKxWfq
LnD+/ikKjheZPfmF2wfWNZp4kTLUaw6gyWrPwEOdXqHEBRgXXjv+r2XoiGCsJ21D
TJ64mMkHn2PNY6qeq5CbeXHNfEXyv3g5b40RZG/D+SPj76AhmoxmfDLxcDBmTMCt
1Hr9psHVvkl4nrJ7So45kJ4FbiCiXyyjrXO79SH1qtdXjLN9pfQX0Q+OiDm0nLPi
q9bGgmxMMCTUtr4jU9IHci4Qmvm48w5070t2t3dCXjYIbaqT1TlL4fi/tuSC/mZk
g1+tgynWRAkxtGW480zNn9YqtnYmj0s4qhwsFCFEmpKBupbe1ogTB1O/fwz4OKR+
ICiuvbq72QPSwCV14Sqh39LLHDVwRDzZNcIbRQxc3yE30VO/4kxpN54eXMHrKbD3
cZltPPpVLXl8Bb8lpTxwC4QLWQ8vPHf/eFGQy5nkfQXZ5Y7Kvi5hsQLqzNQFLmOr
4t4cwxkoJr5OVb18YfuNviZJ0GecxtcwZjabslU2E06747UJ3wYk3WLjQS5qPQ55
OhSQGT7WoMPUCt/v8IjmGuehdjc4HC7CU5N98lnaN9yRRCPV9aMrhh9cI4aXfiYZ
Iq+pdxyqgqtr3TddYSUOSmNfFY8kGeloZ1QMw+f7y+ugz4lchYk5zdrDS74FDTqS
gLK1xF+tvoNNz0mlGYyT8TAOT+Xhq9tB6KOCz44JXUoQhYv/DcFoDcJe4PpGJDgd
NGyPOv2EquVeOyWkylFSQPT2HpmwUOrmQ9U0byGNSJE8kEV6VF1KOT6L3qmE0qIb
qOUVQ9puYczYWT6/db1lI9MRacrWM+lQuWk+s+risLLBbgixw6tamdgGWDLPZSVa
Y2ojL9KlCQ1GTeX0apK3/aVbPZg77cimYXWSETOZ+dXyiOFuTiFkcern2HTwu8Ba
b8cEswAlPEoazfd4x6bENCWKK9R5I5iiMvPEtLWF4ryLIdsVnNhciDkH1QKDnAVE
2688a+GrUap6ySJZw7ZIHalhv+78sShBF6Dw6XY0D+wVD2SwiXblEQ6gexQ3AbQo
B2RoAtxH8FtiApxOQzVCD09051gVNjvRJxr7Iwbj0KQkbYpJMmYzAd+4UX5euOOf
j7Z4d1+V4TDhGMSGnRsmeUMsft/pYfuzGrxRHbCZ6MOolZUDCSzq1Ug5QKJQGUaJ
qFhkkRBCpQJ1bQ85w1Y4pqJwfkwHkEVerlPj4w/lKLQ6157+zvp1F/22E/rfsqBa
6w9h29bMiiU5YR5iuxlQmIbJNBBQS7o0qC26oQW6MnOa76qyy1mi2Ii9RW7LV4Lx
2/7lJRg8TXzi7gb0JNCXWSelxLf9NDlvMeIQtnaKDMSao0PTBW44jbzF2/TMMHac
3kKQx7Eod8PBMdNuSiEAhW1vyCSZ/d+CHNJSmq5aEvZykrSOQwaoGEoGK1ojNVyb
+it/q+TifafKCE/egTuqb+RxM80vGJk6AtOchIgL9qFlxfHwGI589DApyHJ+w4pV
6wLm7Zed7eYFTfNwd8cArIEuZXoA2Xl5xxym/+0u6qeyCqXJfwIgTYj6oPjk0LWn
l47l/ZSEsLfENBa8laNcR/rciawHITeezXud7BmSgtbLhc8suBJUffJG/0pLm4k/
mvmB4mjKQoNIq04FLtsxxJwS5dvLr+srLMcjGODRorc83nVOjgsy42Z3ZuFjiSk4
+Ovms/IqBcTwVZSp8kxkaT2bq9/Y9TRZ+dXzb4CwzlcG1W7dO9yvlUZ1q30vP44r
ipqOWYUxDuu2BKYfUXl1fFZmGZSBF2rqDmNfMC0Ccch/SRAVSP51m8j3YG1DVwna
rh9euJ4gDjAIpHIg6rCehO7Nnt3EiEwPgsiSFykgxzM1yKf3zUL7Y6dFDfMj5cmr
HB+TD+lIsRGxjwPJOgbrokmet66QjjvU/iJ2Eoq8OwA76mpA4nMb/b0RTvRTm/Os
cnLDoNpcha1wD9UflccUKBBFL2sejwbD905VHX3ZvB1lCbnfK104CGRIEBFbIaYn
pwVP8cB/D/LdgTXC8eSqIBOs+N29iuWVYQkbIvyXc+md+jAVXBu4I/MzsEvG0YTe
GtrorY0hPhm2t4tEoK43TBkveEoV1j4vHSOWskZTptL3XYS1PV0yU446htLavfTk
6uMwgQ/CkwNh+67mC00CCsALidJCNEvLde5jg4HMlC8DQUEx+en5hsMv8V0UgMg+
IVzcHK5R8Aj+Q4qLRbnJjD3iei2muut4nDz6nhAL65FAFVRRDZxYzdp5dKU5pG1n
bWyXGtg6coCuJSUKAF5pZEXL9fxOG1oMSz+Rbtid7/zbJ4yoO7nfwxErBKabsI8q
9+FIlMdbP4ilITgVZMYGkHe+HvRF4w7Jhd0Od1kwlapk5rnMuHloGgy4WwmSQdmU
XY/Qhhbnsytg2CyyDLWTzRuo2SqCUrs8VXpeIpuYb64p2JAquKYV3lcyls4R86FC
di2GlUS/5Gl7Br5WCQxYJTpV1hFQRSrPrn4XIRLcZkCNBv1kNlBBo73c22yME7pf
Zz0e278fTeFfqmM7t7rBP5NX2121FKU7EMaxjMF3CvgIO+PiOQSEom/9JlEsgX2w
o/0KuiajQVg0gcI5k3/wHydePlg9ePsiH2+LIA1m3XDImik7OiG00uq1vJp5CCWJ
UxWRJBRw59MCaTbQsFpVlDq2WV4jRitUJuayFYzSRXdcHv7PA5TOfqaR/cJ81IHJ
URxC64GHSzJOyXcE9e2EdL1IoHeMAoNVtuhqQEhiXfVUJ9Ot5Q1hq1w2sTS/3xfe
OlioITcUOLapMe6T0jcitJuKMR32FSkNOt4pSsED+NRd/6TAlMSJ5OLqpdz8nZ9M
xWtjw++xoPRYIRZq6Pv/kYQGUkm0ciSyJguiVQvc/IXkX1glKEqrW++1TkEBh2X2
ZlSFzsHl8XzH46UK6GnVHumuLp7W6XO9LhvzCcXFwbmJKh6g4YyAB9g8DUQpHW3m
HO0VwgnUJLmvcjYff6c1wX6FDycSULCncURzewGWyyxqG9XXBbfxwKEKehL0Qf8F
Of2usXZWvYol8pIbysiVU9Y2/jtOMtzXBBV+xry0Ws2/aCr1cmZs1riwVkEPLgLv
65Dw+Uad7bcdqiNo2yXK/KfaGEyZTOdT7HofCG0db7A/EVbLBRvHoaTsNFAXkOUr
iBP+MEmjw1VfJT3JlQbAUMpC8QSEZ8B78zTjNb0Ji3Ze/DA9Xu4cSWaURNnFZY2q
gaaMW9pTjhy9+E8RP1b/78SxLDr7I8rMKgn3Tc7aDYy+/s1rDS9ALpKdKFApDeow
6UWHxOI+tlaPpoJuYW5EtlMaxqwp/LEx+qg0T3MrKvx/WajGYl/U8wEZGRVJyC8T
0OECUTFH4XtRfrbUjQzOVXstp6WvL7AcgAaLWZct20b5LJB2+HDWdpuon3h5FGMl
9t/gAk8fvnQQ3oB/ih4ldnOGRp4cILAmegU9CMiVJ6Ezjh8qZDYwFr4+eC8YNz3u
fr6sDfSDUF1139hscR9x0JMmFFPrCVRj43Lg4+UinJNEkFqH6kgv97I/d2nJY5sI
Qygy2oI55ZkIjRw3Ei0hzX/6PWZNus68sB9p17H6IZk9Dq3RS977600R97ushIv+
3DKL9JyrZSZv0lA8TtUygbyQsHtif/7d7lsDbDUivHL6hCW3r/Tjz4vVXUV1qNWw
lrYAc/aUGOl1/u1NnmrwnxpG3m95OL2MDKJ2ozyJKjwOtALcwpXiKshVUzEXyKOF
1/4dCQzbUWZRu3Y9bDJubmOa3VxJcKEV/F7GuVyvgNB50GNz2ynBh43R2RRNBY0B
tHxtRBxjn6Re51QnT6Jsw9scyUUDgv1+UgELTp0WxELVBgp3jzOTKhmtatAl/fQa
0CLwBrGZFjH6FtQxmovczzR1GL4MBlUqCrdaM7KrHpqcX+oK70iRVnnx2v2QA9L4
nROT+lT0OvqMkWBsQbgoSbBpHnP5GTE4uX3tPfmLcTG12Rvd/Wxc1lhA0cnD2SMA
V5QK4vzubavN8IENVMRiRHB+p12Ai38EpBmZpsX+uOyJO8pfBmkXQosW5pR0owjl
KGhKIqU/7zN7JRE+Eh8oiHde3VMuDYT0y6cE74EyWVocglyrDMYXxh767w/QOXjc
sckP6OU7F2fLzBGwSPUGzzjq8PF1FYbLy+OW3Qse9SDe+n20ZvMN1841ZROXM11p
l3Rca9ktkdE8eyNohvUWA5GkeFt86aTiAwPoQCXft7a5sxswZ/JiFGqL5hjOmlZu
9UWLwbxYb/QC2XuFb9wWraAe5LhJ4pYECS32bhlqcKd+9QUz8/0Z6+283FUiuyfm
4JCA7Y5BKBkkFYb2e7BZV8LrmIXTLZCNH998rEbxkd68OMvds5muOosRoKW46JV6
4Ob5qH+8HDXtpqltDCz9gfYbsW4VkGOZZuI4suxHP1WsHhk1fayWNdAnocNGRWiC
i4ApruTcleqKux9SOOvtsyZB97gd0lDLgUlYT7UwnqctDAb6IU7GqO5Spoud4zpx
HdSdV5JTCqEssHVQuXQuAmsTooe8M4Im1X0jN6rdoxQfxButUxwNk/peZ0R15CNP
hCRCBl/udTsRx8yGRYCW9nFZ/K7goCss4lVEKsInh9XDyOeSsRwLYAQlQOr+LWqj
v48NJEDAID89Y2a/zJ70PqBBfl11E+kgiC/6bOYuPfOsOtbzIw1EmAAhZ2GIE2dP
5lrx1Ujn5mdU5gOH85RrS0+91SogyJCkbqRe1MdDpH107p2FeQOLeVdMJSmfhCOk
NNxpUnzZBOgnw/irK9IS1gwT2YS9W/zOgOF+vfm47ioC0ERU7f6HGU0+TTLaiH/j
Zwv8YMzdlL9NISjLAQiwoysct5mjzKHUdNj9yJ/mnFWNcdghRkb98zXEYKSAF7Iw
JQzvwKZWIgL1lHMmJV1zb+Wq9xrBBAKvHD4UUt/YxPEOIDjjCHC2H42oaAVy5wj1
wudJHiSnQjGx5sZnhYZ6JP8X8EVvzu9sRry+wdV2RkmsGuCYnbV49HAxVOVrcMPL
kf8C2dd9FGIgb9balIV80ncopVmHfMZ9R0dzXFBfrBrOXoc56ia3G6OPx25ZIgn9
BKKjX8gYU5jSwrox5MJvboKButvhY4QsPsW20gDj4IjEdqG10FXYK4MnVPXFusf3
ej7u9FXt2v9u91MrjQP6uvmKCZ+gsJqf24BEIA5mzjUEaU9ZGBvtcYKMKO0rYmk1
zsq0Vw5Hu28a3sOomsQnLYAyHyBQEymmJKm5Sm+ZId3a1SR6h6cY5GDLQqiq2ATU
YgPSWnDdJMgPK6/qn2V24oXm4cwAVnwmSHbDCa7ss5D0ymAekIm4KT7WTpHUuuxz
twCjKyxZtoflUuGSg4T4ri3NeItTaGqj83rR1mAsathh6h0Xunw4G0ZTI8H2fPxH
u6jQM9oPTG6vRLhvQXNLw2L1mNQGzjp0HovCcyfeOZqVoIiM9CZy7XIRHQDe7fMs
UXWikIBR/ZKi1XfMuW2PMcOK7aq9XYb2Veg/3KkjoCTNG86PHn29Y0Wk9o6BQiI2
IejfxdEwHTzc3swZCoxyrSrDCAg3MzxaXm8YdKK8eUc5QOspRN8sczCrRApv7Aql
oDyysxv1KFUFVauEATJy2zrGv68IgVUUxCE5pt4urSGJmMTtOnKh8iAqbFJkCGmd
sBbFIAyU1JoRIgcI6b+fMJV7v/Yt7rmJmTZBwh8mwerV4seI1fTqMG9N4Ptq2KAl
W9CfwWvMBVOKBjC6vyT44E9LpayrsOl2I7OreQ20TwX12vSsRIYCRQ0PNj5gLO35
6DgSlHsMA67e9+dj6n6f7Hzkc6GdSdZdSd/s5XUHqZktraOpmnrqPctXYndx1El/
4ouaN0OWoBDERTx1o0MqdTYsraC1eZ4KxKRPVkIXhgiCiHdTAlzx5XNduSedFEpy
e6L2BPo+n08gTwjteAtZ7A4y9Q4x6Yo+Iptcsg4Qc4rttSrEuoKYV62kUFW/lu7W
cMQX7A2TgZZYhyVev2RUss/FX5dItnQLhXPWZOuq0Dy4GktEVc8/2kRk0vBeOCIC
5HrrS1h7y+Gz8EnTygmj+8nZeG6527rKmNXOkoYrV0ho0uO+1LIB39gM+jPQJrcH
zMnl76ixJuowRBddbViEmIWr8tD+YqP0JdsJzF2Id81g/5koJ1uHbHsPnWvSe04I
4MeWg+uyPIJhF5NzylLpfRfpHSWffXB9zCb2Sn/8HaQsa12CyOyGTffP9vYXj/GV
TWxpGVRW9vd/78YHdOXPaCLuacnPbSpsrdcMzFfOuW9YqUH4bmRtTbIhB1pFGUsj
lD3+XMiPiZg4kt3aAm1dDC7CektY+TF2CEWTgQraAAr+iv4bCnphJbWmk1UtE/jX
Y95BgFSmsLIkv0mQuZWyep3RiXCJZG7YWfLLBPA6HQtiojbBHx4x3+7PkkRACLl1
J4RmXYOzrQapm5f8YryFxkHONq22o3CV7oNoWD6eGo03uTx6FoGqnlZ9DMSEoUtE
fM3W+8VUy6Y1TKCqFhYAcVVffOwy2geVPjUX6DpdWfaPz61GiFjCZ3r1DNAQ1GYs
ha1VnKg/h9gzfPrDc+C0ramZTBZk4SMpuBoybqZBISW9Z7QLvjIKLxBg9g6A/8NG
O+FwJ7EBikCZ6SAqx3xNq0JhuuGPec8bofwVELArxw5khqG3jKVMP+aQqN/H0djH
nxjef0rM4KMIi5tLrznraY4Gw0ta5RYceY8zhcgoJ75zQLEIbDSR7gutw4XINw3G
+l4lduuBcfqgNbex22NUTyJKfeAyXJKW1ZF/r0um4g9qC3X02B1I2dnDReOo7YqU
rH6he4wM/KcF3zEWO2pFO6CAlWjl3lFY/GFsARgfkEOWFB269zJ3CZI/wmeN8U16
vwQWv3YXGJOfLY9ViNjbtcvBuMZJBsqCES4spgMq0bs2niwdyTRKjk0L7hloePXL
WCKLe4zAtj3fvkWhI00V1dTLMf+eHwVqBKn0hWWh8NCdVgX36N57ZyUg6BnVQm2C
h/z3+/7zMdMi1m3Fb7iyB3Sa8z9ZSDIdkUpzk/GLBv8nkmd+lQwIeDPgNzauu6wJ
utVxTCU/X3s1ygEVilCl9gx0H03R4DB5e85CrCzwxqvYX0YJe3oeoBqf8D3j9q9f
4GeF7zSQeDTDGHsEf1f+zJ/BGfuIaoSrMBQemSsxscJw4TPvVfEAfUtikkCJDUQG
gkBYqfZ/VDudtROZ2BTbP0afyfJ8NrRxCBhT5dq0K+twJ60hyNgEb2GyB0TsKkmf
QF9IlzElyderqBgw4BG3Ag9/e3iz26CPYlucHfRVUpomG/SIbOp5m91ESP6I+6RU
f/DEoRL5S/BbFtt/QNgTvUVZplymZRJE29Y7F9E1LUU+TfSlbfDsa7/eUvEGrm7J
BWEBPSzvEIVoixqf+GxOE+4GDhGPn4W5MZ4UcXwhTM8QmvczYYU9Ht5ksi46EicS
eXKKWeOzFaHWoUOL7ChRx43FohpP4cJ4q0ojIO7vQ+VFv1GG7q461/ie2B95DGoi
hMT7o9OCHXXdxNWEcmEIeeBgsm86a2J0A/ZTYzkVyqQvctAOzMghPFAU0OmFd0jZ
1duBQ7qaCXllmhn2Ro9M1i/M/eOQ4q/O/FXc88Lc848bBtM4faI8yqpXu2X5ZVOZ
vmChbJ/n1kyj/C5krke/kU4x+YiOqe/zurihuezKOG/UR2HzhbPlQQ/EMoBvPrS9
YXwFcEEJ8ig45PBMuil/9zrlYVjmQzPJr6YHsI+61LNjLGKZsbEQ4L+5lQKgk0wz
2FuW1k3iQbRJIAOnDH7qGqT0vOaSyH/hW6dYGB3PdKalb/wpX093y3N/gkEEm0Ne
SkRsAM3eX5SCifw7V617FiQfpL4hwnV6M3kK5S1g43NLrKNrvvPu1BHqGBmEnpfq
Pg3amtCTXB6jlV8RlipPUJb2eg48WqlUDLfswzdu9K9OtW920AI5oUVtOcx2o29n
n6D3IyHbPcsiDXqIT/yRBCIRAYtShilD8n7ek8Faa90L7kZe2HrxHsV54XUJjn0u
aJ9b9ljy6AYgpnf+Jfu/QyfwE26hhhtX8V+JSaP83bXyi0uO0dxnkFqYAG5OwFUY
9Mvp9299E6yjDYFW4hwhnAKCDHlIAB4OlHRH0CKsaV62f9+TcBFFOGppunJgXbx+
4t0VGLJhelrmzR/sr7ZpqEws+AntXHxM05FZMDDIYr5hv6a4eqZm4jcASzRsDwn7
A1oq9Bg4fiFS91M1KhOlt7GlPTzfTg+bljJ5NNaxkvKZ9+qet419figmjBX8+vo4
okl56jULY1fvb2l+zZK4Iem+DZxc2hBvRVsQ8UxFVAYXTg+rrE88ttNdrEQkJSsP
3758UuuEomI1o+dCZjqOrNJoiCP6HxWvdat0hIko1yQsGe/n4zPx+tzNO2TDB4Hm
nfS+tlA1WJXiNrD0XJxCiw64ImNGkbEcNW9/YFpW920aCrOf/pG1tJJdIgkMzgvP
lEmkDP8v8/t7r24bA6TvSNMHBbM3WqQ+q2Z6hHEED6Hb2V3ii22MafhF5hJ9lwKP
s4hG5igY8or71UjZxW+LYNWM7UoX4Yb5bOqXjZ6hXcBudHt6uatCAcQNSDpJnwjF
MS66ZgTPDlpzpMqAPWcVgMZJha1L0I1oa8cSLon1QRQvaxBitJNx6t//L7CCBGRc
mjaoWSHbV0Xgq41oyVltgCX3I3eAsR45gZf/RAv9TfE5kLDFguwAgXvWZtK4umwL
WnRfRRs2kQ9GdOraaosNnwcuVhH7LgaAX2lpP1azDsNhxrtZBeIuzw2kdFs/WJz9
LHc/whi7r9G3T9MO4LqI7nB5KxJkSPRQnDaTzvhOfWyrchYLjGt3+Tc6rETHeFzr
zZAC0Vj1TlRH5jrJWSc177EsgMGSStAI/1U0loxvdvmuhBRrtA9vfR4ALs8Gv89R
ZrKEuwV0H87qFoSrzXuAn2M97UDRINUlDSSD7lx3Ji6OrhJVE1OOHeULH9ifUuzu
tKolhJ+XVCOEQOr0n5OTM5TlyR6B5QYoixwlRfBTPM6JrRj3S+LKfDZn+CgGJfx3
lyBeLGJIuM2WKBoY1z3e2+zjwHBgWo9pNLN2hONauuf5hN9vp/PUnyCby6UVgDEn
2SB1wzRzQm/9ni70Q9mg3OtcVPJLYum36qvc380rvFmbKSa3YlIA03jXXv5ExZ3N
jKjnsUQZ3S2sVlQW/oN3Uc8QLxpXTRphIPiqUSGe9//molLF0W36IOPjs5RrVRB1
8JHahAhtCB8jMTge73FbN/0eAPbOVDBaw7T2uvuGXJacXLbGjoSmd2OL9s+dzolQ
ZvReGmCfymDESrI6xD7/yTQioUsKbG6Z8ERt7Zs4OZtpzELDyY4j1YbQFdgxCRWk
jV6sA/9FFQI4z+Yy6rD9mYfqaoyaighklqimOPEdG/3pw7ZYmmEnViLqjQEem7NE
O31CkqAoYSKJEW1qYT1iO2M/Np9Rif08xfrGCm0dIeYHLOF+Sg1QSQOBU3cIzHd3
zxOeucxn+gsds/UP3jg81jegniiavH9d3d/IsrQZTRfVR2Th0lxgheL7PfPGHGyH
KrHm8FYU/gQ5D8oshlqqszSLT1FBfqCyiBcXg/Z3fNrvM2w+pqCdElWXR4efkETi
T49+5UzZQud+58gQtcY5RnxlFz0H0hHYTPEwOmddar83QtZcF4eQMGMGjjcucUt8
c5YtyKNdw1CsR/2xFBA8lqk26eet38TXcHdLyr+yTLm68rZoPOMmQhf4RUXQqjMD
vctLCt7zBarDKcbvxMfXADyTad3eUHSslJtwzCJXOsqKwUwM8fJaZ4X8/091pr7W
J5JRkpCkR4okzZfrfAoG/nzxpv3TS090h2CdrNNQNp7Son5F5t6eMDKBi+HSEE8p
eqS6wioy1Smq8yuIfLEtT0QRqoaffX1xzLLmYDtRjkMCNkP17f1H8/mCVVvjcKAB
EUa2IFV/dy03dEmvKMqRuXycWuwmN3e7m5ur2RDpbmYkSHGnU7hCisN9gmSkFbD7
m+1KjMRzPXgN+LUR2lEOP+0adxYGCM6UX+gvuokSLrhsflKXfZGft6zruThCywcS
llACBtLL6O5xywHKoBJQU8qORlaQtTmGvmDfrhAKFs153Jy5QgJMOOT956yu7VIN
+mJE6UuiwfmzD9h3zHL+mw//xC2bEz+SG8JuwSXINQRtlTVhPtpjLnkITBPSH2Kh
wy9YKoHXTbEOvrBUr6sq25mPnw2dIGJcR9OSWlKg3pv69rlPPlkgvnyoF7K5uEFG
ioThClYHs3zmnbkfyrVluiKyjibwr4/5d4zRzDkdKH3/0aRtyofufMtexHmUOLv9
mTO1TTVV6N59Z7g3ZCAh0fxr5TLWhRg8Mp/0g10h9BTr0cNkl7CB7UAbdvhQoaX9
Dh2FjiY/acCT5yMAFzHbg7h0le38xgH7Yu3w7xNugzc126H58uoMds4qIscQjGzn
37jXgxiY7soyeoCqBJlh2+kyBEU/1v0gMizXWElsljqsUDh4OMvFbdrXgdaG2kvd
AS7eQkNUXhIySsI9DvIbyURED+gwUoT3DGD6QtzLpShi01fWAmb1drvT5K/T8MRr
sAarY0FG3kRUAK778ta9nP/pT4vsSVY5FTFFI2jV5WqwxJllQy7kUS0ejxYn8Fn6
+1IHrnKUM9FTrTl1NTJ6uIFNmIq7OpdpOe078Kw6nW6whDsFcuMHX0Zo7pdJ/sS+
tWDwZPh0eCHtU1ZBCgo00EsbdOX8vP1mFTDLlrjycml/ltLO1iPwMmuJeIkGZwNq
47+nJ9PFE+x16WeU+WCuCwFXfLLkUFU/roF1nnHDAcwhUi+fDOwKYW3FDhMmDfez
WW+jOfxILD3k+h+z8TaUoitxQNoPZuQTdcHRSkKB4nby96x/qjuYqlz0hrQUPwAX
o1qXnwF8ZJYWrsjYMzn89L954UEdEISBiec3DEV/XWuyy4sOP4wfmUtVBdZbbEMR
91FHvUv7nuOfcR6cXnQ8YujL/PchGBIPAqEBtXwg+gsdGLbxVEP/uZpd0L4UkeLT
G3dWT3n/yW5zoMvIVN4NrP3Uq6F9F7tL+QcZO8W3Idg8B+4S9/RZ1LTpQ671cmAA
gdA5qKWE+K77GiOwDZUFtWK2prZkFGrRFL1XJsPvCLP1MYEbCHi1obxBzLVw6Rak
5XsRAjHPQQkR0J57va0zaAAFaR6o4ST5yXLTD/lLRQesfc30gGuhi/7lABwKLf5M
+iLyZMBMqBiW6Id2UG9V691wxF10H2VnmfGmUOH/9GCXeccK95JX1vDoXC3FA3dO
B9P4olxYP+j7Som+40zfk32btvAOaahKLt+zKya73fyvH6NNFbjUZrrzzqSrxRVT
AS7VEZ+Zm2IH4yhwOOOCyJWLZwApFy8eJ4uhUGBKvqnFSQWEiLHszvgLY6dw+N/K
bWA7szXe7nGjK0HfKHbjXt9kerkR2FfjR992r59E4BMnUKXg6GjmER0m2VGWebGY
dF1jgOjoNtczDx5IpOizqWuWVgl/mr6fqibzxZoBRCQT8f7s8GpVvnLW7ZWjUJV0
Z4tYj0PmST6ZqRasAkzKliJNmKl0LwD2s58kv76z2DSjIe6jyJtq0R3tYyBqHsQp
NVg/d4Cfj2Ny1k2pNLZq7frHQMB5rMNMmvKl19nlHnC8e5L+GfP1IvI6k0/HyR0h
Fz4oPngdBBzzxyRkxLVlQlmx5cg1bjp+R867Gs1Q24sfrUJNbkPBpAgRAGM+Armu
NMMHVTDI6XzRHBXeY43Dd5HWGntSfYFeDIaXf4Gn9IZGsJW1KFMwD9rnK/O58Yu+
7isAz9ZO7AkwL3lpsABEeIjhIA2naO1qXk7KKy2WCqWZ8/xqIdocC8vGOSkDQVRE
z+brrreQJMylxwPiMdZgb659Y6c1ytQ2YOFsa/FYn0yWZhC/vBOA8QNJXMKXkF5m
CJGbKA49P6O46EYpmcVzC0dNgwTcl3wXR22mRrgkT0qWGh6z9dlhHghVMw/o7BKl
uS+++ZGAltA31pC0dPCg5QYYaBBWJBBzLqB6SyrJRX2CRPH/zGMNVHrUL6JmbO8h
ZihhaduM9X3yGynqhbZ0HAhxA9i4H2/AQGFkMbTPd/nSQcuLKfA9D9QR5kMqa8Uh
AF24uFNAeLKPGEj7wrH7a3XKhW1FV/SUu6czHi49SAUBjg1/jWU1fYgewZZy2N+/
6AHP1q2K4Y//jhDx4xaz9IHg0KSRROK3bjuxMghhCJh3KT8UNAcHf5qKcZ4Evca0
qnUk0weB8lJeWo1GhDqxHbF45QHbRdWtNkiolxmKV2Xk51GExxjdmo1TQ64bgICh
5A6d3ih5Tip/UL8dPawyMhaGdhrYDL7SjTCg/FPyfRwTtonuucb9MP80sQBwmK3b
NTNxf9M0XHnhe+6u/Hq6XehTMAm9nXjnOd110/+cGoiT+EnpepQSZJP7PAqfDJMt
Cs4dWtUwPxOC/P8BZbuvGWRLeZqJymiOdxpJJgo7wpNzoWOWnsopoZVoTJKQ3CyG
mtvEP+ExAVAoHx1goSRvH2rs9H0DDVEOYwRIgjLldYnlf8wqaC6j4vMwHox9rdYe
V8k4Rt4lWcLS45PwQNKLbbjSbm84WbMp8p4du30Kfe0UPMiPLZ1z9ilr+JrJ9/ea
H78A/kryduj8s+0pl1IaOOE0oGgKsy3DpJgel7DQSDvnPP/S9cJBRVUSgAVee33p
0+iXBFTT+QbXz0RO1MNRoYw23dc3Fr/kHB+SxokCs436rj1lS3dxfs9jAMRe/doM
Hbu8HKBOTRNMlh/V6zb2+rYk7/qbqx5zFiAVL52I+xRcNVeLR9wBIPKoiJsZ9N1x
o3rGhgzOVnNy6dPNdm+7GF71rblnnJq5LOeXVGgYKFZfvTDl2y2c/xD7gh1L/cYX
rR3bhBaj0D0hVUychJm+6HzKgH+OucJWepzAatK3jGoH+agDgR7+o0znv9C3N5JE
hPGlSIxBBgwIURr1k8SYaDVcuItodHiot8QmOUIZtPg8ECuaR+yVfkqFGWIrdhev
4nm+yleXUeEqmqC3Wpg0dDmvgUK4oz3m8jmUC26Y6tkW+6zJEqKu30bgjANKdFTp
ZW4P7tjtatQ4aE0oO8aJJNzZqU7ojX0GOlf/G9myDYDtCxHWbe921xif4Yq/ljTf
ppETNGjl5YcEmRfwYepDSXSpLL9WfHDeK0Mpmqjh7BLAauxzhJEpTj4UwKKXuKEv
gn3u+OqMuezpW7qsmB1sxrvb81KBGTnxMdaQ4Hk2miTy0zeMyqa3X+odd9JA1zT1
YdY61pMIYufYRKgC6sxa0vqLPOn1CvgJX73LKEYAEHjGujpksX15rpEKsfdZMMfA
GhqTXswTBENbIpGhODA98S/hUSUxj4zQlCad+gdp81sCZ1YMcAAegYEhkGvdmjuh
mCE785nR3BdwNCY6Y8tL+b1POXBmUFl2yoS/IS1Q0/Gx1YqGl4E0ArZz1QqO/EzY
izPqBGf4/qsNj8WfK92LDFoZ1PeyUwk1hwOXHiRRSk55ok8JBrzXRHq6zwOZZsl3
A2kKhTLmS6SgWjVlXJrm+ps5Il/irwBwGDf5GJtkHTNdV91jrqpwBqgVz2pTNLqi
lcH0X6AHYD3G0xKbT6v1iYNZ/UBn0W2l+OO1aKBetDgLtuAxoZSWAOa0SH3Oq9RZ
/t3tPcgz5cO5qdkjhz2ljXZtQsRYwPRQGy3iukuuUEKI1v837XmDbqAyWffo9ayO
m6sVsp7XUWPdIYHw0wZfhbDQncZ1+IBu1Sy49a1uUsM7O3FFxFfbNY0n982wODCP
GlZuf9nAslTZtLLQyqJeBGSLxt3EnI3chQVtVJQK47CTeSC5MWApdIZQNyxt9we6
JkctzjBkwEGO3VAyH00Ez2WJSF6NleYdpa3YwYZokmwjoTC47fwJh/L4nP1TXLDC
ujyVznib/BgUYhsAkoIWSftEXWlvOa/dMic1mHR9BcwwtSKGoqEfIMvbroqUtJtC
NlA9wgucz1/6q+nPSqmXmQUyMhlcI9EVEHfH4R2dvlnTVplL7h6Y+pUZaAfm9xFT
yPRjh6mA2FwPoSgOTdCyJ9fhAskT0gsVqR9NTqU/HAfz0jzFtFkHbEmPbYWpYq6G
fCUFxpU5//pPF/RFq2z5/EyNJcL6WKGvcpPg9hutA+d+ixBrA1twQmd1hF/I+PNL
CgZ6oCwAdQFSKk0FrtZ02F+o7LN5Y/coVp2UQxMeqIN8USMiJ/EGGehsJrctSH1b
Za8gjlWAPa04h5iE2SCASyNv+ryr78kx69LjjxUkDENmm6GscsUC+ZTISPzGUxP+
1SyHCtjZEaJjsdJyQ03JE9prBA8+7rCXcsuy24eVcnjw62cfoo2NSXcUqhxINRwv
Cg/lwcK/TrIsF58gWxyYKscnQyHrUnYZCRQu3zqd3UVU4Cc/pafq/9dcIQeAxEOk
8XJiJdS+qn2Itu1v8ha49ZfCij7lAM2yKHT2Y2KrJcdxY/48YgXgUFzXixd4EiNc
s4sqDU/QXv7WeQch4QAj1LLdov5UUxlBUG+/fQwzi2L0j2tP1Ue0vT6uFeUymA1p
4Rq1X7wf7D3ymGZ3z2xtk6zXH5bZNWZ/bPdEu5C0IJRRVF3e0xvYJeZdrI+iURY/
NItduHSdebe6GDK6IF3qvayutyWd/A0G1OpU5KNfoTCPBUudQ92X7pAo6zvDf5bn
MTTy+4IWXWqoEfHQYyLLCX6qFUdivUdTtkf+cOhhXuqt37XXypEhF2YemgzadD1b
0D1q1nnoA4Lh2Vsk4fQeunP8mj3br0SdFrusEBxbRfJFuYOjWoMCdrDJ5CCy0Q9t
wB2251JP7j1Y0Lj8JEN3XKKqJnT6f0tEvnS8Jsuzn7iOfK/UYQu2PYxq7xkgJvCZ
ZllTeV/IP6YC9eRM9LULwbyln7KbCb1Wo6j4pdR3VWOEoNaOaWUS1G6rPGpmCp8a
HjVbQo8B3G5vipwjQG6zel1DZfJbo62682rzu7UYtwC1W85oWpMjekcFB3OLdxaW
BZU9mXsI/XkqzaUIFzEFVqZW4N5k8eKnEWUd4cYYUL51p1wiT9un/CTEcjKC+KE4
83MxuD1P67enHs4nZBgQbgVdgvdylx+ruFeRCdBrWraK0OaNHCxN/cm916UTe+Bs
UxX0YAYFZIMAXIrQErH4TUarzqwfOSSZFn9UILSb35mNAOu850m5fjRJwXoqVfWf
VbeJiPoHhgG4yMMrmq+sPz89m5zwL7AxQvo6IrjJXyEYIHQhFsgqG6XGuUMJPtiP
qPAH7C28rGBgKL+BPa7tx1m4gaFu84XZbFSOHveIHaPnNEIKPLvLipSqNEPvmgp9
Ptul42kTX3sF4YBXP4rXVFSbpxlfxU6nr2I47v+kScaj8xZMlQcUIDw62iQ8+VzT
BTuiFoZs//C3vccK2SaYoatvv63UR9faOcgqkkgr8EopuNSUwD0n3iY/tBT0IdeE
z6jseRY4NFEmCGLhA0eogcw9lR31o9XxB+AcGpxK75Enkn1zADFhMXLnowArNXC9
WuqLIJ6L7OfWh8st9gHUsDU1xCMkpL1ibuUuAxn4U0a7ZLjXEo1Dtv2PYtWfd2Vh
G1UjXbYPMfoBqkohuFzDyknjoVELONfUz823u8Hz06D21lheT9AxxBr/T8pzPssq
Uml0vHOgaO62dY5stb/pIHfS1dn2vpkplf5R0FpU/Be8t0P9HTkLECgyUr6/9mtw
ZNngwj7Spa4/86zXXTRVAmg8MdsE0+q7wtPzfneNzvPf6mLAHO3jKxCP/Vp1XYSO
8/WDDs+wpymFg6XGyYASkuLfPFKHoQA0llNhMrFvso8+fsYAkSWjxUmjXKer5TEW
krf+jSdYYyrV5AXpp3QyqMbjIr4UWvOdcdCVkB1T4RYT/zD1d+q98kC4F7KtwTvb
DYcqh5jvhtHIvhbE1PSi9HbrVeAfxFi94KCm3k69k5qoqLCUXr7GnB8OokyK4Fpy
AOFfdy7EiXmj6gSXo5qLD/hNRXN9XmCilV8X2ZXUgNSoM3FlaQxya2JWzIVECb5s
OIHW2QxzyMVDgLu2uNwZmvXOJTeqZVST1636nIw/rqauxEkgPruuelQ9xkqV5GKP
DZQT08Xye8QDNs/HBjbhYhTIJZOy7ISGtIWQhpkPWi79i3kc6J69VtjJgzYE5DTe
y7L4+pvRa2Osc1b8xborVmKanOz2uepGcEgdeyVdU+Xnil+pEM8wUQpxmnX46F0A
7ASKb+SlX2vno/jTE4/am/ED5PFdH0bWZx22clLovegWIMMiCfJrjFEs+Ia4c1SQ
831thjNLI41veWT0g4rzzs3dcoV3/Z478qh/f/9YLrkh9uO/UGWMknJ3Lx4Ye+Q1
ROSfY3GUVK7zetiQOXY9vQFfTqqN3Ipv1v/OScOm3L6vG9CR2iWyxSlkR3fTGZkZ
wydqbscqLpOpPhiyNCr/B1f+A/ZMwdN0o7PDGTPPIqYm77GP0630YiFgwcnPJLr7
MYkr9WFHl1jE9dSwIs9JlrkFtLENp29WGytRWp7mvH2YanNOMGecqEJeYS+2ifnh
fvzwOxjEErUiOMufXLysMtNZTR4qwBEGYR6dBh1tI4K5HdskIF8mRxlIH2gxdBpq
Di8N+AF2P+LLqiZtPiE+3gLd57UfOJvsbYMoTpFHrxFjPFnC+SXqbS4ZV8oxNMuX
v6LC+gPB/L5ueSNwUo2og1KYbIapXLQ0opVwFws5747QSGSoLlvgl0fwfgnBhEqD
1wMYN595WZRFrBOgCh76OPGg4SRHjzXOufyWEHfSUwRvBbpUd1bcWcRYm8UpfDNS
fvTdXiRc+TAddtAJftaQm07GkUcsMj3Uh4bc1+QaUV4OuhShZZzm9f0dp3VBhIVw
UwLH2iiMyunnCqH43Srn1uCfwvH3rc3C86EmDklJ2E4urNpAiIEcejvmnqo3dMXU
LX5/Z2wkh45gCTzBLbIf+R19HDlhWdM+7kB2DAlouH4XFHCclfgKUi2Kd7kSDORn
i2JLN6Fyad7gahcJJ5iQQTISqctXQcFn0w/mk3K38/PV326ZXG9ssOKclfnFUdGg
pVbdnvk9OkK2sPhXW5zzq+h6khtRgyH3G8xzd6qeYD5JqCOAxZnsuB+7JDNC0no3
K0THjX1sCSKg22h7qGRswigmEAYDPFoUtF8UXuUKX4nAroZaIlR9XvKCJRs8M8+I
jCUq2gHZ1ipDoG1HiGys++9ub74ddtMb26TabpMhTuuOHTzci0/TyFjDmL3EBa0h
KN/gIEgAvjlVNARPetvUCAn5pvXaRtOiTulGNcWT0nlvcGxgBalcyfa2nLTX+rXi
r8j1hUBmQtJwym3I8sRZ8JUH+Vb3i6OiqeTyIbmEd3Mk6PE9Jl8cVhqwxGe7dRrr
6/Me8+qErvta01ye7D+76rAzeJjw1vsHZKSwNrngnQBmvUzKrDoQkv5DzQ4EAKjw
zaT1BY/xdjUznFtUjDzVDSe/w9sJigWOkjAbLCOqxpswGGDEOU0fke1eLv06j7C/
HfP516uMGtL4aar2F2fzbpn4VZcnG3wnI+SCgjd/u2QlLpzk05pW1ds2naHyRQ8O
G28Hp4l/cq87CajEd/QP6IhCuaMJ2U9qWDLQ90NuYB5lmACxYWPxoWVNoQD+QpWT
5+MaNV+WVCEu+qIm4B80mt50nZqp8TUGWDndP69ZCcvskYj/ZQZ41nbgkwrrcnXs
I931ayIUUmd5AtBoopXdL6Bw+gpmjBOMRUY1YEgILKQLplRbDf1Dg5/LHecGPdtY
dbZSzJUFKrLG5jQtBvlL7hvd4hfFc4sJFyLuctze6SEBNXoWUEBjkevRzxHyy12U
3Gw9ke4+GBkDQA9V3z2RCxu7sHIHydhk1MXNlI7uSfq+w6KVsFBQYyQhVk0YVbCW
dDUrgePgP5rZGNsIf4CLTY9NbqUg7mXPGo49q2EXtc5hr7Kt8t31H5T6j6coin1H
kxcf+qMTWUp57xSWf+66xMnIdJOq1xoKfiLue+zKTl4yfCtQYoLc3weoz7F2WWNQ
MB3zHvRe5khpH7slO49nArOXkHXvjo4WP6q1CafKm8z0P4UWR1OTypt1m6TbuWPX
wOwsEoZYwfnTyEJjefIPijZkMSp9RDf9lEncFYHSfXNwIEjAI+nWRf12hRzV8tNv
1rubk/GJq90ag81KAFQCAe112ROOFQMEHfftOlSNb4NIB3SlKQKtJGrlckohi2wp
B6wv8ytWBRevaeATqK73w8VnW7Od3gLca+xsDjt/6gJPVnDoDC017Q5tc1VtONSI
u59YnldicKYdpX93OtzDiMMUcWnbXRb2mmH13I69JI0K3Ro4GrXsoVpHyGM4UMqr
q693Y/IlFakt0KXVnrYxdSaPtsngiqk0Py5frLRIznZbR7bDbYJwDh0fPjSXfTiz
J4bOWDTP6A/eIfIRE2waLhFGO/ebAmuLjRqnTRkLSkiz8YDS8NX0toKyz+YRNnUm
L9KRvw6/2RcaGcX6dMpwnC+3wzbAB2CM0XXPFgQ2yjJ70pZK5r/U+efOcvHKbseg
tIFFjout2ZdiFBl/FQWXNOBSDWs3QfVbWz3ZNZdpG2QWY8DqRK+b8dlyDF7uOyNc
fBqlKXAMm3vYJ45j8By1TD3jtaRcQyjLZN9OOhBxbIKHGT8AAXpOvf+gICUt7rPK
DGNzUOe77K1QVkYKR68G0nCJfwdvAC1PfCu+nZbMmHXAlgZnxA7gu8mGfJ6OUUic
IgXaFnp/+25FJEzhB+0ATzBBRovbsOiH25xpPc1S1scOVIRVu4TZ1ngkHaShxdbs
yqkF8K712RUPPOi8WsWXpQwnIMoqJJX5LM5/CcCzyct1ZPKbtXgWLPDUaFIAcNYz
Vpy5I2G+go3y5bLxwp+2dqmoq997QLUC7eB5V5Ez1vfLyi4b+JAflXvD1xmIyqlq
ys6oWTohl3vnVgG4pnW/BQaJ8eAT+usnAPCVJNFnqvnADhS3CBnbEHQFV7ZvqUxG
Q8X5wOssgWgNBERkn+ypXEdTBOJeVbWWKaw9RSYPmU+CxuYkmtIeINi25R0PpSVb
8FkVgIMX/EYp4UxkjnNMln8236VDYx0qox/PvLqnJtY/LAJq5R4LwEHt4Z1u7BQ0
72/ClAl0LMCXceI0V9k2mm0gejtTRIcXH94gxIKU2kPsQObQE4SFgnN48HfdAnKx
S47wwdxG+GQMOGpfqu20V7LocixpLgCtFOG/aYlRecO5i4kaDx4+ROKsmtMkLq0m
J97lHdyNteYG/laNCCLbb2s+4ewJj/WAFt76wLWPh1x6zOHZpEiyySdw0gOvivgU
44PVv7beHXu3J2TmPpLy3aT3ZJNGK7f6YgXuGCR2CQ5g88SzmlSemt7OEO55ajbS
lcx673Tv0j6WOZQGpJzR5pdD1MzbE2DDZvIoUPbtVO7it8S+nMK0HiiSK7zOXEcB
QaRsDSklZaZ+zwVPccyyi169szusAVBp8jzLufS7vnKsdjfNwo0eCiaFWlT+/LeB
ESK9P7lx8Te6cY+Z/+4lvfAoTaWlY/WGdz3+KpkdYVFUq7vXPAOdZNLj6ewt7GBg
z7Wh1PjcVIn3xYyXIGwfiRJwVMqBmW4GJFyzqj9X6wZlurVj73A82fdIluP7oEBv
VTeXR7gIDeJobi4rr85g9EnC1SjxDokuF97+rMiK/dLFDa0W9ib9KLbMekI0LkEA
ccSVbeEigVaZU730JwEvblfeJ7j0S9tWmHzFUOYi/i30HhtH9XC62ldcI8d24LXQ
aNGrIa73zcEOhMDcJwLMOok+qXhOLhgY98cr2VblyVOsKFd8mZOCeroVqJIN8V6n
x5yCe/sCfImW2oNISmt/lhUSx6mdgDxU2zRQ6kRNvP0PuIBqkryNCFo05hkjmycP
W4q7g5Z45aP1BZr3vbWYIlkuC9dZmFOfCdECFe8Lncau1GwbJlqlzTTYOeTtkJTQ
54KiXuf+4vsoMHOWupDxSSaod+8LfR0p+hM8owRMw7JWClyo088DOWCu5U9RsLRW
SbHu044O990CQ/uUcQZtUg3mORQ+i553AmXOSVbIvs1Cl16Va2gbtXduloV/ALLo
YgLxWd8933zZ5gQ53V2IVzKLyUwxDRGXGONthTST25/eKRH0+UVLWyP4OsOvJJlM
zDizpAD2MZeJ8DEAxgy3Tlrrtr+a0RyMxHqAKod4mUuzQStZt21ORAS3WQ09S9WW
e0NkoHhdmJoVHcu7h36+NHFEKcm5yeyZC9YZOj641e7IoEC7tPOgiXKhfrjMpxp4
w6eo1T72bO/J9uLMK9PhviVHk/S8OnvRcna8KhUwK7sOnvaAD+7jsjkfbNP/J9cj
XLOJopdgZfaR+6VMtQg6bY3vVbNOUZCi3LLO573ZqGOPolXp/sc6lkGVU64gOJYo
wxDiuygshezhMS1nwPaBrHY6ueuvj5RjH9EFN8fFMDWMoI3P419j5J80czCR5S6R
DRJnqWTX6YiTEHKuSjqY/JFBR6ybCOUIYLRU6OGMXJxPANC9f0XGasGMl+F6WuCY
nQ3jDSY/xA09jXn6zDrRNDuA8NfGa5euZu4KzcRJXi7MKHXsS6wWkdAn+PD9JE9J
3Ja5bUOcl1rAW5553VmzIq19+nTH0RFxBH2UEPX8zYG5cXxfJYnAfZp0zY4ZM2Bx
25Fhc4ylqQ/lWpE94mSUuUVG4ZZEZX1DzCXkh6mAKJ3nLsE91HkoLviKKTVZ2Lwq
4ZTMHCOn2NKsmFyhqFRbo8i4sBsXe1W27A5pALtdJPn9TsNXEH2aEVQHcELPSjCD
aN9mB088XKoOqJT2LQpNuwKLaTjHuAVTqRH3HtqlU/Umw2mXG09es6opVF3uWU6G
C43pgHn+K70CGqIMxCuk3KtDWDEcbERLCvrxn6NBFK7tgE0szyw9mGpMhiGBxPEK
wnhEMQkwIr/BxSg3zX1GKKvmiRne9wH1xkxklX8vlhwQbDznFiDoN7T3LGwIoKCR
IPjjDtH0cnaXIyj8qG43Gor9NPAD3xiie2g2P7neHCvN8yizrKfk2naQGDJ+7Vk+
/Cpoz28rUnMkQwbFiD3x70EWgiNME7sByNhXY8Wk8zZ/0bxAHnrqrEd0xaEy4MQa
ZQ4G0g4tay119TSdr5Y/dQTPWlK9RvpV3iHpmE50MzV2JM9bPTVkrtKVmF/q9PgM
UETuTz5v37wvVZ5+dzapninlfkbv0A+7Hvli+S7j9YPlgSoif/Yx6B95zXEyGdSw
Qo0WXmHNxFQLRv2uBxMM1IpZJpwWjyV+40QAjTof38cksSe7Ioq4yVstS4Nh8lQd
6HVAuXLIjaZzjGMpdK+TNGUxYV5wr0FLaaaWNGKfCogHFLOeteyORYzEhBPACf6f
rRr2du4tUuJmmC3ZI14oT0LYZ/8c5u9uETS75PCQ5S+7WuizRMrtUvADVQT94nKP
328U72IhjEIpRXufpkRcMwJCIlRR4ymm6gJ7yVbq0fPdhLmIMXJYVGGyGfTCi0wf
tW86r2JdVhqTa2hr+NDAC7UJin++D9ZP7Ozn/xs77l58vVw89RL/mzAnlO/CYH/M
UTVcT9ldtZn+mz8067835rVsFkeaNTSRWoHwjrnCMYhAr9LxpbC2eMsB9uEoSVzc
CuPLMWHVVE2lJ2VPO98J+M8Rv0Jp5CDMghSwJ+djtnnDKp+CDM3pto6zEleSABUb
PLoE6a4GLl5qkHR2Utly6TbfBHXFjEKoX8izqZep33NUoNxH0UcPpsec1o050f1J
Cy4TQ2BK/r52vTprT8fE6b6VHXWny5y+ESdoKIJLzRsufe5G3mBY0j0l5VlgCMcF
ngKmmf0WtR3KcYt1KNn+WETx02tlbIbRW69obAUZYghWebUMj/oa/U4FNGuxEgaO
rZE0zGLDQnCkTODivDLuEj7IFIUMfzoRp60SZpdLK/2S1FCP9iVzvpyqf7XBte4y
+J87UeOPj6q4RlqAMFRTQXQXEMDyLHYxDdoKtQqPKgMW6Nrrl0ttSmaIWnmAdJnU
HMUZ35QQRax93CBhOdfS6CzrTYsHWMY4YwGRguATH3TKzZoAH9cc+JGDZIJLlUf+
yPf/8SAifDPHl3RXX+MeI/uwKykv2QSAkbR9VBKmlUr+cr5ZWvp728h3o7mvry67
pPNLM0HThLpd4fLsEUhACXKiyIyQBwCE3DEpv9p3hZPolWDjUzsgSejhVd4r+WXa
DC2ggGQjtmquA80opThd647JFu6JYLfcBnB0OzjX7eDYXc6C76gGePT7S3cpippw
f0oS3A0Zirxc5Zc5XJwelj0rRKq6EsN55ABTWd5E3h9C3U2ZYqljTMYS0Njr0CNG
89FoWgn0eTxVljyzCXVsox/32gyNYMJkKbjpfd4axrqfaNwnM2ys3gzkKGxqFNEL
3995m9kSyMCV3VvSFE4X3kgxCyDTu15E2ROR3iYjY0A9OX84Bl5B6WAsWzoOXh9x
g0VVH4qgQy3gu8mX3Ksrgin3ONS3/n7Hdfh9ypIynITJ2NWw95V47V53LjsR7Bjt
JvSbf64iOzu7RcSpnkBzpTHa/xtzg53/p2FHkaogwb0aVNE3goJIMYO+4Wc6mw9Z
+wzM174JbiOl3nZCSwoawtnEUW2AzYlIs6aYzZjeZiqn2L7HWNE08y4mLn1yH+6w
YXM0odaB1JpyXun8+TP9dyqcLiDkg/Omk+oHj15uKjXOJayGk/zkudKx8yeBHLmL
im2o834RxDmug1AKeEqQ31sRkeHvBWWvBvVuz38DLtBoUr1M9HykqyJAJo4pAZSg
YPObRi4e4/vHSAKO2Bps0xo9clDJsjDvA1vSk1Unor2ws1iEy7/URaSM5x622wV8
n7Md7dxFK4NZpsreqcb8827Ushn6kLnQJGzHvub8GtZJqBBFiT6yfPHDpzHKg70H
NMNGnBoPe1jRT3CNYWbKqRBQiMB+Ak8g7oY2Ai1a0zuKTHyAjw4imCk6YMoXyeZN
TL/uk2KOAOyIYzZq0XeDnBSJ5vWhXyzv1z9DCfQ6Fes83HoVlCb9CWn6yoEe08Qk
IxEEMElj5YaeUySuTW5lRkOYZGyPcZX+6BzGg+g8aCYmsd4HaUXeIpAnGF2DJNkv
76eQmvjf39Pwt1Kj4jd60MOh5iq9cLAwh5VHUvLGPi2O++bmIF7egNre+3C19iUT
OtcGcA+HZJWtiHzRlapcokyGUk/u81yg8aVGiDB5A417/QPTywkYhb7OIkSA2xin
zR8OhgHOJYxFPufHDPWJXkvYTriMpyb4q6Gua/9vKFwhhVAmReWZ8yGmZWhOi6vs
dn/8OZqXIMizXUPZfxRo4Uj+aUo3EXQwZa2WhMzcJ+HeS40vveDzxQzsJSjyufbU
xzNpCcvt6oAEyeQ3jfVUPpohgWKY9eQpH8SM1uWcH30e0WgOAaWfUCePkkuIXHJr
q8/y5Zgs3iFH65hb91AyyF851FdtwoHPifBLIa7oqlTSTqEnzXDmwCQ0aSH47Fzh
UB8ZvOYUuEaDTYDD8VUg722Kjtq/j+2xaX1iSzlFWIMIbHfXQg2rdzeKGsN1FLSZ
IKs7TlUbQ5OztSmjebJ/er0IBDPt4K3D2Ibf+hh0udckO8w36wcJHUTUedo1K+3y
FSMUshluelN2bZ+MFgbpmOYajP5vLuMLHnB/LyH2jwGBvdCONbdBozzINgRx6ZyP
ZChztnQfO/2f7qrVd7A9is0v4U/wCIb1C5OEqjav5WCojAWXU2M5v0daw3Wzqt+R
bBoLXwehL+Xdeu9E639BK+oX2aJQYtZOX7EmR6Sq/ZM3H5f5tMDv0cG+iDc31R4z
pm0VEBSbst2jpFKMkx7yIHPrmWAlKIHiN8h9zNVucR6kbKogxHqcZaomRUYu6JdO
PDd5qHQUPJQGlRBBk0XYy8UZ2ZO6XnEBUlq9Zjd0eNfMh1G13qHGcAX+3+2XXGVl
RLKm/0l2WUFnMPKGAE3AUjnduxUZ0Od5spFQRCg5bqw7JJTkJF061TKXHLSmYzxn
7qkk47wWfg6rXJf6JpRmqJ8SF3KzM0vvMnnNzSnD+YTfDZLrhfaVueeDT86do3Rh
7YDa+wLPZ8EFIkSYRUQbJvppzs5d3t/L095FG90xHigHytxH70eKlwM2/wNYjMI+
4pvFET74tgxv68/y7SJA7p9FWrsc/uqf5DgYXv4Jvc28B1uAIXeg0sAzBGJk0Goj
6qr4r6vn6+MSp73DQd+nQP9nW/8tBOoedsD5r5JfqCSfN8t5y83jDzdOpzkbx2HJ
20ondbOsqUaFPImZjbS0ilHcE42q5dvNNqFm/6LkxdkclpVgRcqt4engqZECCTdu
dFF/+tgfHgX9N4D4rnQn3W/iTnRwuyIOiqPQSj9yYuS6LjT6XLHAGSAvysYDXkCL
DmFmRGPsYkgpYPpqQKDTVqx0ciqGJdDzH+8wgzVsWT/QIhfezS11S0FkDJD7rD2p
IFcYfuKEDAoVdun/+m2i1CRUbeBC1byakb6yI4+sXopmoj2jKLOqIMk/14RmblQm
UUMllVmTWjrRrB6/KX2c1yl5p2PYvmo+nUjAWLqucrql2X9hJWOJYCupXwoe+Uvy
PddgSZKcZtuL0q9poyzEcRpwaEBskjyIM0PXfO0gsNndo1JW7/6DfDaEw3eJcaYL
XfUqCZ//b5jLlaVC3ZVTvymoJw/mwAqC2AxGNh8VwhkMVO0HuliqDlZHyEGsk8q7
IQkTYdv0WKg8Tbst9uNiqLETmUz14JMous8q+piAcwCI8pkZ7XQEQmNmfdPP7Af4
VTd8QsLBX6kzxRsApMphv9TlUaC6ej8VTflJjT3e/JthvzCZMY79lhYcyO9kx8hO
28SENaBMZMcBOqW3vT69vbfvdGNyMODdJ3oANP8nQ9+xGmSRKV9GrWZi418eW10U
zwJkPbZlqTHzzEgaXUJNlMrWxDDo8fKYcHawWIQCEd6+5HNZDVufbZxueTXsT8Qn
GzUuh4eKF08Oeqeocvb6Ah/bOCrsR/AYK8IH+dtIHGCoV9FaWdkNFXBzNR7//tx4
zshLJy7mOSsPepz1sCDiN/0fJabquReVEoF3FSToGaa0ISH/fR6x1hrwHlUPHfX4
djxnmbrMOmbkhrkfrLGw18eBaUi2M/HFICcu6jcwHRabWSE14WybDW5Do90gjvHS
3u34Tl12dC2sPDokfVyPeHXLWusaubDJluAzxFkGM1vhfz8xepjO7tTjG6cWIW9k
SH4v916K2WfbudJpymMBj74jci2yYC/B9xCWi+rfguIpnh5qEDQgOWF3pIite6fO
FQuNbBzo/fysswCgFIBXIgk/KtEW7TRpWxrp+qQGdsqNc8IXIde3Du9laCjS5F8X
yFrzCCYvzJqu9uWlHJOBTtgdbCJmVwYnnIQNAYeFn1dUaUCDuY0fcNinNpmtGw4u
+b27RP8+tDS9QTr8fBxM/f+z39nzkBTMARi7YnjY1DG8hasNfskrAiYMIiUnAmjV
r5T/CEgxzRffkZX+X5f79l/Be0GcWv7HkH1WjrVO8+UuC7RMV+AUSLyavUnWFUKk
A5ZdLIX8Fw6J+GHL4qfgBxHQvWL0Z0huoCj6GCCldYcvwAs3fL1yocPTSTlKS8n2
N6whNhxe8SgYRO77Z3MNQZtY/rxoHSbEUSfivARtwFE9sg+aUHoixaTqtd+Ah01w
4hm4yycz1kBiiWJOUFtTGPcgy4NVUFS365WNQjARHLxU+XrLCeToHGrryJ8fmkQL
+W+NmKWpzKeaOjNOWAhvDsxO4U7PwQAbddi9+3FLpvvL9csVLp5JUTEjPiAbO/I9
y3ufYujuhXG3mOSvJLkdRsqQNPIsuHBnWv/LZJQoEs+if02TVeTkSiUIEjZTftN3
Z7z5LYk/1C/VdeoUXVP9GiQr+fUz3l5CIRvtXELlfZNsDQ4AaJzYC3Teh+W1H28a
fA9jbPvUQ3n+eKqgLtXvJoeKBs7qAi6bTpZoR13VTTNbGKkv5ZXCvTTGEg8M2f/n
CJWIOtZZUWQh/eEIJldt6R8zuf3lb615YZqhK1T51HTJGLlhGF3lVY+xeaZauh7Z
dF6EdMX5Hp6/7lAGvFYUsKKxKGRNUJIwojNt7Kn4xbxzHozXYWM2e41ngABr70xI
eASXEhJj9cNVDTUpO6YG3MA4T65bTAMBqNO7eUqGBINT9BAvS6IbMXJ5tw4PzvbN
M+JE/oVGomqouZoCSjTgWpTyTdPjn+bKxebi4bzexkQOT9TxGtiCpJJsrXAjIjhv
CPQL2DZIXLn9gtBjvPV5IQo+klxvHD+GVtFlOiCos6EHqN+2OQCes5k8gV9VS5QH
VXMPMjXoKdKlLVH3R31blHqaV7IDEd/N0g3DkNJtkFxy5v2cWvd1I/B4h2Zx5QFm
BPKuXkVg7/kJGK1d4eeEIhz5LarU8vXrBmiDfeR8C4Y/9diddMi9RxaLpyIG1Av9
Kq552Bj50F923+lDcjTEVDNS7HpEssOL4yFjWdNaQB1HMBOvadtZT/pVgMTUhE9H
lVZCwAEqZLBzAnkwYk60o1THkKZd07G7kNbP5+bpkYFVt/dlR1qTXpua2DEtMREk
z+i14gn+tnhtGXd6u5sIyemuoODglazXzcPhUcPbXYsEJEX7rno2X6Q3cP9aS9MA
5PF7CK1JM+GeLG5kkrNoK8p6RvzyXwGnKhhLZ+TvDMa+94Ro+eeul8bEJ668zLo3
tSJxS+ThSJyuoTpEUWLQIL6j+6g6P5Y6yYBY9F2QZDyf42PC+ami5vwL3FgqwIO3
6zzKzChRvjAvi3LeIy5IB5akn4/cUKcNtMEQLTkY7CY2kPqX75f8T28ariMQES0O
q5Op7tXt3lNDQ4/lehLgoQOfGijKH/+wwn4ER8GIPjarYynhvlJxu2oSxzdlm+oX
wXMkaWD+ou3LX5lWW4ZgFi0v204QACAiJx9pQ7h2XXcgis1He28VylefEVlKDJUw
b5o4y10YEyk8SrM8tQNkjRHL89e4F2QzZ9dPDeBnJtDyJYnWYHVNQc47hraOexYY
kkP78YtVmqouqH3FMtV5N2ViwMxMtwl6/PSZsSLEhTAmPnSLHw2xrpRLpUJVRahi
yW5rbjtHEzhexjfJYuvvH4q0hfp1dZXno8UU+VNNYbuAsDPe3tiHtCC6tSIlXlZV
v4bYQhns+CyqZrlMiZKNXPYotz+HwsCmbHR0HDS4C3MOQnQFJ4Ipo4q5P5W1FTGv
j8JpK2FOfQz6mq7VC/lC2BDURTh832/UfoDj99CdXXGxLbJ0oyVG/4CGz9U1w8+4
hBK72RA8YfGEYVKNBV62tIlz3jSquQsC0hEn82WTyUZOiodrDRNahxFlzFsYRqUM
35u8OEduvI7SKR2m0qjmcwL19Ub7hTEiMFDrLfqkMGuF3AIAQ0p26S8paKU9k9Pf
aRJUrA9ju4KjWITys6spfXVHhGidiIRTHyvDvWycUq8AS/QRZItU+urdFg29vAfj
6OzhngOwxdSCXyNtyY5C/ifi0UPiZrUe9PGjna5NWw87SwnAUbNR3Nt99Anlv67t
dPG80j+5wRbZCCCV1WMj/H9y6lQQB1UA1lpjUAgQf9QdmSyiMa8/dBz40RiMLwEy
OeKNyM5l7dQrak8GZY8imuWFIwiyvJTD9X9GYfSb9OudfYhnp++3oXYpjapfoZZq
SVku1xzrhdrSfj//ojFsBQ+iJj9YGac4XAy95gX905CXft3L/BZFQFlmsi/bAM+4
kYjBmiKL8Uv7i4vt9H+5rh4yY6qNrbbrD7Jkm4kSurCjRXPNUFZceOnFdSM72CBf
uTkK2QUlNuWc/uVbZ2/vN+5GJaSTmQUoh7OPaSf9ocfBuooew5XzH6fWC1aKBdhh
73AToi+UNTUN/ftwd+CY7ANENqbHSpuDlFsrgUjhi2+Qbwzvj1wPk0WuM7S7qysC
38JgcjUCq7oaQPVW4rQsn1N/I4VaZ+6cbDywsYCOzznj17urOJ4x1EJLUirSIOTd
EHdOFZw2/cgO2JlHuLHFrQ/kb8eJrx79VDMK9zWcyby9lGbA/zMdM6JJFGWVEMqi
seSmSVYnhOSmpVO+rF6JD4nRDGRltob1BsqBdzvED4H3bOjLDWvutNkyDXAx/l+S
PqXIp8F+52PmNqyF97JasqsGvuwXCinqqA13BoLEikpvXcSsr8CzYAGBYN8+J+3w
kLowuy6vCpnY8zVVb/uZyxUG0m1g63Ys2otuEPi3alFoNg6dbT+c/DrWfFkju5q+
qmX2a3dLd10kLf5zkMDMEz2br8W0adLncivbWvbmL5qbI4SWhJ5iQ1Tf0N5W45TX
Hp4nlvOVq3DfKhXeoK99S7aanoiglAWbmm1qvw1mvqyTf+RbVer8Qwk7duhInKqi
ZYN+AsQy9RzHXK+Pr507O8XMqDwNytnXWkah3juBDzyVPi2UxkOzriHUtqNSQppJ
MsJhndhwpLpQLDubZ/iAE1HxhHTKNL62T7qWCKjk7UHhUyVNWTTdLzKQqqA+vwZS
WtyBag4K6dTkmMn15ZK0KORshJVlFYtn9o07KMQt3jhrtFz+Xe3PjzNsCVnFC2dz
4i9+f6Zy/UZAIejD6dEHL8aqRb6D6HOQiYj/Im5pdhKQ+I4WdUsFwwz2nZHzcazu
hj6ZTx9lHyA0UWtKqpKoesLRyCGwX7rCmrjRGAmdy3jCHA2r1WmYW12K/QqnEP6w
6eVNKsoDJzQ7wp2BpbmyYbJlFULJUv8BFiXEaw57HKvYQmMArXVvomIyCNjGyKiw
BX06+l1dp9PsF5jFaGsBVFfKarJW6zvPZhzaJkGfDzSgXE4H4hWt89nXo4emXhgs
+xs9IMFbGouagch6np3EIdxj4GGOvpApHJhsZHVPXYMC7mf8bBuhNqy4RNeRMpls
3Xh5PZ825rHl991hV3jOWUtSUn/lE1oE6yCrmacI/tKweWzTw5fYHKceyDZaAjZB
kGGfHJfyWny8zoEuPVl+V1HnM9e/URfRl0DhrY7EPrZnjzDnDpZeaX72b2+CHyMt
/C4fQ1qC01u7xXRyN4ZEZNTjmq0fWFpBBWN45HhDlbPbH/unT0yo6AB6RxPPbWHv
7m1Q0fZT6tvYqbtOFSyAU1U360bZ9K3fN48BMX/TEi7PuHGuI9P/ybpvzO0rFCIB
sv+RnjVqM9riDi+ZrJrsGxFkZfAOcxEZXuLJ/qkWQY9Zb8AHMJLYkm9hOPPInl1I
M5re/KkVhZWgkOWIOiEoIkNmgO+KFLiJut5/4xIHUEQX993YefAd7rPPEy58ryJ0
4UumPn6kqb0M+4KldbdSl359ftltFpUNN1KSDf/6OJl3wsm9sAXaRk5PIPWxWUt3
H9U1c8QMMvpIViGO3j9L7kMaoZI+JsjKDLiUAnIkR6WVZ0o+NFv9KsoM5n/ehZsb
75zXPdPLO2q9973yQFpeYwbeaNMsPHhEfkNk9nkJto8lE1CU6XqIbK7MuwZfFvPM
ZkkYjKE6JHFGhTF4+gvuB28k+D6ZsXbXq1lzfzlgQe7FqKsMdh9PZFAHNpPvBlN8
PQi3mQYQVIhZ+R8v95fv6Z7o5fx/vsbL09gdImPGGbd5WHwTRNiAM35W6V33BrO+
ARGueHRy+62iaAeVQzwWnzTZoLQZ0GmzwjdQBm4meQ8Iy20BD/gth2GJ9WowlVKI
ZmojNfcd7DTFpKHA4ENqbDRTxOFgoHxo/YmZl91bjzKrlUPNG6J/F7x30I0LxHKB
CRLXqWLwwzTTob66DYONsOeEBsjCXGNkn5/X10MW3mMIubNP4MeKK/nlLDQTmMp2
aqh3aXtyWCuSaA+FVT26GAc25zZyWK6i5XZKYuUm4JsCU54wZaUM43Oy52CyAZt1
oGKyIrIbWIxTofOJf37549J9BXMoxsqbCfk6Oz0oxPshXkcTuPgWaW2P1+745LYR
/IByofWcpFohoh/5Vkyb3H9E5WB6i2AbzFlYvm8pUsMkk52giNjWv4kAINnbOyvu
5Iyv9sbat/wyX6bzVndJVP44WaYyMLIViTvRd2s5Yq2/mrtKurcXx5GBrz27DU0j
lW8bUnSTf+50pNJOYKpAYylwtOf1Xizv6mP5T0dJOku7GqXQSIfoFx4bs4YL8lTC
FlxApCZLjpJ5NI/HvWhofFPMcu6yao8UBJPIHDAFDXmIXB1sZKDXuAvzfda3MFVo
8cuCpbQFoMGt4jYbFlA6OLPp7MsJ/It3w9AA45uMRb+Vj9AXVbX86HwJzYX6/hVp
UPeKYyhqnIQp+JWLanEgp1nFbAbJ13n9A9tuWWBNzT8MDg7e5+nyg+cXIT8vIi7y
5leszN1YgrK6GjeA9qoPlr1qJAsErkSTBJ0AGSfFy65qVa61cXVSwAxi6OxXFstM
StNtZ62lPryq+1L0hVhqkfF5P3+ctTK9jYbTdlzaE1rLLjncueBSWWUMALtkUl3u
WDnBlvxs9v5ksrnhAtYi5n8iNgoMsxKMcDBNZpa40zC+/NrQM2qeVC3i2WGmJHeq
eYwset8maWKrDWTaCii/uixGWNyvXIZwpRjZqBldXF6mxrPkwDWW0KW6NXyOze4s
1nyiHdFJc4vfRIHHR22q1fYaE0YKRv3PVgY9xP3YnXBbwO5DK9GruLLNEa5ZBuQI
x6DPB7dYNUaI22yhoOpxN3inD16k7RXN8MBBA+uZmzoUgK8oxaAidw7ZF54bxM80
m9qYXxHyArQElhVDa332VmQ8UROuBCjEyKCS8NeBWj6CW/kr/wyhCDTsdzTosQfV
x39i7rt6W3F7qVTT0x+nCRHr4bqFolx+jFbiMLqRql4VBbsRnMRoNZubuWBKn7tN
f+26S7HPVtpie625xI/w6dDxhCChvK7DlBWp5mgoX15TzDWCUlR8pNKTIidRhkOK
U+61KpKYr7HBqVvJX9Lrew5EVKAmH69MI/XkfG9lfvuy4kmCYofAPPZwo1zJbGbh
yf8h50VwKgMG36IUaiG/uEkfdLXSQo/mRJrlIVdAkyYc70kIX4xSxXEUinJN3Qo2
pkonqq+YUeYpXT9k05EQIOkDOSC+rwm9FkCKDZujh49LXGMomdqwKYWSxet/s+KW
fd19DKO0gGtqfPTSkh7TdDo+6lFWTlrzLhlc1Ds4h7L+PiLO/cPRKTnYtv42bLHx
xjGNLTA6mULFMhhgJIMM4mi3pfFo7yAr7+D0lQbTjk4FK27jOO6kjtNAqnHNS23E
O8XpV/SY9bLnhjfUc4Q1KMhvOs2soevLjakroiEQSngauIEKr1BjO+R2CRmYh68M
XmmncQxbAd2rA+fFOq5OHU6BpwaIy7H8whAUU6aiLzbUb5qR7j/+PaOEoh5aSbtX
DvCg9wb3dKnbAumbhc9ZKknrItDAkIIDhLLwGtvYPlzl2hW6wGHEHmFAi4RIlrkW
RTnA8+N4k4xRw4nyYIYYwyh3/ewvHjrDu40AckqYSSu+o5q5ulKMCfVjHF8wEcdE
BF92XMGsSZSlSxBOCucqcNqKg6jDBCFq3grQDwBr0fdBNXZc21JE9ZiVI2vD4NyN
bsBWiphVcTR6FIOIgmYO1omPhXIUAqjPKVPP1j6Nozy5obT2ABE31yRJsXF5DelC
ZSg9xDSIAGLnIx+k/1IrmKRLoRPx+71aJmdwAPsZ+PsWT0OJ3VdcqZWmvE34K+9U
IPhppSNXRTVSGt/Earkk8/JWoIYwyqHRjlWy2SzyLzDtaiGEy796jhueDU7pshBL
wUgZ4KDNNLGJG/ad0I1NHIfQ/CvvgVaQLdRk48Wj2PS5zxSwTaowxwwhaTuxiI54
HmoS7VLiCIW++8GD3BAikV+Mx3PW0ZQpxGKeYKOrZnrhQdbazUpE2zpjnmwGur52
mcOJtjNy0OUvxpyr+Zv7gdpn/XBDUus/G6OuXuumXnTKGx9thgja3+qFzReM92ma
Fc0Shax/oRdVpr+ZFd5pOnqETC9v+JFGGiCjbQ/c72Y36v3PoklbsAKjBhqNfx79
kE+MAkorHPisX/sEhrvxObUpFHJCAJbdqqXC7rIC2VLhQBRZ4BjYXOwSozK234hy
pI4d8SP/yqjd4heAv6yGpRApKSeFXDnQJFWhbsmGO1p+E+9K1keeaBXCrymFoLJN
UDmWtNReRgqPMDXNbgTzfObBaLQmOhZJMIymtdptw57hxXb64TcHW2MAw8HWylmV
H2QaHBXBHRy7wz9ma1+5J+SbHbQHf454wYYR27jz0HzsXgtjENxXb3j/ZKl7Qw9T
8H6X+gLcjy8j3Wri6W7IxWuY8UiToBnpdjRuanr1lmG153WSbz2dwzAmjDEwlKSW
8qQcZcazP11YfQ7Kc90XHNBNxa5RKLJEJvP4ULVhcQckkYyN/A6llDNFr592t698
0G7D0Vdfo+eB9NOn4S+4IeJ5L1pRw5TQCOtdQ0M5zq+oSxrLipu/IGOrgRqb2M6I
UXikvAaZW9+RjynIDBWbThG7jQlBo3xZxGxuOGSfAar2Sv/BQUcPx0tO1FLU0sh6
bBYjf2V/Fz7aIQJaRzFo0tMCxLIAV7i1IwDyi1j3yNkISAxRN69Y3Eu0jkCMtLyT
tEUUVTGjhS15vOn+lRpI4FBeGRuIQpbRb5b4RToPY8GmSfbayEDqrNzUpRge67P2
C4Q4a51p29G/uM2kmwvEka2ZassWnVT0Ud6VX5RNQcd8qWoEmq/w1fMLCzyyJVDB
8Wuga4K/erzE+C9JDnwudpl0HSQPDtfUfVCZiI/qHxj91LPhFXPd7IWu2Tz1l2bw
x9SjCLaAaeUna/laicM9YdHGTwNco5nG+DNEHDCbhouBt9Ewv9h4i+JMMwO68e47
WAXqBrvSNTkEmvDpDt+ktr7nz9UHXlgZM/wRO3VW8l4NNGiCggpb5SEyr67lgwVv
p6xZV8WGjQuBWH6J4/yudM8yg3UXec8zkAMRcE20ilFa1wafTRPRHUj251g2jUHs
/ittmSTeJq26Eujeqi10lgEvBTjGdWx7M/QZtVLEidNXyuq1opCW2LMScUhwLaZ3
Zd6WxdmKTu5oxhKkHsIwN6weCkJFj2muPX9LI/WpmSPwtOEiro/oDcKpFeq21frK
mcTnsyYnvd2NPwnoUSTgBW3NeJJJQi3EZ7uvt79sz1ArhMGBUZrZuWT9EeLUaRg1
M+I69Rb1KUuXmiCPcA1/eJnkJcTxmx0A1h3bhSGMQsTGj25P7zNaN/AhCyyyQdH7
6QXCGVkyOUoctv1KuJwmvo0rsfokR4oUao0kZGZiHdYo9zKX2tqMyEfeeVAh0AIM
bOOcEJ/xe9eu9p+TI6FCqhITqBJYZSVN4WWmlFhiklK1CMmJdRiJFAUqL1z1Z8jo
OmR7AUzJtCDXWItxKE2agyZxalgGFEHvo+0w0vC+uS00sxo6uiU9CpLTe+w93e7m
5dn2slTFMvnuCyFHhbX/8/N+WhFqDicNwacefDGAtLUgTLKLp/Yg7mK2BSt7uJMa
OryMtePUSvGY5lTzPqVY4vxUGgoHZauUR+chPtYMMZlwWMBlrfk/XMU8NpyG3aib
V8UYh4uQgJz97E/ntQt5AxLo4mLIG+SJr/nfL4aXjzeJVoUW2YREuTFUbjtXiX5I
bmn7aYqb3vTA7L1JoYxStzlwBggek7E9zt03tmnXySfgXruI7SMjSpsmhSwobR+Q
pN1WY2zO0HMQ/pnjcHCOISnSrhwlMrH2Mngo4BeY2VMfJ6HtZiKdjrWGM+u5uEMo
r53h6Vw6V/G0nwN6MZu8ENeHbAa297XAWeE38RieYAjHzBwptq31it5bn7yWP4lH
3Cml0/juYW24wH1Zhfq3vuGE7xZI7Rjds1kNYjFC8E+P0V0xK9gGHJc5CBr34O+p
vDKmrtzukqAIRfC4964z2fo6Z8l5+zNJ8hXuLpgYubUQNX9ll9biwHN5EoTGe/Rt
iM3CaZaL4tRWkya9MRfdXo09AkTkVkxpFoAjzxifrm80DCE1miwbu6bKuHkS76ip
i17NqGT9TWLMzRBUuzC/XWKLkk9twsyVKbTJCMaNrvbX94XgW0aqDmQmy/7Mywvk
boHgb01B/JynrymSArfmrhAICojRsxGhmFrd88sTCIvsQuAwuAxi8okp5+79gmsV
1PvnVFO38vdkR7XMtUk0el3WohPUeH/4zRhj0ippK7H06isivK2RxhClOm8f7X4T
oj2s4dfI8ziV8CJZOmobLLZbQU+KpLtzEAUiBfTiT8atK/BZzjOOrp+cc6Ieef0j
B/JVAA46ngYfDeN+rg3iX+gWwKaaui9kiR6ZejTwCJYy+nJVllVNWRdq+j6G+wRr
PR8LatBxPHEI9G3pjVwQpm91SB3f+iPyxoz2YXzkp43L6i4P7DaKuemabncXVi1q
9py/q/T858/7fVP0V/cOar2kFE5Uv/T4pHcaClpc/f/v2mJcm2CacvooxZ5eRjPs
VhZcFKyz04pmOZ+QRI8se0xV0Erot03lrQp4vfSTjoBYImicF6Pv/A81XEaq+5Bu
mDqtlnItIXshw7z+Ba1v/Mf1i8PYbCdS26HFXO89VRuT4awQxnHa2SSlcW5ChDI0
ob8f7GjK3sT+p7ZZssemOVj8otwpvdlLZ3urTCHH7U1+LIH9pQ8qI4Em+/EnH3QW
hC6avt+EuDwUStQ1bHNyLvl1BtFvJEZRv5EFg8ys91WVcRaUMaBQw7RQHev9+G84
k5kPafsAfTwDCl0tSz9ZKV/tpXoj4IyXlSFj1pgcpEChmm9eGTQsccXTvI3IYYJ/
HT0nV5M3QZtkeSF5tJU6QcPNa2mXjpoey2ByhK5lY/U/TCybVReKsf8OoGFltr0a
zguDv0HgvN0kqBV7XlqIaG7mdhXZcemRhTwqR0Ic2wcEjTuwACqUqPvYvNs1cGEJ
9Hr/ML2Kv15QGebXGMDlXAqt9v5QT7fSJBVXPF11hO2fU4vQ/JNCeBeOkEwoLDTH
rzWejUiVqx3dA29lx8E9wDtV30s9zqmGBtF7H7PlctHprizZtosTAgj8tiZV7QUP
p4DXOvVl7YF09uE1oiG/FIBq3FrXPplAk4S06mNKUmHnmHFm+/I3L4rvmZUN5BJk
FDvpcT9yo3GIxagyCSnLrg/C850I71RlYG8GBSwRnsJuAlyemja+KEWjV7ad1DlX
m1VKWsGm4RqjJ3jm1MWaNvoBXLCatryBWpTEIeBw+LEOLL3fUOZn+5iIFC6XQ4a9
QEriSUQoeB+O1KGKYC+aGf/G/v24faiGPEfTLpdMgRb2EWRtua/QtmHp4qJlEPi5
pgMjkY12duHQ/rjOeZde5p85cmLJvmJEhuz2/gEu9gYuIVQKktgVbaH+jEwLTUR7
XLxu71s+fhGDtM0yuuKBSalidPJTsusqycWEUd8EUBezJ4l73bLy1FZWQTbtLWoH
ClgtesgZBe2OODOCi4pDaAlkf54jAda6NWqZ78O4BppY+jQMYmwPZXRMH5/13OGA
JbqOEJqXydJXSokRMjBnnBWC/w5pafgaK8l/EWrRrX7l3PalLbK4rNL8UKKI/rSi
9odExo2lPaBpT4LXcyOA9MNIqEQZ9OQtMzsaJtRkom2/BkDVnlb9+hOaipFPR+WH
eZQz2s65J0IwdKeK3/2asCpp8zuU9S2qmKZxd9SlsiT7WqFlo0u+qIME8xMLsh6Q
/B8ks994StOI4elqyc5Xz4AMl4PqvLmfYwGi5bUNoX5iR74GsIO/kQ+qqwKlCSml
0xgTmHhNNZ4+nsjYMTt2v3KxS+i8hfwVKEIyTae/pufIKF267DyydopbxNmAfity
dALicoiu2SMkYmsIaJlNx+l/IJNfQNb/kB97gkepKkYV3uZFbTxYKy+eKFCE7322
08gOo7/HA3qzm0SHzwGIrE2T03UVZUF3kW+0bU2uwPnPnhhIv1W8hKXd+QDQ592v
Ee33r4a1Hi8cBpJVnogrp0Y3g8bdsXdzT+jzfa+mnIbYz/EpP7o62whx5ZvPzs4e
qs8mZRFDBek9/CWtBeF5+vZEAkm6qv+eFYrVmgamWqXyY+xR8VqQGeSlhyKf3ojI
BKdd+xXj2wLQZYgCCUXpmkdG51qxWSjuajOrlxkgDBCpvj2iR/UYGw64HJefNtzN
s4t0D4q3aLJu9gqh/dLLYXyd4ZPZO8cNH3jf5xesmdabcSVcW4C66s45w0NdaNNv
UTE4WMdVWkh4tQ2djH+7e5Ul93Rll0/utMCS/sx6WjENWumK+FXUt6jQU9NrHPN8
L+FSbupdduw3vLIYksa6oc4db614+0Xf9mRcf46MkQ2Ie96y94+UCUKVR//6P5NY
rDGFoCu1UruJaes0frdT7/C65odgBlZzDulCcgpkJYstFZ+/g/EBnqnjqFcYybRF
TKwlYZPlj0vInowdEyFeEtYevvcJJGmj6yIlXTSvuszVV20M+n+rdhfCTuJh6P5N
RmEd4Ow38XiHne2vtK4YLFETTJyFKXRoMDPIDeGb5pChIGRC5YHXPBL1W8g9zUpg
16yiUcjqEPyice5D7xcrLEciu1npFKSmQyLhaHBQvVl6ZgEdBfQhxQZ7YdAnrxXJ
bPvQkYQMxxedN7ncz8lI5tHm/EbE+MtSQJkYqXmeVHAw5WHQfYKnaLd0xmS1Q71a
cpT7yU51XaSnp9nmyGcZLp47hjPxD4tMdhDOH0CS8AhhaJ6aTixow9niWd+Of0cK
BG752AvHfyvwY5+HFzr2JkVihfw8puEyfzpZF86em1dwX3JVkm4CWol2yHLjrDmd
pamPu0jIZhEfU36fmOpODql0mtudaPBuI9aWrz/onuUdnlGtPrRUlyBmlwQtryOH
dKgBtfTQyw4GtjxSklQiwbXmmnMuJtYVjjuPhkV4VdPZRUfOerE6gxwxeirrOfS/
EDbMaoqQcF5t5aoOydBYHA5tdWyJBvUpfQBCW2TaJuPmKxHsVB/8iT46riJG5tEB
WYlLQ8INauIMUzBRrLz1T/NQ0uTdExnWvE5ctJasKm4gcuPMMWakk35cWNl263TG
LGGRNS42Ogxlc0LeLwNmhnTeI/VlyzY+Y1wNTzz2kYcucnqB3MdJpPKtl8OYoAW+
Lvy+2NGRnM+8h2aNlcwuYjh6y8UVEFOwV56d5gEla0d9+H9FA0XppcSDJ2I96tLR
O39fLdQpn7JPMVm6JOkcewbMM0IsjPuzRNM6oBkpYKPcalK8vOAm09FauNip1FFj
lhpdcii51Y0UPXjH7oIMMbQClDhvbUW5e8kmtFquBhdtugsLuemtqvBrZ5B0omPt
yewxcewsthiQDor4t3Bn93fkHUWW3y6LvduzS/c2FTlC/pXSlZrhpmqi8IH6L+Z7
nnxUEF18Zv7+HiGluxamjxp83K3OkXd+GjZJzTa2aXf9I4ppmSu+7KK5wDrcy0Uu
VPTomWFgZgXNGFn97hqHD0tw/62XE835kkBvckS6f/ys4lstS3Mjg97cRORM13kR
Yg0uwFMs5XRFa+bkHA6Kljo97aiKSAPTOkS8UsqZPTzisrWb2n8+wFwLo6j5u7fk
nrGYlmD69Mz6gp7eHC1J44kzykITk0PSCQ1qLeVRyKPT3Ois1Sm+INtQO0vXlaT8
nFDgYjZITWCWn4tnnjpQE/GbcnzSmwjlv688tlR5EZrJM3n++aiGBrG8bRKN2hOc
X75otcZ+zMgnBGTAtwFw0ZZ9x0c9cQSl0Os5r+3mahS+Uymy2W84lBJAGOliqY6R
4WxIx8UNTwDrd6yHqfX5Cioj6P03XnWex2cnnjpGcw8FnSnbrSOvAmCJArGPYOlU
JMsdDHUnHZm17r9nl6RgFs24xRL4alXb2frB7cA8NUpLEpQYDN72d3TX9nhHpTG2
QdmtAWUjrBEAQW3ZYBkXOaVXODjtZnxyjUok158I4Rjo6k4dVukVrWOeux2l10Rm
BFaN7MV6dOVyCu4mYdH3zXVLj+87rvpijR22xsNA3xVwhVH86MtVscwk1PqfzD7K
epKT+614CwMJrwyF4oOc8RTAKdL7ZshmLR01G0fxctJdOupcK58nL3xpDbMB6a8q
fpQR1/rXsFKm9g7htJ03OUYJKGOhrz+E+34Er9ekdZoVs/B/0J8EX9lzfJm/o7pP
Rbdjy9D69rO0fi1rHQKzN5KKhUqsmSVMGs7ulFS7k02oXGAvUamivVjcC7rBfXEt
nYvPfPoUMp6v1a7ENj0KzdA+A1b65d53e8/yMvLq28twlFvV25Q422gXDlmDwSR0
46rIfQJtWgRo/Kj95D9A283Ql8xJlJ9y6ntRdgkg1Q5yRHqdd1hvhdgKuqR+1B2G
EHaX3ndGBX1Ka6FK0+FD1qugzVDZo7e1s1Nq5lHULU35Jb4mnmx2zjv1AkRUZemw
SRPBcZFW/XICn3AgQZTTALT/pvW/0RjKAlxHYTA/WMJf78nzeeO0D6V55lX4vDIL
bzEXCivWApLeAdVT6tdch6tVKxWWRsfLosLWWwBA+6IKDqUubco1+T81aD3+wJXz
ylMBc2t5/2yuGclk49C9lIxrwGBX0C1xBu0ak2VwY5rQVGgKqAXnZNFqnl3R6JsM
Wns8d2rXqhn4hpLJ6fPlFD9nBo2L/HAlf0KlzLH60A/xiqtA/DaJucGzBBGlbwva
OiUzctmo5DTB9abnVctJcyac8BLRlIB9/79jqX8QcEP5lvOWH/7SPYFcP74xJ/At
T+NsKG4kw2n/oDQZpi1SHmBQk7yYH5RNDyxS8aQP5jehEVdYDui0dMjZfawRRftc
KJ7WSdMrGS8qLyVrNZP0qzsPuqG/boaQ5M25ERZ+ZNT24u77u4WLd0lSJoOaL+qK
f3EGkC7E9PnVzGcYobMPEn5r02P75VLODgs4HxXAlUaGFnzBUOixeDl5yh2w/++O
tjrc2GbK1+tr+KKzomrzRhy4rhSdMxZXc5/yO8yekIolsZdZ/Jny6lqGzuPZRjrC
5tRDF6L7w7La9Nd0F38rrUXkIGDdUQKG1I9ifs3Whx6oeNELkM60EqlP+0S0dvVu
xr82QJaseVqVg/6MSkGyUZizhLMzNZa/d4vYRiI6cymc8QRqo/Vo8cnGIFkr3/ul
gLZf19RNmy1x5aLLHkfc35LPajK/Mg/ub4reB7RR94S8sfD19W4MgVYiXfo7se6n
wdxEwESFwVqT9k8nH1V4pub7s5NnVGQKETesD5pLvj5F5ZB3tXJGQ2jVSiZlCf8c
voJxo/WNEtW26UeOWtzLG3C93ddCPYOMCv043Yxz6v35r5si3YQFiO7KcHuSgxHo
4lkLX8SJBZf/6utPu8vtJwohzAp0XS/aT0IFKUPXrdpYOFRYOXSFUBYtJ6wNSb97
cz8bysQ6MukKrcxy3Dd2BqMV/nexZIP0sw9qSJ6y803MYmgq9Ysd2RCeZDzPHW7G
9S9kWXKXYYiz6KX1MUhjndPbu7AnHRCRauCYcqeM/atZNm8M5x6VyD4EimT8L0yC
hBBXPsfgp69SPHEX3DJ4mqJu58Jk2HvxqGxZOxeHEnfQJs5ObB2Kc2/LmVnrDFOc
b0Ov1AzeXaRPJh4joMd/gSdbi+ocmivb/RY7HkLnF2AlZOJk8z4kiDZ8pJEEKJgA
SjHQR5aF0JauH0TjpHzTjtigrJPpzUxfVMy9Z+QLoPrgjcR/KsKkAcLV53P+WIOh
a9SDCWcDdz9h7gVu8C0+f/NU9yrmYIBurrzo2Fv1GW1S4aj62VEWWkzvcq9l8nga
LqfKht19GOxb9G5PVxDVTrQnPzWqQddFdnZfnmXdTWObviEG5joWEI3y1HVPaNwn
ocCVCWcdqZ121f0ES27KqKiI0k2vS5BYDEMw1fADr+FulRvjhA8+pe5t1nUWraTW
50QoDHdcju462HsKp8AXwIs+T4mJ8wLK7B+xfJk+JQaUy0drhSJsZrumh0rQuSnm
Pp8rY36DnO1DG9/f2dwYvHNDMqU3HFTe5KlLUDvP2fkRbdK2QccCmir6Gu0YVqgt
V19Qo8wPYL28soe/9DRS9RvZmQLBMuwSO01Ghap0FX+A09NVeatJRtI8qRTITYMU
alI0q+o8gUeXiJ/IFbtP3hh/JIEh5zUCxZye/XrV73yuq5bZygxecBcdpEq3fU/Q
/vDRDq4k2MnmZKJ9Vvru5HdL+K9orRR0WEDyWNlwNHNpbWkuRd+D9m8crlUewgYk
53ZvDnzGMjatgmbMiLM7YzUao3zMa6F7cvzoiixkMVGPWm9T/yygNzPn5rs1BfeS
DzM46+M1YvnIqSXns/MC5y4/v5utS/Qvrr3Gjmt9p5c3HoIvLSEbZebl3VkVv+/6
1PTQqeKuJ8957m6fxs315gBuJyR4cwZi0ZquMbZt8Ic/L8HAENGejfAnCqff5UVI
ljFvBoee3CpAB/4fzyRBTKMisDclagtm3+dBgIuEND+3bkMKOd/s7ZHMJgqTWuRD
xwb1ZjtY27mKqYfF2bo0yIHQpaIjbHPWTHMZ86aK7a2J14Y6l42+J+6g84nF8z4s
VpWxYrMVzqQymCzRGF4Pf6yS6StXma7HfLQ2inXfcNmy+ZglLJRL52Pct9bg+UcB
W/WA/L/QEi1TxFgf9ExBWQ2NNha4aZ9YKA/OoVUnSmTQy2UbTmwTPaZ28cQsx+Zy
cEi0d6K96c+AzYQHUEoVdhczN4c/WyjpDKbl8s4Gmh1BsF4ghlfP0rdu6xvA5QbC
GOHg0MZ4qTJO0UOBtNfpyp6bO3llRmjV5MI9h+stAKAfsxRU/yknJZrErYeE+3V3
Bu7BlgOOR6b152m4mU3krzZibh6yrzRi9+jI56bG2D4I4ddcRUAYigKFJfPpZliB
+4W1FeEUhHNOp4jMTbtFFljZXFyGbpDZMED8E9xUvFCR9JEUmq/1TWXiJyouLDJ+
oVqmI3EOd7XUDP2sPvG28XplwBmWxbeXxrLoH7Z7siB5NOV2OVSCmU3qH/pG1xBw
A5KW+DWs2tINss1IAPpbIHWs+ODZrMUw53WbbVQDT9Facpr5vnlnNvi4Z7lPGFLq
sa72KnktRDQzqYenfFwzE9WWsqaNpcWS6UV6EsZtHIO8tGsC8DLjpO4qvGw3kdJ/
K2A4PhMV339YOpAduIPatoPguGvrlT6sXm3D7szL82kBo2NssMNES9SYnIv2NFUV
r0no63XYJC2ZOj9f5cjFwmI9NDzEDygVElSNz9ZobMVPQcIOczuTESp4P6kR3WEt
tsn55LbFwjeLd3dg6y/D75jidi1T54oNPEmwKaVaL4ScMUpGjmVm1hgM7kckjxWR
WakTL2f0Iiju2ZK15n670ZTcdIm1mfDeHjzGBNh6CP/2cHwWGmCi6kFaueS7pcTZ
WPWfNsi7p6NgpD8UngnnEdFUJjLVvu6NzMEGKsMWr19GpKFcmljMNI37FIgNaKZb
FiN5Rzq+SL8s9y80vgXGGnbeMhZ11FzFDYWUKawM+1x+tJwlB1G+Kn5WP0Usa7gZ
TY/Y/megDSk2XfCcCGvM8djyq4/dFzzxQDlu9vMpzOouT04KkgMG5Q0YXBPHdTFF
tb6fNmd7BpRX+Pryn7H01qogTtc2bDNrvBjAGvz3RHXzxJsj+QNQtdidtjXnu9pN
/AQ2A4jcD/2+1hVxyCfVOn/GXz9fnNaozfv9O0KCBXtjz91JseO2vIIFO2uWIdXa
z+hxCbZSVKqr1Bcjl4uR4TrRGU+nX9c9s1FoHIRmq2Bha7RqJc98T2VhZjCKl+oY
t22icb49J+WB7uiWuC83naCzUVOa2QVktt5GYEma5VddBhm4aeihmyJO+GHYCCNY
BsAYNt0B3sUhQKhkUKoNO3ausUYGuT3ka3HjgqkigMv4rutmIJJP/c20qgZ5qHaj
3y3bB8FXtKtIbVL7uqT+aFmRwM+7Dc+3ZVKuTRC9IJoJOtUp5tlGxfMyfhbKohmI
5zBuplIiQ4ajvfFxASz1GCEtGl8v4+ZOuIZrz1TfryWvmy/2dRlV2Ljrg+6gOat0
VkbV7onAogAqBxJd5EUQzNlO41NJDu9j+eNwG8olCp4bqVkzFw9FAUcHKRAht4qB
Jon4XyiwGpb5r65ZIpqednjzpf05DdqkqQ+tHFzHzoi3ZfISKQ0fh4Nvv6S/33GU
c64kIuxvmcGmCPv/0bXgDtzwy92hCVaBWuxn3MMbYyNQmc/wphKUAO13XxYMULNW
AVYTFCNBHqWbT+rPyIjFPJpt8ITd8eTFeqMBjHbVi8WE0icO4uL/v+lB8X23wWsi
Z7+DtS0hMRLXIG0gAdB/6X0KS3FCvf/i8mH59B9qaobJhjdZt1LasK5v733+TDv0
muv+MNbH8RLKTuq7DkDTQ8YQFtnVE76Jk6zdLIHF/5nVkjcD4PxkKFykChutJtKO
2E9bF0gi736ZtKj7GSTAe09z5wIwQbypzk41yJjyfcQ8jx6Ev0yOUKhrMNR2UVPT
WaDh1wFDiANh4jCFYHd2T8tMPexb0rVgVSAdfckngeNpKit8LtiyxW99xkZnYX4q
bjo/XNrNpFexuLl/quVpqjL8JAw4F12/hHdt+qLf8AGvDMJuePXJTJjcPWjaJiZh
yga2E+cRBCDN820IBGAPq5C9ALw8fu2+Dc5rIGqH8S7dsPJIlkY4j+f+vtz+m1SM
evAeyAfP2fWunmZnsOZDToDGYuJ2WHW30eVpq4zghNKNcHt6k/UhLzH91wOfNDQ8
F+5t6IuMVpscYupIkswdAN9MXdENYx4C+vRKFb2793dLOfaL6e7mB0vfIve0Gz3N
GBN7MKqPp4NwyNJ/TiFuPNp7LVAth8E3LL5RR3lnBJ8SlCdgWnASN70fQ4up6npU
j113Pg0fHUTjBR/0h+gfrH6JDuTwB8sVfQ8nMEY4BjSHWKU+bqHb6PONFdBUv4Ov
FxejytMhCuPq7rkSWISOWQUf1NBpxhCAJT2TQw/ptka5YIQTfYQ4tj/R+TwD07CF
l6uqGSveSfVKwRxsipWIK9imz5nS2RIuDkR5vKB5IkSCliA4cCSaFruz4ZYEHPps
w0MFFr4q9EG/2N4kfuVXKVGxoPmJa3+R9FCOt3KAILZpmOpYPkwol918I6P9ECOd
dAgkZJQZXHMqvIXhyZHAo7C4ncg9Ew2XH/sbeUsQET3tTXDPy05+KMhWcbLlBiYo
zAHelDSvxDcXtS21fB0t0fOTJhfIWtYqEE2feUBYo5Cgkxp0fi6uZI5ONYofBBgo
qvxDMTLLhnRiR768pOo8t6FVe0d3ZoIjkqcIZqSeNVzq/u+qPVvb7gQNly1pXbsI
WIU7GxGQuFA3dTHh6wSB2UAn/4KVmhvqMak8jps8YSoi1EV+9kRXW0lqQ7q6+EM7
Wv3lFHgsm0zQ9UPDVhquFp8lotvl0RLQqpddZtMdezrIV2RxwbJ91Q8m+NczLQ5V
AugxWUdttf3kjGqBnznRDw4G7ysgw9IyN4Hc4o9Hmvm8UQJmw3kw87ifLso2FmCm
JyGsEto49L0gReJZsAzhcZmgBxLXjSOJz4g9go5tXAm0ApeFWHa1sT5Hvxafsde7
FPMjOcDxh1Ys7gLzUYHK4aV6pky91j1q0B++Rgyd3UQAzmHbvuI7vuG/kbfzoa6w
f0mBKdJmLWKC7qLQ9LhzXbZM7rO5DidVrO940YDoSP37cG7P7rOI9iFKTJoU3Ddw
a+Qe0T9Cas5ouKCkYCGC6ufESoVpbqTCmk5K+V7z/zmkzJZpHG8j9/JMdMJSnijl
Jj41tE3i8xreU88tkxMi/GtTJRoLYiwXQZr4m6aHq+l1ms0Hn/1LhesPP16/Xaqm
1hUeirSCpt8UKkZKSIieN0GmqxaghYXWLZykKgr6CS9OT7xTAay426LsKjsvgLDr
WAw3Uehd7qwLGZeKgHWKr3TnRPzv925396aprZyben629/7KoX6pSMpeMKrHMqxt
F2Qx5s+WLa2/bxMPCfjE0jsvtPqdrU6YUwN33ZGWMGmMFRxdxMJgUomhmnzcTdzi
sB0+PoRmayigpB6qHvcajDfG1WQR2voBui3VHpbHXixJnSoj3Ms1cfEd2HPBCa7W
0RqQk1H0JwBfCGwE6goQUhTV/py3H2YOrRFdPtOgOXAtrjOicTx/RxkvMtRiAQYa
cv67iYZmnSbLZihdZax8ahGNcYi+/QHxBmL/LD98sFuMqbnOwkyHfnMtFJvOg9Qg
QwgBKYmiKmZPejNGyNBAqOuJ5RjFdcK2fe0hZKk4RY2mYmkHaBEtZh9VEieqUXtx
v2mjVfjGAmjAvotVpLleszwgc3hKXr5ZhqJXQxz5/bZbl5vv+grp/4i++yDS+9Fq
P45JAD2+FOvzyt/piBmQJ4v3LUNUxDMyiVcvtPSH5gEu5Mwq8ilyr7x18mRpnlVM
A2c+W53U4e02br1iRxSku1hSglXrppDWdunV39PiKik4R3pxUArhdmIGrxmMCBpv
eRjgdrpCex6cLwzDrR5ypFDstgvx4ON0tN+G2S/KsqMrWCrghEDSVRrHsREfxwBP
HJzG7CPj2zSASA8SaAtaYrh6ZYJBV+tT8gWtwKeRy/S+4v0/QwSSO/hfQ2UwHAkV
cREbvfMjCLgi/SX2prMKW1nzVj8QQvZBeQbrrliijxQL9TS4fhjFx6RQVf1DcgYZ
m050AXHVXNncTNkHU1cGsrUKWEJabktWC5CUlzkpApwt025kOw8XSBtGxc5BAJAJ
vp//2UNp3hJdmMJVONHCvYWn210USUxbEOlEWMxJZJLB0Ft9izl9DAZPnUUKMnxz
RHGpssVgPiB1pmvtlZtUTX+clvMClJHA0YCTanVXOPvGP4qkN+eyzFwYlG8q9K0r
O2VFbsEk0ZLvenFHvaT9ZDRTMc3DLYS1J8voPF1QF65e0g4Uoh7M57U+0dpbJ5vJ
ACidSQ/hAquWMhc2jo6f4ZVd3ISIrR8G2JwdBqkiJaPj6WobQRv1qdSsp7+A3B9F
Lwih6M2IoZVwsmznQhz2t5L3BuwMuFZ0BcpVVCW01mVT+WXl6qAbUu+RZ+MkDOwO
FsgZwT9erixidF5ZAJQAiFZ6PkWopcz0kVkzzPkadoIytXmVLpy9nVtSpazjK6P9
ocsAKTHfFFx1enGyhrNWDnbGEPTEYrN+TYlm30KU08mqzocN6Z4TjuaEibwm2wv+
+4IlhmZPW1cSuHGZ5zcimxccLyl19u2ttu14f6nsyp0V59kFb6Vn0y3WIK6QU/Rr
swK5VQPDc7k9pOU5jh0uW43CjoYOgEtThzCYdl4i4sQ+2VsB2pWvD+aX/nSAGxc6
rQLRDrbEtFQkrvT8qSK9ZGt/AZYwm3127wdJk2a6hGowhuTawCCn5k3WiCeXNlC8
/ds4lJmd4ule5iXEBeZRj+637ycbPBthIG9gtd1bY687qLMgE4gpPgqaJ447RJbJ
1WzHhLKK9SreGHxWGf6NIy62+3C8VvgURZy+VEzVVW/+iyumTD4i1N5foKVUZKbM
0Se0ATqQv+Rf2mIgkr2CEvLvPRZ685xlldnk5D14JN0Cbt+33LFbDD8LENrULQeI
bXx81QGLPJNAXLCt0o9SqzCGl/s0wMXgwGzPnmO63pzoZZqX3pg+HQSo1XtTIaPr
P5YhGdITqa3FNDSAClfs9h3OCoLypHevNtaqje5wi2SFPcFk4Qb10AIZk7WeaWBt
4CCBOeWI8WtPJj5l9hHNxFzqPLXSqIoYfuvX5iJII6wctgerBfH8Br/j00TIaN4L
4FMLw4Nps04Bl3bHPkZkm/65egWNSOA4xZ8njfam6wmEYIX/qIjNm1yBYbzSv+Cu
kM0jKEm7KErNw+oZMnu1BbSdlbCUyKAFsNUWjOTiC356sjdinJdKORoNDnCDqC9o
20fk45lSBkIYOunbf1RnxW+0NH2v/uZtdKhFgiEp674bfqg+CJAp/okUiLhyBKB8
jGRy1XTaPORUNPB0lUnTpjWZS9wzWPHIUX6V/eA1emmY7ZV1XcfemxVH9MBP92Ak
6L2ebIVIQww4tMnVBchT/LNiFQgS46GvwL1yG3VfUK0hiCc2E8INDL3yhtaADM3b
fPFlpAlQQkrhutoP4R2X5Mo8avBvp/nFekDlqn5BDbLstIpPbREp1oOEJa1sihUH
tDncJbLiwxlLhrMCBhfcZOsE0Mnt1OWyst8I84sr2i6HVCdZQPSHsep7Nc98fJi3
yJwQpdZxUAbQHgiq5kAmhCcS8MWQxL58S2i5MJcq6mo8dhlcUY+o0evUz9x0vKcP
63oXJ8aYKC5nSEAQcccHESBvq/3+HCk+GVYk8nRLTjidaxWtvmk//MZSftA3fOVM
6n2spdb7WG5LB49GvZEBY8bSy5L6QzgI257pg4YG5VQ=
`protect END_PROTECTED
