`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TSGT8rRNcbcMMqRTJt9+WJrpLTU2TtnDvu1CRic0iBVQlEdb33skADiG532Xrkd
nOhk1cTX8HU1AIXvWIsWW2D+1vBVqjyXVrYPFw3JYBHfNjF3+wLANahzrlrsaQhB
A6Ut43fQS8cVAbvnw+xmZS3bxkjrw55GO2ovtUAjZswF9v/2S1jlwz7gRywkYHWp
pnWp+jQG5hzZ0rE6OxxAADUYXajl7IFgC81qs+luiDoDSIBd/erhMJoAsm1fMujw
zWDLzEHwEp/PwYaXUcI9C1AMCy3i/VIbGqyegSVBNTg5hjvyCLDzAUX7K2wIlXzT
+ZSpvfzSwPR26BYVGUerjgxUJY1eYbwjohEhdIvIOWPJeZ9LyHcozEP0Eenmpvot
h7wKt5t/jY8e3DWYxDONrEthBW++MOF46b/RQPhOajGP/L0O/ieCYUwoaDYM06Fz
skTAT5rFnYtbVcVP9Phsre3JSIXqXfgvskwIyfvDIdZJpjDyyNVFffRi6mSds4Bh
RX3lxax/0oaCwzBaE0FCMoenCo/pbtwxCNGxM7Qswb4IIKoYAB/F1Hnwl82lOPes
hJ9jYXhgzkBu/S75dB/jtEUusF6xlNlyZO0DA7wRHP7Pul/3dcQbBmL8jV0Wooe4
9Nsw4UI5A65fBh2i6/wB5Q==
`protect END_PROTECTED
