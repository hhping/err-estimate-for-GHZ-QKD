`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnKmIz6MZPDx3nUHYPLfzckwRlVzs4sLHAxFH/Ij0Ie4bdnHstbMQDRJkBF8TBve
kRvuhQMjerPCD/g0fv8A4OH/OZYdHMRGTE8eXQBYhaLEWXfqixsnLtcQ9nbSZ2M2
7fCYYx9EXecK9jO/+KYNI5lqq7LsiNuVqf2MS9rCeMtmwAW3i353qwW2cqPoXMxm
YnMWTxQhZR4rzVFX96NZzFZKHQJkHtiwUkNy18lfPkS+bbFrGUrwJqtXvcpFmEYE
DdAZoDUYCaBXg4ekEQBXbYT5t20nhpFMzWskD4Ajuul1McFcztdwqfwmekBvuq0S
T77GrI4yMXfYG5/yF1tyLih2HArJPBZeBCFyNi6rDxWiDp51PoJNyj7jQeLh0J7E
V2HkUCQscBqq5rqSma60PKqoX1TSDCcdJ31BdKJ2z1vt+UvTYRs97P8hqxD50nfv
kK5UBBJfVVNTt+XnoC30Ha5kaHYkRyuSv36L9JTSg9Pa1Z4hRAG4j7VXKcpi09ig
pJPPThUNleOt9mEHoobFWD8KthcXI0+Mh8MyatSZpHRAZQXUYf7oSBlvzc5ovShU
hfpCDg2JJtegeA/jCMQ0QUICkGfAkeSGmNlRLsIUFuvQ9vBPUNzK7bUuBn1Q1Yza
sk/meUGZFG6pPWtQjNKVlOHiTJnYh+Al1pPdK22W1TKAhQlOWk2G+jQUL3RhFhBK
yhpkqp+kw7ubnqD3vujNifot8CkOEdOasmlWUj2qkKbmNWOrdjauVH2tjkzWlzHb
H+WnGFR6rD+tx+Jplc2P0bWCPS2Qp8ix5ef58fmA0YDrwfqtkiHK2YVz58zj8QWh
fCLgqykRriOdEeHqnxcLMf2y659bgsQxUgjQ7YAvq9LJgOtdK6gqxtql1z9S7azp
ZmCVgtq6ehG5xLm0wV59Isd3LDfgT3XefBWAeDuretFGBZRpFgYS2rhW5cDhX32Y
m63aPXC1Meh6XYHzMbNOVkNivONhTEHQj0NEqrVw05gNWenP40TvoVwSuw5hsG0c
Mt9jOuoqt8LAMhXdGDu0S8i5XYBm9ZPPsPfM5uMOltP0SKb1AMD9/kfLY+cOVxeA
R0TPCthiguSpwDApq3uQeK4Et6zgjQ3TivjIFdIt4eMj1pVmfv9P8z+bIVN/X7/a
e2/NgbFQz2ech6gamjgKqfOOhv7SDkEAZskLz5dfBpx6TdxpmdmiGse4h8B+52hq
SZ5pJ3KeOA7XCItzGZw+XKUMprFKJx5JDdRBPQPNE6UWl3bfy5PdhRGC/gvJ7Z2G
JGG4Odd3sP6Vcc4q3OBrIqfu942jw7tYxb+VUdkSSQNNew8LZj/YYD0QN4WmDMLJ
rA7J6hLdS0usPKH9DIphuQVhKM6cj2pwrJOn2vhLcdiKcZH2HmkZoVDKaxa5ji6V
eu9E8sGJ6aoyxqNO5Nmjj6VIZRMpRmHYDRlDQXTB9SrV/w/LeiAj11CeVuvjhrpU
yqsxh7fA1xsOi71BxBeZV0BmGz+/P8AREDKIXAYZa5R92NJY3QoEonjckKJw+B3b
wENbHicJvtqIgHixQEW7pCTQwpvcpEO3fTVtfVZ+ICuGjygYtrFIy571U/lG3mg/
85H+68qs2mBZmeoygeylABD+0NiOlNd8yaRsr70z+ave//sg0mn9EZbZ1++eQ1SD
oIRm7iUJF3n3mf1ZE3Mjcl0Y5qkz1Mvak5eGq+2p69yFzWeKKcC0UedYEPf1f0CE
utjQrkVKzPs4YNuouZKdlI7MgeBkLgh/BqYfYsgdCFiuU2INMQ2WitQFO1donr0u
6XEWq96fUpquhWVqeZkUDvdxRe2Ds/AQl3+lcXsF2hlqR+Eqt8VYq3smjxr66Nmd
RcvciHescJTYxrzKnKfl8AesJJ0PjrueDdsCcJbDV/ukFCXNstq8EQflM5eyILSP
23IerpREBt/jKLBGCxaA9qHnS/t/lKTy8BnttTJAk1+njeXWeIU4ZVleLqrzt0YQ
QT3u/Fyt9hFsw2eOWBQxcKiuG3uQRKh2T7YrKTHzIbeAORJB25A8ybr5ZXCj+S8S
IKRJcJt5J1GmlgxGnyyLpnXJcNjKoZHzJsw5iaCfjzpdYF6Sqm4QuKRXOLOc66fb
ubfIIl1sE4fHkBH2E5gdU4vjAQLJ3qFD/cV8+em1Mjl8gQNWNHQBg0dtffap7rtc
D9bUBEEGj9EXVJi0ufNWQXsz/siiMbJPtBB4qawWlAZtCvjjETY/itSstQHOE6h6
HPyHFtIIuN2oVmhiRfrXTnHvrhd7PI2EJ7AFS3W64+3jx+lq8aNJemk77x0FKSGf
/5PoNERRbiiwFlJ+SxKevoNVQ3wEk5xcXClT26A58O3LSSAaTML084oKezpKgiX1
sF9HO4O9gd8qDsqWniT7Taz2WAj4/Cx2HiPfJ11E28dEnLjJBE/SRca1jehqNmIj
WkEKDe5zZYX1kUFhagdQzH+F/K/0P/cg03yIHg9U5XpFbCeebg628aV8IozF6fGP
iytjJUHUaUJ5PpNhirm3+WILNRhorprt5rWPCJWSL76oZhuw8IxChVKRhTd826jh
HZ08mNgqe18oX4YhaW8C9IqVBsP60PH2ZY5MxYAZDfyqnPw2PSFaiIp6rAbkmc4j
A1Cdf1CtKnW8xxuNMMnH6ekI8E1ogwNF1UT3u7Db5H5VXXoz63Jukx+Fv653Fnvj
/ViyuuPgrGxE4dW3BHadPipYrdHHtdmZYugJegXYAxU9X4VVZs3NOdE9rEvvdh/u
LmqFXS2YwhjkEgyDByNbK1DfDdI/oHNcT0ozIWMtMhjXose/yef2mD+Q7gaVXY0H
9zmqDCBbi93tfOmXrMkvu2wyJcLiyKNu8/hK2ujkznAexEL7e3RNpWSbxNOTlbZs
U7imJld4rHbA6oc6VxlWgTbBIcH0OwBKBz9nrWJUTaLK/u/+UOpwmqYegbaFnref
IZt/+ILJhMxlnRrXo7mj5mSny94O+lmML4CQe6reHoHg8MniRrtaNrdxg57qOlMb
R++0FCXL/nkxpCqondarpJu9iVGLs3fadpCOvo1IbsGFxiQ5bKf8sHOm850o++M3
xZGhEOnS+I5M1qjaT8Dlf/Ck1lMj7VjwS3g9xYNKWa34aQji1aEWytRmdEaQnJJf
5ZcC9UT4JaS4Fcd/3tzF/9ZlZFnkzjv1sJtGVgTBV+qAfTspfkYtLxUjzp0qceFA
vVVWJY0XHuAoZWlsR6X5hOP63q+5tv+ZI9b3etNvJjsXDHhqXOgTk3XttIjrJ9ON
leZtDmGzltvZkXdKCmPwoxn0n2tAmfkqTxh7b3kFSZJfK+gSQ58f73uVX7nCrGGN
beZWtCvaiZhV7FRhI54TN3n7bLMGSspHi7baeF5kCU7uRGZJLQAXsZyjmMEH/Xxl
fwVRS7G0zbmfv8BhMxLUmJj35cjyZlxaVuZ5kcGO48PdvcRCMLya0Q0Aow4wew/x
rom20n4J4Rb1c6DEjYXQlD/N1hqtUhToymPskPxzaHlChMtETg4q6BOg0mMc7B1D
WSTxIZpWr8xgXMzkw2fczmLTCn+LHVVlFz27lkS6YsSckP1DhL8b11fmZYrHQQmC
tvCLzIKgz/ipPdxAAwKSAqs3hwBWs5F1/Nbe5X0ADYJG7z7CVbviat++6Ar5f0h0
A/PLCktBaBOjO5u1Ve/nzfMsXc6hB5ZEpMJhuaDDtw547aVeTZicNDs52IwU+uA9
LQJU7so+Z9TqOhNHSP0rue2shy1nvGLqmTguM8tVe3J4d42OawFau213UpOFf3wZ
glnfQ1bFiQXTQgBkfzNTFwv7mTPSR4lJmDVHiVEoH5S8508A4ic+me/Tisn1rUSG
NzLnSjFZ2zWaFzrD3toD/A==
`protect END_PROTECTED
