`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Dq1hXge3VdUH58bOQU+IflFWm414xSXKH3xGu9GFXT1KsnyMdqHbhmgZPVRmhWq
BlUbbCSFBI32biUVXGyIWGqvOg8iHhsB7GfxfW8a67XBtFN9KUNBqX57SheK+jJt
I+wGUq9QfS3TMYJNbuBay0LuzdTqInRBVmorHslB39BcotwUoAcnDm1hATsZ+5kS
OM0wumM1zl01Xjn6GalKSU5IIEU0NpLn1ZCBtFbrJofiu5JBhxcS6XCBPExQKoNg
ev0BbtWqu61K3rzlCKGYvkttRBWn5Fdz2ExYO35WZtw5svZd8w/rrhILeXV/BOA3
Br2GUGVdHgjnxvZtrAtJFOOLa7SVSt8x+jnkY4D/06rhYi9zmtRkEI8P0IYAGDLR
BMnL3FucnIswM1JUFBt0PPtRhGab2xSF3nilW0Tz67s=
`protect END_PROTECTED
