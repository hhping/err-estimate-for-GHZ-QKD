`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYtG1S66AQ0/BcVECPtPSUo3SmfLVzTIn+uXJPwfPuHElsvNsM9jvxYuEtqMm4oU
YF6GP/9xalq993epThVTBZRzjwcshJj9qFMvGLHHewzceg5rUl9KgGkP+g66RBJ7
yBsucJYH3O1MQEcrdDxR25Tcdt1WBhK5xONn8Z8QWOJ9HFxyXQf8DVIybZzbkBnU
UNFJ86DFP1hRQZ4IjXqncBUhjinI4XjyJJYt8UVhaJMt8Ax7zEnN2ghABbKKyrUL
BMfomsDjaaig88B1X16xoqlJwqzJNXSBpeVc7NmqdFGtuNUDBQMFeBwjN/LgRzr4
5LJ7wdfGZlRWkC+ZtekWgUwPpTwWFrce3TlaqpdO86Hn2dTS7dlBtIphklKwjPP/
3gJWDGLNnvptE7Ca4OVQfFoPZUoltcobeXJGN/8T1lqDbQzg30mpy2QEzbKjvIWK
nG37whBSt3PqCqikiBV/3PQ863JSqFoMJfzC0Nh1m3CDEXOmyoa8YPt8NeYuon2N
ZyRYOxBqcqcjk+tQALIAYKdt0ZV65CIvuyM1k54D1TiN7FI6XPsOrvDHaUhHOYfl
cV6+vVGM0gSeHS9lfOxSvoaifMZCq2717O0IcMPdYozOyM35bWknU6NK4kfSGHyD
kw3LQRZlRkmdSziTFh/EMw==
`protect END_PROTECTED
