`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Uk0DNJrzPz+pRmqUgYcnjvH/S3gaHP2JqXKDcoIvWkyiZCg1XkbEcE49JfQwTf2
zwCHLvp8zQ8VpmEHeH/qVExADafBT5jsjqVFd9m+EQDpvXUr/p/15bE+7GGfyJ2L
aUVlY6YnVwvhrcZr2QM8euPnfjrNDzt3l5VInczk67BJHtoBmI92J5bzT6gvqlRI
sG39L8BnW7kdydEh9f2l98qq4zprLxuafy/6lgmhkqNZ1hrelDJZ5aYXpvJYUNZi
Ow5v0+gUb3wRR8US8gQJxjDvpowHQLf/NvxWgBlAo7gfAOAsU+8mnQEoqZnflEXS
7Cl9srhcrRK+9PBt60S0KrZ5ml6sW5+BHWJPfFgmer5OMvagNYhJglxoaVuGxe+m
586GdxT0EjYNsRukt9WIufr1g8Zq2alY/IuJNXjVbAnKmYPbQL/rgKiGDsR+Pzze
HpsnQssLKrOYeaThXert+X5T+fF1q5M+VIeGPR7awjMAjpwTBSlpDdgDMeiWkO7Z
`protect END_PROTECTED
