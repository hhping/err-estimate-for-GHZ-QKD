`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8ViLz++Dyp+/Mv6j29WvcnmZtWqT4XLSGZORquQjSK7t0U2oVoY25gte5d1JctQ
hDN85ZzKaKWat9la4gPMV1OINLfHmHz3sKqI1RtSzcOfOtVEPfZdTt7FFfQ9LXN6
YJKoBMKst5+feNcE4BS1unvEaNhJhTxkllr7uEN2FALS1pGUzPTPUcyjpBSbJUDj
RyWTTyAzZefA6zeJfZPNfmAJtWUjbY1ICaq62vCgCUaR3l/WZYfZ6acMkiM3zCBH
e0tLtgitJo5zrm4t9DOYw798zBznQ76J6oDMRk2/OfEuAtZSpM7/HZizW0KPGJqJ
SkOBmay46p0tqqRqdW/T7ldUlqXCGqG46t1Ayv/0L1A/Bk3/1RitUXvXVCFUtItk
tDMB8cKRo1NsNyshaQgPx4NnhCBqJYf3GgLNgAwEEcEzuqkFmWVV9TTMsSJNwXgb
wbIGeaY17etm7+tmz9eniPINagEOC3YDpUyhcc28VBRgGxDvO48gk9bqjbhQGSM6
OCH3Wy9C/eWcXde0VOAQqZgWnlFoyypNmAt0L2N4XupHXZZ4SZhjY/kQQvjcoZJo
N6U40IFTetunI/VJEVozzNVbaKKmxY9k1CdR80lShyvAl/xyeusdaS8vQA96ngc4
CZxjS1lQKWDdBfpKRSBmnv4h58u+vIuQ55G+Vnz6HcLZPXaTqkx2GMFawkobuFnh
IWnHSycvicnneanOkteK7mtg+VdJDYQ5G4Jn5lkANdPyvLSPlRE+LUFIBsuGIyWC
SLPtscYnDlJqgkqfhkPF0J5EGMNu3kLEGzR8smOmQL06vk+Ir5K2fmzul8/pHfTu
Eup1sCrNwq+4nsE+b5TD+fX9er4YC8D0oF+WJrb1gFcdwfA0ZqggaAEAMmEEoHEo
r2U5sC81J5MJH0p2DXh8tz+BbfBFpuka4GpdqrrmtYeKAWtSPjDmqKlBq3DfV19z
IALpGYxtHETyE/pXk2C1p9a7K6G5skE/palXkiMmh1nDD+XJ+WDf/D/yeTrDSqLV
Kb+dbcdPT7wOBs5MjWoTadlY2dKgSzTKIrxGbvx1FDIb/8OLWd1LpBCZh/jL+jXY
q/1ulK/bp5FhAQG+Wumci1w3NI24/y/bJ6siS4krkob+o2XdJ4dBu2/TRQYqeDIZ
eM7qivr9zCEFOjApEV8+QcUGmUHd9/7q4fdgty+6EVCYT6vvgetL+ujBX78Jp1jO
9WPbczOJ7D9iWvC1rVbvaqnQiJJdBTMjgSCHjm3+OiBKplg+m5WPVVVR5vbw+Ytl
x86698IDzk4c2hE83xIeKLDcu8PJTYZ7gjkZSnJbuCABFL8WbvGkojZKlLTenRGo
8Afv0qTqrN6SvASWcSNf4ogt2wu/E4zbo5YW0YCDRRYkkrG2YzIE8izyUorjijrb
vTLO6XN4piqVFeNvbaMxleRl4iH6I7rKieqqN9VLw2ObJhf+RnVCbYKS3tKd2v0w
0Pscz1Xp4itIYkTckjeZacFx/30SY3NeNzn2qc8RZDk10jRz0MIXIOnRf/aKOFsI
0rmh6v20dyUlig3lS49isrW1D1j55zVFfy3LYW2qcnKTJ3kWvkC1Esm2Bk+B/i3g
CVE/xTSUAs3x18H2+OfF8iy2cJ6jqbBbdbm1tdavcPRMwpEViVOIBaH5+w9T+UZm
CGvfLjLIilZzUMmqQNfQGMIXj/Pk9jm+9R1cUM7mPjNZrnsiUvW00XpTWM588Lza
cRiyIVm3M0JdQRxsvmVg9rUrCIs/jtPHcomy2JGyIkhkmJadWGcpDpD+hW9HIwcN
Kgt2W+8PM7Ru8Jp5HJtvckaVal5l44heDSPv+D3/ahnr1V/HzAPWxn0UbVnxiHJs
RtUzxVzrwYsDFBS+ATqyNWi/Dvf1SqyqS7WngiYQy4GViiDD4jEwqJqye8OU83hW
fau+5JNtRhvF1hA/7dOgHSoI04TgikpfeTF/aN4eF7nSl7dJHIsmcYSyXWYqfy7I
g8JolJULcUFQJcxf15jd1s5pP/QwQqm4oI/PsvelwiLIkbVn56gHtnL3ilYSLgTN
wMAlbPOQb/vEgK6EEYgf2URLMjaLncrPZyS8XlT9ZyAnqyTToPfcq+oc8pO0JoRH
7oqm/uFYV6V2c+6mmmlDfyGRiaRUuGAl3zYiFK+j4oQIFEmfTlsBzWpqqva55gk7
Xh/aHBLZATYoN2enDnHtM4jvxyyGXKkL5mHX30eYyd4Hactsj5Ini9xWFXwCk5u+
2cEqULvzvIh7qL6US43pp7OdMLvP6yh2rVm1MVkoz2V7rFQ57wRynsRN5TsNISSx
9RTeER3hz70LMrAC09YCiVO2uY3TqkNObjXwv+cghprzKImj4cWkcyI8yS4MzIG2
3skh1coFCmhimho2JzrrczYZqSVngbxnwObU1/JN8xtBOKG7E6GoJ4cMaU89r5Wv
LSRPrdfltjZzqWDBQcWz39UjJdtF+yJYkNeHOWHaIHHLV4YYsxGd4VAfAitSyczH
bU9eG3fYE9OjP8CxmaWDNwLeZzrP0UCzcEgNQ4t4P2wxsWLfHxQYgSUY5Y9vvAQ2
cmWXN5A8SpJ+dpckb9vJXCvcUaGX4znexUjX1WsYL/i+1cdejm6tgsAqVvifnGcL
HuAhwP5yxYfkypDwOixBP3+T44D6a86YyfvZtQQkNEqItm8Kf/izHst7m6X43udX
JwSYOsjXtgwkR/EjVKyWwcjgWYsP7mr388OsqmeYble5Rrxa69i0nBfcBfxwIWwn
+JuNpz8VGU/vWyrFTTytflWQnIGWqGVxDjgCfdx5znsP7qGGn1dXEITq3BnbqdV3
+Bp5/bv3Yol2GaKRR06zTt7d/6vk5MFXYOn8CeRnG1HenTmumzATHWjincNlgdT8
NYEapnbPQ3Jnj4PrftP5S3LHbuHpf/KxPkmJc9siS+Wkns0FpRCJc09qim4vYxK8
KuzcqwxkKcU5gIvrCC/oNijq07x3KRSJ6k5yqukk9Gvo9CHtW76uA2H73veHNPAw
UqeN6WUaW2lZXKwkkZ/74aXxeyo+xsCRuVnnzW2C95LiGcF6ODzJDn9yTXY9TIZt
TmZuYNUHCh7LIAdLr0HPSGp7/t9OhU0CbVAfXAas9VAUGm4bp5lOONOUfvK7OOib
jErE+x1WOkUp05a/vGF3A9wm/OyvHcmdTC5XkWTqjMD/8ZtFbFAIU378RtA6akAD
VBoOiXQehl+9pD7OPf9lgZl8DXq1z7diPFHTwY4bG9Gn3gzdc28RxKE1tXXcittG
wVQDAJLkZ8GQSCUwxCC71BXV+mwJp7odce7NUbXBOgJU20vmxpYVu6PfpEGzTKmi
XrJ6gEqihqP2aw+rlrW2IvpDZdNFWrposOwkkbUuI1le6e77xG9zcped4pDObuzv
nLsnLB7nZRPcQxth2gdb3w50C00E/dNRvmH2Kgq+jwrdJl0a9EG6/rgVdvrorH8g
NVekVyl6UOIR/eKtSvWp0sKR03MVb2tqe4TPnxGFQKImGGxUo3UiKb25x9PbQHh/
EtxOTp5daUlcULenaaiw+7Hr+HltjOtsPbulv/nt6upxy+dJnYzGrlwH9N0ivK0F
if8yLfz2ykvNLnVCMWCy4hAbs8Nr96Nt8x0Fvo/UaCyZvKQDP2+MxsNN6WLMjsmB
UHW0bBM29a7WBCfG1hsqdlyrohLjvNtELU6JFDgHqDGOjcavanixEwEFMbtJDUjL
xWoXy5PDu+kexFMbij3YlzDuOWFk2407ybbaytr8oHS/fN6TtUNIoPDbAD+SlzLA
CPgAo7QL6b7G+Pky+owDu3Y2nUWjkCfoQh0xAo/BiFzC/3Ji9li1MLUxLJVIdqxz
/6G+BehaQjNTi+S+T0MwCB1XZBQDe62KQwDXQEdly+H/4ujQz7PxIMKrIAfUg5aP
`protect END_PROTECTED
