`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqACXaftYG23iWGJDebI4D8PWhlCwns80TNP/rh3RAQWfz6eAMgBgZiTex2liCQY
pCZxnVhpCN3o5ghczeCYr68T/ckco6D9Vu21aN+eY045q8Ts+2cN0es8ko4ueXoQ
dttihQJBaxT59WmI5z4ucEh46xufPstaGgCExyjrXeIB5f2te8ChpyRA9SI1f4Nn
Ecjp0w5DnFFgkXQxZ8n+SzbTsSjSVDYC8AnoWaUDXw8hUyhezaWZzlBIBXkUK/6w
jkzOnz1RZ8So6fscfvcmMAlTol6ssFyFO30NLkCJbS8mAo1CKoFpzMx9W7daljEp
9+bm13AdVomBEvv7ksyj5HN1ZZ11XPOkDqjgwgv62lYSUz7cVpJYhrAO1vFnrkk0
AlOTcRkBrz7Wxmbi9Rl0iciLGE+WUHsAxhvdBSqqOt03vXltAhkCYVCPN4xo3eq8
2lNNRaZJjqXzknX8n8wHHFom5Zb2//oXyXkb/CoO4D17xVoTdzfSOi9HVb8jcqwM
PiH5bjltdeEJxMtzUq/z8roZpC1e6wko0ay1fQwfFkgnG7taT6uGiM9F5I3GJcy6
ENUlcGrJzQzYeJnoiSFza01rjeuKeVLLFFy4cF2OL6vQaRwEPrHxrIOP2eauF6q1
H1G3wwWSfotIWW40JXLAxaAkTD2BSxOMZwzglyu6+u7U0gKmkdxbbsweA8hzI4a/
a2PKIb7NHBcl0R6XLrQpQ8AYLibwJbUVchng4WJk7X+EfRQQaOXb3ysIG1mwYIUj
AtkBU/M6QbSGyspORp2ZXKjzIfDERoCurlY9laW15jaaGQCUd51VG5PLSGVKiGb7
LhNkyAQ6kDw4skUNoeEUJkhb0p/4QutWC0OgqQCjkMj1pD0ChQRQMTaLwda0ZvfR
ffbivlpBUVbOLb/HyhoH7UhJ3bVW90ic8ia4Y9eOv4BWu2GeSemfZZc2ppkc1FnY
5aTGlrtMOze4Qv2J+6n7AxHkKKeDxmEQ0VDqgmg+8O33QfTC6x3wprrjazfYXi6D
SO9+G7sDeVB+p5Ywc/U3OPFbQ3pQ7rDyEhiQ5/yGdrDPeaejvQQm//f+WW8qONsx
rPyxyMeo6THaGIJ6hfnzD5++o6opO6OidSvNM56DRHZ2DhBfmcoJM+VviT1Mg4gD
AdwBlfFmdWpnNGFgFF50ODR8gii3Y8LRCBuU9MKeIKljbQWOfGeiEIgwrQ05fqKF
YJLdsmJy8L8W2/uKdVkN96G8mFdRTPSUFStF16SDDF8W+REzYmfAX5kJNV1tdyRO
4SnIdvhBGFgFe7LUZhSPBHVu8q2+oC3GwmLMNsIlGPF6qKYAQLk/yATwqN/j9Z4w
UXbdVKWmCGOSzQGv68EaO+1kPnlVfn0HuditG6/6wuJSVSXwXWF9bww2TY3Ohnpq
yhJwcj2xD0ImgjWkxKw5+krtL2tDDR/j6npYaQwSr7XcJTIapdCo9SQeraI54icN
FujpdM2GN/OFuDk+etRknf1tjlGjKhDjPTJcRmQfg8zmrN2rRPaG+CaQfDnEPWHo
1Trhgi2RG6xEOtjKVZeNRXd46sb/U+xT8P3pAmY4SibvZcgkAKp8iBhBRZYvr+fh
iowGRn4+a1j6L5X2e2Fux0+M7UCh91BT7KSq7YkJfwLXBFacwHppHZg1MeHHiQnj
VbXBKCZISudLItvbRzooTsJ9XJ4tDPSpebhBkak+N5NXhqIoPsvdov4zYZx3XjSV
zogKjyyX/C/JcjB2S5s9317hJYKcal0S2azjN6DWmLgkboUa6t6SwyYNb6eCp5F4
1SZmQ3vXzJqazHqaW5AECioq3oFQTTDjstyTRD4dgcuwth0xqxp3MMrZNPHwj4zn
H6B4wZ2fbKRPyhdZyVVBTfBt2Zxi1yNMbBLPwKC69g75z2VRQKyGy7f5xj27J3GO
zrxrNFncoKdfdY06pggOKV0gargLotjELUTKnIxrTGjLWqYO1cwoJ3/jCN327kdo
qvjv2MQHmQmysjNBqyG6XiuacbBvE4S689JYFiGiyC7T0SI0kPVNqmqYb8uG4ZU4
tQfUM57jU61aEkBIvdoVGjAxGbcHLYCpx7/kQ760YqtWUESpxJUKGg4Ai4LkyG3q
FABejS3BZLDJwqd+WzXGyTAH80S7ezhVE8Wt7vlS8w0265VZhIF/c9dZQFpeDog5
dcihao52RV8x3z4fz96mGeBGK0Jekx1WFLysdz5WHA74G8eNAAthBGIwAkLaKBdk
1MKsNPG5kxJfNzN3VG3YybnVfKpevcDZ7zrG3Ix2lIpYTR0JyFIqFFrp0pdyYT41
fN6zbo9thNvtizmEQYQIPf+PSy5Yx5i6CaUumu+W3f6Ac5TGIuqfsYu7qUuloEIb
8jM6ntb5JgqeMWyF3VIY6pV9IwtiljB2mMlVkH8h3AqktTjaBkef3ltkgnj9u84a
fw398dy6SawLSZ+K1uTBXOObwkCsVRyX4jaowPnOEj5jn3P8Foz69ospkaq4DAp1
`protect END_PROTECTED
