`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOYmAY4QlIXekgdc4/HbzPiurxY5j4fbReAC9nMeBVFuzs7DMH748cLEWgTPRmMV
MPaX6PlCW8vIupAkrfrrn4XIXtOFeeXIDzIAzQwM4Tr4DixWEZ4uuG4c5omI0X7l
lniS76Upzi8V7YuLoH8vZ4C/V2YH++zhZWvJ4+/bCbwXiy0EghKKQWS8J+Cd2g6n
oYEsbl3ERPEede+1GDAhrpfNehn5kk3PQ3H/auAqIHz+z2nYDwdpN1IoR3TCRodC
mfXw6ow88TGTqtYxxUMk2VZDcBnN9HvCOcZBkaUzcOmFmbYcsYq00RWkUn+HmKCJ
tdrPJT+sw5b00oicfNVmV3w0jEQbrCUmZBmWO4rsTlFKEC2Wb/tpEuVyL2J84yr8
MXmAHbrAUQbhoVYHrUCTIoR0r5Q5PiUrLw8hniIREk7eJAOfW13C9mV4TOT7Fq3S
J1KWzXVfEuKMb90rFIxRi+w5KpgXiF//h+LYafbr9331Dt50tDBRYFpZjQjYj9kf
tI1ZhdByy+/E9FUwV0tiAUxLCPjmBP3BAY/KbHFzK1ZoyYKI3u1LHO2AvEEvNT68
hFkFQrxN7Fs//1dHeW5NbgG0lu9H0i3mZsMIsGm683VErSPlWbNDl0BdjZv9a+A5
O1Qz2L6QjSsC2XDQprgrAEQosiRw8Yl12aH37GfMpeBDBllTk4SXlkeE+HIEsl0j
LFhQhbh92oezr1MPavizXMR4mpH4jzUC4D7uKFBY4dlSfQRFUuxzqqwAcjkCixIO
DU/7qnB18yaLjUuB9rSeWY3nMy5dcRptWu6VdRtk9j/dP2hRWsnLFAtuKY6MMUTz
XCBVS1AKtytIJoaZojMyvp3jcPM389Wh7Z7UukvV+Ur6RYW6G1oBbeh7LOTzy/Sw
ryI3eG10+/DqC0BhMzNjGsh8iIsI4zxe/aRG7JvDMADQH+TUrlp3C2Wf/a+8Fqs9
qCTZVtBEVgpS0QSnkInRbdeSCGuFLV3DmEQSZRuPgq6Euvmm28FK55fXxqV5I7Uo
GmTD9DgdGyV/8TXSgSKYN34uf6Dkrtm10eJAhad3hXK/2NL3QqaZhpzADLXWMEn5
4jpo0+aHnhcTijmrL5qhQH9/8zetgyVzGHrNwV2pp3gFsYCnTjQwXL2Z0P/L5OWL
`protect END_PROTECTED
