`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rbBNuHkfQaGcaGNszniqMOBRaIs8uZ0QXyc/idSA9zuNSgmnXfz02lsLafZxgYpe
jmjX719X27ognW4Fie2gs3M81QfBnzjRVKeiYn1gkvS/6/YKfDSRT3zSUJKWOlVG
Ld4t97BxXmohFj66mErNROQxTSXqD6ieFtUU2hQ1rnyksvN7JeDd3G1e/aWBL3D+
wG/9gK146MlluWOAuqKstbTENWHcim0ub4gMxiYtJgpQ5mVVZe0PKyOQPi8X/v+R
flJYDr9actSWHUhe1/h/BbZ0v/xLjZs4YPJ7+K9UaeSGqWu1V+NVkgsYMdWGuoWY
z+guMyH9nVAXEE0zkCH3VNcmwxvb/nH/hGtrg+Ng2j8o0jfe62EMMzOLWqwZtqZ3
oWWcUlCHhvF3NaqVtzXrm4NbZs8NbEeyCjCh6Ahyx8f8dcCBGkMyyR+gJRYZaf6b
NR5Y/qTlRLFYdibaGN/imZjpN1PmLMl6ztT59TerUEDF2LRNjcz4SVtZHS2XqfUp
gQ4YkAebGIW+SmD7O0ogyvdTDNLaUlPTLBizufFb427zsFCeX4aMFfkjYbnwFGtK
v+mZgMXG9G5Cu8TSdqmcPS2u25JGwEcB3aWOoJnpCLVxzTb1/9HeqzhZKS+3Sl2h
Wfa9uKTUhs+g0CePBAexJF6OussqI3BJZgCrXOEtIg5rxx8e9wZn6+Vf/6OyMoAp
utFKTehLxvby6kWt9VSUjE8L7bUDjiubjbgylGZtDm1Ias4pPt8ooes8M+s2qukw
sR+ybQ5CEKrg5r4EjeDrTbZdCfj3GpuZH0CmBDzOdL3YtD73KmcpAqZtRToF3Fw8
unWn9dcWtfDncoRwy7LcnR5D97DWiIH4IYRUbXrzBRxYujdHRN5reHJZhbUd5KK8
miwB+PfgXehWNlVvsmAdWsNZLSW5vrvty8cwuSkN5dZ88wxdXKyMUvUlhsrXz/vL
wDqCsqqiaruozhsXalC1uvb4VT+tEzrAArD172SYH2B2sXmUcoC5C3PHw6wMwRNV
FehosOcOuJHrXouSfKRBAQYd8RS27f2qYsqws66S+nodOaMhXZmJmrZ2COt1PVhH
ZWa1MyfN08Px37UBWnrfLGQp0EUo3+qgYg61sfr363s/bEl2fsE/USj8sNU4P6wq
WgH/TzhKqFwwDIscShNr11Bsf4/BsXKi/VPGfbskGoa9mimWto5M0alGP6HG388y
ZEBPGS4nTonuBnJxhscn28tki9BoVItBS76sTjKJE6Cd1mQ9/dYVPZx5Z7s8TDoD
qevckGxjztyV5uIuojCNYA06iQknUrveBziqHj5nVfOIqr9MbCeg63rlBmZsnP2V
JgmNFht00r+o0XJdML+ycXnWbL8WLjFrnaormFeftV/M0SCLgYsZnkrmVcvn/S85
1Gkksq466lj78eIZWFHvKpG4HUD6IzQbFEBv2mhT8HCDCKE4nGIYIfDefiJlnVe3
pchQszwWwOYXq8tIdtdnUM/c8Hxfdkm+T38KP8UKma2fCErVj8EGtvMN6oexQISy
t+hFrUd5TURuIgKoA60jvNojVKW6yIYVexPiu8q4kVlXz3AJE/fm7/lpdfukkNHI
OG7USRmy1r1zLCdgSrHP7PHpGIffYR71IujPXoD42+21/E9wPWSA61uBI46CjXQp
l//9FaPUiW07+qRbdklBjKPJJLIOuhkH6td9Dm9dI1J2Kg4R3w8QnDXED3PIJ7kY
RilV9Wq8V6PNE0309NIct3n6tersn2dFTBD+SsgpnGvy+nEhghIPdWMlXcfIrVl/
hjKu9IhqLOmNuny0Q7F2lW6iVlNS0KPLhOOzgtYma5Zp8lZDOBqcZaAUWuwn2mMc
JrySiFXNembjeZgA6LxAE2z4G4GvGX2VomW++GQfd8xbMhr3kzGO75FjTGxSA0KB
XLgcetqw1+CLbX43y6pHI94mpyi/1bCn8k+K1nFd+L1ArRqA1YXJrNFylJH7Fh7C
QUaDKahzXN1ZzFs53Rf1XDsrrIT3TZxt48X590QrvUGUj9TBg1BCkR7epaxJK6Xu
PiaPd/Eq/Ezw5ngWN1iFEsanhcfBf2/n/X34/m5bGKmoye4WAWepBirjalP0i7yC
BxVcSNafB+xNmc66DXUcZOkoHhk5Z40o0IxCLadL59rIhW3NBNyxlH8Vz9jgbGPc
yqBIVHGihvWAKQXBYSGpsmUOTLTD5W2S3j5M/8bPQGOJpDCFY/KzgLN+XY74s0Or
U0oofwoRuVLVqoUYvq/ZX6k48jO8auxxpOH2mVMZenNMsYdtRSPPl5V9gd49m1t+
kaQ3GtO25AnL7Wr0SKS/wiafGtBc9IcV/GmC7FwCUZlSWdv9zdtNZWRjVzewA85J
ZtQL/ZrJRr2ah3ursVnjn/v4QvPtg+9B6k7ICNHDJiCBvBMQJEabGkjI7RZAqEFl
VV6Po/tZmTvP1e6BEKlIocyr68igG35CuhSUc6H8LsdZYMwfRExsbEVgzHUGzUa2
56AuLJlt6Jx5RD8tURkiY3+tE8+uYIkB095szBvolXNFPulmVwsBj1RI2eRJiXJp
9fRFG9hOfrdBe3KMGhBii08WPdkzSRlN43bkX485kPJ9way1CSB98QEFtI3cobkq
bg6ygZT+tObWjKelVOOsfovbmXBLllBAEsAtvGWYf3EOkBk1iPBaNBB58sONIRbg
IOs0JOfdAe5yWRuVACbE/T4KviVGS321kAx6ma1UqXJPN7GvzsK0yGV85WvzF27D
QgppMtavMwDEyJjoHjf/xtn65FE2gSIG7NQUBz0vMk5fPXQMpWP+3IjANnDLIPKI
Ni96NyBOGdFVfGCVOXHjaZYP8ykv6lG/WzXWeVCLrRwZ6jBRYwpuFbnsRLA6e+A7
g/+UgwCaNsIACTpQtHxWNUBizJ+O1NI5vUrkymBdiT3n/OQRF6gRxRQno++MYJ7v
6gAdQgUrQqKg7K60dI/4Ivn86j7H2AgRx6wY+0VyJaPqyGdPSnuo1SLudEIa5Gjy
/Qc2+ztko5OE2sp9vQQ/eQVY3YX/49d1WdURIXZfoEH7030R1qd0MN5YnVteqqyq
tIt7Ks4MWSPM4xBsRhmiieGYUEikiTiKRgeWRVgNQXSOzszzMiwVeSJTVYROzb80
/znGqwym8OvPtBe/mwpIjkxFfF/lBBnnd6ekVzJmJjFkvcvuvilmTRAUFMOwVBdQ
C+yGX85gM9ASuG4cUENKoRJm8qBEhXvm8Z818AfJQPBn5zt0p1VjXU1f+ojCixWY
pvFpgZbQdq2uQ8kMSwWBGKIzSZmSwZxYg9oI277h69hhfrU1RiZ2ybtwR/SYbMOK
40WkHF5Oq0lNk8bLjdtk83aJ5Jg+onchwqs3XZrJMqEi410Ls9OT5S4r210YuXqK
W+oikCEOWBrnAvd29vtnpuh8+VNarkpu4eVnXn+ASIb5xxKdnKCG19pFK862TgWZ
ESp4cr3wgNgZFTe5UF8Aj2wGJk90blii7hf57/5vyoYqPos+9S+jDJlPmYvUYK30
3KW/17fFC+WGURO9nfl7po+sbV7l6cl+VVrkzDx5hYjnX7yjvL1uUzf27FUJGLkv
nciCo91dAzDm7sKyRs1A7rrgBWEjxdY07MohNmDYILih0YOzXKifXq1ggJuw/pb1
fuAggEHxHd6+IFjRUFGdICU0/sIQi6AQa5NMwMKI/JeUd7qPBWetrWlydU6jHmOh
/qLbWLuuBpBOk66rOx0LRtY9dIYWlg0acvUBU5C2jAOS5eoKYP3DpMkiAnKTCgVR
K/tNXBMVxwFd60mEz6F+NoKaJep9KrxBlA3UEqnhY5rrtz3lwy8FAvgT59FIfjRW
jAvBvtyKm794Y+PR9H6Li5u6SNouZUu43b0WasjIZ/XTCQElwftFQXXmnlUgLFxA
lNoJS96FPlJvV64jCZz8oRzkBDiuoP0i6B4eBX0Ti9MJPTP3zotzWP9IcHPp25s6
4tEBU7W86SF5N3IEKkdUsJvGYg29sRgVvysrarkWrfcQyHT+i9guGpUSBQue3pwC
okhy8rP72XiDgMq8VQ7BUa4V1T1AxKy9ddxYKMJwMYfMnM34K7LbIvkXzNq4FPwN
6SxXQSpkcAtXdWNRwiO1mClnNKj+wO5eHIWS+2DS96EMkkg3Nxe8/OZpKkOCZPTY
oYgTS2RNxfvHRTUewzzcSj/KY6qIohlGj5ro4Jl9SiqTKXmDSzRCA+QHE1RpkPrE
4VMtscOvrz1CGSuTW4/7Y0Q5BgflBUnFlTi5+NXcAWVHe2vPeeu6hUaX0u5JTM88
E7s/cRE5z4TaXqCXmeim1bLo74vrRmgSGopj4HU5ZDiMd4ZtFhwXCMrviYIxPvmT
HV9MpwFatb0d/pXHz8y1RJgWjbe7hz45MKwZbvd1qOsW38gb9vuWhK5ANewghqTm
ixVTZpOatx9jBFKIPg7qOyCVU1q/SdoXDJ5d0syxejbpkOIVjeNfkCv8ClPF8rPl
yMqb9NiaRGTqyG3aPvnIlMfBcXW4UojDQxbg11suCUDqXs7LdUTt6KknUFKxOxuc
a5q2b1OhnKm/i/uOZJMd4oXphJNxa5qT8nWLNKby7ducOMSJnK+NmE2zUmdx26so
vBwjPRwI5yKoMMEuo6pTawywhDmi4xsXJAQg7J7PAgjHhjBL4WNbIeuFd7fSfVI/
WZ/LQng/igB/QsCwXYkVcv1DpYTGTTeW6kF2O43uJpDzicNkFZTLK9099Pb4rY0k
ByBYfk+zO7uIhhOyULVA6gWxD5r/Yb3Qq1RkWG97/Up2R1QH82ZthSxr++kDNnAe
+7sJovLq3eRXFdPT+ebowbaRddjZiKmoBEwPX6g1q4Fdxvo4pTLTBzD0AXHtT9vJ
RVMED3acrg+QIzbsyVxl7Epx8KfOfSHoGsHeJOFokepHuKm3cIDCjeDZLRf4RII7
On8xsVcx8jR6togzFgh+mvDAg/7LunfHsGdRYLBfY8Af52fTA9w+ojZrA9pK05lO
x3aTWaulZJkMZWZe1pzm3DWvzjRYo5rCRx0Axmx1dxUZhYQNxVSIjjOX5b3FYsCE
OfrYI6BnirnRLq78byAeImMEgq77KhfAOzqpL0gZ6pnonPpyt/VzgSD2kLYvviwq
k8akS8Za4XnhgN+iyb3Ckq2bRj6Hi3q77wDYMmBXM6YSHDSjviRitHqCkliiPmlg
kLcZ2uOerj8aHcK4fhO7/8yrGzazdIqbogW+71mHBcjYCxPURq7t8GrXjm05CAUI
V8c9dGmOJMKrjvdopdSwX7/E1ghjtVjIsGKEEa+uB4bbjn8H/FHZrSam1oxDNA6g
otNEerc9sNu3NVTvJSpvNRvFYK892nwhUXiMBFzh54VC6N6YGtwPxop0WLLZ0p0F
Eenp8XfPEcmboj2KymoUtkGBwhNNNOQOos/WCqkyY3lRH9yZNzeDDi8VxNqZV+Ya
xH1+WMhNu2t2onwhYTPkiztsfYyPjSpm3NZhg38nAg/Sj720i0eOGxsJHW0fqh93
LOldlVtVsupF1UIaXdGdbKFOt4w4XTjtUqKan0lJyonNceIPrz+ElUUBF165SMV6
kkTGJSuYdMP81y3nnoLjKgRPd/hKMf7ME2mf59lVjmAAB6mxj7K30+lgcKtyFnLq
NWpxg+1zRyCZqkWm9KCeCh6qJaxojPjq1KkiL42BF1+SFz8dKgwxmP7OVdFIuLKE
R5YY2JBmbmlu+mLFlLmZHw9Ufsc4G7hs5vl8gR5yAc0kLfCqqPrTjmq9q6uoQRl1
8Hlps0eLRZnKQEO4PZujMrp1PIUqENgOPODNhd1QUqcJgT9qRLr1UbJlAToZkBfa
6vvl8R5p6TMcEye5Yd5L3Q==
`protect END_PROTECTED
