`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Gj/GsL/jEwP+/g1WoIIrao6vPj12vIhpKDRSXrqvNZOpolcf07GyCxBTU/UvHv+
/IaCn7sUce1Wb+wmA5JMlWY0mDnAKnt93PZJtwWSXlROTYUnlsx5mFrH6JaGZgwl
5HxLU3Sq1NPaqTRm/B1HnLHpvfNeNJiDU6wT1RG1ynw0gaVc43dTFoTnJktZVroU
KrXjenisxJo47k9NPLyo1Xh6YzU/sxQ1vHZ9R3cLuX/jcg3QQumSnLM41e/KIK7C
hv8G1SsDokfoVPsTJG/xecqSQapSsCVDjnqPiSHLhrvXmMhZdrKn5P4Yre0gX+jl
V6GDT0xCpmUCfifAEkbSQmaVApwtCH03uxVqObBI7lLThO3C57UONGt1CG/W6l0v
CZamdpDCyIyFp62A+VK42sqNyARAQIMbzdRy9guPL+xeGQ0SbdoKtFsfJPtcgl2W
EiFwqjt3djVPYuY8G7NvI5QSsp85sQB0Au2FJ/Q8nTTEKJYl9VW0KnBTVXnApW7p
WPhGGgPivFvYLfWNGTFwxIw4uiDGYx5tSCocXzHw7KEZkRPTRDWHnYNc+ym+NwvR
DBxcxyzmAzW8YYQCxTdHfuhjTQQjjWuMNJ60mNRtuxjRO6WkkCocvSn8cV45GWVR
9fHytTSaTbG52i8FCwSqH6ztkYdM3RI372o3FHH7Gix0sttyBwNqrKAN4PzNmIwe
B6I6OZBA+BjBLmn4trgK+r049e5IAQftZsX3VbArJCv/GjffBntJuYfJ1g7GbzB2
D9+zMxv6mAH/sYuwZbOE+rXT+eVdeAvtxKCGGjPknyh6ZB4tVPXDOzaigUZmygxK
zP693qWjRDjYGAQtD4PFJAqzO8Kx3NWv+RiIKL/XS/5ickh4AzjAI0zDtx8Fiu2p
SmIAnYU511djw6/WZ1nSG1lkhxIWHJal2ImqC7zT12NGSZYbFHWlvnWSTld8sGon
F/h7Zbb5Rj3EjHjhyqz7MrrLp6oR9Wiojdw+8wL7xvWh8IDhcGCLw82Ya5J0Bp8+
JfLHQ6myXsn5ikShonCMWlOaTKwXqSH/KI5MchjqCHDuSXffqzXm1CofUwpKEUXw
VSrhMtUxyqTYNYgQCVEEH+UD30hVaEJSEgJDfKqyYq17CzJOtdgg/CJRMR8GjHHN
RCHCe4DhFOM26+8Vdzm10Q==
`protect END_PROTECTED
