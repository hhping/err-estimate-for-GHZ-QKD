`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BM7oyTNbdk5wxxRldTOXINLf9dL2ywEAOl4n/CjBX4C8TFoyZJSM6UWGQcl7kDpE
A3fu/oe/LRloXxSgyWrVx5uSYh30FlCZfIlt7yPzs/9XZHa2ijKf5BaFI8NiVmM8
CrU3+sQVpJSkog8nB0KR0/Zm2ezUDgSLkHlf3QUeRCnvP+lGNcNeT5fv8PyqF06a
eNbTw11cCNyRLAH+pal6xJdTXKnbOWCSCehbGSJbm4CRN247n00uVJ0HmQGZSS0q
BH5GPtDKWrKSd8pyyUvIGiC18N0ocihYjQTkn6OJnQRlkVVzONuavfqmNd7/xkxG
tHaGe14PbQMar4yY5qFRCWvJR5vq9C+HxCPRW05qcaBhqFlAFFl+PKi8oSRh61BP
qIB+ujjVaadubAF49sTbTjr/LEA2c/WXkpLAXlU6+N03Iu8SE5IvfymNggU2mrvS
VDnZ8cYWh1jdHIB5uMqSO6KGyd1QIBTHr7mli52C/PQ7HNV/bQ/RusJytLEUJvmF
2oouHrM0QZnl2CPRCMW3y4V2N7kfRT1ebAlSaxtYSCxWugNRmK3HCV3sF16qhVS/
vPQkRb5s1WiVIVewEN8RGMkHWv+FXq0/OBI5wL7Viv8cWr4JApMa8gDvt7x7Gf+Y
yfM8TtaA9gtmJgRqJ+7M8prRua9FtA/3BCfmSr1b/KpkwFZPeDO523FrN895Djef
fR67hEZAA15DZnzkBzIhgUmNqOumwTBgkhljMmdbVc9Y+Re3l2n7MsYFFybA/uBS
dOZVzR1/Adcm/zlc9kePKg6gtvSw9b+tZMB1OpXodHTq7qOY+C6xsnlkYPsLbZTf
T/r9OPSf7O8JxRLt/amY8ArN5acOVBrilsDfwctHwCrtFsft2eMA08bfYxGFOj76
`protect END_PROTECTED
