`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFiPhqOJ0VN7ZU2ags22NGJ56NPbAN/7rWfWndo7YGQPNVC2/44srFk07xVBdgzj
cuixUvw8bE5htiO9xGo/b7BR53AzgxiyKu35TYkbbmYFscuiMqAYBfws5O8jADh3
qeQ5QCM1Yy0WTUSAwB1c8UlOh/mue+/AX4YhCKBTerrlq3mfkaGOwiS8KlNIMOpX
F1L+ZVTscTZmDgv5dOA+tAqowzq3a/yFGWDukdsU04Qd/3xwOtJowHVU0ICJRTuW
Rwy9SlWB0R4i/Adiiwi4jA5HHS7X22PcCWwkqIqYXVYijkSVD33YIFKL6MiAdPop
+8bZ4qRWIOX6w5zQ7iGq0ie3fghdB/9OyaKMbkJ952GL3G9u7hGvQl6yfULlKn4T
QLSY1T+CFsJNiwIn2dOCtwFPZIUyjcg6fouE64pe+z+qHQfTHExtqr7IdjYauGQp
tB17vcwqJXOQFDIySkeqEqzeCtqEywKGEXJarjiuKjIHEMoxF5gDOQJ6J9JkpFF5
pvE6b9ZbUo8mOSa1AuLz02qdCkURg307v5jB9MJqMIeIOtj8biYgerbH0WT6qjoy
0burFbmcs3HbHlecQenJtTVmVIkqHIZkI8uQl5nlefVa4ZjHleWy0og7Xhpji1yb
xckv+cYSjR3XTc0cUByvcgCwqxvs9/KK7kAG46j7TI6bVH5z9AImxsALO1zcd/Kx
DRHip4Gg2xstim6KDbhf/gemz/OZtz2obNFeIjoAwHb9Ew+LLgCAtFTsUzULbx/M
YhIz/1XIVTmwRzA8zKuxzDLw2XGQA+UCbNNVCR3Pvqof8xL+u0LSC8g4NyJ65eB8
EdxJK4ROIQ4nFjC05gTAGNYtz9yenTbltAvWOOESzKe220NMH/dWb+s8Y9QsEoga
8TcG1xdiTTp3Ar6/u9/Qxjz/EFWYFrF0EVC/P5ivaoY9slTgtZ0FHZZDAcMvm108
71vN7VYhiwG1EkORGaPx+oiFiwJdNWMEjXEPogdNzKeNf1MJS6/pHmuYuYHdTiuT
rjSn5D4W9i1IwllDue+FKkP4M28dsD1hr8KyTTBj4dCEIlEWxFAIoLYRbv26oCgV
34MRoNC+VF97/aREAtsYhKW5jrQVxc8oD/nKf55sN5cojEMXy2qy0psdDU3vf0ht
ICBP0a8qU5u0UxZ4+NPDdVSQszREPqb/Pj6MRE9mJCsdwujF3MsqtwIKJVPGg021
EwuSy6bhxHHA0IC2sn6Ok33etGwPOlwH6NDQHJxeIUeFYibTDa377EZ2G3/YN4H8
Gdnyq7iih/xt3fupJYzqlrrAAom1vYAsdM4ZsdkJdVowO2axWGXPzuhYSNxzWu/W
Ww9byd8H+Y9iAHQsHtjJFiLKDrQf95YeAiLKNToVtg00METJ5G2SDR9axc13a1yI
Y5cwDfAOpN6QU/jyOUsbvyyOKDDMUhREylTR0idD+iKikYmOXUaeds6998hrfUYS
c1lt5L3DIeR56GRNo8D5QaLNy6PaHZK83ieExgoAvw8nslJsGWynatfyXvXHMOcV
AsBLDl1zWpp0tuBJdql3QRMzkD/F78PItSAG0z3V51NjSdmw/mYY7eLhFjvVrAJZ
LU2pMRDqRtGRLv+1GEhBC6olfFSyVhNB0FcPMfe3bmMpj+Hhd9LyZVl782ZF7wgX
fcuD9fBxKZfn/slAkoDVxDVGKvYNUSpmxxKoI/AH4Xp4GDe2E0hsLVJyYwAqbePy
BKk3h1av81ixMPVRNvjNk9howqW8JDSBoIoX2Fu/czS/Pw59SJcu8h7P/lz5HE5D
tF4EgaCqtSegOiULKrQDGYOEBikBomfVaK5ZI67TJu8BKSHwdoem15AmVrgDFTFN
RgGMkppObIxKB9pbRjx6GpEEXH1sfSl3hAAGnOgmviKKLuDstmS95cO+WHK+C6R2
fVnUk0eRbZidQF0exOJcSraR8RWQXikZa28F1mPj0l/vE/pgcHhUc/SY58abAQlM
15x5oRqYfazGadBvqDP2WRETnLAAWu0JxHJVy8OChxnDYjHGwoKpcWw0bPJ5yMpU
TtTspXMUmPjOtBFQ0Z+Gj6Vma22uXUs0CEmBui37KErivhXImjWAFSr3gZO7d8Ks
u2YEP4Cajuw0sry3pVK3stGGyY35McoyKjQrq+cwpH+ql6F84OWxFua95JL+0CWR
2jHFevndbVXWpHVMNdfE3itTUYn+RZNSSlMbNctA/oxCcSPeSbLxbMi1vp60KRlF
bVA0HuOlxBO5Yxac04ElP/bEX1DTahPDRwpkJDf6cYf+zCrbK3RrUa+ffSTFlmxp
2kpvCw0+huhzbQjfxNJJAk6/fd5F4bvrb5A/Lcy/KWyzGAFH3LuemXZptzpFfA/f
mDF39u+1ijrumLu6GEumKCyGEgfgAPlWT9HFLK02p+OWjU2GDi5+xgQH1hdvS3b4
xSZlx3sEIJt3grcTZEN7yRwVfvz8Qk/9QMniZl5XXqq/0i5G8PSxrgZ0EQmfdyRx
ZwB0NEpHLGSqNQyM6GM8Q64L+w42lMSka4kBGpdUH9I5BtDPKiF4V21k1xiQj/E0
nkEWi6jLg167V71wJGAlZMkctNM2/LyemPRM9+qqK0rF6VoqLpY/apP+z1kq15ip
GuMtchPzmm7nf/CXvHq6hBEI737WXm7wjt8+b12kIO5zcF3ENfBoKK6GeYZZSWAF
H23pcq7XfwpNrPy36IAfTYEXmGrpVHPi1xdYaoYPbetu3quUpWXD1rHExZjlgMlA
GmW27Z0wIOhJsA/qUAIGRLqVN1+x20SHyBJ9KCjm8A/69QrfCzIwk74++oZRrlAe
ax+q9eZaP1KM1s2vqsh6ds5HGMAKwYjTb16YnM6XSNjUc0AgRxRFQguj3mkdpBqX
1Ge4e3psVw/Jl1SXpdHv/lXepwC/S9Wn9dRHdILHGbkOtjET17jX+3Btgu80XWBB
+VnmoKyxrPLPwSAs61BCNQihU+dZXttAGlBbkS/HtYUJ1xybvQJ1MHNfhrXtlTqp
Z/Z+xBtOj+gWu1OUhLLCwxpt8hNFyURpQ++FcsytJ9pdOuSTRS/15e2+JgNWzDkA
JztHIi/+FLOg3qb44AFU+Tm5w4/3BQGjUeFMw/GjiXIF0aAucFI73ZaoCwmR2FKy
yMAVmI2PI8d/i/re0QEMFD+hg8nAmBquxbgiTlocwhlMmvrrTshMlikyoqrO30/A
shWHU7u7vi8WZsT+yJEhIFii4PmELTzA0m3P73/InKdq5cL6JbQmHXTCPbFP1Ddd
YpsI4QLXd6AkYHeOmz7J38u7CuitYCLLCNePAMfCUd7UIYSRz5j+hqHKTVJHsb0Y
S5KFLmW7ItUF8Nrkqxr6RtgB8qYMptI+fuJQP3p3ELhpOMpY42J6qyu50V8FoByd
TPGNVrQtS1DaRnl12IkwJu0mnehyLpnlmKTS6otm6/n+DMP1nardeJHe5lWqFIBq
2A3hXtB8ni+TketkESIIYTSuzCu/VQydcQDElbx1s7aot8nPcRAstfZ2tApvmUDr
cO2HEyMVArVBMbaTVGUtFakBDUs9RwC9ZsUCZjVOw2Vl4A8BA1D2c/3uzv34MLbE
MmK3daNDhOnqJ1nkXMS2604TN5C0sUUiKUMDKUF9XFacb89kOZdMJkEmobJTts3I
U1IuTq/nVpMSyCaDO1mN0EA7yiiWdTUufBOl2s4RXFRUTtLZUXsk3Fa8mtI9KXZ4
/DF4O9hBWS5SaAf0xW52C8eZQ4PdZ3sHAgqLHjG7583bAoliiy+HfuOfooEwoFCI
MXkbMuiYhCfxqtfgd7+FOHWD4FGKBYJYyRmsvJXv9SU5ewBpSOPyKHY9PpdisQrT
9H2h2iVaGh++1jPR/7SHBCenqpjR8SKih/gBxSlo9oTeIh9mFhbpED7Oo/B3v6sz
NTlHnnCHpfezjT7WFF2JuuGSY/QQ3WdAY7IVOxlKbQwRzmQDqVfchM+aV+xhoqMw
QsgId5UV9i4UHRlsVv+91leyFPNHFeTsuU3XgJTtGy2f02mc73UTPzwYPPNQYgEu
x6l9raH3IrKiq4JXM3G56HrbeB9hHeVK0O2CWjsv3qcFPqT5bDgLFiu78AHrGLc4
OZM/QZmcAKb9XGZme8kDtL0yYnhb1Zk/BRY5IFtQgxaVTvX55azkXN0hEDdulhNi
H7iXj8dR83BVZkEFK94PKSEJiX6Si22Gsgk6xwkUS5sp6/uQ5a+v5h4xtNeWEGj7
7jt7/cmbF12cRSZbQmGg5q13HkYL4A6c8+5YD2DoWDx79rr8YqpCc8tu0eV9syKt
OE0jJ6cmhTFxB7LohrhMBW5iQuktR+UEXzsXv+aVjXJk+PE737DhXpAJxpPXau+n
`protect END_PROTECTED
