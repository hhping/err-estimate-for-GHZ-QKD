`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUbXAohkMpYz9A4qLf3gGmrdWOVAeIcF4gVKRoxrNHwcPw2tFzSa/PeA00+65qM+
E22ZhDKeu3a5uRHECdQS2g9JaKTJru1rvkSwwXFpR2iddUcZoakniccgOvFZzq1B
miulL6FvWTc40tLnU1rNpK5A8FYGzFNJstOUpLuHYq5w5IwQgZjwuROmSSxaHhRW
MLetrQZ2aM5/BEg8JySkXQYOcl5IIuJ7Q383D+W2GCYf7Ogxv5g5sUzQKHXXHGjF
/T4mcGw7gk1ASfNV7RESMPqy8df5mB8crhCWm++in4gwOEYmgxk2/xWKLi3IU6SW
kIrMoB7Eg6K75Z9RF2WWNiI0ZlIwfP3f2RsuehlG1wT/5zgcUAUYcFcOWLEQvsBm
tvQZXKxdEt9yYe362V/5lwd288fSBEEuusvH01RCihDQhlwg9MGb0TnRGzJByMwA
MhxcaF/gzu5ONGPX66/Hd+RKnMLaqGwjjdGCo9DHfd0HgO74rx24xPKFmq3jtfoP
AmryAPb3YLnE3dNuXw2yo85iBjMG5+2qYmWdlUfzYkClaEHFZ+3hQX8OWbhF37rW
ZPCBofkPixALGUMRVuB2TB3FkLnOIKhSM6aOCXFbLtOtYnNlRksNZu3NcgpVyFYs
MX/sC6IlRErZhrD0Hjz3f5q3FnIiS7h2CTssWGzjmNb2S/bmm85XRIffcf/4VSHH
XX46y6670doGH4WkEPGk9gFm2NcPVJ7x4FJtKZyw1bkMn0cjuYDGavC9YPMeiPHa
D46E3nNzXqJMa83dxK7GQSn2m/AfpC8S8z7X7P1fuXlv/Erz8QVqtxQxheDg0nNl
jLko/laPDcCXkeXNAwSmsU32PVZC7uNje+TyqSFBNUUCLpe4qI9HVX7ZUFLntoxS
ragIOh/QUuZDnDs0YOhc7uxIpibOYa+5FHAbpxUuznW3r9DU8aZwMwdTLgHk89cO
GoV9Q94zi7P0XgdE8e/u36UwD30BOOAJU/moW5V477AGWEuu+uO7eTjDBgsuAtrC
gPhk8oDKzq+oy6dJuPdkJNnRUvLuzeuv3uQQfJyDT/i7plZsHdhgwWexKRIi14Ik
oNluQCyFwwfktv7jWOQu/ylTDxcluIlNMzZ9xfnf5/RIgqudtIxl8Wd/dsiZko6c
rEeAk6yXk7Ly4ePnnEJnX/gCjxmoru6AAhj/JW1GtNY6GjoxxZPEIiikF1hhIwrN
oNrsiqHQCXE1AOw+ClWdtleJiGjERqLUwzHPvuhasmLOtbval0EIW5J82ACQ/5hq
a9vfhPEkJC0k5f+Ii7ZjCOERNTnGeL9RihArFkFrtsPSiFsmHANfBSnINBi9qzfv
T+mvGkhRyygCoffE+R4E8dB5aceIL95jJkmWeM0jtBuFoI/6YyMXk2xPkso2t+jD
fJet97agjdSm5YT410LzL58+Lsj0UNKhi2ph/mrGpyMNlT86QgddB9CiRXyEvKU0
Y2WHwjLVPiL6q2Qti3/PyVk4tG7Bi3TqnZIHesAc0rc=
`protect END_PROTECTED
