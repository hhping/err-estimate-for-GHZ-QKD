`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bm0ZMQEFvz8sA8SJzo1ofStfCS7auIjwvqWxNwtP6BPR6alIxBG4NVcPSWqvkKxJ
vB9oikXBlCb1/Dj2hdfaQeQdRH5c/7x/7qrFGO4XSPX8CEgeErR4xUqnDiuEd9Cb
vMNiW2qEtiCCXxkRoepMZS/f+HvoVhp60wVnEC/rr6ugkVOcOedRg8c+EmRRjHLK
GEvKX7TqhcA01DxTFNKFlifXxN0gnSdekBfc1Q3uOvEVvKGu99utG98xWtidhyTM
/1TtpPpsTWb+srMTJ4TOEYWp2vAnB35MMrPRce6cHywwUbgyqy/wLEo0AukyTnDU
DkaVTes4fBgQ6BrgI54DGokaj5SdmSzlAt86fYq1hbgXZnX57qTNkiCF1yP+CTG7
zg/AbXjinu+xPXUewsTu9xe/J7dOIay3Xf7EzVVvrJe9Y6ZLbXf47+GnW27I9JDZ
8pgGLBI9KY9tzywH3mgk9To4asu/KC6+4rUb5mv9kzsJG31mZ6MqlpCaLgOb0m2j
KdhiRbhvMYXbQr4eXFNqz6P146pCUH4cB5h7V8zxLp1zv9E2WgYJj0LHSx1vsw22
Lttwk56/90bMB6mixI45SWeBmrAEZ0vlxYjp5jzXmasUgV8vjbV0Kj+z+Kl24QlV
9ohnFGpHvISArLJbWbgHemcQlFYH3y3i+ohRKRpHCr1QBUS4yrQSI5SAaC/4rUMd
tCZJMnwfucBQgvN5tuCi/vCvka5yF6gAKLu2E/+TdQn5vS9ORu6ozzS66IeaxZf1
fd4HPFDlj0wn9cE/1vZYzcRpApOMHCn9tL7fbyGdm3Gu//PwgGvbhr7PdT7RwVSu
0Jrw7n+x89jnys8wSvZgDXd8aX1Hh/PS1pOaDLV3FIQS9I2L7WYOBta1xdjnS04s
mHeGGrQb2B06LryEsdtx4k1zHNqAvjQ0C+T4/k84Nft1fWO9FcNaHFh/dHPEmiiw
6LV+bxV1GcNeSaPcfhjJ+QgYJG+xmfITwmgVMFEcnb8whdtwJFxtU+S0KQUpd9BV
WNB/kOr4scpXUR6yjsD7dNTS3/rdj2BmuiP/SLyPl9RdMrhMAcV2yVrThfv2dnfx
WNtTwg/awhTOawDP7BZjKj/8L56M5zC3Okt5KHy+RzQxuPT9AwJigR0RJQNsqUzQ
xfASZBpNZ40kQgKluo9gJeUCvNaTwcRK6lEGt3GcSrgrquZoZgMBDuaj7n2X9Uo3
PpXOZyAA1mGWAHc4eSzmiAUVLxA+EVpa18tS3MdxTyE8CcStGH+IP3DGRKwsLLit
`protect END_PROTECTED
