`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cv/ex6FLigalG74Un2hRB1EBgR2eDKV9+DQ9GMwgcMjkIZ7J1RN2IhWXj+VhRar5
i3Z5gbpba8I2pDoD6wc4iKyataN3Y/bNeQ+TUGnvt74k9HHWdxtykfuSPbLiWfHa
/QDUf2hpekh/RVP58QDxUVVgmJBF5waETllBty7hWmP1VdJt5U7a+issVbQaU2N3
ZI1joN2bsBYE/siLIAmiQ23Dt3XIGcn66+QXkxfMmtGCfeXzm3PGEAK76V9Rgwyq
ytKO8/qehlrCjCaK81tYGAouvCIPAb3gBElvD8W8cX9u4ckTa8uX57jJQsoxz0nU
QGTJgwBCEjokUFOS7uVhs+0Wjz+EWgRfQpzEGqf/OE8UfveQLO6wthCADBSrZFKz
HlSJnjXi6TZHqARrga0d9G8+CwwGN3u06P+LUWS5z10tAgGEOC2vwvdSdguwJwoM
`protect END_PROTECTED
