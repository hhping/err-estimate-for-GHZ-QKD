`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YEuZ/4HdWwTO4vX6QsSOGBw3xJlwerxkIB3GshnIQPtnTx21LVCJoAjFQwpxTcO4
8tr13VgchAArE+WBsS5svGoxbFxZARlksZpRt0WUFpD65HX7QlaKiWfc4zjr9QTY
h0Rv+Xt6pxHwfJ9mkQonokAIPwUSTe0Z0VldsbeoGakr2hUFdQcxXKpUQyaTAVJH
JKosCmTnIjG4r9VNB7VvMk5BWNBCjmt6ChO/n0e7Li2T/xf7o6m94IXm1E3fOF+h
a4lIgXJ9IbbOGpQvVlcfO0FkJ5gqRFQAlE8HAtgTWZq6cJ3A3PLnD3WmJ6tPsuXE
ig69xWWwDRvhPZc0MDdEjICyV0O9EV3p4PjeXUhsl0Fk3cjnV7P8lmkCu/GryU5d
0J7dsqbEk4xw+Sex8TPBF7unrPgTN87I7QeYIRRxMVjlu0tMJY9SebSRyRVMgmc6
LqejVrZLXKHIn+KKRhiE6pM0uJ4mP5mnOuEiE8V6nK3aR8EI02hWmGduNQ/Q9DLl
mUonjiNjHmk+IQ1VGPrWxHLjj6SJgYoRxQOIsJGNYK9XF9DDruKJkHK/wQOnZcHy
XNeCmdXqkiKgImaabtD3py15kVahjj/6KRPyHG6FlZLAUTtlPgWj6NWzymli6Yek
qgYKQ05tOQrttuzAWoa5kMIfHETrPWNcQSVF3UqoyMZez10bgm9dZe48y6hIQjzv
84junCZWSZ2pnQmp+1VK85J8ew8ZVU8bHgYvQVndrmVprZmC1j9HcqgoSWlAjhoB
wu1SkoELFeKUG4ZrTjnGpFPTgMMm7rVunGUH0VER5hfhBzZjYuw1HlrZ/0CDPaUw
/6/N8+V4eJFiFNJyXGGmmHbX9IlQfC1mpob+501PJbikngy6YX/27oqO0K+vOtYH
hn65UGXFpxQW2PZ7zCGNV0gxjy7w5HKUsjDiTttZatEKlIYHq5PEi5+Syfcmc+R2
y9EUxhtv3ny2mfjP0gK3axFh2W3+dVXWjRn+GSVLDURkiT7H0T6NwijvFwsBK246
1KkUUEwrIFEfEgWE58a1DNabU6QlEBvF9VG9MT0DiQNjtVD2uqh4jmu9pQk7aYtE
kqXEHx+ejLr6SQFwsSx/WAyHRpjsM2X5UOMU+Fayh7B83Kvlv80h9R82gHeSnAHr
3FEVVXIOPMS66esnQIUQrx4DsI3Vn8h6dtc0xU7EW4hOFTGOdxnQpxneD+ZVamB2
JxLy5DTIWCE/Vwyw+dDYA/6ybwMoh3f9zixmIzNByhPrQJLBAlo3c98gX7PMc5xQ
RoR+FCHMjAYfAVsOS8DXoxWDNAfeJHguaD86EU/7M2U8WWQ6onUJ9Ps3Dyfy79I5
0+/QWV55ghtxLd4zZPnDa5XWhwAEcVqcGjkqV90sELqD68FPbiA7yUHrYigpJFOi
3fEv75Ckm4xQQhN/KXvKAmBTGoTLys38+udpfCJD5jKQFKrKt2keT9PnhiWv+Zy0
e+GZaYEp2WA9YlK3YfNWqd6A5S6+qtd/VUg8JxiH1AGQGc1p+2Na0cSzH3T0yK0p
dE267Sx0AiUKWStto0geG06Uswhwu82tMDgscw2qV8tm8hKWHDf60n7uJZV9f5ZJ
QHu7RRsycceYmwM7T8UA+xNvzgMZmkV2W2QarcA3e6Y=
`protect END_PROTECTED
