`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y9z+LaenPqMQwQX5dfgfx88JXUK9DAZRJfOuofMihNyzbPFW6zaADeBC2eC5N4e7
xcCVm3g5QiMxpZ7Ft5KxxTOSUCsZkJacU3w2XSlwtWpI8ONJQERo+Gw6P5TbtZM5
7u6kFE3KU3NHJuJlQOnXjVCERaS6xdKTtsAShZiOg6W23v+7CvOeCk7OfW2EVzWh
4PFkrO9+Psw+spI1Rhi1DNE7HaSCRnuBDdD/tSufXbQsUSrVW3my2x1ZZe6Ds1eg
YYz1IedTTSyxHmKIJHSXKJD57J0FsT04G7/ViJIq0xLnfb/6c/hR8Mg28NNHy5pU
NmEpgmFmZ4ma9O1Yk/O+JAEX3r8QllJGHdy+9IvcwYsFB2oXcv5/zw+m5dk/e2H/
7mO61uGNhQxyY0JU4Mg2Ji5aazbZuOocCM9bFXQZzeBjnwq2nKIkQFue/FWVQMRS
avJko4cXAN6DMsAsEUV6Z1+SaXs8wFUxcYIV6S98WgSal/FvXOWMQUNmTrwZxBPY
nJWzQy/Zg5CNxeQLIOrWndlBz46Ze6FB14maRoFx/HTo7Nuld6pJ4SkWsRWZkVZL
jC2qlQdziUN0F0LGNbEbZiCjFyBHkXWk+RT8FV4RCjZbZlrLQp5rAtwaud5pFAnr
QmeRYCnhJnXMBkcxtKRA9bleeqJBXB7kYfs9yHCqk86j3iGXGm87L559Ct7Pj2m5
0qBpytHPGjC4vgvvtjD5LjXsYZI8wF31OxG4f+b5dJLUdN0Dh6gqFYwXafof6jOS
tK2h6tBGsBiRmYAnK7VwspKFFkSIBf1QuU0h77u38nY=
`protect END_PROTECTED
