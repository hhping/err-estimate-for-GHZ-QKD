`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2W97H3uNfItcaLNvZd/FPY0VQlBJ7TpZMM3AqlddoWAfRerttUctw1xK8E4ewJC
l2WW2jVdXBvu2aJ2ucwzInhd8xSjZAz2FmA1QaeCmV5gtNJ15/Ui9Om3c2aZmvT/
bf5ufwMJ8N+W0d2CATkxt/Wmcm+a1kC4eaIiyga6ngRsGDHyyzu0pt7tke94Phjg
vR9PFqyhXQqUrRuq1QrKmUz6/VqQfe8Lw4PedjWQ93T2r8frkCZ2KMabY4yAcOxZ
DYxCM4jhN8S9cwCB6XuspL4C2xEx9i7hXQB+gSoozvjZxzCmySIAxftjjLYDwBNF
nZHgaKOV5wyVFlxpNK+irxf0cAYLCQcDWz9bxvr1tJry+X1SGdlgxWfS+dQafb5z
7SYIUrpuz9D8jKpuqjaTlQ==
`protect END_PROTECTED
