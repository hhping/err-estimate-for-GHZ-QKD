`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
szr7UOhO4ZjX5fsl5afKhtfTdaOlT1X7AL0VukQpB1Xa014+ByiofzUNsStTSfW3
a+qQibv5dokw9mkKHMSMIG5vMrluMFZLd99dSGRXkABJvrsCm2FI3TkEUK3BSznE
BG8UWUTGKYNUyN6uREx9oO28Hv6T7eB2EektHCIp6QDgST/2TaOMHiFSi0esTTma
SbtBN499bojNrvJCeYuMijV1Nm0bvTTn+oCxMK67Gec0natNFeBEi6TEUPXHOnQK
4zK+4EXo5HSMi++pE7mlP/S96TswUZxNuan+cWrRqGSusjfEGdZpthcaqJrm+eoU
P1fWqixkeiZ0KoZNzEnotKGNMBdHZdxKxH0bPnOdskSL2OU+qScoWlnhSott9wKi
gkPLcqQV9BnP7pWXDAW3Gt8Vn86cYEfICEjq+g0NQah4k5Z5gQMMhY9S4DzOMzKV
KF6nqctW/IH33W1ykQubwnhGWdggt3Y+stbw91++9oTIX8vWwZJFmZJa41MffwOZ
Y6o9rXpbvtHJx4LIgVdS/3YjfYrbPWKj/q0UdOEjWvI=
`protect END_PROTECTED
