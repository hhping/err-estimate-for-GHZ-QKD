`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qiBuln/55PqUTrhErwp8pR7U9X8ZtUr+R5GWBM6N5KwSyrrmqzUlgLdrQazhLuEk
BMpmYxJNKtVQ84YVMsiPw1jzeEbPzUUFKc5wpGqMclkOEftg3c+7BW31y79aDH7Q
2b84rkfrcM/bQdj8+xfTAslvt80eFSEZPK3ou3fSLzsWLhIEot01ammS84KIu3OV
uGWXIJO6QlYQE99Xssa35948TMFtCrDOtp5LnRfZGQIOIi4vq7Zsbo6cr+hu7fBA
oCwmEfwRHJtFe1clxxmtoIbk7SL0A6gR78QEiSPAXbIa3S0FCQtpSPOLRmrBk3GH
SKIjpkIAwF2ybO74jp0iJcERduKAIVkkRjwpfkYtZZ+PCWQ7zr4ihJb9wnfB6Uq0
8eUw78O12VCrRayhgweZSyhg0ZMpQxfVUF5CDT95aRuauVPshSR6pTXahSF1TV8Y
FreHVk3/ynMdZFgNPpHVQb1pvFk9xzZ8vN9fDeJUpQqeK9vZCa5mblmwMWKVDkk3
20wNjIK0Bkbxrv4+qxsMpz/KIgrs+cHRY2cm7vJltrFJ0LxqGs8KPkhK++OCuDJH
uvD2T75cfUUn4dBUY20QsHiJf+1CqpX8WHPronNXRuD1qgZVV0Z+CgzXB5StfII4
6JvOMbsq7IpeIRREAOvUHfvzRtuwP7j77GHYlMwjqRU=
`protect END_PROTECTED
