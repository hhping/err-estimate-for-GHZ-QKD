`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HLqSL5LcQTPWYW8DgtbjRaLHYkmbaHi2z7L/mtdINCmH4b64O+QaeAgZLgDHvpr
Ui3W9YrgLp4MepZzPQp0p/JpftHEhRuPpUO1OC2WWKA+slrWJkIfrPxIlqs/9Mce
VdbDJVyTqy5hFxdWHXns2ijB2TqsBLzFPkM/clrPbgGqndYUCN8I9w2DO8X1cBpX
5wcdjm8KjS9zzvj7LyLEX2Ektfg9zNJTGdyGiqK4crMUdtJ8AS+1DqL1FF9BEt45
T/UKYjUzl/YZaE+VqFnZzR1Na3SSBf+lSWnzXjtgA6qDFPPFXz4Xa/RNHNZrliCn
5NnMe4As1lRHfBwQeIWohAScANHeH8StEV1INIZXyiE2XQcW9hEfiXPotOGPo/m1
7zA1eevrovOReKzDxkbk5WhmYYb4I00gktKNCMP3vyunvtxd4H6IkP4/HAwGUaie
59BpiALrUHHyZSGPq1Cgiy6FcdqG0KO+n34FLiW0KeROtYABmhoT0JxxIlOgDrXf
8TzLY0yZohQxcY9I58PjOvHoT6pclD4cjnZWHB8S8g5aH4e7oBv4oGfTkb87jLfM
cb/gzt1K3B9p0Q+4HEspfcR4GpOYy/Bn7qw7TVO1DXMhcRvNfQcZGGOR7W7pwepV
XbKb0SzLYV/c8JEQcBHLuXIZfzwMHHoY8IgWOildHGWxuDnI8uXicx04nb46+JGO
MigAZXB+IX2nZoORYDIoe+Ji8nR3jWpqtNS5M5vqpLoThosRT1hwNsbXAcSKqzNM
Zl31UnY80yqdMXj2YXJV6J8tshm8tt92jkL5JIZ3rtp/mZ60kx9M58S0PMINJewx
ciuMQsJtZ3/FIQHfRC83AWMXajPuWF3Vnpua0UeIKtZTyKb6puFXhe7xT4xH26NF
STBOmBv8D7qWUjUSiLb1vKpVjfObaYyWSwRO4pWgJ3BowshMW1YSMtXUH0i802kC
6IU8XscnmFjE2KKos2D05EM4QTg1FyJTZW8JJKCsUH17wJoj+rVmkCql4iHa0m+0
mGJ60t26Uu578hMUDE4auVXmZsD/d+uxHoi6LUrc4Il5ZgFG7sc+UFVCWKoGMYy9
ys6x6bVJ+cpNdp0rR+yyf6VtrIW1jpQw+vIxmPOtUnrrCIYjUVfSC6OmEwZLZJeE
fwmpKPMLii0dwc+8CnQgQiPBIPe5W79W6OTU1bZ/3ulBsz1xtbilrznana97EBaj
K7Cd88b3ql5lpWnMcKXmctqqMUQ2Dt1bshn03wip3+nxpkfmxH4mp2D0MmlZN99f
wtXjiLoBeDe9VYrlhOK4pFdxnbjMoCna144wArO6hpgMpGhmu3VptxDtQocMhCO1
TW5ZLqIjEO74D3L3cAne5Hqnd4pD8YMqnC76gB6x+zSPXUV/GWAjAVlNjje9RWnu
3+RHVKxwdNsped1wcQIB1gS9T83u0islA7FEH5fbS0b45TrQ3xzma+xkmMXTTBMK
f3BYOoGfeV3s70VV53viBz3aNdGQ2FeHERw/KsLC7a9t/Viz8IsdIze22ZBFelD9
r6TU4DXsnLeQlECn3JTTEQgrAqHxgRYYPYZRCSQpWln7AOxgzdPYnpRNh/wayE2g
2LG2ZuFVKC3fk2FbtUr4lONvnBhzK6Tc6fjzBHQYmTj2MGzKGum747MiNuL5lqDO
ghHGajNnLKxejrWlNVxQa7+uCxZyPKUljwnmwgUw2oQtXpPChry6u6SW8bypFl+T
mJKd9el/N9X/DBZ5QoX9pBdPhE9LThm+Th0TJN505xc3kS5Zc0MC6fNYs43F1VFt
oQuMaq83+ZJFB+2o9zGIuhm797+YfPMMfN3L5Whcxf5B6VzsGYajrS/idFzTKZu9
3mmKtNzHPdfsqcOgXkRsmGJRqZVde3c6Uwd5SQDAlCRcVI3zQtPhm5cwkl3QFmh9
FSutuwLIv5dhSqrS4TL1ZlZT45S+2RdPjIhF6yRSWUw0g3dTfnIpOBj+a2yMXnyp
TmbWPzM4H+FADHHHv3Di/Sl0DK2AZgRzKVycTMych9e1kMPgbwb0BR9sMLkhnr+i
XDkICUGTKxn0Idj7kd26ArvD9nmC23kGOn0vqtfJoA4p8L3tnm3WMc13rAsxcuYr
z781vjmsCOIe/xmjdxQG2zGz+PxBHAPAguo5tJI2mG3NcflhUa5nv79gtOl9xEOC
fXqjqSDGf3MtdXK6KgXm05tUbykH5wtA3Vi+8DyCBkYDn69DzUOKQynWufEPalMF
tWDz+m4f5D3JtymGNf0YKhcqdHA1X9AWN1QkztF90oMlt4zt96aYRt2Ko+32Medi
wFF0UO7KwK+YrThBzHnKGBFFuSqAhqrypPrajSqkiBHLoUgIMwUllLYdNQmRV3KE
AO0hQmmhRbTo1RKKypRUW0Dr3fY8N0dH7NFItS8SP9PW30UACxj8Zcu7qcGpTMyt
4Y3XkElaCLle/tL34FhjUtwTd8jCTQ+A8yDsEg5p7t3I6/xvnUKrXMNqiKSvpCFK
gbRR/T8yKXZGiZ8sxVAFnlMGDJA8L/AB662eCOF3YCkPz+u10rpJblnAZyzXWnyH
Nz2055Icdr3LxOiJdL0UzIG3nj5rEYdzNcWU9E5PttRgQVflJo85a9oyRnGLj2gf
JrCyMrHJXqbwckiNe7AjlhJoEg4VnEwCJfEGTMhqUvPhOGGd3h/tuR4ZzvlRFqEn
2ZFQGGy5Hz0zjt353M7/fb8ZQ63E31zSQzME+pP64SaJlPFbClaaoI58NCebzv6Z
dIL6uGDJEhmq9nEkScNSbrKxhkUkBB1KJc6J5aIZm2qrNFjS1d5kshGHr8iVo1o5
+UjjKGicK9ev97l4tYaIowSHodzSIpZ2j9ekZDdZUSiwVk7E5jVlP32ByluRsvHs
eOoCzxkxRlq8/iFogZtHbUFaxdkNlOEN5IwhSoU44rMCXBiSizGfoGkgSFLmYCEJ
MTI85gPmG+nq2gE4EqhlWZxVngdTlI2vXM8PmkX7g+U/SZKBfjkua6Cm6J57PQzN
jz1W988x897ErHnsBaqG9Yj5V4rEKbaEfViFCQYsVq+BrwVTEUGhyrI+gDqjhSW4
hbAqzSRDnH6RgkES7FP9W2KJmLThK+xE6gn3xNn02rY+eDt3KY4pIPf2mZuF/4TV
8UBM8J0DgE3gcU2Lp1DpTa9BfiAKcQiOHABLLtJIPc8hn7dne8zTOR+0T5LxJfLJ
afFRSMsX0eAikcKBmvuuDQ==
`protect END_PROTECTED
