`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hEurYWtj0FKEYXzDi4o0mNYPVNAcfNVHQURzj18c58GinBU7sBI59L6yxJggc8AD
mP1WYYLb0H3R42YtAhIyk8xs2OaznKPkGW+l36TbErTgwf8wPzb6afG8CxD3oPpe
LSiTT6EMvUgA4DzzXnrJe6ysHY12yXpinDm0aSIwcns4U+eSbiiD6w/98Knexgv/
rUhbesRDIclbyAEW1imkqOJ3Pa0nXFJrTg0JGcJ10lwnDWmvalkII8x6PYPK3lCv
rp2mzuOJ38/HOekXF/DaAw9KkGMsIY6aOH/x3fbso+svveZfo5mRWc/LkxSRSght
ZS+Tp34U/fFyXVpV36/rD55UT5bf/eqLYaO4eGkUXQdTIanND0IH3YoPDrD2tLZP
IaeAO9TeHZGKOI18vKILv4263NCaOsqoKb1BLp0EuIXrJ4P+3L4V96Xt7OkZt5jt
/XrALRoIwpIwjCoMBEbFHLeIiVTxn3UpiPaElgaHw8Ov6WoLd6WqAvrdcFDErAAt
cnY6TT3JLe/VHEJ3JuxRYkH7c98r1d0TvSzmq3rbjFLC/F6ewkblA4rKF2e6Yf5v
fslIJjzRgzs40W2lEgnmgMFo3WAZ0sNtheTcxXb51IStjROabSMRJ1BKmy6MIECr
uoQoQbLUIZAlAIysn3tt3BPlSe2yZegrmir+fG2NjuKPiSZiDEbLnfUNT7GVskVQ
+xyevoqd9uS3w1TD8jOxybVNLTE3PFhrYNaXg2lxuiYDCiDyQ5qaleAXhZ3eWk0W
IFyvogeO0N7iXd1uCTk+Vi9oOjtg50W5AQg+9E7+dR2gx9al4w+e28UdKsBVvfkN
FoYJgabDIeQmY0YKBcWfy20l51SvEDb6lrJXPnODqNNSE/r42YpnpGPNNPulXkZx
1APen/EXV3FsRDmt5MKyavRbNnUw1zVd32+F2kexxzH0jJ+GDS8XUjB7tOpdcASx
iLPsz9wVHn6oN2on9StmGg4G2bLCeXFVcsYpBOlzcy1wG3YCA2i/3MG7GdmChALb
xRpiExoVE4V5JLYGnZCRkr+IETzsGYO8hLGB04MdnhKa5wQ0Xp2VCq0Y69ngYjbK
8V0m5RCW+zJeAAFTAwd/K5nNhf6pdgSCooGUCNdTftB9SWGgaSOrEWGYm89+PC10
GH2nQktQ2uCjOnG3TMBGzF7zMMrESmJo6xr2f7ROj+Nrg2fpWO/c60PBBH3izXBX
YMg9aSS4wHT92w6iTR+tonp++gBLpIMZgH50OM+VabuwI/H01hRlYWSbYbpf0H/w
b05DUEZ5hSBXuGgwT4ZahnGGC/A/2gfY/PThEDVEk45hE+uWJwevUTNGwf+hgmRk
zPVOnZQlgDlejrQfvE85UP7Lv2nqkINOAZQUrHGpZI6kt7tuGoDAV8tAxbReWVzO
VxVQs5eIrmnOq4sFNVIAWvcIGDjueFZ0D2xW5jMH5CvQAZ5xbYiyiTy2bDVeZwNG
L5xNtLzGV7PMIiQlLdRz30ReuAyMAV1var/vV+3t17g5JlFMsXYPwpFk2dsk8Cpl
BRLtBDAr1MQhKYbqUJTHxJBtn0PEYOACBUSczRwugCjrp3vqXOgCgGiEjUjGW3oR
ZsnUdfVe7Xm5VRElbmnOP4qC7ioSFvlaBgSgG+MOpFclxG+VfgmoApYfQ//wLF9a
E7Kpo1sEpGloA1mJFxUIfIMuw3r6m8/e0ds/nMsIVRIAQtg8ElwnVoRasUgagsFS
fXt76mfgd7nkYD6+zJfeE1rd7SCvwPJX+67iwdQ7gi3iDbmIry7Xq6pa7Omf8vmp
5a4l5s8mtVrzXLDnGb9zeB1+UWDTKFDPWxTt0YBrN09A58y3gNmIG3vsoUnZpjYM
bQVc7AtIb3/qnbExjRULl945pxvYts2nvSVxW0ZupGeYBUJaqJS8/du+sbMTIXwr
Pxe5p7i8qPF2qKS0TZ0TeeR1cz+eAzaxvdQ83OdANLZ4H4CQm60rSx9mJItSnYBY
OQBRAhYsaItQtwzCjEOZ0qnX1AjaA6HWBJ4AaHTUgLqwauvYFh3SrtsKuULUQ0lW
XaesmJz+dZ2g+K+wFVc8v9FBNSbGCDMysymKSZMzPlzpYbcrIyLtfU3/URKl/vWD
y4NlS/r0Q4VebAM8YP3QuvtfpAirql0MsLquprI7Kmv3Rqp2Vmhdk2D/U1mcefB8
7a2hxfB+g5tGj+rlnMDblM8CntTHmhjbXhKwXRi5XVJbTddi6a7yosWY6+CRUSZB
/Tl4Z9tvoiKu9TTiGDztnil2KFUsvya5PK5OBT3M1yOnxCfmbPTv+Igw2X5lFaiH
lAn10gjrJdng8XTK3sEYNC+z4jlcxQjajR12m6yC1LSZMIBVwM03GBM1hvhSb9x/
UTpsgDSMt7tlTA3vUJ0CMniTkrXtrWI9TXDWKWLWbq2VWo2O5GZfQ7v9NkEi6VCw
j4/euycjTFQXIOrDJ3epEsB05vs5FnwNY3pNDdn4K5oLhMpicfmS7dQYB+3NSx12
FWq0mt4pr8cxgx0xsVVkWNE5NCZQLZXnSGijhhE6UQGkPc+zCAPramqUogtM18yv
3e0DguFI42rRMULaJpktLu9beFoOfhqlSrQMo77pHj62cNtQgvrnoZz/mqfYd2gO
uc66K61IIAjlubmzFsao9p6dHM8onrHfdJedq7T83OE89Xy7tRhzrHActbjsofkB
L1HBf45GdluHSoBu/yDqeDE6TSnEOsmCdmqeHNC+xX+jOnfdfOUtJHgFlz2CocVd
i3dWDnqzlFMIrxyTITJpSXtsPGGcK837xrOD0iDU5aEPiumKhNrLIVW4Ypx3Z3/Z
Ulimf9kCkHAM8wE6HTGIaeI4civiX9oHPTtVeSZu42hRTHpLBQqwqyzMCr340XaR
glkgBzHGfgTphJPcEKdxWR56fOJGCbsk7BMuN/lcVxubUNrGNtq0Ok/zAz4Z2iUy
zfhf7gTr2NGw33BqLGhTJfiX9JiTjdhCug4LuvnjpeeNp4bfuTCA+p2KdoYd1nvt
9CjuUDqitJGerFZ+BUYISa1dxqQ6WbYqnF/OrDdYRsADxalcH3eAKH7OHxppTHKN
zkrtrC7Er3FniXPI/+/ZZQDF6IEWjP8tg+1Zm3GaD2TDIJaLsxPpC/ot73/rkuy/
Fxa/91mJfEjKGYHAdYpki/aZchU8yT1zPDatziut3jQFFKjTomawWeSsYEUfvBqS
qZf+4fYomWvXeVjA5u7VcqsOJ9ERxlCWmgs3G4B6Jqd5WeQNbycq7cKqAFT92DFD
buEQeoFbizTLfkiYy4AaFJp5FckPWbjTyGKqqtblZWkoI4B2+fpSS5PdXrfhkch2
v1Y7mDS6dRpBK5t2hSstEip6nH2PO3WWV8JFPJXLmGAj6IqQe/eaXOLZ6qaKmkN+
gBiJOpUcBvozF3yOMpWcfuLuCnGmLCTDgikuA2smhHWGBCeJXv8vCmLQG4L6BLK9
bwZEilXOQNj7sXx+m14mLa+AehAVLdndLkD31DADfCUuIi08hppI7BtjyUwlNg66
DADQLW8WgR0HAMHYO+73N4L8ZdJwHzxFu+wq+32RfIykr94eetLtVuY890C1mjaS
B0cGcGbikbrZB2j+t4NLlmOwjAd4/dmwQCxEqHT98tJvmwqt+m12BVpc50dLRVRL
Aa6kD8dYS7YFtCXxCGE9r1cNpm3JLWngcpkYKk1E+A7Al5ZuwID2dnq261/luzST
VgjavOs+qfHaHGRsvRELIBnH4VbYqRlVlVjZEEmJmOQu+5mcyzi0ymjD+cOFEaSJ
3+u9uK53WtbohuZnCX/Zy24beGveQTFqKlvsRht6yQKZGGmJUh3LMGr+ukuFjqKS
KDGhnsuZWM9+fHc3q4Nl1Mgt8NnvLxck5TKj/iNsWUi+3VGBmW4U1BNnNMEQFEDx
Jd4NU4oMPfEUWzbNWy8HEjrVQuOrUNwzxHZlMz7MrEOANXPTodK9jwOEevNekSuy
o0E594eZY6R55X7jtzP8lI4DHQPxu6KIRIw2XFHYNUIN8k5ZldC6VlAKVUn7yPW4
ThqgDhjEFf3eCI3N/cllgRZN/JgRS+Pmtx2JT9J6SH4du/WX94vFrrOdAYj9xSjk
2Gba471DlDJsftxTIVQLLG+Y68pewNiE2PJqKOU3z9R6qIuMqMksa9aohFwIq46c
I8kCGv2PvRbxt0MWePTwn6VvDIqO8UnStkxHqZSFKPC6KvK3s9zSyWA2eTT9g3aG
byfX/7H5skriwR4qjdNigcAHFWUP2w8JGxPOMe7O5pZTKj2f/6sqqdi6ZyyLxnOS
cpsqaNNJNBVhZOkabZpDZUkaD3ivJAgeH2SxrZ4agsBJhxUFKiLa7obGEmZD4eKS
KGZZTeKrmZswnRMT97oWBJr0mj0ZitDit4FdxuV4M8FV2u/UImZuPELr8000w2XY
zEwZBZ28i+4AHxvHqmOwT9o1KhVJsdIzwB67o28i1ERvV4JLSlHr18r++9n8xw7x
NZIZ8nrgo54cfs7pbwn0i4xAe9L3isnsRespQeNBWHnglvv10UrfIbLFeRlJnvaq
PQp3h79ciKEV0wkVYjx0cCZkNIO/bCco53ZA32CDVv5QpY7+3lsyg+DILvdbKB+b
42z2p7iKUd5qHjGBcI15fNxkNuaBg0ae0Xhtb1/c2YH1OBqozPBZKb2uRBwOFqUt
6a1de8IX+ydq4islQO635RNxvgE+Imy4Ix0s1Y+WG6JMQpA6n3JHrzTJOk5M4XgL
NlcDo0fhmWLGnH9BWX1xZ20mOZiWmqv5w4Ad6SjLMInV65FW3rJD4FWZDVuGXzC5
dsl46Jw6/scz/Q5Keo8C4Uf0CJMd+Iza4XpuneaEBHogN1x3ZvSng98YCu11UG8o
W0WkoaburvTPKYp9vJ4uF4gDPt50W7xgjkkjW7c02s91cA5du7310SkV1TYTs+yT
XCY+BDGOpzL+B/4puVY4BgWB8Ba5Mpm1fsDr/RnC4IZb/RWlv0fF+JC/sj2DovO7
3cTBmbivFCuyu+UHF1Ntq+ox68KlOpAKoun0zMAnCT1/dhzbefEAIrsaTK7dtHZH
aEUP/UfPRf85Id2/UonYrC3OVxqSJuafQ6264hWuR+AXW4H9uMtsGdfib2asvK4P
5EsLNnukeuGX3pDjLFyTFfX4hcOWjHAb3ZOWtuAN/kx4/sqoXFUHktWONdOY12Xf
o37OMuUOTtfpGAo4stscv4w+OszkQW+9wPHmBHG4oXjd+z5XrQ2qhQl554JcTdzU
471PYUnnrMdIFfg8ZsM6IQKs45+VuLOlfH2G/4BC6pNLPgPSZmW+TMhR9clYCLND
VV9qlegu1HM/OfB4up4VQd7TvsPE8fo0RJhOelz6q97MEhmSznT3SjckREOoz5PL
0X3ar63QCZ24Ori92cf8LAtKJqShaCF8z9zydu5Q2o2F/vij65Gkd5PgrBCmWRTr
h9JsiqF/ekiwM6ydeDUOPle4xc+F/tZTMcQURB8x9NadnbaW8qxTLRVMB72Sv395
fjMiB4Y7vocbZ6Xn2SqFlKOT0YnNBR8ZVJ+35HpxHMywWHpiwrVEsADWb26ynESR
jlo2yN+3iCKhwARi6KFrak4mzzJCt9tr3bp4dx77r3adDiulIH+j18a9207e/yWB
Q6WzrB8kHpwhg/9IpEFRItprLRHHp1//BIGU4RaAGzGHMPzCycVN85LqAQJSi0oY
LTzxYAxF/CuGZmodiXeWKcOe4iee+zucTjtidM7Pt8f0ndtaEgRskE/GHNqJOHg/
MKUhSUtMJh8h96IIIKVC7XvCp4JpniTuRwPjw8EjFIeXLhvkfPXZyBZluG0J6u3u
EAZM6EH9lrgWAc6V3ktHCf2VdknnUP9lRI26xRbEu//TXqJwPpy3KBrYYJRVwNPx
Vl1PsWb4d/0Xfci3YdbBziqyRxQC7CcLWEuYF1xVpL2aR2wIzvSsbucrgdaMrpH9
B/ItqEu3nDIrAWd4e/RI6tLm91havGlNLzhNXMiz8ryedM7S2ToN5MAPCOOL7Xxc
awYQeM8R3nQcPJBe11gHFw/+pJVC7qcAdXm6avV+3egS5/57NfeG0CWQTw9DAWOR
yRtPftSS+Ry/oDhIsqMhcWBx7GOCENzD9fomCTKhFlgSWRY0G2Cv4ThN+PdOHKcR
mpiKj6QUEnnn77gXVhfe26mm6D6xniT6xuh16crcA9ZP6MSnZBSnuGlGn8jUvWy6
0DZrqOoYWurhdJk3TL7/XeVXShwI1QnaPWolVq1wJHCZ1hvxf25tZrVp1qQzwpKy
fMLgzfNLvt0TKDldO/edhINqb/9CUjRRJT+k11qW9C8h+nwuECxYpXhGyDf7a2+I
Il1LsWjAW1RukModndR6x2Zquj8L8gptMUwbA5Co+uymTfFgWyUqFDGiLWMA2Unx
XOi1aOYQ45PRYOqLIL2R8iD0Wr0atjqUZ7B+YWnwY52AOpOfsB2bVmZYCDJEnTUJ
r/Q9DylTjrksFHa1qCSIYHnwLAbNXxl4r6eV9DmPpp5Lv4LZ1gI4ZI8TJ8/CSRHf
z9KoP9In7AlTsM2YyX6DJ25M52PGeNAsEpPU3Z6OUnFccBcXLmpn0d0OCZbXHruW
DZ5JrdNJfCp8v9gji/fw96JASG8FdI0Jat91ozIeSegxkqkKlLZBmeLArMNJlXJQ
Wg4wAXLm0kH4EaYSNtYKIWseFq5rupXSmTarnV5coPr+3OtEcDPtgx1PFnoXotxP
+y6zELHO7nX0dnudjge1bdXy4/x5xO0uu17Bcmoazkj8n4S0DjNIBe05MJkgXhZs
VmX0CYOwYFzr5mGTwo19flaNwTs767SAQu5fbSlTZbwBDmcuXJ7SMPpMBm5cn+Cx
KaSEbgtpuICL/ZoPmsYTAemINl4d76GrU8kNT9puXLKuMBJLlePZggOAhTrREgUY
8X93butAjN3xbX0x3buZuqy0CvTpa60unNmOBbF/DrRUQ22hN5P/hmELrBblmgGu
foshxjRiuFWDJHmXpoX90Jpy3xe6viFT5Aqfymy1TinIlDtPSBc7aTR6pS4s/c6x
3VG39XINZzNxGNXNO2h89lkMrQPh4sEd6JkG2SOE68kscZ3V8FFL1+TLR/KLzeRY
dioz56VvzUYfgKdGaHgJuu1kqs7uhgbVQJlaZn3frJ0eGmw+PaFq6xzpWMk5PqS/
niFsXYMaNHa+KiwfOJRVDgSg1St/gfRCxKDyCQqKLRp/NFPpJQjuYAV/1wDPPSWr
RWFpY6ZghItUE+cfI0Wrq4xaa5OCXSm7F2z3qutlm3CySTs+4TrGZG0YI8QbyLQ9
fxVLeUhPsLSgGBYiipPhNrt/iYB9xEeSAij0ioHfnhFate4CK3qsWb4Utx2hr9MX
dmqXXM8t6RSL4tJAqoLcE8uEwmP/Ir+rVL/bGoA/0kCZTaR3aAkv66WWOtUM0/sw
MqkDGSjUAFCt85ldL/AMZg3bd3S4bQlmvnsB0k3v+2QpJF4ok8hONHAc18JCfmXS
6o4DC5sdLdCRjUhmxPxdiYgJ4l5/QZKUb5cmnpMdffhvEhjoKjKCA0bxygTo628I
azjouK8FQ9Uloo5TKME/BL83aa5pl1KtYATYbX3MGjrqzwTmaYaq88OUFfyMFEOJ
bDbSHJtdVxmzWxQIWNiREQHJq9cmMgFt59zIepn2FJrC01BTxWLN8+YuYohhF+yV
KNevr9aKo1d9T5MKnLI+fQo7/7g7DX1iOl8n7CaU78ZitV/HMHM1RC1IMASDT5Sb
UFpbmFgyLENsz+6D8AuJApPx7PKO2ld8/9Typ1eXPNZgQZ2uGxhlzk9K/UiuFDtp
dnQdwONbTB5waW0kFKitR4w8SHWnDv66RdSvNjfoA1UZwlUkkNeKyNfQJBseTy9B
oT33h5Mapd7nwJZyp7Hz3O8527shWxqKmkGmfwfyr2bbpErp+bGOa3V5Z0zH2ZSh
rY/fjWT3rIf4ONyTJ4oBcsLPDU2GVLWBu7NYPGAoG9Q4gDaXW5gGeB7Fb+TTXJMA
nybic+RbWASaMcaZXEAu01/zWTxe6zTaPnyMEcUSAjLeY0F+KSAykMybV2A+p/eO
Wud7Mz3C+FKpgnQqdXfYU8GRcDH/mhQrd4kJtmwGXxRsLoH/NsT8o9lqXY47PzFS
QBuXxaOBCx21vMIhINoAGML+MoGV+P/EiNU9x6Cxc18itu4LKOTtQyuSZQ4zG/nk
kYTadSkOvzfKZcX4xqYb3NQpydtUg/o5dHthXCmmqiS7pZ27webBlLUkiC9QoMYT
T2K/BJ88lYguHhkASlG65MrNm3Jx5sUG27F+30tB9A7g++e34K7B2ThH+3oRKfu2
WmtQcB2rL0EuR12Me/VLkr7cyelZugFpoybD8F4YVX/eHYdehAbl+x6pTNn8H1dq
QhsWbapYcH4Dx/noU2XnlLZ9wz3mh7mnqU9foYKaqsQmZFcSP0tGHWofNkob2Zy1
oDBNeeqk/Ynla+Xi/fcQVaBqKeUZQevDuPgn2rUecruSfe3aawEzmhrgnGwNlbPr
chB6v1kZOTymLhnZSQmfxIdOniUW7/0Lsii6DVu+Bt1ckaTmm91F8Luk6QA21lpA
8QKcNZeHoywRvomZ87PoKzuTeACbIBHxPpL+F9NRkEtz6pD9XdTE/vN3czvC0OKI
CwbdKHbv2aK3o5t0MHQN18mg0x260lDtU/B9jM8wh/OPYbbthYglS2qDJD+y3hct
tmM7F1QDQ9o9waCj+TTxYSRTm+xPFY+Io2bJwpAOE0HYBBBRO0YddQVjiQ2t8SJm
QWKS3hfkaur9tYTDWeIgj74Y7WL0ATlTgQYR5B3JnHESQmCWKHe9b+faRXvqdiJK
p6Wu144PYPLYBj/o3sRZZtc/2ms4U5PVjTYG7E+io/DPCEQGxw2p++QGsgJt6JEE
FLflxilvK319ndgxb3iCshIY2dgc5/kQR2SAcZt2HMFO8rRtgwORObeuMKUv5/Gm
6f5KSCG1bJBJ1LgGB7zE+SdpHjwDJJ46woQzF5VeJvtqpI+W5gU8IuwZcX6ROMyf
XWkzRoLo+bWH/d1qMlKAPD6IzJz+BhAT+IZf9DAJqfjfAUbacyL3pS6+N6bw+TBB
fOLDiq3PY+5IRTS+jRkaZaJP7yOV2iAhespowrGCUxrZRiGTM9RaHyG5QOyfWLpe
DJIaDYJoWjBiuLIYQ28L8vlFGzq8SkojRmU5qpisZTtZj6/lYaBhWDBrxy9iqX6i
j/8cWx7iUXHpDoahvK6YAMfG9Xgt9Y8UncROrmVYb6aWP7CnuE+6iCSDcyUWsTw/
DLrYhoX5SXeM8k5lwabPiPYFp3vN5LD6IirL1ciM50bFmbMDBBNhK+rLD975Ejy7
ijiToyrY4Fo9kZ2OoBYSOA7KM4vW/IWtjg48iBxE0krNknE+tn1jHhk8z0EVBVio
20rG9gQUJdj9+isEFwLdc1mrtwiBAlc/5PwNFoyJBcwGFAqs/jhXDdj3QQpTpx8k
3qJ9b5mQZrumGWdohSpiDIX86EhabOsEi/3AZ3MvuAk6uyw1Mm4YaYKq1U3r/FLe
AaI5FVlwvxdS0ScvmYFnJiFNQVPKdX7Es8m4d6AbRMncpWxqhssoE6M7IwwS11Lk
pFDQ/sDMzmanuPPSzBEeM8Dc/vjCE255TdrGPA6qJmbieLxQ/nbwYJajcq8k3sSn
Pc8AiyaZKMtIkljB0mYTEvFPKg76PPETvRnKRlH75n/Mnt8i0ECu3yh7rQXBKHYc
SsovAbCWtR4sDSGdNcfYM32/td7wnNOfiBiFnuKwP8s8R5cLs9pMi41JsbqtvTBB
1TWje7leATycShrPsGKbDNvIdVZxfOau3IErJt9YtwbXvS6WiDacbfmdK0oL4h+Z
pFcePoxI7++DcOL3xC3jai9r3dg0Y6NiawWVvUhfBuAO5EmUk7thATMaB4Ezmkn4
3tuqz6ttREfgwbbmp+wPu/f8xGZGtJJnMS7nmOmr1H6OL1ydUl1rB2KM+Eri9jUE
yOTotkD9Up3NRlLqHt8cCj9l032WRNbt/ywwK7HtoHAwftsIgkIz/mfA0VCdzooC
75mXno+mqIQrdLZLvWDVkOXinA7FZp7GzfERS4WvxNqiVvYrexCpwq1f/Aj4DXO8
UZtMwrJR1TW48hfGqRIQy8jOWqvV3Ul7OOCMj955lZJDQJkyGpLKAuMLSlH1tV64
0uTIVgnGEy8KfXWvWk7INqBnJwE3eBJ88AHRH0QId2FGHrFjGtWVyRxC5Duw7Pc4
c0YqzL18wBN5sFkb9ORyejZdsuOebyiTBEitksZdbxweue3PqG+oHAKVri7S+h+Z
YFRV8uytDq9uUTjoSZ8Z8Bk0b4v0e5q/BkIFvIfx/aUNj6HkBVUW7YBiJFayWLzM
LKf53xglZ/D/EKZkQPnuvPsGb0jdJHBUpm3OWP8giGURpo9UHxTjKga4l1Ref+zH
DQfXtdP8TPz7X9gJuYXjJrcvD9MVNf4b4S8jqr8mnbh5vXBbY8TgOXvJ/vkcynLQ
PjFGiZt9bc9TuHnW7s6zgbGc1CvnsENPRfCzIbcLJ+tuTGBHEDr58Ug2H1hAgPWi
+gGKtHqShCLMNtZUJ65mod5tNN35b1VRZC1xK8sfS7BqWZZ0MoCkSBbEVbKOU8c6
DPzUj66+L/5uio1DifaMPs1QVYBfgafmw0ttmwNk8kV2SJPMBADOmDfygOGwCjL/
d2kSfeamWbJi56u6y0bx6UB6Rt+58s4h6Gv3hEixQShvDIIMuUkhgsqR6CsRWqay
2jOxVPyOKhJVUuAc55EiWiswJCiTdkicVymhDrMxPdUG3TFCABVRjTvPokNYhnUC
KGesjhPg4e5PccgMr+QzSFDljTvqFCNCHkHNHJyT6wi7jZsxuLlG95rLGFynEOXe
jrzovV91XJsTkYJE/WUzS9Ism2RJFyCnaM+pQwVfYfVfvm4RTYD26bOB2dq6t/7b
rmuXpC9ulV50Lb52rw30fhRAuh4nwkGIBZWTUrxq2kVvAm+ovCvnQHlQGRvGNCig
uEY3FOgmuekb60/9hWkVOOLWC/yNlV402a/cINvsbSyKYBJUJF+CWf8+o4mjrY9l
acxCYBzuOU/RhFK/iIAhARrfgpDW2iZUMh++FKmSh4My+VOEFtg4cKqS5kwd7fuE
dTwIs7WlClmxCt3nNuqD0n8XQWooaSo/X+xr1d0tfDQ=
`protect END_PROTECTED
