`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YfYEf+xDPV4SDwSQTn9Ep//dsHiyS4OHxsniKk1g06KuDonCge/RmYVJED05k9M
txb6PmRrPJZhvntPqMhUZbQ1XVvbNy7BHno+ZbfaacZhmkDe61+dsjGRwNimY/Jz
YxhP3rJmABK6W45V2V+paVJNlWfTkUoQuMBt9+THiioKSnXlb1pytOiDUivLnQgq
291FCm/ZgXHu0LJSN6DOWDdOOgOH0TkuCrrOc/Z6oMbiW7nn6ZppJxWBuvqm2e//
gK1cDfciU+xXnTRMbaesCQmkODBc/RzH/h2alno5FTzilJBsGB1Z1XRproB50UPh
MFBs/ylg34qYdG08K8zbOu1C8wE5qyrRS3f9h9JcylKid5joahKlF8UZngJtJOJ1
hnYzG4RG5z3ybdnZ8yWksw==
`protect END_PROTECTED
