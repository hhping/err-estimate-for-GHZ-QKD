`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAucH8JOPmKqEVQNFRex7SVl4qOAJi0RwZqgVrZrvFMSf5YFQUpByRQRuQzg4oLw
/K7+QcxVMEgWLigsUOfogr0/SKpp9yRjRJHzBawa5KFOsw53ihtqeDch7VBgjpkZ
5uaimeuvP2uKQJ7ulNBNSNSiqbQJ25nDqhbjSjbz014lOvjnxOubFDiISLlouZfi
53RCDGClIbPsquXh6W7xeW8KijxmkqG8Bco3edlskB2bGCQocO2lTHYbaa/oqqOJ
wN3uBiHfBB6Zs9YZvE/q644f5l88rdVQV1RQY63T8wNQaCDYmQyZ/oS5P1c3gC04
WFYCIZnDRM49+KVdsiHcP7SvKvU7JFklpGTwevjbLFfYYlqJ4CrTlwC6sI2zDQZd
dA3lRbTZqmQk+3dGYgEtmDPBMNZVWQGOq53Ch9LDa/IgiMtDh4dVBy9LX8q2bo3u
d/BTX//FeQsR9KccuVIzZOI346nUBlRtYrvzV9fRcIrGGi11fJGXnnHtegnKtgan
Ik7Um07RLeUvDRd6btiR97wW+9HJRO6NBM7gOlc+RgyUhhiVUAxPP9kzIEhf53c4
oC5kNskqLxc89XrltcWXEUAB2YQ9kyuosT7k7E/2ldOFdO6Hl0bI4f7AFos2EDgH
nDq9lxa013vHgElC5EQCra/XIpjZowD3mciRv27vqBDrRzy50L0Qmw/Id5bnKkdG
F3CEjyI51VnCRznhc4E/RgXDTNyoi4etlMr7A84YkeAvjpoI+cOU18AYyC1ZVEew
HHFQ1jLJ0YbFkXeJSeeckqQNLxCII6AinvWmfWeVR2qcNgd4zy1XJXU/oOO84TkJ
2oOzA2jPHOCpe8bDTgV6esW/uQQItWUgNaE69foCDYD8ZVAth/wq6SI5JmyC22Pi
71dV5XeHXdzLZpXx4J441Nwdl55p3wA1l/HnydgCsVudmjEfUY9TFZWGy2+/yaKE
ANih488TdukPrAyPJT7HMTfkryzRn+W8kZYK1dGUyN852QjCf6pTfKzG7pe8rPY4
5Zo9orI+binY0acbW3fSbhNQ3IemuWN7T3yn+mLTwiOD41R64hFrO4e9NJ0fnXj3
Am/ANM6nM6cp6G0xjuLiqgLc0O7ktC5tBinz92xxWaKJg3B2raYz3z5fPrR0t5Ts
XPkBeARiE3dOoE13I32V8SSkMTe7Oa6S+71XJflnEjI/9VxxfD961IX4uy8Bjq4W
u+hL6hv4JCf7AUrl/f965/sbbcgpdWZjKzriqhxuBoXicsfBXez0Ss7GKZbCrz6h
3QnCN0+D8s0CvDNUsv7w3Cnuyyg4y/l5nLmShNmU/9wVC5dyz/UXXZ+e0lmbK/Xq
6eCxgis6zPgYQ+ezN1EAyIKFACyeoImwv+0Ge186oQj0GgxTXQcU1N0ttcS52HW7
j7/iKGq5Dv7KDJnkFh3V0e6fjkow6KctEiqUqrtURuflUwzQ2a2NZxF5AaxRRKcR
`protect END_PROTECTED
