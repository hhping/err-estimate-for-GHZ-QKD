`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkDA9Z38a2k6MvQPkT7P6uqCGafdXVItvbKsaa2LJE/msscY1DpYbwNFU9FPrbSb
/i4fqPUrSqFi/xqCmd8tUWd1U7WCyUCnJJz5oPmwuUPs1laesVlgw2lsMBune1eb
8A6N5hD/mgKl9MkBBw5I1Pbm9XoxhWIfL8xgmmj/WAKoIqqMewPsZczj/RNptlW2
IzB0sE+0tVVHMoLrW5lHGW0ExN+jc4VV82MkIy2JCeyLIC4vv3OW7H2VK4Rltt4L
OCu6LNvWEEWIC+aWZdnpaHYO6G4nzBF7PSyohRTC08tydl1qkoCSBqFnQl0n7I+C
SZcz4aCW6PkSe+Sb/6QqlZrBHJf2zJPqZmh9cewIk6faHu0Z41NNsq38RxwHAlHo
UZbW010g64KuTQw928Ia8vL0nmZFZxXbWpMbdPVr8N7UoDwAk4yDjQc6UGAJZ50t
fYDKD5vl5HE0SW3BB8ycRaGVU7Brn4jZYPYDq7Kgsty1P0uF5KWPM5lNr7cnJGXk
5K/TfEDvnQPukJ8dul0nnFiZxFyiCjefECI0yw3jkcSPQ0ywqKT7axDy8HRMcRPy
V2HyxTV60p0Zm+A8bqhuZkt27Ohox+vGbSuNJE8/NeqmPlvgbRWelvbu3s5Pq1Gd
y3KZ/S7jBCxsAkkS2ycC1u38EB2433ugT+NSSI0JEs9FutQQ0wcW637Ci2YEGxoy
J1bEJyM6TGrQuPE0NqQYqyfqSNJ0h6+Hu1ZqEZ8feutwCcXlfs2dGL53eSm9AZeq
x6sO5oi/H4x14F8wdFGElHwT17qiRcLnLRoQyVJdtva254qkuvjOvq+GDv/M9Ie/
R6DdVtJg7os2eeJ/CKrxaWNR2/BP3ImfNlZL32d6jGB2Eod8K1AfK2wewoUtl7XF
c3yCrXEg6wcOiigvg2wZTiyy0n5cugFh9h/6vZ0pHsOuNWNTHWwBckIEcf0l45KZ
jbyfJWirGJyhg894+BSCcW9xlzp0ILpJB3qCKBUuIxJ62xdLL9+Bkvs+NnxvKJvo
PfW5UuG0+AkKjQI7DG9Tom4QRqXdoAvAH0Bs1z3sni2AQQB/T0JVPRnR9r/iw+0A
x0acphDrc3C3rpvvbd/BDsrA6qKw4enhMyvWnSVVEA4k/sN6Ts7Rv7cRlRgdnjL+
nMdwmogziwtG+oqaOT7Re8GQ0/z06NiMT4FpAcnjibOYMEMDuRy/+5XtdJTgUCWK
tqkjHcOBmc6NYJj1tpP0BHNm2L6uv7gCsrz0Lpa8VpA13VQavU6KPnLlBw2EiACG
+txynLurKCsFoKG6weqa6mY/IZIyfsmWZsiHd/q/iSODqAeELpN/Dm5j2RN21CWY
dwn8eJvlgSO0kvUxzRcCjgFA49HCRUMo+eFyUxXWyMaaRF5TUPidMorUJVP5kY+N
PMUpP5uA7e4btx7jPm3X8oQ71oMKn900+qINV7DglaQgeiixZtciH4bLcjCuJD03
+MH9nbEruC0L3+MOMloytg==
`protect END_PROTECTED
