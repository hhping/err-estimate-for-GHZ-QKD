`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6fV/0ondgKN6fL6hHzwe8Do1tv1UbNHDUaXVQw0Oql7irHutRyNZmOIZiAzVpEt
6Bjx9da/vAQj8ZD/fdVR/PkHl3TceqL/Mfwi/5LA8ADiFIUu3YuvCpYh8no7936F
idq6jebTMx5QyI6sFRzIWjFF+lurSBX0dSx2k2KNHKVOh0X4aNMmdvZs3+M/sDYv
h2sPB/V0480BU0k+A6SAm77tk6T9K9WdRkXZGjRmQfF0Ym8fPgZppJOuIlF5yL1a
lkhRWYi3eUTglXBiD+PxEqqT1SrXA/GgW1Z20wN73+1sPkwItjAe/8wxsluWshIi
PwD3VbkjXTsF2hI982pYRUxdtVgeUpcI77m6fq7kruyOk/FtUCSibpgLdSw7Wyq7
cvfJONMUiK4p1txEa423sA==
`protect END_PROTECTED
