`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YT/nqEeX7R6TyVthj1/FmlnkDC7FLQiwLkjz3U3o2ifR6n1nlnI7g20tKGONiKmD
4LQPz0BiLLEBqWW45eZOmUHbjtVlK1jFTwcdx+IVxDx7pwp573rkm+8/xyon8pXi
oSPG5YIniW/tHqSWBMsTEFkq8sNI0eDPl0BtTkFbz+5r0wNtezJNh0A8dEXkwb7j
x+5wtblU1WvBiB/r+rm13ZPHFjtPUW8ziUMAaTfWF0OELTFl2rJsTrnNtwXDWk44
5+MXYfkH2Gl5b0M6nzit4XC5FEvupeqrqReMpKMyrfQ/cBErbnupE1LpPxSAAlhf
zVHFMAiuIunjYnkU7QrCHCuF2wcrx7luOYcLq6QhwVr26GATpnEBciQntbSlo5Wu
tNq4wrTB5mvNisJk5YCHHZstanFPoY9ztEMBj/x6Q51qZ7Jv2y1wJt6PHr+naxRW
1+CUdAKBtJ0wFBLrWHHkYaN5fzMyOvxJ/rGO1OVLkEanxHgp3mje+rVUGD44clht
8VnhGCwK/Pxygsd5UWdwIj3SQ3pO6WGI3wZc18GUnji0D0VsKfgpMx29GeHJE6tA
EQkYRePy4fHv2kETzdUr/NZor+DG46E2xP0dMCotsgmFcJqPC8l5nTihMqF9WiBK
2XChe2fhqXd73UD4eD8ws3di4k4gOxyGFmcvvYa8OfgK3Cl18ObnYr0tjbyipiRA
I/XH1qOjd7W5CWYYaMfNhU++4E+hFhjSzflxNf6xX5WFe9tZ0WXhgSNrpiiDinFd
5l6dg9JWxBJL8f0Yi1It0spNyMDu/09DVAL/HYHjfQBg7cKcyf1DXKpCcxfV3Mrw
ZSQZ9XyzejfFZrxt7xtWP0IpoZclRRXOtWvsD6/ek7wcEBFnkzNe9Zd0QvZUDqa9
Ej2JrPgRo0J3y5NbUwXJL7ofKZqALVRV/XGAEzcu5ZmuuGgdQAUKOrM1FCvVvFr1
Nz9BUn106z3GSR3U3K4Prq6lqmu9cIkyOKTVWvp88+R4XfvQCbsNT5T2RcZ5FtqD
ullVjUQGDdQUkRsNzfDFbdSUgjeXFoEFeH2ix/NFYPuP3a2yNUor+4TChuE7Gi66
436xLicBqxVY2FYs01DZWeVassveXrjSw6c4KZUMs+aQL0AbldkE4PdYpwG6ZiCq
Mv/kO2hMn+cogETAhaQaELqMpZ6zkMn9KT8R0DXzakhWPm/IW5mWCcFurYTeeB4z
97eYCbV4avUdw2d0JHTwUOOxP+pEvBbN6fftCxeiXbmcGT0Yht9TYcvLcN6xMN9Q
xwNDIVTxL1nGTu0w60F8KPeVneWtHtPWQdT0vvQ1oda8+8fh3/LopFQjvh0wV3kE
6DLB1x4ZpxFNSuHk1OBELKGwocs74HI92xlVLxHhH7o6fJfI/KhzrVeVN2+bGjTJ
4obHjW7KOdCbKSa9YdRWgkVYxPTKt+QwM7AxQ2IIq8IPml2kDQIfXEVJEoV2if/+
noqIFjaRQ52g3LOgTpAYN3k4yAwegsoYK63lgsRYHlL601hbL+AzPBuIJ+8yxV8L
mV7xbp3byOacoXCdfmjTQtnr9JYJvKmbZwW0RDoiR4uW1CCPq3hmooOeU6gJMOQJ
3MjRqIRV/FfrxIERbbqMZz0X8GtEuiei7qq/HYb0o3jdV3a0bkEYFwfwYTEsDtme
42LwadVUQZqJ20o7cXB4ClgFu7RsPQTeit6LxE2g7Lz/jdrTyg9Ze9QpZVniF81w
6aORw/ONO9cBUeuVfrtaHs3x4ZlLtLzTC64jTkmF6bkhrZ9Y7q7ARkTLrnajC4Ln
BDDA2E9rqTCoEEw4AMMZ38RMbJj7WggfHMtlqrzlhnvpLLAWeqJK2q/GqaNtq8fV
apEIXivzCfTnvM7ndf/v3zFkELlCKK9kOSyVCZnNpw4FfYnsfxdbvGObPpacbydZ
JXuLffJ9TISDmD8W3DrzHdmfyM7Ah/A+6p4ww2c4PPk0uYI1EDzeIyqpTChkYpsv
LeE3jA302ra+80ZELfwMEj4u3CWi/pV3FkFxorbK1174JF2bxRa2tK4TnUkERaTE
lszihrXivJds8+qtc9lbJyEDgl8gdvNETTs6U+ooPrM0iTplkNVVpyIT76Or4oVE
arZPRlIAq1rwc4YOfWoGGsxK7RiEsA1XwlHgtTB7+gy5STq/x2zwKLwKd6KTWNx5
+lg/OYBY4MZ1KvMCMNx+Yv2ehAmWXowzh1/4n7dGz1Qx9N99Z+jZFZeSspa0gIwk
/HfbsmzYTsrnNigP5PcFIs9HNUfgql2W8kMkpNpJxL/LGLdtM2m/25pIm5GUDtLv
Nqzc4DwPsLRwuaS6q1w4MJjnUf3XJkJigItWqFA5J4qsH6z5amaKB2HIfoMze8ga
xevAjRuni+KNJxnOjXY89EaBh5DigOto7p/NPsk4p2oXDQu4v5OXjm5SlWyNg7wM
UckhKZJNh/avKSvhaajoSXK2ficCFr1PgFb+/CQqJB1yOna7k5E/y73IGYS+B7h8
pQIIB8ZbmjTvIRfSrMTeOxr6u2LBkRaujp+3Bu7HuothMvR63oahzqe+0n9ELrPE
eR3SXtEqm0ve++f4EM5wt0Z/G+RqP1dmlSx+CjJ0OJGBHoAUmsSOodO1Fa9VB2tg
+cYqrQHnH70APIVdB91GyofJZehHbY2+j4eupJG29ZsubIqx76zbDdQunMPKHDh/
NpK2QiuW+Dcbca2wcYZHAUSDj4h8VJLEWGZT3FJRJYF+J0d7CcHqj3+xqhTqLiet
3zSetntwlSEhYT4jcKyBHaX19qix+OGD+dVv3ZMsKbZ2h/UjnofCometdI1xq4dG
WQMWuWmvAlej5lPaDThk7jLCDgbg5e2qFbXdohQuaJSDARAAh62Gh8mQX/hTiCJc
lLmSVw0/UzeGxaz6HzQ8N5fo8+l9gRnlsX4jjDkk+318v+Rbzv04qOtsSPjIDaQx
ML7bpges1i7sWX0DEuTx7zk0u3BCEftXQkGSwTreDA9yLXfEKbI4hVXUaN5ngBTG
ZXSEF86tyya5tBTVXpx3RLC9xcebEwdRpngPJSukJ+Ehe+rz86nY1njD8z404jsu
hWxfMAW4TCABm9gYuLl+p8htgmZwcy1BVzTO3HJ2CO4g2Tbc7lBLD4K53CrRlA7w
k9EG87i8bECiFKpe6o8mGHN31dQ+n6VreNzDcqG7dc+5CKFa3bO2uFLMMlpQ6Ba8
z+ZJkvOvOyV8vnL+5vWl1XUsdCQyd2yc+OL3sY2iI6wv8lgYSxrTx5oIBu/quHaN
hB53uI66THlozy1JUq8zpStNe3oaisaet5rHPa7iViOvNYQMSDzpbkymgCG0jgGA
fdxxVXUSN1fzf+gm1LVlwwJB1uOyn/M6XnqdxHuBpiw3OkKY5/5BnInRYQ9VcJC8
XB57/lmpm3V9+/eH0kT69NiD2Rn7ZacXXEJpU9ZKyXLiLOs9JOPvfLxeNA+TaHbj
FMAW1K9WQqz+WPVcWgQ2tGiCJJd08QIG+ivD/FPsvrW3hNd69wAMAf8Ewvf3RmUw
sLUrvyxT3yy3/a6bdtT2kXaQVNEKvZNGynKqzpO0b5Nj31hxOhRl8VvPL0QOwf4V
YzaqMYjIys/vDpVeQK+Xde/hCfsMAG4gvwSEuZU+ZCAJM6eNfJ+zj5sYK9r6Hqa5
ASGm8+Z6otIagatx7G/VTJr4UtY5XMMC1H2HOqnNlNfgwOG0Exe9ikdw05ypq2wN
bNFr8XeFvBd0gtJZZpRywT5llVClFImR3XcjsvRtz//Haszh3J1RVqxNv7anc7zv
DwCvPiOPysMGsuNK84jUNseCyMKiNcFJMmAt5BVbHE4ozvIXD5FervpnGvknYyky
ySbcLn1R3oaE0WgpO59OecHoIzprahTd1fC1+FOQWdriwsRLX91E1SdttD6jdweT
PX43GuX5iM5CN7IQL5mzkXUr2k7XO8w0qv2LN//xqjp2g03Rctj/od628PksWdxn
UpGQKpETJaZSPo+DXq+ahAXWjQb6ol6wYOdS9SXFZ+A90Ov6Cg3RYomB6i/e/wAW
x1LQOgHzdz4s3D/LsGW+itKsJDBqr+z6Gk+2iGmHeYvSFr6MwY8T5/Ms1VlBmNQ2
mq86mF5dVE+3Z9LlYGah3/LD4DV5ngot44QGdFjp+UB9tNslkPQU71fJIVF4Dz0Z
C4nuc38CaA1weFLEL3gkvPFrqPBZswiZZsS9e1BDXwUtyuUUBBafnXVNSUFmjQiU
sbaharrlY16KZig1ho2rejOUs81zXeBEZKvh0zv+hY+aCXDSedgXPzsTIi6XNtTH
RAow8xrOJpy4iglFMVeeURrw+cvyhhv/fku7typxARhmwRpqRPaOg76l+G1944NZ
1WkkFpPG1uG+BTP1tggITlcRpiUKBFTdiNL/iYcWUAxz2P68cFPphEqmNCQ5l/UU
P/xPvdu87OgBM4LQiDlrbXHeouvJIEs6Dj0n4bcm0T+2AgtXX8bbvX+PVl0X0XN9
l2tqG6T+MZ6zHy4PgFDXGmKO1fbZqLzAvz+tpji07v1Exi5KBXwFJJKNdbP+g4Zn
NY4nRc/yYTj6qYGenI7xYywyAQ4d2UyL3su39JsaQM4wS27KcW53yJFeeNIzUY24
ZGw94Rnvn7lzuH3/dUoFasc1dEjwJ2J5WTpIyfuI85w=
`protect END_PROTECTED
