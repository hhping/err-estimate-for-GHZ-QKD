`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MENLISfIau34qzSmJvfFfgsxsjLCnaU/eB5L9GWzjpXcEjfIBFHz1S5XlBaxsrBp
u2gdMl+CPJSMVcpPNvrmj9cNpN8judIB6PkNCaDp0BCyIFFfzlCszUYxhYI/SELe
BQAKGgKDQeiTI3IcEZPCRDBrquRrLrZJhGtnRLxzetfXXNrZ4xYrAyrQ2cICA7ry
bUpF1r7/SMqHWmKwWljAubaMrH3886jC3OmIEisF5YdcumGy+qjVz6vVznA6xRIy
RFKrRO4vbtWliL9Gfdmekz8GvWFYwwhH7P5j/XyD8Tmft5mQ7uzshFHHswQ0ICZb
+fcAAUxFNxiBHNpGh3WtOCGNpKr283HkVNFBaQEaPWbjjUkxMB+Grsn7b9+SFKnt
qqsgEveJ2WwuZ40PvcMpYyuOqXZsLyE2MRFBhEEQu9dbDt6uuzR+DxMH3uJjyaM2
Jq2U3PgX6NBB+CcQwo3KeAe0HAYZDI9oXxrnM8YHFxh2JLTLL48YziW3WCoD3qyL
8IlX337KFuS/UGUEszqt8g==
`protect END_PROTECTED
