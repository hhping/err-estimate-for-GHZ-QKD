`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFbG8X3Kl7IMSUcvKrDHMhXr2dcMvIXOHuodHDRhpiANqQ/N05v10PLKXKnm0mmB
CzSoCDSZpB2vhZv+aHgeqs3+XpUigp6bRTcVlBTB268SO5qKbnCi1kbdU3d0nwJf
7ZSImtX3QNWh/tEEkIdx76l6EHl7V6iYDjU0MvmYJnRpgga/UK5UBrNgydCoHMA1
zJWnwUBNW4zZf/g1ZsglnAMrP0kuDrMB5Zdd3Qq74rS+LBWHNKFN8pEDq2JBWQm6
7o/tmhSywvRfCZnqAh9KsQflWbd2gNwYAPkB13sUO9ZC+mNljfeV7EKkzeTVnoDH
lroGt+TrPowFrMscz9HFKM4BQ2roruVR3RWDcszewCO9+XUwPqTdl36u5xprkrIi
TFDd2miU8qfrTAsMBWPF5nbeRisPl6SjuyaD2vwaLU9cFv7RQxMSG/azFqhjimJR
Lyvl3t7P1LstmiEG6/Bs/e6cONYHMbcf90+/j1cm6uHYQqPebtZ7VpzgjCBIacPa
TSVn9QX+1zx9yE7bZCLG8L0dsV6iu0Jre8hhV5/2M01HfXIQuwDssUhmy0aUziNz
XL3QORTfGLlc2WmNpeFA7Q==
`protect END_PROTECTED
