`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRE2Pe4mzMWu2hdJEMjU8dio3XTZCDZ/5nnSPbTHmNwCCTjNVZHJG2tof55CYkQD
o3Sttj1rNPSudr2k3E6MyHoUt4kRIS97SvnsRqYgwCT7IaujgJJNWJVM38LWAHtT
+n9gnwmmG9h01kbo8Rca4a1t/VT3P3dC6rEGX4q57taHzejx/Jm1/x3xXEi6QguP
2nxCqP2aPmuFInTC/hihAXh+ElGQAQrC+6+RNIXci04VpUcWnes4RWIFdx7BZRt4
uV7knQQf33EscTejD5TkKgKmV0HENQHoyo7fuRwEPlOPPFS2bEdnJj9KePiJmIb4
P8cLO5q5hu/kvnWhqvrkeIRVSu1nvt+UMw0ArYz7R4kl0J0wUNWA1TAQr3pArPso
vNiYpVSLh9OhgQ4bv7ej40h4KAzdqGHAhT8nNEa9UGrxsrTJinDyoou6K9tG1c7d
xnQyX0FTWGI1x+rFm+V4vWwlCWaHENSFt1DOHxqMYwGbpxzB37XomWQSbQFir6l6
ilgdeDti3q8AypKYXUKxnsjCnhC0d5iViE6TxBq+ZCvE4bmxupLffgD2w6O+sXdf
zfO2/tAR2unrhLAsBACH2CojQLLmmeW3sqRPVFK2wOoURWVIxWVQLTq3FKAiKO0V
UsUt/qVEOhj4hensRkMjU3rjvrh/dbFxOBbBqyhArFdDjd5nKHKw6NImNSHVAMV2
zpvArfbR9sthxNLpYOrWOol5ANt8POijVW1IY7yPCVbrZ64vuSlSf1O/sU4SIXMD
NiaZdzSUTv+0llyiUvRpyCioSsbbLDLEPxrFHw+GRRJMvlHu+8QSUgsCcRwXZBWR
nIDK5355yZdOF4HUUsq6jVXQXn+j6ypv0qnQewhBHxRo1UgaAVTNP4roOQAL6QX+
H9UYL2ucCr609GRSszbn8U46dn5+pfAQ6dP718E4V8RUP88CTWY9ftDy9jQ2uGV8
k3vlEj6PzlNs/8IaH18cZ8F75U4OfHbiIumrBT2SzaqnVLhNMpgWNHiLf9DWNv7w
+Ap5ypJ3u20exFOLXhhaHKxTPqBzunoIMm2xBOGs2qzyb6Wwaexj/jm1H192v5GW
KAIA09NdHSwoiLP+eIMjkQS1s+sGsW4yIaSBATvMkeCmPkplegJxjyZq6jAFKvyy
ZNCyNPqPtevRPtBMYKPaJXlkAiM1h40M1AKfToPoue79FvzCZoah4Sj1bVT8mN1e
buWVhdsVzANGnZFZp3DaOWiOCbx/iS+URCgzuEsJB3zKd1hluAvO48qsDqUXkXnm
y6gOs5x+x76Jt+Eee2Cc/4TV7lx0TaU20ZTr8uDylXZapMq4rjUeQvERVNyR26Fb
wn0DNgU1o4RFEfNUMRTnleatrQ6wisr/pAE0yhAcrx9ivLFA5879FHhQntD2Nsie
eCrKYWrO4t8x1XLvTwYJaqopnmq9QzAa0QUW7L0Oc4c5huAiQWem/9RSSC+h2IzE
iYNFFm6uMMq6oF26CH8Vqw29Lh+gplflni6h0+/E4s1OmuGPIynywD2CXXp7V3os
1d3zzOx+PNoNKqTQFl60mh8Im5JWiiZif8zUaeTlWTq7HoPxN3C1OZ7HI3jrD7M0
kxBZuLu45ZCGoFk21xYgmRVpTjT/hM0y31M+YVGK+OuKevuwM+C+9Ni7+j9uGmcU
Ky5BKwUINpdYG2zNHb1EdO7M0RzoRl6ljIgKKUSQX6SumTJ+IaBkkvIzA2wGFDbl
iURmAOEr2QW6LXkcL+d1Y8MYut6RadWavrvHuu9X6qP6Oh4HEKE8fn2mniW3YW8+
6UlnUxHMwbf79MLdcIAKiaGgJG1JvYDFL7NTCfJiWrpAdCamxXoWOSjJnScX5KZt
kKGs2auvQdsWDotgJUMSbhvIwTsTHGw4GG3K91e7Tcsf2Fxv0XygGnDZltsa099w
3ay60PKxTPC4ZFYjbUrXbUmPxciMX+hwAK2BW1RmnLMI8yqR98ENfYJlMwuh0H0c
e580nYz0HgEEK2Q/eQpFlyUijEcenMU7zrww+8RM66rRYgGWnKaQr8G0JvzF6qTi
ECjGwKLcl0IU90JPISDNaJI4XcPniUuJEPZvOm2KsunZvtE0gvBTBqY+HKXffcTW
1jSbLYV2YQjm0d+hwQ8qvhU6BVITQVMTiWJzOidCWPj7fLR0A7XAt7XnjUxYUvK9
j8qgxk1zou7mFE14djKsYQk0R2Qgsr5f7zhrIkbt3oiCLSSTJlTACWDJU2g5MKRk
9T4fxIf2pcqXI6yksADNcE+fiRniuwc9j5EzLGPLit0EYHPsRIwZSLJgwWd7CBCu
LbT/T8hQW7fYLwS4HlBlLwqTCAGBBtZK3IvHCopcK7sgogZ5EAasq8q5PUKQbu41
066jxwtxVSTWm+ymBhIokjOJcdbB4MhLeDcoKovOeXh5olMTdpT98YsUVR3sZ+lR
uAonj4fhRQx+SDwY7sBAmSITBu9HNvMSEI7seBfvLd1r+3sLiNOWIXxnm3XnnLpc
0IkZKYBgiRj3e+LXA8Q+8MbzoPdyB4Fi5sSPVUoILmVxjIExglI6E22RR57PrdOV
LN5B2wsRytoVjAavnAtJVeIdFdnVHEE+00tW06QPRzX8bt6PIHqqWNlrfCKxe2ld
fRpG3oYbwUnreu8Y8ayOP5b9FqlseQ0cdFOyXZ/FlEDq2zDDf9rdGw/s/l31M1jY
DQizp4b+x0gTzSHUnoA2mDXit4/ZK3dxa4Ko5K/+jpSAh+3ViV/0d+VjjQo3Yeoq
NjUIHSjKhuqV7Ri5bbajzSdBiYk5EQatt/wq8wFC3r9c7SMxrlYtC3OZdnP67gDY
3sGGn4hV0NSVy52B8/3fv6qcD+Tt+BF9vd8HZgdKPJRJk7IPJ0ZLcjjwe17HF3DX
HgcARNV6P6dEVyoX+ukEe6Oap7VccrqIGdTfuO5sKA58NoxzQlafA/v58xulwGf2
PW7RQOD/BCBVwiYa4+yg3oIHgGKsBk6Qpm3+c8GTwbPSTQUMfwwpe559m52Z0i5z
b3Hf8VwioqgP6PIPRll/bgvzrKHmHmXS6Fm5bveUDe1+qWQPyna7tUhpLLVpW2bx
83d9UJWS2WBAylVpRg8SoDHf8Q1RWgMkCjj91wjzLDAHI+FIAIcyWqwqshd6i01d
zXdHSc5B1/E0TkppnUr6y2qiMUzaHmshdXD9WQfew8DjdbkGIOVcG63iAlzoa0mM
d38d0myd0dk0tKwQiIjBKMYTuiocx9GERTgm+GIViYin9RpJmcXv9w/3ybVe0ZcB
bwNpfO5cOJFz9MHvHhTyu0tWJuRFxtLFueVPQxlz8XvSEd/OwvN26mNzIfIG2i1p
GpgmCDECiP1q8QIetEOTNxsnCe1jLYB/T6sYW917ILk=
`protect END_PROTECTED
