`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BV2uHIGY+r5/JPryg3Jy+uIcjsbLWGnmJJj6/j93mu78k6abG0T2trtvbnrBm3yT
oXr381/sl8V902ib+Zd0u5Nk3jHgAVJ5ObMuVa42490gm6LoGhiZAFBeIZ1oUew0
JFa0ec3IOA6/Imr4czxyStg6943eSWiSbo7a0AACdEb9NLzMS1gqdR+SLMdZjfzx
5HG0Oi/sRCXzT4LXQu2XEPfqUZf59x5Z3XBG/G+b9jqbRIh+hvTQlawMywJcrVIA
WJp92lVOHPawR8GGi11EMJO6XcnSO5ZRItPJixkrTINUWj+eMj7ypoBeyAL4GotJ
HRJH4K0822VUuv92dBmHRpTHpPaDY7x5Lp0aIX8bLq+2dQmZYtctLi6APrRFq7o3
g6ntegTuIF+oQxryV9P3X3cKorctStfcCaHU8Rjv3FPkdN8va5COToIIDHcyeXk/
I1hLZa+h4OPw5vjVwSZH/g==
`protect END_PROTECTED
