`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EPsiKdqNXj0KojRKFo9U6zU1aos+/P2xikIlqf30YA1+chcAh5v96r5jSs0YdqNq
pygvIFCwTSP8rxouHa5FOpGK0kKqxQuNZVTgywly+UTLzvGL5zMp8Cr/bRPc2u6p
vGW7q+TEUl3OD0wZqkWEWq4GJ2NSj9YNoA15VOqMhGyaGSw6zPlAKtC7KLNftHH3
9YNzPveEFshk+xOklRNIeess7T2DDK81x08bfxZ4CXUnIx8dYpbgrmhWtSmF04ex
0/sAl3UFS0d6UnkN406oWWiI24SyAprc0it3fKx1TehXtgz6KAQxA77ug/nLK1Gf
qtZbB9WYjtepIGUPiFvPhjipTG7GdaLjDSqKUVmviaVDIxatiLCZz45YrpPK01+0
Ve+eQ+A8oFjseu3WwTIc5EIY7MsTzGNZlo5Dmuzptk0Uook33q/EZKPrttelhJAG
5GDehg4uHs1ZU6Ooq2/SnWandqWuCRzVMZkOkTzCIrxK6jYA1+0hkWVkb177ApHc
Cl8j2BISAOUpZqzimEQ//aD3LVKVE0NEF7X3BvC2M8UDUIbCt8nTWUH3TjfHN6It
`protect END_PROTECTED
