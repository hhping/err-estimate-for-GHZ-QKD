`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8xpg9pPXkcD13OTBJDN8PQbb8a6BEgW9KnEpzuPHK/L9hwivUtKjk3Vz/GKK1tG
9vBC4grzWXY9ijsd5rlpNhoGJpjxphDYpLAvN4hPST7WkOJ/HTbZaMbD9ZYL1ynY
Ir4/HD5vhYx5b5HPq/9TyZtgGiZLSN6or3EWjFUU7TOzrPrDb/Ps7u/NYcgadBxT
RtkpZ2/ycv/+PhQpo5GzxaBx6zgCvrB3HJszVB/cgYBrJmnqYhgiSjt22eXGc0wD
77HAXJ8J3kJsvKwP1/iM+BoHaKK4HsMd/8Qsx5kdCLw7y4Qu7m1PawLyY/SWNaod
CIL8SF7shWE8iEgp0mmz3u4n9NHB0X09z3B/QowwUex05OPi9eE5rO+Sn+Kdzieg
kUPfeKUQx5MKwG5CXlv6SOGm9T5AePYUvj0v7YJ1uZwnOHLFseltPZdUx1PWyVGA
SgrGVY9axi0r3F5LWFztg+x2g2sm6p8n0TmqMveYxznYDde2X4KQtAu9zRLl18lI
UY+ewZXQPqwh8aXvKHX1X0ch1vRwfH14jSJkxaqpFuCgHgZs3y3D/C8MhaGi/7hE
b7NhY+ZG1bwHFRUsfPtt0eTBB+CWogjs0LUbUXLNX5l1x/0ryhvrYSlvPDOxEoEy
/HOkaw6i/v6UkpXBartzlWAy93WKW5mmUdCbhcJ1pSjar/+kVRFIHoamcHyrvo4s
gX2er7Py6r8E53jU8AgD2hQX0Pyuylf1o1pwH565SmDmrUHQ/y+MnXRSyol8UaJl
zXFiWXTZHfKIDsjCeevFfAuFGkhpKD6qiWEHT9+o7vQzh7zAWrCtw6i1Y16giEsa
GLQwoWogL6mxbPxZ294P/ZLPjiflkS2pKPYSnM4LzbqRAg7An8C49+4ZCbQEF3jh
/CNR7JQkAHe04cnyE6cKsO2fVXcy9i1GzTRjbgwJSv6Hd8t23eGRY47LQz+nb/ku
3zPXWYBsYHAJNweqTxDiY4GEf58foWxXGYuXunFzYke4xrNs5Mo4b2AAaPF+wIuP
`protect END_PROTECTED
