`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kSJUvjgli8LS9TIvpUPlfpsBetKmMpZ48vpmDxJO9rnzF30VSwQNWoa3P543FSk2
U/DRVqp+DbT7oqktERaouyNfIaHKZVVTLgN3PUTPkKCwC/ExvsayfY7a91JjtiyM
aei/BL445ARwKTV/Mg4LPdLxD6iDnVWGcpXL6zj8mABVtEIZ8Db3MZLzkc5i1Obp
H9uHaCk/0XKQeberyAsngZEWw8uxaAVSJYVUuHWOS/XhUJg5oVzI8rDyly6rEsyh
JgASKinnurPXJnsmMxcBwuHumsD9D6aoTqYlYTUpmX112WAdOW2ViUBmKJYaU+FI
ZMdYjNMHidmuRonrg37omvziggsczFeFWV4MKIOOa1jwrwXxNywZTBCXIHvTessz
huYH2lxY/HX8GZawlawxVBc6Z+0zt72Y5K/wUIJfLWAYxhS/cFGKvWgpcq6wskAf
n2TmUbLdUtwzB00KsC+RRhOpa0oSXjTSCX9KKWVgt/Nc2eE0taPrQEiaFpTc3AAC
Dj1fEkhnTcSiqGcy2lbhHT2YO1rkztfPTDHFtDOyFETDwY8QiFR0s/pOEipmvY+m
5Somn+XZPurwzZs4LuKdbbWNtTX3x934c8nz/gI9nPa7zPeukdd9xAPjqY02VPJt
Ckxs4v2UTGeKXUigolOESErJqXdM37plY9NaHJO1jCb5ThzF8n8nOzS8YVZFO+i0
NSmomc4yi8aFOBSx1XjIJf/PaqEDAGM762/6sMZf3Ac5xw2G6UcTk7ouNTGyewg9
iQclyyqfniqNMDxQIbRY8w1VOGpl1C8MfvAV0V9Py6ZlXqxL6DIw2VaExW4G4RDs
n8X3hhG5ErUETd0A7MsQlaHfBbeu17iM+fAp2L6+XUmQkSKoROQL76zOipxCrXjj
5XOvXw/taZbtYtW9ayUWyHzS8Ij032JkZWDPfZg9TD0bJ/cNGFUH6GNiBT5QRNIu
KG6rL11h0qbDjgLDwJR+sP2VbfRYXXpMXZxJvOlNXJCzNmwmC6Umk7haCHeV1NkF
K+p4H3kkeq0okv2Go5/1pzGlvY+F9/MHvde7kUWbYlwKyTrcn1dDoIQpqnU52rlX
Z1fpmmjQe1Y1ihWEAkPHc0HR4e8lhjMnbvhR4/HCKFlFoN7i3jxI+bqKAm6eP2Tr
JM8obfJ/T2czT9NAYeBRGon++1bQ7EBfHW5qqvRyqszCCrOKHgTzjjZdVmXAFHhg
grQmRsm8Jhrt4RUO3CPi+Q15wJihzr8dan1klxj7rbhd4EM23pPelb/kQvAX4Nu7
NKad5OKQjM0O+iRt/nOYOnJ0dcs9e0biC8P6rViQLH3hTnJg76I8oc4AobZo8TxO
WydsaGGbjisz8ZC4qMI8/SgV4RsyiZ719m+/rrrxW/56Z6GuXPmQIRBo33fOiD4S
cp+p5CB67z/dWZSrSJ36uSQMfdjpsTsNM0IRzrpUkD+gJLvKrsg4FGB2Ax3ktBZE
QKH/iT/eV68rTQcHnYo1D02LUePlI/w3kgCZkTMMaRatfTQalHvZ/pGloAKVjEJv
cmjVEOZuMPw+aL9tbeLs9T1D97UAeIgKUVgn030BygvRYjU9ZVfOthS6t/OierT3
9yybfbhfkvgofoyqL7GhhTfVYIeO+b39izIuA40M4WsAK0PLi2K0XDGMbDY8y/IT
7R0Sa7S0Hq40UedAcQpG2cwj1HKvJxYjNq6+TyYJ81HB4ZTakauD6c+p/A4yk4fA
LLfKoVQ8EBjTHlxoid0T9ZduWKjU8Ku1fb/y9ipLjmwELggxKoCq/oNKxX8MkAjx
XWTXoTncod9GdYGzeNIi+Nds/O4TlQ7WCEBXSb5U8nXwna9QlDy2cGTvIpeDKlE+
wJ3CMuUBCW3qWrjTMVLLgA==
`protect END_PROTECTED
