`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nSp+NTcNOmivRh+Lx9gPy7K7QTP8LDAJqXvc+Ud3Vqh6C1oqHqy6hmfwrst+IXjD
OJhxjvgTqX7PcTh8pLnPbEp0e58batfEjr/2avUilb2m+NabLr/zn+5rhVpS44by
2GakiWLMTuedaGYfFTWroHcQG0ipzB2uvY3J58Nj4s2Z4zJjQ/cxCz+DmQPf7Nz8
ALbPNqh5uzfQcux377raeh08gZXyYyDUoBboaep8bSsYM7jN0BGEc/xxTLZSU3eh
5svg8/AEYL2gtEgTz55Y3dcIdKuy4Psiz3bLAZ6I/kOWYJ3AIdHV0Z3MRvj/yzoK
/+H/GJMH/RKaBDWYlJeY9FgUNKjn1HG5epzKCRcUTHmCaPWzaCqVv6/xtg06bz4+
dUyomd6r0GINRkI764InmbBh3TOcjqv4gjpr2ljB+azdNjX5JoLkrL/psueYDqM9
UKhh8jBPDOjlaJ2uGT9EitV3oHqw70jSrtXbbkPS+pc6/XnaPdhoy1uutLMElyYQ
T/U7poUQP1HOqDGPhv45F/CrxwVtU3EoBDYKGXuv6+ek//T+/au5iMgI2hPoWjdV
gBo2i0yea48beg8ns+/gEi3HkvCwE6tW/FencA+yRzSiNvNxgcIwj19+lnKLbp+w
IX4coCoYCLu9uLidy8kOmKXFpwer3Mmx5kReW+bONNjgbI/hFthv6wb7lYp+Mri4
g33rbtrK7YJFiHPCSM/PNLNOdcb+ppj1avVA4q5zyvh8hyNXLSSsy0Sv9ZpongU5
mzAM5jVm4cQmVlY5Oj1D5jwUPIqOG0v8TvRNRvGGFvth9Os7y4iAgvOi+TE6FHwB
sGdrQhiBcg+V/6ZqWqpymc4Lx6tjyiw+jR2BLJHxb7gTL/uTWBallY8mpPJrxfa0
0EBkZDXQldC7IR9AV56HUg3OAo9hXiaCxt1W1mzhi4Iau9CQqKctmwUmrcbc0JCm
mVuayb8hysWdkD/BOm1QHqE1weyQJ1v1cRvi0gbIhX0++9jpJiZD3KCipx+MZ2dh
rJU9ifjI4LoUaoLFMJumEk9QpjAIugexRrPvbMi+96Y=
`protect END_PROTECTED
