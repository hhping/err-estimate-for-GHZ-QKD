`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gT2YWFLosw1A3epG3vA7nOhxu0dOwb18tAjDyU4VYJeU/+ub7mU2avOD2F9JfxbW
XnbGm2Qmgs6EUSHdZJOUoB/sXQ04TU1pZrVxECx4jLkhhpEk3JOqzfmDwRddw/eW
hEfrmMKDRahXf7hjVNIvzueE/ejkN6OKOJHI3mYtIIGiAywI+IE6cgRIahnq26UJ
jaGd89bdZF8g4HWFcwRZoheeGHsOyQSvVpCV0jwvnSJwR+sUcCqz/E63APAjok2T
UTlfYdXBsX2inRpgCnWGoRlWwqIke4ZYMp/2qBUgyBw=
`protect END_PROTECTED
