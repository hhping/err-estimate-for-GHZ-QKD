`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rEBe7FqZuTer+wzpa0vN4kNL3UfrSFVZfnTbdgtEVX2MCmI+EYu2Z9iyfvEtnCfL
V5MWS+87uX7YvsJslNxl/rdebo4LUNu2djt3gwzvaZn0sU1Qn218hiO99OKSLuK9
Pg+UTYRbGEsRqLdRETBohhsQbvd95qmwecns1m4MNMbcrr1CauCcdGfeQ3hlyR4G
72FOqMVyF8A92nI+EklAOMNVv/0sRsja/ZvRP59OWyUD9zPMRbf/FVukQfaTsFDi
0FBoLBCSImwjfIYrVTDTVRtMLB5TtGUu4g10chNk4AGrvu/L6uwQ2g1ipwQMriQy
eeCxpIKVqPviqgnfmf1/8J6kVjOZEa5dWfyoKWl4p1XzB1E/pl9l3hrmLLc1/EUr
ynhhvgBc3PQWCBqvaRVTxzQDop7M1qj07KGeBsVx2gjQ2H3WoOeQ0VYPruDph36a
ZqzkG+6k1l0qULX0NQZPKA==
`protect END_PROTECTED
