`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eM+lc+UQcJ4lJRCYT88WbGAvBaJgylb8KH2XRQQ4l/y1iRqAweydfoDIzf1KeNpO
MGVF262GRPkBBNNhJUvGrw1FbOfFY5vi4rd76PTRT2wVIHV1zdk+8ImdH/rmCo9x
kYJToYdMmscF4SU7ye8h342GyC6QK2bSKDeBCZviSCvgYmPBwUiQFmjWEiVII9+9
q48FpWCixlGO4KrZ7qjgpuI6cYxQ9e4n48R7qB9ToMumCNMHQYL0/UT6ZLZy2BVe
vGInmOGejRWX+PEv0+qO6QIF5SIUXlbf9ZTwGhz8nHADNJW0RvgZn7ubub7JrRYy
+LpMTTf2jWUN8mTiD1spahnUjwVBBeQs4pOiT0g1zCiNCB1iSQrnGPwttIYE83py
rMYjKVwDVhuujhIcwGiLX5WWo/3PbZkh2nCQ4DBOnS6/c0yWmcW4aPDWsfB2x6pU
Bu7w+O3p4nINJvfA4m65tM062uj2p3elwC9Yx3LS9rblXxA6WQ5tV3IG2nS+FLou
6XT1hFsejz1uEIPi1sq1qEoKgyWkg8kge7hXk9qXNnDhvgwGZBzOgBs+BopNNPFO
045UMij3/nZ7Mo+rtuIgJe1aPdPuej6N7ZypRHId+vr7CXNxbzW9980Gy15xmyWG
1jrEz7036lKqFMHbmlU2q+DVeqmPM0+g86W52jcDai0cB4ZXnfDLSTxti9afIdQq
4qKbpQl4ht++JJ5A2CntNXbQoqw/6G8I+sWpo+yby5sWQsxfC/jSK8qsyc7xKXRH
goN9k3lp/E7NGsOQQtcbhQDx9GYno9YPVdZHtI8Y/daSfQp0SNC6R6/8YFU3XhAp
nVDmIlpHvLY6ndwUVaelOLN7IwehmXqhZShT8iJIdW5bR709cMgnBYJk2ig9nVFV
PSVzn6afiJVGcWkbbCUlPKUW/PZzKJRFuIVeVAuZ/vv3KQ3aNP43GgSu+yStI/Ho
K2AAjWRSAv4JjnvODKHBtVyc1iL3GvV8KbbL6/l5csh9k86z35ajF0qqS7pT7Xob
G73QCMnM5iV2uvV6LSCXTbQLnxaGJEAF5+21/2T9GlNiuZDOHIUoKrzhnCG9N91R
AA4Quf5n+2O7ZTAHRcFS+Au3M7iMXPXE+DZH9KvAqUE9pEP16s6kVI9Kf0EtPKEg
ozfIxTkpT1x2cFbjwjMVz2FJF4GLG5K0QSrPDDc++Qjdo5xzRjC/6S0OP6Lz4DB1
lfXhcc9AexM0JB86evfZTB4g7wUD6Cdes+PlOuqqF5pGAf8cUvdXB376RRWMiXta
y1Exe37M4BxPD3So8SCMivdrwbEzseF/wq+XN4Wokh3XDBp10PqWYKLVYD17K9zy
sIcVbB7fCEeLTCZDLWCxXTYNuhvlj4fFXFGwZyksNCE5bdKraEBK4KOmguW3DqaK
CXP4SLH+FptjRki0hY0fJQaZ1sp9Aty42wx3PkuG6Zh/srvf2a99WS8A+fKMZKIr
x22k8rpYEvqcK07CmQm4zQ0Gfqm4hXWahig9XHqsDE88Bl7RVugeYtRofBPxaBeN
Ur4EAlidyjCwrifuYxPQnJvMzmzNmapvxeukbZV7cS/Vpum2AzEIXwzKMZb9m0W8
gm1wpg66nKQobrzVx8cA7KLyqd1plCTGUiAAvWx1EF+0klzK0Nl2W8LGStKiWUC0
We8vkNeGLwAIAtfFLdTSVVh4JMRN/ZpbHBcIN8eJLGEVABxZRQz8SVq+k/LquuQC
c8xfPypeNg9n89cTVt7gLJXnQMcOITKqW2QKUeQ4zei0ce4fiaGQdAmk3OLVhshT
`protect END_PROTECTED
