`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwM1w1h+Qa/x7KrBu5gbbACifk+cuTIXYYwgc75gA8FfgFfatyQuVAWphq77K77R
i7oeyVB2JIzxf8rMX+V2W2QVy4NMBN7uYQ70IpiCytCCMWwzpVjYtPnUH/tyA6Ia
zm0fx+uuK2ZZFSpgQuIFBGYEutebvC8Z1HZRU16k5ZxaDPQtMM/VcQqo3ZHZSzQr
TgTAqUvcBSMk06PBXvm+8VrcLznkCYqMdnk4tN5L3tgP0l2zNbnS4HW5rcw2kWog
133JWn/nzLJUqUmby9bGz8P95p4I/9oCbX8yNmZl04iZyuRvZB/UUlnYs2E68ONd
WyJswf1m8b7mLmlce6QbCW9Aq/ZV/XL36y9poue9a2ED6b7nFbR2S3gbx00OmXig
zsIOLtwZzPorRFCPKk/bUhTjeR6zudMiELVPa7LRPEQmXN3PqkzV3T28StF4wshu
SD18CTbZz6qNH4J7IrkQWYTwkFa5+foy3FFWD0sjzN1/mk3zYNYUJx0ACgBigAr/
RuFGxl1MmXabT5CLKdcDx/gtV5fJJkVr5FQhjIqinBWHOv4KxxtraNwJ7H2U8ow/
4RM0mlYT5GQUmIGSUR4rDUfXJjEWun2U4MV2jicRqNTY8yDaWYWMRMmVIWfj78hz
bVQfxlMfcpO2qqy79BbcNHT0Eg0iypWL/zcqUTTCbhJ1MoRy1iW0A2n7/pIzBqgr
PNLtLEDRIfkUMkYCbJxQ3jyOrpKH25f/zdCshK0IWLEj/fDLWRz9gkIkheWgv5JO
X2GONKJ5twbXqDgJnxO9p1EKUfMJVds/y6krJYZRUgvtfX40hujh0145VfRuKSY3
BbxCSrnijYwOGVodEqYMwBVH09ifHUwA3wF19UGxUMcJDmFlQKbVrEZp/9bs95G9
v3XbN9kpsz4BT4xmdvC5UDCXn6SRW73U6dNjiDAUlyvUfBIATr0+gHvW5fuv8Cs+
p0BX38urH6BLfJVbDYHuTJfQJNb2vnh7C9sPuczABsAHbT3EnvJDXzCyShYcrgHa
CLA2VTZYonPF6M/cfaC4jOd1lCRLx1uv43TlPn0IZvYih+7G5ItXPTpQsLxNiZ6v
XAD+984l2GYVJdJfxSCroOIYNh1j85YCD5phHpYsv824l5bOMnV0yGqwZL0y+tuJ
yfFIemhXXnFtaObEx8Zt80A6gHy7/VuUjNs+asIo5m422h1bpPBvC5efoTBVQ4Eu
lSG1xXJKYVbTiZ0vSVFC/EHRtQ1auQtH71+7ytbKRWeM5+WZrHfY9SZnfdYJsnFS
n//cvUDfaV6w8qNeP74ISfm/tqnrI5gZEB2367MEf8oEQjkMosKlCXY0OuicuRUH
6rDwTGJzIuTPXSjPF2a0RL8mTag7ANRSHIGJ7zSrm0WNbzlnF4LhxPdX6i95INOq
G3Awpm4oKUQBL9ukoy4NC+kRBoe2Oa73zF28aO0El5Sqqlg9IMkTkE8Vewc3p0tk
OfT54OwYtIgMo/JmUW4H8pJOdsK48UXFt2Zh3VLnSVYl2M+RyskGvfw6WmKMek8M
8PJKy37gssozcpoZIuD2UgkJaltyOOaZHrL1MEMc8zbe+mqZhPt7DXWsLXl6wQ3z
TWgNmqSBTZ4BllyW1r+hZzhPU53K7358b3w/gYF8u/AWv6D8xuJ0vQ2BQkIvX7Fp
5myXXlLUFlAkA/0XyUDkpSHq8EdyAQW5YERpKWMCRotkhlX8aH66y/LRCZDSpMCv
qn38raUvmQvAwGSGxmYXKYaitwjOoCSsR+iDTWajjYoRXd4hK0YCFzsXEcJ4ybbi
x8qJmCQXoFHLS5un0KDszlyPaESXqPHTc6/JfMqP7qWrKfQ6268+iq98clZa/bp6
4Zj9gXtPdleoT+BlOuKQ/+AqAZbjwPimJthTlvS8L4+QER0Ss2keOapp3GdbzTdI
L68tR44P6OarRlUNLxEtueec+ZA28pXoikqk/aJEWbGbaFyySTbBxcdhpHfS+Idj
nFoKfaWse2QlTAG0XeGCAA==
`protect END_PROTECTED
