`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
No3YcQlrNBk6jF0+M+1o87tk88lLIYja4M1HD3g9DUFVuX51piVDYuoHC958V/9J
XG9yAdceYRFEhMP5Agt5vsY5+An/CpYVHAYLxqJ67LnVQpU4qLUC4kxbbN7THE6l
RdPbfKERCrttOKK94L4apqAtFQHT2AZXeivU+rHBvrIZJ+Q4fRPlpRSVI+RCgha9
I4vSKfzD3QJ3je5NC93Rq2Mu0KNLfbz5g9gEu04XJmQyaeGm8SQXzY2535xyM2o5
THSQcOaI2fu1+1/DE+O8IJ8sKCUEm7+hUzFDfd6W+ms9//pHgBVH2El9Myz35mwG
v4jpVEEl+g6e3egmY6El9c1PN8Kkt+iMjcGly4aNeVk+DyeS52775Z5Urk7FUOIJ
y1AktHTX4j+T7IgKR6fmI+dBqXSgZOtCTsMeEwfuf+FlGXviEGc7AS20Q1XpLvxd
W6o8QHHCZGmrKKNkWd8jjXTEehfoLktpg9zEaogRRz30xFUUfb+soTei4OE/JoRV
wtUm098K/B6X8EOCKcU71rFJd838rmm7PZNy2LNs8deiqz8gZ9q1unxOzf8E7oxz
w4NPL35m4nFdJCEwAkHMXkdm99i83NoA68dpDKaO1cduEO7r/Ok8qtlXk4zD6lon
T3iZtBQe/qUCM4JIHCXVZC2+47+ybPH/T3TRt59kwiEE6o21W9xmPtJ/EpIj1D9p
pwdydcFpbkZZO8bK/rEPBYNT28Kj8AhiBGKUFrpd1sOCB7cZNgD0ndqqqGAOfI5m
fThRFtNNLH41e2RxljboRPnH0TlUhQr2qfI1UW3GbU/h5NEwyyWoJ6viYDiLPKk4
thwWckD+Un1ZLWf9GWEOjxaTb34rr51rkxMeXlhDSPzHXJEIA8REJ4RGlrTBsTVa
5j+z7ph2vlnn9X2yVNkGzeBeEDDnXFzJ40NXfirv96icxwge0SS97fSoWTtNoUiG
wGDZA8TMFsCXwEREjU7RdpTukGRq3yi7PGuQgGPgljwZ5CX3Wglq6KyKaShI03Lj
2ZQAc4RVThNk13dN/noj1cEe8P3x48nD+tgx4vznWcvtbVbuT4Ae5Tf7C00JewMD
Mv4FsbTZCQ0cyIHM+CPUkwqDVNu8e6FduNHA6GZXOoWekncAAGQuxsjgXMq1/Hhe
tjJMLyfKsJinuUGONcZseS1Gs7P7xWXtsdp7nSm4LbRT2rC3/Hn46pxU9ZJSjExx
UfnoqFpRMraT2Ne94K9KwZStO6J8DL6C3oX93gfonJxawfOwLiKJ5PpBtOQ87MSL
Uuke47FzXC7wEzXGpredUn4XUw52pGsAIbdHlrbHjA2RLHLwDpxQOtbpcfQ8aw7o
oW81ifF4b1tZInxvhc7r6mtiGjiaqdln2M+i88AeW2I36Q0db/SJIpXbTyuKqJDC
Ref/v7JJscurmxcBnqHSDyMG4s9lT5cZlurLjj8YMucN1GTZixkUakVAka49TuYs
w+cWOjZSoQzj6MJRWUxSw3HJE5SALR21X+YHNHd2+E6hfPHS3yQ2d16O7idvYkL7
MDZ82JnEmRTPC7B+OGDUi0qTAqDkBvLFYI9x7zetThynK+wu9i54LTYdcc2QvRK8
DV7m3MY47YAG1nsfoZHmXzPCi2REeqIeUc7y75HVxmVEHPblTFJtQatElaPzwlwD
Zn7rk+S81Q6Du2O5Mrz274W6+pqWgmrMkBmJjk6cWbUmdczfdv6r3kYbn9KkqgTC
owLJlUSJhMCFiqFF5fWZohHma5Dppkg4/+bQn8wDBnx/5eAB9i0VcxVCfvFN6zAU
0TB215+ua8tkjn/aYmS1A9jD15URFjHomGvu+pbd0oV3joOgsPMxQ3c7eIUuGkxd
GEkJ3gJKtTOIqSAMF3KpSutznSkjWrSeXk8YU3YIsFoM9BelUljlnVVj1+MAcDhQ
y3feie3b2AzJvrTZex2VmIMW3cxti4lMb23+gsjamrJii8zlcLGoi7qXSYaQg+59
ogpajIHq80y6bykvQsy+VdGXDymOWoQlin3tt5YfLFgesaPr3Kc1cdFAIdu0ivpw
wPpzNxSbE3BQYSfqbZBVNAtgs9vkvtYMNa74Fry8OeLfLFCHAbGIl/G6eT1QntRO
mMFYlvr2eEhW07MMzATtepJIKouE22Y4DHxXpxhVjwG8lMgmqjE5fqq/ujPnUeGA
mFgrTrD8DcpoAwfZJ89LlUoCoLM1qZ8z0OZ+jqG4PIJoB9rx+tjGoByvKYmOis4U
hdaSS7uPo+8aPrdeNlyoqAv3LeA7+oQgfgN/e+nCGW0AVvLF+6HEh5erZFryVf7w
eCgXlSkgBL86Yu85MyF13JY8629eirPlrJU72UV4Fd6o2PE1U38n880rXWCnHFoE
81kzC0XOITifK6jLkRIAU0mtIBUkSCVto2eMZvNA+fwzi2JcPFrMX6Y6OM4B4x27
vIRK19ygWh6cC0hyZJ3E2jLv4FBToYnOhrouDwHbr+fBapbwNi+ZoEywR4CaTrCM
G98bM/ZbzDqvuw0q4pU6Fecf0LYTWGY6QfL9l8Pvd/8YTD/5GklO1t22HSPBbmWo
egjrutX2P9j5kMKVKg3ZWL2U9g8ZhEZkQbFXI9YqjI5xCYG0qi8Xn4Xoz/6hueQx
+yqd8JKgVCwwMKcn38CaAJqehE49EnTLOx2hjVyWEgg9d7LPTyu6ykpqZ9H4az1Q
Obr0CiCZ7MY+Q5DFoMYPXT0uMVyrfA1YZX6WoZ8Ps7hUhV3AHH4a8wUaB9fEidpW
dMzu9EQyrm8wdtWcS1WUxXwbbaZOOkj8II/es+/99BtuRGZuNha/3Rk4UulZSHxw
9CToktnStBkUD3GVWgdVh0RKMz54231JEWgXEYOnPWoPBWzw7v+c/ADDi5W9ylWA
btllCW1tv1pfHP1HWR963tbENPZ26ExCBsC7JyJ2Vp6AFTZE0xYfipPxw2uIu0Uj
h2olfvIG9fjBtVQy7qDp9+iOnVPF+vvBRjd0N0OenGPibEEIOKNgVffoIeVxgmA+
RgbUKqeB2sQaUR8Ioo8O9kdKsq1YRncsXJ95wOQYONDMbnfjTzM4ssENBz+ZwRjd
dy/eH6RNR2SL+cYzjw/zZtfefwPCsCz9hOIVMYJNdvocHr1C8VLfc7rgk6YYchyC
V35OwzOsHJJ616UieVaeIuNDA44Mut9lCCHXlLbfkyPYc027sHosBfT1nnFQJZpV
cr7psmrAcwO40aHk0nI8VbQ6NWxaDCZq/WgYwW0j1yiIIJhBXSvWPFMVo4oP0hL1
kfMmDjSROhwPHAxqnkTXJEsaNM3BYEG4ACjP0eLSk0nBDud6QI45hEg2d5xi0SqZ
uHpQtL65hzsyfMd4IJv5FoFlmvAJk9xy5qRaWok6X03VCATFFrKk7X7FvryS0jwf
WFXS+z3AhihSogKhDGU+zgaDVDgTgrgs1pPk15ZLaoe6WCFkugeXgD2P1j8RnZ6Q
0kY8/FAUI1iBr8Ca4DEvK+c2pbjEvV8cLhuiKl8sYYdZYrfaQadLgLDiUsPBTRFx
qeMLzuE3/mL3i/zbAJWw9A7NMl0WimIPMLQ7xet31M5D7PBK/ByM3aMaWLWWZfxl
muFYA/dchV22Zac0uI0179wY2jo5VgVtOp+ny/mdwzVeR7ag3nZhv22PnTD/6r63
6Itq4GC/ivrrimrdyPF0dW5I6aXjVOIDY6KsZEigS3YxB8TnAwLxtFgOhg/hkARJ
2VN53/vn+Tb7ovnmGnLMcNiFQVvp6VJ5MLATl7Xfx9RzothRvsj2vlCB7dXZfLkf
XU8ppUiy6sM84wf91A3qgCzvMP1rYBG3KNVyW3ow0YLLZ+ho/nDdUNw2Kfnf85Mr
6EXxoWq63G2iuo0h4Ottw0/I86NlXpa6ae86U9VlK0i0H9zdm6fYrxOrwj5kKWr7
5PIy7KDC7Lxr0sIntbBc9B6wEXDZWX9wqSgSM90BpmAArJMc28IuQdU+/xakG9BP
q1hrmWVwKSc0m9XOcXFbSju/GYm7jsDiICMxrH2jigY5JN/QGxrjk9himh15f0Ro
HuFTnC9MXPWT3f7mE1/64v/6nPPxyQqdEfHTVI/gQHXq1llpa2749TLLhuK1zwGR
Mf5RxruUTdrhQBMn4hcE8ZXY/5BnkQUyHs4cuoxEsmk=
`protect END_PROTECTED
