`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PMdvGv8DnQsQhgoQ2I0rljKgsqPHiom8rLdFPHKDiq+Lr+mtN+wJvJrtQWa2luEc
6+kJDQkEWBUvM3FPXsxn9ue1+ataFCnem9+5niCXj4mIXHz0o5/TWnt1a9mv9p1r
NxIGQuu2XSHSFxXs0G20O7lulzw2XfSUe3xSzFXF/ODbWL2Fr58457V4Cb63NokF
ETpeucIJ2c7ZOlEtt0cG/S5RO8nDYKazA/IwxUW83Pqk1q0S+Ro71pgwpYHzvusw
xCLVtQvxPsraOqWL9XuBoN8Mn7gMwue4YUufAYXfZbEn8pmYIDzF19GEg2xEczWM
o/GbWBQsDhXmTYJW7hMtNtZccIjW7ughz+eYHnroa9e3GoTUcOHNp0rw6KYeEsNe
Yr6Gvk7YFOKQiO1ph+mZhoXfCb5WYYUDsY996vHUbsDXExK2121SLfjgAVs+37Hj
LYXVUv7L74Hj/n4mpmWZextJSZaA/a0HYsBRaN4RVgjvR4v+fJwJZr1OA7J4Scjv
K/FME+TyFptab9eqsny6ILjkM5S8loX/6HT3c/2JbR1OfCq9EHYEMul16y2MN/TM
LXySoaBzLGNzs8BMaoBoO+yMDXlLYOaFmJpQcO23ashtfMozGJk5rNaoeY2oUQWr
I9oET/zuMGgCEC/yH1UWzRaOuG31av12Dnxx+Q+Le2jVZT5hWpJJ/faTm3EPlTpr
wB2X8g5a8sRVuhcgdnsE1nYp+4kfNKySz2woCrBI9UZogS0uh2YwmFWzGmmys8f4
iWVZEWOteyJOAa0uZC2X2zS/yuHkrG8Qpp7jbVKe+B/ySVPi8y8sY45+hmgBYRt9
MGG8vSsegzdv7vxfuNJKqVy73f8WyCliuf7gAk9mj4+rI4FO2KPks00UUKf+M779
L4p4zMSlllNGotTPbau4Kqu6FA/UvNVfYeYOougYhWfNul8f5+NjRdYGBrtoAa+s
qa6wmJlmId1RXfszOudoKQoyDH7AHHVs0/yC0M79h0R7Y0okBSq8VFc3Lsp38ayG
QBgzvSPFzJHaaNhZBYj4tg==
`protect END_PROTECTED
