`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ABVhBHVvTQbg2mC9bh9fGZQiev2Pb71rJV4MBY1AT4Wy1wnguPoc2ZFA8knqOKb
TI1seH7Gf+dc6FSUege7AzCK19MUPKqgXqghUKnODXMWGFWglHA9z/bmcbNNFJjZ
nT7GaaQ2seATVcyXNJpHG+AMekflH8+xNZwmBQ1516cJbnHJU5ygFnfsj2THwoJ4
YYs9oO+AsEsxt9lZPkNqodQwUQcccOgc5XIOLYuSOhsjUeEc+Ej+xl+WmtaQ3KQA
NHl8F+QlVQgOq8YTURSoFoXjRyAX+qQOR6tVKw4FZUYIpsX/AsWXiHGVLrcXtOKA
tvKKSASNBZUdiJ8/K9tXOzZ5t5NC+wr3UiGcyixtWZdIroNba+C5lQ1wH4jiBWry
BaNhD636+ZBo/PzgMHo+GoogkDy44hC0HRRP6o1uXaJeA9ptnMkBknk3LNxTlmNV
/rArXxpnNi1j0LSk9QLv4HcOvCUBO6chSksNp22GNvuZEZmS8vwewKI+Ia005qwM
dYmfqQ/YmmcAh4X6F5AT2tS4uWm7xdSVDf6z9FTjKYMRAbAo/Tmky+6sk5dmlekL
svyClYALnEnlq26uKTnw1GmT2kByYk0d7FejnXcZ9iZIUq2dGSfuG3IT475N+pOR
wJhY08qrGf+rmDRrsHaQMQxgl4dbk2J359GLSu53BwwvKfQrZwpMPTy2SbF67aLB
c1gYIqKKSnMKm2OHGD8R0vH0l2T6dbKxI0ByxvPzNV7b5gOZutqnvbgjrR8k72Hh
Cs2V+5R+a0gVBOD4r8c7A0GYeDl9h44wIpmTJSZn2K5ioBKuzor3CDrUpSjdOEJv
0mC98eg5G6gue+/Fnwei3bsogUlO6bGCZrTguQduKN5J0j5bL8ynlca5jIqNiLbq
dSrFD8EOwPOpqi+3Q5Ye6zjMSEbcZGWx3nfc3zMGScLToks8yK9Zv2Fn9QjVbWjA
B3qNWtsruSu7nxQl9V6hroCwE4YVJIidqw+z1gUw5pJmcN+Cv0ERqHak9Cq4w911
q5dmQq1s2/INTvUn/Qe2M+b8ptJZVLNLwBp4D15w9jSdhvKBOa7CUMq45m7F9Dyl
0xvfKM+IESl8FUznVOEIpbtWrZPtnzmR7uJ+MXFBsHCoFyesTGxQZQKEHX1dLBoq
521MRl1RWLE3MMGi8YqcDXsa9tVK8o//0967UhFcyoVojELRhYSOZDaIcwLJEQqv
KRjcHtUB01vQ8GTfqOVjzNbnof3lmZQr/Jud+d7ARQOCzHA2SBPIy8VzGV++cajE
MNTudFDNj+C1Jv3WyGBC5md+04HpS53QW2f/IF8zAHViQ2pMDGffmxgtEZR/S8Ou
EH/dpyN/wet3SMB5jSOhAiSZXPFy/MfqcFGHlDJe9uKRUOAW73f08r5cahpgmx9m
EdlOQ/EX+jr60EE9fnIIcSUgrCxFKWNRnci8JH+m1JU9jN/B/Vq04grKyZc6ZPW1
IsP0Ph+wz39PYoOIA/U5Oc8rusFwM1i0D4vbgmxykEY=
`protect END_PROTECTED
