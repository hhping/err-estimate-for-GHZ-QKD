`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SW1VOwuVZ5v0cH6bXXBbsKkecG5xo8RNTsYY+/hAmjBPHOIdhYhdqrkEjPCjMMXw
4HIaB4w3k4xOm5/mCpCxXBibd7vQl2Lhm5khF/HiqSXA04xNzrNEKnImbEG+fO6P
+CKxVrkCNGnrWJNlrf2/WK8MzaiWnwYB0s6jWR/TBPsi1ZpVApTYxqkhK423Y43a
2r3wOaw/nzJCVQVU7BjjjM6Jxj0T0on9hzVdL19N/ZcG2OvAigCGol+ITJt5z7NA
nWJOUDxrRdMpE8lG0GPBg+7s+AppzaRcueYwVdmnHL0yIZy6jEhavy0xzVNXPpZ6
9nke9PHSV1aZ4zMlZeiL9GAb/8vTyIuGs1nBKNfYLpjGqRewu6aIEVaJmdAMVPxl
PXYi6zGOXjTpG6PzYGcUHXlvWs6tABWQyYEnLLNRYZXOx1n6qWVO4WzriKL42y0D
G7YuYdkhxA2dsC+wsZ5+VZer4HbQchnz1+vmGOrOQvSsVb5Yjx8oH2VEcQlKsft8
NmssJXUlxm/kpNRyLwPQY4RVXEjOgl1DpuzvbMhQF05cgSduPUIUIJs5z9Urdh55
TX67f/V0r7KDsRu1Go0E8RpX05rx/jhvMOI5A9AFwrYRXfpUwGo2M56MrVlPDR+/
UqrT0oIUeP4MPDVk/VHTAzb1b9vw+vhHrmcE7QRGojGnj5iMCzmHNC+626d7mnX3
KKDuKsNmZWpfo6xNOdQ3flVqk3GajT/Qzwq++X+pblDYxQmls1lSTH/fBwGWM0kL
5fKxucalQjUgomiAgDPL4Q==
`protect END_PROTECTED
