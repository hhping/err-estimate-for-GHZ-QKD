`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+URcdcVfUEi7mJVRTQd8D2do0K5CnWRe2M3uQwejAoFr9BXdf0oMyhLhpFNC7IC
EfZ4zbp3Fh/HEwLWVGOmqJ+Kyq9+aUg6VdiEpg1YTiRgp1EKjfnbMsEWOS4i4QBV
komJHBSPBkx/yfbenqhnxj/yV+nIH60rh5JOgMTkqRPpJn8TBUpRi5e4T4nkVWNb
mjalK4WECB5sE0F+73F4iqrub0vthHzdwJwNia7sgfl6k4s2TY+Z2lUXvnvBnkJ+
hMrWSlznv18Y5Bmj2Vc1i7O2sfiXHrcasWyX3m+83IQxXzvH7RFdDwVrUOgLjtRL
ygOMyO9cW1jCZMdwWHUg61iyCSCHtallaqwJd/TpjmiBIYIdfb1Zd0b7D1S4uIHt
3cI09pRXd21LqRYtAvQ7so99sngQQWMK4oh9lZcl9I2e3bxhyln46fPCmQTYybtO
15FHijPvl/FhzDpZRdsrbYUYDW/5bjeaA0vv/edkZfjtjiX/hHHzSghlfyiCVfz0
+L+BEYXIhZ6Aw6Tvr9C3RT3OLuUj6LTPMPt6hk1XXu7BosBnV4wBqwdIRUxvZvRs
u7PzAQlLZSke4LJ2HCzqEJSapofCcGDCEDVt41igUdSrdRAHMuHlkF4DwbFzu6bf
O3hjck5ap1T46Md1PBwymEod06fLRKuCRRASAo6Z2jj/rEBH+7nJX71oZvhkqgM1
pc1Y3UsGJ091D82pyBd5ikXA9vKV/BgPLdh1Qae64AdfsEgT3UM8ifTSFPtKSlZK
W4yFrnUbEfZMRnOAa9GjLYJgQafsrPKhW+RIQK9DxeBU30QACk654VR+3GhWJexO
HBVrdriNa49w9pWd9E0VY3h3tnMSvrDVosFdUYD5YO6+XbnxqkWZIr4EHSYfltdg
cqpey9cBQEIfBCBgQ6csCQ==
`protect END_PROTECTED
