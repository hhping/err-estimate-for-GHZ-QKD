`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHF+FD8ZJkv06V6pnb0g6P5KGwdeqKPmF+6pUjHMXvdbYGURWXPi5IjcAR01I9fn
B3GVchBdl8DpbEgBUIoCnTMiXjv3N+P9j6fM7DARSmwfxg/4BjM/4NVsdhQZnHWC
jwiNC+oeC4kn2aWnQ+ZEO2AlUzcUdcpVIh1/LdeGw68a7J76EiF8rCULtrQKSTVJ
ISeTQd/APe3+wZi/5/ZZgV3LXGX9LpmcJ+8/C0kyVOdqvLw7AhJUu7hLKFaWA1sn
JuuJBZaNn8JqyhZ2sah6ma9WDTB3bPNkfUIlR9Db3Usv48aWdAZFNqBqiHCgtdcj
RgDWqmnpnlQA2EN5CX2zfZz8W4ggNjDbJ8Dg1alLosh6QutF81HqzS6xTTZ66SCG
+sSe/8gxWOwYGIud6v3cgINCGNYYR4RShG732MzGRDrMOlsmww1qXWBeKNaBxiBD
rSJb+JEs1SHnPTeZXyw3Wsi9X+/YvT8Anp2X6T2Quk2i4qoN+guaiPFQJNUGpokY
x6PwkKkhuBy+4gXZ/EqVq2Jtrp5gC4Q48KyGtn20PGja8o2KJhk3L8r+Xv1E1GF1
aS6DeR2E92viMJTwG3j7KKVMpiavnr4uipMGvTYcNWlz43/uQHt7ksU9/HvzshgE
T1hrOiPPdw5F39fd+EiewzE2CIMKbrA3Cy9mR3VHzXTAP5nJJ0ZC/V1NOu4DqX2v
405Un7vXxJlzlxMkkZQ3xRURk7zHJrpoMp6iZd3heOjyJwzKEhrM+uhPGYs84xW9
AuUg6auhXqW6dwHTtM9qiCGW9vzSpEZOI68EjGKPfnMxJ9Ad+fWT3jCtnX8V4Lct
9E5yDYV/Y2493Oad/Johx2IMFk+6u3njLFePBKZAIRMzTRz9AE8JjM3GZ2sCXXB2
WmLPQYSIHfSj83Q1vM0E/KV7/Wt0MxIWrE5yr5YfQykIjO96e2TUkCaUC7FDloUg
rUg2V7KeTl/WNZklYlTOQV3/N2f1xq0mFjwkybGxJZQLVk/exJsMLfsw3EGi9lqX
I+MHAX6fHC0qGTBiABFjBF8ks+lDEk0hfXJmeJzZaKfIsV/BtEP1F7IIVvVgcbF5
9dBTausUaEn1OHWMHwfno8kAnfMYpV0QuCXQF++Arb8bPbuVfrq63442eRPYMqZJ
BOErLvRBqDbaBGmThZEkjT1qoJcFVZROGwhSLgZ2X1m8S9OzEys91MjMVsPP7l/j
ewFqQQlJxzrsD7VotrZv5NKs5TSKwD4o8sx1g0/cqzMLUcqKyEIsqwE8VUgwbAEq
iIm8wZyGD1tkXq4SAHwvJ4KO+YZn6KGvPwe6sSdh0vw1ZVvuMcoe4aTAZJtYxJF2
Cggm0Y0THaoswEBJHKhJnq4hL/G3FVc/Cz3wP+fWvxO4VKDnIXPBHxUD/PFD53O2
HeIpZpsz3wp68djjPx1F/KSYzlihLMZocudXZCsTxn3O2vSJ3X3GjIRYL4/QAYcz
Au46rMzC5skTZW3PW8JkDUqb1Ku376mLjzhD7fAyRu/zUb8EstlzdctDmCfr3fal
V2IauhD5EcH4c/exr8nIrjBc1Ppz6H4YFdOT0Y1hZdYxkNdgKz3D2D4BEpmlk0H/
IozYGgjWLjsbPPouNR4ERUXfe/BLp28kRVqF5VwjothmbsG15RaPJlH6NIWAJ0pG
b98abvLKc5jHTs2UmNBF5fVI2y521fqTva2gOPFlycmYAo1lWL93iykMSa1NWRiu
WbN616ky7y/s3QdhzDK8MUt4zGEa+EIDiAdlw4P4YLA+Eb+rVXmUD1qioBRDRI9S
klCWGUi/tCFjOUcl+uFCPjCHMdIJ4ZEFCNeAv9CV04qWCmgqSvCL2I0IcKOGPi64
vViN4XCRo9Ctyo1ppy6Fp+dgrU5Dmc5u+7fxNDjzAqLmFtf0VYzLvj5gIHg8l4Mh
WWaleGVL/k2E+KJ/sl2FnpOltiTRt0AET+a9COeifKcFbrs2lQHj8bkc1El3jEup
NKHJQXvPLLSPgUADKwEcNkK2+p5XxEoIAmpBLt2BCMB3WVtgMe52cVu3hlKquE7H
8avG9dqlRa54BbzdIYghAQqR1KKUnBHiVyujcq8OMaSBkBEE05+GriaMfrcSX1EO
bfmnhHoSIZ/HQ+DxYxwE1sx4mRX4hakxMIaJ4eRcb0+pvmsPtfhdOofPeFT+QO2t
HOYS47K040Cljl6jueLR/tnDKxw1oor5+AkrSMxuBmOepqWE4AMINyg2mm7ey08c
IUwNd90ddaWp6zfwr7K1Pg==
`protect END_PROTECTED
