`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/voWALh1y0tJvcyB7naB56gx/ZDcUnrNiEzxKoGTR7q2o4uq1uMjzLSeWF2NLrfJ
NS7dxcZd4uv0KmBwDN9UXPWseGvE9FImrEDL1UuRhsZdSKeEvNLhlolxJSTfhYeb
fbc74P49nyTHJSn+WmCLnZM0cObKRAfk1UwO55LPJlpEz2T3dCeKr06d2qoYOlfp
ThQwbQYOC5XwCqOnNbHlT+tAsVT1zIHddOoo9xcp8qg06IY2CeaO0/G1ePu26ZGt
RUOQuZBxF03dCJqxQTpl7lEv2ryKMmRZQr9J4pE5H+7ER9lslZTUVfeAJaqEPwUs
8pFLh28G+Jb6mZMVGSzd05u9YIXzSy1MSFD+OFcUJxGJm75SIIeMI8d+TwUNP0Tk
89jAUu2/TgpfUnUqzciFx8koZf20uxttS1Ks1+nhYO/3oGK6zfgyknx0XHoWdtBR
9IhDLqTOiXZf0qgKxa+XLhvehPmNlWKW2KcRNl5OzXdQUncw94UjJqAlatkwhOK5
0ealnk9oLutborHt2+6CscGCorAV2+rmv1mH1cejb5fURiVEB0M8bu3AOOIuPBrb
tE5Arr7MV2AjsSCKi0kxMpEl71+QIpOEKIcL1evPIShHY+QfKb5EMM42MWzU4YEV
F8Z2lQnWYdkDLJnwFcViAffdFkZNOomtFeqVMGnBnCz5GGTBUpI1GtxBX4QOwsOm
+5yOkeAwEuUOWyMcbuUVo7Yp5gqV1tS2WSy3lJ6MbukT00tlabJ4HZhojTf3J/yJ
jUhifMI9qm6lqgRE0qw93gDV1hpsx8nHhjGoaziL2+w=
`protect END_PROTECTED
