`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifxmI+z7DITB70gId6Y1bbLVwdkrQWgNsrbbljiZCMgyGMtyvtyv9Y6Ro5t8AgBS
qVEJVyghYFOOU4rhXdl9MwF1KEDPxgIhLuxgCpZS/YS1tG19oTRxARJJ+EROXQxj
3esEng5iCor6xMFLzlGAQwwYfB/mrA5ifsuqiQLViG2SW7k4NG+YnUQnHI35NU+H
J/lgxY913bc7PIp9H6wecbp+8UYAEB4belpkiAoAiiek8LWLWtnpmrPN8hDqCwt/
9ypaYR+NcSKhncdMGrj2y02MCCxN6/nXRlh7FUw8/3vU4DnalZ3b9wIBgFnIP34+
W/MwKXgizBysx+ouJBNHysdrft9dA3vYndww1uVJi1I3kfrV/Dz5Ud6L0s/tTjbM
BfU7zGqhXjfQTBlQ8ZX6AUGPNmipyGYBy5MnOyX48AKKf2l+4ICsBZ4b3xhC4D7q
A/GIonTk1hoIo9KgfJ2NJpn8azwJkU40aqfdveye64K5uaRUnoqVaDdHTvM9ifkT
yXaJshcwsxYwGcO6l5mtWls4r0V9bltjtuNMgIV+9mXdbcgHXksfaccVQWGC8vr2
5LXEdKRZ3TPf6LBqHD8qM1B8Vj5eJpmze9IvXqtcOa3QRCBglgaHZQOgn1U94zwF
6FnIsA6JnngrsEYDR6kMOqNxXJI6eecS5A7lJRKoscXrfOOaJHAOqFQIyh5DRyA3
lq3eAzKUypxHD/lWTjtxsD/05GmCRw7Zs6/lHbJL2njhhIPsqAQ3RD2aEFAvbAaH
cCLrosY7i1E3ARYWPg5vjpvXaoGX0LoaMdFsd+/UcQcsLPPUOaZ5v1L4BGxukDh7
RJwtcS6ISOqV/LKoUT1PRVxOBV2vUsxYT0QIBD6WTPUTU3v2xwArCn2+LBj6INgZ
5sFL3tf3eNPabxWf6wUvAoKSVACLmvqnZsepAxM/hKT4mrBrgAofyHgM4uocNELP
v/p8Bs5Ik+ZoxJmq/mYTStLMoCvlhTNTVUkBmdDoA+QBKJvVEqaL2an4HFrfo4Tr
`protect END_PROTECTED
