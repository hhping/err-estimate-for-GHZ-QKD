`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q2v5C0LkhPLB5Ff2u1/zaAQQFv/vg5FTri+KzUgQCqWF7/WBzdc1jPrb6pWZVJzS
0+13PjzL41ssA2/h5TmKLX4WHLfhKVYqE+M1GF2LzN58pJyYqL69LWqYxkeoDeqS
AIXz3RplvebdIl8vM2fAWGorpqF4f/bloTlLiCYpQqqx3xuWfsUYHWbBo8HQOwXH
y7A14pN7J2zPVun/xKOv8h7lvoPTW88WEX3jsWyclwRWDpH0PWy5c2dazdEcJqqL
twe01P1RkMNR2AkiHWyvAOuIQBmsDvlPOu83DsBe/VYWD9//2C/MFu4xQO0KRx0K
9vFLW46CtbZRNPH1wZil3yZye79i0rL6kk/7ZjtSL3L3PfLmFBWJRKQjBCc3c7db
wqJbMFMh/X5czuvoR+/OXlIQzf7DehNeoFq2Nv9moKw2g9L93rje2TY+DCJcjSxu
5IQEzUv8RaxpOovchFUGNo1JBTKmoApnCaHjFRxhW2eojH+hjB+3xx2JP6s5KbJ3
fy5bIDriPKjU35S5yex5pKV+vXBB6u81RSxsu59hLqelTKsw/UH6asml5xYaXR73
SYVpOIvJ3EHpZWaxp7750/6XYdY71NaYevj8OLgJn200xw3dHjm0U6COldj5QtGX
q2CfI2zNo4VQ/zhf0pHUTZKEw2QtiZBpTuqAv8ECgKeklyNDD8O3cYXiOA1KNeng
0LRt1Y8c1Cn0Q5K00c+TNViZG7ihET1cwXBQbNLyGk8BfueTUI/KsB7eKBX9ajTO
P/YRQzSvnuRi5jFHdDMi/oj8eBZm6LkpLaiFpvvbCjc5yEJBp3WAnPJrKBkpJwwv
nDrO6gR4CZRoKlcAu56Cp+rg2n6ypDH3itwgHdGgQv0QVt5tCwCcDM95WqDvHNtZ
OBIXajiDzkuigFm1ZYxw3VdkcnM5ywM3jaUHTC0r8SUkNK44JGePzwXKG93hYPZt
z3C1p8da/reUN7gOypKPLVQ8WnAV2Aqlrmk5uFu8Zvv2wkdzc/PBdsPiEIF1I0l5
sAZESu/Q78EOTtaZFDZqiiO33dX8tUJV0Ed62RXHz0RmTnAA53hig/dS6nlEWE2i
hruZ9WDpV/PRjFsv5flJTYPFt/zdt0a3DErq+AsTHHK47Hn21lRLb8t0Legi2LYG
yAX6ZMROGuuGl9TQXuWrEI4tx39Pt8Jxp0Ks/GRw5f/f1oKcVlf8v3NWA+5FgLiz
ZKV6Cbix3I+Df8cs6HAsFoFDzaWBTGr2X8jDzO8Uebdz6cOJ9ds6VuRvNaHcuIXi
yIH+i8Vu7QGNb+NYedzgBRV/gbqDa8zYWPsrE2uIhwYRpqQgQDtA8Sg6HK48PRVD
+T7HtgSZWzxZnrbj7nnR/wtTFye7Mje9SRmTfrtIZM9dPx8GirarJCIYvnzAaBoV
OFBwgPLwb8NgZ3fmOs64Ntaa+Sc7IQVhCZodMxLif+Nt5dh+tY/8+7Cg7LAl2TrZ
j9mR7uP4h/eV08ZJGbzNnHsG7rM678lsbF6OPaevyse+3OatuJVHsTgtn9CYMMM+
SHEbVL4t8jLGTEkrt36UWQki48zQXDzDjv8KtIgEkTRw5DU5iGUYmXErnque6w0y
ym+RC6bNW9zfHsf36zLWbyEdYWPfqE7mfP/Z+d6PmpK+tYDO2zg+SJoi/8qlMW8B
dczHObkgdhTtLR3P4UHUN2r1xisEWRScOVZIGqDUn3DI6l4rYwwoij3TU5DwIhNv
6FvJTiqjYpgg+Stq53flf5xSn1TSid2CRawqY2bwB5Jz/eZCb5W9WToIb1e9gG96
lLY0eEKa/G09EPU2BaOHVp9iNxgfz7V1o6IHYhSfzYNy03YFnnCypjQrqjRqNb+8
14fdBrXtOE30nZetiO1L3eYdBQLeKTcVE/dWow7f+vdNHuX+Wnom6o6AFNXd1FKY
TKM2rzBTF2DIVOC+nJKCBZwj5bEgePygVfWj3VfmUAxNsXQ9jV6Ynajbh2churUn
pHOO6YRIGDNYIS/mo9j5mJsKhIF2wd+KHHW+tbJ13Nd9bkOwRL7Op6uRYSPRIhXS
4sF6gKWimeoQ/8kkXxaaaLeFNmDgeXALqaS7Kmv2moZh4au2kSbbaVAOPUuZborZ
LonkTvOD0PXP9siPvEEM5bxnYGYgPWI0BtZ9KaHJnhUAbr486VyMEb9AArgo9+N/
h8nxyiLBdNmqViusYhJVWnwlBDilsu7paQLZcobAqBrxgmlIVBxZSDzwL8KSUTif
NJdcFQbHcKZdz1ToZcrlMDHx8UkcKoONKuXFgmAqDO+WYq1CuC5A93Luyu8b7qLm
jFhfkVpPZSNLGbR3OTitYJ3sl/UMxoyHx9UmAsyNCVq//8M1PhmcYQOVN1LkMZZO
DsLxktD5Rt3+1OFKTbmSqrtO5hZ4756hkiH0ZnVTC0MzLKrn69tUFVqr4E+PksGs
dXHVpkqJIbOVjmQk2mCXDLaI/fEDezdDrqF9CUkemX5h9OP0Aoc0DfoMaokK3KOp
1UiioevALz7Mylm8zf+4moxFqPJWTYQSOHErb20uIsRDvqwGKfrsAeqUHIWeYvpR
IvpuFGibOm8Tn8uPu1zYuz8mBOKh9Gby2zEAaFjR2eVg6EbBX3RyXSHhvsiJnqRd
EPisI5bpvrKO4PcFqf/nw3MmYTCabSSftPqqNLk2+ig2UFqdcsiUNh9OP29h1y1m
`protect END_PROTECTED
