`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zW7OD+fiKmkGc9SJQ+DXIlMhA5wiiLVgefXkwW1xtz2yAItLEkjouaEwwfDx+j0M
mxth6nHuaSJyglxR3CvY1YGTeoAgtwQme95wEnMYFImvm1e9wx+nul8TSiAlqsdg
6iiBYbuVsA7eIEA4Nx3Mq64wIo1wixMqRyEnvjFBvXc0niRpZK0eLJOgXBphUOrw
/pDeaFclMYECN5nT3fv+try8Rcr7/Rpl+w222AB9yC24FfHW6l2U5P0RTrRLLcI7
NE+LpbqTovkMt+gQNmfuGGfDci2TLCaAx/xiuOVoE5uZMvLJrwq64m6XFr9T4RwP
DlWCMy6kQ+6w1kjuJ/nDfLGtq3Pl+i/dhGqpt/Gr199vuFLeGKhkT4/hHs49/gYz
cLPpS3kxmmE33BGvXaCL+q2lC7SP3rmCTbe8fh2+29d5H/WXAubK2U5cBIE6IiRE
vHmDe2alYk1oDbFJXJhcyNu9F3E/S7CSPZlDt1DmoMdQQ7zw1xfW5FHJUE2WT5Cl
fEslMRix0pyJcUpnNAEr7QOFkZzAxbEnZMDwN0G6ymaC69McaQuEqgeNlw4ZhUEI
Nib0hSur0WD0El3efHuUT6SfeujA9EyUkXXDMCQTpxx7mbckVUNLa2W51zhY4mY9
q8L465ilTOLSrRqi1KZnGsPaA96POSY6xbtzSRLHhfdXeOde/wb2XsWgWGM+v3lu
R8RPvP5kNULrTsNU4W/W+085Q6gdfmyRC+fpzkjctL998mYssiGIgHv5Z9yq2qrQ
QPhQQDrEFpqEKxk3XHaaWzn2PIgjjTLtQdqS9uy4XvaL/U0LYAaDWU9VFvn6qHrp
Ce3YUT+UAO5ChKpOrA/PCh/mfln3++h5Vdh0q7waabbBgiyw/1IeimK9XJQISNjh
RiFJq/8nd8Qt+0Ey7Rk5vvBoWyRjYlgdemM8eVWpe3axKulJjm3SXbJg4/wfeoPN
zF/3izJeXRM9OupkLsl+gwErg5yQItS0L1xBuJYiGSRYlsaW8R2iyqVr7JviqApq
XB0hZeduCcmrKbwURp0M8MfZv46zClKyDQ6eGyXSeMhnNoCruVBW6YmCM2WTjBJp
zIkfANuOxH8+uI6OoJmLwyfcmrDnhfF3CxqUVRPsHUmJokhZoU0jDXmLFQSUY8iH
z9wmIj+GOu46fAJHFRQNJK1hw1JFJj9DdxtZonCL1rStjiiOhl/Gz6HKAinLoVVz
iAtjiEEGHx9enavGNcXdF8hNWJplAZapeUPKeoy9Rw3uEh3tmif0/Z0+/0WLZQda
0NdjblfY/R4Xy3BK/voZzKU4N6fTCpElctzcgKfaLsf/QsKmeyZWtQ+pMIpsPyqJ
g7SwzI+DotUXH1gUX7j3XX25mje5E9vI92LBqmUR0FHsl715XtSrNMstjpPDa/z+
d0K5jl3fjFEs7idF4MGw+FBXkxvqCPBUsmhBWjLv7fX7VXzkuu7iXXjMuOrnwMFP
LWhsesWMiVQ6HxpCvzS4lQN70jnF//emKCYfz8lWKNhFh+AFDyEYENmbWLJq0saF
9GfROhhLZPJePfjR4c9KsJnkAMwWZ1I3MSDhHYLrMjxmmiop5NwxKNMYW/mjEf4t
nxC/3lPuASpCvxgqE3fpxhGbrcdVtjsKS6hZ1u+Bz/UulEj63yPV8nk48f3SeDtS
+0DEUAZvPHy/K3izOpFCFszaQ/OPZBgB7FfZ5N4gZFMltmZKYH/5vJqCNvx/Jc3Q
XbyusI8+2JzNih+fIRmHlh68H7C9DD6tAL/rYwLLLfZPK14b0P+TUa3WrhkeGquV
NpXUYILxlYrAHJeSf/JTw+DqgYfHyD6YUmqH1cHE/Gqu4/e7mW62pGckhtrZ4XmZ
UO2Q5wveRpAhkV9ODgDxl1NFmBv+um5o4tr1YLbD37JuAyM9UKrx9YGtkoEnQD6j
Pl82BRAADorn67lAKL32TsMP0BKffbp6xyRgM0BvKXYOE/+sQ0YFcfae/LLFCvq+
f2EiKl6klFpvHS1Kh3IF30xFcWIcK2viq4QzZvazS+psx3zopKYr2wQmILQ6D1ls
ojT/V99RSMoTxwNdCux6oIejKCWE9sZ7CL+7hvdjTylVLu1jEKIpm9fudbAhdtfV
65Xa/OPYtPHAkSmCk1Py0TKwofjFxm6StwgMV//3PtTqPfMj9f8HbCmw3lZ25f2W
G7P8RUbI6SjgD5735iI1rX2dvoZZTQ22lZN9cQunhdLypFDtJTls/xflpbn69JfX
BfXMIBcLePrOmj8wHxH02Vh9/UTkV9wERv8xG7xGiGLhFk4znMSF8MkkFGk+c34g
nxV+R/u/0ssZhOSRXtFrjIevaXu4FO2T/R+wepcwN4nDHSkEt6lboTItQxPxfcn+
e3aF+JgBUYjd8OxiOMiJpbdg5Jh+IaAUA6fyNd+kK6EFBiYVqn8hM0pYiv0bpvKT
EuI/tRkoEn7YuUJDpkBM7Eizx/mNJzS7Uw++mTI4S/GRqcQXDaGBgyrCQi7RT2yh
ITADj36LJZ2J9SvbofPSnQ7TmkojEIgd79rmsWikq5sNYixeC3OsfVz9Zrn2CXzQ
wjH9DZBJF7w3XDl/TdoLIzZXavMDq7MXdfPG/xIEmAmAgv3gykM/In/c+QKiaCSS
jxepbBQPxpSQsmrvU+V8EJNFT/osr/ddXq4FXLt/JubzoggvrnddUUSU/NsmKjyG
6UEMIJH1rHzt3PWws9K0y5EXSuVTyJtMGmJqjQ7foPmbqn9enpaYmui+MOjDjlMe
UVAqR6+ttKSW/IrpI/XkpsViJXl13XW1PmfjZHLp9wONgaNg8rSF9rC0NfZ8E80H
xn6S+sfRjIeU7lyCB2kyDPbR56fI/MNA/yHG1zD9goAY5B9dI/UxxD+qv2E/Q25v
jDKogz0HS2a1rFDDYjoXWAEXcZn8AmYHbreYQyF6Tkiy47c1vpM0St76Cl65cH9h
++hnMmN77wNDtWzrkn2zRmq1EBR+uPzpY5x1ld6vY+zRfnDY1+YWxR/Vouh+smTN
KfRVNPov7sDcr7FrWGn7+FnB0BCS4g0oEOgbySS9xWoR4xGIQGpik4DoJ9zGQOGX
Ch7kOUqIwvoUtIMWH0aKysScnxrsfx9E+oKK3NV/FJRy+HZYarJnrKVBAjqp+3Kl
SQvpKFaj1xYKbVjIofMJsmYC21UZzohAWKyaTydL6DsBX3ocZYrZWxumXdQpni1e
3aeM+u9XYRgcwo62vXyqgyGmC8ES6fYrwi9iJYacaAoqUAhzSdkxBDL2k+MVfNzV
fANVtHfuflSgAVMcIBrN/zlNhYhroLezUBlxqEZFdBVVsMEOXTOZiSOSGsyQ+Vyv
M2DBgrVulFyNR6K6QbHUSASTq19MvZHaitw32FaWN2TynoYjUotIKwkjajFiyIFO
ggizHE7COaIBOeoFdmwhWC++SaS9yC7TlGyym1JxGC1zJI/96ImmUn+PuNZWdSfj
u1A9svRLUReAqAdAZbVWsFyuMWpuKPrnSDx11uTy9vIgQIwfDJA/YzDo303x0Zm1
o0kgiMD9Fppy2jlYjbS7e9R7uTGY6GW+AbozPmoO5cqAncQgz8+IgLLi5Ezay0Si
12p7RZV7MAkUN8nqopYVoEsTWpwRBLT6+O4zH3m+6RghUi5U3aqfzfUuTekXYvpx
kKs4h0jIqdil/CT68PTG0NbWxSz/FmbyOTear0U0HRTHg4ZKF6VGBmN0MHN4AZlg
W0W+ThuehL1L1HlOS8yFzGWvY5auP5CeTBBbyfU4x6jCBhIpoLh98Fs180sfV+QR
2y7xiEMzWkc6vwE0njKql1p51wRR12kzzaexouZ2iRIvzDW8XkNKueopLrf3bBAw
EibKBIm8JxdReqsp8USeKWlJn0zyshjr+PVkv7WI6CF7Qzk3yJU1/WofbeUlYbo8
NYfWz9XUXbVDOIiycsaJBHAvicDsVdq9Zg7xChmHHERIHi7oAvmxuQhazQCKQvkt
OdOMq97wYf79uAHgGOAZ5lRNBStBSPjb6dcvtrjHb2kEWWANvzstPy5DBaC8HUzy
lZi2txWNpC4YpI2OpxtPOBxr5wMQVjtEHW489Q9396Sptb+pznRVD6oF41oWj8Ky
DRjgB6nnOqDI4zBSQrS+G1qQQjZrwsK2pCADJg/w/Vl+VfdfBsw3r0QGHJYn7Tsr
kAJ2EpuNRSBWpOlNUhaF2lnnOg3DEPOqpsGmzD2UsArPYZ0uI5r4b+C65JaEl4ay
3lVbYSV2wY2pwZwalDK3k5cWdk1bo0NkMsVoLZi60LN8ACMFPwvaS7vAz0CT/fmY
t64dnq/HQmXT1O4OcnV0OlkZezej+Jto/yb3nRpQxs1GQgOstlddMUNVyV2XFGiH
4JKZuTtPryvUBFq7UHvk+hPmwKZUQ3OqZSz08G8KHazuHyf/LGdMuGDQyk2v4aQe
RXlemiItaKYjqWWEB6TfhmUTj0+YqAev+zLOB0R1cxxKdtsaARxUBrTmlVzhLhF/
zyyr4tzTaNrh94mzuxlfxpZC6Ey1k4OAp/fx/TDk8+5UBo40MmUVQQ8orjKUDs9u
yZ+vw+LKuMI6j/BzbCdktShzcyodtNRn9EEt8pKqb0VuAQ/CIs093kdswYXWky5g
7kijoP2FG06m8UX3xGln61+jvm47FW9ATbkcauS/6tw1JtorYUVxc5Mx2OefGy94
zQ1o3uqFCdHVlgDbLwRJ93Jzls7tP0virlV7c+xM1LK2uvWqBabbcM/jpwwofFt2
E30SyJjSbS0uu6hwazYsZtI2DJpnUXBefPtj68faWbAtV5DDCLckeejdDCkfXy0f
KrRytXdDtu3K9rq6SfF6325lbCnKCdk6saSXpF7MIr0R91E0LVUfAGOvjW4WQ/RG
bzTW48LW+F8AlGsAYF8lc1vziaZQxf0uATjShUCgYUZpkx6KU+f1h95/keNFqTFc
ZboIZAUJMRpnuJA09a32q5pJ3AhIFN6AId5fB0qPWS14bdThMshqywnkZcjMDyre
IoeNH3RdRUtx1chxC6OEc1LeaznAD6VKwGIhPTb5jET10d2Gik31XLzlg5Va6sSn
fElhb3JzuqdlD1Un0v7ie2lRVLO9iShpL1YBqS0dadHyMl5Cls/B5aNvRDjgP+Rt
juZ8K8U/oFjoWvSBat9lfuwb9vEjpBZFC+/2vtcCv+UeZ3rYNdy+fM2iYmhkj529
Pvje8r6svPi441BeZaxFaYWLJegOZ+NSOoI78fA0BcajZ8r7ig9eKuUAWrYKMwBb
cgcEp8/DVEK8IfpynAelQU7rFMIwGGbUrSbwivjOSo15mTWqq0l7f5WKCoyYXyoA
/1+8nl/Kvi7g5JVzMrP8ITCyyxI6zpqy1+Zce70jXWcOHa0ORuYW1/u6szNFk9Wj
1LT0UNdEuclHf/13RjrlKdYTlvc3xXxjuRlT83tVixO2jcEPwUlTGoVJE4/JYwoq
UJ2uerJdraano/HNBSwC47K6MJT/UUlnab2DiCj/L6vReAlooBs6P0rcLDtPbP9d
KlUchyvBtjm4Pogp72xjz9RnovftMDCegrb0lYLZgUYWJ+hamJsudec74VIHV//y
/p0gkRChyJuSTor/MwH9As92q+vG4uQlh5+clxOfKDef7BgtvULu2bjR0x0k/NTP
Pwekgx9ATFscb+3iRu0wH7zC1j6vaRCXhnerKVS4hvd9J/KAJHImURR0SDmEpG2v
k379mED2wsK4k9BrROX9hiCu8lOntR5gqdFnUmT2uftBTfJ0gytS5jaL+SvbYtNe
ovTYDZOWmvuCD1nnWJ1xMrq0JLig2tAaXQXHrVKFgVxDf4JosYVL8vlCNCi6ACo+
VmLZSagXfCpQazT7CvIcgj22f107klnAqXw5d+w2mnkPqrbCsbOMsL3fIEaOPjdp
4szzkqVanKkq61EUhZVOXl8K1S3CCH8HF6yJBHhsSnJ7eVKLg+B0y7qwhqbITrzP
y9g1TW1Qy/8VSk8Dw1N0XGESoZZTBal9yE38cXR09FJiOKHrrHf/3J08ieBtTwiP
90/2XBPCZGZs5vgZAS4RpIsuuBX/eQlhDelW7TI+MbMdgV/K6au2qbZ7su2Qtuf9
aDOpMDurQ0p0hPAFg0pTqYLzd88N85rMLvnwtZwxMHp0CxLzBkssgKBhwqdLxFTZ
aDdD1TKRZUtNhHzchgTKHDoEUiiPw6cfpZYrtRa6JIfkOiY3QAIViL+fWc/iFcJF
Eu8S3TYXH+riIWuPjSmylXXk/oXhAXn2msiHTA3lRZ46oX1KRCKEKrMjupPm/CcL
LfqK3AsEe8dZJM6YHFPDmfECoYiKOVJSQXODDcn0ZzYS/uaJWsdOwxEwiNN1SM3Z
gpxf2t7kIzwKxbk+o0XmgCGLXA6Ndo41O2LUdNMKY3tonWKB1pSrrRziIzOwDwu3
ww2+gS/dSN8Jo1PQxtDv9SgMLFbR4sFBoaLBk5V2OmkzO4KtdK/4GD9K04uHyuWI
tQ7hPixEEetKPSgSHHVcYPfw/628gOc/OV0a/kpFQ2pAP1/SZNQxJi7S51dH+e8A
o8KvQh4O4W/tndPjgfon9w2KAGtqYq2MM7d2fn6iptCdPkpkg0ew9cW5vwe0R6Zx
afJzFtN6cGrf19g8HavLK+htxCFhB3pxcgRRqFspN3lySOpqoxpgBfyq9VmaXgqj
lnPX7DMFMe1GyYXeWAEn/sXqnZUsYnciIhJF46lHf00GJYllot6j/Jpol5NkTdn8
EA0zBDQmbyTYgRg+ptRsmhRfI3qi0nQR9/wGjBmE2M7h6hSOI0qEow3uGKCo4rMP
VJmfo29N7l03cX5fJxm1ens7TfUch3J5SBYVCubfAg1guZFqydlJA4aTOLkyUKIK
GQHZIpvGXuwQJmjcU0bBB254VbR9FV0ijEko5TSy8hVaG212K4W8tFyEpCLxXFV2
F+JUwqKpY7cfbuYoed01nEYZ0AKe1koNmj/Vi90CW48c2X0iJOluV1KPioVGWuWw
wZs4kBW53tf6j61HrFyBzo5ODjj9t/2qctj5TvyQ1BtlJdcwPw3hQFhyt7wFJfgG
5fZFTjQ5sK8Zw5jphzCeSnmI9P2Y7mA6uIXi5gFEEWD+l0g9Amnd5EJon/nGiSfH
DLpPwYfQizVHXVAYcvSFjJJGC/IqYeG6AOnSHp7YTjRoEDgxfBLjTpeTNBGXENUm
A3AnjlWJh4wqsA0AWkH/dKHeVO9cSaA89D6fwlNXjELdWxvMMn4J2N6KpyHUaAXY
WkdDN/tf23IjnTKBO79tm5SJCeFBeyCn4rH3Q4O/qvyb7EaypZDB9PKygbra2M+I
uZbTQxSR6B2SA//Iq0tVM1jf7Fvt4YfDDF5ZM8xl3EM4wTgve/Hn+nX+asApsqnV
EOTxvJUdn3dZn2A5ZjqXv9++wSq5dR1M+Cx3NBai14xkHejgY192jnrhDKBpkBzy
cuOnTK6PYAMhY5U+0SWsB2PikBUsS0dBpHKUGmeNcd+C2RKBEtInW8lnmhb/nLd/
124/q/fTJbvspFv/Dy+PbvVI4WqySo2xzwsQZPJYVDyefDxZSIicASLBuohx0CVJ
5M+hhwYu93+r74kKTRDJxPrDSmZpEElXkGanPpY8uOv2k3HE23PGNZU0ocOQchjW
O9TwPkhzGcG617vVlugnBNCOfdC3PUNSS1aeLYfHm+RrWxnRGjCbRruHjD0gxhl+
r6nah7uCKIiE67hIgr8/pL2xhscppt8Ds1ldBN49vAPavPBLs9jS97laFxcsRz5M
r2e/gBSmnGABRKeZ3lqCp9mrIYd/euikx9NrIlOApiXj4+xg0EyI5CKlyLlQXPy2
dJEPn3KcoYNPBT9ta5TuU+wc9uNKV/zDhWCM19hq7e/fAUicKdeZg5vmbNvw5Yi8
7/DYJ3tTFqqa+9tHe/bhXTpZyja87nleOsiFIKHDN15bhsN7IyzUt9WFE0mN8Yv3
RnJ2Ipcf6/YpHXpkvDvjCUnj3LXvkCOqxh2gGRYfh9KESK+CHca9t9Vik1AV1hh4
oz3OPMdOEO05rDrrK8YIHQ==
`protect END_PROTECTED
