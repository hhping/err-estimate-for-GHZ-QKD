`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zspmZXL/TjLW8Exr6Q0e5WFppzhJSn+r1BE0pds5DirrqSkXcwFmvgSMAyFyeqJn
ye+GxDyrFCe9LLd4rLiTywFN8RgxvduZen5vZ/MUAZeeXUojZrJ6vj7SYbs42T8A
KNLvtH02wpszzEGgb6WBDZVmctpuiOnLWYAFS9tUb/5RyJ9ECgAxC+R09p3/ygwr
at/pQNXVI6yQIf1RlEWzGr6/Vbpy2SIwNbPPsUJvAMlUqpaJGvELCUcjeA48BDeP
m3ZHn7nz1AToNuMFtZGDqUlDFh6BMjHbDP/wb6knO5WwUq/GuqhyL+XVaQdbr7SS
4rPN0FCJPp8tmLG73prN69mOm6GJSVajbnVfP1KOWk0hMtskjpdEhqYrl1Uab0cw
RxKe2nMWVKE3Nc/XXK43OWW3mb6HL1xf0lQVs3ZEQHdqLFZqMFFm/s5k/PAIyKjw
yCGiPhPindzzWZ2mhDk8UJaV6LMaDr/k4CVQX6zxTZyosd8mVxY1HL5I6hVfT5cQ
+WPKcspu+IMKIAAfanU9bPm27OrjpzKvzrOnLdiJY4qUjjRCz1iYrnWvANJp3ByS
eNdLjouZH5+0guYSbag2sg==
`protect END_PROTECTED
