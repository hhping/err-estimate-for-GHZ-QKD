`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aiK/Vsnq1ZHqSRDWJjH4rpFqlklEVkkhtcw+GTBB+mH4v8qKNQxiP5vXiBX9AzDp
ceKxJDi5+9HCdZ1ACP7JVICH2YignbgeVMObmJZwYW5XQryilex2MzX3MGKp6vCR
9Rx9GJHrZ+6G3oRdkIAJyje66h92y5UnE3F52XzZpNn+la4MBjNg8Xm9UP8LZsPx
JsFGTEKdc1BjhrpH71zec5GkgKcnBF6jjVkc7j/TJC45mAqyNTDLn8GbKaH1G2/+
hCj9GWDT5Bg2Ha22qVHEjMw3aigh41TiiasIvpb025sw+tf0bObIiST9jrwZM5MG
cqVdPFYmJTTIc49/8XOxfCRSe71JpvKzZUyLXWhxOYc59jiej1U957XXtDIFJCeC
/gYNHeSGEaK7zigtrMEOpGfnRuJtwUazevrP+MnF/oHmE6jmS+7YVo1Z6Le20l1w
AvfVE5VwtQD/mjCBMA7Lqyi3OK5wxsMbwj96JfAtctSZZCDAAdvJ4qdwHXoztp02
c2VDLwAJt6SKN2Ml4gtSSHxwD/wouTEc1+5bS5OJveP8zUye/D7gC8Wy8HeBQQ74
XuKZscg5WkPZ8+M81dS/VXcWsT2BuKNw83F6Fq/ibo3QO3m3l2fARI5Vz+qn1LDq
ZeuyCvQv+C5muKmIIx38gyoXCBbLqauWEIwisQMPPw+MZNxhLtyhrCM5I741GyDQ
jRRmy1VDqn8B9OQXG9q8LRztwWmrb6Fl17kbVx/N5u6loUZKOnjY4hknrUWudsh+
LptJtWkkDLdTPhxyHs1JifTRl1DOp0VEBAg5gH3ufw5IB/CVxkB4woDUTd7gEZ3v
9wYclFu2w0IUIM9yn4GRHw==
`protect END_PROTECTED
