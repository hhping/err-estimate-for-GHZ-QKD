`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBzAL68ELuLPTqdh3pev2Cg343qp7tKjf1QRewd0aTFjnTNAvZkyXcJHl/7UmZdq
Sfx5pkjifgtTkZl6roa0xtnffd4PWA0smKilYeLB5vfNN3RlSt02qUx76zJGODts
YzfK5yIpiU1jx9+9pH9stvyYDdgXpHwArHM9yv+LeGO1UScBTpk18yF3AbC3pXCD
xHHohftYfy+iyrq0BzI15F8mErHA0BSlMemP+CLkw0QgsHwvA46nGfjQPLkvFIEt
X2jX8xf+cT/rSSs/RH5af82yP1Q7kw4xTgCVYhetk3qAT9Y6b/MYIk7N9mqbMZwK
za7amb2K8O0lodhLEIAybhiNEZ6TO8jyxTK6XBXFHI9YwJbyqM8+vTEQlSdzAK34
F+3k2e0RLDDPzSL0Sv6oLWD4yDEUgJxG+OGyZXpMRGriV9gS8OPQiVoj52NNdwaM
Ze00pS3p99deyCPVZZax0nYmqEQtOaJ4sKMPcIiEGLwERR9W2f6PzlVYrl0oEr+9
sxoN6yhVh3TV/v3n69LIyrmednsIvepEP5Y8g7ypUExm56EjX+2y6g4NFY/AUrlr
gdFEXQ29Nio9nFW7/hJzwQ5mOOEZJXuYb9Qrwq/bNA6HDMrWw22aD+VSyhjQDkmv
Oim5m/DpNZMnz+6oyqX7y6S1v7385MAIQT4j0kEGYkEvV5H+oVs4bE4H/9adGeDR
OghW6oWuLv/JUE0sjjlNnVRQCG+/yHjxFZlGFo3RZia6SfhohH9DK9WdqZ/VYWAd
p7I1MMQ6oHNRn+L0ZFLzWzLGXwQAJWm1LgC2sCX/LkpULC+4F9gJZVQBze7okfyB
70thvv0y8B7aTOFwKwHWaBs3tfxXoW7BBztz3muQW0lv2xAiBO2v5iQdKfPSbYYv
98UBeQuGdWnoMfCrSdHdGPbRcrvm29NCo7rBaMFNmVLe+bJvFdAE4G9OKNQeTSeG
+HZNPludAD87lDBb1R+iCj5D8Kni3G5P2wRrNwBd/KSFV5B8KHik/m6HBoiEiA11
fDMag/xF+MVAQg+Hh586M4sGXi8a6ESDChxfrnE2njRsi68Dso5AgXUqSG7pSeqi
0iTpm1wtwa160RRxAn4LtSWgmcGAfxtoGEpz+F0tGS0CdZ4da3K/YonuuuJRAw/S
yzOlnOPTx5N/RNwD6BDPMwWmlmGh8CfBM8sgmdZQKot/Z70a0fC6sRvfaknB8Bh+
y1v3RGI3142KefeI+xAOku3pULaN1Gna0CC91bCHueqDNKlxDE3HTNKRgEldFUPe
A0i77LxODMNkzs2L2Vy5c6YYPEq2wTzNnD5K9x0JGu4WXsA4r5qmyUxfeVv4dYgS
0fFauHOa1NOoy45wvFgez9D8/o3h5ouPhIauOlw9VGxAUVWS5NiYiVuJL8nUhG6p
CKyTl5ptSlTMKDF65uLNdaPZU/ghYhcfGeC92N4+XJPbNN1nCUGKJNGD2NWbA28W
90XTKfHRao/wgE+9FF51yntNyJkNsabekTtl0Cvoa7e/DeW3dgUqlqXQXqss3yir
KMWgM7ZbWd6G69MT4XxzbjaIaAUjT0mez+oIM/TGg8xmc0UqjSVNieI1geWM4Vv0
0RE3EN2y1oay0yrmw5DKFRdJVcczVcNjqQnxiNCuwf5k6RzY5Z+DeCUdAFwdI//H
U1f41RqklVMmC4NxIpL+yfZqTkmU5YCMopUueKei215TdkJQWJgeVDFyQ4sX8s7D
FsbcZQtQtMaBZ8DbDYq6VRpWkVeOHlv+69EL3zEbVLx7rNADAdnXzP0L7eMQDVIs
77CzI4f5lKJeTaZMzW1hW0EM+DkvRt4ublgafYrcuoWK+wcZj9T9+ucAv7LDG1oU
tCeJnIqR2oPdtOwe19sFWU/WuGKDV/wFb38RLgUYRQAg44wEJJAajfamGaiBIEe/
Uhto68c0HEcP9mUIoBlexAJvw/EyiansMV6Sd8J+3OvL7Hku52xDzfGJUcEFi33Y
SmezRt2hHJ2XjXG0F43s8vtdclJkvPn3GeKVJAuZSOlmJx0MOSmcApE0XkfZbHiF
kgj4+E123aYVV16xSwsfkJ0wzQmrA0+m29xojmOD6Cwef1TsK0WVDCoUPkQ/SFZz
x8AQ2OVT4jmUSx8fgE5/pWcOUoxscwH/2AkMoJxgYcJuOqQmOeJfM465NH0TJwjy
3ry85LfSgPiHF7QeLH0+M3mUD0Yi9IYhaXghWm18EUlRCSlrQPJc7iULY6NQ1GL+
3Cp/vKhCLB5cBMtWwdlelSsFS76So0hCflOCJNAtgkX7ACX22o6+CETQTy3VKVje
Wz+R7dfjwe4K2F1ZQBv8LX5Tz5+I4wq8rbqcfCaBF7D+glzwTR4QPCdqum/AojM7
mQKR6Ftn2qopYqYHQRRrFzF6gGv7NxteEys1TXEPlJ6iCddQ0dh+fh8yXiBimmTW
090BHnqHvcfXTwwnBSy3exfUR5YKmmyvKpiC5H/9XbYFrArvqjoAO8tQlDN/sfI+
J/x0N6d4tTVf7v6yWe2uRSIpE+JWqWLSsl6V0Ji2uBItWoX55pm69eMUAptB+yaC
P5nlTBG5oerc4MzZgAhvJNahhaSzBLue82Oc2BxHB/ayEgvFTQmv7gjjcYrF6jmQ
5A5xeh8/ZVmkRKPOWKLCcvI4udnNLEo1TWqL6B2HI/Vu9SjtO4dDlDaaWX4szQOB
QnJktbnAdXdeLPAUPn3eBXor2orBJrGL8HKAJNPXrjfle3T8/Cm/DFt+RH4FTXQS
+DLS5H19uY3zTf9ImQl2u7xkw3Mhe/tsg8t4dGPPOXN/5uVv2IPoBEZKAodqWxcA
1MG7lAXMnr8fRP/EfVXe7RZ2QYQDB1f8wb4wzwL9QxONqFHcRPdfzu/L+ONUa7BE
4BYg5DJhgi6lG8g+Vopi1NdJWTe7IRqLvE3f+Oki8govOP0aTYd5Fb87R1J8IJZK
CY6mUbcqzzzjkWSCGoQ1Qr/XqW0Yo4GXu4g/vPmDkbHKMliBp9DAmCPx10LvzL4g
`protect END_PROTECTED
