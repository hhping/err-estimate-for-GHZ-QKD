`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1//vXbHpSAaxUU2P57YOcZVr4TO+PwLyXHvkjbiZOdRxyYpeSeMoJ6yjAd7+JDO+
62IFKzA3L/eY0NvW4lNGHXtfyVXfM7p+5IrEqERer1rc8ZOGn9mIfWglD9NsiWqz
vIv4aJuY6fPZXhHASzNmUNr4TOAUxycnm+yXswdUFefxWnLSt4QwSs0dA74/pPaT
Vn65hmpMnjPr3nQAMOzjJrVhq0eaRL88b8yvDcMk1vydUsOYoHos0jdcLfliBgYp
pIrCHhyszQY4Xd3tyZjsFIlSwIEyT8lCJWlh0u3CPD6OtSwBSpVH50yN4m9zBPNP
dKIDsFkfyCh1Ci2ybozK+v5WVOi6R0E+Yueril03qbPhG2z/CmNhvjkJvza3qu5P
bOXEmmBtOCt7v9/+Jxzu+vfrHVIk9r1qXGkFiyPwYoJQZfv0b8gyOesk4TV3vAvK
2ptkYNtdacoGg6Hps5lnfsi/2uaoxFYGqlqAr27V1eiRjow5ZD7Q8t9FD7h05dJg
D51ccEng46VDWhj+1UfQD/PyACVHF6tYZXFQYXWt+80/ELvfKXAk8fbrK+g1uWTV
YNNAFqVlXPwbvOlM4f2UvlBEgK6nXglG/StvElQ60rg9vqHB/YTNCaBSwEcVYdnp
Y+eJ1llebIGbRB8mlyzuAS19sYs0tb31CcJaGrvVeKj0HF4Nb/i7WI8GGjL9REVY
OGdLgOQuu9OvyRTn7EHb34LlfLHodBWcIzhZrDSSUDQZsSZwK6W8y0oB7md7bpPU
Ym47icK+Q16wNmXdnHNYieBB/lnZvGdNlVAj/xvdPddItXjJJmQrT067gTwXZwQA
ZWgBsFcFbqRjSWjmngO6PKCeh9MBtQETqtyOuGIlvyIEULv7mIuehblY8uL/ALbM
r0y/TruiQDNy5nPKBA8espFexe6Fr0OQzT58ykqjoMYalpg7lZfkzV4Bivm2Y1gN
X/8ohjbjryPkrwTv8VrnQwhgYvvPUPOexlqZVyxwx52hLr9CaqLX61VKMUzLyxok
XPy8Ofi4NJH/ctSrtm7lTj/tc4P3Lad694QZc7rLP6B6gMsJyRTaQ9W8cK6G0r3I
Dwi6PBd+hklFnJwid9DzWqkvYeykzkckWRGZceYmTtgWwz5C5/lcG3ikjx+irFb0
NmwK/TId9yFWuk/gWmBEqznEOB75jFOp/3Qa2rwQizeZKg4StzKAHlWpK75YZ21q
+it0rbnEYsAM/e+EAVWdxvPCXUwKF0jAX9REDvyxFgp0NL29VzdPtVzf93a169FP
mqnVK307bCbaeeLuBHWch43b6NPOpQYLtO765vwcgGVdmYqo1Z6KF4k36DjKugsY
6+VyO3NQFl+mTQTo29acgo2WwvDexTWCNeWp9p+OpQH7gSdmXmPcDAQ3y7CU0ByC
4T+XxpdOoRsOju55+dnYM/ciAa8LL3PFgtMqkNxJC9bp60IjjjW2Ssc/UnkKeXZw
vQmhgRla/amZd4S09IiOqymg1jgEMwO5hycAkQMQiHT26K8rz/YIj91XIUWRz4gZ
w6YaiY+xvrVfrwD5sO69iHtfKBKepI1wRjkPYrs2DGhmkDEEH8KTxxO0cwq3TWLZ
UIm66fwBpnLZmBGiGEMEj2z2ghhFmsclIZOEuiTQfpaXTtl8RDK3ko9OBJOT2GLW
6Mw6BsvcezNpKtKVkEAeRjsFJ+78TmxSmx3x4R6I2HxPWHUym29W3l811k4tcEQ1
lYNyzhvzLiaJlUUh1ViSd51SbOTcRnb1QWvtTEkBnKDpESBAGpJ0IwF7FyJbVxUF
`protect END_PROTECTED
