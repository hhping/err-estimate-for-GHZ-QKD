`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8s527JAEv7YfSkMHVENV3XEAyGU3TgAjkVAgVM2vkUFbxh1rPOEQdEDGOQP66rc
GgDyOrxuSqQBYFLjF8n9gHanTTIbZssWiEXg9HaiZrOmnUgnaiz3ODNNlNRD97qr
SK1IXFrT6aw5TRD5T54++jH2dW7nkEEmV/ZFKAE0NCma4lM0Dxfo/RZ0ngutsUwC
hJFlVkmH/MRO++dqydhWlZ8B7TDhaBzQcy58Fau6hSnasxJg9tbdH5H2Whw1AZuw
J4m70zo8Klm3MfXWjB+e5LfbuOqqHdW+q6uqLD9s8rHAtwArJswVxWLB7XrGQYpm
+Y4DS9KAc663ZzW9h+X5L+i0x+sLyRG/ujDLbWgS/lea9JvwTqexPewmvbpzjRMM
eZKdrfOuI9nA6P9dyIBw+M3GoFh7ewr6Y5jqQqWlZGnd4G6vK0BICrgZbB6aAa2l
BBo6P+zKaaX0Pj+6VKRBquApyRExOJ62+lVp3ka4FeYu3iexmYLucdGs0r80PXfO
DQvB94QIO1gOXLxiQlv3YQGlh7+BsDivqcFZ7/Tkwwr4xuvOgCn9GNBX9fD08njY
S5ZRPVufqhxbplVQBCTGmU7+CSg8TOdu2WG+iveQAZ4M311HnK0pYwOsvgcWtnP1
8kCV5mwWt51q0tiaJo9UN4ThgHTiY+iNgdFiWEyMjxFMC3vBVwCm/yJkKafUwwFi
qpqseALt8DDa5fMsQVJ5FzsnSD3z6287eU8ImLIPd/u7Z5Ga8U3G3g2ViQuyppyE
97yYkNLBQKzJpHhG5MeCYriVo0ug/N7eJFVuAKvl3oB6YbcmL5xQ5VDadCuzKrqu
ADLox96whoxNJ/dS3LT2eGnh05ZJzxaf0Dpw1KBJqCMzXglPQ7xrmUJjQS2WXo03
vy+05nnXCr18PLOL9+vQ32BzxZ4+awS7fhfJKlRNxO4O33pscJc8oepGgwMXp/8n
VDVcQMjzF5lB8dsV+o3IozXG1zjPmikLc6J2B2kGgGA=
`protect END_PROTECTED
