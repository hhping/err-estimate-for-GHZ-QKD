`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wGQ4/d6d/iCNWjLe4D6nWvVlerd9mSHM1kwFkyiNbGgAFKz67xUeAkk+MM4xeqJ2
QNHcA+lDZDCh5kd4gfcWzufMFtNFhaAT1iVtIExs/yPbvsQlo720Hhj1yGq0Wr05
5wHUayAS+repj+mURXHSVjWoV9SMB98q1XeH01fI4cTOT2MQODIlh7kypdOrl0Oo
uatURQzX43ajwWUKhyyCumP+74JX2OKAz4oadfSTdClbZmDMLAiIbgxmhguU6fOD
m95T4Nsx2lLFdfpR6XMzqrEhO4boXf70Bprs/RTSOI6nW/Y+Oun8hRVu2xMUztOB
1pax+jhNV58PwE9CQrejJgEvwa6XHeotCWUOj/b1F1CHCI9uY4WkkfDFIxBcPRWg
KrBYDajzgXYoCjlzXPFM4fgbTFV4wElKKR2kR87qe3sunH8NnM6z0Y3dmHl6wNon
9cZ7UP61hrjwgMxIaIGS1OZuXQt+GaiQ7oKOu2fHO6JpSZqZk1owFBPi2b9rsZZf
Y7p5rCbWZ54E2qMbahnTfTw23pbsoYTUHmrmhDayAj59Tc03VzW4bXDFGkzju6Ej
GWk9JKwPNDGuFhfbiBlROGFHEhzuDBgaMGmY9qesjSmRwaPfCNlMpqsCQiBR8LuJ
gKT1fMQx+dt8BaA3w121BwXlLsmCJf7+QCKQNBjL/Ks0vPsr2VKS/4TeHR1N+POS
r3U7LpIXz0nCHbDNetqaGwzRkSFtsPlF+ySTdbm4+SQ=
`protect END_PROTECTED
