`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkbeNQJ6IJmGJxFG3KnMG536zQZOMonuoK6cKBHxHTI9kaGmKZzxCGw32m9t5DH9
FisNzfjr2+rzB28dS1VdOTrowqJwH3JXmnECJvtflkKI4XYP+R0Q8Aurtac4eag2
yXuCJU4VNh/pnh8zRdP8MKJAmS+5YS4quXcU/so7HbWTfJ1F5FKdGAQJSkpORjNw
tOW+StqHS50jHG2qijOvExUFsvxLni/zeczItWoOmEZSUUt4ZWH4Y63Ux+hqs/3V
DfzFJiaA207IWDkEENlOmgFAhccHFyFj5QgoDxJcUo7HdT+VLUas/6P10H4CJn+1
DGSsXOxZf70gcFQLxWZ+iOOy2cXgpdyfYA1C3u97DRa3MUFTdQvzLFUtpUuMfeZU
IsMju0XCIpbej5cWZEE5ljODnMRqNRWqnuxdFWMbYQKwx40RIaf3qPuWSMVoyZxx
Q3qmHqxgbF64Umunp9pITNudSexat1vM+qpYA2Q4SJQzt+Rnx4VjkcFM6DUi+bw1
QtgZoes8ZjqP4bhJ5/BDqEkdI8GIiwRCAT7sgi89kQ2Nfyz6zQHpCIqyZlRPdvvm
Gk9n2644dZ+vvsN9836P9oVlwVchGZ5c22ph1Ru+KwSjkjM6yaYXrWKrFasNRQIw
/XA1V50yiiX1oLsyYy5+WQeqIOv24qhb0Vt4L0JrLjFP6OA1kQ/o/6NY920l588S
klQMtEWIsxcn5ZC/XoHcVko2R4/NWl/c8SFYo44SsDAdYHQSZ9c8KkLFTfsFhugs
MczKWoYqUr5rHTbkEjK1TaooCHp96iNCdNm4Q2eeQ15YDqom3OMltytpHMLO1xfE
TgEI5YjffJRIsxuX4jXTvJCw7dkfCjGtNHUljIBuDUk5XLOmQz5oUu6GgZhgbLmD
pxNAY3Y+rkcYqyGGZZm2LEov2n/rNyG75OWQes/e8lN9+k7Dngzvx3OjVvrYmJ2m
weKA1hho8oMtfY0HJzGPVBDMyNPDWIUWTpwGBRXVshblUoTOY4m3QtTUQo2+UWgc
aCC4qOu0DLIFbx9DYQ9oaETVt64dA5YYo6Df4+XT7waefTNR1vjZyy4y57tIexot
DHO1neeoxZi2jKs5Twe3EzV5b2uDvFpzg18ACyBk6ktzRno7iqwPojWniC7zwIAa
/A1XsLve07SKrE3OLVBNG4qn0zzdWsIx9ZXpbIpxfnFTNqfqbq9o1xW7naQxP+Gn
+kGAJcSQVT+kqJps6m1O6leH2I8A27EBt2L6DVnlfHWgWxGqXXpn1JZIWgL1cp2j
Jx1j6wLWCfG1TSMie+XuRao8xm73D48pb2D8DxiZ4omaAwIe14eUS48tLVQfxGlp
aSpLltvR64FYZ4zGNhQf2KI7oz5FC/epyaU+trf4lRFtAoYtPGi1MTx/+8Em8LXQ
0pw5UrpVpblpgm8JyH8xvQdbDh2PJOPhvEYguACjhvRFKuk10B3i78Sw4dM6Uq7f
GEx2cFISTjD5v+IN9Zmf5fMufgwrQVUubaESdMWKgNI6P7P076YL9LqMGq0eS1IW
otcPvWCLjHShDj0KBcSCdnFZHjRoupciRfa0tA01wN9jJSBbs+OcQYPRJRxiPKiq
a3vyk08TDHZ2IAtzpWRDyeHPDY+fKXP0CVVBRgsELg/fq4cu7LV6MElg9ty5rCVy
+KprjZTHdTf3XbhZ98tjHw8krWRGt+jvSh46ei1MID8DtBRGjp759oiL0aLrH/P7
Dx4ro7KMtr1DRMRTeSfmf2tD2zN21Mr/tV0PAK1I0eXLmXb2XCy1EBXiWburWEQx
qJBKx/iWVHyQGVkdM+w9YS3sPwCyEZ6ukCUftAbSnhqovsQXLai+gjvlwjtdnMcI
BqGEd+OpWdHj9ZJLnpBqjX1uGO3vECmnNAoyBQWjb31iB3TIU9yti5LrVfJVu08A
G8Pp/T8AT/OLqtviEQ8+M9nutI22r6BW5ETyh+QopfmAhsJQBcA7MBpu7/DyyqeU
KJMyeReIEweocFyqIk9UllcJbPBu2GYEm53f8L/5qG0F2jkftTgFkWGiTXzWZips
INosFDqANsv4iEmE5Uf0SUUaSOkqYoE+JxSZY3KdBodCBiopG6ErzD2DylAxpnmW
ecBAXDtRXRjVq5ZLaus47K67jzppQrJf3I5u56aXnJzgo3G0by+VAt/lKO8m9fg7
fWCzpx9LxaCxDnijR2SkuRDQUVXsUDvVxrbYxVg34ymBq7UK4ZXCJV7eQ5PHqS7O
dshBlopMuth46DtsAxwF6QaQjGqvKf3LOfGZ1FGwlGpOnEW00k5I+1Ada6jokapb
/KG05upFLbZxLp2KL/1fOsKs4+EUOF5Y6zAZlERMyPKYGvwgsMKHdGwkJL09LpdD
SgJP3gUifQ6xb9NX7A5fsx1RQXiboeuHg3Q+xVjfbsYJGItaoIVC6CGjpg0dDFVZ
YibjbMYXKz/UfpDKV22Ts8rwI1OEnT65KuZ0B72YniOvqIiRRK+q9S6O5KvGxxp+
mK3HEOe5dU8Szyu3Mrwnmy346XhwYXN2FAgzQjHZIz9dxyt4m3eainZDhhSwDg90
YxXT1sars0OA/YprWY3hmT6UwEkJ2ReTTj5NSsI+72PWyQje0RtmcjSyI7tFfy1r
M/4xqP3cagrWyTbAa0ZMAgEy9B0hOvR3P8m4VxmvBc1eXiwQQGKePTf9tI5COqkr
lXRq0n0ph5XXzh+3CPQ1pe0Thlqw+AmZGIR7suVmYv/4vdJ1YdOpHtEt87qGP1XG
uLktdMFGmy5uIyNwrEh29o6OMYSaaeAxgaklP5Q1C3jXsohEEl7xRQ6U7Cy9lCal
QJK061h21bCU33bNcG2Y/fsO7S+ZjRBLuJEHoWGGbX9df3u1YRCgXZTOpi35Kf7a
ZWfEzexyag4L1ttq24qbm/0divbwjVQmmaJJazkoWVFwQpffygYlP9n6jVvgzKtH
+bWlAX5x3nieCFcbQtaD6gxvJFJSGktj8GWanlxN6fVwyNE5QFRBY2s937bCKkto
htEwj85RFS8tL0VL7uM1N26LG+9uMWlqTr1Qp/bB8u6/3ui1nXTzcmhwo05RuNWy
Of5FdwSkcHb7dP6gtymccHDy9tOeaH5lFqRKLX7hDxQgOVkm90E20REKyf7J7EGn
6ii7v+E6z2TrInuK1/sfzlDyRjtgsHBicnsCvxR5hZDf/JTUU1N8jTNQ3rBd8csl
C4rG3znhdhcT8NvhDmi0RTmgA57ftfdADVOHTU56iw4M4+bsJj3O0KwQUYOFOA2S
N5GwpnS8KA0BtAP9pKOK2ktyTGtaE2MsNVNseU4INZDMsm9BJU5TAUDWEZK48EnO
ksRbKT1AarCXC9sxVmES4s9WaXP3UM3ofk463rpQ+7CMA3ow0Es6wS9D41HE8QGK
yDdCoY/ajAf+nM20Nh5ISqrtTo8SsDibyCLcI/zT14UiATSecpIrt02nuQS+xHKE
dbt3i0VDtQnLr+z/dmPtHnfh9+KAbo3o5GwreRiagdw+VYy8zUwyDkxU6VEYGS8S
Uq8pmtCnqtBlTb6krkmfk2vzRhicYMa2Y5DsppaV0qHitQu4/8eYwTK04jmR1uZV
gr7lpMuLi4CL6wXlyjUqKxPkf62pUB8Rkod+gvw/iqwTq0+J546F7NdpjOD/NZ6n
mfaFoVDCvWppPJxB+YzbQc9VBCMuKfbKVgleVgpP3LQI2cBIlY3PXZvi2Q9lnV8Q
Ubb40e4OPorGRM0HzxZt1V+zRFBo7tZCDWHE0TCHSEnOic/7xqK8XUYsQZBcKqz9
Pj4wmp4Nzb1dvKhOCsp+SJYNWZxWqv2vkAmKLWThacdDwnMVD+d2ZSse6QkM/LbP
eN02/S0uTJxpf/VO9gApgcvAMGFyYRBqkKmq448i2p4qihrc+Le3DvuOaLFmcZ/C
yJh2hV/F4q88UlB83t0dvTwAMr7EhnZYkpj0Y9cGoSAFzJQ72bvuIpvgeswsjDzE
YIQCLIP4ZPRWK4GxQO7n9vtEq6SFTC4FTS7qR71H1XeYX4VcT8pnYdLqifZpi7wU
25SsPbucfECCjmbV9eNWSj+zthqjfq+DXzsBOhZNTpelgP0x6gVMUN0847J+outB
nSM83RQ+XXVbGovAVUuHmFVlGnzSdR4QYmCSSMDDvahkKfkx3MSQAFtk2r0VJLs5
GPfW8bwozjkaWFEfW7GhMMl476c8mryb3HNc0j5vZp3hSBC3FyiI8zMOJ2xS6wXH
q5sEgVLi6mJbtTj8W1ZbmUhgFiXsi30oAHmtGA5TJecZ1/jPcitRRSNj5zVnwF2M
9wYQyjR3vgquyqCBUZCsFOM3uDUWIStSkcqTLBlL+6P+9YEcXbTo91iixyW7wLBZ
VDXUdIUg5UJRNpqphh/gRkVSVu/+ifnubBfmgEZGCcSZ93IkXcqQKw6ktkKJcqXW
G+4zHw4alfzn1NJ3WYM8srCxnzaBof0DmjNPf9Bo78p1N7xo9CTwflExyG6JO3wr
SUzABtCPvme3E4rEz2iiozCg3NeZlrvdfb7GsZUH8WByJ8h2qQKvwTquEsIhALiN
XWPONFUxFwy9tENvI8xfZXbUmJvEKULpo6zXP0R4GV/BrXuATLQyveADF7glVJ6v
SoWrXeatnIdEXwm4QAVghstOO4GonOnU5RIEOp0MkPBS5L4zJaLqa8MNt9+7Rx+Q
DG01UOnNy9t5z2QZMHv/vi+IfOe/Y6/DZxq9zu997B6deb3A+BrUZDQhX84gZheu
p0mC7d7DgTJouOAp6iNrcypy6CjS8vShaEieKaX1JLvZsX7V+345GBh1riiCywjm
tFsGkgbVSCC8hMno1WlTQPzaM0PWKDkZaxAC3ZeU+5bWslb1Y31Sf6xOQvOW8t/Y
oSV5R1d3i+BdqT1MrU218BjQMyyEtN9BhgdmhViOzyIzmlbkeVpS9Xi47oqd/qfS
3EnCxQvaJczyoeKkI0d9NIRGSAwmi9F/q35smxsLYiqAe5tk1WxXa3Az4qSU+0/h
sIb2F8CBUFRQK0kYf7mnOSBHBLHcxMN+W/RatDpCi0X/GrDOh/GuWHv4EqwQ7OiC
AHVCVjZ11pq1Hl8s9qu0xQmlt95sTXzKI3kKw+r+vqdWBVe/nlycVfZSJ1rsWfq+
Z5HAQvqAINQPVZTmlHcEQLPXYf7RbO5PerI903V0VsV5ebxIejkgI7w+oAYP70MF
P5SDIN6QMoeR+w1sx5M38jwT37r2FIp1dXSx8jxwNY79IJphIEQSoatDjNvwHh5U
2o4jNK8iRsEHo4CN+ISCBgj7sBTOUUAuiYTIGSRyxj3mVqf8BXEIJk/SerwA1olp
FEU2GIbEpJG3ejSm1Be7JfeUgsk70B8gMGUaPtjJ7ymw4HZF7dJzckUzMGcrWHcg
LfdhpNA6AWH88Ep02hW0axSPNmHLbX8X1wXhqWCF2Hf8PWLVBEuv4ORt0zCCBWiZ
5ePavJa6w/StoQoZAuIqwUqQboNKqMaX98RuX42FqDg=
`protect END_PROTECTED
