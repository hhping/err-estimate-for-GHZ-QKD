`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jnuiaGWZdSb7ZUys1ewwN/UR0P8HJTkoBfRey1HvUW7nd9WFwpytk2nAIEDlfmy
FKLAZQAgyrbcMChCpaXYJsxAhQtqN5Gm9MzvaJFGdI+dIL19wMxgV1IjQKdy4X+d
dLAkZPDRjxK4CnRZUoAMJsN2RNEznrjCzpdXQKtW/JufhG5XCnaKkihlUmnfc+ff
pbcsrJTaMRDEcQulFBoOjdHqwbl2sDXya0afNUC4m7d/eVj5jaPho+DekVShN8eC
23+sPohClcGe95S5ZKg74HRiKTNsbAwhlneJv/XcsVC0TGReqWZxNy8d4/DaJDzy
DbuhwCD/5Fg3h9awL7PLuQUpGZ4i/SqPLmPBKr1vht6PdVfaXL6Zffq4bgEjSo52
bFmyQWvV0p8CCLFL6fTWSlZHaaJVjWR0UNRzhyPEw7bfJHiBE5KwG2VWgnUHsfPW
ngZmNODu8puVRuF7c3AQwcXwHP3GwniqSGUXHyRQWVaTTMwkJ27HsG+mfBkUhIV+
IpegiixZbXVGH6ODoTjM79bbNu8FklyDXEMicpLjRup7z/PsabMtMAnbJt9erYs2
dG00gU68bgu+GyOSl/IBFGBNpTLgWLtbLWjXz6T9Jf8FRruAOVDKkQkuJieYZS1l
en+R3zU9njYvATQBnw9djoTOCnU9/4IFMtJCpPm78xjZI/ef03jPDTOOKQB3XVu5
ws+e9h2xfa6W4hWXfeSyvGqH3IQ97UG/asIHqZJ19/OXeH3gUHG6AHpigGv9fej+
n2QUg8V72CF6+sjTmUh5sALrwgi1tL7FOGRnKc2fZi/127GZ80sEVgvd7Oa3j1DV
ER8WPf1qjv34+1zsdHAYq/YTus0RlfzjChM3WWjdXjP1B566U7x3vKo4EAmrq9n6
TynyJailnyXMW2ajg+gZ/kV3TamfN8MqkUEyMlq0LD4ExCyJF76DFIct4GvSaooO
0KgaY8bpHBUFOAlMkJ0nTGILMsVBb9JjTysPsHDsSxFeGFWGy7j8sUfyWNyk6lGJ
eXiV0F1JYNokSLLGixeqCRkB9Wrb9xd641SkY7xdmUZM1OmhI0DZ2VQoO5w91yTW
BJz+buv4HOWEPm9ndXME9k1dAZZQqk7UvLFudQp/Qoyr4L/20YkVouXgmKMbNwt7
4kxcMkqleGdMyFDUxVNKZmn/WH4YpMXNW0D2bDrF3CPZeBvCzFYsny28n9lkvkvG
vVgaICzdjMCcbpC6JVvnkoiOkudlauOLAKcDhjvf/9PZmuEXEXq0xAu4K1j3apmo
WaK/PW6G59DvCGmdt5LRoUTwKSu3N8k1o7CPY50gQpHJYM8X0kcdvLOB4BP2NQBe
RHTe/aTVKF38khMW2nuU0EhgV9aJbjsS4ieHKmfoQqF7m8SJDegHyu33icUzeW2o
i4XVGuORqucqfZoJFJbB8dvx73DCR/VZM7qMoyA56D42HLFwKuxqYMSAYKQG2tox
lo3JEgsmTRA+9Fe8piiEbSmUlKqIk+oHHvV423T5Os0z02aYaXiNFVRlA/ndat1h
UdNyoIYPG3xvR191sCv8U95TmCE2TKU+T0t2ghDUPyJpLjwhCCQGYanMtLLmaq29
d7CMYcn86txi36RTWvMHZSMzs876mcjJIGOuwAEJ5dlvl+qlEIcSudv22ATFe3Uc
tO/yDxxeR5rU1//ttoWyfsrRdn/AMjKnvLNvhjblrH9hr5FtK5/nNUWIzLwKDutE
FhW08KEDX2HaOvkHZnxv5T8XXE1ZD+RZJD5NWJ4k9YKcB9GKDhVc26n4gfRFif9n
weeaE0hyP+qy8AbSULY5eyPbaEMvbpMySj4N25bGPvqvfB8M1qHZqb+6EFKMf9tB
kbOK2r+saiE/0q0K4TDKQjt2vZ8cCNzQUtW3aJeBZJ2ZtZyW6aYBZn7LY44NJS9W
evYoJETLMrJJo/inlHx70+3C/gFuXorebBtWNFUXED2/zY3BW4VCMAmfV/X8esrU
GekrxmQjjRK9Z7VuGK4w4q3eDag3Zjkcf2O2QeloAr5KeJoZ3E/WH41ozhN/rIRH
3zl87u+oVEVlCw8/SRngYJr8TBUKewpMqt1YZe9PX2yAaTHTXrcoy/TSYEeyUlew
bdpgbhBLjCFyDT4laPXjNLX84t8n723advpNqVUigyNwcoGMP8GAWk6d0fI1vWcv
o3HBBPJACP8RqGRIiF0z9xJPBVK51rcEUHJWBlSCIliQ8+gUr6xxFhbzHINM6Rc8
bW6ryPYRwb/alelGaKGKpcxG/NHhsNitT/VNXS76bQBZWMBZXiZx8IxwDIkmbZrD
FFRK3fLEbQNnZ5+2htxq+TG5hqQA3zMsASxKaUQOk1w0I4bubCleR5xXbf1n8lzL
opsJrBzEgeZWrglc8tFtTGbAJIMD90GK8luUWb0yyDsVajnWj/Ykp+x5kgNq2Eq0
7CZpjiY/B/GdCqWFeS/7VgTsOEJKjNWsEhIxITIEN7G6grbB30eIdN6w2SPtX/PQ
K5CnoHlOU2E4VE2ycihA8dCakZQuXJkyXlsHlveiaq5i/JKNs6HYym9KoVpbBFwW
MmThrr1uDnWCj+mDcG3m85yA1k38eMhehCROFzKclR4O9DEA3R6fJjijhmZfABKF
A5fZ4ao2BPNkq47+gsrZ7v7tRdegv5r75ZM35y5OOvxS+2BMcE7lGs5e51nrUKmg
3rCPShxd/wkyJiRQb5pN8oGm1tju+K3mzQewpFiNF59gFZZbxEoeBK3hAGC5gkLD
xcjnp7LP+wn61Cy+oDK9Ye4SxV3i0UUe2mWQVlbvNMlXKBHgV9nA8z4t4zKI898Z
ZgeH2b+bTx9d2PCtHQCcv2dj07KVxoM1Sw9SqfpPg0U+3Q0HxTmwE5TIxOH09gqu
1lp262gPUhf8UVKiyFVYsNrjZLL39vh/6R5mWs3Ck2IZqslWfIgIqxIYrVH6AYtJ
YeG0Ubbpynk52x7Lk0NG+Yy94IoTdgJe9MbXYNgx2jkxZ2tsEKENxuZ7J72HENTa
p+as9+AxVxfgGez2nJdoPql4zIsXsGdYRx1EZ9w9Jn5W5BTi/ZMha0DTBA08V2+i
hTqIuntuwJKwjBaLirF9eg156XPlp60qBUPgpGT2wohYKfnzYWMXmn8Z3YvDxCvc
ZUeLR19UNzUlE4UUunng9fRv6GlttFm5iwavWhOeG7wp34fCyngLKuQirNvgfHz6
fenx8fvXlq1BtCCy0408VtYJtLk1GF/rkU3ZzwkbQ8gbx0YjYExdO4Df5XVXZXcm
0DC/ZVZ42YTMglH0xZbMhYn9cf+1UgHOaQMt9Ey/sRKO12Yh0s65jZS7IAh7A0KC
11FjMBSikmCGe8cuez4PvCRxMEYLdD+PR+sqd87tSE4PzpCQoVMfbe/29LNbTuzR
iz3ynrmSN7bEvfemXOJW9E5EgPvjxjOSFF4SGpkzHc2nuNBlV90Oj2QwNfrWR3YC
JEiWkSbPuULGerPJktOTulRIdIpyLkLEYuWScDJJnOQmGhYSy5C4F4uXbnCgF0R8
8GUmz5doKLbFnjMZM4WKnjygbscreZdvwW5XIemVI6V+4VSdyyb6+uAp0s8vwJrn
52b+koxc8Y890j2G9az3uPU79gSqvrgvhm1lsMnnklpEcHoTMqgLMvMCZynlyZWm
d5EJRV4WZyxDemF/pr1seWbb5M6j5INOPBwRl72mh7wZP3BNl/M7C8gu0ns3qKT3
KHlyu22yCG2H8EprjQe6k57skm2KWybn9SCzOOG3a/2AOe9lUssTUOkaTWa3sUte
aWHGntFca6IV03q/At6CHE6sxCCZoPDzzWlahhfHmOf2UcTZkjv83CRs5MBAoH1Q
W44phqASBtmAwTeEWc0SJSCm5TrUd9l3aBZQYNXtWJbxTzDAFNbLZSRexVMe75pS
foJ165UfJfPnJbRrxCRC2htYjUet0Sx++8q4ee8Jm0ueNjnZpucYvpHTCDjgYSsZ
Hvm8thYb7FP9YVoXNoXqMwLaIurqgvFnsaDMQiCAATzX5RmMNy4SY65cyc1SDRZb
13NSvClJ64uy/EZqO/j7e/P0wGzC2zbTiTrlUPEGTj0sh1N3QaCd9bkbK4l+AKkS
7wYsmn+50CZZE5pOgHQEiR4ACcbj8nzTTSNvQ0uD+ulQ7WJK9BK1csF9ZGqJFoWp
klCtAFfeWzuOGvW8ObF8oMmGRHJT+VoxoguRix6O6oU/0adP0QMhS+Va8zOXBJtk
p5Ah0AEoDNODFXTB+Qye0tHJp0oEZGGAzsRqryQBGMG6yGlnRHPrpmvvqIkyHErI
PRjKR62NTtLqr+CiMyY0Hs0YVt1CyRuSIRrKf9kTP8yP7lleDSpNfoEpff0iEQrm
dKyLY9WluDI7d8rQ5TzU96DtTtCjBeQJ5/Wk6wyTMLvXMf4m07ujGuJ13KEra0je
bP3020UIKAZpcsY9f45yag5rOIUaolKp22iKnnYc2Q19nYeQ6eBSaXxtFcxaA3BC
cwKB179sCd2myYlJO55xOB9v94CBAmAwppru5KnWVciw/5WI2m7iGhDeNlH3HH2U
eQdTXNGkNRPeWdqfXZXO74JInCqSTDIMCmicRWdEievZIxn2Dx6O4uHm64yUlu6e
SFO96Us1b+SVuStZ4d8KC9DRxHbjFLdGQL+K3rq6K0958AYcZSXE2YpguxjXeJvr
vtLj1qo6MgL4k4wG2P0UFMI75xGjp6v4HAZqUamw8EiiLY5tcD8CNhybYeg2VKB8
Ah/HTmlVnLbWnUKdX+YkcpZ5Ng/T57dGoBRoam825Unq2aFpeeoqBiKxDvne+eF+
9eaqc2dXg4fUIFyOsUePlPAMOksSZ0UQZYtr7CHVQO2lnYU+T8S44ao26irUnCWI
77v+2LQ0u7lNiseVIo6Xwi5psNMM9zp1YfFNTwsUGXLcvAPnQSF0N00DcikuKQDb
9sUjRVNINUSq9vihRRt5OxKkumiF6a5O5/T/Xb1LVxfyVJ99xtc6EdDVPmm3BzV/
yUBJqSjgE18X2cxsbUGnVkUjM3dRBY923kDIOG7fmSFbVA6G75xkkU90FvbUwqvG
VEQ62OJ57hIIvvax1U0BnUbKg+6f20Vjv4ihlN0RlYmu9LlEm7NYXC1x90ugWgwj
p6mySGHPYdxIspUTv82vHyzTiGQf83UUfKjaF0TEG9gL4ZTYFumeVdVQnBTK1R8f
qw9tUzQPWy0U4GEhnQ3gJdboZ0JEFi+tEs49pPgUKyIgIUXh/wGcMAdELjmWyJWa
Ai1l8UG+VqbftU0p+vbzZgPirMDh/LLTB8X44VuJ6qbkAVTaE5Fw3Bi6Jl3y4Y85
vZzz6fP8cHxgMTDXMBg5Km8sjdqEoQAscon5x/W4Qx1FLTP8Lt+YqLY+VyQBfTur
8wqUIik2MQK0uTtarxcH+TEpn9QULae3UJst5bewcphUA6S0Nl21KXhe6p6Gfhw8
gOt71WSsCdhWwW5kpu5qr32zDjTzU64elvBeNK9//Ze/ZHfxpQhRz1YCVI4fLdYK
3mS1GTR/dMbNvY8yptUlm1prYiGpbvZeuYY95D+2Mb8p6YF9lDD+XI51/RgMculn
GPqwWXQ4wd7JBRYD53DtEM+fKDnIP+/9yyg3iebrtAZqBzUygyV6SuVgKN92mwPO
pL5vj8AiYheNC0CqUmkxchijIXAJmi2gHgPxnp42h5/PCl0DND1gmVWyZEj91c/Y
n8fIiPtxeqI/w0Q2lfHZl6GhJl403QHK4A5kWwfhEcWafZ2jfGA3zHNOO7QJCofL
I7hPRMCU4LeLRFGcBrBnlCVtj6SPMKP3xfe4/eiG/e5jy+DE0MvMJYCnrvinibiY
9kmsTl04GRr0zmiT13m6wIXXU7W+3TcoCHBs5BLrHTqHafYECbDlN9cCWD1kA5m2
OeFfVz/+GfrE5NSDM1yNxw==
`protect END_PROTECTED
