`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXHMhGXwE/XOLEBrvghWbVgREUMdElVhkZt5cGVyGF864QeNJAqx/o5L/MxXZqCQ
GVW2dtY1o/KX10UEp5B731LV5q2QatBB7STiVKDF6F5NhNVLB1qTx8PFiSuQVF0P
xkYBXgBw9Y3vClmF33hmmeexnHep8pNnADsNT9lBqqiDE1v7AGTV1nWvcYSpdnKY
9CjDUJvPCvQ8RL5txe9kwekMzi3NWA8AMHyYoW42yO0TQyT593fNgS0sbv8kiRwC
ZHcUG4SOaEUndO+mLpVLUlwOFEmmjRGI58SU5A1F6a+2v8SabRXFKl1I2p3qSEWY
D46IRjaF4/0ckG9Z1fBOYgWMT3Su8KTrVaiy5A8QMBIff0mECjfNGK4fRbQK3YGK
L5nJ0WABs8OP2wzOMtnmNQoW59vtBNpVlIXe1OsMt2bwWWa2M3cQaUU9SV1zNIRG
gALLObB8NOXQD/eObCMafZfQv4qJzVky/BtOHJuGR7UwkgjKUyVsrdEd/sh0kiHv
wMFXeh/WIvq8mQl9BzuaHlJX+EIfF5Go4tHGv+y/kt9zc9+fqXe96/AGbtAwke5j
5OE5qLK0CYLvCV3sVmIgylS1Mrgi1e2jhxF0qHzZYADyUpeWdVmZthlXCSNiLVCk
uLocQSH+EmBTl3HsJrltmlEuKhub9fwOedw8m7CDtEuc46jy8FJEEZyHC9sbwCNL
0F2DI+yVPoUsxJv6hd4yJKgRrKqxLd7lzzo15ytThTY=
`protect END_PROTECTED
