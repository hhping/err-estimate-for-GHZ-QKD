`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20FjJ6+NJhSgVTaJixhX71ilcLGV9BXPCsFZHXTXcWOsRvzsk5rluF3q2h79mGB2
0M3aMyCNSM2Tay2FngXz/fxymf5UgQxPg56xJzkL7JwpDpkOAxrPqNd6grmn2KJQ
ZZkq3scNJQHLbFE2ysbJwCkb0NU6VxDxE/ELOFxWr8Ie04lawmPTCHIPsahc2qPb
IZZA09sRsg7brj0sIGDCyXdfEfX+CDHZTlqYWmr8NMVo6tJ4UGsEJnkfbXkkxFSw
ZOxtuBQx76paEZBM+nVbsw6RvGzHuzV47Vn9mJIowZjAEkQa5pV1ASkOw/VMZve5
9mfX4MJT686D9uPYlHPK4pbvhc3YlyzA8Twt9w3pbRwxujS0kskLj47CmpbDelYL
l8AITayqBvY/wxtDJ13hjBwLLZax79mAQV22nmhqnjpFYHNwGYvetEQpsIWgB9wj
nOSCGbu5zMEV074zp9WaGwWMEowmIeFLFpbv8lH//dyC9X3d0pu8TTkK+FI4xeIG
/P8x16gbdPL52LGuaeA6z129V5DqwqC4mihfkuyuEVOPdHBBB2PkxKtqIES1USWU
rZsV3uWCUozTET6vHGLMT4nGNyQHi09jbfGHACDxKfq/UMN4EsTiuzKJIZnufIll
Ei0lwvt2tmfW8d7lhAgH131tjEyS6VCr28x5oZANH9WD6CUjzSwGr6KQ8xr7cU4H
IDCaJhQZ0e3K18gnnV+Npgzo/Wqkh32l/yheyz0i7FpDAaWYeEij64nw+xinF9d7
LR3Q0VP1NHA3UXwe84CUnTYP2u6yWsJKtIHdYuPXmMYH4HnR68PPQZXjAORbOEKO
7QlaTNroNi3erQvGKiZNTLawr+Qhou+9f+tTeOqVJALT33skoMzm+J4okSaUIGAw
t9WoiB0cqc/z4hh4kC/gSSuWuGaxi6Kj6C6gpSqIqqaFx8ZkfR8lyFgLxIe84E/p
z7rffGlXUUxT6xd+1UCZl+ihHn1L1xp6VQ9x3wvR2z6UlWcqDseJIovAGn5twogb
h9+b2NyZzCsFycQ2tR5ZffZaysJhROIAoAf/sC1m/Pb7iwIhgEeRQ8q0Eso7N8wd
hq8vTXjHMFkSMmkzvXCcVxTy43CGfMghRoxPRysxdK147ZKEnaKY7XD5Zkgti9lX
I7QggdqAVVCjO4HHlDgncjuQMkJUrDNQdGpwdKP6WZ3AOE4BaUDzKVRhN0h2RSj/
egkjEGEGf8CsNvBGZyoafTTJ5Kko4pMQd7bUtNkSFoTSfUuI85T8lv63lepdTJqU
O7lc+vuVEdPf9HCoQwMfHLAmJ8I7c5NfBhtQaob9sW2ryEmSkrbvnY54XYlJHa6g
LR6JH891WNjURXT6tGFTf62jvuX3Vaa7Yh1ciulgQtwKPczPXoSO/o/LBo7Zdwuo
iJ9i1/Xo8g9tlfHi6IpsjCLNBPa6NKvMcaPhr5XVT5Si6kIaYZ2XdHipK9ygSqP8
ftpPSEUYHn7fia0gGoe0kDk57qr0nDpodb59bLBPuycnXeh1y++zcJG4gsN25JzX
oXe4emKJ2dbMPTPXtP4DvHSeu5CYusKboo0NBcKn6RGSUkeSwqOraMSw0FjBfMPE
pY8Q7KuzarbNkMh/f3M/mXa6dAk6MMgCgylp8R/q6gghEuODB8Cd/3l1Z0hoheTs
/G7U3NMoh9lbtsrNuPzpZlPV4o23fC07LNuM44r6z+ZgEaG8bu5cg7aD4F9RXhd8
e0hzJ2c9ywEvDLCQ/6nSpz5cQk478171QLlkGWKZPC7Lgui3nm3ElcbnZ/aQy+IB
h6uJDKtFpWWZtUkl4X69z4GOXaf90r8Fue1zHiTW//yKZ+jOAzQkBprzkdMhNtjP
2GN7VsxJld/D8vO5orItjK2LwjVEmfFn0WOJ1kYjdp286L6Fp2E+JlzEnCRopozd
bSJHbYKPECtL1yvl/moO20vTe/YPvpJExnJ851gK3vTv6nXsk5Sw9BS4SP4pOSq2
zgv7MA3XlZvm575BalKiVuqCz1RpNCLHXwId2AF3SuhDrKEMbcIOJ23yVAeD9C/u
qSeGScgsNOChriroD1kT4qNKfn48LHFQuIo6OsI4x6yV5wmcuXPOkS98+3ypu1DR
D5JfjAFcEQGhZ70A33arFxOxSNIy6acZDAMtBjblbuZ/HHV8GuV8YFsbbEgpDCGB
EL7mruPIUC3oQz5MIu7Rz2v+ZUNCsOhgf4oKeBmdEi3Vp7HHSqD41KAfCrIwWIjX
CwCAy04xl32AgAlgsIs3jCZdflqdy5OVzfYDoReJbfG3G6qIl/u6q+EJXDTVy9v6
wCh78uBq9RUJAoAunh8Y3prI/m6c48eyzyh6SJ7ty1JwFNxuP03bEjzBdeG6HQ/P
Lx7hL29/GaFohe3kurCbpjxTo7JpZRnYf/dGipPDy6NSx/KojyGg1Dw6MNYjNFw9
+HZZLxBpc3uiUYQUsYQl2RVuO1eIvNTZXQR72zQJCNeHEcEor/85lg2lsbTqnaEs
IWV/9beXyzKefSzXcpT9OugfIwqc7me7qNT49GnoiQ2OwkB1oG9n31Iw5GWIsU06
bYI7OiYrqABix1l907vPeuEvRvl9hfOhY8+EVNOjcqWCkYXHyeQR0+h9XHHz9GXf
HQNj+EEeDslxbrO/ygS9SNMmBersjPr31JwDxcnJ/MHobps7zJn57KJ/WbzA7Sq8
HfGqOKnilF43uiTuIyC+Oqw/WlwQv31hJ4GV1Qsmt9nAXR3pP3jpbhqSIz4MmXZK
JVDJF2aJn1CiUBagKiU/437i8CgZKuyakSbWVTGlSaBx5+wnU6uYUAogafC4hieF
hJ9cMNerH8cfPZn0eJQHH5BWw6SU11NuG23KKNudfmz4caCUGCotl5NMnjcQv0Zb
90owsHPdHuUzWa7w+R67sBnHeZ2R4OIPuHNyLocCSv2mc4n8+EAg7R/kuI8uYTpC
2YrEqh0454lkU1QMzyxtYSNCxGTEWVAXSpD/DBNYQuEn7DL1UCttijFqVzT5iYuc
HxyXuBWxN+Jd+rFKBM9awzt1KQs5zvZqLqocbazkeXEjcDhVFiS2ZcZpwhMz6ACn
GzLA0DRR6fNCv23gP7xfBUU8r6HQk9CpkX5RicHhCvn+Yu2bOUbQ+N5aM04SVry2
4Oei0QLe7ZORntpOBzysh3CMiuMCP/5S50JMj9D8ZUnIStY971gQL38whfqUfsoY
L3lFmoNqqlUvHWa3yrWnK3vXxwKI4WBHyIHc41DoHhi2Zh6Hk3M6vYLqvdRUiiN3
qgrovlP10JNm5PtJdafWJRF3QvOzMX3zK7nh7ccjtzybzNzTXT6TuV+DPbzb3DkO
7XmYTVsTv2u+8p+jwxzP3+pyd7byrSYQRDqOvvQm9/k3t4Zqvxi3lJeEwJRtGjkz
+mdh36IlbodBc8nRbY3WQeNMd6DjeppgbFEWeti4HhRxWCogkO8E8zsGMC5Adp3f
75+bRtyUKtBPfp7u4KK1eK93LPU+SLtdq7L5xmotfC1OVq5K8iD3UNB+pSnW8XEo
DSPA4MsO8NX7f7ChNCfpXVhLB1FDeNMJ80KNVzfBNzhZoU9nze4VYZHalJ+01EvW
g0I2cvXwyIrXIPcM6JkgH5HWsR7orIiZ3DB/Q43TLswQaysVksn5MmW37dLBVwY0
t4DnAdbB4MTwBN6NW/2ryR95De7/3ZRXFqVc3xgUVb76sch1NiPQqMVBig7GpPge
y9d4JvKVGiiOziL3zZThkmrgDLq1Rc9gFTorLCyLJeymX1fBPu2NI1BG4sgb8GJO
rt4meKyZfQa2t/H1UUmuxW1ydjQ/xNSSUNdxsEeJjptuCk1W7GIOQtzVSgOVV8Zh
TyxJaOiXlgZAQB24BlykQzHh3llov2OAFUqCfeDxwUgkaglo3fuF39FSTXnyil83
Zpani2HCF9pXtVHD7HfGsG8KdKbiBA8J5968yGH5l19KF5valE3+wxzQXk6a/jQ7
x5fIkeMvXf/YyUlMWKRNul2DI0RiwLqG65a44Erchi5mlzRQ9s45SGHJDNgMh6Vc
vNYtuCAz4d3uPWK1nn+wmGLPOVE8OLtQ20dwEQLZ97bSg40Pd3NhL6MNabe8RfVl
geVTYMUykerXh/GsDFfV9JWoTORhFcgo60pGqr6frnMCiNUIvOvN7LbafrpcE7qo
hLMa3muOfZ0zRfa7J4K697zEbIOJVp7c5IIIpIsaTTi8ovhhRYg5e+IN5Js5/e/d
BEkdAF/RUvW3vd+/2J2B4WjiBt6bb+6fwnoB3zxzwxAmHFLj/IV2oGD8YEOO161z
4wVdMwWE1aFqQ5Ap7cWMHKnZoWO+c4ioNBGk1KblTJULfxzSyycl7d+MrX/46mEa
FcctJRa5K2HjB6QsuDxRjXcVdUvtar6eJOsJ7RClSHG34cfN8VaOx9gcNx9/7E/G
idrgde5N0OlxcEdQDsdO/wqqKXnhR5XqISF4+5OTJqKM4SxeGoVgsbPl69ihKfj7
4IWHYA+z8LLmRVT1pCMu+efbdM4ZSOaJvu9XE+sNACeAHKYvQJpAgTPTGkwBo4ig
at+C7Xpdzgmd7A6/vwWyRI5zjOp1vqbL7JFOoGT2TraJs30GlBiL0+QSGHId5SPM
fckLcmigesqg3baO666VrxYly+ll2EsIsfbmF8MpFFz75+MiK6pwMG2XHiWX4MBX
zTck3GisgnyXCqtvL4YNzP5rTBlcMvWDof1zBGRhYbxVlyBmUCldIqlPMuhZUxr3
F2HtIz/rqt8W98ErRGS+Jg9wVLdQU9+nvE8EnA298bEbkDrL6hkyfonxR3xWeX+2
Ggao3J3MqI+ufUCLgz7jRejYmq4HrB//RWuO/rxvM51caVQkYyXpHVidTDmvYZOK
xu0OrvXF5FiaCFcB4oCpc/cVy1gtMDIoqgMV/pwEbdzXgD1O6wkdQkHDlVSqrdAB
L9wYAzIYb3adqH2Pry1claZ2vB2tittA32IA6/taQKdGFQQBQ+z6AlNS+mvVVnkj
U90VGTyOLb2DLhB4GomzEJGfLF+vgoJNGGIVav750MsiR1YmNE7VIOcPYhu8tRxX
wGFKynkhq2bVBttUboEaiNw2WshdiGY4w6SdfRWGiJiwqHg81hKT7U1EJ9i/GEtA
qYpBSZFdC4hhuBIu+mGEeP1LgVaLKx4xTIl+MRPp2nZHbUX+Ve3awd+Hv5JoRpPv
te/vbROHJT9/5JcXEA4uEOParVXuN4Ja+Hg8zUoTYq9NFOUu7oi1mLbDlQbzP8PG
9JMhByezEP2jZUfUjl+9gRIqC0wJmWal+0OMDuTi3lq7bR8TLFaXaKYerOBsmthZ
mJ0BCieQ8dzKLPHsxiVLjMNG2aU44nEMFzlnfjBBBLr9GsApIH1T+RAvJ2WgZ/WV
EIhkHN28Dj5Sx6OdtrhmoVfiU/spRHT4X5kRE9aMONN6aok3rMYaUAjrYVapV645
XsuGoets3iqrcY4wh+q0iR1HWj+4RkYFH5MX99CAsPXaORfjPNtBOq8pFt7hdk+J
DrfYgJd7VEeHrUSutc0ZtmLhTx5Fn2JmpBOp2s7IlZNmc8Opsr/RdR5jM5YEYqqW
fDgju9QDmnlrAfOFlo8t6venm2n40i587b88YNeUCIDZvLd/aHKz3l44yLUYtqhq
gbxVoPCucu9V10bHTJe4CStEZKYFNUTnMY8jnSXujQZvsrdUrQwbCl8w+KMHoSex
Wh9iOEbUJcoPMPKUG1OrKFY2Li+JgHuEURWgXQ6+Yh8CN9+FleSbz5LNMUagDzVG
TK1J6m61ajz8qrQ4/mHPFMD7gaCoj0sKQL6qgqhaROnf99MtyununTmmE3lgU+z4
tTMRy+ppydfY1vlVPJKOjDDyRf09i8FsW3dLrUw8Vn22iupZkL0hvx06wxFKHIxn
hX+SCNnRizhfvcNkLZ4UTVwAICcnQNHY8hDeAC58iFd7Rqj9IOwIHaxxy/Unz4TW
88IPIG/VsZ1DOJ6YOc7NWIVIAbHHJ8KIsC+UwXtzgeZ/GFObfUrQEwGA8EdHA9iw
LbTiOVz2BzmqH7Et7Zs9V9TFUkusLO0beTfOIQ5dRHIU0t/mmY7Fof20UMtMKbWz
z/Wby9qQni2vuI5VAHid36Yb037hXPJA+3Ui9oSwtpnwK/rDKp1MbVxFiDcRYnqT
`protect END_PROTECTED
