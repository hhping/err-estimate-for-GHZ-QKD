`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/v2Cq+jKKwqAlpXr/0UL5s68cw3oSr84yZSv30Cs/Ma/lfnCOgbhGiBLaEo8mLCW
kDHM97duDxEcTqjO5S8H7BAg7kEYvLxhaqhRu5m5Totqa1xGlGsIWoN1qXZhyjVY
9hD22x+sTv2X2jpjkrgxD9EAZSSTfXvBQ+B6yoKXeyOT6rcWANCtJs6UiEwyBQ6r
PRG7v+nrd7mFmhsa3xSuCL4QOxVHFY9X/ufunv6lMs2OeZUb6XY3sZilTI8STwle
TeOv2dnvVJX4f/BbrWVIy687y9+eCrs+xrOAmvIfJUuI+OjkyWStyvSxqXo28rUX
oD8h8h6CvUfR5P4do/zbuiIHFYUqlI88Eg6Pi18if7usFz9N/nOidQsoEKk88kvO
Gd1BJvMGIdaDJ086vqOgDOYfMh1Ci1RRWrM+MdbrPcwP2lJ1G8FeWocoTQv7mnci
m5xk2Id5cVNHOcsVNoNy0zxFzanqG2KH3zpFiJ3m+8bS33ioeu4WMnxwhQv4sH8q
`protect END_PROTECTED
