`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q78kt31ggspbsUIW2ORyS2iQGwjmz9jdNlBkAdgadGQSX3WB8Iv0RjoJl4/nmyb7
kDF0SZtpSY3m9oPXV1I6VUN5a1s+SBevBMfYfZpCMJ+2cUOPJJGXJpE0TTIj2ya6
pP8y0vJAQVibfnhGgfZ93qvpJ3yJkGyqzIwxbg2imGOkGmO2x8qoZ7Ls4uPuZF8n
FIStMSQZBsW6qAtxBJXclo1SqTVnst/tXQV5vTSt4V35X6aUJWTca0bh7Ok8/C1l
x9+Jaym0pKnDf9bkYTdSQfoXcQDYCP2zbYlRiDdLOkzoIuRfaivw610h/T2hFmAf
gdu8ZoLvMq1dLxLfXwhYvb0fubMgAAAfQIWJvhTkU/1dbzP28UPQjRLTTF+Pqr4I
H7/lAxuaQLBK27Y1bOBqTJSTCJ356D+la+kRtHSPdN7BbI3jwLDdTGrDALY3Ed5W
ePDthz5oePJEajYk+XJhz07OjUzvtwTx60WITkjAi+W+xgZ5avno3zwYFiW/mJc7
AEGFRddKfqUb1qo5HRqVxbuxLPIZ5qMg5jGckZndSa9umBy4c2xhwz2zWzl9VKWl
6INxlv+WFGDZjt0/WeWtrS4MDvPrAfzuK0B/JRZVNiGg4s8aO2IsHUql28wFW//P
NRM4fHl20xQcHcxu3ryB4fUc0ySJfF7ONmnwYdtmtSgHKiHHvcPCBTTy7HmADqGd
`protect END_PROTECTED
