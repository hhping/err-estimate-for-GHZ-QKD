`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLorX7A8eY3adAmfhLkcj4ejO+pCPl4NxMUhBMUQWPsEk4s8BITUmqPOtV5RAiGg
PVwx5HjXBbWhtLjfnj0WR4cM7TpdFJ1fZqpBAVXFky3fSzeHxql5t2abwuQ3A26G
MFcVI4jGB41BTrYZ7s+AFNMMWWNgCdYsJB3ByvqpIZv77ELb49Zyn9laVPmwnO1r
G+gssm9v9ayi6WWCmqSFYw1f/fnVvJsOgrli9+j0os7nJPQrdxwUALOXwIY0uu9b
Ct80hXn82Did2x1CRCTd5wJgiAhmgkA97nAh1iwe8cOfZwXTwb/xdS98Ql2Zg11s
ylejK004ca5JssiIoYcyQva1iefsUSrl+sAybedm/sCFSzOLheo1OmZue16B0yWI
0TcZKm9l9yVU5yBPCzy/pR7dugO9EjOfechSnqeSvXo9XxBFBfyP2izy+/A8wtol
+yTjKxO6APamNLLVIq/Wql5X//3k7BsPKYqK1Tj69m7772/lSImTbEiSZDSeMukC
dyEVWFp90KT4R7NDvuuER/EYed7DBPb1L5+r/NgPTCfliXZ6Y7FFUwbK8bXPcck3
3r9AmB32KESfWrjcZR13znJ4t+uHElFcQAPWNC1pHvAKULLppxxhFJiCDsx5+pdF
TERAD3WxnAqhwg6dcqZM8tI9p/7NoX4fsu0pqt+CiuOUMEcJNgVRvmPT/uLFY2bb
/r2vR//YxRyu9r7r1pcHgmo+sR9O307Qg0F5N0b8wr2k5u2x8qjYFgJBjnjOCDY+
25eR/ONu/s5Q31d8t+rbsffXN9oDShzh412GPNGkN5+du70FepNHyjgHlxJ0b2dX
KIj6Mc11v6jyK6ETA3BQ0pErp9Q7SxK+grrNClw4srGxg1ac9LAmYqDf/hXWVvbr
TPuQEisbwSjPJtkuGoMxDEjDkQTNjNOBem/hQbaysNy/3v64VpX7Cg/i4k1PI1iI
d7jooExiaGox33qLvkt1b8fHiuS9CyT289FicP2leOTm5abHVqNnELlcv1kuIhK8
09df+HkMD0JcvNpj8K1V+87ayLKObzD26lMwZ5K4Ll/zOyqq3VxsxilAP9tHf7lD
a3zBfE2AGMdYG3/W4GmS9UCCMimnIfsN3vz5X/d5KLQ68wfAC4TGnasQvqLhBieL
nBc0iI3L/yHTzpCqH43y59p3KLf7jblyU/oW2CqQtTeLaUaRB7Utsxf/kTlwTpKN
e7GSFKLlCFSP9RFTOW2DrtlZsmkqN0OxXEiLSJx7nVnPG5SO0+p7/2Aa3QNKK7dR
qpewdM4tS4ZpuB21h/qNHCz8LqSw1PSvrN+aI5BG7mvM9/6nHJ+xcFnQLIufqmxp
pnvrRRk1fWEPXsiaVEDIXILonewnY0XWnXi7UfPtsEJszmqNMcV+SiBBYTA7GP5D
xui+k3xfsyH+vMCizHXepYDw7qo+3KkR0iANL8yhw4a+N5Rt+tyPooXe/vzjb2VW
t+tBj1fe7m03JKpXJOkVAhv4j4/PkDWxWcLmHoLKXtfLxfYjM/r4wk7iERdjdW2p
THxSN/z1j1+NvI4YMS2Is4iHMwPw1WcpFt1zICNVjZDJ7CL8PljW7OxCrep3VEnm
x6+hJdLnjTWG9bIxnyl/d4mfUyZwrSswQmw1rCx7pTfuC0ASvYO2wjwlqPlbvt9f
O+IMtqZsQhCoW6ZV8iHX/Mo9ucNcJqIMIEKloi0cHvHtotMAdJcjADkJlDmE0Dzr
MSvfTGcZDwzAaChZWifPLni0BTCXHfpxEWFUlUngvd0aWBKYmJLc80R3XBT/icj9
pGcOLrqUJK9PMcRLkVzSjQvrRCYyYXHrwFEDpgjOlXn7nsJ33mvcTyiQ8dsQuXJx
KOzISr5UDzAsq3IyDW6xLIY8BAH0F0X1jEGU2VQ8krs+pz7XQUkEtbzR7DUeU9jL
RFEUnvjWKsM9DhenYuo1X/t9EtDxO4hKUZUlS84/HRyh8FpE1Ml4BLroIaVUyFS6
2lZqLmKoc8e4MTxF52Qof+7k08yR5OqzeBQ7tCQziDZqCWsivtrjlqzGkDzgqmeg
RzbLL3y9YWA674CYGEr5aTVnzZz4e1ukL+Uk5Hu/VPbJn5dwD/ehwJeRg5eEjQ7Z
SMNlQXXbYRZP+FCSq96XsBi+rCslsrVGgd3RwO8fHu/W8fzGSULXbOiCdCuSDzzp
vv8TxQozrUCCqrW9Q/DAaz+KkS6RdAigRK/2qefXkWSZhl3WxFLGBmVn4BeTiiyV
NGMqmBtfjyVH3vuw6Y2kUEiWn+nbJHgF2biB0X+1jg7Lvk9x5lIme1bjwKv24Fuv
Pof1wCGaejPBPAUmPbwnxxpmZbbbrMNkxqINf0O80gQxumhapRzm2rRpyaEDymgf
xBvclfaMsHKrHZzp9wGqVBI1+r3h9+vuj3r5fYakrAOZ3VvXuqFG4nVprv4iTVQA
zBYJ+N26eyqfAwun1Djj1lVQEcpLlMVXZzkdS4romwxaHYs+9WIXdtB9CBKxytjn
DFe0/PweQP5WKOFvCeCLSwPTNnLnk98tQ71CqV2ti/goDwecyx4yXL1TWf0fbSlb
eE6UXUR8iVY2tX8ssxZC28QE4nuYxlCDf7YEoIOi/08kSc0QK+YGiB81VwCY7gKB
M7OV2LHuDQSjTGXozAW4RwRAXC4JEOKFn+TagCr+v6jj0OdqMbFjfIzFgnzdZCF8
whQF2z1LlAmGRWnBMjXEI7ODBWJiBsFLjiqU4guPoBHljjBJhCHEHFXal+C4Ha1W
R15utSPg7773ag7kVV4fWXiyAP2Us+hu2zguZYAXbCnQ8emqqo5a9UcwuZ3qLVTz
hU7n2VNZfEAIKJVvlI/hZ7KkMmsx2GrqOyW01n7PuKc=
`protect END_PROTECTED
