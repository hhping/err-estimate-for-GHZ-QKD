`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZT/i2sM6jtAU/C2cyJQN6cWRcHN5eJ88zwT8+FTjF4LDQ6eG3BQ/qhai/TzWZ8C
79S1wp93Uovuadu82We9qEH+2++tc3XB9xB4wmS6+lUTPLwDrLVx2xoeCQRdM/H1
ipFemsuRPyYOxEU2CMtaxGKv50pocMowP0Bo57nk2mkKX9XcNhvnyOfBiPxx38FZ
fIJgomFkyMR0+fOPoYfDFfkMBiWrKof/GBuYMBoMHOsuScMmtdEeuIupVE8hI44q
zFh2UIFhyAwab7SUwW6U35CeozCT+jFhHoIZirSmxCGuplRmrdtiky3ZMEgwAyjb
Plr0Id7T4Zv78na/QJaEwt4/Or+Zyvkytao83KS4C2V48gZKHwjCyR0H+ZaiEUTs
czDd1XenxRjIvszE8QAZyELm0NC7+EDN+oDS942E1JcAj+M6aliKvdgeBBYss/vB
A/Br5DYHrGwh1SQLP3PCSyaEcEkxlZO5gowDtV7Q5tVLd9TFbwaqnfpyOPQzOjfV
Q8ZxRtbdlj5pTiRtwpN+4VdJMSSBNLhOd72xLcr1U7BRgRBzj3bXVQWz32f9uxlZ
NnDGXPWIiX2LBgY/qbGB/O6B2dBnkLwQDGC3MNRs1HSrWrQg7IbLV1i7pVGOrnkQ
/sTUScvD8qvI2275XgkvUvQgXNXetzBQWIdAKxPTOdu7Aay0uEnn3eZ+ffn7y5Vx
x6zcqBD1+6edy5hjTI1BRsN3gxqdKaeH3Q0zfaHnSpMqydwKwxUrjMBNwHDyrLyl
6wT5zn+MHnEpedFrljDCCf9NpSBH29VaQX3Z2UrDg0fK9YQmP5xfIym5Wy0vQ+N/
If71mCpt42FA7Hob9eDrYYztDV0DNZR1zc5cWBQN+FceBCuGFAAtFVPY6dffCcAI
`protect END_PROTECTED
