`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GxLwc6Moz1tyl0x3hirwcymiXOy1gSzIWeR3GsQ2Pp9dmLRVCZulweeMl9R5PtsM
ENcu+1YJ5lRi0b+tOJ8zdsZhSjrTKcOlOa829At4y7PjuA92FEGri7BDJDoYSlA1
rOPuVOhKaiz9gznR/tGUwKgjWQHojoom1+a5AeK+niLwSIbzsA6vsK5XsXJmKl6l
OE1IhPOCMcpupgk1wCVi4XZ5BYjRUCHkyTwnCvEpOA+Nb1Cy7KNAhIwgRL5rB/aJ
jXSTFjKw9QRyfuRTV/yuxqOvOfjQJDUmjOvBFPjrMtahdhodI9HdCs5TfBqI48WI
zy8R7zXg/o44JHtr0ZZYcVKnrbmPuizbwoXvAjRKoUqSMz2VrR5xL4uUzYkWeusA
MVDSFO7HLWNF0JeilRAwO0AZt+a+lmptcxoFHClKO4DTA0GZs0dlvTIjZqEf/Oxo
It1bIuPjDsjYh1jXJoo5YtmTZjh5AQ/Vx9umvbOcYa2baorA/EzDgObiBuvFJI/M
Pr5dixwgaJmbbxyUaoNm9WQP4KtaWXSaDyQaa7ZGcC/uxnytTRumSebduaQaSlax
e9iT9QW7SBcnysGCOzipHlEZfBHiMgzPBBK8uYQ3npdEO8ZdCmlIH8bELCXpRGCN
Cx0fjpDu8+lutb3Vj9+wxZQ5U64uUrS2ua1LsehQIPPCy0+ADVWBp8aZZh+H3+ky
NIVC0kcx6fKGQXUWNvW8ScOBcjzNc3aLerFM2HxueS66uE+4JMLi9Hy3tOiAffcj
/KFVCFIyDBJDqv39/QFQGuOLgf3kHHhzuPqDs2Llgi0LNZYo+xCXU/xiHm1Hhuo+
Op9Q6+bxSxZeXyB70YsPzKfn5DwuRf0UJmAGnojATy+Ls4uJTIwZnAwKPF2vfIWz
ZixUUbmFamFn32ArVarvTcrdzJcGRKw4/B6WCDa9z+um+l0ShHapYeE/R658WM7I
YLHe8Eazw7hITfNGIG/0B9VIde+Z4GbaGchj94Vng3DIOTCuN/GH31SEke35VAPZ
/H6LmxzEVQPkNeJTv5ab/JllxL19y7ON0wFJvb8cRuSGG9paDj2LE6Rxwpjrsr3I
AQSkgYo9xPB4ZbFjtxajC49pd+e1w/KH7e0/YWQbNnpCZ5j6ZVDfad2IQtEkd/yq
JUNeiFCkwCCk+aFWLqPe2ayWwordD0hBX8rG5iywndFDX9h2odtIiVWDVP3ZUhaL
Od/5MzOpBRqhpbnxDDVz6ph4lNyAM+SfTaPK0gb6M/omUckXtAWbWxRYuTZnHjBp
jciObWzv6zg3VceimMyMWflrNtearleesz9EbKAkeVLk+t3n9noldFPNGiOx6L2O
AMqVgrDSTIRfYrzNjLFNOqPB26AdEZDft25olLiX7jaQ9yXUNCWR/F7FIo1BgPIA
NKWQrr+GQMcRD7A6Pyw0uGbIfhDWhjw/45OMutJmG3D2CkeSlZMGpmBf5hzFvT2d
`protect END_PROTECTED
