`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65lQQI563wvO64MIGQVjvoihqf6UgUdp/gueXjuyEozVK4j21/WJJEgbWhN9rFp1
SANxmh1OzcfILvC94OOqR5hE9uKOXSok5VWblUjV/tWgqY3ED96cuN77WGT+IR01
UKWX+JnidX7r30BtamrdmfTM7VBzyRL2OL2VcRuI/lWSVdOSZ0H+k6TiWan5/GpZ
mt1VP0/mO4u778VhefxxCjErKaOvpY9fzix6pxZM1qPPNbvPhzBPlTe2hbiU/LFF
6TOm0zMSSJawYosrOVGNMp0qHMUNOIkGqi8eR0uJV3E6yok/FdrAU9gNUz/E4cXP
6NydIW0gMMEIAAQ/z5Qm+hlZ8xsBtsBhzmq/yLOMGYzEk6nf7euBevoEKdnvS+lk
ebc5mUEGXN7syuNlOc/nag1mkxhbtCsjHQveBIKqUq/OkHUODi9PqSgdPSKxRzVY
5WeZGaWG06kZCxdbnJz4w1cKqpPLFvLQsvpeWHzwtPN3/mr/9V+zKkw4B1ZX1adE
1ZEx4gqKE66Yx7oAZ8FAnWFnL2pJEIiWHHUv5rlzHZ2bbqn9Hbk+AA8ENu2o7rRv
rOX6pideW0tWPuDVD5V7I7lK8iMJQMEBRqdOW29W3devkOuyeivHwwsAwUTJ7amV
/kTYa8enTkc1m+NgjVojAwHlUDtB17EQzM61NMJSPr7Snfj9zzpXK4rIbntwBJ5M
ipwoEmK7qzUbfP/T20XOrCNKI0mqL+j6FSFqRc5YYuYLHIEBpLiwFIeyect4YHLN
SHkIajDYEbr6UO4PEECZ/6tI/NKtc2NtxD+wDmZ9enNxCB44W7MN3Oe9O1siPlZt
/X5zkv6et21F+myHn9JomCc/X3Z6gkDtcfyOfmK4NQsX1uRLItdzB7dH/LSzIa+P
BMlobnzot3uPR1mx66JyTV/Ceb/qHIKQTP40nE3xy+GqxafETWr3w3ykt/b5KO+k
oGBBBFq4wMB35bQwMqpnihY3CiGgtuie0Ye8n2Hi4Gan3YD9/p2WCnrOpr6JQ2ON
WEO/HYJ/M/2FygZA5DTOqC/Jj423B3HGUuRL9UBecMXAIsCeVRBjjILiYxadGhOt
sXpZszAqjaTTo5Kxms2uzs3cQTd+g+ENPTvmW3eGhQGg0pK2Dz38/yKH0Nkedoyn
HQyGYk1ZOcHfxRBikEb0G6FBClqk4sGiE3u16GAbFyBluo36TmoGM03TpT/4rg4H
R9739TZVJhiPEfGNQNf+rU1UUDNc6/DmKQGJ0HG+gq7BCwcROMFSm3uKNN5DMoti
0dwUcaSew2GLhwJ9T08jemTWj+HgC+cMKkrOLyvqWFSTJ9so6aR60+5cn+2mVc/D
8dEuZZAbcUSO4RH7H2NCLNAh+FJXPc1Gl18buZWSV2FKt/watt4Qtli6CwDzgE0/
nj+1m9+6XyIUHrKw3L2y7v3WQiKyriyaeDok86ExJpdk4G3qBLZqDzge+bGQKPRF
tz76XngJXrIcPq3X9aVfDaGeL2s89QLWeGxVof0BPxoNYqLD4QYpJsPinJgwbXpj
H4NujR9ZoHGFBp3OUuZ6WE3A1JvhdIpXMBQF3nfe0Eo6WjGWsD90vzYrKvkBIWCc
nUNrMKQYEn7vkIcJTyUTYjI4LRf9vrEnVmZFSRiZQss7/5xaGMEq3on0Gdw7GLDB
Rhib6U+rKCyE3IJ6yBXzdzDFScPZJ3HcPuu/ItgWmFLl6QIpBKQCfVW6WbZlCm24
X2P1fFilbTUqTv9t8WAVklrYVjqWRdKaLcxUYuZINc/cVzZiNrZNM9SqUD/UliNz
/EMl0NN6e6gjkF0+c8takzgUWUCgvTiidxYPQUgGa3enfqkPfHuYz3GOS5ez9OOh
4gyV1qlC2sSyxUj1Dlbah0WTw+jrxETOYtILQdIPo5qstGXbeyW/++/S0QxkZpRV
PYEY2hPoIKrMMVI2WiNyODn+HbTrTpOlAgkhb62CYEBTSPDqoxVDNePkroGSR1Eq
bf+jiwg3gmmGVFVl5TbiDISWGhML6dZw5oaQcn7fv4W+zT17kmxhgIikG2s/tMAP
1ddqIvsoviS7VDeEDQeJmEqzHAdXDhpuldovMW31Bus45z0InUu2LQ2rnrYKygDh
4iO6thmBhvE2K/xUgA163av1Om9rULl7yPpL5HUMMSUM7J/CAPaV0tKCA5rD8k5o
JGB4NZ16UxPlBN9rXKjG5mdTWVSvKpFZeNJj4Inkr9eSoN24xYFNtdrXjm1xYo36
TSlk5wV5YszHCQAL6OejBQ==
`protect END_PROTECTED
