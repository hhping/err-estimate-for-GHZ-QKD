`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBVGv85uCIBCxqzs+n5oxDAfArtvLw8DMN8EHFko5HjZpS7zxB1/BxIQfL86lyWa
bO2cMxqPptHm5kmkhTIkddaJ3VK0xHY/h+eYwvvCbD74bZPuPOKr3f32ReEUnh1l
WedO3viJ9clVdHAXWyKl1ZTk0qnEwSbOlYXB9JZw3Xm2rJ3hVUXdVGuBtypNdkR2
0BJVjSQuBN8Gsyxi6OWyOqoMWWa4T1CFelg8sA/9RR4bxCuHYvj44PKpbhgVj/1x
dLuiWHJ46MjRZGne9ewspd66DBsW6VHuAOPXjqmLIokOnfIoiAn91RetNOFg50w8
j0fbI6hsjHDeIkR6JR75uiACZuHpz7okKourjt2fHYiYtOIGcU55W2Yuf5JDVfpt
q6ogC4snMWsMxDYx9B60sNLsb3KdRTmQV0qFLeYvr4aBJCjvdF5ooz8DLzQXdRXJ
pX+EC5+AsLFeJWubLF2si2gue133/B0JguzT6A0HrDoIM1e3NFjnLZ9nAQ8mXd+n
dZWC75denN8FzeSh9UWsdGd9/NoCucvLB1zGtRSRxZPa5qj0JEIS6f3NjnArEefm
a4KQytUFFsWIvjXu8kkVtIRF3eWkoH0kmK8uV2K//EIR1p5W2KDmzqrBg7jAVuvZ
A6edk9OJyru5F4SljzzYC+mU1kDc6e3zPc7rM0MPdjeRuRH8xF9IcL9NBMzEu1/G
LOYFi6BeQuwte0ZZmboXKkp+e2HYKCnWOgqfuNiQaU9/ILzqyhSvMjq3cg+tM4Qc
6+LYUCpwEKO5FgqU/m7okbMwaLjap5aLkjC7epo+MYxDS15GTd5OlpUowozY9zAl
iYrvpRq78J90vxfjW6LsnDikfPSLeRpRrRjJl4K7Cz3CUv+jLnQRy3T0ITbWYFoC
UALvhmO+MK/RhAQmCy1/ktc4q+jzc+li1qhQcc3vso670c9hFMfw/6NVcYCJUqLH
teiAVDa0Jlq20riX6STuLDk5LCGKqW36ek3ux7qgvIdKsZAnerTH8BakPhZXA3kU
A3xdXxHsyYTHcvQ/RtHQbX7dd1sBhKzODj/4Yj6AGRgLCQPQ/3GAxt501+yHorlX
9cij3ImVYQqBs26JSxk3A4mfryWvaJcRwvQkONHbUi6/zOSM5R4Y4KL/Uv7OKyuU
zWYujXsq98VMvsBo9ki3SSKjxXoq9gDxD4Xd6y7Zbwey2akoXWPWUhkFunesXr0J
UM5pO1RfmVOyzoOJjBCp+j+6R34oqchwpSm72xPNE4WMyvPUSRPXymuy14GrH5by
auoF7sfeuDylceT2Qch7HejCl54KqbHWaJ/PJ4Ua4vH8vcayViplAXC0epyhKCJU
AvQyveUYxi32ZKcUq8IDx1SQ40DdOHzDoeYEPoVoOoBowRXTlTsU9POf4eTg5Fsz
lO7l3MnnBJQoL3fzGuCYoTWB5nR+DxG2Gma59nlc6XCML8IvF5DG6iula8/tsnYl
RCukpACuEt3/8aWEU/eHF6WHm6VI9BjYywJswaT83bTYWdFsIUEdpAsKnvp/bVeD
EwAVNUHz6hNZnbmDC+QTzrQY9gXf4kG84H6GjYd6dz08YaEWf54PcVj5r5Ou4jHi
YbupzMq6bBYW7/byHSkl3gg1JyhMng4cGXOe1vrc4fZCupHieRYzkj4OZwY4bRuj
W4XhF7r6zrwwtDJPwVhlySm33Ke07qdvh1r9mIG5QDKH7Ouma9l7+zGOd76zzmla
3z8aCjlid22gAS/gI08F+F8Sn40Y00JXNutP4fJ7VRWrFS6XsjjER7i10LgbK2CF
ClzC8yxjUoXq/Vu9B6MSX+eZ3VB7qg1ujMeRfztO4MeFOxQxMBcpb6XZLwWrPrID
kFRBtXh3WZaXwOSPbdxfFnnHRFdUR/N+kz2dUAUpGLI08+r59bVAPURjzQ5+4woO
1cxGRu11B4cCrAAt6if1ybCmibXLwpy1pK1zyshRkaTzVl+lUH8vpsUBQOolbW1e
4/XOyHWj9XTU+i+zIrsuzGcLutl4XukH2JdpVB3JRqJiwt6oKDqFO5lCSFSNRTkw
/dmD0PNocRSjZziRfhwUFn90wJJDqb3Ofj1jAVv4afndYpFLRzvW8a88JjQjoJKM
T8IP5uAWR5dz2L2TL8lbPfVDrkNrcgR+UJKQxjeWnXSqtY5P9JT54zNA89EJRnnd
BPclvxn9fBpcY0JPPNlPMwvvnluhTGHgAt2z5rzEINV7vaRXcb9pbkWQEomXtVWi
sqakTzTfRCIeNvys8mAyUeDunDQ5N2LA/yAw5N8JpYUhbS/hySdGHkt7PGHChnI0
B4U/sFQg0uNxIbh/Ci4wwJ9MFXZiA59oZfvt9J22ts3eF2Ih6qbONvD7fMpYzOUD
V11bAJaz7d8slqX8zwem2i9IDz1j+oJQPyDdN9GOBC6fLHGKiLLk/NyP23NLbnEr
Rdn0yfMyoISMaROZwKC8zBdam3lgQFF2zLnN/yr9kAmbppEmk1LTyCsEFTqxXm0k
nVU3zs+SzYz7yOrP+PpEK/nRFWZzkvWzDW+l4V2M+BEhLECnRIUi0bOaJYNDGslZ
mWJO6oDJFCiYIH/S54vzn2uZLOglioLhsNt1+ZRUolT/4rHrN8pBoHeI6FlCeOtL
bjv6g41CqD8vxT23RXSyUElfGXD7YtfsfwNIeI0lwPoE/0J7ijvxRmiKDs6Xbsgz
1Qyx5aq7a3qO+vdpENc8RSPTu3jvS+7Yx809x8NvsvzmKKrpUQeHa50rpVvjFene
7LLxZqAUXA5KOfx1k3BFsAZ23luxZIqBYxAbSnSZiKtq4bAKyO9PxnzBV6b2RW8J
jbM+TRJcOYdrJjjcWIVMn1R+YmcUa4WROswfwBFuih0LxNASyt037Z5V6TpFJ0VO
M0lGa6rn2lCySqpZ9vX2gegZP19cxpqROLsXyTTH1DKeu+G8xL63P3OzYUiOLKv0
eY9tlGB79INqeIg5wmh0Xh8sy9C5A/gsEqViWwQGeXbUhQ69iizWdYbhs3ASkxdP
UEqFY+bqEPZyszHwc6cUj0j3zOEXXHyO2R9H4y3B+YgDjcF9FXZA2pgAB2HMbpBC
FUY2zG9Z6ttt5vlMUfjlkE7dUqKDpgaxR2UPoUZcdvOu8ZDIj4VIiDw8vgI+8VQr
pkyV3HuaTrp6WlazP/QqcqEBIa0z5+d20mQevy6oBTnGcuFXu8QdcDZK7S0L+VUb
n6ONm3frhjBsnN6SyoSSUePqlu2DMN9XVAIunAGzX+dqHIGn/EAnRomfE/murC70
g+8BEAsUgZ3X3Lw6/PUBqZWV47mgg3ZkxJiwGh26iGBkfGIzu9WA8v6NxlERNN+t
Menj60O2b1RtwczaUgjCwH28et6SWn6WDJDItOSW6G6XoR2nlGPF4v2DFUyAsQQ2
ygC1pM3at24HP88yw56qpwtkT6q6OycYooJX7RSkMEHkvwZp0RG48Zgw1wh0kwTF
oPcgr3Irp7w3oVA4fMWAX8W+Mzj24HXPIEpxLw3IjYrar3yHR1tvZ+Cqtj6n+Ku1
0dgc/5bYYSca2+e2uTZcRDE5vmPu4HUZKgHn9UNGfsFWK0w3FFeSnhSHl3UKgH1O
TbYAG1M6JxeuO2hJv7hDf5GHiXs5fBD3jYUcgAx6Liz7I+pSkvFtCanPCrHrtv7c
qCHJ5k5Bcq/GDnCO5BUH0L2nGt+SX4G3aaE802CTk8JoaivLxvjE4jb1WUWpjq3C
69MvWdBnCasvwn6H6WzE/dRTtzlagV3U74vzbpN2AXS060p5rWLNj0RgvSRmfOTa
+hGHp+AvYcTwSboi+gZy4oL4LiSEMvyIzeKU7x/HjMpKgkAWEVS9XYaGyxAZ3v2x
Il2haMU5tSBMGmo/5qWqx6o0b6sL3UFBBrxAk/PbnrBeqnf5OVRsayxrwIiBT/M9
9KXiLqhxjCG6k6z1J8Ein/pfy0wfzsat3v7rXbYTHmIOEzvJvkrBD39WZxxjHM2L
UsC+abM6n09J3NpYTQUNJYT7TV5YFnqeR3NLfuj51QH+kRNU/5fgbRsfVYFnkX64
2Z9ogqF2yiZvJTOI7B0vQ9WcMAUxt5ONyMs3/p8xC8W0BSQ0Tqn3GCumwqEmg8ZC
/ux96UJ0uyJkX0viL8CPciUnrYIfru7YDvvKdY+228zZmkSII0yJjrr5f68D0e7n
7g1b4DDY13u9ihxjBnXIwnH8trhb/KkXhKRX8DKgEhWpbmXxSeP6wskIQ+B5YuEe
j60YWz08yM22fgu82QWBMdwDlUCHWvjxZudWx2lnB33g4SCpiBIGomgf7/PFCCoe
W4NPexti/RoB9pk1EEJ1T2ZtRxY8u5X/4FVMWDQyCRY+CSBSX1PJhBtVTyFNssCw
4TuKaGpR3lqRmwArJx+1a4RqinHAlWKDTqNXUaN27aaGv3NoF6XtI+La2KK2DSeX
o7JA3PCGJyMMfRqu4q6Qz09pxVzefp8bihihGpnltQFdWWGS9u+YvpH/szmjj7OU
4LIZ2Dszy6Vna9nTNv514XF3TsUGyaTKlv4ihLK0ijMsHV9uIw0p93/DtsEdqn70
JkBGdP7Jp9tGa0WfhIj0a3O+rCj76dvCo0ixkhBsIkwxJ0NiDvET8LjJplsrmwbs
Uv2Jzal23MkaD/R7LMEfiHgP3wiqTeYrhUhEvNdJen5cJaL0gW47Z8ybLJorpktU
73CsQeZ/K+LrylF6lGYsoHxWT+O4HRPk+GxIjxHgkrUcDkkA49iuWqtkIfRX5Gba
fR/jMuhU4S3NQQoC9oqtPxZzjwUdZRYjnUeu3BVNZus4vs2YIYrC7KhhQYTgKEqk
l6JXksn1SCBCx57CraOGk5lb1uh2+DVDiCgFZ3I9FyIZVxkYlFlNOFacAnGGiuO2
y6otDW1pwmYVtNSAMwXCWcC8opholyRYCkZ9GufjUwHxRV3kZapHLRRcEcSj5dEe
hK+KOjCzAUDs+szncACvPd1bU4YRpZbB+6C9fccpKCrSj1ZQHYDBtq/mg06y7Ld+
PxyCD9apD0fyoM7HJDOKDg6xgeoU3Iv+FipvuFq6u6kGdoeQR8AQ0rmysJahkaVC
ETZYAuWtm67q+eWjWCUK1FqydyG5heYyOaeVAKeafeETG6uFZAtHVCAl9vtt+T8u
5LU1snBn9X4Ykrz3o8QdYG/JRqhwZningEDqCpiqmrfeq12UP/sIhu7bR3cE6HP/
jk1IdtDFRHcgkeAp3WacIQq6s4Q3T9oglBS0x+mOq2KLFHDICnTz6vkLXV68fwAI
WueekcyqisB3MOXNToM8o9o+vm+mcORS988030KB1Qif0Iaq4XpivG++G0MX+pd6
cofmxnKQmgMQ+bIuccp3BVZqjvJNUWXGL/d8RbeHP2tI+9CRPRz2wZ8yWOccxpZk
Ulksr3a7ky0h2jbh5I1IEdwApAdU+ikSgIX2JPCZwVNGhOKejDl/tWy3uSX9uNDx
ulXCZa3sYyj3qIt0B3hDXfNko4XwmcrmlebDgzpd0Wkbh2OwZAF/91zJw5FAoYyX
W5wPrMYPbIsscFYnmQU87zRqAMGQ+r94mb74ZTLZAGQJ0kbXepdA6hfXF8uJVIdH
/2usQIXMXLnysTM436jwPDkOcrVX2VbAekOdRvETEAg3bkYCllyZ6rIkVIAJDNtR
+xINm+88v9VtMhWm16rnXEg/t9Ja+/PEiOPzql3cTe05uMhDYZM3pajPDnx9x4fi
KolkeNkkL31WyKmo2AgAlxRb6P82xHn9ZZgwpGF6x04kmSbZxFQ0DGiukYLbnbb/
cmg5M29NgRTYawbM73UBzuMj32wHtC5+wlixZ4uzVO+ht65um3e4P4hDoFzvrsO0
SSA00HBIVarNpVlz2nM6iwGFTQyoGLAfYP3q04gAQw/FGPpzxJGaRtd0g0pkQWhi
MI2ndVhrHChki0AABCZaX3VK+OFVOyJf46J3Muz4wM/HvwHYFXXUfkMNNESyyDsA
qJfED8Wdhq7eoDMkN80D8j2cslCvS7LqnJOS3h47nMDgcCkJ0CtFLPFHIvVF4uHm
4Iyfi9TjsXIkqbF5hAbYi56ahOw9r/92eLZNqusWTE/bJi6xaI6/nsWpFMWiFDb1
cLRUZEIc2hreE46t++eUDVu5CerMpnhLBOQ5+pss1nHEZegsGLaMprhC0cOGv5A/
fr89RRrr4T+Z0FVPVd+njw==
`protect END_PROTECTED
