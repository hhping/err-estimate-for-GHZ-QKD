`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FiepKSVvr8mfylcmutkZwdREsmXPbLuaGqcPFszyJ2BO/GS+1NTcx53QPEhvhAwx
RckS52qv77hz/4eiZDRM7mmWRfCLgZCdPRMQkwBYTegq7igTiA8iVbBqdfsyLWfN
huiKC/xvMf1vdf2YifuXc+eQfkY0R7IdwJ7TM7iCeWIp8liMIz8TiKvaR8yCIT6N
HVuX5M57jBlZcopvrMFEBzqaCWRcQhsG6CsFX92LhTx92PcdqCc8j5O5J5SHCsU+
bBVxZOrEWevSMTtexHu5F5tDuVs2WzbQlOwBs1soVQHlmAhg9jT3dZCtJ4J5rb8U
BJwpEw2SKDTG+j4Y5GvZxxQH9mPyyspLf/IV7zlFRis0RFtVsmFgB/Zakr10LHgl
eTYHXp8gIzEvkDWRMIFd8FnHDQOU4uoI344Jg+AdmDwoScQLOEjz66iRouTkOsEI
+lMFNc6rXukj86b8TaLMmpyilOJ4jR6Ho7YMT9Vc/guHJqltyycBubOA4Uec043y
PEg7KsSK2oyS3ASep45J4G2Vwsm1HyoeBpM55I8YwiajoLT0rtHtVWdOLM/9bcPo
6DuTe7ufEHrA/0RttDGbKTk1Nmq6kW1Ax/Q7kh4ubXMJ6xOdBfxCi/G6+2GwTf4z
n6ppgB4eVBVM5ct7vwdrpjI8SdgfP1CaxbHjsgm2tNeYIOQWeUBgTI96Blt194DI
5WcRMuoCBYDVcCFnC+PeIsonTRIP655TPvjEom0sieTNb6I7lVEPHg9izV4LXA1M
6vuIqsiHAotBMET8T3dSlgqckVcVnj7rbRDw2DIyXz792WJuOlvx8Xa8mYukAWTk
lCQaOFWuZBTepXDtu2gbRfYZYZeG7I1fowkwGMruKIA=
`protect END_PROTECTED
