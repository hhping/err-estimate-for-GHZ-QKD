`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K602TXYziXP+vPGDhmlDbiEyO34y+AJNwFqj3ryljkeuZXWXElBhLmE1OztVpVpW
mjYBFj0Z+K1SNfrHVK2Px2wTAdloKzLtpgy/ut7kIpCqelUUZPTNpJVK/9zlQILQ
8HloT113FTwUiB/PhiRWbYwngx2LMbm/tRO9KxQbhEpLC/IpZGkqVep2FmXmIYP4
Wl89ifGKgaITXtTxYXJiyU1osl310DlTnBcOSK/t68wphk/9g67pEaPZVhJnI7c9
jdvy8hnZa95cFWpaab6ymRU/3yy7rHLdjMi5Ln5fQHvpYgCricYcJU6j1tMnrGag
`protect END_PROTECTED
