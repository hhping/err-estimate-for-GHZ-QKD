`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
45jlUHCB5Bf+NLs1yJIBIgV8yCz1qOIhNdBtVzkqpti02SnBJjMfr/UmsECrQQ8T
XOuEMhurWyXP5Hx3DAr7zHECyHRunolAuWRdFUDKlLVaMdfal1h/39f+2+iNkkSf
gEEDAUsu+g4UbpXlG30tMtfc6xk6wbVbyepFOxI5EX6TiB29Ee+hN8yUtZc6L/lq
PPc5tOQShPnrhVtxFNpx0lxcCnMDiP9BIKZApR1RVpHLwUpQR+LyuF3CIooj7u/a
AD5TBxzZcSVd1CXJaiQHkT3Xz1yhbsOPQWN2nxEl5Uk=
`protect END_PROTECTED
