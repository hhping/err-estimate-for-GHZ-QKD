`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LL4oIPwdQiJMzgQo83DBUf3xMzpJyRgkiKeLtM5pI9PaOxunuTXIIIoVtxXmj7tr
6r1DumTu4I8/idj1cGrNvoB5X9/S5M0MXHb6sEhtH3TcGL8GU3J11LcOT018Ta7O
zekpDn8KXrVu08rTuAEK7xKdyARWZeU8jihM1Tsi4qxVUqs9N4wHj/ML0zWes1/L
TaIKyXWJY+dSrv4RnSJVc1i5XAznhTwFf+8Gl8XUJwMbL2SHrFyn75MNHyTQ9yN4
sUapORlvVRlA2BLr+Aq00UlJparc5uVhoo1CX623DDz8JsOn3HbGfMKzv4WHF0ru
Rwjfda1JzX01hA9eBuE/CKfT7w+sfLS510t88os0i/MIPKM65Wwy+s7JE5/wWo1B
kku8SDIJqOnbVooY+aV9ZIQ2zq61e2flCzuKh1bo22HtDPQ1n4+7JKWdqEu3yeOm
2YVGEZ4Xy2K4K/Sfr9G7dSDocnHmhSXq9ACnlz0m3lsohsSjCfo5ZseY9xq4Y+Ga
H8lbnx3v9Aa62sUAA0EIHt36pV4IuraQt3wJ/LOylPzRmpUp1NrU2jshSplIhY9C
mfwHyjnYZp1rQpC5ngVmnJjCTgwVbhMql+T9h+fug4jHcEKel1Ih+50lPQH3QCAR
JWV+sqMK8H4wv82xzW1+NhiiYMPErP++nCOsbZjUmiflPWTkHapYGyTwkpd4wgu3
euMNV4oYZTL3c+uvxb5mCqcba2vbEGG4JJQ9SQpaQD2rcQySGZG8/2azkQYKFQIs
5EeyX9w6aF6lFflDhIyoytNspEbY8qbI1J7FL9yLMlTDL1X0wv39PIqmcLNUsxp9
/cQN6l0Ente39tCYMxlt8rFKCXb7RzAUy2BSQr8pKgGyhmNgJ4z9MhdfBr0vopA2
+xwXK/yPyrs1/eEjqArLZValZI0IXpxTghteRkFK3iKaYy9cuZ4adFeyyJA0+b5K
CL+BUWv58ss9mwrneusf/KFf201xu3sopux3Gh3g4xbMXGqzDlvX3vK9QVz9OVZY
Hsz8onYw5cvCBmexUsjA+j4U2KGt892YcZp3TXyXh+IJ/YenY3sklUiRVgNB2a5L
kufvuPPTZbCdMBJEmkouZl7GM0Ieck3jeppeBezmp3u29UM/0ONfh9hohBP2X38E
Acv01Cq34u+LX3VSsKFCS4de4f07EeUS7SSMDQByc5XHzSdR18q1NeoaPp7o6eBm
6HsIF70Sphv09VlgeTb8g6m1EDIB6oH8RLrKPwJX7w/seoU1uv2nXiRImS2c2pVv
`protect END_PROTECTED
