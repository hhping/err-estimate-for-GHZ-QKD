`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lHryuvfTi1nVbxs+QfysuSXtb2a439o0FHe+9nWykZ5eo5DDwzxnRfCDus6pq/4q
x2U1FBWv2O/yjvIFmtMu/9BxDLHTBL8jrpm1KeF+2v+M2VG+dK4bAbxB9I2M0rkH
aZn0YSkMVdjLFX3F//l6rwtR6jSoabjN4a1WEbuVWQupNIyigW6a1K9boBU1tAvQ
MMQcLfXcox5rEdZc0gSrxRuqobY1+I+6ygRGORhJjIbeq33cmLAahE2g2jhvR3bK
NyAHrhm4GHszb/uBEygb4JeZ6WI7Wg8VoRXzNY3REFsPTzul4MS1hb7XQ4c3Quze
VqsU5HZXPn+lqNTi3KM10/WvM1VZiyEJCg0BHCMTeIQ+zfNE9Q8ooSpSL3uK0L82
xYNI/a7mw6ezLYrl/PErjg50PYV+IxG2ybYrzgMOl1QyvDtTm+eC3NfP+Bkze7gf
6JNR5ZqbgofadMp6hR5wF8cJ2X8GYekETKp6/84S8JE2jpLA1VsWAngSbcAHXcGi
hJXVQmWTqWH2SYVIhyrg/xj5DU6+0XcHCvOBjvYl17KRokk6EZL5PHOJTjeP9iB9
Nto7nbbKOyniN44Um0gIVKf3SUtfpKBwLFvNwonYOxlw7JdyAuvl2JhNM1wVwlZu
boxPob890x70PsGIDeL+kJ8JzK4HiAEO/KRZ+W+JOE8MjHnut804bflo5Yz3qGUR
nSK/1UA4QGwNMqq9uLy6elBgcv6TqAs4zyqfFmJmaxhlHccHpLPYm0ornJXm29So
MLJ2E6T5ybh5o5UP1hm4ux9s2G02bo+lBZMY2tstiPgbW8zXQt6Qqk/UDW+Wdu4M
mBk3I3WDgVeFkjSa+XkrvGoLREsiCdComwXOcCL644R69sEXpXrCwD7ZiYAiFxrX
`protect END_PROTECTED
