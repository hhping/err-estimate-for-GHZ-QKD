`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPA/xFT7wEO6CAYGtTYOrDxrewJM4ruDssjfRezQtlWSHyPtI5IDtXJ524U4IFjs
M9+kPbGtY+WC7K6uu7PDDj4DHj5JXOvf9lbLmD5drkad5wM/y3KNg54Av3olBIHm
TUey0xmGTUvm6pUduAhktZmmqzrjfkWACBOquxgMgVgy/YiASMNRFDbN4Y2rL1ZM
FrutNfwcuad0xbvsH6hTGySHo7iS0RBTlZAx2Al4S00Nz5RzhO4Gzes6Dg+m5PoG
X1Dra0f6bhbNUkq4GlL7e5UJvaXmZR24NU09RLRQcu5AMXnoAZD9DdSpORNRClRf
owaPMJa7ZL3EdkBILmDq+kxzDUYY8jkousxvmQlyWEYglwGjHO7hKQ/HBedJi+q7
KhiWmcH5InoRSpabwgLYF4Rs62l5BKAdoubX9Ef+kIxVXQw4BhUiTDk3QpcIExOS
AYLO7b6fFl0vhWVzRx+bzwSZM5/bf4DC6iEhAo0OhizzTWets1rLRkH9W7dBzZT2
8+FSEjHBDCKHfv3bfOXJelWpuaRRNdR8Jzk2IJbUMJpe2xcmfIQ9l4jG99zNi+e2
9YIRH30JmWVCHM9B/l+acefVEgjTPNNrK/DotXAUvyCzDDlfZyqNT/tfyIDll2g1
`protect END_PROTECTED
