`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S1onC+VEGw8egYlhn7GRzFJPWjiyEllCxhYUnK/DF7g0oQqn7m5AB+YpbZ4+JZ9E
saZ2tZbttKAup+vz+7UDX/k4N2d2PLrjWXd1FuhAD7i7sB0nRKVauap+Pb0So+Sv
1jgUBiaLuPEZq87BdxyHv29ZYgAwwwczGzIba7GZgqdrVmZQ8om1vl9t5PeCXuD+
rLMlo+B/ZWn7qFY3tOtz4tCVDsRUw64WxUqAsLr6PKy/eDsYbFQyjD56DcwTFbae
E5emJVylKcYKsdO7Mxg7Zqwo8lY6ZruIE4VS8vC6XUErEMPuSG/Am4zb6OIlVvFP
7f+UWekEvgKG0skueuPjU5ediPwOg88j2/CsqD41Sz7AdClllTcYrVUwiX1/g3bh
y3XFeq2D2kbqHeEsA0iGXHepBi3pYIpiPfX/5iYgCN/3UT91HDCs2BuZXRrLfSgo
ND5ZVsKI4SgED67OJFXZy4i8z1C4Lpq3OInicDz763QJWp7/FcinKIMi9i+ZuRHC
ermFpsKbFqdNPtqzEaFaV1ehfj8BS9ajg/I1NloEteIBlJUMqGfLUp44qwGrOOkO
OgKPKcXlxxUynPt+ISd8S6351BLbv9oVQNrTIX5SwsDy1n83pRGG3tIoQQhSQxUt
4qzK1Ro+zEkgBK8iRHAk2jLJCQ/zD7z1ZD8bt0Qkf/97ZSyA+RCeRgJTw+DhcZev
xkpStKC93WeGR20pS1iR5nLlpWu3+01SZylowNlsdwOtGCSvJ2hpJU69v3UhHHo2
Es0pPS7I6kTRC8LDBaoWmmocRlmomXadJeVOSWqBsX8XnTgYWQUlOpjUn0H4Y5qs
4OkyYTIvTYufSfNhN6+Io3o8FNi4zKATxBcbe+5yAAUkHME3aE4/3dMAVnJFgKHE
neLBomrt3xtfqbDU6kxLVS1HLgZS6nmihlQ7EQrpGLpHLKLLB1+5AneVMhqrrHTl
DqnqOuWrGH3J6/hfmi9oqBKJi00sxXev+b2izDOttZ6lfIPvZihdzKt24ANzjTQO
+qnMB43lryGNBIXggsUSN4RwmdTi6Zyy7HYUHTBWcGBvnoVC1h2Sdx/5XekZqYJ4
sLOrQxtXLIvXyqu98usaTTaHk5K4lfU1e/Jzvitn7MVpjRQ6x0ANRXLqCEIipMfu
sBe1bvtQ7FNGolME8XcT4KReEmLLRw58h7PYjvUhEezQJPgCXAHWxouPjwGknrjL
L5/sOaBasSfIvnWC74G3nmgDCy47/gTbq07H49kYRDlBzmp632Eh7nCEPJ9muHc7
hulWSB1EqkBFPKnPAqW8SVmheY+VwQUnfIWHLho6cOTAh1QYJ0IRqzakKk4Dqfmo
V+9I+jlaX+lxGCIxh7NZ42Ti3XQvMjbUpD908MmDKdl1tLjwL0jmcOnN7fgRPram
jBWsEVjzMBIp9zkHZe2sf6df4V5kyqRmapRLzuNrWEAukFE78LBecHnG2wXMPXrg
xm6bn2sE9nXWnUCijsq55NI8u8iSnA8DCRlYEimMgDZf2eHDTnsx+U4D9V7rl9vE
HC8XY7ouk0J8k7lUye4f/w4rU7NPmDWmYPVPUT8FHuru6eSV+oEc8Og7oWIU0BIm
qoYtLLgTWsVzWHn0M3SxmyKyIN9w3xFjnF0VVom+Zq5rbOd/jsYe9MiO+2FP8fqj
bFlvT+8XzhrWrZ2IwZTxF+3bc7GXhkgtzq8gX3oVKOfH+U9Pwojq8poByckFXgwX
Tpy6+osQw/Apudc976sD6//BWqF3f60hJgPDsw4gj3mdbyq0A260YDXAvdGXPi95
8RxBlDelu0kHujmBjo4AAp7vsfZv1HNBXoTzi8TdUJvG7+m8RQHjT+EZVIqbojyv
ByBQLbvwt9yJn/fE0rsfNDlrMJXrXNoRTM7dVUa9lnVclNw5gosVNjHIOcd6vQFV
buEwXEacYYK9xqTRVf6qeZSFxCX1+zEQvqptHdtBt8ud56oe89FfsVdHuXiiwPOs
a5SMiL1Z3Zvxx+Jrj8f8TF6GtMnzsGkfGySR8L7jzgbibvQhYZZfJy8fIjKpEhyW
03bNsC9v1WLhYrCfv2zE4SpLOOIDJclMctcLVAl9Zy9XD/GpDb9tLnF1yUyKX2TR
tq3+W5APscM9oCbW7JG75FyhiyAokR62phs2micd74EI/LIlptSS8mqLlooaKuKO
iy/P7kEsITVF5OzGO3J+QBJoWhB1XXI1L5JUFAbR3koP+6tKT8x9+p0rEO0JgH6l
/rQPqy80pDJNFsrM0PV0Wg==
`protect END_PROTECTED
