`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QaWM72Z8WE1hip9nLXJRRMZdSk8rEJaLaE+DkMBbK+FjgQXUPXN0M6GJiLYp9tJW
TplJeJbKWoL14CWk/hSytGXy70rKrXP629ATBEmB68lpDGWX2/JVktw+ltPNbZ1a
dJMGqvHxCB7vPJCP91sFWN2k/UYxZq/UFxcvkelxCqLvql7wSw8LO+e3vQr1bwMk
pjyitWsPqBGdZt3nfk0ta8DeQ0mrbGncJ50qW0W0mM9h1zBPvtAUB6wOOz9WbKCN
5UzKeK6GNXMmCA63rCUWWdBk3vqFrVrtiLOlqQ4bGqxVS64XEaWiW5/o2SG/iKG4
GgfKy6mnybZvZoCY23briApAQaYXGvZpEMiXZptFAYwz5kFBEQ3k81bIMJUjAEyM
G09BQ3IYVztXvzBkE654WJDXSQUsXLCT4PnDWNUHcE7Y4rZuhq5P6laLAwIbvkTY
2c+cYWFtdcpft2eB35H2BbTZmeEHerN+PCyAL3eSW/PLzcYmYPigGkzxGzgVkty9
tp6q1Sg+1h2Iyj69URsv48aMlPj2cBDI5Ccus+n5oM+NoaPclNVz7xfcQLBm9H/Z
C5sjOTIu+r9D63+a1abEUV8LxzKOhqpl4ZzNq9EZLkTPSXuvym+hktCjCIEGHxrQ
trBLfYHqL7cOm8KQ1hclSVGlFIIn+t7IaqD8A0y/WINh18Vb6aNwqxfkh69ZkDp+
/xTH4WLc/FevxXGoLghxGSkd/41YbyMDumBWymdm4RjsOxshFAcLGf4RXWPcYGZ7
IWRDfhOwhSVd1isZTGhu1Dubgpft10/xoOFh7Y5O/LLX67C+Zi55prsyAQXfdWco
Q3Z60H+wlFvuu8eJHkRp5CefeEFqs2eBtYcqj0O5qLJZ5ovDsQpAZaiDbzPeGrgi
+Fg6Nju4CkdZM0Lg0UVm641wz6LrDfpF20D/QTD9ILq/YpmquslAIoKJqjiPm8Xh
G0C3VQU9HME/ytnYXOsGxtwnZEb2aqLqz07IFrTng+rzQdSDqWY7Tb0k38Z1DP9H
2q6tB+bPa9iu7SJOh2Zk/3fKm2JTjAMyiIx2oZjo3j8Ggm8PoVVqA4EExCLyo/gm
jn0Thda7KJf62/iCJ4zdizLjBvU+TmRkIhuMH1+QKNvYctP7aL0mvH+V0DUx/75T
xeUzWuSlek9IBILQ/7sveIRjnxKyf/YrerAqW5a//gMyr7QBdtTQ/lqmbsxB1aNA
jkIDzYYhZwp6rVayvsLpqLY20t36GuuGpAxAG07ypRANOboR3wwfpceret8uHNOk
X3StgzoiY911gQ9jVjB5ISQrsCyhc1e2YXyy3rDKeRjTh8XU8VG81B8so4KJSPtB
jMo+plcnoRAddpxzL5op8RMMGR0aYCgMH4ncb3eZh3kFn+xW8s/nOcbq67Igt4iX
wfaR64fcwivC/6yeNYVNZdy3zhuIUUCyQHYdmNdZ1Saa28iq20XeWvrHJLM3AV3t
FzhaLUGiHmisas2Exxk5uiAN5Cg6n+PtvIAoEB5cYM18ZDvgfqwBI0Ul/wpsEJnu
ar6xkyE/GoQOls1Jb2zz8khHE96HU6Zq6y6JdZdwbkZI8uapCMgLJPiowq40l8Vg
DVFwm5ql3fAeL5ugcfgrt9D1b+7jFdfKhEq6Top3NcEbzaSofWMSCY3mO6afHNFG
kn3R+g2Lbv7RKe+ErF/AXyV2pEOriFF71NmLczRy0j4JQlg2L/GTAsLmmlMblnfY
JkHMAVoHpI2UBIPO52PpWxtQJAhSI8XSZlw3rcDvMWxMn67Uv3jQNzrb1yZ5JZ8W
rK8cl4+y+udeZHFdZpOt8ZgidImJNkMJ0NcR1arbvJ12TGgOjHISQkHnR7LRFiKZ
n/J3y0MQkazzSKDm3BCYbvIbNvDLmaPbXPvQuBZfnOOKWAudF1RndApcIFVREB66
Sg6qGQ2wrCMj+KdtO2CuvNLkYoSMEKsDjKM/V/eh1pHEpp2+qXO7kdSxpBPnBwmc
YUAVKoo+JbvZlWDB4T1gkaaUZetBaZC3Q/eY2YeGS9FgiPvRcqEiTBqwiTf3vsyL
ZqysPnWR3vS02tPYDW5Xt4Frvzz+pXaNlzKgX6sjtJgtkWCOeIY7Nmh0gjF1WtOo
`protect END_PROTECTED
