`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJHZQABdA9p5VpYJQuRe66ZWAoVQKiQmmviwfIpjENVbJRvQtppdL0Ba9/wTYe8i
ZFznoFXm6U21Cm9y2JJDyPHUPhxZyFSNr/uL+alYBI5LxVgVy4fxxxh7NQNCQz6o
R90MtbRkzoiqk2/oHMN++Ddgf94D2PJ+EvDtAPbZIRoSw2peS70xpNzB+/Qgi9tf
tWqS5ZpP834CbP04ld9y/NuIsjQ+2w8Rx3iZGbARaamOQ37dgUFvjEtw5gH+3kRZ
ubndo6E/JVm3+nY5HEnl88lo3YI7eIzGFDvARZu7+JsdJgdt08qL2ghxiKJdQsdv
xewYwswuopbkpVPkTVMsCSYYznAmLu7NzAsmckC93FXyi5WmyPT1QQ6MLpo4mMd6
5aQTTcTfV4XY1EhsUBORwDyKc6D/n5YiuJ8KXpqAcK12H4EuWnSNl29U9MMiLZOo
h58DzWQJIlOmdtRcJeGmyPILHHPXsOAoZZAAWJAo467k15fdv6okuW/8q/emCw8Q
vDXPuRs7jxPyQSACY/onuxvof3orxgrjihoowBIygTMiY/IACCmk6CBYu1zAqtpm
ZKEC6rKWTkfiiRDJHtTVdFzJIlztjPUnB11cy2s+vbVC5AuVP3ULIrshs1Wuddyg
GWNLmkIspKXetjjPDO5/cHGFbOZT4HvjWlIIlOaVRuhohxXRWUBQTVL7kbJssJDc
/YT0Y9gJcuXufND6NjJujB7+BOMGxtsBEY0gsGIEzARNjoO2WlWAXx27sMORH6ed
ud2aAnpKVcXoNFT9Xj5SMfSxSzaF+Q8XSp7EAYty4pp20AbzXWHawrt2k+4AStPZ
60q4ZEXXauleKOChP1EQOthnh1pZokCWyRdMMUcQk7+lrW2n9crX9mtLajxYiIEa
7LJCi4epMw9gsBczbSR2tYhcNSn6LBJl5Z6n0D0ebWr1clbcnQlkFAJLZvJD+nbi
kiD+uoG9FurLCt61VUIC52k52OtfwE0zF+/fEco8SkEBi2A8vq1C9kqDsLX/fCxq
BJbyQ7tyBhtg4HrZFmMvvgFZDg2OzWP5df3zpoEoVgI6Xw0fR9mZJBEpnD2Nns0H
WL83vgE/1INwo405DGUzNrZ7wvNWpVZDnBYFbMvZhcn8R9Yj14NheE2NEAay3y/R
l0Na/ua9TbUj49U48fg2fDBEILmQbrFPuaSuTLkcimO2cK06IZgcHNhULyQ5VM8f
ilVj1YQZRzuwpPa95Nhv8Nn4n8H1eTv+rPAc0kGJb7+jax6qv7qH2HbH9ychA3Uu
J8cofkDe+5vqjUB3wKCgMZ29RA8hRVMObYJ06xrwIBKTRi7BKit+BZMKf6FTQWAJ
UZs6YWFAAzErIKsbVJpfYABTk/dl9QYUsEbwjx16O9g4/N+YcJEIffU/3DbFci57
ktxJFDDeBKfuxmq4sTOn8lI1VKzaNARtI/xkXBEV7f85N8iXubqPwGlCzDOu0+b4
a2lqBeKXCQlvArd61X2bI+aj/+ANqjjGttaLwahIZ5s2+ji/zW/ilmEbjz5AyTq+
y+sTtYv/SA5IfqomaXCrOwsOUS2akV0gAe2mnOwnojYUMN3x+OEpOU4wHvzB9Dd0
Sk9ixH23yIlCaF3iG137BfrJkoFZ+5+4A5LcXGtytPa6mdIE0k/6R/BmFF3kl/cj
f/JVYFmuJ8eaVIHhmji6B2S1R2CnTU+//tNiCaDSCoTE+iMnwz8mDxmnyEhjnynT
dMqe0qLtQZqaul0eGiNBRjOdmeeFy8KNZrhoJX/O5oJMucLeYNYux8+a8QsywrbW
UMd9kZpiMkMt+3P2Acna9OXzss6D5eHHzXsW8mZmINR0oqHiVa1uyhyItdm90ATn
NT7q/pRg2HKtH7MEWEnF2MmlU6y7byo0IAXZtVV9OXDl1tSG1VH2n8mL+PyYOBG/
NM5VRNXwq5FQxsqVlltf0buNABBHTu3N/URWnDgVuDhbPG1owrU4bR6/blHW5NlL
0f4kTilBP+nKwIxwVdGvmKI8FjHXFInc16H2EoukQq390THbOmZlZ9jShGpUKgSA
DWuTWOSomxTVV/+bAyXzP3MM+vf+K8ptdFtHEtNIw/4MMWX5NNQjhWRsv30XnQei
9oPvzHrzPlcQQw1UndD3yz0hdclwtasmUJoDkjp85deRTrutFKzcd5EJzuWe1/RO
JLGTjk+fzHskyXewIvdyzbtStLk/LVUko3+nwn1LmoEDivFhQHeVIZ1kOseB44g8
AYNWMUWbR7RT8/gKexaTXNgarN4SfjF6zRt3aFuq8vzlBkz9RGoVDBivzXxbmDSr
Z1B1H9yS3RUOOaUD0ESfjJGVoRqCaLOGBgLdMPLSgKz8YL4QZWkIG0Tn3deRbiYo
TV60tiNuNhQFXnoggm50AZkIsUVHnlATBc3hCZiXOxqs1SoyvZN5Ruvj3gn3ePMZ
IlZNVffBxVPK4VQ5dtVFMwTalxFMJCJ7+nRmt9t6IK6/fe2qhZi9aGIh7C78WHcC
T/M7/j649aKWsggumhuDmlQCG8hHZsKmUGE0y9Psd3zmsa2kTIrYIu9xjyLrLGDN
9ZlQyfVgMLlrZMlioVlQ1TKLntlD9j60Vgkp1IFyTLbR/CMHMgVwPqmh+wYRTGDb
JjW2G1Dg/ILcxyAJsu+qizmNZUU4cFD/j2MNBkFIw69aKOOnut8uG8RAGIh9nq08
gY/WPOBVGADj0Mk4ofbCuzBehzC5R9WaVwkYy0zNHGNxunc3Wxo+g/g9a3sKIhRC
fhRmQ26we2lsw9x82I8NfSlGEVLu+jHh2szAGTS9miRwAFrDioCGXPgn3KHn5HC8
NsWti39a5VgNCfSdB85UQdd/UqyaN70RWm7gRWei4JY4aLspHdBND7Sn+FrqiEeR
dy7aBUwHDRgJVHg9/Nfwieo+nNrub95OHAWPH6lW2GY0f2h//ypI15i0hHheEInX
28B7L7XZdlcQKBKKT7/biHGgud9UVs2t9eNOS854dw2Lakr3Yc5+jCSi0kwiLRFZ
PRtVbnke93V99AyEJ5PEV5DEOZxgffrnDZaPRJyh86jREQkCAEXL+VecMjVfrG+6
U9omyFECtP5hV+mZYORiXjXdE+okKLd5nm3gjx0tFTDhlnwhMcrWNwfxRiczBCWU
JTM5VT71JEh6srm/3ID0D+I4jIaViyCi7TX5lXURLAMZ7pWnR45R/9QD8E3n0FJi
r+lN+g5lYeMnSpr/gkMbCpNU3DTdcw1UgNN+Bf/ruM6RtzKKCaBLUo8SB55gOGDS
qNzdC+ys2Ohus2ASPG6WK2Ve6TZD8XEtcEaTPa0yfSc5F5VQMMy4ftasRJjn0mMQ
gliceI7bZALOkF67Nqpx/rZ1yYCeLlDup6e48vO+2MFp7DhOrbY6Gf7uTGWWrXiF
kK4jtSHj3inQw8Rg89w3T2zgMCfMWiIUjxYPVvTIzG6DoS01KXBnqccaDdEGdhtw
6aMDErLvt+5USM7drqaX4soEi77xTm+KvPIjA9OjEbNpk3DV7jROml4RAKck2mm8
24tyFg6RrEfASm+xF1BUE6GvJQ5iYnkKFvIg299Ld33sxA/GMV2qiRNDR/lwY0kj
2vE2gtLHKoeeZ/Bf9pc2Kv7K1ApzKX7Bbsdxq+NN2bcjsjVbPMhxm8YTpFYcvBeZ
K55GE/8+1ZK7oA4ytKqCwZH582BZVVS6Q2IybwHU9LwdCxFwnbV70WCLKzeIAlj9
+OPPOdAPt2u3mlatUk/i4gzqW7ruDdYVVlXWUPoT3T3tqRSH64kJs3rMMhg1ZHz5
7kqi+Q4VCdnANyWzkGXXp01QhGi7uSOjKJn+mvWtsctSjJAAxz0I8UHx5cr8PfQT
JZRpNVWhO+amw1rmqaMIUe0NnXUZMRMu1Av8v+NP1Ev7GvmXxfdSNuWTHlN1bAqm
SbYvFn2zaatvdasp1QEgu0NwUrvXFLxJ2fLwYxHJrSA4R3FSXsFAfs697cJ4/jeu
bv/i3FcHn+N6i/utDbjUOn+94rlEOnC3SJfNvve55SgKg2HKXUlV/jg2v68DBs2R
pb5dvsxTB6v+xbvOqoYk7yjmUic1gYFQ17+2WZ0DhIAPrhcq2VEh5/9nMjtL8Y18
i9E2npez7VRE+2Nd2bJz+LDeToLrAFXu96uP2yyLnV3S75CWpFwSwTkiXcpxkmwn
mEnHxpaTH7+dr051DUmq8ykhowSoeTjikAo33RpPMas/eSb4LDVv3AYKQ0UkX4j1
84qiUlsNXQ7Os7Fw6ukQMf6vvYjcVoM1A9em7BbLXoe4ORl1aX19Eizjqiqcd+go
kCsFLqfUflers1XCj487dkxbndgZufJbrBKLFIXvPLtL6BsVA0NGmtmk8LcNdrM5
BwjguBmVrxEr2BppNyKPNuUYfllFvo5mPePKt1/AiD+NY+6aDXdJSfyAJn02VRJL
ak3/noK91xw7/kPHJ7eYDUVeHSinN0ayTMmZPgqPjsB0DLr7HrEZG5VBvgt+PPWQ
HwJ1URh4G0bhsquQw5KXaJI02DcE+kilxWVKPOl5VE3ZqyQgq27KAvrzUunXyZmt
tOcgcBYgHNjuhV2/le534n1+4LU2kG9M4s3nurYjECMPOAhK6l4+hVntwJ4GBklW
HzwfJC1UQse8sCzga5lQ40kGswIojPaB0IW6assEzPbOYRkJsyyAhX6ut86DBSa4
uPh7YkJZ/rYJBJjOIBlSuY9ox7R9mymySpawQ4LKwiG+ICWo3r6DzVrfDBroKZDF
sw3ZJ6veIanLAj+QZbIVRpqy0Nkho6CtD60Vi5iKshKnh3G1Npfzpa3oZ9N7t8xC
eS/ENIJHqmfh5CWrl5+BRZncnTkXkToR2q7c8Wwb9VZrkxvd2RS3CtA7JUfo6EGS
GdAV3KMrcf4wdQLexjeXVPR2DNkKem3XXiSFKCp0M1A8zYs8HGhsuooQtVCGbilF
11skj2ColRCEk+aU0nGHVhBBOszAj4Fkn2zO+eQ1dx9KNHZPVY50o+kDw4kRrLNl
xgDBqkwOt/snKHrejvomfwUw3Ba+YphofdopwUQXceWceRFA/BlsQusTqICA1bH3
jTCGnQ/8oqi8ljZQVBPnvHaBe2TDl2BYtbUSMJKYIx/Rci1Ff+GOkyLbKcTf5XzW
DKKZtew0TR6w3m9ptvRHG+4r/N+pIDLNc9DL9gJNJVll7bqNYKE8+QldcvLRqcvK
gBm2ZvJEDQYdX4Ux7iEJfPwKZ988+4DnhT6I/D/U2HxiClyVYY/lESyqZ2w64wo2
cc/5q6YtiCf2aokjL6nelmmpcXTIHwB2Xuj8o7UjzRSmdyi6Rl6QG+A2f2ZI+m1d
e//t9GlBJacTSQTg3tlH1u/0NA4e3btYZ4tiFnR0p115ggkWP/+Q/joBoJhp140F
lduC0P7TP5N8zIzt5HLWJ2F4VopBeZpFA7C89sPnaeFAkIQuxKdoJ1gTtrFeJQBT
HUeUI3cZivRTKZkulrccI4NjhL/mBPNK4uyMiBvxuoZ2N6JqmG3lETR0evI1knyP
HL4wUOgIDVo7jJUy7ME2o5LDqbu0/rcF8rHUr6oXiF5ZsO1XRDy4NlC7aktFPYSS
GDJVIjMC8n9Qf79vD8x73D71VCEuXKGefJuiubuMvWnTogZFIAjWFiRQkD0cduar
QPrm99qy1iiLkB/XOK/W3dCFFWdIYSCHXeZjMyq2sx5AQaZ7uwv/vbJTnwDSdccH
9mZYUg4llfIK9kJRPwAoNy027L00Zi6owlYMJ9uFqxNrhToP+Myu/CnpdfRdXDzs
XZ/nTbt6Bl9mq4ASOXpta1iAO12KQtaxuLo25r6iNK12DQ4lhNRUkrOb23MzkTkQ
ZqDJra5RQBXVFRtbiE2ntVwgqXWjdziktUHvrJhogvny2OxBLBG8M6nNbOxhf77D
HTkhVap6WLtZKnJmimRvp6yfOF/SEZPxwRRCCiG34QkhQZNfQB2dCasgmdBRTB8l
4iw5Mhp3wzbJ9l/D48LndELH6hqNxPyRncVF9JTQsWGXZ1OqYnsDl+X99Oqfn7aS
+uGBedd0k6RD334w690D8H6i4PHyW2tXkjbJFaG9uzA1eI351TutHlbWVpZ4hmec
B/oVf52UnuXdmteBA7Ryp460h3CczHWwMIit7kz7N6EDAN6dQ9aM24lZ8TKULFPC
yBEXkBY/L/G4Vg7KPH0rxlE9fj3Fa/k0CktKK6TBYF0DKOPE/94BXKB2+pJBJ51g
UF1aklT6SUbU0rnY6ERiPIImicTed+dC13xccBiuaBhkbeNj1t00s46ZLPOQkrRi
Gn/8TIIovIl+SlL2+g5bGR+EHbD/LwwxPiSNhdZtEf3tAjw47mcExFqBmd/5jN8W
DwuhAqoPQoEyVFyKq8JkvqveHzXjPaSwWh3QBDSP41CcLFZtEf12ah6e9YQNL92t
6n6iDEOZBLJv+3HJn7wsMO7cGjsR3wlnGp/R9ABGt0to5u3vQbVFzndXW9qKNZUE
921QIm6ZyZZLTMW1IUFisEEL0QPNjHPmYmpbINXbTOlaSIFIEVmJA/pPq290a5jo
4CZK9RjRTM2C/+oA5ZCTc1iWygRYAO9gvPuauvIoVOB6USIC7CDK83Ietf/aSxjI
RZYi3yib2wYMHOJOhE1GslTdvEazVmfmtPbaxsTPiKbWEdc7RAXz1uTYFpKYooFt
zMa1QP0LqKoRbcqg+5RYhJQdCLirGC0K+VgFOY/HVzHkh1SVQQ9jOifkplerrcFL
6ckxqYV432kCujzmII0ButV9hlR4vbi1ee4wUL5JBAMpMCBMSN2fUqpVR0QX0kcA
CpXtZQMZ76/69UjAqtvxo8tuGmcoWamKoAYsqtpr/msgplDwqUTB2hBaKfr++PzU
3nGd9RzwwcndfyJIK/Pbh1JhqP74EOD2BykE2pjTayeX/INfpvIiP16iJv+B9zq1
e99AoHiAF2R18MCXemf2Cx1LFr7oEUJNAa8Ml//rFmIvAZuSUdDLxrWoOE8Ar1Jd
3WCwHsjukOK5VBcyqldeWB/8RANZp5MYtTYq1+xTHMsQKvlTuKWXjd+DBAxmAxn2
iKUxtv5TwRsTLefhwL2pEXGfZx7Gdayy0ISmlAQf2DpqsnWnA8AH2XoARtimO3c/
cKGDJSoAasb1OhIMnA8NNECUQRt5F5U9gxUoK9w2PbVFZK2xFSTMIkRyVuIInxpf
vizWaJPUEefMLiQsMNFDw6kVbF8xhzWru1FLTS7jTMwVdFtZlw3DfTkuTsizm5cQ
TclYKunXwohAdAA09yQhaEh3YVy2KGI9IETg155ojGFuyRqsD+Ujk42XIa0HHbNi
G1nYH6rGIKDFNXJQp3D/sJofQaUC4Gzet3bFPtB0AIowzH6rrpMjAFMEga/G3NfU
RLxBsS8ppIj1DcXbpfIqZkxsNvQZcrBczU1fibQ3ra8pegNTmV6PsnulkHQN/imR
t2Do5SI6PZkhIUDqgJ8SJJVZ2FcVDYZchDPiUKoYoytd2wD8xcHF0VNS9HuppHQz
i47rYg7TnS4au2jc3eUtwH8NnFFgA7jHNJ9rojyWGkALqG/9dqtL66sIq7e7W+EL
zc8UXNem4t9PacZ+x3WKySzZ9mAFaukIKz+RaXs6MocAbeA7d05YpbW2dKw5FRT/
fPdSXB7GG48EtYNDXng8uxUN/U7mvmN95T6iZc+eNPHMmhrPDynhy3Q/QNIElRbA
hINmTSKwxRFIyOt87b/kJ/pg40uaWeL20+8W2cuQdm3x6tAL6LzOxiZK0NYSX885
+aZF35HaejAwcTshb1ExycOy8AnaXmhw+SXUqRdecwzIdakDy1Mid7tP7r02rCTO
Gw1wsZSmlxqdT0LhByPcoLecs7iP8RSZ9/JYjWFhv7m0wNaawGLj4F3FKMuj5137
D86Ai4JRGGuXdP3B0xWEgajseA2QoyHBv5sOE8mnjKUJaFjeZ5t9iYP5F8Pv92+U
hW2Usz8dpUUO86S+4r1Bjo7yMpIQaaQPW40P3YsCNmkaRokB12HI77u5EKSZHuPW
3JU+c2r3GGVZmCsaUF9tLANwjn4wD3Yza8quMH8S7MS20bEf4JyovIUqJ/3PwPl1
elxsangveBzLeZ25sYupskf9OxU10tlpshX15nBAV6UbvAtZfP4OakEBSC8Zx+/y
M+TBBy8C1HzHjy0b39bsAuRyNhT2rbmrgfWBYZCD6Y6bfgSikXGdADQPRSWtr0/z
o7BiBFaUZFqtXEpanui8v1loj6c09h9v5Yum9rP4pT+piyishd+ds+8zCdmEhcHy
2PUk4hi/Khlt+BGZM32NCz3/JCX48T6VZ02vip74JL/Ipc3Eh87FevM6RMl9IWma
VCSuZQJF2gkyFUnHz7VFnLk51d4SyN+75ZRAvpvcHUoGCqsdHCP0yYiKL8hMPC6K
uAw2jdPhX6OVlghG/zNH4LUvmzIqbyDb+3X9BjsgKEQ8Lk04K6LKS0bHflTWNP0Y
VSK7EdPT6xg5ycAOhZ4Qeup+4EUTrFbbgJfywZ8Ji4Wc8Fm6KyJtQuyOyjk6ywnj
ziEsT3sPS/qK5ZzjkyGq2FppZeVddSg8DJ80d0KzSVuxP8nwRid0/jlTeelVudA+
hlfxjLud/u5gOvP6c0S+S99fHFE3GojuZkiFdRCfX6zYw9fAjnkmXQ4BL3tBfGou
CTwUeFzABYofDeUUqd5/KkHGr6idElCiVqhW667QwgySY3Y6SQgr3bsHkgbgbVKl
7XZHRyMMKVborkGqTLNDnNeN1QIwZksbfp6kCowsrYKtMKKpwZr3tTdl6Iq0zh7F
zSurgLFPa6R6cfotoIW8L2+yPwHZz/6mRhKcK1sX/Hi6YkoJ9cQqCFfHZ1kLuBEF
NoRTosYEtOJwvrxZijm7pemsyf6lhozbxsdJ5ImUyrOaXn7ZrZ2OhKHnec7SLdNn
xYIl6FE5LjfPUOqK2tplIfXQFjQ7gRCgBk4d8j1gfnFFcQVze02zaMZB5SZHQMF6
+5WOKsCMBLrm/b8CuMUxtqO94s2fcHjN3Dtz6hEGR254KLmHEXvlZ1BC8AMSFi9D
/M+loOmYLfDWeungTsTbNNykHIlUW5LaPdtW5LVjoKvS538GXOo0scosNHWkf9zG
WhlolGIblXrceE1bIGIv/9yKFNeZCf3SQP5vGjwE9yMWzdyHPESsv6BPCgAQTKHD
KyEod68eJ3YSgSYSxwIrXqporG42lTEysbqwqcetHx+HADSKcTW9zUW7wcfVhH0+
m12F97G5Hf9gDHWll8P9qXU7bpDArj/+AmnNVH4s2oJT9ZJ08IIXExhRaxgHiqht
UpO4tSzcDXC80BL8Amm/x5xFZ8bGzkruuxyvaubusyJu8EFkahSM0agAew4Z3Ajm
huA2DP3D3+lMiv2zozagaGAg5ikpsBc7CZVxOEym4zCeLJA/0axTnHEbGjRad1D6
PANQQBUBRoK6DJ2k7ysSoGROPuuEQrTnoZJCqlZ2gXSGMyNJ7mtHthNREijeFM96
iR3YUYVyUDtcE7cKkxHtf5l+rA8LR0CfYfTU8Vbu/QgKoDdFbxsa7/+hrwOg9mYx
v2PsfunrQiI82ajbEfhqOE4xDUQbi5/JLwxv+3hGnSgNg+ndHCSBWn5xCtCC1fdS
lkV59oqXv4LwzPTn1ZupcoiI/d+gIRFYb3e+urNPGMOrXRcDpThVQEP/cWqeVTnk
SM/X4mXpfOvD6mwUjaeA/+n1wz+DA2ZBhMFsz+d0kU9knHV//8pwuiTvbwd8u12Q
+gTEMZ4sRFOv7stOnt07Elvt9DaL75miB+fIaKbD9MeJjyvQZDXACSqJvkvA8C7z
dx25pP/ksSzAlbXf+3iGp1KfbA6QYiGrVkObqBe59RGFkps30mclhE1pwFjdrcxv
m/L0x8DMMJsHOdHYcRgYk0VSRhwPGP8SsQmmh2Yy3Ux/9XrbxVm9uctpQfmKEkWQ
hL9MsvyoK1Pp1UAyWcRbe/K4u/w34PK21UqFaavx1ZlFOglRpT3hRMGeySg9ekEy
3ORiSvBwIiCxb9ul0WdcOao0WgG8Urq5o8SX7R7+mRqfVxenItx8a8SHsAeB05Kd
T+Gf1Rl1biHyA4yptnJzeNCkJQKhTTyKQjORFD4E1yatEPcz4sPtpT0SyCowzgTL
2yWg6+KSwgKv7O6kRRZVVVzKmzelJexypbCaJ/7+EYozqmDsD1fsdY8T7BUbWR+F
25BLj4ykxa0AinTcxbReTE68mL5V/NlKJ8IUcfHw6eNIH0V4sprAqYT+t7lK1CdK
qc2H/sk0gRULkFr84Shcqf4dCdmMEX5IJvnbtjUqprtNKLPiIrdn0apyBXLBymXu
2I8g3wkmgBzXqGPP88jyNGj11GOtP9gdSW/sVDDT//IX8MIaBkTZWOVxfz84uWkI
NWlVu7TgDbUXUZCvxl0XJR81Z5XzLSFFWc+YYHxSb7Og+iODOoDP6v7iftvel+47
CPusmKsNhbSurUpOblD6Qg2g+tQ+dChEluSzBnK3kaf3HqDSoKuXtYIlWKi3V66C
jBQCkRAku0KWQHvpyCe9fH/ZDyQVdcmC0uW6+weljgZFB4p/fcTViPjhMn0OkK3e
PoEXYALGuo3lHFRRa64MRJYnRSUnLiALWz9DtlBA1Fr5hdiU7yDm2MZyg2oREmCF
GMrnMHhLMujM23GxuunUvkoiO5wZkbhOyLR6UKu+Pq1NTCFSD93rIPYq7OcWzq/9
s/b8u4JLWcnCKOaZtIxciBH0taScGq7ly/+lYejGb2F7jAOS9q1he8yY+YNmXbgp
ZiDC92b8FDXYbTST8/yJ5WAv7G3ZYoHNThlTKmFE06OkDWv9hRksVyivJnALmklJ
831LlQwmOYCV9jSYHWxtSlPP7dCeh+9fHqHUz3AdFOJb506BP3McjYreiaXMiZhA
VFVaATrJYShsIPB2uL9ZBiBXdAFTZbEnN8IazPCPxUUqiSW/XhewquireycpGDCT
Y02AQVIvi/LDAG45i4CskQdOE0+j1DUhqZXJNcwwgF1Aw7dxSpbD/Cdx5FAJCHpH
XAmxuJKMiWn1PAOmP6b8lvyEnjM80H9EXzzJNw4adDFefuVU9zXXZfGh7X8DvHfc
0yKg/7r3PlTN+hpwEwbFuRH8uA3ITd+hS9Tw7NQ4AJLRI6huPODxMzIY0YB5lsRJ
0OIdx7JJbBO4RIp251FM9RjWNIRPGZLw9Z/vtdS/57KSuDWzJp6sAST8LNVyT7Ir
W/LyY9zMc00D/oC6m5lr3utDXuUG2FL8bj/K9HZ3nu3btNd1QkZ3YHP16WVXp3Q9
hQc+Q8k/+P2ZgmLL5hyUA2hEgYaqADgvmfUCjjR/JxKwV9yUMHakJGEohoAll72S
HShysatE0RcjiQposC37Mcivhh3ncKeZSpMt1UN+GErcs8KO1w74WqMMamyM6zbc
WsBu2lbx09HpSDE3PaEknE2BqHOzXzG/gW6EKInOE9Ka6rf6HpufcV3R9H8DR0Vs
CEXffK+JY1qQQfQOxpvX1uQiVCgSw87pLYBjZh8KWy/2RM973mdbre2hUuJUJdSb
8+5SqE8Dfh2MrrqQc4Axtj/oKkIhuGXpx5eYz6R8PEhN429c5ezNlag30CSeSmaY
t2GVCPGbKAar0fx++IF9Gsn7sO4NbrQWLbox6Uc2WIQKxRdmO4KLy+kw+labe4Vq
AcBp5eZDs4rru9SRLqm8RRsA9JgTFCDQSZ0OdLF0pXlwF/n4/izSBIQ9lk3eira/
7hejnq2Xz1uUCXb2wN5tJf9ZIQK0Jrt5akh7VHrPcCJSWwKYCCpHB9TAqErjcRy+
URxM/Ab/b9ypBIzZ9xXxaNBgzI77MFg4MwThcdOniOkxbG7h5jm5rIFSKZ/ZAC5X
+XMFIpkIhB/MzBZGxplj6SvXn9xz/Pa2YnVMGyl+0NtKk19f/Aw3FP+zhPZ1LkPZ
oJrrY26Snzsv6kGpRs6KoVvYCGbCqe3XMTUKguO46OyxK87+EfCTw5olYVvEWJcm
LVUXB5dFhtG7tb1fAeClSoit2Lo0HxdBxztLF0Knn21WgyGR2WaU78mozJNB7DbR
mGFYoPTP3SmtFy7h4Werj9QP1R5GQye18kqdN+YCrZ2qQP08nvweQOBpd2Y2Joh7
W/h55pRqM0l/xBXquRc5mU/QLR4wzN0xGCwGAZDvG7YmTFg7wxY7CspTHPnMeABD
MkXgvOlapxLPYAECA/tXPM/rRz0qU9lI8CvBRijTEDqefBOKBhMH6twhU38XnBz7
sKIKEH8pO9ESiFm+tt3mXzUxab2zHilXyFq9VlcaHBeNgMXZNN08/TEmwKj2sT9S
ZcPy2fWXVcazuKtraQ5TtsewWaDC1GiSPZQWOxn9YaJI4sQfyYLGKj37DECBBrA9
s+CvLQcpQo5rApYsMgZEFl9ikTJZ9ukXLlsib9UDvMcj5uYCcsqCe1Crry2n4a09
C4bxzW7eLuqkpzuHXHlMjWFXk8BnUbrUleGaCCLymUNmTW7J99oVZEfRWkNgxRuF
mdrRHYS1y7BlaTViuaDzp1hj3lWgdEupsjOk6Kaao/ux2FMm4gHJ3C7Td0lTjFnf
0fDvg3qJRwLNGshQWSLRrhL4A+W5sR3OoQunCiGtRe42CLozL0kBnJkicSAO+Z4g
X7+eVqzw/eh8UKKyaL6HsddSPB5RymsHAtWrB7A9IW9E9cp3BFOQTYu9QNPy/seJ
QNY9lmCxkYDdyTX/BMrpeD+DwBMcWaIsmD2uXdvCkAbGXtJqIGICKotzX3pLQagK
38s5Rk47xbupR7+IBaLLHbyvWC/C+N+q8wb8BZHvUVZzH3LAfgpTrryRSmyRB3+r
ZIhxBxRqulsnAUB/coyMxk+2rXjQ4tgpv/530mqv1JBYZxIirE3FFFQ5AyJHSLQ8
sA0MaQPI9prSOKYqsPe25ly+5kz1dgphuGvGe0OFivdBYK3rjkw4kQbLYpAto1Vj
ddiECzxcUgM94G1g7Dw+ZoXi2cR26ujCExY+B4sKAA0ILznztp6U1a4wzUHiqj+p
hQ4TH+TUlPNP5v9EwmrrErUn5Ldn1tGlRG0uV7iN5Xt4rX3pwPg16CBHskjKeA+m
n0ygv40nCyar4ntPX1YuRRGEeoF2/0qjTdSd8jMeNJQNMieHOzA6kPCN/SQmb8Gm
HSzkNwOucq7HF5yvaGRkL/OJFWhA4305GaJWGBXHx9UhK419e2f30mda+Y8HzrWj
dH0jB8tcy3wlR7tYf8PVZqJsVm8Sa8/T668Xgj6l/mbxayXYiuNocx204lnSxA1J
UXak/nJwxumzm9qEl6sKqZQBmV2MXN+Uiljzkz6gZxkJUiGIHaEtwstou5ZPvFsT
vcxFK9IPqYo1wRoe69KeW+PYTGarZViYE7qJz1yiSDyVw1WhaSIzm22/aOuKBjFw
S3xFMqkVtEhFNSMIdcN8KumFyM6om4tTByON/dJVvqlsTGLZ0Ch9gX2RdOEZ7kBD
OZrFMcsB4f4LUBRQTp6N6e7HxXZWc1e2VI5BJKN2c5si3qvUhs0UXj9VeNgihSC5
t/VMknkt3fINWeoseptMP5bAvMH/XUHJhOk+zc4ZcS1rNkKF3rCCIIYk4KfJSvV0
6MjtopA2ho0GJolKE6bHueAJKppzyujuY89CbVAGOxa/vLYuoqufay3Hv9JcslSA
CZHsrgrEmiajS6pwSDGaNxJflUwxl1VRNoaySxjBGlUnF49NIpzi+PZBqxge5XaL
Na5CusPu/5LJZfvPR5tiv1wybfiWJrdjz4yG5W+FvAepH667Z9nXoqnVBDHZvx4G
qngvdCCiYVsHkPJPTqLHYI5Q5nZa7p4p4QRZjx6g9pzqrH+nDcqopI7hcIW94kCy
eGHxFGNFCU+75cnN4ord3WwvDHZhpI3CGEffXVJYVgwz9oejR/YVO/VtM3Ia+SZx
K0EQSwpY3PGiRsaPPQyvuhWIHejxBYhjhv0e7RcadXlGDCsTbV0W3jj6X3Y7ULLg
+MEbuOo4JnoCVMPA5eAi059oYgZHB9x+ndnVoa4th+R1AeNKFxiVVLikkWTUajun
5r5k8/HN+8okkDgR5D/gNC1h3RJHdAITCxJQlYBZ84skmd14dbPF+95Xm9ivNgVY
ZpXp/hMNQcLOYvuw7sQ8ltRYxAWfiA/dEn/w3MvyQmY4yG3vPCEn2sjShpDiN+/p
HcIv9gu+7wT//n7muoInS0MedcKyOwPvSal4HfbGJitq6Ni+HlmiDWHuqW7q2ZKT
mQyc4xsq4X66r88tUhLJpvyFxmWmBsnWkQ4vJzWvfeQ1rYTBWUg/tQLk4d6mt3c1
IJkmvFqYr+Q9RHKwr1C6aUjQL+nJ7C0G+qWwyHBQYpPmw3GEvMumy04bB0SwKUrS
SmDLYhJFaQ1U8fiJfnqQ15XRXqYF+fhe9D7dV6NuO4shkFdSMLA24toyCem4EdNB
FjWLbTBrQP4tUeww/rV4DpMUa+Ma492cDFc7l3cLqpGCkHzPdzksa0MMmxanEE92
j6N9BWqk8JwjCekAwI3xtY9fdFDcL/jSt/EuBc5wPPzKfdNmWswLW0nEorFpElXy
VCIqCN5135k2VwPIB7IrtD+LCBB3G32uPYfBjI+KapWU+sVxMb2kiNHw1oOYOk6E
6qGIFVBsKuUeYtNxvDRaVM89vdQdNuT35FztTGTBYUGHhndle+xyTa2khXPRLCKp
v6AwNKPYvnJ/fXPFt9w3I5YEWUDMu1DvSkRs1D0ngG22KEmyEEosq4V2PJiO+nkf
qTAewXnh/mgsYpP7DTb1CpReXKVMalaqR4XHbrhOcLd+fYZvvUM47RUbM2AfepLr
yngt6/TB1M0GqnIX5Pb7y9OVHItKLb9u3RS1vLfWVBnMBGbDf36FBoJ5Mo+wWQCd
R+tjAQQEBGYn1919fBUIYEht2jYZ2b5tkg1Q0w/J3sSgdLC3WCJW1bzX9G+i3j1K
zg8G1NajSKyKusHz0NNGS2qWJaELgr2hzM5fQn07CFhVGyNRVmEm7mze6SbLvEM4
21VSzTuyJvD8hiHMjMCYV9PJUASSR3Oq32yndqQLTi4zZfyxVZNxSB+ytjtC/Xn7
twsURWl0CfFm0sDTCLjfCvlaqbIUaWqLBayVeIv1xLPYT9XukfvVZPZ0NvZ9qjAz
rDcTwrVxe14BbTeXeJziA0pvcYSG5mEkeSdzSto6KTzvTBsxje3J+Ivh714bdFmh
bphTy2nbwRPalEpPwoUlUNfwE8FPM50lWU5+dTY7Ysw49NzgT/KHhaqm+9Ju+VO3
nmeMK+SQX6Bfiw6XS849c2Lo5g3r1HPxTDcnbixl2UPVBye5oEhayefpA9x3BzbU
VmheirzumIY5HSKV+eIX88baE3mAJQAJ7dz6GVCBpQkfJDoth0c1irg/Sp4tgfVR
0K/cXln84skcqn69Slaks3kJYDroED4XoesM5dEX5R7u7PDO6h4hViM+t02YeXUQ
X3Mqy+KA7PTxgnMaztniydf3V4aNx9x9LuQsFmrwD4hMKUy1hiFB+EsU32gGo7Rz
rpwT798du20i8Hrpd1nMu9c/Dr5nDiL3afbPass0WaFyJ2HNCDBHzm0Qg7/ggmw2
2apFDuKXxk8mSl6QBkTCbfqJIh2GFYyeyVG1PWmWaRij5zB61vsRnZSzWqH+IBVz
Q/BvqbXcSNCgXrGuOxV5v5dnsz6lzCQGNvc5D2TNmyJIPUYdWz/ICsZO4S7Ropw7
zjsdIt1SU5AqL4gBUo7X5Jx0EYlc6BvEknb4yXpwA4WQlbxmzGwljN2si67nWEFF
/6REBWcfp3OY6/ZOt/c568q/5Uvwg+kBrbJVjP6zmOHI3fCDXVq0RRCuvISXYG0J
uBseHXfcJlT4tpTcEFR/xjXrfvJVPzkOnQiZO7bzcAhUSN9MuGpsENbncA482ivI
otHqf5SfigqFSysJ2IhiF24Ezs+kRNqrWKHgMAp9Qj9N3lhAZzjXfRNOe/wgSmdL
VGuNWKKa2IoS5FO0O3C0mRVdN0rbc+77UD/SQrjJqEVHFuzjKxwtZVsWKVDm+hc8
STuRrsd1X0yca9geeSPRmo3INswUhgvM111CGFpetX3dPJ1XbRUwwr5qiePbWonG
YuKlTmck9jzgAvIpD7NMPGR5uWVPxCJoKPiIMV/xpBm38GoO6lOXiG6+aUBpnx17
vwAbt2wkEO5fQRPEu8XYGRVY09Y04TAgvlkBMloTr+d8KDK0HyTsa6ivDHD9taKw
psr/m+FE/L7OnFl0NEn01WFYVV+eSnEMCjec8DBaHLxyWCFgPDxw9vCAxeOak9uK
ln1dLkKM05nWUTmooLqj0nfKX+X0b/DRkd0GZ1+vq7oBRVSzc5ji+fMIOSZfRZrU
9qZNxmYD7VmZkNHTLS5aIWJmSLcZwmPkdNNg3XlQrVlz3JmAfYS6UKB8HxzAUX62
nvXQFzsbu4+e4vV2mXvD6NHIJCmDAKrcVHavSlrttO/CgNAHddwdYd4qE316dySV
zGbZotdMVHoAPAntHq+3d3DkU1KTXQ36WIYbJn5kLfvw3TNUT0dcFKXF3iXq0pt7
n2YjloYRcvg9QHnezPIl+kWRcyHw3HzTXEXpx5Qr3sHGahOtt6yhiwkB6XXv7ulv
DTooFAX4CGMZZJelxsGOleprTBVTdq2ZgwuNs1xVixDtPYSKSGPq3D6rCBCz+44Y
ayQSQ+pSOiUtoTimqQqC2K8vErx4DD9s2SJJcLWwHp5gunVsg9BZC99FpcjUPfiD
0OityyclWfBXr1beaYm6nFkGkWEKvmLItccT5uVZUdvPJmD+D9skx2uH1k7HjR6P
JYi8h7weiK7rzGssP2PzebG3PhfdFo4mMlbiCvmTTQ5nIJ8VGMxQB92GYwrWX87K
bsccw7Yfk+ifKNeTqUNNlFZaRzIgch8pMnPF1+X9JDhr7+bGjJzIwRVu2iGV+3aH
Emhi1a2BfflV8P7B+9gIKt72KjCO2ZY+azSIO5J04gn8HIWD2vSIfbGFCPQbSmLF
CzQ9cn/2Iy2TaPNnqELLHPoT6gOYQcsmYHNOBtGjnCGVXH7g/wewa0ueA5EMHHn1
edfROJuOYboWDeQ0kJxRbB63uDSgJQP4/BWeNN4oyO1kq/miKKOBYX/Zaa4aTQHE
LTLeVheYejPjZBvIbpvjoqjsirzHkW05N2Ph48bu8tN9ocRX5rdd9RppID+kUV79
GdWgnE5yd6GwK/GL9G2SV2mXx6oCi4UP8WzZfA7EtmMg/rcluK0KVs9HBRkBCqF2
UwLag0WsEFxOWDfuPXSLmrbcT5UmlhbGrZw9kEmqNBY49y456+21aW+LcGbpfVqh
9LhWQkDeEEcQan4VT72LEsC9luhanm6sfO7mgqvTqCMdYEzPYDoOBnRt6atRjSA0
Sh7PYcZ45AKlDv19VXblafrC7PjAt1hp80aRHmLd8KAap1fzyu08x08XkWfDAGCt
tuRi7UxCUTKzPlXIawCjB9PLB9IbJCGeKcEl1vDsmlldVPg2UxM1pMguUgzT7KEH
og8fVrYTG0ySb4T1Qm7QIc3irfkUanNnpXLs14rXPTRuPaapoKuh7CxG7DLn1GpT
qGKvkTqDOiL0SxKnXYJaGIRvUTvvNurjf1/5MKOPb64exNSP/rMAZJaUCUBeIwOj
AqJuyRN/Dcu6EU7c97UcKMiM6kAjYawPMkgHaxuynGyUhe9BNjMFpGYN8TJeOKR0
2CQHUR/XVB7nSvd0G4LcFoJTBNSTfsqgSUXNUqOygjWISCzXP2HhF5wNGvPuq01B
nMP3l1NqH1j/O/msGldrZPNnekHx4YGe0TIkCwpU4EjJSRMcgNRxHpVVFU2s9Y1i
CvmumMcU9AuxUdyArq1oW/sE/xAHT1Elxmt9L4naK1MzWgEsaZzdmZmIe4qh+tat
oQbfs+cKHjvC78opYjtuAC/ij81WKp4fmw8OMBNGnczfzmzpVjZraOeE+TiyYzMy
OtrdfNOgztGx+cKnNA7KO94pR8H6m/EoEidvgWLHobKlJz3RWjXdI8cG1ejrtjFL
475K1DSH/KN34EOWxUPIQfmSO2mgdn+Q6IWUZre00MjHS6I6F7Ra0OiKH/1toxe1
yi6VfkH+VQ8X/Lmu+CSfzBjZHsuRFHwkWJ65Z2qe338WgRC9lelv+8scAUdjZ0pm
xoxAhGh0kPOzzbJBSMQ+mwzjYIo7p7l5vXBnGmJLOfyZiiXq3QM9BNbcMn/7ghcn
WZWKKUF040F9elcO9agYiw==
`protect END_PROTECTED
