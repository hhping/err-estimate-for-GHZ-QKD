`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ercXKNk9yUD7jpvmZByULlElUwFz2LfRaqPSCt/0kXTezqF/7lp8Q/fw2Mh7WeIG
egfnZr55ua6vdl70vXJ5yUSXbd+ts2Mc9zl9EL29vNQsCn3p7PFhiMYfi+B1yE3N
spB8KsRiSL0QrU2P/bGMasxI0BkndDbkyo4CRye1ND0WLkpqAdx4rp68Rtsqk9Bi
iGXuB5rbcS/vIbb9FU+7pPEd9idu6TmCrOhiPNMiILYcDYaOHr29FJ3mNMCjFiqM
eX7riHgiScImhujxDxgQ8D+C4dQzTq8mG6jvYL1tbZhylUaeIsszuPvKplk77rH3
wh0tN6nU1P5bFiuLcY/GVKMNwW2yWS5flgqiiz43JZSpiD0DW7o7JFhNlat3u3YU
b5FMycMsozBJ2+0qjr0ZPbV0RdCA+zDG52HK23CcC6uBYFe3KO2F8fm67L8X4p0I
AHexp0jqhgip+Do0J4cTlm8/zoxmocJ70vupq1MykkEHVYv0xTpJpi7fz+ikdVzZ
1X3hzyYkG5OCnPou6dkSywdUDQBMtMY2Kh3fKS/VgvLIm9ZTGEPd70PUMCZis/WX
Qh9x4yQ+n7RomAb0k5PXVA==
`protect END_PROTECTED
