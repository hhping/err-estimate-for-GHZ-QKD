`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhcZX52gq0aylBNhmzhPIZ0xI49Pl65u9z+dPJFrJiyYHliO5fsY/8q2bkua/4o9
nlsUL1JviLBbn5Ylf9JYSgFUhERm6dPVFAY4tUUdt48sswIpuR8P1mueXe3vyeKH
KQdXgWfPuBTuiWSlIyXRC0wsPxedqX8FfYv+D3X7P+RoyozRyr/s3hvOpfKEnpoP
XebhOWMlnSc3sWY42y7nggwbtmhNb2AvBwJKxDUnQ7m/gnBkPkuPghMamWJidPnb
KExSC3r/hBOEVofHA4nqg+eWSAUKrqekwalhj5wwhNCuu1jYFe1Hne8T/6GOBV5Q
oiJ99x+fDEOVsMn57Xnf/f5PiaqdBI9/qcL7ySc9rHOqyT4mOOMkkSLK3y6NV6qo
ArmDGUabQKlg176NsEgiFbrlHrYx7UYmSPmnJwd1RM1Wau7GPtxAtgXwjaSW64Aj
5mN2NkEo9q+isrwVUszRflAvyNqzn+SVbKkzmzpYn5e5SqnotjsKUFfQxXs3HQ6I
seDQtT1O5xdtRuE4YUKzDB40Vt4NhJ4xKW9MWiqaiy2aZJDA6tdhoukNET+FGpmL
q3JRtSArqNW6X+R/DSZbZU1UewdwC4MFNg+UHoEGMpe2nayOyhpzC9KJWlBzj9Fr
QMvONz35/1epvj9chhgj0MVS8Y+Z8zFvZtRMi3iYni+sKsuieTNzmxhrka1rmlUS
NYEv3FNwmAhkzpYqeCJd0yR6K7I3oSALJaEETdaLJfI4ctWe6Btb1ZI0qlHX3gxB
/fiDv6CyKKLjKtZ/43qYAvOLTSGGdyavviYAIMhImwiUAWNeUD5xm3NsAJVxLt+r
IUgBDC0TBt9rbYxddtT4ZWZF1J2N+b90xLTPKJVt2KMs6dL5uVrHdxfc7/IZeVbO
02kJJIfjrZ7Lhc50Mcx/rfgOYLO/ZNVJimL6uGTVa5VWbr1yUJuSdsDs4Folcvde
QryB5LEck79GUUGQQMZMeT2ua7ObJi3qwaKm4I/1rwuOdzPyUn+bSOjncAoASAfF
TWCISQDj9QnHFvUjeYSesl1e7fzBp0rqJIdo6mQXI8GKqjohHv3ZG6E+XAblXtto
wfwlTXa9nOUvqm63UIT44UXW5ZtwLB0GBV6tArI8wTWMACuUkITBMy8iTCsQ9P4d
jD/mqHzIKRYWU5aXeMQz8skPq1sXQ74o5ePsARlTHz9wxtdP5yyYgd29OR8de8s/
yYGmRkdLSyAt6TP/1DOtSQ==
`protect END_PROTECTED
