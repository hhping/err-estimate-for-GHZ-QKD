`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2N9WUzMIQe9/pz+iZ7HAtoEnzmSuKWfH6hSixiCaaSUbqgLEstB/FYV0LE8rFyp
+TbQ+WpgKByKtLwu8BdAl4ggwulBBgQC91UkcF3/WYHV9WuXifUGknHm/343C/mG
Bp0ja7GUA6CYj8NCNjSSeF1FPSMHIWA3aql69uJmbIVAT1Dn1fpBtzDw1njO0qKJ
qucoAqQG/8+ETtV8z56uGNfqD0aLIrL0b9bneXjoXWSffWN3k88hcsBJ1gwq/JW4
kBtbHoHa7h9gcdnfSYimuDHJqyY7cggkJDGllEZ2RojvO9OrAh8bed8BKk6/E4jv
V635N8RppBim7o4qlR94psL8Qv3jF/t2q/kQuNUtX1IuonxNSXzf0v3IXXEfVtcp
OzDHWInpeVEhbUbG2QWHDVC7XqJFxxW/4r0LYIkQzVUlU1Tu5s41wdtazX+QRyhA
U9Vktyp8tj04HEJgtjqqA9T29//2xG/RLQR5ptNzxcfNwXb8MlM+VGpOmXb8+Fte
LP8R/ws7KxIVOoSHNNgO0/mEywqhE8sdLVz2ZHn7ficqYw9wtUBiuo2z06MKXlnN
Z+3NZDlrrA+FGfVxhZtv+0zWlnt7GExqTHnn7qesnMaLdmIPGJcs+foAUmd+F8lF
UAeIZJQO7yyW/cV/AAhe17cHBJ8nOCiQQLwToK3wkak=
`protect END_PROTECTED
