`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhLWSmFAFYtf8Nt9VS4OlqsaSNq4w4iBju9MYaWwLioVv2T6C2GCaafC1COxYwH5
dsWbN0uHarMdkWkg7UBcxXw+brEnKtV/n/upy3Z4I5xiZfl1yvrci7aYO5+mfZUX
oKzIjqCINA29NJnskmqKeYkZUIelklAXVM5hbIV4H4tmsp1XUTUIp1pAYHzbpK0E
9SyRZLRnhK6A8Wh9efOwa5g+oNV1UJjNlQy+b+GP9XCzvq1ci95lxh8cvriEOgul
1WRo6HeL2LWiTqahekG5DJCdrCFzwfLyPQHcCp0Kb2pi4kaNUE0MuNcH0dcNpduT
YxDWrFApIa5Aq+bekjTzbcLQpp3YhEoL407PpYvt1jwiPeR/sOrNWPS4PpfMeYX0
Plkxe9pwU7NSZJ+LaWB2fTXhtMJJxm93GTr3gRMSZsOi89Xk+NBY1wS3EWut7Yap
2nEEPzfWdxAvvs6XbkRb5YWiBDO1EYUINdovYh7HjQjOvr9Ox6Q6oI7xQQ1CM1AZ
`protect END_PROTECTED
