`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2e22SkSn2o3Ki7muSeP9i7eigA8zSvhPzqs0kXXPSn5GcJ+DfvRGECEPrqDxsWK/
2+dCRkl8rOU02iafxe6BTIaU0n2pB70fjcYg1dQflRDRXsw2Maw95oWP7ukfBvhU
SG5ZKxHgQ5UsNMNAVqBRABV/X57J6R4zm6g3Im1/HS9hbQLwFNiIt1kccrS8yifl
/bYMJSgx8apCDkEEVn6AfFOYW6L52ASyoxBwALXLlCEIB2wMqey8cqUck7kIat5V
RqEnpxe/7VITEFJG3rw3FWo7rsEoPOpcDRTXa4pSlF3BveSxVtmWSXgmz0ZAjlw+
rHO4t8qppWgfnzEEKIhn28y2yWMF4x3bADLgJIbSTHL6t6Idq7eCUIgZxjjgRQJU
GuQqXEbsm9Fu4XTB9MhwMcpx5m+mwaccUCZNmDxao2L/X5sqeFbcIsCwNQKr3Vc2
IekepYoo0lcVGGjqhihLFg2uQwaIc+/YSmn74MFf55NQhiIyuLFRb/BplLq+oCAR
/ODJygzwEYOTauDKuyjLqG8tDk39HrKabDJpC1KOzsT/0sFLEO95YTuOtY/thJnd
kDPfHO+v3ckNpZjeXkCRG82twJltg9pMEJXIKPTzWVjWzSC+t8YAN8UcYX2xR2Gj
TGxz/kwPKWdzOjlgHUHBteqyUFvOqbiRXwoTpAG8PJuylFVdnWSyRfzRteKwksFm
sXpusYDCTeV86+JtDTza2J41IvTjEW9yu9/p8sA2mhS+XXAU791g4pWTi1VLY8cO
AbTbD0Sn7NA4H/lUjqcgNIpuAcYSyQbodHO3h8TD033uTGa9eEBex8+FHd2Xtp+e
vt8goZ4+ugAWxgSb4w90SVLb3JO1tEaM6B1Ci0uKYmCueZXE5j7/lrBSEumq0e5y
Dn9+bfWxN0jqrviCbX0YG/OZGWJ6rpCORVFRss3YHkHhSp+dQ/5lMY6z4c+DwHuz
+VzONH+WIm9X01xchd0NNxRx3gGqGWBS7az9Mjn/OKy3f+7zvDHez+T5VHIDnWF4
DeLJTjs8CQgVynyatiBU6UPTQTa/S2Jet6J2MRSunpRjWd8s8kFs8gX90/08LPXC
RPn4xv4izTclPaQUliDmKJYGsPkmTu6mG39tqTadF8LgZemSOgsLo//eKxb5V0Gv
dvv94yFSo4Gs5Fy42Yi6t7YaZ5DiNuThN7WTZ5fnlyYhK0sr59CDezhvsM9mShtB
85U/gq21DQSfaiK50o91gdPIZu5pdIchIQxkLuP7kgor7CJzI1zIa87Fkz76qrJ4
PD3bmMXbFQ0NLDLSvDaY9WpGldrJ/eAIB6o37Yiit/sAHFGad2316BUtywJWCrDt
lzX4BWEpj7SMHJlIyRNkS5YC1qF3KkO63WVXxxNHtFoL4T7HMmsw6VMxmW/9tMgA
qOL1Ue2Lj+jQidVcWzGiF8WmaCb0KPbdpWGQXXEyaLqrz7SsXTaOYUo/h9Bh3tNk
JbO2CqoaM9/qlJpWMXBrG178NvrH+koO5D1Pop3r5G/toX3MHwwHEwgIHsai8LhP
5zCtEFpYbT+ok6iIfLzqf7nuHdUenpqfdvSk0akOo9LfjAewLCO3skzi0/ctCr/3
jhqgW0humewfmgDkPP1+s4/rAl4MqlGqhqEljDwbByTHLyEHwW+ql1h3yAFXAjWk
fjiOj+nRCatPFbkTV2a0N0hZbg6PGxuqHP+OwGxigcEd6qR8CmAjGENf2MOV6ZUa
bdKsuY0T3NCKew02JbDmDwZqY6RMsWWMfd43XTx2JAqvsYhD9AdkuWaUToaEHgZA
/PPNIoRTQEVn5UfGTyEXmg==
`protect END_PROTECTED
