`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1xy/713G2jOpLrtRRIDhziBkBkkMHEeKkYm44BNYBHWMPVzdvDGqcD5lxiPkaFj
TPguCT7zMlLMZk/fr6Gy/dxt+GpzGCwNtm75q4d9lOox/b8BgnNx4wjy297GIjRK
2g1swUIcA4aEBgWRa12GQN5DjtmKenMmTpbhk+mEDTy8+9Vyxmr8bTiY7RqYjt77
SVxnSjBbLwpShU5wPIIvGPngnr9xrUwY48MkLdGty/9MsYrGwY8/82nvcsvDjof1
Mq02Rd1tNRSOsPcf7xEtx7Bwga/SHBEU+AZGVaviqD742a5dS+WnLGvWkzo2jW+o
yJbRt5xnS8ZmvVcJg8NXZKRjkmkARiSIrPp+YbKYMgHWTHDzRfBi9ENtFL/Bsqkd
k6UiVedZ1lvt3Cm3nS6VpkGxDK8pkIll8I4XGNzflaj+Ztjv8nBRNzKBPLJ7XRPX
ddkEpEpm10wV7xHcbVI8ab3BKWUIFjEydSIP0QXQyZnsLMI/yv771J3hE3TW5m86
3SgioGIe7J8xe7EussQK8xmImuaFb61g+H3TF6JEkhhYuLaVVdx5v2/sjNJUNVjL
CE4hvyPoS9NRkFTVdSvvI5GKRpKGVuz0efoQoF/gTjkOKTv0N8qj28+18JYgunzR
uJECv5BGAD/7r+arl6JUyYF5cZGZKEikj6drfJS9r1eqvVPDgLxXVNejFN3hBGSn
aPVX4pIkTpu1K1dyiP69XdmduyXXHcAhqACBJMDOPdzspr2F2TinSw3zGNGJoSCx
f73zZjP4J5YEyOD5DXkiWIgQkexL08RNT+ZKq8sbTP11eWIZQwJD+fLoPRt0EqbX
knEqK6wi0JAV/9JUWBS+/AJF/qg84Q6ZiNm1VGQsQ13ZnENZynsMUXU7QtAMAhFO
xuIKDmMMXjjxiACx+Uz2fzObnUuTX2b7eI1yjvbCzNpnyEXyen89o0JU6PkVmapX
c/ChGyraS3LhYstPTE2dqS+RxncuP6Q8oa2m7IpkC57Ritjjo660piTkk4vAsjTs
bjDPgry1PWfl+R0/vgNGhfUvd66hMx35ii7AlWKeUbb8Ji+7WIXJLgKwAXYqJV4K
XEIHNK/uk1bFRHZN0zgSrmwBfqODXGgnRFWy9w8cEVM2C7LgI0shNDVZfrGJDv3S
uDEejt/ciT08+U8ctDqizI7btqJAh6NrDQUy4glCE80OUq+ivqOrBaAat5Khp76n
D9EPjdM8C9Qj1PsLKGD1/0ff9OAgyHdkxUzT3Ik6P3uFtB324uwTnPeldHziOpO7
3rTVtuviIO8ZvNI1gGQrOvJ+OEJ0Mm14pxZTLD4DGvjXOQpCnvsCUqCKQfUAfUKt
gq4loBIAMH8nfA+eoq5ZOTmqW4kP94JxQ630QEUm37RiLl6RIHQ6xXsVbw+BMKu9
nNHKcvvTcsZuZL+QNRs60gipAbSJ9G59VOYRbUy9ZL9fdXmfkjhsEJVLW32E3pqH
DxGlbX3sDPsoEVz5PsrLiSQF2Elz50ckTDuSDk+iufrBrX31//mRp2XGmw/R8NCQ
Xl563pgMZ0f+knxYd9HfzVq1yUGQWKlfDbmaiLl0mASYz2QnmdfggJO1h9wIDulc
ufkJ/JMWIATc0xM4MmO+v8OW9kdOR21A4E97Si5iHBLutc1hm8bqCo2AdJqD9dME
RWWKFT/16421WA0oWGxj7kGpfEY+0MJ+WmKzGPssGrdQc3pO+brJCOEd05aW/cTg
YaETalDUkvxKf0AKf8eTwvZwqZN7ybGCRuclPXdvkXbauh0r5a4uMi9GZ984g899
UK2mD/eE2d/fp5rQaSzUHHUa+vAeTCic8/UAFYbo+dGYZtQr2MfW95mPL60lezxB
8ZFY2oVxHuwWYDdLAeLUcyf9TrjsFnLzhNK9AX9kqx89CsYpZwr5hUNtGiZMTXdo
MkPfd9xoCf0unNPJ9KIT4S4GWpI2gPcFP56m0RjDTCK4u2hGEGFmcTpmjlk54c8o
ojK2pe7oic+DFn8yNuZEumi2+EpWNsz902b7g9T8xO18NAlhFAtLg4XeUvVjIz3K
vW/CmK9My4pCOLsMbTNIpVIawYiRmw+utmWMxX7i3ky6Px5xQvFk2eUw+zh3Oe9d
Ed8H9WyxnMMGXy5JZyMOeHhq6FHqalZDB6sn5YP8+ULeroK3xcDM6X7ad23GBtxd
kLrTk0nPsWEGpFLeBJev0Gk7YcpzLC6R4uHuNZWCFXE95btq3veFWm6GlhOfBbce
jLfcyAEVSKRPhJ9nOqqSzQy1X19Q1nivZkmtE6qGpdm63/NUEYlci5tzRncBoBZ/
lpI8oPsuW1YChO1oB+mJjA0FinCovxWRi7Djt2JHHJPBjmPg4MOPAXeMJ0qZUCKd
wOYA7bEgeZbVVfAFBp2EaJBBP38JqLr5ImNsYzKxeac9e0oeQudWAYfy3xt57lMN
IGYLNzRom7utOedfU37BWvtHHoWf6iyBdMn3GWNcfl8DTqCtx8JrXukwWeJuO744
VTaYIphOk075ssO5xLCQXThfaIf32RmRKL/SyWHO3+4qRQo+NyYiR1+2kHaFiK83
zi6wC4ma2SFGBr7r0gjwUlrGgXJ/6H46RXBAkw+cz4keJAUmrnusQKUYnm1f4Hkw
Sm+g3vB04jXN12LrDkyJfLUKIFQLPrHcIarKV3Y2Obnfgar7DrZreIDKUDdoQ1Dr
kPl+OkM+liv5jkTnYTPyijzzcySA9iAFTngto8RAomR4C9bCj+8q27LQ1NutYXOW
RBWQO9nOWZIvgudmJOwSYWW2BwXcrs950eDfEX2eiJbPg5ouOTwlZpOSjYM+vU65
tlQCz61gHyVZB/t899DT3xQWa7dUOhAN+rV2QOIkm9fH9BaoWBFJnP8vx6MVWr9c
Tvy9EOfpFIFvTziwkFbyzko6jLwQmJpxzcO7EmVa/oN6tTZDcA3yXM8DVUMCrm1D
yH1wwoi1A7xr2lXw/FAAA7HiytJizW4YvllViBcB22tgivj4sTT1UGWGrlPD7Jl7
rs7ce/y+m7zAtR7a52Nkjbtg+dRiYgss/sS6ngkq28ODzdsmcaK2+luViRP9I4mG
VkqiZjzh74F9DUrl4jp92OazNex5IbbOCD8sGTShP92it++5RxXHFEURAJoSzUWx
f9DKlmTOkM2VLeohvYV/e3j5M0hwcTD3VNPz+nkcwtdlY5jIA3muyVVlVWvaMdRy
/PZD4bUvWvCHm6tRCB55ih5ahVaFBMWOKH6tQhl5F4HK354KL7/9kJ9FIMRkxBJt
oKrAWvasAeAuchN8t3Z7kBNorK+HTm2qnkbW+KIjkd/QDP1kCGy1VrO6hnQZaiZZ
xbtuNdenU7nC3njBiuhAvIG8DNtMRFCelUNj9r771Qzk8FYFzvLbwH1+h+ODXBfI
l9m6dIO42bKoG6pJJRIM/6/MKCgtzujq62GUn1yHdF054uZR3URowoE3ZhaZdE0H
0v66R2PSptjlgzcSDNMxrw1pkesQs3WVA/jHEng6WvW8on2HuiUgI3UynL0AqJHR
dZcVQoMguTXmBLLMHCmXMguGob3e2/5rCF+jc2A5dLvub6p/jUrrmNs4eHNtHdbX
mlgz/Zr7Eulx+8abYRLYlCuXCandemoxQuGu1zmntyeQmz3wS1phHWELGqm+Ne1O
MW5tCWrwFtSHKXS272XsYdJWTCcIZstvlkDhutwiI72+EF3CsOvcxrFq3QXummKU
JUF8eU+RZlKmcL5Wau7pmPN77nWxhABbHfTvEyT4trxurWtBSISSGoAd/qegh70k
YKOZndFBWMVv6UEfwP7CaukGGP6ZTEbIdYbz/h4Fg9c7zISFHEbxwKcBvmN7tZ8N
PzKsI7GyNYqAxaSmhn3xtu+pr6zO/0CnM8nofPPwROiFAoJXtKCmVRys574cKdZn
BK5z7fK5zP8YXsDwvQsYufHehlKeVfkZJIGln8s8eDVX9x4dSIfg9F4t3WTEOncU
AwCMQLbzCx+fwo5vz9OU3eMvXtbqs2MEu+zS7dMKlgxkwAUcMfKcFZe+AIxbJ81/
42KLkOmpWsNRWBHnxV2+kSB8K7esH0BCzJxssBO/mRtuAA0OZs9yPxTU0Kj/wNvB
zhRRxx+8blSxLUzFGudUSBCo5DK4qkuqWZPQKPF3//AS2G1DEr/WiLcg5NVEdjpT
4KYl+hyCiS5gVpQeUnTtb12PyCICSQ9PhD3pJcokh257tWp0uETB7YXY7s25VKrn
MzVwQtTYUMsFhWmOaFiFx0WJLPFcS72m+aFI5S0C4aI=
`protect END_PROTECTED
