`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdxSnPh9g61T/slmxzRvmBuQamOQ4WsQzpFQNh9WMOwwoXkA2fKACOMAo50Ac0bp
ow7FtHOf966xfwNJjwU/RvrQgEJp2pE+zrMMEdfkiMKXmENmqgdIGAddhqIsV/bk
lAgXv+Mq1kaPQJwnrGRJ4pBZ1NPaeqoxXVKkG3ESF4ts0EKUXhdFAOsS6b1x+YMZ
eiL//61nksEuPPgSvXr+TRCl3veqhSf/Xw49iB95juXQ3ARuduW06sdGKNeisTBo
Ohq25TJT9CN+Ci4xbFT9pfw4tJs94T1th/GWIiZXUdwXj+2YSuG+eJLIhqoVJ9po
MxxcrJFEW1z1r5cl3E5bXPGoTbswN7rJRGr6zoH9lUG/6sGBQfQCkDDP3jJsmoTu
T8aJWU6l3gZY6K7f3eM6gf50rtWMSH6mS7My0QY7pNlJPZeK2zK1NVtK7lwG/U1r
Fl5SqLz8W0zUkpUf+9hm45B9GUtgywIgnxrwHA8DNpRk67kBqYuPSxYW8DlsVJlz
9lrBquiq4iJszaqHx6zgVvHzgVXFuco/mE/WEVEvD/bigNtNilN6U+8ZBgJAQc8I
MA821SEWtY3uKpwC+o9oiqd7jD9nR8Oz5aPv2xDGwuz4nkspwIfh60Hy0L01d9lT
PxwVh8M20nFC/HLeo9vmaBl8jbaQ0VvFFHU1Pioo3AEEqtfd827mMpGhke1tPVZP
RvnCHkAu041tNQ4j7n696zaY/nEl/cdNMS9lE1JYrYOtv3Gitirxsp/jLTxsyyro
bsjEkf2hpO6GV9vdDu4ucR3FKemtDVI48O2CvIRJMO+VCF6zda95YZe4FzQD7ZvV
i0ig5UIadDUv0AJ6cdsJ1eg4XKRD80TpFwbc3k19nbjmPluFEllK5dB/3vrXwNDX
lTdKn7AlQksWzMG/JromWvyQcB0/0thVoJ7a6EAkI0srzy4MsU1hNGPlxUdbaqjs
pp+sd7K97uK9Zcsy19yLyeVRj/Po8a3SBu2u86DhrnyygDK1ADShvh1uYrBGbC1/
7mYGEYvDvMQGnI8bNYMQLcvkJdPnvS7PbF2xURQeobK+Mzf3XXIJrGZZNVnv089x
9kcTMGkH0Wz8wkSVrGU47G27pBHb/GEcGGCU+3SthLEHHOdE2aUvRf79lrP7/WYJ
ryh6i+OQJyp0AxQUMp4hHMjRUMzlEyFL1zIWWbSmrhav6tJHB4+vWNonraMQg4WT
lCwNJzwAvvsdnoRdivc8vRZxsS4Mz+FIFUuUa05FZhv9ofsuqKxcnq5BuO+SPk/n
UCkEZAcgG21eqNzAV9GBONKkg6cfG+URWV9ApPSMY4RNjxzmO0OJvM6UyPoJp7UC
oCU1uXUbSWmyd00IejkTrH/cQG2kzKNxwkGmigFgxRzUigRindyim+k+joHQHbzS
11cQEcC3tRKUboLJoRkc+ubaNl384C7SLnx2Q9cWuSK07nG929GdubviaQMA6FaC
uTo+6iH62fPBCZLE6har2Rd6VHwlByNr6Y02D05nZF29dO6ldGuxTyXlv/72812U
Wtqacy1IbMp6IKrffCHb1rnhAxui8QL3VELpaDDIS8k=
`protect END_PROTECTED
