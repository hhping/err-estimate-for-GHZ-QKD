`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VR29icvfer3gZ32Y+ILiCHfIoCdiWmR3/AMGzFYgP6r4mEE8r8blbVTlnAWDrFPV
ppJ/9mw3O7Xo+n1RwJhvEdklz5HJURVXKUz6E37X3Lb4o2hCVYskKifI8GIeh7GG
dWLzrc/9ZM94zUKJIJj5I2Oghl9QJnO6vSPs2VdfT/74LOGf66jyx2XkBZ2dQkRB
rFj8rHp0DFC7giHCN57MAr+enzOpPGEpF9JKxug8h3CUAC8ahyU/tZXIw+L+vSmQ
2sVYOV1gZocX6zvfSmS9z+POuxTQq6jZc9TTp9GehYq08YneNkDKFimojQgUTlsg
UsEaD1l+Hxlh8KnXOb05DllTS/Yjhv04q3VOChGrMdsZjpQUdGlwDURGzIF6Mgo6
RBGUVGoC7obmXoLWnViiS2iJmthc5GSYfHiYaWOpKrjYGMcdbuQedkWLt9LEwf2I
FbMU0IKQwo4C5+ERCjatDHVXzstIYsUsfKv489RNeqk3H+8G/OvhUUb9FacNawCz
vOKAMLUKrkmy51ymF4SGVRVer7jwFBRw6FnmXDKnIj4xdc4ADm14ywLyHc1bfttG
H+xwLuKAtFM52kmGRdFKaj8frX68JGHni0dNrfSnTY3KfroJpUlCJMA9GIiyd/n+
pyB4bAukB+bb8UQKtBSkFkACSOiI4rKAG3yIwnDq17kQIDYoIZU4yl2F0NsDVjhc
JmVFTikQqVYTDoQVcrqkVQmatqRjNSK8MlJfytgn4c9z5yDGOfq67wMefbFn0ax2
4Vi1m17KzCCzgjvGnMzAYnwFVPjZPMz73VbZjhcC1W8ydANAPIhmbqMpycxbZGsj
+o5XxJs4XswTtFyrASGnEFxc6YvfQqzqvyOLQd08Sw+GJMPDYivc44WO5yr9oq2q
gol8f6KLinrzC8eOjg8n8dm0gCtXrimTmDhuYzutvb9EO93OhqP3eo59NYUCpmQc
O/vYQE744tHc4NrNENmdPTKNlKpnrTJd4TN19bmuFHgZ0b42f7HW1uSv91h0tFZr
xuOQJg8IPlteVTtFZ2ksETP8D87aYUm0u35ekBYxxwF0/Mv0BuulNAmGDAg2xCgW
axzyou/69UaJlJlksFL+FnRn72G/1s6I2yc7FN8HkdHHkOOq3qucBt3bGacWPWk+
xhWgQLu/a90R8LHsxKR0sKj2BCNWf1mFmYopJvwbDev9TKXv2GynqRzy9Ol7/JcF
ga9+nWsPVzIhJZypmGA74VAAUN3JgGSYJ0XiEkJJHUxDLDrPlwZlTei5S4grXPQV
E+i+nWkgIIdJJW1R/7iRjfNcN6ZQcSuoQ7NTIlW5DF/wgRtveU+tBpXWBwOv58A+
5k3M6KcMuC5pakViJta+g6fTooCqqGfpmDFNF26E6H8nCE7zwHE5O4WV6S0wYgZ9
hrPqi8bMco67KZygx36CzC6melrdCS9GA9bXZ4e6CHaHI4c72PvZ0N517G+D+lEZ
IQcqhjJhtGLjNzlv+sds+mI/QwNLaEpGvtdQMxDonfMCH5WsfyyuyG/YxMpM8tK5
A9uyMDdzyLTKsRZhtkSWC7ahFuPBLoNBKPFsnYrEtTkdobnWAbOjowuk0J5qVLU7
fujoLWaqqz/QmAwLNUGZ60iEFgj7AtlI4GUP/TcecFlp3GJU1ZtTKT+tsd+kSZW7
mY2UN08CcaMX+uorzIqiMFAYJ+i8QHg0hiJwrkOPGKQuKNzu/WMiIEE1fW8vREw/
CpH2iwPGXRnZX4H22QTH9zyWfWxXAphUDyufcLu4dNPSnZTYHV8ixuxS1ZRSLjjA
bHe/KycW00gkz6dRirblgY+uxyV0D9rURx+2m8exbpA2mRoLSl8LmhObGanlIlGB
koS02PKE7ioyl7DC6wPeOta0LCxQgA8nTkMXCt21n3LuSzhssutIaPnP6mXQtDQ9
KcrMPIpCwkOWieOm3kXlRGnDriPpjCa0K/cUWLfruE32OJI028ExVEisbc5q3/HF
xr1QWapjZCSu8FV2q+3Msd/6hVlmlgVEvEDZtn0/iPVKg0VETlenyRWuf7b/Qfmg
YM+MgxFnBsNxPPKN2ASHiHWXPOM8SAOQRlwaeId9r8OCJoSUDkZ9OdHCX04AacHp
+0czpkOveQW/e2LkltI8VQ==
`protect END_PROTECTED
