`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PshEToBkUB0QlglSYooK3C4clpdHkHjgEQvrSGvjZnTJT+sgvXEuXVxBULf0Tp1p
aC/iyPe3WFNch9dUBP1KnWX4daHCbWYfFValwsdMR3iDsf8XQMvjszUCIul+n0pT
YDR4U1KuxbJQFneMy1hOahbC0rYkepchCWPigaZ8aejKBAI6+VsTi6Q3F0/JLLL4
IuBgWgcYT+kQ2Mk+qNqgStSSDT/DtAl7i/v7itnJ7zaorrVaCPSLqNR8c5oF0pNc
SZOXcph7oz7L5bc7kbfPErcjj64YcjOC9lj3E/ZRqTbaHHumHcl5OHBWneLxZbGY
x9u3fdoTh0fFIHutxD1naR2JnIwI5jnBm+sYsWfPT4AxNlAJHAy0Q4pIbPSD0C9m
MaxLCtwMngxOCska/5c+eDlbVVwHXMWhyHqmLAng9Lpv0nCNsbL6lokk/pTfltBe
Jw2QTvR73NAs7Ianjdvs8RtNN/rmR//5blKR95uEb+xmqD12C+Avw98EK0fKC2PA
IADQPzInGBfjXD9K0v6f66TVExlFZ98Qe5/Z9kudxMZ7wEQgY0pzDd34KisjXy57
VSffLGd4usRBO4zb5I+MmNrqQ5r8fy4CjmgcGjVz5FFuDLN0H0EUtkDaQZTGUycK
FVum7yz1jl6WNgiDqAtI4KbzNMT1YZtVjeFYXJi/U0J0WR2QiI1ow7CBsUBabnE1
olkEYqHZkNcHnM/CkJsgOIcB5tBK3xvBiXFFk3qMSCHlgSbINVvQJsIAh/WBOvIF
gXunNL6yBzB23DecFT5RfyuywyldWh2vvY2rPFoUTCNkWzHNsND76CYMCpS/qF0/
M7TftSn+3PSzfDlal7P3epjuPvhWIKBPcQoADlhWkqouSwkVCi4QvEkuovur1kPB
Ezs4MfKJNLIK56aSmr9ZB2qb242DJaBs3VgRUMpgaJlEGRQlVNjK+fu1K3Gb2sdy
kD4gTDaWo6mApIm5DgllZZ+dvtL8nJGYOK1qdULvM5oT6N79MAEXAPED+hKlWQmS
Msuh9ZSMJ5UyTF+oGt/GanoHM/l0/NHo1LjhBTgWcZLQwhb01mys/NKDssKbp+oF
koLU+mS1Tpz8agm3EtN7Aw==
`protect END_PROTECTED
