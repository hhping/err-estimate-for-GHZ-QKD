`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4AWSt36cmGl6A3C5/8x8Hd/TWh3c1zrfQkAfs1rfwb9oyb2k7LYQIBteK8Gzupe
ZOusK+YDmMLDTZU/SuulspwWaiy05IsQsddI9GvcFB2wbTrWBEl+Y7BNU+FkD3n9
HoY4vU6rkFXO1xVKnhh4vfY5td/X3Xuic2QG7OnE12jQ5lquMtlTsvmKfmpuGTSa
ebqGwZHiB+SB5okVYvEXTMSBYPS8SmXlWHh48MkYSNnahNFbrMG+6SHEKjjWaqbn
I62o7qGuSt6BdT/3SZaCPxbEEoS8fBdsqooEvTB2dCdyQEbJ/dZgG2VQ5pjheMXL
+vq0Bs4d4DGwBq+fqg1n92aCOArHusrboB05jF67BIqj0RTvXuEB1ZTqPng/EbDj
fRG2w23hhORRjfW8xm2T4eTVDygJMgtNNEzxSC/yCacUaz5V6jrPNf4ARyyBEXkA
NakCcyht8XZmzu43EFwR9S4vFez1ul1AWdzbMHDjGcIzKKxtwv4Gp26WL41xvgMG
H2sGCfKrSpHiv6ZxBdQwwfz9TumpDUBeYlClBKfju7iujPEdWpVbEuWx3zCmfekc
XcJMhZiLVX2THc5BOV1fPLSQm7+K+2eGQ/bFUJP1ya3otO204XDAucsihxpoo8RK
EGVmPbNtwuiGpMb2LHA542sWY4KCmvAP4Un6curcY0ugDk6IkayNRRNwzEVDobNT
Iqezlmji+2b5kK+H2ONnuVxr++gRdBZZ/Bps3UedNIml8/1Qm8vVsXWsWsBbpE85
xF0KLWVU/JI9syGw5LmEp1y1pN32SdzCoF1t1ZZWXaIZ9+cGaBx5qZZXddW2OeGL
oEmSTSebhwTjKbbHbsLZy7MSp+k+g1LxhlnX1W4JvZfS0Iq3Ag3dbDxKmf35ewka
cJKYmIuAPBzOG1zpko+zS3dm9FFImVNDGAEp4jZKhK1DRTQeAPK+fYcFO4CJQzbM
kJEivgLyxmjVvtuuEb3izeIPVQJzLGTZqN3CYWMqHYaRswCXL14FtmLELyFSc5RS
/5QN21kDSht547RaCP2GdJNa6St63rFbOac+xAH+GIzvWfr0aaKi0etDcZ5wcjsp
PfaRlKvnhnzvZBsU9vEuYboSasWGBGazrt4wFK71+NIkdposXEdZZtre81MNr9Hc
xbpn7ie2bL6U3ZNA2fBVK2A7by0HuDm13Q0VGh7Bdao2qeuE/bIJlB5RnsX3CWGH
t7M10iqeU9GD0SQXnR6mBLSYQizZsuTTpCQO1NmnlwXBPmlGJyvGpGMFs5LMw5BV
MAYt9NgUNnPpoePD89NXky0wvrT7izajN6IkRgqiv60SXrK/bAlVE+VObuWVOuzy
EOCyPTFuV9dqB7c4KOLKzmnBTWyBPBfRFWMt95WmaJj26oji6ywJIDf2xgwuam+i
9JcvCgSrO7ad9eNZZ/RC1Lr6bw5AZ1LUVaJXaSiy75+p9llkmQuuoCZ34WeTk+39
sUZHq84yStBO+CP4iUm4ZQ9E4P5ENHvOphSpWwSYtXWmGUr7JD5r6COGBBnd9cB4
D25ZLP9hgKAk3p0rszFWFp62mY7ZBvxpJR8Rn2WyvJXzPmChCQQBr5slJ5qCstq6
oS0tNcFak0DdIrXM2j9O4tKf6g0O4cPPQ5MC8UPiYgKwcPYarNaY3j4CYM6H0NPJ
bqJpLtgQHIc6Yn/KTc1jumYGfoXwV8qCsivuo8uoYd95CFVBEDOijZAh4k3StNZD
a5S4i0oMWE2bi83bmWdvt/Xvwk0TAp8LQWXfqqf+K2zGmG/iOloXkN8AJo86CyPO
tQKVqSdqSUJ2bt4ub9Kcl+vXh0cLG9WMrnHyRUUEyQfpqtGuJmMIQlViLcQ220Ll
vWx98EPMe+zLKoq4XYrt1srXmam0UINJN30Qds1tLRQyXd1GuvIAb/QiRVClduo6
ubSy4GPdBDHOAGcIZBm4rgA9HstWE+CIeDHOJpSjV2Wpmf30o3QzVTgo5YVjm20j
4rQNNQI5gdy/TiN5UXac/TjLYw37Mtp0BPGlVewy9hcKhFcRx/N5gnhDH+ndcsnI
XLG9FKLtXTrsGgumsYY9sy3oCGFKvs3f0Dn0Dksmi1gQL308Oxjxc2/VyobHdbSV
WgM3B5ZuqGIv95E/GoYhEjpqBe9l2ZmLFzcv0jLhCc0aAOs73/pJFIjHsPyA8LPy
6zvdNOiHUTYa+eb1VetMjwkyCLcdKfqmmltDZBxyDXQeNqCTx42ww9wQdKGuAwLu
G4asGBBIV6Bicl4COJjJ8zEi9HF3g3A3ViUd0sI9HF/k0A6bTJoiL1ITEmdR8Hrd
rcic4kwSnN3o7VeI5HrDJOW+J20V3DBNMNpG5SNDCZiQbikShXh7ukk19ecUH2iC
2D/RVMOLEIo/pWugTyHQMcR+7IaxzyNRZrj9xURcUGDM7jxu+h4L86UL+50wYOfr
F6z2pEzNlmCIZxJE4GZC5CQU7MnduhjudosHkp5s0Iagc3sfQKLSESfBClQ1Ikdw
R0PN5AcjXKWy8gu2T1C5ZK43Z7mwZsk61KZheNV/EIraFibVqGi+jstAe2jR5PED
otZo6BXoFogMYxi9pmLAh87TEnLXr70+C6Cf1gguP11DymhVa9ZI6gdqvj/Zw0lM
/BGr43TQ0E3XrE51VEotao0ChSQ25V1Buvis6ycIuQCZKcAyvl0d8yqVngKRCvYi
I6CRmPGXIm/7zVJNtoLofRxtm+0a5Mqpuln+3X1zX6pxf5R6FYKsG5kdZPWYYnZj
cFc9uLPvb5sgvyRkTmBf4aMmhot5i7ZYibt6zqfqHEvn4N74Te60HuKOoMLwiTiH
utGRAVHw8XM5khoDVbp6DUVkBjsXeGbt9GgEzFdKeUj2PsNcwL0Xtx3dNgeNF1Ck
8noY+x+yYrVsZUWRBRL1s1GYoLbm30IwxBFlkvfOlmVLygAq1ErywgrtEqmhXyqo
cy61IvEqaMX2poZwKPLfUJ8MqSxZ8t69XwuxO8HhoAeNstMKJisoF+dnd52pDdNq
jJPMOBhghORg+OCGY/kPBtr9W4hLS81TG5uXTTgh/UtkC+EuK5+t2yzEp1Q6TVny
RlLkS+ONECizeGzTWPeEFNAWbTZZuKIWeJ5NpvVTwQ42DBUbkeDaF51MhAytJ5Ya
D3YecmtCW/XXOdKeB90rE8qdLpT4EssIMVpcT2jibqrX4KHx6xRLugEiU3lSQ6J2
QisAopvCMFcg6XjgNDNKvBS0RrGGXaQdvFNn/48X41n4w6kB59amh9HE1fBytsOP
DZa8ZLdxDKwRIZGDrZzpZG2nPDLzByCqQql46n1693NRGDzuO8WmPPYc1twBeCkH
2p45xgy31szGeYiY7nMxoki6tfJCFqFXYAKs7b8qnROnZrxTwb+Vva49RAs6eLyP
ItiCnDUQpVo4YBeLT8KmUNERdFlAsdjOiDYDFURtIQ1QdU2E4ha+FufhS0HMou0X
Sfi//nphBH+G6vYgocAUSNV00Gke9qNn9nalI3ky/50bTYgaVAmu7grA7NqdFUuY
z/ow+YSThYmm/ldILAAPxGEbpP8bM/UA6gNVEPKEk431ooz8r0EFUM96XSp6f22b
IbJpcG8AQvNV9mr0bsUrx3lYhHvXFo7jVE2MLZqQGUGMpbWAxN+XZ5l10LCQb9Xu
eDliRzXWeNMn538VpWbXtV9OeVeojAU2qSPjHNBSewcUfQtnQEyh2vfORO22DXMR
ONoWlttT0HF+k3BHM+/IeH9mJAsQ2vpiMNdIk5nkmDgpcTTt6yiPXAesfrdEX6gp
oKiaSsVK0zNgr0QXJQoeMKdpvpUCeDPWJ5Oceo3Z8KEX9eUetMGPs1IjyWcOiDuz
VqpKLFg6UIcOWwNtPFDNlM9MrB56mQ9wUlsdryaMABs6RjybEEqHlxfUa4ELiDvP
IuCG7YQqamMxdrN/OHLZYpUBzUJsSSlNI++dd9Ch+lYWThxLmSllKXPTZUFeM05/
TolQBtTG0ybDaliTE1S3cF+2lyki+nGekxPdkbOZXvco2Ty3ZrZpMJSaJl9yy2/t
n/Xa1FDvVPUsLEvwR6qOkVvDOKwdzG8lMPwwwA6FWAVoGEIwZQ1X3w7uVZ67O0G5
cFgbA+hiRw3v8lMob8BEcg==
`protect END_PROTECTED
