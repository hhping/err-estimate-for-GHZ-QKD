`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49VwdRJq9Nq9C3+7JA00YEm9A1/KelCCz8mKLR7hrQr0AfDbeEKAYEVb40lkNgeV
Iuyp/OhT9P5fay9VGoI6qLsP0TJJCV529DBeeLYGfUardCZvGzyyX6COCzDSStJM
x+g2pwJY7DELMGmDrdZ7AxdaqIcMa0Y/nyr+Fop58tEPupV81AA5z5AHukKm/D6D
B7kz84eujLosMKnQZu4d1ojkDQ4sOwdRo4PkBWtaUvKO6PcNH7yrRd6SAl4RwYm2
oe9YrXzwfODYTjdF05WxGLV3Xl2ArXnD9NoM29h7bv0KTsHAwBPClL9iUhV66j32
TeRW2AxVB8IOhV3bU3SasJR45DeUh2jydK9FUX+n71GocAYktLNVePT0uMYsPmut
JKtlcQjISAMhUJMhOiwoPlcQSwm7jaIjqDdJsoncIeoDI0cfdihDuPxLwKehWctw
i861APBs6QyRyumeAMPphQPb0f85YaGvFuPXOxzrOgT4OfOU2Mg2xsUfsYwqrCYe
YWYgnxCixDzM0Vh4etnBOk9MqPLjKqBPWHDbVJG6NoKKXHATnJXpTCw0N4JcUfmT
JWjLNyTRaCbbRYyRItNbcLmifrDrxvagrvSrlbw1+3cnqFGuh25TlTAGunHp7Dyw
JFDx5FkLPXRHeovq/orLGPuYZrNCdLM12iYpK8PV9wRvd57vLu3g7DImlktCXnJS
vqxzt4ggqFU+G7HIqFXLeWpsHU3NcrpkdOQCk/ih2FWOnySLHfa3yzCz0oC6dZw8
+1n8sB6a/eIqbNhfsfYxpw==
`protect END_PROTECTED
