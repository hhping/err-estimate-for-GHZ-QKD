`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlCY+NZevgvvJrr+kb5QIdbNZ2IXYzSxwKS/Pen82fW+xwuuVMvn0LysRlNCOFYQ
NLpfNDvqv+D7L3dBhYeCu3aoVKgYN47qCL1q+s7yRJsPjJQ9kR0DE3E5uuZBnPQc
2w6TaicQ1B18dNUV1Fk6vzFWR3K2L6HFzdOGirsO5mktgtwXdcv6dGGFzKXHstt9
E0Apvw8UfitJezZKY82Y/kFiX3sBcGsifN5F3L+zAo/OZXPNNLh2YvKNtACSbhuM
v4BQ16HhnZyMo+j7Js92tGN/AJpcoTT2xrj9vX5cwcTEGVRIikjZ9SxfgPa7qGu1
OizGhT0gXGRahwzGl6p8ACq5mfO+kZlciTjGee3hmBzdQDgggPBfi+3PSPfkMHAp
2PiIUHkemva4Mez9rGIdF8ExDPdjbIBwb4LfHXjZTz62wQiYkYxIJzTIYApEcp+a
8m85oMJvYPdjUfcbXsEtKn8TdFAyFcZiiihU+hSDRz+HDVHPgcjDadH7GMs6ioeR
2RsWayRwDY7QGaGMVUMEaUXTCZPR3X7aV+rxCgtbtVlEVTGq390JZEBW0/FRyT9l
0v8W07AbAIGV/DijakIa/1NTh+zTeGxe3WQQ6cCUxUFAFlfeqwlQgYEBbsNnINc+
pGQbk11X/GglilmXn0YCojCzSyadpfgzTAvhNjFarH26wNAoo1/BCOFGR/gqNdSz
sxg91dFZwFj2PZDfHsEuqd2uEtpNGlckKjoKbI9B6t1TCRMyo8PI8z7uUiBauFxU
urMsGSREdHIy29fhkxz4lt02bCaoow+9OVADb+X2CBZf1tWjTvc19HirqeS/xqYE
58tPLD1X1KPUu1ShQ/V/fSDgt3N6RtlVNftIjS4dvV4C8Pdprsbv2U1c2njdeWne
hvDRfZjrgfvnHqQhCk+puOg+A7ML6s95HUWo1GmjJCdJbF0n/hfGxhNV/lNKZSwc
2tR5hkms8P3e4j3N7O5kKvqOdJC+S114CoCyQtYMEJ0I6RfIQgbxwzuqkxWqj4Nk
OqAoU/xlMxSih0oq9rl0eWGeOuyzLCRJvdzXzjL3OJkAWyUoQ288nwJ3wuQnnmTb
RK5kWIlRQV3lCoZKHs4AFeK9d9lvxAK8oYhhR/XvXW7GxRBu3cUQzin6pax2ZMxn
kzseuJ31OlJfm9nGub/LB90GaEGxOXjm6sylo6x5hIZ2rpYBOjEQBLMO3GUFifoz
ciVL2zw5e24Kx9UDMOWf1r9pt/Nl805FGilvdI+glzCAofNZql/DEpwCEJcDKeJq
i/+bLZjq3bifX7mNtVoEShMaDctJd7xLx2cqgOLp5uvvS0dEKy3J0BQhbkKKC2BK
+Cs5sThHreFh3fH6VQ3W64y1coMe1knO3X+1GME9f4zPTage8S6PYzEjRSfGbqlK
geAYovM+om52cQc3SadbaH3g34w/is19j7yWcyhRFguZYHPTfMRyh38zcWSZGx8Z
+xujGEEody1kzm6ZldCHsvEtAwmAxdTlOnG+0/yDPUYwAk25lTg8G6d29U6MOgQO
tT8xNCcdtXZMlGD+wu8xRyGWT00AGzkcZlotnPOGc51WMuycOR7BC1zDq/CrgUAs
J5jP8TfYnGCZEJJGVebvhSoXgpE0geYQjOjHitZwGlt9dkQVF214PYYtu18GU0em
bdvZTBdtC2ebYSNUbi9u58yLwDcwBWitQXeFspuyFpP+O8hr+Ezzp9bGXU9lWLqh
/7DykiKmptBiiEPzGjmAV7VMWafT/GIxvXrL1+4G3q/PT1XdZsWKn6PpiPaBIUoK
8RyxoqZU47LJV8bruogK02JFzDW6YV0aB84xFVK9IFcWRc+N6qxBgbhz9EFMByzz
c9IRotbxvCnlpZ5KGhVtC2lPtTud+9ij88FR+y567viAWmJXRvjhyOicpsLhW1Zy
vmT8T2UFQ6TyykbjBd+q0fUnq8s9CoS4wmXYqtXD0BsyOcZ60S9nggpLzn6WUToH
wQ1VLKz0KKf7iP58gGjU/1tF5UpwdzNLNl26YeRh7WEgVZNiv64/U+9cK5EKPfCw
s1M98y/7kX8SW3NacftZBIeSj02vuCc5CcTsr4MV4QDQfvCPwEbGuVdQ3R9v5a+v
iMiC0XO80CdVBAgEvmrpjgLsz2GGc/ZXVmP77L1VuQWpqssdePu0ECXAiju0DUHp
KytmfeaJr29mmKduh8oF8hvgsijSVpo77OHnBQa2BvHBkbga+e0sJJajcSbFflQt
5iwkEKoHWbWH1ncidobCARvvSAlD61UwjWO0WHcAM9A0vISk4zppl9DJMR/TdXmB
e1fV5TLP1YAnTdSeP03fGo86Al4gXrHpxEeDdz1GTIwmXkjPfwrDFJypKLTUBZ3B
E5ihx8arXp6uI+i1YkIOzD7ZFpp86/B4m5Bnss2Oh8q6vGsP8K9IXuBCYza24/LN
UIZIuw8JKJxqpWNk1/I8OUnNYcykCfdt5abAa4J8RX02xSUNFTVGq5o9DPKAyDSz
UAao9HbMVTx3ZPE5TuMW/QGvaSH96cxU3cwNZ1ZL/mjqz5gR2MxAELZ2CB6VhQEk
hdNYQXghJNJ7Ly7qBm2OsDG28laQg70ZgT7Ye2ouoME4LVubqpr66p9ArjQO3ASv
OaRcvmkKKe0C5ytfRyWAZx57NFuTc6UyZ9MSnH70r9kqtfvx9Xp0mEV9c93+V/av
lHhs0Tx7jBu9SK2RJiq3FxpHEqpDoH041cfoC3GsNR5mBlLIw2NDfnfJ0a90D25/
7ts7D8exD8x9LiYqHiigpmlIFF3aI0DVzSMOlAxHlb6bvTk8+Jo3a/EezEjou8UV
7CQ22mvnlkmbMIXLDA0orEQg+0+XwClcy8jq8bNFlPUcAuRrX2DZbOwi4lx7ih9o
MioywLKKWkTVt9i1mKXlW2vRYesN7RA7H6uJDpX6CiZp9jjQpz22I8q/mVox1Vue
jQ9nM9/bSITOqdeXqSrZYZyNTWcbuhUZZ1wEfXskf91M2/vtmokA/Pcpn9p8/AzM
aq62yFl4tr0PFyz69DYwDDRDCbfTGmeq0jm8umgIMKEw6ley1pPn0lVQyD837ASz
nsPC6nDMeNmndgUuWhSynVgpZlNdYPDvg6cSPfBRts9urFCGA2xfRwl9CnRG32IW
ENu+IT71PRGsDYv3Rz/COsWwxiKn+rc00otxnp2XmHYVZY1eKrxPxIoJpDEf6dte
3E0XdGVcb1RZALasDQSgAnBTltroT3sBkFgR19ds7NNq08MQpteSzCZm3aOpf49o
IWO+5YfHHrhzQzhS6BhkJtmMpmDxgaxTzIykMRZ9xdkuZP0oq8b58umy/gjHNXx1
ZC8S+3AaKc+2BxfBvQ1S6d5D/ohkel4w7rrH1denDI5LryfPxkiM8uCvayRQoF+A
+635Q6XGuSBty8gwTRfK/qviqV5jD+ENec9pW2d8MVBJ8HXGrfYY1e7E67Z1SEin
q3p1tvLtbGZwCxv1A6mkZfbB5yfNjyNYuhq8ar36AErzJrCv6UdCVhxrHrNCZxAY
yDMhmPkPYpqCb7hRlPmB7y+tt1V4RrvOH2aEAP72MqgRlbBbmwUg+app9xLX55X4
dxH7GlfOsL5hxydofPM0e9YydlxIgQ+X9I8OlHXliOgj0zR/ZLrY/o3NI7R+Ek/h
GDoQi1CO+1wQMWB2I4pma+s9MfTRDFlA2IMJdVKiAWYm4J2ee/jKq4x1ddFpV1Qm
inxsO9HAr7YKi/pOhNgelhnv6VZR1LMzj3l6uYK8lzdNRLSQU037mpbKIpGpPg0+
nTWi019AIUnRSZjbq6X2+0uty4svYRv10HwDSDgR3Te/SkbNcyXFyPX8hQG9+W6o
zOYO5fr9/o8vjL/0vqnKW2vg2qdm3MipzzM/48OkOOD1T78+M+tw3DROO4Jq7ULM
HYarFHEFisC03o1i7NjXmZr+wsFYuZNDZP9Tl5A7YWNIIoXZkL55KSW85O6UlIib
tSfwmLH14jA9dv1/3RLg3TbvgnWzG8nvMBUONvRw9oOXHbjv2JGHPEIxVP2ehPDM
IGyzluAAsxUPePnxCLh7bMcOwfGHJjzMAOcrST6AAqbASCipb3ZKPKYTnVFHFeaY
IIxteM7jt1lp55is8PVMpDtzel8CxTGsxJZn0duqxkhFAu6L3xH2OAue3BiUk7aG
3w5dF3f/S5+Zqb4bZV4nNnOl26sIWwGPCIdNgcA+GbUwMzTfbXA1xmAnYqt2keRA
zZyMYB+oiTGRGQvyu0RmbVmQ83i+XX8tAnQZQL85B2o+0lIdIhnttecPhrAbQZdl
S1ifPkLK8HwEzohoUIlq76JXlLc6XUjALINLZX1OT7s9RHbnHnCk03N9+pMKbgtP
Pqoa1b9dHbpaZyIpj3a3YpuO/6JlxXqCNpivMVMxIrvSEfTmbLUa/8yQMXMniCWi
zKp2olfJghK4m10EF8ajj4W5ARspTuNVTVXD1u4X4L45ZWLf4YhGNL+n/2Y8rCmf
ipi4iu5yv++9GCAkO2Kya3Co5nHImbpYGpD01unM9wSlfbhMHc6n4d8pWHir3UKN
HwtvTuMDjGEbYn7Wixh1CQAiwbSnpvwvPKk3HB98FIPTK8/l3mAF1C5uwNFl95C7
hxg+5BFgWzuVb39LqC7DldTzvoGe3l/vvXrWhDXxR0w6VUrsA2UfjFzZ6dbzprzw
i/miNfJh4ZrEN88Ig5u1Fx3dx7eq2yYF+JnA5bVEoUlhNkybhkwOBZhQWZFpLd3t
ktjWfXOFv/RlER4xR/KmghcA/6GOe1J1LQ2RlAiEtVGMdntlxzed3yPxpAmdxfWp
KvKqJaobliA8lDuqA7urM5BxtEOqUG9/6/I5rrw5Xl83DXdbTFJPhBFvp8FKTDPA
iFlSjEfIkaGgJ2aZ+idiMce/2OMPawXs/uvEfNQl5y88MHhop44karR3QPT0Mkc3
rpX6hxMlvFevVjPmYuBPoCMIuAWyoXtRPttq7WI1mruYPmpf1RTOZs8SUxkBACnW
d1Ia6l1WgTc1Pzx8fVMKiTBRkfsa2+N1Cd0UeQNR9syT9ucsMcJy3XGwYzy6QX2/
x4SdDrRB/P4XtWx1sEQFx16BxA/fSdDKuu/bRaKsTd7Tb0om3yOuBFAtqSQAL2Z4
tx3oOnN/sUJINR+f+3vw3juEmGqImembZ2vJHf/jqO5F7qBxovC1g1wBaypW8guZ
ZdmdXoW7kVXiOlst4cUbmC9pSxmjdjfrFHlSZerwBTgkUU/PDT4i7km7j7j1eCft
0yA8JGWorrU65WBvDsSWKLt0Ryh0i07EOQB4irD1RKzKnbSWftOrr+ZUh9ubNMqp
ynN6A8RnBE1+k5bw5g8APg==
`protect END_PROTECTED
