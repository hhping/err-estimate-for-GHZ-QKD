`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hu49+phuUdjBiCH2DCOJeWR8XD0FotF7jRfDbmfjoz+8VN5b3sLajpuhtsKx537f
gxLw7BGYnEPEYpkuatVOdyAG/myBKZG0IT84HsxEZdJ1mJ7gUiU6DfbcXmHyxQEG
8zY4CmKpWmj4ysXG00mdtzP4iJArsW2kgBVPaR000IsmkfWLlfGUNtWBnSTFQ0vw
odaG5rkH7UzSA/JOy6HE/6I15DfwwcSGUtiAc1+cQ1gjv042jlJd0I45sWlNT9Nm
cAqck7rUYFk7G4PoRg7YJwq1kvqm+j5br7oaZPpyeYGJuUycl40meEX7pD56ApzK
ZT1d8zWu4QMC7qIpa+vA5DXllmCtCC+0fUqmXwbB7qAuuESW1IZl91agj9V9Ju3o
EC/YrceqMsy9yTZH9NYkk2vGLJUGI3cfKW76+JdUHwxOtDydeakO/4jFQNcJ8hoE
ltMy7rOb6XhVGhFmyHkdcGPSwWLLWZ2Z3/3aqEDtL8+0mpxzGu8n86B+iAP0gqX/
PbG7uLZ1jaC5QVpJ53DaZaJ3635Hsr1rHTNybDuPyspJ7aY4327MOGUZqHvbLpl9
6uVnRicZ1JP1CByQuJR8tYEEJps1WOp/FhBAtyKu0RDp8QXaAM7RTEuWpVGp1hro
ysSvRMGULVxO1SKq3QcoEA5cpwbaFc40rhDR22LEEqk=
`protect END_PROTECTED
