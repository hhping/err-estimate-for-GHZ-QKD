`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpFL6qdmP13Db7wWhEQxBxIuZsa6s/UVM8+uxoBBqmICcG0gTycDyp4hFlYMTHPW
Rxo4l98LDiKT8UwSIebZ4e0kx3yxEA9XXCTxy9+ECxP5WQDN4hNn255ey16w4M87
QRD0qsr/l629BH3CDxbXTCU73O3kqjnVd+Od+Nc64NhQj5S0bztyUR08pfaxZl25
2M65dpzbo4eRCQEWeazy2RbOCQDYyWiP/h3F59LqgWdUjCkVbuxl57/1Ofon0gnk
mDbVmGOC2kekiIkPGEur+C+HxgKBgl4Lr70bo+8nEtN8PYWQMTOIKcUWTtfJroMs
tEeUx/ecYgQINsoJrr4/f7Gtd7vZIdUE+Xtb61DXKUyyNxjCrj9s3/vbpsJtcirO
Vh7WoSqduNer1SKH+VCzCxNQfL2jDaQlb1qzzZQ+jGtR/Y8xiTYFHgcQDTMWAC0p
XoUB2WG2yBlvdIyl4IucDBtDNCpVMhO9qXDoB/yz7Klev974vX2cmaD45FjS/Gad
dgD5dXsbtMEfd4RoOyWHVSaUnOnHgUEiurBoUuKc/3B5wHc9UTXyS/ufVe4FuxHI
eS6zbAEGiP/OJf7LumoeH33QuMCLGgQ3MDAbb5TpOOhLXREX8gvxUCpjW6V26ATw
IUQ4H1sZhx2vqQjzul7wu1GJrWPgM9xWzfhvmLIy0fOOhTxHR5JXUZgIKqJh8rzz
DkO1uNVnIlQwn4m1bDelqMpDg0IeFeZr7Md8otRGmA1S4CqFOXP+cRhGldhoK2+Q
VXdSPYP3xgn+2gHRf2B8r9G3aVMcGg6Et+2kQ8UMSupfTq1oT4+V0xg6CfCqgNU2
hzAhM47OYUqWbTMZiPZ46C52cyS4N5T3kkDZKYHFvGXe6Q5pqyv8PkizsB0p31L5
1o6i9pRQ65Q0srphokcCekKl76KUluZfRkK+V6CyM8OyXAT61SCDqkeZRGopOBTl
5/FqCMOnT4jXVxpIL0RUqzYGmpbZ+SjcqT2t8NpLkaOLeGDnZL8+xOxTjF9uQlMz
tYFEFRa50XuSDFXXqwEdNr9tlwodPJCcRd/8rUEJa7IktKn4fMRzVjvlyVizKQyj
x9R8HGls3oTw8bHVUrWNbAz9P7H2kdKsO7cMjknhOG++LnIf3Ss4eTPW5ADSeu4S
CScKY7Diw99izaTT+9tq9g/ryMYpN5eOiLB4HFoztRyR+yqecTgkY0gGprDLFxVk
ktTB7E371Jaw0DmsWGcqzqIz8xaw4f0Zs9WxSJE7aqOvOq6yZD9RNEoFsDIy4fQw
jNagaiAq621eGK7ez/9MAyvehi3scS3bB+Ie1pWE47EB49nu0/TF2ogjGjU+VxqH
rQflQX/ONcK7xeEONF/9XZwR47bWrKZj3PToHpO5vO2fhCRaxTdl4Sw59F2TPXAA
0WMDvDEua/U6PUfaVqcHuw2Q8jnjiFgPqczYJZTlfMUMYKaOPxAxkrRDAjWQBor6
DF+6ONIZmzv8q0BmKgW9zaftRyP3gDKEWeoNcLjygASqO73d7W4GeaDsZB0SgJOa
giH3o0QESnpVYhHnoyIK/lNhKa8WyDYM3aNdA+i1EY8=
`protect END_PROTECTED
