`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXlVB5ilHmaKVRr743m46F2R06nbDXveXHQp6KyoVxqCR6Zq4oMCfSZsdDnuzttr
toGg1T8PLJcbJy1xc2CsLtfcQqQARmQOltiLWrcRWB33xDG7GSxN4GnhDFKlfQ4K
1IdklPPbx5k9fUq2iEU0PKEIveSlqw307O+oixQNmRFeT0Rq//kCCEeGgQoTwDiy
Ff+o4wl/ncwBVd+c/ot3WzS7TWfInjbnYrV5tXJQuwapWXuq3kk7cO0RypNozC7y
O82Vkp4+vbc9/JHivhm25KRfbpma1tCgHm5XVz5snaeeKwrxgJWKXu9gKMaSH433
Wm1oaxUMAh3ZoOrntJvDZUXHkkMwghxX4LHRW+58J+kqAMEcY9Y48crzR+JZxNex
f/HW2GIsqnK4hLWA3rxX6BqnXf8Hb+YR0eJfqIzphg6u03MzeTtlvftKjMEAh5Cm
InaV8ekcnsQZe2eKdg09UVJQD9BT6i8cgAe9MzmEVYQTptmnP4IG0swtk8y1QKs4
kd2IyzFNfu6UN9CJKAdNSTm17PWqdQYe1gsSU6GbIVbsgdDnth3Wuc6GFIejXt75
rdrD2z8CVggWcxIqqm5kWDbOMyJf05UBILmqYUGyk1xTMyokuXE42RKwGSdASgJJ
VTMZXgVrvCvv/kLljmkWRN+g0fKsRbQCDtJ4XqsEsYTx/F1C6Ls238peR66RWcww
FikwUr0vMKQauHh/KWRNo9zx8Icp04MSD81q5qLRoDWFWSUUnxArZ1q0GSE5aOhl
8uRSC75mX6hWEaMIdiBiSuymjcMHq3UHWJ1lnzsS646byicbudRbNEIks2L5d6fF
`protect END_PROTECTED
