`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpxAxGDcNNUhF5MvyWsuXHEaOVSZefj958czwIz619V0jB5tCD2PjWmaSeTaK0WT
MkKARoCZ3reKt2exNPTFoMjFV+BevqOrV43krfenA+h50WA8BB1UJ+Z2/mlgSOho
J49fCAVR2zGj5YK8nauBddttKDz2qMUAO+lWaY8+5sDzt+ia0ss91axt/LohAf7u
O/y2vnNs3T5rzG+kBcRIzK+uFSINT9HRWQmWOIKklhk3LdKqmOl93El4Z0UDHRV5
c881579u1ks4ke9ykEOYEwBGhBvQ/2xdvFhyrN1RAMDb849Y+tQwClOPH9kBspl1
INjxqA5VaekvIYE/M+A3h972PsD+SQGf/qvlOWmfsuyfl3xgsFV+6jiy1twBrAgs
miOWLzJjy5VziNywU2imH5UHL9a4uWwmbCsGN2GikUeHAOIMkAsENSDbIcl1iZdM
WmCMXcNeByGn8O9k0YbOTKBYTeoAg67V4GSG/QV1LEUVJXi8UBTZ18dQGfafXrBb
WmqAMHweAgMAJa29DL5IwSri8+fNi01d3QsbSuAvtPPgC8K+CG81pu/ZUji4JeQg
Jx5UT55FYq2dytW/TxJG//xe6g+SRi65NAJgxjHuNKZ5H9pH1I5D4wPM1XzK1Ia2
fCJvP2qP1M6IQdPGZzPEDhM2us+TeoGSJUOMCpydjOcnibLgSN3r/Q3lhapH+Foj
MaCLn6+7fW+9CCZODv+QZWkiB/o9PqHZRqSCC88n53EDGj85zLu0ncbHroaRSLe6
ptpIaQrJMKh2X9dv3wTAnPimjxhvMeaMMRawxPMvvH2Xxe9f0GsrhvjI2JAfrsd+
bVj/tx/XSqTxH8COtJmn7PMdIbPPNeb8lFOCrL4vH4wio88pI8eot8dddn7Jgf2M
MBHrTxu6UTBzbSbJF6wA2s2BmNMUHrqUvK8heS6+Ae3wSfwggkHec0u8eE60G1pX
rKCMP1SCOCbG0NzlMzIJf/8XvdMH5doL9SGMNhoTmAWGOnxvdhfv/ZuoQdNWs8iZ
XqF8a0l/zyTTdFYfIhbEdbh8aywRD98CVnbWpsax1OoulON4HXudOWtofDtjBMzo
EaBB7PFMZXecJf0rVApgDyOLlEXGj4tYsbPJjCHQaBzGz0R2LqiyLnCzq6SX6edl
Zg30AJ1wZwyT2NgjiyY3zN+BujZ8eOj1nYk+pjl8GZMjeQ6q2mo5rCu795f4ofFy
hkdswxe2XkuROOUosJ3MJfvLMRXAEMSmJz8Vk0ScYjp+4EflxcHPFpgHLSCZaSPK
VVOP9fWykkJDoX9JFM4cJNN+DrnOVTO3IdCxSwjUuKPLzgM3mfDJQa5KmZKJv43c
JIOAvSnowsWMUUa2UaZ1A/SzBCWXlAC91fZsdBcysEhKTdLEYV+XsxCMzjWY+pPC
e0rGwaI4usSm3Dx1ZhGLjFwVYHjEdp+RTd/lKgORTmnk3ZJ6OQr/ayQlu+oHGldb
lDpOHghxudOEIAznU9TgO6DX9iAWt15/HBUc+iiD2yaGyBvcMMLHpZWXNfhUnLew
z02q4ZK1tlpDbti7AclkhF96VJVgClJT7UwvSQfPwy2zJ3w3CfBKPw1+h2qk9OAT
+q0Zko8zlRctHOqIyGPdihFFIOAOGBxbQg1sIVv3quF2eT2Mk+C5zVzjJ7thtnhZ
icK21OjIWocg6fnMiGbs+SI8jqp7NIUUVLxJYfOsj424T4fpOmy4IssPbab2HyBa
hkftsdB/AwtuTWdNigPaeIHeAgydXjLFgWNubFM3XaggOrwAt/YCxAHsk2zte62l
iRYObOMZrAxISkyOPuYBhngJlw+i9SalM/AhYQsGVS7MOMlHb1UCe+Yjp1TmIs+I
i4APWwz8ZZfsHyP0eh18+O9boHFU8VSSU60Y+2S+fKh6XyecRCDsq/M0ZSmx+Qdr
lvnt0krGfQ+wNSnHa8CYkyWRA8Jcj5n+tRKkanPzD1stNCunBB4ZuUsMV1tXN1FQ
TQ3POQ54qu2ln2NiiJKa7j56dTEH2Nw8HffZh3HHvufO9CwYGSk3RQDvH5IDQrdK
xv+riK84RBASGsxJyewF8sTpgB0moUNYKL2ZvnGNsRkEnN6oScc3WvxcVDPhttjo
u9gg7eD2jJYodpk4V/wIQZMSG36oh7lSjN0OATWbLDCkgcQ6m2NtipPwuHbO57PH
b0budya1s3bomuq2GOtZfxirR61DWpck91gakNHYOrwEhaGKWL8nfOhyTOVe+Lwh
TjWg6nkR4zMnFI4vFibxzvjcnU8prPUEqCs9Diww7udiYfUk4aXT8Ba07tBaP/8t
GdQ3d09//X3DU64nOMhkUtuRvBRWVZ6VlmNf0FJgNT8G3tA/Ym8OM8RBZLnm+5pu
P0yd+Uh5xD5W0yljgXcjKNYiIIFj3O/I13+su2hDsBPcc4kURpUpvOlEqlPmRB9b
YdCsfzSSRLxXlgFniBSjoDLpK4kKPDVRKcsMbIx+FeibZdDG4eRsVuVaAQR5Wfah
CA9tS7gui7p0DCDWRCHH+hPmDn6UTpwSLI3rtnPutkfAfzMwQm99b8CUpWY4ImW9
QS7mCwaCBN5ZpEBiIQ4icI+hQ1Us7sKvhYonvROtEf4M19NFwC5X/9THg3OcGR5O
ITwTSuzi5lGEcIP43KcSunlEzJdwnYl/sdqZxhllysb3VL9T5tE82Zqu5mIjqsGW
7+UwSv6ti3F0UfMpNZsOmNLmPCL6hjjamJzd2bqA+VVmb9uxMTwNi2K02z6OzmYG
R5KpxIM3FcszmBqpwqpDpcaSz4cM8dKtJkuj8WC6kCm39nINkAEJCyXy5XxgZGjs
DeXLOGOnyBIb0mgol+Q3qHqrO7bTUQdN5HT2wH7dmFx2HjPqF+qAT+sSUZL62ENa
DFfbKbvA9WPfQRL6eyNBbdau+/lPH+V/iknKgOp3Qk/SjGSM0ukZwdj1UxJ9k7nk
5/qWWA4qyDNjb8H1ybZ3kBm0cABII3KocPOzbqobuwZUPZ30tMZS0Lz3EDtY5tli
J/IaDEVwQKQ1nIGVR/Tmw+58SWOiZV9eq5D+Eby+gIM6Jiqi/nM1PXpuA6K/T74i
y0bBSB+GKblWqhehZCckpDZJIHcMSxk3B96KDItYxNH5uHHDoBCI733DoJhhDto1
wFCWr/9LwLuEXLX6VLxtS/vEGEh98DaZ8gVS2sw5F9Sb1Wn7BUh7xVZ0QkLlqU9a
ra3CyDGmnGEmHCiJeqtpEy4sc1nSVd49v1FaouDFCsjIg0XcrqX2SDnP9wPfftF+
RrtEe3mnJ35Mw0SLDLr6ACs1fUP9WI6PWx6NCt8JIXUuDYfDDg0edZlxNWwHQ43h
MawABSoOfaOIXIwiz0NDjH62r+jo/eU1oBzqBsXc3ioXLGi8W4F9n7cfch2SoE7S
c9Bnz2Nznl9jE3GTn4y9e4jljYl7D8OzrTAb4zjj6uh+qHlwOGH5oqozN3NtMza/
0XWZUe19uNQJxD8LaLvMTttIUgIO/RjiUlSdsKm5Iv28oMZcDEMjJrccOwq5if1J
vBrqe9eFOdYIfvNYylDvTxH7n48t4VpWtn1wZykrQ18tTVf2ltwhq+gonQC6epJS
dL2Jb/ENq+/rf50VsDLB9Sz2wbIL37Vq2Jynvn3/IAE+kQ/IWZP2GtIHj5wT8saA
oprbvRteB3RSj9Q8+ZLqg1CsRO8kaGc9rSS/yQx+JGhHGXIpRIH1WJnrPmBfVgld
I5ouquj14SEsrwrwIgRb1GPDL+raRzfJXKhNDyEDWBZEGJ0bu0qDaKG9zxqmaiqv
OJ8U2UjrUa2R3JlWJj1S/EnUKLNSUJqQftibXb4UHmRipCIow8yYH7/Ep3uA4BPR
7VRaAs7OGnE1sLLWLX7kVREun7/nK4ZwGkmVSL/SMamX1910tgrkEsFbvgPWI+FI
uFKgu+T0mUYq6yldvz/y7cs1O/vtnHzn+BvFPCDUVkbTQapwWl9VJ0A2cBUwHJp+
wO1OBo7rd6wCBVQOCTjusndfPDm1UFG4sDkQDE8ZrB/LqZA+MbypgzOjiJWwywVG
it8aSMHDw9Stk82w9i2LmWhJnxRdE/9IyqrsScXqImjNgk5o1tWW/T48odM5mjKh
iLvVSYtEgjh+7zYAOdPp3QLTHXsTfOxQ0cROTBM3rrfbJ6hOVXm/0OLCBuk9eCEk
vXki8V1lp0N4IOJpCn8R5gZ190RQEREroi2kk2wE4OV2UhVYfZCmzlPjzZeBpqRl
0enb3HNB67tjNGoljnwqlYWaaLA9YKmqpGdbhGDv6lWBa1ZeY4+4MM0/SB++XzH3
ddPG6numjCm0OKkzrVogLguMNSVMIE7HMa5FQnUKLQ8pEsONUfkge6rzk4ubt11i
7a3JbuU+lyvdL0ECIPi8t76IxGODvHcl79hYqEUf9W9LPDRgEuKp4YUo8Ily1fd6
lxneWEwQ71KLwaoFUlGemSnMygk/aY4SHLiMOQUipVhzgZP86N69wHb2l0pQ9qtE
HHBJmQeJ6ifKlLIGMZ+qxkI4xL8MFqIgI/Y58G2Uv+VbhyKbOVL0F4UwpJAyr8aS
Q/uqSgM5Jl8YBD61t9809Nv//HSz9glhBEjpeIwWYYxfwzlSVEW5IIbCTV7a3CGc
NHW4mwjEe0m5+fE1l1iaudyL2jBtTqi8iZXs/jieZQ0PQ9Ldjh6rlvoDDmxEi6hq
/B2M5/tQRSUknB6H2U2r685OEJTS3q/7r/buzjRrKcXHV1CXCmlBfzKCAdf0PfrI
VUY2LpQO9n72EQqK1DwWzfQ+tIWVKzR0GDvvPLHRY6d8PkSKvWw+yVnIeJ6xN3j2
dRxYlwe1sLSsgWbSwsYW7QytlSrHOHm2Rl3gj0HYainmVWdB2vK6FS9JPrL20X5V
OxOUbRPBGMxl2QlqKaKC9L4InxC/m0tiSsRZaqNIBlHSBZtKq5KxiHT8Nym7G77R
NN7SIDCJq2opl5aXhWKTp3kWR9tZ/1tEY/CdiJG9VtR0hbfjkbiE49sALadHGgi2
PlBx6Ea7QbAiNDSwU+toG0bjnQSN5L1HbZBMFOMBgRkKF3VEfqoFOpHWvVTFFfsW
80xfuAhP7PHobcf3ZeMXGIq8c66QBJZoZadRcg+yZPkJ+b9d9ih0FuQDGgrq02tU
Xs2NJ1cXPM8Anz1LPeKGrEhfWCtrXM9tWZA+Zo+vqWQ9m00rmPXhihakkTulHBxi
6kpfomig3Y76hpc2g4kn5JRfRP95KNX3Sg+WLfjyTIMeN65W3menfd3qPtgVzg/f
xpyr9UJgeH2/BiDg3z5wYZRMnjzOik4LMHmFD6qgkhs+MjvEuqoQSeyHV4CxVJ1t
RAP39SAMEYJu9M4LlzIbVhM7fcDW1aNbeYfEAyoPlrirfk7GbsNYwHQwGrbIKjW1
coTGtMp/jz/EWuXMn9BOi5m91xYlFJFqdZuvhXBcvsNC3bIO7mUW5KGWCA3adfy+
aodoZsXSmmk3+yoncVUC1eUeijbLrfdaGvnenXeueCqXkwpjFWy0YYqlWeYdgzZV
XFETQq5aDvDwE5iq6n2yjNTBiAfWQ6GZHD3DFGOaIwqC8IXNBJbs8g8aCU8PcGuf
UJfUPvlkgByc2pcNp8sTdSfI1o3KldmVEnhW4KhgUff78teXB6m0Uy82TiW18pHY
c7vBTMgxCae3G6VawzcUWO04SIGy13s7A4BEjwTRzNGBPoKyNvrKWQ6JA8sXVRDU
otItIWIZbeKSO6KhFJguN3mny3t7A6BBRBNRFOAI5wKmnTHnR4WWFLm6SH0G3VeC
NsDx+jk+lrgLljliAP/fOwyNfCzf8aMtKl/EG6rBjHXC5B+SuZ9vgWpSSYDvae3T
n2EtVm2VtpCelF18dJiMYlgbdWoEL6Ss3lVdgcG1RMApnR147t+F0Ll1SOTS+/Wd
neYq7XfGh6hsYuS52V41nhg0H8CGodFtA0bc9PLjfgnHKMUQ+rxCvfto73CY1ZvS
cxMu2PnGrtd+X4vIgbsDIYWZK/Paq4Qrrl/DsOx8fRh2fvmfRof+hJavusjotuyM
sEUkSdLjs9q4uab3O4fguOysTsef+dWRiO1LPZjqWDFjL1n0y/qG3jPgTZQK8UQ5
uiQRLZtxsHY82p0O+qLBqnNixwXzlqTeaVUwhM3X/ZQuGPWAWV5oUTeaQkF3QxRW
4uDdMoERXrZUDEgN2qkJmNK76x/aO++q2HiCJvPEyGn40v40cPc7ErgZqBYE17I7
/KLj2ps3aRSpYcdNC8Q8qC+43JYtX09JT/PPQrdH7R9lk/rmMFa2bFCUEecOvbJS
X9qsUvf4I9VTkZaytR5AqjpbIiJj8vPz43a/cXEZaKRftCAAI1qaCXDvZOaeWVN7
teeRgGhk3uFHK7ogb/LsXkyYODKNiqGbF1o9/1oFtjvuLWRKtDwAT4E8LHhUCZLG
t5CfazJFHMyWE9JTdcmtcEdcyGARsaQldoEJYjZK3jAx+NtCXD9h5LAktABmg1km
A+23fVcmg8n7uofFENPZFn3fO0of68xlwBnTFUR+ZJZJ7ATonVTFb+O1iLw1HXUP
5faCFAmrobudyf/WxbEZ4Jb70BBoxjE8W8+Zf6zEX8MBND6sVnK6AYxT6FIZwz+9
+Sh0nIlQweVCXS4Z+Ra4ANTteuHf0vhEh1VKt+t+MZr4XkMmT6qT8Td7hF+Jr1lm
ITvgcFG6fs960QgdD8wIYwloj2Ji6XK73RBtk11WSQUnc0xbaYiw+uDU9+kDlaq2
6fdzpeTwF9o23iIVDWMWS5hwDG0IQFbxvFIJYOmvSCb+aIsvWMRPOPmtbr6Py2EN
Lr2Flt80wgkUQl6ZMAWn0UJn1yXMMTA7JycEXO9+TqDops8TIurxhIn2ne2LAHfH
G0Rbsl/fNESTiXTwBYXuKm05XEi7AAybLqIlbRctg/C5cfeNm9oWpDD222ProBf/
HEVMLrotl4wEVTU0vHDy8dHyOldzgTPSGQ7Um3w/vM9o/EAHDfdZtpafhSkvb9LO
JjmKz4SKNsVMMne81HBRg2f+X93B0cli2OgazCYNlMZj02scJjSgTXosG1tmol21
Uu0uMJKKQc/09N77uUC3LQ3v4cBtXRK3rO6lz3LHwKmd4yzumzTg4vjJJPxUEckl
kN7sHE2Z7bb/Fp05psZgn9YB6Mz7MLWpsyUh0k+NnuD0+rXhqqiD+KNyEQWoRgxN
h29gpIhB5F2DynL0kE58sx4Eg3/QPVo4IPat07IK19fMlO3rM/gfnoUTH0QIZY6D
qcQ92m0G2Gnj/f7QqqtCIIO4fVQl2MVCZKBLFSvGGs3aDBzqUJYZ5/E2NK/+xpQH
UQZCVpcwmk+IB8OEBYhWoYhaLJS26VvmjC52bRRylFCw29GP2BVuV9ZmO53i2wck
GOmTy7tGOcIT9/TQjbvn9MXJt0e06ESXkt3VrA6Vk+wy6PfhxZna/usV3OEWsEv8
EecdkQuCRXKWLAKeWEulvya7CofTmeO47xsEq7LgF9S0DBUqrXKttAUZpA/Z7Udu
Jy1wOL7Mb1MVDfnf996OpxTlJ5RfAZ9YVelfJzBn52OgRzJVWuXfPi4dKVeeFSpM
yF2ans9UkZMi8Ci25TKiDhQu4kAJiaTHaPeI4vBCmN7q9cPlSIUPI3nh1ZkQxGWx
YQ+XFn4seSlBj7TcHINI4Dx3W+uPsteM2tDPbTtasOzcE3fZmLjefbwSU+GEM+aH
gstezpZ578nGCPsZqFfByDHYgs0ROABC+kgSElGrGlhD8yiRKupmOeEwS9JlCuhJ
J2qBfL2fsJiILpnFuRHZjRx64SKiYo0hoikQn2lwHWie8pPXOuQiMqjLXglwsLwc
cbo24ahkNoMafel3/KtwbmloIAX1KOBs+/SocQ6fiz+xpqrPjLBrT8zWHdOMoIPD
v0h5DFie9URKX1eplJwtTFh0fYlGY9eNAxHAp58IYSoue74HC1EVwefJsoGI5piw
0EXDCERMhFZZWNN+dfJ4HEdUfxksY6CUuZHmzKr4gtwa+lGEvZ30A18tZYoAEhiN
XA357c3dLacicHD9zIQml/a47RrdgqjfmiXtaJgTOTie+/XZB/CahBCC8HpoqHEg
vjM5KBhgdzmrreg6mFZmvXMOZtdRiPfJWsoPeMuMoBh3c9NVONCt+yCrKHE3SjQt
d/8YGWDQjcU5d7RUdVN4sMr7IVGH4iqYWmHE574vJt5csC+dD1QRE38FwEEP8pLF
kxHGpG7abyzhjyRh3DBAzFtEMeVyGRRHO6TSzKNo0AN8l9gkbOx0qUMW80/mU/KM
IawDstM4UE3Nzs95paQj3SBKrWSpxSzuJqbDGWT4j8tf1hRgZS/S4T0uHbanRRe+
R7tDmtaVYiivXBk61KiH47vPV2pa0WjkHFWOI2WcF/VmpvVrk/AxraqK34MN6SDu
WV015oAyzylN9bx8Y8ubbPP2473ptoZpSDfXEE7G8ccsBNbbxUv46yxFIlQT/xd1
T7TbrqCQDwg+X3i0gadkPbjHo9DQXL/YAYnAXMellfXkTW0n7GllzdkSJKw/wbzT
SuLgthCed+vY1Ad2xoC4j1F2M2+Ln6TzO4h2OZ0YGtLYPAiDvGP+oo9c7SCdnYWI
JP84V9O2LbaCH0dIWgndFlBCnC3vt+R/eOPM9vbn613ASduJPxf5p/VDgM7yoFu2
uVJq/epEFdm/Meea4gqLzcwnr3CbBl0gWIg3KQ3iWn41jz5WUGz2Uhj7Cmb/SjeD
cdWv4gm3YzhCyLrnxynQu9yHTTV0/ntevTPgoi99EN+yOELRwr1aZ3uYy67FUlls
XxZ5oIkMQ3dkNbQwHvcq5kXBfuni/dhqEElYUrCavv50Q9k7wTpPOU1AiqlBiCeN
FZ/ysYvitF3wcGq0L8yC5uwJMeVPJqXKQW9a5CeZNPoQxtMBlW2TlvUJGCRcg7p5
ftCCmovVQ1S/4A6GVFQjE0BAYZYRRbm56ep28Ub+DtavSgyESuD5HzPLPZjKpolQ
SgAoU+LB+OeypirK7fu9kcaDO4pXixj2BKr4iY6wMNGnHCHEW0KDTsdjp+Ox8z6p
moB9pk3BU16XUq93imsncPJgbJ8mav6tVCiL7CroqE+vGJhmETTK/G65DWZQKjag
nWuX1cmuv0nfmvnMfTrJ1cVdnM10X0Bsjwf7pCoedFAGnz/IltmL8rZBw7Sy0ffS
hVfn3R/yv7f/6PWOA8ll4ZzYra9R3Ah07zGQOUMgBDce47wOao3OAzLkXXGDbl5j
Or1YhVPFK7BpNREA2EMza2LpZYFUtHFky9OXIuOPfXVqgFtmhC2XCJHjd5zJMtrX
u9LAD32zyf0nsdFoT9pw6ZDrL50emlUDuxeXXUgf5lc6W8Ds8TLS62nkrKeIb1RX
BQR1S8A99WPjcfRFdlb/4P8VjVfGm4YiUYCPR/P6VpbSVO5lQhuakCf+FN3vZe68
Iig+fK8PTEJq53WiyLrrcbOt8X3TRKouj4zRzwmQidWIiG7KPNBE2/50hpOXl1+W
j7xg8i02RsAZ8v6ecp2utstxSvxYQo2CNDGrPpTY4QzcIJ7miBhKdvXeaT9j2yjJ
6Nwg0nFfGAGsy9JbNoUTYbVcN1S3g1s7T2+5CRC/wDAi84EuLCo4uqWV18dMbSVk
BIniTtZwGF7NcmAkQaHuxBwh8NE2/ltnbfoj9u8OPOVB9sNWfBqRNM883lolrqYq
X/nVjjiok9Kwc8HvKi8zGp6lSyO5BVbc0L9u8BmZNcV1Uo+JW8ei2PBod3sYLsc4
fuuwbasEfVw7T9avrHZ9GSgJvLNNw5x7MyBvGd5XvAyHIR3M/mNSAgQDyc5/IJhS
lri2WAU9DBU2OlxjwZWlx7hts+3WMYXYHd4OpX7zeyIkOXf98nfye3tf5Z9lVYYa
ipWO7k4f4K8rzFLBNx1kL1qRgbu7IONl+vQSRvLHn/cILNhnupJj0dymxqGU2uYU
kSmQmo4+9Zi85FY7EkAWwzdIGeSXnFGmd8HcsjjNk4MmpfK4mRTETcIGXVsZRDOi
xRHIfxiByvkpsqDUwbfhr0XBPFI1cnKvsFpAiod9ISP9p0p4OuYHc5LykcPmqKZ2
4C0RHcSlLXb9yPPBSAcwxxolB2E6a06/mZvfJQFXXf5ERCNgH/k3pzk2blV3LHNK
Y9fC6QY95zmD5Yu5oysdwVsofgS4J1MCgG8XWXQYD2QNlp29oHzNdAQIP5WfiOfz
fG9enV1DGGRMwV3hAz7MMsIY9mb8BsQyDxXxKeYYmj75fvm/vee5zSsYkTBhDd6T
wlPi86NB8YQvK3QdT/qhE18fT81DAIkwCLdygus7guWXmkNxjcsp0eWwLrLrn8Ay
qsN2XjaGGHtJR+YHk4daWSTSm+JCY/DQDZdQ01a0QtTuW+Z6X+JTlM6OC5qI180L
xBIrtU0lSiBrnT8BnEfKUniFvtB4FxBcAXXB9ETENcRmy8QZQW8BK4fbB3W5vsW7
PGzr9mdViEMoEhqgLfOSdgtzpiOHMO6bDnLmWmCvJW+tr0NGrWs+pgHOCQv5PfZG
rwhrtYoF09lgzve42it4gYKtBs/2k7o+rbM2fRb470Iv0YFTkNF+6RiedmUNyDtW
0Pbg+keGv474bDgnP6nylM/k/uwBsO6y2XzmKG5IwGxJ5dnv7McWHbTFWBul7nHB
GA4fS4BGwES3vGlA6RSnEJ6r//ckAw4q9vogXtkQr/FJK7U3USBgtWXYVSCk0k5/
TWX5TMagr8iZwCTb/hYSvF9HwXRD2xWcNlcXDu5Q7U4t1aSv4p+nh/CuHcANn0IO
cPN7SLJOLDgIhS1CXUsbtoqZuvLWDzodygnQnutGualtckwbqiCbtiyijLCZhnPL
++MszlnDAyDrAQWpSSSrG1YzaAa1mQWpSQB+/PNcV53ata3HQ7v0pP3v7/5b7zhc
WTAp0p0uOf6OX6Zq6cr48MoD2c+jemVUXwiJtCuOLBow3rND/gnVkQWJrP8tZ1xh
tWOrzj85DBBZVTs9KYOotDyn3EJDnijNke2aMe12MMLh/hBOVQUOAYsJleBiqi56
DvYJBi9+zJrFtCm+oMkkkKGjqC8eYtfyDotX8sx+zVC4WV8Ln7xs21oKxOkrv6my
UhbfPT814Eli7IaR1erD9sXxl7nLfhVMsgLI38X5fSdytUGaBn1PKi9glQNmipIz
I5qTahoLVJb0aYECsvhIGHbP1biz42M9NNC60gX7u64R5kUif/ZC0avIK7z6XXqJ
sAsf18B9kZ3+BvSjHJYsGzN8pLqQq4l3YUxcXTrokfs8qPTxe0B6eAKw91Z+Argx
UdDjzvMZ9R3siJ9CvE3nybpeKJc9KVAIwir8ou99uaFnYSxp4M9AbKMQ2ZDu7bBW
N8NPOUDtskYUaswwG5U2p8PbC1VMvBh4+uT1koQG09P0DS+MAqFleSdQmHNF03K4
vaAd/LOW+SQgvadMUdw5Zy7I/OfptEl+1wd9SqeS//hxm5ukSw/wiUARRb/YX8HD
6/cKUWMI8PVz2tsJuGZlCcLe9Yp6hz2fXnyxB1ldQYvQS/PxDD9gvRLbG8ayBOVa
uonUAyZQtgY0H2kdfeMFwge3hFExxSPfuIm0PQYsfmK9J+FdSSV6g8QYzVn6AmwG
quW8PEjkRvPvHiSHblD2Vdq0nJkSUbd09qyzrY6xOkWyDz/Tr4u7slt42vyRW6yr
E5nBbnTdB57vF48QF2jvklLjbfmybd11uyc8FqwPNXwIw5YvgKNNUktJ8TLKHeFF
OmeFjRNjgu8IticM+S8osW3FxridZcXe6DVLLcVlowHuQplceTQOah64V1PY6t9d
9fCquBax6qkvynNn+rIQ81JFV/aHaFeasV2CAj45qgjyR4OxwQJZ4HU7Aw5XZohT
FU3SECYKFaq+ZbDr7+SunTcT78v3QA29i2p5zp+4CrWAJJV0l58MW6RDbo+ok4hB
y8PYaX6t8Lp1mwHNh95N9dRr09PbxSJmH9qPBorkFuZKjGVe3Y5ujuCxV/TEcHBH
mY+iJH79DwvIqktICFQBSlggniM9cZ6ADL0nk7tF99uCtmiHvvnwhZQiLCMSPuEI
dWP2yIBHpn69MslU89XgWSR2XQukjZcNeSbla/MIMM6jwVWdxwNNYmOS3c9cdF2V
t+fqg5HyzMUPX110mZ08s0zAAHQ0Wx4iI9M4Ft7fPLKOjWLc2ssHOJhEG0MrftOB
kEOAUfl/sz88hVKkneGVAz7t8rixhuN7wj5YYaKxrN/zlPH958BjWMPOmTdV6fny
mhl0hwi/DS+NfbpTVKBEqFi1nLg9FY8YaMHYnXlWVwTHfK0BPlHHtX97ntTmMeEa
FCkEKK6xCZD6NR2WWDuuePzJnREhpnNxnn7cLjhi3vN45dZzNBz5GiOrTk4q7J32
RbeO7cEh4MHjIXRbW0Ikx5c+cKBz39vVEA89DehTMXAHDjTTo4wyKa6u9XTUN81t
9JbZ2eEoLYjJgbfUoyaNkzcv2qhSurEdAhFfchyX+pLom0CYtfGDpGHn2Iqw7CA5
Hcelqwky+l/zv98FX4HnbEIsCF3/0Tr4Xr8b7PbGt7zHRORrxxgl5HdajXFLMvCI
H9QE+HSktNPSzvqGPtMRkk1hhuicJtX8dMIXe6gVasbE8JhtS6ZPsxXxenmlh7L9
nmxBuMrrm9EXYcRBfVron/5iDw4DVBnsyVGIcH0ed6ovWF4GCOpL4Qxjn4x8lF8n
PCu/0psy9oG+i8txpaY2/TtkRFAy5NtUg6EZil4t4x0bZbJ1gztZqFg+2DWqv9FP
ovavFhQfTsF/7jyHgCNjvteb5Uq4YruaQXwjAzYQoZAbgsfEwpgbu+aFm6apMBri
YnFiYzmVFVtIUrFm64+u1fi/sOkTk6lfjw1zbbjGsbEtVf6+RKSRnuSUq/ZUFINZ
Z/WVreeOqCofmEUE+1G17jKA1ei/WuGU46GCnK0uHlrv1DaJfxMIz6sLYExAK86j
YlsqRvNfXJhqFwa7bqRWjFipvrA0qmaq7GAUdKbZJf/JP5AeVFVoKEUT9luKGT2E
QypU+Tulp45cIB4TUddVdjlYji2s54v1qpZLNIbxJ7EyEouqup/ocf7PgjvUKhFp
sp4HTfWQeOjsSacsDJBUtWjolOO50TQKVO2NRBqUKhxWHEOvc/oOWAe9oL81tsH+
ccPBJzNUlVodVBrupxcoCIt6fLA9SFnaCcGAUmZb7Gwp2TDzsO9lGw23iSlhX0L9
JeE35YwKKo+6dw11xMRmtl16WaL6sxkucrw24HYfDw5ZhHYpaSP+TOGJtY+onbCF
z2TZNSNX36Amg0FdRRP/hyf8jlD/70ErQuh31Albe4qVJqTcichfjV9TeXWzztpv
yXR+t2xGj0rDpeO+fUB6a4JlEw+3sIMS/+/Vvifh9s7wJKt9HzZrOc3WfZjs61ts
ZNLHnmvQUspGkWwlbfGxw6xOGXEaWTBVwtF0LvNFjueQACK9xt+saCQRVmlL1Y71
jmV7xiQCYr07uoiywKO7LwQ6H77PqPsrooLgJi0CGV6X0v4qqk4P6TnqVPFQrJ1n
2/iRwhuh215zEdSCdyjJbx2BycZSV+3i0tOwwBnbr+xWXczmF7vixUcMzSRpoixy
PBs33Bt6q77vS5SsboAciuOMih46wdw/fyOJAKBoBF8qEjaI4bfwT4Hnnt1Unb1o
S+EwhwDjcS3Zqnd7WwvvGM9bQFw3ZFhH/pdqTDjhzRq7ti6pV+rHcekhSt/QZJFZ
85zzYAKyQxPe0+RQ5WlALU708VwbKEMvBox+Amo49kejdx5wK9S1l7R2mJoS7YPt
WvhWz9AJrArbsbjgf9XsP0ap7qDo+Dmiw0xBqGg8HK9ZEipXeFvrYRkkgs0b3YD+
RV6QZdw64RQYwYE4p8UtAjEzzSKZ+PgKKhjX3T2kvXsZgqwU3qo3RoABxOdHhBG5
fSLapOPf/8nlylBBowcHPkl+TBQPXJHqWzW2Z54eMJeNSkzeORKzHMNt7iyqHCGq
CH7WvxpjSk/ImcTaWGkAM6/gC5REEycLFQhzYcbcQCDG3MX590uRQfipENdVwjC7
45naXVBTlLvRcnwU/D4hYjrQOhn6/3HEkZ4/cXPkSZNMnoos2koeynyB3WxOjCg3
4XiWnf1DJA+AFGNlpcwodv42veejplr86fJZ4yWwTr7dfl96trlIzhlX1126n4WV
LbYMWym8l4+I+xuNgsZt3Zts7WbqP1w2nviyTSkJe61H98Wv/5QiiQHCXs55PMtz
eqwD6q81j9jQdvJuWhW/Rr2keTZPE15qWd0GPLuWy9e69mFhqBN21F3KgIw3rYjg
LifgTc6UwEyxO3z9c+9ndh2Ngxf7tVIxAmzBmNnf7vxEavQ6SgpKcq+Flpm7/NaS
2uxysi8ElofYdG2LvqQebu6xDdc20xoRXlnxbsej3u0Iw1ZPBuxH1jJE9AI3XfK6
AWYnVm6iLX11IKiVweCOYhgBXHh+zpjYIXkHKKMCTnlgVy1ID/bYNlYzkMSUSpUy
Xo31ntKEPYSB5WXJD4vyP2pUG/K5mSvfDTV8k5FqhyMVck2s9flaf1wX1hKrIcwa
N6JDgaFKKI0cqa7pbs2cQtfzqOC+EPgZKbxmc6JPBKpHHsS3KPFbdbm4ph3ia1IA
HEJHo2Om0cyUtEayWbb7l8P/7/yS5Jk3flsyo9UdOXYNeB2KvFPwp9flB7oUs2In
vv4mpe26n0Nu3qnKAdKEVJUx/U7qPyQeiWqGJRsr+Xr5IFkJtxWva2MqiPWY0f+j
+hXkyct219dhcUjKB8zcZ9mpI/+9vLAY8v+FIwx64zTJFIAtYfjVfWnR9ip8Q6oc
L9J9HPSwx/4Vj2l3P2KOtlLoKgbrEh7xOEC0sFZXbqtKBNyz/YEJanX1WzAC3h6a
UIK62/Ey53t82YmwhyNvXLwl3LohWpWrU5ncu9mXB67WiOjavdOnrw3SD95iZnxO
6DwGn/Sz1lhEhXszwN7lX3mLQtI7gnusgViizwe/Bm3nMHSPm6exbwJoxOg73MSB
wAGC6NKvdZOjiH7+SdidC988nbTPKLHvMNey+kN0qxDNbLEdRy8zENWNj45SlEZZ
qnXrGLuj5MsisdzzP6LPBHZB5TLJqy0u4UFU31wV9K16BEqw6GDQqyOibFq0+XUa
spR5yjVv/F8UB+GJ7oVjBcwIe+ZQyAsAzABR7UhrvTh/KYL49v/kr4qkmyW590OS
HWpjqTeUFiPyJ8+GqzHngvpgAKbwUQJlDnL3yhBEPp2rAOQKWGdnQV3laAbDTzx8
rtO40JYYGioVNu8GcsaDys/rJfuuPmA7YHNRdZGIoQCDUywuNMXVqYsSi+1e+Dbd
I1NbIfCfWSN6jy9MeUWj0kZmYC7wKiyrRdqH5Juh+Pyq30QMB0eKaleM5a0CRmXw
OAbiuXXdxgBNip7gZQ1WltefATn6C+HcFWORUnBYy9EMITGHoe4d6n3DaLPTYnaE
H2lNypqQHVBsCjS0xMuRLEs9UJT3aayHVOIxtm0MIgFjK9Shu6CwSDSMDpEQAap0
08Dz6NQ+/3AMvzEqlz/0qU8LOAGOjguzEmHHqpkUp8gMirNOt5kn8J5d2mR8dxXn
v8kAIpUu7Q/Dp3kmeIHhilhu/pdOjcsXsuzL32kex7RcLi6tSzXJHZidCUYEWXim
eoigK1++P1q2+u0+XQFxBE6tdZVjg3ZqqQXCquDqPbagYt1ZfTrwVH/QOf0W4ZkZ
bShQy1gEhVZ5TOSgWt/MHI9TZLMuEaQmBwJC7M53s00U2/GWfrX2aDSVLzoRg7Zm
ZYFzZ75caKln6L24FGgeEMcVuYIw6rqJNl2oqMKPcoI66k/FzpI75lNFEXzTc7Rs
ijXW7i3l42QXD2gxt9wILfG0rXjdrzETOfBRvXANQGlEcqZX84A3KZv7jPdL4S4N
1AVczYgE13rcvyyAuj7kusDalEdfRaQxd7zMkeZNbjGY8EaLQ6/kyWH7IK1LDo4W
3iD7Er8oJ7qAYAg0gULMzAJXBqPFxsILoYpcbAUacyGB58Km7cY+XUHHJ/KcqOQc
A8keRIvBSD5G4PPTQWM92+AaNqZ5yDjZ4EC92irJZLZOq/gxKN31/CIWoeWLyBcf
zCeGRa7wLOL8G7iz7XiP+3xYQONz3dBFMZzNh2TA1lvulJwNN6WhuD+bJNicp+uG
zLgOz69uqYjG6kROqUWCIGQtnw6yyTX/U7mfZGOsu/WX/CsEJLP5VwydymeB6r7s
QVruftVPuJFl68r8joz/hN9QWJeej3Z/hVGjMmdllD6JtbCAi3CcwPamXQehNelx
350H6VJACo/+HgsbMgYAU55uosZ29ZJlYPBRBalBJlpoTm9cTmjzSTYaQWGVMLhr
WV9XPAYkSQ1BTyRGUME+oo9spr5pX9+YGv5SyAkLKxpRvB8lbbZoXNFWLmJAORMi
WJp0TbTJKYRD46/zlatdnRz+jtypiOU9aU6a9sJQgY+WufLMwT7RPFgC/0gohtE9
st6bgfPlj8wuY847AxZg2r/11o1cT2Yz48pa/LO9znbRzn3uPq+YDZekjwnmCYsy
WIZEahKlWAO5cUeefhRLGdlSEU3mjtgmpRZfWIffjrGkOZ7L7JOxKAhi3cq/nDyd
idqOBi2jPh6NLCqvyMrCHq0pyH8t4GFMlg/ao3cLt7YZ+F4YsJevQ3mU0yMgE1gR
SctTc7Xmpt+Gtrh/lhjrAWXVxRSL3mw1gQkj8xBhMamfq68wvjZWKE0GZkd4kHtL
8LqbK6vygzVsfm+soR9lAd7V4arIoIs2nJlddaZyBPOBnbF00LoGGtlkTC7LcvWO
NJyyt5jeoq2OxVJMHHMsD6wztSffXxAO462HV/Bstr0XUtCVrcqxf32gRAE5E9f2
Na9VGF3SSssv9z8CzN7p8TrQ3eyzfmpchBH9yK9TqDF599D7JsRdHwauKqJyJsIG
9Yh+z5mDHN15S2Je1YtIW4z3S45lmpHrwlyB3vIr2HvdYJ8I4qePar7gvVdrwEor
OggUybbHVsZLeeDcER9YjHsITmLymmuYi5CTwUoMz1d0HwJLlUFWrjUI3Dbkqiqd
R0DTviZ1Zhbc4m0vaDbyHRpsdUSujXJ9W2sO3dZ0E6fNEc7zISrG3XjXKWvQY31B
J41JNAZwOqhDItkORE5+Fx/FamN06IPZK6K5F6wlxW79wj40gRAtbE8S1nubnz9L
UixyX2zZoeeWNfOQhe6JkxfV0dyluvMpSgLXGE3wSJdl38Nu+l8ig4Mk5J3Wx3rO
QcMafHQzVIaVdFt6XGnqaW+3lI+l1DENIYXu2RxCZ1QBn1zn5k8HozVmwWgDxkya
NtHLB5acwmrPw0Jg9jLBtRiRBe/dEi3CBMSx7XMMtcuUQpJ4+05NtF3frKFIoOW4
S42RWUhJWdxvQNjppCVYMHNFMtZA7vAVm1Tk3/kDrfEsY3XZl8538IsKa3O5vzT7
JrDa1mcHGdGIRt6vZcUwXrxkdzlE7XYHaoRQUNTqi9jzUzay1HorxO3XeR1dkIm6
7zfwbaonEIgaVG2bUftFbHn9uwW8afUa8y3jc91WpiOin88FfGwPxA6jjHJ3XGQb
bI/6iwB4AjdW0VwFN247FlzljXQoQ7wB53WeJIZ+N42VDaTACZZvon13a8e6+0Rt
SlnupRMJLI2XegHCUrQyVItgaMJq0kTf+W5IT31YK/C1uw5K5Oqh8aoGTlpZVlXB
BmwdoPTSLquDBC2FmRmc+UnNp376ACTW3vzRoGM0gtMqcQLuoH+AKh1CJOMN3OQI
c4bIULxpoSW/JpDQc1AJ4Vy3cXn9F/0riYLAgr5mLT+3zX1/3TzqAUBv9Tmzyn+1
p71wYY0jk4NaB6BpPSxLKfT4dzYkSehjBSKWt29LECcuGzV/rVhpS2+3ZsHil+z/
OsE5v4Kgspco0rtl311CWM3SGsmOM0fMCS9jmzhnnNiB/JMF1iL7/GHM2aj/So7T
cO/gdKHHiJXcRI5NC/aORGj8rBwiSZHQU1w9nBqFA0AVo4buDWFhIlxLxPOYQ4sc
sr/AwzfnjfS5KWYiH5THNSN7X98YYWrmGhnDR8uJdB07G88eqhnefDpBPKwLzApt
3CrqZoVPeaX1RiqOY441jibkkgCVoEtZeldbXs3pvEsG84C8z7oxrhQpT3MINpYn
tm0OgWZ8HZJRG4eNMplHJzPjrmUqeaES4NYWujEUNEVxgck+4sBnboBcPtBYj9cp
GGgsKgJu7AXJSd7mPOrL+5LrWk392l8cM+4+19Xn2oOcEFhKWAllWrYVZI2xpPOm
UU+UBVa6pKKx/eLFOeFNKl74gsdFCPV9J8buA92uIXUiK8Rnb6dU9nAEvAV71r/h
23qWaackSXFoJxAUB/Y0awuyr8/qOVVJHZ6CeaPf3GjqgehQjzTo1C0mrereuMzj
uoha3UJTceNq8JT94BLP5+9U4W+Ip2mjrZkD1GtCvWowuh+gl9LpRbxW12L2hvzL
digS3/xKRTELyrXYPv5Q0uWCcZ70tNdkk3eFQT+7ft/ibL4dXv9C1g2QZ7umZRv+
JW08gjwV3sWrBU1VWI6+Jz7c1Oilh+FJfTPAvQgvU4EJ9WVePgI9G3DKbUUMfqvc
ZlsCCI48qekCsj58mY9rbyC4Z/aXcr5K0Xxik6bLsfoHkLSHuL2yd0EwZSNrNRkW
TbSsU6j5gglRGr7GtkM9+/z8oOthWvVlVonp+X+a0y0g+r6V6ndtZZagkQM2XAyT
UO7ibSESROMR53E/y/IdcG4cLhP8z/q9cnN94Wpomgnk+cCbVBfXfZzp7lZwXmRA
s/nJKdtxTSgbA2EzXgDoZ3HsLbxlg6tv2Jbl3X8eIJm3OJrBEOkqEzjRBXn4cRnE
AsG6qEGRQ34NiAL1/4jNhiyCh+wv1FUbcCrZxAU75gRUnnXzBkk3fzuhPVjxp53u
JLjqtnVGaq6fmcAjfouQh0/BLaOc0K88k2fC16U0qztskzzZDDgG1/VPwXwrjQhF
U7bgSJ1LvCgk3gDjH02PLSf+lMG2LJn8SS6JQ8WY49WLxQ0lj6MbtKRuwEJ/RUI8
NZ00A0OOtaHlD7x3pq71QZmLmBODpd1F/rmXPHHJ5ZcQ9r9JEjfWQwISYKYxb6u6
nGz3z89VLY+mopeOy5CTQS7/K0EtBBP85sJfGfQUQMiI0qiCrD/0RIrklg4/x0+f
U787BJPVPqKtn66E2wRfY2uOFwJJ7FmmCumuIgN6SRkvx80lvtDMgMyarJ7paO6g
fVdS1f54kPcGpC301O0v+e1AfJXFDX2nUkAGAqOcF83GNSEtpBHtbVPPgskdBkV5
lMmaeGQPE/BUgKccMeUP/vNG5gVrC+uP1xU7w+N81vwIznS2HhwqKJXnws5gsG43
TCpfsSz9rkBq1d4aUR1M+bUqAfhtP1EGaY9QSRemqeNx+tDcL6sZFjij+M5uXPWk
1tA+F+gkGFRFQGgApLogi7M4CtlQ0iKDaTu3l+N1+0Ju5XU+gdVKhGFagYLUVByi
O6/m2BH1WD2PKiNGtFfjedNRxjBhviKvHu+6kC/jsJy/FipS7nWbVJreRO2Vmo25
CY9oNwrEWQMWu1L8sCihmNRYfbCm9/O9nW2EkHSvS+7OqDzEgaBTVWDQR1XERDr9
GkgKjmje5JpNPynZFyCCGmkuY9P9tJ5ltRMM0Wysqq7Xli1EcCCVz8H86dNOZVAF
iSJMOZEVW0Pfth0iWnsjYnV2bOEKdQBMUT017b37tt99kP30tv89KRh/UGvEXGyL
3HLU1Qh+DMF2xazmrSd9jowePYThXfE47wXhZmFUrqaVPjSwx/nLsd7nEGyoaELI
KmSepm6SAWC8AK09Heac8VgQf5Q/+4qntU2imjMfn1OuPBxTkPl24TQViY1EES5Q
k6VkEptmgnCy1XkbHPXlSxEmc7eDrbdz19Hp4ayKW0qjEGTZGXFmnQPiIsb6CU5k
vvB3OuoHt9SqShnC3i0MOsfiVly7ugopfjLUfF98Fc5VQ3TERyoxW6quyUIcgBt1
I4uuGvoHQRsJ8KEK3BGU/rqAdHSnEYM6lMWu7REEu63mGkPmgcg6oPHRMuHDYTQu
+rCkwookKcXpTmX+gRs9BpuXnoj5W6TUdJ6Fza6qgCdqsMx01DcUK1cuEB0iiap9
F4D0XGiLvFJSI4v0yft5aqswaazJ2VA/HY3ixNIfnF8eCyxCXQC1T7O0ONbe/h/5
0L4egLmb4V76TM8mzZ/HdS8rbIMoemsR+IOtS82f2Mdw5CtrDh9ozdangVJpoZoy
16TXsdInubxPfeiUPORV0m921D2qU/YXxTWn34Oc3OZT1cfSrD9KdgzlDCHphhyn
5YaN/Wt/PfgEl93LRpwqZ098CJHO4w8eCMNKLBRE41Gas11QrhXABhFDdYQNOb29
I2rn5RwMdcuFHXOAaha3wvg1S+3KRPNc7CpZSIQy+55QCNlIZaBfmzs9VZL06FGK
F4/d/kxPK1TUQ0CAZOWLj3dHf03TddzqDiCue3ciBr6FyXHjYWskt4ZH67G4Q7zd
740998yDaop+GS6hj4qLddL3cP1XIABoEC1tlK9h9IHyqlN1kaUfBwKSnp1TepTE
0JAp0gG+B/qRYOonblC9KnsC/fXMtsnGfqwiktQ5kbOv3DfbyxpmHKbPzSa1XStL
WVMifuCqWjrSmWTkyvaUgNaIgEXBn+fI3uWSlCXfgwJ48j5E+SLSPFAodtemyvKh
dm5XwC2pcrDsEySOmC6FjlWXeI6i7AVDxeBRHysaIf+b0E5Az2vLYaHzpF4KakjW
ITEbubRO5g1AvFkz6xorUq0QpdJ8r7VJQr+jldb4d9XWSnO25rGs9haOxx7TewQ4
+wviRbh2J5vDpUc4zlaxb/JgZazi8Z5f6G6AM8YMZI9oJW0vFq84lsiKvbkzjxuZ
1/HQf4IXdYIOkT0di2lDmP/U0F6VswpVsDyOmWXqxugYkS44PR/w6d8P1rYDASh1
G0Slr9NZjq64UzTWqdemfVICXrOdrXCJw2r53hnv12tqO6xbfJfgomjhqWEykuUp
nN81T9g5S9uiBa4WUcppBAGbLvbZChdZaqKY7YbDp5rmryu4RoPU0zrt4tL0xCCI
u0Qf7VOeF2Jf3f/gQMVn46q4UgWisIImd+B9r6H67WuRyYyoZ8pN9c5c/j0tKH5D
qmtxxeM+BoARJdQ35uDAp54sy7f0OszvGuesl9UFL50XK7RtEZ11WBWr/A2VoWys
sn6Ox9CGj+uBOv6/OC3hQTSiNT5jb8fd5fgkAm3J/NBknyZRjLE6kppcQzrqq53a
FA/e8BP+qo4G8OjpFySwmpA8FHu5dHjgzQHF95WOtYcJVU1cRzJZujXIlzGGt8rP
0zjkf62CXzgbCjNW3ijTiCDRbyrF7b9yMOF+EPKkUtPVx77K/Iie1VdsmTtclrgk
R8t3Nm1Hqs/lsaQMcdnIQ7orLuefuiHPbQaLmdlk4CCVb6Xl2oQcoBFu+t7ruQQ1
QNjgc1jsSUHs4EoBoKkoRguXb9+6rSTORpqKQO33ZjNXYF7qnq5z8IKJFEYeeMyh
euR/lQBrhpnqvYIuR05RMaQaW1shIL/e2qcyAEZ+ZL7iv5oFtGF89jEmwHi9a32i
jJk6VWD45snSQEzbnNEOie0krVXAGHN85PNrI8TMQASYQaDnZFqkhD7d8gBsVwR4
vaw3aQ3uszJAAFHr4ZTD/uiNWgErrD/08PNd4W108ah4UTCBHV3LNiklsyfF/xgc
jayKzpcMsHSJp5nxDne6Z7uGJCBO0oHT1ZqZ9DkbbLfa+lazjBti2RcQFDLYmeVD
F/hoeCwLt1GUHI0H5m1VoNxUwma8EOsXMb7H4ZjZVOLSpRKwuexc73fsnime2H0Y
JHrz03dF3u4bkpRT2ui9grO9OoKZSmIo4weFk80R9xuKO/ltc/I67fbb3hO/gYYC
mYAnNzewGRk1hKIKBVSjnrn3genn5G1GlueioV2VwrgY+GB/ryboaSOkAHvqDbee
x0n8WCL94w/71eHLTfEmQ6hDXjlwwwV14KvFXDEod6dm94Vh7rEfvz/F/CRXBxOG
8uXXCEx3Hk1TiHXdBbjUbTWq/OmXMlzetO6bLdn2fDgwfP4WMvyobqV58w/qaPFO
A3Y2OUCe5tOq73Jz9S0paqVZmGj0IbwbSUjuh6YPhY9m0hoP1zLO6mzz4HZM33Or
yKVVg5BmYNLSKMJh5A6x2CErcEdtVm4tYbIjcMe7g6Qq7nnnBUhbnuCMMRQZbvP7
hlkWgMadUkTn/6+JXleZHVALi9+4FGHC7ACKK7l6O/RdwFBuwZ6vN7HHxDP82vIA
SHTCsUBZOjE9lLOpq+zUfQSYKpnKZiuNrMx27yB+Q6zNu5iVTSi0DJ64XaHHQyeb
113+m7S/tacwlz2cs3fcCQB3WdvbskgK30WYNl35Dpk2r6TCcTe8bu4Mr1TL/RcS
lgDRmXXEc+P5s/BvB23cFNW5Ijn228bGwZXOn4VRj2YTwoN6cvkaFKZPCMD3uPP4
Lv4ROiyP4Tl5a6+48zrclEDqwIjaE5FPJBobIGRMcZNVsekN/7UIkpK3HHS62vZy
9QziKfr2ZjteBUN6r6ucx7JAxtg0pOiX0lPsNTnNgXQrfNQc71ymWndg9n2L6C5N
8QwMzrZIsOybQ/N0CXUtkNWiCc8EzHdjZoBat46pFp7A2uV+geRDF4XD7+ywO7ER
bhVLNh0nkoi/lqGNKQudYE5P3cimglGIJeev1ILAXO+GiqgV5s602G5jI3h1lJnS
CViaf9YqBIGrUjKcCEY6o5KwwcMOGNja6rPrpm5s5VwyCFNWh4Kdy+qtd/WZvK12
Bb3Pn4pbNnKELwfayh6nhmcki0lUntRgUvoTwjuGtLgX2EpcdhZv+d1CR0ulVgwn
D5rZIbCltaFB/WZxQwGOVasYQR4f2W/HtoF6lT877xEXrlmAW4FX2vLq4PqAQAh3
DWWorzhUmH2llwnSMMmmRd2YaNAFjVC5LlzdfBYvqKdfFfmNLPYFc0mvXhATdOQB
gM5+x8VNzOXGQOigLTGvr6Oj/Gh6fXL5wbOTc6+aB8oqFVihV/CcFqTqw+Hv2Zvh
pofoHFkNYlXurjr+IXBK0SEWF3JomdmjgVqihiIkVHzvIP0r/XhUZ2HAzn9NFdCq
HrsWnqq8LFqzrqWZAIU5TeSv7ZRpnShDxot+jsVF+6kgtFv87FPNIitACe3oZxLv
ArsSU88+/1MD3dGN2jQcw8bGKU83YjQWQPH+2yLboQFmPKmpgda+yE/eZVSUHzGG
mReXEZRjVoy8ob21T27N8OVwd/Oo40oocLDlzpbfXEOtsZoZm/aybDS4FPvDZcLu
wkGjI0NV+ghfkFEXS7a/LSdfseAvfnPVKIhsJeRGrroLme+kLO/ysk5n+JILPz25
F4o/SGwT3wf2S/n+9r5mER97NXNtEXhjhuqWu3/W515RxlPLH9X3bG6Sq7zMh1aU
EmKLM6ozB8IWFdIlE9Dx8uQz4nu9s0MblUrbCpTvBUWjVi8rPcC1od899N9/UaZO
9a3Yy/0qCxGEFMY1Wtl/YdINXSSacyiMhy4N/H9F6xqA5rh0ljGC/fX5ulA9LMJW
UrA0oG95Aoi9e9C+mxh9Bd7HEkRcc5TFBhhiHxK6Y2/7IA3bpWEp0yFa8eYyJQsb
v9axvaZXiFd8zW2ohY6Q6xOeQyApC6EmrIorlSUzgpEJ6diQu+ET+IqHazFtDQ1X
U+PbSU4aonsM1I/j14Djv+JmIwjNlY4WFabZbA0SOTJdcjK58rFa0xkyDRaX3g0N
UFT7ARnWfP236TQH7rTDIRpa0z7+l5gXX/PPzlijTJ51UawZJfm6gZLDmM8Rq40j
sGPw5HgIIk7BFosaTzNmeE8erne7ptNbiv3BBA5L6Gxz+cOE/jYU3AaJoAL5MN0y
oNste4K3kasnbYGO48qwn9NcFXaDYIWSGaWUutTXmAADmRK/TCfa2S88RFupDaQ/
cjyTZOQH6m9QFDH27tFTnuZp7i9HTZOA6LXkQ3XlsqSQpzG+Nx9zppLDA0g9htq+
g3xbnSer23op9kD65Qb+dSL8Zn4TtOjNl+Hfl9GVB7W8RJOdcHVNEpWugZkqkfm2
2jfo8E5CD/zcyuCdm3HzkzqT3trK/tpOzid8/R6cHJ4wVH3BYifo3k9SFvWUUz9i
vRTOhFYpV4l85ae7rJ8HbEneDm8r13HEBkWw/JuNaD5WYkOFmNX1UvWtX+cATiwm
e6eaeimRdhcQBnsFdlR9phNcl2fI9f54XajqlBNPXUTBVBLil7Yp87Ubo9Xkq+C1
Nx0j1ozhefqWCgBXN3xz6UOtF8P/GJSaQ373HEvzdrqOHD9Eiy33Uh8zoLQ+Oddo
dYoY2XbQAQ1CODaalgJu8lVzHqcEklwUFlkrDS44+Ru1SwBDqxGzDRf3eEo4f2/T
+PfvvRxDYwJlDcJoucAVOT2mLuNF9eQGe2nXZDb5RCQuw7RO9sLgteGWWUfJHwK1
qYRaWaZ/gDLAHOsJPy7b9x2lmblfsvpQ1XJKqGYmDPdhr1in8h3NLtNhE6aHYLx3
sRIwrtVaRRKmFojjy81hO+OhjW207n9K33s2+82GB2BUeJiIWyqJm7Mwvq9akv11
sWZZuLmsMD9Mfh6gvONrMip7wfsJqVNm2L8bLjPw7Dkaj2VHVaqDQTIzN7XxHVjm
lgdKpSR+t82yRKNngJPPV0wqAhbA3C2uVDjr4t5ZRkIYGY9/UklAnLKdZoKCtrCz
k5T0CjKEmBU8h4ofhVUrjddWa3D/k0zOycdi+CJWglMotxX6V1LtGJy+vaeloGF4
G63bFSx8LgMg2wb54on8BhTC7D3tWcPX5Js9yEX3NoNGO+Ltnv+o63eCzMBl0fxK
PPOV+WBNVvfohJff3EGB3QDYPaYce2znCIoxPdrS2LKYlNiOvJCsuhMxfshh/SfS
DrFwTkJ4nuiNeg7WeIN0D0ttci8xXtmRJ8b2RGBuB9H8652DB7OcfJGeRncme9+b
1Le3cgFswPXMvOHUskUezmgiYbENLdwZDWfzF3tYbfkymclBCdRwPFHoCUmrqep0
5GKQVSu5yheUbg3i/dlliGcr2mcSk7REmjxVEKA4/pmETY43p0mzkcn1NWbBdJfH
nj32oJ6Ul6r/+Rp867TQRlHwF+bpzz2JVk9lOBpjWZUMe+Sme4rhZI8ix/cs3CiD
YIfOuKXPiAFq4GsKKFeumTTs3AWPlQVlJcoYMaDE4NqPrhmNi4TG23xTYjfUx5u7
MLlYe9lxeRLDY2TFxdn42L9Aop6W5tIbkZ1f7vfD7Hw7cAnNoFOqUoj2vLBuHbkB
J8l8kEkkoYJwoF1txwN/hoNhMDcSJU4IFmDhB+9R7UQFCf689o2onddE6C02zqRF
MqNVyWIHaG2/Fit5RxbqtmPRd7MbYWZjGBTg0/nbiqS0vvZ/uzngc0D16l8GNv33
KGacFJquvt2+lXDofrS8bFikiePNI9brtxnK40FzK7hjsxrpO4enASbC6jyplXZw
LJrW96u6XjTOVDzgRhRm18bDP7iPxiMeLXbYO415BtOlYqFVbj916W+S8ehN+IoI
QDo4bUkwemHfkd7zjwI1ekjzbhiBv7WMPd/3DZQDEDP1Z0RNBJtzTgnmoskzRsW2
Np6WJKrlmIJotUt6/Eq+HhqIZqM96MZVnsvLOpsxnKcu32eEz2LqjH6nAUxA35t7
twSQTx1ssLpdcyUxaPU3dDZ30s3EdbW39pQ9lnyyRejN4hBzihwR1W+G0vwg+UXh
AMkzdehflqkXdBNwSt1BghAS36tFWjL0amB2uLeo49DCAz3/Z6xJyax3r1H86ZoH
belxg9hKAOJEohOnateSuvF4g2BxT3h3SsOOWIaA8tsJ714XB3kGl+RPicTVHz7A
+4lhrpyJHx0FvutgOt9eLfiDXr4jKoV1WA2ZRSOcW47JqDVP088unlKp2bAu1c/q
l0cYfCMRmjB9yanstHIWyZLUe2E6fU+T+jcyAhBOb4MsUfm65xbErv4BWokMsGFR
7revuNrArFELhLD83JVSK9D8RwhXaLW2zbZKHTV0Zz+Y1Nn+bTIbCCfyLTomj3AP
44gMGZHXPTVEDrysKKiUz+S3wRmUHlJqf0gCzY6p9bNx8WWOnUH33CM5lFMfaxl2
BGs/omVrfZOqkP1xNKfk7Ftz5RqBftX3vtGWm5TbULQOrLD8l/wuCofTPYJ3e0BB
fugk846Q5nORgYuYxZo1S8p8pwePkTvdHFVIzy+zqcG8uSop6xfnNLZZMfvyE29J
0EXQOputwKuV/44fEbDaHXP+XfardnA4zTB/JL862OfbMQGkpzfgJHiKUwC+uaHe
Lk7DpKQQjwD74Ze9KaovVINucv2U20gBVb5eYT0h+k44415PoGAVdlH70/k1f/ZU
p5jUnQyvlYR7n1MiS873jaoBPzEm4LfNQVRtGvMYYtTZSdXMofKCB4fjGr/PRW1M
Lu0QYZVy45bsuhCNnz2mOBb3inJTcTBjmcsm5eWmn6tX1cn2Az1uryzS8gq6RIrK
ksrmLdPgUq84SMs3Xre6ab7SgpTtUqrYo0Lda7pMhHor8u6nOGmkiVwTramTmD9X
6Meme+3+jlLVUsH/oRDbQzBst/d2MYD/YGj2yHLvkWd/bfDImXSQeBrizFiFohwS
hwbEuLW4JcRXRo19WHbHrvMJD+gFlZ1icsi4Pl+cEOxIuIT8hX9z12b6KvSRF8Zl
+AQa5H6O3yCZ8sQp98Sxg0d+ztyrcGGs/k9B8kgnB/J0atS9AfUPPGYvzfKwo/pC
zWYFFho3iPhS0ltvPL/E2a9JntIRfgT5c2Q2egH1jQWzGrQKLXUWINlS45TPLJ9+
+a4OlJmqrxzy23Wvle/pgK6dZD5kjB3kxRUQZfLvsxQrp0cfxkIn8pW6c2ym2bhY
vV2o7Dic5++cckYoaw4N8RcR4EX/XY/LtsZ7tYbfsNTwBqKh/6ajvJvhjQqI8+gX
16njugXLLbYsxgiA2FG0Us+a6rCTBbiI5KzT0ZmzQO9YXwFDKQ49J5GlJoLHiPn9
ew9HL7NiBeFP3jXdtRkfK4cc+URrbkSpg8keGd2G+iuJkj7/KDIumcaCZZNSxZLs
HlCaWgZoakarJkFTsYGBJhMy0zTf8ErA3a8m7kaVB6DGH1/31BGhZKGrW2amn7zs
TkILpNY8ZiMz8PG4PKUnJ6XbHRJaqhDcXqF87yZ3Qcqg7wSlqtq46dSc376IJBVr
RkoP2Ftobo157S5t1IXeC1vkZw+HHh9HASvCqmdd+po/AruSkzLICMnujgbYsXv7
r3VQFqsuqW5UI0tVT3W6yIFkzo6uCgOtiy3xIdrWcQCQ9oHkt+4IFR3BpcZuxx6D
oYzIgg+0JvmEyGqMuGECFdze6+V4AvaxPNTwypNNWpKqYBOckCs2qCNqx0DdsaFT
tiSmLboBP/FQjpKbU1JK3KYh6DVosoaEdOtCB4USQt3GSaaByWro6J+ejZzrNyNG
JfvDwA+segrhWZ66eteJ41FWA8vroNwwxlmoGtv0x1YOqDfvZVqm64QSpCr7pM03
qXBzj30WHuJ1i29LfR83V2AqpMN3SsHJ/WMwDyv1IRMZWakZduYqPBUlKmoHzSuF
w7gVgbxhykYx+8HYA54FjjEzBhdNQixqnIaz8V31P0JOf+YJxdAfVTpaZqNwrGlS
26xx5qnKN7rehw0pxU4km7z1E3JSpud2coq7Iw9FZrHQj+GOF6yS1ebwInC7ELuE
2jTrAFc5NrwsiNvv5h7h3pv1QqfLJ+486HfKik7evTdPuH0KqSlOZFD4+fX3IjTq
gX0KVH7FUsC2lAUa+DxHVnYP0Xkju+Uaei2woSvZsGG2LvjOk7yHflHjiKsOJFk5
yCBJqTdweWV8RVfaptryePsBe9gmgbQHDPrFVo9OZa3MeDY3/viL+Y5ipsz6nMY3
exHEGNJa9Okfnz5pupIbcDw0LxRI8KjQhUXlAYqaBImUSkEjkCrbCwu6l2Ov+Uqj
KMlOtnPA04RnJF0vqIqKa+ooINeQfEAFIWrBCVm+3qLhzuhpaZdtje3n9LK1fOt3
/kkuL2UNYGb1F7iDhZ0fv9Bgg30qHG81r0X9ooXYIsKTRam+FMpe8YfoicIFQ5g2
Ib2t9m3VKMgEea3tHcCctL9MwrZsv2yDzMAeafIY1jHjwo1ISP60V0DJz6yZLYyz
qweEKEI+h/YS4nCjRUTiRfSg1kg2rAO2jrp03vZXG5cOwnRLLlVh4EFRYnOhEmO0
FZT2d4gCAp764YDHi8vJywc+iQ9KguhcDrqtEBRph6NlFORXQIBVL43vvw7Edn3/
Ag1cB7RQi0z34nDgrOsJF0ogRMalyba62FgrWHi/damjSObGo/Ra2LlmjOGwlgw/
0kHub5SLG0YS7q69eONQpSE56MgxJjzq4RMqgxhFDdEWjLzqp9uhwaY/670ZSYBZ
vQ37oU8VSgV5yWINcFA17eJGnsIvhjY/A526+JCgEjVfiRNpgyfekaGZW+wvp46F
EjyQzzMQdGQlSB1/F29ruPZvTcB7R0G57FrDIHXEejISFg6hHnuKrXkmLtGdtAIk
A9BhOPnxaqYyQTzpwZhvcV/gy+1dqzpK6WwnTXFSseDcNeMdXgKkHqO6c+htqYBX
75jap3QisIhT0sq3c2ajOWYTp8tKEhAMZt17A9I04u6i85FjX/EVvvKsz0UWdlut
mJHWq/1H25p2PqI3lf63FXb1DXJ7xKDPe/ZwNtPWl+3eQ3eTxsNoXttGbYsrySwh
BRU5tn/B/aXNGF5GJON6DqK1TEd8ALDv8o+ZQ8tGGUPtjEVg6HRck2Nem9DKReCd
32MvMPp5ue2QFctKDdKX70D0vKk6QvdCJYde791cRszyOlPtIdOCVfvElhkp9tnd
11cplEYSnQfTSAbYvQkpIZRUf6VGXj9rPWqR9GhVoeLfqh16n427cVPtaMRC5Txe
EDxVySPQwfuDuoRwIGfH68BfK/G3S8gBMteLS6u5uG3SuHNJ6rGwMwqNZNRSiZfH
S8ptgVk0/I2mF3YEAbTaXZv2Fb1YfggSv/qEgna688aLAROEtCR4CL1nI2uAhUK7
S0ZdZm8iB+vxNyjWDhVgUhdYP9zdXupmc5nF7zGL+7wJqkcFz4XgVqMIo008vfUa
/1RluAY0RJxh/Q1iGBWr382+Vv5hTNGEpDyASPzN3vcaG9EL8vxFnY8xpO1Ouw+5
mgBEW5Nkb0OJC1ZjLG89MZfjPBgOxQVGRAUT0FkaEzg3pnCRXiy91tzSUhb4+qXr
Nq0rgbBti55fHJyOJnIsda+te9Gg+ToE4Lo75AZ06wRr8pI7HaUnYB+3GaCQxDCg
k1TRCZseyx2q3oe0ApzLbWGGEfoimY3GLICedU1CG4YecLBzf0s9Jw11zoo7qcB0
u7kGJBv3Qhlq6w7baOUrLHTXaDsl4gLCSZFuAieeHttOEclHXNUcGXCvSpnkoNEH
sHPZw3fqoUIZeDVONQfR9wX5/kzUbS+bE98vBrfAbr7RX/ncPrvIdF+X9Vn3DW06
wPLEYAUFa0xGVrDMUlO5g9F+DZshqCqM93n1PKZKpPZoXHI8x4mtv9I2QCRsgRVT
nYyMjegRzmoITHtW2rio84y78IwF7/xMwiF/xL7WNesVZspvvZ0eALfEcI+Rlvvw
oGuX5vTnCDRmqk/Xox8kSBNNmSLEChS7J5dSimOzJXJ7GsbNPQB7TkD2ZbMZDXYD
ffFI4HVePYRUrhNSErnilY0PwX+z0Q6yeDzDQqz1xwiLa4b9dRNbfCQaczMWpsI4
G13P4M2k3HtKFr9+bjdfJcYUY8cWHvfc2/kDFudfDok3LDDqlJJzOGoBFfIO6gTs
cl0pmOp41RttFimF1a/+PuBhxCvHwT+Qw22leVOKmYBa9XvmMoFJoLyUMx403if+
fcNUyrPsUIDCjQkpw/psOW53rT3zALLO8P4IBQgds3MkQInZcamhuiM5V3aaYb44
Z8XhlmsDIe/3Zw0abSC4jfls4H1mZUYkc6AT/R36oF6/IqJVv5OZaOUcaqEinxUE
bBbcScmtea3kXUTZfiQjWHI4uColk0NwuOGB6iGO2by+QkCF28ZonQ4oGl1UypSZ
h8R3mBa+uCR583q3O33EfrkT5foKPQ6hMmjBYtn9RLtbV67vWfJ7053d+2ttjf1h
dW+ilj/B31A7wk632zXAPEzflm19X+TEiAj5zlBeWRtvmo69+RyFOA/SEIfOugv6
K9i8NYUiQi4ijuE7C7Cs9LAY6mu3JH4sI0IN5CzC2r/kfNW3wx99LpPi5DQoetA7
hnOo4EzErraA9UeELtN2lJ57cvyvajqi94lRJO6XcAXHQVH+zR/qCz3UTMnWxTMS
AAWO5MxdD7EB9GC0Bl2LjuuQ2rQgv8QNRnRbCBTBHaHz8221pNgHY7ut7M1qgcvO
ZyLWXs9eCD/eV8+qbTNKF+JQN4w4hwThp053pNmBISEhuh0oUR/7cJwBgMmZxCz/
MseNWAEzRc1qhIwRvtgKCr6i78gt5ip0K9urfukSZn5nvNB4zU9Omr0PoWDNcGTl
YcTjzb+lODhRMZiq93B1ZW2gXc5GgaNEoE88CXpcF9zgYStNht/Ko+ieyF6RzvdY
qsfANEiJfd1d9LVl8ssZ6YA16sozzpee8ekpLQqk9uzZtM2RRB2UtWxq9nL11Ehk
KBzPr2p0Rb9Ap1EQ8uJMIudfhrU+21qeuD1QK9dzKvrMAtQGbPeISeDY3Q9SO1u6
kWFa3Aadjcn8/3vme3UneFqhOfPiyoh/6eNq4m9EPs5XZ1IcUrx94chD3gGSknbv
eJVuLtmUKUOePDeKvvoRsBJjfnjYgBwkoEf/7U2jaXf6cmM/FKDYN+FsqvadWuEl
SQzzqyH9k2RRa7IzPp8V4kgX0FDoeO0xtUsakkSrKx5z81kedgk5HG4tVG3E1QYR
MsQihObzujpzcUdasw0Eec1PPwOmPu3QcLWq8KJG0uiHdGBGSzAKRkwcOP35W4KU
gfcFgv7iBRaf0nM0Y4fclz3zTA5OOxiuyopGGjbuVmWDRouAIVPwGt8DflhMHUw5
/qXe3oA9qE6Owgx85dieNexKaUduIpKcs2OQsyJFN81mBQamygMN+3xC4m/GTelm
C+qeUMpH10EiDiJnmu0mdIXbDk2d3MuylBYRT5zuFlcXRlBWHeVRkMh80w7VbVmB
ekrYyScjWQ7u1QD1MxMXnvsMqKIZ75auxRSEjnwDEyluFvE3Ku0i5FZCI+fj56U/
jmnvXz/AX+oLYLMimyqe4VZ1SYjZAK8oGaXYbxIYdrzaz0KvdtlcYRVgCw5/qI01
SUyC7n/Q5ZFS1HHjj/y1Wig2xQ3vOoXijTxb4RYX7HfA9lqKlv84q2bGg/apwBPK
r9rllbj9rIygktmECAqSigCdbIlDFaDORJiocZTY9NJg6cCNhHN93pD5wCFZsQ7u
SAIKRVTragstjiCWjgLaZdjKwOHOw87YQpilD2hwwm2vIsRbuFlaaR/xYSqcu1pr
hIiS3IzZQwRdPr7gzk2Ocuz0EcmFogjK9O34A5xwEMg8O7MDhdNOgWARMzt8pSAh
G+79yEGo4SV3VtZQuHyYXfvL5Ap20dS4KmPKc4VkYeKY8talUiwCCNTSWzaGDuf3
dik4CkE0RgtBYK/3RD0SvNuulg+HGECMQBDBto6S9sOd2PxxjAPx5sSnHCyjpdCj
MqdZuC+Uf6CqoqmVenDBHy7Ex0erF3uBKhIy/P87eQArJfbJHRsRLrHSEKDLp1c0
+1hFXCgfeM2sFIxPL6WWAMnuBY4o8kqP4EnCUHvPlGbv/5xh5XW/8Fujea0o770H
BAJbnTcxqBdKqETCOt+tqpt/qf9OOSKxw/6jbHi5yotitnSGe8X+vbCGi6Qrhzgg
U+nd4i8oONW+RnKHVlPDcTeIeqWnPDkd8cP/7qPptY0G7aYE9FK6ye84CbiO2Ouw
qH4QPo/+u6uq0tpzmiiSO6OVqqc9GcfB0xZwKrJGSnyb8kXvKDGcPX/wFjGKlOhz
GpJ3Ju0cAegZof600NxcDDsFqqMpHNO2De4RirTX4ArC8bir1u59VnadvhCx+ySo
p33TwgEeLegj9PpitheV7tYPJPxvF5W6ncc0SY2E0zZYq7vCcALDUTa6bqQTFc2G
RB1dvNIbBVHG87zx7t0DKvZTCOuRyklliLQiV/PJu3lFGkU1yG/oqMZ6I5ghR0P+
mJZbBl4RomzJ/Oqxp1Q1wjaJqrYGN/v4jnbud97/iOCUzjIJoXcHCJvkA+y/gvfm
y9zhR7EGVADWti0NbAtRtdnzrJtL6O2j/EsfE7t7+KstEOyrFPeGn4DUggEr4/so
50q5DOHBaOTuV9WUEcVH094xpXr2iI9RA1kgwKXTKddiJQuBL2omC2OmkizAt4wA
YtPuq/6MKoe20lHdc0R1rLgte+VEeseyLMZ/UBAR/BeZGFzdnu12CPIlIdcq8MlH
dWQIs/YHfiEqNTGt/lQtkjChRPzTTaWygyKEmR2fQzmN0+eh4lWFWb7Qtg/jEZ99
uqgeOAto4SOTi38wYFHGnaWujcduvC70hbKWgC6TVR/Ut2rZJAYF0d9qcmJqeQiQ
rbuuYnL9QvqK0rO9fnnIxmpFq/YyjZKpk3o30wwgk//zgldEV/IVpSUt6LBic8Pj
7lJBRa6KbmD8SyQ4uLUn3fMGTncqhYoiNneBoLXH7K6a7gkAAKRjjIzHoaYbvIKS
AMtlUl4LzWw6xZ+H4Ip5DePujWbhESCwRvRZCrs1EMXR5ehfY1vpHTuiCEkcueNC
wv26eYpTkOSDZzXFgtlUBut6DZx8lPkAgvA7xP76CKSsdqvY2xukp6csicMsfeLa
e+G+8b/RVMmt64xhKJzTNFE7ILdoEcNhpn1ebahYePmfY8SrRYRuqEYO/d9NLh7V
jlCAWxvHMPCT9CV7GtQuOrW9H+KCNtoLRLhRPyLBTEZuLMvZ21oJe1BgTjMOuNjJ
m3qHIY3EG0yWnxEQajdnf1Dsjxbgr9o1pKoEvmtuBZ8aoRvChWA5ubl1BqBznwab
da/RU7QdtluSFfHi2nWqvOCBjYGlmV1b7Rw1UO1ZisDEPw5ymjaXWj2IeAJ11x6I
YBjOczh8uq4OYgxoa0RvhoHrWJ6V0R5w952rDpGmowdPb31oCh+zc7+smmfpCWBB
jMW33PZREMoL0JLkZaZfvuqDDsb+XGdYv8Tpjm/PpyfmhB2HdNjwuy3fe2QO15m0
LSQhx6dQ2w+HKVxvMQ9c2BeV6NxWaKdn3dCsAmzwjXcy++6eYhiM5uvxHA/sj1OE
H8R2hY200L2is2P340ynXgufaCX7B/+bugfMfnkG8NJG2rFGm9OzQBAcExkpeN4e
0fl7gE3eLMTCKO2KHQQqYMACR8mEB3tzPjnf7jWMm/wMa40mS7KW/xA3UrnF8ux7
6nj4qildTo7tbOZDir9QyW6ecx5oyrVpZHs04x1npgvncyCGt8l4VoAxbaBmK6dY
o4KLAxpjbQuZsLf0C7zxAeUCNfvLFCoOwHT7hOXsYrTS9XCwomcVpZuJr9aTkTTg
sPhPmlJSnUpVyNJoZmVx87B2Iwk+QRTI2YnnxTzaI+K9NWFCPNQBI+bOwbCB0OxF
6sS/H/NBPmrpXSsbvOJ5OHMULdwAtaNUWtBoyBIKxyNxTVqF+9n7WcBd1YzbM7CF
OnxBqiZ47GY1GRuqerK3yrTq6G7XKxAQnfViRwiokvdeEFAPLWuRWtjadk3BCY4W
RpgOdgAtPLHgxxAL/eoBi49ibJyK9e0Qsme0x180giyvqBm0+/TjJnlQandsCGnC
FfGL/NysZsWOxKXHEuw2TK81YzUVhFjmK95eDR9lpGOi+SgpB+1JQOg8PhOt/5UJ
/o2M47Xs679Mhe8yDuI6/A6PDqCgXO9afoQ1SxUYWNONA43yGe9jOoeEISCTC+xE
qrcUJO8rmhIGyaO38w4Mqfm16B5AOyu8h0n56Cw1voYxbak1ELpNvbkwNvsT/7F/
k0L1CQpJKKL+0cPPIqFVO5tFgXmNJFJU3x8bz27rKUvThrZs4msg7I1gHl3YzQPb
NECigTMbNt00UKfq4o82VGr/3W7K5xG8MHK0spas4Nmxj1Xw9kjYhrLAoKw6i17R
tsGB/bmydbo99D7Kq6pZQuguYOPpYLwcxJbwcXDC6T5dlCM+vNjVY2hPmlqXpkgL
DYkPXuKrtf+dMvkU4ewYBE/VUkMTaQVOR8r0hxSj7M9VlBn7wxqf2TeFwr6eVoCy
6urd/KEyzdYbU63YO0XCH1YcA8qxLr/BQuvy1TwzSPyqCbSNMNs+QGWPdiFIINUq
Hhyy2Hq1/mM4AwVPGWl8WJQ/L+Wcqzl4iHD6P05d81HSoxSr278mR7ptJ3uyI1Cg
ybg9afVaf/Ty3X2RfytHfddh+l1acWO+c948gH9lNfZJ+vWRztmy7PBCGHa61zcO
6I7qQa6zHA0meceCUYG8f2TvIMlHw4/sOJT1uxe1l196UZ+lsx/rY5UxylNYETKt
5l195yXvcUxWsxiAdW4xgCSq9eszimgS8uG405ZTHXRQ/JPvRZevYC3SlPhaV6CD
CgLC4N1oduF03Q2wK+8a6PWTuWUVi6Ua/6/CVpzFfj7oKXHGzddBmhjaN9vIIkOX
U0p8cLc1e1zQDYT5lI2iizRnMbQljbJb4nNrIqZ2ZcqdlcRRCJxcBhC3ZLIgp1Xz
UUfPTUzJC6+nLm4tJYX9H1ZzB+YUMiXdyF5kTsdotSw/x/y4TIAdi3VUF3Gm9XuK
mBgs/pKvUZnt0vSbdT3BilhjJON0OI4787wct1LN+s+yVxcUySoYIhKZvlwarMRi
Q94Oyjf2SMu0twLqxqWU4CaEvvma1Dz7gLkjPP8s5RsousR9JnCFLi1aAcAzaE5B
HxH4Z0UTQ3FCuFypmlyL97rjLMTu8u694sp7m34zzsifWznlhON1gEGK4qto9sR9
PCjgu2Q20EN+8RIL2CMuVXSoeAWh2oiyxPngS3iLvx7zuHAOrmKkQcKNTiYM4qAl
NWMtX8NJLrH6TEtS7nQmjBNLFmP2Yp7sFsAGRTqo4KDUW9bXnQwiRVtIQkZdUvRY
wI2J8p4xmLIsVRickiiV7K2p6SEj2O9Pb7CLSecdxoWNnaDLDjSzReX8Kj1/WGge
drnPaR3bhEMeM3F/TX/367gO4HprpmcITMYd4EdDG6pfE6mACeRGSTNL1Bj7/rOs
RWDNCWXV5RhZFTJ3NRrBRcZc36E1VH00srZI5fMbg8JeNAcZUDFvG6dBEr/NO4tl
tBACHa39O74Phkl8DJRwXz3lFI8GyQLKRYTYErXcW45xW24I2A9Zj0uTg+rwRokz
gIHI64EOmYnCLKEPxvKzKC3nZ65aFfKoxhwdPY/Lt4ZkZhEYNr8SEtZJwcw0hio7
Tmmr0GK7s9PmJPmHGJ/2RY9yDfx75bhrZh2Ac6ndh7HBDr2w6H2brMMEQgB9WrAo
KIXpj1Si1oXZ9MvxPs4A20+pFSRSarKKduS17mK5XijFPRd2m99okjHaovZxB2hm
gfta1C1kyXQIUSyzxf3UlvIMfUw7Ud6GzS/T1hiLd/vqHiNUas838fNw9nx/Z7P+
3uymKfsPP/uwN11ZMC1CQU3eAV/LDn4gdXIchTfQZFyN25vhFkQByukCyK5qx9gE
/dDLxJAkOKvDPQ6bLkz2q6vfPvETFRYvEK35KTDrkZvNWA+bWgIoYd+JQrdTes8x
F6o6UJTmwjEcy7RkF9ViH/15pNeCzmbXs8VCIQF/WqKI1pOV+Sd1XN1KZQJxtlpw
qjwnfjyZeK2HQkrn21rFU0yaADqtqx2sbW2IHdEAUqPhQQ1L1WTn9c0MoojlunGW
mN9mES7VJJJGfqN5/MykLeos1xulq7uDhT3QlLkJ5me2MPPO1e5g5p4W4HL720t1
KlRBob9TFH6F0iIc/OjLS9pDz9vLWyyJ8YKb43Uo0hjXwuNfzGhiMf/KiggtwCUj
/DI8BB+SFXtLCdZkZ/cDotlXUZDd3P9or4gCe5rRwthRnDAyOCgcDzdc4A7xUb7e
q18TFr97a2JF00ki6lRWBk4u6EMu9XXI/9wN9f+wxYk1u8pGS292rptHSpAfC+iI
3DSThp9EOwjs2/XXfpSt+5jXqKqqMf6qDUesET+LHrwMps365Bn+AFnDpia0OHxv
eY7e81qFSXxUoD9n3x5wrl8DyKBFXPNW/28zNNI2EwuBtwkGKNszpgYfH8VsuNED
V+Gok3Lnn5wvup2ZsOiQ3ibOPG/AF2neYIz/RyxUfdOwxGDyyzqNmgV9NCGcYWPR
+LYGb0O0ZKQ/IhDbjTLPy48bIpJqedbx9RMOkbljHtl/0VWc2VNtXDMb7LI94cVK
ZNyZXKuPn3flORCEpceXgiIEkISFsYJzfp52pE38mF0CI/fcvBt06hBJcSwSL5qN
bjsOq2oLEYXxCaMcfkL8/LPiJ06uJHvpsjkcA/Snj8IuHvCqvLYZanVe8yVysJWG
XcgnhTQXuTUPiDqCSy0Q7vFn2lH+7KNYDlC3j43gEbCwGXjoVPzqGIg2T02cSwDB
O43rmHzPXgL+w71Ewhj5OBwCt1MZLwsdCVGbDn0WwD8VL1YWSQdJX38J+GN0eIVI
MxSDnNZjGZMx/RDyFlZjhQzCL8YAzwNqyj9clp3dYgQPg3JC2NipGTOYZjxBPxvD
Ll6rDzrv5Uub9DPa2gq0CXgtDMtekmtLCRS+7f/MmpLWpB9+2vSHo9sLagYgPjQX
cv3cVZAUjrQ/1gUmEZY+leLZuUoOTc/CpB3El8RUUH0jko8coN70h1nt7xNOTSrl
ILAOOj0YJd0HgeQVh4LNne7sYPXn/g+AMxT7BjBJ6BxhvLXC21GRjOJU3BTLiK5G
qKOKZ/0/Sig4Qonv7enFWPFrD7axw21svMMpMd+W9Ql1qMBHL46FLB1/TGgvmcS7
5W659Ys5kSo5/69p1VvGA7j48Kw31rxUUBa3SIrmMAWc1mf2VPDXq7/zJvrIQdjU
qRfzj8Of5N4l7wcLE5/QWAkCiGNZ48Y+iCfRo+ZhMLiSorgUA5XzjpHgSHQF6qNc
muugYxcS6na3csLyQJssTKL7MgKFIVHOgnIfzWmBzME/Gt33QwA0XphqUftPM3ea
Cn7AWHxvjFNJ1ejlUPaJEPOyF/ofWrRQILm8mfIveYKZ1jijbBkoW88sikqbY6tz
t0sFY7DyAKQNWVxmOQDKS61N7lBucdTUWbZ1wzIoHS2g0rlL7y4LbzKpkBtMP+H3
aCah9Ii4c3C0zIwLpffVV/+hdvavQDntG2+QhrVqu7uI/NnEIEDRKWlNl7i4HkWM
oAfcdehkPOajFjepli177a9UaDuQL0IqwsWI7Q6hDj9SLoiT87g7WjjxLAfDgIaA
zC4bxaypHFs1KKGLlZAhkW+N935Ql1aed7uRT6UkQkSUNd132y+RiFkQShNuqxS7
1BwqZ5xd8LBXKFn3nrS0pek4/3ZVssru8R2ty0Z83r1831LUHFE7yhYqEGf+YTIc
+znvbpjhtdrfiymNzL9RQEp4R/fd4u74obhCI7q0M9KzEbokhMl+96fuD9ddHVNF
7zUmdTvnX1n7t8j3U3E9gyOzLkROHToriSlcxt8kTs1BIsyJMdpcdlqI8xicLp5j
Vsk98NhPmlKhNkjhUl9S2znspDTJHh3YapRtOPBs8SWmwuo5aCKLxvq3j3Go8H4e
ki8GyTo/U5mZ4bdxogt9vpDpgEw4ELmZSzWlyQSuyfnHuoPNBSFksYYSS/4DVkyY
ZGZcbXFDQs937AAQqKB3JLgf38/QM55RNmV0FEeJL4lLSytIQBUTzDTDoBTJoqO4
/xJhELXTe+j91CytRGBU2nyMDqu6+tzvWRRAWeiEvE0/UHSyKUTL69a4zjQwccLg
t+UUnTurasaMH/pwbr7/BP6ITjhMfxBUX/I3MquNzvIlc2h8F73YPIkyR83u/ZQO
0eBE3ksylh3WgT2j2bEvUVCglnXJQ3wtnzcSGXzPLnEoo0qap33YY6WrX0DpnJfr
9y6bw1sF4fdBmuVj6KJU2pnaF4XXnR4WaBBR6v/Wd5ww3k1TEcJg2K3m9oB7A2hW
Sgd2v1cr2OnKwkgQCrRPqtR1y5vUK3GKV1WKoJSVphXiPhX/JL0XUIVuv424P3XR
FiMRPuGaBJp/qJAcsp+Mqu2azDdcbasNxNIzpUOxAev2cPCszLItyx5GQLMoCat0
IzS8WnZ/7Phjb83tnCSf89wepJ6Q50TakwA5jNRJiE8gycZv9te4KJ5aCTwFzRxt
XUNs+ksQkqB9RZAEW99A827RsprmmwaXlVAxB12elrf7G0hDakVfAE2SHVtFrH4D
mPaRpf4gKQHnNp23I28uGlF0nh3SG3JYxlOpoTakIVrRi5J6qATNtgP1adICzLAI
o1qoTZ7RPrWAvWmmcrE+5AinoDgCibyob9vR/0+iK/8uLpH4+sokbZD5J3f6o54f
LMgaYs2nPzGWt0wF/V9u6u5Z/GXP0XcP2fDKAU8bD0rs+ZZ+S03zT7R4m+gFi1nK
ND9yfJVbnRBsBU9QMa0moit7n4II2yvA4quBywZDyMV7MhnygsLElwu+xPVGW+lb
fXVDiSUAtKG3lY0ft7o55h2KzXEfL+D7WdnJ3SFeB+hR+nr/TYEk3Z56npMBNpzi
UmqCxuORao2bfq6Wsvw9vF5asiUUm+Li9O94uZcVfLMfk7X0I+VaZlqu6WhproRe
2f16h20qnrShcHsWdpdO2ltFC63nCojaZ07iBmMDs850GfA13WJndcSIiwVKDhRy
ms7vE5RPBc/GMNiVO7ga6SdnzavLQsTzM21e1JfPbf1Z8sww4KqokE7koVRZQrw0
zCjlHSpxH1iLYo4SWgR3XNVOgotQYsk9xyanVj6+uPb/wp94O6T3+jUnVtro+01m
IH2PWvdLW8YmOPM8h5hNTXc8ld2gubTU33M4ALm4RpgTOvklyDs+idf2iquXzagi
AkcBLvh5DJ1DrsqAw73/Iyfplz2cefmIoLtEJBg1P7YlEMAdA8rnvUpJ7Yr0lGT9
bkuU7P0i+C/hGNV2UKtP59AuwxHTj1TlJ2qDe8NGdRtP0JD3HJglo1b8fbGRDDzb
I40niCDSE5pC+N+/PQUFqon1MWOHCl/ywhgfneSxzR5lJsWiiTpsYOZbZRo/Zif9
YzJkGLJmw4xGITFaAy0aQ+0h7qQ9jJQU7s6K54X5OFDhJRXB3MnxHaQPfIqRf4yK
DhdcXXtlbxLi6VS9X9hns6rNJFYWp67UlRGzUiYO29GM8f3jDthqIQVK8N8UuEvp
Xd7lPS0s1Ek5uNlXnEpE03v1gXZPUbteCye4V+Cl95VDdw3gn2s9GihSlyA4CNpl
xSrnvi0ZOAwBJ60EfOGB+xlu/UGKzm4WRRrjQDm4aPn9BBIvhFIFiGW2pKOZJIax
9qcDbwh1JoooxEhcdO/yutS2pGa0YdCXiP0wPbMMTaMFBrpFpxir2MElFnQVYvBu
NL416y0qIFymquRycxWjy1mrwn8tInXpBnU8Vbgll4SL3Kfu1zfOVZFKjgpDYEO+
BrvU17ONEl8Lj6KHPAuITuIHIo+z+yl29ZE8IBXFX3gKJmVkS41YnJfQKTv4JbTi
V5YAfwxxCl3muyC/hYO+E6c1MsW1x6zUw3xNRIx2s36yiPHZhnZqUVg0hCAs8tBY
aI8Q8KJvb9ahWs1G29NSwH10RmFNOU/x/QQpv/wtRwtebeaVGQhLKNkSctVSn++S
GYfUUvHe+QycAJCcTE+ETK/rFGRCdfCnoeezKEudcL2nNmK3ZqE+LFA2Zd2VXoTg
VrJtXHsUvptp9ZuOVQ0ioN5Ms3NArYk5j8lw3Y4MN6Fe3dRj5c7A24ELvimmviAw
Zz/6WcXE6o0YBYV+G+C14t+i7IMlgkPoeLCTWFpyqBiyXBFr9n/qfCSar1h8j05C
Vmf6SroDbxGrR2Ifk2KK+gdgEMv79L+0bUT3ITuQzNXRc7ABahNhfV67OhKoUFRK
5ZKiGMWL5rC0vn8jGfutxgKs2//VX4bVjx5+m0FiKwDqjNGzYyDUnNeSMChZSDxp
kb8H/q43t+7mQh4gSdEmF0XInG+BC5coQh5Z9yG4zoNNNDvkm2VYLIBVqydbnLNB
NZnJFspLHi5iWXGUwZi0nKaTGrQwoMtGnB4ZN4nvSaVBk0HJXn353MRONQhZpVuL
IiV290bE+FYYS/nkrNVKAVOA2vfpg08E6XeVEzBlnNwTjOk0A0FtKo9jdUA75Ahk
Q+Ay4u1Mmwp3dpWW6Nap5mo2V7JNcRMeaUFYAZg4+xYLcXr/aZi4zZlXLCR/C6I+
grN/M8lUzkAUfxrC+rW63n5A+7VGqlyg2Eh6VfPpE2jH+wLaSt0YeM+MBlrU4Rf0
cREDVw55jyl7oZoDXGQ6AUpgAxDbVVOLey8I5NWl4DeqUWo2Y9/VAxdMAT3PDJ50
NGQzAysxIThdvZbyu/SXhmGu9MEqGxSffO8dS2i7dcgRmKpZh8Xatt9sPLRR9smN
nQMw6trpP7XwampmRFt3Unt7DiH7Mg5SCmYe8J8Lm9pJzA7Pa8fnT2JuRpBOnAdp
lcmnSYaRH/pBjwDJwtP8bs+bRqsNIBZdKM6skahIj4HOVSqpo1ajumDz3FXtPa1+
xr/vEYeNFObPEIRQv79weOph65TBuKePe4kL+WWYKDFRCpVHnqGmgJ9aIS3qDeED
a6SdyEQr9aJpVWkOf6UwPM5xUcmlkkaVeN8MJz1bXvxdJ17qC47YsczF31v+P/56
AEKLqTVzIgkO0EtmlZz+5vOZgkmwQpcnTIQizm9pYt49ZjOUCY6iWVDUCj2QAJ0O
JPOYDDKDtpsKAJ+8Q32Wrwna8mwUmv2Hk7Ak/01awnCFxLVET7KY+WOKIyLSr8vn
E9yzjZCtfH/mPz3/aGtVD2Pg+hhKr4rELdyVKXjArDbpo2GPHG9NpyQcl3uCeSF1
lpGexGZc2q0QBfOvummJ2BiFpEm3pl5MRADLvLaof1bzCq+XE7+rVQEUwZH9J9hi
XFwfxTB5NnOW89tFt59gaqXDtB7U9Gsef9hMK9XnrkAXaYSgI5a7M6DYK37dZsXx
ICf7MWydz/2sYPyNQbUzu5cUlFS/nRtAR2QgI1SmKvOwlz5k04AGuvDuTz66rWKu
osyhFLWsxeMuujTshQCu/Z4Cg/SjhlNT4N2sfmwE+MBtDB6NTgqSpZVn9CntXEPo
bnkLJhwtgw5GS4nQqEJHxUmaBI0nqFBvUBXZtSbTJNNYr55nQFbs9/p3QutQdiPb
0JNUAtml7TUwMJxVRNmgfjzGeDnx9rX1FlRCbm+YI3/znyqPB7y12/P+WkZ8I7N9
rOlW4luxhB7AH9doPKKFbRAP2Mvhtos4JWsa3UfvB83Kcn4oZfnT/JUs7yW0nfSh
DeQKaCfMwhgTwu7c4RMjqg67WIGv+sRTpnW2e873lrVt4wWqzenUPKgbZz5ZZ0tw
+ed5q8+4A6OCv3/vh2K+8vMm0dY6BIMrfmK2qh55yW3p3WMww+lPP+HxEGgMGrSW
JOnx0TPw0+cLKrGoBmPy/7ZoU3Q3MV1jYaY87/0Wlv6+xkyDOChWSZG3uXOYtCXE
bWZlbF9lDeljxFT2q+vQD7opWThdVa/V1yu7k9ZrDnmZyLHX47DLjx1pPA6MYqF4
AX+w6edjgblGfyAHKcMs9eH7t9KhvYMXybPNczsGTv6F3Lf2jx+1hbA6umnmpLBg
LKFcWrThh2QeYhjlmgpzHtkzo+24qzoxjOnYNlq0sOdW8yJkLBiKWFCJwUV+o3vq
vkqtOcj7bHYDXzuP2rqs7GOTTOAbNTPmRUHq1BlgxJLwTRytWD+/F6cjq+UoKs1/
S50b0mXzuvIbmEF/qPOnl/YpNzRAeJrf5959Ob9d75qRCTYWxkeZYvSilzG4kfLs
fTRJj2L4hjGlHq4qG3mFycQpP11ai4BO7GG5XlZqRZrRf+7RpkuZi7HIERM1a4L1
duwigDNRr+LDokVpBiJzF60Gv0N35IxAmrFNRgui7SEb5uy29ASH0gwRW8EXMmSz
nchvBwGBRuaUbXeYR8LRiT3AuGDeTzKZ+eb0QbN/qjAW0mbrTy+NdWW8U/A4pGYu
wkZ43E88+ItxTvERUZd/UiAQgneHE8pyFsWtbLf1jQOddWQdn2hX0yPG7c+wfQ9E
0nYLOpD8E/Xig90w227Rfdl5h+1glWxIi8Rn602EvmT5OXbKzXK57w+OYQXp2j+H
1l6Ro7AmnLdXK7JY+mWnttu0fQox8WC4iAiRTjKJXqnQip8HB+qZgQjrL1gkQG7E
peKywG0Q6t9pVVfErizLSlCEfK3CFEgwtoxPFH6fjJLOEkHL290rtE+A0l92agAj
2LCF+j5kbGM73CPKXKntg/5lSkFIprSYxMQ3B6pmG34Da3YAyZwc8nvWKFyUyGPK
FvNczKGt11kPGhQ4TNaScKB4vAHRTgeJ0otIOAs8eTKssOeosEO9ECcjHtNC4rY+
uaNISvYSyFQQHLLpFJyIssINRyb9AnYSUYKZ3QBdSlg79G4hZfqa+gvgFkKPB8Z3
r2tjUAoVK/AGpxIJApFd78iUvLakGqjyUfeH/roMT9V5djf6hS54QcSxYux+vdPm
VWIdNbNAvzFyd8ofPj0c790oWE7DrcZGO/TXO0i/w75n2FolJTsxh4LqdOExkaUV
McqIX4OfNFz8MtJbptzCvfhWNftjPndi+dIab1oEtGSmZ6Iipfo619wqFJA8bU28
PyeKIyAup4cxa9wktUGtLunhMvY8VLUwV7Ihi080m/wldfcjh6X95dNiXpHCqMCt
vz00RB8zD1w+6SYBfvsWgFdIlIGd9YcDApGzPy7ye0/mFQW/yfkxOgrTdZmc3dtr
quAisfdSPpkk8Zc//Lbn3ULUjr+4BepHWFJeTdF8INzFH9GQM1C8paM4afTq1FZ/
QPweSSkBZ2wcwq+WtPY+oRtrhZ16b4vram+w57r+D2JtgWtDDZhDFJgTdy8to0km
jwWIY5Pbx0XjUytKqh8dLz0A9ez+DjVmKISrNnCsL3Np8ztkG1PKPEdAJQclt+X5
GMM7YIOCAHpEkNOxC9UWgJpb7cQ91/IcY0pbWfAsbQTHq0Nb2RnJhhEtbSMpOz4p
GaErPpZZ+VbHYccbHYHR6sanInja8syd5mboSCmLivTUv7nUaUtBSBr9oSRmjkX/
Q0SOa2i2vkfq+5z8MRE8VBEymdSkk76KkAirKf2ZaJoQxCUKdI+XP0dif3xXKUSF
/YUrqlJEhsPid3bmLkHOdzICu/7hhaKOaOwnhvOvf3hJNOfhYy6VFwCiYnIPqQ5o
O3Q/YrdBgRzrQ1Tw4Hk3rqrsVPehdxvPwrJGNK8AxThYRRIZEBG8UvBxi95bNgYZ
QvnK/pRSjlyn/hdWgfa6tvWSNAliJuFKuE9R+nP3K4safWCK5jklsQSVmfUM2FTR
AD7qP7BNzWZKdHYoTmjsSxGO1mbGlFQX82uCvfow9xMom+QFZ226rFm4Jv/5CRb0
PApf6m06lfmYcRbUUxTsoQAprLGjpvjtLCsOpbV0QrNE6GQrFlCX6qnE6Fg9iFhN
OvbajIO2kxzx5n6q77LMaWONZqjm7eFEm4yCXkxHs7GGrJnVS7s5hFY7GB9sSPrt
fEUuDQKrHKWKbQy35KQdz881msff9I8JtzSkU+dBWeqCg+MGzK8ONQBI8DCDDy9K
kxrNSRuzURVMyuiBLgbNbXkkHI2QztoxCXMQAIVt0O725KLljEmZFrcHfwuBtk02
GvncrhDIzh0zb8B8UakS4cnxRTkG8V1oRgXXFaqnzyKHFFWvGglLoWg0LG3fvir+
1i4RAUIcRs7ecu7T0nP+NlMVIIWKmalwR1ZJl718uiRkKHB4I0+pXOLcbaUJHFAi
BTRTEapWdOA87KGIfC1Pgs+aJ7cNUFzf/kcpkVqIXH2ZwUsFYK6cnLRfj6sgnp/0
qeCRGi2FKgm+yHntwfFwPa1YOMtU7MtT9H8K2UEPk7JU2dOV/iN0IFeWawqWsc+L
xbAN9WgN1oZAePEID6SM/NJ5dmpjLjWqn+W4ZIA3iUss6HigAD1oJIVmZb0Lq5Fu
Ou7HLxlOK34brIsosHZQMPqW8gaNYpzJhHaTXVvAjPoGlsZwWYkRHS1QHdMOiO4N
mCI+QGuptKD/JaY6bfLLYXvuY9oPgm7VSFhrQ2D5WhbeYRX3d3fjwG7oZRrspctM
DJ1KZTgqwQhrXcVawPc73xQ3/lnEhZeRM50/icx7E1r3vKc3XSM8p7GujrwcT4nB
S44jWjVXR6IP0u4PVqdn18AUn/kU3+3Al6wmMB5sVhNZR5YvHTHsrl6wof3J9IKY
KINWDW1AAZ4lxUCe3esPAho3BJs/ZXS6WJDEUZFpN5XHv9COT1lMN8hHk/N/hcNk
QGTCBIB9bnvUhlDqcoAHPTD21U98hWIxKd3VGxF2Bgw85GWP2LNSLon0LAaCUkrK
LXTRLaHv/cRTmJUqBAIHmCqn5bptBd+0u6qv5SYb+wyzSzcbUpgPVvjeeG2PzN7U
o8PMS+GJlzXh/X/lj1l6BMsnGIeqgd/i9hpR+/AN0c+Uq0Da6GA5wn5UvM+1Qrpr
zEE8kupebjwhCxBqn4BJKbVu4EvRjQuTjyCU08jC8aAIXT8E/08SGyfwmGgK97yd
229Yodai/9LnrJzWOmLHsY0kB+vkvqjSd6LuyK/Jji2vM7wpvTpS44Tslh1y3Czn
G0e0abukkbwzLaP8ytgToMgtQs8NTnCT+AwlzUGDJAEFdQZIKwI0oyAMxYNAxNpg
4ePCGJ9tzIeKaFWYN1HEL4zJYIvy+Zpi2b81FCFR94Iw9s97MN7pCaNHXirmcI7p
442kbO7+gJHJRZYoC3UrxYoiULqugjkv66+OyCu7qkXK8Mu0lXfHRX7mnRhwTgcU
DOxDlzMua92ep0ebBS3xA/taPFoV9rpIiQ6hvWb73tEQCNCprFSem7Km08RVnYur
/spJzejy++gi1ld6tQtfY8P8rcTNOaaZnVJakXoz50Dme7+9luLcOolvAOzUlUvs
g8FD+Q51evfX8MF3DI85IKbrwawFaZ7V21Xv90PdlGdLIivhIR7mlT95F5FcfUQE
vgqwSQIbfDJF/zrr4YphRhb0N7Y+cLlLU88s5OldiDQtRbOU9+9zAuBDHYnJynzt
AHdVwfhmg6kv/rGtjVWU/DuBccPhcoI8GkMQuPyMAdGgtC1e87EDMpreI9RGTOAI
wjYwRDvJbpHCtL2XLnM1/U6lKlo5Zw8M/2H03dAD6BvWsKU3N2UFdssnhbK14U4x
5fy4p6M+X7SJkS7u3+gbgrBaI91VFgLGpU5b4ABWFsC0+OUvAgQ/iTnNDAVfMEbL
SqkOyp84KeEY/euovDqXcIQ0/CnjdeU63kQ34O8m9tUrptOaMOZE7biYRgTFdt5h
WRfNIR6FCMYqI0X1msHBTm7H5VgQGy7NCv/aLsbU9jef8v/FJ7ALAyhqXsgtGOgt
VGp33pzt58HyGDBngD2Zh2n69a2P1CDGEZFM3cWkhU1Du4t04CrWmELZQMXLS2bX
WMWkpoYq1+XDzRUDo53w8j1aSs04Ti6/1GNQTjUfGczfWng54GXjjZABYmL+ToJR
PV8mWYz8ZGA9qfxiJQlURlh2jwNMgvakyhv6rnVvx4ApQ70Y9mETRL3Oz4Tb09iQ
AQ2xUWCcp6ARFFeHYRUWsK1Bk55cII5dMTKJWY6vXwjDGl1lzFCeVC2UWVS1acuL
zDgWiREV8mcalYVnnTwTVb7+gNLU/4hwjdydZwuB9Nlycnc7o/X4UYFRE6zI2ITH
y7FBZF9qsRQ5eBrly9DwZxVM/C22QNDQmyqQAFwQxH5aGvoFQaFRJ5r2RnzyBeYB
sgkPLLLFb7Cobp88pGXCzY29HqRoSIVMVjdQFatshYv7hPOhIbLWvsL4pVfatfbo
EWpru225q4KwPLji9Em/WKx2mzdJtokHnU1Z9rcB5EJMvDqzX4QCLP58YOdsfJqy
dDBaBpnf2YF+5IA4KUSGbfM6ywYbw47I6USSZLeev3oUE5n+OaqWQ6oP2N4dsHyv
VYgaQdxi1LgYuX4ZWaHcjYHtAeKhwELKrDQSsMBjAhyAa8YPbdzDrE1uBx6nsSXM
aq53G4zQk61qeWvcrH9CSxvCTZXyLAhHDE10wbPjuvEksfbsDElPjoKV8LHn7jP5
vFO3tCIvd1cyqnjHM3JktEM+Snv12j6Jvg4prsKs1T+RdJbzeA/mpwa8V76HqM78
Gt8pkqzg4NANcGSyGw2j9bWg8k8a6i4keVyF3pLVggmsXWdobb9fhL0u0sKA4X6B
4xfYw8mLm1re9yk8iPbWkgI5UyPIuWaGrjHbeb+aWoPI4b+iLXRZmFk/CR0CPNOK
d1MqEJZuKRCkH9MjYUnANFxedW/4tBhBhpzFMaTpz4Hhvu2u3NGzUvm2rDZUsC0b
RyBNFotewrpmL3gMfF2En5mKmBgMC0dlvxgf2z3xzSfuGiockORWMuJpb6FJ/URr
RgNNUT+0TVSs7eq6JxAoY078i5Kh1DGbseVKuFNeIOzjybdrW4xwGk30ux9IuSTF
TpRwzU4O23XZA4WgqYDwc3xaBmvOQE4Ah33S4Ttt76oLXU7hO8vRQpZz8IaiTW5s
Dfe7auGDeHb+HAoRTRHDQDtIJztuvNNIbAoV/GNaBO8CZudO+bk+SBNb3HodNYIR
8PafDakem6sM7Hn+L9G/jhJAZ7uSJI45T4uuc5QX45boeiCCBdvz+iNknmFMyg/A
4wGbSYbNxWmNBmM8wVMGp6F7OpuQRdZxOclvf4nJIu3yNDH/xuh0r1CW7leWRNX2
FOiWRZ7SzK0MQC22pDaWRGSEtB7uP7uOLiHU/cipB3qQccHqEWkCW+z1niKGmuUs
h7FAgFjnxGnaRq3mudMPAjZPJu3tSYqHyqGl2GeV3T6/1/Yw0zV1O1i6/h7Br/On
NnbV8tdaM/bed/KwRLf1Rxm9u9al6aJ+i5mFikh4K2F/1O9nZCTTrDbrMuII9/xA
JD57lxoZr79R3bRmgxRcarnjSMGD0mmGKLil1y5CYKCURgYwpp0IeVMnVdhSpWVf
145JiIXKEsTz7fZ2TVaStFH3pWDsOijxuz+Rd4CSSvKSgdR40xFPQ+QAaCBWvRUz
SJ8MhD5afTYSM/J+Nrl1vonkYySKDV+vJffK5OZMTdsSZ0emWXC2r/yNiCPIeZWl
JWOLO6AJP4MqYPmyDNX2Ff/KCMvXmOUeNVmLDnM0LvXJDX+89mpDzoJYGFb/6Ax6
vb6rapFGkdb8pbs6oEVVdrg5Gpn1RXrDEby6LBa18YOdeDKCRxmqvW/Ksu8mkLOa
dxI7x4fVymIuT+MJhR/qG8g7wJoY9clL7eH3jZ5vnTzapii2/JtvcZ7sgGZJnPvL
dBqdK2Gs6wda2SgTShl7w/kzYuWqyDnEsNJsVBiR3ncHKoB+SHMlFhxh4p9/niwg
unskZihH1ukcfdFIDszHvM14nRgLqZJMUF359pCi3QtpX5SFjQ2GJNA/C5wq5zrk
1theuynoErolrl04BrEk12iwlWEty44JhxUmRv2ftxRQ0mjaVZU2H32LQNtpe4/h
2V4wO/7+FMzF5Vv31aQ243g2Jx9VsaiwczH8jf+5ElVUFzzGwAlTL7Fs6zJf/9tJ
2DxHw9CXygGtXp1LQdf+rHopymPRpl3rV3SZVaYlrURoBcERpV2CePGjNoVO4DVk
XlkGcPFt3Y+Fx2mtgn/dSyY0w0R6oz3I75tD1WY7QINOVXH3aMDm7LEcjjXkhQBC
LjcMsUy8b2Cy/HAXIY/gqwNEMHjn+nJR/Ap0rXGflpR0BtqPglXjve9hIheLUeuS
1kDdRJMkp7VaSDmSZNBs+RsWUgIKqz6KyR+Vgtduz2IDwHyWhLb9fN8i2Cv10aCE
2VhfqL0LyQ7j7qOKN8Ftq5CS21h7+B0Sr13U79+clxyKh+VJwC8rw62ObMUTC7qz
HALnc+4XvaHU3MnQBPW+2MHYzUWvIYpJtpOQyzS45VA0PT2WhBZHoQYCYDCnFgfw
Vs7YvYdkQP43KtggprBBx3KqCLc0cpyQB6ZMlGFY6ZKjx526YmXJecLD00RL+Ik8
+uooLP6XI5OVdpl99DQspucsxmmd7AkuhGfaVETz8/YggeoMzLKgspxqzGjptix9
purfbbnxCidkqSmIybvWfPK7kTVKEP81HSnI6/95/EmqkDg7dMywIqzD9WAwidGO
Ybbkt1iGTC8CQNMwDzGv42O6DmxvG3hmYARo3Nw3tZZt1ScrJpDATu+qOxbwyFL8
vhanOqHGyeY3n076ZieH3tAaJiohuq4SJzBJbl0qu9qbj49lRqj0eFcJA8iXRNds
vC2sQFzgcjZ3MIWSeHvSCU4/HqHg5gwJf3skdAhPDBrccGpBT8ikWvkFqFDBWTII
03easOBv1K6/1o0BG0Q6g68ikoheLBEhshyc2E1qY/GN3F77nGviJIjHkvK2FU/F
xiNkYSK8egGkZ3MxVmh+1dkEW0Nzz40qFxHMnIkz4mPknq/oXaj78qUBx0oryQ/s
gnCbjA2Xv0H60riDfGfn4683JA0eaIl9uxaTFtk+XHiiyg6cM90NsYNHpEt//a56
ljf7V5aNQFdpblnIIP0St9ao2l89Dh62Ej85nzjKAS8uXeAvdWyPf/4v4dlxe8sl
nsPDuTV5SHallbGIQqHn7T9WOq6cWHROEghe3lTFDO7pHUWcHGitfHUGBYPI+xdk
crnXaq5XEw4bFYke6SM/j2sshhGrnU68gjehcnX2x9eF+qGfcsB2EV1MI/H3G7rH
HBCAxXqAq77G+Pzc4IhXGinxS7FCJIXDkzdbzK1aXDnoEoGyaj+sx5kPxLmm4hsG
pDDMW9QWcziAc0VbbY9a7r8BkhDsYpw/PUpXzlIc7UXit9q2VmaPMyIpRWsOJEXY
deYpvJMZdNK2AbPOyIjHVf58nMcauXJG4vLFeJuZusgxpQFdmtjrOGeMcoBjnPkS
FpxLjPbR406bsnXWR2Pm/PamgS+fTmFcG1z4ZyxD5D3acAMWirRlUDEfp17V8ySO
eKwtM4Q66g6RtLfzPsMBmE4HjefpYrLeVmbhKt8rAMwoNcYSZkzqtl/M2kponWFP
8Z18Ky/CGGvpB4zuwVbhcXifv7jiTOzCrYK736a7NApBRD7G7XR1AT0dcw9WaNjd
6gw34eG+H1dAI6IDzk4s9RiG0FvBm2itcnNAh4g7h/3PotT0FWv0O/O0icKXZKLh
fQiYRD1NCknTVarEw4QTaPBgnoIMNwiYX8ip4K8ibHFPOTALuKya2pdSL6+T5SX6
u/GkVOJR0pvDMAaIP9eQus4twvT3lGJUT0Zttm0FlvxLNB+bPEIqjGTz8mz3ob28
5ohlno1s3yKVYxnXs5WXVDwn13wLl+fccn3U2r7daSxLp6OC/aIbVySDpucALv/D
7nlG0eDHkz2NpMuhdfGXYIBU5o03vpJsH+ngaNayhXBukjOKWd3Hal/fF09SMFDK
Ot9FITs4Mkr1S142IIyGHGmP2N0oHyDD8Z8rcLoIMo8+f7nkGWqmKe5Q0P8G+qu6
ELDLxknJRlyCcu2YYcbHVqWfULEZZx+PdTCtTVH2cx4LFcC5NNWdq2e0U8JDr6kb
X9jBrUyoq19m9IodZFZSrNohv5FTWt+8PKlBi1Pu7XKFD6fsy4mLPP4wwndZxHGR
pTr4g0vIas6S1Sgl0i4AaEWtbzOfIcPEOQyl5zEOtGIHTYe8XqstTxZ4LFJXOYAn
KXDRE8hS/mQKgFgsjQAEkiZQlexS8BMkCB31AoiEulBNa2Topz86dI/njvfzOklB
LF019298cTio6ymsjaJ+0CC4rxA1t5Mg549xJPwFgnBC8vMiNAa0S+i3kT/+VovY
q0JWbnzcrnyHSikHNwfO58T8P+jC6mxgdIcUeyrIMysgv6w9qwvTesTQ4I9rcATA
BY9PaMCDjF6npmEYJyUjN1/zzEE6JNISUMJ6WaTHprKHPpPIDRS3Eu6a25ICeYaw
JJN2Z+BIbXh5UBl9GroJMpOnmPVHnBC6WCUkHB729ScVAjtvWto/3pjyTxxXDhsF
UVV+3GgWA8wnm4B7GtpijAVXmArhn/kSA4mgHSenVIqX4zIsGo3P5QsdMqncDnqS
uYBPP4mbNrxmgW0fblsih1lintkJ0bE/T9Ms5wo51+kOoatEF5akY2RV/51P43qj
NBdicnIvL+dCMqJTNVtjj7w4MUSSWrfWUy6IGqPVL1dPE0S77Cphij6Y8rmZ89xt
noxZk9BH02MnMPAiXrqbL8Vd//r/t3eml4cPP0pman2/4MsL0ZE+9B133cDBEIdi
UQcBZs/Fvhf+2pktavDocO+MO3FS0XegpejPdgYj0zSpFY0K95WtddKLI8VQmmVc
9A35wZuMMvnXYpPV5plXAHY8/NbsE5BqgG3cyaQCSLTZY0qFriAx4zSp2j3S8tEr
c+Cg6b+wbRywULFiRviLfnLcweQfZJ0V0L/0kKYdjhk3D0EpExIPQwxxKeSL713K
oe0tBvQnnasZtxMOuEwpemG3Kidy+W5jQErd3fXP8E/TDPJ8PNtFpV9pABZiChe6
CLbYgpYTZFRr7GpK2mEDsfgI61PuEeno2TWVhw7ixXe6Y37si7LcxtJQ9Vl0dzdB
mVxU1nKQ7L/nP/i+MBbYOHh72ycaEbBUxJS36OWd+sPlskEmN7006AhW2fj32IRA
gsuYJnulY/k7jkSohQc/MlOHtK7QbTvW71gstejNqTCxatajLLDlOykSLyotTVD6
5c91IzmGuth0LsJeZOvpxjBd4VZiaWm0Gac5JzHz7OzBrNcTgZ23KalULrSWg+nN
eEOtPQfE6fKZHMjbwrMcwkS0V0LXG5NAcPLPEqmrrBUqfSZjZElCNXq/zJAeskmm
QdI0ESPURrsxbPJEnsJH0tvRGMLY0Aiq15VFFdpcUoiA2MqKyIOBJDojb3YB/xUU
rbn0YqOolyrhc6c9Kd8x8TqyrF7BTDSWdguswb8lBTJOdzQvG92mL7/4TOzLUahY
5F3bsQZOhceK3Ib8zWhzjUrrBtc9T3onnRzQTJys1Kq1Kr0FtJ7Dp0fXvwF/6czf
eH9RCrh9KWBGw0KyiBUtSuN2HrdD1sY8P3BQLjha5u+Vvb1Cf/U7U7n/msxTNOF7
oX+/a4VMBo0Km+yrG4taY8H+PCe1uSXTPJltg3wIxgLQjNrtj0iQ4S2+4K+lVk1L
LTD0AQ7/jp7cQ/9drKg+ZhxHeaF1HvEpoQZPgZeA9+AUPMFMUUY8U90Wzm0E1fhq
2YKvExbME8IHEHX8Wu9wKWQ2tH3yOu+Dv+4uDYRTa0Kj/Of8QS/34nvDMVuQzCMD
3bdStGQngzlGxbZ+kzuE2J6YCDpbCKIfhdd4SQxQQTDMg56W3PPBJWi81ozj3Lcn
NRCQrJKMdhbecFL95LMEvvnUKWDg84Up1wzyDtVCTvEdkVmsQHWwxv5M3mC9IVtH
Lb240oH2f90eDi6hka+gAsj1bG+3Qp/yQwrGQfvQdlLCQ/7UmIHNVsnq43lGy+do
Jb9WrVPokammXdvfraF1nOhqfJoY6wXVHnunPN/hUgE/YeDyc4XDb2+p7wA/4yzI
tiaHYFQEtRzA6esY11nregGZ9vcFgMhRAuE49qsyay1u8krFrmMrfojTOBqAli93
llm/3JhVrSaipWHi0xPIFzj95Xq+DQioucJnPgvlYk0/BFlu5vC8yXTxPkq10ltw
x3YXw1tv/DnW6RgW5ctF6tpRVeVQinRuKkwndKlv05HkaqazxSnYbpPIQBPy1eme
1YJDFHHpwqec/UY6VVTMCQg6fMCbae0zagEl80Bk78BXTirAYa6DrohqQtvKK3xn
4D6m/BNXAa7EUnflHQklYR14jckSagmsbG6YfDE+j+cOXnHBpcrnYTIQ76N1p5+4
YMcH09/HJDy8Se7Kvqrup56KCALuo3iHuVvlJT/15d+RSg2GagDX1rMjmkxuAvEC
kZwIeysqZQV7V0SRFE2sdhKZLUJd9QwcZroEQWK4jPwY4qzU+mfwxDZuJrRoGxsY
FochievVOTwynSvmk0NTndJ1PdSorlbhmyw9gPO7lNLv2UeqfXMxAnUzZ/7qkYQj
c3qLqJESDOpDXEffMZCaU2Xz8j4aarM0cdwzYLmyA7Knbd7+u4hRReXThM1/7Gfn
hoktnKIRJMhBk5OGPO7RcHsXq9pgp/MiqMwUywV3Qf25CJNsTBlICrTrDp+Exh1s
WSo6wgqipzw4paWBK0/x3uPY//Id/P4z34QtGxpaZXuPZITbovvApRdEBZFbtzVw
ZZtouCT2q5lMIF/x7O/GcAAm0Z8iU0AiDMXpxb7dxIojkCcrJLNQ4jIz9eSs6VHw
cdQ3eJRwtycsh+0x2rHwqzdvXDvpHo1dIb3aP6tM2+SIGM3L3OGxsjwj+nEboaTo
g1RumP519n8BN5NUR6gIhjKm6B7N6cgCvyvaLmN2N95Ta6NAWwjGpNUokMQSBBvW
YvBWeZ7inNqF6YRDwesye/sXl9WlQNFExrCV5MutN1wi9/MZjSMTpL02NgOg1nQI
P2Rzy+nzHEMJ45yAcokkwy5eGypjB1vcS4H7TkLGHbgMTVs27QnhJkZ7mB0suuXy
xamCzSbkGS4CLlJ8IxrpgNaD8YnwUz07Oh8h98Aj/glmRvwJa5fJXIJAXfLLedEv
ZE0tTCKKynn8WRkw2xHmUG6+XX6YBcSo8qmDi5xISSz4DzJj0zCJONs7opGbRtQc
pSKOfKQ8vqhqA4ofj8Gi3uJLP7AtTvWO4mP/RYSQL2eldX37LTmXkJr2J2FYf/DT
JivOMRnYxHvwDyNalZEPQk3iHq0qE3I9jlolhZUrWDcCeakIIpRP0+fdBP0KlgBB
UGJDUPz0ujyeU2NYPBroTjk3bGavkckvKkgjsh7GgXTlEFMbZgX1ikM1dqdjm545
q/motHh3Wdc7FKCEPy+m2mFGoIGTRUJ//PCtJeFuSowi10IFUF6bWsVZ/fRH/0NO
9GsL9Rd0uCNwzLIhTZjxzhUq56+trHBZ7vQK2aVASY02H9qFcIQoioe4tBA8zEYW
LjsJm5kxuKOJt1Yblit87fphYDL39nxM0sYamEh4Yq2rrtKIilEROoZyVb8zp89l
XfQIfxaSu67F8ME2xNTUePR/V4y00WqDb/rQvSIVYXxAv+NDl/XXa9PQfhgUgeCP
kFV275kV6mTXbO8hAdW+XQpX+QKVeRVgRizrLZT0TGgDmMu7GPc9gqWSGylNkeao
opyL57212OU4jMLOHW5w+OWkrc8ymn8KyyjFegN3vdzbHzdA7sSpwQ+fdPjfDCU5
SZUpv6I8IvuPl6EUYGnb0LoW6+iTne2ewfwW5XOLhQWQjrrm55NYU6NvT2mywFm8
DfLbF8oN+6BTn0mG7/dDZQlA+ZMa44j1irGbgQZVeMVA1EEybeklH7Y6d/4ouclL
jYkPgbjbFtR5teYCLpKRZsfKg3gkpluoOxp+8uIC3EX6SFIhtpDmveu/kWI7r09E
l5Py6WmgMyofZ/tI63Jj0O8149/USFl03z5O2isWcmnDnp+l8NMPfEYcwdY/4Jqj
0aOjJbv8cdOObOVEKJpXtoYyyzWyQYkbFP9nBEwLgQBQpHb+zF028cSqY5+Uv5uD
Ul6rN1W1VQUriBsp1+eqp6EHS+Mx91JYkx6iMiuF8irUBIW3n03hwoCV61GM3Ta6
eWlSSlQ2bxwWWKkVomH7ZwbbFnys68SMy2gg17xrAC06gYDcVkoL4jjnWOC+F1bp
n9Pyna74gZF9NTZOQ2dInO0sShswB8lmOh29YGMcBh8dFqaZVBVLer1ph3/Qz9q4
v+D+X48yVYCzEpH/qkMQV9oZxJHVsb1r5sel/6VKab8D/zrI/kIngB64cFx9e0sx
/+AECdoQ+3vrVNBCX9Jr0xV0GbGyfBQBfZsZeyQusza18csWZzkQIQcBAse5vt+I
5eM0Rs/muyVFNptaEaIIeGT6Y/tgksisiKdLydzI/i/sh675iCU1J4copIRhlJDI
x8bDBtRvk7+zh85hR51tNAM9bblFFqFbx0diyON+siZJjC3AYBxi6Ftr9DXLOXfp
BOJ6jskK8KaUQNmu9g3S3Y4EnFVL3AvbNXNeOJ6uCPUlBB772bTidSq6BMzjfjSL
7JoMhMXjSuC4xmPSXILmq3RTXEtp7jcRlKjwxSAtzxrmsTTI/Dq5sBgvLjxYasge
FdiIMiCF5SwbmmRUiTkpriiTe4Fky8N06ma9EuNvc7W6rirpXLa+iURfJ4aDBQp3
dIiPzpifihFbDVqBxrxs/m3XwvW7+uYgzK7RKNJb8lc0O1nAqWrQECQUj9PHVhGD
f2uf9iD1ISpeIzfvNeDNa+OpAPa5XVR0LsCbgZtl8pLQ96TYD9pSP4SrSTTMI5sU
yfOSLvd+SC7Efn27dt56R6FevDofB+p4wqlfQhMkIgcbtIR6nkdaReOvDQzwFKV0
PO3CQZDnMvNXpM5deN8TQwKF023/0yoJnFS5fRuk5AcO+BIjDJKP5GZ0opZpt4Ph
ZRJbWp8Z3txoxHqvpr9FjQe/1r/Xeet38dWtdJ9vLJS5ewHVrQalkgdlT3leTHee
yvSYnR32q5WxYS/l2xcotHIZ86IP08LozgvnlV0j3kSjyWSBsiFE5fc+r+ZHzysh
sbSO00OZkvxfy4BWWtJA2a6e8TJAaC5HjhR/G5Z2fxuYb3M+lfep4OxfPaAl9akK
Zp0ALkumx8SAemWo/24jSXLHYMKFQR2Hct0Kg/94cI9diYnvtCVfVC63MMEW2BSQ
vOgVHpvq5+tRgGPCGfAURmAuyt04firAaWnvVr9DBHgIJyJCGS9VK6E1wgm1RKiH
XEMTx3lGMqCjv4Rve7X5fu/q2QWrRN/HCIEe+S28y2KU4BOb+XtRbTjWAaMXsuYL
gJmGOxjAsAFfLyE0h3wch+PAXLZzVOkfRCNevkODIq9z8FkCzSUk7JX9reHS3Ub0
ZNUOQRUnDUJ4DwR/8qFW+fn0ekY6QjwbkmduYD/THxG7zzrSKLt15sLG8UBjBol5
/s38+HHpD7mbtnnn4hJ8bNoDtqbul8J1twg0nxpRu0uaygjZ1eHvydo8Zmz/3j3t
wkZ4dHbdrI14fOFzq1F8eBjlaedcxmKlNqT/HH52zlUnUa+7f08fdBPxmD+9yzzC
umj4Zf1Hv7yUQrYG6bWITV1/VpDIyXSK3GAt26jlsH6Y3kRyZP9WVfAn5WbnBAfI
lKOEKjQBK7fbXmSXLN+YKliISa6Ahvo1f5PweOpHmPJMSnZmf5x71I/oGXCU+u3A
66IloNFozLyk5eJRltTB8fv9R7vAX5hE0iQv5ij2fy0yFPTrOh9d0ti2DB7h/kLU
nTcwqPbmiS35URz2+dMcAVkK9q0y5B4UyuleG9fBo0CpWY7e/l59wpE1j+gQ9Fuo
Ql5VVWsy6NF9op1T19qW3sVSj+ujYWPLKqX/puiVpiKEHMFjCGQFRw844XGxodQ+
+N+hGrlWaxLWBiwud5uLCxgSBO3PTE+WzkpS7YW4WJok+AtvmQMQghQCMhTwenvH
AvBmrt6rgG+Jm0JvyR7JSgF/EfHPv96kIyNsBALS+wN/91dGEvkLqf2tYbQI8SxR
tgwTTHTPj6JVMldaYeuL6zMYJbr0s20Y6j4b0Zfym/mxdHhivTDxdI/lRnXMZlrD
HF3KJGP8agYlluF5308bUHoQTGDchOAW0ByPsCwxaxtEQf5NJOQluJ7PmiJGc3Fm
G1QOB25SHl6C7iSJ+17vGcEejZN1mmTDdKkQmESKDGGqcsaecJsRnEdTBtbgHOVO
A5QQ+KWcetd37ikcSIoCbWBWJsUm5Aa9+VltE9hRkn5/JsUftEEMPfRmdacI5P1W
vfEPzYyfJKcQu8cQ+21HqxMvNjPby3xfYy+Ut8Gs2D+XIBXlBnZ8CpKkfAiwBVxj
F3CSLIIOYVzqHndLLgXLYXg1ekaT/lt+SiXxVcKyrmPHZxkFSh6f1QSLMfH/H0Cr
7flkmLxUNmpauYQ1wNYSnpD+QngIzibeHMPWSRF/QoDdr7znLO5mj5Erf6fzSPkx
ugiNvMUJKjgMfMziKky4nd9ebxZC0sx9WRMTHkR6wroRwgLp+ewbnSFkQf4oPRL0
GL3MaUrUKI6i0TnWJ2TVzAuEo156g5w8XBnLRCHNA/RafL/2Ix7WJ20/9I/vnZyr
gq8LdawU339/Fvb4Fw+kW//ADcfcWpsl8FZExBLuI0F/aDfc9aqCsxbgncx6Oqbs
6Y3EIYDvuHk8O8guZmoXDJYW1ffdvT3bItaTubPdHrBoLRro/skbHgZY+X1XLmxK
cU9y/YfEAuLQEeF/GYzu7CmFGEbx5NZ0dSYJkDPKcR4NWKtMpkxPKsnixJ1I5D3A
mGVTKhxxhOr7G06AB1xfBxCeIhJDPRiklU3b48xz5f4j0RVV1slqlP1MaT37sQ7z
OsynQEsClhrI0DLNVQ81boVJ4tSQ6tBLORSg8ptRNujsJd3apigCuiPzosc1LoMr
iJgUzjB0wqQQM16vbzkbRkdGkVLKMYvsVK1DCmqCSHVhGrzGTJgC78PLXPVlTCL6
i5GoDG1wbTQucBWmQqDur/4s5/bMQbn7xhkYs3F29aRzpG5CUwOHhezqOCWadC/i
RvkEgYijIYupU1P8TwrkjerdqH/gsJ4eGAPz0FMQ5lkf/IuZi/5rhkMN3eliGWjw
m+y1HGz+1E+J/75TwMVnSUIrE949t9CuaBXK3e3+VAvvkpGq7c+exRcxtKadHSsk
StwUyVbl3HKdoUjPLInGkGChYRKM+foWHFCU1A0ehVNnlIsYFun4qc0Nm9VQnyCG
O4hn0cnD/crwX8SEZ7ENd4K+vRZuTqUdMBYLy+nn+Xo/OoZwoYwsJ2+5NPE1izN/
ECXxLHAEu3qPqQFiJU4ONc1anBRLGo0zHL7dCBGtYksbl9qi9kzR05g9po6+9XpI
xd1mf1FllJ/h8grrlT4zGj8Yv+w7rHxwEl2UlaJRjXQI/mNUw1qmY8bSMvtlqfW+
BYGhESVW9C47Mo+bW0iax+8HUN7dByN6vwj9xkn0Qr97UXle12FlZ653pZecEt8O
ZXcy6nPPK+C1d0aMYUihISWtDn1L0eP7LS6NtrHd8qX9y2hSiiciclMq/z6qP50R
4LLZEDHvIt2zv/2jiT6/jxLvnq4gaADGzmB0jOwQn7+FvKAw8wjps/bdYgVjlj3q
j6Pu34kwnmg8NRtOvdHr6XVsnUPPpEFuxBYN4W2pa25jF6tzOWiTb6qylevs9VWN
E51wOkKPigPnl00hCs3M8wV9xybde689+ns9s/cftzEx2G7gE1knzJteZJ7Uv9aa
qjJF94z+KKU0f9RC0UKKU+mREO6w69vYUlnVB+bC2K7S+/4z8tSAvgXxbq1lwOCh
KKe0/ftCES+BxiA16KbvZ2g0alplbjCfKHHopsBP+pA/W2a/J7HPzhnw5tFQDrGb
M9nkMGwPMqKPJl7/Lx3R6VOX/92PH0ySybyzteseZ4z4FXQ65iAAKLcIzvAVS/OK
wXxyMyv601AjLOTCbPYdHdbbzGIVoibBWj4r3F/vHRSg1jEuJ2AhpNZSkL5CShXM
blLbu9X1f9bQfQt9olQpYLst9eYY7kxX8Fw7Xq6FQigP19eyIUNR5x5/HL7yRjVc
jQDqIatU0kRXU1wIxD9eqIV3TCUVRVa/t3znWxUVxov7AWFXe7GToGdA6AMjjkLF
RwiIyzK4oDPr3of0qw5OzrM3RZnRranSdVIegLO/eatUXoGrtxaIS0RP9X2vK3bd
BBIPnLEZDVN2vGy/VPtiLyrw7A24teiELBZv2Kj9kTiLzAECwFpQE93GHMZUeMKU
fZDNi5XqMXjlo9UvPQRMD/1AwkQJeHdkQUAqN0hsmbQuJ2VDT+uc1mvjjjowUeBq
5/kXm3WbXIV9yoNTZox8FOglU2STypcl/psUH7VyosH/eZrTrOb6fs7UB85fbnce
esUpmpUQHhBYwy3rUAqCPsgzDitH2bbXFcgLjE7dH3/i9vD/F90bG7Y/UMMp1XVI
FYrUg0Cocm6MD6jGYpxax8QKIQXE7F22N51b/c1dV6MW7NA8wA0GJGuwIFzZTie3
pVFOZAgvgjohPA7WeYRQ4ag0xunxFQgyUITsXQQGN7BaNJbBsCeat8JbMuEmsMHN
HFm9it+quqDcFD5B+K/+jdHmLXfqZ292cLbwLjgoL2cVRQAKXN4fToOeK01+VYhq
p44yI/5braegLE48KD2YMvPBbzdjtNUUe5kkQ9FQcBGf3asL9jW00kP08XdiuPGh
P0CxmWOEY/pkoQL0fzjkz5bgJGhADeHqp5w9Xk/hKC279wB/81FDweA+XAoMyMwE
jCnVEpIW83O5rmX7oLSKxKXZv6CXQ+u3G/LEXc2wAye2jd3FrvDDyNrZtpsBVQ0l
Ge3qKuILBo5PttAPRQ+n/YGMAtKo8G/O5/UxcBTTHJXeY5JVBfLJxQxQmcelMDKF
JtHtBYJ7Fm5mjevn5Qy10zVUC0U3rztpv6q0/sNNwy+fF4eqflk5IwbEiE6/AaIm
qPmzy9UgC9LxP6gxOfjWIW0Z6fNB5s3awixYw7W1JPEj8DL6jEW+MQnugQV8crkY
nXTsihJsERqr6sn3xm1w8jIqYTHbtYauB/YlMnahxPjTF+MZXojkek+9tGdsk8RO
Owka8vGwBiDMIf0P8PCmy3jC1Mr2XTqe0U7mpUlFR7nA/+dw4rDCi68CVQM1cPZ/
PpCEIIauae4ZSgSjxZ+ze7g40vcFerXrky9sVNE0sLipPOzGGIrQhKesmGVLKsu8
Hbx3ND/7Yq4t8Ge0s8ZxhgVtmscW7WwDlsoi0Lr2f3HsIcV4ZfRtK5SGltP0q5vi
2pw7Us6bKvzNwOldbFzMp7yhLoJX5QvLsz6Iez1MVKotHYxNMQcUFEN7cRipVr1+
47RydC3OWGVHLycghkl8YtuwGdkvbL7IVx72hfk+0zxM32Yg/rXu/Gebi0Q5Eg61
dG+iCs4odm6CLVaAyJY1eilJTME3mtUNa3KxCpZNfBH+3a5y56pr3i+o/9TygeEv
DE4r2ke4MrSHRLtVf9BfexiFHhrfD6SSiAxFveUut31J67HoKilr2ryFAULbEoNA
K0Tv80KrJiG7rT/DHddrhcX5FAq72A+drYiwCnhWfeHYlsR/vSRKQVnOtWVrjxOO
9lRw3NDstm4tKZQB3jLiWj2TJbCheqMhSGTnB2Jk7WPwXOXrWJB5q2XcXPMe/Jfr
4ximwTM+9l/WYYj8c1g6aVo5RvXTzWej/6JU8KrAc6i8VKoryyf3R/DtgMzeAyKN
7oLM6JXGWiNNRB9fJXu0+bX2ksSYoegFM3q49M+T0u+IRHsZyA4oCr57A9711Unk
RwNQyPPbYVt3wSEi/cNe620EzF6K7QpFRHfWaypGL4chpl+VxzYxs+0JthF66ZiB
4ggtY7DIpDOnc76AwOkCMy0ygGHK0lVPW8XAAmh2wTmhGfRcvzVzQc7ulWxE8H1o
NQULSOZPcYutjYDhDYit2hcP5UbJy292tRH5QVwMHVExArh2Ez6OzBQl5Td3mzvw
FpZRSqadvoyXH205v9jHVB1wCuTBmE0maTnQXGQz6qU5AawEM9FVaK4zGJNi9URD
SsGO7b6VsxobWd3K9Y76Xmea40IKGPkgDbdi//OEGx+JJDikRjuxdsng0kk1nfEB
DmvOJQjxS38qEXVL88/GDe6Sg+XhSRuOJHuA/FvjzXqlbV+SQux6mKHMFQzZsmrO
gOXFMY3K/BksfZtnPpT1LyqXel0rmko4XHVpuj92pB3H4Esh3jouGiWj0LzAny4+
nMZpT5Mp1T+AE6sqX0YRS0lWtjZBg04w0tGTlsbRYlizv64KJ5JeRslJwK7yliQk
Mkrst1E5mcoE6j+jRaKNc6r+YcI2NeeNQI4MGj1e1gZFUiiMTk+QrU+s3lLkvKNs
Fd7+sG8HzKuokz3AzNHF+6L2dA3KK7Qgcl3XFnN6K0mpsFipV+jRHmz3ZNg8RMNI
D3tf8iKz9JgEsN3lIE8KGjmxuNJxkS299B6CYkTK4+POZ2DC6y19MLlTJ5A2C6bz
HOovll7q1WlVirkfrqSFlQuQxXR0cRIWF/1bOgBDaqKM60AR80hyoAhAKstUnhEC
uhFOnDRfnShOEyFyxL8n3dtsH7RWrop0hofOcMiy9ddreLlcBCcUSylQernaZJUC
Im2TCZJlvdh/u+DTMB47CnZUSXQLY5zRoVtwUbWVs2C2n27KzCeZC+0Yf9H9M/kZ
XI8C+ocPbY85IPKbBKSZiZ9gOg5agg1FhJClCjAOY6S+a2qxQrPFkirpec7vYL1X
OO4Ys1Sc1idCv6yTJnWGjU4LFJwaaYjg5AgyxZI9/zn1dynDsZmW8IGCiKQdnUTf
A3LXUfY2Xt0OI0lSaD880fvDt+QOc7cBJEqVmz4w3Iv+tQINKSTxJvXasBxcVAXV
Yh47EXMQj9zppHje/v5mlmPm9syyBw+LrUPzMz+Snv+mRxVAE6IJFHlQQ9sZW7XI
+bwEP3Ll7Vxe5W3pb6ma/oqhQ1AZ4WxXRnnS/FJdPNc28eA0aAXi0FMvicoAvuud
83SjlGKITdv39XaAskaJadU/XFx9nusXnFq4USIASFUS/vk5kIde7kDWRErtaefW
CKrx30gNq17RZRYn0TFsl0wwOtZ1v9YSEi3Q5XwYXli3KPc4TdNegFKVOpQqR1nM
/d8svae5VSv2vxLH6hzunHWTez4lN1G7k668aejbaRGoRk7xRXSNlb1o9IO4jP5T
3vNemTmZ/+Vszk+0aMNBNvI5vQlp19j+B1dlwLdX+7MuhOhVNFtTk5x0vKobZfIa
1WBiSZb29+Gcb434RYi6vtgx10WlFIobasIGwUoQd/PDAZAM5QpHKw6Fql+JfROU
ste1IxnHIAk9uktHdTHq6eTezjNpQL7oeIHpMV3X1nyoRjU34g9iarMSbZt/SYSb
VR3qu6uTq1/z5AOE6nUKoptf/OXcLCl7VnDURJuFpMb20NQn+j4c596r5km0WBFP
o0efMrfZopiImi0HEbDQMSi41uyRiQvJx3fwkH/eZtAq8YDxG6tIHhX1gzzdiIn7
vfl4A43pgbQHtv7wEBKtRc4k/710vpTYxgKLeZqWBkNy3l9nV5J6isKIft+jDYq0
smdctUq5vFDC5zYQQTMbcpzo8KKaZYUq4FfpYvHVXSwrq3wFdDZunSOLmVE7kjk+
ZEJYVztRR33mtJsqY5a09Yl0L+VlfFeyjMZNmArzyoST8BRn4TA41Htu/lCXC1z1
2kwr4C5kDGWJK8ENzOo0HmxEbqtIstF569bZFU02LpE66hIiea0NYoZFUoQIPoca
a8/aknaac8phPjvOkG32VWXU8yTIRadPNoIZ6ccedcregLKvvUWkm0DwwQuOBx+P
jTaiMA0KiISA4NPu1mgAzbkq+96JHoy7mZ5iP5QitMqVyvJx9DQt6VPp1gJuA1t6
MaJe1t+hEFRq5VLHkpr5t+E9z/+R6CpBpSPu1s65LIKazr0xZc3uLI0yZhKU+fFA
qQRpVqDON4qmHDqFgwFWLgQ2KMn19ux52Tdqv2tHfPVDEcuYwx3YSzpFPkUmDlCi
RvDQcZeUL9vEkgLP2a9XTba0YV7CyQc85nDdUnfgdQ0Gsy29aS4KFwMEDu0Sn974
nZSSwaz0yWuwtAaKjuqEbJDoCoO8HciHLz22gK+RdJPkUTCsLgwMx9Bo9OWL0L+Z
HGNwAuERj0T7ij1dj777hxE6XOa7sUaAajdxuwiz+uLwzCTDItS4mlzRm+A4M0Ek
nduuYOgUF508V5Ro7UOFZKBNPhfb+b2eZCgOAjEVc/VG4AiPDdll54AO54XGoXN6
ZTe2P/z1frzjN3KsaSE76+eVGZ/Kgc3FnvmyR36LkFRALQBlDwthloisb9VH9G85
Z4SNQYWQ39MflK1fA2Kj2/aihL9rb04NUHLxNZSFMShYWnPGDkx5QnDGxb3bnsY7
gG8D6eY2bW2ejel1sXS1ha4Dr9TN6TZMtLNNt7+OfJdNSRvfgosAT2vLJfafglEs
FWMZGC7lE3NPaJ2TeIij7g0nMEy7eFkTctlgO6gCsfQNyyOYB+jHhY9S4twAVcpI
JxU2YCcg5ORASYBB0lc1NT+PTKv6h2F54ToBSpuvHDuvs5swYcaxdXYazu/jO5rS
eklY9wRjAcKdPRxussda5xoOjwcgdzBNSETsCHPADXJcZqIbJw+SDmH3we6FvEh6
hV+wFZUisYzqSUIQVFrXwLs6cg8Vx0rEyiYfcj/Gbhy/wD35p6Wq8uOZIBuzEdgU
5G6hxMYxkHkTUojaCdydBT95mar/EcQ4k+xuad2rGJVGulay2YsETmKof1NCBgV+
a/jPNog3q+XLXe/7boRPWl1zOeJRwrmMsWyyBwdaXIiz6+cKZzIdFHBTGj1tg9GV
lhVSm4FBPSmlRJuwjZLwTO5vUlhhyIDd9ILJX+3sC+4Y3PHhRQqBDrh2BfgVMBEI
GxhHkuz3Hete4hjE/iP3AMCqGm0l8H/sgcNqJ592THtnkjc/OwQrNc0Hit5fUCLP
I9C3UQHGiwpMdcnccsisKZI4HU1YE39I70JRcZpaYBE9a+oIrU2ShAblklgOlBMb
gysjO4Jngzvxbn6vc45Dn8pHOUQSsAamwwHTsH8ihek=
`protect END_PROTECTED
