`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPfCTh562KVLp9g+GCqIoJdkEf5R3nxgwKjpzHm3hFq2XDTQ+D5U1TTH2ZemSuZY
dBU81Um3svp/UKis8WlcpiANZJAbkLqfAGoV/t2UklBeWBRg5zZ9BkoGby3pTAnZ
dJGB8TcZwmSWUvM4ztFGr467fbYSyP08RfH9lzzOkldJRqrCednqoPLQox3Xg1cE
tdvOZYNIvG2/Yi36e641Ep2PloRbgZ35GZqSlq3zCg3uifLHvzFcdte1nfFKnZZf
5xNhErwFd8YcrCcaTadEQ5kFdjFxxRMaCDX/OWjc8vmghMWbp1DxFpJYw/UAVOJ7
w0YCICVT4NPPIO5kJKdJ3Nk8B9h2qj4Q6DSQSAYEDMpBPKRMsFgGcTgzSQcQymm+
17j4+BCwHFcaX3oUbcyv5QFgdmvqOitqvjWqZTtGcwk9l3YF+WIDO5fuj2Dw4Dlc
zpJKpt51JK4l8OwZMZESY6COUHzURC3UWJurt/Egq0BStpYc49g4pY6rmM4cm8Eq
iwixr32YhryOjuNcviB0J5AhDk1TPeVoGXTmRCvfcESPDHhUxIs5wslr0fCpeeX2
s9xA5GfEFzRv0DZeeZz06LFHDrupZ45/PB40n9CncIKrej042R1qnhzK+ws/LwKK
0+gx17Ycak4gtqJigRgHUJ86xOQt0L+3wN4Xpl6KVSyfxSQhZ3x9svY9Ciunvs8t
b6PPTsNUPwvpfCeI8DqVQo5xl9kBKp8je/GTMBWMBTJljyZyouwcC1UsZHwSn6g5
LEd9PmeSquuEpRasiE843jy9zV5tBj40VXbim634SIQmVyle29WDoOsuMQbw/39e
b7eURSB84o7Lo74TLH3Ni85YRFTDQhF0Otw6cYPmWITnu+jbgdh1n2W84UlDejPB
KmJodg5Kyo2Eicdx+KffObkvUWbCr3XHiCdSq8qwIcfRmxMgzpkrkBY1lN//XvCL
+hKJ3Y9MO42vjaayfPV2Bi5QwlIvj6yiv+eftBXMpu1KovGB+Un+ST/40TwBZ1vS
/dUxBMUkoAvqBdrDZLQh/ObTYNNESnN7JhWKG1l/Nw23ZRGuN9UPjy/iuYvZjHK4
3K79VA6+HowK1CQFZm4W2uS/uy8Iq6HH0w1bf94VY5/oqnclOFyFEGbqk28RHu9u
8Ql0taXGbtg+qK3K+h+rzpme2dQIaMgjENBSH7grceY/ZYb4U3vqdP59RSTdxufZ
8PTMAYBhSh/T6XopOHOjSQklzagBJzo44AJVt3CVNfrY5xfJ+/i2dlpvUIPWSysi
Z7qBqD0MKvKRuOmAQlpVFjC7QdPWt19heWTeiNsPmZXt+LkJ/rhB6ulMnx+TCmzm
js9HJ58hjBePk+ft1XQkAFFm/b8ltAjSGG2aTwaGR/g=
`protect END_PROTECTED
