`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/scIEfNzt6kt17VkDTJwkrdbMSn1jwc57F9Glc55HSTszSXl1DfvuujmPiRpEBRP
IgirvuYA8WMSNH5jlOtO8nCPPidtCCEcFDxFoWmTPFTXGsby9FS3cgBIil2HwhkH
orhZHhpDqo25uFanIb+TVyV5EiBUYHc3FRtcvzsio0UpfKzQzyMnNjLv5SGgx7ZG
jm2lq8Chqroa3eRVWgxBTvmgLsSi4X8iTC5x6jYUKZpz+rwPNii80xzA4XP7uJu4
vB2ze2yo3H58YhN/IPafEG4RdeECf/VwCViw+IMGYrlniWIkbtfq6MEauaVv5ju8
yQX250F2Rza4Np7gZkdDZI/fxpNvy9qlcOi1tlEb9C1+NUu74UJ0hoPY2Sg3cIgF
Gd3fIkoHNTBcbfIrh9lRAKdOsQvz4Nuqa7qglRHdhsHzVbb08kPkX/Ub7humjdyy
A5DPj4UpvtLvNfkHUqFZcm0j2eCjKZq33IYuZXvocOSmmqi19IWpEIvdlNo7tW08
B4BojTsJWZJYno8EsijyaB6kEOoL3NvL6xzRXghay253SRlY9HPIoirJCjxPFta6
8QXlLAhLu48pnxl7rGBHOAP9DofiMRFoBr5MgrSfAvPB9pk/3+SkvufWauQgdDw/
O+ifIkZ1MIk2oBlykF3AQRYZJ5Npx77G0ZdI1GCejzlSmxLl4mGEzHHTjSaYHgfs
XJW2jNrZJe8kne3Do+qlLZm4xI/j83fLhxJcpFH8xEr7RQWdfJMAynoRkVUSLd35
Ua6pK6PaObl73Aobkq3qt8CGP/mJY/gPOj1MT8kPPBWmYx9lLY15xkAsuCfqMqOy
dqElgHh+RnDhjXEBctXkvG3iKeIgQGiqgQ4/HfuREv+oD9hIWqjAXMWByGsaDVIw
ppSE4vZwSiGdILKVnpnRdrGwfTpTxTaidcKsgmahswxH305PHE5VlyzaK+BK+PMy
2jPxwIm1eRsSGQHq134Mx7s/G7tiJEprKeHECphmMEZtRLQdOCyeoleJwiOFCzyI
JSVYJy9mqPSiUNUvtywTF8L2c59w3++RwmkY8FzTZSoWcu6c3yG/nvxPNbbYRoyb
kYhBYhFlxt1ABuCtYR4VAYLzoYKGLTBU20kPC4JEetD8gS5A74YAjEnw1pOa2Qi5
8gY7xOb0I6lz0RxWacYrZhQMc/QuUN+OwoTF8LH9C9ntCoKaDuzHOxp+BQbWWvGu
qwg9qGeKxHnqRmT8PQBtUj/g/w/LfMkFMF6cxE97ITkYt2g6Qhk1404FXoh1nr1F
eoL1FPKIqxpLaDfQm8FkzWJwgLCrqzNjAiHwL5H9uhOeNFUmr3OEOBLPXscXw7O9
iFxw17UowrulfeWaWvq9NzYXw0+INHGaBQltT35UPQH9ucMG6gF5A9pCpMIEeP+o
jN+bv8POS0H1wufU9b/IdvCEykMjCqc8mWQ1wE0v2zlwl9/oQd4GfwYwjufdxtP8
M1jg9jBVdK7yTzltyUMQ5G64bPGyU1QJ8hYRLCu27Cuh1gMkpWqSm6WFxTVWbTFX
oyP5kYUex31+MzTGkx5iWguXhG6jLy4rvTQ7qVqcMLEshsHaBWebg8cF7mEKYCIo
+ZtIqiro0hdJb4kx93Pvca55NAgykSdLXOJ92ZwTihtsRUDZUiN8Vz6KcBsncuYQ
dxeZZPXUpmKXtS7JVRAc8OtMqBafokesvo1vI4bJURSOrlutvBaBYTnLgE5qGYiF
oXI8ZEIFIrN6VenhMZnjASADTJJVK4pfIUzmPKlbObQeQ8nBMECkWlDnnix6PONc
VcThqJYtEzz7Gvqbppn9jVfIZlVl8RrPIWfxTevCNndXEfkgQNjJPzTzz0RTtuYL
Nnj+Cqd4mWROMRNvIDgTbDb07/SJ/VgHo5o+tThOTLtyFUR0dedHW/C3+gQv2ZJu
PiANDCiqxebMTkp2J0agrPvx0a3eS/ww0Jn+/PbP6OxMgsdteLneWJLGhlyX+lWl
JB8EBu7bVQGO8+40nEYCQEM5zzX05sNb0og44sNHNKmIv3bCWITujQKBb4/LE0f9
oTDf3tT6LRI2zUATAxIV7847OpCdCPZ20/s7DuaLOaO3E78RwQpMhgwjupK5zy5d
L1U5aiv2Bxm2YXXH/SyeJ1T2fpaoIHkHUGDWvIN//B6DCMPpfuZp172WYcECErqv
juZx8fk6kxIquPfWrOa81an2seQHSoomP4kXHhbWcuXb02/f67d9ONfOG9mXAbXP
aHZ2OaEml28fq+xlS7Uw6kNlSRb5xtoRQeRN6fy5Lr7QLLI6zznjnTeScEO5DND/
e0iYezErm8qcEcm4LvF0AKjr3FeBMGr4P2wCR9gYV+UFU/F9tM6tJ3mCNjEblWJ6
QCxM62TU7vMYt+kNtZ/IubAofVxo1zwoNtMt0eTekRGNvhTZBExW5odW5h2XAddy
OIAI7B+QJLDTBfvQ3RO7q6bHjC5wXt1ZfRLeSEMztFlyOUJk1NYi8/2xXjxj6wSe
cXa9xBWXfAGdxpi9m/GcxK8JPCZkbSiEfy2dq/NhYZYJdzw+UmkbrBxF1h5OUBll
+EHh6To6N84JPZTtuFFGu7XYgdUrO8RrN6u7617Z8aXEFupHpDuP74GY2pMOX2kR
7pfwwv60zk7HeID3nZZOhSGKmdnS1ebDh7/kzmfhNFVS8/SOqappQAB1elxNoqil
1NIcjcPLlq1X+WUJYUY12sogQ0tywivUtCaleDzYCVBXVhS4KNG2IaIOxPzo22MC
vhLRbZVj+1F1lrfA46alBlEloLfjzJmSIwhJeXLlincTlxlWH4BCTM9CJf6CqOIC
7rIL0NgfDxjQE7cwGQGdYsQYJnrbja9bq6ZOWCANFuh2jjLuCzZbFTPG1bphk5ks
EHBJcnnxH+wLB0Ffmn9/zrFCkUAmBB9mJxPApJbUCnkPthsZYy6/gLelcvv10Ob/
jQIaDEdq6LD86rejF7VgaDR/ZNp6yVRCNsDQt5S1rPMz/IgnG9NTfhG3cxgIm7CV
mRg7CHRrelpXGk+NQ7zuknwHhJ7C/lnr+7RVjHhp9KBJCbvLHRO2jr4dujGpvaST
W/mPOCqBqAdrxTDo6LwoPKzg1KBI7AAxbbyRJeLQTOeiSXwbWIvJynpGZx3Xdat5
14qQY8cZhZ0gXBTWFeCyFYanfASuzRSu9C7B1YvMHpzSl1PYpq1gyuR8EeqfuZHk
TReCLc5U2/4T80ZQWkVqTvmmHCcOQIvA08N5UmjkjWJS4hMIzIddj23FVQ+iuYXm
lrruVzdv93MLxZBYkCNK3gbDvbbGgKHoxfBiHgtAE/ida3v9GgvS3wt+5QMb4u7B
VvRQ2I6S3Yp1FZTQgaSErAa1szyCqK06M9Q8ozCnydFTrmIKWDzwORw+agHGfFTb
4dolQBaiwXZQNw6wORZxVrbsEXDOSTsgD9uDFq+v+IZuZKAEMp2uju/vHU3XHdUn
8hGD/ryVxxo7kkvGuYrKJad3J8oa7RCvLToxdlUN9CkVg10NDx3bs0f5VzCEmRyx
BEtVdBEYhfGRzs24iaHFLePXQaRGyCjuWfnVdaXHtPQ3zUmX8G3s/i1YBGWURhy2
opGA3v57Yp32x0UCANJOFMdkvn1yH9/Fto1uaWEz2xNGxNETd6jKAkLd6FAkIUuo
C7bmxGt/XVJSEEyIbYYZOtpBezRKOJr2xxbNOLf9oNfM07O2CicalNGYZiWVFvlT
ZVkUv8t+Rwx6vncVgos6S48K4wsvxNoUxoTY0Ft0UPzp6+2XI33Pb+Rc/7/l7Fkn
IWGgfV0lwZLE2XyKJIexPbMC6PT10wZhTZagErvyzvskAiGwbAYUBQZ8w8a+7F9N
cMtV1SHdiTk+fL+M7HElvKcGN/ViO4UMaxOFRMDITJRxCUnlayYFwYwESD1FhfGq
uLioJ3Q3xk4ITV6sL15vLO0nq3MgocdsesUbcMwFHydd7y0jDpqsjEB3sRCe6B0r
JFHAV3PkkqltnhgYRVYPZZ9djWYaHa+XgJLGOpogXWcFrde6ntqY/Jw+dxOx+3xA
rrBIGncd8o4/ZCEEcBWpyrkQ7VyNiWHBw8MwFChlSYfKCw7hCOABrNyZM0TRDjd4
jdcgfCeLQgYJQkVXE85G724ISUBjFRdnfcFMWCL+EjeQCJ+5pkkBWw/q8nIDXYCX
vPOTjz3mkc7Cg3zZnZi4FHUJUCBxHyD6VWFap05fVxfl8u+rHlU1DHQJU+iwztF/
s81ICe32jI6DOpGHVM+ba7/EHMDBsHupTTtercKryXobL3oiUvMAuatFe8KFwpl+
IKNEI1fJsbLxw+AYQDvfTe0LfKMdh+i5lBpgI1FRsRq1AohRdw4vgqbWUMZdPpgj
eI8VD0HeEoJihTTZ4+T7h7VAkltUmJzWMbfRI8RuJtdHmMM3cmK9VlOOTxqLbS8z
CVqrsJ9XJKLmgE6L2eHUTPWI3TMcKDofQxoW6ecZZQeA4M1r2PQZLMfqtsSD356B
ImNk5W/oGtZgCMALeJkTffmAXF4GwRBShYxXcffPgIJ1AniaqViimxl5mrttc4Gu
YrleftSsts5AetGxiXkJtOlsAP4S7odKMpP/oqK9L4EaYWmXcuBzrardQ75mCB2o
ia07Vz88bWtH48gUOfidXG73Kgw7Wn1b1rMKZAhX9qX3Y94sq8xpUJZzhxgb7QUO
UFw/EKstHb3Z82DayYT00U3VhXBmbLN32apK9jfUeUHB2Lqr9DiOlHOzq9VQ7Gw0
djIpNlkRUrj/+TvUPVmCW4yfJwkZwL7/uUk4NxHtPJrbXdxH3XLLD1RlpS7q0iyv
m48Gt6iEpxlN5VHVpvCcFGBcGvT413Pu8nvYwxbbDxxW+3ruzxN9W6m5KAumjmsa
BIGtEXjTtcOvTH97nN7hkcRr3QTvJdnoOmQiZmWtwNpQftBBcJH4A3pLavZx3a4p
aqUTn3/h4dLqkCMXNft+YcjWVdsIp5OWd11n43xU+ad9DAZAj3KuF3Dg3iVCXDoI
lbXYgxO5WDvXm2EEtJUczdBlg7cktXMi8zoNft2TH7a/0+3VmOomHWAJBIrmtj3d
Zp/igM1YssCxaqdFd1xXzPOI+TLX3zLL53vW0vWSPeMJ3jipFPnYINSjr71z+2G6
WWTk4/Cc4vMdtfmeQeDpXpYQiOcmABYq8o48pnYIXPBZ0AkdPglb2tGvBD0TUAvN
HzCyx4r/mnxQOJzsOnS3ruQS296RJQS9gC1wdMjvYj3lvOJzWm10zffheenkMcgL
HVXgOHD2o0ocibp3b2rNeeTpVYSU/2jabg0/vjiw22CkWgPsdfRoX/fLkFxI6C5o
CxN0s+4DFojsTiLZNawJQG1/jM/Dv09WTOLQH/W3YampXOIFRD9NpmpyfpQLoKek
Gr/QPTDxGjItps/CNtZo0l/SBxxhHCSOX/Et93bLs8ue/5ez/mI8//xFnJSp0chN
ApgvMeERy7lXxPv5hLJEW1A1SybNadCJ8mVWBuBcfTTbSe9SxmrGkUvFPBTlTrJr
iUkSqm1hzUWZzU2D7jFa6aK/hA9LWXRJRp+uUCoxuAPK7KH8nD+7WsVQnRsdY41c
lAu8l3qEggTUXx2gznUdY0xKiR1ewyiVPcKzhhpNJmSGhwJ5DrnwuGj/i6I9ZhZk
dLT0vkxFF/3BlZRPoSAGtbPhoO3n9pc+RvlE7GWMqt0/KNHDwBDSQ0KIuiWURbzO
Ccy8wuaaeGrGSEz98t34R0PA9F1F8wcjGh3/Nbv98f8QGI6vJ4XyQfpllTtxpEJv
rRQdYfffQn6zc/rdl61hfXjoFh2gOuJMO7pFHgx96smI183tRYgBXLUsNN7E+JWT
VzVNYWh0bFQa12MStaBQlRTclohN4duGhvu+2i92YC/iiZu0QVllyFTU+EBSQ8in
s9eafAxO2e7NBI23ru6MsdsjQTyHoVHG6BRk2ZJOE2hi5//m0ruzizr5JnblWQrV
RPzc71/OKvHGMjfqSWYYVL+xv3CCffG6Ftn/mQOYnPU/rj1y0tJinjMEp8M7LasZ
+IwiVvffggkImK54EgG9Yi3sJYMVOAsKMQE6B6Cl4v7ujY4avhzulXzWGhT+M8UU
h7VDGfJRlWnjC9hVRgIqYFcv0slzwZ41eSTRPhncm1uJl3FywL3sNY3r03u4+xnP
6BXN3rgMuoyQv8pbl52zorlsZRJfXy0tupr8uZOHSEMybYpTTsWYGD7UzjvMa1eZ
DND7Ig+ppNilK+mWs/6HvxQoTQIzgbpxpRgtzi/xUDxXEehDbqDetRUGNOKPNnP3
Mor1A3yZk4RJrPwkgZRjPX4QFrCQdvAOXeTbE8jpjfRuKATPWcJ/jKwxU4Grm6CI
yRb8dVhulC9b1iCQ7rictjRfuXYEeL5xBjPnqukVxeOzvbuFLM6iW7KqJ8d3Ll14
ptJ1lAUx8xxoKpbiTBu8zDmE/f9sGRMymwW/gslFaHq7ub8DO3imzk+K9EM7kEz6
eIIzAnH2Ev361+TTYBhj0hbjnTipY6FjBwqAie/7HIRG812sU5/NQp+gexWUe1Qr
Ev7/Ue6Kg43zU+Eo6kL8VPXcs0gEGFMR1PGrrnO5VH5KWF+XwIAe8dgyzWshdfMm
Pkku6+hxafS5Jd0PP0l6QUY8eX25Wv/n0/ZR2u9wQTaIw9OM7Z7qG7ZtAewNWeHC
Uh7eQIe0DT1IlxZnCGG3sGmSxXVSdE2gSPnaKrzd6YYehody5mMuiryvwvUgc2ad
uSyoz/tSRjerLzWnF9iykxusZczu8i2r2v0TwtP/eKYogY6mYGMXj7/e44ee3RJp
Vd+PG6ynhRZrxY/c2niFrXHe/JpU5WsBTlElmBsTFFbwfZSRk55pBE/FJdKj0GLX
XaguP11uliIojf6Ym2rCM3G6TOIpvYqG5Gcv1iHJFmHWb1fLwmknM8FXy3dsZf9x
ZyzzmJ41rJmTzcu3TbIQqrUeZ+YSsSZuA5XcJ1VsgzXLlBIESk2srlqRScSCABDO
QLQSKbbeDi+CrwHAHg+9VDDfpOOqqoEGu4i7xDBvor+9TNsp6kMkKwjeFVCYWBhW
8V0JCJ4IewGl4OWRj2pQbXYEARQKqsSOvfKqj1IBBMlpD7HE+5j74sFcXy/znew5
KkWvY4HAo+mxYTJT5Sw5iwOihyKUvNxsoNiFDYHEVxXkreINO+97dkBDXtqOvnZJ
cVLNspbUjkLihUhjsEnCAZjQkuozATYPHJlQQ+dsjhTzDtrBOlD/KKbgSk5Fhpub
fPJEqKUf7G626BioOBtW3nWWNo4j6BEvYdaIf+AyYYQnRTuZUh+1ccqXiyw0lbfs
36HLDOd5/HQp8miN5s5UFhGHH+W0TUw+fOZksVQOOD5jqTs6cKy6q3iu4PcYXmV3
v9vqASDi/xwqN1vqO0JrphUHB+UPxeisVFrNTQc1WnHVePcgzwVniWZItqJ5BBfp
sgAsU0+YY2LSH5OhRWAVOca2y1MTUeXGzQpTTQV/aRjhMUA5GCHzjbUoTCK7Zaii
T/MqANepxorf4MD6JwETOYHAoA2wDWCjDegIJAX7D8HUZdPgZTl0ThYKBerwfzgh
wd2OCYkxVWGLxEyO0VdlIHhDzsG6O0d7mlll7st1UXFv910YfRdoWrGyx+WcRJP8
3HBatswal3Wa7WVW2Ybw7gEdOIhJELrCW7Be5y1nQr/xY2r0WcrSbruacaEKtzcF
3SaXllvQwGdh9cAyLJZhnQQUKj8L/PJWCfAruB6IX78kt+vScFTTEkbZ7s9AzmsC
wwaGbpQzvbG1xHYOShHqSIDBGm6LnEdzhC1WLSzubo0kFxYpDIPnlcJ7f99HApmw
A5eY/ZGGNyRGfU8sfWfmLRbVKNV1pxTX60EPLEFr9Yk/3n4xTgHKXBNfTRefS5aj
aRMYpeFgoFeEFR2XS3pwYAgoj6NhJU22gK1sOdDK1gDL0UP/FtTk23paoBYAZeJ9
fdi5K3Rkq3Ex3m+a+E4rrgDe80woFKFuwukak4UJQBkRBRFfOD5aD1YLBi+13rXS
CuWO18YL/k9Xj10kMwXafiAiUOibiQqrOYrNYbC8qkuVlB1/ImPt5VbqIB5CIaX5
WkIjW0Kth6RejetkX76Ar+9FSmFkJyaVU9U4Eb69CM3vXbX9Bopp1axuAEAuNu4I
tqnZfganjzbQmHCmpMzkNgqAjROrvW9hymhlstD6YeqpBahyV/9qSqxz2shTp1Vm
p1wOAlqdsBO64YTjNHUJJ8OaGcXW9qXPGIoeSNRQAS/wbwjyaNDdaqd85PPs81SW
SwQhyEoNc9Lp3xu3cIK3DKXB/aTUIazyldH/X4cwcHcYVJGPSFtxw+gt9DEwPF9K
BCZw8GVFLNk4V0J+7pUFw1wIa6xAn7q4pHyF2JR1a9QOKYpq0QmxMygT0lCf2K35
7bH+CuP2I/1gwKK2gan0+v0kY6ia+iyAZW0hgyBL/GCTaompSPacpbOfdjk6tZzu
MIyY6rYNexn/IK3mHzBqgJhin0Q5m4O+iXIg1Xiv8Yud3ay3a2AyqkpzCrasJXOc
gIF5eQb0sVACRhGlt3G30piFw0Ii6uIIfY1gNmMTj0IGqD6BCBGSLVEdYc8x5hEN
g6h2lHSUSwnKlIwuIBDDmuI8yY1PK1wGCiOMNSPFbme14c0lYD8oVWPTzVqCkjES
pszH1pd+NzLcGfOhMZIWnYPD6GbHihgtLg4071MUbhyONqO+CnIOfPpukJp817QV
MZnlM8+CbV/aC8d08WLQPOnXrKc266rp/XjUn4zdTIwb0FksZcqRbbARjG1WRhfO
XFCs0y4pA514GZZJLdmGLw==
`protect END_PROTECTED
