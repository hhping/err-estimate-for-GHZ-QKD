`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/d6MgzQuwR77xy+B//K/WYx1heUCy5+T4Y0aZOzVHzDXJPJfleF5mHaU/opkIk/u
hXBbR8YqI+oI8/LmEH5n7VJCaWa3Ve2c7i1lPoL2/IjFWdUGVK5CLRjGi13Ig7QT
I52C6JZadW2UgqaGyyEljUNqGsgbjcKG6EfogVRkftvBo/IWLPKAmiuSkDnkde92
C63tnnR8VwxWqbnd/O8OESTeHSR6u1DlJoMPqRqMDt4xA2QdaSfuz1Yh3c+iB8SX
FqWXcdTZlerp7nZ0G+yEuj8dHGAXXAdomxhZXLOfRArXm9z03DTfKFq/kPUBPd02
zrOvYf0TR4ZTFLMagP+qQMtJtlTLBL9LNCDkbQ+cDREoi4OkZ6tddTF8rqtK42vS
0dLXom5MbRH5SCpf222DbklMU7Txam1214pELCl2RiI+0Q3mgmtvNpY1vdENUqK6
opFpa623ALnKf6V1raieCbXJnwc84MDQcIq2RfcQfOEXJN1SUSRFCO94xOw8wmc3
MqQHCMqqwxXLQ1V5K8/oAfaqugwc4FH4zCN5S6j9SVYFmyOH7EmYBUV5pmI01GJN
qp62LHsKKPFfy4WJ1NehSYKjymOYagMxuypy7uFoQiAzxcAuxNfgastP0BlmKF/s
yh9lreZ2FGW1r4V9QbG/jp6lyN5pntbHtaNgaYZYHuo5gfKa6iMfryqLpAtkOLvf
+4BKaiUXvxHalIv/Up3dbh6QBhfZIrjgAvrtTNYnqs67d+hrl6xcMQEb0XGQnJdc
Zc5fA08yFDmtLWV2z//m26/VwompNVswXlQc4J9TDyWyO7XjH7ANpiPSvvTEIA9G
q89k31CJbW8SGonRUm9woP8Ejq2YS8xYLt69z7ENoJQ=
`protect END_PROTECTED
