`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSh1qd2Mx1uR8OZVgTzsUhz0ZINSGW3rL+9Is/OvDSekHmFQ2ZJ9C/wIQzMGXuBj
NbLb0JnJLNYRMMwAsI0o65oYtPZN6R2syg1kYqFxwSOVa9gVjKdDvKNYNprspaQc
9gdo1kg+Aq9j9N60aZJFMF1Ivk3wBwouXtqxapwlewVPCq3lzmp362IMP6SBZZXe
qeU0n4ivLTybcNv4qAfoiOVTNuuTOwOJCUUQjOkkYIoFMnqdMNA2lvg2PBsJZ2RS
K/QO4rwpdPt7dF5/y0ojmlRTO4Jr2bZmHLOVzNhDr5g+UPIm9AoBKsEhwcteJW0c
dmwR4HpLmXxN21Dqd2CAyOc3N1YyFc1J7EAv/iZemS0jIbXCHuvXQK/laEYK60Ej
EtYmHMjcLXRTEFP1U9tF5bpVJqpA7FQMywTlCRZnL7x7poIlrRdRzswCn0L5tlq1
cTCkyYwovBLbAsU1rAIfK3aOZ97TjQ+atYI92cWWpn8crVwIBxEZ30lpv5jYbxkW
1I3qj1KBY6DAbtOZA20rP5VpM8KwMDyC5rctnXpSkaXr3Hhts7FhyADxjdXCoGDj
onwDas4rsh6OUwnT1jbeMmw300Nl+Fss9UXUDCaUJ8qKjGagznP0D2zk/8aga9+9
iGKOl/+ILmScc//zxphijPyN0w9WNv0OJvcgSqi60cJlRJcxRaQ4U4Ho52QPQICv
kZru2yp4SdzUUVTMuY+yURt+hfhfO6JOq1eH9bu3obd7efr3Sys2ugDOsuIe9xpp
heIhw+jxbBlBxxFYp6DjKCNCD2AE31Ra6ciPGMcSskVHnQXY+4KXpDkeDGeTqwAQ
imbUKl5qG72aWMNPncvghUDq5b9Km44xEybH8nQd+8WypllqXgHZS7xBmN/fsAwW
aANUYH4cWE+dLYPpafLbWmvii0hPYzfH/+yyJFfaDRINVz7szkCqIMtUoRQtpNAr
29MSz3x99DGzivL/FkclUg2cR7PBB86FrDGz3I/ht9qOZg5EIAYSNj8qODG9wIF5
rVqJAo3YJjWX4vy1ZKE3amQM9H7O3WIMYoSG9smZydGImr5b+gyzcoL+ZBjBoihF
Du1fXkHtDT/PrvkiAiYDQD3tOgp1DOB+SY7AnDQV+Phm7ttGVn5UBEsD1HHz6kwd
uGCJQ08Cfy5Lgn2oPpmWDelbt0yeJkS3pwMBqISTDUTmlk0bSfoUaoD7erZMeHWr
4CSOp11IqSKYoagxrq4nB81iFh+CUh8rixYS+n102MzGsYdWUAv1SklHmfJO7/D7
TTtSAU55Drg8CzBIPwsM0g==
`protect END_PROTECTED
