`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMthElPsUXTCNvja8OlYGCti9sjrbIoq2B+LR7plU2Zeb6AWWTQUcD+61dgFkZiy
QnpDa5V7masKdNs+8rWhPJwm+2DrD0Epbvlu9GvK/+sCGNS4VZFqEUz2fBQ6gST1
pzkv4eV6UX5tbYn34Jyb7HhzOVVnBcOSN2OjMu67kAjyzRU17Q54KzDy6WiUhil+
wx52ktjPZT78k8TZKfVhYf65WWJkK6xYVm0P3WQgvjHj2AG9GMvDwOzG0PTjIdgw
AYsRaSlERLEXr9HD8sa2jifUkV9AyR9F6FhhREJ6yzCieqgUZ3H4z/qHbxTW9+ze
u395vUVWQHQGDkdTwg1gLfECTq3FeLTSkiXkQ9J2DWADkK+uTc17qug/TNFR57F+
x4FB9XT3LSN6sNxlmSHcjNU73hzZ0q5TLYLwZNLFfMdSjZY2SDBXLNZVqpYWMWc2
YDmLnR41ON8K6c6bMrW22+DOGEOxdYU9B7B61McbOs4QlBdR+TZnqfnwTdOxVurP
mMXgSX3oZRTIpjka5qlhCDNqBNmMxrWR1iAunmcZUbjqwK7FE5rLb1tIhBh6XJuZ
s1Skjul+dXUzywEfB8vhKQ==
`protect END_PROTECTED
