`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3cAThezu1Np43oq+g/AMQzS5gA1sugm/GBB01xPnLux9VJKRVtWYdWvtB7Bjolc
1cggeix/lgCF7caB7hv2FQyETMEu4mpzu/Iz03QMRkmzc83xd6nA4Uidt5Fnl7fj
TA7a3my1kGqJboYLwqzx1bJTmYyisW/rCDMjJ260bSNXCjHMNSznyc8RuSrQdjTW
6oknjFL/gQFzziInngAWcYasuG7SshqLknr4pqrkkoO1JprkDoumvW9B9E+jy3rP
Mkoo+CFzky2PulPNIE0uDdk2n0pLZfzqFdDq+NIkj7ThiIjd5Cyr8BOyaYV/Gzhw
1usrmdDZsFaTCdE3NoKdwTOE6hRu348r8y4oF9aHTrhpIa4Z+HKVq1Gsf02qi+fv
lGe8OxYAwGuaMxemgJB6cKhRKo/NxkyOTZnnE2goCeNjoBnPRhi2tiKoXXG40mrM
kpdQt30UmdbUp5EoKYzu+ELqc/uJkPCOImMOI+yb9VShZHkavzx1+At5yH7BcYD0
xhoquo+kJ1rUSMpglp0C0XdKOVMLji7UJYWpaVEhktaSLnCWZzY9doHNGcinsjTn
Fjf9Sm9+BQRra+hIbiHFm/EZjcSiWGxtzHcYjMmkBR/pP5kTjHLo3dWP1c7N4KSy
3btdglsnxF7jtL75EbkHA2Wyz1H68P9Resl2sZzFyOhb+fewxd7LVUnJ8EquGwpn
CE5WaFPbAoeV150coxGPhwnW03XuHZrDf8qhscx8CMoIZBmnQSmY8ombQYHvJujG
dZVoOoSGkPEFkHlUSovVIw==
`protect END_PROTECTED
