`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXNAlCFcznzUIZHPppAsNLhwO5+xods4TwsN4hfXjmG1SASc10yccANiihHvT+mF
Db3uC6WVab72fEDrH7UacudHWvE+3cmh2GWMpmNa9l1pdYsroSjwqDG2+f0Chw8q
k/TokIusyF6PineRJH6h1DZ6YRZ7DWXzkyvoncup2gGBozQqWoyaEzHKXcXC3i+V
vl5fRCB0Jrq95vOmPH3blELvrh23LMTW0XVFqFk6cTNP9umq6cDvaAVwcJNd8kkm
TkSD8W43ikCT0AppO6Ux0ALzA4ZKZdrtl2ToIOWeRUuG843Bn2dM5jm0cGYv02VA
+OI0HGsVTnVFE+QP1W3vU3a0mEBz5iQxavu/K88MY71eh+aEFBLX6EAYN5WFFIvp
0ErARltDUGpX3pvhacM0K4SmhLBQToFHXVWz0butVUr0Gfg9usxDIOA1ApjrFBpe
BDAJRRUAdq9euk+NI7z0qs6WSW34w9Be+t0xswOtLbyFmZlpuDtEATV1n3AijcQh
g2uJf5Sv5D41YdyzWHfa3nNPXPJKm12Y1tCIcEuk+j4r76cS6xkJHzgZLtuuNoR3
9CcF2BwoKyUJv7JyI1rVQ4AS2Ik0mPdtblivhxLYtqjvhgBdMefztt0ojdrxZ4I5
Tc91jBRpKoHUG9cOE61JHD3eF2Js5mfyOTMO4Hq4zwdkVlRs2CbwP8Sq7/iOQ2/q
y/8anasECa48PtQxzhx6dRwHTSnx94uHMfvie7NlPjJN3WyGOUvo/2Sj20T99PFi
/aqAT3vLiQRN4kbBWK9genETT5sECSBe3gPkQx99i0je57C+xU9JJQi/oiT5jgde
PLOQ4RrqhL/TuQyRugv3L3QzGRWPrTSyyLQlsFACo/QUa9fZYVv7At4MYVHlaU//
6k92jIe6ByXt0OFrblW+CVqdvwLZdgQepaGbxwIgaq4LZCgELpOUU8TKfvVBc771
kG6FHpa//3EOLxF8ZOqOC80NOrHRneA8dh3UQeqpdfMlv6X5xP9HNbRxa/RJkpY8
KD13ycF86xluHU43EC0Av4zBb/j884ckw9cUdMjRyTBragRlxjddg13sslbhKsNb
Hkok7LWTs4b+JgIrN+X9ZsSzPwyO/j4tzm5IVNO3weGNsuAtvg0lIgBgFD84vEq7
051j7n6S6IvnYYhRp4nSd3lCPyv8nmod5ilac6P0kM50fIYJ5HTrVpeStlsFYt0e
fmZxtDdwbVEo9y8S04YOc3igkBCaJkqUULAO2SCa9EFaYGvbKFdgu4ywONalV1cn
BKPndx3JpiAJZK88MEgVVLtIecmmcODiEERZ+WkmqdmUJXLUQS89LJweOn/G63hH
wjxy0l8/K8OtG/TFOefqo7KbpIppBsWilf23ylOIFRWmkufShlGxFE7FNXvMb8pJ
DViMwEhNX+tZL09i1SfMyjEv/ckCJrL/vLS7Zp+oaqRrhqJV8mKbt/pPZ4iuWXXi
eImZAuKmHmHgNQK2jaTOrP964+mrFBXoZI1dxdm6JjKWt3SclI2b94JegxCKu0VL
cd/9fc9zK8fs91nP2pAX0QxrJbjsjO+KDlLQCmWguwqGldZ7ZZ2iGM2WTcyZJkX7
clDsFWUUg7yGFqcJege3Ttb7tbVVUXHjGeEMp8rOyQc=
`protect END_PROTECTED
