`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zau9XE1oEcXCpr++8YJJVIlWhMzW/h5RV+NGMCmwbf5ijH97FdsTf6v2SuglGrs6
nfCFmS+98PlYZLkfo7TrVItRwFXtGF19XV/hMKOtreFngTi5ss0xO57EIhf/wAby
R06j00+7zIc4jkaqa7+Dx+5KwZ8b2Ev2EDjnvnF1Cu6NvzZMII/fYQzABoEzy79Y
965XZKIfrKqpy4Bh+NEwA7epszkS5TLu2TKBm0bvTGXEoJU2wDWF109lxfidbuX/
cYIauvPIoPiTMOnAyarbwCWF1OHKbniupvHz+MmTGNHNRx8k/VV50wO14DGxDOxw
2qGnUqNripbdZEct9kup+qsfTgsZkf45tpw/tBrwdTT5SpmErf542Gdh2B/PTlWJ
P9Ux+nv7pG3cn1UbR7/VEdXkLyfsY89F37f4RZARD9hXLGvRJhFocTEQdvaLi/9e
OvU8wmecr0xTbswSo3xy13Xq79cH+z2/IN/Ai2IxHqh6Mt0uRg6vJMkSfDTXXsrE
soHqIRqf8Q5dSRXVshu2jHxORpBfQY1c/jVILRD3UYE1KabdmfJ+2aIYvsCl7LXe
2yX2LR4Nj1SMEGm9DDunR9kscrFqKyRA0RJKKOXCldqOGl78Co3mbvar3KdaH/Ub
/DVgElmX9+FOajE1QNvUav0AXDNA6n7W2DI1rbdi5YB8Bn0DgEPdxkLQSDrOcQ7v
vRUdRg1cHRsk43F+AQHw+rMIMfAozHwRS1Qvs8FopB77DS1oDa3BqGju70CM4uyh
pGAwYbzeOIMxK0QDDM78zdmzJlme+mNTQ4wG7HSFwHE62rG+X/ld7yWvaUYsQ60P
s0Fpq3gssdlq1tWNbHhLuIa23uJP8NmO/zGbE2AzMZtE034XhgqnqSR+AAl2g4hm
eoqGP0tsZjeYCzyUPuq5h64JhI+UkAg/QF5Hu0Q0nTPtB8lqhWXf49mC9dPpvtu4
/aDIJljjCNjSgN7tQL0MApZAwG1kAZe+vy0WjflKoG/ZPI99RDxL4UTvRQEz5iRE
Mw152gFopvIjZgvnoDLJwEk+lpoNY5ipjPsl8IR3CJr1IJfGOd+kZXtDUBftbd9g
Suk2D/xyot3+inAbHASlb0jXhOe1owaAv7jbmGVuSP9yDovnvCvbdCzjYAHPYNbA
L6sJ5T/8Wai/cmvdDrSrYgPQA6kfN5IjCVUGaLRbIfYBpuvWp+3Ip5RQwP9CWToD
b4LkBU6bsDGfRgVSDD+h9vXqz+Mox8lighQEh9A4pGepNdahFpLw+Jhesvan7q2a
QE32/12Y/XiMjUFfJrCX8kD4jC0rDrHbA4+nqGWuDAN/UrekzQv/uFvi37RzGlJ+
/aESYPy8iDuTXGlYt8F1FfOGCmadzXMmb9xOzlkltMU1xmHEdWMCu3HBBhv6i80t
QUIDG/xZ+peSTaxbfy058mlEY+pOcrbsP8+m1y+fjsIJZvpRI+iVOaVdu/te5usW
1U3WdBnyqcqPbhApeDuCW9hI13tsm16axeVjW4M/npjOm2Jj3zRFyUxbgpHQsEbN
jpOMOgJzgXLJ3+Y6qcBfTaVOQWdLhKvgG0zqcopAxF0KtYZ4sHCZunvYAuw09LGc
YxMyPfe0PcQAGrZH1RHWoQpgvGfDtVcamS9bOyjVsPzRu2seEw9OOH45euHA+tR9
vPxXctx0wxeSeDgtVBV+7y3HRykIkXbw9BveOnP9Rz2ae1FRk5KL15iWyNMzzqN5
/Y1C5X9Sh9r3G3/xPdqrd6XzN6RWb4SRyEbpHv0UK4Zc021Pwuuh5bsO+m8bdYWa
UxqY78e/oQA1vMQZdpNhUMbeBtJFktYKgnUQNLV8Vkmn67Jj3GrzDGTpNWraRBYK
JHlxbXgQO/MC+Pje+XNktaBYWx2BQHyMVOrw6lr41CufWUDxU6P5u0uoHOShrJUw
gfbVFeFkAhNEUuUfHvKbO4v6nqU4LJJfT4LBMy4BQ4tjISswZG0uD6wqFN7XsHor
N7/rK/sbFwMdIBR34gv+mo2eFIuo4KPGG4FG8YKvHjzQszaW1ciZGYY2LC6OxvCg
hMc47rH/W9kMyhZi6q/mzF06KAbrnYpC7qI0qT08Z+TuXQmHfjGxXOdkOnyfwD91
rZM6+No9Yz2Z8jDH4hcOooEVtLO4frhXMkdunPot/x3NfJGDQolSKnNMbhUIRpw2
imMWyqrdCurw8J7b2OuqPsqvT4pHc0N0ePJlcxdtsNEeD9sBTxFd7+oNpTwUo259
Bzbx/5ndj0je3WOYzmajEkyrRFf8GL5pFkB07b6/r3ugx2Q0QeYJICp3BiL2BcQ7
c7pRsnLwoK8OFhw9wTVK+08SKaPOev7H7K2cuB7BiCxIEeabSR9FHu9VYQpqrHoc
rGM1RGDO3vJqhNRMI5ERy8hOxMNypzhN1beoJyDKgPoGip+4lKkMNnpJM1el8bPb
AA9MwNUssIvGUYLWALK1T3QF06ChGFUi5iNN2OY564R4SsRMDIbJkmlR61Fkliz2
6hm7ZxWcO/F8ErhyYLr3xyokBXbSJvDyFsjGWWZIO8PzYI86vxSHP57Bxus5Hrgz
3Q13oOJhEkayM9vxxyYeQXZ6IKKzR+SRnQmbh94Su7Dw5rXMfJmGUcVH87KYwZrj
g+K6Vi7KSILM5nYjj8nHwPlLewINyVzekz/4EAHz6ntgC1/SpL5VLnR2/sde6j5w
FT77Cm27zzyfjRgGWFs1icgk01ieFZyQ96yZb1NgnOOYWx9s/PQuWOMrKglHlLcH
nFGcCYNhhz+flt/7Ra1Wo71rCZv4johFedGF4D0MNTwLYBNlgPnuJvQXHfATusrY
er3gz2/eHGUc8dkJePq6rNlyWWs7uY6FTKNoP3jb5+bg/9md77lXSAUHpxXuT6l1
lp6GbF89ssv7T7hqYNsOOo1SEhkDzQtsgkbu7LCTv9c62TTWxq8NoX6E9LWP26qj
HuhGsmhiZ1pQem8lkrU2CAP1j4hJp0kT0dPMFe0PfNkcD1yxzSZCC96nCDvhm1X5
DIz3Y/bEHVks0h0sZO8Lreg/lq5w6mdqmw9cpSvqqS7PwsUPEbb+mu7vv7lyzIo3
sWPhTct+ENiflf+d4U0OgSOUJwpgwgdgIGVFPw3nGjLjC7vqKcqv3JClh/1rp+bG
LGI3d//3lVNjA1PFijuTPRDhULwUoNFg4JR71Ks5Wc4=
`protect END_PROTECTED
