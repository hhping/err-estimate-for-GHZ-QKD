`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeeqQAmqrVRQHa0iICjn/lpjRrdmBm9oTd+W2b3pqAtEhHOGm55/Utbt8BK2VhYx
MVQhX3zfDEAyG23Z2w2wZSjXBo7TwQFebKOgXcHTZmgJPSwYnqX+tLkpBSjWYVV+
CcQwLCY1h3A2yKGPvoGRoFnUiV8ehf0IfFz9r4t20oR0jADOPWUA0iOSK1zsCWZe
5q1ee0fIYHD3NnforqLsQysTxDvPharpkvDZ8UITkLQgpWgm8knbYuTOLYLAVLFa
ZZztcBNcoLsI/Dtx49VW9D6Rl0mmBy17+jp4fjerdW6v8p/X9oDHdOnfK+bEwJWT
LIXsFRvZPTdlKkXINfhbZ4kEjwYM5dKHsRkbKR2yaL+ZYzwsxN2Ui8HcLnGg2gz3
jA9y5FojNn6HCkSOuZ8lz6zxNWllhOHyue6iaARz6wWEk+VzKhihbRZlt90wRznK
n/BT2MltGx+T68T5fJTj8fIRPse0pAlch7F4nzW9KRLW8GbNRppUO4LMSOS7lSPA
JEBw2o8e1mqhy1I/UKR6lDo6/evinXd08W7FdgYDNV6iYp2gHF/m9Ai6LRVMX02o
3Enfg9t0wFTnYOHUuCpvwLBxIJx7IsAwtrTRG3ndKTpGgDA2ii64PRjx2zWhEE0r
Y/uHNyrWu78KxuK2ax6Zkhh/Ema/UuPGgg/IVciYapl3sS9sD08A+x8XQQiZDLji
`protect END_PROTECTED
