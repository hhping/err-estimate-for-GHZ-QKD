`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sz1xP4biuWpz7nCkfIFIR/xHftv8jEZ3VUSUH+Lg3vCPDiw4qeS35aQVTFEJiM7M
mVJzueB/4vLnUyDUp7JNIbYTTtmXqzczzLDqBdNneFupmTWc1z2aMZBH3vl0nst8
lD1JXVYrWJRAhnI8GXILXey96AoYE+EHAMQujM0M6kwHjFu3eg0PqhN2xlbhL5C7
uTskXfa+CDLDyAk7zoF/P+CHl8oM0d/tUwX+1dhi5A/P/pO3x371a7pcyQrZPWrT
w8CuI+fCa074jguc8CB5+XVg6Wq7h2bisZKOxNTHmLCUyyCQ5g7SHEudbzMkbukz
hDDwbC5iy6i/W7ELKynLaYnGdtjC3jYRZ+1ec0govivinz1fJXhW4TEAJcMsskWs
xXvi6FH1GtTQBydNXggWEb+u2AmCTdm+LtMUc/Gi3Fko9VRuLb4HfVo+fzT2v/Zc
SaMMrmSvVoq54mbJV39hIURQrC0953wiXZHV+kQ+ig4a38V/RjPjL9Ky6dXHs7cP
+GO9OqCJ/IWdJ7J7ZXeeiHtA+nRH1pZLL6jHqj322wTtfZ9IgAObfBAviiSPZcZP
49a1Ex/g6rKd2MO10+gaZuXbJmrMCM1Hj3tlTL23kBi10OJ6DXT0k9SDm9fJDJfv
TeeXgwGsYpzb1e+csWd1JuHS9mW/bfv4Z/kzVTQYAuJuhdJpZVTVOIJBoCWwneLo
KoVDDuTUq+8+0qXaRk+Cv8F0DG07bHkvG+yx4mgCaCc=
`protect END_PROTECTED
