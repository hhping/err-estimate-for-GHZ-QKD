`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3WKxZWqQeKgao/TeeY/HluIwI1kgDLK5RnAuXTPQ/niviGvvlCVfIv8ueicUVDO
nU3iSkkESheh9jG4UNFP9fhUKBslOygOMTqIyWGd7wHJm2/rTzxIMOPWipw3VClE
65LcZbqScvXKLir8HI8pHgklAx7KwYM+PuXZLVgIh1VbrPX18VC2TluusHy62GCy
SWXVOEH5Cn1iHQP4OI2+w1nUdo+54k3PcVp+9HN0NTPj6tufHrjJ4vNZ9COvJTDI
MC2XZgElicQgUP8tsKsYOa7YOZP6ZHEFUzEaZX9EwxO2lgh3zKHdBBBuTP4PRaev
U25CU3cIohfExpyolGpV0SIDyexQyu8/19gdVc7JBCA3Gu61oYBNpuWe/wnv8+ke
9XkQVTSAgasbAmxouJJ18VTgrdt1CbC77NLV95sgl/0emFsjIHDZxvuZjEbrGEtP
sZ48NUF3Ip3RrahnH/pSWwYTdRYdwL2dtmjxpuxQX0SF0+G3OxV+wZIUZ9V9w4WN
n9uclmP8zYEwXp+fDGMDDN38Ll8yCeOi8z+proCfFQ8BrteCM9TfY/Gab9zNIFbQ
lsRs1WICP6LTb1GdGhYobNMxM30nYlVl3l9mJvpw895eo5ERrpn3cyFJ1usn+aVn
yV09R4S8qrTndcyY+1ExbBHCyfcnmBZ4jiTUZaODvo4yVPgpqR0NxeD8BR3/fl65
ATLcj1l0EHtJBX+jfFS6qdgs6u+h5j3tScGLEA04jdoIp7Ubh8MhzjYODtF54osV
JjxW31n5v8p+GpVoDKUp71sUBglBnzkE+W/MgAzFHlx9k3jNxCJ3KFqw+rwEdabZ
k/8O5jYcNnsn1yCca5iUqCA1sF1vlXcRzYsN1hQHWa2SrmS3QVwdBbu184X6MMk1
mywFWdR7P5zrx/6Qtk8vhae2QKHJ+ZPtY0L1UgKt+MXmSdJ2N/l2pBkuQm3OsFXH
uECNrO8GCqIDNGngsheeCmOFwnYGpvs9jKUFszIbl7hC/9wVZ7Z4GoN2cVtMlQGP
79C9nyg/zc9P0BCA30qUvLCDOtGyNE33jBAxLgsEJVRuaQn2CshQMedCo6iNHwSY
l6vgEbz1x3w12MB43Hean+VIy/k4GACVs8rU2qQ3gc9QxS9HUxCc01DqwznetfAP
P3++GzvIPjZM0RhHEjDy6d+pu4XOVUXSw+qMui/q5c0=
`protect END_PROTECTED
