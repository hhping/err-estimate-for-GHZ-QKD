`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMyQfY4EeV+GwEHCFBgVhNZyQXAO9a5aHHcuD3PakbQnicuVbnIzAUuI818Bi+lr
MOt5qPwDz2/Kk4H14C5LeVEDZZeY4sM18VT6153ODS6oooXPzT8yByURzUAHe3Wo
vRvZ5+avhfN62/3/haeNpa9yUmSaNKrClgStWYaFTT/HX8KcxbtO7wdKJlHuzvci
nGFq71sTgRXuXry5U/TEK4WehXBeP7xEWcV9EhgqIJ4N4K2lfS7zpferUF4ZbpZM
SdJfiQ4gZYwOhuEKyLXlFFaL0itUC4WlVjwNmyWEJUZ/ymEUlnaEwmBev0G83Uji
GkK+lV8xq3PJPRtGp/qjP9jYjl7xoJIbrnNJfg4nn/c26ZBJ981D966vF9DpG31L
ueBwRwm4BpVYZ/YQUroloeKveLRGtdLY3FeQrWwJ2fGgtAJyFfNvKC9eKtiiaRos
ST4cjnszQuGTVah17z7h1Y4S6hIn5lPmaAhJ/TbsGbpmW0WMi34f2+Kh/DfKXiIp
7XdSBVv3QiBYM/JKtQPTww==
`protect END_PROTECTED
