`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKlOEflbPPOP9xYfslmTVsJxye19tmpxhMw0UPY+OaB74ywJsrBmDvgRl5LSt+18
1e1bx48N85k7rdVynFfFSV3Jv5xMmPCCvborqa+5r0dvdOQU/86r2LhuZzzdjd2Z
39g31g93Xev+o9EMABhISYIg4kYGuk2Ozw7L5WvFwE7tRMblh4QJRGHAUctf3S0F
qYg26izg6uF/mC4xs0gpbszrSpcjUrtJBD0pjU5whURBH0f3S8EdQsO2t4SP5Mww
7tS1Xwi+fZQIDSb4Cu9Iq29vdCY/SQEna1b2pKW01+hTeWA33XMA/9AF3uEhsvyu
PSbwRir2vhTzXl1jhDbgt04Jy9ReHZSW907I02D9pmXg2Nl8bZKVQ8399ZQ3E1Jv
LH7DcEY0192VPFG3wQb4z2GkBvH2P8Yy2D5vudy6/jZMv56rBuMiMHc6fVDntGrD
Y0fUaUZv6Zp5Zs/AoMejzjM/Q78XrdNv9UdDhv//lfqTOHKQVzn8yHq5c/giHHrM
yAuDxBfNj9tVcSC/6IRa7wE837826vKY3THQ2jQHDB/RITYj47UqeYDdXsjs6DO3
8ZJVAldJxDNtq0BvTvM1LKfx2ihKKAEvs6wVrz8rI/B4B7Iq9SBP0uD8mr1PxMfs
JK9OCuFlkFn3A0xhdkdZeQGC1zt2SHagNVjlxz+BV9KwuxQau0D0fxrXKVJ4oGNK
c9XASnQkt4ThwBdPW2jyPjp18h1wUwXizHqdJ66KE0hRvSjupUMYTJbEWkT/zLlq
1XG2SQ3rPC5jSkeSDc9xQXdGoF6Ea/yPQHX2C5cKL4IhEd23dgLeIOWejrRbdhyP
Mimy8KXXxFa2VQflEnUET4tR+OmU3fPrR99DKWgxBQD3D+MMmN68GB/oTI2wtLWu
L96Ib25XY2TxKSdDiw0H41adBypiB7UJ6zSWrjH9VlO0MPfrGZ9TdDvJgM1luq2S
iWgh0Ib26zRJQ3cZhRt1LUZgeLsiS8ve7v+V/xqaf5oXFUzf/pjqOVmUmR7OFgYb
SSfTfjDWUZ34J6eiTnQku2Ik/xLoQ+PwKWB8va+VaWA=
`protect END_PROTECTED
