`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KycPjLKHhGiK4qUsPSLRkj6ESq6sz+ybhZFIzzlmOXMUpZ0Qp2cqi1kVxNkVTUK2
sSMCB9oeaqp2hWl10EhUOkcCqsigU3sqJ2G8HezA6Gj4Y2YrlVgRzJQ18fE6H2DU
SyEqHwSLm6gOax5pnOfUBamEDI48pFjt+FpyQAXAHI/YNe/O8EjEC4Yx/Gb5e7DX
xCREt5mmdOJo/aZLWe3usxOEdR7uGB2wpBasr/Ls1DwSs6diRUS+IfCl8maEbxj0
XjAbHmCz34DOsfAaqW8LB2Jq/FIqYOzZ0CEH9GTPGOl5bj43k/k4lx5rB14SB3x5
2GgSh0VZZ0BoSB1vxKQ2HApRohMSTlpXg/BxdMfOOMygvrCuX2VbGF3IQMK89Twh
7mjLt2S+faA2YX0wyb8fUBZ+VTE2oi0uAWgiJ6cKT10xdF26lN0cjLaTNM0Jcber
IHYxRGGe6zNVj33EOI8UnO9cGL0uowqGdTMVpBw12PElDwRrEowzz+448LAeYww4
+nvEJ7qvNTXNuEM3AhTPNOVlo/tK6vAjlXLC1vN196IUuYFcQMocEIpj8e7Bqms0
16eK/nBm6uApV17SbKwmdNTDtlDReRNAY5XvnHH7DW4cM+9SDe65MG4U/utmRSlo
5h//Y/YrEW7fTZLKBolWW538P1ZstbQVjePQAXGdK9cHeXahsNZByUJGykLUDCIj
0nePvIZvMN0hdL17Ghk2SqU0y98RPqFRDsXm5A7G3UB+gHie9yCIoTWdXT8xC/jy
jArzLDe4/aruVS/ikxbsDDx+IFeeNzK4FBI2ZFtzaLUhgdvaQCaY9CpF9TREJA8w
d6+QkYfqqEzmZknl9f0SBQ+0vLzboQftKPcCE5VZSqCcKRoW5YOVr/u6NvM+YMfm
aTT/M0rLMaqHB9W0nZ1XPHGykegrMhwTaVyKuU8jya82tk26CFfmUt8Gv9E67NZY
06G1VkqshGJiekwQCGAksxBZae5ELRlRJuwcPTY3xiVCKyHphsrhfqTgeV3LdPHG
eyoFcxqLg16dRu7GpMxbqYUCkYJSXg/Vcdmk/3UkgVCl8U0zf5hQ4oM4zdN7dFEp
hVWMDdP8Ow4bDhE3w01+Yvbvb5w7QkCrGzkqQhZOyUXPtkAep1ni7fUDpmc/PYri
cL2V5Wk0scHlpLnYQkvfSNY46iN5o0Bd9K8PowEdiv0OsHH5OcgsKdFoYC0u/mt/
eDy9H3YmLKySiCpNzLDtBhxQ1cTMpURES7pi+erkqX81UpXqzBSDnnRj4qAqRdvZ
2WGzR1SYM2FdOxAm2h2OZEsnW0YCBHZ5XCHmCRkKeQ/wIU3g1zi4VwcpLXn27Qi8
qGj/ZMF9riG7TQUZzHE8Cj95psPuYknq3MRS/xBRJKEn3J6YBZJWdRl4DO5igJuz
cvo2c2/RtOpK47KcCI5DUfLDKDE05+OZZ1GnYH8JBUj0wal1O+O6sRHhZEximZ1h
P34kR6TxQZlckbHpZPZFtnhXFXhtDlW08K0JMtM5S3Y8L51hIAQ9TZkmUnr5VCPE
JV244LenfjXSxYAw7PCLwKKJbl4eLc4BRIApVjeXmsnbhLvTfD5qave6QVhisNR/
xTVB3pVMJefaQLGMf6DldZvQ6WZEWIco6tg8r3Y/AH/GHaImC2XL2sxkvrOSLmm6
XwbEIVfBCQ6cNHYKTwmwUQMT0zsDRZrDFIBgeUCE6EifbNrWDuaVuNITRwndnXd1
FKKt1iOluxpvqOMRxod8pNumql/0Dt5k85dSjTXa89qypXpIZdyJyosGdqZMh5Js
imA91hqNYJ1ubw1EfqP6ejIaC0v3Dayyhq+7qwr11OToXr+CLcZtY4QvVihxW38T
v7L0fEQxx0IzfPQrvcJ8wsuu7TmdbPV/zszWYsCTyUwaw0glAEEtcfmKT6oyjp75
PmKcIPXHbvJlEdddj2ZEkDORNE/R3ltba6X2SycVs69HvYsOvEYtlw2VlUDVj7SS
XAdlMq7sCF42IMrrTnhE0oFLD1tWBNLlR47XMNffGWmbrW2S1RDbfJYPLcEbkHoI
jqzWgEcxvJf5dk6A3iFf/Oc2me4DxqyIw8lJUzuPWe+LMBRC3X3IlcW1ceFRf+i1
Ot82skngBVxCfK96cIdweHi0pN+6KGRK2CgF7TesfMYgSYKcAFrDA5q4KO4sWrDR
DOIN0VoGj18tBNzxyTypoLM3HVn0ZM020KBKTB7UDd51jRg6ixBtBXLYtKcMQKxu
rBejpThR+jdOfvieUvsQKCBwMid5jvCjnFFXMcT6g8MZbGZrGAkm18VamL4Wiu0y
Rtg2Ol9o5DdYWRO6bhQmpkfHQTZz1y+Fa/mf6AMfK3+wOEHRN3q69Ep9PpZQ3mJd
oDQ6wAPWb0zf4Qafwg5rnY4MJdIgtuzIk7CpWR6HR83i79d6RnF/fNvHMHufUot1
Cpfe+bwbW3/VXHnjOB6Fp6zKlalb6R5bq/Sxqm+gQtgbbh8QIHnG411LgqX465y5
AsnmgNKtx6gyUTbpbyhZtl/BfE3USzWxTanbovFBbHPE/lJv09/IZUymRpYjSjYV
CxPJCYbvZZ5rl+xwHW0iJUH0Ii1bMCQnnWAn5wPq8+2x9dW7iR/SK5HDYgRJyjh0
u0PQaIcdXL/MMH/rK0suXmVcTYKPL1Z5t5ynTxvnK3/OIWz307PeqFhCOSd+TyJl
3NoIOFsGRSNueySrTjagnwKZ2LQJr7Ya+XdyTbnJUc75tBCQTq6Njx+K/mQ+zHuY
hyIGGmRH3s8eq1kVtjBWv8sDev4EulPVdj9cPwETf9FIT97n3piZVYvgy13PNLZJ
rCaDr6pG2efjGwDPzN8NUUquI5/0JKPAZtrMfBXEqtzQl0CUDjU4EaIVXWws9YUn
eOONJMDjPV+hNLfhmwD1LI6oYOTgDeK8UPLktSIHJTXelAE6Fo019tYHNM9jNuV6
DSUJlGc70p26KfDvzYnKUh4UamVYZFZf4PV49EPK6Kjlhs2nHSUh3GmbF59BEYH3
T5mwJvh0kg0ImwqDx4YN+kXtC+5RpIUpjYVTZP0nYkqneBeeVvuhVDM+Z1w8tYB+
/IYW1LxmW6QkNcO8rQMFq9OI1xseipMQFGfCy6yQJrALooz+t3TsjSLtWpJlC4Na
pzSpgw6ZSRitSL0Zl6dfescs+UsndQ9KT5t/KIXEaVzpN/kPEpNokYnmk/jEmUph
Y7hn02RH3wXS/ydY/xXHPpI/1BLtN9zSZzYgsxnpri0FPqaqgV9LzbZa1HKEll+c
wJbKeMljZ7c/JxC2UsvjHuHimZz7XmHBrDBTe+vJf4sUp2Re24EiBESNqH8OEZH7
lHh6icVNd47CE6PvEwuJ56QfZUKyYER++7LiQh23k97o00JmtNoTeGDw8g8Ipqlr
Vj3y72TJfQ5q/mlGsFBASQsP0YDFZ1Tlk1WMD1rbX8w0LF7jPCLPq/aqmZO2B5bM
FKMKcvemrnfdw4nJHLf9n7YiYXpFfQKJpYfB2SAxf3SRlsFeLa6rugHuA82T+OUh
LwHQ/xivFXVapiV+cbd9RGe+y06z5WfhHIbezrqfTWsAtFhaWcCoCbBoO1jE1JZy
hXuI1KgUQ5QmOJDqXG9mEXq7fIBGAauQpSwLK+5zFcBuHfK8dTJhF1ZZqGPKYTTP
gY7g+Oz74Ar/+Tt/uoQo8CEEoEWo1ovhtN5I8aKOQClx600WMvs7hV8R8xbRl+o3
bCEM/9zOLQEU5yiA3U5B81EWlvZrR1z9vhr0OFyRp/YlIWaC4l1xWegspEEuW1Qk
XsSXG670Adx2P8UYfyfI8wXyeQyB5gB+/fUxVDhQbEw6Ti8f4INtIkNoHLhr/4tW
gsV7VQlay4h2piShoefDjIjeh6quFkUVrHGgYiWHw6Gp7CDyP2ixxbYP24BCoAu2
QJ0WOEyhjjgjbKibILWKIfJASoXFrWSrCrsas3QZJQObM6jzbzfRjwZDgv28mOrp
D8V0F5zOvV+JJy7r871DHLYua2py4gG5sw9aDI5P5HRVzmMyo6rmeh2GkoqgAxg/
oHdqzROdX/Jlh2InzUDB4r8ZxRITewQVpx6jYEp8hu6gq3Fv0iYqelPr3w7PJAaR
XvrvJHSIyp56WvWuJ56dMGrJEc0jnoN1bslUlqANhMeJMzx3pOesnuFxFXNUYBxV
gmhy8i+U8kNDq2vFVwqt+FXS2kBdD4BWGm0h7X/qfrD3H4570Wp6yLWQ8GiX7BB7
+S/Qe2jTjPL5gAQEcWINiynoFdnEak3kY0yCvjiY9MlZZVllsatPEKgwoYo69Kkm
A4GgNrVt1w47EpdlzfqefNn5s5envuBsACY40RKNorMuD1aXIezmKqBc5CJppLVX
JMuy0ozAui6Z+rg5YIeZCUvBcAECt9gN/aaeHSIfEmceOu4cZELN2BL2nhrvUQ07
uEh9aC8UGNDuUrOPoBZ8vUhpg4+aCQEn8VvTAnDr4SaoYez6CioW/dDlqauGqrnG
yJZCRlbh1+LsJJBr7y3BpRHOJmfapZ47F6fcQhol+53VJngIHSyPD+AV7eJpPQei
naH0P9+XMDbOxFBpTjo0lYSZMGHhCAKX2efyWevuw5gx5Fj5EYpo8TuF4emZavOO
OTyByGoUfY33O4U3aoJ5clBm9ShLdWRAWnt1Y6Swg4t+V4CisvkojoJ3Ek9G5E6Q
F7OC8JD4+R2K4D87+UL8tEAIppOK99ls6Uu+k9WPZ1JfgXiQr4W5gRTcD45ytu5w
PNNGF8pkq4zYt5EI69a+fCm4pmDPqITCcrMBpcGhH45vVS/pSSBtGtpB4vRaTw2H
9jLUrG0Me963U9F/8wCvNFlyIo/wnXCXMCTEMmIKaMwgIhyQ5bI8F5rNnSJvX918
eAJlQiw1OFWlopn1vsx7hd8527JtYTuPgncBiRDx8E/CDdCez6ShlD/QNfSphr+5
b8/0DheDS7Z3XjqVrdbqQ8pB6kL1QrdQlxVTDZw5eZGA0TVh1Qv18V79eSMROn4H
FJlvjqdHaW/1wnOxUMnMHmhGg0nHbFQkolbT1XOzDjWDBAQgZwcjCscY0x4K/ZvA
q5ESTjJp2rMaPn2eyljr2Rz8yqBYRCiB6gVt44tpl87C/kzuKVt3Lj1y/4LS8ZYu
HvCTaFYHfDtGUOW4URZsVwV3SjU3PCZT33szs4f6ckzM3wj3HBScGFgBMxwEnYgk
FAV+lTmcJWQeQEvMknxtye0VceWFNSSjhDdK1L47DTqvgNhUlz2Pdl8+PGgfR15e
H6sRRaeUIqBF+tR8TYV4Lb4/2VIUG5UXNF+Dos1qlTsqewnWb7jHMEFZ7G1h8gHw
edGuR96DyqXDsvr7INuOC5ztNkySixiW/uQBa0rQ9X2SXXfH20BiI0kvRBAp1EST
MVOXFVKznJd6DhwvVe+LY68fyqq8LorlW/TCX1pkfqGvhXmemmZ99vUStidOdfLy
Kcjab6LsR29L4Dj2UNwO2dqsqf3CloAxfZ7AhBgGHxJt2J37VrpWs28WDjPDhoG4
ubUmu4xk4qKkAFziow8AsHNU0rDmZO+Wwf6yWP18+O/IizVpabRsxapSov8WdIhg
2UMpMnp2Ju/EILWqgv7XDDIgrugRNWZ8PN5V9eb15NvCtOkpBuz3H8YgifGk+qQz
8DJ58c67q7tXvxDg0PHLkbWME2jN74PDmT0UWScPwcnce1936jUWpjnJ7otjMW0S
qmHOg/06RZXg3BO4aIMNhjNVjyEBbXOWfk1vuMCSoHrAIHOfQtV/o/CH4y0det77
taXOmupzHn8X/l2AF5CdrNlXC3FbjwLgkzEXEKxMoOH6PExovkFAVTYBnPwwQtAm
AESSxnMmE8IYFFJJHHRgjwKvELQf2MVqpcfKHw+L2QvQE1v563A6xNrfJx+txZ6q
65bHUmttFbteBxle1tbZfcYNmd4B7P1Cy9NCR8anZPpWpQuggk8hjkGGqJAB39Ny
w0zuJrvaJHx2zWUavrBWKGYOv9r+PqJqGMEeQEyVkQirnlkJ9TYgGJbOQ0WU9xEX
C49hMo5+RRgp19JcqxKbb9HEB1z+RwRBmY868elslwiId2OOKOKCedpGRDcmO0Oc
xWXRwzLyT76CupD2oWTcaQjI1jGUFVvy/qWbWZekNxpm/7whd59jr29JyyCbnZdg
SG5yr1l8Ua7OIxVug6wPUHlNWjcve3XMTbIDZr0+D8IuOsNElZmOy+TauAeyAepy
URSnmcoW+MU0IWEqoLqhYTJ9fTgt/zmo6YyaD1fAXmt6RtMptAk1PcUsoJ8TDfun
EjjFK8H0jdsIYLoVQxa3L4NWzT86ALnG+lGYTKXDm62hgb3P9vPypqY4idTkCvl/
LjFk0e0swDsSqjkujRbnzBilfR8ATQvC8oGDM1BLykHPjGz3pLsy0DzLcxwChV28
pGBTtmwKeSZ0d2A83cqCYSJcD2gPsy7mlOkXtPVcHbvTGBxKycQ1UcCofbDQauuU
YGnpbFaA4vAHKFqFOQsH+O5t/MqhDGGSR+9JZLjeh/q8Ieu5e1a4/n4X1/w5LI8G
EiAUREstIWpbYN2/EmrMACLY1eKwUXNdCkYD38GMVcvO0TeH+nAnM89DjQsqxRQs
mzJQ7plVu6CRrnGNMO/+Ctz+eo4cJG4Jgbsgesn/37kwtvso0CrCUyABoKAYqHAB
pGJanq/ma24qQ+mXTArnAWM9WAjItxtwWKlAWg0gqVVGOkvKfFbEB9xdoRwHTQQA
W4UiSSl/RgF5jDAoW8k3hcOCg16rknm8SrQAbYK+0ocj0I+NRGbD86ay/H1ezYTm
XSAuHsAtZu09quqqG7D6F+tyNr9Al1NUhBHkDrck1efS5XOqflPznC6V2lT6O71P
tC8uC7w4Elg2VBqTmYtHFlYyx4pDtLF628m7bFDDdHR3ZBpuF+aexrP6PV98oi0F
+VWcW3/hhh9tnOaSgbNUqbUjwzaJ1ltBOIcO0qD3HNd+jwtFzaqSQs9CYjYHLEnn
1c1B3yKx5n4ODlFlD9yi9N+ORBuMrSUVSOBczZQ/EEBTd4nUAp8Nl2AVB7dq9GIG
Zp+EX11aGMr5SDCAuhGFcPlEuT6udtv4ph6/hcrqDl9nZxAedDMpd2DsB0h5dzx9
5Wrc8O9NCjzNdfYzhTwYAobZctIT2/Lr4APt+3MT6Bnuv6dreKR5YDOqorM6XAHm
jtBQaPIQlAbHq6gQJKjVhzpxffP2FE6BrBknlk4+N8dqzLZ0K1K0DQwiweYlTErq
JzQV6teIGTkhxSdwhseCifaMEzYYh27+Xh52hIi+cQoe62NKXEdRbVDGmyWhWAer
E5xoJtIRi8xJW7za0Gk4wSf0pQFXfOusSVkh808f2fYOInuZVPSs2vAAq09kWC2D
KpFa3ipdr1sr9H35LPJubQdDDlKpZKVKkYUUwubU8XcdPXgu0h+Gx/anTXrVLHoZ
22ejwESVC/WArG/CfebVKE3imSjdU2YqB7CCPVo6Toif3c9aVRtUJTIi9BHQEHLQ
XXqxpBT/wBfbvlFhPqJgFOx0IH7tcYlX1VQuTrGnTCFn/hdWNM64kqV996N+vQEN
AzgPSLC7du93TOi6kRoevDP1r4xhrj3ZWgZL5FQLlA/NwEsjF0S9k3wyODzKKqCo
pu8U5OK3Bj7Qkk3CraamkvSBS+B20FgAR8li7t0LsbY8kPbOe9Gx6+8q22h49Cfn
d3dnsGobkJGPfD2fTaZz27O/sTMnECoumaUeDqbedRqs8oTQEz2zSLIOgWC1TjZj
wkr+rWhu3x9dgJ/W7pEgzrhiSSmVBlGf8AGUGoNG3zYFcrGdtyylmgCJl8NviACz
cI0JFMboKfIqSlI6XCB2ev0o1VYVv99JOqbFWseQ9eBhV+I/g3ks6DBp8JR8TcQh
GXN2NLjlmg6DXn5fNYFxv4ZNiNTveQw3ni/W0dtvGL9V8JdwKBV7sNqQegdrQOBq
Tk+YN0Y9Ps6vLEsQwNNyyXfUrKab9G068xnfRgaRpy034dZCgmUWMJrmwVhiNu+j
MXz8lPVcqDG2BrXECa9UObC8hBEen6s/WU3bx6w7wuf5rj7RzMWs0imTjbTGNFar
LSrgjyaSbBWqUeTXkaWJvMwx9Go8mQzJrDlbCkqIc3jZdRFj0jwUaFE6e0Zhs36E
cTOCMhtIy+cVU2Y+2Wy73UtZu414UjaxZ9HtJ1M0rYrF0Cs2i1ys6xxdO/WFUOgO
iF8sjeIK5CIzOfewWPilPV+Vo4mg1zdxx20KqwPngYJSzekeRmrvwZhFAY4ceAlb
mTUL6vrh+se3ExIK8HiHEr0dGN3G+HpdrDdDC8ZT8amkraCWURkfwUQWjrINqsw+
4V79KDPfde/stMVWOGHubP428SB9ilGMCneqyjl+/T8gOXcL5U+OZIO8i9VvEpsU
51ve/gQERTTWHQbxUkt+oddPvyuxHN5yEL+S21sm57nLsCp9lzGDW41h0yCcOE0c
77AkxyArD03wxVIzNvUUY/KPxoalOZENXA+3guwuj1+r1F/YXOOKHYc8SHL0EuP0
WNTFwvmz2ItZEFaKjMF6jhgtysWDHVBkbXpwrgY2kkFrD7KbsLjpd5FFqUrvbo3b
DP8J1ZiHDc9+i31K6YaZa2/b6exqvfnp7jbhmXGiKW6wK0RR92Q9ioeGt1pi2lLS
d9NCz8GXr20oXSxks1YJEEM1xkAz/+iatp7zOuONhVxe1nAK9R/3vahBMjZINkCv
zdPZ8pncY957nsVRspLZ593m7QoTzfEqnhUxu9Nukv2hsnisWT3DbSUp5TTM0kxs
k/EjpsC8j3XlwTDDaufuQHB5P664IOG/nGoXAezMRctrkQ+9sqhhfryLGBx4Ko+W
dO9ou2zhDUl8wtWHTsPWBEafaSkM55u7JbweUboFj8AOYQZFBHyGvwnRxtXgJCnW
cEXM+kj+krAmCZaEdiJKkumWVwp9b2gTteZMnzDnRUMs5EP9TZeSE8IwVpEyDFQd
/Bi/DCjMGiHiaWeiSqf2S13zdI3pdw6InTiTbKcKe6ZnvwzY6EiZEOeQou/QnFnN
7+R9GwJ1WMkRdX+FBt++pFMad0m0XnRm5zfY/SxosHBwqtdoKHp5k5r0IgPqjU+J
l02Oo9lC/sPOfRmTy/uBWcPWJghy3w1ssDhXLTDdCfrj4nr/5dDtxUJN0vZigI9r
BRzw2WKETaV7hPyFidZMZSDkc8tyJsjt9LsYLf76rbAwg8csZBCz/uPjJJOH9wXi
jU6roZE61NHye7MQcBnYQfy3AH+E7JIDUuNxHCfFU8SxB5yJ/n28Qu+kvzvZQdeW
GxHGLjxpHi6MVoF2gPHMklAX8d4FiyFoK6xHdazp4MFmmBpJk8foww+mpSfE3z6/
d+6T9jlMF588JJ6BWCOWRjnB17Ew5xHeuX/FMw/+t7rHoG1RPQIjMULIID9/cSXI
JLOTrvm1cFpreGm+YHnrE1J8zZ+L2hSRq0784/l2aQy0TlF/pubyblEUxck6KbHN
12vkbZ83QcvshVKXIXabPfFRQwGmNH1DhMtdYNWfOX0NVUbSuKGCoyPc25pm2x47
QGbl7d93SmfhzoCvQUe9VzWn0a9tOsF4OnoIPR5voB4G5XWauENEWVWS9EgbUrz7
cYI33rSSLlEfRlVKNIDvSRi/GjcFXTW6rAmH7LqSjgLLnkkddyJiZ/9sD+0EcN4A
wN7eyBWbBbZzaMfQeuAenwxlU78vJtx5vqQs/VsTl6QMRDOIsCEqcIC6003nw3KC
Ccom/XoZywn6jdUsUp0nhZzLJI4pd9MTYxMs0DV0+77THZhApqmoft3t5N9cNgHn
G4mD+AcsMYitRq2wl1F2tduiWWMyavUCdgIqMzt6N/hDvbF73vNqWal1gc5QXFis
Dl0PjyObn+1qHXm9i/34kMlgRR+hp+r9Q0VQursOAnRr8QErCsg9c5SurHXZu/mJ
IstywsJZ5F+dTB1hVCe0C2wiZNfahBCku9L8Z7OK687bP+i+XK6Lkiz3Kf4v4D4W
tLfdi+teXUg+1RQ4TVMIdg8UZXLMq9OxecEsbA1GViX6ejUjkXQjnDy1VtRGnbvd
bdmQw5Z3VJhTyrdWRt2CJ0YXU2AfHdTaN176F8m7kx33oGNWsNryppJ4pk5AfN1c
CiSfFOBCgtKNrKSEmLg1kb4yBqLALw/R5LDuDGxtIS/2saR3opHaXtPlR8EaZlLA
TOwtg+hBQTIFH6gGL5IGuE6TWNpLWUggekd9/01EVRTJ4fOjvF44kQT3CjoKeVOK
t+hMIhKS7mJlvckau1Mu5b288B3ADujBBZ50I0BCZKWcGquUXRx8yiE64LQyCjti
Wr5WkRPe7TdOevGRWf9jM0910x6vF6FTanmNaqz09m9mS3VPp1xwTcUmgKSexkIl
JBSBeIPFWOBri9adnEmCNZ4jw+jXKr8Vot3xO680MX7RNK+OOR+P/G5dOLdIC2WB
IfiU72GYxNsQ+ldFWodIxYUdfhF3OI52nxHVUsyB/lismPQ0ShHoBI8V2D1GFAKa
XiyQoOVylNlZ1xk7juOCcfVboEZnzJK4zkLBGxOrMk+RCS0wBTcQDFvo+cAwcPnX
nCpN/2pALYsZfeMYWDL1nl5MNlyWozVAwM+XrP+Kb6W5WQOw8mksVA1rTY6Ad6AZ
NknLSO9X/oRGFQ4EjbDHK7sMNEq2c2cCv2V/ulDMSjU+Z8wb99U/DIqAZXnVb5Pj
w3H47xBnZQgvHACVx65rFFfsUT16BxSkX/19VaUg3ni88hOSWZs0NN561Zn3YnkD
GNutBbNvwtR1ZO+Tig/MNYfxc6U8rje4zbNDt5b/PBR1tk/Ku0+QeqgXwWfsxNL3
8U4iN7b1XF7UDPYvxxLJiopfG2CjYj+TfzLcapWUY54E6bIOOOAtTp8I12ZIv8WC
eI8hAJA59VRbz4pntQCSj0LSJGsikQq/lzBxoxdJUzvMM4wEzXg8kvdBrRz7PRvO
Sx/6CZJ7Vuo/bKYREzzai/y0WB/AgDclHAyOx+Qn0kLKVx3DMCIr/Zl/7ctjUpvu
ITTT3rQ2qHk7wHkvIiFp/l2aJTzllgnOZxxkUN97O8wIt9DQalGflS7Ex/vP+lSR
PT3YcEXb0wExWBJM5NX0eG+cmt73IAtAgQvlIzHvuMaFAHBx+JDrSjuAdFo8p2Dy
xS82lpp+t1L7O87+Xu6dthESvfjpJFVqe8oUskZqCTKMu59no3eWPoRw/O4gUHuM
9ZMEuJuPWzgFLfB0jkQDgdpOV9TGhsYFvuvVJObovct21fJlJxw0PShxLkNoj/26
icqERkplkPw2JENFE20l2DnJxo9IyhMINtAv3W5qx4Eja3fPyBio/DRzrdPuWddv
f23azsPwxbipz5plHhVta1BZAYdhci8CrQMrxsn+vKMXvqamoMEN0LFy0X5opOZr
/2qHDDY52Dmcm97IhZo2DHo9yDuG+HA76AgimXWQhzWYqjeqY4oexwEMdAmn+uDv
lTIUFeG0ExZPnvq9PmVvkV9BswwIMgQPhjHBNUqLjt64Gse8LHrJSdPK8WdSedsu
eiFMrVnU8bz/HoRMT4J8VOXYq26/DYP9gzzGViPWulsYKc9Q5xCAg4XdamzC5Eyd
25WnQud4Qs5Yi3rNJw6HG4JKztRNz4v/UiUtlCFTJPmQDWEwJNGXxVj6cvMhtcEG
XFtCbtFnOcU/V1oVS2V9JbqnELlff2ZMppDbVCFPfiN7r5MG7wrjTAti7n1+U0yU
Y9y5FEyzvrhkYbM9Svp+ADbZL5rvpnfv/hpWXBqCKmlbETaDKanPo8orVxHmbroV
mSiVHOFh1Qw+buizvF7uJJQm06d53CiV7f8v4AKUcKONO9uIdJLWjwC0QvCSgNy6
xVdwYI+F1xCQbk9GSDvlfJ0RfgyHA+YDRPKON1AdrIFrDRXhisPjZXZ0iMq3XSdN
2Pq9CA1ywm8d3stK+OT7ckLe45CmNGxCN2eJnzSWfc+n7C/UWEsgDkx4ntGTEdXR
3GsJEyRLEj1i7B+13fkdjEYpT1phRUOpHpqlYUaZVam7ZyGnhScG/HZ77a8U+URA
6IdpkasC7phdWIHcFi4zVerhhZAzY8/xy2WxsjQFguU4HzOJBWNLI+W3tu1I6tjY
X3W3jr8zVd+UsdylbS+HV/bSGCWRMpEeVxpUpxRRREikO7bwPvv6kAXeF0akZfZe
LPhYit1pGPrJlZyRY2P0xtqlFmPuRb67EGPshxeeyaUn8FnNhDJh8e7oYz8fovJe
LRN+TucpzH2zD66MUv0ZaGIk3Hf4sotSI2FchUWy/8rN5BVSPPO4G0VOYP1r+xj8
39z9Pu1zVA68tA/vq3hPY8R8FN8fl0VELKB4bQDJ5+S5cCCJggVmb6MCIQX3NPBu
FyAm680oCGXU0Hr3R0XYN/gzPue8sFx4VZ0CtV/BxqdIlWkS44kKjxDA6J1A+FXh
CRJZUz9kmlDVHptm9sJRRtzNYSd2kkpgppk+veZO/H2IxGsDLNm1UjhoLjS2cpck
kZUy9vSWHF5LSJHG2GiC5cp2DgfybGSNGBMdg6mmPychbObmhHzpRQJgy0FQiRxY
3baZZjble9w5hH7r7xZpp+qA+taeK9AIrHFzyzMlahyw4HcF2fTD+I8UfOmX+uRY
fjI1VkCXLuhlzroBKb06KzNgymVlkhlY8ul1pZM+EIb9Q+vZU9asahUsTzmszUKS
j3Zb2JMwtjqKKSxwMhfrSuBL4DOb3mQyHJIyhBy0jb1SpAB3TL2UmZexFVRmD4sn
GzbxQktx0l8Cbeb6m6B5aBzoM6tLcZ0TE0A9lARjrQ8wibFjIxmOvUo96oZym19P
VmIz9ppVF25FhO4iKFwtF1XDAd4FrW4lQkZ48VMczJz9jByPlBTd6KT29oX/2cQQ
DvIT9mlDNDHEWJofvYYKLrqJY/wRa6rzwOL90uSFVgMPWSUa9Tg/SXG9IV8PyDc4
xp7nenoWCCaH4H+l7OEgH4URw5eTnFSJ26nyxwcJ2JRrKYZJLnF05k7hK6w1YjM7
UdsBsFq1srAeagCOH1pm9cRl/kn8pQ3T56UBy4tDprAfa+QvcI04Op/6t3/A3OQ0
yaJ2q+uq6q+Kfptnpx8TrCTkOg75/TEsx23vkfMqhRuJW8NluhJ6ocu622ZZyhAN
X/T++he2TCDz5C9dbtfz5mzJn9lkx4AiO9plp8L+qgUoQxZEpwOIPnrX8xpE7yFm
eEUOLZbnB3GxRaka2eyb9gbaj+IMY1o9OjbYS93l+J6nKQEDDKImkQ6kC3io3oAO
`protect END_PROTECTED
