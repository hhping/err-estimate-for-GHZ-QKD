`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rI0t1yFIeKzhp8rDQjy0Cb9+mbrBZk2d/A2UVNDb7ynSisQg/uSRLjCGuWlwh993
A4Xz+k9ZrRv5vAL1qf9RJmyfnlDsN8MYDN6FHsdzA4oStbOb84E3KFuXh9DldAFB
m4fB+50jmMCR/Z3N5kdvnGIItgIfMrJvbLIuVx6u9138RIDc5KSHGRQoF5gFKOeD
Fgm/TttKK4y7hrlzsWcKg0BpNzZwv7nJk+gwnusJG/dZSOx5DUZuajX3XgBz+63X
N3Irc1Nyl45XhmaxUv22bTnQXrpY5f7nghiRbfXKK330G4g+YgNfrVQZh6zbC0i/
wINb/AHRwicyUZ4pvCYiTKsE3NHWTelyHlACGTOQ+edP/2yvNj4nF/8+Z8A4loMr
E3CbCcggdXz0CvmHO2tQOke6SqpJa8+u7w5CMTcu4Xz3Hj7xgSYbeVY9x32yQYu3
iPcFO7kpiZ0geVjH3aykab5wGSOmsmsr6CkjKznKEWg8LY4u1ZveKPRGQ8+18eTW
p5PP+NLoV4GuwgILh+u5NXL/8xMItQtwTXSVn38MqUs2R/R7oU3PW32+LZHE6DQN
X3gafiBbCuWxC5Br3PkgsNa5UjpHdEFITscxINQ8S+UX9EwiApWhWv8u8LI9PwaJ
gdOkrRM7wiJpdZnVdQXq+fjM7NIjNBBJRJgADu+Ey027Hhfxe8RhRePsxsQSB3Wl
nq51pmlHyxyUYOC9Qc8tRRMiLLcS9+oUmxL8Hs2DxYdpYYZAbWgmV0OMZHf9pYdE
dVoHx8CF9SrwcTbfQSpBiZTBJZUwByP3+YxMLtQ3elBVvQIckiW25fA3iL0oF750
7ELqHSOt9Mr4VcV6dTHAuL78aXsCjQNvvv7yeuO5Gih9g+Jp54MakgoTy6CMR9Q1
UtDY2+f+gMHZwUlpWUf0nro/ecvwTR/dnaDumYfQsjJcZjwH3kDIR/ZXAhNdWUx4
3WZ26nT9ESWuwd+8NKST+JOM7kfjNvl2Utd7dGjCx1f2VWzKVPG6gbNbGRaPtNc0
2jkd2PNs2KtPZ4b6ZQ9wyaTaf6UQacEcc2UkzPLE7c+mupyWR/0SA33PLWWnTzJ8
iVL6yPpOebLcsCfuBX4VP6s5+LRDxZbv6TH3/06BggBTVglVxGXWY0uPMDJLWh+L
32FnW2KPb+4PGLU06niHwi7dgKns1nMFDWqW+eMS0YCVyErCG75EsYjR9JQpQ1Wa
8Yl1g5VtIQLAcUoOGyukfri7hEdOAQQ2dTyiXEmtkvZfDyf1395UuKvg+K13x7Zg
hayQ7A/uo0oISkEWoIKCXmRaQlGYn8Kzn24WEy4VHOD2V/EEb5IWEmmrELLgTZHF
+JpRJnrXgEaSHlRTX69QgcW0Q6A2wL/s6LC26NqoAAEulKvfY7T1Kl/xnqKV7vmN
4NMiWZxk9F5D0iRIdN6hFiJZaXKfGdOl6fLdxv9zs/OJqnGaI2GRorb2pYR3Yv4c
azyBaNNLex52NYGZsDKVvtDFhngFA4HFiSNqtdVylMTCJwy6Auu05KS8VaoBQyi4
SkXQ75ly36n573WTrcrRysVjlEKX65jQvE5beYVBpvEv2dGozG1Nsb7WZzLDlP4/
uBAucMMcp0paBQ1lnr8xUgbfl5PV/d8mqg/WgxFEDrba2rK4SpKGNAHBBdyfCwfW
F6SFALjufwnZdOM2dpM0KVinRCsZM4owp3NW4YRDHhKaJ+XPB/1pl/PtQ4XpG2Mm
5kRrEYFATCyhyaqI6tqJxEMhDUczahgFIOW6a4vUn3yN5V0qry4zZKm8tfQDQ4HI
rgdkQ0MMc5pv+r7QuBVI7Bc+RfeCF9wEaj1U+XtUpANnLBnKLxKGMXPhx8iYuATC
A1Nmak6x17zS4bDalOAY3/4D7LPS/H+1FmcYcx07Vq446qg0kFg/w+62SUVXtuaZ
aY9q5tNoWIUZ9boMnoooSujmYZPn86mQyRGF4gB1h4IQEOyQsNmSvQPUDeSEicn/
L1vUxDgdq6k8kUtM96zo/EmUio/TPInVaw7Z7rac256k0LVOyPIBWp+aBCbyadX6
2vy1lekjV/ETSLgebui44RnlXFwD0u7MMq+0VpTRua2XnDovjfHeJhevWk2LcjoN
pPFP9wNAOWnNGK8IkakE9depuOvh4V+AONwELTUvy2h30LybRvAnhKsetQf0B3Ft
LyJII+8jBnXbjd72pKAlyG6lWUaVF2PDS2GbXwOvT6Gop0Tfg6GbzJwINaDoCyzK
GuzC5TZqIv9kC0hToQAiC5rXyLfizueV8LipDkOzJnkJDrYexIxU9PceolleAY8L
sA92uyM765t6b47l5CwevrgQt1JY4nWgDJ2M3KWlYPwmQ6cnyjIcrG8EP31kj56Z
u+QGPpgZRuFwraf/IpAXlViY/atEL1K4E0jylU0USEvBvovJtY0QA9grFpcWyqOV
hzOa6UxXkaxbmhaJzq0WH62KUqcK9lFl3HZB0xp1V+KBLso209vQsSOPBiOsaFFQ
XetWGWeDmiOmUY6Bym/Hr3pOX0uH4JuSYlyxAJXXurXpai2QSRRXOH5mxlLPhlo9
M7mAlKgwWKC2r7WZpJpGmgggDpgyQiHqwY2/bl3d+C7+aRzhUz6puH2Wyah60L3P
fwGLw2plP7WO8sLlsuMcppAOGDXsk0XaZzLDKI+8+TNO0aeg625WESbeB6RGCpOM
7MXETNpaswg0PCX1fWYDRVkZbd89y6ERGLfGayaCWCKSa4zJhjwwFdnpjyRtFR4e
yF2bEl/zon4Ch2PgYMS36Z4/+P+cAzH4PH0zSCU8df6juuEWTR37K46Gvv5Pr+cp
3gy1j6GKrXAofKS0qbaeFrCuPk7IZAgGY4V2oYyJwlB7KoXYmA+t72tXbpiivrBx
iu+r3ySDihV6HG5+quqTNG9zNXxXUDaVG19x/EYBAPY6wOuvlI5rmMMbGNCQVy56
hDCX/mx+giauolwqd9xN0w4DyPBH04BR0yJ29M8McoM5TdZckPu6xRlUjB7pIgea
ZtxPAQORPJI21asAXMHAC9yKcOUmLp5y2p+BsiQ1JiRXj0E9qZMoxX+V/XLb9Yt4
bDSTxHjcNKzaY71Or3eAXAUUzxpYMIfLdAtOsFBp+B9u3JKlIW8VrmjcVCROi4b6
A/9BVhOtI89etBbhFZ44VtHco0DrW80vzF4IGvwXyC1aV5VA7zvNmZMg+diEMo3B
ynnFtENPAATi0mhk9zuiNY5n4V7vdGTSkGWnNWuF5X8VymPo1eUQ9Cf4zK9zEXBK
bReEGh0xgoiWnl/uVk3RgYDSPmJvSz/BKWEHiBZfu0PnSayEYwCniGd7MdU8uPTy
yL4mi+eR3D+CKU8FSPzQhO48xluTjG5tuBa2MRr0VAdQ/aPrzcwfcHVXSz54pDu+
UtTwmHcLDhoM0M5WKGOOM9MjCVKK3pCDKhJBHQEtN+jF1l0fU8emoe0HdjMfl7z6
1Q100eq5JQA6REDMTQYHesKANY+wQBpnOGGonhstoSDxGJT3skhLoXXRsf2cGe/N
/t5mjcjail1MQu9IjSh00sJO53ItFdCHjSD6R3FOIgEfBb8Pf0XQOl6Cpp04eowH
freTioqAlSXQZLy2iZFl7fVXy+q324xCXFhkEQPHGKUSpGQKGvHVgRUkWMnujgUS
GaWLSiw5gSgb8be0Szul77/+tZ4+oNBJgsK3iVWga+DhzSNHE139T2KqOFUzPFuM
aWn79MwA+ph3I6GTu1GzM17vvVM7ZceVl9O2iVMCkRHZfAcaLlqV3kLUVXjEE1r5
W4VWUj25dlmiqSxwOKnJSHnauvHyKbnjvimrfAKW/dYH7Qbn8iKanAIPKfjafkOm
hLeiN4NwpgtXKUkCww48ICh0IPDdUoHPMmAS3O4s8oGi7v25oaYmIMwEKWRyWmXV
7819vWi3jRX/HRNbriNnKBCeF7yu5niCkplbePjSPXLVg+5aNY4n/FTiRGUn99pW
TEwkZRjjDg/nkV75In9VxNWoxGvmmw2jNZ7pcGjgDQrrn05o1dbdaQqtpqmIAYV9
vqRIWnC+n7f13rtH14W9lCdTj13gwJP/XBQhz3ZXegDjcmpuT2JFNmqTUr6Ctn8n
Gb/LeFKEDpNmj1iwQQNFWb9hEcL7ur7tKgXejHXGsuj1FjSoh/a9701xUSL6rJ7j
U4OSkDPUMmzDxQ2fmQBdcrAftjCo6dMaZThZtotEaD+rWmIIzCKhCS/jrULXjVr7
KuMM/4rIsPZVyciIRHtolwIYOATLKdfXBrR3FyWiu+/lAlsCiIX4pZvxTVee1tN9
Qs0coEgYmpW25+d1f+QA6oTIv0RszUU9JsZ8QbYpG/v8VpnboShSeX7A1l+rs5Tv
44UBW6F7U/DeIDWPdOdZ+933v5g2kB+IeV7VFfNHrYJ5oqzttqFBzpwegeRYPU0r
bBCGPUl2P5zmcmar5MG8iVm6MsEdKK3WkWE/FnahQ1zajBFbsRY1b42K+wbSZQVm
+5VWEebx7XGPCcxql5hv/tb95WFkN1dVMYMMZ2ZbUYKoPEWwh3tAadP8ybfHefUO
FebiuaB0sElwa85b+invqNAkuNeASlo0kQ8MVq2bR1lfkfCimbLXrU60hSLsNf1B
zggZSHoQxW2zgTk7HmglDpzxx1WQGNS6LVoMxTcvRA/gT12DMbVACgA21IjBuyx+
/49pnRhfGfHj93iacfKVwHT7xZy6A3UQJCHoqj6vr7HpzIdTTCpXOwU3WGD6jnP5
H8a3fNfFsG9a8oASg1TzWkrHoOpgtvmNmV4MW1jeIgzyjwEuYeSzfD34xF+oIoeP
jVJabZHgtNm+jcR+SUK3CcCbYTUYmVep4N0ST+4oo3rqiAlm3B74lyTLiUciQNmd
UVVvSGIiGv0phRkFPr3X/w2cDgzonQpuhJJjbsh8Y9u0fSxrIUUkDNnUrfI7mTT/
grWo1DqKtvey/3HG6uGepmrjibwMZ6Do8l3ptEG1duL23pIjtqg1PBKjGjqNcZg/
dBGtWWfL6tmm+BlcRMKjmFsLNhji2aIJfmp2NhPp1ePMf9QlrucDI7qHqZtfkvPJ
iFwb2JMI/Tgh4S+9wd7+pYrrhoWWPkP8JwUukOzhZl5FhxV5i/KBIfmdtDzJTeWR
ahtOp/5i3VpR+JNTnry3Qr1WIP5movKx4sOl26fGImh2LylpVESM32RbIMg5ZpHl
KnZjOieKggVOqbDCq+XYhnef/fJkiqFOc+cPP9aU/+1IXDrN7cT62u0Hjx/ld4Ma
N4O9sys1K1MRBW2OnE6VtdD9MhGYY6OwTPJ5uZ+QLIMxbQJYDz/RLrZ8gvUgB1Jh
A6oWaLL8fUwXaslLskyOs7la0EQK70FIAeb4CFBd5ye8+KScja7uKXBbXWaxHlpl
OfPV1NUpeJ6k/patvF6MABcj9KIfczXoJpbP9EqEMEOwXbvULBzhkbK1IMnsZJLf
OKmB/myKgOi38IbpUqX2Xx4fQlX5KTgrbpVdA/6tlKeime4SW969NlWwEnfA3qCa
lsG7pUPtmrxcFEvl9nNo1qizX2kcW2pGzsKV90SrbBCSUdoDw+owH6e3MUIxB/ko
BZlWjY1l3zElounmAiNL0WbRAYz55LSm9VmvwwKgUnOlOvg8RismXKSnVgNx5gce
MpRENtLGP/bHkUuoOIlwxk/+RQa+GapzKpPiQ3bpBOpxSFwe0N9SJleuuNpLpOJl
6TzaATAMXpmori8pICxw+rlzo9E281j9q9wvfsK3oZS/rvRzziYt0JXQOmpjs7Ye
GgsW0o1sQiEab96fkMLjLn2ghOgDQux5UmHeUA2T+DhVm67gOJx6wWBvFMFzIBeE
ZMDrmx7W/EEWrjbxmaxSgus27k2gETsqraOvOi0YCUkXLZz3SoC+GWMPX69bk5Fy
C7mf3TDYxg4FYGtT0cAtDNvxJcvBovlqAXU+0tt59hDZXPCYUDojIk0b9/chrbVh
hFBzucHhKCosg4/qyYQGCUJSq3TgulAxiy5SytZkKl/sRiHh2HETr93iKdmRmbMx
Iko7Y0cVfUF9Fr/jmMkWPWRnFrN5C2w4H313Q0j+tt2w51/yHth5Pw5qKseIfQRJ
nb1kk7Fp5vkr1HUFAY5/O+0hlZVEVerCqmjyv/hA5NHZIVXDhMRGKGlCHiDwAWM/
RoLuIhHWYvuCJ+e8mp/vj9nLBHS6Gwf1b0qDf3/KNKdu0HbYPT3W9SvonchUvlYI
IJr1vN5w+x8ByLaHqJQhrDKkPJ+yeho3sqZQ3xn9q38HlFQPZXT8ZPEdVrfEIsPp
VfTxOHUUvv6KVHpwBo68WcEd8wkh6h0QBrWg6X9yHqTeBUah0vzt/B7KkL9CaK6x
KFPKdJalUrYb93ye20WEUsynO6mfO/OuFpwT0D9oSVsOz6TOi7OBHavM0Hqf1Rnm
tNuHEkLI/xFe5wbN3aJCGFD5/gLRAXD16u/iab2FehkINxVwkk3AKKUjLHH+4jh3
6uc4dVM9DYPna2yW9CFAiLNurs2s2yFUh5fsSIiDTX5go3NFqiiz14ItNnvJhdsI
Oszm6niw4UQBX93+MnATE5Cvz2Uw8c2n01HQ3ffL3LQG46UKqCgFZu5gOQBAfM/p
1qkMG9mFQ/MbOdPHx/vjrFhkkRyuXkMVKzONT6QDGDhuVLezMEfFQH0ikIhxz/7i
pO2GNntnZCbZQZO/771SN4frAb1Tzcg9/WnWYFNdZYblAlO6azedS+eD9+K5pkYO
c+yxEvKtFZzt2joFZIlvEob3Dg5iTWJSGFqXYFL56DdAR+4x8eQMptFBRbj3L48k
OK5gOnbxL0jjKooieKV4/parAW3lyVGy9sHY7a1qYkXs7SMBH4TDL5Q01+/ZsdgD
B9Wyk704dO3+qMbvfGIEpYrQvk6r8MTMSBQ7yKNAUTxIGqtIvaxAXinuKwcBujYw
D6+9D87TgRFpKt2hd90vxu4vXWqSFJ7QW8n80Pw/jeV76nVqVWuFiC6r5mYUjD70
qt13mAQ2AuNSbJcX5PRJZkKs2xrfR+tMjPF/txIIMr3pijRz3V0G+pczG9H21VCj
skbyTW8D1yepAhiVV+1uDIN849cQxZ90GiumsvOoQFxmCBB82ss4FYTnZjNsZkLZ
8tdYLB2pbECoNo2/pU/s3N5lst1BX/W0ec3RApAycPRRVCZ1wS7WywCCesvYr/2Z
5T7Z0Fis00lXgjxitn6QnjL0DYDQPQaksAp5zErPWkKIcw8BU32TC4/zvSC2lYS1
S0W0uO6nGmUDodMdD3Me47RrSItM2xieulPxxD0PG8LvkoD0ijiZCx2mzWRes+ca
sFCT7SI3ausl91beVMR+sCN1gyDNwX9u0m18Bhrjs3I7to8eYSkFTQsSqw6g0kP4
ORamT26SJD6m9PR02ccgXY/YCxgCyaWCguhaa+xD8kmyqnKH+LLPhetxJb+R1az4
AAkz/4+1xMKanXeCe2H8h7SuNOCBCnHJAPBA3EhubygStrl0avhIWYegoRG9nVHv
xD4k61zjJaNHV7gxK7rq2bKeasyoGFKcmMTZYCEuD8wKk/X1BOACuoT/DAscb7FD
cXp+aQTtHAJVuMnSv2cDbiqWOXH/uw2q7eKUpEYSLB7LIEHaZEDxB1nDRQk61O0z
MLIB+UvZVeYFT/dbkVo4Jdp+5YyE840CJGPbdSJH/BUjWjtfd8VMH2VxfhIEDiO9
j1RoBnVBheRXt7EtYNJPsZvhQ8yzhnqYJ9y4n3lfkq9y8zJz5WDw0Iv3B4t+0e+k
W/SLO+RqTzAPKEB+dbkF/zb7apA1zYpwJxL+3C7FjMIqkcYw9+SNETzEBUyxNfTK
qIaMKpNR+7Z66a7mOeq0bKn9AZIE6kxZWyRp0SslepHG7gDQbyW9sfwRTRS7zBtE
WYydhY8xldemQT7Uzowzr4+gEq1aLTN9IBI2fxpNbBuGE3dWpSk3IZj0c9OfPwcY
f+JwBom5SANxi9fa7dALfYo7+R4MpxiPW5UflgHpuE+iTaBprupTkq3042PPa46s
PUUWPgQtDbFzBAMWRNsnhSsMRvrhsLjaldcxRjVY3eBzcV/rODoR7atcM8qbQ3JM
5AWUHYQg9iddX69BRG3tJQtsNpio8WvET7rCzmIqAN1VRg7g7XsasFYSyrTHQn4q
ohr1IZcrdStPFlpDxgWIPyaiEsDLxZss6AsXkTgcnkihX7IraZIlJqf8MDsGSAO4
aTBeyIrIz5cG6Co1vPNmLu/IctdmKSvKBKGENWNk9A8wTeVYcPOqH0wJLAKSJPCo
saPlCHE/8+TJ+j2TdZw9cat3RlOA/9BZqSOTwyKZlrdJfJs79eGQ8dHEquv3FTO3
uZKl422DljHVJeIVl2eQ/ZOrpsk0Vsej6b5xPmCU2YL8cP5Y3aCCZBJqRY4UhjGI
6RJb0dCn8LL8qhZuiKwRg+6OjzhnvWNXkuM0bo3yjjjbsfpPkTNQfE1F2Ci7xFEC
iwAxuRJWIiPIQP89BDv3XBvD/qFkdIfsBLVP8b88WzKkQJLAsSt3FA/Scb5pxxxP
WGmzhxxXL/BQQrrJBIr0EW+StvIgvVRGKlu938sv/CwUR+AyZrMTYlEdbaq6ER43
tm7sqoKTa2RsYCRDD9gqZTG9QZJe5Bcg1TAdHfyItH2SJdI4ZAkV7TwP0cf+xr4I
8mi02Sxn7tLSaIha/ZPg9pyB/xu6YnsIUyp5lqupG4MUk4Z7FpzJ9TvNOFzJ6kOR
KEAPRxBjLCAM0u3VSHKWFtrBJCKQ8i3UgMa8ux8mdzExvp95uCeB8wU4wvYtNBg4
Yrrockqkelhkn0oLB1Y2e0mMIT5Bq2YnToDu5dnzD6FdpCLJXfAYuk8qGcOqUErX
MCzSdcsawi06U79hP9Ez/Ls0or4Ju8BGGOQ4EZYr3TsV+hXtFfpNJ231aMEEsve6
+TB58aO5FQb/sA2DM2bMjh9J9d41JlSjrBxw5S7f5d3tKY6xyuUJG7CEnd4flLYQ
asbH4do1Jp/rjd8WoTfaEF6kJaHXAhSpnr6N0dvYp/+h4ciRP3kVI14Z4cGR/kQl
`protect END_PROTECTED
