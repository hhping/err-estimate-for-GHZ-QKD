`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cH28V69yF2/dkANPZgIfnesvJpygQQdasQiXhtmtIeYs4sZ1eqmICQQeLAL0q04f
HVblxBOOje0hnWaW1Nj57vqGSCwUj+BbItGqlhGVFSI1nx0J15lZnvqX3nnNjCOs
Xi91YkqLjU0wmYAqmvnq3LGshNI17qsfRBIa+xMHpNn7uAqPcHMF09Kf6iNiCbvC
V0MdurvEObjxizZmtUm0iIkJXXKfH941F7/RmWLTcVtCKP6j5JbM2uBw/AkEeZT2
KNAVJBjpWaB0F2i9ICoZLMDIHcQLTIlPq0g6CE4LOhtAYqt2jiQqK6Bm/8L9BP8O
b3/788CyL8KrhpeCEoJPZyVMumfbO7kjSuR71RWHxCJu/bZwfAje8Yx095lSy3K/
BNbWjjsnqD9ITHZFkhanWB5JottAFfFK2NG6IA/aZFHebzATBszyGT1D8pirtn5d
LpcSTGAXqHJkUTiBWdLEG0H5Muc1jGp/K0udxHYgHO/6BO0vSQPRKVYZR3rAbXXN
U/IS+154AeHsPH/0aJHx7oqtsuCU+hL6vhOqxE0bkskUgOWsL/ODegP0yCDrB1S8
nVmYs44TQByfXyGkIUcqL1s4b1Lq6iEpLrkEQ1R3Q5cYshsKv+A2B7OezfwavlGb
9BOUivwvgqGWBqaEZ1DVfmEgfk0prHvXOvR3XkKDJb4+IyOqd+B50LAvOyZXMNnP
YeInHF/LQmC4WqV7PLrhdv3sGuEv0K2+gYf6Xuo3fSjGqiqE07a/Vu1rYl0YIWU7
4AZBWiN05ruexE2wDLAlFzHq9/jyK7tFuV+zbjwjNhTdP3zrwPr6f5vsbslpcF2J
x56tXpTQjW9AJEazuumLyPSu8lX0HtfRaIqZd9hXnu+aCQZjSkZGcjWVjIHQR8qn
oQodkDuJ7+tYrDsPj9RBbD45+MWZ7s0Sbw8vDHtQRjPh5g96TtHthatHXCdf3uVU
nOKZ0t3Bfh3M8AGn8jfn8Q/v9R5NMwnQs9NcJLs0bKyf9RiF4sW4EaUGoSSdd/f6
agpw90F+RQmdrSCCy73rSpwfNV+WZRmG0axxmSuWbXYJpDV+zvy8MRdJlsvSSH4R
I7oPw2txWuu4NxJ0i/5/EUtcmoZzgGWMedNCdc+XhhoWKl1t7gcIP+DcqsG6ynha
pGcAXVRxcoOVPPQAgV+UIiNv+N3a2cqHjXM//GFIOHRm4R268x7Z8ngZ56H9GmII
QUvDFRIHYTyMR1huZDhdWBlFdNtGhJkxS1Be178dXoayqFC7xY9GKujYxIXwY1Np
rCHqgSQ7KJU039kXLYgFHcWpTdpqExWKiLcXgrnukKljQuPw08LxVkd4a4oa7l1o
1t4CVeaxcDBiPGMcnUm9RqGRivT+xazuOsRwlDCB5w6mxV+jM48+b0jGSIa8kJkh
3ozi+Wf2k8OjK8utaKEUtZ00acjvoXd/xsItsB0xuHx5QS3Qua/G6W+ZCLzhIdSx
BT8rXpXxmBPcMoI8mE0abe0Zg5YanxB2C8vaDVrMzGboxaLCcyl2/CWhOvIWsFtX
cGCinInrMLpmlf9bJCbzTBynCLrp6GIEF3gdRhY2WSqB4SBuGAFBAGnqxqkaOrWs
LqWiGg4lgHxq4xuoN95h/cwCeoLwxMMD6Azw/xkJ/XHJX4JdjaLC+CfOhkyF9ysq
7jZkBOt6+Kp4RRvMnX8oRVQfxAZLifN0vvjckDjcAIGQ37YLfxKk2Bt+eR2YNyW0
EAWmMKmiW4i6ibJRQVJuONrNEtQ4Xs+xHXdixYzPkUEWiyPulDy4cxT6swgFt1AL
T27p5dfjTLyyeyD8SKoMa4Rsn9UtiOTYhmKWPT5/RepPxBm5mMthbhMLK5EcUYV9
Gj95XYOzn7ytnVUs7Gf0NWzIpmY+Up3A+TibB+UauBnSeYO2/oubVVDyY8xAs6vC
vUzYdrs4I23pjl+h/LzAHO+3FID///18G5gNY1rrCURLlIimjF5+FKeqZCM89NoI
ROltoPA6AmgUcN+7703bNq7hUtMi6kbzKqTsosecuSog5A7PxLGZSaDnlIg+DnV8
wxHd89kcf5CSiPA7LvuALsRVB4ugBC9LW1nX9zhaIJ/80vPS5pBeqNxD2UFIsskk
`protect END_PROTECTED
