`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmWdwdhPSwb0ZrsuKCKbOwJEOFlq4Gi3YoAoT0Kpony7jCTO9u6uz/aYKsUgjn2i
B2dtdxcXAdG+2QS6Nd4izgNUZdCGPh/AyDmSPsdH035uQFm8uaUUXjlNTMtMMrTB
EL11jYnmGguWlS+hYhKkPUCUuZ3bBZfTfTgbbxqsRK1CwA8hxqRQjg+/T3i1QXVe
exFbbcDfkD8RlHwwirzlVZC+w6kmBJh2bGho4TOppl8DNuPjqB7QQquDIVyJlgHx
fVH8ysmvfKhYVkXZLg14WXms7xw675WtXFbzdC7ws1BirtCzU8WulQd5b6Xci6pZ
MGNPXgUcao8TAkGEmZoiWXs8VsK55RL6y6Y9h0iliWUSopdok2bcnUO6gOwZY7gY
hEs0V3hBnwQY2NEh/Pd4oLVSE0YZlByIDCXybCErgTgNzGgewpugfwWfaDpgZgfe
+MN6cQGt9uENI0lB4AZ7e2dck63y1uw6H+Ie2c9pTfApZF47brN7TsfDH0iuEJ4x
UKoSWWD9M2Jly29l8KruUr84Wd7igED8eYfuI+Sn5lHDaw20Jl4mUCBrvRTmpUfV
fkvUUjh6uKHOWQmNii+6yk7Az0q9Qc7s5kzhGFnpimVkqiX6hVn1Hzuefd74uyYC
p2Zd4xzQdpm+RbPEZuEnFVIixayGJ+IRFD/36L1ZTA0nHmPxoH0DARsJ3Fq7bJsu
oxHQqx/2mN5HuUzxx6oDuHvAFYGSAdm2D0LT0yX64WMj3qAehgIJjnLCFQJ9jGkT
S5Zc9TFB/NPAQLbPVJQT7UVxULLu+66XH7WBotMb0ynz5rWC6ct0dDH4AuStktGL
Etn+m+Lh3jXMBb4QXbIvrMHedS9q1NSjESsO0w8Ny0Gc1f5RUBeIw2oftrDFX7IZ
YrcBto91R5QdiUd/4GM+YtgdbijzygmBPJnh7l1YnnUWZHE/qj10VV1ZrpGcGNR8
CMaagQKF/SVAE2HYlxnPndW9oT0W2PhuQcB3c1HX/hU+uQsAzv2RwtmPi/PpGv4Y
53+fr/HGFi6bLGjF0vs/hCt6RaQuobM/FRgwnWXqi7hK+tWqWZnVXjuqzmbY69D4
pRPJJjZ+/qpYyDZnladFim2ihbsJt0ajl48sy41em9KTaTuuU+VvzW8K8cHDwyVh
3k5d4cARy18awNuVsVzi+orwh04ZceKRWJieHDOEBXFSV87xqHVifUTbLzieuqNY
S7RE6BEG3rBAjmX22D5LGfXig89egNnWLC9YG+2jsJRpEf4V+g3mwE6NptUhrD2P
VKQSkw/+r9tmFdNfsvR5F8fcb0aIX2uj4abknmXD9XczflwLoWF6ZdvULSHyox8S
0P5exOAEJu4T1ZU1FbdbN04GTQztBCiWmVo2GpNXTWCCM3ULmqZ429IpyNomEe0A
pXkaQ78W1EXkzMMTLCj7JqZj0pPwnax5p8NGux39PPQ3z7Oi9cr3uLpw1wcOgXqy
`protect END_PROTECTED
