`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QQFOgpD/RBRKP5Ko7a9PbEK/7f3dbcRMMBDYeNwzAWK0AaBVjkTi9J0oRK0agkTl
9lTCz+TvaAVQA9tnaIGInCqwkaxN0q71I+/zaCkvjOAtI3IUze6oP2nAgmAwXFfe
Ig9EDbAu+LNsFFKHftam5vIAFjAfVXl0rsRzUXowsxuM0MUoo/H0u/1DegpEFA6o
F10Fmbu0G81BLc17svalZXUfUhrOzEOc65UjLtTLf9NuirFp6EqZhvX5t2IKI981
qFllv+z8duBE3l7mXYVCXUyx0Xekibd2kmdxy7G7EF/DfMVh5wS5oLw4qpFgSOHO
wk3FzIDD3E7j8VSPHGfft6xWrHuUkaybce9FSTToZHYFEdavefXMD8r/EDAWSDoc
YWqLWsG74TRmEuvkkh5xtXnc4pfaLhhG8VwD7O5jUGQa8qH3UekSSAPZ/ymgCuM1
josbIx9ZEPDoAP71Ihq2hyO8jDCFd6WxAtEJesnkg+ztVZqunMhmXpMt0181Wu6N
3AWgA8k9KoGbnPFooT4rnPibco7p5liW/KqRYGn1UnwvFr9CSafcEeUI4/XzX4yB
c2ZesDmxhWKqp1UcE6TiJl8L/DJhQBlBWrNeE/VDD4HcckihibXFBUJkCGvZOr5q
pLdY1wLJe1VkPzplZ2fs/6KYPGb8AqeTyAo6TnHwzx1ApHC5IVzlCbhduG4UeZC1
XGGkYZmIg5dUyV2jNFdZXVtRR0OCTZkxR2T5jZsWLAf9eWTpfIVRLKnqmpkewcCj
15gqBe+mnXN2r8aUMP65wUXfwmAoHcVAaELzhfNM0vyirPyT6Q3FcGtksrowZXSs
2/GJ2JBAx6InfI53JCK0VIa6MJjDMlxBgJrZWJBw9g7QxUUG26KAeQehDboo6eY0
6odaL35GNcHSd0fXXSy5kLrp6YXI/W7WUxR5lzVs4tb/3L1WCTpeSju08oe1sRlJ
FrBxBfg8sR8wwWrBHFK6+mdKV7N/azCnkAQE+/5Oz+OqmG4QT3rDNv/qBuOscbtA
dtyCF7BvC57oAg/LJ4Ni+3DKNEOwWQuRX7nfR1iDypRtBf1IH559w4q6a1LabNzK
0eeyEpd4/Y1hqT+31Sg+fMefs3xn2QXA9grjpavwgZyS4ytvNXqjN6iV6Z80GYRI
8kyoJeEUSd4gjLvWqlWUIwghQyKexl6BS1fR6PV0wyuJ2FXtircRvYH4i85aW4tp
uvv7UewL2Tjc18CpMgLeY4+juk5FEzCBrS7fkEKHQgISFQAs688O5oLu1n+Ab4Cj
2dDR7+nP7nArGum/QlxA8lLteUtewMEInxOMNuIf+ZpG7LBLr3WFIr7IYU/Xqdwc
ECOSEuGxWAYbtJn1Ner9+q3LME+fy619+XVM43qtq1WQYfpMC+Vn2KAoUP1p8sOo
bMyA4X8DzTiJPnpJEDA6oUhCaCfg4mrmA76Ux58PLWLNcTtmitSgFAdYesDoWNqn
uCqemn4rc6XqlFw02/2GxwPQVp87VggLf3CNU66d10lmlYbgu7sYC/9UWcWqRFmP
sKiOdIbqfr3/VQK9FxLsDmXff/TqZGQeam4PxLeiK5uiJW2RtGzcQSb0wCcJhD6h
5sLfyJrg88HIb7+6yVVwZ0nwu5UXZ7Bek/ARjbEzNMHf0CJVcs2d0EYCPKnPx7rX
sKGZu4DUERchUheaZzUQXuJFhwbp1P3IwOVYnnMYHQ6NNcLhA6V0bKqDwfCc+Cdo
F64Jr007F4Ry12OaXxmKW7KCLLSJr+jsISbwQbgc5asUNwlbyvtp4Rgk7W3oSt5S
a55ciNGr0iRUbv7w90U27zkQeRMMoHm54DykZCSekbnJ3JyFyakUo75mNxxIER3b
Gr0mgu3u2SmXIJGzcytmtRj0ZfDumu+G/Yt0FJ6lH5Cn7c8akD8xyVwIbWDQdpod
bL1VVt/+3yNIWYI+WKgG3WCHrYVXTeuyd2g0suoDu9tN3wP26vAOIWrIwXkGWxI1
sXiHUTQI/In4G60sqt8Lgg==
`protect END_PROTECTED
