`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJENtQjVxuPWYoz86E3D/XQstBWHdfnr8Yaj5msufNvDz/GN+9LSex18ZLrdvg4s
HVcttg0v+rbHrB3n6e60+GAhhkIi7COYe3FgG30ZlFDDivSvLLaki9shEqx/Eluf
QUUB6EJ+kQULmGdnhNjIJrfsGcvlu50K/smhp50JzLyCgW8XyS6F6ug4AojRqf3R
yLdS3KBRza32pme/BwfggAOPNARyYw3N3IaGeFjx66u2qymmhAKjuL2fovMh40+G
utu7g4iWg9J1xc6Xokn43DBQx5GSdyXt8pal6xnyTXcaUkVmMzoE7imM8ulnmVWJ
ql3cUYS9EBXW3LFvfUw9nX8pdYP5LkYKtjFsdGvuwVPVeyMk+OMzhjZicx327yb/
s7wpALZZE33Scf8XXCrl0C762Ct6+lGoNnJaNRef4VgQyNxzGssEHWBQut+Qrl6B
fGZNEsNkNJqR3xFuSLneKObWsl0bhnK6qbJNHMJMH/3sVMSHzXvML/LgpACgtaHM
qG48SwaAgKI2IHEM9wY2zgDlt/UNhx78QUEB/YIhCXdFnrQ1uRomsCi4h7JoEHy3
F+qqlDtxbgj/0zH5uUCRhMORk3v8IuJtAk+8rKqbBNQ45RUO2x+CkkzeHBSXVmOt
ZUjFGtEUeMSfogOe7qM/2msKnFSiJwCfX6vTu9Bbzw+i2KYaz7Qv6s4nrwP8fgJU
O1SswfeaNhCWG+yx3D1Y1Zx3gjWl0zSSfA+HTTMsAPDWhLu/+IGTq6aDsctgkOAy
wdy4Wx4la9sIYnt4dYXOnIFyjVA9Yyjo3w/tpM6SjIsWSRHny01iEA3/ufgNg7e0
w9weDB/3z4OsdhsdLR/KePsPU6uAJCPuoyOIWeoM3LQ6MF1UKWFFdXBxn1xloQev
Hn4oN3KD5KDA+NFJeoBcvwEtGekNXtYY3ezlbIwt8iNAW12IXfqBUj+lS1f9ggZx
NtfH869vefJqpbG5TOCHq1bPsBDe1Vi8hbfGgYt8wdWq2PidkQ2EQAbWo8nlepXa
42bnR3gfInQWj2EP9i0DAa1MrZZP2qjdfCL8ruISGgb2dDyApIg2Hisf2ifOGB4W
7NGnquK82i7ugY9JPo90aSkZtH0c506xXpytKPt5AiBhLNtsAMWA0U9HEbaul+kh
jlgkZBBPrwyL7pbsnHVcYQ0W3a1ycrnQ8rMB1z1+j5xsP2rG8J+CG22Rz6BhVFIG
Hmc170mpT1mKgClKqJa/ReLZ2udQiAtMk2MFVEndVKcoAEx/5oVfG466bBcRkRcx
+IfxxeIEEJqbW6YGCbHjmmW5TiJEIGDfsS6k7yqMP5pbReMegu1TeIVvD0ZxwcPY
jQMFVmQyU6hzeJd2PD/PFZL6BsPgHBqVwvFwi6aQ4uyuEjy4CZaK7UqJyldN1yW5
cq0WZxva8Me3FP4nXhFQCzktoc8m92c3NZUBrRds0fkHbtuCBTAQrxw8CuGkBfGQ
oEPNfff7mh32pNf7XCm6GyEV4LQgMnbC8bRpLqPP2suEH74C2aSg8y+G24AXl9Ry
F9SItIOQCwPq/CaLkOfTJ6mR9TVByezwIl3yxzj1AXAhCqhxlHFY/nRg16SOQCll
90EevNYaOv7CW60GM15/Upkxf78T01cFdwxekuQ7H32W0xNmApKMqjQn9iF4CfL1
uCJDJeTDRgBGSDj+rLPzkxwZzjf9vS+xQx+tK8IhcZcMinJovGAUrldARErvowKY
ZlQunRqgbd/Du2z+HBdwNpW5Nmcu3x+RzMe8+/NwWBIfSMZSGv+Ra4/3mJIYk2Tk
zNEfIfzq4opX5b8D2P8mov9i5RsspSQ+ADlVA0tIx22bq7p5Z1lwYaY6G9AeQN2e
04AeugNm3JuZV3o3H0rrzT41s6hSALhezjO0q2RUT+vq/V7l3MwE0Qn7eo5F9Nin
GocJMiv4VJT9CqXPyJ4bunCMXiV6Sv84xe8+tFY1kPN0g4gW8+IiMyWWFh142ZGv
rpunl47wOWd0yYgwjeMi+YS9a89UKEksvDrsMPt/y5aGZucho+7iaxuXwzeRACXS
vfN8OZBd9cP0D6ZmVheGdTOMTi5rnaD+DSpBfd3MwiS9tYGPbEZT/xsSMa6A3+tI
XccY5OSxfdFpkmma699m6BOyEgSrgVVOv0jTet25xlGbBQqPDsar/UFfc5cwD/Ij
KC9yn59+QQn8IImrEci4JQ0ebG+Prvg78VEIEKYvAaQB6oEo00WOxAcZMICI0Axh
z/4XfvjANXDcH9dx66TNMm9AQeqb6NQM6Sd9zQhPVQlquuZagBu9+9IttMlHgkRR
WWWquFN0HpgRvLrKgR4jtwyl7Jueh/YZCY71XUAptxLZvJ2s79CES6O0MsrDww5w
8XQC6n7Aygrq8WnF4AhMgr3pHWmPob0SFfV4OuHDW4jxaZCEzK7BVq3btX9gI8xw
enY8BnTSv/Ix0OHPcGHmJPXB8ijfPf4OLvA8YldcBSJeWkoK+Oto6vc1Sc1Q/YOf
IvZeDP7mten5X5Ux/SyhPMfHiuhmLF+BdciH+4mR2P2KgbXswX/k9h/hYuHtQEBJ
12UjF2EVo0HvJIhXhCeSYEzldsZxczQcxoPRD5aJ65vejdM/I0Kv1fcxVHT33Rmf
G8Kf4LRNwlAIAP6Aw2nrVZhM+BkIIvgkxf01AREo1HnW3ohnliHBuf7Af92h9KON
Cju0YAKjhPGz3tY3n+2n6VCXFrQsvuzRk/MdIx8A0y0KXqSz7j0Pj2X+eGDyu6FF
T+9T9lAdqPoAaN7iaHE1CglfeMFPH2VIl5hT++RMUOBG+lcBzIH+9Pjk0j9KN6oX
upJEbrByfjZHvvR6EK4FgWBZKDF/16r6Z9zjqsv83dHBKkCG8MioJ/vuO/nRyHZA
WweQt5cPwlveQVnc6mQPCeGntsYiRwY/AiWKZsEzNYQsamXa1nBIPB99ZCWDvgs4
CjCTq476jlkckyH+yu/8U0pR1ettmXyTyleZRESwdAYpX05C62SbgfQ+VN9r4RH3
eTpL3m4TqjETIphL2FNVG6n0KJpWSR7Jq0pxavcmfhNHUX88MR7+IG+nqI5b23p6
ytGBdZi8DcZCHBfpqlkxa95o/+ryt3MlFyA8pnxtuvPX0usCihlqHuAiMJbIMhfE
p6fXHAI1sEuVzxAy8jhIC6qQ0xQrGxQmYrWlrzJH/ghxijrBiG7IRpuIZsj9dtCb
ikIp95r0Dx5frWkC/eVIFg==
`protect END_PROTECTED
