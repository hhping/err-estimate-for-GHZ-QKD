`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylEVYJfEtjGRTH9dsbDU86rIAitSqPhsxfxaDBBfHsEQ4fp8u6YxCOSRzzdJRzar
gTl6LjLhBIp3YWQvXX9wHYhubMRFs/4k0Ajz8LXOFX7TwS6mzqTdp3KRE6/CtgSj
RKUIQ533n9Clm8P2V0vEgpYZpvWiEGITEDBZydFsCnt3bbGAdodUzeMIwTqXiECm
CuN/7XUgCfAh9KYxU9Ldmr6xOBdmk6pCVYY88fmnDvKifuPWzkSnkg4XukqevvjG
GT/O80MH1qVQEH6Ix/tbk0AVf3f9xC9g+mnv0UH5qzURgeBUX/+VIyrJS1IOOTdA
T5pz57PV2X/s5KfmvKQ6ORdDlsJ8pJl+OuLb8orkJmjKj8nnFtU1N2BOnCoVsRGN
hjEUBJ12rEeKDo3nUr4HrIdi/R3DuWR2tT1kE6oR8e6EO1yIAbBYj44FfR88LK9j
Vgimvgvz4K5+ZWIVZ58AZmMbIz4GTgX3YlF8gY5bEtY1OReJEfqGh1a/T9h/M0ar
ocIASwvzeOZofeI34QLOt4JBdGJI8o29QuOdDDxHX988mwzr7wnlKxoEYXMmEiPq
1noXsPfCPWU97PYfNOPoPnT5aTabOq286MufUfM16utZUz++AwtPTFQDE3cQBtda
61IWXgvLptRLVKYyZpOS3LYhDVOgwbEitWyugWAjS4LculxkaTiiEJPulq6/zZZz
7fGUgTAsn+voLZ2lBK2wnaO5qMbjgkz+1/aPAjXYvD4Heog+bYwbHcugG/uL+/mN
r2WF5pZJ8tfmXZnHJVA4SVIYxjSa1bDCO+B/C3616iimze1EJyQDhdbJ5GSbkzk2
upjuyo/Qb4Ormpg9z9X4LJRCjVknXNZLLbD/rIEWbQUDasAwjNEQgnLewI5Stcx1
zqn4RB6uS7MZ0pX3D72dGhhp/pxWNXBHETIEt2UCQfmFLAeul8TIs6fAzsubWX+J
aeghjqQYlzUC2Lw1fLoEr4PXjRYqUkgyaWPmly3ZGTG98NugmjmhUKtMC895nHsa
ra8its2tuSficz9KKHDyPW8uzSGMTKUkeLdianWyHd5+PMD5ixNUUDcvjrVABSfb
HHiZCRPaGNw2BaDDxxJ3MNEs2gyBgeZePQllEOzyIlG8ysj+rX8qvIXjBX3K+mes
BrJBpos+FShK5lpvgXq5NiHyttaClZcQ0JMxkGyAOkaRcYE386cm9mfFmZBMCe4g
0/L/A9JIyYW7NrOTOUzbpUQqz8K08ipT1AeAkbZFOLUR/eSSgvIcpyB3se4VFPVP
MFQqcdymScSWs7jRH7zreYo/KW150e6xb4kre/c73jEiM73o18DlwRSaYrIpgZxS
JpwC7OCKS2cEUVLOWY6Cyp9pR8sFQ+n5/vKoFpLuARq3PX3jVIMWZgCUZLw07rLn
T4YmZNf2ED3H8YUzZUPgYkrd6eIsNcEGBSuD+Y4fmPNFF7MPWrvjPY18ysXsqjnb
n2YJorQ/cgjmK70BgWHP43+6gPZq5ontYwWSn6MHwa90BWyT3Yt601SucNojJ3MF
COfpneOyjHqkVYDmeQTPynmlAjMMF4zYRtNLFhRaaDBaT+/m6TnQpr8tz+olU9o8
UnAc3B5RTzR/U7NDU2SkzQn0oAtB6z4pLNzdYA8Vpt2Vhrzo4wJDM6sImibdJNJE
7njs4F8t5R+w/kz/HjtM4QraWYiToJ5iz5BtRuml3cBHy0FuszfbgehXuezAPSs+
CxJeHI9rljqHb57XMsEdcAiL/yDQ91km9O8FhKu+cyxayeSiuStOnmI8/x7UlZpD
dqKiT15uvo7xDcVLIFZ6H8j4dG6JEHR3Z1xBwjHxTFskSMAZjaOj+NhToWdAphGO
3J9HFcte5WedLIGUWI4keunIS8ZaP0blsCNmtO9o/rctoAV5Og6gZrJI/ZUljlsw
E9FwoKURLw8I91pSaVeOtBhid+Nyla11CS83UoI4zmkDKuHlsplthyZhmhCMXTr+
GRjd2kwaFrRPpR/1ija0a+kqU+N8bErdYZTyso48PdKN/PbpetSaT/CUZMqtnD+E
N5utJQF5n+F2kLXReAmYVm+BUtQltVBcI3IIltpa5EJ8GtJ6ANZiBjDKxJi/fYOk
0+2CZBgRRv2Ckjm8jOfrZSVeaILevsJwilwKYiOYThlvxV+4ODUQ7dvAkq15x2Nk
wo81M7+fYBQ/S01XBSblxhXzvg305w9o9SaoDA5eKf8vRaEZEuQGPTBImoSghMwE
IDA9fn7bxvgA4epDrRzWAjPiPO1RDQDf0GLOF/iIH2U96Mk8BvYXqFhv9ksgIA7w
/8+loHHmZdh7cgOnV7e0EN6i2Rq8xmZOHC+HbNE/MzKXBdjSVuzZIqBwXWj273Hd
TMVtkiW6RywZmczU0spb5+u0QSjh7oFYqTe3OBgr9Ni6WVfxezKFD3qT/UuJ/lsz
Bt1xOJF1KIEKQs5a713Gppg0/yDEXaefgVD/D8Wzoc7KqjyjgHejkU/5/6RyDSqO
UH3KQYUOILmnCgptA8/820ZM5CMpTC1JY6KkdO/EXtMTgHhk+F/qjBHehVinC62C
lehkGzi9Q3MSSxRMICwgB0dVttRaqsqiouGQQmIoefqWKiBOl/9Aqe4HvLLocFhY
pHMPtUr9uiaBZ73VBYHG5ZIp3zF9x6GbyfiMo3M8FrBg/QlyIwrbhblJxaKVO8/L
QVoaBatgFpKdSg6uos5BkpAsco3wpP2+5T9JmuRAhNSkzhfCMuyb6c7xVnGI20Ye
CNnA6lbWEWt6a9DnHRbl1Q+RJpi9LY/TWUhNtz7k+bC2eLaeCyrdKnUxJPVkwDvM
NMEOK6F/G1Btg2DSG24RkdfBYWt2l1JhdS4nV9Jt+RNbdXKUQXEGHK4lQRAnQuMz
WkL4+3l82CV/DepqYYAkBdOiUYv/XPzxGImqtIy1U5hqrU8Q9OUOCw0MfoBfzYqb
JDJuus0G+mxx3PgDh3d9GMg7cQxv1F3GCZ26oGzF4DMK/dI4Z0gHq4c3LGCvuX0x
ekiDTWlwouZgGSQikgvJ6aKoPm9miyzFunwqbL8ZZafHrmMTCqJkq2bcxRPr/40i
zReKcIFiyabxK0w7dDzhSC/IJnJHLn1HxYu4RaWQsQD6ZvIIy2BjqFa55ZjBL3va
HKyTFlPjF6RrSW70zuzNQDQtOq1Val6S/+6DxKzBCq9SGDK6n+tRnda160XcGDcy
olEZj7y/QkP7LBEC2nuK9n4cMVswWG0XjJS/W8fjg6T91XVFkEj3xtD8wDBVrIjA
mxaXlPBhlT9qLirhttutu77wXdX8Y34bGOmgKV/d3j40xUpdVYDiStcsRlvCfOgc
kvXa1scmW0ToAO7OzDWFxavi3gujn/0658PjVEgBYQIS2+Fw3kDeZlKJXq17tglv
+3Uij1hfOLJPSkDCm8T4Fp1dSSgfnaYMjtFkZcM/opGlcd21OQqUhGMWt5C/OpmK
/gQ6OMuRtc1fUrlPoCYIUKT+sba+A0y+csMvZTrVmGUke9HwzD6s6y6mZ4OJenem
r7z9EHeWgiMNHb/plKSN6lkxePtg7dLY8ifXQN3A81OMmctWdzJzewgIMD9pUY4R
AgyvNGlC5/fnuK818aDbiTqRGtNhsm2cffWLrRWK5m3OTPtbkMYOhj7M1JYSNOcN
pn7dGohwv3wIojA2XMZFoip7TrqUN3WBbtLbmMbDNhlRxOasUWHu1BuiTyxyMJFI
5yuvQBA7hdQhJEaohD9wUpte1CbdDMsNniml+fJO9xUrywbVBqeUwHJFVffvMJdu
mBvKO6HAWHs51Ds8USuCsgWTI0m4poZ1/GeZDkEG6tVAa8RKDyKt8bRCa0+KLd/F
mdVKruu4EUN1MOHK/p9XYot/utcQ0WGtmbB/NO8iVUJCHK4uT+WBjPi+XbrXU1Px
cnABNYQGJEWsdukIpx4kEWWkefYGmPQhwVuL1/eFkZP4WMrmIzOt4NVbY2KQRYqm
mdeEiOhjwGDHFc1C690n67JpM3x1g2gBqQC4AV0SevgDNTIHPiYCKiFSP4m5gd8E
wTsmWhsdnk6Mj814P2LF1tj1pCBDfD5Bc+bOi5mGxkQI0QJrYK1tHC6REe0qFE/H
7GeLWfDzkYDC+d9Aa8jFm9XucBhe9Ew2bvS5PnJ8RLmpyrN/QAMlUqy0hP5021Vq
i+su9DBoEFdPGSWxI6aLHQwlhgr1hfWHfqUNIsoAVF60Mx5sfU2Js0y00DWCKoK6
u8wG7G16cE8cD0DW1EqJOYVCNOO7/GpJ2DVTFuwiiA2bMuQPLkr7NTVvsdtbHj0t
r2G2okgkPR3lmtPFMrH27rta7NYTJ3rPFBTfi2tri9CBvCMQ2RRVmb/RVOCjN5Bh
05VwRDfM9qxKJYK2FOgPc0Bh5mY6SWFFxHA9iafkeQHcrRbXCUu7dzDinhgr2KgC
vIYJq7jNUIQS9Y9s+ze6c+Ex1EuVU9H5W51DtDRLHZsdlSLJ2sYmhyk/Vit54el4
8gDG1/ioIRNIqZt++chjy7dEYEqqWvcupY//9G5hfl+y5kgICSdfpUgbA8dGHky+
HCYZartZFRs2s1vO2J7cDVn4CJUVgi1mX75jT0HrnF7JPMquxbQ2qJZGzdh2JSdt
qSkCu2pvR/YGcDnCYVPBx2fQ5u5luDkuIjXNU1qU5WNlIU6+ORnlQGbuGrGM53Cx
KUJ1Uv9Y7voQTaPs+wp8di+oixoAJ3OZpyaSWL4IiP9vP44hXCqepRJGUMo76HX5
rF34TYUXS8JwGJxwP0proUHxEtTD9ECDvuC8vqNtYQh7XJbuUmvwXUrdvSGKDXq0
FyDAQvWOrkEThFvBfJIgR5ToYfLjzsWhZPGfZt4BaLF37DiBT36XkiuDqzxs1GKq
3ptVYoIgRu8pH1D+jKc5VMcnMNi0jlK1ve78fS+iCnL30VdKw5wXJVVwO04ErPGr
yElk75rXL3yn2936mHiG9S+bfj7U4dlcjlQHRnqEtZkGjPzQJssy1+A4AKnUgG++
VBc07tBsAnE3W6GUl506NitGmj9pKf3dmOxf2EuOMpyRJpce5MaLGbW34osOp5YD
ce0y1cjVBM3Fb218gKhcsSGhpCdGq1S22iUuP5X46q7dFJTxR6xfl+f9elTK8dOh
IkRK3N7C/UzxV2YrG9CMvpFNx2q89DZ1UTWQz/HOkeHbC1EXcbQWkPaCUKIkSPEg
UakRSPzRFTti0bGDUoqVABqLtAuUaoTMxp/fVYynI2HgU4psYFt48daglf3sFgcK
oB5WNg19wfIzdPdYJkWeDGrUp/IYDB676RPH4/WS3lvZ/6S0k8fQdvajrfjvn0xH
uZOf7zglWSk4La3/R7d122ul+WHtpWkXdxdzqSV6A/jxCE5R3ch4xPEjHg6Qydm3
vE2+Lmn+UkTC8Kd6z1q4Ow6mP4ZM5hzB2WquRchnrniKsPiPJUDWm/WlKED4nVWF
AerPbb1Ew0TAV65vWSJBA30o81n97Tk8Z4s4HmnVGa3+HK68m+gCzKeldxYFJt9S
cr3dKo9F2koICvhL+v3iHc6NLfay+jCC+YV6eA5Qb+UC11jKz7sYqQGYJGEePIg6
8+M3P6ICi7ZOCiEAWiiJHxwjPGOoWBR7k30xz2zZfSnXHU4zeIS+yhwJtCZP151M
zicQhwENCMTEGC7luKVBt/WxYwPnKvaDLflt+/0Cv9fQiFaSx8C0MMGOB8/HaCu+
oMgGnZFQXxUtq4/0Ln14V2oyWAjzZUtr3yT9LPWO9yizltaOFghjPJQzsTqP9rFN
OA1xUr60tRcU+S5Sp8ZV9yxJegmXvvjzZHvTZmo0/8L2LQLSBwMOlufw+cwziQkH
lvj6IYGfRog45QUthR/ULJZ2Y0B2JHOkNoKscXun94Zxa18lsOR+UjWwW+pxKAju
7yyjFKvmGPEE7iKmELA26XhlCX9FYOxqxwnFEg3qoMhiO75fr3ShmxnHXM42P/4o
e/vWpDIM/7bGbcnOMm1VVInALEZ/j+IWkjxdcN0FiuSduWNaVLfaA3zRW3Cx4cbr
292nty3Ka32lf5KO0kQoHPhKwrAp3dFT8CvUZtyJ0OmQwlE3kqcEPMJX2J9HWwHo
5Gc55f2PgZZl8EGrXIQVMujX9l1r/9TePv5bfDEEKEt+zlUucfu/ZS/1Zv8+Qwxo
H4nmdIxU6YGVlif6JzIMMEXolmg0dWcpHANgfpvF6NlgKGLb38KKaUJc7pjrmLxj
miqzrU2HJ+U1MQFj062BlDpfpNVmsicTUJWmsU7YMS6nBYk2KzlyPAg1R8/2yQpp
3ObCavLZpIaXyaBoA3rSVk2NzhIU7w/enR9bmwbp53D48LT4tuNpynRKdlGx6Qgb
3zdbo3KRcvm39RsTrG8l1gljvf+rXlRLfZbLnVTl1m2ZYHfTe/s5M7fpVDcmefdv
7UcUjo+BiqbAuTP6MZ7uwPymuC2qHJdZPRH/EiXKw4jObYxZC0dc1ZJdIXdBnAFd
bpCee055zcSG5RnS3uV7A6wyKNd56WGXkzzWxVQPT8uyILAq8BMlI3m3fek/Fg0g
DlXNDNb5lQX5EN6bpSWYmEIskaY9qR/8nkoCEq85QKefnk5a0VumkRbNeyv2ogK/
`protect END_PROTECTED
