`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YuQ0QGkbHg3jR2UuiXve1Odgvlj1WEEF6QeeWh/DC+J+/C0hvprgSocz8Brqa7bH
/SUKS+eRtZ4+4fCp9FYonBrW6SFXnee22ENg77Oom0/kc6TnHq82OIS1FGWmQwT4
599r8BIlSbRR29r9K/7nltwKqqqe3d1JW37Z6TVfy5fPZPS1qBk5Hf8V6rRjXK8g
CFIe6YcxKkIzk64J9qfIDQdJG2wnVHlHen3sCHq/X8D5JxkVs/iX6P23H3k2pPPv
Aygv0w1vnKm2/+dU9ZFvVOZlMxQEnOPH7jFJu+pooNZVDtmwcYI6hxX8j2HTWUas
0pzpOSrmts5puz9VTO6SE84v1v+P2sTzwpkYmZtiM2nIVi7mxuDBG/wV5haDdffp
mADShZ7wVI1rl+053rzZWg==
`protect END_PROTECTED
