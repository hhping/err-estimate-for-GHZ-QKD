`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXW0z+xvs1aPz/Eh3KIEUUFwqG/Cw2VEe5kMgLYQJcgcQto1Io+1RVO16ffbUh0W
4UifRIUTbMn1UfhSgfHtwsmWVm9IkxXmDVKluJw6V9RvViwr7zXhHhu0+jyncoYs
kA97oCr2Tbr3Lvxk4JMJO1Tlzf9dOjXTkSo8pzCXJiAsVIaiInM41h1K/1vMtiLN
CtfZeqFT/VxO0c2QOQN8dsewp/FCoIMGHh/CcFtMT08eEQGjxP9L87vBOwFw5+7J
4Xiyx/RRuHTUYeUkDuz37I+d+jIqPEeEPJ7ii2fi2fmjrwsRHgAn1LX6NwSqIXKE
9wwmBiM0c6lF5yJJoBQIoN7Y1VSJan7CTYMp5nbIMM24PvuAqhXJfu4scOKKb4qw
/HE2AvUVF47MgpPjlxlfoXHcIhhXoLNH1/jt9aDp6kgGV1h8te0J58Z2ZL/2j0Zp
I/EgdFH6lF1e5OTuiqkooFWYQRvgbLospFQhpI8IlfNTxJwejyi7CVvIf+a0D0qp
W6kYOD3mukB8cqw+cERHqFzLV6QmO2kJbgVMdwCmNvAGkVzCEnxb2WG7iqSbONEx
ppLQLmdaBAsOYEr6pyF7ZI4DcQZsxF5Ncw0RBjn91B5hnyxrr3zcaYdQ+OnMR7Yd
knPkM2DKOj1cFSEOfxsy+aFH9zGS+3hKv+PAQ47+HuKTQf4BBPlPUBORKxgKHnny
ADK68HsHtj0+6DsD0T8jho+LEzESi+4i0jI6FjCqipy/3qSuz/b4UGzXXMN2OKlU
qYqIFzSy9zObcfHJvkEECZfX7DXJeNqwIyHc0PEnVUuxaZKyYXFcx0nQIsY6thYE
A9Fed+Y6UUSAtMW4r23kwnjZxn/hqeWgy1eNj+CARR2gyD/inoOiZaMay5hEV1bd
WwgDRBGWNVeuml1RIJehSLLPPcWUYiAiHem+O9c+SzUMYlgs55M9BIYh75zr8j4J
/5g9RiV90ECijGfaqlykXphv1H1VKfLmfLMMe1jfMeC6AxqaqXY9F8F1jjQ3ESSH
NcbgFi6b+afsiucqtkRKa15RPgL2DcCO6qpfixZFTzu04IexEexHHfpaqdUmDcMs
JXjKtXzydSmFS2AJKS35rpLg8ZGtsIx3pUe1MWhRDozcpdtZDetibhc7e7OG9qII
EcpmFWAp5lV2RThp5PM3l65Nn6j/TMo4gBB7SueE7kd/DgTKjy5zxWetsv8HQer1
b9RiUrSMwD6g56Y+XTd9h+f1eSv28jny7+Zk5IL999OeuwtkFi/YU6AVwMqu0KgB
BVWKDC+xeVlWbZtGgrFB8JLzlz2UTtOtZgMNuxaOnakFjnK0bNHj+Z/jBfxCO/lD
R48ZkxqNv8Uo4H8JV55ot2E2bGwkXVfH0ulztCTU2HjzjTup2JuGnkQAWAgq/zdY
hI82xfw3YvmHzQXvPCGqAX3FD9F1XUGYb6fXJNmcm0Y9kNMPjTf3gKX4co33IEZW
NADOuPRfKHR+uoMVH8mipQyfyOAqMXdjSZ4IZVB9T8CbP2qTorNO3N96PXVP/7GR
ZrPM5+h6U3oOLA8EsyGPDldRCM1BIrkIkibyvRfWM8+jgoB/5ukCHPFEZvI46F8I
yqRzBDt0MGiAIydC7sOLEOfcxuvqw1xD/kHa+cB74/DTO/OTxtWEBXUHsQr8RZ8e
S7u0SePntu+TLEl7hv4W0O7OnuXtMraP2cPYTeeVZ5+rp819pmsc3EOA2pSQVkJI
jZJxvSvN3YQ0O0E9z3j3fbs9HEGaH9ktezztzIFFvt/vjAKOCMtCLierZo0wpIAk
JOiP8oDUM+zs8NdBF6BNasoddv1brchEuonQ8z6jKr+APwNi9KTsZiiDIn8FspOr
g8PfeAIOrN5jppx3WtmOMq4QGbF945a8dl+tLSGeOleRKWzqXIbgSQSDz+RXeKIW
RDln8smYmeTEwptE+BRUr/vbdzRb3H3BqqaxHL0gYD7fdeBpTzYoviX36+uIqiak
Q/E+wHtc0NkxO8iPe4Jf2f8CYGZALZHLN08XHkI3PZdSJugRAB2QY1ksfaxnakDb
MFMmlGLgwIGc81k0lksTxSH0KELQU4DmBelCOxwVKWz8wqNscAX5zIFcPulcWb37
Wj5eoRaFMnlpwL3LTim0bTYdt4ro9lqNXItm84VJh/ybFvvNG9Sk/3jk4Hd9BgCv
3L1hhjUESO+Gcy9zZbzABoo1FjABC7V6FDGj8v5wkGXzUA79jHg1arN4fmc5vdMX
fTl4MB5OHIa/GpM7TRISiMXnxQTfLB4LEciqp/MxiYDoFH6pzaF77hflS1LH/A0u
ToCFpgR3EimF3q5uOpRauC6xv8O9IbK2HvMqQq4465LL2Anf14hJryk4nMImqWOD
G609XXPYc8JOlswThHDKAiexKTcbSket4+YkIkOlk8z7Ekd43MBv5RrIMkFtHWC7
WIcEzHmZShUF+3gFt4tFeRrKUh1eLjvBJzS117PlN4x6kusy5cZ9Tu3R14hsgDP1
2tUUF1h9m9+TYNU1dMsYuD/pB0jD76INCpUHeEO/vrrw2ssSk5Ok+B6mqtvNpUcx
`protect END_PROTECTED
