`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9lR/fajRzYyXIH9Gj42oxrGj104dv7nAVnyMCHqV7euCq+LbT20waqBtwng8bHn
WUnayM6e5cTu8EKVwHcTUu5uDBzhK7YxwZwm0HwRd/z/isfE1zAIRgE0DE4ewNHp
2IcpC+g9nm+3dtjMXCG85t+oDL73xilDH8v/F3e9OGU+cTBNr16TcPWJT2G2Lzun
/VUcjBqMX6+YVKvfEEdzmp9QbwaL4TKHzMvm1eadmGf6G8q7LB6BAI2vUHopF9Q+
9yuZ2cWoatwGq8/lYB54GlYU2kXUUeKVXJ4aMEk/WgPH9gDXVmxIu3o+8Qq0KAZE
LUZs52qI8yE5m6SxLDuAwAF5Wj42+iutF/1Qt2xBM1k08fYb0XG3CgnJOREtmr07
ZriJ8ym9oQv79FW1qPe2ZarMmoiMGN9qe5yrv7eH7l14xjGhSqMHT32G63LoG5n/
ExbfOL8m8at6H1xolYrWuTmAsuek2jpac1osE9oiZrqTHskzBT0Keddi04pRmJvQ
UeqMSgt7wdtKEzqMWEeVO+nyXc8rAZEUA3NyyH+HAzp/atTt/iyuPHALQxXnGy+O
fPJwA9mC3YU/J9gE4HtgIdXhWR9GTYayLPaw9gYACPX7Ck2WlA9dGLaPiyw7R20P
KsByPfDQeVuD1PaaRSS9IDp4CaSLD390NX3y4t5Xdrjc/CcvIDLEV5tX0eUV0bhJ
sClIHV4kRA/FfR+CA/XEkQsSWa5qY/QiRA92iFsudUBLW3Hdfu5Qybwrh9FeWFR1
6uFx1PTmCGzcOiMASkXw0A==
`protect END_PROTECTED
