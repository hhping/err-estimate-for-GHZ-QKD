`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yVKpwiixlB/uI3nZUUm4v1kedK2mq5TejZ6+IYj28OipnlwMVw3UE1E74p2gJm1t
XXG+zJ25jvVvscTTiUGCj4+DCu5BlWxAoH4+uIGWz47Xf3XUb6WVhLDB0r9ApyB8
UoQ2bNCUX24shINKDdu5+NNWknL+JF36gIDv/A/y9ffolLzYzxfW6Th8HGoF4zUg
QgRivDV5YPZGFNVjSW+t3/X5/Czb3+ZKtUMM/8KxO3ZSWOzYVj0SyrJYwkLH6XGY
3Bri9jaMDJqaQ8gZtkj7mx/Li4Vt5xa4GJpJrljkPuA0HH3U12kSJFsYwepZOj/k
7CQyTfeZafPE4ujjEmE3BA9V2XWklW9vA8MAJG7jmW/hEU3JaTzgjpslEGWkIzV1
LMK5RF+GswNrElM8I4T90k0pWbAulJ+gqnyvOkx+cg4GbFjefQfiohfU3rwwv9sI
zw1s2I//lBywIs31KMeqe1sRjEC7vGA9pIY9AO+JZclUTzbG+75IInk4FJrxSFTL
shH7xwqCxNZlc5LrEc7pVKxpcebm5NcWT+uxNuEem2CvAORU1K0y03Uq1DJ14fBL
Da9WHuWt0gOL6FEc3qKTBqIo0Xw092JgU4o00sVJwSz0vZ+OlpJqHWeomHvIWsGb
OPi/gMdSi+8op0oao75qtEbzajffswsxGa/Jd9BylA2BN15/LUESKCe3fzQ7iBJ2
DuV8KspaSqXUa0Ox9mjHjH3sUkg+JOXRdNA9c6+aDwpUwtWIp5LiwupRvUroRS0H
6yDlMKdT+Gyx2XjqY7WqS+jGGueUNwKqLKUBCx5h/zU=
`protect END_PROTECTED
