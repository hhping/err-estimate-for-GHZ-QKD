`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rT1fRFbkUb3hfVZEFcP0WdBGXrQJwnNjHkjMksDdLtUEJfkVGWixx5zZHgIsmlvK
beie6hSgYw/LVK9uaX7eQb34Kgq1n9jEvgTUbqI4Tq5C3mks5GC9tG2BlRNZyrjz
+IPY1cl+AGHKrYiXEG7RxJu9gTs9t8b2JwX/96IbkCbcReO5OS+6Oo+F7T00IL0k
ieicHIEbembCWKMormzXS93s/Jxo5wX32H58+8lMoLwydmSSfW4g8U5uiS6HQWKo
+PGPCHrHKpuOrzWrG0i1VhX0NdYP32+E2UkAv0rTpO6qd8ohVnDDM8iGl2T8DoVB
yuTfq6xUTEqDV5hvc3BagVSMxRY7emz1mjLpjVEbJ8uSfKc/5PP2uS/S4RWufwf6
B9mtg0Li6LdFvcQedqCMe1cCFtkkYpw7/Pf3ZyHZE7ADXXXu9bgC1TDLwt38KVp7
JkMFmioNMeOqw2K9iBwPT05ZSfBFrlaWFrojbd5YrZmeHVxDYA8OYDeOLW8g75ip
Cwn+c/puAqpYeC3GLGwjHZy9vqokQvHxqEIWCzX+l3cUNwxSC+THJZ+Feiwdbi28
DfnN5KJ73XJ2uxUeBt58+pFRXfCJFjFZkjUMH7GL20ECc3XI/xjzhzY3y42Il0+i
vBciL0lpUJaDpdlpq146e0dqvWFEZRzbdQXvyZPTgUlompTBAUFzt1KHjA2Yp8Pz
a97VYqVBHtKjZyMEbZJYe1dsWZq7Ha44pRlYw7MAOEcMpwTXwcP4ODRg/yBT34aN
lIpdLWFhP+8VBIu66EtGNZ9Ehg7DFnOzVKJxV3jpwCjBWFRMDCUeSuc17MufhDd3
OpMCCvQlU+ipz/rTMVlKOy/wj9JIrsCCQoWj/yiTZCEOwGj/QxtvXROp9txOT+/c
lKI9uY+AH9x/vg/iPzhLUjIWoscqRs6kDj2vW786zyHpPdI4L6IFXs1w/ShT86vc
J5jwkaOKpDFw40E3ZJHWMKzGFnCmyPikg44xRrAT7DfmkVaURfju3IG7UJAyWv+i
/ADcP3nWMppLUy0DBG1/wfzKiMbHfTS92tfvRMjnJzK5dsvVqxuE5acTT7Tcu22z
EhYEj0tpexqe7hbf55pJjt7bJsoZxO0HEXS4U5jP+E9l6OWQl8rryIjeerv4upW0
C27HvtMumYcRIaZQgd3ebNTEs+eZhESSbAdTRv6YZU/66Mhx8G1L93gjLbUKVPN1
jE3l4m1Ad6feJzeAoXlqerSUWPJ3yqiYe4lbVXoZp0xxTezBME/5KdzyoB+3XvJm
iQtm8WhLTGLMxl1VhnVzY1kX50cCdzs/2XYWkvX541G0AJtatu2HABQkjCTNaeA5
XFeMwp6iBtPHC2S2TnvTc2+vMgEVURyoikWYkEZ74X5ofowmLj9gCt9alDyYjVFI
M8+j95A0FxIwIlQewEnvnUIj/n5algBVaWCewsgUMrTPoDK0UDuOFf34Wr/XuyaE
UHn8dUIocH5g6FvIjWm2FjsD3JTjTzgxSASY5FvW0B1ATeXDoEnZ+4Ph4t3v7RqW
JEnNctrgqY5/PfmA3530CQqMffjpjYXOv0ss2z3jQjKamHnqG3/CK4ViNvOQ8DeM
QZNjtuHVCiGQGoQssw7yphFLpVwIFf46A5D5ZlVaX7/bkM0dtYtujyTaDkleDIYb
461TQPFbgB9MlrNhnTbOAAdRXxjl9iDnTK2pWePVShmdu2HOYNRHwADD1EmeNCBj
A2K3mhn2Hj5aQBZrLs1G7K6Sml61alg50PzN8RR1b35kc5x27xTjKX1d8E6vYk3O
YV1UqHLTdDmEhH7XYEcxpkDVjPzhaDT/hTW7C26oNkQUsUYuy58NJo8GvVBl9UqV
54A5JdMH3VorNHOjMI/YqnT4hh7iMacVpMXMqpu7qPbkHPTGwzweKS3DP9Lw1BOL
7lww8JtqKZM3ZHgJDCE2JeHEfqQ+02WYAZdPSst/Xm3hpSrHHV06/+FbsKr+5GoY
U2MdVi9MPj4VaLQH0fJ2m4cjrfEd6BuzHsOEA/kx5ym0LwTH5XrkjkEv1QPMCrfV
FzVJV5oii7D8LWbiPVFHWMze3zWOQ/wEUghricykq5RAlgvUXwojktSLOAYGmzW3
yMuFZOQw7toditdI2D6vgUWjQLWNCI8g77xmjpCOtL2SCAQfWp/I59FP/llnGRfd
msVI2ftPFiCkUEiDTWVoS7mxf3CnJe3hCjJ8gS9phQlLUuM3+TZegCJXYQ44bUEX
crnyiqgJofdHm0E+m97LfIMQ+WiL1GlyBrk7lUIFi3LXZd3lpceMTztsvTl5ZPgH
DhoJcc+faWGWbRJ31h+YlaCfJN4JOWetqBpW4t0pfIUNjwsaZ6SoWcx+zId4cmfm
3XhPvKiwL4GpU9iyUj5H8dNPhqOM7iPeMs+cxPic6QqZM/rrVSOAWN4lfgh2QNWA
WktanL6A+6Nz3c50zVQEW/AmgQJVE87QqNs9mtynGJNCLBZafYD1DEGQu2uLcMWM
nC3WQ2ODrgj7mpD5NwtreH7V538ICu7ta65o+l32v4g8nneO4fEvlvxIswfo+AA1
KRkw5INQOeQDWD2on0r5AUh447sgDAoNjeuLCz4s8nRv6CeJRmWlqStUaG9t3RMP
wuvGNwuTwXIF9oUG0n1ZR4UkOkzxphtI6Be58jzjZq/qGUZw5j8mMMLi7OEyK5ao
Fw20vBb9BO1itTVOt2eLpvVBblKI+4OX+pQgJboxENdL3lx+wo7brx0GBhgCVLwq
7X5DQIq5a67TRuQK4KRIjw==
`protect END_PROTECTED
