`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUqAfJi8XLqKAPmUVd4Rwm6A3eybVuHLzie/BZJW5Im//QzYh+N5X68Zf+SNQWnQ
VztaLCYYD146OdX8iGqM1/9PzOaALSTmtEnU68T0Spp6XwtFY5r0lLX+hQhjPBRL
MEyAQdcM3UoRqEIHG2e+Bb5TV6CR57qoLe/rAjvJ7UbnvsyXYOyULjjcHRKFIL3E
iEm7rUF/ieMRx905IHQoQZOyVgyHQoyun7g1OqsuoV9mIYEbtk2edQ2OcnvMzv5e
xeKKdCaF3AUJr/jv4wRVaK2GJ6hGYx/Zr4gNrz5XEZZyp7tSQ1xV0y6n3gKB7OJM
cQQmetFQrl8fvJ2Lfzr+YirNavj7R8nYRQG3lyDmSffcbeBpZJT1XLAjPV/saJjs
ZHqxiTIEWOunUd5DXSyjGd4qOEUjzy5M6bu+RN5vrSX0gUa03QCvuTpwSd5joAEg
Ejz5zhBvFRG2JwDVRmIXYqMu380uH930YU0Fu2O1UB2PJSaH2DJrDLnSTY1Cx8ca
ZRFSkgrqdTj8qqZEUhjaq4Du9k0B1YIc+gj31sQvX42mVCJl0c9RdbBrletFH8GF
wc1xHUEDoSXuUfkUjs/LjTnQif1t0Z9NIAglZbX9NlfHmJfrcJoAOTpeOKAVI2bS
OJFEr+53PKANCKaFjsGvlD2otjyeBaPGq1v6EgiH0nCsaKNEgyRym3eV5fAOeYBw
UCw3CHCgH8vt27lxm8VfdjU0P2pmUm0afMaBzOciH5ZvYGUmm6fEIC1E53nxbV1d
VGuWWWBMg94NHBTz9U/XukWOiruf+V2d408OZQvEa/v6ma+NDqLT24rik8bW/f7B
ApuaNv+X9NyXyheznLY+mNxxHBjvpjVqsBn4fHjPpwFSAJcs8PK/v5dQ2ApqDXS3
6G8620sLJcRngMnsfDZ1ywcOunAowGkH2laIUM8KQxPtr7TkGZgpY5ivOG+a+oia
rcNr0bIu/LpqtyrojapwB+9Vkiau1jN7NnnfI9Kw/PE7Q3FkyhtTj3sED8sM4GpU
f4C1Le1dEArl0jOd/n2mkEiFw/pDbUjelSPMq4fgXIRMVpczv1Nwv2j0OJyM5Q3l
qO/98jePtb/aw08Xviyu8HkW8JifvGOcJyg1ru39R8siyh2/bdNpWd6TgIQP8peR
Qguc3OPuPh0b0VQo3krUU2kbYix6tezC95HPy3Q9oNL+qTqobzUNLd9JHlHb2w+6
75PMdu/F06uC7RJV8X77Ugj43y+Teauac/Xr2Cs0+7y6FkZC54NJ9mSmafSvx4lE
noM5cAdPH1LUopQ5HsLwYmBiT4zVXCE0cCz8dHkaEx/jf+jv74zuDY1tqAcPl5cE
2t1lFTDo6HpSC4yVulYRQyQfQjP7Tw21k/Woh86lyKtEgWGdS+wmJzDNzwNdv58o
grCb050V+/pkYdYpVhuHaiOZLE9Mdh8vWd6FLw0shhnguPw8fdYRuLnmTcFlSahO
e/oZruvyBglFEWdYsDgJ2VIIRh51Lx3F8xg/uufLtJ3XT+o7pAz7TZJd6ZVxAl2O
KCs7tMzFufcIcxhn4FgxgTDGGC6GtwkOAetazz1s0e3QUrW29nTcv76X+dQefcti
QifpnHRFmSUcS4XcKLKzz/7wyUjXbYyh73XcFrCYobJBtXbUhCdhzrf74qnjaWLu
o6jSuTGGo+RSNCBtGtiTQY2oOpXyoFK6qL1rz62ulz0=
`protect END_PROTECTED
