`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sa6kJORMSbdcvo8X0RBO1vm0Y+h6p0PRsM1eJ4O+GcmAsRDgHgqcw980qcCrT5QX
62QvAxmgdE3sR6pluCCLVhuTTM+yau+0vCREDstv3SOUCH07q+BPwYL+9kdOrxdZ
Y4Rqt2Erd39nTDmEbeMNlVQpXyffr+Uihb/HpuuZ7KU=
`protect END_PROTECTED
