`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRx96aAiGSgSrFW7/DskCvyCIzpXXNJux9YDa5K6vCI6BW3lSkMzaO6ptCtSqImR
0nqC9ZyLTDkULXfA7FXDH5bkUOmE6QAKXngWyY6RUwwBrIj47WqpEC9xZst15t8b
SEjycCHRlvabnFjvM+cduAg0oVphL300N/i4Jrr8RZNVT0U9zF5q/3HyRn5FZpgA
u7o/515XxI2sRtbv4l2mys8mJtXAQAZsPRMB6BenQAfNmFiA6cEI+kC254Su1eoO
vyO2Gfb9XFTEXYlED0trfSxDe5baGQJ4OppPIrKJN3uSiI3l7WzdEKr3ymjq3dsQ
zmENISpSWimTNCMJUj9CbXCGzN3hXsyNpkDLMHf0zH8k/zxr4ztkOvM+cXNBylKZ
t3yvRwSfddK1IfaA4YPgm+t0g6WnbIHXJcIlZhnFs0Ck8abrTLyd2yzEkvOQJmWC
Rlv2nAHTv/UYWHmszPt5BZPFr97C1HhIQjfA4YlZV5XxY7whZcycLhjJUBvYLnAA
+gqYZ640OI/ZsnLWI9yCFJdxUUkYlNasT+cDVj0snXJEWTaxigaMSyVUugyXuZYs
IMVdClm9MoNXoB1h2Zj5BOF6Gyy2RbHx+4XGzKWfmRn0iI/ZgFAKHsHcvvGCkOP+
Nd7FnjuNB+y6bTPDyJNr39QPtDXQ9E8+/Yks1nTfnKuAHEqy+WujJB4MiXs+i4CX
K+8l5P0Khp7iPY66pHlcVb64rCFc+fvshCTMuWRxsGJBrPMSOUwSVYIFPsgtE8OG
mx8pBSQszdKlpf534cS/WtRmEgHNquNHS6aaDMxmqzLZ+NejJvojPbhTsUppuuZR
JLVkXnNI341hNVrVy62AFRltWyIUhwNYcfFo3jS4vv0E8uqzgaOphVFgsoPIeAa6
lwJLOgOwHX7PUsoMYKLQl1Q9G/Ia+TpyVnSyJxK6iG5FInEGajwuRoXrH644Qgza
jxJucvj1FxdTQKHpFgDYhZjn39di68AmG5oCloA4itCw8VM5p1v+jURD7vx9q/Uc
D4lUAnSZLBFhnCLjYm7b2FWHt5z0AQKm/eNZIePy+Www0CBRTQgLBaJ8u8l0AgSu
FAvDuey7ct3VH8W0uf89LXao6W/yi1TbAfDpdDW6INtQ6L4f08MWgXawmar8FPA2
3c8+gE+JykMIYiTheIbZtuWZysfJboCPPev2YsuV35Rsa/nKu0Hu/YhbD987uavd
UWQOB/KA8lSE/sZASj7Sz9Njn8pAzBRvKFrcDVO+ZDbOcyMxK1WvpmTo6MLdRrj9
byQs5WlNl7yt9bLDomrnQK41wf3AD2vTFqPUaPR96AiITs16LBNhq+8E6dCYoAFj
ijHsyo5Iljk6JaJDSFf8WAf6R8yOlClQT6vHBTWxp6U4/z2/2oi/z5T0ZN2J74Zp
YzDnJU/OBMGvbBJouCu1/vNQE23ewnc0ojZC6XC6vJDtwoo52xIAG8zHqvXHwBuu
6bEib/UQnyqk/fvGi0iiC+iO4erMW1HXi/n83VRDO5CKc/3QnuB57ZESSqV6b34Q
6/JOmWtCaSGUt5Ua1nGR+InxpQsTJ9jajgbBBLmSXPmuq5Vae3Xqr7T842pEvZki
BuHaNf3lOQxuxb2Y6W4j1AffLNq0sfqzrndV6O2mz5pVl/8IQq6MM4ARH6tChxsd
w/+SwxPFtt1ZiDxmLY0rB8jXtlUWoUV62nEksK7AdYjyAPWFOqDfdLclUsjs34CD
rzaIo5G4cr4erwWSzDw8db01yhHU/23yjlLpE/DyXn9tLemu4ElVJqHfkbSbxiXS
fzHiTuX0oS3IFPVKnPeJxtAoc9pd+KQggSBOCKw943PmLe3Ct+RPB9r3tsbN5JMO
vAzAWqSx7yetdtVhTFA8FD7Hec/8D+g6JKGj/MkcKGZTUGqlGDbJ97JnGTfERomR
LYycD6aBpvSHuZsNXSSZUFJn4qNTTrh/0z+1pQa847mJ6bxkqA0yRhi3YHQPj0dj
eVokJzKNBU9T//sH2/jXpm5mjEVJGrMSHvO+aG6+reZHH0FRzscDSHwmH2/MutrK
lFGiU76ThqV8UIeqR/t6tgUsouNUCYdXQRsSDY4XifTWB06jvAo4IsEInJFgkdKQ
lk8JmKXIQC4VrYgkdW0Ypg6+cfw7AWFLfUvrnnKc19xxbGL1E/OYgnk38PM2xG+t
hbc29iLq6/84BUi132i5pO5/L1pKWJkAe5l3/CxrVYej9xdh4n0WqoadYNf6cK38
v5uKT+f8hhb2T6aKyUv4TR02IuN40kJK6PWJLLySZ1UnpCAT21kK/zCvzcFl/N/c
+tutSyHfjHScw5wxfgCb9TGjySiyWdMlcAf71mdKRcqqP3s3/Wl0ZJyH5MGOMm80
KbmRd/r+GLW0x2hsjZMAf++iJ6v57EPqc6WMSB9py+30ryfBtihPsoPKhOv3A7Q1
Lvsiff+QKm+1uV4VzixHKtyv662lH8HuV6gBZy+wvcZYTU38YwLXYIltpJlhuYFG
KlBOdtC9vChUoQRxpqglR5VjT5YUVw5tLeG0rqx336RE5iV0eeSs2uynek9723EH
MYgVsMNLKDjmURg4ywAUHUwB/IshQJDyw49YKXfmhOb0ds1F+hKuknjoLwGmOgsG
kpoE2+HxbqRaIl8KaiAdOM2XaF8W0V0iNNGzLFjWyyLdOdDd3rlVVtS6bmMRZdOr
C3CaeUAIVv77UwmVDSctjRWflsFOORoBN3mMFztI5CHjbnggomxKoTUlCmssNuGd
dnbhCb41/tQb+rtk4jQmhAbRcz5kIPgtundBjxhOfctrq+RmsnALDJqvkmMiNVR2
7SASGskPFVTJoVuVR7/Y8s5g2vHBZ1MDOxaGaVq0Lg3lXuhfxC0KE+lU7aIonrxw
1zI+fPk4K6iNLIX6P1Hmq6eRcv8dzTBnJOMCttohInAglguGUoDwSi8ZYywct7+j
qJ8yhOm4fEnWx7aNtTshqVIFc4dEtnRZ9AbhsEor9GTAZIsZsYnrEA5GPt/to1WD
pJamrq/FhZidM99qVWr0m6HINk1cxc9tdGuIK/z0t3Xt177vqHoftNZFrsLFZAsT
alUZOn9gOos0TQogDxAq9+6jt/3a+kai1niVs0GWwe53yYqekyPU/mYUtSD6Rr4L
dJ74tgurlkp4VKGrz8OxJBR33w9FMBpc4i7HuJoVFHAHFWiWURyIUYmg2Kz0pfxP
PnCC7HzFPkLNlAe08FaX2s/Q+54CFkXIEOf/G8H8JCcgp3fjiM33YRaEd1zmoun7
wBn9UhfMxOFOpeIO5s5YFP6x4gvTCnds+4rTrSQMuQjlKpojWxbyszPKUbcwgqRf
yGCnE2Jj4zJcJuUeDqaSP74n41tYbBis/+lG8ZzmluUgjsy4yTR6R1LkoiPXO6/1
ReEZwFrlqP5DhgdgeL0H+r9wmQFnwOx2gm/YsVoEHGTmL+s/M8cBPxJhVEzVc+Y0
s9VCYK359UQ+VjuG7NipwDhly6EnZauDeYOTSH8syGjVo2Bh7Jeso62Dba8VRJjV
DmwT2rp2HAWK0LLFeupsxzKXyaTTbd6iKGxYIPxOUFcs+fOukYceosEx57ddovwc
BuixQn+gtVsLOSEwf4A9QjoaV5h4HPaDQZeg4TSuMHgzTz7TIiKogZF3RFrh3hFk
F4gk8stV1zRy+3jbWgpfWBEXhEkQiFJFBtRC7llPhYWeZGv/WKfPnCxsDT5QJ2Q2
zwLcUatp9PD047rlNW2wqxL8Hb+1Dp6A2BZsGd8nq/Yb2fur3bOx2RX9qGV5jpfu
QV7yqJjHqhTiwA8ZELULmLSGM0kHLyjODNtPkP6HfSEaUibU7MotEmH8iyCjh1/Q
/iyMtqdAH8NT/Rw5MFrKXnjfp2EIA+61gIHmk1fC27C7tQbSZvDFmtrYeLRN6bZ7
rN8KfQ0o1/qSYmjXjL+byeOSfdrS1krAqhyEZyHb2S9QFKlTfmH8sGmbHQa+IYNz
9EkClWFW6YkBeT/pj3Otqr2ccgCePL29zC7ySeZQ8cG5oP/U8PCzdBIH9dAjqInb
wO2s5x0TPV3b+PtbkzbzwDH3I/H3QiZuvpzCpjkcjIRAcVpEDRPEdTHKXGL4uhUA
QZfcU1hurjvQl00ihufvcrdJ6CwL6NbtnIHBPiR3dFtQZdBgtWpk5zXebgbOLNXQ
odNY7/lE/KjxuOtRD1Wdad2wo+hWQqjEDtGQ79xJ5RrWkc6Nbq1USDAlgf5S3t1V
25ve51j/Yt3Mw82QjjO9PKOAl//upCoFb3iRvkwZZTNOfVwuOMPKWn23DQf/kFit
+MIuypehoFtblOlAfP9dr+35FfvDCDQbKncUDLsK5o1MwMs+xCPVmHIWyWXozndm
PVZPg9q8RMwueBa3mBr0URkzYVWXQKfXkQVSbulm6oM61hTweAM9bRkMktFR34ds
tcLKzizrgFLji/dyg/qWpY978+M2cJpmbxfhG41k2oquspPddExrNwjW24lv8IOZ
W5yPO+0K+znAAigw45zg1qWdNCQsA91dvbtDjxDELK+NYtqeaRhXOxKdEgO2a1u/
/AmHk6s4+F5oM9IMld+pgdv37mw0i4eRJT4nssaogMmWWfR1KPfXOlwvdy0V5VpE
JY8eKEHggzMmQpDG0TDavucrFl+zLEHFDNJEvm8mx+iOB729O7HDStlsnZmKxRET
N7exu9lQHsQdHk3ar+hs5xI5wiRlct8XYf3ffWjmYkEzPz+jdyIJ0nz4lVQwfoEo
SDJfLJQ2wryfsLG7pZVUMn9GAQCqEFY6C3hH1S+67ttXgPyQCF4WSmK8MGgic7FP
50P7aCBpXJmAIwbC9RJWJ7trFMBnEAWE5shrk414y1mNu2wm+64k8dt0d+E27eqJ
QaykqysybHz3Wbaqi56aw17bZ4j08ku4nqK/DUZREHP4vUgnjCW2Av47T2M4BVoB
SQgK1v2ZJSrbfpy6NqS5qicdGM/fSeIJmg+GZATiloY5ckaewDsuUlLMEUN64/SY
Z8w2vu7qzwjFNaRiuXvAbRyAi0gyKLytHea2R4Sgu10ipJa+PUb60oVXG35t7DYf
NLI4kQ9q6HlNZYN2G5A9v7Vg3c4NhSXrdOLhYkZ9hjvN3OgBqp7/v09r2usOsoDR
Iz9nq4TXBGGCsJuAKN0IP2LQoPZPK+xc/WHrL0z42KrJ/OIxuaN8uICJSgNT0ecr
oPkTV7P417VwOaE98a2U1Ru/Sf4r4laRXMuvEsmefDY4waGpaIft/uvx5mjPaHQA
PpDL+WyTQ3lNJAWh9qe+FhS+oA9Bv6HuO5I7Ht7mW97gg9MVi0Ie4xZMvaEDIEGj
MoO0MrksRd4SHleB/cdwacpMxUJ06804OMlv18+iPoF9OHIdq+8KLeK48ApMxU/A
DARVX8J8y+xRr5solhBeb9cbD5U6Lbaxfz+vtI2ht++toAGKg/3w8+dDuFN3x1ht
adB0/jYS8fFSu4pgcfks+ioP4Qb5Gr2CR/LwpR1OWlXHdfEPyEP3nshj1ALPFz4B
aYm13zq2Bx7q43w9ZyCb3Hr5CdssHnVaGEX4ytWcniKh33IRhXhklrJe+1bDKnEV
unwvhnNrSamXLuPj6sR1SWjRHBq/NtAXguLRgR7YI+658/4KFiZuYo/jePpEYnv+
de8As40BmEj8KgQUbCftid5vhUEqI0GFkuCwUGPU017VbJWk6b97IiykVGZW9BAx
V9mI7W+a2phzz5KNdiwD2PQGpDZFRGxxzZ47bozBz+x4XZ5Pbqc77LU0qUdtIhOQ
ajM9zi/Kb5LqS8WKoY5N2SB2l30VG0++HTThuqHCRUc1GpUWQDrkehczxo95SM7b
0hI3l87Auw66joSAiGDmC/PaaoBCYEcdqYAqCkwKSySqNvgzPUGWiYn27vlC9nqK
1lTGTvRftOoHlQVEmTL/AYIDLV1NQjRFbn1IBQ4sNHr9KGJk8m1OBuNN+aOzj+J9
BKYVaGqlOqguYVcfyiQCf6nidGL5m7xBLNrT9hwbB3ko//eejwAUMaYGV0C1EAiF
r3P4ZZbQmSnm1a2D4Z0ZjJB0A1zLsPXeDI3jCJR66Haj4TkVTCYCF81cmVhfAJ4U
URkiXJrhjTa40/Zhu2bD+9DbQlaeo3L3Iasbn8lHcr6Ng09HyACyWlfB6FYJ/Vye
CpvI0KGksjPxjsTVywfxxYbcnpSaSs8wp5CIgJKUdeW09exKmSRa9Xt9rOztzr9b
kYs/1viNiCDkQPRb5bMEm2mq839sUQwMkBn4DbJuajnSzI/d54syvYxIfP/dqZAG
gei6Cci919iSuOK6kZzxsAm+QsH8tiNBn3DCCajnSoegr0rLvE+32RWHMoXlfmK+
wj9Pmlo5RVJZCTGnls+P6iUNyXVrtDKbv+EADcrtGfW9n+wvaXVO4y6wQqXaXRup
jdXQBBN3KJErFTDeLUT6fW4ZuVRmcmpYYHoCyD9Hf770XHY2Ix55RQOXLJd2FAIl
9Puz2nfkbqVInhGAByhD6JYRo435rV+nzQvFkvP7vKUt6jwxkOxMEMnWdREfMqUZ
EPsdY0nToJlNtl3PtA+1SghQXu21XVSIgKm5YUj/lepz8zRTayaFFfzSDYLvlyfT
/CerMAHaBMMgeSP6QQ7nU8h/y1lX2yfmfObaGBFhMiGlx4tTXuYk0pz6LRWwRjrv
jczaM4Mnm42qnO1SmSnIARMEbBVZwsDLOw0j+wRVSjys9ORbG7zuI/j/ZWdKp8Ls
f15msNdmFV3CMlXLZJX0ReTnsE7zdrxzvVmGSzSs1LIdUUCgIQfbcYkm/sClZeWU
v0/GrTnuvRhumPWsDcpAOS9CGj3w8+CPhha4a+jqRUKaRSLRJV0xEanQdA3qFyhf
cfhHaOPjN+WZ5sNd0M2r9fTcd+yu2N84+bbbFvK9A/lCsiROge0xy7OAjmfK4U/E
HBvHHXywduuNqksTOHF9hfPegI4r7/cKt6faeeEvRBud4UOl/RAgagmXWbn4hSog
uMYW0bRygqkKvLrwveEDrcTIrjtWefEvBORkQL8vbX49sOzQVxPp7EL7C0zEP1/w
UaKFQyxNxnH390tJFps8l/vvEm3HxPdDFGhSj/G0JYITBhXzT31pJd9Zdpj60FkM
weU7cbrunNArji4YSYVZPYBE09xdMnYrd/caZgrT7hetQhE3ye7uPDh2KxBiDwXI
4LdwfekE0ZxmCWzGWA+ltoda0Nvzg4p8mB+rETQf7DWqSXtchZS0wrSTXhJQz/Iw
u438ecDAoZjyRnkhyBHJkInXq2PUxTKRo2Fm7/lTTqVzosvVzdWCtXce/mS5xUaA
yib9/djjs89qBvJM+KFifHXSLeEnp4QSLnNLblqc3793wVdAwonJue8JvBcA7f7Q
+xx0tR/wJTy+HAA6Aog1hsAZPiA9oc4CkZw3vd5E2/aqJoCfOkT+ggj83K1vCij5
/9EzZQIDLHSfH4BDM/3ZowUeoaX0rY0RkGvDDz/gv4lSxgCLkG76TrvQCeEazvd7
P1Ov3pyx0qWPQw6JHXMjZRlg4XAsD4JZFjNr0ksxIE9uRCl8Td5arOEXD0dQSXeU
JTlkIlBdEaFUzLIua60PBOtihZiqH+GPcqzclv+U3+DwGUkpePHPdDeVmZr6dYcH
NBw0r+MWfYkHDmfjpksmO4cZI8eKoR2jks/BJk0uLDQMjajFwRKDY6ujnSF89P/f
CLaD2sTzkQbkb0N4VFvTeoaQgRnsg2GqXjN5u2rLIyy1zF4jjFFcRK5aVVOcnu8H
trghs4lhnULea/D353mPZKNbFfty3FC7pGA6KGOzBhCxg/PakF3+fw4xR7WICj1B
mxRRHHuj6vFYcrJh+92tmkCV5n/PiqmN1E4LGdID1bLa3mhZihVf0wE6Xdjnfts4
KWknqU+m6LFjRPrPmOpcHh9nXcOurszOnskhTEdZdh0LzTkuC2phxFzH/2QLs9RL
4yymovoYaJjblt3eBsNXv1A8mMvobSq7U6UBSeW1U5yh2QjqZSA9ZpPUEuX817C4
o7oDs58P4XcbKyngdC7frxw4lDkmFuCHA3r77JvUea5ebDLpf8EebUqIIjV3L+HI
z1rSRaJ5rt2Wvsa+0MCTvaVEi3ZFtMpT/gaRe0DzqqC6J+ZVgzfmOT1wHXEU6KzU
grNf+wzw83wmwp4rX1yt0aMN4LC1SShHsFHcA6hlQTwmK+0t0TxpFSRWHi7iC7QT
NwD4MpqveSQ00WNB0yygaVJTm86fK9Ft6hva4MCkYktrev2uxce5mewWlF/hE8UG
uxsHmR1WfnUmG+G2Jh7QdK0PPCL7/bBpDUxulD0c+p5wPFHNzoaADKGF2vPHyELH
iNbja+QyrHZAqa/BZYKlcPUMYCoETi1+ecL23ZjKN9baxEVbTH+LV1J1CMblGHKD
lcGaB+ic5jrcaz19Tb5MdVE53dRD2cNA7jlJpngB5IUEkq60GF27b590046+znBq
UmOZa0MEqgNb0srfV8Xrr1gbD0IMcSKM/vK+pBUxU3avbUFo8uhd2zObxljvmBDN
kYzGz59mKES7Q8l8IjaxZzlDixZ4w5g7LOh2c1XU4OHG9Z2YIC08HFRqqPPAxdUn
8tSj0RqFMg71Qz+J+8vEH6eVzKXSNDWkfOGpK7idbP84Lw7x+Rz0dAdLx6LGBLOY
ZAfWNWT3tk89ioNIugtM7GzX65kmLzGBq/T7tgZHcSA+ynTXRdzmhhd0MSRBV7kX
g9j/EjPlh54h9h/EKUQQRXyNJnRrNtLStQgwToYm724GGVYzQkonLpmM73as2jB+
nGYScUXJP7yC7TCOlPfxm0Y6RlUt3Y0D+7Px/bGSp44vb1C7rwgt2kdKOdVsN03Y
RYdgjysvBD3A8ej1zJs9aqo6CQ+TsL0WiLs4j9lweVziPzL18/LZi7LXf7+sO/er
ktk7jo8OPKMtV/IYCm+I5aHlwjGSfAhsDgyx45LB6bh6pAZW40fWkoCrjd3tZsvx
26W458EhY3NphJJwyjR2OMIX2svCBaxnNjjK0CDOnDxlBNIfSrSpnihNIBM9e80/
2Xcey62P9rgUGO+p5JLTiBusz6csZpuLTpeoxmRrGVuglazRm0GsvmiuGUxjs1J0
56exzHQbv8H+GRJgeEaPlw/ngz0Vp+fzl0Wf+gyEaRe/XUFfl8kNqSSrIu+JCdOf
pqZEa1m5KwtiKDqxwS2YiyFk4TaOIYPCQc441JCzvXp6Z+QI8iGEMyGjByvg4387
priwcIJvJbqyOhD6QOoGHp4e3gC9BbLduzZBtxx3bk0iXM0LNMMmq1fmViLLvcgz
zv9ffseRiynqWZbPI9LxojarpbSZZ/BXUczDk3+aSNb1GJnji5I2Q+U//yB6RCFi
xNuI3nPorBuYxSoa4DV7QM0HdubenW3vxfUj928kqoddQDX9aiiw5ez/u3g0o00C
DZkF0Yh+1VqIM0xSf28hNf9j/I4pqhwUmB1cuiN5jpdb0eAyMPQumdvC/n6iN+D8
Zy5vVAZfgrbFLC5KMBLionH6Ev/Xc8DsZJm8L8Lb/3u7fGpbYQZ09zW/j6UzLDXr
sa+OgHGps4s/+oSyCk4R149JCWhkSwBR05rYr3I8+vYidKqIFhb6bmdLeXrQYIKq
u4oDzxWCQ6SQIzqJAdScrfLR54Ef2Vlb+bXleaMmC/tgsZGB8sG2qTSCFFY2nx++
jR21jIIk5jSLKIwLknbtZHYT4zKNOpqhee5Er/hxfQOlhYksDJSrN9nbfLKh5yCA
Kq14rDJ3BVS5GD0x5qPPvsV+DlFJsIZdp6fkoRtreeUFEXRhG9KefULbTEhjWDmY
FmO8T+YU+L7hxnREarztVWwC0ykIq3b11h/D3LHBbAg7gWnYUvpcxT+Nz5JhJ37O
yudtOMKMWen5WxDPD9JHRhsalxytNqZsz3y4eH4JZzo3PMpgNqwatlZZXPk0XAto
7nPYi5O7ggUy+8qPtM8ACIQxgrpFt9LO6ivUzUT2vVnx9CgVu37eo8gf+51G3BHS
4j12+ra8mGBVbjl/Lf0KeOm7jlacpj2pRSQ6H3Y251ZXw+/UPoHMr+Efu9Q4T/zH
QILQSW0YYjUt7gr5+L4Av25lELiSL9cy0alVavNqQhZJkLi+1KBPhTY715DfTOe9
YF8I6fGDzhthiNjp10NiAVtjwbiSwObyn17WVjO3iD/uzCze9eaIAZ4wL5/CXSRc
JteMJ20u2yHJPrDwtvdFFtcPHzKDTWPoZSLdppS84PHYg5Wd9BzMMTBnYK7Q3CV/
XzvQiEmkmRPXjZ4OAoyJgfbB2ZgJmypgJyeD9CApk6N7Z4Agg4JW4FVQdMro5emQ
0NF3OKCd0rDWioGFiQcmxVVkspYhj8LUgbqjrL5DZlN0hKBX/zrx7Fq7lMiO1ODt
CbWjtnmv1FxzSPEdHsanQc8Rzstk4cHGWdsHTKl5SuG0RX8QWMkOKd3eGGSqX6XB
IAZHgw4rTMvDHmHE4Y1YfIZFPUCz6izPTCKppRaAwmE/+YGbkXd5aA8A0GZ7IKBD
w+BZ6BWlnAvU7bSvVA0vVqb/ZfvtCJBJ/q1Qwj/BPASi0qqb7wEwe0/X7FKRDg53
ybcX49tnDII5wsg1kFia5Ibsxp9aw/uKkLLGb7+dqMLB0llJKGsmc00qSKdsW6bF
y0lhFZ5ttRSyNIBIVU7wX35tXvtaQTPe4jqeeDxGUyefJwITKs8P5WjV+qR3re8B
hEA/yLmHFoLXhAHKNgQ2t6uBJPHuPUaoOxccvkk4NWKK4NiIgx+/x46MnYPPNoua
S9bYpj4GvaZLplT/UCjaWAOV90VyWk1sC8pwAShXa83xxRVd7W1QF9q28ZqQJB2F
JWeSlezmZnsnMxrTy6vSIiqeDwJ30ZPmz0HT3/mzWpDuTbPzw5MmA+HMWmfrhzJI
8nqUN4o44p4SBoHKcEMo8G5fIQuNgdZX1P7xqi/fW9nmI12OjGrWMFUmEPalQBfE
7QHhhwPFlA9hzzXKKUQWzPL767d/u/U5e0TVb7FRy0VxFZozch9c86D0mb8HKlol
hqfNbzZghl+0ezwu3mRjCVSRn1vQeLaq5bOU9f7+wn4oxfUVn80jdt1rLLYcATyd
p92jFCnpQ1SLaHjxacTKlAoYmrVKXYB0h9SXGliNRWXSOUiKz4lU1osTLl1mCFC9
OCdcQI+yLf6BGvWyzLVgSyV0vdG55QV+F0zzd0pY3sbvsuM5LRSWdqatfMRgIGtB
+sKm5WlnWYhNRc+2FHlD1YAGmwp+E42o8C1iIOuotz1hGg6i5IkA/ipTGLExs1NX
aHjHhWBRD8o2RCqqS7tcxfVi6TwLuADbPllaOiqZbMehKJi2fw3lW6ug09cwyv4D
jZKZEWm4tpDLgrz31a2toymH8W7qv9zS34pwlIPlT5+yM2Q3sBStHJMp2Dg7OFNf
fRI2CoAPmg4scEo+LoHlALjprLXRFZ0il3sXJXvGei36vRH2HDiOQ8YCmlfcHMJT
wPpF95mcN0u8qbugSIUalDuRFXdcBNB4l0cUmfj8SBTSlOgHxZHagdEs36fVgOFj
iHimVe54J9rLj5jhSYEvI4E5fvMg7Bdw13AamF/btGPgVrtZbEmudS92sDDxadb1
YpO1XFkeDXhtCApu0Rmg9tgQubMfwCVeCtjb2gpTpRAaDt2hrLMBNxA7Tfdod3Et
G7NbIbOGIogy9uuoy4fgbHh4VO2avljFmrnZYPVQJjjKdvcb2ZWYawKIQo3FQsru
TlO5kHaC3YxR8f06evPGh3eAdCh0SwCvhz2Hfk+ZjtR5aMj+U7db/W82S4OIOUtX
iLRzB+BMUFVnyTPfwWkzuNK3lNtAiUHUVflAT5dg8oT6EoG4hhzsiy/7U3OIwphq
WzK+l+qQHPAuAmUvHJZkp0SsfMf1U2o1zYkgBbzXHOnQo1ixjJfzsH4oFrUKIA87
TQAliq2MzY4KrfvPyaGBQopkPBpIAnrBqDZi24zO8R1jiQ5+mR/DHlQgp5Z28RWI
QJGmWu5C8NZnmoKtxj9lXrNjkRQlLrcjJEhSaHtwmiDIjTPyaxDBC3NDDeNWs07/
q4P0R3izmr+6bM7moocS7U2s9o9cnqh8pg1NPseGpLBNRmlkXEk+/ZSlJUTeDRai
PTVPAQ0sPTIlKa6H2l8G7e5cWoIs3+9MDarrX7/3OFgVVR79308V1lQrM8sMFx+G
7uBejcmq0YxbeW/kau7WHUx1k4DAOHke/e/UQjelQrHyZA9BfymORjNOLr7KMfc8
Vpk9lTKE1uFgOhsPRg/5vbfncjLbIQ7eNyPwlGVuslLviMwnPPzbUuKkh8wdTRPZ
mc/8YmmlCHL1ZDpPM6KPLEmaGmJN8uO9xPUlvCdbQErQ6b+ZPyHjdI3hB7OziqYr
iCDlfTxHr+hfgHp7V54hf+iWYYgtHmBkdupN6+E0sOOAGgtOrpKjC69ckn2xSbUf
ab8NSlJXB2JrOE4z2lqAOq+YbR+0b3yE4nkJrbp1D8xOIwTgJMRceHgaGqr1v6zx
ulqk9hjKEP2XRn6T58VIYGFCBHKG2QHV40PKFUz43EjIVY51blxqzy5FuOjXIU1P
bwoTHrPyhzz9Jtbvodwgpd1Z3paWl8SUaqZO+1TqE37OApE+Kw87U/O9YApvRr8J
LKSD1GoAr7KdZkvxkwuoaq2p5lT3WEXt85ZemkagKCwT84HtCPmf4tyKjeA9MUUE
lgGf1dR8ScRdGepFOBsK/IF3RynHjKf78iPG2Ra7XifC60VRRpxr02V/cWjCjRxL
l+3aaXbssUhMRP0GmPEHkov3ck2sevb3ZxwqAwzB0SKTTnJQ2Uzs4t21G5VVXphc
0KjDfyiebgEAg2qhJnrsIxXOkI6hq85rczmG0lJedSx0BUldkRHEcF8uvBe1wCCQ
vf1K/Qmfgc1XSG923YGSB8/23dAOx20tkAhmSK3gn3xYAsr8e5z39RkBcPat4xiH
OyFfvgQUV6mxtalhmDR9d0JCZgPWeRpM2w3KbH73vfUsdNaWzCOayc4yujU7botL
S2AM6hU2F4ozhXw1rdsxAonC70PQhJGmAlLYKIjG8MeXFEELVDFrsKWC3p4WfJ6m
6Ca7E+1M+cM6EA1THEpipbfaWhOXHjg9Yvod2iN39cOybDz/fKyGfBy+2RmelLXL
1DCMUXA5qJDobCNegyIM980mGj1dtbtflq3ijSXU1lvrNtOA9l1vKfqZEddM8waP
Rn98T349DoC4GfXTe8wyyvqRRTNULVHuxR6wIoI+Q5XC+mxF8D0kqjDLOQty4w5U
R9iHu9RzJQjY1Sp6yo9Q7MNdkHxWDU4Z/y016LP8mZJ1jMtSrMSEeuPB04VOLMzX
KG+VhGYVFriPa+K/mjjdqXTqbHp0StMB1JNoU8Ye0MYJdAFrS+KvKyQ70Wn6vfZP
BSFW/n9kMp/XVyJMsPfBk1edIn3+P8GYzEJfiwS8XYbiGVG2uEmnDeH/oeOBBjxe
RtkLrZ3eNr1MIFNZDlWSqnHJWkmyTJ2ml820IiDjlNWA0LaoL4v+9tKlA/0IGIF6
k2LsmaScXz/Ig8T0Uhx4T+/r3F7P0pjCWktvGcZrMlznzSGsY8uZ2qpGWZA55Obl
sfjcP+oYfFKozhc/M9IoCXNqnsHT959xCdJWupqVWUvMcH1AT3nqm1sDkVj0sq/3
YyBs9BqOq2zwCfgjmYADt5rDia24Iwb/DFxYewMdUlqCCESo58rG/gWDtUxuR76z
psIA+Wik0e+uMsjpXhb/aHkYRvtBJjtvTK18TALhaTzcrtaj7R2YJxrID38F0XDs
7gu6s/bB99bhmKpchsD20Z331v6FsNaOcBE9Jgz9oEbaFOYXOf9RZ803HmA0MnXe
NWMT9SpDKeh6PjBK7jevnl1AU7zcxWB7zGGGNjIY85vrO9bpmTcj4mYpVxE6egAK
fBvyDsxwBmV2mQ0nyt5S7Wjiam3vGaGYCvTqk1XbVZXiZ90jbC7sHjKAE0jxClXD
zWS8pNwLKJQ7g/AgcwSyo9B1/857gAxd3Dpl9axe5ag0miykBtPBT8biXCIxuvYg
IoJKEcYpVKukJkVUo1ypM1/dzF2q/0P982o5FXFDe4aP1imfNXVWi8SWxREmq2+E
lWzYG7z8vALwbINv2EYF3fvZ2XnI0Wr/f3x5SJKzMe6fc/nb6ALJrovbD0Wk+vHB
DAoScGMXMwjs74JD6vUBU9icmP6Z6PCmuLaCC0fexwcBTydCCHjJqHdnGWVC0cRr
ai+ZhBJ8l/+YFlzuH2KPCapDzsz78UfSgftGBOyGwg/rm4bJ3RBrS7GTmOBU62W7
GQb+Njl0mVL9jEefgkR9JLVrqmnA2knCb9AagmtaFnEFGc1HlYkpqkO5BoBPTexR
zG4et/E/usDRocGIvDJSMIPuzVItKU3lea9drQFPKxrpPI1iQX+5aRFy8/s+UBly
Y8m38QltQsTWqsuxqA6cYMEQEcqtGJdKrnf7yYLXqmnhpGcWyd1T40A8Uhc5y3hl
wK6CSumR65okJmM6GElRtunG8OHZEoy2Hn3Iy3E9idUPfkht1sw9TknDK9oXcOrv
6HI1KDJz5euuV+lK1ymvxp22lyWQKNTOAwn7nLWQeII9TxozlZB/Het5ahwcnKga
ZSA+J/XpAxLUm42p3eMZh7U46iUuqMKIJAwfjcnO9La1dbsZVtqqRayYYe/1LQEx
DgFwzPq2c4Cu6GYfuWE821fGMoo+b+t6DlLYQQ/opMgGl6tvUFkT9t6w6cUzQubb
4yGYRBvl7cDFWZM71KEi4NUhVHFQbohym8ozTGYezoTvF8tEDoBWO6sooYxCiyVv
jy4y5BbhnSgIhFqfhPc/fjYDKNtQ81qUHSch33zAcytNEgnh5318yqARybRvo4W7
nUJ/VXe4CgHWkk0x0nXDSmmRSOy8ZLlJFvMhiX2iz920UCXqkwuXa3Rg2+2T/3g5
LLwJZc/3tXlnbvfEucsgmv87aFKtgK8G1fTgctJy8awYjfKEb2LAnc/IWhJ2CTBu
++epZL2Plipmzxc35/hlC1KhP/eoHSz+2CtoQRgoLphWHZMxaxzvcor0t6jrRdzt
j6GHY6+kKtBP3he/NN/tLmCV2Cd8QlV814eQON6RoVfeCqADz8dMeuWM8TcvyZKd
XRYXR8FL+BUuWEKQnLkj9TW/bjP83FLZo5Tqf4y0cG3N3KhUh0Z4CDGeocwg8QH2
KCA709Gabemzneqi/i02MXhTmbgQ4juNRJ7TYfS1wMn5iYfO4yufc8wETRVirFm1
fiINyqaYjMAxahD9BpQlHAfhAlpIybHO60tpwAzZCSe0UwEhH8oaj68ZBRyN8Hyt
zekrC/eohAKz3BK6FA8kXn9Dq5fNdakQkS1on8T5EUokBfADOrKbZjUzdksgGON2
PmlsrjjAnoJvcoCplsyjVNSj7JhF5JfTaz/L1sNOSQI1KPNpfLJHEQYMgmetxxca
yxDhzAypVfuktCzG2jlPJl3Ks4YxLpjFi1XaCc2JEQK8AQNiAgYdRmg85i8cVCGB
sd9r/SSJ9j8q4oldJloVnp3HypykoY6rhHSAXmj+uNrUMBbdiVk7QBxhPCntXHTz
vkqhxn1Taa1XmE4hgW6GFNORl2gz60cKIZrArPOc/uk9UcIYV0DlQkgBcW06Gb9R
RITw6Q4sXiCSeJ2g6S06cINJUAverDLhffewpfHXdcDDqBtu6DAgR4b5FrGycD4d
dQ6tKa7U1lfi7Hvreow/swoXoeli/S93JAieeSvx0FYqIYEVnxX9/mgHvbbrHnm6
fr7mYwz0RsEK1SmUxzj2q3I201EmS4N4G6QAiMj+f04peWikTicWS+LeZvZPR5Ls
V/HQr0ZyvhsqSJg/dE6LDxM985ult/S+oThcVUpA27W5uJH4ND04fAcdeLlxczj3
spKxm+w44pW701gO3e4TGqfp1aEfT6w/xMlnovNOTnDW0rdGWfnWveV2pRWMEN/d
bybwTap7AQbLxzs03tv2Klosl3nkqcV6khkFgsKvJ+h7c6ow/NFrvweez7taWz73
Qm9Xf5oEzowEG9gdzenAm1cUe/EfqqAHgXhZ4ZgD64WqAJvb8HLke2mfqBM4p2RM
FZ1j5zM3b3ADcuxkN5cfIStM5yC9U0ymd3iofezW91sIqB/28NY5y4tXQitL4QnD
yWEQlzey5PFL/d6Wd98AA5YQ+8aqSIVHOx179ujUZ13y7mOo/n713gHIF/6LAyQ6
BIgDeRgolWJxQKxK7WScDlvwkB/y8NmOeT8ozf9ssqLGMyIBeUtwHGLm8HNMFL5u
5sQr2EqJo743Q/xsDafG5NMmoYCYLCvaw17i4e9pYBh14kp+9aYcge4tBqVn66ru
8vZry6enTTQPRJxQB/YRywwlrdyfg2NexP2Y+ApPrB9wTswVgcObRmsL2vOvlcLc
9OE3YG8sq2BBB3RZwjC8TSZKIQOQINwcEaejtPvp820TCoR8993SEBwk4AFiW7fj
2/SgPleYDU4lkC9GolubnvC7nZ1wB9YzNZl1FoNrsw26DOWS3VqdoegRdBGnBScA
zZbhKpp/EVf2JEIhcbOtX484a0pJVImLEmYBnPZeS74nvZc8C7/wr+6B23t8Ne1S
3utVBUXNn+okKM856HnVKt0HjKpgoYosMPCv7jNNU2uM/E3xMIyEsF0/JzrJe0a1
/P/B76U2F6bfWRdsQ0F6LXzZZ2r2RPTs36Rs/RTvcDun6d13KEVlZW9vv6VSRI4u
KqLKHEWtUSbkRw+BRGqrUUPv21jC1arn3/CVbtIPTe+zs6ZYs6Te2ipdlKs+2pp0
eY97Q4gOVTbHGmBgVZi1EM5xSIBuNa7oibcHhSgr1l+glWqUrH2rML+Xen3dWMDf
DWPbW4Ntn03n01j41+i08GDcXKAy4CywoEJzSZP4PZ1RLLcHuNuo6zfcJQHTn0Wh
kdF/DT5MrhM5lDn1ke9jBZ8ACliO3jQ7QxBPqbIkNloZBtEgCI4pmtHdVflhpHKU
9BtDUKwmBOPnxz0xmTByaq4OvJR+vsqK1MClOl6g5z0P4CfDtuZWGgSlsnrCa3/t
VQg9SyfvUgJCegi6QPJAAax/n+Am5fMxgQ/bBrr4ZERfBO4EXiciPYd7yhb94jtL
lKWQl6SDIdcPU+d//MGfeXfAOyQ7qT95mNj3lfAhU9Gm2xyyU+ZOPCx2Q9bLg3lz
6soVkHmIZArmeuND+FhvOmxZXWhfQvD6UlKRZrLYB5CQ7TpWughC8ou/Jz140X3h
fp5p6PfD9jnuZ+wwWzsxhPDXeZaztAQJRiDAv8U48cVxI88kCkDGnmkqkNvclrdw
5AOTeZxa9zFsNfAJ7pzcK5oIOKsVbg1GOtrOZTqFGVRSKGmxx6GE/gwk0+Im39nM
dYgB2i+Nn+HPzg6tz3Zg63vBpSRxMpC4lPpmPPmZon8GCSFGZpqoRqijMrLzG+OF
zqB1RdB1EBiQORrduDM6J7BbUarvPFIVOgO9HlBdZumNN1w68ldftHfzrg1WlISv
64Bxkh91LtU12H27kQ3MghCwzdh14RqUs1cw1cslF4ipUnM9IUWykRWZkwFzMnDp
EXHPwgQlwCH6ZbOGXHaO2fV9rkR1Hb1oswUeTl9y2xO7d2lB87IwL1mgzUVH/R8w
5w5dY1xfn1gDDRxJyWiTpvb2D3h3ikMFOP+oLbCq6sWC9w/F9yDftfuD1r9+G4XE
2RVk0wOi5IF7rFORM9HDSVKhebkv5E1m6LosXBXiomNbU67y4wEsRUUJJsK6Bi2g
rhNjMhYpjOhcxsRKzDDYwy6LjTcS7qz5aMTIX3I/jM3YCdRgvXfQDTCpSz7tzclH
ztxwVixAeSa8ezSZUYEt1+neuRRgzS546A01Aq7y7LBcmuYVjkKAlOd4KHbhHdV9
9MMFLCqqicgn+fhO/7ZnS0RZlSqgvatUWL1OXWaOmdFnIpNcJvRUbSSPOT+hUxv/
xV75vhxOrpCwA2Nyh3sqbOk4GqoRJi/2MzV8NI3wzWQG/k/BuQmfADScnRewNwR3
HWREC744Zdoah3rJUxxvrExXebMJclU8VdtsuGmasJzFP+4fmVB/XAX/APEfRZnY
RRlawmgPthwkbdl1c4UTIn+XbmFbw//DfLVxlSqmVIf/DTLUUY07a0FSabeO/ub+
sBwQWwu/m0gfWyXfHYrx9WBX1CAuUuJNFdGAlW4j6FXCJGgy9o3MrJ6vkkA3cAQN
/2S3N54iEhEytsNzDCBAaw==
`protect END_PROTECTED
