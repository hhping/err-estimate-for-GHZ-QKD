`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dgXMsX4p7GSrsQCGOx0Zh1L8lF3Ngog6ZyKvNV2b9F5fjR3EBSWD1fllpXb8Y7Dh
8aS7TW8m+nlVOqPqNJa4XySd9Mp4IJvpCOS5IIXQCwVUCtzwu4WguZwOy9eTIM//
MRyx7QfYJfRCJr6isB5hUI+C0cKm+EdzUbHMHDVC3FNzVZJh/H2OVBveQNK5vcQu
HOqw6xqlDnfC8aNig2xWPD52J6DazU1PNhlYd/iO6k+lQxY2SbgFYRn5cb8Kj0Zn
xE/ZOzD1cjseIBcqL71uLpL4b59itrFBHMKgpwzwFpElViL7voVc0QksL58tcoJ7
upvaMzcZ740qz/Wm+J7vVkz2txla7xUy7YuIRL949urCQM4Cp3uhLK2R7t/5DnDP
5WAYO2CQVU+rPth+F++Q+LDb3C4Rt/McnlBJjxvpGodOuaAia0+CfdN8C6dOX23p
eDqjOddn5wroSRHGfRRPTqv8QF6M7q0QROjrCK8AZ6HjRkLcG3FFu0h2slVGion3
LhwmLYx1OgChlwUZqYXWNRLfKf9v4B0bGGhSaEdkG6y7p1PbXvxWtiy7qIcIiXHl
7wQuAaor08NjxGFFFZttmFL9vsXYnsfTKbP65/5hO8IPKlM6csxYgiTkEeKkZqlg
mogwS0ABTKbf9/ylj+lLkteVw/OC0ey7amL29yfn3pQtiGB+lxTJP77KohfA/cLB
DRMX7DwJIPGPxxqiyYMQJ2tSP0eL1ssjIifxQwkIj+2Cwmq8q9AleaBM9si5A6Xb
LK3i+8Pu1lbGjBTpydvscVUGXrgHAe1nzEiNGxH49CKSYsdvXhVgHz3g/dpkQS5a
CYW46J3rYBIdK0eiiG6ksFhRBI7BIfwy9njMwJq05nAj1i9ICYgjBmnAqC/D1HfO
BXypw+3cdDpbazn0T542lh5y/av18EyQ7dA5ryvSd/rKs3erVib9Y/aSMPsyMNmI
QdwKdWfRkvxjOkjqzh1stmY+TAQyMHUHG5kRDYLDUstVCXavx3Ag5XbBOY7+hewy
QXmJPpe7i+zKdXKgp2+flEam6FW3SRPCn2GH11b+64Y+Lg7wUJfI4ES1puYJ0Ma0
gMnqZGhUGNbea6SwdMvf35C4h5Z+yUUwlJgFcO7iZHRqG3r0nJ8ptIwIUQz1mK9U
U2GPT9kmGxH0PU/g4n/yyFLW/mRunU92768UNsJeTYqXbZeOYlOWkCKjPTkrYRc9
CdysDU/j+Zyv1ovQACNkkCACSm8pZvFwJOaZ0OheqRh/+F1x8NyMOy23NvT7J/sy
v1ec4GJ0ympIzFXcqgBm1nu72OazP2dc4+L38VAJbtqrSDxwSjkpYkjwV8Ww34Dl
5x9g0iLTNqm+71FuEcTocOfGQUXVyYcdIPcvSShHmB6XV/ZIshYxa2Hp7kX9Pq0o
whdfX1B7JTYNELwoM4IzBYKKYQtPaETJFUhdSJmpVpkKbZv5Po9INVWZGcpgQjLL
D0sU4GjyPcT7mt7FP8OJRa3seO/hsKEZNo63qz6ganznDHofFnpT70UToNFk4yGa
UilS2E352yvZUK3dMGxRgqFdu/rldIxkBNxFBRQV1D6Mpr2V2Rrtl+bw977Tu+L4
E03E/I6f7R3XUfaMiyBTtwHZiQrp7EY4yLY2EhjTyEmFP8UM/l802Ewee0Dt6+Lr
CubRsFaYvp3+B2f4rzknS9UKtUE3Dpk5x7e2MShV6x4ldTA6Sfr601UrJ0MteqZH
+fC5e8HaZ4AUY23S9xGo5H3ucdjHn4qUcxznj2MXFvqis6FwYdISPOSyRhZdpyGK
w2SMnsTRO4qnxqdStNF1L84ljGmjBej8xvFDYsT4NEDelqt+7kYsQvzxtCdbrztL
nJZ6ZNBtLmCMei0SAoXKroHXZVcjmhDMkZm/zMdhqJ3TlGbOQUxprH+EXMZX2IwS
MyY71UjU6c19DEUGgIx5QaAu2clpgbohBl9IOJRXN2UYBQdO5ltAm7AvsPu00ClN
zq5EW2LLCPc6saQANDBytHJGBtuA71hbXmd/H7gPCDkrCFQOu7HKv8QYE30wdnYA
vGzdUmduxo80aVFmAXUhQhzUYdynvKCHWcDJ5/isbDjnRIXwT0MWZTG5+H6IsgwF
ijfudLeDk2KnrbdfwvFIEN82xrre33SAiM4vmZn2vFczk/ja7ShqqOoUlW3RKj9B
gyqbwaQrTrZ2yjVyGGBqMAuBS1fV31GnBayJ0Tv7y5QReKksGAvlTzJOt+1yptvJ
6hUVtjTtuo/hmS4D/dqAhAYlHtX1mhRyEYst0QV+HNmAktCCnSMc6gJewQzsg44X
9dwz/V32ZliezxS4zJVcnBY4nx7gdUsCQR+zNHVsVB+pU0hGuaZWQ+4PbHq+qukG
d1LbYckBFO8vnkjpdawQzLAWmAZt3Ql0d8iv2MFsrJBJHlwgDm7iJMvX/QAhWd7t
9mZTaVYOkUOPNsputJlyCFNQ/6FE5UhdmciO/HyqQ7GiOBU8HtoNdFUUj81DO5CD
EvWGaNVazg5J0LZYk+nJB6TKK/MFBcRKLEZx9hL8TkQodgZ4SYGIVB4Afxz9NPZt
0Xj/Oblxs9EqrOm3n2LlAUbsS6//jz8wC6wWGuSnXo3vORJk4h7Za6Jgb8ff3mDZ
7kcY34rUv9juXm11by1Ha1P5CEFGA1uTQ1cuqo2NnIXVxj7f+UVnrOH7yKbLmrEb
5NRtc0vtzsOGwWxLEQcVXIp19mQr0yrZ1jgI5edMPBfVa6x0UbOU0Sci2NBBMerV
XTqSkdrVrCtXf4bSZ0nywEe5hIRoMucH6yc4BDuMhBUf9QnczCVi1oWzfA+jjseR
Ib6xSePyPZNToxdVQ6TNa8CPhr/34R/0GxPNkOYU5OSp6rBa+9o9XU1AVfrViCxQ
Wplw+dhavPZttS9oMhDwjqgcDaQ1REwrDp0enKZj0HKzbe9W57evRkVzWz5d/nrp
HO9Xi8ryFVSmQwkkpFcCES/DBwIZLr75axUwdQVwPJe5g4dLBE/Mmmy9ER4s5xnK
BPvr4irjcZ+zZdgvaGb52CpXNP1sLP13D60F9h5iV4p7UOFMjEkNrgQeRhEvNYeP
jCeuTJJ/gX0Z803rmgK6cJpPoTC6j6dZ82tjSD1QiaE4ov6aDz90M1lcLVaNtEkp
iRt3vg3Ld3sXlbfgaZbC4H+o74d0MCJRrGRQIdaXk0lRYTZFMLbEoAWqH55r8AyA
2h+eAXmjcdLMP6izfZ/ZCTvgwqlRSkTY+ukQ5pPnZR6N0QNH6bODC4tm63fyuqYk
2qVJGMIXXm5xsA9t7OOI6a9WCxs0rcHG89a8hcbeBd6F3aUKIfJ4JWV5Pcx6o4rW
uSNmf/ZFxP5BWyJPZdIeFbQagH7gKiydJ1xezXkzBiGu89v8qj6qhSMR+qbyUnI2
9TQIstWutsOd2HhIJHrW3stp57pfaJV8NjtqV7Z8ID/fiirO2T8h64I4kL6OXSxP
042apHNwSkXUL8xnThnXwEVqi6ZvoejR2m404YjCeqxVmoJuwrGL/H+vZjOwgw9y
w8rP6dvt3qTB5J+q487Njj2hkTqNPcdAvF0PloqrVstA+tiG7WfuWD9N3CH9Syfo
Rdve3RnUhIa76vpLBU4yG61xOv1bEOMTfovXasfypw8qJQLayb3CiAkwG/bxQTHV
xTSbj4MeaZNtTm90Yo8/x+jNeSA8afAphyPuQjZdNVWsgmXDLpY2OzHdpG2fJqXr
yoR8rPJMNwnYHRm+7UiqQS39e/JrHSO/ZqzUkP94cfAgTZgF5U1HHhtFjqQeGI5D
ilrutpIepJfMGKVR0peKwzQVDQUNyn3JPjIoJzZsJbu0yTw08IhmisJh+rBJRKxh
B8Wfqb/uRtJBNgAfqa7gkNgWrMlGCxKpmBICWR2eXL38RYpxQxg+6CxG4+334rOy
L10ZDSK9dQfHXxIv26iZmYpJZsAgaDcRr2jujI2jRspYS3Q9YndmnkNz96/YCbBV
E0HubhGAl1otPfBRjhcwYNnDeraOtS0As0UcsJACBAib2rfl00SZKL8xLiNlJEZo
zxM3GCg7dApHnnhY8bKqK/jv8TtVY6KkEl3yRQ9Ajm/GnH2bCC3aV8WRtVQFXCgx
dMCZM/OfqnvuQLTU7G+sgrvhxee7IVflI6nmv5KPa0d1IZRyQIXHhTKpgQAV4c3p
qKVwwPvpZF7ihqy+bpT1x0jnk8b1aQiOaKB79NQFikJ3DECRz+hJuqEgNBIInr34
mC7DRppXHV/nsWsM4ZmZny5GpmSD11hRr9XvBPYvcjb3rCtFX3G8YxqbazaL7jB5
lidWpiwsBSjinaahSLo17E82nJObq2KChWSt4YhFQ1FT7UoVRDuHtIilHy0dUr5u
ZnKSQgOjluY0XjGxYnf54DGIgsFIBTsMUtvQ8jLipFawjsPUorwnzwA3jERdSOyA
lM72oVbAGRdpr1+BQpHiojIO08UXCiqZjsrnuycrKkOhTM36g7PD9sVi60IaYi0a
RYMHgLzGDT65YrZy8fvnBPZus2Ww/B/olRXgfM723cAK4G3BFn0bamb6c3zbzvDv
GaaY3DKR1M2QVGkbpSdzJDJdPrZ/+/3XJ59q6h8pisp6SlriccWRDReQUuAY2KPr
JwRh5zo7+kORY29IAYOfeXAw3w5YaTK+oXAjLL7FroeOvD7Mdf9nlz0IA90OhwrR
dshWBrcanmYOgrGcDU4X4bzTfkEOLkJKdwZyfK5+oT5DKhlZjI1lInloDmDhIeWl
55RnrFYTNBC715tCeI3w3JJN3a375BvNwEWbhlly9xB15cWk6Fyb8PDFxF/mUU2u
wc7rtsNe6RTAxxJPh0eGhFMJehngiScWeEnEyRl8WGhA51ndg8JzGm7ps525BX86
igmKqYXmN3M4akOsgWXO0T3mz8MgHQtK4RAjAf/m8KsnlPPd6deaLNltatUo9rHN
XZPyGFVJ4f6/FjXvw2sPdTrqVKlifOBaeVfqUMM0RyLoF3nKUIfvlNrEjqPbO4QG
ENHnlhYgaziLr9yzf7c/6zfaw6tLp8dwTokGKrCzkL6XpeLXgzIqQj2clxGI/bZU
dWMhyqnwTMIwRKtkQfUJeTPwhTpuOEBQSxEbUb88HF5jokv++SRL7EprMr40j9Vr
G4nx7ZEwOKbwbRH8Fv47t1YSGfJ4dWPFZ+/SxXdGsuy0wgvCBHxXUAkcPuVnDMQo
ev5xHfmoBqgxFURmldfRxKc3Qn4MlfKcVFU9DFspembX8pLDgHsvDn1uZnY0Weec
VtB/FTe7F50ix67acfU7ud/NBBoSvZALvRMFtPPbTmtuSPFwXMVS3Bt1N4P/z9sg
Z5nCDFJkcDrSFGkEV2wmHn59t0LvPnaOJyKYI/+uQaliZt2l+qNvS5K/AMoBic5V
+vkQUQE2V8cK/l3AW85t1plCXyHfTiOGvCEKSCIpW3l3Fw6W3iQzy9kG+/hHF2uw
X8hKzKaM/BY2cefH0UagpJhWV9jatPQ94yce7pkuf+b9Gej3tIsyeB8axfWvaIn3
3oD9HrPgK72yIMFGAWpMRD/7XkgGIGTG9l/XtIiTFPKu8RdXoWfgWFAXjBovhTl3
U0On6gy5Zmmj7Z9VFEw+qWtf7KnPQ/EMfUPx0QA9KJ835FUQNNiYLUU4IzU8Xb+N
ewHzU66hAujKpZ9tqMkbs2J5cQTinV+FKAhkhPO+/iwCh4J51kw1RWicbSCDYrRz
nBGgALnwKVKMPjXdrgvGH8z168+WGJB+7dzXn8XzQgM7WKcDQn+nQoeaDuFy86NE
STnm365/vhuJWMIAsRRNhofLxmFrB+Nv+ibYn5+DUA5CO4wKzuwGNEybDXVKwq6H
tODi73exEXaMwMfHZtpQ628Md9rcDIW1uCmaHCm5QoC0Dn+GJehLiWSNjqDYpTvl
oMIAeHNLMfY8waRZdlQkm8bIbEpm0X8TiTte56EQdW41iXiC3jTH1s5BF+0D8ZaA
IuLt/Bx705KeHU7eKB5OYCuSWnp7u3o7PCRI+AhoFf/JBEl4ZncMXClnSD/p5q1H
PAqfk/np3Wdgxz2aDvSOlYwSBrgNfY9xubELqBTJ6Nt73aqMLp3YYqhcsYaV5sUl
ir7RVIzVxjmPl9kNYFYkDfE3bGODCEptUHAxSOM/ctvIy3zvYRrloJwjY8nhUkmM
vDaZW/C7+vO8CjG7z6Ey2k6j7mgpY3lLGH2zrUa606/dnfI3t4mGwjOFIYJq449l
STIGBBS7Hl1vAkXTr0HUZl59TV4tp0iaoYRBx7/p9o+kEUKUqsYW85QkY/8n5hDb
0xxMu0fj+TRVaMWGplVn47Lq3EtoKsYQfM8s8sT7AXLU2w+//RZaf54b1i4eO2CQ
OCRlDwSMF5JQpB9D3vTvMKmDws8D/7p/Tpv9/jX5fYobKoSJNeYjdB7JTIj71+5H
nVIO18FziiIVNAc/f1iovm5B19ecXl9/o1i2I4nwXdtQC4EnwluX+WWUECaVSfhq
y4VNTPtBFbpp7pl79NUMW/L7uESKsOOLrx6Zvipf5zD+bR/NDD2iLKVF94z3Ahvd
OmKWwCzCD7Fyw6o1iuy3+MWOCPfTRcn2PaYB87N8SB084ArwlFObgz0+2KhWLkeb
03HWkC8pnyGp7haK5n20uSL7+1KKWnWzRvX++WaGxbRsJX405gN3Yp5tolCg9vOK
3L/pVKMmYbp2zV+NJ9L7vJ25sx7yEJUepzzkVBYmecM6DQP+sDXePXwKEh8UYQVv
Q9jPVBnm83PHGa9QR+EdYbRN/mGyIZOEHGft7+In8oOM+p79EdoJ+vdv9lBAC4Rz
LcC81GX3FpvwhjQhbLF1gAet3Xk47HK45IzuthFVIRr84+vwO9dTYtoKnF3upPSe
ULsIRT18pvOZCZR1kVZbGRmxUya7J+8REeSm3LzIimBKGM4yCrnzr7R0KW/1n6xx
+bpU7umGV5B+24n651fLcOMTNQapeK6vzG17TCH4mk1slfiwmGoe+6gZNqULSS9k
8wE5uT4WK97LLkcrp/LMwgbJR5gQak3cmpI/Z079VocvGOrmpUG4+zQ2v41NhyaJ
aH3MK8Xqb1iWVu8y00KT4m+DmSW+XYtJgbR9b8N1IgTyEwUWDeu8kmH6CNTJ5GAu
P7yMuqyZD2wLmIsSSBNEjxpUZSJVQOJvXvLDMPtY1hzheCQ1+Kif8Kfiw0gBqkV/
6JKNI9o0GNGYlQ3gxXIxZO5eLZCUWaFK690QKTrXRnXETevl3DMnvajIC0ptX7sl
ZRmogePSzMft9akrkX+lRXNTXvUc5VtlTckSHSNXlmFmm6VB6o4UN4ptfbatIkvz
tI0TzkLNmExeVj2GBCaaqo52VzzeCRvlxx9NKtgYOuVYQYmA6/KrrA5XI5FlO0Cd
alaRZ6c2yvZgLOH4JYUOXLnl716atag4i8KVJuVMvaGjOmT/BXqpgEzcqgz0c0KK
Jf4mypObZQEF2oVe8ttmMZrw0F3N8Y6Z5a7sLGGqlI9QWlcLCP58pp0oo+6iWC+p
IzoHSkMdCIxT9ccU2f2w/g1qNMspQwZGDslK/+LqLQ7acBLVSs12Yx4QwV0BF0ZO
6PpbK4T/ymTYN23timUC//y0fOu/Kh3LI8ppnTg2ZI0Vw0ozJPM129Qq8OJW2dhI
fZagG4ZyOcIawRDqQ5v4DviWCcVvpfOodzEUdpgKdahKVE6xdnbB57GN0FHFihkm
ykOlESzsafrDWfKqnl2UA1hXAxkMrfp0JDkoIv9ElLOQYsQH8AJIov/zg/XptR9V
eqi07n5tkz+nNyI4EuSIul7NZnQ4/X4g2INqrXKsdD6PzPsENdpz4s1jxVtqnYHN
rtuRr4N4RM8IYdbMClrx+Udkj74SC7bPSUszc/+PSegLKLuSbDw1eh0pRWs8DWHU
z0cbXeV9cSix3O41l8IPHdZgUR2BMpA8U3rC2jVUhvk1ENUS81AAeZX1ENUJeESW
K3khdq/TABdXpO03cxj6GVZjLBduxj4KoGgOIst9tetfsWTQwUjQd7F1/8v+pAFW
kDlR/KZbT7b5OwKHME4Wb6dPqm4NB0Z7TAA1auA89lhTYSp56I5w64U/oseYWS7Z
Rhtz51VB1CWQIKODuz/d1YYvDmWxBhrZlLYMcU4YvArcKRm2m4ViSy7IMjYFplL/
WjE5v3go/hv06/7kYYa/Mj1LVaXAy77HXd/0tR4uWXer5crsQ0b5CD/YdJEnoz62
urShxj+lWc00hCRPDzOhQKyPxD2lDW8bYLch944woLcbZKaaT/5Pvp26z1m+Va/6
blMyjj8jYcAp9Jg90XgkqvQ2La4xY4VIYtWE5f50ZP9+X8keCgeSvDEKEOdb/9CG
PCgATsYrGjix7k+kQ63Zm5xE/C3rWiKs7/nOe2/dIg9YbzamGTkYgI4ml3c//dTK
aKOry0re1+0uH8Jb5VxExvyKC3WOTKeOVBN84+7BE4UzWd9ruHaP7tPN/yIxtbD5
LO345JeZUo8+i92YeW0e9QwbUaAEZu264Pr9SO2gWNItC3mLof3Z9UBpL9/2ghFp
0LufoaL8GfqF17kRPBo+4N3bNJqWnTjaIjWr5aEZMloONhfAuV5G2ekYzBHz/CUT
oPxP8QKCzbs1nppuxmHka2jvlsVG0QF3Do0XQNw7tNcpj3eKgUhGm2RC0wG4yJop
nQjsT/nW7J720LCOzoi232gvisYrHykh4L0iqLxZeJ3ONDSeEP19C+gdCYJcU40L
Y5ZrT4XpDAY73B1CQqgoDiBh4NKuQZxlMPKBWCU0FEe4b4cEpkM6Ah/MUlkPVtJT
QxCXPxuaFna8RE3wvn9mZBcomMMihRIGH90x0a2DQbxojl4jRNYYyCv3ehjSdLON
wOOpFSx9DLaTCmVp/miR7mkWC49AqeRGssvBZFYbPfYvtOmBnTUyapc0PGsTr88F
MBb64xdC7HDz8e6hf44Uf9BZIVUHC4Et7FCvKn9dife3h+Q5ZBBnA7OKklbkExNu
WaizqKTzK+z2ZfO9yr7klqLO60YxB9MQRUKo4tQYtMQKKgQS4KaLK+YKRr2NFJsi
t48fjZqlxIHOW9XwhlsDswtxVYsRaVrVwpXfT//TInPx8Pla1uOIuqFoq3tUokbX
jOMxIBDlmYWGGJhk0yPKY0iarTGwvNpCLiwmEIV0iCzFmoBVHRX1jsOI6no7SfbZ
KKWYE9tVpyyyvpZiAr0vYpY/GJdxRUIWMwLcJm4jzBqSx9+nLngXcQv+03liYNKI
Uqt7G9fIkscIrY+UZLTb/d3ESoHwmAkwmx6QcRWT6WK29RlT70NMJqhOOuEvASyS
gyTHT2ruYeq/34fpGbAWUoY3yhSUPU3nCFMgNonng1R94wCnxjb/opmhmh24csgL
hac7buFaVsWnhEtmLqKNImIIyXBQiWw3M/+JZWt+ENNtNloXXpY8mhp0nYBE7KfG
mUwpeoGb2SldarPqyxn6XbNZkyanArqhMXREY44z9GSfhz6cISza6z+0sxvCx+lC
vvhaC+Av55+h1za2jTiri9JkgQ3iubXitE4uhlkqGl1nnYbKhz6bwPHw1Y/0Y5kK
xtq1DEUbNFA0L0g2uL2E4IP2hfylpT+DUtx5JvCH8/iYny2Of4NZ5E5YAe3U4rot
AEK/zKtkV/B58qwx2unkT/OBsKQBplsJcCrPWwLMVPwf1i2YfZxEHMt9L2IL34bM
HmjMY6HGJY7y608p5qrcVrB3SM3OUcG/znCQK+ED/0v1WQ2Az70eSOpyW0/l3D5G
WSDIOMHSz3cgEh//PD7m68YoQYRCsG2sV5vXWHPUbqltpMmc6q+Yth/SPAAi7hlm
5yjg3JaRfp6V04hcgfD+8UOkT8bAP7fWiMfZMdY6ktX1kA+rHoeWA1X2GOZSkAdg
yiBXPCqt0NWjJisH1fSiruunEITIQhyiR4WZz4OosZ+k6YRubjone3WUYcAGxAyG
HmP0BSW63nkJAWrE66MfKawGmhk0oGya00QPeOIJzBu4YVPBjNojyObM1xGa/qs3
vlsM3l7sfSK4nZN/vbOmV+880cmp06F3wZkiwr8IynQ6l7i8Jg77CO6KZ+5CYOMA
uCgnV6I9T9Afnnj25MNFT7E93N35SoSaOOb5JdAtFn6OdQT1Fy2qKZ99jUAnLdmO
lhhgzg2R0p7a262htQsBJawUyHtDtjkPfiRO0VNMvOEK3Xn11OVs/qh8U1u8m+aH
I+hcCj998fBesvlrIHj0eoNCLUtqR+q8A+ZVRtc6nZ2d07qj454DyRGlGvUumEVs
jUDLOKf8a9ee13U2TViirvJaPKfoLuaJ1zTIhUlDH145rB67Asywd1jsHoDEdv0i
zzsOR9m99xE7n1ii3s0TjMvDJJjg2gqGgAMrq72FjaLz6Gu1w7hNnxMANfL40ME3
T41eZZaoJSXZz80AQ6MuP2FrkaMA8yBtKffAhRccT5531T1mbhSc9HpRgEY06Znc
oiWYrtr4eqRi3y9cDBr3ZOalLG8OhC5IAUWRT1XEW28fACosC5200p8mMavhMUPa
t9NqrcyDQ+1L3lVlXR5OORr+nyWqvqojen6pTELkOX++VgJZY0RWjO+yDbzPXj2w
0/QLS55NFohXmRjuEcnsx3eghA3xF77iVKkaW9l26klepbIh3Hp3zRmaqsrO36/T
Tq4GceQrnKRbfH230vzlHQsvgJZHRli9oKIeJkT+vtLfLLRmWaRD5UCSb4P20uEE
T4txuwOrC63sbRS8SrUmW8xuk6sxSGXXL+bHriL//O9B6hKiu8TGv1iOGWvTQwfL
ZK32VVkZdQoi1xRAsYB3QSyRyR/RTqcgCL4lZp+cR4u8cbnJ2M2wQG+NKCEuT+Km
X88Fmjaw/Gu6+4pQjdDRh1HeVEmW419SdLiu3PUfx4nNNn/y9AUs4KKLR1HkGbj0
mQe+RIOJO5k8pfGJ87i/JwE8pYzlk84byVgVOOTTh/NgzeaaEWHVxCtu8sEw7X1t
3a7vT2c0ZK7x35Pvnvqb7wh+eK33IHMlwZD8lMTXAfzsvjEssWRQkVJwa4YTtO9F
/J7fPWu40cCU/yeV4oU+I3QoWtVyyApgeCwT3U6cvYlpk43MQXsqcOiQr4S6j7OY
8VZKKYfWq/V0VCVobKUrNuAubXmBZu0WA1HWCRPcYVJs4MDAiO/xO5yicKt1HRvV
owyRo0qL9kNV34FkM03My8YkbA3y1jZAqOiVGSEREjcMvgzr2tg6afIMDU+jSZLA
NsbjqaFoYbK4hOKHPnHteEbpDK2+ie1vhBUmI27MqH717X/FtSPWZ7tSZy3xw6eC
96dfr48XOpctRkCPFArRmmL5gVeMNm1Qr2FoFhGyoi0mKxEz5K3+bSudcZEXWi4z
yQA9gTIIgdFSeyd48F9QpH+2PvpxuKWB9AKV2s/iQY3aUnsUKTB9qf1X325YqO0z
z9EEKEMnj4+GLato7WiJZkgHfAYV1IhpoKF+ZQa949aKMLZZrvIKQDz/9/kQXaJy
B81ln3CcW7m1mJAfqqYzMJtqxRRoVJTwbSjaNT3V2/l7s2NsU6CASnpC4D7zdqkX
9YGE0ps9a8W6vUuOEy4rLb4CFtYeOa6tledE/HiM+Nnhcj7Otm4Ioej7BP/5nACK
IdKjFtW6XJamrzSdeMfXQxuf0XrJWZv1xIQp9FA47vg9uEygHEwvUa009763rM1p
v7L8T4rFb48g1IIWiFlSv9HCD7PfxY0OLq3+Sw2OVyw9DagXqO+OVlXWEArmb07Y
IfCLJH42QoRlW3k2ZB2gAtqSWQnj6aFEI/k//eU0f/c=
`protect END_PROTECTED
