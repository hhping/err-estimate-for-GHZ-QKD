`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZ+i6BECzlRaQ1riJv23EiPRlQi1yI9a2AmcCpoHzG46C8u3s72wDGeI8pe77bLk
6krF24gtaVxrbgF2CiqrVMaF9B1d/kwbD4cG7dZVb7QivJ6DPyPqM88rYaxdAtpT
1C9xnlRfQ6Dfy6+QjE6L6uaPgcMXxaEYGmoeG07B3G/P0KEpw9dPAzvNyVba/N4H
rZCMUGAHmmPODuB3k7v/3slH/lpaNI7RL4eeamMYbr1Gb27GrCJ/B0WNOHYGaMvp
khG5laWcm0wu4oqNjEAOoVuusAJXepTb3JFR98bhjCbwfs5rF40Ls09w7mP0dqC9
SOadjxxc38Cgxodcvcl8CR3GKvDNHpPT1YD6PiXrYCy/j0dSefrgKrYx7ObvD+Ji
455oqvkPxIBnBxbduhTc3G1EWFBBb+W+850PZKv/w2TyacRej/ofZYXJZ2TWfZ8V
FjM8wJrPw0yw7MY4MQ0vPqR+VTT9Se2kBnR30nCik0u+LlPJDgrwWKrj0K7gdWW1
JsI492TetVX0e4xW7nRbCbQyYOzApNNvEidJGTswy80jUyZ6biruf7FyAv0rCeYA
ZFtcIFWUWQoj+DSWTmBXtm4F+XheZtfQr0m2xzvpwrK0zYzLi5XVG0CopMlbnB5v
zySSJ9b3/Df9Vyse0SDQUPzqEPNIwBSjSkmR95EImr5vZuMixwx6Z3ZYKh3UDMWa
q2AL2ImnGpHAWcIC12XrTHvrHUMxDOb98gbimIbnszRkE1HC3dy/I+g5gl/swPMw
ZfaYoXV/3K0OptATaSlHpygbeuggsYEWs4g8byeQVG9jq4lTPMEJEjgwyr6Vxeae
g02DJX2JaXkAKOCLHbjDguO7KG06fmrhPVS/LBrR79SdvGgZ6adMt5ayZUukvjJO
o8VIIRxO7H4gEYmICWXFPdobb2c+FIOKlkHA0dd8OoMCxIBR1JguA7J8o80GHkY4
/a2d1Dh9u28P7+Pe3zPgEzFC3OyWm7g7BaJu/tgMkDbY4Jnsy6C7GXZpoZEtpIAQ
AVb8OPtzOxx6FEa35zTn3wcgR/3qGO6tw+xRYk4hmP7GbsntqUZNhZKF6sBa4DHA
hh7XcFD8L73+Zm70igndmOWZBV+CQ2MJCgW8ZL7jlEW2ZrosiWMZeywFGjB6o4Fs
1Cy5VoE7crOM4j3VO9xY6muCTgEVh3416vlwIvx5Dq3IHPqFF2djuGt09Kg4E08E
COt9hMh2rdSJULuO2B48zUukJ/UJQ1jTmSfiZzsPeS5o5HXCkCIFLXOvwGaQ63s2
Va82PKlLpTyZfogP5/uyzQs1/+CREQ6h3EY2XMRGH9ad6ubSfXihmP3de+MdNz1l
MM6owcHoNhFt26xfmpynboARO+2dZLycaSiy4zQGTkyE+dt0s3lPorTcsnX8Hhrg
BVe08VPL+TfkjxLHpG+Wr5Y+ruLSJzH3FaweUQ539P7DC5RnXLV2ETB32Ydw+zIX
La+2ecBqhbheY63XmYT4nRcz/otJgj5zvQGuws1Fz642kU8+AMrCoDhosk1cbNlc
IKtpW9dMBxfGZDiQqOUlsVJqprNf/DItUkFF21fc8I2MGYoSQ7ouaRhY7uAo4tPT
5FJ3oCYJud7LiQy9snfDK8fDqdQXzoqCigaMw84rfyLFO9tAg5YSH6zJqYvmg791
zVeVvwYMs5kxdjaA0YHcPwFixtI9R1/kxGCnq61KES5vovNtaM6FI3zU0zDZSRC+
NZAoH9/5XpQDZmgLEbz0UlVRgGYhJHeQoqCoJDSSTaxeLE4I8WQ3PxB1drKdqigB
1wikpoWnRjUYe3xFwWVEphYjU48skD8N1d2AkrFj4dFcf4lUdTtqdUz4dRi4a8Gx
WLVWlmOsDGVYMrocH+I0ypapqMC9GhASHzPl/xnUdU2hCJffpImlfJ+r9qx0LRMP
bbSeOX+PPKw1eKdI4Yk6giF//OGnzNaVGjrcHjNW2BPk0J5HwRV6coCfHn8s46Zp
nU8S4oabVYxXlwxCI4SRU0leZTBDaqhejVsWnIlgCvGKYlOTaR7qMBhCikRBLJay
o0bKsQO/VVXNrzhTOPaq6uZhNONnzau/h4AHQLNi0Vp6nS8slyMUi2G14rKZkIwk
/s95ZrIeEncHJm42cO+B7o+ab45drBIxpJpVLXKcdZjYfghokteeDyBnYvzAsDny
pmIgiAYOwx7qKJHSRJOSbtI/QAcrkOF04UVSqOJ878zKJHDFXSoIn26J93O7OMcf
4ZVdROkMEdpKuzhXylBgig==
`protect END_PROTECTED
