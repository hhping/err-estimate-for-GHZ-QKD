`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AqJIrwKsAqs+94FKemeBXpDhNi2leESUMicP2tle2fzD6uogdxb0DQ+6/F20WUyG
YJUIxE0m5UaqjhCPzbwccnA+6bZ2/8mTWu2nLfPVHsgg2CKYJAYqR1IJfMbwxS34
UbujtLP0UNimWFCW8JGlWjnb1LL37+o10IlgE3TCwcO2YDVy3QoW8U2sy3f6Y5Xw
LhLUrq/vzfxyBuc0/LBwOnVz03mH2jLR9kQogSB5RktLwwy9Jkt++PfXxwQa38z6
fZtZpeBTlYdbpzyN7efLPz9gTsojFx+I6OjjnP2N56Mvx+LM+hP+3X1DM6JJpkqC
8W3SayR+gHC4uQWJnzJE5i/Z+sbHG+x6H3ThevLKs5gkyW4hea2fHse2khju/PgS
LFVWzwvhqHEhFF0hug5n9E1eF9z/qH/pwngGXPOOJ12r85YIHr6vgoveQDVsL3OE
389bQhNhI4BuwJAWXymwU7LJcTzmuHheWti/ZG3wP5ajfC7qpoQ4NGb6pT76efbQ
w9xNwTdycmS1bLYWUiWz8ABBQQryrvk4JfubUQ0SvqBoD8czpM25cVBayOupc8s5
Wspkf2hEr4N501aTJzI/uYHLBTNMu+j+vZDIEaJ5XWXrfwwG/FbJfixhr9wjGw+l
ZgDFvXnfl2sJIvVcowsed6sr1NGzVVZ11IsGasld/kirmpyYQ8ZQwyTgcTcGVwtM
7pyMMNjPYv/59USDnwdBHbUPZa15amNVW43bbbud/Mw5T6EgkWWLISUIk4mSdJZD
sMxP4r8Q12hczBX1lXvUfK1xdqutmUPyA1ka1UPOELY8XPKiAcwUEua7mQuU352G
cTDcuB0qNtnWgLmXbhl6YYNfmi1+5e/ORgIfKiKkU6FIiTkuJ3z5eSbewuQLac9j
cp9F6WFPwOUKlSZYsn9ivfAPeNUnM5HLsQxffjM2YZ9IGX1xQNpyO5aoXDFzD9i/
JYrcaYXln7yVheJr7oJgMtwFTTkPDwyAriCpEIjvoceIQN7xLqhBFlSLTrOg+1jN
IOvAi8d2WVOuPtb9dUI2rJuYhliyuEj5yKpVF40Ux5gVM9dbR2WL20t7i1y99SG6
RU3V8WD7p+WNsTj/Qu9q6yyxUaF35QbhdAgcUldCRXn5pjjkJ1G+CUVBZNjUfrhF
aycwH2NFXkltYaiHMgXbkSK3qByrsbHEMMucAt024T2lTV2H4iSECekWnAakMF5/
MaudntD26Q7LkY164nz4oJ3yCOs1dxgLxnq5THpt4SsX9zVzCZbuYmL5/17ynpoc
GBEmAwY1le3CmFwYkaWLMqcIqIBxYsRinHctD7Uhjp+7uEQA8xt8ZuLgP3K8jdMW
D5mIIVNOhj/f3We4yCDZlMzSX7vtsEBo00alMvuVWkB+8l48Z6HA2c0Ew3QArZtV
9f/AKhYceeClnnziT2ooDzR//g7iGCnt98mTGrphK7jfYZLcvqbiXYNmqo01VGMc
`protect END_PROTECTED
