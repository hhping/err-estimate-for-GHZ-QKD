`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJBIzH4hQnS1XxJ/B5Uehqhr67YFxQUkevE4B/IVJhKNpXpRXGXk5Dv7B8hmMYrL
OVEuJT9RgrmpA6J12kRZPmRlcev8FxjwRabGRc4WZi1aTc5Ox7s2RjFpKTTQqExc
4nx+eD4mhD0fb/aUT4vQeF6v5peOtx6/f6ZXecBtj0rec1JV8XtKOAr3C5jBt8h9
JpbSRihZQxVi4oEoRSojXrk9+y9SC6E04bDwH0C3bKLorkpevLUYmaTL5/4cpHPF
Yc7x87AHMcn4tHmLBoLgTfMWcGzLgj6KUjoZe+1581ilBpHoEq7t7U4BhnnIJH0X
KhO4A0HSVRaQbHQnVEDJinDPySlgNfokdC+M0HoS0BrhkgPqX3FnkfKOEFiySv6y
F4BIL6CRL4O5b3MvWZOIJzjoKE3OmRt+e7B2TOLcV47jUIOjMLpie6A0yro03kkR
j8+mVFgjzbuA4mx4Ry8ybQMedKaJyx4SY+geU18RRMXnBCdShMs6UueFmWmNpDuf
h7L/Ir0iiGbGQcmUQs9mjPWKLUCbZYoW21CACKOKBG0BUof0+eKev0YFzB1C8K4s
sYHgsoR4cTbHPH79K5bF0wpa076l1Lnczut2fV8uPKS5j7qmdYvxxDr55mC4sIHF
NprNLaJlI9VyNJlNX73QEqrcJEwRVIq1jmYINEUavHG8xGX5VGvN1FjbhDzFtQJG
K+8CtvuYkuFzzakO+WrXifWrYRItjNxfJn+vtFny7MiXg3EzpF1AaB/+8UXC/3vC
2b6MmshD/uJXadqtTkqX2tStNc3jgSS62RgzFn9PdEdcT0OE9BZ+Du48/5fDEYva
t1vTDAIPZB5mANB7NhqJQW92pGNQUikzeLCYnbsi2vpnCzyA+jN5u6b/VLmPZAdY
xWqmzHcwc+FfLao7GE8v+zmtoA93zZZCjbdPKnTW2ZjkNlmZbdNiWlDF9Ehzvs4I
y8PlQuwL6eePscuE/yPDR/lXZlYqUPbzJVFD3iG3Ca1NAQUS+NZdBZAEysxHnNCP
/3MStXSzO0qIIwrWlTkgyUU7EPBq1Z/h0Jefsssv1bVzDvS35RQ5n3UYcBegX7vr
bSkA6k4s5VWbNN+q6TDWienz5WOzF+NFuuZiqKLS6CmD1yAjatQy47sKg6DZ1uZl
oO4xIviwPzRGkVtmfOWey3meMLmteISyQ+gFydqPyBj24pLDKja25hCBQeBhDly8
WZZ511tpDdRCbekg4i5Ra2958PnE/skZkhBK3ZGGXV6vymYDzpCZjGjCdkue+d1S
sa/XLvyd67d6dZKDEwkKRcgkoF/hwzCjqLsXSOY3H/4JTUTExPGdGAFA09JZ1PxC
PZMFShXsUa+1IzTkIdgbkMNcNWk0KguDIdjHJAcGs+2JiwEc7U7fhMfLY87GuLeW
ywWY6ctJOpNVb4L5P6Jwdlgd3YJXjWmj3yRyD0y16QiT0qds6fPAOuWSJ2AhuCNT
6iVSH0D77TDaLGbSviIrdNfg8uj3hKRD4LwheWGZ0XzfMK1ZMT1KCl7dK4B5abuC
iLAs56nI/ZO7eUPpRsKc+DfTP9Bp3DGT/jQgFAhFpv2ApSOFhR6Atj2vRZBQ8i/P
I63Zx+j45Hf3i7xl9EWtyObCj6IeGGSGNQO0Q/CuA02us4tlk5idC4EFwzYqOpzl
wSaXWTHevRlOCc6vH9JKImeaKXyuWPyHuvBEZxE4j2Cu+CYnO10ABkI+RWjk2f8D
SEIfC/tZPpH6aTpgkAReUlNpItzOR8WUCO00dmltihzqCwGWO6Xst87THjDhNb29
WOhAz0qeNvE0c//jrVbTsrqcrkkSsqeBe2gD1xETdp0QbP0SiTDaocoaf9TNNhe+
nuBnVzo0abxriMub7brHJc0igpCAiTBiKJvQwqf6RnQWSKwmx9HFE7b195oKXTNR
ycMfto+OtEkPD1Sm0PQB6wZSfWpWQegyZL1F6y72g4uwrVAPBTk5DsETc30dTplF
CeawKVaZfDXmrQLIV5aE9PjC50Z/zuUddIg2Gi2QRwSrv9LNd2wbBawFEkvEjFKw
dc89hdGTxmF0GBltoNjeOBLzrBfATpWZ1pZKqdIqDNw4NgKLFikVkQ7M/M+w2AZB
pvwkr8HYQ9E+oTUnmrx660flZWNS/35gjySggfFcX6moqsdKP6cpyqbPG0htwg3O
e+fTgYh+8BeP9PEMpDQVsempEN191gd0K2WsGTogCHAqyIuY1YacxgDUd0iAjkRw
Dj9HQADRRFIundfGfIKoKTebgVNk8b9Rp4rpY1swMIq57JJCTjytUHhc4pThN/jB
tQ0NMYuLlOLTJkxvzNZtGmieDkRKpf4ZEvE1uHa+WDwjSQWGNQWxlzTKsY+cxC+M
fz0qy4QNYyM8qALD2UfKh+cc73VBTM6TzqZZHkhKXf3kA1UkH+4W7d/grtX4F9y5
ZJZ6xX7D0EjW2ESdRcjwWXRXjjin+T+qTQqJ4dIx1afuDkvxTsp5y0vUu9WWtsKK
Rcq6XFhPGYs59RcSwTwKEm7EyPQvH+3q/T6Y8Ij+iiVIfrRRX2hGfHWmUKJYUe/2
KI32nZjUqCLoNKAVBtLv0U6kIKrbQHlTzy4v6EBqUA1vlgfPWVI0WFYM1XUXc9R/
69dyo0g+hCbMDUCY6zwk0qE/obCYe8vRvEaRMUv6OiEa5h+qkQCOT85GYByM31b8
vDRd3pRGTFIUkz8wTbIJLT3XdIuSguz6f3is2krc5cLPGAtVj4bSttxEQwYQNRdZ
6ELY4oMW4QYKJtn/wLs4nD3mJxc/ML1lRR73G9Q7iNC6+trTAnAvBekAPP51rpU5
M+I7Zk+kGlD//AdsV5Tcri3HJTsr/jkIwXSoy6+MHMcJPYQeDaaFUvw/BWP4c4jo
IRQpGYLNAENRQdL00iH9mraof6m2jGXrYbfyaWI8goBIuV3dyv2k1YzMGiBZ5sfB
lAl78JllnuifcNyLdBmWS89spwzi9YfwFcAVPcoDqStGaHBXKXvWmLybT+uySNjg
SG8uiXNg+y+HZyXZd1UskUSPIysjzzOptkX6jdKkjN1h1RZu52N9yZ4TbJKm54ZX
4GOfqo5wAzIukw4WNQEYFS+P1z72d2RFe41aMdPO/6ldUXCw4lf3U7cDMrp0Q0FS
i1zLJBrsXxvzI5NLzEPAbs5xntHy2CZqwYTWMOkbc4sxhdLq5DSCe+s6AQDaiuFj
hpvuz2wFg7LaPqFFN0sad7FYjyLlkZnG1BRMJeLl6DQWnfh6rM7EoWBcAY/1U/9B
twvqet9xINaU9fVrR9Q0/DQVDyhwbdy++xa4viIorj51r8TegzLFbz6FEOqhUAYa
xCXRcSuixSFmN4HDzCDYaDSKX7aFtstKNV48nis/JDo6M95QPDwSz4dEZ7c8Fgpz
O7lmk6yCFRxjfFtUxEV457Wn6C5vQZLmNgifElZzbdVB2vrLqvdCK15AWraKVOfm
KnXkkPIRx4/GceFyvG8jEYWtAY+BjW3g/bI5Ywx1gqaOIobmRgKesyOpo6j/LPOi
eZcCfcUBxWCpCj09fs8xPa0BRosSGB3YtkAJ8UfJ3ux4zeeExj86niTkQvCb+HJ0
qv1bLciMup1OoF8WeferYGXHK4fPTIDdEko5M6broAw=
`protect END_PROTECTED
