`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wkWjwKbRyyV63GeFoLkyiNAQmKPYt+ZOtCS574wLpIU84C9mHdXbU1pxccS2+rHG
OIGnyBvT+lCspN/lqITbuzJmbxIpBdIkiLDukV7rj46UrX+tPxDdioJl8CFV3oTM
3Tlx6HmUUUGHH1onzd+YZhO6cy0oClQLtNOy9fqZur/wynSAhtNYPrZrPXXCq9pq
NXAy+g9y8iB4KXZaSwyUiDflCpWmMDs9Zc0LGLFDfHJLbfT8i8kqtcS6HahZUDEc
8eNYY2ZKogLGssTuBhLhpH9cLz8nlH9IRXWdRLTNN/ZsXTknXggjHVZvEGFYBxx7
0oZ067vR77UarXZonpjX16Mj88V5uwNSR9kBuzIKHtZ6DKYqEN88rc6C4OKs/1HZ
eOO/Ti/DatJ2gRKRz5NjEdsYQlesFG/Va93Sz8Amv3a4Zfp6CQeo3KAr19Qj6l+J
uuVFrcQj+onwp3cQZD+ADncalUW91ddsLdppq5/zwIiYHXPPusS/Jy5KHwW0sLVn
OzBg7hgXXQJ0dqxzc+lxdAvlEx+d6tKnIDw0no3ycEe6zYcf3BRBS1D1S9Lkh1jO
SSmd/QOnFsHWbLY+DjTPF66t6U5riT+s7kcXftGN1KWLN7v56a6488t7ThGvtQhI
7nQgjr6JMNht8uD6RLVlahCxIPrZ6JowiQfTLGOvDYc7ETJVHfb+C56z7G6YXMPX
bnGUS8G3V41egmGD8RCLNzWmGB/0rTavKSoNZhU1CE2oOSIcKy5lPMTcOjWgskE9
7XcfPYfthiu/gGXmWsvOCHUNFqnL3WuS1S4YZ4juUmNt0KngTajl9roDPS/9o/3Y
QLG094vTe3k0NK17wV1qNA==
`protect END_PROTECTED
