`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olUjdDGTb4Oc0+KEEy44Jl4O2tNBdYH7xnQlj7j+FVD2oQrIBK8BxsBx2bY8CYGl
FXrmHF/3IGKleS+UaiCaMGWv+UQhCnuZt2QLuKxv/DyNQgkMaqbbjCXtqvw47u9+
D9fUVm/Z7ZSoYpkLPQCOge+8fPeA8jrXqkRa4QcZFTNbM5LpbUdKh1BazmZBQNjJ
YaIlfSg80Q2sErnL0ij4tcWXjeV/TK7HLwbxZgMOeVuptEL0mZbXgg72WgosdK3L
hLv6qzvte6OVD3NtdaFsSHO3EKWA2ivTIPhZxZI8nH/I0rTHSc5z112PA4AWbIwv
XrMWqXOG6eSUFepEUNGngtAAKZ+pWlWHShwDYvn4snkAF/6KufhbfWQKTEk2oTe3
jf1/JLgu4lKyRr1t3XBZhkQF+A4++fY+9m+rWs7UxloxpZtpvnoJgypnOsGSPieb
H/kJ+OBlmW1/sGk68zPePDQdE2zGhGz8WojzVPQoyrJgBEJF9mVD+J9jDdaDHJBP
5bN9TSpTL0x2zv2EVmE+GFu9gBaUeuKqsZjBD0a9fzPn+rSDRPHon6hiu/QFEtez
26jLupJYndoIJE/h8WXoVacqIErAnzKPl1AEQlg2rJO5OYhtF7xbYqsdkNW24hv3
uT+Vq/+BagzPIk+ufEAN3KWWAzr5QwaOqWGl2evTZW+/aHtAJsYCSVHQC/079RMF
N+t4/7y2mmcQ3q0QQ79FU2i502wUItlguldZc1J8TZ3D/VTrmsULBsmTKO2h7tcj
xZUy6e81NC0GfRZWw6oXwxflkHPqyQ8KTq0NfyRpIFOHTJqO8VfeJzPvNaYOkZoU
YuE8UxKJXHj4YL+N0aBcF0ud2DLv6gWEs/AE7CnKgJJtoyq6eUDWWoFs6pVBRInq
hxHLDe4xT5keHN0OWp5+VQf4keaTq1XZMjIYvaqDP9Aj+f+EydRdExxhK9aMCww/
Wg/C8PYKFnrsTTdi1mSnxOXWsFYm84G7FayrEBVoQB5Q5XZMoOlzX3eeuo1oCYnb
qg0IroX+KflTJrcfPx+0TQFSMKi8wFldByyqQUjEePQv50VDqgcm07lasoG04e7l
yo46Ob+eFw22trIp1L0L7u0W/a+QGLhwxuGXEf43fB+4rNQv7lJzZMZIQ56cq2uj
IpzdCc494XClibVd+ITXP7Z/nC1XXb2AgReuiWaahE3snEFjnVzlfIj7K6stSM3a
oy0HwlrZU6vinB6y2NQbsDpnreeLwWy97R1QsXRxD68yLJyUcYrmC0ypXs3FBw5s
IxQpDT6w+H0DjwmE/3/WTAfgb/Bnut04GYTxEAdNr3HD+pqKtdUg2SeSjyPNoO0N
7P6XrViC/bendVh7ECVOyvYjXKBeTPxB4W506hrmGgIxKjzCVE/QO6gzmPDM0hdt
nu+zX7aXVhHJPIFLrJUm3kQPAUZYSnUF9WQBQuAQHFsCfnG4Bp0CUpSORuluzpnt
pkG8Du1mhJXgoK/E1lGpifyyn7arMJylFv+hIV6ujeC7pV201k6KaYy90k6jsGLG
XkDOLiJyxI1nKfXf9OwSwCgFxoiq5uXE9LT2YEtcXS0tZuLjrEbXK8/7OLqc4a2w
CiXh21mPUmA5XepJvii6lAIbSQS2c1B328cgW6xTt5izEPyrkjwHD37D6LHkWxBO
fqMVd1xvgJqO35wHGwcy7kVwslLPi/0JpARuXpBGvAvSUB2mOl69+RIxVwKMQQKV
52w4PtgQGJiVvYCljqBa9NEJRXok3TjO/G1xJHKXriLcfr7uHaMUCMNnr1hDcSBB
c1pM7cGXX4zVgyi+opywRHRFfR5hir9Dj2/NL8z6O3Va0n1a8ep/Sbh+hf4sroGH
I6SvIAPwNiYgyrsa4ZlwP3YsItwyK6WNnmnmv2Syu0o10aLUGBV4sfMuW+QoXfld
jHGyMYH3Pu/lb8irV0kxWh5F4BMJiGbZkPlRbVWdGgPNu3CmfcibJv2at3j8umET
JzpFBnb1vACsWzvYFcJRuJl5jvdGgWKtRYu5INuv73hvJbzZhaDBgchZUyRUOpQS
1cbTmCU9O/iM/qJKReUl5PuwApma5f0pAVYTGlh7bGqCQ+Hmc4fGRnPQUX0i+0Q7
RhITwl/UNmQLaWs4UbFqi9r9/zWZEmzHPv7FamLO+dWVoxBJFfCIM7chBpVS10Na
+ph5Oo7K5k4Xe1Ta2LpKKqDvIMiz/hrqxdkb2KUHu5vBpbXyHMJU1bWE4a7WOdX1
b87AYvD08/f19FdmxW12o3gU0g677XLaRDZgCNd0B+CP+pTa9WvHwgU0yKEZWPUE
JtkQwI3uQw/NPbIV1zeUeDBCOCUkSjxoywC7mc4L/Ir2OUgRz8aQJXKs7DLDk32Y
ct93tmrNKWekpn8qCKw1nrS/8uO6KcEIDp7mByimOwsLh+yLqN8VbgvafWIgzVjz
7KFu5rFiEwKwYPbFyKCwRmqVYhlS4/KU4IC6RpIEM5nevBSqLPV2M3x9oRVOFLh7
GfKgewgqcu47cdtzuNmqMbWYCNIFpdwY2zj5pxKz+4NTozpcc/N7psrMxcvrflsO
VfPiN7McO/qZRcOv+ypKIr/FFOgHQnZwUic1YKGUbDstaMPwDcRideX0fyiEy0rq
q1kRKtYGJsPCpmdRkEgvJzDjp/4p7/vJOgpr4/8NV4UV9g1i9/+V2Gp6NK/+S480
dMvgvFP4xseEOPrlQodqLAJG64EYeBHmwXr8qdcxl0pAptlr9z9coalgWhtMYKzK
5QsAO18UY9NAtLur/pxcLGQ2yGJKUNPGxcEvlctNZDe58e9mxKduwOWdXa9NJfdW
5y187hMi7gZJB/4AvPojoxTKr6aiHYhizbngKZXB2BpCtRkbXJ0QGzAjSDQs9c92
9YdaSWYd3JRA2gQu6VfXRWe0hwUU2byjzkmqNhhOxLOD0OwJtPPakq0TDg5+OYDB
44LDQxdMgXvUcgjfLxoQFT1bsI2UbMxGLceuIwuCXPXHp+arhg2SPOh6LkhaySQb
cN+p+GtvVQ4oiGhFMb30KvJGyS4SzbwqHNO49vZfAQIQuUZqcbQFsRNcUOSHmG+m
5abuXnDGU6MLflzF7KPzDHapw7G2C94U8kGgOXzUimNm6+8hxXftjq36mzaDSE/h
7ilbBl6cAvsa5v+k3FFJuFbd1lkn1M+uGIKNMFfaIlTf8xP7L1smtegNJ6Qam8Re
RSPveVQmp8jNa9Zsyjp7Sz1nZStFLt4/Fcsyfr5cfSzA2HVGBpVzNOMxSfvi8U9Y
fXdSRN3f3BIinFRtpZcmhcruks5Fgy3462x8+l+umflvEhvrl+5XcnWXLC/CAIaJ
MVZATARcSe9L0rhR7BLfZMLSI28FlWDIoraiavgCns+aFzb5ZaLjbuFUfmqa0FTW
klMWMk9G/R9OouklKTv8gFNORabtB7IS9OP6A0ZA9ADrDR5wPyl1X6VSQc1IwQ78
HCmrDxob91nGWA7WcOK1AmxHqp10u+k4Oj5cuOG2W8HJ4+86Gcv66c3Hp8uQQipt
Gn7rbpylkeqflaiB5fFiuB0c+LHmvDXfbVlVF4k+mAjSVC0HatBAmuR8bP+BCPm7
7Gd67PPrVjQgoubO8Tj0gw==
`protect END_PROTECTED
