`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nN24l7OA5TilSwgMskpvI8UogfTLneCulfEabvBX28Arpi+H5T/YpR0hHwWgwGLC
zwhkTq4/W3O+Zx+/EtkeBOmVB0mC9aRaJLHCidsEKexP+Iin3/tUDSsOZUFvjpff
BuR+GwxovqKtzqSTMu2Fh3I8Jpt38UOK+RbtrFsdSYVV5F+rz2hSqnd0wwToF0ne
HEjx/EuuuO0yox8do3JAUt0g5u+1qIrZv3AXUeNjOylNAK6mJnww521YnTVhuvWC
KBM7a2RFgTmoJDGFujmdmk0CvV7T98einWDv4zLIHolJhFaA6NM3bLEP8qPvOPoq
IXvSRIiqRcMuIaAZqazvb37r53GzIvPsxAR4VKYmy+mOIWdR1Bhs3yMykDJYZwzt
lzGePbEPJ/MFeDSU5+LAOxIzNkHgy7+OSo0ZS0texnfIuqHOq0nk6J0xThgoGdut
2fi7QDojmJk2WOMIHjXp0ZLtfO+TfwM01NyROsx21j5pyOkjHMkytR9t+NSuiEq9
LO06168TAhXnEWP1De9UHUfM7dEnK9OoJMo8tuwBA5lB5BpQTyzHfhuTaA3Q0bDz
nYaVGI4dZC2GJEuq+ZecV+OwMRV5UZaN5UdUhey5BFT4JqpedVmGQWJx0M83OGBV
q2kl0X4e9u6s2WQlUeyJkbSn6K6S+431/CQeFDqnr36T0yJWsTXWC+fNs27McjWL
9Ta95nl0c4Q4UYk5LE1/38Z5ygYk09bj1QS2mVOK4drI3rKSMaoVWuMDpI88f6kX
TiEWiUvpWn8hcv7elWtlPiNH1xNiaH28ItfDnvbYZUmjTa3jfu/7X+E1bPYHGogn
gR+dCBAnpAd+tWPgerzCHN5bG2iJq3RCY6KlHRvtmoBt3/nAKQkLGlfVkouA/RQx
Peo2dA2Bp9LQ9SZ9lkOgAeRexb1xrX0On/IdAUiUTXAzoXiJG6FHsBsetklI7/v6
DC2yWrALpQkLDj2yduQAs1Q87HGraUQquFUX8ML9fUwO6NQhdGVoW6PBFVxc1BJL
InHnuMllhQdGFMazi5Xjyy+WQWVxme4xmslh1S9ZIImwTjsjDz2Bdg3+M7i8+jfn
`protect END_PROTECTED
