`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X6dlyTrf+Ht6HpooZpncDvJO46t4CvotAEvKU4I7NtxcfWRYpW1Jh1jARLRVwHqE
NlsAPSWpGH4urmHVV3mIocEKceC48i9B7ypRnW8/YA794NfdGuMPhyQbnRAe4Je5
IO0A0iktUKuAqtPeSlWKWoF7cz+POHQcgQA9TBZ/j9Pja9i9uM2l72Vkg84iVg0r
vbOX8MN+JvQyfFWRzASBhKiGv9/+1JNlbwpY+75K/Qyc+H9BH8ILWRBJcYfCGlhU
WRxACePTx83XWFEE32o/8kozSaczfydeqA6G7vCZW/SIBaYkihNXBOd8fUdmd4Ij
cwVpXKSW4+G9V/KcUztbVmcKIfDc6xwMfP0EqPzsCL5PBe7tIm1/HQRoPAnVKrFG
L+YxCCghjr1OPmS7jrtDr5yxvTH2+uPPLIAK7iTg4NyRmSY4IKHQB1Fh7tGX4a69
zCqytsVA/FRdCRuKGeenOS7d8x3XlpsYjPcmECNJ5zVH6nPMoDddiZtoRi8lN/zg
QHzdI/TRs9CvaoPRJHbswP8P8EN045m832lYo3dQTz9dmbu1Rvmi7dtrmuAu/IRZ
kCTMbRpwfft/FBdyGh5Cbhp0c4F4kOMxavy+ZqyJ9BEaeKLtEcwbceBn883vUxjf
nYUugO0Byej645ZI6La0nHWXvoIUASby8ssKVsT54/oZ6fOKV4iQxsfzFi54oqQb
aUctbsqKspgFlQmll0CarBZQeXHn7ewnJ1v1gagtgmDkXKWsxOdV4ZH4hY3L4qU+
BIDJ+0dTP94Sxd8YaEPRlbTT4hzbIA4O6Og2CSrqFEuBXesSuZsDW+F8udTDxRdn
xuXn5bZCdfTTCzxiqExrHTtYXPi90dikVdHVCOvIU1GOI4az5Kxjx3YT/h1efLEF
+0GEJ/TmJh8rirndD09oPOkywjwfmM40FFAsnCf0j0DPid9HyD0+qVsNG0icpm2R
l6V2mKU0m8j+PWlLMEfVwSSO/qWwd3GRUE7uOC+HXo26kR5FJJB23Li19gFn8KMc
azFU5f+LQeSlxr/qKEarDfCswtLHEtIf7lk/2ek0XfjHbDWp9i8r2rXsvDO0zw/M
mNb63HodkaCF+ENhmuTjWQ==
`protect END_PROTECTED
