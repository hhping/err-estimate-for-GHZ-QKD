`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3GAe5O6wL7p6sc+0uWBq2KUK8MDQCq6+uzBxdTMhaRfa3c6rE8V121wm6gFGt4zk
50h8CsRqtoFKW1blLnPBnjAMjv5tSgkKC+KeDi0TedxzFH45V3huRgJXnfSp9kzx
8aDS8Dc0XuO1l6WnDv5HiZsdiS4lr8KKjPJevhKK6nZRwch3hWyl5lal0HIc9AM0
yTaH9lLjmV+Y9SJ4HlJqn2zESKDncoqUmVzDWA4G8USic08HAKCtonThB+tRLyDv
2SMxvIOBX5Z1zdq9QRf7LcLgsx0LGSis/rjs5JBgP/HXbk+HZOd9grfDa88X320o
mWuXEXqCA3lO/dyRpA1sTFQWNhLaruJ4X+GSfQAIj3YGX19zSAsbcVZA/2yRRYvD
G/NkmzvIhpSCSDAJLq53rstUh1ZX3BSRz38PBBkGQtMtAirdG7WoI2TpdrAotYsC
ec/i1FRhCmk/tpNhuAzmo+813SDxm81+KUp3d6R3wQ7xjbYvNyQ5YQdCscE2luoh
VNCk5CzdTlWS3tZ5D8tghXPLpb0wDffTVeEXROn7AfeW7QrawEXA5XiEt6ulcgu5
nZAvhfi5PfeH7bNORc/3AxXbyixji/WX7GX4vZWJPyzBwcwAzYZ/jZSHuZQiorOJ
qCR6+UKrGtwM/NdWNlwAfkzLrQw/9f14eec3aVtS4nV9zd1S0SRBiny9gpdSgUdy
RemIa20F2msX3H2CIQnLLZzrhyVu/rMAjtHE7dxb05cbHJYIXVCr9HoJI/ymyobQ
BnHz7cSf0UMY2QOzzwQwKwraapUPqAyhG5wBUZmjvJQt4fEOeswwH6H6Ojdg91ET
zzUuXvQTezDlMC6gxWda+Q==
`protect END_PROTECTED
