`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBisIJ53svHmsf72CySX3fSJ33HvRE1YRjAUPdgr6hjDqw5DrhwmOG5lFpIcXXdT
NJDa3Bj36RP7bBh7NeAuW/hvT08M4IFX/eXN2dOfRuMjMAxYAR4QtCza9lQj94po
qn+W3F9qFRgh6MI05U8N2hjcIUXZbdd3fBysyf68z2GzkFDAGiES8QoekF59fidm
Xlimb4A1dOyLC8oihplIE6L3s4SLbEcUpJd+Uy+fZvclwoXSOos7DgypMIWLpPDb
RMlJCSPnFIHoCs+zRJRiG1c5fhIE++MxSOut8RkN/KKqwSDAwdHAELDh34edad2m
teHOu5zsNavJmd52J8bIssgOKNvXBBYCfLjDHHOujYDyMrBYhBvifjOeQXdOHBEZ
pSJ80vVj6GSxevRQWmrvZ9T0c7GQbvGzzRbY1zAEmFp/TAby10LVRYrR1+4JUgpr
oPRSZfV6jt82mjP35S2cyZQMtIkig8iaUAgrzs/3I74rwJHNIngYrKeVKd6/2NfB
c4S4eXUrs93rEYbB8nI0AgdFgISIasTqiQuKad5TSmuG3rI7swN/mKkTEyJfGcT8
kON7ymy9wmDyu4YPLAAaKviwL3LAGoQ3jBM+v9Ppocxz84wEmTUJatpbsWlMoSKk
tOuWKk33ENztIO7azSIozUUWo2G3mf0aWcBqDhs9W3oBh1KHPW8ktl1gHx/f31q5
6V5RJFNfhV/GY+tb3yHXCcEYM5qCQKSGVoHOHR/oncMY8LGulSuLPQZ21JGVr7Rm
bKP5rOKwFHbS/4KHTOqtTU69f84NaycUsnDzBPXcYT8FlZ17bKKXkQF1e2gvSL2z
TkS1LD0Du04y2+skiE9SxkF62djK6Ex4aIlqqV2K9kxnBtZol+EdbjGdsubN66G3
4DmWjqNq2JwXTXLSpRS5FubtVB9mLn4uhL6OXcjp94HS+N/4yBlrPSv6OKiqd0Yx
Phhlye8+m4ZMJBvo02PV1+eGbhOTD/6YLnebijbRY0QCV1mZNLadpN05lh6YxGzz
g4KvnJnIj1GJK/6eif3Kx2mHliy0nj7DeU00ujYxZaLWELMmOGyuG6OVOr2Xhiac
6msBQNX6VFA7YGhpicOLbNx8lSqK6ocQlc/zADG8zRVBTJVIayE1DVUxUA5Rcq6A
dMTm6tGiJIVRzNnKsbKP1W5zmtPaP9fYLk2P9MsFiWXwhKxdsXfoonNSdZhZAgyR
fXhGcTDiSGnmWJ6ghgRlyv9goY4D2ZeX9nxzbgaqICK/NSNEUuqVhGOfv8jcIX+z
5GAmophX3vxLdpBQFQnDlEPgj2YgdWjLYyalfN+IHsEb2nNeOYnqLlFALGWMZ/FA
mXCycpBq6yZw6RcTRIh5vq5MLGTWmItq+sY806XRn1fpgoIxtrRJnxnPqij/mrMr
PTVMqK6UsFcXBkkkNbd6hOIBkaWIF5vu9vbJ8vFDuydPyvY3hdZV+Fr4Qb7hQjG5
7biIf82rrTfd2/4s4Dm3aN+46VhlQT0k2iqBBHA90/D1FlBBIDzpzECcrXqqAbSQ
ODwATqbFUags5bYUvOUQLt+jHjNgaKhFUftRNzqUkRQU0iiCt1HKDq1TJ/N7ntv6
2LAONeraNS1BYfR/pwB1TFtXHYKGpba3EOdfr47p6lWp3F5wHu3wMgf+8Ni67mMK
gVMzWAgEdgdDtom1m414ZhrXOF5Yxxx4+q4P0iJkhzqrlfCqYkwOeKuJ8liO8Heq
XpthDh4zSfGWGiJxuPqzZc0gcwaOazFH1Y83qrMh1JXitQm7d/7GRWJIQGvZe6tF
+uRNlKnZsh+G5VW8sEPDISihg5ade/giUWcBJyw2cL4NcJ7EoSpFfwelA1VSF6ct
QGkIjZcLpUo6/LjtxfLs4/Ejc8x6MEex6EMqxFe+g1fACviFOJWsB69mEUuU2WKa
LfcRInC186OrAajk9DR3WC4laOFyBklZy2k6WlPUUShzz16WxMvcfNjhiVXx/V6s
`protect END_PROTECTED
