`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcoe8E+Cye8WRW2v0g1go7R7ZM5smkhLxE5tUgrLSQkKhH9UtFWGzhfAnYUpo8fG
E8wgZ5hMM92aYUY5b/SZxWYU40duuA/l8I2apVdPKobcEO95a48zQSFZn8BBhVI3
QaubWH8Vdm08+II3FQzgGMwAvO1HOR8XrfuFPCkKVcsjH9gvsvBrsR5719jN0k2u
g6lM0lPfLfOP8aqqQymA5aqAzctPtalYByDyPIYPnS0miq+ULM/oNvxeb8Cmf385
jyVId2xLujjX6eTYJkUJWjlx5OSGLVV2dhCodpzqI2rmNn0VWo0MzZVIG2oEzlmG
QJbbL4eymkgNGZd0ZoFCmFJMgY2nfRN0VAKagQeGG1mmNaGe7ZWxqmd7KsDUWTtt
cH6vRkXFUjBwj/cohujzlMT/cSG2NG9bQqRF14VOwUbBGLpNHmUoe2l4Nyuj62q7
MA+IHDm8wbAo1K0idc7GeHA6Os4w6Ochdbq0nMT0187VpMJa+XW9ODQNS9SD39CV
Y3bIQvChbztNemGtpTMXIrTacjOiKrvoedlnibfRrhnT+t2fM984EsZq5soaS7jK
A5quY22sB9qHXKMQRCe+hKrSVDDwgC7jMD9OAicnX0MDHEhLvSLZu4KWuY8lrviL
5THkawAnqNf4joTriQOEKAhQTOqey7YZ9SfOufS92PlWrx/Wnas+RRCqeWEAuBAh
dihW4/sF6tTeuUCRHdxBrOrM+rJUR874e1GMyJk3ZahHTcUMOJ6VnPidiJJCXua+
CBFCm5qpAXEnrlWFI1maHyhp4ZNINxYgHflKgXLaz6yLW4Nwy5PQoDfAtoU6RrNf
NIB8YEXgoa3jt6MWTe9vL8vX2CK29V+0PdmZMM6SmiwphCCMJhRMoHm+Zca4958B
vHSrv2a0rtGAv2dpCWNsf/C43tjCRV0A8G3my6aNChXJk8j2lidp2SRgjYWrawVc
BwH3SwfjX6x6EIKk6tgRmSaA2NV3PavlzN1d+LCF/V5tfpnEy+r35a9Blbgsmh0n
nrNx+Cz37GXZw8xiRmgL9RFRfQUsYxruNE5nv7gWKHumP7uXHpyk+2wakEv6oR5W
iHAgpIQEM0ej9XvlrEsZ1q7GQO2TXQ2kW+T6VXS1QRj1QIOKfSTj2GkuB5VzUidX
4GkuvMnvlseHuznhyInlZADsRcG4HcP0BEjb0X3UaOlVBe/HKwwZDJQ/g/XtFHz7
fYdwfb1BiWsfv5nYi9UMszwt9ODVFNhHa6/DoE+ZJwiXprifsWzLSzcZDcbsNddC
xSjIeBZYu8uR06ODPHaQD4GHHapGPdSs6/tHZf6W/m57YGB1UZwCpwzOfGQmSqdk
V7/NtIFfEnxutERFmZwZPQ==
`protect END_PROTECTED
