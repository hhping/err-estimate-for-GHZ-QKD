`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzxIp3uNKdz4omsnzKVG0+NmAYKfVxijv7xM7B+m6gE/oYjBIDzv5gjxciDF2zzO
fWtoqr1N2+7IjdayuzMZBl+C04TM8tfm+T9BzKXE+YKsqcRTtiUuEzFUmeTtL3Id
iROdN+knaTpFE36J6n8T1KN33lfD777kx1Xe/kyr4yxunfGUtE6QhdmM6bSaKs/D
fl0D3e7YARbiIChGBLbM/2jcGt6awM44GmmBIMLo9d64UoPuwixicfOw5KKzQ9yf
9y5VRHZEZyrZO5bANEZw325VLnTXs8qkgA1sUCBpyzgMtEWgrICPuU9r7G4On0vj
tRee4SOx9d3Z+Tjc1l1aJg==
`protect END_PROTECTED
