`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/EuNsvAUXlQf4Q9ZgxxHAHHSkBUhl/fJE9W/rjGGNtMBDEDwrKx10yR0LHG0VHj
2u0Bh/KU91bs9CnEgQeR6vAvRHu/wz3W2IrZfumjIyol6+64KZbUEG9ur0/JmsB5
CRTs+hBYkJInUsO6OIk4hWsBHl0qnQ44WfX76LkU3geKV8X07VMEr7ppwrFqrT1v
EKLKOMgi75Ivmj/oZUf38NoK+rbrN6VDy8E2UD0KZvvLfdQ5pVVpV94Ljm3OSIDc
PR9QTw60PkmYl9LcTdaeoOvnHZso2vkxdr+GplMdfC5yg2avWTUQ1R3n6Q3zIC5E
70aev7niT5jRV9Wql4oA3ZZOpmBP/rKSNvT1kCgEZH/itolLh5ZskCVmBTUgdCV5
VswspRAaJGlUeWTV+nSgQ0t9xNlXo4ChBm1FsLYSsh2G1g8SiEPSQmmY/cMNdlZN
F8SS5yh/LWt0gJs+rWrd7huM5GgAVyzCM0FTuBERnrW/RlgwQBC+vx6dymifmV5x
uHl22t+pBA+m59LgpkGe5xnR2zC12JdgZw3SVdmCLk84v2tqzMOEXNJi3pOegLuo
3blZOlmNTnVxqpusFpTxIg7jPkhTXknooWo8eDHD6svXFR1+GMywJpWrtPMZE4qR
5vFKHtawlxZbOb8r86f7g0swyZvxA2Rv9g9qiaXTb1Eb90aOywDkvqWJsU0dy7z6
n79iSuLmUzTVdVT357CMzRxFbe8+XsQh0YoQYIJUoYdsmIqe6jesYFdY2b+gyE1E
VYNkrDLwfOSnwUtTz2uiMndTOHOlKnEtWxRIwt4XPjfICEdtsiieWd2/4DtWnUUV
CQgJpBcRmqwLqfcl13z5uqB8rGwVM400vllL+lWVGTcp3l5FPLi/kiOTFVu0Uj6N
cbBRHuHOQx5jMcFlJF0mEYwRzWPJebvqXd8HczxEP40a6al0xjYh7NRrLBm8eCs8
Oi07d77PmnsXsaYGaEDQhDejgSLyDHYWrfi1hwU1u5WQZYlBwKYSRVsJSiTnEJuk
ez9I09ou/Jlm9gkMJpiLhNk9FlrNJ/JHvYtNqJ8yAjpMdOSr7YdDPx8qaiahqPHI
7AbAaVz8HnDIT2+kUv14esaIxWbKmfS9G9TD0t+b389xF/pYklYdGqnrOfiKME3Y
81UA7OsVf3LQD4nmypX6B4agFTWR2qxy22sbdWTgda2yXzJBTbxiR1MRHkPlJMeA
zYlmq89bHwYjCbrkuCOcRw8wrpxUIYnYD0SiLs2JnIVVJZ8lyDSZaDRvTq8jDybn
HSxIBoUt/7R+wjzzy30WULdtIUAlCHupW7zFjx7plhXpMmVCGG10hvEfYwPOZrTB
`protect END_PROTECTED
