`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGQImCU4QhuerZ9tkw+w4cIjOxDaOH/z5Gpgj3beD1OOZ70yKwtTdXWqc7HgjpEg
oO8ZokTL/DZfvYJcJ2iozgpy16Gp8WaKryIUTF4lIMDlNgRcbmpd1UkPbVOOaH93
2r2DBbQcYHHOdfD2P9q3XogSlh6quzPxU4lnRHFHJm2rj79HA7534RBrJmdnbrwK
RlEciezyt4zvm2uUglGENZmKBPZ8PY8Bu4ZyfDm3hf8IKZkt0oz9nDR3FFJFOWZa
mWsAJLm/9GFJlOYsAwJlWTdXv6gwepC708fuYcgeSETdNG/Gf9MWJrifrIlV42pO
T4JKAzAXkm1MmoxBFETVXlCikQMB7xAcmc/POMr0iP1sATocJ8xis6XSs/rt/Pxm
`protect END_PROTECTED
