`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k396aYljpWKbeCxXsOD5oRqhgpvUiCNy7YFUev6I039pxVogY7dU0M9dMTOcujzJ
s23IsLHAKUwZ3Y1csAO1WXafTwHZ7hjhrLY6aPnABY4qv6W/omwqKiRw2LxgprGX
lUG7DzyYyddZmZYHBtuR3moXgxxiDRvlU6ZAC99w5BzkqiKJp9RKosx5KdBJ0oS7
FGq2hcqWy7rg4iYIxrf17cEnqK0BQbDL+r5XWmi1P7cQtkJZQWw2WAiee4aO82Ov
svi3L3xMSxkeJBG7MD38cVHdP9P5C7CRvBodq35HAw2PA7Pv8ReCDz8EblaT38o4
TxO2Y+Ip0hP6jOKGkL1uLz+823l+jV62KjOyMEVX5LA0nr46aUwrAzBxfjURsNhT
SWr2gaYpnwBgPUZP4UXGKzM88YfUoxLmciAcwGkpXeOh1ITZym3SDG2JgDSdCJ2d
AxIDF5iJBN5PN4anWN5uC1aUETC2tYupibqvlmVeq827V/N2AS+09IcsMGMjYPfE
EtGD9/1GxNub0iYiuie1ZqxzYsieF7GFjxQFrtyVhhJ1/ZYkc8AwIqC9dH8R8GFi
hiuwG3Lj69Q2Ab5Tb7OwVuxX9RuVt6WDKLFtUaa361DTWmb5esA+1PjLAvCj/KWm
cIZcCg1gGmsY0ittFQRdyjPkA3LREnAZDaHQ9yzylD56cwn82C/vBQfU018lfyK5
OIGQI8NYGohfLBArwe40NqzkdAZa0ovsAsDwJ17FJcKhF4TjFWpCL5V9WWgKeSlk
7u75xwM4AvJuY7GCgxz46eYZd8HNkjU1G0QUvQIl9DE1tAc+PCzG7PpjaBQ1AA/d
GG2qGeSmVC1K7hbDHAN00QG7zcE3iRuODKuBaobq1joAyNnAiumorMZ+yHoQCOID
xF+G58XO/+xtW3o+TdWKXUT00Qqrm+fjmK16y+/PLp0ZL+o4tlBfQQ6nXSsbAhIQ
274+6u9IIPRw4KP+PtzxZsqN58bfeCI6o+x4HjbiDlxor9ueOmQ4z/b4z/nk20jO
TVGzWraWKCthC08lw06aPLcpXoZgOoLdZzpmfPydVKeX652KmI1dVwVfbYWanTyJ
I9eTsNHqFQd2yIE/edx7ROAbhWKCK2PMiImsvzcYonJlE+R8LiKikZ9w0G3kc8mI
Kuhgz8/ca4lF0L1Swy4K+inAIh6Lx/QgGs0IPD14L5K5vhGvAEAXw2yNFQRCtHh9
DqK4Gz6zx7+BpFtLdGgNIXLnfyy7S6kXFpd/MRuwV5BOhbaCfFkKMVj4ShAvmk92
Gx8pqrzlZz2ff2/IEV8c+w==
`protect END_PROTECTED
