`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4kAwv62y07Gx+V3IKx+qaEy5HoWuRgx0jANLB1/sybFAvHknW4iy6V4P8AjmrtSK
wN+1rKTIMt9RDG8HY0WUgYlgWr/qoHw8X6n/4MeW8k5ihqSVNctjvTC/pCz9/VqX
+X4cMbixjJGE0kurwmWgA3EZtopGFXZnafp//WW4UL+gwroM8YW2zpkbsEkq1bAj
S0xZdKtYRbLASM6meqQA+8C6fb254SeVSKIB+b0e0x7ZhrJ86lIGt0+hwpsLy2+u
m3Yo2EOFqRhHJwPvkKr/dbjCEBTUU9qC5y3sy7MdRvcZykpsiFscIzx0ACUIITXx
eTh1b5m1HyIxOsVbMqlYq++4tQPJtvP8aE7k0dIpNykMGxVBs9w4981MYdCmzEZ2
hC+CEO3z2qkGMwvHsCuinWAAbGYEXHPSgTPiuGLdZb310JPviSPEPF6Cl2byn01h
7GyRp1/ZFRROy1UCtklbl4o68WBCWHGFNYTdj4xzQvtDVVmI2vLg8eE3tUxKbtq0
vlheXlJ4jCkJ5af6BU6lOn4rlFhhKp67bhJ1zk0q3BuAMQ73VPg/qARaYk+s/kkQ
7A++uZh4+kT2Y5IMsuchj9v4QG9V3Nyu82Hb+6qpmwWF/KUZlEaGsIfuIDEKFT+Q
jyqfPAyjpbXc/NfYRPtT3QQF6W1m1bts7jUaUCa90fWWqMU3z9J3R7D9T6uQMp93
r1iy5XQp5mc+DkkgOatozaBqWf0htxO9qaL5VSSpRHH/th2n4HQnwg7BJb0b8oPA
2ugbcF7a+wI/vojdlXU9KkiqNVPTcih7qwcuU20dR3S/puCksYAlT0GAyKoSDlye
jt+MMlWTYUt1LpD0KIkxHN+mkuYbL0Itn/ZcD7LTulvGMXmVCU/UvgvsIPxUG78I
9fDDv83jT75fsNCF7Q5r6CfySX7PfvSJOmxW23C0PUp8e2wwiaEsTCcznf/JnYeY
mY2dzzucw1z6BXFfrCQZQfEP5XOWzsZaQ7dwWxSw2MX/4WTkkQ+Qe3Yv3ZTKL0gc
i98VlT+oQe+DZGcBXzqSmr6o0rT+b4J2C5qDw+L2mGcve3v2QDieXk/b3xV7y8n6
2U4RtCJRSkBPJW9mnoiEBQ9YER8uQd/flNRpAPty/ipGplavhJdxSLk8IwGOimh6
FzKfl6k3xC2VqrjLnU5hmJjQLAHXpuYy4/r3HIdw08LAlCehvJdYMjrtceHHKqt0
mG2IGjFvJdarh+xv3QM4PnaHs8L224geQmJ07s52CVbULOpjREjpEpYNO5kndIv/
`protect END_PROTECTED
