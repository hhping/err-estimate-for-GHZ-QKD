`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ERAN1pOBUHmuWA1kVbNG1LQNstC7q/0lUaCiJhLxATg52BGWlUFIvD6ijE+NIdhn
MDXM4IQBW5t0Wr5X/JePVSqg+DqDE3r25eS4zfLCKQk3oUcN00Wq7/QES5uCnDhg
9bm5xamTfPE2CatXYvYM0V8BoLv8+FFH4gOZZruP7mwToEh5clsE7e6ojIJfbICM
hEyuluKqQ/00nZnkDWT/hal8GZbjLrJBOCC1biAX431GAean8uXfAZvVonSZBxSY
45c5SdE/crmjUtfEfabyLhMPN5kWJljil55iroms9mNrPFpNSqvIAZG44MxbF0ic
aLB0avpbaH/TyRpn7j9qVj+91weOvL7CFxmFZunUsTs9iiA2OVSppIvo6yMtUk9c
eHQXthbGy8b1VnDsXVqtb3yuFowbSIEMDfJhrV2fO4g6TOvEyW2HC4hy24MQRu5b
BhqyRvLEeTEkQdW0k9M98oOVLuvo9RnkEhtXfnSK40ZsNHhme7yUp/oFvbhuOgFt
kF+o5IuT40TEIn38skGe5nL/ROY+MrV3DpN6udkIOt4Gy9B3zmcH+4Jbfo6h91XM
2YL0sd8ZROSQPvjmnVTA3KFP3XxQEJQZfaqj6XlY611KtddPDCmaOAAV8tPlD1yP
+/Kd5z3HpT9oLzYLSvdUgJwBwz74MOQTOyMEtfpe2OtomEScENkdh6a+N9X1+726
cJQLXB28hRjCK8plutb4d+aMKZI0h8KejiFCe3yYgX6FhmQNJ0Fqe0KYfS6rqyul
rRCh0WzPspz7V0pSrPjsPyafvArBePP8MITngvFezi/+7/zb1ARrWmWPAPhA5kxn
V71ndsNN9RSPpC0KwmpvKrIYgXY7uoT6MXN3fSBDdyu+lCGL6r6nh6Bf2MWOydue
cgLvvUL33xGvyEv7EXROOxb9UqwdOnFq5uErVA6EeFsKtjoPB1mhh2iFf+Twq0uk
S/YFm8L8jpjVd91Jryr0wlECd3AeXNTB0fnzeJbL+TLWe+BP9t4CPwCur++QzUVx
S2MertNrctE+F5j4QWqD+ZjTvi1YtGHHdg6iGASEBV4x4M49dt/FfJF5fn/Llo9J
hRbm9V0J0/aMFzCCSTHSmmX68JmRJYqlumD4t3ti+dNZyrlEAGg4e1hY76naq4O9
gYnNskszHlsCW7JUqoIKDw==
`protect END_PROTECTED
