`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0I7W6Ibt67HlGGW5zfjV1AncgsOw3GWlCdGV5WNq6fwxUarUydpRsFzeYog4HNw
/mRq75xWVUChVBhLOOQ/vpjgNCv/wm9UWzPfquhh48Mp8BnhJx80F4jvENiIN8OH
HGvENCLiRaUWMweWTWI08292Mn1dduTGdChM94JNOWS+h2bQyJmOVzwTdM+Y20JU
MeKODLI0gY3RoS/v6eIYCXBhxIrpQqF5LMJDyGRLPx7xqpSOGSSQ62QwBRass1HV
0pqcNuW+dWs5HIzbKZtLYXDA2V7ssqaUM1S7Ze1GcpNHus4xslDWyQw+BttnzHnT
Ja6wszCz1N7xL+vrOVWz9eDPMrCF4fJQ7Js4+CpOoa+hLCsENMWUFQXZQ4M0fLMn
U5Q1YVKUKa3TPJR7f2Air+ug6zUOsgbIculDDGf4EGnMk9olMZDoN5c7DMjpg8xW
UE5bplUdvLxOoRKA5yS1SdJdBzYBU8YubtqUhyjE06/oZLX/DOTBAlmt5q7Gfs5f
JogwyVareN+vLK2AbVCDTOGiA9PHwKGudKHU9qj8/QTrxsVm7kUmoDLTROleG3Ir
7cvfc6Fp96cEsd3faZe9KaX2rOXFrJOQkHXmEc4n3VUM4Pa8IPmC721/b75ftkkQ
uFJIxhsoJP9FaQuMN37a0sYR+N6HjYy+twFAmleywcR7jTgi14VgJwkRKYOWrUS6
guyAcZSWcwq0ZjOl2gI0fY3nZPMTSVeG5EI8VqG6GYoIrBS/4umstkRdVI6tlNDK
VrCEfu5jeQtH0JzqQnabO+YMPU4X1fXygfSswQWHn0ESinGXoyyP2itKReMoi5ju
KhiQRyJNwmcqTeIaGuQckYf69nmE5WDYAEx4Wo8svebGM0QjqUxG3p96c2htxGzV
s83GAosXqwjOXOvTm24xibzaksd5rG9dmn7SxsvH13AVzEoAlMkDZw9mGM1k9iGo
w21fTQlm9zMze00PZtxXD/PTUZP8EWigHmeJd8fHvzIzh77n46mm/qp9I6JOVjcB
g6iHT5pYnjqGeLt3pjc8ByEMDarbwv53mxjjuVcpukZ6czT2MQErCGpiO5+beYSL
uZ921aav6E7eMQzY3uAtNV58/O/5+Y7MYBy7BqfYv88kbX/NqH5437wRwbLRgYac
77UZepPvIxPnwLIV9GGoMP2RQL96iAOuBzs2ri+vXf28wkH5mBSNXD+fPNwilQ+m
4auWNUYyd2h7uS1LQQ1FVqUByqzW5WTdpZRs/PHptmcWE5IOULkE2mTOZZxwCU9V
FhapGzNms5WjSJGYwEvuI5MbbXqsryg5GabxgmXWU3780J9LQ6yPJWG7r7HcxH8j
pRFICjTKXc+ZFNW+UU83zZWjaMpy1AfGoJSPPEkDQBTfIdcD0Y5XR9kQgShGcuGs
dpXc1BfdHyanOHCVwy9XlMSV89/tE0kbq7PkN/UppOXFFiSE70Y2sZ///Uroyc+I
YzYXP1qpb/0vOHkR/BClIBYpGiNowKdlIF9D11iv55+zLlck/fp44boFjEMtVMAx
NMtp12q7CHD1WdTotZt93vofUyeVewbW71qsEYXqK8KvuCDGIkCC1OF1oo/j28NF
LCsTj0QntfWqfwX2lKpwRJWvXfEFUkOJZKWbVY5E+g2gI/R003u0G8vyS/gA019D
axA7QcPedUVPz/ZLHUzxvxz1AEMT954bfpulTb1pZ2xHKC+vOV0Aa0ZXWmrATtsA
KmrrIxLt7/3nT0SvcONool0XRkt28VczS/MN/0gim/Ajcv8Wl/snj478n4nBt4fe
6znEuLAjNz8DN0u3c84dag4Ytwe9QbhIdrU6m2ou86DOOcPQy6mR3kRALZjO0u56
9s/9q60jP+VU5cT2L5eWZaVo+DrWGNAbCbUZSb67TGwV8h5lAj9H7/5HlFutj3Fb
yq2TtVIpUAQm9LWcxNFOgu1Fk0omv+3rOmkv9vE4D6YbGHYISnxkM2NmYZdfU27+
`protect END_PROTECTED
