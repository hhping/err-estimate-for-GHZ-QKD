`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKCqZTTP6FZAbZbEwIAp3+vo0IgQgFNnvlHpmnTC/h0Idko8bT/NQLIEIuWkiYbM
nCqu5xpaV5rV6clKw8RxQdhGp0pic/TipngyjnKlj5ToQ0GoBQM7+BQiHYMWDKU3
WRzCXj479h+dsO6M+pT1w4KAZsHpB23f9ws2oCgUWBoLB+Ts2Og3MOTmAtBbEmMv
E3FUwgB3pTZBOOxK0aqvYgYvjT2rZ6Y8oYSksIAf6XNHK6m8HCzoe6Cr1Do78Yc9
WyM3pJEjFh7MFFxZcGeM1j5iunJpZjbmtKnI+lkADrQ0MbMc9hLsCrkFmBUHLUaj
qiM5x6Lc+LrHL845d396c4Cs3ukmNA/XEk5IU65crUgrd3W6o1Ah3b7g3JUtP+lX
2B0ydQq+8N1PhLHexU0cvqXQbcX67uxAHpxVQNxaIR54ZUF17MJHvb1Dyf5CouME
BfnARMzLNolOVONbZNo8eqOCS2fBr3Pxr9ymdnwi25I7qmDiRRrE6o2uUcfqAJa3
/TFJDMDlmRimR2zY1t/4S0d27dZ+Fn8jtbtEwvRrP6vaKatWExI81bu1z9dPlrnX
o5Kc3d8ZYO5gE8H2JiGqSXT+UdpZdygH2xh/6Q2dQsSkT2NxTQp88P1L5b3J8WH7
`protect END_PROTECTED
