`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8XpOfwi73rrvoaN3UDnn2BB1XkkLKxwUsqrabFI9Rqo5tWmOONNSX1lz39J04Hq
R38vw6IaKamq8iecuhmAPGOiZoh/ENWAEQto1ODSkmelz9eHuVuv7GEqcF87M296
4YVw/lQTGqISCnhhkn9/nKRYYfe/PrsTlEqIbMh8WKu5uDXELfXrlkFFRqU93/yz
FLvBrWZUFxzohu5qR14cFNAPZRwRZKYpTWk2H+VdJV9COhSjDzQ7vADEjtG1hy0D
wousgbLMpYe0/BtJCh2IkHHcNtX//JOMsLDkh6J+oHpSe52CY/f8FZnOEtI0knzJ
OPgdwAWPQd+6l2Bfn5c4Iq+veaEPFfSjzK+NKS320g+vct8+udZDQBkIV0r2PMsG
t3/mzvKMec+R8rayIEzVuzQHRioN7NgPN3w6iRf+1kbphg8USwj7veOemqb9gHyu
zXbPQNdNbYQ3VPGzoBqDWRe0XX1+2rzxOtErt0E+YC+ZvKPmcqE4MsEtsgDDn+d0
8T91oJMdQHk+Mr7KfUaE+bLZFSAEA5sVWPUeS4kYUP1fx499G6E/JKp6+JVhf1NN
BIDJYLU00zEJVPOXAVlvWyv+2glr8bdYPmJ9Tq3Lai7FeAJc64CFQQL3K2EnlB0+
jDFlv0GjjxLl2L+jesmULQ/lsMyMGnQs/TfzbrOQjEqRpDCIcMZ6dOU6+Lng+y5K
11O5HR92CnV7RytSZ4kNJZuSW7678LmW1H3qS5nfBCzD+rnGbDSOMKtPJR/e0nwO
rYyEfhmcATPejpxJjKJNTMLfx9D1ICoAH1dNRyRi+NBAkVP8YRtphNYOnZfdfiMM
ekRMixk4r89btdzV0lwpvU4uXCnqz1G2TvP8L6ySVqvroSeQXc1Uhn6Rk8H4YK8Q
sr4cjz6KVS0owyr8se/p+oyCNiJvhXNnxpcw6zjxQUQ=
`protect END_PROTECTED
