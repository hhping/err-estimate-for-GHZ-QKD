`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XYk29rrWHga2fLo/dP2DJ9HqHq7gnOz90v+Jp3YIkeLxKY1rgBfcXY1xyxDU7F7e
XRqF86sEP8R2UBArbexIuy0jKE9RlSaDaV25j0OoZvqUHTwzc925W3I29wdmtw9P
neNvyH5O/QUu6oq71nccSok2KRWZjirGHR+oUJVZ9xgZmv53yHM9UT9alT0kOi9i
A4webTsdUP+N0XKErb980VgApGnwSkKnFafH082UrsbsZ93WETxaR5xbaIqVPpZu
3f6IRCdxtNRtuXye3gYAH7kh66Idt0UvPqmWd1FjvgdMPSDtWqGYu6VddsxWMSWb
HuY68neHJV/pyHODVnFd2Ucgi+IGFqkRGAKz9oMmWMrFZeeCB6udP/nGJg4pN8aB
QXLkQrCWZKCbg/STa/xO0h59qWLFhTM5VNNn0vGjeHWdnvlELUk8O3KvxmycfUL2
waCt8ZqipaT6mSFI1fa89Vz5YanIAMfDhX6ugd1gdSbZJvYIT613gsr+HaM9Nxpd
fuPz5j/99SqNHD+nJzUtwfKJcUu/cP6QKsep5H9bN0UbmMnW+J6LvydKpu9/8jTn
RDGTY+RjtfTosTJVdovaVwJmmmkG0ifTE2oaV1DSET+vbYZEsMINqHGESfTVTHdX
CrAY/PM/qRCL0OiuMoKgeX5F/jwSq8iDZmc+K8UaDbBE6Upzt45JCS3B3hSKbdPd
yTxRXhaup+xFIfAo8qpHd/8ziRE5/Lsic8QxvMDl/Z0lbSElSppy6fxmceSEArbC
8655E90sNoyU90+nTLZv7IYlm8BDr253wrZlJtvg6WkURaZCK7elt/bwVqJ/Hd7m
ByHOGeWxMpnagxx3ZHwejwUp6IQ5KrAUJLYWchfonmfVPiCOx3mB6v9AXU03QMAY
MXhw/LHK//jwWfW8VdL51DWe/Uetw/dBpwabXVF5OCXAG/uMvBUjE42bUoqJXGob
HI26Z4wNtbJNxg8wcZ/Hrs2/Uu2txbJM8hTOHsp37cEapjbeMvFcFHfHWFCNz/iW
XZYOW9h+6kXg3b0fbSE443Sj1JRjUCx8RaHSoAG3enjxu6b9kx5oW3b9irgrvq2I
+mKd3FbHVoMV5iYdXZsVwL8e8xKg4tOi54MHJ0ArGFS1WHUvr3zudoV8dD2tdAj9
RcwrzdbwtF/1V3D5AxjbvhjXO0sO0G1id32T35WtZfmg93lPZW7Ou0e9bS3fOfez
zMP+ZKLjPRUyidU7sm3NnLAPidEdq/0h661COfTpbtvz/VguXs8yWyaRhFVLN1gX
n9nEnjJRf44zxymHG1IDnCVJEak9YTZhJ2b6w861/kAY8qRwmLFtXgUcVb1BI7Rl
BqBj+EHRTMUAFWlU/ht0PCxoflUct22ZKBWPJpfzV/DwV4zuygTb35Wj2xIYL01c
vr9jZFiBcww4s69rnKWOpUQaXOuWtci7EBwLx1T61h1H/Zc26flpGfWI07VlLtqG
cEEcWJowQjhCtRcS8irnvxBknvnLY92vOsTZg2NaZoLIlM1o4HJ/3SFxp8sSn/Ky
J85/RVhRey8IUHCftFTYZabML4H+ZAyz1egxE0vjXy1VRImHLdy83xIQnOQSVwHz
MB3FElbtN1W2RykevYRWzYjm/vmO5XhfEakHrYu71Q4R7bvCEsofnzbPJgsiejLL
2eoWaETmFoos0cae8HjezQ3Ltz8zPn7fx1nRYu2NDjg8dllNcr/CPIj1Y6Ss61Bl
bFp1vcIrZXdnvzZgDRAZ6hfcEkl1dUV7+fJOLJbjz4wnJ8pj5pd1IcPo09bClAGY
tDq7cM3Jz8SEfj2V78o8F31kccwfCCRAk3mSz2gSKrsHIP+tGnfv+iQVU6U2BJfw
o3yrM2eBBBhhGtcxylvQyyWUodrxDn2ZlhUh/jO2kWs9fSpDOaLWlGJmdpoEis2N
h+SNCNCiMNckDO8zopG/3bPjnGl2n7pgbZ4RvF3mSQgDfRXgdYsVzmy4id6LNx1L
rJmlLyTWey6fZ7u8hwhRSs53mcT2n5xMjS4XRLJJaCYmMKwMn3Wfe9ztInVGnmwW
`protect END_PROTECTED
