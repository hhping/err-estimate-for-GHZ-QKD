`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wO3DUwN7SFfTsacFZk4aja3xCUbt0wrcTKVa6ZMcYeFw188a2WEamRu643Gbsela
qIxMB1qrYO7KJw7VjDjfHxwPnzfofqvdGrrqkRKXbDk+HoRLjg9V04KmDINNEFPJ
QpWSyTKps9d1O0KHmicF1MMFRLmeZS86PM4rw8QSjPsKg4m5Lo+WsuSjTyRknexM
cHTV6+5CS5nmYA6AAz1wFiwNFyMnQlNLcuvLcwtuxx6N49hS0VVePvoFkISqqYl9
46JwVUyCU1jeBbEfk1LU4kBibxp/Up3vJ21wgeeuJv61tUr8MqhAB0PJFNLvLPEs
vVlXuQ5BfRgRG1M97+HmpzoL+C+A8Lx52GsPxyiJwqfm/hxDBWKBKMtPI4cDTVo1
bSHLDQ3S+v802u5hM/b89w==
`protect END_PROTECTED
