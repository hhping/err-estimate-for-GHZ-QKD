`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFpoySOUSN7d9hPNQt+8kfTcuxUGB1uocc/0XKR5FRV+pvQgdGfHD7vAYAFWglbx
vx0CtqeOeXI1qqLKhqHuD3pee+DaqqanqzsFTscW4v3QRuAZmZlwKy0eNocjgs5I
QVNIfWON3fqTH3n8dJOwCFGI1uOEP4YiTcvPD1oaCTWztr5fGvWjyCaR9rYFmV3k
St1KyM7Jamlxw8Rdhsn1rHvBZ9WeiuQfUK4S7AfdQZ52E4SlodFr0jm7mnaC+nu9
9WzL1B4w6TYpjT1FpTP9imkhjjch/uGOuQVejUvakKfQ52zY2JiaBVtCuK2CTgww
VwQmLf6OdDJJz1MSpIC4rP579Pp6UFrh18yVFn3Si1+AyCHTzUvMNVC/Ywtg7BIS
6F/5nMt0MHvgxGeOHUEG8tv3j+qLb2QfbpheAfY+KGNbH65xaKkPT3y909tfFG1Y
TA34QcfEAU5+QdW3uosBSERRdIwsgIRdZvFZokAMGVAuQYk8MT+Ej6+mTvcY9IOC
`protect END_PROTECTED
