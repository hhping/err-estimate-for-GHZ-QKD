`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xi+YVjTHV9vgXMXH52qR3WDknlOhtZHUA/wyCYWfMV8a7Z2GT1ekJgromxfwCnzd
biwr0uk4caGxXbz+k83Im4YQhcf3d81dV9izpW4BvVT34dnFa8T64wyqEFoDb6Fw
BnkRIToT7UGZrF4tZ9QAx4ux3GIIWq5R1Z1MlKJFVuB/2TGrGU0C9nHq+WZfJbtK
10Hd1vZbfZSy+FmK1lbAlcv6sFsW4MVIKOrdJGG99jj2OrtIvLCRrtNt2jEzyAvN
RI06aPdQ0Kc9NyzOD1OD7mejvpRP6z9JdwXXmkBPHajH+haqmNkDXs0V7Qe+Xw+X
E/D1voCJAIHQngUfnDmHkI9/MElYh3d64HZrjHZHkqCfMK27fcVq++s13ol5ZW8b
c52LC1bXVbRdZPE6SQLtAQIMXBsIh6X6D4vHiIPF161p3/xBC27KYkyT5VEsBh1o
VF6vpMEDk5YZo5u7GRxkXPnat78DC2OABAIQaqwn7iXUFKE8lk14Ovg1eXBBeEmq
fZT+XtNhb2St/dhPZ6FInZN23SWCXDonj93DL3Y+dyKGKHzuV5+18mi0Xb5WbIRa
xST7pNfCby1GQdY9/kwytQcw++jueGyamU39OuQ8su8XyLCtejf9FYXh2gqNuQk+
EFZ7XDjmrYbr5gS1ph76coUPuFKBUQjk8AB9Nm/Ox4DLqvXSIrXNwukumiGqZoEN
Nq9yjIQB9fgCQeQTqFkDE+CaRKW2pp4bqUnkQW5iiF4H//33ZhGjy+PCZjpCrehK
AALHCIA/YEfCZeVwCic3eB86HoBSfzkt6RFuuldLl7ydbRG1pgex5yHzfsT7IfTu
cS8zDygY55kkXULKNMGe2sOVb3zfZrVNsWX0oXdDOFhPhadYXVh8Ls4b+T7dEmcR
r30q7aIkORhRiq4V6+tb8tgH4ZV79jqEQa9AG/UPfap9BL/PZRYRuweWk8BWnUfS
x5x0G0mGgORQQCG87tGQKItuhiouOFdVjgDqzOoa8AC2Ke+KR6uAcFYgtOr9zYsC
EPnEhoStxKrA7+jGY5cqkde4uPM8Zu0X6G+8uM4kD92l8OxJXKEUBjvhmxkvraBF
PmhCVmYDqXGyO8B8m0CYw5DV4pxymvEazMLtdXL51B/3nlOmRs1umYHbW8Uxo6pY
tOia30zgOAb4F0TT+4HCwHvgy3jdPOEtbJBgd7X6YLmUAxjj8wNJ2JdqTAE5JNPE
gAJQjDywJsNuLQlFJ45vdaJiQ+upgHLfz+ByUUTWc60kZg3T5TqzbF6YFhOyhdRh
TuOnoop72zDagwhgj8Wtf+c26t0EEz/Lt74kmafRqxq1PMTsZIRwPmnvnDL+AoFJ
goQXSwzY8wHd+9TMJEWUxQ==
`protect END_PROTECTED
