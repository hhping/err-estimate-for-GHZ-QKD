`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evUoCMD7iyKU3MfLt+VpDxXOERTMgZbwWr+r3HvENDkzqPIOGGokxKTXBkym3Gr2
S542XD9I+CUjzFQs2L9fL+EAm1VCrsfEvZcyQYhQzCPMXsUwe2oFs0g7d6gmCezG
3ERcTzvaX/rjZfVmkanR9+LzHPyxe7LnKn9yVr3yNc7NBfQGcLqS4NsqvWoHBiKn
LJcpohE3N6+BR5/8/ypCjqf1hTf8eGnGuJFWRBcKuM4s2jlbSzDK6UF+1bIiHshV
/gE0AIfPqMEtwk1uCt7p2xIk/+2hXPKBdiiXq/vraiUp15CIALsjaRrwbMAWjb55
j5afCS/fSlE4u9vatucbY4QquspuxYKF3xrrVwz88wWcFTuBRBxD7KOQBM62v7xE
rGhBiJo9GL0NQT9p8fIEm11Uj+fa+CHmoS2xUKNJOB3opmV+PcXQdil4GcmQJvW2
ncP80JZOj5hg7aeLeZb8VkY9E50WbUajoGXOmc/zeaenoEX4I0DT5np5kT33ANFg
wIP2w5LUxziqV4a2c7Db6QsK6i7c+0nHVJAEwet8evbRiWsXvVPJhaIl3g29Gid+
OtSOJGQrPZX4wxS8fp47t53uldedVzwMJnj8B2aB63a990PtGNZ7iUUu2Zcs+SyB
d4SK62Lx30qPpJz+uiqvYsq0ftfFBZEoDxukLjam3FpMpbd4gtvNKIOge9zn8GWF
9yN7fbDIJ/rg676bSk3ugnXqwiLqhcV88eqLJKILS2wpRsqtfRZqPyogDClOorEd
`protect END_PROTECTED
