`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMR79wSp5C/f4p+fvu11JMIG+sDWA1OlJImTKOjKlaxrAKV3CMM3Z5SQE0kMBST6
6jugvqpjo2H7u8eKwnF0K6sZ4gCuk2stLFLv6piHqaP0eqcuPCJBLkYBqjKcYVNb
vr6OQhm26OUzOIzVAq512Oy3XcJhYRzQuEVljLzoiWpnXSNkA+SFttUUHhC+oOYT
tQl4h649/4MRd8dLcsLjJha8nBFxXvM1RbjHIraPUoWVxvwjdG50vlBRIT8m52VI
2d55CVlDc7LmpETvcy7Wg4ecuGp0ROLR7I3tAjJ3A2tI7N0eQffwrBU7rUAsdE3n
TealSGePFNj71KcmxJ3ZjTKu4XMqhofLZeEeqzxcxcKyV1lDsugaz802GjEqZZwo
OeMPy9Vt8U658LnDTd4LL5/Ak1ESbmOQz9iF4PfwcNb9YApI6B4550bp2M4kWVTi
IxOzhcYMSC90SGA3ilfCJ2D8nZreIPzaXfg/FcDUTzrfmhM2xrEmVJ2x1W//MMaI
n/nwUYpf/URAJCFrtWgz69KUgbx3ct9rifvJN8uYaLFqcU7hxtW2r7AyZ6HUUsqQ
ErQoxv9Q/DhgP0djchpU/ImgJQCQVi4SmgHFBkNIvPhGwrg82fs/7ZI4QDS5jndb
ZQMZi8Eb2M51cbG1jTtGQfbhkQFURnkICWdrqlQQvb9A4uekPQN06UDN8Qo2RImr
N2PPXwn0lhw9gVIn1mc0iQhaALCPzUdlAfGZ1aQZwyMh4s4VyEwS07giLDvCOTrE
PhZNhH9V3zbDH8+VqrTtjzgjMDVuMS2x3KsA2AZfpvR4MtRxNKIT7Cvne7OCsuvf
6xjw4cntgLdz3REv46JcSoeuiqfCSZnIkGVlmYq2b6fq5oH422kfsJ74+VUHD6gS
eJfUWJ5VhrgWxHwsCzb/42/a7ih7CmXsc1XrLScm537PC6vwcrSOiA1i3WGkgagZ
MeA2z1qFeRh8lOS6WP/lY0Z6DENEU2o6N3vqQ+mcCtaqgSDR/pvHCbUWWWEi5iPd
2U+RmUlT8M3oOMsiGYgZD0kl7PXBAWD1jMda9ME8gfpBaKsDMxoopPJmBHHqjIp+
OUKygivA1HgRdxU3PAcilhjQeSFdkEoWxMcHzAR03I6TbflJm3aOHmHXTfVzue2P
cli7tTItu/77vw7CB2HvXwgodx+To48r8sFEIhCblrSItQXWXWvlC9/uewYLJsst
PsXllmDLiweTWSb9/AKlXxJ/bku4cs5pRgAVraBaHgF/JgaY5z1JUFon9XhPhPVP
yQkNYAm8f5wfDSIB0QnnL3Pqsyrk7qy266z9VcZr1J74XK/WhRZ238GxfXGIVjfM
3mWGs+XbmadDlAkn2nRO2m4voNz5inOjdzKknZAC8tnT3FkeEXA6oJ1WltcdvVIU
t1HDIjvp1ZOIW6D13AN/z1Kxn28H+atK9k74Tsq5tULpoYKQsUr3CZv8NvWkhvv+
ITeJ0hR+1V2fgRFl0CMf4Q==
`protect END_PROTECTED
