`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G28WOmaGt40yTqNZzFdgRagSjxCo8H7axHc6rmkeCNSnbkx/3yN3dEZD+TivoDKV
GloXXpt7TKy0b+d1L3m9/ZRK882yJtdQtD5ev7bl4EMGC/zMUi1WMnrr4SS2aBV6
gL5zwwkvASZiHiiooPBaxYJndrwrW/3XUELHJ8C8q8DfuDbXZ37a4mMu9EDryGBe
I445xajwpPt3TctIpHtr79PajakLFHJ3qlUPxC3WnZkBHbP1awQaRvZMW//1bkR2
9OJxcgbI/wkAnBLvb89hfp6e7ISt6gPAvF/QR40Zo1g+uFv1IhUWIHZGCI2zWj3n
8+K+/nROBKHUnge+yEtr4cBeAz1JDGuFZAIVDZCjj0bIMbLLnykkIX522eQR+JYl
VbhXjJ/+BEeGN0R/VyaRMijA/I/JG3ycOD4rSTdHJ2Et4gSlv6rPQGRNorGQcEVz
4XGXlvGljNm7PJ1k+IluDJTQcnBhRF8PQcwMZmVxEeEVGOISK94zLyUS5NB9Wh6F
/s8PVRWjbc2YGZLP6+dzD2CGT015NG+kl0OdKU3yoO98q3evOGk95wm08BgRSwmL
tZDaSDLNcizOmapAFQZHXNqpny/JB5vuGjKYXLC21qMfSPwewOdBw3q9zvu2jVCM
xk8amEFEqlUuLI9LR0ZwbMpLuiXkPb5wRhfudedS0UahoaOu9EaMlh8DUimo8fFP
jmZ29MTDmNjeeLofdlP2qiWUeqzHMYY+XthoPK4S1L3C6tyuJBBja6oPxpox1i2p
4d6Vtcu7eC4SYhpMKIIWu8u6+QkFVtb6BCho+S+RlNrl19kLv/wiToItXZpZ6yxA
AzUYbnQ+7q6FQ4zAJH75IMeIBiaZVuQNp2gAfVCKol2MfuwhSUcJN665u7dr831a
U4PNNfu0dZdy1uPLJz3q01rapuoFA2ZRxd2/KJWdN96yxg1k738nosgFg+wE7Riv
6UkmXuSiAmFuzwQSCzVQDAM8eGRh0ZxXGW+t3lOAqI0CoiWkY3YElFnIWDXWhhU4
niSyM4AdI9N4Bcm727pGUDNF8Oh6Kc6oebfAkbmBQNaXtVuzIpT1WYgDYH+ia6J+
eKhqfp+q6fHa+BGHfEjFpA8EKlw+ZqYyXUhH0t0FmJgcVX/pyUKcbZKLNIfU3MHx
gWwBYntnHUSo7tfXJMHdTn5T3cgmS5K0nzV7BtUeZQp8usBgtue/2be+iPMhlOyF
JX5kXVBQx2z6vB+SMiINrn/1BPxbQjHxsL568N+RA+7XphkjF3xTbyhJHq2bH9MX
FvlOyXGHAJV+vC4g49lxtqDJQtY4H+GkA466duOdH8uNTim5bSEse/Hl6llrQttj
JqhkI98LP4e453dEDuqgaz8XziU00BeRf5RLgK0R85SHRW1O66+7oY98r8Jbr7On
dzoz0o0qiGnGXfrr7EgwOsdPnvMsG8wzZHLWmGAlUljYH28cbuExF0KxTn0wSUsA
Ya3BhnpwLPb6f5xdFbcC3NaOV4nElRTl/i+DVV8LIllP2hA3Lnv9WOvjDCeTQnj2
Ej4Tsg9n6Ax+UJSvbJh7mdTGe1hzDRB3NMKvb+2pudwal6n+g5G3DZ/oMgFq97Ze
zaPPt4OyMqoJuyh8GqaW+ZGT1hy/pU4FCv0EdpIo/01gMDKbeR3Yumzc9D9fiUEf
Lsb6OEGdMYvqG0aiQoSPuOT7zRC7nxCVtl2mP6wO6h0xkwdowYSQ4j3RUfHArOtX
l+Pz7lfPLVDq5niDuIWotM4YYEqjgWuLp4KKIqRayTfOoJ2ZpupQ2+1dOYpsG+Pb
UjeZp3lnUVi4zyJwFNXRfqp3+3031Xrl46/gD1+Lx2KaO3wH8zNsjoIDXqM9+u3E
Wbr5OW7tbfPtgwy9svIhAmQpmEmfxdht4v/haS+g4vC3f3LSheqnnwOUkf8Ja0dj
l1Il7ajM6g9WkS2acpYwilNdpwKJ3KvmmyxWl+6pUiHFHgSSlpxSEZoMknTH9Dr5
+VZpvC5Q219cfpQdRvJsZEEcHKN8JAYFianaaULJ36obX3F2Uy0g/T+Lkd8Xwqg3
yT/sUf7galoScT8kZJBw8E1jyfR+/I2QIjy2LsTEQeRNICQ3JnForK0XqeH1dpwr
1cGeKMBklK0MK/AppAT7l7qWbFcwK2n4DW9IWaUzHbblGkO9DeVzyR9jFAJg2yYT
uWmk3+JVKMHlK1kLvfHm1Sg6OLKN6pBZ8ruuFHwShm8s7lq3vz0e8syoZX5pnqyS
gVEaY038KjMSbSjljc+agXrabzYMXbjHHKab3ECq0TzdsF7Fp8w5wvVkrDMmh83f
xYOj4VgpjwOeLf4REZdPaCcmtIXbRhIkBOxxisSxvHEGc3yFrnUlDaA5GJ378kUm
xHN4bmLTGvj7/Rdrum5rCLpBvcbVBHZIDxNo5Jx0+24GRhWv0KOJ6QqFw+uhdyJ4
AyEc/S81Hx2IYMGLh3UlcccfiAiUju4Y9S5696sT3xfnsMAJOi/g3oOGhPyJ2TXH
bQzaRdyGFQexmMY+imt88UHC/KJ9htQMcJkPc+5R99VeGPqhVDmcAW3V/GG+NQrK
taHOPeKbetqWndbBBUjSA/No4JjnYfRGjEdjBM0mX1cw7pUdxgGWDigoLbo6eDRI
vejcjKICb3VxvIbLxd78TcF5npeJ/bjf59bJFPYApr2F83aR037rFeJnY7cGJebB
GIEQDFRLehe+38KxaEJt+BN1VxO0dNLkxeRg//OF/LphZDAdk/7Ti/2e6jCXXJXk
ePqeHxjMOyjdOQi3fMjXQaszyPL+B49s7l5EakU8XKArSl8ynii6T0pgdgJDV9CY
PdgUkSc4yrRsVBmrxg3Yc6f3S1Aimkawdq+NPRkRPRsSbMWLSXzC5RbuvkxPzE1U
Bpa8B4QoAD+RPdTsIWWdTQ==
`protect END_PROTECTED
