`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qzQZ6KCsjTNQYfKzhmrvgcjem6qvXsjIg5WvIcykLevkGzCpAYQXyX2CNMASiam
EB/mEEPMlUd2H8AoiyzOlqR5PeBl4dm2Zv+zTvYC0TFjEbSdKaHJqA7GpuOYVc9p
tXGK5QVyCmdxMtTafMAReC4aXYXmXdDgISrpcD1mi1ABKLV61E7D7iyIvmfFI2+F
SHi98BTBdLJg2CuHNzdLixM+ff0ulF1ecMXCRWXZsyYxR1FQClXkllhKSaiBWzGg
VQiYgbS/B5Fj/lF/znoz+1H8WArPTgx8npg2XAbewW12q11UtymKMgUuP1GpC1+s
oAZR3j9+AKGiLQmk9XIJD/Br/BWa30BTna6SeaImVs1DsX65KMxTAStGuTo1MNG7
HdzmxTa7rVvOhNhn26Nu3+1Dn94QyIGM5WoykcWjbDE2W4nzu8Grkbjq7Z89xRCj
AiV7beTzdPpNe3aGL9mEDJhjxb+VLirb2LvQObpvUBFj6GVtaqJz1sRWh99vGM89
1WXo0ACR+HDjkcj3mokCB3EaAG0pCA3zocwrDlgC06eqe5aMKmwKtcAOOEaKRNYF
2H7nIWvKBLYxLtgakNEeGR9WbuwqNkCsr3ot5x3uIHJIhEMxKykrk09QAoRlncXb
Nnvu6+PmNMTgjEzpOr2cXBAVRaXs3iQjbVOePJ8vOHnWLT1KrL0bJTqV0bxqH0xN
0Kbv7V8QMQKZNPdQxIHmPu0QmBs8RwaTamz4g0i6ETKXjNT8GOhehft247uUG1D0
`protect END_PROTECTED
