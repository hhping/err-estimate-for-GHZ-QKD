`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DnFD0TR2mkxmy52RsR9j7Qkb14kPRJBOfspS1+ba656OzbMli0Mn5IsqCV2FE2px
DHzGnWCX9kd695s3o6OBlkQQY6k5UVAsEhWyV8mDezAg8b5Mdx1NGAEJ+JpoXFgh
SgM36rDyDnm8JSUbAYCnV9f3RekkaD5eN2x1K4z1YkM5LcoUjzU6/SnEu0j3PKhO
7NF6Lr35fvvXkRufqg6K2wIXPXtWM2A9h7BkyBC/ZuKXbEVm5Lsw6zEvG717GX9s
mXaRlRCn7AGUne5jW70lDog1BrXmcZypMVH0mMgcvZbtJIEwLaW7CrX8mfDqWU8j
7OgV4p7R0FT8KzkQip5SCFQcDjuUhKz10QEzFYpsVqmw1JOt9lO4WjW8cUi3c/tF
p7fsrIfgSUiZR1FH8QHJ/zoouLdFkdKAHP2ya61HQ6D6v6TS0Xi+eoC2uQK/fQVQ
n6u8ucnrfkNi6745Ic2JfQyS9FL20Bc6sV4gPHUEhKPTcEpiNiF113fxPRvNhwdh
TViwgbJrJ4NSOadUJRCyesZaUfQGqgurPi2BhUciJ3bmOQg2Zzeupe3zz9l+v0V+
POqn07EHyFIpKMeA5UUD2gSfqyzX8f93CzC7diUZxUNDzjwSlujssEXpzCJMdCtj
Av3V7FXIN4gHC5ueeFfaIIn8CSCaRFDWJjFMLi6opX7A/m4ekbgGjnqsj1OSIDi1
w6T5WHL3VSv5v/HKwHhbrDgDwCIs7Fc8RQTJ1KGaxouZGaQJ/yNy/IjZ9XScmBi3
pJpKUtQnCvyY+lUkWf/Avwt7VZNKZwW53Y2NG8xCFBiVUrSk4KbSKah8yhfIxdTR
m+XePNM0A2lFjsOAWzUpLe1UlWuwjbKBA5ki84QhUQK7USfDBc6M0GRUyq/4kmoR
5IB4brGlvXEFb8SDhgeCvNGvLTOo5rD8sI8nmcw6fRyMutUhwI17we4IRHG4QlSO
JfIo5asvMPg/HA1exglvN+So6cf+X2LtVeHy2NaMgIeoNd3K9paJI7kr5mynDSFO
7paJ0B4yr4WpUHV/Kvrv4ICZxY7tJMOGOGEwD/H/gCfVeqSsH8vlBPQgqhc5ZyOG
CH/homM9Hko+0eFUZEdQfJ7TVmYHHJXe+Qpo0EMLpyOn7rFOI5pveH9RwBhZNhEn
3mqRh7aCwPIpDPCUklMnfP5dauyYrHIYC39SUH7QDeJwJ14t7DWVMOnYEdM6SPDF
oqdGDbmEXLj+B4JW8WWsniL6qwasTB8IUGLVjaqGkUoL3NzTdXCOCPIRO9Sp3DM9
nsJjWmdiQY9EWg0VKu6LvvSKiZvLfSwoevyipD0PfMSxk7SPaeXBFicbcZebXVDZ
AkK10hl2h2nqmpkg+Vc7FGsPsUB5W2KHNkkTko6CBirLKGTWAN9MC95g6e7C9dWi
y/QYS5t+LX7GM2CbuCOXFRaIqj7RqNveOcwySQ6l9fzk6rJS/BRvV7vZb5Tj6Wjf
SxzN9X0MP+NVX9zSNi8YEQ==
`protect END_PROTECTED
