`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iVHX5useMyIpSeSyHrpyh52fvzrpfG9dOvE15k1fVn75u/45/ydkApf+6b/1zeyH
WQlJ6+3WS7fzPg5Fn87gVPmYXAxgANjBJo2cjG9egvQ6pWFRbekCTyI6/ZJldA40
Jx2iE9UxLX5S51MHo2wuDWwrgSN8exzVdjHsB0SY1BAbL3LjOzFQQJdjpoerI3cP
r/0k0lGTpCCo01XeO+vZJcsdNvEF4iwj7SgfDeg2L/FSwEutNi3dRvWmsswwN446
rP7lxYYF0V1hAOJppmBdNQqmjIHtNP8kCWQaiGqnk2KmDuq9rOcSyPx0jrO9Cc0B
nj+ZnQRJsbg8uS3PWIxnikqpFIKsa1Yy5n0WhUSy4tZrsHHDkNSHld2p1M9mQC8x
E0sGo1ZHOUjspAPfVkEapXkjdtePW8gFZypNRwIG7XLFrkqzTKdhff83ZLXKGlrx
WdzV4kPLToSK7gIgqtAhkjqQeKGOHk86z4nl6jVKpOdGvRvg9Ncs9AliPLoCZf3s
tLDwXl8ZcnjxTHlVor/JXdCZUsYHumWEEdZNnxt+vN1aGif0gY9A7tJh8+3MjQsP
4Ul1W6SRlG9XkIqX4cpoQh3A6LdtVDFEQLwNO85k12ZjVnPFwQTBM0bm3YH6nuBL
ObQTqsu7ovNzt3zTT0SZoeGtZdgBrjeCmoywxAl8fNQHxZCbk6zkVJQZW3bzEf06
OUgPH3f5FGIg6ugJu1u62Mockk3GbmY8ipJfXfq5dWlCxDY3JVdewS/wmnS3C9pJ
4jn7S9SEXIlhlFDlJ4PKACMAt6zfY7f1TXbrsRGU1Szvb8nD6zYkANWeQnTo/4li
Ki0j7yR9Q1vFRmIC0/rgwh634Xb7TAPShYEdG5NntqZZbx6pPjFIyjGeIUEdYM1P
l3IbwmBT+nuGMn/It1F5Du0oj8lCn48QdijfkCllPtZKTSD1IsnmyjDVdylol1LI
fFvoMXY46RJvE3Kl9M/+xkNpmlJktjPwyswZEkZqAqFXbzkdZGVXYa3F8CARHpdZ
HgKNvplmdJJdb1fgsLpk/qNcNjhK/DliXpEEBqeQh3FfORGw9DKn/kAu9mW4x5/a
hwno7VLP5tHv1vV+s/rkl0t6zBskgPzyEV7pf7fxA1HjbhgDlH+JVvM0kYShOPnj
tD9yjUafUMr1ismLfD3bhLfc3bcTFbR2MaHE2YdISitMFzwS7I8aTQtOILhnvoCX
0y6AfAS7SF0UtPCl2lEe5fce8TV1IUUYb+cZzgWd3NqwZiZ3nbzspkkV8xFW9tRO
4SMrOGpzTW+z93MRDh65HdrMAMv/zOpmqs5qjQEsOq+Z1Ey58rwzbW4JqnnP7tNa
5YCwL1F409r++FdBieFv1ccNlrSSOcez4YjydUNjgHTDxJWObBgQBNLurYbsGgJa
uDZHfkY9PsVojsn+hv0PlRRuUSdRUJQKunk54QBWJ0xpDTAJG7nEyZC8nu6XOgMf
zGv/LRiRQYCqTnD8N52xEtov42QhYjQYy+NkM89zVkDBLyYtMSeM58fwm2bgSTne
27Lp1qhcYqEskKoRohg8IInlml/Kfa0GgdpusCu9wAU0V0sRdR898XSoadb/loBR
tcz+096nfHEmM3lO41zre7Gds9Jtv3c55YxbfolfrvNDHej5PNIYGJB74Ia9jBCx
C4lEd0hCVsBTSaqObPmISrTpyyalDCiYNLmIfFWVCCXP9PLP64GXkW1qopFJ/vKy
IeAV0gf1vxXTGmkMeLRBdl5aGDrk3hg4emitplZ5p6UA0zA5uVX1zrZnZjlhOxfj
ba5nrPxHSheui9asBlcBycjv85zEJnGyqd57PdHQjJ8LFQ4x47LaZluJrFpn497w
mPuQpEehHcpgq7p+vn4LQfnVroFN0HP0C4itGKsVUJXSntjV4fZbPri4nw/Fgi/+
d8eiJc8nq1/Rfs0uf8O2ewCf/D9waTIhqAb1Cp6UQOTqQhoTatHirLQnbGcbWcZa
vI/Qf8k/4O8aJYUxjk4bBuhc1SDqGC66n9FsVvbdM32tbeobQNUQbWEXWZaQWKkC
nfsUEBZQan+gnJsRbDylkmd5eOqZxuOG2n/YBvhLmw1ObPiKWmibYyvqVMd/SunI
+PQWH7Ey40GoG2nmW7bJR2R0B8kE+bjdgE4V8ELC0Ca+5l3uQhHlt7kMhZEv6Khn
pyXN6nLJ5bat9JOgyQmySZiKmjHUNBfxPfsbm4bitvOihACoR3QpzhVb1kc5W8nG
CwowGcizvTQFzd5y5A6FU/xhw/yfbhkeVDR5iXspRuc5jIgLm65a2/Z+8Az2jegg
fqWMX+V3NdtioOgF1X4QeyX7kcKMLaxQSFlAkBkFantpNJPennFF+7NzRf1sS5sf
RrXo+rI4sIq6BKobmA5naotB+2tyac6M3DPJzHSEBhHnyDTraQSAJR1Vi2NHFGhm
hzzjVifUh6UAx3m16DkhPM2L66Svq4aa5rGsk5J8vtvR3osBibAxsj86/YdioGZz
WFPAxrayWdnuMLTiBWx7W3x9PT4yokbu7iuJcBJGMPIMO5CCC+q7hImlG7mhcLjZ
wmNgygYJFm/d7D45h/KVEEAjYv8y/BZfaCjtPDIRRXWXXMS6l1/1pJpItXRjVpBO
838oOKIp+IFLmF3RX48yEdVXxUNNrNTNIAs/vqZWwI2WQjRjiIIIRv9hwG3VLPSY
g7xftVBudaKHOZI45VIv7/7gCT+oQdnw79tUzcgMWdIjxwU/E2N3jwI3J8pdYG2s
irOOVm1cTczfOqsQLmayGNBfsv60vsyJ9Qurtr/1fiKReS3G9lqMWzOUdS7BIyia
Yv1pDD8KfY1b8NOy12AfhQtUD6EGtFd0oGPXisX3domLQuYp9uGmKBXp5GaRRjn3
FZM0okcw3MsE2A14ddVwcu45BSSbCJY4yBASpf5qisQCgsENFicsAO+T8t2iDwKV
sXCZ1k3xUwOMmlviojIUEIoBrOBEAPaWPfd+46pbYT1n7rpdsWkexZgADsdEJ81M
x6k9dnGBmgAYvYCG2swEYkYUogBNS1oO437X+jZrqYw9E4OBjxlG/9W9FPmtEeLW
35Djea20j5xE0Axnbn/mJ/KMn36Yf0YWo4Zp4oKxsjLFEHcKBCUvl18+2B3cMTeq
DpZki0OuSwqyvfTE1YGx3nhe4BP1esgqT943rvAe+NISSoXQpItNPRQ1Fmd4m8kc
niUAe+1gWtdmbz9jm75pbQYUrZDKjBbjKRecBj1kB+0awR7uuEN74HdXbGFxp5mv
4Yd/ypLx+ugx3C7VLmZFtES/1aaaldK4dqf2ayQB0tDExa38pcLm1ECzTzH0D1J1
PfHCroUWcEhWqlGLlFuT544pf/R3Ybce34w7lnnfjt5WxhUZoq+fuT51CUPQOKUf
C+vOoL0b7i00PWYiUFaYhyZgV4yC977rar9uWbLUyZeiXenj+LBO0qtVtBpGSniv
FRaimgmKEQ7SVstZDH3iwrG8YaimmCJEOKJwdR1ajS2TloEt2JfdiTiskweQ7oQ8
phxHGvPcfXqZHSSSWY/b8wBde/8t6MrQNjag5/XvkKa+gzruUVgegk18jZT5BicK
B7tjVeqsby3hjwN4BpNuoCTe4p6h5MxaXZlobqudwNTjk6vz9zu/tJgBa1SUiriD
vgl7EUOHSfeRPunqfjdpsG+xjDwzDxO4ClbgfvP1VqqVRSthbdNFn5CDKk0YqBWe
vQcny4B8QqEq/TTopGZ2IV4Rx2ll4EHMP7UFlTNMwWaUzoXMLpX6A5CVecynUHhb
vOaSl5/odjmYAopiQKhOoqBejzP/7novnag2V+OeFY12mGwrSHI39EQUJBTBHxY3
PgzgClfNBI0E9eugGF9sVakaD4i69K6QLsgPpQXaiqU7cdjcHndRn1MyQsqayh6I
KLRANmcP9+8nq+hyVuXozLMXjrNomC83yLk5oie5flJbgt2eyYAMlDfZG2u98S11
9JI3LaNJY3IvUVBWMkbb7nQy0kKTa35i/OFqLOe6GmRcpltY0DcEeZSpHCnFzU3C
xbTEOmnS0EWBGc5Torf4nQ9fgxqhnY8pKyKJhAdYe1N/dLKfmg7Hrtihc95Z4kai
Zxy7k8zIVIO8MpX9S6Xf0D33TV4qsd3bRE7D368fjeeO7jd5K6kjVJhW81zZcKAt
pI5vo4vwUVpVNTPBkcCF6QfLPFg6GcBHRqc/FgdrhPOHbsW2rdTkQRo28gAIphGL
U2NKMJCIlZy7vkruxmZBwEPggeO0/tnsU1kBNtD+sZ3gNFMRV9aZP3c8JPS6iEn7
607h8CLvd/QJyCaQoqMjVuyzYSEhnYpWwXLCVC87kt5sKmYezsUOvMrYSTs8KYpp
azvbzz7uhPxXeNB2GGM4SpA1Irwt8T9U66Dsa2X6nV5B5NEbtp41u6gjKYyjCbHM
9HKbH/wGiZjXshhebyFNF6eIjlsLvu/UaFjDbPnqHVhLEEsrpD00cTwtlj2h993T
CvYmGkrSCNT2mGfLYgcIJXkGstm7ayJe66xSAB0Er6zpDHm+e5LWeITJLlBf0wZZ
Ir15KOQ7HwGDx/5Fz7Bevsv239ds9oRFgilrD6s0T+WAYLrQaETjfEVpSZ4tqnRa
lmwtCb014wTiCi53tRw9yUHmWxrxiENBqFw6AwSP3kCe+reVkChTPn3jZMZ3T1D9
ps9QxlVygqPM+NcimIj6BOSokWcii88zrmu+8FS0db1U+UD1qGwG871egZub87Ej
Q1LtEh7DJMvlMOk7rZzXFp1CXFUPKVVOaL/3BJu1Lqr9FH3rNYjW6aUMT22szO7q
UM+8Qdy9yYM3E+Z6L9u67EQigoW3o9pNLe6bbE4RBEpaTTiGD/8xBcO07PKV0bey
yew6Vp4SP7HbbNznoG7Mj5IfE0huAnYgwd/MBDCBurm7WhZtzXlTui97WakPfvqo
rk7otAv4kr9fvYYqUhTurQmc/BOEF9l2h60fhMNMJ2aMkUN4q9IL7Ox+cOufOOv9
s6EHnCYFcfaGrO10uhcPbtPiiHCkRWg+32FVLmTqup6fsi1rw2Sj3UpDIzxGnVd+
oxgKJhgolsbJluCO9E6fPa479APtsPXSPIKtsWlxBYdx6VnntpZ1ruNICqUIqNiz
Os/z6OuXluiFch4amBJwXbZew4Wp+Ka/hhDj0qS2lbaXy5pu6nLEN9I9eo2qjnd1
vsrsutpvUTxWoen0dp7Z/M1keURrsPn3QtzGLKJSuKl69JfXurzl9XBNPBNUBHGm
I0PJ0ijb2ZMYO/PvuT9LiIUbhfefSa505qHcNfgtvWf0dCrluzz7jsa5wNr5ImQP
L1n8O55IbOUTJqs9JW0Q51HZEb8Vy8LFf8T2zutSDTVs6aZnzAqVdDouebFUqHwV
UQnCH5obAMsNpwtotXh26jKHbDmLsfZgdHdZaNAKS51HteCwNLOikueJHHGdUOPA
5J6tkH92WRhu82WYdiORwhUsgAHWSsPZR1WaCdiVcYxaal4nM9QbZ8kaaPscvKgd
rjLMhrZVBgH9M/keFmOfctm1bIPXlOPSvv53zggHLw9tq7OvTmHHpImEG7LSuQje
YVtaHNvwRX1bo83ad0GzMrBLmK5PdREDtRbG/EibwymS8mkkBAfiDSMUC4aAfqIp
l6HAieriTPXibZGh3r7ytKUs37rUSGDTiG6NZuy3CAGV7d9KHVs8hN5Yrq8xsX5N
NZjQRMD3IUZiogoeIpeJfQs32tcEmS7PoA6pj8kMEBPWOP/9MkwDP3+FN0f9gL39
eQAJLzKr4tZNmx62BERBBMjoZHy7x5/fViS5HnvlVp/oRUbrI/EI5k4EMngZL2Qn
VQIU3GQ+jYheHm7K1eotBARLSvwkC2HIduyFWTjHKrFQgIaFUf+pyI7gpUoFY/Cc
5khZXfI/OoYs4TsR1fZpL+p5BOHw1oyncJUosnkTSf+0pFmPxkmqOB/TiBY9psWF
YNMe6wFEEGy63ZSqXr/qdPWNZUNYYk4EdIRtNpFGDbjXnCxQ84ICtLwx76h//25h
iq0R79KPjo9kfmvTrVRPTckJFSkWuJJoRfuj1YtFgnLDeXb5yGaYFQtNqhSLPMnD
sfcVeZC2tp9zgHoUDzIxprgxJTIc9C7CxLJrtuPArbkmr7Zwm6oqx1mDofTTsSn5
6taVeklZo0qDky2pt7vRTqsIsdX92IF/VlauFTTQWUXdrr7tE4glq8ITYIHxlab1
XQEIIaTKwDO8LkB/irkgCXxykbgRBQrNGlNardjEhUyqEendbvdpWvl9p9lYecq/
v9s8PJFLHNXRHRoTrIAZtjR8GH3ZfqWUw9pfrANh3g/oDya3vrp3G4fCZOuZSpwV
0rQykAwGp19DVsmD3vFMM+PFho+D+psrqkRuCvhZHAo6SwAamwpKF/fsuZSU3Lf2
0uoPpjNSzq4QloReZfbq7tvNmTq53bM0R627SrLFHrwsq5k6yOyeJ+OisHVlmdE9
T7dtvH+w5VqxNOduTKxEJVPYZXuLi3c5U7cYVkJU+eA4luAV92O9R4yeg6OjRGpE
rvlqB6sIl0lN1apx8tLFtQB5K3aLcYCRBTS6TVKw+vqITaAJJMIFbYG215o8VIeD
l3tPHCDafv3lPItP1qUTJfSKUlm5Ol/u3za5x3xBom3Pr/gkK0a/Fdvv40wnQXJq
RUPFoLgvhhIXEdgnSgS3vGkIczXVtZ2RIu8OONSoJ0isubmxU7ac/uTChGigWs+K
SdEyRr+Z0DCnh+2JiCFc9Z+Ri5blg8y9fmOVK7+SCp0Uio6gKMv1k8p+1Q3JkhtJ
W3iiWgfY6epzwfmM/bPmMOfF3g1LWW2TimSDZfEgmObQceNJoZwrm3TiIy5LANZk
6ii1f+t6qzAC8VPI3PebUcCuEun61MzwEurpxauBipYsgZsD3OpXD06Ev5A501g8
pv0TRKAHwwT0q6Q/Sf91MI3aJjLMZHFcRXw2RNRkGOsM+Nyc5I4KZBiphREikMuB
aRsM4mHCKSY5IHjjq5f2NGivCX5EEh20MP0GJKi7rR2aezxb8S5vz7LYIcBLZE8m
2i0qQqKuOYTgFYKEmve18KlQrrAHxpXFF1v/13g1DH0T0REqD6nRGys/iNkopwfI
9F/Gfy2GFmrtZHWv9Uoq2jDWUV8pr5Y3y0ndMpDpA+rP2gCOCxflt95OKtE1SY1C
vYsXawnU6KTfKvvEqyPhNMxNMBoeQ/3OsKvy2uijzT7EGBcxRlJ/PZujFnKpAhxS
FgDIWTduescSjZXN/KN0LIZu+rptF6W2qy9n0lE9TUQCzysDOEzisggUdFKG5T3g
21GQirDk31r25srjuq2mOyMdZ52aigv1jG1eyD4v6Tolx+YpEdDnLrW62jt7XT4j
6mI2iLUqOOgwH5RkqP+11mqj4AWZMGcw2CXav/BE2ghiuJpa1DLqFWJt+02l4o9b
LWhJyCaJrBLew6liYfrEKIFCDhourXd3ZYQyIwDErb/9TsaeZcqXaIKgt9IpOk7o
7XSyVNW9R60+e2W5AbWVGOSNsXTXCwnl0UZVtEMY0zEbld8yF3NgQHW1o4Qvj6Hx
tR1vWR3KWonJ0zWncZ5QdIiP908eYx+ZZLQDREMPihQZL11r9gvdzRF/YlVwxH7i
cND3fY1DUTVm6vDmYILHWWJxSI3PuvsZBkTYIIPtd54QTWsijqwHHv/Ncoa/kcxP
Sw2I5FsK8wqimm4ajlMAyxgQeUuV85EcpKucf2D+TcDiy+tniac9Dbn4z1BUkdT/
dPS3rFnqVoYvWmX6ka4DSkV+OzN5kN3GjV88z2h3ErcQNVbJgkzDG69u7pSX01/1
CzHvL5rwHrlpfZKDZpXUxbWhpBzPTyZ0CA+buzAQQn7o+4oR7tE6+vQAVKKO5XSv
lP0zKl4dS3SonEJyAeuZG7OgIPfAw3mSGErZp7aw+19TLADSd+O9Zfl50NeZAMZh
hdzrZWJs9925ovpSGRfH2XQGcD1qLhBdyx7w2hMluPybdd+64aGestshALe2m/JL
ZsA8sx14N9M1lO7Hjayr1xovcAbzIL6qqGTzeFYT0Vvn/gUdk1K2Z6Bp7DM6zUN5
9vqWzvn3PlJ1E/9h4e6u7442TE0+H+gQdfuP4MiWC+flPTN27zCqGydGokPHgJoE
Upo5mWk3K6v17FXYL4FRuF3wpWMztv81mj9MVRBQaYGcixL9QHFQBUtBdyfsTPM7
YZM4dJO0oolwBcIOPzbctA==
`protect END_PROTECTED
