`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pnv5gSKpYl69i2IKuI7zUHDu12l/c56vUneBW16KmpWOUOjdYg+/A2NRW9pYNmrb
iStZ19XTQKbaobLKV+XyNnK1VeaL5iLS4DWnBFhW6ywrYhJhYEJwOpCepbQaYF+3
9U2MPojCSMsEuRI59b8qGxCf2REfWQYOv8bD3eDN0mkd1LdMGOw025LWh+EbPAsw
wyNklFnih/UJ4w9/+H/YEwEGWGFgsmgyXlgNTjkWqRd4nbm1QZeE6jTOzykH46Y3
j51b+MH3+fXedp+BUMkzyAFRV/uw3YVu0uMi9e2uLdCkq3xJS5G5f/h3EtcsiZma
QPtDOV8oLc5EXc6cYd3aM3tSFYGEJ+Mro+qmCZboRl4Tx6MaEaELnWVxv/F+JpZg
VnblWJ8i4DlkycUpgqtTRbpkXBCnN0rhcqQyny4uhqE=
`protect END_PROTECTED
