`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1IIe3pFs5YxmxHGdkqKehTHbCp1HcHSCK9a9laanJgAwXuMduw5lzrOh3d6BrFn+
mQVQf9ObnW6q9hDnNBjZmCI7vbAhuwtQ0MsgI1iPYAgLzfBizf8T9WvUyPTjYuaU
OqFEOcisrxTBlOtvCQOyJCimkAInlayivtOYPT8eMdOBCNwKbjB8YTvSesn9dvTJ
lukQOAY5cKuXxTuvoCcZg5ced937K1ya0wTQKDrLtLOXzqWGAmGR/x/iHxwdf8gS
VfBWlf02IbJN4V1dUTYtHc/KuudqPDKs8UD/5eMzI7atv9XjsGGO2HxweCXkDcr0
Swa36YJJl9u46Dg4ZMXDWtSFjN+VH6AUZvV0CvipeKjmQHgBScEzh9VDe0pJdFiH
w1nlllVR+cvKQb46YQfIYqrEvrq7GOzqeEs6+WyHJzNM+giFM4C2T7Vqw563/K4c
QaHzKLB2mQTodZ/uo3SPEYFIWbXCbI+arfh/wXBtKcw1Inwp3vjj6Cf2FcauOVLB
Yt9cfMxnX8XOx/yRAXZe36oV8Slx2IPsRmnN/tNJKELVmfi95flAfKqj780BRnkR
T+RZhmQTDdaIJLinFiiTKevk2HWUJCZyd9ZbHkljDtciFFkZDLY1Sk05Mygd7zpF
vUjwOI4OLIx5hfJhw36QKzjzzcVqqewYYZUlc2pn8Tg=
`protect END_PROTECTED
