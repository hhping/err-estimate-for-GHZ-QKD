`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJvme05qt0PIibN8sx3eEVhmXpSQgW2I5Ci7C1lDetTAc8j51XyKS4qINodcRGhI
BDXhrNcWMpph9SLJJIAbgFpaJ5u0/TY+D1jsvByx6DxtqbgQnsTQReVxzjSg6PwK
8ZJUFR/eyFgQMutngZ+g1rXeuveJE97rpMN2ylChJdE8co31Vn4bfpclDCxBxS3N
Uqm8p8d0Rk4KpdjLVFBKq16y5osmLyMwP8sf1OKf+cwW5ZkvHaWU/pTfAsXCQ8JO
559u21vsWOdoqfOiW1jmCtg0jNjXBNZ7yTms0VunVbTTqkL4rVaIsyIJmDB6IS4Q
VVqXLi6VM0YIZxE2F8jAdS3QXMKVQVXyb9zfCtuNgwM9U9prhvjAEQimleSuyG8X
7O2krJXxT/IDGDqFuC9ye1455njvAgVB8nzlI7no0fNIuwhoIJQOjGQ1xG+nAsIZ
ExxYQ/16Y4r8zFUbHFr647xKkFFSJYs4J/H/0YbWmT5RevndWARx89qRP7IWt/R6
S5RITrs2UPyKJcVdRCsGPk8BFtipf6Qk0axqUNY0aN8NyrZuhm4kVKw4bzC5LN9F
lnctnmFmb4y16DslKvjk7Uo/TQaLP+HFrS8WbQPCQ9CaDL/JpuBSL3JGJJ0+atVq
owQypzfD/u7fVTy/12I2UM4njIWraznkffNNBz/sQN3GWlAbomYKzJXt2NyX0rc1
1EGwnf0d8mwQsepmthdIkxp6Sbf4zbi+de0BhflruEE=
`protect END_PROTECTED
