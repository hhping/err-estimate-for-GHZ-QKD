`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tl+QPT4sYE39WnexH6n1VmfNsIq7vXbOztgp4g3BUNnxFG2S/sPCmokNHHRWjZTH
JORgoe93EauhrObM8IARnroaKdiOj4Pdkzw1xjLg7sz8oWnFbbv0w0Lgbfz9y10m
FR+/VpTco3/ZHvFzSSq+rRRaJUq1ptnBP4ewyZxKOa+K932OSqlpfgYQksNsParv
iY1WouajRuT0Muyif0R1MLyI5mTzPCj7Xxx3VNn3vRIGNQnrZOyf8sk11/zpqYMZ
GjprRle///9Pv77f09hrPtVv50zZSHxi2BD6hLGxp2ZrbMhF4yfjWmtTmun34XWT
Taem8nuCQl7gBke7ZsOf0811x0Fv2RinvQxShSqM49TC0D+veh4pin8KvyllWimD
boKx7HHLB5ZWZk4cdxLa3xpfPDSnW6rDpGvwwOmsIAr78m+tA7erC8bWGlMDcdrL
VV0PE703R4nTTbemtlPdQ8BdogQqJ4llOsGKL+VibBoBI5FpcUlqMw00sx/qrR35
JD3P13BfKyNP7aTqvJi8DN4A/dm2Ng51y7UFls6TuLkMyxfe3bftjE7rGEqHFvGL
e+h1MFT79g5wSM8rE9GScenZNnUnIP7MN5xWWfESQFcMCc8/4apoDshPQ+l5kkZz
T2qjdaZIut7ee8j7CIWCcnv4Q2kDQxxJhfs/9zUKjIqpdB8oug6/p3ZfAnrkZNGv
FV7kwtQ2hQmfUZtqFg1Lsyz6QfCzbmZsCRatmmQiuQvtu6rkXWzCZJ6/jrx7eEm2
we2eKBrGaRLcWAsZ95E6jjrRPEC3awzfGufcw9Bz0zFd/hToFHluVxvVdurL6j5L
`protect END_PROTECTED
