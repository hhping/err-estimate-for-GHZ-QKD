`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJM0o53G3oNKtJ6zJTi05WERHIAMcVZpBFo6j4SS3g56qfCnafqBSYKpB1BrHnG6
zN05K7E+PRTiGcFNqas7Z8CbtgQm0o25ApvG58M6qUhm1Py+EZT7CJpiE4cFUWa1
NZMr+LijdrbYxCWuitrzzqUiJjs7YXvMHYWGOQrAgyCQrtjugDoO6Mswli2bUzgX
cOZptlTNBkgCTmP0ZW1h54itquVE8DqmP88WDqPNAiAaBu6n4/rC/1Fyqz2brHZQ
/Av+TdyfVttCyf7DZ9TVmKdq3RB9VGp4w0HmyxqOfjDC+zIRYE0lV9tB5IJ7Gp1Y
ok1XYwiczEd6lJePw5TP9SB0WedjX9zqxLkaZdyzzfhzmgOoUuATramL+IdShCjs
5waYcHA/ItWsG8A5c2OwV3VCYpUHmwCmhYk+HrGzNkZRP9H1D47EoAvPYYSZsztV
fed9gwQnJFlEmtJvzWct6hyEtUG6TN6LN38aTGYb2V1lxQ/Yy346P3g9h3kfBDfR
wH4wZJjXsIQKS4vBOKUM+pDjfxptI0bwWvlJ9xShpSVc0i2DugidIjw9dyWYhx3/
JlHka3C5ibFnaFSjBhXoG1YITzUjgKWImHjMXwdd3TIdfZ8kUqIQXyFKxI6dGCzf
++zMSRzccJE0wSTtH32vr9mc2X8HWmhS/5lq+qdW4FXBs1XdXvyj+uXk4k3e4LsB
htR46JHXRRlxKY0QxxEWDRuP58oMglrYVmHHtoFV4xix2eKWKA9yBZn80dYUzXxb
U/LSABVUZDYJKF9vE5YtYwa6ZJljjm2rXx4KXp9OayTZYu8bj5c8rAlP52PWufBq
b2GUiMluifg1D102WNtLDtgH1+1mJ0/ru3P2q+brkjYUk1nemhKoi/UDrpn4MOLd
nH5VhaC/rf+yYasflJRnhwQZDztt06w4qrOTh+NeBAvEGsgA9xNA3K6UL43C477n
WSxzYH5rMkr6svij0zekzhEuVjxIdrdex5zShbNtD62dilSRqMh3ldumzbL0eQ2f
trYh22uHToKNDNdfhmUeq54K0e4gY4NCcpumwMTBJcooGiZ25QYzg+BpmR9f7C/D
`protect END_PROTECTED
