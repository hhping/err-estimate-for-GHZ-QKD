`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGmIRjm+xt8CNsmmYmEwrX/PSNlOemwBQRECWN1qEpqKzxXIHgRGEC/uDC75lL1s
TA0ex71b4+JcalvTPbtWg9YRLOaVt+1Rp/yjNDWh4ppcHoSCHfrfexQb93KQTrSq
J6atcZNclB/JbTJg+bWbCkRl9i1lBdD0YPE8Z0a9Iu1lGQdpkB70rol1msf4jSUv
0BE3Ccz7amZohYPZEz0hgOmkzvkZrvfGJ7sHpTLb95/LiAfkFcWEf9VDNBwgfbck
kdBuUZYVC8yUsW0jMkGiq75j1YQhLrDBkZlQhVsw1fPQnc7yomMWlx2qjewWS9WM
xewbjHLmCTBdEbTMiFjoqUwMAGxjsEPR7MFIvMV3yH4ZZLJNUIZWFzXlnd3LH8dy
k4zRd1LykghdNEnhqpj81MBK+EIZASZ/pYDN9+NpiejO6j/5yeHMLuxI5QsSemBZ
7IIJiQCEZ+ESi+cFNTGWH9AMlEVlCcpMKHOon5zAvAjBcqipYUeMgrRp4KSTvdlh
QpInUTDUBks/Q0o6Aift5bCkQQtButFMsK31b0QsG+0O+xF+nGLhodvaQbD5ntev
7Z9Q444YJiUmCB2VtIcH5hVLc0yKJ821+hgZK1iW30zUNKGBk60hqh9mKkD6sBdT
`protect END_PROTECTED
