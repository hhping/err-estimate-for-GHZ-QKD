`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTIARzfgKuYQ5qm97BlWY6Tv0dp1jOJvF8JlGi6AZOJeML+MagcflAqoegDFwWgq
P/82ZrzXTe6QoCb0Z6KcQYo/V4CgRYZlNwH32XPyrCRrAleSwLMUEV2ApRNyTwrr
0h04zmCKMQ3kqaTPBLhz0jg9/QzoHl4QEk1hfFZErdLnMvHFnZnPp2bKOTmHMQLR
CBUHqNdh2IqRWBjXltBVJpR8kghjDiNcd180rKT3/y+oluEGlznZfqPKYCMmQQ7a
nO7ay3oDbeI5n/7SjpkBOKTwv+00ZCTkPymejR/Oo+0vdJG0GVg0dEldJL6k4CsN
32olzgm9XeCWdVE5c+k02HC4Wve4QQZNJuR+WBkONltsXWdk7K8Ytf8ZcBFFdb94
Rb09PePQaqFQQXLMc3bUPFkNkzGkfFNZLl849E9qyEBEddh3LqOJIH5H/OD0sq+5
Np3hf5xEFP1mtKgjLgx/cW8+95SdjYAEGJR8blxzpOYfxeKUXZHpIeq6YqcsFTgk
n+ioGokZMtPCi9SeKX0nl+d2wQkg4tEXWIlkrVm4cWF3ZuH99UBtyE7kIhlNAM/4
EvdqjLLU9AnJxAoo9pgZASJR7l4Kuh6ZK8oYOmJtHfon2uxxDQ6y/SRc8jDqSQ+c
aZ19+O4ukUS+Xyrj06Ze/ilI98Xu+qzXU7wLG34g5WmBiK3uEcOF/eO/rxz5NAnw
HRdTDMnf3Q8fWeKLKcP/ew7v2wg1ZjEsyna5iNdwLjf7fhh7rxW7WhzF4TIf+5BS
PXbkTh+IVDYQUiV5TCH8ejTlQILCaMrIq+2/IO7W/m7ZK1xXVBserMgAdnlMUSxs
RTGYui4VThPwXCbeUIi949wdJZ74ZyINaaD2EGWvfG77PSIbz/DKv9Tak48Av/A7
Djx7wb2hVwYdPtFtQbZ8/oH7vYqTEP4zj+Mt9+Ztgy87a1wsrtSqa3SWTxM1/DHT
kshc+xcIOG0CmX+yroIKVyuvKsEyT7Xp2uT+fshBLsOkZKZoy7iDdpjoQMOsze/k
8bb8crU1nat1ijQf87g4Z2rlenM/rKgV7qTCDwgkKK6KBx8MrAnamIooUQP4hd6P
ei4Uk+famBeqziJ6g2hVpgnTkol0v6UrgBwqcHZolh05odS/xaUPSR5BIbEC75Tg
8NoX2NtCgs4w4ooPBR61Hi2LDz4yf7onju0a+K7mfG6FT9wa4UAnf9y9BxrYi8FH
G7NSXJ/5sZzjC2OR/ycDWIF2wnFiS6av/JQblP6hLz6yp3/fLMSao+itWIc5/sw9
`protect END_PROTECTED
