`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/GsbkNdtsAENpK5PbJIyX6D1G+E2myWg43wsMg6WOASi+zPGs4n8DjgKpqz/wQL
UL/jHrydTIkWm32eJoCvdTxnhAev/rU7qkx+FYAaSHP0Lu5WXLeWsOiTk6TwS2RR
xoaKZJwAtu7r2EOhgCYc4ewqInfwHy8i7mp6Sy5KicrOvkBVp+mozBjjcvlX70yH
NooRbtZPmW+0Xbn6hSm7m4VKWItHrFa4N5jAIfhgtC2l70JAdIcASNq/omum6fSX
Yopvhdb10XTqvszjA0AGEgfbnDERL2DvGVKyCzjst8ZZ5TfTgGw7fLsteM1iMT5N
oteD63tUDMBoyE6I0/xIZMikCdcV1xq5C5GkBy6owpAUrphnQth4ayC2eUSyjVOJ
ilSVN5PnZ2R8kgEPErfB8GSsapSwOpCQ9rAcckmAYm9jPm/z3xq673hwE7uxCghe
HPqMCZkFgD/Yu3QdXHJhrMSwYym86qI165tbivMkux92QCHbfsUuR73gqStG1QFg
f2IA2M3sN2JP05lPnN0Yc5xJOwRdMKWQ5kPFpVi3YFYlV+wa43CwnAlvu1eY59xe
28efWPlZz6dCI2DyoAR9fQAlOEhCyEIAEoV52DRbV84VhOj9NVkz7darkEHrJzMz
ZHU9ntn85zqph3mA7E62mGB1jc9KcJERMSJrDtElOWk=
`protect END_PROTECTED
