`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eEK2Cq5yRKns6ZARqjwKL4mrx6SV6EjdSRG6tddp+CgWXrYQollUpnfi7nfk6yAB
aszZErKpkRIqcAySan3n/B73oSeqlhUATS/ksdjJY3OQwt8i8He1KuwMVn3TdWsL
6t9IMHauiqrdbklH4hJRZmzsR1IFggVRzX615ptrYYCCP3sDV/PkSImgBZPVMEw9
/cAQmkiMWIYd27MGF76hEAfFpLyeaI2R8zBjB9xDJTEtiZQJEKUZ0jBcxJ3f0Ka+
rTRtTgGN2nF8LxH7WwdgL4foWwq87OnzOglxS5MdbZMNmk7xPACWLYc6Dz9MSgvQ
Ce0880XOgqwkAMFZQv8v6+P9piUBwsSBEZWFVYRG59SufnZw51XMUKidpttUu+ef
GXrn1AbK8JbQuDXznp+78JtOkr3GR5hnewH4jwW+Sopj7ik63r08c8lPauCkctkZ
JSLart0h0d/MdLh268se1plAJHtLd63x9gXIljYU8h6ZmVHsMDpA/Um+8er80/76
C2do2aBpA9bCjqhjBj1TFb7ZcLrM4ncjCGHJolF9JAQNKu5oqBs+x1Rql7tS4ZXq
8tnCdY3/y28yzM0QzQkiXUA51lkj5gEWYjt3f1CD7im9JWdjCMPpV8knRgcAIOuW
jidNvBtq3LdT+PboiIXgugU7rTHTukD2ZYe7hHeKwUwCnqJQHngHxAdZLDM8+kV5
RG8aEiT7io7U2A6z1dvsL2k9FyxAQ3+GFda+qONfvv3u28KqPMWo5RsVQ2RcYnSl
q8kAVXMKbTqzweokHdRje0ciDJ9moWjf5Cy3PgTQHUgU5UT3aBYyKIAQmuPeGY7d
SUDpa5Iltrlf5fWMdLbkF/1Dp2E7WMRX9864uA2kM3bk2jc6Ds140zu0+ThPo66A
xT34SehYAR8C+nL7Dw5+0Yg+kYktt9QvXRjN+xhpJ99m/81awGEeaeKzq644KouK
txjrhVE4XMwXRw0xp97SVIvZBOn1pM7z+Hu2eCZK4/MyBmeNZSXtcKhmWwWtKohX
xvi/FGsm2h6snvj98gVo/4FcKP3Bl0LkCF53gfbFgU0BAfQdfAHdYTuw0lxX0e/8
1bLZKHntZxHGgMGFYipb7w==
`protect END_PROTECTED
