`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/i1yvo7/58gdn/uwYyJZyyzqX7hDkTVh76o6r55GTvYkM5UKl2LJ2esuVYRvknU
OqoYp8czRQ8yffVNScqOm3Sw7dktSew9qTeBH0ASKSYuxzzUmvR5tH7nwR/Q72f0
TMM8qJGsgS18+yWYGCm1hSPxzp+LDh2XCMUNnpJZKY/2EMwxhEQlC9Yb8PSe4aDD
V8i2541GXi+lFws+XwvwbLd6aTuGJsKq6fMNDP0CgNwXhahbZNXdO4ZoNSdlCgpW
BAD4M7st8BTFPAMMUaMjKUIemPKkdNz3FkknKgqONOLpIpbzZMcet08OMI+x45Ld
/BkanJWhb9/q2LX++BPTsf45eTjz2ELOJ+QeS6QrqPECNXrmqEfWXN8J3XEjYGaB
N0xUy9mTTnQjBmqIzERJrDEPtxbQ99YzWpKmWm0ZjTe0HqnQ24cOKHM/NP9uxugC
Hddsr7G4+bjxUStzy9OKnRZ20OmFqYHqxLdWFiuLa/wtHmVV7V9owJsEHFooeXjd
UdIunecBrqPOyKWslmRY8mA1eJxrYfqiFJW4WSG+/+tyWyvUgBbkx0b03qyG0nLq
Hbz9xgMlJP8SJctaY67sUOq2GBopt6EZ0eZlQ5fxcp7ba0HKR2aA6ap8XnxO+653
AMArlhOb81zQKYe2KCQJMl9vJAKNJNgi1BpWBVPdjt36YPZyXph8m4Qal8nxR6XM
X2HqGdhWomTx7/xk+6HxkJavQqEegxLBM6HHSabwTxuUT/IlTxkeEsn7d0tlHh0f
nCKxvqvdnFxBmP0vfNP3EEIuvh6GOvXk03ztggDA56aKTs01vYKi4HZZKgd/TfMj
ej6Qdv2rG5X/p0RkcalDtKU3whpnz/Y7hnJAYPAazf+jOllxqKvh5lceGUuDUURK
c83Eo7oQeEqDVltdpHC01PmFX5x7axY5x3y0NeijnkbOMBAzNH1dwbIDSL809Gj6
mJV9LTCkcGGfoZ7Zhr4axQBn8gyqwYsxVvg7WID4wzEq9eouu8e+63gw64D0JPXi
cN9e1QcBJBqZ1Otu25DKIlDC6GKsSQ+5bfq3hjM9of5/BApZdrpQ+BfOjZjVplsw
vRDbfZeF3HOEpmNPvzbQTk8tS2kcgJZWDH+CRQNvT+r0SirOSWKxlVCC+S7Apra2
6TNuu0q6+klw9/JqCvFztou2KV5KouMFqzIlbFdsMWRLDfgQtj7fx/+Jsg1cUh7B
asC+jXmOiEinA1qoVf6tQrOYCKYLv8i4M/OsvK5HVn6aZBek3vXEkB00HH1P73Uf
gm4l9DoOxSJXGkN1Nrv0ij3z6kUAMF2wn0qVmAVdOsZaHfUIoA51VuVNWXj8f3Ec
2HFbaiI+bncTTweZYRE2UocrvT1o+jUTcbqNgjm6BMVUZnYkguNKvJmGx3dQ5YLn
ioDRAPKhqe7mW96KFVNGqn9xtFYIw1EfdP1T+w3Zn8I8m+mogluuJrHTw4CNHhoI
ReheS7R5/v0JQtJ2TZ7J/yFupgIknsGjBNqhvm1MvSOe1aOYsiK4mxF9bnFfuiDe
d/X0UVQJtcgtiLPH0eVnJjSGUKNDWu+wIo1ccjDJt6EX9RTyaJvXU8GCCyToa29C
CNB4/26EJTQa6IW9sH5nDrI44qv2+Y0sQU2hx40i/wH7f2GWplyhpDLq/bwHF+0I
4dexeVBom5OAY5t5ZucmM1oObwhokK9NxXvYUem16alvDlGXH+YZViRsVyuZWxHh
j9DcQRwghowZ8YDYTzEdrmo4lgY9Mvy9fbS5Ip00FWYK4VKWPiT6gdctTp3To6XZ
Z85CUuk3On5JXoUjuiy1aek50qmI2TSqyr/Ej5qwaGxQO6cY2PlW1XoM1xpwx/yz
6Qjg63mzJsDh+pOOeaDIvqCLXprvwcU+7aO0HEs9gT7NwMiCWLli3vD4igdjec1u
1YShUjHhko4pbeisU3tKLVyLTF1zE39j5UiZYc92NlrnblT5hfpJVq2GFRrx3z07
yW091YbRjJIWLX6WES6cxqalFj6BXLBhFekr8wW65C+men3lJxVjLUjYn0NS19xO
6pwSkCAMzCziZNZYMGuDz91fm2dlxCRiBBplUf1czKlKZJGohbYspVEnEJRw+KFN
z9Y+Dr/r/dStON/nsvlgVp/xrvtTUIjt1tjunUNhiEJEG1zls9LBaQbmq/96s2m+
r5cBOWxD30U0OzxOFRJ5r6zwZIJyAZWnYV0ybIo9hRDjIpKNspiJZ/cpa4YGrnLw
YWqwU8u9IhanhtSYYcSNhUZ/8WlsY5TGcZXUvYNa4RZtrc8PKXHt9GeFnKBBbRr8
LAj3t0wFNfz/Xuuu6to6C8GNqIW+SSaQYwRQgwh+0sUqlBsrUMPb2iRF956Fi/QF
lEROOnJwvOIss2vJBKO0AuAp7vAibOla6VzXja9HBXTeBUq2KzhQ9K6htRRPVVvm
InTfOeDFl5CFIgWqkV73Un65xZeE2Lx5Xgg8wUHL9bYvRqFqT4KLTnRjDEcrokWY
YsYBDDkUdPaWrSF8uYNly3i2Yrh/0OBXRhj5GR3DmjhxnuyQPwSR8WQl8LrXOP02
y9WCi+Y4P3DySGR4vmvSrVRofoBhOj9JR318ALLRQY9GklmeElEpLopS1uV5Onu+
olk2PfDetwXEMnTaT1ErNOWriq29XkT9+R7Wf82I+TxFZzoQDfLjf3pldpFIiT5g
gBbTJpWw0mFIBA4SMdsV10gcVLp2g2jXNUCbClrzcwkhhj4+9FGGAGYESebYDO0e
vs+wuYKat41OR6Uy4o31AGsZghRVqB655DI+Hz1Dojg9HjEt94Bl8XOqdDkYTa+7
kWFGTQmtzSnlbjXBXjhnD7fJyaz4j++ze1huyqeoYxfO116c+2+Zh49DcxYdGRpq
T55uumtkhTg9vm1zpC1EkJ2+c0PwGT6KT3GmM8UYfddlw0/cNCL9qmXqMfrilYjL
1yoAZzrpPDSJa5lrV57un+Qt6b3bXD68LDkT+nqO2M3ZFsJofgvlGt/gRzXJpPhM
mRWDmW3ffr4eFoW2cP79WdvmIpcr8gsbK/8X6MXv7Gx4PKwq/lViBS+WL63aiZX1
OlFAwl0Sh2XJxnd+0eySNR9Nv2lrEWas3XIfGiRG9PxtthTVPKZBYcXmlIWh2Kli
2iSm+kIx7/s77IsMsPP/iGIUvwDltd4P82c6lUFKK8B05XX+bkrw7gdh4IhPakgw
kV2uDZNNpeWC3kzB3ccPRw9ZjbJLkvETnrp7B+YHe7pbp3priNKWOfBaq7wVUQaD
YQgIXCatlIkIZoZzdmIbM8/Qx6mL5SgJTV6ioVNoaUBmChacXWfv4ooOT/yCbOfs
YmayeWvd4oqoAOKGlgG+IL3fYV2Xa/2V2/jRMyOlkSaYdhXHch0iOv50taABD+5E
FinH+Ve5OdgHdFfcjJqNGg==
`protect END_PROTECTED
