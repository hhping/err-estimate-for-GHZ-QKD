`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJEiqwenxnRTymvLrOiYsiOcJpfkZwcTXcPX9OnbnhcTe9RdNM5OCCbjRaX8lBui
MOrtXbSUVS0DFm+nSUHOLFZ+Bl5u5nel0qRHXpegAFiRWc5O0zZ3k6A3PyRUhn5N
IBjTTPpq6KddTY8nWwrSBKrgYT8GUlyeo4B4JU1rYc6VJfbwZD7KPtfqy/tIOhMc
6e2nAeR/IkiPpHWthqcDmf+dAkErdnt3yU6zwxcGRRUiHZW6+rqyDcsGIhRDQ7f2
fAvm+mPGwieFobduim/w6mhb/Vxm1hb4R5HLcx0lcORS5l6mHXqq3FQQ9TWE38m3
qD18H1YFIuazdkbhqz04Ov/X/5ybHrJgxVVqGXWXlMIGZ9kWbJQz+N2mX3kqIcze
f0hlM5dcrfp6NAYTVRDP997nGgaZ0JH5YlbaMqPNBn45v0+LhXHqeH0TEfAky1Ei
10jb0VuDDQJYTfs9djneS7vIKxbRf/H+yAfIVRvSySIpkpKxrFnOeFwvkZ8FGnRI
oiALMXXjeCiMgKuxjgoHyBk3M9B64Z2lMhy/Ufkr+MfESb1z2DKY9+BnryDPQ731
GnQOeNy/BuwBts1ajDhyZRtVp8WI8LgvqiCoHEvZC+GiO7SNzmh2tP0DUneRZTAh
LKlZ7pvKCeZ6tUFy+ASaCgMsja40qTrYaQa/WxrtfZ6hmJ9oDYIAVpvG3q0ycGeq
57ut0WQqxmtqcGtmK4qHM/TQjsQTC7cLxiQTW/RQxusgRaQvlet5zDKIIhU41MYI
wNF9tUjyp0PwrZ3Ny+32c5paJyBeGeyrK8QcWocxI0A5VhopVnXJyfiP65Brn/bR
DTAUd/OrL/UA+J6Asy27ekL0IofqOcxxstT8/XoAO5FRTluveE/z9WeUm5ylcrlP
y/uhGOrX9555FTaOysbCW8rtv4w9PRvxl5fZL5fcjoDf0c2NJhe4HQhArf8rjD/Y
rYkhZF4HCh0aPvkAKVg7eHcDtTopi4WVqQ9FrPjk/lhT3p4eMfm5Gw+9ZMwBcBzh
VWLWdIELGS9GNxZ00k07QXxTf7V7V6uJqilr4A61OAxV7YtdebzxxfVfv/wqBKRG
BG8nC/ryHedAgLc8q9chajUSoExGcueEDg05t7P2Rsqm2+P6ocFqQUzUxbFdpstI
HO9780579KFySWdJ0+BJbzwk4f2E8nHnOYukNO4E44lSvaK61vpFX14020dESJ06
3YrVvxb3zLAUbHMogUuJVhwP0ls6fneYqcGuc5cubO6pjGp1iW6SLGBkHzTzsimT
LspcC6sZMXezOsYEWojWmnynCAPG1D0IURLrHhpfW8/FEkt26uPcS/WC3cuXHRs6
HuL6/0Xrhk29JxU6TS0jxuBxIWkovZ/SQ+tVVuzF6zAycP1ZTuhLe1yrPr8RP24J
eO12gwY0cjNyjjAqB08YEjlm4RCwqUSASUeQEY9EGr5ueErUer9H1jiuRVJj3sAm
xzWA7XVMfVfjzB8msN/nJAN7npSJtsmNYRzWo1JKrATb3GiCni0frlE/UzqRBS1g
yDKoUGq4f+CMlxOVhxWbfiOifsvY3xw+Rz9x3kZFDb+99KRP2uU1B6fZ+lWhMhDO
u9nIShq6/AtGsIo8FQ1a6g22gtS3+mM8dffn+GA89l0Q12u/BFsNGR2oVW9LwLuX
x2N9DtN/qX5ReZ5df1M9O7pJjlsRgWXddlrpzChn9YMnakO0wftJB8ofs/Fil6TS
586Q1PRXx16GSCei68+V7+yHLSAQhjaUORZtmD3zMqP54sT1s/9PxNEc7NnXxuK0
MFKEUbrCLc+t8ForaadP4xtyuQY+4OvQYxQWVRlXROC9a4DtAy8SoGtvByz9d0/N
3Keo7/e0mP8yPXNnvgQEC4FtNB9ufJZsy9yqe0LYAweYEpCefrWbH+VNiI1b9JuL
OwK+5zkk5r+sSLTnUTLJpyqmITtwnHyEGXA3ZuTq0Jhrc+XTam7Nu+fyzUkiCG4r
XWkAEp/XOVHo+4+VgM1U9wYookIeoEyL3bDgiLC8/aV+Nxpxx56w4kZt0YCzrRH5
OEXQ4lOzKvQ1lMPSOjMP0Piy7EoBhUtflVA7A4qJ8xcSHtTqbpzuoLsPbywuQ8Vr
vvgKPsQh62pg5WGM6GgeT5iaKRurQhytdUaDdrnGA4K3h+fFqmC22nfqUFK2JK3a
IFUYfYzA3+xrTgQmo2sI/wwowPrcVJIvDkMBOg5jovbdCF4xgkXYpQPdM13btuIx
akD30icnNXRIRdqN7W8KmiJLP42/8jDvbkjQZhnICJ50E4l/uPUhT+hhmcUlzXUj
qPfRwC0s7kZ7NWK9O0UQhwD4h71EMPOysfBrRhWdTxI6uA9VVHgeZUT0z1DCwa6Y
4zzByhnXMoP1R8e+p06udGcW8D1neXfFCJ5DunZCaEbVLeJormwwf+wyoCXh/Ac8
v7mOk4vIK+lH5fpWikrQGY9TVAEK+cQ0x/Sd8pMlreTdgBHMWmP2aHO1pbJNLH/+
rqDiDcbshp3CU0EYdVHav4TZVuCQc1G18idZT1OkeYYoapZLeq9871Uu0LSevHAp
WG9/ERTflZabTVPrdG2dT00edo29UTLTvi7Vvb0DfufpTKj0So/DDcwqNn7ANynW
2E+S4COKbM1v2nH3luVBAJ+cPxT83RhYpzde2jn7WmKjf/A6u5COqQU4FpIvWw02
vk44iuzUZvzek93hpUZ5X1+pQ3cN0cbBy6ZQxNoEphvTJ8XJBlI3iljI1eNvj80V
bDmaQo6FftIs+ATBDxohIpoyJ3655mQwKJ8/A2KPzoPxLaBwVYrjbiU10jXZCzPu
PHFGzrcxQ0zuOrD8gCJiRtoQU0X1sTWLuVQ0oj4M+XpLYIxSSgRpTItU6+dWWaHR
614PaZ5nB/kU1u8ypWpz9POfsWpaBxDhAD84ixISOcQ81ITEcVy8wgHL9OkJPQv7
+B4ye5gbvWtbukT6rNZ+fHgVQazXv82ieMGhNm3K2bFmJKdN5j3jZdlYxn7vnE4w
oWR9a9OmesKuyqm/6HTcpbgSFIy9n2eMy+P3FsixikYCo9PZAVSTPlVj4TUFx+Nu
nQIEC/lWI20dLVmax5wNblMTZ1lfpcuZLDMavUq4DKimI4fR+Hr5SmMbwHmgPreF
DPMCW0JRzFdBCT38qVG8ogK7jsaFwfvdJrgLzoBwU/UZvNbTru5wfCDnGVyKqxGw
Bsn09IfiLgmPODcO0e29OzU6Fl3b23dt5WFAkACCwpyKciylEzrpq0pqkB5nYe7P
RhPrLYIcRNL4XD1CdsdgsNK2eVSiIj+nU0BQ541KXIbPyaTe2IrPeOh1dEm5n6Ul
fgTvxhPYY8Z3vNbaqRx2JKm5jI/loiBAB42Z5/+5wCrVsnHSuxpmomUQFi9Q6JW/
kiE9oPSIDUU4D1cwOAKgz9ei+yV96hA4kfRItESYPJ2JSrVGc5lwia37OjQfKEOW
dFHXCBA0gqZuQky4ZlV1wbGxxczb7aBtm2OBNdrnKvwo42EKhgEqvNpUHTzMkOiN
yBjbE0/8nURHFCxoCS2jd7Dqn83f/BG4P1U5Qbeu1by94lWXYx/OkcXQIlFpgMmS
sOZlmnnX2n30vAWNaWEzpYMUf+WPQFkjXyPJpDgeS+ao3txqJ/qgGpvrC4KJ/RQi
PuFDcKzlTwJJr5vasTnfYRA4o7BtrSq2AuqjJqb4uGDTC0q3+VAF/mX4xlnWHWZm
13XTKIiAyN2pCWh6YciF4BFbBUvX3r1Ymyo0doQ1/KuaCsnlz5VC+LCQt0tEx+2E
9zdYmo7eXl1Bh/qVPHrcfapIGY6vKffEnRU3G3PZ5mAOoyuPQPgOuOr3TRqXq/qZ
Q3gQY0kcESvnPyQ6WxvoAEehojJe2gND6m1T/makwCJwVSUKvl1W2DMKmSraawhC
iqMxQhQ3+WQ0FR2SGDKxTvUjIIMEX/RZrpQNTrmYMr/8tttxWeo+JUvl8+ahnA8C
RBifmLGaSyq47WiLLZobmqKueU8072ma3qIa1FnKfdVdnqNZutzuYGols8a5vXmj
wjWDIzUWFfJD1Uoo8wWXtHQwIWz4znxmp65IBydnRgIVhaEAQYWgQaM08qlfOKRh
i1WWiiAutToZWJCJT5zNzexkOmobJpcRh6gPx6BX726SdQX/bkcncFS/lpGQA9bl
HM61fknb5YjFDnGFInymR0CZVS1Tpnscytrxo3/KWIx3XhJYU1EPPBUbe/aH00mo
PhRQ5VxOae3/LzZ5PQFQy9lsImbhRrclG7C+twYdZorQ2Psu9MbV8AKiUpuVj476
NkJfmNivIGr6/6oNtqzJN1eXjfZ86OnkZEH3G2sKwyWilbUakVnEf27tPLLBeaDM
QzcxZCb6P7am0TIbLst7S7iXmbKy7IosUG4qiXQTzpf+3/kTVf6MHd2VLYURARdI
4ocNDmwQp6lwPpmAnRQhHi8ZjxQVdRalb2HVddxfS2McyaB7EtmMW+UzupiRhl2p
FFPyqKaNvqe3asSjpYJaExnM9hqagYVzkQ7aJqnFGHq8jj2tT8dZf5VykCUqOVrS
c1jDF27CQrMdZsLuFmo6qUQHZlwdWtJ7JLqCxHVtBp+e4AVhelZtgegNeqAVYT/o
AX/tZg5a5Z1QXBiv0cl/zSdnbviV9b99PVllJdXPkK09LxQsVYMitCPq/n9dIW6+
e7rWZ1AhpDbt7G0ptnh1pAdIKPoCTA8VcP5OpT/SPDBes0pL5dOuoU/u8e6Qw8m6
zNwLEMQkhP/oHZGf8K5SPjZTr+T6RtxBhfcv23qR2IqKajcADiZ1z78K5a//5d2N
Y5xRaPGTQ2ztrdYYxAFO01wjIZQm/TGqnwD9tJSpQuutxcfBOFXhQa9liRChtceK
PIiNlEUgd0usxsntAd40amprTxQxZq6XKWF3JLO2Yv2XRHt6zspGiBGmTqComuU7
wh2tTkrgZs3PJemHfsbNauUAVNrnyySppFuf3Yw8KGvgTwzs9LAIm3hUrScJTlwx
ruxXDdUcNXjFJFAN8eS1Oi2fplE7i63LFW95cGVn7PL1mPCNoylvOZ7NnEHSlB/G
D/koDq7QvITTzrc1T9S0eOf+7z8MXNWp4XQJWx7U4ksW+Yim+8R3BzjnRoD17L3/
+L1xfir+DN5+8a0bslhxhpMPDVP2yvjCmslKncksBEKE+rWkdO3A62WDSrgnxmKX
GiSQJqW5TxEGHwZ2AFXRWsooVUvVJsA4evbcB87fA2f4MzO0BxeWIafGC0v6PTQ+
5DZnKOy/dcVUnRjechQz4sRWLm30SVrNiRB4atX1+SqZm/9DvfiIqZc4kv0VYA2R
Iq2qRBmzxQH1440uUQrbGmepKN/6IPeCMMkP0zpk4JAb24zop3m2c9wFs5TkQudG
3sGQWRnEHH/N3gc64JIADAcqagSMrpfsRwZltJP5elpGbgTDjUFnJtCyZZpsXU1Z
U4HMuy71VVQi9h0MYYhUG34OHaNz/6G9RtC6P3a9K5xvfYbcd+Ar+8lGfMkiJRNp
6IIc8aXhrRaLYGsvBkh9Qr8vB3DBtt6BtPlHrOOWegauGOdIYpyN8E5FistdnriL
ccpvS2A7usJGo1w6DYgxTwtQKaCpSfmWd+qL8DcNE0fhRxrZE6XyilPxVmjVYihk
tzLG9cZQanBoBCA/xhBwtXfwaxUGG78kmIdnu8jiyjhNivBGiurkiJHfi1CNu6nO
j2cvLoKF9IahUkhgBaKwRyVR0x1atCHZCg7QnCrb0DohzyfHaj9x+Whhx3rU3G9m
cN9ylnPRqPyyxkaeDxxrsKB5OsLNMgfV5ecCyQnKMXzOMbcgUf+spq3yzb9nTCqu
UPzK7PKjStt8U2c8C4v/eMrs0v7hybyGO8nH/faJUfjQL4D2gqzLRzq5Cs9/O/ti
k7zqKBpWBkBviQ+Owv9JRzc1sWJn5lAkGnJw11JNhTALBEqkALDRRVCZFD6OR87Z
fWjkAC/tc1uakETYuR2D9hXuswASMV9/cYwzkNs0j859LEknDKIheA03e+isu15r
aUQGqdj4La65x1oJuKZLzJ8NT8sgNLnxjBOXsGjQmottEra8pnwIriBxMnlxLFBd
MnTdTUIh/hDanV1aAZa23bfZl97xEwYCTVryBasUFjij2XAW5VGSjj3U8wKDUY2e
EHCF/pLb2/8Got6wcP5V3m5az9NY2TUv6LI1Weh1jM3EPZ1Nfbm65PEhsYUnM5+Y
/Lrmf/lmHiWrPOnegvV/6IHNwt+1hHzuYNdydDYhmmwXdIDqODWoruZb6FZX7Iym
I3TlF2WeNwtFqGG+t6DF4kqGPw4WIfwRDYIrx3nc56jnrmNRG5ie4MgvgymNyOoG
f7AfUSQSL3dZiTgct6vMdIfRylLsZoWL77+MOG627L66uZ0tNsXd9BXHGDIRz5vx
NJY2PuBjtpZlZ1UJSSXuwC1agNNxYJhhEpL9176tnf+dl70G46U5RA2XhBfOSRM4
vTC2JwTh76fnO2t6LqaLEOCHQXOrOao5SMfoAvlcRuv9sXIoVDKMjjoQ1voCoBhM
9T6V05Id7Xa7Q011Gd5WMTWukQhWatgCkZoHWUDDdIAvnxcoNXjRJzlJMLK+Qzt/
`protect END_PROTECTED
