`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxxxgQXSNQSmXqeKQJsEpNiyZrg9Wz6qeu41k4lXzHayU8XeiVT1XVDFSahHIL8W
PyH3nihqUFC+d0SknWgw2DZRVbk9xHY6XCr8GR4ZA6AlNhUvRJWqVboSW1LHgt5S
aeKUXCxH93eiH9s1KMBsVtCPIHCzUbJOZ0nQywLsI/g+N6D3p8llhHtKJ7L53m4Z
6vSyxz1uDwCLLDF/U/0CF36InAVhr+Oy3SMfX0QdJfbLAhOPMsgtPy7kTKL5lpVk
48uFLfySvIk7bT6fHR3BoebmVGwUv+nVLhD+PYJsjAm5iZpf4R8wtaCtuqFfyIB2
NVJnqKsHlpsZht8yyRiG95naIG8pEvn1seSM9jvCQlTPBVRVKjU0Jxy/2UAl6j1g
IVMnic4KX2vdgidLpZVB7v8RLPWRPjHMCBpQqNWWskAafW3tPBssSk3GdW2san/g
KAgRPGV2IeyWRrHbytkGngiuWbmMNxtDIqpzd5K/nZoujBq+m96eYMXeLzCJhD30
bQjl+So/ad/fGo7CM5dGTMNDH2hkBLuMqKKBEN1gzpfWhLc4pak1lh/GbMsdtG+u
AorqD25Rlu/B6zyF1jIci1zoc6kOCTxis4E5s7psSB3T7mhkVOJd33AfgPWmgrfc
MORfbRl+D/P+CxGZ6B8Z7pmEWj+cEab2E6WKq0WeJx/EmOy5/7OPCfANYKv91Zrp
WYWrtUmtZiM+xQQikAHubp7RcjqmdC4RBgpViaA1hCZNDw1TzmgnzSGE99sYvSbJ
q01WvX1bgJQL6miTfD8Zdz/YRVaRyCxcND2tmW4Iy+OS9kk3YblTh8BlEz6/1mBE
QO5UZdjI84qfwe3RaZTnDWnnCi9bJxvp28G7K1GeQzzTUClQk09m842DPFH1Qydb
PjuMuVvCL+KnG/RTvtidAI35kHp2YPGDFsUQRZ9+DOq2CYJKjIOEupLqXZ1J+GVL
FzmsqE4v3HUmEmQvBfamNutTyGHT/ztuQAA8Pp+cVi4+1gME7cdLw971f9J4a2Wd
TgRsS+Dsz7fIGrNtK/UF6Zb/YtDvwSG8sVT9MCWIVKgrcvvfYWkKSAioFVxW/eGv
nVtDeq87N4QlAx3RpxbpmgME34/RFj6I5ZBBRu5D70FlMiipW+vP0jls1KvEHe3x
gpV6rCMU306OAzoWNWoMu6eR9Ok1UEAH9n1YywNZbtP1MSGHE3WnC6JtwSvicC1n
dkS1k+2ZqubHN6ENDba0fdc7+OcrfHBIXZJZI37clN9xWNxdUC5x2UkDwVtXwf4q
+DYMox/KyBgC+24e/LzBbDS9Om+OgRuQwp72r0+cYC+7FV/QtyvO++kyzryBw2do
wzHTSEWyURQS5AmyvtpmEC3PI+oZep7fDmgIU8n0rVlPFY5hGA9xrRSoawP80wpr
0Fa8XJYi0t3dvuv4NU7Hv2sOIkbhDWXTw+XwMUmrA28mv/Ast5ak2ZsjO01OXTmD
TH2KdMhUkLdFZ8AJKOylOg==
`protect END_PROTECTED
