`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mfDtZ2tsE6n1p/BRKuRpxTwgRDgW4dUY+CCDK5qnbMdx190aJD86aJWL7/M/hfZS
wPlCPd626cGirh71A9V3uo2Nl5CIlcGLoHPlLuzvLbj0kFTQ+QY2o1WOi99HFkSL
jzH1JpQjLzVIB02CCP+DyXdM1z4gxTm3jJJAD8h5lT4JmaS4XpSt24vtoDWHQ4Te
4y0w1TacBbDcw7pHGoNE3FoLeFeuH6sHv2peyfH7NRCDfWv97JwDTYA7apWVgLvp
o+O8kseOgxi/4pbGY0IiKPd9u0aHmYesYhWojQ2nG+GwaWxQCGVN1lGWD1zbhSi8
AiMNazRCr1ngjsQMPTe8hkFtSXk26CMoQQxiVRQOCWFa7mctUJXSoQ1zgMhFceIU
Khm7H5rRwafnGvWh80+qkdVofCVvyvUFZYHzUllgQzlFRkFvU+wSwQpZa5GeNCOH
pXrnnFITaPBi1FFoH3vwrOTK5sOwyykcLWgIau7iPZs5pyzafAULWurchAG4c+/+
16ckNxt90LBU6bRTfe7eJ+GC1pUrRBX1uLfaA7G5Ebp8eaRnn4Nbhh4f0TU88HCr
AZ/1OOJNOVR/Yjf4bn2s7YD0efvitldSUUUvwF0IIP2aTMX0KueWo2akd0SiUzFV
ZugGJ00aWjMnJYE/cbGtxDl6mAvoq8T8i2Kd3UPTEufCZbC7ncIyRyaumKxzIIfY
ExGP7s3XAzZjBJnjB+/hGfWRm4ZnLDx9vkcc8iv4lpav+DVtWStmHmpzyoWlzknw
X9nT+Z73PgW9sHtn21JLoJYYRznnXY6guWYL8HyBRsmb5TpEJclRiZxs24fBguWk
YXgQoH8YN61KgtmQSSOkOgBbcvim1j6MNBQy4/aLTZlZixNFKGYGmZdW6+Nqhd4y
VVkne9kW907ekwIDf9IjDDkWCiK1T/67/ue+oZJwCySrrAiQkj6w3Evjj1UCI68E
UkvHO/TsuWW6LvIE2EheiRcjVfXGYNtJ79NMRtR39opbPNqQcK9UI6P7PDjgiJAp
2KgvjJ2BmNowRUg8Pc8wq8TaRelVEZQVAoavG5i12s1H92kul+51NXj2B5fdE+X7
`protect END_PROTECTED
