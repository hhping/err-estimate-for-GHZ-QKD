`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uPKHwzAWdK3EOmRXoIdu8HyP88a4ep6wb+Ja85/byV+E8fCB34HwefCKnhW0aVPl
FWKeaacI/rAi4p4nLxK/JqwS3SWcYlRN4DncQG8KA7F48F16tSREI08GFZGO65tV
NgYi0AVSDWCaTBMtKXhBheTq2AHO88htgxNfN5byOosV0D85EyDhLM0XV98yMfrX
i87aeTxtyppZ1vBr/buA/49qrzKUaBzIIzmHwuUWjPK1rXD5pywEKQQ0EliU7p4I
JhlPLHOUkUInrV7EUw9lAsOZIOdtrsdQYZs3VJ37OfGS7LufyrVBtgQpUdO4MbnV
82Ye37lIDMKuNJsukO6c1sB324/eRHYyY7mSZCSTgs1j7oRzQqW2rybOxlN7ceVa
oaqfFeOB8UcpV5dRu6r1yAF3mcNL7MvHhX69YiPV+Os=
`protect END_PROTECTED
