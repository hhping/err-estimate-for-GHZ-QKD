`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNVua5tBEAViPqYaoeLfT+m28uVl12BKRi2aFtuE30+esuseL92t9U2xA1umSMdU
3VxkfSwKPstP2+BvKKxfTizr3Zn61g6t+dznf6JLQxS51Umy4UUr+C46nt7DcUJD
AJ9iC7A7WbtXB5JM5zhhvjian+9WKknbgVhMrBTAa/H+FeU/4SE6w05ihWHPoOVg
4KEnOvMqxeC5TwSgDTTGd5Mro9dYGZea0Lwl90H9SNd5Q56y4HMIa8gm//jg5HKT
20UTAalbXjMkKmovBqfb0sCTqAPcCYOYEBSYkjVc5NP5JsexUOLi9TXRTVVE49Jg
wtzZH338DRR9LqmTIisv0UtaYkFHYej4rfdWia9TNjaEoSfgn6yGHrG25ByeIudX
IKvNGWuFDJvePDwv4/ySeu2CS/9SSJDH/oggTlsqWdO3yUlrRz0W38L6M8Z0Buvy
R4laltdTHu/wIXDyrXO0RfDYwzGO+Hc9ST0rnu/3YG2173upafVmmscrBLVal1pb
eEuH2Xxz1oQz8G92iotnaG7y2uHtFsdGaxhsxkn+YtydNV21CFIqmdKDIearKmUq
GCaTlYCUUdpmWtvjF+jXjlaVZ9t4zg5I5Gq+JZFh3PRo3KHqNijNkGmKbZ1SJ71Z
xfJp9ouBGtJwaxuq510CCkK1s19Q+kwIPqy/CU3xhyKEwBj4Mf23uZtNr/rvcHOd
eR5HpTMNhXCJR9l20JzMcy1mVgXN4hKHIlmnKBMGyH82OBTbh5h8m1r4Na+Py6oh
u0INcKLJItzPG1Uez3GRomv+HGSaHoz2wje9IwtEgVrU4Mb/BkG0832RUbjHpBTC
R9d1NkzoSvIisWkdvLTQVy8Jcs9JXuPqyP5oRQ5dP3gYOsUyTsC40grTKE65HDTy
mSp/M4SAIPRlB23GCjAiKwSADKK41Jn4JQhycI81eo24/C6WPmArV0QDoFP0di8T
BlAO5Nhxz4Mn9DY1IW7y4cYxoMeg+PLASTOYmYoCqyrJSRxLnCqpKQfT4FsgjJlY
tm2YS7ZVTLTvd6kBmmwNyCdEJAbRBPIkgtI8NsOUvofql7qMdGs6hzuKVNfb/Q5U
8Wwi6nhMAXiF+jWZ0sSNS+MYvUGcOtIk+0c2NtJ+fGEtG6ZxYUHDSzYgBvLKAtd8
CG7iKrLsthE5WGfFnpefhKWXpJEW+rK9sGVh1UQi3ccB/WZdAxwH3LkR3Z6lieSl
ZwV5ovKqtlP1JXnon+pCueA0UgUA5oMW/OAic5xhMzeJtMwNenrQFUTEn6mb4GWZ
D/SUqkL65K3TFTd9yYFx3W9QlguLdKENHxO/hTXQCxMUoPrMj+gCUgK8XeTvFf2Q
ypF8e+sb4ElwyuuYFV+gWturpKx6FzVqhT9+gqyuues7+iJmDbMKbRnR9P/dinYr
lxe4uqt722rMg2MCCTJ7eQxeTkrGQWR8XG2tTxi9j9w7a5VfNJycIJMhD1Mno3ob
eRbFH7p/75Wvnz+RKFQTrqW1FCXNXhbDU3cFID0KcgB3phLn6teMaEGyPL9ADRDc
o3g2YB3kDzl3uUGRYxqBwgTD0neQEfTeYxIY0keSRix4PsBwlBjNX0hsO8DwvmWD
u1mY1/MqBmnirTDDCyA9tm7VDjq2PZzHkw/zTp8M79NG1fRxUoo2IuLs7QpHIX5t
kvXQn9NF2EaFTS/q85bcEd3PbKk+wF6RxVsGbIu/pRyhNU0QKwvSgjwu1P2oOhTK
f/P6CHJioRd0iWDkIWTj4TGHjFOe+Qq4TSpo36dZNUY3Oll71XyIMvOematdgWPo
R+nCJMlJLOUfVqRda39L1ng/482LY/epJqjy6VH7TqaaWQb1L4QVk1Qolq1LSUlN
9jNmb6lb/OrVuSMSq/2vJ++jqgO8nHFu2htfnzhaklcazXkoTVW3vKrJdskYGSzD
eYi4dihOS/33FGjD+CA7V+XCK5HOfo3o2JJFdZa2xB3ec9R8+8MFgaQT0OTn2Osf
ulP0t/kKYMeNGaWEXH7pM2Mwg3OLs0NHCKyl4O5bHLEsmQqGpo43yhwN6R3eoYzF
62+PXgMDQyr6qOyVilmxswz0zoKIF0/IRwSJnqc1FbTNhiV+ElTXSksvg0rvgmKQ
zufJ7aeSiIG7UD6DlqzCVV6SvH1jNz1ZPyt/Rd+MIczmumxnHOgyweksNmSOC+Dh
w+HQTICwo8cLqYNO4YeMvfaXCFI+VNYyjbv3W75eYZgQKtfb/HLbXSLI79kiFgUq
+iE4qOC+LpPiWd7KqqN/i99778tbhd+JiLMobH07ljNpwW0O9PZccV360E6cnNBl
rDoNe/JvLck2SxzzmOPjyhj0/15jKAt48zRxcKVl8yfstPYpQHIMk6Do1T7S36li
eOG4zZIatsobKGUW3J+087DzOoO5LqpN13pKRwm7wg1CNT8lIUOH0PVBKm3A8lU4
ZNsqJyiNKRv4UKS3DwRFsdVHVA895DyMGODNnM5Y/3/YEWRpr4jpCoEoSEqkZZvw
XqJq/xmEjK0kfLEgKYwfmNpMmEkmQ7K822CO2H8tnfJxiR5zjqG4HQVuqf5yoTXT
zOJCN1gbaSm5BJ7sXUQ4AuguknKIQcUpws+juE4GdD5TwG/qqniVz7/W7Pf+qprz
zvcLnQeGsQVIqjK1+l2KtiSOIqkd63sgCSVU0wtt+J/XvG6D73ECkf+BM/6z1pFf
QzOnDB0lUI/HR3rRI/aqQylzvJproZycJf6NCYzO/FtEo3OfFHXOjuAg7M9sguce
4//kcZ55TTcbkItEWijAOPpJgI8VJaPiEc9mrYJu8hsteyNJTnWOBDTKa/+sap9P
qBJpyrDSjlFF3S17l1ijPG8j7VdPYQc1YAkPQkcah1hTXRLLce+p0XEnzWiKZwA1
hBXmZ4ZIggHfdPJNaQNQnKFIie+aTCj6QcZ3clJuog1ZyqYGdyPB54WMjkEeHwCe
dVswsiCASrgrdirSyUvFPiGn4XaYaHcrAx5C3sgut+3Mi/jyb8g5jt1BahfZHNi/
AJcTPHoOkMvxcbxeDXsxKAaBBbOMdKCI3+t8F+3QzqhsXkXoAEjpJ4SoIWixd+CC
NO6wE4yeGurq7AHb2Ws7lY2Xv7qIVZRYlCA980LTBON+QELrQQTOK7vMkwuO2y3n
2DaUt7pieEr7V6tJ1bT/HpbMKmlyI69PLUtuS4NmpiI9wrIWpQPahd0Vuok4FNLt
hzIgWsUpWaLpQxmgIrFS0g==
`protect END_PROTECTED
