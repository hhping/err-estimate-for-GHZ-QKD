`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wm3hu59YsEN8VcATcwpFFrQMAia+33GRSQHb8fHUYMHz6epkTFQLcesgSiNUf5xU
e6EDGs9shKolFcuJowisaDFwzXOWBZX6hSkEfjNSOyG7H7Vf9l0yzvJ5uAnCNAJE
kPAnNMTH7CUuRoK+3em+ujjkOof9Zd00fRT4oXzLhaVGdVnBE7WbIv4GxRDhDAWm
P/fPOflN9ClYe3FxRSFico4X1Tw7SmQ9DSH+fsOZ8vVgDcfogUzri93iCBzbAlcx
RVhhM99ZaFmS54HerY0tFk7lovZh413xA8dGJ5jg1Nw2Qd1QIXY/CGGsu+gnYkcl
cMKIbxO5hppjM/XGoJNe1f/CORUXZrVHrxdgF1uZ8tO5QV9LMpeVqpRbM9MXjwuO
oj14orYOGZH89FokI9N7eFk7KSek74/NN9DIZwBrZ1M0LpO3epqdjTAjpu0hk3ZM
5spowgrZxPw1SQl4znruoeK8SmkQ4rkuCvwUglQ01gU=
`protect END_PROTECTED
