`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOLA3g2arZTEnIX/+EJwjy0hAxCBVv7wsAxQxC/pmhQw9KtG5WNhewEiTKZvtPss
2LD+BfQSZ6vARtQd97sKMWx5fHIQdg+PH8Y4n3VyRwBWb8cFlBl52jlN6S/9M52J
4E+rTPLnfYaqZgCy5sremKchrkZ5IJOrHLgN81w2VqYHe4lzoRQ9fCMyLkcqF4ZQ
lR6/hMDvwTizpT9zqiDgJo5aBc3gBIZRKnnT5raOiby4ynErRBXMYwGJaPf7df3G
xXqifNuJoNzHO7U+HaSLmDpq3sseBtEbC2nWmPmwEdihqdyqw3wSTJDz1hdUgadq
s+Rk83amb2Lt6R2Z8sfUa+lKOHShWS3xQeDU2KBmThp7nRJlU4+HEwNmk74fjvTw
fQcDa+ii5a3UI5g1fpRoMRPxefp1UzJdwoTMrcd26b/uUIK63p9kSq8bUU91NO16
FY3vBBdSA5akPG+hhsY1Jx5XuQXHVwVyo+utLHhIUSgcrEOvY5FH8wXQWuqUoAuN
3cbY4TdxLFrAk5/Tv5u+UXjV1sD1YsYyPWImmqPyfcOWDxm04sx5O0FOxvbvpeV2
Gw6I/LFJT50gQjvsVCBcTTCvtKSmuclwvgn4pUjIUfJwOK16VeC2ql4T4Kk4xaUF
0GhFyJAhprA5kHdZSJCALsJ5xpVT0p39aHVU6/ATQEtHyv5Ybz5Uj5jUdIUrbouN
xz6vP51lEj8hRV4S8RDJvu/7rR9DqK8crF8UkURrChPXrPGpdIqFNn9Ke72Ojl+u
5EK06hVYlzVQqRglYadICbf3DplesmAJLN2RGl/32qs73ElssgLUuGBjqVqIQ3JL
IgUV4yqE6+lv6E3NrwkX1g2hoYOwd5X6J0YUY13wjs5m4U0uAbYhiWPoBF+iE1Hj
5fbHPUVHuBB5iSzGqqu0gNoqnuz2Cvp7GNzgkSxp33SGGBnuyOpKq98jGN9ShjYA
UK0QS3OXQjROqGqsGftj7JR281j/S5ZAJW0/O+k91B/fQZ+8TUv9Lsn/68knSb2e
1UTqV5tOmG5pymUmTNFkVQK3xA3v5M8hCRjOSni05X22ZeohuDaWIuA7iMZlDJHa
b5y6Rls5pYuAQBNxm9AX9N+iUYApHGlXWuX0mHlkvEWOY8mfQbs+inD37fziOMjz
OxSzykAY04wiHLLgox4cJmliWQYRRmasqgC6eFiSeN5SaTNABdo9kNX1lfXaGFll
Qg3EqeGDi80nhCtLSoLOd1SqrW9pHUeKpZQ/dWvk0FoT1fhzWUVPvhO7TwyfEtUD
KOL8RSfOfqGDdJVIIQICIeCZjdh5Tvo7BbhQaA6ADJU=
`protect END_PROTECTED
