`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4sYtVnSPANYJvpSvjnYo94N6hcgH+wOpCKqdnVzo2tENm+gLJ4saW1ke4xjs9VX
dfMi5/w0E1sWgdXgydoEAdrmUeGvIP+KCM75Gdfq0gH7BphfKV/Dia3XZ6l5xoli
QfZ1b9Y13tHyJRuWPN1Qh72KPvx4da2oGIqgeB5R5So7DhLm++T+m6qoyEOrQzB0
UJ0LvURqwbSYXMnZH3isEGbiZk50vi6yecefj5ttoAS/vxP5eitZeOoMQkjvKrJf
vbIctt6+FXTR0nw44/+IPKpZJwh/o3ZIbs8XLzKE7uYAxuLIqlad5Wew1pFb7N57
cp+Rmb2+EW6nlvqktmHcC7ba4Sni4pvUnkinzUQ2WrVuu+kaC0iyWuVujqFQkSOD
Hw0OiWY9YFd0M9DOzrjD5UW8/t633804jyrHuRoJGCUrznu7fD0eoQAiFidr0HFA
Selu0/gmxCDogcNK6s2iUSq8kYF3uheWOhzaRKdv27iWSuY7YbNSE5EPEPEllTou
WKmJjhwEJXAI541ufTozrSYzElIU6ng6tMH0QlbAB/rx3/onGj5WvbIzIU/DXWOj
XFFxbcpPlmo8y9zmdfrwehI1U5RNjnwMja4VmBWrx2xvAdyBDqvMyIoXqgb6ETIr
CZ+qNYzyfIk8sF8bbfdRjooayRgi2YAFxfDhmVbkoobPenhWEd943t/ZQ1TlEyyg
UpKmHQcSgYP894RKvYmcZBmH97Ityi8FmkjUNBothyiTllydaFNdM8enNPMK4xtj
hgxgdWOUO5AYL679esZJ/C5OMM2LE+67DrN1fPe7xP2J7sg2H2b295aYr44QhsNC
gqrJ9msLKaN0NESPttEX4vv0pjIMMRrSDeI6FBzeK2WHicfpS7ynlqiSXM9zlV/X
klxrFOeEAxzF/J8xb9uOTvC1UznIhLJQv1GuDFKCHScYC+JFdTIiEEzK0fvdvHlQ
Hz4oVd8yDcU1zB1yfRiT4m48p+aprU8uklwvR/MDNVRLFXCayOZ5sMhh9Sp/zGas
bM+pkz0lNeDpXbXNIpF8/QDVyrVYTKjAK9jGeVrT5PabTyD5hbSnI6P3g8UxDOTH
Rt8nQi55AbxhX4wD4nIoGPeG9QWNWoy/HfYcTHMwVV/wCIK4zgZ6covzdb81L9wu
Fto++uZnvd6llVlT+7pNltl0jZ8FWOuvTyXG9fGpseR6cVV5gZlIZs8jSKu8l70D
1ZH51Czbm4vjpaj+F5kyNB/nyeyF1019kio5Wk/DWDcfmn+dkyXoJxW5yDy9yDbw
gEctZkR6gbxI9DLpJaRbXNRRpgoCXW2jhtLkLECM/KXSQ+SLMcSD8LPMBpgdfghF
gR00iySyaLD4Nqy1jUPw5Gy5A4roK3svLevjk4Jffs/DTq0eSppa/wZ9IWr1+fAd
lcQRPDv592DGsgsCUnHeqco52zq43rPTv2gEXCWCS3PFnLvFQBAQwmrFhjqAV/0h
RzBiTTGWVeq1Z28L4eV1PFC4eo5H8Mfyq6Dw3v/V0MTqEMiPSL2HW7kbl2Svr7vC
4e6Q1XAIMJkNjpKhJn5SfOH6eXv3KuGQhmQU7O6TpHhuqTX7HMW8mc1Ewk8H47n1
/jeKt+tT759sMugsyv4s8lkxZv7rBRsBGP4Hmvu5Xpe6F4QLGbB9O2In9X6PORBw
Zq6Hx1D4Ps5jRIOCsSfN+k1P1lG/zreGGpQaXDcMgwaXfaAuXFEXZ3KeZJLVMrQG
/sfu8p4P4pGPs1mYx+DULDtdHBUbpFGiTdzrxyyfNErZtgg03ANGcWwJib4cSpnA
fOEPBmn05U1rp5yW2LjKHD8flDOfLNXP060nfDyHn6YJ3B5TqJYKAiofgNt3jAtn
WENxNGOFJZFHOmXkFcVET789kxCUf6VfErga3NAh+DywO5yLlCAgWDRBE7j0rG0Z
CFT8REec95UdW+oU3xDdrreq7SLvmHRoIome5Eh8iBHuWjrWSmcsyrplTNmjTcsX
CKVPNimJL7jrLtX+4BE4SKTyLqKAtsGz5yVLLOki1E9Z7poE6JNe1m7SYkD7cF4P
ilma6AL+ds5YZc0MgESj8GMQ0PKW0DGedW7waW6NJCBU1Lugv9RrQ9Xt4UEBMe9J
uRYXirFWzbWhKCiiMAQEcE54V8CLvd+CY4bNiIGAVrZhLGamPI7iiy1i89SHE97h
7w+YbeT6SQmt/qqkBVNvOHU8B452zRX0L4HI/52T8s0bXth4helRXv3NEYecpOMN
YXYEGs4u+vrS/MDsZque9MInJLv5Fkpx9D+vAVn88Ncof+6WHYJCrcK/ym3Qd/0r
yMr+vHfEq40NW1R3kF0D1N1B9UWPCf/ZeYnLbW0MlukeNhnKDD6DGqXatsFo1nT8
NlQMKVe6aRIbytC5FHk3tN3QkMCBo3FIeKBy/VgLLcG9FD9Vn4N0Z7rQIfyHpL3h
LTsJoCvj2zN/5WKnYV6RWR+W/A6fGHLqZ5X2Du1N2lewXAY+H+udNzpiUfN0vlDr
Oj5NOdILzQnsxoXbxw4WbcfiDeQfjj5apP/QVPb7Vm4b+dELCTjYwcZJJi8azInm
EWGJ3nHxiPZBIbWajSFM82K32FmamOeIcsp5uwa91Ecan9qkwWd3XzDMb6AZpcMe
+dea3AfLpbd2Wq4TNIX/En8RO+WsOUUVQGLk7c0lxQ54j6WUQyNGD+dFGrg3TjPI
1v2LTJAW7L+uas4XzD6j3rCjSjmFoUJ4blA4ogrF3RA5Kef5Is/DyR1GLm3LC++T
9AJ1QQ9i2Klmt3F2XS0tUH6rk/AbyM57duSvAVaXpY0bTM7KBbCgjCBMstW4KJrY
UjQMjKbHr2YMAibN8BBbp9TG4EkffXfzE52nQUG22kIkMDFJeRAr2JepYEUDBjMA
0XdeBstd/5z+WF+5S7ye22OR5hlJJIWw21Q3m/TGxc0=
`protect END_PROTECTED
