`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ar9oqTNAvmdLAE8TZv9RVwJSk/Xd32o52SPFESmlqtZzcWaUnoJ8tVX1j9TQ0uOh
oH8aVUZsZKFjjjj7nbLduQX6hdPovW7CmYsk7F+bl30u6DtmMCendNji43zc6Moa
IPcdOtHfkKdpPDmb6uPOVYNMcGA/PWHjhITNud/Rq1LNLwGsQvXKLes7ecO6nqnx
LeDRoaVAvRbvqQDtx3doTG8/aotnJKTKfa1oOf/h1IAMOpNTsgfHEB5CiqrbQeMQ
4981S7/lZuEkyFKtxEXpJImS75U5V7nj6vu59KpMo0OH3GRYFyLJ/AWpSYYPVqaK
djWbqgxTT0y5/+2spnZdualrsvTjXDtAeVWT2GouYAfAZYGZJ1HB8k1HIeJcAGjq
dJV3gimLnp98yWPNINF8BF/+i6ISMWr/WUC87fKMMaLaKpudpkgLKaqFdGRfl6z0
+Xy626rAZvPeTe6lpeWx9Ryze5ul/5BDX3DMTGZpGW4M8h4OA1J/Gm5f1azDTGgL
xDTyJZHbiIFKs5kBsVvx7TUM9SHRJGC3tgyf24kG8OTOakAGEeOJRh4YIO2C6vC3
afkUnDlbY0GUgjHfEqSeJKzCi331lo+0nCnihfWIA/RtJ22PBmtgRV6x0pEPBtol
cti2Gw1zSlxm93jdAbmQ+gPMLzLh7Hr5s6y10SdOYdVE45hjUUbABBymB1tqltnM
`protect END_PROTECTED
