`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2qr0q11gI7aZZDnH8vULrBxvOCVX4fftGwh10tLV1HAPhFwnX4EuX/p81iRdKSp
uLydd4e4HyhuJaOWve1jgK4fKBkIH4rhPl8dZ74apAcXfk2Rb7yOITir9uw55bCd
Byvpx3u3uGjSEaVEqCYnI+qiYoQCrsjhGa4+nQya07a7jz/8Ns2UoCyrBZ9PqTIk
4Tc7VLCNoR+GAdvUpN+oYkFneyBbIYuZDm4fGDwO/WpVfIsCC2Aq4QpLkX0jKScv
Ha7RMJfGyr32QSPqh3shfv6bI0NbybtzkZCWUdLblGb1c/dzlLcVpdheExo/gnTu
bALw2lBwdlakiIX5dsZpaXeqZOJZG7T6zyAvIZ6+utbtTTmCAFRMTx5Y0U1otpvv
xryuegqtiGhaDj4WS6SJLuY8CcNuFBdVKg2xTy32UGcU/NMikiz/YkfLbTD4ixhJ
OlkyxM79lNJZvYpUg+7GfTMxpngQ9xHv2nFr2geB5splHTVnHzgbhR7fylG2gx9m
N12bbz6+bwmUy9SjDMtNSZE16tLdKU7Ai4T1mkB85F19EkIWcbsttrTm5mJrx6EK
Tdbwjj56B/uvr/+nf8vVL3gEX01uGELbkHnCv4ZN2xi2DxX86Ke+P+6XuXJInXd2
4/+cf2jOIE0J20yQCel5cNlyRRcwTgUEERNx4JkqXxubMCqqZMpCwtIdCzrAJbYr
tgBLocb7pMmxnlW845XKoY8YOGBNCqakECf5DL0fOmmFQGG55DMOBg4XgsZnTei4
S/xzMzlrDZgPm/TevQ5YpsECQlYCton9su+KgNZ+alDe8BPHhqTDhgX64rVqYQCR
4/FkrybBPMbAKXvTXBRMiuzi3IsdFBq3jyfft1w9YNn9iuv9Z8FIU13HMKi5nfZW
LSHc9qJrqxAFPE30z6pna+sY4trR9zmpMX1Sgekb/zwdbRkqLRnMA5g26xkbYpPd
do0LdrD9BUucPUmJMWt8JCmgte4J7Q0KgBL3mzC8mfMFB3nPjFYb1gHcfOuJf+ju
lqFb8Ak7smqxJMn5jTUCunzcFzZj+AxkHfwh2/k1/N8Fyn8YBaUsjL4L0UKcUMZr
FJEkgWvLglk31chB/YT6ivFvrRUHSTPF56q9mFANXj8+VEiXzJd+2SacHmav/mMW
Eq7XS9dfEUywK4J+mRiZWN5fMOy362kNmezp68+IBD1X2RuQNOoUPFivI9BZL4Ij
Eey9h7T5nPpmmh01Ysi4vKcfE0rl3buNdds1IEUdAk30irXiC2WG96RG4OLWov5Q
lmvQLIkwKoJ79v1O9fYLcAt72Q+uNLsZX3STy7ztfFLZMcSgD1XR4S9nrx7sR804
zNkg4+oKWuEz2ohQNVvQYIperqzssO/uT3p70w4jgoJc7ycC2zGCPDeXZtzKHon/
JBgUNCHG08FmewdrE0lAWZ+2paBHPBh/9Y/V1VgpeD33pgAoovS8eUheMIG2Y4U5
La5XNU2dBz3yQG+o211vz1QSo2wrsiH7JVM0Bdxxy7sAsKhP1x8qngsfDr/SuueB
jvY3uW5IqWszUIFs7fC0jsCEqwo5ITd6Vk/xagQzjgsB/E9L3GSusOePtYaHLElA
lwwUrNyY0aBEyaY99o90uTCobZeNiSdclPI6XTGelZ8R8ofwUwzjPhB46ePWMw3B
wKCQY/mGw/6GbrvFoLyBUihkQ38hCJhdapcLpGjzbwwtf88LkEarZZENYlktHQCc
dW5f8zusX1p7E2h7gLRRoPwub2UFGtK8Q1RRZPRDYlW88Dc0srjhwMP0Bh2uo99F
1BS3u5NTOgew18S+I1NEM02cMoc5FpOYekdFONP2IPEY0gptYOPA0oL+SDe+7b4v
E50Cq1bF9wJ8sjB0T74sJgB6GbwRsVinC6Nk0VjRu4nUkuhQ2t2G/AzdqIBT7rYP
dAyvWe5TzV3RXnkud60xkhSNKFOvnc8/a8GCVffouFhCrZfbOL6CGiMyotqnW1WX
gZxPeKVWfaV0o0HjqCF9Y5mGTEgXbcFoIfB3sff/ZVj2jRji85Z1IsFuMYfU29jx
fkX7Up6B+7ndul1q17uHCdWfM/WknGZHbNDt8LkISPH3WFllZURX5FgKQ3QibiAP
HcXj+rCBo/yJlOZY6EG/ylA9XActYirbks+nXiNiG39BEsiX6l0ZFEMV7+CzA5ck
joUCRe55FCtgf/9sZwRvwwGawB+VkKnwt0+1HdfIwYs/qtTdpQkXjV3U9ZqL5EwE
aMZl3zhKjbGghivZxpq2eJQF87GpjAHQyC3y6+kbJO7Y+aw/BeBLo3ofJSiVSpL/
BgyjOFs/HV6YfCEgG/WVWvy//0UtMFG1jpbWo2yqOLxY33ewTExmcSZ7l/vRelw4
vkETyjK71A/KMcVIymgSXtxoTCxeTI8cC0ml9HpmiiG+u4vUYhqFAZBhEDZsOusA
VRbtHdpvfzl/y8GC++avgoLzPg/nPkQte2hU0GN422egAIBmnZTsCp78gykuqKRb
p1VJt9HgdeAhFksMlVSROMZ6rvB+RBU1zqouFlOwG7mxZi8Ma1ZYdh1oL+uWRv8N
p8WHOvTzanuUiAXg/cW8PGL8WM66Vp5zGVsuKm4HAYxwK0aJhSJY9ni1+vbo5/tR
stuWe5wed2/1+Qiow/RU4qe6Ek/qWIIqGxStljz0Opb7/CEdtlp7hYZDYQHXGsa6
Q3cq5z/JAPye9OiaF3Zn7IG+k3UHZ2YLEMSOjTuYlZg69VxxnMbq0kY8J4mY2EZM
LV5gwhMrLR0+SyKkpX1sm3bfbVkqCy+UuulCkLfLdmtjpYCEvh3y8MoC3F8lEGcX
ld2Z0u88fS1TEioGEES5oywlTKIqTG8gI/GzlYhArmPD00qkiqQWH+7A1Q+I2Hgl
2z56snxrhpP0tKfDSWI5MZYGMcAQv23ckyPmDUn5wFdryDBM2S5m5x0ReT9iPKOA
BELUBuH30QYZ3owF6PiIRja7MkhRV+V+FwnzBtA52Txir2cAd+NcNDAQtwHlUVEq
nPdMyt07Yb9kWRIM+O3Zd9UbzYOdGdwKtzGDrtg4J0UkKFxX7i5IaprxyWGinEF7
IWhwn7vk6l8H0Er3j7s7ykgDU1MB1okXGTLFEDe/QHoEGbyQb/qIUlLzd7v1Cwq8
xk+Vim+0awrI+fxpnEa8A6gvY/7wevJD5mDlmB4e096XvwHkCkU6+L8eJWS38WAN
+XMuvRbe+V12LmQCK2h3Y4LSygfSjEJ1l9vdiNt2AD8hagOEAPR0Domq1iFpT8lP
erTrxN+PRw13bKFVLKYBaQlIRBzgOzt/zIAgMH+MpiPm/ulri8+saqNI9a6r/+Iq
tmPBtrxAKr5MV4gz9H/r4FEcHhcWpYCc79fXoVguTQb9yzJiDAhABVMH1GjZiKQp
deFs+3orj9cSX9nMbrIV1coWuM8hpfFeQwFmeVctWsvJ+/37g6za7jB8YtXUQhtv
X6Nn2ejGlzA2tBFJbOSk5WJ7LJyOTi59kRpbIa4RZQUf43lujBDiVYGIhL616I+c
lDefNwZuYMAmtvi7aTfLZA5mTp0BZolF5LoiMRw8lyheWjCcmvkQWqUUZ+NyzNH2
ExRdaNiwdBH8nG6HQm6t2CwBxev7E4MwlC02Gw9dqFbuCkEwnkPLmkdgXNEYmujV
/1dZSQF2NFQl0daA+vvZX4jnNd7nq9f4HlxgIQq9cGJxcmhUXNmiSoAk7sYIULMJ
0WLgIuFPNjjIkY2ghU6SH44xx5yqaNfReuOw+XqMGP2aV/Mrwn+KSbf9cPP0C7Vg
IDXftJNYWECy0QqRg7IR9cPXXf0ddgIxGkmmBBIbgUy6jGnyCpMCjB0gHlkPrXvE
ZMkCkzJR10bEM4Lr0+rHiztRzhRMmDLavUYgTgfoqItHNYKshEGGCQkJlxDSsIwh
uXMhpwqcs3c/3+aWfedao6iNT63Hj5DwswLLW9G/ieZ9Hmd654/qUfGfHC/auCjq
mmelJFq2YnzyVTXlJc6PniHAfXa70Gvf6jlJR1dN2UycAg3xIKke/VkM9Xq91u56
zJQyxINKnbf8YOoaReIQTIPwojiLHAO43UM9AWwQWAbNET2NTEm66rfk+VZ2cCro
F71npNkJiL3nWf9FSkI00J9EMnhaJ8SOrLR+ni5M4zJIttrZ1/s5q996bX/M6gQg
/4fTAgRQnTXjl/obKaVctLZFpbXchduWw6R01/tH211yZJnc+t6SXIDOSwzJDI4v
`protect END_PROTECTED
