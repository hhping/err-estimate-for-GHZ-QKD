`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yttEQDlQ+q4w1JQMBjhjw7Rs0p/uAkWuhuLrH61XJtZVFjCLPuFFx/1u2o2lzO5
VH+hVCALK4joGRdmkGyvNBRc5RkgI8ZXnC7fkwfpjltu58aIJlJ2YHN7f2QYY+VQ
LkT70Q0AKvzsUQnB0SMvRkchlQJGvLM9xDPmMEjmAivT8dZucVHHGm1iY9Pks/dp
lSj8Qb/GkG7Ic/tiuNrfFsT6lRCYuzZueNbMKe884ekvLedUljHshr9Gs9haDq0h
R/cc+dZN4SG+PUhfCq0WeZug03AKXkeZ1FhW8xBBZFazsbAjwlgWdDCmVUfG5m4g
pZR9HYMYkxDKt+LuWOQBxTavzu1OJ2z5kS/dhz0zW2DE6Su7I72o1EojdB45VVDC
7MfLkpqpKh+8M+z/31iQtFyCt6V++rowKEft3d70/fWuzVHhjjSqpGEiOWv29oh5
cKVNbAWva32ku1kqn7XDymiYEEVI7xqXrrfkmyGqqrUoOokIAR8/8v9s6eMnVJFZ
/Id7JXhhectAPKvrqpEMdAXwmXrnwMXlKaZ4OHuV3Cqjjc2Fg7FaadOgIT1L+3LI
DsF+aRqYbaOmCBzgdlMmnKrM3F2P4neczpp7kfNA1hkLLGO6++H6RMuuWgqQ/yDH
FrdmGA12YpESBCMxvLDIlmYC2DlYyFthMNoENKU47vo8XGViqvuIsPUGAQquAuxu
Ud1fANjirpqW3qUIuJqGQjp8TEoSYmE1WrYk9rgQt1tf2NMu4mfWnmztodH3PgqQ
/QoA1wJJKoxC4VNxTwEWymXo7knfHpNz4THK1UdyEifx1W09UxQ7HfXq50nLwjgA
aLem0pFmWQL/N5ptd9dJRjCTPkIUu0H/rYkqNGfG5d2npcrqh8YqGd1xMB9CJxzJ
MLFY9vVj9h0CAfb8rUVW8AYwPv5yYq9U86vPqF/IjeUvIwJHhm/Ftaoo6392xjeF
GEFlSP9yR7D/DkEIN/Kzl4f/MnUG3tr9hScK6Lg6dzlqRZtsx09XQ4jdTwA7ipA5
7mE+fHv2ia6nIG8GTRWZ3nq5Jk/MLYG7twctNhJfjvE5WeKFBIfAszIUJpYBOwbO
Tpl/ldUAyEfdXdWcGvt+qADYea3mP73yhZpEvGW9Zd5ENbAlycTfbR/lM8cEZwZU
OpdC0Zwu/Xx0EsuCCcH+kUCnw9WJLzgfs6TJJMqT3fmO9LL19bjpDTLZHB0dh/T2
DgU2/D+OBfxa/f9Zyu+N7Q==
`protect END_PROTECTED
