`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AXIPzLVaqdFUVrh4M4iNSslbtcYH4dYO0O7Dt16ko8ZoQaaZAk7ApgAJlteWg5C9
tGDSpjYpmNoJpHrJzE8u0b+5gMZWg1NxM0THorDwclPI/XWXbmJHmLTYO2RNLG+7
CSQKIeq84wGNtWgRTy/60Ie2P0oG8U6HcqYG/xNrhS7l6vNtPtk1Wf+8ULFfjx6I
CKAH+MyZN9LJdqUVceBReaOdy8KknqO4kWKbVSdoxyt04TaVsvHdya1hvSLk3sJU
rRYIpFkRrHgo3A5Fm6KHmkBDmqBQtnw4/AHT0AVOEKSmVOOq/yIJPVYZbKgal7pu
As88MJ8vuLug9AMZBkA9yk0lbzXgdOayUlw1wvx11TelqMP8OTEF47ZIdxG9E4hc
HwdSR3K6QavjzaxzehaDPkZ/npjdC4AsqPEyOWgs1w4iQDzqSJypX5YVlmhrzSNr
FKE4W6jJvaW9yG0tBr31R0BChhZbXAOw38dSH3DQ6GXK/0akDPl7yi6pqoAUHI4R
`protect END_PROTECTED
