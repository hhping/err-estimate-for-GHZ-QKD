`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lhqzyF+CHPmuiVy4BbLZ86KssDLRJHUkxf3lLinhFEeSOxNHvuic+gRpUTPh6Wy
AqAUkqYl7FSbCNBuPl00g7KgIp+pBQLgo+d8yuzAtcsnZHvNDJZflk30MsTpkNB2
2l+J/t0XavGWTQzACCxYdLxoySrvgnelhnzYUzDaKFeuSBhJGnRKkV9FBhB0LzWw
yI0QBgsoKTMFXe4spFVUo87OMmlSrYm6QdexAckZimC2SwGPcfcgC2FwVg9VxF9m
qCSl7ZX9yBYGuo+YGjCV34tUhkTQivIL3TAeQyEf7kCYiDqq16Wa1OzhApnWfxe2
p8JfyeQ+LIcHWRE0rQWad6bCbJo+XYd5FV8XCTg2L+fFdoYqhI/oqaXmXczU+oup
O+miI0WGfyWq0APJQbyvUnMgH79Hv9nClUkw0SE3JStnsqx0OFa63euA8P1k/fG3
3TTvhMzhCWPVyCk6v0+dRNfOwL25PPM8dpTsApLvcPH4doihOWCpkiYKPj2Ar3Gu
l2yAU66ubZ7t64tkGjfJ49qtloq4ihEbLG5ze/K8FJuxrWvxmCBc8VRjXu9yrAdz
DJzGvhT3aFG3OZFwxixgeXdiZ6V+PSRCUuRQOPj0cgPrWH6KWpZSIRGLHfKhPvZI
BYZzjUUYFWh87Hmgp8S4ykJJGstcd5p9IjWNlSi72Mo20O4t+0dmiOqbb5HhPhGf
+tegLHB7qWyC78eOnd2OCz7BZVwgYIr541CJ/neBGi8CzOA4pgac6g4/hTqawmVv
552gxSau9UU93zJq+aF/KS5gQZ2RWDYDTHjnz/8cznmdLU7aJGp7X0RY8hQrNnX1
/vUWKlAuXYB+Ogj/TmcyT+ytricdoRDsoKKFPIXMjxXadXS8kf1dnFBbE4XeOQ9/
bgfyPRWi0umUDtLjyMLzG2HlLBUFIvgYMig0+EiieDIJnw0oclRi2KPYmqwMjlj5
EuOMjmdsG3JeGF43w9u8rV8bkCxophLnvftfh1wdN0aYQbUQeOSyQGhHHeiMZCEN
y1kUI3GRt4xY4J3xlJpQrIqjTJiX8HNsdkM+LWOZD2N6Cqt2q0BCDuqT3YzaYse+
uQ3dQD1I7y5PSwnRp8DwFVCbVCWXznJDNtLppfkdamCvP9BwKj72WrSaEcIaLo+n
zKaWzMO23bDpWisuJccZxfBv6tqwJjVKMR7FgRDVVe1TFDkenasi4YAC1af74B3Z
nj+eP7JblAaTcibs2hP60+HCFYVbmEq0EbRk+hk2Eaq1B+29Pj6Q77IoTpevPDVj
C5BpSapXrEQHy8kk0cWD4gHZG8OTxNTk2dzKJQ+Ly8lkQfmT0MMvvmOS/3Xbvg+t
HlMNNmSNuyaW58FKNcjl/4h+LJg12xGm3RJeE2HR4j5OQNWbA5G7vCT5b2cMhagy
pj4ShoB246WSwATttE7TGmdpnp32KOqK5dqIwnsSo4C42r9puFbHgGsbmCK8kZh2
`protect END_PROTECTED
