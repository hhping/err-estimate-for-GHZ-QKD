`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7nVhYII84uVqplC2Gxab8IpnWc6kxVHaPLF56g1j7YVNe7Lqd8Qni3A5s8dSUwo
hE92AhHHBh0k456Ylv8uNcOZxuon/MmdU3YLpDxvr4Rm97tK6YvA9ot2kfB+QbAC
8DK5G0bxHJBGCmsFsAO75dDIrt0rYBi2uhbZbMSAnpkM2Wp7yEJr6Fkzz8BaXxSF
woZvguYGBNsuipOBKx8LJoD934uenBOMNdLgMuK5i6ztLRJzSiXyMRyi9yE7N6ah
h5OOS/U/PnRWfGO/+EGRdDQM0T/I9EaamuhqeEDp54gjxdn2V1SdkRSGoubfE89I
zh5AdPBSZMDOYJWfgvU9hlxWoM7rcuLZxwvnN8oGAZTngpn3UblRregz37Hfo4Ti
+uHHlT1aViEsio2rd2BTcDciW04R8ECrypENH7JoksaFF/gF8OWhmYUdXnP6YwHo
viwsAtfUmPRE4ALFN4W35t6bFIz5zXb2qkGuUL2ggCjgt5byZMmheTM3yfDkH7LU
IoXKjN+pHabUpxtU0DZFPUPgvdgngaxtexy8zYeT7fsUcgeWPMZba7symMwoVHQX
Zx0Y0J4NI4Ohq83jwIPJy/Z6FYQOAvqR8l3crdrWcoNV7O/3msabgB6b/pLvDD/i
NL3J09bGPNHwd8hTwTXal4L1OdOhmC4SJDttNapIq1eRdeo42vzl3snUq/BM0JVC
bi6wlkKTFbrtPwIntEseg1xkrgyIl2e2V5xpf0CQAj0=
`protect END_PROTECTED
