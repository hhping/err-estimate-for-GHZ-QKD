`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxSi9eFsfFxA/8WNdNf9uDNtjfwc1tmKg9p4ckb6EnZW4dUj0r0kWF4tw7ABbFyI
My0zDTFMH+P9mE8auxJDKrTV+taiFHXyBdL2QLrY0gXaOmA5WFKBdZto5HNEUWmc
8rfugJsNVekVQDIxZgpu3MT7PuOAO8n/to44nKM9IQLaQafKkJCFrLP2NNERodRR
cVlZEV3e2GP1TLaRt3+hjddwsLK93mjXH4t3TCxzfPKX6An2VGvA7QFtxu6lDfOv
XXRif8Hhjhmwfbf9qdaERiVyWAxGSnVvNef756Y0IjXZvoQRDsO8hABJg4DN3Lzm
9Y7HAEA24zzs1Et5OfjlJsu54ZZTYcM9be7x748HT33Bym8Z39yxDoiWAtsIDY9/
iwZCCxfR9DNBcPFWts51Cohv+mydxfWecGBCIOQWORMa6YdZY/fbnhp5yklJhqCV
1aTqQOOWKsRl8stEvClMu7IpSt2MYUcsSuEWukdxFxr/LepF6VjT6rrkSwXRfgsx
O2XQeEVwmrsA4+F8qgtCOp/9EvacrBULZOS78h+beJjVdHpsHkOauDgKZzv/3Jb8
MS9MGGBuZGOGFSd3u8FvxqLxjIHB0ObAUeCGXLSMJ5Pzac2VO2obbC1wOTybu8q/
zSD6VbviTn50YJAtfDj0Yjll0eOi1UAiWOUoqVvQVoyWQuqZJigTL61rLpg4V2m6
kcfblkuz+aQwDCTkuPeagOiZqXS1+rwyfXZBkVVCiEIUfmyDgXdNcQxgw4uJZJf3
WXRjXkm8X/bURHREgP50eA2Mofp1pS/qc9BSTmMMB8s6ML3TVK+j2r1EXLipAlUt
9sP7qdAlcuCRniMeMQZlsb3ZrqFZn+lcz01mx0Cv0Zzv4Km8h9Y18kSv+KjFlpu1
5mAH8NDu1upy6FtjZXaTwT4AZG/U4kLRzjkzlybaLqELfvnM+N9GNQsJsrSJg2YZ
8Uk6lQueawUg3GVWj2w4pimBqOnS0Buwbrn64dWAA+fBvmfGCNAuFmHuyk4g5Imq
ClPsTWQJzuJlzMDlpR9XZrZ1yLUfVODG9iTHj4SDCilwyx0P/Bz1fv43jW05VY2Q
oDqCH8k3Rl2Wu+hFMPwgR6vXxeJodNGPrxT7rDZ9tIf1jXLK/VN0IMfjegQ+TX5v
kd+7jGXNY4giXqHijUrZK4NnhgBN1QjEMdT99NcnKi9BKw6abVMkyRncDm+r6HwW
SSeA07VqOZQvQo3gaXoI7F9/jfLtZDrPMAdJiyVy1qZy7bPQji/YCyHXquq8ZVwv
PX+Z/5KnK8Pv0guwZE6A4cwY2dW+/bMqphFRewQ7CpUItRAxZfOpvAr1z9UMLgq+
gfkW0/sjp+QsYPAWb4TBKm+Gju3JerhN8dd7UTAVUcJjTSGQvW4cCuZNjxYvxMSx
ilazuWNiLEpZbBdsSlCpt95Rdp2KCgPo5cxcmlJ0qKCJRDq1Tm1pti098aRcvyqG
BYEDDGYP+wE75VT0wpzT8o1s7ZivwDsWp3qdSYv1GXUvqEe6d8z2ojyPclSTTVff
VYCgBzuIsi8nsFDKhjpmRyyFrAe3BxifySOwQv27xFmeZ5ZuYWO49s0OrWqDCQAp
kW57KJR0wl8f1acOZNiHCci3mbNDh1viWCvDpjnPJ7ijPe7ap99l8egbgp2afA4p
DwYD2LSkEWtqL8pOfw5xpiMz5rRb2JbHm+fPYqL7Q9u+V10XvHc+T2+h7E4m3xqm
h9pI2ruzQmIRbaDqq5eJVY+P3fS1yKrZ8er7PMF5UDpGf2iXGCelc58nV6csNiYR
Ydhrwv8ypHOvGlQx4AL4u7S5XcLupMk+8rT10zpfzK1cbfqmctu2Y7ZcXjFSkZns
YY3bapcuL+x/+ktYMp63SoVMzcPoAKY9Mx1S+M9dB21U8adVUSYjcoI50b6nZmVl
rRyPyT0fczpu7xmULhyjtbw3VD5IuI0y8rKOSFSpLjDvHBUXje5QGsZ+ABw9Z18v
OykoRIOStPR4iWok9eWHcmKN5wVW2wndNogEUfEjkiOWWocgN6uJ4NGT47CFHx6a
bQDYYBl0gmSwYG8aok9FOU0x71dZJcpwc9Td4hDrm5tUHpDp0pux+61F1vLv8x6P
9Dv3K/twOoxy3HGMY+9ru3RNNFoHYLaWaNf0m3HFkGsjLFLB85xiN7YwwbrKJhjn
XjGn95l40FmBAZTg+nfulZrfNGChWenHli8o7J0jyWko/B9baa6FzspPvxnwIrdj
E4RspdYVPTS5IRueCma1A8zifE6Euhfx25jWHmNjqR3INRpaYGkjoowynd8EACkP
933564Gcez9AWe/zP3qoLy+/AlqefA2TVK4iaHQHEYHDhxiEK4LThydjNRGEWejx
WCe+nvbZ5Wt4xo03XBnqcJ4Ezh9GM91qmjU89ZBxCvY/h0kZypYSxDOigvExoKCm
rbN28/ypbJwaaGInm7g0Vf5pvkflQFGDIQFYWfJmKLj5xap1jaIxDNVG72ZcvyDS
MISLnwwEOupCIc6PY4Lf13ht1g4S/zJMvWAbp3NpRsTNZ8VVgjg8DVCFA/B1Mowo
cihML2jL577KNgl50PqYyRDquw8bfaVHh7lvQBa4pXV9v3eaic2kzVsmT8Sfztqm
8cuINc5+ZBP9h/g6NciBiazjLpGGr4339eEuiP+jMfdgiOmgYSqaY0E4TjibSW8R
e7k7A3ncpFTZDcb3J48TpnvT+5hbiHgumcRGEjoEtokxgpXObyYKo2eoxTWCoC9R
rs6XGLZwF0snS9apJrQ+nA35fNNvJVRcrMHwIKkGZNdGDplyRSIziHbG0ErE7ly6
q2/EkqFpsPsWEKujj3qWH4bArMkr7+DQJpW7W4bV1QdvgFr1MU5ZJAZL9U2x3dDz
rU4umOZWW0FYRLoNDthCkgiW9pES5XXE9VtidRRpMZ5qGcUMX7Mcgp3qz8Bcef+/
qFEGfOFlHMOB1fUtJgFXMQq7VqjutpdeAuSNDmINPPNtn9fzkQgNhElgNPbn9eKS
5Ryq6BPyRikhzB2+UGV2ZSotNorYgNL+PDxGGFbYjuKV3sbzTvgZZ77RfBq5p7Jg
0kBwijbN+td8vi5l73OhVVP4/vNGWaeRvbJ2kQ7z7pAQ56U5xhW3w+QfHt5vEJK/
lyJAxwUJa7u6Pv2xJ56+CyT0onvSOo1GfmoEYo177YMk7Kwc+o6G05sTi4VZBTx/
cgrnSmA74yZlR8Smso3Bsg==
`protect END_PROTECTED
