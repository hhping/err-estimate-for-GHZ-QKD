`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfhjW/kjKBMZESU8TOVRHR9o6Rbw2vYdGoA3O0PCc8+hAKHaCqhsvQfMglsuVhPM
1KhkUh/BLMhtrv+7tAcQIoY8ufR31m5RhTnTBAyn7JakdMyfSDMhKHJngFwJhzEQ
13Ksjw+xriPMmkaOpBZnzwColoZDCEw9tmEeE0a3vw7wtT+bSJ77i5BH5S2FuJRX
psh2VvsEFs+OxXFdxPwTnnvpjqjsPtaAeubqBAeviqTXaaRHH9HcQvIobFNdEkyx
8vJXCD5T0HpzK42OGcCn1w8CPq2/Ci7BiBYy5d7iZdK5G0JtoTDqwpKzWElDT7Ck
CzKVIxVDbIFbodzFG+qfewhC2F5K8qERFHZYqrP6Lr4omLrUoMZFMK5JDAPON/nO
Tnk4OkghdDFtZzrW631eaw77cEiBXtGWncetfuws/y8rLAMb2RK7MNqL9Vez5kg6
FskmMJopWyDB/deBS4mmTe7mW1q3yZWbx7GupHr63/SIxWbvsatJpVJ2pKxzmLgZ
NesLn+dCATwm19UKGDi8DKRKHrjbe9+xOOUNQ2Zm4lLH4bH3ErkhJIXS5E/pPKNL
TmQ2OqDAqzoimWxIStVNHyDvZG8N+dN8SSLN+gaeH7H+MKag9zmhoaFqZ3mSnRLy
qK0upwJdUlXwLpwrSmNjOSl/zZfQCGxaEoATNTF7fcHnpy0ITA2yuP+fBxrr1jGa
jZZekikV+dHBk+wqGFUOX+gd6nc7a+M3r5fJ1PBIsEVJKnkFR+Df/MZqY19lyLvz
p+NQ33ItuTnJyzu3kO9B9VY1S4nTyzerdl4nsYBVldh2+xTe8TafEruXUvl85xnE
aqO2Quj22RlXQbDQLQIJzxzors/zib7dve6I0yqnY9XRsxuYoBtWxcf6SuJJM10X
AY7foJdVtUpeBgZnnMieIA==
`protect END_PROTECTED
