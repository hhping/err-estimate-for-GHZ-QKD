`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eS6Q2qnB1vbpPhAIujeIdblKzXl3OX2vUqdx6ekDVhruh4Wk5AEmhbdFVcffmlrN
8tyAlLqru9FomioEzfbgkCxvpsCalaslB4ZxQnMxbiV9t7MpYLqci3G6rHt4OS0P
0r3/uaFKSKQhTcxtnP4INx+80XpczaKXDsigfcyNjLE9F60KKwcRXp7ZyUY8V7qH
JfeSOmmVxxf9mkX/EmXd/QpNKaaEOrpsf6Qbc12dx2L3q5RNcTOJR+rU3HSviXUB
l83jbUltzAG14PFeee6OZBWK2+Wx4xb/XM5g4xzkgDECFQDXVXYaUeMdX6w7tU0N
S91xlXRtyOHrsGAal5ATJysC2Bbt7Pq2FrsEdMs3slmNog2WdDFtdOjgUtticcRn
ZobnoexuQ8LQ8mu6YQquRWKkqW0Cyg3cCvB4cXyqMCpp7UlsjGvk9YabUUDGRihv
gBET4wvWe0hqCkzdgt8JrUFXmSlx7KqPtEVamupiMLjdgWXrUkE99Bq+1EbEcT0B
aKYeOpi/hYgE+BXiaXDS9kSj6SkGuA+o8fHWDzbpiaHEU6JaG9ETuwUsoC9OYKXQ
cIqcrDdtagmXhNH+a7bXexlH40QIM6i8aeulLHeFDSongPxA0Iha1eU7pPSz4nXW
CeuMNkXgetq7TAtNuIw1qp9C9l0ha1Z7JVuqwEgeWO6ghhxSyupH2j6A+DQS41sV
e/omCsOKJEbgoMpZZ410zvdebAi54ItrpXO4wMU0tZb/Zf9O+zuinMpZkpWIjMFp
xF9puNoM+paa7o+8NaYzm9v4VT6ffh/woLovvE6VMuSiZF2Qnl6OfcDoF6P6dgdF
YW1lO7vUn0r1Inl/DmjH8wePXwPs1wtUnO8gO+luxcRZtFBs4GJu6dJ2rOXTnp+N
2WG1xHefW/C8ljtJimGM8ARo8ej9ld+JFMUmQTOWoElkcl77QP/UHB3RaA5QQeDg
wWW6TyFOoVaupZvG6gn29TB4Jwz+YdiIFOxkXJGgiUK14qafubc+Y/GCqZUqWdT0
jmEcOerACrdF0B2jDPnT5T4t9DDT7pAFVn1wzoQp89crLPWZV2mC9Ma95YOcOxb+
I2656fwEUIGqQRqysIhB+HBYOuqMOgSNlFofif41V96sW/c1GJb4IdILElbtuO4G
aynjZt4IiG8C1Wyn0ngAvW3NMVf+SWtjsTHa0/u0E0ZXTTs6jDBXButwm3itPbuF
/YOiHKADZBqonx1/aRNNYKeC7EDZ9CwAR0NeC8/JIOEMovI9RMp4fx8i0rQ8CYS1
g7PPC+5pj1WKHEqmkIkluN9a+08/COURSo+Hm4II1dEtpf758hEKtkvx5i9eCmJc
864to3YwioZc+8QU1MItnORYAB4Nu74DFIgML0hc3T/INS34k3tW4sGU8LIZIb5H
KvJT5e3fnjcRvzQ/q1zFm0gtCCUNgnl6mEbBPtX8FMXAnUU0WdVGwb736pkFX7fe
wzP0EKvVzCPjne/wGNtZTh1QAZ8gP021/H9OIKkDeJwlbOlwZgSUq6+q79wsoox1
ZtjY51Vsyh7IOlM1tMWFhTOTLoEZ/ee+2p2lz+pH+PxW0rte7V9rZp1otJuHKS3m
GlBAyV8Ij/m8atTQpxYtd0Nagz2B2vlvdkkoBa2a7cm9HJUw0PsT6tJLSuXKad3I
6IeGiGz4qxoxdMt2KOP/FJiFqxCQdefwsnATpO0LPmo=
`protect END_PROTECTED
