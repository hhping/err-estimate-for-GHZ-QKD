`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmYfXu9O7eWZQHZUQmb7mNCjlrGn9nfFmPbLDeF/9IPmEvDSRDbaBXXsDoTuOhPm
1sftgUgIwd/719XVBzobxXxOr2MS8YECNuhd3r0z2BkgW7onXL2oMR5zXpucua2v
ER1uYnzXfWTESkF/8KSHsBSdjPCCOSUYGVsJlXj4Iequgez946U+nNCU9Lf8iZ0G
UDjPR2eQ0RvTiZAQhB4uKvIrvek3y24qVZmKhAwRPEuRMbTAWZM9lLwTdh8BuBTZ
ScYCDgZCjktENqdJ3ODPEj4Yp5mjkiyhBLvnpUYvIsu8ZISLEO5IabTAYHS7zurf
N75+mJbJBsi1LI1E2qNqg4HDbwQUMwiSpvdC80H3Yc1Mj0J2FmcrB3IhUkb1dnJM
Jq2rPil2JBGb+DZ3FpBoORESZJcbBn5S1vcb6n05MgvbXj5791sYfdkmYEdCozpZ
5WRLgZGeC3CSjySI5iX7aZIdkq9+hMQCAa/GRxy5xROFwmL95T9IIBQfNtA3Z0gH
lwpNUwzO8Hnt/tprhMea4MdDDLekHKNBf7you5ES1PnYjFH3mgiWWx2i7ctiZotd
28I4/kcZjdfxmPkZGuZ8BsIQHoVDQXrP6w0lcrlnJIb+ObierEcjIB4WICN7KDJm
/xgjTNXe9uRlNqkLROfw++SZ9MWEpI+7bK6HJ0UuSUvQhcQQsk+NDqSNvo2SNhsG
YL6ibXs7LpWubPjQFHYsF+4Ik0vjzRYVQmbgRxQhr/kWF2D6W93ILo7uZahiPo5J
MMutoLOGa7Cdb4JdMzvlQdh7Sl/eLjzOyvjNotVSmNTne0mhTcOGMFkGZvJtf8X6
6nC62JDfbLSsDpAdt8tNj89Ru9Q3131xa861YMGG3MZb0EL2omqGO+ft61abPNr4
VDfYlp8EcyojiGU/8LC1OffcH2V7Vp5nXuLWuUnlLAe2b0O3X7u5Knk+m900Y0qH
JatDY+C5LhRVovpaExRSjIHsSgTjUlSQpyCHqVDisIE3ocCRM8Y06Xx/6jPcp5WS
gW/u//SYHP3/00pWbSAyxKgsO6x8U7H9iRXjfmLxf+35G7dtzE6io7OlVp9dpZFc
S76EX3oF04jU6x4Q5Cog7I4OsoSot6FF0e8xJQNL6ZJMCKQNArchRCMCP+W2Vnwi
sfIGHhvXYtLtS/6yetEsYpdmGyd6B1S/0os9BZEwvS+lYu6Q5+iJM0cPAR9phTnD
r03gWT2Ik5kuNL+TyJY+zUAEUnM/Z+gf0uNvJNcZhCVnAhPpdnfugelzOqdssnLl
v6P4BS9X117sx6vbPT4ahV9fuX+JR7q/mOZhrp0iPjGMFBR0akiSZBRV3Q7ORX4K
MuuG8orl18q92Eh4oMQR6VuGqhvX8MFoV18HPX3WHqirQhIolDI0wuodvKUu9UyA
Hh12QqnsEe/J5x9xVElnjhO2tH1SKgOa5r20QfUfT2ngYMret3bwvvzkdUFm2SUy
Zrt8U/iPeUVpKJVvtrmkrr4ijrqQ79S3oxouwdcy8rHGPjxZhwWycTv5rlsz8blW
aKUPX/d0ZIxHYZ13ewzBGW3GvzvbLfhx91PJHfIv6avDQs9r4sDFd4i10OrLG66e
bXhdVnHO/o5c9dHPbHIz+es3buAD2r5Btmn010YiIs0Own4sYqzBvlwQJLrDbCQl
Ue10eWLTebDsqEojeztom7XFGx+jgOFb5Av2Ql338SrD3EcHJ1kNcrGtMWs64w7S
PF/b3MsgJZys86qBa7VJ2zP2x2flvkodKJMiYFDSNiTRRbCvjVVYLlpmpC3BOVLk
fd3aaycYqaJD4psZRwO8POCz1S6Q9BDJKY2+pi1rYRHPkHmCK+ZRH4FHcpd/iowR
KGdB3JvfFqgIDilYcOGkziTxpexf7Cb1SK8e3LW6osQQbPFwPGscvhgyhhi5AxZz
R6ns90S9iEgkX33Y3zxOvYsv5eG5YRxv4JcPF7uA0IrxsKxfwpnDNCDKxERpr7NR
+VnrpzmHdmT5Af2WGgwlO7bjIt14LKr3lizzC6GP+dSIBya/U20xaM8nPix/+u9Z
5LshX6DJyBPeRXrhKwAwf3Dkpje/BkxhMiU2koFUOPSZAtt0Mx1wAvu1qkok9+HB
kOHMV+ruzrTkPYh9NxR7Et3+TUNVqxot8/WiU4XA02PdjwLUB3iieB9tUdndCZFw
1LE8uAtElAf+f3klvpoKjEiZfKJ5Qt+rBMEIBIfoaCOvxSdnUlNpo/nmeQWwp/KG
GM2q9EJ3SaNJ64sdxrI52Tgt5SJfCeJTdsp1ktVJ5Lg5Rj+b2dRa6P8x1XGe1Sjt
tLhhvx7wKDip/ABsf4EmuH0c/S4dJxymCTHnSxKnmHsS3e8hb2rT4UlD97Wr/OVq
RWIkCW9AlMYXgadKDn43X8/bkX8oJWMCuSDBdb8abKUq+UQwhoj5IFaS4OfiveZ8
NptJZkfe0DFZH3NLI3uO6n91ueoUKc6jxbOoP1cRXqwMlI8ClGTAzABgl08e96pQ
FTmfY1nHtZoaup3HlVpxzsu/WhGe4K7HTQaHjJGAP+4q9cWU08bgeDd8c7z6cQC4
ZNwego+SlbVObv2IWlEdIv86Ijp5bi9WZHRsaKkTQqLACHvogL6x59J7SYxzf8YO
ZUmEYu3Zsv0/m1bJ2Vus/aQ3n71PNK6PSTqOh1Or3NC1HNnTMjr+N3OOiNTPubbT
L+LDoj0yz46tWKnjS8cP8JxF3fhRuT1mOT77RMTaOQhCtM9cUNHt2iga237ReAfe
Rwb63eDfWEaCsyKUiNYZFV0kYP6wJARG5fa7jSG/neOn8pin9nWek9E5dZrXn0h1
fkPb6fC4Uk7WTCr26P9/ijdwkynq+hwSntAmi+q7RAbKD8XfCG/7J0cQ0xxRiJvx
m+AusDAI54hTcFn1NClRi/NZAE3tBiCM7mBKXSFqOKNrgLQLRsm9I5HO3I7ihf0Z
5AC+Ku0OwXUusWQWemJQke+J8lrxmtzvdNdE++3vzvLw5gOKnIjhquP5sQknwLLw
i579aycHroDSarnvIIb/VVemNSGUn3jngxYcvXNmmM3mtFIG4sZApxM5bWMCCR4B
XXFPd10Ggkk2SlRMNtx9u4wUOpRpImeDnz3cKm4uRuVpYOVbPVjXKjB2ApNB45B+
Z7gB0vAYT8V7wO9lexmXMFVZJdiq/DgPdDPqFKo01QeaRIZ/wwpiHvQtNX99hw21
dZ401IBkY0Lup+vwSdhkJOyGhHRRp0XuhWccezet5/rKUAgDdBzZw++H8DKFWDEl
xcgg7WqKhxbw5OCzW/lwlPas7CbuLUf9008/Q1mQEB+xB0up1LMfjgQ/V9q8YE6q
zfS+dcynHSqTW6ZVN58epDZuK55PD+w8aKpjF7UQE+pZuHwJ0Pc2HNcyqoQ4N5GK
HGcl7YS5HugsY4FNJNZ9WCAe5eij8Wd2q7rkUCZQN1Vg2p1N+rSvayInd4D6lGYG
xn5kY4/HxMYnsyGMw4KEKsv2gk7e+IoypNfcLoicUN3lV6N0E9fBRTuPUi0fwfKT
g5mdkVvVB5mF5sOMiUnVk2MxPX2L5C80BXX76y0GWkCZfWeEh2nVjc1Y+NVbehvE
W9JICMut0UUTUMVveQDLMyl5NcBDSrTyH5Y1hizi+3iQn4mGa99nxg/onRDDDLsg
vRTMLFFMiu0hr66xIvsYZq8G4f1s/P8viEQOysCyrbZskHJdUL6WkuslCoCshVS/
M9g5O6LDC85BlvpQWV+qCdWERLT5zXSqnMqrLytMoB2ZSksbZuenbTIM5zg5DLe5
NVPwHNCArKZz7V9WOzzOKazavlWFWQEF8I/0SZujBBVD/RfD/eaQ57vuJnRjrL/R
uirZKiYplsKwAGhP+sfJ2/8CgXYvfIZlzSaPDCsnVgG1424kQiOWQ00qy9Sayz5S
vNZ0INChe44b45lkH6pYvMCSdFPXn5LkHpyIsfH0KEmhcYX+IWGVBy3mEeGcNVWQ
S2/Znhy9jOMqRTntz8IoCi2OwMrHXKsUp/6vBmsjB78/tlCRDHjMftrZ/BjOlzd8
5pKHqw7lplN9/c6SNK0cobS+37hZflmK1E1qSPOATtnQUaIy1tWHX4pM31IzAos5
+mgzygIZMGvNGEZyxgn04Q2HbTqRe7Cd6JMVjWeEGVMgjCqQ9kOh7gn6YM2qBnS5
5Ggqu6nlZPJW2D78jH8Zc6qJW6hWJRuZuszRxbb5yqsGA0I0BaahkcFnMimpghmp
fBGc9QztfXYXF2Yya/oyPZL9550eJ47kwlzsFi5qArK3BsPuNZcFnaTDRKBzdqGV
/BF0sDbvxn0y7E/p4J2XtcpctHNX927kf3xPfchXVEefwfnzNbFoPSkh4Cg3dIEx
`protect END_PROTECTED
