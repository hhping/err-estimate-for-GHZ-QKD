`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylyV8UCfXGvUDn7LS6vuno5zJzQe77qXC5st/4B3L3y4/bK+2Js/OHv3H0/9UfYe
KOdwRO4JI3GyvHyc9yDZVPVNNPOH2zRtQ0c8d+SFOmNfDLp4kqtdqlNXR3k+dqyL
xCoksPO7mIVs2XYkXO2iaxByQwogkUKXYLWD3HmWFxIWe1V0YkkZLgkItuAyM/s6
rQNW0nJJJ89nomspwJed6731P7TUDDnqkXxrpzXnaSR+xHxuafOSeMoATnhVRO23
jsVcEybS29pBEj6Oed28XPpBqBebbd8/l+omai5jpgQL7ZAG2FD664+irHBTlHEW
ly29T87AiC6RMYSByNWlRXTbXW6iTPazFKKlnrgjmWr42kHPQSScHt3/FBT2CJu8
jXs53e1FefWJEaMpYwr/FxrM0FTyfHC25w+OiR43JX+Gmppb56V1yld1xj8r7W2T
rVzhsdCEDKKDYW+Cckst1JpOzKfWTo/t9Atb4PGIExBrpc1/pIqZY9FC8Zgtjq9w
5BWl2ApBtb7h19lgxOA0Ot6oP/PBMHYQTihFCSuznfqmPR/F72EJMxOZidQwdNfC
colqCJgU9yunhn9mhhYv+8iWETcDkBqPG7CB5VHMRA3X9b4vfQReNntgEjiwLb8O
jmMl/Y6+p52iks2dRT21txTXZR1RlDiJ5D5/wnyWQMzurq+DNvg9qRegQTaqYTOH
m8UIEFBzADWILq/fE/ps9twbKPJXD0l+J7JulCuVcZ6w4sb2DE/J6510Kpdbsfjm
mEUfHz05ZriuLtYu4TGK9ER1LUz4ffbMjG5xnjRAPIgpPFICH/brJgySW56GJmv0
g4H5UjK8SyneZclg3i/bUATvVOyYK7ul1yvkLk/bmAw9Wm0DyLwJ1gqFAbUTHinT
N3BbjoEGKbDzzFBIKuOMq6+iy0ClvhAJ/Vjp1+F1IFcIGWBBv5TNc7oNDBoJNKDm
Tu0H9nROnalUWBD4s/oEdLFyGdvf9FVpDmvwXwZl7rIJt5cfLe2bP/0bSc2q4YVD
jG+CmvEFyiQf+ZZ7PMXX+WYwAIpjT3AIVp4L0YCw2XTYxmB3sjqDE2AlSr7c6FEg
//QnmvO8dt22nIj8ugpZLzvqGDnhNs6X7Flb+13gJP5CG6bgGEaSxnkd9BPsj90r
5B3BZ6YSH0Q6yyVWGFP0EOP0SwZ7/wD0woByV1NgrJcEOxhh9DNpK6s7VRY96Pni
vnV/HBGScnnt2TQZIOr0N7hSBoqC93K7iTn5rY3S+xHVQnqiNGdeXjgyMRgNuqhz
XDQljdugsX2kjInrOhYZSbTXbK/0C01yYyegQVOLu5H7llaZrmhburO9lJfLYU6j
MyWYEUGGDUjg21/vs/Q2stoFr6QPsL5r5t7+Onakp0WYwrOSjajgQVIHxvcgmvcQ
tkUdxsxS/45p87pL4GLxX5stPw+zp/fPT3lpXlHGqLd23aVt9/A2Qxyu8gaJshCv
z+K73SDjNBEwmCy6OUAA1F+rQiBbjqDE7E/wrL2M6tV/jHn+TLNy8q7lcJW+WVb6
FQXnlgtQhHyt9G5NLjFLLLFpsuk+8Os9x2czpe6NOFF1cshZR4Js/gjdP7kTzSvA
mlkIDoRiA2kJCAvcvwK8asG/M1U7XUwPzT6/tyLn5AE8MNgE0cjVw9nHyy2Jb3Y5
1IU24qaVrBJd2UAeGew1lpE7+KKUvPSoXIyIc8fblnUR7M8QUhITavaKCtV8p0pM
NDtSgksZE+ccsbcouH1RNoM9+13ZMOFICH7VsizJdbN6ILlPHe7S1xKPgkfucpWq
nYP5Py4wj8BcE581ns6U41vJkWtw4ShY6OkKN/zNAHIrMWa9Lx3jqBZca9fymZze
+7TlLOmZ3C0Y89oaNkVuQv87e9XliFHiRM/b/rnjeCYZM2KmNVUArL1hvFhmB3cz
p3+EubktlBQMFYX2dZsRqam/uOkHzWj3SUx4lUPmJzREaR8ClhO8TBtjOZDPK7r2
hIGw2hc/6j+spzXe8FPsEE/6F/d2eInJJkE4H9c/JGu3zC1huh+aHVEaCm7uWRMK
Lz+1oYFAxnY0nHj+/53N81on7bajSS4bFZFT3BKUvsD6i+e0Ebvsg1ZVGkGotZRk
L9j+yfhoeSOrA1X9AGqvl1XjLna+MD+wWGxn5jb4YxmcQjX+DlFy9lgXyYggmN02
TCQnRcjs8qq5NZOkyyp6xoit+nNIOM1e4NIJ+9OEbsoezKszouxbNDmPPzFILlTR
SlE4dFYd2+D9QX5+WleQmnapeJ9CbkKRCw5pZkNJeqz7vH+MJQy25eWn0tHI4U2J
vWC2p0+8fY6CXmfSHqsdbUreDoh7OzUkdiLWHDCzHtukWTM18EiTHuTe95BH5q9T
f/RWHVFyS+yjcu2iJ3nqD72deaUh4Vf3lNchoVKVMgChdzd6c/SpmKB2SCUdp5MK
itaCAsfiSjiFS/32qh2hBsI90wp2+BfCp+wZaigjCjKjYGVxRQosRrsi7TIFlaoN
ezXoMeZyZtEy0dgGhqO2fYaF2pNu120iRu02IyfnlkjtRzQTOi3lag5AGhxcxdu8
YEjO/i8ZB8/4KRR1i7HvqIK24hz/ZG10luQtN46ZMvoakivzYKDf7zWnxwGkj5T2
z4PxkkmmsdgCLyOz1QpQxifW9BmuQpy7O3uE9X9/wgasE58hZeoRr7QnpDgoAa61
sAGZqVwRJ8WCchtEMdEN9YnRkhpd2Bz9tQeLl6HWEDlb61QBTPaqB3oBoczFimae
SbqrbPn885cu4WASDjZR5HpfjO1UD+zmigshQUF6fmVh2TcsybGKiCTQtpqJ9M+e
TzD8xEaH31E7cReNPrDTRLnxQj80g6Gml0G3KNcgKOXVCd7e3yT7v579+E079Cf2
qVZSWCWVTHAij3wST4sNqItmgVzy/LZXjFcRoClqTN+Q3eFP0lecIolJldFsHwAi
aWuCPLw04N12V3+ULo6X2fM9QkKv5DgJkRprFOpEVkX4B4Yxih9BPhSjJspp3Abq
DFMMCH0qFUh+/u6xhWK0p8ZopDJ7SRJ4tqA0VkiETdquqQvtbu5OcJOvuG/dTfWZ
MSuQUiFC5nrppesLf44/KBV/P7kuixS44FE77sllNqxtgOCqb1AFNOxTqOdXBZ+o
Xd6JbahxYM7hzFMax74Qjji47Yn5Y58AWJPmAAZY70k8TcQ1x1PVonicfFEZNHc5
nZYtNs8zD9N3asj1OtdBjqUog/S9gQLa/wIseLhjHSnOG+spxICAo7LbXvjBnXQL
W/7Aj4oHxWpMLvHN4q/1WmO5zPxhW2cmcGcqVTDlC6kERuVQt4dgYLp6IvLhPPwa
LJfmNG6xrCKtETBm5ZcPKoEshcT/q2mKf9O30w3xhIG+VBZ3xDlrHqcrM51b9LFk
/qRisaYNKhFVYvJ8ERAcm3oJXxy5B5PlT/pe8pcdQvhDNDGMTeZeQtas6VgcEFor
uAmwkP7Oc74zRk/bAje9j4sbhVpzjoxMfgVQb0pMAfuYCyYqbHvTbDWzGuo7AYqO
f+dic59A6FLtDMXX19y3j/3/9ZLArr3ElAqRe9PzKGwzMVc5c9ZdEzUd9Ah5j5on
AF/Q/H9geL/yPOLkW8kBR40tA/IdQnRXCe0CgFngYoTWKdlv85oDC1BMb1mf7QDS
iDEyAESb0NRoOVqPMdILTMB2NbqniJvTpQd84ahWIjn7HaNU3c/RYouebhyCnrkG
hvOA+UJ9JTWrxL6xvrYVgA==
`protect END_PROTECTED
