`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6O81JGTS3OyrAvYFIpAqGG1fphA5+N6vKfUdnT0nH6Rn/Q1UNU8yMSLLBU4Yq11V
8VxGjLLsyFcP3J58jMnXgdWbBpqK/llmHcIshh+cDT7vlzNrJv3Y1CEr/7T3ST0k
b8J9cslrnZpfK7YbHrq/A/NvhwzOiQTNqaSrkCM2hpAfDYLFJPspDdeSoeOyfEiq
m31n8AHYcyVmK3Nq9LfioBM/qqcBxIkcPfUI5oFxeC85sELvSbVP/7K2TrZNbCJ5
ZtnFJWMOXU4vn64pGXYkK/qJYu1gAKOqvQml++LIjlcg84mqYw8v0z1vPgqYp25K
m8gkYNrJSLEwo7ibx50VQ5RgR3gyG47ymZOS1jAdYvTg05YTg7vWy5CO+MPDBUE9
Q4XO5WW9r6/Lm57lnkRxslv3pV0DtnC4tw/RZFZfLngsuFMWBh0Ag0xVmXB6YAPp
Ot49lHLHseFRuXT2l9TAE9WG76zOkRaB5RymyJ91ypS44PbTHJZcDoD4cy3EKpaq
blWkLKpIRMcVapVkNzFsJkF09PWDd38kyFEnM1sYNo4EJqf8dUyXhBKhseSgKIqR
0u6cG0kTBRTFpPW8AeCrSASFK/MYYpKiliJn2xn43yruyZVQc2fkDtdOPxpCcTs+
uVnbCt88ofwrOdhSAgCgGYBC9XGSUAVekCvGA3aLe/3FECarde4sKQ4Gte9d254s
r/NYWlq9SFmQ2prX79B1QrXCBui+go4EurtzYROqVBAbvT/DJ4wgSfSBUEg7ZYbi
`protect END_PROTECTED
