`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWYEi17yPQwksDv/oufk9jC3rlh4QnRpUg/aNjHhYxECM4QT/FfnGGp3JYBgicWd
H97r8UB3vGEs7jQvhS/ya+2SXEE7CYHX0ytv5aB04LVPAHhaKfNzT+586cuYKyGy
BEVoTZo/duBKA5aI+W6s106zaFZINA52l/iv0E4w+gLmwt22ehU8fyTpdRjoKPGR
wJPiktuFYNa3UE94pVWaWc3/yKAN/8DfDwaI+9aUoQwmPnirH2WX+LYcknSuk+Cg
TeEyrLiiCWi/p51GsTRxWM8ExD8or4y8B4xJ0Ql8at7lSq8G7xeL5MFySym//+LG
jXoyBY3g11hItWAh5WanRLGkT36DW5QMbKDkfvaAlFV5Zf39jAb3jx2EEvjVN0Em
MrMzAqB0cSbE0HczoFW47UV+InvcU+A0+lp3pfGsyJsZ66Tqj0tcLpftj8ZqImYF
4OtxYvqibKGQaVLsE8XrXkpbSX0tShEXPOckbCd1bilL+pLREwJvABPJ1fFwJ650
QqzWDnq2ftL3lOIPtgwIZBgrMYUJD9/T/BHI7aAq7kMJ9/+LjeYTkIiFJccD3G3/
SjyGJr5BLfHNl2fzFfqrMOyCJyZKC7TfGf2+9o7mXAU1pv3IPIm5F3TN74TKARzF
EIQYcMhDBHzwYiuPWnacwuX0xtmUEA0V2Fp6JhpY1dNiOBZbWv+XXkSWwTv4fS9l
OQsF6b2bjJq5UZmkRKSzPWBqt3M7GYbMrtGZ6Sq422RnOGJiMfjQI1m5E210bfD4
8BO6pvx5oNi9hKano6sJTxRYh5mnynQno87NkE/it86iv7yqFWXI9bFfb5dy9M8U
yJJKtIwPxd/mo0yktBpNrnfmKNtrmLftSIsVCEja1tmhlq4MngdNRuM6myYVY3Lo
yZzLxi4/iiqUzSi/Q6taOduo9b7IrJPEIdh2qgIJtj15qI4TzFRy1c5H0MAV4O/5
jijjo3sApLjHELT4GwfYBZFVgMb5i19cwSc0TBxKA3cmxsHqudYBLhAwEG9yl4Os
TdYfwY9BbqgvEdMAhkMaznPT20opdVhB86+19bvXTNDPIYwHPsxllI4sVz1Kdzje
KDyOHi/7X2g+8GpJFr/STwlKc24qdwSatDVf4pScms3GQBN/FUuxaovfgu9BzWI9
4EMESEn4jOnlafsT/tlarwxVwmNNvbbFYCF2zyfRneKacrAmHyl9DOw77RLjDVGU
3knSRPV77AXD+9TI+28v5uFoolxdF2R30v8EMUm25kgdlMjmUBVYh22fG/YgPepb
MZMKs1azdgNrVSqK6Cke6RXhS+eS5WhtdgdNMLtfC9pdut59HI97jjiW5yNRbaKL
Okj4FxWEwUwf5AwhHM8OEBgKdaD5G+RdXGAFO4yyhLR2uNgUYHqQY/qn8N2z4MjT
DYIOkJWCCczyKsY0n5v7uQtdPFuLnBoLx3WR4jmUQlo3qJ+y+MCyX4zfCAjCe987
dUXX4MkRd6Tgwubas6hY05HOBnyNMMxv2NQUqpEqLMrYRZd0CNp4gRol59RnMYYC
46oZOUMPQuoTvllsY939qDh3Zjb8X+c6K4o9lyAlDt470L8wvbDlPcZ9DHZlxq2d
WyW36GAUbrhO7g/5lZrwC7o6Yb5gCSyKOujcmYWaaj2JvMUrbi6OUlylgUg/FWLM
dSQ6ox5dIk7C2yjDSHm4JTwK0Bl6oSIH2NrjLqwG4XKWE6/+vuR5VwmGRTqu05ct
v4gcvtHYMTJg6jAD5/Ydle9DQqiUUW4v77cUeBXmY5/5TRTLtjQDNN9vNt+FxQWQ
SeEv7WuYwJakJj8Al81Ns/oZVQsrpVnDtj9Sn+0kwiqqLSjVRQkfbpr6ndPxsdRD
uBzSKUwq1lJejwq/NcItHUtQhs/4kuzeqzWWhxk6hy6Zqm1kL2CIstGOVUiNxTWx
u9IePDNmsxj8+ksNZvw4rb48sBas/1ETjZ8sdJEcw+dGoagjMhd4Xxcrhn7jQSlS
s2y1o3+S42YevB5QxUreF9AbV5aIimtDuxm8pcQWxPFlqI3LpqFKI2qJW9vZ2Z+n
5CR0vTAjOUArr4gG6A217Kci17+CNH8tlhy7dpXMd258u3hEKYVFNHvx00tEOeJO
3b0DJ/2h7Uprp3tP5MOLC96ZdQ4DeA1gnrwHpOnj8wo5rEJ/R3KNH/QYlMk8b1kq
z0yYD7VMYB/Wa3A6Q8zak3sxtEYtGum18DUkmCwbU6754KH4CyFNGg2Iqm986VI/
RIRS7RF4U0hIltIMXzABEqnv3T+dUsjPAmWBkCY60PI7RhVHvnpvd8MbTe4103sT
cKF22wa7qCtFYehJX5GLeg+39LInfGPdi9WwIswbrjgp6VptxTYtFjeDVbpDhxW5
hujFBnsuI1mIoLNXWhGYngLFI7NPO9s/T/Wpm3IdrQHticqmNrf3/TLq1apmvn0Q
HTGTV1VOmCIHgf0mKOk6xIFrFkfMwDWBbBgZVbtS0G5LE+ff1NbPKHSf5Yw5/dJy
QUiTHEoqFcgxN9zQ2mNvbNlQwCLsWEziW9FPM7ltQWtdCjqF6565Vb9OL0xM3cfV
ZQC6+58KxWJkPIVXFRxPFraHB7ZHc5g0lHGRNTuNFfy7BDRKqKj6F2RJD7jXASID
KGfikWn+y/aXIWHHzt5wdd0P+zU0JFpD8BjNAVscU3Ketmtvi25K1qsPLuyi1F9V
+M15oL7TgK6BIH0XBvcdOz6+znyTRA5c9tZa1l8OK+aRhvjTd/yvG3y5YyU14ENI
zMofEYxau5eiy/F+cnZwIaUMrdBFEdrWqt22JlRwNnfHPD8l/+8nTRevnQMFfQ5Z
lFs9W/1KIEbma/u6XGgCffKqm3EgUdas6JpOlkna3YI7ESHr0D3YsdZML+1potSn
M6nd6kIAhqa9Dgf6LxfKr0BCvJiNGsIqZOSZyEOz2f7MsplXNpNxdHSUVoLXKc1g
Je936m6Bdvttao0fMx+uOwWIc3rUyOLd3S/EAw533R+vEHQpOE0jc9EnYs5wIYZr
X5/hBfwRdjVO4WjLlhXnnKWWwqUEv3kmS8DZqsUlLhLe41Hrqdd/OOqodxvlwbPX
iv9bcESr+X2gNth8W/dzexTkD/jJBaxAZa5PYeL5yy5mogD2VNPK1cFvG2yBjn+r
swuqQCEhsBkBT86INftn6ZVReKgz6iWLJw66i4FDPWN95vRfe6cKeK9VqWtpH63K
iBGzkibsRV/pQKyuut/3/3MVx3/jlXSOe2LIcVynHaAh7PkoZMCZ6ITTvM6Udxbv
Y/yinn3I3gaxTu/lzj8/XjdHU5giEDgxLQOzfxNnE8GlzC1P+t/wLc56DerRjLFo
iaMYkHOlQym4PUaVu5Ypvt2KHDJ+CzkjXTgWbVr0vysLZ4vjsmpksaEdeF9uNVAj
7cBBSouqhADjV0vcJXbKhiI4LJpLezK63NHT0PjZY9F+Z5kCm+ULh8s91MJDd63z
v0sZDqoWlGUB+jbSPm+Ut0flbMWA99sq0Aw752S1PKqE+V4xBVCnPePZm3916XNS
+tI42xY5rPPY69HanuhEiUSsIlUtFOTN7OcbXzboymU=
`protect END_PROTECTED
