`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dEg++/w+mzuluoXemaj4kodAFwmLfDdVxgUEK6isx4J9hyCmxUhQVkuFAVd6UWqj
SUhfsjh7eJqS4zSJGBK4maZMziGSMQTl/zZ08nTFRc7b9KRKjuI3v/UcTEorrBLh
gHxJwbfiMwI5RbzOgdWRtlmDh9dJayXKnDO13nAZLotvnk8VA1NYAxQKZ3Q2VDRr
LO7irqwpKsRGlhlSjUhIV+AKAktHmzSAYpYVDCtX6BrXHcuRupgvgg2kKypwZteC
dBMMWQ2dPm5m5+6AC4FpOrb6/Iev1IsOORMB2POXbhPWCu3d2fbmTGCdCBK7hutX
RsKOqFaxc1/UNZFvmUx/kLpN0hpyWs/GBjSh40V21XQJOjsFdHKEVjqu1Ycoa62I
QRj+cAqnfipf+9u4fl1o+xUBw291qz0tTnQUbVhI2bTbVY+Dn/tFWscsi0uM2FGg
EAx3obJF7q1fK+L6ema+kqz7tF0+4DSYV9N983Yr+z+80KGwA56stu0Y0UdKNaaI
QaOREEbkflpD6E9yzrMpHeCq+NdicJoe6YgLBnOj1F0Lev9jTXhiSrmZv8ND0VP1
owAn8ep9o/4DKXlpn4fQUYx2gWtQCpVRgCVgHJl/dvHLbVYB84OriLu+HCTI7u0V
mSOEZ9agrMzevmAHB6fSZ/QtsjGsCP3MU00hSdaEGy79it2PRdluCUyxND7aNOkO
HONNeFq+yCCUzRVZ/OU5V0Eua2e1TKrhuhCOmYVoMgWqdj8rAy1zqh0Ze2bFEarm
9s+vIcCM9pOFg8AWR+Oq3QoTBiIDQED5EOxOQQUc8ee+h0CVw5btDSnbjjis5Rxc
p9CoOUnOVU+fYfXAE05wWUrTQEs8K1ZOMyD3kr25gqb1PUbGlxAm3//5eh5Wdlrk
P/NZdyU0ScBVWAmNVmX06gEb4zR9D9pkQb+tAlNHPTylwRxg8AzVHsGeMtXJTnc0
+HLYAmck0jS57Q336z1CEG32ONL8njBtI1X5v4lfvc3PHVGf7GKFqJw0pGRRepdh
4ilYvzk9zZPFd1cGQV4bAqa/SyNONVpSLit1Q4DFXMDDrpdU4XMlUCmJ3gP4L2ct
6c3nBO4KwtZ019LAymCepguIh6M91Mct559oUM0+KOYXL9d6DMV++nhX4DDI0YUv
pV1rT0mE56QquIethzbOMr/939NJ+Wn8pUcjBsDCRJTSJ8IPu84aFPnkPIskY9N2
PspLMI1UZjEFDePe4XGvKqMPohsrdJty8ImN2WnZTePVnRHxy0MGOb7DI3XRu/4N
hWbGPQBaHku3qOaxPlAoZ6PvYU/yz+R+YXQJ6bdl3mszcTDWa1O2gMzORXlRagEy
RnSmOn5/81ot5lQvhovvGy6Stxn7s4WbxrM6Y4c7CHS+mhpMQmOaxGuw9hOtEc8w
QnwvUjKA+wjwkIeC6K6Yr8d5yVZp3CVyKh+WBpf5dFSXlaBhoxFnWR217XBX8IRs
koIHiJGy2O56MOQo9DVJ8D5uKUAdP4s8cJiD0oQnzVPmV7mpTmJVAEg2Igb8b4kq
9dlLbJPuJiBgWCGhr2CClWJWvGb1L2o1U91UegjRLOpa857vCb1HeiuivrfPKv+e
0HSDTQaE+IxKJ2t1PO+LUuy0VR2DBYARHd3+kx1Gf79NuEZU0Um6+C8XXlzLJuUD
wSGkGmqxeMerKpNPIvc0yXMt7/zLyfiZPfFhzVYS9MKOQvIO2iMcgzDpLt8nCJWl
JcTLr9XSnhMT563exw08qJJ5N8KYJV8q+VTaZ36E6SLtDqlXpKAMdmDoWzd1S0RJ
9FB1H5Lk+pC/vLg1Bl9YzPuXK3MQ782YtAoZD3AVtNZLalCO6TksK0wVoFUwvf7O
XxjHjKg6rtjkMfvDt/B3Nlx/tH7U42WaHDLvLTjg2r8+u7kEpaZuGXWFjhGz5laE
KjgqgojBK0uFBsoqicUc5s7Vs7uBNoR8d7QLdPi4MFdQAdvmuDWakDT9Jv8Izsae
uKhT5mBT6qH2kp/XwvP698O9tQA5Es8VSxwxdOqloNw6FCi3GgV5YxFb0gODq7QA
d3fcJfiBB3yh2rlV09YYCccUaqkycKqn7YI7SSei1Jhk0tht+EkCRadCIwzDp10O
bYcIZNbHFvD1al7KYaxuIGo05fIdzaFZ38JufHRNWuZe++YEwUiEGZPp7jsN1ofX
WkF+Zr8bN1pkLRrBXWybtjJJkHNtF5K9Ecp4C/5uCcJLGnqOqP9jIhDOQo3VUawj
ycgoKf8s6AG7Jlkv7F9dmSOxjsAB3hk2SXKtWfI+XwN/nwhwasxhqkZNfj1ok94f
IAaxmT4OvBPacYcYpPaxxOnMBZhjS80VU8r7qbD/qWIqLH3oPvKCdkh+tjnBdk7Q
zeQhMQXiEtjsDaUzcwVkWrTBlGqW6b3mg2+PhjKnX6NUDoZTS5O+FuHELqp/sSis
JPb+ZfSlJWym7TsMoi/SNf1WDujAwmI5PrBTkVTZJrX3APDG0ANn3CBLyhec5V52
o8RzTACQ62qTW08Xz/SKu/QlLSsRR7ikGIHdSMysycYkqLurOUw2kRRzMdRT4drk
We8RSuFpe0xGSgupj9gtASelUWz/BRF6YiJKlsM0hhbmFxfEajxEJXLJdr9rZElp
wtsTX00LdWGacEuB2s+B49djp/bdof3uAK6S+Zs4TN7xTtTsVyjGBqybKhnVYB7l
9B1q/dv9tM1DfxywsKXc7wPLGAnmGHw1bfSFEEU+FciMZvTM6/ELcZdMySLArC0s
hcuPg3fNOba157zFs1SuPRTqMwjkGHEErRDrr+7OBqKSsPGGaH0cCxB6K9matyaj
BDVeDlsLXSHDm79cdt5Zj/fiRrQ9CqshDBXY0vTH7M+1xrvukG+7IFgbri1Sy1ux
W58gLtvXr6JrALS/S8oThSSfQr3mS2V0i3qPaYxxiaY7xEKutd9jCmNG1CAw2gkO
wl7o4YBPjRS1VryNmAl6/LXH+vtuYdYjf6rC95tWaoK2oDMihxBETYe4yOrmBeYL
dFH5vfkydkMMrzJ9PslTJevcsG72kfQynt0R4Vg4PVDUz0rG3Izm+qbKbgeuX/2q
4I1xdhewVWhd/xbNCWrQQAPEC91pyYdJVLyMP1OJc1OKJbD/78SpaQ7+bZ3P37H8
+9NHFoHxKSiUobYJ9X7fRcPdlgfOHbRJC7BGi7TLX41t8QvikOUn7G9xZcUH8vMd
uhLoXDaU1K9eEhhdVaNIy9MHU6i0Q9TYLwd5V2qwPbnrj9+NgLUGuCKJqwf1gens
cUEk6BNT6OIy+scrSaj5ow0xPD0CVjRkWLKoLYtsn2AsoVzFzajxjEYw0245fylm
O+VGVipt6dZIEQSxWLN8E6OS9vGpZPBgdR4CUNFsIhyKS9OYnrLbgqUvcPqrW45m
t+6hWTCPe/TjDNW14HuGP6rKFu7l1/fyjg3a6DJ61V4YqpQeilESMi8HCDtwE2bf
8sZuzk7Dm5lvC5a+X4xH9zdNn9oPzqijYe8ZePmPjv7POYjaXkwbOiw9rdWNdVPE
ppmJj6tXrBY7k8JIxS6RmnCwBSkc6WbdGexNFzQAGQHAjUlPlCHdIBUVvrKwFmPX
TvS3SsGZuMV1byYNOXqSRWvW/ynDTpqnyHM6yemBbqqlUscNYtytTvGwgZdiFFH5
ndzmOvj07Er1itet5yAwy63JpctCPNMD655X9+eJN9W8UtqiCuCY0879EwzrvpJg
+qJkxPDvJfw1gNbYxykRaNhFHhdnpn/kerki/oqh5Y6AUmFAa95LoFV3EILX6gRr
36kSLz1uhmFbciyXjf1TVwqo5i7xBc9BCAFn42UUXM2JE0MUsEG10HyCa3I4eZ5K
beiB1u7Nlt/hvou35P1TQlJvjZ3N2rpCTF2MPUIMcIGg8zs2pu/SHuLpNuAWVGVW
46g3Q3USb3pJIANz9bxpJrFfFZ/E1EUl2r6p0Q4lUQydD1fqnN4t+Nt4l/FzPj6b
SsP1W3plqMDfGm333Kza7JrUxDOnhKgbzUWRrFomGAVWDKGnZv1fs/KRXB/wxxMy
V4sBCv5+ntNhfIElTxn/6AAnMvt/HnmijQmnPX+00+3MuvDEcs1+HRRlTnPtc3Er
OVqHJ19ALrXPxJFcoJBa4cViItRuD4hqReiRDqXcVGyWluaRnwspqRlmdOAh4ElJ
KEbnM9JFq5O1SDgthW8ZZSOSR2aUEQST76H/zZ+/ivyDJ3j4zyC6TbBuZkjmLXck
WvHJOKxWGs5xYJ8nIrwJyBIMp+Zfv9+i69t646/IfBn+Zb+eRjk/p2LsSyZg9laj
lOVfumWa1SXeBvXA09S3yiO7N+DSlFcvKghsc0xzXhqr2vWgUhQO3gZbgQn2MIMW
EyLuO/8RpzeMDf7mGxqy6ng2LdY5EFsiOQtea7wwBEdkxj4ewqZZgt2MRebPt4lL
mkgpgDo7HDPonH5OIfFGPTTFH0spAJknAgU/bgnJEf7xbgKhQn1D5tlLI6hmXJ7i
bUrQgsTtjG6FodQJvE8Mw9hMdv+NHZHeD5zyzQ0OFOPL7GfzblEglo0W/VdvJyJ7
A4nm8QvU2pjoFanVmfjbY3EOijW3M4+2fncenPDkE9C8kA26D+ydmy3txBWLOFTT
oN3LLcl7jdxNmWBf2KmTt7bpJA+93VBspCQqf8qkC6R7kDguPNBdyc2SZY7yY2xl
wvAYGErxh7UXr6iI+RLDYJ16TnpCN6pMmM8smUOWWGIoU0mBtJvvA6/81CDdjjw+
ioDQuk3TOHmeX9HB4MhuiIkIgfDOCjKIWa1uGguZJVHu1VTWBl4+PxKEdY7+rY+V
WoJBSpfKcRm3nSSCK3/JTbeZgpXadIBxekwIP2bkUTGadcAhJqy/6jejPASNgoAX
/BkegwzqT3mZT5hVG/OvkCd7TTIY31gnlJ9wle7hmwqm2GDJjqFWGxqcnMBedbma
+Y1jgUCGK8n92z8QJqS3XoXFfrGWjXmtr3qQhHPNaGSbiKBqKKCJ/lJLX1FpnEDo
lC6v4aNOwlhkM6zUUNW9AUG7bysOvms4Wk+fATkSFqQXMW6ZniEjJm1g6UUBKnVj
gHPmeehz+WUCXPFWaKXitLECiRmuWTlzmZN+8+dMjiIkOCpjKafDmhfTwG12EJkZ
vHJyYsrjUhbDsikVeah/+arvHZYPnotMiPxcMxGcvxS3UdqqJ79jYPKQxatxhKX3
EA54PDE9vqvugGAk2uxdwQQIO/Zh7NKywwC05uOeHhf97WO6nZJZhz4VmviFJVEI
sbUxncYK/ItNxXYf4YvHB/qmXFrtsOUAzIVdkJ+18PvxakFOOrN7Brb1e62feqwj
fSGZoP5KJykrTM8MrI+hsUwicM1Slg0YP2c7p6KjJuBrXZWrS4qmCFr4RA0YTEKT
7oANftEt62/rkyZEkFHvsSYbOaA0kvqlfrWBsmTNymSn/eGxMHDRnL21Ph645sLK
1ej5qeLsI1h5HXzPxRrbu5p/3jYh3rE/p19QdZxD7bD+m/gWsxDim04Q4+kw9xxI
xFmYQsA7B5LpPRsBJtwIfnrWhBKI7/HGibeS/tPXRa0Vt1Pb5jDrYNS8QmJa0I3D
ucOKtITAN0raRfjOFBuKZoyl6vTDq9NbSuq9mdjqKq1aC8EP17Zv6xOlTGLn0zz8
31c4z6Eid0mPWqNL9A0kzDICgREGp3bvHNTNGhjIDh33cVEcAHOUe6caycYLoGcT
TfqPrKfMicADa12/wLyZT6J1Vs269BXUNFMxVwvPUHve/4sgs0GKMkit6pA0xUZp
UONHQa5UrHqCyeT9F07gKeIqE0EMMzFJ7MjwnWlSteRcqfAqoQ5gNMLkZ6ETNMcY
VRyyJ3YzGM0sutTQqJcePuaM0X3wrDJifuMqH0n1AqKxOetn9KcTiiBSxSqo6EQp
3Aeh5xrg09TXHZVt+TXh/nRBV201MrZyJebOSf+bfltcjCXD0JTiyCdATli16dnB
2ftBNxGcYEYhHh3uMgABrmRid67kVJFadTKwFJ0/+dguNB7zbnn7LHcRfe78mapA
0nszqFOEnYZ686LGKXbqh2iEoNokzG/napHHJMCtC837ewb3d2v3UAQRFWcnGW9R
cxLNdwFkQmOi5N3ckzKr+Ma+CQG6rJCLsbCPzMsgasa08LWOI1eCWwOydXAEISiM
9Qh7h3t9GTOzQKM4uhMbqrjZAvICLGSIjqpfucbM7W+f5CwBhp0BTZRQeWhTzTRh
PStMjBPtUWJLC0LsmfOsojVsaOIU0FNxkF8z46BmEhVlDDnVSgjBUX3vZ2T8PfcX
/rmk7IHRYo6sgvTZ8nucU2rK9YWQaRZZs/35eovtsYr3RJv7n+VOvwUO/2JFJgJK
dOjX3xzxsYdKZ/bVcYgmBFrWsPt9C9DYcgriowBUryT0yn8DR9JD4nxtdbbtne6J
7OsQGKOT2ToLYPacAbh+nk3MWbXaY9PEX46kH/dx15Rb+7u+KyQsNrZMZOo5/lwR
OQMKRBpNawXk31Gn16czMVc9hV6yXcWDW9hjcrBRjV0PPvs8qLkNzdcOnXofR6Bc
3irDZhSC9qeSWsDh0T82rPCYGQiztBl2JaVVEaNDZn6+znLbvtf3KbNcsGltM+1I
Qt7BSwtXH3xE8DS/rSFWYtQhFOYF6ipuhMaPWHXkxf4jlZaJTcufiOTZ9KrXiBYk
dDqaY/IYL/1tq9RBJ5T8OnYm1fTGnA8ouYo+UJiYqI3j8vvtuYplNqMbtQPsyITg
2RBDJd0coTa8NFIIsHhq+M71sTkMOdNAvbYEHjNCs5LZZGvEG5Vtv6dOa+oNqFGZ
FX0oSfXAy1o1lLAILnIwTBQTa9Q90PT+n5Aka6xIEoYriYSy217bDFFH9gm6sLKC
UUgl8WDMuH5NWEjMXnlP+GxRqWCGpifSae+eAsxyvd/8amQFC8acSL4lafH+lTkq
doNFfu9NpQZlttEbaV2ugbMiD0fFipdh8IcNsqfUw7FNsvj2MHtKyQxfvtbQC/Xf
OoIs8XA2v4NuioJZgeetkdqUPCLlCOuuF9t2vIz/gtPTybRLAgtYvM22KEQegrTw
Y17U4yjQu1sKCApaY2imG2T+valWP2LT484qzAzuaUiWnG/q8ew2CDHf+yuGu8T3
Eh3WVpqYApbnynZjieVvYkEUVu48NLGLdQG04u71uu3pzIjg7GxfzbLW6qv+eZZ/
TTo3vH7PCHpck2WKLz369hbdmU/Y6FSndtruUq/51BYPO3/gna/HZjJcBSBMs2ph
ssHX/kEC5pvds0GZI9iG6Z+kTAepObgd3X9TOHPLUHy6Zze5Uo2go4ZulosjVaN+
74qfPUugBoCxydALLqePhNflv4uleX0JHn1+SEo+SpwBaq4c6JDIg6uXulq1xflc
mtg3WU3n1a2t+fxGKJ2lxF+sIAEI6XyyoD3QvULesGJVsL0aoXmOKR2rMnhwxyye
IsSHVfv1pJ30a4O8BpN6SfjNBZ6x3gZGKcEt7OvktKILHpcMJ+6Gd1hKvHY5r6fe
nlv5muWAEivGaDvUwJC4leyL0JxrWmDHwg8p6camHjQPWhylW/aXFWzm5SlzGYbu
pUFsae5SKQ1WoApBvUe/RcLg/O9yIp2TA/rlmm9W2Qt7fMTaKkZGPI1FScAkqraE
GAHV3w/NfrJQ8LcTicKycjCg/xQLQq/NjGKpgsagHD928OaRD9S5ekXSBH0oZS4d
13pRzaJ5PZftNg8KfYonC/+w/sEdLBhXHqbmOg4CsNK3o6J7iHG/yt7HMnm6mt4T
nc9xROSKmkL8aUemq2rakLuB72zS7NKJ5hZFDbEXFQLGcZRlf/1icFebc8YeP6Te
3MFQrNTsZl9KU3jLnDI80CBQnS9+N1WDbw/sfqHeHrtAvhdj8WOwdvL5qxXBaPzp
iDbz5AP4zLqYERbefwgkbDeY/GN+WwA95co7FoNt0++ZXAYkAb79naeP6eY6Dl0L
+2qTI9oude3IOArbHaNpCAn98gwOHHUIQWoMbU+oU9zq4XwHobHsJqqnfnvkBd7b
afpvKEkwdM+aNBSdKwV6+Ai3B7zUQQNwzqAq2883msDY0TKMsb+rWdjHQqBj5KXW
snIZadTX2vx4uxpt9FgCy8nHQ4EnTXj0tyJbnIkH0EH09GpBC5Gw9YapqUQ3SIlH
yV+8fbZRIlrOdFrQsjbpk/ALQxcvr2V9jsh3nWIVrGI=
`protect END_PROTECTED
