`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rDot+abYEugZnndWXOnnVElvj16Nf7o9xfSg2rs11AU32R3kSFXG3prRiMl1/vY9
V05TEA4LUg5RvjtiL47XLubXEt5E7EdQPSMdPbxxGYaog0mSENT2nhEiFuHw9VX1
y0fZ7wgUjbBwwKKWwajablYVEeV4EXlwcLvmp/m3Siez3M+33Mnk9rWNyLYOMYNy
xiZKIjBG4m+HBsMlDjwzuljTnQ/iT3DAmZ/H+LewiGPdo80VkQXBwXARNLOYqvf1
8h9LPJoAnYGacfEW+ZhwhCxPfh6qjkgsvRGpmLfGSuwOThg4YTKenZ5Mb9jL02RY
nxfdnrRNk3dRojXcZaAyRziuzA39K7DJII2/Nv2bA/3i9Run9k/cX2v1jOj+N4cX
NmwnIjFoqfOfJqzCU9CbbTeomRZqBoEVbF8nW8m7VslRmsvoifHSqZ4/pqhyP0DE
cOVhEq/G/7cwKSSl/YMnumXTnHaoRVNFvlYe1CcFeypudh6fF+IR/dYlizXyl73B
Lgrg07zg7Su8nU8Sc1C/U21HO+QwOXCs2fbf3LSAPDR4EuSjVMfy+vcNzM1uwTyQ
SbVqYEafDv3y0rfzWPggemH91LSGRJBG3BFG15VFYVLxaDomqqNkk71A3flLYRqP
gKo5zM94Kb5jNehk3ObTbSgG2hUrpRaMmWbNaQWibaSiXvFMFjj+kkxOgnXOZYjJ
t/QaLDO/+I+hhI3Kcx+e7b3u52Jg6ZlEgvrl+rlbvZL2OMRBnCNJYBC154lviMZU
QewFdnhF/lXNY9N40WYGA0tkRkbH7IdHSP1dir0WXKPdDSdIEd7+e60IBbjX9XGY
+apgXZHB8TAd1zGitePOn3M0UJauNTLmXs4rNzGS9dukA9SghBwGhsGcNack1cr9
bMWuZC/v8KaRPk32Vcc5lcVM8DNRSePfjknxXrLO0YWtkj0HiDUJklWCYZfM+Eqh
gMg1BJhRlcscuqonR2omRsIwibOiK9nlPwLqhCH4IiRYl0t0Um9JGYZo4nG9EMYz
xFSPRvXWpG/XN0si3zSgUEwH1P0kfn78te5IVdTxfSvCwE3d0qQJi58wpsyIVgwO
PexYMZEaw8Vdo+Wy2G8NtMZG1Tr1bGchhsh3kPZdN8IB39KS07BX6uNDg2NJneRa
9KIpKkZLrxf17MBKSSr6bFkDaBARdztVbYiBEXQzEmdysAf0/skA+VbFCFEyjQah
DQOnYeOSIojZ5gGFhPz9dev+mWpcvCVynbgcoxdaIKeYanmI8ZiOPzsEYoBFyE4i
qRnUhRPlyJvoX0iBlXW8S7EwOixDpu6a09lnXHbxVXK6qMfrivco2ZvThIxlj1pM
MUk+hAJU+vukklKMEq1l4qcaC9j7FC7iRxqNJ0EUKYRHlbIhVsY3J3asrGYJiNt+
USzN/GSJVROLTSe+d08dgc79AasxgtTxcI33Syw/HYBcZ+lKwDdpWuFjh4fhYiue
tuePMD/0hhxnKIdM6rhadU56cQSfP/O15kj4u3oOYEuZEGOTOwO+Y3jy1FD6B4Gx
ZNXA5Wum26xuFkZ81zCqIq9n8ah4LCyeEQEgBZ/rLWOdVv1KLbc/Da4MGRUMrVDB
FvFbc/FApSxW55Db+ok2egCrz/w4dwelxUB6futvqrqVH2YNUY3e7WN2SsTxYd6G
zpxEfMFFD3RKXrj4D18MmocA5VKEXuBhNvvXnjfwpnWbpxMR8NOXeHRgiRmXGGn5
KreCcN1/QeBKd28R362foLhYnNTZGmDWw8f1tvbaxXmxShmLyFSt3TpukxvsLdT8
j78tT20d+HmGGUVxXJqVbQ/d0rK2HyVGtqTmYYYAMuhlY6vvWjApROSE+IjsS7Qj
yxLims4CJ0drrr3yMx+oh0bTUIZjiL7oDnii29ic6WnRg9bE/iMY+zrd1Of5Opwp
1PNT9FV6o8bF1u/48TLyw2slWzoYdBZ6bO09BsJac8LotBA2yZ8LiLNlSUrLD9xN
KRk29XSDLAgPmqPt/xGFZojAfB5xDBFbrij5W1OoWSagyt67UD0mW9NcrDvS5gEO
Z07mYdfU8+6y9wqRYd4VmzMd01qURSifUutgyxZ2aEsieRWS7c6qCrVMfyaQgrAY
QVD672bZz4RB/4BPwrtm76MEAHAt0iHMUCIZN+ADSqeV+cNqc1POpVEgilvMtXJw
Odkyail9lYEPe6md4o4+soU7BqF77Ooaq157IKhG2SSZk9GcLvpyA12Igtmkh0a4
0K0aJOHPmneV2b1cSGi7qBulyzKahXioe6ASzhos/GUSe4Cv5YU83RvjzRKyjBVM
7fAIrH6AApCZl3ThucpHNlLBpCwEMp0NdP2hpo7bdWtP6YnDIjro604GPcRHwJF8
LNg8dxIrudcnrCO1D0XkyIG1kubIEaQ+vUH3uR9vsx4VifUtDIryrCcENWGoYOkA
EM4ajPbIwpGl+ORy8mnhRZ1FU9FLaFmC2ZR6FknOCUjAlKCEHqVWAVsKt7NFxxkS
8X2iUODrfOIMZsGbMvTO6mDJBNZo3pLH4wAftGruDIJfvFpcjE+wlF7Nx1CwCFSH
m0Mic8ESSdwiYH80BQl5wQ==
`protect END_PROTECTED
