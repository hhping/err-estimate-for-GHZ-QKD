`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5jLxLebg6gYI7p4tsBbj9Kz4WVw8aeodsMit1dOzGvMKsToHnykXsuL/Uk64f6/V
p3jP9tlVJVp1WQTfJoZN3dHAKbaLg74cmKZWqHdpEVuBKQTXZMKBbFGW7M2ZH2Wn
W1kDhAHNJ0rilLiOYgyhjhpWAYh4FOwRe2C6Qwpolmnb42VXrF+vdIHgIE2xNg7F
HcYzYEwrWXTVXO2qC+9O4IHC6a5tSiCe1FkNy89oAarZvKWtUSCBZdHNTCGsaTFu
U1ucS6JkGP8KT8bk2nRiyZPjCCqS+azvOfAL6FnbCS8igB46xya3pXCxWS0rjukH
jIO4BO7mnfzt4pTQ44IqvfD2mWZ0K/JLziAv7dVceNwvkqMFCz/ZwPchyjr8v/d1
jy0DLesCH/7en0d+uEaMm7yyJXTD6dBUHLF+1EnZ5ouxLdDml0yYhzo6oQr0bEt2
oloJHqUdsywp7T2DMLy2mwMFQsM9wI/Dwp3V/xNLm3Auz10RpEsvKZdleHfLC2LY
gmR9CVbaeobTFlmvY4pHytOUewWj4EPf7hkxnrdhBaE/Ac7z6PLEdQu529viFJFY
q3dzdHYai1k0I0Ks9GkFOax+lkw4/ouGTNUEI7YB4D58cXqf0s+tfI4wNVs9pYhk
tSz8odP7+9ArGXbm9TLBGA5mSaLJ8pGqksVkG2MmVdNSWiMpynmyFBITDQxgM4Ry
qRGkkAeNpLiw7PxbKHaN84XxcZnpKcOxJ81XCYys/AA3ggR1ym0Y/yO+eZ2DRaeW
hCqqOlRIwy80Jv/eVquyI5JNmXyDDBKo/F8Ic6nNWE0+D+eWq8oQMSJQoc8P1a0E
/WrXIDJxlbLONyCDuznbXNO3+dBem0JV6arjk3B/RoZvR3SvClLpehZUJbl7NSsI
EAPAGBYikS6c/0MTtNpPbWSSM2ZD68Jj23I1ynOrT7aA367HPLHVHvqHrK9BcK6i
iBlPf2NDkZQKlqjHAiauhNmCpgZPvWWLRcmPtelHJYTdakEL0zwV2kKOChyiTOlm
jf+LSiXiAmL09wFmOtTEWwVBIdw8dC70VoZgXuN23gwm84mot8jpEmRsgtkFA3CH
u5ii0WfusCRdJ0/0Vy3gy8ofOITHiKtvYu1SuI7HRF+wwwceG9Y01jgusfff5eY/
OwJTJoCV8hqvPZvYiC+KQEpwwGCrrndv0HOmjcELvjqfXhARnJV9AYRNYzzGB3f5
WZkg9Yx14rSKJkZSI7sYLi4hMLbNsR4/CZWcImKl6fv0VVhBzxFPwx9ShUhZKBhB
wq4mh5KjPY8CcgOuyPY11NIZIOT+ueA10pMqX8qCz5LFtx6kIvxh8OaTZDGfNMyO
`protect END_PROTECTED
