`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGHSU7nIngAqUiwpOHzxnj6lPLGqpaubfLBjZrg0duRynhzRZY6guuTF+p8H7ASI
oGHKzwbP+tqOwBVri7xm8dR3gM6mZ8neToXy9Y5dXSZMo6fcoUDzU7zIfpYGcyAP
QjowM8f62koPl6xR41jBGj21FOvHFKOPBU4XBrskahRcb4ZU0HLy8EHSS807Ax46
ZXSaLfNvR49i/IqNr7NmD5Q2OALPzAWenCIGaU201YPlwaoj2Lt3dmW9e0eYwS6u
CJVxsgDd9StNoKRdShTPJKOm4i5g9cw85CmF7p2LkNDlkea9uX7PvRM+x8CignlP
TVtGSbNcYOTWQekDOdMKZIRC85WC6urW3lml4foX+2H8l78E/orVf+Dro8F5XxQg
LeZci2rcbbc69UTnuR2zxIK3UpULZM+I5Wjn/jVVDCHpbzTn0TushYpixvvTyQW1
bo2PXd7F145SHOHhhkhBcK3ygI5STFODMU9nhCryEZpId9vc/Cwe67sVtnCyF4nf
TTu794TkesVLbAoskedDWq4JYe9owrrJ7kgKnXq642LExcuyUxNfG23z+4ZAeKeb
ticVZVGFNcq3y6XP2O9jeLJsg+NqZeX1E1HdA9f0e+XcmU3wHr+HFaWegYexX8/4
HNEggvvq0AqQntcE63lMyx7qTmYhwTt/UoPpC67bFEQpc7pYWpV2ibSD/XL3JofQ
svDmjjkmZ2WtR6UdUhrliFFXaj1VUZFnzOxSztIPVCSeozg2QbBFx0Pya3Qqm38V
74g/UB86p+ejtO1Cg5LcjUdWNtSU8R7fIXL3FVAWmZTXeJ0DaAklGwwUUqvDLw8e
t7RIP5AD77L8twOlnxsybtHn/U0ZFPKcyuX1b+E4IOK03k8umztCbFcrm1Pd0k0X
vkYrEtYSrUrSACM8fbFJdrFRj0FqJlaOX2WR5/4YQ2gxgbHA53UPv5dW9al/5jfN
3ANaR9+m8W8VffpKC6YipfJqzF/BgAcTTlQIO0H9bCLAgu9z0TREJ0Cxbgd54vVL
8KDUqg/zDUtUq+dt5PNWY7yPHeGBQ5Inb3VwmWJ1SzPwBWB++m6Es7MmDvhG82d6
uh6UOxOAPKnyJTU9eiqZJALCuCz67SHT6idLqlNBFLRTNcGtGWAhcOuok9W82d1r
Xcs00izbL+FvJbsaMlZ2knjnRzTiX6nn9oCFMzFoHKlfruPXSXhJE7s27nZ2Bh/V
9wpoKVg2FapjKEozSAq/nOIOHveAVx9AFtyQPv2HTYJraGSTckz9PCkqZt5RYaYh
ckYOggkb0DIY6fd/fDYHw3WL1HK/YUFVzdiion+BlhEsKXZpBLdV/Ivnt0ZJ/H3X
35i68xFNP4sgb9jbIWPgc5Z5ljSXcM6ahH0KRSgS7BLzhXLBRqJXn/JpTUiNRdvU
Yln70Gn+aLW0gCkcnmCmH/AEyNVLAbMD6VKHH92pwiVSU3V/C7fbCXbHss1p5ydf
q2DzJFIyVznMy6YUdDFls2Teax+02x34jB74/tQ987r9t9eMv5mIy3manm6tjYDg
lLkW/GfXo8m2r0/nhjQhvwcM+pG/T2x93gdTflAjOUFFkmpM18r5cxa5q7rLy8KD
/Y3yGofeDVfeHqErxkp0De52X7YOjcDMJkzALmzeLNPEIfzL1qkIt8E7EVDvMJi1
rc/RuGHCnzfKKZVpOJ4JcG7kUwrxdLbIqlKEzMiCQKJSBY/esJTVSjxG9hJ5hM0w
Kj4FW8Sxch/CHeJajQtKEW107GE/g6N46ogeXZXuPRpuX2tEGLWU+FWR9D8Ns62P
IRJxMivmdzKI9M8PRm8mSEBVfwv7Dfs8p2Fvoh1AfNG56pcO1nrHdudKKh/dlttC
HyzupUkZdVHW8TOQryBF8zMTHx5W3PFey1C9ExGoRi6s27BHdFX/niN+AJgubYkE
xlJ6DMBfJlAoyyZuS4x8UQjc8IJF9k7uZTzegYrZrGGY+IbfqIs92lwqtQK/8dy2
bUO6F0lOC5Kb1RzIul8aMg6ZkZm6GpxRNIJ6hbw6/HaY4ZgzrGArbig1aoRpDSEL
laHIRmar+o1GLRutZ13ZjlIGUEacamOjIzrW0nF9yzqMhDk7zcFw8I4vThwGQFIa
W17TGq1cY+5U1QShej12e+UL0QXbCi9m2Phb4+QGMepDk68ej8YkSVbVvdSYiqsj
3aZfQz+zNUwZkK9bVSY3dbqyp+oblERwwAJPvUdRY3Xgu9oNaqJM/sAFK+aYMlIJ
hu4gjf5FtaGMNvC7fQY+nk8keLRzrjweqkOlPqRoyxVqVsZAgFRI1zspAtOvqyOL
yRpQ0Gr/NpoVNbdAFrsJKOBbvLkweRPxWgw7ttDavigOzDCrvyJmrqrZlnvKHv+S
QeJyCxDlzAv0A00LmdwTMpoZn/BOd17IE53Y41qWgiCVsRPmSjW1315TlsLyc8Qi
LwGQu3snHfjtboqlf7vtYg7dinzM+xv2LxMEf/Id0X265dh42U2P6cWky9ynskUu
P262YP3jDiZC9cIg+kgAWnJMjx7Hw83coRzB/PESF7tDbTku6hCs0Qyg/FvOjGKa
X7mhWIPSvV8FWdjITKCb4N2uS8fxrdjLhAtHRxDLL1W/3SkqJMQnbuUl6y6VgxCT
dK2WGL7D4Nkz+jF3/PihVix2hJe8pUS/ZtaqOBCeSrIrx04l3UEyEGqpjyAkQusm
pCSG+Ih9dNYX9bocpO6NqpcoZf5nxXffbue7JKLWWRHSg6lkHlcdJCwX+udglZnK
eGGFXf/3lN4ywwlLM6SS25ctUSM7dzkFXbPGROCE/kHqawGCbxQ99jqX6q3q1w64
P6JsD/e1wZUxTaBPIzCs29XrvzEMoo0ohgFTxd1rANmAWFv3knlUWLHb62AIf49d
XbvvKVS5W6OAAp06QdAQPlfrVGNVRs5IlEmMLryIS3CuKKNEL96120nu+QhMWSpH
dNLEZb0UDzoVI43WuRN6o1jycbMeLCn4zAuK/wU5NMBsYSgO7+pvRMelGfoErl28
b0BJ+pFp3uPo8fs+eiuK+Mqnk1zokEdcX6A61Bx/gshPhPFYPX8eh53UMAIQ1TzU
`protect END_PROTECTED
