`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRE7Pz2sLk8EefiQkU1QU0iQLe9KrMLHGYFh/ZcuTbv5IS8auaB/GB3DQTZH31HM
BThw5d3F1XIEYsqRXJa8cxem+frBt41PT9n66OlLfJLRMwVA0DfU845cNd3nrsM0
5CUVALzSjkvuwPKBWoEgiJXrYmgtmwgQVdRRWm4k+3/oZoZQdPjFYtGGT8UGFBVn
3WbmYyYxeVDqiaGXBUSsKRDkuGMi0sBrZLbx/q0odaNTxvqRYYDgssDuhnh0XURB
OxElmUBKNO0lL+ZZkyV407gR5qxrSHfGDaNlB+9JdoKd1J+uWuo2cStSNvPxn3lE
KxY/J+0bdZG0R5u16F2KBBiTZVpmxDLO3Y/6ISVFOjenXlyOAzT1e3NF7Rm4Lzf9
nszFO2mewQ1nFlqhXisIyeQv02/az2qXwFDS+gbRs+xvOt67l3pSQDPPKk6qcmFn
DEEnyYlxjOaGkK6eogBQwotHZMUBhnx42w1+s/YGg0Ai34Tp8f/wexJtG7eSFDEB
ihnvyvr1c+xpNpOSLa1rMLdI3FzwYpIVcsvBiTvuHx8LFgepRYI3NkURkUxY3xwP
mtJi6caSb28sCEAMHv5IriezxiiuIcSagTyc7l+E9aeMw8aHnhp8nJ3fE2ZihDJM
ARdPV4oWmQpFPiR7dHYq3uXKzL5sMYQaLo7tn6uFZgP+VZt9QY5M5CY7iQpQdB3t
MM7ohXZYAn4miyUBJutoeyxuwx0xdZo4JYYM8EuYmRBk7Y5r4HLNyd1ch7UP0RyI
BA/cuT5O+J87Hz/D9+irv/c6u+Iz9Tg4TNXQmMBp/ai5LQH4elgWBuCGw1oMSUQy
7xl3g0Q0r/Bxppj4k6WvBpzhSWaUXVFLp+u4gJJQhoxPwrYG7OCbS2y/ViuPF1Wh
LtHmjv6jcfxwriRuWcRJ6BmLMPYqKgznhrz5IqTvXvbQ+xN5puRAwI7r8j5+CVNh
Eo10YqW+sdrKzVj8+3dylrXI4hdbo/shivlreFgscx3+Rr+wRPuyX1QPcUkTxvB7
Lrdf3S3Ak9dxj9G0Up7izb0D19FwiZAauPhDQPdhDP9Ma7vELtjDiE8XC/LMH6qQ
pPjhuWROf3KK6RYCrvZ3t8+LfMaTjQe66rggcwbOvnGl4d/3ZrbBMXDSPJGnEaad
9D+OLV9SQqblnCosV5MOqK7zl3imadcxBKMR+wczMMqnZtA5w3gGuOTBjdRXO8B/
lmUJwOCcYgBukLro4nlDEt+UFA3kf5Hd6mWkYhoVXI2kzXHWH34FJ8H55BhEp5KY
iyqtZLQZvBbZVd1eGJ1HIZ2m4KgSzJaDn91gVs4hudvHwbWbJcLa1RHRDGB0P1Qx
h+ZaFKs9/hyX26eI8TlAyOg0TKaLYelFBf9Wx+A+c3vTzOjH3JKP1GfpsgEqF4lr
ttg7o7wStwyZtosGH2dXjA==
`protect END_PROTECTED
