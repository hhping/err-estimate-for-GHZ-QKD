`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kalkrd9UX5SOSBVbgUbCwQyTMpHefDf3XZMqGXX8rXgPWnHfRPVIJWAjE8ou0zFU
9usVKnvMYBSIKW6M2v2mLQuhtwAJhO5wijDXyoAqwfYftOUZvQwfIUEW7f38am1n
cEyJnbLAMPI2W0y+b87h2nKbYW57kX94pHVV0XecnHGOVh3vjQVowkGpV/mCsYwZ
DVNaZL9s9o75YY7m8oZV3n9ybrUvw9+i1Pd0IokrZGLzQSFUBr19y7ZCBDcGuXni
CsDpcltyLjBXBjBA5fUyNNVCICS6cbo8tFgIwJ9Gq4fnPuj/uU49Mf8lgprC/Zf2
CrWj0kFqqhtWiVmIkjGZHmwq4n+jDLsnPfHJQm3/ch/bIoGIQ9/TdLIEInqrrDVS
65bYt42C9xbFh3+l6f4ahicpV9hgKijkQZMhsmhWnV6WwDBalhzeavQvDZ/fqhMi
HiQkDm9FAZbJTbXAF89KFADSCeRUDnmOaa0vtiFr+eTrZ+CkpWoMTTVYlhLqGQpu
czGAr0KyQdYrfJZrxjinME7Hmur1pNDl+PhUSvMk4rBgT6wdVn5tY4XdaMX5f/+5
7MShI2mZ8CFTsWWIC+ufdL60wcdEdYSoR6kg1TMY9zeTEK0z5ZWJpLTNTMqJFuVj
Jl+fMbAcSr1QhnAkTSdFy6d3dxZimpRkU+ecIKdC+fWoI5eVyzuqcVRZASTGs+8a
kZADP4797Q3bSNlnE5IN67uG8JW0Nom/5RwSyxh7BrMuLWlKdCnDRDgK0bv42njV
dXei8p+5AMRzocJGvF+Syw16y1TnwEqavaa4jBoYYoFtpeng+Wr1J4ctGn/qXaXE
Tix/0OVIhnlCwqy1UZ/aYsBmC1lKDT3FfYWcmyVE96bncD9d56jBjwdOzOWnsuQi
VsQvKXby67JYa01PM3FAZRzDCJtX1iCc2+89so6nq6QkJhbU2/50Xnu+Pz8PYbRv
nIRX3Dk2N9GSyjj7pEVhd+9TUi3xPnJhYATn66TMqYAT98aNaBOyjG6xJVWVjpP3
ta8asXtYLL18qM7cAPQyx52EwY9K9Wp4EmlHZVHayrIvXHHBVyWxvDUvSjyQQ17F
1oOIjogRWDn4JiL3caWl9g9yAvcTAvO+0Fcb+0L0xBIZmQLUWZHKYft1rSY12tmW
ntii1mrtKuSmvsIW4RKmKD88bcecOQryC52YENfShSZzpK8dlOGkF/IBFWw2UCOm
jsjGwhwF2vvY0wWvirfKXmYoNmI0uZH8Xa4df4jP6ILZq3GF3OIOhPE1yZRxeeup
Q4xHE920qa6E4NkOQdHvVhIGIIEZ6V2cEXHoYJipP0b/Oj3kgymy6+6SoVmPEeuk
79WQbT7tBOBtxbYuoZZHbbgVOaBfL/n5VCtlb0bM+h0QVp5SmtMqMCEEHDzpWhZh
iVqOtqhWP7pCcUyfwMXG5zN5trFXu5MzMeZUhysOwSqQr1c9DOPnN16y8UfFnmar
9hIWqEgHM0sVzPz9f1AQiJVgvkKFSn7FUVPYCkeMV9VX2zPg0MnWXxO6VhQYfknU
8+wIhzMBDD+dH67xJWKLrnnRg7Wq68AFSI2SpXAm7mTWaX9K8Bhi4VZlOBLtBZJI
ns7OHNR81dcr2FawBEnuXle93tvZmbTBQdJ4C7SJ36QfUYmX0SZYJkKWxfKcPdRB
5g1Pg/XDD6Shs2JUp8/Ek/uKAApSQ3Gr0l/0ydDoDuyMwV+mmGvp7mqL7qehJD+y
hAXG+6PQCSf4XlkraHbDQDHlV0zMWoA54T0cjr2xo2+rMNjdXsYbB+mlw2aSoRtz
5GxGEMvz8FXSjyL+3q7KiM+myV6tjuiRl66G/t54Bod73XCvs58Gxdy7srWAHN3S
pZS9UOcTEca0bkkfVer3BXp/6wUhXGgZJ/HCf525Yd+nxJ4w+0OGWTnalR6mndi8
RZbXHTweqFmAByo/eT7yCHzgTqp+XWwvWGDJemb3w+M2ONQXi3DgZdATyLhU3Yq6
hm3Z7pKLHG4SG6cpk+sWvNlbBk2kqWv+h8PVVacT8Mav7oK0zkCzSuk72HnFG+md
Tp3RHAawnWLLEBwS3NL1NrhVrMnG4CF3ksu7EVQw3ppEhKsvgQzPbG+P2yq7Kl27
XSP4kKMPUbhP0f/3kHDuiZTBhLJHSBk13Pqn17c2n2FPR0qiw79wb8gc8hY2JllH
dCxbXNRczrqWtqAYllKAGO9rnCoveW3Xgen6YTkeCHU48jDvpYUFDMXhtX1toW/9
7Cn8OmKDT2akLWxpdZFuJl3YaJJ4WJvdhU8ezjqUpsBLvxSr9T9N9Osi4KzalfJo
P/Y9j9vBOkgH/yJYZxRKAzKEsATViAeyCU2uEzUe0uUt5mXzWaOdzNoSdm9JcORC
fgvzS6vtlP4+DFqM/idTIRE0t/eRIUKKReG8X9kwrwsnu4X2xqmEVwyxhc1XJUrl
eXLuyfyJraLNBw/K0jYw2K0zlrnEsNJDuMxjHgoYtJPd+M9jzdKum8hdS7n6Q9Gj
V9GDEtavzmM0+sezossMpQOl0NwNPlD3AxCndcT4HVqQfgTfcbfqV08wKkMvJtzW
AMiT2C/1prnQ+Mlg3CCUGHtK8FQSxiFaBdLjKy1gUx7qxL0rchbPP3d+wX8PlYFa
Xz9JcG5ilQLkhf4n8y7KZBPuE2D0QhPROflgOs1L6EJNUTFbxy7FLWemkZwxA9Ht
/dBa0QF9DW1at2eJ1Bt5Ysl6fs50cic27GcCN9a/iATVHyMA70CBzbXvicoqJJhs
A1Iw3LiXtz9YjGGPY+bVu6TDHwnYu0wR73w4GVVwZze1V7g34DsdhvvUdGbjR4ft
RB/t2rLFcdjLBBpLl5GExzDspSTCksA4AzIuY0zW3pVDx6ey1oA/Arl7bUOaYcKI
g4TPOQLAGPlB0TZY092h3I7DHZJopmdeCn9W9uNJABeXrO5OGFg7QMiHelQFCDy0
EyEVm3S/iTC4MaoNu5xhcX7dKuMmKnmmElU8CoEFFMThimTNXB9LEP0Z+dNWw+Mf
hoBECFIR/dolyhgaaejA9mMOgqknnWg2HWFWmdq4Pv6gnj6PxyZD7ZUtDUAVzNNr
MEFBzJewheygJRRgRqbjUMOT7GE6bx+oL9a6CMRuSm8OOFi7rsyIkLL1n1EpG3zM
97i5lqh1Zhz7UibxCKknNj/ZD2uJK+e7UFMlO8CHPxmBWBAMNY+0/cDJ9bH06/GC
dRB9Rb8Qbvz3olbve27PB/gAiQ/y0cYMcj3SYHsehYmPBJswnCi1oEWyGL0Ojyuu
OcOi8lWuzOrWdHGgpNYsgYQVnUo7BtwYXiNHU01WciYoVSYLN/QfpuQHcd/auSxq
Av67WQMjoU2Z4yuo6eOJjBnPxaLAwgSgZs1637sL638Xq8X6TpiwdnM0kO2WL5ul
+KDbK3FyGKEQoj6A37JRRb+M+bGbNtZs1GTlZE9ACHqQuq7tCofMxntPQg9tWTzt
mYJ6m1sFpcANXJGQ93PhFeDKIEZSFdkb0tkF92mrESDXLc+schI6qZwuXi4Zb2tQ
BFY3dd3k2KnDZiS8fCWEdRCx2QVlo40mZ1SOHZHxSqMWrmmR6AkR30IfAqKyaj+7
+tNFEnYxRHYkcMfBO8MVyXZTq+5nhqSGbN8F1objIw/vkKyNQqx6o/cl5c3OvbDL
pig+kpXuqBFHU7Jm3LSw0i1EbU9yuv/pkJeJmbrwq2fDC0W0cy+QliTbmYtVmrCH
tQHlsnMZXQC9BLCfkljQ1AfcnhrzhSXr/84wCEMY6Tsp94xdAn6nVUuundhDuKDg
Gkqmbes6MijUbBSikJj0V/ZM5BK8WSPZTWScTEK6Dtgg2/GGEAUxDPpvbQg71oN8
DNvuuhbW20WJEtmsGqzrZ2Hmqxn6/gT+lJ0wZHyqCRWLjKgWWtZce12J+0o77u3k
+IgKFc+pI0eo0oc6Adh6TDh9h+D0+tEekwdGDiVpz9n2w/OV63MQRwkxKcnjVcR1
KO7hLuiPwPtdsc5MYpGMvG3pGPzjcvYzxY+RrylBZWg/HwkShdQRmE5GLTTCEjRo
PfECGXT0HNF49qHducbQqd7dNxWeje7ek7+6YQ/dBo1MjU3mtXpKjk6EfXe3tIvc
jHFIe6IuHC+lXO/y2YWA6kxc6AQFNx2Dpr880hyN9kk4zCaNry3rgU1hPQ7+ZA/P
0cmWwn25sr5EeRxTrTUx2+Gp0U4f6W2q6GXMX0nF3eJrAO5LdLSVhdVaNkmafY3p
eI+vDNcjuOyYiF5LKfbAVE9/A7DjU1yw7BPW1y/kaOjObO9/+CYI7pC+Defr2IR5
LaQPGI27tSG04hlpS7psRc8HeEK4k5pF2z9iAjDVYYK7+tgnOk2yAlhfKbPYsdrj
l2NyOiRdpuWupiGcxy96wNdOJ5v5fZLqVUJGZog6yIdc5YTbiMeoGVVrNZJktxrT
bba0ihW1dBF/sIt07pjzk9ZgsraC0wSAfReJSfijqnaBfUhiBuDQ0z9FgEPpYJjD
EqBiEGyYOV+nQprJBrVW9hcSOXj/lnWEKQ3m0KPoyn78908d6M4tIeJO6D0hLSxl
UXjcy0M9Cm2ju/n/PsL5ICLDCZ3wbWKDGFySgVLZ97Cch2M58wya4pE5S2EpLF+G
IQ8MXxufNUpayGGab31cyJiRh32i1FjkjBSQkUsfJwiDEWWIxJCRXKnaCLAApp8F
g5FWE7fjAjsGPYln9UDrf09SVgtpw71sZGvWKMALCxoi+576/nZVJpn2Hed6ibXG
95yLeDVJeV0mCqqOiTaNts7+ckr10PXVBv/FQ3ZTpetd5iUBH2is/0KOzgryx5gy
lpw66JKbbFxLRzjphTPcYn2fYwycRokiyruvJGdoxpNKPxuj0YoV82bj4VpDUhoe
RmCFY8LDSODDNKyqvk6OQ2wJrAIFzSZBlzPYuuk5K23bB91B2URyaJPq9ErLujhO
GaJ5Zt6jekNvuvX4/7RfxVHNrOLDeTcl6U40MbN6pxLqA0DBuSc+v+zB3pZUYUaW
zDLu4AUoNog3c2n5HGmFRZ25RG8YAdeOmv5fuDRQ/t2EIxgjYtd73HEhF6ksvc/i
pyhB2222qpyrJjhnL6VukjrweBKiBCaDaHKYYH6lHMnVMkkk700NdmUQxE5DHchh
UtXI5wIvG+P3Xa4tCZ6emo6tPh7KZKgyfCn8ra75MW0l/K9SrzZm1MggZKUlSotp
SAB6mImU0Gbm04N3FFNG0tOzW82BcYv9DDD7JXZlClBz7RXpSlMv2Ruv0+3PxNzb
XHqbCqJuuygzhewabGOTOyqZ0k1NkTXpPKeL3d6bpno252HGPKC3ILwyQiqgllE/
bBVeFhn3Ib9okbnDBnwDXUAYKzRHYfSC0+vxKdcvrg/LMJBr94qQyi2pxtszEPcX
gyo2o4dsWNX2TDmjY4+0wvJBEZLkbdXGWpZJGA4K4eV7lJUqWvyXdQn8Dpo5Sc0c
CD0480Fj0TSFIfco2JXM7raD/0jKF88RCiBEhDxrmRIgBRcg9FFxgqHCmfoxzJb3
QZcnpGTjbsFsaYVaTdR253+wzA/9C4BLQFB1FckT2l+sVKS+5Hy80xuVMa8ckzoN
U25ZCjG4pMRFRftGNkvxROxbWULxrJikWRION4MEksm0T0Y4VR/DUXzGU5EN30Y+
Zg0XwfVPlGZisEUMNZ5PbDfDaJ7qzZi19GxgCKAys/axlG/ReOfuQ4FFtLM6HEus
CZLVB0R6tTDRjS3Y/UH7OLkCaGGcobIYssHP5wjMJfqOgdKsbXB8r3OA/9tFY0A0
CQBWcX22owh6vL+UhafGn0cBlZQiDUIOWAwOjLTKKHoXYu397psDmsEx/DbWAIdT
z1l/30CZ8p9tBTAVwD4L8DZ9x4bzWZFTllrPhNV1fJuf7UTcD6pnTHe4m4cRHJge
llObCZJp8q6YZ/U0VJpyZeMlc1BJkFXbY/l+0amtFfwZirIYq6vw0DVZh4mBgjLA
WYFausjsy4SWNTy04FbuaX+WfQxNBIUxiFwU6eaFuKXEoqLxNWA8Cew0dOUJY4yR
RGiomZCYftpgoIDJdCvI4xVgCDc2dUps/rYMG7LEagx43dKBYd+sgqEPTBdbrm6Y
q5EX/7gqXk8UBScaxCBw3EhG/1CosK6U8+b+SCvoCa272gKBY6XEC4bbbJz/RHJn
Rf8HNjrSbpyOVr8Zh2oXrxIfJf2Y+UgUjq3lt1X8tU++jIcZNILr9BDn9/6r7/lr
dwqv22fg8t2Lm1u7c1ZZJdwxeKVIihVSdiryLP4Ic6a/H8MK9CLqzh15sxKfnp7H
6Afbse2JIFHZPiQyTS5OxvZRR/o9fJajL4TPhJzNANKV+CCBvKYZaCaYMKXxQnwJ
7w6Pn4CiCO697WSEnjAwGML3qnJGUHAZJIFxRbtwBNUEZN/oiP+rjSUYmplo1avf
CNoF9cKwS/h5X30vSURNO0OTTyEGL3JuTCV3n6vpsrSCMiIG/cOyfWXQtjPARap9
fcWQhQSgcDmE2mxef0G6JxwfRTfafVuE0EdMmuUKCUHiF+h52cZc+1mmJyd2B2uG
778LtiFDKLWUfkRPJ+cPYhvWj04cCoVhGSYpLwFQ56M/OXiBCIY9hbDb9zGojUBn
6AieeYubeAoyEAnCT4zXKsw7pwcAp6CTpbvJU3YPb64xcgIN3UgMIQW6VOHggo49
W18svyc3zuhJBx1qkvpremkGJOExk3uTqcKM2WAbUnwkniBkN3iGOf6bb62c0U4v
XFxQDm2LcN2xOSOnaV2XSWU4qCA/qpHFgv+yMFwog6QB9EWGFF6M4FppL19kvO+M
+1xOB7xbOHLMfau/CY1XcOxYSkeGj6YI3rxjF86BeJEu/Ialvi7FGLI+9ZZKSzfU
ZVw5K1NcdbVh45+Ofu9DSw859lLByMMwfFPG7tOnzxQYiQwODBBARxDk/FXliRB2
2BYNLfPLwKsSGLKdCDr5pU+3XyjoCq4KQ3rOD1qnmQbANTgCE17NSX1SgXgwT2z+
jECRWJawje4BarMdZ+W1f4tVfeIQGKtRlmZYwR/RKciGCxUQyWAUZdcg6aWIaeEI
ycptANjg6o3/WF10bn5iR/vOF7ZTXzpZSh46sqGwQ2QW/Dn52L1McW8GxBhOZut5
W4r9U2aHMna9TdxhISWfB7bonsW3+xnBwpSBwTBP5nFRUcAx1KPgQQkRDdXllLcs
GkJDz8sRwjJjnMrnxIwZq/OoVgWggxjYAPQpKNU9mNY2lxZCLolqyCXCTpsTSPY6
Nav8S9rPhHSFAlbsCx9PRvEDiKjSp0jnQBRx5vmF3euwt665TSI2xQy09NttLXpR
pRINPPbajlqD0NMCnD2bI68CzZzAsJH1XXPPafl9WGtWWF1NfO9TXFlLtPFAKSF6
JD491R90Zhmw0HxgYqvhZR2sCLfyGgaBT+Ku3gtg2xvc3RdPDVxupz+MfUhctT79
hQPXuWLdZGZmPoqqGog134qZWmEW4UEb0n2mWHuWKdNM/3U7xj/DIBhARFCFM2Ke
mSEHu8pYFpnXlfldce38Gl55aQmjHamvVTw9aQ679bDLTRDjIYa/xs8LS00kyGKK
cUvIcyPHk8fjny1fA+NYJrSf7Zopyap62zVVnZlQfZJqRQNngpixdMJLwUKiN8Z8
P7oibPtWxXeCyshvgYUE5dMNjCSVTipBffU0P330GXUb4vrh476O+C1pDsAz/YTH
EnzkQmTIWd3EogBFW/k91LxYOBYpUatgNQgWuLg0CShZXKL/GXarX8/McrtTIdZX
OAyaAuO7SUiXrroeXvGZ6gjfr2M7DgW3UWTiHq2RHvuQRHCM6T+bpgRz02ow/9ND
8lqT7I78E0lIL3GmpU6+2Narcgm4u5Oymg9DGroW9XmvtsIK+fZQe0I6OeUaHYdk
OYzXDtOa6Jr0E5IpNwhucrVTjFnQkFpa9ibzuswKy4iWVwsoEq3gz3FKU16nDnKO
PP9ugt6jEhtiJrp+Gcet8Ulk4UO2828l4I+jwK+NAEoejZZSTZDyg9H1S50bzt+l
yW2gbq4Am89PQ6Wh1W1EdMBWgawhv4n15lle3oeBFGwgojPqKur2TxNqqNV29mK2
OEiTgQ8kBRGyL6xZdCIQ78R2ctQCrEF8QmdbP3m4GGiySxHi2BUIbnSex1yIxPu8
jL7eSuNdZECAilp1W7inMeX4vmqZfSucgm+D2B9APpz9+WRx0x4oel/TOcHiBgKl
v8W1PuNxRnVBN4wzRgA6qi0F3FOe6Faoz/bcsKu+L+B/RWOAZyd1othN1XI/gr4H
jotdsmOxCxJU8hVsn7DmzLIPgY0ihk+hb7Nvbci2aqRl4VrJ/87cOpzAi4AidUwa
V3o11bKMagDOKINMSEd1ztT+i+S7lB4L4VS8xi295Hq7xZ1As0kVackRP/w32szz
tqlPIdX3/hE+afbukmsqnFKBQfisitMPlm96TTQqC3PMN20JrFRCf8AFQJJyIxwl
AotlUTxSAqDCqO+M88fCosJz8UMAfF125NDsmg198sWyyrLjX4u350hEUiYcKBbM
wUV7fzWWUp6nC91XQclpFbtDzPzy/aqcJOM6k7ba1Uh+2JX3wr+NFp3mgBO9hv5F
Sq8L+dDnQpoEPORRZFG/3k2YGK1Fe3iBJ2JpkkapGQh07tAEQKi/YHOycySaYpKl
4OkuOoeJaGb+L46AS49FnLoPMDdfzx0vWJQZC2Z5U/4H4RYZnN5beaOIO4RIoLJQ
Z6h0gpZGuZG1vxBSC0QTndr2jrTlIM3A9UE2rgo/sZklRSrCrb9CNwMFd8NzjMfE
Vn9oRzCeH+MbRWmlquZ8PEt1Wuz7vdr4III2ahdoAVWuaYzgsqqbNlD4SM51Ftpb
+kcZhTXgSit1+5Tg8zAJLmPmap+H+WZ+05EeqfCm6gM2pPjtDkyBlrbwgYaVP3ZM
/TQFfUILoXtSVyR/3KqxLzjJJontJW3mc9LgxA8wjSs491MqNXWp4J0X3qFlxfEJ
wGQGW51u52fVh1AP5+U56gn49SrsTIo/TRzb6oTmMJECCl+EN+Hdlpudge9a8ic/
nHjds+ad5GYuacy/4A7r1fAYpuUp8wumukndmX5rJRQC0IIlztFdJi4NYbq4/sBK
kGl1txvyfEbou9T/4XMZKDL2HbNvRkiHyIUAv3DACJWnl8c4nxb1UigMlCS6bn1y
wtdhvoX/fUE1QCNj5p4z5iJTz6rpzvM6Xc3FJibVXzgphTUcp5Olcjur30dQ87lq
O7S3PsE9sLKCyUjyWmrNUsUj5RI1Q9w7UyvQlcUPPGx6NaC7qLj3Vqgu7ITq/ce6
i+dlOlJLDslYAwcGjrldaMoQ7P4IU7O8j6kjLVMn6lqjwD1JopKGix2qTl+asM9U
f/R4Pa6EyPE1U/LDfjO20WA1Ovattue9B9CupzBxmjGmZMSKgo/L2DkuYOR8Xx6P
6k6aPuCmcyj44IBb6V1yDkazGkSMC3AJ9BfqHerbd2ctVj8EsFlGLVf9Mz/Gi7su
IPVcSjzF3GYa6fm4wVYCfN548bodbD98iL5w2fxFwYxGu0UIuBovGe+PWuTo91OT
6vaWEYYvlkm/Bha8MRb4iNTugX2A0Cb199oo9ux7RutiZcYFz/vq+nxgALrnE3N+
BJgwRvILhz3TJQNEXHvjpv+f3IvoHK9k11cEzWKTS5xQ2bRE7h1u66kq+dDGr+mI
GIzI/ze15ytqyAx10IU9RmrpPDvkthwSxj1vcXOjSVf3NjFwDGMo4t3Qmasj8rLi
igO10fKijXKLcafrW4sgPmg1tMhDxdMBBeNUi+WK3JQidTSL8xVKO043OiHcBe+d
/i1qs//vxoRX9NlPGEJu73l/7yeautLF8snlsvpvACErtIIw4YgMp4hFe3TYIOnj
uXvm02JhnDaSNr/vWQBUG4x4xZTtAV9A669bXNjfosEKFP9BFEsXUIAvO7JHppOR
P9kT6ksYb4q8Bplwt7YllnqXe9LjWwM/In6zIOJBYqAWVcuuAcIQPgaUnOabS2kY
UWG3MYm9eZYZ8hjaBvPXoL0zLQ3WBMlWC/R07YGfpKR1osa0zHa+lRD+b9Tkl2ou
cl4En0wQRwfFvHTiEyv+ozTbl2Jx5MZttN131vCm9IWzi3wrddnu30yvX1QrVcNa
CGVENOW62a9uT2XnWhB4Ys0v9aazKffVb3WdTiy5bJ9QH/rnudxbnR1V8h5I3ylk
mpEXXQzr9XDg5HR9w0JzdiahVjCFCyHgTRyHZUqnVcExGgIwu1crGJUOgXpmDDJ7
3ZHPlXc7kOo5fCDLdb9eewINiIxqgoQYhzfmHvUMmKjMI8Bg5oWHDBXDTFWaQBbJ
KXLuUyux9cpktvmRN+NS39ebv8IEc/a5RrcKhqLMFdHzPG9/+iwD1e1yzO5Tn1IA
wwfRGmFAZKFPnt/cqtYheufh40e3Icbe724INGs6G73joS1YQSrAg+N0GsFARcGq
lysJ0ark4p8RNC/9sQjQFyRhEwYQXeIZZRwsKxykmAUcTJ2XkapoDCjPE4tafwlt
ece71m3ZH/qkD5/eM+Lk2gDrebHfT+DVxxXRFl8YEVNI7Tm3EaWHhdj/mPObJtnu
Wj22MfmPMKG3K/v+ZywTfMZZE8vg6SjYiqhwJDSSyWlEqXx00diCKgj9Sx3wCeQf
4tzvBkV0hrUALQFkXndBXXMqLU4+nuu2qwVb2ac++CRxUsTIXuxf+8NjVbXlEI3j
/04U8WWOCExX8JBefZbvjVokBeh2MQNeoDxf0LRn/dSOx8t3vRyWcAFmnOmYt/Ku
S8RNMTPJQ3sCapq67jwJxuFt5+MB4SAclIHkJmplfUUdT74W9qdGlZ+COA9E2Lu7
YyVshaqLmTV5p1nWvHe7O1XC424XmgCoK7dt2+ca6pyVugSM88dL0BJGjPvOrd6n
f3Fj/CoRnxm31s7zSnaD+xxRFm76QDO+DZfTKbOj26dq4jYoPpANlJevYeUtCyO0
kQg6BSJRTlTuXiZfWUa4X5MSTlYSLgAQi2ztAgCveAfoLFF6EwfMh+WqbthGw7xW
7zYSW6KZYR2QZOzEoKy8KRWYXQaPDQtPje7NUvUVVKk/meY3WE3dduKljFx3JTl0
nFYDCmelCAhcnLlaFjCvFdqI+kjHlontHjQDOjE/zVUFMxo+4kIARLjeYmtyts2g
XF9Y7FSSQW3buM1Bqy0QoC3Zygau4kvZR8+OCeXubKWBIO0ADEV5pW6YqXb4aVEU
mRyCGT+vwnjpYhnscnkZQrZCxmoVtNBbWWg39ORVX9UtFup+7+sRLa+OalLg6MEx
cZZ0WbjOEC7fvxKGZMaDiCYxrLA+BQxFk92Gul+edW7BVPYYV/rsDecy0sf7p3z9
RD4D/NVbvZHiZFrzogRiitl94EiOvOURzgvPhRxEQRDGhRWp17NSJh2ubaIchMN7
X9L3p98yN/OxKqZJ9OqfuvRS6/LneID6FaLyO/QWRNRXSwrVv+swq5KW13togHNq
0CYaY/m2AT6Ezej0sUC3e/zI773UX8g+6J5De5iGAbkbnRU+yp79zI650rpHHQYU
PvFSoz9FQ9q1GvNzfZiHyLoivH/7d9biYVIsupJBhuXGgiQ0MdKRMtIMShWA6cpM
pwRBCVM52aKEJsulWzbUso8Sn8CvAFqoyHzRJASTaHAt6/8U0474ypLEHCZRXyCQ
wjTPAaccBI0K23eTvT9BLw5pKigIaGt/kB5q9YG9JIaC2PvGMgVwhYvSDOQXQfvY
XENkhIx/bySgQ/e2OoDxEDozyoQwuvp7OdawPqBvLr/5pZiCBCBfzyC3Vb7WspAA
1FP2EfVunG2s8xyfqe8RgiJ9eKdyvkGXGcQ3S+kelrHpm4VwZ2jJ1xvgsvXUeGfq
73GV/xcUYXvQE7heDCwbyCQqczWzUlbcQatClXGFyRAIEqKyj0f0FKn6BjJTCSAx
GLDHJHInnpm5YRAGvSGtJfRXZDH9ZXhDDpD2A9iJhsknoJXjR8rqcbwssnpw7h1n
s3z7SYd/SFTG/ACFfNZOvW2gFxBe7E0B21pFBa0Fm6dPsxjY+Eu0WQyfMCp+8gGw
aLjj2JCk6+YeHZaAJsrJ5tBa1Kg4gMnjuRLLnNseizh3DK34f0XYeg/kzZ0IaX0Z
u8QZ41a83MWdX1VY2sYIUyr/BcIPXjvq3EPjWUD4B2yPnV+5pzI0CcggFsaXH05Z
XV+dSRvbH0rIzWZdkyvWQuPVQ1QHYFqKLm1LLvMMUowJhjbJgLw7yrGdPDpHVT8U
d6BHT6Bf6FAVrzVRamI8U1L1cDUbDk3mU66sqnaYRv4Uf32oQ1Cyq3fvmGjl1VJ4
9AwqNPrIFB6mHi2oTVWxsVZqYIP/LOeDJB0pK6bLmgHjkI2kDvu3RkcMjiKGrIW4
cqK4iFICBUuCblY1wXcNWWIRHR1jn/cRxTv7wj+U5LzlBeWTy7LVvOoU86VhptxJ
PgFceJHCGKGl5CvyGdtJ3Ax+CgUty12dTAHjvpXm2xOTEFlRScsqimuQH4E99gUi
dRuMsPWMwBERR6A5Cpfflt2h1wBv/unFyKSmPWxhlAsq/HFT/UThgnsT6b1ROG9/
1SUpnFMgfdCpZnxklZdoxPm7w6dww/sS+11kNoquxy4LphqjxBvzePW0mJbci4Ev
m4WuYJc7G/1a3srGsvXk0XAhoprNi+Vnbl43VnkcfptyCDL5MefNNCsTF70VMhcc
d2MRfAnJ5WIvUPFYlL/fc9ocng64UxcF0amUZamTf+y46tsWXxONNJ0thocR4a28
MIlCqXS4iZmu2iFkMZFwsq9Q/qLEjKSjimtnjCqBWqSQEtf5IMkXe7Dh54IwpKMk
tYO4GvASUHJARnZdddDHJTKyPpfYugZ3KRsEs2HmZwamH1iQOuG7R8VrjmmGHB8T
8pG6GWMeS18A2qM0bBZatvdJGYZ99UgcG/KF1jnNhZ5UIDKIn0KNNnQkQX7fBZYy
cKm2afPAf48zWPrLSoeH2+hD2zGWQjAAd5RyWi79MQRh3ZHmKrSjzGBFqypcl1JE
CA9o+iEf+Nkg2QHJrsW5p1MLFEXH9NGglKpL/62A8yjTm83MbYbON9JQo0TSSJI8
TcnUsgXkffwcpj8ycwsNU3ARzadYAAzhiLiQNLUGqkTAWl7TX4VrD5GDocUiPBYO
r2ThpRRCbMMgL7d7E5uowWGF86By75TwfZ1Sge97U/c4FAAxG7XruQZEFTKaOf6q
ho72xGvDfSwTTOsKrUIbIzAHiQXCP9BMddK0vla5+YO/KPfxuELnX4fadS6JxlOG
I/hIp170LZIHACBMe+fkWUtsSOr6eWK/id8c2kDeBXlFj8lNEQm2NBWOFHLnqYcV
x0m1T3DxhtwXBQmj+6w0hfo5W5GbJd8UXLelj1KngxlKfFa4TyqT8Nkb33V/Ucip
xLD4e1rzD08tWrm9pCfhWL0L8WCkJvPiVGFRUTORqO3WDuOlnADvnZhFEdDQWVDZ
Nq5S5ci8vpVQ4+U1E48VdGv3zQL6j8tGudm0S8kMR+rMHhfZKX48BdJENqZzB954
AW21UiL8ivRk73H5iihx1lfVzLL3TUsc57VUNqf2zQcTB37S11FmfiTnEvYR0Kp6
GH0CME9WnHn76VcbpeZqY0uPFZGG/KQ9H+bUdGydOgvQCQlT/7GJz7FrZHWviUmt
K6AD9ucMZ6mfNBwmLRRG9yUEjFSzo0oFKdbdA4rOL2jXJu2aKpzHblZxkmV6uQwN
eKS6jas+AycJmsp1Nel9yILrcH3AZ2YKjr2HTm2Fg+1wTbcOC2xxJxiaFgZhYtFi
yOpukkx0y/8z4LSgxd8KQ3OkYh9ozelemmVtG4svp4MiNw9cXS6fnHWEEv2Oyv/1
ECY62agRBBg3Ijo3KQ69bPH0MejA3hpNjBkfE5pGRQAabMcpWo+ro653L4axqdmk
jZ6+VaNezkRxPBz0nzpk+6UQGhF0DKx7gseT7UwmIDY7e3mpjWDOLoXNMw4I4ww8
XV2ppWGrUbP3w53HM1ElpuMSON0sx/1O75xpywC7OA1KPzvuYscZFK25Rn4oBSKX
okDo9sj1Hl4pBbso+5aelAhM7SmcLTVvqLDYW8Ww7uRuNsadhvzACO8kHkgjGWWo
L9Cf7PBJIenbvFpQM0T8jxAM/7XOiu6syBRuyfwmRAlI6/RevjRFfurKqim7JR8c
APoZZ6e8TVigRxKJ1agtiCzWmoKMo7JdK01Y2JUb8uq4yYRtieAS9HjFypYcV3iE
OLM1onGMOE6v+5ct+OWo651PCGWCU3m+Bvrj2ZrtBjlszm+REgFgE9iDxuK9+om4
TBefmcnK7hDRpQmw+ckC0Vtt7w0wn+3QkTV09LQa5N6cdNBWPotqE+wcAxazjvPI
LCheqvdXhG5pbHUkjATQ2WbcA2XEk2qJA+XJJbLbRf2qE8CfKaT4/cc4iDVv80rx
8jTypMd89J75BIhsUF+NyH0CkKjLbEKInt5guiDakN2e6MLYJug/veBb8swsNJpS
o40O61/SUGcyn/I0L1QGh8GZrmtZa0Vob7WXzYBwm7I36XleCbCTWvT3rHP8ln7I
Z6ID+nAsPgxXY1mnLQd9k+Z497RIrEWxP8hC1QYDWjtd37dpkfKR+IbHvODGXHSC
taIqrgor7wRt+Gl+Y6assuldyVWVMdUQ78OygO/fMBkLY4dSlb7j9ZNFWJcoonPR
PMc/8Q4m/0tt9MtF17zVMExGNDYJQ01330WZqkpjTlVI+E80uDCj8YfCNaPg99Gj
eVOiY4WT6ywzQJPrrO430JTLhHbSAyWQRsJqrACgkM/Ctn3SFiHjGEsbCXyNp9P+
/jrdwMdUU+XlLzSkPSaHpWy00hkHhrwc71avTbYDxKk3VzLIfsexgSw6BMxijZ/M
f7zBtAGN2YTaroap0LQfrUN6Y1DK/njY2b6HYkFZ3uB+Y9dCaxbNZKFXoR46h0W0
xlxkBi7zOIFkut/pI+OrgZSbakWz0g/B9fnJc6bq+QJ2OuIRv7v1/IdvBEm4NRT7
VZtV07ZWmVCkipyeCu8A7/EJBNCiZi++/wMRBCs+BlB0QJc4L95JfKs7gZz13UbO
CaLClNsL2oKmTORWw9V5Pb7ORUIEfR6JIXI7otp9gKWwS4+iUoXuFPkk3/UgyVrH
qG8OrRuzzpaT9lbTeqnrF6f6fOISmQVmXsaHBLO3bKMtqSg3kKzMaD9Lir+iu6Yl
L7KB/rd1TMulLbBPYkefiCmLkm3VBjSmMBauVitp5YA8tiSus+ONgxt5kTW22aEG
86JTBwHYQk+YOsqzpsOxdqzZosb0L8BUcWUQza+AyvZBzBMtywo3qpldWvThPfh9
DqUCejljLr957Y7WTwlZxA7sI4hYghMmSDBKuctuLk+T4mWhX1p71yTsO4KfwVvj
kw5rYGBIo5d7KBNxpuTriYB77/KHkIjlDGC6p9Aqq6cycZRD0KsHJi8XzF2YaE7m
G6ZUH+6chfHv68hhibercfpnxza7qBfqSBLHfCx10k8IFoSA3cxNYNOHsvoh28aX
XT79slMIPpk5sffmahevWK56X/MNxFnepHef/4eWaodviGLGj3txJTpfhionEMbl
+GokZk/WFe00VSU31b4M5HSz+/kMmAscapb1DALWXaWrcHnxflV4SK4bnebr3IiR
EeSUVxsPDq/kGPU87dT2+Df3AYqon3t/V2xpoCpkJVwywUgKw3Mqukq+iMOSrvnP
tAIJ1Mft2hIOHMa30UnrwceAwiJ2JEBgZwu1l75Qh62nr9SwTIhE6pYw/Yr2ZaTm
BElwoLFJD4qTDRpuydpH9m6tQx81TEsRnggmrsNWucRgPckyOZdsMe/qXgiTXKQa
scg2yWZIpFC1DhgA5WPpLEcqsAI0lf7Cunz90t2X7C/oa3tgOfWn2VW2ptlsvHV8
Gc0gdNI5Pn3O3aCXFEyYgTh0cisTEAsmL1bLwbNOkOp/GNjUSNqmQ50Bmp/bf3Uf
M3bOLu467WnrM7rG9QD2AQelXMWt5bjOqA0yKDtwOdEES/P/gXLPRp1dw5zVb9SV
/xZLU/DxXqi5PeBbbjOOo353EaQNO5Sza+A4G/0cGbuSIAAsiYokel82eoBy3TJy
qI/3+TvCbE+Hxl6cixzn+/rlUVUPBZ2esyrVr0BA+cwX0w7ujKTMWyak90l4k6Ay
UzayQYX63dklxbkph48jnw/LWSpWmKKiC067wSeHBruPxdBZ9K1fJHMYq/AKKzP/
+3KbSlwXUwh1ZitgWtTgm1jl59czWmYWtZSEZkhfrTjL2fCCfKwVSaFla8hH5Ymi
e5fdopL78lROAYgNdxmeWF3sWZ2nxviXl9u/XhYrXqx6tdg4MjKm+Q60531PS3NT
wwqFiUHSNZkOCAHcBupGKiyQ0Ssd0J7CavxFJbhdq488iYeJ+SaeL0v4/01vDeHS
bAZrZJ7fUKH1yFC+ZZGFSzgD8pVP8F+ZS85c8hKopPDe5mNByBvcaFhT3GFTQO6p
YR2glqoGub37tuPvU3FQNU1F3ypUax/5620jk2ABvZEWBXZ1QxR7maThVA5qv5Q7
NQvKkoWGfxU5ILOT8Ll3PRhgYacgvPivC7GntTFyv5wGAoeF8GzxK+RoZL3QX5s4
HIb5Y49TXSHGhv8er5Y3Wq/NtTvPC5MrNTAXnoEn1t2RUGjym1GzeW+U3cV7hvHo
gjeiNlmayadif0aC4sCyQvMsT3N63GZt5UFMa26g8634eqQ9y8FrAJz4ijsB89Qp
0gZD5fBEDTQuhJLPIJSTezftrFjhhVPbtuNDm+KAe0QaWn0ZJx1kSq/fPCvnbtLU
zV2eiX1KqRupLV2ycuGIL+CHhbQb+me+iiuJnP0wLp7X4RGONTOuxL/YC7KzxD4b
sTNk6WNrx1QqvbylvTWglVzcESsb9dgMfA3Cgsd2kBcKCx0EMTXXVng4N3VOSKfl
zHWbsLiK+a6UkEWngJFpvfx/8y0kBO9IXw76oj2Ctr+EnkUDCP5ZIgU4gthjfDhC
hNRY0XcHiuw+cwjcc4PCIYl7iaHOEIIQBma3QZle1QPniq9VW6+dogjpdgx1Yrmw
smu1cHUmohKSyphSITfnyZEUjI7nyVuIbDyt6Q7gyq7UrHQmv6/gs1F3Cfp9eT2T
WNW/9p3aW65IxGyEcaPG5oCMiNNq5azbpFsMKQRCJK5I4qoSuzrXOShdQ3gg82ja
X2YdrawOHw97CF1IRe3gF+fMe5RD764ZH0AECusYlGgR38Jy9TxuWRmu7qtu6+1G
jQ1SKJW0R9qzYOjU2Mij2Xw/o2qqe+lEqL94zQNRR3tfWhO63eHVrzapY1ncL+Gc
rbE4Uk6tZWIWmQE299nAkGy1SHu0Szrg3gji1VaFhN4VAiC3haLRVTgMb77jEp6s
/cvWIBt5Fml4crA1nEZYdYGG4sCJZDq9z2V6OAoolGED4tnpQisXDHYDFnrrKXb6
DT/BcZOg6CeqJ+2Ri2ULrN8nHRU5ybIDqJkO3K8trJ4g4OHTgqrCJC/io+NqZbJM
0IDB4J0yqI9befQes0T9XZviz5quy4u88rqbAV/jnChFG3ACghFfiUWpKYRHlE/I
ByZVL0yTP0v69GviE5FqZJsJmVW89dV6x6ZEZyUULzeQ8qnMUdbaiz0Iv3se+MqK
DJXfaKjX/3VO/Zk7xyqYZdEwXb3R8gyHcpOEojPOqm1kvZq+d4kxSrDyvVSTChmF
LEUM6BsFiO6W3Hvxl98ZS+2TlAa/8Nfi5l6Cj/xB7F8ciOrczVmqqz7LqAa/loTC
maCQ1eLXgVUF91qkE6XrnjUHt/1QbxxsbPW1k1YxI0mFCifxjpInc7dZV3+VUK9U
TXnOt2o8VZlaK28y6FOgFKi04P8BGK8jLWmxkOzRzv0GQL15SRF6HzjBMrCAR9dt
zdR1TZTuKdB/aS+qBCQrme0gCBoTQzRgHsAUuaQgDmyg+FxJ8nEAXmYH5IqbYEFZ
W9e7trwlkP30FSIi43omzOyqXX8PBxXIVAkLo3zJ7wkCEXZP87cdMBkmxQMV/KI7
ZnXEMp7YjEGBdctJ9LfhhcoQ2e07K00CGnTUMVn9bKjMbhQ9ZPXR4hbu/9CHnVSI
72wcc9XROwHSJyufpsURbknobEOD7Zz6V0cesPvfOawBJen9Ik9DrQeFU9DJd50Q
TNRkM3CM1CeqSDJi1GpdJnxJrKy+JchhVeEn/E3CNXQCB1Zdmq5fTwRrbytT4VIA
WHWt3f2UuGyCR6iFzVTZgS7koQNxmLg9f+CwGjKQTONmnSSOUH0jQckjXGE4SNt8
NlJBS9wlueVUKMuR/QOdR794JGtJQ7fjA6Vc3y4c6dsHARJujWsRDu/oIl1Ft8/U
VxZw4oD/0ndB9NExEYyoXB7h56dqDZ3P2MRL9Jm8+xXXB8FutdleX8VwoZyVUh6M
sJS+qCDXNUhamS6jMbZisQfseoidfolG3CfX4HF+ImkrYbgiu6LYtebm7bltctoc
qKWRgBu1YCVRsFJKCT3EjUuiiPkVhGOKIHQufpCI02i5/VwWo4fLxPXpTLcLsADa
l0vQnRik9AsBjBDkCJWYgDD8Qf2tEb+8wsGTL9jWkXmStTUV1jUEpiLSJwBKaajs
h7UkjIwXWu+rHkb/cYJWUmISQ6W9AiOnQJlY8DCQIqG7zYnq4uHErlq0A+dmObcM
ckv0eetRkKRmx86GzdSJWUMrTVJ9TQxltgdLROD5+NYPbqefZvPmqKWsYlqEwBU4
n6+wq0R5KWeK5y7vn0Lka7spjIcuOtr/mtcV0fppw2vMKTZvPBHP3Ep84Wpg5H6T
mPlas0m6Nl2DwwIlfJMc14vMrFgSdGB1ahiZiap9P9GXyzWOlg4y+zYhWBMDnbdz
tnNz1KewAASQfDIF7YyAkUFbPSdD6Y3LXb8Nt73n7FjfwRqSj+bh1cz8gKzBTnwX
YzHPB0cfOMZJmA4a1ZfQWkQ95tPmq1DM/eFVWR1AbOjCOm1t3Qf/3n9AfVr+76pk
WBACiRHxLZbjmuYfR00p6yG0FFqGaEOzfByBfxeUcy0DlNZT8Glvu9NUqrSIacxm
FfSDofWBAGuhadqjUULXPnIceYpdjXH/qs3lKG4l9GVYm/zF9h1eLaTW7rO6pgFm
/Go0Ttni8UqnITNCyG+YN2IAm8FCaiUTtAQR6ZtxVDr2MfZFyo+TC4PzPPCRqgCo
Gr4S7ikZOp/ZOxFKb94zpfNfcUdcFINtiTK6QIQEn89hIYMgN+DzRcsNfegmNFeR
lgdJXW8/HrbCr+oi43M9+HO18Fh5vxwCepQcMlFa5p15hhwJsPuqtQzga4F5ahjE
dbrvORwtrFx2UFoRzBiI8xAve3NdL5Q+xp3WsGxim1bRW2N5jDKXePXwaDJQC9hI
rgHC3eb6iD4iuUoUo+oRsUL/WvwCTaLowN6/tak31f+57XnWD0pYXB6CDjyJclE4
rGmVyw6mk1yWtcwG4jb/qkmz0L1wT7w0sHcg5fyIhwTZ7OSDHbGRuVMbCLSUJPvW
5LfqK9YKI5hMmsHrpjty8N/hKymuG2ZfEcjVENlvGlMIVdSSlwUw55zlKiW8lpFi
bT0ZA7Z/f/zxlvM0hDTEinh7nWKcpQLtmON//X0T+gdv9LdX3Q+G5BdKiEdXWBfK
j+I36exksZ+kkD+B3oKEZ7xVCXTDOd1nwjfBLs0UrIJvNd3uOhgfOz3Lv9m5Q9gx
8P3AT56RoQfk7kfkeGyoD+3z8LxYcGPuvHzij2WhFvqufoBf5tWsovFlFot3BjX4
3lsYmlKWPPW/gGLrTvZBi3SU9fwxsPhQJmVpYZuKPz8TMfUX7l524cLTG1odsv1f
ZXwmUt/BIBCP03TsGSgXYLZKIEr3/4XVfXAazpnO/fwLQKV6Baxp9sU67ygUeKPX
3VSscAjsyygWEfX4dQ4tfXluc7OJDtsjzXiRr4R1Xu7FFad6/3bUvJ0QjWtyaUJG
fkKprIp5qfsMSZ52GQOcAniQ+C02jEkL3vcRoP0Hv5X9UKcdy6tTUHRyA6DJ68+p
NSSLYv5LWsGxj21/Y7jCNY2deYsFkbsc017MP+qtox7e95K0/glG8fatRaH2640z
Wb1/ciIMqJugME6VM1i+sR5xtBlacxFZn5SN81gGgD2wL8+S987izgci0OyLMkRS
o9pC0Gblk9rZeW7bkLEYzr1lgpK3vUog+8U/VM/0dAkZgylNgxR6SBIHVA1ULz9p
K3G/yG9xJjZLdhapjyHsUC2faJNM0Xgahc3PCno4Xn/JmXpIl++VPfgpNrukKxL0
ZuLVg8+/3CBI7xFGKVFDetTVlclsVUYESHilx83wxsfKy1msqrZKEoYt9DN+kQoR
h6kKPeLBPBUF4fYW8xPXiBj6rIgX+UzNGVuQq0C6T01YrvHvmRT501tuwf7g/71C
SItEAyfa78XZelRUXAkdM9prhT28UZtDxQMzJ74FYMyxf85f8JY7PEjhu/mfSsoq
DBhXSnv7uV3nRZZFzPZyAYvKyjlvEFV0cUPDR/jZRHoJtp6wKDy2IO16nEgjbAC4
2ypnQ3Zgr5XiYPRvtUNq2xMo6bdJ9VFsWObcnWvsFtL3AwXU94sHQUyEj+vtOq0R
uwpJFPCEfOyVTtRxTyw+K47pSoLX4jds4pneMkK94QybrGzM4M+m4OcsTJox0CK7
2wHW2K0MROAYBYYkPDNebzVlJy8ddAwcyBODedAHzVroJbmNc+6JZvyYFoXIJQTn
YVO4KXKDAN2Gz8DdoGLNvEBxrIec+ekEKX+yuq+Qly5SGZI+U/0dO5elmZUiwXEm
76f+wKiwZZhpWleQhbFHHi8OnuoqJbkgxb9mgAvTtbFSQG6mVsXMU6vFO3Q5vB5e
64ipKimZXSORvkQ/JWgzTPQ++njOSO5RGkW1deDF8QLTpd5mZrf9puRrCJ61Sf9r
c2QVCHE2Euqwf6oVQdeJFzWqJwtfig6eGKQeVWh9ibygdTuzxTxk1vMm1dQg7Cqk
kgnXzK7+fFK6mcJEy7Rz14OGuVLUgkenaPn2YVE3j6RaCXzV9KPQNRz7jMHEYknt
RbCY0c00SMJu+FaMxrJDH8QjYSRKSZqp0kkxkOdL1eC3AdM0HzEwa+3knZbc0No7
ZTSzDYB/4dUz22f+xF/avbWwPixwXRZYnccTpgmeJ9WgOw+tFvb2hMUBHj6dfUbp
QJ3R6xztklNzkyRDmLM85Y6Spa4ybL969oFmjttJNNIzkulz5ulDIm/Pg4NV+u9d
Tq7AzhrD7gm+frTXAtJjf2ksQFbny9aeDBNJ9oOmtBrwYt7bAHcYV9i/dx2dPFon
dzD3kjIy5qc4obYHsfVNAV9RCtq9/FX1tLaOXteo6HznCrr/0CL2I/0ekG0wQpal
XIxEi/MBgTTfVxWkFMZ2uCDjkoqVWkFPtjUHXg6RnrBpHbc+6vqjocNi79TS6tXx
FuD8Hs2YxoTP/w2tO1y7vw7rEbUGqtz7MvKlFw6nSA+Lt3MN9A9ZCNsqkB0KkWSm
iTeDnIwQAZUp4SZt5JA7BrQtNWrsvzQCYw984lAkD17ns4TvD5lJtIdo0EHrWu7V
BgCuDpvKrrMQ7QXL2co7u8ZTu96UDSTd4ndddFtLFvbffPKwbr21pM/A1LEF9ETj
c55WmqsURnvtSAPFMuC10wK2QsG14UJJFjX8aoMj7bRwjTa9x8S2Z5PPJY58yGAN
V+o61sscm7X2xoOKqMXTS5IQAapybLlB4O3oSLj7eIEP8dejP441lAkQssA936pJ
TDBsu6vd3roM/WEH+MVoC+ZOsKLo+pVXnK33tV2dRCGVwe4CGzvf2M7UBv59KW+U
cgYeOInANDgfh/dYf+JlIz2wWK1REgeUvNJinTTcMMr2Nq+2fNPOc1jihFvUftHj
j7s0Ws7Uq12tz7ZxmkMvBDVZ44OCsaMJY1tEg3WHwel8wrr1VU74Phz8RfSYQ9Lg
C7tOCq0cGU9kt4GsXH7Ew5vow4sWbYleSxnXvmGgeTJxPZ+LylIGsEnQ9PpYB925
7QFPVSdFnrcg4fuVA9AHgiBN3JwMGLPMci+ViCgbVJo5DCIapgKXupXn+J3GI0eF
S+ZiDqnV2z3Rj5AqTeGP1cxmxsn+zUWohXFVnfKUSQLhHvn4HnndIWQfk3qvYA92
lm9e9KBZ8eM7Af6eAjKYQSf5rFIGwv2tP4qw/9ljkLt3TEcwq5Bn4/IaJszZAIAi
TOauYSiijLwn9b0MlLyromgJ/+6raAnJt9rVWm3BOm4mih5A9vW4owbmQsD6DDX9
5HPmHCZtvn0KW+8gmFniN55xHCA8oW52a0wUExiBBHtoC6nv4x5fRRS9x+66Avpk
obdSqihywEUjm5Ne/1Qu9tLtuH2EK6bBCpmwxnl7FLobbmAn2fli3mTdGkpu8K8m
VOIx8Nrvd/fneCmsQB3JFOyPNHsozBZAMmfQFNw7coPpLIW8l1uR6tzJ2kcmxc9w
Z3f5qnpApojftSpFuSvqmscfkgl2apGceMry3kcl3Mu6X/26LaZ4Zkdj5uGjK+/2
PfCo64/+JiHOhYlA7UHm4RbwW57NcrCEDQc16BQumWWwkSQOMn6CBOFJHkOLZctQ
P4AyBDqv+3rvEV3RHosW6muywiSFZ6JLAo0SUQcA83NR+xF8Mlue4/ZdDSf8YtIx
4CZVjCAcHyV+03lmqcxBPU40xah+oYalY3y/KzBpdtkjVwnsvsmBIYae5vO96EOP
nHiy8me3JFxSR8nPF5Y8CGlzMymwoURmlUQhaoiAyEpjf/ylKvZZvmhM/54KX4ni
9U9ep5ve9Tl0znZpPcOfzQ==
`protect END_PROTECTED
