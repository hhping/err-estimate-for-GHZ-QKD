`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thNhm+YpiHSEs/86gSuoEaYhwaFe2NlYEY08qPwqzuTbSBth5Xpa6GNLuxJo9MGZ
7TnZRfeCiauQ9itI8xUsXQJdNGuyxHMYZC15q62OfFlzor6KQSWWif8asRVE4DrG
zMwo0/dl+r8RCD4Y81wWCYWF5BuZFHBnuR3141NtzFqFl3iTVVcP0DnD1wGp3X2X
XRDarzkZNMR6B7sn81eszRdRZBNtwBsGAqzMtlDfUAKia42hvGBFRYPE2rYE2x6R
8za2/CBHE0hSxlSxzOVfeziUpmUeE/VSRwuG4wLiQ/i1Owm0xI70lqW2NJrsOG0Z
x8CRxpbQlpsVmUHF8/UxitEzYow1W2KU+axudVLyKLcxYGXtvulmBiu89QX8jsJJ
q8+Dau2ZgVnjcHQNDyRzEJ+GpbJc1RHAi8c1MdEdVTsq6DVWj35p0PFd4qD7I0+G
WqNmkiWKa3iggco30tz115DE9O9hDU2wtujAbHfvHaBoP6AOksFiCZ1pzK7U5I41
e2X5/mPtm94xC5jO1pTqmaA/Qhevv2GBN9aXt/zNZdcNRGWG2iLwIZ8LqiaTo+6y
RKh85tPsfRA6t9qHN+yH9OkqMY1ePU75/wmrcaS+xwGHgHvV6+TXYOx4XkBd0Pii
4Ucoo8FW5MCWbr731HnxnlMYUiWjBopLqTN5nGpHzaUxRT8b5bvKZdOS5b/OObSR
YXWTotFm7GjLddClBfbaZ7G7SDXSudac44Ss+EVPScrZ4oNL6csPXTOl2eA4m9Z7
J5PepkO8BN71ZmZ4SRUm7oICYnRg6/7gCU1dEIjX2AJfgsbO2+jymNjpktxELtdA
svVmDDxFNB8acO8MoM3GLd9NYymAAcoEjaZrtxi6ZSPvksfFeE/3nnmBJE0DP6SB
UrNRN1tyOwoiMcikqR88sIfZT3Kd3DIeoLnZ7AkqtlpB+dIo4eeKLGObaf9FhbUB
8PqePwK7XBbKUxkcermdPErtjVRnMBufIwSNBcUBUxnDYjZEgX+4Em9hxlZK/Nho
Hte6LixwNRCgonya5WX525hCheFFPlNF3cSG3vWbm9eXXLnW2e3M34Cffj4roiQg
oHw6KQofYX+fQ/Datrvps4CKwHHFaATsJ5IN/ohEGgHVCgH3ie1u8eOYo9DY/6Ih
3szrasUMRvFFg4RV37ucnLT4uR4dFdOFFUACRFNEizmnIAyV60qlvgHfrZfeKUqx
lpmEuhCBm1kP5R80OK25oYPO5j8WAgR+n9vwrrgCHad6XGJpghmIdw9ZVID4WOC6
1YJ25iijl9iH2TSwOkW9vL6Mj9PPjgumoBUqlBWexEXVlekSc37Q1FjUmKYPAeJH
t/VkR69yReMvH+1p7WlVkH4rTdWl4D+hTyhPAIkW0ltSoENujJcRNOylsYk/PDfd
QS/ySpalQIPPjOe11bgoTbO3T20KNzolj8QYucLXeBMiQEF9f1QlFqHogq6BukS0
QbTYF++kv32YpDJstZoJ3tsSpZf8sxr+e9CW9gC7KjJCSHI7CGlFfp10bVr45DJW
3/fqGpmOIQWS8ywpV01koQ5CAGhE/6tgopk9pRmquD9h4DVzLbwUnY+kKEot7ixf
5spoMoZu2upFw9UYd7RLQ9/mUxHX1z5JtMxniu2mU6TCJAPhg4fiuFYq1B4/DgyP
DKVTkc9wI8SnM4OK1lMYk2hOhBUqXkcCHvXC6KO8Qwo/2lazT/cAdIhJBDKBDlDw
VgIcY73VfaSSNTLophwL9lMGjtJqCtQ7i2nQJnIVBwDGx+iCxzLjlHzf2YIN/lcB
BDdTgBoT779ISM9o6TATsVOdBzSmM6fBYJWt2nNRI1t9dAEwzddtwltYqIOF/izV
bYptjIv7ZknL6T2SjkkHImZEelKl+nkn6q75u1o0szeBKgbcIWLPRSNC+joaJ2pJ
fR+FpQjFOhxzRph6/xGIDyEl1CKm+IUC6Od4E6I2XUP6MoQqQDdBvHMD0Idcb6mN
P5TkjJc0cXvaQRphwlj5Ey8Aocb3x1LikBeDSg+lzF8OfqGuT5F83GPZLOCYW+tj
GBUNIwUFlhlcRttOGOAQLKbY5K6W/sU0rjD10JEH57JgjKHdrjbu2WtY04mLLA7z
xjdPFi+ppjbNoDbtJOdtLRRxr9tkib04ylIYJL8BHwKFavMKb9OG78Wz1bc1LV7s
TiuknwFcCwHzQTZgSWBmAi1LI1JYfuwDkXwGazggzmcgLVoHKNJe0mDc3QuXhEBH
pFGQBut3ERbGHATgdOp7HtrCgljGLCbDeY9KUInKE1w5euXf7BLgMS/v6UNaH8YE
dAzOB5r21BBiyXxaBWVI7kL+N0VWtQLLfkAo5s4AP/fdfmJi0Cu0hCjSPbg7zK0B
vpK+JGAVy/oGwgcWLlLHocb6u/YW0+HJiOuUjZSstKbf9pYlYzlHdWTzjcV4ywKR
R204fFLDK/NGkumbOSMJyrDBOOgTwHNqohvg1WcseIcsUyPf/H8m/CLpaBN04t7j
94TNjmK2XLQskrw5hS+PTrrQYNMWGEfzmETK4Y67Kql5hyB+2qFQ/8W3gS8VpJEd
Uf258vifnVnXtth+ep6AQgUd+2uo4YtjRzUbSd4FB+xKos0L4o45C2LUqsf57I4h
`protect END_PROTECTED
