`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dr3vEyhM7ovX1OtwpPfc0LORy6vjjGGjSpWgMwk39zVIaUbFcPOvv/2xYCUn8Aa1
PW/9ALtz7q3XV6zBsYRDBj1X2hXKJMce0th+EcZrT32j198Wg5J4qrxQrRGeEqh3
jRw1aRmV7bvbonOMPNdH3Sa3eQIuIL51NgH1dGZ7849FzkMr+j5BkS8JCgP6OkzT
q3O2co3mxizOd3lOQIpSwnSBjGC2j/gXSQQr31wAV4xvuiJtBKT5dyTqPHDqwzLD
GJqUFCSiLYKAaopcn1MlsWJ48w2El3An9kduv/y5ERsWVvf+AkHcPdoDTq3TaXS5
jPKeNnWlaY4kr2CT2a9SYqbjHYIR5w7I+3zDnQhmI26UHMkjwHxuXJQdFS4Wz++c
tczPh88dlKnY+rFztznnHY2MBqmQ+h+IKnntfT+euYFNdZtmbw5aRmL+43lKR3H9
SUD4FThwLmi7Mybq+C1qK+5fBYFjMNk88UEsJ7E6WRF6Z920gIgrQTW13soYTgcN
XjCojMuCilykNF5U0+2U6LxQYDP0gyPP9oQWqNx4X514BrEIzG1fiYZWya+pDrmr
NBn+iNcTvZ4tKnZQ4bZcFxgM9frLnOgIkdDyD+tXfanXkJCTl3sTHH447hjwk3k5
wvlaoPLAFqp1NO4ehyH2XtobPxtGkCmEZ70c5wJrB1O64JlpV2vxZSCxohzIMHCv
P0JafsAilHKH9oXr1MPUanIf3iFnBUuuHl/F3Ky+MX5Hdx/Gt9imk1VGncCQYp1t
uXvdqmx3tbwyowuI3YzXlFyCBrbZ5/cGnqh4zwofv6qjFqrWzcWlWm1KyPwPrLnc
AxNpnyelaC5Bz19uNLSCJLNRitaGZeYAYbfZExttbcA9utvhgkzTlxnGtW2WX8AL
/Zpv3eyT4N0tGLW2hu02l4i3WyPPO7hpqwReZDTFrrMrhgohzVn7x0M3RCKbRr8F
M1J4/7dvzmQNhBlTTg6zA1pF5p5pMrxJ897o0e7UiLprA5u9mgays3y/NHUQG32e
asQcb5lLDus0YEzZhmjXOie1SGPRC+jrJQJMD+7jQJgA7Mk7FJa2MXwkdl/ZukBe
5phIYQoSCDvPx//PzhiAxAEKolAvZLm9/YWo1VosG7hWx9q+6wUPfhGyC1fUGO/6
quulTK6s2b8MSU8O3R5RX+xKKR6tLNL9FP1qWijDAIcItWz/i0o5FS3zaiN4AyWR
/yLabvpbCIRMIrVN7VbxBbE19beJau0tRnBL7rZtPLW8fWIYiGBwcVJdEl0lCVuc
jdMwrot32XoZ1CS6kos/fgBHAmjVE72hWt/CF/WJckP5veKIMtnIVNjO08hhWP54
TMW1dRhWQVY7/lIJ6NhNs4wr76kI0UuZEOrcg9AhJEYI8xBk8XTRGkFYlt/5SBS+
FirlPJiotwfpEkVZRC0fw2s6He2JQVIyX+dZXKXPZamaUhI0jtLYbGrYlL8QDRpx
/SDm1vg7I6AchWwP7gfJBItacp5ZQdWtkbdSjS4EqLQ1/oBlQd2Cm1fK/+kMPDhB
e7q0QRMAW8qMxUkCD14HS6roVtOjU307ZrVejlTRA4VA43KcE8JFcV4oD7Q3C2Ns
3oHUcOToSZWnZT1IkIXG72uRRkl5l8DDc4tmj6XPL2tPgjUtYtuTX8fcvotYu3tF
A14fand0xa+I86dirOJOnQHGIxgRoFyhZ/vtsEhC8vE=
`protect END_PROTECTED
