`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q47eVQ7Cjs9q26U+lkroQGAC8hJPq9ZCZYnzUVmK7W9jKIZnOYD+1CVgaDQUf7E3
YMc/tGtIwzc1zDyLfXjSR6L66zz3TMN2YS09zZSDtI99adgnm+ugAkrOwcZuBTX9
xwz3ejXmvChyQCMbC+tk7eqlEXFu99UVgIbLrIo1spQz/cewrt8YoRBQEzfsCaPd
KswFwr9nIYOtjrfDb2LVH/Pa1F6UVuBs6Zk41htH4Vs9XHckspAgqXJOzpoEHoxB
1njE332YlY5v5wsmaV1Gj3D5fcn+Etu2Rm7vzr8go/XJ9KtxFhfNff1gXHAuN4GH
jah8cosmglo8bUl7RThjCxpe9r4P8jabBpXuW4RpHzaoepn9P8+wpjhBJdJEYAum
u4pkbbyqKl5LbyFzZl39zrrRAB//57dlm4ikU1003b4l2qltGN7hTHDva+KmHEBW
qnhP/2hqUH31gqE4W+Vtxr4Ab9eeX+TQLgtxHzEYSaWpQYTc/bIa+EnBwfB9CTSy
`protect END_PROTECTED
