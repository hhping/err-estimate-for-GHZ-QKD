`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Y3hICHlDfSgJk6/rHKV1S2db6cffgfn0iDG6joS6BNrkZwNu7y38c9VXWKbz+0u
NcheSG2W/n5PrdsTBSMamZepHsg4Z1MmrhtNWPR191Dihi/CT6AghvWMjhwKDyRU
t4jAFUMRphS5ThBM5OMl1EJO7H2S1i/8GZNrs8l9y8Nz9iwu14g5TiJ5/56Da/Vp
MzFKPwDTbiky/m78AmHCA84jplowl+o2P30tSK1qOFEb19ewFQylvqrwX4KBGHCa
0EX+C3AZ17PkOpbd3QOG3fFi1IjunKffdEofAjMtKUuVpXZcHTx1rma/QBclGAZ9
rFZwRQ+gby8zHkNplqcUHYhy4ueuEkfuI4OM1rPgHGOGTzMLpF0cw/MnhfKh0d0B
95kFv66neM9fvW2VUy8nGHiCiBE+ACCL3WAR99W5YzFE4CVe+p2r3bCK31n/5+bd
LnY/SA35ZTD+Xzmpnlm3twP3OtdvKgUCr0gq9d3LKNlfAh4YLBeURBTjsyTc0iv7
f44kxmkmpuHwvaLb8868VCDwz8gnz/fRHtWnnlNJ2Z4Ig7H4z+89LzAwRgojj+vb
jaLPq3h29XQbZQsweVQvJ/FgQDcHHOdX3OpW5liXk76dzNYg2f0QoZw9BqzI5/XU
gf0BahjWudNq3flTfFyRH43Y2vYUu//1sBzhF3934y29BLnhHuIz1Y9HtathohcH
tx8XPHHPJHlnKVzNFESE75lGz1V4EKsSFAD4Y3G/MaedKcZ48pP6lX2egGqv73D9
ag0IiXsV5xPQ1K+ahcIl8bXQ+BNrOFO57LkEBIbNSv09aheNz2igcNtH5ykFz5hx
lV4A/l+AXez6z5vJLM7BiyqJIfG91ttVupJm/pTFoqWJJnvadiDdu7go1ZYabVjl
Bm+6xn6aHx2EOLu3mwEg6CEsqNCcGjGbLUdK/5cYUBoqiEh5unR4cZt4QkIWrpTr
Oqd+SJ1r1BJChWoOzuGSgTembd/6hRzXpOZIj/vSYnvszaMl/c73vmNrVskBdC2Y
WGcyfHVJEFGG1+s+NRkGl9/zgoakSd+OgsLUR5/WQrBZmcuixtb6aHpcifCSJKWh
YTaOvZt1OAFLrmxVqA2ynAFWGsMEEgQSz+c9mNp19gS8bixWaLOQ2j4VXpn3lZOa
YybOdkcN4gsiu/A7FskRVJgnTULLSSc3aNlnBX+tabdpNJwY5ung4h+gGZjK+p+I
2m5332CG4/Xrf88asBnd74bOEIjvrY6ZqIG+/SJh6WCHQoyhcGiF8iZneGyhYfDs
JfqtWvMiZQO+UxKC3xqVXrxiD2cFO2RTfRydUVWUcN83Gfm50P4km4YtC/szxRf0
`protect END_PROTECTED
