`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHG0zrOBk7/QKotZF8dX3O3Sk7zSmLCbFFqw24T8ANG+yUqjryj5AllmkYcrZ40h
ZdQ1XQcB8+sBqEvku9x633FVS0tX3IvHPKlD2jC99UTrskenTGr0arSIm8aoLjVH
siBAbNUWw0M/lWGia/y2QNvrPsQcslC5BVTKZZnufRcqo6+HjUx3Btv8Ii2jBkvw
5vANyqFgaC5j2ODitFVTi8Mkxuku1WkMBbwUyEf3QKR2iUaqbYeNNtXWCeAXoZvx
U1HeXPQr7JcaWAL+pM1MvjLWd5VLXG37QafSUcbDnY1NUoW2ikjaCx1rOcedL8vc
BfvN60IO34BHJTvcB+FNqJWNTNWM5YWTTxRBcF6ru2ARq5fO3zWkBWG6Av13WzHO
R1iJglRjsUZ53g90cJUf3MnIawY1eQdM4vL9J0bolpJPAqeSgN5qvE3Z5mEiVm5p
15SfXVUn0oYDSNE7+gKS3FQk8AY8OtKYIBsGqX7dkXOtoAaZKjYTdQfM+ASEhGqZ
FcK9wqItey7lAojDRo62kRsRB5ZRa8JDB+J6HttztIaQDEnnvvlv3pBLKV2Yqk0z
d+VvoFxzcLA9LLo3FDrigqF4IiPX4jPEsrfmL8KW7/MX6dbpxwTovRZy6OXTw5e5
greTgU8XfqtFu7KeK701L7NgkPrj6Ts5LD/er04xz0tyetO8hkH2Ew3YQ0+ar2d/
/50fPFubi1ECovgMawzbSEWqhJrRW+mnvWhQy84X70CjJ6Fse/BEUcbOH1C2R/PO
/FpBM9k1a0syvDr6SxPD7GGNhznPeBLq73DRY3tnNcaMLIoBdMDHeUxgkToMsd+O
Pi8UgqDNBNjZdeza3wm82xG+bYSF4J20/qPbbaQDMyXukV6tJ/B+4VFlPpKSl92E
eJaRX3yL4tAlXuZxQ+zomAudoD9O4EYq3mznBKkn5YBXe8ETezQ9qiTCD5Mnso5H
D7fWG9yGVfRYC6RjF3jX8qyVnUCfCLu2cLYcMBNwbtvoXRErxDccirAUmdYLxibe
7Lu/QEHZlcxMIYmCnxE4NmabTTNWtCwHqVdlh2f/syPMAnCmBo2jZzqUQQMvovYm
tLxuVSquAO0BR/QsEs9eNZby/s0HVLxNydO+470dWFi2FotW9+waTlIhVRQZs/ff
Jh9/bTCMq0R4KZ/BsJw28g1oCUFOqwAUh7zXQBEV7Ba9lR1i1aAXfBtLIYFsaLVp
bU0M5UbV1nauiBt7b2lEf6doIjGeoYh0oBTssEN/2GDwb4LCNkc6rSWoR+nUgDXF
QXh+tGPGRDBD9gNOSeYBC9ML69hrWQRNP+Htb0+t/Gwo6T4Ooli3E/gQH7iZXhz/
vRjiXgxNLObo5z/OY5oYaspZ5/3d6JvPCUxxQhHuJkhqAl5t/BJuOEGK51H4Fk1x
xaqY+D9tH4E1gL0M/3Dd0KewWe1NiPRa7/PtQBLSkArOJTYhtnxoIC3LhiBLvZpW
vnisOwdJs31VkB3sZ8KZDHBA6msw3w1q9MV1QND0Wu0HfnoN7MunFGiiuE0jfFgl
PKrYnH8PB5NOmyOGup5tJQZGWezaSCSF/pb2zeglNd5yZhEsaAlx6AVkgEdvjSD+
PUTFl9mldzpKAglBMvxgdtBkCZ1gTqQip0A5W+LP/jt7d9Uyer3hYvlP+MyVADQm
3HbRed04aSTbdBcOOgOlZKGxz0cTxNvMcgFyjuthwt8vBDtht1xLjUwApgnLRjuV
QFfyHDe0Pr5ex6zaoiPBpuaqL+rU7B69eajb4yVI/9ooyFF4lPomBuQBd4rQ/J15
5pfhslOHAiRmOJ43cr4FznYO77z51BO/3TRJyDclye3Nsf6aMbRKom7tl+k0JgfI
htjQ0liUmmNv/bdB9imO4soBOAaJGDy/g4/VpL7w2rTa45p/eDZngo6GymcI7aJd
rMCkFHdqkCk1hZWds2v/UQSJrnP5rsk1r4X5tSH6ItEyNEKrG9UZfUGF0o3dcCPk
XC41UXn4EHwyRvd8eoe49GF4MCs7thk4yONUL1g4hH/CkAS4veQc//JV9t+i5wMg
K74FA/7xF4liloYiFIbtIxrrWD9N7ZHsBwcWClU5S4dQxHkpf7WJCU2cTxAwkjXA
YBslukjkGTAWW+f9ob2Jx9Xu2AthNBoPbUGhqh8qm8KxDs04XDNmYU+pdqU6uo0n
O4F+QXxcSZ7B0HGkgK4CstsSbVI9ofaRcdYh9r0YhO6lIbHABy7Er2BsTSPHzdOC
yefu3kOwmMdEVn4v/2OljdmsGNPT0idueVjiyGRbtPqctKVNFxF0hUurN70IUATD
YY/CDvfXVEnOYet3qFySKw==
`protect END_PROTECTED
