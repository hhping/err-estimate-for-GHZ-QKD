`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sORY5kd1FSQn82H+ncyv8AEIHRksYy8GxYHc30Eq58IBT819TkxypkMZWJTikio
neCyOWyoZInvog5Nt3/CO3zrNxlVwo2BIFLqxyINavvI+2aKBsygDIEsFMw9ecsq
Ety0nfQJX5czLJSjZUhWX6ppa4fJoztwrO3xYWHUBGloupSq2/OGoS678uJV8HEy
bWvOGyOHAFabqKydgrskQ2XwGNGEKoyRMdMlDBm7rYhodBCAdEubMdMh/wMbX7+P
EMfXmo2cD5QJJhHKeh2Okj3BxB8x8iajw/3/Agv/Manu1rnZBndrXnvEIrGkIJqz
9tVd/tAfKNyEu/+e6cHp0Ebhz3ILust6YlCloBI/C1h0x3h3bf3wBqvhBwJ366Gf
eXmq2ByoTwtzXHjpCi3y4C060zBdI/Ke1nWFZvZje+/J8IELJCEFDgFV13bwc8XN
Hxo+Mxr1m2ZPMrb9EH4INOnj08ttUzM4GqMh42KLtTS0Dno3EasGTYqORuUnA5Vp
04nGf6XFMirDsRVJ2BcR1PLXzzK66fdts08B1REBy3SpcQwuNBkza4HtXwbMUV75
AbI6zyfUF4CG29ALXkHF9bq+d6CznaT94SZ3FNyx5ig/wMtlM9RVuIpWmkkrQ8V0
xKHvL6hOn18YAWL7eNgkBi2QmYTUa7YLIdJKJQUpWAUOv9AWpoLuMSKw1XF+C4SS
P1qCH8XXzVj9fk3QmIjIURdxvnGTZvET0wAh+FO6DoHNSSyBiKqcPloR67HUDPQi
xBnibArhmoXJ9wyUicwxBg==
`protect END_PROTECTED
