`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J4nP7ss9L/gPHb34sAoTsAYOlmiIhc7SqBlEE5CHulgXEINNnC3cwj8OtUwixbSy
UIrn8aCuydb3t28BlT5rAMQXAdVa0/hGYQRFcyog75Sadt9arPO+y37NEp2V1Sp+
lHRHS52JLQLLPWPJDoW5N8Mmb4KhuEgnYS60EuWbl6fScGjIr4LLpf5BhwB0aD1/
tjapNNrqjeqNcbhfuY1j7t5w4AXikkwoEGXYJH3D1jPXGJ0C9zoPHaRLxZ3Y/VJK
bN6CzGKy59Vcw9rC7XHfqF81MNUitIrglv35EPPcogkGoZXzEQv+xaCmtDCHc6Z4
zY8zGeRcikyXO7XIm64kVFL2H8cjvcDCD8uedlM7thVYF/+blrR4VBqDR5HQUWmO
L+t6Orq7Jd2jdeneCwkMoiDm2Xsom7QfqS0lvr65EJXrpzGxQA/X4Zgdt1oEhklN
`protect END_PROTECTED
