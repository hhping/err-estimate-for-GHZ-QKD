`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbJMGgeOT8rQcTZ23e50H+zgsdfg6dukX9sxaJz5+0OaJAjPialNNO8N/38/OHTT
orpcu4FiWk1IHW1iB6oMIiOOFrAIYfw/dpXgD7oh2SBZ60CbEcRjzllYhGr5BX/G
mdZd38ChIyMlny8u/hzruhjsbXt2ig4EvLY1+eTI09y48UdMJ3b0/8Vk133w+vSk
Z4U73gzhkoWptt9vcrDuymvTBjNUXdYBznHPQDjsJ5lo1EaEHREhROmlnWevwGIb
udzJ0Peq6ZIvP2L0gj6Ik924QjSeAIcTahxF+RbSPXXhW21NnHSRPdT11R6H6eZC
op7cU4XW/Z79e3Oyp75MYj7uQkBMgEjqwAcmQXtj+4urYXZdTucCeoL5TqPLkoYs
i0KM6pk+KeJLXh4HrYAHbFlk1vK8AWQsOZXdRS1Krts29h4JkdMMR7i2G+mAzApz
wN+x860TgeKK4JgY8wyDhYxfypOn9kLj6isvxpsBf0zJV9JFR+MKkWXkklapZ8v7
tCq8PzRkNyQanvNBUJwbDMrMShWXqf1+MnHhujCL1bgJlbJ4ubakIa01jg9PD9AD
42GrufoSjqff2jg8jo4UV/m7gc1yFRFzzQQxtphRHtZ95oI75ud0uYzw6mwJ+M02
B2U1OKoZHroL0TUr11A/vEChyDf7UjAMJGagxsF7ek0BwCIn/37NoypzRHMHOEob
1QwVkUeel1hb4pHN1pJmmIJVF6oxkPdx95BzMITGlL44QHta6S717mmamae7ABHc
`protect END_PROTECTED
