`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dx59bQl/arDDb7L5hmmKUEW6BxnOF10Ijeo2NVaqZhmp+spkzxGR5yF8CJQbcHNP
EJsheiBSI9vuVsRUcOsyBG49E2GjLZZ1whHfGkZWjY7coXFYdT67hiUSTK7ueZpy
OwuiweV8S/aNLo/xsn5TCXcn0MzcYl8Lem4nOTiJN6GVZy+MUsdv5Vt6pJP+3wK1
7jVMzrbng3KUq/Q7QDRmlFtC+W7DWOH4//b4YCUiWzBrJrLRkGKrPnx/wCvoaXVQ
WPN2fY3/K6aIlxoPK39vEDHqr9J7On24upbpsvN9hiHhDLqLkzg0DdxhxxkHpdwM
1OhXbEfJU8+cW42qha35BtVt0snmg6T7WxHWQTAqClzAw7Fwa9gC8EYvGWjMfjvM
OCG3/D/UJubhauOHsMJ57jUkvl09ghNi5rMJmToCVfn51EnsPMzKDXcBzODCI4fD
mmT5z3mI+q6AQ5OYzwjfdBnzv8rCySfXGGa76CHdFv6nRZCZQeCqjMngcWusGNZZ
XRIRGN21iLZbjORwZkWAi2CcZwNfyspR8NiAIrKHBP+xcx2JTxlQkRLdbX/U1Mr2
ZAkq0VkGJSjhE/CXKJrRKZdsGQZ1/+y91KIlBGVV9wU4UN+eq1eK/YzEsLoj0sHj
QwMgQFPLM/0WAR3sy+fZyde8xmZu7FCKqtLOePtsPrxQW4JzAXeaabmUb9TccdSk
I/1Bg7iVYLZqrWsICgbPD/S30XiR4NEy+xg5zfCvPu0yfMdVo8or5HxUSNb7MV2E
F43aYnKpNBY6XvA92RNVV9jtp6LedsSAM2H5kgYTXD5T8saD3k8SLOH+3ceAkijI
y3NeFELAdLUCB45lTgAERRk3FouyCRNI+jJsd1oLI7a5B9ppaL7Lsvc9pYOT13it
6ZmZTeIYjdwKEDR/2Cn832yQnqGW+TClcD/NaKuVGD+P/i1sGa/x5OVUkLQaPYdt
/YI8+3NgXOGJM8s85nc1PiE15B+2zit/R0vwVLLl+E/h5VDD+ObzESMtfQs6cn7C
bVmzW70M/jaNOS/Wn1YyrpxdIMAK7gYzpJYt/uYxH3Ol14WhXIrDIu6wwWglbM0C
gWsfJDhyETDhyofTtXWiT41xz1bx3RFj38ZnD99brVgvaGOFUWfC5GiI3NwqxPXf
00NIqJab8Mthg+Xgd3dwyrskaFIjsvWOdc/2tzqcWH5Z8hTJQoXJ90Mnzd4bVrPx
wofOSOa4QxTH5G7nb5lHi7es3jMOA84N/UqnhjZzS3EQ4b09YELeVTVKm8JO3IxH
OTCnikpi8A9tyCqQQFJMgByiO3deMmi9ePg0uyzcp6k8OHbJ5o0KOTuYC19ybzL6
AdnvyvPTKzOyfZ4tSVMXwq6Lzz/2RTq1M81Cxxxc2xCBT4quIE8sgNjxHoBbV7Fl
/4GWPiq2gBSjz5JoPLMz4T/OLVZ6rIproZG/epg7uwdDBVIryuvLvn6FWlVimfxW
F7DcA4+lvLZZFLiye+5ReIIQ8fCY/aRPjYz4yoauYGzjgp7dzMTSjlbOAriX/H7g
qHRVqiyNYTh6AE1onLe1rc8XhF64o53lU8YjgTBzBasEv6NKb5D3rm5apQ7uiLy4
0n12ltHIkj3ZNsZHszKacmG8lrQa00/j771UkkeEGcaT4rcQ3UgFIR2gq0V+Irn+
fl1ypsBU3Td+UBN0U0nYkYLkHzLWtgCgoOAZmsEmxGQIPOjLkKk8Y/yWlmXgpDXh
9ciysTV0FGmWtJ1TSe9jFnjOVKZAQ//DJIpr7wY+6S/OuRHN4F/8xHeYPr+LD/V1
VpATmVrqq1BQ+7rCGLHkXtspnNoyZvRYCdqbloS59r/9B3euqd+C4tCqoHlGFEBJ
NTAspNR/E71WTmaS0YR6OVaRDMQN8rFcIaP37vilcNqXq53m1O5f0YSxTWA5+zJD
aoh3tBy6lwYiHk0YMi0ZmDauVSc6QVPHZ6G2UkSEvzXstaawVdDddpT1XZEz8wRR
GumiW+hkiAbJddrHeHjQmOkz7cxWSK1ThqkSG1VneqdO5fGNkVy1DkaWNE+MQtvx
1HD4Gvud780Bja/YCm/L/hgcd2BDb4R4dHi6nX28Z2NzdFB2rYrrwpOnyG+D9+2/
xA94ckLt6fcMA6nmy64dgDDNdrT1NqPwXkOIsFYPxPqA8uGUa/SeFRjDBKHrhvYG
9/OBitjl4U18a/Vcv71OAlu5xsbBQJlXDr5VMYWMQooz1pZOdcPDSKGE76A+ySU9
xuaIPb80HUxBgRqBppGNbhb9aGFrsRid2QRl2Z4Q2usVeFbK8qDd+80GoSJ8VlMh
aNRB8+Gr9DuaN6hm0vbM0+XkR6B01blckn8vuHRTO960tDlTY7Z8zPHzxwgN78B8
k4TLuUX0yndilEjGGnguBy/4viLe146wKEvTtBllosopP9P+pgzd0XwU1Awj3ISP
Fq4KkAkeAUyIM4T0oqqX5pnqk6Whiphj4gLx3m0KZZO6Taw3Ws6jj2uNS/pEXkh6
qHaDdlzw6GSzkPUbzfimxtkPXYSqGFhQ6lbETKf4BOSrvZsCxglPnHN9T2qSj7Hn
rRTcmfvsj0slyfqF4mSarBJcAIxpu7/QC3nRE4gEFQlp6dz4pt4bhJwg9oQgZHDe
VXn1s9+pSp3kEWhmL0HA6x+KJVl1kaVi3XBXwsIVnr/WZsZo3et9p3KNL6MRo0K7
jesSrJHOSDMEjgU4iihnAK8xBA038PpeQwIYiHK1S+PNeoS42lS1AADHXP73oVrf
KFNyCy1Y604xoN8g5VKdiZO2O074nUrtZHJJI3N5Wdl4t2MiX5vd116ZLXfy0m+9
NSjRBZXvEIvnqNxcSysPnEI1/dL46Z3hgBSmDYcKKsnNvIrc12cx0HGknx2WwpSc
IZvPhRfQyMcSrX51cLW45cCVTfOS6rCLQDP6WwY7ys5SkMCwY5zRmwnBRdQP7ljb
mFn3BIR+t/ld4GbNQS6I+RGlwB/wBmXBWW9/0TRdbnxYqt/xdyPUaVZXzaMKU+F8
VzJmM8M3it+XKxj4+lqgPL/RTgEx0B0m6KbawJXyO30=
`protect END_PROTECTED
