`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmJ/RXOM2+wKcYMXfrQ9WAeghzuMONP36DEtPYzrKBQt9KkzNV++tCHf1DnrdKUZ
HWcEkOGVKD7lzwLgHquZqdSGNFiKCwLfajfFiekJKlRvXHvdJyErn2sSJu4Xexs1
AdCnofpzRwxMp/evsMBSXLay6tsOt3hSJglj3jdzsVWxAL10ngx2t5BhqrqxF14J
IKeqXZ1MkmfmIgE3T+Hp0lIrH1nKqL6ORKgvp+BcCeqG8ViN0TSj3CAZVsPrsb+3
A09F+JB7xkqTCuP33VMXbw8483gJib25LpWBLFFOiizcCRQu3WZEM9WVOgU+zqqw
TfzWWFDaQ3GEWutzI8fv8Pq+d7D7LdsYL64q8NORJnDv4CgTNlk5MnLA2Cln12JY
6t3H0le2eM5Qyw+cgLp4kDd5gmM6H8E5HCtK3wvGg4hTDNKqnYUoITRWetqDIGHa
ToEuWhEkpygukne5l+zuBqgk6c+S27TNo55W2UsJR0zyxhoxOABoATnIAOfl4sKw
cmmUCGd9G856JuRXV0IXOJr/FcqzVJWOeOPxawI9aMKQfnZXi4/092HbqJYQ+Fos
5GSCFGajQKW2Vp4kxFC3FgZyE4nVCHzlYgXov9QM6cnZ9yyn7BqlNu0gDNyj4lVq
YeBbr2nZayIwbzYTyQSMN2O9EkKKGfOowqWqzoSVFWlreAAVjmIiV6NOsZdwpEwT
31tR+K6H6g9hSgVxwLmXV2tCiC4nHga4XYKWHbTX+S//n79hiEd4z9IywbI4Bp/P
EY/X5vmllGDQ835Hm+RM+WbZE8NS/3HBY/3Lg3uF9NkbbE/v5SNjhjAKGKAbiDhq
3lUmKykSHNEfytDtOF7FUtkkDEFrl75N3NUyu9ylz2hpQlO504yS5yGN0911yQ1a
5cXfuaCiMEZNSuEaTM0ftxKR813q1XmyzDgEUG8R8Wk/n/QUfPTHsId56gaf4n9J
`protect END_PROTECTED
