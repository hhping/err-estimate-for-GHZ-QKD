`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvxQuPZGdYxvVp78krTxUPNo3MTtTnduiCBXBy4iTSsh73uWPeFn8d0bAT8Cwqvo
b0gfypCG9rC/iX3IyVTOXtwatvM6G3THTAPosdymQzuwwVs2byg3E2uET3dSckQ9
G+g7XOCmWmwOp/5caHvWqZw0Ug9LNoaVo6wjm3+zyXbLPKko4qO3ITNxzMeIefZg
uSVWlvMjngyfld27XzrJc4V8aSgtxFymTazv/611NlIoCjZcM++61CA2wUQuPvnc
NEwsfau+BmB2mIqChgEiER5z/qeE1emueDeKQ2x/X+y5ZBCQzV7jUq7tjHjED8te
Qkw8cxvJCKcoViuXWbV+N5Zav8iKcXUk0TRiynRPWUlqAWnivN3XJKG8N9z3ZWeO
/bW80YlhiKqbuNNF4sw6+Gm76NYx/auxm96q1mPgU6fOiYi0jbK9FqGZiC3iV1CS
5EXCCoVQJtV6azE1GL1F4z/MdUrJacYImBoNLzVfDyprw0/H6llFwI1h77GnJL/6
9kRatCQ6fjI1ptFMdxQJSqqRyDc7EqtNZltCvyASYCDG1w4aogHCHpfWCSyHnj0v
sXMbNDCXyiKeeZFxGEEgKaxfooBDfOxEzFvwAgO4OmphUeCOi98hQEGf7Z8UDqAt
Jxh5Yt0zy1TmfxwDv+Ss0ibR5hfQSpe4UEn3qiwhtVxsbzhurRZXRoAxXLRH9N2+
91u3rfIovPIqqlA90NPCVQOOB6VOWdIbFnj+ujbjoAsFmHBdTD20koJX7kmuAGQl
/hBoU/qJ09G93D4JDcgQ1LqTsuLpcnhHHm+6SN4ioBxHys0yhJnF6R+Uzogfy4Z5
g+4F3zjsHPrrdAxZcpfbg0u82KwCi6Re9rptF9x9OGGzLouWPF+Lx71IpD3vf600
kTyUf1fjoDzL11Vp3hUTIKKw7+egiN08q+wVe58zsWPL0V3A/nlO7jBDhl6Dh3GH
YST9e+CAnv6vnv+N77vO+I0bwVSF3SPpcs2rVuBdidP49o9EanpojeSYRUXeh12s
pWcmvmwEtlqHkLtjwS37djwbyt5/qMIXBOeuNPS626lKjDbI2KflKK1yOoN7Non4
ADq/sIgaPrQMWSrvNNaV4f82xZCUXmVvD3vv4A7SVsfwoaZpynmT/G7CGcYcBjdl
vkXXnXeMJLH1cvfOgAGe3YOjQta/NyrY6uqCmRDFag/Uedor1k0rN4wKRQaKBYXT
QCm4fLRuHJrOZzEIDIX4H23ZrY5XKWTx+kjDfHevQINV7zcfL0Z5gLZ105rmzHcn
zEI+ZUL4WJ6tfRhR2NLLom86r5RIEsb08E2QkOl/C/Fr4S13IQ1LK/3GHfSZYOzR
0/2lFkD6DtmAx7ZWkYl5KC3Pkh92ouRsF7956j2u2FE13Ou1An3BOkH8ulB4MJSj
I+XnULBugZaHNCqjYnBYEmLf7wyb9imo9JqHHhs2+rCcgndhnKJSzBk4nxfUlMAs
KJJh3xt6sTI9qNWLbaQGzC408GbSKrx3j/e7VRYxaXl6rRR2Zlq20BqAo+QPmcLT
h8HqeA0bs78dyt5l4IzMPVdO509a1Bhl5ThJ+FgN7Q2NPg3ysyiSuB8/ZkHIPbJ7
fmHT6qIJFC638gCKX+TpWR5NLuy5CCNRDvPPDbgQK4hYnhIUqFnAy/5XaFgPEVRX
lpKsNDiqhAa24ffgwpMyqn3Qn5LxLU3CjTk4UQkUaEZcukR2LcywavYsiWB50uWD
qUDJucXGO3xYaD/kO0FfDeP8CzHkJSsHG0/QVpmnkgx2nyPshyhdrhR1/qSVYkVX
VQQpxaOLdcVdA7Ipd6K349K0xzz9A3yLqyE2QwGmeeMKU8zdZOFcGoyRBLR7YWg3
tvjWtvAkIXYUDv6F5efwRcdUgElTGC4hpeBzAczqKSEzuc0O5cv07BbY3OmkPM0a
xa1DQNInoFCZjjx14NQILtQlhYUE1GJXsmg0eCgv45RKvRGU7bNfpTdWXmqfGBYa
7InSauC5bOfG/ku1SzZbe/7lHEEjjW+Ohat4u+OgNfhXsaxubELO9qA02R8ZQHmQ
eXeURT/ue/XITbe1Z760KoErSukYx4wJYDelSIUu5jucgBj6g3BtDUQK1ec7L34k
93FcEXgxgEkEu46rw+gYCLA4dYjZUB/x93GUzGNMbe2ZgGvGTg7Iz2XVi4DynA11
MRGSj61Ms+dOn9Xq+0gD1rOio/fwT89ozffZGaYc/bP6IT+IDgCUwpjOO7tAZjhl
otr1u4MQyji1O34EkMj/AHRY7d3Lufj+9CEHIdl60an6lTlAdWYVhg4u1nq3+Epf
2Yxtayl3wavaupmvjXdGCBNEODI/mjib549P8kwFk5ecykgpp8fJRQsOxJhnXtTu
o9Y05DT0UaM2mrcCFOXV1KLU6g8Suk8dRfXnZFt73n0lze5yGUfBR2K0KskzEXRt
lxM/yZBpqBvxx6zaNso0EVArBJxTx8Ue0veDzSPPTsQY4qGuy4pZRpcqR9CBHTFP
JaJzkOmvz7LXYVYlMxJEIIzNPXOQUdRLHgvXz5oQ/nDNfSQI9r/f4u8+VDLwi6m0
ovGnKpvRfhLDt+v3RwQDB0HG0wuPbVLAHZzoEicuVEZj7v4ZhARZ1QeA2DNHmz3y
PfFqblmK3ODNmROs2aVLg+XcQF2+9w96JPyTY9iGI/1LP2zsXinHkqM2YAdjs9lF
ZQ6DhT07sSL56pzZZ+z4fT3vC1DOPWXSv1Wumm1w+Dp83BB8Pevb3cJxx4J9PYAB
Uoa0B6F0/yDuwWyUcv5nos3OL53cE0Z6da1cYGio/3ILoz6rRRy2WWY4sWSBkXB8
m8jN/WRfblwnZQydunRiYyrqXLV/FQhb+rXk1Yh86Pqg5UsNdx7jgQ1jvSlc1Uwq
07CC0ypd1gkFWyj64Ogajh+3tkquYCsqIvmh7lxxdkxxUT8GJ5itom7WQIC01oqI
+BfeteJUwu2VuQ31PP0ZRg7GC/xRKP3y2oUudzG528ZYK28MymUx/NLGXh0KMBDe
ouy1vgcVCG/jAY16XIgzKy4wHKfUh4X5u9achFUf6Lw01M5oQWsQZPAn+Au7bH77
e3Kd0U81kwwmC/iy7m/z4EaqU/5iL1n+b6sXDCEnFtgKeuIfGKgpGmt4Wb+zNcoZ
Iy18wTa6wLGKLCZmKTljBw/x6VyosUwq4gTtCbOelW+yFfm7n4pV3i3XHtV3+jYo
B0qyXdJiO1JkDNxymfv4RxR46m9bSJk/ZgFnlwA3/Tdtr4shI/BEhhEIdjDuGS6r
OsiXDW9SehxIjKbIdN3y5AfCWNrVWwjCHOrjvHH1OlxOjb1vECb6M8onlLnH1NWp
/lNw7lKkwsATzv84o6So9TmQc5cBgmP30WaeuNb1+TV0hwOK1wYlrlkl1FEySkUG
LcWUCmgJva4js21ggg3LbzfJrvwFHnTMC/A581sy4Z0YB+Z9X5AQfkLbZ4hFa7aL
Cnk43CMGaJIObgSwxcC2+iLv0tWLfuwKEPBoQw6omIY03nk7bIwnWANzqty6T8D5
DE6XBoNonxkYy7cRJl8CowHMlx1vwQn+XZs0MdEp+/z1vipx4kIA+61+7JrSrFBm
DFyTR7Ol/+HYDSACYjCduangxDJlGW94MXyOkzvYl21FCUrwa6lwstoIkLd6skjd
PQvJ7uLGTT98nQHq0AzBM3LOXBxniNjZ8AjfVZwcc37K1+dXM43Knyw4stdLb0IK
ApkgODG6W4AqTpoD54Jc9x5gE58354EjgsMPBobzmYp41HOkaRmgIzTYpXOQ9fZY
sNUD7TirsyTZHPsXlqQZH6xxAH0OTEaCbdDavA8uhGc3aFkMeB43N9GfW90slA49
6ArCqo4anZ43sbTrDkJyuYDRk+DGMVFJn/raKsqC+hySe/zn5D3VL9hmT9D8EDqZ
LC9/8aGLXhnPvNh15/OMRsp0klbQFLFqCF5UBxhXDvVbNpP+XBSwof3gFEQPlVe7
+qMfcz1g0qERd3XQQLOmxZAqxiVdleMKYulIS7mBwcATYBDzrANAA/XaNYa1P6YL
ocgmg/dpJQf1c/vDrzpJP2Lmgoz+2aJIYfnmsY8HFm6xC7MoU7DDjf64MXECMeuc
5CiTJDZ/2KgJWXfb0He/Bokbv28nMzLnYSosrSHemcytw4BYbh6hi65JgKP2urz2
2QREbfnqyMYQDa0WLgZwZaaSx/2cSM+9EibQqayQ+ETdXxzsMCOftq1W7hjDrb4B
1eeqzkcuxo65tJjARUy9E9/ec8NDI7djjpeNT2rcZf3J4pAKBZLumJPEXfDfzjpt
0s3ad6Kqu0QiYlIQ1t/4nfW7uP5AyiKV2sIpAI/wsOUzISND/yFNdoF5nuEDa9Hh
qGoJxfl48JyVQKtoW2pAQ+INhQxJ0JTVuyTSvai5K3/KD5Ava9I8whAggZV22Af+
wqbhcz3IijzdepVWOAsnqSCYDnZkeOWZmwLGp4g/RH9fTT3o/Fci5GVF7IFArzH5
rgwXQsdZVNhQa8YajsiNBbtyi2J4vysI4IGy684xl6WAey6Yi9N4sYusrLf8Hxxa
9jfadYnP92BF1JMEj2iNzgfBX1/6xdkWDIWjXu73lfdoXAT3AGXpdTXw9vu1dP9s
Ka7wikAqxRgjqRdhNJQBahWJ4qTckJG2odp+qGWls2ol2h4atK7M+aL1EHbOWPkB
BGpSKGZvjOvhzjx1f/PJp3aOdDpccCiq225m0xs7mBifbRMQELUfp3SCcQxtdCdC
GGIyYDyXJAtSbEVIIaDDnLfLKv8cvlfCq0PrE2NOSi5KR1MGfBwO6HWs1uoVb9+u
EGCj4yr+AtM01U66OxTo69z3gAwEwmRagUltJgDDdsz8nymE5G3ZLtm16hm/Vd2t
MqqeoKtGFz5RNXjruBfgQ/YO4TnIgN2USt/25YmL16iEXQZLcPVhWiPtXbkDEf1s
GZALuJgAgQj/PgGRLMnwtKbIXsXkYmynBkz6I65mqa6AkvyUrAcchyF5UvT/Ln6Z
y3zGaLpyGvUA1NQWeWpBGP8MVxEnjDrD2QOdK5rUhcw4qbNLOXxOopETW5aJnmn6
fHpt7fho010QXxWhhVNO8POiA3tKcLC6ThF7NcEIwiSZCLsx7nPceGqMNYgjNE5b
ReOd+CgbeNB/WiKaP/BPtEePOW0qPabrlPCOg9b/GpLX7TrQuFeQDmMFOR8yeMUi
unb7PCbCmv3phYizxr6A5SeDtWoATcMqcY+o0tjTuYZhHI0eX2/9uEcjTElBrd07
w+ZpGpAm1mGm9HARzeWrPV3vWczdhr+MnkekJRAiMbmIkN1S+UHfEOYfsT+XgAtM
NlnoHV7QsL839Y47ZJeLK3+O8yc4K6kzHaeqKJ5LLc/+6/YgPSxcZou76kTh/LC/
e5zN3LzG7xqsBpKqih4a1v0Ty6Qax7PgSCrO37BVDx80motpuKukj2P6qXmcpiFW
FewOU0s/eBI33pRXKrht0b1Yw5CeBHuF8IPTyUVDh36uS2XVodGByUFtc8T1ynGW
hID95V17xF1nYCZ0CZRSuY0/54+kLvey/pTbmGZ4bCjkqXypgI7ZeRUVgJSM62yn
lIuRzj1D2AWXco4dsMA+yXtCDB4GQOCPkF0uNBQhKgU40g8xXwAA/98H9ZmR8d/2
TgL3Alq2sNq/K6kU3KcWOXvLVceplv6gIEKekdbPE1NmIy0c8ddaNBaT2BLzQIGg
WrUQQywOWAl695nsbRr61Xlm165dcSKVvD1nDz2xG+xcz7qMaPNXO4gsHz1YUoas
QYaKe9SDRbWrMRBY1SjrPpUaMqLrE3ck6OwGb5enwixN+ilBoY9coTlUiQy1k9WH
Ghjy90yITQPZ59RE0u0bgvsqJ/7eEjWD+jn6qZ00qXzCrA0yPAM9wA1yT0Aysb4R
kNRg3Hsr0arcym15JWBWHKJOSJCDFiC8wygHb7Sj6LQNzUUAtc4pxxW1H1smnbbR
4tWPuFgCORtgQqYvaH8RkG8sPgsZ9YzkSeB5z+5zprwWTM9Tkhs+Rq2NQfBnLnjO
bjhf9jUK1RutK5c9Qh6gVZFxgvHRCjUY0GhCNLMHHGd/B9pKsZRAl1LlJTlqlp+J
4lpH+e6IuAMhg8KYRbacoh0xP1o2YvT8zymC2ssmxTmiWWRFQMwTR9fPoc0VOTLz
QLr1OEYAhmLg6Ar7XFjQlOvWwUMqSPwjkaLCoBsneKPCDLCj6/O4Yd1GYOaxwvO+
TkYTbsGyLEeob/MZAnf1k35hX9y+FeojA38OSvFFJPj21riJ40LL72hNHAOXU9iI
BjMBjqyCR1Rjc1mmsG+SVAS/zkDlFm2ZRhsAkvAfWJYcH/Trqt+SaTshiQccSsfo
ZzMF9NqF7K42soNGL3T62vw5Cpk9BPG6vbMetPn5eLVgiADuimCFEroFGtRxZRrF
y3ss93CeeA+YFeHNQwJsAkHFg9QP/nBvLgiT56YbrKBnd3V3120gpz/cemzk4fo9
DeHMZKC9LnId83wsUC0sKTDkNwLtAM/tXociFPTdCQyh65aE7iTws40wIMk0W8t+
ZrytoHPeK1ajpEbhLxfGJD2z87wnn6T/We4Q/pZjzQFlJejUzUR1RL6cnhtferE4
hROTGXhZJ7GNi845aYco/SER9ipwjWyslXwHgV217OLccJ1F63/YhVsonNoArpcb
HfRAD0chUrCHRvmhGoAD0IvkRftvokHh5mObcvf8ar9Jatr6CSDl4CiVEDVInnR2
x0pmKjXkzCg1qZhdHWjITTVz0IukCK4oCW9B1MNbf+D2JGbEmDUYD61CG9TvLAva
ee9Ktgwqy500Fi0f67e7vpI66xNabcMJCn/hy5xAkSbYjoqFIrrRNd1xBXVZIWa3
JHDJffvJCTRW8lKYZBBAiDYnMMwHcwNgn/4ipRgGsznZbb6WerEgkGEnYSh0za6p
Csa/Z0rE57wSjOwvPtfgWKO50RDt59wh3H/TapslKg3RZMZLj9e+mRBHctWZO6HU
OCISoglHprrBVMO/A5255Nuu121GGi90yPDUpO8s9deiN8gsrUwNrriKBeG75lHT
FIeSEC/rW3MDZMqbNHiReTuFEvF6PZ9NFr9xg/CLmxQ6sc1u610V2BEMy4p6ZA0I
ISmaOoR/tUQNCnsvr9Z9HVIrB27aMXMCznAvAUrG+Im686Dx8CrcK3vHwhbTGyAx
pw0IYNGwlzmgDO+X3VednfXX5xSof8Af9hh5eDbkqhy+TVkM991RS1exP40Th7se
GpWyDjkZk/+uQH2mANZYn1TWxDCqFgdAGQD3YoQYCEc=
`protect END_PROTECTED
