`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1l1h2Iu6MrtLavpiHjHD+JxRXw/BCkSqt1lTFdBbbK5Wy39sHxS9XdriO6RaCrg
NSuPStEF6bmsQKnDxFva02iDPmgygRNO+012sa+56/k2k3DyU/plShXBBr1Xkf24
BZXWsd/pmzv6f1Vhz4at6xD7ayumavMEhzRumJsPrEasQQG4UjtGY5sONWVA8Ret
bj2lCOuBnKuArg0YzIyIwH+utb9E3GuOEv8NCMcO2awl3ToHmpMKe9bG99aBbvZL
mLzYXI6OtfrQQlT2eh067O3RgZiitUXct4DwqArmMDqyvWtemC5uDiobkFBkzBBk
yjG+q1wZBrBjyQ+eOZnSH3pmNj0ZQ2PLmo4DxpXdGoL6s6h2tMg79GsE7mm15VqX
6B8NhiEMdlGLBBdRO3ZTmAHGcXyJhYmkWZUTO8tOhvAbKHCv0bvZf8J9KWkoTGM1
2LgG4wl8RsZfqcsKAfH8c22rnZXV/FyALXetelZxyX+ACR5xcaAYyb+m0FD3cUWa
29VE5GIB+KXor2L0xTXPQqwS+QqBUonhjO7O1LDgaQ8GcnfT5MhW1gQ3gt5zMG5E
U3JwyjBIjz6gGSVAYqlfGMiscCE7IplDqOHCgg+Pzv2UFY3Q+xTip1UZNFEVaOCt
yI2lh/9SY1BFSCaxNJeEZlFmdazSOeuKE+5zmD9BrCBKYzuieujDYB3g/XoQr/GQ
2XYavU3uB8KiU52PiZRaZ1FKjUpdK85MNr49LSMjxQFY2Vcqi0+9CMNKe6pFUTU/
Ls6tfaGClGi6OEjn1Kmq1IZIXRiJ1cC0HQDrQU5OvVHfd8ZQl83js2FkuNA6tS/V
/9bhr1I4+lRsQ+BQrDrbUl2S+0bhCdl0MhltmrfEzrLqEc01CyMPcm2NP9RiSmbh
fBlOCKLc5LW0KgyFbqlxOlTZeTW/xr1yB8xsdZI1YsmeeqQfpTNk4ASiZa4IwW1k
Id5d/Dx6lUn/n4Jk9p9xvhfPEmkP5NZoXT4IbbQ3lPqACmdAXfV/gDN6XLND/5pc
y9hM4HAM987mevbRehIOiYaP9Jwe0ziF5g088CkLpCXfofFT7Mu4yDCJk9UFCoQh
1ReWAwZx55LNUMlAnMsDje8zGSpxWt1fxE4r7VnPQVHkRtqlh+JeeORnoTLXZ3gd
wOY+3DZmvEODP2j87fiJEnWgaIEDeh6+QxYkx+fInCVGSQFrlxdDJMaTzvuS5VHP
bhtOERZWpPN+ZZCpI9kMahqKCW1+oSs3okrp0G3KRXU9FcyyWJ8YodW7ZXzyjY3b
SYlrIorVRpglOB/v2B12ip1JRiqsjGqOtzH9TwYsTiUn+Arv05E5eWgLJaTK/bGQ
lW9I07sR5vdXSOPsu8IFQYwDllm2VKN35KQMcpnAqmxslQxnNjQUJnaUEaas6RyS
qzayU6G21T6zcm9qzF6tpamR5h5J/ZOGjE7WT/PwTEXYsvV0xvYfadeOEJs14YXm
8R8UlFW8xO/SkrOOBdhS8w+jqZ3pso0Lz62bdUAd4+aluBHxP7dKiUE33eyXSo2Q
`protect END_PROTECTED
