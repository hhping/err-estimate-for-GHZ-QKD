`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdCla1S/qepb6NLuzZ91YsABNZ5ZEcalagNZ0LG7/ghsnGA8Mw+G7CD9/O+ZlMlD
LOK8O5Az0Q19ac9a1nF5vH1LkV48aBxWLJrI00FS4AKq1FMjtx9ho8Pr6Vt0B8Ye
fihG/Lkr63ThlkLOremLwDD6FyQtBhwdome9MutIIT5uzkYUGnY4CL0dk2l65/xu
TCPKQFvkIOKtDIRMphKCItYRjYFCCimL/xOYGv1L2MEwtRd5fhXo2V5oQnfi9CSJ
E0Goi7qeszFkE2h1qo1CVqVJqOA9hfjPDemCt2c5ekeZrCneEfiIk4F7woNsOSRa
CJGxLIPzVRXQCteUgVCeMTENErqxX4CZWXi2kNHcsUF0poJp1brgQy61jvg2Atoj
YNVXqc8xB3sXwCVfLj95BLn0Jqj7GyQhSS5nshUqNQQ/wygCGZLdvwVP43J6m1dw
eyZEKV5hdYYCmpmeGqWTYsOhG4JCBiEEBfp7LxWZGIEfMxl6rC8sgOsgtCZ4Mgm/
E41ANE/mxAt+CEZmvEAMEJkWUBID6xJpaSyXgZLXV49cK8EshECnJW4a8GiKYmg5
2oZ9MyxUw0lWrxkrj8ZFlBh22SF4I3MhGUIlvYacxp+78hJsah7+YKhG9QxIhQ5l
dNXMB73IiaTf/mIS/qr+rbB0YEkMSEU+c6oks5PN+ly1dDXpJL6rhHLhH6fhTQL9
Fl5N37ddQesd3H1SF7D1TK59vYzZk6lDcCuT/RVC5iEmvlr5ktxK+XpQ3gFdBGR6
9Hme5jKwVSN22Dvfqtb4jqX/2VmeHHiQyPQst/4tlcF9dYI+wI7ND/jt0Wtckn7g
axCOqncL0XDxc7FEHTAwBTBmgadmhjHqEUFmBUr6sDMUAftIfEUzWkBN4r6qSNT3
ozelI3RPpPlZV0p9JmFoKYnfMi0gfzxL2vJYAbiM6d/tI+Q5WlEbkwURQK7M4T29
m8OhxMd9rIJtBs6iUBoUDgtQdDO2p+9ReeFK4ekBQN59NeINcIxleSDkoCxYLyo+
`protect END_PROTECTED
