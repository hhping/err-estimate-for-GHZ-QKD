`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oIbtlOTZY9PsqXJhufsCfmCA1DVInUzAcoXd43L8r6lvSlnBIibsfmrdM1x+Io4
vp9qiAq3tvLZKSakhPhnKsBZQuv0wBGzO5hjyt+Dd9MEqCvVjIKcM+TdjZtQ59cn
QlyrAYiGKhOahL1AC1b9zwUNNX42ZWCgvyVbUiHFJhYNXyhMPTNDgnxheNjbmxHI
HVMG1zeL5ogEO0rCfOqldjOyOllocKx3kbwMsu1wkKGrBbGIaKWxhEHJoYgyNiyJ
cuC5Tc6iH18fClAQKEwyvfGBtsA85GjKvbEqiTyS5Jt5+2vr+cPsjMDxgyLS36ux
sFHcpSf/mhngCpCdwYIsQNJ5q04xqrGp+49wJpV9Vrv6ERb6nuIorjSx6u0o7sad
mVS48qTQpZiS2TeNmUUSJKkHWFFzoTEido60Rn65ARKcgoMTZ5kifLHDgshi8xw0
8JDmEUdyHR3IFw60xbAcsa1SK7E8K8+0WzsdgTQOUkAJOhMppNSrrrjg4n6qAWXG
ASqhtJZOHh5s7rv13h0FklH70es5HNGlKryb4zO04J4ZBwe42Q76omseg6u0DIe0
kzCqiCX0Q0Xin35CqjLi1zfDMIJZ9/oDiwBX3kyrgP6OEz+JoXfnjGKQ+veOdkjx
YEb5ty32WolrYskjv9z6Wvx/7Kz9h11Qrq2RpjN0/8IX9RmGEw2vThx3BGmLg/w4
WvnglnDv65r7LzXqfkoiZ8paQqWxYFsSKvYGnVIMIjfQo6gihek0i2uEnkgsH+nN
fu+JClI9xQxamg6EDeDlLzckQGRDe5p5hC9B4npukMhGFyY0HxVeqIMRnOhCyAb+
fPQXWWbxeQ5prsRry97lYYHKaFcAvEXMzpZuBnQMT3p1jYJPWr2PyD945dNmNlwm
kKyNUZLwAhKZYseJc8J5cUbGQcQHb7ZYgW5N7b3z6Y2SC+wm9WOZYQD6jHUmZzfX
wP8hPj7Cy4jR5mItrUTtHBBlVHRD8GwId/wRYYjcZeYgWnpUpoY8s427V6unUG8J
Ezc0U5nRbJ4byjvHXqz2cvP8p2I802/a83o+/kU0pZfHrFQxN905Hq+EYAUGRUSE
2FR9xEnF2uE5DBidIKQpRUYF8WMb4oVBuwg4SMDv2yydvutQXeiU0mrdTiM08c1q
HTHuVQYVoaXxW3Dqey1vHA==
`protect END_PROTECTED
