`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nwm2gqjoSf4Uy5vC5X+RNL1Ln2Hm2g63qXDgx3/VH5MEyhT85ke+Zzw+XIrVGL1m
t3pd3s9eblDUzsZjXPfi3OLud/r6sZEGlnqjERTwI3j25J5v0m6bdJBarCRK4s9i
B4M/8D+mx4WMpzePvrjnwlaBI4gGHhFW9g713HTiIC9h+3UHtFdOxApspgmp9azY
6eB7IKyfUpuVM8WXemTfxkAV4844U/XWxfOzsnpcFGoZrQEXDmX5q1vf7F/gVz4/
ZtMBf2XLFHEdoXHdhWwEHqp9EKx7CbKpM4MOIWso8/RXQZjFk7qmjbOSwCTuPBnp
hym4fLP1afQWYVbGHNlscEP0J1vNswsdLxP6/FwNqp7qelr6Q0No+beTQWFHFn2t
vCkGTLbe1OzmFFQD7Ai9WytE3z0xAPDSkBfxjE+jytDKRWPEXq9utiaTvrlK82wC
tPmdDUA+BQb6zg30GbdzfcfHor/gmTwR9CiFuhNWXnq8yh9vdfZn8+LGcarygw10
g9DKczkOdaHnQW9WMWaiNa5mnrpyxdwnNVxz+ardz0xZNJfkZHIqNaWfpGDfDPY8
M5ILw3CqNM7yo0sW8eYp7PeJW6mdPyLEcGUhk7n64avu5yX49USxFUBpZ2AEL1jR
aSVnF/S61mOIDqss68zyrFBOodgJROVBsvgHEYX8yB/O2xqwO1+cTtrmt0alERd3
8+YI5bsE/jdLBgCPLYYTFeoLKHzsANNBT8/4cnmxED8KlKxPG9zWQwAYDYTGblcr
GZuSzahpFxiJJieN72HJ1qBtLT7WOt2W9/e/cw4F+06JSVWFQ+OxX3repkFZ0kWF
eKgZEsYo4pBzg+7ifSoWDvYPIouvS7DQvijwRXgDmOahYSli4WBOTeGWiBlkkwh6
uZ5/lFemeufaBya+7SXKx1/IaPByYQSDPb8lbmOU3rLsuSf5RLeGqP02uLU5UZ5b
GWg+jIkrHnF71dqB84HGoM3LbkAO0zk8hq5dWCOFQgRsZmw7RmljfL2ufA9UCSbQ
M5derSScabAstp/+0ySLcQ+WeuAc588JSQ+d7l9vIcyGNRPLckOIIjnnspeMg1fy
W5tF/eZwbE035f+whEtmplBL4teh8iephVxOQXswfQp3BbVkkm97LOppBG9GWI2M
ZKFzq0J5pw14e3HbG24AXTWrL6C6sN/VYTPpaIMDWHQzVZNNdu3tlvPtL9D6CgIL
Mti71ehpGq0IhnwIuEL4R2kAEiuIkHRPcmkGiylS68R08ObME9QOwcLLcUvx6e/Y
7jXrV4LXNCWqp1Wht/X3RkVHiJ85RXa3/KJzeSM7Y3alhYN2EbdPqBVofZAUKNtk
f1jcVH/HyxvhEUMHt1fTBQlryBeqo4bdOl91YjwYpZp5kfSRzyCTKSoue3zo+XLa
g90qFVM7jnVQi6v83YOjVEvX0nriVYOmVRoQmjBbTHWMOaF7SfptsEuz0B1Wt7RJ
S2HatkVM8Rm3+KOLromu1zqAO76M5LrrB+a7CcYm9ZiUK1hezJnNIXlLu+XFvNgG
E3VnWljNoZWxlsjhDgLzy2Mo5+faAKSyxaXFgkW5p82V0uflVPJH6yJeE7nwFaXV
6BdXQMogERzL5g2GA8R3xq/emGsYSzuBYT/A0w5Psw0HCXE5GV+1jMmRC2VI3tc8
AD+IeUW1dF0o+4Ws4tizcy23zdtjigV0BqZWVSowjpmml/r0S7elO1Wpc45b6RLi
ZpH0xTsaJ3qrOxWaU9YWaKTTr9q+5SfoC746/t4wcHzBExvAxEwiDwUxsI5UO58b
aXON6p8pUvB2CMD0oY4PGJlTAmt++VewOuKpNcRm1tTD+cYTHd0xQotwF24Ww8Xj
ObddMaJ5cPn+cJCNcX//k9F1RlXdD6T6ujEwwZY8sdzFuQ+Sa4/4Xc2LfL2vC6Qc
Vg9aNpBtUvr+anc9sqshg2jm6NXd6H2rUfIqFPm1sDwdFQOmYwjiECFJm8TUTi8I
sBxOADCgIfQ9sVh7vEwjLULgzYgprcXF9j1cawziB4q4LLU/NOVpewYoucw/Sc+A
2dhMyyPuGOXE+g6B77F0htWnrHydFZyOcRQOageeUoSviYB4lkohzhLTOXmdqDqS
DYgiC2GCI8/SjtHQBJz0HihYyQC16/e7neq8qHdhlp56ErnLYblwiijVw8wwRWjJ
Yq+dKObkda02eeLanaUSpQS+J3N2FS1Qf0wAfRfA22gQ7A9KTHUPuBfUCmvbbMFD
Z53pK0iX9yqJTNVNkV7Ragsk0hgy1WrrCPutqQQcwTWEznT9UJX/HzcMeUeKSUAL
LdxTZCwmKeLLXpsBPwB8xql/9VGP0F1+eS/x5M0QkloCe+aY4O+8BjmybDyR/ZWE
eBboR7BDIPTW1OoYfJ8czfaneQA7UnaqMnlJInEnUSbTiWyVjhxA8wWtVw3Lx3dJ
`protect END_PROTECTED
