`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjyJyyTMRn/fUlNDDTXT9gtwaAPrJaCZTO6GGvPw0gJBKdmQO7/smdUYwrvSD0vk
t90oPMtkUTePPX3+cXHZ2FEAz5GE7OOMN7eLhqVoPGujtU4Q24UygW2dXd5IcPSG
rr1m3WDLQQAgaU77pPiCA5CK+c438luHGJbO8sGOk8kToLc501I2k9noOFczGndo
KrloPsyz2NPc03X2tPbZ7W3ZmYenKEg3RltOPUIhf5VkmXCBzRMUjnpnqhMkfTZm
Uc+QI2NRTyB9OGRUMh26K6GMgWa0pZbfwqYX/5SQUjMheSPLdCQPlGKH4WOJ1mLL
MHV828gGjqEMB338iS2Uiv8ZQkay2/hDapnQ2FlvpeCEplxA25NjStX9wVKN/D88
`protect END_PROTECTED
