`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6a1FbrLgp5uHkA2VgWGA7JAPBn0Q9/t2DLXOdaCtHUtrhI7kzcrVJcwIL3e6fnQ2
pyZvJxFrX/ciJtjvgioWiQA6zsGrfKqqTPz1p8h0CUZfFVlyDMqH7oce2tJXu5k9
oSRxaHHD/qO/7EDYrr43DdvHSdtPUoc00XlCYV3bmndwqxDUSNzceh5yoUUycCFJ
2+uP0Aux0bPcPsoKNPW3GF3/p8Uk9cOvWZB4sDJUJ1bVoRt8jzAyo1iw45GBHNC+
ubzsyXdIUKLobAxRDsY972qglkrakl6yR1DoAPo7l8NErwz/083gPirC2B1mviCq
/57CSMSkEOpa/TgTzk5hLJxAtBk7SlQGKLw3sNg/y1NtHDWAU9/DzPefT0RdqDnl
CF2pLB1QsaBDGIgLWy0orl0kPh0Ee9LW2KqQqPphOBLndnNW9o7MjNTNfEx3Dw2G
`protect END_PROTECTED
