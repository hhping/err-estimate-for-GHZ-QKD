`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1YWi0USr+V/hs8RR7ZWao4487bjypjsmubewDiqDKvV8l60yUHAARjcjfGXdM4IO
qhQ92RUwzmHuep9C1uLbA0wZZeNvl97kaSTXYKV8L589s90xUalhiPDPdi0dwnN2
vYrmaWLDGeGDO7b+zZUl9fag6pb74RQq/lGlAsj78KSAPF5wh2uqOOsVCfcAumAU
xuHsMP0H7Pd58EFVdPNAWucWmWPx0p2l0EralTyMS/6AD+sZ6vdqk2Hl5n4EBHyO
/TOIXg0NtwEMIOJ03e+CS/GlOfEYuyr4ZhumcKupcP7+iOIenZ4jM/xir6H7QKhi
iJFVo4sbvumMgXrf+VzTik1BfpgZWPLzfIX6NWjLyDfm5Bnt2iCEEtvP9NtG+x+b
azL9Y3Xw+bVC7ccIHQSs3EMMl3BIPrf2yqaiSs70uN6OtoeuGNIaw8Z6VV6RfgjQ
9y+1Xk5q8Xa5VtfLlcr+vvkTwSNIfF5iTozpcSKNSA9sB4zzLkJMDa34cvNbmbuJ
XKhp2qAHv8RXcm4Y42Jv1FvWhrDjlf5YyH0lTO4M83hGADxh8ouduZgn0+9bQ54X
CSBRI2JMdYkK8sYLdLwWgvUSnzjWsAVw+1iurvq6OMS2N+jWzq/khcBRJZqpmcH7
UvgRFOqs1w60r3NO3mWJPZjUMgEhEnMhT8TskWtLiOd4ZOl1fGxp2FCTTNToqS1Z
gGSYwPbevFHtd00b3KfP4Zgit5oE3eB8qpckC+vRiwZ9TsJ26yYA3kaRlFKXXb0Y
7T+UPXepHK14AeUj1T4e83S6wGoyqd5qZFObjBdc+8y86rWzw5Boxhou+WH1HyvB
JQGQGmG5+KyJwuovqly+fi7OU5cs5meDSnVHWFy5c4mBI3NEsJ10G9GRIi5Sd4Ko
8gZM22tJXTU3nUsWLBPng96Lj03oPd5Lro4wy+1LadjRwM354LD5F97XgWzg/rgr
k65yujoCIGu6391OrAqS29Gc0t8IvwjE6JjSSRQRVWCZXcYygc1X9IoIu+RCA1f9
7qbHisq9XfBdvneTxQ2C8HIQURPy1m5JhTOcSNCI+uY=
`protect END_PROTECTED
