`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDegm2jdO4W3nd3f02TJhUyC84Tl3vNk2OeMGXxql9F0LLx6oK2pVT+A9V/1iVyR
SMamKr6M3Z+suyT01NzmFlvNLcblz2t21gwy03H7b6Ry9sruD9u0CDpu6u+/iMxY
y202zCxWJf8O1RjUftpuh8dtrD14+9x1nOOexv7Ps+tzlJLD2OVOfC4NgEtCsEok
PFjaDUfRkKUuJKXFF9ANmxLEKxk+VJ29QegitxgZ3xeWJ0qnCbfsfAMm1qx6GuXi
G9k4ApvaLemyPVkNMHtYH+1b7/PNPgO3uEljTjCa95hDQWQkI0yx5BVOglka4Ltg
andk7aTfrh4dRt9LYQ8mkpwO4de1eUoMSCm6JnUcQNIfx2fNtSpf3+xILtvoD5Mj
HlLLuZsA2pKvPfpyKdzkh3jl7HQyxVI/lJePToalLuNOMJG3vhHDl1bAOSU1OFt3
g+RqfbmCTph7Rg27CWMuvgh5mnwKTLXhkghQeplfq4h00GX6nO0uHbXiZsddK8LX
Jsw3H9LZIRxhhnS3opeNWyLllCdnhJmQ2CXCgQPa/KSLcHsKTku3IKZ+dczaAnSR
bIvfSRSGe/L196E9nieEjXloVSR0VZ853YaJEjJMlYsGhJ204idJQfvUpnX0VRB7
xJbdfsn299fRbYU1+AuZ9WsewD7ebpiIiCzi+SQte+Hrh49EXRpiTiUmFaagwTtG
tosVJoSBCVmpwhjphtNn/JtrsFtUwuXDbGYu7+N0NS8AytgkKlN/0JGu1VAJoTpB
H/QqYYwem0ZrvnEJkM4u7vhAptK0+34kxkrxA5bbpHLXyfbZY+VXo7gxUfjKWnDC
B8W4ODhcvjhCkvJK4xFyilQR43JG34jt9pQawRzJTVeD0VpJQTEACiHnBGSxhc7W
w7rmqnAAbrjZAVoR7bG0F9yrV7FeNTRNpYzvCGwodQ7b2NdjgvNtIaZZhfFeI/F8
hkFJgy5Thr/K1W+BJcYJ2vS7aLowDDibBYxbJTaaW3H4roHpG2wKYro4lEc9PuS5
7dW5N+za5ZXppBwWuiTNiEt0J7i1cwoA/QL6lehMrphi+ZikG0ApIjnbXOXBOiFq
wwiR4lEDFoPFWdce14EygUShNCbLIIYtEzA24uavdNVQzrYA0tOfUOtIL0yWIQDB
mS7EwZ+E3ubuEqJtiP5cNfAeU86NI9rtFqiC7ut/0riegXoeiPBLMBfjhsxZ4mrW
zrjL5T7IItjRXMnMnY7CUrDQCQAYrHhsXAEAQuNCK1DnZtkeVrdi4LaYqsSZaKCD
8GMjihpl5628wB3+ol+6934bg+YRgKAE5gJcif/dO4IQXJgsXNHJKG00foqIdb9w
hFFM7nYzB0yMaahd+mP0mzUfxvZyqk4mvP/fSiSy2EnlRV8Ic/xzk9BrbpSw1tiW
7BnXy4W/2Fxv0aMFsHvBJ4jYEgweskw395lYpmd/urw7ks3xp/hOtOYUS7n/YVoZ
DGU6eBH06yjZDZFMbPCFb5RfdVgHc0+HY8gXmNVcovxhmRzO00DVfovGe+tPh7Hz
HrGogm6k8ddVVo9IO1lNYlfnrFJ/QSgEqkuLL4UVJ3MWz1V5pf+5a2XzcplP+2ec
CxZQsasjI2Da7z7fuV13B6hlfwcgJSpUdNWQ0a7CF0g7qr96tZRmrv+X6lqesL7T
TxmSWo1U3ZLTypAeOz+2v9aBRaGoOH8xuKtYgfeF8fBh8QLnJw9mZmUjd3gTK7P+
X8fnWdgk9pG44R6lIuUHb1sBGIK2RqeIn599FKn0z0G5ew/o3vVHeptPBv14FFhq
I79aijvbbU5WUpQ8g/OLPaKWdhcNpUGnK2Y93btH6FyiE6FJ2QFXnhq/6COhCAv3
3JwV/qxRJidE2Je/zkT1J4te3uF/tWfwRwX1Ovo+5sEITiaodv+GK+fHu3Om5nYE
a3KFrpOuE4hAFUCaCFU5GNMiglPbtG5Hz5NV6ET4TLJRp3JsgyZG3i+8cd9ujg4+
1fzjcFt0r7VVs+Q6/uy2ebxL+gQzEAalBep9MYULmkhvYFJ5a/ScU8W9wkVZLp9G
2K+NqB3ClZUogHNqqC5Scg3U7c4tvcvdQ5uh0AM3pf2i9bVHFTGy2z/41pw3gO2E
1qGQDnBolYR/TDF9uAB0Kg3SDw0HPQUGJ0A8VRn/t7/jU+cHt+M9N7j4qStxgA/6
p6Ggs58lvs1AOaP4V8624MQxOm90lUaogY/ZugBfl0ew6mcS/qjCvOsccuUSadtP
uCIZE6ExfFQXl3eY+HhsQ+jJ8UgZhqZU8yS8tEuNVGuHmGkyk1PHk6fPGSXXcYaR
r/DUPhl/3XOMYhISlQxuHPfh0NyYjEE9AHrjkfSVM01/90ROqTZ1GEhp+M0EuNd7
hX1lwAgWrRcjy7J1faT0HitPjV0zIGfLFG4jtI9VexUESV4IN6u1SIGnhD4alyXz
jc3l9z47zBLjvGQtLG25G0PlYj3U5MQUJXic1pldAwwZJNVDhR9iJCQcYUmlebhV
W3Qpop/0mNieplkZnF9JjB7u1HNQTyaY1Y3QntTpy1y726CWUyjdXN1I7X1DbjA6
PHQa5io/Sgls7OamxpRMdECFpJdFzojFCqTs+rNMlZUJw09q0EWfm9E+x4OcBhnF
eUY+geak/QIyu/8kOkg5wRCVIap09wtk/XowE+vCRDVMCEz1riwM83c4H2IqTOIl
pKaqAjMZiTSe1pbY89R/nhzECGMDv/aSjtiFE6tczYtPD0Ip2GrTE09FXTHmw+tY
9lS5YaPCYZik7LKQmmY0Z81C5JZU6qNO45RjLFM22HdrPdsOI51XPEeyWDZBemVC
FSChVXEv4T33NwgSnH0BGbCGSnOAJwIgA/QWKP/AepRavaKbvdeCMMB8cOLR49KE
T9fIKuZ8awLABpNyPK5tmRQPtcNx+ID238UHD2Qgf9htV5Stx29LKw8DnpJE/nUU
yy2297VbgAXGA0AZlUlB8WqgMnbpe1q5ruzbnJdHKdzlc6WNhc+xPzBG1SP373tS
5MloZ0YPVIrFBP8spLuf9mvups+Zvz0nrNTAIfI8Dsv+sbPBaNZyKasYKnt5ojIk
ePd5gt5uy4bysOwHFO2Tcaeswco+nqDGEwA4+ytl0J4ystqNSVEeBbUtfg/YzQsk
CytEWXJC55qD1EZj/SXsUKGYLA1kE8BWSB9XQHfaMsADp5Jd5GAFGWJGm1aAvjWX
WYhD3+1Jh331qydIxbXFIOEu/vyuvq4nZtKKY7kFhAVPN920ZNfgfnK94P4uAIIw
xcaIMPAAArIn4sW/XZJZI1mvayJu0DPbbsFvDC1n3bnBYw1emi76yRg7qMvsG3/r
SCH5P91Bz6KjTmCFl6Wbb0KVnsXxtAlUnKUT9jTQqXIW5xlfPOwEW+sj92cruqJI
aGF9JdZUkzM5K7S9M3Pc3q1z97+6BupKSwP2JhX+N9zOgt+aY1mwAcPiSdFikTi3
zdZfhuMO2mHQu/dOuJxdkdLjoSAkzqMae/KtocAPL7VFBxpTiNxSvu7KIyU5WV1q
KThOBf5JnDUUjivdT/PLMZ2fPtYwnA8XoxQ7hIlCXC6QUfp7QocynSGfuD3/JY9J
ZCCwrerOWZWkg5UiNVi2s3w2OHBPaB9i4WU2eLYg0Ioov/Grf612ug4C8bQzwn8t
mfBZUMxor6agfgyeAbUhB8zUXgggKSYhr/+vvlXgHbGWvqXRh/BVukwsmQCsBWK8
4EmeKBoRpstspT9dLwFZjMjT5/GzimsVKm1sgUEKHrFRVKjqjOrOfyfpp0PRgdV4
zFxrQNl7G1HWXyAOhlEe/XZEGpbnizl4YNVFo3kj9LYTmTJSied6lYJpP+6cZCyd
0+1YOO9WCY7lctOFh3fqpKsfKdD+tRtd9+IGhP1NGi1mjGpxeIHDBfTLyipu6YEX
nnD3GA7lF0oYmu29Im5+lENnRKHph3QrBjeed11BXN0bisj8Kc6QQoYyvUlu+2bX
j0BD8gCn2TlMGSeXFb3CNWhJ4MkKaeLYBpRwawv669gkTkwOG91fLepmGBOW5Fp/
bBPOP2veBD45gYmlx/dlEo6mo4AMKB0PYEpcqWrgOv+dXN53mBJWujDOEiSMCySg
USW/gqA11H74j5St00R7AVBikJnE8ux9bPuRg/ulrpkMOXAFxuIWz7+7V8zbt5mt
b3Pj8ARzztw8dfVBAgE5iWTjpePESpFMEb24uAfijY8qmwqzgWpF9Ml5U2DFOFH/
TaskOz3FOpa3uasXx/2EKhukSf0J1wE4+6kgYNAvL9Rw28e+MKPsbVUBsjQuwGV+
MeVHebks+Wl3rnqdNT9z0i7bXO92elyj85jIssPR5O/ymKBHUmiqa9Wh5Es7ybQ2
Idt5yvLQLRQjq7r5zhznsWatj1avC/bXLPZZ3NizjyGkCkheIPO330J0YcnSLTGr
gtYqsbDNI7OPH/FNVDn06sGD2uZqG/dzZlByOzANt5tNS4Y9ExVfLhVx97S+1Hbf
Z22FRPCgQeFb4v1YnQJXorhWW9bdNWkBcjv8UbN+IazJ1VMlqHWJt6bB3bfYQmGi
W+5yloFhrYkVcetvrt3UbqFaKbbJpd9khs8GrkrvxNwN5IbVJ0vhJKNm3K25s0wr
67fTR1wrY+Ib97ASsRoeg3zSkmEX3G3CfxZQjVbF9a6iHPCi6i89dYd53zylBZBp
Qiye5gGpmVyMQmJXIkjCzxR075bG2GQHb+uVDaQBGlIG3HhfG6ZSSzL29OuJ+5//
+etVO4btWv0vehj/acstxzFEC2ZqY1JDdx7WjSowqkjQ+T6YZVxAkhRR4qiBomdI
mkwOfKos8LEAIZzS5Ip0LNX80CerftNfFCRAeH3HNgBEeIukKdra/WsAz9OH/Nxb
m9SPyv+30XuwwrKCUXbJf6pBGcGgLjHBdOZ7a6HeB/vOFSkNjbh9lwR1fm2ur17l
jdO3u/t04j/J7ejgewa+QrEyeO1IlqE/NZR0/h3skGq+dE5mYqfhVNF/x6rnafvB
nO14VYchPXJPkmUwpRjB7bWXeuJv3SJ0e32axbMh3k8hzsbper2daOrkHQYwm1RX
Ijj7rEd2CuFCH39kdIaOPcs9bUoPbBeOuBqq+zNWD78QBKFECPj3RXHZAOTaFH7m
GjFIl4UtG47R7uKoPBg1sSsodyoN70y9kQipEjm1rIgqip8K5e276tcUKuBTuuCU
x5JcSWfnrH2fglD2F0EtcbSFvAqKic9aHcqZx4+GIGVamiIXXIqc7iiSHS725RF7
ZoUkIhWcD8yrHZIH4mK26BJD4CiCQDxwLQB5befHbbvT8i3qVtC68pLZNUGKHNUf
ccLYEM91zcYuG/TJaAJ2s99F2Y4L7phNWTont6k81p+HC7JDMu7U5KrKl7SEauZN
8YHZC+27aKXHwSsjryRL0/2JOzY8WcaXjhTw1ZKciAGcYDdH0I0IHjtNBEqrwQL0
m2m29y/kCErBFl4lnVJDN5f4y12/gXzVTq7ssp/+iddiNinvm+FFLPy9xAsEngqe
zHwKNFHv0Vxv/uAtwIJo03EqkYY2xLvpqS5aQXXEJjLdUrCCcYNIlcSVb9ZBfkF/
+Ut9UcC9QYb3O1VbJWuSfyKwJQh/oCptxi7gjeL/kPQc6ab8ubTP/403ujw74Ivf
Yj5pH/phMcVzYaxaeEvLFrGcxgQbvzTjIOQqWOQmDfJRka/HdH+1G0jZF9GQH0T9
MvmeCQ2cEMO/FyajQvhCaJ/yI9DC/IMwci4NHmR5DwMcZa/DiMfJoZuyO3NI7Yt7
GeU1ekYKn20Ntbe/UrUrYbCMhu0RSO9XdkDBATIadxNu2LlsO/q6I2A3KbWAR2qD
7+ihBDP4RSdtg3Vm6Iym/U9TEtPLxKuBkK/U026lrDFjFPe5zH2/NJPSl6HqHAXV
zeg352jmsYWvovN4huSLzHp0JDYwKZBzn0nJ8kR+l78UdifjoIIxaDQJfiQtyFK4
KvtmvbyFtXpTwhi/LSkqCGDVd5FW8WqY13FNF7x93gCsH5kR++8Aa4Wfr6KIwryO
R6A6NBD0h2XomAXnyk51plf50AFhl3K8zvAoa1lE+2Z8dRarQnmttTUczWtOm7hN
r2HOPe7tnov/SvF4VTGdvjGEX1k0vOVhzeABMQO4j2scTBw1TtTEQxwasVckpSz2
FeuKvg7E6zf6kM4wZuJP1T4KshrXsRhACMTrpr8Q1Doze+C02AIB5gYemTemmmHd
cXti8i0fUEHoZVi2UacF6fQVkAgk7VkAUhmpARmjmSF+hY5aTdAn8HMRsCRVnRvD
6w/SM527q5ZmLqWaMjY92eZ65sJHoc1S5Y09fENdWLceIWetIUX6oYcdp2ACG8Cw
NETmZsza3BMaIkXuOqJWvk9mEUdjBLsGu2yTELYUcUeuwpiH/nX+eB+pYhknkmRX
agn9lFeGjrQkt2Gtd1oU/iNYL1Pusjw52ZZ88eSvtid1VWeXuq5bNJKNdrPLUJbb
ndr4ZP8mRoWYFMVEK7eTBf1531LYkzU+iofSrnHZQGb072fPxTOvrFKhGBFv753V
svdqP5MI/v2kL7lF4uVbC0RVTZydbmt72zhrPUZ8Nbfa8ACdUK3vJUPhoebPGDu6
mosTQatYyB4k+vatPvsDbOjpfrz9aFTyhNVO4xUj8hyDevzDU7d2q2cxxW4Tl7wl
G1rYeGym4yNAzlYfj5ezkdOy86BubBMxpZp5qVxmSn9KSWtRy3lnjiFfMbW9BjXk
uCOge+/o6d5uvPnFtd1LdzCzype33h/xAyanXEiUAFUcXe8K05giST2uP5XtDgLh
ODWqzNy1+Tqp+XErmsEscQBfBTOgN6lACgbqn8aGYBaK9bA+0V3lh0gqkLgxH0MZ
Qs+h+knfCksv94lFx/c/jOvGuPHhy4gteO4BQT6ulgSSFdUNJmAPjqmRszIZeLoD
BsdFZgmgtsxhUIpHIXTa5sP5lQPooxqItuUmS4x+jfbIBSX0IPlHtgE0gTys4KGL
dBjgCo0WTj+SgIqTimp4HijeFQd8fYbDBjk+VTYyFioGrgOnhwXmQshIpw89W0u3
XNkAZJ7irhgDvNBiVSUtY9yncuOEZFRyxahI7Ho+fkK8tpnuKoz+DHFtYVa4BLRR
McDxhTXOIwT9UtGtMuu8GnD5vwZMwBliED0tRXE33o6ka9QTzjGvZfYhsfe8HJMX
/4c+nmNvcfyA7pESGQkAdPs09BR4YCdhQ9o4n7DPu5uE1Q8+Fm22CGyHjkYDuOrr
cMLu3zyNVYr8bEktuZvn2zWrlFGDtfbOF6sTm/R1DSgakZ3yGrdKnCcKwGVmz30H
0o8xymG41Qu+Bl6+r8jYpEcSinXmtWkw1qmEwhdm43Y9YtH8A1mhLoCPGYr/xzOK
jxLVfXril9+Fev9n2dQenkKzW/tiizgflzd/L2PmVSdopUY/ytEYRIpPs81ytIAa
MqmuZi33OwXiIy/6vHfRlukzLvzu3w9Q44RDozPlNpTI0QJIbMoU7ICmMPibJ0LE
zf54BS63aiCOuvGlBsrhdIcENdTRt79BKDanyLnNqJSGvzNNyvwQRSf48EOCRAYJ
bGk9i+Hb8QmBlW2oN8zIiYiU4guuJ/yOE0WESg1Ph+gumIigEW6sc/U66M1+jgL0
ii9HJlWW5ohUJYG590NwB9x8i5k3dVXRSadH5JBM1SNicJmtZDhOmhvP2KSGr8g3
jB7n7B3a9BmnMITf4lWapKZkGAKBQtj9uNNq04yoyQi1sakR88edtiqorasLZsz0
bgS2kj/Yygg1fY1gzz7/g+0+zMX0tHL4yLOozQo1WwQ7EsmbYvVxp/B7X4sAnKpn
35I/uJxLWJKS7zFaXzUyVeQsLRg/egZFDUGwN9+VXaPBZ2XzP8IXwt0HXs2qvtOj
r0BgUv3rJrWsOhlX9Ty8v/ow7mOGnRCsMfguHjZlkZdhN1GlJXhkYz7UsTzfJqVf
TD/vlX3RLDvBd5LNCwnwDse3hNQmEP4bjrQMchEfszY/NqSmQQ8qSgLxdHRihhad
Ck7w7BwvszfrxCoOCWA4EY3sSbWwX+eWyjcz4FYzXgHAu/gkXEgFGybtPnWO5/cu
atyfDR5yj1Tqli5PL0s9QxaEiBdZvA8xv0UI83sl8X/+xJ3uPv0GNcaotjvO7QO/
dnhQl2AMJk1Fe7We31+X8vzQ6FdCS8LELjdNvOiOw2rCNris+mfeMh2LwYiZX9KQ
e9NluUJ59/b3S3wM3K+7gAO2NuYSGCmA4eehXTZvDZt/eSngkDlwGCftYAJkQ3iP
hqmhfMxVMM47nMNWxj8ZZErLxROd4HE/5qFZkZ4Sdqkj/qxsJRxuP4RF6G4QfUSm
yv/LuaddB8toZhPufGFW8TqrCh7dsFJza7t2U2zzhyM6/MhLjJbvaf0dais164JO
9L9i+GrTtkbmyaqhbexd7zpJqPTbfFyZZfxGONcC8TOiyZXxCOAXQ1rlk7vxgw7I
j47QEFNBvDt52wMZt3SomE5/TmX3uPA4pfc2+4EWbBUQyy/iGZgsB5kWuMJ3jXKX
XrUbOwgwyxgqvrGfk25tUcNGPxigM8Nk4ayUgB9mVSICSwHKDJVzX/tCFo/t8rvT
1d1jxmXympR6MJciiMOQQZIfjotNqryp0yGqdgGadclb2DkxinuMLj9navVVpd1R
tQDHydCTXe6YMhupMbzL9FjMc4GfvheA3mvaNgiASDXzIBCch4Q1WyDz2096NrPW
jaF7H7tbCZhpx150xoZuw0gMrCfj07PeeqwfzXd/aBbdcB1xnaRQUYkSCrNlx33d
VG4x9T1MXscQNsT/sQZtp1/eJ0oqo7UnrcQg3czXlA1dJkOhSr3mGU53pClqieIE
O/kurxDSkVJiStck2xuHB4AH6yeoU4Q/W2FBZ1ZCJcv9g1I9qm7u6bQCAoAlAZ3N
Glu6CGcZKdWN27g6JS+v5Wwn7THTE7AeDpVxCAow8sksOuCDnZ8iwegKRRSuJl91
Qei2M152aZbcYftAJOa8ZcbA1kYVjfPLzjBSh7CmvXCx5j+k7lAL+DO3YCfvcN9t
WKJaMSpFZSl0fp1FltzCQVsyG5uf/e8nVNmjN1R20wIJGckIB3FEVlxlIg53itl3
fxJEhz+3aWu/skQwyWNgBG+ImoPzP1oTr+vAcaxFonM+RsLC88qGKd4t7lyMy87Z
Oz1wTNpYcAf2NEv6Z7VfLBoMzx6KNDqM9ig+IUfUWaKEZK4YLWV5CkeM+K9MDOWg
sAhIfG7/lAFIc2+vVcVlKvytmoZmUMYUeoGtpAFEMlY4iPAFa5tgQjvoCL7fxLFB
qZOl7SmtXfO/7XwA7zEUYmXn02JTczBNSb4V+B0Mr9aENLR8QB1Z3EFHRVoDz/HT
RHnuvzTeW2Ue0qkqdD9xgxwHKDQk2mMZX9BscddtWXl1aIXO7uI8+PU8AXcs+J4L
RfJkk4xuwkK0Fn5efnV7rTIjeF95wnsVv3Q8av8fgakG9QDmiDLmpP0DQKVHzzyM
5wjRElC355FbB0OaQ5KvrrlIKaFRrBiPXXJSPevbkw34Kjj5FAX1ntSX8AeI8ifP
Fm81zvOvZR0D36Vt7HCGUrilJFt9NudG1BlRovR1xezcbwc4z0GO5WUROj5GeIdI
YriAD5JjfP1/XQNLupRFyBsBx/l8x6RpEYB3b0G/aXZEm8jLzLIpk88CT9WX7UQH
4G2v58BhZ66cEneFWo+JRYWz+80jVskIFlTMm/zOHTt9e1KmOeVhhqvTit2JPdLU
9vZkXVgLj2ilRfMUIH64duxM43bPLgV+6BF+Yrqptt4MLBRn+TGqHzVovlzecKHM
Vbjq2xVWeiCsqjxEcXiyyejteWcFHeeQlkGS5H1BhtIm+m+81q8r5zPPuyEmevWW
o80+yrPoh0UXvPgeVEXqgOvw2izx4gBUeo8GTGSTxTb2+VfGzswmiehwGWneECEv
TkIiYqTN4KOGX0OyYH/7JSrZXkTby9dbKv5SK3keTmd+1eytEzmB9T6FsOiVW/Gq
ietGGlz1R5CH5SSUKdP7oSOdyjowfCKxr5VNpuRhZx01c8f+8kVZMRVj2Vyp4qR5
Qy8rXrugmsOoREv/Lla0e1JqLn0AWGBmyDLOYUp3pVEO5+Vrb3cjiBBznQVzjX8Y
qSWTvENsYCP8v3BBwl/CaBuNICUMUnrk8yAjew8Rej/klVDwAXxzREOVVdCMHApY
xMxEVlGrSEPdL6uNirDYV4XoUZLzzu51tSBez/n2Y68rMQGqF7HtXZmGfYmDtDTx
yPqZkMGUtrv0Q6vFP+atdKSZIWIXf2vFgp0vXDr0CyBzJJ64orhP2ekbPBsg9JTJ
w2Ya7NXYPDn5aursGcmZTr8Jpi9YyRG0+mIqFfvyQj/7Rl/hmt+TiPdHv1dXCXgQ
PGrmSKk3+/AIXdaS06Rm+s1zTJgo0UKbv5RcLGkLYPLsuwzuUsvBYM4Uiw6pDg4L
YpXHQyFjGOFm4cH4hvwLDKLFmb8TF+LkJkTThs9k/0Twea8YsditjGrv5q+wkGAf
nuMfsUtbnNWSwrDPWlIH0rE1Q/ymzQEeawUgjI2ZzXYrHiWWBXutnNiAcFVfarlZ
670EgtO47DVw4C6t3/A/m9wMj5EgGUXCHtGlCX870KFTOPszm2W+oT5e3xYpS5UY
jd2jJDh6wwjsI1ThRTlEb248wDe6RWL3i+UVrhutJ4Q/O8t4L8m4X9R0kivprIlW
clsm2CP4o0ukiRxVjW65DewUJ9zC6Rqme6S2vTwdPRF8SsMjdKWYNcMJGbcBloo8
TNyRx92WWiD2zBht8ES/Mf8UlNM4NLqcrVgPfka6Wia5Rr8h+zgT+pGsxPK3yRLT
OjfPXc0pfq/p/d1sLtLOja1wcMeE5jBgU7Vb0bIXhEqDIkwsluExZtldwLdN2VX6
IH3Q8iZMiK7q5Nap4mgHQIh6GPd0i3p3ftlfz4PoJ9zHckTvrp00TQigp4bTAKzV
yc8eeKd51VcGOBWAPNUVkkBZHJnusY9pVWENoJjSF6HnvLHvcq1ihnK6JMUqx2OH
5k4ws1rN8dTB7O+bYycQKgM+IaLVKOKQeRD9ZFQK9vzG2DlsH7FJDjZ2al+p3OQh
lL3Yc0EPLzH8H6IAKffsQqeOZHptfqfEpohPqI9LsZHRL+lg8Nz99ZfETthr2zFZ
6A35S38Hj8BVq+ScnBQeH9V9AzZ8Zv81WaUiRVBumVkZzSN/5qSDdmHBrKJbpvwf
OnAL5OU1jPqna7nl4vawKrV6dutpj0b1wbK67CiFzoRtm7vEVWi9OBrfgMRcNwIP
gvmW7ti9n9EQL4qKYoqPt+fgg9hiaMG87CrWQCGsMAaDwCiB95P0Mq0ZzK4kuTCD
uLWI506+iq/tU/5lfBVkAKCwm1kvS3qTlN42mDEOr30j1zugwS8EhBcxYbOaemc7
HhifqpQcDUFIA7xvxcQQaCNMVH84KVuITT4/LvgY100VFmeGZ/WjZ4HI0d+4phXf
sAw9P+VVKMJZOyes2MbPeU9ipNaPOZnYAyCHIWdx1eWOMhT6OQSJdDXO24roetRk
bZQSilQHy8ACKTpZFh3w4KA1/mK4KDP4GSYlWZn55NMncfPPZYVEOLDy6Qf5zROc
XEb4Rnr0ZjMPWNDkAIEq+e19fIqCfqTSo4yQ9D+Kn/tFZZVFqnPNh5doBa9mt6y/
rLj5dW99JpIBJRNtghbKYvh/aaKeAFajc0GkO3zNYkz5Qwcbu7+b16n1merKEhXE
sy3EKOr/oGyeWVRK9ElJ51cJOjczpfNc9mjIG1DUi3W+Zh8HIz9qqhBMripVPZOq
kBwA8f0Wy9bycXrY9kCAO8fgHeSjGA0iJRVUK//ikr0FqajUms399io9ktjW9XLa
KSJc6+BO9rUs/NskPw2L27ypSjBMjoxw874lPUFZ4pIpGxtjXdoW4U67vYG8sstA
A+BJZHT/T8a1lPd+qjxQoQmosYq70FbNcBdRudB15BYm4geVuhL8g+OyyhF8qpuz
FZ3D/QGhZcYcMmyPV8hosSbX/hMdEvVmsINE8xjhRkDJsIY9dia2I357MB1GwUng
HS0KhzXWCPpw2tvThOaslAu1eiOtG4R9l9FGg2CjzPRfMqZVArncyuK0x7Y8o1oz
VcMXmkXI8eCsobZ+SFomo39a6XjmIHp5UthVARht0YXi4atH5qsHk0Sm2u0O+XCI
0V0my9Sa8OnV1LiOxPAYuVWGhyOVpFfpXmSEI1RV0EeM51Aq7ZeW+iHXB43V0LzP
6O2dZaoYY4TgxaTqaf0Q5X2hZTjI6RXurOFO6GjhlRk3aXlpo49V8sd6to/QU0NK
wk41sWuf6MNVDi5qoqjf6tFPkmtb1GlaFc3E6xFAmBxzXdfvn6Rt7FDgTIRXImZx
ufXrZvwShlxGKF/jzfjPdBzhLk8VmvKKq7ixStDdX7tH6JOle4cQeEzrtw1cuBT9
vEAQyB2Ke9O1BDFTJxbcnV6xN/8qkN6PMBSln2Dy7WJsstnP97PIhnh5yvjHo3kK
5j22juMz7cQkN6yOq7IL0QQ8457Dj0lzwfmiMWkTi3AYjjTtu9qtJiG8HorG71u2
jZspbr37m4N57yWmvIbHIDNVVUV9DkdrSxQnlubDDph/EsnICTSMPoLK68Aks2n6
Ad/66u9kD84LdJ6p1UvAC3W5vz86TO6NrjdWqLeP7+EKHCvH0IgAFMNunfLe6eHw
yt1SNucKFjuiBiru3XzLajlub9xpIsSfJzp8DbhGKiWqMply4TGGJjtL5D8OTNXD
d/M7B4TMQS0Ih7hScENrgyIZRAdLUIWNS1iSITg8oq3fkePfAVP5M1QRi+oS6Fea
6NTd/riuiyi4hQCL6+f/FT+URQ+3dpFISYInbb2FNg4PzvdmfOi+s3VIs9NR5lKd
BafBfV39xQwEAFpf0917GmxObOIdiP7CgjGbWARWe24+H/a6vx/OC9YRoJXgVCeq
gHAh6CwVqSpaAlIvH3f+QFfG1dVzC+xfQhEFSitJmCR56adRKKQdyjIBbzUOVcwb
o/vLV4wtveSBHFOWV7QyAN0VOQnW4NitgDRv/t80aUKc3ntlJkxG9Tr+ml0K2Z5V
KXVDsuU4oOvIl6rXPZNFIKk6C8VB0O7I13F/lmwh2DUO+9C6qFrW5SNZf6lbNK1q
m5aPgu3qgrwK1Mp5gnlwTn7Ijl2i5btZyuzHxZkTMHc0Uaw7elWyHTLtXNSXGrsG
pybaC7NdIUt2LutCRKDyvT/Lm7jbj9JtOXfeIqfv2SnZ11xMX2KXwgxQcqWPgKG8
AOnHCdIJfxpHoWeDFNZf5N7b0HiMbRzjMp6R+PvwPtgBuB8EnbO7H91PKiNUfksB
OfPQHfqwqs+qusad9i5lH+oyduzBYbbAqU5cNaE9zEgagiExRYtkBy071nrPj43p
VHdSikHiUwieJOa2usp2mS9C0Zdxcz9ksybZN/SsXEydNZMZC3lEMDZV61G6FN8e
0Ls1IaXw039HBk+SVjV4LQKBWApWf6PzEVE5YGIQAAHeSr32srKlACeTUAOnebru
6EmHeG0SBQhMyTmffkUWwVPAo+FoPKPo3YKou/d37FFXh6oKbLj7eFGbv4akq8Vw
5Fbkyvhw3pI9V0AQIcTKtE+Vuw6P9RPI2H7QoLlQHpHbGcqDWOw9KtlWKv4eJRpI
v8RBfgR4FLdFDVesQEiw+Ed+IOecQDYZMgyWHdXdjLXurUMJ9chtRu1T+fI+GY0t
h+BfkRsTT11s1/6Elob6+bgSmxogLmnhqVLfD6+KD5KlYfQAEBbKClIA1NejYzmX
aGOn2J4przwjmClRbrLAy8//ID6Smm3QVF40UK9amayjWpYeiOyWFBZu6MAIjiSC
CIRfpS8hKfQfwrjyODWE+QBV8C20COnP+Hl57SYfwXhYz2hzyeyoNjxGyNCj0IuV
kfS9zJvizJEP32q7qALdlXuzwKkGYVKtTxZyecRTdGEz1KyTcCy75ntMMiTd7fjh
gU/lLz0CPJQW4udbwzLlxS92OT878G/lib3Hgybw9xdGt5qjjXefsnvkK23e31kA
bnQCmtxUwOd72lGb0p7OiMzsaqXGaMyyRR01VMMpk7lMDssdqo/YGCJbKHCUHAz8
BQB6uqoaU7mZEEgpooBsQX0Jz49XrLK4Ex/eW05myU99FZiKgODTpK/0tGY7MAQr
j1MAF3bzmgVQKQiAEZWDwtOQRtkx/4s0GvrlNXMH50D2Z8grMQRSnES8NCYg8XmB
/3T2Xojtt/mVri2/tHJY79T1v9qzmjfscHO+herNGaHQNfEq2Y5xsDImd1Bw3W7G
Yc4R9rNBGPYTEf9MIYADtgc4sCt4ck2+cNSZVPaU6cNmdj4QzC3oQ4I/bXg7QRmH
wPubn1GhP0mWDsmDn75D8X5ktkXBARypQ2BFwA1il37ITWXRBuYrIazOzD428lN0
B7sgpYWyNOokm7O3r3IjUFqXjo6mE3ZauqMXOR7I//71asyLh0UkhD7p952pUdpn
zKGcNd1y8pwD7vsI47F37yeH9QpfWlVcOdIXXZ0bfnX9o8WLeGihKTCaN43Tidcd
ZWR9tFrCO2gXVPhEg4HaTr+KM9GY3ZUIYQgeQWAZqwv+/8GUq7x1S9HbQtYNrVC2
MUXig+QuqLv9Ot0YBxKgxL/Vw8MzSsRoBqg2h4JfNpP1opddjIJYSHVd+y9AgNsr
dvFhNhe1u7BOaG4AwhDli/FgHv/1tpFSVBWg9matp53GEYL44IvGrUOw5uFOqBBk
byHv4qYN5lySsKvRiViargsQQOVntu7Aid+gGrLVhxvcCKWqSJbd4ZWDh60oOvOX
tJ7gPv3/SHZDv60gZ0A+Uth+BJ4KPY1+O9gWmd0LIXR63r9/HPYZfZTKwFM6HIOq
I4konYb52GRMTy8hYXTHKLpqA4D4VVNpkBlRGBr2mRfy+4/RFoPKdgPbRdcToGXn
M0y7ODHYpT6JLL6zPZP2okdVcZWribwEWiibtH6eIVGI7YsuKDvxGNvpRY8WNfZO
0NZdtXxuTdWYXMESQQA52y/rjTREtkshWjm6XCeUwm47eB5QrCrtO5MQJ2k7/8K+
jw6AKD3wwuRb+WChUMaSF81iw9D7CtssSsUouMoX5M5SJZ4Y26+ZoVeLQkUfPm10
6E134NjOZ4qUppHWsS6tyEAM+wwBXBU2wPdGVsNgRxyVyz28V0bzPTm6SdLXKQjv
hj2UP//W3c2W25cu2xGSr8+ovsMG4pN9kYQ0iiKP49ean7a135prcluPH9OeOFyg
gTM/uHKDbL1DvvhjSt5qwSKRJL8mn95kjaCb147oYXXE/gMKoNav99uZqMJzMIJR
e5pL2mWuVJi0hGhpJEi400FRc4nHU/hWyB8UsG0XISrqTMR2JsZnIsyL2V/BwUWe
Vd+U//YUnreOiAR5SNaTR8g/L5zHrfjS57F0nqm0f0Z0GuiyRo2ZM+esJ35LCrR0
EWhVD6BVhxgDM5di/vykYJaiMkKJeP3l4D8FIvfZvg8aZemEc8eq/kOOKnu6/NLS
OKQYwyKrlMkUCPsKm0RXuKzV5umTDGFoVSM73Pj6B4gzOC1/QrAp2ijCD5QME2GN
xFXgVmnWPGz3WBZKol7udDIISdQfJ49BZCwuVjMSSEvkQHZF6e+GiWnOwxI/AHQ5
JHWeI5VUSJ9yPoKm+xf4CR7t7QUciILgunjPwuc9FtQinXHLRtP4sgifZl4j/jgr
fAbebiDpR/tLL/crgYoQ6iuiZ3PDE8nbV7xQ+hmgtSu6zsA+x82+iMSpBtP8dckl
UcBXHdeaqOlFt3dNp9iWFHpZ3sLIxIjJIs/Ct0MMJAlpYvtt1GduEPlk8azZLBkD
e5wJx8L6sEyd4EnRnyyJIs+fUwYIbVEmR8y6NAgr94g/yG4xkcvmypA1zYkB2sTY
zrVmH3nJw3JxVetu2Lgsmwo/Du7ZKf7snIm5ozV2eiEUIwrTczF4Unxo5YQBzwcJ
kmZXrlhtNX1TrTHAbEnJtaAqCAguvDZeOxxy2C2suIE+AgH1c58bKNWwKls1I4hB
6hK5wMKkzyGHECtqNK/L3J5nLb4RKCLUJz6JWsH9TynP8n0ZFSfuxQa2PwpQctf9
39xCptEZ7LYq0is5dcQBpEqmbe8ug5NGFb4bIoL+FDL6E0nQl4umV2FJv1liNQ7+
S635CF6Nslf6WOg1X8ixlWbyiEoIFC/Ifvsf7melx6a7QuCCh7lW1VcirJQMAd8o
LXLEDRLCRU5PtMJvqtfV7vYJRxUfcpgHiZWmwZtyapOKqPvHimZyZOUdZoyNA3sh
lUG+K65Pq2x2CBMsecdPmPAgWsKJFjH5b7ah5WS72WFIjf9lW6zeCEgr7ZfR2+B1
lE6qreTXuIkrzegw1wrXPv6iSzj5y/fXqyVHeA8Uoa6TWlNuEqm04S2rx0RcGS0Z
9uA4VEcr2z0amPoGlEFdvW6UQt4n/AhVPA3Rf94hiiTdIBlAoZmzPZmo+HLC9kIO
LuBiDQ/omnOZXfl2xVojjNMVBJUEmjD0Tj7zxi+pVhIR8A3SFLIRULn2WqFcdzcN
jpfUmVjYTTw+TXc0EnZ6AH5iHTINVwZi53Bq2sYtpUw8HXZv/LNAlR5GaBMwgQev
lgcy/woE8cmm/9ny8suAiGApFBXMIDWL91nOBAw3aPxb8mYoHN/UZtcceacjWORI
NkIKKYBG3x2dwEHYmI7jj1DH1LyGilT6KfN3r36ntSDRH2DjLUoQA7CrT7ERZcCM
ipnOz3tYx04ppMg9XUDgG5oPJtosV1gzsnvU+n+khPGkLVJU+l5173CBmPaV6kMt
uUXEOmzlsF2K7i/QYch14byRatQYBFPN19Ndv5nQUVKwMOnlJH01VQ0RPKpBNPC+
tUwFg33nHbZlVJ6L56jN597TQOno86xcgXWbSoyKhmWyjE1Zdhtdt156dAor6PXH
4AMKIE5x1YA8nY8C3dgSYWtOtyuqOsqAdjAD7Jg2FerN5NUI9Je/rnQDRGNO17eV
3GVKpvZFo/2zyfplxn6k7ZFARYMKIzG04+am5q51vAsXpNh4XNnu6wIu8y5EIxkn
o0LjeaVWXqMWz8erMEc690QFSWZQATqxUxVhhh1z7ZAyIUX5wwWg1hcPS2UjGbaO
BjPsvefTaJC5C1t3c0QpoK0kjgj/c3v4ZbQNyMor0IsKVLSbwaIRgVhlNMKLJBAw
3qUeTmte1/2/AlUX/EbncAyJmY45Ej5WHnkGWY9tRx4V9kroTws9rZN9JOAO7fbj
n1SVok/gMWFKk8itr9n0w1wXHm/mRfemTRcBkWhJQRZS0tZaNeUE32pn1zh0EQw9
nMZpVrtsRghkOIwht4OoYIZUFIn8sE+lNfLmwTG4fLE3jwfW/h3iCEezgLesCfyy
0EDDDKBmSXgPRMwYUw9evMpuT6S0YlrDIE75vLLaJGw3+EVU1PrOaT1lUnXJRnj8
+6C1VCln7kuX+2FEQxMDje9paC2y/nYFWYErufyt+6udiXpbRhZE32Ud1HEA9tIg
EAWnLQUIMj1YMP2Z8tOlvHyuZuGAaROsquA116o6vPi3mckFWeOYz3DOEH4oJhH/
mHEkGhRATx7yQ+rYz1dNAk64voDVV1x2O3rNE1daKlMrdp4KMDptSIfSAl1u+fn3
RuvnPFybY4pJ4Igv1CZW26aTyjAqS9JJ+WV9aWoZEzlIEGfmtwyOn7mzx9xQ7NPM
omqCx+Qc1w6dlhLf0cEy2nJqqpmwKNj+tT7Mjw6UjYh2bxtymanIrRzeOXHVPj9I
S0RYrz5fL/zUAd7W3dZ07R7BD991NUj5ORzd5vOUKTW4q1h8s0KsllOmXY9ajJVm
sD7T70+9DWlFx8vjooY5ck43oJbIda0V3N6TsNjilXWXfDaCuj/DzJvNiGOB8oOw
0ny/P22YeYG8Wnc+Lv+Sieu2UzhdT+5ES7kTz8rf+gEcVppmOjU6SXDAM9GbOtcb
Fjvs8iK0yz0CMOxEPd8JJ8DaIMVQ8iYa3lzBA8nKbW+qhMw+ZUSUIWzVSPK7b+Ph
l4XsgnNjZU/5ENeQ34dyCV4ckVJ3StQVUgfGgAfFzOiiEE/mn6Fh5Leh3dg3nk7w
i414FqkPqE9jbEvTuXDZm91akGeGqCxQmvMYKYQzg/XkCOm20pvPpixONgQwH5vN
/P+OiGap/CmVuCFWAYiuX5o7C+p2MHlymVX5E8ziTotXKqmKNsoc4cHfPDHMQKcC
vc3PbKn0fWJRVEiN2lFVu0Q7GEcU9F4tcXrhJxpljTAhKOw5mxaL0Sjtcvy/E/Mu
Vdzwf+7EmX/vokQ8GTAH/JF2ANdnEEkL/c7PdGrS359GDOrkfVAHOf/TDlCkD/dM
ThFBB+BE87ZF4Kg/ply9N9vypok/ZgFrdoSPl3LYEH31OWwdtuBcHm+p9jHhe42l
CRR0QWFmjOCoQimj/DykTW1Vkkb6s1WRxZNjXRPr/gLSFDVT64O6fyBftMoqB8AA
kEWL+FlcVhP+/v5NzmSWsRf1/NlRltCrZsqYHE7IxPigG1hWWt1hvg3p6/ZqEtzs
1aqCNDnFuqV6UV7Geq1xQq3kcwVYGRS1Ys2GvHr9li9RXKfVFlxknqbaOFF74i6f
TNRpXCi2D7MuZ0IO89gO/58Hmmg0Bbk/A/awym0WTEgZdRErdrqpfv1FyzpGufLW
pptkQ3hrk/Si2whbNl6Du4xUxEQ4Xjh/OPYnrHoVXQgWa5sle+cvNmur9zU/RcfM
5Y9syVdYh47C2z017j3PISykX8OI1Ji+kvOEmlou5eklWw45k218/F8LWAa8pyLM
IJKVn2Jht4SFWEs6JIAboW1tyW5w4vt6GZbWuY6LIVc9TTIT4t6ZDQOH/wQT2WG9
OgkbvbPwVclwq1CbUBRJ6fygJ8mo6RiGQRJitcK6NQL4QnEkSnRrD23XZW8RkLDt
r24/c2S7Qkmddjp4zIItXgha6jWP6eEkZba/PRatA12Jt3RdGJh8yotH/nphKh8h
ULCyBMVdO1+ZF/SeVShzZtiQka+xuoxLR1wvUYvb3bm/KPNt0GIxYV3aPG+5cu5t
8llqHsxFbtPpLtBAlETppFkXdFzkyEII4jSz6OHJ8ROBDRM+RaTS8ha11gFEHPvJ
HZSlK8ew42vq3asaWYPrj4teAyPVyxVAhBCUNY2saZA0J+v7xvlGxu6fDjkbW2Tr
OzylbgPn05VPLLLUoWap1uO8yxhXxP2/cnGFB8UkirGL8wJNRirlqrUzVrl5CM5b
K6dhj7yeCoPCOF6As3tg6/RCXEKniSmoB0dYpVhGn0GZm1TnLX38SpclE4Ai3mOD
Ij/eU2OqSN/MyV4JPnVGuEsufGVgQSbwxawq5dmfhdslIkMYNqkwUG0m1Lx97xeW
12EWkd9cbvuNZ1/vIj1sLzeCRljkctGtX8lxfOit429r1i0gh7s76Hg0Vxk+fNVX
tDyD04pj23xQ4jcIxoJKmaS6IFjN/pc4Re66UqxPGDGzxh/8FE9WYNyPUSrhmbWD
lvGMuiHT/7vyhcpZebYiRY0z8hK+q6XknTBQGTjuyfV7QB1Vq5cRW5hqtrlttTXn
0qfV1Bbn3ZD9rMEALljSADwz9eNupXJXm9Eqs+KeRk82wwmIplw8iM7TBFYDnOaL
f/UUimy+X4AgCDM+99Q5Z3v7jXdG05KxYMrAFf1bAO/VcVtRH0IoaDXXe+a3ymxG
1/or9LPYVNDCY/zc4V2HHYydUP0JoS5rMyZlFjRWcci9sm991nMku8QlB9+YlWaW
pXkGZCT86cnl3UVGyAKwfkk2k2r34BWNNP4MSYDTcdPc464BnhXJa23FlXBr8FHk
EZyP+j4yDHZojGakg+CPtrfdvxy0G4Wjh6tQwPXCvFH9KeY3fkPkvJbOWTqV1veT
O2QXYBKtkSmEYW2S1Ws638J7Yok6ToJa5oJ/iNra/OBSQfj8nftXY6W1WATM7OHi
i+bvBESLf4AFf05lSvCyg3nj+Q8o+v2h1wED8OBBccUg0McHhxIVfbweNN2o0e0o
hWo+78ntuXb2sQZky6LHFVp/sZYFea96Unhu/YglpoSav9tjYev4FE9ve95MnLWR
VwmMeESjGZnTm08oN6pdN1AhOjNdJiHMC3SgbbDwNJaUmvRn5zaHu15odmIjB8vp
D6fc5VimiHHIhKMXtApPijan/j4/o1NvpEj9KmggeIhnYssxFXs+xkAV/eqb44xp
lMTFe2P8AgY8IS4UCAIndTaccyKyGRW5ymyyrPboy35bH5xVAhf3APGpYidOmuMI
y+09LLpfpyloQwYX9sHkKOCOVqF5qw2+c0l1xrvKGf6wa4CLO1gerEt93SjZRbWU
tOCaQ9WqIShDyYyQ4TEv5enEQlubawhpZw3dREV/VIZtz8cL8c38VZzHS90j7Bpo
72VgH6BQ42thbzvVNbgMN17zqv1VZeCT2xY9LHbRGpmXUnugx01yrkQHUFZiDnpE
HrM+fxKtrMQsnsw8nFi8R9ZT9jK29wYZXAuj7dJ2jBZ09shXmzkBpXIIjSLZRl3O
qa5ektBL0fCowCQXVZjWxTDXQTFJucTw+8XbHy+XIeW7tvwjTLwY7w0YEUVTRM3F
9LYTyndlAZFU8YT2hz7NyI41v3CwgrH3oo8ODDs8dO9YMKTEI7dSH84FBN4w8tCV
8y2XBkpA6yGM/kd94lzcFQ0nqJ6VYYGwKm9/4UJ2VHdxLb/fsTCq265luFlOS2mp
8vXy+Q95E+Iyfva4XM8gQUMKjrGKrYY88FXrhjLAaao8NuT3SFrgBm8I0ehVPENy
xAJcbik7Zl3nkTdkAZRq2ABhLIgC2RvRPEQjH2RjDtg7G629cpqIYWO7aOb93spR
TZJ7QlLktMNgzFKsx3x51C9zhLxWPlI6RbkdNJ48qbVqPxI1OqWj1I0G1vnkYMMC
3Y6xmm0xUt25TFon2M8E0/Rcfo2BYm3CBl1S1o2rOjyvCUV/YEUcwfx9a86STYKt
Q2dvjTEVOfaig2zFrVdJ3ir1meMxtMHEho0hm3mudJIjAvY3NfHnav0c3ptpPtUx
baHgqpzEOoZ5N8ea8iatXUKYlHK+A5KjPI3rc7vnu3Nz4iuzx5/yLYdmLV0j0jiP
ZNeR3v2GXTVAuQ/S8A5qpbooKJrqDCQ6yhZvp9WlLxLEzZiAhYrg0GslZ/EgVGG2
9sLGgiFkn694mk3sbCJDfb/GrsFPtjVA8dFk2nx2ZgYg9jJLRZ40RfgcP7A7oXfp
dEtceb32jigJt+olBmh9MfM9/V3nc0H5h9OTMAt+Wn1UgRlpzxF++HVDbI6aF7US
mwWBFKkKrIGHtt5X3JmW8x7mmcbqiUMKpgLoNvFXR9hR1j9e2fM91H6aiwPz4BCN
vDs0ezL8hgibeoup5zSL9nj0lvrbunRdWV81Ee0CD+FWU/vDJEnVbzgwSkBlMdiv
VNVu+acww1OJMWdexRsC38Qs4jflIU3sOyVqZbmDm0UE4Q4bAT19ZWtk26yHp6Jw
SYQ6E8q0cBxLOH2oC2eCBUPKHr3F6qLB/SCHX3aLoahvhZB053KSmCDY+v2ZbAIc
NjaOVlGk/3tWnve7D9/sQ2eUPKem/yGYdUlqNvplNIZIBZNRA4am4WE3oi0lgcfm
QAHjCnLXCRhLLNqjmbqw/bAEHJ4mSFcMuNQOWGT7zPL6p6eEbSKJcINLtTY6xpJt
IQCdBBGnBD6x2ckhrmrhy1ZOafgGM30s8rmF/w71rmOnhXc2gkMc8C1xGAgSmfyb
YN+SBZwKBCHDbC8MY3NgoTNAuDiABKeAWCl8C2NALrAfeDy3PXYr/pNKkE/kdOF0
VAxj/dh6hc5KdOkTe4NA+4u0eRcsjRcgzSQMyHiPFOuP6yESqSQTgzVIlip6Y5oU
/tv1h5xs858rzknSrw8Dnwpz3olC5kDcyhOB0RMb4d1lN/8kbbmPuVyCep70g/AX
e/8sMhC/XQOGlIv9ynUAf6Izm7dVe2POBJhVSvbZYM8JKkR96l+oQjnHrsP2K51t
aMgo4rZJuszlQgqQEdZKrnGGI/Q/2y06tVCE3kiQ8fEYVwrY45YVrMbzvVyALkR8
WAAqIq4+wQjb+kmVFPKNsslMswLd5vR5JbJ6bi5KvlDZhuMwZt4ZIebENltYswkt
7g34ZSk9SNGYx5/Sj0oyJdFMrdXRmMp84CFYqWiCZppqG20sfLXNm5vAi48dTV4R
a6a2wv0Xk6z9JcQSwr+UV3604Y1ZDwR6el/kcJIV1l+pDHhY9uQhkNgTeZhx5+24
sWktjBrf0HbynwvMM9nNHJ0FdKqd9ksu4k0Rf/x1av9upv0/yciVwHn1ddmH/bHM
3gXKW8gRmThGe1XzHp3Zl5GiKRYWlZWbV8rrl3QwEg/TS9SUtySSXn7wjSJReTLJ
a0+6owxxytfGw19lXAkT/hzvNMvVTTN6omDcAKAd3CYErl7GB9mI5fqlppXgMoqW
BcAtaYujBmrF6aHZwIYhIE/5sdFLTjPtTi5tAM6yIdzOiPteHgtqGzSDFSL/d0zl
pHpZosMwWXIbAkU/xINe4zU9hrER3qQ+zmgUzlwPKxyiMEHoo6oCFwUMDj8jGNAv
CxDwor7o4mel60riWTqyUgrJ5IP6NkWm2AsdLG4gjkIAvd/JynCdjHxqIh9fW3Ar
iT80kU5fD+AHmS1wOpG88NtQB1G0yfVeKeF32jycPSFMQLExTrY34xkifh/JlHj1
eqWXFxOHrxow3HS7tDjHTs7ZslT2yHxGcuFFF2A8iUH+d8S4csAqhyczuoD1lhqr
KhpFLkkoWDgWzMW53FwT15BrXqbFKiK5YDZP+pwbnxdv7NJr1I+7fxNjlVj5VoEO
PkOhPN3akOT+aih6W1rXQb9dTeLvpHjqnpjmoiOf/MoVGC0FDo6CFdktLUh5A7ZJ
ilbr5YUNeXlFfXpFAFnsUsDaXTcZWouZFZoEqpNcr0JsEWtxaOEquUjd+0ThQfCl
s6shsSxq7HJIhZmzc8FkGs6gevjAKZHkbHwFnPB0rmuVHF7P7/7q2Cv9+HH2j9Mv
aQwi9FWCd6AL+QHpAl3UNlBTc+zWLTdffNJHFfPY1MhDomuiq3ffkgIdzJbRA079
OcVgqi8vZI4YzElWDanYIxiPtPtnVRKklk2OiisaM+U8nr/L6my8X87vtN0S6njF
/xfZD9XRKewKtkiJOYN0dwubUp5w1W8nhKjdgkCM0DCneAQcc52bzUz4ggRQIrqk
CyxEqYVpRR0zILaNf9oc0Tr3F0OdCCZu541mxkZlRhknbYrfXJKMD4orRxYD1nZF
x6qxZEcuYXEVg2Uw8CYkqby/wnztWmahL53NbvID+mAZGQ4wapEcp3yL6C67FDCl
R+98Knt1GPSUkevb9ZdpFG+PKVOZXdmWfVviYb0P5hFOlXaINeLtqxfg1BX43rUj
wngpxCiRfqe4GvPF3ptlwWiUX3JfcwNvD3NX642ZfXc76CgRK+zfgLonUa769qRe
28QOqUsdHYIlThd0/HEIXbJNTuuN9ZGwEVCV5QKu3Zv2+bzDL0AN0V8PVxAwhaLG
CU7ey649TF6AXp+deZIZ8qtLSSxFUEpDGXFZ90cK9+VZMgaqr6Mo8qalxgvZHDK6
fDkmL+n9aueTNWdDNh3gay9WFnOSGO1paaFzSxZOxSs0YtlgwHTX3s8bB6EBiB4D
Lem+nqbXTfxbYmEM9XyWSoZWFKCYcUSyc2VQFt+rH4VnQBj/mGZ70FJcf5GWNqQX
AhQxR2kLPui00bRy7oc1OOJ2cEf2GNqFn0G5tJRWe2UdihOxb2riIpvNeXr4hfRo
ifFMmajBObjLY9Gz3XYGFklTTqOfGpO+FkVevHrdGHP2reO0RUzqgH9mfgdkUbW4
uWrykI5vaCYLACl3iRqX1/z8+TUHBLbERZ/DO7/SeOyXvkIKCItqIP6WLRC26B+Z
oerCBzH+CPdc8LA+7rofAPoDU0eP3OHN8CafYH0bEQ6VADYibkvDCpXwI2cUkOmr
B1+pTIzxNk/S6dgPt9K6+Pdeut+f4MR8lc73behCVsbSCwHjBQa9rdmz45arGgR5
aOLR6mxnkJcYcjKdgVD8pXulwpwzgHf0fV2Ixpj1qFIPJhVSMQd/vsF4M9FpdZ0P
54mEP5gCjycGeCzdF12A37QCiECkzYfOCJHtCaHT4mmYkEos4ByhjmsBo+wDT9L1
2xDYPU39U6/7EPPtVL3uzGzJhX5sjctAm28P80q+qrOrm5n3GZpkYToXHt0bsYwB
0WGxNDB+LrF6aj/HRQ167xiJyEF9THpBWlFwfvU6mCNDN/Q0/08UYR9Eqn1v9QkL
mqOqZBPH1ahYDuRWhLSlfMAsmmJrNe0NVWkmgr+j1IeR9GJ3ze1oGz3Iot+xI2/E
exWfmNyGhRyI9nBWOUGFQw6Xuf7XUTTHrAXWL5TbhouS12wUsH19O0R35NvXsdFs
M+PRlast4rnF46f9V8uJH5O8HcAxjYHS/orY0TxkMedmq7RLjxuIzYVGVo6lJpmK
VNwygoSK6amyKcqaqPr7y46VD7+4q5864qLLiVuFa/w5tnzlmTPx9gRgbpfWQDnY
ETtP/5ppWsc59AOKD9QCCv6JQO2zgB4t02T3TPatPuxkocgJJ+6Tr8E4U5R4FpST
Ps+e03xvt1Eu+jNFi6NZIa8+I9mJNqKWI0xAhBEm8gxJdY04fj9ed6t3lMOWRT2o
f9Sv4Gja5sLOPdFzUWn9g0TThcqCmwjcFM+Rzz08gKaQpHvhaMrypgvpbXHtPKC9
SO9KpGv9TR9DOad+Ne978LfzJ2uGzVxe1YdtKcthw0QvkKNrpjws1EFIhXo9Ts/O
tekeGwiHWMrpmCRTEls6U+GsM9mqEC+7OJgqNrIXKWjZdojhoYRCRLSBaPyDNUw7
WjLHrv6sx4a/a4K6kTa4wC77oimjTh+lVxrVBpO/+ZnBIsN+8czVVCARdwgFIJ+5
rzIAqz2bXno8UXrlpsNzRg/6vB2ZmwZj41YHJR+tKC8ai880RO4PMuTxWGiejeVa
m1zYok5k8+8n9RLzTB/tJ73Wj6swI5HwCGxCsMSPLveMnLH6LHBEe8xrRONtJHXU
/n3pkYPwVOL1megjJ9TiedU/sJWcVDVohdjlKWCJ11Fj+qWdT81lqPbGRCSxCSY/
XhsTDUhZjgvARPenW9r8/T+hlhpTe3MtwlDyPCJlMjx2mPdvZq9HeQtE/Aurcz8e
ts39/3pwyhbz2IbQf8d/UB63beij8PG28X+kxAnuFBh0qN+13uSrS+RaqhU9azZ4
seYI2Rg0D1gq25wG7+X8jSkkMqwCnFZTk2BwtjPoibLl7W8APLzZlpEgA65vv9qb
SamDtVX86ZvM28pdbgJEa0C0ZIXSh/31FzIp9IeQc7e7oExL8TBF4WJg6F/8bN4J
eY9YKSf/zpgAjU4gh5iWxYvEuBAjCSs23yvRGG2gYnKcSczPS6wQvT13NuGPOegc
xyogrOlD80IkUOKuXCVeIbgB4CmPbSFDGWMGmPUipTpxCVmnzMz6NpQOfBzu2z8m
57oPxbxAXp9FpqzNdFjvPUvc+LY46i9/CiMY87dpOIokmxIJYOr73DsyA1wnzXI2
5c+Rtac5hTMgV5sWyDnU/TRV/LaQRWne5SN532frjXxPw/Xeah8Hz9HaSCmlx0Qg
uN2glBaxNdHqGWUNwnMcK5S+MS1JJX1WpVQoYWMcxsGfzm/Bvz7JO0tOz3kEiHoN
wNKonlGomDtnYBWWVmoHhi/Zu+uRgizu09KQ38Q6ROiZZC3BEwbEbQvIeD87HwRF
reYwwOfNvaOndm9dMVfwxsG+EknolwmY4sNxbhEBItjYJ1710XDn4mn1GFlc/ukc
on/g4VNFHeC0Q9MlbzK0XyX5Hh6ZuXkdG/AFEucZ7mG4tQFe/tzTn3r/SQz+K20Q
oNmG1xCIHnrfb8npop28+j+wf7lrEC0oqNLPgkr+XBvZC8/DsKXI+qXwbeV6RLRm
1oiwAHFCfeKAk7dvE43WSLD8Xv6tXBi0LrGnqwYzZCdRpxpBz72pZ5erWPY8kDnb
KR0SeGnPi2I+7EY5ZS5pdm9hCqajixS6QvXSQMSKJuigAJ27LMqSIacBSNlR7KNh
PtL2aV008vKjRXJHEnUYgvAWGACZrNxb/L8Ok25G2oWYYNKXSVDpWHea+8PvrJ0f
RueW5xJE+4LSnMh8ddXZRULVNYNm6Qt24xKG4y5mtb9KpJ6Bxf+mbEHukXaqscmZ
4NhyPFqymfS1nyh2x8LJVD8f52n2NwGo3ZxtxwGu61O87tJR5jv35mJOI9av6ezv
hgZWlRlylVtkd58uF2vU8PQVoqvryPbxn7zIzsjCtYeQDCqMFLYVtSY4mNk9hQgM
wSyn69ey6EJ4BUN+5ArwMP9z3+qwXQqifJwn1UgRG3jTqTBVslkESzf9or0LoV8y
7A+D+4K6gzxrjLQVOBKiEQNxCozJor0rOVN1pfE1pdzvFMsfsnstm8xsrRgtWN++
648yrElHjIpUCbTuAoJ4Zw5COiqUU4p2CRqHtgl0HTOaRDB7J7iUI4RgTGBSbRBH
Ub/zaMwNJ7t44TH3n7nfGjHcsobSONuvPwuXZDGXTOOXoqGhD7s7+1ODEbYoV5d5
C5G5bUH4Mnbj4IU7wTWIgDk+r2CS4xFNbLEf/mC+pUjq1RTRaTeDqNyB9db4W26I
qluckzUIGuP6ZnlN5Uc37cE0mWgcqfkMWVf5iSNbKMF0d2+/vfWD5hanHRBNJ6bb
fHdOK2if43I+Hn/CdVzs6xr6RyafKgIJy5xabN3ptl10iKWbEzzJswg7UgIQ6krC
PzVhh4L4J0KXdKzJljwvgR6qZjPYg2sSiwZ9E2p5fieiswz/eV+pa/wrl8WIxbp0
q6Y+/eBYkkDgRSVoq8gCnVrzEuQcEWLlxbv5sb4ff2bSWj5U0n/xXCaarelifAeU
YievZD09+XaJ2zqn6jJgmJ9BCy6kJB2wwHpxx3GlzfT1z4cyvjKHVs2iU4GZxmSE
LBRY8vPzCvSgo9hDXwadDQrTRNiegRcMyaQdcp16/hJrqfmJrqlaIhnUun0dzYsr
CHqDD1uI03qZK8mOIY4EXkoQAYPXWmH5tA/xyQQi4DvfCsmmmJHkjotHN/+mO3Hc
V6WmERavwMcFZVf4Fi6r0DUZMLZjg5OooGC4UmDFDT3oX26Y2Or7hP/e57IRC34a
8J36R1Gs8ib04KbZB/x8UhYc7soWsM2DZH4FRvUtAsUrZ6qVWgUDrfrHlf4AXKJX
VeIWqUG60e4lhQG7u6Zl61GT1o2lxBq8QN9DGtsjX+q93mPfnbnzzkwEkVaYKOwq
f6DMFM3D9vJ/AanZAfzion9dg1B9FvCySX1oilwZPdtQvdiJZ0DGtICHCN8D+peE
a9jvLtdlxVZriNeH8VI/231OoWIx83RNYzGUe9fmYiZDOtwBFEI5G2JTT8A/OQjA
BgukKLCsos68XCCHuSWLLK0REdfri++AAKR4sEfCOkt3NpfGR1Zo/eYM73/KmVbD
RVgMv0vhVqngKU1xO6eQ1VvUOVSX78sgsPWRsRd8PI4kbcIvv+v0Ts04qHb18nI7
+PiTyf5V6YUweP2P5XF4YQmg6Rzz6K/KgPT5C+RQgShdmedBrrPnu24xcLczktDn
MwdeYcmkkGpX1a1UJB6W9kynva5F/m+19BdViNTGwGxeTeHKL+JN5SjB5QvFw8TD
CGdVxsdz1UPSSQVZmsFeNRnZmGL02F8m1CSS4gBmbuDNSGKm6zTnrg6XMCGt0eFL
PsXX0MCsVk/mResZIxSm+dDGzqRB8Z5tlIfUoz8L+BKaTmUr3CQcRuse18IPNHYe
LZY0iX0Wht5XvQDeyzx3wfNap+KOJz6Vs4pClET/fRLC7Qof/CbQH5xZr6lkGHP7
Df7KDAX+PvFH+yYcZ186APSfCLnMVCFATaSK62PkceHyo1ZpeKWHdwYM+uDvIRx9
ztBDx5wQqpCUd2XmetZ6x1npXd8Y6ZufcLoAjv6rStY2sJWEslXnjgVBhQ2d9mTA
cj9mhZnr56oIY5rgF1Li3lZMm5RYquXKFiQNxAOgtpZsBMxdvV64QUd3vob62Uyo
LZ2s3xIDW1FKZ/dwJMc1lmXUmJWmKMYNxEEt6J4J4xBvJA5vDSiuj1kJq9dBgWkv
+vanG6M/Z4BQO6hieQJP9REzM4u448nq0ix+F5iNCqR0d9WOmeaQNgHiVfZQlyYO
2n+iQ8bkj7g7q8072vwDRUPEwxOlNSiGvja2o5Z9dYXXyfGk9y8TsYqAq5fZBgG1
FxKjVbxu78fZmAvd7nm/jknFU1rJZPZNO/VB7hPcmac1rVwPXlcAM+HmLW2TWm7s
t09FyUpSdecMOhtBuhi3XSM+siBi8G6T9zLzdksjuY3Z8/k58YEm7f/4BhIdnlOV
2UESC1kRNzogM/kGUgrmYqV3X9gREBHPsd7131xrmLVd6YHgB3w/XfDkv5ckwrIM
0RMomsbmPawgg16RlJnltqYkpNO5qnW1kvv1uCZcNavnLOvJfKuQbmWINhMrG5yN
qZ3VV1TJt9/LKCdQMXoQusvPi9JDKt34eGeT4XkbOmbJUAqdtDGGtZpA2vI2kh19
7QBQavWgq5tethJRuZSWQXkTHw4LgWuT4YjA2TNcnK2LAnHhH0DkBd2F94sNbV5p
vi5XSxH+SE+8sbpHpuOoJCFaR8GG2f3u8bFHB5d1nkaI4fzWzgPakQ+JArWPa6j8
lF4+YFsF7ekjQkHPuC4AZu/KYqhfZycDyZwRaNYPWohX8/GQhVqL4PVHHtsnITZP
+L1QzG1hNDLVbPvuAjBxxhcpk4v657cVpzgRV/LikBHOPizYvXL1zTyrON7UP/X+
T/IFNcRn/jxZIlnXybF09xZZzSGtEQAByYYoEL4fRMZyl3HhZwT/C5bU3YsTIxs9
A3Vh7cmgSJLFyDYd21fpcLEPvIpbRLj/sbyBwutU5lTifIRZ2WY4ShZnP8clx9MZ
eDkK9cIChIy+H0o10yZqp1gVNt9en/eY39z7l3Dbc3np+GtCvn52oZlk44S9z91h
GJKi8U2k3ja0iMR2bVUyqmkZqpIRHFU61npM9Ma+lWrS9oHRJn0//KdjGluEWanA
kR2WsjfdvVG6VP4rBKXC/SAAhNNufqVGVHT3Dlsg/0dGeXCj+y7Ru3Q0zmeeBZqa
CGbGKiGjQmkjFESLRA3MU5ARMl5l+iynjT3DCMUmRqLSFO7OHBmW4lJdAscgctpq
k5yCNEDbsluSDLb+IFzMHgZc50UsgtivK8U2CXHE5mx2irjZVb5jS5yBaRTSS5s3
vdWozLC+ZqHM3gffRIGIOQexca+BxbR6rI/8hFLewgXcxd/khhdDc5tNyMbIExce
xjEX5lXuVl8IP2pK0RckoQv7ZXa5heQHJmb2LYI5DTwA1x40u+n6x9TzDgCns6uu
+HzKSR1hWiMkjFzaUImS9Sr9Rnh8POo6eKof9+dZiuPaSJk8yXsh0XI41cjpfUi/
XA8QjTD6HnMpCbsh2D2eoBZPhoRR+5w5U4bQBBWJtZjy8SRuz3m/u9XRJE4xOm48
gmM93d6WH5CD7fWlQy/18xxsgTiFYkZ7O1u5M2ZfLrg0oL6hzRMBZ5Ul8tdUc4bl
YTvCQAXUA+OZv/TO0VmB5I7rD4+asa9C1NRY3+WV/8DRyaXVPwGooyKxklfPDvOD
bY2vvcERMHfLN0do3Jj9MikaVKzkddLV1pJXcCXc3+HqKCo/+JgqvjK7RDNo4fvt
1aqwDw+HVmxZ1LMQGCxZ1Dl/0yoqMEHoNk+frsbX2K9iVgxZC5dhTh0jAq5q9oei
AdrpP0RhUJJdYznjVuRVlUkdRpKZ7UfqMpYH2OtJ4EGtnhiMAzd20IuTH3MGDEbi
6NH9Q05Hl+rIEynkZjHjiDlgEVPhdqhy5UmJvXD/rSrra4moArPf+v7SFWMY9AYc
wLrpDBIDVlzEnGbSNY8+23X4cE3WBIcfHdhqwlqeuEJDDYkG4h+g5kqBzJ8GSHx8
q2BKX0vjRteNIc8ehfKfUf4/gD1c+oESSnNMBvrHxntseL7E6txX2JE2Topnye+l
zQXWSmJcZFuaemq0LtTg4puHJP0T+xUa+/70U71EryRyb62+HYERrc4hg6qG8lGE
CrDGA/8On09xt3vR2tBSyo344Mijqm53kUWfZCh6CxQgQ3/+4ekeImYVoI1ylJcA
Yf5n/XEWlcuNaY7ryuGedLa+j6lYd6NYd2jHGvCL8V9tCQugO/iTcUHu5d6WerRf
m92B+hX9VKmjuQ1fyy3VzQVYPhBL+nkOoyBqoM8qvX7Kwc2Ck70Ul5gMXweimIcU
eAlFSOyhnp8DSCQF6NGsAQxWAmtpcOE+/bKkLg9eK5iw3J9EmfAcJuZ/bmjn8a+D
hXhoMQmcDfz1giQk/tKX41DXosXA+q4eiSUWIPhRQkCD/K0IJqs+PMU5Sae2TCYo
SBPTPnr88x2s7Cz05bCBDNTWRPgbX/ckl3wXXf0U5GtkdeMoxP1dNI1srgDL4s2G
RUs5Ga2+sRPfMZviAoj1w3qO4DzUn5gY2Vx6EhivHhc6kg65J+ZoM712F2miO4pr
AS7clxI003rGj383bp73cB7w75H/iDMQ1qD3rde9Y5hv7fQk+KxsADHMvupKBZzg
GVo6516cJrbDwU7nSf1RAg5jKAN1VP+GlsZNkR494HmlrngdNb7cMnMEpJiyqyrQ
EpP7c5YmSoYlT8UwY5KHsmDOU8kBhfUtAH6eGgABvwI0nRxJhyfPnehFOfgzlJHW
FSB8xJyPn1a898A1art81wXN0Pn83HX7Skc77l3JlBayfV/1KrtHQvimBL+i0SOF
SWE9omn0L+d4LihQ9kon5R0da3HlYgdgyUYlw5lyFHfomH+plHSK+FCqSMeyEArQ
7R+3Nv3vG+DR8xZM0JImZ2GsuWWo9mV2pbU7TE6oR0GotSOOO17V0fXCkA68NiXb
/Ah6kLj2+z+yYtdRrlG/qx1b08io2E8Iter1aB2iHICDTr0aWQ7QeHD0bqNlvima
NOWlA3Qyam+XcMU+41xUmefWwVqMP7gNxSW4/4h3DFdS+0arKpx4evR9TQy2uHgP
hdYQiNrQzOibs7F+Rd8FpO6iF3eUu3yTPFy4g/9iu8CCTLZFsXP2veinQ3uYzCFZ
vafrWg3xiXNLuhdiC+y1bOCMgq202kH6oWvDpX6CWVUsxsVOl9JDTm/IgbU/OcT0
2jfec8PxO5IUBe1t+YUSyzRHd9/KrShNXLXXO8zoTmn+max9uqkXrGPcIoq0X4zi
OE6ZoRH6rKs5YhMszXYh0OH9Q/fBIzsxogaF7CRUpn/dRY0PRGtGdgfPxz32oSVL
yRcDfRPz12qR6CFVTmtpYQiZPmJofJOvX/iJaZDCKt67cMD/gUfpbg/pYmXwcXgG
YsXQvewc/f9VlDm/RFhe/OPstxRMfT3S0NN2+Ho+oUyQHOto2eEiA/2Il70hUvXF
Sp3QXPQ9GMqESCdKVV5wMnr7KW3pu0E+r809bHifFmwn6usXO+oJp7kMnXcW02HM
tCGqayLo66Acc0g2Oia9QMfU7AzWkbFLqrEYm2UpVtVn72uvii8NljtThzgWmmu9
2osm3E6jH0aoTwF+/MwvwW6PNsiiCzPoOAop0gWsBrfvm8axaOq3889cZ9Susxzz
489SCcQcEnWp/W7bJ6XaBOp7C1ZzAXfLZ1YDdsqiwJoN0HJdCA3pCrS/j8Zyb4R7
B9VE811zJ9pvgnrVbCGgPGnsixJgpWQi+tpEMBSTlEzG1FQnqgqxym+hF7RiwlDm
kYKwAzRrhhgC9GS5pVCLx46aFjgDLiPVQPlkwrA6mO1S2p+cuLYIfxS42VD2Iha1
aFmH9pHUglJ/rkaczWSjnN4EnKj0FOEud0YptG8XSQnZkt8KxlpLecAv8deLFGLN
0J8S4B6DwmJYqFXOayZUgzLAoUEPkUt5z0OzbNYFp2WCOGAfYoiccIUPAmX3Sv3X
dTwIBjGo78eXfvPgVvunx7d6ACDVOpOfMoHP2CKNc/PmycNFvnAzOYatdsTg0Js8
LFqbYA3HwcuL+dSfrqpKp5O1TRZvxbxakjDMk/RBMzpG5j+Fh3yCFVCbuwKMg9l1
WQeQy5JudmzA9OdoH81fIoRG+KJeQaQEAHh8NBdLvJ8HSZ7xfgxtO+CuLeuCmsnV
HPKmUvHouxQCiedFm0RjsVAtq/uITLKytsZvJedqaAZmRgDHN+EpP8m1KhKAhZD+
1+ME9x5c9W2Cr2ypQuozH6fsfzU6ikv4BKUo5wFKn5/KejRCBZns2cu6TOMSkc5b
PPCL9tbLLNvD+WB3ulL0LTj4+5zZ38I+FJY56cZr5R93cY7h08wXwyPQClAQ761g
YyCJCktj1JlZlXEwJMHSPrc655S6+yI63NgAoFrZ0bgohtq/51N2fCyRddYIN8HJ
S1esW3EepjgIXC2Vu3D8Om+sgOjXKIT/FFJwJxbQZmWOviFcA/oQEjupCtEXd4hP
AYDRQjEIjsRIL2V1mnpYlrbSGW5vB+mPPp8swuDr9k/v/Pgp8Hx/Y8GanaTyH86L
KCDbghJo7xM6/9ih4wMzrU6H0/NgNR6uR9yV9fL9c273KJpJOef/Fsd3jGiVjwK6
4/10EjR4ITjwh4mEkpPXEvCRy749gBn/B4cKYqi8ADvDftFkzn7+TWu5b4GrvSGr
znd86ixlO9zrSzxx1PSgsupL3/P3s4/TJoB+4C8cnSTzdCR/ALCfwo+H/jr5ZJjD
gesk+Epobzlxb+L0qtzkYl3R5G40wOxp/Fbz1xMfm6yhU9mw1V58OrVxsfl7d6fU
of0CE59Fo8Q4d5Ub0tI26Q/2FX03htvB8athPTKeAXZasuwRrf2YkYqPrT/jswqE
puqB9iSmuC8ngUQ1EDHDaF/u2WNceFy7eGqqzJVM5X5oyYiozeCJMfYp2MyHO9jz
rtJSNP9ZYiN0kqRwAAxWe+pc97dLnP3zkkcUoy+iZUOS1SJbPLFOlqJkUknrjXjd
wgdQ5ddxWft8AAOvbZoSEfNrsj6ak6Nk6SF/BQu4aFWK/vMZSTSKDSxuq8ej6HaP
PVR/s6BRsbD2o2/qmjzmXu3XyS/heoTV4s7Xs69/Kdded4Uzl7kwB8d/apxUUzDu
vnA3r+jy+yKdcKqfglA+q+k9YdYbD7iEFdFDmjRmf1SwO/8+Z6YCMVLGb3sDUQw0
IFYVsXLmUIav7qpcU1VySr9l269svViFZ9R3VaNOpFYV2xaCEhF9VtRJ3O+fQCsn
Yn60iVWf1xxhMH6VjpKAXz+tloz16xVRNOLjJ6anVJAxFS+BM4sYJFBCjiVME/97
T7vibXIu641LPEplBtvk8NedCCVqn6rN0T3MRLqqx7lpaLTwEL4Dyg//KEyVTAs2
/vItsp3rV4OVCPaSS/d/RZbbFjsy2Hx5zYt8zn6t/02//o7UMvHtggTc7l1qg1z5
Zp9mMObn8qeKCZslt6A0X1kDG1sBIr1phqgLDT5Vw07WHKJjnBoTAzCot6ije7pe
zOkfq0WqJcb3+n8hJrKpU/2ap98BWvm7fVakea8ekXTENBP8D630JYyQwMd78+u/
4f67sooK7uLERzf7jABOb/OitBX6JOwMLWsxmb8chqb1MtAhvjxRQLGOy7yxYdtE
fUCQqTsKrGDIhXFtsZvxRrH4YhF3FC8ugIXvD6ceoF43qQqWCfC/iHPbJKqv5pet
UjY+iWpMv+QZythZ0j2xXnn0np+c3bNDkWmKoB46qMvxmG+rxwEW4jTVoTS82wLr
MFxH3jIJVLZrHoc+/KQ8bhUHH/GTvra/tL6GgZWt4okwmWzmsq47nkCxzifbdjkg
GZAQa7WUOL1SvD2inmBZrZZKYIrxfJbM+XbW0n+3LvVRE3EbvpNWsw/DDwcUPPGr
dqlOCjIneq+/4rKXzwU19IkkGWGv9o809KyKeBcBkFnu78V5JOGJz5IQfciCv8rw
jQ77RKVfz3CFbFcYWTinO8wx3CSQKe2mcWQ2patfNJoesD/xqjLIub6YY6j8tBQN
0F1de9FKbkTRpRA3qSfku1uklZNsxA4ZsgaX/o+cJq7WBRlhQjPKYWMn+msTr4r6
neLhZQwWEg35ziCl+DcMwrpnl49BQKxxN1En+EXApgok2D+h8Sj+3XzFFqdIX3S2
/FERzP1hZm06CH0NNRB4fWnE7bJUzuxaa2iNJM454/qt9PUojzY/Gq67HicccVXJ
uK7rDMUksSmFFZKybOEhGllO+MwMNzJiQbeOCUKbYvnyhoIB9yxWpU+IRoq+sIL+
xxpVpP6VuPe70klIVSMplLjWWqsN8HsZ8mWutlR+omk2KoGKSLDArz7wh7SFiq5T
kmV1IQv2QZ9rSJHvOF0KNtJBwQ1sPmEEVb7U6NCijUGfVd1h8lkHQ8zOQvRyB2K7
o9et8LkHenZTwXqfgDEotdA6FcDN6AW/33TwJyY9a4e4P9SAdhbYgIB7LZ88Y4IT
4QhBcwUMISpLgufbCMBWdeCJG3VQklN1JUxNUe/+SwcM+q0/fr4M0OJoeyODpfwt
KEGnvnUKmHg4JxkG4ARfu0jhk9s4JfEtl816uECwipt5136it4Zl57re9ZUUCIpK
L4JvyIHNsPH6XhTPOhxgikOZwxzxxdNJgOwZMgrrYDixZQ5JyKHBb6Msmp5oJrl4
3ku75yPjJ4iHUUDI2A/PPkQgSu2OpnzjVje4pgLeBjNYhTk62EQFAHVwZ93pB8x8
nu+T4FSAzTMW54OZOB8gBEPOXCLDfYtNi2UGbxf6pQjjoK7tAW4XM4PRb7aGyjmS
YQT4ebZ7r+3w8228cEy4TobfZk3NZOpZSfeLgi0KpGaffqOGQSaKoH3/1MslBXI+
OZn1UUlhJcK6kqKJHg8IjHH6B5em6UFvsy6LiEAuxuxJLbv7eN4yg85i55CCILdx
WF7bljjrwvrLJBAW4hNKhf9am9SR8vKN09ONNomuVz9oaYpHw8S4wqO3hz4IN+ll
+VSRpR8FQacJTJ2cox1wRtWf4rVKYps1R2rcwb89GwcAjB8DZYZmqpR0rJ4zSW34
0uIVPzpdvywAuXhKdjl2cCHgrxrRBDD9sgP3PTyCLLlx7cqVT8b9HwetLYdbSsjM
l8t51lFL+fAKuhR3Mkyuq816nNM9Q93ZtkRlU5Q6ciAQ/oU0TvvGcXDFUMOW+wAA
Zt5CoVton0eTbXAVOnqiJ+Sfs41Tliaxp5x/7ajBQQokRa9l5Rpai1gN9NI+xa+w
qnnYH3yUgMdtk8jvGkPpLM7fhUquQYczX6VV6HNtJclSCdH7RZUyFX6r5l1WSO7J
VhMaXmsyw02bttYrsX2DoUUkuR0/2cnsF1ftthM7k0zpaxqed9VK9wUHNzjpdcQT
MC8iCEeoj/Rfhg2PlMhmHneLVWK8QgZZEGJ1KLZoXFtfiT7bitJ7IbGPY5VQ2jFi
ADsdpacYMbKIqaV4oiwmvvFn9wVS4WscLHTOREBQpVsjRP2cL255ys6ttXC3PXEv
HhhdAe5VEPvGJCzCW3RiwhyO63hd2FWzm3FpkNf/NHRTCP5KVkSNavottACs+N/e
emIJ4uT1FMjToi/uf3R85Y2RkVs10GMS4TvN8eags0g3ZN33b1N8p06i/HW3Fpy6
Rmfco9Rvo3R09qY6b+R3WpWoyJYINDQcDIiH4k3391wqigiU4TG/6hyiUFo7l96I
TY/U4Yo1tHGmwYEyh8WPBxie4AMRWxaGfpkmLMs0l/kfny16UMxCw5YDrZS0CBA9
B+7nQMs3KFD4T04w4xRrPZeKEufd26lj0Eli+8uxvjVj3Fc6G3ZIEXHdQPAWIsf1
9j3O2uuXuy/1xW3z/XiKdwukrre2jNUJir/6XHvw3aUi8iP8113VnFtDR32OLKgb
QgepuwqDlHkwLx+ycNFJ2T2y4wwaFVGjNg/NSRjPBqVsGJKbwZ3p2R4dQq1KDTGv
I3+k2VkzKOCHIt64JaM+bzBxnIJO+4A5vD/tg+YMxjfrNA+nvAxFeN1KS1Xw/0KY
+w85En+1NAMQNhVn0uGQNpm0MYLDYqSbN/gElxLUXYMPZtkE49s8y3/GhByU0zq7
mpXD3/ulb+K3ql3UbcifQBkGrYrxGVEbgb0oqPpk24SmXOE65zv1OuQGwIoq/vbD
D1dmInxRrmRWHGUWWBMH/7t0ATCjZwOm3FT4j6WR8tYejPUxm51Tb98ja7dfcRat
uxhW1wx1xWNZvL2NpxicXiu19SsFhlhigqvq+W0h4bFhuC0KTBULx9biSBG15bcw
+/0DIFOrX61fq1Qt8edtpiVvA6X0MB3p12N17uCTBKk3PBwm273t3CNZZ6QN1Ogr
e6wZbW4xNDk8uA4wBBLiWqCDrSTea3zGSV7RcECwARmwtAgA55P2emhXUPb/EYGN
R37c6KVjNdAlNO5l2VF0GzmlT6u3MrBF5bOONdSuea4OKOQwFqpWS1J6XihsHqV6
PvJDDvhfPlDl/kF42CqA3EX3N7ZcOFaCRyv03ghSb1iaST/OizWvTwyBoLFXnJ85
EJTLnt8dT3K040kyTPAlJ4hw+2f6jyfr8ZVQCtRKvkxEYNCR+v6hGJkd/FFMgeHU
KQCRKGL684sN8xwqNHq3fwObES/A5PMJQu7nuIegO0JU97ap8NxolwUqrT0pb++J
9SPAHZTPw9g9Q/qLbls7auRQvpJnBE1Sm20BbWD5kCcVcX3WG6PUl4GogqjKKcvd
Jtft/55RUFkvHRsWj0DjW7U7hUA4mVgTLZEMewG3DYtsb2eUhMH0ccLN0mtmbNG7
hb2MydMg5ZxrKJCvgOBlaw/bFxvAN7us10VMKGQ22yP3WkiwbjAX4qKUvOuQhOdJ
FCqcsWyG1mrDDrAHFdKV+Smocfog47htfmFDMu7SNyHVPOxxArw6JEsvYGJHmmJI
nyhTj4d5+x9StDJCSHHNbwDyLyO5icaL6JbLFoN8i2jGgIMXHw3Ve9pG7CK6NP15
RgDNcBPlXpxo4EHJR3OzsqMYuvsCQdmjOygG2y8CuSMXvy7yVYtCXsbucHSQTCi1
xxBIDnhH1eLQ2Vsn3SytpkGCCXq/uXjs+Cqexs35sfHqK8M8bI15Bsp3Rps0llgt
J+wFJXbbHn/HHsaEEdDw8DU6kW6kT2es0+ioAPaRx+6A4azcVnbxrSDvnhyS8WQT
y1KqaHLjOcMtt4HncTIxYGhEyYF2H+NAcDuSMmlwpuwyos3forkXqV/OYByrM0l/
e0LyU8KQOdT4C0F386NTw2PmQcmWhdFlqjFWfBj/4v6J1k5/a+wdFNnWtW/42acm
35T72dPZKqL82ff4lvq+mJUnBOE3vp5rgLMmSXYwG9V1yFygCNEdmqPFM6eptmAd
zAc+vQbWC4i69MUn8m3cVX1Me7/gUHcWTaR2TX/0JQh/7rf9OD4pU8oKEntTiipY
LHAp0H8Ybd9UKp3Rtc+w8aslky/6wmCLwXSxoVDx/s6Kyz7pzrsdJq7Z12TEUMSa
WfaJI+gDrO2xkpGa10N/KCOM7jXLzqXb6sBqegT6dVn6jjNotDS8FBa7itW6sjNo
igmoSIUiXlb1xCQ0WR+adbuaeSn1QvCDoVyR9UPAaAycmBIAN/1k+N5Wp3yfAoYc
EvNokSbCkBwySudB6Nul853Za2CQQpqeItanXFdpSx6u3wgONZmxI013DzwhH+BX
kRu1AGmbJreawTPGM4G3TZGOHKNSx9MGPL1uV6FEflowYyDTDA1PRc7NTecOaZhF
9dykfHH2g8CmmaERbL8t7ANdWef94u3IAlXpmioARdmD57NTd4igxctpsOK/zssn
hNJt22Y6s6vjZ2n31tuVURPmf+TNjfHYFfx3PVx1UGMNpHNsRpLjIWcmSRYiPxkK
sK4DhXkLM2bdgxQFYCSRHuLqNYii5jIqMi2f6S7Kq9zi843/zTXcRlgUs2jCO79C
ziNx/bjpbfMELW/EueqFKhdLYWbavkx1KiIwZpjSe7sRbOOZE8hs5NWztQ0u10EX
X6AwgxKyubHAhzeU381opR7Hm6hkmBubJx/c9AtIdZHoegcskZ8rYIc4pFaKce1G
cOq2PZr/otl1jQAgK+ETq6SNUb8Gboz5gIF30dZEr1j8KbXQTQmCoWYuEv0OKx0Y
4/OQh9iJ0+J+Ztdd3mp21SLdhFNEPdqNfPbNK8ia92gjLZ/l/XQ1cZbLCyiAHmLF
Mc3bkDSmD8RoShd4L9sudtW66UNmfKVoaoWHE3R8hRWqdpVfhaTeENFEKPwdmLD3
xx5FjYfmZ4loi0dWIghayqKQbAItDNh2j0MBeo5q2qsqsymVWunsdVvmW56Wxpp6
XNZuLqyuBVmA14+kJnnXeGlxZ0r1dJaB71xdgZdMG5o4PkWoNLnQWxDNudIHA5bp
GZ3oJZA25KvLoHBTUZZ07PDauTm3W1UwHh2QYPiOQExv7yUJvYiRun210EM+G6AH
cp3PVSg7dvvdj8c/UDVfY3lrL/cuSlh7AQeP5py4YsxH2DmHrpuG8zrg/fedNhJq
8+QdFWfU++bWRRdppVrOFdv3R8g1IZy6muVl9LrW8ZKx1SMI1YzN9XR9JD5ietYX
Wv89zHXHK5+LmauAb1Tu4S3BkiyrY4PjmdEI2mGIx7qp6yV2t3efHSa6ldSR5n9X
yhAqHmXHXE689k0EMr5mHCsPjgyke68g2T83yN4h9ix9eKez6Bf2jrzAO+3IV6Gr
zlLOqImjRkMZvuCGt3iG1PnRe6k0JXJ6uiemNTuMfOV5lyxq9eNlI4Bd6dH3Z+bX
5X1p3ZfUVt3zGU/YcNT0xaEGEgsxcg8RGxAS1Hi0wXjESox+d+8f7oFyFNNa8L+A
KmcRqmiI0rxEL8Iy2Aj829SWqWSMOVU4RRY/WMlHxp239Yb/+wF+/YxUoHv3aOYX
EqYirAjf5G1F7BF+5nSWN5DVVVRdZJGcHms8RhMpesFClaOin3g1tR9ZuNo9r9r8
sOtE4f8Mg2HHSfiUl5vrRd9Aj6XkMYAoKpmn/mYaSBj8ssAWF+/AJEAe88bBA2LN
t6GfFzG9aNF9FtZe4VFXgae674gal0EErHx8aco0I+cCC3s9tYqI5I9x8vGj7jX2
Kl4q2w2EcrprAKp/wehg3KoMIdSlP2SBsE+ro2Gf7cLC013T8dj8Cnmy3qjxGKFC
fnZvxD7qZjBWfy/OeXXK9NuHPco5Uni1KxNAw1DdMK5+evhtRitc4tUmgnquiQJG
SMzgb3bpHVLc4bsC0mkDdDagMHvLVfbdKfXxy3LYYl1euYDOeY0aRkIZETsGdS+h
ydZXmSG3lYvLpAoBD6Lwl65oLmbA6HdBiHm4K0Mq7UJ9T2suNgl4WfNxNdW6b2iZ
0+isVFCDIhpFY4U56mXbxxO5yKS1GhS/Vdb5aDAw9y8ydyQpBMuOa25bWwYNLa/v
qwI5dO7pDE8BwmEq2N5XmGRvPmvJei5YMNeOJqCsNwE1aFCQ/9b+2hAf2v4id36f
2EWXRw5MatJNDF1ZLCLhiRogv0SaZpPcuWDEBlt8rtLrvJeMKKi0tcBY142RMsqD
A20zKC0uMrZCjatNVF1v06hgXwg5Fo1W3NJ1PeOc10l+Th+KAN2e5QvLDSiPaxJT
0xNWzd12rjOHYB+e5pkyoka1xg1H+DXYQ3VR5iDS1gGG6M1lC/uCFCel6VNLilm8
LloJ26s0chGGPpdWh7Ud/UHXqI7RclMOqCn/Zk5UTQoa/DlOBljmaklPilnxyRtu
7SQHnApd/IdRlVBsWLfr9pp0AtkMwqWvGQLUBGjPVd49XsADvk783fB0nB6jb4EX
Hh8iRgaw9Gvha7+1KySJkwzUn+K6oWvexdt4LAoRdQkw4NVEl6XSE88jgpl5IBJB
xpxpdWa7j9k0BMs6RW6Z1W1Smy75UZq1mggksEjJ2dH09vvRBK34cG8RuWG3ICXU
FC1DWlVBhllWwv3FsHpgLqEXU0BVtsyZ4L5sLXApFIMzEM0xX58MA/2x7h1+cE4k
OtQfhgteVzBgnhoKXw511p9Mj3X0Ymfy2L67Z2labxR298AhQMlkOV8c1wkgm8qi
n36fs+IEpJs0VqgkuVSgIyixV0rnY6fk/G8XpqDGzjMne1Jl54kzlb4RScyZQrR+
FC/dweb/+Azt1VZgNMPiPTE6uGboB+V06lpuSOKhYAqIqqYhXaB/GvtAQzJIbNWM
EjqasaGX/H82JkbcgtBAXUCkFJ+nmurYzyQZ9k1nTv4Xa1RlChtwbCNivsQnT6vW
1kFKTEKPgMngrSNCTgBPTcYzEmvHIi3tTzjCbqD5rinmKiAk4wMb/AimuZiafLnz
5dqaFb7jkdK9yI8cmRvWj0U2/o4QZZ+ei5wSf7N1dzakfS8QmNLLM7P+azlbhaXo
aDqxjnIuB7+1pnVjyewA+eC0abrANbGRxkKiseh9PaI97O5WhQMXLbgHNsgL7JQU
mrv1GsqBOZKUeW1O9HPswbcDwrb/Llfa8nlGVYElNXHs1aXiOupcXEFBcPhJ4Q+f
3zc3h7Tft/oaVt3to4iqG0+Hsh6eoCyXtjDQN4o7jRiBC2GpKHDoYB2YdFmmL55a
rSu6zkJ7M+D0LAUyASCL6m3cjK2/30vBrdfZSM0kiVEDy0XNvSzqqNtbHtU+V5H9
erWx5HZmXt0vOifpsj4fwwi9KhX7Efe4Y5OpOrkBIenYXtM34vAm1iLwiF8p+8aa
3RBJ93zsi8clsfOGM5qC8vpBNuTpOhMHupbaFyHFIima2V4+I7h5ds0NqdeY0yes
bKnFfM3sORdjrZpTyA1q7humjLbXYCL8ff0FxAZ6YAwzQTPKfHgeNtva4qD0XCLY
tncNtUdvNrtU8CrI+BbzeoQxY5LU2ejkcwA5NXX7c9JVm9/QlidcEklbdExqPYrO
KiZl6RNOXs7AK7Cm2NXrmW1aaMAqAo7JJSoUHZ/YIKV4x0D8LMK1K7rAnFVt4IlE
HSEClDHK/nBEl7DORuAwN7sjFB7dU3H/NaPsBUL/7EzOlW4nfNdLZGARtotaWeAf
grS1MmKbAYctl8Zbk/C/b39jjx+dj2pqpMA6AW1/wOM63jG1Y8Uw5vsxlCcxOaPX
NOCmy1MNL2EkgYKZiqNJMhRtk3EiHl6Q8PRYqjaie8Ol9rSEdrkraTk3KxnjG4/s
kAcU5tZ3i7ZQ8Kf3Nu8grqHsSk8QW4vj6px8a+79em1jFwZY5G09+CUWmqtbhtIL
xJdx0KPAPyncdinCsKjMuxf1zqjEaluQF837OzN67bqaFeSKYDt40Pv4iSe2h0Lq
fajIB7BLC09utZ7fnIl5IMKVoM+G2A1AO3JbhqytZCrmQL9aBQ1KUSPXBpssC1QR
0Vj+Qv/mHNxidnf4o3keKHxie6fvtZBzkv4h4i9HR1gnZWC+cO3UJzo5I9MY4VEn
xLG1jxtfQuDl5m6AiSem2VAc8zULwQD2/ayalLf19b8gS1MNgFygbuKiEKHjpn4R
lezl6HcePL+xCHfd7loTLvrDWi0SsjWTtn/WlYHXKzZhvo8kqaODr3YO67aTybZQ
tvWVuzD85nfd1OZmhbTl6K/FmV5F3LBsLOuncpQsbeuoObE1p+/K1VTO+F/3+ka+
bnMOIiYu0dRXdbV6NMGXLt2C/IS+LS9eoRKcoVvB0gynHbPXxLoH4ZC6b5YliHG0
DiTCCQuPAwDxnkZu2p1s0ThNwc9NLgAKBHeoHw4LiRey/EILd1GS9+R3RtZSXLhD
rXParDQcVBeXVl4PezSKrhtEt4pa5e+SlOABJ7/u5LrO9NnfHZrNtb588l00QDwB
Pbq1TM9yFR0sxh3x3aucO01hMkGs4j542vcvWH4YAryB1ThWAFPkPJ+t85OtRqHT
g05TLMTJen1tJB06psKIdww2olla4qeg/l3OT57qF8nLA/yu7OiIyk2AbtOUaa6o
AyB7xJvY/oaYy+3L0jvbhch9n78WZy06kulUVfduR6WacOhYOTq2i9RsVq9lKvlO
szUQsxBcCUB00PhNOEwDOXjVbyG6FBIJsZX5wP0YW2l2QFeuCM4we/CRRBoLRBLe
x7iPyOigjjDQLJxYNucFQeRlmnWXCdExksS2a+xL/nDJ3+VlrHKG71tRWo97QP23
wGJgIjekXuFXSE6qnvB+opltaattGENN39M6QhV1ZDqNet0azpDNV2mwCfVvOEBs
FE47vzLnnx1O74wLHhjfzOZIA2nGXhPLTSCu5wmJqOlkoSUY7JehAqXC4qmkOECc
lgEkGKtXLHQBRZO9CmFcDaO4vNBE9OwRDyzDkhNRqxDwyHJc+ROnfTeE1Vsj8bnV
gzOfr08hVRIy2gSJqplLBdUJSUMf97E7+uBT2bKBSG6QAE+sPDwKHbpBRRgTa+gU
9nyruUoaktjC3fKRQR4qm4oSChPSDTTvyUl2ZD4UtwUZtv27XGa8oXMR3G+yG2Kp
V4ulpNA1dqGjEbQytvVOjZQvKCKvf04OxuuANEE3paA27OWsPEeenZE1aat2X9eP
YFXSFwCUOHAnTbqBqFHQIsEZhmX8fo14tlLsI5nQq7W1ybI+GKWuVmhqKOTRLClb
jGKg558bEj1EHAvuGQbj4eE2SS8Tex/tC+AdllHvJi4YqG9J3AY+4lTvduKai6ae
ua2KEsq0thE12joJhu+er+GW9C4GQgoOx2p58W2DZrxO3PEgGrTp+mMQ1U9Lqsy6
lGPrvRKKzki+ipw6zrRGiWoVU3ARxwmu9F6gHSJiupu118nC+KrAD9A1LfE2f+Hz
ZsP4VbKy/kjKT6l85FJnLcgXIf/t/3R1L2lcxxg5xFiM6vZQ8YfWv9z3zeE0GL7I
xw9K5H2XBsEiC3eKpxrkNG69Jr11KOGbpo793/eTI2Qmswm9ViixlfMGX+WfZ6Kd
RQlz0m8PGBq5cTObvGyqBkqIdOmG6PK9nMIURUJKaiP0+33/lbszhk7NkLSajpg9
GEAkCOSK1TSwnnKNQRJkjWeKWzaqdUjDkuCvJ9DjFu9BhvyT32N6LIA8UMhBGQAd
LGVgFdU93ODNxYmowG1zHPTFsTD2KeC1sdBoHAdADSViJT4O+lDhAx8P+fyZ9wEY
qxDkgddVC19An04Oj/6B4+2bytc3u9jtt1cklTIriOI/oCVD2s+aNqIWlXZv1vFx
dR2w/5Bo86EfCWm8UgOXXx0M5zRmpg9iLpO7kV49BKjswOQtfzhKG2HanuDg9MBl
KFWgiuX7flkZZsBGmri8YZA90kqnJAI9aiVc4xHKwj2yczov7Sd06QN3jM6CUm3w
kI3lEsD24gRjIdVa5JpNhQSbfwfkrgtFEHryjjZXfF4+PKcMjijFAAUzo9d/1T4u
z+S759dem/o2pxfb9l/7QXBT2sSi/+5FDTmdgYihE5tkrTMKK84QiFqQNL6uN4Sb
QfSGCQw0Mz3LYzVhhaRkHHg6LYnx/YTYw8W3D8+Qy+Nd/XRsNdOqcKnFSE+SzlQi
lSShwqGs+akhSPRQFiPQ0NxK8W8sWVc/UQp/KStOEilRPOnvMh3xRI/B7yIpaQ2L
ohGw/jyPEgCVbgUFTsoA2m9uEQTKLUJdeHz09/0tyl56bJ57EU6m4IT9FjmdUQSc
/JebLsIxpkTpS7UnpsR5/jPvrzG2JuBVTYC5cVtYHTqpuylzhk2jzG8Ug1aS1yrk
VTHNRTcU/ojsGfQSLBS6PJNmQSdZjdLwxSU4RlCv27f/UI5pSCit+NLSfNq7IEQm
XmaTDQUJ6gxOA18jg2nz5JAex7c2nYKnS+qp/Tgmvv9wq1rcbUbS2gqQcLPc4SwQ
yeh3YjtsoqW4OMB//l3wpOj54dcZ7RLD8LITkn0S92M8IjMbMsCBKuq9ZI7o5l3b
KzYPy2jgOQOPaiffDB5zhFQmvZOmrk/3LWihnD8tPH2BXA+EB3UV43zr4hLDxYrq
yLq7u83gRs1zujh57DouXzF112HJkEAW5Ua+6MT7FcXNF0reL2+e27o5011h9wOv
1JOANQXyYHkN6YC3bmqww3PlBhopBSxHgLUO+5UIAnPJkOzzoZ5S2MRNUawm6hc+
1RMfnkYmj0qvMgBoIplUEfkYWohnwHzsiz4F4GuYYMn5+c2OZe4ojMneXTpLsnQj
531liVqGBSAqK3b2HmPgK/GahANGr8dsjGPjUJ9i7HAYLaadCNA21cf/9o1w5HS/
l5fU5lA//xxQBTEGaZX+Vwz6DarY25SxczjI5OTonKFZD2Nri11g95whQf6z98Qk
AfWOkL1U4tmE4a2uj9NjKmgFkq0ubL3skJy9JXYjRKPLQuG/XDTGca2dZUF2Stmp
7CvpZRdM+lsNOCMqqye3c23lPMDCu0Fd4PIssplWg8iGmpNlaCUL7da+3WE0Jl/a
yDUYmXmfwRuX0xLEmdg6TUoLKoX8QNCwRQKevtO1BcFBHJ+D9kpfIOVhEJSNz1zM
uZ8DbqfYTENkAQGUflMfBeGWOGWEkqWNPqJFkdqSZbQtxOripKHp1dAvmGNSdnlN
YdHLGhTabCiMUxEqtnZPI1sYXCwGGl5LPPWz+t1TFGSBod4BDvAr0kmosGFHHvhS
DMrOH6CKmZug2eK8l8bdFximV9kfzaidRmXh3T2YI3jTDhl/Bx3BnANOaMyNYWKq
gbCeuHCqS89mpvuwfap8obiPWIIEQmYKtZlRP14rOErAXa9631Ciw8kVVT8N09OB
AgtlsVEOkXxBSgP9VIMreVAuPCLhZiIptXNb+QNJQF48edMIX5M3SBkMnbFzEKtq
QnzvZQCbYF29eYfjCe6jLWCMSw8bnSBQvqS9I1Mu9EaMkkxIJKYQ6FFTz1ZDJ2d0
cInobL8LXkH6Ml9RQ4Jtmvpgi8LOEo/CkxEFCcbQbeWh3WHavCYsZKdGUXE628V2
87c/MlEbfvMgEuJjnNcGEmki0pZHJqW1OrZkBkKaYSl7NnJyYfciDq+ZElWHQZKl
3ktdigzWzZwDzzg3I5R/LCuI+EkqfirlHXxIdVbrQv/41uKyWCJ+xf68U0XK2M4F
MGc1ESQQcme6njmNaX9ZpHAEOgzZYK3HWYY6eJ9ociSTu4nVfIvM3jLi6te63Z3h
pR/7EVjj1pAsunbD86H1EJ8jhOhapNXRHlGiBFFmxec31HtLAFvlmT+mXRL45Fei
Kh/lx1nGUWpKaa8/qg2NIcdLW3FDGfLjnsU/M8pIxvnn1b3qFrZG5ouln0/58Mah
viSr8FHTXiiTggvPAWLbBDNj6KdAVWeaqSpajxOA+fxeDv4AIrUtSTl+qsD0VKPY
odWCeKODmcbHgiCpcfx0nIV/mqVX1kvaV8wDFojjYJx5UlCMSxkIq3z8fKVSaLG6
uT9m+7+M8r/H8iALAUf8TDdWK8gL2Hqxdh4v1UnMnSe/UVw41OUsx1xa4DGm3QGm
+D+ABmorkjYZZA1ZPxyx6ID7Cpzu5oldIM1tvUgrFbTTFkCjJbQQZto/Wljcy0d2
M1H9Bs89L+gamsaGLxOESoLdPixBvN7MtjNfEn2KwillX3RyGd3lihR4fZ0hkKsk
JrNZvCLfPRI3OTtKZUe7Sx9b2MziRsZmpgAiG/6WSmfA/2roiT1ew1U4F41CpN43
DYlHuLymGehej+LaHq5ALfoGBVN8d2hNQXG30wfy5ih9fnZv9h0ETFoFz2SE4Ohr
/F8cvtdaJ/6vWzRHGXPENNVQUw9Gllh6+jBe6k640CXMWKmFXsOe3a8xeEbhksqU
s6NDxGrFfPsN5WVxPIvqtgp0xvKEkuOtEHvf31ir1JpQejAhNck27DJoHvQ6q71f
S/pOv5EjRaBMBnFuwBO1Vk/6a79OG5Y1GUClxbw5/A8YgGKzTEPPctdIP1aZ9qLW
hinlO9f/Unqs+Xvh/YUWyEJ3HM4PRgSD0o/Byzt0X1Mb/36W8onw08TFLzUdghkx
oNXtsr78ewreewakVxiWcB6K8CtDKt5fy8kiy/m7xEbKkyDdN3hDL7XkLuG4Tr4o
qZ35aS8Cp26Q3EievtukqKNM90ObSTKz1zgyb2eyQFfXJ1Jnd7TlF8s7Ee1vSkne
BfBUoO5dxx1lY4WkybKs+/sMdoUi+UuHVloEpQwcnoRR9l2L/FpQqA0EN9UtQOFi
MecEKRykyGObj0JRnQg1T/1DZc+yNGaOqrDBniJqTHwQrS+R6nLz0oYkgprE2N68
uLKUFm6EwwBJIOv/Bjf17W1zKYeZwA0k+pfCNBJC9WTrr1Ie3/o9FGC5phxl7816
M3wGfSVwlNopJiqp0Xw3X4+VBRldN5MOBQ3Jjs1RYRKuyY2qAK9w2q128HcaFxB8
pFVUXiOE/uEe7F7BmGNFeLBr62mAP3MKM3iNkg0TJr5yTogKtBtKnFtY2cJ5qdeC
yOwsp9XS3l3HiROjP5cwfswixu6OUnFPYWUGleDhMQ1DpPDEF1Eeo3GZKbV94Laq
qo1H/3rJ/4FOQkpbaDCs43QQ5WQyeaAXxVqGxrx+w10El0vkY4l8RdLISo6A9EGQ
CvSbHl/dr0txaKvbSUp/n/FgtmjVlH/Vu4h8r1V4zI/njei1hktRvs8MBayflNvR
NKfTPZVVBboUsrnpU3kUDvbtNOcEh3WvIWX91I9pd4kc44FSHaY09JgRnvlNTxjj
MJXYsY3gGJbPEGZlq1RBrsbGOOu5XysiKkWvOKNEwpJ2javJwt6qGE2oXxDC/LRn
7wHehYafIVUA4GCX4K8pYA/dkTrqHhP1tpqpUuMLRtAblcoxEY6BIOPHP4TnXN7A
DK6C9IoX7N+Mt7N10xCwPymh0XyOLi50KWUHHc3qyMDswqqoMmwvbPjF/RwNfBCu
jSVGC/JHR7eKHS8fGvaq24zk8QKRQ+yuBJynEMCkVcDi7V1YSAfsq7rhE0Luxon7
foEaQclGiHOoqpN7mZb2kBZnKwx8lY8lYBJ7Jtk1RrZnOtCV6zvHBlgaM/ekIqtz
2zXdJxCV8nD2Mu/q9HkPXSAXSqT/WcagBXVEZXv/3ndio7KfChU2sb/+ZkrLXVMX
yBfE939pxAHwoyrIQeDlAVSQquyNwjF7oI3tzfZIuQVe05Xj/IZuvF0qcMwqCfur
knH98laWFrK5PicTdj5tPbhsOiZDVzZ9wx5vV4V20umc62DxmnridE5BkNpqTF5X
WW1WYq6NrOBKRm0nnB6FbQU7J//HnpPpytZ123hpx7k2rdAyxOEm+1zKCV7MzQHe
SQzcjXwBmtuA8mdyhlf4D8U9geVLYSDYPFOvzENccOlC7UE5S17Vz5nOiUC78LcM
IzctNpBYio+ELgNmnV2S+zlUe5ELNzw/wi+fYnFWmBOyOpK6oplEJ03K20p4Atf4
HclTKO3br7qMhWUr3tljczmg3PWP7I9+UCAMPCLurNu+QYk2+AI6tstCLjyQm37B
QxialTTd/BX7vV2IqIQK4CJiQm3xdO1U56jCE0NdAtEUB7LZEsr9aWiTPOk9d7pc
w0YRE1jqGNsyh3qz4863YznwdCxNrHhhWsisGz7JpvBdD6cGYfXSbISVzC5mygbM
ZsvaFEY7gx6OSIgvR3PXms1FUL2v/+8KVCmbzzsBQbY2REVu9eQzLcFEALZo+tJ4
REzqcjx7ujnRcFF9FdAoMbT5Mk+gsiPc8d1ipkEyyw5H/wSNSeSlDCbLrbM0jRpt
3A37Ps4D+GJdqUCRDZcSwvRcdtZCmPZtixhQCeJXdErNPLiUDHXTD9bZCsahQKsO
X9ZEvZe4iygNMdG6Pfykr6NmC/Wwt4uF/H4e6e6y+I3Mt7rwIM4AQf2qcwZJRbcs
/I9cFLrzuLaiIO/EAcG+lqOIwCnjJwOxMyz703A0hAVfmsgJZH5W93Bcd+Mr8wYJ
X7vcfKgDLDa22j8z/4BSb1MUzMjYp2bDkDyv26lE34SuwcHI2iNQChpbUhKazawK
nRG+uZV2OQ7jMeaXbr2tDP3x7eFx+UpZbd8n2PcqUShfalrUWGc2YDaKjNJEvH+b
bczmOKLc4Q8nJ+DNsESq5bh03CzjvpIQtbzjkB+0iNqxTgbcyljBI+DGwHZXpT3+
kcsWHdNMJH2qBC3RQ5nHTYAlWwdNHnJhSE9y9oeR/ckRMUYCuKhaF8mFh/NoqD/C
Pr4uXvSVFSR0WuGg2bet6EKQC3RKEqkmQMj26Ks0YCn4hIaMlZ85fSPliEPtm79K
4oDsvVnz6dDlBxVsTzFqOYAPZqz4Ycy2lG5yos9cmFSwYW3x2nd9YR5nuLUFMGtC
/7N7llQMwhrr32gnEcAXUyqkSeJrC5uPnV1rzOf4oYZteqF4+HmtMmJAuJ6kwPlR
mY0CJBKlZqdr9GFkZwrUdJzdjCbfFWel8KwZrzJFnGPDj3naal7uWL7eKmviXC2d
9SkHtGvn0DOcLhre4tn1Z9xu+CF8A3NMiPQ6M4U5RCdpOZguKzdN5+B1f+CJgGBY
oPOGJZLPix8U0AEg9DXZKRWl10roQvh9ksJ9jyH69yQkpexdCEGnJ5ZwCRdooB9Y
eEGKnRTBBmrjCowkQepUlDhh/ZUto66N8pN5CrosjDjp8HpZKPG3sq++hfgCSI05
L6p7UvpC2I9wO8WEQdFAFnoQ1Q9dobiBhGPSyUMxZlaRvFBjCoclH7uTWIQlbBme
FG9aMScmuKyAL10Wh51QjLh1vw8BdCbLieLDPI4oUGS/iCqNHq71nlvT3BvsosVG
Qoq2e+/R+kRM1GiMF8qwrvSbf5NK3nCkxq4YGjJnk5Ha6czDl1SeovRDOhTnEyBC
pKNVj49WUjYi9kY42AUYSMFn/zbl4UYoF9KpvqFX7DQTga+/oMkLwhAZpnVDIkWX
yQ7I8HxSDDo3oto2bE+UkjiRgJix7KRjIq3eewOby3YFnggDjFR6BqdaIL47R2m3
5v17obvTl2Aw8EpRLe1P2/eRVRH9HOukM9tdT1M9fozAZW5orAjWjl1wv2mGme4G
qIpocW0ZkiWWrbrcUBefeq5SHyU73K7i9AaeZZILtJ+RaCkjsRMEvjMucaju24JM
F2Puw5/iivvETMv4QosiQZFr5h8RjuH+VjhU6chhS/GOMF6zYZ1/f6+nC4PPiylL
7KJHXjwPup+TGMF2SjoasolaXxK2vJZcERUIWgORyq3+KY87A+cxjgsuLEavUSdB
+/cSMnzN4Uaip287j6C5JMAWdkHy3dE9caiWWnKk8OBDrtHo+3DxHGOxFvQ9uUya
5wDxABdGPRhEhbsXOQRsMM1I985OU8Rr+8iyvB2lzoqx+4RdHDvXx/usMAfrksHu
7WS8MIZgRUZGoGnPTtRSOgkwsn32Ae3bjQzK+9nygJPPLhrN6iq8pOcdH5oM3rah
OaS1uztEcimhwL8pLweE+/OAbZ/dxu69lMRaS6rsY5/eTu62xU03EoZ3ZoYQxxfp
XHZEUvypt+SjV13yMLV9IWYV/xA8PIgl7+lIgIEPhZiTY4Kis0KzV8Zul8LJYmJG
WLHPK4RWWsVwvzlbclay4tR4StmsqmsepyWCVsLXO//5rFdhYo+zxcuin2GaBeOU
BztKL72OuZ33roh6qJ2BsYU4SM9KxCNtDIY7Rf24n2yAQVsJC0dBGSLyf0e2g+C9
XyiOgdAfAEDyj0UpNZG14xq4r7ipVMumT3oh43s8dAIotQFNa3FPVN8nFmGfW9Ru
V4VcCUeXlCA2qQLWOGkSxuCPvmupyk1RIwHRARXLeRtpUaKAjEDdUF96mXmFfxWc
Pk1yFm7kIeTDGOziP828t8cm1SjSGLHcqe+9fz+Ax3/xmH57iCXse9BjHvJN7ELc
T/8SwJQPGtU/NkzERAekB8i17shIByB5kRR37CojJdpEDYxoaKIIbrE/gsjWYMnT
OYAAETI7JEj+Zs17vwPW7NEAjZoRe3ZaCz1Lo6iZkR4OaQOzFgEw5EdylYS54VZe
29vgnzn3rDnNsMXmth3fub+7Ch8dtxBrsJ7Ll5PABYmlXEKilBczszi7okCLAkyz
IvUPziAAeqm8t+01N+uQ44hnh9GKxcA3fjy7tFDfSwgV3aiK3GhNMKV9zXHd3r5o
rqoeoCKbUzv7yLGYAmtsjol0hXPnUbHKfCXG5E0+qd2iaKRBhcXk5qzvkecBIjl6
ASB18N+pcTyHPSlJJFmjrzusyeAU5AwLVoL1tIYQkVHy2t2AjNZotZ0BQQVTOqYS
nCUpagfscYG/PfL5eQsfNCQYo4Int801h62+OrnV9rFfPvXLT3q9Nq0UtMPH4aZk
edsq5iDyeSlajW52mUydYETrJgdoqGBuqOwN2kCqAdOgU3V1Nye4BroFClicN92C
4OMi25M04iDJ1vmIdwZMxxaIYMmVcjp7aD9kMwBy/Y/PP/uVrWld3k5WJWAkEXyF
VfWYFjOwM5J3/TOEJ57YW/62JaP48Wrhb4GdRh73DfliMzU7hX1iiTrfd1a4AcLL
mGL7/K+EowYgYk3rb8iKjws/b9fNWizVwbdlVkitGbmRLWGREqXTw/TW30Kx8ps8
29HoP4LvJi+uxL/bbNCayTRS+WeNls5ePEVPMaVwEJF4fWk2eVAaiK8lNvD/Da3B
MB4V+0mwUCHAZH0Fwr3YsUyR+Mg58q9XNkpOkvQ7aaCTcYd4M0GDtAvpIXZBFi7q
N1WGI5aIbeVYVOoyXyEmDy/OQkVdT4nYZB+9bxzrgyr+G7tf4yMx1Sj+m4tH3the
/2i8rHHWDEqFXjBZXzc5axFtIAXbNPxdc3opgCPON/Nr3mZ5ieSvN2oxfk4i3EWV
KBLCD9PCALfCkHO/DPKUsDa2IQmO5H1Wg5w3JS0uhvr0CRCJmYy+9FESxPBUFquN
htvTNs0AHPUAG7TM7BId17aeezlP5Y9TQIBpr9izbx+/dksIL9Lk5UzAoWsGRVIv
Q2X2axh9odY8RKaIchvfyfZ0SIiJh5EHhweDfJgr54r4r0ujUJkFVaHDB+dHfCJX
QnURIp6ARFJpsoHQgINVEnzON+IJpINxq2NP5i0o8uBbIbX/W0RRgA0sHd6hpqA7
gwK7cSNrh1XaPPgxkx24AHcggpatX5GdFk6LZVuFJz/o8YXHQqGAGetqC6NNPQ96
O67Fn4BxBQcPIV25pIQupXNOC1apjXYXGm1Ok5WFVQFZjiIVGazP7qiX/f2oz8Ux
wXxR52E3IxbySOod8iDbXFbUIcJBS5YCnpc/LakLfyUXoW5JdTe9iONFSRD7mqMQ
SH9tPiCE8YFGkBa0DnnrgNDajjxe0A/PhbyyOOrGr1PlwB+m5X/3+v5vE8ah7iVd
mhuPL700qVgl184lWhrywjyZIgZGwbpQd/k58Uo06PX0U55S/e3sVDlSSldQDH+9
LNEbBkg/rqh7oTrdAMR8kJiFDkr7BC1R8tTlAL7c6ofF4DjW9M9w4D1lHKmwkYRZ
tOnVsnMCuH1RaweMIiSpYjh/lox99qvKVgiSS9DVVxFz4aydI/rzV8QX8L26h917
TYKJwfZVk4R2y95oEXWG2gYz6rf4EtEA2qbQ0iBMkZVfAB+xKuu9YofVP5kgxJau
hQG7zbdguUg4vBnDHuuYN+Yq9T1VgTbJhkI/YRTZq/ZjdcGJ37YWBbxaZ0Wth8Jv
zFCqqy36a+MEVnqGkbU1censf6c4vqRrsx/g+w4fiGmTJrLCGTxo3XWGdoVe2USh
A9tFEeoGDNahpLfsBFmsMkXkQtWMmAD5+d7l22tAzhR9ZuqLueW3CqQJxiHAwp41
Ayis6daumVwP0QzSEooZ1HGk1abCExs7lExymEmNdEixPYm6783aY6nhnLfRfO+A
JDe9ev9UE+iqwYYW7jm69y8YYZEsKJIL8L8mCaMaDMzF+Q6xDYazf30ckk95he1v
uzoFBia8CLrRIk+Rc0WaB0nAbB/BbBzKswVGXwAw8XubcsgN88ZUorx7oThCPpKS
xpOY9ZwqXOJSr/w8zjDSoBkO2cbouk+9nNamwr3j9gmfvW2ud1NbRx9tRT7V+HX9
3G2qaX+ew2iBWtqA/t5PGcukAmAcPi/m5tbBRoujQ1rAAKkjYWJ6sxwywrfPXbrq
ScZ7mZQNV3WYnU2SquQEEiFo2eB9VAlMJ4fS2SrMlE2XNDFOvSiYoX2BLgkMwdDi
OgbtXR32sb0XUwKicdyQPRv3pDK4ZvaklMjVIFCZG1lhTiXM/mWnV5ZznMOw5SSu
4jKhUSMfOkVhDjE40oPkdQdLa0ORR+6/ysaDCx6pka8xSvPnLY+Wa1GteHxkG9ZM
TOwHrnhxsFDlUXHGbdgoUl4xuW+gGZUdYdJpUyviNZp/iQyGPm8oKM0QCCgtFT5P
1k1BVto98wjOOhNi/nZ6XBhB8Yzl2T5gZ5iHg60IbVtoWCT5fPk9GHi7MyWFiaFq
gA7HYOnxFg6wpKccH1oTPgHNeZgA9FwYZngL1DnEyZk9Fs3o9Q82/su4HcAeKINw
10CMDWv76REPh7l7DmclELLAt2Pe2lt0LRHp9W36mwyZVtUzFVBCQJXp3aU4VDl+
HJX4ZCTTysjRN+fdTWYm2SsD4VAoPoViXpX/OWyo1Xrxx2vrmMqv9oKxoE9s2uPX
gEG/WYryUKKqraMMHHKRVxA7SVsh0UShc57mrgd4qjCwOcKv4140mmOI/UmPwPap
km7RYG6ysJTJlpD+6vq0uKJZXQcYFMzLO7ANjiAVyyCLlMuTOhcXZ4kdBJq1pKxy
ucgqDwYZ24BfpEGyJqJKJfjDGTCOUSFHmO3UqYcwaH03TFbsBSz9Uwy1Aa9O290S
RkqUijhdQnojKgvzfb18jqNXTn09dIZaWNKwLRJ1P8ZnOdql8Of4Se+CZQVncE0Z
x4D0mFAceC2R2mKxzsbkFOIBCyOn9qpjvn3b6ZCror/OA7cxu1oPiWo5gyHhCd37
OegIVAXoF9TUULCi05b87l4TRar1t6RIbO//366/1GA3uvOMNy71yw2BKaLZBujO
mROtnb5ej5RvqZVg6oiDP7/CEebaNHW8gI+6pO4RSLBJGTW6jalodn5+IJR3kQSu
mrX3c96uwsPLcYD1oJTGWN6B0G0GU/pMk62WnaGQ38B97bgnSgD4yplp+Br9txPv
dzNv0KlNhX3unVFFghdGNtvcFu3diTGdlhHJ66I54+1ifKOzjG9pno+DJpRZ0Xll
nC36SITykbT55stZbwjVX8bimA+SJLgJDj0bMZ94daLDSJfsnozxVY4yvjsL7kb2
NB5YCzV78dm7ariBAZrQbHvez+5zRi1Jgv4NriUVCvW4LlQuXu+B3DtuYhf/F1Ny
yPJJtm9Nk6XSMFbFgDA3fPZqf2KOdG/zE7HUBN+NQkijLDBSn2arG9i57GsYzDca
fXbMaiXuu5QPmCpwhxN2zWF+mhWoD6vsygZl781/YDHU8FMZvzeT9qhFJrDI4Qcm
jJv01CftfJHUhkHJr0dPAQWys7lE8alv9N2dybq4MPnqX+wiV289NUaYWzmF3ZLH
CdEAKLDj9X+gsxZCQuF37H9tYn9uRt9hmRsbQwpw6JsZBRfntTEn/t3qmfc5I+hC
9t4XvACF2x6erhWhhJWI1yS7JncMWwmeBFMK0uPExR2XWu/RmdNH//m6KKm0iEfz
vG7IefA8sxXuXFgViLFByzKusXIp3Y3F1n/OMF86ymwZU5djTE2ps1gP9y+hg888
HSZK+5FCauxuw4Nu3itnxEldS1sMWHfpcBluHRRUrmQaDaP64K17S5h6zXwMGVCI
AZ1GRE9f/UefyT/XqWi2po+CEJuzCitDEWAVto822/xBAdbpRNPiqTX6CsjmsVex
/fRrxEdfJHKkERH67u1aofWRBLfwoUzirZ4cxFU+ILa3wrhqZyDIBSVrg2ZJyARX
veyiWnU6WQOLl9xPzoCgtYu3HbKH6s2LYp52mJId+djQpiQRnqYRR60oWHC8xtj/
2aEHiGEugM4SjVE9zJOEzFu55LEj3sUSRDLcQ6RO+rpENkgYCHTuXxYaxfh7Fr5G
HzFtfzZPbuPajrNIJwRVjVS8HVYsDnBtlQG27ox+8DYraztSHDge6jPQmDakm0ab
lUY3lw9qY/2pyvSJjhI+4xUKu/aQ/re9vOfEknC1YyGTsWguE8TFVA5ijaINRSxz
tB7pinCGS9pDgCArS0O2N2g4bOVtLb9y4r9AIDyhQxUkawlSeAd1yFO3MixLbPDa
Q7Zj4GeVdl7v4vQUsPn7a+wtCqgOZKODb0JRhCwA5NIhAD+61+/25U7cRuzuV2rl
VMucMSDu5QBApWc4nrTcdTIn3WSz9qHfau5l5RAuGxc1H2AzTw83YzlzuJnBqPNW
SvhcA0fSvTkj84snslTo++Zp9YZOfSlQVsJUAsOiPf/ZdHbTexo/uAGwdxxq4Agx
Cg6TyoZvYgEITggo7LVtIXETewb3M8Li+g60q0KvtAGJEcNCIQ/KU8gtGUsqjFaw
epq5ysFNTQbQZqmMr/r+z9RfycSb6QSKVUwI4QnRbcFlvDi14FgJoNJTkvJ3qSOG
pYIRgb+EY0tVrdu0QMYHSqf57AzrPWpDe/LP1d+4oNhrU5g8+rF5cxatDEHQHMF0
p/kv3XqluwMWUBirZYLO5OXEd6RcVibL1ZXtaml3F38nx2qYXeArUWpbhbP2y9X4
ItIzwK7KC65eHw+JjfdeIRO6OVZbGFcUzaCXm9l7/W1pcSIkuKMiAATJKhNKu9Gn
vemnQN/x/1FaMSyr6kvcmcy4lHknCjmWhB0gC6E/EMND/XnTwFRInAaD7qAjs4gN
cSpEB0uq70XcIw6rsrzhcFs0QSHJvmYcyPk1dGPivNU82pPEowRStFrlbE97D24f
/vMsxRWwnSTV6K5J/iTVURbxXJtn4b9o1kaC0dPYkRalBIxyjH6jikY9gEuaVlKI
wd2thFzBnLRdsMOT2LSOORC0Vhq1D3R/Xcwloczt9iHK71A3oUVShqDmCwQ2ruzG
O2CUT+0JawBay2sae0DUz5MbIFBHH24OUmd6MoL8Dtxwp+kuYcLV4WZcTmexbNGc
bvtJxgWAZZkUDyoYPSdrsSwhiHDhIjuvftJDqTw+0THpKLTudSlZidunNuPF2QNV
rxEUcHL2p+qIU0mkONYwHxA0kN+wpaXJVYbcPdYHg00XICO1D2NXoyKI6vjI7a/4
jb80ZWNSCoCecdXwCl6829DNH2LEXoX8/tzWEDFdUcG4Bq/vX20aHfj0mXylB7Es
3Xxr3Jlq4hvNWR+24MQuwwVr3nYvR3iqvkSkxzwlwoslKcqZ2C+RnRmqm6YHhCp9
wLhcbJdFHEEGtvIskCW2vMqs4oG5igM8vueZX+Uhd26xrjbWaYs7aNqxnyqfjvXT
GgO4zwZOrJBP0j3hG3i0YcF1gyVGxCgRWtNmHtWx5QYhL+PcYGw7y5ygNXeCMMvG
hdpAJTvonDurtqjmcn8lTewfEhsyY6raia/sKJhLBTRpMgRuYFKC82J2XgvXtOcW
FfTN3ZWU9m3lYid6k/IebiVJwJLjPuJDlpoLmgYQl4GRw0OMKA/IiMEZXefvYG9D
AfVFOaaxIKZYIr/O4Sx56CRTXzYMpj9DP+LqaStLqxUdV39bWQ3Q2ce+v1SWady/
J+pk1A5PEN35uBWQ97Tm4Ej+xpLK9RV3U0VV/9LR8HoCJjuGOMZG7Y1YfjVCNPAj
SmFZri0xS+La05NvXg7eIIDBEMvRgoXwYwY/gjLW0IRR4nY5fNL3nAr5FxNluu8U
0uQVYtN9Rbxg0H0v+oN5oYtIip+HqDU9CkbCMHbJqeNJ6TEHuatzbGUtbh2nAFdE
KVRWIl8dRtEX6kcszdUq8Qi2jOFm6KvTe/1d1LVmaB1jO3WyFrkyUY+JshFvo2II
Bulhlst0wRC0ewmv508bX9ww54PNoKBzubS8uGnMKnLoSEhwXBcOlFjW4GIvt2aC
nXCx0IAX5PKCokG2tu4U1t2Xxo5a0laYI1q3/dGzIUK3n3Oy6IGWfU/KAZYIsd5l
yoCplQBO93hQYDRy9qrdJaKjACpqqgK2nBENenYpKvuM4J6xkuFypY3Cpd2SuiXV
MjqYV64vIcu7QARMaNKnhhM3R1+dogEsNoew+yxNMSwgkGQ61KSc9tcNcDHPhqdR
p3/nAY8utGuD+MpnMGu+rSHr5wjBSAmhFRFSFcgCFgPuIpw+h6LGPmCogHfdqb9i
osQk11O4mys2vf77oU/GglrOH0jSfFXKo0NFFBix7xnqFV8v3SOPU2etY96Ezj0V
0TI+XV8zu3xMAbejNTrQmSTrLsPsX2Cwg2plMm6YGoA1ZtdKn8sY8aKdiSxdmEhJ
PA99fcxzeakTN6Re3DI/w6T5EkExwJ2wVJtmSG0Mupq6O3TEPtQbuePPQTBQxy5b
M4Gnc/gwFC5OsXSvPEQA7B0YgDQswtAiuOpkSDzexi9K3nQsxLcjT7U9JzXEDrSf
TyDlAaH8YKF3V9yv3rzWb5Pwd2sonJYGuKDheEM6X8fvhiH9tpVGGJ26TRn7b6vs
jqiMVoJaAiCpznwP5oF7LgHDtTCYSQwR8tc7QzcFKQA9IqTJFLlUk2J4wMgupGXa
wRXnf8kz41XT5OfxFCBquF6Q/IKC+qwxNNuew9tSxYc8fX13FiOP85x1TpOYwqVk
2jPA0JTUNWbeKkmlbV3D3WE5iuffYe90v13IDDI/iMa7A9ax19PRb3Y5Keh2rQ6r
mQz9zA2R02mR4TWNIOX9iVRA6bj9GiEdFYksiJQfV/05P4Z8IYZQIQzB3bd4ZOnu
p6LRmIuMtnd8s91O5+P+f3SD/esRFAomO8Yp72MX3m57fNl6SHdagrI2l+lrSfUm
pkmReTfBBQ0L5k1U+cRzXECh8NKpZkacKdJKQ17j4+qdbEHzGVYkDJ4V6alcL50d
/9XfdA40jPbzLPVjd8knmsi7OJeVYqlA537K4VdxTdTXWm05gIr3F+TFX4WA3BVL
wp2cg6BcZHSDhzyJu1y5XMX1YJSAFxC7UbwnWlOfvXAyAfpsmZ/uKmjHgvuY8Quu
yqX1sIuWoPbLHWFUeBfbFw3UCptc6W2mTcpqu8jotMbynntV/0IBlQLQzvS/kgPy
`protect END_PROTECTED
