`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txPd8wnMPwdfkuoc+jv5VpHV4jV88GDv+XnHMaYeweFhC29GqEb6Mu5/Mraz764z
G9guM2GJFEnAYGeEfzq5jcqxlNCEv7XgtPpugMhmesvtMBLyNic/8faWtcfn37+C
Vl25beq5xw8uMnDjTI3NdqyXdRuBu8PRyMOAASgWyJX8NuRRn52eGLJgwPgslsOs
mYlMxEng1je/WuTN9McV28fdE1ts4P/gnu0G74xqoJozDVhjBKjvr6bUbDykyqdk
4kyQs5EPvrSGGxQ1MxuxlkhyCFOxNMNUFNl5HL6NMnY4kkWs/ZakZvnmgBvtdW9c
srYzynoSthvZoVXkVP3G0/LasB9RDT/C17UuFpHj9gyv8qVUj4z06e+bzbfC10vh
9yV7do9ZROCvNee6pe4XZypeSYZaJp9HTVam86s847pJ6bUHBZKv1YQRICz18ixS
qFyCdLbkUMk2/gaqCE9Z9XfcdoP5u4UcduK99WMz4Ue+uKNNERR0yVe9NVs3r2fz
qx4t/soXiDtvn9GL5k65bNQlY7RT/ca3dkQcCE5sV8BC9zIvgAXKiEAwDG9/vl/9
`protect END_PROTECTED
