`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkWdZYBtmOFMt2L+Eczte1sOej7pnHR9gjwsVw/gr89zbK3aYjdzQJ0XXZgadxbJ
3UMnsG6G6atmOJ9xcnoa+h6SENzu08yxaE24NFzvNlqGZQJXMugfme3BuE4rPfni
2XXR0Q+W39oHW/ftHbLGIQaHF7MViLNN7W7nO3nISSoFtk0EObDuShNOLbnHyJOw
WXTYdzykEqC8rXt5a7j8ao71+8RFV6tPMByAAT8gYsxQCSpeB05iLUPzTrGYUnbJ
lM/0p/1Semg1fU/jmGcVrFIcKCI01Sg7vbP2+YjSE6u6LRMdIFnK5aVtZ80xicAJ
SA3rxsH4sdpboIhQbGhpWVmgJZFMCZrFWG3oVTwMqoyBj+6kCody4CJ9NLVabOpc
cnm0KGBat0SH/YfzUfZcgukbjl3bd+WF95KTpHzi8kkhzCJSzVRPlJA0p7tltWuD
WGvif87GiWA67un7U9ILsWHW1jqG43mom2JIPz8eG+DmBpEIIvfpb1RSA0+YWX++
xUJ1SZIZfhpclvrA4ITS4eZjBPDltHOK5H+oS2sh0eaOqm3IONp9Qqo4a9QfYx7c
77S2BaXRJRvID7grvEW5bMAWIcJvcghtlxIHz8KyH1PS/NCqNExffpBJt7mYnefw
0d9rapFkwF0P51vMLs22kM3ehNGYmKkQ6BhJMAJX74EN1uNx2RGsuSnJ5rBytKTD
4ILCRHYMMegg53KSbI5AJuiAPiaSz4W3UcnF4qB3mYGKrl0xYr3wOnO26yUyaW2t
GJEv+xrCxYJ8CkRuJ9g+KahaNq3CgrHWfDExBAWijDFIGRudjiEGHjGsJr5FuEqZ
hoVvPd7Y4MuoOwthFNd7xc205FoIlXPDPqsiZKeyX6n6HYoxA6vCDua8LWbPqPnv
lOAcjsbujJvax5b4HMjSoyJNTbtzAdSmUoCAvOoKtZnFI8Y9P/RN7uHzR/p8ylkd
sCKngqsWL1ogeESAcj328ODmQAloY5qmEznhhlibpJg+R1M85KLNx1JTrRxgXNJT
RxDW2ueaCVCtWH0PAdipyTX9wHp5Xrg943eaxfjTlUJz/Hz3i1r+RVvzk0rjw7P9
EJphb/DhrIovNibP1QA4hF9/T70+claGwHcLPIiAdsexH8+jS0P2JZpf/h5jK/+t
WGfucVdRnkY8mmkI5ak11R2lhSDW1jTEikP7Jjdbb8V41tA2nBqpbtzi3JDpofs3
Nn11wRWhXtLv9Yc3DFvLEKePVsv2Yqbf2b+KhXxdLGDy5vuTgdPGpDW1N/5hU1GM
f0b7cewZZnIB4jHSnpzvlNaOj53dgF91p+3QvmyFSBfF/ZgWNp/jtARGygEWj8EY
yd/SKYRSKaicHSQIRVqMooCyJ5wyo4OJcHDh2FHZcBhxx790GJfTQ1K2+897D5B0
EAHbOi7BcaMbRVR6W4pz8w==
`protect END_PROTECTED
