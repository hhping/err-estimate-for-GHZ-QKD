`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0h0qKbLS/E1KC+mcVUQvSzYOKXWwB2fTA+dgoQqD0zFVKvkeEXM1fMlHo7YtgHtV
BtnosdJ7Cr1nSl/qJJ04li/NCSsTwsUHUR3DbkGsYSwNFIPLGjV3Ody7IA1AgQW6
SKJEilBRRbRgsWQ2qG5ouNki1p9TrAsEEg30ErhE8RGyqfTETBhSkBfM2sLkZBZj
aJxqt8VBjmKdqpHcWQ16M8zPmEYKuSX/lWB6WLDEFczrTAZHO70qJ8Ei4ngDhQE8
/t/qe9qy+elm47wEyYXeZchujkQXiS0ayjcw41SKl48i9VDSdPT/uqc7Jy7eQKk6
fMJbNUZJcPXeHv4Ei1aOA3AJSM9LPRlVqqMqIDrfjQEfyfvVq6LewwUYpnpJxUXe
8zcrGxiDWc0K0+qfdzhFYvrxrMr8dzgepdbhI5TqHepvkeVIQB9hXiag0RzO8OT3
j9h3PiNcVVToWIWLpw6uiU8yA/PG7jqiQ1G2AZuG/tfdybXQWqX0Rd3w1YR7Fg/8
7GaXcdBD/dobmhzcDmhWdq5BVRxQWS8e8srIkBSWNbG0ilIFy8SyCtQbVaMys8nB
FgA4SIksabz9xVrBzLbRpT39qCekRhyVhcXfrQ/lvhg7GmQa2dwTVF8zcWyH8pnF
9o22WjkCfo3qePIjNxYdLO9URLm3KtD1cAWzbAl+Bwmrx5KhLbeUg+NCAF+R1cnR
jpxLhZ2Fz1HH/qxS1eocq/z8wS8BCsZQiLVRvlgtuLDEbt0XRLLG9RJKHaPsi1ja
t27V0a9kn8M+V/MV+/xik3P4mVAxHTFOjk85WLaeDDShtwc1E7kqlfyIxM7ELZ7b
IIyUYrLGuyXen0HE0EKLEJ3f8YkpjnlFrcapRDJpMFKmeqcy036NtGB2M+BdADG3
gLX8AAS/+PgdyRVmxcMh/s+3RWALLPkJDP1Ga66QDRAW9K40X5LgjYjLvhW7OM/Q
PBdSNZDKGEEG7UD9pzsAFc150/ldPrUZEY1KxET2ifcqzlyA64yq6OCRoXaIynuz
+FxUQ6k1LDlr60hsFZ6HGrLd34wxL0CviPvhFoXyO8MFepUepxo3nFO0h5FLb8gq
euQfySBQKnrwDUhTndQe5ZTczXFzssXPUUAQnw73ZAYE74oNQg3bLeQTJEo/co81
mZQmRGwi7hnLGakBK6fl/ZiOoH66bAI88w2sJ7X7TnohVsbnSNM1VRaL485NOeK+
FA+BcRjUywpfigUvkioznzM09RvY8C7MzB50MLeu9uwcqQeoDrAcKSTmxVcJkO0x
x9TbAiwHigN1HgSjnB+etAf2UFN/qu3DmoHPTZ5BtIQTv5UAtpqsQho6y8aeMHuX
mQCRSoEcKhq62esr7NN+oj6jb+8upeiUDcqIJNhWSOgGi+lLOTQ/dA30UNNyXesK
gR7z6ne/8iZhHhl6eUctaUzDjFcYuV8NB8PM3qExYpvKm4UY8y9tstaxIYHJjp57
3QOeciQcnt4POSFuSj53XCGLp666PcmE3yNOA0ywTlHvE6ktPLig9r4rvGqJ12DF
kTWguOGtbT1sE1mfflDP6J2UuyQKuasFz60K3ObXclhyhKhVO0DpWXi/EYWeKRNM
WM41cKiko1wqPEEufTIHzx/yhYVwdmlkcoKCQpGxv7tlsyJxjjJyBc0jJhVub6yk
FUIpPTKq/8aeevd4ZpwXhb1WYNwCi4XTsXSyQ++MFTMfFZj6YYesAbr5frdx0LE3
Xq6ifAu9CX9wI55pOy0tduaj9b/eDxjr3Bfxxcp+mu5Kb7MgFJdpcb61jnIvmBZ+
654nh/h1+3hroTGCo+bJTBQAHNQfMAwTUN9tp14GLSvkgbzCaKTqfcx+Nmb5EnnY
QtPjEfoaQLLf4+8dBEK9puCAQPZ/saqsoF//I5fF/dqPUrDFjOdyvLZSc1yv10eO
y64XXAWCO8xBQouw5dWOtXL5YASY+qEbhihS9Wu4GUpWM4xxYIPnr6/dDxJTKnIh
7fQTriLTAMg3cr9lWdlkEy17EqbwIOEuT1/HAwNN7nmdG6ViiFstrDHSB6W/XCbf
pwOj5eGcpvia1+rekVObzSalqyrqgZxHlJUxlEQet3MaBM2tM87WuaFh6qns0AoB
wQnt/ooqLyo4z8Dh2QEHkxcQQIYVazh6tr0S0xkRYL9qAfHVct5vttam9uTmBYmA
zhoKh8tfO7i0QAuTCjMJvD/iD1G4Z6JQYJxw7sI6yGgkWq0Kl8hbfHYyVXW2oJyJ
2OHn74n6gn1vC7GRRUyqQWOoInVfb3Qz2/qFbIQ2eM7kJk8utzC0NInvtLlcd6fd
dpTxOF+gSGLMScsi6wytdK+eMCfQMYtRudejy020i+Cs0L//6YjXJfF8oWIHmKEA
TQOvciIouSLUZ0iqfi9ic2ibS36PQf44gp9DuqXTlE7qeyJnyCnr7qJZMWgSjEE7
Zzd7xVyxAG+WQvXrmjX1wZmJLabDQRz0vu+hNS91kQNIZB5JNBzVJdEMZWnDhz3u
lMygmBEZ+1/xYWOmJD3I6ILS0TcWYNzWgexsU4ygN5JtVRv6VI8U0IMLzgBCweqr
r1UAXqyHHzpj8RmgYMlOzmEhRXnS3iaBbtx7LViT9VwJuBs4wMoh1ZK0kaJN9QTd
Mbq28Hca6bI2WS0D/seRHL0hv8Q5EEApUU9O29t+JdRY6juvHo3JLwSowgASfHwp
LQuJaaxcah5mZzoBiIeQWsHsmUn7r06rWDu3pOlk+mVRbnayYdsIZbEXUom8XL0N
Iu7rEV4us3RLN7zwqBzrtCGuScLkqpIyNQkHaOFFGbyYypL7+6Lp2GJdfxztslGd
N+PkH4fOTk2TP1bnoZXfdeauBUtJhQ3/3HO+B552+4NotNnnc2BuO0DreMVgQHfW
bg36DRcS+p5HquHc4yOZlXpDzghmLcdeiKCzWE700hdBC0iEm0es1W0qb2cjXK+N
RmAYFi5b8vAnt67s3MJR9DHZs2Uosg2MyeXATM6TCdGQPSc8ZSaF1Nubr4XK/n/K
SS73M16qMqla4gx9d22EmIllJTbKsQoc0BBC/BEtpTCm8B6Ct1gs+dApPzqtHUvm
RsFkl634ombENj/4xnRU3WeNdOIvzTwilBRoacYD/CrPZfnX7m+ETjU1DaE6LRzI
dyZKWdY+psduVXQv/8+hA4D6nFJZ3ThcLYQ7ElhThLDlw8O4kP3JOiDPZN7zljpu
KG63QX+rsHCzGeZ3QOpa29NFBBsjyz0Q3ZI9lyyJq27sL0vCnAgVNviv022oFQGm
LPetCI8ib5ZNdoJXu0LPaQkrkEMcRAbXvV0S+WhzXTadDBhYjE4b3+LY0xdm1pxP
T7+shqVgKG+OX/iMq6SYJQfTpuJegv0w0tjjTy16eSo6FH5cI8YJjxPsJxtHCQwk
c+nsrfTyX98Qvj/GdDGICD3r2HOq3n00tZBHl7M3CletQ+9ZyDkZZr2f5tO26FXO
lo8XqTECcVIESEGpj1t++piZsugdnNoiPeqp9vUhqrJW2Trh2hbJRkTRx9KdGNOQ
QhN4tgGJHW1O4P4cu9ru/zGLHJdz+JV/KRuiXvOGNlxlzk2uLd9XEz9tiadzdXPK
`protect END_PROTECTED
