`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nQUT9Anv+xL2ZDmAK9Lejo0p/dc3rir/HhXpgPjYOlm6ydAsqPDsduK7vYzHzM0
r2yJXieDO9utgSeysHrt/VzoW4mV2WQpnXYwlTsxglHTH7fLLdJbxfQhCVm+fanV
RELFhSNo/Pm0xnYMWP56wJcciZtLXr4r0J3bjrw005gw+G5TKxjWbgku60wEmUJt
o+4dFmh2dbaQQrbFj0RcOxx0vR6ZZPWQSkmIPaZooWBOaXmzg9J520oPYW2bEYho
2oS0rlbpKbJijC0WqkA6ktMsgSBggAJmksZ9BucbYPOxDD0ikgEl8EVNtFr5bMh0
eARJehrbpNVvDSyAv65koZuSSlkMJZ6PqgtBqqdpnPxS/gLDwI1tuF5+eSrLrSLa
IkIKt0IPtj7kMs8uYOi3VrffdYKfxsBP/1ohJZmnMj5GKEqMnfvvMcqWeiydB+ta
TVSz3Sql7IcewMsP4rzI8jJyT/DaZiGkCEAPpUEv/7TFO8BfM/zj9jiKUJ+uliAY
wAYVJ6RTjLzf7CVDDkc4GRVcUHEG1GxmWZ2KtuCgQM4p8UfEDAf26e5mFPWgsamS
8dj4+NHqe6Gzr37kjIaBAfPCnPGznD12LKF8zoIDfosHMfd4CSika09n8PbW1Yky
UFBynuWiIuJFOWal5yHES41G/jp3eCzb30dmBlYtKMRpeGLW0nq/S2Vrcl3pLurb
3EzcfLDn6TgwbPma9c4DvHKJTSIX6O3fBqOAQ5JqDYqwVQzqRa5nu6FG9kdwD8z8
i7YNWxD8U2QNQ8J1tFBwpKMV+L5WC/NWfbyhzSHcnKpR/w6I/p7J5kzoGVpwHD7e
N5A+EP36d1wVnA8YyT1JZtxouAwPSQB7P6MuXmebxXGApQ7CIq1qGB+mmzU6kaYP
pu1NeaZWzF6upiwis8kRPFOBQ0WpRoh6gsI70CzPprfUrTDWjdPAgGz2yy1udrtz
fskJELUor3W0+0zwbjdGRhIt6rLVArcAYlUP4xEGz+kKtBY1mQsFlB+BtUM5xl0w
9eS37p2AWZUc4KBneT/+0nMBoAVXDoUpZUJr1CueZuCSRkZfQgu9D2y/vLRJLegA
nAosc5EbPreHtRvnBRQyznzBlCXuKp/M0PT9uRnA+OB+WqyUk41kTsgUVkpIRLRr
Hr24Zv29lWqKIdJ4jdJT1hn6EWZShYN6akfZ1pniyWy3KEjiPR4DXR5IF9vy+6El
oJxklz0ivTZNFroBED8zZXHlHgzWP/+K9tOCmMrZpjuZcC5Kuo7BcuVpL0nT1dky
2OF0JTr2JWfmQv7U9ivZ0KZ/tHUTckDEVfI2Fd7OkPLDx/JnhZb3YLqTKs2yAk2i
/FanwVGjvFRntq0bAAdejKMcBxybMlPzkhZhTJqqIfwJSx/IAHPkSiXPpvX154mi
zIpcwtCwbNZ9PmF3tLyiao/JHdW+HOrSOi4f/qgZGpaObeSObo7MDpAW1SaGCrW4
iA8t0JHjCP8PW972v3X5u6t3nFiiIWp4jBaGMt4Q2s17LImota/0WUNCZ9mNOoPF
jUGIG6dijCbAxUA995DkHK0X08VRtk+xxR20J1mScDEMgY6Q7yoLLrawPPuiL4gD
ChY6Tvoi3/LOpxyW0+tbO36wjLjwGX4XConG2B+bKMN5Gok/eCMWQevt1UfyHDG2
TjGBAB152exhnER8N6NXaRREx0/J9M1ea+N/kAQ5OZnTCjt7m+Iti2y2TzmIs0eQ
`protect END_PROTECTED
