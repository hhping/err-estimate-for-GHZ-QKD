`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+BINbBBu2L6mlpqypjnqIplewVxBNJxyiN5LT3a11DLI1DY9oh1T2vpssvooG1J
XucxIbb/wkpkoT4IzTByIn5PBIsU/5W4ihG5ycHemC05KwoofB2bBjJbdV9y0r6a
g6CccFv7zuUcbgHQuH1Tvm3pw4oh2n4YWgKth6izt9Hd+8dVPXCg0HxKBLCtK+R8
B/Suc5uPLghQVlrijp6dHt1URdwrEtIRuiU1dXk4puX71n6IRCPTYJMrjZxkWoMj
0jP89x1KgBWzw4cHzb3yr8KOPWYGPLCtXt7jGNd0AH00dqzXmX+gTF9OzLBywm5/
3rjnQ58a4GbJdIpddqjxa2Ub8SuN5c2LtpBTIWDanxRXd5DfiJ6bklDkDL97A0C5
KQbmQqS0GTyIdHXIvUarNc9/KQ/LR7VHEjPbVpcV5a5io0PhUQDG+8YPmFeZiwZl
n3UWvyuEbSjdRmRw4tzwUnTOgRs5KYVgcr56wxc68wp40l1kqPBoeE1tnxdsB5Du
dVRxfM/NV/fD/7lagyjAUy+FVVOtKCXyV496n+L90Log1l0b4+aCOQ3ME87u0r48
VEwIiOrstoxZZX9FQm5tb9eb2uUSEu9fC2nazI62jPLWHKeaY3NbgLIBuIJ52VF8
ZJKYt0pWuQJPt31f0GN4/+dPq/KcPaT6rQzo/pippBfWiOABOAro59oLPt5AFMRu
q3Gb4jiOFuSsn0vX0DSW3KoerkQN4QEglUZBnHmzhf0REcqK813rksOx3f1IGJ66
DNTDYAAAj6HPdGu0O/yRW0f+WKFph6xPTvZWeDpwfkp4dERfO+ozqSNpht4BG6Rn
rlkzHbwUQT5U16dlNXqDzGOF/hrm6GbxCOrGlZIwnvbJSG04PRq8eV6OaPQbh/S+
FtzPKPG4JlLJ3G1lOwD9RISjYNyH+hCYvPmOlF73xU4rgYh887G/E+E7TbrVmyou
Gbfe4HrdkmUhCSxEFqLIMU/JRfYxk9X+sOI9WgaKlhbF16iUnblbfvB/GsnuMZJB
QKa5J133iBLKch3NyFCJz9ESBkAqHJI7zi0V2tcPqNXgTMuGQXWLgYkxSDay5QHc
TBl1uGgaiiWZAllGc2UkB/DodYDrzkIoY1y24u2Rfprn3BqVp5aB/ktpVmPbWxlE
VfnupLqpUjlKeAx2Vg0oq+gO/SS0ftccg22l3E+se/0t6DdasCk5fwA28BSGoGCj
tDpGvZa0dd5fQCefKO+mKpFljEwgqXd6LZpX45O8RDuq6otd4afNn+ju1uOLhLn2
HKSUN2dPU7Sj9SPKhOP4KZij2x7Fj2TxDfWD5boFxgnWhttrpPXhedHuDy3BM64r
9p62G2yeeuYRiiz0wvzq1Q24tQbLZhg2oCag0nSr7JEcq4wwIP7ymYl26qo6wCu7
9w2Vn+noFmBLQw+ycjqDhyXvfTaSekfZJhS5p3Xj9r67Jt3zaI6weRWMpq+b7cXX
+WHIn1jecXiJdpG5Rkuskga3PBOC9HqrrWqePqtHBpAKrSWMZ7AtDqXq34XuRm4P
+/qoeDjDvRAP1NMtTf7oLHGMAm0XqUO5sq9mjPH1Fyasd/h1EaEwmiH1AGo950XQ
GsTQZNECaxl3KPrlINeN8R1agfT6x1WC6wFO8nhq1Y8Czu7lOgt729K9oAk7ZPWv
IeSn5MKESkEnx8GPK2pIfZRFYtTsEmBcmL4ylHIbFaKFEqQCFP3dfroxviB+P74F
wTmo0DKhM5sIGel0saFdAtpEWrhcXOo+HyEixyp0PFGG3YwTk4vMJheU9BnGW7cd
dHPOc+8ONrUBjH8hjKnVuFauoTin94BqXAVLmXVXNJKLsfOiwbKvpy5JCMghaPIS
PGzSQQSPAs+bOaKa5cmvFIvOUEuFBuXvqxmjzVP4g62UJu07km9+EXSbLvLWPM+A
4AEwkDWtWKHALLxj7GsTd3C1Tv4eDfXMAh//RTJJCncrJWzvgH88LSiduQzxyLWg
PXps1a+iilm1EUYTuDiItQ==
`protect END_PROTECTED
