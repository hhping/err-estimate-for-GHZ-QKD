`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAsOESKXIriF8uITVKOhDZnjphhAvc7ca5EvDEqZz3ZF269Cmswr2jUgSTrwEJ9W
ctwGKtQdi0sAL55gcC5bDk+ilA5Ajf12iyz0utRXBX8P0g93qjVtRiQN5IMF3PeO
8BNs7EEdyEUx1LJHsmFqerrPJCbtYwXHAT4aNa/dduFiA6ihOtrvgJUAoll8W9wK
C53cNlZXrLswwH/CvJZn6b0QoGftLvENTunbt3QrpeHZNVa44stj2OlIUIWT2afj
iB3xMp6zD5p1y7+bzwzuTg3lh4MDGeQEQYW65AVPeNGhF4H77YEekte0kuz0/iCt
MKZuRz5bbifsy2NCHpLsTmOMXz5di3gHHCj6i5f6L1RPGDgrqFuzf3buSxkeDNOs
tNKnfJwLWjMKQcR0GBgwcUC1Us/zk4A3MdrfvO8oCpWwj0GuvteynOP6guPk9Zio
cUIMIePdew/zFQ7NQjoEGWJwzxY3/RSrndwFF30Qhns9RVbyj5mxYlxXipAqMHm/
5Jux77PjjQNOZy7MuG687JOCr8kQoXn8pvByKefLERujLxXyWPEQw/sgow3hskM9
CWPKZKyXnHAUy2MTeCv5tIg0vxaMVD5OflfxJnZwXO5ExR4IvSUCtkWKH/zBHPBV
DfLYKW+QiZGSm41kZ+hyrEzAaSJz7HaSqzqx+HQBrX2GH0SQvqOzbih8yhZi8RMY
aE9kik2ioRaYgE9fp9zejf+J9PIomSVmgaJkKgj1ZuD5/LJ9rLrFTelqJHJGOpdZ
FBNow1DFv3dyiC/Zh84kqt5gMOtl/SNFL4HcTopxZbQDdDa2M0LnLIOJ/ooruIto
TeLGZkqZxZVqNhsu3195mT9azWBVluZ5Mo+NMadQIC96nlSWwUSXrIsgfMk07Lye
O/daomhYM4c+vgsSP7eBwCC4Ax9bfL4f95H/ez5c4kp1LAmeT6XzSDEbjUKEt8xz
vgRM98JlxSdOfsgE7uWyUQcfO7nu4hAt5r/nSGbKP6Glqm/2XySAsm5TXB9R+Wvw
LnLvhoFT27iGbaWLmeNDNyQW1C1i6w30H/qc6ze42O7MVkrtXtz3HKqZHeYQgfAY
hJcsHMAi/LohTC8NrpjCc9qTXQcoR56GPvTbH5Td+ZjOshojGNWC51J47wbTVN0O
MltTehrPmtxrhuaLkooPA5O13egCbKbFMBz9WUSQOt0eBkwuxg9uN3pqsPuTscIw
Lnq4Uv6gKpB2r7R02GGCv8Gxaq3B1rUAOANVCO+84oNhdM18k8bEENazzijJuNNg
lhVmEDjVlYUbR8UhgEyoa+FBDjrIpKr8GPZR3P58mB9kn9jFu+lTy3jQBQD62Tet
exx5IRYWXLXR84GpHnB6tfBkJi+35pvy+J2Qby8IsmeufDvWOcID0jxewXgYLL2K
+fZLyJzJE+g/tQnUtLZNhwvNOFXDLBs4Rw/Zq35U1IjLy2MzJgIOiK50xODVxu6s
8pB4gKDeofdn9riTjk9BQlf3hjP/kwrzQGcmimkj45fphw1iej4J0AZpDx+BNCKg
2cKkwWhR7BxmAUQthxkQPL8qQddI93VyGFhD4dyMmtpKAv+xUr6e5FTMPRc42jn5
vCloRzL1P1LxZnF4b1HkZibJ16k/Cg49ZRj/wbTfahQh2fu7KNJDj3FSUlt4OAl2
rfSe/5UNrRH1KXcJqmYkR4BFWy3J2I14zw1RZNRYTmrAY1L5xKY4k/pxUoiaP6mv
9/nP6GJTcp4XsMqnm31lZINjYQ1sf956iuTLa5HCXWe92JZGpFibLkKlsxVimd9R
0MaVSFZsG/qba8FXfO2y1gprgHODyPofxOoj7NjikL1/jPejQhtUUqMJWvqes0Yg
Kk+yD88cjKybTZ/+kEdSH/3DZ4lB7Vh23u5UXkOJBB+xh79F/m5Rcd+Uz80d8aIN
lCJg3uSSDaqrYwFVhE+6LlBX7jROAWhHVItoRDoIzWYxJfNJ6hXVxQP3NiNYJZqE
TBHnlahQDrZd6sye4UvbZz18nOPKt3ScpmE3KiCqu2/sYdnPrIN5KoQ9enf58Dto
OGkCe778qi5V2y/HfRJbGt0VDfAWN8wzkghWTbiY35MwxdiNkXmslq4m+tOT72hQ
ZRv5U4fXDZi4eZ13XaqQTVx1GlZwaqrVzXazcMRz7NUDb17OiEcKA+rX+vVcxl58
pQQ4q4JGyPiG89464P3tNhGiI+DtoB/5ELvZwGHpqplsf9y7UXke6O1tF9RUfcCB
pB9V+DG2g/4dIQmoJ7hQciCda6uBopIP/EmI+FFPjefsLh8/F5o4jo/H9wjsnXyd
qmSDEBfH/YG4f2988ZjDGsaJmD7D9Uzeq3byD9mdnwqgKsKQ5iZwIEGlCyDlmp1/
c4QN85F7iwQE84wc0AI91NeCEhH4FmkaGKUeMAd6LxAmrVxLuoodTCacpJwinhSs
d8KQZQ9d7aqleT1bMYCiHqaAI7BZkRBo3e39tUNKnZNYwSLK32p+KdPYQTaZkRNH
f+7N6wUHId3ysw9NS/Ulh2qeVg6U/YM7rKENoRvdTcUg8+5dYQSAqBrBdfAxW1lt
3UcCcC5xYNXnrgtTs/OrrS3iuf7X5u9iNcxcYaeUETp+8hb72wkgu3T0dPLV51+Y
JqlVDQdOTMfB8eKN426MigSlDKucClP6Pvs+9sQpYVzyEOEyfzD3Bc4FPQadz/F5
0sxZvzuipM67BdpyTez3MV5JvySZa5e1EwnAE3GZdexdXxQQhQ7W0yFyCtJSrtsF
/4c5tGINKVWPkr4hhoc6SbbYHkxzgLwhqr1QWiNu0UE0LKSN0k9WUdkf9kx5AR1x
54OygTwX9j0oijpbNYd0cXKLVu0iTDxNLKz+PFzmJuLQsVT4fvBDKSwJREof35iN
rJBWqIFxPY+rd1IjkEqgxwh7WFOvKGpE5oGBDNt6ysQ/0/tC/vzvnSMpbS8Yo/In
ts+3+0H1E/G3jcRS56Sq1To/1YiGOTWjebs5pYhDnFbhx9IJnAW/+wvcMRZEcvG5
Z2Hrc2FMaPsubDPCPufH7icmTG7rCCyUMQYmYDDnjZZuMYx8hZWKHp0FsckugYC+
fFECOzkvcRwDz7UrL9l8Zyq/BECwFHc4KuwqdZSFBgjMLUYJ7/qYLgyU8dnAhy0a
MH3QL9Am9dCt8nfrJmjU1vU3FmqtRJYa+jGqnA2f7BSKU7IzAG0jaVsJUepVeRWM
AFEnkWwocKNyAeVFv1qiH8rkS2yVTdpsRQZXhGdcML8kp67SwhSFlrN6Ffspoa1h
+IlTrKA6aGVw3LGgRQXOyDwRW/+An2rsHHUVPTOtBIzHffntYvdOJ+/QQEYZVeh7
L9GJCB3E/UJuAw6Jv+InbvLvs+ZjeHZ/j14uN5KLrOQ0sf+NXTENUZMw5k9U0S8c
4xk4sQMmdMijFuCqp4u05L72MccJsBciBHSbYlsFG5Or8gfZ1cin3rpUeiJBgY/c
VoXgWBaot5TMJOEKaNmT5ib8f1/OB/gRN1sUnagEVNHqOWl5EZs1vTu8WYI7wWr9
lor4NeU3d5iNEhfLvPTBT38ZaPftM7qxIaS/Zmc3Sxw+/Rh8VEDs8iI1I1FKn0iu
ByQg5Jo9CClHujnC0JmpJI43dXHP5fXTYssXXVcMhdIIz5IHwKagJdQFw6Vd3jIf
kjQJIVyRdRAO2OTZezHSu3klK/KVBlAd5cY5m3ZOLzE7ntO7LbUC4LQP9KqyDWsB
XTnNN6X7OSisPF8mDQvh2Sn4bmoWzvc/+rLXiKwxkXe+LQFThitZJLdpDFM2gvnp
J18eZGNyRtvyAdoZntu8hNTPOAqx0BhBpXOX7+z832KZ8RbnUwI9nPPbCxeY2UMA
eHUlW+SYc6TD5WPabRX3bLrWhH2g3N6xovoMiohU4albzgpJhSS4Hhxz1HehE5Li
ykcg6nNN1gBXoZ6LSE0JhWWviYqI9iAip+uyCDkVbQ7DCsjsY+mJsDrjeANrd1AS
EdpNwHVtpEXqii7IA3bitUfT2VTPSsQybIa+iM4j1Mk2wsVTvKt/j0pLJ5XkmpVC
ATJ3pNLy+/AGIFNjp+bKzV4uN6fds84S4Czd89DWcTHcm37516FsMm8l9xGV5CzR
YsNFQmElLxC2C5U5XhSB+mwebfvyXNv9vvSoWRRyYEHL8msqcpEsIKSFZ//Z5R7t
Z3p1LqzrSwyDCGEMNSiTp+yZ/tuhv9tuAVzVKAQ+9a2fNwD/k9jbbR/lx1S7tPSW
tyebAAjmjMyYimHsmVoMB23C2xOEo4BpKu4XLt6UM/JXT+FWISuf6Nm6Kyviv3zj
gCT/BRlT8D3NkJcmb9mTvBoy0fCjKOiFaf/2deIR+UpVaVk/2ZCSecxx14ahhwox
6FVEAIvJPvjR0TMWYHCleduUZ/PYLnEtvYKcLtV+L3m46MpFpczbjlzk6vaLavaf
5c20Q6ZycvEDQz+CLzOH3aFHYYR1VtB2qmJl1cDr6vNRaWrxscdyx/+ambZxJEGE
zg9vb4hi80GnOHFAJg0+sitSw4mgh5iqWfxkw2HXDLMBrZCxa9vePSHuEf3Wlmtf
iCmWBACXsCc/UqBWG+K9PLCL2DNvkKS3EC/btl/R0R6OOIh/N8HrUTkATx8OV31K
aG9WhhxgaBLnVj5RLj9FV6bxDhkNE/TSRlj3wdtOw6+48ylWS3lpClEtc+82ddEV
X/D9NNOkRidpoavy030O2vt5C2rIQMZLO2tQt+L+LSi5vk1z32NZHJPSzFSApSdb
2fbGTH52yaOgrUXoTZSUk7I7cR7L/B5oP6IU9gIpikRAFkojG0rWuXVV6iJrRoZs
p/+bWJkr4ROOGl0AODniKzHVy+8v6xVBY+4pcQgK1+KSymvIHEq64yjCOowktMh7
O0E3Ig2QgOhaLhrSgoZS0x9i0C4hYq3ZOaaBerhZhpJBG/5KKMckZaoK24nAq+Ro
7nwLIKWTVwSz4MNAsm0u3U/qe5YEyYlPwZ9buNs7YIX5bfgU47R5h+hUVYie/6Kd
JSd+7mAlfaxBD8sqKBjJ+on6kceJtf4FKA/aPvkOfa7g5zhGz1El4v+rLtozxxAs
xCpygOhuUP/YBf8uRrpiqALIueqVxI+DomPGsBRekgPO+rkszH9aAV+5kWHjo9kv
ouH7OhgJxhRCTHaGpTqcEyB1aNP81FQ2u8M84d9EjJFsiDoFvZD6hpNlPSKVg8AQ
KbxBktrZMoOhWiWHI0vYrBjhsHdOSK7pnGg/jQcwRZV8q+Y27oz7DMtuTOM5xK5W
uU8hoD1EuBkGMS1FSMVe1IXsKfLLQs7imBq4AKPVB9DdKHA5eroLfs+7iyIxHJ4U
HNOxVKF/H/mKEBBFnblP0y8BsxI0/blU59ABKYQMVmkbWAiC6TVMpBtIooCI2sGT
YNWOwMQ0YGmLTUhlq0IMrYTbJTxTQStAawSkHopFXvq5B2Z0Q8sKAxIR8Lmo05Be
gCtraguGlf+PPaptSLhZxgap3ZdWkox38fD0kaz462V66mp5oKEv99kcDU6Wp/yW
EWt8kz+1jmSCZecIDRsOtU50IyUpf1bOOkVgTO4o0S45TMiwuPUJLXdpFhHyF4eA
8I7Z4bpJ1YOpTVyETw4JXRMSJBs8LmIOk9ZTvjnl9RZK0GNkvfMr5eVTd7OK6XoH
UwMUIGi5LCWz4q7dUyBbPIJQ1XnkZuqOg7Ycmx0krmYuYFQ1NsijwmFa5OJqMq2M
0ywjAMgdhZbdL0eXvewSGgKv+0IFqn5UrC9TW+Wwn9/fRl8+PwUTMItmuqhSe7LQ
wgXPbnmjiLhGRaSu+ViDCDFNYSitzF7TTfizXj7Yb1/+Yk8UPaXOuZ3ob/113zkX
JZmjM3At5amLDS5T15BroVWO6qpVwtZxHOlvscrQkC9qfJ7gjebjJQbJKmWbfF0J
7HBK5h3JbBxCw70YVRu1l0M9/MCjO6BbhbiJdMteqE70/PIrHHPMD0Z9E9VPcM3T
iLWSBS9v1PMKTNPDg+VFcALGSL96C5hJh6BXt/0WFQWYHeArzAyCKMsqhBtg1CnY
gMW/qQJILnAyCWrrTJduAgh686itqELs09GVLhAU6NpjgVKJ6ykNYSWyHOOE2Pio
coP+/wfWz8XzcEEfPPfyngoF8n6jriMFQ0vYEV+wiEHJSNvCVmxLuDPVqrUj29jH
pwt1/3koa3JvPb229hcqbevSNCbqh5Gpp2P67Xos3RsgcQ5eBXFpsLQP7HSUj7kn
iKNMNQ5xSy4CzCJndT7jeNFjLARLh2XPixPRH374DjeFtBVLG/oP+dfD5XnFFUY+
OMDOlmIiFlk/ilPdfnDlThUfPAzEpYsmi0hbl0pMOKBOLesCEMkM59tk76GuhNmY
1KdOkiLlP/pTDoVjWYF7z28Z92ib1oUKxic6sqUrb4yJMygV09wCgTZodmH/uDs2
gfKynqID3A4/O9OfPLV2XD0B0aMP8uPKdIYRLuP4UtiYUKivh+uoFXBnhew1mAOq
IUyfr3mmLi8XN6hHxwmCwfht1E0GMTGW8HRWNmUhcmdUV/4Kv1/K40gnGvGy25RM
lOzMkXhelX+NwcCOc6HxVc6Vm9pfGX+IDquoUMUvCaaPapeegcf9B/VC6uida8p3
bhnvHOvlOAVVzjl/INjyX826fjW/cmA1n/pELkeVhzdmvlJ0i2oBJXvoapRRiRPK
GGOyaFXoOLfZ4GANx7qZmM2CGWQfrg18xpJLMI1iZA+vimjO4iHmLIwDfaKHbNS1
/boNoVERNcX1qFS9bHHWLf4xUKVlMFnmqRXrsp4i0hmAiDc7H+KZIa0MWg2YW+Fp
5yArL0g3hv2Zk/+1GD7hV+eBgsSBlq5pCUbApzGYcB9GPVGp161YbfGEZCVrJ2nC
DVxa+FlnKOFz2PThjxjy49KwygPe4tXkCyryO8M16qXkQFVVneCkXQshZS4tW0kD
VZLOHHKWhLOoOysNkJ2cYC7VKEs6/k5uyGu3EKBJndMaC1Lv/dc95z50LtKk3FBE
yQtvieJnSkSR+9R8RIwsNxxgHwGKmJ7lzgbSLdyhdnYLRG3rCAKqmkIX/csasz3b
lXuuYtDrgj90kRXGi+PQpmoYdsFGNJgSz4BBpzF97RmUb9JTNH0NPAZ6g+c3Omed
j3IOmXQx81pd/l231aoqj0yTONcPTwiQN9he4BG5IgSxDxm8LzwSINpCmoXW5mNK
HArtYYSHR2y21QksJfo5RPNikqwsMOeFpO6rVeDexLQge7T6/G5zNAQW/Q/J/oww
is5tCvNc7V2KSDCOeHycQz1waquZ07DULT2Ita3oQodh9b17ch4gBYWM1uYcBE2b
vVkvQUR12tzhgvt8cmwWckJS6ek9GgINT4vFR19JejyVswVQUs3rnXxU8tYJ++E9
iZYOP4AvSfhhnq40tvgFXO5FjYOLJpjZZeqJXuIKF1A5F7N6gSs3mq1shuMZTMS/
vmqUq7o5tPieq+Kqg7SlA71O9Po7t5JN3TcnJwyS72v+ctxfP3O9aLDHuwXZGiP9
bzX/0D3Q5yVDCDgcbk5fLcfaD/Cv7JaTPPC5TlBfoBwNmwlAt9Z0VMv/33LGp8FC
G1FmPq+C8i6Qyf5C67azVNoT0H0QSbUsGqiYiK9Gz9SwvTJtxervYVJQJtUCjkjA
IpVKrA2ASJlcg+d+GTGwmEIBHPXEOdknU4JxPBeARpnJqcsP4wcC03L/IMa7mfIg
N4A4rjyyJgVGezX5Qd0n0FaCgXnKLGJ6lF95We5+HOmrMqXxN7Ru1LpTTn0bgJVM
6wRr7T9rsU5WWCjYyLRt6vKSLQVUcuGdw2cg9vIM5Ma3/luLdbXN2a0KNHGr4Qv5
rwwYMEmffuW9fKAzGvPpn/ulshLDYB9sz+x5gCRjgGGywbhlz2FwgpNepCr9L8uR
x6AUGzNSyqn+BBOtWJ1ZStpZh3Qr7mPE8p8+HA3l7IJI9tnRqj+0HWKOUPGu8ml2
d1AZVNMhnNSZjquv6jU53oggqo+FYCDeU0awXTeyHelyInnOs4dgdDH5mqweKshv
FLXSpVwlIoxWS+6jHbY4mGz2/zyisa1y8SqjXdf4glmgClSTTtNj9eQROYEW8iFI
xcCkHVc0X6iGsMVBp49BM861JBOeBbWE1mP7MTm0GYSzVpc/Y+M5X16sxOC4sjCW
GhsPMmg3aKZX2r1mNEP3ns9wBmG/I4CCgh7ChQrLc1+eabMfS2Rz1BpbyQe9VTmh
Vat6xlyO9ieudhITLSostXikjIinq8M7CJ/lqxhQa+4JNXSarOTnoaB6n9F+mt7o
r5BAiJBMx9wA8uysowwslhjyJOXPrXcuMJgn6pK5JySJRZkQ6QumpnS0qwLf0AWm
tq3Zm7oHTZytLSBxMLrKNJ4U1yxPT+yf6DvOnYFsjFDyFFnZt8iFVzJ+01ilZFd0
O9pBPsOP+J2W8ZZliv2zPCw592cDSUGblmWXDxE7QTfIs39jQXFCntCB8ZOtPJlI
k21rvT29VetWJ+A0zNUIB3UvVQ0QfBfMoHyfrqwgUE7c2QdPugZgH0HodTEcgdPR
EaD1Wqw0mBZE1w4EsFwpYFzzyCGYXJIostF6C00Q7Z8VMznUZ5S9VBFDFnymijOO
P5YEV9ppbTWwemlWGQ3RroaYgEMPeQ/arBYCR16wskPT6VoGY4YkOJix67yATQbJ
un3tuB+NqYhtqDDd6vuPFj6pIk+ROQuti0w2NwGxW7/qXir6mHUd3eVISS2/fN1/
JZ4PGeyzNb+vlTblw0jZkrLf4kldNIGCiDeVXVImC5XsKoiGIFNNaK2zu4OcUCcV
/Nhq5yOLNCrWCrCUf1mD2cudR/9zJjpNqB/ZPEzC0rPOntQLUusr/BUdOws0gabe
wNlgAa7LmaP5kR20rMUoke5rIlBknrQevUCZxn/RRhElZ5/hNFWO1kR+KdjzKmdc
YX2L1lLGmkJ7PwHtbdX6+slKfDXPczgjBd9qGl53aAJ5GYItbM7OEX6/oDNpnE5M
MFeYk5HHt7k4GauWwZ7GQJdloMwoH8ayv7Qm/oDHvMRlnmnRgOeFOSOSA4xag2tw
nnbbzTmgRn3SL1znm0eaGFWAgufNLbZsec/4UblWuYy0w6SxRt7FRY3HSRaBll8d
VTzd4pwxChAQeSOvOvibucjQbwfTEC3k8Xo6axlYkl9tVQiLKOQ2zSBHJAgp2gm2
PqU4LvWabrcQnQAf1dG4f/HuX9XtwoXrjO91ENaMIjxkBWr4JuTowPkz1Sq1tLOs
6qb4nu3dOJq7ranuA6GjkXep6lgNfFis31ydML+2+NxsbAHpXQbK/8raAA9RT0TB
VXIfv9p9y76BTISfiHlNbB0qTSbCtD03eUVDVzbw02cngg/68KF1al/RDtZDBP00
PpuSmwep3HlzcNkaqZj5SG5gir23370C33TvWTzSa9MPOUQfbQTw6ED6W/q5+fnn
iIca02ygaOnLGq6Z4oCnf9bQyXkn4Y1tRq26HZcbJJ+9qrM4+04gW6Tffk/ejpKi
FF+PmGfHI8vqVtiHs9UuLWE3WT5YRpEn1evI9XdigazUxspSzNAOhVWV3gMCMos1
bOVukIII/KxrtIlZtWLLvYF/t48oTLpn4OG+yfkdz5AsSWv0a4sr1Glid/iHpy2y
yU0qi4HUuUWfx47vywpBOHrFizheVgqsONlZDZaXZLMxHT0i4fEG+YU7mT/I/aTq
pxA/EvNWoUAVMRg5pNo9YTNnlaDPAyv0QWKY7h+rPhktqYba3NZh7nHBUaVY1L0y
Y9aJLqhiuvOV8HPLcdJ7X1O3KfbDjAjA7g3UKSwHQM2TuJRSuuCu9KrJou0Y5QEU
SH6VvGzrP1yEtamyxvOcfa7Pf/PhQqu3003jo1Z0ho7kqNFWdCPwxXexaxBDCcgF
WoE6nmPHMh5hnR38qokNAxd1vkatF+AKVZIM7nLfFiT/3Rz2/h9Q+R6gq4XexH3B
8Kx3IN/9vV2v9VNpVPFSHMkRPIipIPr9gQwcnudbR8OXjeOlFQLauHR6cFQloQJw
WlxOmnNQ4yadfwA9u7RNgal8AyXsuVnrKgdi7PRVwwd0K03Ira96TOfCS+6+XMFy
iW8dNBRSR+G3pMllSp/xGppBu1TdzKC8x/pU1eTBVpV1aUZ3zXG3pq6OEcAI3jmR
BsUYm5opTUgtiI8vrSx81Kubxw5oJ2QGlIvPAW0vJFCRJ8BqRk1jPWKwNgkOKgt9
Rt7PVAA0UYHXF/ky6bq8rvPdbyc9jhsxL8ylpL6eXljKItYdrrh8aeeMv9fWP1Dm
ExXXKeWomZPSRjoumhABH5lkuvXKOrGZIM+fWW0zvzTyFf3y9liMf5N2tPQ3JzUH
P9pFYBZc5xi1weaabEcpyJ+LA/GQCfaDDnN7r5e94hejLPupvmPviumXd8TMlrqs
XwsYj4AGZHWdmJyga9SSxXfz7eUl1HkZk4zIN2u1TP+LTnzuKZ6t/4P0WyIxUoCe
jcyBAMdGYLXXteUCiYVlA/ZMcp5gCTFZgjMwy2zKqnfqK/qINQZrj85FNfC4z1eE
hg8TuUWWGp83Wc/+BZJLr39U0VK66m3BK33XS5MzzaJurDJGToiglH7oDlI1u+Mq
Dqu4OE07KHsFInsK94/N17NP0kES39IQ5udZXbM68TTWhnch2bXc+VIYMek6m8NQ
KaiO8r7dI/OH61p42md3cPcVg1CqbzKWdRsO8zFzj4118Dqcj022UueZP/SYPx4K
wXXd94jZRgwI6SK5drT15Ku97jULNMuyN6+CeKu1T/RqYHnm4ffkLDRVrVPhgSFr
iJxw9FhTxyj2qLtRmCe14yIoMALzVHndc9ggkHrwjgylZkbM6BHZTvgtIJkcI0K1
/xF1qxcJ9ilEjorXpfR3k21w/NQIZGdkmCCQYa9GYMMyk6qe1fHA9qZmBHV5Hphk
kI8spCOEvb1UBDvH9UUcNEAI7Ln1lqYxqZQcw0vD87K/Hf7lIRA8IugnYf56bg3W
5UJghx7sSO2FKF1U0Lq8NwFWokxvyjYqgupnygK1R5ykPtyLSCBFmJ/S3msLiW3W
rJVf9KCG40xu8+0HymNTs6bGnCzH15tB70XZwgXl5f0PA+tF6wvsmI9CnOeo/5Wb
HAQNYVJ6LpxJOJQbEcxhtjnF0q7xDAHtNlTdAw+npxFvxTBPQ9dExBhVTSY3OqhV
qcfyu77BbffVkbCA8YBqKWqjQAqIV+3wVBtAj1Ky3SJ2XnhHPkDU4k01c0HDuYjc
xzPqSWLGC64ABOiMMXh2CDMwIIcRibcj9vdbOrnT14RZj+IXHMniaFbpbIRB8egI
1zdhgZ3aKZurCupAlr5uOZmlPgAUdlFxodBWD11aMiMrD+PJEf9lDpHJOwghjEWP
Hors2eSn9LAWxs3f3mVEWZxvu4zqnMCTBxY5Q7FmMrja3Gv0gK/koR7yPbxVxSmH
68JRKBV4tSILvQo7HnMCGDUleUi8sIT/2D72AGfjfALcv0NljTEHOiDqfcNZ8lj9
TY3YUkCQ1iYd1ulpv/qhtqapevnFKGg7E8ZSRvDzhCbYVXi9k6mN+4+P6cpSwtB+
tn5V32ZctTqO4jMgPGwto2SpvOGCBKRcG82fkDWW2Acztb1nKGFhVqsO50zXJft4
8e6KuZvITKFl7tvAvjguU5F0xG2ZiwQ9rNdQGaO9xsIXCxyTPRoPMUbZXU8zJKOQ
Cqyg79ps5Opge9Owc8l5yil3GWffXjUt7Y4LWPV185+R/WTBpYxkCDxRfojAiztC
ERQh61mwonk876zxt2xLh4JG8XntjVFMVZnQ4dy+Ae/jOVvLrF34STNCBsWMG+jH
ESfn0nhPjKj7SHjJVriJEopl3IO34rWfQORxyskLT8BAzXMbE01UsBb90cuu3CEo
gPM6Fa0lMjPM4GvpTUuNKFItNjLJBnZQxaAT92cUdrZk4YqWbuS2SQp+a8k3qWOw
XoXMRPS5H3i1yV9yw380eXzGoRGOWMFY+fKBVocUyw8JorbfAQF30jAYWjjXkImo
QlTndMlaP55KIk6b2NjB9q4vHGfP0k+FBCY2SgKFSQPMPV0BwDfhp/sh7qk4muzk
kok5ujkpkYjmYTpNEN/MGRnkafYixRIM9gjfVcBQ+0CtFKyLfu2mfe+vyUmPXAHC
MxZf+UCEfgrKoe0uCVHSRSaL/xHhQfy+fDWvHYXhEDv3ZZ8Dt/QsreEHWPQFS7zJ
GL332VtMweGW3l3wNZsl42222OAHL1zLnsPYnoTh4RjrqYAZkKbUNnVS5wGJaHVd
6/zHJLz06KsExkDsiaEtmg0ZFnPDCUT0oy4GD2IlljWZA94DWUuZKGqGC5J9Hi7J
Wmsn1U3gLbF8WwEdl0h2BCJC19EzNaVGXDufHELHP/6YCprGSXVEYC05aGwY8bZi
E7F8uW+X9JINaehqZu2p/g4A5b7ROihhG/nsaQGPQoGHVM6/yi5bLtqivKziDfA9
0qvSj/mNYaXHUfvYj8I8z4fiMzUN5+RNDFHDQx2ZGQnETujEUjiOUJAnZUH6jcKv
OKDSaRq9qjxm3ZNd0zrY0B4KB2OaSKGxlFPM1wGgWDaqxzgwg0wvSNgWKWQK3w47
q3WPEzeqFbsVHnieyijypUulq7i+eXduoiyFJtW1k+EQTTFdg7u6ubUJXXeZ1vk/
+7Zf4O0G/A+u9xc49+MlO/P2hu3atFa2Wtje6sAnZqvPicUOA11jP/W5XMJWB3mO
pyx/Db9PUgtsgRDCJx0AWRg3Qnr9a0euYo8XNsrWzBDcZxzS0YazkR0ORnc3wq1J
uHzPBJ7MzcM8lzhEVjfifHDA5CIE82rWNFzMdHhELoGyZc6OCkbISm3xuRb41pIw
1j+SJlcZVmLgtZSlD63KwkAHbEMAs5eEmzdzIc0rjBvStsfTx3FEKnk9PdCyiuuc
CUIvaB6e4HjBXUCovYC9iL/v5D857QWIH7e0jl9FRM7l27PpbVY+YL68JOaE+Lrc
sGpC/U+od4hsnt/pQUChLIo/JMaPjMZZDcLgm+iVAHH+uEsEiGqDDRw+kqS/p86u
5g9nVlpuEbqLi6m3rCaH6LQuWO8lBzj5uJ715qGOmag=
`protect END_PROTECTED
