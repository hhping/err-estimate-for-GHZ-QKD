`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjPT8HFiBguI46QelwwZ3oVg4K2xV4XoJjvsz7BTMG3H3VhbvNjy/q8ZCBtLS9ZI
f7GwsxoXkaTWlO8CGo5nwevqxzmYsCvKGWSfHtypwjxhJqeIqV3TP1oBoTT4TckF
xY7+fNzoKEsO5NeySJoWnnR3LUU5RANzBU/sq1QxKvug9pvdMokm6xtqyGOMxnM+
RZnkVc4OAbZn04AuiBmzqnNiAT34K0G3jzGLFLbYsJJBpkqLbugf5II08MaqHgqk
H/9HPY6KSBO0SiVPXy0TjPC4iwd4tKWNElD93MFQsDsHK+Kup4y+z8s0HvebIw+3
Zy8QYCRFWsgDvM1hac8X0rW4hWMbkMwKXBaBBuFNoQQ6I3Papf6N8YDau4dbXDsA
Gl+pXOgj4umWDcAeJXwHe4yghVYMKqOU2KrjHTFkSX9OFSguR6LOAVyu4x5E8Ctg
prDfaCHbSoVwfO+gEj4TmNxQxfNKK+eRIOJGP7wsL3M=
`protect END_PROTECTED
