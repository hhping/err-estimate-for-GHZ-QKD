`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asiUgqYu4hFy7NBHaVbZhdzW7A0SoKr+FURZB+EaciT20d0h+QeypOfcwv5Zdsn0
rO/K3+w/mjaD5GK8MgNgQ1/M2iYqgVXASSUlVQnnQdiQJDFRMUA0Q2WJScI83l42
WwVYw1aw0SiS0vuJjdR7i3Oc1e03LneMSna2TfWp25FVZTX59DXGpitcg26DxFPW
5Azpab96wDQujrQTS6rG1hmmZgQpv5XEo5DSuXlMzjnJnz5CFAhFyBwi0eNUiZ13
Nr7xmY32eUamk2hprF2YP8N8YRjx4G7tber5u7+5NumH6LtFIqHmuTkFW09s6uU/
COBbxUIZipYXqTunv/MsJaA3QVA1qHQt76swW51iyQoXxkP4rRwUD3eqsxsdTCZO
6jApFNOEA5TdQsVN80W5Pg6HmtgbuzohyWOaco798uoS/3qCWGrgX0rcWysoi1Nl
h5bvdk/aznIGszdjVXoffcJfg+alxDm/x/kX4hnosdSRSAs5KgrIEGFP4N4QGpGj
IOqlLK7+X9lZA/RAYnF6590zrrGw1LFPuqvegt5z3jkvOj5s29S+QYBaVgdZMOgZ
a0HJVVDNY0srT5XtK9QM0w3yrCE7N1zLhge3xrI8TO7cFc70rgTP2DbfR98wWVhj
m6seJ/xZ4y6IwC7a/g4KaOVXjdyXbqQQKrkJ/jCYP0vW62up5TyS32+TpPFMrfnG
usLr4GQ5g33Ihu2qxYTfFjO6HkLg7tEJavNVjo/NU3I6XqBoP3tOknYn4HImcAuo
DzDpBOwRUK6ekiedMgDpv2t23qvlcfMZcTnj3CI4ShnQh2j1rw+OJIqYH9Uay9MY
PiNNIdPBiL6/yh6cu/zQzPueu8tKK9r1gkTmltTcXcd3GQxbYIvy74V8KhE2NwMI
QeXIoTjG3kiNRjV6q5tVWW/GBk373xnKWN1Ux8HvFLTa/FfWbnsxoJY2br774VWX
Vs2t2uvLTO9rxBtoWpi5iby4hgsgPGRjTnmhQ01QsJbL0n7Y5pXswUF6oX3DE8+s
m9h3TMQbjrHGzNHC1s0gFZQAhATdxt+53ztgbJHoyvN6ealiqVDVY3U2QTVttury
YJ9mrJddDWdRVYKzFMz3VYKVVruBC52o9FNKrNxQeh2FECHZUf2fg+IfMgHqueck
zctTPd19uJhlSsZoT9kiGzammZFnKykAza9GW+47Z0rONPkmks4IST+c1F5rydwA
jvUm1YkSPk6lAY9uc0H+uFjrafcEsmMwwlhXxYjbswTbYrZJjjxELRNICQGrvSoE
B0YiCvlQY5qaMMJ9O4BQ6xUWqUEPgr8QfM85H39oJXOxC0l0xUWIK96SSC19umja
ri+w71jJ5FKgd4NQ1De1UZrOd9aGyz1rfN8mL8w04WI4Uutb4s1Ld549v9GI781m
4QicN/U3fIWm0MgiwBYaGkPjvl6jrvgvHfjml6K8CxeZUOfbxYB6oOHhCUDh4Mxo
z0pODjbXor3IHRnqWnTUmOYlywOsPvI9olLAKAqQXgbtv1q0cnxCOEVGaeY1iLz+
LQNlaTczT04ce/ZtVE9rpJy4goeoQA/fj2uvEXPH3oAikSwO30eQC/VBvEokTH/A
XHjSCzrfHPj7/WvZzcy+Fbfi19VC4asrSf5zbiei0TAPleYuzAB6ec8bs4Hux6ff
5llQ6YjOH9oBh10alaw/2iSzUbMOIYV6HDI5ATsfmZt/ahi9N27uudwNA+LjrBE5
e8ii92209ZFIedfXpQJVaVCZJXUcIEBKAScBRB/H9DB1pPpgeOZRzwksK+4K9wQb
NFuNBE19Xlqfj+wTwXaxfZRxMPjVBqdxY4VkgcxFCPKg9hoKZW3bBTogdYf5Nayu
x7gsN7A72meW2RZ9//TUZ6aRoCUTAJlvrNgXr25isftCSDwV5xXv9puuaIhNVGkb
GgoyKxOX144rBmIFT8nTf161lNKSiJZCODDZJuQ+l4BXpjtMfXWxE1CSgQYy4hk3
YPBs2xblWKMQYgjSPqofzKVJbc4ZHM8Rng9nVWEZNxGdqeKalvSGiReVIDtIDPEL
O/NDEoM4CRBy8iTRTB/X0i+eEySylmwONMJyVlU2EGJgkr5C5pMpGwNWt7IGDx5a
qv1rqJfQzHHig1LegWQ61a46vjZdBeILOeQh1zP0KFd8TfxYgA/gt35XJw5KLBBW
HCLcIfv+oaDHqXke3wtqT9UEZKFfKzoc6N5s74pF5b60B4FApRhPL7KM76EwVAJR
zvzqj0PnGE6PYdfALOpt/Mjx73QU0/Y4fwTPDvaOrDBj8bhzgFC7RR36WNBW1RnR
ZrVq4bLlVWMuTT0UeX8SgxULNMuSz4IhwLwl3qYrY7l0Ac9D1rJmm9Aj6pdzw+sb
Nm2R++nXGfmoWE2szns0vt3g4PbnS6Vxe4sH1mEtIyJ9cPERkoIHi8Jz7rUC3Vsi
NtRosedzVxjHQpv8mIT3VZZPvghNNO56ucg92WlDisU=
`protect END_PROTECTED
