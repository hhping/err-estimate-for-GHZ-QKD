`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNJFcI6JDLlqZEwfMrGFlSF9lbyM+Wenmwy/021RdYjtCPi/vRNczX2t//5JSC60
CpBC9t4nGLvdpu4MqKulJLlzjNxCwNd7w7fN1GMb8LmOdyjrRrqajw1Mh2d7UpUu
W9cUcIO9IqZoZY3NvP3d6t7b/aSdGh2yvshvkzfF4nljTxEYH5oMAG+Yu0A1xG7z
JR/7ZQWXr4UdlVU+uKxo27mDhBJZ5iMd5xZEibEnUxTdKS19Woh1oJrp2aWCrHbC
M7oL84Hbr3HXrdc+4SBVhWzPK9sV/hjUixmCp1zg0iohddqUJsv4U4HI7CD5Klph
lVA0g1o/OG9BKauTQ30MoVme4kWZUHydrpM2YfJ82M4321UbK/hEKlEMOIYdTbhc
mhhUuLzuBE/cSBPcvK5BYNv0RcM7XAM3z61LtPLFA7fORph2l8Rto9PPlBldVrvP
gv4+CnAm14W4uEG4AcGq1E3M1p6vCY0aYgGhEU4Wp0itsSzRbfDYFkJfhDdcIgem
PoRg9eWqHDgZJpj2EPpknc+kxOzWaJ+/CBcWLyANILzGbPFOSQRdoNUsczsRfFGw
+s0lglWPP8OgLgLkYIsrY+nzV0sCmXGgXb+F/OzAyyDqgq2jCmNDSeMbDoS+PNfG
e3ajlR+y/RVaVWt77opbZ5ypDYtsNmuBtPeEMxM4baWUcKyDg5184A/7oRiCDiEt
/pf7HtZrplCcypTEFnhxxpJIah2HgNav1KYCLXZ/XKhL7oTDwAXkfbQChjL09JKY
te2AWf72sceI0slX1za623OQ8LfaZeod0TCosGX+o3EEBJFpeW7/d+ft4OlzqGsz
Ur3Z7VywHSiBRiIcHKle8ZVnOJmWyl0X0ltvG43/iuZlkmPaHQPzUq8+LtSZGcxU
3FRIld4mKw/u1Cr6YhtzuYFRClaZAfuYnrw5IpGeYsaXwUWiH31juUalBK1v5N/i
4b60EwN3R6BqpXSu2c7t2ms3v6Y8SgC/O30FEJUoLOlybNkEIG8HYabiYpil/yH5
M8NGzy476UiZnf4rVm7HpfTIW8Y/tJgn1eljLMR5fW4ovf3BNqNn1apB3/vhmrAn
rRcbvtkiA7ZxE7p4+FlqQv9s/lQjXyBYqL8aP29TUh6dOhr2lUSYh09ctX3/884Q
4t4SVupq7QQaexGw/kEqaQdcl8f7jtagh9/ejFNawUZzQF8wLjT+Wsg8Gj6LKv2y
kljsu576FgT38AIJ5w2Lk5yJGZnTwPMKAXXXOddEylJ0n2HrL+eDueCfNrj5QjIQ
Aa/J1wobl2J2GI37tG2LeaI68Ej8QtocO7iTYQfD/rE0F9yOq40zGzknawivbFyx
jR/SY579Mehsof4nREaRmJ1V+DjmPE9pEcGUQwQ0szq/kXg6c4YyZgRkaP6Q+VSv
nRY9MZsgLMEHoEuRqRLTfbVHBvlg39xKKirVlbVmr1FC+92/HwNQE2iqfUpWIV5j
o5/UbYZ9VhG3/122jFIHOoKAMRX7SltNTUgO9dTnpWjbpC+Iim6XJ1TLHUE9QBrX
vNKciKvyfa1cZOQ1tmib9Os/M/oXusutGS7v2df75dar5VZeAvILG0giRyDgl5Yq
Q1/dmvUUBJRrlYu9ZlXRidHTIxjGEEHK+LxCjT9DjSqlrq8NyOtjn24/aDEn5c5M
IyJcqk7U6rw3PToD5Gb0fGilp2SE20bOpLOXRbbdRkSF72Xl52Ozzhwekq4m1gmH
EdkdeClndktad5GFfkU5p/myeOOMgy0GRlIDtsBc2ohh2f+gEK3WeTz+bTmbK8G3
mN1qHHP05/Mduzro0rHLo63HiNu3sbMLb2976xDQHWGlF1MpXkPe4iygEidu/btT
TmKDsLWxUz+R6odkbtata2ShFTUTZAKLrJ+JbybbZvIeVxGuT6VG4oZkOpRqOmIK
FCG1P4kX5L2DLwLWppPFNOAfVqQRjEPQl96hjsWuxWnre7XuAJ3TQhRl7bfwfjRs
OEm1aQ4RHoZL6PzGWwKE2KWqiMnqpjlwe1b6H54bia+y4Wo5vq5NNctD6PCOp6SB
6KizkNAmRQUThUx16bfMk1IYBaqqDAl0llXBKQun1/NrBuQ7HLBnI2zUMkE0Qt4H
+/qwjpzZiMBPBy+cyuDPWoky+cuYlE33mwbfAiwelRhKS1EuuAii++MYXm5rUDTu
sxpCZNsTNr/CwL/Z1ven8o/9oFZugfNIuQWdDvSZC5VLSHLvCDu5jkss96AT8RRJ
sNzKGJoMg16/EHP99PQMSI1hKKO13JLJJi30U4Y5UNr9ZXfDrzDylPKeZ5wC8Urp
qct4fqs9Tt3NSCCyKRXjE3QAhkzI9DXTG8JiZCqurWmEn0IHILsuKS46DDQaevsy
SaS/TUwOhDZ2ZqfjmnCudob/IN17X4a4epB3uZa7GQPhiWPvz9xk215ytlp1LLyW
1npnIv41VZWl9UU0ieKjML4Xyy8J+192/l5Tehp98hKgd0PYKXsVUi54mDuPONqV
yCUwTp9TVOXsV18Vk44ikeS0lGzDq/B9fbXUEphoBxacVwrG5rdxPJhScTuWh48k
itY/HnLQwSYDdvyYknLXFHBRTIGrtcVdkLUXnfey3wrnXZCfnuorEbcRnMrZo12T
7imdwJ4dpMTy9A32SnbPYUsoDqrLQRhSNidK2a7g+GbvFSGR3KJ8vXI4NsNUn2ig
4EjzIwXwZUJO21f+N7+Mzo0mChTj0vqCvMmTBJpwKjNzmjouXUJHUAjtZsvFcxSr
LfzsKRYgi95yp4x28GaOUkree1eKGZeYWceZqJMIaqnhugeSjNwqJRwXRtuHpZEc
s5gUo6Oihr1KoEVUtJTNrVjXNfsIzBXDJv4bMuRjDzUZMUIODW0NKLc7Ka7xY3z4
zHhsFQ7G8ykxuyR8ooL8x/st9vyl7lrcR7DJ71OrNHzqIpYQWsE95gCDW+VIuDWp
+X+pzkicnLTnIlN23xEif8KcK7DqeItEpulNXYpROx9bhZCwc29X9kcJIL1a/7W3
pHBa9KM4QM3jdNxOQkWQgavIcUqGOWskPaKSLW8yrQ3esoRQd+5udw+zzqsl8g+B
U2bjPzdPsdTBbzf6h6vo9zePIxrveJaXk4flvn2/+TkksmOnIejlfE86D8hvlk/l
2ZFUJ0QMmHL00wjf6+lYPpr7MQPHDFKlV6E4kijX7w9TNas35tpRSP/NXarV6UdS
F4j4RPpenqRGzeLsMp3F8AJoP6AnTEJu7XEvFveuBd8WtddJmxNVqglzCbZsy2TJ
h7swdaBpdEtJd5k1fwqoK+Uhg0LWC7iEyLBaqTY3ItdmljFL8mJFU47UtQKd4QE+
meK9z66HRt9e0hiMI0Ea17HMVsocZZ4GNnPNVLJc5WHjtakHyeFgZCRHRvo3d2l8
szAxgbss+Gctrar712evdX0NaeTTeQ7K1bpm6XIT5gD38299tg80DT+Wh4Tr5d+p
TiPt9R+vObTlyvEH0J/NTOR4z2eK95cyGq7dqxVfhfnip+BFfRoMUJqkVmyAj11Q
fkYohERbdaaofS+Parl5nJiMkk2499f/gGx9HLeijF+kyobc+6OEBvj5Q9i1ltRV
/71YPcFKmfB1utfzrmWOTc7tP/bFnaYkFjhiPCLRsQ8+/OJWqsVnahcInWyJTJW6
57cTfBXmdRF0/P1+BpWs/d45MmcxGoR0P4X6XqWZHadJxebz2n2zi9B7Wrk9uUCw
yLTBm30aSyZWaZ2Y5OOgRoxZOQrgAXSf084axB7P1WOTnOavmZq+C0NB7NYfhjeF
pcBAJFSb2q/y4TxzddD3/pIlL7P6IT1GWkT42CV2/SDKuh/oeZ2r+tkq8neQpZzo
3OmriuU969RkfceJNQb8nV3hGHplSOQxdyUQ4uhXklpPO7mgI3uKxDEnVGVQR6Qh
RAj40BwbDnqJ3IbNcoJ4FCA7RvIv2j4ntTFXSohQxqg+5q3bB3J2NVeovDN1/QNJ
Io1/rp9oOm0ZRESX7kVRdK+mu6+aXcveM/1x9AVtHN4aEa/6qs0k1yj+OPby/yF+
sJXXAVe4s96Id2vZJD3rKL5z3ROo76YbehegZzfeUOqd9SD9FTl9jUHsYQedQDm2
HeAhXBPYHcf2OJeYkD/zJiFnNlV16GLvyXfnu/ceQQtnajq+wZ/NiPt/4xGUE6Ah
riQp95UScXbt2b++0aATDgrQkzjMmjjpUr2rPV7BNecF8z8J66PdfiQOzuWSJvht
66nc1wxiAmNJSHnD3Jg2YdjsQwI/kGDvl2lVOYYMWp2lMBCyLDyDRRQOTybsyZ+J
0hsXQyKAydwT6IRDu9Arma34Duy2VoU6tEUshmtM941ZpOO3tKIq3ZLo0nVDyoi6
zij7BS3w8wVe4WofOyJmxIn5us1oiBXBiqpzG6aQIvbK8MoQAkXnVNuxMP7tFzVd
dMGEDJQ6EeKPMw+sn9DZJTh8e1EDvk2gx8e1rUktL1rWN4pgY/HCVsXDzJLgYii3
BDJ8JNgdhyDuY08HGA1E96ocXDXhyD2BKLC8ZQV2U4lSVpSZ976DdPCHio5+9W2R
asms1ENLFsxP/fE9x7EfTbeQhGjy8Xwc1AvxAE4iS11F5+r5hz7U0E+GBVOoSWBY
eOxmIy70ynC83L5Nnja8yoRdR+qK8Tzvo/1yOLcP+/ZHOeZnYLGBM9+ltPQVLnp+
YPHU36akEIAcfMqbpixzLE8YWh2IQagzKil0t4tyF4P5hb7zRqIVuIdYyM/ke2rM
jpv/ngS5a4I3tleU3yD5u572LpAaod8IXKlMekafNdxHW88nxk5bUTdRMCyxhuJW
THWhaNocZVfFyGMXbfOtJgaynKA50x2wRAzhkUpYaUxvjL3UH4vO83dcMNCA+qz0
T/gDTOeOW7ShgdObMGSYZOshQJ1R61SjpxOseezmsSrztmtFbGv07m3bFiCQ8uns
LoMu/LfR6gJqJWAJvNYTEaYqnneb6lXIYQGV0yP/jlX7tashvMs+CulR1QuwKtB6
c4SWRA+yfjbN7JWzZsfd2Nk+nE0thv8nMYV9sTAi6AJZW/se2T1JzW88H7EdBwRc
sH/o0csMfFPwOFVgrqVt4xm5TZW0oIQqZgAL+f9ug2u0vcedvYCvyeB00KNMhLD2
rv2Wkfd44MVKCHKLFJBHnGxny5/7g0VGwa25irpOFBrEj4P2On+Cw3jceJIF7x+d
BEMLND7CvUQzWn9Ze6sY8GWcLW02wtBv883gqWVO3MbTf1/m4tDRQhJetOOuYue8
1e0YELcgZTY3HCUCmyK6wSbIN+w4WEhqFuRMjiSWa+bxtVMcURtNWa8l7q/Jzq8j
y65n+YoxfQ8egYOIekxsH2Py669EHtPToIZT0iczUqWkEMD8iZ1mGaPL/unbY57M
ixq8HaGpWStq56m9KE/NRjjAotc2Rm7/WPMfMZH9DhTSrtWliKyzat1t6eIb1RYZ
Sp6bnG3/JqXeRCCzdI+WVx/eUrfm3awUf/XXtX3Jzzx3KM2h9LU6hhhOFBPkquN0
p0dRloqQ+OyivAzH1YTAMj4/ahXIMgrjdqZxtA5020kgr/JIgFu5AfXMv2q0GSXq
YCC5TI4RPqcvFTAy6yq8AwZ088crx1v18KPgRmaYlHRQ/dOWVHmV2YuOBc4/AAf9
mJo+ZESHXBcEolczBo0zZrm/ZZAv18dxSV4YABRbmzAV5YAyXQqdfG+8wgj5Kqfm
312Ni3AMr06Op/lCH5lgSxRL0tCoT+Rh8gfAanj1JOmlEU2nJZT45Y+ImZtd/4lp
BjV9irSLM0kbYryb0LTbFvtoZeLdTjbyXG/gCZC3OXVegSedcfg8GPVhJjWMYM6R
wtknZVokmmhubD7GIML6gtQXD0Zd8bt5mnEODjDCRQ70w3LEO/E5/LPNjT4GWFUt
hMGg0iu8/c5/xaWVZTZohpKuhGoBOUSOo2IHmBU/bJuwJ2gOFeX29/TTkUGquQ8g
RaZMcQ1K/wha7VmReb2OKLSM0ZW1JD1iJu7mTfFJ9ovI5V0pYw3LXKjevduOIhZM
JV9tGE/xMOeAitO9Jfolpds46xkumwpYjoV3T5nmDXlGygD+wlb49+Pfny44uL4l
OkP45kRBA+p2qasULcd4FxdrENI3YzEogIpOBbN9+yt31UpFiGvunJvXrybHEDy7
pzI8WoLwqUE/IV3PfMThzC9edJy4IMXhBoWKj/PCDW1Hw98kIMTgB1BK0QLnOsLd
Y72NoQZYdXdIvvlnx2Pn0AcrlPC5lg6r6Lll1Yr2v4SpNeWAAUOoN9L3DIDVTMc9
HpeN61lqy6HYoyqMkLLfv7xxDP919N7LDDbJDgrRrC0FarHK5gaMyH2QyiskaxV/
`protect END_PROTECTED
