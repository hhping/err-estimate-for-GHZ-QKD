`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IyzuGcFIWnSvEyh1oSIXOcW2Z37+6SH9zMAUAfu1Zjhi/UBnPJmLYav3PW3nmFb6
rPxrlLo5vnYnn3Df5G+ucwWbJRzCnbCojmYw1mkbIIJLl9Of6GzsTMPKsNqzVo1K
yr9CpGLqdf97lyiIWQm6MJ3AsFH2gJp/it9sb5omkToss9pOmx6HzDGOXV2Yfzuq
sz/ugAlUqntxCGpAIQeVn6Ca8n5mCic9ukWPrpU5/of+CRaWt0kUPErcuoutEL8L
5gfqVfpucHyC/tfwarq+tyF//d8F0ZiYK/Ql4kyLz6IM9v9VxAUGLyLYDQdUL+w/
6kR3C8li70g9SNmT5c8R4IHULvrIJqlqYQ1u6kiV2u0uN02+yFA+YfhjpLT2RTrU
IWsFq8VpDJvzXJpup1GReaz4CqEpWgGH9tJGRkrJACxnBZFiSR3URbEzJ9FW06w2
I+hIHwaP5g+M9dvyW3RbjBvqqGYM2qc73Sliuvu+Jvc/odVrywoWVSOOF098088e
HigvuBt/2oPMa70SUzKe1lDwOBfMiofV2pk/uF+UQ37WMc7iGfsu2KJOegU98t7U
oa7UafJ1D2asGNT3uoZdSWmk7JItpyQJHRS4y6F7nXmMb0A3gPT8lIcLHN79/rS+
GsMS6zRt1LTUzfTwzjb1XmWRDlmnxIysxZ7E8KbVfUjc3SD5Pu/ZzRArQNUlM3G5
owtbPXeRAsV2+E7FL4SUzfB+8Z6n8GjUfYn/pvK+oUwJ4qh0XEi8VRm4E9hwIkGg
VakLxkseK2dd00pQpDSFOHluPXYjapa9hBhGfBusgFFzpyFBdckll3hxHSufTvry
TQcxs0aSttm9S8H3vkC9KVSLEmvNC4XohzvurFe9DaIBJLJcRzpZbrnph7e3ABFP
WOtC4AzGKXqGZFMsUPXgiF3u8iWIfXUlgKxGSyJCrr4g4lKlJ6wfYGmcw6v225Od
f9IR3ky1YEafnyRhS+8Z6qia2Cp3U4zII0WN9nVi08h7tINkdXe4skijhsysfohz
tqRfTuPePauj6PRKP6yd6cU68DzujQkWRLDBhaMLHuNkyI5AJGwIBkGAT5BNcjHD
e4BKoGtUIRl1jBzov70SLSLltDMDDO2qC6PWt6qJyi0aPNYJqVDJmsqHY9FT0LPP
Ri1uVdZXSanEA6KwzdXHD2f8iBG+MBARIEohGj9HAkJnfwjQvlxoW6tkoEwkXJmi
xdGHqHP2+OGa9v2kUo9gHjpwV9q8Zfvub33p784B6nPsEPax1R3/uLHArqi8TlPo
TDn2azClgcjz8yFZadmvP78N0x7EOTW5Y9gZfQ8/KyHol3HMKBv6jtlXrM2U1P/Z
hLukKWKgRXMDXlfzk90HCLzl4qsvcpa4u7N9GP2EQHUfwHvchrjAqr7e1+RRsYd4
UEK7LuZvMM/wl4A2d6gwP3ytZMwGWh9k/ID1/BpmjxZBpwvDedULX6fuRen2zgUp
NgzGmi53drgZheEtIrzAeVcad2SKJdMQegiCv8BVM/ZP9FfxtsO0L9R0vfBmkltM
Sq6mYrEn3K6+N3otK9C54Z99c/LAJNNlM0apzKyculV9kjakZJOZUbiku4e+q3ey
hBvO7GsKk7iWQ76IkPaubVA+6J4OrFEyMyE7tUeMurykSi0C079c/ww9uQpqB+v5
Td70qc1gTMcLOfvnJys53dRHDORMpusSmil1NqvJAvKyxwIWKMQ+nlcsYkEPecXR
CzDsefGBrEqsFPbpeLSYb8aPvD8CEZz7Ooc6zmDb8eD40X2CHdKRbCbM2i4Sda+I
ncVUforTS12taN9C4CJYAw==
`protect END_PROTECTED
