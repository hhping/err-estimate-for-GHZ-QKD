`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4M1g0le0j19moYytbTZ6hb0p5N8vRshJlieyLxbIySIfJm53njaKgE/1sWSWXCt
QcjvfY8tcGag/k593Vno0Ec+EO7P/cKLnFcBdeLRMPo3gVVWwRnRI70yAPjbNBtJ
994REkNVHuT2097puBxDYLnvrkC80VnSUYRNSmInNTaLxVmhCUGDmM/PLwEf/gJB
DjZCu77JOLkYMEXYvkmw8lgcErFc1WAXnMdWxa3BkqQlusE6pq7PHSm61Zqj5Yt5
PmniGU/FeIJW6d+1gawDmW9chGgnFKJio/xDMaFIpyi9kXEB92QHwfA0voBhRFC9
fO3oXehsltOES1Ib+wPh27kdHLWUsw+9dXYenN9Hoe1vfmBkRioyJQH5SBfawRRI
I1L2qb+7mV8izKP41jDuGXSPGQVVjrmcVF6MlyIl6rUIThYV04tyqq3M+WKc2hju
/vHdMtoBCwqeskNC+nEtvetSZt9/37pnwqlJUiVfJCf25WOONgLpdiSBGk8Zpho+
vvMn3F+I+wTAkwffa++1XiWqD037hCdk0h5t74qxRxnrCcHz7cwEekvsvz0LkvBB
iI1TFOavUIr8HHMiOe6ja19WVIGaZNb5FZi9ixAygb/355edLPMjkhr2A/13nTh6
40SDkTv6TmIpCvUke22W8fFSdmIt4awb57pKRrxNNp+BKMKdw0Ibk6dh97063YbY
EavjW3Mdv0tboRMx+oYDtHVLJpCghz79B1MugDW+wKfqmZsQtH6M9KH2sv9tlLQj
CChJLFQZj8/EmILexRiH/dMQKUIZkON2SKxNDWRVHCbllRLc2ye0P+umLDEwhN/E
mcKCHAhM3/9ygW0+bRqzztBcu+X/jvayypgszOV/mgPHARbxneYqSIsQvw02+vpQ
WKa05JJtn1JZ1wnCgL/9cjDNYjrBNxTRJ6+weMMpnGkkRO2jITkdjPsCbXBjtNDC
IeG4wE8/AG68ZwxRewA3WlZLJuOkZmVjnTUh/O4DyQUMX4UeZaAdW3LGXTRd4Dvh
dLNlmNtD1tdF5Kc1xsG3PUk3pIRuSGxxG6lWpaKj6lAhwQUp09xoBU3xzjkcV6j+
Iv5e/qTliJi5T/An0587IYKDeQIYE2GqwqjoUAtWNvE6y5CvDOfH7XXhFNvzHcRG
bA27VtPJ42bGaLRNGBEO+lOdl4+lLgk5PweV4TRAI6ARwgPPMSn7hElHcE4JOKod
bSPvDGi9G/aC6bSAjR+OERMClhVxDpqQ2TtYpM8NPbtpSpq5znmrZmKhDjzs0XVc
qHPy5UkuhqsdJ6yzAYjbaOIoyHs8ix9QAd3XMEAq/MX9Wa7rEw0FQH1kvo5lq1vS
psvU9c2q9b13Ixa6BanMSYTM3rw43hRZLAm8J0EZ5p10Y15DX7FNEtZ6EgsBH2c1
WDM+qGWWlIIgEHAwsjXGsZ+SkWi17TZ4OaxwaLII4mDpMHwW7Yusg4PulcAHgB3h
0ssVrEGNJxcRyW/dAT4czldaxN3fIr2ybi1I9XSmITGw3N4SkBognt8JeQAinYBn
RT/8GJR/9WWlc4nawSjulUiSKRVTJ61R+U1R0r1ieZY=
`protect END_PROTECTED
