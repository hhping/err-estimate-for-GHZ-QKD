`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ng1TErBOfaknKCTXCaPWOVktwqUcgmSxXHwd9eFBL2hoRj9ZWXexTBc3gEzldI1a
+9R0nz9MTswuaV54brpCcpAbfa9eE0o2kmUWQ3Wraif4vXg5k9p44luME4SrSHGD
4LJGBUGHrzJsmKRqCg9fy13nV8kwIu8+d4Hqap1aXTo5AMcO2Yl2QbJ/SzMmbZha
SRuHCJ6wdzHg/1Zry/nGTo3e8iMLo4lLFTi5NVMm/pUPA6wInXs7Q8NlQ7K/DjFe
pp/inUr6IruCVCFyqx8CO9knS3oQk1V+t8uTdnADhqiGt2zZ5Ydi8NMdYcyscP0z
8uc8VFdf4Ii4rO4fqyPvd231jBArb0ZW+khZT26k1aig2r2YrG4q5STvCQkDuZ6S
zFZRokg5+dIc46OWwpP7bkqEh1Br9d+GBwAO9+ZXaNLPnRXxzi93zLA65rihX6e2
SWTShJYP1grU7A+gm5nM/B+dQjTnG1uhyptnQzRyj275n179uRhKVhWEBQpx10pH
LALHh7BzAdkO3VPmXB6piILRZoneKVJcobxUpTRC3PXVo9X9yYmXbB/WaRnv+Kpg
lQC5WQWMbgGlZyBdjWpS8naL9cmgRamCbaD8R+MqxruSp0yDSjEdfxOc6Rgfhleh
daC4Kkd21GBZAzs0GC6T4pISqjnZC+QiBA9vCa3N3kLL/yeMdYjwmfLAJ4ltf0Gm
`protect END_PROTECTED
