`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1TuHUOlUSIgqHeS3oO6wDkCrnHj79va76XPxO+0oozwTCZ5qUI0rKw+KKqJbgNot
ZMnVNX3QJ7/V4WYDvunJLhthogQk9REOKGVs4WCBDh/OJndUMW3JdXQLduj3HbtI
dasmRK6ccI0I8KQq2HtZXZGlp+o9TbSvadGhJWInLeFRYivKAioTH1zEuOnAG5cN
frDIsaydpYyqhIybegotoNg+KouXQgyTxTG5LjPYYY3SMPzL1mknn3lXdLLBiNK7
hKVcjSdz1huXLMaM6F9yIZENP3QIOLzJyQFHSIZZ2fbfkSKXkHt5ObhfWkY2qCX0
4GPOlwyNa0Fq5KlKIzmb78mB5HkXQCWv5METN9/W10EwpGnYKgsqGeKp9rdnc7jo
m2UJZuh3/2S6JyvU52CziK6PJ60VzctTpjt2m8YdBydYp/tHfmUyPIbt6romGM9s
9C2ZcQn3FrCxlI2miuUPd0I2KQOOF/U/nkGqbltPDqx6ZRwmbNlSeDin5cNA4N1j
mIMCFkaEBLyjchuT22OYYSLGcpe+s4taPL00SHhpVowcB8DZTU5xmvpBNXgqeDJ1
N9ru/EeXS/YoTnHffQx08ew5HSuiSTGFYceup+G1BHatooh79c4mX1Wgcqq0efyZ
4+A6Ky/51IBWjbRfb42rt6SBoYDV3LtlCxD+mQkq3aKmNId+mgBZzL05bK1sCtrx
a63H0H+X94nfLAp7TWnmQJbDFaRlnGfH9wB7YwQTmz5bmGfrNSJCR3iPZSEnAAFS
oTl71Obp2nJq6I5OaeQ6nka5OTtehLgkOoaPm3qVu1x+sBHvdfllkLkFQhyMP56F
3esm20Pa5QMtN8ng0RpLqAGg/nYt15PLGLXkqNwxjxdDr0Zp6VE4heBUZ1E6JrMi
Ns8ebGH46d151fYdZ62HGWao16MX62MtOmzUlI2OA+HnSAKoSipLsGSZAujAO0jr
GfpZWEX2YCb2umKjT1SYKl45iQv2QKGFqKGfHRlxFUSJfGoY+fpo0oBhIzEkWNsp
7KLIzYA8P7JepxV4Y9JREOJNGORc1dQLugFm+h7Xhc9vYGbobn4ph5HjA8kaZ449
+bUkxwKZuU12N8dKV6zXvLbzAkoXK6gMNUw1t11GQxC1hg5LQEIdFbpEcPCsTY9f
QBiDQZYai48S8bwHgNA8B2xDv0J7xegenwT4BLy3eiDmTqEBJAJRSvMy2dxe7e9L
IhSyqIC3EsFyAC/sXxRbo/0bsIqi9ugY407G4xlC1ZPTSRFKRMx6WYzc20hCceoH
P1CsAnJknT3uQ3SRDEp/CwbvIG/uW3jgCkDD9aYozMYmzqFjhFFdbWlGFzC3CDUz
HDbLOiQYBhq9mYzXtRgqAzL3QnLrZyQdhpr3PK2DCgkaK1m62rQsBTX0QRj79b+m
CPORNiq2GcT6ep6F8bY6XWYC/MkBDoYv7mNo8llo6kH6RODLpF806oU3YhBkgvHk
VtFI92UuFsVFpxIFrms0bt0np/Hq9aZVxsL1TBmwwRMwcDqx9evWeeOv4C4ysFl/
mfLNd3rI260ULnut8NSQLvjp6ovLR59SMxhUpCrMBRdPodU3dGxSaIpvr36XF6aM
6mJ0Qi6zOXuYJe9GmLH+Dg4UcUnwIf57Lmk5UCoMo1W440mQOJqG8SKD0LNbxFdy
GfGHeISQfe0ezBsUELwHHq+sO+sQ23j8qZgPrwnTZDmdH5GefqJyuiiUFH4KDpGO
6jD2Pi6hPWUXxEOsXCxmvJsiIJjDeVGGLX5BLtwQoDdG9b+gXMpwUlKlvukqexXl
/lkpmywPiVHjDVe+8P1cHGQX3pd4n1vVGM3TKQs+jT4f0Pdda7I/xbJWVbVgDDOY
rYrN8gWEKvcshLF4X/5aGbfGO/YTaHKzkjB/B/KNW9xHT+/4QRuHyahWIiX+GRCj
vuENgecQqA8UgqLjt3CFVTAPFYYXQlZK84JgG6svbGQT+RdmzGX2NABIS5XEej4w
+772g1FdPoX8BEFkaO7oj+lTV4NZj9ILRqEgEPhiCLkMLK8xW9HW0rKwWEwjbpbu
cylF0WZM6JP1kzFjnDSR71lBPepjb4rrXgnK1FeFIoWS40CC1aXxsSpJCbYoQT2w
TGdi7bareKqMamZeXrMQciPcDU7ew3hHXxyPOeUq2GDkdOVnW5bVQD/Q55sak8v0
519+cuf0S/+HjpEQS9rf5OquFTXmwFq13Q/p5eDKE/DZZGS3mweX1TofynCuyoLz
Ivo/yp1j511DD5UY0OZvrX7LH+v9/oZr04RLSPh9AWLQTaRgSDgFTw0UzeC8NS8E
EBaqvbZagi9F69jRcN+Zmy1gZuO/pn3Sewgt9fsA6PjImT+hAcbsqGSud8TVCMZT
eKSGDvxCojvUuiLExQdVlXY+bhF+AyHM1f38B9fe/zgorVbsff266F96tO0tgY5v
evAubRvHUI/7/Yzzpr3uJ3+rcC86NW+gkxSvNwPiP6K8wn5RmtUDsQrrdZPuDdis
GrmMIty5CDgVJKLnIHONKpOApD+WQcElmqT3dVVRJjvlRiPp7ZTfdI6GUszsk+Fj
pCgXDk0akPXai+ztV1+JEBq/d3Aotfz3lLZfZ+xuSQPRwoKh+d2H5XlGpQ8aHg5m
/QnjDiIPWCH7kVLSCq3FYdNEmYYLxLiR5+/J42jmheM=
`protect END_PROTECTED
