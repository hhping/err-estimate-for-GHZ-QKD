`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
px0MFNaaPQLHYObGlF7OJMCfvxv4zVG+GfbvrgXTIUlaePtMfDQmp1JF/pVoajhq
sXctVwtZw3VjG0+gUHIwft8BdcySSzKLwgByBqTHFoxpe+w/K+xG8oAvOoO//wFk
vBIOy0T8COPt7K64iKmM1mhN5t68sN6PdeQQZtQmfXMQwtaprwShxbjTUVMN1GGK
0DZ7nocdgC2+Z7OIwlVMUh3F+AMk1lkxlqPUR286R66rhUCaaX02mlflkd8b2bmi
p1e1eQ99GSeepDWfor6F+R5hUeT70PMMqQ2lonxfnWuWBZWbpKeWzt8oAzfTuuNz
OXU0BRUTH2l8kYnSyINwzCsx2qWyUQ63eJivCtWgPQP+wBM3cbtPZtmT9P5kjIxt
XlwFGXQKASMldBNJckQBpQ/kuI/uzQo78X7+MfrJHYeASwgHpYBEbWD/i9Lo9Rlj
o6Sbq+ZsorYFzf3dupkC/qb9u2yITOJKXvtWk7hqlIJfXcA7gFX7sb1+ABn9KJkC
jxZy5IBV1fXZB9NcJ+8fset1s4vD+zZjsVFdrDcaRMSZyrjMNvVdHYuQKY63KXuB
wZsbmAwIard1xzw8Q+wDoGVXpnIGPAZ2k2oer9JcAl0CUkYDlpofAKiKwPi89qea
eADU0DsOLsIgYByaPyuo5/CAUuC++orWK6X3sVmAuyKKao+P4Pu9CCJxuroYSjbP
7vbiekB1gj1Co7QL/gnAxAo8CIOwGFw6WTVXnZ96gemdohqH++Ybu5oqDL/j+woQ
WgH2Q0yp0Tnky14NO4en4k9oMOufwXGcS63NdEcfjmvLmMQB8E5NqchGmp+R/vAY
A3fTOKHwNxZ0e7c/3H1AjgNjmZrZebczeTXsIDwieVf35tKObW31ag+xDFzFqqSj
fVSwutILPkLu7ufCy6lzIz/Huyho3uP91A5BjcivNB33CeZj1bw0eiNFoVRlmq3q
p152+joSKRKQ1Wrr+YaUUn16YLL1LwtuIAww8XWb5UVVh3ZWfbx1JO6GeHlDlNnt
3edxEEMRlxoJBz0RvqB3FZ5XugG4Fhe2q4/+nP00SG9+qGudMZjk4kFwgy+Sz1Jr
xK/bXvDyHdlQmG92x6aYaMwlor1/ENDA/jJQKz6cQb3Sj752FekrPZgBj69Z4rH8
+86KAGhRgtM2pDomYI+zdyzbwYzNMD7A6n1/4TRq3sA+3a5wUbs/lAa0wOE7BWZ9
De6OdWltb8H08YlY5dIqVFHOWjX/F3a0C/tPvbErjCOzaypqhCrgOhg9GBU4JclI
X8WnVEMtr3vINM3qEVwgqtTFsvWJgqjJFUlddtChzAUMyGomUFFsL6ET6RDfZCZx
yj4/3uAupjgJwpl73jb8CUgqRXgfj0fykPQ3CR9cxxWWjA/BrdNhseg707En8cZ3
m0FXRGhML86IrU/TEBBvU66lcLcm124e8AxjE5/0E/arTYFncZk56hhu9FBRq55h
7mkoegf2FAWytwD/VExFIcoSiTokNA0KD2aVeWQ+sxsYBfgJ2dYQqqW/7S9Lyh5j
FCWSyaX7C/fhSOdjfkL8H2yPj8wzwSJAq7Q8dkMSPJDskWPy7KKF66jibKJSdrEf
Hr+SvPHXG9Uc9dCiqY+np3bfLxB9VnLAVxpD8LkFRovXvT2vWPg5KEBfSLZjvbwd
7GU6nst3qNt+pMQ171LLUMlwMyLoAaXJeNPX76eVIZ1kKC+b8OjllIOsjPy9ZjIk
00W1QKw9aM1bIQn2jLIz/DjrZ7RCCs7UY5q99csDIiYYnA0dnm9+qZqULFSrYCgK
PnH6rsttafKLffnhGYr/bxpPOREp8JWl703MmFjO1hXKHdTAakJ8/iUwTRsZ63eL
/80pXSiOWhFmZetzyX3DAvIOxQWvIMqBOwgplmtaUyoG03rak45On4Iq9pjWi2hU
W/5jdapcaYXvBKhBhcu9xG8UGitLK7wpDQKtClsC6PHDUzlBNlDBJna/j2YjAWhH
3/PqxCoNh8JS7NRZkl9EWA==
`protect END_PROTECTED
