`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gHDMjgXxACW5Quu0xybwf6lk2e2eQdgvBWPnoMEw/RVS1OnmizAosX4cfCdJDuSZ
G1wfagwuDVrwz/e11bsWmfKVjVC1Zi4lT9QWBfcbCsgIOq9OdAXdHXXHKa8diQOc
+WOEO8Rz+fd8Hk4e7RTfwkWAH+UlGV8hXT3kVkgOFF77FYroD0PZUC0OQdLdBm4b
U0z9Kj6fQ4BXcBKwxsdbYLNZrpnaErGIsE4TTV4smHO7qOTCsJED1m08SDkYTiNM
0QK66jfHqwVB8xh31Nt2iJWAKEnvFvy1+FrRKYfLcwhQtJWHYrp/BjWQ7NOGs9yi
2i1F2lJxhbd8EcZsFJoOeoQ+bcpLXIMt3zjpQgpAGud4//kEjJ5HE16Gmv7wB2GE
L8WcE3rodFqV1XfF+7CrDLATLpf9wZKbnPpGSPG7jSFa/dJ3Mdq3Fv0eskC68adi
oSci/A/q6ev5cHymXCF0DzbSJG/+dBBp02cS+yXh+HEzBRtM500rzngxzElCPNqR
HD0/Bam6LGAjnjfEIBmDeYZhdpupMtSsBTV89t28lARNV+LfjNM9ZKFJ0vryiblx
w9wdEAHMRHXUw6NKFzmxATj8rl6H2au8MvdzGoAw1nyuExXbeZcxzipumlFTJ55v
gtcdxRCWaWFqWV9U4RtG5JfZw02P+Vw19Oe7rP3VYYda8S6VEK4UM6YhxZAj6O+v
Xd0Dg23FTxWHUG/4YbSGoTOelzRSQJZ2qeuU62r0s1Q+8Ivk9JPJdgtkVczZgxbE
+weJLona5Gh5nIYkEbbK8TXXxvYT9bmSVPMEPauFr3F15oA1LqPu0UrZ5rVzodic
FVeKTdIIc+RKOP62Fxu/8uYT1hVIibHWgT9v9zBtVWV94uTr0e/Fj0IuQs/PGmfB
8JVQX8wFFT4DLqG8BtcmToE/eE7e1wGvH/MztFDxC4fjncqbjH2E0Xxs2XlPCBeD
lOCFVVFZttuHQq8ehLHtNAY0JcH1RoBUOOnalTj0JGWV7c16hmcjg5VekIhas/Ky
9vwfvx43RBLp8plLvePyfiwoTKTO1XPBqkxdapfvBD4f126OkwBtCt9B8Pc0YANk
YeUJ/AnEIMVA6lEoAiX4O3du5vQOztFfKAnapM6ze3WJqFoglzBCn/kzUbNgBY3o
SNsIBKp0CpkEZh9DLRhxHIC85lWydfhw+iWe6o43Lq5/iG7CAOPmcbR09FKMSyAy
HPOympcd9n9DvUrE5IGFZddkzRg3CnKxWv3k72yHjv79qSCcIxA8oOTkPXQwuu01
7lAMJgWBJ26I88GIDZf3FaeWz2D1naesOzGEZOFD4CCh84v3npmcjTdrTCqBQ5BL
JcZIHijSUCLDEQUjp02HXDcYpqXx1ExiG5XoNJdeteZIiu5X88Z2z1VbMah1KIdy
DqUTaVBU9sJdI9wxhVjywxmsBolEmiGn4p/7s+qGh6fAFAJ3Bx0tIyrBTiYtL4aw
4CIISj6LtCj1KN/oTbhEC9TTP79MnkeDpjws5Eznmys9uaz58hJOfC2ARxTPYBKq
X6E9gflHocBhwwFCqdjzd6GPotKbIzQMbfJBBH+XgHJCzM9CEx+v7IpqE2a1VgEH
UHCPASJ3i8nPDaYENQLb+xSRqiqU4R82khuorbz9JvHKWhpOQ1UKraHVbpbTtUg2
QRZWeEQA8dsWGrUxi0bkzqbDRFArgvdV8onCYeJi4Wueut44KftmZS/5a+xXOzdC
4anG3XW8dVXsMr8rtRBQIGVJao0xeMYG39SiYJ9hMxywytP64fcbLZeEcP+wDcfq
eC4RRKp4L0N5g+Uzw9yAj7efco1nhRNYu9VX5tNGF+nAYjkhAlQaKJ6dNY0LZ60h
EpZqGL7oeDkMrWWYm/rjcU81NIcHdimD94RioNXyO0Txc0EujA7EvDzR7Ksyp6bb
MS+juG13EZ0WgTKaS1hjpeO8GHkFqr8IL+x0xBswABjk60W+TalEVIiZmDPOnR1Y
R8a6xky6KklxV/3sOEdERvTqf0DaLeQaHseN8YixIj5NfQktLson9hIo0hVIGhwl
gg5zrbtZ7G07DbqfFkEXG7hJAtjQn4+10CemRaP3JmmzyDQawIE9bvMTHhz7eRYY
FO28NimqeWtyXIjD53M22GXh13QkPnZyUnyFAH37Si64PHp8V6/9J11fD4k50hAU
jSXLRWjxb9pvjBQI5gOlOwEwbT5Wlf6tWa8cfvLD7lrM5bF0rWK8WWX1gDCc5Jtz
4haaT5SGe0YKRzMNZcnZUC1skKOfoxaaVtZo1NCycYnM4xMD6Wl+ToZS+fD5mf4n
1PHsaPN+Fn5u8hT4KIU1gP5pcpioMIQB456LvS5vVOnCSxefIJVqlC2SdmSiN4H/
5xh4NVeNGYwLYH7Ru/GoB5fjC/ANhsQ1Cfpis/jlX9HYyWnEIzOn4eehXeEjpMC5
mcYXQ2iWg3IbqJZMZr3Aw/9VphwgfNdDyiw/u29MmJa6F8e9C86Xpgnm7/pw2xte
H9Ty+nrhzv3HrDUnOvvXvBbde38nmqRWw72S+0CQ4iUcoXhtHLVR5AmvKymlIzgr
05Kw8o3oSz/nZRxSpza2iuth3vteVvfNpts1nJC2q9xVjvP3mH9kdSewaM4SLlu2
lkLKkOYZK/9zwf0CX0+r79Muq4sVmRd1VJNhXsLE5Q+0bzeVrqd+kwfD5cEbslFd
gp9/+l75siXSq32RbHCZLsuuo4FmG5ZMW1PLyuMtvDyz+gDu8i/R9ITkSmxo94+m
ZSXKVO59iggSc2JXwya2tUZtCSDF41/qN1Mlo+UIjHyw5NQPMKf1PNM667hQKncm
F0HEqapCQd8+iRKTLTqBlxqXRthPUIxJyUNPt2zM464LXSbgS4mkavZFqUNNLTph
tm9xY10h1cwSY+GgKavuxMhI506OuAgtJtmriGBpqOIEahoXfwm8WiDrrki/nNNC
jj4+Djl+IRDLVtor9eninV/u5IuSpLtt00vlP3nIpStLwDNrMVxVOHs9MvQv1hT5
xJ5JtJmg4wmy6Y62mxQm310mDFHPbj98e6a4F64u0nCeSPqa7yLbBn/nRQmemGkP
k1xZEF3nSF+GApJwBC+WES2l5U69NAHl9Vr0WM8Wa8nXPyydKYYNC+VILA95dREl
nZUKm12kfe0GbwIDvjQPTbXL0S5ZgvexvcuC0j8Y+wJx6aegzi3Y16dABc4YnzlJ
oTPnXnfTksEHo3ZRXe/strbYbop0WTYzfbcKpX8cO6GyQzeH4I3mvoG5j/AU5tua
3naBvdlR0/fzjUAkImn8O190LH6PMoz9XscdAF+6IvuBNvtclVfEcG8FXEdElE5a
SkfnBWnR96uOzZtHvcLzQ5YBH4nhS45HBhzX/027V20kNIl8EJatOW8C87VyT1eK
9MyS/2xGfcOgZ2BqjjkrqaPgLz/ZrywcYX1xFIupyqplkeGH0tXJU1vkAaoArN/X
BnciGfKs9JwIxn2vKaCpydQqHbnXHahrihF5Pr0GmbTvJuOtpaDgHrktrmVncH1O
D+MF57diDTtk/wV7GfXVC4xfwvIfeosmrkOuh2q4roCtKIEwmR3QRbV+3eJWnc9d
OUcNhu8ju/dPKVjaik4mFfI3IU62nn2pkbHJshCHsl1I+cI8Juzwka34RTrzCys6
yBZnw075z2WdyorX16z3+g==
`protect END_PROTECTED
