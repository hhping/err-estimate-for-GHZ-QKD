`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4am+0eUO+P4d3UlHKSbQdWApSZVjkYtXcl7l1vRJuSUE0lzsHJM/yrlhlmfz4Yhe
D9Gn3kDKd9o04OXyClQ9Suhhou/YswupQS4t7DnVc1a/x+y0iQaVGMjNaDKNGtjX
O5vlKJlcQMyQ6XwjIJ1p87QHnyxR5e6clNZQYcWCpaXMX6sIzQAuyqXMQCD9pZLq
VaKNxYBJD5A8/eWW9Pz8ItVbiYX8DZYygV0sfMfRqe+yZWND5sC/61XUekkBw+0u
ak8Zui0CDeN+/WgmWfR6eFRXUcuoSHtsAxJokLYWeaQSjDraRCaeQRsZsIgh4kFq
tEvSR0iJxFKW7FYMNKDQm/l5uvZD5MtLvS/GR4msOlyTqMHnQ09akYBkWg8IgkrU
R4SvqXkiwfjUPtDsc8+SlFD5BACrauYIESUpjcsbbvlN/41aIZqwktAIWpYOw1sY
VrWLaslpioieYOXB2sZUvFYzT9I0Nq/T16I4jAaIb/fRRPAaMlxcPTjJkYjXAoW1
x41UZX8xz1V0mo3jiP/M7CS+yAd/NeRL8fSRoQ6sQerGPTHUi5pew2JJcLrLicVW
t+Z+ZWu0bZjHULc5hvLNlpvXIvqCkMAXKK955yeJckcs09pBnRvAhFUGd4sfhYoP
56gnhDrmzAi+Pjts7H8TVVQ97UU6+U+a4ULBDiQHv8ssI/pvjaftm2sRu9FV1DdQ
bVFhMHy7wBpx36t0lfp4b9zOryoRiN+S+AWW/Pq21bmcElTckWVunMX1/SnBZiQN
Got3gi6TU44xA2m+Pgfzb8xuCfE+5aAddSpORB+ZSM0zksRB+YI+0mGTWHHeXWBw
0CJ2+43dc0EkvSDYJ+WFx5/b4BFdL5GBAM4Hv8DpbGdtLVUw7+kBuyTqb0kNQ36K
dlmOhBtVXWV5BIRCa97oqoUoA23of/22Ahu5q9G9R0T6P+Ts8UnYn4Fl8qGKnpld
yq2EV5hIFqfJ+xCo+aHeI71tsTEkLMf+JYoZpTbnlGtJ8PuTvR1W9u1o20Vp73VG
hO04f4bj7nG+vdHVIAim5HV0zQhzrXF1HrxOO2AHlHVZZeKo/AxoLy2T+etet37B
dzILQ/TOQgWMN8QryBYkMCGqc1ZWHfw0VZQiByzr2NSGYJwpKkPClhYYmrwje0zj
tVUm+M+B85wX9/rc+wEhYRLa/MOOb774AKRitJS2gKY4UB5xU93t9M9zEYRQaq2a
snpUlOzmauaRInjLq1wX3y3AkHQWxsC+yTDda1SPUV0p0oKKUZ18DHnsqc3DDm/R
yiAm/7tss+WlJFqQ49n2rYmbv0POhTMGOHK3PoDA8MgFq2OPMFO3douNFhLApviC
lWNkhoA1/FPRSBCNXsUx6vvruND94C1F+UYc/tLcUUZwMhMG23qj/lxVXog7bKLz
rhIS/UOa+YcMLvH68NGna4Jex18gjpE2tCqZk9RxqzSwJPvcvVhMMXOgNkTUgIvZ
UdyeAwfEpfN2b70G6UeuhU9DVifXbW2sgmmVRgpsxLz2f+V65nL8Ke1AZ2ZE/ZZk
cCc2nhHuZ/BX8Q5R1rcJ1qxTW0x2kA7m5Kvowj9aI00qb9rZfjtB8M6LOO3cxdEI
9vM/pyonME8JAPWnDMHXbnBg6XKmVLNd4QdqIHTN9vqnY2x4a53Fd5SroGUuhWOW
EWJGDaO7n8o+ThnumyalTHV3dhxRK/gJFnLCPp2Pad243uJMrdFsqBkpmDlNimyW
issEgcm9YoObeIUWoPnlC2B2vr6SwPMJo4WxrIe+RZjbdrwN3eJS6s+0wKQswxZ9
xm6btH8EG2nrZijTnv8+ae5pDYOf0mEWSxViyujbU8bc/nbs8jYv7o+NN/qzoMdw
gF83Zbhahr8wQ9n6j9qm9Ab9MJWrVWaxeJo6UrL/F8t2hYgd+r2iqNNshZCjai0G
PdcZnILa0Ttx3TWJUQo5p5MJudvUbcDkrjK+UruJJ+rHdskkEVZm6qsw2MlYCLiO
7iRGK95EN6fENd751q0r8WFqvT57MphfKI4VNvEFlzdH3504Q/0b+TJdNXCRhaXX
KhULx+kGAoMHdIeE16hfamu6bZ1J4g452bUpPPl/EAyziyj0J2jYUtXwicSNwjmv
S3RnD5GvIGBA9kYyxOiT2VDNIdnopJfEHWK3hjnn3q1FEuMv88fGva5MODnLsa+r
qbWzYyJCNNj9CD/YRGtFUpHJstUu5QwYTMgQXIXm38P+UvIgyYdztBhEExB83a2z
QVUODD4eT6cIB10O0/qlhPN9jeyfddq6s+h9HzHsrZH2ov5MsbWmzDSbemo+jhuP
7VSp2mm1z6sB6cuM7vii8EEG5j95Bn+LjaNVQ/eDm0aI95rUhgcC0lLq5D+mvfxA
jvWIc1iMS6rvLJUojSIte4U2hXovYzJAwqyZkzhfQRAYmF5liYehXMzput51TFxL
pS1EON9vwvp0welSfrN7raHWwIfQE27SOOGrPBQ0H1B7QnRCLLVJktfvCfXpy6cc
C3NJeD/dQVSoylcRaSdL9MDdU4SpFSWavMURqgsfe83tSOlsyEM9iv8EwpyxePDu
L8N/qLvmZLdH7k1B0AXb7kRrws+IdsoPC3B7r3PLVl4C6XebPHYx0wQ2n3LXdmfS
selGtWP5mAAUg1Xs8WTGmi+anaLN14pDE3IqYkFwU5awudGEPJY7qAE5+FkQ9WMv
AnBMM4RdzOJnxR0aE9X9Grk5bqw69S7wfpr8MLZK2rvPg8se3rM3DtmnzCSu/GkD
zjc/gpeNP6U2rye9b7kwG+ipRLv1s4lpe4sgPP+wwUF+1W3oBn4kPSzVPlaoihYz
a2omhiITBMh/oR0Xa9scHwQCu/Jwb5u+FVFXAn0eZqcl9iiAbcSPTNaYj7NINkg4
VBJWj7eWxgrXwaKB8ceyfecLqMbxQsiRdfgmOAbNxC4KZhECQu3QLWV0JiVgRILx
YiGhpwP77vB4m1HuRZlQIqLiHsdQLfOZdOS/T+7w2XQGIyeJZZKYtjGYCo+YmDzH
rGEcxzimwCYi4yojTuxTFrwRXo9clax183G4TAPq7EgaK1ihWs9cIgAG7riTokGn
kh2BwaaYJPbVvBP6YVGyJhQnom8q1oD2xyYyxEeqrq4LU2EXECohUnv2AgkfxsTw
5Ju7D0ByaEWh6qmvgJ/r/eVqeKObgzzyS8LYqAOoW2XKgpbafBAcXBskPDujIZY7
aX7vd8j1iIOFE9g+1yC2vg==
`protect END_PROTECTED
