`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfbWrQmpNe4a5LyVYhuYaGYkbZO3GB1L3/+pw4EaaTpQGyGyjOl/hG9BOu7FfmSS
aJinomTMgLVv4SGig0lsYI77WdqTmWKKm7K5Vd6YdpD7DFL46kYx8CRfmq0QvzB8
GBi6kCrTaWKDSLHwOEuu0iY6E7NqHP8GwL00JyGAvCYPyRsritGMiyfGx9Ht+DB2
iykmqFqVt65W42LJw5YgTuTMuoArR4zbh2a1SP6H+jhBEqr34joxNcin3I4DCri/
FznuP1QT/NIIbOcaMhXLSxNaz07ClK/zcZc5uQ4wDw02/JmQG0MVn3X5vGNykUbY
CSg/4rxVBYStItPFSgIMNsn51wVsrt9YrABPt/t5rU5w+/l8qo5MaaXw7Su0TwF3
jpL2bl/+QP9ME1M7EgFQ5Brt4MGvk90abeSCUxJ4hG63j/vXK6rojM856fHCK6Te
V5N9WwJfEK6xN0rJhEtCJdIYLX6uPxqGUqUEgkiK8lCI9IOhFpYQmvR8NYGEwgka
ueJTI5O9Nh5R3YVX88jt2a+7xADgT1O+5F/q1Gj9orInbRsVAefPh27vFFU0ku4c
jDVw2jA8yHjHPfzbRuolubw8HNEfJMTyYDOzbqFuWzXF4o1PWaFDnpRuVuXDxdtX
hfZ1C2VM3JIQyeT3JJdpQ+Ea+ZlPWRnc7IA3k2wEtT2GnlBrTIcq1COsB8ysVp5i
o+Ot4VkZss25fDbr5YweKkvpYf+OqAdvpzIbhTaRyiLzg4kNrgQuAFyCCXitI6QO
JYROHbvlJ/pnQo4B3suF6xnc6CC5aodT0F6xuQKRFK4jtP3j8wE4/F9LeIfSIDwl
`protect END_PROTECTED
