`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fO5SNcLgQpRnrskLkj256bU66bV2bK8mNKFxC34NhJJXT6SuX8XaX/dod+tVxYLJ
y33XYO7jTtQIYNg/SF1w0VrYwhLljeCVLXB1C72J1qrlhQez6PWhviY/z2ruG5gP
LG7Pc6etdtQx1kln2Vdyrik8kH2LyFf1wpvw2aj48GbF8hEtO96+hhD8uw0JNXsY
6R/MAR3esZByJ3Ew/0rWRCdLp/p7XZwCWV8pxb5a2rfIvuh76LuLl4WIkwWouT09
SgcNGQYd0489AVIVJSxBArnAy+LVd+QSTS9iKgVkq5ZKc4kLIwlLsPuLyc2N1yI2
cUqfswjP1kSFMnqpVOQNfVmn4mH1aBlb3XFHup18PemEJ06eLZvzPJfWa6T3H9sX
QvJrPdGKUiN+NpI4PdcyqrtKwLZH3KmZy1ts7t6jcSCKl7eA0q5iVj57yXnOkLij
3wBTm5JipYZGBEbQMjUaJSbBBOj6aCOyltkNfb0h22ufvt5hnaILdryFPX43UDMe
08jWMmArE6Py40EKQQ6+lVI3vCF+QqbxbSkcTmXl267m9pNkiyQYiYJ75dUfjkIr
xR0skA4FCgLF9GGVyBHU9iT+hoEwt25nYmV39TbSiLo3jAJfu4wzmlQPD/MHK4qU
cCtnh2lKVAtGxtdinSRR2/kZ8tW9KXkv7IEjbhfzP9ftFzZAgNkBJsItT20B6lF2
eF71MlZrH7VQj14+XJ2SaOQ8fB2Amt15rXDAcpuCIl/wU2QIPdvMQzJbe30FnPax
7YTd6CZNyUKzj5kVk4bJHEb3A4cQUyWby5dxghF3DqCLX7yAKlpvtV695CuYjxP2
l4drH5CnDBQGQwDOwHmjYLoAnaI2vb6SBhaaMezKwFxifMg+cTPsg6OBX+He53aX
HJaUhZz/rfmD9vo5H7monWABzyPj1Xj1tbKW69cRxmJ4JtV/AQjFYecqE4mCRuMm
qlDKq3g/S/SD5KYQXCUpFEdaEOf7TQ/wKBlYfXa8N7pn2yp64vJ6RgfhwUZtcbBg
cyA9MGoNtd8cEBcDrSj3jKt/QkZaURJoSzSAjVYsi+fGfS3rRZ0+f/bpfvr2aWa2
fPg8Khn4Bm0okJc0xzWimVWiN954SvMo8v9p2Itjvn1MG/gWbGTJ5Wn38/RU/7LJ
5jAHc7Nm0ALmaU5bF+ez10DdUYpK9mDSLbSDsqT0zf8zl2DU3YA1Hn8Rh8W39b4P
`protect END_PROTECTED
