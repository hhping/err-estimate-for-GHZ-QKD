`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLk0YWbj7V7t6n3fYlNBCE9rNHLVWPW/y21Ah41DtjTFuJZV1r9KcExqQCvZ/X9X
ulT8o9ZfVRvLamGWlNBpWdIXF6miF/HUH4C8k2gl6sRjq+LLAt9qF73EBDQgj1ed
Z7mH1ZAYukHmfX3FV6SHpnCTM5+7CAWSFyzP9tqL2ack4+o33JhAImss2aTiW4ZF
F2mDZYjc+9nrMR0cDDU3tbGSa1LM7zFy4lqeCHUtc45S/6mdh4qxkOT1FZQJPLeu
37GL53PBmwl0qwOzDjWhaCZW+62L4Z1Avu6GNG7XUr5MPUl7QltdDhYPp7TwQOlY
Sw8aQP1qcNcu+fROHZK2SNfgz6ykFquoeEPM7WZqSZeR0FJruZe0A+wDOeRKsMIa
3f6JlsOOadR/z8A87afiieFEkZa+2CT0A9PFwKZNzkA3ailQldDOfZC5KfJ2Qpj8
AFlLogJdQ4WO2rSu04VCuI7q1QHXEZwO0fDZY/FygVA5LHpooQHKGN91a7mS9wpQ
6TMSUs6MS5SdXlQr8TbcYr8rQ13q9yxbunA+oivUl6kRPNzILfVLOHAhvrmIl4HS
OmeJOgoLFKPXaRbHxHzsFhTfpPU/HDNDsvoQEXAQwC46ufdX0R/WlW6Sey0bv/99
GoXOGMl7UI4hMO1heMIuKcPi9vR6lninnuXsuI/epSdMvJ0P3uOIUPksKf0ht28U
UX2TeyaMNECrQUsNyguWtxQJ5XZiXe+iTxGfOJcaEeDGkK89JURnM/dn64Qaqctr
zKSAkQrP7CuQZeypOjWQT4as2bVw/BA1VwUEqmfoJFDlN+H4L2sb3KX2/evw4cDj
mJBU4Mx9/ln5EAOsieoEXHM3Bcvt41pvcZMVoDObXVi1SBOdY7XgGBRpIiJl8A/b
cKDqLUkPJYjSFW5ALc25v31LJiwAFW1n4GWwud7b8U8z5wFqPP7A+4uDwFGq5jtK
23CDeh2KBSRFHLStv+4A6JVQRhfT8zfzIxkgaMtpK05XIGIjkr0Gpr2WhVfUOKzT
dS9LsruFgIOyHm/6UI4FzXYhmV05syCWPG0c4tu/EEsMM0xaq+RWufUScxwZKNRT
`protect END_PROTECTED
