`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDix8GdWQ4m9QFiVQc/ptXT6QdGHHB5O3QBagH+Y9K3xHJEufJUFIRaIA4pZBkRr
afKv1/TENnXdY9SapOVZner+eIIltoCAtgnJReCKXvlaFctlaDC9DRSf3esXEsDD
4kBuVzC7Z59jwtKJI7Yq5xUW5pw+7VxhrkcnLcaD3snLW2eo4ohER3uEeizp1U2z
s7VypMFrDXpptF41cv8cABo4/mVTRcGlAE6/DKCpVYj55xZuU9DNI4cxGCrWT+WX
Lk3xDmMAPjbXbuatWQd9S2P16rwGG7RtX0Lqn6MSmJ0zyyuZwM6tGHz1tpXFaa0A
08tikXzwYFWbxd4WpjcLI8C6mYHWh7wg1SoUOPgYmQEnlUA6H33Mm1pxxBwSxe18
`protect END_PROTECTED
