`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kOJKpe1Ea+PzbALuisoZdd9XZCsiV+8uOEZAjQWFf84oDLGp25pdtZXmPE4NRLBz
CeKtrIpoMqTWZcCx4UVQ+UFt2odI76Ie8IG2H2nOh6xhh/WHQO34oJoczv5vY3Nv
LFAr5ZuQGjVQMEDn1GguOJzOkk+UWLotthAGlj0nIGdXkITnKK7VhmGahZdgWJQJ
A5gTEcHK0wDltPYbw/P59qHjh9Y16qXlHAUHet82y+bpg38SR7Us5Q3DuGnEOttz
xzWq8fxfEqx22Y2g09DYN5OxBlGPpvryZXH2UKYkx86+3r+Gq0VSApSOxJts5U44
x1ZG3LSy87w6oMoPKNd5qTZLTafjvg4E7izA2t0fcZJDwd+MBI+uT2XMcIiP7FFX
5V+oJ9xIFNz5r3USpEJhOlJghZxRCal8XEosH3jPytndkEX7unsbR7sBYi4Cm0YK
3XXYm/dKH3eOhh0tewqst4FTFFRivDU4Y+3dXQZB5PuhD82tqkcADIpLKAAipp2z
mWeTMT+aBWTBy2s/PGo4Ghj+i5K8Xa/fPwLfZUhgAeyJrWSfqC9ku1J7sYcAJ6W0
`protect END_PROTECTED
