`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47oiRbxFi7lH0rzIEGAMxeFs7Ueet0ZSIQbTdRJ9LQVZ9T9Q0D4nzgAwk+2FYUpf
yiP8tosNpDqkzX0HHzRV9sFtz9kpJm81E20mk4TOockEJ4uvGvXU9AdLvkURmriq
LFBALXRDYDBbeO8ruhfeqP6ytS/ukcOWjmzQP6WMuTO7U5yUI7/0lUC3nxBA3GKF
+WLDYez8fAGwb6MoaU/znAl8+EaWcE5V2ooZxILZi9lxdkFl138BJ6Y/adrz90FI
+sSiLtQ4nSvRTKsu+/HbMaJHgQVW7Zh87hVaAHGnLk5DnTRsaMksgR/ClGW6wlO2
HdPzwWieSZIFLTlBe1AA0/S2OJJ4nHt04IkVvAnRmMIVnbwiJl5O64OIci4Pl+gU
FTcgWRm2rovSOf+xlDGWmv+3VIvVnOER3voBazheqa3BrQfX+DYV7mYsbMmsduV5
ASBxj+K4HxXqs/2F8Ukbt3gcFNTTpPwPYQkPYVKOAGTh8lt02yHd4FUUFG3V40UB
oF2FqOFH/4oS63uSeyMvy/d2hsY9pxgftHwBEl8bpyR8CkJasoAzVA3eecpYjJ2Q
fcqFVXjhRlA5PnrudXtR13bl5jOtGUPt40tA4mSLip9Oc05JA8pFvQYCOR74+YtM
4XZ+VGTYO4YHIkqLYTuPT5/taL9qqHdYqsxXywAvC0caKpziko4I+4CGLfYpwKXQ
0kuicOk2QmST5sr/ffFbbyg4g+O66y5NLookjPys95xBcZPCOO5oflfbTh8/ZIEe
us/8WYqs0i4deNmdiz6OmwDmJ7GUnz5K/1Xth72ld0TYnUudtwdg7xhmcw3+1ugY
scF/tRSEk1X5+4lIhwO/RiWBgAPohg/nD9rpwDF4uWwKA22nx+vEfs/ZDta0uviX
uXS+ZuGh3S2v25JPAKLrx5QFCN3tXUFFwNefhRnb7eB2vwIhxL1lsGGtNnsuiLAq
O4L+w7i0Bnh1XshI2ZeH3yMvNEuY4vrbXAwGpzJxlu4rS/VNXuXjQEqgbD0zt+Wp
YqPMvEqzavr7one2eA9TCC/69JaupKUd38Ido3sMZeGNbCl7nU3cPPyGoHDtsZPL
DFNRZu+RJXzCHA1jEVlm1qMQMoIi7Sa2HBbjUAEB1H3cQ+4/ELpzo0Gkb6DkkelQ
PWFAzJCpZgNo2noBBzyoinG5RIRgP6z2kfe3J/gfR9uTqvbIifCWH7witZfWtvWG
j8edoOUvuKgYe8ti2k0HrnAQqVr+pg8MKHdymUfBq8pMCEAM9ttyBw3hSg0I/Ffs
n71Ph6sQwtxnOEjH4+HHvpDyq1lgwsCWrb+eZ1OQVKKcR3xwkzne8AmmUjExM85U
3zyBBNfvnSuFUIjDRyCvqR0ZxDvO4HPETqFeoc0/nBcnUc0J07yzvegP3MtnR49y
L9CSbXCK94m0Cp4pNhuucibs2K1SQ564A7LGAbMt98q1FKX4DrN1el4woCYi5e8B
/HxTu1evhT/qPzWNoeMXkitsATNSMHzXiHPzL4ZTQFMpb8AwVjo8Xk/UP09lzKQ9
Qj6QAOTK59/dM2py6EmEbLnXYPXB9iWFw/n0SqPDZO5LyZAsQbW1ieKHc7H8zTMA
SE0lEKfVFtQbeLbYT4wGWRX3+WB3u/yFcraCabhQ/kSWR7DeHNG+8/vdkoaorChG
8z6grKKUoo5/9j/Iu+M9n2z9RAA4QF3zvDPv+A14JZneJoMUR7KrdYegNTaTckuw
NhXWx+egbtnlapFF0hlJu9WHeaV7m6MYKIae5OZx+f8=
`protect END_PROTECTED
