`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCrM7pec9012h2PKQXkho2GoieTdOTWKbZ5scVLEK73jCvc3KOZjkU/WfJBbmSNc
J8TUFIdesWx+s/GHP2YkU4OZxGhq8d1BhCVOrQ5IVsYEIskOw3eMeBUGZ0T3V0uj
dzicxz6HAf0Cd4ne9bRVFiRUGdX3B/NGkemy17+pvgLGZf2UXqT3QJJbBTklDYIi
WZ0wh9RLUEiG6jFsjwYWQQWLB7XbnBGDeyC2ER0kxDnEiT1zo8+AdBTyERHlhA4r
z9Wk/AEULRyVcLnDBFDJg+jIb4AReJl0QmD3qn/veeuJaEsx+4yPog3QzfbB+ade
mIztAWydOvhzrGwdWyh28h7hn7ppBDapvszaXK0i6Tc2yilsu+wFPmgWdSv2q53+
x5dyd/H1d0OF2ar5vue6w+n9SHl4LiKkzaGrFKGmZ3ajGaiB2MclYZkIUqclINw9
qBSzfE9nTGz0iO5cz1GVVjFOwifG8lHN0VlCRruFccNJyF4x6dix00ZkyZy3zarT
FTT/mi2amWGyKvA6SqG0E827yDW1CaLPgGIeump5DiK4XXvuR4Itpi+dJLeEpE7f
AGSsqmCs9xRN6QuEZY+U9Z35HqI377vwKI+eySgnv+jiIvkYxVMthbU5NQyEZeu2
PBsX5lriYw92MJK9BiGjaUfKPh/gC6THkfAXkxS5BYOvBG2nmLbtC0aObGUfxjfv
dG7cOJBYdu8ztSsyBvfRFTfWtbzXTfaPsuZRctIDPesiVYiyQ8tcY9tZFLVc69q0
CUnt1yx/T3LpUFBJfn4DLPhpIRUqcpUT0S9Feejlm/IbB8yo3U3saiuVlBNVsiyG
qE8W06yUCu7RJRt6jb+CRQzTV3E26T+yGug+1sj7pYACSv+mrv3N+OqkCIVtpLlB
xWBMgXn8f8Y2sYRIhrj4p3ojHA1KJ0mO/y+nAWcASYfA3YMKhYFTUmmuJt3NCJ1F
W2HXpeQYM5Xn5Y69KAcCLDmT8BWlCJtJ7cYjxg+PUJqHCQj02OYE1oOHZPq3MnV6
JC9DiShrtkXio8XuRDm5M2dcCsaeXiow43JyLKmUj+zKU2UZ2TUXekGYGjpWk72P
GQUoOooAdFdx1W5MOVKZOrOYtoCJea0qgAnlo53Gh1967b98uWNULrEv9IT1r2U7
Z5P6dPTVp0UG33whdawypJl6JbArfDXMwz0CtYseITaUQKz3JUCrjWMotONBJjYA
fpx/0aXXRhdmIFU0bOvU2dRmvtaDA3yDp+KMgHceCWn/XfalEH9qT+xVDTqbKifI
1cTeg0hoe5kTZK7t0Dq9FsMFMTqvWI5CDb0Xpo8nChGHQx4gXQZk9eHwg3YUxsyw
OPH+qHitgVvIliAQOU3zoUR7ympS93sIyTJw/0VNXTCjtcsMh9VXJK4QtUV2m0M1
duRpwGh1TmLEYF2CIC2aHggiyI+uZur4ilgM7ugNb3/6fptNERNWZjnqjj/gqAIB
1KxlZixFxAHIv+pVGNK5hQil8BsqGmceOaQx58H6ydGXVjHWoOlV50jSLcPFDWfF
1B4DhHWqS5nYiskQN9oVJDSlR/gyHWvkw+WLQYSnsOyS89lmFA7rdgJUX+jtyGVq
xdBvY27Z/LDmcLa/NMJsKKDktdt85iIgNAFq+McRz07FwvR2kUw72MHsWGzWT//0
BbWTorOINzUy37fYaGpP7qCZPhSm3V6/SyKvW4p4RXXzfzhHex5suSeQVhy0WN0k
WuI2yXqLTmutx1NZg4i1ay/pjdraShCX4AbyakMdWr7Mn29/7QlaAmQi8zt9xGDi
`protect END_PROTECTED
