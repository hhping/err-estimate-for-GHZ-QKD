`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsqNtZTGh9f5ci9qUUKl9HOnltHlKMjpPa/RHzxh6dDZ0qtpAZ5kytdEJMe+9tCM
Zq9NfREJAgIATztoCePZYBwloEbUjv8+WlL4w4wvpyb1lea7O8gkHMa3FJf0C4BB
UIkV5LKzsyc9Vza9rgmoRjvJawDDQUqFwBBKYZLpCBpyTglp7PzNq06xf4TMc7Rh
1hgTuefqRP60TEgKLniC6CI2pNvszMzHAtDM750bcRZ8UGeekRiv13ign3Rk2Y5j
wM835MLaK5hW8a6RNZ42tsQ1qfr6BJZhJOY/SFjkxgtndPBPQlf2VI4q94UQuRrC
G5naT8IW4w2eQM6o5uD8Vq/EeTbbv/QwvZMRp40ox/urLiG3cRq+1zgYmTH+oq3f
RaQZBLtn2P1mmPfAW2pu/U9EzQx4olZ41PfkvjdUrWhkfTJeNaZTN237W8y+V73c
M+yH0q8TrlpujY0lJlFul8o1liQyaPJlzbKbAkXeAoADzkAUUtuHEdkHAFDYmGk2
joapm2nBoSIOWJL11oXFcv49CGjJ6w59Ry5NvkFTW1BnXDzz1GXBwtg1O9aFAq1y
QJsyANFJZ6bGSYaD0xPoUQJH7exnv5kRaTjFyyjcgK8JtE5EY6AYmjdV/KKTakRs
ydZwINrbR1nSKOaZkr0nUlaLdtLjU05CE/cyyuMtVXCN3T+K1PhMlMMr1EejKk2x
1enTDJO4bNxta41b3fZIDne6MRjSQOdryMjV9kQR4uQ4vHaGWdYYrvEC6E0FKvoN
i9sKd7DoXVffWyMNu/9kTCyY7gYkwi4pPzqL1KGBN8Jt0gVirQoYsc8yoq4Xs7p9
`protect END_PROTECTED
