`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XxQ0hEkcVsxu21f2SDuA721mzOK6MF4nb/CZ52JuRb5hGv+yC2WPJncevOcNxRWS
Jnw5PZjc9cClLx6IazFaJKQMAcV2HbNT8QADN9FdPc1knK9Mj5aNpRpNYx3zfYT2
bmozcjFWekayEkRaoyWazD65ay/wTXbuCy8LoaO5UmBoyArUcGNNe5jImVz9bLOA
/TpewtrPGWYPHzZRvxMzZ2Cpiw56y3Y88MyJxaQZ0NxHwGIJl9oj/3X1xy1xAn6j
Ht77j4olyKaOqaTpq+YwMXir7F2sqj/kPu3pSjUbmiCOtUQXHgZLATmEjVuSDTOV
NEWHN6IaXBY2FnZYfTbeiqkQPU6KltkPro3bIg1qusCc/eTzFAAmy2zXAbtdZPO8
SYwSnl+9l/+YfQ6SWclsmiZAuWuTfezpi5C0fCTotC/crvhOgUNZhEgwPHMQq1/V
lJf+HbR0IbVmBo3UG93PRNjIhU/BBW/2XHBKGLhYIon7hjmjLA9F9bbCqnDi0elF
yNjCIQe/mOo0oBVGO0D70aYniuhvi8XHrAtUzjyyCXAp1h5A7XqrDrVqeX3RkYrS
Xpq913U0R9MYKTKPeB0+lx/qGCW+CN1YkPBZKHcd42mQIvl1e2BHG+9gtxboUCK9
iKZqRYKZk1c0wtH7vd1f8XyfiuhIoYvDE/u3oDQGStCPDh5G9zDjlyC+oml5donI
66AQV05OhzpClOZfz049dE16BoGCmOoiTWf0gaNK63J0aQTc4HLvyzCcb/VMMiB6
xD63EVINMq/MWW0kpI+4DDZZQfRcB80QrrnVBe9ak4lkmbRjNjwL3RREg3+Dpa/A
6p/qILhvyQmxobdyw8szime2D8yQyKpLfwc2bXcQ54yBTd8spk3Sjleq817QP2Va
K6leOHYNCrkD35eEcZ/A6HTQ9GtNZM6XdWs0UWOLHibXzUBXFdaB8WL1RI4QULXo
ceZQzZ0+IaOMxc2jFYkttFp9v/K/aHTk3ARgffIR6WTyRLq9WFFP23gTf1tH6/vc
mLfl74nXamqz+RGNIIIeRnAjkqks5Hg3MlNMZobyC8pxBQwdPJsATX5nN5MvjIsK
lhAfCbFpbbMyUaP6zGaYKUFWSW4P9cTN6SlXfNR6iEQgVOOcDNyaGc2qym48TRwx
VdRtw3V/yhjpmeiEQNZTEFQfnojWaosaVnfbFiZTFgZGD6aa+ZsklGZIkm3g43qY
fj+ItLl2a6cDmOrJFzreCCmM+R5xkNfkhkYeeIQPCqGCO1coKZP0rGgwOI01z4dS
jXa9EQybaCqeWCA1UzqqTU3Z6ML7JvIiauI3tRDifsZ/ihdezjZgZ+34C1OmISt7
ZTNvLSZMIDfIigrxA5C0IIW350j/AXC9wiZ1P7ZAW5m3DWtFB5OSTQ0CXAHE5zI8
qnD4QyWhmC+oO3/NcN4lf+3nMucetSdS2GF0WsmbZYjW4jbgccjSVgGx3nBh4mxM
D2CYrOTe7vDloAdRk8TUSS63j6jtgXYQtljj+z62InMcASrgLWB8bVeyOkf4lSFu
fkpQDEaQuNGr+59INwvTlK+wySK0p6Lt2EdJX5oPXW4=
`protect END_PROTECTED
