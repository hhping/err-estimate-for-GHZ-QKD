`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3kfn97cXce4SjeC7CPNh62SSl3hmr6aFU7+QJywJnktXw3z87ZdCO7XoDA034sN
FKpQR1u6hQCFI4hwF0LUe979r5qRXFIqekkz2cyTjNGK2dtapGQ/OaICsPnowMpz
iZYKR3SS5029eKpxQ29agPpaM1DaLGWaX4fPULwJiiGVSoMG3+kh9wpelDNeOhC6
gVc0/f3p97p8VY+ahoGu6mJpV+VYCqgDPqru9+1MVnyzX9dFdcRJn7oA+/WN0oOy
pM4cXYKwD339sB8qAGvBtPmLG2cl0+qoam39AYBhmHzsswGiKXCtWK33KgfjPPAz
lYzEBQe6HBQ5wtXJZHp6moJa4a1VT7NLl5DU5/Ublu+GW9/VVLWBq2kEPWCNZilU
H3YWyoK0Ks6pdNu6pDEZbAfFmm3sG3xIdmohxkr+oGoSfKDxBy5g9mgRZn02CG4k
G2NJqQV7jevzQhketahlIbm2FhZmntVGMrCqZeZ1gn+HOV1vp2tfKFIIz0h9Eqpa
+QRnfwYUrqchCxvGsBRJlJzaZC9qZu/2Jfi/4Y7ha19Oy8TnxDf+4X3C1xkifZKN
kCeoIZ89tDzR8UxAtFxQyZ9/6I3WXQzpIREtJtNXHIMrA8cS29Eg7lgz6ZCUBmJn
xdpIpWW22wHO0KI9IE6PsOABpdX1M2Lv2CAlZYma2Bd/CiryiJkOH8hhh2oFoWwA
rR+93LPzUb/+vKOCidJ/EeVVepm89v3gR8JDbL9ghd32URe6tRHFdOlb4uzFPDDH
lUugT5ucNumJ3Rr+ZJ4MXtJ8WyqKlELeIZcPcbFGevxBWpCrFnX7IbJIkLXuaB80
4sSjOxH+KAZrLDXTks1iIiMzePQi5995PsE7mtMpj3jkB9o3/+zqn/iZDg7SPigV
lqxdUS0SlmFqy+KTRLtkfLooZBUad2YW/9zcaDLDsafDMz4nIeFM6HIWPMriBuTy
a20W2r7u7lPE0QHb1QTPQ9Uvkne6mQle1ec6I6N+VqCNq3F6qBvnrWfFVMJsy+S9
CsaQ/xpt34Lx1X2dfjjHfEjV5vevyw/iiF/794AoXqsK4J0GXGdOn2TqiymETH4L
Uyvp1l/i4dYWU3tWfc/5HPvdE0DiE+p9u9OzsaZ6ZRYeqWqQEqUmDppcJCd4Yarw
UrSGt6Vho/qRcD9BDnXCz/nhskcba7Wq1wbjaYjeKtcea6t1YlglTXnC8QH2CWhh
Jmr98MuH7PseltLdoy1NCQ+1R2wkRiNA1vc5mBHgndpbE2CaTTkOtdLO9l0DyXEH
PzuJLCjl9U4XJEDw+LvTAZJL6fEnwQggrIZ1dCH7Q52yj0HJPBV06Aa2z3Plbr+H
8VjSnfbZiizi5Es9IIk+0TAF9py7NIW1QPIOmBvxwugJBxaBY2HkKMsUAMh4l8x4
26LX5+iFdr4ncw3YRK5SULMTpiF7MtE7OlC/YMPhsJcB5xc3igNXnPxf+PQ/z9nO
Sl5I2X8Mn/j8EDG9l2j6QqJ0/+cMVWvteFbMFWm7MJivmZdr1qq1oeoWDrCEYvIV
XUC3IZEPtfWuMPiJF5rQ30owWvSYqnDjGYkLmBrExU6SEHG3UzgIPVRgX+FuJ9d5
AHlhyO+StfEXSQma9vdcdrUXHyMz0JLHYM6XvNsK+zNiSXCZPI2Q1saZbbdRQgUu
LZgaNPrFs9LoacPXW98nOteZWNTICsQw9WTDUy9UTVGIAyQ8A1Sy4x9ZU2Fnb/Pl
fqYRObD32yoHsXWRRviRzwW4TJqZkaUNrbgMYi19kHR8Tvm8+vOMVbZakYu2VKWC
ocgdLCAo1Yv9kkxx2169ZHD9JCLWGhpxKJBv0IvLzrWjKDNhAGXkdxA0nXM+GRMm
L6dmZoySLdQQzHcwiaSaVIzUp+wc5crQGGt+/PGJPjqZ8ae9ywWhNiz0ZIt0V3wc
Aq2f0LMeH+ZlSS9SCP2kI8W5wMV86TYxlOv9AMnYn/LwVLlI6GUCI9gRaxeubCOO
PqHvI5PGCd/kdetg8TWP2GLgi7Gyp4qlZRRZLloeZmIlu/JqEEMTwZU4IWeoLn3c
RUoVijV/5AlUL7iE2v6RQCGWUFKBZrBHivaMC5g58J4tKxh/Q86KU8VebhMo7da1
ntJp/jZacswCpAup+ifYCw7/CFJCowK7WDLTEPMYHRY58hFtKD2vpkeAerutOgDS
sD3rGfOT+/isAFwgYNk+rVK1JKxcHHmpJiQYO9U4Kh9IpzMi1AS9sFlom9iqTOoB
cEai1oC0Kth5z1PBzxpxyHZCja4qr+J4E0qORUawrxB5Rws0iWDLkaxXTFRCfP9t
mAiG6tY4kMeygHCU5/kXnI1mQfAA4/sGcwr9lgb3U8Ody7PbfFanVIvrto9h8NhF
wqZrPh3zhh/HJTOLDjJfxdhm2Pl/WHxpgaCL6at/j50CD8QCEe4xMI+2r8zRRh9k
Xzgh5YJkYot+17Vz5Mexk8dkR2NmSYxCa8ahkf1vAs8GUaObMDm/Ery5+YzPak0/
6Yfh4e9kGJpmyuM9ll6T+7y8c8XocNceJJNwKQI7ly5zC1qY/izLeOyLB7dBjuxj
Huqg/OXaa0PshL0XI75inueBkEfFaPZFHEpNJXSDVXC2zeHxUrtYgbmbDwEx2QYA
JxwMCa8infrsXmtn1l2UwUKGQyxaYnnBAw7wiRf9gpjkc6d4IOQioq26b6NVgosg
EnUUbOlYcMsQ2FPh64cqW1IsvvdKf+Cys6O7z4dHSylifloaQ3PWs0YpRwxL+cY2
Pij2xpqdTuAdaD6DaK+RbmI4TqeIDPKjDgI9mQ7+IaVRZZmV3ER8zO7yzjcs74hN
U4u3OS6ZsJgboKbjL2wfOVXlvj67LKrcGapL8kO9/xB9zutNJrXIGegkAn2lL4Yu
FoEnLSt6lpGc6qfZEFDHXZnXsBELVf+pe4Yc7G5nFk0Qse2idI4SKHvrgvGC86G5
mqMkvCvmJinyRSO34MyjVhFuwkaehq9Pajdzsn8rZr3s2XhOG4+uN9cqIyXsE/06
h26CsUvXLoRXNrPoAPnzrn0+/1uFELx/WAegUh+8+M2Vmum4xNq/mKooyKjp+Ick
hZJcnKvphEbk4tnnXZAncDfaXv3u1Cf+81o8Ibl8yVsABqWp3B0KLr8/uahEYhAp
gahkzCGeNuqD0vXHah49e6G7iTYPV4p1y7sdr3mZaEjH6MCJxwlXnNNxCKX9LTE+
EzfYXiilLli14gLj0R9Cp92RC6ADW2TyRrPEExkeHPiKpcnwCNjG/4r4ou+ktl6u
q5Spj2JF43f8NqseCkKeBKMdBhdfbGzxybBpFgIkAbmJEdykmAuIo3AwOInBTHCl
VTMfRM6rNLs4LHEfL8DoQZJBK5dB0ZOC3Ln7cN49cbtQU3nqQsLgCCDhza+y4uo+
yIGIIO2sFKVPJCfa4/ke0Hvdku/c0nyYpoXrDXvsFH/grdpBW7xala3uABj9LMwd
lWX8C53Ty8anVFnQ2JpZULnKydUEel7bN1mDG5LpO8T0A4m0WxEOr+trJNjcCy2R
pFa1PjWggQ/AIjJZXTu1ZryP4olStVMd+V/iHoL64c7Jr55QIsernIWKo1hY0cGQ
N9qCKgIQ95x8G2NWEDGm3uZVJn+9norb7jEKOokRqqTvdT90PzNHmxCv0FTE1pCS
fn/zv0j9IGGlIsGtvzFLQlcK8YKdj2mc+D8Q8VgjA4V9p2r2vQQVrj2+0RZNVEU5
hwICf0+emYch007N9v+XlZ89w/Z7esQKkwjx2eO/Gs8Ae5C+XAm3TXkeSA27K+Vu
hHcBedoVRAV4lJO6Zolsmd+hQPw/ul6nwyEOTuwYPaBrjZxuokCJ3uDIumC3GSBK
wTy8RQqP0Xrwe4pg9+955cgdMdz1ayx1WfSIxbZNZ3QV66XpEG264mbKo8J7zW9i
W7FAvqFQZnvBfHk0RS4K8o9mP9A4vGNiyM/2denyOZtlMGS5qcBugWEcMlIPph11
DXMM1SqxWcbE9a9THRUzYh1+ch5nYK0XQFkqS36SkTLniAWJJNDqyAKmSQ5e3Cwy
17A+a+/UPV/pEBqJLDMH8LQFEkt0psofmSzGpMRjLYXuwzaV3FOYDr9F4mqyrCG6
z8B3nJmCSB1R8FoCt2ZxgaemECB+IYdCcAQzPW9MLTWIldNnyqLj4KmBXjFh+N8q
P1uw17Sd1xlhUAO3509hL17p22W3+bBfPk1ombhC5vTvE/Zh8jYsUrS/zG9/jmBV
81uv2BUH7s7/dLHspF/PbvvIQ3OiUynhpKE4u0HU4xywShI4QdL08KB+4sGuesPF
BbrndScH+ueXMfpEfl//lkt5IEDIe+WBhkQl/D5ikp2CNAJBhNN4dui1dF9zfphq
JgBsXWxRwoJH8TzHyfAswGHCRPHb8ilC5fYxLcWVq1nv9PgEbXubRl1FyqL9kUrJ
WBjzkChQf5F1vVdXajXD/cOtBjZxMhXZTlLcFtmkZRPDHvIfuTHw4DfF4wUyxoix
DaBVWyabp4bgt6vvn6N4IGgqj4XKESjCkvwVapP3mmhfW1JMUFXEUU9BwRLkJjxr
WKEyUOQE8fXxhFp2zx7x7DrnPqjBTVsGp1pELovlunCfKZrZCrj9tJKGx2NF2Oub
5Ufm0Zp6ZJbXFXbxqXU4Rl3YWeA5UVny0/wjWISKzhCiHy/JmtiNK++QIJAt2cDY
2uK/HpTuIqBLr2GscX4YKVfPDfIBcNaMOZRy33TtEaOnBSIMh5FbuJtZAC2ztijm
0LVTXWtDaR2vgskaSWEEcmcSMw/ZbTh9jU1vc5dPkm2r7qnCK3jbNJFL4sawogQa
aAqE1oNeKPe/+lnSrYTZ4s45xtmOotOYRvm4sVWKxljyIAy1RHeuf9Od0nwZsokO
JTmqkBLY55jyJWNvy/+vzf84l7hly9T7CT+XHErc8Bx+fKl6RmqApHS4HPSeMe/9
BBZDFOD6TK4gt3MP0bLl2fvehiYjl8k5h7OXN/X93W46PtcsVXV7nSwZ74GEET0b
aL2eUanVcluavRVga7L6ojEY/9PVH+5Z1hwE3zEjRypVA7ypauHA4FO72ZTRl6Jj
6G0WkDO9qujPUneLNdyxaTXft/MqTeFRW/DQ7CxlKH8tvNljWtul4PVwgA0OTPzb
WgpcCMaEecSOmNCqoWYKKS6Hxiik1/PxS4MadIwzOM9Sc9omhBzjG7i/4OmMwARl
fobJlIEd5cb+vB4BAClVWvwPa+LWiVwMc5HoFvACH0NWaHVnEBC68PcW+66NhR8D
Fo+D1NW86issgUMi5ZNu2Ukdnwzw1ro/wOF/7rhZeFBgNVta3RvesLYAFgZLcQ1l
phb4Ziu/QJZ0M+zOZbWJFzLgi8swFgtLN0yBz/6IJj29kGAIX+S/AQr9VMA7tdKK
iPRWVD/IOZsYUljBNWjkPu/RpsbI3fg2WMcRsroRHsAYL3M/XpKjvMZHQK4+O+gX
CQHnIQQPYWELbzJQ70qlIxFo1Yx8jmtdTX0QOrOfUd+EgPxRGiyPB7L4xDK3AKYE
DITMRzBNv4m4nFAA+FAkhkHcl0X/ioRXxIL4qhX6mc66FYGiLmP1VEmjpcr7/gKw
cHtqAZJToqmgVqz3oPlL6iQsLDHwM0lOLKaRxcn/ycCi2AkNYA5wISneYGUJajut
M4eNM9tLhPHUtKNbZFCAc3KhvrSZP6uAx7P0ryMnik7B+7sY6r2ip55Ai5mWR/W+
5CTSlxqo+9b8xxtYjkox7RtLMjVt9vSqgUqWhdzL0VWg3y6ooHhe7n7b3pOB1sFP
ymHvTxjiY1zIDZqrx+0o9eGyKydrQ68ArNfThL7ChZLTkbm4RnB5K5xx/E2o/qEQ
tVY5GcdDYdfIjfh9xGq+EhSXR4p+zMt6CMJprkcMQedrnS9jQKik7QM1LSCBVCNr
iisEYxKLlnlJMeZzc+yZnubWqJJTol3Xj8vZsziL84zWTDIrFeWuQpCzHh5wUW1s
JHYWDXrD4FD0l7f6EpFetZ1bnRGkkkeLn11MZ8SYdeojOhf4uYli47ei2rFbJfDO
w208jDnKxCIUFlSLLzSvBprzbyYE/XSTYxU9Iu4uy87QURwolG+WiPhOYE0UNfBU
IydFkWgPwA/9L+X3ZdaQED98UOWOJwGABn712QZqkIkeOm+DIHlyFf5xWcP8lE6a
SOGOSuwRjC3aww6l24S/XoghYQb6L4a1kqrbrTKh0sj05QSg5cdt8rXG9zZd5dkd
tGOwelem1aC6IObhoB2ziMwdD47hGVtseuZHh+qoGZqLOb9LFQfQ4j7XFI5GI8Tp
VfZxnkSoXZuxVXaJckE+cwK14qBXO4gRFEOfS5H9KuTvwHz2CQw5KPWdaWfEeZAi
4q5jMZTVB5LHX7jfOBizEsYbAI5awN7HOTACvtxpqiPMACV31CXJhVZmmRJzB4j0
tabZoHgkqO8ikm3q4w9G8ykdFAQBwEWvyDSFKGv7J7QA50csUK/JAhE1iuYDnf6N
0Lpkj0yMQQ1SzBLb2/HstD08ZCFlu8N35SmZfDWS3FvhNKvc+s4XiG0prl/Y6V3V
Hp4N3WWyKtBn/WHBQE0AxWm1KRy1zn/0HrZQxpsUgrHUM+lmUhGhbvjDEQeGaFKD
j2t7LZFhu4RU0pto6l5tzwmwx4FSCAq7vNSXCA+AHlsGRg9uIH5F9Mn4uBy7W9uq
siomD+nm5Wo6la6MSaGoeCP2TEGzai1LyOcA8jB7mkHQNJDarKuz6YhXiMkBBdiJ
ydNoWjkxmDhhEqPbIv3VbJUcmUUOTIjt6JBRFAa5YZztec1wdRqlnIsNbYZTmwWK
pVswdk4mPJbdN3Rbf6VAmhPty2P/NrN7aYxYNFCp1J+NPb4C/5uH9FOGOXrIQSDl
Yt1DpwBYtrHv75Mw4f2ExoVoew42N08HxAIWX8CJBI5I4yi33+WtO27S+8GiKTab
CZqKaoDCS7A0LQkTK7g7uivg+NzuUtp/t8mPF4s8hr3OEIrWCAeyqT1l5ZEptHVh
nhDK7wqtLPUM+kZ39B2e32mmSvKzcaquhqdiNVmZvfzlXeoPF+5r9uTOnzlAG/5h
k8MMSqMt6jRoco0dCj7U/9j//ev6yppbCrJx3wG4q9FNDqv+EwL9pKd934hsTSFQ
GjFyXSlcJW0tm5dfeQBbfpwE7LJUa55t0EAB8QAAQAIifk8YoYtjZiTdltSJhNjb
OFc/Zz0ubD3ADN1xCN+AKu+8NR/09G9UPchXdvqRJYROcjFiRCF0CXWXij1/kYdK
MjCqFId7GUQJq1KsNa6pzchkQOERW00uvu+8DKyVsJItmJ9oJVvsIKHGFkEyF9wG
OK/u59wkX/J+8UBW75Pm0pWphE3CKP5w9JfumMJ60TO/sbuy8yzIkUv0FYgpcUY1
+uw1/n7F5QqEc77mFCP1ZgStn/ankL1AOhnWjxV3ofS7DVQh7cAInj3+tgSMkH4c
nwNLDOjIjNRWUQxgQa7NIqDRVlNg/cHt/Owz9ggotmCpLz8u2LSEarJAIUHtkoKB
aFJlvdn4UVFW9XeGuL/uW+BlVzO06MFijQ77grulsPjnYboeOs3PFaEwI7e1doZ+
prnmwaGYqG0nExAL81twOjZQnykGQiRNhcj2l7gwM08WoApmPj8xgSv0wg3pnebB
X9cr3j+4BKv9FH8fnFGrRtmtb8JldQdcNZcEeVJfhltkSzc3Tvn2JrZY0NfPeoYt
bw77YgCVOXpq3JuHZSf4AB4k4Gv0U2EGRIPMeeqks4s4uH06y2uIUM3Bm0q3biRm
Ore61ojE02lCYpihJaoAM/KLq+M0CIdLSKOfaYMwZ+TgbVn17EeLSIl4uLVHQcwX
WQD10laJ/rKbruWPLb1yVsHYL+/l7ONoPEXBh4ZT9r+sbUHx20Fy2z5XRIGlGBVB
Ajll39iUbNG1remeuO9PjWPW2SjhSnCEIQqZPL2kebrd2J5AKcK5uWjZad3u2pjW
dlN9YSDPhQas5eT5SF6tqUQcLqiYpRLCBXtFVhEQ7Wl7vgyPngzx6cGn2kqUW+wx
VDZPqgBQMhkdwrqoELNM6Zrwm9HEQTmMMZgI1DemjjrHlzKsF79prtjrSKqTtLZR
PtWVU9htDtNyxw4F7GWPg9IT8M8TyYmu/HwBz4TtYlAM6N3CLxFYkDKMHPqQH5cw
c1a+ewR5TGqU3krwJlSUHjTfSsfgL1yogoYE+FEXf+HcK/da5++XALuH/Z2Q++q1
IJB6ECSXKrF0Xqo8MCml0AfpVf/FQYJLj9N5bRMWrFUV0BHm+eO1QxGwg1iYHN2c
5eCzVgcVNIuNwNI//6vtkK4WR+LTRAYKZNyolw3Q+3NC/wwrIrMWUhh6YK+MVeUS
pZf+rxAVOvLXpqEVXvAAvonqPTW5BKlbB6O/8jAFTs4vXCe3GALbkVMzair4YRfQ
WsCA4C4huElTByo36S0vLX06zWJYpFxgEqlzZKYST40d6pytCgSGBzzHLE1CSeR1
UpGBrkblG5bIeuvyZrtV1MIF+Ol5Hv8UXZZ9fIPP6hjcStvOPbhTdNGfOOKCU0Pk
rd9uiUUY9+ZUJshKJ8VUp4z0nKt1Mp+YmbnCCB+MgpILhnJ9pJiJ8gY/XUONcdme
3U4bO2mIqwuHQhZKEbzCzZpgeHiWSvbI573h7hKFQYUEGCmiHivrovhbx/o169TC
j7PoPD1QnR2xUYU1Kp/nxVZnkWkwlJWabfB9zccBlqEdlLLCRM1sJrhTj9qp8oYf
M4XM3c4/nbyUZgPjmRSG2AcaGuJoRwBqBg+GTx19iq1fRy0QQVhX/yuPgi3cuE6k
xVin2i+Remn6aquO8qWWT2ejACRu/Af4vL2HB9Rniy393FznhAGCnMZ0HO6Y6/lU
768zGGBzW2gkIpQD/zRzC4H70ipGKjaKcBJkeXkslWe4JjJu+8zcESQlMFFRNxVY
AgpS4HitHvE9y+y3wXZ9uqHNYJqbOvnIKFpVsMSiZxmkEQPWFXZYuWpNQqM+3NGO
DXgHZRGOKNlBn9CoZZedeeZQTLZ+c8bHcWvkrp9iJUtHGKds+3Rer3BAKYLJO5kx
5MLPVNHoeMbcAXpNJuNo1JhRFwn92A5/INjMaf2ifumfUdngn0p/InNe2GT1JaCn
xqvyelq/4wYD32DEp6X06HbP2gWSKCXX81FRkpssfRexJrpyFwPW2ZP/t1pjTJbV
+lE+dNHJ/ln2B9cKb620UvPKc4SxkieKsMXhYmGu5zJf7zqvxlPgWQWZ3xWJUWdk
5lZgRYQ9QljcOO7AuYH1uBbOMDcmFmLH+3SzJinAFu94RCFYEaQZCefnOSaIHyS2
fIK/H14w1RTIeyZynoOiJLVcw1xN7qFfjPswkt0Ursxi3UTCNTfIeTfhrTU54u8G
4Oo1bjELP4MjQv1Q1JLw66nmO+0uAF9ARXBb6ybU5KpKfvtT3oNEdJcDiPm/GDS8
xwy6OU+SbL3aMFNzRcUil4hVorESYRi5cM8omXgehjnCaJL0ZuvKx+xMAcB/fHsZ
NbxJHgg7CwO3/CRvVIOYb/orWJ3aPO+Il/w/NAfYgIITG0pzm4Mx/VkGXc7lkPub
KEONP1kG42PUyKjqHqJn5QF9BC436yiLGpRkMbJ3DDoYvHSytKx1VuDoXXH6G2RD
oOJXgQCTMGdtKhFtvLa+LtXe6n0Cwlbmh7tjK06/4fqO3bXbu043ukCgFpeUQkQL
TT65pgDCvkG2FV9DdFk9hVzYbcMw0wfsUcyRGYjwc+WpJJ92nvSUgrMRGtKZDxyr
z3LuehjEnt77zS+BQ2eCamSPaJ42jBqtDV2ARM9/ScX556QSKftRVe0irlt6a/8t
5zlW7WS9oh/T3adIxV60eGj0bG7lj/W4a5suW8/xSuslIAPqqfRJwbDNYLF57oDP
eT/YPzaXXaF6Yi+2MvB+l1xEXYnDKdPUP75yCqKOpa1ytBhoPEy1fZoEDqciEl8p
jjS2Yfk3C4pRaYropZ1UTJ7YmmHTuWqgnJXhKa5fYDFOzIO155Vk0cpTEks63Q7C
yITGFBMIlfga+z7lDTbnL/MlbPuHGP/v51uXJ9fnLRX1s8924MxOuLbM8OpjIlvH
KJ7paC7vX1A/yjkUuUuuTSVR74v4/B525jLCXhV1GpYnHGzuNGaBk0LFOA7iRNP1
yh/cvb6P98i5bZ7ePwmQ8KI6pTRdUbgLHsYJbjz8Iw/u3fyY9oXVbIgibfL1yKyh
N6rrFDlH31Z3uSjNuJPJ9s/VaanBMDj0DsPFcPIOlgrzSHE4tan+Wy2QrKyWHV0O
rZclLFyfQltiUIafrrZpg0Tudu0D+A2QOBL+wi2TiT1iRozd3+2SV2LUe5dpf/Cu
xuyEDYM0TpXor5GaQVhY8j8vIUITAlwJtB11JCo9X0N7ZZGF9qcB4Pk2O3fduL4S
V0ByU2smgYuM9yyLn4Axud6ORIvP1dGV9VWa35u0YyiHHf8Pe4WOZFFwqJiGYQBH
rLX/oSu8yraZs79ycQFF995mOz5P8iLkBLlVWNLFxbLzlzmxsfsfVmWOEqOLoRTX
yQ0sFWw+R+F4DGd9uLjpttzI0hHedQU1V7jOdy3J6ZztnjFedR6GcfisUYdDBHCS
c9rPl90+nocfVJHhylttOZVpf6Q9Q0EVecwI3LLWVEjGX63wUWBWmUO7qmkuknXT
8GsFIZI3NCGk2D8cFDG9GkADQe72sua9BWe8Mb5V2/OUxwBIaFeYWgyRmGAZzz/8
fXz9xq3rBD8o0pGx8uBoWNGAMJl1LYo+rbgupZgJ+6aecrHqKlgXtygolv8MpvqF
jVvDhCPm3eT7It/Zhv1/rLtK4+95fSHnp8TQbF+xPq3Pm7XulwmkoBAjjI3W6iv4
B0zOcjYYlANyxcneUAevex0SevaqsgM1dK8oG522gZAuIKM3in8sW+x6Blry/vSA
6LQPW7ADfmOiLheoeaSA0w+RQzjLcDZvsTK1E819oCQ9JfrC1rEvcrxb5DmoXiMn
EQ1c3t/qUgjru3V6+mtFPE51umQSL0yFDLRbPWMaTpNiyEbeI6/UEWrlOpOsfXjV
FxG+QpBcRviiIN/X7be140FfzWbepn3JaYE0WDgNXPzshb8OLU0nMklwCjUTIrhB
lb69xjb7AYW4nA5QWa5B3PlwXQslRqcrH9C6G50wJTSQ4jfIyp7gKVdoa3099ZG/
+zAiHrNQfcLNBe3coyiGa7bbkDHkpoIn8uXiDvKLFIPOtUB1EoJw8KJCC/X/QC1Y
z5M/kMLKkUNZphWv5aGZixWQPwbUpSSJzHGYqpjsvKWTUewLmcY/K4rM6dP+0O/7
B/H9DLXUI6lccGaWtLdAtDui1fzeI2LaBXWEnkFLtHNsjGc27ttfa6KzV9jw05YM
cABsWnugwpyGD3T7Ubwj5vppfTHhOZ/nBZvs5hxdF/45QSIEzm+qFTkH0yZ2mWTK
B3TYooNNVzllLNhnDfDgElkyYXlDOvwwSXbpaXcpyKU9IMzcSoP4o2rrgVBJHTFO
UzfsW2BX6tpkr4fQMSD00K+YqwcBqLKDs2JTV0CWQWyEjOqCRXPO1I35yE/01bNk
+eRiGxeES11Yx/ioYBjW60mr7d5bTalChxnYLLDXZZyWL5XZuYvkWgA8Jq1BbDw9
mBFNnTeKJL99HPiMCHedYsMAYoccT/Yl3WuIBY+9SG/lbWK5SKc7O0CgGsjbp+hQ
8W+QcHqsqrA/4co/620sV37/yT2SdtKlcIe8QzohzaEmZyrZ4IiSUTkbvX+4yeKk
pOzWf1XpiSYdtvQFCEp503vYWDFTTMxf/hHFJ1dIM9xjPuI1ZeSZfkQwhOJi1us5
QnHbuBFzYa3rUZ4e434FmbpN7Uot6shcEygIJOcl8MoJtNbz2Y7z9sskDUKVHMuZ
Z2WtEm13ELTh/S016T9Xyokja2ffHYVMx6NVZe7J6lWQSmjzk4Wwa7AWoGbfqOv+
Sg7669OI03dT3HjQp0Nij6FTCTuL2xDmqQV9RoU8xanDzztmKYqVqKXD8jRujPRi
WFmtr4J9Q6N89iaxUuorpyjtrsuExjZ9AelvK5aK1b/G71AczRlIIeV8k/zeGkLO
bSXBI17yNGUmoaNi3mGo5p19oGfjgBWMdHANLD7snNFxb3WLXQtBbs2EQYmJ2ND1
3hv+XMXO8uN1/sZjmjebuHnr/tWS35vajL6mm0vUcuuIRyoaAAASWpzPKqc7Bwsa
WUnrLB99OBhNqCyPa3QucoUTZ5eD17jgh/Evw5r7odEFD5nUqzEZ07AhPnJuVfj6
7uj7nIChusuEdtCjj1Y+JBoQ5VsdeOS26H3O92Rf9gsEd0m6X6wS9vCWzqVyYWrM
gYQgamQLysSy1m+aQ10v4yZa7lZUjBWOdJCS9j5nFjL85uhqggo9dpkxSslW5IOx
yaQSZRq1MFK6NBuqEnpVAtYH85uvZN/QAI86SbyRgcs/LngoSt2H923zjFxqIgMT
T9j7PK6HU+Yb2FnjeWcvDBEYBC50c3IwPIU2wxZVQvU/gTWcIXe/hTXS6gFsNng2
imUfVq2CvLfg9mMiDjbQrGF86kP8aBpleq1uS+GtDMvLziD1i6JD9Gzo14YtXJG6
Zrr/wcSpQjEq0Eo/NjW3rxjyFI4wDFszHYQcQ0a3TblSxhxntEl2m2ZO+E55J3/b
Cb02K0+UlquwOdRNs8QqXhpxy2KCbBAQ6RS16vVIcaweUUc6br2P2aYyoZDFa/u+
QIHl+YJkzif+0i0pFjd+QV/ze0sLEqyJaa/RcbcNwAw/rffZFMUxYPwc55JSiN1G
mhlTl2oY/Eh8PYP9mY69TU5TBG+P0HChDtqIBBopzA/6hBDBXTy/cv40etfFMiL0
AA+AtBEqrJcrQEwzBwsBbsI8n0Ed3Ymef+5r1pnANCd3ETggBbu94Z/4FpWjb9C1
2f8fB/2fGF+rWIyBiaa48LfGEOgaomzAalDb6k+ZeH+7yewnNJr4Napp22pxd/rB
j0ZkFLG1Io6Sfn2DPqXMQWFFLUTlgN8G0CcJ5863NKlz0NLocO1fVqsAgdtLhSWi
ga2EjZEF9T+yp+Wus6eILif/yOILWOg2v/FwxGVc6i8S8GXdxIfAJTuAfbrILxfO
mUEehVhMKpNvb5nc6LCeeFU5CDy2Mq1R9ZfKho4WXh2/kaMtfuEhykweJJMB1ZLo
XVHtdN7uXs8z7l+/57rGZaDXUSLlYsD7pkt4R3k86hlPM7N03ZVjuCJA+EXcQ2ED
fx7iKtfBLveBYchdkDgaZlnkbHkC2dzonewr/DHcXwfXUXHfQlA3x78UOoiu8leY
qcHTHE6VhVoVwvKAIlR6N6fvffO/dAqjJN52JxK/9PTfUW0foyzbEIpe864/2Xqm
mt10QRUj9jKTCeoEfj5rGb9R58NYFcoDRBpU++7o/1LOilR0YjPhjiNQo/REtL1m
RyCrC+F/zF/fh8/el1msQQZ3yCupcXbGWbHA2q2iz4uAi5rbmUtsFMy2/Yb74HaC
sQSsVi6/JW+6azkuQ5NdpX5q1CFVab7Cu6EUMItZq3OIQzJzV/2egsDv4aeGSbvD
eeDMTtnz/5YfNJPV/2C0tfPjgcsBrDDUMoC4+g8RWHD5q85rbhF4xxPe6ykGIJYU
ZHTqu1zEadFOKcpNIVkqbUiea9bsPPFxHIq7JsH6vYhBpYizFX6zA24SasVVpCqA
yYRFAYfyeQfDY8wt/unpt6yzylpNkQnI9kWkpcWJ5QkcEBsc9/huIaPUcKw2FNVl
OvYw3i60XG+TJHPaNJ9agIDl3WmX3f/+G3yQkgpMNCS/PLCs7v7NxyT0Gg+o9UYS
Og/oD345m+f0dDrAbSwC8Me1expS6yt3ljQSpIzOs5gtTskn1eBmVt+TfYRNMMJo
O4eFqWOQYctVn+SBDnQ7/H24lrbaVnbZ701ko+NSOR2f5Qv2yV3gFxCShLk3guIr
Ika7uwAEqWqd+7e/fX3f+bvCsT2H1l1pSTyONX5QVpdqse5vqiKQyoEkpQUdX32O
22Y+uv7Q5BGrqSJsuSb00SYDTjbblkx+9HDxg2UKlQxRHZ7ifxFtel1tgpEk4+iz
Pi/PM3COdC22SJaPKpIpcMhoL4rVASuSX2KF/2VUYxzuGXtyjDza8sfkWwwz7U6N
JDgeYF9vibbUGTOgS6QBW6ErQCb4LuoL/jpEXDyzobnt02nRZWd6eMQFMgk0Gst+
Y5ysFL9tXHT1k7wAQg8eyAR34B+eNFb9H5h0bDCm0TxOGVekO+EsvQG2HSgSfFvh
wO4LG+xaLjCarVNXlLMbyK4I01nf7VM6eFCHZGXEmgugAzGD7VramhSFmNBgS7nF
DfAga4y92FcZPMBjSsrIU1DuG6/f8F+WnN8jQYa6E3lNk+1pYqqOlrrLHplyyCCW
ATMw3j+xsZCbVopgRaPYj6koL7ISYOBdMpbMFfcjKgHCu03hxRvTxWEn7zRBxUyX
psAR7js9LoKTlABuV/88wwKr2Ckg5ABmRgV/9weAByPxswgmPrkNP5wfLTBzMWeB
wWctgxNrsS/vPpKHGwBl1eNGLCLdNK4cscdlHLHXtHj1HoYNaDM7mgZhBFYkSdkg
VM/8Y4ml3zxzwHxIJcEur34fcpSnt6RfUgRRxTw0UDvQZioGaoKdWC8gcQ6gAkRn
jkAubBel6uQNOWP4lGNemRzTQOh5Gj1NJnmoOqOTHome5RoDzZqWSxHXcJq083Jo
josHLrNrd2L31HqNnhXC0QYGSFAxegKK+CMXy213HyHKZ+rIgzltIKmcsTfHIvWv
dlWWxW4V8WSd26czrDzy/VAggiIuhDaHrrY6Ot2mhetG5H+p+FLMcJbOC4SJUzAP
BjymAmvyFHG3KXTg+Zz6wceZ3hFSd/WZdFksqw5mteHwpAFe2cuKlX2E2ODUmcji
VH2t/hTBpZ9v+iSsbJD48m/0lUPqOguL3aqv3O5w4yyyqbtIbFKjIUL9x0ybKhV3
9dS/62t6xyvYcuVJpNDobCCdqx/tWxRi9ISthSimACAex7YPNn0Etoq5DaDZz/xF
ZluakCAAxraqmevPvp5wD4UrdjK33swHa2uoJlmIj2KWt3Z4KGF0MvUCOLxDWZRh
uE+8979jun233RmFTTMsYEkbfTxjfuXeGQS88LP4JHQpm9xF2sBzJg9MN8SxMTg1
NHdXpHqz3KvZQ8Hj5r7RnfozmzblWVbcCHYBUgtlkpUqcF1UzjhJvbADhOXqydTJ
n7Utzlh9PeV62C88Ntr77Y1TGUZZLF4dRgLxM07h6mi97mTotrEYxBixts4RrvIk
gQQ8+NSbKYSv3SiRT4HD7wlZxbAHAyBspA1MAZMSExG3wtQkjLIUOq3QwGomkU/5
LHVGJAxf7JC8zin7sOcTuPPARjyxDmNrDzLYgpsxzQOA7n0GznRDwHwCm5VeyPnG
Jl07Ff3IFlL9DqIGjtqN0WLNFKnXivIDJPb/aYFKwtorRvIaOVHOQ1EUpccJy+gV
Buyx8e6XD1RwQ0DRIAOEUeTY7EH5JjrQJG5yESTPcQFk3kc/Yp7mplZVAgqanD4i
jMnttMrpc0JYLIu+p7bqUmYpxuLoQvu/6EKQY6St6SFsS2NmQ3fJwXD80wk70EJ3
h44QwGcwhbvrUvyDU22cs/jJhziJwixu3YSDvlHNvTvm9h22zbIBQF6e5P+yMfiA
PlABfBEpB/GgsubvGbOyVgG8NDht1ix93WBt7ZyrrIoWenSSlag41hc4teAN8CR2
T3gw4/dkMFuOLgTimztrogUBmSI30wSL1jrfsOb+z5G7tmFOpXXTCORvv+eH5SI0
YFr4wYy5jLT7b9ojPhkl4bxyw24MhNHRcjttqz1wUhbKiZKJnOKoLjJLDYtToEEL
aelvn7HQprpSP52V54D3xsdn0yAGT6dvIBKXxIab/KsGjT5xc/+8qsnVVxfh2bK6
pUyEDH4YakSAWeg+nDmxCNCj4ut3vjlFcXsqyDBDbE1u0+okTb7HP//IIWjFGht5
ESp3Z4K50mVlgH9b0DqfWra8lxdCJl122o8kZXDHuMghU4JpJiD5z3QEs9zqlE2w
YRArBIfjjMFwIbKAM+hn4uzOSm8LmmH8XOdNf56WB2wzvhd6gGz8y9nwgBzegM2E
kTgGfr854ko80LmyTsW5IS2ldIhHnEN/4DIx7d/OaqqqD6u7z3caPO1ppgoQmUzU
6plfc0RDbyXIXfxVFIjMJft+LVZdByXaNJv3fF1b7D2zBpinYtyZasyNZBI/7HqZ
hH3gDdcdgv4UstvuftSOsNMwFKqO7w9n52cF+ZCbnj5AeqxQXTDgYa4VNmguqnDl
4nTy5fyCMTZ+ynI2Wquo24AxBYAVirzWQOXSWiXTqH9OFeae99NWSygzk7SP0gAi
+h4SvnYpT5rNhDJgc1SRaCTTuuoKTxVzcZ/+upGu4Pw2XwOGSNKRy8itFvOeyWQf
Pov/ZSeDX3f+Z0VHEHUq0VDRmyyMVVbdzUl7yvwlAHfVugEBexAW1uMQNLRgfYu2
gvWuJk+u/WzF0gqFzNvA85OfLMj+ydFFUEinnrw0Z+Wq3bX/ECQMDR+qIAucIAnJ
AYOvz+1SWGkfdEeDgCezpO/oMxHDY3ww8/RXOOk0TBpYigCPA/sHnpicW9ee3kYd
bBOlP/J2TCOTatyGExVIjSeDZ+z7OgHYpHbLGI3jsJjYMGCXMHQIj1h3U6SZ0SAi
JoAwvUld9isn+UZOLoPAygy5HwbXHXHyY7AYO7q38UPc6CGcSkwNGACNsIPCyDk4
+1rOQxpvV7lQEmCKUHaqa0lwHr1tdkyblG0J2mHzBxxTb5hO2Ld/z7rPYXXV+s8z
yPOYM07Z2fXCuDdJZsOOvSPkAHNxruHqROuDD7r3zUCZfFTuhpziSUmBwBAAPRaj
v4HqoRR3Tcr/upbtG2BV4oj5xVo/ahxNGis1MwGN69gyc1MmJr7FzQQp7icbACdx
VnSxJKomF/vco0YV6FTEU2CXMep/gxfGzJNaFt/N+agGnhVyk8hporh+qSGRoBzF
ZjJ0+qf5/sm+jnDQR+R0jmQ256kDXiEgW1apYHbgXrtOsE907E4lzcZgAabvCJoA
pGl+JiYKAE+C1rM+2icZo3zKBY+M9vpwVPXqLuqV5dDpkZm/IWI6YEIlW8cRjyqk
MYH6XE+mM+tBArLA3if24f6Su8Eq0tiovHmnQSccUUmg1q2irghj5DwXgG9Y9RC4
umOa16OXYQrPIvpfFBjl2YOIrmNWUsDaPVMQ+rNjAi54Tg09PvVsbnu3//ZSribS
PQEYpoxrYrrkEjAqNZiNs7s5Ff2eKLZpecuGi3pNbDlYr/UJ607YSZ4Z5tM6NZ9j
diT86ffSoPla8sGf4BlSbwpwTG/WwGUHsQL9bWSZyf20jgsTemaPhuUB4w4c2EIK
DsTvuAa3FGZhBqxVjOqsYK3tn0VtXAoACGki5CG00D/5NVaBjvDiZL9D8WWZG8/f
lkj7B2fBM1rFHKWcUJNVC3NP9wVJvxMjmOuJ0G01aNQ/N6d3dvR746d6LsRSGYvx
QC6P8zsGHB+9hsp4gEIeGaN2tD9+p2a6ck72wqBRygME6LZX0T3Tf7tF2J123rM3
jxCrdO5jbpPvkkZDFwSL9xJh7fTyj7ZYvIWCPGCSWW3lq4ZEOLxV040TExKs6ovU
vo8oKD5lsbsf4ML1/zPufbyK2ooPQZeiqJpRwGg+ioINlcUYK4hIVAC5cr2j6zP0
HXvfTQcvJaDHBiStzDf7NtX3EOG3ydmEexr3U+cIqFrWdMpr9kt3nqJ532Da9nmV
KaqhFnUpbr/1miJVvPIgBQB3laQibfBHvYSktRLZdjhIbAQ3ZlG8vUiwbm6Ybskw
wPjf0QzXQUpFqDNDuWu1EYOPkrOAObLX0eXcLnVB5IIJFXWJ0XEm+HkyBgwWJ+7K
MS8qnV1rk6A5D53z0u9SNEGoGjhSgeTFsig/hCsItIDsox2hpGWv0j9CYa1iZo0v
OVmhYNV94xUCFE4O5Fw7318jMeP64sutctkcJKnyYJNy5bMDn4eI+kH48swypMN0
MhV7X+kX273CKZSeMxcqobJSSm1XtVXzYJlkVE/mIPxYXzGFSa3tED5pvZPaM7i7
NRmUY/xo1CeFzlVyEq1TA7jhy54rrp+8aBVVajWCdnWT1W/nfWokob+hXjqDtVK+
ShVSUZqPaKPaaowDD8/OtckxlpIR8ya07bg0l312WWqEgkPwTan/QtBsX9Br1Uzj
D91vAPTHIojxdPxMdjQ2MbkQXe1vzyAZQcEoVtyVUN1plcxMKn9EfuEERrM2VtYh
u3y424oh7Tc7aFhg1iJHhQkwGoxHZJgFxO/4Kudnsp8BUvdowuBx9BDDXgjnBOw4
pQmqi1CCBgiLXKaT5KSrWkkfP80KmgDSmD6YZkfZjpdz1r10HN7Jh0PLUHlWguqc
SCodOzFTZiwWwgbVMnnI1s3lMhZpspGK9WQS8I3uVnidEyeFcH3p5sEd9FFK0xj0
PELyQyr1Z3JwWvrlqe6Wp9SaM6bPNrATherqX/Yyx9XXRY5DcirUYVUd/pSutzy8
QLx0sqobgakB1sn4+X9mUCY7t4p7J52aynuHcMA7CVUqymdB3valS0y9wuBlqEfa
AC/zB52xVdugy/xFd4ApqyTfUOxokfWXGbyUdcPb42Qmn3vKzOz4AEbv82HhqOtN
cXpCPf8lKGF/B9GEZziYOtO+KMG6ZEfUIBw6ub5YR0ezN5wcnbXsr+KYheNPcBAT
fqomfKSo+nZam/TA1AnYhKeaJQTi2IRRQ3ZsRlLoROskvgsglBW81s2BjRq0+pJ6
zADL/6BcOmU5oB21+DshiwOAZVRJMiFxGfJqmfPMwwXzBPtK+r6NCu24bXVErL2p
orz3KFAfOzzG5/42l7JG65Jw44GU1ccNFNHD1/wwzeWpF7m4JtLHdASNRxAZxjZ8
Z55zPuM4buKt5ZwZU6QGWThWdOXBvlhuPXtXL6HbBLm3lHb3f7Ok/kgrN7dE6pm9
q5N5vklgwSAUBZiIrF36pqCElZt5QdxmeHw8HvhNXPHoYg4AOeyE6R6uc9A2vWd2
/wpk747B5nI2cAIdTuFhquS9DBOpwW/bP/g9YaYZfKMl6QVzIO+xfpFvweK9dlAp
yFijkFK+czMCSMe5qKE6elSa7T9fktZo2n3PCe589qqiiZ8Z4pyLsmarrln6qKx2
XCPWzl1seSy6wcRCOUJyQb8ywUpKPqLnw//GOhKEUpX1Y+NIm8r+dkMClSR+BqU3
Y07DShRwhSIEJ6MhhfT07qlKAUqVNg+Cw1dHrZ0M4l/v0T5K5xpxd8fDmg9t1YBl
HmOduXczPFnZI1w8kT7d+B+q2INS7DdFAUuCU6cWbyvktMJq4Gd1gFk4CasTVV5k
K5iLpDqaq7OmgSDF6hPYCEE/pzJezmUDFg/Mu1wzUXAxVnCVy7tor/eLd2rFlmsK
1t/gprCHXLjDwU3CbzD3ADn4YJQk7H3/VELQiGtOwIBvNPise/h3wq5LPBUHJB7r
eymzWgFmzbeP1SgxjbyKsEk1CyiNsJRgYjxYFCwEFzv8cN/YfQiX8KDZ1P/dBxTS
Zz8wcQD+JM/kV7NctbzR14qqzbvbMzvNM9Uit54byn1W7EsR8pTiJq+CDyQSuCQX
6JTHuiDNEnTFBQJum5rps3LIMAXzzofdZHN07NhXYCARYg8ZafQJ1STtyc/RM0ij
fdAZbW4IccISOuBSfMXIY1q4p/NCaBuXdS3uvgcBuaDQPL+MRedFBRQCMe9rfL2R
asJoXvoa087ZyCFHun4F83Y8Mu9peQgInK8qjTXNdkr/0NmqoYwOG3uA+NrrTpVQ
he6LVJC+R3NgMQSBMFqwLslRL13AXHaNHqQY/gk7pJ/370Jb4sLv2SQOPKdk6h5Y
dBtyO08NeMqNbjA9CGi0laxBg4ukTw8QsGNH4Yv4vyIoUUrI6xdDEZTJHe+TE8SF
zgVHqKv2MOLLc98RFxu6FlxKOxXkrjPiOZIZGmG+OYHtAO+fLWxngHBVPHQmLLlE
r/7lEuedYO2QM/UiVEIxaWhNpQMZ41wQVO/g89Bkb0BiWybsf1/eRy/uba/+NgxM
dTeWS2bPUstBWuwkpJdhWT91ewmWnFTvCJio/Xfkn9BrpnM/DfCSF2FztTANl5s6
QBhyWbHrMYSodyo6giqJX4EBtU5Gbvi9Wlb/+Evo39kVe4tgSO023mKSOWSJWX6b
i0SJVq/lftrLXltkv1OGoYftLQqqku+yoUYH5yJVlgnBzln9DnB3In+3rT9KaLjn
Jff6Aj/8lHZB+7lvK4EPYhqcgNV/iNhTgVrVADASc3X6R24vkpPMeZ5exK7I6qBo
fNYnpt6uIIkP28kv1fNcedmH3xtMzsfFK3+sxahrXZ1bds2pPcVTw11BGMvxA9uU
gl2dRuIQo3s8R0hHGqYjipUyYyljL/BOg4MeEkoLNzW642NE5zxTv/Kl6WyQcQcL
QlvXB9bKPoGvx8F88T+c64eVoaVphJbR6PeCoV/1sYKCdJL1JlWUnD2AOm46LDEz
sOo+5/+h1xxlexc/+dAvHUB1191c3N6tr/nnJQT4ct0kxPD70aQBROHujqc3AmtJ
DYFtEjqvr1awksH1H0dwtxf1gNxTdjxypXpvDR8riSgCNYHYNfbnLiQCm/8/3/lO
t7+YEW43OsWboWtk2uksSQpK89GULEzG98wQ4v9Vpaja/8TwZZzOOO+sF/u8EUDg
RGCH9xa6RtxNOkoKgtrKZZXTDQW+SAFshswSPnzexqYe8EZ0GrG/DWcha2cCzXnB
xBgBGfi5plcZe2PtqNTWsxeEP3ON/NHo8Ng+xm4kVDTb1jTjWXQDDHbWh7xh0Fwp
KmFHPgXGvBpTGdy3KlxqivENh7gPwVWZjsEn9qPicU4GhX8hdkH6yhxVPjyCWi4Q
zxuJ0HkAJG2LcUchzDKtlotvawwt3jwYeUty5dSiTj/XUjDXBHTp2RJ2XknwNFIC
h2eR/1eM8PrVrK7soxmY18jT8ikNlWh1hXjnpgbAAwjJKLItpM3JxAnmBnxWQOQN
WQ6xQk3jms8DmRMPbszSAi6IPs40F+7tSaNgLaPulKjCH87FTgIojPJMJ5upDtsN
MKMFNrLX7R9f330MZ82OX7slNoFBKk4HHmjjDF1sRonrUOCagHtYZqWBfjOClgEU
wWR4jN6PlED0YLGiXbUmi7zJ2F3EOi1eMs7ufgBVTbV+S4IrA3no9kce9GcCUgw2
zhCv2G9FWkdDx6Np8CoQoVI3aGnXGxhs1SzgyCZDCfdypImPHfuEnL3HPFpHh0lc
kg/P6LNiSBFo0kLLftbXuanQuvy5V7YHG/7eE/JggCZG9b+iqmiqL1zGapyqiMtW
603ekSPKd1nxhFtT5MhpzkG5qXPMgQlwYitDA338jD2PInIkkvzHdD3V4JrwKA4R
50Cl83d4xpxMNmdq5rfp3f3YxDi0ShBg6PmbyJyHVjjmAH4HXy0cDZzmy/fhQ49t
c+6cpjsXWp4/Trhi7yKG+EJYwxzGYS1EdjKY6YwDiPP3xA+BVBEyZX9SmhoZKy1Y
7QwuDocYkjiRho+J92tPbAUhxMGAoCDoOpNY4Mhy3MbVwggXMMPd4qsg3gzvqcHz
yBcml6LpU5Fv/k4fhxrpQDtju9M09i1Hy5mDxAz8Wrf5FpD2VfoinxhlErsn1JYJ
a5UZY5U7yG/FppAwdXGtsAukFvo1IC2L2YfRjLGnaQd4ige9Wzyrt+4L+FIihCu2
stuPjFe9CJWGaGLLeyrO0TskB6Nno6OUCd0hGDAtw9cextcVBlEIb5HTzV9toH7U
vkyQWRHi8vGf2bhtXSUfXT2HrYq1nacZauahRNeUlRN1KEMR/uzJMPtdCh5c7iu1
0efIT5TryK6K0UobucIx8WQGwu4BLe+T435ZxyH8irD90d0nZM8uGWHkxlqMgjkg
hytn67uM7uTecfdhSD3gsjN3G8ARMKsjYOh9TCZvl4F32VSoXIe604rMLIKVtE9E
CVBOuqOEqX6xRJvOQ1b6tWr8L1JiQ5vm1N34n3VqD4j8ulwavDgW8wjex/DGg8JU
iElV7TK9gUdG5RS1PYrnLT0B/afRdZbr8pFnOJpLbMiN0cmkNo7Y/r0AcU0MuibO
jABL9jHiQTxiYA3pa4L10asLSW6cN05q2kkIOFh3ZGyqNIxevQEtyy5igF0OGCY5
e1mqxOUuuSKPVNvmhGxCgJr5tOntEUK+EE6SWrQjFV1qlgHjcAvhzN2XRoZIa9l8
DA0smDCxc4Bhad59hUQAR6Gyw3EusrSGcAhwTMhdcX0E6KARQ8MDHPluiwv46IHF
s9E1vqncj2X4+7cJHwnEjAfL2RDKxE2UxTq3fJuZ9Tm6BZJ0fOA5GOBMwSN190I8
90p9qeX+StnZmwT5g+cP0J+io4CM9Sh6OVhtPYcYsCw+sXSxXnr4Gk+7OLrYybHR
JWSZfEj2fBZdEA9uFfhBGVtXegjATV7anLDiw+bf+0+CCE4dZiiWxtHqTqsFykTc
bDHVFYDMeyoaQVlXjY243P/EQKIGLQXIrSGwWrH0MsdSSmXun0zIk8iCnQaoINcJ
BYnsn3/2WdDM1PaFRAQ1GJDqY8pGJTGgPcBKuowtfEndltBZ+aMu7kfiwufbij7/
Bo6s7CIZ+1lc63C8Im91YiWBGcxzi0YCqRVD/+j0RlM5CL0014cPwEWnBO0viecP
O+T+NvCb/pS6YiEefpqr0ExrOqRdI3s0M2VQbQQdZUoWYOWbxTjMWv0TCYZiUxDT
rPWBM6NXqsPd9/v5e3MRMKDII2VWbKFSMpGgruVeevpm6QE5Hs6EwVEREN2aTs6c
3iIjtKq3pt58XGuaWPLacM0aPFaf9Mcf50xmCcdaYriD3XVd8R3eQgZQw3lVTOIu
uh38fkuSdmhfySO8x9+HJIXPBlRWyH05iWajMDomJaasB7ZZdsECIhSGFDrzfOUX
Garq2GuitxwGZOVj3jwTTo0LJMG0i3WnOS6nj9AFFyFaBYmDm8Vy9yHrNPH8CC3+
jYJjMO003+SGy+82FCrbEiitOOGya+hDoZm3VcbzYMIEcJA4Rogu3M//aiHxpxql
k9WG6yuwG9FS+8S5R/W6DRlK3Qst6hzQpFAbq81PRsdejX5ovz04wCNL/nRHqQ6T
hM/TuvGGBIlnF0S0Ii24lyUslyaexC74lQ7tcpESo8Q7ehB+CM2k6SKtXReUucqS
H2keNtZ4JbaVGOK+gt6Kw11fv66XVqaPwsnsx3wZkglt8mjGo9HKzdSUrLGyWhN9
61P94QMmR4RJ5rQ2Qtb3DoJRaCq684XAUoEJOZNJGCrA1+a2dc4KEFGKhl68lkVJ
p2yul4anVempBJDNjpZvrw7rqfPrhGPpnW8SgpzzbdH6ediUmvyrPw6rgfnfLSQU
M+L4WnxlHPTWwAaLLMSr8JpGBNV7FnJEj+YEB7pY/lgi6R2pw1t5lUTe+pa/vM4L
XYJcJsOTAfPRFh4wTN1Htm92NsQWgNoRBj02RVa5V/2dlmP6YsHHhj8sn0ZtYC0x
Z9fLr8hKwSPm7XSgBSZJEojnGNUzT9t7fUZRVxav1VaAs6IvQ6NOAsPSd1NHUJmQ
ttZuhApYv0mbOkXq3S+2G+qE1csJR47uPS/gBjOCXF2JZI9cA1GXixcHsx7grAtp
cPL6klg4/m15yR7zSJlk6e0GRo07gKomZOHnkptT+T8T/oTN80YEtNYavvAxVlrU
TVefchDIAYYjO/9jrM26KHZTZ7Gksmo5NSf1HOI3scLgE+52vLUWbElu1luItgAe
6a8Iip21+9q14F6mzBA2tP6mi3wpPMO+Vdxvzsipim1CJ6rOpouS35r22OxHqm2V
crJ1/I/lMrD0weIZyyMntN4GXTl/Ulv+Y0jyFuDqrD4a0DDAl0cKZg1BA0Klc5KR
lTxbKx0we6WuHK4xX6h8hhabWiKshoIk5Y99ApS25X2LeGb5ic3AhzedtWPSgVMB
AJtu/cmnYYVIX55dPH92il/torUUk2NhUmwY4XC/m/Zaa+jfMl6an1UL4YLnuYUT
MyCAJqxG8cedq8SDpEG4z3Ri5lbvt0R/3H7jOTFnFfOwuH6wRFhn+bqT6Kooxi9u
2+GIID49PVeYONjGfmyruXZ8j2LtSqWszLsJx1V5uDN/kjm2//8KzYb/gyqDk3Gp
81jYo6qAyjmqx4Pd05zyu8rUX9AUDwF3E16l1JLI0VMioDw/46zxWKV1Ob4RUdrG
UDSt8lvJywe52vobrH+jXuqCdmqmsWIaSk9vvYBuvwJWKrXtzEf6EGP5UA3U68dB
o0MDHls3h7N4HLWYqg90cAXN9/rHCf78VMP3dkTBod0zzy3N0kRxKoaJBlBbJxEG
VupKdcnFo9FpcFEI7lbPcInRHFg45+2BvwtYkonZierATA1O/63tiCoZNDTSCzXZ
YQLKmtIGzruzj8CLKQBugmkrk9eBKbe2Ps7v77EHQlyEerBGlLv0w+D+pmqgIQBB
s8yoNj1gqJGwChVPSFME8ya5W8YIF+K1VdyXo/cAVD4CQHE+z5BzfmnoO2kp5O7t
WH6aMhLMvYDGq1lTw7SudVO0W3cq+pYFAALuQ8qiAKTcEq56mIAArub2EPFoRTcR
ExFiKIsUT0lUm4maPr4lB6cuUu9yzabcGxd+xYrvGfQxFnvJys9vG7BYAZCjZTgb
suPfOU8rXnUxVHjUadCDFsqhg9GEJG7nOI+Y6Ww3yjYhaaEEDdZx2b8SJoUD8kZe
ytubvTsOcsdyovqUu80UHpm2XBMJIM3nltRmTTkNfwTCFjwQlOhse6nfum+bWBz1
xLnWrZ7HupeO1M6pfQgJ4Q9ZWRvApPJ5Nv0Et4N91AiErfmwQJ+Hq/VARKMb7eNm
n1dnyfgxtpPtp3PPMiYwn/x8mRsAqejbl1OqdEWDLRW/+UP48LJOSIQpaUulDY4V
gqfQGN1JJt2Twb/JjQGwhbWXAtQ2S9fhiC5N+CS9x+nuaOL0Eel0jKzPtxW4ph8A
i4C/LHKM/FgC0KjQHnD1A4XBSmkrXBkQvOA+cMGSYgFtAdBH82zfh4l9V0hbsrzd
q6B7Sl0DxXNEwKqqPeWrIE2/IjeO5ORKNFoLFrfFR/BpipGQVLWC9HvSDQmO8y2Y
DW2wr3P3r/Dk8Nvd5i6UukjsxovRDLAdvkMtvwRLkvcq/MaEWKP++WSbfAksQC2U
F/Uk5yt2iH2CbuiHZCixhNJ5ag18xss9+q7MAKQx/Yww8XXYISRDx+SHLltP05CO
ffoIHGNUkYNNVi5gkuYRFI768NBaXy5WtVcWh8Ic9T54SKFB/mXCMWXXyFdoN163
FPcA2Kqy8XnOZ2/voXQfmyTQGUzCObgPdCF4u5fCHWPamSBNrvfYkIegBRsQB5qA
2d0Je3dMeHzcO5HGLLVZT6c3Gv1nSxTUocsD38CdfGGgk9E0kLwZLk4XJs43qnzP
PeV8tcLWdKmyHKs6puJji19f+dkiLqNHZd0ciMpe2B376gbEn5Y/SzrLH96rxyBw
/l2hLsktfK7WG/l5Hb64+Q3yXibrV3Gl4v36YinY/oZgBCfQ7VNA7Anuu+yehlsQ
cbDZFW/5eVIIyXvE63wVy2XisWem8PPfBg7xmiaCgjlyWLZ/qImEpNTN7pgE6LCv
jELNiVMkqj+FSqfQEsZ+LuUBEb0W6WtQeD7xQhNdtxEMxBc7FFK+C2AoF2H8Ln+N
YF/CVS971E8LiTNNuG5ePzAQYb9EJgw5gQkXQDeRUAGriRr8o3ye2MHmu//9e6G3
BsrK2rXpVW3UPTFgNosZ6k80k5ykQLk5yG0UvVNNjdQDJT/k7oIYyl5lfvZt/V35
Ortj9Hks5XmdIFN8l4gsLBzIAekwxMGBQdpc89k5qUUoHnOSRAFX2LN8tETswPH9
OlPnz8i1Me64zK5HtGqZeMBaY6seskp/mxWAAc6IkxTWJZ3mY2cBGFENdPbkoMad
gNWnMoEdYAwUwWPr++oiTAnVwBFXQmkF8z5KohGGvNYfgufT3MRyIhfngrg9XyVw
zkCIVbJHA/Ed5GD8ORThN0UfDvIUsvmGUNEJtYqL60nUi9HchTGJc2yU7hEpjxci
gU/9z5nMMH28DLbLM6vztdZOUng6uWcLPje6o77He3szKFUcxXDz/PHqE1R0Ehww
w9DqzonB3kzvg6u7qhjTcxPriDoaSzFue0ANxQXcTariAlqhIZiBxYooqd36MPXe
l4DWinnSaX24I+MGJ2njXaBcYjMkV1ad3FUioyruXOHltmi3rRpOwbPtgnYrS1j6
6JvY6i6wz+OAaqwoglYa+RMPehwzRrB1hb54lRp9rFO0yWlrwu0ydvhN5FnG4cMe
ckRcW+Py68/oBmRYCDggz38UXVHlsL6P0FPx4klJt7ldvlhIjEQvBY/0Ij+2hAMU
1DXb7fV1iV0aG3njAr6lZ6QQ5nHgnU5TG7g7buT07RM8qFsXUelc/0JvpkmU5U/H
ZVHEqCqf/V69quibhy+XLLlGa7ntg3RyspNmHyzbUqInQksXTJbDZ7l6Ff5eFGlQ
BA6fdagyXwye7k+kUGwfRxsqQC2yOM9y0FUwLXkhe7GQ5nk9ZTBlPu6Vxpn0l/8F
z4hxUAT3nbEWsR0fwuXulqvWN6qvJwqaJ8SXkVYpGQWinaVpCJIBIlrROAJZSKRy
eXSq030UcnJ1lwpXyRwF6WnydvnsMM4cSypTJeR8LdvVMu9uAVMuiZhTvPJDwN4Q
ccC5Wlvsie/j3/exxIIBXHrtD/ofmmWdlPz4dcSF3BlfLqDwzwV13Z09HMntkRXC
iVSOiTmK4waAzHq/NNf4GIqALWyQmEGuC2sTa1TNMXFFhlpcXvlsS9Yoz71XBpb/
R/8ourE9O/l/yBIZ9LK43O6uXStBy8CvLZzIECtw7Mc6LOtER1fJYzsVgn6aEhXi
dGHChr9XExF9O5wkT+KH3maiursr1nPjVu+jmR2Cgdhi65lBC8LlKv2oX5rMe8Cq
D7a1wdQHbriqF2EZQlsVGvzeS0dR5gZQEi+wYBJYK2J/pevRp3qYwGwwB8CiC5bw
3yqwVBgaxnLAGsCLd38tVlIRoNyRU8y1VUVRoJab7Kc54ECRJ5wYRfxlSOAkQALc
PdvtbV6pgriGcgvsT8V3IabuaYDKw1DHsX4BxPTv8mPGViOr0SSyg48P7pJGhO7x
vdNxkfBEzoYZN52XqMrGTDWD4Vfr3FrqoPc0tTxBqgz1J1ngzThyYOiFSe4kI79M
7zfj6zGLwPmmhBEqba/XUS1TIRhtc79JNqBnX70TXbuvYmeeKnncoAVzpR/goOtq
aFFQSuBbTQf6JXvprgkFzVCgi7Cvw4eXAjgk07nXyLQzD9jcrb3KOgK4i2G2sNbM
ga42tCGRFe0S+lazBpmvyLV3CdUJmaTEq0dLKz6i+3fDmA6ji5gHNd7fk2pu4nQd
xJjFguzSXb6ol0b1g2wQXe87foDGXnq4iM4BrbQOQG5g7RCSf4muydXfuLA0tcjL
pD+e/MuCgT1A8WyDI7kPOwTsEAwHgulzzrSO31g0OsiidnLHz2GYGZ6+eivVyGAj
UMt3ATeaz46qx02mkOnri/u6chSzPtY/zunagQg5x8ie1FZ0+sDNEUBQfnb5++Ol
iPXV46u6+gN71+1F8CdH+KfRClCzs6Hc1yvS1dqcLIpON1M6KwJVU2TDeA/nYT0J
ajvnofYtGMzKZDLWHcu8dc2vsZuYL43jpTTG2jCAXO18dDY14geo/Gn4WrYJNMi1
MVwv7dcdxD7LZM5guHvXuA7cL886cqFt1Nsl99cqhEOSraib7N7xrsPqNc9mlbU+
t07sDm6pgaTumggbE/khtkve2S1sd2tFHYdGR4Sid+CkorHpSKfBsjYo0+pf/NRN
cLhvdKZtFLX6Zz1llHHwVR9QyCA/H2h5Cjyuv75iHGVp3Crr43a3qTcDi8lieqWR
Dr5RQqiyD8uaOMCC3FB8oU9HJi+h7CJ7BZrpEg0VsOBIYJyKozNsEONiOs6bEpoP
5/kmtfbJo3GyhTY7CDEPa9OY7O89pb3JT8iQV1eoXbaX4lsVQaJCaxtq4XaHlfXz
Tb7uQGL8b+TuW5cKkcbuJuTLN3xS0kuJIggwizQAgDjRghlw0g2dCYvHt6BfImg/
fqBpUdA86Cpbs5ZvoM+xr2DpW4iWRnYbMO0O9AT0d1untmGdgPOOZNv1aNRrU4Hc
7zDYYyDa8TB31GMFegb2XCgW3Ihu9qkCbWodOBRP5xcBPUwPIqIectOTOXlPcno2
ecYZ7ha2SmZ14NFgC7dZyJVfKo6pBTqcoKX1Bz9LiaOOsPVg/Pyk8zKJIJJZQIQQ
T5tbKFHJsZJdf0wfbY+m5Hp7QzHnVRZK/6lRVgQirY6UdidSUXu+mfi0yhkXmF09
Qnk7pFR8UgBblk5H0TyfZ1LMEVy2vcD0ujsAEuM5T/Yg5YyBELECjEw7tBOXNrkA
KM3BQSR9ArrBICe6AWKHMz0icLr8iKssvzReFbGdnCwxWVEvNGnGu4xWHL3xH82c
IbzBhOos8IPGJ+vEPD6RsbkwlQfPSPAwyNfpkgo9QBYTNFXw2M/3xkeJ4myezWlA
784glNOJc7mUSPFKu6uJKgbsdVGO9Zk+lY3P9IQkgQRZY1MQYyrO3GdumNkFJadL
oD8F+YfjnJAFjGJ+yAopKgr7AvPS/20PBNK+8hTckeG7/6r2HknJpuYFMPCuw9G6
0tnb74sXWPuymZRno7VgurDUu8/9tFwJ2zu/1AzT1DhX3Cgb0mSJH8fW1keGbx8v
ODw9E8RXFI/F1UnWEy4zDtd62jAO5LRmEtT9HZ3jyi5hH9+O5TutC8m9NPsR/z18
sxzfSCMXOric3yUq+wO+/8sgcPG0jd1Kr+VxRdhfpyInzr64HEnnkXhYP/G2/M8M
Jbg/SPmWhHEKLms0hkaF+7wNPiqe73xHyrCj/mYebuiek5ztyNX5q3NHFaa27FJu
6xk3Dq57w7mAtq1YM/f38OksmokNgyIZ74lDoKfNR1owJLbf8GHhNb7EhiEcWWB4
bE15NtmuNxGwUG61ZVi/61Ql35RnctYTsz+kQHXqFVrIcj+SGwpTFjjbNCZBpAmV
7BaRKGnaAkJi7Eu1hfZRMgyXRz+xWtJeXlPx70pwUlP9dKCns/w9mIFFYnKOXOaN
9du+5sdBmSeeDEPAc7F4AyzKqeDdKs9lrScgajmSjYl5vlMj0pFF7hhQbX63bFtm
GTw0AX0HGevxKKnVT/NjvCXBXKIlR/8AW0orQIoKFiYrYoMtcMUhqm80ZnYWLKpe
PhGXpCDVMS3saaUEToeLA6vnaU9Yx87Pq8VtxonXjdLISA7vl6amMQB2LSOGSBmc
dQiz0F237RWdMWzVe3BPfCl4lBT1+38Vc3YjemgOmh2EbrB5JSgqHMBqYzOCpRmh
H6N4q9e9OI2r1kD06Xc3QHsnR0AExPjRRTkrEo5TUwv/xQ0Xj2nxIC090gohXUSu
0XwLCY8b1qt4VUJtYW0trMMxtidXGYPpROgXh5YW0uacuQvgvnKrsiJA+KszsuGM
WXg5EeszvV1/porxKg03nFNZomkItUA+BQcMVRvychMVxkhYYnAxXcBjjod2Xx9/
9LphdZWBx74zwqTuTVZgTio9BNL9N66Ce0E2+wCQo5J43cCVJSK3n99iEUqDRKZe
/5DwKlQ03k0yna7oZNzkWdFwR/JaxbvGCZ3AOKc8IbE1dK0VjsF4gifOKYSY+0yx
atj7knzB1HfRWLLRnp4ni22wjqGPFUFdnJqpmUJ+zzF3WlQvda2A/3SC/LCjC37Q
0i4BT/0vgLphhTQ70exdd5NK4A7JYxZt5lWaRXoXv13Rx/YkYF4KB5J60Y3pBY88
3AAJg77tlr0DBDVPAP1HdazmTWh57VyDcoPITDvAO9x79lRHtCb8nXySe9EqWDXE
jhqja8Yx2wqjj4CsjJIeNtkeAt8s9lPeYNLJ8Kj/AuVr2RYCwBwLd4J1gtj0DDFI
cZqbbw+6lAx2ghaa0skrd5eHad1CTbIPpFG63vhgcXCvY0dJoRMXgN0sydN7iw1V
arUj7J2uAyJ3E2lNX26HsGL57O/1PhbCEiUqBbw2BFG38O838iMKhpDk/IyCdHnF
Cnmx1wcSxnunmkCZiNSZSdJxko+Nha9AVpi8UQCM6uTYhqIDvdf24MN3gAUg3IQX
AdO2V/pZ8Wjjaoo0kHpznSZCz0ykE5NUmq9GzzmLsDGXPRc9vc/sIDHnr9hSg4K5
6GsOwbiGIVM6cwyE6hPeI35KfSXNkC6My4QGa9UcsCsiPeC61m1gjvZyl4Gt2/xl
1m9JGFDrchPLzFWUf6UK6u2RAlKH0glY7OLocxij65qkGGYmMGd/1Hbe51jn0Emy
1LKClXh1kfrreoszVaouaT1YIwkKivsj5vp18ZffzlpZnM2DVZvBXc2XjtvoE3LC
GKfSHjBs4oe8xTldO1NQ3hKoOInHRKnE2oJobvB9ZgmOxgsksJT+S3ElRFaVJnta
tPWY8/1zTmNC/JgDgIGU7Ply3fnMSUzoc+VHyxtwuFqgkgFKSUKlDWg6D10iVYHb
9mD4ucBCRYAkBx1dxVxrrUxGPOOGF+OMA6snpXR1DPyGQwP1nA9JGuIeNA1AEOlv
fl+hKcLrLECAwhWBLvzlyAOWdCATYYY/RRkeRDXuaUcuGiACQaEHltvZ+tEzi7WO
YFxEyKP8qiI8ViNJggosxFhU1Y8uBArqjrfYaD+PaosGhYY84DHS5Q3VX9is2kNr
x2LrGI7UQMdTmBuPKQh9RQzr4DVrj0cnmFC7AGnLYbPIM8SGMTvOEy2b89Ab6U9O
mrh3O2TRv762WxXN2pbJgJkClCuo1Iwnkg7l1RuzwfGxPclLHzsbKLxBIifcdk1E
nL39lpp3dcTlGx2aNCfxDQNz+LeRExQOtwjXm6YkLTpbR42BNWAAc4e+ieCiK3DX
utjBnp3qiKODbLLbpP8rMsVDsShuMijlZIisVcZaPfMXlNY3O8EEuVSWJikIbswn
W0DkK0eQnkt5yHSPTdDwz7+cs6V16I+jzYwUocwevCTZv3X31MYzdhKy2k0TD4KW
e7WyCcxwvfpDhdFKH5+1UzrXm059cXtYZVTJUVgAB9lS4q2twhoCJBa8wwluldSV
pqbhDsCmIo+t6ICQlBgvIr/YGl96q4sip2Yw2OXj8mS0a7ANfNUvG8biqkXSuZGw
fN31gbredHWf4eM5lNPa0QRLiP/dJI8KdHV+0QItuZaI9eJNp7wgqs73jdBP9hTm
YZc97h6hOVIrif/BpDkfx4Z1+J9tqQLy6h3sZtZAF79oDrzjS3OB7JRsxqlA2O50
Q4rk+E5YLtDhlx9RFV7rNL0bTDmh/+VxNemu8J/Lp81vKN6J1j6KgptsGIRX79aD
p86Cjnt5SaztJHBayNTDkNP+l41AdOh/mNtUIn1/YQAbzIqD0WCFSp3gEzz2O243
sCKh7HVQ5XQYiND7fgUKUi9LxPBizZJiU4YEIonIHZIWYjx+GLvIW42ywRSolBYo
s0P7RNWPhL0rNA3lqfifPkGoYgV6eJSnRws7IoKMc64xPQ3+ObTClCA6bjhVCGIx
5sQ+fRp7sxYaLMCPcjLlCYnd/SI6KHOTO26cdKaWXRzt98f4dl6TEfJlPWtTHbBJ
pg31NWjxj7gDs6oMdQqhn000IUGhHXQ1TUNyiEUc8E94Y1jz8fXh/cZ8NMhRNyCP
I66btvkjg3qoYCsfvSucYwZLCwyif7O0OKoXKI1h1NqHUHMnwzbAHTsalTCrsf+q
kl9JK2we+/s2dIYhccoFztZTpybQRWxBbx0hMnYhtV7f+sLZUkrQeyfuKnq/eTnz
r+7FfLkXYBdlJvCKnnXG6BFMSTqmXm8LzhDai70ciWg7cjPx38hMSxMNQj19qcgQ
oU8aYAHNj3xqiJmn1S5dgcHN52Mc7RmNW5hGTt5VA9otSvfYsXpipGao67YH4+fN
wc+Uq9dgXNQO78wsrvnES2t5G4OE3BbOb9il3WrR8TjYnqfvi0lKtWfQ2WcVIEMZ
3xKvUOjzXdZ5PPsO4Gtjt0QbfV/onwUJLG7L6TxZbBlsHFXRAJyr+MoUTOyziX+j
NuV733VvF56Tl6HcGjpPPtLTqxAHLBZZ8Ft6s19V9TnAJyrrHV3Vtt2qiPZKKg1Z
OA6cm36bFOC/rkUSmb5xxvBRgtnyiFTXfEHt0OGJ70mYVlgJ7RuslRY1Sx3k9mmy
lD/zskRe8Irg9siCRkELbkxze7iTGD56EHRl6RLvABPC2KWpjE2ujd1RFICptSL2
v8cTZZnHJQ+1wC5xrqBui5nwzZgt/UcWonf4liPBDHcOS9MMOxzWvIO8miTcH2wX
tETtUbU73DuZMfLqygWOorGlf1E+wNaiTPm7bS+2omZakXb767gEuE8gLtpTkLHY
RDxWb8kiE5Kr0ugoQ3xbZbWQXmBlxDUb+w1SzbQW0uzYIf2Bc56ND1Vs3pIPL6/5
KE+bXvSNdTCiLClxXygLuqSWKJ/cr7a1Gcpg4oNuPUAVrdM6TbDts6Eoqiz/qxSy
Q3dB031G42uW80Nl0hIL4kC1Ua5st1XOK6nOSmTl9vU6TtmfEmqrtjwWhHOR4odM
CyfPfm+V6gJGEvp/tO4u5bnt24suThlQ3IrEYG+Eca+wELELqLuFsLfX2aBuCzeq
/OgHgcJEmAIXfThfx2U93T8jR2NwAZC5Tyq2DGloPRwWHowOXNGMUrTQe27k0ssu
PKybhFoew0ne/nnykDeTGfZWu2BznJLCoXQstWVP2Y8Z8jrGmS/BdYUu5/VTVlEZ
z6DpNxFQJBrsA3nUazkX3lXV3aK7qSWPriYYEBpjvWofKueK3amOULpBh2ZD3/ri
H7Bc9pL6LDzrgiyeyFbgBaia3lMnu49Fg6Y8fGIDDW2d6JyXarMaR5Z9+Psv72SI
10MpieIJcJb8HUqb3lxT5ocfDd0eSGmEFWbNXPhnEtPLVYw6mLES5ot/qt88CyG2
z+Hgha1wb/hrXeeouBRZEY8qZjDWGTMj2mZKLhptjMXGsNXrWYuzxCoDO3uGQ5cH
IeF3fkrHNZfN2HtvDJxlCntIwkPDKS/nidwM8Lons1yvJprAqzam18cGFnXM/1fW
f4aXUK63cbyaDpOZCebG8bRc31CDJ6WnmmBUxR8Y3ewysRgtRlNqIGP294gLUvgS
Ip0Wjq58qQnkPal4yVY1WeevlmgDa6pKVaZKEVO4EbCRSIAPszr0uxklm7BefwZw
jEC1RkcgInvoU+FjAppsfUUXmkrpSLbYrtvK0ltn5wBcFz9olJoP98kHHYUHBVOQ
fxZyPVCFzeIW+iBD2E2pEV+ussTv1icFUP5+/6LAQDmCx7bCBFgUo8tybX3bpzNp
Nnk6L6cGVXeE9Cvenc3oOph9TcVwIbjS4OTGbUfRRBqvGiQ+r6N5Nqjyy31c9gFr
qoKtxGspLihv89KOoxI3AFJQS5SDJUPXVMquX6jqQfD8EPrdvpGNJSM/vOiXdV1y
KE04mMo3f0EJou0X1RJHMxnCXoeyZJDzPh73t7Pm5v96l2rbbgkRIe0U+nO8f7mS
CQHg/apjHQ6LFJicO4fCeoLkgMnctxYJKf3e9shDu7ZeS5Ik58mrNrX9KUsB8GsO
W8cnLrVpEf2rTr4KNDQVCVSY75A+cJCt820jVNMQRUBtzJp8yi3gHEFMV04y2iV4
fVVQ6dHOD07ROgtOXUAx26FiIKTB5STKwoGnAKYP9haE61FhrOkMVHL/a0bsWWAn
uVQSEQfPAfZXOpuf/L5VV9oZf8U6qOTKUt87Z6tR2QPu/abetamJ5rKP21DttPmd
MiQrkZ5NzmHRqBX5D4QbjA49pEQHEux7dnjhdwCfpGOUUrhyMLnZGaJ81JPypPuo
DtrqnLurwlQIHYt38rBSAwivx9E+FmOeDZ4N6CQhDOiSxaDVc1IAUtOCNE1AyiXG
Qe8gYFS5Hj70fxSxDJldeoqnzrR9LLtZyIVpH90nRLgyI+1yONxgQn0pzpNIGWiq
C8szeAp1njQsWccvjytiTDYMZ6lCJa/+yhhCukO+8qFGp6FgFYMatlvdmXE+QFwn
nm2Ge3v9exkWXIfR1LqPfYk6SK2GZfWEEhGmEUEcSzrMF++1IqGwIKZtJ1ghq0M0
uvrPTQV94dvYmCWRUwYfGf4xZKvon1kWyozVrUZCauh3dQw5PArZMZ4MRcGrvIMA
nWtlmJgW1vSWRMN93poDojKmphpS+mfNlMZXKDXMW5vFAXh84QEoy/knmyiYjQz6
LbvGgRqrG9VLLlm4r9oRIAtbpGudOd8hFuiRE2AyNTHGTN56V6XzRK3MODcOzt2e
mcXR+sLS+ZZUN6HAhc2cNcdFHDXBVNyWOfi7aaZxWegdENr+VmEvuwIgtOcDUNuj
8ufSWovu6F7+vxUBP7b5G2bAGPoiznWXnuv7Y1xCHO8GPetO+YaJrXUQjpXAhuJ5
PH+cpYL4zuBq6cFk+hbv9ZyiQ3EbicSOFBwE5ndFMu0xQJay1TfYnJU0JZDX+8s4
hxPeDOeThZAalEn1gY4x4H9lya+6QvMjTemloyrDqma6OQc5KXL6NdOlFys41R6O
yXjmPZOZZY7u7NXCFMomKzlclfbRezQ1+LILG00JeFM90pHoNc5tlw1ONW/ZIY5N
tnZTltSpV+Mrgej+471lMqkCnx1Cfav7Wb80gtQUfFtFi6hWn3m5Ti/rAvJCv48y
mmpY6DLsRmz1T0v4fjefHMaKP43yZectIn56vTlzjysJOpRRjwquaq/7xirehXUz
XLQzhrkDCK3MD9nkiUV/V7N1Qs3U1jHzGSEU3WFbn5CE6evj8cOi/YDSZnigRKNG
5yyN29KlmPNM5e3UXHjTQ93Lo5W8IFch1FsvDH+iU6zIy1uTvnoIbWzw65k3ssO7
1bnw3dyhCwhClVstRGStqEq6MXi+Qhdh36U94bW9OAc89LjyAiNrp67D5JiWW8wc
KAFIvwB7Sw11auQ+VyCmbO+d72rZJethrwBsHOD12SHNWyAcB+rmD0iERJFhrBcu
+FZFfcxwG7ugh76l9iwPdEoCS6TsM1at7WD9aMECsjuPSrhH/OBQpduHB7i6bpvX
3vgpvAeglbABXDvEoL2oIhUpCqy7LnRdxyYd/cUHX+0QvHEESgeWaD/CLRgI6XAE
OPPlj7AS4162BjW3hM28U9/yfaOHxokxD1HcPpaZnGgj4mAvXK1Zo/+mNO4lSLc3
y9SW7i1E9C4IlLD3QPAIQPnInHQkptJnx8Lo1y/1diUK8kmQCGXb3JQxnKAL3lN1
C+ZwScoGZ0nd8AD27QE1uVHlX3+sBJeQuOHJ53qEP76djjEfSt0NyavKLLPnJRIy
XuRia62FVAN5NKraGBqs5kOiEX92Gh5S/x54dOXzJs9aooBsqCvd0oOPahAMoxP8
SCFUysIfSq04Hve9Tw0I5xZuh2ycxzs1tTmQpmN0Arr1/2fRI+D/4UjAujJ9zQ+/
5QdozSuhm+c7Qeojka5bP/8VoCVXAJAwTJ/d359gx+96WpVaosfXndwFbMC7SayP
wQbdPo4OmXUXkptGc69+z4JJRZtgvHUZiDr66jpNzwL7y40x7Hcwvvr3RZJADxZr
k98QGj9ac6RO7WtoJAORHLmxt9adTbVVxHRYguCVNeHg2A9cgjePT1cN7l1m0oka
5ITqhtPQWu3TEYD1gOPZ1nfWvpMNNHu0suhAlhSeQ9nS+VDaladL2h+8gJycUAc9
synDEmcX2ck3vyWFvQS6O7lji0IvnJXt0+5aKm+1+pw2nJZxYdHZdEpeWT4Sv2XV
ojWm3fANsOBo+6yzeT98u868PNjU0WXv32JV24fUyhT8rOKZxy+OLULSse2rUgrG
KcvPL5l/+zVVATZ6vtvcul38MBWr28DsI9vKgVqLkEmf1Nkeg5M1jr/bFiETP4RG
fTr7MpasatMEr1M2QwG447k82/trcz5Ktz2xuxvBO4ccG+tpUHpN+1qU5j/PZ46g
mo5ZyqZV7mDshCX59WUvfVTXJybmn2dE5UDOPszT4PPa4QjgWMOojPSIm4MakSaQ
YscWQZjvqV4QXON7iMAhXdjaj8OK3bcBhdD2ojICFwlT/2nJZSCuHukcW2dwZo1X
Bd8gemuRLqEOpwJLLLFSoW4BT6Sd0F8dYe72856pxCzWu0/wYQSdgxY8AI7x/rGR
QBrIA8aTQP+mXJaWYIe73caxkhyxRjYyT25YP9XbIAIpMyQobSV3ltlVWQ4Z+vNr
wuBrcdovvAGEPbcWfKVq+ec5jnWDGXXcrft32i7mDvnG601/sg+vNhpJmEXnermh
j2/B/pLX0r7rA8NIfXzjkfJEQdp5Udiezp0KydAi+3+OLGO8U7GlVVJGRQxtqdr2
V7jGe/QL53IDSeMS3t3hRyvkVzoGIhup849PdMz1V8jNICzSiL9EK9Vq0kfWNR3e
TdMIyGONNzjMu9U1ehTLo16BP4fwYHD5BhhlYXtSqa7tcrYGxqsfHy6Ua5AtDmr2
KDe+yWlU2IvDf8G3Qbl6Q1OGeqaNvY5UDHnk8gcCGBR835FWxtkVdSs/HElmOSz4
RBejr709DvI/x02i9uoc3W1nA2ixBnncagCsOtDvs+EAmOX6ZIau3BtCxykLnw8l
B3x8bAZ9DzlQ4uZzfHA9H5JsnVW3Ybevp6BxJGrAQHcPkXhTMmL+c+wHkbk8Tbbn
d/GhLX5QWYOeobJhFUi72fC8V6DFEyJ1nz1SnmkQBnlhT7L+wCVJT3ADZ5N2Sk88
DMW1MJwHmIY5Gor6yOMg+X2xI+nNkjT+TDqxMJxgmzWRpwY3oshi/n7brZjz3HIE
FU3EkZvGQKR5Px4nVjbPElCOQN/Oa0yS02FyhHV8/XtBisM3tT0Z0FRUWEETHNd1
Gbbm/g/P3oJ40tOAIIirdJGqH3adM+4lxIiRFRG880/bXN7jo24glRNfb+/DPRb5
85Zgr9lYxIVx4apwATkq2a7sTO6AK13SbU+L/YBXAHqe52phHcb4ebkr1rOnZRo7
cp7/PGhvFhiQAhr3yGPhRy3LH4oBe8+x2EeJGmrHDKuR5HBEIS4x54BnbrOJhJSi
jFC6Y8iPlHTJTg2hguiEM3ubR7MjzPPWxHf+e+XXEB30F4nltE7DZAy5u0nNPbY5
klWWvKypNIvRrGdu2J5rOsrSUR1mfBiE925mulx7W40keqdiNzooneri2pTRYvnG
5Xuo9DDdVfq1FfK0i/uh+VEW4eBHp8/gXUbjjmH+lYR3wW6b5bVxDWTy1lmb1PeE
u1h2DTnpLgJXl0hQfCmrcKRQ8WUF6yO+pj/cENzDcgt4txc7EUb/v7h7veExUE7I
4eIB4E8/0DbSr6r8ptceHIJPvC0bs/eG4+Ysx2G/cZUWfONlu6q7SVIEfIqnu+k+
9BZkA9DnJRL39PbbdvFFmEeOgl30Y4t8huuLJbYUl3z3A0TOmdlDFw83ZaRx2SqC
8ja+hj8z7ykoVFwPSAXZzpWdFUW0tfNIN8jkXyuXybvVQJ40ClQBR/QJWF8tegtQ
jF5L9LrU0JiQdPfnXQFvoCKrwOp4J7sFGe2nSCoYVvAFWsBRNecETEoSxF2KS15t
q6utQR3SMK30TV9qoso91SPJJc3stmOzjb9SwmoNHGhtCq07A+q6JrUlH5WvBQ8A
cy3uci0nwCF59K4DTUILQNbyK7ojZWuX/+b2tmSLGTtQaYsmN/zu813N00kMC1FV
EoYVxAqHa85Zt6HpZBqknDk7xsHc++pVEiHoboTWK+E7n0MEp+AWaIy6VeiYDSWn
GV4PR4ki+jKjcN9VdwnNaj8QnE3JdEII5uhfo29Nyd+UJ8vDKli29xbvgT1SspRk
CZofOsVW+ARlwz3fbbyt7MvpnlSAoSCEk1RFh9Gj7gRyYPs9gC6vfioVzDZXVj9g
9LUtBhIbKKzcgUmwv/osvv2jh3L9uivrAAR0hDvBbFYHvEeDjKgYPgpzE47z5kLH
O3u95XnL+xg8pFMxYdAasWBkaGyzPj8csXS+tNhy9UhvnXL707vB1MqRdN6C9IjU
Qe3TKNf7mZptg4MCoCp/664lR78tzdUqEc5uTGuRiKZadFm/QuuliHduQJgevxxi
uMHeZzTXBAsnev6bw03hagOHLM/9fO0/dLaBlCN5FXKW2IpllTXiMzPQLnA6L+BR
UClSksuMBd6atRqfuIy0DoLzzPg7oPOE0++VvYbgCvh9vV+ZXwHTKVpTKH8MLmZw
/wOAoJmb6Ylwb8+u80R5zLjsKHrozGbMVk6iJzgOk0sG6LO9wC4v5xJzYm6MApEf
dAPwnlqbRwNYx7SrtUXZqNJNLp9EX52mYkujj6VRu+ZCpTfyoskG/hDJtUhY48fz
p7SkKlK172fiUwRJFgkIAJtAHXVVp/iBsykGfukAbwFuHlSn7Cs/PEG1Y8aQjhrL
moeiAEHLpFmUT9kyfcdHp0sLmaid7R7yvY3z56WSAoJnWDDa+B9/2V12SP8OhWC1
YCC4P4yJjE9qXUxKrhXMBbp1ip9z9JAHNEcxDTYR2NTezH5EO2J5fWVBca21jMIF
FZSw7G0qKy84QTQ/RaRVn0uZ6HPlPTrXJ1ulLiiWhYP3khLrwXo7TuhudSb2nJjw
2EJ+DBvzFZgmt4fF4dCL1HGYcLGMC4D8qb2ALAqK3mbzCq7kQ0YmT3Vlp2Hfd2+R
UW2Kq0Fqv907N6mJfl5bRkP6BhXsCNhtpGiHir6UZUN4GbXzzqL14AI5DHDo9l/b
337W59KcgyqThhLUSZd3t0DgMI1qtrPAdPiEkVcPTiGDmrJ7EIFYpif/21cls+hd
7AQCBMMUb2gklMKnPECZanX6q2aG9ALW6QzcX33Kn7HydsezbIJvroqDo47dwqBt
KZiUK1XhO4wokD1UyIxOnyT+VefAWFb87Jp373w68IjL4IjhBJXp0JwxkB64X6AF
RTthr6k1fdnN4ian7KIDB07muHYWWFM769lGOQ9kSJAh6bX+FoBOV+7XxO3f7Nie
/Ur66Lw0YeyI9qLaqmNzi3RezbTFnwsEHgSHVugKqe6eTX/ESm1QM7nDGyhLsCsF
KcoinlNTB7wFg2XTPFrQZMTlxEBFFxlTlv9OOeT9F/NLnbAWMADnNIH6OJ0kBgGz
MeA1+XD7OkihXRmHSN6Ipfh1TiC9pAo+QPuxgF/ZzLGsIwZC8Kk+hruEdh7lwz67
FKGtJradA0jANzlJd5mr6HrzmqxOERpkuoUCJhLJwXONO/4pyqZxtRiG0UFvjl0u
ThRYCQyVEaJI5mCMb+76emg7Kp7AtOQFmj1j1JBi8NO/FJKFbzcd/aoT4KqO3u4f
Wq2N7Ob4LFcFO9Sq9SuvRuvz8Gk6+uFGKbHqfq9jfGPrQdk2p1LhUcsRr4i6fBPY
X3RvLxPtExI+KjqqYfVRPLfxx0GOqVIEsW3Yo2j+FZuQIpi7CnaqyJGrDv6bG2Ac
IgrmIVFcM7NgHG+gbrJlSeeLRr0I9Lc/dfmRHF6OfI5bFdj+RT/wOauqcrdgIVQr
RwdkldDFxmM7KxBwpoQnEP/t1ETQ1fNM6c6/gzGE8MhHxQNN5kHxmKMNWBZ8VLOY
fKDOwfksMTC3jJIqb8O4rKYMFi9PdrsO/XE1kLJd/Gq7OynySxgr7L5k7FBCCjVj
w30FExTYUGU7iu+IF2I4RpLzVMKcIzr0YSgFBi1kPzfTVQjl9tAag1wlNe2T2TVB
UM9sNNDykfcEV5Qyb6tjVwjw7ls9mi26iP7hYxg9rXFWDFpgq071YaduRDkxHmYS
bZfQoZBnENS4U4uzlyFsR1FO71aAx4Y3TIYcqx5DuTfPXBnTO2P6R/xwb+QOYH0o
qlfkkJF53COmSCQ835Q3o5xQJ/FQh1wTu/BxlHxY2AvHwM/cMQF/gO/cpq/fUMH5
Ffbvj+27wSj8ts1hPnp44+cNz1FJUNT9ADCKBrBqI2cWKJo3UQOjsuNTCRqQW4SR
84j/cIDDx8OCzLYQaFITkZZ5p47zS05tR8POhDMnYXSckD3EzWNN6ph4kXa5/XxA
YPDWVMELgi0gM68uN87jTJl9AxMzmEBFxus5KjhebcnlW0K3tm/VVelfaDZLZxPR
5j/qP7GfFV7BFOKgaAeGwW6pyungWut2DlSdqhjHlACNBBErHnd4XKQahdE2bOF/
GXzqYFp3EYgh6B8PtBe7zsc6EXUZleVuouOjXW0CVnvCO3O3s4Q7DF5F7zcmfYeV
SRO8DtXrZnx5bL0bkRakGDnmfP/t3JWplx6U5qe8HOuQay3VATa0YhC5hYyU6eHU
ytVQAPvJvRPesvVlDdN8eKo3IxIeUACiKoD069CHxhXNg4RFh8qtE0yQqpdGQlVu
gQGa9VvVrcpkuevVGBkBRQbTEq5YW5zZDJdujcfk5x5+u5FDuGWYEs7jFuKVOqm8
TbcFhDbXopxtiV2dCfqCJpQPACDyVMIwW97ePcdb9lDC/4HUDojkAyta3czWrdy5
Oyg8HTgowklM9BMd5feqa2iyBUHx2nI11eJL5y93o6ey9DO+HGtoQd7G4956ptwF
+FnVoqzqI25fHrcjVzde5lzWTcrBHVatdI2hI+yfnUDSQuOeVIV8z/eiv/IY4No3
BdZuzJADMIVJkIcb/mbOIhbfQefM/T11zhxo730Zza1kNnVZsrtGpfjDZMNd3vTC
2CnHEMOWHrHj4UG2WoABGoU/CJbXFCbBS9sfBRwYfdfUwIsqCoIXhpyyHVZ6jO4B
PMS5tY3UQ/OWmOENNRFNOjWtEWx5BqZQzNE6Nk6MaaUdIwofXMQLQlzi0RycY5fH
lojieq/GGVZCmBIfp4td7yfy2AgAIHKyP0iteDCBG1zNPkWsJYctgj9htd/d3bHb
8fFtbFkLNxHPlGYqfG91hkJOZzcUyILuq5jC6Gh1b12SWoojKjPommPK9dwEZMZE
f2eKzEAy27vr62CnsPMs23cge9bIStHigJ69gCF/LkLYIGLy+3Ksyfku6JRh31m6
9jtGhook6p2waBmAggWIlzjGEqCG+I1oC83lWuxhjcoK3jFEV2bTlwgOAYRnT+iP
WJyyPBr54b9r7vw7gO04ec6OAR6IKJ2J2fJBcT03RxfAA0b3n7zZ4BXkM80NKn/K
eXTok5xf7jPCnBW65NKffjE7igCa9Zgwys0uk9A6uJbGanb+mKgILVWwcivWFCDa
ErxLDJAQ9FLlI3khmJrntcFxUkRhSfN05c/V5+JiTttzIwKi40VO4GEKNRTeRQM6
GmCwkSvl0N8nFcHXqe2f/i4QwJag9bXNTnVy7xBV9S9MUeJ4SZtC1Rp81jSsf52c
nHNKdT3isf6h+d22hfah3WykrHPFvz25mL/Ok1SByQV1GscmBfAFE5ih78I3jTCO
rtWskFnk69woFvGfdHN6b+8XL/ZiJe56aJptT4aRvgyduKl1omD5E+TtyBDKaCPy
9Dor+az3b2hzKP3OHL4Z0Ja4T8vdGFjU14i8DNTdFwvhMwasuQyQ4MOVqTs8RT3y
X7dfvCsyv6TowlwNGKXGRNid2inizsYMCdSK3IL6Hsuvuye5Y5nyfIQ0yh3PjV/5
GuwcgKU75I5UoQzIPLiXcVIyBuJUzPe7LUE21zqj6BZxc3joU8OqbyClbb5Z9BzU
zcudh2HBNlojAn8iAUxGCoq/FX5gXZKHjjtnmMIUfl5O0k8dpCelQG8eQ8kL5xWe
LrFcP7oY1BE8Nt7QuI2U3FYKjAZVy+hCJwfZcwEbw+cn7EvlZ6xMSuY9CdEsTTsO
JSSC2pwaT3gh8GnXCQBTiRA0IbR1f1EE3h3rJbZB4MOjH/2wqvJ6SqAxY+UBp2Ju
bHTpfV67qUsbIfZx9PGwT8mcXAOCz8xuJKlk/rZbdw2pYe3bHzdFbhhXn90s4uHo
yjccVRsMBIpOgN0dEV37fg+g51ooi/PN6GcBUxASSqQ07ZK75rU7Lg0+2YU1AJ1f
dDBMxV//t78gbkpEvvPnY2e/c9MhmK0GoALYjKnqZ+bRZSJx00XYBtDnDY4GCyI/
K5Tc10B66MNmizbUkmK+ZGVNMDb13JAAvnYwEZzWP2wlC13YqTIVDBBWru2O4Rp6
umNkSZmaFAB+2coL763IsOGgoY5rIhXDGU9a+EK3gSlnkIAunwgvH5u1Fn99lTbQ
4K1TECw9BEzsoxHfENeSzgfdZkx70zCTrFeOllo4Vv1veGfU930Gr0ZFbHT5NsGw
WnSGGX2K7PexJ+ikR1356nJW0PO3B/4Yej8FuDmaie7k3zhncbrKkD9Iidiu/sTA
qj4SNgfwCzoL8kVGdf1XpDfTrVcDzFBGXN3B83QGnC6S4vCboLZ8ChZXK2XYMKE0
6pfxJc35VnbIUO6pbob8SbWGn1Fqy3xMBoIZtCBB3Ncopzmn/u+BVNLlPoVyVgrr
RkcUW8MmZUaHntPsp2c4p4qAHHZlhZ1xnnFvfozyNEmDBBJlEzVZfA1PkA7ct7KX
yxmtwWAnXoRbRuPo8LY3jfhtngzwdiU1miPov/GgTbxa3hEXzxjfxJmnyfZTcK1U
Y9Ay6SEgaZq+GNC5E3/8st8PYla2eG9Bc9pstIOG1dmytCuYaGbpJiN3qAuYPHwc
iXNwCgi+hM9n4a54k0v3UPscKHz0s3amPn00idZAQhhqFc9iA7HqNMnwihdzIpSt
drE3DPhFqxBjK/BtoVsIBWz693KNBuCWxhJF6P0R1I3nJxMyGe0tRKDTqvyBFZrq
0BgUuk76rT0viZtYTba+u6U2dAEbo0wpvfbky/chLFJgC9N14DYQTOS8gXPbA3Yu
fTCO3SVAwy23IAtN9WUQvDKQApAJ4JDPJGup55wz5B1FI31qJSSWdgBk4Oa6+RC1
iUbvQhUM+jjgABHCf7pFVclkVbYiCGIJvrYge4xw2SKNKgAuar9ZCcI4n15vVuat
pXSvBALr5kcUDIMc7Gw8nuDJ/GrvksR/hwtAWMHaZwsKmdTn9DlMEyGK+ZL9KKsz
0S2WCIVrNH/3DflrwsaGNqVAUl1U4Vlx1zGtWNbddEY6dDoCwisdR6uvB3GCwnJv
TR5MG37mz0vjUyZrhH/tQhjfhA8D243yGOHi87U+xtR5+qX/GAVlLfhEd2BkDB3T
r9AC03tuqVAX2MJ3BNOZWbSGoFdphbF1FDkivHLNeDlUYufAtElTYZjvIkzC9ETo
z2OBXX2BnEapHgns6PzFhmyhA131GPWy03L2HchlA158fzBVWoxOhqZsBUQXhHoT
sPqB39Ry3IywDZlzmrofErllWbzpulhzao1wZVoNDLb6/nbUtduoa3acvff1UIEX
neGQGXtyDb4vOVl09vFyVPG0Oercs92QULotiv9Fm6M8ZNwh0jemQCHIsfGCJ3zZ
7YZFjsqIVFbUT7cvRhcwjhQRMWrtVK6LNsJgdKFOQp1+cUeRs/0PLBSI8DDyAtms
8SW6IZRO9lkHjK7kVZH+NiE/coNCMroBi53tXAm+kEGaxqCDn/hgFj3Rj/jLf3ig
VSVqzVSnJdzdDvESdMpjhIj5hxJR/o8n8IDpKl+cwDJEH0bapqwCiZWh/kKBe80H
NuZWdl9iESstZposfT1eFb28mlMG2B+jpon448qDkZomU6+StiMm1qEsfLJzTsja
E1bY5iothHgC9ZC/lnUmc/9DTJ9GIzmOMtQrVdDNZae7efcSNdQk8by1Jlz2wvDI
V1CsNWfH8X5xEnSS6TlNg6oSpN/xWd9tTi//fKr70rud9sB0rLMrYg6nZGUVrjbE
0TA1hR4cJlQZLQIR4SDKIivvduP23wgF9ZeB4RKXEw9tqI9uXN3uXpIvWocAVLvX
5Z691nkM3Z89honbydmZ7/yxjx+nsGLrHK5W3aTPSsRTNvBQY40VfkaQREiNhXyh
r+ev+4zrPvUkeixERRafqkzDRKaXWv+k+51cUv61sLmiaMIxIBYdQbugHyVsmbKN
34e4+n3r5BRZ8GwcbMuVMnrIdbQHPq0JDO7/Su9hZ9QMvc49N40a9lqDslnznYQ8
gwWRmIXbJ5nBfSvUjSu3Yql4Tgwif87LuwxRiygAWI48hUGFsv/HYW0bh6pJ/jvP
sZBqtJD7ZT/UuxecGpPCbAQFNUBEKRflP8e1Lm1ZIeGgVqSJcYPRdUsnLNdgP47D
xX0DCnPKqQvRPtpgeW5EDr0fFa020BStHNHN7Re+g4xH4ZdREl1eJu1eRLlE1hbl
yC8bJGheO8vngd69R5o6Ohbq5BToNT0EblMDR07klQn6RYmnIVZ8C9Ujf/Y3QLUp
niRUDck0Uf8MF14OTQK7YHLP2uDCXmd0pYe+BlQWINxcgCGtwQe1z9Z0lFeLtbYd
uuHc2frzYk6nHU0op29cEDjyz7/pU8iycLrp733VCFChuj3zNg2v0ukS7DT/TsqY
HlD/ltnyvPeZnsJetZicUCq3Q9PCN/a9Mkxz0FgXrhJMtXWX31rCwhlrTmjemHgQ
UyQQt0zLX86tiuxBUhL2XjYiaymrBaqtEZ/CzpBQCy0aYQBGMnf/ZhMZe+y0DXDW
qiL1Omc6oANJwnOHMQWKwoGSv62RuW6c7TohJJlB7sbIH5u2KuQ7zrm4n4nUpsa5
NxwDGbpmYqJQvh0FIFZZynpGR83q0M+zw7dwIriLnGOK4vCcZAYa+SHuU7c+A2Fu
Gn098+AKgIL4EWpFIjReQmif5ahBRu9YSbiTwYWpDJROunJvs3vW9K3lu+6REeoV
r9JTGk8DzFt+4LHIMfLiI2UMFREkXjf3NqohqIO7U1YYZtVll3jbLt5UjJe4Xk+G
bZ9a8KwuYunesOZYm56SK3G57w8ZXSSaWZeHkCkdjhOd8PKO+ZxabdNvLHr88hms
qZz06mFtcW3NHVxilnmPq7T/1yHaAgKgHp8D33KRZXHZN8h8cpQmv1wJfwKvb6aj
xZhmR+HupDFEP61F5qz+I1KWdAmcbW0oLMY9cmd2hR4CDxs6wgU9xWFwqwmLu5O6
XIKDgsj/Jq+eBelYJc4drLzw3x+LPEEUHJybPhS9NYLzbMGZMuh70hZP85SJv5+M
Py0BKbXmdHWKrqsK6B+Li+3nMWs2Eh+pvurJj3r3FSmZ83ZYF5mLTtPPag56PsPJ
2nPfHd4EoKYrO7Of/Gbv4wqNzl9ifpVOIivRhWhpUEYpe5uvbyHK+yDy8griArgk
3P9VMMo4AljcmyEJuSugJKRGIO6CSKrM74UMcQXSCg3AIlj5EcvuW63D135OJF+i
oTjEyKSKfL8QlxMAAw6XsLlzCVOJLRplFjXXseGpMhib927zqjkuOdvMmzz88lq/
wxMIMdjFU2wnhg+nzmx/5/nA8/o883tJ3KfvSCHrk3v2ig2BumX0H3xZ3p3moI2Z
gi7xxxyzizdh5w1wjZdCyQ7RA5036ZCDo9pgTlfq+k1HuwH8BZqM3+nkTv4h0Yyx
biHVa9go1L7zrSRkU46/wud1gq1IK/ttQoTuyWtY3JOO7+7QK5iguauLBC4m6iEQ
EscutL/tLMYpd73DzvVELYd/e2aYyTd30ya6WzJZUnyAEPHqcN/7/lcuq0cGXfFM
2NDnISPpTzPG9oF+ZJkJJ91LI8UnGvXJYJJQt/QbP46I6RXP+NHDvIoOtixNDhPw
/YJhvcLG/G9Q1L6PIm9V55QbOrVYJYPFceEvN08B87lxMJEL6AQv7bAJ2ismvJla
gtXfuy+HC9s+lekuKamQmRj5IokoNclYpoAgf00ALWg9W67X9daZww44wQpVDaGg
wa1eEeS96OYDlcUusO8fi+GR0ph+R6HyO3LShP22Db4zMPjMuJbpEBRR1cwJEoIz
LJKeDDskF7bQA1SHzXDLJ8eLONLzAyxWvV/k5Levi9uPitFNh0PI5oRvehE9F/WR
edevdWMAdKByTkH3eWrme8x9QwGjYOjOekgwqDsozjjlL6lXW7uPhw/m2II3dQDf
YDzvk/S4cyPMJR1kmOSKsa6dXbtz+pzo6jispmUrWP4vHorlILr2FalaiK2QSNEc
qNBEKwz8fxoqCQR6bbefFT1olVlATlQhgZj6UiB8pbiJK144EiL4J7eClPICl8BZ
g3hQNKSnN9rWm9qE7g0dWyS8MJyFL+6lGZ7Gh9PfiKvYy6Sab8S1GqGUoH0JH2CD
34Nd1G26RXM2bH0UhqlbBRShO04U5O5g3oo7aFqbFxePXo4jBpzn8ZatnbYM6RTa
koBvjChcVyciCX2MhvcI33t1WTnp6DFZGOYjw7Axd9NAulhH+jWEZkhMQOr/Of4u
LQY5EDEy54evl1uLBRKNrf7CL6RtI3Jd6dMh3HC4AKqgjci6Gdzz/M7C8ngrU2ex
j03+WEpWU0gXFXBFT6zNvBz2K5te3DixO8FW0FnbtYnEZkdoTePZRein+lxye1gz
UAFBnbfUO3iCTZXKhisZyjricTBur4QkT7A2Vz7SpsNq0qr1tfhcw+iAXLK0yJyQ
u+zvGToRDldpvuGqx5gczIKpF15nnCuLJ6ReZElx5cT4YEBMcvbbXoKqtZWC14d8
HtxX99mf+UiOqMLvF1hdXF06bwp0ChPjWbQZQICh9FpW0bdNG8UKOe1o/trZMIUp
GE/TsfGOYQLRRjTask5I9YY196pO5I1sxZQ9+9/c9F1U9SLLhrLDxJTyG6W9DphC
FY7ZG+1OXsL+XWMpHqYi0TIxJJdZ/HAw3VqZJG8njXSsw3oy0FVBC9KqGnOjVwu6
P9BOR+vQMzUVehmmdtfZLEmLqfzygJhbkEPBky9eLzquwdh1P+v7T8Jn2zPfehdt
t1pV9FXUuVqMskvUjl5MSjwvVrPOLsJ1i3tK38fK7Hoa6szCojhjdcDwROnr3B7f
JSbyeoRBT+HOkTSy6uY8Se8S49S+a+qW2Mr85qMYaQBROR1ZFmpwN7tZIYTAMAhH
hGbPPjTnFnoH4FFKfcGasfVkofOLjj2SSgOr2hRPmiNEl2MosdJgubvt0Q+jFelX
3rnLbBjuZ2JfqR83v3BfjDgR3sWUB6+WMPz8hLHN6VlSa+JmFFiXif0HadI5+wqP
zsUz8FLxs9BcolFMkayEPx7yQOzxTU0H0UhWYyrziPvEkOg5ACWnA6keNX/vPURD
CZnjpjPgvGK/+gsC6T2rHpGYaiBj+mqz58kJEZ3Ltlq7a6vNAjqekcL5tvFVJ8TT
LDQHRQdoHc5SHSsSMh91bx0qmWhnajP+kiQaL6yg1NHZ69JAli3y6YuCZ3ahLMDo
DQvtPx+pVHq0zyu2+fpkBFAqWL+MflzxZIru0TAMZC531cCrcLsLEpV4hP5YYz6v
yMn/kgF+YuC3x6Zj4na66qWQ21h35BKIiquRdYRxDb+5ODwv3k0kkB5gK2sgrRBI
fNOzzFHLc2ozWmE74DuA6z7D3SAGjifLGecHu6hkER0kTmi9hsxRYK80/WwbsxAb
aV8cW/ot/mLzMp1nz5jVoVULts47oLea6cP1qDPA62Qw8vJ3FIHTh5eHSWlcd79X
H+6msru50rZjwP0Hjxdh6NmTXeIt4B3rf5DXdpplMoA4NMi4o5qgbhCGDwhVS+mv
3VXCN3I/fqD1rN/ADhcZ0KynVdI8xCGpREp31hdRxqp1GOODTsNUnZ7CDrmv1miC
fQjsVnPXMaQdFpQznMocaEYZkAiDXssdDMLiur52B5AoFnZEy+x5NQ5iLIaELmze
8JxF6PE8Gx/dpEpFQbdHtE7/y2MGCjJ+Px8eNFz8+65oj3fD2EOWLT3zYoDRqbTr
bFvC/KrnxufWrg09q7eXbWCPvj5PID34NTUaWwSb1j8Vo6PC5+YKu3GPa4iXhqdS
BrhUHeS1Kjpe3909m2zq5IARZ/w8RttHUnE/Sp2ophtMAXT4+DtCzi7tArZDDszF
+KKSioSH0Qmq7WR36bOr/vRj9iWkfW5SgMw6O/A421fLSEoGkh0GFUOzUUmr489m
mG9hVUGwyfvmWr9tNOBBCkXavfRiholXJNnGzUyYdAw0ZERJnKbXl3TQ9gD3WIij
eQOw7C0zLkd6tVs2Ud/xMrz/eXxe94XMUT/VBMqtD6xWVeeQAznpgrS635XsMyX2
6qYdF8qHtvvc51pf2XKtV5sQ1seIAylN07DfHXlC+BhLqzY27saSucHFSfpU/15T
KPkrtFanWdVqhHzZvmctEkU/Rn9bs2OUJuXKpy7SJfXQdGDTzuM59sSvQceUHCne
pGnGTUXvsAP8EwOusBKFDnnVI0nuTS8m9JfJWQxm3vnbxpE9GYwfaDXLkg3sUXkP
1vW+Gm+S879N8FYT1c+5Y7U0iJ0e7qs3Gt530J8zPatgzaZdbQ/Zv/GLRc05JT8b
SMAJymb3pQDXVq499AWziZkOzlakjb2NPQv9tfYg/+K3zdZ/c66ve7Uv1ERz2PwH
zfvOKk6MJVJy21ugomjWYNR2Fkmu8rsn10d/62lsdgkh83CqvOUQ0Tez0CESsok2
AcXIWqxXFYHIPAdXsiBF1FWHaIacJP+94NjHvRr84Y6eAcdBSM70QCpoq0Pn7WB9
Bflns1bDFsDEixJwtLbrGTEOcu8T7H4P5ZQlSWnJ9pg5dhX/axKF66RQyQTXabeq
fJlYctMfKt6oGQvqsnWZxYbrJemZXC1HdhVIVMNTLeWIDRTbc7fNLNX7AS3Mbd0V
O6spsbA7/xEzWILFycEPCEIvgWG9PlaK+tRH7R6p2epi4g2hPj03s86L6Oj1tyWU
U9bTJmINKk6NIoQvgO2RM6SSQwjm/1ZThWmeweeXWFfGNOWzuZ/qpIN9D1RxDFT0
J1/QsMgAPywn1ZFunq1lT3LALUOVH6kYowY+OaHWphM3nfM1PFTDVWwiI3pHUvBr
vFbOakDsIrcC3sqrO3MBr+KhDC6XJYQGv0jXZdDL+yrCwORFWaEN1884762NYgsc
9HwO65X5nUnx/GgfbJ7f1mNdfGZka3/Z89xClcf1gwiDpdm+B/vjtfNTjRSYYzej
7iW7FhkLnMhcjtWR4mZa17HT2hKl/Gidv8SEeV+YG16bp+9k30HZc6zNJlx4G22M
STrA80urIgrzJhVvAPmNdzA9LIPdDiAKt6RVFR8lhLlNPSkUiJ1Asrjy7GcxveHV
glj7YgfIU8IXBoFAB5do9vDwmxd0P3ARJfi4dGmPioEH0/1OfT26+Gahlp8m12IY
9l1rabpogfO3nnZbFxzf0kojJYBtAJiNfyHbkn+rbyGACDRemvLlwnDMzEn5cxnm
bV8qoeKqQNL5wYoxcFjF2ZZmK+FImTrQ/v0KbaK9bRN3GKSTf8AX10Mc1VscBfD6
l36dK6TUYKfutdNkr8WjyiZHQ9qFmfBsFiGYqPLFDCXNlb7BTWBjVPXyt4a40bcR
Hkkb7e2xqOx7yK1Fi2S5N+ij/LkheEmfVJqiWqfR34fn/Ux0qSgXXUBImTktpTu9
iUv+rSJ7Y6rMxgW/VO0VpcYHlZKjbiTQUg+0JRql8IWXK0kKSkMbfblIaf1NGrxZ
9UTVyCbtWom7o7jHSrd+5KJ4GJAx43MVsWEAXcMeOtwtkk5js396rc7uklNiWFxH
D+IHe2q5DRRwgyw+2ZsO+0rv1EZafpgOx1TYXsjYUB/Bv6xX6+Dh98diqgNSjqHT
fu8HG6EJBmJdaNexz7XheZPPXxr+pOT7oHqYidHDdo17StejaiA6TcFAIZw0MnmG
+tR/oLqOcOPccTHgVTFFNcdYMKZrybCeex+IlhCrZJK7H/MVGIkYX3lN9JDRXDbP
9lPFSI6mcz0lEbBER5veFFChHB1ICInilFUQMzAhFcNBpa+QqSX9MwBidwt7x9m+
vdItmR6bnDItrfZivXwX43Jer9rGRljX3sPP0BJWWvv/ZhB2dXEFZwzFCYlvPwCD
r1XbkG9r4th7DltRrDoLmOoRqGPjIfMyXlJsiBvWzThNDLe1mNT865vHjHu3mUxa
kRZC4fY7bLJZaBY3AlGzxe8sqPBgOLsMsCDnQmYB0npv19llakeTyPWjgHZCmadp
JYWADi0GrGpX6Z1wHc1NJ0KZnfTK1sIVVswz7/RBZ5JDVC94uXNTs7ob8u6pjZZr
PClntirXUViUjrK2ZjAP0FHYQpTD1iZLsJHilRCu+wLvL/MOWAwtDF86AGFW2n/y
XY4/7lxCa3T3dKZhVNRdv6JKYfFBgkEWfaLRhtapzMHyz8knwM3RkuMYqzref6+4
/qrPfTG1KsXfS9a0JZe87JAjvc3NAPSvVxkGK4naxrGg/ro4HvfLKRBlPQyYnYeO
9yOyGUMvBhI+LFLerIEqTvTtHcUi5X+maQ3AJ94PU2OWTtoYCmbW6SaNC/dPgJcm
Dp/JBfVVh5qmUzIKPQGFUBc7ZSx/kd3KJkfrADs6nI7A8Gx5S/EQ7b5OBIUoStsc
WdHnWqcAi/l3vLI39710E7IBZJBk5drw0pY+HEQDqM3J8Gdm3jffYI5merLRnTfd
MdOmHZDEzTW1sg0hKEU4Iu2R5sQf3J778syS+osgIM9H85Lv1zsbTjAcw36XkXRz
5MreACvjXm5ex27v+GWmUWEY1GGg2TH21SqruZ0DjhNQhNQIAcagRRkZuKd9k02y
JzyR1zaCDPgOCBKAAdXPKto0/GkP+xnuYVRWKfxecA3FKnckwlxZ0d8bw44q72p1
aSo5TUObB1CvZHNWtziwA6wMhfs/kmrUSCaAI8Gd0VbH+JcsRVMHxgZfBwbpmEm2
rKeUpt3J/YBWl05fS5yZ/AVzUoNKKkwqW+scrogp8XPmiksqcK+82yqxIkQbyZHx
6JxhXyG/IjFyeFKUToO1QzplznzwdbSzPfXpTZ+98gNg87mjhutP8+B8uveDJv3+
7bFl1ZshlAqBKLEMnqsv2EfvFRtHVCCiHlKhN+UlDmOVHWmbGSozaBA7U5j+9LB8
+tGIKZG5h1apuxKtg/vaf0KdImek85ouqPOC+kaJtXWgeH4p8XIo0woUxK+17hTY
dD65o+RVt0t1GVXVu6dp2p31rhwHXdlPs3voOsO/ZVZ3FTVzqG5UKtOEA/e19MtW
82lj0/baP1PzkCmfVgeJYM9AZs0xV0CDY4gUuKcyQejp8/UUJp817+uYVyhMgWRO
gv1zsBysoSOoyr113jse7SrxnSDloPOJA0VTYSN7M4sBqjshS9IoG09sYWrcHJ7Z
/HOUH3UBOBLHxIWpr6yHApMbajtU8iFeXb0nNMqvLSx6XA4A92shJUGnKyicCl64
QK32SVw81UZpoq3PRY69F2l54QDskbZPqGWywwIjUdI1HgqYLhhH3UweC9J/YPzz
b2R/4Nm7EX5U465Nd/Ot2Mi4e3xSjukvNVJpgPAo1gvqmxx0jvbhNodlBNsnbhZ+
T6yhZBSKoO336nyfurs9YpwbgmqRcsqMpTK1WcEgqYMkZJbpcpafSymbA7kw6VxH
JWZ4nkTlWFl+4sZFhXFaC2jQBBSBNbtnhl/RR0uyL8d4ie4f4kwQxFC6R1SnQHuM
Eck44EXdqhBJirBl3BWnOtmrHMDTxItPCbr4WlVfKRPQWYIpnBfR7xnteSpv29QR
5/hiqeM5IGsfiIRh3oVUagerC/f9USXlyB+9HzkPeD17OuwyhPB7cM93saAUamhh
J640+truDsMmUgRN8PM+sGNhEMUkgsfxN91XqDZ0vX0bpzo9ycdZaa+nw6pPIYX8
s0pPnw2Oke39RZGHi5oc0O0k75pzRr/6+ydd9ro+VLQpXDKIXFOStl9wFYTTc21L
TWjWAG5Wxe0EmoQ6n64TtWO56EzLAYy5bh6MUqu6kxp9IuWP0EiHSh8yPn1QhOOw
zmwC2i4tntEf9PCGSMHml1/T/+2ln+1XfPCSAHf0xIMtWKxyTtJ+eos8PcOnL1LF
UipZHxyAjMENQ/S5wb5qmPUP9rfpuga/k8ljZAzRBYct54eb0C/eO38039HOJdB/
nX4nxtvhzGBZPPB6ffvF0XHk/Z3lH/Z436Ns7VtyMhMEr8JlYJvRXJrMRiFQHl+v
XTFxX61tiZOLYWaephjC2iXAiSM4uW3EsLcW5c/NNt/3gnIGX46hzPkvbosQwSgk
0tQyFcwnJNWkdCX4ueQ7Zzx9TfpOk6S8iRS0JCrZK0t7i4InajVkOmEEdGGu+8ZX
iiW3lkILAkIlGNS/nOe95qlPXbJAyoxHY51+Qu9PkCOM+jzWUX6e8lfuOof0repK
/aZ30LU7O+1OMb4QJOJQskpAGFERdl0XjXAueOxK3dx857NGfFiyM/Q5HFcjowYK
1iK0dwmyE2DaQnRT+CBOwelWpNs4bT1KffAKs7TejlrnMLwjjQir/5ImKnmaTk31
iC2JqB9cWK02YOMBZYF7JK7lAqv6GN0z9/CEMWIVzzzkEpv0JwqjmxSOrIdidsij
PGJs35C2BHi0q8moWkL14fyJVgYmkC5so+TwmCTYW0vd59z4AR6+HGmrP7ZrSnJf
ZpyuCfAie+gcobzHzLC8F1SburJurTgWNxA7zMw5NEkOUf9mfvAsBS8aYxkuQbfu
k3Da5mS1nXxCxYF927Jf5aARcZXP7nOESUnvTn2gCk37gpPxCUDLZEMHr5x7iHGQ
rAtU1rLcrlcINdgJC7ADPWx2mk/vJQ/xW1Z8AawFgHINeFUtTfYogrwcPhvgbnPS
4CnW89mC0JZld4qvtuHKPxKpjG2K2Ti+dmfS+nSZfgDA+sUM9aukjlquwuKWnNY6
c4DJ/3d7AZnpvEkfFgr/Eq8AxfjHNXANRSrBNtRKP6+1Kyq8OBLCtxSi/SXO0VyR
070rsMtz+70yx1iCtSa0UTZidVYTkyWdUq+SKiyOO1MJNJAupMtVdYcUAIgUM6dj
K1QwuWBjT6mZB+a72X8nS5/YMyKXbHrIWf31UowdK10Jr+qttqPpksaNRu40hFX8
hxfoRegVFkkbu1ceiMXtNUIx+Grc+uLUxSSQzWrDSHHhINQgikFObDn0ZxBlR30f
MXswPsRl5XyhphWV9+Q/FYZ5B/6lEPXjzaGnFLHZeZVhxVyz+W9yu4cr1xNatUtN
vzO8hz1vVJUFcPEQeJQMlfwH4z0L16brYXsfrVW3TRKfxju1pHEXWX37Oq5dyxYk
fUcNDxRN2sa1xERyr/iMKOITKpYA9WjgEFxuzX74SMidy5TeijKxCI+JfFZvFmJ2
d004EVLO0rrI+LNfqvVxzLK9xX5EA3mOGHfLsl0Df4W4WqvKPL+Nn+wI5bIKTXZ1
7lYQq/wAs63/x104Rw/h3IIKfUmaUKYNDZx6NTycBSrVgXb8p/C4J2E68MzEUkg7
LL2IGUHYlBecMfZVOgg8prMUDUbOepQeLaYacQIgnf0IpVDqBZ2vjJoCcITfMNZs
plMznSzqIXmqt60cAzwo0kQIQu3pQAeSLCLRQdqIsWk4+TKwj1THIZrXezr3NiP0
pRjSlLOpOhMTXvthEBU4yH6KQPpF6WULCl2bJorrIWaroGG+dUKbl+onrAQY8cbf
noKTpXheTtTI0j4ycwPT3ovYEHZ2GtMw0At/kiHJdd+8L3D/J2GmHCTp9KHfHdYb
Eb+BtaLwLSISCmOj7zYVXxMF5AfDWggfKP19Peyw/v8BDEq7YA8+rYATUCgEDOfD
ammnUzxSNxjtmf6nlkNY7GUKJVSVyWMqDB/16KDC1CMf6v6yOFoeA4zC1wl3BLNq
iflVWqtfT26RvmfqDisL20CD9vTT6CaAxnYppif0cnLutvAZAMV+ZpLCZovpF8O4
wjLXatjey7PitSZOkuXVkLCZkB0jcTLIVY6wa+9k+nJ5hwfrJHYA+8R339C/AaMj
tXYCvJN+TjyVmr7RqGdDT8vaK1m8vJRLJw9rgdhs304xV+cuCokzt6sWBFtvPoRg
au/QhlSUKuOi9p5iz/1igQCxgMAdVTAksvr4D+W23UfkpqDowDAG3HFPlztxPATv
fxwbU3m//jbx0amsrmWISQ3aBV7N8LLeF7p7C5P/6cbovOZr4QJZWRj4xxi5dnQ3
PkDDxm8uySOnHlvrhDo0krAd4A3P+go2pR6A3p6a7j56MYrTrBElwOcOMn1kCC0d
oBBf+hI33xLdZLV12K51q/lJjwW5EtfM6+YQ76dADEM/aRG6+892rlCbqM9sgjL7
RWk+lQsR4Lgjmu/fhiPCPn5kNbR019Gm3WuDr5ysZC3FJE2IPDh6aBdjqcvfQVSU
zDuHEkNsEkeJkowvqiNUhOBcKUupNzviZ5Ve2vuxSRnHRD3NXjvG+uy8jis8zPip
i0Xj8BXoegKMzImsECOmy6hAtRMQ6UlMgZV4xT8mSp7BjxmoJG1OJ2nuXifHH3TW
n99FpfHJvfHMk60A65FJJF+UPzNJhPd3h6VoDxwobDcMHXNzEtMIlh68jiKuUq8x
LRZLswnHVL6MogspBF8ya5kpQFu8Q31Nrb17imQXwukIka2ggxnigQMS2sQq2Jeu
/Qq5siC2RHbo5dYID9DrCo7By6CLEwFGeq3E7+iqif5/XH8mUPQg1smB9cb/1Pos
7kNuatMgxPvtkERnqr14MEoN+irs0Gik3EBv/uRRmRw6YfdOwrt4inMGnYs6MktS
7+fK+pFtBkliG8jxceW+VRgTnZ6I0/H381AcdrsRndLXknlIFfsCK6E0qmGru+hP
g1omhT8BeziVXLSA3xI7LgltYECpNSkFK0Q8wEMA8PScELwcUyhWPczyZ7lJHcRW
LkzuygBkznvELXgUhkoKKRzPI9DbWeta5Lb3pwXmCmGeTuJC7DIe4Ui1CK2oPjPt
qXNpdyZeX5+3Lva8Yx3ieCC0rBsqEpTd+8ZWdIiZGo1XJjxN5E1gxr/hKsM07aI7
rNouFTfpFylL2NBQzh+GmU+uk4Q4weKBwoj46Fo9uPKwj6Ia2jJ+C/sp5MhGZydY
Mk5hmfgX4LhJbSv/53BWMNeZ4MYqL4ELuTzKQdIYuLBs7DbLUsq5A3k37lsGZNDD
MiKY5vNJsWrdk1ZrKRaSbqMXJP4B70qyzhFDQvLKuZOYhcNul0jE0017o6q5/jwc
EcZUjuz7a10H/EYpO8B6lnCWMr1Up41atw2MOtUeePvgtGcuv9Vckf70pw2p0njN
GFEtq3Ck/ftime7LiZo1vOINCkSUSqecU60PnTF7wSNo27x25RSnCwlRyFasBqJn
5d7qBA5GALG04E/hS6n4wu3v7DtZivn7b9udYmUOZaWIXk1Sy5I5bpe4CZgMLK96
j2XfxJKy0RXqkB4Cl6XHdwfOzuFFxk7D6uKYlL2gVE3gxH53RjjwQ2HyicEeXmbM
n+9X0xPmbDDW7gSsUbnQfAwL+8O/J5jTBwQhLmRoBiaELWvZMdxEaaM8osymJ0Rk
vF+9ENfEjO62QFwR/ro1NCiwhDN8PxAQHecQD623fyirUdtsa/Y4KQAkiH6tR+3Z
8Y6xBnEQSfmtbQkCh7EfOZZZfMK383icMPWeOmKBFyEM2QJ9Nd4qmL9gUxnaLgQA
WVfnfLUZabg1RdwF54iOyt69IESvCEe2tk1M3dGzyX4P5UqxxeVrhIW75hGWzYtl
SFs/PmqIFjzroXUPW3a5yNzZnLB2NRy6TOL9cRBJ+NMx4Qi+CV2eaywQD2mOzNuz
Wgc6F/eX7vc+awdRwefuW7szkFNEwPBnhBYiN+1A8aEPSmhgMdGhsaKjhEYyupYq
33HrTLD+9C3Lhao3b8povti9BkfSwFqLqtylK46wHnpLaRqT8t965XaQ3DL+H6Cx
jhjPKroEppKCw9aGVWFMvFtjnwp09wqnfQjgzGAsKdtbZcMihrV9WQ2R9iIb0nFE
NkEXC00ZeYLL2Y0RVefRZ320YOpJz0sAIV6asKjTzV3uLKd/XUkBqNcKGp5U8XIz
wZma4UrcSMjEspYE1bKzJSwv4KYkbQ1cTv/sQaK/oJWdROp0dUtSw1DQJ2aGLmLN
3SMIpBBTGTfIrfVXXYVq96/VH3KUnzOkGlSoYRMlyUru9dJ53dSBowFxoO46Bvxo
pw62mO+cOSR3kHok0nSO6FHzl0lAk6z2GYaApAzHh4aQ7T1lghVTG5XeyHatsXId
k8J54xyoM1Q2O4UVAcrBgHztk7q0JYZM4uRG2DogR0OWUQ+p++mUo6GynNuWd3vS
AbImR5z8o3NVRSLFxNKTBowhLwitbdi2kWqgjfFm62fcqvtoe2FzsAcwid5o5ND+
5HvCi6/8K15+Ryfjc5JYCtnXilVfRw7DLa4lnVno9i1lPsGiaTpnGOBfrWiacxuc
QijuoPgMpCyBq0tgFQ97nM7hiKXAHJiLjawL+Bhwid99A7W11fk6SElT2iMFyAEA
aXlYmFEOzNpInn85jFiHZX80S7+RzG1K2gTeAjuTE6lH2g8U5UGOOm3YX1XgWUkR
zJcwueJROtjNn1Bc22jjWSpUO7EAyZ1MtQJPTHYRPnfTC4DZ++PKQip+Iv+aEBfE
mBvIfbqyCAkOCy6GlmM8Tvq2ah/uif0B/nQKbgOSKbd4VVC7GImcXtLWpb7xpmWs
Yv5dVzn4SepllCUEOc807geDackuHk7cBinNRCkhO0v0pudtE0btOSrHwDtKV0R9
Ylk24toV9AbnJJ6uZlqQy6Vfcx1bQxNeaYwOAG9MoBZVxawoQG/no/VQYb+2Y227
9go5CMkqwkPGipxubDpHPVTEO5KaWPBx1HgCMJJjxM01G8AnFvDvFA4cXWchs1HH
ugKZu6TSSX7xTwi+BUw6WU3BxGzmdB1AWVdicSJJTIKpfAQiYVwnnF01rEo+AjzM
sP1zOEVylfy95mpvvvlsuc7+Cz229YkXzx/DoQItZsiX25cSvmjz6IIT9B1njUE2
pj84tdC8Hio4/Z5uxjHCt8F9dbx2z0kBdFTssHvil2nmEqvGnVSNMbT0ptk0RxsO
U0lb5ZKgC0yAavsl3Ur3L+us1fzyDQyo1rMlHdQhKqUaMuk8fCvSty49aw+y+GcR
j+LT2wBiP+hlzCeTOali5bL9fql2ly+VWYWLVRoZ8kwO+icbqrRpcEDV0NiY+aVH
wgFEPAPfGFbuOHI5bcFkeKhJNf1i0T9uk/P61jpR9S0983PToLhmnAKRM3wvf3mG
LsPY8mxHEkM39RDE+CvCI1EiO9NcJjUs+ogV29PPFxF/W0z1H39x0YYsVdB2iqGr
k+CVMBWdfl6S2YRFbcQ/hqD9LVZqozhrI/sE+Wvr5RK/q080uyZ1sjSZQEDRY8hH
5JmkWFr3JlM03llTztQkmt1N4D1rKlWvWy1/EPVQgWfXVABi7DAmy/GXFI5IDRLU
nYBcm2sFvKyWlXPfRz8nDaAWQOq9HN6nAUoBRsL8WZ4b9UQePiKIfZoSA8vBD3zH
Ql3deeoHbhmCAhKhLeFbTShiSNiHsuPa9+TQildAgd3PHs5yRrzijQyyt4vFUm92
C/khKf3xqZbufPHOWtSGldvz738fDEHdue8XILB2lDMk5BFL1SNLQGFNU1Jmwyuw
X9QTyE6Vd2JQ2Np19ybSTRikeMVXwToedQ4g+STvwdlhWzDDdqwdgOP5cT3W/A+q
8qzsIV8y3IJUf5bN9zKwihNI3WojsOH88PUHbUgc8PNnZfxhPRVMOO0QZBE8vbjQ
WW2u/mcSprZalIaXF+GGRHFMGM6e3u4rHoe6AsuDE/+lNFr0uuxHs5y0x/zA/isY
XUR/ge0EOYvc5Pwzn/Io/e5yvMi1pYqUuwVlKLa3Su+g+IzifrYvgYBVygRVNtEv
GVAY7UukWhy6cL1k/ZIRKdUInFf+8k2PiwXGQNDQoruU0e6Ln0ly2d7Dc34fKzy5
dc1iXDnDvfM5VmU+yHw+lkE7O3E+mxWk0QQ7/iSHiWcLjyuysiTI1VrZMs0LAhor
y7s1/H7L5sfaKPUqMUa5iHDhEyKJrBzTxdw+TC4ZoYO3jow4dc/jorlucTJ74MFw
iOqIJ1ohsW6JOFcCv5ixClhtrmdIygpDyhzN2ZEPL1KgsP0z3vhXi9ay7iN9g4U1
vW58Ue2qe/rmbKfti5P+vK8XOTHYx8Aki/NOWXL4DLCSypCLf+hatF3YCxMtkdqq
iiqNShEHPiMgvNyXqhM+Pb745eVB1ovglkKrUe2Wt8cetNRy0N3lR9nkysCVxdGC
0LKJNrI2O7aXQbEAXqy/jWeuFUddSbtaX+wKay6QalFv2J4jb6Git6spUm8/j7Sv
EgUYasW1B8HClmXbfv53G3rCXJgSncHHjXeyxF6lD+P3YX3FmuTF+zhpG5Eq9onQ
z/ZlUJsWD8X7TAo0cLA+ejG0FNKeuMJYgEcbA48yWyH+Ba26PwvdTGXrCMgaR+Dr
U4Pls1ckIZ6cZD8ckLj41BCoSvWswET2RoA3LqmseRbMGsxDGwg7xbczc1nXkCsH
pNB7vgyxkRuopQ9DXEyzMcHQOP6f9qbfT6gMH9tX5exgUFbXrHS2xfTF5+m9s6To
Vi40T/mivvWR9yEUpvjBeYqfE7cuxvM1C3EnBV1mhvJHvAnIRI5dTGZaTt3rxJsq
KpPdvBpboMghDkef10iUcAB/EyaAopUUoghfMo/oWnDNEuq/KwnAeISs1WsrmxKp
eu46FeStavBxiPWyG+7fCuob5Keb4f2XWxm+OOBGOdDmlT2giZRuEgJDd3sGQEww
0c9/y3paeszAer0BMZfU/0td65YUaso2bKjzEs2kZZ93jAX8rgMYmuQhMQop9XXA
grcMv2tpwfr7PdMMy+cI9zJlI2ej6Vrr2ZfX78FbsOnMCbHY7Y+7OE9aF0BDz7/g
t0EtwUIbGQVMs1Re/b2xFiIebxKqnSsg1mCuU+u3bHGiuKX/4PgQpAe20CC2Fy5t
TLFxG9FKKOlJxx0llRu/h+f0l6e1UR+Lqx4iA94U5xqZYFHQdAsEZgsxmzxYzvpe
f8jTp01LalAKqWYSzAcx343ui6rwG/6LeO2vxi6a8GdkDdUCIwvZUJKklKEw7Fch
A9WJyFRY5nWiMfBm0Lok/D5SziXhfYSGKfm63In1jDmSeZ18IIho5ZnTegrdkzjc
aKks76E4FJcE+2AnuFzeV8POOZqdwssV8pe9DWRN8wCloEDZmjU4iH/nSL+HsBdX
/xm+k8E62WyZ2wxv/hgRt8xu7Ap369/adL2DuqJjxaOrOQG64N1o7BvXOWhs9oF4
m65YI6lCL8oV+KFqqsvWauOfmmSrlik6m9LRvyPTE4NEDCdTINdzMvTYGTkfCYsy
+vonmijR+ARF1aiuGCKAF79aZdjmSUzTtLn5lV89H64E04dVAj25at6zHsaRrf5i
0nq7Lw5FjN6+8dX96aTGtpPQEitIEieEB9CvPJ5G/IOz2uhZ7jRWWaCPjx8IQ/dy
2yftdeskxm2qM3n7kPUA+LOZ0lqAPi9Zm4uNZvXvq4C0XjmTuWDqrHgbA5a+kN02
s/toN8IcMsSP4mKCvLHjHTHtNuIVEeRZ+j67SovLCkqfNXpAI1HeHd/LSgH60i/O
Ws5lqq678AMUZaMvMWGH40rx0a/w5HbruZFWS7UN7mhNoiCoozviHB0xpKPy78+0
n15aKZctTYMhOS8JVCW0V+vnHBe8P5JOliBrUo2DKpl+UN0lWWRpb7eTwal9Vws4
7HXbMRLTpiCYH7Z2rFRqRJxeX1zuECvoVGFpHae+i/Cmonla0RQZoWq2IY5QY/bc
66cbCaMU88vYUszAMNsGef85R4lwUlFqs41FZIDK9IgUAbJmrHN+GEUoH+RDCA96
Gj4YCz8Wv24E+cAxFJlfVcJ6sFJNYAlfW6v7AHnBrwgEYNSpdd5n0lFuty9jYUSw
dqLDnJpxbFeMkFIrukPAVdo+Us0GpoGmQopd3kF1sXYjfUXdVPRg5X225xxiUpqM
jkjYd4g1KWwaOSAE8xVy2KIEunPkO6nmCOtJzRhc8miTaejAvUudBew3IT0B5dwZ
YDpvE/8kqr7d7cyWdhyPMVYcM5npWvVsmf645LVbMiUcr9jN1kwqDQA/yHMY7T2h
cuaj9jsY8ddv9XKNhgBIf99UzFxJJdat90zV6g24B1Tzx1O639eS28Q2Wv8LF6bC
BM5lQHhQ4/QbcK8rDaKrBsriaETEA4hlJQL/Nn5/roJMu4Hb7JcoshJLoJFamtfX
siyumibZozkGp6SWBxZYzUxG45y3bK5cLY9umQ1ZmWkR7HcF8FatOkjjoENa6v/b
ldKV4gejLr8J/ZVs/2Q3fx4nkam+y849t9VtQw//2Zwhyi7lcLSsEdSgTCcBC8mA
LMiTaYAUEAYSZdoWtQr4n3eFVeXQ5RhUOQG/t+jfU+iCw+DWZtlQcTuDNVVlqxQF
d58k/spkBUNFPgQAHg6LL7bOVlqjZbVlKiY7L0gJVRWpfUUu6k7Lwz/c82OdHM60
5Q822af47YV2LYfboMyVVxvBaF8h98MoDmR6aeA582IALD0vFmKBHI+Pa76EKBaP
7+yIlbz4WGOcAzWkq9YNoDERVcvbT62Y4eR/fWq5PT/ySf3pZ6GGtlkafLUKNN4J
YBuafSrHo1N/PinVCKe35l1bzCMu6b7uMA+1IR9z5g9ekpap9SNF5wbAPkhe9eBe
NsSsTg2ObO4WMty1rwunm2uV/t5A6dZs700WV19joIuMGA3Q9qYR0PK/qI0Wd1uv
efIuSwLVlLouUajP9jGCaGfelpHe7QcePxTq0dvkENy1Gla3WSQwF4kd3ZOc6a/t
0IAgYevy9Dkrf8J/MkMwxalk5rKxM/UDvH3YPrE6Z0GrMZ3jLegAFwSI4PdDvJUQ
0kk4uz4chzbgR5KMyNyhSuTd+btapGciUAfUoW9ozrITKdR/ucjusMBhv9s9kXPa
0Jrx2ggBeiyG6ionw+jIuwA+/eMPIaWMDQA9uVDVeHtV8lV2Ycv/+W0s5MDviIQn
czFv9c0jHL9i2mffJ5NP+A2mRXPUnFlDzCg577VXnh+8z8d8Or926k3ZqKrLd4Ix
R+UTh+qIzVsKRnJfj2hnz7yctoSo1N6IuzKwHHFROLCgbqLwcGhYSXp+Z2oJfhJ8
8qvt+UKmetKASk0FJwPBFcAJy6EsGs1Ybg4eFB2EqD8aKaFabiKh8qNRZPPgo4Ka
oSrhhLhENcXFq8DrafVyVjoZctP7q2DJTyMpkgTZMI43CHQpOwAb3zy21HPjQoWj
WzmsW4qYTQVUAJdhv7iTvqv+5xoxvmjpf/POtsybeUFQpMMEwPtnJ/DlauWEAVkr
/ljyucFAgywMtwaY/D9OIXlxlYM8P9Yo/YZ3mDN11j6BY/8/3AxQY8lVuhjxR55M
e2WKBi5bQG0spBwwPJ4bqIbZJFRq+N5By9ecSQj6EicgWX4n5veq/nGXs9ZEHAdk
HrDJhUHeabQkcr2jtUMK8PKQeOO+utX2Sn6SfbbE71CWsddvd4hG5pQxojoL/RZE
+NJ58A+DLq+21fhL/a7ZsgZyRLEk2ckh34ivyoClUBWDnrHMEw2VJL9b4wXATX2H
H6Kml1oS38ETQbcW2bXmHyVrss7APj+9POwt/V3l1Jz7WwPrrSVr5IulNkQ4+UC7
tJsuGeHv15WNBdERVOoeaSZB/JQx1tfiNRQGJRQxfoen6Ml3UD6eLWvDJddKcfrE
wzIVcX2WS65BE0zf38ZTMWXAay+h1XFXkuxfRJoGh72lx2DohMsUWYJab4r9mJUj
6vZd+qm+YyDLK5PpW1IQlIpNDrbop+u7Pd6CyHH+K3NZNNWqMRjFnEHxvFIQz7Vy
HsBlC9zijCTG33B7rT2vHJs31DkNx3aDb4wYMgeT2zlQmB1gefUEMnWPgEiUO5vS
wdKp9dTyEjtERjlaOZkJ3qPDr40oNbG5/2Q/5oEnk3CPEbzCMmiaGGNcG16yCQsf
KHUu7OKfOdQ5HErmvPdKVIGlRG2JHSgv22l3Mp8tNyYTR817h3+f1ZgnzEeq9qSd
hAR5hWfd8/oHvXac6tv63+8dFdm/E37rZj2fRaBb1rNJhsTbixjFvqpS4cF3RN8w
kYV0lJkNrckznwFTz8fNyJIisbK4xKkmC6xn85oXGSdb1P6j6bx3dIJtXvkt/79s
Pz3eiVGhNs4LR08PFaOZQPWJ2vPz927Zuzpf5D1o9hC+2IKPtigpqmsLUAtLU5qN
bElsN2W8tlkNE3Fyvz8v1UZoJ8M7xAQaYi1dBhfJ/p0ljNw9//7DehSlZWc8ZkY0
Rq8u2gStI4P3x9krEqlG9mXun7wnXfgGF0xKu2VDZ/jAU1cxJ9Xxg2y/uGXzAgjO
uStZJcOMWv0wlPauyjIeLrd6zr5eHSal7VIXagQLQfXGjYv/USA/mjKur0kF+1xb
taXrDYO6Sen3+E3iAd94T+HoRpFDXhFeYzBgC7htWmj2N976cJJLqd44cjemR+D+
1IU8m30NhxMVon/LwN2vbQvg123JztTai8pDlysUomcZn3NsVrTSbbajbMfOwGwP
EknT6iNNBMZppZbgKmuDuu4bslYxJUcL43Odqlv9kat7davFx8ddAdyHsIKCoPGD
EuV8UkEF47EOLBF1AnrlHNANXwUnMdZrfWt17euv6UEhud0BL1kCEjbjwtZQbITL
inUzir1lnbv+DDvFHynTzH20ZPEq7NsA/xgXFYxdhybb3g53RhU51vbzZQAiq9uI
ZGdrBFIHUclBaEPTxQZsJySEMNZCK2XSd6y7CTckG86OWr5m0cm8WVD0H1jEaxS9
3eV2mX9qu/itnrICjOR7wvmaLhSm1Dgs+vRsAmYTQ/tKo/O2pw6MWli0sR6JIMa/
/O2gbn7wW+lbGzGfAIoelZ4BgHDLfmTu4sqhJg91KUQ5M1OsgT5V8tF6Z+oNz98Z
odsmNFF6d1XFkn3oelKKjVVUxrWxRXFZ8XBLaPBWypDqLYrnUfbB0crKxPNOWnQ5
nkOxUITcA4+YuMiiLC5nXW0bF81mXQuXY73PQMEVBeB1JiTp7lk/7P6OtuSnmXBv
5Ls492JRTf5yIz35GCJSO4eIQeP6tXbNIRI+7Pnl0jQ6FxzG1fEo/gcGhylBMf5D
Xh2oxtfhk61QsMl94OcQtcqDGUw9Ekal/OPl39fCRVH2YSeygYZgcyWBAB3INYSj
unwEK+RAoSgXs+oOB1MfG9fsCaMPKfqEpWb/+a5ywDIYrJkd9qoZK0T/AWzs/Jzh
movNXUUsGjKyYCXu7ADsccFG6+xJhy1k9kMIASvdn5pL5SQtQ8BqsQ+9CsapK+KA
3Q1qN08FeHmGQZ627lf/2xc+gZZynTI0AUD+on5Aw4u6ZqPU+gogTeASRP8qdbIX
H1ncSV5yS+eVrIdhRt+lvun2YBYM21072PTCt8P5K+NN0pDII7WGsadMbJ3LyUvK
zzAIicKcyIV2A6gAHaKblODNYD5DIejB4jkFS9Cv2eY1qcDxHHA/prQ+krVb6Jpp
wSuGKUtcZKVv3GyPRsLnenF7UW7LBMH432bnFWkjmVe3+fyp1jqyyc5RSVrG4RGu
+NPawhtMkWd6uBSLsomWnWWHWlRCkJAyv5Wp9pphRy4NTeKU/O2Gmf43SabHfisn
BDeh71bgZPSw5bHYeKf0di31cU4w97uM47MK3oNi03T1c4mdelOvVaGgvagW8mrn
cmFr78EDc3B/I7n7XrHiDfdzT2nBMJ8iWlLOlyrHEze0yoOb5nyg2raVeeE7grJG
f7j/kcAogntUPzNvyPvyhZbzwNSvB8pIKNAQZyqA9efmIWOA8kC4HCUjALL2dZcE
OrCpJgy1t1qQuHOCqWpHImKtAI5/v2NE+aeroSFmyOGJ4gsAMnVXo3cq2EMSJaxz
CVwPRU2fcXqh/AHLG5YWl9b/mkzjSZwNXwFT9M1MN7Fw+wO3WUIbT8JBV9iAQmcu
Zp+c71W410Z5uphoKMGHygpR+nTqxnzniFlL34pDMVGeTaKe2g1E674cpXvfl0nd
EEjGTN/9ftYXo7rSq+ScE1kOxVRpXV33/MZAmgQYN7Mf2XJr46EZuocbEgqSEfLf
tBoN+B3HkETav6zNqwSAekLWfQxTdOy30499YYP1yJy6U6jWcDRSycdZCUB7nrgy
tf2hB2RvUhs3cHCbvkXxKe/jYjJ1C8zv+pRNyIoiGpaVb+fBV4TePHTqNnVQBHRL
35DwXDlOSbSiu14cHKrgw8mvAKdjXSqqfmdtqI+XjjE3bdaj6656GwLDhbPrjDAd
UMR13Jj3tmXex8heZkwzRO3s6sKhNevy2qQMUJbSzbFnzPAPKYLtDCHaL075rPQN
lbv4ECaOK4ZttRvY1Qz8rDiI74W+USdLRbILu+rzbHjuO3TwXYALoS6pqsj/bgJj
CHXd2nzqPG4KINJdzDB1S+z8ELrEmUvk0ovabYwbZh6Qp7ZWQTBChUvdn0+qIevx
XiwcHF9crcvwLK6oV6RpqUzwTw6/zJZNim4QI5KsrsUyf+tFpnK58eE7RfrMqnn+
xkCQAMjjwYIR8zNXdXa1X6LJTw2/mf/TQM1GaIwgslSVDMuUZlvgmeVy4Y0RoAbi
8GaUEaMlFRnnVHsgMZ3aWjrQQRchHFtDFyaS3GksmXNRH06aYwIqLBEzJ17JRcDp
iY6QeP4wI8Ewizx9Y9vLt+Nus6Yq8fP7b77VPzJg0XBed6TKxbtKaeQm9tYWMukD
T4JEDspNy1gCqiDexDvyXndwdY1trf+ajmRaIcX4bSsMbYy9T7n33w6h1Zyj+9o9
t6b5V0KwPy4V3ZXJ7pF9KLB5bsbo3gZaV5fqxypP//T5+S7Cr4JiaJHDTmu8atSi
clNSQEODaNNwx9W8ibPzkGfD/5xWpYp17ugHETsRJczGy7fcdWcxj5Z7tn8Za0ml
/jtcZf2Sr3USzra5f8g5iz+h4YDKCnScuoREIpfII3QdzduJd1M7UNAFUozawiKM
HNw2fSTtbBMWJ4EtKcQOiyn1CFOTHnqZ+ISyD1wvjMPJobTFv0kHx/pAEbjV0upY
eDvOzcArC1A0xLHsIds9EzhenuoloIgEyPhrENFMhbnRWw1NNenD+hOYJ7X/aTA0
RXYLYOluEsM4WWimYRzV8FjQviu/GSK7uWjY0oCGTUKH2J53WIsiJqLfbrfbK6cf
nQVpf5oU9UJN7wVxX3VxLSaPl6NGq3quZjnJlMcFgS/cYldUU6v7CuUAhdbA1+vc
ZavVeG/YBxvyw5Gha3c/FI3/izjBXjbI+90S4v5CA81evBdYgg+Ha72ughBxIRTq
xkP0HR8wNo4XCtB0UD4XHNKt+8M+aaZSgJB2pmHuscqMpLyqbWpd/RoohdCubLHy
1OONk+aTADYaqEB+jQc3pX3qvjaf2iSWIH19QCPMUiy9qc7+cZmc4EI0YPRhMHce
YJhDQIcbSe1PeVYg56BC4o/a0xszOPlltJXki5wOvjydNk9MCqXpMsEfjsMnSvYd
6/aRbvQfUQZeNgp+yuZ2C2KqktHs8X30G0MGw5+cxT/M9LlbqPt6aNRYwozc1EPX
p+eIZSAlDiSpTM7bWm+tiyItXd67TKCzNnU2sjTYJpnGdyuCDLP3l+zqcvLEa5ZJ
`protect END_PROTECTED
