`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohb/5sf8lCS2YsFLCweXjNRXa0v/zpBeZv8yR3H5Xl4FYvr1AXu+3ZfGTus9FX83
yEC/V+kSfKmd4H6sNiA9RrUZ+qe5A7RPWrPzVwu12g16K6CSyK7qrKqjVaSKv+bL
5a3eSfuZQXhNX6gWPIrCpTR6SHtw+9ACuwAbAmOh+UyHpeOuc1w6SaQ6uaOZwoYm
TcqYNEt+PSoMEm/7Fud6QbV3Nv6KYHbpRdAuSQ1UDPu40oJG2doN4eSx9HacEBFj
qGtAGkshsxDy66W0HOUwfsqljoUGfnik7CYvy+4ct0iN3m7xkVij4nm5TwidoSpa
UNouEE4esiU/3ahGaRqX0uUjcnEdqZ9UIKXnKwsgm7clvE9EmWQnvE0zNJZW0ZHh
`protect END_PROTECTED
