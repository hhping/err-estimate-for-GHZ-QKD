`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WuIls1iVBro/ArweoCEhhoroC5tYlI2VgoB6FOC4XKbV3VY+fI93E+TsX4WaOABj
JbUwRCRmaRj+OX7EJuw3fgOvGdrL8I7x/CBi26cT/UUSx9SGs+I/SdhB4hG40iTp
MxjkN26qAcony53nkdD0xBxDv2y08I2OSE/g7IwUap8HhslGplf/w6Xo/SIFDaRE
8ShreOgYgu4fqfzECB6zq51qXpb/Vd/NHH9yuBA3w8AMeSipt/bnEqd54KLELeHd
n/5aVEjtV+7tgHK1OiCOmmNEWHdX9ZqOUFJmB4AkY83fpmjEnGwKvlx4Qy0t3F2s
g6GlMBKaAxwYPjU7sUUUCKHh4CUwI489CmdRTFJbQSyDNbYWO60hVx8m8m3DrFcD
X4GSBAjCq+UKEwuCBah7J+7bTPX9u0sEYJw+VKztn12mBP+T0hzQ0Shk/J99WaLM
9VZlTSXxenPEhy/VJnNyLR4My+rXGMutjVqI4d0LACO4eZCShXRp4K25y3XaI1yf
25rXkHrqlBflX19Wqqbk7Pr4HmQbpjqSulgNBFPjzOR3Q8ksmXpZc2ae43hcIrq6
aWVlBED9eAwUmlJDEI1Pk6lYkolmIJzwJkqiE9O0BgPW7EwYgsj7fEvI/0vgzpgP
X4zHwNPeO5smovuYPdkr5nBzU258wS4YG8D0AFIpxYXI40C6K4YJc6S0ldQXO9aq
CjPwzIzYxxFqYdmf24pcKalKxErfcKnia1vdddObWSY7i7+9b4rmQTFcX9GtjmbD
R4T3CPdy7MNnimY5quMyPI74HkxqChpfHTh166PQ1Q5cSaZk3yPgNYvI/sGb6emq
8syrsvOKZ7VDhF9QZm2x60DkY8DHIdOMcvfoaIoKo6V0kZstZmD1IXtyRJaiQmYN
jiZi7jnp+bGCeBWE2ljCnbvPl+SaSX3dSwJ6III3wdKBq5UycmJ9E1Kb5YLUVyuD
DzB10/Umqsvx/mOYptsYB2JtPVtF1ZsnqpvPsvyTgSMH8jYAbEn8Kg86CtWcvj96
gsdHtIntDo79fGNPcJJ9iKL75v5iJWDU3ZVxXP9EMVQlXgcIsq3of05iPGvDybiY
mp65G2moC85d6KJFteV6XOBjlpPNTM8H8SMkZwFIrJR0IE6EJ7eQ1bjQR6gnEVOG
d7HerZLr3u6SDH5zAPcbZFdkf+gutkGZZ4XHrL6GKgtzEOw/syUkkXMjZhotNmBy
HKFy7Uv9Gknht3uXfnKMd25b5+6qTxFu/qORzZ7rrE4z/wUWPnBP3MJ2/I2idtVI
kY3J1mQhYTtmjoFoCutdVNBwphwGrNvgPhCk6TxJ/B3y/7dT7Y1G2eD7f1qAUWbV
1QRN7J/Jk8ZVq63QrykDjJJ5yX1LVi8a52hU2l6FpwxsJyZLu2Gxvd2HIKgA42Bi
ZyRFYi/a5tf25mBlmfWv5MU8lslOEkZY4m1fE1uXJ7PvRaPNA6g3CI9wm96tOfJM
obYmKBeUCVxf4jbLpnrchoWJsdKvHZCK0pQ7XX2FdwT+SrOvnQ7O1nSVdTpsJXPG
HgU/WM7VNv+SPANwEKhDzj0STKbudcMOeTKmiZiX37eBYl2WGsxOUm2k8434oHhZ
uduplBH0cb457GY5LjR1YHt3ddbXkzo1dEiVdIo3/7CduGLI0JcyEz3+ZSdRKILw
`protect END_PROTECTED
