`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
loPpD3ExHDkch1gZxszIkIreUPhU1LsNq0GKn6qBV/uWvdJzxKyPOzfJLV9pHPe3
zsIfbtNc2SOkRnh3eBrc2+bEV7E+/baVdqF0mQnLqBl17uARFckL2rdG5l8mIwYw
Uh5tlcqC/xEZWhu7AfSFYGTwIL9pM/Js/LIKJdGKfWnMYjhWbk094kziNk8g2Zw8
3tA+7nTepD56vcdAeJaoMYLFlm4cJnx5eWjRL+mPtKM1Ygyk4pHOJ4IopE/DnhQs
w5JKC6LRfSfuLBSzEteVaLC+t/j3T+mMaRdbfMFJ7xtUnq2oRF/N/vg+2sguFF+3
0a5JVc3IYKDKTCcVyxQg+d9r1TTkMXapnGcY15xKDoqANDS2Q2AnwJfLK9A+DUb9
SjhxBxiq98Uyd9xA6sH9bsuDagFeVPYKZF8zN7pKFnikQLotcoORUM9GwqSaIaVR
ner8JR3UfmkAePnTpHf5MR2c9bvXFnfpLS4TQBchhuZP32kndUWLfre+Y5OCdpCe
LOC4xRZKxmXyeoIxowl78K4Can8NrR1FlXrzmUTZCW2D3iJgXVPLkV+kx4OfjN7C
B88OkwJZBbOYi0hNRHksPWVNVJ55hylVvtwol2jz8fe3ipV53L/C9HxxJmS9qPkM
0FkpDQyzJoPnKe2HYPuGPnHt9Y8N/sI7bthK4em6uo1qC6sWuPs5INIS7OlOxX2W
3Y6AnbZzbmT39075qpwifdruUCLtTGUI1n939ueIcWvYNkxBSMU2S+uS/6/8Nq6g
OoIqN+FUBwBuQ+GBijy8cRsEQUuFPJvHSuFCDPPQJBn1qj+72oQD5WnJxAvm3YSK
HbJifOi2XZZZZq7KpQu+3hRChjyftYSoXOIo2Z5d7PFqMCgIFvppN1TE+ecwjn9+
siapfB6mgkyqWjxaXWb8JlB8WTIx31UXEbdtnvF7ec8=
`protect END_PROTECTED
