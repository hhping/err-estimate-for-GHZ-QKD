`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C0AA7emkD6MhV2eOxErKeBYuEEZjVTHmhzHtVCfVbT5TAYoGGDBQNPYBQ35/TAUc
s3Gsh2iu45qrzKKR8HEUDs6tn0SJ7Ch1QjzIitFgBOtYoTKBdCAZA5qt6adgPZWs
68mi0uBMvX1I2k2LlPfM6XTCWOLodqokFsN/NZFNaQHKF4JaUwQOUo7FfX+H6WXj
fFVJb0K/rf1RZqEw2eEm4IJVG1aEB9hwptRHjZH6cMlSnOrqHKYJjNqk62LaUp9Q
nycsOFHR3nuRw8PllHMMrQ+hHem984Vx/tH6Zve+bSOacf7nCl0PHA7ROBImnGZJ
p+qizskaSGzBwGrnancqgBVGiZFNcxrPjS1mr/HLcZO8ba0hsXyXf21dQIWmCOM6
2RlxqJM9VkjocybV4M718qG6+3YWRR/BZnMz1fLh/zifktI2UZGgTIRb2fTsKoko
DENO82X25kp+gpfTiEgaeg==
`protect END_PROTECTED
