`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbVa9CzuGGbgBXvYJyaFjK4XhMJ8+xExRxmft6aBU23/Pl4FxGNc0Pbl+0wAm7ig
BM/X0lvHI7WOkchFCPVWn68dxVyNkGBP0xuxT2eVQWYaBEL1G1rPx0DJrOjXPXTp
Eo6bhE+IT/mLSe6Ld9+InVPe76RqZD1e4bgJM2r7O0heDiLS1prVPrAqlXQmEU6t
KK2QAhdHpbcLmiv09BONEiTWYfooyuF7ku1ncnwsnTq/7sh+SYzR/Cicyj7zoeVl
HTs9wA2ZxM02sEeOqM7Z4JIGGdo/8z5WRGoqw0GD1z3y9bA7BkleEiiDuMEGnN4C
eix2bo5iVb6unvdfFDBJbFnbgwLdlkjBeKsTVFQLM9dyrDjydiQ2dwfD1CWDW40+
fUnIJbOd8ZpnK2QUObxqwbFcpu2Eb2qQBwg+PAhWpgdmOobsx+DZcPlOcz9cPLlH
rzTiNDm9U7cC3NVd2AKSP0xe1XMkama3rNy5HWZ6UKhe0Fh1xZsM1dz34/zl9dOy
8o04BGrzZ4RJ6yyWPYt9T48vgAb00azRpcQkbIOTgErrwkQcz0YU+ysuS//wU9WK
YrBxTd84SA81NkF1WHhwZoboOXsOoE3QTJZKqS8Qmkz4yb6NQfSiD8OL5kw7t8Cf
+QsTlYVwxjVikLvyXk5S9DA7PoXXa63D3awyBrNb6K42dB33D7NLn7dnqHuSyELd
Xli20UdP6Glp3S742imF46c+S/W8GlpYM2cFP0H1ab1AdlkQBxh0NGlq09kThz7u
pSaa3ioZjG6F1GeNiF7UeXCaYhKxbTdR4eSQtRNDLTS+7kuil7ZReJKREFJvn5Ao
1NWixde2YsINk/byUeFV4egOxyQGW8xPQoFQ2J7hT4gezbHnqug7P3wzOZ6/f6Gc
dOBk5X+3m8d/la4OKUf28ek6/udbVG+aHKwIp6pWBaEB2scO292e+GoTibngzlJs
Ed4ezo36CLR2vdh6lqpVFSlomoxKnXEjKeFC1O6/NpTBhIIzmec/Jrki9XOAvkiG
bOUN9ngI+++ntc0DwnjYc2EfplM7gsDSM0Nr3VnXgNaRvTl/ONalYfQyKsXCa3RW
aMDrKVr7dxFfvtbVJM9WQ/RO78JFFJAy9g3g0OPLR/964xaxNrVDz2QmRvoj4v1B
oqzVuL1ls2NCuFIROY9wzUowjNg/fCn0tu2XJE68nbj+Bm6pyPeYtBn3RGq+ivbN
`protect END_PROTECTED
