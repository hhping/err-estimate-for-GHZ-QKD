`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0rZhvYaAj6rq/LKx0KQFqxb6RPOJ/F812fi/tsKADVZbLZ+uMVgo1hP6jAYP85W
J6TdF+J4s7cpaauHBV0bQ7Zrf1m9xF/El+UT7rhFREeJOtDmZkpHy/6RbVXUNxbO
6PeXYG8rPrHKrbBJuypkah6g9V40AzN8Ir7peOmQRds1P2EmbGWiY0tj47KrkwdT
Ud5ds+xZiSUbrO3D7gnwWrZS/OKoae+caIGqyNcuzX4Fe5CkRsZRcbrnAe8hxK+9
Ox3MROjoi589hpfbNInG22VIXIjromomqqsFBymNjz/1Hj1TNb2FTGW1wIuGyPbT
3CP0Enlo2EBenKctjDMZmjvOfYhWT/KdQlpxsksuygytIbB//qoB3RdTe79Nilzt
kiZr5p3ad6GB+bj3ajTOOg==
`protect END_PROTECTED
