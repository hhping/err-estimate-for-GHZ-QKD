`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8S8yl/RPAFOcLj9TBmcWjfzxU7l7ilvDcAPS56Qn5mpOvpTUSKS/I/dCcy6sAkSJ
wDkpA/4uJc+tILDt1ED8Ny6EPRA32D8JZ/8jdpTPzPwjiL7zodpkH59ZEA2zujNH
VQ9PPiKY0PQ3Hj3dRoXC9ln0sOblzJaqH2HcBWXr31SO6JMIqot6f2ZH1qnFBh3y
eNh3YO2R87C9UhxoyKlAyohOt8PUDR6kSwJyHAFuEFpC0ML5wNgleEwz5FfVveki
vAqzCarJMcj12s2/U8oHr6muUzXNOBIjoNHIKgocPVsbrFuNRvBwhXaoxeNd9WRA
itN4B+ilgwIs5vEUnKeLTadF0oMZGfFFWFxsZc/X4mSHr3fhGNEmKbVYaXHqy/8P
W9B1VHARg86cdIt5IoYjmvh9CceBCOu08I/C1150SAvb16GIaOe+Z/ekM5DN8bZ1
sjAa30Dr+9Fwp22JUYeOgCdkc/NfTYg5+O43yMHrpnckn1NC25az7dWSFH5bE0VH
BiXS0cdIbEiRFGBwv1PzcYz2zwoK+pVGuupFE+jz/z3CAQoWvMr+Uy2GXbW1ooHo
Q2TrBe1b+JYR/qYRUJdCVzD52fbU9qXas2PIHfweVlNUB6mLFJ7fS4d70G+UOMjs
eyhBbNjtFNcHnilhbr2rEE754DqbOhD8fKFAa66HcCU=
`protect END_PROTECTED
