`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlEP4WtX1GtwDplgVKXwUJV7uZVUOMy1lrtgczZ+/lfXjeNSzIUejCUopDRtaRQN
Eb5zonZuHYsWg19N+343zSrE2kGsb68akO14/qxmozzx5hd7xJi0HVAHLc6lnJPY
45fddJjRQYQpc064QMEooB9CQUI/rwDQDO9CQQ2geDa2JkZn5ST+Zu7JPp6iMUil
RpPIzeQ+FWH6y8XaCEj5slnqmABFsONpx8bzLm9IRD45RcMxA6+y3SLJhADgk5W1
3zzha2dYcAs5gTfqFCDCcths2QDmogO5fU3AOox2EZ7luABlAP3mPkmy1CvnVkKD
0O6s6Q0yN07u9IOY1Y8TCYZVxiqndVW4Fc6VlpLXWGwrmQyWxte1s5DjGZR+sAoS
uFcJ5+sR4uaNyz3LwQPCOKdcxi2y36E077+g75chZtY/dpLUKXaRbI0u52PqFG8o
xUq+V8AnVQ3h6iNqoi63grGUSoleq6BMAugMzPI+KlU3FZsYlyXGX/WANvviZ79k
G2JZaBuuiOHcnff7NgXiUpNlSj88jmYkc4D3HXTQUAb0jUOyeJS8I2FUjLZXEx9K
GfAiIwQuKCOf0dP8P00TFzVuPWMe6cXYX4z1OuxmdXiu0q69GpoRrP46Fv4L7IQ/
z6Pxz4XbNcgotOl6nDKr1XLl241z4MFZvahvJMspU8NPRHD95Xh/1jO7KtxceHX8
PljGgElQP8MBM+xyc/RIaPEcOh57MgyKhGifpgkmsZ2SFORdsWM7sLm3J+I9tOtQ
Apzq33aBdIFzihNS4fuRiPprrH/5io8yaviTWESw5xYwsBWKHFnLQCKMZTF9e+q8
6/615rcggqXcHBbkTl5qleymS21vjNLbZfeCfE5VPr5W/mRpvw4Tm80FigY81fYu
7uaKJfAM+kF9+BjTaix2bewnK//qXADjpCRB/vRb5lpZtrRO1T7rVSFsI0G8yEmk
CGlXhuiryXsrnTOGzWyG4XdK8ePJUKJ7/r2MLQ5vm8V9ZbAFvj/CPfqMUSTZkKM2
UIIrNx6g8jkwmBTiSVC5RELBOtYSL/o3klpmyQ8/G/nAvW0YlTXknpW/DB05zoiF
O7mU3S0EDwYxctf2u5hw0UFWHKVlU5JiLAljcxKA5bDAB3X5cZGjLGD8EHFHt8G0
cuj6k5CazWmCj/vDzFy+TquTJXd7ZtN4WOiHaDFMysSxURyzgjgs4EBnRSIKKWWS
Q3T9J+z/+twIbbRHtGhofqZjmKsa6VvwDQk/zq56/RXIBCh8qyNvpFalN9wzG1Fp
We74pPNyUdOp0XkWOIfNG0R8C1DGfqRMrLXx/zYOjRs7I5114j8aWqBBDcAPuopl
BcDdWVduM0QSiRlZ4Kd/jz9YjqYOAeuvZr3chGlBh/nHOu0bYjZv+m1UHAmGS+hY
v0gGWZ3hjXUCrJfU/ATB8sYHuqfA3677eUY8QlUM3kJ2AlyybRj9QOxvHtG6jFYP
m/93sUDfPGJ+CSDEufkdTmwQXFOteZEwUMWZ+0+jJW3SXd06oQYKfHEfHUKseVX4
CAbcmmr/mthyPov1qjvjD0wI04omuBd1DMelBbNVvn0GNJCbg2YuhVaaQBA23a85
4aT34dCeXlCZqSqS5lUy/BIHKonDpfG3Gje96DytPhCMGs3iaHqYyE4PMqwLlWrd
z1Fkl0EeRu733c2zUWdLu1Ge7jwT5vPlTbPZfSZ3GB05WT9WQfERbQj2s6kC70oe
QYLabLl2VKVLcwffyrc38cfjcRqA3y8QSo0okCXy+QBk6w4FNeWKrEhOLtYJfGDB
Z5D5k7CZDLV7Eh5p0Pq2KWaYn/h5JcqdgByC8/QKj2n8rlFFwkx4eulJ4CDilQx5
0gBttuz1r9M/Ke2EOv/+6gocdMQVJrJ+7fNZ66d3pDlLViOCej7xMXLn0JVFQDXS
tZsZHI1eMJt/slKbr2QkTtLaUizR5SkdIHfebDaONYvdkXPak19ErjpGYRe+ojTZ
HVMUVDvUDTqjvI6MLQ2KfB9tbRfIJ4k0H3Jb4Z1TdIckm1A0hHzavs8hAmFRuHB5
8d3cALnqAoQgiX4lmdXqug==
`protect END_PROTECTED
