`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0GXxqbQsWehnEwN+yOd4MR4CIjcWccYho57deji2pwKTGn1mAnKc0kmr+pHJGV6o
IVCdN0oEAX5JLkuyQzVhF1RgDx2YekVJ8J05gKZmOI02DO4VPSiINZ2RpCRyf9wq
wUitVHLX2hjPgccroteRVEa3HtuV5prgYlt43LRFyJy8bGB2aehA8bHe4ZzY8bRW
2qZyiAlbrQEVzSmnhJoWu+4SmRiQ/WpIeHMFa6l29u6fvr3AH7ZosoCjftAHnAb5
UcsIBLOzLdxH54F8FJLWm6UQz0m6gerKM5btzAc2v8TAwc79Wa4EbtD1E7Jbihxr
rDjk5/ACiff8GcwARRqYCC8BajAlwo5opyzM3qKcC8hrRhz+PEdCtwz9cwfi8ocg
8QpxA4kjBDht6ASBgxl8lFy5rxSXrluL2tXEoDkGqI0HuT33mLglIlq1IDxpI3S1
dxYV2bzG1Uahy9lxUYfMHe61/AUxF/9rOJofvvcKowdULcvNF7jWlk34OPa8aEy5
ell6Q03oxQDJKhg7N5HiwRNcPXrvRVOU/vPMzNSFqW4AfqaeRws4sTJYjUOGDJeu
KPS4+oN4A8ElT2NSo+CoKAc4QPvmNtsjCV9+se5UD28V1iT6HTay2Tm0RV0MhbgV
aowDXQtAZmLyK92KtLcNw9paX3SgK0+izmLeIjojliMHIffWysT/1Blyi8en18ES
3B3lS59Ml501P29LXCiVgMUCrwhmnIAq33LWM2xSH2Xdoqb/j2IlPRrPppKgCEob
LSBwjefHX52aFahOeFfgtHxolOTlnpYFVxtk/EqxMq60cSx+ZoWmoPXRO7fFC3A0
sy8l8abevtTS0O21U8HkqgsEISWMtQyq/TNV3DZTjgIH7N0n3HbuCWMUuZJVbj0A
92wp7lWPNu7sLOV5YcoNkAGSscz4oM8bdNGLlZhDagYoAYHwhQGpH5wJBfMuV1FR
wp/7Hqcv76jVq+RaJFk/Rjyr2mSIXvjAXcCqKlNIP72y6sHcHbFwNDqJIbiCHf0h
o5VAvBnk74xGOLfH1rlafmPJGZ557iXnso7eY4IFDfkSWUEwFeycXhojqVf2uRlx
DfTqMByz4UxqB9QHOANhZRkqG1/5oxjH1F2CNS3lEiNBFoJikYGtL2NGf8+LHlA9
n6X0mochWE/3z2F/t/4JJ6dJRh8kUG/5A/dqj0Zk8YaLfNDOcTHa1AD2m7ZBUYh7
Zz4ByC9OSaOTkgiNtotAo1q98N0zwRAwcdPBcwN/r6ZdnywYYzF11qyCjPPMPL+w
CbSrAoFl1MaNDaculZUwsWY3c6etYwZxJcc4kaCk3cBEQgcTY/1GBiVtNAkceysg
DlfuQpEqANNRd+WyPrpm4l6rW6Lz3/VpKoH3nhtZe939qtn4nKin54H6BhG1XTJK
YHC7Zcm4b8OqAXDK1GlZ0yJerln/iS67GRTu+uNEGSDdYmiQOBxqyQrZ1mqomE2o
6AbZeHovEyFAYC5dNme1wKszcWbfiIqvfrjzBKZ+9uECypZ6xBWllbWFi4wYar+v
KW1pmzNIiYfIbwo/WyZafC0iN2VVTXPIEKBJvyquj+YZ9I/fp9eBnAevnA2aizHZ
+ZhZW3as6fMbUw9plpEwTwb7NfPhKB/a5s2R3UKhYbKvYkuhtm3GhiU2LV2CITo5
3l/u5KXO/pl2ekMHSQDymZKeYJHl+DQT7Fw9FGgqAPDUF4jmaBHhd6pg+b8eCnFI
zwf4xSCpJ2p+5ILQZZrf4Kr/92ZIr+rRMQVDU2bsKNkndm0wz8fpa8xi9zOtnsAn
5SIFlT+Oll1uSzDZZUEhe63ZNsoomJP1fLz/YNaazjiwIyie4Nxv8Zpzs3nsB8aG
McKqYYcq5FGs4UKgbk11E+07LsLAdHisQmthJdnM69CdLzRfbXoMedqD2WU5Yzc9
2IWb6t57ytoqkeP1IgRYAjjUX5azPWVtk3Wu/XqANrZNHNGzbUolUfOFxmNIp5Fu
sRr1jsAvNop7kqFNg0TPD6smmZRiOGNoLazVoZ7SyCdDr6GDK1VHtVx2C+AtCO33
t1DCiqTiY/A43MwlInJQIW04vcUr60C3ZxU/otbpTikuv69wlDIU9RjXtaPKjspB
twJeeUOfZUeRhz7s6fvDg9xbcj/pjRi9QFhPwPO0BtyCLtLQ8CjA2NQoR3Par20z
No1IUoBR7AVP54uK78wZtJHkQtBew/IXB8iM90tIHLqrf4BrN5JslsoL6NWzLr/s
H0K9eiODzgXNAZjQzQycvaCB4nXWSULm3Oqi6u+EHCDaDcnUh1GbCdbI7gUUgZHc
EI/OBc0NeWjk5udho4AMp/TPIZdQ00MGO9/BOkJ9AZSKmhg73cVvL5sWcHH9Cc7U
bPLy6AWLbc0LQWIgjmYDDL1jCSv3o8fvfuOT6ada2E4Y3JHrs23TUinkP/WS3bd7
y40qc9Vw9dWZxiNw99IsV9hY10YYM21y0uajyBpNR58bcL1XRXuxILo2i5WPbBsO
jQWbPT0fQLh20MvIXuG0EJR4a9hqK0/sewOLSzcnj388MiubIsOvgwQunJP51Zzf
UgzM0Y9QUuJgYe9NfcIqR0bAn6SUBj4NM55cugafyJbvl/K9GQb7iw3FA3f/y/el
lYiVtn/WeIaOI7366oK29xJ2Ozytshqvo+29hxjLVC+F7aZSbEfF5W5rTD8rZ+8b
ixMjtJSX1Pnln8TZL1WipNvLtFyH1rL6mcdfQD0gd3fpkEFGGmmqDJKqpawsfhPG
zDpOtYPLG5DtmAprgjxX18W+mQjK1SwGFKyr2NmH0/5ShvWpcWIm9Gnj0Hyknb6m
APjLp6aSIPn02Oduntw/PTiV74lstFaNN7Dax3WmnQvBxPLijJXb+EPFN3rNRJ4c
qzF4P3kmk9T7qAJHkja8thU7dH7g2VIoHjs2Y3RpCzNbdw9Q63fnS9CpiIoIBuga
MuAq3os0L+0Xj97lYbWY+dwYTcmlDgb6ge35rL2vWky+y4ZUDbd/aLysvPQq8qRW
KtXeqqL+etrmmBAbM1eQxTVuFAE6nc5VZzqTCuiIPDVp76KlwvAtFt9CwTRIgkRX
8J/GXkKF6+mVAZk2uJdmPltjTl/FRme6xWZM0n2g+8N+aER7GfEF/21lGJEgr1In
MsAPUUCyn7mJ0htLlX/5kaKoE1SLdZZOlOhFKsq9wxuhlQ2RqCs9SeBFbd0sV1eF
4HIzlTsK3HKzF6pWRgmYXcsG47Ln9NTfeNCV7wKkVjIALUH4+mcrxJw42+Ao1eh9
0HKkg7TJXd6orvrsQw0YmqQwhrwjmeBbllrvFLjIKOHUcC3rVdNUHoIT6BUKU7IM
hPbLjIc6CBmzQSaJcYozAmVbCyU8VRyhwp7BbcYvnRiM+3woBRoMugn24a7+uM2i
DeT7JbSXjIDYJMwQJxy7iPtxYKtH8mJqyx6yhrb7VrAIgT0dnVKLOw+0kztLgPpu
1yBLZl5ry7VuCv299xEL1tosUcFhel21C2C2wlETmNFoPmwaGYKK9G/s/xvJXvSk
O50J9MzR5uNuyQ4e/F97j+1pNVWF1teazhjQpwP8b1QwNFn5ov+OvnxEcff5BdWI
sRGfQ/ZebOv+j9ifS/BOF3/V5YGz2mVv4AxM8tl6N73bvIgb30tjg94q/kUmX1E2
crQXLcWxV+/TMQiagybnxr2c5lpl4bPx5i98T72gh465y8zGhQUzOevx8BpYDU4z
T1M9zg2nhxT8hYofNjFfQxDz4bpWrSSTp8jmTt1pvgRhJeE4++Jo6Qvpnrt5save
ghjU7naRoIMQEtkoFOxgoxJvcahZQ7rv3e4fMCCZeIPt0qrUwJUqvCaD7E135IE+
iKF5LjBT+N/DWRZmsnKllWE3a2hqdgwNcLM/JzdmcNevxZpQclHZ8bpaMKO6HlJZ
bvoVw6wZqFXXmdvSHybrhLI/Jkmwk4fhy4zd1T6GQaRJVCTn7s31EStasgGl6Wcl
HsPVhcqBP4MI3G367vdN8XgEVOHfuid2JEhkhWbliy7LbO451xVhCGw9tGGf6W5c
gwjGSF4dfo3p+eWvbMwUe+HogKKJ92sFjqv6BewEMLbUbrld/X3GLeZzgEkpitRa
KhYn+BFQri2N37zKNmAv/Lzws+xRlHU+QqfF8KtDbeY+GBvPrHazRTlVRV/MDSWG
ohg8Hhn9e2hGT/tdl1+N2MFxmF+zCB5F8RKfJycq1Y9SFJLnxiUfjBe2rrUGZATg
`protect END_PROTECTED
