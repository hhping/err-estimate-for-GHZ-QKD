`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yij4FL+BwM62J/hyTdCu0FiBDhJzb6uSHmH00Rcv9/RSurch76Ct6LsAZfG7qkML
I8E1LMS0UQngKuQ3iLIHjHWipzpocaxxjCsxacOqjVFaUbO2MrSOvYfHR3VxMHct
XgW5Q8t4sRFXTrU9PlHaOALqGwVAzPcW/0LIExG0jTthvn5WOjze7XntRVCElLFL
U79YDqPZ7dQj8gmYaSNyP0vgSIdMtR4/HHAOPPn5urQYgdWmZTfp74kG2THM/LnV
g+haLNKG9RsnloSKUBgdFeEkO9V7ma2D3D86fjc0m8suhj8xRgCUJ4Y/+TRQjkaw
BIu2njwGkfKSTKFxdWecswfMiVqm0K9F3vxQJRiGAloUE8nJOIsjbzrcl0Q8iOqh
JSEn179EQoFA7xSQF+5AhOdewrip31hQOeKbqz5sO118v7uZd9k/1talx9yC7Fua
dYR7nLmJ2BvWgf1PQ5ES4zzimZxlhTLRQ5YZKDCJN3FQ2VCwE90QAiMa58Rwb/Gb
j+hJWxVVPOL+kjJILSpEjkuJZDyRBjQ9tbjftztYSwTa9Yo81U9BVT+kR+oUKh8+
jrPe3FG+TPsCJq3QZrPZ7xm9v6r6/IHLG4T+0bn/nG2KvDgN8Q5Kzw7t2YLLCnq7
93+Y2w5bV6R31DXlKGu42UFPHfxRdGmgzu+KwZafhWVMhrsKDbbtrgHKIsWDZkfF
VNhit6zTS/vSUFn9eg3Cc15I87kfWAi5U8aMG0oLwKfRjLHnKi8nbfjmCvU0BwTU
yU3aAIIYQribEXgySbp0MHkYoz6o/kzGG5Stclv0rvbsbEQ3e4yUlN96ZqVZetbl
JDWwKFnzAmovC4nWDZmOGrrek25SzwV4saKGUi4bwLPIk+UoP1PJ1wMwpUboVLS2
ZUAc5ruzivCBuqbzftj6oqFhtz2oXVJjeuSQFNekLxcRust6YRDSPTSMj1eZ72PP
iTBoRLizUfbTs41K6N2aSfGtjHbibM2vYBWiVmvpRgGs/2uF6oxuQSQl1Zx2vbOV
VOJH8gsb9bLSjvG9x3xXw/jY61l8JpiIl9n9SkfVZxyXY4XIPPfB3HShxjRolmvd
qk4O2kY+zbZ6p8gQb+4hzJ/cZxMSWdF+Z5sDzf96oX+7qCMNdT95Mhz1K+Cu1h7u
7RYXJX8ygedLDNqlUzaYzdu7nvhq/OV50OtReMVXkNLvJSRv5z31IQmqpThVBa0g
Nz6+SPGdBvE4NKiccqPpEAOWjxT3x1qLpKcNOhOmkK9M1a8p2HubDDwa/l/PH4NA
7o7pKL9hjwgvWaIY+aKjxpWjFBKtEllqO8cXCiej1Enn1+VQ60dCImQoCbuVH2D7
g1gTHba5kLXHEZ6aUT9OfL2W+vW59bRAhz7/TDrktlr5OFtCyZRKjkirEmK1aDDX
ngf284lt2FFulsaZdRajsO3J4OeuoQiMdSXboHDOSnKUL3wIEjvRl2bbu303usaP
xUkx2ZKrWV9YF9L6zXOYp1EWB79YLM/WJbvtPhJmvxsA+JbmQ1xGG73c4eThQR5K
nLAhKu0w/OJD7o3CMzcQp2K6UB0Njmm+8Ed5Gl4Z+c1S6TalODyGPCqafcaEDyES
C53ECgfq/uMVLiH0e7fmFO42c8r02ieJ+ZEHRKgK7ZfM+e8p8cBeYAlL6dmbb2bG
3+mjUZfCHf+VsjvNvZ74IeDuUGn4X3wqkY5CyvC3P15k0sjIs8CWEQLOFHPxQxU+
ZtSK8dHJGsG50vrVcI0bnKlBXJ1GzDttiIC9f2IhN/mM9ni52TNPgFN+TQ9HTEAN
mqOZrb7xlS3U3xGqdOL3P2q2JluFctKDvvWMBe2/21zhjWi1QN78GxEMQWSHKwy9
kvbDOHzFUo83vW5yRFRkLoxasOk/RXxEu1Yp9RFPH4hc9F4RVB22+d8CMN6w07ba
VIhRGpeZOWXoBWM0qwNPKqee1SO7IOxxxqfGj1a70CV3iqY394af9zSAlRR3DH/z
9RJ/CdgcW1otdOQZuKyZxjKa9LFe7bn4dX2kfpBJgcmhgr5IQObys0t3BG/mSOcf
4BrvtHUNyFGii1eAhrHlPdQ1nWfwIVxqw45JlxpFh/u8l5rk1ip2MP5UF7WTGKCr
pie+r2vFQAhxA4VvX124CTh70q/wpHUvqiCaH/gsg2lXLvfFR5dsuIjbz8fqYtR0
7gqt2ZIDNfxkKGbX3lntXz4I147UIjK49K3Vmkp/I6iOd2TPFUGLyvmaULCMO2xt
Xk1+OxwJwQoCFZdFNqKGiAZH0iwcIN0dwt9wNpBKm6SkizN/fSGHlbSbRt9M2PTl
gdb9JUSOZ6b9h/9i+5fFzx9mRzS1e3fb7no9CYlC2RyvdYc7dFFM9DQhHU0F98iy
faAFq02VbOl6QWUW78o4iy13IR9gUGHoaCxtBKfKffmatxn+XcnDgaOkLnr17RCE
KxU4KR3r6mR/VSODPZduggM/kU4YorXDz/0SD33IVW7uyugkB9h77R5TOQBKI8Uf
XX/p/ljyiGE60r6P0Tt3+ooZMHql7gjHn7i4eOtyOQf9RsVylSW7q+D7CuXlFZn3
hNVJWCrmVHfGF4Ilg/OzF6TKzMeV1G8/kfEjU3k1dUbIhXqf1D8rRJubW3uPhXXb
c3ZPDY3ovNTL97oQ9fy/c5nzCTyU+70kqnap3a0Dz4FeXdQ53eGSq2hsrxzPfcG3
zdDSSnVrffvmQzF4mT8jnTtdTphfJzGFcoCbWtrJ3ybQrTq2j9muRUzUEXwdi5Qf
IFpizAS1CmmnsOCRmm1Ts0Yy4tfGWADZgHB0oJsQbaHCm2b4wi/zVtpqLKTParKh
pfF6g56LzUq0KP0vj31a6M8o+wPVTg5Q8vd2JpvwI64H7ioAennarrwCgr0wJAAn
jLjHgXAYMoBuet69g74DwNZ87emkadMm14wvm+dwZJ8CDWFl6LwlC0vP1mQ6fAXj
LQe1KmliW3Nfz3UROQuLIuWEmiShSIRD58KN08WRY6GxNrI2Dc2j2J3TE6Tn0ePu
86i/bRCx2B109zg+mN5sKITmPuIOxHlhKGKdh5GcP5sValV6z6NTwuuRPRe/mB8u
oWlcktYkWdJoivnNXtUg1AQtNYXeHLVtMhGQuYMooSYXJXg+m28b9EF1au5Mr559
uB+3NmGfjLC344ed8D+CQiq4//yH9c+QYcBydPbxRFRYWzWy/Um7RzFtjPBDhxfH
d+Jl5EVftcaP/Fy89ROvUydMlKTGuzXJUkxSn742SFPhL/d9xQR0JyxmEY08M68g
RJrBh1xugAW/ulqm7On4UAdgrDQb/juzXasklVpkuDPQ2vYSSsJ9hDJgCn93roPA
`protect END_PROTECTED
