library verilog;
use verilog.vl_types.all;
entity ALTERA_LNSIM_MEMORY_INITIALIZATION is
end ALTERA_LNSIM_MEMORY_INITIALIZATION;
