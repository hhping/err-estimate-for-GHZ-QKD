`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ocqr6PIcztdpniJQOTlGRkYKJqcsbJggzdXZc4t9vZFa7L0BdhXb6OZFIclWzX62
M5dsXJyrDeHxfuY+2H6fA6l6fpaIkYvCf8O4ZTN60rm011D+J+2Nqo6W1K7/9TRe
QaL19g5iYv7k7LMRtNdw9bqLKUbp506E4wlZSXD8m+5LTTFw3IoZYSN5si92bg51
g7rMD5Sb8GBnhQPckpDj5F4Fa1keNvlvQSEkc7oOVPhNkTX3q9dqz6+0BML3SNxY
nHkO6H6hh9Y7Mfqe2PNoI9+cbMX/PrtxB759S9jzz3FHYwDA4zSaKvJ3HycjF1ve
aw/515E0eyggWF0tqNhwcubqe9YNq3xXpauYhxDGtEooJNYExk1cz9DFdXv0EgJs
pwh8ZoJRqHFMgg45pWpy1l+d/AC9e5MbBVhHMtGspC4JhCmSbCMHLo+9T/NPcEvu
51+8SWe3x91VGuBR5hDR2MHbF1uzEPHEek7bLlT9nRBCHRBtZQ36jnCQjdMlprA5
lnUPvAx3K1NjUr5eioseFm8TKOD8OVfho+kEu/oFzK/31Ui+2+ouajBzipKL2r1F
XDy1lU2BI7ZXlEMi5P64Po+jAIJ3ZYpRSxmHe4TecJaApCk6Soks7Yqf1z+858Kd
GuLlV4fLVahx5yhRdY3tmVIfbruiiAZw9lPuXeUZaxQaUqgntOadNIoFCJSVeoTv
juyhk1ZANAjHnCBnbyUyOGk9u3IFmrsRFtjeGc6Kc6FiUsdzxOLo0uzC9eY22+gl
KImd4mdi6Ayy+rhM33qEONf2w3sRbIKAGsWSN6WPkf0RqieGFPFb5pI05wkk88Zb
5ZDSu555Ms8McdImuJt6a1pqFwvgei/QiboAwU5M1cntbR3J5W7eU4gZaxSK8xh0
sYKwtz+YXDcDyDHsUhxFi8/FuVglibRfWa7t5qrj/SPl+uzjw7gjCgivdywV0Vz+
sYEvSOePPbyEeJwYrpISieAs1n2ad+ODc0vddJiNkQk+EsL3JklnrYKm/KPw1JNy
yNbSZNOzSrnLk/yfJV6tgv0kgYHhsADaahrPFZ6QSAN3g0tziEYagPFCQUYOh93N
6Eo+WeWLBEKnvhrvReV6/oWZSvzaLA+IHJzVnMFEMYjE5Yjh+yvL8QV2Y7VsiIsL
lq3HKL5uBQR9p2+INPJFEmLIuqeFvZDl6kCANjGPOLul4GRFozpVSY2Q13yWg47M
CbUP07gr2Zyr1yxRusMUel5iQwjVcj2kjmzu/XFyO5lACfa5fYXyRkDbIyhxz73K
+cs3klaPxF2nM+AGdJOOCLRhQxVdV0U66qB0+p3OysmaeSU01zOR7w8PjAsZV9RN
+nw0KFR/56Yxu23R4gr+wohhkSqydH9gfmkKjHuhZewFEiYYM/SJDjjJVFZu9a+K
R0DGmdQoNR0DwNr5JpGmA2qhwiTo0DYWmFvgvIccgo0c6a8OyMm04Cf4cHpUrkOq
9pabglmN/s2wOWJwyi3QerSnARkiJ+Ay8QHc2CnUCpV5HTjZBMKocGtPk5yspDV3
AGc43Amm9nTbyjtUzN4p1cWgMPw4i7Z2X1LYV8ozj88ippOn+kAfLH5C9YfghxAV
4u+H64AUfsuuslpov1upzj4H5cd6edrlTvZmEpA5NwMeaHlgdPPXY1SFLBkzJgHP
+JI7sCrOzH9lComXEhkd4BFTwg5FU1ydv+7NkvNiyvI/lDjmACTsA3LgoFbMUVAX
NusfD0sTkvJc5B8pJyjRDfrSnFRbv9PuE40m87FkvfEaN72HlMD967J+uZQ4EzGY
VN2zeyidSOk3S3UoEJ8i16PrXj9T2YCPUdI8Cqp9NikIEmcKz1d9Y8wxHTlJIfTD
KGa/Iq4jN8grW1jRjRGGCBh/0eLFF6kS/WmE9bkYkrmdIPG1xyzLeyqd5+mXFkN1
ejRUyPMfe3WOYiuzOducnbweB7/fD1YFZI/hA/iCGDweti/MORxEypwf1vNfHgV/
HDgCm8UeHOzEYE8IBG9+vwcn7jfjSZwYbr3UL4agXTqvZwXOZiwYUQbzpmCSvrs3
tmcIFe2Jo1b1h6CUS6QO1/tdT5mhFLdvtmqM7tEeh5R2Z/OHLE0BQtnQThoIwe1c
vWrcqkUDwC56ljgroWxRTu15r+oUOME27uUq681Bgd5aGwynI3S95cjMBRIBH0r7
ucUS9H9kVmH8sKuQBz/Gu/yZwQ0GO/FDnZU9FpDQ9SuG/C1AzoTrWMgNVSIiNAwY
Mq58fu3vRrUpBgDWu8XinEy2awIsxCk7laU/x/QGociqDUZfoYFHSgWn0Z04aHp6
g7Kjoy70JOcSaO6RMHQn42KaMsHZsIgnHRvoZOUuW5W/K7vQR7Tm1dBXwGKlibMy
F0hxiV0EIFKtAyhCzNUQKWBHYGxPvg3LIh2gnwS7asA=
`protect END_PROTECTED
