`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
baa55XdYbNUX+2IaICtQq1xpZRLycQC5O71QG/8RxYE0nQfa1c+XtQkofw3jxBUJ
NvCxfdn3VUmFD7dCdJOfV8n+hFjQF6J5u9N/5AoBh5VEqPmzVF1iGcSCU5mMQLPG
iRlcOC8cag/PAKHbI9wwyqeRlpidLXoHQUG+JTjYP9P9BJJjtfq9ov7jG4B4indo
pEnnqcf3vl25fNxM/eARlGOicS+BkecPeFWgMDQ06uI8TO2ohkjvlEcmzTiMx6UC
dltJ7q/wyobhszjBuhpLDE7eJRqOqfhX3bk0lsxlMzdke27rF/KgS5oOue8ZbdeS
sjpeGxN+9/Fdb/6pWzXawmbk9xYePpiVujISftVi/a9NZpavWBZcnUt4QzV/FzQr
pXQvm7SEdWmoWLoyxA9pfNl8OWFOT09euAraeTe8/qrxEkXRQX70x8cgWiJJQPO2
smfUwsLCoNITgJsy0XI28/DE+QKPrhaaLf5QYHyL7vGjl2vlf0Z29oMUfzwN83vZ
wwmVpFf0t3pA0VJbtq+iOeU24T82XZeZoRZ/Y0Q5P8mfmrh5EBHg2hSTAKhIGlZX
M1C188KKCGM57GIAWuSiKHEnB/byVNvT/6/h5i+H61JpH+2ii9rufwUNXN+SXRoq
ClKYqaFm7PkMCrEz/fJcQa44zRznxd4+7T9jEz2pR4vRPFfLuruEthdIvT5Y3iht
UFpGAiy6zrzcL2mg7qDi40pioVIaLf8ymkCZrXnSaJLiCB2Y8NuvAmjYZYL3017l
LHroH+D3c7s+ctO2jKjQv/q04zmGMwOdk4RcKb54Ak/TEP4OFmh7vgQTG68KxzCh
Cp9JDaVUy9vW1wFReVP6VdOMmwCpZG56dW2qJHkmjW09QcsIWOmNuP8COtl464Rx
pI4VZd5qDEMweOCcaQmIKGOlwM/lkyftQgSFjnjvwhmOO46MfBEfmthZcyUIGUHN
cxiIXfgRyKUAtB0RZpghNxfziSJ95srqOYJU+iUpe4z7DTqtWv6AMjkFQzbRkomC
q8PGdsdtNIuLrtwbVyzbPyesw/skY08+zUwUnnHWK1gUKgL/3tNmeQef0MTxGSEd
luWj9vQxz7qp6ALYh07tFWC5MgSLGa+3xNebq+n22ow7GJjqcMut1+PJSuj25h5K
TiC1bajOqEJZIAvQ1eJLCVtccFmIlxITMsoskKJ5ysS9rQD3ICpW3mx/Rwzf2yc6
VQhrerMq28L+x6HV5Zs8FHuNaPUFRh+RzvN5KYKw9RzAXnhOqKqPan0BDS98KFVN
qBpGG68p27MsZbJGo2ZDiy0iy2kgUfzqPKefHYu7dq6Sac6qPSgIUvbA+oaofpdi
/LlFuBzABO4p6H+aVseMbJTLhhfBSHA9KzR1By4vw8xwF35QF/gHJfg4TZuw3MBD
vj/uSc2oNU3WcfJPLFZB7t5R1t61aDFRz7Hi1/6to1KXD9jnrZw4K7hmGxBBurk1
cR6ueCQ+eeps1OA5mViKTwHuw0ImwYMQ6QSXIsio/sqRfgp1I4TFYFjIx3xZaNSs
40giKqCZfnLW0djdfoezS1FjcLNHbxPCjAtP+O7w3csVCdLW+Igd2Hy+OcROp6zh
GxLGfM0KdjyA1VJvFJYfR0sSauLgU/wd67R9y5GLxKOgOd+vOlipTigcVeZ4KdCH
CscPE1Mtr96F6LwxyK2iBn156yAExHXhFpNK1gBz7vH8PuPdxV8BfUd1uKw58XOJ
56fXZbmrCwPQ7kRaDxq9Bvqrow1c3RqdZwi8yE3XL1o/Lx1qk/UhoYTr0sJ4fzlk
Scao5V/PFrOS2Yg4PhsjfQ==
`protect END_PROTECTED
