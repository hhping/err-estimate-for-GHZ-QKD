`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjTcJCkws19JmW9mOPnAuRUn7HC5xgUQr96LjN8CRfSssL6jC8Y2WjWq9Cukrb8/
ta7GRC9fI21ILHmcNEY5Jd/o5+IMccS2pz2Rm2zctqqKRQj4w52NSRLOR5QxTgLy
HnvUvpbqV/rtVHUt0VlR6rVSh0n+14KfYI1mmzk5mOE268xaTv06cu8l8ItU9gEn
KNUEGT4Zy451orIPTfusEJSqp0vvVc4RTIH1mxFPqXsUAXVx2mQlX7cU02gQ2I6y
22Al5E8O+qR7Tk2j+2MoZlh7E2mmMDD8wEQDcLeVsP601N9UnLlzkknOI9l/fpzG
1i80QItKY6B9VIXyYinvYGtNl82xYJuXBTLKKleTIRK5KAeQCguSsBkSK5rNO5B4
Z2dxFHsTYOvUhfOy/RNIDvx+brp++idvgVUQCb9AFHwGxg0kSyCNXxZ5jXfjWO08
xHL7fZSYbGXQpmjC269oqjV1L9WL08EmXAnxijCvxYd1eSrT+actQRgl8HTNFbDe
AJyfcyW/ihT5359WSLsuGRPjCGkge+iak//hWg3ZoFmnoVWdJnrWihCbcHyTv/Tz
Tg1DY/qp+SaPacg93b6otFPSoqQy52krx39fpQFpGNv/MHHppM+rpkBb4g6hv/dB
ZKLN75vG7Kfi19ka//YfZTmqJotkwAl4ZrsKpL2eJr+iYbyXWaNxci+iBVVVia1P
2x7jz4Gn8QNLAzeYSOAWiKlsZ7t8YofH/b2LIiQRs/aARddtBrtsqXcib/NtLhyV
YyDz9mcjFHKaZma0Do2DZJrIpFjSlqJDmguovNru3+Gujqp51kLTtZ7erqlx8IM6
K6NKyw4oSdOxBixl8qHIYnqt/IRipmwmA7A0PBS4nRVFZ1MIztsETzEfogo5I2qJ
KvSqdUmP3xt5hmuBa7Omha7t/iwzVTZ58ysSLsEMXyhgbVtr1xOrwSgw0s8djz0T
l4Wtlzjza4JQsneMQnMMO+z10y3qMcyFZ6sORDDQnSaaXfLYpAzErWNfTE/jLiip
EDpCcW7OKl5lQ4YHIZ0Pqj5PayjU8LuCmTZsSVzgAYNHqDCHcjg61zxhHp1+5kaT
u5PCpVcs9NxLENgN4xV7PeJueQU/FKrHpzBg65HF6YWT4caqJRIO008JbxTL170w
f1tBhXxaaqFfASQyVecPqBYJftlKWvWNU2RVLfXtdcJCG9UEUkRx6uAEqc/TCByv
4n5JOBd0B+tjaUWKA9Sx9dH1gdcZtdxZORHIqWuvhh7BW1eH4gffTj0t4HuP+jZb
US1uu7bdSBRGxYo8mWWYStO8yVe+bW5ktRUxowJWhOr9K/Cmxp4hHs2m9zqcOB31
IOQyjL/i9OKKYsfLAn9Mh+kTRynSBbq6kFMZAPbQUbittC6FylsnHeGDvrNLaTyk
QRTD+QruI8ZmajRYvi/p+AoswDw8DWjwNxFAWNcwrTk13Da7sCpHXexp4V4FlEp+
+4fMjuIP8Hoe9VXCeJ9JvgW6AE/LNLoLb1n6BJBZG+fH7Wv1iWqsEYR/WhsV2E8G
A1FysrIyVKer8CT9uDTWvZ/WmnD2PX2fqcYzWBUhseKzsToVtlNKOo+pBGAe4rA7
fyX1IqDmWgIuUQfq4FXqEHfUoH5inslUBrpLtBbmVaTbyZJtpgv5oAupxHLUzGXQ
IHLZrcLQVE+3J0CraCfTfJ9J8txJeurAIVTNw0jpoOob2n8+3VeucmPJzLndhsFw
EujLuq+kemUoit2RK4Xem4xSwfnkFs3izHPKJneGfwLquAQDLVdexV5XZJcqGqpA
umQ1SBrMTpEQMWzyLmflCYl5Uhh9QnaRDdIp2CjuMxkwDB60RwfsWzGO6eNp+6AK
qJ/2UjTN4SgmAyMQssBoIMF/0FHM/qWC5EHvcEiJ8uSz062+ZJyeyMGo7ae0CvLR
PjjKSl8DG0Gy2rdnJrhwKR5li+0UPHOsshQC88YafgQC8QD7jqzdUCLrZfwJSX81
VQem5vO65TuFl14Jta/72d3YgnG7AsAXLXrG6kJDs5wXMvF0P3G5AuYuFFGSgRRK
L6oCkpUIwCMn9ba4Zh/C16BqoJEIG98iZrS5+UJvhJ4GM6068MNMlKuzvmzB7zSF
55NQgouYkPB1XmXJ+82MnvIVDOXtEfYBLyMTCsAMIvlFCqDc9ij04JFcOS6Qixs7
UuF6EUGtwSbyVmRY3PPPVoTszrTKRUy12F431nVxim8S1s9IJO8iuT0fsRYksgCy
rXVxJjb0KbVbSKOhDjnPs4C4x4CoTWmXVHjKql6jt9zQ5FxGXs0HtX39O48rAz5V
oTU61p2pDgnPBYUrhMZ5jz9cfcHyVsMkeA34cGbfRhY053Ia/DENYOnAO/FSZ2M0
DXLxkSKvIR/1wKfgWIsFKgLelRv61VzNSlP/yDCdGAmR2mqeNSSUS+G0LWkFTl6w
Mvwec2FOhyxMnKbqGfVsO6bsUMKaVm8qL/ktk7sGztE55fsSAIVR0/fYCUPVXecP
WurjfnuwOgwvZDLJzb/UNJfzZyzt74zoeejxe1OmxNTp5Pn9lGuHKhKccOukJtet
uL1jvBSXKBu3xaFOBI3MqBcFBoQiqo6IQLh/Z6sJu/H48M93tlyi1CtKct5zH9oP
6g1dHtR/dKJNuMs3iZgUXBASf56p8Mhr+633rCvIbIWXq2h+qZwtjqudnc2QLH9A
jhe2Q1mHGGVPLu7FGM0e4CJJ5AsIRaazQSlrgAJqKoNMe2FDCVw6L6zz/mNZeiFL
HkF82csetYa960ntU5xi2eGA0zyOoEXmn9MQV7ZHDMUBFsv69bXnfyj3WLHcLnev
wJgPisma/IvvtGQkXGQdBByNJuvccwnwHzSJdm4O7TcP8JSgUx4tVRzy4wfoZJst
JkJ5bKb1mxtJUW/Yxb+1j/bKj5xwgVk+fOk4sF2lvk1KU5857O9/vvBh8u14kFCD
`protect END_PROTECTED
