`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gaK5KoYIbrTa2yCCsf+lIm1oam0MIQJGim6zSviHcSuFaJHAMULVDCsW89EkAk0
MrLrXpEzE3Rj93H9syoyScZO6dnuTlmzlC24Lv0QDuPx/dktDwbvRGuAoQyZWK0M
UXPpnytswvVQBQf6iE/kydotuyHnq63KGN2hmAbTHVzZPqk3pPQdYDJ5ZMd407Dk
K8vD/2K1R9ilAM7aaKAIsbOw8eM1ojy+x8nMpGuWyzGu9nD1LHHaMpd2Qb2++36E
iwdAe04TXgMccnJ5hIRqYzTZbqC5xdiWURID4WnOmQCMOZSwsezcQjOSHHnbgi5r
nHPlrpOsfkdkdGi+QlITulA7Wr0pNwAVP2kB8jC4R1XRn3aRdG4kIviQ2o8noDyo
d5Q4f3534je/t8Q3mlZsiOShzsz4cuyN+NuJXDVbgBRR78wELitlUMdKAXhhWxCD
IGT/Fjlsq5Mj/YCJsD10GVyQobh5WQqm/LpdhbhPz+uRq4wjN/nzepoSIH6Mp/p0
hVTRHaZi8ehKFc/5zp9qrB1diBHO91Z4zoPWaX6mbZ4lDfo+WwR0dVYBvFKQAls/
z0/uzU6CTtHrpUnqSCntf/U89B9EFmmmjI1tmGEgsrgM9tsRELXLmr9WgOHOq6kZ
8QTd65H3mu3eQ7xkQIMzLQ==
`protect END_PROTECTED
