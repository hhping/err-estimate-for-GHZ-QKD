`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9TbfiMFQpYMAAbl+QQKB5sY1CaWD4XTcPJ31iieHRaylJXpkztQc55lgVvlZzx3
Xwqc3jYEHFCQhidF5GGvcAr8C20lBVszlg1w0tAhyOU8sKuUE8aIIWqxFEVF0PtO
EAR0Y2SLeJU5kL0wwumGPJRvQBdqk5+5+hkrhRGtVoEZQQ37zS1KQWPj86Y1XJU4
9CqXr2ji5AImPGhYb+PYca14kPhE/jExzH+o8afOCAxWK/6n7s43yCFCirNTddqo
zF3+7+5d79NJFwM2Z0ZJWqINGZjhPM/r4M3SMClkct1U1HmkFWA1CwDfd506tso2
QCZSaaHwLfESXDMXwcePJ1kBghf1IEVrTqY6yWnQ8JSbLwJyC19PHPswsdVzoVk+
ElMnQ3m/9aPrA0AC49ovc10+3Y9fIMBb5LxoeRMM+PmL1W2qnYgxtMlE/0+YHM0V
8+O9ZgMTDh12Ddgkmr5Nohz6iUY0CLZsxxPGWCsyKWjBNQmfnJI+7sAkTvxJyC33
AAgWKGBaPezJsoAc4sRLT7FSaCQD1luiqRg4HfRhV7lhumh6SbITeV7FhuGaNI9N
ku8Z2VW4NDd6qyZbwdWniQ==
`protect END_PROTECTED
