`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKEQOwFCif+u6RwnUUwdVXLXzYeRJeKTWa4DYVrVfGZOOp0hkgj+XHmz1zFbOlFf
5dqkweUfk1jwzt/jx7B7poMhni5129O3UT/vH/vWsiYCJLpD5xHIgnjEBTno03od
TjMlYPT54KsEkzabTNhADZClShqpoZmCxWLLHVbfitvLh+Pt17wbWcJC4QWFBjQp
7+WpKNGGQbasmnUyoHiEz1ma0Eyqp+jm43s4Skq6GRRiQ3GiNAsFtZ9rGGn+m6/l
VwjMM383fMfKYDSKCIanTgTwN7ZLvd8x8mW0TaQTUBVSgm6xJxWJijHeJVET+T0p
mXvsgZQgY7/THIrhmsEDKEF17n0qidByaTqjvyRCvwnfTbR8NzkDUZ5UkBjY9WLQ
pRmwkPc5qaajv03xL7uyBA==
`protect END_PROTECTED
