`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmIzaumMsAGfIHhet4V8vdZoUe9i10xZ9HhE/KxGEI4REmpkXbXy79zOyJS80S1U
X+jyYH95YQiwa7Bknt1QIQlC+c4lWMQL4KKldOIAjogealinhIY2hvY/ut4c/qiS
o0LXIXcoHbZBO06r74LoURfaGbGej1hsmeO+ZK9JQ/7xVgG8HzkBYvwye4qjyXYi
h8EDGDTU5yVOnYCwJ6yygGL2anO1TrwPwKfK8qeIzExjHoR+r/Xjf3swJOD0o1cP
mIyzHByt8vqknEPJxiN99iogOB7GpXVrCgcOUp5a4xNMyJ3HbFXlHKCSJTln34h0
Jo5EoW3Fgs/WJSno0VGWSgYtHQ1TQTserb50UHXheLFnlTv7rESKZR0EoZIzYCyU
a2Gotdi4bRdYOicyc5pFiX31k9NPn/FmdnJm2INQsXf86V+S2YVa4X8lSuGrAp3k
+0jStbYacnFEldc4t6sFqDKEr7orVY5m60pnHgWkqA3nShTsP09orv1fkyfkPtGk
jguvF4aoOHae5QTtBnUETWW3eeFZldGxCb9uvC+BpifhzkWDrHsVvX+unvIPtG6a
oiTBComeMT4rel/8i80YYf6JfZ0aEep4GFyjlTN8kfmLYGF+kDak/clfmpusyfC4
r8cfETnayeZH554XPbsQvWzmes7E63new0odMY5Nz7X6Z613+1PYkpTjoyNIEZH8
SLUHazN3TjQLebvZYVW261xKVo5Zsgfm8McFSLN6RQn+j2asjDtJXHHhucDd/4B5
+w9VJhWpiJz5uBaBwDGA6UzNnN0ufLbOMIkVIuMkQy4pyAj1ARKyIfWQHLCl99vA
9iNXJezMdMUeNGhjL7nYF5DzIIc/1feUU7IjzSDDUX5kZ3XdJScgLkIO07x4UJwF
mkG6Hk/D2M/oJYqYF1cygrBxHWPaY2yUnHZI2U/lQ1B/BO25cwTL+k4eCfHJJzDl
akBELGYt5V+N9X0zqCgfBaosYUpmMelX41FsYlnYFACaMa7T7FaYg0T6gawJRfT1
O0g6OgUerlQN7yMqwyborzc7VGSNjaGeOt2qi7ixnCl8gYFDlDMbJWGIrofSFRp6
IxK+X2iKsythF1ucFL01YPFciBaPICGnpEjGQL9qwtEA75HDNynhLz0CKq2DSBvn
8Ejt8juc6l2EwpETAVfZewU31S6EbKWyvKLIm/2bq9I4DPJBPJoVxGwgxZcv5PLR
no3HWqmkNXPZyp5H7vkeXkUYsFwi1ccks1MbSqN2sCmMwR+YbGx6dm835rxOY7Y+
P65ng/YiSM7N6ZlxiCFNpsf1pRV/ZPJEYcROAmt9ry0Rvx/AMXhwLWJsq+PPuSVi
PTTRNh9e/7cyYtnROSZEYH+UtJ/pM4yndESHrGTpr+8Q719aUpmLoo4iRKRovzx8
grLZ7LoeRV1zcSiDYaIFU9ipwA+fX26KZy/Yb03+WHI2iGGYWmmnT6+k7D3HRg2g
V9nCgDeZxurSkD90hb0tLFozNktD/kZfOIamEWYwGR4TYdwmFJ9yy+YQsGe3c3qP
56s9r9Idrn7l2gjKjh8K508XJQ+9keGajBz09TqGek5RIQM1FLYLLkAJprcWejUr
K98zLUde8++e9KmyBzjIs83dArO/pc2OL/Z3ErcjyxlUdyragMghRAlXSP+J8uNf
`protect END_PROTECTED
