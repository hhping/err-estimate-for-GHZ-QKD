`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+sXM29TDU0l/egQhdIpVuMOLtsXYIgCbKNrvqpl/yVyyOabIPX+CKc3gRI187BU
aRE6kvuKkhyUVljRXB5wRGvb4r0gv0b2cgXkNt+mqvZu/AD4//q0eDSM4G7bdlRE
wVVtlvxEVt+8FX1qC1+8NeCYVN/tafeV2xdXY75Lpbh6lu/+1NZBgmhqKH7xjvxD
Uu2bsYN5EO23Jv1nPRrecb58n5H5mjohMkBOaPw23mVDM1E6ZOqYP7VJyg2068Ag
iK16KAV9p/kqXIblDWqYdlcqSWiYNvuf/R5jiW9FONhIF24oqm1ffHobn3qKHsur
PlKBUTGg49+YpIDA9M8CMnkW1RjvPDtJ4YBA+Ekr4Fu8zY/UUlEThvIYf7qS6Ahv
xcj4/UiWNIOMh+YFHHKDhdiTvg3dAjYmZb0bwgRGzpnuu2ZHP57aQQpRtf1xst+1
1Z+FToPMCS0JH9ubM899WTYUEhlLFlm5Flw+p5NxySpYnKw8gAu4msCmgWtsG0JQ
wnluOx1/Fqz+rMUkfVfJgDcdDl1XlQMhep9QO7DOC0RaIQ7byClxKquDA0zq3FSJ
RUwmzzbXGkVQBz+9z86AOsZ+bziVtx1u+nqPXoZLqwPsS7QkscULs/xGi1I+1P9K
pXm8ZwtdeD02X/h2gPnVpJiNsHJaJGS+VXZhA8gPp2M=
`protect END_PROTECTED
