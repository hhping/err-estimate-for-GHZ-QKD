`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOHdLB2cqRZO5ZDIYZ7zJnDK78+LOlKnCyFtCe9Qca9+5o1cI0kw7EA85/GV66x5
AB8Bfs2PCJeWCDIBbKHEsiI56xvKwimGvDbykDmC9JdgPXQ5TP+O2Yvpp9GM0Hpx
zOuRt0Wt6OP/xs1nZeTdVIHNTC3tA+Y/+riT6Y3j3ibtEPHvMGOD/vT5MDgJ8E70
1WtSoAekKk+QOtvqxM6xGXXqYyKEwzZBQdctBy2miUwnGYrm8F2QacB1znKjuQsI
D6By5kv4Kg/CJV+sUZQ3KqD944mCyuCYt5WFQS0z+W3GKqB1ub7SWMN4TOSm8JLy
qeXcywhgDJuNt4M/hI349scHPMsc+peLUau1Pxt5dmFJ4geZgsG1kNYfIp5DZYz1
oQbqlSXjq/HI+lRuNvFLe7+DwkXeSPGloT29FfV1U5Gdl3ZMTrz8IZ0z6STLZfo/
HL+U2yWM3ZJQKcOUs0TKApx/3Ykst7b09AWVTHuo5cl+If+q/QPG7KQIbKlJvuzp
EQFk+OVbL+x5fqHsqrlPAQ==
`protect END_PROTECTED
