`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtPxP50tZ6PNuM/PUd6epBlLWpkA8TMDWkMqJXjqOpIIp43VLg/inzl8NhUMuz6f
GBmGvpVRJGLDR4xEZKUgIDcJ0KmUC/PeaFZK3OmlDmklFAFpoGcxgmRJcyblNZ7T
j+Q+f4X0Bid17p08LxJ3CWjpvfSWVoYibKMy2XQnviWyf7JMzQTgWfpTta3WA2tu
kouU2LGjhT+5X9Q1cdR6m67eJWlKTyvWZlJ21UtCMxDVXuc6Q1fK58gExXCkC4lZ
C2LGk1boJYmIpS9eWHiB1Re0bchYzHY0TFeByuN5WjeWPhMG6VCjahFwgafVQ9I0
FzVkmHVtiwlzcqwpQ6epmRPjkZsBDB+93DySuGoCRdMSDpl1NCa04joWWlEB768J
XgZnUe197GBAffQieM+MLzA8kkxFQ73YD1h1abnoZnmEeed1oNt+/t7x+Ij0LgLe
ePKApwn/g+JOFLyjw5SmmfmwjhMthgt2AdQHiNK7Xb/yk9PYGmlhYxITI8j4Sh4g
du4/yT3sjLGGTPcQoWe8MWPxJ/LkNcUPos/lnFuITQYs3jft233yMCmltf551+ec
/uJlt0sSqin/KnRn3OhmxO8Ev4WZHXM3JZnm2iDV3lWu9mxOSh2iDgWRNYCuIEa9
AkSZhANVo/8O1+ndnKDI6hg7R8IRXzkHTkyCteP/sKkrbcMo3z6oIfZ24ZD790rO
l3clIu4YrDJM59h7OYTsJ3m2nmsmZLkd6rrjRHmAw3JbZ4kB8S+lGRSJpHMUJwOW
CBiauuQ1J9hoy5sTfotbfXDcP1PtsIXXj1N45kNKBa1RUO/ZSAe8WuxC3ZMFyiUs
2sFl2bdbmIGIyRcyOCg6dyjTOA0V2c6ccU3Y5AkBxRaTYVgkQmGiniQZbex9Ohwu
3JptOsu3J9LpR9FgrESxMpxa9LJNqkuJchypXS4U/0TINlrrD4jeABMXE9hAvJaG
01BH2ghcdAhzGyvxeAoZSLCv94r7eKT7fHsT3zI6h7jL0r/VnIfDOdpeEaTHM4y8
bhEVgBJRato80kqkgjQnJPSznQP3rCs7Sk7K5vlJFSuHImr9gT9CxhtAjt8inEAU
7NZFprM9Ncb5FXfeWtUX+yEcWTbpDJJjwSsq/2OsYNTUTUK2s4jZtprcewnCW39g
lRwvakKBUK2Xkjh2czeGfWEAfYPbc3N7uBl1Y9B8+sBRmNqnzhFnOraCz57EM4dj
MT1iUHjBlgWU53IEClAldiuynp2NCLnSoVXCVgVuiAVshDj8uQ3NffbXgcp9PtPd
XNuDaNbZNwLkiPfJolP9MsLDmQd7xen14Q7/Ides+q+19roVOQx5Y53G5T24MKLG
REo/tKv3C40u+icDWoltsuKQL9wH9TsSRxRHafkuAgdE+bVWLjF96wm+uBWqaiXw
QhitZkVTjLl9TIj8KpQbW7VudAuSKeKe3+14trAUjXnN5F3ugYyPET43gKEdO4u2
GhP3/1rPhOGtc5VfglgLTPKlp3u3sg5Lp9ShvFRpWDpcJsmdMs4bpJQNfSQMGRxq
a/bhithCRBeN+0vJAZs25pR1OmdOc4FcF0EKt2dV4Xmn+LI3xlLgHrFV3hwsxJql
UV0/Ak6wYN4iLev3PU/taxmtPU1A4mb7qr7NKBPqjCbFICt+1We8ZRzSUci+/I6y
mm1u9AUhlqZPecQyHYrvIjeC3+qNgTBD5RkI9LcXk9I=
`protect END_PROTECTED
