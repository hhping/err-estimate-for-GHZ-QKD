`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGdDZ7l5leh0dTGZlDhab15oSPkYjbfkJwUWMqpY1M5fnOUiZGgXsfqXMVsIj9eh
BGU/KaMHNhtD++qDreuBXuvYG7WR1DJe4AwnQkaIQxQBtFPG0FjHP9/DPzbEwi2R
745ufSPnFsRVU9DFytDvfXBaXqtierjzaU4tD4/1F3ummdeeDElclHodLyoaKnVF
hA+Y8M4NJsnsiaGbiJuhNYXwd68GEC3kSVpO2truNq5ZUGtpDK9SsoOllHyvsgXV
KHwPat5vTzQ3deSumVMp5uR7Q3v4HZItlGZ7MZqbDrrYALZWlyfkni9Cspzc655w
xn7Wv7P0PhPI7ruND7N88O1EO0bhRsEI1GOaw7zcq0G/e/uKuCe5m3MBNvX0cpRT
vQtMaHBTGKVdMyhV8+3kAL+G++/pmzkr7EXV2XkCyB1h2sIMBoCaFuvF51I7Shym
lw/4LWyXsziw9fx4XzzFrOT8Pl6BkEyj1Jz6J4pw/6XW/3z7YtNr6qJne3K9iUqY
Gu9a6y7woSIksJidxzX9iQVtCx5GtuXmcfXMnm339NP0xuKo9/P+BJj3EXLuqQgQ
GnsW8ODIhulqsv4MI4/FhaWfZrB7pPhWuVv4QkfWobOQqITCxkvA/RiXtL5UB8VJ
FrCNylK2KdTcOPybMzWhh7jgvYPVYWTsO4aQmmmi9PzPKx+mYlQ4YHKUZkY17Vsp
I0xAZvK4vSYgmU1J5XpUnrWilPSmCTz5tBZPA5A1kOE60CnHSPeEkT1W2OKxR9Qh
bZQPa7A/UnZ+73d2PsRewu6S7Hd1Loj1Hlil1DsDpMD910WsXjetZVZYW8ckihvW
LGCh+wDS5zSmNSJKx8W7H/t+zMjMUIV3E04eK9IV33bJ+dLwl2YXfER7aDJhMgr3
v/CD14Eb+cZIPu5pnRH17wnFaJOwltEocUWvFGTv/Iw=
`protect END_PROTECTED
