`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+CO5yV9pArcczsj1q3KMx+RDTRyMh0F10L1GfGVkGFt4DgNlhf5VpcAJWhxJUav
cniH6a8lxr7U5V71Nh1QEYb+Yqg319/GVUoRwQdOjYa9dkO8PDONuP9A6rHf3Vmp
SNLKUqQXBbG6o3mGs43yYOHNoWC9R+nr8YnaLUmIzWz9bzCjh3pMulBBexSpEVfS
7Pr9IgGGEmmSsWi5QKccWu6Wioc520ifr5XWS3HgQyKsO88GwjlzeoVigbbPOSc6
OVm4X2zwdjyQi7ZdYdE/ALBGMPnNB4j3xfjM5oGlteoi+aKAqa8687izme8gbJ/t
nJ4uTXYQ934BixQpxI3yIwP3plz8WVxgHgfH1NqanGkpjBzGGNBxj0YKTKR87xuF
poGxRf8potAP+/3+sG6GamWijo/nwdQC20umxuk1CnbMJ3KX8lW9qQjTJjpdYsZX
qADCutu5Mud7ugUJ76jT2k191XTbuoDWosrVjNvK5lv20aRpYT53H38xVVg4n4dd
QRjwm/eianQ+V9ARWRzycsPGCi+YTjkfEqYrFecg1MXUCjEZ6J5JSvtWoFjHLT5X
faQBSB2uX/PJjBwiwx6q2dDe0Fi4tL9nhTiKsSDE/heqGLofE8isCLewkzjG1Fgc
MRX8RL1rOObYZxU5HuUG0fTfParaKKZYsmbsBDk++DpVV2CdzlsItCA5Y5IDS7Ad
r52syQ2yDPHr53mDGff0HQuiGPSMg4cRGH87u2gKF2/CESDvx/XLZM6iQoktpt9I
3yrS9Fkq3/OeTDbD9ffWFXYPDFQjk44Sl2KX/XKRGRS8353wcBiwIS3dmN1+gMYa
kelg/Y3/PIP/T+/cMf3snJx2NmZVpUkoNGhi81uIZFl4EqwUr/6sS9byBaql07WT
dsjdpHCCzJcieTUtDXv6NAyb4BcZzi58FLLtphfC1nzy/6TSYyQ8mgx6+T75t1xZ
qSK3Z1i7bo+4q9k1M8ooWzDu59K/0VX5D/tQk2T8FQyaR6PlC30jIXYYpxrIYYtU
dizMjVGU0w5v3a354EDgzBL1l6qQkVcChVYSAPqx3KSPu0acByk9kDOWLGNWVc2J
Y35vH4EsKtaXlSBZ3fjz2pchegvsxwTKjenecu9QNoF1fZwsjeWagwle+SIaBnYR
jkCQgq/qSjXiFa6VUgISNwTRhiOAg4saR/F0vQE6P9wx0vhXe5y9m2iBGDnShzcz
BnC0k3JT8Hw8R488EZrGGJnHD8zt+gfkeC5ZC5hAl+49iVTE9mdWmE/wBErhz/kr
1+1ANwaw5jep5lXbJJKijBSLWCfeV8ulqjX7Ats/qZOmYZIZqG431Eaze3T9F0he
yMTPFY7UxJsIeslYKO6jXYOZ8iJIBJ5+/PYjhkTiQnbFhCw9ja3jnY06VyAkcdg2
2BLnoqihpOwfsYcgSB6CJwmQEyoWaid0/fbpHnxcsEfgXwq/crkQDyO2GWqKehN5
wgS4a8ekdBVnsN35MJmiSAGpUiEPpJED223GB+gMvQTUP6OGnKBLkN4ExtgpU0EE
6jTJ8B3K6wX1pAqCBP1GVXLg9ItbOUh7IOai8jMSBeIzywFRsowYxu2IikVr0ESN
gWfk7dlorz9XNqKIFNjjGrbxSkmRiDHyqQx2b+Yyq8WKG8HCZq6fVZUQekScXY8g
WoFQwMGKHbGP3JAc99RLfvekl7o1ncRCP8XTwlswztdI3byXQrSxd5gP9eJwTNiy
S1vDASuUt2jErLVre9QqtskYQskjl4/6/p0odIir9/rflcNB5LqW+tufKX3NWzSV
1dxKiWg5EuKW7MuPK0TLpB3bMSa8Xg1mHu1lwrvxTah2ExXOpbIyCVAoM3l2Bi6G
UGgEz0qhyKsfs5ft2aZo/ENM9MfH8R6gOK/uz932M4aVgijPFtHxt2AL+P3+MJHW
t1rawO5pmH3qls8un30ZgSKp+LJ/57/BSlxtdNFltieRDdENM8ZygwVIJwaGoiSu
XHTRX+RgKskNVvqA5c0LcO6FpXJeLmt4zcoaw4WvdMsThoef50QAbwKxpP4JHHs7
vrFh6kCBhX+/EnYU3gcCDEhd7KDIZZRu48RtC1kQcUuYioCr8NK/RftLFscYORfE
j9UhOfsysyJmcIwlQQkbEB1cstB3xsrbmTd7huZpDa0V4uUDZsmTKUFSHUuf8C9z
Lt4TfYzvhFOelHlzOzmLQLYC5qfr3VFEa06WyF5sz+AoqLEtp1UBXS5Amg3ln+M5
9aHJQA99tKPRPpmmbJhV29QL/hvd9Lwdh1d8f9WdeAVezPZHVkv22iA76aW53XFm
yoHg6NO8Hj8dbhRSPeezY6irPjTBNMKjHy8fsipWNLNQoXDX7SMdvQ9pBfcJmk5e
8NbfBSC8ysUXv+FM8Q5l9UwnZckjlORh6N0DK9Rn9uWlhMY6OSntdZxsi/OKyMoN
aIrrbb04qkfCs2davrw+bPiTNltmBX17aIHy3/0mshbOn6KnBOPYAllWfUAigJd8
ejGwpYJ3FUQfd1EZyKvX6apqt+Le2d++xShTitY9zDpeGxgmoRpCM2S2cnBaaf5L
LZMgMJ3FI34ck8iRSzX1rAgUZwKeYcF0a3fAbgrcl5ll1nsPmyL8UYcYEh8GcG4h
A8QkDsnhg1rdFulcGjM226WhQge+/Yr9EEQtlXR0u2qOpjGrUAUpBmi30LqI228k
EH4HL4B8bmjIcK8hfjcBj0vG2bpy79HN+iNOSXpdC6z3fc2x8/3tW0HOqQftWGQr
RCHKqgmDXezRkgV7VZf3clvQDN9W2jB8Mq8vn5MO7DIVfmfTS7Xyw8vHlmgxlWNt
CZPEGjcqK1oMExpPYwGBr0fsx3O/4SCuzcU4kLwDVB+/XtV5KtXNnC98ZQSby46W
sOnL11Vr6G52Ih2t48AF+7XTDKU5tBnX/65Ai0iCUBlj73gBqeaGSLZfZd8wsRV1
g/+L5X6P1W6+oVI6XhLoWEs9hLWh9Tu3UNaKVfiNnz/QSy07yp0IfrtxqsyK0nhT
LujDKRiiHLfantiEHwEq284iPgHsHX3fC+OMdKnUFDS7c4xnepCNvs6v5RO25Dws
gDW7/EUz4AF+2s/xbE8kzZK6LcBM39avJ/D3YVg7VSakRRFb8y2OqXbFonVF8VLq
jP3CJZhQdcDiKc8go1sqLehitnR9IOIxPagAhVZ/smxUEHz1uoS70RCEJ8IoCD1W
hSpNqaoBcl85o8o2qxPJoWFnNbR82/uwq09thPIVt9Bi7vwZKS+KXV4dI+jPfHk1
Xb4Y5jMwPIUAF7+tj0ZZNjK51tZxX7gUOKg5OQNwKZauOfrRWwlBKOYrjR5YFbhX
EFXTUAnkh0axDuSZZmI7TC9uLg2+jFBP/rn5faunC/O3rEDYsTdgcZbP1x7ADXyF
dUrKK1wk8E/NaKLcZg3jL8QLMmf0PF4aLgAJOm4Fq1qhQTdHncJBncb+nGYRYBer
8fvCifT2Ey6worEdanRRKy8mttskfe4kT5yvR3kT26gppzUUay274Nj0wEkHr8CQ
PQeSyFOyiwWjT1nmzDPyRsSzzl9sBBVI85KxAutKD3iQ4hN4N46BicuHuV6tYtBB
En2+VevT9QTXFmYvLsecbTdH/FjZ5iWTSszsN1jt0zgdH4tcz6+9RO2MPUGHi72w
Fxj98Pen+tdnW0h2NcW3APAWM9MS6vjlc53AnKvjSJzrW49MvtJ0d5tFZ0SoTcYd
JOJMH+kmWms5FlJUS7X7iRIj8XBIQdCkW9JHlpbIjOVTmUUxXkuubvvN6kGYMJv1
Xo4a/jq3M8UTuHpH0L+p1ErpOUwdzmkWDRNmNgoeH6W71bzRDzIMoIdaQP8O8wGH
5+oNBDR93rzw1eXxRlyy8yXz8DO4VgX7Ge9Np3zGCDIpVFep4NM01iGSoPpcumg5
eBFanwXB41rWSDfyrUvi6T20tvU1+UmftfkoKpV4J1y8Joa/k83031zCON+sr+lM
hdREjItjC5FTG0U/fUk/w19JcGyUqN6ukQylE1RDELns5rG1puJP86RGJtQTWniM
ejAJOArJSWeK2dRZuwOtLWQGD/wo9o9oZEgWhMVMGlImjCrKv502qOWBGMbJZuND
skRrEm1IIRt4MV+zDORi+7YEJZOG5N4JU3p8JaIlLp3w+HRmQcpJYGBoKMn4iKqy
iWaYkYtP0djGPPp0KJX3cvbKYir6MwKsjO/XFz/q2lgSGSgkdPwpviCxNic2G0pH
qWZwEOnMoRYmLhxeYXRV3mUlVR+PMXfv95n6m3Kxzc9o2POhhwoBnbwyjK1e0jJC
cDu3x2r5SS5McbI49GvfaSd5hxof8GW97eQPDO6F8ExbHgrc/wovay6JoIfqAyfp
2Wyh6gcQ51liGVoyIIy8looG4a/+94SDHezEIXUbh7sWncZH0PVTypMhwcRcOCbb
9H4wbug1qjwfDxNsthCb67RHBd4bBDnf485N3vOmD7jzeXm3JzQMdRPONxG0SGTX
UaFQjIK7SdeKYPOKrBh8gcGH+GAU2+3a9S5Av0eRYHEzCAKw6yLPR7T/rHujI+bi
6wcQFzQmD7jT/JNqbunHEsRciToSWhBjDI7HzUfgDgnnZhjo5Qyte2SFcfJI4oit
hcSOt4FwGfVLZS0M6rndI3oHQxTAmGPtHMD7SyftgmisP5ml4VXcfqFegkie19pH
k4+/MvIzVstqbu81X03q3nW6KKS4BBC2NLMgGxxHxeWzZE+UdY9RSqjzxVQMSv+x
DLzKMa6kz+RPPHGVZIoBt3ZQ37XT2tRMjkjSD05vHzOwDX3WQDazijw+ItydSMhP
mx127rM0Jay6LUtkHCzzfnnePYBpEMzjl/ZEs2pQaWSBY3j892diidLbrvr3WLr4
QU9CYIzx4RW4t0fbp6AdoQWxxKrrlk4wHBNC6WAB1zHoUltNfHD4rTPi/llHkGPY
phthOrRHEjCMu3x7b+X7Ou6yBD/co25Uy6J5QegsP8KSgfHTBccp5rPIpdduiLCc
R/oyH7N2GpfOqCjIwOWUoJRcwshV+2gvU/8x65D2PaV2ElAtHHu5G2w1WeBLWnt6
UhS/tZoWjN73hL9U/p3vOCI2/tT25wVid16JBKybjgeZgwhQfT07Bu4nG6RLrWsV
/v8WFjNGYBQxQIo+OYFLdqHIs+NVeaR13styGNkD64shdES8JkKKeUw0Mc4bmbaX
tkUb+U3GBNvehuR4Q9JO/C9oOkCXmgO+MfjVNWZefT5h+6Gyv/CaOvHKBrMgM8Pt
0G6ovwt8JKqs7+sfZlS3D+GX8Fc1bqM+/2t96btZp+fJjGuww5ijKtmOhDzeg3GC
kvLUmx2Uqu4UvRNdcztwWxmONHCSO8tejml+WGSSzBJ0izMIsK9E0YWwcXF/HTcA
3zyHThycs1r90MoePaekefHIC1e5D8InEKfa/fDlOCqnH3CCsa815neXvUfq/m9v
9vMO8eY1lVBzRaEZC+rAu7GHjBhvVAkcMTVwJxJhFdD15RIAp0/2O/YdsuCHIW89
83WHj5gS3QxfVlaUfdYM3eLtvUgwymNtNG+syrAF5mfIA2J5g57ZX8AMbQXftZ4s
pY/qLxMCXi2wvHT3LZ3cP2eP28bPPazQwpcHq8IgtGHWWwtQwkQNfXOCsOWwoscd
XZca9cvfeCtoTzTr7dkGUiSHh5XQ579j0Q0jadrYEBMOlWcD2A/d6W+mZdQITk4k
PbsIeS1jIpcQMcGWbHM2JjRIgUpBHyVuQA807WO4oitXqFZvmTuoqGMdutOiGziY
xGwOKUuwDI1caPrRv4LMH7ihUgAJ8lNnr5niRU7ay0Pob8a3TA8/WopEduWyAxyv
Az57MeePed2NvyPk6WLbuWR0L738s/uEOkZL5Jx1FBNrKJX1YE7I1FmjJVGGtmpP
7vlOvXA+/ZatzxTlh1Cmfu9115LI5ed+w1KYQcUMXEQP1zi31f1ku6tM2Lo57Kdh
MsgcH4M7P5NGgwsk0kOk8pFwL//FTSCmt+Mq+HxOU3di40qOOU4lf85DGbZj3iu5
tZkQU/Htq3VKp/7oMBbRrE9TbpYN5KhlzXfL7ZV7p9qBrZ7+393VilmXHS0DBMVd
1TZn4YLGrbBZ9RX9An4aP+VTT3oHLMPa2bCWNYNJRMrtehbeC0Oi8z7NDs196gRC
LWIO8dzT5+uA+wQjlND30i6rBmD1/09OV76VEfO7lajYaQGZcn/ds78I5bvATRsv
dljYCJVyCzNy0rVWrvu25X+gzkrDg4kwUXQZibDylMZ/4hTihVVVkKnYmLRDZEw3
aYHtDlV8ppIZ9kKP2Vrw6S6gZ5ZUl83FwZN+1JuvVh3nUqBN3bhkSMR7rV3924+l
YwvJ2KH6fTQvo4PWHc+cyfmhajhzUKl6NF1jjLtR5mLpLnkGgHnJwyfg+liyTXEy
gRes+8UqpK95MWEQH5X7MhwDHbreCh00P+bpxUttmJ0DvyZmVA2q8RNAqvIZ/z3S
wNJq6T3qsCUn4wXNs2KAxeAJnzRnpEavIMfSL5eRh5nqMK3wHGdbmWJSgUPnLL4u
scGr2h7L3yXzK7kuCyp/3jaI4UERXqGjRVEuMzGvHDuEsxkY94oB9pjS5H5s3rkX
Lf1xTkirMWTgDd1yq8Enkf/cMUoDRsqHy6sSIvj9ifYrMuP7YRPvYiMH4+NsQksC
vJMkpp/hMrlGLdzSILmbLi4xSwPJow1IVg6pyIcBLH/DREzIh+yWaD80VRETfhYi
NOE5qSG/a6d6A1pP9LG7voC65j54Yp6H+Aw3Tn4YPUd+l4j+A/A7j1syr2s+IzLE
EPj0MBNAyCXccNfy4KlgbXfFx9ZYhSquhJaOL02KJkseH3e9slYxqrTELoaHAxtX
oR2pZ0OOlUit1dr+GF8jDSGvcHbNyKsbJ+AYxZ7P7dezPm1VWyMXPZdMUNEBAnfV
iwKIOCIJZXheB6tDD8GoEXxQk46AVhMtou5c/xYW4XEg4rGDCh9YUZyw3NZniFA+
iHRneRPfTWueeZnUo04jHM5PTcNdzi/nSjo1ucY+E4iz7/Ebr3W98FdKgAdApekk
0mQvvQt6Ix7yO9q9dUKKnruGnVM0Fyo+RQgsAtGznN0MtXmpWVtq/naRUSQ6GkOp
AHJP42sYTSkcyPvmRtti5z1OErpffGOjxIcM/200rJlqF10+TkC0kWzHruZZmkMd
VA+oIIv9Rsxs5JQXMfqpQs3UK79bakxSBcfhwCuHwuWJsZTuyrwtNv2QyzV1+ZmB
TXdNxmYm9Z6zUNqAKy/t7QaSBV1QmnKrd+Ah1Zz8icSetUC6HaQUQCXfzUa51GBh
JnOLGUgcdLWqBQbvrCtd6IfKajyR2z5hOAbfNbKQjIun2G2XvFtNR2/vN6rkZ1gO
4g9FwkhiHue0Rrf3bqsIRR6fbiDj0JrL7BaBbpbcvIgZhbPEqseoT/XVD2tjExC9
9nsQMwzh2dtJXAEMZSOrVmXDK/9mBkY/NPX7G4E0sWOA5jeNuJJw5hmBaQGPUcAj
JbxPtqvefooIFH6Ik/mA9cbeAUi5trnqCm90KBOoJK4EI5MOrFCasAj8UkXQok8W
Rq4yUN8Yt5+9jJrMLMxX+HF4d4pzud/VvceER3HAlD5VqmjzBab576jCM0ikeHVP
J8nc0X6d2vidWL/XDwT+h90W0LZ+pzfRJpDHdkAzIo6TNOzXWYZWlf6bXBkKIn9j
tw9YAoYuKnULP5EpYGwA/K3uUFdh2zXxLj5KgsURJ2WBlkbipgxcj2qxqWSPI21m
7eyCJ1VtXAOufNPL6EvbgOzyBb0CrX2pBsfPUmVRdlsh8aacq3q5m4QBbHaAJlc9
qE7mlCYQsxqLyQc/xrNW9ZuiqIE7HCCbbw9wLE/Pt8w71en9KpUjniJSxZ2YEKIm
WCXSi/bW5UIrnnMrRVJUUGhNaUA/2QMrstbPZJ5fhwcjlC6AzzUHE1wMmwLgWDWm
mQAZD10+o+IkvZeEWLIE2oInYgwLHyTtTfYH0yaySlP0S/25E2FvRu3HXRUg4Ae8
j5YOn1Ps+gxK+dNoDaJicDVhS3biZWRunn70ET8r7Om8+i48ftVebEF4+XGmDHqZ
vXNH1RVpwA+wnMLKl9jVp6mthjuz5LQGUlSDMzeChDMeJReI6DJDwqAZgYhI7iZr
b6cDI+qB55gQAoq4HFb+BKpXEaHwzVLr8FbkFkPGkeZFwodvEc4w9bjfeHX209lJ
/wbalBHvfNVZO3vc7ywduli5/mti5Lbvl1ljDkZOSzZr5k9dj1JB0Q+XJyCGMWl5
tYMCWNhDSaZQoeX5gGZio3EAzqnJFN0PG++zGDEQeye+kiWq5uqqTSoKBvLt9DS9
mStNhA1CB8VBsQQOr2MSAqGJRaAVInGqxEXrTmzwxSA6qsKlGW8ZTIs2imohuGE7
UZl8rfdIcncr3rL7Z4nrYIzglcYr7EOlLS2l6HfMZBbnMcHA3hK3kBstqMUVj/9c
/7M+cyEQH3XmBRTlCoyDP8hC9t145BBJtaZ9izBNzBTr8JjSqmtEhGowe92NQ7UZ
Z3cdwEOAmy0fNB0ySkAv1gtdT3AWWjDVt7EgYYEx/iaRfCJHr8izJQZZs6RUa33U
ujoY3a8sc/8Vek4rlEBpmFAuFS2+CWpijeJgEsmg5JiHQadEMGF8QIKLogOAuDIJ
Z+Lxmqg4j9KhpM6l22rL4sgEkHya44GRxxExN86fOFokQnVj6389/+e/mjANn7aO
Dq5RQbyxG1WQ1jfpkxHYrGL0LAuJnGWeZMhEBOsf6nGn6cratkKy/7oir9PbU/Tm
BXyEkzbOUrCHsCQ4aUBDfGRyEMM8w9ddZDC6/W0PGDgg8eGrjmbdxfnbpy6pFwc1
HOtb9MnsMvohd8AHfYgIUt+byAuHfOdEkFJ7uRPNdL+fjkGxxWcGtVLVBU6BewYq
OXBq39GJR8N3JUWxnt2GtXggYmo6TltordiLmVxDKBvyQCzVyNStq3+pfyuXPUas
UOciwa8x41mRKAEW5MO2NV7JS9HYCDxcRXVXksODKB5JW3e5IXL8eVubOTzVEzau
qck0S/sjJC0UMNg1RaJLgP+2b89ZAsYeRIVTHnJhgk9BdvQkSRctyhqIpbwOy+QQ
TmJIslR9nxeUHdyI6RYOgLAykCqmUZqQlBi7vunr6MkE3TusLoAHKWcWd/ZIT1UX
bDfiDiLet1vuOhply913Q/+YYVVEKj6wd5mL5LfPzGeH851cdYjgvcExRNIAHIrv
eACl1SNZlspzbsEPpFFJ0u0DF8n3N5PPj8E4w4KM+nubMM54O9iJ/L2BYgEzPcCU
HJnMUek1w5uJJStjsnlZ0HnF/OimkXlqVKYpvJa2jmRPhZyTCU9k25p0PebTJw7t
DhcnqCOWUdjTTBJR8pFdijoT2CzfGiKYMQaZdCWotxLatldN6hvPGROy2wswT4DF
xuHXwim0uMxYTDb2LiUX8QjDnUsz+jdT4p8z0nh0q92T6EgbXY0rzH2ij++0gY2Q
/wwhzAYtYImo3WMOjOTHWn2XNQ7aWlZg4zAl/hj5fN02PHQSn4JP/Y6WFuG6GzHM
8fbiVFQCpOOgxAcW8q0vALcdMxVkqUzHW1uOU+77lZGUL9DxabX2hUM+KK/jOMz3
KcOWBRdoMC9TN6oY10y0gXzdniE+Bs1Nn1ohKda+Y/6w+pCOysmOOZ7uFgzM0y/m
qvvYTzF25JtY77ngdb8tA91tkdF2jU1W+p0WiCUSroy+qBJKd2aVCpgpDwQW8K3m
CpmmVJjZiL2UF0BqgPsZ4UaUNJvDFa7a8wkIcNvggY6fSPxcXtrHkKC1XWeWyGPj
l8cmZs94DtixWVnQOEuR46n58f7bgM10lVeE3zG+Ek9vk9qfZzvjRHZHVeN96Upt
Tx/yV85tJEI8qKO7D2xfdJQdpYoCZ3rjo4MwlKJ7+0isuX3tHjft9jmWt5xt0btl
w2oEWv1VxRCR8XvQX/qcse6GbxqG2lEl2ExC63ObRKSqxOYu4b5CpvSw6NaazfwQ
y34DOJ6pnv1YOFILCZUjV61GEyviobTffHQpWAq6Vi/XkWcTzJ3ow1yPHXGPDapL
e74DmwZY68RXROZ2HpJ/8jbjvE48KKzbaAtReMSrIb7eEV8uhafg9W1Mk8mgNHA9
m2No85rVtEL281HSC835fR3ohP1f7WI7UoaUjx8rQt1Kc0DSVC8VV+K42OohiVxZ
i66hQtMR0rmZua21fA937jt0eacp4i+S7L8RaVjo+c9WMbSisFNDKdbREtxkhD94
yxnpgGxDwT+fHBPAC88ax6py/XYgmZSyedkhYZYGyJD7FQyKFU4DQf4ENy6QEJD7
lrYWCmuRfUuFG/la3wHH9DoeMvi6gXC8zSfLl6RQ4i32vFjP45O9u6v7xiGZyoZA
3KFAS7ol0d1bC8+KuQEkMKBC49Mofxg1C0KalmKpllMI7A7DFZyMcgyVv3iMZ3BE
PEjPQIaHZgI6bsJvZCG3Y35moUG6e3BcCMRjyvS02510P+CaVFrO9wj3F2hStFok
1zgTAxQ7tYzAKizO/XezrLTgG9+ZzkCkt8m8ZZUuHGlqorUbwxOLl71RVdpSnLGb
2HFjKinIktsbaMdxFYG2QgOSMVJVayFi5Q3h91XZ+5CPSmFkU41A6y53iJzelXyX
ABi3sFG6ynpp52CwzzQ0H68jAlvHJ244IWRH/hXEG+k8WgneT/rhqRr870iKQptW
LtDORuvYyfd7W4GInyJt9z3dvby6QO9lL9oKHggooz9GVqtdmPlKZaKy/ND9nzEt
JxmtWKoppCSN3jM7HO1sJykz8sNU4DdAxsWsVio4skSpcr7dZFPWyz7MQ3twwx2C
hIBOo8i4eae7MSmMgDv1MrHdYoTbBVFjWN07czlI8Ox8PXcRaV4OUexzOeCAduxG
Bye0yr2jsPvnt694qckeR6+Ok23OI/Krw12mVfynYtabGyhfVtAwGYMrykNltaAo
hzqHJBT/zwlBMD1ifk6Yx1jx2F4PBnka81wkXUND6oUy3aKM7QDzpvTvznx/RwKk
dnGwPuSGzsznKQ1BeXPGpRnq86xg5MXhFp9daqfxMMUm/v/tnT+fpF9oKhMh9wc7
c2KdxMDI6HYNDO+SJo+D2GI64xfgl1tQJQn6hKc0c4/CKX+03NOWLfUH4CsHfMe0
Re0eMz4JMRTxnRLG9JakzlSan/WkaV6ew40nddV2oUjWFyso00BejlmJeWDZOVWi
k3TRYHTR9zixIkCA4TFx9eaXuQ3PjbtBbCT5dprH4qC9AMNESq0VsRGiGiYw5YfP
oWeff5cAGnXsD6lzL0chF39o0WnY1iRMI3RLsTkp3IEtw2n1JEA1q/QBtPxhMwSj
GzRizx8e3YKFpG/23Iu39MRmPLxn+0xz5IRwxPYH1VZ4KsL1hgwRvnr9BlqsXEUD
wkJb4eOpwh5JvC/2Cx8QgvIx4VMY9Ru5wlk81tAmmpNEqfDpPaw8WF+KyOJnwBSh
4sSDVGtd+qmQ19PEOlPnVRPa9UPI4WBiwbfxpR8smmuAclvazDj/dp+9Ve5/32EI
M4rKqK2RtX3ekVSWoYOvFMJHEvCTK9vxJvk5kNQ5KiEgT26IfeMMckzNoTPGz9vi
vEPCnmDlb5FoYCfAImB6XnDXO9FrneVrqeR34oazMeoUHzpW2W0NBW6rszNmrnKu
nbTp+Yqz0n8RV+wu62t75/n48zNJnJgtvdKIIajeaLJt3G1pAo4cA/dk1sQ4C1mV
4Gz0EPtxPWXBWtmHZgZoy0yKYe+BeJXlTsAYlyfwgWVuxpcDlgFYjIWAuYGW1uSL
chVJ3bIybYWMvyTj1G6jikDLj8zT3H/5K8wlMWhprHF6fIZj0EnztcaGXJdHt1gc
Shs5FEslcT1GiO6zc4RKKd6zPRji+RqDHZPkNKqTAB7lROxEx2ezW4/tQ7kbcQQc
gZEEX2h1bt8mf5fc3gBt6NfoLkxV0ly4AfhiNWSPE+EeI89nbhAMYIzamXASeRgO
UIa+V12s8DcZ4PMxMp8+9xFKwqVeGbRALtljMkneuWeIv+lE18NT11KrF+W1e6/C
VVISiJh5cDjJ0XdQi2h9evHixg6RongOlABMkd09054zmUiDwgPyPt7BPF7lVHA/
/sLxq59oU7shoSN4n16JOwvFGEaKm4nCuhiBR+G+tCjexG9+4JYWw0TiCZdPXhX8
CTLYPXyu9r2g42BJ6T0xp90+QMkbxVC5wZcwv+R5G5/wzs+CK7uDbksWKjfiTNeF
NNr2eUmBJC+u4GuFkrcPIc24bZc971Rjz9ZJVWNh3sxQowVjWNUEKC7GwAYakS5l
tGIA/ZHz0xOTX5wTjqrgiB1lDSi376+daHbhvnmrLZtwAS1fDa88NckV6z12+9Iu
HjVXXO0xCXx8gImSHBKCzwWfqKcZ/tWH2hzv1aBgNaqotuaRsu6ChHLVSRO9/n6K
S5ju6hu7a/TAfx2e7dczbZjgsvy//8wZGShLRFtWxVPLkIQRgYi5V6CGE92fN5ue
wTBtRNlqLOfME7wnEU8gZF4RpD9ZNxPFrbREJlNMhtp7bdwu7ATFN2NlOtSH+Vjx
DKB5b7egxxFQkDExOhUE13lF+012nPr8JzBjuDeMDYPc3i5dhdE0bFzR4W9gmVQG
MWBh1wXDNzA4zxp1j3m5TZakXLSaT4kW5RQY3dcuO+mo1X2w5KvVrl1ZN3DWdL0n
BZfz6G5C4gmVlFY2xtY8icBEMs0VnFVL6F4bEHmgW4DtPGzU8zs0Y3Yacr/azBgz
foMkg9/+Y6yk25pXOWUGmTNXYaYxBgziUBOQBWArNaD5wa2bcg3JqmOF2wUsjj4N
HnGGjZvkRcA3jcog+OnIMF/StW48PTBhjuQnsLbS3nyaMvOVbXviwp5YnGg34SH4
eTwI0TZ07WBJHbK2idnzcvHs9KWYhcMyMBueIlL+ZEjQMiI5n2s92MtOvH72WkE+
6+0o2D2vtE4wDjrOdyXXT7VG1i/hKZVrdkEGN8JVcjDncVlR/DDZaKRbME7NShdd
UpkjL0zaSWEI7bLT5lXke7X8G10DJuD9gTX8+o10KtPQNQKwoMjZ4cq3NqK500JU
3e3D0kunVUjnYjR0J4nE68QIFnqiS68FoZksdKJ+x7xScDS5MOHRcB52L5hOt7N4
COKiF0Gxkzb9SMLGgZ4LP6cvCVu0jk/lmEK4vPXa+lIphJOhCw+tfy6QvArsHMeO
evY60j7sWTqlELbkroT87L9aTmy+Ib9L0ihbNPzukl4o/25x6juhOIZCGAn6f1Fk
w3b9t/W+PFb+aY6rvXi+cXexkrj2GD8A6w7OsqZ4oMFGydwV6AffYs0b1bmlPDsp
45x74pilWPea/sKyt4r4oeJmf/aPkVp6g/yid3Hw+cM9gpMzbRvzp62ZFPR4hmP9
SsFXe2mY7/pA7ltd5ZOs9AA9PbyJNm3KqYEbxgT28ayL2IjR+isJsRZaNNTVn7l1
DfzPFTBifVlDvDXDTt/C5xnQmovrXtn2tweKQREzUNBTQEvJEERqA1DOeiZO/AyQ
TLjcNxmCegSJzKbjmoIOfPxg20uSQdmP9uFkL+gPADOUmsZ7tdW5pKfA3eqJHdQV
L41Zr0sds/KyNdZ6kfjAih9SyHYKQwYAWytEKLgUCYMWgdTe/fZquv+xh4FlksAF
VNjyD0S/dlEuEkwUvqU4rXIraLC8P8+PqZKRsYuONy6QMo8T4+lc6jOTXtvnhyKQ
O4xrvB+KraJeXoFbReT9gn7rhDWv+cpLsiHaytEVsRAWxIZAfUVb1xx7x33A5s88
V4ht+CGitC9NTLxrL9dXWrw9z07RLfQvHBJBSiStiX0hGMQdCDoq2JQcGedAtttA
BAT2qDU2Cb//CA42inqJ1358qFdW48MKFd777oBFWki+Aima7M4SCCDChNn+qS9t
bGrImnDPQcwzvzreCtcKvyoIUtjozjsTSnd9bWuqOyz32MamKEU4+hcTJKq1Hjyg
5nGnCHrAtI2E5Ae3zfNxZ79tX+iurS/3mlUxGujzJsnZV6XkBlln368AHHzdgaRd
mrq77kO/QaFnAsLT1hTmHVImr/leaXvkbrNWMmjsei8ukLUhwEmBBmcNRqiwCxFS
OPhdJjaHmbNmfcNHe01hT2lHZ0xce4ZacdkoqKIfK9ZtKMb4moGczz3NQKvLHp6u
xbq9IIkZx5Rr/LmSrFUtNPl8pTcZtz2i2wRHZhHnGXaXjsFq9a28XrCWOkNZ0tVO
FzZZ3LH6CAeimq8sbP7re7x5/qjTlV73vWzCMrgw/Z1sR+6yjJf4y3h/26BG1P/D
7MH2BBR6T34zUAhKAjDtzcOEv4WPTQe/tNEvr1mEME197ryHEwSL9iepEZjGZ2EM
1w+/6f9FuLU+VOxg8P43jICYN4xptVMu/UteqnBeSS2b2GLDOmvpQchvod5jETbG
+mskt6RUW/yz7L5b1PITPZAIwxDHyyVJheDh0CwUYsao/A9IIMjBtVUs4/MwUf1W
hiVqwHrQrxeVmNRL1txyDeFMKcLgsofYWr4ZwW5/wNaubIvks6snFQPUGgT3owvA
cNeBLw8BXDNJsukxrSbHyLfTrgfFGJ+yb6lFDmKdBj4TkLzykNlvBKGRCeqRO1/A
umASVME8Ek9AAPcBWBwNJuYwRtutxVE+7BYPP3wDcUAtVg33R9xh79KHX8BqsIPF
Yy/qyldN8fPjimcrIwwRkryZPtIef/Nlc+1p2lbC4cwMI2o4bBl9yvFGoajjA7hv
v5dE2cpx3bo5J1MnsMpSkft35DDIZ0HHkYavGOr1JoZ6qewur/V7SW/JMlKjUTZV
oKIOdwQo3yDkPz0XRHCVovlRIOW2jnTwT0E/z0hXqh6zU6ar8ULmsgJnHu6aZqPu
JSguuWjXbHZfeUtUNzFtGBQMRSK8HI96+Ar+KcdQSxgr8kBwcnSaqSOVE6rHNPan
JPNHPfgDz/bKZiVjHEqfCV7GS76+Mn8F/1T0/sXijoK4usZQHqGXE3MzlX54u4Du
WuxkqOLrp+xxeyIAkZgIENPLkPME+j/RL5llZI+o/CHznF4Iz6VgzKgfEYY+Kzwg
HzhPuyIA0k0Whs0WEVGwIi9kltkkvu6hKQQuRuD+CUFCKor58687fNKBYdIg44Pd
b+Wqf0s9pUJMYWJzIeo0Mlo5+7VS+vXXuXjEDJaFqyv1eNbX6XHWXTdYvKZ6cTnE
lnxCxGloGwbTWAyGND/XWE+3HQr+suq+dC19mB2KKBDQjNppBeJ1ZDnfH9lv0f8p
/NWPigxWj7y/6BEXwkoxMWYMHaVCX2yDZDv/2CbE73YQfoP+tV6XRIaaANlGc0XM
ix2wSeL/3aZkPa6lGROWTRlJhgzVlrw2THz2Rw7jbRXFyXs71QjnORtWTCP24D3r
cblrufyxqt2l5qRJ5ppKVDLvJJjcYXn4qiecE1RxPCVxs5GCMsWyzCfXLdYsnPOl
aRK0qatXCSEtnaxZ/uPLs1c51T/iLEGhmk0iEkIvxUSCwU4EmSFmR5PA1LeQgVeb
CY0ePfZoRfupU111WFLrQXTWSQCh15c1LlDHqK/fO1iFCzpcLRMncxfsYk1FIqTl
IQlRhAbZbnDKxuRQ63jq4+Hrt3hXl4dqxhIQNwPsDCbA5JCEUbsd6XoVqoX48e0K
FixVMFIcgWZnJjuktAbN114g4OTBYfT3d2RMTHHORBxW8R17cZvyL+PKIl/MBI2r
Dsw5i/x1HnVQb+vBA6dcJm83U/LbJKUqKSGTIy6tSyhtlTs7vgLws6FmKxLdxMBf
o0DwbNQFlKCDy/EeKHYUjADciBRj89U81TxicahGOjvcm9pP2K8kF2nr2i4sxnZB
nJxy2ZTpYChSLd/f4e2OU4SE5vCx2rSz3xsnfU5+b3gHGcyYa8LoO0FWvV9ZHrEK
+12a8PnQ+pfNU1IKVTi1QcashUJPsIfH10pZLQFwxMUNbGmD2YbLqGJJm7+fRbZ5
CPWeEB+uTw+/jhaQDdCxCWaDnm8dvObrG0I/L6xP1gyEbbkbYLP5AA/sX2ZpmOPC
2v+tAsyf+pYIzz+5AwnVZjRRgpTkVBw8JxXpQGgSM4CA3XP9YvDCgIvXuSozwhmw
k0VyjyeoVQru4ftPhrKwtKyt5DWvTryzvxieGWB0UflIUolDosfDT5abdNLJyote
PKQJEGWaQ+zU+UJgjy/HBuqkChcq7c6rAYkbXEiDsEwHeovAVZad3pYArZJJ2Hj0
DA08oSg2ZiR80iqlpsyISiwZjzJywZgp6QcGD28UdbPurc9ikdamDgmB+wxLqZfo
NYVmEn98klEXGPdhw+ssL0vjR20cgHvj/A8ZzdSlv88MAkxv7WTXInQav2HV31bY
rAaY/AaJuhhUK1Uc0rtz7iUGAtidk4DCnuE4PzPWnwT7UzdrSOMa3ZHxt/lTWr/P
NVu0MrV3RRI7JeJNPhjs+EOC5XQxzJqc4FbRJbTTZ9vd/ClJ28DrKBQBXroP/5By
1BIuDFUXU06iSobQ1LEjM8Qz5zeKwrHgujcv8JEgLsYwFmB0l5A3Ll6IxmN4LZPT
WG7+J+yMUp9jepTZepHJe2IDFKIEfyafniw+px4rTkPbQehaUyGKtcQTEgbxq8Ym
IbkJ1YxV9SQpWZ7VTgYTUws03ChQKk4QHf9IPcZNCbmVeVai6rmgx18mrHZ7NNj9
k/Tq8s+Cq35lXZTx+boo7ZktZ7QQNwNrk4bT4l0LHRHVr10WZNoJeJRihio4gHV3
USUfzt/vO0ROL2eVQdDunzD3FEY2/glBIk9kGCYWR3iUG6ZyFSHpzkm20Z+084NY
Wsqdp2QCntG94klPQpgqb42jw2T3MHQg//0zbu0bhc7a3Ag8E7tFB5QXTzTlZruZ
opBXxU20kSdgzi+EZ3Hs4QPWxBys9xpYdPtYa/MH6A0ib81SyjUhFbnfOfECkL9z
d3TRjhTU2izjHy+Ms33qHY7xXVpV4vuPsJFyu6/nKxmouUw6VFzTGgXi9OuYR48A
xXOXcbqiSIoZFzibjiJRTmRwUNdq864fveRq2BPnBAGIEfDzraKXk7oWZHu+RIN9
0UaKwWRUq946eO3nHY5zt6l/ZB6rsU3or1KzWc3P7tW8/leyBp9LSOwRKNOe7WOs
SUHudBRLav5R9mmqiXihkg==
`protect END_PROTECTED
