`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWtgqxFLzciOOOLtZ+aUevVwzVBCAMNvJCpWl61LyYaadO2Ifvw0jyCqezLUG6tE
MBcUdyL8FbVglciXOd84ymDN7ysIdkN8Ra6M+mSMtISlpM2ljgLqys3WYfGDTEfZ
R8HDFLGCMXQ/rm36bSfImRz+nlp9U6OHagqQ4DA7YXGXWD5PGqmTQw8Yb11VypqD
XRgiYSejkmRR8WIqu1qlAOWTgkGklxpI/60KSSHchitUeIOasHbozWKsM9MnksVB
sZD1BuGGKQEAHiQYnsOsf/bBHqgRVLhZP+fn5epaqnUL36lfDValehrUUBfMmCVD
tMU4KNNON7H9XE8igChKR2ejmGmMFlG2c6V09JLQnQWHzKCogxIvSLI0DoLqb524
hvALukKvzkZE4VheKeyPg3SjzXaDkVDeXc3vtR8Och8J7k4qdxajRvAZnUiV9UbY
t77DZadDbFN+XNYJP7zLF+mFlXwiwqn3Kr2KZxGzVTgN/n9RtP1aPksFD5/yacWK
gJuQEgI5pMWeCX7zX5aM6+AIwjMOQ1zVLeWJJtT/297SkHnoBq6067GYZtB0qU1J
EJlgJVB9eJTuG/AT8IZcdA4A0idW57UwoAPuLnpWBFzeNej9fcj+2WNDjBn/hSNb
4UGAJKm0YPqeM2HUX9nzGW+ves2zaEi/3opjpcnL14FxnsA8KcVAHY3qBpiL2tbN
wrMK1h81M8uJ6Y8y74WpmYy4CS7ywmdocvVxthbctgYtyYI3vTJ9L7MK77+CnUD7
lTm7e/zBK9SIcpGr46jtwOocvPFDDXrc6MaqLYTxOuvfOPx8M3Yvk6R6NAM3lKw8
2JkDh8ZF6k8t5lZVzTx9EsHWfx39jyQLaeJsVY4l7rXQihgS1e9aIDAxfjdPYhKt
hT7rZO6HGtastg7zuHf70reHLAwcQ5ToLeCShBepQWPo0+XksLkNsiAimgDqM2nA
6x3NRjdoGsz3QrGG6ihQMnzq1F8XWyfxn6cAFY19p0s=
`protect END_PROTECTED
