`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1gv6Gpwn4nzfbRIIGdV8CuVYKSJzg8rBoviy7+js2leu+aZrn0F+ngXnmABcB2v
jQict2L3JKoUkw/qn6fvrfQDUs46tMozu7nUCHcgd4gCgPxJgK2Af1e/SN5N1/YA
AymfDJINQlQcpQnluKc7Tbced2osiEDfntXS99RP9e4dHaFVdUbkST4+zP4m9Qx5
50QeSrIPEWS1xB8nQ8DQJht4YKgcHLHk7jDOf/yhZ8FcCMUcdAu3+5+01yWz3LNm
jT1arNqEV406pBjpSO/k1bccAtQide1JvPtuaVrid5JnhAVhCd2NQkHhe1bqmLEY
+sKvtHGrGc67p+sX1V6ijj2ktK1lV293p4e9XLyOb5vDu2YkkS86qS30eQ1vOWfe
i7ptPePV31uQViRT8Y/QWkq7eYzu374umSyqEIKiLXc6cnsDH46jDUOlQ6Bh+eKX
BfFufYGkq39eA1ryJKV9ovNbIdRIJLoLLLXJVtkWSGU7lwpzLv+yMDKlZrtVPKVQ
HO0h8f9zhw4OHCGWUBUsKNqygZV9eHq55hUA5dFZBnVWw+u7MIhqq2VY1VLiPyR0
jakH9sg/jaRFo0iuL5ANu/rjTLbPU9jiFPwoR2efzqwxPr2tqCywcoXG5uK2rT32
hHqrScl+BhheMQvMHLzQorrqwYYBmrEwfuhUQNtHi+Dsq94JDcTXsVxBL9UYj12I
emiJMGidGg1u4HASS1HX8mvybktl4oqhptd+rkUxzWY=
`protect END_PROTECTED
