`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EhJM5eZcGZWSBVto6NUBycXchSySxA2YtvwAJaGrIgf6ycaJtNQs2nMloTyWpqSA
8C68YhHCJETC5iXAAUJxKOeREUuldeRZOdkClZzgoOAawqgzrKCmGZcha8WKxM9H
0XQTJRXdeyq1RbKOY3fDDuueLvJdi9+/FqJhllKYg4hkd1dxPXLGRIU+wVzbYHo/
nHK+8D9MD7lhjVnqQc7qZd0pp2nbas27UCyaUYDDybzm0S7Go/N04B1uZeh3XkCJ
rcxj2rYqBLtkROWid9fg2Tg29ZT5Vydd1IXsGAKU4eW7YpEFsx7I/1cMIrLYVOHq
6zCnCgoKD50J247HBT93RHOdHG1ORQH4k44OJ7rNc2yZl3bz6EeLtUa0GmR8dzCq
dBdlq751IkYxjIh0TazkHHHhtTnWlBjJIVXy1SeAigYXqnDjftNT+n4FsT5VDwnE
ke3rhUqJRMvO6Qly0+1meRuwPWagv+WY4NzmwaAGCmt94cc/nXWPBHW9sz6BT9X4
UPJkqprnOW/Ho6IQADWEuc2oQ6euRyrpGr3bnkT4OnC2107xRLUF3wl+zkq1FJ5r
0fG+Kt7XijiO19Xor0zUXn9bdnmypyw2tw7DQUYOj5CPaj42545iEzBOoFgvqUoB
IsTV44eOvoNgpzmKiJStHZe80YhfcEF25NBkxOHZN2k7ZWZS9nHAJVi9QyEYEwQT
H1GxbGZ0MsyNb1tzO+TrCIXKE/1hDqZnWoAblODllw47z9FRcAcgx+Vf7Dp4CSE0
TlYHZoQe0S1FkM8sdcjAzwUhVP9QMRM0fzIcB+ZbfKU++PGDFU/b+Ap5wcbPV7Ww
KRjKwLyNJiojKXJv3TFbBvtSYVN3Z7+/4o1HYA/UGY9E7ZPLK27fvm71V/Z1U270
DtvGNAWDYFa9s62cPZ8WI0wmRomMdByoKZzNUZgQKA9SFuHURsdKlBLqjcanpOdr
UgxqGSPxPBFXw9VZSDlr+yAhqzaXwdLJIS3LUKPKO7yXdUeSZs4YgEKg6+OwozOm
C4lRzuqUfmbrX0kTUT09Ri+3s6krX88C8Kps4tnEmreN6DtgB/bvwryx+JUQPUg2
`protect END_PROTECTED
