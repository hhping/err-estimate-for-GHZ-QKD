`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVCBULZXRo3n03MrMk6MPPgqgplRgc9VEzdOcbkbfe3Y8NyEXULMU7RtRdfl2X7T
JXUhCWEry3/xOsVUwkW0cpxeqWnIMVv9csavOrTw87wFqOpWVbYTE/aXretl49Ip
m7ft29x9VIU0+ySS/1yNNvP7zgs4M+aesvv9A2/1HhucTylNh/Khcbt5U856ghP2
6oF6PNTteFURIJEAHKZyuZ9ObhD2VxA6Hww12b9OkaBAWfLqt6n+ivYjD2uw4wZQ
EelLzb9hSepi8RFE+umx1zFVw34FBWwkjmyXeXx8d7VnUQziOZPKZQ5vX5QfJySB
44LfJtEC6Ol85yAsD/3wjQyPU8iTIJZW+dnBcNLJLrVPsGQubJRvQia8vWoS08p2
Nl4WUU+vimAyAkYsDHH7aJy7OZeFwHTdRXOUmvhBaXVF8/KmyalRAuEpMN2ItESu
4FrDpAQ4mE0mGI44l2kC3GcOBE2A7uNOdYrEr1l1K3tsJCUQA34FpiAWnuERfKDH
YH9+WPjNTTRY7TT3ye17cTXhgHIhd/mFyZEhcKwe0yjb9a0vf4Ot4P3Ov8WWRcvP
fu6isK8tM5kTNDrMbR9bvZLnHnac5M1VrVLcE1LQjR1NqsZL5mMMZdFX4GMJ1faF
aTulteZMsPjumL+3wQEdWzGrESn9cAF0yvcwEftdw4HHZZ/wfko9/k4AD7zV/E2M
81LiiphL+/zxdYWPhMp1de0fmXk9O1fRvd2w3QAW8y1P59AAWVY0Qd/EIVveJr2V
3VXfPwU3oCgtw5MBsgITXUdbXayI2iRhA9vI1cfcL+E=
`protect END_PROTECTED
