`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mjYb0/WcEO/GtzUqXB5nvnswDavqaFWMmLxnrQTLmD9jYQ3Gafn8LGU4bK7kfFP
jZUdwGQnTdQZXajuxT7BXxDtJJTuOADXuvYmod5Du2xzvGnWW60a0eccz8HIoKvZ
LvHrv0f7FgUdg9gDWPTfV3n4AfQKnYsnevsSnci6zMEg70iqU2YQTua43fYGH45L
GtgE98JoIuB7j8homhOpqDl98NZW4V5uUxetuaThAlYX0d03zhpfkKTy+oiOdZt9
jKMRMVeAwgEyabyZvwaky3O9FxHYd7rG37WS4+lGJppIWRWSlDFvrM01cHrVmFVV
Xed/k6rpnMKw+lUwe8ijt/lMkgpJR2vLRKuiprh9H+2CZOQQk4LEqX3bU/E4U2Sf
ZUq2j2VvhhaCCWbhbGRkYSrq7+llFqJZtnloXeXRSAbtZoZm8LQUn+K44uFTUTyg
fPr9JVQpakTUIce4LbCoQbwU3n/sbAwiGz6qv4SI8IXFIujVsaSAhy1fla3p2krS
AcCKYozfgLi+3oW3HFRyDswwpu8qpfFyGwQAl9Aq07gucxWcbN9cpIix9acoJU71
x9WXQfuZcKIQs7tTBmILK8qBCN4jUvv/wjhs7PTCltx0o2q5HGuOSA/9J9+ODgoO
OPRwjyb+y7tYAqW+DL1URQvgYaRr8pqcIZaYJHh0V9i5B6UuXxuY/B5IZqbewkHo
jOlran8b7U43lNgvJ4P7J4fXLiTEtM7QfltbeiAO7Wso54FkHN6hzkCV9ph4tcuc
SYDJAtE/QHW6EddBvOn46/6PrpGR/1FD5GECCDKGG4ugHP9AF+b9ALFygHh8WKQ+
7HlDqTfdOBWD8QoPXoH9rtF9KFZGfOTE0HSwPYb2M06yQZZni3dH0/zKV9ucTZOS
2/52GYEc+edycYTshUMgv0a4RwCjWBHtt5b4nn5l5V6KTymi/IuqAfaWK7uPNO/Z
KguC2j0o8s106nUcq5hYefPwuSIBqnw7USNGUJIptOXgnBbQbwkdnLLvkM/BZ1lN
zbT15D1a2FIH95EXBfZ9a02tGqSW8SjSzqwfFETPSTfHZ2lp+5CQcZPApWrcinq7
G/4Sy7+oWn8HupVHxf9YZ/zgC0+9jDm3cwquxbIPeL+yGgT1Jmwe/lKaxwnV/Sri
Aid6Rv+AnbunRmcePreWEnX95QHPhqw9g5hxpfeH0MKwcKuIcez2Iu0WK1y40yiW
/D1LjQbrTzNVckUjvzCRH/H+ZYg3Rl45TT04of8YuaIhjTMt+rTGzOpKrhHyhhh1
Txj8etI1XNh890hwLz8X2JdoFv3SOsK001hERwMVQ8m8MDibB+Jdl/iUejcura71
SjYeYBnAn/rr2J/LmKR6gAbjKSSiHZbtH/z99hxXYdgonIR/BxPtVatz/oDJ8AEN
8STDZBKuDD6YxJNk50LAR3VObiGqDslqEFfo3HaCuYoHwzidKIFuloxgNtub2eJo
dU7p9bZV+QA8cnm8AHOE/M03e9H/1TjMuOYCBCQuE2fgu8kTVqMaIupMDo61uuUd
6x3/Ex+T98iSMyqfHwsPIwSAMHvSopjGGZlGVCz+0E6GlSq9FLzJqY4epzKjgVr/
DdeaPk2gy34IQ5W0ZFjBVS7sXA0q3+GfHipkMfYUAFFNp0i+x5b/a3e68HbrRQ/e
nMoH1rTQVysAE1pVVkDLCp1aWk93X7cJUwR2yrI/LJic49va0GV/QhRUCDBVpJHD
1n4ykS6luod8ey26v8dDhtxa2BTsHyVd3h4DVGqtCSdl+pwjb/GZplnxGjuRJzG2
se4S7ceXOls5Y3sltPpySe5AEgr+Ur70ilSnb/pzZvYEHDZr2fEDh9ZkDVOb5x8r
8vbQ8kAUh8pk2c+JkVwI/4VLDFa7ugLu1WRF44/epCQjMrbOCBQgFDd9TTJNOuDg
3yua3gMqFyYBygHXcp3U7PdUNN+bPzO6jD9fyJXkh7StXwLrpI9AfjQQ/WWF3WRw
/0LTcX57RJE4ly39J6nV5sHXbF0snwXh3aBzltE8K4SEj3xgLjSCPOs1aHrDe4zO
S7OjUncWdbD8iBl7Eti1RR5UNmWMyUxHw70sxw/XUwuM64kZXGGcx4V2lzCHqnPb
TpoL9PWhpe6ptokdw87QlJK5p1SyGaA3D80Al9/fpEzDXX/ZweCHUJj5mgTx8CxD
lA1h1BbLgWdNxTHpYccW5UnMW6ol5vcOIO9KpQY+CoJ8qQ8TXogLGblh8yy7+f0+
r7/+27JzMxdSI1MwyRjDVjoTkQCMdapwI//AIi3W/f+x2vH0fzWDH560KBUVGW7K
9XTN1i+T1H/UTk9Ria6Dxt74LiZXpq4vTkipf/jDwyyhXoxOltfSAVkFZ5y9eTlS
uOvagWjEL4+lIKnk8RJmym6N8wbIxnT8yVGfzB787N7CoBRpY5WHNkH8LqGHL4db
jlpYltxsntkrRh2HZuDZnnd3xxkJvJ4mSn7XYbo6ISz02oVp2P4gPuDpq7oTdh4b
pgV9vDgryqA9BD7fT3lZ8qj4wGm5Pixwun++ukwpqINShIkKlxbc9ya7S2xokVcl
KWbRZMQ0SxpHZwSq0fUxNhoEGP5dCIX9uYksTgIcSvPRXWNnzsCy3n4nvk+8nVeR
WXUv4bcaSKo4nLM2f2J4zSxaDMhJUsRONJ6vDEq3qQ1JqnHYiwkosO3sVhgthFRQ
YaNp+t+Q7hSVyRC70gj1BzSeK93Z/R2eSAFgFJ/ZWgPQvJlova4a0Sh2rMVzIEj/
Gb2ZyziR40j11Nj3CkKFx/aTwcYzLOBUV49FCXpyRMIfnZjQZjdZXFwFlRmNJW2/
ZT7gPHl8LADIMl3BVrH6O+j+uGq/HJ+y4S0ctS3L9Gisp4FPLkqmTFJ4mQEkGt52
ZFEJFHHQbESJ1vFEmEUPhsSyo9Y/dHBS06N2qjfRzHgb+XD8DYTPd/xIaVQ9yKr3
cyxwiHaf3UNINgIJbI87f7scjdu3+blboDg4SE3wd4EBBzst/CRr+ZDsuoUwPpGA
WPS3d0RLaoMUa/SMTdSr5kQGBzjSvNz9Wjmp6hbRkPkVgcs50+8uDuHmds2Bjh2E
lnVh0VXVoMNCTEVG8JIMDalg5clFPVLo/tPRGG2K8nB+pN58XJPDEyD/QjIrC4ga
AP5PXzJzpDgY1TIgumCfmMPnokj122IMJ/fdYe1Us4jLrmMuKnKQyqyxzciJAVig
oBrF42IHTlw/LbjVS3KZwX46gARwniL6O/qmIWznZWWgHnI4gmBTcH6e3bANqmEc
h0pN/oYjDowp06i5muhqsdFmzCRwKuwBDU0eYSaKWhQeqbZ19YXq6ZZIEKsHt+B2
oqBMTZ9FTqkppad49cLsYw==
`protect END_PROTECTED
