`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9hcuaM9Xu+lrdhuAtCtcoYoN5LQedCZ4N879aIcr0PkCbHusuF0JsKD44FsK9k2G
E7pdkalLgWqHLQW5ETpm1jmUIWF90HdIcujlh0uzq4aKbEifhxVlC5VSaMItTX14
MpJK51XooCfUEqBD2/Hmf2Z3ETwrYKwF94iD+xpgcAncTBQ6yYltp7ORLyNijtm9
wZD0NxZFdEPjBSIanOTbCKPPUZdqeQZKj4jB2xehfDd/510b3XKRInDlQw2teIA8
Sw24EFu1vwq07aJnP+zeqF4ISrfw3KO4eYsWZflhmNqsTFnXOWsmXokPdy2rdynh
KXGOlYbEzNL2UW3B+q5muaq5UJCZkrPyscwHuWNHO90VqKQjkHbBlEp+9bbmSa/z
8WO0rYO9Pn5F6bMy7ynIi31uWkmX5sjd24N2GYzcYUdDm2zdYE0uNnf5EyUoSi1H
278Zqv65OYwRC5OfngbmYPPYKLKgjUmrtHhTbIKQ8e/ABhCqqbMe5+vr1xwcN6Sb
Fn/btmnMU3MeY0+OL99ImzWqG7utbCyex7Hc+SiUpAg=
`protect END_PROTECTED
