`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6d3Z6tmo4suQ3l/79VP4n+yQ5jfk49h0FINERwB8FcaRVspBAOiO3kEwyG14fFvw
qg2z1q862vyrKifCABHl4FqPx3Ogmf4KDp87slG0lnhgQJV/dSw7INjL6FfGxaZ8
iqSPjQ6uBw6mppDwXLtbxmzGzOyXIP6JgeUsnDiuTXFilH20+jJH7RxFHmXkkAb9
AUkoJ+dV9fMiTYJ7sN79tf0swDocG4MawB2Dz94liGI+51/1yQ+EIPn0DKfrb16d
n4uPryQXHgQ9Y8dW4kWjqORB1VEGyzqDJsQcnCSx4FiTNS1h0Cp6ferHfw4OUzdA
d5U2S3ShDpAM81pSuqVbY0eqVbGNBHqIv++2v59f5sGUCnCtwtbxIMQrsMkg7sKF
RqDkyRyCR1dXy3ENE+J/xE0RMzwqUAa3oMiiC5RBfaxpzCTw7PYNOSm0raAb/5pV
Q9yLANwXSjDkL5rr8HrWnhKWd7yXe0FLDWPIuKiQZCHN5g72yDeytPzkSwLGWoPT
1tnNU6B0vLZlg8p2z4F+nz0RGLF4uakhSWQwAwrYQ9j632QJF8WC0CklmkIGgZvR
lQQStnwJbvCre9sEVq8XneD9iOZ7QFC7cIxXFiDyU+PrYdiL9PK35Z2MtoHMUaLP
QFCxyk4rBkraKDSw8V8H37/xluPmcX9nRIZeahI3HJYbKwm3IaNRohosKhfF33xt
BExea7QwZK8D0MoEuh6gLzX5jI/NQ4eLwyUeFoMxyWZ+h1v9hAzJL5W/rcK8RDW7
9R63dvMIqAXuVnYe5rfnLh7qPwSL1XiemSjVDVxwS3zOtW9AIXF9RM5vcQ7GwTeT
WMRonRUZc6ZpQi6DPAXuGQJFm1d4LpoI2AjamsNUBHH0f5+wxqJbzjJZqjkAymH0
3YsbKlTCZ4uElDcAWr4RaOPjphkD2agOWrjjRRpaX+cj0S9Y5LT2IqbWRFZsYIYy
s6eotXZvbkecjzH8roQlj7OmcDng4aXFafT+WLKlxoASdoGhamyOZeG92KjAa0Sn
TWoijxX9/Mx+4cNGQyeOKCH4O1MsVgY5iTob98PUNj4otVd8beaklz6qyMPKSnOi
gJoBfMcofa+PxfQh8hzYg8ZQ8bBrR0/Jc0wGJNDW2dy1W8y4vYlmaWlnY2mzcJpH
QUro8hRs6Vtw0lbbB5CIDSXLCEbDM+UMa8DeRurD13hNDkacQUIg40wt353BZFAP
g50zfIzfvnKZABUosVWU2FVa7JLbmtSfa+Ih4vVPcMthjvYSIZPOLoUNRutkARE4
GlPMW1sVxFPiSE8Av8kLNQvKp5O4bzqogiCcM9konF/M77rccOvsRQD+ndj8RN0K
KV1ZL/uGWAQBPB8QPd7RJcRfxWjgKos2fydRVj1tyjCYV6Usg3x1mkOBeBqIMU2U
BWkXUc65MKKx3H6H/DxaJahHXtPvAp3THgRLx6lcthHNTPmGtzjGN67/Qc1wapud
uziMnekD1UeoIT23a4wsGgPv2ur87zggH9R35AN66fXcTh7QP7PsBll2iyQZX09M
sj+cMNXLyL9HPFxs0+oRKYomXNXNo1HKccCs45ufhJwlUEqkFC8iubZwMvyQcy89
qtY5ucRHBbCu80em0zWzj+gTqEk/gRgf73TDUgAPEKa36q9QDweyCfJFM165Kd+Y
YKj/K5mze1kpg9uI7JaUnyFSzksEr70bVfDscJyQI6Shz63rn9w6Ax52d+o2WGIw
6yPewCHxSk3bGsMCMlu2isI14w92FLBdA2x6Pgn8M8hyCb9ukS6RMapwa12Wln43
oyK9UNZ6SGEpUw9Eee/29ZQyrbww0rpFkKAf8TzGKrNc4fN3Jb4RMIEsLvTvVybd
hIAbJ2bRBugxr7USmFxxSNXtKTCu+AHZf3izfgbGDuDXPFLozLXb1ZNIjNV8EjTw
S7hQuFHhwcMDt/ZX6QmAHbGgWlnjiA1f7Y6YihkIbAS/OwjMjVkqBsSxSfhD/GcR
wgkHyS0oyGNNT0j6RQLiiAqc6YVuzeaTu2I0yPdeww65a4tpNJfCS3hB01dVe0pd
vm93y4pZO1E1BDr9EaQLdplQykntKVygMTqlmte6JWNqL6y1tf9IWICiWywZI27e
/jBwDaux4nORQbnfOk9MoHJ18aosAFXQWuw5SWq1BmELjN/IF0ZKip7W8RLoxwAx
fhpbCracdep3FX3dejb3514+cOv1aeBrTfJb9KUlVYWgWEn4Y6MTtmIr7u4PQK95
KJ0ESOHTLEENk+b/04Mni8Wc+b7EqvoRKknluyg9ffEHtAbZASXeAHdNlHHvsNtg
jbbyLRiqTEOyICq8gsy3cv8HHA9sXi3GDl6356cQG3tuVTvc0+O6GkMIasmrg1ky
GHnHZTSbmklk/3fZgsTORNK+W5fWhAmU1np71C6AUf+Ecv9P+rhd5I6L3A0p1I/6
6CNAK24eCk0ckiOINaufBqRAAhp+x62nld73H8Y6kzMCWYXySyxCgnHqUo0i/+ft
EvFXlTN5J5OswV+G1t7XpGWb3evAV4yGd29SnBs3dqAs01M9pNaVNvQmkopu9rdz
F45/JRfKWP9XTkA0TrwRtHTbmiIAE8ShFWQtkHr83vcvL6Na3uVV7cS7TEQTW9AX
PJLsRoJD67i+ZyiljauHLpG2w9C9AoXcmEeMZ+9f22cf0slRZIm7wcnKRliRZDAq
QBuOMx8+z36JyTUzt4WCwnDC6lt/CoXuvkV3Xyc2mrtc46SeLHbaPZ8+UVGM+40T
1nY3caYckAroBwiic5tIJEJwapb/rcumSFeOz854WU/AJtKAZujwD7KYoS1nKkYu
DH4K+cF+Vq7FpG/PJcGgE201Csyx+sxzQCGjgoNYASDT1cN+jtinoZvkv8u/Gl5r
WhlOuBTTaAV8sj7jO3f+ijxKu2Qj9IUA3yTluN3s5Hj6zyef0S9FcZuTCuSidGqZ
LnmcYrT38LZnK2Or/xqbQdt9u9Ta2EQXw19A+JegotFg6EwTqdgLwagaosWaDZs9
9Q9/b5EFX4JSux0/UNE+oifOiABeZvXjBCtPhmg44RCgzWUmhvmI03y49V4SInvm
R9OfEf9V4/6e/jks0/Dzw6LQKqSGd4buh2+ZuIX2HLIl+IsW7KpOVeo1Bzc1zfHx
rRohaT7l+sJA/9Zmarsdmju7PAwoe81bLhC3bxkBdSxCFkzChrwgF7ZCkoj+UBlc
2ywRfDGVtPZtOH/BbmscZloW/nJBCTXiPxLR+RIteVE3FD0c3yEpmO8Tkik6fnFB
9o7gtIaFh12IhLDedcVitHPZ/b/K74l9/Jb2OX179OFZTib1IBbgE2ITO+WjLJ0c
5e/hJ3TX5CF2SrQKcx4DLBoy1AovZXqeu6xgq8RHoMiw7kvf2/qJuQgjAzHnobzD
WChNoLH18ZY3tw7PmwX8WfBuUi+qaN51M6t4h+rW0McDyIWI8uppzPIXyzk71YQ3
l7/BIYs1IbnrQwC+mHGrHp8hlkU9WCjDyzWimjG1QyUe9C18PAdkQLItBAga7ZLq
5+fcGTPCAOKoh2+QxSPlx9qvUpYdUjS5GDV6xOnB2S6TBIweu/9HvhSMF8DavdJL
bziACYpHP/cehJexyonSTpFEY0EZCJQB71gHSgJHNndZcjfAgSMFZHU0OdGZNjzL
Hf5uVISVuarW9Veh8FEejRBK6hZAVrDVcb8+6Jh4DJ4ZOfhQWOtqq1nIg9yvkj2z
mza0i6M+VIpq3TYyoL3Qan4AdRAZ7RqQH1GX3UQ3VNrgBS5g0nTOOfMX+9DTBrgu
idPuKEyWr7sbxNu3NqGM9bpdP12We1RUhZlE+t0rM6YgtbIAJ6/jfrJBJxw7NUe3
37OtzCZhA1q0wNXhV45y69D2N0y+0GhuEKvoB8SYNISQNjdyCZWVtDza/YAdXqIa
wLQiJa4hgijeEkhNnK11+ojE1+0OO6P5VMk0RLFwrg+MXXKzN9xBBftCeHwCJt5t
IIvIR5zG22/mn311bl0+CNUN86ntATIRZcLSU90dl8hwvHjmNsjThisk/xBGfQPC
o6pY14PmxJ0rB3r/Gy2onPHdOMewEf7qCcxGeTm4+9dhtE3RXxGwaVTIxpDVz0uB
DWnwfRaisV+PnxLNqkgNr6XuVw2cA7A++8DSul/8CTWRVXZnqTdW10+PQ+TM2sox
0d0HkuxM3HpjFut28picCAZVRpxZAr4CVYcHPvPUe1WKzI1xoPFSKNEAfRRVOoXK
jhFAmIEH+QtO1KnCqG2ebi5wtHQUJ8FF7xRK11oArX7KxtWt1en+ZeYC77YmQbiW
zGpTCZaIFANrHiwl8Hr57VDRElLyVS8kbZ81d0CYeFoTPPJ0QByBI+cNgJHht+zZ
e/dILWxADtWwdyde+awOJnsV6EbtgsvJLzOC5TZ8yBtJy3cognQq5KJog8DKXS2o
YcBafvbmDWryvoTErK03vY5raY8TpUCHyb8wUcrioOmOzM1KSUSRaseQ6G4wuogB
`protect END_PROTECTED
