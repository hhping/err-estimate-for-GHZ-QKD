`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5fOtk0D3sVvjrMjnNpfSnkv1XKTCyVzFN4GoPzlM3ws3i1rOUicDRgDvhhVAXMj
80DMGhV+vlwSoLSjdH7eIBSTFdiaOVbxWUJVnFeARHbRfY1K9BJku/9dC3cP9khc
SbyNjij2dtdVV0e49B4c63w+fQJ5Y+mCKcbwWaNAYEjy/aiNiTgeOUvmhDkWnklj
5qBGf3rbswbZAcf77174TFTdtZyOi1Noe23nQgBPnPUdwgz+R/9rZYvdhefstiVN
AlHjh5AyhM4yQEXDFKxhrYraam8hYyh3AyZTM8a/jbuzAyvSUd0m9LRMH8XAFLqL
+kw/abKEzTzb7VFGMckhGHQOGcyJG3EFaHeGf/vYBG4YcdU3r15bFpP1WuMGmmWc
QVj1O9ls/f33YUTp+G/Z0nI41lbyGPYOQR+4BGG0LMLNQ1GhZZ1X5ipCHLRD7cKh
V1noPLI7DgY+X/AWCEhAOWl4XVDSUu/oM25J0k+nQ1vAB1sduaciOUtMmKzzue/+
ZGjhs3vZKkKZemqs9zkjzLJzUuWAkZzh4aRADWvRnd6e3bM1SRdiv5aR5AwPbfPF
GrRnQ2tb3rQUz/racR/y9DuhFIGa/DeNcWY55pRkt7LcjJ9C4uzJrko0alhIRrb8
kkFKV1UWMJAft720k3oRSUCwxV3ruqCP1YmoNIvFsD8a4qN9K703RAB2eaS78+Ik
7GKdhgDzjk//gfQZN48okqZCjA91GqzkUwmTdseQkAlus6NateBMX4UG0Nj/Y2oB
S2FBZBx3eit6IZe+jE1ymTRiyoEeJaX5noGReUmvECTtYPiQtX1Qkt3GvjKikbnG
`protect END_PROTECTED
