`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e2jgrXgLDEL0WSrxLItsWottAI4+hr3AFSzexJNOGJ3WERhGXrh9Ica1MTW47ML7
OTygiGm75IudnZUH/1MAkLkfQPKZ2476TzbemDBNt4ykwWo5hPVRRLmpoW88HG6v
bbSp2sp0DGzYrwD1oiuq6BvYg+AXOnnWlyJXZlQhpZHLEDdiH+TfCGpgzsPUzsH9
pNB8x3QCNkydG8cej5mJneZJrp8S7GPIXm4MQPSEnacvKQH9bNseSoodLHPBlqwL
nJMTXWipvrbGxhEhPrbfPUrSObToT3HmXTjVd9PZuH4P4H0a0OWvtSeMoM20YsYD
AzNdxyyaqijysjvWpTUMFNmD3gKyIA2HTzOYLuUKptzHf3+RN7R/v87GpoFqulsj
RA6ooJ3DFklo5Tdg1vSOWupILJBlMgTuxMzs1odh4Rg9kxUQBJZiKyFiFJ0I6fA+
oeZr+j2fXpfZ/kJxwyuW+0bS1+27vfjKOYaPB6hg6hKEPG9W+x6kVTu8lV3LN5rD
inpbtnbUwycfkgdJ0Bnl9UAfFCogyhhu28DG66SlhxE3yNAsXIDBwbDeNXqwhH/S
1jV/QRZkkGj3oAjYyQVdYDSQHcwVErgbD9fODNQAoN77GqcO+7qJvjZqKGT8Fzjm
HsRe4m7TUlcUOAT66vTFdPjkXbb99lLqbos+udChXeltMM0739M9bRObicBRrZ1g
sgX2vDCdU8YonlCKUWZ2BgDfRQYJCB2K7uVgqvJKtHTxsZCPbYEaukZh2T5KIF4t
nYih17/PkOueLEu64NXSXIXi2QmU9UsQOyMBLx2lfFppOpAsAcaZp2OoZp4uXTqN
eE9sFOEG14jk6gYSgtEUECbTGaBdkRDOotNSRuyiOYJ/6P8BAP+aIj5/KhjenoPh
B8GCV6n4X+cMtmfHDifJCrbN4wbmj7aLf5RSkIUf9Jhv0K1SoUx8GL+VdlxufV8g
twjqU5sLc/iW+Ndxz5DKtAX0oJwjSJIiNNsuLeyVtJHMBLosF/16OzQ3YU7OVxTW
KadfjiiWGHSIy9hEwpp2zcJd2n+1+DA8JNaXCT98TJmNO28ZV4diC29hAepHm/Yh
DPK2/SA+H+d/OhpjPs8GzHcy95lJOZ2GxA+DnyFX5/pIAJDNIiy1tAbhRb6NQ/fh
unySPq3uSvTV7F9tYcGKzKqr4XfQFubq92eoiD6sW6EGRlm/VXGCE0Oldxk9FRym
Dt2um1c0sJl3EfFh37+2ml3+LrU5tHCVpIXTTELOHdeeHGOVdEDK4gzkrV6RGUnk
bexLHrX2EuVz0es0qj7umZyWeA4gzXrw4EibKZOCxZvwpqIuCaQo7O4wdzt2Akey
WprLBGcrVbPSDTnMebohCur8WVUkfDNEPQL8ezAeFOGLVi/pR/RXmjrJI+fr3aWU
oomZEeeAlEXWGqtU2SbydL24nyvcgN+OguuTZQHO0pMbWrM8yJEtqq1xZnSrXECK
q6tvMV10FvZ2A+69tt5rJV8fH0ilUqcy5Ek85+ObBpxzAIOfHkpEVQwZUpx5gz1F
2d9TuTLrtv0GQEZYTSCZ44lnx2yOboDbKbK7Rt0w/C1Vxa+ySCKhlCS6y8dNsU1/
HEumIZh+092br8ayl5N27ydwXBDBFUuSb3ecY2XugLAMhBfiWGccbS6XNzDvsNmx
6dwi/pvPd7low882jBxYJCAKMSZc80FK0ghXy+UKHm6hfQfxBaMM+SCiWUiijK3y
7PcbefcoCjcUOLt+Z/HOIQhYap8keEt0yc6JGWWuKHHF6dtFF+U5gJVdsFda8YMy
cjIYKlEQpSU2QyxtmokmXfOIW68q3RmBIfgZgWOan0zrOdrpTJ9+zO+wj4sh/kOW
LBbYAv2ce1jEeC2PAiup3BF7j1MCijcAxZGF8Pod9Nt5007DWD3w7hBOrbmQt/Sy
LCSlvoGfX8+YaCA6WACdGS3sKK/G5vrMWWXryIOSdiWGpr3zIvauxBfrNpg2bFgU
pk4OYPdezqPGzGb1prFFzf2Aq5a2rEpLKd8BTxKDGbPHe2WZSqS7gzQo8ZhFWHin
midwtOjrnQed647mx3EkaKK8INMXkWHHMUBoH+UNL9ejN0WZ0QCvb4kxSM2mlKCK
C19H9m/bF8AvBQCi6jXyLBkIx2m1ZEWohWeSO7Sm0jUTkYQmLaOuL8mBDTkGqgt0
0FhB9StyFbHpMr9lnBlq5NIMLF2BvOkW/6iXZ4M6npeMroC/Cpdy0cZbQJ4381WN
1CYbfxGCQ9yh96pDRsMKomorPKsKpYxrTEZR9oIFtSBl7jNJz8UtuooGMGd4IDIZ
qea5tzSrZrvY4AVhd+h793jw0N7VSljD54eBavVuVvErhnXZldLXUN06UeE1g+G1
27ykDsmTvP8XSsPzt09yahT2sT34k0yKlMt4Z+xbCBZ+gffSV0T48Vak7XlTh8Ie
GAVV0eT0ouHwHzSrql1ou0UFuGnysa2oFu0TdLMnQXfmY147Kpxp3XGn2nk8lE+q
lVo4+5OgGjyScC2CjUhnNuXRAAuqLE2Bservs1kKd49y/bx6q4JzB/KoNs9bayeR
7fnLZaPkUTmLGl0GyscPz7VtJDCCTK09G/7KNdJJ6XJlBadJDb2KGnfJS5DnNpVG
1liX0uDOawSVtqD76S1mIod7jyASsRwPWiIcZXv7YKqeJvODKGpjD1XD3ZlzE6Fn
pdviW06tcXosQuWQiVBbJQZ485CVTJoA08bn7II1XatX6NhOp2Zyw9ULqEmqm6lC
ooJb5+bG6CN7Z4gFRg5tPsmqW/a/D45nsAGWhSGAH1fMUV6dQZh/AnWgTZgbr9QH
N1P9iDV+H2kWSDn5rPBoNw4tTfinos6sl3LObp/l358qCUly3d4rCgyCSKs3lVTK
Z/osfmLNPHY+qlo8Aj9YBskiaFDudu7cc2bSczQ2c01DTouwgdaq6BfQ6bGRzOFI
9y2wbxa0Os9Hi7/zHzjVlBWL2U7o8RtEQZMwunTXHvSKgEf6mRhXFYW4RlppJle+
4jXm0ONEK6xA8Y4xmj68saKR2oMw/JTHbs0plOmf4JlM77NcIqI51bickohqaPmJ
6LzEinieOA4E3tIw2GnKdeOfbpQdbFi67a/QwHX9Wd4pGha9xunOjzr5VvEiKDf7
a5SQvzijlA4P2pV/zRmve/Q06rLJU2Tg2oBpZ4ulysjvsYZU9sIxJT2z1Sw+Joo+
tD83ki98Zs0uLqM4z0pKShDROKDreBohwnYrEwqXkyenf9kg9W8NLFysoFNxNqFl
dU+K8nn2Qw4VD23JglA+6hLR2Nu6UWa0VMr0pltCJOI17geyDCi0ZM8L9gnkqc4u
RLy0WbL4ehsINnLSXpKmqUDSEDbUO/Ji8e+WzQbC9qD/0fYyCq/wnjdi4QR93O7j
681Act+lc46c1NHikDi2FS4P7p3/u/OA0b0817damGShcolZdXf6zAZDQ+tLp4xF
PAHr5i1by8g/MLeBj4UA0WAzwagqKjeKPk5at50o/OJquSY8PeWMnmYaE94XV4Um
R33QEHmFJnO2Df6wln7mVi/7KqmdH8duldFV0j/bI3QkrBj3bH5C5LUklWIXkHmS
o5mY6rHKPC2iQb9cpXBmTjKh2Zr2jjVtwL3V9LYnanH5hLUlB4MDRIeusIPGtbrX
ThzcnrOJbO9lLbehpxexPTHztUPKcr86wLNyQC6q9D/ojfuF38+QuErZd+c6HQTB
WU0zzj46SC/AsDjRUaYAeAV3y7yLdNJVIbcfT04Tbyj0IiIi/4whWTLHfzKYNXux
+9KBQtdGpNcgZODaNFxIMpS3vpQNrbmNbeFThCIWaQlbjSBC/zWThRKnXFRCxSaY
/JluwUQ9s2pb5nGxj6Y0WAAkRBjTpqcfAxDh9UsAGAvwbvAvhtIugFlLEgHRGX6p
YAx66c/+hoxs+iJfZaNBTec0kKhAa5kRiwHInbGQ+6ccEwIaRhpoiCHEOjD+Iv2S
Tmq345sfkOV8vMAqposxKHIdNSu8HMLXCGeWItry8NXreUiCiYGp+nicwYUY1qht
tj5K0ZiCO98wl/TzY83gYiYw3kSEkz9ezr3p5nWRaSYfTFU9ySedYeHTeeXXOFjP
MqhSu5z1S7aKH2iTJdtvxSY/VFugrc4wRlV+FFP9A7CMFBWX8rAzM8LECoLfxN8n
V4I4xVON4+oCdFYYDR0o0opG5TT6TmEwv4UIqh+NALmUfUacO5DUw38xcK3W3j+u
3b8Szs6gjKOt38UT/sFqcc+zVuf7sPlYOt1ZcISO+BSbaZXjzi2AnEnd+TtuqhxP
Clj/RMrhQOBhqFxIGqEpGxpnxYCKIdw2wQoOfY3XqRrMAwvx+4z5+VLoRvewG/A6
Vpqh/bVHMSwjV4rFd5Bp7AkwHWh9VZWqKKeYy8G4T6snZIspRyeQI7JySoR7LgZC
XtAODRqPXhEB9ZBgczbkT8JR0hYWG5Y2h72+w1NpYbyy3ZGFI0e+Poj9KjE35HxD
mw1x/vhDh+aApVbRwrGLRAkRsxNZbSv9xRQsnggUHcd+wYPyeaK3ZFCAfogKdIw0
u/ydgwjrgP8o9UMVJrrrMIFYbQtrBiIZb3+cKW7Xd4Hxdcj//gcqA7qpBFKMhu7K
JZyXRb9rSilbWdI4bR/na8B/Kdg1s3KLljd/xWIsOHJA7o7BNfHxcabx+uFJ2+o6
qbXztvcjlwyfRJu294tvb8+4Fsts/PC+nz8QeHI4T4DLtkGNLqfV4/YR5YHSOOXO
ZMlrWEqoG2Nsb1pmSns7pU7DRsrp+0eeYqq4gsqJhfOezD89T0k0v4tiCEWjDJYY
3pEfrqBsqCfQ6mgWrE+ELrYBiEIHdxF41CxQXiVhf0NqJeON7mIUzvUAkBcOBTLZ
Fkt6Xw8Npn8AvjDTtATjWn5oMjE44D0Sj/UiIgIf2fe3hjZ9SIhNx2cuCKOnWumr
jAC+dhcrhIwjMZlJ0mgH82HYZPIMyIBaprCQbryNWq8lvYBZS2EZ0qB3oVAwWm+l
e14vw2fQoWe2cqLbqTskO1AFg6Erzn572VQailw0BqSCuarEaajR1SnpEkkXy6mc
+/jz55FjLMo4AyQJP2JdelaouJlZq13epSVYgStqIWgMLeX9C+PbuYf29JgzFX8k
qsO6YyzFDpmTHTwm2ik0P30doxfthNWjx1jGNm35/O8yhHfdJ7Y44qE86gwig6eU
KTC0ao5tadB8wl++h4mHdmg7KU2txb1EFNQHlYyY+IXO/OEl4RT+JJIYyB7WWVkh
lh+avdXHZsfAVqsIR0gtaqXYuSwhjYZvNDqc/HAPsUF9CvENN4qEvig05KIbmvJ/
T7my/Qb+xXKsGIWy/qgMHGnIVj6bNlnGAKWQb53CaxkYMOj5hLa5yPpPVR4Umt7Z
NYSlq5V5ro2s6HZfoZ4QFnWX/YhMIwbc9X4GwmceoaxV476Gm6xYBwF/LNwFho5Z
12StoATzHAwd1MrPcOgE+2/yEP/dEHRZEAffD4k2VmkC1nuUJG41/EmCZnuuM102
AbGvCtcIScuiwILWFwQRnWXeFU00NCiKv2pqtLUCB6CFzhdLaSecwI1yaW8Ey1B6
SwPgOG4gCg/nLxpox0OAAwFYNDkz19UHy3pZuSpZedKL8dClAXnvojw2r7oB0+pE
3qInmUifWslKNUVLaLLZ67SRzqQyAC0bM4+m5V2xE36IPYSqjy/nIm9CmAwfE9O+
HnJAYc1hREvB9afH9RdOh3SNcmyK2R7tU+JmFl/5KkhzkKTWpmeaKZH83o/OWOFo
81b3KuzzvO3u3+85QEsf+RYxoS1yRCCzbahnbNRWMND/cIvNEtpLeKHW/f6UvDFO
SwPi0w1RTwqw70SZL+Kj7KFeBqBXDSD3XA2KgQRePeOQngWkVmZT2ZeB6gepTpcY
fcfKXAHVxtFZwLn4A822WjA4f87Wu2hnG/6cQmOGQylXYJvLZ6BrLgewadiLPqLK
4Vx8cq4ShykNNChGsDU9zbug9ayrUUpdJAvq5VZrkuv8kaLMswcTeBTt1CeDkEfv
Vx253shnGwoFqHLtLe7UMiUOcAbL0Ozf5VSQuAtU7DMd23T8kFY4T0Un+5vsRM5c
kVc08V2R/o5IN8ppi8F7bfziu1eR+0HyPOyttYJVboEO6+5DIBxPSFY/m7v6Ehvl
35R3mt9V1mV5vKFksp2Yt4494EnLuQh2LmF6yBx5HIsZLj8T3mLzzg1wubDBSOeo
Csve1GdNOaVwLQ6MD0jAHoudtw+j7heusgMWECKNj/a5Ro/77kzue5Qub+YxObz1
AIndG5uMLdC5fHl1PkHGvEkAYulziNDfc3olcUymqQn9ibkuS6iRA+Lw06wfIXjS
rk7dCx3pD8L2w3zFJQCmmIcPXh+uhASTHQaXKISa1IvcD2R7koDtHHjSi4SIWpe+
lOrgH2aoWyfPDjM6sSrV50hA0LX0bx7qgxTgDSRQp7JIIHL/VNTLzhdsOKJ+MTv5
lhjpp3BDOHCfZGpCOEDg416kHxsdMjlqJ6pwyeKD7epCyq9g4BAnKvMKF8Pwk7kX
LRGxnMp0s7u9dfDiICv5osJER81Fp2NgcfRwJxFZRRJOLSx1Y1S3KTEBSDQzoZQe
5dvdlLyJ1heBI4757eqXTA3gv+MzlxJpfx7plJufL3LN/USoJWWNsnI0Eeno4iLS
3zcN/YaSbRt8ICbhsI42foEWQK7SWqQqdQpVGBIyCe69f3qKQ3C9/Kh9wsVS6XOz
s9B3bEuU68+U6sACIMuwAIB/dg/6UjH8/ooh7Up5l71pvQ2y0E4v2/+LnkGD1kdA
xMTalhFgM3U13RypZrDnKH5/NU6kKoc73gafnUAO+z0rGalLfD24zdwqkWndwqdw
h81tyEDE6r3QxHkUGPFD9KCPnLKUPPkDArKObhNeAL+SmiXzBneLXtcpKbf2njU1
TQbBjYpphKFdeW2vTftxltHxXJ/CkoRW2G6Mx9aIHivyh9T4ZcTiFExluDTPWYjw
8nwIbLvWL3NlkSpnDAPTHTaHwv9WJCdcKO32f8iPQoYJ/18FS896/To2ER5jrZ/1
M5zJ+tDaPMYBP2kZgSPg+aLJIIImiWf2GKaypGq40eF2j7PUPVEV79KjgCez9rwF
p0mg+W11sSk/DE8bYm5ciumZobXyfqKckjvIwN7n5Cc/8Ck0pOG17U0uPBTjyQju
dILA2eRk4I2PvvIuH+BiHo8mM8yuYEZbUIsQH++iuGE8GgKWmhFxEWq2d8ZhUtSk
mnXzzUGEjFubRISeXaXaVCvmw3JWvJJyptSGQV+8dEX00qODF0HWhOmxx7r5nHmU
TdQojl/OnqOXTzoxAT4cr8S0XleQ61ymEfbwsLSMAtahYsgxOPxoZSvG3hR/m9Ae
gqLD5Ati7nYZqkCPcPIOawVj3R0/Q5KxDxDWJr2B5M31PDjPGdymilWemOzwRkvM
lDiv+xmoGYlhxU4NXwPSn9/lE8l+deWvqG5mO17c+gG79sDHQjFFD+idqsi3zSAO
fpfjXKiyodCpGRxI65pzB6obd/UWNTzkocIQ13KdCG6tQHEThAQ50zXDhViL4Esf
rjx+pTtnhVpPi/F37vRxTSwkN/YvNHHPWEDFVVTWdqSOggPrzD5sSMAaChp/8yvu
sohNO164NPFyCrCkvgXIU06SBXJJAq+EMKFPQG1qmQ9FM/dkzoI7fgMvo5vagNpr
5auynyyZydTAh4z0wF8XQW4keDbuqUWmM55SrIgG8NS/KphH3VWejr7AcaSIEacM
PNxUlij88X7AKqsMVtmq6fhofTUe1ZOI8sKry+Xk/WdwuA42d1aASVFCyY20Qho8
0T8D1hV0XmoG6uaIccrtfxgPwYDEaIk+5yVsV9bpcNztJwN/aJW0AffPCTI4CAg+
U6a9s6azkwqbd0dndnQMxFCS/hGW+KRkJGAnQ65oDNhBjp8Ke9yo7DwnWFYriA15
ojJWwCJRHiHyR+WljJGziYKJjgAISWdHYkMWN+iQQrgeBtCgau1tEudgpM3J4HCW
hvGwbffLm1uFUopE20sL3DyYgv95dIYg3Dyc9QStUwpqlKCeS61hOBwlMYkHXzLS
8UFuWwv9lAW3fW8T3lSFDcEJKgz9zu5it+BhRCpxswev61YeMHh6rXgeacb3YLD/
9YnSZSIJ6GlP1gdiMCnqTe8uX0LeGMPDUdHwqCb64kr4ZaFpZ+a2d3zMZdg76bkE
PxYa5W7y2R6GzQANIGyEhsi9qe1Q68v2WWRpW0Yzue0GAICjrGZ67JZk3s6mr2uF
IxTptJLTJAFWZh5p/s5S4WU0cgPIxEmQU9FrdHvgix9xqU0F/EfCRZH8a7cgmhVE
47oxjfKjSa/1isGGHLj8pgCmCyIEKrGrQoJ/PbS3x9qA4afKLJPvVHXlLILzXlkM
L/VG5XQPz42RcGO2FAz5uJWRRLOpOq8hpRJRRlW9uqhHOcdqjF5V6vYuuxEHZzcJ
mc4e2jK0zQb5bSJEyPdMLKcVxDT+Jhc1a4veP82gQgGt1NBRGDZsq0HoXGFTnV75
l6C2BM7wor/oqmQVAHZP/5LBngw5X0P+BrCP2kPEV6ZzDn6DD+RLdXo8w34mehjB
3Q2yKbu7YTreoeGLkkSeelK2yU12Vedam1DUL+5KNle0Kfj3B4bwkHLQUIsyT/c3
hhh23KAdgBfM2LVgiQ+ejaMQkatJlkh1uxInGeoTsF5K7a42atJF7bRcatl3Rhxr
9SMPrDlquQFVjTBPFmo/+XBMSjWG/Xo666V5yA4sQED371c4m2/e98Ou6QmUhLRx
R6RGLu5Bb6KL8TR4jTVGm96zf+PlTaAjFFURSxB7pa4O9OBfe+XC9o88Kv/sWoBI
7bEIWVohAllZHoQpxyc1OphRv6Ylfe7DxfS7p5zfl+5E5VBlczhKmm691aI603RT
/yw7hgGvbxruDP4p8aCVBcr9v0u8TEzJj7S1Zcb4U5QwiQyeibrDlXQtdcXxiZ9f
faxOyzHw1L7+JjE0P2szu3vXzVGyhBK+a1176NsQGC6h/BPKdTtcv6jTToynyVWJ
y3vUzH6HYDLk6iRTztJIO6TCGYa5VQW/7XERuTTfe63wCk6iZwy58M7s5N/SKYm6
vxKENXLx7SMQuDrwKLKidBCg1IBw1Wrl1/YewAAaK9jMse7rhI+21tgnFxfNsM65
o9QhgDlR6BhDa3wAbz/qhoEmkewq3xmBdnQFaLPIha27z4hCwnzB8f2fMk+T/Of/
69BsrFzeF/5pYGFIq8LIXD7numO3SzKRm5ToPENxB6JWr8g7T63xTT2N54C/OSLs
BVY5cymrodN2X3ufLLuGCWuOR+Fn2vx9oAHtv64qAfhezHp32nO5tOvDyFzNPfnw
j9nvsF6r1X/7y492X8mTgzTRqt0m8MT6HeeQQNOMQaYE5nSZu+Vq2xvF9B9Yt+1S
rbSuij8g7N1mPrQyuNPjXlghbaq3bARz55h7OU/Dh6e35vUnzH7SJIP1Lo2uSwAe
gnXZPaVBuNA0VkYHGZ/24etOVIzlEpDoVbogjdCdlaQdvV64tmYskrD2kaH/uGmq
l18gWovISQ3flnIkoT7JSvBJWDkhjDqx1khQ4We7NzIwn4ItQYr5Ed51M7WfcLzJ
MA28VvREjvOQY7zjbZT46lBuCr0Pfd6SuVkmHsUlGEFkLkqAwgB173OcPMCZSyt0
xGwlhhJLk2/eAO2leHRF1nDZxnP2yvZENKPhgQ0yOX9updWFfmje+uF4i884hNG9
H9RyKWmX7WCuNHJz9WUm+jnfsNMUGzn6uGXZyghrf4E5Vga4QSWHoWISbqIV23vt
IluSeQVyOCp2ggzr4SMjyR+X5/XIuWasbYuaj7uOdvyqob6yX2gqYgQhwiw/e62j
uBzTca4IGFIk3M2FzrKQjvNsqDJ9xN6/db129668AQwwWXqCGMqqbOvis5BF8oEz
AaMf1iIczCmtF2Eay6cxzhLXqcgrpVYqDVbpWFOVbvIdfixt+IQyVrE5qlyWTGol
OhMTsv/rZ+hojenYewHq+O6wR20cS3/JngjC16DMvQNuvqmVZJK6Mx4y33ttijT7
/KJTvmyKM/3YKwbVoZirss0as0Uc4udl6ZMdf1Xoj8YUgvNj0cno9wyrSdVki353
HaOXoGlreJHmSCPdY7rzSt5qOtLsZ0GMB2zHrIRqi/I7LejOOBWZ1rOL5HoeLYj0
dNOKzvVVwXB8LkyHI5ziwUfvKdZZYFmE2F/4x+av6m2sLfmmTFQZUswJW61Ms/wa
zxeHUoIQozt3JvjDkc+P8Y8X34JZZbmxkE0k1rgBueuw516DSSeYIIM9kVbkgbHF
yRtGb2W0jvArWTzr473U7TGT1oVokBVszGnFOOxDY4J6UWcA7e2+4ei5yIstBSGs
d+JfRYwUGcF0agjUXRfLZPp+zHS+OqzfcZxtXxDXmbwp1S1XPDMHL39Bah9JPsXJ
p/TaRfNGxUXluFVr09P7S2ZSLmA9pqQ9Q2UXxdmUQyAjQzByDirmDQ6w70ULSxuo
QLqdBnReIRtguaI8+apek9MK+hraxaBvZJ7B/4LB+Tw98tLKTdgRfS32qm9S8fc2
Ah07HcAVJA7TcbDCV0RYpDcnBHuCRgGn5TiWbYxsKBSvt8KFJj9y8K9gOj2xlbJG
VarxXxn4hOt7VvimHzWx3XbyLIG8MRGEQefufAipz6j+y5YF8GTHWGiqYMwvzsQL
YeKSCwfhoSxgJOkLy2NHrrXNbKc3vOR2qWC9NbJVjlPXHCtrHj72HvZI/YhisGAy
yetVI+NTyftK2fwoi/6BaR10eQNYHrGFhPbpQzpT+DftxTaiTbMdli9eIrF3EFsg
EQPpDYmwVlp3ypsRR7a/BxdhkdngspktTHs1+xtmIKM=
`protect END_PROTECTED
