`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZ/ZwC+nmTtQsIpepiJGr+owL01IcfVjgjao/GaNoSnWTbQV8uFxsBPZsE6Kc3ri
8kXguHTnDyGIv815O2zXrMJq7pM77PbgpWKQwuuNDKzb29v9gx1PoeEjCq8ptZnT
gJnW371Dvumlm1qM6RTS5bnjBP+PsZ/bWzYfMTUmwIIb54cwj2YJdlFhgKdi0Jcs
x1fC5wwhyj7aEvFGGd2QHy2CE9zpEXxh5uCm07X6f0k07m6Z5uELRTklXoxmCGZc
+3zNpR6yyzLasqlFFciOI1lzGX9NlnHbEXoAuqbtoVuG8fY8b/eh7syMG03H3eBy
MIeKLkFfGW1SaljozOr5FlEThdRXMYDbBHUt8rrPVdNnBmH/cT0m4g9+B9t3vIJ5
xzRbNWbFl7/cX+efwZ9EM8NHFgurmb6SPESBi2+i4YTqseiGgEEGsvBIYkhKLZPh
T57fpAI7IWNVobTNSyDgAiMJtOcmMv6w87aSRfDMc646Vkb4YaR5YbQRa3iRws8o
Upw8UfNrzz21+WQP6JY1as5ybSJh4hp+j3SZrbgNki0pSsj47s4eN9cOgl5bIdbj
oZxTTOQsuQN76Au6y2MUQ0uPlcaClgr2ZNWE9QQjxOiPLr50ixYi8ZKSZxw36IfA
7iy+JUbOhRv0hQ4lhcWD0NChOM51fRwOJJi2pK7npOght7+mMnev2jr3ZEZ/27yC
s7NnHrFRIoJ1dweQWMKGnYZB8TsDL60S4kRcZ2/oOmc=
`protect END_PROTECTED
