`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5yjGMmuH1K+W2LLlqlsuVyb0Ii7ggMGvnYQiiNfGQrKSDfEsoX/8/7ay8LhUoGv
TmdM+RacxjSBbDY4S0gXQPWaUVwmuWbwODcZ54Lr9fGxgrOh/y0KllkqPbh+rvOC
dEOEVXpkdwwKcKBhIGxiYOECm4hS+XMVMIYevmpwCwZ/RVC5CAsWDabzJyZXX6I/
EorNY+xi8wg3js+UIbPq96OGh621ePxSl6GeYhUsZLllAtLTg0bWw1qemFRBzvYI
nz4DRL8Nz7etLV8EVmKWb3dzTbUMHeOeyp+YDDyIt3A09kXrx8uhyTTtuh0k1BGK
Jd0KVdjUmMxmMROKzHAr8KxgeDXna16eMD+0u1Ni981xlvrStTWKkFUI065Zoj7N
umGbw6YHSvuY8iekB7F6hVhpCcg+EC9J47Le83b+y1T8BivA3ZVyqufLB15Igddf
wSovopHuHfupsd2xqweLcDdf2B7LYhp1drZhRhEMAZM+kPnMw92IBZL5DbLtABul
d+atfYkACHouPReYbbFHE4LKH2P85wLSo0jadzUDxJ6OmKxy36g73WCdYivdreq+
c0Kb3P+h+XjumJ36cxq93UFWjVRrMVCnX+coZuf2ZQUKuwVg1wMwgcNTEzh7iSeR
au0pv8pfRysn6oOs5uub7NVi3Be5GCARDqOATBBE05EBgS0YYPgUXYCSKGc2Zd7M
doaQYuR1MO0gmywXU7cowDB1w9bBADkWkkL0Sz8BqH+5SeOIhzRHJYF4k51HWDVl
uFM5JRrDh3AbLcQtKb1A3OwuR4XA7Tlme93JzujwsUu/hNVfmu890Kjfh3qLD+6G
7lTAabD62BNYww1NEZrYmPwjDtHTCxjmB5CmzvWEvZVktuWPPX6ak05kmBjRdnBh
hkbQ/ylOieuzo5TDO/qx1vZ9E+/f5WlaM598z2HmKjl2bR3RqR+ktVRdD6gwvzUG
QEqDhWUpns0Ga6fKyElKWer0dxDv2p5MzmOekfCsIWfBbSo5jM9wxKhhGVZDIOKc
cyWM2xKFSTTwzdAW+y4lYgC+UyDP4vVkMvPtdbrYEVXpGRIczFfDH7k3Nh1d/UqM
/VheTSuEU7kqN79bv9bbEfNd2GIXoxObSZwv2BdbTXPfR8UlUsstJiiqlFtMPt5j
L/ZTtCfnEgumC9WbsX30XAojygaO8tkWXZ0pTwehchHPAGnukQH4HWY0zck6GaYP
C4R94DgVwAHARdRTcCybIg==
`protect END_PROTECTED
