`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ANKRrx4kyz96D39+Y3kGjxqK1NGu8s7GacV8gOtt45kjNV47Tj8O7cl5H8Hbyq7j
AUzWNtYuxxXOS7weXiMA7t9LA2o9ptNPAAeHFYbyIhlQWGjjHYilqnpuYONxI6P9
sI8vOONUsZCVfbBsWE1om1hkXOWyEHbTMVQ8HwKg20T0NtDmyXZtt8hp308TKRwO
6jCKNjYpl1cZguRF8IbnfbK6xHC/R+LsttPZFCTvmp1GQvssjMqisv0oKkPOwMjv
AZMCLhtL/k1FU949mL6Jmb17VsYMa/7upTCFE/RhWrGe8BtwFwcx3czFB8z0X4PP
U8WVuwOp9JXc3a0jPQZtBg87xUVsMQi4gClsbYvo5YoRg2csVtuINpZnjme/AZbf
UU8BA8sgLBz3/qsPevyO/KAMV+Y7KodPLlJOG/Bp7CWUDvxh6z4fNNZkaME+jq12
qwwVwIZSx+0H7XuhXFWkSfcU446Lg7IlPYZpg+4oxu5x1gdHdmaBhuh/JOxbVKs6
lnmZH24Wu7iBmMLpbryWBB5GtF38h/VzEBK6awVGsRDN+9F3lRIPLQSQYW4Isfil
P6neJDqxFpF6I+KA42aGDXqaU8jOxOQ7STcuK9AXYT8hA/WZn0+Xlg7cYjmnsEHJ
OSz6xud6aYDR2mM6yoJNb2I+8Pmmev4pfr7nVpLADGbeJXs58oRtGF6PM464EU9x
a/KJf8iPvm+UOqq8tmjo8cEa68Xerga2Cq77L3gBP9/6TtlOaJ65ryccPg/jXGpS
c0JYjiupffCod2otFLSpTAoK1vlWnpuoFlU72kvtLSoQCqKny4zuOkY3CZ4CU9TV
/D1SH6xMnka/eh0MPiS+EkHGaGpAxCHUCJdHg3YbkkU5wPiczu5lcGxmzncFHEc3
RpwWpMiUJtRDkSBtvyYr7WTvQ2OXbGmkhtpTo/l56lBvVsSId+duLTOmrEHrSIPB
M5YHcjxsUspywmZgz6d7CptjQQ2fZHYmkRMzK4ClrKu1kffoN+txp5b0wMyMbWWa
Z8s8pd8MEnWZ3JXozKfPvxa+1gCM09ZApJP0P2b1M36hJLfb2H5b/fFCrX5mtz8D
MOQmmu6269VH2X2kTR0RCyDCDv2YcK1sVbUtGqS2mAmck9Mq1O9lAQa/OraLI2Hv
5PFBFlBY1mdFyH28vvA4lwCfjHT7z0+J0RR+YdtHp9cFFWQMhuKYY9VOvm4/1ufe
Eo22ZfIe03AOOIl+iISw/zB06DmlemfXMUVEfaDMbtGCerR599FEY+nnD1S/5pDe
CvrdPdU7f6g8V6ZSYdwspzlSd9HRqb5KJBT0G4bhsP65CeAqXh2cKdD3u0KHLH3t
9eGS7j45Hr3QEKbirkU0Lg+GiTU49OL6bz9SsGDtLllX7UwGpNFKPu6Gzpf/UYlT
TnUs/sefC+nTPulP20Amp5bE1IskbTKhRyszuoVBuqwExDciuCiucpgXUepKtkFs
ZQyGfAzzFBrt1rbrbsHQlasK0U8h7xgpsCxN9rJF3iDTkcaUG/sFGyjENfEHAkFE
o/cjjcGhTMATd9bINs4mdvxzYoKr38Jg8UltjZt6HRZ8oP2Z+KNmsWvDuYifGMaN
iZgVFKM97Jff+rDZwXuI6yEyTUBZJk/YDwyYjDAVd+xp0xcjD9LIl9xUEZr07zvJ
KuwSYQSO3vgWaqNtvKEd3EKhjZ3L93K5aZOwMBEJG7PR4YY+DHfJ+QvklybAtXSl
HJYgco6gYUPeKrexpXXqe4QeyOdykn3rTLBKSEVDUW/LnNWhet6P/J2CSms3IhaJ
8mAeWHCZLXyYjr4CHKEwXwNiNB8864pFBERKxM/MWFwN+Q/J6G9NpiMWvqtjVx12
GU++VTtx2uzjBmuUB9Ty6c1hizHLj+UYMF9QmFfMi1Pl/iU4oOksGw0gUpw9i1yo
nBwyC8WFSEmJfUf/wi8bn1u4y16paxlK3bqtplIsSTS33bY/ZSDVQ1sR2JVOOpkl
xMRKOKfAjYrvI7tiY8Tx5u0d99HNN3RWf6p0eV8ErXnuGHmIK718hiIfS5yMz0Nt
ReUddt59j1AwNnjTL9GC3xc8fSNWPTGUR8UQfgoNTcN0SEdeHPj40B+bl0CGm8Vo
zZ49OV9xK2m76l7CFM3rjA5+ls8fpBMsvCdIooD2zRU1r8aWm8Jh+wrwrk0Jn9Fq
oay1c6i5hn2cxtJ61BH3iTnUgqamTmLuOvSaaOBre+iqb+aEpkcysG5sKEzY75w2
i0lrUFbmAxJLOef7fA1cMdpnX7jO8A4jF+7Bt7JKNOcSF+hdsyCbTKl5AbOAjxaQ
RYKJxP+dUKCwWxyCXMtr+H3NMd4NJse9L7uGKTjsUKBNtYVQrtGz1+goS5oYUX1G
plSStxcGBwZkcdhA/jaEAt13wEAVVYeN5CDlztKOEZZjhHVaITHIzqgKss57vz2i
IYCKSzvTp7ExhGj02aKJMjyUaP19mKzPXGIJpcSwhQwJzgC7ma21kOvAnoELQiQa
7uTYqDOEh0fRCVLfCacrBvBNiPu21RoxHbsRHmkdp+HfZA+qMGmkFHZK+Hkg7lTp
hJrvOpgGPfc34gQlwugCtmwpxi6CqpQ62dMPLNAfnypi8HNAyvJ4+L5pIH14cFHP
rQ9HA7/jizUekxdktXSMT9xsXx6IK506rNPsocKX5Wym/r2IqtwWAWgmp49ve5kd
Jz4TWa+Hl0sCiRwhydhzQTXYTEFaqh9E9BmwvxqrKSw4v6ZI3EW0DZeev1QOojOD
Hpp+0gKAkgx5VH489ptDNAAV3JQOngKqm+ZMNyiqAv5gdEOOVSBYdlXwgKueRMpC
he3JAWgOZVjQLzB/JIE9MKHfDDWG44vxNFiRhVZ11si+jQTBFEPBFEOHU7GmJ1fi
abk2TDerJYmaIBGrIwSROYoUSpunFTOayBREK9p19MDs838rg0v5qbW8VhbKvJkO
JdyuFCH9TAsBsa+32ZGU3l/I2GsSsYxeBcKS9t7vzEjZaRs0UDstSlD8rvLZyt9M
QXLmTgi7aOkCVNHSCUd+KWA6D8hesSAH6yG4aKAm8OBYQ9jCGrrMwt7pCdY6VEWL
dh3MSnV32IeRBH42Siis58Oiil7xleA7t1LD/LGHrc50hXG0oqgaFajBBusQmqNX
h1fUpSYPsAz646QBpTA91dR+patKDPlJz0KQrUvk4iE5yhk+bwZxo4pAReDDmjMX
HZxYegplaM7LBWmhPOsgdqWWZ/CJ5s/FY9Eoy2UhRN0wIxJQykrkxlV8ZIuBLUTH
LPskBijAlV0MkjMKv1Ln4UEAHSw7EyBp7PH9myRcd4tszALB8Yi0Uj6gXEeFZtV1
yVvwLWqW8KpudHTNcjft/QEql4iuAfyFMSzAJmcBIAF1FNSxBI+Kg69DIlsHLxy/
F34CV4SpsxQMNjpTrqAd4obIVlWmaZuK5Ug2Bw9XxO2U60i9Iw0vNIsQwgNNrcca
VYzDvsQHueB2DG77r1qaaNFco0eqlJFoT8uyvDwLigh+/0YqaKsTbPiqUXHKWrXH
skhEdpwonTYNQM5E3a8Z2XYiOXsMZPIzAo1vpmUGRVYPx9w9ueVNkmd6n0Vhx9hM
ylUrZ+IC55NIlFYajYyfUefeFHo+3qFmIiXDkot8wYf+einmKeSXTB1/kSAgE7yu
/DPGp+rYl4mnprNiKpK9MEswoC72aWPyM70Bsbu2HndykdfHFFxdHsUblz6rdxLk
HW2154hndoipK45k4V2+zXrAlvFKlE0Yfk4BoUpogVWcYrPdTckRVRDLvFIIIs2+
iHSCHU260KPE+tRYW3Q6t78PSl95ZlIRZVM9CcjBKIVEktYU2dXQ10Gs7zSuhEuH
wOHGTdLAAPEhWUJ/9PBlpLcR/M6BFiMI4ky3Mp9eu4UjqV5EzdXYJ69KiSOfLMZI
5CXP7MfnakrpL6RWHntAxZ6QDIEIMOwTZFkpQt3TM1AmBPnTzr8oPorFS2TaOkU1
SNzqifqymuT7reLuz5tSdRILCP6hLA8FnIcQ9d2spggj7CYhb/Fcgk94pXKg9tX9
ejVkdHpqH1bREikuDWtGql0OK2cCX9esdEAqnjc+gSBU80UloYzOHldkjMBViIJ1
+1r7rgetUC9/0C46Ho/L+QPmQBgMC1AvWUbTx8hWQPBCrpnJltI/HuT/Gbit/P66
4Nv9vY4MdWDdMwtEIZKIutoO9XSTQyL1ECYA2JYC4VhIFBTxXTOLAiY5vk8BmkaO
7imaypmie2NGaGTYFxTCiT+Ljs/hkA9UlLbBSLwt3wtPt9SbwmrLLoYgkw1C5cOm
qInfuQGTEHgBt2yezuWmp1GLB8FNGU1UtNjmeJ0UdGkGOWvyEGXcatnAc6bdiwk0
zpCYRKWzHT49jTk0ublXNS8Mu0BfWJpH9FcZHdPNIL6LwrJDLNOqgXQ2J26EtyzZ
vBBDKWemJ+YxysP09/e51ayEM6j9HrTxRqDxZ2LcAX28U6/VhUsp2x1mE+drsC8M
rKxSoXyVEqWk9PEtKn4z1HuAY8QYc1xWgd2/gSSCB/8cqmRECQ8J86ylSojT5ClZ
jbygLXmyqoklXWcJFdGno7cjYC1yXy8kaCQ16Iwe5Jc9O7SH5EqsZRc0OBMhoEEF
oRrSBP8DpxQ8B0mqMKqNxT58EcEZ7xDobge3dz/u2rTU0Cug2lwx70EaIxjataDk
oHJoxVKKB84Hwd7FhRjEoMdZ4mwXEh55gulMxouHZn9YeZoVkHWlPu5d+hHeID7j
lEfkow5jZ3HkP1Xk/bijHjm5bhpeKXM1QmWfs21kVrHW+3uYXhxYpSrNUJQZjUBg
sQLi4zNbBker4j7/FOaM8QFS92296yFPMTB7Xwyw/7ZGTzsi+UggPJ2/DLdcaV2N
Ezcf9KrX28o6vMWp/WVB6cDKsChdz+Ie5uvyNY3CMsP8VhRbraW+Yk82o6NF4cAl
oLrUjMJPRJ497FMlz2triAILp5g1FNDqN677tZXiX3slmsjzdq+dWimx+nHkwumL
Nms3VNr0uao3sRZ6XYMQns+PuOVBdhIQp930PCocxU83QwTqIwLNyXoM83I8oWzK
eJyH0ADO7yPH+Ghccni945fcxIoRN6wcOAqAXUyEQ0FEgGRMzSWcdbdDYRQoXXnW
bdIgyQPgSWUldMOSJYjPcvbJfsM77jRFi/eZCTwnRRal0Kdq61DE/xbufhcdcb2u
AxRTIcGGQVUXBR4AY7PXS5zL7qS5C1ZMfkVjh4cqIq9hXwnfAGg8cESj98Ykz8Gn
LGvc2H814cfCA4VgJl2FpPDbqVhyTWeU6ns9dcYi87Cflhb8k+PsrBrQ5ul2KZAP
BNHez1W59p7tzo9o0/yNBxvtwYyvUNHSg4vkNpsuKylX6dOX4+5MwFmz7fqSa3LY
N7eqk52+0nMSM5mjp9K4Qgn+cTRFdafmGiImQYDaQTvCiiMMkJVHtnPOMe75Kmjd
K123XqOvMSVF2UbKW8JkPBDFfsPncCg8EKRRtnG4Rc9T/ibarDg6nCxU/BbUrrBs
85q4adiSoa2uS0gss7xEUFIae/2yy9XhwjsOE5gB5sjz1f/20ieABP/bfMfYVVR2
e2LC1yjlqurfxpTcxRAzm4rDF0ntFaYpSn/lrqX044GXtAbVO+aCho3hXrDsFtwS
Sh4WqvAjUITrbGFQeTVXMd5bX1n5OXYuNKtTgvtCqVQ=
`protect END_PROTECTED
