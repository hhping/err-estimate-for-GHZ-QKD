`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTgK28BhHsMfQfCm+KgZ7/v6V9RfQq6JGeKoNcqfiW/acJuV+On/xlRSQYtNnXo5
c6hzYE4Cf+Rs8LGNkCPVM6NHzl7xokZgvEwwl0ohEPk4EOSc4ayJmSzTIt8PdHk1
7hNX+y9GdnuBEit34eIzHaFTHkp/zy4Wuly0l8vE3znicCDrJ72psA6HqTsw1IiW
I13F82a9W5ijoq5emV+E9ZEkxLCZ/YGJChLKj61vFel2pIU3KEr78WXUkUAjyoOR
7b7qvh5wWQFVx0BVEh5NHhWsEWpe/0EYz5cZxzmU3zaa4wHPqx1P7opD+tDYyj91
7l4zFmiwjsrxg6jMpR089kWD9irwXYcOyycIfDRdLzKI8Xt7eV05ecd8EWpgqyAq
oMBhBSAzjqbPb0QIrlTAhkCP04/lLytMr89pKb+48mqQABSUIFaAZODD299V3B1e
TrWM+ahouebaEoIIwVU9emsm/4yN1UVOYoPVSo10GBscGJkMFglA9CzyK69MCFve
facU5Hnuo/JP9jHkZfiU52P4UF8HzrL/L5zcPs4QMagSCfdL5gN4TO0sOMhZB+d5
SiGrqgJhjL6nXNMj3CXSgkR5K/mI91D7WXNBJXl1ru1TbO+tEp7NJbIym83VI3ri
Qd9TIJTL9bPP5I1JQn4ozKEkY3UqqjxH740dgYRzGjPhtdb9gpDzeC9MhRJ+X0uS
qrPMxem5UBl3aoa0rC0kxX97JKWBK1heoeXDXTqJe+E=
`protect END_PROTECTED
