`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkJZYi4MjBqoJnNAIMAI/aKOfaUyrbBIL2Xk7QTKoyylMOBjWhAuFYZ0o7sSiNfI
LtIZput9l/wIu6tt9W6I708D7Y50vUrWxxonA2zMbF+MOQrIxx/caZ+3ivO7Jsfa
D5/b5PqmBSUoDjyC66Q4bICBLI4Gt+cLcBynZdEyQx3adDDXVpEbarLE5L6D+McC
Tq+VJGyqlNgiChqFoyNsK1iabgbFViGLfgVrlwGo4ioOIgftJOXGB415ISNHSJTJ
wWCP8vESHGl7CT+2YzkGQHuc2PByeNerzzKoFXdzycbsr8p9dtw/cTTV8RQjoyEV
TAEtXkbxtz6P4rixBBNN5sa7vFPm3jt+ezs1ADnMWApjNfv8pnhFvIC/cE2/a6Fx
6FgkbWPJdj+LceuKV2RnLTKbOexmXWTKr5SUrX2Zya6Dc0oDTGoUMsDWxv531iCe
HxVon2GuKaX7ulbsKl35n4tufq2Tow3nXvyDJ1Ec5AqncnyQYF6R1jWDSxpTyqmZ
/5YzS92E+6ggz7rDWIWZFPm3jKkYz1Y8/7gEtMfpevpzqhyFXaK4MgOz7rTlRBwH
yqH9OVGlQx4uD3ioxf07QOhlfSekG+mw1488LdOA3a1Q8EUR9xT4iP1uxewL59b2
zBQVbxF1zVOWWWH27TWU1wffuuzTpzrauJM8urWOK9gnkjfBO5Y5AzxeRzqmO63E
yUuadeP+MYxhiQPkfsElnUm76z+6YGVAnhvK/k0eZFLkQ5gPE1lnoT8t36346wlZ
QKIqXwIBGWGWThZfbEYLq+l39YcUkJdkENwYOojPalXk0J3+QnDRNyi9UURyafvA
xrbDc/ZYQliXeTMIieawNDErJm+Z9Z69cMqcmcRMj7ou1JCrgDHK761lhlDK9yKE
JYfWCXmMRWYujB6DSf39qjAl/QRZU+2kU0ItuV+48QG3ajeMW9Bwwrpbjk6I3zuU
CAyqBuwrcK45Q963YnyMWIPTx8jY4DEV17PJ8ilsYlIeRZvGp6BcYGU4EsPxdw9A
IXPg0tyXdAhdLvg7Ufjq9VAotPW6QoIttqzqACf2ZDYyGEO6bZgYA96Xn/bwh1Zi
f1wBDBWPBg98kkttlgAII+MVBbCzLneNVi7T1SmXYJfg9iKdUPG7FeDT4Wa6vRaR
NHMkD04htFG37pFgDlyjCqVsZeTdA+hZ6hFMSf40//SMFR0d3Ygis2VZXYUAVDS/
STUw3O6G+mEIKCaoXtOFjv/rO4+0uQNq5vx5tCp1pfO1BcdPnoSn4fnTNAEVKuAD
sh8SdTTjYv5i0EpftfCI1LKLey8xgnytR1kSdFeeFHZmekOqjkxLakA4diqtKjJq
55wFkgdCoZ92xW8c0//rTJ8zMVe9T5RCqnb0ihlpki0D3rpwVyHhmYR8tTvojZjl
b98gUfsCh20yDtKLAszcFEkIbtwWMscOMlmHmUy8SH2zjxYtkZgbErLFTVaBt7CS
jwohHADLl0I+L95hWEM5EDYRbKoJu9dQhiCgofS+gJV89Kk6fIP4fKFoIRxuqGxC
R70YYSQd5RcgbO9t+GXB7IV7K8Q6hUEGSZx4bNBtkZRmYV97hcW6npScffm0zjaK
vgxP1u9nUO1Xrl0AoOfZNK56ZpGTsBjNgzTaVoMMEhDEIrMii8wJQmwPbdqass01
VuuPcJ2GtkTiLl9dEI/c4uAPJnSm6FQHsjNqkOP54HYQ0IZZ+ytLNZ13HpukpbVl
Amrt8kwiOlvjMxUCWAUTr97PITt6u1S3VLyIYrVXYnf5FKA4khb6OfrXzkRMBqgO
KnZJt5veIOUnYm/jhKXO48RCR/N2olTF+KXvIGbFTvOpC7f54YTq4KNVlP+BS06z
2UpgW2srKnNBdoznF889WK2tjtxZ48Dv8r6tLHn3Z9u8d97Nf+lwTg+iydjOFqVj
pDv7J91odeyJHUnux0tKHOVUjiepDi8kvGIyfGbAr0rSbQSU2fLnMWIBUVMwSk/B
Aa1FNtAONtmwvzxovVTq7s8/SFUfsCZVqdmZtSNdwOzSxiNW4aT7VZORizrrgIfa
5kTWj5M2TVGbZThzNcJr+7bJ0alSxUrPD/gu0h2VUMrArgqtRfa9mhS3jhPHjo88
JrC7/NI3RC4nQSzG9+h7CIbRT0Q/LOGS8QpuIuXAyrxSpHLREYR0EMS6I5tHzCco
EnBlaQJ546kYe5vfsIRTjhJZt50ppKFTZOldmg4hkhqqDvhPO0npQaMdpFAWWGMh
9/PIgSF5wbLlEr5qoQIxdtdLwxxgGLa3dqzpn85simQbv8vifvZuDqv5B4DiLAV+
0CC8CWvqsYc8nAYq4pdm8ZRTVP70Aje02+L5uaanA6wEsi+PRmtlA6aQo98GP1dA
JHwTBxI8RKhGZdwxmck3OfiG4sVfCeMs9CGt2aUP6IU6WQ6Vq/M737owoVR8ImnN
nw9+x/CO8d0URxH1wb67uUcjkQKVQoIppt3LNrFhfu4Fagn6kuvTY+wb1+ibW0py
67kZOJnMS+99NeCRe6l5KFWo3ymnFiwApQ1uBjdWqvGRc9yey+LGtFAGGUfFaqzf
X6zuBBLw/iGMvEp6wwE8byQ7lVz+5mYtst6G9m3qzEdQ7xTWt8+5UzGMTioPfjJd
S+1AcSwJKP2WxAoCUVsxsSASsZalSbkbNnqMy12+cK0Hjuvvq3W5tF8Fqjk4V4+Q
HADejDH8f5NbbeRzkRodPf+ltQMM2+oiIVDQlrxVbnf95mHMf5RJ4VT3h4iK3ULh
g0lqKVINt0wh1h3nlOSRNLKfv7ZjuCR4WIz+Q0Nj58f2iPeUgcrDASu6O2uOGjRs
Gb8odGwNat6vTP2EBrZQsGgPdVhbCmMRLTpH3TJsuJZD5fbAeBrIGOl16IoKIzrQ
8zTYVvLSIunvwtdzf8jJ3X3yG1GlwsNiy75Zzj3LwBWz5wPE7P+4OtlLEQCK7wiN
iL79Hh2LTpYWsxEH1aZv3ZtZGBtAo1JCoNJ/AnYQgiOdkkeANW48HsrqtaSu2HsM
LL+NPoYoPCLlA8GtwJCrSwres/hKFcBzQ8QFuQj7Hycs+O0n1P5qqmTWQWlZJeKh
BCkQrPKak/cJVm1PtTjyz+t/8dkZP7rMkDxtej+/gMVnT+XaeJjVtcStc/hqXUkr
HWJT38swtGizABVeOaMWIS17QTkmY5+OYYUdj+Utj3n+ug7SnleLwUsLDiWFQ1Op
faT89iEsdtnkxxBIyjQ/0h12wDBkHm3G1DtB+uXnoJ9P/M1zdbiDbtDAYOVnFZeE
q54steCjPtogbOxruJZLeHpA+uiDW3O14ZgAnwo8Z6LykiyYsaHG6xU7iaGfK08q
8pelAf7fZAtY69sW0pj+QWQnPBDETVp+ITNDSX34CwhWgV52iYhLFST1H3wYHLor
GDjwHwDBBiLeyd//uCgnYYRLXN4es9LKu2qyWlcRCOn7pj52txUHpzzOYfHaLF1X
SWGkhFPvVJEYYD+tALgRFsPkMkHHRUpVpjT3r2xnCUj+RyxSc2XQB339y8DzfsQH
qodhuDCi87FffQneiDiC03njmky4ZAnRnWT40JslfvP9wmiuLn4JmUmNlc55WY/D
1avVd36+SLBnSFbHO1Sf60hN3UVy+I4P4eIqo7eoVOFBpDXvgGgH4SmQ9Y3FoSZ7
lsT+u+o3OgeMKXz0j7lxVvHabBiyzSEbX+cwP4A2NVJ8TE66X0TClTwXtyhUVkCz
DAkNqsdUPjN/R+Cu4WwFLgaD1848h/bPpGK7V2E+5lWGDe3O+q/U68Bn1prTBA2M
PAa98CDPR11KWgWDSlXbaMnLWsSiWzjDG4ngI67h0aPdRNQVzfuJkY+QVcQVvpdo
pcdkqUh4lb/l2uKryZ/Jx8s641PF9O5qWh/Ca0kw2VBKumR7WlDcTKMMXFTS2/5n
kUkEa2lDQw2Q0ykTet9n6vtg1GW8PH58DH5LTwnMv7rv1HakHBXFkH2PX7DBhBCr
iMqNYNca+PZk05Eu9fvBxh9jsGFKQc/SdjsTNGJG0I4oIr99zGat7IR/pmBI493k
sO3VhZZdp7pHZvsYUoThsqM6w7/8DW3LCxkTfQD2Cso8/40VNCZRwU7kUJePNaT9
9W2ZoOEL3jgd64kB+hHsgSjZ5brfXSugTLDbyDVjRVRbzRpN1f++jDDtOTDfrUSA
yvbz8s9V7/Vy1N45v2WP6b7JuwolGakVKYq7Tg9spxiWPWyrXXZvmkEN+5m8oD9t
mjX+JeTOFTt4YOX7DHyDQaHaAAcnI4Gs0iBNYuUHsqAbXyymwGUOQ71jCx0HbzzJ
L0/lfyBeAOYK83bjNTr+JeSkyR6UAVHa53fx+JpZKfK4+fc1GgAUfefbYd3N8RWY
Ri5fn+YQKbFD0NuGq9C61ZJBbWOKCxPVD9BpSuH8UZtrUc+4Ur5KVXr5ZoXC1Ke0
F0lWP1SFi0rxX7VxoYKHlKWQk8ZfEv6MmyW5d5sgVHsnWB8hzoWkDy0XIEhvgNPh
DATNvw3vCc0dEVItY8m9601Qul1omlWROvq4s44O3HPF9QNT7UHdnH+aNk6zO79Y
N2HdEBOhnsPXZfmlhuRfwIC30Jr8LbqCTVz/Vk92FBGz6vO4O89/DNBWWpXDdxYg
O3g63ix6tGnJ3szGXNKu6CxPBzf2ZgRDf1qKMPf7LJA7rSzuJPAXjBaLJzcDH7j4
l0ZKSCNKgNHJQbJS9PeolN0cabOoG7ra+RheHkUhelOvFUd52v263maPJCvVGRYg
zgMOIVxSz5fqb11FN5j33ejd+jB6Ppx7mYuAgbuqFSdTDMASyDQVBXPcuTlq3z8f
rhTGgx+pyIiFDWqJzr2gjfAvgiP/ceixcfn2p5c5E/fjFKujOA2ZuJVELr178nhB
r2OVFzjILzPjRIZa32Xl89hnYIpM3LA0TR8tadJjuQpknF+W/PjHSmv8snuPDi/z
wDhnvVn3QGCCQPpXuItUS3lE19JtiXRdSEcRuOFbLaAlsFDzzxj0xjQribMEub07
H6vd2V3LwftlT2EJpJAvchnWv2GBPAJkGICCSl3pW1JoB9NmA1OtSzWEhyJZvmVj
1Kozcue/nejQZ96XfIYkNGvfTY5SxPVfVmgJHjj2FTNIHdP8qr2FgxFfByPB5Eo7
guClby7Wg3yJLoLs62EFuvAfOSyAipzE9aonhzkhvWW9zEBPnvgt2m+NpScJM/W7
nfzvGj47Yk5QNV8NqiKl946w1pWC1/5CFl5QnUfEWhUJ/DLDzyTo5Mw2woAFccOr
LF+wzpbhBuNne6y1i+2qdVFUY8Yr1AHE21pUnU7U6RzkkYE+7C2NlIX1VI6loY26
eoBwV89QO0co1aM+drUxRnm91jQt8QidJuz35Ih1XUekSUITasUy19HVhbr1ZuC8
JCozHfN1F2aNiKzji+o50gnzIl/yRiHaHor3o7qGaUzNwnZqkkhr7RYWJqy0lfq7
KRaQYPBYwP/e/rlcItYk0aRw0lKcACEGS+TF5F7E3l/CQBlDjwWr20pSltD/Hu22
5/hG3L7sEgI9YDe52jaJ8JzDXJ5EfNilJJQBwlHRHWHoXbAyJ+Pcgy9GecSNJr3t
ySieyW96nVuQigk59qRgmFuREO6hJ/0OyDoc2ro4jQlIqpBhlU9kcW+CZzwxci1i
WoUmZU0rteVAsA3qsP3PsyyM5W5zd/QyE5GjZrCcgKY14KEcDFlbbTnYGb72lvNL
c0ehptpMa0Y5p/1JK/OpFSfcrgzsUFgU/NlBk2ShmOghWlVr4bJfQcFae43LRtrl
6iAmkQnuX+1EGa//B6WF/sMUr9uvoVNpsvQXmgow6pt5IJpqgU55fuwxFid3dBNb
B8E9rWvC4bqnlGtc40ll4Nn7eqpbQDZ5yNiJ9gYR99JV6NJw07z98qlo697nRNI3
Jdj6Lz7f/sbDmsN1BiOPmfW9sqbO6nsXD2CVEFk8zhdjXDuRtUg1nAMtlsL4lQ2F
kqgvqndlTv4tLe4o++/lOXXUVlav9JY6mecEHhD8o3Z9egaRD1sslEnoqEfVpn7D
S7pemZzF/T9Gfq93dsRO98iqzDghl0SDQKA8+E0JoC/LbVIpqQq/nAe757QTjZ4n
dr0xBOPlYRtV/073skalAtcIRq09grn1jx0qtjs0ieR8PCcHdaeQNXre17vxhhLA
d4JS0zYUa6R1glwRiELH1LKUda8Ii8R/OhVvQPEdWqCz1pU2o4ypV2/FyO/Nm+rk
QmYUrf5YvyLZak3sAa81OZ5O6RxXkqrDCqiLV60BaJ/q/atoI73nf8mIIcK1wC0m
/NJMM/tuSdv66iJ6bs4djsTqMYXXl2KDj+E/OAfJMivShJouWIbh8V2hRhynis4o
67KxxEAgLlY4NrmjG+T6MndeMeNWqizRBE3zn3bLIqYvblszymC1qZHKC7lzwKNo
mk02M5BbRR0di2PMXqfN+pUaiCpWVt6y/3rH5YDe8WfA9gsC7YjqzDTD0xiHMpaD
M7G83tEODTxIukqQU6ZQDHKyVsY4gM7z+LODgIoLA91KFoT32xDwULNTofJebS64
pB++rR6qLUn9fF+wn7tl8PCaTHZWoXyLynZwm5yOHALkBJll5lgCaD/agm1GpnHS
SERmJqQJAqJP+eAPJ8ZfgfpRLXLIi/cYUSJTdZa7mGGIgSIfOV1GtvR3QReNj3rz
s2m86XShDLUhD0PxW2U1hhrSW7tF26IIBryEEE0jn+Ud4NzfkP7mOJeBcQoDfTJE
pvoa/sIqFv1EwCu6rU/9Qw==
`protect END_PROTECTED
