`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hBmokc4I9Z3zinDWbNqFDANSDizT8eSYHV8BB8i1bWh/RFHfaOUdX8El2Y5EIb5g
2oIqQ7dBNJJyo16O4huGwOpRncDD4WNU5sK4Q3Ju0wKOfdhdWfi+TE0niAAjE7Jl
Y3+7xeSX5LnSZB060cJZG8gANr9SERrKRuoeZE08MqgEj3j/GcfFVjkofNsFgV05
0gS6N1TXbm1kZcr8WWROnR8TFwmYzsZaPJRxaH51SwEeeBrUcW6fiRHGqLyzF0Wn
EnAdq8CNS3E6lYQ2JPTRbCGZh4UA9jzGXdMiqIf5kW37WbnOMjQDrpgXVh1q235L
qANNXnqx0pSRi2BWIjo6c0F2dUYvtXhYHUi5mYVfz7VmNib9eWazL/A1qnRfkAqD
kdRUqBdybwJ6rIdJAVCIv91abKUN2dsnAGuXuNRLqXZXFBrJ227W8QDyPewujuQO
iWj9X7vgTHnaZLqpecXybjbUIkWGiLsDAeBodurm8owoFfdQ7Jd8J9KXmcyPra4f
hR5WSf+QL0Rr2xvig8h6GFtgnCVNGgxlpot2kBQfOu9ORvQTPYJwj4gvbzhUiIlA
K9LbrnrmR0SI8lTId2ACSkd8mGCdDAwLhO+ZH0NzQmR2Tzq0LiGNw1934Tbpyait
s+zsTrEVHakB2xrf/3oU9ETLq6g0TsFvfnTdtpv+fq0ZkfGzzUTmqiaFN3hFPN3j
L9+F1buJXPExNJA3HubZZu6cArDF1aPlUKJdcFm8HK+QUa736IkL2WturmHu1ADJ
AnoE6CVXTCQigKM06o4iIc1pW2h130iMG3Vk3tRN18G8QkMhOP4EGDaQbBLrMZB7
qiVj7o22tdw+Hwl8Ncp3bskT//NNMgiarvQ2a5sH2JdZHnfxR+jQJNj0Y6oZ0Sf6
b5g0KTW7mwej7NSt7NTPwwEJ2YuGAe6jW0Hnjp0UYjyYBFKv/3oGLqR3AwWH04fG
GCAA1UGKTHic+oBOCBhBxicu1qVnQOd08cmKq7vOiBUX8NJDDaAZ0RH9nMODE6uh
q7L+RFYiWCpX+Yzgl9GtOSnnzk5BR49EnO19C0pw5O+maDh57+KmHqG2XC8WTNMV
4wICjMbN8nhxrsuhWBbr+Z0eu9AbaaDZUEoymj9iaJ7oupqNBTZ+UvcXMBqI5R/l
3/4++PuK4QI1Cq/rsUoLpAAcPfpPSiqHI+0lFoD10JDnGXcOf/KhlUN/SoX4Qb2u
cI7vXiV5Oh4/Zy3cy2efqBdAEDLzXs5FnkuqXF+uMbGhp6q3WPV+GU0PI7yy8eEj
XVdf+RsoTf4fdeo1qCAhN3rgfCmO9QeRCVBtirT3hi3yMfaVks40Vo/T/4HPq75a
dDkAR2ZbJqhtOuKKQpZ6CfIbxwLDKOZRsUujPxO3ieSkwLHHBhvYuMOqqmldmrgF
9kFn9oBVkBRvO5cGUSrBtAeqXbnxsr9sibac+UpffWomLL4sn6SvpX0z3z1Sm2HT
MlgRvLWdMio5FB0whTLg6z4u8kZnc8lIAp4edpVPfrIx+o5q6o5LdZ8s0G0c77FX
NLaG3eAP7aXSe8TRXRLyQVtBcM99K4f1uLnzvrIWnJUQHJ6iTzdlhCctZGNnRZ6Q
oSPNJ5lk4eGhKmdCCUjwo51JqBWrdGwqrpzo54BNYbim/KYSD9V6OprmuKCTLPX4
Vp0ir/ct9G6uaomUaQ6REeqcZnghp/omJmmFb+3AAKPpiA4i+OJr+rIOpP7Muw9s
dONtrt2Mrdsv5H/3AQjjiqpBxiMM6URj5ifoDrfIHuig4KYVOulUKnEO6cq7n3d/
Jf6RleIKUfPV2pEq/gqQydnViFJVLtihnY0obAuSsb2E7eoxoD3ujdLh/mCoF/YA
jBYpiPDpQsgKCfzulVDNH7HCmlv/+rXPbFFSTPaxzKuY9FJ1amBx7z6SGr6h9c9H
6BXpHZAFejxeUZ4ahBGpfFQA+6N2YeLjn3roeaZEpMw=
`protect END_PROTECTED
