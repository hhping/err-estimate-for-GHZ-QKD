`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqHR0ScHDp7X+amBm1ekY6wrSdxCG3TnPpxEI3y+ZSzagovSGBtvfjL38aL3d5US
ssyWwHSHO3X6UhPRwcexKBAunMLebmg238k/p4w+b08ihe75DeDMW0HfMd33LthU
1+YjfA3PMvI6ekXF08MLQAN4pbI/lx3/xTZsWGyi2AR/xBOLJTlF9YEpWmJkpiOF
l4m0Pcyne5s5BxpoXdmAAAm2EaEaueXHAstS97is1ykIKuo9n4EpMHvCpzJJ9Rv9
coIZfAt3XSNDzdrgelyDOf+c6zeBB8j0P6wlueYpwzD/jMuCGABGbILpQw1rPldi
MbxZ+P0nSbV+7nFXLHEuRwrYYyFFUKCsoA1UO0K9IO+v87hcQ81PClsDn5tIBWn5
4EoOPV4ypIuUA0P+KLbsxgaDzwi4SphnucZD4kCL1uziChqF5677Kvr6B8+TeX/w
gsg2us5UlnubsGYdul6pBwtMgQJzkU/PC3nCXRJ+rEIpDevueptvWChQ2hErGJmf
phxAaaf6JJQQdsrot5aTpI1f/ieQJlvgRVhtJbKsb+6pv2bmhkd57xV4Bes9iKPu
YEik28Gsnr7Q/XpMNKW65Yqb3e9UOEmBtTBIdPiBJdtfY0z+fuUCu9bmnbkkZWW3
27Yu11KU5g1jGso2xlEOU2jzIoiz5RKimJskxQaf65nChL4Q/L1Fq7OSQRgSpw7l
0ZzJeMuiMqLpgnI9BL3sRuUbz9DHgHY/TtQxXyN1I3qv1KFedPwA0w8XkQ4OKNbJ
Ogx2vz53qBCkmz6tPhMaKnWdHNvsAxEwV59q+oq0h+HJWDWDAWpYB/cugFhD5UQo
6hnTizNGJPztVF2mJnFV6Otw3rTTpIpc3WEdLHxFj8XE4RAZqwWWm1WnSfLFp5hc
l/kjndK0hoqQLQ4pqsXMHczgaLs5wX1HEFqAmEzRs3P6fFl1aHJQda/itG8VL7hE
OUSn4pyInAa+s7ynsroIupNJhUvwp7qmEP06HvpdttBWvr5ESow4krQkOaAZb9rq
DOQTuau8F3+e/XfHBeAacLpubuWixEW72fNK0GZyp8B7qRbHijpAQxgvkjlVi3Km
UUsb+OiK9A8CGAaQtRPSTSYj9Cq0assn8dxydO9i1A/Bhq98M1daN04B7TzU6Rh+
Q1GrlZa3TM9CUpn9tqYkdfaqBuCqHkWYKE4j/Cck3+isnbXJTDe/sjzurehOHi3z
1DFphEj2c6euMK4By23pIIiZ/A2S5LwzlHdAYZgtnjqIPtjOibWaCxnjbjix+p1A
ZAIcwwkUYPomGJcUf+T8Z5xMj1ky75k+raqKZu+PhLpk3ZuZj/lw0u1k0s+SYC3g
DRYRIpv2JuVgwQp5WViOePseulsNJNf4YIbd7OSFRJ7h5TPu3mNNgzVE5A8HIlhp
UlNNw2WB3XvM9K1Of0fmGaxyab4k+t+GcaA0Gf3SdFfCtDX0E/HYh9ws+IXQBuKg
B4xmJufuWlaXTTt0R5poaTa5TeTithb7BpRPTpNAA4iHjYOBWR+UEHS8Dk3f00Of
P52jf5A2oK/IsXAfwJDU4zEiwtCa2Ohwa+CV1K1Pi+uh3nP7I6PcBjpLh6YAZsHh
mbuYHLzpSOOpz+oZlHoZpgmjCufTpw7OcDwvPm0uyalq3mfMOj9P2nbq4Wmcj+mU
eIPzRkp3EoDB9/skwHNOMw==
`protect END_PROTECTED
