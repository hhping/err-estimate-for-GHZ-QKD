`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+f+Z+bCUmIzuKjcgfKhCjCsMjqBw4k1wRPWhhHyDaYtSSTJEVrbUmAzcqhTt5P35
DGsad4wqiz2oHiyx18Upj/SUtmOdcpmwBdhpV2gsQYfp5QnzjD8GP+6w5nlG6wcs
aioqlxH6Z1SNW+YfM7t1oJeZObsxkMQfdwfygNFOksrRlKncn2pJ2DYqcfj5O12k
PFvFrq77GBqzMrWP3TqV+cciCpShocl2F0i035h7PhwuEmSeM4gZ3Qp0Wkd7aZMw
MlFFKt3AgMlNQQv2JaTcCRfMaeM/HCO3fYW31j3mU/F/UIM1fweKtZ9il3JaPGMC
9/9MCX8s4hoCYeWX4nrS8c7SDNc2Srs+XbDkLrKtmlhgNt/XlvaQdmwvVG+EXsNT
i1LDTVl816P91NPFO//cvQak5FnfLuZ8xaz9gvpVf2zbqj53qAbl5uoP9iO8TcGG
URErJyrP2zntmIXAJCDtv+X5uI8C+7npUPI7Y65kgR9Z5STyi/sYKuSLzJTt4F4E
WzTKxWxAqH3Kw9aJ7MaY3b1B+zuSpT0T2Ny9712nn9qsukmUVTvgiwMwDq/Qymnn
`protect END_PROTECTED
