`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rbBI6a1uPXft1Sk20+ATs11ybFKYN0BxIAg/oswETmRndqjs31ryobja6CT+7bqM
B9jM0JBlF/39yho12Xxiy1wfbMWss5Cmb9VaRWJ7Qop3lkahjDlhLO3iBtaR1FNA
dENel+I04VqHhsq5B/Bpr6kJ3eukg3XCo85/kPKX4ghBWVCKgxmaoDC2W1d+kDOS
0z24Un+dnIgn1Rql28N6emHXRQj+nHZs5sCPWRsKr+kGaqPMV/A+t1lUDvsQksKc
pnO0TtMhNHIuTz53T/tFobw+lNjCj5Chshq0z6uTM98IwCCR1jshRruXTVNp/bDW
462aN2HyQ/ZhUNk7IDv1jaXUcDy+Dndys8bBbSbnkPQ63jDmEEEkkHBkVf3M+lNY
jSNiDTdNsaZuHjoMfiJQOcIRqloyzN7SrjVPh/k3r0GIQSU5iBb0Xhj3j07Pmuzz
llxel0hO96M2qEjWLw+GWdDQOLl6TfwwaYgs97o/5rPUuvrYz6ipZBwcJBl7ta3G
p25Y37oYODPRheok98wCbj38h5E7azCKqIdpMudAGT9OgvWD1tHVJytRHESFQ651
3yrEwWNN7UQTrY83cadzE6rkTvEpPm0BZL2C6YMle3mqARJ2vSsO+uNhal7zEBxk
zKA7V6wd9LGX6aX5Olzk5inmIZlRpR+7x59y96MKwRhp37QZuiE9NaKVzlAFL/xx
tK3fw10h7rYV1zyno1QzcMXjSFvJKo4jwJIwcdPIe0k7fMS7HnPPMQN8c7oNY6Nk
zNdW33DPzMd4X1uACJRDOPPUd4qoUe4dAUbscfqXsrZ3mJw1Jlpjc4ETouuBsy2F
GFgcpUbg2cHKCMx62aBFL7AQPGH5eXHXKzSeJsgw+B4qtSAsOQjI+8/LJzhB7yKp
X4aoCG25qNzFsJShe9m+GItE2eDOb50dZ3QOJr6SRtkX7koDsSX9xaFsg/8tEhIs
OqI6yQPmrdqETIYKgkc66flQV7aOl+deSFxlCwRUA/2/j+Upi3mwcm+Eob4HoFPo
5uC3/R6x3UNDbBzz4ScGTJdqMOtt05T5qZMPmWTvLNzzkkg/KdBZDKoCHvR4T1up
00rkHHpno8E5lGRcc9XI94sb2eWS/oELXeCpPjSVYtotyv9R20OSa8rNkULB78GX
/3heZ0vtQItJauNUojrIovtcLIHba2bdqkgAxMHlhHAxuWlilJnrbsi/7I3AEile
0kwkmgqiWxlbZ4CNHEOTvN9G/HF77K8aKt1DzFBTdmql/3/lmXngPHiAHl0tyedw
bU7cJRZj3Cv/s0m1Z+uFCZAz6oy1JP9YGU+ZOxHKi8Ok9bbOkgUepmJRPsENBM1g
D5omAaIUwoAObhqOXIuPtUEQEqKAeq+1gxcY01SYsQDRVPruJoZRymnLamynZJWO
pEZCqHPioA8MlIXZtSASj8m+8b0adFDhp1v5ZJFIiUFbGvKOggm+8U1b3cZJxtjI
v3twcCbj0KjD7lbkMy1sJ5459BLnWGcQR3ARSsRVDbRu7SFdGA7UyjoF3PQNEzQy
rKZ+qheZn2ljQSYgH9reqXypylgBgbct/EGo9PCxq3dmo3ONVgtG0YaJfOSeyZ4/
2mKBpww/nQRFseXMWG6VbY3WGUDtkcqyudsqbsl1rcNm0fuWEo3b1ULG5UWmfLY2
KRlpy/w0YwzABBQ+ItxA8qsmezSMAq47/S/XHQur7KGxG/pFe3BpHq/vKoyfu9/X
SWv5SiLn232svmmqAt73um+/sv0Op69m/6CcLZ+Vdpe7KdWL6RPYXqVS6NMaGfeC
91KLyLXX1ZBWLLCYuev3mKhHHXFkD8dMbmbXUQ8oADxUqQS/Z62iE636B31FFmw2
oAXnr3EBRcQxwAwxsweAW1TwXzpI1vwc790CP0BedKupYTdvOyHO6Rx6W07Vpo8O
VLMB6HJr/FDvOiLWTWdLezo4caYWT/BCSlCRr2FDg8heymhF2F+WJFloYX4vCvo6
g4wjQUjl0I5vyG3uSM7OLtKDfF8e1SDcq71WyHfnCNnuj3kjVqM3M3FCyl8v5fRI
w8ycMv0NrGWZ2vDZzOwqcjqG39gQlwM3LoY7lNTGlQD444PNngoPDaJUZrkFzyNG
i7VhLy59sWEVL4ytP7UMnUt2q/5K3IrPU/cMpmc89VGFZ5ecldcj4V506wOW5Liq
qzMpWzznj6W9COEpeuhrQx56fOqnQgwpBmu91444uYhMqBi5GBs/CRSXqCajhSkH
9IDDM0ffPPblX2QCMNKnRyaqmkEenvXWfSFW4t+BYxkHk6T/lRGw6FtCbiUuTqIZ
VDVvoq4d5UCcr3xA0CtkqFMxdQiW03n49lQGk6MtVN+fuaoOH/LIK2IQxTyZPHge
JmCGdg6Ryyxv7WsGB2NZ3moVvZ97AVJDZCb01vwx3R5rcL9y143H3As9ZERZ0C03
0TCiLScma1MW6bM/C19FaSTR0FQL7OCy5jHCcM9ItwMgElz8pDwA11nnAPkLC1UJ
ynnhh1nUcEiaBA9hq1AbO6ynestSdNNKDKTY0ruj3ErOE64rGZBkA4HeQl2mG1Y/
vrg9gYcRZtQuRspZrzeD2NXRUKKnviREw4AD+RMHGkL6Uqzx2uKSbUgVvZRGlPNQ
OMEbdlTbnB2rXF4mF3ty6kWpqPEnzMmjAwqY1SgqRcOiH55abDOThOECfVZuH5d8
iZsijLcDyAYvdc9aYHsaB47Asr2hlNLlHsK6IH6g39x6W4i2c7wV5l4AoBwxn3B5
6JIFkaSjg0Kqsh2ucQD7Yv5didzqT9VWB5Erf2GYG7vkLRx1y0SMnYCinPRlvlDd
Pe1vXQ6HmKwr1+2TBOm2Y4XGDbixl7Srf8iXFEb1GErfJY539bRWKSrPi9THiMC4
EwS/6jyQ3UHxtMoou4kI7LXnppku4pp2nWtdHtEJRDXK8Cvh+ofFxoXG0NyYTmG6
JkdnCX9govtX8z/FYfi+uyxY4gN+adw+m02gvzP8uv/iSc8PFzB0zicnyOIwPP2O
EZTzXV7Q5o65WfEMjnY6d/XmdVz20m+iHI10vHanhnKMRv2nnPXle+uJVyWWhQcW
Rp93zRKRvf5ODMQp/pYPl7tK+bYAgn3l9t7fJ6zjojhNgsPLMszxMuEnjthBNbji
qe/CVSl363MYpn524jWS8W9w/nSaiBWGLi8k7TsxMvjsdCoy+ntlza6VpBqRi+cQ
`protect END_PROTECTED
