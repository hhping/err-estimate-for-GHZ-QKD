`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTCKrOYwsP8JZe8AuP1pDNsn4jSjqFHW0r6TkvXqOf49KDU8TOgleyuxfwV7Zx9K
c7H6fGFzC4/ZBghtKPkdRo/B5y2qbvg8ypgc3q9ZNNeiqw0qevtV1WVC9qN8OZMl
cuJfqpVVDCmGKX/lASrZJg1WBUG7VJWcNV2Jx4YbENqAiHXmEVZi9pHrXN72gIoh
MbtrcxFniCdSWnYnapqKYcw5Pa7fSsJ/y1UDPoMJPlw7ugC+E9SdzaMJz2UU2Q63
P+Lz5aX0ILgri8LjcACCFCtx16xHyOsy4DJKMYdHn/GlHqtJb1Yw2/HGX4uNxP0R
6zIEjm28OtXwHMTMOtsnxpdlg7chX9iwQCmR0kyEddSW3fY8AgpS+M1QidQ47vaX
rGRzgeeEzEiAR1WvjybLDol9R2RjGToaut8MLskIUO2sTpimn/7uZlLbQemJlqx8
N0CwGVEvwCa9brOJqxy/eoHZE1dj48X2kEnTcU10UCMKQIMRKEGhxdmcl6jpwsUq
BHX8JoiOHsf2VYhtj8cLYBoaBbsH5FtCbOwfP+1TdWuadfQnR1m0Q6rSGjMWG+7o
54iKSerKWs8PZsdbDTkbKh25ncQWh3Mog8e9a6++RA4rBftSM8RU0v89XLAQbbUk
GKIpZJaK8JM5QN2psF9i76w8tptdYPSRoiB9tAZHBolUmxQQro++ScWXX9k6FJkE
o2LPqyrgJPg7EVPYibrQJwGrGICkUVvaZwpuvg0Md0W/ccAg9euOpLsnbvjtX/7E
dXg4RPyYzaSfGpxKl9XrU2v9UCjmEb5Zwbq4cK/2liVs3BKXkSzzgjL+EhDm6IT/
LZ0eqbmoITvu6dWmsFXk5vjopoA7xrl+WA7u8k9Nla19eVF7Pzdn3N6HzQl2NcUu
ORL3zTsoRBzcMX5V2+OmBl4/G2LNaQV4psv0A5yv0ztsuTNXL3jC+PHw2stNEWih
MeVnoeN8Gc77jlIsrFrRJ7Ct/WJdLd39kfyZnafno1SC9K8Y76Hb9S3XW9P4/aKo
25c84o3GGl2CHcKrA26CGFXXED5wNEp+eBrE4X48ND5rS6GckwEEICvgywg4OpQ9
J1qkEeGrW9IU1ln+m+O2ot1z2rX8jT6ewrE7Qyp0FzYs730BgFChNqjEMngb04ra
KHBDXpptcAz+coUDfJpzMgV2z1XqI6vGYMR8BTQx9cW1E7UdRy95AZgt2+1iAeot
fA8W39s+eyydkORO8ItYPeujhdjMNNKWujgb6LgCAzzQ7ObhgwqKPh3Kppkn5XFQ
5hMoVp7XfE4nhDXrgWWI5EvkfXuvIgocNlHujoJ2PXrrL8bTHPXOdexW804lOR64
vGVhADOQGEUCysyoECrj3MBEiuW5l3FGDi7INZInLSgfTUzNEU9WmK5V4Pt2dKM+
SxLdusLf+7U9Ucq2+upl1dTKZjtWV6iWvFhl0EOGJEBA94cCoGDzAl/o/hPByzvU
hPWiaUPBwK9Ii0ZGhpHHl5goTKy1KJIWvqgMPpo+aBYzlLLjRg6cXqYknY5DVHmR
aK1GJh2xLsAuYEX3Arc7S3sZ6+tp+PzLUW4LnK5srjCDIrO8D9++Jtkc53udZI5J
J2r+jod05FDFd1BqwmmuB6Y/FIDGMJZfW+q/iBPg9BEU3MWVGjyCvN9/3TIckFax
bHlyxsWAtwryiVpw1r08dg8o2YBBLtCF0yZIHIU3G/aKGc3IMwXbCFVrIgeiqd1f
8HmG/X7QW/z1CtMnTbve32B/pxmz0XiOzHeZz+qdSueU7FEsmej8bqelOV2VZFsy
EiD5lkcOJ8wmpIdDfjgGzfV+djorXb4pTtugkE6+y2evHc6O2/TX+1qMbqSibFHP
FxQSgemIxDy2qMU5tocIbd6EN2Xf2XwtYY34MIlKjZsefqVIB9CtUQJsc0vwPK/+
bAtUsDqo7XCq0O+1EgTjKPwL3gKkI7TOv3yLpwoytF5fCWoHDj9OzbggRNP9WjgI
hp+gyDd4PGf9Slf1kMlrXjt1Kd9fX31Lu8+Yo3FeisV+sqi7dpxxEpJbLTnwFegP
h0Y2Ye99/fVbicdgux5DUi2ct9Kcz4JFDULCeujuSeuOI41QXpwGjp54lg7szbu3
3yrZGS7w4iniqbA4aXJVKX7NUcfuC6ljNaUs9oI7pnG226myQM9JhLlQ7MpvexRU
+hSs3ih5agnfyyRmV3Hn24zZz0wkopVvyObQnQIr2L6OoA8ybo6nplZPHqKK/WTE
24aRwYpdP+F3u9WLjwSfoHG7OtG7/tV+im03FrDlcdX8eGEW39CrZB4TkaClFReB
16IadLvbVJ913Pue5aSTE6qrVXs9C4idROaUwgFEizC8mLkNQuWNRD0m/elQ/Exi
32pzd1h8nD9EEPaVSieoXqE9LXAgbZoSHcQwEfWu7VahNmQyMgqYTRnLvo0BlfnK
675SG2yRGGhxZW9au+lElk0NVtru4bZA0C82JZ2GXHgQ7UWXEKqb2WnMTJNa4ptL
tMhvRqxstaRfFs44owz6Z5FZr/zRqCmRBY/8YIBxu/ZrEU7RPkm+gIRBMpEBR+5p
nxSPz6uup11Wk4/3MV6kIukVDe+iklhP0nQX6pPeNirQM7qIyBwZkAPbuASOocbR
uei7gYWl61i6HgHOGYT7YLWYHe+EfmEwJU7wLXmcj8vimxX8ISc2rY/tUoaOkOrg
YI83/S/aZXwwo9DNcqf4TeeZlgLLdPADuknLBLwTv7xVyu0FVBFiRXOdKUXcKTK8
YLT/ROBqcV0pmlWJ/7wgHXRtUHwAMuPmV/6sjeTdBIAMR25tLTLl1491SInn4pKT
3WJTuUvlbtGQTP3MCSr45xQ1eaCzYWZfwt+BC41d0rZgYHF2HdNQfV9nFUGXSicd
Pzq6lrLTu5UzvLfBmIOySx/zV/aUcyZUcxo7grWGgOz3La1mzkTbqshM8wLmk7pm
nXxKiXzRjaPH2NfXlzHHj3wAemUyvcW8XPYllsMeHZl/lmtcsJ4PaLgrXCASZPmj
2J75sPpLyJpdcGUQhiLzvGwZuYKfN1Hq+ntfWMbI5KVjjfOG/30KG9BtaCgqrQqY
o2O/cYddnt+pbYxMh9iJ0wQN8yWtlrVrCBBJt0w5AV+72tGMVKqxeq5D/NvkD7Uh
9NVG/Xts7gxekANbg9y0ctbDAv/6Zs+4KwVRmELWB5iZItXzR6h633GMW4v+7f7Z
Igw0xba/dqSmZO4w/SLH7F1ySLZ0yPmcWNhFr+HZlZuw4Mgk4HzAe2/brziaFdY/
vhGRcpo1vqQ58JrwDhVG9Eiq1M7UuFDU0lywRFFfKsZfNItUKCxTpL6WK9BrnGNv
p7SohYRzyq0iZmC+MgWmFi92J+PGIm0Rpd7lIfKrrl+ynh29axPo39pYHOPVpl52
llTl4b8ecCm7lY/Cm5TrveMx1n8HLnWD8LQsxzw3quOr/buItrpw7B1TflP1tMJr
MqjQPVf355Rzw7fD1SveZ6s7hX3mn72W9VAr0mVujG/D8VCl7IzBg9INsvZ/fsGv
+M19/18e4oAv+7oiwO3fkSO9CrRANg/TtBenSkTriSQFE9oXFesk21BRygQPL3cq
qqA2eNCOll9iIYKN+SPgbp7Ly8rZeFluraxArgdfeuqKBEtcJhs8eqf5LUfstd3D
bxoSoAo4TW4Qa6S8W9Y/W26PMqcRHbqrKFcEXaHlRTNwrU0mRWxYbdBrhMLEJerz
uIyak1IBK3f3sToDbfK9YoQ+bhwLWOXifQG9PObcwO5DgutCRlLE+icZklT28WV+
3jPBrbqmIeyWA3NlXmAHRhnyDQS87wKP/G5daPPFk0uEj6Y29ttbibMVGrBImRjl
FgecNXKvin78tVnrRbusiAHOvT00Nxk6pV3pjyk0B0j6ndHdz576QRJUjyFGiBAI
ap945n11zr72JH6EmI1ROBO8oVH0Mkau+TtKmqb8ikf8Hba27Dhg6LWKKgdmLnyf
NQInn31kEL+6Lg+owqRHjuJcjSnSzH3SW5FFPU5wBuG1OTuc+ctiFaxq8F74O8+a
96yQTxM6xpTA47FGQuiKjxTtaAImjyS5Jex2DMGow/dGKBAr4Cn2RXbJ3mIxl/jB
0Oj16ulMyNGMu4r/Ycm4T6YwX9RgoUvjLwy0bfZEg66wvE1FkswnN9VXYyPTSAlk
MZ0KlxB54Uv/IpyMbSHL4Ab0dhrEsoXLSERIYArsJDKX104xFlFdzJT1m3IcVLI5
rAdE1jrXb0HwNDfghzpof2THZpYIkGm+gmTDPGMld8wxheAqJD6EUvJwkfDFn2AT
MejpfzoQm3uLv1ECWYgtPtesFH17N7rNe0hh3imoYgCaTQyPYd9yXDXTiC1vR92Y
826hfAdA0bhxlESgfz6biik3Ee2lAkKHKLgKzWZZEWSyZe53c3oAj/t532cUNBlc
qOmYg8VWFweCxYIEcAfD3POYUzJ/k2vnp7z/urvNAAx4igREgnr987PQ8jvCGvBJ
VYmweC8tFg7mgkdf2we8X5Y4zaonVQ90UxcjXHw1+4drHf2Dl755uKZ0G2TfAksn
ACw4NfaRAlmdK8tMUyPlGA3z7fJ/wTEU6roQpMu0Xwms3UFOmQrkcGLjJFPUs6vJ
ubzGtUPJsYMoTvoOoJP5TNh17XL2SdzjWsfkF3J0JAjmL8f/8X99xXCyVtp/jBaO
mXNt8NGn1vAdCo7OkJRihpMn/ob1LW8OTS4c6cpe8OGI+41b0aBpm1jZEa/DdDUp
b7V3/26IctcezwECZDVXCfr+cm1iYi7wSmb+KT77nSN03u4jYguGMtexZj1C9mrV
fpRHmOrQkFRj1d+hroDi48j40FL+RF8If98Z8g600Mk/m3kJKUXHgvzzUkR2ZFCQ
ig0emfwVa3AXTXsXVKg3pl/L5Ba8A8PXXIdQRuclR55How5uXkv8RsPHwlE7OdB/
8M0kTh84NxWyBPtqngxOE0HvZNDS/27JrWRILxA5ZbTSXLE5wfm+MgBm18qRdBCV
q5sSX6EKJxHTslLzmAqqaY+IU2QlgcZDcmPkFaDR2lksfe7iDUY+nhyXPRNVPLfO
Kcl/RYoYbu9jAghSNXOwJsd8rJHnjHl4NxgodHD4xbLoXvlCR+CdIjAVZxUKuYaq
4reY2oKMAy9JriP3pnJ9c9/I86equDRIWSdLrKrfnk/F4ahLg8MiKfeh/pEtmfSB
2pPtd9nrubBFII7y2HeRDuySExo9EtpD05lKEFvyR1kKKa9/MxpumWcY/nHns5jR
JUGjtPJ+m8Vkef8JZjc7/hpHC83ioNcLD0zA/b2GCe8qjuyAd3R/wZflLOeftaYd
IPquXLVEzKWxTQifvEE1V81sXerx+xmDm1ut2y9YQhdzVc0WHEpjf7aO1Ltbpsku
ii70ltS76yB4dFDZlWTI0rrMbjhlZwaABKE0G5u3abHEhFm0pb/J4ftf74ElytKG
2PIrW9EJ9lX4peN7l1uJ15zWbwDBsdgvqiGlt7AYP9OOfec1MIKCCkpEZD+OPP89
nTvNCG3BVHxS9YK9TwJY4acKUmSxXpAMsNYg3iSDi2uv29FffrSRh4xlnX/VABEl
1ss8NsMMZA1FcbUrXvyZxuaC5pMF1pi28ir15UunfygV2VLWgUmUhcRE4JweMXKw
A5qy8qJaaEn1bvCk/Tj85VTSzc/pn/G9hjaXWGQlB6FclZ7lh890VNb+CX9VCJp0
1OUx3Ujt4Vp7EtubiX4O1cKIT30XNtDlLz4h4NP9WHlqeZ4nEl9VY6DzUIDIsrlQ
TxPZblenA7/TVhZ1JdqjdArmCJWWyqWD8auzHdjOvyyrA8x4rA/PaHOqHCSLTSmb
kiEZBiedvsWGHnxTQJwv1jIA/C3ncRnYtdxR6HHAlk3OPevAluxIKRTBHPtbhvcI
g8A8KW4zEzpa0jt5SZ8xmr88ctc0iLhxGebGnmTVG6qN+bnTHFDZ+AZuCDJ7LDuZ
fNwaLJ6LdrzI8WVkhfhobYxytlkXseJa5Ql4wtBL9fpyuD4nLNWpzaNz7+7RUZD/
hKnpufZ6dTk6fLkR6zKAjPcHApPVOfYN9LI7LJn8lzqXnqNeahAoWGHLTQ3eqc2R
wDXQgp6C4xjpDFV5Yek9tWdZZ8qiHiRoqok4t4RmfKw63V6CHeO29CotbH7jJk2x
GgfMyEQbd/dwBNswLlT+iCwZCTXsjmqYszVNgKGBn+TiGQw4T7f6nkPgjc5IUCbV
XOLXdb1djGaz4ROvajn8pf0kHzvRLYI+cWbPCab3CdliRNlcYGz6roD2EEaOEtNC
3omRoDc8aeWZi4v4TIsZZ/goNPo6cRAnqecdMHsocMN+nS4EEmauOSqFAae9oHgU
rVPNH4Ma+vnqUGWKSojsLVkh6BP++0o6P6P9GXCzhr/KRaCNmOaer/S4/vfsLVEy
fohaX9wa5d5HrctpRgRf8kYms4F7v87utCwAQVJHI0FBtcXMCkzGKHNpPDD4aOTt
2Gy3veHqudCMSB4evrA9u7J7iuD9ULF4V10ZJDd7HXkk6pQ6+Sq9Ql1/HqP0UXVs
62XQtQ98/edC0enN8wROScWrkwLhSZnC967zGc5p/OR1Z05fLWjjHMq2YqnVOq31
kdKLsIjPRdiDcv3eOc23szCWp7JDWZI3sysxSapvpdCXMgLozZfo1u7L90czDIb4
1YIQE+e28ZHB++4LTFYF6l4906Xep1SsSVqMFobuScLmRehbhkxiKgUIcld1M7AZ
9fCefv3l6+rOKlr6lSxxdzHaQD7Pq7ebcYegDoH2GyDgMLRm3dCaOGXw4UrzJmNZ
rKnbVYPAtjQruPTQomYjdNW34CFYjklsb6x51kUlHn5c6e81Aim0JP5jueqCa0Jo
DNXF/8PDl6V6D/WB5cJLDkEoSIrMsbLgJJkxQtHDDdTFVPDPcvFhyTQb4s3kvPNh
LjAo2TcK9utJ0OncidGHKY/23zwoET4zY1zTtNm4diAqZtP6D/srqVeKcIqaKaDh
PuWy9YNjZ0xNFwSptEMjWigC9RG5VhYJV1n4FL+gMIy7LHb38KU7j3smNrawhVV+
GymGROP3nmemaLbkXEy6INlhZgKbU8RNL7qK00mqIYgT/apoJvqy9RdD0ERk2pSu
FeonflPgTC2mfathWNssVMwjtWfIFvcgv2mJRLhsccWg6u5hZnN5Otbtgruk2atc
FIltXhC3lj66Fo+iybRnu0bKE7iRWBfDDinFEIEKgXPdxdRJvj58UGbh2C9JhOlg
slMg66elghUGkEckjYwClwX9D+JqopSEzsAYD681OJBmMrizEr/eX2wh4qJBwRbN
qIVk42k6rGLp5orcoQPgbW0Axnu3ZAKp1jlHGcqGHn1DSv7O1gJGg82T1kqBMKky
5NwfAGX22h35y71ciVFrn48Rwd/+zubzs+qHmHpvJKwGy3cKjE6SKbHLPSShOROD
o17vJuYK+CmKJ9MIdjNfvaV8kMbznm9EYaM0+0VlJpY/MT8rTCjVgRk2ps1NjXy6
vBMQ3Nz+HL3IyxMp0FO32SOdF+Uwm3Y+16L7o909dSJIzDfyPR5gD/UySiOk1GIJ
gEs0u24SoeJKObaSs1jGkvPYA50vm4WLvmyxjA+sHHxfMZr5md5O+eT6nuG2DEu5
YUy28fTjHX6irq4DjMUTQQujRMT+4D9EUJnfRKWtwLXXwrfTaUa/GmoBNBAh1coR
hZhTiujj6k7AhAMZ25pAOVtj6RpkImp2eRunGNNroQEnxXw4Vogm+buhjkiYxcve
bzRRQhARXhbKdCdZ1+PUwYu6ZMkGoubE7dWk0ElD3dMGHGK5CUs31odeUst7+UOK
uLmFvX2cXl14505900CTRM4D9wnRnUu2QSV3i4O38k2xNZX+/5aO+/liCwrvCAHt
bzHLMcGx4PpFr6wgvJkGMc+N43V0EHwZyb+P40uXKRmlFR3O6Hm3H9R5Nd7vXq0o
sFTiwi+nz56Ws8z0pqWvqIxOJZubLa2fAa+TWgSEnjokRvBE9dfR5h4oYk8ilkgd
+lNCtFS+X4qbNXkx6WsA4MY7q/XaeEkLo5i2N6GUxIlcRzm14ocCfrYDFQ8Rszva
hsgre8t/bGu72xYLlZj0LbicOWuVZK/Gd1jvYijwR9yRSZ39Dr/z5Gc1sVAetVVw
wUqvlLu/1QkHhQKuHkkGdQqSOBudnVOaOYlutm4p+maq7sHpE0nZOrGLtsmVPvGz
TnQcarT2chl4KKpPtBkz5LV4l7s2php2PvWLJxOqICp9dOWb2Qz2sfw/yX9qKC7c
qD4RodQfWA4hOHtdDfJzqaSq0oQUMInS8dTW4GUu4OZAapRqrTmJHKPawwaDdm6R
f05Tn1tgSyPjXR5f2ex8pvAXD4FshuNNl7t9afcHLjtjsorR6iXmD02FPLW4/ce3
dHvZcxG50d/w4UmNqhVnYUAbTnr+6faBNnf2WyexHUnX3SJ+oioH8pqAU3vXKRjv
HIQrLDcABsSvV3e5eJ187fPo/s/R7TQoJwGmZi1ge0FjAAixU8Pi/9iFmujS53+X
s/JCaDo4VwRUuuoPd0+KE4KTbBDIOmK+qnoldYQ9s2LM+YFdio0rCVeKPo8+pFOY
0icWdg/JLjjsZkmuHPBdFMGgPFAsMLKWn2wjSj27DiDFDzYDdvvew26ae++2lobk
mByqDEHdADIBnin48Ff00hXR9KPwWBuH/ChsWktZnoopppiP5iNlVPS/IlxMKx72
xdwsnqOmyTtlu7wjIu4XM5KB6njP0dXij0/abo7fMlpxhhf+X89V+UnP5HQcEitH
5kFWH/8ozHI5j5+FZLwhGGa97Pu0V+gHciFxBbPWKHMx+CZjimjm/6a9JtmDXloG
MDoQfiQMttk/uctWewdzQy0PgbCM0ZOVBnI9uLxMjGB30SOJQOajYv3+Og99cgug
nrUVaHheWo5yNEjcJjX9IC3uYE1gjjL6EdgHJ9pMGLhTodTuWDESjjE5vmxvuOB8
TOCqNmXuscm4oC5QzEr7AVOgikOfUkSRW7FehN6pug/mjOCBc3ymKFdPAo1A0ck2
iUePNWptcP/wJKRYIahG0MAAYJt+pLR7xnNwn7fakEttVtTH4m7muyFb3tXl+cv0
IsRswl+D1ION7JL0ex8VZVXb/dZ47d3Cs33AM7YSeCsv5NcJCxmkXL4fEG9frrTq
8HEmLZRgHP4UlkUdSdp2AdjsXFfjG3VOwP9u3uoKwouf+cLbz4xDniI/6xYa9u+p
yqMUi8JZ7o0UP4d0Sa8l2RpzSvYX994KvAvapPDfhRiShq5u6rmj3SmIBmbwQ5Fl
sL8LHEfey4p4NfnBG61ZF/6nmqRqbrBenqJ/b7jiYqsuvv08Ec4MhTSf+X+FAwNv
LciLFKxRu2y6WZJcyWh7PVyyZdzvLMaVl0zADSQ8oMtZex43DW52n0VjtJtZWgmq
ZSxHc/ZNz6Se5XV7L7qCLapTZPy4PX7F0I4nB056DEjd2qJLJ6WcI9tvsTeOhkWF
8RtMdmUVTOWPJFmJG40hFa3FCNQe1GRy2urqlvgJlDKG96HvNBjeF9XRoFDvGTcw
7TVDUxGHQ/5YwDeGcC14h+J1nng0VPChxtPvuNZhDtGW2ZnU5ysX0qjVOSXeK+9p
F0PMWcF6yp+pGCCdmlHuN6Yi7HPYEaqltzN8xYPZv4Aan4I0xD+mUWuJZP+RxTQD
vX/PrNbQEBlgVZyDySG2Rx1XbuZbxLZxpzBmLT9fTIYnXiMykrwnpkP73pOa/vWj
+hGohBXN3cFlU4zFuEsuUQklmJEdbEbE7k/fRgl6D+KVwZSso93rhszb/rhczbsH
YWZA3DwnyfPf2YewPzusYwKgG8xYlCmXoejtK+0aBwTF67mxrGhos1mIlGH58jHG
spqgcQGG6yxzeq3EjFynhc8uZOW2zjO+ctYc+EeV93UuYd/XStb91lnbkPqXN9Li
zqIZ2RnLfwwANB72TDKlgkoLei0jiTsor/C+3E8fDYnCmQnzuVjkHCPpLDalrkNO
KPfYtq0eubyMT3M8n/oLO9Qitu5MhNr2kbPaknKqWZRiyyRwErY+YdoEO97t4nJM
byNeFw1zjEuQ90t/qoq70UbBZRmOAuF847VLV5r+/EqtD0ij9HxWoaqCvcM0XtdN
TlLyQ5npxg62hLmEtn1m5mNyTS7jWnEfBoEYUZXY2+uC1Qbup+M2a7r5jzOmRbEx
hXmze/Il4bUqfx07/TZS0VE1AEo0bTpsW1XrbbQsTmIN+0gEiGQoKgE8z6vBi+kW
T9qoW557RJnzyFJqy7on0OHAxQ6vJAupRpVjXJusVUQsz7vXjvl640O84QM7NHN5
5ZMrXipQpeyPk1ls2T9jpoyk/kgwJDT6QtpFEvC8roq6bNW3voJecGsB+3PdWwYm
RxV12MksOmQnRT+phEckB0+9NOO14AcOhKb51eDsjE0QrQ7/sEdEON94YwryAMJN
q4aD28sEUdLoPzd22glbADaVjBSYMXcL9yUJpL8uDEcxJrJP1TRT1gsL4PymfvxL
oW2SF74zcasQDVGUjBo9KdMl8SC+5DeL9yVAWOoQbgqQ/uWvhJyxZFegH5K7acas
le+M4qussFQ/ocfSYHpZFPpbB9SbG/QlWDHYD2VWYYPTQ98x72hZg7IdC6oZAaI/
tPm+1eRdETlVU3a1izCiGmQgOzIofHCwCaxN8aYfGeiw7v6PKUCHxQ4CkUhgm1+y
+c/EeFP3+0rBIWTbIp8eshsoJ0Sv1n3OBBUWkRVkxII4ZevXLmTxlK+bqJeKODjR
Ghdua8uv/0CbE/AnF7vmzDNI2zuw+uo5GQXeyAW5RAAAK6ZufADLShcV9Zw9mrbQ
s7/1u0LMZRQt9TcAG7Fd0hMMakOSNhTWhiv+KGZuuP7Ndz2uuIzWUT+Tpz80UOyc
dIZ4fXV7hDEeg5fLE6L+zf380r+wXABQ/vroOXSzqkOUzr5pMwoGJ5FXM/IwSRxM
wvAUQeuPmXqJYtwYMKeWyXVW4MZ7p3X/tfi/KhZhFPCU+w9FOTnPL4V/tLTHhzjj
lY9Zv7zCmKphK0NAGC/aKLcUze/GOyHJyETfhHCmSXpYJiYAUtWvzsqCbxe/NsPk
MXuV6/ce1EFDtIKkwrQJeaMJV5SyPFCyieTf5xM4dA7luwwauHtrbrpdS7Yn6gUX
WiOzARsrvpeCAAtl1/gcd9J4DsMbpsiE+h5TTd7mAbNIB38NLS6tzvAYeE8j4MNd
/LLWvGBxAncttxgGvK03voNTVcmEo5jEiGH3qVa9At6qh5qB2EcWs5KpkEDGTDcq
z8rJJCPwp1cx2NQbo8JM+NjD+NXPdh4t6erHgCk/0mOrzjG1yffJjj3vJbwHPDWN
d3pCM5EOs8B31bgH/5NMULJuovVpA4Qj/FtGC4tjLq8SfrBd/iKeUL04+rDB5Qd9
vSOacR2Q6DMbP4YvS/4pWEAtmxocWpduV3aoy7kxAZjf/T3kZDamd9yAt9B1QDVc
rluVhbbX0OrXrOxV347mxOoAYxriABNkiIzyIOI6KuLUHb7bket4q1Hjxsj9NCEO
MzTZhqf4K1gDxtpqiFB7Os9Cc8axF1Y6IKm/gq7Aaa6DQ0hY3k8ccnqKe8Vd52CL
gCmBaP/JPeFDTcsWcLnZ3U/0iqCtL68gjmDYuAVNmQoKtm1M1WxUe7U0HZTlvF4B
LXx1kXAM+P5JWSOVd5W3SZv5hBsdbZMq0WHbjOHkQHOwVy1RQ9lxTwSXLWbsnV3Q
0xcYPG+L7C3i+fvjAomWhsf2Zc6nPjXjQnQb+4EqYZ1CtU6qNnegupDEcfpX4Ha5
SOAWVPrFkT2YUZco9fsgoYacR9M6WBjb01N0tYsuQV71i5w3IjaxONgemd6l8S9y
pFTg21JbSt0Jn0rQU3vPuEl9IGNahmMfdAlGuBFNkzxakU5SPPKI+S/x2KmbYIfx
CiGdrIyQxneS9z1RNPA+J5+N51VM1vpWG6l6r4g0g2Aio20x/uy7QBTjBWFGq9Ej
9ZT99i2tVe84tdjRgHpLkIOj3hVpuBDhirab/NH4f1e/HKW8gWeEG1QlHdyiuybb
pE7kTAQ17J+gKKyeXaitho6siLEkg4Jk7eNFUeGsQkv0QfRBNxMHl/slLZeYZ7vL
HpkZ8/4ICKghXKV9OoT7PEZnWJd95ehmqH0F5nC6m2GQfDixp+bgb4IKap3xcFP+
IRYVGaW1hY3btjWUKhRaAg0+FgRmkJAhcJhHR1UBEpbSLbnJJ4VyWbsrqxv4CJoP
yUzm/qi710Dr+BmJQ9gelhzH3hkYhS+LExM1/fBU1AlJgQu0w/msnPpX8wwC1+op
OIAOCV4KyEvN/Yay/+NL3uvBPSC3EJZl6KUdULjj4JutIt6OKiCRnmcrgNUdxQsv
IwiDwRko8RM4/Q6ppiClGu8y2+Kj3hDPhwuMGq5VNKyL1nARB2/tMZyOX9/v0P54
Oob+PC7p1W6z7i7ZnzivpohgMEXkkUWoa7Gf+a2oaS/+bInprB/Nd6gRRIeda+wY
vwV1AAOrPThLOyvBuM4oa99Ll3V4zt/7KA3S7h3BDiPB8WGAZIDVh7nu56vqAKFj
I7eL4zmsCBKxSTjF6r2w5yoMbOhlJrzbFfyFBzwDldR4QMbvCn13ayDmmXOZZTvr
ad3H2YDJp36iMiFkclMego4+LUw5gGH8DHpCKwVjPSgmn1JqRv4+sqm5Wz2Cr7Rr
JHls9GRMY8rMVFkjOs2HBYA5SMcOgVwaJmqp+U1Swq0ozOTUULTSJI30ZYg9QIIx
YnBCcVoQUIYp0H9DnIXH5jOHlvD8Y4CYjRQYfifay0A6SWlVZpNFNkPecWMPrcl0
P3deB7grAUWbFjuG4qmtXRmB5erikFbuT1gLG7sYqay15oiIUw/NDR7wMdMuhI69
AgpXyQscfQP5HcXV8XZH2HB4Z349TMOxRCUmd+DdhjFT6ZK/YQoHzJQd+7yVGzD0
6zX5zVOmrPx+vDHlbOfWSJOlp6xnIn+/OZV7UcM9k8YTncswfhgbZWQOVD3SBgiJ
ebTgmQG3GLobl2aXGlttJ9KoBM+uLKLpYFriSqT/MV6h5OiYEI4xeef/3ddCvfpT
fhwrPlceBK9MpsyCBNSwFPN4N5fTqZMb0i0qca2H1uW6aCljOYaS2G5X+vqGrnwf
55uHI0XjM/7Y2XxZffLq6GkGDxUqgWLPAF8Q9+25WSZYPwXd3xvMutTFTeGOGsrH
5Is516b8BXBqV3vurvV3kzfTqQ+YFfE3ITSxNu2OSy7v1M+R/l8vPMBGe5BSAUn2
VNJYxj/7co2yp3j6O4mLYeWwWxclENik2t1jOH6wcnwkXluUAQ5vGRP96emueB0/
NOJDsqgIpXuqDY7ztnLAO/S0ISMMW6FKngM2wHcL11+hlwgYDGVgjyAtLeI8t4WR
1c/omVIoSUFnzSvpwa+h0NYlVUT6rbo/jAAzBSAJQXMdc9gOu7RP9cQNtRxDoPu9
8/ALtwh4KAPSXk9+F4t5pF4pQwaGiPnEZ85h5r30a3W27tLCBR9+Cgu8sLIfX1RI
Oqmx68JYWkSt6b/2mbcIC1hk8WC8DeTJOxQaR0cwUF03pEHAbv/V8TDFGaZDq5N4
ilUjfR9x+mRXsRHtdtSnAd0OSjXlOfrjGax+0ENVsLb6xJqB6hFCnGROLoMBtoZf
4k5qSPRTboT9O8mcVlsIc7vH95uhaYLl+G5PA1KdFqW1dqhMCqch/8PTDCRcEOpO
y+kzpQdiW2g+68zetdH5vSXAB+d32HcBOPUBn5KpcRBKF391BjHPn/vNbmgcESNZ
OFmICMyHWP6+oJhfvWF4SzkCb9FWFKhPQ01ME3JLZCPsa5PKnvkQ01QBtNbOtn91
lzT+eHfItVVvOtssvHESHYeaYBOObW8dFnt5iHA4j58SjvK2UniXz1R+20naYX/e
SO2Gkb4HNhWzVNuQxpTn3UzYhaeQrtoldaj3d2Cd3Ut0wptAyCBXZOg5qHSoRu3u
QHq8owdtSxTvQ/z5wXk2slLOEexhdqrwJmJXENVvGfKoUQc6TgMIDJdViTD01C/E
uONnD9JSRmPZQHFvz86kYZvyUwAISVDKbgGzY4omJ/XyAMu/k4T2NM9KVn//8r3q
kFjGY8K9rlchW7Pc44b7RM4tUA55T2lsdta0u75xMuqxAmJRYq5lLuMVqbyVR9m9
Me8bsZmq193msqxMzIbt/j2/uLovNncHlKCEqpE6bgKH7mOJCSzEm0clqnw9YQ2v
1kYJ172CxS60aUyvK6iFFd/w+bCbHPdFH8SdNSBJkvDBjr4Wvn8jE46pQHh0N81k
xYCZIIUKiO78x5m1MqmRq3YnYr88+sMPMfhAAWrb8ypA7kOI259FuJ+bYPCacS+Y
aEv8mg3flzF/w8GfsWzZ/H2eP3HZkVt7oMS2kAT5aM/CC8XDsUCYGiF63GzlS2Bd
oLlu8Tjai+xAEQ2ec/kSJHHgBu+n88Vb6t+2xbt1BGZK7aOv/O6X0cr5+Y/hbxr0
/eDP8CkWbvspat5sxxsRS8tBUGupncSfeSsEF/JOpOsJZ0HS1NXx8ToEL+PZyOTD
egOAPKPGBpLcTZyRiQ4MU/ZBMU/uH+8J2swyWAqoKOCaX2U5PbwcysJscWldWgPj
Z5PhZv9wM2n81dG7p5wpM0JSb8ZMJBIXpss6fiRSCuM01khn0Z17kqBC7IZdE+qK
uhHB07R18C8qqcaGTSUAtp6sG1jYnKtNLqZTuVXFRmwtq1bGSvv65Y1WO5MxOzLc
2wdHDSWKHYZpxcpakDmJ6yx1HO4RhiFTnrfSmXSAxW/oolc7I6yTPsiqi8rbFij+
nnqOvsoRzNQZiyf2KoK4c9ZZh3JSHp4Sq4/fP/aroq3+xK029tHENbozktW25adK
2yJJHFyxmA9yqGEH7Wyfz7jRZdv7bert2uF0+6GbfJJx/6F5p8yRcUCRneOVstDW
u6yGURaSM5/YRvK6992txN/JvPcnkPUEz1PK9j2ZGYbagMg54PYpxIf0xo2tBId+
RI0Pwu3wYCp4P5sN+zlNHsHcg8p0g7VNxET/Kownm7y/oz2NC2t6Z3SPJYa6CTkD
FSjNLEWM5N8aExlCSbVSkGQuIJfGwMg+YleVwoXpWHjfFaxmjoOKf1D7uka8owPo
wIMHwYWsSbEoKYm6zATAnqoJsWlzJVavzWv9ynrRVS+eaIuZBPHUkubiFPon1m/r
S/lQiZAvWaUYJdiIeEkT2OTvIgOmoovWaeiJ8bYiaYUUO2xEkd75N2rmzEa0rC4Z
3oDzDt2wpoxkmqi1TdPFnlA3lSn3rry+xRl0Ie9diElNM3Jp60SxtZFsBnXGrV1/
p4LEX/XjsXWhVy1dpFBwiaCBGgjr9LAs3BOT6jA3HQu+gPK6NcMYOK5iobVyc42B
KeI9378VCFvfwdIRzWIS+16c4KRENvvxItnBo7yrmOB78VwtC5YqMTJYtBvoIh7u
E58XR7zWIJNQnSG/8M/H4uuHSmV/V7kE/Ct1LD+/Mw6dWk/OKLZ0vICxNinOI8hx
Br5iXAitwcj47M/AFd6fHI2LCTlKSpDhkPJO8nx/ZKKkLf7G2GVthfr1qhtiy+VU
mMtdk0IAYaqSmjCXa0KW5Rl1Tx0CiSfcAorY+iClYWdq7bOLRfqLBWverlxagh4a
KcZmID7mSR2HphHjD/MlKN6Zvf+fBCjNkCrE1ZXUw2AzJZk7VVSueLNKE5Yz2QDu
HrjK6Nwef/M7GG5oxCkg/r/ABlcUkR1oW78gQAMCdr4+f8s9S1lccgFXpH0vaiMv
PRlXdmjU2THIwaEXwfsnFOwnItTTwWzisMgXR0gjIsyMdKxke/EJkcQngVjrHrj2
xaMmt6v36iBtRMdwRaxvNAxNlxQevv8LtPQBwAVAEWng3Vxo92iKMUtS9hv47VT2
+wPwpNeIaaRnnQuBE0gT1chE6y3AoApS/VhuSTgIH0scp1R9LC+KoTLp40vZTGNo
UYXQX8hk1IS7w6uolcIyOaGsSyFtSLTSmWKBM+u38K1wav/aUzDBW75F5oMxoJAu
ml4SZ8ZVRO549PcqZ+f2857ALLkLkLZOAlyczLpsWSyYxjXx1BdIRJfOlOYUUrWH
FPbQtdhqW1l3MTtU3XF1S12VdVn4zc5JNb+YqgC+KZ1hIuQy7e52QHWIJmFP2KCu
SNPFXDkihy+DPyZPYG3WAmEPG/u4LKqNMBXxmMlbTSntZnCFEioKITvE1kCfZPqZ
b5nJWcUIRAnVi5SYnz4dUzbNoGRX5S+ooMQ9MBwxpUTOw86PYzKsJrTTaNx0Wzyk
Ewo5JvGB0YhPxl1WDZVsiEeT/ZFjlsrNLplOqce++j2SDVubhI2OwVo4Gw/x8PAf
gwuIQ+yaLesSWgeunhTS2mgooYZ6r0l93zI2QFvBYweYik8s7ZoW+B5Kdc+cF8VW
HR2nTAHK6c4llLFgQ04e5bOGeg9Z5FWZhR/emPZ8KVDac0+6agauJvvA7wsKSwDZ
hcmBW3VtZVQUq7lsrbMdsNU2r2/lAy52Tu95NEvEafx1KJvTdYKX5w2wzHdP+Jz1
wQSP39UW2AThVQy0+E9x2u1VierCWmjnXm99hNthA3nRNTmOqEdBaSvkTX0R7TMz
LXroby3eoAkLFMeCcRp6Gjxo/3UCmJbV91iaW49Cjnku54LFoTryxtgoZ6UrHK8z
0ToEV1vii0vv1BZBOvuKoajP6/E/ffKtX4uyIfq5mn+7ccV3CPFF47pL6mvZ4/cy
oQdPsIBu5eAA7hQL7mUB/Uy65Un851MeceT9M34lw//c1IVDdWZpAdXDUYO23dI9
wnDAeBPSuPi0/dhEE0jg8jeNpzdqQvxDoUBGxKdukKOoomuK5Jck2g4rZGW/mt02
NjBni2r77f4GSYntMGXJ5+W9vLKSa7MD3R8LzrQcOBnTCtspW92df0RMYxgGnoAo
HwSWtaRTV/xzQyvY44gsiNKF7yKEdbD55dpov3OlgipV9tnZQ1u/FUiFetQq0wYj
XPScXDC9Om+euXutGwWu6HXcF1p4Q2uWnPZ2qnHAM0FI2YuluiOP916e2qmQm4VS
jsefFyHLofTl8rLlBGs1UMpHp2G8ZdKVdOLUEDCEZBmo0wlKLPfId0uJ02FCYk2I
0MDx3NQPoFpSP3lqzXii4VkGzQBg6tpI/x36va0425ScfCTll5haI62B2mh3t0cW
MZ9/ConxjmUOXmrvzMBFzEQrOM2wJrLTWyb5Bo1mIDGm4Yc6NQkkA5Jt94JF3Gxw
81UxMCAotJA4N11Ye8YTygKUmhvCi5qtr9C5lQAv1Fmnw4zIPcFOHgBpvgFIPt9v
rn55vwQ0AyHNFsQECTDZZDxbiCaQeymcjP3xQsWZajsA8lnK3LrXYSFr4urYLLkB
3sP+YDvffKpXMcFkq6gitaM7oh9r4eoNJV4GcS0BIl88wku28x9SwSOBEuyTdVGA
Ky1vAnmHd3pn08Sq0WwjoZzJOHqB3LGFRI7y6MfjliSZvKkbb2BwyoTZnT6XiFxw
pq86c8u2SFh/I1Uv2GTBS8P6DJZteZ73KHEIfA97/BUTtKbdEbcLfFUdqho8t2vU
D9buiYduHAdeCqQimpHCegYXTbXp19AsAyXdlai3MkZnTM7QKbyiF34c1VnnH+bw
5Bt0xbTTPBMbSf5BvQiEiuHd5T8SBtG4lub0+C5YXzOnWeYhq2lj4GIIS48ojTFB
hFR+KjoRy0zS0ASYP9eeUYK6YTFAwVQnqZAkIPzgb2SpUeD0Tv5acoxz+1CS1E+R
Wr1dLkK6FjVF0O8dssC+4oKbRP2s99xLKHlYiCbIgS85k3uDy+PImuqVHUcauI5j
vaphlfdetF9WwlcAUW1XvaNMeiwJFkes+2E8GAQFyhavjJs75DGvHPC7qdHoT3Jg
pLKgenRR3WDhytSyAgbWw+rdx+pfXWKLYUE0TDIl8POHmY8A2vlH31nCm5sEnjC6
12a3Bu1m3sF269XBK3Kt7D1pxulnUjgY8psH444wM+pVJZiJepKR6Bkk4ET4+RZ3
xWgM9k4J5xoWrJSDBY8KQJ1oF406n4JTvXN7sddj7P7Y4V1Tirxcze3IdHfM9ja9
WXXoI9YsSc3HOjj9g/gF8Y0a4PZ3OZGUc48DQ9S82MqNdvtT1HXf2/dxKXHlcMjs
0zIHj1k+f5hmG0uHZNpOe9o15ru1x7L+rBFyODw0O4f+rwPo7tl9/1tkXzV6+CyF
umgk7cbwg7kQPOciAp23QF+vkWWsa7K2D+R++63fnQGiHmafin+PV4Y+avfQma2q
+X5J3HsMizfMWjzJSALgU2bANfTIpo09OOlraq+gynaMZnJzxLGqqQmREUYAv/42
l3Xf1IWx3sd1i+LLJpRYzJ+pSTZbAWgvzdPTC/SHov7ZJo2gMoawJAvs2IQNqFLM
6Kw43XjKa1GxiUy83emckA2+bmjtzBFas1Mo8nkdY0pvlaUm1itUKuYZYtsKayqS
J7+Hl/8QUIjbNAdK1Oq8ZVt5GMuE1cg6kK6gy9LeweQx5IXoVQ4NcHLpxw1pwjk/
IDo6jf/+8g8NWD4ie//u0Gdh7C54XhGNxIAvu9EMnINSs+7Z4v1JzfJd2PsDlIFG
nIEIAfiYKaHQ8leOd+6V6EBD+HcAyWcZ+aeQe7E/Qsy9+Z0U5GPFKSB4ZsvPW3um
YLj3OGFSGQdl3WeSiFpxYP/Sx0Vt2Z552u/cQlxEDigCb6tqayBeNW7vVnwsOrjL
l7k93NeYRnZ73JQ2ljW+mM1Aq17znyOysYT7zRWwHu1cdOhSmQYc+Kln6Y8WE79D
vDcyKHg4vARQx89yennuk9LE6Ii71y1iM9nKWVceJeSIsfGdNfshxRcVNHKInGPG
K1nNwY3LKw86PTTq9WV9Y+9KjTC0z9wnXxuNoSsOOn1eh7Tq+8kHe3/h1HUXxdup
d6gFIQiNMyU4qRhVTC71K92X0bnR9awHIzY/+yQXWHvhMfCslxBDvAtkkCajxbV5
OlYXkd9YRB/dU1HLP/Pw4N9Qn/vaQMEytwIYIvGTVC0=
`protect END_PROTECTED
