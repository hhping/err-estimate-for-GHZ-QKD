`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFj/uNbzNqt2RFa6HPsWRD0TZ+A/gOMSCSLbh1u2WC4iNZbxufrKAsuDXQUiEh/t
Q7npW+7xsssc9nLj23pL9hudmFHysaCiMNdgqr6NAoAQaudVEFRF4nPe8b7IoEiS
NnLI0mNN3eTCpHxtq7dcyzVRkQa5Zyi4CtnsQ6p5k/hr9SHDXLxZjz2Y2CzRWK6f
CvxO3ithxS4X41frxtLNC8xELDXy9XewDOpm9QITmeGruzuuEtP/J+srU6EQMFVO
AeQQFT6IILpoyi/ZbAb2VcKrn717bz5wKji/11/sikP8RfW1sNspcdwmZ7rNZ76G
jQ29kyToeQmJlOa3xUsKoP7rKclypG3evYGLIZ4at46il/lMvJ8qsDOun3nDzNCR
mVgPJMp2s1IDIjAy9QVAx3ChrCzXdYQxL0VkYa4kGc5+eKjwAAthp7VEGc0IecvW
uLx7fs5rOoh3kgtrMnwzQw==
`protect END_PROTECTED
