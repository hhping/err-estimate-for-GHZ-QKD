`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QI31HfNcj63VuLmlFPC9ClwgXoXW7WWO3qjKAv0++PXm/y8wmKDiLeAd8v7On/yE
G2icdLy5UGlDqE5GSnX+MFaQWONpjBL9kJpFIRvFYm2K2dpUUkQCuYxzlo6lqGVE
PgBaqL1yU/nLMPHvxTsOkRIDBluMPnRmHXdGu/y5IZnnCarOosyFPq5ZDG6JfkdA
RCaffQYJjACKOvYESBtR2K7mACV6Dp8bEvSMeS9YuOLhATJm/zw7GLzC05/ye8Kn
Ml2NmNEgYtEMJ7mnjtAFzSqUYAaEcOWQazz3Fqb5lwyk9v4HvxZjYI7UCH5wnaaB
GA2mE8dIRkXJyFYCBtJlDvBUAN+YoFBzE5x3K2hsH/MCiyL142lBYxkzlZxMxat7
D6+f9EjueYeFVaGMX9CK5mSwcwM9iN/PxDzuNXG65cVofSYDwz4mEZdcjKlFCsmQ
XZtgaRMWMQUcn/5TIPRLreLDmzgjq3zqUa4NnE47YxSHgbft2qHE9SKxaHMidVNV
`protect END_PROTECTED
