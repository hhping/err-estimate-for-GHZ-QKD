`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4XTSUSUKo77+ENbWYw+OmD25h4RoFbSODstoyGbWv5SKQKFrhFe8b7vNXDKFh8y
ZM4n2DPpeTMfTib6jZHBtSF1QRKPJS/7iipzipPbuJNIQzcWXVOsygb/wJcbCWgR
bUKQiQ1fqHK7IKPJlQAmzE+iab67QbQKdU5fo9OqZF+8/Gd44FBQvIJGQydal+WX
pGeSlWcQm/QUDJYKkq6b9NFhevRk/rhrU/0vUB3yTv+ceuMt0qnI0gdPjzuaFlly
k+KrU5as7II2+zNqo4QhCwg5Vy0X8ZukPZgubP8vVbthEODxLrIM5LnmdXv7+XTk
C4R38BLm37Ej5WmEzSeHjnrga4GAvTmykPhHMcJ7ZnE7BKkop2ucx7BE2ViTQ1rl
2tQCIpnYOz46cGZqXECHD/Dm66bHLZ0eS1HyTuccrPDfBYpstFea8KR/E3b50Gl/
LBY0TZDFNo6qYsJbxXTkFHgKWSnPkcqOnzHljuJfHTqoPKNBe/6M7Yd5e2kYOzjN
hncZFSXnQTU/vtB/Hs9N/69QjA/I+zhLTL5tDfpAxncwbRM+0UddSNGHVCFMQruN
sUh4/oqMHod+7aJq5TKWsHjucjfyA7DvH4LVqLmz4HtgjYZAwQ4E43b+iNxOc63C
9R64KX9Sk8MdpcmnB54yaxCl3bwahOOM86v+w8auoCDidQE4S0/i/uisSHjB17Om
9H72s1VnjZbermXox++DwgBT864m5WJjn4O/fzooZ+MkBuwJkm+RT+qf58A+sRaX
pjXb3frOY/vxF4DlaLRDcFGd7Zkotuz1BgUV0JMITTjYDma2QubvftxAmqH3aJAB
ZLE5PdipCP07B6lXsN/fZY7Lb8LsRctTXANW8Ymtoak0cfdzZDWU/ocZUGWNw/TZ
8CDwwDqoYe31CKTXt9neH17fj4KP2fIXNCpJp4MQc2bq1mGSezDGx/NH3/orzm7z
HMDUMOv9oyfcAke5KZN7GsiHapvYapD6Dl2m5a8jYyyjTiRNZ6Py7+pHnR7mPK0U
Ufr8V9D0LYzKEuXBjQWMKPDOWfaUuHlQ8BYJCN1jCXUnY8F2RPZf07f+2g/Mn2lo
7IGixQK9j6YRgFwqUmE5ByUgI1928aojqThfCPe7GWnCOWYu3dSS8U7x/psEMjSU
Z2ZnsnLHW14FetJj65cDoMLh6io9hiD63lkFbdnoVtrflIIRWVZOIQIcL8+d3dvz
zJMEPdzcAgWf0zMvYGPQ7FSKqpc/4LNnyzz22svfSQh894Lkgvj4dzy9nDKekBjD
0qiezUkLTm/ireiyKBoJKsetlBKlsAH/7Z9P1SQXBH8=
`protect END_PROTECTED
