`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGVImb85XONTbiEpuiteQq4uN1eIOAGYZo3IyxRh4mJ/JBoDJxIhykbwHPfvqRqK
bnTD3OpE+G3d5q46O+Lch24NIKIr8OJfQ26vjogRiWHReF8WRs1XfBu2qiqu/fcc
D6phIl8MDdJ3sdE1XVK2CLoVBViCAuebIODTvTdIbjGb3nUy1B9PIgUrs9gktUEF
K/6rclaxcmj/adgtXKDlQ1z52aENIMCq4lUOXE078j4KvENtU9TqtSwDvChkaTRH
gEr09uOtVkVSf7mYkEslod94yTW9Dq3BhOoCOpmLvPdC9wHxscfU/A08hgNBhLU6
dngm7B3xXcp/ozilpVNSfoMQA+sVfjSEyFDSD+VKNMK8oXqyhEv+wRI259gBs0zl
XSl4ya5o5k6eqq6GGUhMZNXKvxqITC6SvLg/8+77iatLU/mawh9iVx0KKR7CHczE
O9IygKpaUFAzCKyYJ6h3bxF4tMOZ42Su1w7xI3FGseoK6eY0K+AT3RUL67NFyDd8
ViEDFTgrgngW+Fg0iIocVVcRo1upEjKCUAMo6ZdFRxjCcaY7U++zQtvu7RIWsosp
n0zj93m74+xw+97d14h8WF63JClyVGnf0Xqg0bA5Ixg=
`protect END_PROTECTED
