`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YqNQTKHmYRe75Z0PAWp7kSM0jXrmEMlJLENtyCKpCmj/RbLT64z9McbdDKkJXajt
3R/Bp36WelOcfPPmegn3QJR8rHpYj9yVhy9aainMs/j6LtnfRku/bzYULnhBGmcB
ztEXZAD6t59tvsl0ERWccZKHh+X17Cp/tn7eUqs9d9BEhoy0KmZvwV0jiYDH4Ple
J/twSa2OMLL1kYtMxDYRdqxX87fr9MUvCqWvOXGuyX/v1006sVRMCiICG66dqIhX
wxuVJfbw/5+3onN6uqP78oqDIUu6dEcibU6y0UTO0UDO0NbY90FywFkrviBoy6TH
pHKotNOmSxgHHXZBOe1Av+g4y4pfSI3g1ll3BFpiL87HZse8+hoOFJ9H7WftOxLp
TKB4BfLbzDAVl9kWqlLQ+pfwYz9LUFnH4vM6XIrNQFoBsej11/zi1OcwH3ikmJvA
uYfnvwyf55P2fVdO2Itexbhe9m2XeuorAyZxzjDvwM5R3+XxcNYzvWDmfdhbt9Vs
mTAQtEl2b0ncPNh6ZwdtmcmkIn42hDGc8HCALdYc30PnYMsy2BNfmKQu2l5DIahP
z3Tfx1xMzv303TaBDPSJWbavBERTPjftmUZxyXb3aMpaiJ9616mkgPoSjlTjxjBI
4qfRAOY7vhh+fCUl70ZcRz3gf4orz7Gml1F/f1Ht+jnWMg5LpzolRdnLI6RXE1KM
awK707Wtz4CakXZj3qVWbpTgnk3HnAjE7mWLUWfP07sSkW9aYYm9hjjc9iDd4LdY
boKnOuyuzo2gSHcnmsHQ8qScs7oXeq6JwTgzIMGSweco7pfl8++7GiN4rWT5nJUD
U/X05/GhHXM4cYo2w0AaR5IvvNwKNgmcONoK0gJMW1HnalzJOoXLumyx1g6bTbIK
pOHxVJfyCBU/PC82YRLZZQ==
`protect END_PROTECTED
