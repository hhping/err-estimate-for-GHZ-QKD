`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCzJTN93DYVnU38sfkFeTRFV+MWmrA460aKM0Z/MG3Eqs+dxYV4aLfU17Gi7uVrb
6q6SkvcUqHNcMDoRzPn3EilAaAwoecuzdgkFKkF75QSdnmKHGvRwTaeENRW6Qvx4
OFNvrJXGAYwdd+DDTstJyBHFkm5h7ghTUMGeYUkZdco4rbZlKfs0Uv13JzuGx3GP
4Alf8xOXDLOiG+OeGUrA6BpHl7prBMtBYn5Glb9S6wP2umGIA9tCY6lw2nqkX/8o
LU6A67mlXDy/X0V6kvUjrw7OYUSrwaF/hN2I6wS6m5FZryxbiZr8RzVEE1PlX7Bu
nMgf8H+swVHX6hRYo0t31A==
`protect END_PROTECTED
