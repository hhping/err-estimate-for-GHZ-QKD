`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hQgnr0uqO709XcHUVzhVbvjl+kTnfNSQbhrOI6gWXNt+qKjSKGc1OPLsygeyG2ft
60/8sEg8ABI48n1PgddasxpBUStvIXvMx4zJTOCfw7fCfcTy7vNHSBiCo3RLv2lS
ILkhxJ3DAN/DuVaowHnfjNfY2t1R0wQHxoHnLJf3Z0gEiSe/N4JICyOmLGqRs5iz
30YyId02WDTBAmFlUggua1bh8se1MnclUJA75cL4bfyQ3XqC3Izg1c2+KD9W5/ft
p81LEoANTpEz4jnv6xggRsPST+e5+Iv/UbVVTd3VO8UlhtG+PUMROyz4jgpP/1gg
x5dODV3sOjb7Rzq8I8xUecK+GyrE1TIlN7SlO5K2drfMySH4cr8iHcc0Kh1IhsPb
xT3LYMaj/fYdImQlmH5xnrryXx9najhJ+T1Msfm4U7nKV1eHjHbgBQOj+2KE5O23
Caq5B5vyrI//7YY33TfS5PYnTS6apBzdtenhHbmf+Dmg4F+aEatpgPdFkE1tUqFw
aJJeT9Pszo7I3I8k5+OQcF1dc/dQ7dL/ZJ4/yn326vMj45jqJF3JNCWWpVgwobyr
L9ngte26vKb6g/8rmP1Gz1uKibWVvVy5n/Gu/9a572XCgHeWV/pWjpSwMhChh5Sg
m/0b8tIX+WdAsMfLoj0t0wc0RbFQn060zTTnwluPTmv7UI7w/LzrcalyywXLb4v8
GDHYdTK36TkkYGsrqCTo9Tqte/6sdditdd4+ZDb2BK3ujbkrtb6ggnlC7ZPfkHJI
1J+E+OSxsWVW/jBz/HAdC+XUBWwADOwrTZHGV9NGkyDqXMQMvyRnsKcIOMeYuJ2d
WWcsnGHOANNvAs/shJ9Ralek8oDUjovu8VBeLKJvNLPuIWTJFRhSNIfJuhMd8dOW
WnVg52SiqqVGZvWsXOTVctUc711s2doO9t9TLaesi5o5xkwOPoNZfYSZwnZ12WjJ
5OthuR7n+a8e4rXqW0IhUy7G3MPbMN9fhoNNLhnKlt3AL+fncBr4pR9hXTIirgBA
FWhVVUDpsRc0RmqGE/z8EZWOjyue3EsB8Ulrkhzac5V61Y5ta+o4SGzi6kRrJ6aC
WSRFudxruWxO1BgrAFlCXembNrSe65K7gSoasu5N2fzwh3YNC7g+tzYMJiDB/tGt
cK8celyMV2lLLSKzW2EQuQOKiz8D6Pc1YQDnHnoEZiLwn+3MeSAJnwLc2H1LsjcH
/++J/F9gceRCxllFtxQuVwwKkr6Tf/um5WeDdTiU4LHHKfhykwB9EngJjLukE1zy
FRU3BMJEE3LJQaeh5Wu3sWtiUXfnr/XtKm+JjzCZpemqdrBn8o5BtOobnvP6bLz+
Om+nGxc0yPym6LS+ilcdNi1xvE6+ASAwZR98mCsymCLKYqIhAnZWlb9XD8//e4zz
QO5iSmrYByK1VK4j5zePiUaQQIi4xRgOS87vnp75pRb1HPQT+wDFsbEaHXW2ldCY
ra2oKDiWe4B8xxnkbzTOxiZpguizLmYtyJIvtsndTJ9eRuYAQG3rRC5w8ZaeEepX
P4fcFFOZUJSjRHb5cWfHMDaGmGNmv8ymKAZbqdFW97zt7X+/oKMN3tivcxT8cQwZ
QcVqpQ7R30HwYNlcL30q/+GwbKq2NQulbsSHfv8LhV/1zYniBS0sm6VVk5/+e7a+
SdLZoQvDsHc8252SSy4TDOMiFK5FbZt+MFjsLDYLLqY=
`protect END_PROTECTED
