`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/pH087J05iM+jP7Wuqc1u36U7n5c1J/vAoXBzbGyz5+Htv6hCGu6yiM0too9qW3x
vsaF8yfwt9wTKOEZSBsTGEvt9QyDXL4IIiP79qqA+mjU2mSMd5QfD6R/VAjMfVsv
Lq37k3CROQDg5dU8BpRHq+p++S7TVDfpVThG2QvLwD8SlTJpAkW2msHAlub7w26+
1Kdfx5joYNDMeM6VU68t7oivbTg9bTjzvaxwYIL1MDVGVQ8xxVoHG5C/upCCylSu
J41C717mLWMb1+i+UocBAxYXzWudAcgbFmUG7avbwcE=
`protect END_PROTECTED
