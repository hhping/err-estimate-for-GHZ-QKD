`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iUa/RsxSylJHHPC7VuVnktbWun5PsT4J/ExPydLkDikz+ewk5jTngTcqU+mfeSa
7P2b8PnWj1XXPf+sNmj2Wlxm0Dc0et8Fa5mDfMRAxZfQcA0jwTBw7hZ01SVJVpsb
JaY5Yoau/TesEZ3TG3PmCSZwcOtGkTszxMcVRqvlDLvnCuN3Ja6wMuzO+mDKzDqU
K04eSHY5Lbw1dz2RYkqNRAIhEjY8rOHKiaQkY5VY2gWWY4L6dGCs0MpKXxz8j82u
dp5rSdEFJrE1MK+2s1/cOdRRZypcgnck/9z4pDjrVcmgWPWdiFjNHpGE0RvVj67g
dRcid5PgFvCz6/5RxIwXT9L1042dR+LTRo3Tui9tt5VNgnQUdk8dORzjNqqtLiek
kZjjJejaUhSh0cOJX2ONbmgSS5KDszHcldcfb5v9QAlMNJepnYkb2ZDEQaOfa20c
1S/xE4TY0K70eodyANEQcR2FSiKn3AG4Fz/lF9ErEhZILZIFSoxJDmO4CaYEGyki
`protect END_PROTECTED
