`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMivAmbOTpvu1Y2RK1AUMQAjIcjoUGusz2ovLdi1MGApmyrvTyGKO2dbjgnA5CM3
ccOjNWpe3c/MT+V1tmYakH1+xA53qo/mOJcnGkpUeKPp517wgstbX6o0CdxB5V1M
6SG2HMbeE4+wYzV4Kv7iCxV4RXOQ5Lr9zrp6/JW5AhuW9zHTRX/B6S4QsJIb8fQR
ikDPNLKm2WBzlxe7QbhLeJD8+kaDrHuHUeKqlPHoYPDAycYnzZnuXZuIAjYJS69J
XxwxQpt/W3jDQsSYGe4078Q2BMG6Qy3X7RFNMId/IcihYdy+7s/zX7zTAX6pkSOw
Przr7NicSTUL+Qp8cTUcGScNv8aygIHn8VRc7m19a8nF5R6Uzp4inc7fYM6FUJB9
2KJr9V1GhSFvwtbi0sAfmferWpdFepvQdNHbozVTcYon5aAFjURib3OHbQzKPJB7
oGZsHdGlqpP7K7VA6HN1IozHxw4Z74w5SJgYRmpl8JIwUdbhf4S1+o8L04raTW7z
/JG7B+Nj3foYLGon+N2Uypq6MW3wugc8sXttyqX3aOHPUY30C2xL9A3tzQvyxidw
4Xmt0jGtk7bhpLVSAq7xDJhmve8jclaVB8FXOMUmrjt3UEDvDdYEeu+IsFdsvI5o
`protect END_PROTECTED
