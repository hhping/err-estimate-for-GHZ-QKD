library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_rx_pld_pcs_interface is
    generic(
        enable_debug_info: string  := "true";
        hd_10g_advanced_user_mode_rx: string  := "disable";
        hd_10g_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_10g_ctrl_plane_bonding_rx: string  := "individual_rx";
        hd_10g_fifo_mode_rx: string  := "fifo_rx";
        hd_10g_low_latency_en_rx: string  := "enable";
        hd_10g_lpbk_en  : string  := "disable";
        hd_10g_pma_dw_rx: string  := "pma_64b_rx";
        hd_10g_prot_mode_rx: string  := "disabled_prot_mode_rx";
        hd_10g_shared_fifo_width_rx: string  := "single_rx";
        hd_10g_sup_mode : string  := "user_mode";
        hd_10g_test_bus_mode: string  := "tx";
        hd_8g_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_8g_ctrl_plane_bonding_rx: string  := "individual_rx";
        hd_8g_fifo_mode_rx: string  := "fifo_rx";
        hd_8g_hip_mode  : string  := "disable";
        hd_8g_lpbk_en   : string  := "disable";
        hd_8g_pma_dw_rx : string  := "pma_8b_rx";
        hd_8g_prot_mode_rx: string  := "disabled_prot_mode_rx";
        hd_8g_sup_mode  : string  := "user_mode";
        hd_chnl_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_chnl_clklow_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_ctrl_plane_bonding_rx: string  := "individual_rx";
        hd_chnl_fref_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_frequency_rules_en: string  := "disable";
        hd_chnl_func_mode: string  := "disable";
        hd_chnl_hclk_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_hip_en  : string  := "disable";
        hd_chnl_hrdrstctl_en: string  := "disable";
        hd_chnl_low_latency_en_rx: string  := "disable";
        hd_chnl_lpbk_en : string  := "disable";
        hd_chnl_operating_voltage: string  := "standard";
        hd_chnl_pcs_ac_pwr_rules_en: string  := "disable";
        hd_chnl_pcs_pair_ac_pwr_uw_per_mhz: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pcs_rx_ac_pwr_uw_per_mhz: vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pcs_rx_pwr_scaling_clk: string  := "pma_rx_clk";
        hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pld_fifo_mode_rx: string  := "fifo_rx";
        hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pld_rx_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_pma_dw_rx: string  := "pma_8b_rx";
        hd_chnl_pma_rx_clk_hz: vl_logic_vector(0 to 29) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        hd_chnl_prot_mode_rx: string  := "disabled_prot_mode_rx";
        hd_chnl_shared_fifo_width_rx: string  := "single_rx";
        hd_chnl_speed_grade: string  := "e2";
        hd_chnl_sup_mode: string  := "user_mode";
        hd_chnl_transparent_pcs_rx: string  := "disable";
        hd_fifo_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_fifo_prot_mode_rx: string  := "teng_mode_rx";
        hd_fifo_shared_fifo_width_rx: string  := "single_rx";
        hd_fifo_sup_mode: string  := "user_mode";
        hd_g3_prot_mode : string  := "disabled_prot_mode";
        hd_g3_sup_mode  : string  := "user_mode";
        hd_krfec_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_krfec_low_latency_en_rx: string  := "disable";
        hd_krfec_lpbk_en: string  := "disable";
        hd_krfec_prot_mode_rx: string  := "disabled_prot_mode_rx";
        hd_krfec_sup_mode: string  := "user_mode";
        hd_krfec_test_bus_mode: string  := "tx";
        hd_pldif_hrdrstctl_en: string  := "disable";
        hd_pldif_prot_mode_rx: string  := "disabled_prot_mode_rx";
        hd_pldif_sup_mode: string  := "user_mode";
        hd_pmaif_channel_operation_mode: string  := "tx_rx_pair_enabled";
        hd_pmaif_lpbk_en: string  := "disable";
        hd_pmaif_pma_dw_rx: string  := "pma_8b_rx";
        hd_pmaif_prot_mode_rx: string  := "disabled_prot_mode_rx";
        hd_pmaif_sim_mode: string  := "disable";
        hd_pmaif_sup_mode: string  := "user_mode";
        pcs_rx_block_sel: string  := "pcs_direct";
        pcs_rx_clk_out_sel: string  := "teng_clk_out";
        pcs_rx_clk_sel  : string  := "pld_rx_clk";
        pcs_rx_hip_clk_en: string  := "hip_rx_enable";
        pcs_rx_output_sel: string  := "teng_output";
        reconfig_settings: string  := "{}";
        silicon_rev     : string  := "20nm5es"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        int_pldif_10g_rx_align_val: in     vl_logic;
        int_pldif_10g_rx_blk_lock: in     vl_logic;
        int_pldif_10g_rx_clk_out: in     vl_logic;
        int_pldif_10g_rx_clk_out_pld_if: in     vl_logic;
        int_pldif_10g_rx_control: in     vl_logic_vector(19 downto 0);
        int_pldif_10g_rx_crc32_err: in     vl_logic;
        int_pldif_10g_rx_data: in     vl_logic_vector(127 downto 0);
        int_pldif_10g_rx_data_valid: in     vl_logic;
        int_pldif_10g_rx_diag_status: in     vl_logic_vector(1 downto 0);
        int_pldif_10g_rx_empty: in     vl_logic;
        int_pldif_10g_rx_fifo_del: in     vl_logic;
        int_pldif_10g_rx_fifo_insert: in     vl_logic;
        int_pldif_10g_rx_fifo_num: in     vl_logic_vector(4 downto 0);
        int_pldif_10g_rx_frame_lock: in     vl_logic;
        int_pldif_10g_rx_hi_ber: in     vl_logic;
        int_pldif_10g_rx_oflw_err: in     vl_logic;
        int_pldif_10g_rx_pempty: in     vl_logic;
        int_pldif_10g_rx_pfull: in     vl_logic;
        int_pldif_10g_rx_rx_frame: in     vl_logic;
        int_pldif_8g_a1a2_k1k2_flag: in     vl_logic_vector(3 downto 0);
        int_pldif_8g_empty_rmf: in     vl_logic;
        int_pldif_8g_empty_rx: in     vl_logic;
        int_pldif_8g_full_rmf: in     vl_logic;
        int_pldif_8g_full_rx: in     vl_logic;
        int_pldif_8g_phystatus: in     vl_logic;
        int_pldif_8g_rx_blk_start: in     vl_logic_vector(3 downto 0);
        int_pldif_8g_rx_clk: in     vl_logic;
        int_pldif_8g_rx_clk_out_pld_if: in     vl_logic;
        int_pldif_8g_rx_data_valid: in     vl_logic_vector(3 downto 0);
        int_pldif_8g_rx_rstn_sync2wrfifo: in     vl_logic;
        int_pldif_8g_rx_sync_hdr: in     vl_logic_vector(1 downto 0);
        int_pldif_8g_rxd: in     vl_logic_vector(63 downto 0);
        int_pldif_8g_rxelecidle: in     vl_logic;
        int_pldif_8g_rxstatus: in     vl_logic_vector(2 downto 0);
        int_pldif_8g_rxvalid: in     vl_logic;
        int_pldif_8g_signal_detect_out: in     vl_logic;
        int_pldif_8g_wa_boundary: in     vl_logic_vector(4 downto 0);
        int_pldif_krfec_rx_block_lock: in     vl_logic;
        int_pldif_krfec_rx_data_status: in     vl_logic_vector(1 downto 0);
        int_pldif_krfec_rx_frame: in     vl_logic;
        int_pldif_pmaif_clkdiv_rx: in     vl_logic;
        int_pldif_pmaif_clkdiv_rx_user: in     vl_logic;
        int_pldif_pmaif_rx_data: in     vl_logic_vector(63 downto 0);
        int_pldif_pmaif_rx_prbs_done: in     vl_logic;
        int_pldif_pmaif_rx_prbs_err: in     vl_logic;
        int_pldif_pmaif_rxpll_lock: in     vl_logic;
        int_pldif_pmaif_signal_ok: in     vl_logic;
        int_pldif_usr_rst_sel: in     vl_logic;
        pld_10g_krfec_rx_clr_errblk_cnt: in     vl_logic;
        pld_10g_krfec_rx_pld_rst_n: in     vl_logic;
        pld_10g_rx_align_clr: in     vl_logic;
        pld_10g_rx_clr_ber_count: in     vl_logic;
        pld_10g_rx_rd_en: in     vl_logic;
        pld_8g_a1a2_size: in     vl_logic;
        pld_8g_bitloc_rev_en: in     vl_logic;
        pld_8g_byte_rev_en: in     vl_logic;
        pld_8g_encdt    : in     vl_logic;
        pld_8g_g3_rx_pld_rst_n: in     vl_logic;
        pld_8g_rdenable_rx: in     vl_logic;
        pld_8g_rxpolarity: in     vl_logic;
        pld_8g_wrdisable_rx: in     vl_logic;
        pld_bitslip     : in     vl_logic;
        pld_partial_reconfig: in     vl_logic;
        pld_pma_rxpma_rstb: in     vl_logic;
        pld_pmaif_rx_pld_rst_n: in     vl_logic;
        pld_pmaif_rxclkslip: in     vl_logic;
        pld_polinv_rx   : in     vl_logic;
        pld_rx_clk      : in     vl_logic;
        pld_rx_prbs_err_clr: in     vl_logic;
        pld_syncsm_en   : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        pld_8g_wa_boundary_txclk_fastreg: out    vl_logic;
        pld_8g_wa_boundary_txclk_reg: out    vl_logic;
        pld_bitslip_10g_txclk_reg: out    vl_logic;
        pld_bitslip_8g_txclk_reg: out    vl_logic;
        pld_bitslip_rxclk_parallel_loopback_reg: out    vl_logic;
        pld_bitslip_rxclk_reg: out    vl_logic;
        pld_pcs_rx_clk_out_pcsdirect_wire: out    vl_logic;
        pld_pma_rx_clk_out_10g_or_pcsdirect_wire: out    vl_logic;
        pld_pma_rx_clk_out_8g_wire: out    vl_logic;
        pld_pmaif_rx_pld_rst_n_reg: out    vl_logic;
        pld_pmaif_tx_pld_rst_n_txclk_reg: out    vl_logic;
        pld_polinv_rx_reg: out    vl_logic;
        pld_rx_clk_fifo : out    vl_logic;
        pld_rx_control_fifo: out    vl_logic;
        pld_rx_control_pcsdirect_reg: out    vl_logic;
        pld_rx_data_fifo: out    vl_logic;
        pld_rx_data_pcsdirect_reg: out    vl_logic;
        pld_rx_prbs_done_reg: out    vl_logic;
        pld_rx_prbs_done_txclk_reg: out    vl_logic;
        pld_rx_prbs_err_clr_pcsdirect_txclk_reg: out    vl_logic;
        pld_rx_prbs_err_clr_reg: out    vl_logic;
        pld_rx_prbs_err_disprbs_reg: out    vl_logic;
        pld_rx_prbs_err_pcsdirect_txclk_reg: out    vl_logic;
        pld_rx_prbs_err_reg: out    vl_logic;
        pma_rx_pma_clk_reg: out    vl_logic;
        hip_rx_ctrl     : out    vl_logic_vector(1 downto 0);
        hip_rx_data     : out    vl_logic_vector(50 downto 0);
        int_pldif_10g_rx_align_clr: out    vl_logic;
        int_pldif_10g_rx_bitslip: out    vl_logic;
        int_pldif_10g_rx_clr_ber_count: out    vl_logic;
        int_pldif_10g_rx_clr_errblk_cnt: out    vl_logic;
        int_pldif_10g_rx_control_fb: out    vl_logic_vector(19 downto 0);
        int_pldif_10g_rx_data_fb: out    vl_logic_vector(127 downto 0);
        int_pldif_10g_rx_data_valid_fb: out    vl_logic;
        int_pldif_10g_rx_pld_clk: out    vl_logic;
        int_pldif_10g_rx_pld_rst_n: out    vl_logic;
        int_pldif_10g_rx_prbs_err_clr: out    vl_logic;
        int_pldif_10g_rx_rd_en: out    vl_logic;
        int_pldif_8g_a1a2_size: out    vl_logic;
        int_pldif_8g_bitloc_rev_en: out    vl_logic;
        int_pldif_8g_bitslip: out    vl_logic;
        int_pldif_8g_byte_rev_en: out    vl_logic;
        int_pldif_8g_encdt: out    vl_logic;
        int_pldif_8g_pld_rx_clk: out    vl_logic;
        int_pldif_8g_rdenable_rx: out    vl_logic;
        int_pldif_8g_rxpolarity: out    vl_logic;
        int_pldif_8g_rxurstpcs_n: out    vl_logic;
        int_pldif_8g_syncsm_en: out    vl_logic;
        int_pldif_8g_wrdisable_rx: out    vl_logic;
        int_pldif_g3_syncsm_en: out    vl_logic;
        int_pldif_krfec_rx_clr_counters: out    vl_logic;
        int_pldif_pmaif_polinv_rx: out    vl_logic;
        int_pldif_pmaif_rx_clkslip: out    vl_logic;
        int_pldif_pmaif_rx_pld_clk: out    vl_logic;
        int_pldif_pmaif_rx_pld_rst_n: out    vl_logic;
        int_pldif_pmaif_rx_prbs_err_clr: out    vl_logic;
        int_pldif_pmaif_rxpma_rstb: out    vl_logic;
        pld_10g_krfec_rx_blk_lock: out    vl_logic;
        pld_10g_krfec_rx_diag_data_status: out    vl_logic_vector(1 downto 0);
        pld_10g_krfec_rx_frame: out    vl_logic;
        pld_10g_rx_align_val: out    vl_logic;
        pld_10g_rx_crc32_err: out    vl_logic;
        pld_10g_rx_data_valid: out    vl_logic;
        pld_10g_rx_empty: out    vl_logic;
        pld_10g_rx_fifo_del: out    vl_logic;
        pld_10g_rx_fifo_insert: out    vl_logic;
        pld_10g_rx_fifo_num: out    vl_logic_vector(4 downto 0);
        pld_10g_rx_frame_lock: out    vl_logic;
        pld_10g_rx_hi_ber: out    vl_logic;
        pld_10g_rx_oflw_err: out    vl_logic;
        pld_10g_rx_pempty: out    vl_logic;
        pld_10g_rx_pfull: out    vl_logic;
        pld_8g_a1a2_k1k2_flag: out    vl_logic_vector(3 downto 0);
        pld_8g_empty_rmf: out    vl_logic;
        pld_8g_empty_rx : out    vl_logic;
        pld_8g_full_rmf : out    vl_logic;
        pld_8g_full_rx  : out    vl_logic;
        pld_8g_rxelecidle: out    vl_logic;
        pld_8g_signal_detect_out: out    vl_logic;
        pld_8g_wa_boundary: out    vl_logic_vector(4 downto 0);
        pld_pcs_rx_clk_out: out    vl_logic;
        pld_pma_clkdiv_rx_user: out    vl_logic;
        pld_pma_rx_clk_out: out    vl_logic;
        pld_pma_signal_ok: out    vl_logic;
        pld_rx_control  : out    vl_logic_vector(19 downto 0);
        pld_rx_data     : out    vl_logic_vector(127 downto 0);
        pld_rx_prbs_done: out    vl_logic;
        pld_rx_prbs_err : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_advanced_user_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_ctrl_plane_bonding_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_fifo_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_low_latency_en_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_pma_dw_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_shared_fifo_width_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_10g_test_bus_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_ctrl_plane_bonding_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_fifo_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_hip_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_pma_dw_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_8g_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_clklow_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_ctrl_plane_bonding_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_fref_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_frequency_rules_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_func_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_hclk_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_hip_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_hrdrstctl_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_low_latency_en_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_operating_voltage : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pcs_ac_pwr_rules_en : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pcs_pair_ac_pwr_uw_per_mhz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pcs_rx_ac_pwr_uw_per_mhz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pcs_rx_pwr_scaling_clk : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_8g_refclk_dig_nonatpg_mode_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_fifo_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_pcs_refclk_dig_nonatpg_mode_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pld_rx_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pma_dw_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_pma_rx_clk_hz : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_shared_fifo_width_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_speed_grade : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_chnl_transparent_pcs_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_shared_fifo_width_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_fifo_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_g3_prot_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_g3_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_low_latency_en_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_krfec_test_bus_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pldif_hrdrstctl_en : constant is 1;
    attribute mti_svvh_generic_type of hd_pldif_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_pldif_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_channel_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_lpbk_en : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_pma_dw_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_prot_mode_rx : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_sim_mode : constant is 1;
    attribute mti_svvh_generic_type of hd_pmaif_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of pcs_rx_block_sel : constant is 1;
    attribute mti_svvh_generic_type of pcs_rx_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of pcs_rx_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pcs_rx_hip_clk_en : constant is 1;
    attribute mti_svvh_generic_type of pcs_rx_output_sel : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end twentynm_hssi_rx_pld_pcs_interface;
