`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlsw8bPP7xUJp8v6EuZQ4TVigJyKiHyFWr6omGADp1g4J2oEeEjLXC3585L4np3o
AyHSmkrPfeZw3NaPlU1ReoCpNIkFJWtqefNsWVzLDrMszx4fI6WdcLk/w1H8Wbmh
6/bD/6PxEUZKKgPTDlsiyTWHaZ0/MqBkzV0K5rgObp/7Ax7AtEmVAbFuaMBWJSwH
Z+PX+op/Eym1gvWhJWrKwWO0thf8ats47u2hwbOQPb7YbC3Wl6sHg8MbVFmGP0Hm
o3OMYG8EXiEpxx65AUH+VF8BAwFGzS6jErtlnxKm0Bsy8YuA96fJknXz/8kvfWOF
mdYzARU1DaiZ0WFXLwWOFZk77FJUQtKZGQsaLOkwfItJ/oK2WZzGlkuUS1uLvUI1
0TQSUw0lNpw0IqW92ZYFzSPZ5mq8dfYP590aZdsLApk1kpsMvAT/eM9xI1350mUF
YjGAE+ofKMPwjXr0xKk3qGY2zp/1rn3W/tjPaXvxpwgkLc/FNOkf2FIzdFmcckdc
N2VYKAvanS5oDdCp6Q0bGxyR5PzfIZfI7BqjILZnsxJ8fms79e6AQax4DD5wJPwb
a3gqn82BLGEJrHbbaQXuXztOIFvyPUy4lJLQ8Mla9rkW+8RJ9jpphonZLLThvIr0
/0CpbttdL8TASmot0wQPaaWAphY7erVQ8867ktrvnls90g43f7jxetgfl3Lp2557
lE2U24C84XL5+51sMlZfX/EDGdVmQ8RzLCwJuWnl0AXsS9NsKLAyy/hliDZGBr1Q
icje2owTEVW9+WgGaFTr/zAPq7qZZZHKoauTE0enx5D0H7RTgVGNKgMC/S1/VmUG
tv98kA+BjAO0RX+x7gLeULpGqvwVegGz189Nqg6NiCb0AYDdEDcGPpxiJI9A/h32
D6y/YxMX3v8INu77Q7seUGcTL+P5avg8NPepjh0ajRo/cRmHCWbkc4uP2JothypN
N5/r/+wp+7b3cPtgbo+OHtzK2x2cixlEg0UOAYOhT1cNWu5gtgmFV4X/P0QR0BE2
`protect END_PROTECTED
