`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3RsHkLo4DvqRgiABrPifcO2gtWIPE0CNXYLF17fMNHj9HJ4Z3Diyb9JxA8JhK/T
VUDd5uDWwsBzn+9Yv8YA6Kw0BCfjQWo+CTq/3g0dhVNyjkco1QzD/FfQpBfqZR1h
vkTb9OXKwhl7HxJ1+O1EUw46MkgFqNtuCKIXlUx01tOEB0CAn5wCDqNXnDOwiJMd
MsiA/W8SnT0aSUrxXQUEY4bt1lcgaM92/5AaBo8RlRqFxPAm28iijuNspX1RufwV
vUhPc5IyksRAGV3U6LjmtFvU2/F4ppYxld6Y8iDiSJqvzSHd0B0vTA+EA7h/XRAh
ruW3Nflra+7Z5hEAGfUYACn5L3Qpyk5IBhRf68oKmnDuw8PyolOGjnVMLqXH57UQ
3cLumjdiBiNE96sWMIdILf0GsjOMTECIOGvn0gzGu6b2xEwNv0Ybpp12iRZYOvV0
XttpDObj84GOlEetFMhsBG5fb7n4PDbmXQi9jCPh+9flqx+BsyU2ZjfiA/6Rooti
`protect END_PROTECTED
