`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLcaL53+zaSkzdh4YmxX+tLaWUJskv4/Suad2nN4D9FDVat/39SlkUdPXZ5gfs7w
k/sUPK7LPvVTLpAt1mLzB9/iy/Qhi/8dg8HX3h09gPfd26hqeyxR04LFO60pWnWJ
oHXzFC4ejwWjpDsukvy34XfPjRk6ZSoo9yd7KFM8mqc+TEkuQ/fd8zQzIRd+8ATY
1d7iKxy+WzoGCQ2OLq7cIC7d4aDf1lTk3AGPFaC33ctSqTzroU24Fbw+gq7T+afb
MDkUQ9WBvb4HZz+UAqtkkoTjKwXP3me45NaceedfhhxwNeRC0m9RpycgDGh22dlH
3g0285btlkfNea4PJ8z6rIsQfAcFUGLcd4BXo4zJlWv5VYWKOCVPTvoyra8xiA0w
`protect END_PROTECTED
