`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFsybkOTXJQsCC4085RjblMDdtb4yDZEkAiiQLrp8gh9KR82ilqbMjU5EpqB2v9M
Erm4jd/oc1RqaFDTP4DjinjkmAQ1H8tpg91voiWqwa4k4+UVE7jqm3b4yrSka6Tv
Lp/UHaryACpjKrvbhmiMw6X2MX7rTeRt8AZLCSwUwb8TfOIpZYffsdZaPRRLOXlv
lV86IV/Dof1Xvvh5i3UubDSUhKfwuKAfiPUudNDS2me2ns9wMenP/iF8KTqw4flY
Ukh+QP8eCLXSVSwKO5EeNZcSkw7h+Lb0KJRy0syPXqc27rJx1Q+IjKTlxBxbZQn7
yAUfHBZhptMvCy7iO5ShneEVjLBpcdlaEr5PvPjwl3+Z2xM4zOs9zpNWOx4ieGB8
T/Wv1Xb2bghrmkqhaIgd45IoJ1Sxgla4tNR3959kQdeo4caGHDSUxBB/xLFLE48o
zvJA3W978Ln4VQhZ9Hhn19nC38NosQztE2Qzfq29UEPhESOL51lAqgKbeptCvNQw
PdWdqxWigcLalYEqoix70wbcdomHp+3+iU0vobywA24cGibFjp3eWXfDDjv2YlAp
GrOV1IBibYrXVDwsT+5mClHc9+BBRF9PPfZgdNNf2izYgmGNRbWybm0Ngfw259r0
D2bKFkJmRXEFBCEx8B0UGm37Be+4UqzhBGxDpohSkFH0CIJ/2JRvSYI4bJdG24vA
agp2CMEkg+4oKe1+mlOybHWJoHXmu8PQXXCM+2ctCfik04aNvRlg8Lt/92yTWOCC
rf0iYTE+E0qw4+7R2fGxwBeoPOn7HFfgCsFJsaAZc4uFtX83wckAewry7Lj6ibwR
oMfelc+JAAazvQhnlhvw4eeKeRZOF0Lm8goTR/x3wBAMpdhlXaJJB+fACJDLmc9I
rLIrHDY+qZRYR307UrGZx5idj9Xj1t/gOQ9ilU+/aOqjQvlBh9xm89ZoEuZ6uPdk
zg4qORZ8t6alm3LC7Mx9eGLuowqdezhqOnKhFGGwS1Z8uBbqoMWtGPKOWULOR0/G
QqtRziQAXWEAaE73xl397cnHVpUke/N05Uf9WajEU/ElfK/2i7H2AZLhTfSYdohE
0CeIx1EG9jffXtn8p/aTMgnzqypFEmFPdkD2b7Oa9fzqSSbhhQL8rUip4q+bWzGN
GKDXFOG5/8AdmgOxiBOSuLPp2gYf62Xmfs33+LfUkoUk35d55G5lrnMiPVOd8xkR
FZLHqMqAQN7uTnvB+UlTTueOlNSXPPsnW3w2iocxeGC3Y0OGflkB8NB8gOc4rR2U
QHlM7CqTNJvzScTA4Xl6Pue8sHAzgFoWrHo9afMt6gTmLQlIOElIpvpUgAeUoHOh
lePmdNdIEzdHkCpZA1ATDbWras7eI/RRYSE29SkWsUi18co6+0RT5RBb7N+OyJnH
+rDiCoW+q96MuKvxXD3Qkl5y2kLDPg3cWtEnrFs/7CbzzHbm8dYzBhlU43kq9aDV
M7OAoh7GZ/K2tfdR2uiXgyIowPkP/4q/YPlK5Sf+7sG7LAkmQm3s4zC/6G2gfLHx
EQtZVA90NP374ifUPcS/WlkFcz/ZokIogFLVDzzfRNfpV7FGh7W732v0Y3bYfm6+
5ocaYPnVjskBB3drIIGLC9He01rt+loh/psBRzqk+xLacjSZnDcdW4a/K2HmR9vD
kR7puOOYelMki94TBVeHNx3fCbO+Z8/7Rbi06vMeUUMyVqJqxKj1H3jIVmCWosJP
xN3ATLpV6JGEvxGjN++tTDz8Qcdh3iRyOtcWUOBxVs6fZaeqa8pgPusaYQ4LtQMK
84mEgoeTisxcMnQvFnLLZNM1lDokYHBPo0k36Lir/jhX35njVZ+p3m50dK3FpwWY
oEmhgaopTfyzkUuGTWrhNak6fbFGjaTCrWMaE43wVeRxv1xDZNUc6gX0bCN5PN/R
73G58Sxl6kBlv6KUlQMPa8/L0IHZaYM2Z/THB4E8vJb0OD9yjMPF+Fx5ehS6Vkfw
HHzbX/Cv/WOvhU5HwhLe6N9O+W9sqn+uMyWPdv8HZdRBpDhnISuUhcP8og6CRCjf
Knb461u5W5x2qXAjLdsdUcuBZaGQYxAQVL+wjoQyaOIRh837PknVdxW+9paMmXEQ
vluNXR7e7BOBVB3lF78D36UBej6QwQyx32/uVtdG9oA3wscBzdhjoK3ZNSXUX2Rs
ZKO84veuauyN/YEQMc2MwcM6Ug+hVLdHDluz2TenC1C2426h5H79hA540l3xzu0t
7/s2LOIA3vwQiliSagiMnLVqyMmTaFcDnYHkdC5C6Yb4KyclP/zEHsVzPQwNmID4
zxM0aLVj2FIoTd+YLVneAdqsWPveTnv3dQmj85wAJE4jpNylWB+cV5UUc5DVjIDG
+z3tsdOC8F1Mrez2KbDHDsSb7uUGZFsrGOnewFUtMTDD8UWtTVC5EuUBQMuwq9bD
RHvBhdbI9rp/71pzLrG30lK0GfwEc3yWcuddkJLyAgm5wkKHzXa26OvaFrCAiJNf
4mAML/oj1xrEQdXKqa5oW9OaGUNbYRVZxS56PpImCR1qgLDJXBAf2CbdjACdqAkG
`protect END_PROTECTED
