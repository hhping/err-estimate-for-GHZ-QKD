`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glNFzVk5VFoZE8Md3KAb2meqO1E/hg2F/HztWcZH/uAKDig+PNddauSi67aX0ba2
LycnfiVf05fDEngU7MlLi2JUcIIxotC3gaPocwo0WrT3AQguli4KpJgOmjwSl26+
qIeU522eJv/sV7toDj6z2j9I9IwuCn7wXxwJodZC3LsS8NxSECOjVewh46EzbcBS
Ew3igbhfH4c+EQjNEwSLNS8n4pz5uFLhqDgriWmdH48hLCyvzIE/ejA03+o9C/SP
Vd4cY1cP0E3HaVQyGjHmm5WV5cosvsZYAkexdj1fYAVvT3gO4We3/PvjkIUTeG34
szO64nfm/1evRjVvV3MdrYFRRFDRWYg9+nRppOdeZZSmDbLcna9gbQI+XmkfCL2f
WNTTi/xc+VNVmjLq5xotqv05iXpn+VPkKiCGmsMaUI7ErSEcD04GVwd/GPQogKDC
emGuHJCQ15Ych5eMED/jOrPmQ30WHBqrtGPFD20SMmJaMgr5GP1C6DsM1IMl4gLP
kUMcJQtDvUmEePk1ieO9mQpbnvdynUvj6L6s4+ekyIib9wB8E61zKAfwF/2X4TQ6
m5ReHEJ7T0EU3WaE+d5D2zs29OPp0b603AG9NiDOjBgTtJ0OKEGPMJdwPVmbW1X7
X1pULPw8+skJA7utqpNnKc7vJW75Uz4jUHG4/NbtwFLBTySlxBWf3Qc53+IiNLFD
PLFg1VLzZNEPnOvADTwq2InC4D978WNcUXFK+qwvXq9ITuDDHyAutmG9e89/x5j5
M6HzBFnucuFNHm3ANZ9Kw+74bymRLb2OxBogwZVM5IiMyxznVqu2GdkqgqC0XGnU
1a0NYC5l0gp+DQvnbLXJQmaGNSgXSd1l5vnByzfH4TxOq5Y44aThlL6G+0HeRdPw
Q+7/NnHG6TfIoUkvUJjoS+HGuZcfG4fjDYoJAN9R8ucEnU5OHX+r40gSjB0VJVFk
zzpH9Ps+raIcihFXbRPWEd33CQlbyBVV3p7t9zAucbVLrhThzNw0WfThFDlDuccI
wYPeOO5Afzq1j+IzkELpjf05JHw+2T0nksnjkJPkQWq8D/EMgp/n78MJl4/O35Ou
`protect END_PROTECTED
