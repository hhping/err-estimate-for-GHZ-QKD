`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/9yNfdmQ02WOQ0ZKzZD0PyabGehBuSggtgXUHu7I77be9YZ3TmTAHxa+VquUVm8
4FuNzALsV9f+nZLu7J2Yv3Oh3ROMxK7W2wFYhOzF2jkkYaWCOGe8H5D1UybN5Slb
a/o++sGWV8zpUGOgWuWLxcNJ12Gajc9IRvwRSnDyI0GR4twsubszi3pQqML+TON3
PGq+Po7LxLRbNdGepNy5wikubNCaFcymg9ZgDduxvkzAbUtBUV98Qx1HRzcdBibn
WwzclC4ZkIw7Kg9riqCKjHOqjRAbWrLrNMnwN8pkhoH5U9sGZYHOf4MsprPHKHQg
YGQE6SZha17cMcvrBPDhLI6qOU3uedRsKhiXrqr0BXz3ZfZZeRTuEJLBmGW6bLep
Lu3i5q1+mQaq5T+KDdxf6bNXhiZs6rmBo0NwwAIv+3lZUaEqeTawuSWKNMlDmcNo
MMfMzlOgBw+xA+bI3YqDGjZsi1yNrvf2jYbg5Tp2Y8iQmr8sYyFh4k3mDb8ZM5ku
QYZlzOosSXAxU0W9PdkqHTNMWzIHXwWboo85YDRhFuBo4H8hDkduE2nueA6OjdO3
2P+bfG7dXz3zHC3gYKPYaS9I2r1BbWJRYzOGVg2TIkXR4pd4ZuZEDcaC3F/CcTFn
hox8uIxteojUdxxadLZIjVprgFl1yQnPKKe2TsYSK8dSXUEzEWT2z6xyACdYgCRP
ELnDnLTzJufMpWxdIp6ImveCipWqppbnQpUH5fC4mKwR2B/Z4bfUPIdkAMxsatwD
D+KthGg5nRJzJLfYoLYQRNFptp6KYVB0OX2wVyzzSdPMlGkgnC7ye1jXgAuR/Hz/
n+zGa5T/vphIYQMLvFSwwbffOTCbtGR6Fxec7p0Sk44Fnm8tE5bdbUoS8JHL+4cz
1SaG160voNYgkfQgRBtkHKNu6xL1tu8OTeL/t1tlFc6S3K4c3F/CUGY2rxe3z/07
`protect END_PROTECTED
