`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZyfTFvwYdu/x+5WH7QehWDgI4DY9s4HTqlMRB9yJlbNvbZ8UAL/3ggpv378GVTM
/7xjU46DtlgR5yY9tGH62s5Q+9EBPuL9PvQ8MzQz/eFVmO5wl+Sy8sRL7AZpqU1C
7xt0kcu8do31wa5+0grsdeCOEKYqRPFww93pL6ArVT/+DKZ6tQ7kjtqBRSD5oSq1
iiTWBtcYAhLonzoXIRSI7aIoSu0HUn/U5uWXLg2jML+yNpHtwbE2QSyJkz4GN1t6
u8TaU0kS1gQi3m789BAy2Biv5CEuKVCjM4tDnhi++MCbGLQ474J0ebHzh6Nd4Eco
MJTbdxVyb8tDLN6FdtJlGifYkltH4dpI0dhaaWj5B4DXnQfTpyiV7mqGiFJwSbEh
s08rKA0QV8o1aIaOcoAHE5PMKZCN2VULEokTG7/Xi1SJlxNYazM39kOSWdzAQs4W
OdXquKyoMySD5QT+ClUScGEapKFgwnBNoVpn2rWOlRJDvnz/i3qqZkFmtoRKHdpI
mNjnICcQuf+ttQCwNpg76K4HE3ycRGnA949pMUzHEM3VHBOFDSoqNzI+hNMklHUH
VaxkcaCzQ5XiaA2YyAeZElYELg7OVv6sFrQ47KvHR5BjX8zcPC1ejx+A1qF6y0AX
0MBzkgFmEdAZ2aA+kKL99I/hYZuK8r9omypHbx6l6gMigzlI/0yABRb7xPnwu7Bd
P+sMAROmka1Ha2byHqATT3g/2M/1H2XJuMRUp0XfIMf28Jz1qLNZTKoX+Ddrpj71
UWTM1FcHZSzsjXEBGeHied2jFjFMSOMRRAz9Lsjl0pvBW2V3YU+WWony0LqqSsee
1zYEnIp8bt6pMYWU9+lhEHveBbAjQOePs7vWT3LGA+I+0zh2qEWCQTDnMxm5euJ9
`protect END_PROTECTED
