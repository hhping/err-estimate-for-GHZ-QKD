`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UqYhWvT8z35EspBTXiB5hnNkn0kPGIOUxlX2btB82y5kWEkcUs0jFkrbpBax6pBk
+A6oG0LPpBAMWItlSUTKuqOeQe+zTHSI89g0nTlP35WbVu2OPwEdpu4AeWAsL/wb
jz1xSVSC5S20dsuSZoFHhEW2UmNzk3AXbMfPftwTMkORdciN6OcMasoYgAz9p3LP
9VHLiQlh8KdWUaGle7dz1+JSRfaZut2uIqhb5a7p5QeT33y6Dl/jFL8NkG2uxDNH
UpWvGUSLZ70HWbPHwVk94wILhzuSt3KdFtYaFsbN2HrySkBf95YLWg6SwzjuyYKX
tZHLFyX1iAfyyvf+Rzg1O0Q/5NzFJ5oRsMhdZaHRJdXWlFpuBUWMKJfbw8/1JbId
2IS+VhHAnD21mkFesG4DtDKk2Fwx5AsVbfHp9CGT/NXLZay2QCSS0KZg7evHJwVk
MODHT+PQ1diQHakF2Y210eQex4HCBdjkQ2iNCz2FYmk2Nea2TxmVFzDg1Qli6jgN
1gnnpJR6tTXF6kgXwGZQWOrRQW6w4ljUgLjlQDX9gt8RkIPFF7tBWMJsQsnAoXHs
e+uYlz/73J2PogJBlG8UmOtBX0/HoGfLkMopPAJ93NgwX0wJ5Zl0Lm3v0PZ/Qi3U
TQG3PczNO9T16Q5Pij/9Y8UT0wNPO+PPykwXArGavC1+lffmiUJb4O09fhsvCbRw
Ag3Johtq0fPnakn7kZDXoLRakF1AwOwWFjS5XoXutoUVvTh7hg5+K4vJlet2giyT
`protect END_PROTECTED
