`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxmHw9Pai5jF021ZkQYUn5fCah5w27kQdhIw0o5KrkJPFSAAXG19Bte0m/R/9s4+
YVicPui/z/EnOldCQQXj1k9jUTMGVS+rR+2SVavtE6U6NGq9KrcaFNW1bTlY4kpp
v6ae/7Em2A0OWuYqTgKLmb8iCU96hNscdc9iEyXfK/ND5fCln/9zGPt871Ry7uG5
f30yDbpjRUR6m3Kq3KfP8fa2jq8AHKfd15j+SHcXvK0b5Ym+SLNcKfb+mYx37ptM
71vKUEPNk0IhWdkYLayhAAlyaWfjzl0G/AElkH6nYsQ95XqrghohTYd+JtRuvvj9
FyymQRHZQr4Jew06YUpixEtYUUjievKnUSFWIz5g/0FeX6BMRkQxIWM9uzwZfArE
JSg2jD2IXTMRbQY0OJo0O5rGrDTaVUCZjlTFbZBi16lyJj9exqoYp71W086a1zRk
1y8wN3hLBnAPk83s5bKzojBT9pVg8g0eEKksLr8h1crPndbjPoaiofyAfzIi1AGa
LRFuOpY1ELfu4QFYrzlYtah9FjzSdlRzVtRemN3QQPPH/BC29aXtmPZKypoPDQAD
jYHyZ4TFGnutS9ddIUKcCTXnr+pE5UanMrh7tHalRiE=
`protect END_PROTECTED
