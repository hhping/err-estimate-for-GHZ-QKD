`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rf+1ZfFPJqzhYQvE26Olv3NbTstBbC0P+PcU8V4vx4in/GIKbybVLVtG+QyoqX0
2mKwe4RoG2g3pIWVXbpZSvlxvzCxfB96bfRXUzmKC+j+oMWJwPbg9MGJBw4QQXQh
XPDqDKuOSs4pmDYjV+H1zZlerONOdbzwciEV9Ovbp6NuFItsj2itd3Sc/9pee935
j19PuGKWfENJ86BJ00cLNuM0APjuMSPvmcbu5C7Ne07i1CcGBL7BNt3ziNlyLdFA
7JIq3n4JYNe6gc/VbMDcoU5Zp8Ace/zekoZTd59N5WfJXf0IihQ9hinrRZ3seVTl
ZqQoSXifPLex2RsMCzxzPt69xdYQcYBbzSAwIaQhJwQNZ4GR7joJtAg7/xSUVQg1
W/qSMhERaeqAKwQ1F2YRYzR8clnxnc191XFsqZPOs3JTIUCzgPu+JgCC+fk9773g
A9bd6mx3HAljp4HDRw9mj2RARvtqhn+ORAbScrXdlVJLQ+3bVtXNUXkd8SQ+sM4e
JcieKnRSJZ6Ix2gr7neAxUnB0BwoN8SeaW1K67dtk8GPBFpfAnBuFU/88Jgq6p9M
wLIlYefDHXrHAinh+cFE+7ZSLC5uukzAh9MtqdPLR/ACPKRztj65iY9MPc5E3SI4
1Yq8S8YyFchcAKzj8A1htA==
`protect END_PROTECTED
