`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KVoAeLnKGOg8L37TbDJ1GLvXpgqDdvl4E/paBNQ+I9bo5x9FZJmo30UqL28YXvt
smNAQjhlzPohTQ38+n0GF2XeWADXnox2gdgc/8Ht0AMBrECVrT6/lcoNfni9+ETO
8sbIEHFReWJd51eQYLUjwpjWRS3tGpWvlpDvr9sIF5riM+AO3+c4Z3ALK+sU1yFB
G1stB6y7SscoZbfJAGRk7stldBpMEWuwK8A0LJt3R3UBwwVL6IO495RaD3JmSBAw
NdH09GcRJzlJxUuIXuWw5AuIaHLIVp5bg+gaucAprFS3wMHnzUiPe+vq/4IteyLi
2OBE533e+UCYo2bQngKz+Wjf9RXVWxPIYRe2ukTZay2GvWnuit3VswIvAdzcmFru
5YsX31VLw2NpMW8FjVBePr935SEP0otT+AMenCAsa7SQI/TarxDtoVc5zZwdxx0+
Owby2oTXXw+n3HDfEeqQLlXUTMwmVf/fFIietaSdKWZYXy+HeUyjktwOnqPYnHAb
MdmF0VFYsdZBhTWVlAjfL7XyNm75O3Q6HZzsSogdHlgcsDSs+rTOH3bnX53ifGQG
Krj5IPezLmxOt+VSlKs3PY2VR9A1HW6dOpzvV8ep0kGoaX+nxf5fyoxnifprQB2D
CfXo5de/kXflvYVJo3peKgoJ7DtScQwwEps5Lyyd8/GJQHxMcoLUAOm6p8o+8mdB
f3Y9wZo+Uv88fYFaxo2FrRdrDDeC9EWLQZG92BsRqoFPhjC27vV8ZReSDymGiO3S
xkhPj6RkEt3U784Gs453rcxLGr3socyHU2NXoaoUY9/IYVjgAjnGnb9hNmbxfzEb
AS1GSGp9bd9BKMPn93wwxGe4gv+VDoZL/1jGU4a1LpFZZrWLs+t9e3H9UlTxdsQR
Gc4TETRm5HSfbkSv/XubeTnfF6rvssdB36dPAbJ93nhcxyJzW0S0NWim+wAhXs/g
YF63UeixWGRPj3/hRQMZ/mpsei5BKxFDwUXdgl9j/YLLBKLSCf+QeOjB5PXdQNW4
M9Di+DQxraRqDcXMN0smBwtQ3VX+X4+3EsWsE/JAnNuuTU3ALw3xbhp2zwV2Ga3R
uGggyouxu0Lc8I3Z0dfOsOdErUmlUBAahgNt9G1+gzqe617Rxv5adUJzlhxc2y2J
SEdjXmezTUCzyFzDjQFN72AaBEfmztxdK9SmzTAjtVzZG6gSVGwBBMc2QZLYTIqr
S7zM1EInA/5fJzFN2m1KDTEw7FL9FSUDNpIDPPjw5waAnW1fFPqqfMEOhYdooUoq
L7hAqSNCcW5pfI59yJyINyNtFCnbFxS3kHhWnC/Qez2lj4mlPvKO0IxcfFMDY5NQ
Z5hlmZnVR14LgBaQusRdQWtMGEFgcxrcShchmWEdzSh1fp6plao+Ka9i1D0qCdF6
cnu+gT68VwkgDfq5mmRS5vwLipuswSkLzyB55Xp6ZqyzzZOLRNBcCiymR+ZCx9YX
xDScY4h526S4xwadPGoO/mLARcXiYzSEkE6sNWCPnW8pT6vuG/O8vY/j31CBAMoO
Gr+1vGLbJPSf4IOm2WryVfIWS8phrJ9mvIYpjldMdifCN6VDc/juX6U2MjApOM5O
I4SyqAh21LHJIB0OlNm9g40qj7lk1kE6j2FE+wcm9iKCb7QSm6HAvhdx8W3yMlhc
LoyU9SYWu/1gxF1GNchH/D1FOcUp7BowNxMnWT2K8FD4NyfN1kr9rRQnhFrY4vA1
K0fqhj7LCvxPGUftRJMHnUkMU2SOqleJd7TzYz5e8pn9R1WF9ddNi2GWVz8rSOcM
eo/WVaQMK50s9uGu7TiVWyAccSHlTw24JE+Ycc1fS1LVtRiKqG6M14byA5tHSBuK
XDQI1H7pSOiatuKDlIRUN8c1OMaWD+VUdPdCCmnpkdU0Zs6gAeNRtwUu2+WO71Yb
Ycro/w2t3dnYBNpNt6PK+Du5tvhcmiiujLQq319Wrj9p7JvZaK2tKTylyjp3bxSd
P1X4xgrOUu/kms8jD5qAqQZBfYatwZBYcngDMqRJMrRzqOXCr/nk8kVfgR87s3Yd
nilPV7ctuL7U/ZLaorDElWvKyUxnomEudEO4O0NgfnyXrE4QvN39RuKlsMlWRnRP
6/1UUlXfU4eOHAy+pOI9JQyE92anJUDzAr6YBH1FC/YSNaa53Y1eGzHbInIApDa+
m2Irg/yduIFDjMQC2HUywRtc15vd0z7al6gv8A9DIj7QvVZ3y6I9gQeYIAbvYHgx
Ul6cjcC5PxfzITO3VwZbrz5wDEahosu0590kJ3+cphSw/Qv5dinx4YCWGu9Szegv
aEB+cfI1T11WntzH0cnyhIjXK+sEahoD9n36u9+BmAeE9A5JTeDsC2xTNUZs0CfG
VkREPA23YOic9MQ/C31YtS6wJXPMVdwthKecMIW9hVZpqi/3N9+SxvgoOU10WMV3
NPBfixPKDXi2Ym6fPY6Z6dDFOLoE3PLWPgBRtdvT02CDisvCzrPU6+VBacpFpcQm
kCaInBgTzw/W2UhXc94GBeIB2gsxqsbcIa08kq8t9JjSpRlW1VdcaSWT/CzKIqgu
lHQuPMN9abBlPXVigQbcDQSDCHK/COjL82qYFzZVFk8W3Ay1VrESC3JIPUo9X9xA
gAjK7SBtRnWvr7OqfdRBgrlIkHd+nuRZWlcoviaMYE70+1leu06qcE61gybiaa66
IeLTqdNF8kTO6ahfSyNVeeJnyhR8y6Xqh50SUheziWwotZH/gqajkld9M8TQ+ci6
H6gYlP3moiN+Kh5RU/OcZbOWTGsOxnzhxQza6N8u458UOJNszTtDIsGits91pGk1
+xPksNRiAzrMYPR5YPGXGQXNmJhahv3lZO4Xj30KBt8qa8LOvjHlIPEyWlAkTFwN
EfdxdQVQnJAJh5OsEIO7WsNrHM8tlQ2wVlyjPBhHnsaId6mgjoRb3MtFFNQGJ74X
pZi+XbKBstN24LJ+T+RmbVBBMr771VQbTd2yKW/HFUVInpz3rwrSUKkUy8o1WjOc
yNwOhAqnkCk498BqVoyENWHw9Wv0wgfYwImz091Fsp6y1TDhRYQD+ubZU5u4R4fK
g4a0GLzffklSxYCqoxKurfdQ3F6OH1fJgc7/wuJEkpIzM7gPF6NsXd/BxYV6Rt5V
pEuLPIZRNQPaDcGR63ZK9c9cGMdrdACQYVdJi4XHG5ZOP22dfNjCbgWfs+SIHKUV
BTntpIsiSkwIMPJFhXJP1okooddcNQHpPCEVgWIAYwkArEeA/XAqa/KVpFK3P896
YLBxQc0Ptf3IQ8P0ftGRJmI8Cs12ohTH1knUZq62Vi+x4y9RFyFMBI7srnrvxyoa
7N+vloX2KSRQQV/KpwGKLfnVIlNM1vNK81evC+kWR/gksetD7eYstwk6bT5jCWOO
hc/oC2lhsEbzimjGUF4iRjxDR4LiRfWfzsfBVehf/4XeuVH+xiqU+W1vHbf1iwOU
qL1a1mH3cmedYhNFJZavBOUgu7az6JCODYoTaXHRc+LqOKrdQubczFvLn2XNRPRW
JOw8ILULKiHkplzD0Gybx6kw2TdVHy0YI2/o0pRpqQZo76qa8jVYO0BDUtVSPXQP
EI8Ph/zCkwcbREmlZAU5FRHPGHE1rwy3i0tYqEWAf8umLn+R7bskJ4I8bOg87D6Y
cRLYgJOS1GUg7XH96d8PZkLqngXe43lM9tlZMNRZ0BTgB7Vxm8ZlWPh781kTeCEw
33fOZ0fWjWozS4I49uvQL5f7aV7dGvIx96hmLM+RHp7nryno/rzAqT86vahObjVJ
GdHL+ddOW5LwogR+J5oUNsb0zNgkqs3AQTn2VUI/ciigNVni/ROuTMtg7roxAdHx
GbCUvnjGBphVKIcsza0To2KAzn0RPneQtY2HoNR+HC7iEEdYAB9TAaPRXKFaC/z4
PzRzoxzEJ3xrCQKprI2cTxR/fDXpRGs4cbdABDbKClCADL+0HnuFJ24odRAKujXs
sh3uO6K7tZR79HrNywD8lrh7b9iJ3iRh6ZfKq2dtXuBBN/pbeOfHqNvi8Kq1Abvx
twCPgK5YRXimZCcPSGl203vCask7x8oEn7H1hKYOpymX6YNANXiOxGf9iOUKcwZy
q+Pq+ig4qKPlvZtTOCLCGbAzzVe92JsVGszk9HBGAmiY3D71tyyEGk0ovaSQAkey
Hdr+DpfawB6r42zwrZaTcn1/RmhhRce+EdD//QIsyGd1ak7HIEpSBJ7M+c+ffTMn
VhrCoPNJRbFJagSyhPm0vMQYo+pBlmOrMguGIuaDTztCerCc4bAe4b+B8CynjTcb
y+xeM0Ifj7sl/YWao+0c4VkmNll7NkgGyICiKmD/ZCrJaaOPYXOw8md00bgUNo1A
1SomKtxcfGM8FW1B9Tw6aPi+AU5wKN33OuXsad7RqonBNBCZDdqkbi9S6/snWPUU
FF8VVR1l06kgbaeII1eytnH71kRzHex1WYjGG7Npyb9jMY5ZGPUePx9UIXcIOl0m
HwpU88Kiprk87ORJFuvY8x7Jj7WbarucwK/7J0yhpffQChmpOFt4Xd5u3uVonY//
0si7GdjwXwUyA9DsC84x0g==
`protect END_PROTECTED
