`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxCoFzgODRwdL6nuyDoBTMbq5w963mV0y2IpXL6IDmhlgIa7F95QFlz5BZt0PmHG
/uXZZC36Cug9ZkBEOaKBbYSUChtSHC20e3ZWKycTQGAc0NP7k565bcNsjOeQfYOf
2qKPJMZIMQEtxukSw57a5y5ZgG1uKgSN1LorLlYOCWe413JtWJqDAlXkBkwMlp3t
m3N5zFlQ6Qls+LLHbAtkDyyi35uS6lr7+W1tbLEgjmvF6g8UzyBV4KuPFj7JFOYc
XppmN7CeAsZwQuTSw+xgmtQcC3AAHVsWe8WuRymBY4HfsfQPtlQZFgCWE3Pj2Xr5
izNSG9U10Vc2BOSSRuSEX61SsDn66O2apcfNwBd6hWs=
`protect END_PROTECTED
