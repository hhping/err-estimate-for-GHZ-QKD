`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xV/logbYpuDmgDbQyaEKbJVKgTpfn6PnWFe2i7anwVjh17nDn32092cndgIi4lfb
ZCBcyU6rcj7z2BSO6NmF2Jqi9KIlIhY72vToowa6pN71NrqUwsdG3rgEztLJMHaY
eketCtop1ONh465NV2dgwIoI08swC97dksghaLTuiO+ZPKemDbYe4/+I3JQLC8kK
5HyCq0y3N9v9nYnZSOVBMid8GNM1ETqHYAI743FXaH70s6pXEwgePwcTNp+ldlSZ
fNfEy52tgybCiD1jK4aF7DIImz9SYG0Ltj6/H00mkhBuNKBM4gtk4L+UnTFZu7n0
qdl7G/cowH9SRsBSiPR32TnMhM9SYap4EFV/vEIfUPLsrGxIACa/qPEPg3Ih19HG
9K02TDBdAY0TUwdX25pgwx2LbPDvD0wMfLQuBBsqeFRZmqG22mx5/cfJVfHWIZ0k
9z51MYS9DSNkwGLEWh0cdwWS9X8JEg6VbQAEMKp0wm1ZzLgfhopbSyVU1DCek+d3
2AfMFf5tq2M/4fs5Ie1/bW1ii6SKt5ly4Dy1W+xOu10dQXmjgML8TuRQdbgFY6f2
H+7c87eb0SOzDJldAATwbw8gg1DiFQv90Uv/ysOjfKN0neiubKVI/2ZW/5RxcQmp
3wld3gjNnazbeXkBZcyngRLuzBPYv1l/e/ahi+37dZ0=
`protect END_PROTECTED
