`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFerODVh1XYJYJNLWAjuMyqz6BgysaPODGnyhAP9YIoayjrP3H+9I77qFiIXtB15
yXyUaYIf43+RtCs9kB2hE8BxkAnqCM9mVtf/hWEKRQYX2i59pA5BM8SS2130wjA2
tay+eqk//IbAUog70f7rg/OntAVlrloQEn2hrCvlEu4=
`protect END_PROTECTED
