`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjhDM0U/OFHJtG3vW2G1wXosmBSqmsgAMIxeFimOYXio2/OGXNPld1iYMQOb3DQL
J8MosZlpDbvKJfSobT0R+Jpt+cz8e+VOpGVd6i2DLFLP5shJylKTuhixd01MB4YA
gMR7QSbVS/BEaUgoTBXTTDFDJon+MtCfQ7Llie9tvSttp2vgmbR9TYfh5pT11VM0
7Gr2fD+FEwD4JKsptSk6ze+dwtZp1T8aOQt4MHpi17pOuUZrZvZRbqR4PgJm/D4e
ko7gnAEBnlDHAXE/Tv/UscZheM5TyhY+f66pwkIyFAitPm/80RwcWwk8Uc423iTk
wHQigqBYtBbZMDf52VpIzrr9Qetkpoz/+HvGl/XA3gmUztsoEeD+SlHv3vL9Mtcb
EM2gOisn8TySOmh8a6pZnlfOVPEUw03M+jPtR7Wvda7ZFUnEhG3XYfXW9RqXQOoe
DRR4wBsnMagTnPRgyraS5B8sHJXFCI9o52XTKkZsKEJnuuNRoVPAELQWLVjgfjY9
uAliMkXblLCVTTp4HNQ/zLrzLFb1txXez9BBVa3W5AOJmOEnjxhocxCPJkKMJsY8
9Vy6IjqEkEPpi4R5MOlzKcArV14zxLo/PFUst2i0r5S1deMYP13OBz7fwcOGFihG
IUpTToGL6wkwu3CGPU5+OGoqH0FVhaeX7H2U+foWpXN8r6fSMgpQxr9x+YVp8aw+
VYWWyQqfa7MCz5CMgyxmdDNx29Bss+aYvQz9/cpq/iUMPKNDxOXBm4MhEPWc+tIJ
foHEJwPi+86vwM5ALS3e0r7o+WondPzYsNUVI7ChFJKHUKcOuW0v5ZLPxBmjemL0
v8Xy0+aJD/5dPX5R8Yi6Eg0scDW8QcT/dlFsSpQ8lXLTTWQh0Bl1Sp8mEy8wKBuB
D/pmpOs7g1Rq1n952pzNWtg91fx3TKsDmj8oMRnU7FlRcyA4CtUJGTrcKF+ipxQu
vHPtjUz8tnZSI6S2aefiRfoShKfunteHa2BqsvF4ZFEUmIOI4G//ruHwSUCkSmUl
OROfuFAhx1rWsE+uZuaztt42pCeXJcvZnNaGswHy5rDqR4+9wG3mmV5Kh6v74lne
ZYoAwzzOvMgv0ZRhTSgttlL79P2vJnsoe1fsy151OPddSHLqY0i7a5HYNPcu0oG8
A5ZrFcVyoE61Ycbhq6pZ3PyDCYEvYGGeJLzL7xKStpOeL44qm5RVYpt7sy510lI9
NqNR2GaMau88eKO8rTU8AbVle/oOl/vMoMh986gyabIJr1oD4rmmfTID/3Fe8nxh
hIXESrJO0ZaAy/7yymEWZdZUFe0G9jXAdDjDI0FxPFzymasnY7uibqPEAZejchou
z+pcSEYHY66vzA+nQjXH/gQhJSqUH7f8ULzSEXYQ/P7bXukl5aV/W3/UUWu+yg3G
b+Mx/KwxKorKbv0MvC2uGFtZ8zpo4w25E3sANXyEDLKCDJFSEmJQfgg2gUiCfsCf
h2Wsexiu9msoaArWVDKXWub1cwUQlkJm4QmIVbC6bMmjvuk9pvUm//WVvbTa+e1o
BEGV2b7FWllwnjH9gv8042RGla99yDK17KmgQP2gpVgwgJUb6IjclAKK5eiv/iBh
oR8/27lkwAWxmzIZrapyaKWQysbGauqhpKngARH3EZZpwcX8mBxyxd0J8ma9/8/j
LBhcHyvaVCO5hl3NXKClwxoq31XocHUnr23EDdVaJYeVyX0M4zjzCFGBeCxiThfa
sSt7UhhTH/6WrbKXbMRirTuBZ144kNGSdgJI/jDmgLZ1s/jzj4tha0rlRExLQfe4
0wvSMbwhuqjMTaDMDDglnZINWqYK+m81h4cVIogD4q6nQvJ7RJjWqARrJDWscj/K
EWO/bcL2xIl/hsOckC05LcufH7I1oFqkmITIQmoSSaypnb1jZrJo/QFZl+ij1PqK
o9zKaeAQO2NP2zdX1MItni1dVp/p6J0X6dT7zjQ+qtxtK2HXO7NsCKmRlrvtGAXT
18E4l2KcObEpZ9Go0TyXeXz37mjoxFg+SebWB+nbhRh/bJeLqLyIzDeBEY0EAKX7
p8ZqTQfXdeAzAmIOAE5OPpQv7PJwbGpEFBJuAG5usu539bnyu8GHai1S+4LZDILi
0i79bAVqo7f9tJlAYFLoImqzlyh2OTG6LYk+zDcEm6hwu7jM1grTagPte2D4cF6X
rTRjD8Srrn5N+hWvIBzc5YcCSVebKJb6WC0pn7xoB/+EryKDNM9yikD2FcNwkZmg
nd6lbmFZIZ4ENuiKsRQnNOc5SEGI6RIa6fIXS1tnMwB1myd9nTHCM4tdZkMfz+S6
so/b9fC7+oD1NHzcc8XVQfvY6pJmgr5pAcDg18Bx1TjVA93Lj7ZDClHWDGTPI0uc
KiOglAjjAiito72J6GsNZ8fjJrqIWn6k0cH4Er+d4Bppwb73MqiDDlLPhi0YwVWK
MPLtiPyDK7tJW9e/yGSg45oRXzCrDPj9GEXD+XeoHVfziCnYjix4hG3XjIva9akl
7B5Q1+KrPEw68Akn7F2F+ponPyDGZVku8BeCCp35EyEkAO7TeLo8qcDHSh0ecHKt
XVbfxxzkrrjoBnFNaGG7KM+7AlkB9ekqOO2ZbpO3RC7sdoUfb1i9nwa8n2CNYQZh
KicDqm6c7r+UG9Z2ttX1n+m7Gll6BBwu2ddedTwl2+pcrtzgcTqc3GcNhcpXcv6A
wo57gyVxNn16JJ3KUhjl/HfYWjD62MeN12qlc9yUr/Z/P9IA8NYSW3stk7BYKsL4
HKrCh+9oTm6L4vAC96bauUT0lv+Q0n1qmWyTf6xyhzitr4dHJcN+D/0U9ceN2J10
r890Z6DXfutq4TN6CHvOjRsKto8cV8cxjWfdTYmb01gyRe0vVMsZdherq6dzDQTk
IAxcBv/EEXsPzsAHFy0w3OG6sD+aXGKB9Y74nHPBXQcNlxaUr++Y0xKkQ2ILBR4G
KZ8Ov0tEHDiXuX7jGiGK/NMMu6fkkYIbuWykhwbtGy65Rel+2spkF1akWpyO3+rK
4xLINib7bOcELi4p/eL7jYQH0uLHP7yXqylaVH02SIGRftIrqflamg9CVaaECMi3
dGwSouMnz2o2Wg9tvR5rxqs+wgBvrmmmF6n5EhwkHQrNb8RoUk0i17yom13SxsKj
gL+gyaDNlxZSoTdovVIBGv8lncjqK9T1l/WSNYu6PTBmCd8N0AL83mhVC9SI8yEm
brbAxSMeQCg5vkmD4W5E49zqqFTEqI88bBCv80SiB3TTNkE8e4vR+tgecgHDRQWR
RV1jLFt4wBoFVINYaWZqHMVV5OS1Qw5oT9tZDYXMTxorJkYH4oKmBqZscWSi8M5h
4A2WAwBNFGINF3XHA+gIHQspikbJmIueeBo4BT9PmH5Aw+OjGcEWRcY3jOijf7tx
aElJIMJzw6Y6vp/wa1JGcb68iW1lAa0gKFoX8OvJRmKJfGgep8M8EHCHsGJ/gkwx
m+0VmjVc0i14ePSHvh4s2Myw3iyrbTtu71jY49uEfVjJamIRHk7LmrwNUdhxQgFM
LaCgdtt74XqWwVOiik+XHfkHW+OiRv2LtDAWJ6y1XM53tHqVf2jFeVUic6h1vtDM
9mWCux+hZr81Ty8qoFDVpTUZ1VHZoof5R3KjTCfwuKmatw+khNMiqozfXoTZaeDo
kpbPoiv+2l1WKaHXTegD2wwW6P0i7ENtpQ7YSXKovlVz1f5+XqYJx36sGr/qXpdW
hN3izAHXcQxIgOuE49qxmZH8C6RVz6scRXZEB3rnT5Lpj5P1U2nf+dedbMIJsoDY
LCnyLVok+3kzuQ6blgmqAKY5wZoEjEoRSdI6eE/1gnomZbedi5EPRXLmU4pjH2dR
+Q5ZxRHhUCQ0JlgN7zD3FkN/B3oqTJNlKG36YqSXUSFwParA93AUtX+lL6JbFSGI
JE3bi3D8NhLuyhMT/7Cr38TlhtAqS6vy3gUKaWxjTXmAeBhyYU79jJcx2WHmMJNr
AkFMat/4cNQaiVfE8qOvmzDnrSoG8LzBLqIj6TQwZSKuU5n6xOX16+ebXm2DvjOE
AuCXyUw8f7/BcoMIqH+f7hbkTmK4K2s9a4LNY6smo6hEZrOoym5SXCEm7xD782LE
IDSBOTn+/Qi00ZQA+R1qhdn/YW/ET4gqJXGIEnlZNO6MJrfyQDdpf5jfMrvPK+/T
3pws8yMroAFV7XsTpYztpZo7WN5FM0bKiU1kUQNw6K55qWrt25w584fn7CZrb38f
npNWpsQFXuRTHhMZ0PpOb3CSpfrV0PA10z04oMDMUpVLoGrL8akkUvC0yJ9Gt28C
ow74LolxNsf+vD7EsPFJp2JWNZK8ENk2HkLeV2eowkbVTmTOoBQyzK4dY5LpYOGd
fjBojQFvu6Pv3OQ8G7e3U67EkH1KB3Fj4Y0Qo5slkrdKXEm6ItXn8vesV/ePyssi
mi0DzqP3Xl9NMBczXPbeoE4r9UiVdjkvS9Xf5Wjo/XdI790gqkV2rl9AW12rFA1p
eZUCT5svS0py2/Z0kAi8MK97xhA/S72tj4OGBtGVoQ2mCIz60N6hqP08nrewoQGj
UC28+R9ATt8IGWq4rOgAbpBy0fhw5QB16Gk5Iu2JVm8dncsZOuLTi73N3/VRc0Bn
8Z/mpQdeWJv6Oqxekunsb2+36nq8aM8Lmjec0muuLCJq88ADLv24zywB1fdOCLe3
Y0BHzoS1kwxEA31NGidrcxD40QIFB1J0TWzsore4SX6HkH9PQC9LCJpwCKB4RQ+e
arsKw4XuQNDpTSjCNzsfQYKuBJkhjR+Ut9A++TBEhdLZpO82G7fcDSiotCZ/PCf1
YXUpFRbunEXiryjvy2QET9WHLdg5GKCxC3M1vGFdRn3bLLJWcWFqnQNErgimCB0c
jESIRACtaJZ/rumgZNMyO6lVMPQZicCSJJI9Saf66gzy4ERwIWnURgnu0pSEYMKx
FyO8fUBWQ/wuoK20TFt2IgV3i839G1IA7ADMILM/+g70Em5GjkxVB4nKdSG1hh6t
4s0z04iKZediwqooecJYGPc4IVYfkZpPwqIXuHp353384mkq7U0SBuQt+lG2jbjR
SCy2MRZPis5/hWEgZtIaXtPt3rypv/FJAROpB5sXhaM03KLwigPU/E3KyYrOG7jo
KLGrRqhkMrJiG8eH2J360c6YkzAiedKX52SJEUL/eBCzliC0AXpdZD5R9o6IVNh5
qgL259DwpuXGRcPZ3ltMJ84GGkgiT/Z0zGU30/so22TzYBYOqc61HqMOZUdP6Rcj
cehCLX8jjMWUIULwgQbzVsBPf8lrGeJK3HKVJN2tMDy7ASR4IMyKQdXYwCaRBs5J
zFJOk466dTiLC0b8uCQ0ytYC9aPuHmXf0Lo5jksXv7QygoSfphqiKPHunaCMavdV
NuIgIxMgbmetGHHDn763Bk8CFKPspW5jPTQK8H3KqB2jBFCb9NlliTRST0aUNIQV
3sqtxqoVAWI7IHMPdd8/8uSI2+d4EM0N7IsE0WYNji4MSea6ELQ4KWlGDzbuvXs8
iuUQyuZtCKLWzzURoF0O1iLQLA6M6RtKU5Vz7opUsKDslv2KjNOonBbDEks0nT/I
lCJmZCqap+Zv0AtMBgVm2cxBIXm74oOFX+9/KK3Tg2i3uuO8srO8DFDIoZ3vfpdl
pNTlxMpCxwDUcc6aa62pAeu5sLKXAYkppsQNRQ4hApX8P8vp1JeZASHDdlx1OL+g
exay4Y3jSzBjkFXepr2DC4+uA7szCvsxFrVmxkClGx6xMUJs/Dq9cNacgL3IzLHX
W5n5YCxHpg8AsbUqXzeVwVv/nJbTCy0VR5CooF1CI9RDeNpIKA9dJoaKyZZORH9k
ydo8hyVMgfy2rDP6k1FPb8drvFOC+M1UYhrTZ+O4e3MdK1u5C22VinVitRK0vBhg
N2zMfIRX1oJ3jaUb93EYpAgH5pDtMCR138q9AJs4JM1xrYYoeA7tvm0nBn6OV1IZ
xVS7mdoDGlE+b3fckpz/l9iF4u7eoBRuksymgIzmOS/eXpdQHzBxTITlwwmxrJpR
sX6p5k0ZPCuABWrnc6jllyrCIHIsvg9U9OLFDTVVatxhXCcmBy5zfGFPB7YgVoTn
IIPX2D68Tk0QQvtc8kxqVpmW71Oh0xqX+uqlvDNKuT29zKyL9hjeWDGsc7W3eptg
x5mUzM690sf1CoDDhMh6QiYjfj+UrT/aWlY6ZHKDqmbyORoB/H3G5qOGilv7M8yb
9A2uyksOHgZxR4fP+5PaYBpX/Fvn4O3SOMimB/cpLV4N805Z8pxZy31iqsp5IEHi
pEJVZwu4T4gu5frfycoyJLWPamKRnJeQ+8o45svqdTfbPhq4ssEKMyjnrgNcuR/Q
Bahlx3zfOoeiMjsdnBQH1QDzp3it5Uxmw55uS+YA8bz6Bzh99vInGFW4V5GtyeVE
ubIna3YZgHc2d3PaPFzSknEDnBbbIsDYtSl3jG58tGIKzLQlTCf+qE7IIVBMMnCu
g0UjdSQEE6tM88/RrnSsSOUgXR/MPbwSvvHXd06WpFHSkFnsh0p/wId+sdRvPpkm
Bqu2scO2Murfe6B2b+zhKzOHZWcE02lTSTX0oPshQNNlfqYTHKCa57p6jSzkmeKu
bCRXypkkct9ACofq4NP5+NLAjLComQR3At7DKBnJH/eTrHBEIMQ/UfNh/d6hIp3F
sIo1yZaH1y+JU0QGTFEKLyP2K1r8PG818v720KQn3Rb+QWK0AOlqW+UaMyifh0lJ
crDhqA9Y4LJ+ub1fDhkQN0+Vb5XV2jGqkI7YqaQ6YXzU46qdBxRmo+4NSTxO6Yr6
IbedPJqHCtm/Op0viO19wphlGWO5dRiNGBunFeI3Bl2IZ4tocRN1+fH19yAWMvob
D7x4HwWxbB3li6hcmuYzrMn4CA3rXQH33CowghaKFvw7Ipm3XCHdcBlzGfkjT71T
67rsF68hoCGU7lbQ9i8+Qcfu1uCjeMcn4rfqvAZnrQOBJln4Wvo7nAH+Y1KQH+Af
KejNugT3GZImYslxdR2gEi4FdaDRXQ5dNhjMR6IePoZ0HYZpbuHIeU5pv00IA+Go
naW0IVQUYRQHmsDgNVAd7G6fG2bf+8Ov8mGeXrSX9vFn91y0qP1JH8VtCPpXsDFp
yFMBK0Yn+Q491JbTg0uuV5rnX2hvGCYPyhkB9GdAADx+EBvyfxtNaRMtIOKZySek
alYnbuGOSGukFbGyu2YFUwmGeFd+wixvX67G37zCvdhljr9/i2hEM9FTpeONLyy4
3AcAsNssZMhLFLQ90BPIhyj0nA9jRp8cg2iht8+Yz9PDZGzsG1KS7AyL0VD98HZI
e2GaSFqpbp/T721s1E4ob1Nt+5YiamuDVmB62nb2xzjVOYVZllRgNj01E2bBzTGj
0SJQkvrQJKlZRQ+tBT8XmngmFVlUgne6xWbWl5/wi5i40bBCBbSAEo8aB0hqGRJd
24Z5igfz7QMJoY2DNZc2onHdVqMet4V+lIvTFr94zTtuP6gr2vHLilGuFrQffHlO
VRWIN9U+jXksw6dnLeSged4FiItQGFwqYRPhfAQKpyujOtT/cz7fVQm5ZkgSocq/
UdpK/WrWBQuBc59lvPIpJBDAXexep19K2HmvyaIAXTucjtwy3OdgXxi8AEIZdw0n
c0cQ8cO+zN96r8wuLN1kc4jdWSGYKvZ8MDGRSWueNpx0eCOY3qpX9tqgSiVnV+a5
6MM+IlEeFSAnKdMV/SakOfViwPg59N9j5k3g201EQX8vtS+jNn7cXXx57zGbLd/p
DIRMs9NvIRD35dZwpqA6SNZxs55cxDF3fs8lc2/0Nf+HUrky2lsjrVZAQoSfCcVx
nlbIZKSdsZW9UOSl4UgIVggVBFs8qKxKDKuhBrTuCmtNqzuYfyHvvCL0J9tm4FkQ
MbL5obC6ETSMm4XPuGF2HNxqinYNINVVS7qW5fNASC7YBOtZSAevcwQxZG/e9/oR
fCl0vB8zSNmooZlOQpQIwJag/faVQK+QMK+eHL86/l5E06SsxjCjBAJ9eiKysSGr
axxbhTpFc/Zy3vX5EVxg+8YolPm2vh0wd9BkwxjQoW4SwpJZU1rmnXpmB+fmVwly
Ox0h0aeN1QiDxjKZONM/rGc4OYnGbNOG6WyrnISYIwIfZKEoqm3cu6uLZklUX4a3
5r9rPCV2y2sBDs2AgDdNX32mpgCX8PFuNPaDQSEB3fuY+rT3qQIfgr9jL6QjxpSK
Vo/yxxSsZHZJ1IXFuDmY8IuBre94IOp3GWsaqkV8S+y3rOaGv52feumh+82jtdAN
FEonOAwKW8E4FKtVBk+rfNvKVGfsjp3IHaWBHZSPQVfwX4pEWeu4ZV0kXQ5c348x
9pJhrDjuvbmWv0Mf//5RJkSe5kmp+Ug+C616kaUsQqFWrnc2r90gIOEkINz9myuq
+xmeukc7IgcRNt5PMQeKAe/+ZabkxHvsrQeXsXq+O1O2ZIT/1dHsXo1BcmqeND+k
OLbsAVHahrBVF8nrdSf4B00OmENh3TXWow2w8R8MGaXKOhXxC+gqgJ4pKxTj1f3Z
xndxDL+DxMOh2rUO4FavT5TJS4C+waxPM4AGzvBD+ATGDx3hZZGfIfYbOCH2ZOAN
j16KdI75wFBioUhl3vUw+m0Seifj/hS4OTIp4lKpPKtDV21A36jVRaUUSqu8FsNX
jDiz2eBQ68XEDJMH06p6EwOWn94WMwvud4iMn4kaR29tK8p3M0GEGxaSMmvpop5H
tmUx+iFY5YGkvNLa4ORWZnWDrOl01N7B0QTftgOBfJeETr+BRzXvXoaABQO9EgGr
tSi/4SWXkGSwn8K5QwcXFzsuFxwriClqfBjk5RsV+38xyg0NX92JURdvH3Fb7yJj
NMLghfTqYrM5P0PNPsUYsq9epNAeJjjeNk4mP1CgrJOVaQSYGsJMEBIuhBYVeyff
tmzyi2efhvU1OB6EE3qjTXmIqtKBTSwwaRgBJi3yTaxGdyWbRIwSt02ZRLu+SAA8
ZhmUPUk798k4RX0qKU8kiji5ztf9rntJ76EeXpPyZN9wcpxLvs0XHJ2O5h4lvHGX
oGLO3QCc1D5EWoUiuT4Mo39p6RkoT23lC1mExSYeknEGifGXJ4oW8aYOeJYi5EbK
c5tullS81YKyrzhQZSbhLcaal9P8tn4P+T8xssb5kIc/onPo28Y8BUp23S9cZZim
ag4+aNpqugaVdj0vQeEq2ByU+GGU4qwog+pUj0Hy2l7usfxszC2ubX4lPE0Ywuum
OICzyIuBs+rMcc27v+oWRp2b22Uvkqq6GYOoMVcan4S7p1B9KCZMCIZ32dLKKA+4
XBPo4zxCTE0BRjYlHM1UJ+y2vqgrDSWcfyrDnrTe783gljrPxN6FRjYgFioYIRFc
EXfJuP2BYAMVcZkO15s//ioxAqCSteBNsTGMQjdP3ZvSPVxIcldenmadnVtEvXfi
f1yB/5qm9RMwMpVk9OZ54GXcwHoU7mgjiWg5Dh4f3KTjJ5AmNOL+enuMI0KJ9EfY
dv5eyLTJfnuQPHsoJVxQCkmZS1ybiteSMxDWOny6sXiFV8hY11f/kyhrKF/QTsOA
pBa9ehtw+l+czo6f6nKGCetafNm69xINexDpDJwwE93KuCqOR+N3YOKzjeuYi2W7
aOfv7zxa/q3S+sOpvXc4qsJRWwlkdnAX69lx46u6iEPZSL+b8XH/hmSqcmXKdnOh
hOrELjCsa1dXRAK3iq2OzA0tIXkRtN2irUFPWtB7686d3gdUSTAcYKjNBLxYG1fw
oEtMwn0S5B2fz2DlUJpfBOObk/kIf7fHBwXTUO/4W114xaV3oANirF9ipxIlHV3y
Hac2TCkAzta54d5lB2bRURDUCByRxP9QRTj6/+lCOBabSd/EVwrqeJlzvLi3Kad3
bJYbnQJI1eLARdJ5M0avgrhwEuZesj87LTcqqWf+u63kAD+27H01nv7DEhjaMRsn
wY9g45BWxuPx6K+ULhnmxUntWRb2h2nqBIfci1OFTQfK9odYtcDBz4qvZ0FV2rRd
Ea33oWYZFiVT6tSraS1zkY/dWOu8dBIzzw78+KLM9+fMBVPVXVDKDu3H9B6cx4N7
51230hZPK0dEcP1vqbEbaBkaZCBTlyzDMR6cM3iwok1jZeG/5UC4psC6/NKad/Gz
fMMQ1qSJyIqF7EFg6Yh0glN6M4iCawU3iuNObuv0MfM5YqiV8vofTkqBey8Sux8g
QpunkRNKvPnCVpxx09SUZYFK2nksLLXOsbAVpgC5tboOB6x09KXmqVUtIXaRuJ9s
88hp7UwtOSb+RNtfhN4FxMOHCxVFLhoT1c3g3fozHUIWmBQJRjadq8eBuGkfQH+3
pmH//8nKEnGSBFk8QwkfLKf53veR/rKxO/IMeMSHMqlPYToNnJkjd6quBg6xJz5C
OyILTsGXMszA/lI5TbHon1Kk6y5AURSXIndOyrM7CQPjdotnMXIzdBV2L68gt726
yI1O7zWdqNpec0kWC2fi+VwEoaLa8lqG7YEDFwAAG5Nsp+SuOo2v6JEJb7uF9Ra8
p4Zpi2wivumSNdsEj9PxUsjLmB4iu0YAcuzABeip9pNDI8m/k6Co6ujhliNfxKPB
Ooe0wct6Gt7ppv4WLeLJFzHXKbjDTHE1nWrY1TGwpZJSKA5APn4Wqvaxu7LwL2fI
CUx8M9gdKB/+1xQnilhAmwdJbNLHLxlOthVFY2vDs9/rxonWb91jZRQ6uh6k95K6
AVHYRKV6B52jhOy8Vr5K9AWCf30+QyTRPO9Q5S6pU/s4l6X1y1RGiim4JIeTIZIq
4u4ra+Q5QsbvIJxkjjRs+ZZziXy53I5Ilm8WtU/u7HJOW6fEG1/4LaS9rmA1vaM+
eeDUsBWGF2EZ5S0JQBRYrLAM0bND8G8npQaNf50bkawjeAeUyFwb4k04LjekS/cd
ljNc952kTJTjIUAiRRd2svGm9CUDOnYPEPSyC/LSBJlRTORcDS1rCC0DLIYFSU8n
hDgmy4hDStiPFMWQQ+tWl7NuV3B3hXMxpWKkDi5VnmbmSmVCBz1D7Lp1v0w3jOm0
6817N49lTWyld8XK+efFi1vLFeURflZkrnfDeKz9ggfUox1K6X0oQu5VATtxdEpI
DBRYQuKePovP+PJgYtZx03QhnT7qNnMXOOp2pyO07ZU7xbqO5uooL+cv30F2Ickn
Pe1ydQAVjTuiqAAnU34ZzyLPEW83EdLjGpJOn+dqNWi8z59n1KpHh7SzuHLOHZnQ
sCyBKSTeJrGoN14j8UYB8Mp3+v1rCMbPA2xicfyTR2/ttJe26DdT9trZOrG3to02
ZeH/aRkJNJekT9qa+BPCD2UKkz/RjPkWaCMaBOrvjnWTSKeUiq2XVoUzM6IfDwCK
0aoc0udjv+HZWiE403P90V7y9Kjc3pVG/+koRCdRbdXifLXu3iL7ldoWCOG00+Jh
yNL1NbcZZKHDmD4NZV9w9FwrU23iiqJqxhni3Sfo2g57T6LDF1wVflVA4SCcpTOo
I+OdHoVh2BdpfRokpG6+YM8+9RJrMwsGZvLSutDm8sBDKjyu6A4/gCNMS/Lht1Se
DtyXOyJIuUxRXwBpcoyKhLvx+7CTwuOO5aOqpZtlIAIt/XawjpWPjEYuC6YlC/Nw
RS2LNHrkv4ZYBhnaNyG00QW40lOLwXHuxEjDjNQ9pPUmgfbFO7DOmqf+kgBCi3wg
Uis2HSWXxWHm7dCndBGcjB7uxaqFrVGDbQxj8fNJqz3w6svWyHxNxcjEL3ysvq1b
autxscAsURb/M5YYI3lKfllAuQ8mjt8zdwn1UH2K4Aix9mO6iJwOGZV8h8Gc+r8c
f7tg6HSo0exZMsl/knA3px1qBJsfnVinGg+Q6E5f8u9KtqDLYQQbunTYcKNH1I0Y
SRSe95IdszIEIopcPEppy6EDqMD9CPUkSdyQdGcU5lWj8UZFwCQRpZuUPRdr/BLk
wLRelHeVcqSR2dRTZ1M8PvAjAovpu9trXPEnxqLp0qwCseFBCCs+njtMwFduMbtE
bGEbd9Yp01q1E7sSjExhSju7wq951jThtVCJx2ksY0ri3gwAJLhbiKYnRA9Tdz06
HycSbuMtRgIf2NzupgvdjCTCV1IVjxgL6P2CD6ozmUOEgXGbp6GNEIjGpTmNy3x6
WacxMBa87DXSf6XOU7yLk9MVXmQHLk2N33ZmmoT4BS9udayIjKtlwJYc9nCFwbop
71wtlNPjjJLFZoEeKR2773B3ljLN4oZBZfxgbWDiLyzeuosOoiL14yE3wNggewJN
qCT0Nwg91EIPOxNeZ1jidrpYbWAGUvDg3SO04lZAFKD2j/o4sH9YHzzlBPNMMu4V
QomnJqKM8UQu4LSp41HaMGaHFpLI9yS5/NUwy/2Bspz1S9DcbbxBwxpu0OzRrvfu
2AboaZpuPwPkgeChzLVzsuhxRIRhmNh7H4ChXnaaCSiFjcgJDzPcCcVs5wgG6K9t
NVzYUj4Duh9fRIuVrTv91xz9EUgKbYn7GUtBOcfradKC5h1ThPd7OGn8MFzy+bEA
lyTUVmHsKHpx0XxyLaFknfVhvbLIGv6jOi18c4MMyJhKr2RFB6Xr8f8uVyYz/5yw
UExjXWKVvfyUk8jSVKeOVXEE27loc0UjIfDsdlnnQJcFxCg9mI2LWJJ50ytXRaqu
lKiKcegzATnCysjn749L1IFxRnf1/6GjfBBDrGews4hCs+39tGIvt/FtsZkNWQgR
TGeKBzJ7miraoiJEwLek6H2ilrMnHM7/yGzhJ9Ujd9ZiLrZKkcsuBGj71sI4rEGF
rFzZVe5p0d8DuQf22Umlmk3frQsiqN5MuEZ0s7+RtXU1LgzSkIwGIGz7/lHjzoPX
aJrlhEzVj175xubhPbfT53U6EfVV6RjMwElv2a0bdHUxAYc+Un/mDxtHhOUt/SYu
bSUGzs2bN41qWvqcSo831pnUviRLQfN7Wu0D7BhPu2gaeep73W1IjnDcKYpcq5aq
1HB6yx1ZHU524t1eVG5l5tdDKSY7OO4BlshDVD12LNfWu2YR9SiklYFEWnDVzrsf
ZyNseE8zYNqIKIca9h8Ms5+eT8+IT/5zUKF2B14lNnnK5To2v0yIaNiEM6s/YF9J
qJhy3vvKYQbD0urjyRw4YV9DDVS1fn3k1wHPipboIPljHIj1CIwUPsmkwUmrCEEg
YjzLmMz0+srM3QMiptjhBNKXnsGBpkqPtecge8jGMExlfFE/c1XqzYTNZoVoj8E8
MPAmSSx/BPLKSMZ9WlHKUGvantIDeZ/K8uV/FURS1qMBHORKEjlR5dvu8uPWxyfK
bV8OSxeP0+3vTc9jcp+OIFJq2iMxA7nnCIKSle0nkMr8IxR2NtSu9sAekqmB38h6
HWqm8QYHw4b21vzXoKU3tHTDFW5fQUOCt/71OhVGTDDc8VPeAX46IHiknQ2bYjq4
xHONl4mj6hQ+3FZRDj547hp9ugoJlRvmxTUJ+WrfS68Cgo7G36sgNSo0GKtcESjd
+lro3VoKThuVUEvUGDjb1+xtRK3CTQh3fUUFS95vQq9xmkE9FuSD7MW8NCKjGlhM
Y7LxtL2iVVN+eHT2eWJjiPK78mQF0wo/fWyd8+cV6voTf2GXI/s7ZMb0NwT0GvJq
NqHivo6heJYEwf7E7BdyRvwwTstHzuMKSDM+S41+lIraL6GNIKkb+eSds9ectfnd
LPIMKHjT4sI0WQhK0etkxznDnHd4qf0grOrIH/IwaumNdPeGrbZmqsktVxgRxTYQ
u9QtV0vkA0X/3uXGaqwLy16ZBFN2N/DoQYCaiX+xjIxZGnStynjXQGM42ULh3gGz
1HUhJjgTYjekJevn1BfVxmg90+kdzIrJLFnLy/RKCQwgidjQgnzMGZ7k14VxbUPw
Wm7+PUoT2BfWwZ3aIrEv433/Q92aAVzXPBcNDz4diNYC9ubsAdXcb4pz353AYgTj
OUdMK4ZTXDeM1OrjyYC+/41sBblnFvj+KDyXI+rpWwhYGmW57YhKPOV0ZfQ1PMm3
3SjlmciKGN/+OqgDz0CNVi8fi4qdCu7uCWDfP7lHl+V20+7PutMBJ1BzmxpACGst
zCLgJ/HptmU88CQTFcWP6zCJUwV7VX/FVcTU4hMQe13mzbfIE/sx2Z92W0BPb68I
bpkyBQauHDU16UAJB7ZtvobIu8Z7RPlzJlHHVTNy8Fph+xHS6KS+tg7KXyi2W341
85xv1J9TvzzGk+LbUutKsQQjDOYavxksV2oy0BYV56TbxEyEsbWN96DUVgBpNtPs
8Lk6LiKN4Ok77OAhBqSJalHOXhQRwSe7n4ouRg+j+bZ4q3QLvHhVUD/Co8Yq2/OS
C3V9mfm6/bsDrdaV4TwUuuBJYs4n2TDYH65AeRqUiAghGrQmYrPygfKwir/sgqyd
1EZCyOZ9fL/rUHKrMWVcIbDGJxL6jMHM706dhAAWlePZEapqq/1PeHTpWlxKilF5
WRW1cQByrJ8yhHzeQ8t68svUDuz1qfCTPILL1iDEChCCGQ8T+eZM6inxbIbho1EX
89iCC1wovWy9kPdLWrUkNvFb5Yf34QLFBKU09iIRTMyDV/dt2J0X8IZ5hL4essMj
Iug2SLFNat7j1sBBxb4eXLgjXpa9+rOvafotxGiCbmnsHClxi19Ck6hy3S/WRJ+E
5MMJN3RGzqUb3Xr3y1ILblLV7QsNa7QoWZaQv9nEHfCZAB453pqJ9ConM/+PaUxD
D5j4mWVVEKWA2ZHgt9oapWtJMjSOS2tYw+O2kdsUhwBBe9ec9Uku2j9Py0SX5ogA
vdRR6td1dDmOJFtYU9mEYdUMSn8HdlXC+IpxelpZDnUj+3eUrYO3G+fkIexzs01J
H+bW58VY6qWBdpkli3hH1lCXZgO4Y6RIDwWfyCQJFgbCDQISBci0UiJ3yJ//h0Wb
fEtiThP1JFPVW9rIBojUd3nNpqNxKngC3pT51uFSMesGUyVTshab2geGtgk12D12
qQoVAzoHJ+x8DUadZha1uyf7FzwMPN55H2ZRVb24a/vimipOvn9zApW27bgtzXwJ
6JZxuJu3X4r5PUIr11kT5spL7eL+zuZhrio+zOfNeu84ILk8cHQC6kM4C9IADF7N
8HNXHfThyvWbWoi5C/AdsM59WNfN7QzwuyPWxQXiP43DhLh0x5+LqxPhI/wnThpg
IXZZOBt94xAt5HuxDTHQxfxJHuASZ1YspeFWjOUiMxPB+OyGaDZUimUufMIpJ9ko
rxx3sEyahQM54ES0shPQQagwxDtYd9uCf2XYak4dQLkD1bd6vI2GohX2FaeYTL9O
MoTlzYC9grAS/UGh6y8mWJ4XwOtte4BLLLQU9BSKBrdy5aaC0/FjXygiN/ngkFC9
TN6F3wJsvu92MkXD/9SfUDizsrjAuRb7DF4ahVVB3RCaqTmYqau45WOszHJ9vrGP
A/QMkBPOaP9f+wkfQ84AX9R4mUF+d6KkAWLJpdNYgecockjdi1QG/UiNA7QDITyN
pZsYf2RmtYht3uCa/YZx1X+YZYsRUdw9c/PdJu+LBPsIhGn0D6sMyv6uLIvZiwIT
zl8SOCkmJMIcxbaq6tMyZ/anVpM+t4bgSvGbDXCJIewoc3DH6LdafX/st9k2q6jy
F5Gpwn3QGa8fJ5s8uMc7kKgpHXbDvGqscs79Ccnsoq11iinAEvnerNwe6I0wh3VJ
YBA3DIJ1D2/2tzb5LLyJmU8BWfjqH24XDQcwNVM6N7LsT35j5+h6xqUJoAZGafFn
uC/PAjFx0LzW18ccWBusPHAJboxfIhy/peiE1iMgHn4rFwiOekqbHMKqYobpydrS
zQ2ADvJMIUch7SBZmmxevDgIpzyhReRODmOBCM4yKOXSLUbAAhXeT2qdUzsj99dI
MUElBeeCH1/QYMu4hLQTHqB+LNVbnpZQPa+QU6elTbsckyrU2ZSnCy10sj1RIZdo
Gboyu/eMyjDT1dvO5mPHK9pWEIxAyBam6WfRbb/ZjeqpoKZK3f8js+VhJ+WaPX2B
V13wrZGXEtuSJUAcFSOpBxIkgfRH72xc1VTI4Jfv1zl0uA8q1L4Vgl41rW+rtOT6
G7BsjLW1J8Q5cl2vaUo1eM1lViGuGaxD4hl6vNjVYUutsqQtXP48WnvqMDh8+9BE
hLBYh2Bsnw8TaDRM1nAh1Sr04bLhvx2qhR8/w46ftCW53cpyIJA/M/eDb6MUwNlT
OpoQHhc6oyIx8kOUaoHPe4flzS7dxOX3bjQ+kwW8CTcN4C2vwfoe3b+I2n2wuIet
83VCm2b14Eyz4LgvGMZweaXgejizX1qgdHMgOLwnEzGJYZkS1s4kQPnI2P4Qtf1B
hAVs2afRzEy7V+V/ls3CzcSpImiatcRFNlEQCIa95iY+84mC+g9wcQdlY8rjqYLu
MML+6BWmMVDmf1ts0DTa6IkQhiPjXK+XY7meTC/r/epg5Y/CiQBRZaKoACqN7PUt
3BZNmNobaIYVM61Rmmq+kBysQoC4+4eaZavMJ6PzlZvUQFqNPyU0VBQRXsbhKOjW
ysP6DYZNor21vbuHsq4SqMzIbBsTy2C/MIlsojYAcpGXy/bykC8+SCSiwz/RIXlq
As8iAsYOZ19wyobXcx+buUB1h86KWIoSmwYHoDtlZBPQ05fLa9w2wFhWe5IOFi0L
lfHNEzaXUKqdhbx2rvbQrt46PZ7ZGzLPFVRbgqwEsDyPJTYFBa2tVNtpLAqWKOUR
fxvdkJ4kFP0omYf1jwkAsALPCSzRzF7RrYbTj55CeWOU5W5EJw/4X+Mh1K0k2oTR
VUi381BfUjDqhVMcjr89WQULfimfo1pwcuTKiCIWc4K+OfbjW/Z5idjedm8g9neU
V8cnYt6tPVJOdctnBETBBhXyxkLgoS1kVLvhEUQrqt3lh/S4trbxjmSW/kGXSpPQ
/M6ASUz2lkMfZ0sL8gmiTyypD1jw4r9yn5U+39SsITYVZmEjzjADhiI/3Fx9g5y/
qP67oT1/CrCZGuk4Pmh1u/k8S23n2Vi6xPHacylXeG8YLL3FLC6S5bZBPX6byZ86
SfB0QPoCZn0vmx1bYE/1qndrUYGfl24jMQahsK3B/M4g27oaEMrg0Ldk4WKEW2Nk
nnTgxQhyHTCStOWb+awtxJ8gb2QlUE0nZ7FftyCial166thwhgBTclEJ1ZFYgE+z
507IbCJBID50u1hdQoIQj8luNFT6srnGOc+8GJBVO3oOspLcvAQ1812yTH1V+ZBj
cqhmQ+e5Ogp53TLZ3VCT81Nbxsoeg6GXdaOMQ2XCqQo/Brsq5RRzun5vMa3z4yQ/
1hLgP9mTgfbLIuLBfado56Fx1thoE/k7UA+JnKkPR+COKfl/HfhO05GXfS0sPNbZ
+rcSGtnjZDOZ65Abz5qJeompFhN/MbfrmdjfXuZZadsziTY/E2ocWaJ34rwxJ1jY
vsZu8+3v0U1rmeC02QCw7bcpb7EPx3xeRli+6Mjfh1zBlXvKRuafcoErm0vL6ze6
Zw5zeRo6FvTlqOrgEzxTGY7/2ICniL4Il9slgFIjaYT3HQhjSb71WQlncNDAl80f
INfiuN4gMFW8WbbvpMU+FXZd7YUXGd5fN1IpNdLVedYHEBBp5TLbqeiSGXu9cjPG
gOuXHPeeP8wbswGdISu0L3xkdqqYjFfE9MrdFRnyQVwW3eM6G/MRqozeeFg1k+yv
BLUBbpqy/d0oTsrSdLjz3FMVVS6S4D1+tyzxK6WV+la3GsGVBXf3691gSOXZ8/t3
xRVf6w2z3if4sqikkIiOFNmETcjq+wdtYcPngIaQdBrUNhtmFMCCpaIpdP5UwzXE
6ipVaU4dvWHM27b34+HCP79pIisBfawt1sPTReHbjci3YIkjTKSS+fTXggRaLGBz
Yc1QiFr2QeZShMmma5SFC/wYGnS18+yHvViRxZ7Tv6Sitpcw3WReMq1PLbT52s8N
5pNUkbQ882rB2TxEVRp2kwVlBpaP/wIbdvseFcsnijZ2oXA4flUMHk5TMtKb9lVJ
ZAyZk7hxGTRinbUkkic/i5tNmqcfwzUJW5WAWJYAlk1rPkWFGNp8mqA1IbHg49l9
4Ka6nc9dl7Kulp485B7KZjl36MiXFgtpU0B9Ux4k6yBTEcnzn+nLq70q8a9L/cOT
dV6peDC5OXuwKg7LKJs76KY6xUiK4xdNC2C5PLIuPBhwpmgZ2yiGOz1CgBpVs6jP
CCb42Z2fBeoOBtxCUgloAi24wu6G6Io6csyxUeS4n34KEy+/Ly5oXi/ScPzqQ/KN
ygqvhJWzJJGYQDZJOEj4C7tsOMAbD9xV0dmZLZA8+qO8eXm7z4XEA+Tdxnk8+IIY
WmrK2KazAkRJY12KKeKyVM5Pnd5SGVBlkwAuTgjSmwLaWS65I7yar0rmAwdSC27v
IEYU+3Y1ecw5NwGoDp/h7Ba+fINOQdwaKusZSaS1PEzwxXZyfYni4KbioBHKqflU
JD/lXGHV/5tCMbCbMhgh8IY8WNJeOSYOpS/EEaAQl+Tk0DZLQ5PtMtQIkee60AtL
OSwWwJsOU25HPHsDf1DKn0A9UMmj3wXJ5EB5k6mELOBpeT26ktCcxv7jRalcH4rh
Sg+t0CB4mGi+GUgG3+3SMyh6wsioA38QxjKTV2Scbt6qCEBS42Ejf+lWuRwtIYcr
7JC+nPajS1ft2NezP2PNYWnYdxRz5QhhcmJ6Mp8iB8gAG+cRZZFaMvGxYXbm8F7/
Ezh81ctfC2VLgTyNv7bub9tgg1M6D9BIMuTdY0GVCsXlG4T2+++XvctKDJwe/UOD
6gHY1Sj3q1Xcnxbrb4ppB2Xmwo4bdjPjzDWk6ZvLXIRn124hD7DF4n6SnJ7kHanc
7nmgK/lmpSp+/uCOixmQOFmoXOVyWTXNxf5XLWUgLSXJ7BZXyu59aRzI6i9JQNNG
20sPSyiVV4R/73/r4icERmm7rGUpivh/AK+98bOUn3fQpqtrBm+Bl4UffiRelpPr
B3szZqJqy1isyqK6kvx6CkDC4Derk7fy1adQbfaGgCZoZox983vj9Y2hLL0D4fm8
YqlG5eAbqFk+g4A1VuTfw+iUtfYHOyEPiYnrCtLhfBzYmg49Bu1+zrbFLqEKvK8i
g2qFzMkBNLNtajZsMhpCpUOHd9cA0NaspWukLWURft62Dcg+XPiKr2PGwA5aeEIB
UqTv6OJM8lbpKpOzOQSShius8ZvGPHv8zoYuMbPELyU3g38+ufz+cxoTZMM98dMJ
laGibpujMZjfOHa30RFzJbNc4YUVc03XDszCVVT5vdK0QOxLwsDPjLlHitzOXfCk
OaIphRQaAeK4yhbmgkYVV/HiHtHR+lclrPcbwHuhOpd8WVkHVHI+KI+DjZZ0vpDg
Lz3AsNpy0++Uuqxo1hKxGu9MI8zMZk6VqN6i64FvqakNRaNTi5Y6xri8gxgLodIH
1c/UwlNGYGnuOK2sAx7nicL+I8erha9hY12bhBMJrCYfmSxEEMAg4QhT1U7IUMp+
1jyS1KrX/M7h8/qB2aqV3Z09alhUCzdOcMM34X6wjEHOtjzMwrrN2TUHOkuIFPNP
X1kfMFfJmBFEp2pFy5Zc8b2BVxU5itWqc1FKvhgZexfwjzMzc3h8Lpwo6VoFPslF
7jluTnbwvffc3BZfGkW/XPY4BCcJ+oSiz9iy6rjbxQcrHk5Xr0GWC9k3vS+vhf+M
ib0LuF827SHxXLOkVDaqHtYioRuotkIOgdSWHfbLc/AZFVsswZPMvjpFZJBKgYhi
IB3XdWtt/cVd1lq/ghEfGYB9YQhaFRXKWPPBpfIRVP1958emb1fb2iIxPtkpDQMp
BSivOYIIyg8qxCE/zc0iHJZn9gUR70pwQ3PpGHEn5kwuVG/wjCF/9KOVxhHMX35x
zz60hML1DO1yqyNyuglgXVb7NJeKHIdf1dYEHoltc4IX8YjomZABCXvWQeAnep+H
36Cl2Fr47GnfibJqAWzZCZ4FguFLoRKb6u713gHfCfv/FEBCHkEpg94oI3Jdousn
AgMS39AMRvecrc19Qsak+12T0Ytrf4DQgm3b9sjc1EnJgVQ4qWZZQLc/tfIZmgc/
XzcbboGPGaTOIBZrSAj8j1LFR39r6W3FCP7334WkzcEi/AkC8BHwZ/pf4cSBLksP
pdGL54P6EkzVAH6QYebZjkSWifOqrtPhGcOPdnio8QrecLv0gqkfHhE0Weq48icC
mUCUDKJDAEEajI38ItqWzRml7v8cy5RYax84017c/4ayaWXoaGJi15GH7w5HqnNQ
DmZKe31yUoY4HQVwABfyhDciYQx13/Q9dN5EgzurLTvqho2Ho+VvewX1tQZvEFrg
iIZui5zztOgXAic/BOtafHzWuhEU6JpF/kTzC1WVSu+A+tqVJLMUzIKj76ezjQs1
48IKItHEUKY7idUV06YWU9J/l9tAqzwzYK1xzoYZxCirMmhoNQHq4XYSREnjHq6n
EIUC77LIE3Kan/4KuBeF12h3Qp7vkYigkJWz14K4QLYRbBxFdFdQY+6+S9sWKsYQ
R58e+8HjuymJFR2v0UbLKCgwjTzP9qDKI7cJZmPmlPNd0pMZtZRCOJvNF0tPxY5m
4IYRm4enN3BgEvy0xHvtNv3on4ya8EWVgsbt4D8hd8F87b9N5SvSt0/RMBCqoQhY
qJOj3tU3CSobNHRqPqHGe+aY793kWC7nRMDBr/HoKWjAkHa0mzhi5LNWrW8rhig/
i/kHomsnLV0GjNbMZadC7TadDzdxE3/5leobeOqWOQtuJOlgDb1/jqrolRAR1eFs
qJ3nB9/s7cMpvQj7JMEBB3Ik3ENQqk0nb9sd6MjA+G/ScZHcInVOb8IRjIODNS2X
f/SKgnXXDKIN5Q+4GL/F2hvipc4OmKyEYPSbP6H9bdc9hmbyDCqh6gx8/tMmvTPx
W3r1RBI0LnxHVXdqKvdCCc2qt4MW4OnxPq+70vKF0vRrxZQgtB4BQn8+oCzG1/e8
8Yy++ZCsvjQ5ejBlo3BCqsWK7ZygFPccivLLDtlVTPZgkk921fJSu+aCUEErTi4A
Dbwu0L/AHR8PHYb5nPUMS5TPgRYDu/4bq+FPmBIPQ81zHUNRj5pEl+nUONF9GtRI
j0W7EmwS33M3+drquj7e7BrqP2qFY1GuRSj96a6xYE7UYC34LFgQFF/00JPN5AmQ
nQ7U7FnT7vV0F360T79wI3iGBN8UMFcs33oS+CfOUcKztToe7PKdXIUhNeViQVbs
tM1APpBW1+QB1cHiVqyRUHBM4lytyBphZxZdSyEEttGHoIDAgibHvcXdI/1M5u1K
SKErxYK0+l2hN1t12dgzmLjMMuvq1WdUJyXCaqFC8l1FvXjRHz/pcaSapjT8W6PM
VTSiCgptFqSQvVKIOAmcaBry3p4nHD7zghlbay49zUL76zUFjugNqB6LB0tSmm8d
1BHahbd3awAwIyunwIfUsODPFxgdE/+sCwk9eaaw+29uiHvdpt7E3hrttYvI2W8Z
lwWOUvZtMu/4vMmaFk1cGe70nC3xUmB+Nrj6Ppwn332GTRiKgXOQumH26rhXJ+pA
J+stVt6XdtKdAoLPxX+TGVgvdKTWts4QoN37Anm1EtC8F4w0NJPA+FfuBOcuB86G
ny2qllI7BTHTLA8lNOHPqs+Q2tgjtpp1Tavng9tds9aJy2K9pvzgzBkgVfZ2u+sW
ALshnI+u3ZHjV6jEVHjYYn3u+e4XFl7uPXfcA3/BH6w4imy4y+KGWCH7A1ZIVPEw
Oa29lxgLUv5vbA9vYYQo+nZrFejMrqTZ5+mMOIigiYlkbD3ZO387PfKoxv6w0ClV
jNnGbQThftBq4sV/b8kTrSekohaAYgW2bMWYzi5ov5mmQ1HnGMLVy4PuY9tfeoMw
g5SiRpZSr9zYDHIFRZo5CwbxLnC9zqubT8Xyt+ZhUkqW7sFoRM2iVNo+fRGWejsH
wxLPvj5FkMZwZgCm3BJ7CJNMJScpNt7J3icd2RCMzZFcn7XTC6yRU+xdZfJXVT/K
kC4e5xwa/rMFjuow/u33ZeO8VR+S4LVhkxvL1Akpik+Uy0GYQNCUmgzU9tKL6CnO
PPWqUPwhaw9I8nnKONgc37H6zeYD658b/S3xlyN4Q6f5Nyb+G2KcC4D51j8umO6O
orh5FMlqVT1GOTuDatJ+RACpcHxJahOlxEeEMcpPU0LzZnHkgEumrprYJF5GT2pQ
aRKLHINd0NlfV++UcoI3zNCxnJbuicJdWOzZUrWjsiItd2zsjPzpz8NGBeOLYylA
LJiPcet/rrODZ88zTJOdE+BZRs3eXD6E1mkngj95sKynDavpKshiV/9auRJRdBjF
x0+5dwjotP1ievizAZMc3+nHkxpdHOVS6noFalDAU+jtis+xEro1UT2ddFGdtLGA
un8jsgN/BlQ+faPunDfDam43XUvIhiwpXAYW6ChHZNPvVo2nVEklTYWUrsUMvPw2
HDj3DOPcqa81wEh2XS4iKCudTQYCp6n+JzF08iKFHcTyNONd4FJrKynchejjkUh0
a4TNL6jVdnSyOvU29LibSzo/85btT6QyLSjmkwhzL/YWMGaJibMLDt07hYCGtbIj
cWRBih4Qzp0DZ3dH2kfbN1jZtv/Ubyzz5f6li0YHzrxp8GTETuuf0gfMp4wehL2A
wnCG69n3BqjxuqIJzxAiZwfuH434pjptdIf3h+uWLEY/XqO/vtaOG7KjAZLSyaow
0HVklFq0dwXABbB54K5HV/NS9x9MMLamdQ/IjxhFtH/lrKZe9GCO0DC7FeLqca5Y
SU8hM32VK0SPL1OJQ5sUny35JMncw8SKz0i+MS2KwrkRc7dLap+cxdJDn7hYbIRG
HH+k7XsE/QQVrm1HFBBcEICMFRQCzbJI51Ng3NUBEeLLWijqVBsn7K4sSYgiWy/k
x4DdOozl6jbTizVaz2HLru0QDhbn5iFfgQZ1vr+aFMgFyXPvLCyCs+8PBD/WBgA0
u5/0+M+W8XYFSbhJvB52BOzAJPhAlw37kVtgLPHwWZXHFhjeSckPFlGo4iL8WRHC
7NJXfaXQzbiEx00XU16tbwSzx/X3KBfoaETtksIwez60Ie4RKphpXrXZWa4nfY6n
0BpUujyI0aieM2mjP4EqOVeJNJpp9VsMEcXwLzmWxKFFrEU7eASt1fs3zUjIXEUm
K/WCKpYp6fJlkXiXbBL4K7kwr2YDa9da/Ve6kg/6R+x2VDwVRN2D4tuUa6wVx8aD
QBMoKAmdZMkSa1cHnX3ktcQzlHl8/ORKfUYPHpayIz6MqIbJBWfaeww5aQ/qqTZD
4pOW1sU+y1lYkk+AV5Aqr02h33BeEcIiuH37DaVteurGPOmtaZUiW6HzvSgVJ8id
O2dP17jn2dBAf3yY986jNeO3SSqAj5ehK4Td3grIYG8mXyAT2D5uwmS9j5eR6Xq8
a74lUXrRWCKX9N59aXv83i6f0Lv+/3E0C1SaXszftRASs+dI2LmoA3Ege3OBlHGB
2gobIBhndXeKcmTOQXRy2pgFBanZhdc+LGa/sARyjvUzyrq0Ah2PQW/uBUuRBOQO
w/77wDPT4N3QqYIRw/n5alpFrRoxFP1A9LaDFPFq7qc2bKYWbEYIRZZai7TMnwHp
7gE495SyUtursH9bBQG9pWFvMgd4aAnNL4FPyALWtf7uhA2geliv0IPAB2WlJyWL
Ah4yLtLmAme6oj+qhqSyrVugAj71Hfhf+m+Gt53JetXaRQ2irKJN2KigSM/FRf0v
/M49jge5kg9T/EMAdO0PHBxjYv4e0Wfau17FXwiQXvMuThuqzVBl5ThC+4s56UU8
sWS6/3K3pQCyNJR66NgJWP+gfiESvAIBe8p3oUVfv7/625oQTFz+JzcbeBX+ZHke
tQ+dVl9w41T5m5IX72O1S/sNanDDj11gzhdYbJOVF0B8y3o8qfeYj16be5T2ZAYC
udH1wQWiUWMsn6QSPbuUoxUSXSHl3AFbuOaHms4IcWPgk4odScjrdOXckZg3Gz69
O+ZLzVOC/15/CAWz2Ljq/56yaMQz9xjCvH1jrDTYJj0NEcT6UCgnr0xNjQv4ojuQ
AEM+FYNhXijdQ0z9Sgl3+w4fcHHRfOLIxTSZHl5y/itFGkbM7o+tXOihhPp4U/Ig
RgsWdLfdJaEwVF/DQug70Hzd6zo1GMNn5ZnXyKyTiowN9gZvbguBbifn0pc3am2d
tJH2M/62m9TJmfBvWzcR3Rzb1dkwTknVUgvirf/wAImelNpMGPbplB1GGX25SCcV
Y28enmzBP0dEWcGqjhz2F4TOlvZx3S4MSe48bnyVbmoe2DDNPP/TNgetHxmd88j7
jXHfFjS8egoPwXfSTSx0c/xUWK//OhdjaxmefIW1f7bs8y2UDgf6Y2qW8sNiYh9S
CZI+SrwplsClJCXpmeU1usKBWY5aREHU44ZsgosWqIHO4eINLFQkCakgUGHiKxKH
Rwv4hQc4aU57FUceij0CmcRBKhr9amAwPk+HmkgyV6KQc0exsnnkUsg3uevR0Lsc
luLBRF7PKsYr+l7FD7slw/ojbBETsyxvlKE6X+5XyeFjGtJG7Lvt4ZbQr76jUTGw
R5diWNcJHudp5Lv2jsTKKhnHj9P8lVmAFIw5DC3Er5vayUnb5ozFG+zzVxXFAVqK
3FToq79VmBY3fJ56v8A+b5HD2YZ2HhCQJAnOG2Us9zloZQlr7GN7Qu7RUnHHHQqh
7clbjN7oJxZq1fg6vPq9z40Nlxq+L0FDOVI6r3B/BXrKvWYBq7cMb2t/0SkGwmO0
lmlmF9KP79zw49ZUuchHiblLvoLCNpcEJjLOwvuAlzFPxWRPRunoXLcYcSyP//KO
pSIITnDpDwaiy7f3U4SKCcrCW01ngpE5FzTVIZAT2q4CeHT/UGgrOGKuEqzr1TPE
OcFdr2jdI0VjpxjY4FEXeQlDFZESsz+Y+PFRQ8HUH88w0ShtCCg1t+SWSOiThGjn
OaTb/CC0+mNJyqFTi1cI7Fq7Xirojv+etNYkKVtjB6XX3rEh6/xzAgLF9acQokAn
sEhrgWTzBdLSUyfBRJCH+VWx04eIi4tA2uRxxsx9mqKmczNSy7RUkrf32GcWtPBl
ft3u0eHvY6lOJl5xCFa/JeK0QnzoPXLMmYeb/zGExDaSCWTHqTbQ4tI9Ss/MfKWs
B5pMRHFy/LrpAaP8IVB4838B0SYx75JeSjXiBufn75xzZskK5ugxf+4rrGuQfsFA
8NON/3ssG705Pcwt+VxEIBSH1O9FwFo+o8fVbKSnz+Ol/MbBOtafLGDUr9DADJUn
4P2PhowGxE7rTIQYNpDY6qVZJLdT9QuF5IECQQidh7V+64peOBAP9ttnE3Honyrc
y086vwqHFrfNdbmJxu03uOaFFdpPE3tv5BukAkEbMXM5LoIFjxgFPX/hJJnXQ0r0
FCBK2S6ikLeyENzZG8ijPVWNKv6ZB92IArtaaYI/ToPBtCcxkgnSaeQPgBKy/+sm
Dqwz6SC/OTNaEWG6Uj6w4YVMnEk+j+vZtb6Hza7xWqRKJyor65uiBNas84ncTTsi
6MW9qt52+CCQRPjBbOKXS8QuZ/9bPasVGRf/+sw2HlfGb/h9LW73DH8qO9VetAK8
EeMnemeM3MaP+k8wzsZ0D8Oznt6qOO+H0tsWXp9IF21JcMeRMgZfFEylUsQkwxQy
vQ/2ga7Qf7SQyvtQG8QGDfJQW628+d0VDzDaxXxGWcu6yOcW12yaWbyUCflC+sHA
tRC+6LSU3kfIkPuJLrVlFYsHMRvaTpmo/4mRWKGUsNqqx3r73sZlmPGwYH4d4UQb
5BKq/hO9qQMmy6tEtiUGZpCvw8QGKFKGQAW6eYR1afFYItVvMVCJdX1zq9KHFYZj
5IFzL4fTqj4cPK1rQSVvZOK4TZgGz1wo1gGzGdMTfpMYWR4SpbdWjy5GiLsUYPxX
EGubI6F8llOpdDm8plvCVxA76pT68+/tj3v1ELaW3kbIs2rNg0UsrsUct0HSnN9W
xSZc3I5d07jqM4uUf3hlNTlKhMTVn20GomHS9G8A+rZpinJAwsPpAee4R/hOZ6gZ
gfreTPErR9jdb2SGNI+nn/P4/vwATTCysbods3tsIaDsba2MaoGX9Kswv2RLDwZ3
DZYkysSrbVDjH0jPyLUmiDTDeULpKRGbJYezDpQxpAz40dWNEsd4FZ1YfqPAGTmj
o6BetS6w8L+r1PSQ6lZX1y5/b7NWpNVtEqCkQeapgO/zp6NRrBfEYfVPEGMYnAUF
zDg9pr54yjQuClMt8o2/CG+osQqNfar5/QAXxE4xoliVkKvYdrYN0Q7fVipqkjWi
gGOJOpizcDqyHazQIZPmuVvlKpktlCDzNLIt6gxe94mDWpLMJ2So5EqM3eVuUAsZ
DMUgegDwKIy8cMBpOIMRmiwAXFue1zmARSCp7J82AdSj6aTTjuQjfDxSg7TVtoeE
0r/wwvkkYfZ8z252M4Lmy/h2OfGFTAxxpPV/5jHkui304Va/Y66Qb0mFpAH+6HYb
jcnxM0jsUyHsxlFtYubF1Bnq1CNOFzC+W1aFvso7z27Z7dJpKD6u08Usys5sagBl
tCp8m+LyBLy4TP+GpTZoLGhs5icBSuh+iNTu262YzO6JlyWsIEwNDoJTXYFb+alb
UFm+kFcvemvLwoPPOYrUbH/AGKVzLIP6h/5TZB7Xwx4OEZ74RtYKaDddVqk99MYr
DZlpidW+FGEGCeByFUxzgQ18lnvPai2Nf/B4LLdFPafWaVxCoPDpzVRy2+lSUGmY
JehzT0GusQB1RVRWKKAuBsnYg/ynTpymZ5/m0jTFiWbPuhwxKLM3Gvu3nkdPOPzU
Whh/5gfHnwiUsIRNOYezMK7ghfEh/HKE8jGS6qIYaHjLvKuNCiMNQYacBEwkPqoK
bueyKCCaLHIupH5iZC8ABIgGEQCHrIqzT2s3d7nJlbSwUEvParDtC3vjt5Cr3O44
nBVO5c0JKCqXJHBdKlEjG/OOC4PNJ8DV/RIkVY0vJccHKtML6h4pWgC+rIKHACS9
fDR2Dpbz/NQoSoWXpctyRrya0UO0An/J2bZ1Qduo9hwWia801cEMGROtxLC23HR4
qwiu0GiAus4OCC25Uq6l1tAZClSPRASnjz8W5+o/tOUlZJsKFJ0l2qLHKRhExCAP
fBbJCaNOIalYcl70/FqxddGP/n5AjKd9EVwlwnUtNHvhmMaurthQptsN1kpBkHrY
0IQm9zbykkf995N/mYvHhjWyP8COAlN85fqC7dJ2AC8oIL65Twis9kVvCtHO5iL1
M08B5FY3U2cY+2QX8wr92TbVzgU4oW/uhUTEqSfyw3X3eI5cz/5jPnit+xfFM0dD
rc9UIgGEuGLrRAFk0e8ji5Dax/xIyLi1NDwV/3sr8mwtI1uiVIFCN9ww1pfKzAhU
GFCPAw8FYMC0GybU3X/sO2a1hMQ50apSdi4PfsgOq5NHlzNd9dAufDOzcG2V9xVi
xwVupHCHsJv6yihfqM/eqKj+VaDn+hgddmLIzX2TJIIytVswCHMCDCTw7UyTP/nt
DYUnk+F4iYLdHUhXffSzOFF2IHNJbADqxmsZFP0JDMFH0GdV9AScbR2KOE3bHRUC
S/Y/poIBYehYu5JqvYWQ4ZrqUFZva0rudC7Y5/CN+AE1UNDisHfyt5GLu7jd3JQ6
sVE0PkvcagbIl0Ij6WzsN608l55vvNrW4BKfxlgj7J6y7BqUG1nb9+0xXEeTGkux
a/htJ4SL5fyatkNRlJWBFaKn2exWNxAvuj8BkqTeLW1Ne1SWScpYxLuhR02TwIot
fBiSsA5pzuKA29cdKvThhL6yQflu/+fB8Ud/voSpElTFw72QCxJ6W5TleC8qxZLa
C2zvYNMfi5ptiLDvsC6w8YpzjKZZ7LaK6M3ttMBBjX/dmr2ZT8nPDC/BvG0PYyA4
xepUhlcBRmykEvVOOPtZMdF61WjpafNNZbJRSG69N7gM3iK2ymm76zurLussnhqR
0BvqKtd+kbwuDe7q2s1nYUnGnayGrnLw4qJGibhLYouHZDQ+SclWywWiGP0xiV4f
C2/SESclTMuejXmMZeEqRtL4bnP6he07yhDSVHXLEJF/Ace5eKSGX7SMNtFHUDal
E+VFrPooajN5knkf464IGOlYx2kA/rvKxLcdDRf5UQWszxRmfT2F4Sn76jpQjzeK
wLZpTHMmg1ZpHjUSLb7lSzBc/+IPsC+TjlOXzRNvgpKYa7aVkFP4un7XjQXtNu55
iNLlgPyXbz1la2tfVTd4zNmETEjQDbzF+7omtfB59iUCMdKzbhQsxZ0ys0mlsBTe
dS2Do991nkLQkxgj5Fkz0iOgwkrMG7UWAuNSmBfkzwWvf95/Op9Wlu2gCxlSQTZ1
1CidaZggvMEmzuHxkAvL2Qi0HroZO/tlezfopwy9WqYoNJE+SAMi0LUf6DKjfJ5l
CFqrs+IjWmGAGcoiYoN0C08mXO3ZtlWpwTu6KFTZVydXCuHhGmv7+2dy74Q7QhOg
AYqdI9++hsy3VGAkYszu565FO8045rg2paRBsQqU2EHMMke/RQyY1AxaQSt8FSbz
7HItf/9UuEJwMrCMh7Vdx3zSvCvfgfpDc8L9pDkr2qKpAjCYeTuwweYMQMNmZhSD
rAPD68Kj9r2DeiG85GKsL/1BZ5AzYndEyMJ1UwvAZ4Js9xiT2o5YB3ydqvIEAE2t
yxbIU52yhF4NUmnimZqQT3kgtAkgMYKtCk/cIUGm8sb7BKeRXve3EsfcPSc7OD42
SeSL/bhWYmqbdzAFERLO/cx7sw1dAyweLf/2SuAca3IHEtMmKgPbDiB+PkdYkSNZ
byv8buDOV9LD/E29aZdPqW1OSVV7LtEgtdkYUpi4puT2rR6ruzeO+EmR+VqXM8Mx
U4pRq7h3//0rMYZW5HBzn0ttAJ1wQz4U6JPVcBKP/wsQQvqA7NUiEpi1IfBVuhRi
aBF01kFZK7cAVrxJhgGHQnn67fLOt7RopEl44BSzbDVYqDILAVzKrCiGOgw64jiE
mKVS4mJhYw3eTpIXCgHg51nPWb2pT0DP6ketmUeI/LWvdLoTqHDwiCn7vSEJDBUo
n8+EWi1V1zC2/pfRq5LO9S3NcJTfFq9ufUtAJiwjFNIFST9lm/s5FWFIwes76RuV
bLoMbiVB5Ll23LqLZq6+Sn0t/ZD/DHSG4ZzqD5FxkVC1dZ9y1rLIki72ZR3EAdZO
aiiD2lmhh17W9zyvXZ9lEhR2jvjjXvlNNHzRxxDpzq9uqorqToZJERZKvYHPp5Ti
MBOPYsFPjUcY9XtD3ueKR331W3Va35fAGbuCV28InEHHwmal+8UoR2x/Y2241iIP
uC0/Fu7K/6BHVgcgCZV1zMGtwfxb/H44mZmlevx7KbMhOSKEIm770/RQChq0U5Sp
7EWqrJz92DB0k80B2xdDlgpGIueOZ3h03eIMj7MHnE8Z96EL1mXgZdX5ert2bI7F
g6XxJ3xOVn2TlscBzfv/B+ljAU3wtTOBFQgqZz8MOcqwpooPkL9fFCUP2IUweLJt
wKfIaOXCJ1B15Q6UeHFhW5IsdFYLKMn4MQp3fw53RYGdfP1L10aAuiLkJNZUSwmu
YCseJq8FCOsj8DiIrzFjGghYXBjgGWz+7L8rHkXm/gA1dIaiHs60Xy8j2Qub1EJk
/SATkmvCRwtESyXG7C0uWv6XvI78Qz7XtGGjAAQTnLxjZ2FOj+JYV4G5QWqrnzxk
CA6REw0mTv6IsdlaFGNZndvw/RRmgrXz20T6OiGA3LELcf/DWDSzs8nhMOmuMOZ8
dUzPYr9qyS3VUBqBHj8jTnZsv9iuMzjo+bLto3J0NUoTqNi3YgLVq7kw1007HXer
+dmtIzFJYlnUND2QzyN63+nk+OctdFSVcQCWCInTfqoKH9rRdNPuj6jxfLuSgVDm
AxNcCfukGrEyphT22yOdlJYnARaFcrTZ7D7aDXtK02IyqtY3cO4QRDiaGShSI9Ro
ccyMPqYkDDiT6VOp7T4S4T3NaI4dKrEGXIiQQ0uBApFQGYrAZ+ibjmL/jQzBIFND
c9ohSmWgka8t9R5N6/7cFndx/ErzfbU3Zo6UBNk69I8IPntA79KhjalIATEN6rlO
0v3xsqFEl2dAZSGF8aaN6Mb6Uv51RAJiSjl3rB/zOCgiAsH/2vWVwomqO7yhVbl+
CsJnHpMnFo/RS2Wd20j4+ZwIF4mHR83XuiwMtDIt6oPwMZt/aS3dJObRUgPDz7Hn
EwuAN15dTetpNeQMM2d7Nk2FM6PaDD0wNHkA4krzSU+3Gv9Bk3buKAFghPzf+8Y/
cO/PpZkYSvgi9pUN9oOjCmEJMyTcsQioLVuLPXD85BJRhMMG7bniUjU3kNle0Rsy
IqTzR/A8ChUavepfhmIDExLIxzYU0HZF9ITIkiqGqhJVf0G6P0zf6PzbGWozAlyr
N8EJfV2JV7u0IGNIJZaoGUeSF8pTXsqe671+x80OaS+wGRhyppgE8l/rmk1mv3j9
My9NXd43nn85aA9GQ76vWSJ/hyl/9p+uxF/nxFfF4y281JspwLtBd7dlC2vluy+0
uC1Bx5zz59j2/f2iV+VUkmIZq80iQ5Da0YgRjhlZD3gYjs3QQI1eWVsRnShv8cUh
XinzMEdyPPwD2//uqQfuBEd60GGUAoEMNEoRZcNgMeNKcTIiiMvIxs/ghevi+Nxk
HuyIsseuTJS++UnoFy48msG3cw/ecYHuyqYuHuTY8qUrN2XMvobrhIrOzvJ3u1NH
xrOMzP9th0311un8g3n/i2LWJb5I8j99tUzU+LsP3RcmD3vu2IYrmz3BjOhcxxX0
V+bf6cG2GV+eTjF677XZKqq3vDiAKuAvdGfaypPjRUTQM3GnWVok2+jQs1fpTPdG
ldBXwfKZKnR4WgXyLIsRw5cfWOVNvjHYLm3Pd7SE6pD5++ThuSejltt8pERSzdvm
BoV/ppCO6tHckbOp75h31HIywlUNDv9NZBWeOyb9gtRvcWE2IVpXq/slEeEWIpOO
HXUO55xdBePvV64eZ/iKddwjnc5D1dl41hyfxoEB7O1/0xoOeOY605UPMdLz9Vrx
wxQ+BbnD+QnRqazWOb38reiDc1PSA07sR/UPimvyh75b2ZIVmbfJvg40aD5INWU7
QUL/CGa+CvXmu+LMOL6EbRgfq3G/lsDevfeUWPonrMittOX6SRmP9R806y9o5NIz
fcWH3ObzX/UBbKn/fsXiBZmAVihIzIaDKvQ6+vhYyyeH+uNdgPy8cbrVAkPT8FKe
4m+G8EQ5xI3zbRXGR+FV2ZW1+d+aaxAh2tdnBvx5uQbhIUcRr9BZe5XMsth5cXtM
atxnareBP12MyPNpmxziufzUA/dtQjNl7PTw4wr/t0k3lvU0aazhYmfZlnwlhZEg
/NA/byFzBU6TWvvlmunWHsZkhRg0DTz6Eh0Ty5QbAJXucEfq+C/acODpEjhkkBxq
m/24+7mkGl9P/IHvX8rFna5Ks6qwHLahzxqFZ3CjkEYepJfscLihcKiJhX+aBhHj
gXFHZJOn/50qDxrCpMbIh7cn2JmOEdPLiLvvcz+sX8i/qypLngMC23sJwVv8J/8y
AiOEnjXQXPphyNQm2PLxL5G/4h9J8mKp1u3V4NQkzsSUYDlWTS0HVyMGe7uSIl2J
Om56aYBDvbtjv0F++hMWIDkmfuEdFq+HQCYlQKsjc8oqZ0bS7G69gxDfDkzTLtpq
GhjAQnLVHOKE7zEwr3DGZz52KY4knOKyJBqp3IuYVRxl7EgLUHvp6oP5stsVZKCv
CLbyrKnJegj07azdBYMrJpe8SxqlEU+lcCmV9yz7QvdeTyLlzQiReSX3v4cRCFjr
DX8xNZlYWDHl+7C+JKHwGlMtlqWlTGKUIZcrgCmVwTwtrBwKgoc/okellqoB4n7M
/iJVuxcrlAVONP3XiQDjx9YDOyDFgSMXu1AZSpwFOsWk70VNnIfF2drhdiVnBEhV
MbhKoHhXYOM5rb+ggJez1y43FWDSGiSjFfCWK6c1v0UpwRLOGrywNsf6r5Ye5SDJ
INyvs5G7VQLyLgoPox9TlHT+Kuq9fG7JS7WWKaFcw8ZXJmDRLpB11uH/3GNbT2gY
slguescMjd16cKE8W/H9mmJSNT8r0zreFa/4EnXAEt3+I+LezSgZO17PiSS2bRKz
C6aVJv0IATGKnrG3aGPtUmwQdNTRip8PLP3Bf9eJhVod0IGk9G5LVcpT/bwtf9DR
8zb6zmopI2RsrdZP1fwiBJBnch1sVx0cjxChlqUKel0h4Z7v2NHIdV3+NQjVHRMd
R4e9nHc2J9hitefbYmmUjaSKIb9cvpmcraJ+1HeYpCW6Ky9Pzqxt/VxwMX0/2fPj
eTqyHO+enHCgg6wg70KLycVwZV4iW8SzRSqL4aYs0GjtQv0B1X5mdXaTleHOzSnp
rUmrkzqMtYymbB1b/NcJqiE3xgHa5CR7vZR76NGFhRTA+XSA3UhdHd2eOzc7sGNS
cUDSO51N0L7F4pgSV3WEUH0BeMpXm54gbjuHsyrKvBCVYHRshMKPxmsWSzSg3DIz
MQcbMzDur2EDsK54Vqs9wBxhGfce5pHvrnWiaoMhYAxeD62HYq1x3XUOmajRW9Nc
MZX3L0QAU3QJjDuOp5Ty7LS5sIUjYe5n5up6vl5N4Vvk0dRaCDniHM0JtXM+/DTK
OcfaD0jxmPvjxRM1nAj+wYD4LiDOnDE6K/XuSoi+NoaTYA2WFWj0pq/2xJ2aKJvt
1fjiMbs8zhbOt8zKLnb/2sYbQoCp/dy/aBjOUYl4Fg+8wERiVhonAYeoVy+7SlW4
sV95TtfU72rGVv3uVNV8fnuVUgtQ9BxB+LeL713+GrG01BSzwYIGkh8NO/U5IUVo
ehEL7J5QSIkgjumvInl4NZmSbWFmFpW3fiYzSD/iWI36LEDQ4p4w8icxoL5L62fQ
3XqivSfBnxNldgO3jBZEcQ8avwGUdoyiKp4Yczm1YwGBhysZA/KJHcKk+CdvOz6z
Fxnz4itC0o359sFV91QZneQKbWs5N/IPMPRW300QJmBBVURwOOhEvIontovtbrB0
2wiSTH1gf0Lua891TFbHaeEXdICGkt40sTzZW9anfPUTOxBmW8+5iHtNwrYFId+O
kOKGSYx4oV0xnB0yx6N/VOEbyNKuyapxS1dH1ogOSDv1iLU8mxn2twxz9CEF+Az0
A/1H14dTe4bGrUm30h1LQ8hTt78hnpozukM5LO/GbgHYfkeYxlBP5T5ON1iQZMpu
dJcn4CqvsauOd4Qt3fCeyRNTWXhXfsXXC1OXWdnr1OJ4LcYI2BL4ZFdAYUiHGxHC
uHGBncMPY2m3s2vaK9DCVpPlxflYxOlQA09KtIvg/gMR5Y0+aDlofgc1u3Vy7+Wi
uyFaw0LkTeOkL58SeaJ6918opkpr/T+6XbETONo89E3XUBqnszHgTmDIKdLggqp2
Y2JOFlXhvJQF2dHbdSLmGbu/P3spjoi1plnMQIMKOjVxgBp1FVdtpnh6EjvkmX8+
AvG+bAoLoyD7Om6o1ZnMk3A3gRGkhrDR5tSDwXWL3iLwoqwGt6xQsAkNQg+Ac/u+
mtJ+uuxq1PDifJHBFqlJO21MMJXt/uS0ztw972Y5NPaOdmRw4Y10gusCqx87N9xI
sZPizQvJcGXL5bDXoWqJrQ6s+mJPl1x0q33FSbs8e6i702g43EjX6Db3oS6Z61Bx
Cw99JI04eW0IlJITFY7EY19o+9+Hf+hoOGBVRu8KuFkIUci8ewiXwn9oapjuAuJ6
BDJNb075jOBinQK+TlEHInzCrenFJCqdmHQKZjOgD0hAZm4wrEXOBri2UNGYOb8F
rPF+FlUKO4w5E1gcsfL1OMEyhewTd4YOFK8hmcxIYOvbYC3UgM4iR5KOQ1jf/nI6
lFS+tO6ONCZAuxbiubeotMhiAvVx9Emc45uafO1/bXXjTzB/jyEfNPFGEpn8zmi1
fNEq3AUacQWFu+4dUhHpmNWy4EZKrPVaUoAKoCwwwKds/KQCakSxwqG+KxWbhyey
Ty6rO4j1EnzPgqZ22AwfNC//CEh5ZMz3TEmnq6s+iVjz9EG1IFncxHM2WQz/rGd6
bGDDFr5EDe/mO7MeDa0MZWGyFOFeiS8LKq1WirCr/Lw26IUM930M8x4kOKFFgvw4
YNPiBptU0zjRLhr8xLRCzyZT/xFOITk7ksNJlJmFNal6lar5NzkNLYhP8y517/h0
fbU8Fidsg2BY+MTpAYO6k6/uiJMUL8o4ZUM+Do2BUWPUMsCfm6VhIP5YEHfz63dx
A/2jFDgj9Hq6W7ga5Xb0pSzUCZqEWuQQ4PgycWG3W7s0jWQNI4sVtM1au3xINBPv
AIJ3F5+rs7Bt00FHWPUwJ6/uM7yBsyE+ZmIIzrQdq8cCFE9KjF2a3eE9YiSxSLAk
i/z3OOmvDT1PqQQW4yWAHi5vGHQZs2YiIzYARNfGRiqSmd97HNLQBPOBTLGjfy2c
1uILHG0XLDEoTtDO0oN3TxD6pEwnc7+a25TOy/gNco8uZ+UnqXTodRRb8cxpAR1q
0VYed2pwTLKbbGjVrwli1jU3q2iAKSV84M2K2Jbf6EtXg+eLEpzrCXNnmpJm/LKx
FpYteq2fKnhp1h6zdjpbR/rLZdQfh3U2wS1qJG+wew6XZMwuGQlB8kUgSmQwbQ1v
DCc3L6ZdIqUZeXTQ0yfmqIl1YxL7leyYukUmYOaKSqiGNVsNzK97yYjwWm0tsd8E
4yEWTFAqJK86hZfVSVnO2Zid8t6971QlI+KC29/LY5aKizoMC41ksZzJeZ5MSbw4
XUWxrLLH9SoFupnwzxtox9s83ztztlpgLrOzMq4zGZX+LLilu+/pYTKLmTZSyPP6
OvA/cknpirQkQJlZAJJgmNcRo0fsuFaE4eM7VNwQQ+eh/T0xurpM3VVS7ctUFM4K
duNM0+Ky178org3aY9TkuYGjMspFdzVQnTGn1PO4yZmgje0Ss8sEUf+tC4qZ2YK4
EYawdLpW7mok3rkO7ze8GApVT3hu4z1nKPK7UDYECt9AofUYClBSWDBkMSwYhQrw
HJoZQ+I2z7XFebnU952MtmG60Oi3wo+yFCj+olQ2rET+/xgVUK8Y2OF5YUaN6EAL
9D08Qrknx5colBOXdUf1N57+GHtz9UK37KnLdm7HgG7BirMb394sRug4A/K6jJY/
P6lN9HJFxq+Nbfvjdi9Dpn5WOvkPg/Rk7CGI9TsXh8Aby6gWGAD4KGuQt1Z1ji5G
DlGIiBtf05muevRRYkmJ0G8OghqcCnSBs0mQVxEW3q3KKHNvb/Cxy242R5t8zsWB
JU3FyvMdy2xnWqaQoGNkVtMeulL2M6zrpIlu4SXXANOZTPKjWAaRI/TpMi4zG79q
/4yZ5R2PX1FN8keyKwuF/hMLzHso0Mizm9l8ga6pFQBMcTORoUsEeyLm3nJ42hu0
2AUbCWmQWNyFAtGgNBftCtvJYLwzbmfacqljC1jMSJCJNBTSe6KfMRRYNvd54p14
7K38jT044QjBgbFWioVQm+9gmNjNbmBJoQko9x+zhhY+Wwb7kooXdJc5VwR69+ya
jzAKvOge1cN9Wooeifm63HWMsFPOGIAWHCUkdP1ROkUFxits5mHCDelzzdpTtqT2
P+H249yuncrXaZheD6loCYTl2Jqrbo5FafrhLz1FyLOWF350nEd6EbxD7CSnEH1g
q7rLtSLtHpOXw0u5curgSl7kPtZpXmHq0ymBrnpVsgfj0zzOgCTWPqhIHhsvu8QC
XutvKWs0qBRJx5Ev6y6QHRiK8hrixXeBvHPtgFllu9vBxJ4q3vbARVclvRRdMeUH
rmb0ZJVIcM+wLKvmZlN1hRwVAm/EAEmB10lZiK9ddg0y7Mwa8opb9nps7s8AeO4U
uJvk07eDF0bylqffnIt6O5/czErcrbGwasY7xH2VzFqPOefllFe0KIj/NxQd6Yx3
XeUDKS0/Q4qoIFfJxetCWkepT3qpKOqBqAuRdVt5tVQMPYjdEE2JyZ+jrgD3GAgZ
/HrgtRZmfr2naNiGEAIQW5gsF29H59dNRTpJU15R7ETQaMKtjF4VJvn4yiRF6xvs
xQfVVGLNpVpVD670iqZ+u1fESy+HVqMw14X7qN/tF68p1HrN/1OmFpB+UCqr5gdQ
fipC98/l/7079NXaqeAapk1Ysk5v/5KbxufDCWTCFhFqeiFr9i/1flZiNGiEmPHJ
gCg+5oTw0gy4IX0Y7elVqbgSyz9TqQddJppQvoigRrKkEpfqFLSEDIaCOnjOtSL1
Ngw75lszplNxMVVI2pa4CcXfdXHMgZ3pK8nkJHmXSuPrZI5CCCs3uyXMtNR0WQY3
gDvMBtEhOxPqf3bBQK/2W+PmkD4Qj/8UvX9qlgUU00oanU82xaoUt4Oy32jnSraZ
NqjZMDIpz+fO9EeTE9RNYwQDOXvP7BDkNyixxcxTVgfDAP5yBkt1xfFYVHEvkyKX
9nLrRwFdenN4/exWLpZIKPVWQ/0+vA/w7ifTc8TDqD41UZAN/Vi3yW8E7BzdcPf8
2sef/PqG/YsrS8hT+waHkV9rAhknANxrnW5P87LEBkXPorhZVP5BkRegLn+AOZ0+
OYlXZ+qEMCg4XHDBDoXBTmEWwlMQKfvXU1e7Uf7EnV6eD+X2vKl4GREPOyZoE2TE
EAo1lf5xSS/z5XJK/6yBz71WOtdsN2hPH7EqvozDmozOoFseYeR4z2yqElr3Rj0J
l7LdJj/DIADkwXREIJMSMfQzbZ9szLCNDTTTHOh+r2npdX4/cJu68nZq23qmeFup
d+LnIzKvRJtnPvNMB0h290Amgr1Xq1CWOgod/abYWFQ8iZLdsdr5saSw0vpa8w8q
2jtB74NbF7oK/JPHp36nFVJGrF4FwkFWQENYlNSyHwnNNer49lJuz10s2vhqytE4
SsLn4iF6Y9m9jpTQhFHaYO+CSE/DD0Fqei2wgwjDTGNlk7caqe0lpR8ptwPpYH/w
m47gKqR8AS2p5pdc1FFRTJ76iLO80TZijMQAuvVCra+xVjrMDpdglap213wMzidw
83CtNQglybW4LBKmAftClsPTeJ0ZKezOisg7Jq4w7pUCpXLn7P3/wcbL6G5nth0x
E1nHcTVVeQXFOJDaMORa7yq4pRkrybsEfOCZNOinAJh0T5sGMtkr78zeSDxskHKu
+ayLql3yDLA9APO/OobbqOz7gbxZ4MdWxZU3wh+7NvoRc8M5CcrdIipdd8uDQNh3
dQaxtG6IIDxr9yw1xi6DM8Qo+41BfbdjHBkGyitR8U4uQy3VEx8JsHdLxJ+epTf5
/a3X4XW26VqMINnprlR6uRTwiZCl28RXtZ9i7h3dntfU9hju0HmQsqepqgyGhshd
9crzBM3Azyuxlc6ptbcy/Sr3Obk0kWG10HhxH7SH82OS7w6mJY3rUvJIWVj5dEtm
HelBP9RHtXdLGSepAHTEMd4aaTYDXBXaQK6OMBGplewe/1TPFjTp7TpOHCbx7L6R
j3ie/AxNv4tNB8Edwg1Bv29QKMY3nOXwWl349L0GNTYJjmckFl2Mmj2qV7t941dY
hmQys47dx8vDduTRTSLyQKO9uyNxpqDC43jwaP1OuIqzArh4ETRFn2Ykl82S7Fj4
zXr8qXF5BQLQ+cl/1/vrf/L9V1UOldThvwhzGzy+R3THYrwLdrA7PgecxUngzZ1N
t3RIXJQgxfLrHGGQbZL77vWjqdjzuZi0i0KU7vtEsN7EPB6+GpbKE/DaQCxGPCJA
Qs5sWUqi+9X0N+gPSud2mk2JikEF2uy+Del4gsjb7zVizhQDKMweGtLhRkoYJrsw
yd3aUb24bvpW7jm4uui+GtHAbkrVsSjo16ol/uLqGy3ks3eMlQOzeyMj64TO7wBf
+EvfNwKpBR34AhG9kQlDuw5O9lyOij9NgAl9/x9BCnTv2pySJGM92oKZRGu+Ya37
SODScJZVj9vAlB9LANdEP8gYLLzv9THnopn4QOOvpHXCL/pUWTV+YoZY9zSZo0DU
t5x6mQnkoArJ9rggF9mebC0YfRxmHWEcx37pVrwOaFptRSnqNlOAj5tMZHSB6Dd6
nWv0EC5lzMTZTRZmjnRSXL6G+6c7woLqtD4hEutPrduWwO/yxWpc6071nKu1lWgh
KAc5UoLr7DS0dVBkVzJ4Smw2EqUjjmZHyx731YqZzi2KMg7oVoMJAP0Rec4CiGUV
thDAOxjuYTxKDFSj3eMj8gJkXKg56byl+DLY/d+Jbx65sBJAtlloodRZIdbSwde4
FRoABCeyxkFS7mBRrNKS8kBzr9t1SmN6EKr9IelGw57NfOmt1BLnUwtz2OQPiOYZ
Tu9Z/gBOTIzracNp0zBAX38tpj8z30LiSKsVyStU489ZOxAyABTVx69oyrB+b0Zc
8OFo4y0jOBJ4g1VIMs9/xsxjG4HJOtSi/khSGToqbjODLrpGl4H3Rejjeh7bwuZW
t7KzVThASvygF9ADT575yrTKlVrRz0O/lZEBwXE6h9gbLcrJyXw6gs/iOWLq6246
U8X4/X15L97Qs3WmVll2pTKi5xq1I+GIu+T1yYzDjnKgWRVMrgXdHcUe9XELxPuj
5nDYVQEEvLoSrSphaAc0+iQjeLt8OYyZpUyFEBIKDbAgDSmYSuaSVCZOy1YlXB0f
x4p43ejp+i9OC5xTcOc0IsbQlCzlL6LnGgDHKlcLAIvY5MtIEmA79T2wSdaYUPJG
myi387UxIaLHOtZ1VKoRpoveSIwT8fx5w11AITSCBwnwYdCdYvJUvWIv2FrC0RTf
TNMXFBFLwdWMv5/ozcaNpaOskfpgAYTVoVVjCoRluLTWwmWHr17vP8X3ATK4YMNx
hwajNYDJbDlPjP1sOvHJ63CdQMUVRplj6luxjlj6unBGTETpV0TLRx1ytdIhcKQL
B6OY8me2XFAonkQYRcJ02vSpcJsw08aGo/68dUGtT+v/UxpBbUZZ8QlDC0yzMZsT
Up73OwuPWXA16PT5DWlvYNkh7KQ9PRZ7payKRGvmrlEzQWc5+pCPc8bBi92CMLhc
pl+Qbl+dxEs4H5iuPhdj1QIEKZ4uhnNoEzFYJpUAenZWNSRx4Xpsk+ZI97hfLkiP
fWGAnt2vRR515kAXFpiR2NEQ+AlmzcAKHpblNRfr3xpKsEzivqBIh+YFnm1xnZxO
i1CcTFRLbVgYCaK5IBMawavzB6VD0/jRfgmQUbwV2u+ded4vTPy7rQWyFFj6qd4R
iECq4KlXiwahBv/XfYmVllWXoiY6eD19Z8LxEB7cxLQ5ynM0xH1dK+4LAdnflbP5
kyt3F/A4nJSPJGee+A86MAdo9j90xbhyiRdZGLanZKoG4cbzsESRbcfwMMWxZSgh
ez0ew2uER7veEqoIlJ7yp1PP8AjYQqUMh7rVJ/Q0aFoV4K/F8yLFwV3xRbjumAMC
ZP3SBUS3nwAIuKcSvKzTFKBU1uJrSMK83P6gj1EMXz5KZxMgjx2lvgruS6NxDqCL
G8vla0Bh5rdSCQ9IDsNLpK4VDZJV/jQZNtsTG5cw8Pz2cwq3FyCQhBSDGL4ke3bs
waFTaEYNFGaGPPhE5+CsFhPteNAdiI2GGdXM7Rx/RQM7ko662LGLKfoHNR2A2RWh
JWwEx5ftnL3myHlFAOSuS3LrK2q997H+8rzMvSGu/ZlF7GmWrWaeC+7TyMihoZ5+
nrjQaL6+Cv5G8GMmBZxXGIe2RKGFivP4Dt+ruqlDCuGBqBzqbvBg/RXxUWfU7d/d
SLCARPbFtEVp//MsULvCcc2fqgaxtaPagjescqb9BK+sIvhJQFAZFJDseXnAAEEk
gBsa1Id99owu75eB5IqC2tab7PFveRp2nhRCb1czRJHMTUzIMgKUdMx4zUWvubA+
Oyo4Dd3gKmkx9zVGBxlAStldvKoQf5UjVV9feza6ENHAoYCabNtdUUo2rSZHHivd
iJKzZb/03+c0xhfQMERIX9gtAP/nEf2jRhl/ppTqS6Ofaaqv9B1jmfHgHWNaMEOo
lxWY1eYNx8fCWcgnmt0lGgum1woxTa2ykXV0pvP2ZPBScimUMFL6DhsR1iB/H8gq
qN64sN+CnJHulo+3ZMytfvXrzqg73dR6r28T3UEEPu2uV2+pGNDCbbkl8rL0TDrS
MPKM6bTDbghMIl6NkkpL2r8Cb+UvOQn+Qf61XQLcOOTzYHcFzIVOgeSRA7WVW2Tv
rHniGj94YXSfY6zI7TTRYg8PemO7W6myUGc3DbFoENSKyxboe8GEbk3KfuQ4xPsG
tdJ8Hb0nBvslVdGlKSzo21AwqF5w5/I5ltDfcPvx+XxnzqsOhrieRrZ6YmS+5xdN
/nH69hnH3BEV+Ow9UUIBFxSKXpVatsBfL8AM65ApOmNsZ9ZjwcmchB3QfdFAwlsx
hEwQPjdCzl3Uo0qOnSD2S4wnqRO44B3wKqsjF7thH28CZj5K5iNUmSiDsd0z9RC2
sIFcCn1jFEPBJJcchQ6uG/igCdWgRoAfuyH65OQS4km7oT1q1zO2eZQfzpQ+UmHz
2RZn65vxHL85YgrbMbvjiCc09xJyi0WY8NFEqN1l5Zorw4T71NdyakgL59Hl1Dex
UgpfA+/dP9tPTyiKilGiYWyoXdqKIwrOBpfvUyOTKEa0NpdLHB654flVJ3IhXtWv
MbbflqcKLqovRtBF04r0l/a/ygwFwJMUI7UTA03HlmpAxO1lFahOV7Z6D8MXpSRY
TUY8SLd7O4eu5UA16mM2fhglKds4VElPkyeonAuH+/y2pJKrxcWbGIz30+Y9cbRT
4X8fgv8FGPK4umcjmd1B5/VmrdGqd/rJDcMPof7ottI33A03g59l8BivkHwNBiEq
PHtiJKRrt/Dia+XJ8TBNIZ4g4k4kPlnFtzP6Yc0ryhp8DsFHESrks60TBemrWLTY
zhndgjtAumNxexEbcz8Cm6rdV2Qbx6gC2yjHX6tvsd17KdYBqCpcssjmNEvDseJM
eLybeIdndWXSpzvkGXYon2iD2WlBtWOSPG4Q3hiklT1dPfkjQ/U7X9YsK0PE/gfj
vqaOMm5IWUOxWdoBhp10YXDXJUvHahWluwhF8Zp7j8dVbKUZOPZhMzOKVLXXAI+W
vP/BVyX3ypXsUAllWk5YrIlnXBpFt2Yv1GxIbQ0wssCRhNeVYlf6ICb40GQgaMVp
iUWZ87AiUdR6hJURfNZWnT09uQCJn4vTuOGNHoi1gyGiJYBlXZLSFQxRTmgrwyyG
xlj/M3wEmH7xMl670D613BqFBY14hF7NkYYwaM5Ww3muCyJeNVljM+Td3s4aq71o
40UNdJTgNmzQfmu3ebjGLo3Lr3KSVglSGwAxAlbMsqb/ZvprZTlOeBVVLfNNnHW2
3jn42li29xT8HKqWEsfvhoz+zA5Hfr6cHjI51C0bm6SP+pKMuzHPHtZfFMz1Zk9a
uLf0QDMsishsZxCbxgDtKQUvbQdUr0mDi9VhEtpYjwSJqY/7L+Gm6O+kHYacq8QX
Fkb3Cd7b41QheqHUbsAGs1I3k6R+6ILhSfNJNzuU5dFm1glWYrDULgHAyxU2SonK
ZRQJL51BY8US863VV7xHldrxuprUIuFCzyJbLXZI3wVn87m9yJ9gA3X+RSVVwHIp
80c9fOIQzYwkDhd2o7wmgYwTTrTCR/xCXOCI17Jxz4F8xIooq7mbqszFc41or8Pd
oXaN2jsvLwWh4/fSTuLufzjTY/pKPKNBx4K/P1lLTG9y0H8vm41giidZghEv44AY
F/pI3yERgge0vSozN/7JzYtF/HHoMGN4E1yd9QbbzP/eG8FRYNB2gjNcHTc09WqD
a+Dmht5mewmbCcTyBlVmV0rMNZn8aOdwKnZV6yxMMS03/BbPBJeJBk8dITPfH+Kz
UnqxsenXj3h4o3c8Q29nD+710idKpDLcCnuUoLOELcANAEZH7VHrCGVczfC1Spyg
T+YZ63El54ETkbPs0K4OE1xwORd3GewDvGuI0rACA9bFJLupcyMeinpwTWEa9nSd
0CMc5OcIxHvWJmnb0IDN/p7cCLrmr5c/7MxSXf6k8lng7o3I91Cxu0BOWkvMpb/m
SluS4jlm1DYxnPEk5x4S0BoP80yIw2ZtTOfkZsWGRzoCZ+b6uYorP1EFTa52Pw5M
kIoks3iBRCybdd8FvYlaZOAM5jXsJeOpydsz05Z+e464pNkwC3dVdEPIJAnmn5vZ
kDAmuy1/qZPjlhPGoOCEWPiKcdipRg5cm4sSfXOQe217CQDGxsq0s5FcLoC4HjA7
ARzN13x1TdDSeaTAjYaeN72SZqIdTMNpWMNdn8IEkDEkwVjsfC8B1MKz7N1A53Y9
RVY7G5f6cIRfkVOq/orVSfoM/zAExLAW+Z9rZCzqVEZ69fFCLfmm/qV33srWpI5d
yLpz9qpjw3Xp1TJ2iGFU9wSrppadqC3Xj76zv/x2CDSoeWKQsEy/ThPYWgVbu7yK
cj86vDGt28O7zQyisYH1nFLLid60ck+NAsSNBqwnOvuteBXfgwDC5mcl76AgH7z5
flOhx5TbKdo2I+54IyNoeMoio8Mn+q8c3xFuzv1ENJ6mVoSKu/ONhhwAUW2ET+qJ
syaxjlZa8OydgRPRC5iQ/GBH1F0SlNB7wFdwW13ImMmN9Tz+i50OqdQRt1Bys9On
M/7nJcMGBvcwLHJO1/spQYl6AdVSHuzqY99VYYg/MA2+deSK/gnYClrwe6Rgc4qV
g2G0IiCJb0Po2JgIOzqpmNVYWuO0lt1J21vWjWFtVrlm8M3HgYNYqXDqwy/GeGdi
JcQZob1TbmFl/wH9FB908nLKnyYWdlEArw0r7zmzXmqtgVwRvel1gKDlirVQ+lA1
T/ESEI9nwhcB+tUU7xNhm/fTrZOKtKS7TKVkaBTy1uVNaBd803wVoMmFtmo/Tkkf
wdf+6Q5aT2GubozGMhNyoE5smFYRm26RYMHhfitLEizNgRNJvJZqaZrNZk/lL5LG
g1IYVxQ0AsMOmaJl5OPmhQkDnMLFaDLzQjM1ElgmDcEjfO9Wo3kL1ip3bGdIMenY
JagdTVpeOawh4oqq3erfRDLLYoNHnHsb5Al2g/GzAJV6iEPddinOdTLBv1Xl4aFj
IbDWOgXQO217h+jlfVVKtp2k+qgLamOBlSgzhX9TM3y0ySjXpQ3LvF5pHl9wT7/t
8LUV4567j3mTd50XpL+MzWvvr3S2v+U2hJ9DJOFhZ09rQr3dhYQvF/UxixqLaWe+
8EnkzVzdHPie6tCRBAYleMubv/dy6nDcmGKNvxg0471aJ5EBzTN+5Or6yvRWuc4J
XYVq7mT0ZYMnbN+ruvwx8ssggCTb5mESCxpi0/y02JMEzEg1BH7Otag1DlRJYvFj
YLHH+gv0jHFRPeNi5LootXuyghMf3wtQcUpyJwvJJWeCB7bynVAsA2SCXA0EcgxJ
Y6e4RZgOZTVSBIJ+SdhcqpR3X1NushcFIMHB3ckteSix4CQrL3ouI6loq1jp46Xg
gJkoJWSMDrZbKGFvuphnCYl84lLjiKYHSakXUPDkvwjpiNWncet/DC7pU7yjM3Px
eBXtTrQZ+WWdkqChYor29YkmYyb+lHkY6dkshwNAlsgRCt8ANjdK56GxNwnsj49x
g2kE7tvRIbCPmzrRq7nVrhRBqA3vkHiUGZWHY9P/d8ntlOKgQ+aDQMvv9TZarJRT
WkfFU1bzTaTrswnWj/lFLtzNLfLAqFIpRuJHp+UEVKz+9NFgiB9ghNg12zJRVQRp
3PDuMPF/600+1/ixhNZSKGp5FPOIP9QaugXSvvVDM//J5lHS4O8lI3rvw5ECt5uH
CBB/UuE6hmGo5hxvIgeo/b0IGkB1jr4p77Zv37R7PT3f0LstlWLL1lF+B9XUk2Qp
+7xnlJbj34NMyy3HP4tDaL8AVgO3Rm9wc6tyjPsSFunfE6ft02Bi1oqy1Sp+bYty
Ed/jNeB9eET0PPOfOuC/fw74Y9ZshNzNx3AygR4/mGbjchp5znT/CVBtCZKJXIG5
CLOHbHGZE8ClQg17YTvRK4Rp3Uc6ulRzayKmDtvL8y9FZd2xkJtTiBV/M7eAeEAm
V47MHmuRzoffmgtHt3G+Ryugt1sfOgVc/nmTPV0rJFU6HermToE4iu7giBgV73PD
8s9qF9rh+VQnF3np1CV26ckn8ITg3500Q/+rm0O09iidfL40X15gHCnaesd1MH8q
VSSCoboOE2u9r2sgQ94a7ZHcK3guUqCgzMvSrKX/kebKon9gnifQJuKlT9ugMskv
QX/elhFExm3UqQYDQDT4q5xc8n2vl1steaPG+Z87BzNFAo9bq0n4Rr7RE4V6dhZO
RbO3UT55DOyR0YXWPCA6MqRZgD+OJFvfUrgic/YmXom5QBPwAXsr57es5JvdEn7f
7kx4zpPKPYeVHRllP8shedlDIO0OypF5RQiGB2EfmRCNziJjEc7Xj5R6HqGyUOL9
EUbAhmodmQ3pGO/Dx81NuBMkjgJdKLd+6t4uGfx4h1YDNRPJSMP8VlUpnp/kjcQf
kXfU8DhuUXwoMgx9Fu2l6skRFiuT1mdmYquZMlMUO0V/9iWHaGtkn2I+sWv4YJ7b
xy4o157WnZTewthuHUbx6eL8Toa0xix1nTWj766kSNcv7lu/ENAKzEVZ53NyweLG
zSKXguRuhmb6o7xCcARw5fMCtPhDGyX1cXMOKpal/e0VdkPF4NF6hKHrwu5Kpxep
SbH4WTzHdLI7oVTklqqH7Qipz2c+x65DPo7Qw+53QoNvtlvXuamCxyj7tr7cwBCL
ZOdbDD3n3NFOo2k1QUTaPjZmHCnyWgelsQXanBmnDQfzy7+52fdMhdhpa5wUR2E/
nnHEEztk1niSmsRgKv0pxAQbodSFTIf0Jqjj5lkVucM2pf3NpU9u7GIlIvyAXzAH
9TaPuQjB5aX+wzSOzIHXLFBoi6gP9xUmYhBAbdLYtUjyjCPZWWkIFM1zkRQbF4xG
PDQHtbKgC7t4FlqNoelr3uX8DvKm/isunT9+dM9/0Jv3d+iBaht0376srRVzHJqI
vHrpTdRGB9SRCRO/xmHR1akPUNeAv61U5lfrsLkG6Hpgkhmo4kWWGVEZvF0UjPIY
HqeDmZ/me0sPxu4WNNqK7fg2JTMl29fd4vRvDyoA5PM+Gcu0u+YYsTvA1dHQLZ34
2dzh69CADi3b/ydT0Y5Q9aho7LVAreGc5wokzoH6sH6WjDBt5qG57x2Y3hA9lYFy
pQ3MSVaCGRVbgTnvfg4xnKdBGJ92GpAZgso1xXuaRTsmJxeWjOlbFgo4g26++Nb7
hhQKZpgE/7Fmt0UzXPMBgUh0ozvpUtY0GG8Kwxu217O6r9+dM+bq2dxjCbk6JjQa
Y0ZqNpUqv/tIX2ltN/1TgKKBvS/uJlCmUnAv0wpEAECmrjVSV/1jqzzo7Wzua5yJ
mLxLrTB4g402NIkmyXs1tWKs8ajghNqQV9JUIh9ywdRFoOgSm2kcWL2uGbU63c7s
7HP3lxhgt5mCgSQseXSUfv4XtD4PePDwbAxbrGElr4KnVQ7xyYBqQKx12jrMrnLn
P8ShTz+Xc1yW+5Yq++kjTVGYtIT9PeGjkBqr0jXUNd/ScErNI/OQ8zGOiCm4t8iN
gVl99uRxY1eU16QHiDb8VwEbWaRxAV1qW8c2BwVx9esnaeCjp5TsCUEFarhXoLeN
rc0NLq17PyrzHjFAxkGfijZ5DzZhgh5TXZnxcm1iuIzWTICJWHIc45Nv4WVjq7wB
mGnVrf3JQkdYolsPJKqEtlXF6sOdAw8bVUWc3HIo+v0EnlT8vltdUQNQKwhi71VV
7Q5iJ19BExQYsr10uWhJyul+o0M+w05U52Nt7nbpbuT8X4AIbAD+GWtuyZillJYK
y8JqnazdkV3HWPOoDYltc8xXIHeyz7WI/+9SItKssj2RpV9Xv6KsrZpXPT4eASeW
BQswXQe9oL3EJRwaWK5bEKx7VWWeI+7z880Nvn2FnYu5lczC4xmwF4R/4bwBd0NV
HvcSaBoTSVPdCObJQgM48cuzTO3DJWl2UwqcF2NtRfKUzWYCGj06I9zMHpPl+wpn
yBpsFj14Z5wxO4ZESeQfXaHiEHMUhwoiFgtNXmzJKnyxJR4+GlAZw/Tewewy3d2m
fhERo5bjAo+0OVSzBwB+jLG5CKo/8V/AjiCJNS3uaZnckkM6jJqXGH+UqkJXpiwR
VBgIBEUQY7VL/21+4BazoDbM0mJRJi7ZVUD7P18qpwJmkf55YSGFHbr1E/SJDOWV
yBNw3D64NeSxkTtQbdDRLaYg3MLvOTHG6m+5GcGZ190hYOp5lQzC82hA5+u0QwAi
CDvpgBwq3TbGnShl7ZU2y5smhON4ZEXEBWeMe6gkKul6bxtBSoPYeklemfZb/np2
oFTdkTpPWjHSz+32ND9hx2XKGf758CYkk0xSO8HMJV9ycpBpfR3Hx4ZCZHiCT3KJ
I6ImXMFfsc5MHVfGcB3iXSXKjy/2B5qvNvfdNaJ5nEYsqQz02ERJbgoyiw4NB+qL
8k6zHPxX8ohDhD6pvT5S1QbabCdGCljRp/NrvBT+s1PAVGxmeLlafscIPjbHQGQA
LkaWg3vDNno2abV3hZtoarVfRY3F8Lv/7KIQo4HjPM8P5mZY7J34t6Xb2FzUmlLl
iAD6EqEpVhxyZJr4kM5VSdw7n+RozXtxnfaQ7+Tv6MR2RlSk/N5ZECfa6EzUeCBS
GKhNqVXMpNpzt2DcdQYJN/PIWGO85U3b6BW23lsH0U9hyEufmS8TAu63MFCUw51F
60f3xYDVXMgOsGzh/uRKDZZdmEV1rJwsLCoAXwoDufFihaHN3hZG2oD3EO2TeHa1
JD+a6HufMGbyDWBLmMXQiFdueIXXka4h6/P00Hsv6ntjmcFHamEftTvmUWmMjcm5
/ARwp+P+RsksdFXWNFz14b4VmJCyoMVKOLJRw/LUmQGBXG8zL3BliH1ZIyUjEJAg
SBbEVGowp8EDl6aM4p3DKh57F1/ibDyzhCqewZ55ioXCEeWm/EyvGEx2kjFF3QGb
PpMUee/uB5GVl6BlscMyqI77Jxx2VPdiowRq4pUPUnH59u91vD0OYrsIoojU6/rr
ff3FMWlFGtrRIiw533W3JRpd69+ZXCCGvkK57KNvACNib+N9YLSRVHLj4bkj4Sp9
fCrWdc/ZbLEvQMAkepoeW60/Td6CVIMX+pCWsjhwktnfxRJCPsali8OJAWNwYkNB
r6HVlziH8vBOcSKE2O/rRaVUpmh4OeoJMYlb5nKn2MIMRGr2LYrssjw8Xwx/FIhm
2D4ECiq7LneUJ03FBEN4TTH4tmqxmM1krzrjNb1okNHQDJoUJlZocTvOp4wOVBa0
iOh03xImGYbh5t0ltlRUNE2ARWrNUZk5r7d6dlJ/7NgtkOxxgcL46R+Ig2g4Rjmt
ym18NTbIZlE5xAln46WFktv+TjSIcVNTqPjM/w7eRCcxjy1uUp05CXBqYxunR1JN
cjnl73uj48JBl2duCe40kgvYV9wDI+6XGcNi0TZZtJwkrmjcRWlyuTaFKxfZ9ey9
Expe15lPYCyLJlq5YUKPH/aQ+TH4bTwcxm9chawNe9WVD4lO46SjW93AeIbfldsa
/6uPJbOM51zXGARMsUYkgVdeWTwUDwoYmL9gzKb2IAZzqyALuK/pF7KQhf3Gid1J
RevpTzrcl6QA8QPyRABk1KZxWv/MimoH8vQxkDMx83ol/h6oA0jLgicXx/czJafM
YtvbEIRaGtivEopUV7DqC7AGCjMjBJ8qIJ/eg1AkpyMI8N0RmMzdlKKxPTFoNEEG
peNgvtSMBT3k8fkN/CdIciF+ce9JvyekVoLR+OClUoE5HJfLK8/5p2wAjNakGXbE
Xs5kj6E2u3b66dHfjLj3cV156bxIjp2qADbZ8FlGCplhlkQ7JCN0K7ym0HEP5vr3
ybYQviL7rzf6GpRJfOeEF3x82li6KUBp198CoPuBOSag5yyUlbnl179Exll3IKIx
+yhJCbdfce0jUxSrtlN6I33IfnLQ9KHA9boT0fAodLQANs+BvELXK8XJg6WBX9NT
SfIxqH0N5GJ0koEPGtgbZ54ntw0/asUpfr2KltNH5wz+oBDT5tr1/WPP8aElxAD3
GZzJlV7FWgIAYRoT5Q59H3WLIAVzK16bPQI9UwI9cTLju3pLFsgHMwZYtk33RBar
sk9BJZwZJTERbt8RzJ486otjXJXNOVaDNU58GEzD+K49+C0ztuoqOM45abNTTi7g
vTL/8HrEiZHsXuclr7Z6qqdsql07jnsOgY+nNvdbTQMu32ogfRpUfMoBpw2qRbKx
vU3Umz6XDfoShAHmduYrCMZCoVWUhaHACDhCSkzej7MicgFSgTEP8A9JYLE4OpTx
6WO5IEAlb4KwI+aeSlQuuFgJn6/EGvfZQX9hly/9XAnwX+9rG6s+zyonnat8wSwS
wiyZZx5NDluQL6M03Kc8jx3btg9CiXTZbNCK2sHHNALFqUMLw1L0lCaLZeOGAWD+
1Q/U72v1uv7CU0cu4TKRwKgbDRdwD++FPrEpev5iyNP3x3Hng68pwRei3joYz3xw
gVH4nYJJe25wN+JlqvNjoie9T44bAhT0XnXMJHWYpqcDns13+UOT27lBtjxmNqc8
I/Raiunbw0ULoYaTm7DST3mWXyNLosgxAUOZCbbY+5C0raakDF/iyVaVH8S92sU5
wyGfQFGi3T/ObfygZhqDfUrVhDLtX7C3mtr28HJmdHaLWNaMMig255xUPCLkNd/x
jnEz8/dkhn3PYRQal1raAk+EOpAiD+vhcRccx3vYSo7GMvvh006w5OZzi4peivDB
Ti5LUZThn5wL6dWW+LSUhQP07Na+M++4Xz7PqX0VIhxNGIKXjwvW+qinqGZOfr8k
Aqov/Aq5SnVSOoBwFf8lex60uo9EQXU2TEcxsfj3u2q6IHTpgXjNT77xr3xBwUe6
bPwJMWm24RCyIJHEqHeWBw/AeIiOpRgu1lpVYOLNLWLHO+TqhOho/lhqSms2YQbH
HvE7hjaLJofuCr3pmYfdbDjSaCJs/E9fn5V8S8mirCBo6AY78IxYb7ts9xfMaRtA
7mabJd4CiNlVmB5bJuMaBC0iVjxq/xeH0YhLFl4qWuEPinFXNDEP0NO5T8c2vr4S
GFFZe7OhhaKsp+J9nLIIGYHNNRQ6gne4EAMaGe1kOs4EJ4L64Jproti6614tjtHH
ZcgZWGGPW/aGF/U8FCBgmujAxZT93f+WGxcUV2XXeJtG0cKX+oPlIKGCFTHsl2Ox
UoX+kn83Rnh1tKncmJtttX1YR7EUQb3oVa0y7tDXL/AmLo086Mkr+k2O0CQTBDw5
JDrUaYWzTGTBe2aaA7snBy4/gYdUtlYuEWy6dmRKVJ+os6VTy2wbRS+1JBzWVFUG
55ErYCry/2fWfiQPYogNzBCSfj3oySKZsKCypRb3Lcje5A8+WLf9EM36BCDo1vgD
FXRhEYprtyM7uLBU0pHfWMO7hahp3ybS2Y3BKZ2fUrws98wmK+o6redIbYVU8XGN
65iQXpA7UMTLQ9ete2uQwCzWqKj2lAgWBTVg1Q5nzGh3tBrQgHwICYh2cEyZVGME
VHAAfVGv2My3P3a/94YL4LyPOdqIL+xboNXVh1lm8rGbgsfB7u5bohmbLuQAtzB4
+QsbWBrMMYBUxG0+Bp6iP9Mbl4iZsILiyxm4vBjACJtI8NwLEyiR045ceT3kmOMT
dJ6cwMAZ4en/Pxv8CvBTE2j2olVMWtontvroWl5zuWRBRLNS0rCeWkNLxfnmF64W
WBXcIwSYwcArMpyHoF7gsiMIYodIramvx9/a3o42VOCiLRiFNxdSDgYVCF4eMhjU
fTwcGlLd+R+IjKQ81Jx/YNnsDWuinYVPHv0q7RxLdVahIbUid/6kMlZweIvuXwlb
Absi0CV/wThYU2/eLnTWbgbEUwPNv0RBA9mjxmHNObwdxzX+oP8hKK2eodEmzfHR
dl2QFefuABFitgeLE7FOyrboIGXN08l4Wwv1BzdLU9WCjQx+EqESO3/+ZedeuXCW
jUf649v0th7FdKY4GhK6IzCxAqz02RU8NTD4tvJ7hU7uMID+lq95LkSCyjQQh3Id
9wP5PcoJ/OW5aYhz2/mAFsrhbw6d8jYkG82QfsyTNbLrPrGJ2nYhArhHRyhaoEKd
OObOclCFybdI/qiqpJxfpLw0X0EHQK2l3PQPvgLzZIRgOecHQLT9vZJ7DVPTWQOp
ucL/NObdv0hrsjzNGTv3Db5HvzF31T4HhfwnGezXzYSIBAWZWQxJ8L/N4eswci7B
5oKSRCicZN3isTZeddrTrl+OyOgrhbOJnSaOyJxyk6lXLJO9o0p8hM4C4tGQWTiC
Z35D259aLE5hfAGD/BpZFQGcOYTrO5od1Ph9Oe81unBZeGba3f1JJKQkRJpJI3nZ
LlvzF4U0WePBXTxjg0Z0s1IfITtb0rudPznMseovNIByYoEq1d+5mXFGbBlKYYtu
komlPouzdV31Gjpuqym1yDWr6jk8ELPfZCJilpiIE2pBKgh+ZyQeNwScPQ5IeQ9e
F8Qk4OtJZ0ymEL0HUxD5XdmG59yNMQLOQnZbWnMvjjahA3pXcrQAhvbes+KgtCwz
fFru/ZH8gBSXARCcG2bPfcx33wf/uVVr7wf37L/WwmreTWouFITBCmcLQptP5RdL
s8Qpl6G7Erfi3+ip4WY1yKIdVpk1ZYEq5/G6JvRGDQze/yfQRp4CJp9PkxPkKQs3
wVE8SZ83iz+XdSC/+cRqMCVikoZu97EeTHvOP2ID1hLhC6LD/y84TdsnZy+YJsxG
HQYGdU+Jsz3qgRr2bMUR2ja4kvnf5wrAPBFr+G+Sp6fPrqmpikAOAr/YVkktLvZw
r+XWXxMkxfoEtewTqHGroZGrYNgAZUmjbqhe2mNPoexgAPhjmaZcSDACAGh4CsIg
GK7HD7Gqc4LQP5f+EI5tzU7DI4aTVkO9ZO9ZvC4/zNh3hHYs21WY+hLwvSZtgaD/
91WfmP0CV935GV1j3sAdGQ3AgUQEsAekEwPNGDyPZxwZPzdxtpDECEq91T7Sf8fx
Fc4cgpWYDZI4k6FPFQFnJ1vQJFJQ3gimJeNNFzCrPWG60XzngI3tgjL10/ac649w
9yJLkhwBEXOWYkVi+OQV3aOmiqK8IwQkRSJE6HB3J4aeWDN/fs1pqqOH95SLPJjd
WkBPrSZlw65lx52NqjS8NzMlkODD8smvM3GHvDiig7uQOlc5dd4BdvN/zLNVF8FD
itJfXHRm73HERCgWSNBnmEss9hI3xdAsVgzkY/+TE2QgAiWkmdDOGvqRKcgn/rFK
hcyDB/bUs5rFiRfgvncUrHAVh/fk6YsZbaSVR8iKhkCr1n12xJCH/MmgXxHz57Lu
g/N+57ggRMf0NM8nqbwq4XHLvZ78R6Fe6X64ds4wv/uMJAZyawryUASbxvlr56SS
pqLwosAg/zclmZiw/Db5AW1Ic1u7INW903J7lA7k1dV0gTsxTO6ffUoYH2ubYQLi
AfQOUaSFcQt4Dy9S/JUf3d6kvBuRBujzNFjLZosoXb6dTUtBnXKpv4ZHQTpCxJEU
pfi09Y7b/t5N10RMzsYj8l5SweVCzXA9ohg8Wk5Fwfrc7EkjEDb+sIKSdtDJhAHD
6cGPlLXBgUtewYzXVFh4apRo6X4uDKWHDtR5BOTcppb1vpbQwndLrV4VqgegBcIb
8gx68RpjJXGCCDMLeDMLlWDMXduVjR/2rQvHdgRHA/icjeZPiNqMDFNvWj4MaOSh
Sem0WeD1oPDQgf200QpQagC9FGLPI5jYpEFBQDqS9J6n1/jWetoDTIgW+avfsDwd
RVQhOn7YF4effPb7pWpcQRZ04eHtBCt66bGUkbdZlcN6K5gEl+KKfPGQ7ZaUDgI6
nSV9VSP1mvjS0XhlHAwz2JJEgeK5h8fZdkGum8meT/JVgH6BY1s+cNq58KnkMEZY
MvAg/bYcfp9M9BwVdg8DNQn810vG4abpmB7MLxALV6MR0AgWj9yd13SIfuqqApqu
DAO5d1QMcnufQaumve4hQ3ntVOGMvZMIiaOJb4qFly1euwYZkx0/cyE03VGVOnZa
L/1gpfcwO+RWABWyl5y1p+ix0RFdg+7MTW+6bryiL7bmcPz+nDGQxnzeK4UJ9fbe
ShRCUjqEZ41iyWAaBib+mO4rz1CV7i6M2tNpdSxoJcGj3bGauqTEd3Wbo8nYO/+3
mZc+xvgZ1gObBYPJTaJwE1hw0AuUfmNB3oy4/ue6dHhlmcMP//AAcAf3hIMWncMB
Ng/WjtuH/+i7fEzXSBCzbii2daWGhup6CZ3ElR+cuKpBwecu0XUdglrDkdyxN0wt
sEkmfHdwHWdboGgi0DmKiQX27IdIfkhcFgjexMVQE5YuXiiuXuLQSjVBl8w1gQwY
oDltr/kB8RlfumbNwAPZAxwGBz7IRnVtahSeEUynfBb7CqqRfpwr2+Dq7vVTz/2+
sg3iW6H2DoKceug8fLhbNzMqOBBzjxF+e0gp2ZINRUNk4mbPXq3BcCuQ0u4WX9gB
5O+RKESIGdixyrY+cPrwfbeQUf73JAsP+XHDCYURDqe0vYNiTMrR7wXd/xkvhoSZ
Emde1U1hml5355JsqKkx8frrUrMhwmwI2W+3G/DiSFHwpbUkMusTo+HkoPbU0h0Q
R8kwdlT5j18qWPdawt5GHZxkfRuYvltis+8SDpoenoeudsqR3/nuEdSphLHXKlFZ
lGFddCyP75F9ElGqT8+YNwdEWeH1410zWVuVJ1k7EZosyxlPooUL1dnPlVb11QsN
QBXee+o2GrRyCXC2SP5IaWWBDFpK+O9KqEIX1uBKYqtfXaNGedgYVvtne+R1RiOt
Gw7iVMWJbLcERIEJUikqw1EZrUz/6pO8AZ8aBFAb8U3V4QZ+Ze6OAXNSCAbFZl67
lwQePcjjom/gZiUqljpbXkH/I+whyIYC9Cyt0RYmUVsVNq63rUYPsX6X3Ub4d8lI
Zl04pUuqGDtuZ2sOUBd500brjjpB9+swjK03lE55gSz5RDV/JyFngX3doRuEx01Y
OCV6WRlVn8ivzVTMHHjWRyECxGWcK7Obgrx+XjpMBz4JPi2p0VbfNlSpQCqYgmft
R+EkyJJ6XkPYPeb+DU2qw5o9Pnujzj54d6JOKB8kUccbDQ/XTKAc7NRujBV5FYDn
A0fjH0IWnw6AYZ3dvb/OliU9fughvxdBMUBmOQs7vo1SbGy2GPQ8yvh0Ro2hZ2To
7aSgUstpaaMO/jtjcHSlfwQDA5Zd6LmqUaYpR5NP8xhOC70audz0cOZGDF17iyjh
j7hUr2db6vx7rzgUIebmH7p16H/w8RqEwsBvOjBm32Qbs01ucUFckQYZPZl1e0hS
yynYWnvJtlc1X+Lxhqu6K0uDjwRB6XRlhih36AOuHMDv3KpfU3YGK887+JUvr4O5
YyJT0UwM94ZGQAaabv7tP99cj5ygHYWkGYVHa+LYOHAc+nwYUt5/I4pM2U3Fu9oz
LB642nqEBDG2YVKJbfDfBuZt6mj4ImRlXbkRLD2MnH9dF9dFOfA7k6NabD3cUdk9
4AdaSSlPHotuUSX3TqK0TyPyp+xGM7Z9eKvJmXJvCqw0YHudRE7Sf4M5YejAnASb
M6sDu/a3G3M1vUfcUQXispoejWSUozqcGlNxSPj2RU8ro8TALjKuRboTv0s8+a9J
aB31QNccrB6baWxk8g1fI8gK9NxvPOMKofmcS7U24zkL5dMSReRHaQD3mbZXX5BW
YqPYSQAfROvIhkjYVmp13eYktkGOxkmG2zwwaUmdsCzC+iHruLI6UblK6c7zFm5i
kk4aAAoDLv/jengsXGSsPu8m8yUs9pzdDo2f/OZzF7StC8KBEo9Maofd15owPMjj
XprAyp2wmIdmsZPTsLGf1SuOPu6QmuQUqGAahLIpczMBQV2oOTssfzPQBT1vYBq0
aeIDhqtD5vYTW8siDz/0CjV0dEy2O0Yc2qxsMhY079KUotQ3+dONJb8zK3sgoqro
eIjACNO2vG2H7iErUW37F5ktdk/8WsHv6D+VPlbTUrdYKaMG8e3Ve9hql5hNlGS+
ulLjukq20z1pq1XaDKmRqUUcFTGXtLzwl7jD3SxLfjETYR8A4U+W5ciiCwX2V6HS
7dhWh1EUZqY3FjgOHg/wtbiotwFcOnHFrSZg3EuIfLXxcpCTFwiLGb8bOd1tcyU1
oLv07lAja30Q/ZdUJo+Ptf/EbYhpxiTjn3tjTIfmEveXi3Aa428k6OiFTGZwYV75
+u7ti+UNS/h4s8sRetNSpgarWsTzL6OyS1J1IqEMYxLFAS5TJcEKjLJcyhu/Flsg
Z/DGnczcHv/zU0unB/Nayh5+vtPqFDDCRzfiCE64A3Sg7la+dJalUjlNgBXSzn/A
/Wk59bhlUQAmGTz8d6lgyuCrcolDtwUDQIEL8RBsar95sRq/411WLoZBvUv/RJui
mnenqZTsa+I+/mgC2m2v6K0GkrGlSfKaN8USTbUcZZAyerxN0ygNYnylXTRROfiI
Em2ykcXw05IWhm54t+JNzKq1gPv4AHcEMu5iq/0ieB2El/nwb6emniSCZUeElByX
XVIJhyxxkfpOWOR6em7EmD0PdIAIQynwB+iHGWt7kBv0WTYCl6hhzRer/vJtaS7f
LC5ZvLDbQhtdf5NRFE4+Bjwc5NQPj0Qz1Xk5QTui2hsj/uU3yJrOG899iWVHR2Ql
N6Ksj0HurggT2fGoYbUadhCJqGINp2h/vySzwhxv55tUjGEJhUAPjZz0/DQXVFg/
kzDUpCmj75rSLmPZxRicIdXkPeKDf4yrXzw7XmMz8edy16k/VAKH7ZeoeA8XiMgt
+2QvH/1HGFHQW4WT2Ww/2/N3jLrd/hltrFk9C4kpuIhTiWKnUde6vkqwb8EN89Ii
2v034XwDHTtWhuQF5uZoJ6n4X3MxNiMrnkt6sQWaoiBYfz9qUgUuxKPfOsu4KOGc
tAXWMmyioAqGXvfupAZI5RDRdLvyOhmaDDFY2Yna2vxZHkPIMJrESSFGCRLttmx2
Cji/dY8IrC/w6Pcsoo2cjhI9uqhbLLO32J5YwoxHs5Px12XcldP7U4rhSaiC2Txn
zbePpzWpevV2Yuqkwcm++42Fma/0JYkETW6u9O+Q9CLiAiTedw3p4f23yhZziAAM
HHcLPxya6TVAE2Yz3n0oDZLdn8ctPLgxjbrEhMg0E88cxe2uJHlgXHV5YdbiNRgN
F7mCs35P/0ss1CZzuJF6RvHrmAcApP0FnjH3Q24y1E9fXwtigJ+bYqjS234rk0iB
QRo2zI+EZy41hDI31Sohyw+bCRD2ljmj+HJsIzg7LIggdMg6CDBoY8000qeXgZNv
rEjXL8TlekXXK3b/v8Ji1QPrubQIBRLOU087dsziYIx708Zk+1UPahSt4/WCEAeV
BlAgId//Ex9nq/tYzNSSpWrGnyzy2bV1TeTBrH2sba+EWadAJPKikyzr4bGoJrZD
mPuyYIcnIvrn1DM2IRcwaAXn94uM8A/c7m8ib8orfXcfxG6of4RsZcNnGo1NB8EY
E+77Suz3EDxV6G5eCNC0qaI0OWkb8mA+1Qa8w9ncSyQO+PGAFZXhrkAdd3BlRozF
mUS5uOqvqs+Gw/GdHY0DqtyB8CdBffltE2F7eLqhoPatFQYJkFYEk1jDqm5+Xbc8
wdAdqHiyLUbL/yvoqZWE8vl6sJRc2kqi6Ht/v47oGnbgWO6eir/eb974gLUkHZIz
lhARYngv2nmCkij+gH2qHHqIzE88e5bJa+CGdP3HOZSKlJ8hFkfHb62KG8P/eIc9
LMumKN3dy/mc0BjD7uOg1BBeeZVmIkYrBPhCN2wi+Dk5VGVeus7Bh/uBzwM0aDKb
rL7QCdyjpwCWzI5CrHqOPwobba86lb+ur8B8/kZjm11sgNQq0jDwMyIFc/9/of2H
qfn7ktgIeBduS03gwPzauRTp8xkR7gSKrKF8Mpr2kK9ESwAr0tEkZZ28tO0e6TIr
bXJMqcWThhI/Fj/o0sbrqRL+gcxqep2FOJW0w/ntbCmlWHPl7CUXp9ovZUrQ6VIS
HnrcytBhHrjdhrd2YlwacY7cyJDv1pa/xXirRALlY0s65mDFYN1/ILn6J6OfPJMP
/8MDyg2SV1x1jVscIyHYIuBNqQ0eUPHve2aI2XgY7e6DsKq8frPR4LVk4auOBd8r
+2upm75YzYm/iQCWiBOGI5bsxQ+5LMPvjGgOmgM0jBcMMXiQuwcjEY3MCCdRlCK5
EInF4F111MXccG2O7rwSUrf95Jn9gMJ8uBUBKQp1kqqVzH+w2owAQKmdRbpYYUz1
E+iR7Yj3DwCFS1AqFPkvW5hSozGFhss5VDiYwgRWusEyR+rDkHUTSAskypjCmNse
JkJqYln4Xm+qp7DLS+U/GVP0bxRWozNNY5Ppr/WjKKuXbSewwpLMUUVvkYGoSf0u
X2qg6tRqHk7iBDoz2G7Y3PMav5YbsCD6ey3sXQYrWzFzIoBa28DvGytqLvAfXwfV
USZFuDJ77a60eVuaPEcbPMdZilMGg6zBkiVYd73HmT9ke2YN7YK1Lo94yOAHvLoF
Zr2mixUYOLcTs72UBWPGO1iO9LsZJwwQnhevi+yxLBCVJOHd3Q4LpFhTUeWWsKVK
LcVZOj+Ii3Kmcs8vV97TlN6QvGlw6L9x3UcgokhlYLDIi9q+PeulcwIx4ghjen6o
83nlFaQbaGdTYJzMf0Te5IokJnDA3OOKRI7bguauWDVXOXA75506vXfwM7u6OiHN
yvACcabOVwGWwC4S0KEp99LoyEfo5vTPSY3tQFZZj1VmtQa0KEgPBUSydh+XenPs
a1p8DgH0SHcJxl+S/mbQ0bNhyMFOg6HTRcqwOfEXToJDheNd2mWBb4I1AwZgeoar
UFCRHSllVAFoI4dF72W0gMe8IlCc1T/W+f7hIYSOJ/ot2Hgelk5VKlAuYs/8ceWG
m+SkEdClgA2b/a/03VqrFHzabQb4gLEY3TvhJTrTRgtiojTQWb8LjApXqUU8KrRZ
pyWsf1Oby9yK+/y/Oo9EhVL97FZKHAyB2O5MMqCpxJ9TAQEKkUIto2qEQEcWbrzZ
ZvqAbP6WwEZYjLNbj2JP2dP34kq+CsIpYEOnk6+0FKy1/3itAYzB0yFSv6+voTeB
cgW/Qxt+EENQQFqsAnIltsdbEIRLWh8rhzJKxVFwECo=
`protect END_PROTECTED
