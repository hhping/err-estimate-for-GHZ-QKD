`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6X8mHioelfa/wRbzpLzHUUotV9YB4GHPWEDC9fkpU7LJFSH/ue886C9ZsYj04/e
xkzoilxy+pGgZYnuiW41DXFiEXeY/eZlXytSnzurRfyHocPMNYRsW4P/CGDVlYim
A/a6arIsL/hnQxoVwabZuy8hjpsCAhLtlvpkeeuTWiSJw79AYrYYBhBIslOYy7D5
JbBFFZUE+hchAa0XNczAmFWvFDSrwPvPt6YDNShjeLw52T6eV4o+6yM3J2NP4Zfk
THwnBNo1t+aYlUMJxKi7HlwvmNq2cZK0ZMF9XzBHK24wKCNt5f6GPhUHccp4cCDq
YhppH8buUcCQAMd0Bv8tLGJae9iADAAHU4FgGc2ynebrUWet116wjvlCzT3u3Wqw
VeU04xO/eFtTmWbp9WboolHkL49ga5vE++Q47X1etKlRKJzLqE58V5xKBRRALXrS
3dLLW0ofcveU1uJ8Jii8bHpvRPLr80jKHyjfCmv7Q0M66b39eLCY+U2ILfnby9Go
A2dOyUtHpKf9Pl4NHfV6OkEi35Lv/Q/BbcDiNGQSxt9M3XMK9WiD+siZ56LiOIx8
JbtGbMIA/Q+9nHHwruC7Fw==
`protect END_PROTECTED
