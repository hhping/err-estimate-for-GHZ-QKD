`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYadizw2nUBqto71CHA4TsvrnUOofa+1Q/1tEGx+ZcQ8iSRp2Kxo+aEZm4M6+yto
Sm6PWqS4JjT6OhF0TEw98Ut1gMULJ9tE8bK/h3XSdKVm4/diOomLbBluHtHCrEQo
2JGzbVeenPAKiildIVDV8NeYkCjm2EOD5MvD5OGD6dw/VY355Ijt4yySU149JOdl
Z4QPLzGGMIGszFVjTetyYlU/svpHJFQjBst054XLkZy0kTMNBN+GER8D5qvGga2x
VozZXhbc8+1xp0uKilU3cGa6okdRkEzTVdRmulAipCvecwI5HFmS6/gAo6BzG3Oo
/ga4ZvI3jhvYRzdLfak8f0aWCFfaGd+fYL8IwcpqfO+H2theY1WxHFhNsjGVi8mV
s2CT1rmWseXXACwJyjR/1pbf0gVQSQIDPWuEBb2HLtzowdvPMJGsQf3fKOCts9uR
3R9whvk2yUgcwcVS2I3kkdKJghM/NF31hgsv5aNqsJYbnlzXufXTHYu0F0kk5XZl
hfIzZbvjLUo5xNUDGmyqWcc1OETDLJQ5Me7tCoabpivX5zVQm0N01xXXB+8Zfvcx
q/IYy8OuCxUtGB+NEJ944VRm8X7agRvOpOa+SpOZ504yMDzLoEyGG5zWqe8zFc8i
dm9bequsGqgkrU2u12pOGeB72oKbM/T3imXIloFs5CZwtQtgXO7dQh0Lj7rgiu4i
UVnaql9MS4GspVBkQlyfSmvZKENsD8p5xwMxAm3IE7I8wKbAfAM3+dBdkcQohLui
`protect END_PROTECTED
