`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwRvsTYAs4i6Mq6Nmw7j5j58IiIdCawXopOLFMVWjL4ENknRi5027tEH8LFn3Hip
DLoyLPBAk5vGpJDBJl7T1xqqOWABZwlyFS0u6JSviqp1gqoA/ovtTpzGto2i5G4y
wH/m/jeoVg1grHK4VOF52nfsdNP4dudWPkoquwOP6totK5INkdsQSCSHqsb3F5tJ
hojwkk8zeyI3C7uFezW3yDVVExxCf0eX/t6/PGCD4vj7yGk+ghuMPCkeTGyl9rbI
oU+RwjL6nNlZLe9mQr03pbNdsua89LJ+gQipv8Shs9TqBNIgk9vjKAAD1VMVR7EG
kNDdALOldq8nT41VLY226t1OJgjEDiZ4p0iWJt04q/nZnQkms4ukzkbPWvyOLWRG
30VapShEabcHFNW6lUPQkuCWXbSvx3noUDAjUnWM95I6H7Rc7XDNbMjaPI6yWpjl
H8ejH+TCVTGtQcw2PL6kGO23PiMi1WCDNhmCAU9xUGshQ+PZ1R+35zVhQr0nDxKU
v57wfDjyzJJ0iWSG+DNd2b51pezaT8h1MYkFFoCvSDQvBmU7Z8LJol55RM7oSpof
YhyFmTkKccT/TLgpwPV3gmyTvcs2ruBvfywYeW8XVuGwutWkFoDmDPtMQFx4MXbH
fWo8HcqZ2j+65qILahc6jSmDQm9hVWX5U3kpCfTwW2tLoRccx6BRN6Ddv6I0+D4m
r2A1GFIhC0CitVU0uz4tJCY5Qca78drZBTyEgHaPvsN/AQKQZmxAVp0U3YiXQ0sI
y4bqeLQJG3qzwcL9QeHNccGbj23Y9cFXlwcRtQhw2Grll/gtY7kv5XvQqPzhbp3i
TFIr2/7id+XAIF524Eyqo34d3MYy5CvBl9QvPh7m2eodHOJiYTymGdJCFAMmb0+t
FCRFNdqEFg9Wk76U4DcQzqiREnFF+gRSCdLB3xnOucbPB+HoVyE7R3W/DjA+PCK/
uCwsLs8PjpGTdwb5qDL1AiycRLtWp1w3NK/kMURcznGr05AEydqNKaf/QO/FnUIf
mkGg7epItr5diEuuypTL/1QXA91kV2blHCVObbWzFOGweJySQ2qXduyoK7R2XG99
mDbcFYqspNVjh+rg3+aha13bMFaPNsYzdFqPgETrKylHQKOHPoWFZauLxhkWLWHq
ObxsV/ziXhzRtpDkKRQSkWfLloaegQ4RLHtW0x6L30waX/EkeggTrpfAAHtDRJXM
BjdTNAjt3+QHo9uJAVbMYnJ4+ydIhgzP1+GA8yT4ec5r4Goi0YmXLO90Z3EqA02J
zqdkaRfqql7234RWiikcMrU1/JpD4NeuxzcFP6bYCPULLhbQLu7iMtc9sJs3Qd3a
qcMgCxIoYBZcBtnEim+i0HPXcA6y5U+B5SzfqBPtcqd13e1otSyDKocFiuajjIJD
0uhQL4e+MGcdpjEiKscJFEpQnpBZ27PLIwui6sRcvSsW5GhDjk5JME2vFHnL+xlu
HZAgcMdHrRMvIraYBvH99L+qmXS2TKzvqTosLh156x4Tbq83nts8jvu6yuo93/Cs
OOdQdjcgLjKJTtEG+OuJN0UJGERZtC2Y/g7z5syVmGMZaNi/5QL1R6DBPd8x+pVI
1JkkcHCAeuSsios2EhdaMYVRNyumHmN4+QlT08pg3ZUsZ9BZrFCmF1u1tvrONAKz
wjQGbxC0iA1g4XIOf9ixIDAkBRPOK2f52teJUawTp0JtT+qO7TFIrctI3VqoGSNn
TeYIjTYMaDIZ3STbNwFEy5e6G8qgD2/AAF5mg42wZb51Ts88bYmqRO+64AYQTJkG
fYpkbOTEJqvfslUqEYpgb9Rq20aZOjZbQbEYmIFbL4aQy/xhokuRGXxs/mH6pj8k
pvaK++OUhq6hI2sLyPOGB0fqPapJp4mkFUwS8WUh7InyUdD628GP40LPsiBY6z3J
aDbA1E3POovnYygggtTceVBszXfcmsML+aVTSkbrzW1jsF9Ffs66pL/AhX0CioCE
T3f7zliKo5FIDn6H3X42Ea3rFmTmU0Pdvtg3RwfNH8b/v8IWfthkYzxnuDDy8SKN
SMcyKeowVoLPMLKJbOI8Hv+ugsMLjttuBdT7OFQDLHI4WmO3z9WD1jSDlPXLokeP
fi3wqsHWu+u0/ZxJiAzinT9CquvxhxMoIY7Kx2Ep68qG4GyEaDr2qFEZnV6RxBJJ
zbNTiFz6PkX5Bl5m8FdiOJsWvkk/PfdmQSK2PGlVhwjHIEuImzjHLSHPsmSi2B32
obA/78k1Z8MnKI3otqhxFpgIW43/gj7wM+5CgPoNkdOa1GuhJpoRCwJfadqwV4U2
WODOmWlKBpxWOhjNirKNNxVtJf8emmPMgIMQDLgit8EN+6EC+94f+/tQbTyi0dY2
ui+Ie3UfF3iwFDokq6GRM0dZ7cusFNY3GUA37PHS+NFY0O7I+TZpurfEyBzQ/8lX
`protect END_PROTECTED
