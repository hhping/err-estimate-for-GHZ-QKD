`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3x9grzEMFFpJe/gRJLNDTl2JmQMTB07ES5o2nakr5fqxcAdpMmPS77MajT7voMAS
EiBYb5DdQOQ5qWfjmyWlO2476uIbuF+TQbbyetDhIQQ+AfOH9lFCLE2KoYzK040h
ukAiMN/A4++llZt6Nr9iTW8Yjc/3+6eu8XNvhYByIfl1evFjJBQ/5cGhopNQQCUO
rxWktUWMISN2mr0XJDLIvWT3ZJDQ1P5PaSMcwMtP5k4StLfPe6NfHqMycBp1LVAG
qWOZnJGPk2gLDxJPPhkck6ZfgYTA2RAXctupR5KNmbLjY/qsAVAvzww1arHwuHAy
XzzCDp5eO3BnPOc0UNbKCFUmatw3SvGqGWrpz5jD86K4rupPPvKXrV4oHJJHVG6W
oSKVW10ssWhrhkGmJWdIt2THNWdtBQAw0RePrJYteDVZaokCKewswJcaB2PfaMZC
6x7LyzlNr3crSxSRxmUXanuNzEq0g+WRp8n5xlnKGrwv6l3jPSEB8Bzu/VhjlCr6
mh+/66QZTHNN4eVwsvyogodCqHyJTXRGJZL87bBT1Pyp6wk1U20Vd8KNyT6vQ5Kv
dVzV8WXP9e5HokdFym++YGxQE6jsd3YnYYiKxD5sBS0JQt8/g/KGbcTynwczWTr3
ESqgf/ereWK7n1TTeipDORGAE4Q7h33ARlWmLJOpU8gnvnfO9+uc0nFClqlrrNf8
ViTOwLtj2Y3SueC/YcC7FzryUOrXM3OW3F4ElCRiU7KW8duBpHIw9ZYtt9HPo8oY
ObjuwhK1ysP/5d0f6jks9YRLLj+Vkc/7Lj/CzWiO42JWvzY4THv9shGSf93jlLl3
EUBeqBUO1UKyeLKdX9o3CY5PjH/RagaHxH4BlKH6XOKoTnC5o2SQAC6ZsIBCxayL
4Wm1QsHzjwSo3NxHdORVBGMJOEu6wl/da53SsMWz+jhh2ATPg9RgN5kYsfWTn5Fu
QjDMnQ/pBjfAWYOt1T7+eOoh9R3qsdndN3tg5rX+F2lBF2iFv12FZTHGmcVyrWYX
TylWcRIEL4Kk5LsONY5CxXj5ifjLJbl6a2FDi1vlmgR6XQTwdRC2epq8FauVyQwj
0lM0Cm5bM17OtSxvotwsDp8DocK16MAt9mnpi+DKU7CyqxV8ltcpWiwWUuf3dVcm
Rphtf8ULa7/f7wglTlUeOwCYTt08nGq4aduoTYRoNNuuISOfKitqFao5fPKBRwps
xF38bPJNKRmkRBvnVllbmDIgxv8AL040Yu5yMEJoJAjSfPTGmGwMHGTudQzhdy9v
DmWUbDvuXxLc8xLRAZ7mqavuHknEHZfH5V9Mu5zFx+LR8pidC/CIgL1W10IoZrGo
biAINBSC9fuqlFXFq2MInwpj6SUKZuM+50uvQ/V5HkEnQZHrYtJA1d9QM+VfCksm
d0Bd3glDm81oHCe5PDr4mvg1fxtm0M+Ku6Fiy70qOYwH1csm/mZf7Ku+6OHcvLjm
4ZIReHbWOiG41Icz1+70rdX/TRjwB9ZEBLgU74cox6/xa+vBDYZYgdT6/1YIqfTO
zdStMNQXxH3f1PREpggAblPKbZ5M3TKtlyix2wt4C66J9rAoOGnm+860DNgiE1rD
PX6LIroKyp5O3hIGhqX1DEFgAMFoVWuVuARyiiUtEpy02bo19TeKJAuiM0ovNbFZ
lkFzA36UUiScXYmo7KFP/RVSSVb91gnjR//IrxhcOUf2t3JHo8wo+NUCCFvflity
rTU2OE9LI6AmxsEAbAjiQ/ZM3qGQd8ZKH3hty6PG9KRd3vP2vtq6fkzkcTYZeNLD
i/0ofRn6RqRhBWDpBfwjU9LvDgWw6quRw4WhA1/Xf5XpXp7zP7iQC8eqKgnTzxj4
B7vmkO+nms1T4T336WuE+JAko+ttM7erV3Uspi9FVSZNy33EqpXa9U/1RZXdizvU
5rM0GQAuikSLfwqHMFa2DIIH0PEXtaU/rWT6k903ukvW/vBdXJPcJwFjMZJygEyo
BeclVr+qlq/FdR34+dy/a2CS3iUpWR5EDriSN51UjmRIGAD72RZIT0058daJS0YN
uJRFIDZT7F0enyznuOILfZ0PpCL0kThouYl+8zU0fxhTsGlMAeOpwU2zkUfFsg1G
DZLn1+UbjOWMlR1fGO25z6zisvGtygR+O/AP57L18wtHxZ1P8J/mlt22DxU97EQ3
hS6Wu/aN+T4ofoppp+x0FH71uPaHQ6QvtzWpjMvM+nMu4qXYU1OUNI2w7feghXdm
BH/cvyrwFXCtygRf21CP2qPgzvSg//+vveIzUmQJUF4woNeZixXCbRtHxdD+dBjJ
95Xpzs8EoJSVcckIfB2xZwXw44CBGvOm+8q11BgcQ0Opub862lm05USCgoD3v5+f
QpsaVgpze1D12xsgI0/gXeQugOS4hKhEl6osmfjwjKwFpXQA4IbvB6H/123g+Rdg
e4tg8CnpwFw4xuDTMlaKQOEAiBdYMsYxq6s1iG2EbEZ73K7O0DREk4FJmfU1R8tc
96DYXPHQHF/k88WOorqfjnn8DAz8jbvJk4VNe6pSznC0ZQwOJesPs4FKgnVvYqFs
HfRSWW4SNb8UiybEryeyhsVlSXZ6sdvaYofmRCeEalCoY+11iILDgQyKygtQbhqK
T/73cP84RiVuVhDgHPjoqSlIzbtczJp/MWQNu98pZ9EWG6J3NuPpqGb7EmV1iF5s
M23SYKiEXxae9g33iX119Q5gqlr0T5h0aLU5gwOWM4khd/RNIGowGM0H9aF1gJZX
5amPPe2sWNn8SZsHZykvhIGOLpIrxakS0plGEsUDdjSCv4rPnT+sV3XjS5NtYRsP
yfHDHpjjd7xKkwCNF+c3w0gif40VcOLpBIEiMhRQLfDLzsQrwYrXhZOWmzK7G9CV
+tD6vFqbYrd42BHnvodGttmGFbY2dj1kY8SR3bmeyQs=
`protect END_PROTECTED
