`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLyJbmUbbdKvKnKdDpzhnWVquCHBPpk7ApJeHihfwJLnkKZvsUJscB14gSdkkBbW
se0qZvXeimO9keqX6OMfJlLKCM+FqmOETPVH9x5bxLynHgXYYp94tn++pNKWYCn1
GpLaHXVcFmdZLkGjZuIO9kib4kefV9XHJ7IXKuBuG/BMSmZpfCGe1vyU2PGWcxFq
CUTAJ+mUae/JzZdejmlTanG5182tA1hK3MD3Zc2wZJe0b6omJzHjnvGOF5Ed4SQa
rmMOB9LZ7UIHF4Wit4nCN7/XiOwuwcqAvlY7ROlLlOQcdoHGmJNDUn1QPYsH+dLd
4Dmk8IcGk29IsCZ66VBhUVelZ09RP0mBProGqItMCRKJQpOx2dQOkBUotFNW+noa
rQa1IwFriKD5+jGu/3Q2Qr+XFR9ClalCl+rrmlai0ygskyTMkH5oKEY9T2aBHksW
YvdwFSs3aHHwH2m9SdO/OMsiNK86XeK7Y+l0euddyDJtocmFCYWn/tW4oc4a7NkP
SbAsnfLouEaKJBwe2hi3EMkLFYz5wLafkeY8rdNgIyG4wHFQHtEqdoLbBePpKLyT
VYtkkxIr2oG1VnYTCbxifX6G0TiDvkATDhjj14AK80zJ+aIbbzlbTBUBR00UajBL
dnvaLiA+iZkoRfCG0FdU8wH47BXTsC62h6/u7o3FhjyQtSfjhELBDragVm3w5Ix/
jA2K0fSaFWegjH/WSRdFQug2wWXM3x6qtz3mJQymc0ALLtMEWqfTxqODdGP2rVmX
YWQY0bmO+wvfk+ZC+PBilLBmddpEhbqWkYoqFCLQ5e4E13mP7Koy9OWXFHLYXZoc
BBTUKSu8m/c4Yg8jfuJxu8CvR33J1NZUilkBxrr2rXUCq4Cvbo4B/eA5v7mQgt0p
EpAKKPMuNyMCQ8fNpK+Mo8mlHGsJm6jXfDB+FVYFPx+qtDdrre79eFs6gU1YIDOh
myS7iwjV0fvHgMSA3Eg2JQ0wVezyn0Jc9JFDrad3c9Ws5aZ5h2w+pi7/bE3vB4+o
2C3hseIA2uLTAT5Of3NtcKPV7QdegFMSq+//iODx3VUreWMwJeAS3CembdTUcWup
o0ae/DaLRKzQEsPZBU7JHocNXFtt6BYTJI2ChQNKODGkss7GeDjPQIC+7g/2k7vD
Mvx9AjK0ReY0MBcmCjL7xja5Zn4WaH0j+PKvB+DyIGSW5yFUCYDp0kZBnOSxZN7X
PyuMIofxjNcFf/58z4GWfR1ZevpO2xAL8Vbgbc3lkn/o/pqCFTxbo8XHSQsxB40b
NrOGzxBy51O2MEZbwDCQfaFTzfSciJU1bypcaswg7jA7tHJxf/32vJILI/nx/PQP
+GFqFGs6uBF00hjPLlZ3YYl1FgTy88DQynEt4O/Cw4/PNnOa9hfSgovKpHC4ko7H
/FN2P+DnxEBiZxvU4juJ6I8Su8i7ZwDQ0qejuknaSksqCG8HTmdoZ5e47zzFyzz7
vkEDZilk+nb5zz02lUARlwe+DhMhl+SXRgsycg+Be467L/EFrQm2RsVDLndV+8C+
r0DZipK1EataBi8NruQ59tutN1t725mMiVRxNx2+4GRWv69MKVrMIIIDVT0Wcr1v
UitJi/eS/0OcG1IhHO+UGPqBk+lDophmaEcp5/483amv4YWr6rAVpDBLc3s8cg7y
0MMv3ecV6pyLNEI/ZvuFFDQC6qchdSe1pifPGlOuiqbz4e5bEcqThtjLMWhzxncc
/bHBlp5juE4XxkLJkA9Zlfv22M7xDWpwEHB7LAW3z+DCFVy7qyMqbPE+ztEO3BS4
EAI4PMHM5cxtJHAXzb7CQmmwypb0KDozuVEXKZ4WFg2Qs/+lOz2EAYkGBiHOkIvC
oNuKNttfB2s9ogDf3VO9lnuMpTL4+9GHE1gG6XjrJ+AH4W/F/sCrr1p6HsgrI1xN
fdhCOFHCxdRL2SWAAlJWjCeJh35yBZNLjeEOVtFITWLorOQV6o9OFBoeZt9915u1
YSZ1RsSckIMHQy/4NUWpMBZpqg+I3TLwA4pHYkxcyf6fZWPwCduwTVRg38eqz8Z8
Bh1qIhCG8n6RIk4dQ1AgGT4pfcho4o+S5C6Dan88C4lb8naU7ZVQjTPaDb6ZgJD6
Yfp11zoK1cLOnIr0cJl8QcCT2QCz2ciW/PbaHaKJHEwvruFtwnbl0adDRcvNAvjQ
XkQ30mQHRivuICGIRM3nVzOLWGfPQRD8xnnzDiIXi0NrCaXXwSZUT02VZ+iPKo6m
y/WRaiZlmhc40FcXNJh19/koEsYCSMCrZ6FlMSS6gGNakgmVnQeBBZsMAP+enIoA
+rA4KNKd87zCPSeoUefCaJfb7vGE5wyLKLjCz4dUANqSzI5Sc6bJKLxGoBjhbJLi
1L8cnS7QaxUr2SdHB+Ml++GsAtjhBbw4fftwYVDw2qR3Kywr3swRa6MH0FBwTJ8V
qBUr1YEDAb0dhHakcbbO7qqBiaBQeDS1G6cKlqj4oK8S0CyQC2rZu0b1GPBjncWh
vE0ivPfhhCGOhLUVcxz8wQb9KnM6It0ZMWrOHWKsw0w07ZeT9LYqv7Mj8/A6zQYg
YEhlzGate8U0jIojMTMBg6BjYgoi6WU4BAoVQQ8v3HPxMu/z81Wo8d8W7OA2tYWq
GBIMmEhqdUqlm0ZgY95sSEuBZMwgxEp9vvcwoS694W7aOZVjzfhZu2ZXX1KZ+GD7
QzcMqIM8nQod4JTjw2TsdjyH6jJG+zNvvEJ/MCOmkMmtgfGnIZ0vR9uTweFBLko8
H4ggaJDxfQM6qZBlZJafAVa+Ed+Sx7TICiTcZaZvefdDMYpMiOgM/2GBQMkRKuvb
N6Qw/kJTHaeWV9IfNlCnfTygwj78QsORz4uz4eb3iSI=
`protect END_PROTECTED
