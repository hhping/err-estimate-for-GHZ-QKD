`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cmwIpxwy2O7kz2vuYeC3Q3MrZfdXEklQPhekhRyqPj1y713iWeV3dbTJDsFmIF4o
sPxxPDKlyESQUVSHNSCw8ooru+vibRzZhnyscH5I6AhPh5xMSuzml9uBefFsVVmY
oX7XQQ/MXj4yPvQOwO7GF8Xv6XXXP/DXQCgMU/iAc9ZpvrFJXxpdUfwQ9rAh7l1R
WOFquRom+MSjcIRUDkhWMfgA+ntGcMtBF6k97DQjV0B9HPeEhIFuGPT8wTgylTAh
eMQ1LyNks5y04sjavaHm1OG3iV5+xUlEJE6iW6Ti2+rLfqti7A9Hcs2CJwcvMgsO
acVtRgSpHgK4LIAxEvSAC+PyDSaMgMeLIDLbXJpw4+8WG+Zdm8+j1HXrlQps+Ekv
61fopWicTpOu42C3Ty3xZFMbCf6W9tjpAtCHsFFOrkAP2Mhvqa9nQf+Bh4J7mlAJ
owTpTbDg0DU7V+V4vcBpMeTto7whvbcjNEh/ApH59x9LWoguo/8hvStA1VBVYkKm
QmsaDEFtXLUq9x74HoCF/qRNPXAg5AER7djw9c2zuNJMhlRLVwFUnfRGsiltxd4a
YDEmBn/d6aGyGR14nT0AQAvc8IAwUccVHqIS640sbsM5YLaOseAmvZTs8tKX8o+S
TvBx++ePubZx7Cv/nwtwcNgAyhs9m+JOjKXx3/lldX9iRxqsjhmi7Eupuugcv58b
XHceR3fyQTksv8AMq1QH9dr76VQ51SAu28bkbob6ne0lDdNC9KH7uZyyiauphhkf
wIVB+4W9IOXSu6yma/jOGIDAmkJ1fzN5HZ3w/pbMR/JpErZsSuBmWzQxCpbVgIwe
vligXBi5EtPendjCL3KvXHCEX0Unl8O7QLab8DTbHvl2sHT4Uqn3XjjgZC96bX1K
pE3NtK/K4b/yHC3aeql/hQRfAh+7Mnn4FRRwmgfi9tYuiMIKLx0IxqJgKTQ93x5N
j3x/xieKpmrn3D47o5ZRpaGfZoWukhTtvCGYb7o0leTWtZ1IusIpEqZ9QCoK0c37
vMJrcERLJlY3BjvEchBFkgJikub0ES4CGIrTAKN5z+yBJ2A9vPRkI+QI7Ca2JRHb
xubxKz5qCy1sA22wtDYkxkf0JkvQxHoSIsgdprfZTlCmlz7gkKEC5bhmo0ug0X0B
VKirfmUsl8LNDNvkbQvSfZEYWb5mjTbSwMKzBgpqp42BKo62kGXMXNgo39iP+tvS
JyiX7mivuszhHBklBhU5uAp/tvgNdgeIulgHWrmJUGTmZVGAvfRMLJ+l3C70OiAq
fLr7tsTC9HGB3YRWbmoSpsWrhZVt4991tAcRkqcg14PQ49yZ4EVqlvTset+KioaM
`protect END_PROTECTED
