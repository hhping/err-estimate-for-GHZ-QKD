`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuQsFmJq6ZQPTBEsk+D+bCPaM2ZfNlua8l7oscpYKN6U+nxYy4lYT5X/6Gx6FM6g
vlQWDuTCcToJyVJgaMNdyQqPWdefBw6Uoz9yIuvgvg2FaR9N+7J8g7t00I9i5/o+
GszPDcCXbMaKMjnWwNr4BIu7u1YKTPaz0XUbo3N514Sj0Ye5KS6oXwXWK75RMopT
+fqc1QdVShTV8vIcpo/ptm9BwGAcCoufAhRhAzrf8ep6AeE3dGrD7sV75pRUcj6H
VV3NlB4j+YRgu99imUfUoo8aMrR8f4+ulmpxpCuBpBNHnF3si8eO06itkfJya7PV
8cOYoklLxuwUQx27t3fPYB9VpQSKXnMxrbcVuc+cK22G08upBwFcE3YDfhcvvKwO
TNQdmc6uxNH2ZpBCi/iPEkB687Vmp3dfFqrxPBOVmCLiFDCfJBdP9QM1YQl8EW1W
ZW6b64tWxRwd5WmGz2sb9L7TMWcvwc6VQBq+Jtrbi/CVhFhgUAH+LY2eTcvsNDSo
ScySx4XxvqcvAYwog7R3rO5BHSXlg+zHzT/crw2LZw/IXTBVzo29ZK87La5S1n1M
RugB3JpmL/eknVjqWaL80MdUQOltjtRuwN1pMPHT/nt40U1rBY7WjN8TRGWpmg5Y
j/CivT696yIgNy7qqAq3J3N3f/pYByyHfzJRCQkLSJc2jrrf+M47IGEviWiLZ+/r
R/akUzdrC39viItAL+KKDh568ZE+NnY5+xIA9l7CdpRlJYTIitSuj9ZeVH4VoymV
TlOv4ifDdMvEAWlcrtBgdi4p5jO+/h3kSxBnkAsDszVO5j1TCKCQ0bpE13V5EXe+
xVUtO7J4Nl9lssVNJD/QGlfmTOWGtnQNI/kjk+0C5s5oxRauj6l9uQ7NKIlzE0RM
oUrxb3kg3yODyzYa7U8Yz3A8UikhBnQ7Yz2DfRdYhha+I3i89lVUOluheyA1SCPm
mcnA0rHT9f+YWC0VDVQ1A5yY34bQtwufrw+zcv2Gt38SkWpU6bQng+67jI8uUWTi
1izeK3+qNlZC9SQzDbls1TpY1zMcENap/NDOmw28Eqim07MOdlOHxDB+1dxSyJCJ
Cv+FzxHnsD0MRVsN7IAY4wpco2QaYIO29M8v25P95RTrRJEGViLwsBPWPWJronN3
/wMYsMvlraoYnean5TI7nAcDDW94Fnw9vXvybQFINGLFuJNy9l38I5CqounXaaY1
fR3yFYfohDigrYgMaPStR4F8cTtfF0WMGx3AaSZ6aGDA9g8fnLUzS4ZCb7mUas0L
U0rk2jfHmtebE++8RK3b4gwDIW0ckkzLcN3knccrViHAuGlD0VDO/ChEUYXJ2u6H
BgbUj8zArPUAVaEeAI3IkMyOlaehFRIutmqi+SW9voOTeQBgqB0qRr7bum1s60WS
2Qo1rY9jGiXDFCrMUkTEtuxWmjwJJsGRD98wjYylagE89FG3wtvSd+YjAxqI7uWT
4/nU6cdjuAjUO6T1F+ZQJO92ANXt5PKHA1qGROPR3vgU/ECfHXmBTt5BmVykRMTS
K8t6gCr6gGpvSSp6HgP977ykh1alfrNo3Yrrfzyl97rXDuw4bei1UWelXRQNcBDm
mbaBMq2gEHizJHtaJe88yzhRMVnSfli0UExrMMnOsrKT7BV8fMt4PVcJ8x1FkSpM
tdUpjDtorltiELa2JFw9TdyHhjc+LHRGz30qp3959uLZRVZ+RqHmikeIucGWoCY5
7bNVrQt5eU35urcYQWUrOluPjDOphFjhHqO2Jlcn7eCCekdFEcEWz9FKBj/bKUV1
IgMkj3kbK48jYIM7J2bcaaxFVxNBWTYp6Sl/Eej1TQjbPyzvCZztUgt9nQX78JP5
RcBk23HEJ2Ez/VT8CuV7K00NzlcaZwttd1H33E8yOh2qRtXJUe/Mho1/MHEuGDo1
Imm62Ok/C0Bf302xEahSXSb8DN8wFxgUm1DcFMnXGkjCbErtM2nXNz7oouDQVlHh
vZNCWewda87kh7VMSbZaQGpER9WIvg1Bgg+BBcBtTgdgIuSSDaTDA7oT53l85BUo
mcuYjQsZcGw9RLEkUOFVTV7nIkC+F5Pqx/YacN8LD4cahTzErVqE2szDLf0XDTro
RsucsTwnS9gpwMfZaW06KyuRsKBrG0vNfiBz7NN4HpvtE3jGhSB00HDpKX+QgO/k
n1dV4pp/ZrNIdo82ZFXvbAowAHLy/Ud6janjSlCkYOq/BZNxLIL6uqo/j7ghGC2h
6Q9UNAYQR4D95QMGYGYmbACxIFoopfsO2fXijmjrFx/Cmljx38AUt4oQZW/Q3D+S
05AYghNnRf/KQk37n4l28aknmtGtOFqoWT3TfP2LjY4RyATiwal6bL0R/LOnF+kY
02Pn3ipCiD5iW7r6kLA5l+gAg87h7jSWXy5IzHsGzeA8FSLnFJwwOve8RPi8PjgE
htWinzlMcy06acpJeSnN1YRlyFiuPcCD4dbmE+0X5shLfKKJTYFZHuP42E7if7wA
3xopAiYu30l1sB1DxJlGx70MQC6qM+zZuRA11WF13DdHuJCqYQJMN8XSH7iuxctI
k38dUzQU42kqgDNrv4cKv1fdOIwpcqmxrci5mvvuiIyQ+4+9C3vNGnheJ4hUmN8l
qnYOTM9tvQ7lL+AwqDgTvG3piezqm2fny1HKF0I7Z/LzHCz9ppMGgBljVqEyihWb
ZKGPpUpA0qzUCqLFWKKJFvYzMfSGCfhWoCiB05Awhad1e13ow0FOiV3khiwVJvqh
ybn56aP8gqz3d3gFsZViCEPHJ5gg356U0pHNOF1O3ZcboGMDPELrycXP32jZK9HT
0F34xN0Lngo8XAIsY+VBFXj5AejcfGD9VLNYaQwMS8EJO2xIhvU6r9+5ZNo1WmuG
LhFBDWfo138BPejQQgwXT3jM5vMGClddqAnm5QHPsfIFAiRrgjc0LVIvEi+syVv2
6ps+skhvW9pMXMfjhPonpuO0iKDNubaLZ2DqUzDh/qQflSqqYohOcyFHw8Tll4jM
8bDf0eSp20otAt+8MHnBHHrD+fkQpnMXi856bPxvfUpHNoCG1M3Vhn7pFy7THXsg
yuA2Tx4bSYfmeSM7+HIRT1IdyYxZu9QuXxXIpTLk89JffyQpJE436/lHs995umlQ
OelT5efx6DwaEtV20gThYzRYLcYGB3wz1yZ4xc4NK3gJr6LzpytWz1jiD+R7pwj3
1KWU0gxZ524MV8TEBzKE0wjNzxlpl5IPLSL990/idk9LLRW0gtB4DxHLZILjG4jP
Lz42164KewlNovewcBAd95UbKyB0mNZpCObtvUL3nwlcSKNgKEM+gUuLU/904vQW
A60RXvpEqYkS9xZIV80sCIyRh9kh7STmbg64ZH32AKllRm/tZRjJGZIG0dHYUulh
hcHMOxS69ZzrziOyskWklK9UIMj79+Mo3+lT/Tk17C+dseGoKHOE2srg6CJ5cyIM
edF2nfnRtxLrMRNtvspibgunac+9Q5EXLsAbICauP7K2Vp4A0H9v9vJVrnohjJZm
xjkZ3zJsOEWRpNZZc/sU3pLErmT/blj9d4RclLI+1VppV9FVztsprdZymyPACeVP
OTapTJ/5Bz7PhwkmeH7iHcTtK4CbPnh21jTMC2/DxqeQIB+Jy4dFKcjyldJuOqmZ
Xfc7G7SOG+cdWrWsjn5nBnkhxLxJPLmmF+srrx0Jshn6q2J5VYZAEbeMfbIA5QUl
X4UAyw8j9DFUvGwd5pDQ61GNEyB+4tbGWYFupm5tD4Zxhi12mZgxHPduFMtYOjwY
vmc26fgHffjR/yK5HLtR0XSVIKc+CeW04+MuuqBBeIdt3G9RPnPPzwxXxktuW1Ga
el0+cZxSV+q2JbjxQyFz5w74k/Zmd8EUfXE/ZnSnK0WP4+9/tNhqFZAnw6L1MSIj
1DZRsi/LeBXKsqqa4/Trhi72bN27iUOfIzLF6HfMuJ+czBa4tvEL1e/DpBCxhrSc
TrRm5KEHAZkl13I5Hd7cAB/COMHLDRHRTer+BDHGa7jnoUTciHPIk3kmUnLsv74p
i1Y4ZsyWznlghTYtX8J1CNFwoS8NLoYRP5Q4YHGDCuOlwd+Bhzq8+oYG0rriXdrP
BX6R0MLITL2/2nxgjXBdfR1oLFxMOCUdOPpucCiZu2rYZrYAF74oWCun+4IeUJwh
LAioRyjSgXHHzIlM85Yb6VCGPNJxJsSuhblruT+bkpnjYo8BO0C45fKrIIqsvizO
vbAzSb0brRpbkHG07m+OuRvS3SrkDOXGf2sVz99YFvGrjCa45SUacEmXcSUn+0t4
rNzzVYl2wx6Qa33Iokbc6kJJy7+6wzTEa7r3OjBUG9Tv8znl84r2GpZOQVzm6EnD
zRd43yWpBupxTu1OGSTK9e95BdPcjkTaCfzBn7NL7VT9zTBsY+4+6SyW4QtSER9F
MBY3fnfwPBXYqYhITJhVsFgKjzkmW1e8+52CrKghzUINkV7T0NSDhfKqu7Is7+4c
EP/NWFR41ppTvs3FRTEt2ubrGm0ln+uiZ4y80Tc/Jy8RAgXQ2WdFwqlV1W2/N/eq
y9Fr0bOx8+5hpXfwfeN/8NAnYdBSlTtdU55lLR4MEkaGDthTFlPi3ycxXdAmZhgF
C0TPD59XwWsCFnbvPd26axzEbE5di+7I5jtm78Pd1KekG9ubZh9qZP13CkUo1VWa
+CG+fiCJTA4EElQLJzsKPisswxuLTpQ/pS79VKvNlF/D4Q8njS8gSf3qghmvxOhO
3MhN5CDIjnhq3RGGQcrzobiIatBypg3dcxwBUcLw6cu1knn8YrQNLhlTo7ya4+hq
aqG9nC4dWUfYjGmwtT7WAHImNmK/ro7jvhzBwbjZl5FaJMt0Mtkq3SKsnFd6JsqN
2vVOqJvnz6965S1w2ogZVkxopf2y4dxb1Oc5eqM22Dx3jHgcO+OEdPlKMoDcylNZ
cjk/ixS+ADFT8r+fpZAlNVrBHmODLYHAUWiPxRqMAEhMwnubWH/B+NMCpEKdRG/7
2D7g+kiVbSNsWVvkS7AnnzC/dnSPa8WYFQYcb6u9/QoFGl/F2u3CWmzVl5oSbjkt
2lyeHSF3dzYP7eEeD+wbudHsXUyly4e0CHNCXEY2+03EQWCc3wgC7IE/IQe2ya55
pMGuULvu9sGjBLLXu26aBCPBChHysj0Y9WISLKU0jTejIDDJEHX+FZK74BJOuvqo
Q8w1wVgKzOQfcBkre4HbGmHUX8w9RiIREzgM2nR8EsfLOqKepSQ1mJtsPM0dM5QN
07JfI/ZZbX7zc7GavTAGuuweJk8+dEzKRyfX+DZ9Rr/55/WPV4774yiIhimS7I10
Wv64VzUwr0QhzNKE8mwHFG7zx79B/ReWxACs1aWwEnU9s/6mwDREPnOoq4QaH1Id
DH2J9/HBdYB1k9pVdR0r7J3Wq8ZJqzCmLXMbrVScsFB3Lw80UfDsIflP3C8E1lfF
MdUQXEdltEkSE3lguvQsHHPROkAa8FoXQUHMd5fzFxJRuj4c7Dg1smqqdUt2mP4n
6Br3NzMBOjonYnXICgo+KFuTPPgD+cEjbTy9QkEk7VVjLAwXq5KSc295eZP0eEgg
a02Oeh5rL16n01ZTwkPhAmSiBrIsTWeXIR1m3aQXvxsY10RCVE0ZPXwrlKkzzvZc
iTa8H1JqRPnf3q96dJ6CmYvxnL6A5np2AtvP6o3OnK1aAmEJO6I4NZRGYsIazf2y
93dGxJAyY0C4vynBuTgOji0vEZ76WtcBOJ677JkPqJuVikXo94x7hNXnGboaSq2h
yBKjXovWBxkjogH7SAMTvzLXIuPRCTI/862+yWrSIaeecuEuKuC4/VXyBPQHe28z
AINQyK6YcT+ujbBaGDwQrS9Ak8u59GBgwLMMQo5im/1et7KQ3LvwqJ1QoON75gGa
8PzvhlXMBTb7SKBB7ETnj+QUhOjnj7Up0n2hipJGc9BY33YGEwAr9iMV4B9m1uSm
lTTET7+ie7xoYrqQ/1uHCQ9AEovNci3uKu5tfYbzLgytgqZE54aA0iyYZscH9F8B
aWWQFlXFsb2Dr7VZaDCxcJixsUO+BwVmBUWQgbOAyJgM0a1faXTHzdktjcvvQx3D
/Veuhsr3S1UQ5rwQkfvWusAy0GQBMnUE2ACGvVzlTJJN6HoocUkt/NXxRQEKFSXO
m2erqlDcegHoetta0sICs9IwuvWcBvp+ecYC8eQtgHD1gMdhNJZ03tN2JhpZks3c
6VwYRGtzFxFo7MDDebJrNQRhpCh81hIujwleau/K2BiFAoB9/GNJXlmgQsC9yK/Q
eUqplsGIZ+4elPRlsdu6gGCVpuAkHBR1dPPKa7AkBH+C4Vty53pXeLX5jhHOt80d
ICyrU297oeSJWhp91wUD3I+Oqp2C4GrFlssGNlxW3xtMtkpLobMaL4EDat8xUqqy
xGBcZ/w4bOEJgdH4kj6fUAKKfy8hQ4Qzs0sXy2jQzi6n0wxN3UaXxizqOg+z+xPg
kaTT3Isvu+qIsYVAdyjSOfJVcrzcJnxd4eN+5gP+CEEaIeHhQWEHYTDlXfAHjl/0
Uvd7KgUFGsRv8XaJZhS75W2DcYzP9hfSbz6tFLonWzzbf2hS3yG0OVfV1cSPT89b
CnWY7CtUVw4WKEBOJBg7mLA5IoGWge66G/cIdY+jxGr9p80t12Z74oZ0SLOIcRaP
MgjBMKw0mZz2YtY79yKRXGz7YgFTxpycJbSZjuyvu23+TQyCbkYhrpwkVbblUV9g
/60taBXGpd+GGXN46y8Umaqv4I6NQzWzr1S2baFkOKuWzj9VpP6XUtDLNMZOeRGk
ExYmAS5a+jnVEhbFjg5QX6LKApvJWFhKKKXSRbp083KFgNMcfJnlk4i57TsUouF9
uRfNlWlmd3hKh+8OS+EWk4/txDaHddxTtxLfuJBXWJAsebl+gYJgKXJ/RcwfO7hs
1h8KKlsZHYDfHKG6MqpiPYL8MR8dIaj6GSEUWFmRPsQigCmf/HVaBwKr0X2DFqe/
3vlxafrnNaX+xm3ThbWD3FAWwqu+vjseMgn5zsZzrfl+TUcZ/Xdkn3WbQ2Ozj2lu
lMZFnVLyZehiZIcPMgZSrz7ynYzkJ8XNB8uSPB8ryDySYfxY+Iz2PmbgsTIXeKQV
6sdTkxZKyeuJMdX+a0f/wp5AJl65KCHkFCJXXGfQDE9JqdVfQXFJbSvYf2RUWcMN
0xlp7iKIT46oS51Hq2GHobJr9zUQzHO6AKsd+YzgJ2sTGJwoX+euCwPMxd0dedXT
gFNhQ5wM6/irOb+tvXV0Xx+E1whsaGurFm2QzDxWLd8vwe03WCKqbtYobC3Yr/ET
Uq2u6Hob448AXjspACpGXIZ8GwLUNHTRqxHS67lVtKFc6wb6aRub8J9fVm6BKd+f
I5cmFWFKzAoQwQNmV9MYq+92XMXCs5vTS1MSsCFkTv0YzTLCLpyELqECYPZnOn3O
3dUsEkTXQHL17jGW/xAPTlNx76Icwr6l3VWUIOt4zpjlae8tG6vXViM3vAxZAdbW
lgrbxPv/4kW8apWa1wrnJMYHCU2X5vulu4mA2RkXMJxrq0SBfEOV1m+8K51mYXhT
mF7XOrWqbJYRhoYcKJY/259Y1liZjhxoUZrGx8yGlp7JN1y3/E1vt71faKPpLhib
oRUXbDQc1h0ke89kKP8fMpPGAJ9XSX2fGX4JuN3U9hoEDcOsnUDLur9nWGezG+BS
tDyGnWLhFdBRcE94KUt66t1aUMqpC/QmaUJgX8SR/V5PmJ0hoUB9OQk0N4XH34lc
sinnXRqd+RHxXh6xCa4cpi53FYBxgcjBhU1A/dxFh0UsAnooDiGhROcDiVncMrBE
fYTm31O9gB/83PdjfWGgdKZmndMxg0S7e6GbEyCyv73GBbvfD4VDZQZ/3XCHbr6b
F3HGAbkP2/ZO90FdbomgiNCpbUnCqEkQ+dLwTCw/azHJxI0RIXKeMMoNKOwpd+oE
oMAtQ/89YyC4fRufj+Ozx0g65Xae0GEn4VlzmsgFT+cil8irOU8CE+Xmuh9hJbFW
A9vcwZ5InqHLzvyL425RrVg45WwFsVptd0cLT33hc4mj3vXnAKuOKTK316ZfoFhJ
RJ7TdGKf8h8SxfBNSxBdBqLIx+z8Y2O6IBda87V1AK3MUnLy0cpUTm2q0QZ7XlMU
T6yKgylbjK6g13xwCLL5Fr18FVm29LdW+yC0+ojOKRAbOJKBZkG+sD5wpmE4XLt3
GzvLW+m5ZvISfpfae6itbDGw1yZa2IiT0UwBFRgKo6hHV6NTONTF8+ngzI+C7PoE
blEqCR/38+A+olgNElM9ii5/Y4et7p5wVZXrAak9gg3TG1tUgt96oiv7XbJm9age
cWRkbH4Rn6nDr3MGGUWlYknELW4S5bg1UtzijrmGUo3mwJUm5XRGKcfYL22pAwLY
MBtJsQOZrQThIZ4XqL7U5NuKki4nyeGEnfvE6XidJOb0Gn6OJS8kjsgFvqOqjuN9
aRcXYjnOMMsHaNqChgPbs8DA5zZ0Z4U/Fz72RZXiWC3FAyqz4Wqru5pfESaabCvY
03oHp38ZlGVemF05cbEbEItISXwyY4H5eNQmWaRg0CQAaoEDaD+cUDfDXRvbZam6
`protect END_PROTECTED
