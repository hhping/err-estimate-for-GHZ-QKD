`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ThodUDyr8rwS+QCiSZifXmY88nCTuQ/OxkLUPwi55RlEhjok6uEt9we2/QVj6Sq
O/YnztbpDwyHueoaUkQFij9KB1U03r53UHlOx+B5Pd0mfdi81et+9aSfq+3xEJXo
Vx0eIIAxbxBZem/9olIZX2QRJvx698HzJjch8ueHUAvWR7BJn9J3hCULMK6oz9D2
PjfoLZCZsgtTzFP7VcYam4uo/9i1cnh9mzkArkt33H4fuNir1I9fiTewVI6R984p
zuvhOa72kzZj5SSZhfig/lshFL4enZ1tkmS1tmWPH+pWLal8ej3+ulBig4J/iToq
m93P8NXuhFeveBlhVXd1624x1Y7WtuX6H6vk+yFtddSBN4pzl+XOr8g5vQdNWeCa
27Bfnjm9i3UPZqThBsBNyBvEnnL5griyjEpaniGyjdvWOSB/Tmq4qvfuYSq/9aTA
8OZNE5bPP4QVuuSxycZulO9gyrXR8RA/Bd77rRLa6l52N5Q03J3hW0C6lD8zXMBK
ofBJd7U/Ewmky+a5WGkQGPN39kuybR3E7ITsjsAJlWw1CJEssJ4V+XZOo1WG8g+C
rolIeWBo0sfwaq/0L7OwZ2Zhai9AZImCk6L7Y/SpiQlr4SsYCNFp8fCM+cx52dOK
qShtkP4hohIsB3yzzPKU8moAz2xT/7KSRRWSPsI1iwEUiOvMhOAg2cT54/fbm1kw
6EhBVU5ft7OE/w5egNPGBdmdtgtcgdYvKQfNUMrdZvKeXcxghaqh6SPgVjejpAqB
i2/WwUfxmqhb+QchJyKraw+Lpnga8711folJWt59MxP5yk6WzFCURkMyBhTkmIJz
d4yCPhxGl/2xkMThPyvlTMlw3yom1+sNOupivHJn1CM=
`protect END_PROTECTED
