`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLpgYWUBVpk90VUvLGK5oU6Af8Lgyf8OpbPQMh0R/2wKv53Jxpt3RkW7SmZ0PFU1
QCE9P5v/Vuh+vk+bgTy50FlrL5zdnEo24r3bjABC8OTPgHAVREevt8XB9NMHctRG
Vf0WRZexedydblLwBx4R0dDRR7E73z37iGJr0Ho7MT2Oc5hD4WWovJaWM8yFVl1Q
yrlX7/6lQ89gYrd5cLmycOaXbD9AaLwgjJbcnwOhExlVwm+TtMWOSODdyMn8Jpzt
zzrnSEK+72jeIjeE0j6/gOK+LPuvXoF7VpW2cOhZLR0=
`protect END_PROTECTED
