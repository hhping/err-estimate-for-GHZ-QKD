`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1nLsTYW9OC36qhUwsg7K8nPS1fXYKS2T1CwQ4FBxh6KOiEztr8yqxLAcZw7leSa
jZkT+r3Pz2MHN8inFJcA89Uwsthd6ePJwgBSxPjWRvd4JYFt59oZcSREuFqyNhES
eHJt1kaaTQhbX/tbGdlBYObrH9n4MShDv3/XmvjM6PS9HrgLBl4remWkgwNHPAP3
/cw4uZzRE/GgbEgVE1G6IWZICRaOuvILdGQnDjTgi3IT+gmWN0ieSEM0lPpYjo6T
lGI8UNK4afSgVH43pJc+TqoYkKL3BR9/5/bfB95RZ6jkQ6ODF47YyXOudcbvArEy
ZY3gMhC9/u3IRJzXhWfDOz/+46kgjgA5Hu6P9XdzRaZwznvwEUJRVPcoRci/FV/Q
5Nqlh89iuGlj9yUAlYLIWMTeRrDr7qMZpA+qvxvvk81nkH4qOpG+OyBDleyQw/5v
cnS8g9ilFnfaSIqtNN1RTDWFdFSDD1JwVVniBDZ1mYvJTqQEiKfQN7hFw40iv31M
8jucmzQvUklrM68Cu4alihWXjc5j1vvywH8etSZC3nW/D2wMELYoZrNAuKU3mcuh
e2KIZQagcHJXByMZ8qH81prec5uhWIBTW/vhJjSrq40cSCdw4k32MxXsFvgbYg6H
`protect END_PROTECTED
