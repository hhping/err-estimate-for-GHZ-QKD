`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fD6inpKFowU01YEroF74dlgv38MiFF9gn+U0G7JeHvK/1gaFeheoc5gHa1cdlJj3
x2RBzI3Rl5Mq9srQc1cVhGpg5faNrlFnbgExNX94pgs/8RYizHIFu5Cuo+qprNCX
5Sg6Tf63qqUNKf4kWkHtjgbmSkB1GwkhzaXaSwOSb8tCDJCRC+AkF8MvWmin+nLj
luqQcJDbsq8IVaPs5LNZzSUG52qRaatwUDd5+ERES6E6X2v4bVzNL89GG2D/N5Se
jBywQzG32nH9L3T6CAfBA+vFlYfZj9Sco/nCAx2gSftWUKFSLx8GmzImLffymhGv
8x2qC/La5/jIaDlLkUu/JfBT/aKmwjpSkn+ExiXe5te6GiCsVFmDTAbKxlt6zNLJ
H2n1cMu9e0r1e0nkiCVanAlgHgmaY6cUst4+FbcpXT0oi3dvcLUADDZHPuOwjuOZ
XtOVS7hwlZ+uHYIRv+Hoc4u/McgitQdizAbEux0oCirUHn2fTBhTLyKmk2aKXvWs
3xUkWUeWisjzAbqiQLfmutq/w20W/ZgnYt8eVMZxihCYf6YjtOek0Ciu6zaW6jUe
mUKeQgAW0vaB66Vy9PFyw8bo+AUBw+PmNjsWNQVtA3OdjeBYhm8GWxDhXEBYuDjT
5JlCxi+xbBmqOGXoJaP/Fc+RrvBtbsfXX79YXxOnTmALF5LVRt3IvNiP4fePfE+u
XkR4Vvs67YIMZ/SCfvpwuGjGkx2FC1gG9BQsns2OmTHC5ZxrMZHMyL2s9GYg5rRt
+Sa3s1+nKl/a3sa8izCQtJ+1Apaeo1n14kOTUPsuxulpIcYj22fFpbPWyrG96UvQ
5d86lIwH7i/1ImTBmXJZIgKoiI0jBp+pr88soRXOCQeD+bl3hDbLwS+UbNxPni4y
Xywk1gtFQSDbghP5l66jciwvZqEh2+Fy6ealJQjrujXUq6mVpkzrDurLq2rTWhCH
DpS3era9pQl+qtlKBPsWQ2yUMG4Nkq5wGIUeqjExWhvZfjhefez2nTCm+2jO8bxe
6dY7lG8+z3Z8TwF+7LQrO1HdJfCPl2zSCcVDPh8cyIu+hwXNfwJAM9HMZMGD68Xd
Pd1ZSVYMDjSQ0nTVltoq0kVT+2++SddkAgpQBol0x4NEWR7Ms/739w99L1nDMEgP
01IqhsQIBNtnhoYKy+P83qqu9u0sxXTB57g+oMoij3siu+hq/tfFf0kjXh17xwON
9QM1JqHcbWMBv+A8NBpSCFumLF+VwRlkyTJFcwXP6jW71XvJovcQdzwuA+iVHR9n
+dmZTsk55v1Cmw8+zqj6T5+FLleq5Xz1E8/785LmCS0W1sdHLLaE8J3NjzdNvy3R
rdbSGCpv1SCBcW+4w22iyfqPyBoj+i6c3juE26Yk6TDodazeQE/A+sV1hZ00RAIS
rOfZw8X5lffhOojsqDfjZdZRm3IdOwqQs2PQ9bKEF0Dco3saFTRf6XNSKsZXxfyz
Y4F0ZBS1qTz+z55FHxqdAYAD7B7gKJIqTX5j7X4oDdFGkRaBomTJe8prGoYn/jKO
Eh9uSsx8pNQN1KPekIdmpMd5EPSYd8jtY9JEp+XTUQQbz3GG09W1F3ug42orqb3c
14/hdQJ77YBxlbYn/QErUQ==
`protect END_PROTECTED
