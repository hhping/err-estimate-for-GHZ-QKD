`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPSQsl9fvnuaW/tjRTQ15tJEY6ryy1GQBQu1zfWJ3PLsvbOHemvBBkxptZVPKY2P
FNgyTz6wxU0XVSAq8AP0ee5oshhwyjdJg9AuSLy/ZjCI+NuJtT5R8GpIkyojVvfG
ymgfCcapFMqsOFk0Lt0c3+GmZsejDdwyoT82jIZ2yuNQj04FCFmOtrPgfRJ/sjMn
QTUVrfgXHX3YOOqcBrrm31jakoqVTAfvb4UdElU0zs4zpEqirzCCLJBLIk4wBg+G
jSi9IxPmkIODzZJVepTPn79X25Qa9b7t/93nL1Jgk+BJj+vdhJSJhb+Myh0xOzfp
SKdyqTSBYzgh2PGTGnI6cAswT/l7o7Y5sBPTL2rAAqzeIOxI7ntPYI77105aAqC0
PTzkfGSgiowcowGF/Upcu3sX+YpBQ48vq95pASwfvO/eBqCBa8Rh8f9UyLUbgJfB
22BP3iDgkAbTfYY2H1T/oCvyoLOe4Ekx1Z31P9jhvdDncVF3zb2eJJOV3Muvd1l8
lKycBv2rgL47HQhrIWvO8uclSdvIwXKVBvb7HcVJBP2Hj0+qVldA4sOyVlG7iGXM
P25NQS0x5t4C/aFOSS6VOyi+yNTgOdm52aoFczriv0DKPldOY9C7A8DDER9UTF5R
+0P+eVKPlXCyj10gT47avMGYw1YvmV77V+1hpK0aJWBaz1qRqDRru90IwBBexgXy
1gDrXxU1bCIFtG5bfPQBldjk0FJ8OHhRNH2ZbM3SxofEVKM4ZEKsm9SRlLm0jJ65
nPdtrQE9RmNad8sav8lNEYyXpwYztBl3KZ1TUYWv79OXiyvw/y40BsqojniDYaOf
HZJgd7maX24+EP0b6IyWvkI2jMR2IlVd0PQxgEbZ98l7kJHtVYEIzlIcfyn/k48g
3L5Mkx8DZcGjDNFFYfxLOIL6NvbfxuIB3Arxv7b/LX+F+8v+R6f7IFn3K7IYD4Jg
pPEuHD1xmILNdRIGCVsFzxlNIG8KdgS256HVeNRe1o+cD+kKrH5ClTkuJNAybYKX
qdY8IPWJSdq9JZwgADSLBRX0f6rGTDpJuX4K6KDRHog=
`protect END_PROTECTED
