`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2B0tKHaBVD5JA95NH7/19OaqeIFfHXdpll6eXE5CK/VwWMSpo1LGa9D4lNc+q9Q
uqLT75y93z1NWEpzsCM7yRulX8BqQUfmDQf/f/3TPlWshtImvyhDK0Lvxo8QFNNA
+eLaBQr0i17M6Db23JlbHW6hco6+BF8V73l8+xQO/JnKA3LiRaxduHpM+qRgvFkl
PH/PpIffd3WMm7tNAnfooMb61/O4Za1k1NZhekDX3PlIhhKLzEpZuWPGwgA0Od8w
6b8gu6qF/WZlY17Mrg+njpljF932Ia6fqidf2eIOenM016KivDAEZq2zXfnNfl1d
H8XQE9OCiA0VBgTbj0FK5wqhkkK+t45Gy9H9cIrrx5B3oeBKcjXTqhRTtkdTk40t
b2qq22Usgc3iD9CDBh1rrBPQ56eHJXS8KlkBwuoB9sK+TwGa25xuhqpZuHhN8SWa
zUBmgWcPX14gajmN1+zSWmo2CZqoIzpGyZ2K13iJh7MbgcH39jln2fX4csmsRRAN
YRvcbaOcDOPtthQ04j9ajEKA75Zwv1pXXyVaY+om65JbViJ6CVcO848wleT7tS+j
Y7XvvZ8//4m7fIQeuRJEBJhkk/BQ7+E19xFNUMUJAvWpJ9Ttqxx/lgS4PF4fNWO2
ild9E2DKDslwol+he3kVXPU3XsmW103Vu93G+QemrLuXCagWb+byMi1CVo62/m2Z
CkxrCevjELIsPLAb7R7MaubZ4aeBA22hOH8Ad70dtKXdxv30ZoUDY7jkJQAdKwGq
Zr21KGiCNLdcKm+OxRHtEE5dUA5yXJv/O+tuET1ygrUx/jj/NhHF8EmK9BuEeT+a
`protect END_PROTECTED
