`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+fjCVjtSbZ9jth3EbkyBG9nrB3FV0knWGbyyrukM/Xye1xp3gTMGIJQz3vuM7Y9a
bXXzLTd81fDu1eW0PG4tJoFxnlZHp4cK3SY76dA5u0Q+z5VYpUp1m6zVaisU0SQU
KNiB6wYwe39oInmIsQHgGlzUrkmjFTOPQ4Qvus5wfKFB4UBcPYp3AuJU+jvWy6sM
RhfLWH1Pw6POmq343R7vGJAxZXwc4iQac11wYdbCPt9AoAWSenc+R3f7RByAm6YL
cu3AqwoeOjxS7TtcJjsUacZ3efqnseBFm+Qhi981IFpkRdQgXins71v4405KeuEK
/U/ve1AMqyDZHZUkrdDvbojSFunf5mrRqkhaZgVOB2m3/XcDinR7bmFqqA3EhtoR
M9e5Ev//YKeSfyawgcIw7gpgbQPLJNNSk+gR14eJ/dsYTVEU3v7U0gaILwEJn50U
JH/wDlhCIBkzWqJSAbcg6LO4n7xCAXKl2T/xMYIGmsAaafR9LJY4oZHulk81Wwci
OugEHGqRpn5LS2icPivCLMJcvyVgun6kqv5YTfsNAEg76hh5H/3/WyZs9fxwgE+z
/Bofh1Hx7ckTriWnUnv04crIiKTXnNI+DVfSlPae5iZz5Es8S4Rn83wSudwkAgYO
KZBLtsaMPvt4E4VVauGnPF4nG8slYu33a6hUUMalFwBfe2HMQHc9n6yhgQtO++u4
ys4RNfdQLOZUcYE6kLux2IKtPOYObSFpGl2aqJDbkaw/DZbtoosGoDOhz4PWK6t9
fkP2XF43r8+UCTWVD8krklKtKkwpd/bMAsPbR1CSrnUmHaHiIOp5yprG4FFfx13/
MkObNg5EKR/+RVUmwv53bBtGJx7mnIb+a/kK5gIOsboxwLSnurAGXBuZZX3DZNPI
k9DPvAX1KlLddjENoRerrkXDQ2LV0JXBZaPve9QqgdUEqGK0Ta0RdYzLx4sLQlK+
BGiCq2LQzVPr65Q0e3yJEbXE+dkTpd4ilp5E1EyAXasb07Ok/QjpfmiVdoYzIPAv
N/BPYCWMe9IzpOd44T+YTtTtSt8LRcv4HFJxtwARUTCvh7UVWQdpup3YtLWN9nVA
qipVpMsAyzh+n4MuWjNPRFWeJcaY31leZqz+UUTlI5Jhn7yHhV2cdJ8hRVODtHhf
6ffu3fu1k6pN3bTtJRMgBSzppZDaLt/JvMu2qW8HuBP59VK96R4Abdp3XuYuMpRC
HniLIWISKI1QlKR7kqRQjlBDxiITS9X/9cpdtwIorcsJfAeec38CVmNuGXmqxXpA
qNQ3GDTyTdcM8IE9XB7QBrfTgvJJZamYUzwByuPXYt+RFvvPiKAhZ2idE3TJznvz
x270l9DPvbdYanUYdSIOFgstypPnia3kkRdO74U4nYOWboZdtsM/2hXFVmN/WaA7
BVgC9NaV8xQQelWxmpH9cBNgHBQVS02dJSNi68iX7n6QlKM+Shku2ef+j/LNrZ0T
UevFnEp/hzY20ZqttYnY44h794B+x/SepEPn1c3O/fo/gD0ZmicWsLFT4Jt/W2Dr
A8WMID8ekq2G2Et63EnhJ6jgrHNWMF7EeqQPNwRpDT0IZseGC3Xb7NLht0oUypD9
8Mu/Jv2ihGTULvESiN4Ygw==
`protect END_PROTECTED
