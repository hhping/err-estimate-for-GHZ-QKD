`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
463ivzB2CWOSeXnSwWpmf/JAy0xf42RPxYhpYur1h0aG9s1e/LTdANDLx+k612u+
fACc3G+uJo8xn4auFM+PRhFxWM057kW3647350Moaj3scFdJqBVixmaBjsimBgu6
nStzbK02Zc1j96fizcwBYXxw31tnYFZNElZ0qNfuh8W136AlhfRfOUKtkXwmkxcD
YezqttUqZlxj9gfi77WTwOLiGuJdo1jbkKpEXpfXwJWKRSxhB+0Mq+1UGp2IdYUc
QwsleJkrGnlOwxzRQL/XpWePsClXfZB9idxZuFwQJyMejV2MTfhGB//qzSyYdnTo
IdNk/uKNV5oIq/I6Dnq0SeFrOER6ywL7asAp6oh+X3axSv8b5xF0D7Y8p+GGOLp0
FRSL14yTDLLzEPTZDC6aLdC1S/CIv21VwXhyD8y6b3fADQFK8Hh3pm8mz0Gp7hPp
I8KEu2oXFe+088sq+33O3oKy1MTWLfm1bQhPrQlTjSTZvcObL5MJK8E4XpizXpt8
pO08QhQms45O6Fq4MAsRndxqusoWvJuEAEFqYQt33fR1F0YWM4BSIkHLKhUTW5OF
hVELmWVVKPlLNNWnVqDJbVqtz7TjBEDTCJwT3SnG2kvuo1ALeORap9rVoAw9u9KE
+lx98HhygrRCpKT8FnuGAqjwbdZhuhV+h6jIeih4GaFJdrsQtU8qpDZoJ1YgD1Oc
z2ISBVnVegWHxsuJonVepZ4Y9ZgP2uUrfHceMMBZuA38Q92Hmw4OlEhNUOz2tqe3
OaYZsgpByZ7S+5bi6xXSJNJ6cPNk+ZJKsXVYjuPutWo=
`protect END_PROTECTED
