`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Bu40lXQqMlqTOn7TCHnS4LeDgN6lauD2yya7sA6/RlpnYQ27xs2ffbyfeHCC6TJ
k2ql8n4n3MB+/j6qSvtJNJlGknnPE2AkeYpkWtGbNHV4BsUMcVeR7SHKccA/emST
3XWuSqNw2UH6bwH5cGvOXHY9y7+4gQGK3EL0EFmiB+0whLXGiOdCSi+iGSar+AF/
ORzxfC5NQ/drjiRAAn211cBSE8uS8Cgtuy3CRwqZ9ZAS/tlfmT4VJZd2hFVSErrH
To7qYeABnSCBHsgphvYbjNDuBroduJlqZqB4BpdZiMERH4g30bAnyeTpAqLaceX/
OQ87c+u7Zc4FrUQNgZNv5gwBEsGpdW9hKczhHq5hiDFGYVpNRN7GrXKup55Qje5c
P/+8UAUrEbfES+rlVyyVRJnNr81lE1RzAw7oY8XbwoZ9yt+rvaMrzwwoUkXzESik
`protect END_PROTECTED
