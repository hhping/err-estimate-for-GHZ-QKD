`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aa/Q8osm2PQYVJA4yUrYCtHw+bvuHgEPzaCrGovuzICdpaypdGdklRmO+fLxxV4X
Tp4dWvz3qJGTNBegfRvDyN0xrTezk5aa++VlarmjGHCaF4fMTMmN364oAu9upYMI
4dVkCefnGmcIypZ5oRPTSHYxDlCPsiEE6XnNgLHWLty2nmiV67CqZxJNxvMv3So+
gcTldD3PcVZK/zDolDZimYR4eptTwpPiGylnDha0U9N+Qc1HJYNGgs0OTpLeA5OM
j1xTiXxwkMeME1NxQOrFn8aY+OywZbpAKsGYnxUrF3e2qiLglrAt5zXcsBnsjxoP
Ddt9pJWwyvR2HbogDEo+rvOJGRuNKL2iojepzU0253B2z/WklbCbz/m+8t/c4bNf
g6S/trPtiY1b5pvj65U2PMutmLzVLBo2MHenJbj97Hp5FIWnH0yEjkvo48PLJL0K
pefB2OfSVbobRuAblAHZ3rCzYYgfL6g719j9AqX/ORY2yHmm107HeHUEChsqszEL
D5/nHrv0GDH9huCIHkolmO9pvEs6cdlP9kJSl+Ij50+P7kF0rgOHOooV6iQjU/8z
B6Z0GxjhAbNj0LIDTOg9JdXCZZBR2fYxxrz5mXDgF06SayYRpF77sYMO2yz54/5u
uv+8tDWVLl2d0vO3oxhx0Z8fUN76K1tBoN4wD05wKWLrG8/D/tZWPWtI0JNqIAq2
nd9tbMaXk9GCkOhkc9j08ROcWrJOtL3rps3kQBlWK2G3RFdvKyLnKN/dv1pDZBD9
t88zIdvQxQ7m933qFFvULlBIwhYxXM9P4fluYjULB2qiifnH2GFKSiTrKBQy729n
a3OJgyNrTBHghpcG3JlUsfcjnEiJ01sQwWw62zYa8ycgBQMLijj62y/ppN+KFV1q
5LU7Z4oKbnMfEW+1UpbOo08LX1mf6BTrXrXY4DoodMMDjqNLR3Y/ggdVXVJuI9oK
Pl7RzeGaTsRXrpVZBMeVPq1uYckqUDxqHsNocP/l5Uh6afGDj4PHZF0+87K+50eQ
aXBUXtuBP+H1/rJsU8K6IdFOXa4HnBarBpwYTOhQ5idyPj7DRVxhQa5O1wef6tma
`protect END_PROTECTED
