`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4LgLqcKsR/K4CL5yNZxXMdLPqfsr4fhuVeqZKBnfjhQGeEHxqwX9ie9dHU5AMrqJ
RurNhJ3OHgXO+x1Pb9fJhP9OKx58u+sMcTF5C6iC0gyn2zV78GNDWHFKfv8VZr/U
ID+0SW24rmVjEimTQf88f0dCyapSSlV8Dh/t59I9Q7czlJyBznpqav1W0qpjYTCT
YzHlnBbqC2muRNI4YtBiBmsTEfhykBXPFxZUij9++DIaW2n0j9u7kUsVtqA6jrP8
1NhSDWHXUfoNZL9mH8MGUwRrIEWKZl9KbBkcoeeRYnAEWQ1SYhts9a9piNN48+mq
Rp3/sexbJzYvuVV4gep37apAf6KvnVB4tQ9lrTvva3NQX6S0cNtFJAYTNaROHCOO
5DnDkREgGZ4B4aUb8+1MT72OL5NvljrTvtP9DkmvvgU4dF0WoxWgSeKL3HKl7iGP
EPmzXunDwE6HwfRycWhTJQqCYK9imxiHG5GuLm/D+wFph8dEgLmUUMqhYQHorZg9
pjEN643EofYMzEX1TQk/bKVUfFFNi54B1BuqS8RCQasEAqew/oxDIm16rbxTyboK
y+pOlOu3IbsN+37/bPoxoZ+X7C9tVkdKXYMxuZbHiT/HRSmFaxf/cBMh7lh1U2gf
U7PgO4h+jn00Z5GYsByggavoKj0So9W06Vvc27IHxTRvCCv7TyiQYav0TWFfMs0B
45Q5PngrOc/98hHY2Q3uG1j2LeAUmsc5UAbuI6/BVc9ODCL/vpstNsqI4Ee1o54r
uwzlXkmHI3LTxH3aPvjSqL2ZIEeRjb3yTS7tapsLOHk=
`protect END_PROTECTED
