`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eV953mjJ/FCGo9J0brOsU+YGWAWDIPb+rEiKdzsc+QIXtkdbXCj51KdcHH2q0lwf
mBwZjSwN9mq+3bu6pfH7/TCvOUGaY5SILkrqGSHBRfS1X4OEiVPsc47t2wPSJqR2
0Bmv4YcceTrLWrjpG85qdUJKCVHa4pfqmz6Zma/1F/yBzGH7/YT2pNvfml00uzUW
RDYc67gUfyk315zPSu0MlBaHUI80wUa0oW4A7rKCk+l1Oh6UzkJeXkJn1ZDX3M1V
95o5G/d3U2WmT9nFM/W8Vx0NraeiqesnQJDs97XRGZrjrh4+6HJUvd7M1iTaRyuc
89EiBVni9zkywaRHK8gq9k8A9PiKqY6qJJ6xYwOyW7obKCIZ1oYTiKoNkM+8X3j6
VTotJOz8+c9JTqbiKVMxrkUW5nb+19PRosOI4wtP7tPfIl4Gknq5SSjgN72602jT
Tpt1SzwD+rA3gp/DCjvGiasAXMIg3qv8N3Xj9b12cA713lrvbguAQDCy/zDJnDaJ
nfWSbNSl3HDXNaxwVy/qgaFjJuWAFmG7bjUaLDgEbS126OY22q4nGu8COCu8xZqB
qawTIYDlo3uHg1F0zhc2supdDFm8ot0jzSIgQTqunpNQ/OGfxrIbPGaFh3luC1MV
PIy/CwjEds6+jOjyO4t7jt2oZzRQaAdOVP1EcbP9cuxfQOvwKD0Y/0GEiaRhQ5fW
UBBL5cxCAibekm6zDyT6ZmPIsnN07PsHd0UikvcMCUo3pp3WFGtNVnlkodlVOsEC
wGRVzROFKwjoFl4e4ynadMINRvEa9qLmDuLS33Q71s5nM/ABEJ6huJJzW2tORS2Y
JxSieBhB4xgmFIOBwjZZw/KUxRwv9JK6okdTYRbT7olh6BLCQ9VYmDKa5QwxdG5C
THV0HCpWFHS+WB7xMYTby21z62XAXp+puTYuIqw0ey1HUlP6reloxhTr/1vp6jX0
IMacAFlc8qtVXyrkcchx9l9+XMKCn/aW7OPPycF4JcBLqT1cPJYy0tb8li9ahWBH
f3JrX4kKMKb6FumSv9eOwp71ZYQoGxyvFLB8Mm6svYvjMHqrotrp7TS4Krh3qzDR
j18kwBEu60wD2D279ZjSgR7ebdn9r8h9S0y5K0FLrDXg3vtexVjWSDKh9Oa03qG9
6Fic6jW3RQM6++PW2b/nGoFH/D8me9poiwdItZY9VQYJRzN1zXQR3GTqnAM8rHYl
qb2velsl9Rh22k+C1FKV4lOb2sFUpB7J/qaBz9ktUkHcQqfGzESccxhoHFECucIf
vbLv8TXgfUpcVnQU2FWVVnIPiwwxMKX0C/iNIEmzO3QHToOXyNYNU8w0Q43zhrBI
PTfI3bvDamHL6HbD4boSLzeHXf4LQ/uZLw4ODNxbQGyGfD+2YlzEM7ZH95B0CEL3
NAc2ojMwt60L9JaUJtdQSBlcQ1GIsPzUug0SrxMSZsTHJdxbuCsdJmQhJo/vrMx3
GKBU9vgEKmNCT4FvOg9/Qp0TiDr5tmAHl43JtleBMZ5dmr2nmuFA0RPpDgPEG6bi
yOMI0S3Bs+thHyzMa4NazBkpepzrzKeVFh2yz3MAFH6aUEyssyGjBxBFI5WqjT2q
Mx9zGFYjMhh5t6QUjqN5+iVpOlQ70QAfGFQ7e6vDigZtvK4kYXLi06b29fWERMT/
gBuSfI+qOaKVHlxIwxSMXLP7Su4H8gRg7Xpye/FGkGfvwf8J/k+MR+gj4OX40Wd0
dL5UHgyWZjlippE9OaqAj3ET5Z4wc8UAsuUH32Mk55zPMRnY0/6V/mmY89pjYAkA
I+HlSq+t2eszS37TyhBJKHhzF9jgHluCHxWT4KzUxdx9/wmthM+BOxT5JjdRpJbH
ESvp+B2MT1BRytiKTPMvYvnUAv8p494aB+zYEM4dWBfqbnFbubktE1v6RsdHB51m
1vfI2ausAbi+deOmQkEv10jAgEWiEvS+gDXp/tdNb2B5FKRM+1eyN3eZF/h73Aau
jyHhqoNMY5oXe+4eumZs4ijCa1pBjaa+eQp+cPg8WTPVzHipPDXZHXrPrFj+69SO
dUcWbzbwUmdbXplkSZ3TGi9KoH0+oGDBild3cNBhz4HIKUDxECK/8k39TQju8WaG
pi9sLDlQT8wSBJTEldEvoUUSW+xyh6xDSrQrYlxsitFVintxzuardegN7Xba4pjI
oGkhkAYlZuEthKcJeq1j0otAe6aYx0c0SSzZxyAKe88NqBGGqASPyUbgd3gazlX0
7xPel3eHI5i0zu71I00F4px/asR3DS9zG96ebRY4EjFe4Q7a7emhTOAH2EEtjEq7
2VJZ/WKnb7SiD/lAtrooXLEn9ybDVhlhVguyg6Ma1ftO5DIJV2hnwhD+ujbqp5Xy
cSOyilmpG2QGCPqp4aK6DPZCG51wzHhE/trSX8mBitKRUXNEZ2IhMVqZnzrO9Quf
QyOifojbRlbSP+uXe/mWizGV0j62CHsQRn0oI8LyDkECEas67eq8hAwpLzNcr02t
h8qdLzb4ukOGbJTi7DjnD5TbimKURFPVISn/hjTL7PIR+5zPTZZnJnAoEUbUnRg0
KIEl54syo/O5c23WZ0UlmrNmbAokECVbDvrNGb6sXshE6YMI8rLCARmnu+RY3hZn
ONGjcd2Hr7eILj4rFKvF4LjfUqsql/v1UxOhPP1dPtHO0U/+sGXDBRBjLDInNAmP
G51uRyj4e4tDmgLAnhjBtMhunMBQOdVAeV6H+PL+bXZBsgSUA7N5w7y3sQHZuFvV
eQitu6AyrWlvmY2bMvTxHv7g03Dw91Yl9JY/N5G/714EbwSmvJMQd3M5KvyVQzP5
YO4GObZTYPjXDXiHfz6u/e7yqSWHOP/vWPwmbBmQPtTyHgpfh/jws9k2Q5ZmgWie
exifuuuITg7OdZVCUUi40xgv99icFk2gsELHhGF2pNs=
`protect END_PROTECTED
