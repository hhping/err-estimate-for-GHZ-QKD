`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2H4ipi1GwhJ1nFSZpBGUQfw2VHUcBjL8ILilPVig/A50Ak0wD8xhi6wRWPtfm3lr
SeKCwDdD1Bh8zm2seU85VimVJ5tBiQiUdJsfmIHvrnNeTS/WJzLhecsPKlUoDUdU
E2vvc+8ts5bhTY2tI8mxiY8xfQqnoxm+a/LK/NAC7YCGPCNZyEDzHuivT4UZo0gB
Q0n3ktksbBZ7+hZpclXZP1Var5+0nqNEsyBBAChEWVdXTlSfe78nX/7FzBGjCKTI
UrNFUCfp2t2JC0eVdzjC1C8NhB9hCuxa2tYUfMxParMCZSHQEFn9oubMF6MTHaHX
PYA53pVvgMRPWAK0mXYiXMJvodb6R6OKyF+BrGBhFCMACH7iyb1MolNNhRvufqu0
wZUEelK8NVQumnQHwkeF9VPQc9PTaHj6MXOgc2vG+V8xrg/L9JjZhxnKTSaEh4Og
/MeZbK1alAWhmQwcidMVcsrGi+gYlOJkOd24c4bAOvJ4hRjFJXYCwAw51YnvOG5Q
WM1aLQynngiJUZEqzuxERkyZpvaaFHTnv/0LCUXofxqvznlLHIt2WMHyj0rJOEm3
A0bxIwi9Crkpl4fnJpsXzML8QfXAma0SfMKqtpZZXNsdVrsCl4awDg6FjiaWqg7y
dju+of5jyeQoI0wgevNqTZUXzJStK2V+ArAG7YpdB5tYGXe90XHmCxL2xUs3O4kj
qcLnBC/D09imdZpoDgtsEFeCn2zb6ZKrhK0z4Z0RvT/ud9HmzSEoRYPLDD1Yhpxj
5RCHsq7bomn7KRbUU1f0wLVZaX00AMHodiDnNhN7Dned4e9duOPhQAsTlbRfbZyj
avGmsrrt71zVwLuAZ57yP3ke6qu26y/fz5NFvTyTvFVNjRu5sslSzrM2uHZah0qv
Ooik9vsjKMzg32OZ2xUGYg==
`protect END_PROTECTED
