`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlR/t69ZhlZnY4sw80wcQVUjcD+sDh9quv8ckCsVjJbg1aWlX/WF7HA275PTZI0c
mwN3hHrlUJZidDsctdUUhhbhr0EEeholL0IfUWUAlmDEkPBVjSU+tjhoOR1VlKS6
SV7ULUXksSnPblYZyxNBcQJLktaoDkQ2d9Ywp/5XJT7B3kyEH1rp6fizQom6cOQw
iezBxDdobSoW4M5D76K+ZypX+mLGEGHZNqeowV6iL+4oyblybqDDii4SNo4rGGM2
wOoTqvCqRlChgmDstT6hua2GbezZtBpA2aoXJFL4YpM0n/brwwEvRKYKL7Zj6bPQ
0WTen2EnRNsZKiDWzoHmCUYo+ap8uLz6l5kmcCIYP8qVUjTDUQ4z9ggw8rREzFM/
ZJj8xAxmUf16/5j5AofIIbNnEv/HSiaPyhDrZh3lyPj612vH+KcI/aAkFYquwV9t
API2TgvyUW/HWA7MiVgVXmE2gp5VZWW463Q6UCZcaDEUfmjkZjUHGW2wqizKG+pJ
OtRK0H0dDx63OfL4h/38ylwZPx5DYJw4ryCR6ThDweeskG5RgGBeb83bhZRGdw6P
psh9pow2LZz//lUbl28dn0ejiaXb1KFm95cayA+mNWeSqUZCzDXXdhQA7y0Uv4OI
fgLYWyPY1NhfPbsziAghJCs0BnLhrW0vmNZpEJnOkqiFITJV0Cbh90suA4XNSIB8
AdoyzQGwqOlMs5CUcjCczq37quGvbB7pv6OlOsbk04ZHEQXDFoON8W5nJfDIIJ8Q
jBetYiVRhVnT2Ap6PwwhkwAYnNg3DavW6qYSEmztAImvXjbFGjwaN66N+7svgVe7
lLM7chkkraiR72bQZ3VMwMLz56KOktrER5S59923lMFRoHiXMM1r66mUab8yIlKQ
5zGfi3q2qyNsrfPZWfTFL+nYvku8OgFn+ce176D5yKXj1DoGqxnfNKQjVJXcCAwJ
wW6sPjRFQ9+hbT83iW4HnBgRaCQntxW6fWKWvvs6ERoB6G3hT0WE0H0poeLILaHg
LZH9QntohtMOzb+TGDbT0G15yMnehsVOgC7FrBAITiE41LB8a57rMMScdjk2Wo8x
a7XLcFhgaooAhfN2hKNgouqUI5nVm8k1mVayjcbZjnUHGDLFmO8gFgBZXhDaCmDW
sp/FiatMXDYsq3Rn8T3JN3lDGSh8JaJBjHWtrrXkdK55JgcXmaRTHbWKd2hCvwP0
09oHW0fOL8Ho0PvLKfJFX2cBUYc0aF67VMUMpRb8mSsTAkTm1ahBLQCkBoegQ0dF
lMXuWusTHKdUXk1b4iw0knuC2sNZ9OqsOAdiU4Trt/5MWman19IXVNWHlWwKh5Mx
qOggGxFcMt853iDxs8OMezx4soixZggr4xPItYZR628xoeqhct5gLF6p2gGFo2u6
PsAE9ESkfpdp4s5nRjI8svTeaAY/g4UF03ZGhxsbM58SnE3uaTH4dy1Y19/15uLZ
PywWxNKNzoyXOs7vkpTB5eSBYMBdipwdFnGN6pRyFreEGnHHjFB0oe2c3zYuPYzN
AHNvMCJn/3WvPdknPZQcmw/D9RUtljXfxHAnXFVy6wYe7yF7T49H3YzNqkIIcE7X
WnriMmdWSCsW3Wdm7jfq4EYD1wDo/8AGWUpi064eCQjcn6q3pPjp0UgvaevcSvZ+
imUfEMkKPP5z/VkwABLJxyTvvMi4POMuZKbhUfAV19Fu0v5v1yvHZJLhkQ2Hz05p
rP/vEn7n4T5GdyoQwYqzB5jrEqZeJlrqBG9oFUdTpKbjVKUHF89fYuhP7Coqpt4E
0sskhelBweeJFXWpkVS4UOEmyspThO8QVeqGi7rKYU+GsbQ+4blhXYu9dvmQqV6q
mrihN5HjDWVgIhXReOY/XHOwGtMmNHQwK9JgtVy9Ka3P/chqPPUlU5tYOvHUp3+v
Nraf6+qzkoSFouJqfqxhE0ryC4Js8DrTjHJK4ewh08wAGmm49jE/FR6RjrCHx7cM
dI29pJo/jVM78yKcs9vqUD/xCI7bk1yqFHOHBaExSjPR7rZlm3ojdP5B35FlGUKv
xAKHm4BSt65chUki8daL8707dp0nawL64izGYkfStjIoIdVARSUuyWHXF/sS08hk
X3LqiNIyMaCEwqbtsShKBDDFwlXOusULtpoUubGZhDzHqrQsOvpc5i/4qGaTcIVG
FmEkW/a1sLDF5C6iWH877JfMPystz2iHSR4bfTBhKa/G6Km5/gy7+sTvJJ+Nnqa6
jr5IbpEWL6gj3IziX/YDXnDVY6F5nMyukK2fHoFNXKkUXSsG6QcexF7U5as/PKif
i2wv3MbPPbGCLC1dt9o2PLmXtAJyK9bOnD7htjnd27tdiOiPWfR5I36fxVt5MaJt
rkadQKOwVM3QA1ATBYXzogsjNizuryaNEFgiCVp+EF498kdhfAhBiMRfeUKktQsw
mwFfxwjyVaOS2vbQVcsCm/GSDMJkjzzIu/zthQHbH1t9X3Cx6UMMa0mq1/KzoAFx
7vDQDFm7gQN+ZSn1llFN6wxTZS4Z6MuBieFY9JlFMSZXsKn6wQ3iHWiyaUIE+zNY
XU9pPzOhHaGbk1J3/AjbbF9D/GqIaBEZWjVpdPwDGrLZBSsp+A6Uu3DUq8DLv76c
d2wU22XEoW0RcOPIADcMKF4l2S3dtQ70jrlKeCaToNTwkPeOVSeO5Awy5JhX7U9Y
He6EN6KyYw5WAqGWqOdua029kz1HkwcCMyT552OXYYMf3ZQLlQ1lhw6XV/dNZRBt
/cEgKl9703pzI+w80+vJxQ2CsEy0NGpO80xHdv77W3QvoF36j75qgFvZFLxAK2+l
j5u7Z7/j8qjJm+n1YHzjDY/G/coCn1V7i7ATqg/sS1M3PQhNr7k80GWWjzwqh7uU
pKL4CcFyT3mqny9TljQgRDiLIPCkptqXdzsxMYC9OCRsWha/KrQc5q8j2hDvv4ue
4e8/XeJeA5BBp99wkdPNoYFjAzkVvU6oF6OckFlnnDFNZN6s3XZ74AQ16W1+H9VN
lkRBTqQEywSHl2uBdiJL8D4+gpxCapiwMCuksw6l2lLSjszPhpfmuELYbKkOrn5k
rQf0CjunbG5qfcYv7XYzTidjagsIgHD9TevTEg+IRvEH3IGHbHUbM8/er+fISlH9
B2v29qn7pAatKPU4S/6Rt81tyZku5CgwYqOkB8N/zm6zTYdfy/USiWilc8FxMZWY
rLHNynUaVOKTK3R08BWk1wxOoYlnVrCGGiPARqLbp0C75icMqadaBxhsS+XWPeLb
RY+VOvlJfNqxxPtEeJGVtC1BM4iGvhr5sVnIbGq6AxIe9k+jnclsmkxeDp8/mdl4
YTBS4DvbctZpkxtIH/4jSuyYNs4XvQYfvRqIdm5B2buERO4EozqISOSBJNAveRrC
tPLqZx50h82Qp1OcLDvYU3cqxcqEg4Q8paei95xhWor56PllopMQzHcSR+/SgI0V
Z+3LS/0VoAouJf7yOLqgJq51JDMZOgzL3yT4idU83DC+OLeb/8Whk4fN06YdQWD9
issAwZIkvk2PS/JW0kDO74+rN4agJy0AP2/Mb3hoz3Gx5kaTfwN5MDKEKH3p31L1
9kpexEJMBYD8i+2w9POagDa+y9aBaBnbE/fWZU3RIPitVD+rvfK+FmmH1s2hUqoT
Az+DOQdSDp5bCcjK4bbiZRtokwwEk0CI6zFiuKKuTETUpM46UybRQkllEjkkugoL
ddXu8HEMNu/O7Iz0wnLc813Lod0UiXdkSWlqvdoignkb90fvl4YtQ9IXbOjCOwj9
kAqs2wTgm5K+Qp9io/rwuXOJ6Teod1kFKW65UoLzvmPKMNnzYGm0nMUhUy43Ecxy
LAcegJdnypd5ah7K5oPCK+3QemEm37ROyN8qfRB/+0yRAwTc6PL5mzUeZyUOTMrH
c8O4gyLgGadDd8Snc08so65AKZpjmojUnrL5W8tZWv7iK8R2N6fxDyNFYYWpggtb
avPXzUi2tjt2GFlljl5UtUBACq2fvfSWAew/o+dww/c9F0DtFpJqakJ9G7kQbyVJ
WNDSNJP0AhDH+gSaNCmmyD/mPbJIyXTwTBcheRi9rSxGanNxglAFXivNbv6Elnb0
gBIPv9RCc1Jl/JgIW5Eu7KqydnHqUjPQSvFdlylrinEuS3kPj/oFAjD8BUWDnXXc
rBo1+BMVFOJkU8GH+WsWn/JScqojbn2Qu8FWvycDkv94gzb2xfPVUYVnItxHrJhk
cTQdRWDSF15+4x9wwWfnTmUeJABadl7Jw4vbLZEPmETPCZXXK3Lm9cc/s/VzSyEq
X1s65rPXk9vETpH7JRg6nCxhLz+oq9EQueN+ihYC78EjqRiQLn7+dZ4KTKf6RHBC
V7G7TOggK7LKSEjnACDoFVfwKlHg1TWJg0CSXf8tQTI5yflABwIzZqjlArTzWKTX
AI7ndx1gQ9AwPeioGhIHgOfTpDS1BpRlZHp71D34fXUo7J42WBwsFLfI4TWLBcsC
a3Q8N872tqADpGjqrD8rOOzxFm5eMEwKdM83LIljn6PEzvS+RiefKjlIhuvvpoV+
33Yk1YqHxpq4x0vGtCgfmbH1P7HDn/y32UTrwRI29aeoqcltHT33PEOdCB28/Wln
4Ei2caJ2blw3C69XqfDKP8Z8XYaNrfxk80Boj/amp9MNZFKdvTFM9p4hg8zoOXL8
U167IIf0ehn6gjBNe7q0Cw0axlrtwR2Sw0jbZUc3j4KZ+m5j/zhq6UeJgP6QNNTv
5gu2dZjORAU1HzNlQyyrWfXgvAcEa8g9ZXF+J7D9yE+M8iEQLmJjOqj5qhY5pEHk
eIto/fpR1WYbNWbeLfq693v76KBNgK1kSVAfhp8zu08ZqwWDfPojoEzZDkMFwk4G
0hSpZPEmyrRpSJF7KHnCEvcb2LE/Lws4ydP4Y6XiyxNRG/7lxfZD6VbYF97gh5XM
GkpxGMjhC52gC9NQ2NWwVfbs4do3vrIpISQih4Szug08PEK1NBq03L9vOTsG8Z6p
g3idUaVm0H7Q/zKxwXrVP06+WE785RA/RuJ3EfOBI0ES2No3XqKL5Fv2RTGl4HNl
Qag1q4S/G23eJuRQdjaSTKt8isUnvyk7wePE8kmWa0Fw0dtUHXSW05h/s5mDzHko
FDumGMQFT8gknM7Zxe5QjsUe/FvNFSXBieRIdnb6lysmdgyVz9ivbj/gHvOYjF7H
QYbLFsJdcrOsb3GsowzUsxteNSJfq5cSpcXKYi2q3ClMTeDMb3QoPRODvLePi9Zh
OS37GbbOt6Lx2Vo/jtMX8w5ak5CMQtaqCbK/pJtTol4YsmiOLor0Pk4srj/ToxMF
L+J3DdSHQczYDAuWrp6om3fYR6pTh/RDHm9NfMn0UH3MRxBVUYqFs24YnwbVmcb4
hXNs+ZLEPMsJeeVJkriUjIquEUYOBxC8gikGFCgQEBNxl1Sz+wSwQ28mQBCJQR7N
LagwameykIizULAcKIUZOugDn3YjabcrJBmgnr4Lqt0aRmqI5BGq4Is4CmEUYxip
29LsItdHff+meDWFPipuFi3kAxMQGVKrAj9iNF7Zz792uNcH5LtPjjDNeQ2+8FDZ
OLP1o7EDyQJZvqY1Lx/fw6zobkeVVSztc4o9TwLOaGL+WjLJqZKxW2PS1Z6RBqFb
AkswI1D+aTgbZnxY3HyxSygENH6jbWS8x26tHVTAiFa7detW/cmUqMPkMztm65H7
TyTdfrE2r3CeaBAYs+uQWCJzSlYOcPi87DfTeBXbL8Mj4AzQd27o+C0PSYsyJ4W2
mIIs4QzLrfUolYdxRdIBQ0movdpMiAOeofNZQLGvQfhkksvZdec/tx2ZUkPqKHm1
TJcpdT6oCqYA4/mnPfhLOUGxrNXQdCapiJ+xq1pyBwcnKV8p7ENFgkso51gIXmJR
niCnsj8e1NN1Ni8QYhOgfhjOctgPcJHmmLin/a38FcUXX8P/Qho6Bn2Ax3Bp3XI6
Goy88Q1Goc72E90JpQ1bSnGqjwyKjDQaZcUUlC4R0KdRoEl2LbQM98F6y6eTmLQv
5BF88c8Ka/DC2VLhJj6iBnURH0vr1XkOEgOcZYDT+8ROUHcogoTLiGf1ZId6Cuew
+G8tTqEc8aT10dX5uiHnhtANch/r/DP39wp0wQjB4sPkmNhZdLNVTxuhTqbKlx8Q
SWsz618lxLTC0fUotYFecpILDk5epoRQi5cD/38rm6aeuQKtYTOyBHJSDJLcVlRM
KeSwSDV1WpjnfapbwsBz38QKhgoyW9/vY2xeCXIA3w1MTpsOvrYv0jP7/bH4IzBy
Qkzwm1HIQlk8FTocLcOnoleWqrFh316LrL1P2rXK4WJb/PIm8+0j1DfZr9KPWDqO
iZXhOKGNF/WD7AMA7u1SdSbwp+6SCmZ2qkSKnWzCrZZ2fj+XQCFHQtHaxBkKdIFz
00zLRfA2vbZXoTxsK0GpcmMlV5ePsrIaOVmUPSsgOsaAnPSz/Dknz/dhuUlAPUab
etTncyHHItZpj8DIMMxaMcPfx6ORmCMDVDP63q2z4GUfxBGcV9DKv8yGEMkH98Qb
3guC6/BP0JLnAtfhtbdWQEzrIrzcTslWzDnB8zYSZE/bmWaf24cN3kc5foP+IBE2
q2595/gd/9bSXbNCpy+Pq0HUhUqgof9LTv7hP+V8DdajE0HK+jq+7/CKgG48Aipv
IA4PNdtfd4kKcGPliqBKsDNkha4y4kRdsyS04thfBR7pcvmuXiTtvJ30yuRJ2zVZ
+/35xN9mqIl6Z93g+YsKFPzJVhzPIKd6FDxlyjjFyO5EE9DnUtzbz4qTuZ1OiSPd
EEcWCP3JIbiQJoXUWkF84nti12g7vjVI66eoVj2/HVJjWHyp0g1xynvAJYl1TCgN
mxa5XMJ+f0n5Q9GLczpNAiDFpZWMkg+2j8+TPJohLC3MwcFZah9q+vpfkLp3NxfJ
PiYczNcren5r3Ip/nqN3YWY8SuKPH0dlmH1Aq+AvPjVVckS3qPrIzUQpOUuOFCI9
WLrBhA/2+UK5NXUDNsldIpQYCvoDI634Hu+NxEm9Q3z/8WGGG1YbQDqcpmEEyzG4
vQtk3E4DNY8QQUZJs/fPp+bB1h6axSayu+9d2mjz6yIcy1po22ivbjubNJAcHsh4
yZsJl3jFXYb04IzsbMSl67RxsycwD/+GiHT/EObzXhQW7j4HNm+P0f61EmMn+Mjk
PkgRyMQjjB1DiT/TkCP3RsuDV/GafjW+dXI+/uXZ9iOeoAroTTBqmK4zyr91+dWW
FMEybyVIYbF/PDq0tsgXhknVb4hl+7XeV4zI2CMgjqBY0ya4+2VmJ1zi/Xf/5HRm
4D1T1mhn6Vux3IwpZp7L7z9/wDXz+uEspKgCd8GfkMeYs4v7OeUVJBdqdRO9YhAi
+5+P9lyndCwPSX6PqWz2ZjtsGjWvmcNnLtAp2nzWpXhYPh4YBi1iAEHm3O+yUS9I
f0Wt13pdQRy2InPe6Q/tMmLYoYHO45R3kXPYt59cpl0DDnJFt3Q3vb4JpIvEwSvT
lCfMkJqRACiAUGPfcX9f1Zlu6X4osUFg+j8k6SfUZtDCJanXUxNRtebtyQgsKkH4
+5/mzzr6gVCEuQEuGEAs6XGw7aH6KC0pp5FbEV1RcIulx5Cfm3D3bzvegPpB77M5
/IarmTBYZ13R1AmF5GMKQX+Tg9fHCo7kAxrnopV4YM6T1YCCAt7eNO60D9c+8Xc1
SZhf3+qOsWXQd37Oil+/yrcvpcL0X7BVdSLgUFZqVeKuaawElka+sCtASm2YUmoF
Jylhr+QNC55bhquxbDI2nLvLtI1IybHOEauG+6vNiiFLk9Fa1j1DrRvoLez/ysQK
gGI3YF+42tHxalvnLfmVMsC7pVfQwR3v7aH/CSe/P7rvreaJoV2A0HGoWTkz2lCu
bkHIXVThvRD1+84ZvSU4yDjAd2zHrDxumVlCkXAszh7JnaDi2hAJ4YhxPlDjJSqS
RF82R76/uYWp7MCQxIyaYQfhfwI4NJEo2uAtqhQsOvtCNtMfwyzkebY74f+MNas1
xbwUTRuOCU6JDyEHsvLsUgzdH/rfU5aKnjWaNLwAR6rBwu4mJKirB1BqBWS35B7n
mS3YIYf2TqSC0nuvZwB0hMQmqdGxzbwWAITUi0LNjYetbvKdQfLjpbZhfodW484A
LhjBMdpkZD760e30cmTwFaH6YjpAsycRuhvmS1aX+BLLeXLXU6lU4MFSrAcOjg2g
yoAoakthMJIQ86QPtBphgVUGT+mW45BUWlp1lfSQU4Ysf0E2393s0LwjIeTOtYGY
TfVtH25VFz3t1TIEt4l1SePAvdIN3jfB3O12RHi8jxEXLCjU4b3pfbAlZN108fIu
ZNl61GONK+FC4c/mcXZ2ucWYnLCquDUS8n6LGb2HPRTdrrKpkaNtk+w2EJKKWDIb
b2WGlgXpymFPhUPvGnhlAGblOVil+O/AmRoZeM8xIxvL8GARL0YgOKmU7KTsPPVe
vvkBP0EaQIkx8+xIqZ9+S7p4atA9pI1O3f+Wp1uCPeg4XQkk0QkPXYGPj/E5QPy5
Vaw/MDI56Lld29APPoD4qxWFBrVJ7tP9ZEHh1gbT7zTMXV/v9SLEeIQYEzqBHcuh
e4VAQcxu1eiVYrSUqhCbQupCZXYHPY8nc3qz80bB5/LqWV8nWRKQLrmGvKREhUTb
B24j3uMrNg8a4YcyddZQCnqz9blCqg8WEDr3tckJTkTgAiuERsPMOFgvG7BcGyUP
qHpXF8dX5t077lAOSYPayIxcK2nuBa0+ClPGp6WBsphvnATyksMn/PRf5ky9c/2S
nyR3eryPbc6am5AqtInRmfAlp/h0hp9KQQHwONuXcIxHACNhC3JYbc2esFYqe2oS
G0Tjfq0+I1zYnWYsTUdL+PhCFFLDckqhKFBF9T22yfAyTkjv0psqMYsglL6sOnbn
NghsK+4wqWT1Od4oyK3bzdfxbUqVEkanGFQVCebxDoTHtGixvcKhl9/gl8j8WL1B
Y9FbGmiwf8EZK8i20xg57KrbagN0dPqf0MrHAdw9flaM4MPNH93Galh17WP4bFXV
gFVkR5C/I7BYrs21ulY66Yu0b34Y0SF7oRjMtZtL8KxVA8nSbmvUgp6tCqZj+Eub
vcovI8lZp3Plv2xCle2oLPT1884/TdDsK4oACLyDARSbBCQ7C4QXG4ukfrA8hZpQ
kALPUgu0hZE1wigxH9IFjHn9kiJ7qEvrj6WRW4k+0YnJ/ZGgXL6pxC771o6GKOx4
z+n/ZElNFx3dVQghIj+6UsQGH1LUDJiI37fjluQzqZdAX2mnU2aqydG3yx2eG+ak
uWbUZaoOYEvMe3VPnxlR3Ny5mIeu2CNmaY/Cw/BTWRAjHHOvxNxyEi2whhzCrtny
hPtkSDbE56/YeSyQRuXP+vFIbt4jt6/RT3e8CtoLmGRi5kYDUzyoOvVt1f+q63Sx
Iow/V82hitk8+iMmyixSlMGcVU5lIA8ppzOdKB0qoiCN7eLiIH3vwgjcoBA1gcQy
od+XuDEmRF07FkpUxss93Gv5Ay0J9VnFKWPtU2ru3mh9Jd5zr5Mwl0Ds51u+hOSP
Bn2x/D7unKU956AGod10liTyWBrS4BKwFA0v35pkPBkhCtz9NMFki4kVEmpo3VfS
RsMi812nw4UxVVIDbDCVv6xuSl7lAYrH+P2O80/9UOlFPlmZ6xkFYWX47BIR03ht
N9X8u50KnEvWX0rGAjfJ8aTF9yLB7LFojJGeMYOSqXT5NnkqHQf0RrVi8gQ3thhc
KLxI7tx9L1/uDNLepy87XIjMZjPqNBJaJysrtGKKkDl+9NCpmlj2NtpAX61vjqTd
SFQ2KuaT+g2OIANoHor6vSAHh2fS4splAj2hSMbozFOo9dm6pKQtk002wGcxChq5
tnfukpmIJEa7dnFnm8+zGsAxXCZQ6mB3O/Fo1mww2+jlHJHPc4mYTV5evCYxvf2T
YschUuljt5iQ3pInri1xYbqa0qQFFFdiXq/ZdaN5McqvszjwZBjHxKMkScI+/q5I
9Z/vTAqBAPU9DN1BDUoU0DfvsMoVN9KqeS4pyGMTwnZ08MH/fKqym/hsnFPdEQFY
ocpkWnhZJSSuwzUCbGmiS1FjFapRquslvSilQO5Z/VHUMirVtxn2HvfEed6hBST8
n2ORW0N+q2AmdXFaA1pceE3nftMK/muYVtMrPBEpIB4MRoYK4eG4JlatWjVjUZUm
pcY1lu3Ct0Lib/tKOsi/itkEjaW52y4ULyctP96rQodX6Ie6f2DdC7HRAGICDmPS
dLh8/Unmz/7QRKHJxYFr+ABX6+NtC3foix416IrHLJptC2zcXvoDA8/z8/WgJVCG
u+21Aju/8M4t+d3X2aODFN3kCZqeLvXuXwZ0Z91iBXNvLirn/5ZxbkhFmrH9GvT5
L4qJ9XzNuC0vY2fQxpIZscCgXVOkevjvhMSxT7KU0UmK6DumXTUJVNrk2uPniFnt
MqT68T6EE7LMTZxP8ndiAEFnTwTswZji/5xdVGOXBiNaSjwVjTz+MNpT/sH5VWOr
0x9CqZkIRebS3sztD5AzRC2fW2hWUnKDzRvT/T8PhcOF7xhNUHtR4TuNNO/hrNsP
nmsfmE2OCWcYzzrINrLoBcYktRgnIyTRO99BuQ/OifOqaw8ryTI19oTwTzr0PmUw
YstichHr5jM/5Uy9oaPxJ4FZ8u2JbaGi9fG4JvsQjAX7rdFm2Fotv33xc9z1baP4
MwbJPWSkSTv4FqxjrQfpE3Rfea/ngvzCnBVxVRBL5jbz5jgTdPRGqUxEgWC+Qx3k
0Suj8UNFP9xCOPoIjrB0L+B2pFzeOZDcfPfSSkhdmWNy8yxGilvODnA6AAXQHVav
bspAKykHngowvN/EI4LXnWIAWwRJjGr77U19x8KoPnSy8XsU4/ZQdt1RpelCddP4
i8hRZOzdIAvbAHjbpcd2xFk6Gh+MnGxF/2JcFH+/ErW784A65GEhEe2zHMaCs7bo
OV4OzV3ot5sjPSggYVTnhVc8wMPN0jiV8hGAiyO0YhUXItwUCUIYZCVBfeN9rUZ0
dSHPX2g94MA73XWUG8JlMcZzAjBdwqdZHmn+XT9LWtSOQ+psY92BEU9dYcZMIPS4
OrKPl/nwiFFNam9a7bMnUe5r74pDFOEVJZG48vXrSk2+xTnY50JzrOvuorWjPJBl
P9AyeHVccTlCg+YKZiOwRxcUGU5cIRRKq/mD/pxEcA/1MJAT/eUXfrf+G5c15bvu
M/22rPmjh+q6LTlUOabAjWofj7M1Jb4Q4RQ26iaE65886zstLc33TtUJodNzlud0
1CXtQDzfEqK4zrazix2FyUj12OxI7/pepbT+gVv00qHBgX+cN9mD5JLUT1cr++D0
UyZxCMcBkTVu+lS/l1COMh22xbIgvJM+znigOtaC3RHV3pRAdYM+fc0i1MI6AoAo
oKKlHSF+2mwLSah1UjeXgaMbJEUai4cRSbNDEJuRAexDTiNIhjAa5RX8RRxw8qs+
SPenR1CeZxjEEB8Zr82530i7QG9lx/N8RNvyhzhNI/ucCO3LTbu49GZ7LEirppis
zSyRO2tK2g+RZn2/J4VN7BV5apudI+GaKc6gy4bh/1JqsZmquUsCSQutQGoJS6RH
JgofgitFzzXY8uOolMYlwHYAtQrMH8o57vViIrYBuqq8o3w1SPqrTjc/+lrFGMB/
0N0n+Lq6GqrCoAGWZumm+jvmRAJH+mmAuGizkpOkQeeoRoeE4RO2CrCMw5NyEdlk
9EitMCyLNSD7Lcarnxpay06tPOMN9Ph1I+9B1q+FN4OWFfg4WT8nJNYTAUzgdVnn
VdCJmbVAw1OucCImGYc7qOGJB+WJwl76zp1LFR8uQcD/T8z/C3lyLrsgg5SYusqa
esDgRDTsUEYXVs/cX2QWc3/tfkqKbJDVTN1+oO15+Qr9Jol8qB5mqA+GOR0W5QO9
ZSTbMlGDnHxaMYdr5M1jPD6pVGhAfAirGpvyyTHQ/a5iZ9Ih5EfOJCCb++W8GCAM
IAOXoXJalui1DVqPg+nYKwn5Y2Esph7J71ObMjmurn/OESll4VMSvPOPQVsQrN6M
TwhoeiTK3jeDff7E76T9hrMIREChry1WYlTRB12Gkg2JGrmr5Ufmf9vaJtkRxV60
5Wmxj9cc2OKZ0DJAavmJTKHwVnT71TwuH+p1BJJhoE1phdjtbOhX29oQ6cDrxgxn
k5hmgyyLwtyjpH5OabXHzEciq8KrHJyECExmMtjmhm/BgPdO2BKQiV0dRuHRaE9e
Qezszu9ngzVdsaCrxcUkYiVNst3IrMEcHc4VPMh1AX6g2pPsRO4n+Vkjy4Q+UK9m
DzhcBZnXoonT8OydS3bLPKlIxkVPsFs6+DNGSvBAmC/tgbKQBgi+3OwcGuSMBN3r
BCDYzshCQwEXH7wYNbFYLCh7Dj/P3+1334K1NVv/4KKxnwww0j1QNjaB/Y/jvsuZ
pANuBko+oMb/pkaOmyxYmlMZuq9nC2e2gg4KtScCcwpkNYlJSxhlgYwVSoZSl5lj
5ijqk6Uhm9O8WTzsG9sU/uX/LdyRY2B4VX8BnnxQh2SALRSQnLkB7lIJaKnX4p+D
Cuhmo0jW99Qc8M7sFHZIxqaDaNBbg7esJ1Kx+IChEr3uuadrFqG54OKcjBEcib87
8z+pTrwVsVOGl3vGzBK3j7rYmZEwq8gKvEQp0FjY+jGGKUWvy2zhF+5WoUmCS6Ag
lGGWD1Xan04EQS7ksKk41TkUTn/vwGB11oCiltOF/okMOUnRfVNBZGO2YIJ0u4sF
Yi6Wo66TifYTVVWFq0EErNZnUteK4Jzs93K6KEu+IasY1XDJLvWSLvamsSZ1tHB1
Ltg/8RAhgsDAlNZpnU01b4wDler32rfvc32SruXyNFLdIOV24XD71tQT5aH6GhGj
k9fI4UG17/H4m2IplRi2/ij/9uZ5hzDlQdwZHhYQEyi8EyRN0AkDQojkophCQgtI
tFoBS0ZxHJvslyuY8DnD4xja6l4rEueuzpoynVhN/b6KHJubG5cq+YfirWcvuY94
3l3Sr73flCUpoCTr6BU3f6SFIDbajCleV+dmuszzxkvfShmAoEsNQGctRPGCuNYc
JYkQLmX61hdSDkVJXhC5mbXOH0FB5Lj4ZzZbZbtNCgzAJsxi4o31Z9Xl4W+DNwqr
dPy2+OMgDAvqaDZvE3H7gOGhW+uemDDlGiSglLFrCsVU02nLnduh/hPPuWIVnLye
ufVQtAM6cJBraSDveVw4YpImge8Gh3Ek9YtS9xkfprmiMltZ1GOj8O5yMYCol0DF
KhlstHuCbUJamjT6rrLXLnQcE3zuKLqrHPlle0I1J3bxZtXOtTSs/G0PipULmYOl
La0JTtetUROe0/ZbsUOehAo5qX9iPDs1cdIOKvVOS09sCHNk467Z2LcfkSDr676y
/0y2YzOFoXzPh5TjODV8gSKUdFRTiBLCb2J7PvXoXKljaCcgV3ZXiVSzFHPSf04D
vlXreBK9r586vFSTHzikGDcu0em0e3yJN0OkIaewJbuuJb18JgAH1Tjh057h+rEe
DSJCG36r/CFfE63jff+Y5urAzkk9uxyyElL6CpoTSLquPTkfPfrjCmhBEPWx2jmG
xx0tLHDtfRxRDAcDSuK/EBMeT9r3a444h5xl2HnXOoReCKC9WdQnJSig27w7qeFS
g4IJvAYR142GoR9358HWR2RYQXyQefTV1Zn6CV5PE1PwbFBTIsBBX9Up4sNf7vlj
FO3LHtr+A+Qba394dzK2FhmkvsSZvSAuqwFzn8c0rro5a+DoUv052FEWzx7Lpf6W
gQt9oQv2ce1LRIbklaqwZsP+XUlsGCPoGNbJ68sJBproTrIEPKvBjtjwYorexUsH
O5AbzL1Z/ph4zyf+YjMz2zgqrBc7m1YRL8/sxmPd/wz+PzR+ExC7VPDw6cM/1L+T
WqsVIzknwu6qhiuHwHaY1jX87SQggyWgxQ1+tsBY8ovMIs589RJbBRCNWvNKI6gP
G10AunqhunzClbeNUfA9L73P3MCfUbAJdq7yBFUeHqD0d5H7vOtrYzJKOcb1VTd2
5X86Mw4VX9twBWiVLktXbG8Hw9eRzeiLDN1nAVAdtiFbQkaTITcjE4Ua1aJFZ8g4
kbiSP/UItK5AidkQzWkX/Ur4jPqKn48UjT7C9V9xfCXSYdLI4rwfs3BgXrVYT64Y
yqd+BN4SSAjJSviTFVf81SHhVB5lIhDr3kRZ1twhFj5i0GjwR7SNqpGhoLNljaWh
jCd5kVs+SpX/dSgfPaQYBXzRuDr4mMPozgUaRbv8XLMZeIuh6w+WZvG/qg1QFO8K
Q6/p2Pa0v8Qg8AozLtbU531IxXuXDL9oHnxH5Gq4GBdtqDSBnCT+1G8YLAVTcpCM
6ZHoUg+wQaF9u5nox70dCQ1CTSbhlzoUo+2p9a1nANjZfduU5t7kned1ux+cY8yk
PMWlKBn8gspR3ki/pxysdEU1NbkOQe6tZyQY6RrjLoJYiuDBIuRJGjCqROe4183J
3bMybCE5oiFqKtdFNZFZ2w6dlGrcNEZrZU3aYUY772q8kTfYMo4609vppB05Sx/G
VIDizRt+xxTqcZYx3hvT8083Zzw9t2ol5bKLkFxsyxbz14R2lJ6nRUaybze+INC2
jquJenjtz90xY+ovF4ajaBND3/8lbxTQKneGWGzfzkjOticWdiyp3656YGwJWrWe
HLU5F1a7j/hrl1fccW5SD/FYzzlZhG4yXjhYROM5PWPbXAulYF2QFVQUANEa/ug6
SLjiOkIrugsXDKknzDDCsFA1u+GC1iKAuyGT+aPOHBTOmVTkY0nGysbF+Svo5UFU
B6yH9lYc0BuIQLx191Od3CQfNC0UgQYj5YXT29qd0xecZiGtMOmSrcbHdhVTxcr1
BlGr+gWdNtkGY60MdwkCqwl/0TzMShz/uMutCt++Db3tnnKtUpuYab12wY98tLYk
gps19v0xm2VU8zZzyt3+mtOgJr4ZSgdSaHT4DQdeW2x2/4gEtxp06TUbVvJ3WUQh
UUlxguIj6QWSvmwM3wm9a3id/FeajI+FNH4SXhLQg7S2w07w5rmCfBkphBbk5tYT
td5i2t3rTjMBP/YlQwQ1VpXdKdM0RUZ2RUKwM9KuKdUjZt1c3TjTpCpbzhLZKPSr
pC60sVmGhKoOe0RGh+ZIGgMtbwgH5eQ1HzTyvywGdLZkNyQg6O1cOqBgYvt3HGmi
q+GD6L+mp64CBu7VbmmSVTNCnFPHErrde9TYsp1WnjEYKacrYgQvfJQjGfOE93EM
r6oEj+yJtBwqy24BWxEEuCMKszZG8jK8slFmog+XqkCIAvPPKoQ1ySHlQnCq9V4B
3nI1173OV/NhDbVnMZOrTMNsC2A2U67BBm44ZEGs++B0RF2dKpdj7YFNKaFasCFP
r4HmlEViXNl40WkIxeza9CTVB/6ix7i1ZZI3tzXWXd+o99eFirB2ykL0dUbnSP34
rk+LqhQME6EpgaN5s+jGf2l45b8EI7BzHLe4SuxkYhlzXolT2Qo9dzCJCFgYmQVm
a9b+oH1BL8+DgyElemvK7flgHhmoRjrYo4t8cHNEZgodsGwcUneyW1Aj6DcoltnN
o6JjLYGO35hI7TlT/fDw5Dh3eV1wh3OeUco3SY14k2pSf8ggdBAeRapf6eBxBPxI
uLXlSBgdL43JE2mhyQSxpnO54XVHZcrmsaSlFXS26mOI99VyDpjVT0skSINdhhlP
tuy0BT8h+ZQGUrIoj87LkqRCRdbBJlF+mWWGfwpOuLr9Lqq4+GMZzFl2AMr9QfiU
GAfWGyeQQcED9e70BbA1oqR+dXr1V43tO+YQerioKyUTLzbnQbZLddNABUId30L3
UZRpde/AtYtDBDflW5MQ8Ohr6w72+nnByFZP0hkGk/IbuMkW7bIsjUWkyERUWsBj
MSJnUZ8l8hdVECwQzf4Hbn5Oha0MOLvZczVTNPieNaOlHptu+HjGDDxb5YMOxoLL
jQAb/54lHQ2EgmxHKODX0tl93FXLhC2CV8fuMqbkH3HZu6fixMTVU3Lt0NLlETs9
IrbhcgptUDQQFJI7fVVpiwA5p3rtBb+9Sl9fLsEnUHDj8isFIiN7DhJlr0rmUzWm
xSxAdZuAWmlZdKt33jaLT3GOp9FvPIE/jmE9DsvDGOpNigesRYLWyftFgzwI9MBN
tkI5BAilVu2eT7H7PrWDlLCrN2QtQYG+WA+SP6NyuRvqn7YAButjugbbG71MGYq4
VUvIovG5UUNzJmASFV5M6GprtKgRZnfJgRJxuuSOEFBVR8CtQb4D9iNHhvec6Hb4
NgzQxCLtUFx0aXin85Gx0tCM7E+PYM6ykB3uv7cGVJqGHGSfab0TL24i2VxpP0hY
iCV23OPso1GnpjZRZ/YjM5BzW4uWDgPQC10J9fAnlSvYtDmO6qBywQ0pwVMx4BhH
TgaGUeOSOmZNcolOB5vPvqIb28o1IdoagD2P4rMBCk98ivaN4iE33vwpEnxisKqU
hg3RmIeznZCcTD94MSNukCO5E/kZxNFGBEd/kETbX8gH4Ym78ZDm8+67qNEMUxuH
XBJbTq04F4Hp5t7ukK+91xJI6I0TnmJdB6F4Mk+/C0lm9V1VRmaMvqmA8nj2bbHx
JE5vmr2HEI7YerItaAu0vgj2xih3OyrSX8HgcDKel6a0N4qme92UOT8vzvxqM6vK
5+1/ImOruczCxb5XFdIzfxXappEHlRDeVL9F0qSLDmSd8NGKRjv1ho4jbE1Dv/cE
2dkQk3ujlFh14wTQZzuM8H3UBzCaDeUf7Z0pScSDtRP9HqvGCRc/ZCexlSLzOHg8
Hqbe7J3NCSclmxkw6PsVItDzrdhZfj6NA8JfHGbJoXbnQ4DtbwEtObtrDA56NHYZ
1wfUn5TWzEvwS08b/K5CFOZ+fYCmctY2rbVgT1nditAaML30gq8ckrGts6XvY1oM
FHhAhu/hoj5W5LrmupNfNZ4tsTQx1Gu2wpz9ABo3OR00KUrZjulzUh3HkLeYDC/y
0PurfvkN6DzDPlG8d/uU1EsRXV/u0TCVvhROjxEb3I7iqGzujagnRrCQPrcN3QwF
+Hl1o/ANxiFZH95XLOkUOsw2qqfytqcjc8M6q06OhE5cePyxKlf6jLkyrZ/VzT7y
PhJsbBpFOuGfb+PqoShGzJkA3hpu3NicjDt+8tm0Ka16yXMEhUZaNNAaFq8cZl6+
ypkiPyWHh4eCIVMWj3wNL8syFy2inJyL+4DLnjA/6GTCHda5gbtKyVmta6ri6Mwa
GEneNeFQl2smXtwT3f3EkeYX2D6NnvT+VF2aHsu6q2uP3pSzCQuWv8zIhIhvPnHt
odSon242OzRfhvHn5lH5NlWnLAZTPZB1SNNMuOOizzAQyvfg3nPs0RfTadQkoEzv
sROJhLoSGCq09ixzGMPpLFVCanXNRp8hfMLPgF/8YIpeEVqnbSC6S24FBIgbeZT6
mHUYhbvs/qzQmmYa8tbkI/9V4iRDWNtVR6/8eLBmyM+MxZCpg345BZUm2L1td1gj
LflcAapX+Co/l4jI/Wnv31ayg9PPZErmKYbIr/F6qvaIc3dzsvHQgas+XRWoMyHr
SG7RIxNC9ihGQkscf4YFRYEji6a3+PHjzD3nWU3tbDNmUOHweZK6eg8k8VcX4Pem
nQ2qAC1JKxvDI19eyr+RILyf+LyVZYZDDSrUWYqzkHMo4PoLPTIdg27ZjylI2t64
QXlCiTxM5SaisQX9fXCt2yXfCXdJW4RuXq0suAjQDEBcGaHR3YlD7QtiiOrg8b3O
b9aIRWtzjXUjd8ruR7bIheKwzQkzrCH6txfHhVDer30ofwA6ITqhT6swt0e4EDPY
2WNUO1o6+VYZ8MGtdM6oA2ylu9zldJWBxYAQi9owLA6RXNB717bZyTAD6TLJWiDj
tWJerqh3QpRn6A68qF6pyRrTIlSubDoT4hfAR4fjRUji+oqPBx/G+ux4lB6m6UrW
roDcdzYqpiH2rM1jx5MFBnnGnlmHZgwzGN0iPOFz1VoHOPe/T3OHGRV35lKYL2lp
Dggp8TURDNqrkMwjFzQWvVd6WSeWCSxfUYFbtEiEuMhmiM2VJaJhXitqjCAPlV0/
huNhU5bvEOIhp/PhVMEE1CUuOaVcSaKjJquEy9PLKzapR5oUA0nH8Mqas6Q6lSYh
u/iP8z85Lt8YNKr995wSmwguJPxjZRlKPJBU38Q18TTI9bujz7qxwgs6EaU4eF3Q
+peznWBOMLTnoHkrruqS8NuKpcE+UQ9cgi7UWKH2uDH9KDF7ShKRFrQKIQ0H5SPT
dPhqUJ3AQT82hcOR2oWyWno9gjPsVXui/ofzcsxPoJnjlh6U6zBJiEgqLNVqH0Hs
cdO1dpIPVYKmf2VI6cL33ccCN8eFJdBlPLwW+3da7cnbcnYvKoeY95ASjQKdPzVr
mOtiM8PsyJXLiCz/MpOD0ZSJh2tGOYLN4AkwGKwCPBfhxkgS90rOuxkKkAdvkxgt
17y3ADO4sH50qx51Xr/30/RkLYb5MkSxIxA0goc764g/E3/XW2zyMvCt6pgg5d3C
aCkyyQjbtRaMiMP76VPlfhRIaePeJAZUbLDufgU9RUCO71CXRVUd+fTIiW7yR07s
HRIDUFSE62CfzBAHE0tcXXU8snsDFboyxf8VXq/YO339HvK9mwBApPc33KbWqLwe
Bpybs/iaEKwd4PX54kumN2V1VvS/a/Id+Bm+ivhCL8G3G1I6HeSvcS7GmnKMzoVu
y8J7CoIycF3MR9DMt2oWE6D+co1qzB8GV0/USo+4cSLMX73O6R5iEfEvpiMz7YOd
Y0PMq2SgYglfzaP24yuZQ+3SvK590hjHXD66JpLQFIrgvcNz7cK1KxsjxtWJS+ju
l/JfOhiFHkzp+a48xt/TacQ1ikqtdZy5h4dRah7T63qb8HzACxgZvFasjNH3puWr
p8r8BvIBxnPPckmz1NXX3a8/S7fL3N1UGE1rmKS0oZluA57RneOytmvRP2leeR2L
cL8qzJ7U7iEMGni8RBGFSViBUC1r2i9cN/ruVcprlitcdJE1oMPZgv7kF4OzlDHc
kB0rdJFDrdjYqgKwSzq3gNRSlkk9JLcVqhn6VJZgZWJbKWJx3hm/wE7YXR39ycln
EzaLeh37IE1nxbaLWBrp9FzjpzhFjntyfLCjEIon0M4Q1mmZccQ0LtVsameYANaE
rSOGKDPsZQiM5NW8ByP2+SW1aQn+TNu4iXVpujdJMEQavwlCiUyc+M7mWU0mtghA
RM58vsvm2LJ+vLqrDiG9N+vBLkKhCXt8OOp5YQYJj+24KExMfUMpyEcZMMv/1vKk
iXDq3Rn1Efop1YM1GI2zS87aLpkgOsZlTUTQqS16b4MFJRGuCeNgSEQSSTyHDptj
robzTHmjd0nM/lxWQF24gf0KlYqPuqL/4FHy1CZ/Eoz9glqWzwgGWRHtILYYXwpP
fvq8JQVthCElErmRcGxgzPreHj76jHllZjC1E326d2AhcIude/ZelsmcaQmwXjxA
Ec4p6so2LuqcqTDMNdcD+0wqpHaOvCtXCyxq3mqBwRwGBaE2Iqzb9XvT3dzs0EOf
NWRacJ/5ex1pXwKCvqv3VY6brl3qHOpVTteHqAyqgr1Vxnb5VN1R6K36JeFcVUkl
NBcNcgW5S854ySYQzeCBe5R2K1xymVmOJ704SCVNPomD/IHYAZWI6+C0+eFbXWJy
5BzQcmYPlsVvwWyqrBHWPQM7AdXE9b02oxMtkxcXSi/+Zl9YY16FaHpbL+TUE/sP
fZimIJ9W407v2ucsRSEr6mxiaNUg4VP4qu2f0/pWA7dh9Nd8wv6b+1+pAZ7BFCrq
AStueZYwIrFyu2VOKzCaK3+nvsR6jnztoVtzEV2hw2t4F/xMWWVfV/MQ9PrY0hua
ScK/fasQ6ldS6jgvwaW7vDnKCOrMuMGrXTbEaU4j9aO4MCwatCLYqbGMz2sTD3zU
5i7hbLascWkfxs31t75Tal+BiN6/FV3/0rO82DmgF2YwhnDmSHSnWFv4uh5kC5yI
lYu7skyHYVrB0PF7NpQQ1aSzBtYS7ejqkEwOQbFv3F2zLN41ITj7pUjCSfRgzZZg
XWOUvNeL+qFk/3aSEL23LKVAHUxF42hwyRjksaDLDHwJnZtjk9PrP6f1STQSBoSe
IKzAWK4FLQeao8KJAlKC6ZuBO5+QV34lCoa0MqPN5Bj4AyFEhhM807Fgl3B2wLKT
BlQxSG2/cvWjrfv+k12W6tsGI+drQbSLvvQIhfj60kK5HUkQsQTtIHX6ydCoaa3V
/xYrTyxaVIPs4UrS9IK26MRXjDil8OD7MzfJAbqkxTZI3HgG51e+68Ac7bgTxZNr
ZIKVspW3XxdU49fTToqhs6V9ZsHuLidwbXgazI4MPEoQAzPzVCLz3ka9HSA/+8nN
vjSRUXAUjBwDgWihluLXTGAGQD/lnkt3PQZrwmejH+1NkZ9P+zePRNYysZaPJWxh
g66rsvTrSsJ2McnSFr9zVGMZ7ZCdm8frKJd6b+u3xcbqfO391N95+VJWZNKV03Yg
ZbF/v6oUR4j64op+pnEsUmntvT7BrL021EHslchpR/NXk8ZNwXhyA/cxMTtQU9hg
qyN812fuFIXFLtHxm3S9UD+4cFr/pguqo6u/F4yCDzDExxQlll6zz2Zg76CqFPpf
t76MhHUXuI/cW5TDIZEDi4V5o+f08cda7RSDDXzm7itBm/zEiD9u4Vxma5ioTCXs
3GISax10/bQVVw/kt4IpAPpNPg+d83Y/7H7JIyzZJL3sBJiuIdJRhWCQk7CWr17g
Zr9eBchs++axGiBrKI2JKZQyFpdcitNht1+vHkSOG6V1ytNaMMEzMGsKW7KhyajO
lKaktdmhoCQeE4kMlwMbJCT8/hK6I+eLba+LwHeGK5OwB9yREmyj4tOPPSNUgLZQ
ox6P3qt8GEc5TpUIs+v2+Mup3f/8TK+E4VRtCXScmcCjf3lbIjtly0YARlgl/Zjh
wavhCAvZudFBm9E/OnQkvoXQvFnsPvpSMjizGZjjVDcHhSskuXZZzepB++GUbWy9
2qL8KSeXc/Sccx3COKX+FtpQBT4D4nxOckpKterPwQUUx90ec61BbDApUXK2rjxJ
NXC8PMf+ic8/a8zhBfcQ8L1S8u7hieDvvOJ/k5f0p6Ne+p6vMzY0PL4POjeFJTZ/
CbG02DHDF8+gr7zXz75JF8ugyPrLSfy0Fv4yiLFdLSgnqaZsML1vdzD8CUl2Sk8O
6STtjvPPf2e/JQ5ErDDhMVzzSN3pQDjiaRA6APxulVbtWrObSMna5VWqgg0OoHHg
nknqw4V96DztPlLhbtzqDvAfYwj2dbWK91lA6tiMsWcsQ+enDqIyQr3yWUGMAH3V
Ez4U6SXSxzBUvAdtT/YeA36CcE0oVCQEtVahevS7LK9Qyg3aNLKaVO+jly/pyvzp
uh/HtOIvlzCykU/jiglyNPDElOxPscO3B4OeQRuEoG6zPJABbqfYKAdeBbhzUNvE
kYz18Cd68LzlTzmObjcMqR9x6hnnE7ETAHZeuobYntTbQZz54KiUc5E3YZAEXNnQ
KuMufQWVzn94aPvpgbJ3nqDMBSbcSNGt4EMxE8I5Is2GZ1NmXipCSf7HtzB1bA6a
FcLyMBFaLBASwzNAYzIFJaow5EtytAsv9do/bRKJ6g8Q2Sn2QN90WMVTi2SrY9gz
B4EVwHk2Sp4zpiNdTwaKkw/f0dQrgFysA+Ytgf64mjqouUXpHR3Gvi0K5f6p33e+
2iE6uouLdVrWYIsABv2ls/UUgmoN8//0lMXVmGfHN1c1azQ4uhz/rxrJjn30XO7K
20dyov4wNvN8YHQ9/FNJ2yDmfRGt3vwipyoYIQ+hRYbuG/zPmg1Y0jW77EEjLTD5
sXHK3D/UuqEtHoNVohfbgnFddLLlANX6Wk/Pa+xduRWerYH3lSn5CpoGbSqkPPln
esL0Xl682VCt7aGpgPDGnZsJD6/qopvGSvMnQoVZxMweyQ0c/kipOxhhZT4bdmsr
LE5Au5Wh+95/xjyQ/UZnqopOQxwxpdAKItkOMrOlscXWYRU02lPLbmXeiq1t7Ux5
fudofaZdhDLDEiEwTM6CPdCly76jCi6Vv86tPiUvrC5+EzStttm1CulsQaSV92kp
T+aki185jdaItiWrMyBJf1BncXu/EcKwJ6WNMXdb0anwSolwQlg0cp9RxrHMzwKM
cnog5TbOlwy9gJHWZTjf/HAbI5ec3YOVXgPObW4S6JRfaeP4fvWa7phLJqfhr3Do
vLimfSswq4JCtuIs/froKEhCo4jVYSnponcbeaBya8sarj1a05STydYB6uNDmvBr
6fQ9xpZ4bpbCX1zwjuj8hOlVMYZ1xnunwLUbzQLwqJSbGdwmE0WMQbzCvR13Knkv
POL8XYRam+HUPleQjfnXkdDeIvMIxQOIqIg1Fpf5qYbq82/kgwdsrGiuvzG8jrW4
P7bRGsTl6xXFca/+/yWd76VVEIo3UzZQ/9ddhDRRJVE+ALBgxw4VMkB9RaCVK78E
FsOFL25+y8HEiKx1GWq0Hs0JJYeIPISVAeDjTicEU+eJ1hGrSR4lrdve7tf7t9rg
gcBw4I5i0hO2iFiITWGCzwmmXqAUuBWYJMMqR+K2fFoAl1BskP34eomnfDQZrSvK
t11I/HBH50EVLS/abNaayITDoMl4ki5p1S6gz4p5ie8//o6gs0xKI7mmYUesW/4n
MJRybHTNVEODrIMtldkJmR8exSCkNhxCsyfaNwWAG3uF1KO9zL8X8QoxDPcxK2bb
wX28X/CGI4vGTHpW93JT8cWyLkmlWowrCd+rRE272lQji5mwgS5QTLwOvXSU2yJQ
Ks9ash7Xfrw1j/lezLCLUau/GrJtEJatIs5q/wyd9pfqP52fyCQ8q0+TzHnpoDw4
D7uVHBeaVbogii9qtq0dq4nD7apSbyZuqURn3007ovfko4k1npAZCu4sYMV1VOZz
Qp9UK9U65rCmv4j9BxsJnGb4eAINT+aKJN538NdhfUk+/zBOQBYSJ0IdiJ/QR7G+
vSjb0LAkLA590jTZ+i79Yozj9Ddp0br13phjgogRL3Cx/wSEIqu7Gf9iUuWNF+KD
j9YG/LR/QKW1W/60+lCO733FfHlIwO0w9l9r5fc1Il8YpOoRTVWgXs3IM2Ima1/+
4zMJWu5Ph5RpuujZl0aUlh9dGA7k1OAJ9Og+pxFZD2sPMbkPbm9GdQaAW7WrURul
QxqmRJVqhr9cRnFvYQZVUycBsqlYQ/VPqzotrfgF4CCpC7tHBWlzBav0OTdJtcqE
Ly2YRxtbGBw/ZPJi3dRg6pAuxiffkPmjYxXbHZturlbuanCJ2CLPfsDtRRMvUhb3
qbHuqK3/e/8AnmU4Cvl27qoy1gvuys86ypL/AKDqCgBDTKtTPY7Kon2iv/eLLp90
LNyjIgDgRJR0PfLKczt7o9LK8nd/rH+mvU29HJ2GWwC30rkhU/OmjL3UoXaKFDF+
gb4wqQi4eBWb93nRlqgVnD4qvmCRr5luTUQST5oiEc2C6blAb61NFIfHgss0sIGx
LgdTQ+8qtsA31uZm2AKDQ4yeu1DL1YKRH+H+SjO4RXTyaI1Bmkhx0rLJyh8OfyF/
KoluxxnTC2LKb605dxVMeEOIPuLg/VqYcalN6bvxvcbs04uHka/z8BcvaF07P8Ni
614rgh5SQ9ogcT/1CX0ypBsiahiZJEqWFhsSKp2Coltkzn7C64ZKpGf+OJn+WR3L
ZqcEKt8aK0zoTjCvoqT+Eu5P1SUaqetdqvHQFhDiQ68C+xmUvisjt6/nkzEnym/s
xQaxNEdKcyS3u5lnDNIzFv8i3tpfhR4Apf5/3o3F4vV9i4vBi+/RzacSh+IXpSA4
Iti8rXWIT5vbKMOYB0Gzbouo3coUPiKOl7q3amqXNwuTbnQNmaAZeZT5/+ruCAve
3rQgKdcNi9oGyMYVWUwy0vMc7p88kDKdtSFBx+DEpIprilzwDKkYAOU/vjzb9UWQ
XZzIUeDgG3tZb92/3DpZ7B7Er8fukPySK6URY353+qDIPcylm52OG+GAn6rdHmL+
EacGxYLLuIFoDUz6SiGtBu4fQfwWKvewP/gtjzRFBE3qxu574haLi1vgIpEpILDK
nVoQvI7szpDLcBjb3KddrbAWncJl0tqMyx9B77qEflR98dk3mhULeG/G51zh8W42
RFqXxwXOZm6MD3rtMNPg8kwtud3SQQRdBbJT5OVnhv+5yBzPME21p4/1IyBRuJBQ
Ixo1DCbjGMwq41sEwhVzDnCyf86ibhM0MUKvmaKB7Fs4sWvaBWYoS6+BnvnjFtOC
RMis4KjITLdW8fzEZ7wBb5RkJ71yZc7oHxsScLKQDNaG5DylpXtF6MnZeGqUj/iu
x54b9WnqfpqW8Za+Az954Mu9W/KQbpTWUzPSj5o6UPKCbt3Wpge6FqLk+t4pv3xC
bO67UkUHH1wpvWsiUNrNoZEOYvab5tL8/bbpH2890G4D54pDhd9Cv9M7m6+PP96j
mUerX4TF/boV6AWWaLqURvdjgrO2uEmCztpO2PI4qocprqrem9qNKe03ftMBwWN+
cS+lssVvBM6PLOSrbBwIRsoc6BajVS2VQ5Z14RJnZ8TH9cKOwr8F49CU6/7oZaV0
IXl75lIacif5vFP/5+CcSN0xGIm5kuIBPf3n438oHyc5HWaoSEVLV0EKdDDE0dKp
HPe50Y/XCXuGX4+YP3evdAz5x3QXaXp/XntbT3uoB1197J/HmjQHkh3frfgGjwFR
Uu1jyHjRYOgnXXpM1G0ZwIDa8bN3ABJqCeDA/8+EDom2MP/uN6/E56yMkXIepQGr
jblvJHSaTL0dUqoyLMvOYjTV2WK/puv6KdILRoHhGJ+4UPLSMisSYru8sNgPxstF
OhOXgU6ZC1wFae/4Tg/mn/9DbhQO7IxUVVpAFWGCM1W0BV1J5N2ricSgg0szy+3l
HGysvxmQNEcJ13J0UsQmAnG4hNKrOAh5Oq9jNBLHiZ/u/+T8P5iO45CF48cxKny3
LyEjbXgELYzV9dgfxvt8zO9QUcb/sYA+EjnczPdzqpqJlRQRrr+ehC5YlnGieXha
CjWXgRb/yc57c2Flbuj60TAT560mzUfZtvcXOCcmmD/Hl5qs9ywhy5vpFOSFGIQO
FJn9SVwv8iFjk1sa4URGYDHPLx00Z5mxlEjEyCbfpfedHo3DzUVAeBaFZZypEeFB
sgIN0/fYAiOW386wSoekKdEWPrDZHziwprqTK2mwgsW7h+M0053IAS3aTIlgoxkw
/MIDGKj0E1Drw6Y/OPDSPbv5TI2xC/Z5jqEpuGQkyhmohE/98T4dqrs/QoZcmVZ/
9IDxWs47lo3eKCIApSOQm2f3TUwVP6wmrGs9U7RGaphGUii59lPZNmt4U16q82v4
7rxzmMcNL1vrn5ZrTBSfKynuClpGRLT5vurbVE7C7Vi3v2SHhWTwTdwC7gFMBA8L
p/GrUURDAhs883tDvtUtxY1wtRvnaCnYrpWC26dQ9qv7sLLgjiDE2Qy7wGZHjmyI
LFMWkC2YanDKs9VJmAdFAuNr3bkSjQde3Hs6jIGPagkHE6c7CYQjGcihOgZs0TDn
kmg76UDhv1pUeJFX7B0XeL9evkBlsPasz/BpXqBb2JH5XRhINsutfCsrVm2vUzi5
kZXrUd3JohBBr8CrNpEB76qs2lsxH9M69omG81ytoCqAmdGEiqtblHxTLs1I4UQk
O4e8iISrnnemHAlN3CpG13IZYIkBPPm2IAgaQcDWecbM81xV9mTcylzWFdYOchzW
Y0jgM1CDhYfSf7lhGBkODd74iT5vF1iGNotRUeewbhCu2FvxzA7zE/kcB6APTIyv
G+Sb0rgS6TeoWP0Wj6DnjLkv8Rke9hrXlsTQ+zGnGShvNDx3v4Xv4a9WY4p0/J36
WPJwHZe+I/5NCgaKsyKWM8Gr1lEB641D+JGukp0kEQwbMg0t0SIkBbryHqLAxlRC
/Wf672fDADSouKycqsl/CI8iY+Enw+Ej72yY5zaABocPFbctYYctD1RysZAFmX1R
XtYiz0tcn6J2Jn6lk2c/gdWvgqGGxuvf0sAKfzERW441Q5zE8vycdnwj+9PwMjmt
Dvd+KcsDfbR5LsBnKDwv4LhjNcj0guKPWoNx4e2MVfsEbS3n3ji5OEgHRktmo4ZS
qgZg9aYpNn/5ZDMm/hthbPSmHvtDRMyQxGRVLhj5Gnj57QIkZRjYQR+Xh/gzmT8E
jWaFZ6YJF9yljVjyZ9O3C/9kaM4NgvoYajCluyVtbL7kr8iatvQXe1Z7KeqHoT+J
H5jCFmj8Q4UvLZYFlWD91A5E+ORD2Xd5R1/vc384UavX4D4hZ3MeRyi537IiE0yS
Kbszfp+SptP+VerwzZB7dt1Uwe+SJht3g37CKCIO7f0/4fwBWOHB732sczr2pyKf
jdgUmh3KLKEStsTuFaxqTd692g+MDHHmC4to4CfHB1rNlK62BcK+JlkvAGCio8Q8
dtsuDPVsGxPSxZz2tovFoQwq3hs0zl0thKT9ZyiklHNel6l+N1SF15wFXvasmF75
mX1pLhdhQdFyxBrVN3/DaMDaNRbfekTSDyc/e4ccpqpvpLncORLN2Pj9G04mHPYg
BD7tLhLCxLb/UtVr7pRKzEJRu6GcSrsci/y5Vy1k6v/+JOVuiG0K4qOAFN8C/hYV
lvr4YXp827QIt/Nhk6P59F8GZv/SBg4Pn2B28hdMyjj2bummbmIiO8zG8N77gBjb
zQZP6uxdXk46X1OfNioVOHn+FUt8Mf/He3MMtgTdMznzW+HrhSD7pxaTbjWjLVf2
oL48OsKFEt9oecfG3pS9O0fu+hkNwTJ80eW9MWyzSsYQrwHdKVm9fGwHPkGrGJI7
O5HdvdCkFJMDGItTz2wCGX87rVU6J8xdFGCvzR/1pWPChDFFaMOUSbyA+7Y1Vf20
SFu5mVSTW9fmV3Kc1OFzk827ADwJfzm4bQTCRyNCU2MKahJ50pZgHkzhb2UJVLvx
P9XYcR+rwuTqwJFAbfvJb0N8LomY5NniKZ1dnzQsJGIxngnDjGdZ5IIwIlL6KvfL
O22b4Ad8JECWArE3cTlTu3vEJc0CpoRM2UrRVA8tWlrwczcCfVrnyXUugXmvLKGK
StrARNfm9IRLRYV9qjgmEWO6jQqWHG/t8Wyy3zwIhB3s9SBIbaZtzrC2ZwstgVcP
gc4YQ1jbt4o71WM8llTlVdzyfwrdflcaCFbGa2m5fDxe/DGW/n+2ORROSGMmpWQg
J5QxB00k970vBHZagBz0U+M95GjwoVJSoLUVRBK+u8JoomDkW3PLPdmIwT05JWbJ
Qe36yfzOTQ7wIjeKvt5kwvG6lHQKSQdAtJBMyt9TRL20ET0zj+NvRWvRyIB5TI1I
ZhRgxkd5UQzBHugPM6LpVJKhMQYqLvMCIBRnxM8z/zPjAltoT1NiqGWODlra3RSI
mAdLzuO7U0+zusHv8TUtyiqcP4HfkDEEXH72AyvFWX5p0/MxsEoJsydi3GLU/vTt
/lEWaGFgq447cR7+BQRozSoBznpxRZzNZxflBlnhP6EyUTIYJMJRDEVoMsA/gjOt
V4jLves9iB5SOp255hCtjKAcFcVuDI8Evqnr4o/sO3LUAMziYSnZqhR1MJ95IqkA
taqteM0JLlPgctHX7mTE7NauMcvDJhJwvQ5Brooqav79OX8rPP35/IUXI5HPS83S
ohOzhIFCRXdqpHTzcLvkrqNNc1Xdt+AwtT8Utj+yGLRILHfNQ1SUSYRVdCm/aggQ
AJzl9MxB7BARSXitkhB+uA3RYFFSY0bBjZ/eNXBqEdTyWSdCINpZFVzCX5GIrFxc
O93y/wRYryJ8c5wtM3RHrbI6a6SFUQci1udJmeF17p/4i9crLogGaj6RZy8FXt5p
2NShH1tvvYRTu6CkVnDbFBQt87lAqlMlbneWbBSL8lCCrnEZI6TmiceeIcw87sHF
qjSlqnzRT1Jxcvn77gm5xIDD7SyZlLQsnpKzBO1Hc5jWuNOC4lg+HJOZf4xTYl5k
1jjGcV0WmdPgqzN2epCvfapCtOYeHwkMco9NVHSVI5lEafBiaU4gk2L2DU/Tca7A
2qw8gYg1RX4mPCr93a3KDGz1Rr+wzSwewE9DSLGgYUJcZzQ7ebJlEO6h+oYUvt3i
4eLWJh7qXBsThSkBdqbjWKJtdJzMZdRKxzYc7Z5zCkpfHD8VIGfKBs+MiSfMKcGZ
0O5jXKmQgwokL1ZZqhHWcXPff+Tb88Y1f30Om3GScd29d3xLc/VFzgYNrq71n6N9
HghYJF0QgkyrN/54b9tz/NfTFe57L3+7lxEnmy6ckLja8/WpWbzAt38P9Iy3bLTs
pmRAM9jeZynEDEckVyJncJtNfiJAWmKeMDHB4vHzFNXvvZzM1yA+0JY1KYWrXJAa
JE5UUTT3baqLpql/EWFggnykZoLB201MYyhdnKnk/qezvBRZfM9gcWV4uOeWAwTP
ceKJuG8H5VSRZQIZR/OsYETCO+U3KSECl9gh8ZFPg0N6dLDAlENidxVrmaork+j8
IHq+aVk1VnOOGH0dIuzHvkM+kH9S+sJyWBowmd8GodYCkxMjswvFsr4EZY0DelHw
0GE4zqy+YjCyAw7j2K1hCJGyed2wA5/AR7iKtLFYCPN6yivaJ7Sp3hezCdUS3xXO
h89yF03rXb4CR32/s7kCDhlV/HRHmH/EXvkIfwe07jptN2Xqx2q0s76WJlNbIa6O
OJHkEJsX3BmcjnijsS3eRcheHxdht4xuslNJ2zng8AMuBx77gsuDAH6XBEFQ/yRb
j4odlZEhBgdCJ3zrvu6JhUe4zGb9tfHFZLGhKL7m0MGNnNntxuKl3au62vTgRGeK
YCllFX/zosrXjIpSbPAWKltbgVXc+wBMrXb3TadhjVW/93Tk+iSPB6EL0HGYFzse
zNV+PglhxI1HfU1eLOzI5phBmNspPQcdcxbroiRGrys/NdWmz1Hr+cUD1WeklGV/
lcm9P1lY8y+suO2v5OyY9Yr3saJYOErThxvx4LAWmBt6uXaEj+/rl1gfo5tZ7cHJ
wl28UPo+bUX3BwWQSFOyqUIAX2KVAkK61An5Niyd8s+njDW5/Nfb6aeM13ipZP9E
Zz44teYLTZfhX5AD0V3QJflZiVIz8kuP/NYAP3HcT1qTTV3ty3T6oNnzQuLOiFCi
qWSmYfGZtICqIkzmFJ2ZQLpqseiNlxbTyOP6sQX36u0YaOK6PFfT+0kS9xG+Je/7
a6t08uD9dgGWEh5YXe4jzgYWo8EwwCfLbs9ikEzH2OfbiiM+OAPxBHekoOKe0YtJ
6UyzbzPCgW0nQjlb+czD8CUv9hQtNJtQ9uS7ZN06GZW44HQrmIBQlTiujkTOIJty
dGjLEXDKeqoX2WhT9EDTAg3HhM1rUmQc2GrJEiufOoaniV6zgOc8RtBl0b5vuQVR
DDPrivdemZHBF/BfdZB8FIuyga72U7g6N/Ph54Iug9fo83tBLLAAG2qqLcVjUxs8
pBFYnMtMEU4/ZK2jmT1oCFATInGd0eq7VndKA78VlkLmGRORghenLViwrRYiNLOZ
61XYOhBy2rAeRrXnzLCPSBi8OrXPwIiJ5/JIecRHIA+5uj0ge9CLHn3s4bYB4ceO
ONMNt1kex/Bb75kx69O1b5ma2QSacPJn8zyTr1xTDGRh4x5Bw80l9DqVFNqNdztH
B7VFY1OxtyKVeGZb5ZQSaHsaTzbS8KvznYOYMrVRAAq0r5AiF9iXgTe3J3F+ATxI
L268b7mm0oBbJaBb5CWoAuRTRSViWa6rC2LnkBYHIuL9v/XvLCvUjEfGJYEgdLzI
0GDopJj+Hh4OIYV+UDaegregoKB4JA3uOY7mqipAlPqvl+VCD4QVr0QejVxaeHxx
aG+cle7Y3yiRD/CGZpFfe2+q061E5dvwcHCaeuY+LdE7Ih0Ca4dDiYpGysQxB3x+
KsfWYDiUzQz912JKmvKwIHuDsQJI9huLpUPCKeEU5GsjIzYHNl2AiqWYOhCR05Qx
QOAchj7c3rhMacGfrynADP8yeYW6k9M6VhXC6VzaletzW4KO0iCk2WVyj8KdMFRv
DuboZp2P6tkWGWK1y5ThtmUijx0dbi9gwkeHHVk2Hz4VIJ5ieb1U13WOdCCFNBC4
SmK7x7hHQxrdoBij7YtKCf96f9JKkHNaJXHTFVJUKxIc+tTBa38dQ6WADouhrQdZ
L/Z3uDru4HA5Hddve3SRXFTah6vDCKTomqE+yNKTdq2U/efuGysYvRm67FJX6csv
gMzz6p/pDsp7jlaARrvUYwrg2cCNUqVP2qg9tlWtb50uh+yJDT2g+wZHZi/7siKa
QtJVFoapVro6Za3tZhEzisCXVDdkWXHsJf1jWm+PQVUhEJu0Zbb+JSeHPs5XSfbb
UfFxHasEDyCtEeZFRxdMcnZUa9H+EIhjtIP2uzKK5jiMqQ6C5hHzAbX1hA9dw4k3
M9iLf0mQOaQXoV8k3Px3LEDeLBy8HtLYxQT/iaFtfqrogmafNUUcqPABF68sqPRp
IXrwHX8Ibx8APIxbHs89WX3bbhnm/MmssMBXdt0Z/l++JFKWgpooMcHYOrFYymLr
C04fIcdmoogtwc3M7Ge5GO/YoJXX64k+2sgoQTlA7Uf27ueZPU2RDFx+ztOWuIrw
Wy2OAlLLgge8j2pdYvrmqCXq3XCmq+Z+S9UT2zLpndF5GQok4YyfgkbVr+DSRoBm
WE5uo3h3Yg1GBIkt7YS+iOUvzNonS5LIA3tE8+TSSeKJ95/3VnyMYxOv5saOq8N+
5Yf1KyVEuPfqvKQ8Ogp9PZrhx7iWZ1Ir3OdtzYhmEDtTImokaliN/Q5ABaaTLhPA
7e38CZW/A3+hQJBfLZjxGtkm0or6/4C2urKWY2fuKoh1ynJ/m+MifhhNIs3MyzOu
XdAog6mWU7ljxvRTf8m15OEb75+5Lb0t+mKQSkiegcwwm5H3ts0e4ES+UuhEfKmn
N0NPKGZ5yvGMiUOZA/IF3DNCWkGpYVhkFBxv9ipJ2GsIM4ea5V6wKQuqUFJtJfhB
NBhxVxOz+LyKYVtwoenp2zytJgegT4tvUzEnzFPT9bUxndx1kIGvSVI2SvTbiReT
h423eVM3AhaacXE8vVz+v7ah6V4XjbUBU+MUBEKJZTXIIf3OC87lPCUSltBzk2BQ
LYyt3iKUZbGfiMR2fsJL5Rgacz0/WdKDqfSUEcTXbkISiBn4Vs7+OdXaCXslLNnf
hdHjyAJqlhHu37MWiXxGpJnaWgghUrXp+wV2wQ4fV5Z42mRIX/1kmqJA+1H7DwFG
3gU8iWTLL2qtRojrjKa8L4lWmHkJifkDlB5DS4KiemCUrse8HXplWVn6CEVdDXGs
P0U92c9MngYXV2tXz6jYwmD4U/XuM+LTIY7kMRVyzNk4zOcKyy/bAmURdkzg7OnJ
zjSbcFyuQ6U6AQ5pyQG0zGe5UTmyTnnB9FugVJCB6yos+z+9aOBXKIkCpB2SbNNC
PLtNbEim2YPJgZqp9fD2rHf6yFQJpkaQGy683WJDhWlOsf+zY1nEaeqXmaqXPze9
mV6e0mwN2Xec/23bhHoJ9t2Aaeep3iuu0DNuQLuNm/CpLFMBFmdHhnmXVdQoQm6E
GKCRUPxr8mBQHNG7wfeSZKoddqSqL1P86U0jRkrismzPW/0WSS7rfSQ2HJmeIra/
xCtAGKWFmTObwTwCDzHr41KpACQ2CVCykfcxTwUt8byPDfVSQMgn72EroKio71Mi
gv2PC4oxy8a0Ftf3mp8ZTDqy6ls+U6va5EZKyyG9pUVA1nSAA0uwMFgJJqJvSVuw
+LlbS1SIJv+WHN+AsvECqCwXSlI50qZpCSGJWckv+npxl74tRf7ufvxFNJrdXI9r
lyIt/35XcJ6ErgUxubc3KJsmfl4h8C6b6BlWX4mzLaKKTzvXpk0ZFB7JktS5Pi2O
uzN32j1cH6Wqjs4f3zad2wOwgoY/cc0AYppCD1p1BPRsC7dqy3/zeW6O4Nqm9iwj
hKtme3Sx2tuNVBw7FxR3unsIXiKUnIu2izvPMYIVpQxKeFKy8TTfFUK7yQmY/4Nc
ZFMbsMai0+nXYdZIVIRbX0ef6fOGNlWjl7Dp23D1IqOI29FHXC+awzGIvzYaA54E
pXM1fNt6wxJ3GQrxmxn1hIdKwv7bOvsqNHNAN3k2eh0hJplEBoQTdE11a4TaCvKo
1wEe9bOPveW1KOegezYJv7uAqftswbHQNSHQdHvw/XM0gcs1Pp341qRvq06SxhH0
LiZaoOQZ2luKY4lnBOcUfGRz9xOMQCcogZ5zKAjaltvUEDxj+UDhmUr7zyhQEiR+
fW99tpcm6MIskh8PV/X/nx6pATCgyzCIXHke06hquGGzuK7tPerG6D/pkAYgWld7
IIrO2Zm604gCNNI2ZGAGhp6xTYpTQIb3HSgeSNk7R1m7VCiixc4ITzSg4OBIt6Nn
XWLD2cmai0Jtr5WQphI2rAHgr+ih/1Eyui/nuS7MzfuvqRuvVL3YrpoZRTamUSX4
W0la8L9LO0hPS40G1r3zZjYw41AbQMyBXyeSaovBYBBBKtFeaywRHlRre40kE7B8
al37WVj4w3FF1bUk2hMZjgSibxaiXrwKIcpWQjxynxTgY3hu1Ibx8/gtTp9tD0jN
OzSLtQx0qW3oKVsbPrk2+aISmywRND0BU+10D13ExbH3P+07Cb7Th2gCrc+KIMOQ
XSl6+N64ZkC57HMzDQW0d3Kne2h1e4ViNaFRyDMHrsJuwz4Av05LHtttnzZwD4IQ
5B3sYXS1zEi6J6Vg0FZ88kiTnT7vUGNGnIuTym5t69pweKE7UwMOqbHdEDktK6xn
kCSWoyuYQN6lhq9gDBgpmGrjr/dkcx3qeI1a/eHkHfLFZwK+2wcj9rBw+9Xt5b31
Pk7K4F83bn6QsqkYgrmU6/eOOVhyzPd//fn448OqfLVNZ+UcMDuJbY/2KvY6UISI
RorZ0Lc91B3ifURvezkY0SzgrjfUkZBlf6yX5XfhH9gN3oLFZsWAmxPyXEpFEsik
w4Pl6kP18zw6zQsAFlIcg3UvmltDLrUxEu3vcHClUitPoA4AO3UNLEeA6iD5Pw+5
c4K7o6ztxSo8ZEGi0QkntyDJZrQOw/UcQwMq/PEMtKP1aiDilb8WSAP/BzpR87ya
S+HjZO9g1rql2ec06WCr0jQgj3yUAANriwZSCwJGB3VjjOiGuhgopaMk3d/E/0cy
xEs6oPlJO9JAUY5uuoMBnN7MtsSRBxSDL3QxnVepp5xRgOdy9G9BtU5Apdk4Fike
nWsKlKNDdofqgifGrHoQZgAe6CViTgckALaAbkW/BDrukwINb0xEPiQxMD5hV9L3
rae8CTxKH2DL/R3kjZ2iKkxrgPWaAV2gbVD+HOixpW1vaCpxhfPCtLgIIw8g8dY7
6RD5P978XRLUnYyN3FEtod4zPGA3FfLbA+Br+z7EK/s7M4iqmjX4SFVQzhdiB+QD
VEVMXNGyACRPnJXaZOcpi8IgLCjdnT5GpEvt8ftrqfqJ5ZWg4Ap4mJ0k1cOgE8+S
zFIZblocj+8aYejqSWGSbzwmh5N1dbtlLOGPlBNEY35kiR5KDQZDsAoc61TnlsHM
j7DP3gHXkHOGYGkwq7qUPJ9uwrmFFEGbmdjGc/xIc64DdcAndXMzA5QuqiqNNP69
+chDbQfO4Mi4TkExEDHo3miTtUWqS+62NAeJutepMCweesMQmBL6WjW883c9sddC
mpHqsFeW8TFlaU+hDUvPN7Ta0GQGWsQnRmMqjMuJmfX+NkeZNpXZB3xgOgMXkqKC
F8SPzLpoLG0m0vdZs76ZUQjHr2Y4MIichmepe85uKA4TlVveGx7FfuRlnEpRxxqi
4KInPkzcXiU6XKRUVTi1MlqLOVV+mvBgcWXySA/u/OgfzjRWxncahAkTkKI38RkS
zl8KyStjlCgj3N75F7c7Ni1sY1FBlco5ZkK72pAWpcRKmI4Fyc3UViyekFn+2gNL
tZLe2MRIUpydBFfnvcFKBrF0XzdK3pBzlpLV025bQ9ROUTPIprsHownktS/qQyPQ
ue3SgxXYWBesjI/DBv9S7F1ED8CP9kR+sSSpq+DPL3HC1EWaif1XfI5Pjj0xkWZd
amI+Rq+4bVCyNykc/tim91X6TW+xexyof/uGOiI+jfIICjNBtZ7lxEHpVQzzIVbC
b/I0qQQjDizXw85QhB46qSzLeDPUeZvj0I76co9XJel7inJ/ofNB4CnMS9sagcRb
Q2U34q/OHfTj1mSmkV0R//Y2rfRDF/ItkMMadVXmX5kkeQhjXX6HezE7eORbjXZc
nMWHuYQ0wNEhCV54Z3abEXHgwZtgY+mrRo1jrJgw4oLE9TksNAWgHhdSIWTG7TWk
yfGPFSff3tnzb1fhHACkET8tkMXuNbv8Elhe8UmyYJ0SR5W6himKiQbqNbsjf94j
MKMW0gZuhBX6BajcQ4s69rM7DiGClThAyc0aRMQvpbSn5Of7Vg7PKM2p4+Iyo4yE
V6kJ+C3AUXkShiGamaPw29auMJdXeQ8RiAZOTZoNNnGhATXiHur+0G2RrHOkoGvB
pZ9x61lb0CdU4EUx0nh4NmZst0U+dv8ueotv6yCRB+tGBtVHIlTDFSzVmo+LIUMN
7g/W6NFfDJSzToyhZxE8IEV9IcOqGb/dWy/9n5HwBcfTjpBQgU4qKMWI9tc2aMxa
J4NN9LhsG+qKlBGwyCQTHne60sDcOxyaY6MPaGNJ5MFQAUkwSnw9XzsF+9kC91v9
iaUi3BssYcjtbhgsuo+5pshkAojrir/Fua8wgEIDdNHJd6yNZJySVcnrGoKWX275
BICGnOnTwukBJhUcyVOxSqGNoKKdENdEa0GtbHEMsrrNeaR/yKTvu8Cr9SWbkkIU
sTKJkCgDffAVV9bkpUv3BTcUFkP7Tqt+VMIqUSJzzl8C0E6CZopHDoqwtFfXZrs7
/bIoXEwws8ADB1xNCnAiVsx0cz7UgS/FcB0S5qr/Pcb4dv8cTmP+gH5AYbIJP7KV
1Y77I/WP0k8vZtxbWFZCAAh1f+z4AdcaEZHsFHcTFYuaB+RslDiaKrKtwgr1+rCh
6feJqvz5UcQTtdAQ6oXUnAq4pL/KYPLk9FrL3N3cI9UaHkZL3JMomev5GK7XVOxs
3zwZPJWYWY3jwYL1UDkSb6liq137SwHD0QlMel2dWFoBoIB7OCJfELdmYgTK3hpr
7xA3Y774zBQuII25s0xinfgJMbcY83Li9u86gLlsi7Vg7DTUqni4lMbDaoyet0sz
Jgb8numdE8UzjWn4Imzz4FwiCIvxg9nODDdJTztL7u5u0vryTTk3nOKIxX+NXv2j
rga40+j0Th1/wDso8ZOxg86kSsImrR9zZxGqhbdGShtRbOdPJ/Bape+sGz8AnvnK
IDbVuiqSSspld1uzCnSGYr/g1UL2QfvWvq0S/bzuun+tuhhxUbMh0Hej00JbLomL
q7g2jxdiA1kzZTJlu5rC/G89OiTO/DemraNoY/53t6MRS1brmmH0/htUyEACJaeB
82YfVXJqFaI3eAWAyljzADmPjoeEwQWQ9a8+GzgFcBljkKauHgdMs9Oz5JT49ayD
E8uiO8qIQAd6F3bLzrIdFAWCQ5lYDq4H3kU9UColzmpHOIbL6cNrBwlPdbLqIvVY
cUII5biWRzk1UPghRCncnFnaWq2iA7Itdj45Jgh2BpBHK74n3bRh+eqCHWDQkHJS
2DySCPpyf56YD2enDiPq/6oE3hvv4jo6rwRDGTaPiY5jjKmhlv3wkg9PFIxC6PdN
hlBSw5O3dnaRdckJxoyuP+djKXnrTDXA3IR19ciCoQ2iXrFa2N2qfKud2tdg3E4f
0VeVRdvXXv5bwi3bkn/hpi63S/D7WjYMKQD6vWraEM8kT81LZ8+5cw4U7XWmlrxO
iheXlPmWk0nu/KfQZjcVkAnyXX/2Ba2bjOMCmooVcFKbyKglZ6YeDUSzM5jm5rCD
U9q9YzPRZ+ij6GTnD8yRx6RfLKTCIFPYK3DaAu9s7Cp4btLnaduN8qJTJTmSc2uj
MnoxU+/Zc1ov0tClKRNj3xQfB01Gsrc/oA3wIf/SX2r+icpEuqSRZrK2o/0zJ/b7
NJQTI30R1Ql4sjtUwVAbCpEuw9kxskWI70HcVK3ifjuwSSFhYtug53GGshV8nohW
EjCFiJPDzzSv5KpaEEYTZsoJQ2R14EhGpLsJSSIam7lrx6ZpSiFVm8YNDnR1NbLO
NLqWhEkG2yjv9QgoedKdTPkQaGgIM2Sr1aeq/djsUyxMRw/J3H9Xf5q/+Z9EjTk5
VSktMk9iBPGkKjb0meP7UqFI754be+Pna2lbXMwNxHi+r0aN9Sl3I9soxZODR6a0
qfMbnmCP6QVUsJOt9CRuhz/24awRZiDgXxDmmJ8iCmf93Vz1hc9SeMMlbMW6TTI+
EEwN/zXKRJzwzmdx3kfTmAMgdk+TXhqTt7cA783VEE/vzkOQgt+jkWOgeLEYX0Db
YbJv4O1JO1DE29lZRZakjLrBP11nIqQ469BigECrh0XBaJ5XrNE58HhOzVRo0MUt
k38hxWCEd1EBm5Y3a1KN25jhKmvZ6NQkzjK7wPxOXK0bP331QhzJbyRkSFEJkDOo
puCHdGAJ6Mj5aaRakCc699c0ju4ztfSs9nsz2JJhkWApenRlC2sWuirW0Vuj6UIu
DgkAGdkKPzPIRIT/BUD7U2f1/BaknQlu3h6Njca5lw6/vBosw53eUtM2oQDWvLTy
fuz+chhkwwRR6ff7tRMx2BP16tyMQ5bucZotOx0JYpg+N56LTHIEAmVkp1JTyi1I
X8oKeql6CXvawsueZB+Ib/r/yvpLnqgbw/7DLTMrGWGspSxsnvG9CAgrUTtxqgxI
0TWbJmkYKLBf7o5J28SCCJqXfbtuqh7ipxhzyoqc/M4WXr6PDlC3wzFgVACPkmwl
045Rad1w2RgPC2hsxFdUGLkYKJ7Jg91Q9v+lo2ImDuy4N2k3p01wOwdKv8lQVZT/
WFIwsWibX/II/vuy73+jGYrOFzs9HASkur83+/5WhGi2qC4djl/5mnaL/qDJ681v
bjhUD07MhIbkqMMPwjym5hBJMK6w28/CTll/UL6V5RqltdJpcPZoD0c+AEfRYf//
tozk+446cbzJOfjmvoGK3UiqzR//BplJx89vQ8la1Fx4ODHhEOlYxfnF+wI91Qqb
ak9SfLCMJao+qBCIq/YuL89cMzsHc6TD1jhGztToE9SY3BHMsq2nyUKZTvN0OWbl
vYkrHDEaDOs2ebiJ8XF20k7d6CMuc12jM/BwvMHJgMR4Hoy6WIbn5gTHDFMEqqEP
bh8l78g17pEqJCvvJKfLpMRqI8QgtAPO/9nwI4FtGm2vShZSaYj38pTzvERHqdrl
ChAJgEY62QUK13pDzZAZUkcma6dRZqwGnJauh7ZKIJZIdL+Tc0o4Yvc3JaLi84w/
C1Nf9PLZn44vLu2cHnWvjlfmhHlXpW4jF2GUF1gMv6ueJ6HDYym/ddm/Fc5YjATW
Lf9iwI+9Fj/QRrelj75aEOB3D1QEq7jWTNgv5KTS86BC4DXc0ePVuwHQBMdQGsm/
6ENfO4fxj9TCf6wDaCaBbgA/a9AgCFFqQy3HebmTi6DZUHYtWbwJsELjQwbCU4sc
0Q8tifkzeRUdKCZ/XuCshmEN/DT7icT93eULlfVSWI6rT4AOGb+wEpzwuqxWc21K
yT/0w1J7NFbPtsiHwAXf2g+OsKIrZ07J5ViLRmj88pL5Uym6oN+FZGeQgr1R8Ejc
e4XLvADa5S3DmCi0LynxW0WbVA8OzoF4/vKEZcUc0PZjPw+l05PQdSkR7LA5Q9/C
HW2ke6KrD6dkI2pyMERJIIUI9JTS1T2MQLmMdIhgXJ0o3wkMLFKTcBDRLzaT43aP
+pw2BzKi1n6fRh2RcReveci7//iDD6Qi9wsyQbcWi35b5lpVXDdbHTVK/j+4SANM
hJZgJjKIBoSprYX0kc3dy6itfNkLSDnvlPC0/PQVIPlDdhWRLU0QIwse+jV487FI
evSj2PWwWAzfUZgXJFwV3hNIoWjxe+pql28WusJjNYZhv6uHYvyhjKzHYQvuOKZL
WD4BggurBB9N18dK8k4+aBDFJRLiHAyJlGI9Oo+7Fj0wm7RqFIqLRW3DurB/5108
LeJBHWFNityOqBWXglsIIQdSKGaYUdJeUhdSX/HWjJLvvA/QbVjDHzzs7NFVOL89
NUGRfBm1gjzPclEnSc/UW3sUg0/WwjoNzMK44WW9iJaqUR8pKmlHUcOuXEnXRXjs
/ovgmYUoPPEEQRrG9uKC14C1aIypc7Om3TPo7KYICBoDICazlALQ6TV5Pp9hGyBd
1y7SunU3B1q2MwE0+Ffz4iTiLilJ9O7OfeDiZuwdUFAVowKbsMM/a1/1n4XgsWD0
1sVqNNx235mfVKTRjJowMJRby7S+CjjkNjhYOXixg2DYneD50EO4vsiK8GkmBNK7
pZ6jqi3biWhjYNWPJajLMEkkr6h20O/DZibWb36YYH8aF2gRNph79oJGRwlq7tKl
vs3T+E+zQZ+nluClUDB9VaZCDJNXvFM4y1prWAAZupyyGf9SQQPK+6ADDuKKuazj
WZZlBNhIlzRIxYQ65iQpKl2XCG7k4ykOCWIWPAISocG5bJKwkbc9FegGRufuqgKJ
6g35VmauEx40eOO4bVz2JdgMv+x2nguPMFOx+0uGAZyOejId5A0huRJAqPNr2gmb
ftCUNUFzBeVULRxi9X6s2kMe6hU0/wtMx1zwj7ms6Sd78NtLYK9nhNtvSVET2pNO
AfjHiBFkGGFMQNqWKtxaqwnyrMp5jmbVKT5OD53NJkiCNEeZLgqmPAJ+G15EUQFJ
+UMciqDH90t7KiN7sDJMtBuALX8vzPysGSKhMiDfx/QDin/MGUP5+aXfOgRQYcQ2
0KUEr/VFEfoF8QVJCOng6ryOA1RG8IXi2L8u2HmALXjQ9ZkkAlGlkkNfsiWTCjpp
ABsJpQKwWxNI1L71WP9vrVK6HInX6m/Ii5AErFPhKdnIlYgE0HZ9hdL7g4QeryL6
SyCO9HWEtvqZpojVDKDn3l4KuS8lz+THovrigQq6+0o9yQk6N4vJ6wqBLSKEHcWD
BroIm1FxICkaizXdQAVgY58tt756QnkCr3RnxO52uBGaY+z5zyM0OtZt3Ecd+3XY
CilMehvvwejEeOvjobZmhjWdPenp3Q4cXHea9u13ZCQSIKzZ3re/ABQ/JXkTiuFK
wODeSWziAXLTKP29eMOs9odAvgr0H/qKywMpU5MfM4UrP+6ntYQe0LYxD6LuEP3d
WCbCHpfhrBihVOiSNlcW+It06vqQOWXKup+/xhfdclW+kdt71Sn3o5d+vTR9x17v
EyABMpQ3OZ2tAa0AqC8+GWCKNCVxo46w0/6i4+rwpp2IW1PBI+FfWTsQORWX9hup
elCwGhDrwmXsV890uHhqv4MHhBwdpP5ipj6Cj1pjJn9cEAvJiHH0a8qgssEBBQ1x
Z9O01lsITrf9OKFWldVPvgZiWwPQrO7+b45tScxEFw+yIOW5MD25KFeZmHNrqNg7
SVdHmTNqKnUrurYqj/ap3GVg7EIug4WmFR4gibwXVk3ck7q8K7jJE6JvrUl1HkN+
nonL41EvFBH15ONXcBL5/oPlQwGqLff6/DEKZcf+rX9c9jUfEp6i7vif8cZmKmbF
WelHK+igwbSk9wCR99b9c6UBrsL1jLDGH7jxY8D9mPFXtv2EhfAyStGWmMH4aToA
hH8n9ds5RYY0OZBNcGrW5Gh8DAHtx4oAuAPOBvYIi8+56P3RLxxv0/jFlJPgaQix
5bhCh0Dh4W8SuLiEYQYq6OvM2ylwwb7OVYbxt7LGZM9f548n/7mPrZ4cVmHyX9Q8
h+Kvu2G9haoh7bb4gqGYeyBhMu1voVmzFr4W7Sdd4UjJ1fsuZIi1rZ3+X11vo9co
uY8zf9UqUKE7NwPGtoQoxiSj45q6r4z7TQWm0+omCLURmSDPTOslgGqTViza0y23
qxt7t8TJXcQ5K+gNVU8f/YCQ1gzJLEJLSVRGpG0h82qU7IPHk5qT1o1yipiAP5be
/UOJsNP47je8mScT2gAit+/wnKkeQmbfI4tdBXRrAoNDDm7mzGo5xXsujO8VAJU1
1le0Xu45xbYIVflYB1D3wJuZCBUHD9b9fOjbgr/IJeTeFKIccUF/KWST0ZNThq+C
KrxZw8Q0nNuw7mSPSrPV7CB45YNKv5LcpTPL0VrIfhkML6LwMhouXs5F3A2tFqN8
eBIQg9AbFHWVFial7YFmyTB8roMyjoXGp8dKzbL6L5DYPl+xwMt24rhAG7hHFgDR
N4G/u6ASwa9cKaIASiblWJlEzz06iHB7ypl3Uq1T6lML0/wDONA1CKxkoK8ocEL/
RFhz6J3VBg0no6jlw59lr4Bz4e54Qv05PJuV0SRfiHw95eAsw5sAO6bgJmiuQkD3
4zvjPz9s8SYhwrtdOVv8dwJ4O9sbvBtfBeN3m9Hl8Yu0g7RVkytrxrwbfXHCzuXQ
tO0xKMyXU7m0scgz9q6myn8zgbwiEasrpMTS/0Yrde1UWOevK9jDePESa/dTjAGU
iVvj9UatF1ytYWaMrTqRUxE3aYsOAezs9NW2Ca0K+iaVMtlD2sBqQzvj5vwYTo1z
2g9wpys5VXcg74qS461e5PVj9Qx2dTXKIi4LtQdUR218VnELRWr3s+vzFxGR5oCp
+f5OGVAHBZLc8q+rSGt5v78DyR7qy5/fWAiNja6uclh9rIIRjwlVFy7VLS4lWAOZ
lm4Sk1go9F4SX1Thw2KFb7+ugopwY4e4jp4tvx5XJTZFk+F+YglSNQn9cf/dHKiu
PVHy7MXC6cUlEZ0Ubq2FcCIDtLEVWpR5j3GzghSpDhNeL4cDvNHTXD4ls8DkP0mv
vOKf5kZK0fR/p5HfqSsX4yHNfsYOTs8/shUGmYlYfE2h+4mIClOD95eLUrs2ApRS
zbocSovr4WLz75So5ayMNc+YW5ICnMqWirDUrjwjSPwwOAFjsxmVvukgzPnpe4lo
Uaslmei2dp2Ib/vGXBClogVyTnLo8BJDBxgbPquMP5dShKv/Dv+KfbMhZ1V6SP+L
YW7qF+Wmyna4bZlrLRWQjEqfqM2kzo0/+q7VaT5gy9OVG7AxPwfef/kKsTYLKQl/
ZgsKe2WQLRLDb9wLLAYY1UhRu0q6JAFDxoAU//J95A52VGe7scyXqMZ6B6nvgRij
Xy0QTLunMIPdZ3L2p2pPHzJYGYcpJKpRxreqSQKhXqVPVczCs7wJTQ5dCe/PaSnG
Nrpmng5f0x0RfeCpcFpoiSGqUOpd9rYtVLdEXxODjCaJTBtXnDP/jrC35S5a+oam
DL6SaHTg2EUcbCxhjUouMrWX+S9MA+8f/mO8Hre4ryGcI0/iNmVXhRj5S4/R2vSz
yTvvBxZvZUKgoY4K7lYE61BxFj0GYdGO1cPLIcEx8fBPJg3TkGnWLPu2kGx3XFNX
HRqOHvMJpWoq3az51lQlkVbQuuNaLfmNVQkv4iSNO7rcuTepNRJaETwvofiE1SGX
843woVM8icaHavjrpCqqjf8HC6JqcA2urvVyzOchvDCBsymTTHbHjyDKUm2yxnLV
fFPzcQ66qgEO2PHORfY8Up4Uq8cBduQmzzNPTRo1iggVe31n7yETb4kGVU5Kex5P
rlbGoobxRC5JTTTXZqmLKXtzkvMFZvkf7dVMyFRsjzPk9kkZXTkBE3oxdzHQQJGw
bhWL/QQE4IOflIpcYYfu0zXLPBY6luraMpm4WppuHjiluvSmRRMCkOheL6WP7QwX
JaDFgiiS/YapvjaerHEMnrHaSfucZYuguKWdwtbbDUClClpFN747vaVnUkH4Tg8W
xQrgmV4PiSCPfY+9mAiy4v3AeM+/pStBwU1+gxnXkbmyXtAhjqyI4wNvv0tXGedK
8RDqXkk+5Eca/9FeOu8LM/98a+2iAhY9mmUQLjeDRRuAEGIejG4qG/+yvR7EvsnH
GcwgoQCRKJ9T7qI4DHlm4UiAP0ZVGXzXnFp2uHTz/Gyf7VJgzXNwsNAQSbe9tWtl
wkUdYkDdZa3DzQsKnsAzhODTJACOP7OXkoC3hdtsNXc2D4SNqKCt4eCstDFWOSEg
JdRPIPjWHNBWLoxYMnTrsUyl3rV/Y2Mg2KQ2F2CyJVfPhqaOpIuRCOVaVaKUhdJ2
VNYGTYpBDxkzhdsmtpjqvcepLi5vY66WJNCubY62i43wIOsQBp/5CBw6pCWQF/Mz
GHhP+sYY1aH2W1mAQAVtD8FrcyM19WCJ66beDAS+B6gf4p2KcQd0EWzFkkfNJWlZ
pp3mc5FyburJuqeln8coEGflBLH6gWDcrA74ZaGrkdiPMO50/sD+/D/UFk7yXYak
Gi3UFLOg3FR7B6qbt6oPWRkIQiQOqunMRH/nBggdx3/fcgg/RRoRswGGzP/x8EyS
AGCOWlgDmRIZvkuxBuonNreDinn54shw0SS/Zs83h4+SFvoSv/2isJzPrzj/JOse
TGlZKSOotcEhLHoy902Pvl616Si/xZQt4iRpU+mjePprMSB/al2XPg/9oRSg7XPE
xRBzp8IKJ6kiouhIp5ucsMYZqkGyiurxUp04tBfAmLd8v+E98HbjVQCECBsFRIWN
JvZeIyh6vYS0qLHgi+ZoIZEkIwlHlCBLZ+Iv+ssJY4njYjoiXGm5t67uwHueQWsD
VNfKcw+UrVRKPCGeS0LbQS6eqzAH13ORyDxFmgTIPWoBFOxnrzL5vuUfIWKDZH/0
4hg5vIwKUZHN3vSYTjludh49R37uAnYP6PH9+vpzMvKy9M7d1GrlnpcFwHoBJhzc
gfl6ZMxaY4lyiyJy9NrtglDnGg3Fj2qFoZc8K2W/iJ6WQxZCbJGMpu6eo8aj/XYf
wl4bR5di+ZHdNmHf9dNqFtsaWiPUj5v8STgof8sfjckrjQJ+cjKUlT9crvDhXuB8
ZegWVW//Q9YuGJfdFUH77VCYyMLcarAJ2GtjZw04HbNOo/59Shpf4TcpVFjb+9Gg
dqyvELVZLws3wK3z2rLYMpQA2GuFHJHNCb85W0UDz7MpaMjr/9dwDk7UzwvhKB/I
Rt6arvxmcHVGcF0LuSS/Agi103OpdG7qRqJekUvUor6RhOz8EWH+qbb6Sfl/MsXs
4cIpawJ99ZmcMMyVWWp5sbbdnbeAZXLImPh9tMvOz8hj2BhistRwSgmE28runmC+
9mFgnX8zqs/X/xwbDMANYJCEzlMNY39QA2ZRRnZxIIwtmC846VK9Cu7uPo7ob5WG
Za+xGq3ADL+CcHZA+o98iN64GHUetoA1X+6KrZiEdIA9rJd5wccPncTl3u93Snez
x8+Lma0psUpzF46Ks6JqCvtX3rr0OPboepiewfw1YC8dqI3C5tYuq7Gtx+eFAB2z
A3NegCRbbLjpGOPzhr6RJ9HPwnnyqkdkuX+CBj59Osxck7r8W3shIL4IDuvLAvQ1
oYS1FfU+M7Xu5ShlS/NmoLqL/owAey9DhGEWd1LcLKzhbEseV6Lsg7aQ69M46hNl
y416xJpavX5Dqrii+3T6kSwq9aNz1z9Qf9HcDQJ9b1WdXlwArM6GyLhVzxkXupHJ
pCWtsk4JGHoZqWo566n8mCDn8JDgINn792ETAHzlNeT4LDYhmaK3e9iduvj6Otl8
1Vr31+o5pMjzOGBmDyow5NBxmhBW/3H+Kt+dx6EkD1gq+N7Ok3OENh+bJlK8Iu4u
N5XXtI8OV3HvqCLMlMljqCqxvjNKqPUP4lnuNJIxa38IF76Xob1CCrZVeI646YEX
rTZy23KLEeByksxnhLNSoP8tO4gi82tb1pf04LtdI2SRRy6l8usG5LdBXg2CHmRy
htsfJMfwS/mPaZQMRnABB/D/ndIsnT3U7lX8rCoXiXAFNZZfkT1FdXk0AzPF0hQN
ossg/Z2bDcdChShatijjsf9aoiS7RZLnli9FQsgAwYkRpIlkXenn1sioU6smseTv
RHIKiVe23apevYfmXzaRKHwXgA8hQrL0gA0ikCdxmCnuy1XZPvdhP59xcUntJFn3
BEy2im1TdwKHB506YPSr9HYBZjHOzLf1gw6zm7GJUA69nsw/jvHFAOZI2MmM8U8T
ZjXuQlwe5E3rCO72rQRlgFbVlF8vLz/yfszr1Ugize6VzCFWoq5a136I1Vj7vnBM
xvKsPeZ39FUp76rVsp2EpfLmbjzf+ezqi5M9w4ERBGHR1ltlrZoVUmPA5tZs2zH2
4bty6rX4DhAqwmjAeHB1lhygRWfBq2gQNbZK3QXB08hLiM5d9PPYF9vppXqNA0Iu
QiM91MPJLvUOrcSxySM47d6J/iquBNZoXph6BDct1rCp8mYBm9i70fpDmyEoTRbs
ia7mxvUlQpWNTt780uyoPDPK0FuAs4/QCYWHsVNW/InnPJhuA6zLS7erdOjiPEfo
8hCWCLYvDznluWJRwVvNlG+AiXOun+ApK7h7D45thzg3FJOl+7UuNWxznPjZHaJ0
D0bzfauRvGnTCbq1zO/4pC5oyv6USCJ+TbaP2LHDlgsaKHcFPVmtJ+4evQ2qvcUs
EWX3pTJjSI9gnPSzj+Hkf/06bxvg7ka3SrvjtstR10Hs67lerQIHzQrrwNdxXYlT
/zZNUTMWblW1oYijeeMwQZyH7ld3sKMBxLDXr2Lvosk5MAXYUTsinaWxOp9wZwEe
ykGNI7wrcbONs440b1ub6wqB7al1O8qzebm17dLZmtoCPYwLkhurlyszrHm7X2sU
vjVLQrZ2vqU+gJzW8bmWeKKhWdioM1ZwEzZgU8KlZUnZDbWk42f3HJ76VMEOCGrl
fX1NyvmmNQFeUiMbsdf2d+SmiGkKRgLEKyFISZHCxvVVKAWBXbNmXKLuAvAv/wcW
zl04alzp5lcoNaVQHcQy2Hm3zQMfNnI9oih101teqjSeUjp7NGvGvmGUlvxgtHnG
P2IiLUhRYfKw7u51El5ug7QOKkN743XFgaxItZeJEKhYv6Z1NzSZscud8HrlyM9e
CQLMd1zvTGKvQR3FbUH4i+4FAT9Hl7fPIqPo+g/xSYUiydA8njh4JWWDUbMqmAnX
ua7345vj64tIa350w4dNedX5vN/uDN+K2jDLnGarOxNloG44lEczQAqrYvnQINMf
u7qk7JCdWm6Zg+DnSuPsw9yluIcKzOxPbLs2TYFVtgoeCOe/6T0pWMEr/eieu2Q9
PQfEqY3vNPHWPjtPUFp+G6g2nUAm23gtB1JECEPRrcgt5OKAfZkXvBg60QjrIsL7
3MW377s9GIFJxcQ7HnYYt5U1NiuzftONntzxUKpY4sUb29YdGY1wncLC298kpZLB
PRXaTYp66WHSy6UERRWA5UwOcXLxi131U+I/GrX8Hn9HzlX29HHiQkrsQvEw5HM0
RpclB15MiRubnL0qc3VaKcm5+da47/uj5WARcLvXzQyb3QtcCZLI6au2Qr7xqqku
MYXV+NHa5C9ILQiA+fbEryQLSVEvvW/SR5dmc3GZjTDEBnKpmh1/+GfLUPQUeEWZ
2hGUrGzl+TvZI9OpMG3NQ1FCP8O7TzcX1Nb6BMgEjVKI8aRx1wZyz8YtV9LHT5jQ
4V3VY+WLnr97FAgu/8mpHLiXQV4o41u5LTYPErRLkRd4DTd59PzoP394jBfBOFgZ
cLTWWP/duiN/ubZjYqIwvGO0HFG0XyQShbmUvoJ3FPn7YIXgnRmZRsJRnfh+0fKw
BR/uRKUVIv9hv65TrbbeZYrkxsLW3bghkV2Z7DjfCANJc+L6ubK+BILNDrRCN8fy
+S52biXOUVL4vYhSelH4Do0uKHGNr30peZv3EBeBspOKMR8VWyZB/s7AYjRYQYCv
VhvLnEUQ/LvNvkTl4Ob/L/3jHrGykIdwpPCKsy4SWblsZbDWpqU5VT75B64Ut3pk
puDsIq129bF6bdQMNShOkTbMxRPm6qAc6ITjUfaCTfW/ZT7P8ipWTyCnZfrgN2jo
mUcfFeK0DG8zFbo6w1eVY5qCl4VDaVkHqZIZQYTmsg5V1nTHLTvu3IXM1cIW+cPB
9wiKH0M6Wfu60GOlDvUjx/bBeleyvgw8rquc6T3pelE/7iqQd8JENCf16D5fKSA/
FRICYyEaPgYrl141f/0Tw6YiUGwgSSkeVgUSYmMVTy+PpGmsX5r8YFQo7qrM2gu7
cghCaxdI2VBJFbe8dvpslMpApE3oSgqhWF3uvFq/VnRqwp3/zSxU3WxZ6MMJNT6t
wkySkiziZr2ZU34xlu2lWhVf2nxSTKm2yrYYAeWMZLq6xCgk7E6JJZbSj+9qPkLx
GPZOeC83fcvRlWLSBoaafUfT+kV5PbajpnDN66PyVBPr/KGB/fEXJm5/cVKjK3k1
SYIkZ/P8wiXGOY5x+tLPonKmlnh33n4+D/wRFrcWhYPWeXTRPEeGp8sAtObWlRlm
EPZzdeNgDQFid//QQuM+WIGpGzR342DhEJGmEXGV0kYnoFwbXJlFME3AYksSPWAB
N3/G5upPYZ3o2t8zDi5L+7VWQ1f86Z6s5nvUPys9IQlOED3M7tiH+5MVSSE+B2rj
Lk6R7QOo+W4Nej+TF8IDOv49aeplcsutPccnji/Z0j+wfLTtrWTnihASfeSGm5iJ
rYkv+/UxgLvwTl1oSAqyUIbF9zZmalbcl/F3j78S7C/TVbcnDxnoMXN8YYSSyGY1
A5lYSfnas51EGSjji+Gvqxx2MNm2PnzF/UbYcug2jwuCU8adjbfVor51mpV8mq51
MEMCKdjmZePpY/tRuOPtJp3U1mOntMZQyI6z80Vp1+NgYkfWx01SFA78e3cMWN3W
U7ICVZZMxA8cTCcwknsJeq4fDQxnyHvpjxAqXPwt31rljjV2oP794UD/jvqjBabC
JULfUQKKn0hwIfjdMozUpW9m0yUZNHA1y6K/x+Sr+sgDwmEOgcjDYxBrZQz5PfIa
pzjnn7uDYF4GZQ63mSOM5a1YzepKx402ElZQuiWKUmY/ry+Ts2m3DTFakz0cEASr
jX5CU2SdpyGJ8/MnsmPQrqB8DnXMeHeXqnHwXc71d23SqapFL/y1VirGQbCUIc6W
K5PGJym7LuxxHOg0ELjpaWH31YQboBoBWapzu/zlVslxpUSWAYit8f1nEJd7Ridt
jyEARnjsxRUWATFMqyp3/EZ80xXJ8urydoRTDaqwW6XSAfIBeqI8P/dYEUDtzGbH
mBdJtznzjjkiA4CfJbPeB33lwGkRJjyLWlna55CbsJpToNbPZLwMQ/G8Z9yGHaNb
xsXTu4ls/fT4A1wpO0RmA1tbAtUzvOXoPrWxb9H96HO+Xkngy96MBfSPRkwY1Cq1
Q1hFo9QL5+GPu9SCGzhe79icEWKmUsiDRztCmYDWDFNi9EEF17u+vYA8DzXsnnGi
82dhI7aaOAXiGQfJ53ANL1LYqehiM2y0zwDb5BG/hhaH2caVf9hirla1iy0q8OH/
JrWk+hWdDt7k0pcwhPLySUsLnf7E15btCN74Npm2cYgvZwElUoWUBLJfgh+2isCY
7+LnUwjxXvsRMr2CtzO3DUWjFi9kyoMslUkLNOU00bDarg+F5oZ6vTKWX4GiNaiO
RUncuu/FtU51rDHJJIQSXVFUTMllHfXtX9NlA9ciuw9aJXQMQUV81f17YarS3mew
lMYsjZ+8YHwmNfoFoZlFZJMIh78LNkoJlcFxTsFtr1aXeiBdQLfrW2xLZEv3jNTh
6RrxHyyAEAzqM2ydnEQZg7/+FHzpKhfhXcO5kGeoZTyUbswejKkFHAaIOAF7eFnu
D2jDbBPlEsmPSNtL/XIaRK90FvemBySaSZGucsL3yOq6Ib/sj+fR8ep1x2BF/CXn
w5p48mZFq/oBPa0hamzBJmWkc5+KGwy4jwJ94R4ZBocbv2ZzZ06tbOAJGWQWQo9V
b9adk95t5YY7qOzlg4PmBREW9+pt5DGmWgHSwW1HQeSN0zgSnMMmY9oAy1q+olSy
Ze6yFG3Pf89v+c7pTkFzFUedWGjcCLjsqJeAxgKSzwrhW+XsllY5Z5XK6xKJj7O9
DubOiCacqUnUeiWkWYZx4BSWs8lPBAJOoNXVkaZRm6dkfkaIX1hUQEGPnYTSsmtv
zoJMhtButWHmBvm7XvmdcSDmI5rZuay7KGIAkMT2GZTZ1UvgYZZPajJ5v6Pmb+IV
Dn5xb2eZ2zHghemLyacgiezxvo4Qbp2yN+pgCUqqOTk8mEwZ5psJXsasi1jxcCVg
1qk+PS88bKUu4q/Au8ZNJJt+9nuLKeKgPnVMw64t+GH5yw1yPJCUb0Z8nXqcgxrX
hCghebocSD7SEPAqAF9MvRKq0zSGyy2lyzVhFJm8ctkscUoA8FsfGwp4pIHTCdqx
MgAaI4wxr/cxcsJM/bBCmiYqxhHEhTrTnrrkQrVqa5QnKVAPM5oF42zha8dK3dS5
9nOJDzBPL+FeRuDLQFAqC+liCLX6VRaOYut3Ht+VYX1ZJKRqfl/r1BWGD5QPtQOd
gQBD4iBAsicSjQHVPiRS82EUXVgNwgG197Yofr5H6NtE78YpesGDEKaAJXMicx8I
vOe3Qejh0TM+5hDqfZoVuNvKKMk9+Z9tAvJYjbS54FDmQo95GqC/eB2jtH2iGFOD
udKX4I0fp3KOWWbIPG+0xrqfkbdI3iMikzxy79n24mNP+Jtstp6EMz9L16tvGcQB
Sy/LfjFwOTwxbFL8WM3h/YjxgvzACT9kKmJZnfXSkWV5uBB46dv/vnWzXNWC+uDH
Pmm7+OdkTwGHjesmg22PXQEDgHxHFkM7WiDJF55zNrEq8dIgBz3FeD2bC43nE9nK
WCevtayIPFrvWY26YJUnLvIVqsnw6q+qGmBTGbfF6clNiza7ShH8ToE0lKspPtv4
9gsBLgZ0DP2Xrgg/tUGCSSCHLXhKlOwa6V7+dOebKeDy7aoE/tQ8B28NAytDQy6F
RAEJ25AbMGimr9RkelocA35xMvkEbrqrArQi/p3zdSJ1dmPkXvVXwnuA/2UHn0WZ
P++XlhqWbN+S4LQ2BDqz/BZlxmxI545bnqyYfw+ydJBlaAOQX4nnk5M+9KWraUfA
5vjTqTloAf/UKsLwD+uVSSP4zUuYibkgEPBhmG8kxttcvpbCKPPFJn8j6erLupgC
bzg+DRFW72LOdJbnfGk0ybLsLJv3tvUt9ctnTe6Tx8A/RltzFJORgKUb8lQStjor
6WHVlIvmfXuEdeEEKZkKJVDgILlCJgzPCaXE2lVgpr5T5u1Ev3bJNu6n715NE0AY
e9X7G9BLClkqSmJLdPA+9YYeUtyKkdYQi/lhN6OydQAwjMqynNPNkOzyLXMSYCdN
LnN7V1pdu0aP7ofzLjMx2QS6uSlOFSeDgwFLF9Fx9pjgxtyGX+AWEHjfVhdaMc9W
cHwtP/YmGGqdjBEMg0bIr1n+TwtXAmGkUh9WgU7ud/ykuM5rkCh3XOoD39mJKB0v
R8APj8yjPuTKcWWSPJmTIT0h7j0Ij9vdLGYNBXvCgkGY401bEsi88P27NvvzJb/n
QWCNUQ4h3Fs2jnRAB4EOKdTGNyekIgQ7bffBcd3/JSqd5KfB+Gv8SHBSc4z7FCmy
5esL1qwDH/kG1Ui0G28go0WAXV8r6AT5GnU6oeGBmuMvON+DN5REWvnfGv+S0ue6
F5bARIKw1FvT6uyjzJtpRZtMG0qc/7TdwhiOwDz5ZycRkvzMz8Patb407q4KXDrm
4ApmKHoI8AhcZY98fn6DwQrzJSAxZz3uWcTHHLHaQn+xvcrK+eB2REaWkL7g2Wki
jdaAHOmP7EYW3fkxn0u5YO5+U1rsz7rFZ9tS/6Lrjz6XNvIVmOD+udWUyOR2YeLZ
1FW6KGnl/NlKby2KUEKAeztTMtWgnTauy6aaF0zsAF/HWFuIyKBs9Mf0DecBBxSf
hbKCs02Hn8N9y+JUVFsKk/GghAIlv5UH2cq/DkmV/+TNYNt9uUJTTVUQlBDOZ1b/
csk/L/w7G2wsRa6XUeHoYbCZkvCv+94aV6CGo6k8+vPXgvh0YMnCfPrWE5dd+/cs
TUKLIcJBNDdpt8BH39Qf2alMgFUX20mP0xnpbL8dFZmsEBded6iJBWVvm/4XWvRK
MfpY//i2QqoFtVeKhwjw88EVWIoZquGCTHS7xfgV06cxGHP86i7nl1mehj9DatQS
SzPXS3zYJYUm4MnFmXRzMiuLnjv373sFlrj4/thFYtGDAMfRQ+XIdmzBb1aMYYa5
1wZ2fDuKZ+qwj4BsQ7PBJVI4fs7NcMRIuxoXb+guoZXaohAXNkNK32Z4PjXmSMi3
3IrNBMS6HAfru3cPy1pwdTUqDuyAewRFRhtSzaqfVoKxDdSvWO7ztCG5/mxUT6Zo
2DzEE4EF2wlvlxuxfw/iYu+blPMv0GhV4P0llswbZReIH++K0If4XbrfcboWN9Tp
SfXrasvMgfA1O+tJv+eXjeEXHVpWx1h8cOn60EJ48hKyOVItlE1VNy/GcOt2YLqh
vPYY6YsP8xKFSZAPqMeAcHTX+G3tZTXKcVdpL9NpnrSi3vfZgMZJNVELoP8+DDvM
+m2SKNRwwk//rSEEfs6VLwRba81PdOz8A8JCjWHA7N3E+B7OHwlX1/6o1wO2j9YO
E6ZZzrZM/KSY1nhc6YKyurVF3pUdht+lRrGLIzYYM22zv6jisYqLm9/0535Wap/h
8b2Y0jb5tFvV7ak0c95IDyMi5M6NevfvXiJrT23kmtpe0yH6TRJj4lLLXlZTJ5h2
WETTFJkhlcURTwdYZf6VlKkoPiBtnW0xZ1P5w3ZixlZgxco5iNvYAeS0LYZxCkIH
3+6fyhHWlIZo+6CH3gDJ9t0d4JFU3qISxLPqepzSpVzLwR2b8zxHqUSFNaHOQ5SH
5j5QJddPYraJuh+fjSxkE4vsjL3X22Txhjtz+JOesqTrYAEmrVS5qpkLxxpZAi/n
dayjBkb7adY/IQpEP1ADk4pdDHPOitareHjJIWkiKLRT8MaTNQfvh6hXaw5clOPZ
8DeGocBbTQDDiJJyxgI3/mrThpO+f22mcUzMgLSrm8CBCoDDBBvt7aynCp1/eiU+
QrUBOVqOuR8ACgar81uLW68CEzfHzOrQFYsF728SKJoaakMWGgKi/NV0gkx9UJyy
qs+EMh9eLP8DZfn5pOuBI/0qQh2hdRU2JVDDLHVmS1e2I6s2vCiNE1gYkz7kkD3e
K0RbBDTknYa8lM9eG8N0NSvI6feh4b6t4fg2B0yMZYPTtVIYaG4vO9mFT5BTURr9
P1Nt58oJDPoOuZnczLWZT1lnot5BxT84Wm+wtft5gcx9XNnNH2x/NpV5bVw8+4UL
4meUG6vvP/+Tpgcp3naVjxmnEqqKVCqnWk1csMXQHdwG3yKur/e3HC0ZqOHMKXPw
t2JA0dpcOYIs97rQAUk8lW2qzE8deI6V3JHg9nBkF9A4j56coKODwE9IGTU47EUR
MgOdX3IjT2pi9JHh2A+boXs1nGfs3q7g6EUEy45Ps9WqMYFSYSlTxOSv0wUIlAmn
FoUFeGcjctKjlSj9NXmpWX16voVfBxRlcQeaVsnDUeawelZq0jHeEpO96ZQd0Ypm
7CY70U1DMXQNwoAnCYfb44UTdHTk40DEdXWoEEb/h10vc6RFC4eFIdE8Y5UupDtr
GIZtDku/5vpvu30UXbYQMdm/EkRTfmG4l4eomR8mOyDOKAfkPz3QUztMrNWWDK3a
Y1XgSGKVhuUKuMDUbKRdx3mbWsXkKO2KZaSLkk23FNET7g666FiX7sKPXhDhVzlc
i2BhGesxw9wjjzfhS9ulvCNRWIKGsB1gvZvrwrKSMHnFbZPuArFfaB3koMaoOMRf
/Cfg9t9G2Zzifboi1uI6JdSgdyJzFtOVOGBG99yUVQw7NWcSDohSylc7F/20zHwO
8HUsbtS5RXttLhrg+REb+hoSIj3VSPk/QQbhHx0PJXFkrwcV9tbOLv1gPiRsKaNp
51c4A1VrBzf76t9HA+hmq0kghJ+Exb4aAbV6YzqrwUsfTc1dFwMLisax1/fXZlkV
/n9zgBGTqSnIKf19H/U4AM31a4ArC1qFbZ6da6kuCRrC3/Y4KYtBIgiGLWvl1Lps
NJCoUiHSVXBL+uwEzDEzSdvbcLLhLgW2bjfm07YP1OW9ychiQbKrRukqCYoOQFm9
9pfoSirF7qTHsuqUjrjqxcxpeo5EL++KQED6fUSmKA2PxnlcS2Wl/hr4B3dxdzBe
k+c858HPdNSyte1hks9tE9LnB5O+/gO4UKYhUPJ2c+MC27TSBHyImVbaj0KeLOw8
e0T9FxKVqq3mREylDQ3qU0ssgPn1GjAblNLC7Qld55Pj6Kv8S/te9LCLjy+DJF46
nhprKZElriD9SacG3orDV0xamNuJnNa3WAoiHtG6DjwjD7xRUGkH2dTQhJZEzE9u
1MpxvkFycwSvdHWasQbzEaHDNp9swH0/aHi0Lrfu/hmDIcTteTzkDtX57smSHBNm
Ul1vAU8KjWFD7ZOLRcoS03ppOw6s0J+qMKhL+ghSdMmicj8mCbmOMjl5C2CRptnA
YUqGjWJcvFq38XzOFz4mYbqvEHCGZ+UTKzJMjLAT0GWRt8H3rHDOySPG6lRilGuw
ch/bqeNJjDKa5tmzbjsWKjiLi2WlAvXvp2FMu2JZ+3UoFrIjYpFxt8uqYBsBQ83+
Vd4Dsq3cVcOtH4KZzqwxnwDQezJP8c75Ae6v0ZjJ+X7BbxmSXORqZ6cCg3zzS3XO
yTLTtQffx+6t1U408HLYNv0QejgFOPXKHu55NUG7TiuMyU8jwfmP0cjGthvPqfrY
hMui2Yb/YQ5/hzgSY8PmfDZBvHyauSkSo11g5Ku+wWGlUr9n1kHdx7fhN1XKHE5W
x2bdNqZIN0PELjk+qELdx5uI0vh1YX9IPslg8Fl8RZkrrgU6WBHMgaReSk9N37sV
j60CF9WlNLjxxLQ61ex1UnVW+UECY51HhkAmoL3gMsvOJxxGRXZn4zeolk/MnOyQ
IccpS7d4Zadvi+CCJUsOwkeH6c6wVf6MmXtiD3Xm6itTukWsKz8AT8pU7atEHIxZ
3hstbidDw+avKiphKLYSDA0TbQ2+l12Q75qze9xKBMJ7mV0vwHOreOiC0ndduyZC
lrYZKlM7zdspu6Wx+Ht8+hZBOnoJF0Pty7PyigXnDLIBy7BWsaOvgCQEnTQmSw5J
d94B1rRQhyRzzAZcvpih1y4Ag6En7SAf7GB623UvUaOC5F8LC52XqqDbAzTbV4Wn
kDAPvA9CPJOTq2tCOnZR2l/fgtGVSAKcSRtLYJPadVdOJzmrcmINONKfqPIiWGHJ
UG1w/VNEM8rvb8lOU1+jlpZF/VuGTh3xXdNnNlQV4Oxeq1tdVwCoNgJdP9LG9hLa
dNTkvAfLLdhfWaImNZOjEi3ImdCSZwAUD1HJovQt2Fo16ytpmspF1POpU/M0CzbA
ykNMFTT7KOT6yDfVRKEw7TWMqAjXSRQygpctUMmaIK74az2ytUzYDke4c7bWNlLU
b2DMGcJ+BUVJqZA0NHuA84eWe3068Nlc8zfv84oC7eWMgAhcyM2Cwj+3R9IudPyj
bbRM/EadupPnmZQmoFzogj0S179aKeK1XUUgmtg2kBCu3pU4/j9gyeIOwpPBOeYX
w6LbtoZ+Od8l6LWHCc53+NxoAd288zG1yixTDI4FguXzIHmeaMXHOFtdEKLdw7rU
AWvb7f7hU4ZMgW0hNBc8YrzH4U7AisZ/iinUMYUojQTgBKHddl2ZRUpAOt/DEZ7O
R8IIg6ai4zYZw0BUxF2N/5P63LRxQS/HsQXRjS1HeoojpNXb35BaxdgMKCvqHyw3
3PrbRb2Q7PbPiS5umUxigNqUwLPZ9A3rQjOKIw9iiW7Azsa0PhdZ8gdVXLFz01jN
2N35c5jhJk4BuT4iDpZhZM/kBEATKRQxzq6PZYtqxofGjwBEOXQ9zeEeR9+ah7T5
ggRePWmm/ZfX336LrbrrLxNPeh4xxzzDHiRO8bVP2ukrFSAL16OhIOean2hv95u8
Hq7OcHN9zEvIKlA62y59nB8xzBVllSv7MkzMTKhDxbBFgW0l2wVbp3VwtzV/cmCn
IW6NALRhbWP1+j5zpdeuqqAAtT7vlokmqh/s9QyidpEZe3fFJiNq2Yp2T5+WMp4o
4BDEdYZqx9sE6VA5qvaVmLmlKie464XcIFoOHvJVRzVHko0pxKakqOcz0FX5J5Vl
D2KF8W+7IQGFGRnYdd6W4UYuzyFvTAFCDQSgr6KtVccAGXhtXDpU9F6KCLCvXkdB
1DznFV4IVNxeyPabr0FWfy9aOzyQW/0Igobs5Lhk7vmXlZcnxTm0eW9ihnqLRFJs
lkqGBVPWa7NrjzbWdZMFDOzZYHtwLwhtoHqy4Gqs161hMgCFZvmvmaflbzNAWCmO
LkIkn/dsucce4vQjnYD3euKvX4BbzUjyLuEWAFrRRkuJ9gdHYVI87puVGb9W+JEk
9poqQJvT+iFGjFak5vkqSvarg7h4sbZrnD/BLsjjVItinpQqiall8Zs88FFX3XiM
MCXmZcj770XD92Lw3cYlYUPTvPREvlU57UE5sNQCml4MVfETrDF7ZUXQxfhtas4J
siZSV11vKyqF8s1mUpHZZBbf1d2RwejKi1ThNy+dmyQXBcH0fSeVWMgBDh0yHoDt
MJ3lPT1kPiSxSXi5MqsiPRr0fHFEo0aqMUkFmWJQRQeWYjA7QAAWi/FR3hq7CHPC
Tri5xBWNAqafaq5JW2c7TuHSPk92TZi04Ls+bmqwvGuNQ18uyszXrfRYbzkpTP8Q
0UR+S99gGqdKySBeIvMg2qjnGp8nYl3XLdLuj8pCem+kFsFJY7uoDmNz+lyH+t0F
Ntg9ke2ow055JaPZOt+8ijhXUv0vNKdipXhdPnwJfU4tsy6HSN8OOh3DyT4Fy6cj
Qxq6Z2qW65ry/bQxLavh64mfftumLme0MNtbgcMjvnPRJwBcMqo5kgRsngx8Sr+P
00SCsRFcWkLpvALgItclpbpTg6XCqfw3JuzW2Q33UNoRxqg1ZyHF+ZIhcJV1XWub
+BMkaEAGzL05gp85Phukfft1KEAIp4mZHNrWldJ7UM0PkmVLtGWm8w9gCg5Jxp6T
oE4xts03sGXQpGTaZGP4sQ/WGy8JWJukQ/42900gecLUP5S3fegUu6W7haLUAHev
BXZyD/Zk8CsQJV6UBt4AaVlZi+PIYxsREKcGDTQVnqFRZ/oYqmmtNINsoutYtbJS
e221FtO8EOdyh1tQb8rOKZWVirkvjh6zAunyOZkfWrro+bOy/NSkLuk+eq4CcMB5
3ngDPg28dw7ct0SSw3nTVks3BzkzqkxZVohQLQ1rtjTfc81IT4tNvEO7cJu7Kk8y
asZ6720mpTUQjYWyasQMz6YC/q4uni9FyHYSg750o8NLHF5tujyP8+9MF9Z2grVo
0LorvGGeixz0UJPJai6EFjAeyDSYJW4UffnPuTYOfpzejvPY3+o25kn9gDEh7VTU
5tUfixZuQiNghzSuMtiA1O8mAb9VrbfIMQtgpyd/tp+y3ECnGFcVuJekjee2TXlJ
/BzeBqX2+WpFJB+PPFHb8Yx2pmGjSnHwlf9tnSf9UZ39OMlULn59PKGbRBGpv4fz
CNoAOr6L8DoDrkl+T1bNZYTTIFVtejPysCba3hk+SLkcIdfNcztyMZ4tZbqwNVyu
REFIDKbIjT2lPXjypBT2beQZZuKjigk+KkwSYRHmYxCwg/iK8K5bCEG7T3CHgDIe
Be08P9D+NfoKbMdSzPPD6dKgTLmd1oCWH+kY8kROL+0GWrhthwUOFblaqwdtelX3
Mcq5HrnR/O84uQ+r1j3uAvIi6lRITrsY+tYdSnOdkvXh2PVQqEqi1rpk+J74bxV5
YilZVhm65UY0PW8xADX6zPLZjAvIY/lX1BIstwxakWkRbzLnpJk4nnFYCzcS05H1
GhT2Y5CV7GOR1tjHGO8R//c7OkAbRFMDGEUi7kEBhVUTgsuMPwYWSuzsgLedxR0q
RGpIjAmXGmcKsp5UXEjgLi4KUIyuJjgDaRPXDBxr5kYCvgzH2A/ybb5CGecyA80g
50z0XnjwGmISCRQlvqSV8fDKHCLikwGbHxEhr0LEzxFI6oJdN8DilOC8HJFGnKBq
rTuI1AiT0FPIGoXXflJg4oXE1VXTtvHr+htQmUDaFQIlqRVwLZ4b3wT0PJa9IEaG
obd/11kBo0oPDpDITbRVv7QYNsK0n5vQHf9jFotqfyamcrXapCY5k0aFQeQb68Yc
bfeB919Uymmo944eL4Fs4oP8bpUKizcce6bz79uC0kXMO9jYL2Rm7MPXIRybFSio
frjQZelBSY1dgWSW3d+nJFQKYxoYMWa7PNyTlAGJEW16kPV+ntVvE0PpKdfX4SZb
T7pH2C0ryCwvS2SfVQEKX+rsCn/rvbA/hGIXbzOucw2McTbrUyN16iMJpKc6wtlV
F9s6puZQnpSy7F9watGY14qdcyY5dXksUau2bpQXCJcHcVzbHb786roOLyvN2Bim
4x384+ZQkLn0xPgocWjQSukbTVgXwyxe2M/I+6E6XjiWXsJoiCpf2w5d6SfZkK+n
5pO0l+X1D8zh3oNfU7mL2LiS2IetlPaf1Mrd8Oc+7q6udaa7j6FXHfQEUIIqLDuc
Xle+knLgDAVZyAM8IxODNuJ0FSjrFeHthicpblNnQTmG2TjexozzfuE8MtyKhq8c
POTGaYcD0rHLoiRrTOz0D67ZLHkNa4MWDyrMMqHhZUAXH+u8KWl31OvK9QeSXGsM
VzkID1ZpUg4fUh5IHbHqzuUx+c+wQQpNWuIrUP4FPNyD3W0CI56Lry836G7WPdkl
Mj9tO+3vtwR0EBUHDCEZX+c7lzSCnKpfuHFV0WBCPW80m6klPiQdL16dgkUHAc4h
haRzJHliHcx+hbycBehJRFfOxmMsPgU5hxtPm4hbTx9FwHRkJqbQSVJ80dnmi7ev
eaKg96MJNy9rwPGtVpCTAlTDSmsf0Z6OkOf6I+pGdonxWjPKZ9iL9CPh8birPu3X
QkHm/Yf7KQYcanbJ88l/PlE/7SYvvm5/YrXcVoCu+SK7sOnP3JZfcFDG/FB+1aJa
0ZR3Nr8AV1ltP53ykgoYOyxh3QHf3GIlHKXo1zRZTWcNQxIYN0gXs2TZ7ImRktNS
jTdcqcamMIfIHgLuzPSl+LRSz+QWiiOeh7bBG0CSAvgu+8mwb1iT3S2V+/fkqGEV
Iwa/Z1zlFngBVmLlF5fNEx2vVZ/zYYLbQBnaKSeBC6Du0l6//AnfHMX2W2B9OW8S
mSgC5GHjHHvFHFF5NjQFDTwPWEezepMU/Ew7QOvt4iu/gznUcxdqVLgmvXF75sD9
3XW+MYUiPlceFh7x5TvBJLQgrbF9PqIFbRDdwklamma9jw49ppcHvjUOju72FuPw
Fn17TyyZDkVgK18SaHquGC/6yOBm6+LZNR8KWKMYUEcqtRwfhDqQiXr/aV1/GuVi
pL0AUFSg2M7m/xH2Pfcm1kqQIkMsre2HOWkVwHUsWSus7Hw9DpixowAGylNjrDk4
No4g4J3MllymifXSO0GIu7xXgyXgJcgAjco1fPl6uM4DcMOekoKgBV5ljWmYxc05
Rm3HkhSmIa7zRT8Y1X7gmExoUJBzqFouQGplmWOCWoe60jtsbuUQMmFkt7srRgwl
tOVvVrqV0PeQ/OYeUhfqOUlJ1rDM8ViF9qF0sXoBFf8IPUdKmOTJf+5MLPi8jSIs
2jTFMDNfLJ/8hf9jAWH5NVAoOHv3oTs6+GQ9uW5/jMzJKIH5nDYIvVQcmg/jO2lK
BB7M6EZbKIHZBWOegiCZNNCdYggvfzWyMawTe+kMJ2MS/lRah5Rju11Eyu/lU2Hy
6DvtolGhDBDL63EenHJKAd6lDnafEU2PSX1RvYow513e2c2jZLTM1Vewz9QrB6mo
NCK3JvJU1BiYcsYWmEQmbeGdI8Pdp3ZJKRSdtMdgdcoHdlHa70UuxW6lKHpSPYzF
lSQc0C4W69aqmqhchUPxQf0Fy0QOvvYOp3nKM+W9zcUec4W9aJ0iWRBMoKhgDe1Q
matBcafdifq3iOaAJPQI+JZBfTjwdxxiJ+PCVo+l9p1SuHd4JP7LJk47Y7Ba/Uzo
jl7xc9BN14diofoghi379VW5niCZzZqT1mVtJMhllRbwLQ8fviBPxiaSSrNfCpmj
3KDlEZCoGbzbqEaEaGUP+tZdEi/BQbTtj6WHug0ru18ldRhR1HpXatqjVkJi/7jQ
on4XTQ5etZoXcEP2CkhId6+3GCQvuiVkwJvkBcR3L77QFQOZl/axzP7UWVwyie3w
hF1xskggl78a9Wsiqefnzs2+pTnkUVHARke6Q1F9X9l5KfFyuMjzDa7DYCQUWJ0l
lQWH7poCSgusjhRcTL1Rp56HxeihVIIySGMI327WtTvIT0M+vZgoihP3h8DK+vzk
GoGROCkkHdULiUHCgc5Q2dAYmwZBC2OZe6IuI9QvZVf2Rtw1iH/FqFWvLCWq17g2
uiMyBv5jpTyruT+LcQSCA0ZkLHMjBgFkrgshqBhCD2kqlnbGB00IcQx7akA6bygv
cuu+mXM9bYfpa0hFHeJGsLqdSLPYQPJqmtBucFSIgXK4n8pDmJCfeUJZxZl+6Aj3
1wnSPj7TbiSOz2+4MroMKMDu//1CVkRtC6zSSfT46la/S52NP07p6j8b9reiwp63
7QQeZ7p+UxsdG+uHoCmlzc2m3dvvJGdtLUcOgO6IW6QlXXkVvYTwoQsCPCb3q3du
Sfyudavaltar87QhRbrbxRO9BYE6pXo/cuBThAi3TwVHJSRNJBxh3o7QiNReG8Ff
qtKyyzRJnt9dMdMqLsDI3LwiwN1wgqQzHzkwWvAsAS6GkaCY/dc7AiDFKd1YRgPv
BYMGhgUZefBGIIG0wu5KYKHJin+hb6Pj8KngKSS0kouKVnd0hZNclDjvu1e47C4U
Hbj6GDB9IqF2o8tTwjJTc7Ye6WIwPBM9TlSbuWTjKxy53pVxFPTZuBiBmXPG79lh
91X7oQk22ZOn3b3nDQK3uNDjGbTXeCAREe0xsIzCblMJL4B/rfCE2rq3+EX493wC
zKYxZw2ABXtC6aDVyocxd7mkb63CtbUekmbmtjFTB8jhAmrCsS2X+FEiTGJoSLlb
zhUCKUnweyYTzomnyMCtNSukQaGgsZVY+ABpm07LFIJWs7YmdS5FbmBkdIShSCfS
R90TVcWFQZd2ub04yyEGNxi0eJKjwUYvcxLOBOVBwgSuGoUBgkQs/5jdeNKcoVEI
8awAVuD/Kl3bvc63CZVRAwfNaBjpcg60yBf0ol/WJmPG1xI7ZVISCkYvCP/w/ktH
cqG425as6ZweMgVBnhNYgwqZDHIuM1AMPOo21NIMe6exGq0CRZMJhObnulPb48Kr
jt9BV0hCkwgESgtL7nigAMNUb04MFYNft0zFaa4dtB1EPceTg7rmonVCeWWleSkA
wNJ3Y6jQU7NN5BgMuD8mnk7AMAlKHQ60erljDN4iwR2bAe3Y8P9Bt3hI/2/JdXM6
S+A5qn04S0CVQ6c6TZ20KZIhSrKNhsX+syqeEZb9jWi7BDs9MgIXs+Zv4WUg2EEE
G63L1QLwWrZOrmcvR+XK56Xg+d9CK0ynLg4lN6HXGIw4pjCAxxRk09n5SdV5Hh75
5b4E61Ff2LNI7ZjRUR4BzH+tWhr/1avR8gRRO479ez5GxwwU5X5MpXSwrF0WK6LP
NWByYDm9qZ5YdQGXqOFVSKVJpgRUe9X5Sx8LA0suUxhSAloFFgfK5+nkucQoMKm7
/IRDg3RhDIr8gzNqAwty0xSBmUcM5sAqWQx5YgG8go9pb4Cpjb3SrTqbkqr9UYDe
pIrdf0ZEsSqub8EcszCUy4+x9EdMxpz3nTFlsyKkTTIf+mzp6b4IXDoTo97hZ+89
bEpuBE3JjIUouL1HJM1jWJ2fZRF0jR/G2GaYeDtwfR1jXWqMkT68AuUObQtmgzs8
9UPQ7NXee0dUIp9xc6zJxF6XUxcWR85yqWkwmmsabxjmLzA4RacbYWiwYmem+Scf
adc0wOMXk9iSPvCZ0+J5R0XM0ip2yIJtK9Gv45uzKpqfLlzumKB67zVhO6RnmmB9
TQfIJLh0n3krG7rNK7XUfzK2NR1DQwc1hEqy93T4WN6Y1fcl7w3VmkGTxP4sg4WU
E+lWCijNEJrJvbsWScY0I3rEGguJoTcYjF60VjHqeaaihFwKkl55tCcfCXOqHNbM
mcbXZEGoxvu2E24o2xdPLEjjvJ0Bjm/xWND3/3BWQ55aNcwkS+ihIX9IFLICOVmi
CDTAb9K1UZFPsHugsLQZ7QwJw8xQfe6qYlMHjOhSN80BHDsf03fp0c+hMDL4Z0NA
CDUELfY5xx9p9IN5d8d/Lrtrvdq/mFwDU7OnvI4XcGeJuEhCrwZh68wwmlXGviTM
83qmxFEufG/DK3nckLoQLn2FzXIiohOsuK2TiGb5ALZCbusDv1xnCtiP8ttbp2cd
59yZu2ganmNz6knHFrUCQglNJg8aGoUjAzS+bugZ9+hvQuVAaFCbfvx9kdOl/Qv4
81J4LU/WS4vSviZlpumg/CMtvL3ebdH8obXYSVaHmIuszOBUktrdxsHSG1Y5R2S7
rG+n2dBJTIdRKaPUvMCMUP/xE0FSBCAoAeBL8IpdSXvPlqUkYA8iHxXd6u3yxzQ5
8P0GsqnmdIxCBVNvxZqIYuZw4HiXnzHlgAFQz7TB5V5TwwfdgOwP41h9FK30AFpv
OjGbTi61FKkLHS+OXezJy8+QuJvTe+hD2+WdWGrex+RAyd9FXUDgduoYG4R0jBPy
VuVJEky9BNznF2Q12BmcAfYV0reeXkDBTjy+sMpK3f+hjrOdnJFf+eLQ9QvOuMSE
itZ5sCxDDhpUrEw8CqtjedJIAXkIaX2z3YN5g/a049CaD5Yb0I7aUwAC3w+S4ddJ
3tCqV9PnP6BiiX40R9iUFExX0cIL5C5MNzuFjBq215kXMpIT5CbMYQb4AAvPDbQE
tAxVEseqpFHO6T4rh0e80V4kMDc8xZvm2VVQ3J+nDek=
`protect END_PROTECTED
