`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6FpC6UjMMYJo8um/VMEGnvyiVGGslg9+qhSGQVkUY3VBd2etzMYEg8smdpLZn6kW
eJR+ge/eN6kxkBMGRbXEGKhSDncs6zjBRTGcJkvV6FMURlvnxvGQi26gMKxt7Q5P
Iae6huIrnPEgFx/zGY/wZxmO4zX8KKpxQldawA+7GGyp9mCm0KSiTSZ9e/kP/YvK
vMduixE3j5Ye3YDo6PLbzhj9+ou4wU0P7Bngt9angUQrMxxKCeXWy0pONBLo7XKQ
hQ8JaP83riMOne4mks5+X3/unLtRY1CQ5NPnQthDjKmAHmrgdEhXSHWMDzwsrmou
G9EjLIqI7qYZJbOS0QBM5YGVw83RcKNBGBDFV3NcGLziRXSRV7NsqciwA+auxhfq
A9DCFUOc0PHN4vSWgsPmX+MaSX5Fy8TrrZeqfVCqnH5u4sbJL0EpYdDPu9IbIvrK
iYLWs1vNbEABPrEn1eJpLuzDjlTaldsBLca6wrkIOM1zqepKGHaFge3RmLWAmG5F
QJ9D/AxKm7F3bCR4nFBypRfrh4aZ3V33FT37XZ8Ynxy19ydrl6YSuZ2boydrTyC+
33LZo35O2TRDTsXhuEjNf39n4Vh4B2oNbT8raQp828qSxZ9fxiu5U7xnCgKRTRAK
aJxAnoiGhjpdlVvkYNsEhT2ZFA6be0/2fU+k/6CgYBFl/1q+/eWYYJDbZ4yykAwE
TrPRFZzWkMgWpCfMgGbEAsz9zc62+UvW9m+FIOVmzqr+kbH5zaqS2lES2kCxKmg1
GyqtYQIGWycz2CXqAA2qKUDOs2zZu9bW7dWp+lj/SLohb0Ex4JziNEmzsu/b3mdA
QakLrfZ/p4PZW2ooRtF1d9L4pyHgentVMnVGIF7vzrQhY4/LTDRSjdkZlwpxOGjj
Qr8MjrOPMjC550m2tZLihJmGuxvVn7LUXgwPFxlPuoDRfRhUDhLvg7XUj7xtGlwy
oBwdbl70Ep1uZK7W6hmtmvW6He/iSGgylNErtpr9iaWkdCpXIkQR2XP2UX/BHcQX
jnmrm1M7bB8SUCWPiHZSROY0Ta9+4l3rCwsvcDEhiP1EYQavbJb6HJcBM1aI/i95
fcMMICcJSqCMYZqoHfYJVOI4hADn03YnxjZiBg9i6ZmiONPt8+pfI6c9Kk0jQ5z1
DvDH9dpbzIVQxm4jdzYyHM7U35SuI4YK3Cm4eV/GiPFVTRvfd3AkxkOk7bKq4apn
SNl+AcSJN3eonAmZ7UKc6SMrGoAaldK3YIuJt9do/sBvRNZbRlED7arZu8nQJMj+
ymu20DccpxjGlqST/4zzbZ4DuT/YhDjITa56B4e4OXl/7sICZc4YLILdfwnVpDd+
xFL4WsgEpnnUbzj6mtiVz2NG4Y7UDGh7G4enHwmLaUerFQTqDsAyJNXVsnsVvfxI
rzCex2ixRB1hZKu5O/vPrhL/qS4BUgv7miVWa0fYX0WgzjJ0qvXeGTw2tU0j1sOa
tGtwul866RdzdgFk4BpLnPVZpxoa4cMl+xPdNdDKpqJl/1bqMUy/SOYeqeJAhSuO
2/A7NsLHoEsZtMyVzyFGpgtnfA3BWyu+YG7W0yeM/YnobloQuwsQzQls1prb4yyC
Hkbfamhy2Ch4NyAK2RfIcVf3qIn+hrgXwhhh4o50U9D+0I8qTt0swwX80zLIfAJM
73NLwdS1W/IpmMQPpatW86cOmLQEtjFkDXGJLhDsbngyWRJQ8SlBxKjpCY3apb/E
glDXQlm9QLgHqHb0FHPChJhEI/cNESXXW24fA/IEOShCuYfjGvCvDZ71Bk4Lrox+
Tr13P+TA4Dv5xFh8fFSfOqtGm5fBKB68R94iytJu7JLxFYapq8Yeo7rhPTDT/eGQ
gKlbG0p9NOOKj5Mh3wT93mD0Sh31f0iIq0Uz/wr/x+c02eiTPaRECzVJbZdmRk9Y
N4UXa/sXPTEmXUnkfl6dgENpsqWfTUj+2a+y8Oa1dHpbcwWp0pQa8Hxx/SEp9QW7
7znYCSkO0OStdVrVtVWC0hkPpTll01Q/KqF/EJv7D/AE05VZkLvO2a6NfoBTr5jc
WR7UDwDVe/HqVsPhapm8mZoJmAwbPM0HJZxw5JSYi0MwcBcq6eQoxsIs+M8LKdtl
lo2LKHRATGSE+CKaIX82C3EXY0dLEPt4EAiye/y1u+KK5uMAu/q0wQVlxdOboOpF
YT5Kj1O+KcxqD2vZ2WUbu9rhGOCLhBVeuUsmi2hKayZL4lG8yXM8nnaPVZ17SduI
g+JMauZK5CrmiumlgTZX+V9HYMjt+Uxynws9CT+5YULSCtxAb3Dv/J1Buu5rd3v0
fMOJnBJ21eCARuiI/qlo/k/Ddos5+RpzcVSQyYaeyYww7QiUrT2cgZJP1Sz3rrDE
aoQwuR3biXoPTFOH8Ss5ri7ANSLr8MSN5cPMMNkZ51QviJfouELXQNzlF/wWyTxM
glVb+OPHo8NpD6rQOsQsqIPYAWwcWjWOoqJ7lsMA2dpafmK2LmoLTDXwyhG4Fb5/
aJi6phCx+ObAXQoYd9W75d0I+ik47+ibcydzb/l97JG+WC3v5t3qKo3uFKR1N/Oo
6ZaYPWzTUph+/GHOoFGVxFDvJu+TtjDdoEqDEex7N7U4uLx8pzEuhvS4wnvn0wiP
9854edHypd2E5LMC8tJOIHuNjvx3zpf3i3lYIlfRDoqC+pIicLjBd1sNnKd10tuU
PMNHAT/uzmXyqtVLihK7jcHMTFJjDQ8GxPPi/JpZa1HPJawnXQB/5n9oVk2oWh+l
wkvqzt2oe2Hcfgv2A/XgsEZH5OsxqqNbbQ6YWLLQABEkNJWuEZ7ecTS14KB9X8xX
OZ/wrkqIEDMowoM7RZBhJLRHjGCdhuddnZqjwPHcaa4=
`protect END_PROTECTED
