`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yx0yvbsZCH+CDIu+smEHn7l9gWXUpuGJiE6Wb9YbBOp0JFDyxeaOtJIWTB75HN1S
8+xYGf+C9SG8H1jnMrzNJhbvdYYrJ+ys12dd553qKvNW3KYuXwFjM8dHqooMdPTg
mqNj6cIv/Ko+x/70h4bTfil0XZxFA/G9uwRlrVpykKu18Z+tA/iPMHEQBuyQ2DpS
VE2HiDhxxf+LQKd2CB/jHEt/NvkEeYIIw83z1hM9ZSvF6j3BxEIw7eChtRpJNB1S
kijoOYSlfCq9nWlBwu7xepA6WaQwAVJs3YVm99LAa3z7w+E3J0TpsOdhZm6J1j3L
3IMBgGN31k7L08XoE3xcoa+ap1E/QtcMACXGf+GhEGa09o41nRorKIPLAIqZijYg
4dd1oG9VZW/ATWVlZg8wUh8viZlBhdcJZv4F71dbYCZ5ay4eJ0PvhpvM1izzA4X+
FkKQgbtJblNvMNabqmxhv4oGX4GUU5vR3oZlBvVzNe7y1zYZiRtYFF7I+sygYqDZ
u4I1Vib59bcqpwtS23RF9lGsX5BY32f7k5UIG0NDaP9wEOl3mFUD37qg498xzRWm
KCa5MJ5Lp/PLFhDFpWvpljJfOSGIj743JXqSQtNurYoU7a2nH0NiE5W/lqab5UWd
jtN1BV2JrxOZj7HLSA6lYHG3+jdGyniBnxYZNZaRd5N8Hwufi+rtBuTMNYN3RyKb
XuMt0ht+1tO6AJ2/R6Inw3cTydDqXEPe6uVAlVtReuTGQTrUY7j3/SfyGuEMZ4WF
YmePI/RRPRbJAl0+l2NtPQyplOZ+EQEckAiwi9C4UJjr6pphRcTlz2Ee5DqcVZjT
1Z+jW9C/DEKG235NbZSfJxEZmqWFSnsMxcl6dulvmqexjt768U5ngAR8ZmjK8ZDf
6ppV/bY8XlBgNl65qAq0n99zRip3uQvZs1YHkL1DsSFXctSwMECcWigLByEy5++6
F4tmAphjFB1uUmNOAWzj1FAZkOQRj1ibBFps5pdTcstzQX274H9LRzgSKlZx3nrc
yyHAleK3LCzLcYyvDYLsHPIFR6Fy+p4CjeU6zhzZGnuLBpYdfOF9pDnLTEL85bpq
MZzFLto7eSa1BxZ7rADzWSpwJAhQTTVhP/aWehRAGzFTz5l3a/Yd3g+htb3BhXMP
J+YW8fCNXJN1YYj1giniBg6W2O+1gH9/j/edtto3Geafl87noZgkn+SlooDx03p3
RUgR4Rl8CjEQJkZFij0DxaSPGt81k4LDdZ3V3gfNUgKLbLmG3SZjE+bdVCcl+Onm
CrU2pSK9Q8S+iZ9U7JwfSqLJlutGw/Ei76cFp/EKc+z6BxEkrTvV3IxoFNyEFBNY
4z14nwdgo87qBXR7U0Y6wNNMz8NixYC07WCpTk2bQb0zWILB7cQ7sBg5Sa5K/uSf
0ss31I5JkTXtceVDlIBsPzrZzANKoihP9DKM3BNLTklRBb+BADvHMU4wVqoFGsO+
sEzGa5WJ9+VoFDebO0YzIQ61lMpSzUuMNLNTWUA5royLB77ZZvJe01xcXVV4Ow0I
yuwaNOeforLN3l2Ph3l6PPAgI7Dcysp85RRyYaraZyKsT9shHub7o1IcwLOkEKjd
gOGBVJs/UWH2bcbk5zjAIJG2wdSQZzckgrefYwK7WI8/hjsjVnHgHiMluOOZy2Yo
wRqhu6+OWHjcaTbZfSoR5W8Y4RZuuoWar+pEUhi4NJOlQ1Cah9RQImemNyyxXpDO
xJ2HOuqCY0KzYVDrHsXWdiZ7n4py2mqn/RbJVg/PzlgXnnhDKMQzf4Yt69sxKEpu
XXvKy3O5c47PJbYKG2IrlDi1DGD3ytCEQMTJ1tUo1NJ4sSlAIfWFz9n+dF7sMGsX
LcyX/ZbpA+hy6SHycfRoQhVdhtav8Jefrvpgz1MTumoGD6RhygSZCP/JvizPovU5
7ZzEYN6qQwRBOS5meE4Ur4elushflaE2TAvUhxqypFnM1yTBv/6QeHTHvd+2vj8Z
M4lSyxGw2iguRQxjJ4muMs30GOCFZ7CiKKl0/ecWRIInEsjx4uKOLdlaI6AbWycn
JNlzuozy3oCrxUk7OP5hnfGPWXhj294OadY2DT+8Jr4+fnic+ITogs9nmUu7c1XE
18JlXP2c9mOvApnbkP1KQiOBnWCuhOJvT7ARFztpM8wr8d6ftm8lwlJB7k/H2aEM
aqI4im6WyNtrISf6qFO2ElCWOOHxDXe7w+wNEDlI83INOluRSVXnAGfCLCysBt/E
k1q0ycbcWlN3S+DU1HdTjeQySSAso6HlxiQ2rkghIWK6IdD86lcBkJ9LLR/iZWuy
u99gSlyODAygod9an5OmejqtCq6njOUlxR4RiiUL7W8G66K0cr8E7TM1lP/LuhNO
enZXB8CKfBJzTZTexrxY0GvpNd2qf0YyYUxbNIYEzE2XFQAoJ1Dwt0nuSkbS5XB7
3a4tlW1MxM0ouhTGtA257N2I5QzBbyQf6v40brQXhO4sRmPhEsAfI+ddAUs90zb+
WBIZA0d6deEXV3w3N+AaaOTP4I+YnQhAXUvWMQRL3keWoSk2pXuUnf/XW7bnG0hd
w69QyUlLITjA8UVKUvpQV5vwjNQh6jL9+uzSCI/QrZCtnZe51LZWgLaAtyWwb2sO
qCPJ4oPbpxVcbmTJzYoLS5Ks+V1rx4IKBu+xUTNZDZkEakzFd1nMYHSsPcufGfod
3RJJ6Szi8gf102MwSj/Q1NCfP4Bc4icrpIkH3GsLI2Nt8jkT7CTWJBOy8KofSROP
uWXI5qCHMIJHbiG7Z2dz15HICslys4RpEUz+v449COyA74WE57jPZq3Hl0M9DpRh
pd+FtVeiQq/8QALzDiGuvTUwNQoBL9CbUEENmoV23sIzHKtoDhmD0ciYPAnOFdZy
/J17GiNZk1fP9C+PhqIyfYasAhwx45hCjEGdKhJscWnbC5kPkYHhiUdETfozXUQr
wyUXcF8DUEJmLkGVmFDyTKI4Q99OpOzhCqXqHivFUwDdoPf2nbEve6VWnUC1FvHh
yfMsxnyEg/VoePuObuKWgZ6IpV5eWvRDh5IiKPz9K87p62WM43lm5wv7P2Ta0VF1
YD8WVfWhIGhK9G8hRqw58ubErOS7+4JCFXYyn5VBVJ0+7EHpIPx1qZ6RR+7Tm5nZ
CniUoz3O4ncgJ8q7oUQhNZCINHuoMmIgGw2gWE/9ScezjroDxMJcCFdUGRSXnyTR
K3qmkM5hs3G3yM6xRLWT/2kXqqzOwURI+5qA/gpJuB2O5F4TnejRyYn/y4nAd4UP
rVRjtomdYEdIflRy+8qQNxMdZLycjyS45pQfGQqLVS0eu6cjMIjnUIpvIU6fkXNI
FBN5VdoAMgvkahCD6ftBNGS7iZ7XUWGvSC/OLyhB87J3xaxnSY1AIgF7YPjb07IV
VJI7u4XMwcqGXrOxpxCmxZtUktcZIvHzGzwFU5Rf2nXz9ehqmWGno741Go8UnG/l
fzHeQPDiRo+ar/qh0Wms7hmFcd4ENedynS/Ctqw/cWDurBYcnKBZd5oIHJywxooB
nS6TJrXygDqW194+LIQIwuRyzScY2DwT4679skV13hvFiogHrhEWchR7/yaEsViG
XHPsj2uHXuzFs31nkrtQFd5ZtCAqy6lcY/I8svECAMWxrbc3JtnSufx2uVSyVjmj
4yuIDyX/riz5fNo75JU0w4oZVZ6Tq8pdzDjpIHb9ziI4Nt/sqk+X9idzGWCbOhOd
0ZSdshzPB6AXlFrFVg137DEoy9kdMTEY/Ow4i3bF0ifHBQVVJPJM+izZx3KxEpDE
f+ltb2lfS7PcEb33f+aO25DN/O3ge8f/rzUS4gxfniWq2G0hv5p3H0ZcsfvZmCTo
FO67lDxnhuYy2QMZvSu60+4e/Gvswe5wNITpQkNIfXgZT/IChdNTbJACHx4gz0p9
Cp87nIwkDnm5PJcCPgR41tHYw5oAHth9T0dcF/4ZltkHITCROGbpOu7oA8VbKTcp
XDPiKUeP4xy3tprSLC9sD9wMWSbVAVSu2Q9d3P76mreRv0q/9UMg7b6hB+7SvELc
WYTUYO3C0cNhNEyOlfb1szzjwiqC5iAnJxUZMovZWUBUNcnsxBrxP+6DJ+VEYxZQ
q8osTsiaACDZwgLQEnGLovkgaxptnOINfWeTnUqVPTxE9Y3KohjDnCi/ODhLfYoq
XAnkDXMPFotAGF6FMp1ZfkH7VhYMS5Akh6mmLWhaVX0v/5t+t2a7vv99cl3iC14C
7QdgW7Co5jf9/9dO4VmonoYUsI/SDZvbz1ltHVA4x+053hzm1vz+PmZbFIYVCwI2
pf+V5frC0nCrERlVgrsqwxvm5CaPFZTZzW6y/q9UhBzr9rmdKgK3qZ1NSvNDdxZK
y0hXzG4DPr2Kv6ahi8fTux1pqAegWFAzli1Q3rZ+amrkG11k06JnNfsVM3AmXaGj
K7P5pMl7bd/VLil9kc6P+fGu/Mku1sW6NUzw57uGYOt7w6Ql5gm4RdaG8KkPJOcH
Y5jT40jgrI5PqMj3tqX2KbHjcZ3IvdGDS7vuFCquAcYmEgZjTlR3sYZ164ahCEAR
JfD5Ehxga/pDKcTgv+FxsVU0KE/844iubGqL2tdlBb9d6QHIuWg+0AijpY/vFMkW
7mGklvzBJIv+VWKI3bpstxL+FMXvW6otyFsgz4BoszKeUZYAPMNwKn9GYi/V6wH6
KVcQ1HMBVQakw5xQB1luCfLRnV2frmNLPssMrX9KYc/ogs4ibW98gMeTeUxKX0Ha
LkySJ7OmI2gRFyHRK1W9YxLi1QdUOe3Mr7RHGdbdD/nU+VX/iC6On0B4gXK+MvlI
zKid774KK0BLteednOoGzwFwZ03jyJDVUXOvmmi4SE/xcvh3L/ALR3cQbla11nhP
Sc8UyQe63SiKFwIhCXcTMUHnXcxG6lt+tDYknmRG9aG/GDlYDDoCSeM+wnBiC07n
fo0B7+UzAtWyafif82j9+tLfDYZJy1I/Qwo964ZZkzc=
`protect END_PROTECTED
