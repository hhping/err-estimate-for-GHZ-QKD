`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w5tD92POs3QSQkdu9kkVboTPRjBM5U7xlC2+As4DS+AddinMRsOtp8dqBWaPyE2p
M4XuV7qoB4hOVM4l1tlx0otji8hiGbuvcUjsDyp5YjWD94WXf1SKol7AAeLuApKE
tkw3/TfoSw2Re45FwO8hMxI9B2pfpNCIYcfTouvtKfQXRdOBHQT7EIli8T8wv9NW
O09hhdao8CrdeoQOQkYXfpC7ShZQrhG6KXazxKumbWdREfPENiXSTqFsxqd9kNVD
I5T3VhW4DVXA6hcn2AZwxcpNYBve2YbkhfZ+Mj+/SiYsY0W+J1aKFkHoig6lyD7M
oUP5oXWtPZcOdLu7s7MUl6DQnLL/TxXtb16kTCVV+f2QEenAk3HZ2ilck6Ip/6IV
38IwMWLxbwEEiHjtgUBcmjOyIoNGA8/pf3Kg6mkVRqG51MMKL5V6TcihOYzaqCEx
mh5ud/ZPdPCPl55osgv9zu7/DADoOlpPPFkz7DuyI2T8LKzoVEZ6W/qPEjGQXkga
hsYTka/wW22CA4K29vrU3I4VIAdgT1dJogyyRe8P1LMmuI79hX2dK4WArJyzG0Ad
AoGvEK9hgmKkVNVsjpb4cempQz7k19yZLk9vWtamlKcI0INWs3KktD6BHPQcCYE7
qQFenx8B1A7xU7oAm5jRtvfSoXBgYH5QBlAdpPnm5JaO9KDphfeHUar/zRcElvpP
9zMbx+xnjDvKiKpFKDrh2NkfRUTxgFQZ8trZf5dlRr+zhs5f6u+D+IzwgbKgaWuZ
7PItTOilHsCfB7eIWnOwgK/TNUqYuvkABUkZzkXBveDVjV81WrVkxaAUTW6pYlPk
17/yOC+T9HROFXBaiZcRHcCetAFiUKhIr45hqmhXoe0tL/jnKI2GKYmzW3mBEG1y
Msmmpic3BMprj5dsz3Cu8Q3+rBzf/eM7PK+AeDh0kXLpE33SfrTg+vtikBSujOD9
Yds1xUGvRpADuZTrTyyafWIisx6uVAKLVadTchdhf6d3XWWZrKP83UuH07F0QTWj
nssHMvrtaTMkiDfWW3d4OqRSCHHt5eyn0w9f1fqw15rMmGP/mh1LrTtUa8UIo8ul
tlpl89htbe5mzq60PRPik9DvcEz6MWfKNBViVRL3w1WTh/oGi3k/FXr2FX4nAi7h
v/WpHYZVbLkAHeJYRKruMYaKfecGLe1WGGTxT55+QuctyPfgn2xS289L7VrbXJ6K
TyFyViFBPbQkDrmRPFXMUi7ja7Nm/UL7/06+kfMRSY4qou13p1+FGRrLmMaxn7JW
mTIPy4fpzzJ6P2hp3B4Al30bXHndDi8T7o5bHQRqIioCGc0icRiNsSffU2j8XFwh
rl7nF6SZ74XS42VzM14TtCrQGV8iyKNcii46GuEs8nzY1AMpFQKMzxGC7cEhZnW2
PzOLY3Gwxn9yjLpBLYiEeo+TjemcXY46pny5gk6RtCI=
`protect END_PROTECTED
