`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDBjZ+pV2ezWk0dsrkg71/2DsF6FCw1tpT9DoIqb5SOEAieDxcbMs53KYfWUo20X
JZsb5o76xQMa+IlWF+E8n3r0XVtdIPDSWjRnxzHh+w7aWz1OIAn/Jt4I5anVuZ0O
ClbqNAEUCeEycS4nbbZIzQuHpdLjCSMSA2LCtkESyJ6hUe067KqxjvONV/uI0c9K
UjDRZStR6GgxrL9nBgINt8fbkWtTOTgLdLy/cHXVvIxd4jYanMVTrxfjG5YcTFFv
mi098Nm5YQboIoI67HGU+GhDke22Sa2DjXDEE6ZO/s9KgNigPqWS/TZAu6lvE+i0
NwMbakUASZibOjsvhTC0v6uyKKsOYqqwIlO1Ozv94/M=
`protect END_PROTECTED
