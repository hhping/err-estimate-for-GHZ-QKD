`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3FYxAc4LJUV6cYs3AbXIM4tfwuXwU5K55W4mXkkPqZtojiWahCqzzTWDrk8FC0p
fTCIerx6STvdVT5Z+972ZLXie6vJ6S95kc/HPYUO6fi1t01qyjfZoMsVX5aUBfcT
3NppQJUizGfHA6JUZLy7IYQpVfJvtzyTh00KaXZxyMN3dOAhRnPVcGI8mXwLj2wj
WBDtLF6dHs6vYroi/fnv0z/v5RFW4usl2LXOkjQjDl5/5TTQ7Vr4D1gjLVCiRdGF
8AraUqX4GfHpf8/zfQ7Bw7eZqC+sNm3KAi+OIKzQAndVntv7Rw+RynMAwjm2GiSz
JjWp6MbHwscwvVUm+it9ElgHgj5Um+ctlPDJZdPr3oLmXNBSkwxBGB6QpivUnGmX
x/kAGgicgWsuDi7ncDI7KL0sgMtDTCPhxUDX//pQlHz88aApk7Pn0W/dP6DG7cnu
K3i2Y2ioiTEWa7kXbMvqENJiJ+vukAJ5oFtvmMpCDtNqfYpc17cgxchmS6eb+uiS
Oia9tCM89A99+E54dZ5Yn57RzCRSbMqYmrZkBLtcPVmixWU+unLxSNk/2EZCH0Mz
0NGm8ieaD2aVVTdAqYG1QBgS0RiYkFheLr7laTbvaMMr8jbXjhPoFqCjc3wDrezS
/KHPL0X8DNPmoKZuGGGDqANh1tj+8Iv1uIptPCU0YUBbsQDc+HHEz2+FrHZHLEg8
7Rmizvg+BTQHlqko6bttFSPQgK8/AnpWkKwdMbHpl3GTTpj961pMxwLQo9PHeyqq
zd6qLyG0ZhrhuS9HHEJx30+ijzpCS5NWvxrSSDcfKOQ9Trdw4iufVdpQJmJlt2HX
EGNKz+LJZyEZECJQMbHcD8K3nYmjPXov9obVRIxCfr3FYWeOoK3PEX7/OyYshxck
7CsjCjaHSYsFJYoE1y6L6d05KtHposw+m2cbdpiLL4p2ECJDs8msIA3AXhC5hQy2
oRLCOOoEm3wL8kJwKlTrLBnBKropybzApfqp6YoR/P6OHmHZu2FsDECOzF5dM6PM
+4LoyWgqlw1Ainn08jy3Jn0AdwUFch+IbcK4NbWdOhyldeJfc4loqDApoUIUVxo8
3J4z6lIGYDqHNiXr2oH7Whu8qMG7cyYnZZbbLbcOaw5cpqV6n18GkwyraYdEL4Ca
Ia+jqP87yNOE3g2Z8hCLJe+AcWjk3syqJ/0vdCU4wxHRE70cFUlOuU1G0yMqSg4W
zJfhSyo5yoBjR0KEV03/Tl2Tq3CxMZbh+0wbpw6hSqhpWBB72twY6i4SezRXKZE3
1uNZREoimTOWXgJejVvjkaHp35ky5TiIjf+6sYEuO0yDk/A5X+e8cLzSs7EkAB72
w7wc1661uRbPveVynhoFzRSWSHc1y5bOaOfeL4k96ov4lGDJBDbkO7gakEPsU8hj
VmhRAT35hcRm+J1OxcjdI2zB5BLw72Lhq5IJjDjVzfLipwUjM6AZW7NFgg0sZBxl
gH+Pp+DT1akKVcs8yzGI8rjx48xb/1Jm8VDzjMKsCj9CP0KgoZVR8mGztDbDzDLv
vyP1zBl68lSKHeG36snffYiN1vru9N/wuDA1apgyJ69yQ2/ww72400Gm5zZgCiMy
p8bF6Odzs2seX/1Z62TQEooglyNwQ7UGGzCNM8m3r4Cr9chXeolfKiUHGlty5dNq
IwRgPiclVMJz9eP79xYFwzO1Bb+nsq9MXgzUTiUOgEI3E/BG3q3zyLhugSxejetm
TLGfTajgtjhmVwog7VM+7foUtuOv/Obqcq5f54hcojOg+f7LmiunvQWgIedG2ZaC
flTWVIT2MhQiMvv2IeUupW4n/zrJmRouHnFL03npOwFCpngEFdiqwB+BN0iC2SYJ
wi2dbpHwe26SRUXBmAODY3LpV9lWPVi897LWEvCa99D8odbMED76Mdxd/xq/yjhR
Xq+/qGMdvSbMT1h/TzsTtpYT4mzgmn9FDHPcdEIdkhIlkbBuFlmQeadm925icNcE
a+4u6O3HQ0HnAmyIc5XSBwC7yKe4hVgX0KNU+D/csoRgBJwtCWAo7Qt0o6BZZWMw
/KSEnZDR3nSat6xiOCTsFYka4jEKXHs9iGcKB1JO4dZ1kgmtRcSurYs9tseuKgFY
1JLxIAbZEzpJKyyJ0jEX/4lKuVBENVttcPKG8Bft+bdThWqLzB8IAedO7xCgINYX
bsZYizPOkC55JAv5o74u3anQ+Y2fYySwe4r/kw3AZ61RqiM61ZB+lbtkhVEKSnVF
FwThh74FEwuOSIrZrAAtQZ8qudSGJqOO0XE81AGfvnR0oWLbEsziES3dj3DtmCAs
HbYwN/8/z3aQhadZY3R6klOa+nyXh72xC1nmOc/3exmurWjXrhbFvbORXTX2OHo3
kFG/N9C6u15ury43B80Gi6ahancRdQ3nTTsai2EyLL5W4SEcExLRviKa42zH/MIj
aZCuz3TBqkNopqbWE5F96UoQVv204Jt7mhTMqXI8BeHP9dM8Bl9B696oWkpIo5C/
/u9/rt30aqkcKZcoGh8vNc4bH1l51l1dPWLNZUTnCrp+Y9hiM7hFNsLZNuAiINGn
SMAXtrNXX7K6XltQNUMU0EoHPyeV3NTMjXg1SGNHYiTfFX+5VV1CPEdeYmuqPFIU
fctKdSSxfIlgwmdfh4sGXFfMm2QstBAmRikADTmm8Gl/EUHOq/ELvkwkva++CytX
EyecA1EMeIoMf1DnOthIGv85pGlCCibRL8a17bRZ6pvi+nK1a0ZyuZgnZM2qgk2n
WJf/VT9m7rOMTkdDYRBxhTpbcqLQLRlugrslYWa6BZcnahIFGoT0e/6eUuR3PhH7
AG79vD7fYkXxJ0MDr1gKPrTsYATBmCl12xAPOXp9AVFiE/8jQkGfdlIMn5ivEvgv
/GpBwUyriB0CKGu5SnX3nj4kMJZlybvxP7dCWSD5507kajDIC1yOvCmBOXDkb2El
3TIs/bmkfnf7stTM8oNeR1UPzQqJFy9jxa+IacvlCcNaM+iePFffQjvykHmB1myh
FLxwkzg75E9FlHO1TDjHty4NBfYO8pQCgnXFGN02It08Jd1CDtyepYvdFdFLVr3g
rI9F+uzFYjYUeC5iggH1hmlwvyEURmtI+r3xrkLE8woLYqWc1YjrgJrcqibXH4tV
2/L1gEw6RAp+HnSb1puv3qz9wVR49+PccGSgqVkMQnq8UgLsbWAZ9Nvg5H2iO8gE
/Psa+Y6Qu7mbtF9AdcO9ZsEJnLAOPkU/ghssdQlL9LijXq/DlX/M5+ktZUlATIiQ
5GqbtfZT5UNtyYJYTvBlUEKnn7E84PAhZ9XrWd4tsA+Yt/fEKuErCfKAP0CQyoqr
UaK0t3QYCZQezXnPYpE04UGukyokgRPA7lKMZLGM73Md6ko9rJaDZjHvBkeKDb0I
uYvz9/F7v8cJG3oZu4vjVg4+NCFK4JUH+AUiyRX9rs3Em90RwVfzIjlbAmaqZLch
pO7QWpiyp1u/KScUngLxuhXSblZ3HC3RryDEfv2YKx6gmkVbe8HoXH5CnCcIspTs
f1kq1Bl55GuJrj0a53KJ7yWbJJEDCPVKT275HWkYbFXp56x9ZYqyNoUMYtMnDGBM
AgQf3zf3MZaPSFg6+8bQ7jyFCqH0QJX45IxGPPPnahQ5qMF68pnDMEo/mFSGMLou
NbFiuuMJepY1yY1aR9RFVdVJQw9pnh9BosdsiMH/kFlgb8VDNcPKXNpDUmyQk4e1
7S34BMgLz/I4Ef1NkjJQQ/8fw/TiOuXB27Ytc2tcKVW9R9rGXsGo/9Rw5am6JTTk
n7wDYQ8Wv/L5STCA74LvitklPSMU8oo6GQNt04MsVCoSE060O/xQ65rJhOc3ihH8
i9956MrARFA+s1H1fqtDuw/lMwAR8WeuVin6h/jFkV2LHgVnes0QqHpfRXsj0Jp+
A7P6U+pyItCHPwvEfs0PKY356yM6lQhakX/ovqQ/+91KCSEE90I46uVaLsDEcSAt
5quYg4soJR3+OemNB2v1QuAYJGP8/q1p7kgiaC3uFJZbPZb6k66o/JYfb8fIIvXr
fJoyxMx29LvKGuMpdOaaQc6zPgWbrkddYtltNQwNJIqmigIKLiyOUSTSXxCQcCcI
WurS5idSolBzeYRfWOUbviL6DKg8JriTTuji1/bWiVXyTSjSdzPvvkL18gn48I8a
2cQbCQvv+CCMT0BOtsdPteU5dWhs1reUiH2O5fg5TlVkMzUzUj3vNE0vP7ajRwLl
bVm/lxsyGFhZx9l3nmb3zytI7Qk9fsCsy79PZvyRKYV/qz2aedju14+TJNp/8p4F
z48te/FVsldCueBAGtRjVVHYTPxl3zgGtanRoHg2mrWJHSByUxCpITlNoJF1tNv7
zgQNEp5yTSDmrzecs0L5RjuOz4lY+ogTgHokdE3cw3JrDeDKNzsF4zeqMlKc7nev
1CZQq/MU2AZgdjrsImbrjB/Le9rwpuL90fwCY8shCvwXUKlA3c8bKVGHHOPRl1N4
+61CfjKf0yVq7qoDp6mNuuJwFdDuHYoGNLKM1FN1Ve36rcd1xiwO95oS0XXERX67
faR+sxMvBwdQz+FZkW0arQIs0G9i0vvKxym5GNos/RPvaPhg3gF1VOMePKTV8zzr
`protect END_PROTECTED
