`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uvzs7vmF4uQabuNQvt+mKL4MgJFHRcQuV9aSXJgdXOyZQbFZuA96Ml9WS4nFnoWt
JrzMt03zKFshEkvd6475qgNVDso4lQvl2zeBZgtMjWfIdoYRLKLSUxHq9h7cRssA
mkBxS0DV/itnQDqLbJQ639UJhzUve1KZyveeUvCBVDKV8IGd0WzQ4jTdhHAp4XP9
warktKQC6i0P/TDw3hNNF70ESbPG0SHkJm5hYPKoAKjVMCsEp1nwuIIF4AtEKUCj
yQy+mREDyJGq6X1CXy5DNbPb1YMvi/6azmFuX+jsK+uxcn0FL4kqwBtzmJ9NAMDi
4rpb4lGnj4nfkefgJMdSm3Nd4NIv2DFVfY3yPxPxr/umCQZfGZ6CJy+jnqO9Nwbr
n4MljFCD64KCCKCKk/yOKQwxb6oPWKuu3j/z75a20einov9NtCcbGpJ5n4jwHv4O
WnrJQuZhjhB5zyC8W8qxh9hEfnnARZIx5zp8E/PN/UsstvEmAp2nE1+6B1a2dvXa
ZSx3ZbG4AOFZHTRT4HZlcFBcfZDlKVIflTKOrCOV8wUt2feB++Hxl7xakP7YEw0P
9Sk34vJgUXSsk4CGyuMMEgQWa4v76//bTJ+zHCKR/g4IGQFfEztLogqLp58fWd4o
efB+JGn5UB7ikYSUoPpDIUtxetlv7Jn1G6mTjiF9MjWgyt89873MWmMyEVMNSEKX
2d4oyW6RwR07JrjxDQIAGTzoDvfSW1Wx0clHHXO+mQDtCQ6pPep6eQaLHXNalkbQ
CZnKcsQUVY3o+6Olo1Q+8hVdSec4gMlnOKtEa5reunGFBDh0KaNYoz0ikX7KAHrc
`protect END_PROTECTED
