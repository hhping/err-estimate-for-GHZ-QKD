`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kIL9VtuPAXsSmqxQEOZObtwnSGnLyzNUTvqNajEUESVsMvI49FZOd6PsJhAKTo/5
ZhgKg64d0jy9UHlb5wSw09mXl7dLwscUdREyK/Rcar5YuVe3S6d7GB27dccysd4l
J62QEcTC4lZDKkLMCQ2FoU4tBWcgUZraXdw7NG/hnlb2rTvkCG3SQHchSaDNXicD
u3CKzFgE/K7tFpzdegHU/rS6Qg95jA70CpOQsSpErdQSUrDVtRgtltKOR5cgxNS7
oN72nT1fsgjZUV3T1zBfNJRslW7CbWHEdPA4v7otcnENWewrJgyCB7ZqucZXR9ce
abQeROtmjjQyaUwd9c6aBbRJDFApeNjcN3E6I9bIGrW5po5zOurm8AeU56yNb9XO
/TnmEytu9882Z3MfYjZSZlFT26Vri+73JO16q25v+CFRFRfSKW8osbtM0NoVpDRG
X9guOYfQn/vEatac0W+5WEu50Zb7ULJDmQxpYSJGNWQm8//jB933etk0L4A/9S1D
f8288lu2xG8l9av6BS8J/u/Idw60bGjMibRvr2k9L26qxWngDz+Ig4uJLj9aiklL
6qX533LKAkhn/rWv3Icpjoggy74YtIBr3qxgQJZf60ARGsrPZdtbZwjoUmHHRuqY
cyed/D4jm9sbntlaMwlkEZ4R6yo/68/vqGZ4RezJkn438ZSOz9SrQb6uSYil8Ypm
VeE6pSynITlXqZynUUylwN0dH2RNcnzmFcHTaOeoVjsPr9FOdx5Rw1z/bX6v4ijO
8z69Z9xm5JLnQP8kyq8ByppQOADc+79Mi0TPqciDY5K7ehgIf4rgQ0HJW+l7I9rV
9LTSgVE+0R3C7tLKWBtL5+Ay/ezi924iejTIrNZtW9tICsyakOU80IBQzyhhCAiJ
JK1u3oPKfWSU2d60f3tnXGV3vT1FPrY94FOp6TkRS2hbLNlUXvZq3yu6w3rr9neY
F0Xb86xxSnq/+wyripPbg4SUCJVa6hDDfOgNqhYlRXZGN3SBX35ilcbVd05LBA/z
m3LmQhzV1AZwqV46+objIGrthmhYLGcesjHVAKQrAl39BodfblSRgI3+m3hfGBCz
EtgpxlZ3aWRr5gqOr98hl4aXHAoXr/Cp3iaV3mNKF6c7qEDEeVe36LVIfOUwxPnp
KOF5Mq9dyOMiLgOYfm0uVhcv7rizsbOVhJFcrIo507uuwwncwZkpidpr3lA/1Gv0
hNQsEm2APewJrfYRTytabCN2M0bnqrBW9PZUlzHxZOKXUAfVo/v8a+77vZSzprPM
iRooDS12YR1c+gsdmD06CGbXQO5e6EBdcl7UhWx+jYVIi+4QQCsfDutUF7Ir3Rkl
h0yEkXPVrLOYyIiM9lpb/2bxe+5a3ImRKlI9wU6Ky08dcUVHu9mvNLmleyZ2J1e1
qhGiYkFELn/Z30m1l2M6j+3FMyUZP1ofscEdHv8fOum3TJBHYDQSp3q4+1cVoEzM
yR1h5DZOvNRzlpXpzm42te8S+ufKmaaKrX1H20gkc30+wP4Krl2s1nk3rDCsoczM
YGz7JYlfkWa35EYqcqjNoJpH0lun5QXvRc1q6JEZpa7FJA6TYiR9b3US4hzT1T+F
sMPiMS9g7dhaNk0MpY0T4OdSJ+ivAaDxSzynO9Tun4b5DIkZMKlEiQZw9NnzB8B5
NN9ahFb7cjEhof5ba/XOZUFlZ/Gzm/gx03DstdiJ9larUI4h8Q5M66AmX/E5kvt+
jkC5m/KDm0rQCIlSrXIb3nG5jkI1RQWEA6HkoKcdCYhvTYUNgNVSA8246RrhONgQ
xjWtDeflbjSpRuqojKTK/X/5JjbKaCS9FCdEmS1DmWjlovKk258h3FLZ2JCG3Rkx
ma5KSsCBggXc3570VB1dHy6DNFxxBXto8lQdjZjXYmIrnxyitc4jdgYwrN9mtcGA
uBu3E5zUhQThhwbyIJQJnsdHb6MEsS3bs3AvCJqxUDKcn7/J1loOoPhAbqI5E0B1
XLhyyb26tYDw808hjmn5vRkY9C/Fhrp4m8eA9Ed0l2dpsHMryvSfqAOzxT7IYAg4
kMJ3egUKcUwHxmY39yXUt1FUV3ticeAJ/rzSb1X5hpjuBKiQK986vWjoKL9TZAJr
mZsITwgfBNSWv2nTd8R9YpmgEDLvu1t9Ee5KJEK5c2sc2Mn3zUW3dZYjJvsw5Sff
apfYpNs4WC4/IzO17d1TDv8tXcdhikFgWGLSvlDqzSvJZGnqOhd28q441dfRMaaC
qq1bSRefELGwOcBm2topEhjUeG0LaAdiMgHlwC5F2maFxz4SQ8daOl9+NzOXAkc1
I/fklkhqePX6Ggm/ZYtsICdN4aX2SVcP5fmyFjXd2olgV0C+vVk/UxPSUGV9LrqS
WPD7JfzMKMVqRwV2bxdztkOF6YV638z8U6sJ2kxbXMrFXWQYPP+N2vOUlKxq7MaE
Fol5/JhGsRKnobOVSLj+XnffG5OlgRZ8k/4nwx7ymh/p9ef4lOt4fskFlXI/SorE
ETpAcCKDix8zeH7N4V/myMwjzBY4hwHLHOC7BgizDUufz0w9dIAoeyTe0Zh3q2c2
wcbTy8O3ki/OHYHfp03ANqC+wIDhjx8LmEHe3zbNB8CgwZBzS3cMk3zPiAb0oUAb
fA7e9ePcfCLhqn6cdl3IPus4COrUKIKNribBThnn6/5dT/2C9IiSA3kXbhXkbbQH
hwFsBp1XvohzMMcI+feiTjMHjmv+BUb7dGiJ1prhDU7f1JEYelJi9t14TmuQ8Bwm
LZcfA6e98SuC1sjF3kVZ6qqjZWZ+dyjB8P+wS12WKGWNGa7X71q1VCIGzP3rG8UO
TeDrCeOHvQm6z4VLo7cqkMporoM/d1MfJ5MlJDXCauj2moqhP2SJhQmaDtnu78xg
JfmUtz3qx8Z8WOovSJ+liOQX58FncJxJISkgnGN2ktEBqUFXDfUAVTTkJsL2UZ5n
ykG1BALeXXeETcJy8QwQ/qKo4ZMMZZ5046QZpO859XUsqzscS13nTsBQABJ4F2yy
uQtEMHZqp5SwgBWNqsH2A1ccIiOh+54fDEmZcVqwTQeyUoT6tkCEELK7mgQtqWS9
aMLtWfR2plzE/7ldOMJA5z1VlimLIyCt8FL1aaMKgL+bYxTWbKrJjsIGoYKsFsp+
doK+/HMF1qODfN2VQdGaBa9OZzlNFqNPRGlVbTDyDd3j7wGUScfmqmwOthcWOf0L
llS2A8K0ZRgfdPPxS/6b3V+0GPTNWtx8F5k9PocvHAUnLFKVYcbGFiEHZpbj2wQ1
nIBl0X45SCGgi8VAtDj/TgKo6CGndKnVxjTueVbvEMU=
`protect END_PROTECTED
