`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CslKflE131oXyj6zOa8Xg3WLLOe5Xb6E2ewkWTmp5PfJUBP5b0tV4Atsh9gHyIBu
QtlKQyk5i7sOOKQ3/X8oa0GouUP2lX94z7j9eRhgiiHSrbuJvOD2l7v65gRx5wlA
lcFdeeF4tWwS62mvPE79dcSpbkAUgE5BZZN8E1wK22D5lL+J5q2/FNAzve23YQ4t
tbjNYq3XI1UX3W1dkyZ0a3wDQGTohp1faAgkFi/fZUe4qZGEPRwQBQDGsxQGVk5b
6dotMCmjAxCUdTXpnOuY2GLVjXNqjei5hfM7FnRuKLJfxx9iARJFMrp92G9+ajXG
/uOz20/J1SbFsDWlmj4H5Ybf5Sv5ARLk3NBkYEEMgR2uTrk5o3dtAWy4w8Ax5kBk
EBwV4dcMmiv34jL6TxChFqjnim85KBP5PiFgjHpd8iRJ6vfLHTYAIanNWzLVnuGy
LlfUqdQJmwDwqPhBqItZg2hijmnh8unW980MidA+YDUeZknwJyZzjNn0Jl7OyzE/
dCQFq42OUM4ygqFB5T9m7axf4hk4fARI1B5ytYnLdJtXUGe38vRlXNf1DYuOE7p6
tP1EMxRqE2JBY+9qyd9HkupJcHzLPvl9FmkzgWoypHd8pYMhoJmTZEsXNR7VPLUn
zdIsaKYo6LcNYx/RH2e9gopGGtaSMGYXXy3yU9eXWaWEDJkwseUBbRbhfLRK9Ujw
zZKeaxl4DFSLor4nbszhWFogtZ9s5o9N07nvIjJKvz52tVcYk6c4J2k4LN4e8PJw
LLIRgtfjhR3Sny2i66Nq4HY2bou+A5sA2jvykzhY9rc=
`protect END_PROTECTED
