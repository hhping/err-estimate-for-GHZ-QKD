`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BaNdUVWF5TxuQmYbwDvRFJzFS6U5KqCs8H1tYH+B1+oO5N70zrLpexJZjXfqSw1M
WTf/bo7aZil0GayUnrHjMtBFUcriZ76LaP8MFj5Pqjw4LM8g+RaUgE6iIRmQ3AdB
QGrLIDmqVReHmoNVulwcT4bxjpx7ZggSsZhfpxcTW7jnhc00VLcA/1+D0Tt8sCbu
VfzqP72bHu/M70WE/Kc0MynB4mGLxw5kXBKLcalMa0xHm9akz0gxVmJg8xUcR4t0
qkgJD324+yp8DEf6ZTqY4woAY6kw1OxQQXc/UP0MUUIgGo9ko94vtlHyUnPBQGSm
SljK79l8Hdm9mDzxj2J6dymYarsNU4iFjEPj29uMrTqZ+xYlNQUQrTEY5wp+13/0
VsR1Hes/c39w5d0/7DyTRs7tc6dPLXVhUxGqK3irGVlTDErIbfwsD/OYM2dQ88pB
tcjiTN/fELofQyCKh7IDcP9ZzDlKVObvwSuAK3S7aDX9cgNRWUQJAU6dqPUT2mh7
FH42DUXsDZnoDVEQhbssJHvVawRTbmNdHakyOWSq21CLnm9KBdX0tJ5H3FIwFQ9F
73HyQ7VLKQPikPQ3PRfGm9ydQmMS8dkl2u5fnCzdqiQh/37ldRFuanFg2Z4a8K1p
9AVyRFAX3+lf/utk2vsNL6v6jLI3oSwO8tHWF2qq4iK/tZckTzr45MwdkDlQNZ8s
asSiUO0/+qxHQqVE4tbHcAWycwotpxaJQOu73LZb8h8B4zVm2C+ZW2d3LO2xsXLT
7ju9aoFpR5oDde0vpCpv//DlQ3PdLsr0kvqrXUp6XW8o0CxeO0xL35JmICJ7oVY3
NFfs/fZZM5g+aUwTaEZ9vv3AHFgpmmL+JMUwi1QYKE0D2c8BUjNsFf1b8WxllSFG
g7zF/BtZROUyfLKIjFpnosQP7Kau7L3SVgBzSUFPWGUhnN4pvvSQM6+VggezNTSS
TT9zTkGsZbE+YScOcM3XSaQ01u0pk5RvmMA+TcgH2Mbo0Yw6pxeufZT+MY8AIX5O
w6wRt05YTnKVW4YghsHXVvT8AWIpQG6Bucr+cuILLI6Lngc91cEBGsu0IHWSx0pW
MRLq2uggFqCbws7XKViHn/nXNrZCPJGDxCx5D3LbzeOnfqu6lbQnBC49nOIM5LxI
HlUN/aFFUmUKLf1zvuU6quctJEZ1CUoIvMP5FB6hEDBdQHKKo2GfjPYgFphxqVUK
AUh988uOKJv2GmW/pXpd6Rk9VsKyUsEf+9fojGhCk6+3Vq/3whfowL0TXI2PXYn1
5m3T6h1FghodGcizXIF7G7xXLaPD2dlqDuj8P1hhSzEKMya2rN9mchub3F83rGmS
wz4AmwtV8B2hlsjltbrp85AQ7qMdKgWf1SlZrlCLLZzmNSUO+uZHIBdtQe8IDZy+
QGp0+OtbqNHVaaMJ0lih8kcuxWfLWj0J8kRLGYZbytSnoePTNYit963RI/+mb8I2
A7ZtPNAHs8hOs/Jy7n7ujI5/VzF5s2oTmCi1wYbHu2evsLIagE5nM5RV3CmkfiQ7
UnNni2tG4y+6fiaGv3FYpjwoXfQHVF/W23rVb56r39ykk2eC44BpmmXPwsGrBFwj
0zvPLrKEdFiZFP3KCtQrf83FQ8wRKHEV7zongw950jk4hHc97Urm5Cnjx/VkFjDg
XkFFumwsHCvwqn7W5c12JmhT5y5v3l5LNomM95Qys7wsG0fJhUcAEJvx9fuWs/zr
VJNNpA9n071PFAofNGjOEyN6i1fD9TNGWiKzGvHM1wOI+5OOtDwuoEL6owyLrPYZ
vf8DihZ/jZaeWlX4dk3h/zkQZuXHOAaJ3K+/pL212piJhacdjXgYF9DmhkfKap4R
mCeUzxjeDZnjkoLTt/rD5pTQcwMnTCIfTtGNHJyRUBA6pGti3nWyx1lgnf9zYUFv
+2yjBagszdXLbEDNgye09CQ+W1Tfoi4XE4pJXmhSwXggF3ij5YuHXnnvBvnC6FnK
bVz8S68NbeJDsMVW35dvobt6k+eEvLHBEekhe0ff+IDsb2EVL4G6bSeIb5nSAZgh
rQrt+SbcRIUfDBKq9Mr4TpzTPyNiL3PrSKeaA65cVjRHyUVymYhNxP7COxvAIbeP
NdyRcmPJKBTiTIAGdvqvQefcq6mD83xFundCDppjEiwq4wML3YSHzplGcKqiiPmq
9VlfBbpXiyMh7ga8Wz8JJY7mnHCPZ6KLeu0BpkdVEf6mBbkPODFH4Uwtz4+7wxNl
/i8t25f5KWw4YbmYKSQx8WLf6lLhaBurFWN044yQzuY73dbvxPWfYJF8bLbjB7HU
ODvHaXg+I+zXqTjqub9Pb3xS9qVKvduuZtgbj5aDVrTP7JwDoZhJH51bm65hDUjL
dcG7q97nm0k/icGs7XMYIgxmOHdSBsomJNpaJRy/GVFcnf/Jg4YQuZp9uYwBk45a
bPKoF+zVwECN85+0skNaMq6Gh38ExzjmyTyZHSwVmB4sSPdHQ+YCNriHDrs19x6L
aX4nnIiVGt360/FKTicJKheb+2f/Dfz/i1lpAkDam3L98Q9IPYsKLc+TBg+SpXl0
F/3KmjU92Q5lRE4aFtrmDGVM+jJBh8srFLLxALGhz6YJmttfbkPGmM4s/2dc3Nrx
OIzL02i+/7qPw1qkrFgXpMnrE4faynneLEh6QJ58hBEVYASKCPC4ldAU8Gz/WkHq
52UFW8Cd4LgogdIiPSdaIlF1DrosP6M8Z8mAD54wObaCuM9GbAoBwRIPJNPlgPst
PBFJA/5ieEkV42GNY98Wv+xzRIU/D6+EPvH8PI+DXoKgBQdq5mnYNYJKoCoM/6Za
CL4jxBTK7PYOODH43CiXmBRy1IbWHnmy9Rtsh+fxofzy1+jn7PLDr7LJ/lkm7P2b
H+VmBW7tJdnKVmMrd+VtmmKCjuZvhX/JLZcY9ud6CF4=
`protect END_PROTECTED
