`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RHusrdJ7czBPoPoOtNiUkF3p0Saauh3QJGJ+Tup0D8R1A1SlTVEGY9HgkJXCu72f
Ov1cVmly29RB7vG7hci/egSnYAh14hc6nCLttO4MRd3xmLKikyvnsUTfRwUknt96
fbLRgDxpCEqu7/YIkQZrcW8WNfi5F6ZS5hyr1UxyOGECvZ9KYDJgKnCWsD4T2R5O
qgzTUHcrgP68/zy5Z7gW8WhNgiw51gA4fp3tfibEUnXrJjuI4vOx7VJhvNCzpptQ
OXMMQmj9kDtYrv15Pn2GD11Cop2s/KpMf6u3Uv8oJvPRD8F2bDt7Qwd2e6IEKwmb
2+72IqhTYspGvtSn/zmZR9AiF1yD6+Hnv7Eu6Ec85xL6P39UIgQ7FzVLWOV+zNGm
c8ZZszaJ18kyD5EIXorwpxjMf4KwmLpw5BcBU/f6wYgfs/vypb2OgCmuuM1kmtEJ
Bvcn275U+h6DPZHVfTXhzMcB8hLGz58rgI4Q7sLCKXfi55+3chZaksiWSkrreHcS
YK3LiHPSHp8gBxw2H8sP2geLF+P4vp4TTMHFVn1uC1Ev4Yw7JujIaHUMUhWef6Ei
r4LkgWuNC+GeJ0yAWSq2iyTx1x/D1/rOtQWQFriAsxgEoJQGJt/CyQh/OJHckh+C
vJObUZwjbdLdYw+M7V60FXXns0TeasBggku5WZrReOtWy+0VjjCHXlPQW5taY6ZY
gqBq39QBed+RxEjblRmvcvd3zh3cHsIW4i8vVi8jLuE+SB7+VGilhAryDhKyM5hF
xR9TV7q5TWNYUY98RgLWy9CJTIvxzD8L1AKJypRqJcQ/FUEz02wDMBFiwvaUfdvE
`protect END_PROTECTED
