`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EfzdPPklouWqxpCEMPEIZIzzRS76O63cG+OHxWPeGAJwDVVZKyww3RtgU1AKPcjo
DQ4qZ6eRA2lEYHGwxgGYG+EiFdJRn0UsHSqrSbm9Wom0Ux8nM5bP41o9esw0X7Qt
lPYSovsG06zxd3SpsfuFlfcPHpreQFT/KaL2k7O1ZtsGWSwZ6Pc4oBxQ2Lr7X+KC
lMGNnnvv3sDTSEuoVuyqF/liib6M69i9wm/kJS9LkQIlHOjU6z4zsvW8PkHOQSRb
wxIbFXN/uf2NktvsZKTAPGK1f7JjQhdHkcP7w1id7BFLXOKU1hSf2/yshswZjBNj
lmH5igwPVaf/CjzVfLnxB343N3lTe2/VYQqYXJ+x+Lb6X1IVVP3bt1nOnDkBmCzy
MUaMVTUrppN12v55FhJ/qlbzyu+zVjPOmx75WC4GYidPCbSS9+ky+aWvhu6j00om
UJAnZTsv5xhyDaHLX/uQvAqrIYXB9XD0tUuKJL2s0PJOQCfRT0BsNOoZ1TwdeEiD
bqOsyf3b/X9EFDMs1gva2dToKs4eMg1KeSEWIEcuXYVzDJKFDalVAMyAPd/77Iqg
ev13THu6kUKSYipzPMjB7LBv4Wdcf7dJUJneZTAK0Op7RVSZFCGJLLQpGHgWYLos
mcbwldi8ekX6UXK1rrvuXyFynBJ51x6wVao10XQDm76sDnF/gtgN4zvaLbjPfnm/
tGisWAoXAc8zkQhtcWZD1OJcZTRKwFRPg3vjHHYyh3EQN0qFGC+NJCmSHNapaxpJ
uunR1ZHwCMs/JNgmkwQttxGauX0YK1UQsay9QDD77oPE7SRfn603WG1uWz30y2Bn
`protect END_PROTECTED
