`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epxuHHHYXuCTFVOitMVhRSqR4MfUHslpswd+ZJ2n2NjgZ+zgobpAKuyqGGOptsgK
yLhoAgld0PEmwq2goUCFmvQM7zGRWA51Igz0osX4r7USbdS38rgz+hTFdT+a6WwI
G6ORHzddVPh84yEfLxErhoMxZ4bfrNfIXX597ECLkhrwVsy0cypQvXHC/o1C+9RT
sX21s7iX3kicWDLGh10AsjLkTikbvT5mYt/CmAQaMO3WqWg7ubp3IdPVJotaz7Hb
48xOLJNyX6vOfTjUEN3ltZ7g/qYPFIoZOdS062g8sTE9CWXWJCflRe7YRiMXRDj1
SoZ9upj0NYLSoXY6bmo6bW5aOhCHn2L78ZxH0GGZXzFCKRlxtGsu05hG6KirqMSl
Gryt2CzotCwbWAVWWVQFQ2DyHw7z9NU+z4BEpLKfaIkvQw+Hz52UoU1MfvRPPyN2
3zroajDQCEq1aJsdn8f5FtMFbiO5GOR/FfYNWCd0+BzJrNLOvWX82y8ULqne41qK
jxy9lMzDo/Tp6+cL62GY/Qor70qwrJgtUAan5FlgoynaH+9O0BjJXN6Is6JI2UnD
rRnVmtYuQE2Rbz/Fy5J3u7XXFTF5RLzDmDJEU7bpTEyRkFjDma6weNo1jCzJDdRy
rUvizKYRqu8qcxCy5qVWijrVC+zvQxa9SNACH8Sd6yH5ziItBoiInujpJjQ8QdG2
INoq6anPHA7JN1C6GgvANu7bNgud9TtehkmIVaiZQjMWbLCkeSUFBDjRxpv9Oznp
IOTu/L1WEwrDug3jE46kfvh6zt8Aojwhv54MOHWG/Fuf+T900bjAdb6Sg/3KTbQ5
ENWp4JXWmDXIq1UbJKwD0p1186IA3mJ2kf3IDOHGGzs=
`protect END_PROTECTED
