`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9Bp4rIc0jePXPtx+/tnu+FxosAUVM+FZ2tdw0k3qXG2fRSrURrrOVSlgrV+OmHE
HAuDKrC5gOdFAgIJLmkNA+ppK/MiV1HA8/lUd/N3Up/HwzViZ+Njyfl8Y2OIK6C0
a6fmKDlioGfuxjYBO4w7SRC/DhSqBLBT1LSD95I7qqw6eqIcf+QXQYZ0fxN/+Kbl
hy2lFHoCHMHTKA7p4g1JqrR5zQD+u5vtO6a4UoXalpQM5TLPwXfDYBVFM29mAIUI
h4aoFyt+5mQ1UyLMnml4RHL/96jVuzXvTd4zDNE5Y6/yp89IDifcLBedq8hOvy0g
IhhR30vp1snkkCuQov2UbhSjx8rpktcndInRVWENsIkk2yZRFb7s1O4Rnr7lDfht
Pon0rdX05AKQ+pjfu0cCkQvq+trlNr9wvhcChNIm9tEiJ1J8TBc4M2HXraUoRThN
RdK5RGPoSByUGSfn6hhXSiPmdOzYyTKZ9tWe9RqdGUODOLz5YFD+cpmbKgjt5rxu
wtP7reAlPZLmTSyHMC4cDMpVRX0sdkDrVxFa6cRgYzJrF+MybMfMU1xVf46IRTyt
naTsH5hE3/lF0Yc71GgVyhgFPXTTrJzMNvJpEGh/DfBx24Z89EethLOx0EI0z5Cs
ChbXKZ5nUQcSnZgX8ljzSK1jMAompVSoozPbvnXqprrDCTX6wPIHIOQMY7FFlRhP
9hWQUMDp7NZZAhNAS/eQRrxA0mU5b0TkqYf1YijlSThDOQmXdOoqwCsiPilx2jt4
OUTWHBH5Yf5tNb6vV37kTKGklWn+HnbSQK1B+fMZYn+zqChPhU9nu4nf3vBMlxZV
zNd2NYK2jOx1C76GkI5J0C8Ygr8Y2A6q7cmsR0M0JuQftxC19Ue9836wDpCYvDPp
mstg+tEmu9AlUSnKHlkHvqBdbCqu3QXvQMjj/hV6sglRKTD6brKmy4b9waG0wOVx
KZHAQFkjausUAL/NCNC5AC1IdPzWeY99Sxh3hzH0mDF3FI1z5HIWRjEmP3J9GkeB
qM9efTdjuoYUQbr4nq6YSVFmnjaZk7y3XIZ/Gro/1zTKqRNofjG9EYqeqgL24gbz
50cRep03zpxdOu19wlz2oj+FA4DxWkSxxhAo0cJUX1bULT7RepQSD0l8LH4K44Ey
ZCb8N2mRCWWb7/05N886/m7JTOh01TLm4Ss/kbid6YD6gP7i8vlvQvhTylgDUcOI
`protect END_PROTECTED
