`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQKadCKtvic4bAbP+WLn/sVybCKcdYcOUOG9L5stuaPJeOJeTyB9kqjtFxaWfevi
xIdoDL1LPskbRehLCyok333/+YuIUZfdwywu9VgH7crmNvYyBRoZlL617oxfUbso
QlYY8Z3JDi6OgDdYUl/daReSgv43JrypBTrrUgGjU0FV7eV1JdENQIKdS+YY1jyZ
tlH+1pExWeZFC1Nkp3bAImRXb4eOXflhZUI9Ufjqa0Vwzok30acX0DgL1cIndrQv
zJjDTReKe5UfV6//muj8UGDdAsIU30n1RoVQIyO/D6hT9Rz+NTyuIkIUFlnKBVI5
RBACd9OO8YsjU+G0pciydGWnyeL0/0brIC+IO3o2xrYSp19mOHOUZDTq4fENr9Ul
lsGlZ4Z39KkBmeOV6cDD3pEXJa70HUV5UGQM7Bar93A5ZUvogNk75F35D1FfruWD
F9IncLFsK01zHkU27IvecoOaMq0bmG6pW939eLgk2FuNsR2ql6HiVRcbcnxQOb8+
iTPboakBPCgaw71NCq0oCK1vu/pJKMWxtr4Y3Ylip5NpLWd5NPPPbOY57b+O9gWt
if3Hp6RyRYM0dD+P9RKHVnivQ+zV66fFVFIN1/5DqO1qrv9E2WEbpeXXh0OeVYvs
hmBl7WvVveJf7/Jw6vQm/+l/wUGH1SQsii6ooABLmns50ipJok6+Z6SMD2XVdnRk
dPMQRhX1YUhYrUScNW9p8L8KsbCj/9yMA0edhe3ALT3E0jjTn3HKXerkF0vPO6F0
DnExbU26xx+q7nYets9GXzjMvmLMgXhu3vm1ATY+bIZa3O92CtTg8zeif51zrug0
c3NjMuhwcWlKiqtbSEESg6CREihNN56i50RWa7MpUnkwg8Lyn1qgtvB5SXmkvPLA
9BObmxC8rQ/K+bijQa5K+z+URpqMrJlUnvuvXnRbGpZ3qmqv50x6V407/sSbSPc2
XXOIZ+1zIHlTptEtWlMeyPpOIcViJIXyFg79wgCiPPHQOy/ce69Dajou+wZpTTFe
2ehu/DHy+BNr9+6kVWE8DftHPc4KpnSlBdya0+r8peRV8DUy809K7OQIJIO7HMF4
sGTKoBMWc/g4FlGBV5F4l0rgcAV0Kx0iDASg7nNAKI3aEGPJdkaaoXCBahYB8DXk
yGQEYxptC7mDMBT7h+7AK750Logy72WoW0bTZKRau3KEI1rByjdK4nzN3oif2Ull
t3tsKXzNr7jTAb7w+OSq6UU3/Fpb1Jq+CCJFtB9uS1jEAHRMWcUOhTld3iV0Ww5l
+FQRqHjCeKjKyNBPOTsq/HUYdbDwXWlozuGLVQeXTEI3ekjOMIJTJnIG4f2k39zS
YPKJWyI1HlG9l7ADefj2ul7i3tKrht5Wk5qC4TuRSFuiLDtz+5JHsYXJgwckeJpk
QhYxJEdYDiPnQ0ce45G5hqJ4URgHgd7xCZ3CGyJky1EGVwRp6VKI5YA1Pg2aw02J
iIavJhz5SubaW/vJS5gwBZOLtj7EdmxvDtKb4172Q3yCMgcEHNIPIslTiLWqblze
SsMev3WQjQh4cBMXNOq765sPsStNNWbXC5vpv7XWxywL1eJGcScxnZtbybPpfacR
4CemdtVIO+e6LrBu9XHfBK594ccXo3jKUELKU6ctiL8ceGl5XdA3fvgv19CW4LZg
0TJidiLQSeukmFreebi+sSnHVaL7dUsR8J5bzcrQFjPspm2x4iNAtuKLYokQtuZD
DpW7bMzdLLULm3MFDvF3mR2w8MnvYLSo+PSIeAfHtO4QLSf6NsS2dTA925EI8eW9
ovEhZpG0GxXDuw99CWttGceVd72/2by1jMCpdTeOQrdsudldo0uZAqaoKXxCgqB9
KM1pbD4FmYRYIHrzORLoY4xlhcGyU9gpeaeY1NzODULdKHvLVNsaAMb0Cc4HKYt+
AUCZZJAxInA4I95Afq/MoHhX81CEhOtv0TzkW+idg2wxVuD147uRSuFmR2LPMkRq
radi8M5FjZk1yPANjFaj2tS7r2r9O5bIUrsw/GpiBF3pDscCha7oe7Vpancc/OS0
UbQivIshmdsvL9iabSNT7TflJ3DDLvI8JA28zPw87uxbEXtTBoPrLRx3mOrYSmIE
AddlHjRr6Xf73Zpf3P3ddYBW1uHFz7nYLK2rJTerv6dKfe9ScFe3BLQYPy/VMRhT
6fgaMoVLo/czfyniCxO7rsJwTvMeUWDsPQtUQII/aP5/Rjv1En43lTjbgrc+IWnK
V94LrjmVOfkkBalLY2MHANhSYoQBUHt923mFGTqIAxp779hvMmtKsGpBji/Ztqsv
w4HoU+0PWfFpm/2squG2xw1stR2Xn6PeiXFqiCtecr6xnoxbUFKDaD197/nFdlms
DH1KTf8SCqg1qGbO0t2AeKZY5R8nmEHbX89pfSyzo/j+/mrkXwed87rKaTVzdU49
stMeENC/jiJOQ26qebPYb3m0gCrvOgif+u6UdQWBb5n68lI3Mrs/Sb6+U3C8Ar3v
lPKR5WEEx059STmdbrHxhtoGzD9IXlBj+BCWl/+mGGHkciP90cclMI0jDGjmEjyC
GfPjcwEqSN2gVk0/pLaZXzFNCVJoSy9kZW6AX+HOF8/sPgbGKGAQeQ/lC1MT3Rt1
M5Bh+4NVUxu5TPU+T+0pjWieUnp8f0Vk4jVqq7dw+iyIvufKd7u6eDiryMsm+JZc
OAbJsPMLi4koPwtFNaSSaYIB/R1f0z9JborufzKl7iTzVJM1FjkaTq8vkesIX/g6
60AohsIxfr0A2rD75dgAnOYfNkNSAwNTcmYyePvaTKIX+N3I+fG9trP/TXzoxE3i
7nelu/ESVJGjP3cJS45wcCP0XhETWRx+iyWvq3i3dgCVmsJ+dXClEBtVY3p2ayOB
l9OKogU60+Pd1qkMau1+NWZQqtersa6NgagahVA17xJlDnr5oknbbNV4ogCb9DoQ
+JpAttc+RTqMFOaHf2EIxYkQbboDRmvr8Vg9r9E0TkXYheqWpjN/vsSeOWMFpXRL
URAthBW984z2fqdbIyaNxst3Ht48/yTFXjYLex5r6PIRrqLjE2TxMYSivY73d4GG
8xgbEAvpYFMW1lGajGXQdZtj3cGK7j9GUtoNNNfRN05jrehRtNSR2exHxkOGzpOi
g+EZkBQIPAi3edyz+pf2lD8JL22u+/0zGJMM8+a+3NXW1H2g6KJOPyGjOM4rFd49
Jpo6tfgSOXITCGCLkgwS3h2otp4nkCryGsgypvUxffe62/1+JTQ/0wuYZbV1surn
4tSrllTpOI1VmfpJcxTiZL8BSEweNMyqBbYt40RafO7bSC6dxGd+oZx//YlM7q34
FjyKyT5Gql1mthmC5Na4IuPWZV384dB1NQUOoWEONp8O2v+qGvhzLKPjdFGlpwMb
O8sWzJClMNLNd29L4nBJPSE29BWv1eKkVbPKq8ZKhTJKZFPt1Lh3EIE7WiaUXTCP
i/iits8uoajRLon9eLWAE0VaNHgl3We8Ob+gwc7sSk3F7UWP0IqdkDAzBajJYLec
ROWhfC/Sf+LhCIawaDbclH7Y/xsWPXiPhifr8fvcoO88Y9zZf6WwmC7LcBEQHqkz
FDIIO7mp1egWNprqZRDLC3hYow4COuHQiYedrtVyiJAGGZM4c3KqcdVOoAmbIQBx
+05zhrnAN0z36RA8ZDl61rh4LtaEEun2TMKR64DLI6XyicKuDxjbNE9i7tghdak6
oR4pD+eUOUe2feU3Hsc5cJxoISIfiLOTPeR5gQ/hAmGMt87HUk1SeoQKekNJf9gR
BxnyUaCDExYq8orXXGpbjDOiUbJ02Wh8wEhAV1Dg/GScnXkltRJKXC7imaxz6Vqu
04ZS2zpCzAfkAsZN6Hb6WDs+fVI49sKStFOvrAWgzSe5UwVOiK26rqa6/SN1cr+S
yozws77TdTh7BG/ARsiYRpw7y1mCwWI+7bgU7ZsXg0SIVpoGCE/p+XmOAM0XzXrT
RDKrLY4oGPXyqUIJVBar9qD3Kd80+xCooKzJw/NN+XVTN9eGn++YoP0ntK3jd1A8
+4wft+G5GI4nNhg5lWF/ApzAvG/TaIa0cWzHp8HOpN77VQxQx3oS2r3ScGslydM/
mQ3aqR8Ft4Z+68U0YwZlvBV+HaCherDs957QYo37RdnYE4yo8jifWXh4BzYmbIjx
d+CAQdddAOP+FNND4b3rx+mu5MSDwSyZyW6bA7V3kT9ElzwjDSLZr+kJSzoRMKCq
xFnZUG67a6wpTdVCiLHDeibjpJzwJ7xOmEjpYiMVACeG+gKk0fZx/2+GpHcnF3Sd
N7Q7NnpCS3YwSAgQtIctw0vOO6enLr4F+iBgSu2jQBDFnLo40MdtKbweU/5yg9Hv
hlggB+qbzBcB+tpfRhnuZL+2bOIMFvOhKeE6Y3KsE8YB+9xPSM596ZCBo/fQXykD
SLoDxBSrIWgA1iON1UguvE0mFPsNh1l0amPXY1Cv2JvqkYMdgwXhXddcokrOmGkA
KwJRbBJD7+JqJB1w+TOHAP7UWoKftNmTJZXntvA+2T7hKnDBrsWTRJJxa0Nk/HDV
RiYlnwMWNyCa9TrG+v0xOZmYymjTEgESJ6Hvi4iUMG3gFANDoZlXx8PGHdx08PE6
fzc1zujJKcynXjs1R7O4WQuvlKv8EnrBI41iM4s5faaEG7qBXSYIUE1uTOlIO1S6
M0e1uPuiHzpZvnj7GvTjedSj4Dwr7q5OE5/PawkyaQGdwSdQY7uHc+99gp2sdNS5
TstPlXOLw51pqwN5B/NF3asF4h4aKY7l3M63wnI/rZEj1yLwYsIZQRp77Sos7jMt
yRrU8trlr1sz09Ctokft/id0tbhvFU+Ntnh9HOUWFF4b2A43d8blekfXlqQ7jfhR
nmNTwHFTYG0teGq+hm1/rlvlGHz4Iqf7n+TAkCAmaFH0FZkX6GcGtmoGrjaES4Tm
FOvfXoy8+uHPHg4x5czHeaPilNqvwsQC/IGBEnniGYs/q+d57qDp2yG9eMnb70FR
b3px+09n9fC5Q/eqonOdegaRMZyLOc/ebKb6q0VM4KDiDQ0g1xOx1Bg28KpEbuky
yOt2R/jDotZ4m0X8si38g4igHELLdO8Z10wB8TPcBoY9graPVLoV4jmu5/voHQhD
l6I8HtcZfQQBwMVKvVbANYOnc5qrMAQTntx6MNKAbi+d+uIML/tg08chbILmbchU
okU6w62iHVRXxtzQHkXwboYHcRzIX27cX0Ri5U+Saw14xI6Go5bLcv0SI16RtiWP
upZIhLw2TWk0E/2+EaatQAugXwg/y/5CLGGMlPkbyUTlNatGnggHYQkFGsGPgHuZ
oDXZUas5YwQL/6JumeByqMHOeMaKHmwIpXZB1wD9/8Q3VxrABIwIGvucIexE/gjF
v9gWjElmc3ukTgqHkppsNc6kaOxnRBdY9V6hWP7FvYtPL6+7x1RQ9g9dAz4z6shV
LLPgAiA+VIzljoRYinwb5kDO1yLfWqAB67bimCbeEHBUJF6Ofya9zkrrVKVX8kCJ
+p//od7nnRX/hxW4tN17dZGgu+DMhBOnE8O1zHy2mrgOlq/EGC+ctXTsZiEegi/f
sV880+3Up2lS9r33rLTMDgX1QfNjHcx9o+FQGWpp/8dByZl/7/rtwjkM96ATbxEC
9Kvf0XhuJFqSwsUM1Tf7R2cP12Emp1HBZiWgF2rE2WNa6vNtU1YSyw9ZjmudXPdS
/GWu14fsqBk8u7o9Q9UEOOYBnLChHLazXAbgiVvtyLFd9BsoB2C/KfGj3pq12GeJ
SdD9BzrZbBEaAgLfhtAA4VtYLZawOPJ+Ro3kVqfeBiUUYhIYE14x6yrTS/OtpY6Z
SX2qqzIE8xce+4Yi4UIgSVtNPwKzHV4/msYWjEMyIK7QWWojvOmqrM/DgPAeRosd
mjl3xL6S0jWtHUOpkd0E4jEsxft7ofRSLf44P8QV5HiFJ8v35fVEZk3Q68UTrFJp
td3wUKUmr/vYIPKadrXYrqcpnQmsUevfQm3fBGuzawq/0MAemKMuSC9TllILrfO2
a9UWiECcLoVSBftNvPcD2nb23NXyCEFI199lZBoJjMyZk4M5VIqevBKGrn0azoou
YOUfQfS/KphFuIfglvO1+pd3a94rACYRmmeffUo0EbQ/i6BHP8294+HccCdlHPX8
NgTJEsbS2wUGoXKp4mQcfTScuN0ZRjfYnO3L/xeVYyW+K8n83pUBnPtDFg+7d7lc
LzXLBuBSeMdpRPspmRz8ZUZoaQv+N0SjlspSC0Qha2MnUOefpEvv2wh9cf0VpXSX
JD31Iu4OSPnThf6lALPV/nlYV9FctJ+pylqyN/g//PStd/3UJO3SViGNQuZFlT8j
IVfKUAykx4ePjPa95TVuGx9d+ebavkWLzA70QUYM7oD5lL6EaH4pfTu87hs1uy82
YYhBzFUR3hFTyYB60t9w2F0eWTNXS10VvsamoFotAYhQLe0iXfktggkJ1Vid7yHe
o/JvgU900T0nMvUvq1j5fapfNgTMq0TvbzTLKhAu87CV1upjlpYgq521GYQKT7yo
KF2b7EtIuQbAeW4zsoRZyzxsyGTGKfImW2hY9QsfDeYOtV749YqLvaO6Od5fLs/5
YI+StH5+eYzRhGkbMPmUJ6ykgDJpTPjLLVCdqzq9kfFnXQxexiYdunIJLZhpmyXA
Zh+ZkF5FTyPkebRaMo6F17ftXdnqi5nGM8OAyU1qEQtQemvmvPwSFpEQKKknDne7
ovObt+kNjVoTZawQ1QQdWb3hYyT1ZXHAf/y20mXhBaSNfptso88lA3m/+CNhvzib
D3EF+ryA30IV/TutcNh1VnYz0JQv82rFHywJplH3noHAUn3gh3N6UJfvpzsZAbta
QwR2ihTkeMxdHuii0dp1IqXygfRx7ZtpvkUdcPNdbpS5knp3u5yihTiHd2rRk/ZJ
qwFosCNgxgYWbSe/I/y+1P4j59aPinsXNF0XCVncEuB7OQREyIcPV0y+C+1XqNBZ
ZdGe6ICRGwZGEC8QPN9vtnJ2yd9wANAhmSTSMKq3WO5i4xDjhxIENvHcii6L1f+3
EWEU7zbpCk2+jfd5icCmeDyeLy1RWtHl/ud40KUSmvoKtpwyBqp1SyDrDn8rV6OQ
8wY6IN0GBhwVpfStJVgXSElc1ujhw7liSzJ3859374xRFSEM1e+kteeIb98gs0/6
+uy+Fc9W7MXo+dc5BY4IKxPeeyIT0NsU3NBBnl1zNT3S+Tzyxr3cuAGPbmzUdnKV
SVv8dBEKNl9tpKU82RrrNbvJdjVwCaqSkUGNo4VvI+NWkkb+y2lfEDTiOzLp53uX
XBRJTA1YEAv7Xxo+NL63cVLbcuXBFHC+4s11r/UAMNDMVDitfdhDUjYjO7h2c15K
RPcgvWT9tgoH4SeRcbsfsJE6Aldr6RpX+wT12abwFIMCqcMQOjzL6BRqG4fdypHY
L7oav8PXtM7FAVU+vtt6ANK4Do6NJQezw42I28It57/VKOOhEfEEe1Bhud1kW0cv
QC2ABYRBfNGPeS04FEuf71loKAlcs1IzvGZhVI8KtN6Z4H+72JX34Jr9EBgYtJIp
TBbvhemeAspdalT2KEKZNRjsk5XydJMpiXvjUIAOGNQFgEimPvuSyNjju2PHrUpb
trPF2C57MnNz9D9dxSX/A9KXjgNGQcG/aiJXLV+fzloTzSFCRNghBKHmNfZiziHb
ZgQcHmismbAJfbj1f3/RYYHzSF1xb8KggjquWvMKzFNSxJ+9PSwJmPC3PEv9KrK9
QqassEC3g7rYlcHXy5bUGMGciPmLS+/4yKIZ6XzU6hiIVL3h97ljEWVoPhPd/Mdf
iTmlo5J1pStl5jUFYGBYfiYIn+9N4IF2mESN6KFZP9xJBYWlbvQIxGX5CYcjem9/
JwFl/xjyTs9IsqAmiQeO/rZF8YKjfE4BXrD3jeJyJY1Wnj6txq4ELoaFtXDuGCR7
UsDL/ZY6FM526FiPyPczvTOpOQkhSQbWKK9e6zcLkjRScllGZZsPNzmtPUjeqC4s
sq5dX0LYJ64GHu51699nuo9gLGE0zyUowVMxDFORoFSqrXHumkI3gIocEvBbLY0z
/8tS4wfDYVNcw0vdTOzCMlltPIbvTyhQMobX+COlLK7mR6QJa4MRDqqofRC2EVv4
XbJ7TQmd7F+z6cnkCoIv9YsvwLdsV4h8gmCGbIxiVgJR3XC15KoBpwD8OqdEy1Mz
3ZJnb3hlQjzS1c/gbEEifA==
`protect END_PROTECTED
