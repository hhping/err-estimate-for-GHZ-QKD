`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uv1UiJ5MteTwLC9GuVU88Ki3lqacZtij/oSjZziDwwJmeGZIHNcRz3aP5XV8uCty
P7LAhD+xKJlZJbFiXRBzM/mXvssNaLw0r9SDTqmlK6zH8P30kGIGmPn2sfBtkcNP
5BsAqrGrER5IYGjWZneDftg8G1aKLRAt/SqyPh1eUqYMTCyMh7d6rJkfzcj/Av5k
MIg71m7O1+Wl3VlqrOdvFj1UR3AV5pAfm44Vc9JEH5Gb9gPcBS0Nx7mLN0LDfrGx
aSs4sFC2iQDSZQmWz/hwHMcf2Ne8hxj35feMiAoJUNqNbygjMH8FtAhH8p2v6mTC
gmAJ7vsFkQxTUyJwdsVx/PCOGfwmyPIvP0op4TLBwk7PHbAhJVj3zwpTWgChQZmX
Ovn9buDjf6zg9C1DlrI3cIkl2HO3qo2fHgBTfs7rPWejiFjdaRxJRqzrvElZcDX5
GyzVJbd92uqIua6tmdAEGqlXfYcBfhP7RWEtaJ0ymu1en2NSTc9hA57hRkkT4a5L
YbqEU6PH8ON6GfY5ow0e6LqQEybJP5FozJZFQbBdW9ZHDSifuvnnzPqHiKm7aX0q
dbXp5KPknV170mvQ7VuoIMlXA2uFqG/gfUimCBHtHaCCTmv68tCN694ptpNsAyqi
JFwGfA9CTe9VyeW0VQ9b4bvC3BkmPERzGBI8FCvNzTeqEK4C+29XZLWqpwBBszF5
Nna+5oZxRlxBJwOqHxr2Ue069aqZ/qi0vAArC/jbQd7ThiW/w5GFkqHuLyJhebtE
fBuWH98zdP7jwRRf5NpVRNVc0xNUNlSF2YSn9LvVJRs8yRv+EHPttU+Gem9ddNjr
qe8epySNIA/6DqUT/kz5/D8Nj8XwpY3J9n1TlysCPH+ULRsvT3eufnKc/0iCdlUH
/ix1k33kWjWKbrpWeSqufgc5gVdTOgLA8J5vUP5IBdatGEOSpp2itUBfuKP5xCbY
/vuAejWdomOPsEiK5yKTekMKa5wHpEusxv/7JH4NFWCon0yEBDqnz571rVdICCJb
KyGxj5mY0pRiGZsqhff15IXv+/M1PKVImDf/kmIDWapKf3JOKCfl59Hh0QVer6Ko
5eWOjl3jviX01skwNxvkp5dvy/9YeBQp6wYkTWsgodKULWPWX9nUDyNOUO2QeF6O
4sDR7m2cw7rbNkvpEWyT2ePc72jmxJWfAabyKYv6NcbvgwNWnBoCKaQHKtt/O2nD
8znic3cHks2mQ1492rxMRoj/pLlRZF1lDASVud7/d4K5/Dq7oml3KzH2GzXUUPsR
KnNa+reqRGufYfbNA5fSO8hErE8888BNRr091c5AJF9zl/bp8k9vajQT772z1+qA
0mgv+35KHj1rAAd9pgXcNGstJ1G8JSxdp1qqPFmVuy/naK57vlib3xt0r0/P409H
Nz3CrS+vXadJQPPiD+m4+Bj8dHbjHpSpRq58vp2YNY3cIM69/2TqSNTEy3lWgSwt
dA1+F4Gg+1Q6avxSnj90jbf6rgUKhixQef24JTZdtVi9LvHe/Xu7b08wXcPsTMib
quCbefGfN9h9pHgVTMplhdP+juBGB4X7sT7F4ip/t+ihL2888t/4mJ7Y5K2CnZOe
WxdxKqj3pVswfovlm9ieFybN4AXmtR/HU+MXHCtyXVCEws56/C3Osr8bP6MjJDwT
QTqF11z8YewIHz+Vopc0NK4581xyWbbr2ikRayk6Y+DVsNBS893QYfXdCR3HwE/E
g+rOqzCJ0qphwuqiSvcw0UUZSlYYvsRXV/Y/ZahcWR3AJbyVdyCGMUoiRoKjFHSw
C7efVKIPxpSiyAZ22jGE1h9PZT6B/+glXh7MIby6f/t/R9TKFxEEADoAxdR0EJ++
t9ZtN5g+HiGjC3uZ78hmICS1Wxvnxx3BVK8U5cGxX35FO7FXFNZ2XieaUWEAdYFk
cb9KAn4R1ZlD0DgQVnvOEyfLaJfCtRBN4gAoq6CRpyn4ZfFXtadrICED/UdIX3qO
8pEGBjDzwrRCwrVanOf6fMM9vlsY9gjqApSIXsY8woVibejhoOvyPv4JC/lHko23
C4ZAWARaPmUfhbcpQeuiLrot6LyVbmmPX80g0Qxiy5RmxjtXuHJlCtmHeETPtrOZ
ySPX0wsY0GcktiuDfY9KsXdNX9HNQYkLQeeZy8ydjWATfFHCOTNNK0BexuNbRly4
m5sX2+2HHLlEdz5u1RzHRZd39nb1s4Grx5lAZ8VfPkurMyW69n9pfKCZeGPJ46PN
12NHy9voikJofZYIu/Ihc6W4aAebpNTdlVahV6VTtLvh73B01VlNu0MKyg6eYsGG
gcUXYZoKGHYOZXcN1FRF2Pylqma5Bp+vCCkOp93Ak100k0ZjfrPFOH7mvkFQYY4R
8l+uXahIjdjrpghks29P5N4Ty4jZThuQI0sSzOf7YcVBef/w5RhV6qjNqcZTfusx
a8tS6b+oIZQVcIE2UdMWqQvesLuRnVIIQFMFVhomrzjeB2LWh0QwHAmo4SWYhKPu
x15c6H6xe7JFL2JoRQxSUGO4fHqDWQLQ8c301Okg0KI/BmtRd4swjTsqYq3ixvAL
XoMAfBrLiqEpp4NVgPe2NyWSdSyvc2btOxvxu9+e1NDTBkVZeD27ARj1VaHxq2WX
MryQIFYxx34IZo0xabnbBTHCYKHPUn04yq5vtnBxu50P82fJyZEQB7qFm3E/iDpn
DKyimN2eGECtQiBXZHuOwjkbxJX7rNbHpuYulltyos48WndFPoUMa/Un4PNx4X2M
t2azcJxuizGSICKUc0RKC9sEO1q8up23S7I1mGkGIDjJI7zesh24bPtL56OngcgU
lVECCf0cjHv7v8hL862xbkDFjbSM8IqkJkhRdiYzUu4h59v/maAc6KE5UHj9Vz0h
HLorgQ0Ne3ml1ZUqfxV68YkNiojBJ4w96oLk5SGjVZ5txhf2Dp1nPaff0Y4A8Rl0
tyLOixIRu4L7FFJaztNk1dCZ68/4F67HxRMXGOqrr1qh1+M6VsDfqWCHhvwsNonY
A6oS486G5USta1mN5Vj4fEtgCTvAz7G3YAAwpDgrKrDhtKBdgfLSr79nu13eUzJm
rk902tnqp5vE3h26R+B5xWP+Yluvj6rc58OZ0STdQJcvK9bYit15kvOj2JfVpfeK
`protect END_PROTECTED
