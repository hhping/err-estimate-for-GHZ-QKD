`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4cKkCcKrahegDJtCQM2HNUxB7ZsOt+lVidNF7LxAZPxr+r66UC9QaDula4PJbEF8
cnQFdRSW/qwe/e3ZUhLqYkEmf70+8DFIRCbe7V7EZxZPiM1X4njR1vt1yBSZYbqh
Eooj8ERidqdn6fw5XDURJVcpo9/Q687ve0c7+pMT90Bu4cY+mcj9WiPIbR1bHQ49
RDuCGguf50nAnzkMqJf6oDvxi9Ue1zgMzpEYMhem+XSI9HlD2f2LRK1NBDoypeeO
6h8+CjBDnr37P013qhnYcoYpG8dsXkfCZHAGNqrjfqT+FOHoIfKsKujKhKnUim7C
P3Bh1YoWFebHkMOQMXnue+dYHKlivvKcJG7gAFUuy2M8JGtKkiZF8XjE+uqErXZb
fBybwvnu9jsxLdPJM+cwYBMZWstPPPEkVi03rHv5Kykv5nbQh0w+o+cSfgl7G3qG
ynfeXy2m0OjlUrAP+TzS1IvDu6Bn86qjJJQatP2wCV2vSfp84EFhEe/vWJw0lHxg
fruYJM8Eah3cLR/WvwPzfxbNGvlPjW8Hx0xJKVilF01VuwGsN2pBQdlfVUvkDAv4
`protect END_PROTECTED
