`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IG7SNmzgmA8K3C13UrL87sU0WZ/MGXxpUXzCShNiSDM6EdJqOGgM9KKgKJYMBsqR
D+86Hpcagb2zao+tCs6z0Y/PriGKAykZdLErNaPBhyihjo+pXgN9kScm8AnM5uIU
ZgwRmTcqJy4ruZn/StSfi4Z/doZVynA/451MPHHdfbkFO87HrMQ1YExX9U+oclvh
7kbpms2jGiybhfJqULPd5n6uq53qLWs9DVlS4rAQj9SNu8mMjudcIhWD+4CjNSRp
HFdzKFjP3GLNSZUJUqIK5A74o6SOFGVoN6xACTspV2iTRUnuzNoCgH9XQSjyrGf9
f0TuAR/c8CH6WZIdnDdp0dfmwfDUhsmF5e6PPEf8MJMlgcw665NNYN3Fmk441WtW
88tDqEnOmh22xwtif2qcZnSHjU3rkuxjr/tqwfyeigH4TSQnFkReD/K7hz26LvM7
7qyyfzOu1Oun7KVn91sS2gDNCg+Qdvx2yt0xbCCcNUyYpwk0CI78xNvHBgzh7Ili
gXdAlV2Adsz0Kr2fmjfQIQswiTt+wfLsMTqEYko7Y3ypAc6IookxkjSoTI4vMJ4U
kVRWdbhR/eqL3CJMoND6afriNbfO47QQJYnQijj79nGphFCIvLiXiLX4kEtNchBm
VYVjRgyecnWCIEH2CweGJIhnDtRcZgwUfAMucz8JM8tH97wEm5p7Rlgm/ySa2iit
6foJwrzxjljAdcpQntbEK0LiqF7PPfgX4Ls/GvA+7SI7s9QOzVJpCbadmuGavHPN
g9d+Hb7ZnzdM0+ICYaiOXUahsA9TuSloOfktyx9wqSekQ19n03g5UItjEC94I/aB
HZ/JOKvISkhDr4Gn5+7qFQPb40ynJ/VxJCcFsa6vpjh2bvwenknqTfO7ynassPQ+
Wz1nmSGS4DwYJx2/Cw8LnYBNPwT9KaX+5BuWaFVGC11cNMZqioxpqVxV96vVrG1z
cqMPYyaZlWXCNt3cUm3ubJuayrdzXIKyUVQITic5gRlkKJkzFgj9tQ0KofFc5hgo
OA6Hq9NcoBvbtTPt/0Fc/HU+vVGwE7KcI7QmzBCJFdngS6XhhG8w9gLGe2OlUl0y
Vy3SsAVhBx5Lth9nuhkt5+hHDDOC0pMp+qxZJPBe4Bu8p+oRUcoFEGLPV3D+O3Yg
aSV5O8PnajpFzd0F+/L/vprvWzFRQ1CAP+iQkC42eIEXynteKS4DPlLx/Z92CeOj
1G85S2w4C9Y+rdNs0AtPvVoHDgU2lY5Q9bdBFAynKZvesEqHSvOWShU+MFTZMWB7
xRzzQeF5/+eH8mqW85phadrTiZt3vDuS33v/G+v1Ullr40uiWp2dY+ciI3cBYICh
zBm6GPEsX4vA996cN1BZpXdNbNwL1hzfKrO7C5rCLh6AxA7OQw45TAQmyrd4B4r8
xLJ6Gi1o88J2WHitA6qyjw==
`protect END_PROTECTED
