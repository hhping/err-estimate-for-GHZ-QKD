`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XjXSJvJ9u5ZUNejKtCgiQg4cdP5LkxuiClyEZy6pXrkPrOSSt7absVpDqa0G7Cd8
m4lfiSlOoLeQpRGb/LnZuP+0PitL26YRrSEyJNN9PDhnCA8SkZkCdiZJmEGoQfkF
0CA0pdIb/wvIWZ3QB7iBwW/aGoRdb5K4O6j9ssCB1uVMLdpbEp2WSXhcClEf9wXd
abWhi8RJS+msDgK78uxQoycLyvLsvTKTrCfAIqGdnORN78UkkklfsWgMhc4Log56
zbmDInvnko5lafjHmfQYR4AjuesGwPL+gA1PESY7kNY6jF/9hPwoXWtCM9wPlOha
t4cSHIKeOEBUtfznNt8B4oWHaU9og8oxl90tXmZHdWodKRwML3eHvzTel+GZ6eIK
k3nRJbcNUiePgdiobSzDZ2vt+Fe4+EUL2QSyOH56hsmanEt/I8EoJOdzPJ6mk+wd
qWzDDOItWzdvOHJ4ogHdhsWmGcWAKiy8Y/WrmfYGGRhgv5ntmkuuAwTsAfC6IuR8
gOrSK+aBzLwwemg139gVgO4Q84WpoywrNLmMufLzXEz9qgZqw3CUtNksLOUwzABQ
OZMZKoAE2UriAPgmZt4sz+NipbuFjQyRg/67Chl1fsLwutvuuBdSkyv5W63hmMYe
WD1cei2T2XkJmFwIMaDM9QrLeJ3w3EzyHIP7mE41BONQD9kuYt9hjCR7Af2wLSHu
ZjiCArkOL5ZEP6VMohs1CKul6K9pyQHeDbtUGnnDTJ7fS9acoeN1/VEYIomnEVT3
Uvbu3MFT5s313RbwEw+1SnHP/tHkJdMzDz2KjlSTjyY0SLseKOeVMqpLzD/UNGE2
jK0hKPWwKTTBun0dheUfBS70CfDzQ0AnwZHKvbCnQxjfehG4UvZdSN1lxCuacfuy
t6SohrQP2SJL6ULnkWds3xB0LZvHBl6rT6n5ePzeetFFTIAfqfmV/OF7riyu/jTS
HkOVGWTwgRmg8QdzRIwE+v+hTKoZ1nabNpzJlHdniIG7yY7xzNBpZ30oEwUUWXro
+FYnd9jFoWLSTU16YkOyOI412aO35HprJUNU3Yj2E9pyp70dlJx47ieVQ5JVAp29
505hFxCdjXaTFYHUoXc8y09yYpmCoVOnklgq41LN2kM=
`protect END_PROTECTED
