`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UySgePdIZgfNu7aGkvNraRf3U6x5rsVR9fVtY9CpyXARiG95gp862Sa3xheAfVcQ
ZFlD5DBEOXBo7f8y9bG4QTcz2mFOsRa49W0vrMToLW2BtALfutseOcifAX9wtSdQ
HXdN93PDSABJktMse1ACUJYtXSZX+wNKHnjl7TykcyKNZJFPveD9J44FaSHy1KlI
W0B880E/vbMUQCJzoV4OBN9E+on8gvALeyEghylAknm9M5b+FYxsf2vzIYoZE44U
a10Qj1xk6cTKbByo4pTdV3ERo7YxPoj24gcBiOoztRqJ/avoFmG4LuQglulOsTFt
VqLtFxz28i+/E9D1NfMmYm6TKn16Esyb/6iVxFAYrfzsIXzqPDAcShVfrJ7TwWMU
pFUZM40Wv5DxY8V00PwizYvUZaWwQYaO8Ccy8+9n2OyoopBJt1YsiqZutujgUR3k
YA7JMr1vreHqSRDO3k4AcDkgYs+5TueQHSUeK7YBaYaHt6tESrzuO73xso7eNWC3
K/nTXP5URXK8gb6+UxqDsO+wFexCkXSQEcI5G+/tI6hr2fjUTcfm3tojPl9deTlI
8TB3R2l5ATVmkmN+I3wewkY+0qgcFalgFh+Q6ny489XzAVK12DrUN0ow2U/p1y6d
2NE19dXIuKNFfoFpWnBVKcrQPM4FCINXH41icWL1QUJVvMQwwR60I4psue7Vxahn
u5z1jKnFFzuwby8rkZGKNhFhoBk9zwoHOIpCQSfUHKlXnIwOhlgYCyiMq3Phe1qW
UTjZZGNBzs5qXY4tafK6yCctozWQU5YtFnMB+Rh4i5O8dNz+qxTy1rawVgdjOeVZ
crJvx04pxyyhoQU8/GrB+TpSXTgwGaCM1YZtU0V0jeh5OmWfH/mHtjfz0J+bDwRo
dK/grtLv0360CBg2qSlTCXQrHrlJoejKmwDtH+x5f9VoJ2GttF5ajdLwFf//zuND
dr9lN40MYhraGxot2SQ1N3IMLES1PQrjVbMuX4tAnuvMFfn+zrMGkRj0OoopBujN
p+W04aFkvQ9X7dDlOkgPCPTI/YtxXoEeFhAQ3ohpqb2kJyi/fdbN2+CXkfq+3pET
pZg843jNYB2tnOHsf/+WdKvbRQqk+/u4GkxKsupQIKA2/NYPyUcS2OEVT408R1YB
U2+r25fEVo1ntk/HzhVlP77lD7lReDg2iWh/weOlO/RLwa3/N548yWevhrtgMptr
v60TshanZg/UYvyky1Tc6GSilzcvyJkV0p0ObWpZOL64SfY0DfVF1t6VaCYTjdxs
r7ysYwlQWj5wRPOoEoD7mkrmB2wRBv6C5BKDYNG7GjvpxVzdkdSfKV07/CpecjnE
Ce0ngTpTlCcimIGfYCoCohGHzw4PPk+0ShwxPF9ECAHgMncUYYR8LSYBRYspbOwu
RIb5jTsEOTFqweH4cYKG1OZlWiht3BQ5q7b0xzWkFbFPv3a32fHzGEWlCSf6miXU
3MZg9st/q9NCP+ezsOI3npIWvC29ixbAe/9ToqO59XiSW/3dIvSi0xRp21vwYvGE
r0N09qZS5y5fGXgH8fitmk/FEj2/b735Tz/c4CyvsfwOs1uZ24FndBAIFg6LFY4K
dshWhMIBvMXbDKxDqEVlX2cfySAaSLsdC9eJT3rRkn7TgEtCZuY8zc9rd0Qz0Bx9
Fk1ec6X3kIvXdLQGQEq6wQv6SG8YguBesGxnpMkTktyg+1+SSPfU/op1dH/WX+pD
bcOb3KZryu3F+MWgIxNZ+1917DGRxHbtCoCkzwpO5gaE2IThFJCc7cNji1l035tE
lswdmmRGmkZpKhXgFKA9k+SqXWwp6vHnkrC6sTxr9cDZo/SO4kkKvLvMhehweXDw
hQPudH2Rg6/og0ZetNYDfpVYHXnKy0Kl3AeORSBcMdtitdyqu4zmEnRh6nKHp2I8
wHUU1fLPPG0HpdLbHhNQgCaXvu5Jng4ppjqsgQWz6QHBl6Vukaay+RbRxcO8oaxV
vUxjDQjhMmiqzI6ZcTeVN0lWEHVg1TNLrNCuYNX1GsgFLI5RiLHnBVzW+ty00UlB
tkXKGn4OZ7pOx9GBa1xBHdyZj88A3I90cOXqytm3GdAvoh8HpY7LgM2cbLF6FGdQ
RtlVas+oYj6gNHLAj+6bHVXrlUDcSTJENVqk53iCd5dXcuyrug4KDjOMGSE1mzdP
KUHbwnaBe4sOzJ9sFMzWCXboBnmTfybH/Vpskw7DqAZQ8eZTE8kbJfZe0v+OsuVf
fIWzEBz9gpLieeyCn8WUxImQ0QVHkEj2fCKgqGiHSuF13f8s8M1zRUxuXNyASO73
g9NDyBPXURQH0ZH8sjrS79HmCD6EjdaeNdJixE1gScW4x4xzNEme3+pKRaBJX47u
JB4XLhesgAmYdpORSemTVY2j6n0arTI3jRVZq98+W+cmCI61JC4KxKyqu/kLaI7q
j9Tooha2pWAM0M9LCESzpe8uN4DlmuFJ9A+kaMxAsQUfIFfUYgf36vszaCbqhirt
ITD4euyEWAQIEOfRispkm6e0ukaOApna89be4F8wLY2xbH2o+gf6FiaYXjbPOKUs
x8hgaB7BdBaUud09/Og/WfSGPaRpPIGiZNY040x8acFQfoHrY10v/vMwEdtTYo05
iFMWZ9UvZPip+AWYOzgJqQcm9XbCJaone72BymPvO4MbsQDwEkz1x2WruI2smMST
oYrcMP7posAZmLwj4u6bd7muy5CNquTgUlzuZzpyXZhRXmjV43nXJV5LzBotleqd
XQNsxz768rSZ/3cBn8I4fnvIZxqMhFYA9ZhEdAkrIE4yS1oT3Hv1PFTphjMRASsz
DG6guOWrPigWtXcRNzOeQ8rj26TvuN0I7IiGwX0Ba5MFKNPptrsef+3ouagoSnL7
L/cpf6XPMdkQeRnExfc7O5gKdMM8NslCejvwg7Z+LFMe5fXfpySC6WDR2QFhaQpP
Yy9YADst2CIYSQAq9h7xXjr5VjqhUx7is0HlgBXM7LjiUCJqYMG8sg26QBkrTppM
/C54wSR7ejY2whHHQH33Y0wJqi5kxXEZoTgPIpPskjsPB6ZHqXyKnS6DKltcFj/a
40U88FdydFC01VjJuWcEghCttup7XoQgMxv7mxL5L0ijeDM1H8kh03W28TutqVAa
79I5okDv8pvhhp7sYyTZtFQDy7X+/Zp8uA2YeN2eWRztVkIXVOvArdcCyqB3qes6
xS4ixafCiLJ1AO1eq5pa+6cQIYPE79XsCzoohlmaY4SRsbfxAdSNwt4Sj++RJrul
A5GV7HmzFckPiE97zk7dS1s4FHtNt1lm2RzF8EUp6iKKd588yn2uTOvh21vZ5aa8
qz21fXACJtFWbHDrF1qNe7yddOF6phN8dUwlM7zUsYKCMUcmPVYsMfOhkYX7m/V4
Pqbnx5hPyl2/19YdROQ2jcXJRa4mwdPDYp+h4rhsF+2xlk1KG8WxYuNTAwfFEtzx
M+smOxoQmKgBCi6m+mFwBgITTyQnLKu/In+xbrKrL7Ybfd1linzb2AE4T02vocWo
LTt1PV1O+0vtOPR4xj8TZY0UYm3EVXfz//+72hapwDE/nZEdSYvkqAgEYf+q1C2D
yh91GCnlerB/DXhyk5c7vO+pMBMpeddBrCZBpIPsVgue00vSxTpmMUfq2LdB8ux/
1B7LDL9S05t55kNMEz+nwjZKNbSPzKGsh0XGxepexrNXxVSvkuH+l0Gykcaspnty
H1+41d8/yqzWx6+CG7WiSl0hidE+ePgoYJI0/2YuW2RsGwg2riMyl1U+sK8DQIfD
4/Y2+QpLISahxrpJQD4PfkUP+ap1tpBY6slpIusKKDNMqbv3TfEkmEka9BfR/0IL
SOdsRiQCVkESmTOhB98EeVkAOv13wVdSlN7dQfjY2T2iPeevem1NUUPz5KgVCI6/
WcplPJbV1chwayaWz+sw+xkM78SVF8RxR59FHmtVU9wM/lHxzQ5t4u6qd3Ins176
RbEO7L7NtmagwZiOrNRclLgOR4ZZvHdFXNRwzAn2fskvcd0ZI58tbBrWKitZZSkO
77uxjLNuq+NF4CAjFPEtB92OeDooi5J5ssR1TcywLW37O/VQcUNi5Fspdz02FkHY
ywyu57NSNF5b4Ia+skX6hG8cEE8DzIGfXaOwu4IkV8TZssr7W4McY40u4P/qoSG+
c6XE+0DRzI/e3CBrLUg9CSdWfG2nAUm7j1HQ2IIQCE76fbAVAr8hTYugVz0gT8V5
SxJhTdhTOcXQE5jsfFTMs48XXUrVt7kwBLcG0c2qvU4SFyHDElbkHKqUqQcU5Y54
VY4N6qO+TfkNM1y3nGOQS9hb0qDDbAteNL+RoPEViZxBpjdS98vo8bkHoVLKEgMc
5NGYGpnosV1WQggSPGa7ximbBwc3lC6zp1Ih3IEB7KJ5WF1ILL4O0IDRhKdV4fTM
A/wcdyh0xNBSg3dk9iIPGH5pK5GaGBLLzCyZjuCT5rcs9Hm2PzyhS2GL4nhnEppU
ZPQdS+fdIVoAPivUtVS46Jt5slV2IiDGG88aLbZvWoWlwAjM4B4vu/+M7vVc88sn
38ObUR4NY5I0NI9CQaCm+g3W6vnkjQKXX6CAwUNhzqSY0+LaPoC83UpBq/G+wj/M
ubI44wyTsMJ2eLEPFIeb9bQLGb4b4gQyWEbTM+b+2O67F+GZvOMwcufGdsytXAou
kg8GyCsNj2zijus1fhijJDTC7kXRLhj3JLrt8DuExLvS93cHhXrd6yCCt1X+UF3I
MLPhudIkSossncPFQlmhvUNyQnYoeitnsVYOkkE5OBBZpi5ZauHg0LcUtRANAqSW
utYATgW24wu1RZ+Fg2mDGnO/2WdJjKgco9i83tmZQz0DARinhrXLhbwYcuEmiNsr
Bjpq6oVtjO3FnC59Pb2EOGVfRp7KvkhnAceEytqGMnAXkpnN3mtdpgk595UksZCK
s2/EEhseEOC4+ncezpE63ov7i7eAq2Qnns9fM7GEjWHoPv3AMwkkrdwaBRs7o6L7
P+ogukCFVk0NSBO3Q7ZhRsE8bLUUC15dtUkEn2gM6nSiF3yfA53mUnhDhMFK4DRF
y6/oIZ9F96odCesDrUTgH3A8txBAZpk3hAyzn+OwYwIgYyYavBoY9uf0yu55YBBG
tU3YvC1An9S/u1jhqnEREJodmxiUYY4ChWAPkZajp2UG8GZH2LT9pQ+El/Ms9yXk
5mVrEyHjDg0GOSItMkf6BSbMZj6Xd1MhsgiH4Ku9YQQF5tUVXNfRvlYKhtg8Stju
pLDwgxHl3BoXtr325qJeu8b/qCm8ppdBrq8VS+DtVY1Ke+uvO1L6VnTKll56f+/W
IuFu7GjNCUuvoz3oPkHA0S2uweNGheqjNiqVo6KzTGLho4llgq/8VJDq50kfvlqK
e12cCcaaYVkRFyBqjVf3dHXOrYoAUQGNdm8X1b3/jtpbJkUKG6olaBAt707GfxnW
5wTf7TPwPXW3eoivRqH7gAPy+jGN3qken8Igg8Z7MzGeb6c9VpDeKfOJ+tJc+dPI
n7jt5TZVYN2WZZGfbkEZhnU4U65619zne+NS5IHY49F8+SitCm4JcxD/7GncbWu8
WdTAKfbBJpAAaEEK6xH07zfj7V/opogB86XXXMQ9c2c97nC/zBmK1PAlkvHSrQIL
ASvaUvUzoqSe+hVY7hDAX0Y4ZKecubgYXXhVuT/gn5ewJqN9qFEKt7DWuBM6bq1u
U4tnNRIK4IS3c/3FF8h1KA2Hw4Vwx3ILUQEWZTvsVR5CLfiFaDRShGkFcMR8HrwK
3w0hRkNFDe8lsNxexAMoZXPOdy4lFJKb0JSywxjyoGHWUeEEU+pla5qqopuu37eW
B7VSQWVFUcTKcKXcUKdjs6Z0aarAuITAqZFyUqNTB6yGQVfyu2ZD+ExagFDfyMN/
iTfqAzyUThwhe32G+wKnnltQAheX5bE2KjxywleDTov+O9CU0NLVM9l15KuVuTgi
w2lA4zUQhLXpodKLYh6MdXXcuDHHxO9xjzjcSlM+Fa/B7JkIu4DpoHZYlY9uVqGo
pwzMQmizBKFGxHjpP7Nn0OYczoaokeQEX1TTbhqY8etfLzhLlir7waO06iZWfpUA
U9CHJEcagV0QZzWbv1j2LpMZpXtNXUidgoQxPGgyX/twfCkZD+0/nmP79UrOQN9X
YLHXvLoXZC34YJNRB/lwDvN4KOcnGmEFPnpZgBRbUPzBgQXyMmGrw5/mJa+lQ7y7
PjeEL8FG1xFNHhlvgEHlyH1qa6uuRK/taDO/qQ34qk61/75JqXSDwYO/fDHY1FPh
GK9dygTL4Y0neLoJbldLAh5au61b5Sbu9fdjf9hBLRaqjqy/AIreo47GZ2/kREzU
pnmY0pNEsvG24n8eZiRuh1ff2q1opgg836isd+xTXW6Rwr+xzkKFvRtfZ6NLRCqR
Rbo1l7jKUX/sQwsUpTUk3C9P6qsQoinpAM+YSDhetSA4253ML7OGJZcp90NzKbJZ
ptjhXhvRZuE/bJk3xz121iENISD95lcWih+dyPrnhGPRJUA74D57kZOdqhQUip3I
f5bSIOMVOgpKzgX4RWdfuO9Hu7iHlT52ws+9+aDkakrgd8A1Rgto9ldmglVGEa8z
bOYnNc0L5QgegJ1PEDruHajBrRETEMFgDQywZ4dBhqP9/wlrNf6RB3iQzZR02YUZ
x6DpPLbEOB1t4wt+Ss5ohyadOdH9zeMKzQFoGjkdLVB0CdPaI7H9nny+GkkD/Zjc
kvco79sjFx5VSj/xRgqHy/hP7O9vQ4HKVQOMbJR9qNSW92rcNlRlTf99DpRwaIJg
DoNGL2VQ3dIzEo4t62kt2zO7C+ezA54ttd8Rs1+B5xwMB1xGZezpqtvB3usMqPIK
fRUQ9ZtU/PYQdqnB7yNdxCv9HrP8eB8ZWtcoJBYRcGoX5ZCKsbq60E1NnZzecSJE
/ARifFnr1lb1vvdK5JD9FZq80+k2gIfHJuY7/45pN0zSfDpYj8bXESX0EiNmObSH
LnLrJXgCB7c/hPDwNHvBzhtyquDoQTNzazWvosnrDwKK2f6H0JAtQTyE7iC1THrP
Bx5l62+aMpicjCrTuQR70PBSb5EJnRp8cyx0bH0I1LIP34Z34QPjJNSRzghCsUej
ni6BVATxCUXslPZlbZ90kT1mM9OKO1PfdrBSW446mcStJaBgTOZSCBHcFVtwwjzS
hFIJkP5IJNxPN/TVbC4lx2WjMemJ5JF4uqPxzB2ePXMSh6GaY86NXl8BJKH0k26e
hOnVt9CBMETNoIZZA0hDEXBzEi8ucBMY/eo80l//95FELaZ+BVR8pLBZyUd0jt9v
QpFEiT5nNy2ZhwasTXcg1C42WbHpzpC2VptmI8PJBmsUOBihTqYPuS3x9qxVfN0c
KX1w2PwNEa8SRJFtIJX4avLCbKW8+djwiFiG4MY/YkvIVuVLByD7sRzI4DjiTeKR
aeGw8mfX4Bm/mmp0TdzJ9c5U+631DhSqQr2Rs2r2bxYPWBsi6wpg0o3Uty2uSX3q
Sek0HRSasEGuGBtsI5Q+BZhW2M3PFki7X1763pNmO5TbSgIGw5CASqHUM7TYvgx5
EPagUYgvBKVMrtJs/4ELTGDLeV4BJQwLteiGdJ1w2HwamEJwnZhg8gb0K/isarPm
RQYZukTLY5e3UCplanAbAq8HtWTq4vZm69psM7rGwhyzPzAYovOm7KnETUv1eWtY
nB8eHsAmJMpIQRcbNhNtICMpQ55BG8LtKE1TRALE2kHBgBKgKu+WaHbcUSuYFBTP
al1Peh2WO9igenvTyxWGLgsuEsrCTaS82bbE/lVVT6CuU76Q4RxkXpQxGNBJ+np6
sQ8qomsRC4TUkKLDEJNy/mllVNJPNtydpulTSzGGzaqMuQ3zdNybaesS9usKz5FE
qYfht/BnG0V/SMWpZnNu+jRvgT/1CjtrmON6ozLETe9crPYwOImAoFsy3T3tAlIi
c5x6vLBNi7zHrBY+qRAYq1wckczco4dn3XMGVDt3YsrYWcIwk+guDlKGlXGnrILU
9N+klFaLYEN29Vb0N0/xnohSmqR/oXgNUJEORLhpJH+yLlNuzBc2bVqcSDD6LI6P
cRq/D/gKV1aSgWijz8WZU3ZmEyfeug1jkl9cv2qDgtinqi/m/hNEqd93gcHcZelJ
+t9wsvZ9fNAGsFftH98tbs5M8PH+oCQaiAkZ4ZRo5gU=
`protect END_PROTECTED
