`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewKXY4nW+BtP0dpRsGJmjrD99t8x++YdIkUgzN7zRa8W6mtmohGV3/GHjjMCRnI5
yj7qBTLQNwZ2+I08T4GECrkz3/FR76KStgmCwzTTOn0SEVqsZ/hMpE6acOw/qe/I
ggBK7ffO2bM/CMCuxibblZj1J/Rg/MmP6srNQmt0pXE3LgtCSFofubbujOUrWZTG
YAFpg4on3FZMhqr7iG/SwW5nooPQ/Q8wAcqlJDh9nDMlBtJ45MLHlcpRpMyDbCj8
ovA6qulPce43GrQCw1z9+ZbDBe7zC1ZdF2t8yIurVKAd+tj9wI+5Fyx8UaGEcytP
2VQk7X1SSQ8ghA4KrgqdNMn3qX+jpmQ5bq6ZtgoO74wp4JW9BEXUcMKZqqf2fLOf
B05+MjUcphijZbwFZAJnRrnI7hALKo4LSR8d4gamvKfNcf8jstN3Zs94Pm1pM8HT
i0myjCHhkT05llegBjd3zeBXuGo2mzD8yDAsgRRoh8oCabas9oUfcdfnUyLhP2/p
/4xwLitAz3kuSvKCGTTQmNswQCcn5QcmH6DT2e4ChrVKiRTheeoe3eM/gdVBX+Bf
j4C5gSBeO5GSVhmuwB3+2tg/+mY0nETHPOlZIPL6R5/WyF45GedIsopqLRgxOENh
dz17zYp6JQyFZtGIDq5Eq3Zz9Ks24fWku9CptM6x4nNWa3CQjQHL3pgAkvefAp3R
Oa/r4zvpeNoxDKsEcEGxWTLaD5GINJweJl6WNvNITZBZM35fspOxiqy/k7HwLkD3
nCCK/OSAVHj1DBIDn6l3bmVzPm6DxF6F44g2sGdyMcLBhyKgYQz2I1oyrjadZ8ft
7+u5h5+SwxPLof1NFyHyLCzMM6erTBdFqMBoZMIt5IiXzHSZgS9rOGz2nnP/PmdT
bxiqh5vbZrTNVnUayIbtbx16FdAHXVNsmWy5cDG7hfW6v6rjFtnOMQ9brd33Fidn
8ix+9F5Zeqxpl2TuUMafVkbpGBxtoOgf5XuAM5LmT4gyedrejP7O7gQKiXsBYFWH
ueGCo5a0s/6nETTKOeErxyPZ8q9IgRdOic37xuoPFb+vLeJwc4SRx1xsZN5Kmj+J
tdeLqfK3wQKaOPeP4pSsA+ppm4leu79wesncyFlKdTZBZid3MGfpR8qInNs3KeKi
UO6WXjsEPJybVH4rHdz1YZnOdMV78Js8S85mZzUBgyxrbIQn0hxV6btVhcD6ndW4
5C47DGFFPf5FbgV5eENzRWi5q50+D2AJhZ0MX2s2h4gl4bmNcIDKIlZwURiZLM2t
qCtowF6ZZXGCxnLtuUFVn9BwJWrZP5MtpO69SttdgOgZvnHqiif4BTrsTKUyEOQX
3rgBoNmMFnJiwSZ2rw39kaO19yVFsggOr0PfUgEJ0dTS24y98jVY2fB5PAZSKST5
gGjImqZjXBTQxK1ESMSX03J7bjtTY9GY3XLa1+Elm6AnpAl3zoJhYeOQ7pj0kgUp
ZXcXn8ibP2z5VPaqxcMfJFtmvU07KNX70A4F+7RBnlVh3IxQ9BFj6KtJy9v8oxKZ
1m9YnNOIAtepXqsi9Pf0F44RTs2oHrGwduiHC9gCjWff16ic15gl+BM2k23TauJf
bkoUml7pFO0YjQEJZPXbHHZ8s+IMUL5auj9mkE2BX/4dQUX/GXHz8SB4RJ1My/TX
8/nCFh8ZZBUpPACawX9pm4zrI9n89+SX+JkscHJP/5Df/GwJUOlRKhfVGToR3w/c
LLxHA0cxabIHR7I2JVjVEDnjBnI82Jkx1BWyoCkTCpoMHZYQ+99qzzI/oa55Eabu
2OA5EiTIHukR6PL0leH7W039l8VeIbhgnOw5sgCvNj3Sj2BGJCEqaIc3SNOYwT1R
5WC8IIS5k0tlm6guEKSDug7FV9lB6rmXFW6cWXla+ijZS9f56OF//mF0AWPcbQ3W
FZhgAMOQZMjDimsc+XNL8u8mvpHTj36GXSB4WLgCF55/dDXZUoEqcWF0jq3FyEa0
wfKhrFHnVr2InB19xWCxjCveQWXFBAwz6QHS+Gcc2hPg1ZVnBs52WtCahItKzRlZ
VcYTSlA04uQywgo683/fWGrk0/RV8FXzEqjcolx/rOhHiJOdUS9LxS/AyYfGpJYg
JLW4KcawlCMrH7lMJpL1Vl0HKcAOen635PHzbrApYIBWn+J34SBEze2+eXHNm5d3
3ySPR2bYQGYppcDu75iuBg1ncGCsE60waThf+nM588rR9BRgMLce8NcAWZLV3wqM
0QKJxaoAX8sonq3OK/+bcC4HQjHtZKJKpNY9F383gXCejvoqa1AxgVt5/T+2oHVj
eDzD9l9G7SfPW4ynvMemKYbl/Xq9zYx3P+f2+yF942A434B/JJTrgOtIu7Zq9Z5g
3wEw5L2ouGVqfEBSsJVg1jZe0vzR3HbEqcWmWAokpDBsx5zLt2GlZVWo/b+6JxzL
JKk9L7bnQsdgLOt/iTwwefkZXea7iTxbFV3s1wjCduiI5xzHUjd3bNlJtFuXxfhq
GiWgIu10vkXp8SffVvMyjTTGxZPd1qqICeQqZnCHJnhwxRCUoE0wUto4bk8r0pew
/7Z26MpZwk0VDfoUzq4Dz4VF71uZ1kKTp0ul0Tbw6AFJj59Kxe52QWWdLHKkq9fs
3V14/F/kPvURMhdyb/yadRC66nCNKgt+BlC6r35uGFRqWyHk6Cx/R5xae8wSlquV
r4ZvFV2ucqwW2i4Qizpv9OggRNe4RTy2vjImu6h3smrcJ7hq5WBuea5EMKeHP+NW
o8HNaQtkW+WrgbUSPkGnrr6K7hU9cp+yNbh27p3P3q4GhfJPZeL7mFksSaFOxicw
712MjvN7pDsdvwDjxMDwnUxdcEaiWRZSmPDLaNfO7z0jLInuqaUs9DNwgFB+qurr
GFQ31nA1nC5Ew3RPdlnAwPcPkt/ABZimrGxBzBCTMI67I5ndrnvK6kMOE69iMLXF
5JsHsaM7V59+/2IlQjFR7GShj8R9msr0gzYcrn8iUUr5QLCRlWusUVWGGSRxWkWS
ynfASuAInykTA6c27Lkkk3C9MxSNdGLnPPmN+xipi+zBA1K1Sv1C4DdMkiZcgpLQ
OwKUHl9r8ktiWby6k7gdRO7CBXZUVDzulZIyAYdwxEkn43NH9mxy767AxAAyOuCK
BITlJDVZjAQgs37EROgetTOL3cseTBi7NUHKub34W1KNMXMRjHKbWj0ZEGvIMn+J
Y1r0WHaKJpNZNp3IyhuM4GgVkRVgQ67JS2l44wMwbtAIcAhnD8ipcc13fn4tuEVd
GF6B5PCuMdXQVcHMkrsaSxuIgpRik5CRGkKCA7MLNV0YNHpjc/oGnImmtEh5DzzM
OIeM/CODx+doRctJWlYj4wEI2hFFrsJdWKQTBuaERYdw1OmJW2lzRB7P/+tyHcm6
6LjBAPI9fAq4GXo30U42mzh8cdnpgA1SOk6g/C7OdGxCiNBKUtz+UqKnIsPQFIlj
C3XW6AnShMxWBWx33aRkVRMyMMNq5AYp8Y3sNvtSg5XDKCMSK/k3xYp+3uAlCrsv
fy3cyngImYTyzfFNUOgYEs738qqBNhjJDeHl4QWmbUhih33/hEwL45sKwo5KCnZI
Ylad2/OL0F23mM8CK75pmzRQ2cC8wfEzTH2HLRqmE427PXolLg7wXJ6kYLReWjG+
YEtpEHJfPcQP+qG4gOEejiuC8y1kRK7jS8E+YQrk4eopyP5JMKB2oBUqHlvq2kAE
Ckuahhb7gT69tZjJHCSpVIu4lI7YH8tpce2zkhkR3DlshLmHCphHKe2ebpclP4PE
ZOf1AzI/GUUVspPDAs080ZeCwY49Chuicd33KtkTRpfimqDeEFTeD2YzCVcKNYKW
VpcaIQ42HS/nyhfFkFuh78oqQ69T4VTT+dUsvXs1Ewx8KdkwwI1yWG088+HQMENT
qRIfL6PtkMHK8io6lQJft1RBtxXpr/VswQA7sBsw59SLAdS2yTFHMnjsLsdX2JEZ
qMwdB2rBxD1penTlnaQQEwrnEB83Xk6wuIiY1EF12eQEit5RMSFmbHNbZrQfLOVg
ki+9E0aStAkEw6YPNlGOow+LNObaM2NcphBbHVLJTyMN+u6XpEfYqrVV6XI3Tyzw
b/csmqz6XrPs1EcLjWAIs1kR2MmlTrr0L5O0cFCtBZYOxrCF3/preAB94n4qfpj8
BO2ljDYyQ3HONbuwLUMawbzTjUsARrjE/bFwci7XoO2qNCT0zZKSdvOk8/HiN8X8
iG/zKziCtdGEiec/uwdN8IxbKv39pKbJx6MA0Bgu0Z8KeCHHC7peXuHQpop4hdsu
jnJDI88y11ma3gHop4GKS87Ju4GZoUChsg6QslfXl0WD7KF23ITBUt0HCMtod5df
PMo/P118xweNlC/hvkMLnEbrA0no+Jgy3nufVhlzx226tkwyku8OnwlLSUj3Dka9
coFVuxnZnkQGkFmN1xc9++4e7d2gPJ0CKZKXUkeP39GQaG9wrR4DFbQNhxPR1sQN
6FAKx1pTxdMyC7sghLJ5HkQSlUK256mNaJvm+UPdtsKuO1SCYUffwj4Amq1bWnQY
srMbDuDj36FsCrErHiLczcC1/WGr3mlXBkMPQpKe1WdFKGyANMiKsr++gpcg4jPB
9ubtFHtLvo3ZI3t5BN2rd2wJZH11HMbwGu4YLrjQAdz5iA6MjxFRprYtMVoriow8
iTl2TCpkvcloV2RMIjLH01d5VK0qe+mC13cT9E1tgm7bctwbZ7sOAr24+SYRAzUM
QDLdYjNYiiZB6ByGrNtaKrvFpAvSqu72PJKvPsHYzKh5FJQvaRD2T9Ql35UPDvsN
WnGrs84xCn4hgWIwsFQ6IfA2d+oRqpUQPWuf3fmuVo2NP2MQHOvUAuWPTfc/OmyP
8Xt4rJeIXLHOLZtPHqqVAAH9Zg32dI2BZkI6PrDYeh5r4wRQeIDr3dWcDTFZVaXJ
bGP8Q/cy6EJRBB8EELq01ElHLWBZTK72vfmZUWo/Hr6bGOTU1U8bKCRc27Ah3pzs
Cfn6rXQMxpDobUyTP1KseSXLcPkdLQFU2Sih92n1HqONa69YfM/0kymUCz9dP1Y8
canuprdMpxIsaj1DfG7MKc+/rL/YZqADLeIJ2GbexFeDdIxI4u3jfn1hvaBfWyjI
TG95qjMGLciohSNrfpJDMN68PTnKkFl6zFil8CTCQ5ofP7F1JRUQcg7BOg9ft7Ab
dixXiMxTRbPF1X1sf8fFp2pPmL0o+sbXOMadpGHsIBf6YfuscQQgc9oBkQ847zpg
RKoqevZAyedfPvGHsg3xMDGZPsBWTaFpgEp6dw1eaVsmzqHkHoSUi/DggxYZ6qwZ
8t3iI5MOpdcZ3zBu0gvhkVaC2Jkf/fIVbULDn/la9SWPuzxyHqrxGgZ5HtISlHrF
lm3sBQ2oGKzlmSS52Nld3CJ61KwckA0G3siuTJgrhJ/H8YiGRyrndWItm7fNV9Qb
YubvF6uy5DqLXCJRFkxEhLiAR76NzcaaCb9aJDpHqorw2M22GmUI89zP8Tk2RymG
76afU8wBIDTQgZ90gal45PIMH44IT7wh4ALy0CFEbpY7MUxVVcVTgDRkDLxJLN7b
psNgrV3n+vPX1bzfHlgdI6ZM4kKaEHVIi3V8uRW4PNGJNLduOerOZ2IfS/YYWE8R
`protect END_PROTECTED
