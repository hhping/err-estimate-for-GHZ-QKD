`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJQV+Q1CbzxY8No0TpGzCyjcODiO3o4hyp3+S/ZzvtLwV/qyXkxMFLslyLdA0+TO
1D9vvHdoVaQu8vn/kOqf0l5ig+NVm1vE5GLrnterdOtEVdkAYqoSlqY2xjwD7buu
2aK2Sw3w2Vzk8Qi7tjA30TkXK8JvHQmr2qzRGoQ16KOA9Z0e9r6TjXW7QOmzTtCt
JyNMEOy4ZhjevwGI74t7NB+VESG6sLY3jpjgP2/pDEf2JaikRO5lforsmwFZVt+G
LcLHUtXgYCgw2ZIfnoM3p3kopnOy1FdN4OzGDr4gfpajMGxpQzju4N48CwdM/Hzz
oOYbp4i71hN9A7Pd2BuPaPOKoEOhklm2aoQ1vCONMgtxKhS3ADXNwodWrCO+73WF
OXDqmxnEUYljIZ4rib5vcWCKfz0OUwC0s5uwkGciauf5aqV7xIBD3yXpwTlffwI9
mPPOvECuw3V4ua+xKp71jBoJUbkvPvZkMYkTJkhi1puAyatS/D15eSyCGhxRLw/J
Sr4VgUZGeu9cXK6JXOkSCvhO/zO1P5wbEjlNDI1+B48Vj1VmTgmP8i3D0sho0XwC
/BQUi+b38ZCNJ8NCtc/N6XNE9EPHw1acV+wmN501LnWsCAV009o3EMDZKHq2jp4N
YyES9AyY87+UdvPpaLqLX0nVi9VaDYDhAbzGCgF/T1kqYew692iEaFtKEZrOJizI
GDI5e1jucU8TMzAo6m5hYN5FPiXACbN7T8VfWGFaiMqLfHRJjzYmfmlMiTO0g/lT
OcKiv6+G8iK0t+F13kGpjsp209c2vK/U4Vbt+l3xBO1SjxBU1z6Bs8o40WiKHjJ6
wpI5H9xabRKlS8dK6HHaMCpCCis0R7gHyVkbNKlVxLGSocLtDBrdAlib8QVa9+IO
xxaiNH2MFtxqmbVjZkvsmItCypyaxpqbBkoQAkWwzdUePD5KUYspBZz4xS3wwQPr
EHhofhy56ZYsg1eIYPaS5dxLdbyJAZEQ1rRG/zjJhIXg5E3n+2gcYWgh7D8CXKto
PYl/23hq5ppEizRfkGwWFgoPS+4BKp6pu6aP41R3HlQb7hHN22hPOg3vEjzC8wGC
HxEhZKwpjbbIl0IQiEZ6XxqTwSR7hzUAXJrDoro4pOJOsEGsiULlJHfHOGbv6LlS
`protect END_PROTECTED
