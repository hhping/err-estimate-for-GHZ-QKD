`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbHGB6NPXFWEAGTqcG6a6K9XJ0WDc+RdU8Bym6QDqrJKCsuyLfd9XP202dZcLsg1
JixyUZvED0LPAjVUPEFWJb/G1vPUCzTXoXbIO3En1lm5yvOl1IwjTqGs4tqWl8ph
JJGfjhhVOSZsAMY45AvL/IDLvaRmlUkaW2M4EdLkrID31kiZ2iA8eH9SYJ+89N87
LFMn+3mmq/SGhyV5JHjwq/wojjRcn62LDB7euktOT6myr31znYSyHxFJvsJ/upAY
GriJMh3BxP4OnjgBIYufm3NzaYe8SIfgrL5Air50DM/ggcaHUUjWmWHgtjC/J1Go
tf5cGzrcd9wJFzVEuio3s4MNGPQceCXZ5HwlxXs6gWkc/r8QNr4bDnzrkgfwxB0x
5nJiBFuvHJDTa2uxef9aetK6Ybbv9D10kGWFlZunHbZLLRzyXO5bq/HW/gpgDpRo
6f3hxHBmhbeH/o69TtWmuPbsICLq9Po0juMicA+eNROU/LEf7JxENNxNemffT0ns
Ov3zHVf+jqMX1I2teMEcZ0IHkIpLidGKAiiMPh5hMFSO3cVZamoBgyULvC8qNhpI
tOn/nerGjDKFJWzKjdkLLS0OoeufVdpDfUKTumgYBtqeIZHSt090HnuWoLxHhyWq
bGnE53tJ6dCEFEYm/cYYFi1DNxTduyFE97GBu47K8icQwYmkM4MHO+HcG3tcUc9k
mOMmqT5jN4pWe9pGsZyp3UKUb0dokwnGh+cXA3PbXUYiD0U0z0JrTueaTkJcqQE8
BwaleMIJUkPHD/MvGW9mMfUvwiKulOH5ZHTkO55yOtm2Gs4RHrZotmrtbV5m+Ivh
MlWGoj+335p13HefkMY90qF2Dh6GwlDhC8sZS8duHdmDwTf2y/goOmW8kheYg3aS
m6jIUd/SwqyNaQ19dZEuJBDl4/oxA6OzxHKlBX24T/2CYZWvpkM8awJbcVQ0TBdj
14OR/UDnGggxsJx6PhTo3LVROrXOpwXuDkfs6Nok4GhckpNJ0NPvnI7CWChawWm9
2ZW9NYao2BgN5JFL1mhtbBRX5fUIKbkIZaWSUkROVOc0F26fp0yACYUDdst39evF
d0+TV/Ox8gl5RjxCni1FODiBKOGoTM/N4cTRAIifLDmqKp6yZAtHpTTb7C1g6jcu
V+N2P3xflkYuVjD0Z8EcHQ1XcmBWOQfqRxvkHElsU6sRxg07IGIp4lbp8vQ56F3q
8AGdvWMGDYTnjeB9ntgjhcIHwb2EO+cMb2MjZIK9nBDONKLraTQb0UaUgr12M0bj
wFHyNIOEDLsyoUj3dsdDVaIJZTANwMzZ+sNvMlXlpOnpbmzB2/EDJ6uD8a0+1NGq
7lXRWgu2HfmdVSOBg1Tfcu6xjlLukx75d+S7CdrSGvNUOQRnw864vbPmr+q5wrxS
wetN+XTA2qGuqsjfJQ+uGkPP1pPhzGW4UEaVZq1r6sDUkMqSGCREUfOiosbnecY6
JLUEPI7jTdYjgwG6F/URIszNYC75HJmWQmPCHohIsLmdHTHBZAwABMq7nGAlocEL
oQqtpmN5UvHUTb3jaIljjNGOVOROkovf257txlWpwhSPoTClgIE7uqzRsjwpyHYX
N79e4i6KwrmNDrEI2lZ+UtEs2dYQLEFFsTpl9HcZPQRGSQouzvdek28S/7nuX+sp
TPCS19q4jkTH2KV+TUW6sxz9qLA4Wp+gBDZ2wm768X32EWGn+MU5EaL9hFGBfVT8
sKoDpcGwHTKAhrdM0p94D7mL6oP5qyomGvRvgn1iV/mHUOlOC8LG3KV3vDywLSXs
ArqOX3q/VyGZZmN94J9SUC+qZjmtfK0Sn1KgS919aVY8Va7+l24w+nBRcs+BuXFN
DTFNH9baZjtllNgeUMe6XcpRDoFhkzYaaVL5LJatNNON01qZ0bDhyS1dpEP9XcZC
LHXxeuuLlWi1ZaUAuO/aJgEOdalwdn5OpXxrA4hvtc1h1cyfw0HeEHnT9fLXKkPd
FuzPGA7Iq8fYQAGUZ7JUFgeVS0GRQeUrfqtc2Oq8/O4Xt+ci06RilgUktNm4dNu1
JRK2qU3T9yDF+YXZY92T0mF1A85IJvFv0GvZnp2PUpE1khKn9Gs36eavbwLZebTU
s4s1/RnA/AVL3RlEooFk6/f9W+LYshhkJrXf7vbLCXEqJgR5L0nAlju95ZPlqCTU
OwwtHYRHE5tk/FV2DDmXezSd/+i+hTO+8jQ2EIY0znuvPcjFg3GjBoQCDIL2H4dk
75hgOFyCWpcIdkQg6Yjtviuq/k9vwm56DyYZGwyS8r+P8ktcJS/+y+66yNjxHumr
DECD2zr35YzZqcKL1ib3PhgQ7TSgZ+0YhIyUEpsHGr2FnpIKp+09maxfp1+PBDeR
g4v6Iqj2UHQTve7xgSgv3HEGkGAb0OhZcNHdtVGwmYCmNfvESwhUMitNAoBJ/Pc6
8ieRYBgEI6B9opLnnKW3KB+LNMrOiOpBcDWmLOzoyjSMgYF9GKuEi1NtASKQSeL/
Nkrx8t+dQgUGH18h8uWWJzqJ/PBsVSPtrcLEGYRcfXLIRyxmlw16+oxUEEQVMFxR
VoEDBrj6+oIy8p5x4GWy/zDC74lZ4GTI64ET8l9QfDRDSQZiO2CE3b0gjJA6oWOq
R4sNgdj++CqWMHtQK6Psfn4cD7BBpZ33gsduona89dJboFGnMAlJwAoffkNT696p
FFQAjWqCEmVAyxQR1Z+aeFxyD6ppIqzcwQlgNy85eetOHDFmwrRZ8G7T9ccSSegy
XBxXYRUoGX/4rKqRqACLinSJbKEdRXE2Lfxf2kdNPDifsIhm1f+8HmRfh4n1vwM1
UlBVM6fS96zo0GhOPsLmJ5/MRagPg6SiHqX2qKCl38rDaRlyIohX6KhzwaR3Q6/E
CCV0a3rTKN3SE704zMD/Z7KBVkLS7UyMFEyopYgteTzhI4oxJS0goCtPOWeJE0sI
DC18C1N9r7fz3DIcLYoRHbQoQ02rk1xt9c5FIBL/3KfysLpHJ2w1tAiY6NK4Q2Dv
vOW1svKEVIX3KnYMz9cHsJj+ynd6VSRhpX5BeTkc6xust22WxWK3NId4FX+6tupD
D/1XIgW6FbWWcogv5c0Hv5qrumVOaL1Me2QFGfGAyiA498Cb1NfbY2esCIF2Vcy8
SKK5jzA6b05seAY4VbSECj8tdaqHbgmA3FiGJqtvAZqMbr4eU/0G5jFJ6pzA8o2I
PEF2rGDSZqdJp2LGgABYVSanG2dt7DlTZwwtntVRJgWdEfUgOR+g2BDMLd4VxysG
3nsalO0wn6+Tu2aoPHN1QugSmIy6Rwn1l9OotwOOIwDJnzR2ajBAdaCnr5K0UEMz
fG4XCo1j+F76mCUlJ9R2Efr15YyX9FWMQjzNQWjhh1sOJ5aNFpqHeX3WS3MEx75J
3dxbhfv7ZbfoETXbOCHSSjb1JuZhZiekcDqUE+7iOI8iavJUdxALgYlIPhhhHZpE
GWHGZXZoyztbOYLOMaGqBDmmPsi79KveiA0o3BLz4pgAtx8wD7T9wBI6nM0pj79E
8mVZriPxlexjqLQg0l5icKi6aUI3LQbMqD5tAPM42ujUcUDBlGYYgA6wloIeo78R
T2k+bOzmYGRMjhAkFcBdrO4az5b0OXEF/N/CFRgDDKA6VKKd1qcImvBnC+WxSj5V
ZldeEqfIRqsToPs0y8HAwG2TaSxnkA//SOzRNzK2nE4I2a3a777ioK1ZCMtmdCAN
tjhHwJ4BZJyez33nNfSe+MPFcVXoINfIfExRAiwi8Pst+qPJop0flbSIQzt5IBat
YcvVs2+WEHhik+DfFdyONwgUXScJHc6qo2/BtkocxqKoLyg623XbLl6NydTjCXP4
5XAD7W4QZ5KNTZEwrU0m/P2SPvnjk3Vf66Gbguchf/TukTxQXbq+N5Sm4GzR7cbV
TikTjE7qVSjB+yVB26snSo5JbmVFfnnbXuVdFq8Xt3ETrrZ/LeEiTqbTJNo85lwE
IRaCNpy0VCHnnNAWBrwzueQ5u5Jmtvu70AamYZhScTvyw4RXIjHLS51fgLIa05+X
NfHsPQtXvzek/TPqqmnvI7ULr3maSUtabhpo4z/zYAp2x794Bfpg5lPfUCFncMNT
PK3ixUkAeNq9EjJCMWdGTZaMzZQSeR5P1foUhyo1Q/t+luGovjbFrOK6948CQ/V0
/fm6M05gJuA6f/X+qSnwOmAeYvztZBgLJNRxY9fTKaualNeLvqdG86m/iRWUfiQ9
003IxlfFHVlKHpgVs2cO72XvL/I3VwJEb6b2FrVd39+SUcL3Vs/2ELmukU6FUDCS
+25MvGm1VZ1zObOr7pTwWmmSrTHtcbeYhhq/n1do2JFNA5IcJhqwMoCfr62CkiUx
wa7CMT+wB1VwiWru5EB7QJie661Rx10o8ac1Y2BUfKH1Pow7lhUjHFLY9zBuRbf0
WtmhfUItLmXZmZFVHUR2qKEUqtCnFZtp227g+CEQqdl3YspHxvhKO6oGHh3hGDKh
`protect END_PROTECTED
