`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgpYxuIaz2V8pwJNXKIXV+U3+U2k313Ls6yxCMuyAmqZAV4Sx09IfGMa/g/kin8j
fE+ch9i0s4xmxcoQd/dIY1sipngEgeb/080qiwkESA6WE3qaAL6Er9NpJ32SHUgE
nNXitON7z8GBKf4BHS2qllc/J1ordHvwiKT3TjIKQ31+8ShKzhYWCuY7B1Wc8wnl
eWY2PeWHN3diadpsoPtkPOiXf6qFWKLx0esxia7g2sJ0hZjPDGJ8aVlx0eD/EK3k
A/OljYManutmjIgoMkH+wFL1iSUTfed0QNyIVgBWC/nCfo5MjFFoitFOzdfqLPMs
GGmmDBbXtG0VwUrLEuvsCrQTqfwm6yRbHtQX8OeAxUMN5a89Yv1Ikf48YnboRp5f
aqTcwynDQ2lsXAfNozurE2afezslNJmhnF7y9UdZJNQ1/ozT5WCDVRq2KdHuCowI
x1JHaadMCcOrHyLT/8eUq42FrsBxY1IH7JihS50FcArIkXt3hwlonmo09MQzeUOD
mdfxYZatEz9RAkF8GO5hEOPWmiahj5U8m4uc3D45iuUrE7dJ4TnhfshcmVzTzZet
b3W8zsL6s9+/PmTr8y1/HT9RwhkqZa/YByqBQbYbMFAsFCMnm2P2L1kh/kGkdrgP
erV+ngiAwV0bhV5S2FLqrL4viq+tyCFYFGsochAV2UJgO6FB+chiRpZT5jNSzX7h
+Kk64d2iLZU5uNlHSCgp389Tmof8CLcLSMSXtkIEKHc06MXzqEqBKxvAc/k/bO31
IZVAt7LPnHvEpszmPhWddc9EzEpk3dYItT1BtlGyLo0NtiU69+fi6PEK4U19BBeg
UO2CTHoyktjMbxLlLmn1mqVck4u0yZRCKmd5He77EkEVUOWB0apO0NvNAkPH+f95
+9qjxH+X+yb9QfrPLJxIGCTwbYDtBImZuQFYRNhKezuHGNKWPXVJ9GBp9ckDUsD/
`protect END_PROTECTED
