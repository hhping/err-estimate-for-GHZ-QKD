`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnZw7c5OnQ+MHl3K/DIjTs70mmHnmeltXGD/9O3z/UdsadHou66ipr+a3kvNHua4
ics0WosfXYE7enXtsrImBDUR9CtHztnVe1ju/Ji0vTlPP8z47mPT/cDB7/6VJi5u
yaqhas88GQjIqsp/eG/oPrd4nUUzuI7bhTfElvU6Lq9JsDamGFLkcFg4D32P7mXJ
1PmZDY9hqs/FTstTd0JteP23FgP5lAMU7Hg21PIPkv0AGbgQI3TIraJDdybEN6wT
j2y85KxlxP6vLX8CKQpx9gxZ+hCIwMX2V3RJ5jOst8r5PyPaFlT6yXE3NuM/4qtM
yNvTFfM+Uylacp/0tQz8Y0N0Z6JIeG/du6xTUZLc/cWpjDGNOHNaZeoiAPYjORet
mY9P4nlpLqzEgcA5Ewrm11kFIaA3hsWq6BuqQHbIcBR9B1M6+5H8xXwVkcUtsgU3
8s3aZ2Y7gn3KT3dINx8LrpHiawFD8r2HXu6S1T84vujB3Fy8NOYvqUsulE/8kyd+
iMwwxcbxz1syv7yLax4gPX+EcadgOAGvxszrVzcmYLH1+4SmZndrYRdOklMmmL7G
omu1g6RMN65I1+OzJ/1LS90hInKeyznJxxxC6hhLKezEnYqm72oVTBxZyIiuermJ
oDYCAGn+5lvwZu4jxMLg3ErbAN4pE/pAjUcXvN5qlPz5XdNbCIxBjgk25Tdlw+dI
IFV3LvKuzk90dXzTnDfXbm7hbyyViCL/X4Yf1RhAvxsIRV+Zy273v2x/1SzGP/uJ
UHfmuanxC84GWbSxHoopsDcMn2ixDh4qZZKSPrMr7FOidkTYKr787W9nSgiHSbbQ
P/7f6vMrubpCyaH9cyUxbNRSmZT3zGoTUJXiB5+sLwziYhhmo871YYvg8J0XPMAH
OVJKtgrK0iSARSDy0ALdoVyQIpEC936LmPfovvEIBBZWpAbqQvqV+mGsZDa1UE50
E9cDdCmQ9rKsES17DqFXdbsrmqTVDVgGUzpGF6MdnjJydnW49wPQCyf8J+xNMWr9
szmuxn3YkOXRvAwXo/DqelMAvYBw0qivaKGWZI2lRLIhAXy7Zo+qcu8ZmaPqqiif
lDUf/uYjx7l8o4yi6/ZL6HqSSS1Aw2wzcLxuQX9qkPZwzyJjBhIXB+MLRQNJnlfz
lakq8XmcbcnnjRDgNpRMcsq2gHo5nGuwThZjbJKYrF4RRJNO0A838zDl4LHqIJ/q
hq67AFBW6ab1QFksM46Jp+78Phid44l4M87mrdpYhALalyusctTy5dvt6fyUpGIK
RaBT3JkQCW8bLit/uB9CoSLib3HvpP1ufUozvRyb9Xz/fGlJsdQ6RlPx0PmAkaSQ
i2uT3Ge1JJQI0VKo+jeeUoY76VFYuyBwInom2/ouqwp8wHTjK2kUNYsZZ/qwy/dz
DxkVLD11bn7Pt8AO4tzRc9mZFs8lAQkMTHwmYSck2jbe8LFVCpsLdV56IcA4rbNz
m0uS0C+L/lr/PI9oH5dOkABE3yDuF+GGYKam4AVy20FkqmTn9Rxk260JDVX3nRUh
kMPRhoJM8R50HwvDKVbp2ecdyKp1j5PIcgHcWQtU9/L89hoRUSTrlyMwyPsAOcHh
Sjequ3bn5aefU00QZYJSpGkuMkWzSM/4c7A88+KVg7aWAZIUi66vU1k7qdfxGmeq
gjDP4n0dkeY5lpiO0T477mrmYP9POCZp727BEROt0jgLWsLGjohrGHUujB+1rXdu
kztq5H3995tTUbruBtDoYCaZFjffJOdRA3wsTAV4ItIhZfDpVbv8dsTMHiHLpbci
NqrG0sWaIaeS5fKKv2JW+Sl9iVVMf1hoZqxeOlFyz/xH3Br32agdIDGzWmyAzUYS
G5YJbdVCD+e7e4As44zn33qxBn76PQe4SXu3Q/SGDVuLrOCWUnPJP2ojkShsEAJR
6rtgUxqeSqcAQjM1Jz8hSE9sc8fzIAQmf/UJbbIROZz/7WZGP+/3bAXC1H9KPrMv
5617XWyK2KOV3WBwx60+uBUEjW+v3tW9tjf9UiBIkgqsYLnbkyrxl3U164ChqNAl
BUfwTEFb3wqr4ftXNm28S9UGTsHe6p+8icE8BkPuGrjoyiN7f8j1Rplcawyo5sMl
hNBr+ablVXuKrDP23ariaQ==
`protect END_PROTECTED
