`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9YwkZ1eSSvEfeb0lVGgIWTL/KoioaXapdIx+pAp5xEo5DPhg4JbpK1dom0+V+QK
i0seLSsMUGhORA4GbqPsbkRkyajGFw3NluHJWEodRMigwXApLFosqrES3dFg4Gzk
NRBhqgwcDCzkqJJXQiTVdexQTl/hexR+M/scEpwkzQsejLNSWJrT1L7WY8bcbyHk
9bKAdpzvwG/XkXkPFt6jxN7QnH0rs6jZ6OUf5hA5uvs9SjSolcLtLLIifUQ++0ER
I1RKbh1nNG6OhEr1YsjojU1kHXngN163UaWQZ/HcS1tcK0cpSVBoYeY3+KQiDebm
UDc3pEfMZgnPxbzhR2w4pxYPeMWNgvmJ0GJw8s8fvbI+dertMocyCxUR5UmAnwTv
WWzns5HOknY6EuTd+IYg1E3Gi9gYLacXEes5YoNkRAW0MFmGG8cSDXZxxkx0/IIZ
4P2srFsyiHVeLpQXRx5TCmHDK3rTG6xwPP6QNsr86IC9Sr7q2QOOmDYIx4PLsvHw
tv7N9ubYr1PnDr6pvUpIcoFp4Cmz5ow0GShsdOzuYeBYEnNcMTFGvTLThza6PZlr
BNMZavyx3zo0UUDdR2KavOaii1LPm9PCi7b6xi3lhDssDNbTqcsZ8c4bD4TqfqN1
dXa2ssmg30tVXTVkTK7BUYZv36tGx+TwAK5zq9fIvQNZMiLBaSmkCgJ8tkbcgLkr
HU2y7JqOsdnBWK21nnXb9ikztSrwPVLn9muyaC+Z7PmGmxsrGcI0wj0calDetf/6
7/NVa6MCQHPGlPlBYN55LTI33rRBGXv0TAc3DYEkQU0AjpeN5mAKdzL7XyT/U9PM
pSfjKU7OAQ7Z/H9e4O8pdKk7stUVnmHqb27S7YWhn5Cgc+g5bM1AdGiAMkm0plsd
8Ui4dBsvuthMg/7VEFWUTyJB1MEh/n1ubyzGZsBL9ro8eaI2gXR1kwW1cstAh+a/
hKQM7K5n7ybIUNkkU6dnDP9TCPkP6o2zPPnRYGWUgDPLAr3SebC6SgGo2YkNixTe
MFMH50fN6jd9omvCE/hirgDCrPww+tHXIbNX7YsjzEw2Vl6rQHFpoq+KXcw5CyuZ
w/qSc7TFwHV9cEVM8EuNOraTO3cwjvBnJul4puJQBFKWJhTQqS/lboy/jZQizOKt
qBv+TTluN2xuRXsZUbT2rjDZEafIRxawEos/rtdyLafgzs7XA3XBVz9IXxEbo6m1
`protect END_PROTECTED
