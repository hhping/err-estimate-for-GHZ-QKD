`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCOKNEUT7eF/mLiElJu+msxKXJSw2qJS/jCVtvN+xqJaic1dQrMfmUeM+v1q3uu9
bFHifu3Widag6rX9cPtUt1oKwWjljJaGD9dgc1jUjyCt1XmfADRaY+kdZs0mIwRr
9rMkvWsf5yPcFhmr2i6pnC+LbFg6QTPo/9mespofTs1cDXJB7mmADE2gNAaUqakR
bbCsCwxhA4IHn0YinxstOVj036uyxTmaephdxhTpNb+zoHwiIRoRs2MDrLM5exul
VNIhPCpT1vc0+TSiLO8Vm3ZqRTqzcTg2TZSHsO/9KKgAJFfmYb0dBKoKPug/5uH7
3Z/adnWCBodtTJkuTiMDZxFE1BuAUuwREPaZBelrNsBYC3i32lmIPmfKYRHfb6Wr
zMtRCk47kizC5ZjeeEXYvM8MCSeoggCebSuTpgxOKyodPkzb874G+5+Rvgs19D2k
s4/Pnp+0BENRRDW8bSDHabf0tgeeo6ydAP4M3EsKrxVdDZEcXegKATozi2H1wjg4
vA66l7T7Q5HyApfkF3k18oampTudpsLBhSzdNkd2uPTs5azWEMTiVjknF9o810Y3
gALoWMQ75pw7L+gBGUti/1LbLBOu4wcF5jd9+zUYWNlngG3iJ0QUP7Jhul4/QZ3f
/4V0kGW2xIY5USSeyWeLuCws3Tax/LfVjMu8gBE9W7RfXQJgcYLqsLU2kOx7ekDW
wAM2Dukmn8kEmvme6v32gpLYW2YUSCr08t4NgYxYfwVJX28klA3ZzalqLED05IXo
KFIJwUxRM4BEZZeQHJsIcwRkPnf6TlDSK1HwXCYyZ2WVsbBrggTf2Y76gN/AwRIg
F9K5S+8fEXGrNb7xE+9/YYviOh1/zGl2dN76fCINvJDCcQjJQHjgdWYpM4pKOg7W
UX11TomirCKYUgrCILKZrBJxO5L4bmhRceMw2hCWlQzBsc4ouxUBlTXPlUOXwrI5
rDh+FdklK08aaW5RS6EGBJpWjFYKFaEa91y/kcnxdtzWB2CZnzxPqnyYYkUnsd0u
tH2SFboAEeTRrpEEQDVXessXJIunreWRM7tLXN2f9HXfcLxRontVEh69RIHqyLM4
`protect END_PROTECTED
