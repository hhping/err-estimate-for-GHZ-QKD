`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XzxWEoOHExmuZD20u0J9TKjcTh/8BK4DhWoioSWVfgfT3cERdOCDvUkfJUEdvoD
nOmvoFkCGWEZf8a4ZicI2zZPY0v1WufmH3nf9OiqzWfdbrgRbLQ52wPx4L1t1G40
EmxOCyn3GLDnQTRZfmd0DoXAd4u6YbwsTTqptTaZAAjS+6bwumAn/lfFIsMKKccW
bigfKh9eQ2WsiHeqv2DQWuYTa8rAvZCETBTashkBxhNa6ZalMp0gPWKlx8CZ9Kfv
9cJurK9RUFgup4fed4ytyWoa0Lo+TB6dpFZPMX+UseWULt5GvT/Am9RqHhO6IMic
evZNZr5LlFIrLcDDU2H6zRLviouTYP2GomDhrlk378xqZfhJ8Y/+VWL/MAvchwUu
6cQO24nS58pscLPuWNp+MnJkVRDAnznth1HoJBOhCjroMMN2cWxESHXWbBCdRnNk
1pEubQfncm0iy9XOM8ItE1scQBBAEWuxwBdqWeMP5uk2dn95HcJAgdw0BTKD7j1I
pLLFkzKgz0P/n5kpgrUKDRSs7Zolj8M75K5hzfCQgp9/7cl7F7GilmQzA+RPMdQQ
CZQKq7Odl8SA0OorZ+FlEvPErHiKSBvMWI7CV2Nv6k0=
`protect END_PROTECTED
