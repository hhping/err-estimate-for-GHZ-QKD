`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqeaxMiy2/D2hxBeXd12wSJGaQ5TxNqqdEXYvmrMA023DEte5hQdFukLPkvEV1po
JXl6L7WkNIj7JLw8WVUE0crPGzwhb7AGhbkzOEMag+4mFWrEJq2Z4efxVCVpWzZM
yhzT3leQCL6KPFJWrLycP2BsSOZ+nRk6c/G1hAf4iExqBMKLaRxEET+EEElacP7+
Q3c8b5ZF+yaEzST3kpj/maplYSG9Cf6SgjOxb06z41jqmuAKLSiwewC58V8P6/uZ
sNU27TD44OGr3PBu7bifK81V7Oc1Ayy+mwLSdORY+S96880gllzrt0OTZJcxNsn0
/YP+E6r5RyQgqYNoBTWiHUHwQs3vejDIPCRElCwnDWstAnLeuxnWcRB14ecvHTd4
j2pcp6ERxgM0boPNiF9GPiMs5LYZD1qcmReDCsul9X/gH5ykxViFPjP1/ijyzXWs
LGChVHFELq2JAuNecBrCwtis0lxnh4gtr9zazdv06t55HxKHyQtfL4I7ivc+dkW/
R4XeX259ECitKVtnLHA9I6Irvo7pU8Xv5NZDbsXzUn27yFsUTVrfguvdtiPAcraw
FjgASEcs10TOpiNZ+BXaFrSWN1EMvdj7V8xYPc7iM2hl/Lg6mfPu2qfklpxu58V2
eWcYLbGisIDZPbq6OhwplJh9a7WcSHmZE7Qvcji5AgiXKfJqbdB1z1mouRsu452M
hr5NJsVNHjsAFqY6jkGdgXDJLqgzZvGATDBrGZVRJ2JczwD6HTghWl4J640qcAvy
gjVHe5Lgb7wAvji+6xx3w/4ScE6vHNdW/009guSsqOCb0jHY3lotUEhkTClBWsF4
uMm8MAdsBRdp0sn7oCywgRvXt8IjDzezcow6HdsjkEPEpGqE03BL6kMjgu80KMih
+meiJw7hreDLP8XSI8mbi0Nwl3PgvbaLMauz1DvhyFIDiFfcTL7ZEowydp86X2dy
y0bjJt4CNY67fLcHxx9tTMhHGeYRw90gE8zRzHnZ6Qpt6QG6SRBR/kaHDjRyFS+1
vK8hHBs+r+9B4PKRb8n6jRrcxT/EkHNgDlzmUQApY5tItSV+EYKQEyd8fZmvFgG3
WyTFUHu0b43yBDIX705aSh9DXaYQZgeWSbi8q+9L264zQ2XpDReSZmZyuCR5/v+R
57H1EXqrJt8dVVSPec8dAA==
`protect END_PROTECTED
