`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+wdq0LxC+f4egQFG7dXZLWTaRQVZFJLhs3JMtFsnOb9/2PMuWG1t8hiF56t76tG
a83rvW0uJorl1PwZb+FJUHAgwIbRRUJdyciZoTjLYpQKEWMWGjg51RVd2qjt5czp
c+X3amjcvQZQOU1zS+INIhJmYzoIELsU3UStTFco5X8OZsMaS5osmeWYB76r5Cic
cnfk1KChfnOBf+3XZ7ZltC7nQvtTbSnOxdmzE02oRBZSgH/j159PazMZRY7PpJKE
0+6+MSPNM1DxSfkhhFI994GfdkTMrcyTgvXfAqaeBnHG45YJZepOgz1sVyQ1WzH4
qduqqPY7fn1Hd28DpuSuoVkYRgR4YLriK7x6/l+1YF1cs2A98ocNQdcFeGBIhO+u
B7X7W3JVVIo7PE3+3Hp76UdRZSD4PH/DpUcROpVd0ExXC+d+Wn2WRJFq/XQbVWSD
ubM+mQs6a7Xnk4wsSg1QlbHU7aH554lvcyvfQmIy4mGkUkIx6MkR5uLEtUqTD+vo
HSDBny3Ewj0CKRf9E6Uv5XIIjubP7PSJgMROdAb3NXvhIsnZ2HEcJf9n0BVm1X1N
9tTjdSzXVWIaAOr6Nkr9p66SdMHwdYf6NoL8SW3q8PwloaBZhsVIiXr4GxulJeMb
uLDYc2DCjoxdqKJV1l/3XtXU/PmYjZYTZAlCOeJerXt0T3Mc/GsfX3pei1DbNuB0
xEPzjlftSaV6Zl4OCHVYL3ILeC80ILRKg93d/oRbsoojwOZ7OxbF5k9/Sz/TaFab
3Cn2K4Nyk9Ew6VaijcGtIsWqZ8yamQN5lx6+5ssrsjxsZCxvudtPLVrc1xaZ7PwC
w2e3L+njHgS6OltP8CC6MFTfDjpX3DO9gdOHhRMyeZC4EFLQO3wxta1zHNvpWc4s
FShs6S8Dw2y56UiLzgWWTZcEXew7/nNcZ5DqOwpuOA+sTydyCqV/fYaTZIa5ffCo
HN8iunnMQxrwEn1JmQ/JlZARc4uBKWU7W6wswBrShKQOKNAGmCLqNA8MM0hZaEBg
YI3XGLvcjur8xd3pJoEURCbas6vgaJSzSvSACLy8nHMYhd1QdbTMft4wGQMGX6cD
3XJMeMt8AjQ47mrZM0bciDKIzgQsui8bysq9ya2DL+NgpIbgoxEdZIbmGHG+eYfn
PFC42w4UqnHLqcCD9S7k2yFUp9XWssF8usLDn2RQDcZG6+gU6ch9pJhwdkkmSRRS
TFicvdN36Ph/hbWtyYXuD/6sGL7tdt/4e3X/K5GvkqGNXTTIOSGLjBl3Ol0YSmyF
`protect END_PROTECTED
