`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvtvLRSV39yZpMd6WLX2/yE7zaRE3me7Pvs7obG9XV5RKk8vX/N7065LahbNK1LM
Zp3P2hQGgJSD5518vSGeGdPhECINyHuWT1P2sbg0L8CNaltDOqSkPKK54Ir3xQIC
9smRaSTW9pNt8TgxKFeO728iSMetGiphBGxMZYBj/t9mV+/16a0IIJCDQzYS7uMG
iDnVNFfJ7FazfWlt2iyavz/3FkKHVdcLBAo8H/+wp+49mrtwzufwcDard7BaIG0H
xa4tjPJu6G1fr0dyh8cLkQ3+q6RupFMmS9co2d4H6J/gu4xpz0YIeqOK2EvsEwBE
QIDcMdVd63LYlZsHOlCRKkatX+2DRjo5WMpx2n1yI8t5fQ4DfvVJkoK49uP8jdBu
itcEI20tMgZmFv0uF6F34LWafltU3tCyCE66Q5UQojZo5e6QJ33cmtoZYmZZjP27
XL7CsSyc+2qRrrbXTacc2C2gofdfjauDJ6TG1kEl9zrSb3kKIdnWTRJyJxNgcNF6
JPDQ/Bv6fXwQLo918xiuXYfcJ9+j22m9cW6qP5YaaVHN3d0eWHZn7i2jvZSyI8Nc
`protect END_PROTECTED
