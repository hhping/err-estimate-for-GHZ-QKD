`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zz3wzMSBkMEOpPZVxTO2iFEDvfjmPHdf+TxPI8snPoLPSCqv7TtGabfn4YsAFezb
9U/BQYRm0wtijgq+ek4OEgbOrVYq5+A6mVRrq4YFUaaVZvUXNQEme1vZr4o+VttU
5jITFGLVog29U6z2JoM5wFYvSmme5UU95dwpVABdIj0IaIkwICYb4d8wGtJnOT2w
loLmmJNtRbAQtBXdP+O/VfsLKlY6EHfKi/HJfSqkrpP0hycgTPFwS3QfcSi8QNzF
BI+z7EsChQEk5Cozxyig7/YfWYeSC+Y3GYOsZ6K03zY3ltfyXuV/e5Fi2u2JYEms
4vgDVbWX/6NTikdo2pgsHMwVAoKlwY9o1Rv9ma1PDq+hhkXARcqsHfU04ubFYdBz
5qzC2PYaNXxyxVlAGYGpEQ==
`protect END_PROTECTED
