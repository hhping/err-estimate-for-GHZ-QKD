`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEvTXLOZTuLt0MNzkFmgaFZv9LSpq0msuMOFOelXgHKlGpgDOdSyZaR087hfMUXb
T4J6yy6GeZ+RV84MIsCMEQFySPdNvLXbxQ0lPXZeRWv0jRNguQFHtsOCMW5cQsmN
Rd5nRgB5Uc1Hcpg/I+bSbGyTWAuplLEcYoE+FemiNGEif1nVw3Sn5TaOdA2Ha4SW
AJYdxaCGIyH3UpejW4q/A8FZb14YtXxxZuNMzxY9fkqBiSRZyXXI0hlFi1RPRETO
aBMMn/eXPaR9dgjyXZAS/ap5+HEUjlH3HEz25ZC2na1zCrhmDK0J7fXyu8kvqlR6
tdfRyaRUJvb1bsv16msK/HXuKj3KKBFTL3TJIyYX1rv5DJw5mPEOWsCSO6ekoUDu
7yYZ6nI0/kU3BvQSzmmqvPfDBJsU2uKejTyPTXKx94kzIV07+h4o9gDJPOo/89sV
fnFY+Xb3R15gCbt7Rbqt/eRPlhHZHxPbiQIHU+qJOaOdPtLH2mTQ1/f4e7nQt2w+
MswW6CVPvO7eYIi2KJ/x08wweDBe4RSYwKgqa9HR8PSii3or/uHLJBDHJWFxVU7O
4gJ82UcRsPLlKtnvYG9k3RrFC4Ht0CH4jIN+/zEd25gDq954ot0bqhJVsKimsvT0
sZVAUSAiAQry3uv0qXPGaQPyjPlNO7qRcKCsQAtbk+9X1PZ1Zogic98r+wrKjQ5z
7/n7KFNIAT8CD7RI/rFVIg==
`protect END_PROTECTED
