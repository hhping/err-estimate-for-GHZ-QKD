`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6x9YP/+j/+YwuHuAgsrn7MdYQag7cIFexLczrutcS2a7UpKow+0TFbI54Zk+dwI
sxlortSZ4VToVHnLWt5S/19YcKizA1hawcfPjPX+uZnFAFta1QbC9sUbak+umEBe
ogo9fhlE3Z8N+cdP0Yf/cjFSUdHXV1wyqU8A48z8BeAMmr+6NINd8iLskZTwxSYt
KVpYV1few0EotX+q7mKVcFc1KcBdm9lwJsOZaeT5lmHApqe03EGQhjlnNd5a6Ymy
0HSQPxIsaL7NYJDbj2yxgF1Ntyj/Rnlc/VfsUIpVH9Zqh9X6S2A25TF6lgNr33hT
Ag+FLekmDTyjuiBqR4TTZqSwU0u8FbKFZJYrZZ12dmQ9kFwvgJiI85CMiEfDBorQ
Cc4bvFOrt8mWuhowELxLNtInpBhfh4mYCXWdazjnKPF3dJ/qdkdqs07AYUgpSUq+
beUWiNpS+dVVtvLiSfKB0zfhq4ezn6FcgqS58I5vsj7Txh+PFog1NXyaJYfSbRmR
R9JQfK8kyBGgDOsq6aRV+0lfvaZhVNZhqb/x+pOtPvL+AtMaUy1z7v90dLqANPBX
FWbYTQibKCr1XHhncOXTJMtcLxlOX1cLFJcNdmm3qDGSJdKklfVIkcYC38OFEFfK
KFSbhyOuKlHYIZTe9Rnive2RCWuiBxbgqygoHwsWXNqOvLGwsXsRb7Fv7tv6ATA2
+RBwKwa8ZuQx63UrrA2zNaQt40EWFz5rtG8vJZE3WMS5Z9Zf2I39rU8u+PlHOAd1
VlFcZmMJg4vhPd0eK35Ku8e4sRGnShAFSEZAMaiaX3ThkhSN6sh7y251K0ocrxVI
EdVQ52y17A37RZSzZeYpjP5ZXsKhBo3KELppgcnksZ8wCbBKfsN0smYQxSQnIwXD
3YnUMoD1mbKgn4/Aqs1BxP2WsE94MR5SY0gDhpF3FCXLped8X2w90cdiYLi2zhc1
mfcWCmbfa/lR1rczrDJDpsInH2OrFSn8haMuxIyfPnLmUBxG2OzO0njE/5kDyHAq
+McxHG6wVbcs4bYqSHXz8yhwsO+e3yIYZWXwWOSE6Fxy6PRxstpqOYUir5Gy0e8R
/dj+wkWSSeaMV+eYCzqkDyfHC7RRL/nGR/8pe8tjyYEqZHcueOZ9y2ZfxEw3WeLa
lp137cqX4eHximMEdOVmZjX37YYlCbJDYX+jJOovzd6juUokiFxgsIEGfdYlNvw8
Drdzu2wITrkLdHKkQuQqGZ+H5U0tG697C+jjYTQkwBmhiq8QcYJ0+7cV5O49gRGG
QmEuCLDZictElcMIvnsApihGmk61Ey3iGyN+tHurY2Fp8q+xud5vr5wEBD8jrsvG
m5aJCPyPQqt0FA4ZLE93ZyEVuurcAhDgbXll+Zp4SRT6xd3a01N7kRR1fH0nslO8
+rbEoVMCZxKMLAM7ql7hRZp5Nr6GI8vqsuAaWDgOIjpLrewKHNCG+m26XWRzKzpm
2U8UiquvQRwJUVFQPc0t4664eLJiSiroZoB1UEAmGXWcO5VjN7y10iL8nH0cqNLq
lJqMOznEHLtUhS+HiPOqDge/hgaG9gUmAkDazf/hWbS1fxflgTg8VAXkVSfNpk2/
5StGINM/dBOnAsDhQJQiFOxu8Txug/b8+2juRjHODGcTE3n31CdoKS9kWv0EZL/D
JTOIN8YrlcXUsOTRUqU94lqWQZZ5K+RUEiyYV7d3PFL4biPMfTWFUT0U37lL6smi
HhrqINbPgqH6htUh9p8pZ83RRkbreTdDwOGV/UD4i4qjN3YNrMsB8gr78P/A7pRK
CPrWwTmhiQTIszMYgo25GkZDhSpw8FoLCldOAGkGeUI8qUg2+/k0R18LqgFwPbxi
FfRB4odZD/VFa1wdb1UFafNWMfQjXmJWVn7qIpexEnHFn4uHT9VApv0S5tbA5WTT
hNmkpLJjFFfy1udYKeqBIlVcV4TPRN7n5aenU28+vIdEhMK2b5mXDrlVDwT0crE+
iKMTNTkL7YZqzIzpJoz0SpxvavdM5CidPNvbvFGJJ5DYQIFofsNc0nEkwoF0+KiI
hbrTQhBEd5Bipb42nrmPURUzUPoRUjBM4OwqFDeDMAZwhHJMfaGWptLh0VJPjg81
VghVXkLtCl+jawrcSW+xInfFmFBFeWung/T1qr4ePy96PzstNIzLCOEaZENjD41L
Tfo9OKfi/8xg206jqYjrNh8BhCGouCYno3pqk2gtSpc5/grpHPpY611NChN99CHb
iZAly8K7Mn4A+67K5jHeFFuNgwywGJm8x3sOB0C1UCOv8tHy9349BP/fNRCNClnN
0SCzcwzrOlbg8+Ahq+opMRvw2v4YUy5MoACpaMuvx9HAw9eWA0iMaKsu9LfdDEpQ
GnvfuusTz45p4l2irXufv9qu6+CUCTVKLyCyugtFc4nLtd89lyZq2mvMLDQ/2mfP
8BEvHQnr8FKFPMCoAT7wW91SegNYDgB8OanYvDsjXsFAhSAAv6VlmCpXLkIC+EnA
jAW4wpJGIgaTUzs1G4d25sDCHCYBI4lEVfcb5vxajR70/lk1fDFdGpb0Oiv2EeKF
usVT5a/2TskMI4BP5Dj4YD6AuWnC2yjpMi2PKoGaYmHDwX4AxArHFVkNLFC+aQUV
Zfm0F0T+iUhDljWn2G//InvMJdtVbxSAORLx4N3S8YPkqyWBTrXT7kkP4u5lXlzZ
kXB+uZcaTk+7BvVNxNrT3I2r5QaAL6V7RuRMF+GAGKTpvouLjR2BwSVBz4ocmRgt
tWWRu/poYFk1yi7rFzh43XNKknBmrCOyrwjbrhOJaGCdVIBxnseGYZpbGZovDkED
iQEaFpSnW84chvPO2SNp3ySpGBNNtVBuEwkaTFT4b7rrdAsblNRdVgIgw6UhhA0s
pZsqhde6Z38GecWmloLcc5aCttP2qMPMMwARGGMo+L1Hyz/j6Hq23SxTayp6uDCw
5l4ug7raTuD6sRNh+5lC3Ufzl+Q26JMaW715o6+Gcz+iGOaHBDeS1tRLRZe+oYlZ
OoXka4jttPGgUQc+a7kUMIpOboZxlWw3gAD5DnAFxzBnEZGgUikYOtTCJw8H0mYk
zYva/Y+qkuYVwIqK0wlV4A==
`protect END_PROTECTED
