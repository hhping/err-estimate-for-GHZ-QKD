`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kOz6EfIsfIPSuKaNKZDu1yTA14UWdd1YnMSM8Q795dnMGwqOEBoR/2+6bdMH4HBS
c2Z8ti5d85Ydn918OjdSRCLXi4c8TaHuT1tFyptP16YtnIWAYfGyhovgl//U3Y/s
7blTbc0BH3ICntlrDMFn6RI8Moor1QITM4CoXQOqAuTu5oQ/fl9UGMUBWDFi2J6d
wQ+IiKRa3fY+oQx2EvtM6YRKRX8DK61vRPUEFoocMRHxxN/W9KYfHZC9eLJfSTs3
Eg/gykOvYaD2jRyzURtmZFdQzHd4anqJmGx/SQOLr1FDRZyYZfFme8/N4feGxuwo
uRbypL2joP996uggbYTyMN9BGIbOwiw2iD3WfOe/P5BypkzNPyQUFo9xXzNXNHq/
uR0DDgYIrVAhAYJUViVloKgo+jFGwws5pHaF3Gkm2dRgIW8Eke0oZgHG6eTb1SH2
ZYDuIhe4LeohPqjFWU/gnDyoGmkHuSC6zJbBpoRC9iGd1o9KDMXB1k5X5DblVD9+
gvB1lOAaS3y4hMd2IU0IvYJg/dE5/34yYQfoRqgZtWkQKA1d+uu8KdnQWpU8yH/I
xsYPMoPU0mxZKQrEokp2iIIi67+Wn2VibuTz0J8gRVMMJIkF83PPWQfXGK9Mwz52
z1DwuPBF5/rwUShyqmMEk+U2pamTrZCj1LpzUU9MgR4wt6EW4BuSOG44qFw2Ys06
SkojzAFq3hdRTxJTSX56ALJjPzf3tJvtlS3ekbDqIfByLrX09H99Gw74SSzztkKC
Afe/gg6uLJkCTQ9uCUlAdZI1vL5KpEabk9pU9ZLrtYyzEK/vDqkLmOey+I4Fa0Tm
aVtDyUoxW4N0tz8i83rO3lJlI0H2kCItFyoXMrV3qnzgRRj1RdiJOaDe9esRsgvt
84TGpL1O+dSbMtDbX2yV4GjO61YEGsDwaNW0hvNPctdic9KmW1bfLxLuHXxjh5o6
lmmQaZJF8hw1tSCtaV9l7PKPsYeS4nx+X3v5ConxtVsq+xCJwwdqca8O/9OiqWQD
T2quvRvNLfPKA4XDexIE0Q==
`protect END_PROTECTED
