`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1Gc0RJnjj2iwSZOXIUMyn9YHhdP3QFyloE1Vn+vXs03nw3a6hntRfVPHAONdu99
lGz9VVQforxC3OtzobMAB5Bn9DakKskVif0u1lq5wrQ6pWiVEWIKpvv7YGfQIYqP
6pUrlXh2rAnivXW3YVIaLZby0qhg4DDIaOrEdJStmV/gs/sPppep54LlbbvQ9gH0
x6g7Pnb+/51eQDvK4HK7VgkpG7qBqcywIJuw+a+w1A7BXJuAq9OGc1M71nnnmIqs
SPNK4u+kgzMbweSIzLWGlb5SdaDVTSQdPlYk0G6w28fwV4w10X1QL+sHPmmqX8qv
2E1pCVc4Jjy0GbSB2WqH0NsDlaS4ghwt53NKUcvvme2clRhcXYypGXgAoKuppx1U
UXMj+KKIv6oi8m0vlf5GolxhzwZNtGrwTMPNYgndKsiOIJOKcGdqUTKohwnncHlK
vuN5pdxTykGpbfQZWAVBBEo95MpCnxJARRMwIeL5r9aNWhD76KbEvtoAS3uvA9Vo
T+09ZD5dLBsPhkZvY9vTD9yQullhRR6HmvsQgXyRZEtQzQMBvAbyM5WyV8rv/LgE
poXtcsQhuT9df/NeioUDUnWjD13ov/61Qyb0p0zB7iA626mxIqarRt/w+wMMWrx3
5RwBYYVdYuUNr3AfaVNyVleEgzknnoBcvbn4+iB3iaftIMrMiLufEhXBdPSodUHl
RnMZf1v9416A3k7b2vVSFIrNq6i1qh0Xd7RIVSMrA9Y8A6+AMRozn4s9IdXkEfux
KEbUvPx18wWVAGNmjVsyx+RnYFnUYPfGwQzanDIAwLf9uzxAMBcPFun906UqWUYK
q3Jc+0f2uPJYy6+NjJjACGGFtrNLx9VDRo44A15Edu/RDYCTBo7beoU3xzC9oAyV
S+NZiEcI/oAKlUemDQFPKQ==
`protect END_PROTECTED
