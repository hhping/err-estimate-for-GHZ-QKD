`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBPyqzy51zjGGkFlZ3WYY38DyaW1ARxwPXVPO5TGpU/ZID0qNJ+QQRP+EEZ4TdKk
AmAHfEQBMjqh3ngbYG6hPZxWGYun712Vpg675LaadwGZseBI01cRuydPSN2nmfuA
lI6V3GCie2INwuu0rsJzCyxnWHOHOHw7npRvQlTOwKIBqoedJXnbQneb4hZuaocH
X0ZGJri2tFH7OtaDxwCyYxgtlpRHrSF8BxyKmdqbvW0WcxHE77DI22tkA68zA7YT
0hhq/clv2Zib+NTq/Ai1w0rT2eyhLk0/5kLpOm6ESyj8XPMX1FXkK/uA0n+9Af76
sG1PM9l9zyY9p5mK+1pFdZESQKPDxuqTx362Fa6OjmKf06Sp4Ob3jK9+Oiizh+4Z
A1Uml2b1iUZPZZnIcELnnanGXW2FDxL5KHChsmxTsGEwJd0OHk/H47OrsEtNJbg7
b5cEndsqOCG6r7f08XyquCWTX631yAa3IBbCSDLaMVw5+4AG/d5LDbBvBxJtN1Ct
z9k7as6Jjx8N/0f2hka4BGSyR/zZtysXQERMNoVfgTzqYwV6bq1BU4n62PglHZjx
7CRZ8bnXL80qjTa3x39DJ1eBQ3yNeHAooEuoSboDzL6jj8yWVp8+21VKYA8whHjr
pRmVgBatO38Tp/qK2rZI6t8vJqP+Zjc53rIbYXjnP28=
`protect END_PROTECTED
