`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AT5FW12iXOvEPJUdlcueR5iSIzhWIuQ3b4JzTnxI18nFlhXQ0hrsKs526PmkIfSx
qzp+f/ftUl0zAKr+Q7J2WwMZ/1aLjEEkD8P74Bf73K8TNdwN4BfnEVN0UrsfxtQP
5f2ZjgWh+w0TUGpOz7TNXFzogyFV5PVPN7TPgrVQTdNKyZE0x+NnWg8mZWRAl9Fu
8npjNVJBz13yM4QvLOkiy+4DpQLA5kh4mcmCMLgEjAWeUo2HL7QndbUFKHtzvcdW
NdHXv7EYUv1W2n47bmXq5iiOTQV9Cl+Sm4FSktNkUEDak27Bu1zsAwlTMWpjhyP3
wnKt9o+sj6wKTUOXz9KZQNdQ+pv4i638RZjQX1qU1vdG+o4vCwJ7gOri14Jc1qtS
N3la1592xyV/epuuMDfBf7Ky5Uq9T7J6q9eh/P9gF/vipeqFM119x8Q+bXUM1vWJ
PBZf14XUuCcx+sflnGH+xFsiqSJLSd+S8pJB/770mceosxy7HjapPPkCe2UVyQJC
StTkKz5U+UHa/glfjBkGer73QQXUIeUktPeIQ7hJUvc8hFk9dlcu8MUUimokdl+K
vRJuGFg+jPKIY31NgTY8ejrfOr+I5WIh91LgkZSwznVu/cHf3WNPJ43fKFkGeXqh
eRk3yXAQp+gfS9Uw32x6u7mTHTbOLNJY9qoUJg+iPIZ1INfFMthmNqI8tFJtrrvI
saFIMun3xNwHEJjR85pMVKO02d1TFKi5gxusUksQFf6qS2ZSMlQyjZ/GnfnpIwgk
YklcYgBPOSKTV5IogT/0oSlJqTFmu9XKpI+w6AUAs22pkjSPxaJbU9WkgzJYqP+6
Yj0imOeLuBlt9xUGOg2YEBv8tyyaLB01W1KuQUpnXZZiz9r9mVerNVRFpXRhPpMT
TBirDO5O2oAVs8dy8eNTQyMD5qTsu9032S1LmnGDrSriqwzJx/XW6oNNMvtqtBGh
RgEf0L54MGAesJdfqNhd0ZTVpu/7YRntQH6eMRy5JoWdVJQseN/g2zji8IL+BIun
GjkbiSwvppcsPYzfpTbRjqxS6rpXRCyoy67jKYfbIUIgX8hMtuJm7YnPOPekJUPb
olO2pKPA1m6TgieMpUJLEZ+OIZBdac7mauqOuHmYqwfIJ987PZhrgB8wJ8Qj0u+D
i7gP0iNqo594gIKACh8m32n13eGXJmpzuh8txF8uQ7s7zADt/svPGDsAGUsV/gEB
joKOpdc62SduxvnS32d/UqktilB1sGBayYrKUONk3cc95IJ+k4dZHcTgvb0xmJpd
tOtYFb8QX1DqsP/ttfvAQNx2gKGMdGs0gMlxtWHLat6rOUw3ZYQWPa247Cx5edAY
A5VTlFl98HDP8mQrgRo9xGA/GSDmWJv7wsLBcwNdwiKXMyGRDtvqE9rGOYrHzgnb
8PoXICcrLkF/J4YW1bfGykMV7eIy3cwhiW/e6b0OKoPJCPOFEZV6G3mM5fDgXhok
QKPiJ/9cOe1puI8Y+CgYHLkbcGRz74x9QmkOUuvgOE3Kv0li7lqPcq3z1MfLQH5b
1kgRipIPj8vFVQGrSLmD1Y4e/61nvwwG5Qvf2TVlIbzVVrlYaa5gDjbosfR8StOG
fay8FiO37cW3RBN8Q2D3AxYNBds+cEQGTjbiFmMq9NrH3EUttUkznUSp9aIiCXhb
7SaRL6Fb0Crj/9i1NdTP7oTe70ALNmlY7hxL4K1m+chueNKRKcWupWmwr+cPVAst
iLal1wTBv4Xx7ueCue2OfBhZ1IYYQj+nKGmPZdsZPsie4r5Kt8i/sxUleBwhsMs1
ydXdLlggTfxOFfn69M5YuFB6vAHLk3uNiudI4fVOfuEff413fWVx9NtBQCevjWSu
ZmybIupxYG+WCkZFU2ZCOnPCxbv9St/76wivB7GDzrwycb5jd9M6zNeufsjEGKLR
yr6TskcDcE5RYZsoe/t5go/DgJoWtas1dhe4L9bUHwwMWe1ZdyQp0/eOuVZFm1DE
oJi7EEZ2PEb/34PcVM2jZovFgTg9SegjptKc3JNiF/XiF9aCCq5xpfc2+gjBceJK
TKdnzUZoB6Ew3pFAahghN7P91VDn3DW0UtDVZCrj0NuSuva+i19KWLH3mPaN1u35
jsVWqhlPLQdBXwBBaayJFkuvj8VtNshuEnb2R7rydNjnXoizBKcvL5fznECkbcHo
2UWsRKQOO0r+Jm/SH03rOAcwHzBjzKC5mEHjJ1E7dLutEfboWV4TTtX8CwdODQUc
auwsO0eNR/2D8z6QlmcXxvlR7BBAy6QLuijxzBlku59ybk/d8YmI4zsOZj9gsKo1
LX+mkgHrqHm5cZcn8Lcn3ETc3i6uIiMc44W4iF+650uZvQv4kRmgg+pksJzRB4O3
/RuIJz6EF31urGO1ynBWbkT7LKXIZiG+K9E+XLSPJkYOVSItEWxnNWIUBPu6npLJ
SvE+mTBwVfHagvCRZ+OQbsG1RZeRMmqSBr2U8cXUE/umeWy5mcBA3M59SM8WLvPh
soNGHi0Yf6VrOU4l0docaCRpDZV8FtUI3qJf5Ai/A45zbsgBestZKUCQitTi10pP
ZeclimH8HDGRvEiHLyd7EnSqbCCTkbvVBcTca81aqU73U2cfpU+lzGo3u8KJd/SM
Szu5IBM4Z2lTUTnUiBUKnSGq64QnphthLluVqID6VQINF9SOOV/Rnji5smE3tNVj
RKlKTm6IBZK0gT2aTMRzWjW0To0+GUqfIXb2krf2XooZvW37AtU2UbX2hyQxhb8w
TGj2kvbuEqelDxew8UsgjKr+WJrrNfp4PiWdprcJ2ppHvOTXZGcss7AT2y/YlbQM
GiRSdb5zHq4cW+Y8or8h1vL5RuTaWjspWrnQolkNeLG0XhoyIGAkaPUk+0xH4Lx+
WRCLfA6OLSsENIptgUuSTz/N+w9x6JIS52Q5GOfct/aJIaU4cJ951oYie/5q/64z
zSeds3skxMEInfqd4gKsVUtnfToiiPOcJ+8gi7LWFbo4tjJLPLaGFg6uDQ8DHxXR
byVGL5XV+aDTQTxqx/geCzCi0ACTTPP8DJ0h0hA798ZplE/vSTDIQY+0EBuS+MJ6
gDBqKqybP5gzpAq2NP7Iil494BAFyy5VUXZ3sFMRKPCx5wZOCk5Hi/s+xkTYwdeY
cdHNs2eR4LsCT847sXIaBNEJ8UGE4If9CALvtdxzIMHLEpzW3KZCUN9x2bK4nWKB
VebQlLkAl+D/9pxysGTA9wDUpzUkeBPYJ/moaHJ0CeDay9/KBBAoqY4X+fDV+N5G
ruTAphdoyXqE/imLd5avd5G7Y7Q3tOsX1HdGVBLQcEqB8A4hOOF1L0ZtbwmJ8aNq
SFCKtvuv/psOWeOXm2NOS1KoeejvF8yVYKvSt6MFVBYRdnQY2mo9xzzw6hSk+Mmm
/X8EYdAcCX2WtMh1aQB1uvLRjUJh0s2f/qlVi+2SYxMfWn2u9i1Bviucw+Rl2fU3
XZUwHR9ce4YGvbZ6v9oxp5qJkrjQ5pNFcJEkw7mEscUcW2zr4CC8RVfaSAciuImH
1JbxeHMeg3YuYqAodC4fgRA2CbMZKOJHn1AjZnizOu2PDq07MrC12eTp8PQOJzRz
B9hKmEfMXaf5zlFFft4+ep2TCkGHijgXvY6V60ovtibpyGuFmf1MCbdM/v5BPhzz
1j5O0zYk3TmH63CWJSsnDfKh4b5YiaCRUZkU+UmShjHo0o1zRgHJFG9zSV0Kmbje
06zrKWAkWPTerIR+hw8E0Qqx6fB83HHRLwkL0KrIWCkuKDm9TVt/raie3e64ZUa3
eOuCPECvUtOs+GlAgjrzeaq0zR+1CQIin8094SS5LSPDvMmxHYrnhgslXkLyJjgH
iygA2dsseIx8+a2lOFgdIN5gzUiumD6UjxNcQZqC0n48qyY4+vG2Fh9ASCCuGU2Y
DLXjeDe+JpNO01fymtcUOSmvcDGs49Y5K5EI7wg/9cuoMwCHTlEOnHDxeyFeT7G/
aQhvkEln+mMs/koQqM7PooE+AL4ViKpCcHDRFXGPENOAs1fBbA/CtE23l+pZ+1Kp
eIoaZCkZfZDPxIdZI76pMH0F0eKi29zUClrjlG11+4lJFwHElQESqKmfiJepUPCO
aL5Z5dqZoXiOZ9Z9NXTNtEorcNP9/MnP/fF36xtxbjT8M2Rr32/RsiGwNYL8lYQk
KE+AU4KJwmftn2sibYuCPOAjr1pl4n/nyuCp+mwyTxXsdRkY3XxcnLLNkmW1cQBa
GzUemWg0dKzMIniz6Dijnrg6RMJUkLl2T4zV3EUpR0srwC1aZsAiTr0F3Urj6EKv
7qPD/+S5QUAGFUcrYm+1Wgj2JKjmGOG+bOYgLCA65MGV5f/aCY5qhK4Hi9DfNyg3
I/2+L6qX/9DUTw1f2N7DOPu8IqlYEsjszM2fsZItIlfzEPTNZ0N90aCrFj/+gx/i
z4dUYC+WOkyjncyu+P1x1ES53YZ62FabveNn7wfGUoKL16aBzCPCtL1qQWR3AANc
0FiZqcH6WLlC7ENKawXPPEGwb7fbZs3+KosWMLIo0ZWpzdIcidoqMEiHqHRFbKlG
8MzLqQd4tVEER00xTPeySNMnfZhsR4jkKJ2qo1pr9SVAKblKj24cyLmEIydKYFWD
G1+XuNFhqygG5XcaApGAre/4sX2Blnf0IooswlBQFE57jnXrlSY6qnQ0BhPT+aYF
upaBYpHij8QnBwcbhgEcZxrxlbJHAO8FBxtSB/qkITtI7JKv7w1jwtsNMW0fFTr5
iDZnZjF9MZLwCE8tvDn2ENm5icDMcIyUlK2offrLB0BzNbMEVkv9dBd0lGcRWV6x
C3WqIPP38d5oGL1WrE2dRlPFEcT3RQFjxfFEodaykfzYC+I3IZpve0iuOHT2xCMZ
KsYneJtPXm14zCypySszraC6Kx19WSE55KwV8TeBR/OEgoAD8QPggBRiHVKHuZFA
AeC2YDVcWysllTYcvg7kUiddhwJ9eSOljlh+wcpLS3K7P+jMuyow5dPiMeOsz8ck
/0NV/e3zXCZgHaEXsBoBWcYOlyEP0YikPgXDgmE6OFUhfA+QT1o8DgsaYPCXe09t
etdlFr1yZ9MQ9SQx0z1CrExBJvRSj5I1YwKNQCcnfwqPOV/0hF4cKG0tBUtfo/mF
iTq/7YW9NbiDqpIoGgR8Uvjv62l3bLe2X7dOZ+oJRTYkYnrnqBdKvK2sMJH3jG4U
Gz7rcSRE0OHzewZGFRMi0fC1kZCBniHBbA0WTxYJcOIrDaQJRkhsgrgvad/j1ym8
IgdMTIrHDgXE4hkeydZsOnqAee3ofmBS5sln8D51LKue/oShzuG7r2IUKqdmWzRw
YbkHHgDb2jIt3fUOhotDpulVg0P2IZu21U5AN7ec/hmWq/XEWNckfU9QMaLsmXCr
CEAfKiguTc6QzQZeAuk1zu/b0v/ehxFs7vug13DkOI3nKRKSiMgs9CAkIYNx1LI0
RhFwPlj6uIojDUCQ8eYGBa+lTlve3bWp+P7JaUZyEHS96UDIFOAoqKpVjNAU37L1
UnAOMjHvjGBR5uVeRBfKAyKiv9ExcysLjzSF2cnTnTQAu/YbHQ9aTcN5kTUZ9M2t
1AMv9jGicbNmN2Ioq/6mJghvkrGghabWEKnR00C2u/ZUl6ABf+hDzi2ex4jwbn/q
xWZ7S7eLMbqc3mG9e8RhT2vsZh+k5vJLCOIZ5GX0DsCdWvP2F7R65HZdTEVsIS9k
43DONWWAar5TGdZbRpRmxcvsaxwf44W8N/WvtTiTmxU2LKuWYVV1hCldwXbEZ0oJ
W5xNbEI5p/DDjW0eKCDAjfzEu0PpZs8lpgiGdmQIIKcG4x2pai9yg2Eu7P92OClo
grYJRCetY7IqWYjRoF9maDfTPvNYBye30zSXf9G3eY1F8LeTiehBhUvAYbGRwL+v
XdBQ+ujVeF0QMA//bNUREdIn2tUZyj9gMP+Z2+B4Hnpzk2uhq50FQelLQuvE1xPM
O/qV7EUaN9W98FNPfLnsLK9Yylr88OTdeNcz1f62D+U7RlTmkMZweHP2g5XemQfj
90xKDjYJVBEkYAPuBK5DKZjICu9/weYvBSSW/Yf1mOKjqeBl8rW03880lYXYd30s
IG9o1WFI8cynTm5pC/xDkMlUiZXFbv301FpTGODJ3W38y9T6KQHnVK9q0n6kNbI3
3slQ0+cJn6zgnVmOJMvI4/hYaY6lok9nUVzzJbMeCwYY46sDrVlVSYCqpoZ6yKTU
ix70jjOZH8yw4mXY/swoNbBebmli5xWb+Cq1xj1IQLHdajJ6kmhmCdnGKk6IUbYA
Rox5OR9OnSe1woP0vPeTrNJ1Pn3bRaf3B1VFLbdaIZAtXOyfA1ENNeRZODuZtgzo
mFbd2JKCx5M2pvRgrIOwY3kl5glkE1QXUBkkOzkrLudF7+5ECc1mqjiOhkVeknmT
d0KG6G4nakGrkQMznyv+/RM2vIduIUXqZvKpD5PPQTUsgq5QgI4jyp6p0+jdaMVB
dR1uGLzwcxyy8j9tbN6FVrvJ5rYq5u6nW3/Qfu70ZOV7aYL8ZGWIJqRIjdirXe5V
EOIbtX3pX/6lXcl9qcD2lgoP8TBdSFiVrsqKJ/eyRFeYPLuTSlCBtto6bwmKX6y1
sNYzQOLVkZTbuJsE8N8eMeT4l2DrYt4Ks3s2PfNFDbMNWESMxyYBCIdjfOGb0Xhi
NAg4/jX1b5VXgeTc6Jp1IbHmfOpNpE8+ATDBcabVtcK//Yj6SOk52LTvjhs8cARk
Yib6jiTsu0EPKstrEwmTZUg7qo+t+vIpHqr8rta+3lgqKcAL7xaidZzF5n3hiv0g
q8WwcJ9cGuXo1PexSyzDCyzs8Zt2HdqWQfFBsLwWV15WnssxNgx6yuEV3kitCoLp
g/sTb2LPpEcFfsvxY2xufYobkm4xvwjJatAXPQk7czb5FgDffNeo7BDTY0+arLDk
ZYab5PKH+nz2LlL0GgqlBdY2pIPzbR5IcHEqdvxWeZJOH8hKIvNxibkxO6ayVJ/v
z9HcmeQqgoX28yHR2ozBujzygIXgcPqJyY2FxOSktD6qPr0OdURGO4utbDPmuGpO
nlyKblFbD6a1QceCJdXwW3vHsedIfaM1S5VB5vcD9FoJBYZUXAEEaDqBk9an27wb
wqftRNg9Bb0IC2S7sWAVx1/OEfKBjcV56CFi9m4Oy8jOxgoBl6UG1RCdCDOsVf+N
lrRUcmnr6usTTlduS19HxOtn1H/71UH5TJSCCqnSPFntrdCAuBZAK0/keMPVzHJd
gtzvMucZLYhuuPRQHqXNGnVtlmgKnQ16qHYdWnkWE/iI9eyb1WK9zx3D9o2n/gcC
st/iAzvE5tjfXTzVqFhuluuhoYa83VIC2mNT+wkIHXfUIFU1QkDF6meotWsozJ5t
lNIA2BMJu1hFqhoe870o57+IG7JCd9bfZjoBaEp5ixSJxHRCig/GUGioaBII05IY
/XOxg9r4uou+J9CwFiAfGSBBYuLW/RsMdkGH8O/RsNRek/IFMJRkilLgt+v4iguq
NbLKx6+133B+m83DjeooDdgdO7luPkmw8PhJZJbNXS7h+fvuvqc4kgLXxvCUYqd7
yVRM6cextUfVBCy+TbvxYDb+F90N2JeqmAAktjLfobflwKd9c7OKgcFun4cznqpW
I1EpgFg1S+x326JNeTN0fIMpvZr4CiUVYwbEdZWYJ8uhiq6PNN+xxJu6jDWPtPmx
PN5OMT7UVEE8nNNCnKfoCE8bFhcnG++spmjEGhrhm/2DAfpSmFz3YyHE75/jjCpc
61QRyad/aRh11II5ciX3F8Bhv5kR7tl9qJyERd2VNeauyiLEClwXQiqM9o68bldc
jU9V6zQCyQT0N5+gIqqKBPAz76j82FV01TeCW/DT1hDUwC7NpX5+pSvsW9YXbf//
0wHg789MJ0+s3EPn2NsSAyWBUOZSk+Jk+4uIxVEK+UTOjSQLXOKuH06ifrkp1ntO
XkYuKJAEadln++mgQg1ngN63TlQ8Meh8acdC9FiFkvDAXckgmuWgE+tVyhrOqseG
Xb9x1osssbu9kDo8NZznWYJzqd6NUKUBsqAB1GyNtx6wHr2SWj/NEqybOIiuaiD/
gD15V+HynbfcnBeDYELhyAR8oJjhcQtw0WQykaaruclNQcM3+9i85iLJTyKKY7Fv
wckydZ81zgGoQwz7weaPwvZqRNHlZzFgGhrkIeQuQ53hbWaxTtoXzSJpaZtxMX7Y
FwozR/otybPnB5xBFfyqdD9r7h12C2iL5Pwr6vmr6FAwlCTm8ib5deJg2Qa5tBpf
YtdqpA0To7ctV4T01oSo60Gap+T/mf/tFh4nBobL97QQlZyYIHGeTF5/4pd0mdbG
hBZmfl9yHP/cWADU5hBKkEuDdotpUmbdSLprk+9TcX2DzhVrF/JBwLC8e/9aSMUu
e+jzeFUWREEQX8Hmw1/hswcMsutYhAZfVcsxuAcLZrORGR1OtyXZnz67feFlweIO
lwxWgDy/gw4WdZrLrvIv78EED++c8JVMBFBxInKAmzLRkZVpcczYVHGFyQNvTxfZ
7F5nNvOtZaI/N5FsiHr3wRnhn/LzjPf9180LKU8ohCaScHQj7mSdJCaEDAKyAqbR
Tp9/R+s2CXCD+uj1+kiV6QNvb228TpSSCxtT2G5uEV4lvwqg7faSrWXgyIdNoqPc
P4ggXcNN3oKrBs6NXES7uUVa3iT6CLdIWdXLTCaaeNRKGqen8yfz/bIugQZzDYxQ
wdWvEx1EKg5qHSw7ruuaQnbCGHPDgBgkrAOyN+b5mKyOxJsXdUlDINCWlV71RtcU
JkWM5LtibG9bv62ut22R0W/Mvjz4W8hWrVIH2raeNT6hB2l6nVNoHK977n2WEZN5
+8i5nZV/0sAhf5AI6CYDtNLmY95GGrVW7MC88vAAGPq30GfrmTvy7hS3uyhA1+Vs
pEMiJd0UzFzd8O5fmZY3ll9g+yI+9o5YrAsPT7756Qin18+IHN6oKcQshqxOJ7Jw
JDaP0tyBDmtN7L+9Y1Ue1I8SyVTUYIL2W8l1NtHXYvlfmbba4RTC6+CI/v1QvMBe
U47vP8btilQgcYJvLFEeV/FdVGtuSuLZbyHYGbfSEeawHcRwn0a8gtogLT/4K14h
Vnf3Jw68L0r9l2yWl1rZ7rzkqwkfBpbsKvwkHBnJQFsJylP+IAIofv0AmkOVai7D
XWBLaosYa7bV3WcbeArOqb+ivQESVPBEPmd17Bo9K2yDzSPBBaTwrJN1/yMWUlm2
YOQqAeolH+l6MQNmOSMLp0kAOzFI5tCuRopbAMy/QVpcEx6LaqS71v9RaVFmpBaM
5fDPNJtQolvuwZo2v35SSb8zWjBgAEZUUAKNOb9SLpJIn2fo4aFprkjIzq6XVtTG
UU/0WLL4WxYrOCdM/r5+jy801zSoUdj0DTbp1cybS9vvWOcfoUpxBiZtyT42hDPk
xHXY/wXFwkBrHjh1FFV9VdYCVRvSwelFIRhKsSPAylt4lEs64RoZH7rN7+YWEnI8
+v738W2kc2LEgkkAkREdif1h0MH4pAB5SgNQpzap3rZEtf0/6OE8X3Sguu4KjzL8
1FAANFC6+XfSpvDwK6I4LimP78Mq5/wQCIwaN86lU5TYNCkxBgXJSdrVjRRCygc6
fZQxtoblMMB/oYtnDCckLVZtHCfQjkp74uZZDIEtZE1g5dyONHhvqiJEUQSUfXnm
jK6gYg7a9P+jLrdKbXm46fDNODAkUqMPIvYhSglJK3wyAQXBmRjEX5N0GyY+J3lL
rJyNisfWDxR14ze0g0a0AgRkj9RU42E+CRwxVvaypxo=
`protect END_PROTECTED
