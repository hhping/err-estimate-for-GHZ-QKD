`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxwzoCmTAh/3dT5GMCHg4stqAJH+SyV0eQaIcfLARWFEKypzTsVKpk8NNpkYz+6S
CzL7zpJUXSZ8AatGgVwoUanoYfVOZKkaudMyGaWI1+aHbN2svs643ifm0N+PATx7
qyf8k4HIB7VJpmAbn3iCo4Jl3l7rQdwmUA8zL1qSax4mszdiQcXxvCWs4lB9720U
Zm9NzZIdqPOv8fSuKfw5F18Y2faE24HwlnEJLjxN2ZRTF8yg8w1wpsUtyldtf9A8
EThtLfYYCYkIWiCRKtg/Asr1Zm5FhaH5zJ9M2htLod/Of9KPSoxooYqiIschRogR
Z3hU08D4+jRkeM213GY5pgkipagxPJwtTQPFI1SZLYALd6sZBEypWOKZPsthDllB
Sh2u/b5zat++YQggxPbLpryOAg3CgK3GN9ewAei+dNjlapvkNbCYjsivQuQ0yJzz
1DKYs5ESNrwy1fAAOZZFSmGhbU/2nQuZjtyLK5mnlKAsAM+gcb8PLSAbdWPHBRXT
SJnCjUuZ4A34dOyCeGpMIJIpf7pwnHMF9FAM2/9lslZdtsNMc9lZ4+y97i6bvl5p
s8LJFUHq6wVM+VBTelrbKJnLeOiEkp7Icmf/nxQiPsLtPf2q3ldgqjUPML4GWaMv
/AXGokEQIbOuAUFDDM99iaCNSfKN8fxKQ94um5rw1GLwq4cIr9jxUCZhysC30f7d
520JIBHAwusfaavJig1dFyI/bYS/wg5CEFM0tGiiyvUKNp+fCXN3iRaAF13qCcuK
P4t08to1Yqq+7Bj7fk+/BGikludSbaiz9GLAQmF4eaCwHRAkzhfn/6TkeyTI2uaT
zPGzvZOGKR0e9WwokwWqLCWMZmzoskYfMWw9a+MMGKcYbc7TQ7sC5BknIHvByL6y
N/yoEZNOoINcFM9CoBbIDWoXQY5YVjGj72gGRJN72sjn6tO+kAkq3jOLZKOauzyi
0X5CmwnsYKsnEbIAxgV8vPjFSiY/RMY8vMMJ2GWytfkC7wRTQ0sLcKYkh7B0a9KD
TozjW5wjq+y6pP1LiDJNQr6ezn9U3FBEryouUeLdcOT0UHLFo2VVFvLnBaIOH1Jy
KZbek1ZKFsXP/K0T1LylGBz/KekTj64ZwuVZbrw8OtRXTNBGteSI2Hkg2ppmJuYJ
VNffaO5+rZzyVZtzzIwnnopKCuPOfER5ag5jaNWl7xD5/HsfBwTOPws5BZ0n/9/H
gcHPS21kTrl4oX6aTLYC0TkCt5hBLsfXvOBplQ7iQV081ZoQDUZ7o1Cyx/hTa8TW
ah3KQgLDthtTauukBnukMBshTCkW6HlM0z1RAL9r2OXMDN/NfhRpRN0YZwwaLHhg
Zc4XKbbtnttAlLC1kCSKvCYm3ySFB0rexJuqd2o4TgCmYh2ykc0vWD7ANCuE2OHP
hTNKzz4PpR2jYU3KI8N075E5G24SlDlvWcY+L+t6PxrKg9Gl62ThJ7t5UgBLyqxL
s/33LFpk7dy4JwQqmQsVhCAQuL7bmRm3UrRFNLFrz9uw2jVB7S791rCPzSTJzKX4
XN6VTM1jE4Kwn+BpfW2zPA6ppecj+nbQzqHC74shTsy8JLv90z1uEwTlgFIG43Yf
rNQr2hHo37ALOjebkcKz2/EFCNQ7MiVK8DOeNFeZl4jn2iBgTSHHv3OJiCjRbtSj
vYVun1oOOOF2j/ioWJlf/MUnh+JOcpL4YWi4GcJhFTvU2+h8qAm0iLdjLhA8EkAH
Ph8Cgpd4BIbEMGy7am5yYfcGCFFHBXreg1SEc3hwN+txZBezLZB/8/9ciQvyFMrF
8YsNt7ZDBMN4obTFxarOXuPdrsbBJDx/9oiQrK49ygb2Ll3TkZtmONe8oLmDSDGR
37O+X7qoLO0lz37Hb3RU9nvQJO7OJhDeASEAhyCpAAZvUX0fj9E35bsgFnjVWrqH
KZz2+LryqCp2h/LOXtD6KsDWB3LXSJpiSXxYLT2Bq7zYrpiB4ra4qm62zmtheIRv
rady/kA0oWaHVQoXio+xUaXHNtNX/Pg6fJCfb7U6NMU76xgBM+oQA0ZTSk390dXb
wng61PV2YRSQYCCd/nStf4MBixYMGHOoxSlnxPM8kRDjHa2s/bOHRbqp0w24lX73
KJFu2cYvSAKk3CnkJKoWwT8zslnYjyn6tI/MR4WfRbUEbUFPGsPJ09Guj08SAW/g
DsP2OesbSBjS4tNGZ1GM1X9afsiHPis56CRI016l7L2lOfCsbGxXuRp5GTP00Erf
EYfMMivXN55aEiPH5WIifqc7Qa+4HrZF5Qe8A1eGU/O0/nYJqOFzEUDGlyPiRPN6
ZmfIiQe20+PK64ovnbUmPsHvkLPBKio2L0WFlnu4qjOgLNOjoywNnhrtiEy9Q3U3
nTFle4TsFkxQNyslnin36X6xJBTJvhCWQS6n95ovwt0x/8Sn0jLXowAvDAsasHVm
0kqZXC4DjyxzLVjt4OP++XDbNrGs7YPVYcmEtiMkOKUCCJagtYtMPED30lakbQrR
2eIGXUoUcmxSCaD4FvITVfFgy5geIR3MDtx+FZcxaoJVjbxJvUNqIYtr59lFSUCu
FlY0I549Jm41xPhkCXyS5dwOCG0P1zs59SmrzibFC8IaLSvqjK9Zz3BT7smT04KX
mA7caTYzVTcvNROSuEvQ3BK7I/Z9RaSFSkjAAFnBm3TZLXJfZBQfm+JvFo21G+5X
yFgF/ookrMtQVufVIQWFVKQDb5xDCgeS/7UeYJGxv2rH0cU43hQfmYJyhUxj9aFq
P40nX8p1DGqLGQLtdDj9CtGRVJ9gjXYZJCZNk5JGB+QRrpyRdRxToqnh6mSp+ogy
YjXr9ScqPfngreI0biIKBqzr1Luyuy6EpR6c98edBNagND2FTBUcfy9cILjS/kXv
yhBKIN7jOxgVFVoTWqaRxFcubv+d80GW8wWVbYir/Y527/pPwwKmDDYJfP4kmGuu
TdfizpJWaOrUhy0HgkKsqhWFD0hDGh+eTOlUHg/piVtI1vRC/Aa8TV88K+tO/Kcl
5m1RK2attoUCwZUOqpqUn585n1REoRSIkq8kZGR8Y+jVI4f8hj7s4+EZ/HtyPk0a
EjIkmbRod2kNe0wpikfmHrHzmk2xOxGsYtvIpZpLo5U2VlUztKuG97VzcjNi9oBr
qEGN1RLKXPxQUEmGw5x1ysDhZDwckmDtfZeh9pVrsJHo95keNo4cYzl+NMP7ktKc
mKvOgrFa0S7pOGSyOrs0iGUk0x9enQQLtzgfKwDjBcsG0zrBO06OkxsTQ1Rw68Oi
TCdpqGYZNCx51tV+M5NyEzEx3iZ1H/ztqfD+J970rd54NiflTN+X62fam/NoB68h
g3BKZ6+PG31J2Y5+90U9IGflJGyPLrSH/yitFZ1BNvqRM5/wxkxpHuTWRM9a0EWw
Tth6A2Cml6B5L183C6th2hhGRE+n+cN1MoO6uvJTv/mvBODzGhd+T5R4ekxCt614
n5O4GqcAfnm7NvKT26vSW08zBk8/+7tq6aMU0uH6OlriH4/69cglfeBVfx4Ac6F+
dh0Nu4N5xwZ1q00Mp5oNBLA5LU+UpbXj0wkEUlgqpHhAcUy98gWCdbUz2L8sDBLQ
kof3m5W8CJitWdjwYHK7j6HWP3yL5tRl43ZP76w0jo3N0w0zmUphe0zq7K+UJRBR
ZY6JVBYGiYEzmP3y6Cj8KqHHJukz1ntAw8/RbJTIfDtp2EdTP/vlDyVBjJY/qxR3
P9jee9oqawkKEcE1j5k3bnb3v3AjS6tWp+ktwkbbC5WRrqsJ5MfbljaSwJN8IHpw
KCZo0qSwEfyTy+SNN1pMgJCgKp/+BwwTBb73RHddK0brW+SFjc/nHgE0ahallH6c
s1ShLPvrgVuOtBUHxLnkxSSLXtmSPDAd6Xd7nDyxfMIe/TcohE74Rr0Nsn7QVH7u
KUv25zWPEQK3hescu2FOmwR2GMOjMsRcK3UCIdMrHpTS+MbxtHhRv0Seb4HZFWVV
P0vdVurQv1jjz88/3hhgHv7WP7qMr6/sgEW5cx5s/Kk5AfQ+CsZKUX5ISI68lvYh
gnryLLldNfcgDM28jzAgT8fOJJ3CsG6PPRTXQiiGGBfsAmQScB/b9nAQCe7hPvGv
pz58dLxWNHwpuxa9AGHC1pIYuOV7b8KPbniw0c+QKKHqpCDpRoKaEqXj5vVDUC9c
WCMtPc9/eYL5+1FpoaBDp94+Kz9DL7+wvpBXMOfKXvnOJUdrWWW58XdLzGKuwOIC
Shstt5zqxT0tp3b25A1JxE1GaOKWsMJDE7FLX8qc9miA/vpV4M+g0edfBJCp5K90
ixeFm6yXnrenrhPU5iPr86R4mprIpVSL52H+uB8OHoWugvxViLOk2N+UVD2532vu
`protect END_PROTECTED
