`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjyAyNbMav66ONc8e3t97bvKY0d6iKmjLYk4we8aA6pqYztbYves9zW7i3GV+2jK
MO/mX//T+MJ+uC1a/qIiSoc4gPOjvLvs6/U6Nz/DNHDDhgqYfcX+2YsPcEW72V3/
8i52ysM1ltaO23x3+vCulrdMpOQP2lI/x2sGP7fhxgj8ar1cupb80Isxu/48NF6/
vbdhxgHEELA/581QUfgwr/z6DnCpzE+PLUc1XsqKSDM3DteivIEuL3mAIVZQG+//
Qkfbt/5ZXa8JGabKfLkO9daxmptslKgdoL35jfgT4LdobCqNtDhysf0xG1ym5/LU
0g9GUfXicZWsEbF5NZqveNqHoTuJQz550LHkZkuXNBLpiid7lZwdZMKWFK93vpnO
iTYYQcSsIxqNWEuLIYLkzI1sy8BdNUbrdM6Zu6Ru6b4WNgYW822+GY5I8sphF+IL
4oWj4dLWI2COOoSw9b5zHXpyHhF3IIqzcG6m3yJI1n1Co13UyCQ4yePrXoWEAme3
Ph+z5PbCn3/lPWlDdXLvhzPX3UdOGZ4L0sGDq52kFbf3NIi3X4u5qwJGXC20V+ch
PxYZZOEu9M5/zOw/i2DbvWVVkQSnaxLbnoVfBXhiPO+lp+Np3RIJVoJDTON2S4SL
Nav1rPl1oCDAodFOOtZovI6RPBMNQzrspTl0HzFkRevzqZxKOa43s8hfaNLskvnk
3Z3WFajpTpfHBZgyYHFQ1N0GN8fnL4ut8ygNXCUppWtqxNDWHgVVXcXqVZoa7qz8
NGFpQEoxcGLJKcjz81vNybSfZDFwuOAR7iaNL4LeiN3lz65GgrEBCIoCsgRR0D8z
WQRJBf3mGYrg75f4oL7fFlFyegvAwwU+u6sje97Cqwa9DAQIV4Jk1xyn3LhSCKWR
aDV7UhJiUJl38VvWvSe3UHP/tKkYp54vRLrOVL2haoQOIv4dPXt8DQQWPNuAg7eo
odYtkJYoYs6zweP5Ig8MsKX+pqDUwikEDcutVu11N53L1+42iwGef9LYm3QM1KTM
fcKhiufx4dACcWYcenF/M9pcJh7JPXxDkfmS26nL21mozje0oODOGduFZCx7v5s+
NwQKROUo+d0nNNWrkQ7poWUeSq0rqzBPGtpmnT/JLm2dr68XHskdnWAQ1teT16gB
b/tMk1+QTdcg62EMCixp4iWbT9AP9gt6HHBoZjAYg4XfaX1LF3uMJ6P1Gs9uChmo
Kp2PY9k/fX3braIoU5tNWqUZkQLft8FdnHaDwTqHdxgZiWx5gkWJRi1/MI6zkEqR
FUdrLY+OxlHB6JyYnYwxwp6soTNWA2kwAxYO/nA5E5H3fr4Qb/5nHci7g3ozRWRJ
NC+C7PBYU0ro7UlPottT+uOgMEs5zVwHLH9ExOUBsmv6tGqsTowvVCBWAeeMjysJ
b7ppRt4mcJJJVxLp1EUJBUyTSvBw6gOvMV4cDX5TJow+RY6AwKUGDr6DoK5p/tCp
rIkdal7tGxtrNFTyEjDunQZ5Ql+fPnbJeDs50ZTjha6xZbL2cQjVFh1rS09n1I3f
b+EDtLvyjYUSO+A+Nwbeg+jlFrALpZ+wgXrHGCu+sXjd2Chw93tUGQFWraKACBgG
JwUQd22Sde6uWuZ0+iQ/fMIk+xCW4afTNMMx9ZGDaTVjem9S1Q4oWK7WEblCRF0k
6itVvU86zgq1dAe6DTnDLTFkgdQSCuACxvsiJIWXlogna402+SsaCLQoUSSbNH7t
RB/w9XBky2VSCe8x4qBYyvO7wBxw1+Ohwz7zgJGmOlNRug71ewpu+kLqewNZXkkN
eA0yDu0BR18bd5h8RLvYYW/QDSpzm1oxQ2GgONDA/MAkgrq3Jj5HV2GkdsCC5qVN
dE3GiTqkGJg/erFrrftFUuSywdxK8r6AzsiVAbo0b7uPYijFuux6xWxkj1HvwR9t
J8KCpkaEkSqqRZN0hjMIcw==
`protect END_PROTECTED
