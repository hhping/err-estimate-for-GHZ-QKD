`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lpsjQ0eovD6Jzi3tPgJY2L/cI7s4d7aveboUkKzYAUfKRQTo0vojlfzyQ0KmjSuK
UUb8X3eWoWEa5ZTCGzmgs/g21zjzp4eTXzsj0PU2u0N8Hjl5U0Kc0tx0P++O2eD5
uUN68MtxnmyQGP+Rh2TbvKWmfmIPoUEl49uxdL2QwVblpoZDROaaOpAKTvzu0qBO
aQA+1xAghAJJhcpDxvgZv3IM099wbTPSbzHNHMibrWxHBr38lCKCXMVzR3r0OMJ6
nIm1buSmMQUwLBCdTrAp2lVgeAppzIWHXfklP01yojmBFw/AlVD54O9pvKNY3gTK
fEb8pEhFm8GOn6TRw3KlL85JD1qZ3OqskqbUEWtYiWopE6XeC2qpJNd2za4V/mL7
3QpfbUV0Z9155P4ZVQpVgaSgQuhDm0MfsDVsVIIyU9jeVHtnJryQzLsD0m3suV4e
Z9J8yZs+GQMaQXkMd8fMxcIC7AlcVpyHriHAvt8IMMFEk2p4wHqCrd1jO3xBNb5v
lgAbpPqqP1b9K0ohYysDy5CaWdWmILYq+Gneey+zWWE=
`protect END_PROTECTED
