`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Tt44tQo8zNUHunUxuoJy1L3M7hsMJ/JmiDsRoYLT5+n9QEXU47m3U/zBzEESjbJ
UsDBuubJllfXziqRE2yNG0TJ33D+3Px8/VGRV09U4auj16EitLX1taE789rYGwT/
+MDGbYLIB4UYU2M3mjvd4rXFADNzzKJtrb0NrOaL5baasWjfGbfl9BOhPxT+KB7v
aCBbw4nWXmbM0gfLk7isQR6+QYDC+4MhU6ClooBca3jj2ffQDczDQySvUiLxFDbd
GizGnb8FbS9MuD9+i5ehU07j1Jz01rlk/MmZYzffAU6yDrJatStpFsLTGU00+kzt
mN7LeNYTdzzPeEhUzZXXzuWqZOQ6yJdYNR5s+f1/mZukQytZ/BR7JIDFDYo9gi6U
bhCSgJGYYGnZYINAb6Tn36PHEX1dV/woN8/aSdOaksyAAFL/wiEa/MUtB4zJDBcm
OotrU0VScVir4Uv1VYMcACtMZTesfGW/+ryP/CVsT0wM9Lm9BxgeUXXnl4xnTCjD
AkAvr2rhYoxEh7NhJEluDZuUcoBSVHoFqL/3Vjy87pVLhLLcnVqzeNkxbKu8KEJY
OiRqQQVlAU4jjqZj7fgDM7XoE9FRcfIeJ2txeo6qjau0JOk1gbcchfDMUgmhP0xj
oLV4SDF+DmJ8bQIlmEW51oUFE1EQ0r3sFzPPC4bRDP5wSEGsJMmEl27VZLPykv/I
/SM50VnkhkkyFMSVM9SI+TteKy+z+jib6d23lt9dqAUcI2tGj2oA7d+kWk4kD2JK
5NBIRlifNbFHYzXMZCmuLVEmGG96rPWMXKyl8OiWl08uXO2liRKY0TwigXOwRbZw
gu3BigO5C0SyuE6nIFdPtmsYvLmHKLXZJohpek9WB5sw97hiAipz06rmxj4wRN61
vYORwhqE9TEVqBixR5SMeC4MASFLFuZhL8T4A3gqbM+l3pO6hkuIZjXDmGKXCgXc
IEUcyyWMyCd8cCYt0whasbTvQT67tpsd+10WxOapcIwDIEIVYNTERFLphyYJVenI
YtKJPUURniKb3IANYI09RUcHDP9Rphh6+uE+6sZ76mEi5+A40tc5fwbpBsyFKQqD
ilO+lAN1WNI4uznEfW6zln+hqiJzDXu4X3L8hCAr0pQ56dPEzJpyYH1uJMST15LH
BA0XPR5VJ8Vq2NU0EG5wUB3ct8bflhEyrXEDmpEunwlIcbA49TMG7+sKZLQVWDgb
4pwDm3hY1/WrfRQ7NglD8vByhnAGKTlF3ufsbrM++v5MEukOJGJUUTgVYd8koVcb
+uRfZWdqrI8xPhoRZVcIY21ubDY3+XFZfXNLwsSa64ilv3ZCxt0asMnXkw6zv3Dh
wYnue23/imK2rBwRU1/3KQ4qGTRwrBHDHZeSyUlURCyJqxoFYWHsG/6+yB3JkuKF
FmivYb0KP409vmBpgAmT1t24/06zsHQbV38hkqkmU0uWBGn+4MQxHYIjY66ofz9d
QEzLyeQR/Iz3eF+tCulopDMwNmpbmkojjpQjgrOGXAJFoB1ZcgZCBZOC9BTkycwD
WE2r3/7HyjgnGbg16pkVp3OlrXZXPFkuR+Z1iOzGtQG25df3oSaptZjrjaNZyKhT
rDxBgMXi9dwsogEcLzQNd8OMMAX5RsmzeEOeGtaO/ibvDUUoY2JLv58rvugYfBcW
TlUF6ND5uPr4cuqb419fOhbPKeefhuRB8n4UiJUBKui3iNFmWOBFnFMofHD9ZHsW
hP8cO02yDR1p9nZspLrj/m22zPZ+Vsh4DBn6WdaCj52uMm9vcGCsuWz5/xv5jZjk
WnZUYagz8006lzz+//hxuUT44JiiHP3HTxlwbytIbhhnJ73TXDFL994E9ZXy8+6/
ZR1iv6WulZ8aPGrXxgAL0p3WWKgidmtEzQVmKclpdOHEBehMrdi1Is0lmsgfZk1J
KgyEqJWr2FuI2zfAmYzY2Z8ZZOFBiPMLhxHmtG+9uJfWqe0UPkpdYcloz6BXOzhF
KHZlCG4ygI1rBebLhfREJzOTSfVp8kpn6lqjxooGMjPAcIT30R4d/2QyXJEO/3Oc
j4DXjbhs52PXZwEngzqN1E8fYG5N11G+m0p7YMKsI5Jiq/KkuE7iYNPrRW/x/4dJ
`protect END_PROTECTED
