`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OEfg3OwlJmUJjFSvQcPX8dklmv4/Zg0BEcHyErlZcn9e/78/8Zn80PY71yDYTzx
KucBNB8jgsXyxPHvaJEqu3SB4BnJ1ILqnC5Ca0Cca1Ek4jEvWSN5zBZkx6uEGPaK
5Uv6X0qNN/ZvmQf9lNcQTALXT5+dpQJapRCYSFRTQP3NXEvLGlxvS4hPibYCtZTK
WeglKgF2SlzWe5gbuCcpD+v1G55G5T/F6jWHRNxzSBWOIZ14EODyr6Wh3hXcCQGJ
DvKcSSLhi8TVFYnDPa4Pkd9c2qfbecyei5Ju3aCX2AH+/6F8HWjgwg7z836d0WZS
LdLphKVe9por0yjt2bP/yUL8jamQCiO8KCQCVvIpZf18beQZo2m7DCbhJUZsu75E
itxrJ07npyHZDNth/77lKceVvRr8KPK2VYlfIAvOmi9amsqRa7TqCOFsoGPX4aT4
JGiAoAih3VaaHKPr9grdSfH/qS6xbt37CsMToVv+dmxmYoc3UN7PkcgR3mCzI/xP
n2g2irg7Wft7pckLAbWoCE2qz2u6aDjT6OeFtH2Lp9BJMg+arnrJHR5Qg8FnWlzy
0JHBRMN/vxwmzuMHVeY8DDbOoZLrqlNP+h7uwLglS8d+DBbg3puZksJsKISGISd3
NPM7kySxm8EdnVMNfI+SULSUrHF+vitoKaP3DVLPTICE/wCPfTL2I94NU17+rYGe
YTfq4zjoi3jxPNLf2FP3+jCS8XRuYZQ8/xfTyCflFsMUZ5AeIfy/0GQAu2GNAPUn
1FUi5u9IC6tR1/VUzBCkbxLI3T9okpmwKrrstCZxjH/hYTdsGK6Wa22E0B6nVbbw
JPeQ6/aHmauAg1SM8rBVf82RJJckUnW6uuPbmbE+lw7DTGsSPx26fTcgHQ1ohtj1
UJyndm9KcE44DvViP9FaeGYmrn//lXo+T8zRX9Dyt5tE0GwgxgYN+AmZm0INchQr
0+dT+pkuXdUlrma2gsgUG3xyx792q/yVxKrQFcdsyTphw29l5crIgq5bGsvCS15Y
+F98BvJDRCO4rOKsHTgLltJTjbWora5mb96NnQUTelSGMcquOKw5d0VWu/+ZkiuN
1GXMFp84c20en70Q/YBshJwf0W5OUBbwp1P7U57VgPUjFoOpxH2SsRa6uy09t/YR
/ymXXMB4cK7oIKI2ec2RZnwkj8dU6/Ms7rBOUg7AiS6bvBat4/LUIcY3sTeK6kwD
ZuN1gF6Lqpo3HW9fgRYldXvuN3yX0N2vRn9KfNx0jSQInYnUSd+nASEET9E8nYIF
Ihwbgokj5r5nrYSnT6ViiveS7YcCAf6LR12AZkqy7Evdvuw3aiI8YUvIvL3tDiNC
fuh/50Ysq5TsiX7bv2/+tlPAPJEd8ouCyAXiHkADNj/jdKFa3ZYbPtrmNmPRT82T
jijcQPbp/+bx9m6dm9JChsvkS97RetZM2k/5KOFlaBZr64vSDsDF/oNl0jdVvin5
OFSGR7KggnCEBFIKvevU3Bzay1eNqx7aFVGFOjnV7FlhnNmMVbueQgkX75uwcoqd
TOCYJttVMfYrv37/rNWmPZ0MXnHNBse4l3VCZnxQh1pClkI2Pi4GRqL6qT17hccD
NZ5q8+TcKwrvIP+FzJJm84hCW/9Oh81D274cd4s5LoyuKjpTGvBCtGbm73WKA5dr
rxeumeOcVIcRrCNWKzBIxKCr3Ijgg9c4NzN57oYxTi9qwLKAbjsPGxjo6UKbu5nP
lDUSw3ytaQaWJk8vveyqAG2hMUeHFaHNqgycUJLGFgS7eroohG1jYMLwV+w64ZnM
4O81BTga2SO9w9knaD+yOKD+kBfmHtyXRrleUppwYGALT+Ebq4io8ZU2tz9OwS6F
uYbkp+C6lpQLYu6TaWr/hFxrV1Z3VKMT9VwL4REshrgOaImIQRMDR+05ycVZ1tV8
ViPSlPfbYL6WsUsLWSHKyDEqatG4kl69CFIB3uC0hBQsy7MZccylNUd8PHnsuxR9
q5BceaJ48Ub1arrKbYvPP6IojiS4XWf0MNIFkxd3xEv8fqELqbhRdXo1sSt/Smw+
D8b4hjNFH7I+zyIkaaB2aDG6Jp7TizHnb2Vbhk/6PDfWtz61aJ/rGIdiVrhQVKnk
clSHS+BOHfgCCzXKlNSOF4jyZEfTHROu3PD4Szxg9mTgN9JN2eA9kmKl1KblNSoW
2IxFGa0l7rSNkJVNeiluZOfJPAca7Gm5QOWcmjbaO8rV+N9UX5IrF0fz8/xEBzBe
eQJIgPLl4Es1Ie90568yzxLeJmty+ZSCbRR/b95LE3pMzn6yaxe8l9rdOYO2gJOw
K0NMJ9fidAzFxvvmP2mUnLPMPvzpMYVQLhrsPZtSLRQXrWCgLkWv8iT6imO43Aq8
H42zHbWJynx89g4jOsEhaLdsZAmeN1mSlcOqxv0httfBhHIySiDM36mZhoZRVkPP
ketv9KTbailzv5ETgDBrqvrmHdw4zmdC1iZs9fB84SMNXeHFJR/w4VwtUbm5xQWA
wmvE54QhQxkojOBAMjzd5DE6zMcpPl6i+tfuZ8695FjGvTQncngVtFwcSVsUlEbK
NlG0VfR++mSyBiK+PiA2FFPqy4YocLqP8zBKVVPKws1G9vTfZPstMCd766BZju/E
mKgU6Z3kx9n/xuNxP3qNZTgqPyGIEJ9p3qeR80abMTzP1jguxH0UVnI/Zlh0+QNY
/UcdiA6cc6I2lFcwb1o5e8gxHKIp8zww58+b8IlyNjjbxzJVx6F9MaVw/wo8rdyN
5C+hm0Zl/EBCQeZCFpoRQr4v0B/usyTrnQS9s+88SpZxGwwLkQNXSlQRjjlx9/pz
YvcpRGvhzconvkzt4DrK/aCNXqLz5bqragiIm7AXHCUn4Iy4AwIfCrb3Oi5AlGHp
S0f/g/gKLOfPKulAzrO81r2TRpPrJEVSRrwGMgPSieVvka+N3SJ0ChVae9tfzyLw
zuP1QffQ58/8woRIUP4zLf4b+S9ttFLZ1k47bKDXwbm+BOiPs2Hs40pRgmEGNDIU
u+tlUQt2CvBVSXfqymToNbCDlq04splgBKIMT8ePtAThPUD1+tNWLVJ/B9U+zLuA
aUecP8eXXFQuN2tunDOJXygZ95BTbzwsnt0KGVc5WP5NzkWxhfKmEV3zAxxQw+6P
dkyh2xEknnRXmX/vq8i4aUo6HB043zW1+1jbtqZqiWEU/Da7JRAwW07Dr/6pGo3/
F5Qtx56JvvwRdZ7Vu1yVMXRvYtY3BAXXSSheVWl6Oy8dvRy7NwgwwriGGCUSJKxp
HOhI5X/tjtig5UKwvAOHQaxzvmNGgZS6b+h5oJ1JoRLYOnwR1T646oSt+MoQzKoL
aYDwOBg3VBD5y6OAJJi+PfLa2CvJLnUcegXlJBR6K/06Tknteeo1tdShOOFFvtIT
cdaroAzAZZ3WSfdkayi48K8y/nzTE61Meo0Z/SCRsRG8gjjAzuA7Yjaqlfsr5iZT
7v4YhBR1wnWZx408bG39RkOS5onjJYoVB/SgyXrGbvTi1Y+YsJjQHg/h5kbcpT48
eUZbjxBS2p+hRxPEJPsePsFNk9V95XsMLGZ2XGlDJF5G1+NMRt3up3YDZV2xJVKg
ph7hfyL9CXKhR1qjPlCeVIOxiWGSqkB0//5H8brYn/jJlPGihmknZqw7KKvzDjyg
Rr1FpTsSoArrRU6bcBjNASvqeTW9Nr15bfjSD2lO9vLCN6+ZGJ1CoU0mPHhyG145
eEPDzy7CBimqtKl32aklp+YbPkymDLddM/EXi2PD70oWu4t31dRr9yPp4IbxQhzY
rIp3a/X0aK5ZSNjm+ITSSS8r1BVHDPmyXfh5bndJncr7sW1GtwBdd76kTse6LQui
AvvQRuiNhDg/7f9dn3VZtbHrgiGfyzrWJh8R6lrk0CZVUknjg/lYXtcZawpEtvsU
eZk+i4TEIYcUrH3XEcHk/HVDUmhIk3bj+1ZCeSc7wvEy+Vjwy1b2eF9GeYHgdKcE
2aREF16nIiiWdwqEJKBhncBONqIVn203lzwMFoE3C2fpLSGfCjcTYosbogu9fmSy
cP4W79REi5MqZ6dSxKUJrrRIa82m4ZqIgr5Xs2FMYoX7E+cMX89nlCDF1wWfwZ9C
Z8zBKCR+F9id0NU/UAkQsgR+iFFNDE5pyAGqpCvXiRJ6cl1RVd8Oyyz4scYXvgCx
zEWXZvBxGPxmjvE9ce3LQktNrnIX6DlbaWkmaE819nxWzjSCy7enDfwFV4HyUKe+
7qhN/yYTay0GtSEWCf/H3xqC4OmxByO+Wzttuguat2yArv/QS78KYHrvndVIiXc1
0yvBRZaP3F7cC1dK8qWlG1bFz/dIhq7Oz/YyzOkiyCtFrMz/YOAxP0SbqVqDQoyF
/jphpPys+//ExWVSOiWFTwBV5ApPzdLsDxYWxjsxd9HTn74lGpC1PX01pPHiA0ms
hI50psVP9oJuaXgJqdr8IQ10Bj89+nSR+oVq+2RxTesj7JJsDfhOP3PO2V/DMjnd
hV9k2R33LhOeTJEoG9R6XcZDqfeklSKY2KuaJPZw5rp958uePlC4XDnJ6WZmqKjb
1XnUxK1GhBVoQTLYn7Xg77EiAAoas02x4RGUYtgbj8M=
`protect END_PROTECTED
