`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eeNfdMHv+RHjq+LflbtJxnjOu7Ijz7CF5HJoNpelAZpTLoWFuKnVM9gi2NvoEtZF
IzfD0pzzFC674QYPu+m3vjW5Y9/uQBaWfcMmLVt5FfJhZNRSY1sYgxOwbrl2h29s
7SkiW24LG3RLkxoTObpGXpaOBJ5yP5u/LJ99UYb8tQMmLP+L/SYE/azY3IZSt8VS
KgQ976iPf2Y9qwTZainmLIQQ7vJs1jz1Ba0sdKKF7DzyawFDokUhkgBteW/mFkuk
8zXsU6MjYsYvL7lMHHX8qreXiDzbMgDvHxWonS2hPAQb5L37SiKaeiJwH1WI40sm
q16zl8C6SJkx65vkmhGH497wUynqcOoRSYkzxmxkgrK2pgZ5lPtwmVkMHziwh0/8
gEsrPDJYJnAz2QlgVVyIzkF00zwdTIKws22zotLcoGjH8sEQne7vdYFeES1vPJOQ
ZysVXHfXGdQctVi3DLUobEOBrk4L/KsL3bq2LO5URsldVJaMKysTlL4AMjL/MNg8
VAevcQ/w9p/zOHVDBN7lINmduZsuUCKuMS2yYre4FKw0uEOvw+/YyJ/mtsppcqet
NkGNr8GhRcwRNvGsVG1m/yMra04RCzRSUrkrffcLhUOscPoJnpHgAtkj9yLnia4L
Q2Pr1/FkpPhWanbzdSkvFKYTcPFDBdMc/sURnCVAuzyxUDlrF9UsJ1fcdT1NurHE
MmyPcJ6wxvNTHLFjUqLSqxfaUjrlEUm1zle0t3Gs+JrGhJitKpxueWWrF0BjQimP
qyQHy92F3O9PmxXhGy7IMxcY0AvnrOW6cyaerhfNfJhYCe5UfLsB3kdl4gr9QlTp
T/aKn1mb/jo4YjAp3mjzchTCNRGtUJ/Kw5mAaa+zFxP1f2M7wlvfpz/3fgkcsYLg
gB4M6+HJHVbtxWdcL40gZ1dXP3NsACm79L6t+Pza9ElJngO6O4T0FLNAqVRY8NKu
9hbApxemxGnpEJHn68mhKPMQglbV+vWuNFRZgZWHkKoUwp2EvTAAsgo73zrCrh5J
MRfJXoasoY2sGnv+orXLxgj9ITZsNBS01Bp2aJ7cCIPXFQ/lrRbVeVzI6lbbOECX
KygnYwzOhpZxUbvvkqbLsaq/Ba/U1smPc3ZQ45sqtvYaEe+MU/OEdCVqbp/r1QCb
bow4K7WT/+P1K+7sN/IO6mmVmD09p63y+nzK1RtNL2TqVyAKEJpcjPo+nWW/g7Ju
lIz7SB8dDJ1OltWdu2NEmW8K2WXU7G0v7LrclM2soIZDgTuhlhnZcY6XKLSEXluo
1lipu/3+5R3WCh5rmERAOw==
`protect END_PROTECTED
