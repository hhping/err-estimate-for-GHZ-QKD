`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OdZolyLIzhtU6Hnzu3K9XiRRD+nfz865VChJeVSm99arpsyGOuVpK0HX+n0Q5kgM
vrQzgTdojYh69Up7D9OCb9/XFOKWdm2thm5tsRZRljew/GQWupY3Ke+D3D5re+KY
C/0B1DEG9Yd+TwMQTArPn9qIQ7yimO03/0bw3R7jeQmcLANUZ9hjjYT0VGFa4dmS
ZWULW2AqL8DlbE404HkPijwnD6yk6BGBMkeDHH0Yjt/PR60D68S7EzIBT64Paobe
PYOU25xcaUJcxQy00qatqyvLaEXldRcs999pEuXE0wNaCEsbO+QYxIZbml6Udkth
pqVR8eLCmnMY2D948bWZ+xXNlW8GUNEYBolkGAKpPZ0evAtu2iXcsktlpsz+EnBX
Npszu8I3YzUSRKCD12ERfo/AVfutsRjQR42n6olA4D9sCPU2vROwHYSGmPmR6nEN
EWG1dAlX0gi9Hi2hHbBwD0rFAuvjsV0Et4lTw7ErG3+Bbs58GEKGIVdmzrCJgwvA
4KpJNsouGs5NNtcmmy/QVk2oQl7kWRJW196//AIuaUWJy4f1KtSz0BC5MPbsKfa0
khPQvF9nuwJogtn4CbZlHip5TTll+Fr8sJ4lqsnIN3FMJlTjva5uF03vbICuj4aA
ITDG4l3nmUK41yI2Pg+2vp3jrFVXvlfUgetpjTlu5kfxnYgrWQE7koWQbNl16dJQ
K9hazQcZAF+VI3hk7negitClF7TkFpQ6FgoKwNGWg7ebWMzOYh7pbqhiGq+UC8Yw
nFg02aI06EmB/Galb6TsqTsBkotc8fdIdnIwzeU5iV6/Bx9ValDEzOutLqcIdcyi
lOBgHumnrs00HnePJjTbM3gzFGdxUCaW9gBKH0bXsMxkVhs3zsEZYL6B4GbkogkZ
EXze5IAkHCCKxGAjMHtNyw9olm7+OjvQ5VoE49auGwfDfylteEUcjVusUmYAGNux
eckxdekiMRPRnub36k8nxX5Ep/MlbAj2mYumYk5Q55jRb0RRlkigLfQN8CUnOd5J
nUX44t/J0f6yxtYwZQf9gadISXi8goeIt7sVz3q0L8gCkrZi/nDMp96UtiG0RZE4
`protect END_PROTECTED
