`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KaxfDqePsXeCvvcMKLmzOOZX5Xqz4c4NYYT4Opk8HlEMH5t2YGBS9yDthmg5mlX
dCr3xqOOeChSlVaNwdrszFj7y8lbTeeYMeLaVtTDQmqRV2JJDDmX/iFDunKQZRyL
viqunZSqVwuuSoW8ihNZ5RYCTfnWxMo8A5x8hEE+G2f9WWKUw6xy5Q89B/53Ue+c
TKcMsvmi5MCK2oThLUDFWiQDEmWd8HZgExn5c8ZjvJLo68cm2dqE/I64ZSKG12SW
cmYEEGOLP1vOgZmKrfwb2fP3+mkv3ERbKJgZaaihPlZ/eqQEdraGIzJ0BL8eEKYl
2/y4wBMam/8VFqhD2Rwtyb+5gN7Y40cqfMK6YcKQ1dwOuhbXIUfTpRnKbVV5Sq4e
40yFVygxaf7elIy1pLJtHtcgbBMsm6pkSLsLAA8lRDQh9r9oW9JD49HMdJlj1KKl
TiSUmaJIc/QG0dMpfX7TeVR4+tQrfdePR75s39LvtDco6aM4+EpMqe4ughEw/+CC
0nqENwkVoACO7F91DFJntmHt+tl6154KdAECWIMGQbnRIWRNmO2RZunxhmMk8/mj
FlqgpidjP1qA54Sfr151KP9gPcSCqccXB1XPUcxfoAP50ewG04gxNs1oPZMjifp4
Y4qzGu5E+qvQu/NX1836d2xRbu/9MLQiaHfwnIMvoChYYecp0sS3fyXmM7dlGmx2
fi/xeTjfbJZ6ASclr8pjE4vHZFDTnwpYPUyQo41nR1c=
`protect END_PROTECTED
