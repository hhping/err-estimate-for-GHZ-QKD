`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7YzIX5s3MPEvUJTKQ/AXhX+ro2mkWT7GBJHvB2ZOMVew+ZFtmSvfOVqZUuSXh2pO
F3Stg6FKkUUr7tL/Q9+pO/StBsF96+1NiNiz/pQOekQMr+xwcG3dLYCaj0a9jRGh
AdVzIUUdxD0WzRwICmA9JvyRp4dB0W+P8CdjuZvq4Aob5a96YVE+/yi2gmjM/ixM
ZoBFrVSf97tcNti1Z8G17RBmv27oPq5UuHngKgfuku2lNu4fZ88rxvQ6IGW9wYey
Loc0tCg3SHkVKWs8gAGiu+mc7ecUWvqWNF28LyqPPcdNMNKmbp4OtCb8lrF6g7yp
sGqTiblQYuuWPpmbh/4dEYC4IERe/2Y85oEYw2fgEFWWWKk8ZtyJiGNBVq9H7xcD
WPBH1BALjboOC8oHb5CjXuBbcvKNkvALt3GqMkp/4Ts5U5FrinoqMWP8NKcFe8T2
9tcU0xXIlOKIR4FBDIYRK8aQEDt1hiQV4xDKXc8Pmkef0C/RSMTx7XWNRRRStvPm
/CaVme8zy4xyKpCazqn8odzPBJZTdFHFGm3kc6v4lsB3/lLwWuAHiYypUf1W0L5V
zMg7hw2IJFmva9o9Pf5bEzNhUJCva/mJBJlFuhVdATlwtBYDU0884zOGEGxaYeb4
MTvhKCJ/w7klOKzdlFnW9sdU/E00CF8JKQRk3TAkp3tLp32Kq/iFLfacoSSXf7Ai
v/O8tDOA7kL8Ggs+jb8bgzUz4aN4/w6q4An7EuA4b+w+1/fUzrXggNdINc1qwiu8
28s+1cyTfbeZDpcczOQEn1XMt2vKtiSQYBcNEpvW0gmaU2siXssACFgKOnuPanb2
Dlg+w357X/9fp3JXQzJb+EeNmQBTBK2lSrXSD+25HmZcqlJ31Cwi/xDPy1yzQDA2
VjME9xTcqdQu80wbkZ3HmNqLvwhA/dlT4bEtp3a2a0yAxGCUXSwPYbfq/tBcL9+c
8rrkki0eJywcvsCWwxI2SEjQ9WpNJmm0YVWypQb6i1GSChBaj3LJp4rSBuq1oato
ZdHaFnoR3WA35WSmWbZhK0f+Pap1hD3wKSuOXdO7FG712J3W5WIyqiWm5Dhs1eIv
dEKAbAgCy+QVp4JY6Z7b8aAa+nGH9qEtfzQj5P2N7h3+9a/U7z0BTH16+mIOv7wR
lIFBVRakbKxsTMjT5BJzRwqK/8EaW0pfGkbk4DLFbSfl7KSqsoxLps3icxEOxWjg
pUVrWVuqQStBezRDBp5UAsTEZkrLwvwOHBO3qdADEdgZH/v/obIMFfiWZMJL4qJb
ITH1MehsNOIprGu2phHLBBUHzTQtofvpsq+zbPuLzDIg32ZHjMYDgJ4PZFp9JmaD
dPXlCjHVIut9oWTJHUE5JHgY0fZnjdEQOM0Pxz2awWmcQhZ02aIuwCSc3IN4Y7W4
F9N5Kh/fg37RyBiDL2Z3LF9GXkAi7KVr9/7+6ZabrQN9WBSL6tNlj5KWsY8+8+UB
w3o6mnG82jTuJX8jhlIxr6KuXUAmvElvBd5Hr/B6sx1pTxTYE2FrYsFVNIBSV53f
fefdjpexy+auN7OrdW+g5gwGu4sU+TQ37Krpgdt0o0yAPqcr+Tk+LYOCKYbSMmcR
eYlOqdxgU7s/P+caiLIl93LL13G+yy68dzeKXwdG8WUbxMHO4vWqYRGV7CKdK5ME
lnZe9XDC6eBYhVBtXdVFQ+0SSXr8dSAknF3yPkjuuoRfR/63E3g/zbzEaWT+SceF
UdzqXFJQTDJ8/XskOgNy3/fiww02chcpeX3jf/FrUereX5o/dOIviE3igIXT03mA
dyU2ZiDbx0elaH/6hQKVGlF7Oag6J4VWApBMFyrpthYIo4uqKwUfJa+liRnDzpiM
f1FAVfbyodL84e6tUtcFCUeub0EgYZQuid8gM9jIHbmKJhoeKesc8jDhL1NOSHrE
xnkx8edlvttjW8LMvk321iqitdva5QHEy4E9DhCtTt25QZR2y3WZYn3pzcNsrFjw
gZVZ3WbzarGlNUgCflZ6zBd1BEMAgCDpXkxDk6horNwlaYkTCm2+uTjaobwj4tz5
DEP6d0DxW/AuxpxZHDVo+NeDdzVBTvHK08qSJ4rYOPNZSN/kVlyhez88VwARGZKw
DMpYXA5HMcRiIReAUdvycTvFDIe2x/blKT4KzglYsKN/BtewfXUzBP7fwAWYTXhB
6wM5toDxobxpaPqpyyaXcti7ugoOGOQLcAk1rkn4SFgiBw5CC91on0hXnryH3a1N
DajGdMg5kucXSwO6wCIjKQcZcVzOg5yKaQyh8FHtoFaR9MrnOZA2xXthMtd7kIjC
YGnzkGK8Kvo+az7whWSqIjrDJHrZWmASIyy1ThLt7I6KTQwjlbCnAecsqPnxkSgl
3+oR//ltJW2i+rFXPaCfS3Gae5vAT3kun5iRhGhWkAMGvCY1wDzG1ZHCwoo/M2of
uWkM1uSa4qO5LsLlKHwF2dvYHFfnAQoajuqVvZnmFBQ66ArR5tRpPOitkrC1yjMj
LL9ZR0ijWU0KLIOVS9Y0a7kl3oeL/QWDdT82WtdCE7U8OHFXO1feNmdG7hk4ae4F
`protect END_PROTECTED
