`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tov+VRYWC4mEhRvt4STXNBmbxDg6+bzGfMtG3zbNOpucwN2p86nbPHK/SoNUcI4B
LN60R9+3AsYMZfcioV2a/k9g1z1fwfp5EJtoK9P3HsJj7diEoHvyOBRTNhTRcXax
owyXNcWL2blxuQI3EXSNu4VEDDTlqtgLyvQmIXhhKd37YBf1Fwb9gMnSE9PiJtgH
XcW9o7phnBnkzDkti2FfImbI+BL4D/s0RyOp10JjbTJMe31z+XCcziGT0kietWWq
sPojgiSjy7Xw6V5jfvCqDQU24dxzY58wC6HxNWhNB+ksatxz0EacF1pY18DG5XoH
C6yG8hHeI+szeQRflqyasF8DunOkQEEoqbEXL3DjQK3V75Thso9yjDAYtJRuX1qF
nwpuT/BQdZJiJjoeNj2fwqvXgsCzuqMwbOgFvmw63OArVn/KSGuio9TzV6YJ6nJ2
u4ISMmbWisLFQwB5pdlg3bMUZWpXAgyB0ypg+R8LBp6ViZy1aV2u5AOfgXN8gazc
icKPQBdd8gzsmghkchXu11dhHtpF6NgLSFZvGNB/LBF7VChBWsKnnSKWRdL5YDff
J9WM9PtagwR9pLpgwoZ4cwVz6XYs4ZKjoMKXCp1EiMKPYRI6qAKplwP9Qn9oEIQc
F959ofB1YdiTZbzeSuGVLLKfYVzA64PXrco42O4ucsQQ/DPJCocmeCf+iZFVe8IV
2scgoWLQI3ef27hw7koMgnPE7FH/LPLd0Hm6McqQB+TQrgapYVhBpGcpxJJT+zau
TEZKfeG+VsSwQzSz7RxskYDg8kK+3OeVqwe6A2HlpPZQgKhc8IK4iqvDnyhriy+Q
CX6CK4JXxYd1xTbHhmiJXcOYfvtIPPwAlGDXMHg3FnXW9Y4io52XacINNgv8eKrL
2uzQZvOUglcgqf6z72WWMEThu9CIMsZwCVlEu4v9riZI1rFIuRNgAQz5c1bvqCza
VA3USi00QFpJZfzsH5XbD/geDl+UxsSVMhMs72CkYRWmJxPW37mVfXzpQo+Vvt/T
HfqYACF8xVLSyFF0QZh4p8Yaxe91FXTqYH/d96ig+qMmFZtdCJ6ffSAYYM747/Px
PGfn9KZ/i6uAwAjzr3hCHQydo3mwTYrIjRPVVInVz+opX7jMNJol1PBgfbiYKMa3
o0dwlOgIXpAgadzG3zagzAEd+pzbUyHhzan4p7j64Hc9t9VzquPCRe+rWRmKgMsJ
Ct9jZu3lMNMT3eoq00X7Re58i13+eFPx0oDtuMu2UOZpIL8JYaRlTDul8faajW0a
3Nkyi1L24qlr95ZouyC2/uVw5AGIcH9TtuXcLos3nk2f8Arqwj8oNIrDAxO91gyA
88tznmdoey3x2G5Xop1Ow5pLXnX3Wh32OTE3sWn69kmz5uzkLfltuhRYEIVMOReO
AYxJt6i82eu+znNmoDlvisNw3LHDrlAgNMKFbaOPQKozsoLt/tPckm/FfhtynwGW
VKmIX/snAGs2MiCfUmUI7TsUdirrhJejjq1oYbVlO8cJSIBvI9AoElSEh3p0ZZ/M
fPjN1dMqjTtYQQ1FVEQwhKu1qNfEa/vviDOi2csAkYPMdOhl87uhb+hpXlYKctA4
aO6fWe9AxRWWz8WxQTVBhEnH/VBjOGNQMMdtuQ0blpH16RKy/LTelX5527ay/uae
H8ZuQ873pZzqsNYKxJ3pfGhFA3jW99Afh1RzhA7FAjpWyZFoCIs7EloelFtd4uUe
rOGHRHYY5cRizbIQ+gFgJN4VmxMyo9y8rFrN+m0hjhsO5CrEmWZQcDOJj1RUffVj
fqN4SnqXWjVUxyoSN8uHQXz3V21xUStMrtjsn8vP0zP0W3E73tnuVakaMxH2YIsX
EfU1pckAzdBxZRdlORiag+Qx+9aR2wexHKo06NxAdrApe69EESd1x5+RHHmD0D+z
Vg+2dLxgTstq4+cfWJWlvDomfvgL7r0bhOUgulxXzI6V+seiUuFP/fipKDYbZSbL
xdTQlnUJWjgJCnrlvHEz7bOqw3zgAWtrfw6yFzCn2rVjumX5aaG2Gn2CMXfkDaDW
hfDkvFDj8VhrVbY6Vgv63mYluOuVzKVhV0yiTCjvO5+W/5xnvtPzAK1YkDPWUFqG
Wzz25XORmzSaTVbDc/FQXdDnjPdfUpOaG5C4BAY5VE1As64HYmqt70qZuUsEvvrJ
NvMWZcjjwSP1Dbqnde1Ep5CIPVE40YP3lFiDGe2FDelXP7CSuc8yXCEC/SIje9UP
Ja2Tj6NR6h1fN+jVoy9fh/YLFD+OqMtWIDS4jVxv+UtLERKNcPRioCS2kV4hblqp
fOazlrDe+EYllCr/S1J4hQqYl9Bd4++TDKKQIsbsk6wA2xLwUuWOFg1+6re2ptLx
dK3HGETc6mznT5BEptsK7w==
`protect END_PROTECTED
