`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ImIwhsjz2fL904Piq+MNKuf+/mzeQueUjC1BH6Nf/mTC75Ip8GoB4UCftuSmROYP
wPfN1NiA+3YjP5oYI1U0NVQen6wRVgna6kzkSWyhkHNNcmJMzOZbOvhY+0wmDgEf
hv+WQEkIU2qhAG0KfA+S1YYTAE9ScBSK7ezfzHpIT6mYiQq4YCFdedlzshc3dvKX
86S/Uwvw/JQ5Rt2qB1F5wkCm9N7N5po2yaa226dlRsCKdcKvqhUdYtrkkvRgeATV
3rjeS1kA9khcDdvMrnNHEFoj8z+XQAaLGl6SG5575FnjqQwe/mm5djT1/U/LSl1c
m+VHzyCjY89UrgLHsb1rjjQjjh7QOIDxfN8v9o+34xWXdP/fohgJRTDiuWPxycYF
RpPYGzthMLoXInJnrqq0SoDM2F//Yj+XkTzXQ1Y58g00vvn4l9w+wBeAnZPNnCCm
s3ftpyhOrU7jybsBr2OWUI0SpsbSbKnmj7rBiX6Imp0KZmhrDSHh8f3oORQ/gezM
d5pdfUcvedVFftyxfJel5VPoO7vkerPOh2avej3CR3tsxwsa3Lhmy9B9XIyb7cwD
M+dqr9v7wZLitNPIQmHYXiMm32K0NOzJ6K4CJZo2FCtMwx2drre2u2tAJMk2Zzdm
1ExaRG61s4zIT6GB2RXLSnqZOS3u9/7NC9IuLohfzvj6v8YRvpM80pigg1OQEAjq
lsW12Nlfmwj0l5NqVy//T235TFBNHA7ZcLwq/HWBAXdiTwLfkTpRJUTqGEgykIdH
eEUxZWiptggJE6ylPBxzZZeRn7WDS3YbJD/AIciCD/kaqb80+/mtCnb2CKQ0ncRs
DcBxWbVActJsVHnTe7BmesuA8l9x3lPJGcAaToCav7yGdSPSeGuQROOKHQ3qGyX0
MxtQupMYF+IGYOWZpL3pqLDerb7Y9wTKUR5uLV6W4RyeZPFwjppsDxHOdeKcLuei
Y8Ml8SqRc7UVuCSt/RRZeB0ZXmit22Pq1P+kxI/MLCfYMbAKT1QbrluQRHVRmw85
lJnohbQDU7TuUqzvmZLk3l+DZkGLnZIaGd7BsLwyxv+wigZZERPgZjMryA0ugk+m
DTc2YgrYuYOi6GSctU237h20KVz9v5Y4dkdi7oZDEOvGTg5uO9F490Wsxx7wf5Wb
uXCRHEnCiv97L2VYZFipiaVUmx2jXMLVN+Uhp4qkqjNNeaQRuuDxJ3oC9tJx4QxJ
Ya3XIP/jPaSoC4HMdFX+IDH6uCHPWwlVIcDuwpiEWaccieZKzcyg4/A9MdJggPWk
BDR+vd82PtuGfAWQupo+pGNQc/83TUgk8YUXXtm+J0CHnYxpL/bj0RnescFRHxKC
robj4TpeVY0ZyXXHoy6xWGUAUvQBhGP0Gh75Gn5OiDZnoQXPrgVgVbq2p9mOHOAN
XvcYd2Mn/dqOl7eSQlrBLZCsmweq3Q+ec9ldICRbvi/BIq7PqY/lI5BTxmB5TJMU
YuV3IlRXTWqNe5nt+DtmtQ/0W7ox/QUmFyRxjGBSEwoslcnDa38QoKmIqjkijCFZ
TCEn5oXe4tdsS2D0j6N4YXSJ4l/k9jvna2Nts21642ewuO/G6L5IixaBRzwWKn8G
1VfrhDUo1Yg+wWCCAzbV9lq50SzxDVmdQrR6YV9wRV6IEQ+x+Y3+oBlnbBDJR39f
A2Kr+761vcsdEC64D7nVXc4B16r5fzDNJT6rKmMqS2KSoAyGjSXiiVSV5e7+dU2m
WwbRB7YJf1qVRUpX4GJwI7fy8QeWOudaoFjAws9t+pj6HGrTYrAfWm1CP1+dXkeg
gOoMBMvM46qHJzxPo6lXh/Qfm8KoOeUOSlvlY3hgYLsve+cg5jOZ1c8x55JkcTNw
t46LNfUsEPpugTmrA1767z2RZDm5a4WKYSBRVRiCBpJRDQruRIv56ky+OpUPRNcF
De0XFRsSdOypWKLCrPsJSaQc/L/FL1FX9mSI6FwFQmaSUuEVwFPrnkLziz8Pd6IC
5q6ihnHPElTwQwHC+hktV3xuHH5nc5wwcIpMF2sRcuXzSBB6/smBX0FWgffuLmLJ
RN7kg9b2l1AQ0oq0Ije45k9HHSozyW9N3mYN4pG1UiRq68Xp/gAIaGelNHKwVaDW
Z67m/FBXu1hxOKddqzEShZfgNSeD5pfwjxM3GPWhsD4TT5t/bH/tILz1WotgALTI
Qzvg8/kexrMp0IhVMnqQEDsrscKbrve7BOkAwlhK2u51Cj3JAnnixtQzaSf/T6eU
z+Vx5KcHb2Ne+hAPq+azARmajSPh8qKcS3OFgqUuR55e2yuFTS+EoNt6iAadFBTX
AxmEKpej5A126HbIPzodArdA5dfUNgJBelS+jdemX6orWfgqWC1pJOERBt9kOwm3
A/H0P5h+R1QY91/rUzjw1L7bhDRjEyp1zIfZJpJmoRCNrq3p/Iv5ON+DRcTc4ufh
g6/bgNuwqBl206+FZHTLvvxYxoRbHj5gNqT60Rg5n8Y41zMrDkwVtA6UV9X5G+hF
VkKr3/zjm7BA6xqfgq7bXy0Opt9VLdQgt+mYfgPvyENKseEeba603yI0sJNpAGpa
JyCBVaIRnk87xEFiQaB5zDykWqQAHqjtyf0DgjYh4+7mrI6xE6rkR0VGNpdM5fkh
7J78yZW2uz4I3SkOWbxEWo4brUgQigPkFyGt+6TqF6q0Mk69JwfwXnl6FR63ipoW
HnXYo63/I5iVxYtGQxXK6Q6zCOAS0dZOT8JDPcUnm4w3LgFfpYV3mktJCV4k1azf
RNMdpOniZTpyWfw8QYN2D/d6rTNwjXrgmQryqKC9+XQ4Wr/bnfsbqiANivj/aYv9
8/t3lAPgMjfT1ZmhBWVlk0SMCeaBKy54bzTDbJRBUTQ5N3Lpij5Ri1xFdkYxjD87
exTgjRoFJJztCycUrkq1ttqOjv9+Ui8/IZG3SihVMoe9VcrHo1/3Ah5ZyxAxP2se
KgvBKNgE8g/gp0PpDx6S9F2NVgBhwFztxFOBXHsH4+xI3TBOl0zAP/176sfdyJJf
yBdp96QH4dn6+IoT90XWHbm5jRvH4zn9GO55LZvgWxqvIdCdHbFeumOeEta2bJH9
GttU7GmcidbEZDwCA8tY50DitOhR6TA5qdQKj1dCX3+r+KZjZtfg8pK5sk3BBbcL
kcnQR5n83ROfkHSWdU3xUXjNq1ZYd218RSU8ig5MDQevRyUsSXqfgmgm34PR/bIb
yUdfIw84wBTMjbrPr/x1QnuCEgJwCHQ1HgzFIy4Yy4jPVbpvH4VdvgLNJ0bDuhZB
DIuL2R0JIgCGKNss8ZvJ/ieSDqTrS6gTckdPrbyygsMhILd3+RDkxK7ModFgqhr7
d/BI+yFkvwlwdpu0bD3poFuU9ErrJ4M0negCs/xxU7w08WnTODqm4/ZN48rTll1H
`protect END_PROTECTED
