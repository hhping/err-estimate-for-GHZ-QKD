`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kTJ8iNvprcQuCwJa3OD98UZVzQp4Vif/5pStAutxOH5HU8YeFPNRCpZW70d7WclC
TJVA7xaOj5LucEYi31zBVmGhgjLEE9R6e2/CrcUDYQfaiXnfCBV/L8sEdOQnKZd0
eYASk+CH/16xGpSIiWgof5JInRZwF+2WJLJPLhJPpXgK5kUa0OLgyHiE5lH+9nvn
9unOgr6eJ0DgP73VyiFQ30mB35cb+PL5j8B6U3gB1gbzP8aIJLxQXEU2AvfWt3H8
9jiZ/IG3bhzuqCWXTWXNsARESERVQ6PWDW8faR/PetwnDJC4oDqKqXJmD3ORlliB
UXQx23kqof6XiIIXjs41DgR7qRkgdwHhDFdpCihTqH6n4b+lIidHHIbfL/Z5aaJF
9KK2khtz/CbxYwypqjLYA8qS5ZOlXqafGaMMIM0OCWqHM3kUAH+6CSv88OPSUmyG
AYQUkx2S5DiNRbAbTID/0zY+PpeyX+ltDcJcc25uF6PY/yVfxtrApvZHVx902Cq/
W6mdp3lxZuWcvguJHYyLgh1vdLovxbFgvVxnKol1lDBKDzHjB0gjzQZo3BaezWQM
XmGx9SVjytjrM7ViP/TjSW9kOBfdpfHl3IOHoQPVWVUDs5SvIAmZ0dqRaVQx7m/w
TPbpvIs0UdpRPb3ohc/I2oCHV6OzNeArXj9uc9kWbawKSou4Q2j9JFNcpd2Sj74z
JRJeEUeq1aA4hZ+2g1vqeoUVW0Dh8EpQNx/PhbEu+seQIq4SWNOoWOCUj6NUo145
6vR50j4IvY3vPbromIxzN9lJGi3glMbmKJuFMQbmMxtEfuGaAQdfJ4HbzS2VfVhT
7vfBL6odzysjHbEV/XhZG6RQQph+Q6FYcXx8kOmq4pntCx7QN3UOEAZzgb3liRat
PvPnn546xc+6PaVZgWDVOsGCULidEGqTE7jNhCe5uD8dJColLF3LzmN4g9J60+HH
FWAQx7dOFSJaRsFo8oQYAXh2XzyO///hxOBx4UykqSJaXemYRb1DdGwst8VDa25f
j9eoDTXHPgXCEJSIcfDWO5FOixX4X9KHC1hrgYSUaljj3y317DfBtFXwa7xrHQpe
qu3RBzlopaLSsdTxWMS8nNvNs89dMmFF2MdOT31OJoyIQW+lgLuCMeyezg1OtWL8
7VtZEcmiPkloRV8xn67/5Y0LAJsrSIUdAeCx1uW/PdXF3xXnPTp/1XHfmA7LBcEM
EvQytu3wvmqIaK8y7giUm31bHyivsjSCwrlprUgcfzuRJgWdxWkUZ0evZMFYT0g+
PVn2TvH1Ib3BeQnDs5z7OMehNCtakTEoBVCaxuJmgeT1shdKfo6Hdcv6Zmr0xhzI
Bn6hsGdjDkZ1Te+mYcFyQ3LTmDtId3zYXpiOypXQJYc7ZAFMRaG1VMz/aOd1fV99
NBHFWkvUnbqNKco1xe9ApKS1EbvD5DBQAy17ELuDbRR2THYd/BNeMTGJfI1g/yXy
/A6mF6bdOo0sGkePLW+Ajp23bdF1H970fO0QFNCYkwg+u7K0kyp7VnOXpdIO6bg/
khXc3UZkCo/2Z+s3ZW+ZzFkuXxoyyZqcs3SUiblQT7Zr+L+JuP3UTDMhhUOv8AtC
Ptu5Nvmy10gWPSNms8BlEYo9L14ZrUk6crhSYkImVGvPI8GlAkFL0MoqGsHaCqHE
KNymxzWMUUK1rs1hCGSEHzt0tk699EYUQwCU2NAGB6KiCgdNn3a/En7ggfwH8Fw2
nzuWTOCJw7FtkFooE+zBgkDAANYNEb9EPexuIRHAG62vUy3q7gcg2inaROAQwwe2
iGaOgP6vmrmgvAWNirCg6SXm589ql3SVgzTcfgalPj8AuQ0o5hKulEuKQp5hiomU
OSSkehrNo9+V8igsu1VlUp6EFrF6SEaRlyhDc1dWykgaeZI4svpBDdtv6lIL9Cs+
akcmzo8l9ZO9lIkRktFW1lUYeX0SQ5UyjWpbVGC2k4cx5eK7miNf0T8owW0/8oSb
SxGz67cFsyaqVDxOuVGUogOr5eWs+8pU0FP/uy1EWJS7Xbiz0ZW4TPbizDGNw9/+
OTRtvFw84wAsGJcVdxOZhK1gtpwKQ4dyTzjr0gxXGfAuZvPtUj35hNXnI+nAiGSd
jq14qHSzET+AV3cbVWPi1K08SBUIHCSU/pc7VDtHfHqX+gxqkI2N3tWSKimt8b2/
n5lbC2FBw9JQHjrit6hv/M1Io8PejT9av9SoKJR3gAdKD+G/5+P5xt2mQpvIrst+
bvNTcVN76v6dO6aebzrUUw==
`protect END_PROTECTED
