`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3vcklVzPlPv90wjOFAHg+/kW/Fq+7bOGz3z14/vz3ctkI6Hu6+FX6xa6uvkcSmf
uChhBms753ygXSTvIYilZsCdobhfos0z1DcJHU7/pj0cLc31Wp/ay9qij6UcMuLH
MZvY/yVWKSgRQaxz7B3zK7cZaCtweq3g04jiZuMccxaIwOQdxiGPt5TXscClm735
kZyWCvPgd/UVv/gAQJvdSE2MRveXbvnEaud0j+RGWs9SWH12ERwCPX4gcby/KraV
bAjco+TI82dkxrZKN8mB32dKu+FRAtOmbo+9xCsfBE4WEHyMSDPTkXymoOWwU8Z1
bID2JOcE/d/lSsgeQNc0RdDJMc8L/4fCfoJQsWQCdnTBGHkzV+BUUfYXEpfSdOQS
9yi1RfqqiCuEErura7YTMw+13tG3lcreEjbdAkXOQNkmnFT1bC/94t/td/URukFj
zUFEkyz0wCE+1aei4ziALf/Je/FIlmCTE1bZdkocBxibAMr+PIee64ONMKMqTi9v
bYkY4LCqWFjQG+pXHzm+2aXXIjvD27n1xKqqqs+7/jW7ZpEc3Vd8qMcjTlJ8VLsI
5VKMbOYmQKgINM+sC34cTME6xVn7TYo3z/vhnP0vru6vYS5r831E7o5ul/LdDfWr
qeS+CFs9kYkeSWrwTpPKia+tr+OY3zi/HJDcr1pxfU0IndBqV2Q9bYfjLG006Fgd
vnQh/znGFdVn58EgBX34R36uxIPjUiZGb4N1NnX0w0vn2EqDR6Cw1iqlV0AWvd+l
N0erjFMewmjl9N30fQZCEQ0e9/8zRwvjcLVJWM9xMv2j3qWwKYPCtBRbu64976M9
BdC++NnblW72UVvU+S9nWr5CgFHgi1UUy1OAhCkHWldgl+cmhAmrhQfpb+9lR7P9
covuaY/1wzsNZ721hv27H/hhEn4XlhjQgLzicMUaRqbTN4AkXD4RkrWmVwtYiaPP
u6xraRgHEi6WH2YPaKxepmUBW8M5cmFtNAz+tUPsQfwLSR06D6vC/WZ3atZ+cRqq
6MI6+D6qj2+qMK6qzriRjnDYz1SuMOPUmkPytbBw6SKIl+CusQWS5wTra3LHagRL
ju6LLhzDVDvZul0eT33O33aJbOCQpms+M9mpfS2XcnU+/NfOBWb4Kte8AHpQoM6J
KjpTr/t/QL1BxUnfgHPrHjN7qvsmkr/mkmSPG4tFLaaV/YLxuiOfUJxGtHphiQsF
MjKtEYcBG0kD1SmmzTdUonuaR9WZiG3Rpn3ah7cG/xCmpKFZAVa5f5g8vPa/5yWZ
9jBLgCl8IpBVLbk+kFx3q5EO4fzHhKjTbgeD87knZGFdlXk0GZ3C4h2hGfUUMxaP
jNyOUTiXeW2PdyOI6wfz3pqYpfED3u3ckuXhWn36MLasT41nsdMRPXbDRgiL6ZAl
FvGEF72YPOf8q0z9WnU5J3vWrliBj8nKgTUyF2JKIh268VG5qtWs6eJPyFuJcCPq
Y1DB7HtaGQiFCJGBqzEAbQK4kch5WV12WVnNma/1aJP108o+ike87P53buAC/hfu
QEhwEpa74K0xrU90f0RuoxzJ/xJVUmhsUmKzr80zlMmIYMm93pJLjdUvBPI/PXVc
qUBamGmsbHe2QjUZhtp6B1DXh0qS2bCs3BueM13S8A3mnkIK2t2D0YjfIVsWhH5B
NHG1OaH0t+XLyS+QkD3Cyu3Hvox59HfIrm8ti+PcBP+PJCh2KwDHeVRNWC3zEBmX
GlF0rrncBJr18rsrUAdowc90aQ1jcPiTZXNcCbZDYK+B09QKPlLAZrtyd72NogeF
4pgpiJKY91djbfN7wlLjD0AAmmjgpqYc+RqA7hXIy6dTbta9PRKT0F/SgW81NAfh
Hj/71hgSU4dFGTNpGa5bZ3dIlb4lOBzOgnmnfbYQFgsZXAo3e1LofojNa5jZg6eO
`protect END_PROTECTED
