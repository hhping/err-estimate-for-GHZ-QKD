`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yK7Bbp1XazENAXc+4yIeqOEOwcavKUX92l27OikYDm6IsQS+XQBGbTWByazIZr62
BsS8zZPPbiKBlZ/vFYDCe2Z8A66WKFWTEAj+GZthHgOXRxnd4bPxCQFMMFwBeZMd
p+DxrbmHsbPEZRgr7RE0Xka22AR3gKxbg7SS/6EkWazRMW99r/gOla5fQmfWXTIx
V5oQAiUvLuO8Jhz3rlmfH1Im4Br7MTtXwZNxwhY03DFW/6zDqYmZDya/HPVB2OyY
fiS7AaiEhR+89cqCkrWmNkGcf8uGXcoFRJvGu/FC9byUymm5oahwVDzacM8efhqC
4kJy8615F2O4axVtRVWCGZwVGwlPXKwVypvrMyZntevbUdPclpc9DGXwM0N+zO2B
Q1/u7Yhrz0rFxhk3jG02nr3vgbExmHBTXn/bMREVNHd1p+GMUNQ2Q6fc4KfM6dmz
9o6AUwItGtHICJ8KqKIOJp6p4hNPOfc+x+aEQxwcxIalurvmwYo+8y803WUxxjyv
8LJsystEKlds2T5d3poh3s6CM9r5HxQhs3cuemoVVWIrkYKpKO2kxYOpndFu7Xw+
W+fscQbhBBXwvYWVOFVfFjnXSqJ2orY572efHoWd4aCedD3+uq9KOMO0JAX/KIkM
LxsZWzrCwhPB1RvkDXoTzpGK438jOSxpJsXVwAZKBx3vdMThb8jkgzxVqcN4dGAS
0MGKrD8vR6mvriuESSSMhV+0FMPwCPFAciVJZwMy9ebPj4vyctNcSzX6zTZd+c6y
mBhEjPsYfZ3nWGjL3OFsWrigJ2t+H5DdvOX0TVEeHJghXF7UkwKHbeLv9aZiknW+
xJEOUCsuWzTHFQ9rRDUAkWm+B3JRNxqkvsuUDva+deZfc3JvvMflXHLd5XC+O6BB
TWWkWXpT/NCi7uNXRieFEMmG3gebM/TCVgsS1v8/liKbsj7Lx756VATJFjOyWplC
gFo3bvBBHXdrk+LWcgHk5HSX7SGbmYq2Tk5YttgbsILkZZlHM3g5Bdd2wRSYdbLB
aEErdltBo5t8Ak9VVlruE+kSmBPQnbKoS6FG+Hu3Ow7pIL7j+VZ3jIWu9XBiCQvn
dLyMgeg8YTc4G0/Jtnig+qZKHh/q/i2BdOug882jwGChhRWQqKowjSZ+1WiEfSYj
PLRnk2WxNXcqPodp/4rhcQBYJ0hOx7FELDP6OtFaS7yW41FTSmjXtGdRwZC+4U3t
o4NtNA1blpotSmB6Hjk+C+FlBUZLsojp1Egruc7fyeJXte00lHEvlIHe9++gnDW0
DpsxtMZ1/CW4iPotp2qy7SkYtThAvc3S376Nk0fhNYn/Bw9q0H44/+NWQ1SD+48F
GM5kG7E+FkG1REb7A+ob8JOwZsZlmZtWyPnqFsWm+OHoMbGFHTqc3VO32pR1Ds9w
TXLn1phX9gdjZDH15bexpK4kE7lpAJ57sXkcscirfX6lpCk93YVkUt2G9dbgWg+W
oMzIgzoNrAXnMoShUWoewZPwAI7wcLTqe2h5SmdGItuoqpaQASiSnRtKgVtbEv2d
YQLCGl9oO//6B+EQlj1S7u71ltV0lZDxYf/ki7zA6ydSrchcRaa36EhN1asiJYbG
hov0jcL8POneqYwn//g3lYR2dOh8wOhEz0V4z9xNTaX77U54VQ/6qBTC8gMtpww1
KL9lCsDSW2VaYSih+Uqe94e7DmejbHdopSU4pwZpBxRco2/ufB17k3pAfaw1Gjvy
JsHtPK6Twrbn0vHcuKdNdt2w1e8yXU/ecNbE5UCgvKN52yil4HaMoR9BZYnwsd4Q
On4zRSNHqrL2KY73rca3He9Kzcu1WUeo7Sbvn0qI6AEUfdGDRZAoNyjpCRMRVhBH
sHDTOQvAoum7MaxSBZ1Rl3l8koEnn/pl5/obwn0NWNHksrC2ylyWsbCCST/I0jpj
KLbY5MJLvgLGSHmN8K7rHbTVU2vccp6XXxuqNMSqIES0UcwAzCXB/vbvwztJwS8m
QgHIM/hE1/al/CcpGdYVU5wvcwR4GJaLTlLFkR4HzAlws1+cqj1WkNhpoj5zBqiG
WHVMYlvCaN+xRdoGeP6C5b6qsK3xIYr5TwPcJAHp+9C5IbZ4ldHdDXeCQ1tXhObx
YbfdtGKXzhuG1kGq2jsLPl9p+dQDmouZFiR2D4Md+csfd25oSI9wZ+OhUYzpmRKy
SaOPyV26kMsZOSvjT0dw4T0VMN4biRquAd57YBzOEjtD3IIuEqLg3igLI8HL/TbM
tSnRg6gXi9JSXOfMx/PkWb714HoT05idLD5smqDRcCLtsIKURT+xydKVSZARuoWu
w79hRw0xjSa04m7rjSugVJNzYMqtaEaONOhRguzmkEJji38MN9yPTejjf+GzrBQt
d2dtOFPsz+hWCLG/hCl1Oxj6JJIfwLM97n2MlnC2LKdgWD0UElnnsm7Ov8sVj2Q/
dvKnoGAecnXMJ3YX1CFG1/YVbr5vcSGvgF1CWcrjfIE=
`protect END_PROTECTED
