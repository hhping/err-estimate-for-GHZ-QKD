`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWzGP/WkTq5eTpxt8BlN3IdGnaUHT7gxXYbqhEONxk+75bKJgrz/udnwmZgXn37v
eD6n0+6HmLLVoxZA7aaIsjUjuQ53fi6fxpUuY49T2XwKI684N1wgYFCbRLoNTDVo
xC8P+4MMdeWNuxfkMWxJ9esMSjuSJHkbZ2bU6OBjkM9wa3udqF86ICRPjYre3N6K
dGfzgyt7ZWdQlawfUwyy/VqtbGKv9Gk/YW1MQwIG9AcQ20if82qnMczj6Uya7wAU
hUDzf2UZcHHx3K198YCS0GsbVPi4HrrweqzqQi4OWXu3E0NOvfitNHZPXfOrgVat
jgetrzNFDjXvQ1SxWl1AKg==
`protect END_PROTECTED
