`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5kLmyHBP7RW9BVE2opsu011edJMGfjiHCwXFNf+cbb0t7PFHrMZPNTALCDVFOF6
L6Njx4GxLTbtKpdieN92blRKfTR3Qh1UlbuvSK23HoGzbvpE8X4tnd4TYiCGGbAQ
yswWfkUkiltxa5hFNtFfnIhKbTuXGdIVNYYkdKiL0DAcnpgVX3pgsZ4K1llX0iDP
qbCGSKxv1rbyrzFA6/j4cX3FtSiOCGsiUGpe+l2xExMKIQ8GFhlXPlIagh9i3Tgt
WWoP7hEGHXazMoZ4vqs1AItx9bJyFtkjgbh5gz/gvzkIahkibAQ0Zf6sPfaBRT+a
YGskCa5191nuYGk8tHRtBCuEklCVqLHbT6lWbxFSANN2xU+hWD0qEThfdBTiLSIq
TkHF6HhQcQve+UxTdBAsMDCG8cwYKDTwW5Prpwy/NCeU28HjHBl/ns7o6xVIQvA/
VpIkUC2Mb9BSSYUd4XHEa4oK29eK53ZqXVrQdvNGNd0mPTr1nFUDQdX8HFnqIPOY
Y4FMrsXwuJNoqjGjo5osKU+30aUF0VH+TJKc3bCx1HUxf0nXd09YiR8NDhQZpZ2T
Vj328yNBO/LBu1L3hCMW/uBjOQLS46RyFfCD/J1zshxdZHJv9KCCBVenAAYXTGiK
yUPUfaufcipc9Ecf1uBLzOMusRpM+jZFBNQhAMT9y8etQNqRexd21vRcfFEbTGZz
nmxy/baMduX2yrKi07vjP0B5V51vXB0jAvHoRytRDmV9oe6cmyj97MmzQNFEdA7p
PzxUiSKZ+j11NH08wNNe5VbS3FVzLsG5c8VSVw4jKjHCS1TxHjrtwbvlUWsajdc6
Wn3jIgfDx3QevoIpGLccmwDtTKb+rHN4eVNQ8edYTBZepcMVqDSkkSANerLKm/a8
IE+0L6nReBhKn1dO94Q/L+76ij1sJ6MeA4dJJJ6Uua/HPaxAJHuOSR+K2VFvUliG
JGP5EJFhmFYg1/hEU+gsrwBAqtjEmSl64Y+cA4ktepHpJUSVf8vWqLwbtmYWMKBw
EOfJuI8uQLRNoGSpmGRoU3yXZ6+nnkMsN8Z6oYa4vp6ehfq0VDmvnr2Rx7ajRs+z
3KTQt+3dIE6+Nn90jXWbCw/O9CovMUUZg/gmdP7IUKn6n4Au0ce5aPm0jQ2Gv15C
w6A1EJ6oej9XS9VC/34V5PXwS+ZZxVsrpqd1Fgu16IGWXM0cnLdLb1+whHHakyRn
h+BiJwMI8jvQmvIkQgRobMyZtgfVplOKIeDQsyNBI+8QWAlvgfaHfAhp62MfbXwc
07FstzKBBAXC/t8doHjCBCFxEPa4nyYXF7LtjnzrhRQFzkQEcZJtndMwr9acACoB
A/Bc1xC6CNk2BafPdmRql5P5hWxcEsaK1SFnxnqv1GrOQ8rPHceW9INavPNtbLUD
0kiQpuWIwqfKhS7c7U2qYwtMsOUggbF9UbRj+qxGt9EcqLjRKVAdeG2Quhxse2+0
3x4NIEHfjFBt5djS7UMN5A+6scpIlRE14lXuIg0Jzr3Z5u85S+i5gKTgxR4Eolus
wUSIJYQkEl+IZ1zPSWmasAmSwFADju0XJha4qspZ3YcyAaFk112RRmOrm9XItPgL
/tWWgcfkZgNq+lOyKkAoiSvFTn445GGRT32yw6mK2SyfItHo1N2qOAYY2QH8J3nM
QTpCUPojLLfFs8LQkrg8CqmFBZPT9nD8ouGkFC4yW6qdmLRP+pFYNBdRzHhhTEAn
D8urHWPutOlW0g11fxlhdyK4jpOvy7cnjDNo7Gz5GMYXXOWNGftVREGLBBeXT6j3
ZBK/ABKKnNJEoJrgq0dIrug2oQwffhvPVTpmOLDKFVOVk1Exjo+i4880JstjLxzI
7p1odCuqbTnonQqjADEFAzJZ/ddVnRbxU3lW5sk2UaisHM24vyx3ZoT0bmgOAKB3
+PdH0Z28fNGf5xSn8DP2IlEHsvVGTaKxCvbxmlKtupnDCqat4lsMa0hrCCR3Q5Kc
nCjoKLe4kv6428OyEDSy4XrSubTg+CvMtqxigPkHgAnZX+VAAQcqOxdqHYBIIDNe
0M6TBCRXhiP+qZJz1zOVjd2RrzxL5/GQdf6wAi2wh9d3eyTy/5yRcn6nhJk3Cg9Z
9vwmE/oFHjUUWx9WJS0fLZUdTeDE0zHAm0lD9jQr3bPPj+MkOIDbGN3PmjirmMzp
SnCIaZpdH1DKDv7bXFdzVN6dEPdgJ9TibahAx7mFNhqlvnqTaEjRnG/HnftVLyCL
Sg0nl0bQ6U6DQ4TORUByqCUvbAdPY6sEogXLLFXAeN9PLsOt5z+bKewKQvHTSAFW
cZ5cIJuCQz0XKoZcSHSB2oETNVAGgImACPKW7I+IXWXhXcvLTVIWM+XiBdGDsEFo
2ag2UgUE3ka+3dcO4JcOjLuKahHBRxIJ714PELue9T88XBOeIvgGnrdjHRqOcA6S
u2brNvPPpV/jjDBSKIsc3g==
`protect END_PROTECTED
