`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZ8+dQG4Rp1siAnStDl9EB41gcnpCnyFgpzA3HHvzhzlwNzncWZMBALNO1LUTURr
egfTr7nZ0MnUspsnnrZ3oLQsVNercquVX0N5d/o24q/dLgOIWBdaoFAj9RjjHxb0
zVrgXU3VrOlik/T7LmBp1Evaw7WDDDKwJgMAvNLnk3skcSkK8HvjoTqz90LxNQwk
ZKn46bGf0YOW5+h5U9uWZBq6YiF0S65+Z+yPtJPUwxhP3/v5+EbkXpXa3DXBbyOK
Ry4SnZIZCtZA06aBj9wQtZvVpyF+5J4uvymOqbZ8goV3pUVUqlz1Nmyww8FRfXrd
lr7vlnT6CF41dmSahnBadXcp32zYH9b2QAm9UVOkFAr3teFRXEMqV27nO6N/Fy0f
z93OF2eMZdSG3JdKmWV1osdVYvyQcIKeTab3h2h9cDnyG3d5qH0z6YSvlbjpdS2/
iQbE/vbtVzKEGdntwsm1CjdOBjrXx9FVvhOjwXgzfatRuOULMZs4MkNIf+eZIP4+
/dxBegUO85N/P0lstC5jaCfeo79JGcYJWv/7GnESa6DvhaAgppMWcmoEB8AZM1MF
UIVYecZQxRORTq4xYcVqMo9tj9nMRe7eszyg+8PQseQXuSjgyGL68x+IiKi66xAb
xOl7olOFJa7dRgSJnaVlSVyKPeZXutSgYkrM53U1YmZaLp/2ofw1u4cXpfcr24YU
Vw9Ji6cKdRb32qZLGYag5NWduWb/0o+mZffqhZ8VpLom00oGrXTBE0XkmItIarvz
MoyzTZKlnmkzLsq6OJUMlfkUM/3W1D9aFGEBZuKuw2gz5Wg8BzN8EK56BpUFtlwy
fr+LEEv1EWubgqCD210hVTeA5+t0d1uCbPHCuUCHy7KqzwlNNqJOrTXnfAeuoHhb
XttpW4CkxbuiK3G3RgtIkN77vSPF6LUSFPB4+lLUxUckZLEmGrOUlys0yKUY3Hnt
Kts9ruC5XmRWA39HuWbf4j4+OAbZt8ftKS4XLpODJZ6Av0fnqyZir0Gy6F8Wx7x1
fFi4X4BTevmBDv2rcvtsPmT2BlWxB1ir0zSRjzNV+BH1CYiNah1c3Q8JC5sk2pMv
LulvUSyVBWqe+U4tAf92rGMwDShLCtHqRyRAYR/QYbzxfXIwC3k1r6iXoGIkQcY8
yD18ttdfdHWelFuOiA4XMdhSP5jGaVvylE54YRcbla4MD4d43sawJieLET6yz50Y
7ABq/PDnNVULZ2MAYHWRz51ixqZp/yXMOPc/vgZnjERLpEDHH4dspgXPvIxVA6U7
lQEzk/QRm+sT/sLIiKrYbbmMHGI/nRtDXQ5AIMzCpnBXUog7IJ6tRSab/afRD+tC
u06hwDF+4a8mYEoN/b2ENn9oTfygZrPSueERh0piFxDiHeYxnkEdr0rtxg09+14E
xRt2/i5eAwyApFPVlEkqcJN9+fsQGlUQb09DyVNKISYZfxiyB1/hJJQMEdZ+Jkwo
o4zvCTvmcJuAv4DrXKVnow==
`protect END_PROTECTED
