`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1r555PcZxtMigxFOZX59s6E5FIwt883sDPehuRMIbG4DRyx9qqRd7ySTWY9Vu3Dz
815I2GnYgELpU6dXOVz7RmhhyGgHxsc/HTbNtAlm7t0UEBZQFIHAOj8w3Aon5AjR
KQbUY50SdxlNnWd9T3I7U1/LGeFeeLApirF0HKnv+M+OXyHt68lwBw8K9thRw6GU
l8MeLsCTHF5tfwdyPgLIKzaIME4viQPx3Eu9TQMZharIutQUMh2Hvmmsxjnd0Dc+
/jsOuQFrt+I1xzIkqCN8u6zf0lSdNeBdYT2fDgUHZu481dP8uV7lcyKgBX0nxBYj
yUGJWnI978FkK0OpbO1cX926UC/bKJVDgI00SV1OzGCcsQ8YSkP4VK7x2r9gNTQt
WqKQF7EE3Sb5IT7JGQIh5fUFTtB5hY8Tzb3XXvqQgnEVGL6r3qz5meKJttiBc7Hj
9znNfl6fUivj5za1ArLvTGo/4sOwUJ5MMnM6cNrQdH738auwZwdzLakK0B1t5h3T
uhAWLeQvER3RyVmf5KZTWcOY4O7mzwKZ/odPafoQOpGa5AWecZxUT7u53pu508/g
iF5ZyAie4rlxM+CXFjkyGWWzbv4Ku+zTIJX57EKaVUPntpQnpXvSGpYwYqsWCqSh
DnjME1dJ64XwCJi/KHKzeqg7m0+edhw2mjXbCFW16w36dwicfqUQGur7hMF79CmT
0amP2kt0gWIr3eEVlRMrYaBgzyKNQXcL3fW2WpzWyfMLEniMkzQNPxH6CIGQcuzR
aVZuC24YC+0JzBphw8Ax7D2FcBxfAusyQaplyZ/AZ7803d/xBuz5Kpv1+LPdKPLP
C/20EnUq0Q6pWLjOEoIw+2xV6bYbsB8lIaZA7tT6gFL/MvtUCO/9SsLxaByD00fL
bQJg324/VGmNH4dT1Aqf0udswM3CybOOYqVjNAf7/et6l01Vn5uWnchcfJulADfv
dHmIO6txHEn8Eqx8xHdRTO8b3eMuM938nKWq4r5EImUyG+7926fcdF8v53VYkH3Q
wm/8PIFcKBd85kMzhd2xAY4oGV4bdYIBw3oQg5EeE+PU86cSnvVHJQwe3mZsZ9DK
ubeVAN8SqlFafMFcv6JfJBVf7YK1/7bmrL/QY11U16iAlw+garFUPJ89acmjkW12
anJNmDZt817euZA+FHJOdV5dlloohg1cBppzBUi3ethlOWkV+j+vl2qcXjj7yYRO
3uj99d7wNcnQpiONWgFRogn1N4KJ1k0PIcFmt4hWOdupduWcc6f7VSB5pfTeCVxw
YotNpXa67egsajlEnq9YO2NGz30ss30NryuBas+RK903go32bRxWCa7AyEIhc6ZB
e9MV/vbX90zWMjs4NpztnHJ5BPni0XMOgDT92xXRUyO0qSvmixtFQkaBBf3RdItp
M4tD2OC5BVEe2K+kcrz5kpKMV5kG9O0ZSUUWpitwQAWpv/beYdpP2JuQ9897FIu+
yEcoEK5DaE/v0ugWdtK4cQtv2/CaMX+ZkYtmmIcUp46EkvxYoUZ+NarPoRJE1XWb
l2KJ4c1eWRoufkDeZVqqvBEpHZj4XHw0ucvOXDuqPy+L081Bx4giH9P8zyzDotdI
xhnrF3+p5jTmTYFXO27op+k7RHbFToVnHFIQug41mposSFIpg6KDUqM3svj8FuOM
1VxIxy2a7NnPLumi+tsQjsDJPESuPDIMHOSxIDfNPVnFhcOuMT1UXgeMrAGNbw8/
zbMMXop4HPovdWOdXZVMZPjTiN7pJsOTjVmC+CNfFomoaTlVxfnFo8d9vM+x8Vuz
g8iY35com+4NPv7PQJzId8r/aypmvNTxLU9XepcO8cd2op3BwN8Ces8S341BImVp
sEJ7Fc9/c5wY1cCWJU1zVw==
`protect END_PROTECTED
