`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqCgevn9LC2UgRgLyL7hJgerSAHo5AVvynnEfRe30OYHLhA0g6K6/YGdyw7o5PWv
8LHYVlFbfkL7n18GG9gT/8mWswtqnwGD1wB7bDbSqQz0jo6Sqd8k0vWBZxUtP7Yi
acaRXSCRhkdsYwt8MjI+ORODp0wz71TplQVpJD9tO7ud7Ug5igV882YTptK1FZv/
eMvGtsVQPDXWjcHtX/wIKMwwuSzLp8k4wf6d9p9yjEUD5BEoNR86dOstcGzHkJ0B
R73QmT46GpLYh64uqewLsmwahTa+8+Vj05ryhiWN4dvfTEfrdXAW/nAb6n8OG3rm
Fq2CBxZEZhNWflA8GRIzrugE91fQa+EdhM4DEGTgNh1aS1FeqJylOyvQNUzM1yKB
HsvUQu5zl0xMzvxnPLfTyUNH7ssnO6+dbw+AxMI7g0U43zNK5Iht0hZ4jP1BYcxJ
Ip0rUJQEi3ZrQKbEhjF8bFh/O0EqlDHbqr6PmWf/KYDzGTzN53SrfQVzTdn2P/MH
kp1oKb3EwVyXL0dowAkub2BQzX1eOCtOeG/3W6c6yKdAnyczJaERgev/fwS+8yWL
jmmW/ipfbm1fmBT3q/D9j8hAKnIMwR3c9pzMQ9BOrhccw0Wpiv3t0S4SiDivrPrr
Kyq5qNlGEu7uQ6zUK8tW22bKci13KBGK8plNKjW/5J4AUa7Tm/edxzHGVuGd6YDb
jxQBVC1oq60VA+UF331RR2mb6zqgQobz4v16hV6uxtl5oucbm0cKsCvdm/GAR7UM
p8UGATevxEGC4+QkYwic/gfLJTEQYny+S8DiLjsX1ybWuCf8+Rpg15KHdGCRTy8F
cGcPVdlvxXO2uwL/L81PkKFsRc+UnkB/x2ROpe6mFQYGYWuA1gDY2pW1pu7GeN1D
ZggUfDlfDVy7wypIQkARF8WphXIcnGBpy41vyE0580wSBm3U6vCBF+x21s9qiQE3
+eU22VwNSdiEV6ze/4Nt7ktojtlEB5DH7liLh7Edag6bMCSGoW6cgQbwxleMiJdG
DLXYoqooMyhQSTL7BKOr/uIPS7ebhjEk5X38hDqjD/Y8p/EhQELWwPz/JhCOASdP
LGvH7NHyYFLEm8nPTulPIBIDw9uF0oPDCGCcml1O5joMw7fZI3ginJ43I0d9/znY
`protect END_PROTECTED
