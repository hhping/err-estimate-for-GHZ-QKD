`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ia7DSvy1f3v4m4p/ZqbMnYQnj5K2ErtwUhQab5fyZPaAKAiUttmTAIrk50PP703q
JHOzFi1pNaYyCcpvLWar63Lxn20KB/Qh5JD2KmwJ8hlA8zv64voh2MwICxnMlPBU
BtbZUrMQjHfD6G3KfBSNDi4lutA12Q9CNodE11HNQNYY5yDZC7ZBCQHIHSXdO2Vm
eahRN+LxcrCpSd8nWITMnIgi2l67siLllCfMZ9Cidhqd+Nadqofk6f7J44mnWASl
Fafp+Dqv024LWZg+tHIUKydzmWxMg5R3ofAoJX5Gl0SSHE82iirwGOAVsJIU+BDF
9X/k4sLmYsHxMKnS1IsdXELcPNYqt2owcgVWhFOFUcuh2DZxAZkSxMo9ld46HFtz
oBdmrqxEyrfGtMKsmKStL6th71LNnJnf9YGOd0dFOieyKQKnyq0GJgvP9H7MiX5k
JA9W2L8ycTAeJtS11VOOt9zmGhoJRdBtB8ObZxryCXvq8kBdSzjfrocRJ6YBrDia
vGhhmE0E2KkBryIdLx80H2upYPqtWkNikKiOqXJxuC1Kf5oy34p6EZZbCGylK/RM
/38LB1j2APwCpD51OWA/jyZwNhcMwzfpTg7Q+siRdpiPyQfMMcUgo4TSJntVc4+M
TS1P5PNCSJVfz1jramKox73NK1dnb2lx+cM7jfnc49IFH+WvhKJngvbdBPABPyUO
oOGC3EfCvKRAjmgNEkfzVSH3YjN2lNcDIk3AKkVCMGUkVbTTJFhhogTgsX7aEUxY
`protect END_PROTECTED
