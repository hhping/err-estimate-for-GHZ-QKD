`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXVfB8L8+7gKyFWZLkPtEH8CX95UJYaJGrz8J+jZt//xb+pIC4Iwu8VsUAxDyaAt
tLZ1T8xTVT8Da3bDT3RRbPypYaExLnx/qmYT2OjqhIkktBb4CGzDxXt3FycNoKjW
11m8cJyUYmK+pGXomASaNHvCdubbRfMoSjmnwyvzITTQSPvTBxE9u0z9o1R0BJq+
kALSmnEpxa74sJFjKke0TlBUSZgkGzsQ88HPOzJUJQdC4m1Gxdc00+9jc5waSfvG
faqh78LUbl6WFNEGi9iutDlMN95FpYV4uDNNjT98XSSXSlOJji73PhtarTTkuiVt
cFv3ujO2v8wqdwzM3GjuYyZJ67BetKzpTLwmh79VH9khMaCVRQUecXIHYKQKVObE
WFMVXbqimEJ6iPstCE73EBwh21Sof+OjX3fYWfTztEE2r52Qt5nDTDIOOMzzbBAL
HkMcVB085KkIhX34zGSGPGAInG4UZLL4Csk00MHAeTK/E/Kq7TKpIrZvbwIo0dgK
ZZKV/wLZZwfya4pnId6I3OqxAH/3HqWRM0Z8mjw9Fq5rM88pdOsrEPOF8BoQhbsa
y5wh71oZ88Cz2BpOhq2y88wxpaHZEHx5EYmQ+9ZVaVYvnpUa5FAAKD+yH7uFXkiq
mNcbignV80h8KBu/LCGB1oANiHYZQcslY1bxRdAxS2gWDr5Ct7dmrWd0/2sh/5XS
MDWInkj5CjaZ5TeteDfVumO0r4/DZSebqeCNIgQmYqeONJ4ddZYYcyECjUPTmkWc
+faTcsPQmbZEOrMR2fY9zaO9ty1MPc1DDRQ1zEDRpbxRnr+w6swA8TolmldudxfY
TcbZJt/ttlwaazpynyUsqcAYk+DwpQWxV8DndMqcDknBkSZk7H3iO2w6j14LIQ8W
IYx+qoF4jW2FfIrgXLYwuxGDFiBkkDkRRwHozGVl29/QG52C+7sA1ZZrmiGFhH+y
AsMdGqJDghHVXJHk4kfmT5w7GB+jbe/8mGS4LLh3JymxeCgYfAUuJg+mVaXE+B8I
9UwOjTMpWyj7cOmCkexPorr30s4HsnqauAzGlzNKIW7Op7L9PD5csdtaHhQbfCIa
ptp4bCTZasPLL4xoTaoj/OfM0ruude/Msfjj1eZmIc4PjozBKNW94sv+XuxJ4VtR
PywPryEgf1fmOJI8ikSkfJ2hJQkF30rrDbQnEAKpP/T0Yh6gqg9GxOu/EkikawlH
ADMwO46KvovsOnogJQCOg3LATPVauqWWJZOrIdh9aWIMLym1fImbLg2jsjd8n4qC
5wYExTvq1N0vC91C+ys8E6KK3V22pYbPIE3YF4ieCMEHV2CfjqDoRMdo/zPBQcB5
z3MNTeQ7lhLchKxhX4CNZA6GijmRJy7t3aWnORxzC44=
`protect END_PROTECTED
