`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3HnNxrkxadt3vZ9cziTubCeEHH/f0Z5TM1ScYSG10tDxaWp7s6KrNuty2w22vSm
UqpbXgGIeZSNLZrJfJXGsCFWiKA8A2Q9ntqpCU0vCDo7ItdIfZ1ffR06ZA6v5Ixi
ptDkipgULk5XBGt+HSaI6AweThECkTfkPQpgi4gCD+7EvtmN0/6G0Qq80a1JVdgQ
OA5EtLvvu/e5RqGioajw9zGag1FgOrxPD9d0s3SFAgtcwnSu6hDI3Zgeyi+QMbMJ
maJETfoO4F+shY9TpF01n1TmQQfXo6OQ2IujE9aCWWLK56WtQJSimBPJ/v/e2iOw
ZDUrSy70r7CuGC3rWb1JcrwVU67cpK+FoN5V7zL2GOebzEXmp1aNKVb45F9l+s1j
QaMg8a6l0LqlBEYQ2UsN4E8kcD53DHtsEEtbYWTCHAvt+6hwWdyk6/0J9+GeHx+3
FoEe+9LPm1cwZC68hx1sfLbuGc5cO6rGQ2HyMUxA5NQCCiSUkcS9HWqWVbcB4s8r
MuijDAiZI/RY8b2JTVbqWbUwiOMHyFhLcUlmzWlUB2FbUbUwQmojSY1RiPDmuj9w
yDztP5hoWlTL699KmlUpsbtAvYn5MooN3e1E/DENpo5B8xKKvXSFu2RDqCGElN5u
w7Blz/iUszOJKkQ6o78nGfPGcLA4WBFsiQAY89EeZ90SemtF89+2g+YG0cqp9kGq
Tn35hg0eKYrKqXwcmqpBGTsYfoCe0Jk2F+WNDRvqXg72Y3oH3dNiluw4Z5NOhhh9
cbBuY35BzrxrlPsW0NvkjL72hkFCVvgcb21ea+wPIJ84Ta5oEpbwy9i4WOhw2TPF
eOCxvybPthziPb1SzQV0Tr2C9BnFBnKmYHVYhLuFFNsvnu7FZnjS4JcC2LtxQgGc
JnpN5NUrTdPQeFHw/p5xPHWpH1kMSIyWQM5trYa26S0Y0h355m1HpJ4O5FhOkWqi
9Kv6enrX2/WJfzAmAigjdbEjOP0GOQYLyNKbhuoqitnpDq6hSXPzclhH8TR0To59
+hql77+YLZXHibaOYj8qqJd5D340Q0mZySl/5EHyLD8=
`protect END_PROTECTED
