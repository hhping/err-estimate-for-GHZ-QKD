`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ay1lXHi7QPqyaKit1C4mPPejS60C+sPZHxYEr8pKO7p9rQjUB2obCZzsUdVtUMlI
gEmJzNGXdmHXBcFEPlWwbvynLmOGlNm0FHR7UBIt9wnhrTf/VOw2WVSIdH5V8Lks
fPv7O3dgKILuQNbPTo7aLyGIqDXeHa5iQs8NnNAZX7l2bPIZBGBmeFr3A2/qhoiN
oDlU/aLgXeG1Lcf7Jh+/hWnAFonqPQqLuLm/ICdOFIYu3nqOOg2rWN8r8v8LPngq
ocnOS7FYxIhDRKlMAahycu9LFG5TSdodY0HbpvCqLNnQyC0BwwpaJVd2XuvcpZNx
AF5GoTvsnyPX7n/OZDGNPSspV2beCBheBS0h9+z3Z/AJBS1cDMPzMHX1R0GYqZ5+
U8Myv7m5HMv9Im+dPaZgOWHwA1L1ElcCoNtrJH44f5MbuQmxhp6TsBg71f+QnjWk
uc1hjoB/85dp0nZcD1uS1KmSFWP0i7oYMDfMaqP2kRHeQgs89uW0yPGwyJ/hA4Fb
REP7WOcClRpxxwwznkKq7i7tzaS0+IN6gz54T7RmY6H5durv0JTuReyD5vA2YG6X
8zkzEXF5bLeagUP6VSr0lJdN/8y9oz/KCy4UN5r8WC+bf0XOHy35DyQljvkB53cb
6eo9aQJNN8pmjrXfdn8tk0egCWS1y3jiQyBFv5xIGTYegomteq4/qbz0bnhA7B/s
wbRUW99HA6yjxQzuSnD/1VgsAeJ4fr3xGDlxW0KtgXBsZfjTgssDZWG59iLfpbHE
PamDMJBJgueBtBjAA2km/tUcIGduCM6Np6WnKe2BxwSAWrEa/CAtfWpD0vbCUCMo
GxPMAzRJmV4hiqKoSWZITT/67jl0pg2qMybyk1LVmDKBUiiThs3UES+kHbtEbkz5
v4hwSsun13AtRii4OReO1H4uA/w1gxPbgIDoyipjWQWv2XYKz7SZFWdBOJt2Shol
Cg631RiD4OpBSVPdR5Uhj1FnqyDzDgWFFIzzu57s0cjs4Ts4nr5B1QfPTlVkf5wT
ej/p48r+2B1vzpqpXd9Kt/tSfA0spOT9o6c5xzeVth1dAuqKuFQ0Fqa6GILClQ/z
jTSYJQBxVldQTepP4025ec/eyuwEZb56pQ8tokyNOV9J6GHR6qd/uDrJyqKz40Oe
`protect END_PROTECTED
