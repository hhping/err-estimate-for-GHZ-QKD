`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0zgYit2BxsRoetVySkkRgdS/ZAp7ZkSgYaGWEHLHM0t0eQuYAZhJ99+RFfxtq5C
zUpHW48EyPTIdVmlMZpDMuOGn7JQhydeHzWLq/LkZiQGq6hpy7mM5xwn+fkOyzPp
FJQ/7yky4OvarMNCTjiv+viLLPGAsuscofeUcBp+/hB/33v2Qv1oYpr4g4wsG6aQ
Qg5x+vIbmbIDPQyrKtjDXQEjVMLK8W6fzASM6rzy+eCLBi9bvxTKgmhT9D8GrNY5
5ml/FSSBq0kzDEVorDcH6sddnXLlioJdHeZcx3Bx7584I/yuM6OPYWTuQgAfgkaL
FKDz4VzybvzLuwiSMidCUtgi44/LWMV9UhqqFYYXY9dBnxtYLFm32Keia6oCY0ay
ZcXpVjSCyv5k9sHANsPj8+mLYUWXGOKm4fkdakS8Y2NNLpewvquivXGPm3AZVi9t
pSgr5veJy2P/v/bUc250rTxcN7lvmylggdQ/5Hn7TMucEZq17IVc6ux7uIcu4JlE
ZJ5HZcNRfnh/ZuizVAJU3iqdCfWHXrionEItxM0u26SwYRJ9TUOlSltjje2+14HY
0bIdoGTwV3CJ2z5ZzljRFj9gfQs+++TTtTq3QfpIL18Bkpsk78ZaltshkdZf2I5U
F5DKKpYBt3pGtEGXjU0djdOwATlxB5bOeJrfydD13bXrvxFyyBfIc/CArbH4R4oH
dC0/oFC9SSF+QStBU/cwr1GCwZPGml6b/JwJ3DvWJnNk8SmcQOBAIoNDM6G5Nm4s
A02P8wWoKDkNYRS1KhiWBIkFuNma0qwrC2UzVK1AKbybUdZVHZx/8N+6NxlfO8QR
tDXi3nylARwSdoh1C7hgnxDja7YvJro71BzMXxesD8MfWHlS56i7zx83kefQJJ9r
mSr5Ph2q898eXP9IIKRyU6Vi/dgoiI+vcH/ki6hvEl4=
`protect END_PROTECTED
