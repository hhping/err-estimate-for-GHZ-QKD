`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQYTEXhwI8CzzgE2XkYwS0581qyTnOwsZNk5Q5otmeE0/ZJevGbU/0UMJAVzG0wx
bAmmzdlANyF/DUxZZv188ODZpqv/i0kHsA5KT7czc6kNk6L7Te9lJsk5JEKQinMo
51QIrMDIZYhZePTq+4OVDVkYjthsNNy0P1vov9NWRxIrGu+AJ1FBIv0Yl6U+jqBT
mjB89y7yRkD+v6vaOwTGXIBLcaOg8D7ZOTxVg1PIesTWAkqJSYmDhI0WpCUQ1Vk7
JvQpIvvfFsMqX0a4P+MKhv0TfhAka1YvdmTIXwHoRwVx1H1M2+C1V3pqHZAG++Xp
iqvWWu+oaoAP4+9vtB7qWtgSNEvdDWYzjTGBTc11xUhgd/Fi/nwp1UNBRE91YcLq
K84iorRE44dU3kQs+HeuYd+R0XZV9XqICWqutItjQcMf5b0oHPahrqiptkHaOVXv
KrCkM7lYrLo+WavvFLifpK5ZQfNdXY2gXXfvFzdGeAk1cJ3X8Au8prv0XJz+WISp
V6+BgO8WNCkiA9159iuRpzxzE/bO0H4aZEAWnOavrf2+nUpVAJRk8XchaFAE4bVI
2L+UVoo/eYoieobS82FGnBCQmoGrqLaxfX6Oycdo77rwbc5ejZqMxJ21w21qf1Mq
c1bVdQ5VpSdjYL5nBLEFNj7kBTl8x9wM/Q/Ri8UdLhwpzHA3pQSVj/dgc9jTTrUM
4WhHSDk7fj3Dfz6jood/boDMBFgr7QkJAG/E1RBTQiOXjXGfktdgvXEb3zcQdoRW
/oQts20dW3RNt1VYSz7jzXjEDEhyS6xId6SepBmCS4OIqojO4X1ST/9jtMfMwYGV
RWpYxEa+zy8ITRUEo0O7gWBWVnc43qNLvnsnHjAbuLW1nlgWEjaUO2QOxJRpbe/3
M0Q6KaGcXpBFwwwVIUITmvM+OuLCjG7EkFgB8YopEbkuUxo33NjD6aGlagukx2GM
9DNAiA6eoJC0K42GmvaCQW3w9/nbKbEn2Hx/ogtwUrIwJdOu9wLoZ6IOD1xU97u9
bcfjlEqESrAg97G6RisKUZekkyxyJ44W4yFT2nlrapPQJCGARiFsNxmHk//phahK
bF4n4XpHh+vDRXgyQcCVfMpBF91msbcDrwPV3K+ZJV0dQan+MK85VhqSzZFJ1Znx
X4HzWbPc8uKpUgho7WFY009NXQUHTi5hd3fxRZ9uVHSIGp6RSxivOxQq1gsOTEYQ
ybR+C11TQswzaheTX7rbYnRNb4rXQ+N8sh4GWxkD2TVFGOafljqUfrlwQ85TdjSk
BVTZxkascpWGTwBez5bRUB94wyoUf6TZoKTREmUfd0EpE3PlpMS7IoT0Zc0wLwMi
HETaKEfNaV4Q7AcQ99ykxiNAF8tx6+E64v6yyITB12oJOovgGUyQXDD+DtDTI6KH
a2bJUU4MjpvMDDgRI5l/kL/eH4iLY8TRENfKeUcFcz4TuSyV8BHsPTdObzCfRUNX
tsqN5KTrQBM15eeHhDALi64CYwWunUydZVsv69zlFZOO0hKpS1HF7x2OOjCu6p4Q
c3S9dVjjmaRDKWN3WKOhu3fKXutFMsEstAmc31w9BbXrY418Eu1G7CQJW43TZf+m
hbJ5RYmfGX4c+2IHGFLylmUNbdG9EIokBNEHhKwSPMKRNjyygn91JBBmGgsQbBDA
wXA2fBCLN1X8SV8ZMqn296kSWsUjl0loJDPVy5kGbNhRjeSVxGqOvRhWhonSY+XC
4xJ7YjD/NC1Tf81hQu25W5Kir1asHzZgOG2Nir8JV+25cCXUdWvl87+4AsM1ossx
LTb+Dq1vL0uSfDWDY8b/ieU9v8cgHYqi1LGn21njibDrCiHtR1YKx8pOGs/jidMx
TAhFepSmZ3JMZnrv4sT9K4RWmfxm/xiNAFUuegkE8ne8nwerIM3ACl3Z4t4nsQxV
FEfefwrt6vHDCKVwTECfp5T10QMlyUMZ9DmiBHKnf9njoBSwThm6yVAnkjWJI2N3
zUwZWI3VTb88dNqhcDboA3hFWEOuH3h/I7EVF/mE7L3bu+BZbDPVB5ppuQPcghqi
oPFhSaB6jBTCagNkCYK5z2NxI4TaV/DmPRbtjgog4SEIAirU3crBxpK9vPd//1Ys
`protect END_PROTECTED
