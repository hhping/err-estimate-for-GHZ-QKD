`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eHcW+DRBjLTwyxQ0Mt7rB2W7oVRjsoLUo1r5BTKehDbb7JocNUAc5+P3K+FVy0Y
hPjFWV026gG6EwvTcfuWSPbovckgbZ3Ls7VX5ILVuutZw6mmGT5L5JOcZlt6iwIE
SsKEJKER2qIwTvqDghLNgsO3slzZjdiA+vVeiGqb2gvaU/GbeMO8W+rEnNNEhQNW
O/fqgq6vhaKdmtsCqRMQw6hqq3CsXHo7s53vqFfDPUslD8cAhtGceMxbPJo+MjOD
tXV+zn/hYGzGwMupUk70lYc6EvC7uR21mCHN+FbLIh5QJv0WSKzNVCc6R5SWU0By
3mhNflAWdyhTVsO5K6x9xM7+vfbJvtyITzPYJBEXplvu5NBtHfFneCGWZ7z4igIX
MXiXQhe4yrMH1QCZg3jKXQdYcPACWHg6xBAXL9IAFrkKgc4WLI+/tOEtuMApBMrZ
ABN6kifJuqRcsGx6iHHteg==
`protect END_PROTECTED
