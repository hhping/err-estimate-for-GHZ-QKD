`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUt1D6x3A3jzwWsqbpaRRXYPQF8gjeV0jI8h0nDZfausgHFXoz6Kqya+pssFOAe7
VvrP+xXYGH1rcXIqh636EkSUg+SXcrxOF5PMsihLhHEG9NIe/4TUw3xJS2aoiclH
n0DydLw7UkpW8H7dCaCHSdxz6Qo+P26NJ6gO0SayxjrL45dmjZtnwpz4Jk6zxyYm
gmzw4fiAHKOccobgHJzCHPij5gZtXquxkySWgtY6oZeYBACVd8njIY4s7PZtlxzF
3tn4lCOpZV3Dq8+YoDrIpc0hgDu8apjgKp3gOdrw9oRfXMhBAOpMF9XadrnBJKb/
GLZ7uKnCsX7RBw02uHi3qFmQ8ent9xb0evrSF0hxVcPerrm4jR7TeVcsKksHim0r
zNvjyV2jxjiRyf9B5w8jKMMVqlMzQBi77WxxKPchtQQCUZ23qNAJTSZ/lQNr5lxm
PLB2uPb6eNcQuWwOkTDvddaHwXAfReG0GO151vEwQ1fE7vrhv1UOS10p+w67JhQm
ncaNnPgRfSVyGRxUvE60GOe5he9hjWC+jpcDf9N0CKESKoMprVdPA1Xiba/K/Hic
3eQq2SGNZRGtptPeBPrIZCKbOTs/pUIDi/Hjr3cUTwmMnNfm9F8B8ADhK9sCKpVx
wHNXqI7c+ZnO79Z6SFszfUBUm8LGVelMUD+5WbTH5fW8mnuJySCj/b26WhJnxj9m
1xnuS3zfmPDvQiNfvL/W+MexzxbXouFuLTcDPTH8kNYkFEtmgIZMXnFpdhte6Rla
Fjk3ObgO4WQhkuPXYtMr4JGXMQIFECg6ypLyprCGsATKWTvPfb3u/Z2x3igPFqoH
C0rt7FrhhGdtw3EvPBNZI0XwPn9raWrjRq7bSKLZ4erV6RyzMum2uK+quB90YA8w
JVKeM1b4NKRBFZz93Q2j8Cw6jaXzODSk+pRamwCgH0V2AZwcQ+FkydFQG8BQfKvI
xVoyEM0BaQnRVbUFm5sQev1NKyVw0ycfndrQw1C/THoe3IsoZR1BlibVRWz/LuU1
9lKhRhsYu6WkcQEUgqvntKE82EvCsckTL35oW2DynDUDCywvij0fFOcpVPt61FkV
PXRWdBCcQVEMKOVhzR8SsmOFfbJyGU1ofCyvcslgPd+5LQfi2otZ7spRNhAOQVir
dX04EOYaTxbZuda0QlNjAyhyaJZpdjyGA9SQnC2OFrgmyt7t1vS1zhtC+DTnmG3g
PkW+TLYrTsIEzDDcRVm3KBTKqYWuh2yceUQiCz+kyRy31N6ekUbzKSWXuqAJz4VP
9zJPruXTd9Yz/e7Th0GydA5EJRYp5CpgwSzqNN6wzmbpi1Sbfn47SCIYmhjr1lTE
CLXw8y/SAwGsxJa357KGAoswrOG0cDx79gjny9dHzvmMecGx0h+ilOo2e8xa0Byh
4S4a9N9Zy7e26ubIya7+fMMiDwYtHvwPXho1pG5k8BdxyVhH0c5GBc1BqXaXA4NQ
MgafKJuy1Ut+S3whdFpCCJngwLlDr5AKi6K4hnbQ712ilPRilYN0jNz8bUP6tYtS
uA3/WmxwACNIgPeR1pG0ZJX/jktJgBnO389o/ferIY4f/cKdac4Jfu1XfafCq9OH
XR1bv92PGfpXNZ1ioNkkOKKsJ3Coi0svi/7oXdPY5fGrTpLhss6ES6xowxvLs4y5
0NrHfai08dqlSYpoltzuWWpT+cs+X2kAnhIqAE6ToKETPnzjY0BWqNs5hmblY662
ytGGj4MQjOyq2Ol3X1vFG7/Hv8CWTN9jD7vnexlewe4mhgkayb/eR8sb7S0KG3qf
M8mE6E0IMqYvgJUC76E3POUhPGdnEjFajM8uwIhDL8j1AOsqXMNnCChclCzt+Mwh
ovcD1INkvvvSe01gZU/g4na50dOIitAmyIeciYjcyzsJZnRUyp98oq/Hi1Yqm1bU
LUviD86ffMnkGd6v8PeM2ssVz0rhCsWna6UrwCXDPvcATunFGVLMndlYZyEk1fUE
V79i+lE9QC+VQGdVNqDeM8Wmx06IrB5gfcGvIsg9yH4=
`protect END_PROTECTED
