`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6MgTM9qV6SvaPnNX0PeH0Ta/6dfnAGzyow28R6CVR29BT7v92DPShV4KSSbqpAy1
LGP3FvyOPP9QWuFA1jM7tsldeKPD1iGhPhtrPU7SdMn6gF8o7G3ZLCBBIftx3BmU
Y7rvb/SDPKrrQVUkpobzLYci0wlaxY/TdvzlSIR1EPh5Tp5xWGk+P1YdwYn4tLlF
FLbOUHUzbaqNVY0qmjKGBwHqlAv7rHytGYm2hiFi3TpIrIy/9u9hl99ITglP7wG7
tps5Qyt4PlyRS0EaIWwp17kJS2AxM11Go9rNWH45sJsdArL7mi45zxJSxsD3sSfY
AYI+K02TdFn0Fcu2JLLXJo49OowFsOByGBmhYPyYmSeptdDlneX0XfHDe/oyuCxL
hzQmvB6DI4LZgCIGeLGpq8QsYrNsakpoBJBZvU3Fe9e/TnWyX58jnMBIC61r3b2a
Y7BxtryegzqCcq14lS92+2kpi7NZz6OJEs3ohqaWXu8wu2wvPS7fbNCZcXlKW3h6
fcApQliqfPr7iMUs+ekj3sQvB9ixXuqn6gOlGuAm6dE5CyS0aM23Kok+Hl9oOzTE
NiE2b5y/SDtb21BiSDO9NcRDxZysLucCnnKjdWFsYSl2ZFJxLMVGlhWndmMj1Go5
qC5QkrNT6rVjpFDxfhuRv5Wn7bmqGPukFwSMCaARhgqz73VtqE0mke4QgxeMW3dC
6zT36lFyShjNqrNMnSiLISKoLDRINIGphObhlXCLl5avttr9DRSZtqqC3yfmUsoy
QzwItLBTsEV2+PN1pZYEV6YVN94Ux6aw2PzOMlZHZl0q9q5rFkkytAxog0Xbzco/
gYTlZFNn6NdytTfIHNNCCeiRYcUdB9MGMng5tjD437tkWr68i0pKMG8EvsLjdj9G
uTIultJ38ozg2RBWNnviZ3ziVN60AoFU1LiXDdKu4AT1Uh598lARQTV/fYdy6TEc
kSHEuUZtEL7z/vilxnloYflYudAs2kqj7PJwGYXFKWTqLicRRRo6oYu2gFmshPvZ
iiUCSsYgeIa6Y4tkUEUvtQ7Pcf9uw0OsWJ3VT7TkWLoFcq3EbTiQ3FW//YBE1ZJW
8tPOhg6rH91g3P//jzE/GiGTpcDj1Mu1MEhDCUGWYB7r7RfnNR79vceBxWwS9x4q
QwVH+1mikE6wHoR68uxY3gXguvZQBY1rTM++l6B7ScV7f2C3dkDSGG0chwCiKsgF
2BI5pCFl6Xy4bJVTsM6Ceg7Q8t+TKtyO3BD+yOKcUjG2GcCNX8/L4wkkG6Kn94QT
tHnX2aeaQdF9kyeyfGGOQWpuMhTbYrCkyipPFvRM7afcA6XdENi+CUY6q+hbZ0BP
a+bc+RRbaibY2+geovJw7fyruUv/uHQOxeUuQJwrmtqY/yiqEyEWTLcXYBkh9Xic
zCYB6fLxBjnMpkIkiOO8swDrqbcy6v6e/QAylCY70gLBUC02hs9V1MRZEyfz1uRq
t98n4GnXmNwVMkROvo8D1rAS8u+JPrwMdFMUOwY60+OuEVhhNpRlyJHIxrKMmH4g
vlYS1ZpwqKTNizbRSpRZqV57Q7faQCxjeaCa2kat1k8J/Kk16T5bRIKNQOEf6i48
G5ocfG0tWu+v+JKRO+w/E+8q+rKycowHOhFJkHfikFRhXBwgoZkKjq/Y+Op0cPE5
cvvnLC63WNwIxckxSo2idmJCYX8MLUfs+EtchnXR53GI7YaEEJaEAhJkMxmUHeqY
HegbHjr6ViEF3tIhk/H0OaWz0pHRyuaa4mdA4hrKFH9p/9vddox5cIEJUqPQRHU5
rJKvXpSOGA8Memt2WHqdFBljhiSp8HzN4KI1V1N18knQTgHwPjzTphvxsbFW/bIP
/5sIAsDFVFVvwpQs4IugbEmmd/QPiNh8n5h6pZujdb4gJ/51GoTyToD5eP02/KTT
QDyarZk1NsgFighDJU2FUhAgrB6ucwqJn7kDBXRRU3WQq8qGz7cxz+er8WrsOIOi
QFCQVlOsBUzYEwY11rm/uR/2BbSJc/vIYEAb2tqkO2EAM1/Op2kZGoRBP9nSLeoC
3y03YI+r+sOILIq+Rk901doIdcsFXvzzI4Ij9UCRrBWvGKQag9bgwDCetdKYj2Yg
m5emnzuvK5Lsb7XoqZDfZOrCIcMeDJzRzneWx1L2MpwoRFU2REk+0RbwlFkYoIu0
RAEmD1wEmt5pFFeP9BE5kze8eIJmyPwscjI30XXqHuS2u9PdoFmM/Hn4YOXmHQ3v
uV8xy1C4XqLiru9DM4X93yRMVWBF7VWERMAioVrFT0Usao2zY0/wwIptoOmtEoSR
C0DwwxWRypq6WDZx4wiR4P6wqi8qp1XCIhTSj77JoLpnhZ8DTir45beROyxKwKlt
7P1qLQ59CK+3h8CfSfRxGiQIPlDZlCj49nnYH1UAsPWM9gCab2YUCRnO1joWIWVl
ANgrW6pagtqqJSt9ZwFjDFXkzR2iNI+E0dh50iLJuqdBDiXXgkn1C5DAt/50XYg5
AZb8zMKHmHuRcnKIHCUi4L577L+skj5gdLQAxOffNUvlDdfBzOg27TeoVdul6t1y
/vIVa9kLbQsxbrtSO8Q1OZ0wNMqFbz+hADrF7Z0G0O+1MSnYg1HGjXJJabmT4WNz
cT9DOw5g2+b+Vk+K24ZcUANL0g0XgrUUztC0LYDwBTC4FKPsyNJkME/WYqry1wYs
cSF7W1rRLfEcLWg9SNK1tw==
`protect END_PROTECTED
