`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUnsRDUW8MOZjgL2BgtZ4PYyYsYSniuGOc3psCZYPS4oSsSSkKj5Edf214JUGzcu
0VuqqRuYsvaNT5VKx8euNpUsKL8+yIQPKoLdHnZsdrX0rL3RHEzzeS6wjh94Hygd
jELjdQKKdqEcZ4Rza1BrxgGQvF+yCBIxHl+BnDNd4HqPlgnrYvdAURSY1K3/ysdh
zLRfOAwq5Zed+0W+fwOorc9jtdskfe08HLRRlQpdvwi933oO6UBxdTEXVZE1J91Z
VxgzQzAe8t2sxfzHpxBjQDj8fouB9bSusGuS3R9TKgpUzKQzFraVV82Q4D7tgpdR
uJz3BjWK4rZM62+IYtPBgcKfjvK1JExZ02CPHK68W2TY03uxmO0zwkJ9sVVoeCX9
QqJ+ZMSVGgY0gdIZXTqop3RL1rgSOEP9CzNK9qdbmTXr6OgUacgHLWhbU9644x7e
3HGY4vsNPmympMUOKF3Nk6ZEA/Xy9L6UpMVphvQ/wZjGv0O5hCmXYFymeXACsx98
FQxxGrJKUgLUUdz3YXh4yg1dg36CYSXnSfT3A2jqmFeqls0hOKL0l5vIf9DljUlh
EBG84Ox0HdsH8QaM0VUEHo9F5gYjmjinPaNFab/iqNr+NX1/GpRuFm5YVOpOxgQc
rymV4rETWT8HxvSbigBPNlhGhyEFSYtERIwKU/PB0nulgwctS5PBioHCT3ryYSmi
XBD5kJhfbESTuWxnZvRAB/intqyXON/e6PUQesBcT8slXnd+uPE4zi5WUsEHiAI7
vELOtszTnqBB1nr2wr8PqeE3SdA6PTrUC3gyMoWFmy4eTleHg68GVNLb6AzMF4M2
eo2bhjoUrGJKahLW0kDYtf5wMQC7xdvLGRKCH8SZ0tdnTBjM5eyFlsninuBmJFTJ
4Wu+NvXG+scuogVpZOBG8n5j+gImu5IhdLSu7JsgLRjJTZvBUhGz3w2PmScQKD0N
LU9FEtyGDnD6zNHt2OiGs6fLUDxMcocKEXUbg0HKdzpwMv2f/M/DvxZU/brhJxHO
n54AxqGJ+iRby5dNLLGcpVYOlUe3H5mEMlu3VIwT1fLATEDAvKoed0rnpPLYW0YP
TXDCCLpaPOX+sP0UjSTcHllKPreBPIoJtTsu3l1SfX3P1CUiGPJy42sT9gXBQ0iC
1iQF0s0mv2yp8GIOVTwy8YRAdJdc5F6v+QSmqWxJgmoBFFiGB0zI9nXJOosmAhUn
HLyNESsour2njRY8+H1l+XLwDgEt9vibwzVFW6t8P4LvgfE1LE+Pp+EBlNOBDwPZ
Yh3oPBN8DvrMZCrVTe5ipOAgp+S88vGhJG57ZTiD8sbFRxj9+pfvkHjcpRuOqelz
xK5t0sUm7ddmULwmbaP43i5BTEnVShnn50BbbjWkIKpGEik/vkTstQnpQoocVN0X
0Qg4nh5DBpUfjX1WbaIJwgFJaHx0V88xj4Pc66JlormKpyn4M83Mf/kqa919VIqY
fTd/bP1wpa4uzsP3KuRplDNyrvkoyphfWAUalzoOl9HcQIextbTtBHe/MIDsbhBO
FKX9V67cGsaoRPG7jnNh6NkdVtqnpbsAWaa1W+KpS7ftYhC2/TbQ0zOgDEGiP+DZ
dGxPhiOC2bacxPNjObglio26/t1G/ptKJuEU2HMg91GKitq4H2bbf9EJEn7sZ6Pl
5eEyb/MC4pNKTZw8gnRFOjSU17+VtnAFCuBeL2tEiZ8xbSzX5RoAaHz1gSJ+6esG
0b/bkFVvTmS4sAzTvvgwGgTxfu1upep4TdxcAfeIszJfMz91AGpNjIGqurWSs6dH
LFfqV3QTCdx75rdkoK3xx44wdE6AgSnIqE1BObCavWMyrGah/CBADIMyJjADDpZf
CdSUsT8MXY3X4EQp0Z1mE4xvf9d0oUb77waiW5ewDpjKGTFV+lJBLjaxuf8Sfkxg
vjiCMeLKGjuekJPMZxt9tST/kVKzAf9Qu69CTvhpJlS7wji/76UFpl/fCVFk+axZ
Q5op375SBpbbBz1/aYrPsWd8wNRfe5Z0Yamq2vCkvpLeup2vV8WvV3aGieXgMmOi
IK/6zthzO07St8NvJ3Aa4Rhc9mVJmmQb9P3p9OKOzf756srAFjmEw2yy6LsQ/HSz
R5yB5ycmniGW+h5i31NT6BMb/Rwo+2D8MrFP5nxT8LRu3gWBJWRje94lWwJ3xyP0
12pFGY++yJMP0aLkI5Azn6PYFG7hXF5NFrkehcHQsD2x7FHM52SebifsN3z76hun
qV0dThJNSr/CBqkVr262+iA4mBbcgpt9/VegkuWMeccKMWd3BKYinGaL4epZyLbO
qc8AD0pNczExEY7Ci6JE04G6qvOAbDk3jCRSC24ToUSdmiMPVrXe/W7b9aJfs26L
yXfWR0ggwXX20uE5VnCQpdBBcLC1WgAksRUZ3EAFiiGf5IXHDPTR7b7IoFKeYDIx
3Mc8FsS5Ee64hpD0etHYR6iHgasBjP3H+vtyy9fEQ/rkKnyIJOtZvv34Tr+Kl8YQ
mWpPqCi8xu5AOblSpHk3tOJ8inTJsB/lBCcTeIbJt/R+w9AEv46n4kXSzta51g3Q
sPyy/xBUaGDlbI2AWE6Cui6EHopyYEERcOTtUCE5lmg2AWXiZDRumvTZDx7zoIoz
RcgVtzDti63c0mEanNcdbC72rTLQlhFQjAT0pcdGjxswk50LEbpwHZ+JP4VCyTzJ
xXuRPI0vIidNRdjedLM855KWa5yFRG2f7diFPLlJVZLJeIgezhKxXb4uq0UEByUj
uY+F37hV2C9HkSZLKU+lRZfjXa5jnfHCRW+KwWPhHXA9cU43D+kNVF2ODAS02vHp
+8toRJAjnVDXh4yR84cMZiuxwp6Won+7zXkIjLFI0N1jao4HpN5rELB5pGzmvhP2
BgQshmG3e9Ct//7MBSwlPF/fvejgJ/Ye6JuaJQofdazqfrh4C6wh/6wZ4aJart+D
JcBbvEPuE1gfyUCtBw1bqGOWbKZIM8raIkTPu50yUVvfiOQMqJDTSGgemX5qwWPF
v/Gqzp3RL2YlVr8AmlFWzT6XYznlA2Y9jcY1esboh/UzEZj4ua9EoTAt8n09QzrP
/Gm9+v6Bv473wcodCT9gWdo8hRDSMMJsJWzYnCos7VDN0NAO424MPZycyPJnTN5Y
nfLhKZGZr38SNSBONVtS++o8RiXgdQkBwRp3jI1DfjA8lBI/Cg+XMFSSXteitpO9
Y9vo8HJ0m+nfiO/bs7I7GdelzmwXvbzFEUgtWgMTZKbezeB4EjiufubKnZMyOo0W
AIK3YOdXlJTW/T5qXkis9am/cpjylNF2lLTsPaqxB5kwUhhYbtGl2k7bbW4vYNoN
XYhAVJlfwHTZNyuf5Tltw1CLHMrnrGy9yegsB0p0yF5yLGJfoyxYz2AaYb6eiYQd
WrzpKuht8DqHuGiMn7RYbasGqn/tZ9UfsNcev0VHKXTYT8ZdhZIObPU/S+lv5djb
5g02FMtaGCrBjE9Sx5Zu29hLRCqw77i77QW5I0fj1q56+n94ONM/3oSzgv7ejkqN
wGAlepnFL1xZUE4etqZws9sJEb7tpLi4gQrSOD9sPa5kjOKE8Uawl6ISMR2ZLFli
nb7hmfN6ud7pjyce55vGe2xx+3MunvbyjjADDFPObR4/lyJrIM2rbxnr0kxYQOgz
HnHUUufAEaV1DJ6MlnKGnpuaMUbS4ey69cWCyIhDmVrnqa4QG5XJ+XHt2E+PC+im
BHZahGEQzsQeYUYyClgU6zGMNQJ6y8NgLwwt2kHWCxhVE0JOAXt60ZJ2uXfQh6jo
Qg3L/i3DblG88dOQFYdRkkoaXcn7Z6CbGRCLhoFkrUc/w2B1SPj9ic/95idO/H6H
aE3pm+/6Num+jjKch5HywBwZt2zVkbCcA0G0i7HvQRXgdjkTdAg7AanSQhbRK77h
LBPwqGx16UM+uftfpT6o/vDoQowaHD7ynl1cVceYepsF7WVqN2qUkDtcCmYXjZBa
KHuzRk1Y8KQPgm9IwbLDeO+wCbaWQBpRw6PFl/wUZyIKn+oIt1/RR7GKfU2Zv9j1
1TwzDaPRm7/W+qzsaDTV1KwwBCAtLG4KYGGCLlGlxY7hJ+Fc0FYs3JKTpJ9DjJXS
YC/XoDEenE9UVP24jYUPMHUn5/1o0rGUmel1i7QU+favmZxsl533bIcZiDVjQJLn
5gesBFJkXutl1hhJW+F2OXht6wxDR9QhyCTcZpnBluUXcUAEIHVTe0LvfQliYBKT
2DwI9tdij9s1h0ZAcdmWLk1PQAVJWQDS3gGtaiWLt123L1ZbmzGfrCh8T3QaETUC
a1MflineDOXXanKElqLIcvCl10IIEdJspliVxodbnwYUFauvw+tWZhAAyxr0DppD
JfxA3N1cq92ocFv7fg5D+2E+ggOV3BB/eKHarQuVXEpWHp+ubfCz5AMkiRRB4EHK
NNbhhF9xOAhCWbA2FzfAPGsr/U1kiCY4R1v7zumo8x7cJ3xdWUxpNDVZ9snO1msy
07pRhXLA6EeeKS85SmlaQ1Rg3RAO7nI3X7/Ce+kmTIALzUPn6s7neXoaXVhecXM/
Z4Z+FjOVgyYX67+sMn09aMWOTXQzpdRXIBsNmUsiT9ks5NH0s3PnyWwshaFWilJ6
c9JQtR7FFczsW0kbWr2RuSk6yQs8nS2uUnVf4R/yVLP25yGTRlziQtA0JWg0gJkn
weyACnrgHn9BvE0NaBcocXc3/rzLsBFbR7Rwhs2Hr85W3fQyaFb9gR7xLm/ZUrS1
S0WxuDZjpGwFdT+ZAMDZ5ZDoJK/36lsb3zHqvaLNenERLDN0KwBCe34VdvFurVbi
A2XLiWcPYfSi3PHyZNRkJqGjapcoBpQ2JjMoCCtrHIeL6FPE20HI3YTFIf7NKz5O
dHzyQbhKRGz4J7BzFT0Jx06evj3kkf2N3TKPwq5EKqAHS4ouNlNjtZxMel6qvxwQ
S+CUZ+VyGVg9s+l0POCBMjuzMP2SK8IzBnaQeo0EOEkLInQlF2GPxGrY8mVN02en
GFyc5KUWqx5sS0rMYC65eqhhsmxZJJ4LruA0M7Zfl1c2XDm+PHDG32cWpGyx+L+8
E1VKwyXx6mmK5X37bK+519WuujzmxvIPAJj5b1Kq23ckR3011+Mmcvv9xO1B/JnN
nzfrWHePrnLC4V/0F4rTJR35MF5fuLKiAiLTzNh6lWIqFWDyvvvsLWrA1kxoQgxG
/acJD9dEIhrL2JxVL4okYDXDnrcGSiC64ihkfkTFhuU88HstpgyJkXmBqpDwQs6y
FiM8Dxxt8lkcHWm6K1LeRcCymWnTvhOoEWAD6cqjnYkrMrzA8KhzevzcFFed3xlv
G7Hxhceau8tBrospId2S5bNb/AQWEhBzVYYby/jxN39qeqbaQeIFHlSzOv7UowYw
+lrkbxzT1hG+t4P9GuofWAL+5FtGqOI3vqEulvkJmZora0ADt42Efxz5E1/3UfHE
8YwYK84s3aDy9+VmysZDTAbOTfvBJafCtcshvwXaahuhchiw9gaykTC+SM0MA3A6
0/x2pdSDd39+Mg8bDe4L2p1iPELuZ7s2KYUabe0MUQbRsxsjN1UPsuA2rl4KANqX
MvNiZLeWKlc09KTG73G6mfeWKdVkrWSqK4rqhFVZ0W4reyuhec75lCEDbiiLLibP
hAI2/6NiWvzbnEaTRcer7bMXFHtr1whHjDhBAA4otV2r+czFZXRQNwKR1Rh1hhbp
t5D9cHE3WDQEUO7WcAea7fs53fyt6qEiwZtbfUoimgtdw/EekhKuUygnCAvQi+AA
MhB9MJBlLHTLU/UMfg3DVBFC+gk5VJ6E0qwAGElypVBKAeF/jdmscRVHw2DCNWwD
ypxxwFDY8mrHciz7WQmkUmLptjBWgOPbrO3dQKEqDRCmRIJ5P4wfVzkhFiDcW8tD
htKY1ZqvmG2ycrjoUxkYi5z0EOwJxWdygBsThUO7NeZ7jKf/qSwR49SLTt39TYcH
X4IuG/xeLPYEyOBPaT975OQHPCIu1jM6wgPLOJQippiwLkK4FQ0x2nY6REOrq4sp
xKLZCr8lZYcwSMnaELvlvB4VKMpO42h0txBu12N6tUeDDHqbgztr7nBrCots5yB+
vEPgemsDMJzCgnyCtcBG7zq0l9qsVkYF48aylMqSszemdnTPcIuiYmliEvF8NVV1
AqDgZL+FRO0lBCo288d/Bz9GufsNkSEC+j4E0GrECA/NIWBz2y4yo+cW2zZn6npg
Cu3Ug7+p/3tAevZs5829tOXdx4TDrABigg6BL7VF4Z1rZ2nOO/i+a4qc0oPlwUqb
0p0pju4+drOfcp0o07b9VIS+qFQX8nzrhCQ22lJYaCnMBYryejE8Zdt79hkyul7O
/zyXAwZ+DE4bKNMIlfk+G5TYijAvOMfRrZYmq/TQJjIPfry142xgefJjqA5aIBSP
thmNydXWgC02d5RBJr5nh4By/Nyf2p6FAXw6GTwelbhbKF8NMHfaOhpjEf1U2v6N
6+eGpEmrnaOunhLsXD323OBu8jLqUxrMGZgX5AsJF7rABikUu3/15r5uELoAfcHq
dMR/zJJnNOEmzAsjamvINnmEw3nTrSJaFht9oNFd2NZA04oHHGaBSkWe6rk+HRjR
ul+28toD98m4PexBQNSe6tgbdLxFWtSuk3MNTsmP3ccEsZpuAM8CDjtgXbR/3mnL
VgyuCbtQYrXACgKVZngnz+vINu1pXA4W9n8OA2w3+7u4Rg979zQ+ScIUrdrG1Ig6
OlvG8K7xrQ/0OBeYQ+CwTVBohcz1CI+nG3s98aLXKqA4K7iEXVYFhob7ee60cjZZ
xQq62B/Tx6c2n/0goX0ENwJdRi+zepCJioLLVccfHVkwMIdWYxAgcnOBVn3+UM/m
7jFFyk4VrHrgJfg+W7tFtwimVMlfzh7fXa1nlV7gFJJ0SvJkqGht9CCPDFkEpA2m
V/VktOC8Cj96XS16QQS+W3fNDlAFGEYKWCaR/qdGK6EobKz70YEkcWl8FGfm2Hk0
RfHB2U3jPFZWKg77yyOHUltFMLvEIv56JD1t28qpaxfOVIOTjL9/x3r6WwjgoMCJ
Yawm2jxkR1qq/8rpSgk+7g==
`protect END_PROTECTED
