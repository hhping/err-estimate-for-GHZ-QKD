`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUO7MqQ6plbJbjC7yWHxk3jx1RIQ4K6DWZbVyhN1/OvY5Exa3wa01bmSK82ogHa/
YF83Zy2clgLXKnZ48LazXebRgqAaQDOWIhrfxEH8H7H8fv22MZ7CYGOA9OehBzwO
38NrFjNLitrVaqBDqi4CCk3FopNJSXmyzRjrJhqT1N39avAM+saksVfzA7PJzBna
Zuk6ZnPsd86Gvx1tq1KkTyHcCw4qOXmCiRIIqzHM+/8pVvm6e/9FpB017ep47pQ9
+ZD26paDFuiif3vEBw1H2up/VeSF7ta9aEu/nYUl9u7vosSPsfmBxzU9g767WrID
Ps5Kpz/Z1nQE4+pmcgsSW2Z78RsHxFJfTFW2A2yR49NzRFPh7/Oj2CSbA4WbmQOP
M3uKlwQffP9Dd+NvIU6iW5Y7UA8C6BZcPHQVFPzXGQYH8CDQJqwVXUnVtAWAIP86
151jXf45FQyK+2IDufRaFvjBWhkKzcAPYp9co4rOd2n7QjtZxKe8N3GYqn+NU4OJ
O/wAWXAbpcIAZ9PQ9gURzg==
`protect END_PROTECTED
