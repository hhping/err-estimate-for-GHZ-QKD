`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gu9rIFW2sCjtWmVluRtrIQXgTv5cG8lrmy116N9PYQPkEUrJcp8PZswdqsn405pa
08k8Q9iH5BCQAJ6aHxRJQR2iRvUf07ykDA4iryYQxg7sodQ2HqjK7fKb5lQWTZNe
vVIMnyGXrFk7Ld8ri3QT/1I6wpRF2Yxbn5RheiRmTiaSFa4dkVJtl4EZeI28w4ey
ZiaGi+N6bGLz02dAGuObAfNz6GP0bLed5elk7O+M326CgROw61DSUL3OcYZOynPV
elpO8l8FkPo+isBEYYdKuwb9YFTVpiRCRLC1X2KxmjStCAX4k+QDm5QrlBJNIQTj
bmUDMaf9j4ucLfCHJNFgveb5ANLltQRuQu9hes+4VmXeCNmXijlFiR31ZmQvVZsJ
sJr3HIG0AQjk7Wv54yjggkt2+9s0IsMCwyjWsmzNzxuw1T9Sb9RKQfLcox5UQeFm
wPJWnr61pACEkuU2/z/YyppMNRUxD9tphi7xKQVXAblA+2fDumxmIpJphyR/+GxI
q2ZZFlNTxnIIxDRlfh+iOoIVbbTUCn14iZlw3VzUCC0khhNeqWyqfKPMddo5/jui
weRMyJlaLgYWNJHN5v0pe/dt/cx+H034/BhtlSza+8KPMwDF9bz2fqVOIXV0GfW8
o25Lk/uVQSetd3XT/cYrryuojE3gjcQFldTZTB3ltF3TacevRqYIRaIqWWKetnMJ
gLU2pMClK01mU6DNpdnydEbkGYXQJw5vL4pGZA2MKxXgy6MXSfEDPqFEaV96xE5d
ekXt1n9jMWHWGUkwANuGWd3prAGfOKPHeH4LCziJuClHvoUZy9Bo7E/I8nm7na14
mgaR0LrdDZto92WuV+kaRwb/gVIBk3lYY5VHp0rLYDt0q2K+8UiZe+cUw6iHSnzF
XBMO1PKzvU4iB0g2nbJbDuFb+jKw5qFC5Ep0wN0DuzodUVVKhpnJOlBrni9Y+5Yp
opuAyVnVh0Er+gVxf8Kr/JJr6tmS8RyKNqllywcnMMxsWt9DWED0Hfbd2vyQza3C
YdZo6Ogjqdx3qk5ZcK9i1HnuBnwVp+ab2YFWQtvIvvLCXr083B46pbOnNltBOKUk
BnIFn15kjqWhQTxXSQz0GHfvrpSYP5bc3Qzjb+DIoXUy7x8MjXSs4MRSzMmEUUdH
MWGCQCFAdNnUh4FRNzfZaaTISFcAJFFNG8YQXHeYJfg6e5WKUfA1qgCcEe4Bunr5
jkmX2vkdbknDtypejfSsajLXCR954DKsE49Ls1VTDqOoLM0dn6Ds78D/kkyVCuCf
dSNEv2FBvcmad23z6v9aGgmV2bmZdoBb+LdIZct51TsU6N2pYRHXjrRNp6ck5w+8
AgKxKHdpGrbE/i4P4IdzNYqiKiQbTQtvLCWI4DY1heZRN97QhYfG0Ft77bh4BKsC
wQwkLw0GKpHT+XNxpVce0gn4zLdLwFpXejI+Bjo/V9ccmyXLllhILPCjzjU1j78F
lpiV8ayx2FsUAE9q80zUVUHrf5Yz60Z7OUeJLTdMHzDhMTsRtrW7M7OTOLk0Y769
hqyFQ7DtkOgsSjymUD/785bVM+qoFu++G8Wh5+bGfXIW6FjHoaIH9ebvldDBJCyD
z0jlU1U4aaJrL2In1SIENqHJUr/MeS6uHaFEebVPpaKuuQFTvhCphJ/jNqhJrO+5
woEgOKPVJ748brgVQiRBXGR2Yu6cHNDS7TJYnpmjeUn0P3ggfFUk0yXpMj71Mj2D
I0EsvcFDUOoDZw5CHWstsYe814sNGGeyl4jxJiCfJNnoi0jZyyVXrX5WT9XixBjI
v0xNGIWImhEFA59CS0M/LsECf705i0qCiJuiQYrNZUxJ3LiIWUpRRtQ9M92vp//Q
/ee76+gCA6001ipH93isABv1W0YCEa29WW6T044oRg4YeQhV6bPepTL7fRlAm9Dx
gGvWi28zsG3gRBaC17DCCg6GB4P7mmXhoO6N77LyOD03dPCnfOZoQTYbPks7uLOk
GS0l5I9cYPq0CTAQCIwmwg3S/qtARmxVls23n7tW/sHwJK+TYZ2wXp3azzinVSif
x2aDIHhNacMco4Sy6O63c9zs0JrQmL7GfbuJkyYUh1+1r7AgG9KgKWsTUbXHN5Z7
rnP8GE1BLsB2q9/ibtftNE+MUaYOMQGrkRzhH+G2v0QaUrIYNL8aQZd5iALM6ZFT
B6DIJ7qvBubDKBRkU2cDe7mBJdXHoBJecBbR2xMNynxPZICEkoXZDYyKO18eEN7X
dtzQgBYNCpgup8y15f/GgZlttd4dmjzUfCFZil6tbkiqen5nyoY7Bk0gmNoVP0B1
dc+a2xHRS+kZwikzK36V18b4uTQ37GSUh7hmXQhxNj+XDidPckg6U51zJSc1vTh6
dGYkDXfNF+80kxezq8HX1K6ZE3sHhYE3gnMv/3Vw9I51fyj5U4Na2Rp3YTRRb61p
WNd9A6QaCkCgIZ3p8HnBJUk5rXCP+GKUKygzr3fxh/F8x6OXCPJK3Fi9WArbX4ls
HJRyoStnFV7aT5lGhJIl7bxi8NcUhpxRtPUxj1vfvB0A21whnpm9chEAwzkEKlTf
6OdTb7nuvCAyXDpAhmlIqe4bT0J8Ltk5iOfkoWrzlZpCI2rtutAFuX14CK+adfsP
Sgs/VgaGA4D/G10jEkzVbbQaoF4QM9lRp/FhopyCoInMnx//9tJzBcUc8zq6GiB/
VvlXSgGDu6y909RxIATlpDTWPqH/qfjWhfiWwspEV07tXHtS376gcR9e5/rx+owV
xbaXqdQAn0rjYSJ0/N5QNJlAn32BY0mO5kNp800lHIR1dS4+w4HBYp/9RyBszjqL
TsxB19jJnUkmg0WiirPeZXHwVA0BQ1zsiXTWoZ+hnBn+V9X45490hPq5dIInJ0na
ecvKhH1zpSvC2GPpDoAw5N8OgFVj1DSxcK1ZYZtfd0tI7+fau4J2yzHDz/oDLNny
ARq8PQB3l/5GfRE1BEDf+JC4tvAO3qmr0odljDke1T0NNxSxQGkii+2oHQIFdyar
LlPG3lWrHiGHdTS+QkVyXfl4KCQFECNHyw9d2L6qQkY7oZ/y+WdzemtbAQxkY0Zs
5YY9Ku/4ZOfBjmAE22Xjx6K61tQBt7QZ/dYSeAL5pZ0p5Ckwq7iCteRwOqeSgxYX
/e3/R1TzWJvcKDVrAXhlHqQ3TflB6+DrOrJ5OiSnoZNHQENUBcGzlTbhpSCSDvyU
MrC7r2ULQg7LMxrqURjcXWdexcuzwBFAzwG6WATtj/hHtTuwwIYcTFRLuKTDbT2o
HCwt1M+aWSJT0DOjTsmWdAJZIz/qfuew7AqyQ6pF1zqboDsuZH2lSoDi3BLxLAhV
+14uJh3W81gLNl4XyEAur7MHbgM0aSW0bidwOZ9iJNoHufTrILmkd6zOLHLVuAWn
ZnElJN1MmacxfWEUCGg5YEhki58X8y9IKDSJOqld6A2tkoxatysa75PDIjfH6qZs
D4bwV4jlPDksPNQKyHEliLxHxms0bdgv50IBwhguOHD9+nVN89x8DHJO1rYif6SS
kdtyE4px+IFUyGbFxEv6bvInlUu79wXeWI+9S79U2nEEKNf4pCr62ofCfSJADky7
8xSDSuuZtSNcQjpDgl002T2ZUhlkgJCGqfHXuH/yZ8oreClevNTiH7yrlXHdap5r
kl1FEh2EyYxqEloo7NrydhQGg/mHSI2XU36h4MRYFe24+oEKMTsSuck7a9fnImR7
2s42AUuro8HHdXzgdCs9h0+snWp9NFSmJ8KzREPLDB2zGdIDLaH/UqFkLxDHHOhG
wazLZn6K+uXbhhpVeAQNAQf0bm9IVNBtkAf+4qvgK2/F+N0iiqcdtrsVKJQZP6z/
NPbMsUyEETaMcokYT+PBo9Iu6FX3T1S0hxxARTpa2ZHJb9CRMoQ2DBN510KbG0NO
o3C27A6jY5ElT1VVOgRpEc/qF2tbcI7Ci2RHxSIwg8Fq0EMxU6/v9tzUbBleYMYe
Kbz7nNJrG4V6/l35pAclhVkYiln/7NZDE8Uug7DTxmMMZG+VUNcZ0gZjhYAMaZ62
3zrMKnFm6QgQPK6mST4wH8tnHZcevUMwFZ9Mv1CZD5sLKVG518qsOjACYnYDZIA7
QxtWOeDQmFg6C5bNR3TSTnhyVAShPX20mpESO1vaLxUPSMgu2ydWu5dbq1ulmPl1
6YBB9h9eaePG57ZN9rMvAiuouiw97K2gVQxpR10Ogv8=
`protect END_PROTECTED
