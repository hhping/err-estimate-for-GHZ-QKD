`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Es43wnPttNpqvnRt/BGa/M+DzFvsljI0sgeD3F7+9nS1orzVkGXeyK847whxEErn
itMftQEVVUJTG7ATdpqsS8WLHswzK+EWTcrmCeq4JIKQqlSO5aDfpEpxdggYGcZx
v6IlXZ3n9FCI5qAVRslGzRWmx+XARfj41kCs7uVXGvxJm1Fv84ViW9vookt9JIgv
+64OJ5rIHN7wHBq7tXfpvkdYMgdU1Y5hnocdB6TAl2TRpo8GTH+KvvJCc5uNIFCd
oktFA4tWk4lwe67kmWSd7TigV+A1a7ySHGjMNpaHQ9bZ7sHRfzRDk/ivuh/2UNMC
HnBfWoc+vMCKPXgFObjxjiJqxFnuS3fyccV3G1+dVxLRR4VFiKk6IdV+2B2Xrd3G
UZp4nq/9Sje5WIXBIeLKkxZSSumw5gZtT+qgYpkaxinKCTmhHdQVIupUhC6cwDDY
jVL8r/pdXBp1FIQEM6s1jIB5U8X5tX2j+4wIV68CM+I4K95jopkvKjeVD2VZRAAC
TLHe3C0pM63jkHwGliJzkFRn3rqHfYQkkn2shDoh1PSSkAh9zy2moNbzSccLKpA8
I0wIDCHMmBloKxNEkxmqSX/KMsLYqslFsZWW7IyXLqNjuvBW3xkWcGraMmJ9E8iG
kANhyZ8iMsdCtkYtLqgU2EfywiIngw9yoQUn+YaKDEntyqy4DVF90u06X/u2vruZ
XCP7k9A31LikrJpxk480uN2JGmG0DyIrdJ540qG2dGujCa4xW/yvHsiTJiMxEJIo
RStrSuvexH5qaYpKLm+fqf8txiEJVaYixADmAKjKT+F1AQGUrtl6MhP7sRI9oxJA
iOYwRkMsUsRFOkQF8lpZtrIDlze3ZAp8Of1Lx4trN7U33DYmypfFB2xwhzqq5XjT
NbMFYtw5a3a6QKsZ5xetyBNdk7e/nXeC8Ol8nuTfE2iLSJNfCXP1zW6UrimDjbJd
dDbSW+rw/q5aGudwnJOT0ouh99JqhyiwBqzMw2JQanCurYytWTmY8SSPCDI7LVkp
AMGe84j3810iCd7uA0vMAlYtppXPVtyRrEkhhHkXjZqWPWlD05F/bdPXEMXylwiZ
JB/geOSuNjRO4rXjbZFO+arFQtHgMiU1TdM+e6RLK7g/OtYCYFFGGlMfqHgbjeUu
0+rqRIqBy/vfMW2WR/rMnZiaBbrkr5SpHENui3bVh+SW2911Y+7exZx19Z7cIJ2E
VukoQYDobcY7NYqEwbZDTkkqS9hZItCsFsxwpJLkPNoWekdimE83GYBpRy36mXaD
VWTWfXbg0G4BYca8p2EPO5rEdBX9ttSIVVhg8ZTBr+LJRAfW6vKV6Jfl+y+d6ky5
CgBlcPG+TpURB2i0QE4URG48l2zBlnL320eTA1sbSg4KG4c6+0PnTmpPLvCqqJP1
KX9ty0ZBexzXpCOmfHV6tJuaHIG6Y/BQrTbPCEx7AZ1FGJWvjFu4eAxpEGEm7dIH
ygYQ9aPaFqRTSXD1R/Fb7QtrRzoDLb30DgLS2bN3gRrjvOupG8tr3yNvFR6MI7Ff
Y5JN1+dQlpVZI9orRSB1Xipwq/ENVBJqY2S6fsu0xJ1v65y7lMB1G1fF6ksHBxwx
XCkfCV7JGIX8OSjTBhTTXSOpigJPEUQxP7Lg3tOyPmz2VUCpt62q7RUj2G/bbVy9
HZ/hNAgJZ4KaGSas0QMH/i5Epm6mQOazxVuesVUhI1kmLuPzUCf8X6rZJTZZ1gFc
1Q10dvJd3cm/3hwhcQqch/Gj2HkMqWr0k4NSiRGbgwY5wPX59NK0Nn47Uyynkwb2
The1fhSXtZNDVj7y4lw7MAPqxxGu+UnSZRjax+zAazE+jk3KaZ5IwtQ12kLXb0ky
xyfjpV81e/lzpi6AIayUWdUkWrV/FEOzAEgPYCv0Ae7FVKdWvOQScrkdscOoO+u7
t2TWBinbGZjd3Bp+XEe92VClOW2jIXzjG2eyfA4hWDcIzp8/pahY7uTInTbJKEw3
9Sf+nu3PHfj9dfX0qqrdgqGLTgoW/6/LOOAcaT9G1Te9c8QbdvYQRMIp7ggJbqr2
AhG7R9FgYiekwwKO7MLtHCMg8zf5VY9ynzyTALrGryA8GCbGZm9ABIs85tBuQdQV
baMrIxMt9RNwqUq5+Gr/u0QALXvnef1sI/t/kb29dwWLqdr//BfzmXgmm6zjnaUn
IurMtXsWVHlcKFoicJN105WWWZAD0dKcX7CJ3xYGhyWVpREtNIBpWN+QLaCYpwX7
Ea8qBQ2PMzCs7/i+GoS+swIA9MmaH/xgmBbz5oJ3iUWlPnDkiji2HIB1THaVvTRI
+ycCKJiDAp8G54D8MBA3oV2mlyQThO3xx/83mfAzTgZ3lXQ8hjwBTrhMoNLN9zl8
Y56kYLCQ3u59O4T+yPQ3Ug==
`protect END_PROTECTED
