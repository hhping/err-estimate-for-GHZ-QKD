`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jPqNh4j8rQqCvhleqxRwtsEn5amiKz+012dZPMN1qGw4EMEP+es15ibZSsOI4rhY
vzV9Ys/QTLikVCAEqrpGij9IMpMAy3bRTNyoAgCkh/jrdcDdj35HHaihgqJBee01
cLGIq0/ZzP7yculbN0BJmfC+tzmHimuLf0wIBx0S6kgV1W3aGZmqlORLv+9nvLnh
WLj7Ic7kNehXogi7a0blGdcRqgDuH4mur80WML46jgkU5UPoam++uGTSsaR9/1Wu
q18o96I3vB9BJgfk6R7KEHwjMoecNsciwdPvrKaW9HMH9RnRdvNnIyiZDwgY5mU7
O4kpHg/gJKWqv4n74QQFxts44x9tc4QZrTwT4YGnFP11LHbxLwzJRgJ1DORVlZjm
CSwntk4WWd2mCrtcgjdpjedmxfTdvHnmUVNna851glEn1UiFSMiGTpMtQEHXZ9mM
9qj9F9tnkJ9URb6qI5vHJyGvpMmLD4LUurfWQ+tmjRbkIJFtQ2K16WpTqXg6b2kY
1iX1+sEi4+rUrysWlbUXvWCjN6z64NKn7SKsL5zH/MtP0fKMpDe8CSjWeZB8TBYD
gYIlXutjdf4rozJzZr1Y4RoypPMK4zfFRpC5oXOoWjcaqNchhhPEiQ8NDvD4E0dv
4YjDAk9UKu3dZb3C+5a83lX520u4fpj+7z5qRdYv0UiKTENdOG7kZASymwMkP27m
W9C0m7jJqWsCd6TGJ0XBTPkWKO+qXUPwxuxQQp87Z3Zu2hHWylaldXOBEqypgFn3
DWWhzl/4FTpry3isX7d1A1i3Ei3+rGV69USNlLdeBHU0DKEjAJMuby7IxZwoybFM
+su+wU5Ib9/15TaP7ol0X5bhqa1WSyAQ2oZgfIZ9574Dz2fQ8Pzm6abm+YRBov7v
/O4RI1JhQSULv5aCqCm2FprS/Ia+fxDKTkDLX5rCGgH4eH+zWNXRj/0YxO7AkalR
NNj3Nsp7Y3VKWxrltZvrXhc4e4qEQJzE4uTVFWvWrH71vJB80eMcSWwWWxyvBkqF
YLkBjJBg543dtpKsLJCnRaGdo6o7ujXuOdep2alnOzKqenm67NgLlMmxAYoRVsDO
cNzNqUeGVjX1B5ww9e+8eQVylbfCQPfv6l0x/pF69KTgYm04RUbLPvgbMN96QrSY
O+l5RfiYKVmAHMV7lLShqQn45PKeWnCZ+rMtLSdoGCxFMCJci7Vc4OaErMs6189n
vBLeszPtRoTOpfa3gt44t+tuYt9prGNn9ywyCqB5Ta5Rdd+PW9NNfrENIigl2WLp
fCJWziY8Zlsuw4Ib0/WTQo9/jUuSLYv1AeruJF72jRBc+mZirJVeyZwtCITH8Pnm
g5DDZYhVgCyjiQ+quoe/xMlX08K5rYl4Llk0v1/AwCh/mrDFp/7LM4MvbGrpBgRY
n28Scn7+NuASvUMec3AQwmVchhMtW/ltS7BDR8gu1AxxQ/3H0Fu7McblXgzHOHVs
cIIccgU1yEnqhH1+QVlfarBUJKuOHG/ThOYLT+AgrMKOuKMx0u3YPzwOPk31sG8I
ljjLOzCOxghQ65x41rQDi/fGp8EOX666na7EghKUXaXylqG6AG7F8K2dvcIDRnBf
xyhVdC89C9BB4KoxvO8gM4w+c62fxJhLDZ+aN8+gdN0MIZvseSJZOoDJOCISM8qQ
X3H+RCIgN7mJ89HN2R4uE9VOsGc2Uc3XmBs3LtK0lLJ2tIswGo9ht2T+2dN5PY+R
Ma0DAPFTjTUO6dARFn0uUZGUmWqQRXHYP2Coi3HKGPWzsocaty8JvsYyY8RD7500
+vzKAa1rxobVyETRN9w88YvOTD6yCAvKxgCGi1m41n9SA/YhWRuRbVFEUNFex6+M
rkNTMceG/QTFzHkA19VZL0n/FI1qQuBCyYI0r0/vrzuEYuT816VWfVYECIdqa8Hb
`protect END_PROTECTED
