`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raIClWeLWDbRw4wH5x6Ss5OCcbDIXu+wh9PPUjmvtRvAlTi8g2p0Qk9iu+dtcqjV
VFRPhc1Wt7Lv2rC8VDI1G7igGZk6+4c08TzvXTRus3VD+7IPZ4bwbf268GVxnZog
3NTO0X+eCeRBtLqOS+Sh7FgpMUxvgtta+7EPukYJY+grDFrTT46RiSxyG2YdOS9Y
1GjZ4XseeYCvvdf0ahO4me7i/P1wstjhYKrO6fJmuBPTBY7Vx+vfM9Nb+J+Cncpf
UmoV2B9rnlDPDTpBdTVcxEiMNbNBC1DsYdErwomzccDd2VmEIslG7pYzWdmMcwr0
itkb+RrD8+CofNFQVyeEcX2K+dIbGRbT7zt4XRb72MVUnkrTV+GIpqx9ob08Ug7/
fhS86t+LSfU5q/o+QkehcY1QLIRj8j07I81yeJeZlGikgf0o7xMc5hEbr6q43JEt
wtm+h4se3uu6uGnguVI3HzmqhSfspyWRbv15IN/Pv6ye5NLk9THRLmGsHhAzjWi6
QRO72kch1pL57X/QuH/8m8KJLTVbqfPzVz6QM3fActagOkR6ltnT+m6q5e+zQ1G6
IW7YkdWuHowtv9YRzubC71n28G8olvq7OCkx0nPbl/OVCNPVc66Fs32XrEU1wePa
RBKQ08D3l6L0Y320PwOEB+jTpNUfwJ4+GnLH8vqRrqw149jssFiU3hy1YYTfbM2D
W2a9CpP09ct4Wyy0Qx7wAH8qjE34jVGFpJlw0Rui+wm8qZfwCaSFXSXHiJAQZpPO
mw3/RZ7CgeIpfab4mpTqa4m9DkJ6gW9r7cir53YCYwATy4nQJ2OKigUG9aNf+VGX
5kD6NTqwc1srLQaumUGzbV8nFjb5ygwfYQLA9Pqo5dVoLlxTy9e751GzM/0x/BGX
9i9ASYGJzpS6WIb1Gitj1/CZ3WtjUyUvpT/B/z+z491tF4L+PrlyWxTKDVSUnGT1
09T9dHC2RBv2AfK+qjOpeg9+77wnaO3+efNaEXugNIhogual5axteqqjJtLzE74e
nvkvC7loZsp5K3rq276JuZqBu74SQe25Mi9ko0B9jSR7FNabkfhHAmBPxj6KbB5b
JcApYUB6rScPtDQlMSOUhKL72LoH6gNS+xBO4ccGeVKIrcJbA6bQ967/M+6OwZlb
n8umCckywQ1ZxnSXEJwXPwa+SsdqLuFQRbssL42kN1gBknY8FulsqKUxfXnNTmyn
k0udGu/vtUXbCsCv5mmzEN2ZpqawqMbYJPkqukAIpkpO6joyBMc50lyTGzsbWzNt
vxA4dPa3OUlNOijU0EkESZbDq8r5LIVWWZHhsnLiUUfkrLKKCYiBb/VfCCwiXz1h
QfCvQxYAzEuGcZPK0eAynkHxEmsJK8SYUZJy7YfR6aTyWJZYP7i1ud7M4UyDg/jr
80LYv58xMXPDClDZhI9jfcF9vFOizJzhqJj6NiBRDlqsqbzWwO7vZsQmffiwFsUo
nSymm2g23MYsRc5UZkoThhZDFV3uCQzYvQsvodaryjl/l4QMrbdGrIx8Yx8Yjh21
VJClpkoTTJB8C2hB/j5QBJUrZD2OAlPDNE9gW7YL9FpjBCh21sbpOp5l2vrMjkvz
gKxgrSyDcewqqIWMBic6a0Rnm6ZUN8JO8spNKcBvZuHnRRbmSY/27Hyu/NkwkaJw
gvtPxotKYnX9tAtsb7VV6b5WTWYk0EJ0Yz4WYlFI/1Vj82pdQ46vD2J/MacnetFX
UiDrMU99LPOgrCPwv/vMZZCuez5YYS9ZJwIKCcvxkBY9oDVh2GDEIvR5DB4jTOWT
MK3JSsYtZ8heODqraXkTP7mUzMsWwXTJ6C6E4BUaeNJ3tMtF1CjfsjIk1adV8nXg
YmBIjC7oKOmhFEzT86+TcvjTl4Dipb0g/4UiUeRcs0y2uH+pZ2ZRnhQXzxwPU7oM
xQjOte8E7Z5Wzm39GRy3J0bi7JEi7e6OYGT6t1TDaa5zObpPkXlA2hsR1Ze0pRpl
eRYNkLXk1pHlxeSyuKopY83IW5eNJy+MXKUs+tClV7/e1n6Hzp4MiuieV2agrIaV
jil0X6XoQq7vgykUNk9iaUd2nVrWqLDSoa7vUQ/pdbxmGDKeo9ysZ1peHZewngZd
r1YFEfU2EGT12dTgm9fq+oBdr8xJVgK221bomNGCDk2OJMmEQlfI7PZc8dU9rBVD
97CEs5CzVVBRRfVAaFZsGmpWOsux5JJ/w6o/VO0cq55o+fkNwwuFaKVLqDff2FO0
U9W5sdiKo9fXtvrJALk9hQYmneauFPTGM8AMfidpjfN+KYZkE+y9qSG5nKiVCXLA
mUM42rbZKTFPnFaXsmnwZ6rzDKMqXwH2w9VGflyTDWi7DEbxM6rrmYzS0sKZznyA
m5oFBiHRPWBh+rp309i+50lXr+nYSJi7OgTfCAiHzAa3KO1rW+RZKCRhNFRVTacL
Jo4N+kk0dQ0azgYZweiw5z4a8uCFY6qrLFh/ntOeH9elHuDCNgROnG0pO6N7TteQ
CCUkNrfBR32HadyJ/Lf5lDJ4MCwypPaZ3zrFIbK0A27TN5NVHvnvTpqQaxiQK8u8
HnxotthxZfVvEZlnQqLGqNloZFttqYk4bCr69bACsJEFQvbCoPQACSVJMXgy7j1s
S/QdELywlVtgBV1WL9GzZrmoXHCZVXw2wqWN3bF33L9yCGDj4kAWKXa2EYjy1n89
tFJIbGdKK3qmtim4Q+DewuZOCXTqx360F8q3+8ZhNb3Ue/u5gdFdN0wW/ZYkw9QL
amLsnYgJbiZs5N+tCb3VSobldx21viDzQk+JwvhwKLrJcJ5TvIuceGbJI39Vzxoc
ffIv5r36/bpoXLoqgL1URFv8Chigk62P62U6v3crAh7WaXeJ1UNcadoNEilfX4ou
XAXap441z160lOVaaN7qmfSf6jCz782ev/ADv+LDuHmWWRjHZXWpNplJUvnpDX8C
a+aR4UirVK4VsJU5XG9uOK8xY5Zy71i8llSdsQwEOpQN8t3lTGw/LnM97xeZjhDe
Vw2ZDRjUcry0xahfAaIaF77eqy7m6/RIVIUy0FMfJ6LoAIyxJiVkhl0ukS7gxdrF
9meQv8kWGGK6QTwd0Qeg7PGtBmQ4+x4LROINRkWljV5mbLkQCG69gc7Am4hKzQ4s
kwlHRERWD6W5mjOE4tXbybx1hgAGa7PPkFgBZ8Do443D3AEGIHJrF/Dxc8wiaYv4
nOeRx3237CP2HvDo7ntOa++pi+SxGLp15Kj6o7LhI7jb6TQT5uC4T1kx5j7ydIjh
PuQQnEKqOE/6ULwESOsvXhYeQM0jZzgk8tKfWbCP/iFF1lBRJGvSVF7LlKRKVk6N
ozuk5L49ysIaTcFLOam9l4/T9xX+fTcgECXihP6ZYk7GQHLCVpgNDy8OA/ultWQB
12tbi9LxAFye5AtSi9J6ygxAgWy9SJuO5dw+dH2+qQS4hABJNQpbdpBMy72nYzoP
IZLKNIekuWo4eeDMkJGCFc6rlbVjPlaLkuJLhR9EBAY4R5B/8NOcBrLGbqM4/+4Y
n301PpwgKk506jUxmAx8EOSCN11AggyGBal/JGOUEBYnkVtGo3ckz6RsSmH6w23A
jAj9P/9eYNNEdGCLj7hA8gGX0+Dc/eR6J7SRUjfTG1QFeDduYDBCqkHh3cepB+PW
5+CE5ZmWEq942RnwT2NMHqUN/hLES4MZVhBXR/Vr9MefGwqn5o81CgDz4eMR5Wbo
MCCIPCo7UAK2Eo5TtQllKUACISw0tv6iXREXbqV8FmQXl55H8lWyhqzXrEOmwPjH
N4p9+rmcymWGMhrtzSoj4GK6oK7q5ft3u0gVHr1YfcnBnw8ftXEZ6DJGuLbODIJ4
2mYlQQNASszk0QsAbtgDYzRnTUTAnIcMZYX8ZZwgFad5vFf2CspbVAdq/F+Bhn4x
d3bNGmS7EwVD4OKKbtpW9QxGfLAixkU+3EGZsA9/GXT77HvkLyaySsWevG4bm3Zo
I5q5mOQmKp2kSawuf9Gwob8vt4ACXxC/tYmY9B+EJJDSWV1nPzsaayI44oqXdUiG
Q2umRkqzyDV4Mtp88dFqej0O5sRNx5OGQk4v4hS6aEQEpMZfLfqsv+NTBc7Odz20
GsxV/i1m9Zo2w+lXTrZ1kl0TQ6vp10DbB1+RylPH/0LGkHLQ1HVpcn7XmXHtXs7k
CNnpmDxLuakbB6H3AkHg5GJbtyXqmlrVKS/b8HJkmAhscSd45RAddBOjTMNJ374F
1Og7GHTrsPn2+vLM47c8Y/S1ggKNsCgD4nrWjSpQ96A5zimxKPRuGLZZVji3it9B
78UwOq3t+wc4GqGdELBL5fzuol/I/wY/CDC9KRQK3aNdWAQZtYfnselx43WASeE6
Ue2SA+T7ouJLDQ2K8dSZcVUOLaK2Fi+goZBlfQ2i89l5GcODpvvXo3OUXIdLJ2m2
IONfH5sZXi/y64HsGrjhnqjlQcJYMqPTzSCghFNGWY6UQOcV9iIES0tTqFO2OrcP
W6rbyu5l79ThsgGJgOwluwxX9aMFDBK2CC44Tx3dZg0LLIY65qSC8uG/sI844RMK
YoJCpuX4GWeiOku3tIZd3i9cynlMaR3oDxDjVTm0g8G6sGwQ5YZSVKj25EFs+beP
/5Q8YKmcDcSW4uy9QI30MrNEA99h1ffp7e3AcxcJVE6pxZZgpXAgUqVrI2/8umW0
YCblb+hBiIaQn2eYiZAxT7GVN1BSVbLHvqaG2pwEodIEvNtYyt50lsvyCW5OcK8x
OJ439v1NtC9Chhr8bnDiQ48vcZ2pugZhopNqLOf/rMzraZs4iW7LfoU4YbUhzKL2
3ouy5v0DDeQItqn1BHHS/4o8CvMBbuVBQ4R/zYzvv/EFVa0KQdRcvttYS4LmruXC
6c0L/q9sEqqMssXT1tHrs2F9/reDz8yAkSALClZOdA6qwJQ5O9Ij96qa01wqE+Zc
xgeRMzR0ySJhKJtJ/kuX2DrpwfTdker5GsJHE9rznTNnr45dK/daeIuUJ/UD7ex5
U71Fs10ALRhmGXS5r4JgUWRa4P98KoFhp3KOZ6ByqfCkHMjV35AhJcpik+lS60e8
wnIax0uYCeMQyZGth9MEvv0D3hfgfIfkM0ULAsBfxQDgyJzswwvXlxiRSksULbpL
3o7h93rDXr2B8aubao5ZdY1eipeusdvhb4xxVAiExe6uQIz3E8Hb+1gkVkv/tmQ/
ebYFaMw9h6mjzYehiLToH03jRYRBLOAURRmB2LXpyXWpwstCrM8PbLzIFF8gdXwO
jzvGub3nCFH/pnHwUd+tT5FSJ4D794nHy0ID9o1NP5pgxQ9RKC154lhCY8FuvQIV
Vx8Ylzq1hGMW9/wv2VTTr7vDs918lc9AjKonwgM36EGP2ZYOfIU//G9c/TvFauh4
+MKjPHYErqNciQrn2305QoIhEThjq+K8+I1FmPC6mgB4Ce+zB4qXS9pZ37vESwt5
wMysOlhQKCoiXTuKgYfCiieXQeAUtV5oKQto961wVReQYa7NxEzM/H9at+EzeXAr
BhvKeXr+aBemIiIhLqqR2CRh/fxtPkdNDCq5COQpXvLDCUyW9TjA/F9NTKxj/vBE
wa+9ioOfQ/owhKkDfEVacz0Tco89NIc4mDN8TnZMB2YDpHQe1y4q8ECQmNCZlPYO
9A7Ug/+9BYYShCcg1dOuJy0VQKQ2S87VWWQn8DpyZ8lywpkrqUgwoX40Z5E8hXI9
HNyKHhjWt3YZVk4KI6cSyz31/LqT2KX84LB0SqSAHXlK5QPoQGhsqXeYu0L9A84M
/vFQ55FgMsrmAE2Y08HVnxBqixqgVW/O1CBvJseVUYsrc0mCmq90a66+h4WZ2HtC
atgtu5gBGwiFLKljqqXZeBedZ4xyhpMBthW8yLBs44X929B5F0PvNczZRzRY8+Sy
4uryO2/r33NBEkWRU7ZeHKjtk4SOAB54bjFhlboGUctxEIkmXafyWj2u1fLC9kIS
28Fs/RcrxxSpuUMNJV7MzS0cWfUuT4SB86b0sj4qNlwsBm6ivIpizZFxA/c1dzA5
rDzm/OE1m8n90vflPRe0HWlVGu3Oq2wjneVfhRy8Ss1h9E+z+8cmq4tDeh87MjoL
E0RhclY08Efrvpq8hApkNjDgCBI8liQ5LCw5KgpeLp7MIQsGkqOELpvVgkv6nevv
38vURWvkrCWqvBSdy2dJxJzccMaMnBFeqAF0yfmriPLqe2hZpdqfZeGX0hdOE3tD
Hdjh8LuQuLHtIjknygSJDuudmk3hLjKEZ/UDw3en5mTQX6Dqtjk6gDp8rkUsAVqe
3PfJkSLxrsMK4Q+36OJ0JfvMlJADZlBQRlb7/IZBCdog5rS0Y7wAR4lrax24Aj35
MeXpXrcgPTS8/LdGaQh+m9QA+h7Qu+vP4fUPBlspX28qHKbt9mx0nB1pNy1g3Lku
rPw3NaILPQE7NwxW/UlyyCgv1csNGAj6oOR0ad/O45o5cp9F8rWKVGhZAPj7TrRd
f4IBYErkcC4yr62X2r+GBiKEn4od0PTSEKJA+meFfzOGzrcfaUTpC4ke8kzXsEZ8
BkxPyGH0FPYzciO+4C9h14vIhqXl1jtNsYFYApGtS3WmHrM67va1ziBpYDT+Gu2t
KU2gKqkvv11KtOsWvqQ3eDDDDJs7h9IFugpOGxhqC4fZ19Q6zFHB7vhruwzSuID4
iTQsbM6TEqY41tzkDcNsL0AD6cfEbMTVad+xoieJYfwNo2Gl+GBss/XiqlrXNfQ3
LCTNRsCjmbbNYPJzwK6xNROnkBfNVbiDqJea0xpFuXkDoNFnUvRELlwceF3rWzin
MBefs8/XOL30pO/FvuTRLxdUcTEl43wX1wPMWgYiM8mUjiJfJdJHm3REUgVeprD9
p0KJ9zKaXXTKC/wDPgPGZvpfhZlMFzHg8Xg5dem6m91PRSt23XSPOt7PerW6iSfR
Y/9GfD4Ry+q9UoqWb8lyzXtBEq7aBJO739B7B3wp8QpTDY1YEyl1vEiGlnL8T1xY
A3h8TKpJB4uMWILlZeJ71ddcVlMcUuj9IKNAGLDk+TTxXC+42CAMR9wqJ7JocOwE
YcaO5Mg2HRR12DvPM3aTHkZN494P3/BBvVVcr6u/drf1gDmRn4JyfmZ57YZ+nMtG
81hF15B53QX2YOROexqMr7CVk6q1q8yHcN68AWFQ+ZJrdR/+hZsRP1T+WMCLAhzZ
901GBOCfe3YuXfkd0p+a3gfOLxhY5B5h2KSwwqr9/JC6blbbkSRlQlBRzyHxfyND
OTVN/C4Wne6voX7kpEJnPg8aKnt/QmhGC0b6O0Z63NrdwhOEUa9f9JzrzkUt+LC1
pof3LBr4tcFBXjORjqRqMHVnF1BKmxo70Q5PbcXdAuHiRoVLqYjP/7ERs6qFfC5g
zt1OOC6GkjZ4fOKLpS3B2pc57y5WAxdxE+hfExFXPiJDTN26CHGMyjrmIfw9WgME
XtDzeGxfgBPxflLmqVxz5O5r3UFExEOg4hnm9tkN2Jjr70cCDKw1KNeBUoPlOYaN
8/y/t0M8hkmnFHc3kcYItyVneUmgnoTHDFgmP+fpZJYXiJ+QiZR70ehJg92MkwtV
eT861y7h0sEazPw9oJaaIxfPHli7SNc4/dCToasVGyKQoUcxepF6DD8cgreZe4tD
RyczFYWvuh/TpukqnncDUatJfZ+hro3L5w5KpHUOQugJY4dIMnM71o48KEL+Zmpa
2eoX+djXhdSQvJzOgUHNPk5h8SvdbP2/4tVxW5vXgXOpXdNyMi7fC+5gxPevRNxO
dpiyP9Cxl5dxqTPIUlRkI3mUJSZKAZgClNZsKRvvmOpXL8AyRIZjrhmjno9LhOaO
PW64kO7D9sEwXxxOWqdDv1S2ufzy6OZuBXsdAldn7UjU7bqzyDohfFqdfuYI7B2V
hm71S+xBA+KABafelJmsTzTWSzwFzZHvCHJe/L9X5x3MIbYc3jL+E/qvub0VyDmv
7ccy647spk6M7zwii+CG62vbqU89KU4J+MSoTsk/RcKuLjNjJqTM2na90vMEviI9
mPmokQJb4/KWcJudWi9wKAY2RKRk+GxrX7vHN2ErOheOfJc6WpmQZj5ChwgoBt6B
DS6boISxUWWtSbtp1wZEOxSxwYV4K8lwjpRGqQzQdhYqaNRYL+QLw4v/oxCehV/K
8RbYk5KXoeddhoL33ovBJhYvDiAn674Sae2hFRd4FOSyO0XbRY6yyA4wKfo5FdtU
pF2SyQo9g0SIrSc+rlj5aIv3tTth0H/etAVQeHB6iNTYkjNFrMvT1SqHaJQTL8Ga
3PMbNSGpfV6t9o4+SzVWmVQd2keFmyDovUgW3afwPjjXWYqrrHG75on/a2+H0i9T
cXxo+14IPZE53iyf2lwBc1c//ljv0LM87BMeEu5RQXllzS5QNRD+5LG6gaT+I0jZ
edg5V9Hm9aRgHOmQkSoXOagkBb8fgI65yqCgFLW5+R9mCU8qKdw5dcI64QC3rZ2d
dqqj9S0kiKdZA02aE6eb+UbXxRv0vPE+16l85oD7HlIsMXZI5GafTtcPxfAG05eb
objYKw3fjRF5yysrFwp4YGujgbmS8SDuNFISuV2mGPwfQSWlHzYzh3IU8IBX5oGX
vkKfR97xm856U9BFjN7uejxbFrEwk+nU29GBjMUKguqZAP/8y9KUNzeBnocebh76
5eK3PAeh6UzRBqiBiF8tVXDBKgNH+r1dT2JDsZqKmmO7EjTYj67pi8z3L2lqKldc
qIUo1w0vQjohMB1vnB/+bk9Mn27o7v0DpDVGuycIKfXbIG2sVhnGhe+m/pclJOyl
pxlxLIDCbnn66NSEWisRtVmMXiE+d4qm+vGbLGRriXHtINUNNWRJkiMgBQsQlafA
taNrZJJYV4T/WfhYFB3NVfZh2w+nHESXZbMuG6auy6qW8t/r0HtAdSdTNmlzSt5/
7kVUqHmtRsN1nMnnfEUrKavUht/kn+Xt3sfq+yT4hU+OJUP6sbWLpLek/Tx3dv2N
P+B4WZ+pKkzeG2u6XE3qBVLyPuX0fFY+U+62TzZdr46M0QlAe8ZpPHo9vpy1CuKE
kpONWZGijbo/ToQKh+2S6uaM2LaRcTEq2TtI/Y/HEqKFrDOMDnEqPkQKsEThycwq
ONK0mSFD5OaZAQ2px62d1Z5mpHBxe2/2FCe7bOnwTR+WVTR9iQ1Qpytl1xczswxM
VxLSTNAmwxwRJwGqxI2ifJ8De5zZxlp7X9YuUGQWCgyLYsEZa2epyMPsmIqoYuaV
tbhW4povAEurYVCrPDAVGC57VdXitfoGmhpqALHsuRJ1GmaloYoCXvTq+bM55zNd
84NoRUYt43g2ruYJK4w1rKbeAsaDCbc+22KFVH5YW4I9MLE71AGnWXcb2S7kEbGd
XGlezTwPbbIepvWpTqbUmL5JWbfFmCMiC1h9F5L6oQJK/726P44YwEHXOaMl+dhF
umftBjjZ0zScrJBwwq3/Ltn+Fvx8tVHzD7moRuvXdommMKPT3ueFyiXpEvFhNx+i
lbDvecXJQfY/ZiiHfFTS33KNQO0yFxRKphHOZOGPwrE5ONnbFRH5j58o1NoXOXm9
HXSuXgK7rtooGdUuDYkJqJNqyBSBzOezbVoINSgsLYEYuk8p/QFWkOLMoPpof6Iw
n9mzLWpZVPrUQuGaF4R1cTnKWB17A85LgDNQhqZZ3Uu7CNs+43BYHH8aYEhYSH1z
VstfO4TIxf3Io5dWbWV7qc5z1b9IBb7vF8MOABke6eOyol/R9aJbcWIOJL9r7aX7
xWrgmYRbi3IJmbWSK89oXMc8BSVcm5PCyo0a563+J/BgGAsgQUu74w/PIE7vGVqP
+wanndJEm1B30OEN8RShSJa+MRxM1iDa31zCOvpgRbc8FVo3D4TvRdRkq6HqnuqU
H6SvvhnnRcUANq2F/sqYRYcDP785pXIgVhZj3Pjrtd7q9XNzGG1NBL6pnfe3Hmtl
tay3QqDa6GKte1YwjKhpsdhIP+lvPT7NOhY42vgDmupxDwzknPdzswjtF8eLNJGg
iFaZd8Ot1UyfvmU7LRpR/8VDxhPuoylFc4Qog7pabhMmDoQhJfzO2NPCHgCSicEB
dCsnRgU31M/raxC/5ZTLLw/HaMQNya5BNUEW3mMGo/fCK8s0Es6V4oSeh8veVHN2
2OE3d51jCE8GWOhbpUTtNOOCx5TPz0F7fjNg1L7CukCWZ56msb8ojoE7KCd12TOn
sq/sfmDSnp4wII2XxGH5Ebjd+iMiuLQHR6ZI7BpGcDtq9JsYNSe+BAt1GY1WvkZy
pdVg723Bl4Mz4Yl/cWBRxwd+NI6hEhHtVA+IK+AY82F7C4aI6PxCSED9hcA2vcga
sJiAg+M1ugpINIhsNL3yqTEKkjS3daT+Z0dMzYsi6SwcOBWAsx3reegnIk3v1/Pm
x5d710kIh+YVecaG/xM0H4r+Ano8CKRKZHD65/F5/QRJMdg5v38PKfOZ7TuvbZYX
MxBVzTeuYJvVMekiAGfvVDYX92d2HT3tpPcBn0fHlt68klXFOoDm8O0lBMv+7EF+
fLcIGjawnmsHhgsj0fFO7PIjuepZvAYdYW11q1yReeM4jH0N0+x3yduNlDczAD3B
nOmJtoOIsZhkZiUQhFw+W6StHNbUL1U5KiJI+VO6p11LHNZypG9UmRhf6LOcMecD
fVTC3sAcAYwBv90E22jrF04KTwgocipPb5wQjT4QJJvJifgfxc6dK8s3rPE7c1GE
0cBaowAU4xTp4XHwG1/wYhVst7QyoBYnhkBcTe+mk3RxdROU7yBDmc5cU4wzTi72
Dy9mqsnVw4CwXvhwJaVeRPJfIEoaz06ofrHUpuMprc0RH3CYFz3Og2Thh1/DNBsL
S0x4aLJfQ0G4qZ+lbwj36oje3iLZqVka1jMmtxhsW0+RqzrZMCCuTuZM82pBf54q
eGZq6I2f5sMAdeW8kIdlmgiGPRk/G128Zk4rCgArREu1yw21zE6hq/xzkd+dGiNn
UDQmBazv/Zq7rQPHRt8kGLcTbi8v/UlvuarJMDaHwcKFgkyB+Gcl7LRQFmu7KqD1
MVxbx8qDCB2+RoEaERKNb9vezXDSM/km7UTERNXr7VOKrB/no4/J0fSJ1MafHFqg
I6dgFZ/5A1A27xV8CBQNnPbQg78Wp5uBKohAVOeWUx5GH9zHOI7VHPwJJKjnxHre
vHlem9N6nBDkwTy7Ycy/FoQmky0xlavMFqpCJ13ST7WPPunzNOF0PFbkKP6zYt8L
tl3jzH4dgKDrkq9oRUbZG0By3Rmr64eNSVzrvFm3NV9yyTfd4MLfhKLDFIMe2oRI
xUqjIz3XtpEn19ItbIcI7NBVNwNK3ofWFRZDWRm55V5LJg0TZffuXm8Kl0hWLuDF
vKMCiQaSqBCVIn83zxj7Eoycgp9+mLScHoU21K+228lCfD2AKkU/YatoQ5NsVCxY
r8/YvHqJvNJ5NZRpSxHawGBaO2r5bVylSpPKqU1rn13O4vRhXWyOAh5aDDrKV+SL
igRAykdfi0s+5e7oBuCTpiRFwcNPF1VkGDauJy4yZIT40myPCiyq15iAi8J7x1Ou
ZiRlsvCc/lKpY2YFf/f4/ZLIbpuyIB0AqbUN7coxUnj5l5Q6a5WPzZpwRO3z1/7t
0k0hp6r+lfQ6zDz8UbAaM6JhAeq6vdQ7kJr6fYjupO/YC1f6RiX1aXJPI6LDjisL
cq/oldI7GPqI+mybB1yvPm39tuhP5mGBJ4sHoKiYp1JaQcAYcYhJVqKqWjQ3IXSi
67v8IXzU4kkVVLObGsYYLAUoXIZoXAmlCM1hi+mx7hARNyHl6QfG2qX6S3ZZmnyh
0eOyJntYMyu3A19lLC21ynKQXlJneeqyW2uOhDplEYHlFkEejvzTo/x4lsXYAZpf
W5eIUNyqbqqv84v3lkFruM0f7wkjpoWbK/4Oc0YgaAIQmXLrjszxpVWYHS0vI/ck
QgSvgU5feQq09Pz2IaC9MZZSDAuwutoUEAkyco+jQqoqTQajVp46Y3eUzLBihTEi
fOeHTofyOkXWEaK9sLiXTDBb3FdRzCtbYjIkcAUchavIBZ5QZ9mt7A+cJyqMXlW3
FEgJIcu8zqmBNDe4mudxG0cnG7Fwsjs1YHYIyNO3GfclXY2XhUDYltJDeiYdZ6Z9
m69mngoZ/Y7Yo3L1PDW1vCu8Kkt/ahUKOoy+C7RcGWYMdfScg6oYwtuvvMIc1DWh
lMYqFEcvI422Xa24QetsqXj+fGBBbls5ymA4h6cIOZvn/PpoLfsn5LpwOqH//7wZ
x1bTilt2uGUE59ruus05sUWh2p3n/Wpg5ayHZktqwFFs/lWXeAgQ9zTR5OHOmD0Q
aSIL1owfF2rb1b3GJuF5xm44+crJvuoIBn526gVSwUQfHn97cRbejbFf8fcWcDZw
xWWEQYVu/6nbPQQzF1vxTP89JCkDL9ydtP9wox8cAniJIQfCZJkSaiFgTh9/5NU9
4pOFflcnY4bC1+DBhioWXLZg1ActXIV+DwTLq0+iwWwFpoCvO088ewQUFdBALw59
wjyNwgSKcb+DNsteCrSSNCSjtYtks0uY2e5BvK+7RN0Jk98Xg0vOEGJw0xzc5zCV
Ai1rnMQvAJeGg8rw155JJKS2o7Gijw05T4iMmZXUeNjuIJ4+bAnbqWkFQtZTKvh6
Oqqd5d9kyLJwzr4hpxybtGdw2VPusIHKEollKD2HGhLl23IVbC443p21lFrpDTfM
1Xjqex4r1W31g0CLSjRpz8wky9pQYWy7POa8kIAZgxT8077MdN09CZhZ5xlhlE3h
GcGe8hwTksJoen/JsyFVDZSKXQSdkp+u9kyYDDBL44X7U0Y/MpJ+LGwUsjod/gN3
CS3/+Y/P90qVQpSnUsc21X9NGIxHsm5WHsgppcZj6jkc7R720fO20CFFqNw2TnjB
6CfPRX6FdAyAYMyUiMCTxW4xEItWRTB6ChLLBpok02f8x532iIOrj/ux6nCb/2VC
3hN0/4BMwO6VADcFQLEsyETuhZ22UhjhMY1XPr7m9dqRMtvA5LJqO936kMOYrXAO
eIDxfzkoDff7/NJ84/QDDQLGadLoqb6Y2lNZPF3BNajhy4S7hxBfQXrDyCejJzFF
KHJFWaHKyQd9kYtsGw+T4VLaTfIfcdiId88CvtKSkCuv2RzSsSURPO+14jTyA6zE
NcmFdEG8zB9a0DFw1z24sH25c7qW9M03EIi75E2mezNqj+hbuPnU5DEABBMTmzFh
r+hGZRQekYqS49QG1c9KOFQxApPbXc7AyGa8wrarpz6Gcrx/1+77TBe8K49xbXt1
3qJGTsg61S07RtjgZXJ8iyY3PL4JRgSHpZhBwiTayD5lU/tBBbNeCO16skACGZoc
LduDWqqRq/2CHbpZfasGpFpAQi+HDKwOjWdXwgbWPB8EadXDHC1r6VWy/4EWyIp+
aaw3+8n4CdrZYJ6fhp0g20wbreOOUEgPcZpAmeQXQN8bgj7LO/wqIeJ2HBU1Sm+x
NIkH+0iK2FEqfSHNhy1JFCIlhPrg8UJbyxSsoXPGpF0KrgcBQGy9IA0V6EWg4oL7
gO+R8WQbAHmVhaFXoEfE4IrGagSIV5ps/08ue93aElwythReRvXpTOYwAmklK/rc
uWZRRIDpm3emU1AdtoCiLX1Mg2VKpZq+uJIWjpfUHnwh5jmCeOcj7t9JvS0qEciA
0msO3xj3Z48oK245+WNyUhzaRgNt6ZVHcz0p35OUFLO8wEtV1hVEL/hhxKdz0osQ
lSnl5XP1WWfRzBd5dKTeSiNdFezp3kueXiHYIUO+7e4NexulU4YGrfMFtL4XBfJ1
HwRjPVgnK9UO/rFHKSGUBgCWlaize+b4YqrDwQXqVb0sNQLD+ISXBvP9iTYJSdyn
3MR9BSLjacoSVk2fvTj1aiPrqCPjYyy9Kug5YLAc5IyU4kA/RDx/7HAYZK7tRg4g
H6qXbWh3Odi7Q8C0eZW4cyY5cdpUNtlmc4utlgO9uRrRhsyAVx4yM6ZozCe7RNGu
l/kbRLxMi5r/G6+FAfYmp9NQtVfQ/QrgA+mSGEiOuL9YHK7Jq+KimQJtzxfg1Hml
+Fa5Bm3a0PxhtcsGGptj7KKEgeVCrjGV6jIJSV8CnssLXelPptPc285z/y3rTAwG
ykD7pHRmnnCYbR8pWOGCf+fwwRiHK2vDFhk8Apk9AEwCK/zPEFkU9ZLVvkoCH22e
aBlOgpYyJO87OkoFIUr8eSQKat/19GV769uiedCzEgVNwGTnFJ5g1WlOzGjOZ7w4
545K7fRl+k8M/J1jZwafKfbW8AVr9de4xiSD2NEpgXyQjmRB+h4cshhLYcZcMjSM
sGOnvGc1EMTHsTDUkPfHX9uuQZaWXwSCfmqvG9NVk7nncu4ZgCZ9R6rcMeWvvKhN
nzlgoFQ18crudpeRiE2Z06gEqwirdgdaN/DSiVv647n5gqwnsrnpRdJHs9M98X84
tpV6WAyccEg88VaLxjphmMT583VSrz4lH2gW74l0hO/pNU8MNgo07JxLeeI5CSQT
SIp9Ig+9idplMK1d2MCGhQKrO6ZBj3Hqu8oP+HdEKL4c5GBowqmjXr8h7yfqRo8I
65c0Av8cnn5KwyCm0GjWew==
`protect END_PROTECTED
