`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WbUbCtCB545+3LvzQ6Qf5KdjiNzfKJuAj50Z+59GPbT4wZtOfK77x4cnQxfis71M
1ldKjGgUHBD+NHxhhxCfAwngT2cJ2aYjJ3OY8LRnpmSocGdW35j6a0IIXtIMLHej
Kf9blcA/DI+s9WznKOiVfHK3cNt6lHkIEtoh5tzWDK8tiyCX9zFqkUyXSG3s68kR
Oo+zoyiJeXClP33e14H9q5qzMGVBhgn2fQNGQtZH6QHurWFAQUPOZnzM5Zek195g
J9nc8+ZxPRhc8wt4OoQC6vAe8Im2gxxRSFPe95dTQBazkb4G+ydRbvh6DuJdDh+u
kGdIHe3mkXkmSrH4pGjW5Kcga55HldfJ9EJLMsAShYg3U3Mde1bsI6aR8MZXLcHo
jh45e278dQc19zS2vD/6wtp9RxhWqArPpUMGfC8bG4K3iT2bIA4A6p49j1Z31iBZ
HRMrReslyjGYvvBjhB2+fXjYWci8dnexxQzXtjbyObWXe9rKw9O2H5dpcxMb4gbu
IkFbYqMFd17bYgfTs77dMWR6NIwZ7KhBTACZbUgQur6Evn4uOL0DlG/eVVGzzqht
0kb0vmJZi7ND+mjt5BpuNg+slbeEy+KUsKke7ma3AeS8bQYoiRI/g0LSa+XUmlts
mxO5eNL+PZoq4Ofs1BHWgLPTsZXekRVGHIFKFiP2x5VpmWjsTWCmHrUY1cow7zvV
4jYLa05hC0FZ9wwPiVbIjiY/fUHKjWer7F6Y/ZeO5kfPDrClj4JkwhQX+m3e6vks
U7Y0g73VuNwBkPQC43GZojXdWSiRoe+Fh39iGWKY/NzCKq6sSfRb2glGvkQwHv31
4LgIXS3GgBJGFrghGcpKW7+0E0fafXHVjI4qjayMrbyOfHnvBT/vNnfJfC5Im15T
4ElTbUzvjqN+Enkd9EXRlE0PhzvHOXL5ZCrLQzyHwCE/MZVXSqXF7/smbhAcRwSA
xaa8x70mTPV2G3ufZxJxtGC7AYlyh4f1oi68Dx6LXcYmLsaMu/5BInwuJk/xJzSW
SjA01rW9GcLwS2cvuS5zIw3uu6Q26FSeMUaj3GbF+VMeVMWxESYJaBd8QoTB0opX
FVc8aiDz2DLaY/NHC370+1bzXY0zZJY7n3QnPWHDO0+PhSHG9yVNeO4N7LJnEnG8
Eqtgr/XGh7vqcwQOvhtEybNOmms78vDVXhRbotveyMW8DKf0LIOgq7KDQzxSJvnl
jyS4HOWebkqMQe001U2O8d6nRux7UIArLlQZAVhhr7fhwEvdJJu2UnT1ve9ZkjA2
NVaw4wSLKnnsvZLH9zAeiMdFFFVPYFZ8il+HX0Egv8d4ss+Bm7nfRE9PQT6X8tZX
uU7ko+nRnrLhlfFIjUiQDsFWY7XlBfq/CKbGXDaV/uo1iVsv7QrKIXYU8k6gN99n
gi/WBx1Yw21g9uSC85hxAne5G1ondswYAq2l4zIWmBr4NF0rbT6oxoRFYjyt32lb
fJToQC6cxo2ef1UyqykrKsC+bFFSXLmjQD5zm3YjiRExVvk1eo6B6U/KK7TvQce9
iDDN8fDn8AJJy/cGmnHe9rCGTyTocH8jiUArvt1N6TYNpFHJRbU4pky88RwKW5tC
k1LqNCuoQtyYiC/YJMcBZYvWx2UBeY7zulL1f/Q/qgQuud+OH0avWE+/4bxzJXJJ
GlfttXOcbj8UtDp9PH6gpEsaLJhQHVUJoZIWELwyedOXpT7yiz70PO211N/yO6VT
jliNkz9h4CjrHE/aAlYyhsILlwo4aBbHRWkSLf5tTJL8lWcKhkMVpa3vNXMBdYZj
XD1X0JDcatbRm77lF89cinzzc94E5CGSBZcCEuelBIfUpiRu4sFM90eBfIr4oSZN
EfxYitBHMs0rPfPCfj9mcPuMXr6bnLgCPHD9XBhTNHRLmg7ZmF3lt1/u2S94gyUa
`protect END_PROTECTED
