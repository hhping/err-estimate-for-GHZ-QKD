`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vh981InzDvtBkuf8UVndV8w2kP60wYrtwS28dg2eIMKK603yLmXdokvqk/gqgSIu
+LJ2d92cN2xMrZZvwhfvZFux7TGAlNnM/Z9nIzEJ9F5CDLawhNrfWRdGQ/9dB00A
BK7KyobRJNVcPYIRPQzBK4p87XX1+3p/XMafgftOMvTGtuGwaYZ7wbsgv2toTFRu
NPIqCs5hz1J5Dlxd3q+2OW7PHsBkxJHFwZSuZQlnSR0/SUtCFE+qGmly8ILdaXYc
yx91i9rMFWj7qQV+uIoamW8lhkHnOWY1zIJb2zVXENmfLO/zhFp3tkiXgcilBxj3
WKs+HQDVaYvhDBzDuNZMNJfxo1JPgvPEFd5a8e6ZOlT3zdAsogLxELN0R6BWJbs9
fryOsk259T4oYH2KXSqII3hvdSLnVeLXco6XOQIYmPjaa6vD6O64WXeCi9as4a9J
NqJHx6k3Cen8rI1hDNVvKUlEBmXs1+DOEBWxta0zaA0kYzhgp+G8Bn3iuBPYcsCz
3tPUtMqCXmhhkQvBXc3iOUV6KTy4m06yELNub8z/jQ9r4/7hmtNvmwcfd1OSTdR3
o2vzarDvWMelMVWPr2lOTkKSxAg1JgE1z5OnKRPgdWe3rAtI3iOoBZfGHiUQqO2V
+QYk7s592Ll8vmQ7YrNYK66CvRgP+IHh4jsO0ANXv8VKj14JHVtpp1t61h+g8AyF
3LOuw4198dx+GlVy4tIfgcQ/hjXBU0YUvWHEzJUlAHYoCr3gIx7LoiQLC7Lu0CeK
kuorbL2hBMUHIGpiS3dvEeTtmYfY4bvblEQfJ6BmtvauPSl7k8kK9HKGbFpI0FDf
Dgneplf98GM0rpr+8YW7HN69iKLGVNtcqEN/29ITRkUCePAq98vo8Y9pswPT1ozK
RsMhD41zBcwsCnELoNJ/VYjSxNpzC5fqM1VErc6gmM7ot6WJIyD+NsN5C3rNdNFp
Eke4MZGc0+6kaUdKBCj3XS6pESGem0uHPM/JtOyjNhOyZCCKRglvUFyFn+syIfLf
`protect END_PROTECTED
