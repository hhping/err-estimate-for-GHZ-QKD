`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ST/Afq6gQtBOsPsE+ZcazmxknPTvas2nHfcGUd9hMFElAnu68uVJiyxZTVyzKpui
7zrrMN5RKP4zfiCzwwFfk//IOkzCUDBKTvyEb2N86CkPcc4e/aV1EvQ6Cvi2mNoE
KxyJvjAGetLJ6SmMQmAMzyQQUVNXQ2MEHBM2YvKGi7MGmbIMZKsQLTcM7yFAGTXi
yXpwJ75mG3I1NS1CTOTocNTXbnfqDvWKsfxvjl2c4lcKxjMO/MUf+gRuaKhf9CYx
lx4kpZYm/4g7YpldRC7vIejN26M/Ytqv6byp9UmqZZ+QI39Pc3dvcGsDLKc2JqqQ
S3KCV2Vmg3bCSS2FxUz51LhtIc5iCRwE2myvgGRG2Z9wdgPrR+IwCEX6OdNZhm4F
uql58+0nhNHrCzShNPIEEDIYmi0Fm+NdeEHF57J3MRCNfhPTpSTAbXCORRwYbQOR
tYB9mWRzDn1jbgqE3mP4Bnm7+L+HX9Kz5B02KQBenlJSgevQJm9hKih+veE6Bae0
gqz1aEWygwkpoencZsm9y70ThkyQ1GKKUcFtrl5yXWCsc3oPdiOqmXIhP78efFUm
x5BrFdAq8uuhDFiF1KX67sivKyd12cb4I2e25pR7ov9SunGyo5sPxrrSpeRVS3Ca
RFIPrSTcU5tPYnHjpq4WBd0XioJ5hTlMIbtXCFG67ccovt0a/pgRYGhgeJpMlU21
bCEf7ssTi4YPSB4Q37VVl6J41C3zt1QVU/qrBikJIm1MUja6KdFfp+av0xAoWnNY
TyLdFO6N4PuU2bU9RQIbgBY1jKnn40bt0eXArLTrB+ZESxFwAhiNebc8U44cLxg1
dq+4iGzqErzH51VFuteGf8JCwIPAUFS5rmQr1LZHQ+/zCLMFZeiImfY0TyYnasj/
f/uwXhJD53QwU3jJ/yb2C7+QOM1KtooFOxGzf94N/9wdk2thQuvPhGBoF9r/gYCg
sZ24Qq8a19wiNelhwXS7Be8zVWguX1j+RG9zfM9MZLQ9JysZpon3Xbo/IQgVdXlk
Lt+CDHu2uXu5YbV4aTyuIAeSv9GYIayrq6XTMmKXKndBo+oq2WCXtKIAb8+3m9sq
eo5tVP9hVExOvOH3THp1RWqHpM1tTmNh7aTuD2rRROqwuivA7XM4aAkcYgHMC2qT
ZVE3vC105mSVU6NXASHQ5iP7jQoT+/GCYiukdCE75hHBL4HRMg6VPiEF89ZmhWt0
I1zMCI6kLkUJ8ykbuZXH0EIi7M/0GK2tl8z1Cyfs7eTCwp9VSo7LX4Einur8IRXK
FH4XC+bE8gblo6hwVxiwul/LpXoXnLopzLNvRzknln5k5/hjLuYRjKXM00pd/Vtr
YRKflWQou2/KgGZ8MlcoDBSRSrjBoSZ6/D9G13MX2UZyJ+pU1Izldjf3TokIPQBN
WJmXybUk+fSEnkAqIAjI+3hyZUPXhkcdHspOV0f+9YzW0k+10w0b1usofzFT5xjf
2YNRoMnJ4zSePEL8f4+7sPBkX1d0vF5PsCaXUzI51x3dGGQp4r5EiKXjZb9QHKhN
AN0IpKQB+cXAYKLUKIum2w7C5S5wRSkPgWIlulXluLLwSMyDmW3R1VfDbUs2/CXG
0tcoEZBwzfGvqzbhgz+SfFVq/GNNTWl4kn8THBdRe3Jq54EkmG+o8qd/0FmJ1eTE
pLo79qD52LHpotxx6sBk5R6++uIFEGERkJMPMcX9jFxcOoN1cGCH2jxQLjeyI03e
LUcReb3m/nsXPT+OHh7IHdVmjLKRdRiqj6xJy4SNfSmJS7gxt4PXEC3hdqrXjGLz
k7Gd7/9fvcP5+mIeFk6mPMwT1+fsAKHQhxi9V5IOVqP3snCcFMjReGRImqxo30lN
DBfNJtyPPVz0etF4LugLKNYiyZhbe9LVHPB0oHqRupS4wqWJRcUQXv4UrorDwlxo
VhNdRsq4zQ6YzoUjILOcE8dKqMghq1UX/YXdgdQ8ZAe+ebluqjkmu91LRtwsyF1o
i7rbxRFmQxKejibEEa7obRM/nA3zqv6a0ocEYEacWNyMVPxwi4VN79mRSjnhsaYz
In3tepbt5eg2yAZUlIBLl2exMcr9MMN4ipjGHB7WaWBG4VyXxLGskmTrz4qEi5FT
Wq/vYjAOqNb3zQIyg/t2nqUhrciEeX1IbKeNggk5dHBvgtmIw7Jibt9nIZQG9Ud3
+da2pCVx/w1KhANDoZCZe0l2A2gvWrFyKr+5PwyC4VqgxZdgHIfJa48qXcCP1HP1
8ffNBuXnk3rSItmxr2VBkIfLSwomOew8J+w4DeKCJ5rrgB+V2/5yNHq0wuU98RF6
ob4BF5+EeeQx5DGyhhCDnV04QiYJROXi4/2PJ/p5FyuBkHcT0QPLu1HGJG9DXTFp
jGuirRzJKeK1mx9tzNnO8vUT9J77j5oIQGRDiq0+IDqwvQTLxzD+Bxtjv7R55N41
1gE7HZHT8RhOqzIvGRVK4EJ1SUZAcsdePJthwnZPBre1OZa3nCLdxz1KJhKzh3K4
UhZk7o9fjr6kzx1f0TZl6Y2LSW2DpwQRFgR6u/Un1o8K15kkcspp6N0OqwusFBzm
rApJ7MoSioK8xR7T/m6bHXz9XuyoD4ovwqCoNljlrsatQu4nc+NqA+KfKpWJKxQj
GWxWVMmEZnURej6sNH/g89LgVTooKumg03v3uC6LaKuWQbO5lZryBJy+6BdVnk5Y
fCaW7OMLqatHz3AUDZ5soZhoe1+R6JWfK3NX6Z1/sEogvCKuhImrgOpOMHdiRLCh
NfW7H5UoD1zoaCmGG6apgQFRpdc6gMPFRP8DSBkpoOG7uJa/hOU+ikntsqfAkueC
7h+s332GlNIP/aqeSb7m0Xlgsd+51Eel2It6ZmAZngqTnt1m/kputFuPsts6zVkd
UoH2H1qeI6NqMf9jJg/jS1bbfm+F2H5ixDL+fGfzYmmi4HAQWaLAyjfdsrFqejcA
/sDk4SpZ2McgMmQ+dGb9GlpEW57+07OugwcBG8sBFdyc/fs1Fhuyf+parA2ESZcB
INrmTxO+tqiqWswSpDmLbo5bUQN/B2jRheNQ7UfMzVpimQyFMl+TBSGBSVu06qnQ
4NSZ3T7dwe10hQcWS5iXv9z+76rQo4MXRPaFzNxrX2iC3SGKQJ6OShzhw9nmTlGN
lt8bqfPqVQipUfVFGOd31zEFo7wsM6mbWKoUG3rbaVa4W8MzH1x7Pf4/8pFuuPI4
OEdMW/ZUZKXg4kV+LEZi7hlACupUmNFMfx4NOEBq4Jo=
`protect END_PROTECTED
