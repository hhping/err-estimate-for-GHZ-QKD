`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbsDUHMZ2fc/KSLiwLShT4lUd0U6pO5m8IRU0B1NklcduXq84tsQN3wTHsWC20Fg
mDesohcsUVUCDQKJ8ZStEFQmdZ306fIVIlPc669WQXVxFYOzY07cabqbpqLGZ+KE
j+AlQKprxbZBd7Pc27JKWa9/TlVjhjKkU9ISK5UBPZfps19snOUQR1GkmuoldTMU
Ie5tqg6s2NxLD0U/Jy7/sKKb5ERRtx5THOwu9ib6/r/RviOFMsvPNqiJYlABqU54
xqY0wLz+WeNmiK5I0uHD7zlyz+aw2aWGuSoO556dClIc9zGhCdkqvZ3uKSQHVKEg
usnEAtW2nZ5q/RuZMDHTBZKA08CTbRfWG54KaZURO6tTY6eIiBRT9XZzeYSy/ly0
CF3AKxsQqbQOTlrXkl2FJCXtQ9aHHXqotUEBzd0uO5yZuZV2G3Ex96mUZZvTEjhf
1rDyC9h0ZRknRVKtkEsdfRSTcUCQyaz/pR4aO9oN/gapkRzMDL2oh+fr1CSy8J1Z
bmr2SfTJdx8FtHg7FBeYETklUf6bP76yOsWZKGreIK+d04R9E9I9Jj604kvgamL3
q0aIO8iXdSdfh6qH/U6nF4mHvYPo7g6IFFBiqm1CQrfPrfXxkFSoU5BWpbOOy3Nv
3yH5Si6NKC1KjgLRkBoNKhpk8dBYycHZ4K2ksUh0VyJ835Sllz3XDd6B77AWbUu5
MeGkV7xnjvDM7MRNeg+1D0w1Ya/eOlYM6ZoQL3NWEVCUVYuDr3BbPCWzdlr3QcMM
`protect END_PROTECTED
