`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1yklXA4R3SYNdXBTIZ99Pa3yAt1/1NgA+dkHAYVXq9Ogtbv24nOxEu2OHSjUPFI
g3IvYXGN4SiLejV9sNjAMo+4GWKwWm1PN54FM8T8+h3NGuOOqt9VPXp0mTQukV3r
VLMaUnRmD5wRBPLNK3g1HKxsAxEpik+huqDUZZ+TZ6XlYiaJ0D5orLaeOPslueZ1
Y7J+MBA+FoUrtML0kiBmez8wnVaE5oCSw7W9e6CJ7Qa/gntir62UlkUVAF8ODdhY
L8vMJGFwCBvTISIoTwd3yscer0PyH25owW2Czz7IJr1XN0ys4u7sp7nGdKbGqfUS
OUbGRNrcQ2co1KOZUvnSe01OsL9PzyDoa/A8v0mrTOaHiRsAkblmNpaLE//9AYyv
cNaooNBJcslQ/Q2cNHsEsNq21iQi+WgZIjU4aROZIxSj7zix0DZFm0MI791QZZ7d
r6p27zaAeoIfWOJzGiqnv4xW8kavDr918RpejcBGR5seZWaqOzFm0tD8Q5tLZHSc
IMOkoNHtslizJYNYkAhBZA4spuxFSTPXYbtYOFapjvoM9P0lvU+Fstmi01cGdYRs
TQ4murVEFA6Zi0ZDUbfxE9OJKQo38zYTliRubLcDB6dUN/2cYN8D1AK5bqFo6Tjw
t0D3X91+Mk/N7z3oeeSMaG9u5XtrTGf+K3NeBplFn5XQPC0ucQKdgm84b8kTR9/a
6Rs+dxx0QPs1OiYFgORfXH2O/MThUbLHOOqBXbGVKwgQ1Ng4hBVuyAsd5cstWlA0
gEwo2zqL76Rk2LNakeKgIjPxsylWZNMueCkXG4K5V8FUWWXBVeBWAzCZ/2kh78ol
0Vz6v0/G2yyj1ROQ/BiIzLRqhFeNaj4u/iTN0KDJBvZZTeJKoPy2MYyrYemfkwsm
gOdnKdac6BnKjJ642FqcrJgutyZCAaKsS2+zI+8aKMs+QS+331SjhXxKP9xrUEQV
kGru43YHomMEZt2S7/W3j9oIDOKjlvg4yYTYv/wRGNnudp/fNsTIZXq+iOyd1Es5
oAn6j6IY2tLV/WXrldYRDZ6T9mjj/dXurhKEe1OpN/BkgCcHudunzxLTBxHrK6oE
y81xijOZn4wq9ptVriJljdfvwrLUqgND5jj9qHS0alXZsASBrH3L8bxq7x2MrSzG
qml27gytGTigNFRr4b25LfuCfAeQzF5TJEVNHlJp+JqS4C9MHNEWAaCnjy9yYkUo
EJloSbrCmCCDvNlhwerysYQANfPT/uTFkDNi6mhU24Hov3jGOkoPjVmVkWYosE8K
xLRyAfLPLd0hd4sWeCK+9uUvck2h7woBbuvaxnE9poryFG8GXYx5N37i0YwV90cC
U3TBOnLmIVy5+Gf3FQixKB39Dj2yPZOE08ia7eAmGRdHxCfkAf3aiIeWbkzGNTT1
dWp5AKclN0EHKlqj50TyK7pgch0981WsZ6d1ekFJN6x5rmQAfHbeqosVuKKdYn6i
kegKPBtk1qA5oAS1gVlJMrPFbRyxCGmAcnQwwQN6vwKH4rW9tm0bj4uFiXA7V3lG
s1LestCblUH+sZ7oPKdQwtAhwj9N0yGlaouet1gFTabzBCrngARc3iBzG+NHP4dW
dkQ6x7j2Ij6RrpRc/clWnQ4/MF/pgBrW7KsZl/ARqEIq90XcnmQQhVM+KuFgcRgG
fX/aPhNy/kAV+tV+A7dojBjySkmwA1XzS4nWFLNcXciS4OqI86OSCnuU8lewN1lG
1CGi4F0SlgycuRzjleKAu4rb3vKe10HR22bwCtB8dipZYyoEFTmDqWxDSj2obPCc
H6UeDw/+xBcjDEg1Fm2of0cM1dPdEEdXeYXcLF/Ny9/VHoVgBXmhi8leVEmCjhCI
CvsToPqNW63+xnmlgKPJf2XTmOsUI21ZqtVIEiu4lWwEHbVYj1o8ITlORiz+Hqk6
gZLWJlcTLmUMb2dRFpHTOY7W6m6PHJ6KVsdf9e2cq34ge0xDrzytocvH9NgzraUJ
8aYX40eGIcdpeWSwB7iFHDnV4yFHm3Am5Q8p40F+0KJC67Lj6toaJOtcHPt3Asx3
jsbOOOQakWiGKGIFAKHQctQE+6P9NGOsAB8WwNbxA98eAWKMRmpA664qAMQP8aY3
AUJZBoK0PtlQDyH6qr6Tsn/lStgo+iZUoWF3ydDDPtLwnPJTSRa+zhNtvrPzf9wH
/y0CUrjv3jKA+gG3fvgFLX1UjdppIX5TuiReIQY0MakRtOGLA/hQqJOEJlr7SQG4
fUsTnYxQs2nt1iOJ+1K03VxinkE2lZEp3BOZa7b/+CZxUr86R3FlKF3l9Amt3foD
49Q935YXT6E9qaMzgFOpB5CGxwi/FcKpPOxCdXSo8Y5MCh20585yTxP/sNaukSqA
eAo5zQSKTwBrGyiq6aIrfXB/QJC5NODUPVX2/YSQLZtT9vgtczfCn3RWKEmj1aOA
xVcxyAPHOi3v0cJtwAH9qeY4Jzl+WBQWWU/KlaMYknv/JagphAfxNZwKBJjhXuVv
aU/iNQF79WZ9MEArF9Y7le5R80TovzcULN2zyDrZOwPc6g+rFSYes5H2Ld3deV4M
IuJxxY1QYprj1DNs2H5eP7rw0Yoho3OhpGori2EqNtWfl8BSYCyTgGR9oj1+Sck7
9OGVukvgL0ScojBzjN/CSn7jh5uyb8oiHx8L4E940yqplVdbiJehEnBlKayPzoH3
d09nwN/UPq+453QpszyVqjkypp26qewWg+yXhmUgMn1vtKOLXgyFw3MFluubXOy8
CpdFF06nZQyU38f5kGMOplmNg1eFPCnNqUzSCIT5WS4GPkOWwXfkVCNUoVx0dfyG
QLBzflCsM5wOsf1tB8vSXU76YNTXB9riql8OtvjERCBQD2fg85cBJ9VOLiOc0s4b
lSy+yJFZ2RXNcckYoZyrRuhsRLaozZkTl0tZ/+gyd0zwrqKr8D2GxDTbmhdNnJzp
l34BHCToCjjYiSRJswhIUcjYrYWvYOx+gpDKumhDd4FDAamcXvwwcdUJs5X+HcQ1
08G1ajZSMQr2xILn26RjCV/r9qEyOQb1Sf/OWxCmyNNAz0bLbQVgj/wWFCVyxl12
p6QAlgJhDUl52/ja2JxiMNTO5rZnNoZ/HGiLZpJmjWXJhleArNCRfIm3WM8f5eoE
+Rf/+nYxR0ZE8ODPxgoZ5drQS8NheABJ3vwOOa9Sm0me681DJliRgaatKBMnjfz8
uqxyyFPJTYcQ7wXYXDdCSTvwmMB1xnBYpectEZiOawNRrUT0VurLjcxWW9wpRnTL
4ThnH4rLqPYbjhkSXp0PW13tOmOnjnuA7rUyG/gT2bS45u7P/kjh5mhwZl2jU3D5
gHrHdiRurGsWUGMZVupI0R8N3obgTTGFKjesa0Vi93qyvZ+JsRYVK20BxNmpmcnV
pQyg528ArhejY6oxpS3DKA==
`protect END_PROTECTED
