`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dcfxMglj/x+FYJIHPekpT32ypgTn+TluWlADdvRN7T8Z7QwuN6QqkeHC+k0aty3
QAIlzD5Mn8uOsCJGYPuQDhdJsuSve9kwnaBK+5f6x8kc2r+UUsn5/zH/Q96g7b1a
n1QRBSTZ5FZPiT0hxGyo9hKmINDxDAefh74/aR8X5G8JeBJwA+3eNjsJWN2BOVJY
Qqvhd5gzfmx9ZVL16vUDRr/As7wqrRNkp7OBFO5EzpqZEPhieisfTPSnp3R/LTeK
6Op/ylR1aWTJWCkdAXuMF42lz3lj/4rlGZyfK0I6WP9O8vQs2dPjdg/Z7fIkD2n2
8n558LcWCxPBY4yzW0JFqe88aO+oAbOy6HH6t5cMErnIuNF4IOa6tbzrErUIbv/6
OokcDyCLqhWdJy/3gfQ5xZtSxY/CAltD5XK2wA1pAaqd9EEEFSI3orj0tWPKXX8d
M7k2x3g5Uaj+EkfGX3ma8fekYqasz9L5TxJUJujVJFWgBt7oA9981O08Zf6YYpDe
ur/kBZENtWyBGL8lYj1v3Vc5KnbWND59UHzP5ipt9bLKyuZhECNkPe0eNg+zXiQm
kIBHzJ8drs42Ko9RedvZLec8gIVH5Ifnw4N21r4K34D2mliTXiQrBhfILcBKtDk5
oMv3GefBM7dfLxH74IlYNp3AcBkD18hLcYSItzMUq0V3nOmC69r7RVFuTyqoeYaG
1pZwY0+z/TlMk9KPywU9itcrONnZheOkmOz/Dk+hGhvGWufq5e5lSIOg0FrrjL6d
1fFIAEect8YGIRxLVH9Gam+kV07orRiCqSosMuB3Bxd409JJGBmrvtspadUpXDhI
5JWDNNn/FeIVp6CderMrXY8klG4K7hn3uHKHiferFMJWDaezK6rBKzQqYsZIhzlM
vmt5A9j7fC4egtsU1qxtSQwKmz/Xmi+Ie9Ai3nx/qIErxw9k9Jxqn3lrEwuC+24U
6j8V92enZXKyyavhPmwPYgNtBA+AQwdD3fZHn+W8WXN+YP5eZugECKLuY7KExm/7
g43X4tR7Mo/wGJPQZX5Nb2pine35gdibPC7WdwikDFgeeRqSd4eyUaAKXZVJ/AEk
8aUK9JeSuF78ttu6NaM3lYBvFxv+f9fZk9+oMCtTs8Wi1ovtS7V0SWuuwft8VQv9
JDMFsSBPqqohh66vih9BPUfb6R0kIyL0DNpSvMurpCTNCegpWdmYKkqUDvhqUB0i
QPDJMh5vzmNuBM/6Z3pJ2kuG0LxOhtmCQcklacZA0EEktvX8XPdW7GGqmlZPf5wb
qR+DxHS5JT1zUnTGEUYOgnS3B/ETFyLRYx6qbrhYm1nRd2BNWH8/OsGrfRh8FzJl
aSk//D96t/rZt9iFtm5ubpbs85A7YqaEp5qg428oL94nyOaRTsUhsD29qPys9iOP
VgUUxrWOe1QxT0DAESu9MFHJbjz8mGd3w49bVywYaAQP4+PRe++GhMTUbBvjb2re
RBIyQoJSqftpqpIhWNfZGPWKMFQn03BNscUTseeM2/JHKbcGaV4QffHLm/2Wqqs1
jwhNh3YhkliJyrqY8OUZM5Y4sxYEN+/P/bypnyTGb4xST0eJqAhBjAbbNPA/TWKW
sy3cdT7WJgy2OKlHPHV+WcEbhNTrKuyH0ZHHxOYxRH/iur5Dfj3RbveRS4PTdLrd
k4DoGtR1CUtKjQ+Ztu3JjXAhtq4+LiVDc9RzccWLjMi6M8BiSDoVMmUJcf+5wmWd
iYKxePtlH3gBQaeprzU4ysDXqv7F5rF71A4gf/QASTS5lohVwi0B/7bs8W5yQRrj
bo5aWRWOVSiGeIzcBiwd92l0MuMT5P11F6/LcbZZlkrX21d4p6ie9yTB7XfhNMCO
14W6bdtTaoREhjtXeCW5dvsOSqoSu1mEFwQ/fR7oODOFkfVWq+3e8nxXnrtoDocv
ftfQF9qUcBPpzqiO3bziJnqlFxpQDFKzTuEzAj08SMJxJeYLdQZ5FtsikI8xukXw
AAvoB3wNmS8D9eOkCxF/081mdNxCeZnXIS542+UZEGuosfxKSKRrzrNlXToo/h9o
MgkS4tJBrz7P7KiRB86jdYo6D42DPLPIDn599JWAF56IRe87aeBzwSmc9ttIASjH
oOMJJiIQV5VmBoBujjn4Sn6B2f/N07qalhvJzNtyAt/gm1AGrPls0d9UKljCPlpg
sz3unlGSZLj6QQpz0xW2fMyUWU7yhjo9VQq7TxO38efBpQLbR4TV/g7f1TLkzZFI
c4lvxuakvrmuCGn31OqcKMke8ljFgUrLmpvQGsduRdWaOl8euKzN5mEjWM/4iVue
9FSVkY3KOa8pR1zZGXsxSgNr3SW9N9KsP6nyPXuZVjLAb4KGYgK4OAtL6aE4RPK5
7UnLJbJmljN6cWaoaK+pMjB2/5umpuJFR1Kod03R/YMS92Hle9cxK8/6kGnjl1ug
AC2v5Q5YhOPCeciz8JUKEjHcidCciV7Ny3mE+IhqUu4bUGspb8mhRrXx4oWA2o9j
vjpEe1D5Z78ZWZvT6Jn8eWnMx/c27etI8TAxE9GPXWTgyNCHbDROu9Kv45E83luI
ClWThQ5yHW7Pulm/L8cEIwDkoEDJAzlbG8Rlo5vyhSCDeCqdRD3FOLBqoX5IUXf0
bVme5fpf6X3MEFmhXypaGg9wWvBO5HqiMjju8chxEOCIBySFIPGPiPdq55oT/ZSs
IR5mMkxhR3mMJXzgsHhXIlvTjxLEjTTvZCCYJ2Rm4Gd9AKEpZpBwQXs/qm4mUkyo
8Z9lWmRpCmtDz7gjqmbFj7pUyDm7GzxQlyqI85dD08Z9qIs0wiMDuLY74Ubc+YXW
IMMkk+0On0IJrXhe3we96txR1tdfMpvB/qqmrmMvHGAl7kKD0dcqhFCSTBk2U4cT
i2zF9n2/Bx2HTJniif3I/O2777sJaG0P9rB+rUl1d0MAlQGgqL1lv5itS38j5wma
4Y+TNMDe4rZyQ9JvZia4w4sZrQaQSmHO3XYD4EvWQS8wjrnJ2a4jmZ9W75DzBxcz
PnrhcNaDVLWo1YlCCDYnZI9WmQy4ClSRu73EevYOrbIXtcrQyVhVu0OM6vSn0c4z
Z3q4dZlw87E3IfPTNaVd3qiFn2zRhqSH2q/VTox1xjQS5FDoC5Y5qB6mj94FR83z
5RMpXs37o4drmaR0jsVF7DtA+BImXmqJFTpQlkkVx1RH3egmMp7UQt2IUohBRuNf
6/83DUv20bsAY4flFvxVKvgnwT/rXTZeT5yL7HXg2ap0WiGcjrYMAs/Xe4S64TjD
ojR4w53UOxrYiNdyXThtsrsBPkdUCAWpvSxP9rk2wiuV2kNtn64K58ME3rsbXlry
q/jx2LepWWpbFX23AvJtNJj5ZPep9wQ9W9KsXt/y8tLVgl71GXd5N5GxQA4DtOQg
fYCEV8417kQzr+GuspHMBwCGefVzLcd0QFVEk0m9U+qjrcwuzmJqaEhIhJTaFboQ
9GrEpF8N1MyBL2MTs/vmtfKMMCDNYIveCi+ui3ckbW3PT4N5RybD+bfIXNJgMS9n
aBY1j4/JtlCPj9w+dlcl2wp5fb5rxRUhTpH/IbT8eEFzI/1uIpX6i+6vhipH2JVE
hveYXbs5bLTU/LkmQwyzYmawgcPYQhudEb/zR2ZkQ3ylfOUGHvs8nhI7GQjSvyrI
wXV7NVtotX2ArTfRJDv877nvzyPcaGFpd4Xf+seCP7vSQG1hYkObe3jkN8hyFVxj
gJAHv8Q2aCwtnL7Cus9rvD20eEgq7VNz7crhP6mKtWEzNvB13XSuJt49jhngYfyf
1oW8qJJWDSwTJOTXF3qjxHz+F/QupXxop2uyA5Be0CDzJQ3FbZbKpMftBZJFMllz
AYeKxWrVrhumMYIa4bO8Voj4QWma8n67nDs7VzD2fG5WXcoF0PjNpYvOyDwwwZws
rJCjKvmmdFs6ZikA11PJYIuT/GMf6hDhlDMlftLlmc4NQ82YiPR7TPSEhQHvMyyO
ctJZQPobBAcQL53a96lO6g8oDSJuBUPJaJ/2pve/d1fHQl8npvTYchnmVdnMHvl0
dTbTNsLP+IaB3QytsXHw3LV04eKmhw2USwWZ5raB+K8xDZXCxsxNwU7RbciA9hBw
vFgn15csRm0wNDbVu+5hFRqvS+wk0sMr4+/2tioxXZM6/shNRkUn7XcctIrM5msB
v2iPBmXpsldRqixmXbMem2gr2lPoDTcnx3+NeyOpxTlYIB6lfxZxwi/AYlNqht6+
uKu5nAXNgLoayQV/9tm9e73K4oU2yfE2ZoRhNR7t+P4mm6STCu5Zvz4b5jCuJf3D
B145Hv1dxuoeQrDDnYpfhp8/I7BAj283tklJECiutnp29V2x9trotqQh73c18l6Z
EARelBIH5GKMXvcSvgo6CF2LfXccrYUr6LBfKInUyAsOrq2DBGb75sNlFZI02cuf
vLxlQXn58M1ZbjLRwJZnfhOLuRNTk37C3ByMVp5DDglcEAqJtVwfIAPSE/iuPZ1g
kM5kX6nhxb5CufcxEE0boNNHXbJ8D+Vw1LxSxJaDywGGfmKry5bXyKHfZ65F7XiE
aZ+8v7LvUAuX0/IUWQIDUPzfMzQ6IlF53mjniB9X/YSNjk9ODQcl8Fiwg8HLzpuq
VJChXeCH8N+wnE4NITwVQVJ3+zanhTG6PnpEwl2vToVSKIPcrddzHQlR4m2d/9or
sl+FPCS/KdmbjZUtv4+/WR6FKFA2iwyKDYo7znB62IcCAwUjCEjOyjufqhxmYtaZ
YVPSXAM2jYIwewJMtqAAdkb1fNEElu5gNdQ/LDWtdBXfOzytBLx8IDPrzbWgNyA3
KTs0sSSOEep0+yEZcLqPLWxrn5UCVMOW4f3kdj5ffTnkiRp+oCzOBHiXXOkzg9Qi
QBB09XovbESoPGTv1Ui6G8xK/yKV8mlGT14OuUyApqm4keYc/sgXdKvypaj2nyY6
ETH//i9EcicPsroSiMCtLTu9RME9negxZRDWF3HYuTzeZBvcwP1PacRpUPwW4HcH
/nLC6ipiRTm3SWXCT1hP/ONqHJXYf9HjhtAwCE+5Ec9fuDjbDrIjShf3Php2/vvr
RQm8K7aKLcSB890SChlCYuyXgZiZXwZ16CkEheJsA2owZC7D6IlA2/lOo0xTvCH2
MsHxryLwMeyMStp9B+ItQFFZ2HPfEYL59B5tqcL/H58nOMmKv9Tyu4QPOcLIzMFO
jKOi6jc+cAgBCRHZW7UkIN+C3rkvuYob8cGGEo/2fHg9NqMIZPDFpZdLnNVj7GQb
BNESZOHF/r9l4kPXrwWRarkT3beoDr1zZ88iwHlPuLeaWKmkKgO960E9oDLOJu+o
sNxhspHRiPnllSpl8Xzhh8cZGjLub28+S6h6pZiaUYHZddi8soeXHS/xaYMUn4C7
jj4ppn1BDFGTlsohZishjCjwk2IsvEiQ2TRhDXoJSi6bKi08IqCLBSDxuCHPcxn7
9uZj8VNGSSrBaObP2V0R754p1IV6KMUTXzWb7NwIzQOsV6dSOmQ4Z9vVVlKnAFo+
rMDIhObwkA/j02WqwuhWRQ0Rw1E0MyUfTRQTkEETkX3zOZve8u6WtqHKUsP0AkHr
HMXEGUfN4Y2So0WBdHuw5U0LxcCmfTSay0OKdUyT0qBgWLG5GBno8tPip876ScgG
QhcwQMG8iXf2kRlfdsRgd0vrmCQLRyCE69IQXQhyzslhTY5z5975K57sQ+cppZFY
U8Wo0H85QcsRxiOHvZSLM92VlwJAS32cmXR2ctogC5H7UQd1JtjQcXgvj1/zJIgA
ow4qHUh8WYqmhydjedJydOBl1RXIZJX16KqUF755V52x66bBPZzzwoK8gNmbkZ42
Xa+UfqaV+mFg/WrGdhlEPjdJZJohujNvPUCAXk0PAytssShp5HCYoBzIsJaHpmNL
pUcn7cwBPZQq8bRqldx43YzFzFzo9rE0bThr37WXetKiYFrV/5RhTjmP2NDrawXT
Ghe9VFRx7HRxIAY8zeCmmpICX8H+kflRWSPY9tr4SzwyOjrIgT5sRvJyW/UzXNEi
aDNYusOpNTW2EGr+LoNmdrTim1Q7q8WG/291gUDrDm50UAx9m0UFMaQF51vqXuaT
J5fM6xZeVwBNDlgeaKh42alSc495KXkqHgGkaoX9+qPGZz+00uoIiBkYZiiC0MGA
pNmYhA1snwVOt4jdcNqXMuAs74sjH0DbKSMNNVo66BcAs9EovCfrbw4GZlMBt7+7
MjYzeTbwJABmMzjeopxSushWx5NP299LNZFyGse7MKR0LQ6owKnXFTNT9CII/1gx
FZM7wPvfFA0xFFr8T+/dQB31ZZcDhBipuiiI6vFZ5cVy7k6tswiSfX0RbrD3vD0X
bK2sMnCj+03j65BmPvBq9jw+rsBoriybnA0o1jjiWeJSQzdbHPTa47c8J4WA+RMi
UW/LnjFalVtIrrN/6+VwnkepbvC482FrcIMLN2FwG85LLBT91Y1MKk5D6SbmTG1M
SRtmFmkKeD8ewtoUoJDlMbYwheELMDdGBuz9/J4swHApUlJuo7m+hobWrhZR6F1V
Poas2EqwOhv+dpYaj/1foMXoSDmjQh3/Yz4/jEjx72i1lY90Qr3eZfxSs90A9Med
V6Fci3OsgbZWDccMgCFYoftfIoNRiJzSvTwBn9uTVzA/thOfH2YvSqJ9ew1dASHU
+AQqEKXFsghe+h+m4EoJmA==
`protect END_PROTECTED
