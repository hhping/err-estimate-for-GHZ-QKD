`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpCfKKx79w5B3J98I3J+1FQgzwRub5vj7yIUlJeIpJtCxjSMt/7tkTaGPtfrjOzS
i2FS0bymdpvKznjV/IVouKx1gJjr1d0Y4b2nYKKnTE3i3zewJVusP14dP0gN8BQM
nx2tFWCp47vjhrvwCxt+vvQMBlupxLsrO5zCe3c6mX+sqjw/mL/3zwqO6PVg9VGj
hCKsquiv10ejSCS8ysxvsquKEmqcc5JWjGlNRHnGDXLnn3++vdHRBmDm0EiYlogS
jJlnE5XeJSiJ/iazQDZ1NUflr5oYCinIAqLy6d2pbnwA9DP8r5crScnMH5yE3CeV
HcHZER50IPUNjOn0HSMHTqtpbgqckjrA/9aoJ+bv+x4Xod4rpkVMRGIio5IELYkc
CjqWlQ6umpz/XGwtwkr5ZFo9ArQ6Wn17NC6fbQ801ksQTwb1qn7jzPKcQU1UUKTk
Nb2O2TcuKWiawFtaOi7TAfwnwL/TnfF9WXMokjGWZYdV0Lvuf/RE7Uhqdzrp+qLg
LDsu79/kIijxu+X+KIvXT4KyLn3y6gnt8XjobkV2WQId24JiUZglh12EgtgKgXLa
QN0ZQExdtPunvX44eSYY6v9N69XBo32nG9yq/tYA2g+xm1/Cf6ZdPj6hhCV5AWOF
LOLgmPbhAWteiZNzUUDV5rK7ZiODtYaOq3/24TkrBV5ZqUECCtJutt9dkbs7ZLqi
6jH1uSeS3Gh6wafzbEfBNCNi4R4rVH6M/vHbdgbT0qFK8NmdCiVPfEEuBDmco2fQ
Dz9Mb8NZ0VoYxVY9bsPnTn4u2zG09BertFKc/InwzC5+xz2P33jaA60jezKVuB+J
gJYSUnvBjtGKpCrrr5rMPO2SEXAUdq8s1KH7R6H6bhpBXDscjIKMNC4YJcGzkskG
H6JPIR/BHfEUYodCC7+hYoiIHZDffWZzFPCo7JwbLyyQ3foc3dZzevWVBWnWpwmy
0iWH3bdT2QxGAuPi3UOsGgHL5xsU3Dfvq2greoJj9e3yMqp2nr1rJIrAWakufv6a
1qspKzv6Iydd5Yc2fKNTE1XtdaYGaG5ffw8Wr3v9kgYKHEjtvXIm5Ks8eCSwFNgG
vFrUNPQXqIHrBHN2/3yheddvki40lyPTYSKpR95RudqJX0v5xX16r3d8ruhmVStf
uopZ1VUhZooAANvnYRyq+rF5fuqJRPPww48eRHdZfAj2uU3F9DriQezNsEKKEi0A
mI6Z4tWQmWupjm+zbWYb/WHH0trkD6ybKySAHMP/p91pwu4D1MaxYa/QcwmSdR25
HkDI3Wr9WH1Z2MaVYVsmOsMHWTmu2vduuYL4snROvTJlbcYZWSryJNnqVYqD2Dex
feawNSSw5xOAbYRkCbdRuUXOpX/WoMcQulo7dESq1WmmC3cCZhGQFogaYxabdK0p
j/4fJbwSuYgYgtxGLLd6DvY+LdZwYuMvjH2WzsBIjDGpqIyvUmJbO4Kywnnd57jb
uJI+sVFLMjBLrxI6FkO7aj5CaDJCYlNJxArv+ZJkmfE=
`protect END_PROTECTED
