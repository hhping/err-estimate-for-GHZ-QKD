`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXmLQZoJXFmsGFLLcBywCho4l+YIeRQZ7QuibW0Vw9g70PvdwrByKp6FJ+MWuEmW
ybNhzMz3b/8G2K1JPWdC5m16qEKwVjqG9t6JHsiQI9T9Y2daBbSpWYgGo6wcNBDp
KPn1i9gqwvL/oqJcV03JoxRwneGl7PjvF1o0POnDwMaSews8DcK8ja+xZoP7txAi
tdE2JFNwDhuOMPOkuB+iLx2D9nTduYybif+oMdyP8pEpDdB0E4YFkwrURF9RiydU
XAjsgVvug0P10QGJwzCFeRMo3WUSfBUdSPQgJFlpBPWNzZknbJia/iP+lRbW+vxN
Oq97TpwPmQHevVQ2JDxZowNXfii+a0lM4PLBDU+aCOopWWJ5Cu1gmbZDgRwOjo6C
wRSVIuIDbaoR5jZrqeeB3UiLrijrLVnAS4eZo6z421uAG7rO+vsV/GpyqLi8k4m+
t/kSi+JfsTVykkcd/AbQBiISpvm8fc9Qzwx/AVfFplcpEtFWeR5ARWFjYSuWwYPD
kj+enaF9fG9L+BFl5U1pRQ1ZicoqHZSZbwqcaPF3lELqfe89nfLKazknwW4ITt9Z
WKTjuxrtfLoYO82ae7uhr0p2pUT2XL08uWDfOVxcWl6Mo3ifFw1phAP/uL15mmqB
eulLJcDwFl2D6uU00OapLOCJBOi4Gc44mVVqtWhYTV1LaAdbKI/FBAU71AFHZjee
PYlVry1cXlJfI0D/Wh/AKFgf2Mo5+rh+q2HO92zk+AyzlSGOGdjffQN0z5Bl1WsV
jYGij7m4z0MBHHiPMpC8Mdtcs+P/cuc8GPrYrhOdvADLHla6BekAqPmR+/sCOvYM
+i9oQZP0GtEQtQ21YiREFpk7PVJWOnWyJYXJtENvOYFQ00E6+TBucdD3ghjvNdKA
LV9bqFualjtDEspRE+d0c0O0WTfAW8WAbKNroYjzrnpp6/vrZqJxlS1pzDQf042z
D3LwDXPBBHn7O+yKRK3qSfyfLCdCSWxxpiVqbJ79hoFPeUelxHuYHeYDpWcXQ7Wt
M50vX1NE9ik4AqSFIDNqX6H3MXxLzDtY5ke+3oCNPaY8cFDHvi15JezsA4FFH9BA
evORhhSjki3iQKjR14J0n/xdquKe4TTuUzvKp/Mi47i69ejUSS2nj/CVYseyKzKq
fJM0LFd9SISHtTfPtd3P0kzbr6vcQNawSCvAzfDLQQrM4t7PB/iYJ57ty8zc89uG
UMsDdJu596yo05LOpQ/JAKikkC8lNh3O9cKS+QwIJOH8G1g4MoVUcNmSYRalIEwE
RJzu0nRqyVvZbnYf+7FlRVzH58UZI0hrLWXB0bgwi9C0NE1JVADf115SCVbicIV6
dGooyJzvEAzNLh1itawHu38XWshKTGwrlXIqAquor1Of17bJ+eytDPave+xDYHyX
HDl/ix5htHhfomb066orr0hoiutrP4h3yS0SrzAYM7TEAxHaTTsRcIyN9uUY7UHH
OsoGoeTB5gBa/y6IaiQht21CO0/4B7n3IFvcbCLa6EBQMshucOf8+4vDFuJ6r6m+
3BKTsVYVh1UOZK8cOXOoHGmnPEYxBzzJOJYBZb4m4g0sGtHRz8QISK/zKWIzl9w8
8b21wMHimVlxFxG0G9aRq7ABxbfhCDAbgf0Tqw2Whi8qojQC/keA3odL9i1AnQ3f
iIZyPwleCKSdOJwOUGxPSa9kd3RuSEQJP+nKeY/ZBnMZcFry9avCeRTRCpjr/Qlo
MOiJCW87KQekG20wnvRXb2lw1T7R+KbwWZN0E1mjobK14mr5KEJo9CNApj/u1Nxq
9CbVKgePlQzGbrad2cTkjHu9TkvUv0uBpwUZBwXAzok2mxSoDLz/E4mC0/pCIHA6
VL73FBjheV/4jQkACfR8uzvsTPgw2TujRKXf9q7oW3HEqt7zdKG9ISjKhRLL/K33
ZT30gb3qIOHVOxcVZiO3NkCA6g09FGXZn9a1v/iyVsm9EyGIDpFaa+xr1o+5FeeJ
IyyAlVCYQhyhSSBZpfsuIkDXiPMaw7epVttCoPiLLVSjdO49xgP9wq8eow+aM2J6
Q/YYZRklZQR40ksaQkGhXkNXNN3WmSplXT3Re1zAG7J568DmjVLAY64Rjc7Q2XgI
Ugf4ZMUu619VD96yBoFKKNweu57aEn9Fj1gIIYAOt8Ot+xE8lNLrNpP2wGltBL2d
QMXy3E9nU/NG54jfkT252LSqUYB5yEBFrGdepp7bUNnrcUIQGpYQ/bqNmD2WA2/V
pv4LgLM+zO4BAogvFbDG3bO1zNRQWdPoh0TXa0Me00qoxSHsAjbhA89/2GBzP9Fg
kIfqVdir1euy+NSrdOY/XCm7QW/2eSoDSZMQw6QbumPyOiI/6ltXJdcBCjLm4gd8
LJtq6fKWQ/1ty1Sl27vE3WEwpTaRsbT3V+94Avt8SBhKUVNsjhYWyHzV9LYiFog8
Rpje+FdHx2P8AK114K/fccg1oOmB6VKeYmpAl2t0iMBOfrUx3lL4z+hrnRQKEMor
ptTLAzcXlL3pDxpA3YHTZvQd0FInGn8Mwye6WbucADWibCFv5LAJuvhenS74gzMM
v+JOM83xOpVLiL7TBbjjZNQDGEfAjFmIbnaFba/LDR24mYsmwjxlUKqpp9bti/a/
HflH8EtOB+WuV3Bs2+sbuNdBGvZnAsUii/LszqAvCHFkqj6dBxmLMmK440XBqg5P
JaO38nkZNxDjUxvGvBz0PK9aJ3ccoqsTsd4k+vMODqaoIi5Vzgm1boPQhH0h+L7o
rplbgfTQKbmggaO5nfF6b5yVhNeWf7suwlD2HjrF1D91Akf0OicRMG+jstRVhe3S
2zzNxmp8h4ikmgz8DtKsOPZB8FAxpOX25hY/uqI3nMjSj+6pZvFK8kQDAsd15i2D
UgzVmU6IE30gaRkwO1jOKx9PLiCmo1qCwelij3yUXqZ6vfJi/nVmJvVxfbg2fNeu
EAlvu902fiZAWID8YfAXpb3nPP3nsXK80VHyglPzUwLHNYyATnrGGCCfSKBR/+7o
Qj+cnK2WENv2li96VrCymG7Vddcb+L56HWJzpi2VsKPhcJmrxpuEfl8SXJCKNwTt
02KCAw/F6wEx/oz9o+Pb+ch1XkV8oIBtDkGx1jHq7eYWfVtQFlfATW494N+8Bkm8
7saIe/AZFNBujGIXFuj9SNFXa6L6v40doBlhyML20stRE7RqbwZ2BIFf2UgXk49G
tMMl/4T6FKwjzRZgUZ+UBp1/yySY4x0R4DyrkZe0Cz53o3xvYeoirKjOtkwHB8DS
xGqi3NDarB9pGSd4I4FS4K5823L4OqGJzHjkQ/zDJVGNrgmfBehYLcP3MwMYYODz
vKNzjURfikvIFlUuzz7kWFLAQioLUDDQYben/81IK7FDmnD2KSya/RWPrg4WSWY2
emrUCo7opcGEw+ua1iSna0liofhTJ8oZsXmlOA1F9KcgSkN+kPe5C+K7GuRUnR42
`protect END_PROTECTED
