`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxowJMLRnEA9I/bHsKlIwUPPL1jcxcPgOYBgsqvrW7mlaIMGggJxqC3WzgsxU5N2
zYHBT9TpVMXOFusrp3XdUxY4eIoW5r7vP5jZ7Ys/Pq7Ik87eQ5PMOUrWQdDeHQKi
tsKROGcwaqzL+HLwju6w1cNTYeX3M1bh3ynq+Wj3pdayA4HuXOf8hwGNVfLfZGCM
zkc9wNp6vrERXQnsD6AFWRs85t/LGwK2KizfGatJWfqGqyEScm/fDmBSQfTfAi1n
JZ291PE9NoByVkw4m8OmaGVj3Ud4ae6eMkVoGhzk9LXxsSgCKTiOC0OrNq+bOlCa
Ydar7kyaP9Udt8OE0zS2lzzUVFnHiOifM0+zmxo4Ecq6VdQ2GumuHG3GKGvcTtLK
XaGmymrErSOF99vm7XDohddcU1Jp4o8Zh7Ir1SaPsIBDT3Un39RzkEDnkIV3zE7p
iwACIppTdnZWaD6pC2/j2fou5HTy/M1JDU5VCe2+Go3lZ97okwtSgAd076GR9Pmh
QkMIN6zq3f+n8zrjVm3fxtrcuh8bGebPPqzPBZSrVGXiZF0SYy48ksqSU3onb151
EmXWTglg+dR3f56HTdFrKsxIMi0ORxFkBrEuDqOwVI7rMcrzV0K06+1U5I6LWuu0
j49MlsR1ID+mAmBoktryiU6qKwqJHK0Q/yMvrrcvcLNH46jzfxXtewtCBXQch6sE
XW2LAaR2Gth03RPOjLWnMI0m+JlEftmVVc11ujQspGSM4cMiNBzMzGc+3iSg4iiV
KfvKQcOQ53/OW69P0uYZLSuuqBoS6Mct43Jt8AhElAvipOY/VOKBUukr24nwPVWB
Sp4KpyAsqnL4vDzL1a4X1IbDt0B4I17NxgSJXedrZg1Zl0FdpO+moIxW5Ebfibqp
spAStV4aF7cvK3yT/XvIbw/xXrIl/jVlxXtE7iqfUnKOL+FqUU0yorTNrKv5x/94
aDeKdiDly0RSTfdhZUdCZuP2d+bbkQa6hNuHmEWgNHz/+88aOVVt/x5SwEIVZYDJ
rqjfzVrX5l1ivPfr4yzF8NvrHmwa7IcUmHLi0qbU09qa9/bKI12OWtdr176rxrRv
nbAQErmElNNYBHSDBf6hfPvX9S4k8u1/WJKNUBaTm6woB0N9/HbSBDUVhadIEqDe
w5icWjOfALjauJJhxGpmHxiPqSKtSefKqjNGDhDWUPEin0slQjYQHafZk+0rNW6U
E/wd5hPRfEaL1VpaSE0eoZVLPZ0jL0aIjC4bSbiA+LLmQ4gA5nY2euUKu6iDwvxA
DPvazC5mPU9P9qMifgqiT6o2VSsJyh+lLSiavOKw/wzQvGSuCbWLehPyxAhf2IDO
gGPU3D45cHzUgTNV/qo2KHCJTmBmfkixb0ctHe7gdQv455tamfLlgV+aWPQgh2E0
eg8yyYw3oY7Hl+c55G4vIp/0sIv0ODBjrBPkX3Q5NMa/VHSxNOQsUq420KwD5zvk
tBsvh3hOWOzO2O6LQhwsQ2PL996DMvVHKPplg8UkWfdnrp3nv/UHIyFjzzNnxxrF
L/bKIWsClshZmlTpWYjHAdhAlmF0BeblYsOT3Ac63FtV8MZnztr43G9Ks4xghhAh
BhemOEfwyI8gG3jXugaWv8h3Z1lnDtr2ugHaZmoI8EJO68hsIZLaVsjMzBeZIufC
m+Xt52VcqSzz6w/51HFS01ug3jHucm103lQdl+B9LXhjVNp8g4QOsKanSfbc0Bqc
/wOqeI6vVh7xHgxJOt+jxfHKxB6AJiwwEQwK7obVR0SmugCkIi/WCbld3P2AP1Ms
dAR91DQNMSfvFRcQ2X7Kh6TeWtHCDsMdiLHPR5OgOBbZRbpCFVk1JsdD0E4w4KFB
md0EE1UC+EMgsr+xtBsb6rATXRZl6140+EE3C6NIcYAFLkt1f3hBmtjUxEHENdJZ
VLSf9UMhd1HDIFLkmIK6aYmO+3+mgcYuhhr1FDRxBy48KpmSYsptvECEhJD+/dDz
hkQGJiYgeplsOcwBsNYyewfQLeq7/Gprore2S5/Dk5rAJxD/2SRK5RWTb99kGnfS
CrXVoBDWq9n8Bz6WNFF4dN0V7XkeZ2ct26NtmxlfYAqQgKLLHngYQbfMaUP4zqyV
Xlt18Hfw8F+p7wLbUk46PbX6xSTL0it7CTku+hUuobxpBI+vjWJ5LCbTri1/pEZ8
SuRvVtkPyRsSAUkouAGCBCK94vCikaRGfuJdGeuJoF5ODw3MSJo7KmkpgS79iKuJ
s4g6v/MdjiBiDnCFQCwDzNtZ+SKBMC2uzhuCBH2RaLWq0sLtIINB1gSRAOx3LhAs
yD7uWUdEY3rurzUvIBO37rbBcZ86qJW/e6F3hDtORlK+3GUzZsxxnOFJekfVuFYP
t6zBzxDDov+WuB3jXaRdoD19eXugY2zUPrxuRd9bfaF67Ep7Y5BJ60/yOxIeY4jV
0gGLoG1OamYLnXSN++mvsvIg/VLNiq1KUH7XFLfKODoFsO7uXjoKhx7xqqxeYK8q
4D6X1XCsnaladlNnbNSJAiHN29GFDmZYemngvHiZXraM1wb2H+w8OTUUX++LzSyo
gX74R97AjDAANWSk3OmjxG7I8s+s/McDV+ULAQ+T6CkqlAXrih6VOyhSBpYZfMmW
kN8cCTlw91LhKBowfYoNEqZXdZv/EfMxG/Wq1HXS1IFDrJgeqAGtNjwljkCZhQD/
Vt+z6NWXX6wCqQTy0tPsqPRjhcB9mTDklldHopnyO1yM1vlciv2pwcAFYnqdXb62
vpVw3ehiI083Xnh5T6/HOWE54FjWYmL3K6fJF59vOalS9CKw2znyppmm+BJpobbp
VGr688VcEtoOo89AJ9xavqZcMmJU0WxDIyQ7j9xZNG/tLlS9m25ExQKTf5EqZw7t
8F+hxezMIRUsahdQI0aD6TfJA0sGOGPkoieyXIB0VTJru/6sbiMTesxkUAp3WNr1
WvNCLD2CnGzsjcacDmbZRDuNNAsEUhopWmGONa7+rxK4K0/Ba1LQ21RH20FiUOEr
dnZpYJYDREMll0u0GId6FlgdGiRAw0j4Bpr30zukuN65peznfr0YTs1WD9XVGL5K
ivGuYZEyaNveNoZk8JQC8fUZyvzc9cOYzOrcEGmIGZy1ez4xe3MVZn0CBVs3WwYd
3noS4/iXjiKw4agcMoAm4Fr6SQ5FVc/BaXwbcVvkaRVlOfBWDoPw9NN7R1bspmBu
r7n9ZEHhMsj7sDOp21DZxgPMGWDtnyD/zWOXM1DKSCbsbG9ovzfXAVgTrlYb7SWK
oQlj4doapA1Z9HKdLlMFrh6RLPudmBIbn08noXbIjw8a96KxtveKkOsasNzlo6iB
/Md6wSljVPSfoCpviCT9lu9AmRy3jAfacQKq5TVihmXXtbaexbUxqmtcpfOScIMx
j6RbvPw8odgkoKSIOtq/dR+cZ2nL4N+ZtKHJdbs2B07OOobdBuWFj1gZ7KkEGDgp
nvQ5lfHsYkXRKqQB5thY6qmoih8AIsJXaxz05+xKDSucaG1xSZ78Ba6MbQubE/i2
T7g4huxMGODP3egsDV7XWc8pCurJue9xhLvZx/GDSZ4GTlYHCaeGn6r357D9GBDE
5DBLbMp8mzkQw5Y4XfEQ9uCJSHIAJqmAUNE5Hj67qrA4uuc8L1BCwfGunyRu/9D+
SQikxMlQbWXhjvZeOu3zWBiCPskE/vmnEKP3M8/WmakLkWdK8XX3IXWAzgse+vNj
L2jAc/3owD/iIAVkxYg67kQd+i4a6n6/n2j/q5VpdVn/20BRWMUZeCXEyzOcebTm
GOkQ4FiIdi5vWk5V3KwtOeUFCJupE3Z0RQX6B6+gyztwNk/uMsWsR3iOC77EEU7P
OFm/T16ozhUuE1ZH3kMrobJgZK6rck4WyRj1tXneildvgN3IS84GU3u99QXsBJI1
EBH8S+7VT43Y67YnARaovfqvu9V8kGLl7N4FrxSMXFTXAs63cKnGGRVXY8TjIB9m
F+zoO5DWMGLaESAjjC4YIYaIagPzDRLjNZa+24yj0+pFTQpAPzGtUwbhq9QyGt+8
uKGMC75R3z7+KfYUiw2Hk2qIplgPM8iAArbyMazKsg6wFeeoAlLSq5OJ9G92Nv04
Pd1FykFNfirz59BX9oriYUNdTWrXPo16Y53bLoJ/xiFwIGR1G0xDwwrO+zF6kus7
sScKg4+IPPTf0/QkZGL+1DLXjgSIS/2+CBcrUEWTI4UerCJ1b9bBDnX677GPeWHk
ePU3AS5nIcWyRltdvzd9up5XD98hCh9P/FUWSdLT70lqbRBp7BO05tM/qY2RnTEM
qieY/GBFwtRiMX6W2mkv+A==
`protect END_PROTECTED
