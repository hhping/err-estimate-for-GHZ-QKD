`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+YALcqRiNh65aabomU6ShesPDfNw/fHowuHWu3cA0w9Lmv+BGdijDi/ECTemzxL
E3hzCyrf1zxaZCxqaStmdPQjkzm7bfWBqk516NfVUdHBE7a2idnqYyCDa512zWME
rwmyBzN7pqy8SmGz7Ve/L5RZDRtNAVxyIbnh5NDsNAo5SafSSt9ptdX0AKSvY+DF
Q+wkfWd44d3BZnTFKVhMyNhuutQ0gUqZSrra6jqxcHJPzL3+s6/+wK+/u3lHAz66
/elN67xpe73WGnehd3meiznSd4ENXjrPKQdEzGyWEdfWAdV3eYz/2FFT9rFIW5vf
w15L7OEVESgEILAqI0TGTKYkFQh5ZSWp2Ko2j8CbMMEoNq6+MMvbigrTHyWVbmjB
085oablIF6uwLQYVH/VtMK0SAVNqTJ2SigEAGvuPxynm3s5+T7MBMDvN1bdvZ/Mr
zByzafIx5AwUQ+//3FinmimGCPkdZ0zlNSKjefYnpxs9WJjHUFqxIUrJtBcGCr8S
MWtJa/rnbCArIbRqEAMSUeTKz0pmqT0xcR4FNMsf37bXijiA9T7G+M3RmSHitqgR
ecIcWFWIoFe7p//1VdHly/0fS1xoJMvRxZNvv7bZPQ7rPPPyPQ6j2O7RXhJuleuT
58WVxTaM9a8gmqWG3uz/2aluHs7h25trZF5xBN5nkgxA6BlHC7uMpXJCs3uPdWMO
aAKprwa4Sh63aZkycZUosmmNGIYL8NFo7NKVpqmgiofExX2mHYkePIOUyBL587FC
YR16W/uBb7RcxhcLD4v40mLEeJex6vu1I005YhrUFHsgfcOlMXuHqJ1Z2nJTLGMX
wqQmkK/+x23nUqPAfGR7H/uOYjwEXrk37eUY0JbULoo3GGkYyDmBB8hKG/47HJWI
+5iIpPVeqiRuwpn1LbMXKPIZ30aZBdU8jqogjmXaHyCFnbq2KYshyHGT9YgU/T1L
xmBnmPufzDbqNOAbtXJAQJR8DO4rleMpXdH/SAsr59BBVIff9+vVHwtEM7bHr0k4
Qjt1vdwux54YbbrEz7xEJ7faEnrEM1eexBpA0KxWqUa/OdUrVIZOZ1F6GTcpEsx7
K85sZQptcJD/xkQe/jrBf57KJPWhA+qkMNvfo024NUwDrSxqCEOK8e0vsMavPWMD
E8bs/CoVVtuEnnMziM20MbQ9/p2tiIkNhn7LYpAqZtYNOlrFikqYHsHUT6ey4Z+N
yys7YxQ0X5HtIMZZlUtewcSj9hY7uVwfLt0gygVb/xpWVRd9RFEUJhCKDTfOGtYO
S8c1KX4Lk6m5nq6Gi8pexCbso2A4w67rGsI/3JZM/nAxLdp2j3ziBfhDqNK2GN94
gfFQjlN59pWB9bfxTzyYQ1Gy/rfm8w4tnPoJh2LJn6LzLARnY6FeHxnC6Ti1qWWL
IVi9sa+wQ3UqHo7qqdK+0xF4igHDNYm8MNhdAxejbQiTNlE1cqOXl9/C3xC7e3RK
Xs0EQ/kE/CL+QPjGvlOAi3QutKxlbZe98RXuyyaFOHwAWMYSvYKfKfQJAN0YIilL
Fcg0Hz5tZIWbJlSfc2aurkZWQx0nYyk5CIKFke/kjd573Up6G3TWiaj5Ito4784q
g+zypNggigX/Hv4IxkdOsQJU24Ah0Q7HSX3xtbNhV57bTiINcfx6o9Qh24c+d1wR
7vb3pXjFTlS84gqtbNx95kEVoZ/ucj3XdPjPN3oZPIpfu0ZU4XKmYYiuuBCxreWR
lgbGbJWckYa6l0a3whVODnBPLgQeHM3YkHOs9YGhlRz8QnTD6LRRoxTmD5blWGaB
dpNn+/2TqxojmHpLcODPXeux61f2/9K8J/cKZAsdyoMO8EjbWerb+kFS03KM6EtN
c2UfarRMb72mqDwvCCRVOgyLOc49BXNe0/noXbqXAwsI5cHHW0o7zuirIuXJ5dRC
eoPDSm/jjyXFssDKyM036NsxOS7dRi2pzzOM9+q8JNXYy8dM8RHangMzAtMaZhxs
SNyjBS0sEPJ4ArAFvkVGQQ+UzN0lIFAUq7OLYxqs581X3j+KXFafCEMjPct0JBYD
F2S5U/g3PECbAfBnc+0F+tKWzDUrYVNgh0PQ0yeXOrKfgTeWDW593T5zVmbxGuXB
V7pR0abUvrc2z5BTrAs3UKc4s7cmMrMKtoDPyeW4ERW9fAUMnKXze9RcBPrQp+48
KG945I3a/nuNwM4DaEDzvl80VddSYJYQNvRcmgYMhWRBFWtYzN4gTEGEte2Bgc3E
6oelglSaAoYAcU+oAKCdj7q4R11nl4RAAUAdPsRCyZLKCOW826/KPqz0AP8Q50tr
f2mY6PRx3oVi7oI19c8gs31hPi1jdaZCb/puVKErcTJpgk47EbSQucCdrexe2THa
hgD3QrICQpnqHWJKXA9cyf6IN+MplXhaFF7LQSHIBh11doQwPcm5P2/+yrj5AvgJ
YR9bvMV0VEu9uc5s7YWhhBTnE1/X6Y/de4k5KLOQBhWTfewCNb8GgVFGaNKVC3vH
7lQNnO8yJZ4XqN1GIhHEKpm8Z6Uw43Df4IwQM3cyA8tpfSKRSWGqSWDc2+FNwxof
du+63Hut+ROs6jJAM03Bc/4SvL0Z5UUmMUPN6ew1lgYXv/oWSXnNMlxHz7fMvVbO
5+8MNeGP1Fx7hFNx0xaipI+SrFDBTPbeRuj9Pu8pTFZ+XAFTUAAPbg/j5akp4tPb
nomOmye5+kDnacnv3Yk36RI+mqZ9VgB6CR6PvYP+Vep+uPRIWkbseKtEPHIQQRFv
mtJ6sUwrOt8n4iz0xBU8qIKccLIA/ZGH8TChmyzuHea/jCkZt7raWGyy71nYnClK
bSAAh7rAPSRR+zHyvnIq/UUZ+imXT29NjeR/DwEG/mHvugXLFaOWFjfMpBgZY5QU
CKusNsdi8JW3mUIaqU2uviTSb7TkU3VSIyzPc3XjM5dmj2ecM+t1Pso4kzSVssrJ
pvHQZnpqEvHlL7wsfyJB2Ctwn3douQTalzhlS2/k++yTYRifgRNVonquZIDfUNlT
nn58by4XmqkjmjRU4tYs8Hjcq8zcpUDUfcofCJg4al+dxi/Da3LWjdlMjUrFttse
sXF9j36T4AZ39oGKVScC3YakGS2kJjcwattQDoAl8/FisAD0URdukH8EevzXeYTb
8xmS51eR+Vze+Wau2Pe9vIX6wmVcNQWatNKNbAGOuJVlIjveQiYPbxgWkKVCAu98
b2+2yZ/3teWYIgAH5cC4WcynWYzuuzcf0hXhB80hJ7s=
`protect END_PROTECTED
