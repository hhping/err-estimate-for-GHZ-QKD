`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZvW0Sf8zDnuKmfEikal2CmFsveSDPdlf62Nlmys1y46DoVA9PDbhxEC/gjY0ki9a
/n4cZpWxdcOW87nhDTE3nQCP86SwK9lyVeTsALZHGDwumVqeOborR9IEq0tigkN0
1LYM/ng9NPfCSvWgkgBwpZJMlWn9GhIDlTDP6sIVPGCdMcSyE178B51iPYrjxHSt
VgiBq8Mp/2QUbQcG5h8PhlsohdCW95y8Sw26lT7OTYahgYeUDFpRQdZf3vYAetWQ
QL1dbzxg3rShY3fbpPrNimya7IM7FkNM4bjL4ktqPrDmsUwex4hVY9xPBhBc/Z8e
r9GIwQVPzAIPGb5s/lHwYvsQDUitJf1sizmMET+r9194eLT3nYX4Vdwa3xARicia
BJK5ZGI6IVj6H4iVsiJ75w==
`protect END_PROTECTED
