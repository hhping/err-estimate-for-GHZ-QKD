`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jud02VEk6bRm/GRUbjYhDmNtqQw7E+krDDUBTZTUMW+f9RYXmr/SHOru7MXKCmG
G2VartLLIUImN1A1HLgnm1iIcD/vMf66mk5bS++pDYB6q+qJy+KjW7k81jGpmY7+
RaElu4zt9npCEIfYwuLls84PWQT5chEL5koLNQJ8d2yrRTy4gDbsTd5NO0jwe597
FIH39D4sIDNU6+naQM7Y3G9HBeWD7k0DtoBpg8FnBYqc6mjkghcKZBzk0QD5/0//
wO8LVBBVvA7DbYWXwqiLWnuEP+bQ7XIJqfrwpylnhPBX4h0D52AesuR9VpSF46L5
DMhuxbGu5l0F4T49bVBjRn38vkrsSgeWXKOeGPNIrTHbIxSGt4prvFfp/rhKpSco
Qj45nNOvmN9k/ClePHxuIL2z4mpYQQdFo7qpBuYoB3pLM4x2ui0hHuo6Cfq5BtoR
uWUHBYoOUljcZAtNgWe/UQ+A3ezIcPYB45ksl1tDlQg=
`protect END_PROTECTED
