`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waISwdvGZ5k6nW5lusTZrwtkvSYpDYsr0P0VUX09z9HDdNZYH4ImG5gwpO9EeDA2
r5Y9BVKQHRUBbWV0Np2bRFufPyrBtwTH/WLzX1KCwxmuA7jXTzpAdftKj08miwTa
EgHAF0EvKzng6FACnEGdCZ01lLel8Yyhbd6axBU8iiVf6MNmwOGIA8if+bfT2yJ0
DuGBNqXfvVBR0XdTWFD/7A9jGV0D3RLwhBSyGG2Pmb4EBC4ptRQMhtjOeGJjROd0
YFqOSac0niQ+iZfJ9V5HviisNm2pXHHE9u+OtIrnpGVl7JlJ7mOFLqgfUpr3+ub+
e54rNlfS6fSgKD/QiBIUpd6DB4o2Bf05OKl7Qizx2VscCtqqQRLZDCyS5IOlfHDO
UHC4GVC9XuF/VMKZ5i6JblOI0fsmiyQ3bNBHKBa+05xQjUilvJ0m4nBo00t8VDQF
QKQfcT9zzKKvpRR1W5Zec7M1mSCAkW75KCwq8zpJEg2p9OxHmFssfZ0VMolnoO5W
kllMUnaNglY7QyDba24AO9PGoXTpZFRwdHFPnybsb5835bt3tlmoiaXkyTaQ7Bqn
L4OLxRDSFWqisQExrr6XLSO84tOoPo/fZNTTg+Mq7IL+AE25A2G9eiDx/hEm88TD
rfhWdOhn/Gkv0eDQJVF18BlRPeGoJpvRdzJcIefu1j2nUYuG1CNzwXigL8IOIhgb
h3mZwSHFh4OTYeVD3FGsVb9zK6+qLkSblFPCVMiiDZl1vJn84jmNBewc9J+IheYc
ScQPzHESMMqaHKN+t52vwqXZW3BwuzQEOYNBf9HvgNXbRDSY1pEQumuPIcjrVkcv
jSjNudK+VeB/pVe7fKrWFBHNi+tz8zWcR5JFupjpg6V8iPsDPVBjwzxazwdCFuYy
V1fFU9K1brXcWi+w/NO3fI+rRvAkj2F4qVblTwttxgqiAl5D/ozjUgSZrEtba6wP
ceikKQqfE0aoYvUpi2P3o/V7SbvbkakZKss4bUrgRjbMYWNIrls86bRJCKU1qzzd
67P7qtWrlZJH8BHz6iaDLVj/GDTO2kVCvxw4mrTVpOvQF/rT/EGZ3qOeAvVl0B3j
lbk7QYTtJ5SQks901MnjUBPjj2OEY/Zz6BomgWwdMaLVNDf67r4aPUwNXNXREjy3
AqLljMioBrc5TvxmS17U/lmuC+RIxzF3gzMRLx86WburZZQT/Wn+IQ5n9fKsT9uQ
0z92KUqZ5ron0DlCKViOWO8xJ2Ps+j2VEleFgcl+Q1nLw+6lX1fw9U506H9HQN7n
zHQx8EnfqclQ/y7AZ6819RzyxUI3hVt1mznNRuByLTOr/c53v9qFQuAMZ63ZkvED
v/Nxnl3BxlcGt4c2CSxl7bHJnoIBduCL5YvReLEvEAws1RFxXUQ9V3rIv7/U1kNz
iYm0bUxhWB8pDozvbIpjoKY/8XvUPO9aLd+iLimbo2XzS1oZuwjIQtbtYgBL8rPm
0uc8TnTTfaMC37hz+W0LjmRGZnYyFWGD6upEaSTXTrcb0MBG0eO7LgxUmvEvhEof
qoIkx83yQ+9LiEEz/D3zC2+gLxmh39ly8fIBy69kfEONa5r0DUDNRRMUXpevbMR8
Y/pws7kJIDM6rKAJZq5+QL44vYgbzOqpOogeZJtxqXivo8jqovM9uDRnyKb4HS2Q
CuHp0BS57DgpvVl0sLi6fz98YFs6Cb96pcAyp1h0tfcH1zU/WFu/5/t2u+kaWIou
Sa5x2QVofhBTbxpS82iwuioL5K1kjeRbBA2uqg/nhIWu1UrDczPi56E3G+w24gGn
EA7F4sCY6OS/YbiJzHXSTg==
`protect END_PROTECTED
