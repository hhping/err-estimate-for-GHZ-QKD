`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZiB2kA9QgBOv6S58vU+T47+9jPPnJ9sQLiAOsFWm6Z6iwIslBQ47gHsbj6iDmLa
lfMD92k5odqLtgkgcArjbCqRXuNblBNsZsD41Wguo/1pfAvB8JX7gz/+jB/W766e
jiUXfYMurer3ajXFhnQ+faCBIfxdByvhuecsXaRvMJvfZDAavjgMNqy89e1HXBEC
Fm66onC7cDiV3W8csR11B9xtB/AoBGa6+pX3cCXCVeVq+4Z6K04/SuaBXBc1jLTJ
9YrbQdAOYbM0Eh5cJ8dnj1ksNl8/sawkkElmpifAy5m6VflhjtQmvhJw/4qQH8sv
MRKiEDLGPGQyxSyFKRQgxVNlsLx1eCt2zKHeb2DBVuEsiUQxTagCMutmGRJ+zKp7
ztOherTaTZmoBgLtFGoi+ZgPVVRdI+/2N74WaD3seKm5tGnv5QH0Xx8Q3tzE763z
Uj+2gMlCI8zQZu2j1ipm1zOz9u1tFpyaVQjWOr6UxCSgkY+Wi9jZunTDRPrTeAVn
R5KMeJQMAn31207ay7wvRgWjumxW2bajWH4qKIqXgIJNdMUDqoWoRLdT0TLZKnDa
u5uITafjOLNltnYBxeB7Y1zXrx99Kdjmp1IzPcSPJcfYyv602UVJuxQjpgMhY9HD
z+355T7d+MpJwFqI4pndvN4IpsZSG71wKrN+QgcLv6C/Udeu9BwxJJF6QQZZ9nU7
oq5oUa9rEPKZdxlHKUo2Szalib/jKn8gnaUOiXHfot2P6SE18A9tJcHl0QQKesQr
1U6a1wuL7rXFkOVzUVo9sGFRB+lVcQBbykfvDbbQJd2oPtc95Ou6gms+ken6Gj5e
6l4r18XferS2IgiXi3+iKxa4dZ2u78lXPHMbL9DlfVEW9TAsMKPbsKQMPcwCOVjO
p219pAg0+5pvVOVlu3DIoVSigN6uGfUludc0Ns+OKuDwfUhyXy0cXhC1HwYhtqDn
XHogQOF2N0l2TNIxj1O12fIkOLmYl70iLlHjexykV4gJgqUGGZ7RLIdYQAidWVwt
69Nx6ClpNcBiip7j45Rn0eLJEdxcCTnTh6tdgC9BUEsIxl6l1ye0hFve4wkdxzzK
`protect END_PROTECTED
