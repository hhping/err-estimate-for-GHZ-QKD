`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XBdBd1apWYJY+13PUWUqpKMfsPHxtNe9f/QPggsF3f3b9G1i74g/dqxXRAy09ik
hrSpga9pvY8hASpndy1VeCe+vlZKIEqM7metuo8c/o0GCZUQwkeVyH4tybYTpbbX
S/zrETinDRycasbWRJZ8LcPofzNQLDPFcVh8ti1KdFzH6lc8LA9gi2x2m0yoqV9Q
FaF+uvuFoV2JD+yvoUQ8ESWww8/ElAqXQXihUJKQrgTC46qgIybrwVtOEMHfalUe
lOfw8zYA7E3zCyyvP+Y8sQetuKtjNQyXK0ZV30Mscr28CflKldU87y5jMrP79Dj4
SiZcvlhF+w8rQoC1aHO02YikQjQe/wdxf1n0v57uNDT2pm7aps9sCBt+REPrqGVL
uZM6e6sMRoqUCYJV5sg6kyPILEdKiJIN8+TJasjrW66GmgHICw6Fl9ZcbuBKK8ze
cxOffKLZnlyG0IYMGShXspGkaYEHN+NNf5p3wOiMw6L0e3n2DDyDLnGllC7d82y1
wBNfQmpxYurW0TTt924BiTvubU3+VrvDYoEd79PJxwO4usE8zWCmIJUIzDaitZaG
/xSztPkyU9BUeqPJj2+04uaY5JkNJ0U7q4URA7dnQ1c5ogONsjlBRLxR/GQ3Jjbr
FJoQaJ885bPYjvi1dls04MBkeEBurPmlU4hTkYMl9OlQ0yl+1P1FyYvh6Fx4UxgE
VB2g9mHZmNHwedgPiYJVFfpoS5fgZMKS7wrOgpMpjiscyMflje7qLc7VLDZpBNpk
w0HfKYEiH+vZItNCV1XERevrNpBb6pWFFZ7t1emf7oiQ2vApljrRdZGKhXQje/Hc
L6GDH761hSbWKgcVf2+CGBKd4tnQR3cbecKzMbeu++57jloDn2vBztslH+TgOFK6
DZ24RKiKtYPjoF4ZxNRcTollJq8JH7xnQGpAi+KEFLpzsRswaqQDW4ZmhKTGSvw6
CY2ys4UQ1iAoM+OFrvvvmEzG+GFTYOy3W2T9O2tk+f66DldZkmAvoC2se+5o4G4o
`protect END_PROTECTED
