`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmBN8ZISqW3QVZouoBF5jEBIT8YlF7QhSB+F2dkXTcUKfdrLSTSQkF8xGP2OLAkO
s6Yyeb1dEwVlcQzLmlkGFAzTpukoHaVbFMYvKbqh3wB9JquUXu5nk7dP9Y5sS3HV
ylni5y5DfeFLXcn3HdpOfk7ZVuG11QyhBdIpvTDMvqiSPhFFxchmgCkxUkANQe+Z
U9vmtjTP4oiG6SjNWc4FZMM8fNzCCcrNFAAFexMY2MdZNdZumOuTAP+aLrshHqjZ
N2OFb0CTtp5oy78teRKe5Io1fGH+nC0VtQwLfCGfYP0zjhKRjVXbEUcB3e6dOoEa
eVIygNt/RoruFpIn2UgHkCU95jnw8zGPmKrW/jkUl5wuiPkC+IotudHx/e2vMy29
nXoKbLq4rCLkn0UzFc5Im3n0q1Uwi4+QTqmpEj2bBjfQVYzOXC7952VZiNtoxZuR
9gSmVH6bhRhqjqY9eDVt/RIZrff4gd3PvQHxN4IG+oahiC1Bceukf7f4xUiiVnjk
Dni27byHKDsTHdgJ3YnmeT4sC9QGJMwGfrQ6kP1G67Kk0vj+4cZwlZ+Pft2/WDFX
gVVhIgkEzq9WchDH3ojSpjAYRESWzOF2MnHEfG48HPyFQYrMZHPNVoEaFz8/4SWt
`protect END_PROTECTED
