`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G0iklx0LHKGUXk3WVAINX22NKkMdnPUvwZfPwMqGxeULCYJfzHomap1TsOPrl93B
o6jMOiLhxBfVKW75/BKpqSBSteDjGOg2byWsLcztfcbjBgU1iEks1HgqIVP6P6zN
pgWhjJeZDCxoB9XaghZu/fPX796dDkIUpdWEOKjmn7vq0xbJrmAeM9u2LBkmVtm8
6OGeZbsFDIU05lV8U8etEwTrLCZ23hwxNnXBIV5MkusFgbrodlLCu9m8/kaw78VG
AeL8D11Co1v3otImk0fKZq6e9lV9/NQQfWGa3t9bi24os3t/NJiRH6U/Oxk4rjhJ
gXR55gaID4swXCc9T3Z7oTsEiN56+oX2ApijPdTYtv0hYGfstYCbiAnlvl5qOezP
tZ2a4DQn74rhqbNGXMTdajmonbIuSEBnKS0uu8J7zYXpc5+cI1HUW0qm2PMpzHUk
yivE1Gg+GZFXqMZn+eb89rI0jxYstwxykPM2ZfeUi66jr3TYvJdYN7a++2DN08cy
baiHUVsTk+a96b/eGiWgx9ER94WzKsdhSO0h6A3wOLwwrI0rcMuobxV29GbsT7IF
7MXzpauV8hf+wLSoW+z03gz0DkoVFvCJQNsI+3bgx2Hquc4U1ayVAILWH1d8V5gu
22XOM2bdOWJZjJ4qvnarhmqYQPaLET9AxeldjEswCXGcTPIbySF5pTHI0bg/b+Mp
NJhBZnkZG5KYCmDZhPxHMj5/ap7r/6ysR1OSLOi/c+lnypjhyp5p2lRmqEZ/ZKrJ
sZLW7uP5MFDQossMJ+A4HHJbx/AVsKwJia0f8IlptUcfd5RipyHUXLw4dLj+hfgw
`protect END_PROTECTED
