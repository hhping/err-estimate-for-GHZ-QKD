`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Au46tkk7mi6bKIPJ5lHmYqHpKOfyjvOVBNoD5GHAA/Z1m2skrm0YzGIraJpNjFdg
oqFwYmH37tJvmR3ihNILcwfw2DoN4NgqAm/GWAGVzu2xYD+a2JC5OYv858U2R7jI
nUBfjUAxJVqAG4wgv7SEBI2mt+znekuBTehNT6cE7SOOqE9bixxpHt5aGn+P3hxU
oP1VNbQh6V3ToGgJF5n+KBotBgRmt4WZEXCAlWRBm8BjfKkxdDZ15fQrb3RCPdfm
YjBly4O+dYhbBHHvtSiLnvK/IdR8WV4hC1Tu1npiqPsq1heZ7A4RhcF5ou48X1Cy
tH799HxjvH3ffnw6fV3bPG0/K9zB/xXblJrOYvdnF+GzmOQEGSGZqEKQx+7HGa2w
90S0AuccMG3WqNBGiKFNRHsoGcGtnDTWiRsyTVIkFsZJ4EC4os72xj3LyxLZwYlL
+IbME3vANUi2zRDFRwRsRlDg5jf5WL1SyfkbONOSWuibvwPhxsh15czt4avLD6Je
dF68etv9/rMAu3fj+zmwOKyvTgNOvElrGDLOjLByLZbz307wtH0sOjRxv+vbC+hm
PYftnW0VV7djKDlrMdZTgZ2rywIpaFLOXLxIaiTVoJOB0gVgKTJ1cQghPiN1AP40
8GlHSubPiBqUVBbekkoycCfIzmy5gJpdupYR1gWxOoi3ZcQqoU91V/S+vynEuCne
w97HjarfaM3LJoEjWk7y3u1tWDd0/g7hBqjqk4zMY2ZXdTFOfU7DwwIDSJFHYHU+
bOgqttrAJUbE74f9p9oPCKlTk0ntqLZDBgEIAroLzYOfthdmgh3beYDqzm8mVJzX
+PoRFhSUWg3YvHRK3DJcNKelqPyn+e+SDHAkADB4IM0ty+Oq7Y9a/XpwIRwIb52x
evKFp8j8YB0Eqo4NFsOut/XsfL+nh8RpQDuajdzH0CP8rrlzQScYPsPtLvSSoPVe
yFO0Z5jUodBCvzNlZSIy1O3Dx49JysLh3rCKmIsdMfCWFJ2gy0El0r4KpzJD6hbp
FhnDfzeXHxklJOJPX+tGvXhBEE4llUJgsmE5f6LDqok=
`protect END_PROTECTED
