`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pvS6twafSY96Izj6xjxRkvp6ndTugvSBI1s+G7ZxUQMxekmfRjcA4fsirxY5Tnj
01jSQU8m6hpcqIJ71k26q5lFqFVw8CAS8ltzb0Tb9IJzdE3w++UKVQcG3msj5ZU/
BF9cR6DKONXmbT2pP5t07atTqkw8YaHW3DXGG20K6Z+3WqWu+nwStx6dGhOwjD6r
WGAzLS7LH+rzybgJ3gwJAdBOtgWEOZEarpDB5uyGSDEqbLpVhp9rdsaPfKexBCpM
zys4y/nxnJ2QyRUSR0xFW9g2TWXQ8W5WU4iPN4ychHuXe+chxScnsmTyhP45XG3b
66iGCoEGFj/022LdKf78799ED+gNnmnVEDWrqnL0yKrq8tce4TVurqMwWq0nxTUQ
mEE56UusFf8eWp6qn8jeZjbX49osnlUH6V2v+7tUBYR2X1Qfr9CUDqQrpVnBvZ1L
u0zAJTqBiFEbx5tBMWQgqSyuV579u31v9Q1hRtZHgtqSFU3K+FmMgwHvMYKqLe94
kcUZV0S5jT6J1HOnyFsOUg==
`protect END_PROTECTED
