`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EgrtQ5dERKH8ALXEl2J+yWIRXJD1zf8fcnfeSrM9fC8M6V6IAcM8M13nH7cC6YMr
bpQWqlHL/Hd94wCKUc+TxhyvqAvI1Q1Ig/s6qfGgmezCGZkQpjq6b3d265JooDWw
FtMIhB0MpStWGlel1D1BMtojBLH6ImxIu43kzJEbEZ2cnF092GhKpBymTudJQBwR
USXE4B6ZVkuc9RKz7YyZX9EjcFC8PT9LvmyijIe+lGPoZ+xmg+SuMYm2wK3ldtHT
CSq6GR05kvZ/0e+rym/PJsY5HRsZ9uk915evUjx9XpSzb7akT8l4KxJhNKCNMiDx
GOvoNCTofHbEFyup23wlvxPjM8RlpDRP8JXh+dG4JYl43a+pDRGgKZ+ccdaZtX4E
YBRU0HrM0cMunPfBEi5c3C9QyyRBps5YvG/5EWxH5WpI7p6co/mYJV49L+k7F1Yd
dPOK59xXMQoz1FXm4XzwA9V4Y/j9h5IAU4AHV9N47NHRb9po11o48zgexBI0Ccj6
o1lcuNv5Wkh5FyXFMxp3d0xu9u0mw3LUkrOznWlZ8TF2+jtyCrcZkjMpqr1qV1rX
2tnb/iSBNNn8ZGC+6Pr1UgCWvik6H2npaCa593zbF1QzLJuavMh0quWj99WxdMJT
0cbqbWoXyGPjePETW1RRRcV86+tP7mzbPyAMTxrjb79lKunOnHf0jgkVKJRffpyk
3mBCxsfAg4O4N5TLd/z551Rqxviy9ta1Yh1vZNCgh1MrRLEdpbDvSWsIXpM7ponQ
+Pg+zAITsaPyEyrtJP/Z5RM13HpSZ+WZbRUPl2gUdjbZ6bh5JAwWlMKEXu1XHeF0
OrGh5qeDwgQbkYeQMXm55q6cPIPyiYB5AqGcSngUD0x7NhlTbAa6ooqLCu6kkgRx
NKhZ19fRCgN5+s1b5ycjfta8/qc4/hXmn8shkLD9osVs08WObgW7wX+21i5hZ3Yy
MG4vyp+/kyZzs6huQmlB42bxuK8WOueyw/dx50C3BKQ5sq13zH6g6CpWwEg6EfzH
6SdcnZvKUUrj8XFTAXYtxeq/cZr3xZqKvafgGD/p5CQH9VF5r9KLG++J98qLHbuN
urNitMkGAPGRNeje5XT43XEuJ/pLe8hl+7V01ujZLa3NQHtXHbtcb209/Ev7J+xH
zJp6nGVqcH4tPvkrc4k43RmWnYQ3Is9sysjFC+LDFGyHpxOnfVsy40rmaoKwWC1H
tS321+P6nQAbro2Lf+8OF/4nm8s4DsQeWHQAPBLyTVxsmyi0XAFLnxJQqYUyry27
+qSXfzJFQArE6yy5YakP3TNGaufbB8QxNnCrBetrmg+Rl4C81n7DlBcS2/ZIZinl
`protect END_PROTECTED
