`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/pNJChcLC7sIblJYKNtU0UiCHYX81Taa1SpgbGclfORfSNhUMoI87cn70Ep3gb+
rnAaOeiQmX6LhwE7urIr52atDtNFw3lz+N2EgEQlWiOJ+1kgwIKuhGoKRELQPrKA
7mCIBmSAg55KuU5CkblWrsIMJEufTPfpjBxVM66JZ/wlZf47KR9wWfk5wze2rYOs
I9N4PpPS0Bd9vO3JN4ZsjVqgV7Or8hLuJgbkdzgajCWZVEdbAvgl5PC+Lmhnpmcn
Vc0E83dK/AkETAiZ/3r3+Wn+VvTeZ+STk2XYwMWwRkX6U0/1+nuElLH74frqROvW
art978XRZ/JcSUkvPJMsLQVAsH+BjvzYSpOZ+aQl33luKwcegZUYJn4t7s60QuyV
bN8RPuXMWoRJMucJPJl9aqsh9PVtDzZ3jiJHu3F0l7B1Q7CLCnuVcTQdefY2AfQS
jpuwFuvmTkUv3I8abTxyHESmxcC2rh5rvlY9vZi0jCwlVbhgu9lMGWfkpSvV8sHv
Q/R2fIHtERkmsFLrFw0HP2y7UVxmxesl2NIcmwWFkPkrRtcvUS7DDJxfG1yE8oYr
vox5eqIEWX7nZL9S5Fs4tg12HKqgStzOg6hzTXa5RIrr+/7xzR1QU75SMjF+smra
oyGi8U8E8fHuz+tgpuAmGYahjjFLboTj87Z+zkQUiqy5l0oH7yk2bTIBKdev/7Xe
eD/Hobtx27k8gOLQDMqpVsqfc8sXw+YnFGbKqEyVD2AC6OLElXtu2HNqq5GOTjjO
h8gLTM4cs4qvC6ufq63s9ed7vdmAxsm6kkigvqyI+RnrPVRYGsFWFlQr0JmuzZuO
24UU0o/7bUjInT9ilqqs0uG5aRHniCxmszpWhqUdgjwRscWlgZQyeOLWmxxPSLLJ
NS8vlyswfaXLelHisSbTo1vNVoSAnzmi5tX3v2YD9/zJ586h+KHFvfpwmWYiXq2G
XEtlGgNoKA9EqFW6v4D7Og==
`protect END_PROTECTED
