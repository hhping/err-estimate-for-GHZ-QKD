`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEbRHN9cXHy8qB0YMPqgl4JpTXYfwlzTX93tG/8IbrG1THX95LQVNb0lSyY5RVWq
XPqfaYYHWwDa7Ep7ApCTu0RXLILE1ZzeiMqekAsuVIAdp0y8hXcyyNnbp9cToZI2
b+Zp5uNlrBWe1soprNYP4R3DPEp5q4Sb1xOZGn/zHQwK8kVm0QwyTJ1xBH4OCeCp
zMf9dh1OwcI77wT0WIFEyjcsgpYMU/PMUoFG+EPG+pNFxTZGT2tTFEhTAbG+F5R9
zhD7VCLvG2Lq9mmZLy8YXtJA2brV6HGlNOMuU/W4G6+B6ZBalZj2iRjIwNoxJnzk
M+Iou/EoK5H76Uk6nW+BdKZ1AMp5NzJAg9Ha4N/OAOxbgJsAs5OhX6KLT8gMfUaF
Awh2oGFeaG+sg0pwkzy4sQIlSAiiyIirW6G1y1BB831uU17eDhcIJAXXW69rPqS+
70uEUIur7LmG7iytYDwf7HI/j9A7BR+eFX0ZzWxRGfo6IqWDy29h41WpOeKTBsAG
deX0qPiPeE5J+8bLszGVd3XpOtPBdXDOIE/vwS0HZ3AdC6Z0i5597fvvqjzg24fJ
zwtsYcq4b0L1y05rCUMJHyEDOey+RAaGnCWFLP5SRVxRk5LOFm/hDOCjopENMSeU
8nNeOP2PiqNla9FIRpmD8OlsJia3gOuQK07WFUfMm3A=
`protect END_PROTECTED
