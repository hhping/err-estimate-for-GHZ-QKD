`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMxWHt74jX9uXR+2tQhid9LDxTQyimecD7VQn5R0dKqVyjaVXebc+F7Dg9FtfByS
RvydR6SF5TqoKNEdECECRcI1cDWh/tzKUe82DEHjUJ9ttIbzqoGQfTZHzwmcwbrK
uTg8CvJiUl+PdK3PQ6lEnFuKuX3gWi7+oZrGNN7iRXt7joe9h+J8h8aS199JhXmG
9AZxKWtnKIhhqmcRb099CPjpUZWwOYidj3AC4+xfr+NQulJlWk8Dim26j6jbB7We
qX7lFMkVHf1eCwamFM9bIGvX7wx3jC+yEtRrD9LH54cVvkqZtS5LBjfgLTY38QLw
E+AyPNeouf167soJpdcL5RkV1Jx34emggG69awUv7NuBCAmFzpBVBP+h99EwIOR4
rnBr8npjYpKRrlAe9jsSte23OxIM+pDDQwdbkIv6eDgL5xaA+yw1WimI/8DVxUt0
ZsboEjrtym5ADi+HtmsVcPCWWd+LZlF8vyvxYy0Y+Ag/gDn4emh3Fft1p6XjhC88
7WU8zGA5yjjbfVv8uWUf9bvlkoOAtpHAZ3lHHHRr8sHTJMohQKqiu0T+ab0l5UsO
4nte6W/Bmn/8JydJ0phGyEOhHNfomDS3JF+DZzEKSkpEsYVPxAnmaorV9Fl8DAiy
7bf4nmZW76n1ZywTB4l23rPTpvIYy1o8/a1tDrA681CaErr7NC8RxzEF10iEKa+r
ac+LUBYI5d+pbT+hkbUrclKILxY2XTYhTBBNVkOC1CkM9ilK9KoelvXUXjJAAAe/
ggImaijMndjLfdJPtWyV12FmK0YGf2ya6xL3+FhMDYOZqksgHqSPMVplecICPbem
ErA7i8VG1Z/QGik0GruJhY9m8Fcrcge3UuMyePVcP7mwNskoPq4lAioZPqCKGtp7
lRC/vXGg3V+1+DdhVXGIwfD/vDoXXtn2W8vEVV1PQUodlQ+pEC+g7Dm6v+/O7AJr
822RbBONPx+RGCZF/8YbgM9rjjyphLppr13p2PT6+8Wcpvdi6fLhlbLMxLuuSViA
AC2RACRT7t9FUgYEkHiqWWhaVfhMIZMaXjw2Y7ord82Z9cefE8yHPNjjGPcwCWU1
WuudepcHrhANk1B/lKZ9o8SstF+PRMdoiFGQ5kBSlnQE635wM03ylJ3qwovZo1o0
+IjEUF7lQSI1a8GIrkAKZUBAiM1jLm2Pwp3xdqUEN7FE2O5OAb29cHRtyrSyAeVQ
+tiLAgmLRdVMHBWdEvx+peO+B0ZEmfwzpIlnZO7M8PXkMBoSyp5nl9vYylvYr8vI
0XKb9cT/E/NCjlsscN4iKHcoe05KUV8ePJCcDR5SLaqYA0Zd6B5p5ZAOJvtBVNfe
7HTo+Kdh2bswAdX0opVMt0vfqcsyXx6NlbuZKJiN5e3RUEkL09339MKqFFY6ViPC
E9pdvCpL7+gejNEAOumt8F5SaA9A2I4CmGRnF41Sbe1UEUHY1/pGVL072ThtxSHJ
9TJCN8BKXXvYfAKeVpl35R0ME2vGWixqcCypl8rbP1ORqzZVSLtn06O1+0WPWu1W
`protect END_PROTECTED
