`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+2bHE3aYAFnjgdn1bcOlTF1bLZ2CwKRC6I5jtGnUucyvxYvdUo408wtfrFy4rrZ
qcsK14wR6XRVdAVdk/F7fOjuyfXs40J17ne+AmUaDxFXxmaX6UIKH+ntA/C1DH9W
XYIsz/Jc0JD/Bv+/OrwCVfLzldbaKsLolLx9MTa6Vm26Rs3Ezqj51ZqJM5ilqpAU
RY5ksjjNPp7vxHZanUFm1AHH7z+1hvurN7pEPLbyCWWSYjh1RIPPCcoK+BdKqqVf
TIPPmTzmtDQHeOoPIYOES4fRaTXmYydIZWYVyc6LTMzyG8boiZwLdNEJnq3HncLR
iD8fdXv+Mh5uadYrqKd/O/E2BrL2nU4tjXJZnkYYqz/MIl7jHWML7sJPZ8V3rVkA
Gj6yvFIhC1a0lEUfuRtmoPAxwAOTqh/bOWKZR2TWOtoJuDKuVLwROzA8gOMS+OCT
EtaJ3N5fxN2oFAOsq22es+b5ZwehhQryDAHsoEhMkWhy6tiJaQYPGrj85gtmMmw3
d9Y2lv9pn2Q09SLKL7lSMgu52IGAWJMmNaj+6XdGni0Z61h69ErQg/onBWObJz1s
jiPtbosoMLY4cDR+9iniX9mG4CZNqKcvQh+FM3l+9eHtC32qRI5yoy0nDGKKHkAy
1UzD3x+CjJttMk4cflhkZ8RMqbWCU0NqIIIie+FkB7XlmuhpEQ+RDnHQIQwgNxQr
48Mkt9sb0wey9Pdc0QpE/G9J7fbId7OzUtnY6Su97DatisV9+L5rlOWNkZPEurdh
O1KAACOh317yRLp/X5iuDeZ2fCYEoe3Sh2CbRh+qyhqNeRp4eXAMI1xwYJCuBYRv
jcq4TT151F2oqffeiHqmihDNB4r3WlOhAWUq1maJngRqAx50p7Z5WJPyf/GkGCKg
9TZ51OazCtj47yrzdaLPU6xJJxHEN+Mgr+qaLd55n2RqtAiWE3AXcOm4+iSudWdx
9Bgpg8y4etsYYYmnnFyM0zezg1KSinZaYbo33WJWr010EcCckVdzI+mOT1BZbR2a
3Dw5e5bMiNhdKUssXUXDdWwTfv7mK9LRcyTgFLCsBh5LFWY9+nPZMcca9fQvAAVS
4lyKlaE2Wz2H13tAtqEs3j5Wiqol6PkmpfzDtvzMrOPNn1GDvZydQyPKM2in9Hxo
8hVCcgdO/h3FV/Grqf2ZV7VeYrZXdtFdh5BZUZEG2D+U/g/wFIZckNcsaZYXRl/o
vWh5N4za1uVoCmrQaZMzitQ4zOIyfjJfnblYbuoizSY9vlXyGsqxB+Dqu0q76OIS
iazFVz7dwkg3b7qZOaKbwhMsc+V+dYCk72EgeWnvbDoPzRIqFr8tT0CzDa0WZCT0
GXWK+pt5dumIckwC+SKUVKpsrlQJyyC5+n3ABee+GOF/mK8quExvmOVvLjtmpjwx
+xaIfbfwX882BX/CcI7tftmdidRCwZXjM/t2GKx2Fnx5BE+Xo8oQtNcKAozGFMDC
hTlqDYFCi77e1gX4l5TyIgfDYQvRp0gSCqeSAwuqt3vIsT3d4+fILlcFI5Y/dOr+
vPi+PUVkEEX9eOkASJ8Ex97wsSAkPHYLahAw8V8AqoUz2Q76JiUP5BZdZ3auX+P9
yFTX7hKlSUwvB+7SZMF8pZrZfqdnWMPM53bptxstRH9txPJZkwJ9CyaH1Zcs28Cd
/NbjAoVuQnu0UOa1pw8BFdtWMwzSN7+XjZY89xr5h1+hzX3XyjzNArnW2p7ceSKs
XobHo5pR3RutsLpCgLeq4+5o7KtGoVuGN7niUualeHG7PZGFBds0NtYOaN6i0ws0
JdxvUAljxcCg+TAyBmloIM1PXRNWT0VK02yQPKPfG/0lcqJwQbdB4Ux0/8L31xww
ZBknPUU1pemmvOmORbcfbWzY2+JdAlW32ZNbMWMHLgYfOuvGPg+xv7KmMhz95agP
Vj6wcgYkIzD322+uZZ8PMNQL929MkUQ56p9+S5yIftFQDRDreacB+VZQUwI3PT1l
tdHYR7Yqa8l17dFFEyrcJSOwGhBp/3NT2A4cSuL2Mb/X1ZGmxiGwEIJGEjBebn2f
6bq2lcRuw3yAA/awOY/708TQVReU2qAhSqhr4fsBZOhK45RIl9h7zJqZCpvS2/6q
Ea01lUJcVqqj7eQBoeTk4JQadfmT8yuInfx0acTxfJMRnF41zqS9y6VaQuKZyriP
GZafkrbABNxA7kN8nZGRPbFSfJn+XJNY2RS7AJPvT+VDnetvFhkixyXCH90uhaDh
oq274ECG1Y0spoU5tROB+T5lVk4jWdtI53KT0XfoMgwDrKzL3qIlb5U6QGkIrYc5
F9f2g1c7Q7DREyP9m4Eakze+A0qT0WnbDWAHZ26BdsGiY//yOIwXME4E2XoIigO5
iuZp2xmh3TkiZqR3bM9ra8Zd4GEHGLwjJSbAaXF+j62CLfI65IzvcAQf8M0DLU16
+Wt5eswbB4K+aIoI1tZBxGXF9Euc8ipN85D2/H1cmZcTgtwOoJEDSQ48J/ApcqNt
isA6ZHmCfUoznUehxzZ0Twm3wHS+kli99l6Zlzz39ppRqtXIanFSE4eppIrfUQ04
8Nr5J+NXMXZNowARY5RFiwKgC0nbnWQFpiLRW8tdpEm+nwQtT2dM3vgJV8nqGLI7
YllXqG678m5OsmY84VPHQnETq+7oczxFicsp2aRiqLvX5HaJq00cIRKMb1cMZq2e
fVkRCQwjAnQCjoPTXDuqgV/mqvOK5hTlND2wdlRWRNZLJ4wQQdyOxfXd8o2uNkHI
07qdBgOfvvlZvo8tOy27vzslBR7LP3QbcO5A8qGl0UxVQ5oXAnHTsVYgPXxSLV1H
3cgL0Ir+jsHWXOgyCrml4mtUg7R5GafgBPAaUMAdRChBxDouhX2SFPU8wtfe5Ovi
XDz7CHS6W4tSLpbWRvBkB43yqI94RMv/n2N91H7b7euYeKhRNzGdx3W2+CWh46CU
6PDznG8T2TJye9Pnf0dOF5Kk7blddX39uNbDE3dhYETGdocIv8kDzUsB080DB47R
hgaTBUcvZgl1tPTri2qoS0xb6pQzmIpaDsh8eEeZwA12v4mKN3sfBBUhSgya4aoC
hPxBHnvaLDCswmJKFzNkdg/d0W6a7OtJ5nqaqykK1KszonFHW6U9mMWjAHWcxRR1
t8wjr4IxHD1+s8WP5Tv4LZ9Ja3brCOH7Q7CtvXMj0ucqCd5iRSC5j4NQy2yLvz3Q
qNnYn32dChQ/FCoGo8xBRUfDWNn6kFo9OsWFkCHDW/V2AzMl23grdyebhwpHJ7ua
ya0gvk9I7UsZXoIbLBPzUKakqznr2l73+5ZF53Wo2DUQY0aC7eKf/JECaJRVgcZB
bIM48f8mXH5zyoOqmw5rMiNrsCAfVVFGtoA24uLpC+k5cAxiSrE7MkZw2VR4+/vl
r6ClNi+p+2414f952EAKnQ==
`protect END_PROTECTED
