`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKJ5myk+y2AO7Tlkn2zdVqVi0ahmMQMQEKn+n+m8uv5/yp94iTnwFXY9KSEmeqbY
Xrs68Epx+CEyVA8nANf7MCjBwXrn5rPJj8mZWkKbhzysHMLLTmztEKKdPzWMseD/
S0Wuasa0IsdERjgjChdJIdKNB21aQVen1A/pzt9brmp523sbx8PjsefqGRo+5oeD
cuoe/jVf9fsLtmjIprsbZ2xum+OBhtC33HRtysZm1jiylMz3KAg9J8UODxK7ZAZS
QtxQFxNejFDJIfjlbxlCAq5NSqHTO93ERQU0z+X7Jx2XNe6X0dZqqXCKlbTZ9Llr
wOyf9PlrG8c6LTAYzAwfOlzIw9OSeNAeNzSd8GbUI7m2au54ZSeb2gNQVV/3hBAr
iMAX6wcsUIHwy6jwE7tMkeNFltsAdLNI9dVNyLICAjd8+nphJU/kRBGOTwSfHlGm
b+N0kUK+z5y0+hM4FqrWGRuKIJy0AvTRPMhJWmPc9tMhBofv/OMWtx/h2bbyU7Az
Bzo6s4QN5lrD25IZmL+kvKG5fSB9vBDoM489kvBTlD7eD2R4wT4EURlRf9llyWDc
Hw7cdAlhH2RLduaBvBiPr5V91PytWdTXk/1F+e88YsL4gAOiN+qS300EBYaxlR9+
xz1EQfMBd6VgWp5seVWslhnRN/KaLzNl3TmkOO+TEw3+xj4ggWs7HC/cnypFj4s1
POKs3EQ8S03NPbszRollJgj30Abr03gscDIrwHFgeh1ABnqZcPcZMBRcSpBwWxH6
ewzPN9PS0RHmT0fsq2ujHVwx3VyD3y1GMgNd5un4kIez6b9b1854E+6cXnkVtz3D
SZWhmMiHxssClZO4DWb7PTwwOj6r2mB2pHpLrW21kJAGdEQW0UVSTZMDFyZGu1E0
+b62VdpIyECDtYsV/j8BfQmYIb+NxTBQNr1au3Olz2FCtOdNCTLeYRRoNvWC+RpN
FZxYw5C0J2YYOlElnwy8Ozc8oz3cPEzXf5DHyMjl51lJ6T/Cm3BHa76Oaislf3d5
kQl/dMEpPD9WQtYCo+c067bEC1N4KhIuI3WUAGp612rDpPTZcYKq4EYNKsdd8XC6
YtsROJEUQqZ5IoxPQlmq63KpbfoSXRMz8PYJRT8/KGemH/V/sN+A/+Uzu9Ku9sTn
1z4LJNpatUKLsJeIh0DgtHM6/v25DbE9BdpjSW8rfbtr16b/mn5hrXyo11XqSjqd
upbiJtGvHZtQJ+2vVnz9qEQYokAMA/cdkclf3eDK9o20JdZbB61vC+eqX+t6dsZh
a1pu2csOAvR8vVGMW9eOS40AzYUUrRA1Eqppr0IMFJ79xI/nZUzvFMUyY5n4ZgcU
z7min3Bukv3Tml6R9V7q0+b6jr9MfW7PWpB1N3kOXEWH6+orGvKxFJPMvk4YWc6d
L+QvacDzIOG9yjj2GhlI/ryOg0GIF8pcxencbE7gfRn87pKEZpVqxr6jgJ8rF6in
DrrB56cm1NUSl4Uin5So0jgQokrQolkBWRlLzTTjVlwsG6eTVkAvvd23AEMpZOVM
GcdLu+xNmlx+d5k2mrMWf6rP71psqRfHVIkb9KaVUxAneGc1dA/fDG+Nm5dkyg0A
Vn6sXua46Lj16FWFFV04m+o93ChFBlcXYKgXPdd1PpUynW+79vt8IJraZuZAJ+85
nioXiUHOTkLrNkCYad2to2snCTIDExtrY40MqY27Vtn0hoKz5REt4LGe+sxJMhIL
KMUcH8AuULXPMbc317T1hpp7x+rEhjZI4OX9qhBiCP7xpEQX5m3zmOIJw5Y4/XCf
OHOvJVECIXpDMV36Lul2mJFape9wBrzZiiGtMHV3HsXEPxMFK+e8cgLXhbOg2ICI
TvulTApRkZkTYBMoTEeyls1mc5vLs8CE8AYCPTvFf6ogeV7t8AVLLgISNKGp0XBf
//jGhUmy9iYKGaac0oTs2CTU5+wMPq1HRIK1GorioQrXJYfjWt5Agwwk/JHDRnUp
cX2xnlmXdL74YTKS+25kltXh0y3PG3xRKHvv2TdH42DMXxB258Wzhvai5Vjfv5/J
QwZ4HFenmpac1mSQEa4w3KRMPvw5FNJXSDOzgeWzLxgcgYyH/vQikWEXRpBBlxJ/
vTcSsF6KP2VOZ/az0AsxaJo2HV5fZyZJnABaDA3AfxZN8jD0MN22PPDf/w6FXuug
ExE9ehMQtj724b50HtiZMyViju3GIdBw17sNdbR/mWLvIzjTxWwRmdHZPbeOTZa/
yzfD+66rBQyI6qQhIhfTOv6XP/+8wzsKWaqFDWu2aZuly++S+BxmGfo2dVdBgBGP
jKEWlsGK/yOGbzkHRXxhX/m1G1j4wuo6wTmoG+JcaQvoVRgP5/lIquOocel+Cb/h
iBWbG0MoQ6gHLx2utc6Qcf2A3hPNlpTG2Tw4jlaq+dhsaKe5JHcItuI+NqEJaJVE
Ew5ullmr7Oqtv7BTQQ0m2H0pYRXckTXLnAdejtlcFBRAqL/hdLVw2CoJxqD48Y7i
9h8RJ6ILZJLIxTxvwSMjUmGYxY4S9kVAJvT4BA8UVL3AmL/AR1YpGLqaKtFW+QYC
RllpIVHAg4WhAGxlFNoG9K7A6LRchy8fnTPGM39nPW7r4fPrz+rlGIe3cotN3tPS
QeA2TT6Q+rehdUWBac2Bf5QZC2AdGaJJjSPZlr14WXZB14SyR9pCabs93LcekBKA
c+BEJz9nK7P83WreYkxvzAz8Vpk5nK/AXYonYWJRKNZVa8AYL95nVkeEUDj9binp
5GukVJIY5kWDm34KmaDqMhPwZed/BY7+tDGtvP2kYj8u0INovzjVbpY8lFZQqkf1
kyo+f+TvbabkoHzsV/+O5bX0K+QhrVdTuML1nibvqVvaCfEzzIO1rWTJYuMDhD4o
lLligIscLTuNiLcXkT6/sn1hVvwH7iNXgSx48FxY9ezLuq/5148LwjUx6mFg1lri
I/W7ZLftTZ9hRtrXZo72K/sQ9WGP5mgnm4UTH1Vu2zMzHZ7JL7e7i9d3BcpS8vuf
QPqxLquurA3ZxzJ2xSP60ng05FVA5TjweA6xyW2b5euR8JFWZ2t9H2K5sy9vQd0z
crCsoYfUjJONtdmkXSLkImiT7HJPsg9kkoFyPnSIH9vQ+LpqWcUru19p0agpw7hw
s1+BsxQasXw1SSgK1t/NA+zyBCFb23X9sSTjQXknOU1RQbAV2w9HTgOPW6f544vl
ZSU6uwiHq0rDstOZPDnSFG9RkeW6jwetcUIU0tAQAS5Bjp6XAUA5HrWtCy8sN7UD
YN7Yk9IjeSPPbTZwdfU+6QIIFOhvalKEnG4UBxJi00XlYziuzpAyYw+7H4Vcjb/Z
XZ7YDuRJyVALzk34ljd77TnSv4pZVIWrQ6EZehYAj00Yimqm2fbKE4+bTbGHFQAT
qF4GAFLqWiUEtFBYH+qPzG+7fCo2Q8L8z9AcCct41+a9WrXCnYAkof4Z4sqqBAr8
lC+mVOfY3PSrzapJFtZsxNdsN5o6/9EqxQua8r3VTiD2C0qVg7qhnnJrDN4Qum2M
qf42iz2GktaY3OqkTt/lLhH0cp05FBlXLBk9wvsDXEcKWmGdBA7FRqoer8zfQtCC
qBu3LCgdbC4/HkZHzGZ6LOLfDlRAGz5mzsW+5HTRTw5Ly9m2WbZHj1/3Lk01NXHN
1kR9S1v8AYIvkXlQ3SLcoaYsAkVdQ8DUZzD5TRa0kQX0Sa68ZVfKYStMRRaZP59K
`protect END_PROTECTED
