`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UVzu2mYkzOQRCi7P0tSep++KombSNn9bgorxDT9Ow+ZL6j/lRUYtkKAZQfkP5zkh
HBtsXuOTJb4VfiTjYRYx4s3x4KC1kuQEY6CSGsANUd3W3Q0R4x+iLW62W+hhdMn9
eCwOM/OYQVKw8BTDx6fbNoGoMMCflnQrC6Arvl93M9J3eMl92bgDKN5D44pV3mD6
+ioPaVn49bYb/2ldcamkiEXF1RVQQmgYVM3IY0n5C2NYdGVdFxC+TyIqv5ppTz5r
gxa8uTJsGDDGwWXFGygOGGLsTCu3rfh8uXa/+8t9B9+TmEgQA/8ikK7RtVuvVOlF
9CbXY8/uNdaVwhIbpYcO+pNONTjkb79/1bxkfcmzdDqQ3HaEeuZrAVtT2KsGAuY/
TclyxsqCT7joMlFCNzBqlOckmkHp8/pUtfNKh69D0J5G3CgOpng/iT2ib9xcDtn9
RATncMPWyAAyVamzkTigOpglnV8SzHMHjz1BdTO9zwsdotnjLHmR0DB5Zf0iRz/P
XK+RQxJKO4SEaMKB+tbGplGvPXkHDnNLo3IZ6ZVwILWtTXKrkLmZlDN2j1FIwHQQ
PcZdu0Gf4oz0ZKODPNHGK3fZjXclRojH1bNN0gYxb5vMyyjRirPQ6sxQs//ZTvXJ
KizEgzCGZjxOvJ5zU9+CqRq71y3+8ATnf22cHleJgvxECdpkQgAn+NOcxn5ejD2d
luU6M1fihAquNtHWSSGB1/uURyId+W6rEkDxpvL8iR+SVHtD1Gn4E5MPBc1fTie9
jpNrC7uC3eJcf6Yl+2ThpqtK33P3ruOWaoRhABtf+sZxx0VfbJi1o9e2l0irFOjr
agOpNJnToIPkfIoOYrhbsoE8yslDD2QG/fT/IMU2d83aLFPGAlbAdkzQj0t/jmUn
`protect END_PROTECTED
