`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H46sTwERI2rjmHoBJUBWA3aFcVLZs9hNu9NYeG2s8ILQGLCzRqsta3cyWbELKTm0
VAJK97TfoapxoEZC3+c+DPgERLEpPHlRO9Lek72Oc7cz4FW554tW796Z2Vk+5aM4
71J7vL7PVm0NdCO5eKjz/e2P45p4NcFzlw60izFFNoItaImE1p1DLVjQG21HmhgM
mCARn10FpBtWNYwqSCHSsWwK2TEd8ZW3gG2zPqJVcd9ozcD5V+w0l1P86KX85HdJ
2KFKUNRNiIfuRmNy901+oHidZqQoVxID/zpvUMbwW3vKFgkdSfoOmkQjiOlqpG5X
gEkvEZCwTsj1V1UC6e03WaBj7rn7p374IIdam27rzxgQBVyokIv9fCCj2Mz7UqDY
YWPbnwgQKMKtOMKfgAq6uSC4D3nghxtQJ+I3RV9WacYSVvEudyslZBD+vw0MhJeo
pRGEmEZNaq0f1X1HrWQOR5UcZmR4IEfs3WXLRJ4knqIcJr8CIQtr47hMm3HQ6XNx
u7s+LF5Cou4LygdUDjL1j3qINQvY+OgSCJ8gH/z95Kc/WI94pHVUgayPalll5JFL
i9yHvkjsXViSmjQdSKp+3eSYU2ZfMvdtyp0+C3mXjlGwmWtHlYOPDr2OEwQLibsd
gfDa2g9ibIV5VPIQTp1YLSWuQrNMxSRv/IhC04986U96MSHd6WNkCu2YqaRnRKnu
GxdkG8CPwfHHFfdyLlXqEoyTjsRUZpr0lt/WBIFAt7kVpmoxVUatebmw8Dz+1F1g
1zrNci7jvj+SsZBjdO+D7ccWzBXrG1NH2NyKuoKyMGsnlGufpzNSN2+zYTh56heF
T5mXJxt8wNiyokcrCdH/LTIhDxDixoXO2D/gJTr8+SA=
`protect END_PROTECTED
