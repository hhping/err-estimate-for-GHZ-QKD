`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwChcA8C7wiBTKwMz3NMlokkhcBC5aKiDWm9LaeiJ3rguBNB/Yw9UtrFQu1qU+4R
InMQt6PP0hd16VtXWw+H/HhLuE64/bCKCiyKfCnczxTlc638yx2+/Z8e6OR9yYmr
NneYURQPxfXIucvuQ4J//TjfC0ux0zh2GkTlZgjmaqliYt2Twoxq2FmtdQ2XzG7x
dxZbsIg4j5RLtNecfZMPDxOzc9wqJ4cNxWNOfFX5Y7rOV/ytDEz42/69mGZHWsXT
TtE7BrRINnqWjvB6qbnb4lPzQEMcbraxicUfxBbodE/v85Wof8VpLHaof+mX42h7
EMRBT5DLGPceq46/8V02T34VeSdl54AIwtfsUEwP22Vjguyp7u0V3W1IanuvM8ty
hy99pIWjBA9v8xyR14EfybxTD0KMUFLuGPFwjb+6LkIPQliEsRNThpc6orbMvp9O
zYakHXOc7qH6xHjfzD/T582q5IwRTDvdO+m/7nJz35TIU1V5Tr7SOuAWJZi2qRwR
dB6yI2N0HThpWD2VVPallMLOUAxk98qmg9nabesG635k48Ji02hIsEd0fRj9RlgE
/pIXra5ITdZjCGpdXPDfF5GEd4MYSsXuoJDk3Y7cfw4YeA/akrSEHk9eicbQgm34
3jbFa5LRaFAJnaH4oqLIHh5dwwdfg8P8V/AAWYF73sEpPJdg5uv9TE2lGJC9t8qS
UxQhqsP8iPlHS4XT4hwuBVwHxSkwspT2zMpp4669A6lSsm2tKiCeZdO4JLMZGxSE
Bckini3OX8FoL/ZNPsH26DvP9vaOezrLEfgUs/QCaXDzV+6lWkVsXI0AtJW0Q89E
o26AjkVUAaehgpm4X+iZX8aec26hb7vaPzUcZjnfNGXUbsAI0Cx559fjdakKJSbN
bnE019T/kk3N5eIbF9qvan0X2xTkyEngBunPA8Phq8QSAi/IspGkpp9geCVP+Den
CYTs5N1xEMQsk8Tlz+tbuyckBLz3Ainkj5R4MjPmOxdB/aEeSYIwIVI+Wqc31Zg8
QEafvRyBV0jDqjsT/1Wx/r5Z/hTtUUi8I1yrsZpBHiB0BuAph/H4KFYarH/FwBpG
5NxBzHMc1yhT1yfhyLIUwjlqWz2Io6zlQ/+Kntnp3z8AeI3ISklufyxFb+d7UEgC
fVKSUGtLHeWBn5BCJb4gTT7jmmeRcXmyQx0jyy0/8rhZFQUlvoX4NmA33UZ3eeTe
vp7Shu2kcNfRNq2xREwaHPSt98P7GU5ugYQHlp94giSoUStjZAcuc+OK0B8b7UXB
42t2kSX4cIM2kalLPO6VStTK+p1+T2I/chL2JAYSioOwBh6SddoxcsWv3mShO+n4
5aegBBcW+Yhabbfr1Yot1zOyUeHvGAuBEwsWwWblRAjOFTX5QiI7fjCYXd4sYAeK
M2RxDYqqS6hdxLKGh7AEg4gs6ObjU0W53jCsCDeoq72yoySx8qXxQSRFOjM9QrrH
KgCkRFJs3yC/y1811NtoLsK3Fgal4++2U6UQd6PgGXKM3g8s9CYSJ4Rb1bJ5rHqb
eJIxP6k6UQCUjaZneuim1Qbe5JWT3vIKIOxw+n/2qU6HxolMXa2UA0EHILqX93Wi
J3Bzni5J3BjXeJetA8hyMpjKT7P4b+kys73met/fC+2684e1kFXf63wRbfqc7Cxo
w5r+emYiShSvdbKWmwAFjI5uKU/mFBwOVbCBc0v/si3hBie/+hytJ1Nu+LE1PHZM
+ltsB0q2bWTL/mWKkqUD8q3X94oLVvpoYofwD4dpxdktxmvAK06J/HmOg6led7Ad
Zy0UM+H11KcCTuB+7OheN/CSFj2ylQWM4wZlbJYrzNV1WIdGdse2VDi2MABme2nN
9vi8TEQ/07vZRg7UTIE4QvVdNwU8qalfIddwzCrdKq9cLmdQQNv5HtwdeAsn5hfl
HGpK3TifKj+PGU8R9uOMRqX/bj8rXrP/fppaETmbaD00ifUzg+HPr+ZkaCBNHVk2
HaHEjmlLBl4f4Nssq/lmLCZg6EY6xn8F8iEOJUCLIkGV9gZ48v+HfPxAkTyoLo82
xQo8k+XF/AdzLUGP+kslm4cEyImptZQsBJZGSUePub/qlufp2aDTOKbuQ8J86sim
JJxeVNV8HY5/kTox/hsWwgaU0CUY30Kmd+BXN1SDtN89bTTiMkDmNo8fhx2iGj4h
LlDRFL7lpI7vss/cKkSQVhHK5eBsSLwYTLTORc9o+0nK4mB/dtlUXBrut0vLFjr8
w4KZhPXZBcxCagAFgKTmgAaiaOpsoCcvT6XrVnTWVgMSewaabSvlp0DQxZMBUQo2
lZeTJBgNHo5k8njHPFGCRmSuwXyU+ocdaol4XtUCaqWU3i/aEP2VSJ72NZVk8S0X
kGOz+AE/nty7NT5/Y42HMomugxsH516cpFvEPKLNRQcFxiEVuVSoDuRbRa1jIaZ+
lkX2XGcIOtKhF0qe++/+A0ze+f6nMWz3MIFdJcYohb4nyZVqsJn+gLdkHvI7w4Iq
d04AV5almUOlji7grbrTwJBhyQjl2nT1idrp8toVx8CAI7+DXJ2vrhEAKCFsp0DF
nfrr/E4e926QUuiNaX68yoajlMXVgC8utM8Dhr4nIVZN989aHBTjfCM3T2k3vTFZ
qAZl0xaW9hTvAJaMkj1gduxjfCsufeZA53apeQa9Q7vcYbrQsLjVt+Z7kt7NA5O5
cXcaKEXFTaashmtld4n4yoqUPyEczbudsQ6KM+O2NHlODvSJSAxPkOESCEKxli12
mOfQsMMF9nW9B52OhNsLEeU+zU/D+jRzOoJWIlfWC0fm1qoaJLjjgFIvn8GBQc9n
FwdF+SbFBHaf3/fYSE5uONf9QunqvjvlHTHLjNaopzbPPdwuYm0JgH2iHJDqCEVT
dltV2KSEpxm4GEHlyzi9wHOc4BZoaFgGpHQkQiXWtV327LYcEiVEjzorNuG3kcDx
/OMUUWiZy+xZJD3BUC+INi2eC9JQbTx2VIenxp5jc7UGsoN0HJyetURGA17f5kxk
+Fr8qthTCrKvPqs2eY6kZIfHZne2ljs209rQ3INj+9G0xd9QDkjTwOXH/VteBrcv
vhwd84omdGfrm8vZU2MxfcuRd6Ahk4du5wC9/GIoxGBS8ZCs8rx/40Z30TN0PHTZ
2qCvNpzQuxOEfPvy0mPJ5rc9Q1MF0nmUAGdtIVREGd0tCD6vuFnuHBmDmz880/mT
Px2Q/oclJCfPxJOvx7CbdFE5GWOOrV4jKPx4Ne29+dxLQyz++qvqx04R6D/NuatA
xie+B2g3VZ+esB10cL2EirXj/gJlMMlu8KKFvfxCanj+Qmf87gCifVWdqDGwVOVM
tS/wribcIAxcN7UEKMcA+g8p6xQlZtJm+f8e9arya50=
`protect END_PROTECTED
