`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ScxYLxZ86S5Y0LanRP3rVIC2TST8GIpzAnqex6XgkfqfzdnhOyXYlMznY7KZcfVg
ht38kMFSdTkFPwiD2RejwJS6TyTYhi4d8Pu45CvIpd65TaSNk2u8bF4xLCfrtHnH
r4GIX7qYUftKO5QaCmWYeX8hMyqQhHMwYgM8rKSxNWYYfAvB5q2LtvMiJJCQdqit
U9CtgbFpJdVQ6rt+cNFxuDY9YQgIWpB7szPhtfT1+srz9FXEXVBVP5r3+RLqHTb3
UTuOcBlp/bh0CtR97xO7OLKy2NW0L0srLk7+oSuqMIVfLdOAefub8Xgzg9Z8P1cM
D4hvZ/5yFoCiS9rgUw2stSwoEHhvxfe5wIujliVeZoN25ekB2Kx98mUSloCudmlX
i9jfBIDy+wYxeDlZNKbSO/Y6yWEIPxLCuDBugytNESyuMaq9EWOE0PGj3QjYL0T9
xmZeDd8cr9DfAcxvyj3ijEPmknA0X+BBm+NRDareAZ5ZS3rI5me/7t6Llu+rxa5O
dcCkvzhLyvVAGvdAjJIOMKozI1C5+5ygxV9LJA9tYBF1g8qRCGMyzuo1g7g6kh8H
Vcn4b//iWsGyAKw+bW9q/1Kv7vQSZWRgVjeKyTlR38CYdc6EKJEqY9mSzBFCXH8D
hMi2cDRUjQyBoJrtuvtEUoIH6CeJDz5B8lgy9aKw9Iv07Od/LlWc6yZJaG1l4oky
fG3+anO6ZeYq0KUFobALDB6q0/DPeZcz7gv1s0nrj38kGk+UhP1J7KPABS4dxfe6
A3pnOYzEOgJLUPFRR+ORtj4w3gk677corIafLGK5TPZoQTL/bcyk+KvbMX6fpOqB
qwnyKlTGvBMeP03Tp5Z4Dud+e1kVspe96cErCm+s0kvESuuokeI9lgNLvpKI1Csu
hR/p6pZ8u8KOtqmHpUDbfFbQVgmZ8g7FzD6UUvA8J3WVx7WRBIV9WmPY3F3HcmiW
/O6tExJkyp41duUfYQZVd2Nt8Up62UG8Ju2geTf3cB7g5bflBA0M7W87HP7ZLkCB
VBwMD5cenh15VsghUB3ZpXATbpSYVtpE82XCvCIGxAEDi51Bi8uwfwW97m4XNewf
WCGOgbDTGe4ND8JtEu4X/JF07CeeAFMrv0zMu+ZEaqNpCCjhgIKCAkKVy5AUIFVm
rVsXD/fCfoRtntozCqIQJfy/nxfJhW0nuHnpTsPVUOVqY0y9ecclqddtfSB90b+P
LdB1MuWQLoG/ilpOlBOvgZ7H0p9gQDKIuqOXAPrTEk12ewOctm6DYgXkof7KECni
r+PzyzQ3bwA/PIi+k8hPrJnjQnVD49FxKFCgVWg7303i9gDiOJVR4921yvrotM/x
WIOWMHE/HvAp1uN7SmTK71nVX5E50e+BbsDP7AAIaQK11vHmwybvfYf5MxQljGKo
hgxEgLlTx3hZlgRhCObO9ONiPj7Z2TRH8XDIinZPjJXgJkrmkX2ZseHqA/zwPy6k
/+La+Tw5JtUQY7dGd7BSqshwIicilUh2egT1bb95a6y7rSs6+Q7O/sQ+BZuHrzqO
O9HNWBVerIsGqJe4aSUgPQ7Tb2UtDFmPZbQo+SwAadKh0CzmvrEr8Xu2Bm2eMjQ5
OJMWl/EYAZU8NHTy3fGC8esOxCmZC6LdbCq8AMM9309PuNt5iGY3dDuSG2UlwNkG
0kVurSG8JDtLBwp+paw5j6wt+6lhumIm5hrwbuTTETAbwNqdd0Sps+o6yvU7crs/
95/uE4L+wzlbsm1nBgpLP32erXvMRFFm/nz3a2yf9E1k7Qq9nSX0tNcG6Lo6zHdM
r41m5L/VZ09i5qUWQ7DFDLYuSeoTWeyRQmtaHxn1T6wRLYYvgDDjy9gPGm9/6SaZ
hxh3y87V/C+WvcpyZdpaHEc+rC5pZm5LLuUXxDYgW/fUV5qkJPfqG1sF+wsd3RF4
DaORvIIMH468ZAHpTtr9jsDL0wskP3OH45z58a29IeFEzQ+VMjz7i3mDUiYSKEA8
TxP90o1mZdAF4SmoGg7ry4ak6hsKp0FHNUnVKPMNnEE7l3Yhfx8dHUtimQDHohIp
Txln7mm9XFUSvgkKTirpQjnvMvs7tiKA+sP9MTQaKPTV3ewZMDyE5gv7OLdwh8w2
stkqHQJW2WU6MWRdDjON5M/IDgDbJzbApAnZK/IEM9Ql/YBp6g+V/offrcDMOmIf
+rIy2Fwbq1AwdSFHJf1+KyFodKn34qi0tu7PN9UeErGyB0WexpBFCZs9M5nLuWw2
gNUwMcdFZ8lq7wyML2ENMRu1lVcoC5P/4RLwAUEt8JRNjzRGvvXPWbGaQRwrYEa7
qeK0xEURb8DqXAO2dT796WVKCqf2A6DKDobNKJWmsr9KlfYQaoDqBN3dVmFkP8dc
xXxtNVQD2H+1P79LzPKatXKx9VVW7XTI+62dYLo27EcUtQlcLGGHk7M3e+Z39qkO
F1CYYbtlb5PZIdJDivL6Fq8ZH7nVW/crym+VJr+LW4S3JSMAS43dPurNAxNU0et4
RSKEh3dT0PWrZ1+0BbP4wJuk88xlu7vsC6NkpJV8RMoQzZMZyxwmLIDNwzaSmkpO
2s10K1YHkp6Ez/2rE0lDJBjJxB7tEBT7UvmqCXYIoEFlOw9TLQspGgzyUUgfvhJu
Rh1Q+t8LQOo/TNHaEVdib9crjfFjmedXnAjfHjRCeOnqZ3PIx8wDovt39HUglGVk
tLsZoJgeVRuAfwt6k9dRLLELAcRimj1KSXNX2Qg1lo0I2UxpSAbFFG3GkYscozJd
GH+jDzjMSNVlSw5COD8CSofQTOMQ8+8D8YyKPrH3UW/LXK5LnM0nVhP/X1t14k32
+Yu381g8tvL/DJ2/g8igAwQqU1C+W/eXVHaoaUN7JmZaXgPekcGL1gEe+CamOngF
Eh1vAAibEHAh+TKxXqyMvmDqJZ+BiAo+iBCy9ruy9/RrvLwJiuiidcoFTLixCMfJ
7uuz4aj6eP5j8kHdDaveUwzEP3yoXdtVxH9elx50JMikK3wdvL7xLTVi0PT1LrjL
vghhGiLQlcSGpOW/2ueREL+r/DjgmaHC/lp4rKmTzd0ZTaLCyBunewLXnhykw5oV
CJ+i3Oi1+CA+enljqdlvFFXcobjks5t6yY/ludMGgOprjfTR9Wi0BogD11uwIiJv
eStvsFA43GU6knAFaglKmKCtE8aqkncGEEKAxu8hIxAY6OFf/3KLdRYGd5vz+fCo
z+ozOgDT/Ua+OR6F+7WklLGgWVIwfnwK+8bqFfl4U9sKUY7URSvKqHZuQPVKfKTp
ZDj6h3mSr8ewVNtyPNfyZaRhT4A01jBMtaht/3mjvhl7aUV5+N8RKQAZ9IH93Q2+
KBGe+wkAkK6/+RP4NzWgzu8aqOJbJEoFwe+wj+yhmSkf8In37GRWPYOtQfhJwrez
zPGK++bb03pCwNS1Tq7yn647thiv3+Adfd5fpfsVMZAgCXFc9mRlOuLalnkzycTY
rah5icoFYlf0U5vrgrBJO8IYTE7UOlFfOdlJwtT2bdPFhLvYjcTc7dlDy3zwT2lr
3yMy3vX9drMLVkc2GEEB/YESM8Aw0IXDKmRuEZMXBvYhCyKoPrUhPMBP/wD2nM3h
uRzsDckcmdt+5lk6Ggj1dmddSRvRQqBDE2ZV74QJRHbfRk2UAyLH7anW3GP8H4FD
o7hy8raCpmF7GS/OMaBj+Fx1GoHemNJY5vrQBIj0UGFzcvfePYHogekwgfncY8HW
NObqVvFw7MWonFlyhvZMCBg4aHNzQDgEgmndyNPGacG7dAjIl3uY7dsRrTmFJDS1
QSjOAUdAEolDy1JCDlwRMVX49ZHif/YLSktlSHigikaK9reW9cvhwM0C71BZfH8t
qJCWDWIPs44+L53V1qBfouf+Vz71YzMOxR2m5XKzog7s1MplZ4yebQ4RYlsVTvHJ
0mGfTVRASZN9+C+lJ/K8GqB3aK9JKWuERj2hnbGpWKiRPEx7kyXkjq0Vny2BbSHj
OecY5JaHNqcvmLUTObuYkE4yTKWSUzrNddRdlfpvMv/1exig+dVl9wKQYPmfayM1
P8Zd1va4oOwWJImHvJ2Oh3UQMA+tN/v+acD8jRAdWEGJvTITQYg8IydRSRWHjjED
imSCGj2wywm547qNLtCpFg==
`protect END_PROTECTED
