`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VXRAMcLRTCUQvHJHQ6hsMkkyPv2yL44QdJ2JQoz/YtoWaJEZF63AqGYRaZMw/Ta
+E9kRumPXwTIfHlIrNs5Sps5qJykLQXzNEToE2JH95Px7K4tz+VG1ldKny7rRygk
UcAi5ipTSbC701QSg4+a7t32w5rScq6w0dAadQdk1m/qnfrReBUYuaAjRA6tX/oa
ywe0NdTawxKlTndNBTUeqmx6W0k226J+xi6y+OwOf3D2ChutzCsi1cUEn3Xp9GUG
ZlavODhvpVwWmzVP4oEFlk59GrAwYD0slO8LWWXkpVUt19wZZmIlyTzn6awnkB7o
OwoDJkFSdu0jBGiQuzXUIxGAPY5tVdzoGOI7r/0Jkl/mPlRHEoL7B6bWjEaT9Fgw
/pWg/jJprZUug1a8GkFXSFcQJ1a25D2S37rhvt31f9AZ0ASPIpQJUW6p/fXddlja
jz6WgFHhBvsF+BO0U4lfxAPaXFBtODfMjOjWQKvQuPkFe/hhy99PfR0NFZJQhR0p
loq+hxLrQpTd3zkk3i+i4SLFod8bVGB55FHpSJSokmUfRp97l/TwAteAEE20YLkl
QevSo1AaSFcFFtv9QPLhhpWQWqVIqdM5P01+gM8u9gPoz/y+8iKcI5pfSza3tBuI
6oejCCdAD1/l1b1zzDqmtCXFgdkO9NfvmjmhAssEfhDt9z1/40B8Yt6rMmX/HQ9e
I9GnmbBK4OptQwENk8Yta+wLhEyQgqxlWI6h8ONEX3EBDrBqPygkHz7Rrh5TnOd1
VBHMz3ag/TWNk/17bzyqVpEmgB21GfkjVjshGZTkFYTmBAV4kU68dVNZqFXQxGCR
xuLRrRXG/DaZNlliU08Utm2FXr4OtfSJXNyH/eiWKexmuO0xp9U9hX1oBhJxm3c9
7zbUuDHLpdHo948Dxwz3pcP3CG/uBKIbNGkiqMelon+YKEU1xHk/Jet5VommPxEm
71tLZ95BTlk6tuWYP6qx0+B46wZ4tLoUihHAJ1I+1YLJtAUTvpe4xlsQPLsC8v/4
QJJ+LGfDz5Jx2Imc/Eok2NSbexZY5PSmb3YFC+Jg9FYv/6Sb78RuCwMBrOTCi1f1
+DRwnU09uJzI4qW2C7553NiWklVMxTf86MRttaQFELhEG+qO8qi1jvLX43PYjZqx
LmeXWUwxNlycvRLhCtG0i07yvCnQB+dNeDp+BMfTxdMIWINvgw7eh1kojgN69I5u
7wIvz2swr2hRHw9U0JlWe0b7Y/BxZ1AIxzhcx37EcHXmyGWz9tMunq12k8pvcGwY
GDGPg/DOGGt36s8Uv5c7KhZx2Cbv0hoh1iWC0XyIEkF91mR1PiuU2fmw2ASaYtH8
fVvwlggrxwHcvkQR/qpgGkjguPs8DTGBx6fGreuvsgbzmapqOEJy29LiWcr13FQI
kddmBrGdQ29t/KERngVyEq1DjUzaFhjZ211LLyGsou8rumGk1P9vn7yatK40L8aI
+ynwUzwqU1YduCoS0LbM6ag+5gxyDSH5+nfJqf3XFROGuB17tT4NJ74YJ/ZrAPuM
oTbxc6MemCGjueoIO0ZtEGd+1K6uIQGOwTAtAmqg33OAJs0vnrGxAsz2vu/t+5mC
fzMich1hQFSnLB4+p5QnLzqbtdsZO8WjWTYcS5Q9T7tnJWwUzaABF/hI9sr+9ai8
xZtfanwztCmmZgWxELPBrpX436+NMHX0owf29068Rijve6NlIiswfGGeWhTWhR6Q
G+Nuf/2RMC0ve4BsjY5OciQ4rMM41yIN96NhaW+tMMBuf6TLmohTK4P++EtqRTSE
40YPFiIdbFP3nRvqhsQxyHCUt0Pp35w7ya5JCg7GcCnLzfvrTVT064m60aC4ZzUs
NCDQKzVkcWRWh40tzs9MMLRKgnn8dI1U3Ulv2llhblghjyz3eSmxxsyZ94BoxBBO
8I6K+5cERqKJJc4mx8wHvKkiO+MxHKZLBP+BoC/KTwnuOQXozbB1qSn1qfdwTEzr
eE+Y90mODW0gMLiK8ts31Q==
`protect END_PROTECTED
