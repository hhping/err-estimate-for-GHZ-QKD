`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GnsGQjtWl5Jz4ngeNTn3Xxy5ouzrI15/5tcdR6kaUA8Zo9tKZKARtbRSdcM7fsc8
btYzlxTqUmqaXxQmDrAG859I7dfqtNIHJ1bl8ilFKA4pY71cl9kJ/0Mquo1GKziy
bWadnQ9mLi1xCGfiG75j4uNdiGXC7g1MtbICKnWaCC1tFNulOHAr5S/IPKWXRzkW
DkKifGPPnNW66MECmkfV7upYvaVQIhPtARoJ7niBgldplTQhbzI/dqroDRHiUU4P
YiJDXAwwgRx+rSfNizxE8JgEpNjpUDt3AZy7vxlEdGwEqaW96dQWjCxbBJnJcPJR
R/eQgl2oMONpdMxB/avHb/AaBK5y4IehjscuJAp7e+oEeSvDqVsZpvXSjNBdF7VP
WqWr582mV8TXM2hyxCXYpcWCmf9u8nFfMa2MRsqliW6JflfYAiLWQ41Hq+WrlixU
DtPxgKGzzIGzOhYpcWm6+7HYjxdBoM3fpk6D7HP/r0awmgSm+Z8WVxHMlkimk3Vz
7EKgrfCacIS3GJBNuZ0qg27bxQLE/ZB1IJbGxoWWV3+YXupAwxAAUA4FXFbUG5Uo
siFZAwTt2VYa8a3lvozst/rIDmiXXI3eTcvwjcEE/nKn3L0P98Bcpn7V41TGS2OI
ILX/ru6aN/Lb8QB04r8OvtY4iyOA2T+aLZo97nlZmGrRPpe8snxpGGHCVmjGBCum
n0zk3L0+UUYLlnjxEJzJZAacb7+Hh79ZD5blyg3naLwydIBVwV59P9Q6VaWdPXTV
TQNqVXE1zMwqcJBC/ODlz4LHJLBOMFGVLF9AWqdTBcNNNsQ7hb/JR+6Y8pqmbcKy
tX4UUSH0AqglbMGr4eFl80ChHmEikHPGE5Y/NZKtVqipiCWZwWwxVnJ9DK2//U07
jML2d96ml3lA8/+OGH+BrPFsW9hI6ym5O2pTKWiyFbkW0Js5BG6hzC7QZ+omRD3e
hlrB/v6nxqhWmdJMOyW6HhC0JxDu+eH8bXkPLOeanWXFt5V+pRrwwnmMlppZmRFr
4u7ZNgNgky/x/MusggCmsDYB6P71x/Xdk1y3V82WFOj54CGBwVbyniLU4kypBAxO
LsNGPZdl1WBryBBG1TH33EtgdVXay0bUgHugRbyAqkTwM2SvFyNab21SMvOgS/xj
nkOkRJPOqiH4M/J3Ud0aj09nZBl6JPpTVzhBakHKoN7W8kepCTShUKMHIdK9ojkz
/6BMR6X0pivys6gik6hSK4l+v0aw6uOOzgYrO4ZTYOZPKRSRkr4mrkCc7VZHV4GZ
KNPIpbJEFvMtzQHgziK3XP5eCYV/4Kf53QnH45as1cSg0M2ESSeQhLJ5UZGYmzSX
q1tPQVaXq4BgdM1o+bM7G/nr3+qjanKQxXOM5jrZfDcNpMhIoMKkBWHqc8hb+IRC
vq0enKocGCvctKW8JUiSba8My5ljA3GgdqoX63s0+3DcqaRgmVjf2nR3q98HGK1T
JeXiZLx4y7bZZfCcFsH3lDtgv7Bv8ejqRtOFvYxyPDYsd4WfXDt17g0zwGEoginf
GbhPXyICI8UczChwBysbrS7xXWy9qbOzkviH1g3/OU9tETclp/6lAhj9vZsM2+Qr
E37tyaRcQwCH/OAwIeD6Kg==
`protect END_PROTECTED
