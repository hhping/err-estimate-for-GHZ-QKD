`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eSQR3c8se2FmD+sc3BtOLUkf6/PgNYy0WTGF0Zq41M8KjwtI6A4IME/0g+KWqljY
Mhd5zVNkwHA5U1yAEBfMwd1KDSq+5m3c9FaebfmcRn4+jdRzYVZtTfef93U3+wju
HDoH2aC7yolgJhnhCKhy5bvH0TSy0BXXMlStFZuU0bBKQ1nntAMN882DO7MXx088
mxB97Y8S+avU+OEPLDZ6B4h2s6UbfmPkduLhofpTsHxbSWre2CK0RUfAgNTKqmEB
NR3T1BmDAr8A6lCaXZnGr9gTH+MV4ZvMiSv3ez2SZXJoDx7JFapK6reV9QXUYoqc
8bhK6mL+FWAO8bH7KvafM4dOrqmfPAWfUxPDsUY52+qdCTbI1M4wxvMOaE+E80rV
3VBCaH2bIHvPJM/VG/qilU0aEb07Zqvf1rQuLS1VEyxVg1jnw0m68BoJjPUBVIJM
9S4Pp1hqQnsjaYLhnjaF26swv8HFcGWyZb/jAGAJoZJE99Sf5KioyfXmdChi8vVT
5GZSVkkeNvwTliAIe/nYh1bKA3gIW97lyeaKcPd0YRnXc5y9HZ9puf3R5eC9oHGb
`protect END_PROTECTED
