`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OS6JH3a/WFlaZPzX9Y522xYlo5Cq6a+JbBOEHIAD7zJOOl+mObHJrv9djNhlg/lb
hb6TPhDqMmB+daKhscRd77FsaK7qqbdW6ZXElvrczd8h6xk7DeWnELAtTE0bNVME
H+Q0WpQCFTW1Z069Eip5OBB/0InRm5xYu/HWbf4I8GoU9VAYlf5dQRnCecZZ4xDk
N8565m2gsuWBlBD6JK6+UNFga/tQNF383l7gT3+DIsNaqDcKkhqLPmA5fYoqTqxP
IfyIZf8ZERzxFzEcJn92vCleiSjz+TQJRbzeRJ9EG3VAizW7OjPB/OdE3HdFt709
xvBxZYZNCg3A219cZKSQkKf/7vIr/D+kBpD+B3iZuwUtRmg6/61T/jxzjpvSeGyS
FwHmFGD4tNpglM0/la3Pu1usi/UCCqSxG0NjEhSeBMTerES0g5bDrQsjlEmppM3q
UfBhf8rhFyp99uejLcUNXNgCrgyvxjA1pVzgqg/NzsWSd2HrU6arB41E0e/0geNg
p/WvP7/dtpCgrNnhhVAUoY0yfzddCIVBnTJviXQIEav3pxyv71yQ2ihYr1VKch3C
LbcnCbi70K4lalKEoCH+cVzOEDYS5SBj9D5uSI+vOXsDRKqpgFdG5G0c2woaxVoa
H+zcX2L1OSAsqQ8BDxBsvmk9xmf+06byT8J+Wdfueux8ns0qsSlPDiTXoaLozQnx
vwqPW6da510JHeIzstAhOM/z4V6EMxtftZKTojYSWePQacwQOzGYjChUtbIrK3ns
Nd/vUSBhjkxqXJqGZMVIjW74cdVufiFBJoEpv0hGSksN+/MWJ40A9+yGKl4w6VKH
nPwTPHshBsQJLf7Z3Wg0j6N7rbxC6hj+lpdgIU4WemILadxpye/OWW5K7ydohJRF
RXXMcvdlwj5dX7Zvx0kzZg/DgzxBZmOaeAhYGJIGT9L/nRaGsNFU7gYj8qN061Xp
AiFeHd33yl1E4Ca5x6Ht/YLKEJbW0YbhwONEOxMHZQ55+Mq1wkqcsvEH2pBz2EJJ
4G3drkVdDxxrB8CUgkI5NApnTednxqOY2aAUDvdJkRiIdcQmTcu2OBMxmUu0MwHQ
zvqyVXlth/hfmQ4LXric5bCQNka/TadESzy/QYa0wi8L3t3EZtTdicEDIU7o8aet
UQ0Gpxd3Myx4pm7hi2865e/JEUPC/JGqMwn9zQC9og5VVIQsXqAMYnEULUB6RynY
5/PzIQx0gQYxbo1fnXQb1qJeI0z8TXdJ5XbQoUhdwhBiKwpdyaeVthe20W0QH5Ku
cyFrpNI0z4epeuyDIdWvoQybSHvDQ6XfzpFi8lylKXo41HllXFBi15GQFPvvk3Oj
ljPcypmMLQLJ+Bc8c4DGn9/dok3MLu2FqLoFOK7MqsPkY5TfbNGXn6cz2nazwd4T
7gHMQ1OFQGyVJyVn6Nj/j305zB9dwTsgLf20SwwHx1GwPz0cSr/QQTE0nqzJEGcu
xfy4MULEGihFPfilRIJkLHtHYRU+m8+W3W4GNlo8v2iLTxtNPDj3SmZCYQk7wZoJ
alhmgCoKj1e7RFYpb8UhBVhbKvzsncgOxWjt2eebeLnlx0gdj8bYSJpEhoBcfLtO
Km/EDioBhUJ5Hpk86X3PqNX0pjy7bgLgqtkhwIIc2A5bL+ANSGmUf3anss+54EFX
AjSx7yL8Uiy9LXYduwj3E8wLzwKNYRjAYDXi1+gv6EPdQaBnlGIvEPhwEXUZx3kK
AGcJMBngiQB5P8Z82fRxBMpUaAAurd7wTAj1FV0CfdopgH+l0blEIawDY2eB5Ljz
g1R3bOAmlnzLyMHleaqwkNDJYjmlygxB7XOEe+ZF3ZE8oKnaAF7YLOLayekCm9mR
JC5TEQz0a7alw0NRblf+by6LkVygf74nVYTFSS/v8euieW/i0sG7r0M+Um4RWFbT
7sonxYhaGpr/jt/zkmM2m40aVhZcA1KISMC7Vt4Wyu4sm0lPhvrm30Ee8//L6Lvw
`protect END_PROTECTED
