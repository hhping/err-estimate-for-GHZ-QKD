`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYrSXKmY73/v88FlLbLhqAxGYTsyfWFkxsoAUrjb4Cci3buRrjWgVUp4IgGKx/mm
K7+4mO7ZK58VDGBp4zpZfXRrZaiAZhkKXn07vQbRyxAnfTHh2GAzzh+Su1Igp5JR
EyBM1qsgB8N2r8PFJiHizGMUiD8VgJTpbtteFcQemcvl/c1ipkvgTKP/0NY21OSf
KZGCsE7K2nBNjbeQb3qGogLamFgdfg9lKELmqdw5MZXSiGhOycl/LvGLVMDY4krM
XtLUJ/WMgqnFB4Ju5m5aPt4piE18jNoYdkcw9EDBCDG2QgRBTKlAicFQnH8COvzD
wgv0GdjhWpzTVm0aOP6BCBO+bSIkdFidu+HPeQ1WBF/foxc0Y6Vfm2m38l5zJFJD
ChVFdA3jFa/IMlCNj2kTlCtOIafca/YZVfKo7ELN6PT3WspDG916AnVOulwJ3Zk/
Qs6oGRwferVUTrDtFxw6AFLBTfcQFIFInxPzj9SdM+HYdg1qE9tWRa7cxc5OoOim
HX5a1qospLznqT9UYV2Ym/Xfg2Yq/kl9i4Gx6h0Ww3Bt2v02ogjNLnMNefaS5t3o
cFrFUQb20hpQapIBY8ER6c7UPoJ7TEPFfGWxJoZeSRqzH+w5bpE7Vqp46RRa7LRd
P98KwVu0u9HpjMJE8KiKcy7g+e5YSkl1nf2hNyH+N9LqOAMTFxCdQc2fiPegJm8A
KEr5t76BgTCLiZNkwXCfTm/lf6njR+iE8QDwo+trPSva83uMj4ZWdx2unWraQGR6
5Nv4KuJsZ6m4pDBiUADFuQ7o56p4q1UbnFMnP8ruPmWeb5EtMj0mQ282AlKaOPI5
yudTWU8gtRWYOar12Xd5qho07ENpaegqo7hIHAHD5NCkKD7kghDUznEQwAAlPvOO
xu/c9ao+GgpqBB1fdl+KaIQ0MVDuXLWKojgL4AzVmP8j0AW6aQxypKxsgIXhmOZS
AmvVVr9aVnXDVk3b7gI5Drakg8quJSinKqSrmRqKdjUSzxElss+6YjRiscxKpML2
zSSgpZM7ukfYI4rUvCkIILrGQTQs9dDdHtuRHovGpC1ZPGN/vbi/sk/YesCKUtgs
43lHqP5KgwQrBpo/ZQLO+1x0X4Ifn0GdX8H0V+4YhYPwfOetvl0ARaU38Mau0ATd
Ka8RkCYpwB3knrE7ue5cWS3+HB14fD30tVDi4MDCfKMb1Osc01sK2rvKdopDO/82
/eX8Fk49xdIoJP5E4zHX3+rZGeb9u42CkEtCrrPY3EFpH9JErfcflaYGxQB+pBy4
Ms7l9MWpVT87IsqYzeVthMlH8mqqxjfBh6oECSai7rJQjvPtVShldtf2jezHelgA
k7g4FnabStzp7CjYP4X/vZSMuDleP1LcHQIiCEqRFD+zCBNDnMAmPkmflN4LOweU
9nDXwet4NeP6gEHQrsoPUciCMOxgiYl4NfQvvcaH8/LTSERD/29TdDXDYpUd8NaK
oxzNbP+7B5E4Il/tghZMg4jyaxY6VcRUJX91dHxOIVj2l2suzdjISPJmt2XhTMAt
kIMrAT5cJWQ9adprfkj21uSJzuWYbvtSxp37DHOBFpMDThveIO2pimATlPzM1RHo
7mmuMNZ/DXLKQcpBsN2zy8zyhcBKzUbbQk5Klz0f4B4pWVAV8w0hcSyc1AxOrpTf
tuEqC6vo8gpuMY6XuzUEhIH6J21mZ8Vz0qA5OBkleQO0d+VR2E/GszAmszMWH+HA
8ljxhQ0Wek1HvQXdugMfKbLYTbIml0DVbmVQgUSyHM+bzbRXTXKd7uhmIBpQYxFx
XK9x9phLdVaTnJG83QLmuntM9dap/zpfl8etRRkxGFF8KQYHshtlB2FP1joFuezZ
IMc0wv5j0ENodWn5mzykZm1moF61QvmhTJNX9tkU0ubCk0bHmP203wsNUB4VEcXv
PiAVuKuiKJ3yRf91uGraOrZ1zksqilpF4IcFyge8jmcYMIko8Vmy0ucRWSTeLDhq
cddfiyH0y6eI4580IOGf9Qd3nFy0In+hO8cjU1DP6CQ8cwXJb9gj98QmDnDoQbyp
JyRTsZZFe0/rWNAbc32WcHJ6WKTYsCo23gUoOACl35vTL1ghMVa0pHacarVzSMX6
CR63teMVhsvYDSg3Lvi53WmbmvX8Le4YcS6VYbH4xIXTuA14kJHyTxdbuXy3/1og
AqP98DgyiI2dPDi87cwOTq/BHUWbicdM8yf3hVhUwsG7Evf/xS0doKkBPhDCe3Fa
p2O3A4SBUAcJ2wZ1kDgAq2TQ+HRVns5tQL22ImJb4Pf5edPt1aO2TfMKIwGRFcqH
zv2ZaIjUm5+uJNr7mh9sN4XSsIi90qANZcl7/mt+m02s3gjfqSm++PeTVCCYIPRs
+sN2PoDC7ilPevQw+6qMfDMZ7oCqDb1Rii8rYSzAlCJIHJcHATaOHUh3tRNrZD+A
gHjGI/e4mSzuBAnFjYLMWNTpyKPBFhoX2LiSNsdfE8Dw6F3wylRLk/lZususCMee
iazZED35GefVHrEj1M29ES+oem/fQ0BC90VhtK38uGZojP0blg3neU4UOJxM7Bqy
MoV+/a5Nme+FEKSefrHazHhxQorArF5kHeyTlr9OfYVm0MlJavdat9bloEdQOaW/
3t6fqFk4w9NDlZACJWb8FA7MN4zsZXqbGfWPNsMzEfW6RrbvmXovD5OVO0hoPapd
2SxDvstsyPfibY5dOIglAY24VpgmdSeF0kfQYzkrFrGS7i3duA96WLWzdPYsTlFj
dNptJTBlF5hLCXHVv83jrBXrdE0VFyggzkIb3pXvsZEg76nGd6igovmo0mbl/V5n
S0DiZchZHIHHPAcGvxfD08Hddt3ozC+1ikzm3Fal3p/3om0IvQunHR09qO9hr2pW
iasvua3g+TlHqpCmQPXOK6TGvyIhRJnZpVIF9MnCkg68ZFFCU80X5OAYH7sWHYZj
/WHQgLSAHV264J8a+tmDDXI07HjBb73zwHOZoh5p4H6e6TWtEJ2wQLzxrX5/CUzo
`protect END_PROTECTED
