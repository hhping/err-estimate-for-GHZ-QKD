`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJDVUuqQJiMvO4Q84NiDGINSBDrD1ldzosWnviQmWVtgLWJDUsT8AwBkEFuf1RgO
HitKA6wNmlRzMy3f0RNrhIzMZbmK7tJjoq0KjbV8n+JlIlusfVd4uJ4OWjy40Pm0
EU3X2lDiGk/yHVhTgYrbSc9E5HRAJQrO/LRmx3MfzObaCAmyy9E80lljypAZ6lVk
sOlvOFfGjfvDDfCQyYgY1jnq8Bz01oqfLdVe4qjeiByuMSzFLGPePuXnADStISlq
P0oZoeLaohBa0PlyLiA8dJBdjLhUKCg60TlXoLf3LYO2v4GaCUS7LdDH0s2mDjHm
qlPu7Gg+IJddin87OdU5Dh2O6bw8gfEEYrGMw3zsiaalz+4jy+mTf+Ldl6i8fPdl
IiEhIeMzxZHsv7NHFuTnW+qZPwLTKuyqxaidaycMVk1p8ipjg35bB7aY8R7lqifS
ASUO4YSQgwF+MwmZ39//uBZyvNMsm1/m7adYsM8Tqka0+k+md71RRQSLyr3K27xL
w8kmBTjV+SAxkL5A6BgespJ52SkV3t/gcsn/l+Fk50Ab/vlqdnM1luqUgPaHrKLX
f1FIHCkT3HKcraGQ0I8gYHNm6yjROKNgSineUDAeoEQYYsxkBQMxlSxW8bV2rNL5
mI1g4I2S5LgkZmmH4bwIiVbsjDcX75iaKperUvbKCZKDP//NeKS48hyPIGWHRdu0
BfaLgr4JV0IOtkRmgd+E7FwE+uN4spMTnBVNAP7JtCJG7BxfJOjqilvJFHvXQnAH
yEwjpVb45g5nL1yIU/U7QKSZhEps8KsaQ1IVtPHQTd5/h2G9DTw9iuFwaLc3yzJp
dJyBTUjNdKtdt81Akck73+Ut4ueTsCuBIGGqu8rb8yggqVhLn0KklLdNKTgZ6zKq
6B8kaq9rAFL315HYO2mPYrJJ/SFgqBdl5RZVqj47hcTbTT/eAbKD3tWUd9QOMmM6
zNuFyeU1FOOk8cY4glrkgA==
`protect END_PROTECTED
