`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUZYtLtLfRFkUTs18DgLrgyPaQ70BeVSiKks4hDTwmRb2N9J2EoKTKVeaAWtBDTk
rPRXJLb07r4DKo6Qecyt3249ama/X2GjAKzRAv7yLdvMYmSa4uAgo37eD3YGF4GG
kwlmBU97roYusK/dtSyP4cxkW2MHACdlfZo8e+E9RyuyUzN2ci5YPq3QZoOD+hkx
UhseI2L5Dw4PuzfgZ88nHAz+dUxi4fa/g5guOxogqgClYDAlftUP6KI/TcNZg+Df
j7eqoRCQ6rUBT57da9LRkFuvp6ICunJyU0z/mhTihoGzw1Dov8+r1kl08FZ3As9V
FeW49PLqXDOJIEGcfbgWmNc0YLw7DeQPHHEwvfbahBQqsdyjq5Tw2xMOR0tMFL07
3giB3c3oD9AFXi0ai52C2kGHnIs2hv2GEi//C7GoU90=
`protect END_PROTECTED
