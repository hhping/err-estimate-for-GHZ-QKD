`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpsQDrstQzqj/N3AP8uqaflpKmeUPmylJuDhmfutUCrvB6lrfUguaEEYmSq8PgX6
vCcmQ0pmVmOR7Z8RulAxZr9yGH5kUxWEzB9WNZVdGwSE+7OkzI1cQv6m1v5beK/t
1b4FbpWpWzfCokNXzg7gApRRCH+elUKQl6Xc3mx3wNi+Z7vHGRM6uO+lhwMA1thu
9ABJgAY3utXoNy20RWbjtK0oZ4JlqvEjHiH+YL5PUzBOkCZw2wPpTzN37SjucbMg
VXU/yT7IeeRoRFUfHJ4czuUT20z1cL5tmZYKyt3k9a0AdkGdZx/HGnFTLY8CLeJG
iD5hZLP+THNhyGYkcS5Iygsre/pydKMFZnPoykNkVZjbEdzRpL+1pwahe7JvCKyY
YRfdq+rC8HSxz3tzYk1xF4z0w7EkuwmdUbM7MI+ka1/T3AVDu5byd+6Ulqu80S0G
Ih5flHA5sJnbUWGhmLHw5JUgCe+isJuuIms1GxM8azND0tBIpYfNsMRezOfBcwto
wslSiePOagmHrggAYcelXaHhr4ko+WV60xsfxj0Zy2guxuFDa6cOWz//hl4HKe07
gLQoAhz57aOga0n1pqynMDS45hINaFNZPeWuULgt95Mf4z585KEIPOLK7znynnBE
E9ZkLW2KCITAknui77R92D7MG4wqIl1QJuBnU95iRPhIH2fGS/fAFjMIWPYVBJED
vT8s7NwO8ASYne+RUzfCtyskOz8auHImZyWE0DOShWNjjxqRGa20lLefaDcYNJWg
`protect END_PROTECTED
