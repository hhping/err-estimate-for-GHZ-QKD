`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vm8g/G3G2/buO9XeAIwLBvkuWphmzk0TeDekXBDgBbYKFoQTscqnOldJVJxPeQH1
Y7PxK4nNOvF63QxpU0/61FU8TqkW1oM9Qr7HvSFs97QBYMEIkrh3SxKZfFKZ8B/6
++Z5zp+MNca6x1EzBL6eHHvKgRCI4rjy2VyIWR4OLCQSCaG5Gsp+0sV12xUZn+Hv
xEbvbXEjbDzHwzCkc3Wmfj2OueXLE3Za3cKe597NQiC1Y3sd923jOAiFyLFtQlaT
D7vw0F0/Ufw0vTowrvv+tPri1EvMlUfjfO9rTYCMCNAAnLOSJMQ2LeQIQT9i30sf
abcKTjw5K9LDT+xMykgjk923PXqI4qnTweKxaog9PGgsDRrDbYZqn/ndHFuV5IBn
+JmLvOG/6rFV++hhJ4hwv6k2Wjgg0BS97T0kD33sTKsZ1WzJ/v4SyQFZf+RidlKY
S3MbnUqjUuqCjmqXp2E0nm5asQV0IChqwtWoeP0NZ45p0GL2F/jXF3tfIJh64rNO
RmTLFiZebVFYsEuBbgZavTjDILD6sLD0VKKMAy6TAi7YIJO+JnkMV32BFDo3/A/Y
ecHXN3/1fE5oAcUlyjGqFaZOY2Tw3Y7nTiELwFsSJzS5ssHWaxpaCZTj25tSWwAV
CHMRtWCuzpYDmTp7JVRTYJRfZn/mSKElKZu1yGUQFU7YS4f2r0DajHA8J/l/Hdf3
z7CB8fWUQXj2b0u4R7oBGRbtoUOIMMt0SI09oaRvVhOszj/rMni3611apOOwFjZH
xQ9k4tcOxKwfJ9iDtSzlAnCUorcyivsr864qInJ5hya7qcIFKtXjv/7mdgRmqJNq
LGnxSiuz6KMIbrJcSNUefgniYUIWBdLkLUIkwJZCp1zxGpgbHjLnW584oEHUuOae
J8QJ3apTzJG79+LP3NZOkQ7wyChUZa1kavHG4G1prf2fVLbtlF45zZXarBWwg4s7
dgeYC5eQ6ZItOMyQGU59ktrK4JatBVtJb1rxo0v+afl7NTy6pGQXaf2emmaSzmme
rH2WfwTdpk6HzdjqI5nHLU7jF8u7Zvjvhr0zVFDQVaezxq+8vZ7whRLJOL9PCJll
NbAk7yactNWzrxiK359cdI80gVzL5YbPtCUIreTf+mDBW9UBw6OONX+Omy1Mwu7p
TXgcLNpNSH9mmhaTD1LcrwVIbHaaWHbCCtsVDg1suW13xsppRSLeX7Lf3wwNWTQ6
2Gbphl0xwhVyeTBlXcOydJJ7Z9ZpooirwetEQsHGDVHpvZTuHrc5TTIVvbFJTJqT
hF9RHa2OHofQ+rAbVZ8Kh2Y68OtsXiEIos1cGh8xFfA=
`protect END_PROTECTED
