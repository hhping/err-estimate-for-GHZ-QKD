`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e39QFBEhLtY3HtIRGwqpVkYZ/aQtzEKesXUkL2UN6hCY7Zrx2cQey2tMYu7jypRW
g4xj9DogriDmyr7cFPN7wat9ZQvhayhi4AwXG75reaLi7cRenu7E2h6JlrItrZk7
ifm/EgWfm2nW/EDCYGwowyxGqCOmGYmxxKR9tgk4mFkPVMh310Br5Tx/bxYMk4Ps
g/7oeEkvbw2Qh7BBlOK9wYLL/fRkG1R3mUqlHOHsbVH7+RtS6w1ngiM7k7x6pI1e
OroI9q43hbyuFYxrZ2wjUMi2Glx+3/Xg1xmegJ3fhY0wsZp45loxBAbWFr0ssrR0
RZm7fOvuBLZe/3G0G8LVAhYSl2+bc0a8Tro5dbTxiqhpevv+WDIFAr+3FNXr0ogi
ZsRDdUiOqRL53FfMervG0UJzzojM+JOSpleXTtkScoNrCGjczaYijwbj2DRaRceD
eEoKWtG0e6dkFgiSbFo20PKBwVcLxFPvCqWPLp2GLB91mis0j7bKS6EKkMKCiQdR
3trmj35AbcMSX78SSuXUaPMVAbiCfXX0Vex6HAZwNtXMPbM+SbTpH4ly077S2g5n
`protect END_PROTECTED
