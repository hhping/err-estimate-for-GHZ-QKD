`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e2soyeR9MqSJh56mc8zbFd/Ulrv5lzn1WvOvEFVu4G5IaHMm8kAcIu43it1DqSxH
VJBXv7wk8fo0ACN1JJg9/i+WozWATsu0YIfWp2SSLClgOloZes5BKNr5+8K1di27
qHTIcHRwxu/j8aMRbpFpdz25hieZGfSW4RgIIpyA1P/jRc0phaU7LraWRp5GHxrD
KyTmVPmyddyaaZB/1v0oXP3LK90/apaP4XGhdVdoZNrAwlCE21rJOx43L9lChk8y
TgknvEpRn8SBf6mK1h0DepZoY91Xm+ER7m/IAypRT7vX2rayfqvXvOJXciZb6OBv
CX9fTPGHJzUZFw7Hb/Wz36ztS77oSvZ/hEdmtD9wlaiT1npVDENI1aZdWG1AgSKs
R9v3d98nbO+cGJEwlQdjaXFJb1XXunrm3tzvyVafZZ1+ygwlDXue2IBJkwYROWXH
HMY5Tc8UCjYD6l+Jwyc6oZO4axmk7TFNNBa5LdZqEruTenufcF2DRy2eUlbbC2yF
qXsJ3M8XfPPhAvm+U0F5nSHosLvGe3ErvAFLidkylQvZlrSRoEwAsIJHlQA05nqe
8Cro1uNTdaQ2BVhuKuPBUUcuWyxYpPp2NFF3eWAGIPJzjER6+qhJ2YUvyXhuW15Q
0gY73mq1oWJwKE4BeZatrlqPb/CFpIL6NjnyRZDDdRgI054fEM2OpBLwqs50ZYJO
htAx//T+XUSTjR+6FuV3fnSWAstZrOOd5LW4f9Ol/Rk4+nCwfWlFY3JcPsD8PpfA
8CEjI4vLcqQR1EwrTn5EAAI9xevnh8xE5VuLA/QmFQb44o6rtnf16RIWx51OmvKY
GP2LqX+ezklMhsqkRZAmLjptyvILP4fqZxc/x0W0vO+KJc4f1CZPrk/oBnB8ko0v
DEFAGfuPJFAjNiq8A1L9sWTun94ms82GUO48zVKAWY61y4MaFg5Pjx2diuaThFIV
DImVFq+6rm5fjQz9pXAMaEallJ4zrt/SikPFfs9M0MI6OwY/OnKWCG88iYykwMSp
zqWEuxez/wpX5fcIy0gj3snwHjCRYUWFk+G7InacUmcdqZ1aXvlMnmoU84C93S2a
iug1TrzklxcyxathXXeksQjCKZlYHYUO1jRyynuUvrD7M82zSv2go4qGpzhE3OZG
Z71NJ6kSbGRRhnrUBpJaIisN1wR43k7gwjloZyOXuXHQ0xaY9eB2pNbe1vbTMFEy
oZCnnOFwLIiDKhHGWMS3pxbn9nTT501tE92zz+WKkIEWv2905yXYWERANQC1QWqq
o7t2FOjGsRsiNPY/D75xdb502uO3OJX14gC8++5LrIFSk/ZLIA8eXQb1/7oVzPhn
txaZrf+MDwNyrQ2fxdTnIVeKOI/hGuFPMmD6nSVPjz4w3oVZDrHnJSN9cXP04Mmk
sBhEY9PoMLDFvE8RGY49qbDHg2jy9flzzUTBJhtLhmOP1XhouhErRpdjGylfXTRG
jaBkXE7quA1VWuzGb9R6bPDTA/cxSD0krhgJAaRt0jR9h+YKMH8Pwh/xJjOW32VC
Ps29KyMsShDxQrWVxTMc+uwSDICqchp7alJ5v5kKxg3Kfpg5UKyPcVRrsrIptw/D
PMcwfhrUsfibrW02ZdU547jOg6OzLd43kDTys1197+e+bZA5uXwYbSI7xwwaj4Hu
Ew1xVmLomArW/Jnj1tx1+fCk38IM72or02UzEmcWf7ZDh9f9kxBQQisM1zeQbyh6
ctgBvs6MF7Fsa1PJLtVtxOKU79xo8TZPCL2mnUlmj02JNK0w6juxnP0qA7dstoSO
pkpTAc+oKOGha8YgHVhcAvRjcK5ElS40KMc0mO0rKNApPdCuykw01uhdfasa24Fe
2hmSbqXkIFBUArYV51dCOedg4emSdkGSJGw2EmVz2/yUDYf2eVby9gTLl1zVS9Wb
9srH+AvGLXmCBsKv/WLceY1DbWJwI5t48+0LFGrUCcurN5Gyg/vS8zpB5U5c9wk0
7x3TrCRP3yHi8GcWWnuaARTbkmIXenLW4S6nWrYtTKH7QATTCbnKMDDAGaEccTYv
LmE/JYQGJae0sHLa6LYCtMcUNKSfBFD+3H5DUwG7QJuSdvpioSwrvPW2f1ydP7t/
MdTir14dNC6WcPZwqF02gJTwAwNfvY+m05ZkYZG3fH3gcSZ+GyJTK0Kyy38nAcoj
151wcqJ7zDRYfzL7MIdjLeWZK3HMsimHwkxHL+5zUa09WZn6eE3QW6tJByNH0aM+
NSyd1QA1/bVPNVmL/jTDiyM9SDEkeQcXM/bhpDjEcCj08gs8xaF4STQKWklUTN6a
ZxdmYQEbw1S+RdkusU/qOKM3PCtrAHmNUB21zYyMOPfuAti6PPoJo6WU23t2e/N2
cjHy106fUtWZRw92TRlFX3zrPP/B7IHnm/Jo7DKIk5EpDqhYA0agPeEpH281S/zP
m1/GK12mqz8Q8eDfwJjGXLlYDWOA8Zopl4ML+xS6A5WlRj2vS6XzCPL+y3AIZwcV
FL4WgGWA6x/KzhCTO1u4zK1JfnJHVbNpDQc15qvWRBk80rGHay7NjJJI9w0m/O6k
sq5IH+vf9mpCNCOdZ3iiXsJXGuoeOOQkirYvrp+MWTwYGXd5z4yf3J0kD+3ieriV
3wOBBQpKq/rbnz3h0Uv5bZ0eDrDTa5DDY5hOcOWyfh01NEbyAM0v+4wXMBfvl5GV
m2+c0f4RLFYDgvimnYwg4NvbKtwAiaHSTikwH6qZK5yt3vLtRcoeSZgk4C+uGAtu
Gn4RDTQ/deySKzqPQ5Z9kDzegx4WgT+yUyu2ocMjC9w2Yp4OJsuSOFKMl0gkiTOV
U96zFUMZi+KLJbrhl2kVoJxvF0g7BZYQBuUq7z3Hp7/vt/JoN0wUgPE/IaQpYoeP
HyPEFj1NQlk/m63xOCpWesbhlc6eE8ZZhuI2H2FDmuAeA7SSTFQ33zh8N2SdwABZ
78zcAFqrDxCVh83kWQv2BXBxVbin/uF8GhCl00dzEEa6UyzB+D3o2JFGC3l7B28x
3lqAvzlFmfp400Fot6k9qKLMex96q5NKEARF7FsqrpQrT8Co/OZIu634s14uesil
BULKxPlcdVbkSHFn+nxGthD5CG5GeoNcLcaUsrtLbAWRE3NsohDrBAjT3VN3Ug4y
gxJ1/LDinwqGSW3vcVTLRGTQHmaW/+QJYvtINpV8IVFkc/fNgBhQ32Zfso4+S4wM
LoJukLnUHRptq8sCz90Y9R/KGYKRYiQSKiMDqOz0oKC/OsTB/JeAdQ1scmdrhKP0
2lsdLnepOOyXS8mfD10bJd7x8clY+lDYgIJ5Lm522ri88PIE5yXqTBjouYPF1gnl
lbrvJM5rCEucujFMKXWN1lcCNYPX20q0uoyouXVCvoZUiM8ROZ2rzTPIQlBwosLp
mmLK5gnMhHz/gbs2EMLmYRpZcNQJ7rsjtNUYP+8IdzCerGfvtuRumZ6NERIEKPk8
nr44ESr7jyilkFPzMT+zLto6mmqP8cKywHpLsHKEO9s=
`protect END_PROTECTED
