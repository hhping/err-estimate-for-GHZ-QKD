`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beQf2t6D60YachZX3Qw3+mJD+1ZA1Vfub9hkI1BuKqfiXorxvToV/TcOzHe8hBmu
kOqWm6wT+6RVuklOvc3ga6GGrdor0W/kMwMZjcFj3nZWcPhrDX8l8WtS9dDDFvIW
NI9GOjxoj5IaWfey7DFQRgh6KpFivSXG+t6xobkyZlqApq3tjPRhwMtbGFeBZjVx
mVEgwC+NI2FHHITBDveFn4aTxsaScqiT8Z35kaByqtyZnyNVJAZBPyJeftf15bnw
xGUwGSPbZjZoLjMfwZi6oJfGFdvKy0wUA2/uWsPblIwYVrelA2VRI6118ZFdLNmY
gYbbRC/zOiEjW46LHU2MCwEL8ZXWFBO/Y7OnBFqpbV0Pb/GxW0QnXge2ec/MgkNK
PLzf0m+3TAycQQ0LOo24zDsjq3jszEfDbMaJxsTPK92FLb0KihLuocEZvNxpdkKk
Bi0Q1OgFNWxKdXDTt/q7/YVdYTDV7+TeWhZYJT37XIKbxI56CU1BrzU+j1dQlhiy
erJzAx9ZmIXDzIzdgBXmVGIgmWXycooySyviqt1/TOF16Ro/PPFAzcSISpJWuyH3
bLfw5P4VSqnTiw6FiDMavNzYbmOqB5MP+vLEUO+ftR/bNZyqHQY+ySEYcE6RvZ8O
G7f4NeDv/nV2k+Fuj80LE/l6JgFQtE1TnPMefXAkSyt3uNUdnUms4S9Oz3nOlLMn
S1ghytBKreOJn3rd1on/DJEvQR3Ip/3U9gUczHOA5KQ8e3532kOVDhHyOpX2DW27
etkM0bdxhwOF2120myQFpC4tb+IWnkSUwrZlxmWoegzSBHck6PsiQHpa29gOoap6
+kakLvIQf5lkhLdLVJB44B3vGMMsLEt+6zAdkxJODZ91VXh4MAlzH3/FilXYjKuo
33vn2onydJujecrJTWVBnzemT2x4JHIOXdyu41LuM4mfsOGFqoNvWP0aKRJyFaNO
GyoTqa5QUbjy7y3nA+3t/vkg3dnbtbrd1w8WEDQFbripZmlP7NoRbuKcBa6x5bOc
2+PUWsVD4lqG/tL5QWYOlCFoelUdNWpG33Tv3ouhiQeDcweYnFePQXbkMtzG+mlL
aI2u/k9apg2VKCspVh9U4d4GcXQq0304J/55Jpn6UmpCVjj0Q2x2q5pHi1Sxt9Vg
ZXpmeiDJOPHFMWNoCKXnJdVCs8JlQ/5h9SnVs9ZXMYGU023KubR17h/Jvrt/HBU5
bUjCXXqKmsN2pwASiqTh+rcvPaUe0RCXHzO6ZVhv0VWI/JHnsJhzd1zGaRdBKVbT
ROVyeiljpOLiGGKA8+EOrHd984ngVbNTbBUuLVBl8H/vPBlRpS8bHBo06/Pa6GU5
J0FKA4p8zEJC+IXiSlETs2CY7HpfP7YcPhIbf6E8bvWlD8N/+CAjuprcd2Mi0RGf
432PMfSoQ0x722sUqR/VCF6A1IAixFhtjTK1hJnYYyNYJeonU/txxTJVCnWz7SiN
6+F5D374zqHXMpN2irbz0JZ/dsfcaSrl1vZoYkiGU9AAwSoXFFfIydDy6YtRzmQw
Rsc6NgmQkLa/CiuLlESkHHR4uCyknyhH9r/7o7MxZf45ux5mGnkiopvQBYnyevsg
qJYpeVPcRq8ysxsXelQyZ17wj34Mbez47XATRA48GDRKC/dpUGky5vTic8MiSLMV
Pq+mMAHk3BT/o2AgzyVkEDu/kv4ats2gfqu5mWHH0rcf0cbkyiDeJOSNPjD9Ks1Y
K3iQBBA5/R0h+/XER5MLrClWO6oZb17NBoh7ecenuVRNkv0PH65HJgVVbhRUx/Tj
6Uxoo0Q+QQiWQU7AElynGuauO0vg/FOl4s6H2gFoKcygT1lXuyYdyDXSWzv5X8+R
LD6f8Ld+qc0Ab3MBt100/o20ry4oiBa7eJRt0OfGO59KjWR9PPHsrBS0oXN2l07/
AURi93jeqAf0XMqqnRVy78kseMexo6XCJeskbYtYIXQrZ1ian9+pCJaT4El5Vhao
L3dzdfeAhQER3JWqLShPc+EPTeZc0kDJ5rUxU5nhy3PVh20g3PkGIrTOIi8TOS46
+YzB77w9bewwCrQ1lNXXxBJd0OD97AODMQ49muyX8PchD5tcNHG/2JKnVnpOtOGJ
HGs2ejgUIwgLpe1W+q9kimZxjHeUMOBar67wQXr90U7wnKRt7xOUDqAL2blfe4fU
XNb2X23j2ysJXGdxUUSbRN2YqQNDz6AicYSRlvW9EQbpT+IuGTIAPr53VSt7W9Ny
jabp4yMx35agfFxmdNno6oGmSYckWSKDfjJi9MLOOdZFJY3IEPSdLdM7QpmZNhdX
JelTc7SpiHT9cgd9B4XsuHgwecZEViHZw7e31wckQ5rbl4CPiuZpomrVOxmBoQbI
A4XOnCN7hgk0uHni+oQ0QM1Du3pSkXqq5cLwK0A9z+t+00TKhAEMNglhH2oUshMf
wZYVLZmIgz8Zb++thtAcfVFlKt7aztYaBwc+5o4Huk0yCniN8qFBwXcsTMbYO2uQ
W57hETu6U5tM4WCvKgB3GA==
`protect END_PROTECTED
