`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3026mUo7GucKm8TjqtpARV3JUL3ZWPH7zwTPD0AgFSRU117A2mSanX/iqq5tFEZ
iqAT4eTRXulUP5vT1G8zgki2QaZfwTwhPFWkNR3C4Tse9rL/Rn8mBZeLhsbTmIuB
DIFKqFKV6eWIRuxa/4fMP6EVu/O4QEbGDVU09HRkY/2EYN/4CLJCJOhjsF4ak0PT
5EQ82e0AR8KViVeWVx4hXMn/DNFMI6kcW9zILSJ/E70AmAbfjQTRZAxyGFZIY12t
O05VaPuiNvria/pv44oUeCRzswuDxJSn/UXgEbvgzdO5HdP7TXe8UdNQVzUyH9Mu
0nECYsO7EaIs8ZVboNOoK3c2oKxNEDee8+xEzm4AR8+p+yVZUSL5opTNwsqoCHI3
cwuS7Wx9q++zqM3KxeGxrKHjxEc8w+ZHv0cSYXvWMl1GGXBxpUAGzUDUhGRpPfPS
RKwHEndCvCOCWVZTXjqErCLg4TKVsWnzWQj8Nsiov5ItBpYegY6io34NbtDNG7Op
GYNo7Xgv7M2FtwEEcg1rrqhoGthCVrSekkRuyMyFP6ZbWU42UD7TgR9j0qn9mEdc
GeARyuSZ8a5A3mk3TnAePeyh2zvbZagJl8UqhKVNPGQx2adiyYrFF6ZV7xaP34oU
Yg1AJm3HYJYF28ROpQTJjOZvHIGAk0KX07if33PK9BjMgc5MQis41QGLgz3sdkel
0qnTzmQqJz/58KJM3XvHCPLKjyMEvjcga/xM1JiVu19vQ4M9OZOXv6u7erSIxYV6
ZXnt+Vsr/H7BAPsRSx+gXZUkZmpqXcofzKm5owgwMG23bSEn4F3yt4gkwwxBE4RW
6LHPclhly2tpYZ0lL3qGEWrbuYmB4Te0IG2PbEBpPzlspz4eO/Ca+cINfDal3qdQ
7sUmSTWowXpI0SZ8khqGWFFDk1IacePUyB8i8c8mpfk4YG7ZKQ9qY038R3mmd7oY
0izan1Dq93IB3S2cy3G23g2agvDKbgV4JKbPBY0H7XCIJumI3Usl+Wm7fz7vuQfg
aW7CAzz2OgylSXISlHFT8LYriGwgivb6ENA3v3Yz43gpCgNup+mTNXv41zHn6pW2
sh/1ibFCoGXKnUqYk+6q3rIHo5evlcvLL2thpnOmQarg/DM6I3tEWyg5wYuZr2Fc
`protect END_PROTECTED
