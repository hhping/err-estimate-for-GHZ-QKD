`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBVQW5AZpOrl3Un1dx0PR7tqkbeK6pcd9HE3AGiN1fB+6pa96j/yx0VRQwQWvLa0
aGP1e54XP+fojv0NWQ70yoVWckXy8Z95zbyxyucAoKhseWiwQIvte6bPGq1isPTb
YA/6w1pKxf4OQEE8KdyK6MwQSn6wVu4Jn2JKUg7NykP81h1FS2RjMzhkP8mlDZwX
D+5HU7i2p3bSc80rfh1+962rzYY0PsmmJnvX/ZVcpRGEJJT9HYkiYE0wG6F7EdZ5
irI2YPz/hO4BHLVJaVpjr0tG0O9WdzhGsMEU3X0PIunegVW+r8pPA1hqQTI/lZLH
BzPTvIJuTLBEjl2EsBnuxRGdPsMK8bBFzSdzDrH2UQxMP8ojasLZSBv/YgG3bnxN
+yFy4gK/9jckQsmNKObI9tc42U98rtTjZY2o/0II5uJ1oz0TYKvQEILvpPgmNAbv
2TmcrJxRfhyCHdfMlWng4kKcwLjKTkZrA1OKJ4TS2X1P6FD014jPUdeHtIPcOssA
Tj0MSTy7KBYmLshFPAgtLYPtRNLwtrePJMwJRt7wNqxYUwSpYiyY+zYFDsLPxd7s
/il5Y2eJFGniy+GrKCBbR+yeR1l89fEY5K4gIhXL/8pQ16WJ8zqX6kWlpFk440jv
ppz01X+6Q3lAM29XeSV0rZXUVUCg7UXCdDXRUlxAgFIWT3fslAk0wbp9ynVVReEa
RRyKdwiSerHnFTgAxVG5XQc8ywqh4IZNVf1eMbIMAE3D45L8BIRqCQ4u2Bx37MVz
zZq9XipfNV6rCKoGcl1pJGRejxxhpYk42wtxE0QgSZKhlg3jpOkdt0YrT9/p/Hcm
NIRXH1y3QSUu854QgHoPGIzXGKozmSQrpAp8IH2qEbDoqw1JQRhJUzPGwitaX05Q
ZJKTwCCJp1rHKX5kuXtRthM1fPa1h7vNHr5MuPu+bkX1R7S2fvKlwowFRorTYnDH
HuIPXxWmHP/UVmDVYcCnVkT+DCT4gqsbgG/7R20eILPAuhhpQPaivyD8T/gQHaVC
l92+SHVVJQig1vKHXmYYPo+uixgdJt60ygxrZ42IMg6ZDz7P+TNtNjfNrbB3eXz9
diWRwg93nX+/WJsbncD4Eg9MQE/cvsDuYuyfFCCCBMyLYG4mfyWuTs+nXF2KZ0ea
J900P/tIM+4wLMDHeYqBKLKNE9qOVjb5Gzwe9kvH3TEnwo1OJxz0iAoAUaMfnJgr
6Si+PP5Hupvm2euHuuQJ8OZMTrkxUCm7rxTOmrSn+wbqd8E6xXxUlLn0+sO6pARi
k0BSLNoCqxOJZeNVyTKhl4eELShqNdTMARzktScSrNX3LFJqeLFXoVYMCGzgSAvk
YJEaogn5Qk83E999CAyfSsgL1YpHFdKcLrHQXTuLSfpX8X57JwMxMf/GUL6da0/a
0smOvGh0crSjpX6WLMUUcD2aD/6tjw2g7rsOjK1wkmwLyOSNnKgWPbqL4j4zTyfF
Tmalgg4nPeczVGMfOwaXRO+Lf6P99p8JMjWomurpbZCneRXF62N3Bs9dNHViUwNy
E5NZ38Ewlwcjtz5vD4mYZOSqXAUuUtjkIz/w1G5Kt87zpwmYXItPsPJu/X3wLtZZ
`protect END_PROTECTED
