`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9P3+HQoDoQidx09QPRpIMaDoGh1yviYLHQP7lPjaKhSdHS8bkSJ32rwlPS0D9ONC
M24yUwI3bOfICX3LxPtE+weqWGoCNxcRav0gBzvVITla0qdnr7UUzaJVTKx7zVjG
ygmKTa6L0KMfDXmFL/XN7G85Q4CDGz69ZSjjME4N4T/YAgD2gRDAuax/yngGHRv0
gr9QAspjXwUuWxyTCc+MfjYUB5jUQt1r8nudOivSdQETtUhm2ixw0DgdsO1Y60C0
na4ZueAvOMFlZh/oGEHo1dHrg848dgwYuyOnplO5o7vOOCV2DqPqwnlkHDglV7DR
/lFf1+7hYAVBoYX1is49HlbUu1rRPCMkeWKegH2GdBMgaWK2vf5RAeyoDJPqpNy5
3R9sME3iqCSUz+4w77YCF+TUlTfvKBnV6rJ9BYFfSve7EbHVRQRWANlNLdyb6hJp
V+DzsKK0tECZpf99xWWyqb6Y6hYj94k1H8AZRkBoLJp9KODbJEei963LB/6+9hGh
MiYsJrjRbgCgC+w7K8MGXKmjoPyRHwR8tNAoqtMGBIJ6NuNJ2UNn5lzp3Trrdelw
Gb8M77/z+/nDAO6nU9VJwzFEwFb7TSb8/gd2h6bzPHzMED9OEQX78vPcAVctRBm8
hlBHvxmOV2P+mLiQLdZosJ/dZ8o27cZAt2KKvfh1znk+BIh6v4tkVj1cInLZt+GB
s3FgUEQvmgu0Ch9oGLy6cHr278MZve6TOuELhw8l/OPVlJdolds1Ksl90xq9VnF1
LdI/rtD9M0aLr97p8tPURGsPB8dYQwd6QwnaVtkyelwe2ms30OsxNQP4005M7Y4M
xAaqEiRo9pwiLUnjt0/1vLyvXdbqzCdrgDha2wVVIRPZnq1BUSd3PJY2eCa+eKdb
QInmCNkum56YZciB4RQehyXwHg62ab8/9RDJOQNhgQIxzHRS6TzU5riTS7ketR9/
piZXjV9+O0IVwjqWD88h20INZ83QtYrlSNG1PsXPi3wfU9RjwnEDKspYtTl7FtUG
V+4KjdN0/F00oMg4PJ17mjXLgFBjSwkzW2jwEj/G9qbSFqrqUX3Z1HMp7M6wVJhO
y7WF5JGVlRnEMIFjaPKU6i2yRszCAQx7wHIc19tCN4mddp9p6NWfkv4PCvq/tx7x
nhu0i6ayqT6fK7sQkpi0BD/bxwo9DopJXgtgn5vBRlXbwkVTiLYBpnanSDQJXQg9
jbT8Y50Eb8tK7Hbl79V5dysHYaHErtjtsnMYZQrNtjz5F969+Ql9ycFCAKNnTgKp
Kzh5xW8Tg+MK2WG24J3SzFlDXfJgK/k09IjA6qTD6eugwggo0jxbD4pGbrmHXTKr
YAoqQsMMsMLupT6V4YFuFcE4y2+rL55vY0qDeG773qoWBJ5q2U1ukKde7xJuJrSP
i9fwhM6kMLIrMWTMnoWx0eP+qc4gpL+FrPox/4R983BQyYZCUkVPM8Bvuhftl30B
mD48x6+5mSTlsVpH+xvZoAjwhnkk8JTd0wokDIvPQouQh8D+OAY0D9+iDGO6K2GT
UwwzM3hWh9AT1QCCinKjKLud3o84SlFzfcGWq/oKPRG6Y41v5rLAKJCv6q1jkeTL
IGx92KOvErX2C8FatSwPXJaOdPDXMH37OS0CTVwekSyeStiD/DGo5LzEJdptTxRf
xkRDjQA9R8K4HJUu5gI5JnlPQL7UAH0QRg09BP75yX2TK9+rdw5iTg5lI118Ew6n
RUaGP6LSQyms0SQyUvxfOcl1X//FsCUeHTVjONm/kHBM8dB9iksUgR6W2rrpz8YX
DHYQelmamG9eW6mduKROBN8D7l6rnRKVezLPEVlBXXV3xHcrGbXRvJjZ6N/Terw4
y/cm+ayo7RRgibTWrONKSotLcBT6na/uRdPH4veZM3r4BSvhiJ07cHym9skFmh8G
4fjyo9CqYEZ2hqOUMZmbmWKhH/XI0RgtfCF7knjJ/Fe22cKelscaDaZzWnZ4yyoS
uZwwYxOKFAO0OMP/88K8/mhtm6o6yC/XMzMQCNYGgICOqtvZ29ccyuCs83xNZR+Y
ePQHGTOphrZXq7jnE/3oioy51nHUmQDNJ8HwyF2N8eTvtkYdeE9HBXhZZTpgmrbf
iVHVSf/cYd1yqs8/brrEXs/Ca+tWSTStwN0hFxkKSONniQ2bbFqAHoBAHJrnn7Nh
6+x5l7dDPv+4e3J99GQTsePfCONlpTWbk5cj9SBcz6CL3GlXww0LTVUiR1WfGOnE
529PlTCmESvIUK6W0DyMV2wviFDeYu2HfqCQs9cK66HUGfNAiSXuVuHGHIKZiz9s
4EbkUOpc1EDPCz7IqaQWmgHWllF5ojBNN5nrJs/RKV8z8clHeDeP0pW+oJaFGe2f
lRmTRpBMnpQmSbJmixk6OoIwku91cjUqUfxsSEkkf4JGSri0/nRnSqL6dgTUlSPg
l1hgJ+knZnFxrMDB+Ojp8AS70GTJJ2YjMDFW4jG1esuBYuBeg+dnexTyu19GA1sH
mF/6/QQn3o0R1pUNMOo204nwr+IZCQMB8wR38e15D/WASbUudpQSeQlnxxgha+27
Rv/To6TpCkV/iNQROX0dzUoigoPpp0oBPjdezjAnpBIcktG+f50oBpFMEfCrqAuE
0KXdDOelJzKuzuhiX80eb6MJw2oe+7mqgqqea8xpnMjjMNRVgEig65t0wJCIZbWR
8Kl6aTcWtONTby72GSQhaySU11KukSCB8WDwMCnEazxxzb3wjWt60HeTlcEsBdB+
O8towaaRNPX1NIuL60OSk/35RtH52Fo6srpU09afBZBVtBoacJnnXLBaJ3enMlOg
/hA5xWHmTaEruTUQr0r6zDqwj2eB3aEEbVAUq4V8IoRvPlQkd+n0to4qhBC8w47s
d34tB/Gu8XW60l0sMBckOQZUVq5KDy9cwCTNIeL17x5kPkmoeiB3emwmAQ6wtzrA
vmjDjwhfMckXbQDzYuibNOzOVWwdjT5wxLc/qndOiumVFMIO1kkDtV55FYRinuxj
Z1QiyWhXB3mVPnGjRovLoxpFQZQCG+c4LkmVIU2AWoI=
`protect END_PROTECTED
