`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vlv2K2WLhyCk6YTecIe64UqpN8XIQGxIaRbGN1Xe+wpf5DUmTQl1rs9qPWjEBtGy
YyDxY+FhnXtXyf3/4SSerdfaQYIE9/823y0wmiO82noGygm2RJT7+mcjveEW8Xv2
ZV2gWjgmrmNBwX0GvG3BP03XGcVW68CF0W/10YJM4SBOBHPfAqJKbzyTxH4PjQZv
TxFq6KgMuG31vENzCqyWp/ifKzqzYs3dteGdf5drVqkiq0sCr5xCVDUQUYSITkoR
OeIKmsDll5yvKfK+nfxUcFEKwxCAb1zwNkH11t+1pOJ1pr7si/RRWfelmCM8gV9H
gjBrsO+ttoZkHQPMrs3LVVIqhCXbAyxgO9yZhqVOAlQSIGpwJ/ZRj4i0X1HZcIYY
cppizUUVd+bSpnQExMZGJP0Q0XdaZe+R6E/aozj2dTmjvbe06/nPQlly9k4LkWaB
n1bxFwn82XT7Qlf+4jV1vMYwWmVwOvb1nSxHEuwPUfr/dkbut8Gr8N7XZUGvCZXb
/RgTsOC29ocrFlZenfk4NuTKWzSbBz3ePlpefVNnBxZeaKzEW+9Lb2UInwsBqSY7
4CE5HzDRNIdps/VB5T8bAr1LnlbdwOSy90Mcf5dbP9WYolynmpbdvhzvswmQeHWs
VSfbyUgGmIiQMSEUPFinV3e1Fre9KnjLWrk7L8u1mK/VvfYwqxBv5FByPzN/qYYt
u41A0gn1NVRXFCd2CkjaBfIIKWl2xAuRR5Yg5U6VlXNsaVbNOaNEYbpODyA4V53q
SMQqi+b1i1mPz26zF3plgHCeEFwqzqn1UcmKcdA7W3cNc5Td45ZnZKtefD+WXyIu
e5uAWQnxhvswS3c/55YVuSZuzTA+bHIYi0gSARgeGb8r7KXLdumfTTrEs22q//xO
K+j9/28vL0x8vy0+HCxoVEImoUv/CcDjJw0PQejz4mT0SnxUV3+DOvLOCT3IHQ21
0ym9Rz/WnU5i8w78FBWG8M31ehFJh++19y3ly9ukt7/1vC8jhUofSZ+sgbA6pkFw
sB576GFTN+Ys8q00dGSL/0UOcqegdudhtlmphgubhCkjGgUv6L0AKlBoKbQR8JT2
LyjTZ3naOH1sh3pycGi7DHFo1Ee0ySQ1PRkQpfDa/6EX+uMOpUSek0CHHoecS5XO
8Eowb8al9EEe8kroZg8WP9gxvk8bKBpTAgXEvZvOQSMmoeHXdKeDV0KHSep4tN9W
iQls/NR5flpWmkxYhtzpnAb7kNcVCoOKMlW5CRZOoVZpOpqJAyE0f4xy4pwfPegg
4jFmTv+zrqvx54O2cG6aTUylyBbZ7A0MWuk4+6KSWHXK6UXEKiYGZFh27NMvEF6R
J+QJZJQHg/2NdKTHn+VdPneTautZN0kMnWtpWvT/pxrB1z322KvmDlGDVh5gRtxW
1szt+/wymtxaoLh9zVWf6/sfjzxYuwFMm6YuFzuJWvCaCWVImpH5fe+3yjSsJO1l
kq1VKt5KuGBK4ehQpiP1FgXnFE2Sw+xGxaNClEipnHatNwLYAIIemSsLH3DEqYE1
8j4K0fikIy73I14V8t7hZA8h6pI9CcPe6ih1RAHf6Iw1/dQNPHg7g3ICixvJlEPz
NAR8f1DTiNinozJBEOHdopiD72a4lBis3Tj8k9gsV3R0297KQkiwCpLPv962wYCz
GQ0xKbvnps33KIPnDTW2SL2hVAuVyiYvmQqJkCBTg27m5xVWWjVJsETXuj9IKxfo
5ZF9K9bf+OKvsLfHWUCyS6SYfDYAALXd9mYkLheZWaoVyWQTtjkyOJfYaGLbMxM+
2O/75P1CsO9ejyYFpHcrxLwOWYJOHeGVWTWnvoWDAft4xqgH+phx8M8mk8YCAwp9
pCYIHAdhoRU7RGtiLZYf3AeThgRwrWKlrF0MTMB7gs9cXI02HwyAzGEGTFHpzEZI
V752kfn3/sd2RiKiRWqIw8G+uZrClxzVchnvTXS4YDLehudDcMU41sfAp5FyYuOt
A1xToePp9VVT2nhhVDQCm/yUdYQqmmaMw4+GHap5PLdCllpXDeTh+87iXZf1QmCk
KWDSemWxEDCpZktwDqglQmobylgg4bAsbwAT2R/bHP5cA5QBL6wWZtCkx5eYvgWH
/+4DymlKpt6OdZ8YyXjtkxoWi1BI0KeNUX9D17u5P6j8mWkKTkZiAoqsqvI4JUJ3
PIpDzwil9JZ6rPQfXiJzK/nATAD+9Vi9uFSVsawYUeFTg3PBXEL06SpAQLVrxnc9
9f+IUqlmPt8z4rZgBVrD9q7SiIU7fL/6IN2cYwzDk/dgWH3Q9XYqM+j2Ddg+3WtY
pCqkz79rhDLxTmYbwkdI6eECj1sJmm+tV5WDKnFPQOIIgUM5FneQB2UuoY4Sotjb
RHj2cTl5rXdntMBUH99p/A8yjDLM4HBkftryzJVLzYClF4P/yMokVIXdL626Zli9
QqmlLFarMw8SA/daFvKYBhvdA8REhgiDXcx8h/7VcTEmfzAlPDYza4pvfWiTDL87
qjDAborIkgNmNTCYv4TM/9Ctbp343uYouQv8/sJ6NnZNfCTmKzZxo1kDQCw1gQI9
WIEYsE4gZh8U5Fv+Mp9smO21JfBaQPVS2tzMzwQvkqYcWx4m5Xxp47ZjWN6hS64c
ZwGYc7u2b4XR7C4FtjOX6vzzRMLdcoqyFDDhXWYx3vN5HZuwpcaerEGKF60eXEPp
SKB6LgwOe3DeAz4y7FhUSpXsLQwENZJv8jDfYIpRmsXMTBDB7DKuuiOaH6B/tHDp
BdJimpoAm1l9mqh6mAueFeVZRvrumCu5Tvmvgb1Bp+1Sztmf4/f/aNC/gZ3mvK+Q
8O0jzodQHJ1Rz1gEG+HFgHI2Yi6A/zyYvauEnDmMcUnJ0zsjmWplz/aS5l4N8Dq6
0kQDmo8SBnr6usnkI5ymZgCvNPIjm0HSB+REqsjpx8yolmnDgnsN6JIxC+iEzOgD
0YcavSoki2CV5T9Np2bZaH45BT8FQrSI7yETAnwiCs/gc36Ehi3mW/jamrtaidnq
rXGKh8CkkUpUzpqeNBIs49/5mdDwtgva34njASO7mDgRsV2dR+cYRpQzqHghhyg3
I1++4JKR7dRFsvUOzFN6Hh13tOq6YgSjhselhBKYMprRRIgM/YWvK1XxP1Tot4uh
+cvqVX7wObUFttSNGfhoJyRX3uur2/ydpmwwHkW7NmYnTDRAf6tSBmVnP2MOA+yZ
cSEz3PcNuYklJ5wlp5HcuD4XYBZtnIPaiX4BPOtzTI98zVedQoV0WntIBglBBDoa
XqsZMCdEr+5QJPAlX8oF/FStpjqwhD2pN3U5YDIyRkuS1iQXXpYA92OKsiRjzeCU
FH19WWy8b23kd+OtJ7iBJhnZQgSc6dQ14wgOJLWVOeSwh2az1Ll2hs+TCQckgsM3
W/YtM+WkllXGypZ2DBVDvyQXERBXPjFNe2EqXGF65o4fv8wvmrkpm+7J94uB0bYu
6avUxKwu1V9rMF+QWBmhvguyTVxI/iMVt0arg8+GzSE1K3owufKzs657VyhQWuJ0
Chvl8svcIGkJnV0DJGRjKGO7UcI+CeEG68cFdGw4Gx8hmcpOm7p9kfY9kc7cmUJa
3YmvJJgiNhtMhsc9nzuVqul1sLmMl/jPUEwWUSrWb0cosFBoAtstZ2eHDFLooa3V
Iv6edl16rA0dJE+t5hJx8RArrux1m5b6HPhK7NcxmtGmC4jk53SorwyznpnrfLWS
Xad8WbI8OfYkhXchXQQIMnNZ7xDidJNVzrXzx6BZUiGj3g+dbTyR1lpp4WlW4uX6
YVqgII6Di6NwBqmmkoup8l1dnoIMOPr13Vd2Tff1Vhg4X/dojviDNKj4jIn6mHw0
Pi7vnHR/bCMVQns/c1DCQE01wjivlPxXQlwUYrsMp7ncK9jbJ6aqtFQGAKGNKIz9
DjjiiFnP21OMariAB5okvHTeMpIpTS3GfvVnaoOuzlKdsl1chN4vKUEXydwoiQ39
fw58xwQFyNvy5UYjs+9SsIYsNiB0ms6aS0omNwErkC/sZqsdmqOzNBZ4aqahzNwe
hWY/YG6qvTYT175V85NNQEiAlYC9dJh6Dnc8A6jZcJ9wVaeUe2w8E5fxhB1Xu2nW
i+QMbGsvWeqgXFUl2E1siX61YjZ/Ttq+DX1YOlMg67suEiitU+b2ui97uHn725dP
dCGcd8narrwK2gxAEMv20/k3OvLAXbwHhPTZSEQknYPZOvmHAVX/TEAsD7zDw4QZ
AYzNc2PPdslTuoTTo13K/RyuwNAbCOYIjFcPaD1hfKWNytZ6ZqtwF3oMN5Y5bgc0
APoUH6J6w5bso59b/cjkDFUhQgOaSRyTNZA27m/9+5aVCLfu/lKJK3Ul3H1/fy5q
RUBzQYJKBlwyKAdGa1pyzoHcx9B5X4fjFGzf4c0tmek4LigtR9+B+iWAWZiCofXL
njEzPMgbbUYAeYUx9yNjDsXNVhjrcSahC4qOOKZ/EhSh9XSh94+WMXxeq0Ugwi44
yjmDqQfMctbCo4pCKz2qsrQVKGeiDJfZCesefrymccDSVIaRNZh2Dyq6/8oopAfN
htt38ZxfFXf+eLZfSoWTUeMO/4FdRRNeqzixnp57ludeYI8mEPzO60KCA/6V2ia7
/qnRtbD7NLf5EuB5m3CcWi8AHrtsxwe6e8kSwHSqh8gZmxAfKL7231oNtrs2cYDY
pnZs0Jvoer1nP81qGU2tmtyv6QknI8OXYaYvD0x9NUWnmoB3MNW7NllBTC75QTtT
7fLHjTMmC/AdnUci3FXD0LDfO+YaCEJC9PwAsdaJb3TXQHhS3Bz/AbLvvXTgm0oP
11b6n2y2PPN15Vf7X/rpVQGWsRr2KmrsQD7bsPTXD+k9FF5a9OesHvsqqrXjPj1u
n9i9LWNaqh+DxC/HlN+x1JqKTmzOwimgU1lAR3S/wRbbkR5anVZCtA30qEHkdQMZ
t0EbbsLd351WsNlhWM+2M+BdaBLRbSZH+H6ufYhjMDawN2W0nEx8VZbw+F/o368S
CzBX5meJYnKPdDCqE5x8goa2Eo1Jyz8RqIIzzuoDCd3Xh6b/0ywkTuq0fwT/PVu2
f3HAXlJUjI7sdQ0/ABKQRBqOKzndDueMlUCDlgkekUWIqvYbsHmRFGky/uMJuIeH
CNBd1pSi54JpGgO7HHazqK+n3UuxR0SV2VzBehvZKTaMxSzjxi6aJ5Ay/C1rvf9f
iRflE79ppqJhvcaoL43ounSr8STjZuTGzAG+D7lZ2Nd6pyMZhI87Kun+77l4iB3S
y+iqidVIElJYxGxneRQJ/ZpyCWms3guDYRcMs77rXyIAGUUmAY2ABWAmj+eCbNjI
ndUUONIy4a0uc11aQ8RhJaNYF1l/7/NPvX8zyD46lqnSmxSI9QZ4elagpbCjGtOr
3Wpaq+c8zb4K9GOX/m/5bLtuYuu1RvUrwzbjwqZW3c/fcvsPZZRQDMcmbwJqm0Vv
Y8xscuPWYdCslr1zCK56S1P9dXrj1k0qjLBJiicigL3Nm5Xx5ibGsYDmsSgdqsJl
5wF2lh7cxTkI2ATG1x3O5oNMZZgXlp8B+cmdtlaJi2FhI3DetGt5S8F9hJJ2wMNZ
g6S5b09DKqOy7ApjsUDQn+75MACbJ0VUiU/JOVa3a5qEjghinoXe+6z651aomDHO
OOdKfrMMCVSmNv1qi4rUilZqpk6ig+DlZH8GvlsNnmW7m8e/s+ijcvKUb5kWrAhS
tN8Gw+IfCCJF9eEbnpOe3wObFKa55ka28hCe8TwF1Pye+bdUKdgd7Busug9IgdwC
9XHhtGfeRQedN1yedn80/Me5/sKv43FbHxDhgI4uvgkvs/wuWtP8CsUU+kv6XmTL
pBqb0yDumcNzsVk2IUYmLRbwSONj9TsL8IHYrhHBkUk9H9Evj+DfsJXmtwuEyd0i
YSaa5LNBtCzo9h15/JCk8DKxC2jGcvEQiShUzDJacRkR3DBp28irMSRQd4X6qDnD
FxSLDT9WFQaiVZOfSRdVTSjexSKiNEDrI8JkVxbGqATHbx6WvxQXUafQTjALSkQG
i+Aigy0PuDeThzO+kpPbx2HVYas0rt688CCypgrM6f+16JKAohqYwipUYcXRrGDR
XQFDwnO59C25PwBFH0zBtE1Vr2n7FkC/k1NMqXaeA4Xf4B8RQ85QLQAyUTYyp/kQ
4VLSnrwx/E6oI2UnKgLs9CgZM5vAYAtRhfE2Ahm7y3wsg9AlmRWiEwSlb5YNL9Q4
z70FA1RZzKgr+0xC9SOlK7UoTY9ZhEH/bkdjamwL6FCbLfoW1L2TqUrzglQ53Fxl
6g24As+UbJgEtSzDR5izd+noBJtYCJEllx7uq5frdlMjTEHcH0HygHAuvTTLD1sy
sOkmD9dxxDXED/2M8qaTkMBiEOs5KQuijJIoJdmNkz+IV6VNcbBYwcENv035Zaab
AdzKW70kkWBKrMvwDvvDMtgl1rIEPHE3G9j8LhM5XOVYghMfU13RmLcAn9KSVxXX
iLS2l3KjLCtRcsLyjSQ/cesPiD+XF0f3c2Utx2Pv35Ao8aF9CYvtKociRVQIHizw
tgNB6rhlCDPyA6Y4c3tK9mWcKP47ov+6TW975Z/3qh13oc22gRkF/6yhxXEbe2Sj
GuypCSgeSzzx7+E8X+UjXMTLeculA5zwFuIP0r+kIqRndYZ182uBww80b+HiCQXu
dj3iFwOYlqEWhHxKbQILon04uevrL1ZFNNlT4kj/1Gr9xRZ1TkHXj3g+vGbgzQuW
6bXWaE9RF2DDVVkIsldL/0HjLwADkeZZbp6B09FD/vMINjmnId8SU6kSXjgw32TB
aZr7FZOEgTDJ9rwCZMCEqT7xqDVO6K1V+66phWaeHC128ICApQUVsCuysXv76zwl
shopvcObzREg+OqSr26/uOUYKjDaGh/x9HK+wPRc3tIsNH4JZWUz/jXXTsR6GLMo
7ZW3spbziiWgWMoH/mToVm01WKZks9svSIYZTNv/ARVYh7y+BZyjdguC0HkSFCNn
PMwQIOgE49dwDA8L3H902znqeIGf7NUYiVkraYXVbsH8+/S3oit3UZzMcw6l6929
pUVDosHWNITCSav+w/EjfptNwo5DcyFNoIhmPKac9KzOhn5UzFqxBkmsxg1IkFch
Tz2B7ME/55nsF9wony36pTR0f/toXgNbzuNoLoZt/RMbU5wTsNtNAbbwGSDniiJH
usKUC1ZOi2hVORJsxdf02q+MJmzdkgh/ifkDXSSPCeMWA4CQukkjPk/BHQhRTA6U
UmxB0bDxSZQiTMVyqyThune4JsHJpOc7MftGZuSB/OwKA9AV+5cDQ7UGdFhmL88/
v9VvcSpi4rNtwEH8QsPQmCihIQI9OmNcSSHkI19/GIhSWJ0vLG9WKEcWggmDTNpj
3qwKsQW5nCY7ZyxF2PAdmbkQsEmobO9HuJdEu4lZNVpimOf9GH1dXRcv7uUhkQcL
ac4OdXSiW0+CI3Kl7E5iHmF6dDTc4r9ivooqAlL57HNbOON14XFFq+BiRvhDrAIF
+oHmFjhuMf3gmZVlF7AqN1XXZZm21DEtvH5aTchzTy3WW4uGPMCy7kH/nliLiIg7
NaxDJym1IQSKizJ0YzHHOtSiQNj5hQt29KtbdtbpdIsKcH+ZjARvMmDrmtmur3/W
uOUkN+Fji5VafDly5tCMGalgv48gGmYcLZymlFDBvSOfH/RHJy/kKX2D+VXTUUGu
roozGNneV9MGcRxQWJiHj95wr+aXprJGa2l2AnZ2SXzvH8iQw+CoYXLEnqFx5tIy
3DQZVa+z8JyRUNuo7ltd8Pzk1emwAlmVhJQBxQvYxyxpZz0newj5bVAZG1YbarNC
18ROFFYmfhJwdI7FjgIJ9XhcKalQW1maK7CNAk4Qe9qOEHjnMr3RzRxChD2iNTzH
ftBgrxlXr+HS1JbkEVx39eL4fn90jzUa/8ZPUUZ4EdiwtTgf5/K582LaBqk9zM7y
N4h3+Yqaeu+tmMW5dpnMSE8U7GNnzw/lvjdQKlij23z7RGyxA2SLuXhXnIsEZyUp
txM+nvfBsNX+pPW7mXqaXliyEh6XuMYtr7DjsBA7tOhxeElz8OyW4r1/D+oJckld
tjt+CGdwB6jenIFQi7UJPK6oLoef20sdMbu3jHyQh9SviQNuCFIRwwEAmRt1j0h3
GsW7YGetpsB5U2BtOaFv9uHnvCko9SOTePO9OtzOz4P3Ye7DA8+zTj4071luAhVg
CAnbHYIdWKKbNBB40kg5HtzKxmWXlYtt1bwe9EN5l7OHpoIRAxpLpTYRVjkTx4YK
2w3dkqF2moM2udxxtY+Sx4W/H8ogjBmmZAuVR4Dtb58tF6hX3Wf8LiMUdI0gjYgI
PG7tal8e1pRHEWlnAPCvUZHm4tkLlOR2YTzbL6NiPi2dlpdm43nnSDZ6c9nmbqNr
BF0zaV300UcFaXk6GnKQvytjEjaAjqzcuiE+NSM2T3Nqrh0Zbt4UMvPVnibj8lJx
BvqfbAqYNCqM7m1ZI8yjEUiM8eNnfngaqXfOCiDJiLz5YRfoj2/hLUJ2ONASS0K3
hz1K3ZstgJVCWC2L6awvxj88DSgzYABCMn8P98D8YWFGaKgRVO1khM/dWJsU7FL+
8QIoQZeHivlrNrpNvQhXcjE/iIAScattIERW+sGCKESyCbI9n73jgZSuz2ZNMvh9
evEblU/tUtyKgepaauv2rPRLGjTCTxkzR2j38wq5v8M13bhP8FVbS7JU+OKwz514
5SCMbACoJa3Ij3I5OPkp3Hy5OjTLtIe/Dn1UaAC3Os/kzpOZSbewcB2kwb/aM7De
LtrxrH3iRULpvCSsDW4X6kRgqMo2gbSgeohdB6rJuDhCwl+1cIrzapbrLoec7gCa
S2WBud3ODUP7hnSRFfSQR8LE5VTwdy8ND9vwFRIkq5l/gok8yM8ibmzIVkaQePeN
u70bfEkRU+oKoGeeXThTX4DgKc4Y2sao0LLqpAa16ci1z6ftnHfI1AywOieUUWBD
5Zn4QTdWDxy7Jz1snTbC62AhRDyoheENLVBCQMVGXdfLxap5FkuiczImsFREq9ku
5i2JeWltRxbP7I4Y7YmtlO8+BKKun+Xe0ZCpy9NMaAHFleOS87OSCT370spZkqkr
rbqZKMFsoBBOom92xmyzPuUH+bTZY2TsJEF9pFB3/NMaMzLAVhvIcOqSReHkDJCq
ZcqiCyoSP8VBYdvZkAcMcoznLdfEWk6EoaZlF6IQD2BQ3gUM1JGHzHUq1+TCNLeY
chWD3oRRGIHrI7N4EqX344cxjJsTkjk+X727zyEN2OlURh6Oqo6neGojsN48By76
IhOfFwJF+yTp23GgUxPA9rpRAHJARhX4/r44df9xLEcqn2ZKEHW5hBe55qSzTfoN
2NW+clfj8A9cW/JqF4LDg/s6GwQ0SxGVfscmS/KEi8/IO++eb9CpObfbfn8J0flP
4KPRA1yyD8vzleVkQSzjyoUffcKhazan+VNkLdiagiAIjH3vtfEL7Hv2rl0L7rPD
WZjulBeNCj4le8TGJnhkwu6lK0UHIowdFnrXdez7hSyDDFFnS3F5BWeE1YP7WxB8
9tLOc1bURx9ksBYxr7KuRsfEVaexpXCKaMHf0Caa5hDsHDxzYRjBnzWNMUUCVrSh
YmuSjV3CtO0IdrSpz8V2PX17LN/Chy5Y7UKFHtJ4bpcgmEw6aKDjS2LFPQxe8bRX
O12ritq8qrGAvZGDYW9GuF0Ftruvh1dXBECs8tReZf1aQxZgMU4rDDsn9n6kvxnt
UHCRxwrDN3fDcJY1aueT82JwCC/sCCxb737JiqddcuJ54Z8gVN90z1WkTgMGRLXJ
gWKSP56KmrbPtIylOykK/0UxW4wN4JBrDtmm/RSMrQVR4eMdbbRYoonNvx35gFVU
qrfjl06UoIci5nkJwSA+0UlNDIA0JWB0aDe36Y0Am61dSaFU76cqW5DI1wqAi56H
pxPEkh9tOyWMUqgV8Gwlq6dGORch1Z6Q61xmyvLT5xQAU2jq7quwQ9qngpUM3//z
HDDuQOMWwFitq0IWlIKQQS1MD+AKLfPJMJs6V6wcxMgUydKxT66elywcbYsBRT3P
WBkg0tFwB9Avq+VQ/I5BuJhlCekXEezR9IbPzmaaGtCZPu1Jo4QGDhVRYqkjhxMu
DO3LdPmk5GxUAN3fjXamFc2qUAdzW7r3wqttu6hDOLOCbpnpP2vtBm+Fl2HQlciG
n/lbD5kOXjyIhL86jhu++oDuuZxF/VUVFQA0937JQKw2xGOkkPhGlVYUcAcr/Vf6
WZf1HUnafsBH34OP52BFo+kGClYyDbk/JIbxn2U84AZDxBIO8bPcoOCSy+FmWeAq
6Udk0nsOqa1qtU++xpCx/ZYan6d7p2wKMirzfTr12VQ0knoktWTx67wqyVTfHDq7
XhC2lWWOb/NlG/flvhIbLTmAJmNvN+5aJ5joVFNFvDIK1JrIrmcVFGgEZuFNvqEO
qjx409+Bg86ryhPn6/C8y73ax1TfZc3XIpVTqdunZqEATjRsJMve9nHh1vf7rNjp
bfA34QjgHbh0A1RQAExS+uQ1PNWNrlg6qaAC+maFjbLmwXf9/n+G61tpUFW9gVcO
P+nCqzj6Yt11bfa847mRj+9wU/Dm3DjMcx1g4fIk+b6ee7vBiDy7tGhMayc13fTy
i0y1VHrgkaez0afXvcqsghzfJ1SM/5EtPtX+4wE5ewVmoO/kKNAaHmaslcq66E3L
Avy+tMWU1sSYC2CTczk0c27gMiYA/xvrJEhHGX2+kQySa0WIdeiikvNC1mXY3QIa
uejNJ/V73IETbnH4GtT96v9LDPcVfntxwEQvkWnVtc5OKLY7QVdFKyNwYU/Kz9A0
OOe8j1/8AJ9RJgn5BI2MoCYG+GmWCe5l1bI1M6Cfq6AhzaqEZ11z1yTOomZhn8bX
ux7YpE9YkbTSM1CWeRT/XHiyWuLr6Gj27NeWFlxJ7d/SGAnT0enhdbYcCLN2FPg4
O/V7n7lZVfB9Ywu9GmxS2vC6zFL/+6V1dqzI2t16P/E=
`protect END_PROTECTED
