`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmwkDPbsvoHBtk64VNFaX1cwsGN6JMb5BTCAoVYAZcgLYW/ubkPE8si472VVixby
O3yV1a9cbGyX0rUnaE+cfX89alao095oFdYHRNT7H3K6IVKEph8xmU6QVzT7Eufs
nJonyOyO1RsKFDhaPHLp/Kry4/nC5/Cylu2LB4b7kw0EBdECFpxwQlQnTOSQ3gnv
qcO8/hNTDXN9gH1ClJC3ZtIp7VvDrwfDMPRawLMoeblPbmZhc8aCo8Czs6ckdksl
UVppmekzjhmjCL6/w+d3C9bpimgvvw33vTmlJsBQWT+NuUI9735/1ZEGm2uYhM43
N9LXbZduOII1NM0tP4yoXAz5ymFBK0LOsJ+XryEgdYV6KqxmZQVozYF5OtMWhhms
w+tIF4xpWRuUOEJAbTyFoRd2R71xhNrNQl6g4kC/UJoLG9cgjQZRQM1DNTi2pssk
82mTyXWTrIl65aVUDgvk0u1XqzleFXrO8mPZbe+ORcyCEtBzQempXRHVYLTfyegk
adQ7K2yd15Kn5Zr+2kYpQA==
`protect END_PROTECTED
