`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+U1STns/9M6ksjz1ggMHwiUkAtnipjvQl8wJUYDdRtllj3JE5HMelLd0vCPwbvRC
G7vSb4P/jeUyNuyjeKwHn2zinbkBhK9Di3XenBNG+zNoUSfJ/6vzKYNVSZbd8uDY
HRYf2k8gGwuk0JvQXOeqaPdjSvPXqRZFsLkEDqbXfhuI9Uf9h+0lh1QtqdhkkUIS
dikunNy3sDsw5rmbkPrZy4shWt0EzAcj2DAgNXePuJQi6E+knWXZW4UJeSJwcg6+
aeYx8m4TGDHiU1OcNO54zxW6ZHEkhMbZFdim4tuJTEYm/WeQGmi5XKlFRGHQnWWo
SZd8twDa5Q8N+33fQThipPlvhZ3UcjgXGVwqJfkEvhjTUHZd0mjRs3nsKXklVUoR
ylsX38F08riCLzIDt824DO0G89P6A+6FtVZexNYm+aHp0VaxMGv1hbVNvv3/+IqD
s+Mm/W8IncQevkKKS7kxZatFr/oxmlSlqqmx39nM65B8aUc9VHZlgEckwDJFTj0z
j6+260nssXsO5v5R/j1BXWsmhLJVoIWef65dgMOIr7zHV+fcGMUPVPbQq4ho5aVu
GVslP+kJG5a+9oeHulbm+y/zWnik0YZF5BjkvcBq3AS3OtuNo7LBzITn8bGV+h8C
HDoxh++ABwq2XX+opakQcbmZQ/rqGBv5A2wCxhG7y6wFGtc5KkpQ7W1kZHhYK0jE
p78TgxGBK896GHwCyH5TMLkcAj83o2ynvwYfqrbrxCHLvr52NnfCG4pz+Ae1XBe+
GWXZ1KTpzflpmQlX9eHK4meO+GTWih3bs4xoNsHvlJ0cv3iDSQ4BKvfLD31YeJJO
WvANB5fp1DDb9/EJU4wH8ovlfvhkSizjPCmCGihDXRAV3YW1w+x965Lfw3I+8fk9
Z5m8tYdzX7+km+8jj8khybpTen0anmyRsYZFbaiQKSohWL/mSq4ObeCdgphdR0z+
GSxX0Cndci0A1ktOo/qRxNWBzb+GH07NKtXKavIXcWrorqNeq741cW3WCWMvMmYw
17XFR+JSm3TRopi8sVgX7eRZ6pUHED5JClvSnMUD9iFJfkui81SRiqg2eHlFr6eT
SaWXm1gsJl+8JATKNa2c8ML2W9owyY4jVkxzldjBnIQTQQqy0Yz5L2ZiZsRhOXpH
gGieK5T12zCRNjaoxMdsvTPRWAmwfsZLim1K9kTc/abmFJW97Mzqt348IMqgTbVu
u7dqW5Uo1cPhpBtHdA/k7uwj0Bbd6yrHPN94z8BLf32jQd0e7dft6+lQDEFFbXS2
7hKmCETTXr5We05h4VVxj3SRffJNaGteyvqyBMF3XtAk51e5VVJB301Ny3Eo5+El
Q/Igaqo3NJhG3mynKTMQFeuDvNGlSoq/kika+k3jegE/do1j5DjvyqAHV+6zP4UB
ZD2chHaOKu7big3T6ZxmAts8PzNSKnHr10hxmd7Uaj0IsUrMs0vTCGNHcGHWAlVL
8yijoj4I4+0RIqpBAIuYR9f0I4iJOkrRrjydGqmMyDlM4OnBhIWBlDH5edYOL66Y
VoSywAMG/5lp/u7izX2bRrWWqLROp5Zjhw0kd+ZN3kxFgsRtOto/Lmbvc3g6yB+d
v3ZTAU1U/ajVFSwGsiOvng5TUDg6y3JQ3SRecgJR3qpRYRzj5nZCyUZbcqAca6dK
44G4I5xc17MyW6MMnwNxoWvu0NX7CCAkCDekCACgPfoWM8reCxTh8ocfXr5p/FBe
xWNJN5773TlWMM+DX1w8ySiVDOPCjtD2LMJrZuGhBtHP2BcWONrJ/TAeHnkaOmVd
WSP1fhm8B6k35l37MClw/1yBpWS7c29m0A2vMn5X24bMeEa/iTyDRwzkmwGFb49a
6kuPGPYL52m/Hj4JOjkwhPejOGC63LY5SJxPEancvPSCBOk0GueE8JuVfz8kx093
ry7iM9Qpm7/q81hVS96bzg==
`protect END_PROTECTED
