`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CRYd6UdWzwANne5pIFTY5FLag75iig3JSqOcWX7C3O+44STMqQ7xBqfK30wyPuD
y8wXuGSLzxFT8ZdPz3P6w1wAoKkHyNqLJ6RiookogwDdqnrDhj61KyHa4+ASEfB3
rwpEXeRNj8G/8istE2XoOj3babLDvxaTAIzISimagmX6ILSMSxMbUDbS9VlLwHMq
GnpFcmbJLIDABqvFbqCbINqQ3Qepjqm9x9E0zYUE8Mt79jKdd/THjnYPnwybLWGG
GBIJQj/69lDZEiqlPUK0qmqsDIftMyYw1tFBnaCVavtLANqpwLYM/+HFmSf2Leo3
sYWRwAKvRz9/mW2AB2UA+lYZY/DegaACD5ZRsEDOk8RV5YNTdUAv81CyH+b1E20N
A8n0dsL9wwLnUxIAWRDv87CAPSnUpoxpma7APsYCugEXFNdINdqMz4sY7VgisAt2
c7231PWySjTzsUuDRyymA6woduXnFVA6QM0Qo52RPnJMTcdDJDhtDbIo0FglVjoY
VtIQ3EYRYmu9tKZP6x+RcB1vUMgRawXlaVOO3cJaWt16F2GgLafRsTGEF+z3QuTw
`protect END_PROTECTED
