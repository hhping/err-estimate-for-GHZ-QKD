`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4S0UeqGdhCViV1FfjXWWSDAW3mExkrJDaIhKEz407+TKsGUMBYJgFc3/w+y5o6l
W9tdFatpnZqyW1Y/WXgyUqDKsXBVPHTWwoU3OnTIslraDcFag/9h1uhG9cJOGFXC
nXvvSF+p1v7+LtnmAfZgjWiYSEbS42egz5jJZYRu1SUtFNO9sRWT888TFkxbiTRF
Bsns+3fGanXO7zFRb1Qpavou32SMD/ljAGB+qS9yHwRUTrm8Bofbaqt/mlH4V/L5
pN6dj8PSG8E4QFhlF/qf6E8ZjBsgr3f7BAak3EOORhG7YbPk1wT/gVTBFns44RQL
XzJ1lhqtL2matfxr65bCdYuoiSA42elTtHWtWgV0l1spD0Rwo4cWQgnR76OINPd3
jzzeRgIOlKQvZYVRBu75czM+CoG7Oqf3yR8aDvurloH4NExBMNhhsHpAjbRw6QK7
uxEGV9lymLOqtOCjjpHmILYWJwfPO/F2HINPewNOEdk4UYDw7hbT2fTX8KITJPMA
lOKY+364+pO3P4Kys8jrHQhsi4J/LB5oNONAO7LdJFGF0qhVEVv2RvUC2VbVuC2P
JebPUNwgp6ZYx+B8bSh87CX0M/cjJ57J17RGvk2jMLkwC0F+sFUf38/EAk1BlO63
eXFstrbgLOV89699cLOUz19s6GZcJNSIg4KKDmJplwVoHfYBfmi1qfyGJG2phAld
KeLFJBfWUjbbphhggmAxXsmryD2tTsLdTlU6j3T3QDFOOFlNdEEvJ1EcoKgtBOFu
TstrjZc3IqBY4yropc9z3gfaLEXg0DLJle8ERKJLGLyC8FnDN4qKnN0bjj5UN/dH
UtIF1Fvpv09PYjJ6hkZHh3uddljB82u8iK6+YVExUXI=
`protect END_PROTECTED
