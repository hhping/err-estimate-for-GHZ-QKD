`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOoGHY4eEtZHhE+iGbrNyfprVVUbb/LVQFTrdpgHOUaVGw3/I/1Qw/26oyZUD8j8
MXdno5FEDsBB7EXB5fAnukoDRYG6nVrFA+3hVc1ExIn1yz6uki+xWnL9MtXvpFGx
kPt3OKX+oFYYqKmWmMMHwHLPxtjhJazUOGpqm74ovGWnnRzOpxdu+vooy5a6Ib2+
ZhQm8eLT5PrJbCZbONkKAlNHiYx1CN0WWl8WqH0FQv47aXNxK475QGbIWzxZQ9FM
VOApu7ZYdHv1v40kghm+DL0mi7c1LLZtIFL2nFJUf/nPkmdpwAmYW1eG0VD1vFjI
zp6RKe3moRTDJf5v38SKlwQphLohDa1+HMqNdPSC6AQorpJ/XspYdhnnGtqIku0e
cWouG4zIc6dlvn+QoVUino6VCKxmkoGJAPIZuvKxZAPyM68qigZy+eLbubXm7cca
I5s/fNKoqtng2TuiRyAnuostwDX7/znYOEJkm3QrQoWh/xLMZiyD6QgXxcmNs++/
/bEGDFOZ4IsFXQzkXUnvYgir7G0kwl7xZvKs10J9Y5qpVTe3RiD9cdbnXFxw+xSN
kg/QwbhpdB4kmsjUro63IrQdEh50JYDWSxUkpzzKN/QAokAvj3ge58qBvd9iDCXS
`protect END_PROTECTED
