`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWZg+yaF+Oa0uKgW+cxU7xUFTB3bEQojAhzaYYiZD+hEPHfMYazJqUT28PwRG/FX
cn5EeDPgXk72GjDt0t0qgx4TnlDpJJShgy3oioIKtV6tOlhSVy6bTZrkT0dSyCiV
DcpLLcX6GGPhXClkl3dj7ODZRAE3zmSkOfgtmgTY4A9QMQn2I3TgKvWM6hqru/hx
E9Wm32zzkCgBFd38h0xK6KmzcjqGOcZBuO6xzuuBSyYE8jxYTOCCAgkete31i9tT
Nz+XDbmwes1iIneojSi6+AQlQZ1zI81aHvTjBGGSQ+0sm0Q/+4/Aw47o7Q0kS+tB
eqRkOV6O6CfGrZ+mBuX4rDVXZ68E7tH8Nue+GjCMh8xQfIv3NBSnNXI8ZzJ5b333
YSjWGDhNqWsMY4Z8MQOyoTU7wsFCxuMeaiy8fWOU7Ypz0Fzz3CyazGmMEe11COyK
EwoYoq7q1+zP3/LHd0Vvx/lRrnFFq0IRRODCj+zOTFybygyHrQZ1/wmGLpGHsbn6
TZeqOVfCBSl+W0Y28uhy3idNjXbWE67Rot2VRn7hqyWk5lbJtAle6nXRJFW8HWD9
mq5/1pMdT+98ZTr8RsPibnhx3Flqjt/9vNAk9NqStaAjOhqEk7+en8oaA9KPvo/E
/rVxpA4opBj2RPGjgsiz7Ndp3mrs/7vGHq2eyRd10xShgIOJFlc1l7C+GMATTiG/
JlDJaXpYiikH5OabVIEBZova5SU+NETCPmzuBGzmJ+Lrju4ZluIeUNisQ7B3NvOi
Gsq1sur01tIIFhcFoKornYv7COevRIMcLTS5d+CoNDdjOjPO9dTiyymi5UtEeYri
5CLPZ8OOVaZmrEBdmX3m1g8Uk8AXujqgTRj1Gn2U8oXqbxlxGpo8TTrpfLkxMSsA
CVqayUhVLvNmci57igZf1yBeHtAJoEU3/EpCk4iq99hXfFGUkMjhauE+vdwUc9ba
UocczJLpiIIsyOi/m81bTbx7EbAPTcq+gOzL5cBCpud8z2rK702H7PvPxDDsXwgO
czKuCf1ioGM34zENiOiqMM9P8lW4Xv2mIEptJ8M68RQfLRHsFicL2U/1B1X/QLJg
E7T1fXsXoEAn4In7pd1KuMUIecl6jiFszv5EpQgNCnbMNt/mmooFEVXr6ucHLYKg
j1fCcdqpHNnnZyc3b5v/tpWzv3GmIApz31ZeW6mKdAD1Io/VflKHbgWJmdEKZ+BB
vviyDYpgEktsnJ1y5J2F5jqwqv8fjfckY2+qoTFE2wcdcQK+d0106zZwKb7Tc1N+
XYC4nqxiIDr/aHWBOagAGcmt+ixul/nw4PWZOCoCii/KN/PQ2U28siVkdJyRM0WV
StcafB9gb8q0llOnH54hCEhUX/oyPFTH4ZUxjRSeSlJ3BvdSX95Bzut4gwcQzZF+
vIZr0kldRhrv2Xa4NJ6IXsGWvyzQ8czQF/x3t83HGjcroR7S559LeSbnvwyZR7vR
1n72cn+LN5u3X4zuQzP2KmnsnedTWsgG1FQNRsO9glswwMAoaI/hF5RGV3LSXa56
qXRJAf0dULvM5RQuSbIbolqlhONIF42KcUIqZonSGoDKCP3eQJI1t2CWMYJm6BAs
Rdueu3lidL4kHpQVfHUW0OEJKTr3jEgxrVtXdwtOlzqE4910c3xwOEEjJK3XKicv
uzc5RsgXhBWxgpI9HIHvLV5fkQpKT0rOnqmKadxNCtsPuTHMkXVRBx2mZSdgx1gM
SWDk06mb/vu9OpctyZg6PgINSwS7+gnLR2U5aqz3DXDP3fgpUSQiB/so+8iiws2O
2G9bHe+Be77bwzvIWQsNoxPKqQLoK8zXs6dtQPSR7Q3z9l5YL1InyAiBJmCvsiR6
F+EXkL01OkcRJJeLbEQWL0jyUso2eCPPPwXJzZQFnBPaKZgMKvgEWbdVE+fkmrj9
AFwVQxAEKf6gghrlbycb61XJQ/6zR66OqUttqfA+IferF8CU2gd4A4yX2UY/vccP
v+MzvGteapWEAhSj7JqSoeQZd+gn5ZmasaS2TtMg2iUu7/hIBLSl2LwnCTHxk+ra
vwEBEf5BMJ6aQbI6GOv5aRbcLrnHmC+4Rt5RD+pt5icO2Q0ebxYSgSMNxrgKw6pU
rRbZWHxfYwfgjikyLLeVSpExdFiwMbO7gI2XZQBoRlbB88fZh5N9+mF7ZCCwmlNg
8cK2GOKFhLgi20rqvp46e+JMD1bFVMh6HVSg5XX1MhbmGsZpw+uaEyzh+a+UFupZ
3Su+FnGUly3sCGZabhSBy24rDF4ZmxNYyxYDXys8H9FzDe94KvDe4x5fUqPu4Dmo
BQgw1omY4uAxRilE90Pxb3sGnyuBPS4qocGs+4+SNvlGnWAqv40d8okSdN+2KSaF
DPU0EG1uhlo2rK6hoZbej1phbopFJ90q8Xm0BAotFeibvvcQQBOUV0n59AIqUKxw
LgtnZYHv3IBoG4Ovcu5FWloq0vTJauKxaECnDakoIVmOY8fU137fuOFT1GgMqrae
MNDtLPkgHO+7BGDKR2Gj21qvfTkic7D8MS3xifvBv//6RDs1B9o8NATK8lo9nR85
74nhe0xvPlIcNGkEj3e6bXZoE6bvocoLtiBIr3ajbtnoTwvbyyXrYmCPb45AZhSO
DLJCpmgEU4VQmMhoeHTfVNDVar2obfpyCk1v0cOdC0Mk5UGAMH4QOd/8G3ZRU4RR
O015YeOlAbZgRGIL6OT2QbLibjzlPyK1TA1dyyMhc2ymtGqx7UajU4lvZxdWD+pT
2NKQiWHOjLkXxhIpCPow/nUJ8y2xb8w9oPIzd9RmvLkwMRNq9F7QgKaBZxR2pIKH
+EP2/eMc0oKOS79YkoK3WIFqyJQpphwgKj9EZIswXbX+W6miBL/JF2H51PbZu8Ef
wvuURPf9IrQOdFb16vPvFRLLZU+yIX4ND9fBVvBKdrOi108IzSc/VG7P6nzM/atd
2gcdtiPFXGwp5CothHiYc2mp6+twWvPJ9vlUYR4QV2e1AA1cjWnwB6qLS0ltmIfO
hCKPi3EoBoqKf2TWPhp5Kce0hOt9+CcImRm2mxo2f6QcNhIScbQ8GyxpRge6juiZ
xWU/D1W2wRP7TYiBPkfIg2bQpHxY+uuG4X5GP1S9iU45ro/DFCyZBmQsDmTihNV6
yeJx4ackATRWd9Dr+mhgwOUWvk2iQutCSdKKLUmxUvmk4azKuMqPT8ti1egeYU23
VN+PeqpB67+5boXqzIM1E1ePePI3HcUwPMtEzM20F90=
`protect END_PROTECTED
