`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XbkDkVSvBiEYaWBSXPHQCIPHnlyYARHjq+CpTBn0JD2CMyC22GFwhQs2nlgOUOLK
8hVpVjr7nmLIJyCcyeIdpeGPRWm2EBIEY4HJ6hEjFXwhgnS/U2rL/Dt5Z/E03vKy
Cso/a315DcvHq8f65EWsaWAvku7F4t9wdBx157d7ZAaZgxz3LFYJrUxHMyKRRxN4
UiwyeLE2RpRaUfAQ6R1ylHYtldxg8GlTs1hnbmSEEdRBLb44j4lYJULhk+UBSZi5
Qk9g6FNQj6E++7EgROnP6gqa4YdUSeSLzrdiFo5teGRqFo7swHJVTEdLx16X5lek
eCIHXGTC1mzDml4y8DQkzox8IQvsy9vISQSIdS5ddEHv0pqTIVDCrdaa2VgfHOEy
3W7pSDExcBukKHcQfjKw/eALNsBep8EeybVpsczrwkuJnF0/nQ0ts+z46RaicRmL
S+FDsmVuJz1OAJg8X7l4XvvywG+N/qYefUSIPINW4P+d1zL7MGIck0DA4GiZixek
aAtfNnzAUXdC1umaVNI0Pi08P1UNBi5rXu1ZRofjRuxYMT/vcjs1GP8YPV7wiBsQ
brD3Tgu7VTsSfY6m0Lmgmo1r/TIdjASt667iUCBOqb9BXcFvkMhh596YxfW2NTgl
`protect END_PROTECTED
