`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJ9D866s9UGhXtuCBCz/bgymM5Y7b0Ifr0vd0K+ljhSjL0Vf2MfT7Mr9NIlGsnyz
az2AQEHyRdsannUWw+DgqbltlF1EhhM+WbCgHvqO0FuYWcPiZou8j4whsxSfDgh0
HtNQq5NoM43JqNM0EslpOICOdtmlOdco0khaIdNPTkfLoh9hHqIqTcm/PJVAbS7/
jyWJkc8KVkSADB8aK9vQPZbbnepDcyiQMIyYcQrY0OsCGpGSAFzaOwGVzf9TY6SR
eaWtmgD4Lz/HnxSYeEaMgxMi5m/nHRceLgjzX9SWYKPTZTONOcFjph7Tfa1FjQcX
HPpU8UszjBGG5WYzMkdVHDyaMe4QN8ZyP2PptqFWUH6+CGw0ZQ+D/2guPcaSXH6X
wc+aszni0K1+4gHrvUcKXXy/OnDItzm0d8r9zlmSD0Sr2boeeOya8uGiLb+ZojSy
0EHdXsGLu8BLxeV+y3LtH4+s7JXSGlRPY4gN/RfWCogny0lNavM7656bzHn4xP5N
lgkZqZGULT9NnA+1PbmeueEudHtE1Vl/G+rPouJe17gOqHarem5BldPaGMJnQ13k
Ic5yOsqAXHIomuJw0Z2/ZCXc6P5vj4a9Yg8MxVwa4f9sph4Vg3uXnVtRQiD+C8KH
LWOtkUAS0RvYnulsBOv+TFIZIno+AgLCLFaxDV82YjEHzz+Wohb10KSI7+gBS+Tz
9upLaz8B1MwNdfloJlqi4+VtXtsdHwhblGM17vovO/+Zdw9miAVL0QGWiJJqx+oH
n2yD7cXGEbVYRyvDdUfjWjmAYApJpQu7i577LE9gZxE8Q5IoBg5LVWOPUgeHAJVS
lQ78PidLjDPbh+q1QuwU/d5k5dnAnuOgSILLl2W4TAho4zDaPHVMvUFbhoLrGHP/
LQlINdn0B83AyUHVeCnDzaVzrC0z8v6BPa6YYUglF88zX0lYex0OQQ4XnnfdFM4u
cpE7klKRqkRFq/J3SE59lIhVW7Xy0dksgp+risL+yEJSwgRLpq9QmvmtXNjcRpYU
pKOQ02/ued+O8qf53DP59osZmWnMylJiQZCsdYNn3Trx89Ad3Prw07UuZv86FZPZ
j+Upu5KFYsq83z9jjECSNlYF5xQZx49BvTLoUX8vT39J3FnBVDoV/zionWneJYAl
KLsZ2f/YlZfQlKys1aPs3INWo2WKR8zUaQjcaMQAG5fO/V7hWmWC2O+oSVj3OXkg
FThQT4h5tHUPoPT2g+tBvBnunC5WXdU7P9GJbgO+d2cGQ3HkfR5eOCU3ZMt7tbTs
f8YndDCKpvjJ6rjD/S/PRhxs0Szw/Ep86ltUZOO6NxqB6BQXlkKAHttZycKWRIFw
Fohwu1+qXWXdZeYJsALGdR/FLos8voEiN7TeZwt2Xa/m7GC76GY238s23qe0CLqQ
DqKS8Nds5VSdccWaNTu++jEYjTWLJgD5OMH+BclZqyliHNCxrMPkPEprPFXJr2XC
uGH6v2odclktJ8I+lVEWR3fKJInM9JvglaXAPMgRgvC0rs4qbzKVgM2T5q3jvSZ1
gTr8bOwdkD2xrKNLVPE1j4m5b6MDXEYpC+QCh9jr669g4Sk2kB/8aZwWiLVNZ9ME
6qRCPq34K5WJQn5UkR864ZcjY6c25NQAIO4sxEjmRiFnG8ctvesZ9ljYsOP7hpPp
DTiV1pDCFzoLfHJz/voslmr9T2QJXkYbNhSggsctUUeVCfIA429iMoMz9uhNsgz3
okXcaJ5zG+Bx/xp2Fn8E8CnetW7cKxzl8z/eRqxWWI3cHYk6NVQQ7nGbYAIeleXJ
8FW4D/BZ3o5U15qu6PX5+Yo8Hzj4oYtXaTx7NcM+EHgnUrw9XLdLS312GJsihrQd
sSn1zvkeIVP7Yl1sP3o9K2BQdKn3Eiowyi2m0XHBRWWcgF22YHDTYSbllvCnPG2C
mOhrG5WBKd6/1lQXoZloAQQEMmh+h83ipbx2vlAh1Ax3TnFdHJTNmSOiV7Pbm9se
tW1Z1OUyBT9oj0uCBFIKetdX2Hge8B063dsE9DU364dhzpfnyOYBTGE/Q4BAahpd
8J174mTf6e4IiDJbKrOjf8ByVZoG5cmewogtDjm4AabPyt4seYlitTV4EPdrSG0j
m6HMOvDBf3RjVVcvCscVOgERVNvH3G2V2VeBUqkbltG23fkPFNNbiTpjR0vRHp1R
jKzW3ZM5fSlQvVPCD2WiMdlORhNgDpYa+OTKF3wJQ2Zm6CHP8jj2xqpiFOpR408/
6YJyffBPmr6HTbLO0ybaxIoO+k+fnH2n7YzxJxq+wsmIPE5JWtZGLOZzu1hGj1n9
tCSxmtM/JWP1vclcBvF+3vZb07W7w7zvV2KyRPbpPb+6Gd6+f8iX9hc625ImdXUl
Y3Ypo90QfvCdb5By3SVHgQXqe4non6or3uaGd573qeEx174kWzBfb1Bvb0MPnV68
4C/yR/GkQShyWv2a5hcl6B/GMS89VdxGK74Q5LfBXhxJwLN+tu7VQnU/XX8zNepg
6IXEl+C/RBeV4oTXR/ye3P0hJHclPCpcIJmG6IlvmX5HaQSZZHYqtAzYWZplciXO
DPAzENVvKXJw5ixToRZTeBcPgxi2MYWn9PB0jhvba0noOcEfj/K8Mhj+b2Ld4xMY
t/EMXHdyCicRd8/3n+wAgmDLLJH7M7h9zGzT3l66RuN8TOjEXZt7eyocfaQwBLL5
V4tvPUhgaDhkH2TyFYC3dUm/gUSF4AxGN6IPqwS3aIDgyKjO+OMcvpn2oG6fLEBf
pJoHxwQf4fngmRXgi6Baynbx4579j9gKOqM8RR9+zagOga42V25FrbdmltTNTAYi
LDABpaiwNCczdIGV0eN8zBRS7I+3xDq+n+6ayf5+xy1VKnH4ne20lCeXw8cBpGCo
3GAUylRxYscMcjs/TltVco87QBDRaq7WI7b5A1WdROTLIiCAL4tQv+IpXkFaAh6p
F/79jnv7MhY34uE8nVN3VN+SXzYYYHk+0EWGeQAGMNVtXNV5OQZllkWgCJJDio5Y
LNYkaB9jIuTLbtxUAttUohi0e4oDgHmsdX11Py+BesIzEEtQw77TLFCabak7DTXW
UjaW4pthTjafcW0HK4kWvHukmzolS5OVk7iuBTEPvAs807ZgW4Znk6lH+i5GABKN
chlE0ahoLPsSfCXhSKdJgfq2UpuCQ6L2+G7ObkYtYzZm8OXlxcAFvGbBSqRFh51+
Hk/Y+a5TomJ/1Da4QRN2PKT9OKv86QDZsMUJhVi6+hqW91K/eZtZH06VTr/geNzY
VQcgvX7G6dynvAhzmZimO9KdgQxOGwEVqxW+yjj45uBs4emg8F3p/SyHhL3hpnjh
H/gmY9snOnZsXHFlWy8RXPfJpJajs1fIAm7aWDGKVUxTGBnpzxjd/GHpUJSIUOcW
3s0yp86WpjI8eAxmw/kNEBm6pzmHapUFkR6vKj88fDv9Byhdf2+1YKewEaHsbLEJ
tLnf7aRfbLcKDvALZuTO9ToCwGv1jjpxj7OGxphywU2Dlq+kuD0fUl8s8nCB0aXh
DwtTpv4MRD6y+XvbmLIKAuBQeKGKCRvD/vJ3VLrHz42JAJa++ygE4XxC3hj7VH1u
dweP8vR6DtHwDBsDBG9lutlV7FRvnjwrDtVTMypknP4GYntvW3mrkzDdlZGwDj/c
kPuy2oadOCfRqWH1lz6m9M7cKQuwd8cWdg8kn9fvNRQbm4Jx45QdRoRbXiR9folf
2Pwx6F0wuBwIIXOaqIw8nIpH88OY0XzoP+/8HFopYXvdAAdrODf76xYVDb8grBda
1CInEkSxBms0mN1IaZ6HCOdFb5ekc9ddYjlzK4xAVhgZolhOW5DkW0xS6sHOnetQ
BgY/5ie3hsAR3WlOZkFxjsCjAAprpVcqemfN+ZJn02QDROVmu6sQpApKvjw5+ZK4
KMZgsdON37eXgqbP1nGDjGCrYz0C3dPnpOP1lhHCyWaF10hfbYs0bJ6Rrp7G8V4W
s55DkltuVqsyOLcvQqPqpj5dhFa9S6o6bvR1XPwlj0EKyhVELXkM+s3jq7zAhD7H
RDyZo2Xy40jzUiQeGXt9i72FFk0B/IZVImeJdK3ErxQ09OrJ4giUIZSS+rPdyjAq
8m7tKB1emze0gpJ4g/Fgx5lyBIjvU9iR549uVFKdcK+olfB/cRbqKreFS0/fvuNX
2oXlShjhwbFzq5N3n9Q0+fJ49IDAoHPLxPx1ZI0rBeEYdiVDMmUiq84W/sTz1WWU
PfzS7/jF1FKVj0i0r4jr3lLLa0tFcgIjWeGL0HUM3nmJLOV3IN1JD2qzT3HxVs7D
9zi8IfGre/oqMWIKIwwk0uhmlH2DzMJ40yobzPUNP3f8up3LvKqCVyWYTakmvzlY
OlcVcXINhLiGUP57S3MMHeQj2EYpreqTszAvyNljl9Db+x4NqNKumMXDOVFnm1rJ
DSMOImTPhUoG2QNFYDE+rYCVe0EzReUnfzDzgrxGQFCyyahyeVjXYkZYaNDegsX6
blXd8WL5NjT5BNCieyL1wAClh79arQ1ADiDF5qMq5Zpd4wvPuVOVygcvBCEKuyzO
lVCSwqTZ3J5O7v/PxztjW/cRHsmtLyRGl4XSXZfvA8ZQ9kHO38OoYOh29t5Z+GPQ
iYYG6IyVwUQsJz7WZnsgQXdLdqVXykE3p+Tf4Cbl4TmdovxR/KktbMVXjlMWvFT0
O3OqTAFyodx7/gowGXhIMFulJ0F1YgYeb6mlJ4wMhivouROhYLOMu/6GzbhgZRBZ
Tk5mMCeuc7grJOZwlt83EToNtJoMxNpzEak7G7rAIN1whGLx5othsv05I3He9RpD
8pFy+zQ5dhSL+IFk9L1Mc6ffQZtkVRFkcvPN/oQJv6Ulxpbe8r2VZpKXlAnOjKD7
WvZCRrI743ZKBvA3xTZNVQpH9rXwUl3/+jZCWIlFuIfiQa5FRonFXSF0f4agFs2+
H71cSdD8jTuoKQRX1XY0vrtD5T/gJsgGCtfLEkkxOehg+tRUVzzzUbYvBDFPShmd
Svvrip4wh7IAu2uY8DRnMvy+Kl9DTnkLPdjWTy/ZvgV3MD/Jkn4f/j6Mo/wogaIf
gkeKJ6KQEbjjRNbF1cQGR4sZKIr4Kxh/6fkzPFrWQmh4Ot3/YKb09jXD1f+a3G4J
l3FM3cBPQo8Uz68Szictsu+wCkc3IzGpTRHIE5P0SsDDKy17w5unscMONoKZVUv4
YaZFo9NeyNO9DsDxQf2zYLwm6pzktwn/UvkCWngiHVG3MC5HRlR1Yl1iOmYGBIjC
1DuIQI1rt31e61XzK2PMuh7oILVEZhnwnFzBCLB130OOPYSIQwIPmVyh53FA+aVJ
YiUIqQWv5HPThG6mRUZ6OXVz6dmQXarRf62YGa/h2asKSCXFs2VTqFGPsPqe5kQV
bVzRRhQJHRCQYpM+1zmS/wPk+QFbwxOIj/tNC83/eILDfivqrHC8pI1Nwse3X+sk
ZxVUKgvWFtYtieaoE+DGhJ94avETeKjsQ+acNCozi+HYvh6MomjyL2O1ps28dBgj
2aqzTdwypN1umOCDanNyc0VVwkagTYykYAiAQ/AO6Cdobv8QnVEgrak2zr0RuKb2
vUnhYRwUIyU/rtOdQki4q+S4LRhWz4BvGww/9OLKO6WtyttQuPiSTp56efREw6Sb
FUWtG+VoN6mMgIWO251oPV5icCfY3jYmpXeoaijDaYmeAn6xEFq2flo6wCDQ4vLK
mrhUYKXPm/7nrSpiJR2mQH7IpYoWC36066wL0MSsd4KSptZloCVJ7q0txmc2c674
rRoB6EjYfW2GRMoVPuVh6ZWVUPi0k9vWJawmE+aSYTZ2AWSrvKP0IkTLDd4fPxhS
OGDEB0iYs3Th4X21hHNcpQK/H2JTudxwRoJvGfZbhBpFj9+hTxd/Ncmi9ayM2+S/
nloaEF7FuOW/HUwZqjv16jOfiXRnkG07dBhRQ0KpDBvAU+6bZWKFMHG5teyH9kK7
60MnIU0YbuWgp5rXWo3W8f3Qzw9+XWUcn+qBwe4K6URwCNq0eOE56l/h3HZSrhin
0H1IN3Ms1jL9tAXC3rT8n2gG1IqiPSZ/UJPQb+Sv3WWUP4+LBi+dz7LJJ5GLS9bg
OfsK+rVEwOsRha7J3Ujg4g//7PJjid1uA0pjcyY7O0J4AIfBErNc+GZmtdbXhfgP
zM4Gi/kYf+HdAD8iHUQA5kDf86I/Qkn4s9XFxvrcsvmxGO3V4d+MsnG6ToxxDyqH
x7/kqzs7+2oe3kiJIA2Km/Ro4EyNvZBhCmMqQfX0FW97E1itTPwgYXWUBrQn5WvL
X6gI/i9XXq96C2gOrneIdO7Bz9x9Qogq5UKc2Q8QodUbEdClIYPKzn63EnDf7OLi
bLMsqNn5Fl6HJceeNer1QqU5BJ8rcDMQOrUazbaHQUnC9TECi40uq0hzzSfed5/Q
MtaQIY18ucFi2F8gO/Qutu3RActaf715i1a+AHsRWwW8g/1y06Ahhrco/IqY75SP
2w/ijBtm4t9168D/u7LISlcJ1NlIDEfITF4sIuvMlx3dimaAGJD8AM51eOfWTqbh
wUUgLff7lPj2OQ57eOQH0TsO4gDdwGUQpp7+8MD9XUhRH/A2YAT9VgScpuz209e1
SmDHZqeR8yx3769NtVRlz12Vt6l/loauf2hO0zFPSPMA+WZt0teqjpEsWTc3cfCR
GpQq9dqG/OgCkIrLQHgqQWCVD5OGsErSreM2831DxBC6N/48r3XxaOIS7M7Sxf4d
GRgGi/KBGEGdPfa4VQsFzzVxyHkNtZxF8r0YQIK3UPtokeQKQvau+R4Kh8JVqNSS
aOmUyJcK76dvGlzDlRnSV7c6myK30+KSKRaGV53Q1pJPlzs/Jep7S2hACKdPhVPY
1Ln4E8tsoxJ3P28YNrXep+GyXxAJoR4V2AggJYn2m3cYgI/uhLQtDwGnwVyPKjuq
bhDDgmAviUjqfWKlzINqztoENSFpN74HzT5ly4NpdRbyzjwB1IVzKjEp52bIO7aG
BO4D8YOKSdcj5FuvFyfJ4PH5djDQ7RkKHWAX6wefGRM9XIluFRhGCyeIFWXPxWkv
yRmT/yJFevvmyIfk1woYeWG87S78ipncJkGRmX+gNVhyUIaf9Fke/wGQ/PS/yVA5
QCyA2aP3lGGK1GCjrPoKLjcsBPjhd9nmk9zIDKa8N+KY+Vx2z/0ywFhScH9PuhMm
ymDsSMuJMsUwxuF9m7WVoFRiK+yLh+HoKNcCuX+NDaTXZ/9uC24C8i6p79UXcRcz
cshFhaLGxR+2egkfOIDalOpc3STLNxr5cRGPoOf01o8CJYgQmhsr/mz8nVKEQMew
EkYK+rxHOfWFi2KQC53Hez67P4pIbGalaZ62dv0FabDEMLsbQS+qKXYqGdn8hyt9
tctfhqcl/F1+AcP0yZrxhXUL8gwMIRU6VTcA8ag3ha4b9LJRRcfZpNwVLtVwXCLK
aGHYekzhEwwkOnIvCtt3MSWlReA4hMVYEW4BWOzjHwdQ+PEyIUD0KKK6hxHg/8Bv
veCkgQWn2vzd8IttSbpUCbHN13KRMJisSi02pzzbOx5LZGx6QHb6wo7NCAyo4F3S
EQe4akU4DqUIrP3Txx+1RKWPlMr66nrVWR8+FvC4kmg6c0jWSMInu9hU+PWyUigQ
fW898uLramQT6oa+C9TKwgPVaxHy5S/cE64rCA5IaaIJI9H0Md9erUHuSxZdS6Xj
cH80i/vkPvnvgsP0f1obz6T3dFhDduDfu7fzAVk5D1YUKIMDYtH1pB/UsDvM8YS8
yqS7iE0JB8NF0FV/nzG1HIIKIN9cCMNGhfDf6PIUuaOZBI1UcCymN6bzN7If9pXX
HDoBbS2hIEIa+pETE3aJM8eKuUHWR2VT73UOlUBRHhsXsG98Ur3k4sxcPvjF5m3h
sotT+o+yNFNRpGwm6VZiMivo6b3df5NYrxmaAgbrT2xWKWWZJPfgyoBfrFUXvO3D
SpVaHcQCTz7ETWr1Dcm+zlF5onyr1ErBBxwWU5bUKg5Gmxqt1P0H4l15bfCBQZIp
cWAmKbQmOuPMjYxv93dV9FhvgSYamFLxOkiSfHECRv5IvZMElx7LSHJCMjWgK4oT
udpgm2eUDpRVII+KZro9ka7KxxLiZKpo4tndk7ayqjfM1ZqSbZlt3fhZuPRjiRa8
/gl6RVCuRgxOgaHFPSunSpnchOZAjczyvXf6qtyMf7M/aFcq9So3PUqC9UH6PL5U
STX71+DuD6NqiDnMfVCoWmdbvDahG255ZHJ2jV/4Gb9eHe0IBL5SW16m7Sj5Y6u9
3ZWdfYtTZrTt6zxnr0iaLXfbRTSCUILfkZzgpjQvHe0IRjKnbr+oEQSJRvDRakxu
bgHV/eqv98pa5Qew9c7K3qBIf4UGTJQY/bBhhPJC9SH2Yo2a0sUDzdIH+39o0+WL
IY/POw+YbdmPNOmyFcrBR1fKvjzZckeJOP2hGW2RkN5g2QiowRjxImcjTtADK86L
GcZjHCosZWI6qL5h99Nih2YhwUVhK4BO5ikjymR65eOHh+ETrT+OVWYE65Y18U9h
okdf3LCOnYKSg0dI75XebKRJ9HvAThQWeOjG7Y60kyW2GmJBWMW4rPYfCwId4pGY
8fgqZlN+j5rJludz1XpowFOn0SgOA/TQv9qrXyvi4QPFT7U+uyJk8lawvXK4GsHi
Whd4R6czw3metZZNwxvNLWug+KA8a5vtd6XGK9U4hRD0A7rYW/m65YwU24npgOSa
PQ2pNzutmJ9U+QAbdIvcK40ZviK+NfZlqwNRMCZSriFKx6ePVCs8nTjdQAA7WyvB
qPABzQtgcAzH8HePa8w1xciPdOZAKZYMgp2wz3Jhq0OVIUUWkYBHLEdno3L2YaOm
emUOY4czC+9Awo0ACTXbBdN3qYvWZm/ixeMW2DdF6BtGYi6xUqUFe2E2nbK4PvgR
zaSWf0/IzU6BkXURKeBj6l+a1AVCIZqZstldbsLu3TWv4IJwbWzcvIawWaBReu4p
YWXCvik3zvLojM2Eryirjkl3quT7MXRa2AH5NHAzntYslyISd+4+ofngZT7fuxG7
EGHr2HzG9560YgZ0oPluQJpZWDkG+zaa2pc0671Vd+jBspa5sNMHlbZ/r0VLQZZ2
zVQXz+k3AZC7+xOrQdQ0Zrn59simZec8NacK7/7FF20LjPK4FVfCuyD9mvzfPnNG
GNOGh2oimbhINb7vVy2+2oTXb0VMUwvycxMZEvXyJ4efgyh1Pxu5Pwrqgs9FHrSq
6be6t3xoh7FdB5aZmaaeBfomtoH7sFJ3L1vTFFhax92Qn9YCn7aCFnpJDf9zbeuJ
dTsTPGeFPoGj1NTAdwo/FQv3JFjGqhqqKZ5gAmmHrCRMagkkAfQM0idkILW0g3Ix
ViDGeYFTsVuxX2aWSgtoU5Fsdo3F2v2LqfuolT4ZEqiN7aB6b4mgknl23n+GbSx8
w2lRw/bLAl4O+hdR9LWHaENIR8QlybxXpcfNCfXeq+DQMNwhCSby97lne36c08w7
TcrU+QEcJyvI0N2XuU/HjRrWojTQdGOFX0C1OiXKS6BSu9CHEQsiKpdOBHoADGjn
3DDYn6CloCmjGCegrKu7PQuWTgE15QWASw43+dr9LI0k7j3WF5VOTm3DgrtDQ3G9
VxMGNAaRZi0+bv7HiQfehdkLYAbeRWR+k/M/JTAkBEIQHI4U9zH+pkbjuD9Ovfnw
4DA66dhbwXAqDJA55xxrmWX1NOuILPz+OQ7skA1Xjfj3xL5R+/8y8wRnJ6KxkCIY
nExI9cGmVv9uGL/T0+V+2RNUw6uj9OvcObC42nP7AfKYVgLPYu05PDKLTHZJDYql
W0sErMyV9ozXWFE7XEyp7Q0urUqCQfRL8i23o4l9xGj+xRNdJdjeiS1Fgz4GWscD
dSjw2lpkOSb/lqcYTR1eJskHLDdweuxDINCNXws4ldkm3i6ZK0HaOOwoi9ShlYNq
AFkDwIuryvFYrWK4OjDNQiQP5JlMwqb3R0Q4b7sPETbzHDJo+CIhLKIohcueBxXH
4DLalsc7KPMEW+w5SFD2UZzj9nzt5mMq0TJAy26xTag3xMAq1EkCumc4QS18tfQz
hae+lNp9B5WaV7qiSCmtptd2FBXMLMC+ougYeO3OE+mX724z3GhgsDlxEvnWsCAq
8LCAzgvOEuA9llApPb77O7xudgD0twtml1wA18xmCuMROcAFpyy+yi0Y2g77lKtP
pu74N+NZUJWHFoHxb0Shib52NrMcV2kWy5QncjptwdV/8dI97swF+rx0BfhPYYOi
qKcuSt6AZR0CD2fhuf3h6n3AeNnJ6/bN6lkXqcQAEqI=
`protect END_PROTECTED
