`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCIqjTUFUFAa7onwEMMq0Fh6l62vniOtZxj5bnnOpWRCghIJGZKkNp0go9t3rAXW
zlMpbCwMT7PxMWjKjS6WhIMLmkA5BmPEAfi4aOxnM6SKXiEnYkN/DYudamOs5zJ1
jS2YjzfoTuNmy4UYtfeIANFtlDm6TeaUVNWrc3896ok9wcF3rXtGdMELlMmnzTxG
KZq/UIf/4u/c4tCeWz5Y0nlfKl2nhSUG2ObqHnmvnfFr+mjclO+7TUely2XN9YSg
XiqSw5KXF2oiKbGBtlZ4cHyuG0V/6iySQCjd1ZPPCqvBAhVD2aUfsInBZDn/4YYI
hGnoBc52h90o0Ma1mAQ1BSqlzhXzE0nQIsn3cJYRY7U4utIEE8cDEr3+eGfK9Xb+
aJfpPz0RlgFer5esBTyDnrhCxUGWWol+X/3//OyTz2+tYnZiEVvB2Kb/zhQq1XzT
RWlj1zj8ABkb8NPIXrfwbQ8islUwq26HuXO0HWwk78PyR/Bd0AchWj1y8IAtq7/w
`protect END_PROTECTED
