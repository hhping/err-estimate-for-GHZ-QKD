`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hm6UorcVq5EEGDTHZJdu35mqy7gC+bYN7qvmRHFvRNJm34q0Vf2D2E2KITc4+jV/
xwOsJtxOPCGq1PiVsQxXVzpKeHbZarFtO6C0dgYootLm6wvSkuLbyz5ahTIgIkmH
K6UP7eHqfsgJtVhGDsTmldwjq5kN5NK+zicgk3rgNg1jK56wBcYdvffUWWxzDRPZ
zvuMXHPgmxN1w+iHIwlbMfMYs5Osf0ztBFDffwH+7rHP7r3Cuu96Ps1oxBcDtZu/
kYxttj4qK458jL+CjwRBdIigIWiS7/afzPYrsPThppHtxqI/esQPmm/hOTnjYnDO
GifctiQaSh8M+sqmYZfmVubsV0sNjzP3HQOu8H4sJY8lyK8rzX4WNnBDJ1uBLT1S
MZKkPGw/dt7CQ2nkT3Y/R5G/4unBX9mAjlyIj4/I11UYOLUBgai/grAvHZRX7Y5f
mWmuXll2pYVMnDkdcd9AfYtMv+qdx7Qmorz7CsjysvMsa5i7etDqbdggQdSDAizt
k/STb3ucFU1W14a/HsOZf/oVlOgG1Xdd9YZk7Bq88hutZoxPllLjAxkkRnJmREsB
9PKNdJwZSQx3sT2QXKrQWM2MsVB+dt+zK92GgbPzRTCfW/pCPbLBTBqMmA2VBjil
gmPbm3L0mwHr+4kbopNEPAbHPePdIOH7t34og8vExvvH2GlcvhQFI8qYSMgt/z+4
m1wiMQ5AQ1mfm/3+/dGUG+/uftpvqgJzdbG2S0aXDTGP+vmuMYbzPh39PAhSHPgQ
e7VjBMUt+VmCCWl6QDfR0d+IBefRkAiWdvHRwcLttyILoBOxWqq/JnKZ2DhHPlfL
Ziy76sFYt/wSMBMDFadoHYULb9i6cxcyrFeNVws7pmB8u5Si8YFO21JE4uXTPpUb
8ndF1VRwfsng8Zv+BfGMqNeLJJTIs0C2XsVYJqNTr8EKMW3K+xLWz07Ne9pwSKkA
8Kg1VPnZz5iY/7viCXuFrcDWwbCl4ZycaXDR60U+ziQncOwMFtw76RWTrUznybju
qdu01CD5p6ka+yLZYLvvVV6JhDkOL2FNTg/Zy/LWpSPrnR5824AyP310szgWno1z
QZI2oPQueNrRQtX8CepKY8WDLF5QOR0ZAhfp0DyGOeObNG/KkyaEYjO9a8UZF+jM
IM++oEFaH6Sb3bGFQ/WcXzcPfE64PoOYw1z8eSIHnz88xmyY9t6xgFnwlQotQZik
mRy5/GWCShSGWyA+XSLgRXKL3khD6n5RiCUEOOpjxc/uWBMycNZZfvn1WWGcBGEn
niDciydc5bhbNxTt4fyT8aWJ1sZLwNNggSasLNRR7QUwO8uuTjlqmYt9FCi0E7/4
NLTRjkhIuA4w4A0xPWc7Wr34rg8QYioFz8dTakDqgR+Rm+FCGHmZr2J8/Way+Y0K
CUXX1/rUEhhDAwEPEyS77+YH/ZzESNg+v+3PIa3r8s5rF3sGa1XxvJOYWoXShsZ1
mYCzc6Se5R5+EyKRpCaS9vDcAq0QvAC09k6FAODCGGHbvNIXHQDDjI+33I7z1LxP
Q8NlbFlCdaPBQK+GEKpXq/M2Eg3+9F1KmoMakyosiNFuTa79+9VmovhWYQDDn+b3
89neQZEf/nLMDPJPHQHC++tFEvceNnWgc8HICG0UC2c/wGaXZsKheWDNKoPPjxgI
sLXKoYkhi0/H5vEXo6CcMwywDia4288U2Iq7se9DiwMKTx8f4LK82B7uFr2wCVC6
zU7+qAhHb3ycDhgMG8NM0CEauf0A2PxJuaA10eW+issEVtDxfkkO8KMBCn808bKY
84s4D3GinwEFx4vr9d5DmLzEFi1Cd03oALebg6a21MbEfj7thS1nyIV6dUwVBOH5
n4lcKvydvPnCf3u3qx6mrJLZhjdIQS06qVZw7HQN+Vxqwo4x3LNKNds2DuWkAQ7M
uQywLiIW/k14ZRU03av4gQ==
`protect END_PROTECTED
