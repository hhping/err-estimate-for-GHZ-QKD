`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kasAaBfteD82GXiOHVxWJ7XAnqPG2HAtPNQ7s6qLQUc41ZRoJAE3a72laPiEOvPM
AKgFM/gmIYkn0Q6BMsO+Kj2+fV5ACNH4v1SHvMKzLlQMPmOZIl4m2knc03l9UO9H
Ecu4os/9FMWRYI5oMz63PckajeSNpqEJ5IXFPZU1+KE4G8IKQVLoEVcVh5FAButD
MSW/Bazvmpua2fW9ALKubvxgRThYcjmzVU/1KsCgQVYkjEFLnx+wy0AynnQhAiC7
MyrHJMPh0ACFf99/EU0giPs0AILYGF61Hv5R4b2hQ9Xs2kYM/ody0c9KgP7azqJM
Hd0WMx77arekb+bSL8QfgsYbz5eqKLqr+eTeqlg8rNH0zB3I+mmPkhRZgWYJe6sT
X5A/GCbJLTyQm4ifgEG4qdA5DWrgaTVAAuALEpm5csa5atIBpmRamxXwLTeXdv0a
iHBn0EuXXUaOwff4Zq0iug==
`protect END_PROTECTED
