`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16c2Wmt8YAXtDd+WWu3+XEcmOg6HBJXNBylcthW3Wvw1tlkqvXCoIRYh24YAVL3c
zLRv1Ie0rihSOkI7mQg7VxjWk9MKQDD5zJTCcS+thILa/M3B8VNUXz1scV3WQ3Xc
YfYGeLEdZCnUM0LtZYbZLsv5hQFuoKcdjyUbe093oaYwAqpi3gxLrIOlbtwx2hud
I4vv97ELPJzOHF4xWYqQ9Aj6A/KlXMcDavbXUzVoVFnWkOuLFsTYpzu4KOYrX/pe
enx6hy5gblJh9LgPEotXPwAKyQkZp2FKYti0GIMluF9H3Zwl+sjjQ6glL8s4emyR
a5V4afnMdKc8Yu4v1PxxzPiNJSP1D69h3Eho1+fk8glSmC9a7sgwlWH1ykFkaSUG
+YirfB+zSnN4mzQb9BUf8GrPPG24nJonivSpB3mqJj554kVHhRv/LYBh1FM/lgov
YfIfeh/4QU9iWkYRGNjcSbjq0UYKOhks7ADXh9wxUYwJWVlJ468pKBUcrfXoK286
YxyJJi9UnKZ5KbR9kqC1ZjClU0Wnr6OL8YHfUuUhyg+qm2EDdtCA25SbIm1tB3l3
Z1dEQ0/4FA7x4b2/PFkFgPIwZhVnn/nWyumpayJxSbfdyYMIxNenFo6ALKCmKGAI
BHr4oAAHmiWv2V4JXXVVNMeFX9JC8JS4LCd0czv7IJ/pWFBjVLmp/aUEwtMv9Rph
udAl970iZV0pBzfrYMPkvKHkouySlmpLCv8ArsUKmeLtfJPY+2wQ4xt7YWEm4fDf
tQ5UoqzZnltOkv7wbuNV2AfqzwKzIqI/M7k5ilbL4R6H0YI9QJdxlBjbX+P0R51s
49a8TnROqX6QR515C3BXuj57An7eNsxxABO53yH+LteESdQm5he6ZYHuGgSDM1ON
AdendxpfKyrTpsgXzUpfqSkoaPadinR73U2InAK8Mmec67iK/fd5BlDLI0HCmUGa
5zbQjww8ok7JMb08DSbmVlEmyrb2wcJB54dsa2Pt+S5KqEkzuWlw7kCm4z/VtTIA
7rj3zMyjhw/eH/2+xd7NozP2MoXpEExRpqTtT02/AHNN0LBTxsaPyAUl8QC2Dqlq
H9d9YqzaECDIj+H79cMbDVT3g1SSHUY1YkFAtFmWHfpLRlTRc3+qkSXDP6vJCWG1
S9LKHKk0jDt9XROfTRJflXRWsb4IZYOslx9/+DuOgbdTswF4u/7paZu3MOPxDLhJ
Y1rWboziM7m8sQDZK3Ij7T/BZnzqADEvfZZM8rLxfSUtZCI6ZZomZRSWzoUFxOL7
f/NGfGBzZ8aNEq6wHP13kzNTEeBU9EJ8q9ixt3wcbfOh+T8jOUYOT1mgjPfMEr/Y
ajQLeDSleoc6i1Y2mHh3rdePXYgXXv1rmdwh52yQWXemRPR8xXeuQhEsGV20MFE3
C36/sBcTDdbbNPWGuS/5AxtUANjJONSwPqIWz92KZ+1U3W9sevG2iGHNnudjovqv
Fqv1g17aekxRzCrXin+nIhGZzt1aCIem/E4gCiCh0dPacZtfHkxjX5pEe+diYQP6
`protect END_PROTECTED
