`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsLWNpFGnL4l0ChWtwQ7uN/p9L3V2zFtYaqHXsC2u/IDo09ht5MtQI+9Ti/vKJH4
7LxE25ANLX2p7iQjR4TOKnzU04KU/5UrCHQQonp4PEP4cMxor8Gql5X8SA3yremL
bsz7orUbqVXaD+YK8oVe5ZDU7iJcVVYl7jNcLFUU3EB0YJx7rmHIUZLMXuXnJB1B
f95+4xZQMPyL2sEs9hBdK7iA7lvzxRAdw3QqgrRgirGd4ppNIvNn7u3O0K2KVdKH
gxZMVJKoPasSbUVMwtJF0ZB9pnyLOV+piNeOeYJBJBUZq+eTs0Q0fWUmuOV1kkru
wrHQGLpY/CKzF/AlnCe98seu/r4JSx2c+DRDpChydKPG4TAB6Vi3zPgk9/pouQ5l
FeuGMjmT4U0qU7gjJD2j4XKzuywnA18CBWhjMPfSZ0xgq8tderFGNi/OiCOtxdxC
pSso8+ttH/F/m2CGrz2jxmDioA/UgKdHkLEgM7eCJ6mf9LGLta6MYXbHhiC4mQpp
aVW+eEmWBT4kWSqw7Xe5q8FroFKqeVHR5vSxc2EYzWRDYpALLXLg+q/zMDNwuTGn
BsL4zlCzmby8c8YK5IrnOwKv3Kj+/WCqJFVHe3jrlJc/2c+3vJaHt9tnDHxj2wR6
79QPwEota7LmR6LTt0q4snt3W8Hg/ej5Luim2WSvibim8noNm/RStthx54h1voiW
BwajcsNgJR/0xFF/emElCxcHqCagQP+lb9OJZHRzI/IUKm1Jb9Eug6uapPS1+npY
YmsqgEeF5rd4asxxawIQjEjK/BNhpJTdlfLOV6OVpl8H1f3VRFkExtYDaVphwKPj
YkUluSxJWgW5KqJr+Pp9Bc+T8VRA8BqEtMHWb+zfSc1Hnjpc0wTA3SIrsEwk2EdB
sjMltJAIOTKUPyY3tZ10aOU9JZ0DT/YOG9frJFkQC7TeGEEHjQoq1RHHTDg0ZRox
c7bRBfkarX3FUHWk/nfnPevdDrVsWi6qXpAAZ2H+N4ca1g69Bs2CL2tJQ+pd6tlT
z4E4fb043ho0Fr71TL5wzyt8Qo7QYzwG1b24yoJKgpEmabiDpfKnPdnOq7mOykzC
zwL+dIRaljUZXFFNFT9diuVOdb4CRLM74tzyz0AO7rZyVrxbN21VEKXhFE6AiSOp
aLvg0Uhp6+IWpLEXx2EVc6CSr6OYVzGqCo+vWPATNYUzj/hnnluF3cek0nAgHl+m
q9oNe8tgGeNyif0M86zLTE2bSnASW/l378h2FBdkZ1gcnWRKdKAszQJwIV3R7z+L
9HEWy9y4o9ovfDFBN8JFdmFV2lNWg9ZAtW9cs0W2K82C1w+/c9RfCtrZtw3cHmzv
j6oDlTCEzaW5783cujvgcb5dagqQVZ6carOKOrVtij/wH9Eg6QD8x3BvUSqbPDsn
IR37+SkBsm2ciRCVmPP3deZUeup5AD0vtP0IVrt0pII6uah9pe0Kwh9Cz3KAdxtb
ELm3tilOg1xArKlHR3EqX8cQnEOnA3JGhQWvPoBQUqcZaXbRFA/IoDhfAnh0eI/u
lL1VyLouLc3MoeGuEFink9hHaNw0DTxQpsr3bHQhvCdpsnzOBv2C2xLreuwLt8ON
HJHKNudxgWwI5oE+8cSkm5KQfa/6D5J00WuGNV1uoWax0j6jA7gGc31SxvGTvRGG
syzpquGzj3hQ0mL9dKeTsk31cRIKgtqipJx7JMIO5J7ockP3DthM+BFahubkXkHy
DEhiaEl0L/EnI8Ie1NW2kBIMMy0XDHI7Un1aIV1v0PGgvKhelVYFypDXQJGWf3wi
LEa9MPDN913PcaL0OF2qqlEtEsL8pSeF+8wRHWgisYG5zu/isklDd1saaVjbeX/X
S46qa4bFGYwrVhxvPkuzRxANalNWJmaCsvHOa7lr5XMBFANpcNrdlYATUeVaff17
1vA0b24enBlNhH0wY8HWP+l+FTbd4Lgcx4DI0gSgniFMGh/PcYgna5yWeJ4ABjVW
1+cR8aTpuG+wqPxCUMAMbtaFtzHw5vs1RZge/WPZIlF/t7NlOaUmCJ+VaWQ74qV5
D6GJw/57AQH1jd0xvtXyZZPkzcx3EHjaxshkLiN0cujwDnkmfJgWfBg+HDnZVZvv
vaZWEE/oWIgGULdLycLMLzMLVC7FLgyoa5+AY3JnbCJP5FjtPPiZ74tcHPEecLJw
qVuQ1+NjJ1uqKvVWI1u7AF1Jko59uxNfLcsWLt3GncX2FeEcmKF7t4LJoThc3x1S
kCynCEi9//bMs9nFKX7E6UrzTX/hPvHLWYlbgnXGFBNEShnrLhxCDHkNrlpGmX2J
7JwUUB2DzCrDB9mVLH6EmBbSq9kL7VwKZMrHxd5iKB8coMY51I/xX2P8uJLGpitx
+vIwmEWQWpn8vAJ1REiNj01eU7+vKUiTQrlz1tQCbcb0zSip01QWUgVdxIknu5mI
74jTme3Pw+93VvsSG51vj7aYlPTdipNeEJRF3BWCu0ZlRqhtP2688SNx7BDGTZuA
cJ39oxxF4vjSHYsWk6tcJAvi7IqWztXxqqyVQcGOuoxOGevgncJ2gKBXhliTAd+K
Y7Y9/fdxb4PNrVZykklW8Y2ZnmD2ymovhpphBwgvFbBx0ybHhX/0Rb+N1nK0KMiK
v3uL1nAa7v5ue8hcoNJua0O4VgeNAymTWc3RkJrMZXya89338N4d5d0qsca9TA/8
Zh8wVXaxIhFHCO0BL6wyrP3eAaa31QZ3zblg5xfbSkTy0atPq1Bk+2NzEL34Cm8e
uLX6NJHKxFrGuwk3NihFr2vTmz39k9NCswjXRN5YnwbvxfLeLOGXnK6Zuq14N8dp
OXkZVo7FEnkQIXMuavxXk2naYQSuImYFaFkPh1xVcH6ue0pkAm+E7MhX/b3OCjH/
TYTZH98qsgkQdI6fcjbRlFLVqTxpGYNKIA+2YlokAkQmWuQYfhzJHFw9wODNj3mj
qwF9EiSsVNq/LlMgF70gu+JdDc2jksGnQqiZv0/NLmaWiQZWB6/4Htk27hDWtsRH
iRDEGdab87ItzMRNnFR/t0NlIbRyPlMPSwybYesl3GeJxcCC8h/NXUWCsxEp88/F
Q/a7DFg58K1KJwiJpQZ8gNpScGD6NVz/q3Q9UT36tgQzrIXUIxxATR8t3TgzUUo6
sxYZ793fdWc6XgqIqdn9sVd48PQLxKmRy13SVuSs4tdMAIDDjtpvVqgeMwgsMUEs
D2AOKRC1wdnNTnOrKPCJmD5m2GZAtksfOXlL0B1KbNWItcayUKddD4Vvt1g+yO2N
sf2Wgs8SYGdZRLfluJWN0T8X8QQSYARvPViMpAe6tuq+VgjjN8hX3SBCdTC380xe
uAttmUce8ey2HvZod4VkWSIsdhxmXYPPtXKQva3HIUY/wIHczc0sE+oXPmOqUZB0
/RB6KYvevJ5VUTbwnmHfD4yaKOFNlMOsk5VTpJIXLJyzgfaBiy3twwZab1WduPe8
Q//BYF+mWAOdD0paqFaWTVdSbtSU5leeRvAesAjLn5P2OL6x6XXwTwSylq8jzqaD
PKHkTlJpUSkgZnA4XT1VoX1wW4H2bxmpDOKRcbgpvAU76/esDZ5Qeu48n1rBb4aI
8MnQgUxVnXK338W14/ryJ+3B1vDa0cVE5aSuP6SPNqlifsMdGy2Gd0a1QDNQ/RaL
MNTGK6rgAoyXHJoUBasn1BRHsK5qIVp1oDhEDH6qe/Pb2gxve4LHZVHC/i9zmZPP
Iuj4ouZQfg1d649UlL9pSO9eS82H4uTLqD+M64svB+I57uejl1zzjyymH8SoLLGD
sXhzp4FazchkkQo+EhLH4IDS55dAFn/05Ra4npz13exMGJqIcmzc93szCB8nj7rw
dKTAA397dv12/26uZHTgRBWNXZsZe7nnvYAploJkmuZ9oH5FANelErZfoP7K9Zlg
tDhq2/5fthWoCRaY/xJsuXomOUobMxKr0G4cvVJeKk/F/C9eNXVEr5Vxe0wtm1KV
vPzV4jWDiB2aJrWKOmGW2DUQjcqPVqBre7Xk5szT/mcbBx8GiNUG/n8k6AsRFEny
nVZoqM6NA/r2qhnMBv8jtMjemGEjGL2M8I+Oj01HsyaEMJ3JuFdH9jwNGzEA4I3Y
NUyCaEXrsnnSh9O0wKq7ruSaCS6cmmpSxjt0KccAglk3qlrTsdZK/LqKG3DIkFHy
N9tG45+2NTTVXz0dCNT5H1XS2aIcoZCn/z8IZ6nOFwl50I0f85RV/Q2/nusl0qlo
Dq1Fl0h87OD4yrYUBXi4BahDkqd1F02ukXYp1vIJspd5mcTQZI530Sg13p/MSLV/
STQ3N5pcAr7iD1YrNkCnX9vSXMis572KdOyFGmPNrJYu2B02ZMODcJZ/DG+Xf+uP
06gXO0gaEUvSePn32j4Wy773iERBXt03VEAnlLwGXKw=
`protect END_PROTECTED
