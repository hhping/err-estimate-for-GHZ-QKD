`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DCf+mq9q20WQvS5cFLxVFY9zVcDaWR6tEV73IZ80TjJY6f/mEpD00gTRx8H491PJ
S2Bb25goRhXum+WYRhblL4fXUh0gm1DqcpBFz+jT3ubLJygSSC0eMjRSs/pD2hHU
OpIXJ2D6vwHNxjPSGErOqErUTCk/PEBYE3jQp0CQ8F7uedeBhehT1jIyFESukA7s
yMnmAmbP4cn3jZiprlyVOK68HUbCBYeSFYAQVVJ3+C3es15z93TjtAxcDjxaLgVQ
BB94cC7Jks9Lx/BmYad+hdtSyet6ACtyFTVRgFsdBv5WOroCdHpFOcdBOFYBwdDs
vLL27UfaQ/GvGu8D/2ufYuLNT0/Go9QCHZts3VGNh1+mDgARVUBmGIuQPMFPI84V
CdVppzc1DyvQEOIVgbr3GZmeAroUfooxptKkMhHKXkBFyhyJUVUtiIRceA6E7gx7
0jZmbemgYPnRH56D0LiTag==
`protect END_PROTECTED
