`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQ2zsR5KWilTpaHnVSqkZUWWrOMTHtXQMR5dQFVlThDpyBRIP119jfuBkVCXLBVc
6lRGuq/MaLgJlB7MN0JxRZ5uMmn1HwGh0ssaK5fISsQPnB46AjA923oxdlKOUl+r
bfHwX66Q2RwPy2Oy5SmZ7iVYHCdOAHwPSFCh6Vok312rY+LqmhS/9tn+N4u42J7H
ff9vumiD+ISfYs1hIigOc4N1wwmYIxz8FJ/uQW/3q9WkW6nq3D0d7EebH//J5TAH
qNCbRhPScP4GrjLPc+eo7N3xdrBcnNqhBMK/Dllu7MwgwFZVbW7d7znyza1TkABv
o2TMNw9XnxJi5NhL4cJS6aLxfzie5odJlka4a/kTGa7V2ZjCajF0RrFqoVOlggQf
2IeKzQZWOuBRjqvBKHsxcVr5fxGHBnVfM8le9S3MgIwfVInysbEb0wZdl5qkPxdF
vH5jo+JIMqGZ2DT7QKaQ56iFIaHL5FjRPNFiOuWWgtX+c9MsWWDQ4pxmeVnunVIA
e4/M2Nnze0vW7mJcsL+a48lyN4xlB7dtqUwi9zyZpcbojWbgE8hVteGuyUzbLDb7
GuBOfAUDladYSHOgyvdzRL7QSYu//OevdzilMiZsnGEapwn7b3ovM6/GyyXChoth
/z24JF3VE8P36Ds6TJe2FJFRwb0xRrbQ8iCBKxQ3dR3YYAxQigOnUMryC6uESCIw
Kfv0hv89TxONyDa8q7Mb9t06O2hjbc6RVr1Kg5M7NubqYgXwecGSUUlgXKBk/pXP
JFkfksGQlao3Q5wfMErgjop6czhTVNWw+oZSruagH5aq7nOwflTiXsine8ljLeGq
nhMlo30+YfhOAMyRz/6DM4AfKy9ISvBjAKzT12ZGjvlbefJt0jqTFEHNezrjokVl
CJDjcgnyrWtQY7l1tisoh16go/j6DdCB0wsaQ+n1gSx+fbcbJ+hGpHnRUEbWJDYG
tSJ/geabK6iE4JJA8TdxdTOoGBlq+w3b+PNT9l8b7DChHKVCQwEzex+XC2PXW3pG
bGm/+cPlDw8sgQR37WdOGmPPn8myc4R2NpmyCXnDlyc2WdTB1jdPgRMuNCjL304o
4DbgyS1F10n1BXQx/eOAZmlC0HryiMohQ0QLQxxzS2/6huaZKjxjQ5OAGhFJYh9v
ZMjOYihrVM7HAN6Mvzl7ved1z97DCoY+6zP5AGOOlL5W1kOBtbJSFXffR1XH0Eqs
F360iSGDQKQ8K83ReAIJhuohn+6E95IoArXRPQGTOCCs6FZvgfnaZJQUnOsbhphs
A70LKKEewir6psd07voF3x//T6SYOreEGCGBhPjYIbFMRDzLiB4xJk3ofXWuTlCa
8iZxq9T8oNswUyFjKVnFajpTCga5vUfzx/KLLDLuRLIgMlVT9mgqxLzkOCNN/CcF
9yrqa3X5dQbirdRHumhid6s+ula8eqUf47NQs0Yfs+yUcAZU8l30neA5WeIFs9jM
klsgQxec4ht6sqZqkrePHkX+LnvHY+qfaHxPiYaOLsxJiN6N68olEHQmeodsYd5X
Ipcuy9Fxq05SF+oDNTWTP+v6J8HQIeV5nzEb8jqvtizvRuN0gcTVI8HJIpR4OwlZ
ALHaN5nK7RK4R5eL32MpkxoXnaILD18lL0okXx3hgBfQIXllbDiAJAl2tvE65S+J
NVSpoCu8XlX3X1sv0pSTbUk2D5zwVO46Wdz/bDlI7gcX2ChXg7E0H0pkroW71YjJ
c0TSOew2zG5EvdkhBl4zQdqKBE5ieXijywNFxfLGuynEaNI6N5FxJO+8WeQcKxs7
lBqFvvDtUufGJamm1X+L9M2ZDqvGrYwGqinOTNo23cS85/S/z4WRvCf6qpq1yFtx
/IPZoQdKLpuTHhG1uj39hgPnNbs1KR7/RU48QdK2I388uQUl48Vu8Dy1ZAQ/FwaJ
rncF8vwRBaISTry7SXevRINnGUHoRaXqLoVbpGNhK1vbi2NikEaDwn3LZV5VyHsg
8oagf9qZqJ2tkHM9aZZlI4YoqdU8WpGoDIOpJHskthcqzm6AFo4VmWXtTq+bxVA3
ZNLW4cgxgYtSEwYhF3DJLqRu5mC3seUitz6WBu1hs3zZEUxcOS+iOs+Kip8fVby0
x3MeZL9NcHo+YBer7s8jupKx0f7kvY3Vifor4pc+6WP6r487QJ2V4LHICOMV5yEy
6ys4sery8qAkbr0M7MVKz+5iKj8WL2tbrTx2wd9IpOiVEQKFNltOLciswnRbvi1F
1Dm58MD9X9nfBsiONV1V7DJNajDBXsNE0R5MdVLtAhg2MnN2OMN+rj4fWuFZmKAO
SVW9gEZ8FfR9QDvrte+LHnT6/mIk062Ua+YCSmjtkOAyumCczJXNBQYRa2ZRulOg
wM7UyyMVnTIh1ODZi2WRpjFfOGzSzggzCTCbfZfLAN2x3TMCTeF3LThOAz4Uz5He
bj8zFUUWndA7MUQznK3n52+ZMdWNYFxm2BbhD0PH/CEMcu91IgFnK74+9Nsqs+oc
U180Gq2ITiWLZdH/De0GBgksS2Mf81LU44aPniwZn1tIuofHFco54KBY2rVD7n+6
SELs880l8y++EW2mLAXKRrg6SHvh6ce5J10JBE1UIr/PpUP4SW8YYsSGy8JRjCsJ
eSo3cQCIIzOkUPw3z7ydMaBYaNwNu27hLC4DBp0WpxJkmClufswrLlscpY0DZs3O
Y71hWeH/qXXO4VDXtC5IjDU1HWTJnI87vgIPZRsMyQuRak4Rs/IzvfwQ0CZaI9HR
HBktVrcMSz7hHxUgOT+XylRu6VNhgZtBtCTfUEvpilUDlNJMawMAXSg37xzoLZFr
IM9VFLo1X3pU92z0vD6X/khE2ZvoUDVo5x+8KUe38bOwInpJDDd87FdRaQFjPxp9
LoRv+hQqY01kZ7aHmZ6tR6OYU+h2PPK3doSx6/Jetzb2ErtriIJrFixHIbNQklHR
/eqxHTxBes96AD8itmL8QcoDFgVuFlHNt6KhF2ctkp5XeoRltFm7aKaQhhnEUlM/
k7KJG8vHxIH/oaUjP6oKpVOTjYjkXEGuyKmL0pZPF9n+8goAa74li1tCtsOHnBLV
YEqO2cfSzj1fVu1o641mz8VpiOpps6E6mW2QIreNi9PHpIYVG7gMEHA/jeQItQpb
gnbH6rCKC08ujh85MvZf9h6j/WtnLEZh9ccqzhFiOIhR55WJ0vyazDEqthHMIHtN
5pbm6Ws7hep4UIKQ+MEs6QFlKMEbs7Og2TmQnattYH/7GNNwYXF98avT3IVEP5vx
XmI90MUoI2Wef9pL2et8enFHKLxK6TkUDUMbbq4pVQevNlzeCw/O5h3ZOLRYDh0X
srxsw25o4PGfQ/SOTh7Bc+Asn1/Im+H/BceGeJ4S/2j9UVYNQPx7Qi7jOfg6fIuW
voBW7Mss2/aGhAXAvUFg1tOoiOPjfZJJPi7Tj5+nppQuNyiReWSFvocTnwn7LNuR
zBzUMlrp5hiEgTaJDO6ui9miYAtGRxJhC5RyTSuYYV96IyJ73Zgt0FAjQNLvZT2h
6DNeoojpjLCnIOUDqX9tSIqSvaLdmQIiN1NWhJaz3MyvizT/bd7x/q+8XpdXmsmZ
gtq3hbnIy3zO3Xb10ZdMrjeDdg8fkhcDIyuWrm4R98OOxMuCb6IfgIQSDKlkRV2P
5z9TFcoZdJ8ZC/anPqq81ACyH6eJBoR6pfOZfzwDYEs2hZHCOMEx0KsLBSiHdRIt
Fxi69lqR5jFiTF4kX2bS7q84PARAkKMAIajMZV/B3Ts5MBEQNhDqDiy+gs01v2Rf
KOeJQkC8plF3ug2mG09w1OJFHYnv30NsuTuzV8jiqPArXKgDswP91x+J+DRLyxVD
colFmH9FRg+KVl24XrJBOdHrx70gGY9+tlnswBxfJHmPrsKUzh08V1QNdtkiucF8
R8AMj9awMlo5/7j+x9rk0KGWnXR+v6CuXOsRbqpzZsVw3L01y7JeqkOpGLxiGpNK
uW14vfs6TlOZ733ZNZBOi7468yovRJSkGWBprAYhSsTCK7qo2+3CQ2F+95fA+yLd
d+G9vXfILufLZWFm4KYNG+MhEeOkArKW/5lkhhZGRhnafn+T5dp8MliIua7IFuy9
lR1a8tNMf+6p2F2c+DkXTGsUlze5bvyd4rpnADnwczzD9kdnimK9HArz6nMv6H/D
2HoAcMgAMI7bqXT1g7WsbbasGoHeElaH4pjq9SIImVpWlPAmY+996ABkkbX0QtF6
SwRC1HrqM380A2BdIrsS6SIgG5amLH3SCIztrcI6y3GYKD58kO8VDavar3ELPVfr
/hzCt4jT2svlpRA1ul+OxSKNn246iLEumcetI5hVQEqzxLhF0o4gXdYmB/zOqmES
2rQ9CI8+uR6wIwPY/b9/jSIibxecsuHf/IoWKuHJQgxRzQf0jOWzkxU9YQfeToDk
Buc1Bomp5VGdybhA8HL7niNsPiXR00v36bDM76d3QzqfrIyyD/wFNmGhaLRCZ/lk
Y7k+hmHip8kAy22AProRievHHKqaHZBew5UmjguoIU1RfwpI19k4WUwyHMCAVFGy
bbw8xYkZ3MLfhZZS0J2SIdVtRzNLQL1ngQud9JdFsvqQ6wtdHu8p+7kwS3o2iT4m
6MTInXUMaocnaSfGbcnl+moXukpBZjznT3V0hi5vbPNNSJoDigzO3rVEQ+fg/JEQ
at4cRAx/VnA33bE6QavVEE0Qq9pTXag4ylEZ/sT6hwikGK33k+Wt8JUd++oW7eIT
2ulez7eqkdNwbEUZ7UUvndpi2CwNJCSjltE6TtJcEHGuAV1wgiPGTkpadKvYBQNB
3s/3zm6xVtJgPdewg8KnFeK73zVxphx1/upktAfkov+rWQYr/yI3FySzWE0Un6W8
OdItkMzZIBG/ea5LrPmYGA4+o4oTzWlK0c0O+Y2qcbKar7cQVB6C8U5n0S64q28Q
nfnjjjBsaAJVwoqH49JNgAzGepmCtkvkWUeOm0yXoWSiuWxuqVgFGXrTXvN66EGI
sr4KR+mkZbA7I0P5uasKM8KL6WDwrkLWDEZys+qPNNyNB9gh/TOkdI+P244sJiUJ
5ggc99zN1xS4/IBtnqvC92e7KKgDqbDmkPSvaVEmXqL5781sR4XLVE7CWegBTjo+
T5pFxY/oI5M5oywzz2hbS/4v1x/aGwcxTIHx+t6sQbqJp7K2lYw1AaOALMk5Dx4j
shU4OboOF9osnboK3a7FfvoH8N9HLzvRCHT0lAKHp3G+txpsnBFVAbcr0ww5qKEX
o79OBouPjgRhOAubwUBDyNWnCWzb9ZFUW/eFF2GtKpAaIfRUpBaWN35yTtWUlUrA
dXnzyVfE2dXRMBTa7lpNLN0MTb4yHFfF995KafoFT5kqB9x6eFHL6BSj6f5zIFqQ
2TZ909q+eX6I15APfCXQgUrQC+DMz1mh/stFF3RvI6rJjER+11IuPQ82u5xA2Qln
g71CDbikkg6dCb00IH8uUbK6xSz3ivgkFVnZCiJjMV72zGOC42YUJ1ZQoWAfEuUE
tdFNGxvPqJGEn4HXEg5QX0t0jwjwXPWf/xqTI7BvOnP43sCg7JAj3P0NJ/XDis+o
nCnl2Olvh8RcuaQDI4wsufqCLaa/02wSkYnA7BPOkmGwyCCt1afUGkK61Ojm0rbQ
Nyxa1xGZMRCgDd3Ga+vHtmbwCHrbU3/lIfV7rPuL52R1KeNZq0mqq88//73l1PNu
qYfT46DbUlbVQGTRXz6pqEmrdNDO1+GtOwYU/UAhb6Ex9YLxVBmYe08jp9aMJYbm
3Sy2IrPBXgFldf1jAjkNs7XUo0XA1pnIJkhDKxM81l8iHGYpDS0HTCtvJjBIz0ot
Hdcf2L20PNiVVaQPorcgMYrYcgVIU9EpThhTxlwpKFpUZeooTaxLu8tTLGhsYr8n
v+JyQZ3cD4ZEibHhKiABSVsvFe4S3dUXfquDV/L+S+p4ZKL9UN+tZxs6e6Aotlst
H3Q41YfUcAS4yx1rYGbs4yhhZZ1h0sGpCPREk8OGdakTE9flDNSJm2rsFkYHguVm
fWwZetfoVqD7P7KoaXE0MREJH+F6euzBoEIvl5s8czbHrqc7NakoyaH7eXh90AGn
a9NaX+G8sSQzArqwDMYN1RVumxRxZVhO4CLXgiGEHZ5DT8sZ2IOmWC4Xz1Csacto
0tF5zuJiTv3O2geteFiVE5MaKmzzgQreZLMvRrQd3+TTPFU64viF/gTXp+rE4WYK
xwedF8VPTXhD8caRkZ5sC6QGLepunZpXVCVQpEglZKhZsJ+Fx96vLJGStADlWrJ3
wlzg1sln3I3wqEfKFYMkpwy2SjEAjkTnlIdmesrYCPT9NLtqz3FQBsEooT80vkBI
ECGFEuZVaYvJMp5SSaOTdwZagSuXyvbKmpZmvTcmLb2uosk/O2Dbd5V74YlGid08
s5BHUURwGGmtZKjYX495BOpFoBFITGHPuMCCDgEowRHTCGj4ojQb7BwMtgrK3OrN
Ms/QJTyFHb9gfQ/RBMbsmwBf8lWhcT5kPfzy7qnH6LZJRfwC9hv7p94KvzEuN38K
kOEPGciA+O9lK3hoIKXSyrAqgjavp1IlHyA59bL830IDyPmOWba8PpkBv8kILqBe
1PqQQykISCqSq+Qea5bvQgWjev2pvZI3XrUIREaSYkvIctsPCraRidPvnKiqicK/
zvDF1MJjamdibXHw2xl0xlkm5jU/WFMMCIy6u94afRJ7FBFAjFm5mcmBvjwPwnhZ
k3gsftr6x6Ac8EjYFQlT/lnKNbVCBZ1nHcfdAHIyNagK+4zFRGkVlqus7nLJTmGP
u2E3As4n1n3dZ+UTf3YVyZlenEgyAjOWl6DwNmQQhHYho38EFuKU4D7BiyBVEl5Y
sMODjJvUYVUm5PvyzR617ZiU4MZK1S4YlPnchT1Eq06/uJfpX+s4sbnS1wzmyw/c
HEGi6v5FwHlXJDcsQeENvEry2akgXBRkEIpynikXuQqHPeYKIYDrVwQZhZEStc3R
B/VKuROUXAaGuOsfCMzw5XmCMfet30+MFpifZ6JabtgI3l+NWz3+ublAG+K/2e0/
DBa7sUXHL110VN2pSXAuXr/JYDrjM8pukTkgrpTSjNWr3o7OwcdtyCW6KsbzCj+4
5ljosq0YzQ0aFcjIC7gxVZxmqghB3XknAxjqK3z70/zdsLKJplLBgn1lhVTMwg48
JQblKEMvKiJsXg6FuUj+ZO6h0d+aDo9Ni5ft46XaOBNqmFNhnyXX7RpN9OrJJpWL
RoyKvTW9wuwInpAg6lzBvaHIv+99mq3Yq1gsuhbsaUXG+kuj0XV9lS9LhP7pTEWf
b/GxDBnceUVTI0fo4sYTRiekL7i+s/Uyi96IoXw3Vi64rn2THV9nfiFGRGzVeTmf
GXOJfut/TuDSGGWWC8U4Dz+mBh1O5MgIsp8oBu0fawt75aDslBZpdasrtAaAFSmB
lNzCXQDjq2ctWrTpEm8mQw10T/gxKKhOw9JGdqWR4UDj1VWK/sOOwlxPE5m9n2E5
9562LhFnrgA+Fl9id44ClfvHHbp6/sEGahKBmd1/46Nnh8mctpKvxVtkBdwfeuoJ
ROpKLNQB76l5jZXpamhGbq028kYl6hZOBvENDvozaZgUBFc3TlSux5kfV9YzfYGm
MWnL2zBF7FCKm9rWviQYeVlWOJNNNUe0GiMzxRLp4EoVzVTdUNW6nlDDJNF2pMtq
Dwt/3lTAZjyErUVZoOYJxft+mYFszwVRBMns1aq3cWEAGwSTi0ZU2hVn2g0qpmtH
GpY5kU9tFoiPxH6qF7s17weg7k5bAjIC0zekojw2AACmxZW8lbVG2Lj16veUzeYM
SK58GN32XGVfxfnsDYXNmEB4nRQnNCQUcxB9lLPNECRckvhi4Zf8oT282s51qHq1
GCD7zykWpNYpKuV2bsqgd07has8jg+ayZKvTUuAAYjo+HRBQe2qF6npK14rlOxdi
4j2YhzXw2Q36IE6py4SK0F28oJQJBJ6jRAnNi3VeIA9nXPuerp2AIthCAkUvoHQJ
nnl3+noOGWCU8ruPZUIHBG2mcGnyzCqfpfylEe/HEbbSdKCZus64+Mdroff9HR0n
m3p9AdKj5y6qBRDl4f4NQi5B+6I5qRLt0PaT9fkSs55gvufJeVDOt2szixt4I1nL
tLzGUDlW/oa3R+/nwfwZbSWJntRVomeSr+urDD3SlD+hND4Nboo6n7uEoY9CXGVe
bHjgmWptyIZh+OhH0cl9d0+5W573lxafRXIbOkA7Zs0Tdfj6gIbIIe33V7CVAhrt
4U5zaN9qmhc1Dtg/vnJ1526J/snAMrqA2xIqpOE0oM01CWHJwNY/4bj/D3bQmV8O
xnLET4K4cxJ1V/7K7dovQAidPoZj6QSB6eWqY1iDC7oxThLbFEBoEN6IEvtkkhp+
CuRPl2kZUI1NA6A6T2FHZPr4f9OSF2SVNV9OSUyABndOt8ew05HA2CIv7kHqoznV
UeGqj+epx2pEVwZqR+TYBLc0Dg9elB3d1VzD+LRl9uuo5V6KaxzOuFLljzGXgEB/
50ScGkFUIITF5JEsFnZjqEEhkLXTEXgTLhdqhGTorCf39ueCQhPg3q6ztcl7abln
08AqXrLbv2rN2/mPi85yynbaa34SFDYKnxEuYBcGHffywW1lBQ3J+VpEx5K47RoQ
au6wNoojB6y4gq2TymD6MCGtwFGii183uSnuhow+vR6LVIjQgspUNxFMymNkmPzc
mqSY3JvwcHPYxg6OgY1Lf2xNTNS2BmwmoXvoXWZgAj9sMWpTvZ1BLA7CkDhh+9A4
KFRIRP3i0TFqC+i7IWw3sPqKBwwI8mHhXPtIJbjX2MNyzSKxqhp9nkDJfR0/og1P
QHfxT5e1bhpUNWWfTApKY0+WiA2hnor4zk4uU2LFhOOIdSo6gG7xWag6pXG522BA
5PFpMP9U7/jQpkOy/nlxXcKx0Jwi9bcATVqiGKTi93I1UBlc6Qo6fUAu62+MreIQ
Q2yqjocltQ/wNrXnRLTWCWM7svAOeQQWIDAIO8IZnG64gCnvUjEkOIix5/j4SUJu
Dk9BFoG736i+juR4exv02htTkwNe1jOciQov2ZbGI1KOpbekCdtZrz3Fu7+DQWiQ
7HW2CrUEE+FPv782qsZLyfjhWaiMDEBj2ztds4DLffKd63NEty6J2VxUPhi/O+wj
FF4uCVoVxA053oEoAehT4To/55l5rIhcYDjMal2hKlzB80XKc5SCdffk6QAIXrXf
g9WYLHU8IAniHL3a4/bRhPJ/BSSJnSksvtC31r9aVMxoP7m/ezuZraA/VhfrDnmp
i6SAscTutSIseFJ6kUysmxpMOEzoW1u4Snk4LzBM34+O+QA4utgX2hBkymz/4/Ep
YHNp451LEC6ew2QK/RxNJ7jbWlPk3ulirciHKrr9JVZQ1IiRpUBX4BFXZnQRyJMg
eNvltzYR6/U5H+33XamcQV3bYrd+KxysXakG1+IuN69yfkpDPsVgmeM3UN5xfqrZ
gG/KakhkCg1DmZ6YjkEKpFvp85c9qbdiGv0y5H9ASHjY8gwe0ve5B7eekudjRF9r
JVRpSNfgg+Su2wQLry6Mw8btizTVWMGhU5ziggoz5MKE9oAGy3MBJyUqonipNyYv
kpMnZXZL17XoRt+m7uwJ5ROvQpVFc/GQBSsXQhJmZ5DT6b603MRixmc/Th+NjhVG
jf2nNdAC98OK73nAkHsrCP02cC02bIoBOnBSt83Bx5uY8M/uRd84/trw0AWHxhD7
+bOvi7RyFtH706cIWe2w6NKka0JewZGzHjkrT6tEO5Vu/DTwhMHzQk4ZCywoY2Xc
Fwf7YVfjgZjuQ4lS9xQyAjRcMQ7/G7tqJ1hIS8bsFlJD8t/Ky4igdl8ZgX7rsDWh
Hwe6EKQMl40e6hKsI6hKWu7ZpA0eNnlYJM3l4DLwh6A8ZXAyDhdE7GqWgUSTbjTt
+rR9JPc0D/9k0Nho9vDsOnYQUOOuozhLLmWp5Qzb9n9fDWGb3Lc9H3T2NWw4iOk+
pmuwYh99t8QJCn3M1IIOD7Qrteoc4sG22Jt3DrYUqVRob8bp3zrr4R5x6H3vPjYd
8KZjrmnH3slbVljpvV/aWw0rLpeYM5XmMXSn1nAMCzH6PH1zuzD2lj28ljJ8YyIL
Mn6rQE0+qbVT/sUGre76Te+qgi+pcMQmNvzHqryM1iIxQJbUSEV0ajsC7Lrem06V
qthgoXldPs8+w5jAoJ3WTe/zZqwsiigABTrRkccXGnF8woC9OOeU5h/SKIdl2Q3E
8G2kqLPY4G12eKpdQcTGFos02T1zYfgl6fJzpJ+YwXXs6daeLmM2fysORmXDwM2V
LsWkE5ERD25SALdcRNOdEOZNUzL4dIxSZkVv4mRIMocfSk6vkq2EgG9u/TMdb9UP
PlQFTN6MdUlbhZugF7EfJnhzTcmpz8+xDglwns6PQ7LYI90jrRbbdGy7yhsmRxnW
11kQYtBqUW49B3TBVbAxdlslNeYYd8KUWyuJtQ/NT3Cl4r3lXb3cLPgMFKZMBZJX
ApIwgacJD1s2qqOurZ7+G2p2wuGxm9wX5DngZI3Tvp4TksS0kUP5Rj98zMqVr3TI
2rQExCL6bRnDSLnDmxhQsC6mxffJTAt2nF+JMMiPpF/NB883I2sBd1X9Jn5CTKzr
fjLC/wtiGkgei8mV7IMrbfO3tZH0rj0DrI/nCqZqAy9PunJNfTD2+MgHunrghmFS
KXuahF2GHwWHy+CMr76T1vssMt786tUu8SQnERTWs2g7mDvpAwKwnko12xDxFq/x
ba4lRhFvEFoBVNliwbX4ReWmv24Hy0pdat16/wtzHeN01qOushenj947d9fZbf2l
S1nbxI55b6COAOAaJGfmoYJDXP8DgwvcyXDsq6RVQv9R9IK0uTzSSxOHN7d32JXK
TzFTieLa7fZZQg1m6EvpTnlCjbWRMV8G2uBygvapbGKbdmrIyjSHfgYO6+BXCfUe
0JXxhjgCxIpIpvGK7ZCSC31dX8C9He7W8syr9pvZnK06zeviVxRTuTl+ugUkg/UP
0xxi2nKX8t2OEZdKAKB31JOnmSnKzzn2fiNLFlJZQy5X9lShHU+OZzU37v8tmrHH
v9XVxTGFmpJpbKbglJ74kdqHhYAHgabeSE/JVy5OcFWDEPXks7ziMX0muxkVWim9
1ZflQ+KIZh3HzFvqC2u/gtmA/kM4e6SpVPgennBJb6c8h6Rjqb3r5NWuqP7nfuuq
C3JtKWGkXqaQBorXMHaJDynS2diCzELMDfLdfHTq1XBaT3ea1qQATHceuG2Ugj4c
zvpNqqkB6b8uDfLuTS9dYkFmNh3+y0DSgFnEymo8udJo9ZZ5Qqx9HqZmQH/Mkvdg
Rmt6ZPwmvLo1Gj3GWwhnAf7K5XohgHEzxYnM4dPwIIjkckXydUguv1DRgVpDSlEX
vs2+UR7gGL/J/5Glt/v2i/4tJrOhDypuHPa/7LExEaK4es8Er4iVY3jsHL4ejV/C
O06VBsoiKP0aIWU55Zy1wik8M28BSMeyVd+SM87pvyDsT1Jb5Rg8RovTtr7bo3vp
b1Fn25qeK+/es7idqXA7NNxK2SP+NM1X4+vknVOl0WU5ot2xersRjebOY4+ntRiw
nLLNV7EdlZnGTWFmoMYSos/tOthJeojhUQcCYHBRHQ+diqUlrqlpseYZ6cHthJbs
+9XU6BUJV+fMWVT19H9sEwsuhZuvwqlmPZCwqwJ5a7kAHDeXQSSFuulRAgY3XGn6
81KR9rVuDZyqX3rh9DPro5osXFxVTUiiIlsMHd9+ipmZ7L2gkAoOzNuIxcKhvlZw
nP7LO3RY3/l+bI3vfJE6zntIf6l0PqmRkMbrHFfyPtV8zw4UNQS71LxRXgfopASu
D4wCYScvq0EKpWxMrcceR2Ntaf2pf/843hHluGUYjWprcP4tvShL8AQTi09WCG6s
2ia1IEBzgXT1AC8yTkaSPMRpvH5NsJP+kWPE6/CMdD9i9VzC1EgL7e+guXTgBFCA
FUvCkK27ps6Q2m7CwVX5XrCAlzs1AOJsQ2+EPBV4cHUV8avY52QxFkHtXQ3ElHNf
+FB+W63ArwSxKFoF9gDbpayAK4UYjd0pmjrgVjD6wNXQZtoe65AXgk34WxPaRwuz
GgL2/lp3iQCAAxr56zLqvXXIQiBr1hsesB9QNT/b7hBRQCvjthJZZMPbl/CTAX62
L//Ig0QK0aGeTi+CY9BewEch3ZyCVrPA0mzWkBIhwzaVgzqcmtgg+fUf93zLQ2Vr
3CPKFOWMB2fXlTLO3bMcaZAQEBwJNA2PU3Py+lqykmcWRi21u38Oo44ht07iSbiX
4fnkvsyBMcvq1eptE7wJmzRUCNU/g05zirWXpGbqQ1TKi5zeEodeXtk6OkZF0CH4
Fj+jw+yoKP+kwRx3reZLwF/pn5AEfZJdaflYU30CRXI4qhFmszcvGCf/e8IKdDZ8
HAU1WCFzY6gq+Kfb5O+iOxVZXDhMYrX2xczaOALHPoN/2IUT2Yco7HyNwvKA2kAq
u134002fgCcO5OWS4EHIlGY2QctnUgFxW1FPLwIoRucfIOS6UWjTZEObzP0hmNDI
bV1WcFZzNy2IAa/9JDBbd4B8K3pH2RygPaFy19eBR22xYJ4/ft1LLisZJriTPV8X
sr978wk+Gqq9rlOr6/57qxz/UNi59i7kIIi30aplpVYetdPRkJ04M1qO9n1B6G3I
sUQd/Fc+Y9erekrXuvgiifPlS8sMgcax/gVlvLNDlFyE/Zk/WNr28MpRhTQm8Ytj
bGccwI1pTYp1S5LQqvJH4pf3vd97ZZ8rNjxUnBJI65kbLzuIqa0cdAvhzHJmvYOr
IWhwMcAmTjbeuAN4/SFpo+PnLfCmNmfD41IuGfjSCPywGtcJKYkZE7rCXbmV3R0j
EzZgiCPYm4vaUXK5EcXQgU8ZDZz5uNiCtiInhphrvw+0pqXKERT3H1oqgf6cjeM5
Zfu/j0VrqX9id4UkCVIJ//lX07/pPKOoJwlGQbFnMFe1GNzPJsrRYdvfAsWG94cv
sZROIkEDIRzrgk2qlzzgfnbAFSS0fwRFpjIgM15zqUhvC12eum7LCqPXVJZOq1du
5nfoNYqnFyPSmLejDQEtCy9JMQviCVvrubapKBHR45BoIW4n1lMPFlp2DGB29BSt
X4RZtq3Y4rEFj3f8VteCXLeaPKpdEwCHAJmEG3gdAKwFo5L2uJqSB64X9ONfcOEg
MUiFQz4F947uRsBQfUH/0IkTMIGd1ki3lF5utA7CWrD4e1JDIL5BC9RJ17MExXqs
IEF0bsSh5poyPqj5jfLBhEbuxLiudwtYKUt1cfF5Qnck3WeX5du3u5CQyQH4fy37
ukxkBBVpce6P5jcOHu9RhtM1LS9nD1JIgLitcXxTpT3rhJgy5191ZMio4B0Veu6c
NS4mLb/rdsK/Zl5pofx0T5/BVA4/d8ov7iIFRrieYAI6f4SttC+F0y8Pkm2NsotG
bjGdgvQLdltiWQBa4Ee1YcBsYkzz/LClO3tFDD4IEUXg+AraA9tDRraDi9dDEclB
/H11FiNNoGxQxKwiaOZF1J6/XkAfS2zN6gQPRv1ZgyT1dEjkwbeD5up1zYSaVmdG
ytp3ZouqWnpqGNV2psVjVph9AbP6AqiPDZzs+XasUj79A0r4Cw6KAGwGHVf27Vkc
ZDTXUontqcPNtOv50dh3atWJ4DGcBrTh85zC3cImJvUY4tNlNUHbu8bN6p8l9keV
DyKQ/KqoHoEZPaKai18MB6zXDW08yYR1bm4QDHl83I87md21tp8Y91dHz530+ZWY
GfkhcpQT4qCyRQHEQzylSMxUFqlJ5XlJec6jhYGDAIixaSx/Z2lshIW5HY9jyLVO
Y8xOSToG6KEwDXfIfrKO46dfKkqlGZp35yl/XawsAV5CrCXA6VuCrOTHOBpKet6N
RpI81WglwyMPwOmri1CcUMZI41Kl6Rg9HEv3j08SIH2DQ4ADkMtAewgPc2srD4fF
fVcFl+XF1jxvyUAQEVr9/0jGPcfz2inUaYR8a+GLdcjRp1PPtrhfmOfl8/XcIy/r
WL7EqhkwhJdB93Jb2vnzUL/0H3gibLd/9a1Cc0Q3tXbBE7O6/g0lIBcDvC4TyZaN
kSNsybNUKCD6yH191qHW3VwU9BBhaAc/ki8i8ODUcLYZpqZPCWHd6XzH3+FTZIxl
EgMSOaJbvOpGhCZoHtqg2zX99LFpKQ0jeej9c58f1c6OFQWi2ss/X1fdui1vrMV/
n6G3XSg82txsi1Qj+Hha3aSQI2266obWFmmGHj3cq7NjgEhmGsgifuZ8pFOJxgV1
wvbc6gb09El5c/d/gqW5aLQCYLt130jE6Z+OloxFfFfBZCvXygHCxVOQLaeTVtYd
ZgLLuYOQLNVUywbfbu6ebMjajQwEU3e5qfOLUUnnqVkePZnEJxfY1Rw2Qlnv1DzI
vmrYi7juRjqvwmrqmweXj4TiapvQ1Pz8Syl9uCNm/kRwrqp+NIebH3P8XhZIAno3
SEqM/9Quhv/i4KyB9M6hwmhCS52jrfgDsrGEbxGiVSRmm1ko8x5NSPXtBxQZz6h8
EDhbxUpjUqxqi+37QfwntXsVCqncbyBUizZ2unDbqgZTrIfjoJfKPlWI+kB7PpR6
ly10tlggubuztD/wbpUU171i6b9pdBu0JlLo+K4LrTA7/sbnylPf4CogkFRhZP1I
6W/ISeadl4nmd3VMWuCE56aKop/iekol9ua3FTEG1/AS/QxYGWlQypbU2anld5an
4BC157BYOi6xEFdNFtxQADUkcfgz4BF5cBgNwoww+EITCLqAJ68qOhae/Y2BrDwB
QO69e6mz9H0JA5XZ6IQi7pjJbaB1X7CKqs1gMNshwphELA/LSVTUAxnR/vWR7Yi3
a4Vl7Xz3irrY1pHX7rO2m6gTGjVl1oI+k5DlCfBzhxoyp9KZkIziZfHTTp7KIm0P
eH1sR285AMylsmkqSyPzk7IVj4LWjtM6V+J8pQOeVSz9dQTuixK00r7pyXnG25N0
rhZOhegziaJg7oYx6rwfrDKs07IZsV6rLJ8btHn+bTgGsH2mqi8XkkF009piUTEP
WN1P1CHrb2sz8dwjsRrbn2K5HKwK+dY2xYA482wG9uaa48GwcZEPOZ65qzgdGSiR
`protect END_PROTECTED
