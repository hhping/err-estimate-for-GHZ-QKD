`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IXIuVW68Hf3k4ZFOoGv2ZXtLvlcmAufumMUapYLEEqAAibXddPe/7KoGcWOaOw0G
qm+fpbrfIR8j4Z5ilCQxfEaL8YAtef2OtGoDFFaBripn9K3P5idV2O1/BXJe4j1E
PNVVUCCYty6j0JaF7rgsu0f/uakRfoBsujeM+jQmzrqbOZB9H5ZkXSXhMe8Ygfoc
n+9jS+/vtI0vJsefPHPmXB+q0SjzgwVNmdlA06MKMmEn+0+KtR74Is377c5QCxyO
o6YJnn6zYvtUBkqw8YT2ODUihFfNvs2VoGIdUMMcMwrTQs7KpN30hfPZSQnDdqZk
XlKOMmziKSLvL7L6mwCWP9LpwlEz9KuaX8bBiJGWR8M1nfFhsgw0B8xXC+bMVHxc
CoC7cvoV3seAQlaT+uICsdqUGfHlXbdg4e7yzRhSkS0oQi72LiqNoH9GoawuKAee
nmmV1q8bdoTg/YIhtsB3OzRq0zcykJ4EslgbzDiPciktZINb81M8S3zcNJ/8N8Lr
oYWVkG1evqMKJTJ1RWmvTFMYs73oMPdYiBQCyYQxE/QRsTqEsjI3XKLV9wV1KOY1
cgrjxe37Wtdctwb+ngYlQryu3tMRgdH3WgML6ZzgBlXOz7b+nDckq+Gifmpb1rWh
mOpfJ/ZTbJKrZoQtq+l8h9Wby8rah97UmN3Q/yhzuHjzB40Q4b9yB7cTwfnOcgtS
M6pt9iv4T9jF1ofIO2XbHYu9t3n5d3xSx1BdGpFD1y8Y4KypL5LlGw83ZPKZdQWm
H41DZ2mPSZsAWdyCPAQs6pap3wY83G4lFoYtHbVvB3BuGS0TXMYca8SOwHoAtc+v
kWcQgdwwTaYgC7lwFY+RYu+wxNdUAqYWygfUaOdeA3ZLr8lXZvt5zR4k62Qd2dHV
6VzN/8liJNHs7BzskzCRkKXRs418G10yL/FpUE6Hp874aliPtKHD+o/OB184Ge/U
E/nIXy4JoY67EHDC5nHGNOvToF0Ccg4cKgJ4LyU+vsj+Sw/8xIbHwwFGrvnn2Nhv
toJpNfqkZkx4GJJoBW23aI9FsxF7eqfmVBKp/DOKVAlVwycPLigB+QBNQfYyHN/h
yvScgwJJoykEGGgY2/lxZDItBZNzh0ruFsmDzHYafFNKLrQ2skW80UdD3rrQ5PjV
jql31Q2iP7D6YCOCtWeL5JbCw8gCNUSGoBhqgxjU2QzuxuKofAdPggLg7FwHp5Sb
plLYGMnMN6frDW6BQpPCSJYqQz3Gl/3fQXuCMu4uYmZZ2jfEU8hpgSx4swyFiz6E
SsU25orV1s7t/4uF89vHNihj0EhKKCjuj4zUwiahswRlEI6hQjj5bM0RnOy36n9y
eIucjRG+Bm1ngWveeJiugrHnS/WkfNUL7L4+btuDAbldCb5T7he4Wk9iH6Pe7jpb
yl+I40aCl0/ObsuwYZVPRS0KKF6oMB+6id6ONiswuzgCilajG+zmjXfBj8sEDOuC
vIHejB1htIVlbg0eblIeGQeGR98etqV7Cn4mQrMPe4pI22/o0RnFyPqveE0PRB95
TFLe4YlnBWXuslcfPFDOJWQqWf0atkWfLMj6sthrn/2+6TzEn5xzEtfcS6ekiWNY
Q8rZyioJoZPmarbKcoi4Sv1b1ETkkdOtxmFHNNXxuIR/Qe5lhV8GZdVKUHT5Nheu
RhiEdeyTgLpIbhLNq1VBdTdx1eq9bZsmr052u7DoSVjRHi6AyJOuxj1Tz/KNhi2x
z5yin+lkCcHVkOiDkmHdY4ZHSkmdikCELVBKLwX7XS/NHwxW/dPuKA1bzLbbjCWu
0ZklxkRwlinp0Pg1zP7EzY/oIwK+XS4FMh4pbWsfTuEy1inH9EX1dIXWQ0b7fsid
kdB5smDev7eg13JwhZWjGwEUg5OJBZDhITpUIuPT9y59IYLSOmOGrccymOop7mpB
RJPNskqc7D0s+E6N4s+BIukgXR/mmNI35gM3OsKs4aNOd5GgfyWMF2cOicLbOnHa
DwcU1+9KJLnmMDR5YA2FjtxLl79rBMpiBrj4fShh2ubK1jrioDiH0wUd/H4vyZ4v
ndb6oNb0cfvsiKfCbLnwhSXKj8j6OIUiBwPeZIuQMy1yIpjMbD6ace1mU1I+dOYL
`protect END_PROTECTED
