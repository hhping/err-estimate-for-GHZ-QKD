`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGaC00a2F2pxxvItr9OjtcnmgIFUMf8nEAd+P0Qg+3buIc9ZemPVy18L6qGSTU8Q
dMr3SmC7YK1GjTjWtz4U+kugLH+j7Hi6E1S0WPcURtK+5fvjHxItagTWzcrnAio8
8LbJoDy+oUtwT5Q8FqR3JqYaxkiDyLkkOcZLT7zolmfAuFqOSNcngek6Nu364UGH
nBsiljcSyHFneTPmvZeoHhYmX9nXc1R1mfHFc2jTj+LZ6VFKWxXSLu5xODAAzYn7
6rslQPOn8v6UIiC38zTvI0SNmjvCXRVWiSfZNn7i/YMxalQrsf6ZkbIxXYfTrtHW
29y1e8QoMGeIptk/cWpeqqqET+V3M4XQsi6RzU9TwLVwAtPoofMES9Rjz47xABg7
KtqPLjVuvJmLQR6PmmER7Y05m8h25Y2YWyw93/Y1r94V60sDC+zbM92N09vkP1Kp
dJXwX9N5+yPQp07TRvMCVqmFVqmA/cZkdF3hPJt9Tr1ce3yMRa4ZwrN84w+xdduv
jvMk1xSfry/DdLyF+1OB60n3qKF1yKMfiUoUMDkXAzouQi+79cCKrw7weHAlllWt
5RXOBC4V4oS3Shvp6r3Xk5EL6Sf/MkbB9VVSbQgRboqsLLOgWrl/w8PyUtFtBjlM
FYEDVVbWT/g7eVtjZndmkz2I4rqQudZV8qA7toxvkh45Keu6b/H0yO6y0AQZOhj2
Z3zDTgStcPQG/rltw5CyIMRuJ89bmzFDDRtgjfTdQfqtqoSFidZBhpc0zQEEX/Q0
GC7qz+wuSwHovKjU2xCsS91h+QeHlNAJYDzrHuc+hj74oBgE7J0TiOeQPKxZpsNb
uZHWffmPuN9mHOkKlnYx3nDwd3EBSJdWwd/ypoJmjQzHcfk8fIpg7xgOos6Kxd4/
nB93iw4M1L0uHBC2/WBic/jNo8XdORJ0Z+24k11+IwZCLBiRGTBz3aIFUXen0nvL
eVxF5gWGyFOwWsE5w8xMGnmpzpy5m0a/QW3FG3MeP+cllE4N6scbjYzjYXC5C9Xp
N7dp330soo4M5QniwYLJMic9KjUHet9/F7C61m+lQRyJNClAkBAx+I9xJFolR85H
OKBVjkXWsYBXS0ZTZYz56YB62QpL6VcMXPt1FIHzHAiuTZnZHhHQAXAtuoRP8uvn
IUi1ayQlZHwgv6ZGMkYcB7LL9kyVGE4woG2HTs14WPOzaTzaT2iPSqFYwTL9uGmE
TYVZ6U9ANopIMfz3uq301vWK4yDkuxPj5OuiAdvOVc4SqhefgJn+2DSDucESR600
eXiWRkY0wi3h1TkjEQzfRKU8eGQEzRb31v4Aq0mwI/Pj/ToxRgjiL004p5q0nhdX
k7uo3prqfW2eJluwbKUt84rDKzRPBc3BLsPfLjx01L7xB9lRqhy8Mt5uyMJXw+ST
dCGfg9Vk5ekcorqtckOPIX6bEt19Nvb6yQqOX+XbvDuGS3sePeiqq1mP6ZSsv8HD
s+Vgl+SnrSixIGsNh+tk3hCOm/M/MyFpOlgBHMXD//USxtB3PIxKXgi2qGyqh68D
P60c3PXmIRGeEPCw+irKMisqlg9OLSvx0tMnwI+lE4ud1RxFdKMu8kWf3mUzWhCN
K9F4neH2qZudQ0ev/HZvoJ3xRQkihh7Zx5c9OfaJdP6MXKH6TYJ9UPZGhohLtiWS
5r1cjGYYnxyzv+MG/FUQXn0O5sbtP991XLVeDZsMX2FKMWsQhe02hUfYbzXoX49p
RdIxlnAf9OO8WBD/Vgg6QVBu6/n10h/jwTI8RJ2TGdrJMX0bKM5vy2NR/PTVdgbo
KZT3IYIn99yeDX9jQSF+evZ0abxeCzHCwq5C1PyUrfrTMd/XnRXxMg+yztIVzAxG
vE7rPjnvMOH0rvAppU4VK4rbalaOQHVvqdb/ov+YEqTSs32jNW5QUbFKdQPTcmeT
iEQV8pFHeUOMtPXAXvBoIpBzN7a5k09tu//wys9JAQzd4GGQbPECyJH9mAhpwLTp
DEyj9SJJ95QFSNy3INuFW/K9CjMnKi3o2pjIp4OxDj5FAt4QwYIxBzWppBVB+thQ
5hMEyU3UhaCsCXaEUj8gZxNK6Uiyh/rwL05uYMTERbjfH/etZNvzwVHN05xz0on9
MxJReKPoavL9CYEflzPri9SygbTvbGr7FFBcP5Eaa9/XdKAYef7dUr5CKHChbFjB
BzbxhesNlsc0jA9X2I+DQ4eQPXyA4PPPLoja1uTJ2ATMyfMNQ/V850n8D+DHMLv8
PGo2eqIGgHUKQaZcp02Elk7VbOzTPCxysA9AeKfrIZ5PlmLKrRShvFbz9kTVyIJq
cjbxxOKvIu1etmHH4CZ3ZKDiCbsZ6VWfjAddb/0QYnh9pK7RgX9w+NUpYFrATtVd
aLcEZP9qTSiBNQYLUx0qnHp45EE/qrUnLwcY4Fa01XBWcUV0ajVByvyiMWayTHQ4
f4KINl1DkjUwipK2IjO1/PBAiTwZLghPafztDQ3HE+e9y6FB+hahWi3kfyFVW3qY
Mzywu9bYVxWO5lcSw+pRWJNaLPjpAH/W714xOj7Db80aJebJFTY30OmWjTFYZrJm
rpuwjlb0KfhhjRGUuchYY5pTGH8SxxvU8MSVnzZhcgfFHgaORnGEgJ4D6Pr+5+iW
DG4T4+wQnoEu5zF5x7HbpX8hLTSjRmH/5HA1+s7QBMx9LuOLgqvOf43ERvCWCATQ
6oSfxmkGT3J7bglHpbuBTTkSQL+TYz3qhebTo/pt5vTt8U2mJIBlmt8HoMiYZp7T
vkFp1klr6hBm6WRvcPisux7nalktPL5LSYltffXl5AGuS148QNPZIvGPnEAK8lYW
QszJF30kGzAj98ANvVlry/UIlWDT7+i7m7YzuPOUP92N3OfTLhMlmTXZa3GQlwYZ
rSufS3bf7aSLjt3ADpeOEkV4bF+5qw0raNUPE/WrBTrhtnrhbq2reDsVIwzO39pw
U9DTa8gj7Qc2m/0yteVSP3AusDoTq8uTOxZLDn/y1SMfy097nlYpDPIEzuceAoS0
NZEPt+3TCL3qalmmdLHKAU+/shlqeqMfixevPgY0bSkdCBpUtfcHS1VDzr0yq3yk
3DWaW6pmxnlOjBrPj8DS1nH6mGDSGD+BZiUhZJdX1HIowk2028IhcQEe/d7zdWc8
tIoza3Pjbv7OoXwcFBFKHOXJU5j+To9FsXRfrAFUGw8XbxCb45Xfhp//1t430K9J
7sbMrD9kH+VFE5mbP4m1aV+ncK2/ur4FSUaXNPOT6LC2mPfSw3EFBjH8P1lSmbjw
V3Wh3JdIwQL2+Ts0+ZliuJQdYO+6w7DpuY26PxaWAGBruwGi9OQbbzX437t711t5
pM2BVqdjJCvzIhIfmkPcWp5FeFyfX5Ayv2Q0t5Sp8rOJVxBrZb4OmC1glCxQw95p
j7BtbXW2c0NslCfzBszFyhbMo1nzQFYSk2o7BbCprfhe+DZ3QLosKHZVGz74Obek
K0IYW6ZS6nToIoclzBRCULQZvY8PmCmMfZrWvxXYDA3nKo+J5NX+RvSNVxE0a7nM
SIwh0wSxfjO9F93EygfcuAcYPlSj9fyiPp/cpu6bHgjICXNBYAgy4wXvnUq15dJe
lpLlwIahc+7kMBCnuA4z9iIU+qqk9de4xzlRiggPOVlXfoOhMCaZosp6LDLjJ261
quSvvza0Ztfnr/NIu+0upiFvINfACU9qIREEzTQvEJFUldxIMmjos96ZSiExsT/D
uK+aosNzAllBmLXfd9hUZdg0Cz1k4juROZYLMigP/fk/TZVvEj+FGh92BNdVKGif
fz/8/vedgKLWOeDKNcLGvfw1X82MeDagkF8gOkKuRjiN3DZJNriFWbnFGX43VHlw
9n25NY8rmJnfahzGE749dTpChNn7xiHzGxJIV/qSVRrw/jnK6VL1Xe/LxKvAoJVS
6xDgrHMTt2vI0NOcZKXyPxfXzNuwKG6ulvtO3bTEFcSBoH9141IasBhtP5pRiElK
smg8v4saVkPAObxASPZLpgOOkSQqHrVMkS79QdRndVGBTIKwmgz8WNUsQhCrRHrE
rKon6Dz1oI7CzIq86FBXytF06mAzz2lsRqu860ugH4w7QZgb1Nzt2FKQL9nwQKiq
JAn1LnaHmB/pTOQ2NSqawYafPZsn2hqSAZcLAXL5tG2uJq990XOAGqHPRArfMq0o
CHY4h9ed1o1yu4e9igQ9FT2Uo5CfzvR5sN2C/pGArBlS+fvMxeKr8OeUE/kmiBPd
Ye5ErqDejkkr0DZfWNap5NRSeZzchqxiNZ9d2y+yVdo547l5aOHH+eHH2Z4c4wz0
eM4WLcqqVK1GvQ9TGZA3Rk+9qMbWoBPhzl3fXGDOWuxsKXMfNDgBX1sezKkeLYrc
beVbw2lg+dewB3sVm6W916sdquSTbYke1G9xONeqE0cPLSrt3IUEh2wz0Hz8lvtU
OVDL8ll5jbtMP1o8/l3u/vd0oihtwxA0xZ2kIA+Hr0pczyowvN+V0Y3RY/JVpIe4
ZPgU6wp9S96pq9+7Xo+qSu2y/jMZSqr/oTWFAcThRPmUnff1ZmzVCD7uqojtxTab
7d9b4gp1QeL1XbQYID75Ye1XgZS6CmDEBTHU91Ydfg9l0aDovdfr7O0tGnh/Mwp2
USQFlNjuLr+tqnqgkDXQu1qcBGioy+PCb1pDkDkIZLDwVPLTwbcxco2jbjrxMq3c
ZAap5XmT9KSr0R9r26RZP2IDlhMfvdt0PU8ziRaPO6oqeTAjlPg9d0eUjpV5b/Yy
zdDrzaNEtzPA8wSvpxVcObg9i0Gz/utwfUtynb155iUmWqO0oeq2TFm22qG4Wobc
fiw+0tUhz5Sn02dtcMw+vWmSRpfPuAMCip9B3YpqwJBi0Q0m7cIHp/cjpSh0Qa4Q
qhY2MHfWVHZp1jXpaTzTVUEeYB0HwzmSCOf7N5iu0Ri9VmWWZKo3ETzAieWbvApU
jhk01r9exkOvYKrjhF0djD4AfDT6SUJCJ4Ik/Wyk6ZItwPfbiStyiLiaeXeCjZgU
vvhNe8h5md1MZQIQ3lXupGKet1ASRiGSveWT6RD/mfEn5BfuKnMF9Z90+eU2PWzm
s8A/UuOam15+HOmeHd/cT852bIuWyVaT3CS2UgFeOiiNHB+LOYcqTCs5XZBzMIaB
jUfI60/M/cpmYgdIMH6j46/uA9vZcoeX2jDpwnKXnpkmGVXe4CizIWzj/ntyiXcy
CG9y3ZLA7Xkt/aoS6EydWjIA7HA4++pthoyynYQ3Dl4C7QskYNy+RBc8I/HcRMZm
FA6To5sAgFcAjcJfZBugwh3FXMYko42W8fqA0ILthx/iBPu+Kdkb6GrGdoM7Q7uh
SbDdXMUm1H+Y3j/QFHEluQAQVL1oYz0YXlEe19CbWaCdoC3gJN9d+6prX2aWeYph
GSGHDlw2fMYO8BHog5IQy6R+cRFTxhum5wLn+/M3/HecIPXCP4/FRZ71vV9lWGc/
XAc3ilFFmtuZll24dZFKPhnVbRWDwVsSFujEafVF8dbwn1m36AMsQot3muTkiEZs
t/0vh0euDeyvD+clrjVqI6Y/91QuUHREm9aFIeVPI4y4pXgcLcQLO9a+zow+Nr1c
59xLVujgBs9ZQcg55EN1vE8mJrc3gZQ+YDV+ZLWB/LqXkcZol1tmSnDjHU6Udj/F
z/kcUC6qtlLvDFeH0N1VxIXUe3xf1Y5fXZpKrAXOBwj8FjDKKtugUFEKGWGBL92Q
pfTl4wVCSXqDXz1FV+3cQIiMFs1BApREH8Q/VtQzjpPvqZ8OAdQUKVuKf+cG3qMC
4E3hSFkRSBlorRGCAZMwg1d6mY1vF8fbJ3FGL+G1DllqaejP+dAFdWpLxEzVlpxN
ONGG434VOsOpH2R88s6Ttc582Pu/qFzByV52i0NvhzbX/GhzmLf4fBWbc1FMIlWU
Wk6TyCkHuG/0bPFElAJrqPisppJg5tYG/3v/vJkTP3T0Az+FxYJ7JNsVIU/kHPdn
rS48nsrPpRHMTyT2RktSIQHBjE/qabfMQpYOSgL332uLj4+/G/+NX53ajEgOtYMX
+5VGa0Mp3K86srHQo2kq3V1A7T1pxdzP9S1diY+lsy0IkA90IgnFWE8+4LCHScvA
xiDnR1brsgB5xws/GFfFm/LBdPPDyqwpWvooI8s8HyFXvXBV+zl61llRnGGoYQho
H7Pk9f8OIHgL1VrtJq4w16fCcOuEz5UbOLpdJKOdwtb6xH0zv9zaqB2zRaDdQ6Nt
TOxrFR83uTMlZnhCayRHAmqxeHksMEknG6h5cH6IPtgg0hdJlK1gOrPzl7qj8DDM
fEqKcn4AFmEiS4ureDg/ndhwoFzxJtRPcVlvY4WkEiiKyC3h9K76/5sMqgyWqUDU
EnZ4qOWxr8rwvI3CUwijHO76y1oidvYF1PcgRf9qiqIJ10kID/21SZyROhhokQQk
ImjJIsYKrNNVdfknbsRh+MB9X2jmd0I6lJ3vY3Pbk94IOTrukHz7geY93yIM910x
xwlOhOZdT/CAWsIFB3aNNsiikBmaLH+4xDQ71iCelANEgTBjhYWHZIAizut6ZeGH
BiNuI/yXFpQJlMBzPlkjpQAmc791KZTpH4cDtdpwww0019RI3uobZkGP+D+oCq1M
uFUxJ/OQuRvJMKVGWIScAnTFDDA09XdOPWN7Arzdgjjjr4hDmPV6cmYKLk8YM+gs
vK0HYKWeG4aYIW3UK5Om1Ut3KXnxP7VD9kcBOdvNkrUY0ly3gQ0TY4wiQQbxuhan
SCAZbesGWN9QU2VlcyyuluDVez1T2PbRhiLy46ig00RXiMPpxr5VhaK6fT2YtNJA
JvhP+Bfd1KhHdk07nlLau9DUBYxvspa0oUDU4a6Bs7hJHKWImLVsXx9MK6H9hsNJ
N3yga5/h82goU13yM43uDk2ZuyZ1aUNmBUIzHOvz/9xnqSpPcw+3aqTJIzkbyw+r
eG98qVMcMgmtOdBD68bblBBfxBS/nOzCM6Ll3JbXwcFXFIJpVpl8JodPQ7KOCcHb
17R7hpSTS3ieXhy6TZD/1AiQ9xrSo4svyHcjCkbJdI3Ze8CSPSIJF1CKoPzK2bnc
BOLEY+FOjc2zC11yAmvl4lC3t/izY3RW8zzQrxOXFmPLFkb+9EQd/aN6vE14E993
s+v+HRWwM6bXYpg99CBtPzWecBDaonF40l/mJrs+I8BW28rLuI+pnBh5hjbT9tYQ
yS1IQOvgokVzZRljlyY0g2vBJ+XtzF0Tdncjf/ub36KRLvQgpzfXUn0/L6N3UQV7
/x83OAs12wm5zDjg6pAkNHJ/9iasNIbBnDWn1b3cNO6VacsS//fduJYb05L0i6a/
Gy2/wh+0wK08D4YxIazYX81LHDr1F71rLNWhuqDDkrshAFbYEB5i2aP9Z/b/q7zD
iCRKmLnNFt3tsoRiHDeZ/uuIove7HHtL18J5fApgO8wXqOsuI+mIgNzCS0Yt0u01
9yr9ILuPXPchatYTXyWdnDYYoIg0SaO0+OzvIk9ZGoHcGXEGsedO/kKR0Dye6dkU
KsPCVVweYWe5JE529Ji7wXpivJW46gJrlL19Urxx5jgan1Fxs5fup6TL2bdcIZpf
0g9aC+J2vu7gxuBZfom0bg7YuxpmA3b1vxAAmDiWv3RbSi660v9rdMXgVR2cHRVc
U8tU3eSjk9LQCYMNYVnC9IiN8VCh5N0RrcZ0/gy8snYUcuMFt4y9LUYrBiOwGwQL
x58EKgOC/tJg9q69kUk08S8rtUbf/R3dVri9y3R4M1F1OLAcJEXlf7XKCUhDpFph
2XbZ35MPJalovmugsRkPs39KJqniEZOyE8EFbDS5YTnBSuxzQfmV6WbXfHxoz9qZ
prGO6SWRBzzmHjWGI24E7jppmhv0r7htjGpYJmPjw+oh4BJtQ2xCc8T1MEhTN00k
JUfCAYQRWs1gERXrGKE7TY9lMzGAAfBXH2ZuA55mZG9HrIHMWDLVwayuIKa1QwGx
D4U98Q/eoEt20tLTLFl4CCNiKsY9pc+E85N5OTzl3V2me2DZ5NPgh+pBikfOnHoJ
JHCI21c+bGJJ49E2QnVUyQOjdfYPj4kmOFlUlJtFAM+IsQ1J7oMJCr8cqknxkVSc
UmwVpCUJayBXFcm0Ilc44FusznyUr51G8DyYZyf6eARZCxZxPDzhUbUHEIMdaiPB
JUXvVJra5+IXE0/AcHn4hdy85PTD8MKK8W90XIDt9mkBOi/ft3tKYO0udjS2+hJy
umh0lV1yuHiYAYjUkM+N9Gg+IkJtlpYGnqoPhY94VJDE/abM/k1IiY6HeOQX+s2y
XVVrp0tnUdx4i4d9GoF6D9y0M336aqMMhnwQUK43DOiR7tC/tzaP4KYqAAKVwHPL
JtTrpw53da9xMsrf1c6/mGLuuNzDq/+A6O6nCCADq8ouAQIC5OETIdcfn2VRhc1j
UFDmTS4KDCzPy91UzY9qmZUgqT8xbSAKJOAOE44hgvuskEKZg+e8Q1hI3XC0XEVG
H6sLMj3QPVktmjnfbrRnW3W4tQoneOgLPfKuQTeTfWJVcMpIvIONIywUkPIAo4rI
VkARvsK/NzRgmTEK/GJZ/70Gf873L4+8JsxZAsdga6LDDptzpjlpbyVtj83XUnJR
0mtsYejFajU6e/l470CQatq6hxRc939BCQ6fdJUpQsxTU5FKU3BLOHj/pVknnWJU
0czhaV+om9lvFl3IScOG0K+4lqTSEj6fIzPBnss4NLtIXPlD61Xv86yP7kv5Mei3
JqHtYEn1HvQlZmiUU3mk1420Qj513TfZsOp81tqKSxWZ9NcvN/3VAMn9TXyQSzf3
sRWojq5L8LiEE638zrslEG9qQpCzLpNwVakx5e112cV+Ycae/7K9t+Bz/ZabwTYB
o6vun0bprm1XS3nh6aeo6OHz39h5TvHyYhwfyEctKH39Au7JHuiiIJ3PqXoHQv73
IiLW0k/p6+Hj9Tj2oWYQSTzWOSMhqhju+D0aT/i+pA53hcit4mnvaQeX06ykkF1r
JRMkFGHBaaeF6qkUsCdqA8/BNHQycu2/jZkcYiz94Pe/H7fjDT0/it9TidjHCTHN
AFu1BL+CFe9675979pD9N+Pw945yGa2vtRLGEylJyY9sMLzgTJnTx2/zE/r3dJ6Y
jo48TssKg5NbyVza17uVR+pBdEW9YdFAGw0pEDDE5GCvGKr1A3uZ1D1sAuXkBbTW
giy3obxKy6CFo52goDFKfnqX76gRZC/wPBTavtI432NFrbSrZLz3yLfWk86A7wVG
209U5MYpQyiA+BllPQL7RUxrPOctz/EiJX4qy01XVDp/C3yAaCCcs/MmOq2JXOGy
8uZvTi0Kx8h7SknXEjEaPYl4Gn2h8VC4d5FO+zrRUMNE4uD5TwvDVi44F5xhnrpr
k8Y5T6o5Vyb1p0D17/XPaLdkqGQe5fjqX5jXZPWkhLTO9Sq5ZmVYyy4kvhdE7eUd
Ryntx8w02AIilHX7WY7+W0QsjXPvkjC1uUQJWHDVIpFRtOT1ZrqEUMLo4qy8E5MA
6m/gKBRde+dzg37pWt4uvH5iNPaXAwv6k7pShR1uB3+GTw+qCQ7BqZbogRNY0vWx
nn8rXzrm5PZEPyqUQ6tSFNvNLOLypQ4ZMI2T2ReZZdcmcpHossyWyi6D5K2a0q5B
aOvaFdPkUnXyHJkuzBL+ssrj52KIBaGuMSQDUFeBF0nwrcXyOEMUzjVeAoUtq6Jx
+UwP/WTFdEtaPS4lsBu9VvcnKCdLpRPoSWxLtCtlkMHnDWGJJHNkddG/QWcIx7DD
CGqLCwLNM5UpAS0Y3AvShlp/ZiSC3sCL5tQZzGmHKRceFP1RMFvTNPospr8Eo2yj
V8JqYhX2yT7ZkNKV+b7dQJjBJFUlYZGhnedphmTxGWsP9EaO79+ogelpac0Lme4X
P86c4tSeR4F9JDYLAJOi16E0ssegDW8qGP3WtvIcWSNGllXqdzIeitbTPPGMdWTl
HGcGZrNXjsii7PhN/QYSrXOWDkyey0InrpWnC/ovApNNlco/zN39lFrKftK7FSKM
BO7mduY+kQzJN+9teBkfHm2hYS0wABPk9JCiD3OzEkJTBf/YIqsFBWy4T0SfoCsf
AmexI29ECAKZRlfrYhm1PjYUcVEwkG+HrWPyUHzTv7sfC91JCmvrx5TRhChZZzXA
5Sok2hs20dj03pqleUstiix6j9bYL5mYRxDLjkJbOwdzzz/IJT1x2Yd7fp9oKpOn
FV/3cDO1uBysHb9wIiJPk77UnZ587GUra6hvdu7ekaXPLelsPemuBwG0/qsRgG8d
SXbNLyyIY4rHMrn+znmq7rg06vjfg1j4KRWCBfjAnFkgivVP18mzUZR/pQnTPzSJ
fS5m9Tv00tMN8aUyIZhMR0dMULo7+Q14NT7OzdsYYIkzegMaxUSU++8pmBhxAkDx
DIJj4RiWtZadB0hKnLOevKEhEaT2z1BLMbY1aGb5YL1oElJKz5kAzxD2PNgdbey4
Pzy6iEyXqNTF6LZVjL6qUDAgIEZ5/is1PHR3er1za91Hcnh1LQJf8MZClvcdH3kr
okbKbrzg1vrBm5jQBm9FPQVLZh3CvzjSDqfJDwX9H3UZbGODhbeOZeB+FrrTBHTj
jgsSDGvQeNM3CNrdGM0WIuSQ+Ur/IrBDmzoItUYzcpT47TV1juDBIvYmqgoQfQ3Q
HkA+r8tIX6FkZaia8cDpcEokC/+PlFK0DcA5szvm9N2Bw7qN9FIwAwfyOAdn9eg4
yN6UHWPdlTHSVNF7wVMv7HD+PNV4cGZzshVoZtYySLkEMRBY9zTQ7WvbjAx5rrqT
9XUfb/9+LcDqqGz+K+AjiIJzgA76xqShOEJrpAGkMWQ34FJgeY++m+eE6oDzYpDD
plO7UrzINKhOXLw2ttV/0HM2EoXwaVfBQZ0ULOCGdMPmT9MUJ1AgJx6Z7QEInF/g
wjPZQkVuxye+yUXjuPgGNoksvYqieJn/EBcM0nfHGQ5i/5kHFRyuwNffdjZsax5G
Pfh76JOUz+3MdBsP+CSqABNRtiZJr/Bd6QzzioX1ruKVVoSQ/w1poNTYCXxwA33D
kAXI+ip7aGaBbKeBM++2ecORavlCrLQGihND+VarthQvVqatM+mKzV7reM2hRZBx
Hcefkn1WoGNWTJCfIoX1G4bYmzCsStlcj6OQmbVmbBX8CID1hWflaarY+iIN++q8
cTbHiDShv7sOgysLnOiuaNf4ae8cPCMnpRjDfmP9EiYBtIk5AhMydhm5APxYpZh5
77YhSTqP/GjHebW2HcOxyOgRzun35uJylgUHJvKiXhg=
`protect END_PROTECTED
