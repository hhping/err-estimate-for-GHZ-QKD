`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QL6fLoVIelA0lGmSnxm4/H5l3KXEaPLzzCM3VjvUXq/4gJzpWjfLV7Ob3lHXZX2t
K5Rx2zvSfUBuWrTZ/rqSl9Gx8OkWKX4+d+KJ9wavjErcY74S1JgVTfoljebZ3itr
cGtgAP6doW1fsQnsZ2uWNnz4Xy+rcDFTKlmko7LQUJ025HiidgjwGHS3TepaWO5x
CO5FMKgEQtt5+ecUD258j9fuDiodewqIDVq7boBLI+OCFfGTGrJpGvPwche/2eSt
C/3V0jgyyb8VF3hl2C7tEuqATvqEY/WklXHK5uvTXPzf3RtR4gCJPINLaRhD19ye
RgMB5C9K3T+5HrGR5xSnJrcyf/YadrRPBEnkXAskrE932R1ya+P0oZOkPyo9BkzT
b4S8kPWqa64gp8RUx1lwJzH+4gfZ6AsJD/igMXftcrBLx9KAc+Rbj7NnzyPltdtZ
J9X4OANjF9aWh0vsoIur7QMl8bgHuLS4HYWGHJGwuhgfDfvxPaWjBKdSRiwvhP/3
wt4wtex+yh7YEIjG98NdW9lMJ/Bj3466crKXEvW+J3bYt+MnjjemdYd2QE2VZ22R
KE0AZ0KE0TQ9+uo6etde/MKoYRCKStX0Hr3omN3DLuKZPRl+wIkt9A6aW7fhax04
tx+G3iaPgceBV3csqVejfY0h5h0FuO/0a3Or4uiEMAQndbTVznJ+YFRse/zLk9EA
GXLNStIUvdnWyXhteyZuKkyfdZ9YhTHv+G0CGbTg2LeGSvqkTHsmR/gTAR7vdiZb
Xx1KVOloGhHOVkijzccv1LB7FpcyIZ9qyvDVe5OWkbT2bl8P1N7EbFEKLMKVsS1d
PoWBI6hQIvZy4S0TMvVj0Sve5+XMbFDwEZMy5MXmTHp+u/Dh2ljjgBXLC5zJr8Mp
VcAvJjsQqtZYA8dI+vhhwgQtbyfZPOq2pr91eMzhjh4ezryBnoz1vSrCQA2QQe6E
Zi4+fwPb/Zk5Rr0iZ9gdv15wCN+99BLSOmqBfSNXV4ug2m25bPgKzaCNNsqnrhux
KJ2zFxpSugzuv3X6lbUzP8RtXvkH05UhTs617ax+Ni9pvTZLOm5XSJRdUXM1aqTA
S1GBP7KYnjTy6OkpW3gaIOkgLwdX24m5UFc7PhO86cWYgLq4BAo7xdiLODkG0rxh
Ve8REv8PI4T934QMyNRBvz4P5goMJJyiGwLCqXcEPi4fyQc14JKVB4ZgjBN023BL
n22eurJzcXk9oomLeQ3XKF/fuX0ctV93j2rfhdGZjXRp6Bse4DJ/XLzDiT5D0ZPE
wUuBGUO+gwKJ2PySZ1tkjQfekUL5sHA1XUAmfdLr5E6fk95HwaVXjrZvJ5ABwPft
T9cbhOBr9pGHgBrMmZ9JJzHVFwK9CdvyBIUkLt44Te30pk0jzeId8pAxYBm3dTFX
XWsBaFT94c9gX4YmM5HxIX9nZBAcLndtHW532Ez06YtX08XgD3XA0ERUdgnqyiKl
bgD6cfRjy1dEPZEoA9ln/S2qFRNdguzjq5ZIw+w5+nG1pULvq+xPJS9WG9WWTFUO
X3uDh37IfrlGbSl+zqrvmKlW0Y4UDFVok1tPyQomo7qmQoKXDPhq7gh6GxFz951S
q4IVm5iAryIh9QIYObyZxshplSvWm5guiMLsboxYvBe0ZRN/RX6D6ZKoq/q88nJP
GrYOISvYqeuDM/FrmgnxvL2R0dED1mzMt4GYaCP635iaXCq8+TsBwbrBXVpJwEi8
qc9a28k2gVwGpFeWyaVBtAs/XBk735a9fab9LHsx1de3Y1lIS3/F5uXzyQnw7Q5E
zzXbsPPntRsCZSheyOvkoFpOmfNmUaQ2uqiLPuaVmy62gBJkpfufKmtW+MnE1oAp
DaiRtiJWQa0zmL4uTfFdhLcb+hhUcl8Cq/EUpDc+htI2CpmcDMKOIDbjJP2rYonc
nDcIAO1nfhZlXXN8uRqyWi4wV//7fcmqLYnbJLj/H38O3gp55iApsP5QIhJaDGsQ
SAI6YkpDEtkWW0c3RxaAjQ2hYDi6Sg12/dADZCoZb9RF0sHxol/3vSWNO945h6Ow
1KZS4udiNdpAx+EUacg7KuNFttfAk2V8UW4sN+LXsZO+HzkOjfzJePsx0Iq4nVic
dlQE18i0R9GdlINfvVI1ajZwO/ncUuyoUfgqJHAKcFRg8rwy5KktR1pupo6coD84
eVJArPMprMThsHThN+hdDfb9EVJ+vVNBsgrGTjIBWIph3K+G0UPMs2N1OqKdXc9e
LRWqxGyY78isSVJM4QCPsDfFdXYawty2lWXRv1IQDNeGORZu6UgZJP0Nq/ccuCkC
kh9nRoF7RQCuTkGT/emVBWKQrBfvgqSqqVoCaT7Itc44bGL4W28s4ra7XDXIE6ne
2U+ZTWiZcD7VXtxkVfbYDxDaowz5YE6A43t4bIMly9PwA7raUTE+06Lp4pkm1e6J
wQO26qzI+oOUjJH1/3jISbluaiRt3HLow0/3e28lifu3kbTbIvJhAbvMyl4vjkSy
sfVFAyUgzSl8QvpYMIM+XHBILZdzCIwBTUcGfxswr26sZr5n+L9CyjWaQSlyPNPU
ezgcuhZYJkyMN9wH7pdqG4IzqZQeiE4JEM63256p2pSboyrv+LJgZAZes3OQD7pF
Wh4csjtq4KTXencsP9dOHl+jr3xbcgrBfVY+0QSx+aEtWN8FTlKHvfHxeuuOS4dj
0gCdhob9ciRgLOQoG9f7oAHAYO3lN70mLRGyKH4WMV8s5Zi2dApvJBlavf68HbRv
kxIJ+D8T5xtu0JM+HrG+h9Z+GoSnJZj1iSz1g/Fnmv9QTuqoAChgnN0s44ANICEm
jpEwbU/SVu08GCrvezsJiyMg7rAzrlGM+pHCU6EYujr+NYH3pmMCOZDmKFH+zt6P
aiBDd38XFqjdh9Vb9Yh2rVim4tpy+AQjMPECyE+QwLuQG4mHykiz++5nRyCFB8sa
g6VL4ZvVLPnUEFgb5qRuN9LDT6SRJiYkVm+wjbpi0Y6x2cEOz/tlCfmXP1wV+jku
qROkO8pSBYJs6kRGjVpJhdd3KrfZnTGOzI151KOU3tdy8iJFQ7E029ufr7nQc134
50V0gNmHfVVGU1IT/6oBaysWAT2d+Rgx2aCuVeM+XXfrLOojWsW9qaqk6yDVjBIZ
pnI1iPgdqbux1YbWuzvMRxIiY5237ZK9PU5vPoyrQ7Fhtj0OBiwooxqEDeK78wPm
0VC2SEYWAMoEEbWbIcFuh7ZSUz/xKyqIFJoQ261dkZfsNBzRySDRC+k5OZ44Lip0
lkZkmUR5RXuXYsbAybH7MtHUCKPN4zdBixD6CXE7hGac1/StwTSJ1hTpZqtM3Kd/
J/2hj/5Mx1yuZvObIRNwOyOSvpNOdLSw/S5JQ27Lz3AW/NrdYXbxoLDQJ9eqevb7
Rsitu0TCYslBmEkUdr8Nz5oAurCyyM+KWdCY6VLWBkqf+Jit4osv5fpCp3yl7Q3n
zTfVGHtFRre1p4OWUrc0MJTltlbgXabtpWkE8kU+GbuTjP1G++ubW/oHfuxhlmdO
qUTLpnM0LiSY30MWgC1RnpKSoq4zUQBdQ/mHYW56NlP8BTgWFQjOwUGbHJOPCZXI
lCHKgmYYtpYf2o9DKsF377+EV2i6M+dyBIM9GuexINgmXSZQfxCHzmGvWslntAIJ
rtNIAB8U2+NUZPPOA0XBwS8JW8kX0uXGaFg2ILM8zQTZ8IfLb2xZpX9Avza9pcb7
E2B7dpINino40hYPFnATwVPCeYclEomBnZT0Hc0kqLZcOBaRk2jjORU6cWD71hLt
fmG+1/VLyVfzOVcjN94xJIbIKrxNTfs/LcS1sRECZjfxW9eHWyRD9a8hkHNMueC3
GPrOL9PCoB/CQTMRaKGFgVEQ7j/VXngcf0rd7Qa4fE2acxC1MC9su50Eg6mfV/3W
1O7Um05lV2gTWeo0JWbhzvU0y7/TiWgyg0UViZQSy+NEvZBmA66TTVhc1FTs/Mca
+m5dSnbUE3xLR2t6IcJLpJ5M7JJ5a5Pej4FPu5YgfAUle3kDNUJbIpCMm+EBjql6
l2MrXW3XVgRzP55lgt0eQagT8wu9PM0VXCpTa3WKeF3Tc9eHcdzZheNEUPUggd2c
B0Jag5DcaHYUUm7pURApUCSSDCtzJSUObmzJ4QSW1M8dYvns6g0qtS7SuYrxKbeV
7UWUrKJ5KrL8YaVmomBG+wAfPBwPdXsJvhJsdmUJvKTqnREesgibKcsQcnfd01LU
M+mm6D/dv1dLcyEfEt0FaR/HX7OUgXkIuIMmftEgFM+I2mHeslKX7w4/dLJxOuJW
4EgplN5VYEYcc4IPJIKR1CVHtVJjQjkaRszYsnHY96vzbb/9dhCKsIkV9d2mSVPG
BOi9zvhtlaIClZ4cd73lyUBcUh59M2baHsCDv+ry9vKzwh1x/PknJOcBsjEYl1jn
Xr35T7pL2ixu+89poPkCXr6vPTf7J8/oDsU5XpJWomRicA+SDRbXpQ2/8VzyN9VH
BAw5MmvO6WV4muaCKHpVoWF4f9M6czsWAmFmv1JH3QkfInyJXcliM4FeR/o7e0un
F3yRtQshSBXgIsqyUT2W55V+z0mg2hP1ge7IFB2wzFpSYFL/PHmiisSxgJMMMiHk
Bb+XONlgDrwuUT5GeZcc03ECpybG4Wpy8kTG8PZRmnf+DDI2OphgWfsqBqbyWb6d
kSXi3cHYr7t5qKCNrugXzfNflmhO+NZgPgJoM6iuERaXlc4837ereRioGDE2d7v+
DTr+FZbvqhg0krPEmasZnr/4CpKRU2BSDNeU5pMYX7hfrzVc8HmOSLevz8cr2err
GNQOj+C5ZuwFP7R5tMRWurUEV8MAyWmpEj04jwGgANKp5qcVKsoTDtwRRYmrYN5R
0DWE68pZkSj4s5orprEqASz9UHpULXqFlXAWmr2lHxXSSkk29xfC2VDJUnOadP3o
SHb9RavXzChImNieFfK+qce2dFW7NWIHzUbhWh1PgTr4KDUDf2bXfZnmwEuXu+3Q
GcImyiV2C/H0GtzAkl+2WUeoaIfpO+GHXSpgUKTQSMBseS1Akb9lPLmEgvz3E6d2
wwDm94LMnrgvOWNoUzcPSFJtnf1W1exkjE0vi5irirpCUr8Hxgm7yagYLrGNXVM1
arHNDtE83K701olH8pebngYafR+QelypjdKX+5YFELb8mmlkLfeCVVYFwkvUzqpH
ljZYwOJTY6KcZnz92pNAHeEPw2LX2011ahvHfHLN2vOwVs1D0Xwtjfb6RqAdM35h
m4ayZLOYaA5FYAO22BfukTtMsEoV3nPvgI1Zd6mkL9kEovr1r74kJtpyzBQPx8yQ
UusBnbjXxfZtzgFLiPksbZDxQU002tFB41bJOpXXIUFqUg6hBMTuWlzJYCYv65zu
/fEjNtcSiismcV7/f+fXhL8SoRLOOrXA5v9ui1SgUtlNpU2P8+ZOQcqedUTWjfxR
k6o2IaMDnaKl/o85/O90c9EeRVUQ1cEn3rZZOFLOFqcp0zTOsTbn7ZKjDFwS1Yln
0AKEtLcEjgHlHpXSwCPR1jArWa3gxa0PwmNIsIM945wFxCKJZwOC1umdtql+lQMJ
mzCgEcJX1XuwgDqloz/xtVHCSRkrYmfZAnZMZJy1L5bM84MQAUGjfr1+5Pm1g9H8
yEgQjkLJngD8DKE5340zumPouZKEvlDm0pzudr678G3PVYabeHRrVh/IpwqLq0LK
6VZ66DFefmSaoBIpX9pBORjTN0FR1pPSIRuVvSq6yIFiWW53RG5BqOzKcR14JDZO
/BXRPmoxCyda+JV77cb1qUEfytohgReTewjSMMEOCXgmoNY20JztFIqiQuErYiKW
GYF9URVU0qE9N9VDHzBlBMKpUU+JhLdU+SlNNgRMWlvgf4e30oDgcLqS3/ZToYco
mM0e/5meGuhXJueQwvBNMi+9QOfMuWM690NagihOCix+bkw+FefTpQ6wM+RWngu9
XRaOWPTqb7zjdNTfSVueJHbWtlaaDrxjaCRraaOUhUA2CucTdupVjzPyvKeeluJl
kkDQK6FZ2a2AC9VDpYRz9CuKl0UttqU52fz2I/hr7wfdICMj6XLRwAdsRbTwteGe
vQc5MsJZc/y0TmH3Bx5ljDkvAt8TICqiqGwYaXSwHIxuKqpkp9A0iugJzii5diW4
r9eXefwLXo04lHEafZoFn3oTvkuCHZp/pDn2d9SLmOSKwa4WsbCLdlJ3d5GDDRRi
oarqVxjNPbTAX0AtK/8oip9oPuCxzq9vyc9kUYY7gnLmkpZviyQ04O/zYgTqTgBB
rsBTn6c/y4Skdo5dpvQ+DSrUXcI6wSCD2mmHMyPvTGB5aAX9Sx7mZxjDwxZ0aH+L
QjSkfz69sjH11jfZPYslX4xhZP95dtwxR5Tob5ntB2yQdoMfltaPTlAh4m+nCgSJ
YEZVAagOeU2oxUb328UFxZVyUEEL2vM9BDuD4UUeU/6I62iULnpwDj7vx4CjIODd
5gg9Row3OkiT47p5ElZUmDUEqOjQ/salF8LcKDIbnmcVTGDPlr9iJuulYKjZjbt4
A+cvDkRuAGui4AvGdBbUGNtWG/o8AmV4II9c2QnRxAFPxG+KRXLklJpw6lT4yhnR
NkAqIycz9eg1mXzn7Rdk1/nizA9jsDpfSZwLYdO2/iawDBsjPMufWC52DCPtnsYW
p5KvIT6TG40/u4En4qDeJ/Ks5LSBg0r3brXeCAifVNgKgGoAf5EvZ2SUKMvuQUey
DGDlPSVfhyxmZQCVy7oPB2eX9TDSSF39WImi/oduap6g+zUYIG9QOuRrgBM7XHyU
Ji3bfvwH9k87ofUPabd4eDdN3SX3BhXgID8pRtMNWZQQ+xo44a3p5IK3pJ4Xhny2
mWdztySwX5ujJnMQqxslkv3eFcaXQxYpNiNhNpdz8wkPHO7CvkXNHmhn2+ZKbt+y
kCFkm3SHcuPuSubY7NdZp8QFBfnNQaR6bNIMMKD/svbVr0FT3iD+zdt5t881O3aT
ul1/WE5GClHY9Tp9XxajUo2qZMjU52i/3PHtQ7RSI8VHThx5empZpyyOqtTVuPF9
NhBlsTsy3RVagMyyT2w7hopimraHvL0XTJEIvvdYVUnmEIaMmrbIkBzHpWreDAnk
RUVuGWc0/6nMt1Wx/U4gtqe0sNMuFUwjFK6uSNGNWcVUkRU11PKDS8jIZ3TzML8/
0er2EqmLpxuvtEf4CWVe9Rj2pLLfNDTxMhuUOcqzrWVvkIXf6pK/vWsR7GvHAVY5
hUoSmnH58xJ0iEcNvWrhdR+J5PP2Rc1TCsP0cUFJgTASvSMvQOwatwi1XAIUzT0K
HHHQik3rVyYnkSwx7r0Xa5iVBvgGPVRpHosHqpnV7KlTRNTT/KcamOG77/QrndEE
m3plUexxzgLFxhr+foNKFUWVnPpyXyZvV9ttgwmkqVfX0t3r2rYXCfipsjTdi8bj
GeR65YZJWz6dvhSI1w30yIhyw6M9DbucQjXpPF6IKnCKnrxPhkMnO1arO37/qjlx
NLQQQAVAb5WrD17OeYYcoMmpU3HhYe0mVOEwVBli9aOozi+2igSIHOYFnxHN5Hdo
/NGnlz2i1Fi49ZBOVUHqLgx9I6EsxwrYy6npMyOVTL3G/RG//3oLSLUc5YiwJewJ
dlSij1XAiDj428hGyGmmc2J8utRvwUylw7jvZIOovwuTp4MomLs+cB2orTSpWk8y
LtG/EMSwxDv2khBP4XXQfsBE4kejFPgRxKkhmUg+sOGxnrlTDlzLdEYIpNpB9aFv
F7FMqQ+eS7Nqfl9on6c+01rjvK6J6z7b7H6kVvZOyL5fo+kQP6sqe3mLQtMTJD+e
6ga48F/7lIioEDyaxqpPC2mRRihlMZTX7A5veqxXez+lXbfDFcw/wo8ciUuefSA3
uz3OBemkyQaxXfkr3aYcTLympGwbKkKVxKV3kP0zAYWSFHUan3WNALEaAwK4dYv+
04LirOOEEnhXPYK6juEEf2iexUEy9inB73RN9k5H2+PWfsO0QcmuXRqU1HTGwjnS
`protect END_PROTECTED
