`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mC6XX6jK3KVJrosFgHQ6ZDMO2NGvaa0GdVQNDoBRUrckA5ytQTnjRUI831C3Hb/Q
lbRxoinEAvgGKD0RRB0PTNNzc2bfMMw8Y5jPt3mU+oF63NgREbe2R6PIft/4n08f
csXlNadmIFc3fD/TB7QZlAV0IeR5OIJf49mUu/Ul7Ic3EOjtXgeGkgoTIdW10Z1v
vSd16f76XwX9Vkokw4V78s9+qAkb8haQBl97bzbFtdyVH+RTc0ikodytGZCvUckD
dl0C/501vKUrXbXuIkhyqSfK2C9ry2cBQoEnSTSHb5n2+5BKv/nxtteJcVkn16EV
37gN/y2ZD6EECNDPSz6d4B+WrSFOVGABHpXBWIAhhNfSpM3kMrL9+J+yLKnkNxr1
zoMYWjHYfOrmr96WSEzGXrqhnBM46+DTIlCh0Es21XTqY4b/HdzTA/zSLuv5cCbz
epOor9g5riYat3oR6MwxTvlVGLTuieD2bchyJD073gaFacu9+0h9bb2xDZeqHLg/
Fbvn327czpKX77fKS1dPtCvdvrSaDIzPCqed1rwUGs3tHoJv8R+Y4Pa74yqwXqJx
MGIgxrSmHgmKgrzdaQrczv0nkgYM7iiadAAl0Ly6YUWZRMGjxFe0KIKu2pxa7j8a
BS17c7wM1NSgVDfU63v5cq0biL7Wk7zS5SGsTQmebN1grhgPAzxt9GEuDYj5mkbo
HzwdfA1AXuK+jak8F+zjwtntBaiuOWt1b1G0+kAm4nMId7LbBf4iKO2IdaT8FSos
izlCNNiOZ9XIL98+FKhR0jbmKyMUAD3cZz48cgAWhWbt/vz/LGMbHpronRazO7JA
`protect END_PROTECTED
