`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ydHDayngMi2/1LmyKNy+jED2+aC9XJO+TfVV951DfNG9kzvFB+m7M1o4pYQozz1
lwbeU7If6Z3xupIdQObx4tnpT83/sRWQvAZ+uICwPdKZbTBC9VoRP8MwUPsTZ7oe
pmXGbwyvUyChNW5gJME5dQycbvB34u1kygRyyUfxBlEWYj7CBfv9F+4uuMMAFE/R
tfwaNuN7lnb+axyajBGFHe0kLR/QM04thlbZXt6nfyXa1nVeH9lbn+m01U/4C7/+
iuC0UiPcUAO51CeFEyfIddP3jKKH6Djo0mkM0Y9OfTmlMEKiLj/4yZix+1nK3/Ha
rs5sQOpWSdTj2dHoRTboI7AUQWW+TXp9iwOOICjUqsYyoV/EY3mGCRR2UPFIQcOg
+rI6PEJw+MTh4Rz6Unn1Q8P5IhzSFwIv+uRGGUEvrwuWkQHYV9SIR78hh2Lyvw8r
Rk1X8E4zkeSuU1WmyVE17bR/YkTFjq+7uzpj+BBFIbigmNkaUSdvleeb9Q1E2KiY
LnXbVBebhCEbbga0P/SjDnuVLqyMDcuRkbCUkRprEFtATveDPOAk0aIQAKDD7iLY
XgZiYXlFq4GcVg/qPPiB/z+h/hweVlqCBZ4m5GEV0S+1OeWzhGz8O+alkUxduJdR
okk0mD88g3Vau4oUi8Eq/xzfdOfydZPwEYDhK055ES9PEkxTZQx82nlz4eucUcya
xP/MnlI9Kd1buOq7qKu1O9keGrdPwvlCKRC1XPF0sS5VAqJELN5PbyPnT3tdG5B3
`protect END_PROTECTED
