`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPhL943fdPqRbbrQhcKkOIveOt2ZoVeX/+jIJfBSzChRD3qBkTUZ7pMle8HVOBkg
5JR9p4VDZ3+wC7ohYEJw9k7Mw/KcKS6dpCJp+MA2J7IZZ6BqWsnuNAAaWf86GqVx
HSdbAoq0t6AnkLHQ8+YdbAqcleEAzJUnGHQEIXKNjS0DmdKix/Oxv2JEAMCSqZr6
caqvs7ElMOiSNRoRMfW4D9LjfiLwWZMT2AOqSRTNL1m//T8vJE3JAeHEAFQzABBK
wRbk1an7TcI2x+t+tZLdPWrXmKsK413GSwTbUltyArNdK8VKIeIZlbUE6i4pFQcY
3ngdPTmKo3zrF+6narz+hzh2hus/lwOfybRR8kULkNwN5rZLsB/efwksL4i7w5ov
lNZv46TDDHnlwI0D9EEPkWoeeXBtpnlxcmgJlf7C1jI=
`protect END_PROTECTED
