`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvh7i15RQTrXhmNPS5ln8/FQPUChmLndbqfodAE6MCca+1wuQGjxNZ69cnyELVHb
MxeXgvSV+Os30sjlMlWCTM2+ALm94p1eVJk7WlDcmjR3inl6V0YwO7V2nWLQMjaJ
5gyqekX8hA5Wu10MxU8/Mv0P4qYUBrkscPRVGiEHBwGV2kQG2RpWu+ZGoQLnN6MG
+miG7YIJckeN6ZW7aoZc012tjI6Ovy2Vw9QGzYumgjhhq1oqhprx/y0fC0qJ88ht
tLA6twarG1LgmdoAHhzNTFZtDcm/xJfcdi3pGExq3MenP04J+vRrukuMqmifdHnM
107mP2LvDNcVimBC5RQs5T/sxFirR/ma24qHPULCS/8kqgTO82dtwLn4QU1Lf8Im
r72KyXCjHzIuUfaMSvnqAn7wTqlCYoNYMEM/sQo4tMuiVkrcwA2dxM6nEtsz8jEn
32jA1YDIecWSyQ5bcF82KLElJud/yUlc8g7lq4pXSCdiqAqu1Sto2AklHS4Lixy5
BkuSa/KFfoayRmA+iplLRL1BoOaaMfMzvvm6NshQqlh7XySl6q0U5iO2mLRTiQbf
oEzsoaAlYT+r6jWXjNc3ZKM9RsX8Fj+AlQyR8ZHK2asYpkkzY67ay7uvqxsv5YXd
iFu3EzNEdOg/qzKDluH6CNleB77CjF0g9mCUNHN3IZHDzlzCHEU7VyCSaba/5R2D
mSpYLdUfsLgAhawB+naPb91czVNv8oaIuNfU0RJ37nqrNjsc3PHxBJnFoZjlSq2q
NNHf4l1JHusTQeOmUe83ZOPyrSdfbmU9vkrJUSwCvIM799Y9Hy6dsJYxmy2P+CPe
L/UgjOGYwJleCzEFVcjtvs+0qZ+9ha18c26iNz7Dgz+1eqQHYVOK4jkRmktTPXNz
IaMTbrmGold/CfzgZmKH4AyHQRfmYbLgBq/T/iBsmFdIqmzn4zBqGR4VKvQpP561
B3008gnXt85JJl4bQW6TzbLuTUrGqSwRWbbo5suJEEk5WjqNJj7Y5DEEnJpjRTd6
dZdbPgf65XqPZuHex8JisxCv4xz9houdiFQt7eWbgkFkGxMYtGnV2fP++Nh1xLt5
mnnaNeyc7AFsBY4hxcnGNTdC6dKfXeVFqZxnr4OngC6zzKTcpDTQBbxjOVoqu6Vr
Yb2ZnPrkMc7QibSTqpr2wPgDpz/4cb6snsza9vJfKSgz9VKfGU7fv0/cfAr1tmEK
Wus31thwQCgXAaQr1RU+GmFhLEwANCkHirGB5uyX3YfJ+esQf5A5xPTV1a+Z+50J
ZJHfm6H+Vsk42o5KVc+BVzQeSzCqnaBrKMldeXQK6exwRcFauGkX7SRaxWq1M6MB
lo5SM8ACLU0RsPJDfYX0hUq2mTNHZTnntg2TqJrdCPkVcYYCH542ErVVO+HsxRoI
SH9ztU5FlDTc6Sp1ruN3fHFqvCLTwjvBByrRb6Oz7OVvgcOSVhtfQwQ/k98kNvF/
FXBJQaQcyjMD5G2laULb9S5wthyw4U4DCV0FFnZ0eHRxyXB81Ys/Pzk7xXuzQGtX
4iG4SfevX7balRkCcyZklBBFV0ZGl4jtLdxAbGNb6AEUVuIFr798+YeJaE2juqDa
Nwj+a27POlKzz3dBfdo+pWEkb9FWzzy5QTVhz1udDpFAbMasODKSGeebFCw8uCu3
KX2HrmbO4r9fRRBUxh36rRWJmAlntxEcceEtzlkfIYHDuSGK0nhY0wsRaC7HNhf2
bgxofMZCT4SgtQ3jhPsQ89Wq8Zkhbtk9/1nD8IP5I9FmU1QM4Gy2HbDcPDhL+vLK
EyVsyxBtrq44I9AVYcA86K+P9teXNI+RxG3v7ibc80CXzz97lbMBIzXMOobvZH/e
c0WZId75a0jYZ8lekWvPh2zFN/7qlvh4kdwb0OncqNE=
`protect END_PROTECTED
