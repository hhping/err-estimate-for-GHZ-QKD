`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AP1Lcw3V24eJBLq9niAGDzdeS88fBvsi2JXCcjU3Hqussm0MUo3thwX4/ptygFJa
9d4pxh5q52S8fQb3YxrjIMyk4ikNuVnWuZ96v9VEupTuIWvhpYnJVwqoCrmm6OUP
3GdiLuD6SnMX4J+GIPaNb6QFFmJJlyhxFte4g/bRKY+itVrnMB1eNEcOWMQPDagj
+6CZKv1o+0bPDg9J6i/2U0luZpdyX/hu9/oTqRXc6cLVNlrlUbIPS3es2ToC7VjL
XIEujJgHPf3mjQLG9vZsXCA+uz+F+TnJsJlag7lnxgIa0dnqI5o5rcmQcoNrG53I
JJQzTs/Gn6ZNZYpMAhwZYkenXcT/Cnlye8wnIyBp/bVJHS8ONbHcI0rdnWfibgt3
iOxLMZgMgUbGRieVwfyvO0JOeQ7S89mRJDhfsPoy3GG+c9j5MKj0s7z1sFrCVO3d
bxfMyjxTSh/2TFbZj18MPCnQy9vyhqkfO8ZM5jDTBUJNp45ibRBX6M87JXUCEBhs
tE5xvEjNV+YgbGaLVvGTniJdi96exwWOL9J0TnwuOZ18Ei9ssQxMWeQAYODevGPU
WZuDwlu1gFKyiu39bPdqeKrN3j0xtdPERBcBdzPHXnco7draNXcNCIL3+Atq6ClU
/2v8wiYs9+Jg6XUfRfk0z1xU9WmQ55i1LMgG8XvHOac/hBp0pjCiee8IAHZ1Ict3
MzRlArreT/NaDalcGB5xHu4JK6F9mt4p2gsbtnJq+T3jxkywDV4lebvXnRviklS1
D1Ou40JEbdMtCIGgAVE1MtylUXcPlg/wedqSe4n7aeJnY7DyCc0WpCex23OPNNho
gSSCfTMbYYeAzqCf+UXB/Zw280BIvVyHGabR1zp6q8Lr4h8M5zqG/lvT6xN3qB4j
y8ToHsopE1l2T+Btk4wvyFB1AMDiLuvm+FZig83DwpowXgyRuVN0keIazvkEvtQO
vvssb3IU6Amy0RI7kiI2nTnOtSP9yBBru+nlnBbCod4xWcz3pAAyUgKKOSY50akw
PYSyPYXFc0hKyKRzkaKK2mPkrWi+cFoiF4kGTFzwTN9XtLiPPMZXjuBE6hVWaXnU
uErYI1wWbpl+jB2wpUAnMyWvxZFbAxATqq5nms/2BVqc3GOkjWc/st3gW8RFG9tm
Da161FiFbOVlKqkWTCIIxfbQf/GSLjuuOz9UwXO/dP6wkYcnygs7jyoGsrC/IDNk
ydogJ9Uqcne26iuD23jXkIjy7RGNzxU09GeY7497bxauljcMDt/KBAVNP/Q2qX6d
T2WUahKA0E6LpbYOu4WjGW7xBLOYzWimQPAMjHI1fx8oe2xB7uU248giIkOVcizU
cho6I/3kx9xgsALdJwhuUxrqqrmWUyNkQzmwZD2uD3Ml/c99mzjRxeUJ1jWNESWA
RHbBobXTV6sOTiBj6TP+lFVO9QcZZ7EvXGERxFtgFVVuDcBZwmSpf/V65IhzWkVk
cptFiU7whvpB1Sc1N1pWCtcDTAXqYcFU4D1PajYtaI5bUMZ89zukHqtdFViuVhSh
JlEdT3SPQy8ZtW/7WjIAhRFE/8OJ0iSsaus3NLqyKUKtKw0Lh6M3v5NzPup9pXRt
Om6BvxtaKEz3kE+F5ZS/FPLHY2p4zCRcgNs6NylIJzRIjkSn6OLOY8aHoYibzbeR
rEPF4vDPcTuzy5+xJGDC3H5bV8qm4Z80sF7WATCvVYEHPZIzoReB6seeM7LxmREH
QDZJ9hTJKaIxu7upyBBf0jNSOl1Ke1Tqn6ZyYYcZ0X9rJw3Wu441TiwhM9zsutJB
EiKbwCyiwECY+iJa3JTTt632MkkejN95SdmdQ92JZZPc9xA7T8Na9/nBH2Q3EjN8
ul/o2VGy3QQeb1ivqDdtGA5yb3XYbuXTCoTzxvLYhV2RzITGgF4WCwDRrY+7Zd79
+hsy/Qxupg8DSQ7gv+SypXYKmMkCYJeXqg1otLrmR2/r/QiuE5HiQcV8bLRd1kvi
laejRssHxJLEKn/++S1Fv86532KgD9vTlEMLRLVBR+Y=
`protect END_PROTECTED
