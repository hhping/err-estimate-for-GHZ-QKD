`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7D/78LVM74H0SwA500LTyzbn5s31CY1aDwgIJpww0yYxS6QATmEAI2jcu+SMmQ3
b2jdoShlt79bgTS1tndXLe6tG087N3fl8Cis/9St6zbwkYM+FV1Vk1OvdlNZSrGH
MqhQceC9FpgsEZ2PJ58I/Jw4qirR8AEw34W8RsiiKNn99oiL3xLgcDqqy2YAohYp
ehQQ0ozPYV92/pWkEj3wupoNfWb/tBK6hqegeOdNx56nSmmQJIP8JEjeIp263YG5
mPv6BjZcYvPu/s379bOA9sVsMW/SgyrXNt1CqqNKK5n3D/Go+en8m5vbpIwWNQhr
vjHatv/C316H+tlTfyTQq9hIzdvDCTpe+LhX+97+8IcxpdI7obi1GzVfGlKviMSP
NkST6Ir06uA7rUvhisviH6Xb4avBNtQdZcAIaRGqkYcfsDuKAig/aJGWrJsBSB31
nvnm3/8LqX3hReugxjcpTfQo0tLhZCOjNQJns+Mwp6llXyUucHKO1S7qHYPYPzjI
6ADhtzbri07qWRjHZhc+jUtKINunqagk1mhWbh6Rv7HRzqWRmSER3CE+xdfImCr3
eYSeadnRSA7avVbE13IqU70ytzvZvCgW/nD0sZXyFvHQRzGsnibvCarNWojPJ9SU
QR/U8uIonFPnVx+VKoT8ITMOWVbWEHWPhHCa/rldAry4V3bxI3VjtIVF2MXnL6bO
nUcGBExatrg68nOmAHT69Tx0UQ0Er68QoLg2+iyvwCyy+xbcor2WoMNhJsoXAdqc
Hfk8c6RhBfwImlM/V+a94z3PNQixhqfw0M1wgeMOZ9huzbe9MKimQYyvrVgj7NdQ
1KCIKRU1j+SlxjiXv6bHBi52pTBdL3VB7Jr/DpRzHgtFLHSoAXjmSOLY5EJEXew+
zZohVo0zF7Aj1h29mO585ytbjDezoXGqFoeJ/eHjIwQUtt/N8XSZyd9g8jz3TDox
0cuxLM4nMAgD4+/u0HlY59h6NvQDLJ43+Vbk6mnOGtcexP55rYsqtdG16C4sh8Z4
lk+Gfn/Ih3Sc0vPU5/KTFcXRqTcG5dWi0YE3oyHiytVRpfFhLFjsRROJc1Xffy7C
WiaQ70MWTCa/zUdYeI6ygM659HGh0dAJTN9GL/Tvo2/E27+WZxqiD2ZrSD/+KPYY
JIrPl1geu2mvpRAQ89HweeRA/tuvICW0b8fAB4EKaU8/oN0VItvF1FijVic9Hbpm
4w6TnyAEZTPIUuu9tslH1b/sIsV2U32Acl37by2tzwInGH952N1weNQ9fRRStKAS
qARyR3+4y3hyJybowkpD8Smg7K4fqbfc/Cu4i24338rT2gXGoyYWiQLfnqQvtEHY
uSr8J5hfvzhcicdFVjjEjBU6XfjEgXFljYVIdimTQbfZuhsGqWIctsMDnDCzSkbn
SpB5Vrd1K7TxpHImWkOZtx0TAerV491Ow/SpB5LJCMsHbWzFcZAu5sj5SBDdt4wt
rjoQFh1guAOiuyV7IC3fg4C1J0KI81HF+ka3bEDboXXXZeHutdsBhtij7bb25JPf
XYOeijKwfpPL4Q82NsL4F/DsRfAlIh/oscAI33EVCXGxhYaUG71ZGWSVLJxBdJI7
u9u0r0I9ixAM6Ck2PNqXXl643gaz+j+g0Hf4UcuF/mwXvdY7JE1scuPkrgGOcrHP
Mg1EChFzuphoy3S4wbIxFibQ7jaI5ONgx1ZvYyAGVVYD3IruGoFOK29u/EY+UUN5
Y113aRnje7K1sGYT8H1mmlOhW4I+ezjiqhq0521/K+DG4cWiKYqUhm6jOgj9U/T8
Q6QOcLSI3aAoBnAF8YpPq8pmGO8ESYz41HuTC+nDbfPmb9OoazpSr/zk82G5pzS1
i55Z1yLUC734QYl1PPI7uYc/xXtP+o72VKlTQVyk5pkZlzYEW+u7rxlrvfxtx/nn
GMBNucAuO2DtRJHivV8b4P/kIGzbw7mnvAbDiL+Ds/1NBrl6VT4d7F9NckFKvQAc
oWEHkhhqtrC/VUkSEP9xyrOjEuWtfoREfWB3rfsEuQO3YyKWETd2jaBKQ8aG9skQ
VlQqJ6V7JOo3Ispc1dAZkl6fkUnJfoD9UaiQQzEW40GSdtpsW0zn1elVrePepHPU
cI7vOCz6o4BCioIQEtYuPbvjI9rNF0+InbtsahFrBe2pFtI8u57ue+ul7JUdJk38
LzEtKhkEsI83FhMyMHFQoOcuQ1aDB+R3WmUsLSzXViylPKPCtvoQaKIqebTDjRIp
xTnOS8NulOPNN/3XS7gOukShHbRQuyYn+pPhx8DgtUvCpvXIavl01Qonyu7YSDXl
WRAcwmVFwKSUpqLBFTDf40zgY/63TKwsT0dqKaReT8rHtvyx3e/FaJaEMoh0XSvu
O6py/lebOXegKL1kCQAJ9xYIl2FJVdXJqrEoj6y354YZpdZTVY45UUDENp1kB0eM
djaMR9TeWUq0XWCqr3TRpZXJK0VV4UoE7fXWhrYBZY4VcNMk6JBeZw778C/fDYES
TrKn45whuSHFJiV2jq3A23ysTLHS3KSr3VO4XzjlNKi8j5uAo6legG6Ld6GEchQc
vtoWxXb1F3kQkr8xYDskXw==
`protect END_PROTECTED
