`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21eGW4IExwN5UUMKElY2F4L7RE5hm1x9Wt2FPK/5hgdDeDvmsNFOsf+jwMIPx8em
gym+E9XfK8PSvG63imSn0PzMuouw9vOBNnxLlSzYPF3K55vuvqBhsnA055Hf81UI
cNgU7SAObqnq1KPvNkEjS8zHuscXulceAxUFx3TDkfBfEL4+TVX0vnMA+fNpOFH3
tiQT79DODMwqxgi8u36dwH2oqE1oRM/pNjlUs9tx3WlLHzDEjxvLUcfwgWpJ9T0e
lB8HgRgTkK8rCE+HvtaInGsvfZsLe+xlMZme2SH3g9xoqa0k+fzpsHY/UKgrYuWJ
7t8hrTmVvUjJBGy1uGoSXPYfM2iRwHzjZbDqCNLwZlxQzGKkj3U+inZUsLMZd72X
newiMKDUAOkEuxp802kdID4eOtf7uwcRjkJZREtXUQzpbAHWLlvILk/5F5v8xGNa
RyigibcfvaEUxW6Z1f0T9GNj85wVYMbSdYLYrxv+i+k7Ii/+rCBSMxg698BsKWDk
Kbs4ZWgTq+BrGcP9Tc70F+/8PkkwVv9Y3Dxh9/fJQOHccGezfYzdwGWRiAo+O85O
DmGNs8D7pqKPt7h4siQgEiOtH+iItCmbul/zNsGiCRXppuE77dau3wUd4m/avHUn
nYkpuyg36pTLVsHExbLQtNLIZzSMS8k7Nxh1w0sZvDLO1J988ZDncH2VPiNciurN
JLv5xpZHLph0duPwhXJ+xz9qP9Frly4WrYGh2PK28PlS9NB1gZf3nCWQDzLsWXJj
9xw0opRr2P8NxDMKzbMrE3Nr981uoIVNrq8tyh4y6MRLHCaB6KneVQLED66+qL1t
Y7cY+zZM8LZxyJnsiwGs4OVE7k8fSzBIEEgXlDeQ2FD48TOEjdP8jfsD8GoA1r/D
6kGm/yWEMxIXQ49mNiQsC0FJE9+UJGorBQmkbvKUJk1pAz5frkCrPg7o0SKeQNXO
aJ/+4+cFWjc55wcpwNaxBiVR5QSmjsbEnWZ6CICeN+QeyubleX6M/v3UtYDncVTH
iW6zJJpf3mXASj2EFbXUAlc6ObTZhgfsHMPubR6QkihqYC+cWVQP88hXrfyy/d3p
0qO5DjEgLeWCn8CrXsoj/BPLJB0oLaDb1rGufk4fpg5xxZmNkjwD/ZAzuj09UMQa
PPZqyW7Z+pKmGEcIHGIpfVFYt3j1YOCo4F92RdpKlEHAsseWInBnKESF+KtqjNoo
rOJIPm13/KRkgcUF0tOCyVjdduDsRNykH861Pof95vIBj9JVUwuKFhmnizZUV+71
SGAovvt/1lybKAjCsegP4pzT18NvqgfpXUElw6bAzpM03Ubq8BEGqDhvtfzB5Y0J
2+bgmUSwK4Qar2Lz0ufvlU0rZTHOGVr9Ne+8YKuTqU11mkJVnA3P6nKw+VZNF/4K
EfVgKMXSt3R9r5bIisW6OnbYATij9MGDyWkrRUfTHMCLvuqg9rdDSwDXWtKeujut
H95Kz15nXXyuATTxGlhphN5/EKPUUdVuvEvgAwXsRn454JJ5MlPOyiHAgQimnvfu
EEbI5YrOTVTZwv4zqLX6xHSRreAACKkH92Bh3pSW6xLL6TqJxa515+1NDbC/lDru
6nWWqzxfFXmMG0Z+bhgLpiGbHfYmeOcn6IdNZ2790VmbfxW9x08gNPpS60QyC8LN
JBHSczThs+8cxPQagFuA0dqTrrHMGWUzAM8WW3aLvEhTNvRtw/XkyDPVnytOS0FC
jUnG5525QnlT8b4DgyfxzIsr1wqMKIuOJBS//eKDF837Ii0b5DzKqxa9CQ3eP+H8
ibYwaZNpC36O+ZlRww4ewcrNl83ELy985FBVWeNGqdzjgVO3gFh1C+FFzF/nPLMZ
/EyDebvtxVPB/+J46BhJfdVcuNWzYP/o8qtPiJCkXcB626G/+gAoSb9FLUrXtLVn
65LzJ3+PfjaTWR1hmUVvmtYNVoLZy445gimu6eoLMRADTSfk+Dm9hd42nYGILpYo
uW/IwFvAs2evsifr3FDjA+dxET2VQN/eLGzkuIImo4MRzTU3S4iAXHPFcx5WYMkM
B0RHePjApk8pdG2xdNGwzTYCCJUlyFLpRI6Cz0X5wiXVptBOvy9jBox32qps/7U3
eR8p4VR+ysvHU52bRmMkxuCdti35V/N17PFOT+qgvzxjI0BtMLRFPWc1Jr36FWBV
nKgdPiuqHePZ8QzprnL0TjGCzDXk7UQe9syT50bMgNugpwi7pKGuAUMDgYC/bS5e
YWzw46//hfweIoyFspATQovKkGBh5bAWmzI2RuHkTxCrVteGS7GYd/p2BZ5o5u7V
lMH1v2/J3/uWBlznWpMoENY2ghzcyQ8cJZ/xpqImqAZOHXG5T/5GhpSgAi8Sszaj
OzpyzO4Vn4t0Qf5UlEc2iL26pcKkLBizt9k6Kj3rkqRGpkuIgtNw/wevsscwLH6s
8Rp0ZKUpj0lMJ8lJl+AmV4wia/q3nuQVBghuCa1c8kfTHHWun/skXL7YMsNXV+OD
bx+fzLJDvb2wqi3r8HLLUIFa7VnZ5pLBY5qRbPu4hkMv4wV7eOPmYJmec+0dKyQ+
V+SI8b2jR+lR4ZBv2DYgB4joazOXAJlafvmAI8uE3RjnUb/w+mVBTPr8Vv6eDWRI
q671mlHvtt5jlCVkAlDs4BU03UmnTsxj6Ak2HuLp/yrlFL8u97oN6TcbIIvRv24d
VZw/FDL3cwGUZd1kjHe3mq4zASdT1HI3tj0ANOF3bKe38KHzh5xHuoFRQOsbhhaJ
D7/wU5G6C+IotQdEDa8YBh6wkZFGPF8eZb4MtyWjHiVEZc84rOPg7p9Bn/OLu+1l
NxTXNeMcKR2MaMejULUTVBd0KmgG2apL8aMUcQPyMi1VfNOwD9MJRjHwm7wBfRgJ
NNB+pJZrDwUKoyEC7ALaZObCMgsdcK49u3ja7IkS0h/2RqtkSvL9nWvU9VBUorKr
Nc5atJ+2oYwbt7DGnN8UnlcKSZFOHy6EjUKTx5s8OyuRY6B5iwZ96y83MoQyUv0d
bYLaRpDzw7NUtWAj/QinKLzHDV36tY3JKbvFWoSla2gWUTNayZdppNj3nQChk91f
9Ju9KIiBdsdNtHv7HnHEi7xIN2kMWT3p4IS/KNO9RO7o0TFaIJsRBLx2e455Rs2j
QjC+JUhyyakN2Ouu44MAiZqq6BJZXENcExYbQ/5ppfKWuHL2PmiJsiknH/x3R9t0
o08RYWFFED7Sqqc7JDjMXlFZ/4Kdh3HMfECHrZ1B/45+fjZ67fUoIRj3uoLp5i3V
GOTgf5xQotX0zGhrWjXTIAlispA28uV/psFwWN1iT7T8IV31QDb4kLv/CYRU9qBn
RbYxdzmIP8FrdcFioepGGOfCGmWwa8GOTMJPQFJQeHaF/o4suyOOim0L4kvxdcB4
0aGRdOKqQZvLDWXzgLdWNYKl2D21oEXrkdVdAg7KfqUJk5zdXXG5A6gB9Vm4Bxcd
XgmhVz7VaWophXPj/FitAelZuBF7L6KNG9A/Hoh48xkGKMYmKtwpEioZGUfUxlPg
uKM/KjxwB7TeF6EfZlRc2FepL4jSm1kGu8H6SQyO1Suo4k8pye2pplzfut1QDfpH
O6ySu3VRDeodAjrhxBCIx9DG6mTuRX2Fidn4tqHPog8dYLhLkcxm98jMBEtRsL8L
Ataa82/khxByTz3AIsv+STYAQV2JZfFhMCnaB1pLM2srXLH3pJC3BrpryWdNMjBf
H5NAQtkKn2OdWIgtYSx3WB+V7WDKV5vSUa/SMfeuXuEPQ+KC7QVLcBNdiWfJikWW
U0+kxKPmMGpCmpmDD03CKvmDtOPmMiESxOFi42tfCUsoCcUKeoEmhl2Y3qxq2wiT
syNyt8aIcSSwpCJ+4PX2vs/+jegmW8vCL3j/cVTDSIUmIT5h5aptcjAuIhD0982A
TL69JgrCKZPeBv/0qGfIir1jHAo8R5SQiah2nXTdIFjkcRDLBRqM/vzLkXGt9/am
dnENapxnbHP9HzC0L0In2PF9p5UZqG5bDa67EOpDVhJSQpP7Z1vcyWY+tCkW9WaY
qi6dxz5d4IRVZ/Ms0dkRufSN5CYgY1dLdN/0+IkB5tLNNW6hW9s9TnlEwzInaNZR
24AFLB8VNUACOliJ85WHjP4wKUv295eIYX0p6fE91tbYtiML/ueQRtD5hzk+jVy7
yAU7T9KdFLf3Y8nwhNchFX75w3xfio3ItIGpYZ23RFD8F18Ko/a9vPkzWjg90IkY
VPY4Jh0ryqRyaa/zGkQDmI7JWir3kM303uc/00kgD2VwdKfLdghedzMvZP3TrVzB
Q80ae7BW1ifVltwz3FOfNBTrmqBoXpKDeihWoA0t8MuZh/0b5Whz3Exl6diKNl/7
eMATmMyOHt1ONfzgLcZSD9D5lCl909TFTY0N+NH44QcMTiUDigul56Vmtc0F+5HW
GFF5d3gL10224SUtMxUEIOABmyVIpyk81UGEc4M12S0CtXld6WsVBs3pns4UPI6M
62Flfc3OqMOrcHwOYH44Cj9E3ZfdhELODHvYzFyFcbKlEJiEorMWAvUKM3LURs9M
pOk34QcSloaJSULfEwdg4UMZYAPDhCITj1kHTFh2e/zdn1lGTv/oyTJDnjjaxlUY
uBI7uEh6C+sAQCaxhBLsOJ5KIG+XdhsML2hPjlgN4lapJkztXbnpNN+vf68Ci2wu
URYjodC6tWXoGE0t50u9yK6l80AmLpbSWKOmC5G4/y5SEpOaES8B7iCRBKeWB43u
oUe42/7Ka4lKO/CtW8KgYewUBmKUFHB2Y3dZJ7CANW2pUMHFCuMeIolvLx+DPhbY
6EgHKvJ7qqGfOO5OEPU9uBNh3ngoismwZes71BE6YT4sGk4oeWM1KfaEe3PrLXNU
9Rb6awXwmLp6h8bXPEnX0zPPpFJasZATV1VnfrYUEZjKfyZ4uEah5Im8V3NM2zfs
ET6hTrA4evKcOlQNiJ6W/XQri3Dhh7buxWfE/IdScdnVWN/fuH+mucJN2cJA0NJi
OXY9g3RkhqUGCX48MlY4beSltNSl4v/XEy/xCyYSv7HZQwnOmE3lAomkpHpyS1iu
wlKdfXpQt7hpgO3RaH5PHvjoBfi8FT9g2uZ7AOTlN5ZSiuHz91vgmahgY/gWsfRA
U9ub0aA2F/o4H3yCXOB0S3w4L2Md7sLoP7234vQm4Bdl42rmGb47gKyNFu5fuRqZ
OFoE7+990wHHGS18PnFdS9gMmlgHzg+jOPRW7Dz04OC9xUX1atRI9UY2qTh74RSB
J0xJDkWO3yBiK0bDPw18Af/9FYKDV6IbzbNshMPFHn0AyeOjBCjSqSXr1FzPhmIC
KWxqbFwTm6XVbdC/i3tPCKaVE6qmE17Q32lrzav3KRH4RgTVNfr4Rswdscn98suD
D5pcNzRbHggijeET1yDYB4qh/PHZuZ2Zq2DItuL6nJQXhqFX2+lnBbeqG0LP7Q6z
nVkVdKPpwtZ6dgZ2uJyjAFum3H4LciNivCVsBZ3qpaoBGNx54tBE0b1pMsB5bQz/
GkkEi+pNhoIyU/9tZs1qETMoVgzAKpu2Xkiw55mZzwd7SnKGkupMe/HfGlajO2Gd
XM98LtZA7pZ3OcZ6WOJY3iQiryU4lWmMEutOwrldx4OgBUeL9qa7Dd9jEaGNLgVV
3Z6Vn0PWpQFs9IaHoOL3ZoebEt1eL8LMOKgG+YQeOn/Q2tOGmZndiWiV6ykqIMiH
XqUK/+nO7yArD4zCNk14plqJi7+7syE8aHDys2SKVHBKLlq7z/fUxtlMTV0gD8B7
xVWQ310s7IU2GwvupQ9AOY9u8LT3aIj5csWFhw8UDfwXhkyqC7xXQaBRkuIddRKD
/Qex/fkRUEx3RxpcSBTPjNv7weg+1qcoX387FuOqlK2rorc6TYCEhbjv+ZgRMakk
s50es9KRBjmMoNEUUptk94GfhgCQRZgwaFCW8U3BLrZakIwqhqx4u+LFKZh6a3jN
mo3JIemGc8m4u65iMp/0zef3h03ApnA9/YzI8hx9FyDIXAoCOy7RlguguZyvOCDY
wc4zZw53DE7wcKczWukOgpPEkC8lQgYo9ORmQ+KraXYMWJGpywtklhSxZoXxRGUf
sdPqzqTJUYYvYQpHW5vOzu/l2GYRwcyHzVa56JHX1umcYafXp1k6Z3oqjU540GsR
oO6ItOy8AgpycRhICWEO0ByooYUeWvtgkUloCes1FgIcta3LhuzCW+/E6iJ4elPT
+ZYeiCQqbpwoU0DzhSrJR5grR5uzTBHE3hhMpIi2AJfTvUi1zgBBPHrvN/H3Iy/3
u/G9+YOQz5ZkFKr6TPIMGwVgWA2QNzey4snOJQ+bYg06CEaKMbQgQP0aCCcoD4FP
/dC2jNWc1Txn0N/VWM1SFo2PLc2vxOhxaNBT9Ho3K0dYZXoR8O61Ay1go0z3VRTa
wiU4tnsMVvTzJ0gcu0nRcOlmAuZGV4p5ZbEVOEW5Nf3gNSUj9WS//Bjy66FkmOjg
kla9ycYwFuRSeuTcNgHkVbuRn3zqg9EctTZeLtMz09K0NyvI/cDWKgChaYFmVA9F
3C4GYc4jvX0CUMvnYH2SPwazsE26gjfuDVokN7MvjiLb3PrjB2TUn23Zpxj9iPXR
`protect END_PROTECTED
