`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5v0rdpjHPMh7TVIs5QP2MHCHQgPTLWKiEx78SAxamqMEpfRkkZ7VTxdxoq56TnC
cRhDCL4DDrfhVGEGzDR3C82MhABlrIcjNA9ouIlOSZI62CiNqc/qFub15yiTq5+w
bv+AFEelMfcTpkknQEg5dKaZqW5eu6iLPtojh5rs09JG9DP/VBM25+9J/14eQfaL
3ql6cbDSSaOGCqcB3EGVVh3Mk9SwpJ8abR5cpD5/dY28581QmrT+yaOpB57fjz6w
CjXiabseaKKDkC8fq+JECX8f7OopbuzUkSA6QFC4AJ6N3sWhwUjilFm0TzuJ5CBG
ACdbf+ywdMcBkbP9uPDMzaSdld7YCHlFO/rGVa4t7KrefCI6fAztkV0SjDpj4hpV
6K0cPlDhQNCJYGyUgE7XVr2bg+BpzuyWJ6EaALMRaAsDplL6XglPIRCmZfBUIrwB
RdnySIAN5UpvdqNQe+TQjqCifB5M2yB9nWdaQi+tbVwBUZO3efSTwM/eFOgmsIe2
pYUx1usJVt1oAi9lci+e3sIUDETE279PGtDWYmtNREqKtHlTuWk9+0iFRsIrXLRD
lscSrp3CJtmhvwOiU7BWYg==
`protect END_PROTECTED
