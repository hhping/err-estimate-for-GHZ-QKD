`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R7leGhw4J2eF5R1RyupykzKcizVOOElO155uly8+q1h2LqMWSFW0ak0RVANOexnu
/17hJ0LZ3QNSDBasAE3rrcKXezWkLCqHQSv+moIXpbK2txo4qlJGouna34ylxSn3
ZiZe+3odR/3dw0oJm5r5s0mxlc7RCFpO6nno0ZXKHTrsJH9k8HCa5y8KVXFxhXR2
Zp+Er3TyZlAfJ1R53/+Agv3FwfiETNTElwzCjBZ8Fko97Ldaa5H8nu6hEkEv3UMe
1iqiKaSB79i6/eKbDE3qwa7G4bIIpSjbAFT7MuphONY82lzxqdHHRV0cPBKK0Z/G
03FzMb7nNowPr6utcdAeHhI8VStBn8KUsg0B69u4SZlATxi01xDWpvKWtgHfc2NY
488u35xhrmBD0ZG+vLjXl4smtuWJeVo9hoCD8nQOlKMDfiMWUdEniKoS3PIdPdcR
VQpVOt5/46EZLURQTXxNhLwsjJe3Mmu9Qr51W3T1yrm8iu0PlDGGLMAIkoNffvdn
l66h4CchBYAJVcJp/tBmqShh5VWVqh8NrT6p1+9nLJ/VproYrNJYDqqoJZQahuqQ
Zcgg8SK+MCC14k+tdMz1vzBMBj8FIl1SEQf4zk3wEaPbWynAq9sOtJk9jY5F+BuJ
nZHVZB8NTk9CJ4bO3lkFfmod+OFFI6EvoyBVXCVgTZ89xUOtuy52+683ELku63Du
Exj9zPYE//0EyOikRFl+RMxdzTwqNlpeJAACD7XzVVFU3YwQXAGCykHBIaxGePXR
bXG/jVphQlGhcTmAQlvyW/h3AR0riNxux9BTlrA/5P46DW1o9cGg3WJny27qQzGl
WOarT0xRAIzDaEA7YpXta1JAKYwWUTTvX5WRWrhld2fKyyLuEMdo3zWXX51Oa1Sj
CnVhGRONB/jpWERBbN910KkMalPrS0YA43APN+5XTijw+HAuyI/+J9dtWckI8K3k
U2h7VqKzKGu3UzySffYZRj9YXvLBHnilqi9EgYZiz+tPfXfKNs+2AIDykY4ZxAJW
4qfVcte9PisiD2ZKkW3hWVHqQl0iVQt8XnaCOvx/Kxq8dhJSMccDcgcwKGXUO696
VyLBefDq2US3F8atejYyt3Gg8599mDS5i0BsF0zZupZORgO9OacQS/fWx5vTTItH
9vuZwKPpZYpTcboldQNE4YCW0r3KuWCUWpECUkZGkV7gE/emPL358VVl4k93xuXT
8tss98BhXQZgUfuGpYjnKzG+EjL2T4vd7MYSotIgdxVF0UAPOVhDszrlgrdOBrUy
P/jcD4iB/dSWbu+x6gQCPMp4LfVWXeQZkLrojE0h+/boxzrnIMzYLetn2/pFltsi
WISvGkZ/oEljN8vu2jj/f49/p57/IhzD6vBHOzbGngINIUv7vpxHwxybdLugtbwj
AfzEvgWprBv0ZJsqmijJEj7LCoYRZh2xcMdOaLwgdHQHuiyAVg/jgDIjWZxfbZLs
5Y4Cb7tQWdS8VSrxVJMlaYcPu9PR/UMadXi1tDqBO/suumNxF3YMiO87RV4gI0kr
iRrN6ANSh+xhkgxlKMXnqKlXYASF8/wE0R0tR1/MJoSfVE71RkjPANHOmfd7XZ1M
34PseHL/Z1Jp6GwpmihUww==
`protect END_PROTECTED
