`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qj63gm3fIhXbxnuWACWAq7Wq32y6AKFWNlmWiocqw+pzYwbiEaM/wzQBTpN1QoLT
D1em4LgC/miYGNlxYRn82wa8dQ8pvhJdgqcjikiFJ4V0SlKnLLZcT3NHqAruLyyQ
LZNjr+F+OwaaS+Hg6LR+w98hJsl4n2HK2sGNRE6VzMP0HJ6GcglMmyrf5TrmGcxu
KZ2X7loDjLMqqlEKWvvmlO9zCmWQwjlMzMgxsXEQy9/aCRapOsnv7y6Qnp/XT/XU
LAmXVpdHFX1B4Z9OtDJT9+Yjbmwqfr2QHx2oTq2lhi8nHIU2SL+l60U3XWQGP93d
ixhM3iFR9HVvxU/sxIbath3CtcwULFDbFBxiY/M+shS7uBTsW76aTEyI+fEwbyxh
SU4Buq/fyC+1i4ScB1H2WDHLNKTXqo/Wl7MWdambsWwXZhGQW6fgOTIg5K9owQrZ
zRiYensoyxYpYstuIxh2PNnM3H3E7TNbf2uPk8FeMJjk447wuahtuf62jZytLGig
I6burN1Db8dQtgkMHhtyfG6wG5WHX8VRu9IAmiNaVVYdTYIaw7OmqLjISW9Gg1OT
MFDsnm6+apoGNmHfwzq1gYV+c38Z2E8sN9bNLzDxwY/LpM79HZi07Wrtx/4pulHC
DjmHP1f7bkMOyqoYwj0Kk646Myxc5FMxWYmPPa0pEKIRSTnFLE3lLLuFC/CosEkQ
CFa11fhPCgGdKp5IRWpvOw==
`protect END_PROTECTED
