`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLsNaByAVLAugfBjEYT1US9YbJ2e5mc1PSUCIadH9uUcgGZg98TomSeaBbG+eOSj
4WwVjGKAH2VzxRMkprUfaNKr4XsbKjacxz+gZTQW344mMk9omnOwW1aIPADE1yht
v7YYEZUdqBKSV2hYNNtqWHUV/l9fC378Eh3rrrRjedpuONxffznK8n6m61J5/3H5
FiEvmo14Xlc0//tSxn96k6gYENPkS2AJsKliL7M7u38cZynZVlfaUKzzlchH2YyY
gl3Ntlyug/8JMeKnAX6Utl8nBfNgT6DIaEVsbTJDQuGre934HBL6r4Lv///Dm249
yc1SeO8mDtPKT7vyDoinem51E6pXuTGGnQDL2eL8R36ngKWzPW+zUkhhRCcL/3nR
a+GMmi8gflTi2u1hDoqjvB2ukFks/U24v6KzWx2mAQNAyDKvp+XAPyoUwKbndrUv
7fMHnrk3pmiHVf1d55PKzkFjhF9d+AVv+spyV6jx58Bjq+D7h8otDyWx4YOEan61
Yzk4hD5B8dBHMOkuquaP2IzsyxEcrGOadFy8DnYzqGPL8anqc7hw0JZh5+MQ/TVx
LqDdEiA8ez32Upn8rD3uLNhej8L1LJh+V5s05sKaDnWHq+tBLcSC3dZrCLg+ZJRc
kxRXsAi3QzPjhOS/XpTIUvQRdt4IIFzLVTno9DtrphXm7bOtXW6mo1ZreMX8RfEJ
PCqWCBOjYfFiV1eZNX/Z36pCU8sudUA8R7GSB8UFWMDGqUfKEVM3vDDnvn8cUCw8
0MR7eaAou3OFyavYCb/97aRS6vxQCERTLGTPa2QWn7FENrB56MXVxISMzq4kjetQ
JfzwKiTxMLJT4cuIcuuQJNcZtIJLchC+RK2VQa7AB6RM49AQu8a813ebLEP4aSC9
NdUr+SfpZaIDj90HNF7N+EIqvmo54G4d75+AOwVjmM51TxM70jGHtrpAQfCilvcZ
w5tTiuDAmXH+BbocNrbNpDNUQpJrantKiC5/XwVKMUVFEWysDjdiGlteVR8ZP2wo
Gvm0Bg3fP7TXXwUCmjF7T7SRJXDWMM6soVjc5D7Qb+neRYxrsK1Y3/Vi1sTouAyo
/IeLYa12DbqA8AfN7NqmhTaZSEo+Snz8wLA4KomC1eZh9Q9Ii1UCRLG1mRiZ+exI
cfEdGfU+Cpr5/RsLEhBY8uQvwxCwZd7gzOdSSMPjDylx+sDDXyvNOaz+lzJVSjJ3
reWDFqvSJnfuHbaU6MLq2rFoPRRuW7j/7Ykwnar0NuefaFFF/QASWNTG32HlQM5R
ufEk5QKgOYsBCHgV6E/fqZeYIzZB8e+npE7atEyp96Kle5VygQdFCVkezajAetpt
eyeizivgWPz/y1I4MaGpEaruZkrrXFCx91yVVpjU/hy3QsRJ1G3QGUe9FMZLqFi0
teQPY5u8dcu70Lp5zzUmmk80j6QFFtET+jPHQ3d4Ue951WhrSLD/QwU/MiQAFA3F
5ufHu2GqfSwkobWQVMYw1FrTXWXDYb5owofHTK9y4u4wnjgG03PVWYv3kQNmG0BC
5mjt7yDtSnHPEPzUqIn19RG7b+o8Wf0FVQHBLBXDtlQvgOIMmd6r7/nlFSZHeE08
whHHqpvIjEouhIt/MZrERjAfyBFEcbSuVT6EfeUdQ/Oq4oAZgu0gp/0R9i1J7FJQ
N3skPDD44oCO0bQ9wuzt7e4CloQJVBiGCpa5S369MAo5ZoCew65efmb4tnHS/UMY
yxEBiDVtWdyaQANPtlRRRFHjp5DCkTP5AGYTSM01XhWh0M91GS8iaEoao77Uh3CZ
3s0WMXFKWUT3Mju09SKm4vANMgh9WUv0p+FYbYNU7t1Cp89xvmN7W2hzUD67tN5G
Fy8qxpODz72Fmp7JjmNIgs8QCyWqtSjBJ5enbpZD25CVF1n6d8wfjMx2hjmdxUjL
4SIqysOTktG7z7n6F533eeUEEIUD+kK42Ce5H+OqfHX+S/mAhQu7vhD4tJGN/2Ix
A/9ONEv+p6vWTYAltNaCLbT+qKsRK9PDYiRwUzor6s68HF581kyjTpI2OnTmcP64
wbIAcIT2dgkq3qoPF9WPb0HXgNxC45bwLYzgVrI7jnYt9nWCJ05/1m48+lmP7vJf
xyyVRxxJIqI2GjfMmV7MnBAyxy31vuN7iMuYNRQ5EcmOzW96Up24W+H8c7NAsnil
3aTxuGDEseC+fX2sTadAZ0k+9VhCirgf5mWCUR+QG/MtHPK4MN0ZOTaSFv6uJibQ
gr5CYHH0VpBSC81tYTb5EvUsQ5j3u6crv/ZJ1ArnZOleIZuvA590AXkiMmQGYNCG
QXblaVNNwtP6AUhbeLu9tQsasRdECl8MUXFHn29xvBM1/y4jJhaYPdo7IIdPNAKk
JQBM9kcO31mewjCl0FBtXs9CuPd/7ZR7WpE49sZzxH7JGoowiJx9yE7ppNcIt30g
vsNbPAfIuV0TQIGrdAukJTcnR/FonCxp3rweZUraQKOnFEl2wAMgJd0nQK6hPBhB
Ur/hleSM7Ye7XiLxfrEidyj8VHzurqFQ6YkmctQSzbauUSv+gn4ha3qY9uZ5jEPu
1Raw2WlWQ17tYzR6QpgfXK+md+OJu8u7E3l5Sr5Zu43FSwcymWvvj8uFdQvtQxf3
KDYfKauuZB5UjbrK9zm7FQbbM4AyLZBpJ9Skkft2PXDjcL+h3Bn1X2eGf3DT66SV
jT36lvEvX6eDONqPx5DvNRS6XeeybgP8qlddJSpuaiO4t4d28RUFRepfmE7Px0fI
ahk37rrpehvz0Q1rodvR25h+O0g3Es8fkVDLRTSycbMebLsefVuYI5FYMGEURoIM
R/1K/P83jonUUESU6218LEJJaqNJnhoDf4cIBc8b6ZRBVOOdCYcWR5fDpcM+FomC
Gb+s2bES30jIlnshPl5ir/P3s/vonvYNB6hlDVfWE6uhzkl4uR+atNdAd9wVjUbt
1OfQKaAwxmInLHNbbTfdWFNNxIkRR/8xdGjmNKd7T3VcK9fLNTYR3Ok7+wtdoOgn
JYqNRNLUV0LJmWGZ1fElM3Zms9emMXOBOUZwzvTINwf9tATATpTp/OuDXSQkgJgB
tvhketvKfEQt1EDFZWMuRCVEinwi1btMPedBobY6l+mYOw6sry7yxTYWK9CIc0Rk
mNXrkp5u0bW4enYlLDRirB/ZyTKADKyVEIfjZTMydi4HagI6zVf92v3gA1O4eP+Y
uAX3yq1ck6Wt/BoM7Si1t/NE44NGc6rLwPOA5oD+SPKM4AM/poP5AKVbIv4z11oR
8abwzolSYh9T9KYSIioIXlWVv42+E1h9Ae51paVtf16P/UsORqR3saxfBye+Y+i9
jvK5kLGlGAVYpLTg0pKqY1IJG6KajRDlzUg+aIAHB/wMhLVx4wjjt2yvySPkkOrN
7belYmlM2NxYB+TOvydhYrFvLcq5EmXailjG/2MKO7o9+D6W0ZwBNIoDAID//hvB
DIKJugHj4g9K0k2y9jZN5XzoBzgZjvo921psAzIIGLpopLgcrQshUcXYbRhf4YwC
oiOHE5C1mdTfyN7Ytq78xCZC08vIto/VznCMr/X+gFhbN4qAO5Y6Yf+dp1hCRhKR
xHANr8VqYCDA8lgHLUJydoY/dyznq1kXXBF3gM1lcWRQIJJh4rsN4bmuJ7xpCFYW
uzebce1JLHUAQwHw7zGWUk1PjAlwvyUX52Sb5ClLhrjO5dgWhrXD+ZVW4Q5wZq4o
HJSKNn65cTr4yKdg+tdQ98XraJ2bo0uCJkNL1Q6HV5XciSNL574Hav7j0vTi1Akc
gYGXRTP5bzwaWVbFl4YzK5vCdPgjA31PoX32D30sIB/K3ly7MFBiwcVxaa9QgpDx
Fuk9oQmc+WtUTU1NBZfc/21hqkTwEnPT+JpdkoKLtWqxI3+HxdoUula+AiTeLWfD
4wwKHuBoQY9rVPQ4ZC1kq30CekjFK1IGzFYni9mPKs29yGsEXijTOqYDX601OR7P
FbONclV+vLt5N61reaHOjNsYhXcfKRyglY7K7kLQUieTPhrop2iGH1g8mtDOgxt+
/BWDYdUgei4iA6MdOE6xb3g6WA8VBUFWl1TNWLkFsb0fBfFywBix4Wr3MMUFh3/3
DxRZX4bfspms4IyR6Rx1mLz4jW6MIit6Ypy0vUX9W6LukxPAAZKkVo+5LgR4r/9p
4yunZWXxp/BgQk8lVW6YDusZgXn8szyezfGl/HN8N8oL7t9Lmaa19+x3MKaFPVZw
csYs7ukBzRBgUg/4/qFiI0ymo5M9wVCSqBWRXSScavse8zTqBWYwl2WQng0X1eHc
VFh0Gla60vC6H1i4PlEdipibilk7/Z8HcRJEyieWG0/e/xd4ZUQBi2YPuerSFYNo
7lY1I6eaLTl8HrF4MigQrkfD/B2WasLEM50l+Mb2LurfOa7uT7M+TG2wyyaDtLck
37Tr5hkCPtiX8Wmm7TvijrUotqn1i/TUJK5cUfeP1evFeEyPJI8Urfvl9LN/PQ28
8MywVkH2dmoMr5mHLMxubYg9LZ99XcA3kDEUZppbx7eZe/8Ta9nPAtCPiEzklUrr
sI5rlQavHNYYQIWMVjQ6pff8ibRBVhowU5WLiHbVaIkG1D7Q5hMIkZCAUTAVHqPp
HC8pYMrPnfJa4pBMU+T+YB/nQldlZL05x8BiRKTdgw8VseXsrUVBVCtq0vxhZzNt
EtX32/Do12IXSfl8Ifv72B2CmlArzKoQyIlYReQw889z/j/tzvbqSZc1AKNnUZoH
h64YcaJ3dTuzJ35lXQmcypggJNyiOnAdvU6d5N0mFEaU9hWWEx3hiGz7rIqmTOFi
5HclktT48naCkEPmREA3+gjwdJBKbitTHyXtHJg5MJqQNt7sUeG+W/RQMrT1Iq3+
w3i6zFBOun26MZhz1XE9WmcjQCY9sFuhOSUygr6mVCVvru7w7JutHMg9ow3GDGxq
B+uKPSMc9ngEBnx4eDQzktJQlLqmp04t6i+H9+GDmJPhXVe829xFxYYrYp1ez1QY
2jzXjJHkVUwySV29aLUUc6mXu5sNeJZmysUJRK3xp5WlYyqvF/8tpsX6rH4Y50PT
Mv6iSE0Sm0e5JWKIrxXIup4HaYYwIUZ/VJxBrNPJjgu80h6yROOm5sh4VaCwsWfN
aZsyV5BJ4CVplHB8kuo+6d0qBd3cMKU2CtdQq9Hqts5VQcJMONjOGw7g4SiR1Ukp
+zvWn9mbyjePg5YTZFhQv52GJO1Mee4OHkCwPOFhnQmb1b4Z/1fFDHrAoml5uBwb
NQG5BwWFI9SnButtf/siO+TAKV2W4DkE+mQV/vtZ7nIRLXl5oiQ+Jp0I0ZjtiSVy
8qrOfTXv6yVh0aLystuVHYukTqbhxkFbnx3lSvCgjhPpOTjU3nhC01p64xcaX1GY
vxUDly4b4LiueDx5FtbR+QUUxqawl2J4KkaCZ8iJUzj14D0Fyve2DR4WB2uxmpyh
/jT0hQfdeSIamYVNb4Mwsi7cdkWKlffTZcbtJ752MBbdQ5xVT/t5UOMVBJDyQ8Xg
ouUuHuOXUPCVxNCghjLHNBVllfPveq1Wn5OsiqX6pWn9KAtdGicaoa3ZT26qaD94
12Vf2Enxqcjz5uZYyYcgPMyQxiWarU+ydSfAoax8ZsjyGlOuU+sDBA0fKGYPqnN6
Jz64t4qIcl88KW1kTvcvrkhB/oXIOfbf7BOsbtQ3327TkPsAyca9PpXhMFdxC56t
ZsPW6pBSwe8lEoEnBAn0y/pAnCl/2mSMizL+YLmd02WwaX4Vauio5/wlPFilb4pR
8pp/tDvESxviaB8XOZ8xBYOcS8WrOQvKpEiuh07qQn3kdBFcr0ImM7Df8Vd5m55j
eM4ezcbBOuQaEtHv1Jm5YMJG6U5AaCpvPf8wEf7RRK+qwYzwTA9ZgjeOfK8vcgm/
346Rr6EuoaEejQbWwg8M4rOCPivRfeJupvJrM1kiqmCBJA77gz02eCIlfdDfJozA
V2uS8aeg8BbtwPhSrjqWJ9wYgGWOE/GIbc9vVjxNVZGol5Y7GLEMGlxwza0oNYw2
w6HVzQT1hg78C+tNcdkYuM4PXFSVkBJFDFHIHg8I4VWNJAAUsuId+5QhBQLcRrYS
8Ybw8WhGF0AAgnOO1cHG7rq/sNKV6MrIp7lKZSFYD/SjGTB9Ng/Svinv49ms6spL
yLLT9QdFK+vQLOk/8nZV3sIIKsdjZ8UKbuggcaFouU4OoQqRV91/X6s+NHWWMsq8
F4P87jwSz6BXovjWkvBve72V0U1hD7JsfwVaPt4q0jUN5BNy9jhOcCZKl6hYkwAW
86clkPyt+tmdoFZAml8P7GFp/mRTovyVgCFZYRhPIwGD8m+ADp3hY63CZ454Th7F
eROavKLT8EPGIMMKq/NeYcBOeBHUUCZif0C8g9FQotwqUnsuDV+I6hfWQ3QbfyGM
Bw/uqGsHoekZ9eEktwJsZEm2/My1f62adUV7klDbbz/XM6TFbbf037uE5kDvi64N
DDACWts9k/4ZU2kDtBYllRxopYVGttqansqvg3lF+uTsTuhRSdD1xCGNnYSiVRW5
sYyjKwteqfwUK0uzt4BUjrfj76214BQzzllLWv95OSqhKgC1Ud++SnyvoqUDftVQ
tcYLN8c3e0kQ9WtwGRv9o9n21H+I5TP23vUmR91k/9HQZs3zw2c9g6uClXfxix15
r7y75l5ITT9tWHTbSOxF/Z2L4pQYbAdWqPpQkAAh23VAZh1cgu4kkQ/WvUJtULl7
HhpSrtmA2l331apPtjsjsg==
`protect END_PROTECTED
