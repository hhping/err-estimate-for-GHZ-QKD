`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OiRvlojpMd6TDS/MVPTOfmA7xALe6v3oIw27kw/hr0GWLMZV9/ZSorjfr1AVvG1+
d1Vfd+a6Lw7i5hQ3/hE61kwkuSDzMuCrdz4OKtRHv4iAGGGE52q+Gcn1a4IY5ZQd
jxNkn4rmWJvTvjE1/aa1+SGOyNshO6sUCDGjwuJ7pC+SIqZ/jDXS6P75lLFwMgTc
nYZeRfQIcxe7Dps4j4eKJldZgQVVQj91BizO2j1im6fEC1H/bC6YLckA7ojbV7PJ
7HqM4RD+TNSox42Ku9ETOJsvP86oAcSwC7ihqB8VoJ1NMeqHe9rX2wLkDPDAZgP9
HLXDb8WuvLIMQUyhYgCcL6v48IFtHDBctU5VRXWD+vCVxnX3UuhqhDgmpiAi4I90
`protect END_PROTECTED
