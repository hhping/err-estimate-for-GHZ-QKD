`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6RkBXBuS2PdmUHghJwfSlF/mamsBWIkXgajz0smEZGT0fhenAYJ/dxNgjKLpfn6
0DGuEjnfie0rV4ziUaXd53xbup9WbjQoylFzEerGfl4J/b/p/AGdVK9C4pCiMd2p
XcTHt4i25nPgOkAF3auGnvQhgTWWYCb9AIUWOYpb0UZ9Aut7ZuSmXZfMip7OsWDa
ocjuwhsJkydF/faOavzCpyQ6+rkkdhDQ7uEt8O0/YaRNOSRANsV3UUtxfOHpt6YN
DrO8pYQ33JQrpvte2OCTHyBcXvyYjtvO0pwFIznf6LBCqSoFJSUQLinX7RCWZa0M
hdvWbsesZoOJVPwL8FnhFgR6HSNTt3jdrIy6flZYbWn7O2M8p5reI4XEXWakBSy3
AVdSTjtHQIVEkBFgo0VECPPblyVTug+/mlzRQf2lZo5BoFFByRlAWpU/WvOUF4VE
X+xBMKB4MgFtA3bAXXgkK1uQZgsQpo36o1eKMkt2JgDhMFEj0ZdAnQ0VGbtbPUPW
tg+lVKUVkizE8cpmG6hD/i47L3l8IUiNTLkqjygRW79VFNpLs6uuFZPcuBkJkxbz
rlxI318WJsnpbRL5Jdbt93Pw3h13DV4pDi8moIerBVR9DaMW07UKv6ZuntSLrRIa
SEmgH0XJL9uN7sSfw5Id5AOM2VlvSQ8V8D6j7QnVp1RJcsfN3CYAS39Wy55ZPEEX
YjJ0eray0W65wca6Ll/fIHRNoLPHkiUAC7jID5SQoVRFBb54+Q2us7LSmRP3mrkt
j8hd7Sa6o1BnmryVIDYU6QfoIepPbWsBX7lwBMZaj3z1HvTe7kxPvc/jRPoF7Efa
/uHD96j0E+xSwMkvtKs4Rscm3DO41ozW/r5q0rO+zcbjua1rz67bONKbLF6qO2zi
fxV+tTMXgfgSlSdB870YG3GBvsr1robEsYDUNIyKc9KA9ADSHM5BAvUwg2zQuN+2
eoiKKMcWdhDeUNTU0mYnTOK21/TCCCvs8bnb1IaY0g4UWuchRR8N0BdXddNmeXDs
49fLSEgYonzFSsYbbDTRJuH9T/ojMU7U88laOITsDgTAADeAt1FQ6bgYjPaajR4B
7zkBd0tv4xLo0tga3e1smQJzOAzIrcKFdcSN3/1mE+qFcx1FKVW0ooLlanJf6kjU
7VlIFYxs13jep2W54bbEk5+Rh8b7zr/82uA57RVBKB2NOdj2zH+/fB5xskS6jSh+
IQobUV/s7rDpQr8mvgna8hbffhbrhwunCRPO3kaUNihs5OKu+nloNOr2yuSJ6lhX
eJlg+ptjqfvynosm0mZZinKlPI90JM/+XzLs7KL9lup+cK6IauI5rtSfIUntsDim
NFa36Nmfg5j2rINl5NG8FiwbixcSzIpEaKrRddPeqOUvCiqPbjn1LcKJqQFL/YVE
vRvD0DhZGuc/i6E6zorxDCn+I1pzAs5n9ZPe9t87T5uk75JpGKFXWU7An0XJL9QD
V3SMi8S3vWtAk6haqPx0Lyus1LnPKSs2/PEgdn/NxBEVaWIQtnndr6r3bAkSimP1
C7Zl4oiGJz52tqN1wngjRswhWxAUin35w+Hjyx84nivqHpH8+3Lr86905rkao7qK
EjHV1qAL5yCyHbhaijffI/UUr5fuFarb2yS/YQ+IGPGXCr5DpM0jei3dyTBXbClf
EZ3awG+Z9RcQcqcbcw1Eb5tGvfRhWHMRAYH4TFC+78WyfRfMcDXGfwE0EHk24HAF
TAiaJZUYZFmk2W/dIiB8uwIcIedS4NgziVMoZFMft3UhKxJLLiZPPOF9u1Ryu+ie
LIGux/qb/fzgm4YfbPqBvm0SI61LYGGC4j7Z7wfXgGPNtCipgUElFZg6hs5EajSx
wz4uJbGh5t3C2Dr0v42fgqtugsTuhKe0Hw71mVqMP1qnV0XBBJIPy0JLpsURU4lY
iWkkg07uE8pombLg/fjcbDvMF/GqCkVQyMV+AhNwIbxbZY5GQo1WNMnqwkiq4Qwh
1850WIy2fF9QQm2gqsgBC6/ocWt1jVjbKaUalfTNgSW6I5nsBpjqb/GKN2Y7yl/8
ZObNsF2ARUJZ7aADMflX8Ceeuo8Ye3622tmX6h//d4DgWTOdhz2BOttQ83NN6qut
7hWrKx2MYwHBVz/JvCCXGAHQJdgY56wH+mDEB/Et0OMKDXHBlMzbhYE4byUf+9uK
GU8eiUxuGBfe0n/GdBscbXLKpFjInNhujOn6iE8VIodlVyqz3ap58W0oMbyh0vMm
NK2P/PIGKv8HPrW/sEJZk8xS/nrWkvNVWNXHYNcJQWdYMIbs7SgyddgTNl1IBwLN
bQKCYNyklgOXcidkgDaULOA0CUDCwIocoqThirzlK27dptZGsKIDBLCUr+NJS4WB
XU7RklGf3WZXuoWtQkuTYqtjdejsaOeelH/cjCNWG4Mo/YXh6hVwliSk58+iwGEY
kPvHFpz1vlHSD/TdFf5Lku/wrmcOctLV6cakPjGH0b8MLF5KAibAdLhxbYr/+YRE
jPqoFa5GemIr2tc1YlVE1DA2f9ohELLxm2G8oDdxWElt0YMrPexVhiEhoNTyGIPV
RP16WyxtWHp9A/c+xcNQaR/gpNyJQAVx+caqRhEK29qLqKodhf1+riHScXv/JljN
mxlRAZbhROXPPraPH8gyX359U31DxbzMr3S4jdPX5b3IoQ7R3jAi8CCfR7jH4zd5
B4a+HCk+BUpkQcZEPo5N6ZKDyyNTZEtwcXTj4MLszmng+TcSkbjc16cXhSwKxJrE
c/6jjiHim9bgxCq685imVpAmR2BDXAUqGIV/NfYJhjtl61W64HdaCZ0ZdjPQ1bYe
X93rhL/+DJ2Zc/P0KEwxcxMw7MuNhbmtLOUUHx8BeFNlmxOic6fOl08Ud+7tI40e
SspGCZJHT5NIrGaU5hGeRFRMVrC9MYppEWcSxayDQ2fGiTdx/rpfYMvQiR6p6d2y
H5NGQsX+TcFFqp1JTPdbY9wYN7KSdEJnhNykR8UYivT8l1qHQvGfxf4Ze3rGcV+u
9DN9VxrZWd1aadluKS1YH6YvcCzME8uRziY5SuTL1670uqN0oEbfEO/ZFSTQozWD
dV6Z5Kt6nKBVG0Niv2Md0K0CVXmUfcM0su+8qGSyDNYN5Zz3iq3pN4GXAEKW9bir
/HlzIaBV5Y0MesJeyCMSx3VxV3zU4VAMO/ImaalqOL1rUVIMNpEbjcn/K+Um+Evj
+O8eH0kdt17p6VXE1uvEE3Q5htXkRWNJAfFPfbJ/z8de2b5N86xNsRiNUhRSyeVI
6TUzTtv1TJCTrJ1SzbdfvQYH1pCBAMN9a/8i24qFDcRiLsDtJYwxJXXduVpl7/Gj
Qkc8YUhdz9d167QCUcOWk0gy7vuueI4OkVRcjmgO9vfeKVIGy7Q3Xde4v3wj/byM
1+NKzUNiNk5DZIT0pZOcV9TBMgTDoToXnOHioeBE9VJuw+LznZhcKGoaEnvurlin
//+z7R6Nuja3bH7W4xgz9k3T/9dknzRKaAxTYfmczJ2mef3rzBA+JdgdZJBB8Kvv
MpQmhQP9V+LEMtfndBkkRZcJolPqm8dbjMXpCqFaT7QKrz44Z9AOuboY4Tqm3rYa
xyY18zbxNgqy42AKusNniuGKbJGinNT3EZw9xT1Nl4iyZdc0pDPCOsuqnrihnsP9
yFVfBkPl7ISgJ5uFnlQwsJsZPO4lZSIihANamdyJNfPLU/ghknYn2VQ9iBfSgvwy
GDH9bgeRo8gTc+3eOFSAkLZqIFJZDtkJKiD3PG8y1PxVn1be204o6Li4O+PKNCfJ
CjnW7M/qs+vxDAjyKpPnc2ofs5FZu8yFtce1KQTV78/RNo7Jcs32qEpVza51hw6A
4wG6Iu1iscDnfk9JAjO13OF2S3xKeUda2sZV130cFcfGlHMTFPAd2UGZalGpI7il
JkRAxHbbPYMg2fPDqpLlsPvg9u4tk1rxWDjll8rjNxS5Em2RE3V8u0Qf81QMcUge
cR1MsDzeltmaly7mfke4u6+AVNLp+Tdb7WOswOnda7TBkyBHB4/mgNCASph06OXY
Doou2Sya9DfCHkfaLkHR8D+4Wk/SCvah/k/QqCczXpRSxrh0gldgTuyoDjfuQMph
/qBAgUkW/1RXD6IFWEoh8RK7kXW0mjA5X530/Qlvq9gVBAe3dgafIk5LBUXePhIH
+JJauTsZnWjAd75FKbRCWsaCuAnfTj+FMuVYvDvo68hNenFterY1iKfH/LyAC8Ki
AS8bGu6PXWSXA9lto5S9taULwN+w0leT4wr+h4C9gGhJmL/iyTIuelgrvnPcEt/h
vABUz1bMlbE6f6sJ51S1K7xWEcKYgG69f5SmCdxvRD+NysNQE6b9Y0bdrXvdmhXZ
GaoJXLWC8GHxocR4B/8TntFpP86xeUVCQTl6cVsIMTxvyQdF8U9giNJE/Q5yq8BW
sI1WmV66jX+iLKf+v8LAzZlHxJKJowT+iZ6x5XHcXy0ahgmgl+vYMdOCImiuH5nx
1NDdOo4UNBjVRjS1kmpI0YkuMY7ddO9bVGdz4FnO3RiWifZ++NNNehBn5+/rLAG3
SA0lXbOZnIC7VA/6Lz67MTeDwbkpRXks8kkyMV7lyGDdzl5fiUPS+J3fMJsBo/O5
KSAJabJkNUm8SrIjkk7G4MfoTDoMI7ZlZsCD7lZ+xaZ0dCNSWEMVPfMZNOixHpQJ
TPA2gxM3MM4wvSWdWaJE5zalVQPOC7QgxLsUF13r3AVLq2REQIMOeDaDTpXWDS6O
CELMI7wfWA3x7EHr4ObzcYBgTMJMwOMBuzXIy6ORuhHnuIsdRWnBCiySPnnR0GHF
0VraPzQDwLEdy4yYFCF1kOkOGGD1ZlQDP5sIrEma1AN7aqM2/1B9miWWyebBj3ng
6aCgtqoQsV7TTq4PVbciNR2aOpiNucRfUM3oD49YR1asI3WdNiSZWqqv1gUKqwOG
vI56YOeWRsbokiP794fZh75qnMH9uq8DztMKcyt2VpoORHbcCZFUvbxPYEJHawsX
7w3HzthU4NeQEUM++bXBiadP7k/c2/l6yhknCo9rGBM1PyVvMMNzXqDhbbMwUcr1
yGAJJbYX+tbidzirGtke57/PVDwpa7NGtETLxjxYVLzIz4NFgfZn1zweiEsBR846
zVG6kKRjVGZLlsY1d5uILPAGtA9hc7Ch6MFKk+KdG0ynSjite/ANtgOLEbhRtQI1
TmYfZQ4fsRpdG1IAddCr2R4b8a0cNcwhds0vxyk1Q0yQBZzhCtovWQmULNHtC0t5
f9XWHMTxuD19A73ZmcD07GoYejkb7KLGPUX2qmCgrrxEO/Z+/xMahj/ZqLKJn+kb
dbrSFN/gRH2trpinsKMVlVAtaNglxHnZk/nUoil3fjEDfyfLDZAyOKT7rPxakG6r
AMe7oQYqz8EDmXZLuKwq0EMd1LLwOLAUdjTN8h1hJ7vCPUmlCI/mkFkMesAN8u7a
ZAU+Jsd8/jdxOY7B9AX+xYEM4KCR+0fUMoNEEBvlv83+N/cPAEbfJU1lCCcDTQMa
q9bTxzH9f1/SlaQ/r4EUYQ6HiFawGbuKXHZ5nVZVO1Cgt8M0fuOM+lNjuysAuEbD
/H5h8UBR0KK9RGYc8FDlDUgg1FPdoVA7vbwR3W98FRMDdAk6nqGdD5IicO6OV0t7
ayDsZTcRuL28GyvSiTGx9Me5Yw8x9+NJTL519V+lLNEWGdD1l9N5HIbV+KM7Y1zg
X8HIVYKrhLshVgcMHRNBoW+o67JIfLRcjCWTEBg6D1+QZSs8xFTh6FjoSxwaoFpq
AAS5F6DfqUlPJv05IN3qyDvSCR+Bz5IZkjHsfFDmFdMnVvKcLZJpax5+koyfgZPB
/ZK6+aqA4cNvBDxMcedE9lFkCYgVcWWIgWmY/fvMNssMTokJaNXTlgZK1PKnxA/1
VD61opUlYLmdu1vjqiYkTxOwB9HflqA8r6Ig2mryQFAoiCUeb5r4yr9txc+f5Eof
iiDe9muvDJ9u5joZfIYFE58oq2aQe8RgJI0aMavmZoZXpRMdrZXbfMRiYljR7UiB
3HiMgHx5KCNLmV0sYowlPcmvDhHok4klGomh6gC4VehyKNc/hf5LvhrCwkfW7MgK
wmfZNg16xYTZSzN4q3Q86Q==
`protect END_PROTECTED
