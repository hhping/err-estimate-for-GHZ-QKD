`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzoSqPEFqhnZpd526rxL4hbsZZMfX7gBTh9fJdOOv8EPVKS1yPu/cRC99MJzxwbr
2uz4gVLvaB0bqfiRq6rLsxJkRGs/xl9JFYEjqoTOr+PoMT5eKORnHtV9i3VWI6tF
VL2oW8j1Tj4dtTkrDQO/dARrBP2sVi5fWD/eQJZRyI1wizeQfTlLTmnC88P2wStN
JqpVsU9Gu2OHy3ESjY7y9TtEuIXBUGftb00vNrYOiaE6NvlY2chaEHh9kJi4M6qc
a+ToiR2MzC1kA1FpVIRksiHMiV73nLYFBor/HZ80kfOrUPo9Ui6ol9l7wHjdqWiv
TwX7WjaLYMjNVrH3Lny0O7v4wCSixbqOjq0MhwBx6i/VRSQbDOA3Tq3zkcNoOZ3H
waiGeXmKad5e9fEptsYnWgYdan9ZRod+hFM2/yVuvfKHdNCc1Ihv19/a5yF7oFzG
lim87Wjo/5aBmq8+fK87l8/ORiK8od2XSkmGrKjGqMowoHB8vyHE+GO/Qi8FKcvx
8m+KLOd8mUcKB1OCNdW0jWXFlZHRdJityLnyX/SPx4B4C6+DX5762Ovx3rkQFXjk
LIwF9zczOEI/+8iy5QlVAikwR5TsfGleavua9Ot8L+AHFvLB2KxEpmT0BTMGbqwP
TK3ZgYg+BghWAHv3DCA1Jp7QLTMbAgyYZ3eLd3IawRnjQGOinhKwFG8K3YRosUxT
sRj4kDTCElNTi2fCI8hkNultWqSTFh5gFLoX8sdy2++gjBlPMXezD//gIw5NSSF6
I+JNpAF34Kic5OfQw+yLGq0Ip5CBWRllpJ5CYszYI9WnIRtNq3cZbC9KYGBQJHu1
oBG+1Yb1DYlN3KGN1CjfMgo079wgdRp/gXvM8Zj8czgKmWOpAwBoEUNMoKQJPOlq
0FBAAzgPOINkbtD1RHGQ7xbSyj7AkQezUp/iR14crBp2NHAf5iQaDq96292Wx/WH
7D+TJgutpdPod0YXZHyZesRBUNCX5rbJawGMmFQP8FkZIztMGZv7t9Okf4B8CqE+
mViarYE0rN3V8FyuGlU1yQgPc2y3GcgCsZWhqgleYOXoeUS7rYRYDSbEmk5z2bLn
Zde+7huZQ+uP0Ma9LjsjHD4XeAKb21ro/LbwEHy53Fk4HBHT+kkBFoLVICdGtsQT
JE0+sT6rA6JJKqwKTlpvpO1qqmwXCq8BFW2qpd6L+KKDg42Qtwxdle2qDj4bNA97
lugweQmsRogET+l5xelfpMtTFOCaBXe87wpivopH/mLiOGhs9OykmwEq6l21NRmx
ye2EnS2evNBpdQRx4jp3LJ/lARXO/iQhCRhqkoK5m/kHpL5NI6z/BwzdOu84k7iy
/uXqu3JdsB/1hZxtSuZT3ZPg1SsV0SEhlpBRQNDLP2OhjJtL6+ORIiEuMnp403Al
klzFGxxmyKcwOhOI7o6LnvvWIW6P8bm2EmdcQXlViZnCkn8MgQ5D5tWr+5qYANOH
HkNOdX6wFEo+DA2FgMVAdY2hRFY5NmoDiJr5Am/ZDMxmhPnCA5/G0/By6EO1/YE8
MH5RI/Wadqjn+rkrtzQye5UUetTUnh3+YQHI7pLz9eKpAiyNnvNJnNHTl+f07gBa
Yf1Bh0Hn9JUe1dTbZpcH6UnIbroNnOB6glKsX1ULGz14Ra52NiEqM834vogzek0I
m51iLlnbCVGby1qaED6PFtkrxrKPjE1pk0P74I7JiJwawPe4wACuT0vEjRcxureY
In5IT2yy9N5JuwZQQVx3ZQddKkCseZ/Bq/T4CSDiaAAtPl5gt5CktxQxkvgiKYXB
0qE2ReUXX3ilIfJiCESxqmAZNWZ8yVIxAMkarShdhldfnrLNvroCdLGVDBDlp0Yx
kpxMmceOOQd2JlnPom7eKbmbU/R4XNRIdEuZ6t8NenwmY12glYpyN+WymtpXoIez
W7P0TrIjWIMDMGnzuhT1bfCQihD+RxYGer5J61xKbnrzbwNSk4yQAH13OdtXyzhT
YlQyBhXdI5iiimzHJDtMZVYJdNY3vsc9F8Hcvgg22V3k2rRhOEyiOIiXnKrrkmAX
f3RXFrZp4xtdOCs+dvYTSzz2e2gNW3GYGOn7BM7r/KZk58uxZPPaLnXYR0w/oaXB
2u2EF3nIlr9z3ok+Plj0ghluukUs9LOhUOf95uGS31X04l+lp9iZcB1SVioswLoV
PYqFmGxZ/hTzCA1tgGNcT/EGklOC3zYSeW1rE5ZI40ujWNtYh9l1UnjODbVA+EXQ
LpIDM9M+ZSuqHMJ5SGJybK5leorwk4zHcIndcGU83oZ/IUxa3yrhC5U6yvyVb5EV
dpr1lfQXWfSDoHvnzOQVxcKR+BOBj4H2J+nH4Ba9wUnHcPTPUfEBwMsooZ2BXamG
erKFrPyCY5MCVsNwJatCLzLVlO4+W7M2u4AyGaCWRfJ6vgwO9UeGd6i+A7z1ITf+
pDW3IujmkQkKP646XpPiuyHbPfFqPhXPbeXfVZz2j8EJsZc5kcVIaz5lL4Lvrl7K
PaTPfryrpkwj6e8pkM40VhcnZsQgsT4A0r4gDr/6lW4IsBnD8+8+rNlvJ22WnxzF
23gLo6VqeS3xuVIcW2S6O5JdKePVdKjLLiC3jg8qvCSXCm7rpy0UL4A2QWuH6BYN
SMXwPBEOPwLpuw+c//3KZ+99DgRSvr+dqPo8LHxCYYpbDXX0A5bYe9ZprbKB/ZCP
YgZlsrNDjJj6b9uz4gL9R5ipCZRylICB85mz0Y9kuTKl+80hnBsXtsEu5BL0+aCy
kb5QUdiFScmfvdZj8DrIB5yaeggTaCpld8Emp4m4fAkhHgrOK5CyP0dVnFhOZ3s1
RTDlrDvzJJFGS88ulzaTh85z3iW8DbRjUc27ArACKyNALJoCpMPszJ84oYLevKbM
SZ01XGihvKPr4kdPLKoEDt768ctH6FNA6/kmFqjuA+kWBRwELWcl48Z8YF30fevp
uvjH2EX+5Sz5RzsX/up7JUvrfzD0oj50r29Fathq8cxtA7j3NGhQrFkaYcLpzIDC
ZwFokQT8pRMfVfEWaxq8RAxfP5cjdwzubIZdYP2vIauCZc4SSYCi/o6y9q5jYyQQ
bzWXEc21TG2sEWMXJ02Qg0lN8pYl9z7LEeIcIPW+rR7mK3BKUEYHGbdybUAVL1yf
Adt8QoEcoLaGeA8+bww/WZhkfiKYFUbhRq65cUFDIY5g4Q8FI8pgF0HFUDLVLXXg
70TfHpVF1ZfVhrZQyyILJsCGlrST8ugtMQ6UgVe81zLUor4LsO/3fWmE4Dhn0Zkk
NjVllbgz0tXrwdHT70fEifkZnimoRM9pdpRFvnrtAOU=
`protect END_PROTECTED
