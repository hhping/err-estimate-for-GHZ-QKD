`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Q9pRg3vtq5SlEPTUkqdadFXWP22C1kGmln1+d+9ThrKXGie9iRv+HVH6EK7VoEE
sCax/9U48l56QcNxC8f0vUzbDMjxwvERDnWIwP8bmFWWeGgCVE7uIBf2lSb31Js5
Ehf0VowKgG2fGxi6vAGbYbn51n9CfQhH6cSYmFp6LYjJuwilyuWmq8Lu0Hze9g+/
RvOaWcJPq+z3ZT63W6stby9uyeTbTwlwUB7uxDRHE9IOY7YZ9mVgj7dMCQ2bZiOl
qwFBrjduUvg0Ia7rf7olmKBeeGBKfBY/6AzzB/114GfDxk3hhB4T/MHpM/MaWvEA
QorKNZB1V9qQWMoIyCXX8mpi6tzBLtfOrVSKcdt81zQheIbOcYlZZ5zMhSZXX/+k
mC2p0kiJB9FqaiFr4YE2n8u0mTFNF7zDww/3dYMBa5lp3onaF89BebIgflD3xGVB
gbubGvM4dbmd9yWwDYGv63ep1I7laUN7sdkjAfsveGwNOb0eeLTCwdOvuQOKQHcY
b4wGbvHWK8C+lBqEybT50+TpVir548rOHIfk5d4TZUkSiWLy1+dByPPwsR/G/VCO
AeMopZ6LV4xiR9FfEawXgfzFlDeVooTRRofXf71FURI5FP/XyTFgPmqFqXM0Ucq2
t9p1bUGz3lCkavNemnsGkLDbsebK9v1bLoh4zuGfTI+WHnsVEUqNyVnEzniYDUYD
1tKhw5kj7wPvVRgk04aSybXBvU9vreU4ChkUTTmBwQcF7hs1c3js/TgAgMRNjEcd
91f9lraPB17JxUjlea4ZXrKnwi2pP5TqDPW6g2JHRyS8ShAPAicI5YRvybQs72KU
/ZwubDJxuQgaKXaPirK4ISgP3ItuSennMfJxRydxpRThEehaVICsP/0vVUZu6KsC
`protect END_PROTECTED
