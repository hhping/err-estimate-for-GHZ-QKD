`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qn8MjOxGZh5+wKibtejFuHZMCx9/HTB1+HsTXeqB5Ym4ODrvfE3udPZ/nPZzqwMO
2cZqP6YBli0USACPOun1RETh+JvTDvYTxcEE64MceuKa9ojUtzmWtSTh0I8+2oq8
UDGyKS0fl5VNyfdI9/LzZk94WYrOndNVNprzEMKzpbjJXkoPE8Bgn3SQRPcBMp3o
eScOFksQ20cB4bV7JF7UTTZF/X1HwvGjUxQYaUUk8NXONda4ZNOGh/01AmhXvoBZ
H5IDPVb25jEk02oY3oJO7oD5BV7Zgn7irKW9Pm2VwRGnLfM0y1q7LeCIc2f5Nco5
NXl1MpucX8SHbSuNEORhxeht0WMvlWZuGOkt1rXQCSGGsGjm2RfVWOgHulS2/Frm
ShOAZEQPm0PXBUVFRYm/PWUEOIemTfkPMeb2IFeAV4U=
`protect END_PROTECTED
