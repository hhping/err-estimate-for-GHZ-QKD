`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxVyN+jQyEwMUBHJ55V4BKUqC8JnET4cIHjdJPe9ZB5w3tmJRDwmlmRamZKSfutH
BgzfxbJ4ryDKDZdQbEKJnfU5eZUavISP8VD1dsqkISq0UO1dVIjwXgpRrqRJap4m
lsinPxTc9WJDn6EHeZkmIEUdZGhvSi1YvlQa9dLFF702uuFKiZX0alk3QjqaROjh
ZruD9r06o0Z7/ah+vhADvV71a2zSIOvaWbu3RM9nY4xjDI3gHcYsE3Oz75/Gvcmb
CpKi4yRkLYNIsaJstB5V6hzsrjmDP3sG5B7dKAkiSg9GUL1kNeZQSUfmL1AbiUja
YYimk6JBzCI/pcwr/h1Ddi58VXIOu+CRIoFTeOYkMQUukwxGyi1kc+s8jNTX1HJt
ejR9mJV4zkBlPSVaMb77Xvyq1ghLzWfHSTrN3897XxA7oCMQ7ttIHGwJa1t5Gsa4
9uIy5E1s2rQqsehIdilXlIwqpuFxBeStIDv37v+I2gvlc720gzsGT5+KvJxsN/kC
XGeuuFDhuE+Zp0H49qQfcXp6t/Uk4BImZKgw8fa1NAb5V+REpqiHoTLWftOhvaaQ
V9ajAlvViaJiX7r7qhqe4+NJ05Siuiu8XU9zx2wzkDw25D6n3CywvBFYVgDABAO/
Vh94mZpIus3fFjN2dMgLfZGVDt+7I/nFVTSqCBLupRDIVmR2jTXteRC3lsD1Sy+Z
/l+VKMCDAvNhHog+BudE1RPpFBctHT4Z7mV23SxIMgVdDyjBqhU15V+o3zVSxi8z
Rgo4ievw5fXfNqU763hvYsE4ClsHh+3LrzGFim+DU92IA8YZ6ST33Zqzirfkpr1Y
GILkW4jl02x2F1gLIx9gveKXx/rU+t4pFIz4JryCBgooFucr+ntiqfNi4GiXHAxH
/R6YfmlkmU2mWkZGJDRLMftjlPj6qzZSML36DY2lDhoNzRCoO8Ekl3WIQ5UmrOEX
qkNlFjkSgZvwZUCMFGvNmaeRDOd1JkNWRf+iO3LNq9sLSD8BNU4xfUAJU0Nbu5Yk
8Q7dEnsXA7DYoHGxfR23GaZNtj0ilHqCKktX/KFWkEISHMnjKMgfUw2jaJfdPSae
g0afAU3pILL9jlV8reIuPF9vXfOHlKoiXAb+DClMcQXch+A4DSwlUTcBTqO7GIhK
jXlF32xNlHfSyYB2ldthUplsmkG/YXrMia++4H3yL0Wve330/h1U8UjIf5cUN5r/
zrQjtaZFhaV4qzIDYZ2uh8p/aLUunVhitQQvrpcoQ9W+W9IR7M11xNuoAVkM4uvG
CfpPvWC+y7UJubbNYup2FnZRgQADYahyhUXmELaONmhaQs1pn9dUiyykPwCltKqc
ysLVhJ+1Kjp592LApD+gYjWLSybf+DH1nQAAd/RadwmWNEtoaLu9QVdLdExBlNya
V2C+czAnf8seXSnE0XdiVpc346JWVK3zb96hcqupC5RLaJeZEvBSoTmUq3ZL8KDh
lSYzU4pEBxGEKCsnmW+NXFmcXD+Mzd1en1Gz48iMUQ6QhZBlUSU0BDr7s56Q6IyA
bNjJcV1EVkoOMiuA+gq9kHSL5Wrco3q6KXlegW1+UsReiK7ehGC1RYYIQ/zUYvmT
Q0yuVp4aDvDGZhmAUU66cmkrf83VyonLFLEgbuOhMaTg6FRkwlma6alhHFY3cnw0
nAaTugGKTmRvtH6XSUKHhQP37jjpit/QI0frk2Tg5+BB0f//6AuZOuTXgu5upoNb
vu1VUbF2R7/ZdVk6cYq5dNWFUSa+MWwixsXcfyAJrwooAhj4Qxh5LwZubuojESyk
UZ1L6viEEPkJog+obrwdxT8PnKTaGg4Tr+R07r6rbd7vzCo/8vGJF1L37TYya8vF
1gXJCwqJyjscRFL3NZsRDbXNDG8l9B52o4P31Jjf/fB6xk0eqq64vJOKaZFM9pTR
wW4mXtIWM2leAhvBd2k3J5XJjGIOauff7kUXccqmEvJPM9d3o3FhTjkHRUrnlu2u
zFsRHcOPSFCYTI1B3v/X1IdBHIQUNFtjI6k1fUMplQn82wesovf/PDcL9I4JC7Dl
MDFyN1lglcO+f77BIb7gbp9eRnG35VTSsin4As+jjLLWj9/BhUygm3oFUFj5BpvG
BpQMX0EzJku4x+8KpR1AtFm8t8/cdTb8sGyoY4/jPYVFRXm+WSRDsorEjvAlJVWO
vkeHCpchKYQAU7MeQiIQJUTTGFLcOu5RewvIG1aKxDH1x7/DCHeps6zXY5giQevh
WNQfnudAVcvJ7rkiOyxC+WQVw0/dNuxkKUonLGbRh4uB1rv464qW2U04YT2ZnTEs
+mpqpwU8IG1+wQZzWz3MovsjWvKs9dNieNCFVYYIeTX08O8R9OJyZ295B6Hmi24P
EbPBYtwfW7ecq+vYpNm+7W7q0q/TVz1X42jURbIiHAX1nyOR+LLNA6HoqriIy1SC
enD7euXLI42EwGRk8uJ7eqh4CUPHRobWJf93EoDvjL+dsMqHyVc+aZktF9GKwiwR
ftPdGYYvowrqp7h8RteZ5ycSxH8WQZNWSJvks1SQ/QehCibVzpyYONStCbYIUljw
416D7QQZpbNxuykK7Mm5ab3GWdFWa1NhIH9/yg2mPF6Kd3V3WvIEy2fVW8AdT+RZ
YNq1xAGjyf3V63RJJVpYe+YtGfnlOunH5+0u+snhO5QAh1T/aefpmMDRgLiYCPLY
YUhiGc8lJ0Z9kj8Npx1WA1tBN6SclvnHSIQWARAlJczCnH6WPwLuQGGtya80xSXL
IQDLJ5R4brxwh7DKMkhHSj21YiJjIH/oBwtJfuyuRR+4a46GyCm60M1V9UkpDqHO
jxHCiyB8LC0gHQDLaWhOb7uoOI/jvEenLOdammCKQtIPnO82amuNWmPzjMbtG2Um
WUVDh8jk4UIIUnsO7KwiRNBGXX9kPgyq0ZiJl6xYlCnEtSmgu9qLdclwp/AkiGXv
2mRurPxByMwWC29YBj5zjGQRKoUJDsQqk+wgYUt5SB6gTIfbEMY8AmxRp2YA5L6h
naEztklisAjosI65WDsNrhTd09b1II/eR/T9nEQfM4Y/wVAUwacnctbCwhqb5oqV
7RSCnGWh38rhBQgaD4pUuOpiZ+c2jiyvBmL/p0n0oBzSPj1PqJ57W43YGPYQ8FYx
L6i+vJ8SQVBUWKhG74i9Nx1OahHPb59/xPsnkJgo8bbPm0X2NEMa0XLodyB0v4Sx
cvIp6C1D373/BVxgqQGCXjgRczyUIjYEUCLFonaF0e0hYbkDSolqCS/Wt3QMFNZV
DhsEfRecLn46ENGYkIerRlFAptHZp/U0XYNtre3+bRl6RpiN+3MhK1mu7RfkdSoN
qYqt7DR6SOXnTbfwVYj+epxwchVBDLRIDCFIPlthBtbDgcl3DuxjbL1j+mFzeN2F
CJMJzBHVuvteRQtkyp8KdjwBZ40ZvbamwcHZcaO3DS7ClwDLov33ReL1FaicSIAA
BmFkN5RBJjsCa9DyrPCgXk+Ve+P4zV3YpLYtc9ET+k1TRC0gjRI9BaQyKIWIWZHl
3/a4bLX8jJPYZ088KGt01oDFS6OQVklHzxO8lU05OAr5RfN7iG895bsBYLcWO+3H
M+ID22gT22hAVHBqMZY7OWZFKFfoZo+ANTA60xog9y6M4SgX6qN1Xn7MAz13YjbJ
fr/s6wK+z2AXDaeMmj/IV22lnwS+Av69vQq7MICZqlq50u7GScnR6QzVyQ2N2a+2
mrz/lToIiwUcDsk2W6LAYMmQyVnN7iXim9vA/vc9TNhOoJIezr+57NcEQ/VpbRWd
GLiZTH15ZZ6iTq3QA1bSYUMJXSuqrIyCYrDQLDzcdtwAOY7X1tFJR9g+Wa8+P908
Bgu1GWthDUz6PLGkZ1tHQwe471S3lsR4s/xAJuqHMbJ+geOprWKjhsd+VfM0DLXA
uf/zmE/0WdqeJL7d2Ki52IV8ZCZbJBkO92d9sQPXsWfqt+0mrPKX38tqKWvg3yRl
/MT5/68GMniBI1vCW0/lw0klIv2I2U6X/In+XkKJsv5Scl+4k1NzEHIKtsYrPx2K
T//jToOsIayltxog7PMNn4NZVc+/4Ryy2/GKvHyLwQ+mLevHUiHMg+9W3Us9PpYR
edR0/wno4Sx8uJucxSq4oSgDSQ0W0BzEN/rOlXu58diAeg15w2i4xozrdVbNBK8/
m8OUCEgPk2r/Ds+0ctLjmqMg4L4/XiDVs5rsnwL7wjzaF9Qp5OuydzHUm35pMfSE
n1ZfMdq7k3JiUPben1KhJ5L1xanO2hfvTFkZYFxn5RuZJ3t/cta4t2MXDkcPXlHa
sFwgCvw0u4Q34rCF2eF+R2O7C54QKck8OwnSijo0RuyDobu+Yko///ZppbJ61UWS
95dO4xr+8J4pHQUi+KldyBgf7keItj/0Vp9dAWr8wA3wJyYQ6JL7W7see0HodXBU
+X2dBhb4kLljQRLrCWvYIMX0O6jrs48E3wvrLqx0WkiVCYEq1DtSLd4t4o3Hut/r
NVvu7gU1Ns1Ljttp6s/qOUMfZZPZH6CSFfRBVD52onLA7arTzUi6P9jQ4hWEOisw
zhJrxbPItRaXMFUUyvcQZQhf3a8/EI1Vd+tcs7jl6KJwYSDq1IjMvAUnj74wSmS9
8ovoPv2fpRZaci6LK89tDit5/Y5BLiHbZLKiLTnfwI4RMRoKNPIdNk9t/9t1oyCK
xW4FMEHGxvTxOxYWWCSCZfws2z2ZtJiTbKkLc0Q2wLHgUR5Ta1SzMTrMMxQbhrek
pUuo13/GLy8ha+EcA17I+JrpwmoUZKv41FrEZg7eEb3VhoTg9otmOos4W2aZvZaW
bDL63O8MFtIVpLaFL4ThCY7t93JN3wrfaxyGZOvgqv9O0CSlPfVaAT2KEOalHBOD
t/WdxmrunEzBBgXFpRU1C882DuP1LmzMFVAZ8Gkycx6JiASvRHt7lqc4CJh8W5Dn
UFOzY3gs9ozgdl050LPaWDCOUw2apF9UxlbNf1z9caigbcz+pcVE4geZhoMa37Wr
WAm1Aa5EDPUnSfb9+ob7037NDAnT9htlkp6aLrlgVoAndMhpTXE/HwShKq2q07iA
6tpbzi7nw2XYOvynH51PtXmgnZuQuR2KgSBA5DRX2KNtlL8T/hYvecsEZ7xaQggY
6c7NQCnEPE+79x4k8SJkZhWyTWWYeiVku6Zx74MlLkdxoAjp0JMSnwKbersVO+P0
bfDWVs4U79NyXrneGDfxdvd9vLYTmlWWV6vsfZ7qSx2/tpcwH4Z1bXo2gwqAGVzc
BJRcRAhAcoYZGHeUJDNQrCPeZhjckpZSMsR9Z1kSQWFeAa0uKshjQlWEO9+xpc4a
1CCWzEMnwSN3Frl9jPHvykvEhRXAQrg2DwW3RuSiUgnIpZhgH01bfHHwwva9sUbM
8lnQmIc0J6uiNqwMrwnSbF4SokWtRNYSeyUjIgpxQVdli8xAXkMP5LhVXAgcANWV
mFb9ZfZDBGrs1tIzx3814aPEnx+MQxn0VNYoWYa5jei2m5iFqT3rPOM3ZS72b9l7
hFcriD+LLkiTKcmmLhNtKQ/HdZ1UqnLMtQWzQYr4LpcQEzgU9OqENK2z9gQzNa6d
jfC7TOz3xEviUjb8oxIsGwOgfC2wR7Ps0XYo+wIxajPzsdN3dxMn0s1hSUHYMZDg
dfnFuiJj1XNkGE5LbO56xH3lTscB2AOr7GE1k1QngssZFhEebEMGh7ruiSef22cR
I1Autz/9rI5qH6Y5kx6y5PCQls5wznmNZPwvrOhzStLyBaJoLSGBhxPWvSg0XST7
IcVGlIZgXif5jtz2Iw8E+ZSrfzTBDUbObk2Jdt4O01LtzpmJBkCQ1Eo7GliWAyN0
DFcGRQmj1EVXqVw1wFMic1yyYNGlKJuI+guze6biXl8eh+RZujbCylbVdDKe+aR8
xrNgbXIh9Xvf8TiAbUZ7uj2dQEfWmJM5liNk8ifjPFMMYbpD6z/Fe5fxIY1jDFV2
aK5PxwJVqCT3mWc8UmBw6YRiPTq/ucWqlZlXbyfTZb/ze6zrItnH01p7NXTDuTvf
S3bWamqhUJouw1OCcjxtwYMwJtOP6nHcTigEf2TQVxkKawPSYWytY5P8ZG42j5W+
rgiG2eNzvLzQa5M6c1uC/lxYV6kj2HCZeaNQ+MZyyP7oJb87oIA4n3zvkX+HJj/X
6BDUjKFWtSmkTWPAvM9gNufPNQeLd3j8+scQ87DuMLsfNfXiJ8/ScajiBsfMrO8u
mgzmEoDcM2QbMEI0dgijWSNdV/0aFDqd9pFoSMCJxZfdoZMwAHac+Bso52z/zYrT
wkNus0FvI6ySh8XbSpD2p3eIh9Gg7mLS54QXD1a5Pt+nrZAPx+caEcF9DrOpYdpF
vdsd+sHXLYmSFT93VrT9Ob6DTDWnPrEMnXEGeOzkJa9Jgh3yIpcpxjG/Fevq5qi1
QhurKA3r0R/2cTDSQIb31oFUe+G58djFXqnv2J5u7GKh8Zho4EHdsUimuBna+v9P
mky+rXSP0rhXZvzbDzu6JKXOE2tmSPzBZjasejV2K7PgjZ0nM8TVUBfY47WZeL7n
//F3ZyBVOid2yaIjDG4Dqfq9Wb5qkXdzjcENolJJK9NrdIv3HuPVlPG2ZjF0vMHj
wG0V7GbKhm3KkR6jW4Wv0oEE63UARjBgVvCvD+FHlcPpdJ3GCKej1eJAs5m8DHs4
xDrXZAVXbG3WJ3kAQNTp6v8WElx2eZkhpOB4TbGMnMHDn1lgbL+S8kgVdfXqifWa
+j1VbMlbkuE2Edf7q2mlS9JIxgaPNnaGjrkXHDMwwLM4bsKbQdc3vvSYumhzvMmN
E8JLd9BEH48syMCijnDTfaiQ9+9Jk+cR0FNj5JVqQpX/kcurbn7cUqFgViDhG1tx
`protect END_PROTECTED
