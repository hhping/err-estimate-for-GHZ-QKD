`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQJLIKp2Yj0MXQYdMOGhAMgfjbTVAN0Wv3MXaElMgWo6jSVX708ALVoHVX3zlJ2E
y+3ohQpW+zeSSgNK9v/unH5Yx/OWM6QkRXnzfKA0OfIEjIxLNqWEEDKOOe+QQNWj
IiGlS3zMSbcSb/a6K90WOIOy8BWOSjiL9EZRsZT8jbR7wAn6RfgEkKHzMiEQifCP
flIFgMDAMW+NdazF+OP6nUH9ah/M27P9EpBABcmrC4qtiTa4Fo70joFEylL2P9o0
J1s36rmu5n8uV/nlXPC9eA4Q2SEAHGbPwFs3rJ6UmAGfPhC8NJaSZat8JWqhQVpE
3km0E4QoWGifxlDELtrYViTRpAWbR6YbNM1lhJtbbliuNPk2aLtSr0EV58BJPq2H
JWKmoP6z0+uuwZ1/TsI/Oz4RhGKYWIe/cQ8HCBN2G2HL6nouHTaodMIM906tG9NT
6QOuP+EZG6MAhqJNKdo1zCzT9TXll0OZdGrymLWRkw58sizBE2cNUE9Y9tgeJWx3
o3nrgAR0IsXT7d2p5PMXxe8l2aqR8V+OnwEbOxEyLZXO72hwphfrVvrGp21X1IpU
pbt9K5agQeS8jAGfegIoJ+ipNgAjS5mx0j6YZybgqfcwv5545sHl0U5UNvjy+4SI
2sTDYYPv+doYUkPnf6I56BAd+XusY4H7VZp4hlgngQ8T2dBSfYmDwD+b7+QfKt3b
IcYMqyermhTyajjufqP1ZmP2f5BrXzZoO6i+y3/J6b/AYcsSZfz2eHMKgvoc7JdT
XoHnKx74DXs4DYEBkgr//2T+U8R2Pr58Dyfm5pDIFGqc+EG69epA5jQZ46kazn/h
XOz7/HArHt3lXijBn0mmXqdFO2+utwoMaVp5emiVWNsKK73bykGIrWPr6jk/wIhP
K14qsaEJOcDhy5Jv7/MJhAmEw4kmXUWo2Za/+wP/T7WmBNLJ8XWs8qQmiZIhzHKZ
jfT/1u3/Ffr4iSGVkhoEU51fJWq7FJ1+gRiQP/W84BcOS4fSge6HGbxPtzWBYOEO
sIikJJWPNHC9Hq9pm/OQulKxuXbQfslvLMVLHyv4wP9PHO+HQkS70W1bu/RLx+Gz
JLZYSWagqs2fBFPr3CA2q3x0uA8Ghd0SomfudNn0BHVgsuaaup9zhtlDScM6il/c
UYkKhcc2ySlKeI1xtLk3M7bTQtTVNbkzQ2US3z9lspvYjOrUAW82sLXuuckWUvyu
Cf4uCKqPlfW9U7ALBGye+Q==
`protect END_PROTECTED
