`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5xppBVt7cO5P1avf8vcsfEz3c4TpEouUaLe6+GFjdLlYhfobQtoW95V2zLFJHY3
AtWJIv1YWqDAjQBBUf5zMzIztNzIVeWc3t3aCmUOh+Jdj6Y4U1mIexQldsO8Hxvj
uK5XsRHxSLg1OHH++UnCVb5MdEw9X15KUlAwwUvTs0Y2AYYpyLkH7GqE55NCpmmI
SvoAJCt4MR+RHD2zfOkHQ9foKGECHsPrL1G2MMWUd/r6Q4xnH3ICteoUOmUrsfmo
qqGCd1PyyNaIgSBWPJFR+72TFVgeoMTm6EaU1VJwIjQsPCwNOwq+1r9xBcfYXyj6
lyRbCLKLFwKAJr04eYqvD/lUzJdSQ8dTu0yIIALAqOge2gVbx/HOcIImYE7wk5yq
iM8wMc+Gmpb3h7dJm4tqjln90PemBnWbpwbqsmv15a4gX2KbwYdvLLDrrECjpb/u
yBIsx8iUHsTlbZOnETE/VPiPMwvEh+39jUhTnFnf9dqkRGLQacwweiNZjZJ2gLLv
NewjW8/6VR4SoQMZ7utr24c1Psu5NnO6+l33l6W2qhhpClkZD5A2ybE9AI9MPd4l
+iC5iha25oa2Q/d2pkok94c9L3ydELazb9MRrcpm4U8Ph0VDiZdataUtA3erV/sO
5ADZTnBdxAnFV4ArKiZcWTXswZSIIoT6N+P73gsY6bKdxCpIMMl7mjInqh5vGyzo
1CI82QWsEQpXMbMQauTSu9djMG9NqJxG0v2LUGouy0QvMSF1RH+gLD0XV6kQ2BSh
bNUhbEyP2fyXPkaZHKwsLlOPIqLW2rH40D3/Gy279PN78l3Yek2SKTYy3C+FxU8A
Zky3e2zLa3v3HbfzSGfl8HiIavqX3Jf3ZenOd7qnHCnvMgZ0wpp5VhYd0OXxYfOQ
rv+MDRX3HAwu6qg3gts8NHzHLJ0D00IASF0QF/KJf7RelqTfZlFTywuAnkZp/M7C
c1AlkCyS7xHNVm6sbtVVf6gGH7KxhLOFNXSvytofMVmiTKfoiiWzDoWiiUyNb81k
ytTJE/um9q1yPCmY6k70RjCHsA5XTTHhhMsGXbitfwDbjYNPW9EAsreQKvGZgU0l
FoKDRX+p6Y1YqonMtTb48dstsnGL4m0jNckg3nXAPMvziOKUyQzjhguaqYdCvp4b
MOCfbMqxfiy2lVVNqbQq9Ca0Fz9GQpCge50+LncBwruFk6fW0AGOjBeQl+VdEfrG
klWYR0EXdSpZaSUc85GbDYoB1gUGiraIf+W8nRGnyNA=
`protect END_PROTECTED
