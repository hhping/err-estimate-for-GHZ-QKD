`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0NOfwuQtM7/EHjeqqjqG0idxq5Ym8oYiQVWxR5XK8WZEcOgOzqg5g6jjy+7p3BrB
xYF5acglKV9uKuFPf7SutaNbwVXRvo/Ap8RBPdLkENgWz0S+Qbisi1rHEiar8r3s
GsxjRYL+lmEGBr2ExnSJc+Re57J4XACN55uvupJkIBNHS4TgScjz4u15+fGNdGbw
qTJMuC9jpTPnQLRH/biCunK3rIyWHzcc2g/lYywMisNP/XjT9p0rUyQwkfu1OkCc
z24VxPLDwFrMlnFEzVBI00TDnHoJFukvOj2BNSpVu7StWzy6HCt58Ntiep2yeIBL
Gv46lH8g4sHSZtuh8RIPfy713jdvEr4E6zX5hXbZOQTY2VA70vDpIk4JauFw+kym
`protect END_PROTECTED
