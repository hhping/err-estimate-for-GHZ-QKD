`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k/cE7AvEnPWL1b9Ez1Io6HxFlH2MhY1E9x51HkubEZLPaXWvIaoRSW/PIMquHq86
xs+I4JOGlcLt0dEulrZa2Bd/GczKQPwPa5+r5MpeHLLzkqgypb9TXp4KOt+Pcln3
k5VI5cq+6hAdGsnkG+P5Q9/7LZQIv8Itqq/uoUQ//LjpRc+VSqBwAQq7BtVrMVM+
hmKvL/qCMYXWq3GxvE+EHtQ9HiP0jVi2dZkbTCzc6ka5FDZ9y1xVKdQ8dgrZas1t
hKqNmxxm2iihpzdFvU5rJnYclhsyQm8N+7t0uD9fK8gYhIQJ0tarHl561+4YtNSm
s2W8iQN+UBe8GPB83cpA70j8KGzemiIJuhh5tFYpCM0U8oThqHzV523EJJ8ROb+l
8t+28w0m5SMUhDiqmpValbZt5BlRzF+aaXHqBOuG41vqK3g7rrqsIKpdwB7c4vGN
EemudWxTd0vhxT6tyHy0HAJaPLfI1iYV+KhKmh3PzHZ8OsdLtAakxHK31C/O9llU
Zy2Ma4XZX8slTbHWZ/uKCdCplX6MVapfPK8oH1N8cX1Bb2HnhViDWPArqBwxns2V
qnMJJRNPRWyaMBvcvKbjBEtBQ5gtDZn+2MgMzvJbWI12Xj5XrPMwVteCz56cBBHf
OCJAWKW+uO+r3PJKefXu5cm6F3DwJOwFYIh7tV2hjK1UcQfoYjSBnyC1DXDsJyK3
Jg35mMZuwk6VhHOg6US2ow==
`protect END_PROTECTED
