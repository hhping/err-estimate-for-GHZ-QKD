`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcajKEEgibDQiwkq71XL4osou75rYH3XjXgNolX1X8/K5ZhntjgZHoxAlocgCIl0
Xd0DilX4yEFSD1G4ederwTM5u7+qAibiJlaq8eT70saoOHSjbIr0ex6tm8VIX9oT
BvtwMehikmQrFYUkz4VHeIehdl+uuprDIq9r87d2naQrwNi0Fpczrhl0QLj9Y88n
wS9EOcbS0tVRhGThCl21LlMgrIz9L2OdvDIPpP+7rb+1/CweGgvlAvE3LGP3jRzZ
awVVAIHmBdak40ZRu9O2QvjiHTXoaDSOmU+hUxAoYqPXKOtVTRZ8sY/iMkmqyJpj
vr3Rx1rz3XeTuYIP7FIb772qV0RDhq5OhnZKhHrQ0VpiinubmF6ZFdwkkqv1kQ1A
b9N/ItAMAv6x/Qd/MqVKCK8Aqt3AJ5GhkBW/ygP5mur987VqL9Vx7jgg1QyzoVqj
NaVSBvcYiye3agzXyc0PkX601lXsr7gQhKQYggTGFjyYlE4Xv5NIPqJpD1waaums
k3futDQuco3jE2HS25jbKnlbDxGxIN8YSz6PSfO3vmXzRrBge9i8UOeVGMzkeA4p
v55voZ5P+3MJ65dre4gleXN/dRTGPz9Fo7pj+YPr45H2LkGBI4fXKP+QQqLboBgj
28OoIYCCpFH81LA57w52enGmWk1PoHBIgGCRhAtXWZpCvdoFnow5VYDIAIdF7cc8
Y3cj1FfTcZYjTR6gLCtz22LHUMXtV+ZwlXLbRMeSFqjcx+iQY7LshJIWrQJPYNMp
YF0qykNkx2hA2fx4bXmsVQo/y8xQcwKnSS/gJseoueeh76YP6e17+D/K2I4uoCba
h9BjVzRqL8n1b00/utsSRSPF/7q2eQV/CpUUo2TovH/76FYxEitoYO8Uiu94Rtxh
RPg6yBPtXAPnqYSb9TD8ADgvwjDe3rmR93jF5mWf9M+lVbeLDecA2tWdw5qNfQQb
S6o94G0uN8veSH+U0UzycoKyL6r2NE/QvMAUgtFGrgIyqw8Tsh7Pv4Al0gTWW/ZB
OtIDDOM3tPkSJxqyDmUsgW/TlCVonKMA/rX/enQXdcGQZtpUL8gLTRJd9sbYhnsW
e0V0lA2OmteznGRIFNlsibK/eAMA594uBkuiFTxDRRrq76V0RYM/WYj/77hJXy+5
t8rRXjS4Rhuwovs2kOndzFIRuyAyU49o/unC63/fMcwH5kB8mjq3iitegJLRCCKs
yXcbQ++3N6tAB66IW4qM+C8QnM/C+YP4aK9oSfwk5NRkL/GzEo7cJsFtl0cx0Dju
MV59RMunHEYquJf+v0S/aO6dBSuSq4+YOPDW8rxtGio4DEXJbyYo7Rc++oDMZmJa
rusH+N+32HanwbOLb2fN4cWi1/TsC+1GvH8xdFCMTnsVAzetODbbX6rFWiMY2Lar
uWhzLwi4Ypu2fIQzmcKzBNK01JJsT6s/7vs9qwPsCWzbzqbBFuadzks0zFTJhX3I
YatgGKYH0HJb45E71r3vhYOIZfpW+u6u8IbBKN69XSE802zBIF9gNBY6xYUqZhC9
+fnaet2SQwBHzyhRm3ZFI209CJOltFH6Bp2iDAU+csWQhFbZQa0r1qp2yL9vXigZ
NWrDnywIAOxrwHJ5AqG1ir99hNO7yWloamg/NWAgmj6qYE8e40sZQwFpIYNdOktp
WXINCqoBhpKR97Q99lWSmbBO9P4nVuuUQDYbMtWgq276dbYUl8MIkZqj8PoFM0LL
+GOYgJ1gT9nYPTd9HWjLgvUSH4zenK/UySCJ7Hd03meVh4GcBjHjEU6j1RBO+kj/
ygBVVXGAhgv+yMED0kB33f0AfQ/IZiJ68TjS90YoIhFNZVGHD0+jnrX6Ct5uc2LU
L6Qs96ZnS0gh776WImpbtEh1zO8J4SIduhnX3uENgfPYeDaXXgJbayQpElGTMTib
OMnPbUlIamsSm0HsInYz/Iu+SMPMsWsXsuI8CIE23eZwQXU0Up+ZOl5psG0PUqgO
aw3NV89/zqZ4dCo3tKE9lnn6sozux6ua1gMVgjj0AzDIzwLlEYGvmt2Tphdzg1+0
FUSMJRyXi0/xWS85PsV2x8JqasvH9+Wl+GWw9agsyy36uOvjI0+Dfcj65RknxZpg
KZZKYh9Xa9M+GCCdI5ptyt6RhMZ9xSswZ93voyPKfgLESXADdUYGwPTjwNyB6yfr
1yo6XoJWlL8jSK1RmC/dYm5F53EvNHLcZd8asq32TsrD5Cwcco5gCpm1O7YFQ33m
B0wvoccfnnKc0emSn4td2sFw3ssCQDW11J9mJ2O8Y6urMd98ZNQH2u5O2szSm8+F
fX9XUbPNvdydAMFoz9io92hjgLZPcS1bDPZzimu12K3/+2+SYMPCRBzxVhDywd7C
dLTs9lXFb9YGOBi58YlZsff7WW/YRtckQbjx9YuBSrkZyILKGFXRUaNGz5Lu4gaZ
KAmSOMeFxAuslxYm80tG7j29HEd3CY8ZGO0j9lcxGK15KSBGjxjTuARz8KDP7TaF
pgRfna694pzNDjo2mxKbO2/0lYgkKy/9tR5k1Cmnq8apVrvGdmVQfBhqFtYwpaaK
gQpAQ4CuUCvr9djRBiXxxzHxWTNTpilrHX+bY02+43M4OJqyHNG0Owb2h7vQiHNc
kkxa4eSBQOH1H++gQp71R9R7BbtLmhtFgCklSM5V+p1H7gEwL+irwfQZJym/p1gl
MZyC+mcV1atmDtHv75Aa0wzJD3nze8uiGamOP40UOl40kHfo8Tf673F+gqATa/Qi
9JCTieV3L8BZPBSrxNqMmfPs0DSaDXi9rFeWCgvwcGXR8hbQZvwakt+dS8i8rvjF
VUc/5kf3B4uPcUKd+IYBsfrN58UVn3aYQltq/kkGXjzvUxE6F4T2waQu41koVoYQ
q6k2EnGQF/MZzeB+90epcoxBM8KqdCd5sV9djGRJL/W0W5e+aTpTfShwRHW0x625
0fc3twydxsDikoTFJ/VhhWncbzp7OpWw03ldWBCrl0VMy2mG9EA/fbaz3SlfxxAP
`protect END_PROTECTED
