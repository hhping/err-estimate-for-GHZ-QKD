`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qZ0JO2f4J5rqCgJJu+JpJpNiSWDhBMLe2m0AvvJWSX0j10Ps8h/GlgcWnawbosZ
820mdsV34I2WXBoKbhyczfWZ1FzPtPnExWmKQlTAA+KbHuIWG8tW7UNpioTdcjoy
etOUlwBbhEi2eHuu3xfG8VIme4HngBdpiv18fyjxTj+s2Sl6UPF2f10rTIxmkdzX
9aAdpDKsapUE/KfkfNO5yXn6lzS8K3DbEGGvrE5RaCoMgnqmiZHiOZIc2eZ2W+2V
Mr5Xu3xzQp/yJ76R47Q/YoA/A1ehdSXXc1ZB5euU81UGfLxECurFDxvOplHkLfo/
ozcHegmHOLLqjT56iOYzipFkzGuC5B4OuHlVyhuMF4mkd7yIp1FmexxPUsSzt8IP
bHz3dDnyjgb2Bw79T69p8gQCqH/UgDWNjTVtDiplqgg0QUa6cEJMgasuEyLt1BPO
pdq2z0QZLIgyMbNF0J5aU2ILoiv/IIKuDPS9h3FHlWiBbRr3Kcr29+Q7nruSM3lc
aW9nQtwnV+sMaa94uSOu3Y2wThZN4uZrLpYHWc7LL7RJWbUjiUBIN4XD87BNnKBq
50OFGElewGgp30lQCH1Vg2hHoZ2iZ0nto6UqQzg8oTA=
`protect END_PROTECTED
