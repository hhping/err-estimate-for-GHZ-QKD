`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6iAYJWWMJjKLhLMCie4st+3E4KiYKDEvYr03GmVpFNIU3FIf22A8I+pe7Nl8dzF
0wP7cshomHN+7XYxVqf1ZpNwWJtM3GDx0YZ8+H3vZGAcKHO4CLK5iEuyyL5I4X6A
pPHOuY8cwtm6OKHAcnK9+cco4RUoEvKo6Pcr/UqjGXb7iA4b3ioTp9YbDLdSvTVj
BXStQFRgBk1fRoeE2XgI62ooN7bh7uDsXw855W1jRVRyrg/C63QcEJBcAg1qiej/
cglbtaMG/D1zOQ2eRUrjGdKLStyBkYVQm15JcAslOpFKbeYqR8Jhu6FHeeMiiihH
fYHsT+eS7dpX5/Iy+09rpsG7x6CMdSYUUV/F54/UX17VYjQdf8TAHR4Y4x+1IuvI
mK+ob7+qVEnDm7hM7CFuqa+VRo9fVoXY0xmvnPSIseRvxuXcYbwFxyuI9vF/9Kop
QnBfzznndc7gJlMh3W9Lvw==
`protect END_PROTECTED
