`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15e7209lHbtKVvFnA+JUG10ewXgOM2E8AF45ENESD7JTeOA97gqGCxG1l666r28Y
bzKZkgafQ9PsxXjYi0yxUNiF8ob12TGLvgu45oh6m0hALQ0cgFI3bCFMdcqTKqQm
o33Vm37Lrx3J2ja1yCnrklJSYlsQx+cTfmKPX4fS3m94xy0SWUy/Eu3NHevko2/j
x/wz2RADxqxDQJJXcj+TQ5oY4OHq0X3YPYD+3oZoaAOD0N306Ri+9HkRSF+jnPOM
i+g4zhtzvl84kEaNfWsqmCJl2c4nVn4poGYAyEcWYKMQvMDYoJhT+qgucbcW1j8w
OctLF0l4M4QnVWuwF+j4/Kczi6zQISYDSjrkHcn1yO+OzvK+pvj6m0YmQSRyMUNr
TqxBYfCqVRI/+f0AkeqXcYotkDapZ0fthlV16L4qL5azALncxJ1GslN6QjlSMiDJ
1fsdvm9C9uCPcaz4LV5DFQUDDoM6O5mDxYITXnkj7nIerxx4JZb6kqUB04fwNFCR
OyoeRqIVC35rj11yEZ69mWbqX9CIPjdtMurfAjEnNtdNg5vhPxcAr1UU7LG8bkQp
Xu0NAeDL30EhkXrU+Gqu0Eh0nW62yY79fGJ+/TLruKfK6Ix9yHWdpF8HQ9cbTW/a
alckqLnpUh2Y9Z6CfECbhdY6UL4BIpey/YmpKb8rDmxWTQqcnP8e0GgB7mA/g/zq
loNoEN+YD11SKKYr4YuNwYslU1T7YKVavnl2cC7/EIxESCUNKwbxVmoEScEDzeX4
7G2LdvWQLBFsr4hI/coLPFCT5pvl7wZOzWKcrW8NC6WvaWW2cAlWdQ3oJREzK9zU
20KIrXVRtKOIYduZRrWYSOr/hWmDQNBE8SGaj6+Z54NCoMPRERsFMyPLM8nq06XH
YnuhzrNMpmygX/sFTL2oaJD1rjWVPwiAMcJzaBuOCl6jP2CP+x8sAVGad+AioAw6
JTYIxubqAT/woUpvAvT1NnHbQ88IvuuEk3slh7Bv0DD7YzUaasiaksum+RWvxciw
zJxj3b2bAq6RyQOTACfvU5oDQd9FGpKeE1ENvX+kHkE6IKpToeO7tXzD//fDQSSd
PPwTCuPtnApl0WYiv45tjMeeLMg1BB0dzQ4EAmAWfK4508guGimGZs85y8oGwx/6
PKUesUP2Ko9ojoQOE0xIlxY0hVm4yj+hB9VrBnBkduiYjAVaZGZJJXfvtgGrqSja
ynbxTvJSZ0TerbW0pZwlgmN9eoLnr5cOaWhb8JzprA395Z1XpQVI/+PzLwKn9yf/
d+JpPPn1Cwz6Xt7vSFsjguaxx/KhpGp5Hl6E6x30ve4w3xqYtQQpqFL4Ozun4+hB
ds5pKOgbtgjUgfJMBHMMslItSamHTe/G/wuErX9YXX7Atw1P91BR6LBk4LPOvNdz
qy2JweKN8lZxG8pzf9quxN0ScqezFLn4fQ/TVPGFap6OxnROo/whCWIv1dDBmY/N
+vW6cpOhqYTsqJY5SS1yjTqYgdmXyuxklw3CmLe8Qqi+DMJsQ4fsM/ZuBe/gHl1h
MTVDfE2/0jOtnL8c8UKVdSZnz8Tdaf1z9MKUE/cMreZf/7RK0gCECB7BKHJ2XWgQ
tvZsIV1825vpgr8M+5Z1SO3EkGUfcDgCQEB0RBuVjnctdRKfnSVGapV7Ro6XkfaI
pHGkujzzF0NsU+ND3YXhKLAGQCrC53BV3Taj+MX1Tcj+wsxgyc2X2b7N5V63oC+o
xFCVyQ2VUItsC9vdEPSmu9d9rFj8RFwbKIMCFjCWA6/4W4EU6gY5CgTUFnVulObs
nV4byg/crLPmqG79tvD9Rz5Y0psMvqe3ws/gQoPRakHXCc1vM1Wd59L7HaQ0JIkH
8eiTe6xe9wtSHUBZbF8dBqUoaNYKutzc4vQ9SXR52Qhr3mcTlN49ewztoqwTzeWW
ewItdJbNhShCzWzcPo8GoxNsi3PBG61x9FM6eoEP8GBz7dvxHRMDRj6TdOwRmPdl
epoO2HZLIF4M30WY35KXMqvt2b8FmcOb5Za1qMBI5kDZUNDDt4IkoQF55+ENq1X9
0GuAL/G/LLOLWTZ2JOEMb8ew5YTEgpWmTHEf+KWRUGO5VYH3LajLahpbSvJ7pD96
Q8hE+mzrZAm3puxYqzF0P0KVJe90gvIWB0WCpj1YrLp+tmKRY10oh5+bkfVOurV8
m+6Y27Qvg396fuh8WRTSBKW2Pe07FmmUzA/LFna4FXzRgQiUlnELgzU5rm9eyTpk
FQuHJL1T8NlSEB9BV6sAdTQuGj2acRa9gs18Z49b47S3WQSNwy9DGJ3MV+IBGPM2
3jx3dNC+cMCSRCNvoMA+p5RgZ2oAJT78KYAQwie3uyUaLvNtLAU8v4IJz2QD+XOD
l4VKRK4dWBm9B1F9ovZpPqC9jTavH/q4xgux1YRBhuQB2Fg/061+QIF2C8iiaofM
cUH5thNYMIY6XdKMziTV2JbuefOV92OgBTzH9eyqO+NtVe/dfXrUEiCz/A7a9X+Y
Tpl77qp/lY9trEg9L+VI2qshuZrix8vvqAXNJqrXe5r7TV1XCAn3cXlT2MyWEzst
JBhV3iOtVQvfNtaD9Gf/klweIpdlwXskWRvRdbSA6/O10aRd7WBrSb+dlC/2RFNg
Ti7l/cw2PJ3lIxx9yswlPx8oQEYfHQ1MxZ/BPPUu7kAj82RkM4RSP2+sWO4NbHMl
Y0XXbCuWy/4puCkHsC82Qtpm/2mnH/5P1yGo/O3gmHx3X695DRON+asjuBefYMy2
euI6Of/LBl9HOH8yOYuTacACmabKK/HbEjHS68oj+dLqhCZc2VK3ds8dImbn6Kmd
BuFwbNPRG3wtcjVYL7+YRkHLS82G/1wv4mcyxwg2XfEvabKxTe1Izn94Gh2WPgrJ
7yHjYoc5AyjbHtGtDmjp3lfbwhOSqPUTL8q6DDFCbsWVU4uWrSLc2d92ste842Ee
Dgm4bK2z7Sw/iylg0r/kDZDIY/2z4B1HD/31AufHE+IrIdmapUsrpvTG3q47enzu
eAnXmlBfb/LarAg7keHr2JhBExMHNK/fJk11yiGKjAqKzA/NUFrmy/pueTeK6zrW
FpGYqCoia3KVc0qkQb89ihcvPH45iMlvM+vlVwTOEv60k3C5Sm29IU4MLEFsypE/
Do8i4p11S4wUfoAyfT5wuGakXfxf+q8iiIQ/MHY6f1l7m8ktvnF/mbmyWgwbb3je
1V/RT3J/5h4W8bZY5VrNmIFc8wV0W+GqTVw+5M5RxE/MpV6x24AN3NyN7l1leUPv
1cq9ODGnkkeQlkEPHgF3ktmu7V+2EA4QYvnQcZrOA+I=
`protect END_PROTECTED
