`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZsjNC+g5gydep3GPXaFNXNSkO0SzM5agKyIvCUh7C1wfCfLiiLzV1PclNr46r1tE
7JGpzkuFISIkHZtK8edUF1IWVJl2MMa+8qFWDpknPOBwKQDpXzJ5r5P5o44dUHM+
HgQgW6dHB/5Txd8eJJizPNSOssxACZc78RHd1Hnj1fFUdAelxDfR3TSe+HY4a/u+
/kGibSfxtPtNqjQExZNEmJBlD2PF3SPlwAPuA362cWNKK1enkAKEsHoMdeEM4uos
SxSlgtEpzV66yoSWnG/7bFDq5v9OJAs4V/aPs+wCbBssVW6tbjMY4PSRlewszgRv
Frj1xEGIPLbz+FHQJ7rnkaHkAaAVnOpBKsE4CG6VyyGdb1TNuBufGTT2vDq51TOg
72rVL5k+PajH3XFqpWWKjqECCsnbVtS2P4D8h/l6feBmhZWAtZAAIT5x/2PApa25
McNgFsQRuZi1Gbzi74Y9WZNAhON8V3Uo6LSUlsl8Z+zOIi949hwfuWojWRR/Iiw4
RUzk7NVoz27aTzscIZYoQr5qy6Vr1ifFFIappXub/YV0+MBLvRCxxyQkI20OnMrV
nWKNMblc86xMt3qpqOwteGsu/uclABJ7bK55YFbZduL1Z6ntgkL3cXVTiz7ugT3Z
Iq+tlZQQtBiBY9WCYG94Ea1GbM7nmfAh0bsX0BfDvS5TDkHQ3rAdho65fW3VeEV8
4oamzXcadYtJRfD7nybfWcYnyTGFljQZNJzPo+wHU1EINcov86iXtfjfSxSRQ/p6
3NcEozVvvMwmIoijWySE7YSCZ5ECt+y0pXysPSl3NVIGhcGKasGGjLqZ8EfD5wbj
pnG9j/7OXlytjsir6UqbHZZV5gMvcZCs5j/E0Sck7uURplXmGWvPk5nChrkZwzww
skrHX8f3kXNkIE4/ZqP80/rrKGIjrSMuTCFeOUBV0c/GNWSAaly/ydi+B+Hu2mAj
UMZ+cU2WlGP2YNmJHSo6Dxo30UBb1oI8mrloPtnyBgErDgDCLZHYVayImB6hx4Mj
o9sJ9RpM6C8Qnevp5/ptqA+YNwBPWtSTQPzMEqIBTcg=
`protect END_PROTECTED
