`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/o23yIvG0v9kjpCa0uoll8UBu134jJvt+wWy62OaH72rVwbac+bd85+/J62xn/j
Mw7UFb0UYKVWxPB3/FK8E6QSNZQD4gmRRtrOC8u75aM22qNJpWGjgVp7OGT6rbRI
mtqQEKNJ7GlUaRZYPG1wYeSimSJUxp+WkZvodjEgv0UNbzZx9VGtX2r3mUSfR8UY
Q5Sm7ZnXhuWVPtbjYSF+K9T0VgCO2GfqElPk61nogGLV480bTwRqJg+lxS6y1dFh
XgV8d43rv7JEVFXZr6HhQueqsXLrk1hBlV+KgRdPLf9+l+W4oI8StinaspwM+pjS
D2xn/6DRaAQYMUmhYuqywakjloMxiu+Kab05xyR6O7xruO4THDIiQ8qyhRy0SiJf
2F9VtGZ+TYCJOV40o6rYp+dHzdG/oFpCHtW4vebHIjXLwRSNvKfhkuh8h+K1PqLp
xY33xokAD9zq8jjBkjnYsRkNsh7PYdVqpmwANyXC30ED9+ReWLAVfQLVmMT6QbZk
aw5RDLk3wInUhnkoGOBidjG16p9eCg4+NC/MuwX2Tkb3E0erS4Iknf1cGeORDHT/
aCKvrl1BOZV0FZ+pc21L1PwhIDutNizmyQTiJ8jRF+MnSMo955YEbBEhpLi3qsbU
XFPEvv1lfQgR9WC2ReGqU5hTqhz9DQckal5lOMvbf6bh1h/+igBfAXC3iDv3D/Ft
yoa6M1UJ/0kAN0RJqMBcjv8yi4rr32mUAvRkOsl7BsHbgId4mmhrvj2sbLZm++kP
j6Yy8EHNH/ETOlp+G1dlt07C8ehGSCqdXyYElz9lp/iFEN5pzOcJ7KemcveQGqAZ
MptwGal7zfowpz0GsSnzGGuH2Dl96LP9VZjMKhnRT7chOZItZGRTrAt5xRgCwlIa
JIzs/AoYXBCH1so7L4pbjkdL7tpLLzQ8NRnC+o5UeadZAOAU7hJ8FDi+SWiU5356
rgjMUv9/+B5WhPeuTsjLhMOd1E0ixpUb+BgRtaE8mVwnrl1maqe/wI9FSm9mAQmf
zx7h5gQRXCxUEVSFe+Ug33MkXgkUs885OmX0yidxqDM6chsSe73qw0Y7f+/WDdGC
hkrY70WEbEaRrTjuGX8315pcsCafcsxOOI4V592UrQkplobqgbQPdeL94XuisP/p
LwjU0WYCYupPOQ5t2f7B6VnyykwneJHLn/OQVuKfn4v23bhRWHh/I1ejAazcZDaD
k3RxBTyGzL7bZLBLPRdjbJlVtX2C4DzZmCouUOzyj/uTKlhtglr4Ij3OLHNWntvs
5eBBOwwFhK+M95NfZEl22tke0/FJ01q6+IsMyN2au69TAGYVv9LTBgXPGJdS3H08
ky34uCQm5qWa/t2noH0lESNsH8l5YB73iGCB8ZV+woQdk351tA6dSel9O/cj6o1h
GQwQQnPlhCIvBK1uqFiCRuYkLwDqOcGWdT7wAEZWEhrJiOXRSTmW2vmLINrQ3rMD
doHDDwWFwfcY/Hxgc9PmWVGg5YUgUzY6DqSPWFPA8h/aADlamFjtXKeFPIFhXRmT
nZh23nCFWl+T6LeoVtnZhWaYwGhOEFBiKMoSeHqOrnz3Y3Rt0wVKGOZzwso+r5yd
hLdI/wGfgS9e+U3feScd+eDX2juZqPBDvBxlW8k9eEeP/BMTB/RKQjM0o/17ULAH
W2QstC9sNYUOnDNWtzq12EhEhALA9mVB3b0xe10VMy23+REZGpu3KzRJhbBQmZ3s
/4+iGkm3iLghyduyc4O3nW8oLvesTzcwnVG6WldHQCyCuAuzwbOO8sOxGFq8GXXO
xM7YsXEF3aAij8e1i1viteJwR6duEG8w5FqgsudG6k5Lgu28YHZtLteRf83K4Ylj
zy02FLgF5zu9FutRZlBIaTz6Xmry5mBSEBz/cTxgLLpIMZuWKBLv0H/lKzl3RghG
L3qA1u3Cu7L0F1wZp3dyvLtDOs7tcjmxhOiHtmRgnMPNWSumw+8MTDcqfJx/l2D+
7OHlJmSZTpBSa3E/1NWLXf557p3M+BCqWfFetoChrGWD880XV696Ql2dCkflnbOo
olDjryImoFuStkMCR39q3TDNQipBWM6IdJUOF+qlxrx0PQ0bapMFS0vXMONdgHcd
sMwN+yaUXRCSKAKeUUNsl9pJZ1a6IswO2+jFrOp9Xyq+X5wohBcpehmbZDEPn1fy
SNFLdOhbdq9PyYz2QoRAVyAB8/TdnGh7sy1onXzfIaY7wEiQUb9SkcNCau6Y1r0L
+awzSLvs81MNk+01g05VA1L15L5jhNB1ZlCT5o1M1LuFiOegDoQbH1ZzdPuLSTPD
ENfjvasG90DyTE1Y6UacjlP8XnpR7n8lYbh/4NyAcGet7OJLImYcy/ATbru2q6Kc
v7v45B8/RH0B4/VOWANq+WpfIWogP2JGYY+wo4oEGWvt2/y2lH39/4H1OC2faxkO
hO+pTSmY1fMKDC4sutmdadI3YYvqdq/HJMqLUrCgCXBOjVNFT4VE5b6MJrBCRKzI
Xha7Qy0l6oOAyYmsrr6lW0C5XMpBodBlJNyDftbcQyoQDafH+Ibbrfp0xoDFIp24
ssHYZhLQG1PRvm3Ihm2D4d2+bslrSVpg9IayI9ee4pOVgE9koNgudQJnl7TRN2J4
sTkAYLDWsx/G8/FnUlrUx+WwxDmZRIhwcHPY+EiSw20yYVEjrr1wSwseB/5NDJtA
YzHe/AQ98dkzvcWvVidvGEPMD/cupIYsbzIGJnaJBcIMd6+V9/QWOBZ6Uvu8nf10
Zr5XdKaW75ykZD/LAtbsbeXTtopwJ2/MoiR+j7gYQbTWGzHCjkdSIFI6kjLnLdoc
GHIkbrzjstbv9nqEFRP+IThzj+Lq2FNJHsvkfSWszjCKjE4ghGP10ESpOt9BCADl
LZOPhtIBiLZWwaRnHgR34R0yHAH8ZnilsWu3NEp9T/sBmzys31YCNUJQKpcXxyl/
iKE5MafT0Q0S++LtPMKBS4Hy8Zq+g9RC9/tqtEb72E1PCFRMglkTI+9N7VssoEB7
tidqzuj3WxH53HDvvikhSVADs9vEdb/pqX5mTQcR1NJZic0SPjQOHa992UoBqBVC
IDMyT4FRN2YH58bkwlFLuPnIspjHWzDHfh0bZpY7dlbnv/fABiL1IYqSTQvyXhjy
3MSTmvjDyAf1hcGOdojJKedii+BDdqcYhyHNOC422p8N91Pp+6aHMRGCfHmdghXp
EcTZLot24NcxefBJQFK97YbUEj1pb0tmIt6kOeHl7edggLPL/bjtCe+aQWzzNjfx
zLVxvl5sC0cQRooO9P00FyNP4LH02SanJV8Fn8CAa3DnxPAqT8OeW63oU/mU4AVz
+ufG9/ueODBjf1UeG4fB9PU2gwKFYCFbUOoUL6RMwXf9sRNJLGaCn0rHfUFqA57S
pWrVTHFJsS6xGhq7J1PqgGxi6am7puiTfUbEoyCjWDCCkKrpL3XfylLY77go4ano
9tuQt5TzZM/RdZMlP4mEmLFN8+gHgdnZV45Cx0+APXOJ/RGCcuHq5REOoHBXURYg
xAzqAL5+qJSAX1KfrJ8QqoFEQf3ypbxhwq8tqa07U9GntVsOvsK4IgZEx4XMNWFW
sojPL1gkdznJc9KYKzI/zXBC1ouN16G2RiBRlpEn3ysLPLqV9JvrzgVotFRcIsJi
P7A1EpRhvsj+zonqHO4LtXZkUtUzdtYThzdh5mdbGDBmV0pCb6tSvD+hSyJ5TqcR
GS69/i1oUQpWDRfsZmPTLKljzli5YrDCRJ6Y0e9Pd+IAqc/HuOrpr3EP6zhdEkUk
YlzKsqZnjJi2t0UQVtkobe888DbaoZkanrWd9aD4my5CsxefKwXk8Qyb4vDYWTa7
7rqrixD+hJB6urm21KT6CVr9+qNa4++VlUz2NBOPq84URp+kcCLVA1cTCu01or1r
TRw7ygL6Su4SKAzsiGzAZojX6+M+ayF8gEBhlwCnxPuZxOc9qXqteUjebucr0r/R
acoKurIX7Lvdr7r+QVncSxvgnbPj0WFwXA0QoXQq/b40uyglsdlvaBOxZw+1XBIj
N4VYpuDh0S5opMp15POOri68ZtQXq3PI//Dck1PQrYq+1Orjgh4xsxuYmwhhuAOP
Z4MdZnR0ZArX3iFNCzhw2Gy3vwQdxxdkTlxT9FmlpTwE59RMWMrilKZrHNpr7Gdu
n3GccR/MthCpIuVsIQVNc3B8G5Yj0FU3pYrd3s2uiSFU1Y4pQQ60C1fWG7RQuHVd
3CqU80Y+xOqf+ppzzERnCqd4yfbDa3hB0TAIudoFDeGgH0fT8p7f6rH4x8OGXCyi
N4DP9LGO81/A/i+uog5EWj9qxQuP+crjKxQcvqsy7tgrDET9ctoWc3cXnz9vapHZ
kuOfoFgaWMAteUHwMd+fslwv1+fHDB826VLYdLTx2G9WRcMm3UIIuzazCk/4omvx
/Reg8sm2Wk7YlhBGt1wMRKC1RHSU9mG4rUpbH9p8++DDdwTNxBZtvuxDK6IGmQok
REamUpCTlWsLpsl/Kdrb+QlQrnv9vTXVEIMoIUQF5h8AZEPu42qD3KV2O6ilSXIc
APi7TlDP+1n5N69hQuceZJrEzLVit9m70NTkOUjWR9rPsQWIEhLpoIUDfSee6hxI
p5Nh/Fmp2YeLOaAVcNbJbWQGeJ9pMMJV1RB5DnU4nxLkeyEwQp5YXh3s23/0AnfD
dtEquQ82NMXRZrt7/ySubm48kQ47bb50f8uBMFp4qE8a35zPvSHaWBEuLN5gZVOp
kUPvXb3+5IWGf42hG7uW45iZU5zbgl6nenCUPV6o0nbl6eldquQ4Kk+F9CIMB5sa
ep4V3rhB4DbQnYQfcL3TkVGXyKtai+a/qaRQUkOdCpzWjMbtKclSlqiCtOodE03b
fo3RVDI5LbJ0GhYE4R9ziM8EQ4I8Wx9s513e3HKWEH0T0ZZ9LnnKSC8CNnOJi6V5
4His/TlH9XSAqqdBBaJOBjF6jRzTChNp45aSKzE/O9e+wuMWy44KlD45+zuWyeRr
7SCdo3jyJdF6L20qATQJx+LDLeSFF8kKnCK5/6QRx842PdyDSd3YwWv5ENMdEIgE
PKjkeBLXvxf/WSLlMS9d8w/bvKfl9kkui5XH79Pvs9pUqn7I5bOplFC141GSEDQN
omOHrU3OlKzfTBuuR8cYWOw/xKBulF0/ckctVHGMIyEqGt89ICJItwOl3FCr3bsY
nBTyxqk4SjMGvQqwWPrlfeocffH9UrdBJfRiMRs/DB4DElOa0X06afj8mbLWVGq9
udod8VqyxbXnSblxF+6lqyDWBOhd1RpAB5sZRbKfEi0LvcD04zsh71nerP9+aL/1
RstrqqKaYvKG2ItfMlA6VZKubIq3WP2r+SY+B2vRor58t0P3G/uId+Vnn9wRJG9e
+2eSrNV4F1YirbFkwbTNZDovnf76VPi24J5mDrNr8aQFCKE2vSzS785jFY3Jnrcr
6SV+xMaUfcjsn/g+ZeL+aCgHFN3XbkUdq3MiyTMAsP3+iSrrneVxL1Mm58zKyAfo
dcSZ6xd6iRPjv30eYW576rrlEMUUNlQ44FNS0MtBqsG9Ehn4dzj4tb2cT41xO7gb
Yxp168/fblUPdt8K3h6MnI+U3BaSWa8lxX02PusPUNVURiYW3WMKRNXO7UkSHuws
chm/p4jukSWUUtzajrXsPvDmn8IaBW+xHUwq2R3mz1ji6bRdA7kjbLG/8uQxw8mh
gg2T/cZ20PywEfH6Dh1mlmb7Ea4EM8wpDNONdlouwd52ElbwQ2WaaqEkkkuLVCS+
AiYknzkJsAWy+3RGn1F0pbVkfoT3wG/nOPn+4cfNWWTkIXGtMloF3PH8S5tym9Wp
AgjbhAdiAojv9FE+2GIECe14HQrQPWQsrBB235JyIsT/mE8mTPJvxVSrGuoXqaD0
F8RA+Ytg/J2Zm97GtkWPixFtKMC1KV420giBR+gdrn+BDEdFsTKWleTYGEDJ0/Yl
yjuU2DnJBWsAvRN8ZiRUL8KhGnRRPiTStRmFlhw/We6IaelY/BuuY3UFIHnI+ec0
318z9eN5cRkNyEzma+v40TNAXR1oS7c5Bk6/NvBp4oC7RyqMlU/shxK/MNM2OGd0
eBeIljwoKHM40Tm24hZG2b5PH5SOX+irfYorg38EW6Roco0iU4s9ejqp5pF2NEzZ
K0z0Dh+lkKc+a1sZQ1EAy6P22Xmxvti5H0oR9CYOx7oxnGqWygQngAUI5w3TbFVU
BJ0EiP6qon5VFqHHKo7uWYP9lfw/jYYnp9V/a87dUoIeItaM97mD2j4RnXWXL7/o
b50UDtIlhaITg9Z+H17ePp2/G2uR1AC7pAerPQUErvg=
`protect END_PROTECTED
