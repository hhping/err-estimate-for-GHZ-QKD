`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+rqANVFML1ToRJ4IVq2tidDWoEoafvyiEK9JacRSZyAyFTJGrzl2uOCDzZyuRZZ
p8IBM4UdisAthcR3Wtc7hT3YYYG9Q5efnvwBPmbK6v/hKDJg3xxNGaETtBZ4dNao
o4kni2qKh1/l9eLstQ3T6GtLMny55V4vrCic/n0OypP7PewuzlTx9oY7XKty6fnm
/vnAkTjNJtYtYevGbglUlcUwzUWdJ4N1lLjtawVJbLX2DcLlw7nStuhYEtqzq/go
bLfHn3KM3jvUNmRaPESwkfG3R1PXEhg5DOed20ymE9DM8jrRd1R5r9aEYKvvGk+l
AyC67I4uCo855y2Zby96XLVKy6olNqSy1oYvXNjqPz4SumD2fEXwkFibKv7aQtEU
0IUtsuTHOJuUYGsnVraWoXt3KT2T6F3zCAeKJol4VigTbihq+SpUcCqLP9s4cZaB
3iayiRTm/NkeHH4K1Sta3MseDRxLMwjSbPkE8KwERxMoY6TLNUSKzzZP4kQVTJ7w
zBimTB07gg6WUag9k5Yv5R9hIiY52rGdDxDrpcB58nAVNSpGkx8RSAuYN3tIX9oT
`protect END_PROTECTED
