`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yzsLFwrBboXJAvg/IUBlZj6JxsT0Q4q79hjYBYj3BI9IwuJQAG7L65/sttf++r1j
S2WoGfaHvRQL/gHia2wmT5IR45NZTli5zqImJMZp/7zD/Ri2MvGnYd5Y5JenE+zB
m8ZqUsEadipZaM4hUWKrKseK9jTxJTlv8qaGKGZrYNQnKjpHZTc9+U4hJytjLknk
G9ZzAfFG2NLoK0nmxuHl0LhkOANDiK9Ese1SXnCKZxCLvH9Hq738MU8PnplEZmii
3fcYBFCZphHiiyOewhnXge2Dy/aMaQHEfedW4XhcfVT6BVtQ53+pz2dMNf1zHxWQ
mKVHX9ft7trqJp112LkmewKq+I62ve6Y4DL+SeI9qtrhEQ6WmDEzq2erwlBuRUOc
gXlpcXZGNm5PbWKSK+O49VQhNC1YszyeC2i3xmMFFwGHYE13GbshmcFJpowbu+uU
AIbWd2yW0qOR954H/n4JK3sZ4nabXK2bJLMHWxsJqgI4SQa+A7IRKqiLmkGjgvt+
djwDdmaIQydvUAF5rsIj9CrclX7DQ2YksSIUwzkYPMikJoeV75WeBUvXNXqTeR0U
fd1iYwYk7ySyiPJHxNy9UIOEM5Id9ve1Uls0OAKTnw25UjcwRgakAb99Ls2DTmR1
wE9mgfGT8w8QfKpi8Vexsiiz/1lEClkthzlbx7lu9Da5FQ53+6W0WTqLBGfyxjuq
qx7F0Ey+me8DIsCe62FOtSsfmQbBfE0ADXi1nq6POQSZpiSKkC87tCupkxIbCfcn
Q6U9ZVpGQoXplClbQ/V6dRxrutwwm/LmW63IhJZWzCO1LUZ8d1nF2JYrydp0n77s
1JwQu2BuclamFMlvFr5misXor7WAJg0dv+Bg1/BUc66P6ZxKecmCTE7zu15bsuei
ntKNyNnPlhxPtuJrnnD8zDUSjDluP3hMtWMiE9nJZbuxAfrTJTa5Z1P4cmR9G/8U
V+J8dE3rebxrjR6+enUAqXCxdRBkDEVad/0stdRych/fo7paRwc+B9l/rsPmQt8y
iQB/i6VMSTxr91vQVdkyorRMcMS2TdWdYjsEdhWlkLhc7gq7j93AZeU1yL7n0p7Z
ljGzqlc7OLvmh/Cg2ipK3oAc5dMKofgnLwYjQ/p6UoMEzXPiu25wEorb/qjtXy+z
MW47SpJUiQJCWUh2Y3d4P1KT+HW+sRzDkinnLri94WDfbzio2J//F7F3pGoMtx6V
Hg6fX3crG0mJ6vqkSuEPhnsYS9s2MEetfSsXmtEyGdigkvMyEZQhFvNdCsyx04t2
73Yc5QkNNc80zKiJ7bpA6aOO+i66hYxaDPctqnXZbZEerid4GUzgOsm2+DV3xKYe
r9tv0YRzYStlne2Nc4Iddh0QuVCnuWzq1DhrhT29dbFZg04FcK4vxyIvSh+eg07A
72x45rb7gf2ulgRpnzIJjys4CRPs5mMPC1zMQOS0st0OWcbUtTjLDXXasupqu6Qs
aKORTCVskYVK4XjdIPRPsYzd63+7CzaibCbYFtCJfqJoixDibveJyndf/iwsTaJ8
Lkax1nT9a6VPLz7JXb/8HxR9rvCMo9YhyxTdXUJ735MAaGdoBBF8qloOpUZX1l8s
GQndsddnBa5M5h414so7M0X/wwmIbe55jyuOZ+BxrQg5HG6CV2YaxfgvHKfJ1NMu
7L/emHbsj7L6vgIElYyex7zuVUr4Dm7CQ/z6Q0Mr4OIrekOW2oyHTqiaf3k6bTM/
89bKotAuJXf8aahVVkQSk5h3pZsWZ3MywEdoZMWW1YEU6vw+ySljZHWkDn554zMh
WWnLx7r9AT9AIKpgek4Do2OH8Y54VjsSoG09kt+UJpX+ivmjHnYVnPDy4vPDTSnT
3dd/WLfvewoCYkLf7U81w44mvOeMYnbVY+LfBzZvSnQ2mW5fKW4MM+YUmvZH/Kl9
lKPJYiqRrb5XHoTDkJrXzdhS29qI2Su/dBUUOu32yLM3J6cj/X2cJuFa+gWSfQaz
Yres0PGSPl8GaDivINoEKkB5GJ4Wv2TqlWaPNardgptb3q0GJPJytM/h2t4+pzKL
9E4GYuc5aOhfHm9SYLEndIU7iHJALJU0lsRbn2xHEujZ/eI9Ak16vBwfYl4mbipG
XxyWmaftVbzmqCmN71UB++N/hT3MLD4DNmg5Hd3pkIazjrKmUOF1kwPab+XgRC25
3RY13QMmbTv7gdg4zAHE4kNyw8Y3/+4HQyS0OXLyv7rPL5rMVdzbWBV8QiUjKJgd
F3O9g11kSDh3fnWvvfU0T+E2t9FLOQRLHIvZpREWjQHytOesOzjUS8D90oR/AiIX
nGJBwZ6+bGmv+FjUz3gsTyYsGKeGIch26XQ6vxMdTXk71LDzq9MyzQOYK46rfkM8
kOmiRAv91d+Ny+A5yNCaw/dLCLmfxN/Ewtd0Z+fi3Iki9FL8F9fWeT7bWWW5Fkzt
AS+CrdxW1pXmSX3iPoYeB2jfwDg41lj4HalvbYyHRyoHsRk9DbsJUXUXxo3dbo5K
viMlQNv028Ba1CrxlUxbSdsa0Sx4c49q3XQrUXVrZp8a5YedTdcH+yj9ys/b9UWW
UKRanfLm0CsLi2+FpuqOpkdLfw6s0gv5kXzOQC25pPu1wSqH9G99Q/6RDfV9wqHM
xBuHWKfW6V2j8KtKQDknmbYc/f8aCO6NGay9bMaZ+q88KGCsSYPdJaK8bIZf4b73
pxSpkcILyh5nEOmwM5U+4S7PvY+LLJ4kCRB41ndUDh+6eKwkJu3ZgVzUxdV/X+Dy
8tUlcLKcIC4DTCy7JgDKmbPw+/4uR+pgRo0UQKMEfEbD9w1z/iQBvvTyYq7eBXdX
0xGaqEMnyJLoQP3vDv4B8uaiE7H2GOTsDj026dsPkYY/qbDcZbdasr1TFT8TNNri
gx2xH8oHEE0psBYO0IQQ2Hh+m277YKnqwiVLM182wnZJSir8g7XMoYxH39z6JnVr
RbY/awL4vL8Zd7pRPbOUnlAjOf9vz6ogxGCwh3CO9Twv9ohacPMwIlxCcgQ9zdEm
ltt2t3rOsBC+bEXFLddjRyIJSFQwybPA27eJHkDeyMwp6N9+PwgHME4VZ0V4WW3r
X1jJ9NGHdSRilfdb/SZkI5wN1aqiKLoygIiMvwkyGdfGY6pRLvBz8dn8DDNq41Nj
eCkZNl+b/1gAOpsaClE0Y2fXvIQYfx7AS5Q+FINeZpdQ82EMpwvnbtlWla2nCEUa
+VbGjAd5gKlzAyl4JdimejgjnRpAqY91s+o7OLEspZ+u0pXMtk6gJWpEIM38JoVE
bfJnnvd1jiF8kYr0oWaM6lGT/3kJadbyMv3pe0LWimwEM9TkgDPUEBKvuPsol9X/
If2VZwFZM4zP9WQ94kLb8rBdXN0N4YyBL4/uffkE8YirNiL93kxpb9/OLTx8wYIM
Q+K/4+v39vQssxinPxAlqigt1hgwZ6x5yREdh0VqC7gNbCC8eRvdBgLGbt3+djHL
Ko8J6se1ItAhlCfP2tqS4LX+bJ961H77LaWVCsQw9nCAMRYk4WmxRHhY8yByU4A/
ipPHwVBRno2R+2pNwar9Ynn2XfsrHlRjZWF6yIkp/NkRk08vAx1Wn4psJ8RBfu5J
l0xlQUA6ptgypSeAxVLjIm8ZVJJTYigzBKSyqMolt5FZWSfC4vknnrgLnvdyY3Mz
0LK3cYtJ2r6A+43loSSmGe9vGDe7/jmUt0eII+uWh7RXJ7uOYp/Rwybc2JVs+Owd
lVxUqw0myt6iq3PlihEGKiFGtVJReUVmY/Yjg9+7O5OUe/yuD1ukMH9MVP+UN8L6
xI/rzLs7WWVt7Urw//2gYmcn5BYCknCKN2e9gkpEEsM=
`protect END_PROTECTED
