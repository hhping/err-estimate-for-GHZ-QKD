`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X60DmuYKKEg6u5u5D5m/51jMWA8fx/Kou8TYKkd1Rn9BAvioE4i0irpPjX/PtP2j
G+d1AglCIdwelboHToCowD3dl+0W4DUh8iTOCSVilP/Yl1IFx8Y5Blv5xfal3ki5
7MWu7mWXRib+DsQ6gCnSbRadw2BhcRg1mKJDH4Nc3y5gFImR30W/oUEupEu+Word
N3wXBX51iLUrHvD797oz3AEhd8jNTpqAK/G1cXw9iFhkggqHEB4izx2GaNFZDQhJ
jBhBMEQJNOcsSN0F1Qlza65JeBrFBVvXHvyjxoyGJPfC9m703CbI/pm7NRSJvv19
3IGUP69KbaRCB5VvfNAdBhjCW8WqkL6glh1biWyfoWEZxk3wlZqt6gwXST+5sRCI
4hhoL9qMK3jDdjT6SRrtra1NrUSjtmHT+LJrglbTSV+NHpLK2Ro+amMIukiAnG0n
KN+eRi0wuGOwnNfLN1jdQxLQEPWlfHMe22ckN5D9+fm2Un/RnYFe+JqWK23qYTUo
/otQAJ4Rl6MuCQU+4DRETRRO9eIwjuP8Oym246jaguAvtKaL04+qe1VHHGzIYdi1
lD1spHPpRTCqASv72OqDwIR/i3KtnOg2i1986YMGtWyFq2DR9c8ppMks/XdEdknI
zpL09g6tp509zRPQPDbz0Gnq6T7yyd/nb6Pba4k1Wq9nO3pgh+alnExUU+2mW+ZH
nyAEUUlyiQWXNkdl7oAAL5VfDRFUXIdVZMGhb3Jo12l1hSEIqGgKILuxu/vepxDo
Flle+PPYAKUPneqwjgdHSOkZmjBRayX5odmNcOk8xJ9bNMtr1Cz+lxsLqNAnklus
rxEsRXAocQW8hj5W4Ed6dXhMhP32CICLMGPLeDmfYc5zcI/Yev499dBXx8O61GEp
NR82Kq7STojEwSPIWM0O9tfRPVtIG9uoWOeSkx2TcJzxh9N36dZsZ85taNH46CFC
UnsSSjygejMrw9DPwg+D/kSOb4EwH72vI7q7B4hc/85NrghvGX+FNJsA7+D297eZ
ONUczRFPSWp7RbGLUq9oSMTlZoZ4M55QnO1yv3AAMvNQTNafM1iSLwqwFXOFx/Vy
CwLQpHoeD3FCXMSsTw164HyApmexgysz9dakUu2SzTB4n9M4eqInwtdm6LlX42bW
3tQ+R2Eh3VOFCiSYegJdb0smYHNH/8hRJSVhb8oI36qn+RwOsSK0Hxs3BhHcWqgV
pKtmRzulHuhszbrUaNUW9V6KvmG5XK4TBqup53QLc9PLxJEX5uzVx/xlyv5oT9CG
I/eYiE9kXayRsV6UDZlYWkQqUIYqX/ppILAB08WBljM4aqjd1LqEpnFrmxbbEreI
fKkIFg9D5KJHkzXkjDWAMoNpOU4GyMpCNzf6ubv7vCOWMnszUPnaio7YKLBizr2/
VxYjB+5Eajbnn2Bnm4VopOFbXo6DeBXGF0FvrIJ7KCfrNowSbRlqgbdOpdxRMpIz
DPlVnLfmNU+NdJvexr/XBJAAcmAuvE0LStmO8yJ6SRBXJO+JQHokiWWTIus4qqBE
EjZ8PmnBNP4b3JpSwXY755aBLbmw6vwt+P14DW9pgG/U0Nz63vAb3G6VpzPmdl0R
eL/+TDBT0O1jCFtLMA/1TXuik/rKa9zYGxFtZyhTS+Bj2qf3F+biRns4xdE9QY54
I07NPN2leCmFXQ6d8j7pAKjeOcyrnRzo5NMhQ8+isrT4JxYUxRFanPl4hbFm9mNF
7RFBZBJCFs5BDrofTP9Je92kxpw95m4nf2IDzWQgNs2ADwprruR1uavbLbSjWrtt
muolPFujUd2Ku61GAZ5Log==
`protect END_PROTECTED
