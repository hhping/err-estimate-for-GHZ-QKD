`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfTfaDfvu/oZDznJb2Y7aTO4XE4/YFtowB8dkNneO5ZpaKaIcIb+zCV4kGHtRpuB
39mWOdNABuksifcThh8/FfpP2t5WiNhNmEntQ6c4WY37gBw/mvAqkkNLke4gmiGE
LLwBK5WJ5L9NH1dMISmLf1Yxm5xTIRpnb0hZM0FInjJ+oLxYsaLdXLRRBLU+7i/8
j7oI3AXJjxSvCICuxpK//62D1Kt+sSaGuo4Ymnv8hF/uWJS16AMQ47o1Rc3cf3Bl
YC4ETQg0OIBuK6jXPJmXEdn2SwTjdDrciLt7k2KvgG4dOvv9+yJpJStcktKW/mAj
gV8ose0IEcp8v0LzIK96XKzRuF2QuJzX/FC4X+iUUKyKYKn3edjk6aw0d+ATQYkc
vNq67i36vxO1XcFygGDnbkTvN7kNr8M1OHj2FrhjXBLuDGxD2OV+jXIfE9+zrYMj
xPi8557FQvRAaDhIWLrdS7c3mhR/SwRrX7egGYuDtsY5lcIVV4y3yKG1drrkPVVh
IdwMr6r6jP4AuoUAKxMQehcMYrxxaXzjMtuwoO+qvAiIczHTIWTd19tfZkTupzxS
gWmLnc8R4VwJpwds1fXjl5EJOa0zFO1YxEoEStreNy/gNtGSJBN2ICK1o8C0ZhKV
OACUzu6RqtLs7PEwEpX2KYN4lfk+uuLumzWsGHcYgGtAawZcIAwkJrHoIqh0S8x4
kZ09LtnQEJqlsUcAFVDd11gShm+Otrk1D3roXdJ83L3+/2fVMNEIyvP0YYw6iPw1
0mkTJmAUkHyuZwTSOsN/jfkxYYTDYNqrTYTIEQ/4653mUjOnFdvWxqkrMSDirXnp
VeRD4aLWc6HfhQJA26kLGSMFcucmNRvNHjuRBRQWKWs1/EuGnf9QJmWJ9zww2MEw
/saYpaARXFXAjYhHsYsEBUTKoZUh8h6qGOImrqF3KwzS7VhReb0KxV3Zi0g/oeWV
4MxBnEMH9dbwYWUmUkmxjWFVXrUUMk8ZHsjh3ts9S8x6AkDSZxOJBWeKjhFAwKu9
IJrmRrpnQMYMePTJfSHqjNiDHk5bSSvVPg+7z2BuIg6FnKP+QeRR3lcTMQgTrB0G
31qL6SWc4psZbRmHdDYokFsRJtO5jGro795flgJGDr7dvrtEwf4xEorhdSku9Grz
leCgQ2Ldt26vhIngeZARlN5SHKWl9s/sioBZvydL5rjgWuDs1qEc+XA94jyjCRrw
JbuBb/kmMnUy9/qX//loTYk5FiFVJlQpfu36iLIdJeq0ic6hC9oLup14Nwnnelyu
+H4v5Vlq9KCt95gVGJ8Anat9ZTb1+3GB652UVtAe7bGyRboo59VfFhEdo/O1qUQw
cCDNufgCnCOio5YjU6zIiDNkaxElK+htcsbGNjS0Z+hK51MHHCSIw0Oeaj5A3g2J
5DRpz+UthBXzgCU5Ny+uYX/Lzr/fY84hp05wTfLKL3bXtPe6X5wtqcf81ZroFEin
SBUkwUaZV07Rm6L62ticXibT0RqNzAfcbGxSXutBl+pNq894OtCYI8fcAGgUJw+7
LcAkv/gVtrjX/RA36nz4YzUovD4+qb2xBCk9RveVkNZFzh73DjHG0sPJyVyeNh5z
XSAXHG6N7dwAjqRjNNe+BD+yPU/HnVSK+EvF47zm1Xo5uFwhwtolw6CqgmaMWiA7
tJNsaJNuHRJwmajOrXpGATyPcrBNDEYwOiVd6MDkgMdjTb5uCSr2qeJtdp8MNUxh
NuZ+4Yf07KZVFMb2Pr6WGlq+xiWgF2jIqN39mweClSEaDEbk5otdRuKCUF/oMg4+
BN0lujUECI+PyL3UgBpALR7WuTr3QtrmfFQjMbLEjMdFsziJbk29D9VGmxisTe76
zbIi2KetI81JCKk+uY8eNw/IUE+vhWjQtcSwaOWFBic+XRq3DhkzZPPLPSG+748+
EwJCgvsq6Od/XutdUjCcLyJaKdiLE5bA7lqZMwmVMYTkyVbopYuiCrl13LI1wvdt
H8XZ15TVueZMe3dSoDuNyppgO8ZEcd6v1CZzyC07bVWmPjGG7CYLYnQCMOIFxYLt
Rv2xhYi3z0Dt51818xpagJ9I2xIHvxzyUDSJUKkHKtZdghcPdFUdBFWXOPWrqSFF
ZM0rgjpECLW5RBVmYjZGGi/Dz9ZZ7IVmEMdG0naIH5ODdITvK64hrKBtJDMBplq4
On4tlvP0O5HFOXqW91/+dLeYc1o7aflRSloX7hCbB9brBYEP9tt1H1ouESkMFWpx
3zNriH1smom1rz/ixuE31QApyQD1C+Oer2Exx5jbMGgDsy10BHHvaot53/xHCLE9
XkKL1zpn8iLcZkdmUseEyOJuF9wSFmOCxvpY604qVvU3tMpt9HVB8n4ddznB1PAg
Bm7RAp67oJ/odZtV3S2XnrqgvkCASDfGcuZQKtWwZe0ol3vgKQhfb15ppzVXJYee
9lgEzplW+mWT9hozUKNmHMgBQdsGR5blUPxIJG5kGPtxgPjQi3us8HcHB3343GOt
MjhC5Wdw+QY6GnUGoBgNXcHST0HitT4mC4e332FZuSFEvFBKSfIzCxwqAapzAHPZ
JE2yLkdU5SLHzoXF32RH7cuGqE/KPgWSK6GjOEJaEmL2X88z2nOuupBJqUfgXmo2
f0eKkDq21FqKQopoubGBFzcRQDyo5RwQlozfXDwh7kGTFyMVDH+TnzZot/nn0uti
BY/puZekiON7yseVfGNl+Y7N24Ju1SGa1usQ0Aq8B4X/pHfmwbigEMebCDGSKRiw
tRXRr2Ch6rUeqeOO5I2UogUPWo8SanD/hu7Aw017CkeOYhJBpNRD3nkSwleHBeMB
+x8ZywwuQxvPNEgc+SH1rUXzvhlTCax4cJiWZdxryfMAnOf+Ii74MPRdnMPNDAmb
u+hPRVPSLvqyYsV151KA4mLX+dSlQ6+uQ7/CrdA/zF3jKTjOyOcomoRmDgZ7DkIx
2XJ2hkI8u1+UifoGuqIZFkQR64hTvPy63LZS3tD1PAFGCS7pwkzc16AALdA/BOQl
OXDw9Sl4HQO7iuL5caikX8EINelyUe80rsuUPzLbXTa5ohrzBPGlwIRpE7aXHqq+
Na/3gVEHgkOaxcTVzg/rdz1GNBP2gU4CCDLV0FwMnoi+IqzVjcJqRTK9jsYoOiFT
egihx8v93+iczmVm3Cm5M5v6vFKxF12g1th96u5nPavy0adWdOxX0x+g46NIsYA3
vZ/rtSMwfFOaQkhbuZi1DLcrMeq5amggTcKNZUf4YBQLvRKRpPnqn1ILLDkAcFEz
J1YmV8hZcKYRYcH8+ff74lDPqao1sXDbFp/hgR9Kqwe9sKYcvvgIGXQvoD6wUov5
WcQ7IVdyrVDmfhDu95TbHu7lbDMnrydQ7FW1SRvkiuebv3N8YV/7C3P/8rjDCtPD
kwbK++oTl3ogC5xA8vDP0plvkMV7bzPmTcTApSJrC+pAsI9YKcHE6pJodLPsHDL3
erxw8z6tgVNmNLV+0wtLsye52P2XchSoVc2RfVfKI3TPndnj7l064pGnfPLxV9OI
JM1XElxtVTZbowR7F/+QgsfXBGc50oahHWrLZjPgVFNPuAtPnbN0y+MHaGBdbhe3
6IZuqov8coQnpdLPP6p9QiSR3gy6uo8PZDmkc0/A+WQjL4N8sX8uHIvhEWPopnMB
Tbo9G7vAh5DlEecMGoIL9RAoib9VguHneb7FaRPc5dN6oCzUXOdkToZdJNZ0rRkB
w2WFA3Ougl0Ga28XpbFm3w0FBtaCgh7dQD6YfWxZ/Ls/9UWYhPDebfbhakyYP2/6
FnhIJdec9t2RMAogfrtdlNZiLXNGRvqkMYc6XVgTAgHKP2NaFi2QsqrbtSF+OLeq
VtXzsr8wZog3/3aHf2zbQVDU5rq2g6lknXi90gQP7vn6fKT2ld+AJdTbVStVRg39
wu25CDDtblYAAtXRtjQp4ZVB/7brQ+nStYbg3swWyQv2Kfn3iaO6zvfITLtpG0EO
ZdIBcZNzGQlNydgDOKc+yExliU8I4qZs5gPYZ95jTsmKXbvcdA0zxw+y5QEQP79n
SZAIv+lKa3jEX3Hxoomrf2hk3BvD0fzbjeBtFqaNLqZeVHFHMO47SJp+q+iZ2k4K
ubV8SvKVMrMoAbQI0EHHk+TqvWFIQnkSqfA6EJGlqKNe2T4XfUeyw6tLLwOzT8iR
Zeu4SpQ/OCVVZGQwhlQHzsIBCv6Eg1FThEyzlVcGyqNS31bfuXN1kkimS7s4rmo0
f6eh1dOlpeqqJfSz7+fNqrcaNikcfKmoeSZQddaZjHCI/s/MFXrCPWd3cf8qr7TX
Jt2siYK95MznStSbc52t/otO0xtImUXu6ATDP92K7gh4218oDP2vyfPQcdWCbYDl
0uIngKm6MOsZPVlVkwM4I1gJ9wI+EY/91tSBCAb2Vv8OHQihOQTvFELgbUQTdnhV
bykrrPq1iajaEUSs/aRCuxMqYjJyrcIZPCsbgkg/2pdp3Hj1SH7pgucdc9Qbn8VG
jeai6MKrOajmEYP+/ZGOp+7Dtx+/A6dEk35wE/mI8902xvuLMcQcwaX+L93/mmY8
9TA/KwZHvY2UqlJCo2a4Pq3vXMbms0DRtayPsGwBsq+3wQZrycUdV+0TCId5MdMG
RocZT/OQhDiLga68OlKGldc++tf0UPnaGgODwCZ17D0a+w5Paa0LYtxVjO1fHIoJ
Q8xoJ/4OmDO4ukvweSv86uf4A96h02/vnnjSYt7krWsx2Tz0ljRsIOlC6otHnMve
0Y55u6q5EzIsjmPum9whxD0ncGMDB1fAuCoCJzCkNyPJ85TkoTjqH7wzWQublucG
e4ywNuLwgyBgIqkmwIEGIRAGpyp5to2UPHNGfYZRkFkfMwsVd5VIhG4UHHksdMit
aswPhWtfixnZSCK8tbtdjBhN4q/PzXKL4wOPfEBUVGI88+0ag9Rn5gbId4hDAkcm
HOeI/L6Le2SyiCk0BrUA4rESuiZE2CZBsSZuL6QfhHXFaURqHs+Gx672Rb8DoY8V
gsJ/7VPMtCaqy22SfXYPDR7N+cORPvtBjbqZ1J8e8K3L8kv2khc5Iitc3N+IZnw+
B8bRRqao49MQeNJLLcO0BC3O406Hizv3UYPRZQQErxOgHWz0UnADrTBXHyrFV0Sw
zwFJtKOUiWHIenu4bTkiEg5LyjJMqhZOH6hQvlqnpsGhxn2YgSdSdwJl0CpBwqA6
Gnd/Q2twLHO04NHtKWzB8pPZs94Kcg7hI9r71WNpGYn6WhUV3cGts1ztqPllBQMd
iyT/jcEteBIYqo7HDl+5OpnPFBZF6l5xRpgtNL7pK5rp/09MRd4c/51kKwRnSAGE
/D/Ck3KsU5NW3AXTA/smgwAf7QxcrXBnzXNX3e5uqwRDBRArRk5cvoxqLGhxoiVL
qslHDbVPTNEXt5sZh5ucNPqCBmalFAd7J5waR+RjA+4gGmJysLMIHtQbghZypbOO
nAGP9d9XO88l+uHgYHKKrXSf0ioIaIQVz3X8b3cgJ5MC8IJ31zx70gA2YMpvKv5W
CrSz34/nPsBCBicFqd/3J7QtCJdPK/qlOh88s/64c9Ziwo5Mhb37D322xhZ22eud
LkQ/XYEP26q4m75Cr09Dh62UkQmLCgtlxOUA2JLiTlBGyy83ZWT8cM8QmBevhFaM
M6DmtQow4yQPUOPOoZCvjZ7WeA1tNofHjKx2bzGVdguZgyML23PnjdDYF2sws/Sl
q0ev+n3dLYG0bfjWxS5ggx6vvUDWKqCs6Il1HA7DAP4ddLcwfV7+h4jGEjl22sjD
SS+wyCKBU3U6WasCswqGIC6zdMz8/AKwzxRk5Sg3U3NxqfmcRC+BTxHIzcag+ltn
q94AvJYmCrwF6SyXXrDVXaAG5jAZVNb7RFNXd6vMfAXCEr1aMonqiX5M8fBVP1QK
9GCI0bahEpBwT18utgnojTmYjtjsrB6aIDQ5Jn1Eue4BuDwKbd4qM5s8AQyKJRbB
4odJgjeriFMfzKmw3Oh8GjohdTUUADKJLpzNlvoyXntnxMBlmDbmcF8evpUXNsuh
KX0J7z6PjuvkBTJrKsoaZm757l5eYI7auB5RQuFelpxYYQsB72XGU46WBuHNhw9W
Baf8KNzcs3xVSufo4SCon11ntSraj7CkO4TDdLy6y9V7hbnFuVlQ3UZgrCZrG2Kb
jSWXQ7MP+agfTb+Ue7f5u1caIWxBh6dRxODMZz1PHaSq8zglK1iaQVPr5n9SwIlW
v9MdxdmbSDs/v0ApTFqCDI35OrklZmDqRZ2HzYwufghQJvdAR1qgItWMx06SOimW
KxFEZtNSzIrfY7HwsSaXPKE8lgivonUVaaXxOLNHF1WHO3AvSL8MMt2n9T77tjAL
lALA70S579Vl9x2CevotY6zQJ1J3gA3/7tWU3PI3CqgCv6Zk2CvOyM/CzFpdMW+i
beBo/b5XHb4ozzY5BItHGg8Ac4ieBVTSz4b4IZGGZs9EagDWTXiQ2GsA/1cb7pdk
z6Kwzmu3JFfMPDgsxazjSMtWU1Yd7J91ay1rjDcUfYNQz2rQNAe704kBDzqXTGqA
S5xDgXcK/y9ZIDdAEej39p2cD0gfDWdzLagbrHiCJ5n5Ie+L4uQu048Ggw9gMRGy
/pfD/aGlRQ/31AHlKD5vPaCYNXHVHBKWE6MwGMP9xeUwdKNw9bULbGukRo/X1v26
pris3wODSIyEx7NWTli8VGr3lfKsJt5dWPGaPdz8JtReMc2m3lqMVw2fh7/YS0j3
/B1+b2Snf4epc8wSVyNKae4hyz9zMFDJN8XAqALdxBIu8Frrmewp9Bw/spENOYB5
64vEwDHKX/+Rt3AAJmvxMsGy0GVH0F7CP3pKSX4rGRk+l+7L9mkvlE7aDT8GrBgE
NFpDmRH+JA1X7U44bdu6eW/azsRZRAMbJtzxd0c9UElNaNepjV1Uk3hDv4brx88D
sDp4d1hpM0VV6nNt5j6wmqNltwk4soHU3jn21cKubtC+u8zf7To0l1C7RzxzbaT8
LBduyyKLMpH7UhkVvYYr4y8KgV6/Eir1lUBkg0a0pqdocmMgQMSUGe1xMQ05hGSi
0ZtCx555A3epHH/CMtpxdj/TK63S+T8wwfJ7jG0WAe+pSXr3sMzBq2VlAlM+BJyN
7lkJt3YbW051FOiFECwWZm/Fgq3rqME9tkAQLjj9kDs2w0jci/kImxmfllwPjMEB
N5NYo6ijxg/Jp2eRkxfYIA0ns4kktc/nRL+X72jhKja9m8auBV/ccJd/wASlzlOZ
6sGRSHFulM0264wmyY/TCg==
`protect END_PROTECTED
