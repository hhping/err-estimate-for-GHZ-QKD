`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dVnds8kOkaek62n9/ve+rIIfwWLZjzXV8Swyw7QoV5CpTdhlQsZv8aTXLe9w4REg
XDHiXqT/oEVZlT6ucjjALzmY7nICvx7+J6Sx8rXr2r5bKaa+EzHtO0vIEPro4yZ5
EMbPtM35v8eihzUkpUbFVrDTZaTTsSdezRs6hgS+LDxeuI86eRE9UsTe183XsAvG
/S3EByJVwPvzvnozyDBYfgbcRFFSNQ6oHBVNLFVsujc4qvmeiJws1yEB90C4UAWx
+CuO3mxdtmPy6h5dKr2UmZPlI/c1WtsqoWwqXmLO0S8IZfLz95jmIqgxGgZfrOqH
WYlzUcwdQEAAklTM3kwJj0lOL7yIggo0+S9vMrJVamt2YpR5jJziotC/JmYJxjK4
8HILlqMFrs/nK6CxeT11UR0+NGQmGAo2xB94sCsdea3xRndjrqd17ylRExJ8zHZd
uQOrT+C2mgrnkL1sUnClslX8IoD6Qc98Vm9jUQYd4c5mTtzsb8j/1bB3qWUlP+a8
AQVyN7rf2BDEEUeSMoOIZIGFK34U30fb5B+imca511B9lEiK1t2AuxCJw2iqmsw8
P+u+ypk2KYsL3NL7J/bzgceZfu9Eli8zJNlUY/YX02WrLERubCh5hqcdRB2S1YTL
3fI9v5i/ePbZmnV3znB0CRjsMiN1/R2J57cJKLv4eayRlY9LySAUEeuil5ys2QAg
FAtMiKLtwuqH+VstgRcz5EgtspHyQv2lpYkcSR03UZkDgIHc919oMB+qnwUudk4d
xdER9EqycAGgjDe1ZFCCYt0lhtJ5Gl7rYXjpDtZnfriGbaF7CfG/aeR4rZMm+oJw
kJ59mvBt54rf6gs7XuZuwKn6w2LiBrP97KP7CtNX0caGLZJfZPiHMSdMTXx0UkYq
e7gxBquFXZw7EJH6UR7pYeT+/k5wCh/c/1sQtYDzLs1l87BYOSzDjhwa9hzw1V1m
/TNdslJhPBwz7TS/NNpJRIeSPzP3ESUKelT0zkkEIRHf94E5NepyqEWEZ+pZMQhv
Lyi91BzRaZQoovWeGnPdYcYFYLVH7qG8m+r1VFpA+V0e3SELc6MATDME1XhS6DUJ
9zt6rXz8c2T6dBV3KOmWR6ywkDHpLlcqG4/0+3cG2FTLzu14RP6sPh6a4H2kPaPq
atsMW+oIDxq/GkgmWxun4UXr/vs5QhtEncF2qGNEVy2YQK2yvpkLXpAidKO8gV6g
aDJp61ObP3dfY38zJbRJ5mpWkDtaJk5Fu56G4ptIgVpX11eX3mOFfn2PRjAFEn4W
3Tl3mGjFkryEYTCnnZuvjs7yIHf1pevtOKu0nHimk0ji5oBJ+8dVpuC3j3mggAM3
rNeletjoOlJXzsb3TZAkB7eBXS7vUvtyj5/lyhHmdXMcDTLwSfBUPRdd9l5RA9Ie
EM7uy9xExhh5Fmb/CU6TKA4DDHmmFhdDCABzpXxqdtfFLvbHWEVyF/HZ4DqAJOMD
wMneqa+y3EUmeX9LRyNSBtSo8UP7e1Ws2GWUi603d5wZoZD0dBvc8Cghs2u6D3n+
n3LQvrLb+TEAM/6qpdK/+imHPOnizAk51LX/y09/fudMCOnn097j20pD/qEN7ch5
t43I6c1nw1S2AhsASCE90xiLLFjBYHjttTW0el0H2suSDA/Cu9KY/E15Bi1Ax4T9
cli6BVgqc6gcOpaUFqIBrTU5a0RiP35pcicVowovkLmB7luluCkwTpgHXsr5WWhd
8w3+DnduQ13QxVFIDS9IivCXWfRkl5po9zneqNHzje3mK4Ucjb2OyJHaZGweA+7r
aUHKK2pcWyPjgGYPnHI+RKgBJ8OZCQscIVKCjTF6rWz36+WHEbvQcDLleqbN4RCw
jOhHN17/rHhBxBHl11Gvv2GVF6WvMvt72HimzuQyIp9SoNTVA47TYZ60oQ7CytAg
DbUtRkqe+RTwwbmlmDWP2dPxBj5uE/p2EB4gMmybK4FL0mAieYcRAMReoKVhPXFg
q1b45+bhOfq2zpy8c5HCA/utQhXY2+r1Et9h/ODFipfH5VsUMAlTFPMleuGGMZcY
hZd2f63oBK+wlGbgzqtpR+GBtWiur3vENkbIk8/gXVkWIT8M+CqOjE2VCjG5VvRC
Q/oNgpe0L+SR4XDE4TcN+W9hA+UUadYe/+dTnlz9ZPQ5N4h9SpVH7B2AMQS58Hm+
HuGw1N5TxQFWfWJHmw+fECmMMvqjefOUyoaIxWGwUDlSKWfHYGcFxS4d4Y2Udb7u
QcKj+0jFm7KRSsBlOBMHwrGg+509ecLoHnqTZ+eYZcWwy7uCyFmMx1XLR0BBiFnV
gvd0Xc9C5Viv+9RzBlLIgzVOhznT4HRLYHKRxH6P2sCnqiGYxsqJHPs1JWDF5kJb
3aCyFRze8y0m4bHA8jeJNU2CfJawoUc2hGwFmIBYIEZo5o5KCH0LIuWCLcKcU0Fd
h6Z7sv0uc+On5SzSolUyNJGnLa9J0VMEmNnsmwdVDtRtTORIKwNFHXbFhdgAjxtG
o2Kq6TRPOd7Z/z4hlWUw4jmvAbRKbWfyohRRHmimJFzC0kHszGdBGG2Q1Op2o22K
70GyZUXmQ9DH2F+TpjCK8tGKAiWn3c/xHXTpmH9I7bIE70kUG1i37vxqzvqTOSvL
btqI1r0JFkwFG8qQ7qm+Gd1SWIDL0y4r+wRQfVsFGvb3frYjQmk7ZUMV+DRrgxrH
obukZm5QM+MwWGWuJzz7CcJscQUuR7U4hNbGDJT2QoYxcVQcw7CHWpnmzD2B5HyM
bcjSFjs9Yf8zxdFQe4utXZylCWodx81t9gXvfcQYR824NuTs01zHmQgjrHYprdrY
2JdRLc24gnrykt6WT0VYCnn57cWKu83Dcm6Dul7846CHaiKeluAxsDxfs+rsn5h1
Gk88+iMdIkziQ2dlYwmx3rThwxDJUV7hn+J1UNU3iD+rR2ENXYJEbUIevf992HO4
v6nSWPcCsXg23NUEfd7B6f6RhrCxHQZownqIygy80lk/jsFFqKgOZh75tuzp0ZCk
hFbwu1nkvV0tWrgZH1vx6sPRX6ZSsahExVIxWaRq0ANEKNzkJHcuDc9CkKfclNFs
xTVtdMjmbTqDdcgbkoQ9XS1yojoIbTpI0UD5bV4pWYOeCxmaHdfyWKTzil/eiQL3
hxiUCow/MMN1WB0kDx8plmh0tOHgdoWUAvfWiqlK03mTsopvPxtZxEvgaVLNpesE
z4Yel6tJIw55AVGr0Lr11q1BT8R1d+CzTKRNMrWtxcDf4DJLnyGVjBPgkgt4WM3I
QFcuWAerY9rTL6VD0yrijJ3bj6rkgd7ELNZz4rKPIjR2eoYOZlnNU1uF+S4Qt/GV
oPnIyvdwetzXD7xA8KcTf3d+hx1HcWGKMnFl+KuTYpKc5bou/AV0Zxo5gIBzCwWb
nDOgH7lT68EMAtPIRn7ekYeaL5xwq2/3zDc4go+nvseaTIa7usKMMHeWIFa07CPq
pqlk3tRKjNn/ABcPaJ92TPROLNGQYZqN1Zt3A08KCcpPMuF0UDO9bQZm9h2wutc3
r43cjt7ux3y+sN0xNo7fwPUfX4MJyoji5EbYplR4YAHMtS3kjxDJEl/nh3ZVi1ZW
ZHucGhw6w4koXw1yyYCuqwn3AaXQWtqpvPrLCM49s9e9m0KWMunh9ZX83YBErrz0
WI0U0Cww9wbaVxuMMF5ZEqY2+CZVFVNw20V/agVce2RCgA1HlydSanwBM01QNQ1E
XIkLbEw1ZumowLFDuG4PWPMYN/BNucshz/L9NzHXohjSU9uipr3uCD1/AkM4FpX8
juZb7uF+JY897s0OTSDb2GOyfCS3jj9yIOTg9CRN2NiIYYfqKPzNvLbuHO1JYFvJ
nyW/NgPqf9RgRjG7Gr+ZykB+dVhiEfRNi9Pe27VU8rWXBU/Cv55RtbHy+ecV+0M1
0ZSVxgkZjWrJuYXxkQAwljNfKJabsdTdiFTxZuAh0aE0uOCaJQFCPL4Kq9pb2qz0
xVbS+q7j6B0oGtyvcUjBUrrc1FOpAdtyL1EicyIgn/3974N7cdej1326V5Y2aafy
t1ZqAWaQoKPzmkQM27wjmm4rwhmvtJmZahcZaE9AVDeKm1PkHONiWLzE3zLQcnRV
CLQ9cKLM48DKg4YmQGsScznwkHRti7K/9ScM5Tp0gPKAIVdADSKtoM4baSNl5neK
qVKzdVmf9wn+d1gZ3BL8QyPCNJ3YDqLO0UFHFUqBW5/EBS/SSuAUYIuDnSfad7uP
PMPr25UX54R9KOBrCMvllyulYR33uDsm3PFzQQ2wLw5vOC6Bv1cJR0OxPrHaTAvZ
NJOFOgfKE33Il3JJCU94n4vsb6GUSHt9fM5U/xNQYkXYHv4ooWcwwIdE8xNHBe+D
4rBLvrNk1Q8utu9aU+E5CUry2HwzfIrjPJb33ilR6CBQXtfRW3bO9IxUqJhW8Rc1
yGVaxcsSEU6Zv+CFauc5TgTIxS9Cho7GFx96fgabOtHh73XjcsM7Js8oiOYPvs4i
MB7Pmxr/Awqz7aM+bGfetRx9uAxtN87u8gU6/6AUnSzxIZ7yvOwD2tUj9JuCpIbV
m3TAw+5lcdqUQdEXnwZEakfoq9NmJ2gM6TFsXUW4IpjOCAssQLto9p8G/zsFkEsu
R/ohzKSWKSMvVxJNqeIhz1c5mCkmTcNCUuL5nvcRVpsC1VEbPojLYcwTVxWgN3gb
EDKOiuxS8GP7aiVFfsDw1NhLYeWaall8WXvNKfi4R3a0WYbhIK3XP9/6cBzMG0aF
J414BnT/hQV+NlLRtgU/Id0CXOY/3sDc7W+BCe+1X8CMjGd0Oh1VWgrJjJXw6TM4
Qan7+Y/9BOLVjxk51G6MwSJiezczOUsvscuG2Cd83Hh2+CVGqA2aPRxnT/LxzvJ0
MYMDCseFa19Tc0an5c78tGWHjWGAs7dPqWYFJpPPo4jUzjBSCb7S+bMWm5pK5h0a
OaIeSzJnrx09aBCPAQFCnup92WoO91LIBaKlp/t9eh6Zy3aMitcVsw9Q/KoMZf8o
o2BW6XMirOAilH0BujSEG4SNqD+Y5N4731UMzgJoOyWTyhyYus1TjA/0oznOffHr
eiqcJhDQ8E/NNg8qLrFmmUq7ArSAoNZTQebC2dlEscoSgYZNOh6emgAQXsVh5xlE
0wb7kpmXxXpcCHVsT0N+T7DmaiVV78LG35hvS7BNn6ftCHlg8kySTGLLBTDBVY96
8OPuzH/JPgnCsrY2n2FoZCEb0hpzjZVD+TY0vOF8R4xBpjHgWpsuScvNtHD+YwGU
3eQW4n/YqFdfEy3UxwD2Qu0e8Vbh5iNp1fS01RyYYb8PBcuJzfommkUM8SGEkCkl
/cZEawLuNwdnDZ3/vHeIgS3HI5HFBk+ROd6QFNcl0h8id6cKQWFrX1gaDhRb4Uj4
T0hAGnjl37IA28An1JCWKs+QEsvPjm3mSqc5Il9yM7pLNtGnNDjc+np2r6iNg3n8
Z8yFn1SMoa4XFOTBIKweGphvVGV9qxb5qg2pzTjyeuDc9Zqfed52AJARkW+UlLqW
JA2VdWth9lepqs0Fk72rorODBrFfjs5jPk8klI7piKsFobSvuSIyX2HdudKXxAhK
UNcV27YazMUJDL2zjnCcz0DRLwYRB9tKn2d8oxq0wIkTaJf3vRva+CCd13RzfTS9
ogITKyCBQqJcarxpac4FbXbcbKKz+Hx4/xALNvyqeegihZqFTiS0m9/10OQfsn3D
Cut8CKvCDD1jGO4ZO0TfZqQ/AtBXhukqVm6ziWNbHORBE/iLGnqGC6rbdfSpAcpQ
ApiEMORFU8rBSczBzoo4ghJk4CiIaN2H4aUyZNwXOniembIsdlT1UBVhAfEAkopu
Ah2vYMsdYqXsGT01VX9tdJnEjAUw8p7sCezTESswyev0qX85yh/vGczWPY5TyaZX
LZ16rHPZ1vn+nJl6dQzfUZQk3JEDpioH8IdzMMSCP+9Ku6wiiK2KYtRdPgYyNewj
Cwd+mMRyWKiK4BsYvJc751FJYHb9KZ1n+nGsmfqBMhHa/AppPanLX7wrycsoIzF1
AUyNNe82RJOD/yF4pEHQOpDAd029PxDJx96Gw2CSkVLrFX0lj+Fprvlc0R+zMyAi
tjFyHfZIjMAkIByaye9DOM1wgzPRYxOV4iEu5Qgf4kU5JZu6cIb9fshOfDWWWP7M
ullN1i4k4HXvptQQZrU1H269HoxGi8/zOYgdB8x4Rp229kTc0TwekMJzNQQI5WjA
M1mwh5JLcrPrl3DnaddXJmSWKjZL/Wa5ORl7RnbG/rFzMQzw6rbkUckvQftDztPG
cOGNkIZorxVY15bhabORPVgEGKOTjw9xmsBvvttPexEToTC20Bvmil1Ke/HXetmE
+7bbIxHMV08U3gmaF5G/FdYBZFdXyTJagFyWszzwx1ZbtfgPp9S416jZPHFQhIG8
3YenKvNucZchZtYNzWMM+Q279seEUFraf2AbYEPhWHccflLqSAcZOk6hnUd4igfe
HaHQI3V1coXi3mApobySCYYWkd17OCmEjSx/OUji5s2Yhc/jtulJvpXxXN5jfsZF
mOE2jh+vsZf6720LaqAovWWRvRTefLM1uR62lHO2O2rjEXsh4WKx7vaYXtmMwwKJ
/WcaxQjlFZlxtqwC+tBdluB6vs9gIansJt45aIhtQO2GbQjHoyHetLT1rmklwnkw
gbr5CACOZZC/ldjkb6gMN4tnrMROAph8aZeCadRD9Nk2QCCFvvq6edOszNQHlA4W
dO3kOlBNsyzc2Zmpfteb+P95DKKy50x8Q3OpemXW/fuFzO2haljJdLLMUBRHgrad
FN7M9MqGfpdkDFMGgrERD3F/tDKkiqLSzhbEeC2oGpC/vUI04FjLepJiC2oC4pqm
uFXIkIorF2S3ZHVfdv10hKLjmex6Ic836x24BX3jHcKoyyY0JSb88dcgVOMhwAIe
cRN4Xn34MRCFmpvM8Y4cicWPoTkF/rW9AUfk/MdKg4pwXcDgJhsH5aKRszh5oU5G
NDpvTsTszsWYifYE/5gxbd9Nbyex2iyFXISp2vP2oUXhuALdAg0zz1/cxzTOjIh6
93/Gee+uk1mB2yDhZ7z2o8xoBQQgyGAA/lkG80we2iGtnR5ENnjK0QhyCdTWXZPz
HHFSciZRAJxZY4r9tDmq3n67xSupjTvRFFIEF932SyAGH53yQNrsJZNohu8++vny
rqiSQxDM9K3pevXhxynChFbwbn45fQl05q5I5JpCaNfPiAzHJpEE1OQkBjSvX6Jx
bL13HEQNUk3AbIonJqz0llqJNLDgstE1he+dGFqf2D93sG628A2vMLemSH7XtgUH
hLZiGH/GS+n6dJ9fAHFiChl36zKjVkO6swWbhTsUYV6+I+f/BhMnAT/Cwr5OjMHB
Je4KCWhwpTzlwl/pNwEbctV0+db2Qz2iqWOt97ADDgIeqHoTF7h9h8PGTkVnodmX
Rw1fsS15D0QIszvOMznDAD1EZzT7JZoPUY4b3oS/g9fmJgNQVN7mxB/YD4guZHE0
g1vjfeZOElY28NLJlGNmIMhBrvu8yeJFe4yLboaGRTQAphcVaZ4pSOjvP8gNMYlg
LjzcULpniIyyo3eooLwu3nHamDl4qb89n0h63X3Vc71iQ9G5Gauzr8t8fJdsSn0W
vtCYTToiAN8DsjmE5arL99m8Ld0TxwQT4iM40CA+36Vxp/6/Bl7y9EQejAXt3OZN
RKt+d9N0kawWTxEhycNVJBNLMXTH5DQWs9fXnR0LTpCZ21qC/2rgPFd5DiFXAwCM
P8PfSGLtNYSDvrG6H2qkwkHRMHTEMKbXvhvNaKwcnAP3YgXK+2RpmgXpjlgH4rcn
dfvJFw7zYjZDxB/rydW1VkjWw/9KAsb2Oe2TBNJ2z1GiwtuL6C7KS/MlavbsE1/b
mp58Mz2X0Hnf0NOpBdmGezkRo25M/SmszSKUJmgJ1xTOiiQtokjZHW7yzGkp/cEr
XjH/YQuRUsn9RVU9n5Ce6JFFX78ysF71w3JsUOSJdNjOlMROkBu/6ffstfnJCyTj
k7XYfRauGwzCg2zza8jaNNmiqK4/xucXgl4bD8QdN+IflLgY/k8JBjiHK3nRnR2W
kMofvtA6PQQqNabybtonlpWvtiieECLKBAwEjtTJIS+4a60OxiJaqTn4HMGQ5mv3
RiNU8vCo3uaGZ/PEQ/U4g1j/s/yy3HttKm9y9eKOX05aVnxObunXrft/48I3w/9m
ZISdOJJtd19KcxNV5s+dzftRYSenxbgcT5fsatzhq4kdkDrx0wd8yKzb1qCQL+I3
QUVKrHxQ02+e4lGqOd8TaRg2ru5882ouQMQOtIE9PpyEB2VykJm7vy5NW6l+5pOq
2gIpGeF9O4NU48NXqW9j9BlFn4dsq1rCQ2e+viUUVQlogIO3bkaIc5AsS5EQkpvZ
648BJY7mVhiFGohB+LhGxIEfoVds0peKzzRHol3roIAxSuipEHjJfeJn6Orp30yt
R9vy62iy4EUeZW8GtEUDdxbMrZVAXtD0xU9y2I1hDfVR5innHOEDlLDE/rRGk0A+
k7FkK9FOIbjejywkM7TtzPemTIo6TU33VQgBOsepy9WKj7BA30uhcnO+GaTQypv8
lJC9/i3REnG9nL4DWOmg/rL1pveF/UQXEw8H8HskmyFJMliNs2iJ4bo0u9OI+g7b
jxCT1aeZHRD4JMZ62lNFe2RQmxEmV9xJ1Rni2puXmlgSrG3D7aZYuRBF2ZkpCbcF
VhqYGyk7i1+yhyULYjjvOEdbIusF+e3N11xeVRPF/eHcgHVUHbo7/hfWOMgyDj6R
4aiizXlz/VqmLQizg9kFkOmZiqQuOLHpbACsQrxOny+SxuhCEJqpSjE5MoTAb5NC
/PTHE1vbCECsgPfvFmWVcnT9a6RwiKOgERqp1Q+2CU5Zm7h0JVQzH40HxGEGSf9d
C18B4tj/7TKk1uqZEIMuTtcTHK3EqNAZg2awbyYkRTVjUkuRdmuyTEV2ze1GGAKj
cUwyTIDzudBlkIAhjhRyZkV7X2HViFWUB5zPdqADykPBrJYiLl5zZt8nkE42kljq
Qb53mD9TKUfQyUnl6adgOvZ+tNum23fNMp0xQsY7f5JaDHK9n6GQGqGxIdqqDO2R
nnT6y39WjlgoGVRAEuJU8uy+56nXxX7gLB4RRjDgDDzhqMkITy4iOGX6xiwupl8d
9MpfzMzSi5dbMTkgcHwwGUT+8o8XagBONMiNVy90EFVaFVXiB2ApRnVu9aGNNNTg
KvbVP3W56ZysiOAU1kG+mL9UJQQG0kb9NEM4xm52l7Pd5BB60+5RiUk51fbxecxQ
XeQ+OblWl9th0nGPtBpZ3LmamlQ40zCeQw6BFGRH/JUfHaesULIR84rbo07ViiR9
slcvB9i8/i9VYP/QK5BLY9ACTp1AqOQB+F/opu/NcL/BgCky/XTnR1jt+Mtb4Vmv
70GlhHT0S2uMJvDsPzqxICXjsAJZonaZf8CeucuHFrETdkC5tIwkqkwArJQUJ4ZA
HDZvw82Hrp+YnX+w4bx0/gW3lNdRVUG+Q+fuE/t+7XpTzTi1Hvl+oAWFP0TQQZLZ
IQPzl28bc97RqjCMubnjJooXw4gD8TNDeUXVI88LuxvsOVYi5a2q4WY4S2Chu8zK
wyrjZFGaPXc9v+Nw2qi7C09Wxad06l/dvre6BwfPrZsNF/kqlhyVamkqh1jgbWnF
fg0E5lUwTui3TajjjfB1h2guV363fM7BGJBHQ6cz4Kd0IyXU//HxzxSPEPhODFpq
dxme54WlWpMyIEh/YTuJWqIuv/QYkuMBuXdDiVa+2Rj4TjspzW6FrMPB1T0m6KB6
i1ZBgDcEvU8sa/AWrLubl0jy2Zva1jlH1N5zdHr2Wr6ikt3s+frdMuprP6r4goD8
8QwhPcuW67E1rcPdNmHeMgKRC7+Gy23BMSLVSCDTS07bNyoG5E3VnoNfjfrI7UV9
285PiScric5AT+wTmTS35F63Rw2CmlA0oCqsvuB9QNKV/NPET5uLa/pHGzU0Q7Fd
nm+GMQXe0IihsGHV+QDAw+0Bd8IctHBPcWUefCbPj3RInex3aZkkAdwaKhqdpT/t
SGaPtL5nMXBlley90LZaVSEvpWRnDgh0l7Z+iTJeqqyS77Mm9FcuMdf/vrzF3Td8
6/QWoih+NCz2spH63NjdGN93ERBc+podmizy4TwH4sY+rk0IOWPxFQRBRcWAJULH
syseKz1LiiHq8qmkfUEyiM6vp8o4zXBcz9rNQue96PJXG2qsGiNqB/AJU0OaEST4
fWk7t8YYpw9TTaw/+kSRpLU6rMUTQGPoYgw0zcMAyowU1UgZHbEBzKcx+pyanJbt
xFDjezs2PneMrf5dqv6AglGEjlHoQ7MOIFnd5MVZbR9anpzgaSV6c0aMs1cvIYSg
K+7TER2+rgYjH9fPnUfLIS3VoNMmGJMQ137FWWXl/rSOUFT8S+nQobUD6JADlYU3
PugEOWBxp8NVwKhl/jCgJ3U4YPYGdePP/Ug7GFMXLW/qoeKeeEpiE3WhyTA4X1y8
b6bZ0sQT6ruSu/8RV7L+Qk3xCDlVMPNKY63YxJTMmCuS6NpdztR1UV8nYIxPq2VF
6iyPrIxRkrMtaSHUceKRi640rkC+te1J8dZtZBMaipouEzbIRcWOA8Qimh55Sixd
9PIl6bQvy4w97vzeqfswop/mMbFZVa/M5DjfLOGehFsk9sLexLhk/0UDnvXNwKtA
X51CKX1/a868dIDQoXIWpOim+QJPwmmhAqA7+vbCxIzU/wRFqql4eV5SpZzpRrC6
XFmksiv8R+MUK3i0CaDwl9ENA8uu6jYJCbE9Y4xS26Py7L5ae3+cvvXwlCNBIwfZ
uizdRBxZ6aGNvUt6ZoJxx1jNurIsUnWiynwcvBGI/12BeAcrlQrfxWnp/eVQH++9
fuPUFfzMcSw98BW2mDGFi2neOkBv8Q5/iiTsJaREY+qygkOBGIckTmRlGUN/V7jr
rotiVv6qqcJf8/c2DoNaw9ZYK28tD6zMrflxpzy7DWQQR8bu/2CajG2XVB6Rrcow
cSqT8TEnDWXMT2Eyd3CxPuI7f4LZqRUOttCqgKSKACcZ9KV1sOyxiB15EaVySlD3
JXfvifDr0Pvdk3fN0tTOh7+rZyvNCCcs5Jsvguqs1Mw70XrAu/j2sXkt7yibQfLu
9D+o11ScHMpO/UjEezAxz9lnLCUuEK2T4R1Dt0z68Gd/DfSCOknbyvp1DqFmJC+q
Rvu4G8qeOFQZpWTplNKbDmJgLdsNbicvIVWM5HPdUIJ+sgHlRYnNmYo2/A5WTjD0
3fcgLSdLC98d7fGlXFt1TDSa/iHzpgFoxg6pm3iMzEG2iftnKKYCMWmTIXzBukQa
FuDLI5NjYbQ29B9T9DjL9gIB0R4U+RaFbEebKur70A+HQgSadsNKmYj39e3mFqWi
Ot7LMy60ht+L7hQwvtkWqRQ9wJ2hkHYcAt82s1ryvup2YmlHf8QyQkR50QBjUdvp
862S+yx0oGInlChIiTqrzUYdxaB3zx85UbR9CGnIzVxXze5oRf7Z5fbcPOaFZ7IG
1Jwn260VFCh3eN433tQsJ6UTbrtRoO4kRVZt/qVKroCbXc+hBooLDEZLTgFSsnIE
eMdG7jkBJGKmUZiZM/Eio6qlzaM1o4F9D7WjGTbf2COuCOZlOXzedU7FE3Yf58Nm
4+p22zg0UCPzYT7sbUC3Nu/WGVJJrqaG9ZA7fdVIDrHs0Xq9Dc1f3eurDquN97b3
za/WiqhUI+7lb24HSShhC2PrQ9QQp0cas+Vw4/JcFsOtdc8Rmczni86CWzlP2eHN
HTLrsuevEVByGXNGXz+2riJY7spM0t1tpY/nm3eQfew8PpJcPqZuzFyHQQheOG+R
J+7FNpP8rzKxIbHsclufUNSlnofcEgd2sZm1+WwQ8L6XwcsI5deWdv74M29VDFc1
GnH2fVPTk7rYkH6Y1uVbJFfI+9cE99S2KB504NtJQPlGfhoZNfTIzq5OAwe+VqXJ
essmPPOif3kqj3Pqp90tDGbt9ngYPFq9QSBoOSbXasKYvtrtVCJtMwkQOgHflzeA
TpcuRyz3kJ6m++BqB4mWDyG5zGB8heljoPLn2jBCipncXPYaGMP5vxEqc47K02X2
tm8U4VapnKZy0mxobbhLEdzdz0x3o8B0bHGf2ZVzF33yx1MJpoQIG7S4UH+Zzt6I
Y+o6VO8J4ngbrfUhBvjvKID7l7U8xslF4zJ3yDDFktItLoN41L4XH7Zq3DWEQHbq
ATdJQ8IZ6Lkl+dOaVT1Q/9qzaErpRIwu/4Fj+SvQ5xbosmxz4BUUfTtvEZfMvT3f
ieS+r7J13GJduTKPcmb+306T7f29WkjjnlsFOwarJ93GfODi84z0YDc+4P9H7M1k
mvUCoOn25rxH0gPUqs4BDez8CjJaQ26pm5EIr8lb1HSa9nZFljRSaBiVBDyPR4eT
dcms9pey2IYbKJ9sVYJ9ewMN1ZNV1VrgC51BjyBfZVwTJUT4wcPfkuRVGrAaLE/H
MO8wrPc75gOTeuSOY1KAWtIq5bCGBGaTFBZbyfc82n4EOAqnWuZS0nODJyG+Bc7l
6b7BiMfZQ9VzQ1Nj86e+X83yujMtj/tLHE5SGMhnYb3tzgYL0vkV2bphv/kywHSN
pwfU2WnIcJaeFQJoCEdE3tLPxpfOF3Uibkz0ZXAWZO0JWpMB1V1J89cMeZI1sDo2
XPm/aqaQnUIsfSkvMpEPgo4yz07Bmqe0idEibMAFDRWQ5YfoyY+w8mEl9d9/G2ZV
HAIlcOHSBWoMfuB2hbpmeNqSp4+3VwAkd15oYXgC5FSWMbemqUSg2heEYRlZ3RoU
4y7KwggmrOqaVI98T6LNpP0XYDS6vcBlyBh1ukbP1bW7TOmclEuRmabPGoAjksYt
ByYTesDWNSb852mQPbtSKqsnGczv5zVFN6a6c56J1J9l2sGGk6cqvjWcLPF4LYtD
3xP5/gujpUnZsZuKK/aOwG0LPGNnFHoTj5zjXoKFIKKtFpTqPN4HRZmkMvRvBUFY
OLqZu2V25c/ANmHBcabbmN2HZwvGvk1le711h62bCBmjfBOFE1rXxpb48gTC6YBu
VPPWJiATRBxrLM2SG2WO+2r6q2HiQFQ3PshWFJpBnon7+5GCZFzD1BfP14axnqw9
/Zo/4Vzm+tCEk+L2uHUXkMEwFteM7lXIgbwWbyzYo/9xQAhsT8YzW45VgLDwy3df
BOXUFizxelTIws15dgQB9eD9biiEUGJBQeDMWaoE4CRIPYqe4V1dlLhRtwI2kC5h
EtFyXojyLoLGBDtEH3ny0Es01D3g7eUkWDPs4UR2VAQ9m7q4DZNcNRT5mwA5HbjW
szq6nMpSivw76IvMjM/U8rlqG39dCmDQqcdvCEkT4T7sr40JQm+ZQAqlsFRWPwBw
DKYMQ0MWyaRbT9wlRxrFeubz74MGEMQ+shKtyjIJt2SbxACtds3pzUn7FKbeOUJG
YZPiozF9PHPrkcB0E7ZQBgJfNoDNJiK2sLpaODLJdyeG0yoeXmWvZPXnQF9IJejB
e5mb+AK8ExD9UVKlEVr7gh/iRnY/sB0EsBd5yceiuski9f1ONHb7M4SJpJG5PeDe
W9b0yYhPUpm2HPi2kbXXaoXYP5ZMyxaEWPvZeM9KOw7S6EPQEqJwBznEYkPaNS66
KwfFyQ0IG+Yt4oTMmMGUat9homUJDwJhtUYLIo69wp2Q5g1yA5pFRG8YOfwkSPMm
w6fGdKC485THk2olJofF6c7ksXPllHlvZsmAzmSITFHkAcUaUNmp6hGcIm7IKqLh
4I+4FG6HeUsTCr4JdCKuI56p8MiKNREwl4Mu4SIEFnVyFY5/RL5XV2o2eV48uA1C
DqOL9GN8URzxsTC3upyva+G7LEZdPXv2GKuzGDIaX+QeXZ0leXuzW+v0fk/jIIDj
E9xwsPCXWB84bHkj0JwWoZHliD2+Ea5ufsKn8J2qL2t24vWvPNnrYwOOJR5W1Zre
oV/PsICDSWYUi2C1mRSQ8O+LX1swG/KvtVxI7SUJZt4mewQikUoHunbBz5286e/Q
IwC7EvsrXvpJo0gVMJoXH19evNq5HJ/BdwqXHCAzNzCos4GeGrxrw29X21l1FL2V
2LBXuokyIUOslsBLoZj6Gcs+bviMN57WHu7+rL0AuQyc8ZtwDVCc5hNTK4T6f8u6
CYsVKA19rv9jZMLrkZ84OF9/vCNpqdIGzWNtRIbWEzSskSrI/mNk7G7iRDWBKuLQ
oprKiJW2bXSZlOHNEb5DToJkArDcRnar+l8pQh0MHi++fU0HrSO39lyF+vxyCws/
WUXuGL6rRZLNkwWJN+qUG3P+E4moIRb2moZ5+up4S/Eg+kHvbvto3YcSSOEORucA
R/crjcTcTwUz1GI8hJKagw3tu/rYN9MMrOhI17leWCfGmzbOda/i91/FYSs9NnFl
5L0WQwLn6WAvn5EqsV24v7FSFkSkojJNIdY+u4ZNzDUgzPgLUN3XW4OvQ446kDex
k707UID3kwCZzBEEfRYmeHfD1Rvn6V2G9U2QdhK/tfyQoTCR51ytiFAPxWHK7ZTI
a15m/wLShLfOoIc4iFYnbaPrt8qtvJBhXzHbfQMRql8Q5tOl4tZ5YzQSKu11RhX2
H8oz2e8XQXJuTHoRojqnwN3Lpdt5aAAsh80hjJ24ddZRbUAEqIbLlAKbG1AM+1UO
fr+DkOib8vVdc9XpuMpJn+CpD5A77Liw9Qgb9flpEJw=
`protect END_PROTECTED
