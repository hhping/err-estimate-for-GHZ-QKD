`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uhLY/kWBRAkFKvgz31GO2HtbgYQjVr22L2Epk+iLrtid5F3zMv96ptkWwCwm56i
umgWDfiY+IGx94uYhbRLyQ2+b6fY1Eqb9LZOtac6A/4tIMd79kQIuIZARHi98bjC
HgkpYGE2ZPyYmuQC+VmnnxJRORupNUaleZTA6ulBh1Spm6HCrwszg3WKeUtXJMgt
6A+TE7RfMsxcNaqaSK+QUf9b4KNgBBb/7GgovogE1d997Y/F6ydpYc/Kv9rlGHIC
qo5hBbKd6QxJ+Oluu5utTvzaAcJL9gNEFdYkMLdBcUHkzJgCnP2M2sBKFNN1Uxdi
gbTzQ5hG37CfqzYW/htdIwAqCtep2g6Kyz/E814ArN0gdd15+E6m4nzRJbMc7obZ
xZgKQGj/gHD1ee8Ka+uM3B/KoA0m9+45+ArgjamShMWcfKU0Ji4TeGRgosfcN/da
gfZE4Dy0uiE2Gx64hOyBK4eM/FOKz8DSLvWgrm61etJwu09P6K/bN2yN9srLxTwQ
0kvTXpjoWQldMBBoJ+XjJiCiTEOFFBhNn3LMX2gtD7t4krCzjQNd0VsWaUKhFp+n
`protect END_PROTECTED
