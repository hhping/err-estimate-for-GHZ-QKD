`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKYdoi0+AYyvATmR6cC2H68jpvsV663Ftrr0EvgUJ0abWDr08CqbMPCnh5mlMC0l
ypyqFUN2oPbvRAqJnl92GpNE9IGPnEUDfojrUAWMrocQS1HQIHmoK/lPSAmzrNnd
3usy8rCOc1D84IO+hrKbGunz5J+CJMGrM/MIcN+mUBMh4BMP3/iIXqm6af+NwVbQ
+QRVRne27ZM5NPONQj9MsT4JHXRDTQBJaUHKKER1aoppd1y43gO2jPl4cPcHuoSh
ubikzTISE1TmdCk6ENwsXNL0s4MUMIyzTDzGP39CBGc+mBNTBT3Z7h3OxqjGCf3I
0UGwI90ttz99UcGBRT2rIbPPlYmEPUzyOBX7fQUjADDONSJt2Qv7KUeR9blbi2JX
2xGPipoHRA8ddZqdHnxHHiv8hyonD8L6XMxzLEFRURfLri++s0Ym6me1Zb+Ja+Mb
7qjtzcSzdejjmawAa84fDxhKulRIC+fOMDZkPAMnmJp2SEZ7jrZchIHJnsb01xjX
TWIwv6aoGG56RTj9WHi5QSd/fe4HMLsKJTP1hu4iOMOoCnmC88WZhKWivn1276c1
CsGxGkykrwHW4/YlI44rGBaUI5Rdgq4PKLZZKFnXNMypyKraGFykoQd/OlfcJvVr
t2MZX/502B0vQ9bl4u9K2ZRxNPIcUvOoJUSWUlD25lmaA0RhzvAMabJ4+QmjOHsi
kN6CQMid15gstnTfDY7ll8wtEqOyvMo59dSu7GR5ASG1vEY+mkSuaOT59Bf6EyDW
RO+mC5z2xhwHT0cda0hfue5mXchzxfWcKW2jo6CVqcspH0BJS/3gcMI74VwSwo8G
VdLldWEvlkhiuKWGlV0U0DGj+kCbh9f7xRcq2XrVUfRYlsCiNXa5hrEGuo8dGSmJ
DluQKLorSTt3xDRvPu81TVRjpzvSFmUa6EgiYzFruJViX8WN3+Tn6lbcxlMraxVg
qbHXkZAyCk4MSaCN+9OMX+zbT+9ZPsy6vpKZnw0hdfDWGmhtR0K4LzPqrGxyKCJf
6c8E/bJZdJdFxh7/2AcKY68sSdVeWP78B4+/U7M51mTRxUCDqiIZjQ31AhC4nmDn
4knuL0FICvmGgeTnOhW1SII+qVS6RR5gMCtZNcbNX5GK867zvMfl+ZVhwaAc77LE
ChT6caay3vVAP+AnI7Bx0VhLwvziL/p3Jhbd0EINqY67VSmIq/cAzLouBeALURDa
PHGEZGW0X89xEVG9dpOoXo4jy3DzKRM6stSYX+bTxNOCFMwGTKbhyk6l5pvwR80Z
lTad13uq/98SAX23u9RE2RYWcscOw2kBRvlS/uPG9AzNmN4HTYC5uIMkaYbGs0kt
q0H6GbBNCUuugG+i5LfOgFo9ELsDMePa9NU3JIfTBqC7NS31R6ksm0k1JNcYjq7D
w40sSEusNo3taa9rGWSZICaaKPlIrj2aUPclxx+cYKqWbsu9l1Ivg7A9XnbG2S/3
ohZUnvZspn9onBdNtM1SagI2T3V1swTFthHfP+H0FLlX5JsUowkPrapF9ky/j5ol
0X9342W/wshYg7FPDXELZkOsIZ+qGwRXaliu4SAuGfh4U6aifO8bUE0OjMyYV1aj
RbEoNNc6aiCdXXHGu3Lqug==
`protect END_PROTECTED
