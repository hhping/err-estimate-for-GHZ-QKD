`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuHG45tP5rfBaaE0mB24pwbFXWFuBh4C5e6ZL10XZN+z5IGGLxtM4H03icEfL+0N
xdR7ytn+jEQmKbM5BMOrg8Ev1UpFoWq5FBV8QdNnaLTSAyE67DWhDt6LFIoKShC9
pKboQbwXte235fXngmDl+Ii/xHRXAI7h7LHxIe6YLd2jA5hVDWywmVP7i3xQfvHM
LKWPaNJR388HGLNsIGXUXJHCyuIrHYWAFHPKA0YAyp4UiFOcF0RE4GyHT3L1cAef
Y1opUIsi3o5sVJ6p9YLMbb+cwEtmX5vQaQpdBf2XlhmFQ4lm2u3AahxmbvEEzSu1
GlNpca4wt+0O1ffbTNN9dkfGVEolK3oObYw+3Wx6C5tyfqQlTEiRgd9CK+fXIwl3
TQj9NBpPCi80/Ok6nnGk7SZoYZsEh+JYio5wYqfZHpe2WdevlDildfw8JYozqYlK
eQAFWkMfu2KAZRQqJuzppbTJPPER/GiHY8JqrWOB4+raWJIjFWBVl+nMORndwECi
IV7ITDrAzl3ET7SEDrpLmYr5lK+0GCLwa+cTFrcoCKwD3cAGzxFjLQBZ9TL51LHO
ILNvV2p8RgM3lBx+8pVcmeuQuz/i70WdXe8OqwH8PtvoECdWIKMBSmcMvUu6O1PA
`protect END_PROTECTED
