`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ct42ZX5Pr6EkUnODDNTRS3NJ5P3tYt/CHMPhKGjtYHog0mR/+qwDPdoX99PnBnaK
1cEHJdQmso3Gn61leQOG/pzj8zXU7dukui7vsFmakJ0gplrlWnio/uFamtmIfk1R
aX6r064ObywXG9paLjEZad2Z90bT88tqhituOZGHk2n93pnOQ4zbqGBL0SB/cBfA
duojmI9SxcqRIAGRAs8+Ndo2gc2V1KkM0VbHftBItoq1qeBsbA6g14nVFQ1seRrS
RSn6Ys3czP0x8JI8Z4GrmznqIFzAFNcvhR1lDIxMuWreOuPd6e/FK/5xM27vDM+W
Y/BOW+ZWs1PRw48ywTbN9ZaVd+YU6hxLX5/gfTrWxD1eN9sAISx9g4nWj/SFRzHf
uZDIP9COpTLQvaTrJvPgr5g2sCyeM6ujYrlg6aKnqJGYQkH6rhGlzY8kd3HDVVBM
iQU8OEpZ0nSh2758mY0xsLBEjLisdrjc5Y9W2JA+3eNZOv8jtmVEntZL7avxYrwW
S2GFyYhY6P7dbpBk7s0BI0TJYuziH9r4hFE1r/A0k1PPhTbt3yAxvlNQcCvfNX6f
QPi21eAjwaG3dDpi/pzahM66TNSaftOxZabXvG6/5+EvwQe37kNN3aWnViR5kl/N
VjaynOQVugWBOgw0ZWu8O8SFY/hQvUWBEOiX7QtMRYHULSFujdhSeXJurkwKep3k
/wRYvU4kLq4JR3rlaKJBvxKqBDjxv3qZJs6XnP7lzKUI+2lwjPew63ts+EQQq5VG
NYAjROrlYG707cYsRAjS9/Lmpcf+ueZI5P4BtbhISxT25qJEE/Zp4oolzAb8vpnR
anN+GVIZ/thbFB9479NeqdLrQ2OsqJM6VebVU5ZvUuQ1gM+FPaShubtiW1O0rYpz
TSXy3lQyyOCVUtsB5l+2lCI8knWVRcJY3YyAhvCxVUdL0swqjmSU7KMPI2J31d27
CBNRwxFSHbLI/vANL1cxV7uPzGq+UDHjIyNKmj3VewrXpXXhFZpeULRsDEMCCYED
lA1CVh5i71wOKrwXK0cTInt1CQdKxGtaIPc/Liq1Cmc7aiOM/5SacuW3ITuRFJBS
+4ZEjwwhT46o1HPCgyLho1nCDBgB9/baF1Sn7yqz1bwneNQwlvbRSPPG2rgaASTd
ukuaOLyCgQJ+NBscrR4C8aNeD6mK6TVZJlO3TyZ8i94vN+0FrlivjpD1ObKrBpBM
9qCzWEzbJS1l0HkQgAfHb+V0aUxr1AL4CXS6/TnRJljUzoP7tinBLJEMs2k5ctLu
XA0XoBnOgMs5/MWaJ/1UzPL8tiF1ZZEFUUNp8qj9eCGB0pGqxVR+w5rILQnOBKvy
RBMqNfc6CunQq/T+aVoRISPmKipNo4kkCTmtuBGcKMEQIwZcpossib39jNzz7Vqs
GmMt1+ZQvqFG1liTpUTEBk/1/LAkLaS7xxxusznwdUehZqY3N3s9jgHXFCTMATvU
CCWjrfI8DpZEUXmZeAVy4H4HwPoBqnqONnGuSQ1i/KJZ4G0bDfojy7EmcWNwF1Sg
aEXy3WsucppLkBi6zy8yEWZhVhXO6c3ebwAy0tgXTygTrOh1VUx2OzeS5ffVIztD
FwNtJfWqaA+V7ardWjD/Q2WDMD244wpb3Od+mcLSvTvpKooIGCb+XofTRf5i9Ixt
eSsB6bv9UFI1XxuB8dhRCTEoFQfAR4pPljyTOXPDbc1ydmUAbJXK9vcmmxQ1KC6r
0kuDVVhJf79Z3upQK5iJ/bS5Mzlx6fmC7SEzvFbMEC2CSAZwo2LgSIHeudfxlkI0
/IQeG0RNc/xCM+R8WDKB1uSNmXE4+obJnfDMLkMBgtWH0Xohb0FV2wZKIQVxJm9b
0QkfJXTtpaUP2kcyLak2g0S8zKD2epYOjLOoqSgIYXjoV3K5Tb2nEAlV4MlXZMgr
PpQ4WTyMlHy0SXL6OBFZLCZSl6hqke6r1F3OgcHg1RUBh5kfhEdT6skuc1GjnqHn
tMUL/wyb6kOFpxN5EZfno799oH6QB3uKh3Nt39PUrnB/o+oyQDgedpQmRoYyxyPJ
Xx3qj8KkCDAc2JNjCOO0zpP4xIU2hVXbmxxLIpJsR67b83syruyHg61/gWCJbNBK
T2Vg5aRaL0ggZJXXORmkgpoHFjasEsayF2yDutU7XsxxDLsTHB6bbpMnEJWoW23Q
lAwAT2gdhgJbU5zE+bdDuwOOew0bIrkQru/7ytn4u2vt38fkaCwCslTbs3hhqAGD
MIp3773gVbwiSbN8gSSltm3jN+2INE7lDbRiGIjXjuCH4f+tsH9VuEObTj62rGvI
CCrIt8LNEpHB7CguVXWqTa4yw4RAcKRmJFauL9qzX6jJ+rsOJex/fh/qNQj5MYNt
hygLIcKXrynYXqp7eV1wlyCGdaQhG8oK7L7n4WaBI7K0EO4qPugBcup+E23/Cvdg
6sNmLPbLUJ9X3fhI82f9S9xAkB6k2rUM+MZk9UID2Pdv25/rvL7qyVcDcTcm+PHK
IxC8LUPLt2Inm4rLBFfhXpY/b1j/zvo8JQfdPtFaeOVm4FO7Ifbm14m3p7kiQXlc
lQnVFpkhu1jL/2hrekmKSKtvcFt3fvpSV20V5bQjyfZMoJ7Cc5z2iCBNWEM1o+H5
QP7fW9iHKoq/2sznrp/57twt2oxV0957Mbg2S9FVU3L50Q7rzav8NjiZ8Cwxel5L
sQy2SkbXCMmhxQgeZ1ziTWfq+r8dscaOsDASti825rJhsilq4dMSLBJ8RDBTO8a8
y7GoWilMg5qyNKSHfABpbJHLyC9FfcnUykE3/fwx+V2Cac20QEjUTozJ1g9jxjq5
ngLQpPUh4pUPgInGpuhl/ZJEbVyd9tJLoA4Nib6AOAmRaTRULjoIS5fxjMybzDZM
+pEMvNqKRBa1nLTpj8RbqC1ZWmEENpDBSd/TTctExtURlJIhenu0QprVNWHl4soJ
s2Gs32rDThbBLffr1Fe9NImDFL0IM9lkFKcvWpObmSnFEPOCCqACxH/oWbRyXKSx
L5TRAyqTaRPR6udRC9imJMvbVNzrLh0YQDjL6Iyfp9+FrxG+34Zpyv29gajgMXR8
huvRpkNNzfin/47/8YO9jscp4CI89XAiB8WnBGBjSdEi6pqYCaOMNpIJTOUIkVVB
NmoAQBJJyRuOrTOroQ+crsX9KNim3D8txJznOSMPIvxBXKoq0NlxrurYONX4Zn9n
PCD0gV2Syte5CtmGQTPanAelqOFkletZg0NOMj2awyntgrxREEcTdFX/SmJ1KsH0
SCeSyRL5BTAVJkR/FlhBhpGE1b9hXDGiQ6l0x5xIPAViG745Cf6zdW9RXp2UeKbd
0HXjwtecMwRbFFqHIEIKCd5uwjmxE8mEs9un88MfZ7QPv6UPMS+D8GAkPKs+FM4O
F9nk45gTMLnFF22itnQwOSfNcHO/JL8KvJdyPddpGzgkZehF8gRVtBGCWJMiuH9o
fg/dsNsFlmi+ldcpYfmb0M6DtuQo0YQiCGtN0n/hARUN/T4BW1q7gPfKWMLvS99W
Iz5J+KEGFWkRWbqJ1bEA+WdeZyDu6+KjFxQcfdAGzwadsvD+2ff8GQLjSE7lBXQU
2mrGA2DN6JSP4XFtnkOG/kIs8Z/SKXGEV80Q+6uU5/AElRwnm0HpU5S2hmZc/hpN
6l0/axxxzwuLSESc9KXw7aTbjWcyccpiwSiWoppQKlkvj+fYopNE99ruS5p6N5qS
4Bt0nL9rIa9MvbUm+ERtyTeiO3C6R6MwVgY5v0nThVMa0zUmL65/fLoBL3KzMFJ2
4RMo2KB65lvtIMTZG757aE2ehXQqQOLgSlLEOR0dmyo/gfoVVewYCBwHY/5k+Z2w
CDcWB4U3ZZob3c58jKpWfjFuCOkUNl6IICMegEM7FRfFkgx3YiSjI2B6tx9evQLN
54E0LwzfPAbfipPHPwX28pRv+05a5hf1wx04JPKjM2HtsXveSCBWi0Ap+SyJznNQ
Zk4Qw0gAo5xA2vCZApWB5tChv1g55vw9AGkiZUGa9kJzoFXIgUB3vT3ROeu9Ms7Q
j185VaihbIkbWCRaujC1exgnkM90HrK1hmDNF78icSVaLHsfuBBU5nV6Iusep3PP
A78nR+HT7E3CTd2dMMe2/Zwwlimkl2xKUpqjmoEDeVq+s1wx7YhZpJ9GZ6QV4/VQ
6egDq86b3Bqggo2RR7CwoRg0/iENuJmbs245al1kH9VXT6ldJf961E4hgzsU2sIm
2aSMFK25hlvl3BToFATsNoaRm0uo9CHWoCRi9VdyKitfbC64DvWIftdZXv/zIrVE
xH0TpkJqLJB+8EpPRd2RPCSdZu2TPv5gUPGeK7Ck7RKvPg6dqg8zcddtnaxyyPml
8ElmWYer8UWOJuMp8h5DKj1YTQ4yea6JTlBZhNAIw50vYo5PeQWUJ/SOE9MNIpH1
CLwi/lRnnydDkpQA6BJtSbWjYA3UwJKd/0pVSPh1uFL+HJmMkwXhWTY5kfMxHelk
ueG2Rp96pzjC0X7J/46dsfaQN1I+Ui6J5EaAmiMzDLW0cB8xy79ZhkrswzKL2eUM
prJfGXJ9l9CR+BYNgEOmtZCysFwT2EA7so3DWd2NiW1iHjz2J2vv0KydxUlFvnaD
+8RNMTj6mpOHtyVd7Ps1SUI0ftQiEmhPWExN8iN06c5wevz7jslhsJzfBGE47Vx+
EIPRWeX1UOm2vFkzuhf1ev8Hn6ptBBmFjPvUn3DYiPZabBI1vRpuQo84rrGVfHXg
vWgMorpFilK8mSREoUsUllPiTw3Y1CM+wznUtjB/JD6JHt1ffNBT5DKlhVaxDBtb
mbgVZjAwLOQAUqWsSe7IkE3NvvCUtn3VU3lViGxYiyQ6Xm8lrEJ6dqEUONVAgj9d
LGIk57tiWLX1Ag0XElI0ucsTQvtV7SSkdntVlFbOQE+qBPSFV0fi0CfAsntIijRP
k68SHwOKVwiy3AYlBBQMNhuIwVdvbNbRaA4bHRAQyEGUuFUTtWZc9VQvuml0gc04
zB0u8QKiJQFZp5r1sjkvD4Wb7otD5cKKNYRnc6+N7zURdV6vWPSA64i7sB62HnbF
xj+7vGsdfxg7PZXraYiCW5TA4Le+rvz6tWpmiTqcuhODH17OxeWprOaR6Xp4Xp6a
Hj5Qm6NqnptAHPJOI0hA1N8jtVKE/gwnLwfg9VCqlhW2hUAoTj78pbIs+TN1+ggu
HM+rHXpmNvlGjqR2cuE3TNLREh87nthTWaJ7tP/wfp9QRx06iQM+LeegHpLxIQ+R
LeouhBeSq3coyrWlA+QLOJkOX7prCtQ1HNOPX1xKP0PeBcboE2lbCCEm0TnTMDff
IEFhNW2RThYooYP1rgmWd95i3yUnXnMGXsJTkUqWczHPngY0mAnbM7cwCwOkWpPI
7sVhbBzofhqkFRo7rb8DwwXGDs2Qia6nP6nKzki76+JQX/FkU+4G0JNEXJmRtX2L
L4QloDheAmKQSOW5Dojjr9eOVSG5HyZQX9YvFzcrl0sKXYzbLUlyq79zW55amvtv
QX95whrSs1E0dJuGxNEW5htVFaSikOD7yfoBcWik4tNxltigu5ymvZ8rKiji3JX+
25TSfiLyfto24T1MZ7jJQ9MylwgedTuqSKhq7sNNWvFTBCqYpwxH1gUwqfDZ6O90
Z4x2ZzCDw/ZfjpGFsyO2wlHN5w5nBcFn9ePJoouXFwU9ZTR8dqvmCbBaBiHoCHDa
vp+SREpaOeeLygKr8tmSnaHqrpjqS5eZtzX2jyyiV2u+iX4cvrH0zJmQJm2ojHTr
sFVRYVrPgQYqR0R4P1A9ZRyibWzHAlGsMXCqH2ekZzoA+MukadfrNq7QSh1psxFb
G/gUiZl43ddtCrDGhOf2pIAE0dlxmIrOKRnMZilGgxAXWXOiZ8CX4Jm+JiyzOReu
7ePEbIC6wlUga4U3wa49xdPsTq237S+ZwMsln1xsY4bhdMRuSCM5nNWUCSj/YxZA
03DzMXsPC64HNRXPFD0h/tkOW+Jbp615K4ZMdMrPjMg=
`protect END_PROTECTED
