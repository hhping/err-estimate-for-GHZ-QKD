`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zlGOYrjBQ1HOZo2uQfOInOYoLgyzQxScCn20rP/5iZN/uzyDdMks9mj8aZBNXaN
WIOgzDLn4we8owYWGdkBFhy9HK5qGypYVZH4j9Km6L7DBXoZWd7Qtqz4T1XlrPGT
7y2vIyMq1Y8R3CDJmLj5yP37pRaap/qa4xPNa1kWc4fHYuzVaadGezj/hMH74A7V
gUm9pDyIr0X2f3K7KXUDjlANEOHAju4IMQIypWfwJiC+Hmj/YInU2d4bplBgFLTL
Lgp4Q7c6X1UOCCc3i1Mim6x5nDTQ9FDHezbO77muiIU3TjsvRSpPRh7BTMorn6X0
U3iH9Og0DntVsDyaTH4EPTvCHJ3T5bkCaOYbxtkFVyFl1fQ2NLsXoYDyc4RPYxxG
ymZWZ5refaQP6tqb9EyfiPlrq8EnT9TerR0TaT6ujmh7bT2wLDUrKAteqvWBpLe/
lHnzKQuziaQsIkI+uk6MLMxHU0A4K9hJ0nF5BpxAHkCYzWLkNY5dehifZgL48Wwp
ni86RtHvSiA/NXk1lauI58YzsGCutIlo092UoZk9ySkm9ePpYREzJG95obJktUIb
xRwdPpQxqbnlAW6hQYUTL3HMNB1dzGMzV2HaAhpjQb/j7rflhguVYsrR2YBlyLGf
xD2SPavFYsRypG4xfYRzdDlASju1omES2SEmzPhFGR1sqw9+sit5bZWkxijZ81wV
cRngp1bmVZTHT+MIvud2kEdLm3QlI9ZB60fykeUVTfl8nJvvbqXpK3pYDdbIIQB+
zJricROw7/OZiVOvjCS/fULulXcrgP+yg1QVbOtyOMw=
`protect END_PROTECTED
