`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzDTN79rkbp3x1+tsfTy061EEQoLjCfG7YZ7514TwFdKflSbnK+TYomkrTX4ImPN
P3uoGxaIS/xeLvUSIhxIPQKGbdB9giC4U2XBvd6MFATiQukvWGkQufedFwT3GMT/
c/F4BiPR7o3rOYcfSQBae7Rl0riICLxWiILU1tEBHDLURduxUK/FEkv36Opy5fjO
iBBmqNpTNLZ1NmHgGhpVrdCh8j9vnSv9mudcjn+hSso5VfQR2cdKv4Vd8yEFkyV7
XZxJn1JF+ztFyXxgVn+2dbMMhIHG09zt7897ACr+p8ONQVNWHf4HZxUHCkbwMuXG
RjWQPOvtb5p7AXlOs7Ok6ZPD07J/uCeS1OqX8eG3LAuj2zg6F56OsrILXPWtIwjQ
K66whu+X1I3QgoL1sy5FLWIyVofq498MHnFJH0VdP07V8XZHM2eyboUz5a4Xmjfp
WCkRSGe6vluOAkjy+jRHSZGdICPRIEK3NF5MPKzJ9BICVqOMLuZrNgYzw6muYKTA
Xm5V5aGVqm2+O5TeLPoE4Zdf2oeSlbQppsJy0aR6dmNMV9pTkvpihs4KpKYK+khg
EuRbMEwHm7pMiNR1386mXKl6vUOqXvgEr/S25dHLXKr2nsMVJIUzR14MR7s4DUX8
EdzExzyPQjhz93B+iKTUUZ/TEVp5KOzjDfdwNsEKDY8FoF9uHPkQU6BNxM2rfIOO
7zGB0EmvEVCiWHj0Cg9vp/fH1wgV8YQH0Eqzr3jFyKaoUPx1UB3eT4u8EAP7IcDo
2+gTJFLU14gOYS8qnLYCtX4OKqCF9uWiVfVVgZgTf5yVVLCgRbYUnehcsZN/KG+M
1AWXInr+TkaeOXT739l5c4tNVybtPFh9/sjcreGU8eK+frioXUniDGYTWrGdxfu7
t/PUQJjCXGiyzxCLLLlBDidZ9DWbaFpe/XJw7xQbiDpBd1qaH1XVOBOePgV+5MRY
KFNdXRhoAsN1ksxuCAIR1hmCQH0zwDDGaYw2SSP/1yfN2GzfdqUi16kDQagK7T6S
sRPHXqIom4pGPcJaFIgrQvrppLAcLJoDlLfJcVBUpb89/uHBuCLOYSL2a12uLGmK
jhOIlJj7r69x7yCBihIZv6EiwO/BFzNFXBdg7hpHuCH9NAqh0bhmrm0FCHCvdiL1
naLsAq2rA5MypLsCiLaccFch8I/cYJdJ6UMOrY8RjBb8Pv6sugtFESv6k5nTsh1u
8WdRM7x3YF9erRKnduTgiT0CW5KFKZ9AI/k6YUW8+v+nyBolF41ROEkaTsyyraYT
Nh9eWmnGAt3SdtrWDbj1b9tmt4EuR0Bffg4vLWv3hXRYB910NWELGFcw3/x8SfSe
xj/eAWUFNINghpfCzexzjwiVc/otkLpGTensH4KB/vyDouqzTxnMqahShbdX4iJ/
bwUEUKNQpAwsQ/OE/kqjv28cy2gLbw7MB01yH0pRSwlMH+W53R5tGFczK6aT8X/I
0iob19HmhgtCUngpZ4Gl9fHGqb+ttU8Mz3I0vkDU18fQEKlJ1daw+8tS2sbtYyll
Tgy1gB6Rc4zzi1NFCKwS5MkhI6MYTEi31dA/zoLEkHIfVO/kwspE9BwUCGmF7NbJ
C4Sz5KrR4ahiuscEP034K5XuhrcMmThNsfwhcjZI4beMDGYuACVIkhJ5L2V4IvLg
Vr+JjCvuiapQTw4rba/o1Y9xj5nbrOpGA0jMtNGQxWy4W5al1jc0ev5wUTbSuOCe
NoZdZVLfgbvOIa4DHHKuIUVmfD5CBkttvRFpaKfVVkmQ9E8Up06Z/HWM+mthq3QB
MwVf6un0qv35XOKqOTlLpMO4xU3XlDvOyRXD5erHhQJoA+v9NamlQMSo9TRxt7ud
KPH77UM3WQNtR7tYyTSu+F9JJ9QN1Ez/6Zll5cPucW+WjAXXg3dtgzBCzI54OOBB
4osp6oLdGH5jRUrNM7cm13ZA+B8+VVo/ZqWIPLsg3/x/bgMSmDUyGbTVyoA68lYe
tAlPprCKH3gcWFTKq1xMDzzVNuWLS3JAh69RYsgxsUZ1klOxnmR9tN6FzM5X19j6
LuTQxVeYVfrDoz/o2kiIkOIx2H75fjHZMu+iEob0YRwsl6OBmkqUSLE3E2+XZctw
Z0O/e/Qo2ahKsnUCOTTRv3rw9DT3MDLlL/5Ie/IikXbGi/h5WEHsK2SJrhjwohbQ
OkWCAI6RLlR/4kZlo2JxwyYVJeC/ZbU6RqiiYeq01B8+6eUUOCrDJQZqWoP1tNLd
ZVbHDfPFobP7h58WtyzfmYWEQzkj8FOTKa1SnqI39f1tZtE1r/fBytUedm+aWqrw
db6pbkHT2o42RA79tv3LI+0SvLSd8k3ebYNDMEXoq4wLC/FPXe71MACfY69vYRDj
ATcKNXQJnl6t4SbmHELfjIq6317KV2WstEtopYK04gPJE3EBpQCO9p5zKIaizpy+
gcm4MGiDedUp0MkY4Z3eg8hFqlfYVUMFx3fom5iv66/eCwL9SrzujzjCeur36FAq
UrYH+1J7oWNLGvv0se4ro0r4NEuadnlmzFMzKZ/iwimLxKTUdbnkXVy0J1JuEdV2
r1AJmosVtKLkEiMuhXxnO8LBcvlokuwpPkdMWQQKUjn20vb2qp0HDC42YofqKi7u
kIu92a+RyCF+Om9ivGcT7O02cXdQgofzOOndTK5HSkYTIhMUarooqI3sVLKwlhqa
lNNIJsiiJSlbUad0f4EUWPbsHVocGhFkdaQPGAmLf1bsdazmUB26xTkkjOkcb9M4
oi2AhnoSJQYQre4nriVGc9qfaBmm/V/vuT2ovXMuV+seOKIMRdnBG/H/K/vGg2Ug
+eYj3oVSUD7LlvjrEG0myrJK0Gm1sQTDALYzbDlKXgD/FQPErK5WulbOVJTsht+X
nhUpbjqfc4RlrcFpX+DzmFM7slyhD/PFaRK1Z3hIkIfh4JNJvqaG9WB1nEnKqkot
4T3ZHrSh/+oyzMeSc6QdyV9vLgsAeZNUo5F9t9JRulMrKralKlqjE3MjaD1MB0Qz
qyzL1NqvOuxLsu4Imrom/HxC9DVFEKkwmoOvmYZNgtg80sRIM1Mgf5lVqT0x+8Cy
tjIZNalbOqskhHzI5uojR8W6JPjTJXXRJ4eI4PNGqyhP/WSjfg45r9FyYtEA+5D8
4uZGhybF1/voLxtzD1Xb0DJvw0oX263QRbH1GHcj6+2dGtrTbmdvZsRP916HZGeo
qQQHgeVCBcD6wNzjNP1fzD8eI7PYjGWGj+xCiVwMeJ8y2PHK7uZ5HzTYtNNMquCA
MZiPxCFmcDCZXo3p+AshCVpioxLr6I6ohGix0sHpR9CnEfKeli/8DFEMoHtz8kMd
/w8Kq4FqiQgvoWBF/kDZ4f64kL4RkBHEeH5drR2VOLizJsmLHHQ1d9fEQiN2/MMq
Tm4OmLA9FgYoj5r/ntY3UhrcstZXRUXX4MQo3hELyk2DzZOvtJRhOSihHaYOQx4U
n/ZXf0iOwiTisU86EXj7Zwxr1qzDrGPBlTt+Dq3L6CThV0ssQOg/9geFvmcQpwfs
sGbMb1VnJ+yWSFJVwVRlhoTwj5uH6JguVb0xBU1vLZPF7XF8rV0Wc6/kzz/gRnrJ
ZVoBdS4YKchu93FyIRzqZyCsVmplZvd43P20OVelX7Acu9dbtPsRMpBUwNUwl6RZ
xN2vfCfENZdVlAx/0AeIkatc3GemB/FRazCehrrS0YE9+kwl6MjkLk+kr3ROSvHV
ielS86pORLkXLeKK1fNiutEuy/y0ZQIXaSgjmQfECTwM0qglURbqf2MgfiAulz9h
xmOuc2sVoxt+PTCZNqF8CieroyKyS5zd3FctR3G3EgXt9k+kMLVuUuJxPH/txR0h
rvvIeRz8tfNqIw+y9MiMqPMt0Hesc6a0bXaxg271cjBVVG/zsxXfJ1LPrnDK0toe
Ljhi1sNOPUCMDwQFgERtOekij51CdT968tMYtQwMx1I4ukTG5qsd0RaqJc4ZnXhT
QpfSH+/cddIDIihxC5hH+Ql140Eh8NDeUq4eKP0+aDUFZA0zOwckqenOna1JHS4O
uLVnjJL/lstvt22EHw5D12hCb8svJjE9kPGmrcWOCRLerQqWT+7VBurmgp+rl7pP
+ohsTQAnEqPACQN5+PSxAjKZ6KOEOKylqmSSZlgQg/q5r0ZqEgoBFVKkYodkhlXg
C+rV5JccDDRe6cZ7oz6fq5yn1R7va8rOpPbXlmU/Nc5JtxR2kvOB12e+eTukKNFy
5FGk3bEA1CbrBI4ZBdOf7Us1C7XCZ/xOE7E7TnwrqtfbT+qiLf60v95Y8tpccOy+
h0PFmNizW+xGasIQrdlpcnae/cv89ei86Va9a0XoC/gX09CeFHDb464FudAW9Ck7
BTvJ2MvOqdwvaeeZkmssSJ4xTV+4vTZ05+LExVsHZ4d2/dSeeuwI+pJM3/7TQpOF
aAvCJrXQVr6WQ1XcwUAZmU/2RRS5kQVXUNFnluqQSf9qyeiJmnAQgmr17uTdDk58
dBJ9B/5MnP5dYWtP7LUPHrj+pHzx8Lu9T+cgJYexlXrZGTppiBccIN8xs51b82YU
ctqo6VliIy+67PgtXoFts4UtVUwN+EW1RYQwuUolVx9A0i/+Tiekq4EV+DIw8c37
yJVcEFcpP9k0B7OGKdUb3+aUVfLOpp5ElK7wQx3uowR3Arb++w1UQQSiOIym2ftM
+eB6G7wxXVSrt8vHb/J/GQsfi9omwusAXTCJ5UKNXJFGmjO4yhwAgDHYTU7S0XYr
Z27E2aEhvQEU6k4k1ivoKJ6DcgzvgqgKzOw8KFaCrZXBImXdJ7ymvoTXZR3vb3Yi
40j3WCF/oHxO5a8vwOFkmAMv52I9VsS99ZAo47EjScBXd1G2W+U4/2kQ+CT4E6Y5
nmhrtkZ4R25mgzPZhc6EbPTjvlUFz3/xP+NDjYLPUDfl0VNRvpuzVdsWKpzlTifC
S1EFvy/Jv7uWuTmkwV+Kdoh42lfwN1R/RyoKyKWQf3IRhTGh7cEdiVGXrusK31/w
JQpktBdhL0jpInrPSr0HLNVmvbbjTFsCEbnqgmOTGlgd0F3tTMb17uRApMRjlzuF
33rfHKEcVvxUS6gWyt7lvUyjsGgt2uhyGCTgzmJGN52lGrkntQgU2Icrfa1hBdVX
DtnvOk0ClNZzP7fJ1fUSmwmL8Dv7HcT3l3RQ9FGy8kNrGBnoIwsawHez7qjQQE5N
YUTrDKjQwBpwMlaH3jSAUn69d4XNrLUgntB5T6f3cQghVGWXcQJK/XaJhp0WEu86
rG81h14pnoCoG/VMc5PdpDX5AAf9R7r/pSNsbzwucX+eRLBFrQtWnAm8C84HyNPr
P3aQ/NLenbDNRgXfw72qB2TtTNwgtjr90vVM/XhHAgxQ5NE+wy7oG4Q/EybbNdhR
GgLvlO+Ci3kiOYQAnXuQU5Vi2cPm8btq1LIChL1Ioa+HTtF7j9Udt5yAIgfsNGYK
8R1dmqQl2KOpSw96iQGNqa2bBbCK3Jv7b4qgsghDzLoPsT7Ds71NvANMueMc9+QJ
S3RVToN/yXo50eWtOaYOsfshlA3fMZVPXmpJSFdxJF6dzw6UEIR2yKvRwYWGG3NS
cb1ih0vSEp4rXIGWtnSo3H8d7c1CBc1P+Mjyp2aDNYHa/GzMk3UmGaHXL+qd1BgB
PyjcO1XpcXW6xtea4QEoPgkcmKQ7U2MviBrNZCVcSVzTIgcfSrtMcWye4hQ+Blun
H25rQhrjDZ5sLdozv/AX9iqDvGfUA6+lw9CRTRBBzyJvF7HpABhEKb2njI3eABpT
kyCjmER/igUjyJ6ILbJOQdHRiVntYUcg3sCexOuKimJfVK1S0jaHmFdjFBqjXE1X
kniemUdLxI70NtaOVBDN5mrltWTM3KMEF91XTFKFUjzuQUfH1cJxLLODf0pWamrX
SaHV50kpP8do47KqWMg3ZNx3JlDttAs1BuI4htrWym14h2HaCpIx15x2WN7we4sZ
zF3TCyecSTujrG05kJFOKS6p+hTFTP0qNfmpwnfLBxGRMqf35M04AfU1Vih0yFXb
KqNsvANZMTbOsSbRjGQ5YAOHTBNAY1II51ZbRguvE3t+yavR9WzAYTszG7JR3Lf1
qTkPqWzZYZ/EnlguOI+Hgzli1SS1ZEsnSuJ+sZN8LegtTVoYcr89Rk2pQXmUJUrQ
juh2DpPvrUQbN4a0MNDpgyPQytnQTzvNg5dbFtNsNvbht7+lC0WyeLCsFoxOC03T
8etddht6mRCOYeW7rqH7ktF4BysuKscS2LuiI0qCiyE7HRSjySjFVrSDZJWGEC9/
G5BXLu3uMeauHur8ZSsay+RmntCsR6Duvcp1dASz6IIfyal88uuAHYH3+ixlHNbo
+kle7vrkU6rDLMbM4XHu690EjBiFrESV4mbzK4J1YpK2r+tRhLtGx37dvWHnzZaL
wIbsc2fzWw9K/1lq0rHhT3b8sjscrh78dLnDv/9CxKyKQp7eNsyCPGtQL3DLltEo
sTignwcinjCeP/Flp/Nn45EgHvCvnyECeGikSDPrOkIVsPCHdw9W1sZ/0cmatVLD
iB+sNGniRTxMcArA/iQOun1i0gPomRUCCL6ms8cAJQbLrHrdjpMUGAMw0+QX9M+W
plTc5dAdkVDqn3zUvftdVpqT/uR90mG/MFf5w7HRkOsiXKCYdCsftUX6RiRf26Sm
+CiQkyvuabfo9QbcwTCLNt2izL8Roxt4R0Je4c7bsfSYnAeokK5jArjkYilAmWty
Epr5pBhwRGcRqf4ePVjaMsEq4Cny+oBqrS9/+8WJ5BQb4BDKW+BJKbvhFW+WWb7e
o/IN/ZhGLYHGuz076UPQ5kyqD41E4CpnKP6Ho5cIjShf1Q1Qx2yyM9NKwjvx8eX8
2p2f+GVFDK5bSFlGJQ+9Sf1cZfg1IXgg05tfjlgNudv0CZtFq4EZRwylDB6SE5CX
MleJNXQjYZefmX4rpo0BGcHb/8cfw/l+7iwzcQgxrYo0Jo8zgShk4YxRuCCEgMYh
9CgCC0FgDwcQnSbo1Ge6XmHXyNxLByh7mVzLGJYc/6qbUmPiPR3sP2j4b+UwZVxa
vxybjML67ELKKMZBduYhLL600w6i4XpaprmDet8nRvraPVBrb0bP3F4rWt3mZKaO
ZmTNFg+rd91oyeMlwpi6I+1PPn1OKZ0uA0iiAQNqvwf/kdw09wSSzIe/Tni1hlOo
uSWElCNIVzYUSzPtpnqwq/7b7z5hblk/S56Eof3AYSqKnTrXNGW+yOWFOVQuJIm0
LJIVb5R7k8cBZKtQxPGSJi1emZur1SWy5CfUzAqyBEucskH2OSygsA+empwkLiOM
jEqq15kSZ01tVpm7uMz7cRsNp0N24XiSPmeQ7ITb5wssbwijbyE4Xs13IGFkeyBH
2hcPdj50lRrOmfRv+M+ct9pktfZ9BdTI90tM6bFWBPtLowvRYRx8ZAxrOquEi8vx
aPueRd5r1yoqgZnolmOgFbeut/hKe2MOtZTN3DYJcHb924aCgXZcbBAWW2wqop6z
jm/Fso/WJugfGUzK1D9eKy6bWU628x9seXnaEcjDy1H+ZXz21bkKL9ju4EKotc5Y
TMdRHSEX09BeMGrUryDWd79OBdTEE2eWC/omKSmcK3Vbz0bWI7dHjOXMmymEBcb2
Cf9H+o5rBKL/bfoS94u3IwfRAFqkD1ckkUd7UTmP4R+wxzh2ecPLTYYoiphclLlW
q17LWXPtAq1imaYrOa0eholeQ1dSCKDAePmDlmtDUndMWBztEXXZrtuG3eTsLtf5
Or27SZutAmrZ8b5YPxaeFmzvJNGVil3qIKEHKzH4eF9VS+ElPd/6VJMMBBraufBc
G5MjodpPo4UFriStbbyVR/113upBpX5gmBS+HPwmvte5v/zCDFVlBofP6pXms7N+
KdWgHBsR8Q0hXZ2wv3KYZNu71YoE8qqB/mdkd3gOxpe9uAmu2xBpNuSs0Eo0vOLo
hk89WCUeTFH6bEmKY2Q0R+SCxbXWb5npgDWgg/0YFAoK9RyMZaFfTKSZlMvyPxDE
Hllv49KlyrTFpY8QuZxHfebROZEjCgvEetxx2Vz1iGLDfPUKX3yTkq2ujyGVImo4
bahQNYXNn7stkFoRb6XRopk0123eRrHKElQWUeGCB6ZG7+5PTxrvxU3AfS8zm6T+
4flzNy82emhYi59zQnBFRFW11hLzqMAuJc5sNR8ZCgrWQTjRJPDbo3TrXvxr9VHk
nX1SgVEShsYwlwolni6yfzg4NcMtX+lAl5HIAPxMGCwVIIDTUsA8TCGsi3VQK9c6
wwpF2CS0LMAWqV5ZOZlGhz3DE+YCZPkK0xXLDAHIsfzCh/q1V30xcRCQmXK8+7xy
YETXOcmoHFRhtxKrKRY+aYPBmNlWMptbdHTcjRC8BN/o+DSikqoFp0RI0rev7TM3
5TRw6W5UAlqfLAl+mlUZJyNK8f3dAN04XgnGz9ODx78T9DbmZMINfnwIRnDJp0mU
JFJD8KXxXWetXpwiyy+KVGjMB36Jr2jyMVjbN8TQhemkLd5zJOtWaBdYQIe7gzze
CEUExna8M3JfpLGiLkz9W+6A4ZQbQgdoQjyLE1elGrS0z8YU4X7s+SM2iNZqJHP+
b+UN3WFQaLYaBh3nU1IYO9gsCrY/ACsOnu9QvbuoExadRmHlPcVcIoKISnSGpN42
PPiWMiIhclblBIaDIKOSsb/pAXrJZ0sFKOEji+jQKPf4aZReAcRYnlQT7YB9tEpT
NxdjQM480hipthNB9jlbmryz5UY+AAgViA7SGpOBwEVV20eKspPj+szWrRPohs51
0I+DSDLvt8wWXY6NrGlPaYTy26epsP4VBotDCinFSaoGyz69fcHMleRfwyEBHVSy
yz8UjZu4kQGEG6lewrMvefTQ5KHmcWIGI8op7oxDjyodmNpA5/Hq49vbTf/bvc4h
sL0sImzPgKQ/xviFDdYO94Gx2G9ZvDwABUkg23HfyS3XbOXk71EEcqKY0pDUuxr7
TyhTTl1EOv221olGxG6ypVaYqFawhMRtttkvIDzvpZ4/Mg5PgIQhMbtWmF/MCvsI
dKXPEdycbvbSitP5BQ0VFAEppUu+a7XdiS1PRAgcvaTIvKuR8rJKUXXkUVXgF9xi
1WDs5x72mLJ3+69apDxURydRTVq9tv+X5kyjIkuR12X5be1zYv9AmOCk0IeccRXJ
C5XRJDJ/cZvMeQMS5Bzs8dYZ63U/bbs/C41rB4q6IVogF7acxGorp2IslaMUo8xv
V2QuJLodmqKQF0SN2GmStXZuV3KtJNADxZP45xpM1JbFyDieVforifn2da5UDLw2
m1hKU7q3Wc8VGzyK0fDNmewtEMAHetatw7Js4KXRnGMo1cMdM056DTTvJQnQYLOS
9Aac8/dXUe0A6B9YW8OE5mHBxGw5TNbkbUA0CLxljS9u7j849hNDX7GXp/zZq5co
oJ77NsCpvTo3OvSra/yLhiaTjgQ0yNh6+69ctr8HPI+aN/aSRDjgx6Rjn8Dr2Z+f
uA6NOJqPfB3JGgOZJk6NGX2eEF0D/decFM15h6uZv421Z7UU71+j+OV2knEpx4oM
HM71zZmD1cNogzh/k013c3eqwIzx31TeXTi5i8BfFzISwliTIurLwes/SMOCPYhn
M2I0EsL6MknZ5Fq3+oQ9HavaM+vKG2hRkXuF1+gabaP/Z4cdDEavLz3Y29RHiS2e
83Ij68T3k7+jtZaP1NEvXghT0AXecT4rfZes5ApLELB990HPXo0GA67/yVJupvbU
vjziSvSWDNJUehW8VVehNovhfxkpFrKjqAGdrKBJFNbuBD+NuSL1X+AKnvn2jDTK
DvkDVNIKK3GVD54dteMtJp6Hqfpm8GWYyP9Pku3dzzSazgVmIMxR7gxMS5x7PXzE
+1CIPj+CwmlkcT+8fSstT2VHiCqMfs/rok5Vr6/vRmjjBJRiQQ2/GGAixOQ9PpEe
ROin7fHu+yzLzbgfQ1ObTs7/zXtoCZQjym7UTnZbXD1VRXcxwZAX3+ow2/bxVdP4
8vSNW3fJnbs13FR7ZMu2MLmGlJRcIqoDzsNgr44/z4M7TMIf5decKelySjFmSkTb
R8ttdl6d5WGViPy5IEn7AF1lAk5BVUKMF+/2RShKHSdUK0mkHSZS+Cx28eZP3ED6
1KGrlaJh+K+Dgdv4mEagS+FKrcg6NCV8QkL1TS98Q4NhGZ8bYYJMg3MjHU9zuRo9
I0TXj8XVjC5HLNtXZLY0LKC4+7ZmrnVW+hk2IdCdDwi9PKizEKIhNlPwImdgGhyG
Ar9V03mnCmDVOb6pqUfouni1dpZSjxoPjcSslPGZCGoNqY6K4rISYIgBZptTLsKJ
CLYL2O2frp/0fR/QjD8/kB6PD69nA74u5lkYvHIDiH28y17+36N0Ivif1OffO+aw
RlD5uEeYVLIMUNboaQjZashoPi+m9FBYTDNyh54A6QwWX2xi4IM4qbHTEOJcFBDe
Ap2Z9UOwZJ9f42DkK2NWNIXP6A0ECLqk1zraN1mOAr1U39w/cPsTH5IRw29ZXQCq
1o8v1TXh9vlzeeWIuqueLbEnJ8a5Q3mbeDeCI+1vnisJ41PfFMXQfytbwZPVqmgT
O8v60I6j77SRKO76Kbjzy1QmZ3gqAlCRwTsXs1VBLrDLfRYTSGw9tBCOfMOWi5N8
Ck9JBKSLevsw6TfxCFibeuQ6+sH1evyr6Fy9+GzmvGgXVSJozvYvIea10rNg2I4q
jXOGlfcNGz/A3T7AiXVEiiofnMbrWyRxWI7xitVlbQ5EHpbCVzQrUNG4b3YTj6hw
HEe25T1vaisGgifB4bCUqOZUoeckPGVb3dcawl0tNpC9c9wfxT96QjitKTWRJmyK
W7HieqeluQasXyszd8v88bw9SEVZAJRxol4lSMQ67GEbwHXhEQ9E+gvP7RhFUSHI
Csh9s2hl/aNuLUr7jW0hRagXG1i8QoIct431SVd+duE33B7EbsbWzBENPCVqTFC3
AamN9KS0+EyVSZjFGbMMlJ9ZqW0iURgdDJth+hIW9fytQRR2bltIz368bT65V3Wo
0oXbhi9FdD7zDonU+Tyj1k5SSYDUbK7nUqIcUJ/PoObyNjGwdGVPlv8OFcu0zfjr
TdNpMiQYHVsulco4FnAAfXy/i5hZ4esG3I1StPaAfYcfbEt8H9+wa9jxaiHwc0jJ
SW5z3ONmOuXffv4cPtb5ux3zfTajYLs+hDn/wvH/xhcR5Er/eOGNjMmLpxNSstN/
yFZrzCuoqL2tfBmiYg4jmjLNXrnkySjbgzPCR/XbTQEXz1pkeHeXHLlxJ9iRMNaR
AKxcVH4WLJ2MkXJmCz6EGSLjLcQST8GinSX5zuWCTkEwdYuSWCTzkXOEW8/vgXGZ
MkhDKi+ViiKU3fV7nPbasPCf06DclJ0Dzl1F/OOz4B21wuhmP0aE2R8ZBEaB64Rz
GcJvhEV/ajK+JY6vrNiTHiYAXYSgP8AWR3KWTeFPyRcIk+6n+M471V5CLizJrfIq
5lj1ujcRcIW7WA/wkFjZ+Mp0mHszXlq0ZwepbH78bF84d6zwhRwuwixcLOCEYj3p
yFfLDl8UtVLQ3u291i9TSYcKiNVH8UtoiBCIT0kTlQgC+PQfZTlz+PnPsc5fM9vD
+8dvPhEKjdUReITbcVObBdScCIDWPwBiwkksJMkdaBk9tnpy8oMEueU3yS8YAQhs
MEQQB+ciKagQYz/iBrEofMN3PgKKHIsxSjmAuDgmAcJF2C8rDyrElTHvYMB+6NnI
t0ZxPNSz6L9eNZEw8viuEGdA7K/4NSS2n33n/bnuPC4SxYqoCfTZD18o3SCi7CEh
L4nylYt/A/QuxfIqIoAHQHwqqpLjYCbF/TYM/mCr/hiPzEpbsBnHhoJivoD67kgH
4DrFhY9j3If+xSJhUrmsUOKtkZFlqIdSH9Li3UnKxbYEjVTmqpGvP08HtcY1JGKY
kT49LrtL86LRELYbeKCO731FIWJMNs2zo/w59JJGYiqdq1Wv6EWBz2dRi/Ph0NqD
mTxM89Mlhj8OKbzJX2WxeHEOMSkxfZGNORU48Pd2kK0p27BX/4y0z1ufHiGkBGmR
mVuvZRUBYtgoKtMocEpzAYoumfGZA8Q5yENcz9NWGGAzCJhZFuOl9asmemJjlrh9
qdGwF7PdyPFkHpbIqLOEcWYSJeZDL4RBgYSi97OmXcr+eJipsCvOEOTXKWSZhyu3
4Yv+aOQvg1msuXHHfpmnqPbMV+4HyKsamH/SkYldH9D3SIX03ds/o9MzOV/KNBUJ
h3RI+8jbnZuI060wExviNVphO4wYxXWYEyPvV4u6mwASFQpuYOT1+rvRwQ4pvTNY
wx5ME5UNsLtBAUZSNDEI+LjIgzKZ/6IWGAnaUxEq5VJra3H4KHH5vXipzxa+Y50+
SB2lQJ7nPj+kjGGQzNV18IEIb3wF+WWI9m4wbZuVRQadYe4P97tASp8ouPEqMTdA
TD/kTU6CefCGJ8I62e6EFCg9prBYumkiBhRpmkB+T+ietZo6Ra2glPkXIZ1q0hcn
g8NG7legD370z9XWmKQa5e3exEj/OUw0lQaT2+GVGvgi+vd8bGPNpbv6bOq9AW/Q
aNJT5/5BnA44f9PJx0jZneCgN+466v5fclZAytEpHzIJF/oIaX99aE6rAEoWmEH2
fkJXGkhOnbsOdiMvn2vut8COmCwAkvdG+OWgPKXnFKvk3qkmh5FsIixiWImXIwq4
SExeYv6iB2IAKmupOHB1lzpfuabkjRE8Cm2/aKmGIICSbEvweIWbDsAdL7ON3tww
n4NXon3PpyPS14SOG9FigX0L+H5CUha8Atci86oM0HEip8oRShHuuIFABip/C9Ca
+KneSv0UL3BTbjczB4v0LBZofcOZTwk47FEZt0zhhdu/aeaAsklMiNTtrZTG7LBB
ahwZGxKgxhjhIOscD0PI2DTRAEVQZHljnrtrSjct2WRr0+HXcakRufG7PQ1z360G
XtAIjKUC5+sM7oaep6Ld50lvX8wKcpYZn/TJiTyn48ReZBGyBs0/+1XWlI/bS5Do
qwe/87+cuZNvcO3w8mnTqwS4B7aGVkNX9yTT0nOVg9bqo2xj1OZJDE+3wgy1u56G
jCW36FrtCdikF4rOfbITSQuOJ+feOVzsSYxiy18WhBWPoskiPkudhVr5O45Fftxw
4/ZgUwlx9jel0Ka0TZewAdo4khSdG6cUIbRdv91aGjDpGisy9wMC97g+/UjxzMRW
gUnneb0wru/yuw8BWzNaH4F4cR5/DAyvJ2BCkeyaYgmP4RJ3qzex/eUFaY447E2x
iJAbLih5wNATn9c2tuV/shRA0LDlcTMrI9oi8HPVWJ/A4TXa+sBB8aIPtUXP7V07
PBE8keImL6LJsZFbHeNKBModOcuM6vpFz10PdpQ35utbFyMDNn6wybRtOyopOzNE
NRSyx89JR/8W0qZLv3kn7H6a6uQyyp1w9Vu/xoZMPSDA9k1xrDpHW12pEsj9Ezhw
pRJK0FnHtpk2wZ0lrNikqFxLeQY20nBDGaAAEDvM7ZlE+6yc2+S5q+MnMN78q954
338NqCTAxlMLp+1nJUX/4bLQdzwFVkyzLFFw5K4yVO01o3IMKFizfszpm2NT/dl2
jSYKo0iA0MS0a7zLDe4oGj6XjvHO8XsM1X23jMj5FPVf2V/woIxW5AckpIYaCwWl
54taQLFAVEnwoDX374bH7KdfuOF+GhPRxhOfAmeJ+Qkt5774Xp83YtqDQJeRmARv
i7JTGuySx2Fb8h3gtEWXXS0GkreaThk0YwBHS1RAptGg7pZlrMRKyDgLvF1BdBRL
OKN7QVaJdPQvm41A24isyZo8QcQovWbrW4ZBrr5OneH2WsAq8AXKjoPX0HgOOEJX
nNXZq1f6uJRGXjeXFscAevDnzMH7j63sKebk/d2jXTtDJByp40T1al5SsNCLzRvl
ioldbTMj/UlmivcjMXil+f3go1NdLXB/S0UlsfEQ/ncBMcw7SQ6jBGZXRP5usLKz
atThuNnW1hlondU6td8iTFOJ7ctuG227dSiXibguQJQSoVNeihjtWJhy8WlGCofT
yJLT9rfLN6uWlru4vrnjNDljhxj9s+OviLZqouktpus0Rjn2c4eF2YsuwbIIDyVR
rNeoZUmfpEBs0gC4fndUIAI3ZidOmJtlrTkHr3IB6z61DKbHRKlXhSCUyaRlLws6
QDT67H4qJE2GOXqGNCX1KC5sNi4x0QJZi7TTpKP30jV3O+NQv+O20BtyF+sNNaVu
xgDV4cfPzZvbW3yjYiiQpb7n6JuJsym0zQ6HPylkBXv/8+sTi/gZ/YhB+74dZJz7
ktjGE1wM8c2gm8UCd6XU8jTp2TXOhDkkxtK2l5fg+AsaSrei+2IHcMpmVxn4yNw/
PqCd+Y1Fq4oO7d/KwgIC0wMoyY3JeahrvBaz/rxUQ5G+skxH0vFLHdpb784NZLpH
7vJWjrYU8VChkbjFyqkp0pc1e1J+bGNv1pKFCXarBJeGm4nlVSxc2wjj5ZAUAszI
Y0kd/8u+eBoM0WfmMSatp2yRLml98gIRQxjZS9EV4BEEM40pQca5Z+WacesZzG8E
kW0qzpFvpalPjwJaxQGTGAc6wPD8OadC2elyExbff3CbNk+oPeU7K4828cO+xMAO
u1a2c613KJbyB5z/26CsFyBH53P0JPveQT7BlUbrVkaHEArx7Vddvlz3t2avGy98
JsVK623g4wyGW/Rmj3CFXG6jPmLieM5DjWa5TJ649lJTjIgBsJniPtKx2RFgoWvo
qEXQ1Oaomyr5uxzcDeXYcjFKmNEjaClMwC/ITdbh+KPeSEwILtUj6cnESfHRXEq7
nJlMIskfA1KHT/4ZzTZlB/aQFj3D/C0xXJysNHLZdlFw5tgypgOYwB0/rkxXbGzj
pQWYpr9z7ZOgW27HqSY/2q9bFsxQFXcv2BvFBQFBdOgmubz1U/jnwFbMoIqlNmQ0
AdyQoIB9e5lLxs4LaCct8Ts11kB5miLdepzm5O16ncvDPykSsjv+90uLkJcEt2ww
KgsptzrME+EC8kFoz0MqX18xPOQoOf73grzh0MwHPD+qle+cqAY7SRIkcuP0eKB3
XmZ4nrECUMBkw3WCivsem80/BthipLi8rEUwCOxGdESBF+106i1Dlv4Ta3NHU78+
LCeO7ZTH/dkMS81hiKb7U6ZNPp9dluhz/WIZLobsqR2qQ6s89hgKDyAeW2SR/ukd
JDzKeE0tu71mK8shVlu/lBIzdmgxzvqetKQTzIMpvMD64jJkUjhrngWclPvKw9gW
N3BzvH0W7+BuMztFTtK6q0ll0D/5GfB4/pXRxk9aHdeDv9ApHl0UJYRzZ2nrPbIQ
dE/Hsp2UvAV6S9rZ4hpW4b4Qjywm/s5CWuW3S0u5t4rvT6Il1TFl6IJSTvI8e770
520X1V3NKt0ZE+sfGcQiCgYL7WwMbVO2NS6KuIJkFGBg07tNTqujKyC7mSJ+c0nD
ouAAj9BUe1zW+e+AYcjCxIH0laGyUP6fFHgi82etQ5razOZVQH0KitZXZI6Cvz4P
p/DJqKB6Lk4jR2Tr1NDVZEcCfh1P9o84ENv8UU2luXByAvfrCPY4RYmsxiCZ2bpm
qDdxP9y+z0zhNryMHXnGsNke2vYXeL2xTy/iaM2RRLSkfM91PLKrL7DkdH2Y17/l
MQprxDCVYrplZicpMoDkLExHkrJJYF7lTa64J3gNd+DhmG+T/deDVzPR+iramqwm
EuvRytqb5vPZJEt2Jyn6N1GfmL5UsHr2A8yOJTqyg448pE9utGIakM+8NxEXH3fn
g66vQ+O4W1YEaB/86UGV3AkhNLyWqCsVReR3E5qS0omwfLKjxrwj9kbwF9ekm9En
e/PtmH2UTHDcPQkr48L8drN8QkHPTryleOcPS74iJ8IvWGHwuX0zHFhmWj8FuUHU
LCv13C7DrbfXExyctbzqWD+hLPFei2z3ruw9qAfnfPpTYwky0RDnziQa4c/n14Q5
DmpIxHH4KvsgmYBBqKujvFacpE0JQGiRvne6svHqpwLI4sGRpRJ4nMBb8UNRIdj7
H5tdlNcxjlNCwKAvNPWw/LnEwSJe3AVLeDiPDHYEAmUNZJF3ACFrkQL06RKbDSrr
yd/+yXzeMaD0piQ0b7/nousheMmzw7TLQpquU8mbuOVZ3ejv4g0kCU2C3WCKKt4C
mHWDOk5xxuTd7v4NohLgNIfUXYRvOQjmSSLgudSnIyRIjnVZKIaburLvsn5R/Lp4
vo5KQ4G3CcIJLYRhQyR/Yf1HhuCqyvm1Vys07BTidjT0085qhgnbjAjZtrk5oJ8p
hAJOhDuv2FFEYPdmYzXTNSfMnD9e4Z6/jSGU1UxYhCvclIwHemHXzS0SzXPchqDB
l5gFEH6Xj5BrETLHLM2voa2bpQ08NsdpNAqnlHi0gt6Y5be07YPY8PxO0cjn3YCF
Z4fjqQZvkj4Es1PD2fxw7FDlDnU1geEH/arfFrysXlZyAR3NCB35ZBVb9spmxrGT
ibMqdaj6GxCWgmfZyjGli4AkK8LEBginzQcb8w5syJcnG0LYzbAYN4T2jla1XfnV
bKq16Hizy/iUdAdbAq0WCuzwVKNgt7cvp2hN1ChTdcPd1OxETwbQ5iYeYhLLYtuD
xp38rqxeGrP85IgUV/9+M+IaqzciTVsGcZICd8rk8chyk+3fd8GtZi1dmS1Hnw7F
7LhSSnp/v5Qxf6T8nEVmyYwGXyB0arbaHtUtqGbc3X5p8uMjQ5Yb5fx7bwxj4v7h
2lCmgiM9tvlZ3Q+G0sO+MHaclG7IXOQwja07BWy56nlmUlap5XID1QFY7xifV3zf
LLc+HiKBRTo7lQgKo9GkhLj7uztgvb4iXV66aGR8Kst0nW4WMk6SooWIAl23GGJG
jy6IpvOiYMzv1PrIlAi1us2FxXo3sbpCD8fepsC9lWTU4QjwUYtxM7p73spvNOsr
7mbq4M88fHoYniulUkectbOfMv8Negr8fmgCNU1qV/e38t7NKbxTXfQqZ2OhK1dl
ixZVacDJO8E9GBDBlq/dvpzcFzDbmRFJqCrvEO+nLtwEFswZa4nwnIoDvz4AUY/A
lMXh/CflFNVBIj4JeNukcU5kV605cckeImiy/bYLZKVKy2bJbqslH1j2vRlVUk6l
KapYE+KJU3DD3UoB5DBQ5QFsRcY+vAngpDOF0g5ueZLGKr2eGN2FnZMH4xsiHJ0/
4esQSJ02hZx1FwAVWHlqSt+NRTC470vbNl7vAKVWNN9gktV+nkbIo5wO2i2KD47G
3eUTbg8za14fwU2FgieA337hfvDCjHMYs+PQhlNI3Y3jtdKp8bV4DwT/0ATXvn94
LufJ6/FqIMDGFO3vl3X9zICJa8K4SadcRS/tBL20bMpLujNmdrgCnVUoVQCFcUJO
UiZGh9tMRuZ9pgw1C12rDLeuE89piWwnQ0VEF+A7RO69tM00jSWCr2fPnLRplhED
U17aUWRn8VlRUd/3SliVDAEBttDbMEtnEty5HIcDIWAQWLytZohi1p3y1+ye43Wm
+fz0QEi4nz3DXhbu2ZOydDUTyrao8YRX3s2t8wroDa86ISBW4MjhPfGDWAh7FIap
1UgO46fHyCrrUirTvPfJW3tYyQzGA2p871ToGMGiNtUXnDAicVwjfb3tL1CwPqzF
E/iMk3Kh25Gw+pqMo8Wr+/2f2cgKQvMsZDLK8HGv4h6dhYsuATxaQa9DLRCLazVG
17PWR0t/giMUymoUb/cEBkx8DrxohD5ksap5Abonf7c1KT0ukCfc73id+MFTCcY7
PgFMGf4+xShmZtdE/O2T2PV5AbZERwJd1Q20oMbnsa70HgFGwOYXTtONjnYtw1LM
gORStoolfk2ZMTImDoH8k+CorJfON0NrvIL5ORuKc6GrGhuxAN/Cw19E/M/ZGV97
iFbGNWfEeCOVHd3mLcH824skBMQeO4cXuTIYOAUposSL/L9g6sh2C949F+ZojYDU
Vo1OHq/GDTrHIvT9fgOnWH3Pzq9Pw3d9whqWfkVQo9N123YfnMa/5y1UyugUPitE
3A9SuOQ8WrYYwi3J2BcT/iXVsRHyb3cZw/UJvDMhJ4sdFcvbbxzeDF/RQeiAj97S
T5flkyF2L5GWtOTbP/dtwPr4LFyK0UjL7/zhCeZnXR2OBlt+XyJb++dZ2YSc6auA
jsGPJ9VaEjiimIYEFECjgvn8SX9hMWZ7a4HyLzirScEaU6bfOPR/dyxb5JOeXDPU
MYngrFZQcngNDCeW7/SJ0ZA1AACArlnDerj9DgFYj232zzs2vD4xnxmcb8pfxzuq
PfvEM3fXQVzmUrvOIl6CCkoawtl9KyyLAc5vn9FfWPKvMzDscodUsAycwliEqblI
67gHO7TNt/+Unt+eDcsUZMKW7kf9XhwUDXNvSJMAVzW74HC477q7sP+OkJ8fQis8
L3r/K4o81uMz/bw98UfkEa3k/HLRNFFcs8rU4C6xnQVR8fW/lLz4yxZOZb7r6mSu
AAc+JN615o4eK3MtMqhb32B61FSwD1iNloMmp2NNxxJIskXQ6TovM8wQ/II/tN78
cMRTc5uUxlVNLEZfU+MAXUMWy+Y5j0L9dHbcPn3RaG7QLDnT7f9RkpVB64Chu68I
2lYZ3fUZYbHTdwkjEfq7nECOfZxZDzDiUD283Uw5QzW14LegYyhXnwlBPa68U++E
iCXSDN/Rfzx4pOzrTsOMBLHBCdbzyFVi5OMi6N6pCI04VxMdtPYHgn4/DarLAvv5
FYfv57Rx0KveQ+WlCdMl2pj2V1Qhm1skQeWfn0kH7paR1hwSQ6lQj+/A3sM69Z5r
FERO5KobiHLzyET6DKt/TwRg8q4YqzavdRc0zL6NJBjMncU+2W81voH28Ev9LXJU
3k85PVlK2cpvpOxJSv08fafHjMcjR4kefEC0wrd1AeDWbyyPP4gj/oOtFTKR3HYS
b06Bl5OO6kKQQonA9xY1SwiKn/RoO0vsAz5WNwYSfR2Mues3CVHnjx/M+iW0V3g+
u/VoBVKb3DGq/c2jr2qj/232Ed4oScGjQcQ/9wZ2j60x9hgK9yp7aszfxUow3RJX
EFSus7lCE8OVAwbJy/i26b+DD+Z5Lw9d4SeZFibiNeBGD5d7Wc4gLxp/qnlm/EZo
iCyDlrrGDf5gt/OQnx/Xbtxj9jT7rnXqFm4pQSPybNiLcky9EOm1uO+FM9slZSpI
959xiTO83fUP3anLS2zCeDyyrKdbqe2fRkDACsTrhsCY6M0hTcZcFwTGdL76MrYh
2Za7SfMhw9Aavv7ZzGjYauv0AbVSFTZ/qzd65pjq7Pft8zsgHHPO5RI1ALENvAOW
ETxZeqBmZgIJYXWWCypUGImPEAs+mF4QuxDD8hZXD24tydZNukMtIkkbRAZMGxLd
2H9HJvgfgixl4qEwieo1/giSafPYS8szt2ntXDQfTUuAcioCgPpAb08aIPQSqZCo
i7kSGT8g32GwLORPggDtn0TyX+pwtdT5f6x4KLXBX0LqZMEhV/yZ+2dgNNl2KxbR
MXVhUYkv2qYBlPin+LVya+53ZayqRQUqdFuAOh+JJiq2OQhHC7NhcLuf2gmvDgoF
szYVJ4rz/Q6V/Y0NBtZaHXpcomi7c86uoqzuc9CymbtxEnyQbMCN8hSbPV/mettE
XGK3vSyYQDkcO2wV4PIlQkMH1aqzBFpTyFKS/NkTiUF+PQF/9TzN4j2943HjWbUu
9M6Ti5HlXkd1h7f62x79IARYDOiFKOs/M3i92XdiQ9hjBKl6Qieqqr7xezS/SP/W
VdD6+Jlt7lkDHyVJSE3RcO23R7cfUflKAkzMWLV7hBUyXhHqIOUOKMUxPadWUgZK
dIsrTR5FfdbmHBw+VTYo6v+5C0CLS/f9JvWku30X6WDubf6tCtyTA/35gTjVm6rf
ZlPcOidk4FxGD0ker5xR/y2tajSA10fFXjjV7FEmckQR2IcSEmPpk/UMxIdaUqG3
pz8NnPl234Gsg4wgOcEfT50slsjsn3xEQ4dN/IOAP3AhjTNddwyX2ESUr9h23Ygu
tjCpGelbVK5rCq51HssXFPSVFFCGsHSwn3dL+2kLwMnKlhw2W1kvXLFuHRC3eteL
cWxGP8AFETdroOWnoEDtPcKASdnzxCN8bEcYeq3Ilpwk3Gr6GMM9G2ikoZxBx6qQ
tRawyiLh1TQMaGgS6dM7xo+Wt3Fe7+nCg3+B9bKRjKGr8J7jTV5BoiVLar2faMRr
D9VuRfpo9Wly7YFOQBUFlk1dPq5GnJZ6PXjW43CeGfeNwekvnBLPHb8YPgLZdhjQ
Ni2ISYbpEVJ6wn8V6ZdArSRiOx6f/6RLDOPOndcRr246m4TqDOvY+E3PpcOTZj7X
ziMNU2HBz1ixZaiBX6rhHbDwMda7w7Y1Tqnhge21swdNOWb2NE6qFsRmgrpWBG3L
qiiCChxS+xt5t0x4YqF1Se15Z4cdiyP9DASTVNvCL7LZRV/7I9OajNPHeYdnK9fM
XffsPBqSxxolv0ZGmT76kRZUI5Vd/codFWY2RXpfbce3I0ZATMm/Q/usDgkjbOYS
Dqal3SSLSpJ0841WWFkEIR2kqQ3BbBHr991ouicBsBBZgM3RZGkmBljd2K/XeJkn
H86YXVR/J4Ot9m49KdDgohniAAcIwLOyethPkNt3bXa8DbnJ1VKzpLskQ4kTQVat
RRZS6psUkx+kxv7aE3l0qJI2hTzlCii0d3YpmecQtg5gWv+KelasNCCN8Nmm4CXf
U8HZRB0bu2DByXY+EdtprKPlC7We1Mr7nUSwNKWpaipCxycT8ghxH470jGOKeRgv
AZZDOMlDZ0X2TbIRMOt61JezozJwhxIdOrzHdM0cMq4H4urNh759JeypMARC2y3g
QCY9zsmsiGVmyv+yM0gY9LUuxCFCey5efBiCf7Y3/MdRkSmQPPllu2ZVVqCheuab
6EG5WMm69WK46JPdwDnUeZbWm8rWU8M8EEbEron84r7GuuYAy2pDL+6kIaH5ZXvf
r6P3tqkMBozRkQ0Ax7HGAqoabNrPviDGpdGJQZU6Y44EXG7j1ENi+mEVXQVlqnKq
6IQrPTu/AWYnDppqlbLTNZYqRnDfqJADG3tw2eEgMc8TK4o8kyvDaGDaj+h/sLwg
plHjaxsYLhFfRM9bprSb4yoLAWI36/Nt/z1qCC24pg6AaZ7B5jJNzH9sCSLdxYfc
+3gwIs4stk8kWQGXIIJXReMad49TUNq6xOIPfbvl24VBSwNi7chRmaHwBgQyk+4H
d1PD+hFXbZf7RVu7bvVz+LKDfKXBkKlPDFsb1jMnoHigrsC1xz0YWqbT3DaRaCdd
nwJclBFyd04pvZMBbAxM3fm7N+oCN6zdXkGFlWX14sOIK6zRVpQTTNHT/t67Zkxo
Tak515Ak/LdGsGlR4PdkoO1e2wJ2tegm+XLuQ+k2ktIR9Mk3gZcpOYT9/HBpUKx/
jQFHvGWlnw636qj4BOcVF4KI9iXcrlzuKWjDkTEnL+99WIMzcsTBxGdr1kCgTUgS
nh2qGcVQJ3f23lgaWcY9C+pptB8nuahc03ZaooQH0nFR9Ly0/cLqBv2Fi9YeY7jc
YEvq/tP2YHtc0Lwygkx/qpdqiXJfIuQIUMFGe/MmvucIfZqWgF6CXUhDXUXkFDid
EbxbXGi/hiIdOKALlRe2jA68I5fDezkgweV1uF2LdDRXWjJOOV00xLLT16yWM3lU
jGYcS0Id/vTan1aMkFLGwm7LCEU6f9UwtB6AHqRHQU4vXNxvI+Mj5ojPVulz+yMF
ak3/VyTnEU+nuPV6kvN1Za4TdnoVsjs8DwlDvvqXpzENMyA3vr5tnTKYtYrfD6Av
1If7EjsfNJ1QqFbkJzAgnVeiG/8BWSdgWQdM75W8wGrkRTxFFiVhMjQWNJzLHl6e
cfZXQ9kbW8BKGjmkYJvot/uSvq7DUvUjZjvPeaBhAZoTv0KtCM5+nUKxk5VXWVjY
zdtitA+cDpjbLAAoFxtOUV4xlzMd21HzIBBZO+9eXrC9CHWufk8kZNjhoxiJfW9V
cRq5Ir+jVvW6UQBZDB6fUcpeQ9Mk54GYNGp6xMhFKnGpfHBnPuOXcg46uP4/FKkR
gvGMOo53hVN5jtaqRUz5oBLkYL8ZGYU5oWM7B5o5FbWEIgkK9IDQeRMRxSKbhGzG
G9VRr6AqaNdhZAe5SJXcmR3WusBXJeo8ikTGMCYYAf3Z8NuQvo3e2zvdy5mkkU6I
SUZxuMKykSGjw9yYBPi9HfN2rTWcyFeEMymGsoAmJH1ymJFSc2mekrDtnyViBuxF
8tW8wCpIlzNJxTIzabyxM3BBBK+DpMaPUp6MRpgpF6uB/qzZIeZoEl1vjFxAZQtY
9yOQShv9jupZlFWde0dPExh2d/VBlEEGhDERnI6fygPH3HFpOZY5PMrYLS0iFjx1
HATtCNn16no2k87srJLEChEv/xLu3pl26MZIRR166rN8x6a+s8pa+lpM3jvGYG99
ZksbZzuhsrfp7U2FA7GJLHK6qZ5WcLRVVEe+tAvwW6shAzo85yhduDFM+eKJyHDZ
zdO4j5xEX5uldsRF2EJCanjSKDFQYQmwkLwfAR3DPFe6OQob3afV94aFSMTTeIoS
daBQo9K2D32wPPurumZyjrhCraNmk9Bsjxog/vjpWAEwrgh2TZmUASoSc/uZpYNY
oTiTBpFvaVoYDTlyPxmwwo2ZIEzOmCoRGnvdy3Pjkcff8YO3lE9I2P5pqDE1tjrl
l1UFXJT1A6H/IoCvtpwNnkbgR2tDoJtnDz7AgRNaOzxgrNRzOvT1BossFJiTy14i
mlcUqSSoav4Ik0MAdI/WC1tXoiyz92pZZ9RwePovjYPkRt0sZsq+AHPuOFRr/MAa
C5cMvmV+/m2eQFHfGrHKPlzFazrAfu09Z8YnQCIbNduzdPAN6zpXwXxB4Q05yhjo
hdgcc6w4ziylpBAGS0jUx4noE6RbgzFqQycYp2U56ydt4FV9tEk846VVyTSMPdV6
1tRdSE0arc7nDTcwSvPwZKa6hrpJE07Q/u8y9z3DsqxPb1sxlqO8qrpfmEYIDNGs
F4lVyqXInq9zmYU2ldMOe2p5GiPHfH2NRz+SSDvuntMBSbJ6GN79Ye0FKuwnLFbb
zFRf+Mq31RnC3L4MoyfecU12AQzVageef2OQznOrl3RHXU+Q1yLNvAFNGKai2Rs9
Wxx8ywbNGjDJYjewSx1/eDCmxT/J9vzZ6b9B5S0Lk85Wa8urwFH3/9gdJWo9/gqQ
6rsv1IOMGs4pJVrviqf/YMw8LOr0ShiurS3vJj8+PlBGjUsyWESl7aVzeSWEdoa6
GB9mhM7iHxZ2xfQo1uJ2N93NgBEtfpXWIqnEzzGORw6uBWwjH3/IyXIcd7cHq6Hf
9VFCiwfm/mxZxir3T0r/db2bHnztL8tRvvY1B765MK8wjb42tUrQ/egu5w5SA7Ad
cZN/bgaoqEd2Sd4KuGhWzZiUTqSmQVeNA9wemJbCHu7/uIkYvOt3RcZKoZ/2D916
HKIrlWuxnBPeAWP9o4/gUSLCaI1JLlXnJ6KvAqo+m76mQyGyp7XVj5ZF9Xg0KIrC
ZuaCwSFfwr7/rH49Dmi2oDkMsgTN9eaqCAAUbPo+mnsff7E9B/cLmtA20f7yWP1n
7eGY1vyTwDRszkl/c8rXWqyVDNch4bosHpT4xjGt/YrCC51UGaiM05IYX9ZKMgjl
XFwQlnVQGs2Rksqi/ksrm+KalkiQY02yjTEjXsSVXG36KiFGDjeC0g8ZdK/4LhRE
3yqyVNEU9+UqoFCAuEUlIKkgBJS8UmWkGranfFKnQTjmgva8LdJU2oMJ1Sy+prVw
1+ITXUwWenvAoF9C1qQ8yiwAxpOmsyju2QdB8/FTz5dx+2WU9MJ1fL94g1xfGKpk
ly4GzhlH14GHVjQqHNlx+XXnscOQF2jVjpPBeF91M2fd3M39nuuTK6/X3+h4zRR+
+rF2qeUEmYDENzqqxhT1O3Nqd9zTSUlOGm0odVkcDMOBfwpsNuhEmt9hQb/qkzO5
7hsdmrPKOMGnsbkDccPtLAIypt1TXWsbg73Am1dbMt0/GM8G+b/iCdwBj9TnxGuF
bZqGnE3BJFdmFeYsRHHDNf99aE2j8NCmjPlQltlwweQdjbeDoBmgw7BlkCZcP80C
Tw5tTyBQ/3Y2y6c7Sd9vUs0w8HVVpE6rmbfOZiXpRMsp6Mdne6o/FcinfdicbRRM
a5MmlXrbAMp5M8/cAYklLkhSEL1qagx3nxhBVoZVO5Eztw45NSLMMIyCjNLC4IoM
tH8f61gzhk6GBAhsFSYWcqUNgnWRtALjQu9KwS2IrgAlKVR6mMhQmOCVjw7d0dD8
EG0fo41g5iP98K/1VrTJHup/nJIdLrCkhfiv7RnDFps33kj9rMr+q13f6kiKy+SG
U97DZOY84UdT+SkqFgK1m/9xNJm8gougOfODcALvomsjy/vNH0cAPu5gBDwQu6eT
thn9S9FMbV/66PAoxR8/9Aik0EZPB2j3P4TFGqa87OvKzLMtRZxz8NGX6y1zdIAB
9BBH9XicjMHflyLHeYJ7wAy93dbiDwa5GMCt5c05f+y9f1oFoYrvaA+557TGN5sj
88r22BmvZ4OXv6TceSrtrf9NObuLzfLzUUU7XRZ1m9eGs+V+sbrpAEk1dTy+sekr
0gHEJ8kxr5qD/fj9Ikg+vMr3wzA8JDwwlfwwCCmZMP+Y2ilElm61HeUdd0kneYgR
6gLT5yhAdzAVx9PYQJlfYzC5h7/4jChvUZ6yncw0ybi6r1oTljol8XS9f6Ivu5MD
1sXGLqUVJfBveykhzWbaIw4Toy9kjgccRja8L/vbKrPBU2xkrnM1zEjUwkPXENbL
IXad2lAxPy1kEeqFO6CiaDNnlLC4yqIxW46ZHuyYsqFUXeAxL4wqZjCR5tqv2Iod
DtKQTfifknoPkfAFOp5cK2dve6dkDgmsovqmLb+PrmLaVd2G+S7rd51QkMy2pb5m
k1ZLmHwUFS6y7Di7csReBn4kOWI0h+SD6z3zQ9Pa5uFzocV3fKWaQYS8k7H2AbRL
h7ul6YDxS0fIsZSEmpTiv5xK/Dx48hsaSWidP6znKKD7++Zrs1sX9u0mO8GRvpYd
9lD8IACEQ+MVwBxgIdETnT//IqPh/hSnuEIAol2HcUAK9HZbVwCCCYLEqig3X5rx
3QHlXsSMBDOB8Ge/AlPiXxSUVcCNYM+aa/ydGfmJqJvoxdxKq2gT/ttVux6IeJKP
XAUaYEFiltBJWPFCNmC4pBbLCN4gK7DByG8DbcNtercb3LWEKdJoFIr++LhVKdOk
6/GAK2Gt71U5nX73eha4BaTlkWECov/rXM5vUP7biH8R0TJGKSwhhshpRuyEBiUA
nP4EyTKPRWdzdVtGC5fXyREKTwsfX/liYV5wlPKI7SvphwoINxzaHbNtFaenuHZH
R+8OCDjc2DN/S3L+hnMdGQdDntxNI+nC177EXAuxDP9UmLr9DRJwsHti5iIqdDb8
sDVie7k/GZgrfgPm/oyi42PaVdOXqwRd6ei4JJfJrVpSHPw3E6/Q6u96BgA1Gm7d
rGgXYvsHOVpZHwVgwH4v1Vp6GPiLjm4JGbeiAs+ygoqNb82ZB/8zp/bUp4Tvy5mr
seFn2A5lYQ1Z7k41+4xFTUspYDL/ZYOYZudl6SP7A+D/ct63ANglWhqHOs8HDaVh
qconxYnL//Pf5Ov4Gznc4sPvGJfH0LLaakri/7K7GnCa5T03GFT7awF0WY1T5JoI
hwa/fMCjB8p+gael7UPbPV15SuZWOTnecmUontgHsxjsTvlysCHJAsuLov8uE9hx
Qnid+8XMtxqGyNa7679J/j7/pJ8K4FYWAml59yGTZZRsFWG4YCQKzAe4tBd8C3up
eCu7WreNoR9zA/9b9gfFdqV/GRsakYZ1Cs2k0tBkK6cezDWYZhSVYKhg1vEA436a
s7Iv8IGlGTINQaPZ6Qqk8fgUM4432/nNcSNhKP/zSB2X0UgZzY07BySb6UTqULxL
06bvr6yQRor6sevDEk8yYUUcvG1AMs/FiFOsHnulOgiYBD3FY+LRmLBFOcv4aCCB
TsNBNJJA/3ppQE4v7YSv4l3/x8NIzfmE6VWnquMz4X7B8JBFHy8AQ1/58M0QbFR/
zvCrGL2TEyGb9/0XjtZlcd0DVrHVl9KroQX3uIpfx0DP0yNec8mFFhU8o6Yd7vJE
BzaUuUu4xcBEuiFlLmCa4o2WUFQLmr53rn/8Iyzd96nTDZQvK8SRAs0p0El9nVhO
Iq1BuWPIG6u4WerWvHyYIUo7t07YvZdGwKmpQdKQ0CkQiE7hBjdWHKtHSdxcfGr6
xY/b2m5L+K5Mf9xu8x7HGFttqADAaOcHpuvpWW+IaFEx/e0bUTBvzfXzwfTTt2Nz
EBsGUJn805H3gf4QIfwEPp5N+42i2yH/DrisFSJZV5h/r2biplltlabC24VbnfF9
FN4DjGud9eOsePEGWSo+7bbrBPZQrYIR1HQpm8axnW8D/xLLWnDwfSnwkPysiMCY
LHfP15fHS2fKC+bNcvvYV0cqdblH2Jauo+m5rlB6cUgDTLQd/w/3rVctPW4uKAby
YEX0QmqX9rnyx/V3BuKNwgRtRVuNbZaYCZaCfXyAg1Ro8rPwxPeExZ85hZ5T+ZFO
Sztv94OcO8QeDloKPAwmTo0c9T/Gwn8vz1Tr5T0a1R2Di6E5uuwh0ZoEq4loaHTV
+dIUCXH49CB9rFO6Sv/cBSiR+iF2iLxtagoOlbwSwMcBxbMG6xpeVonHyLwaDO7R
/alAKUMUIU58gJbystaILCHm6SlE8Nvy3YEL0Vv5K1FxcMxjQtreliqhIyONLNPk
jtpIpeXFf08zmVB/U+b+p87dcQATq3yGc2nfSBG48o1Chr8/SSAxLwVj/a6arHtT
DWESFX4ZiqwBcGyrt1+fvnvPXu/rgIpU+p1TeNHWqTPKQkJ4OmaTK/Ybo9MvRHwC
eFhaBBe+KlSoZ+OnxGU33HDaMNJhcVTw1TK023KoS1eA5jLfbHiI4E+0x8awXVGF
0nzg1o4enPOW6vu0h/0JXA7FMwRI2UK56pkOm9V9DXwwERC4M0egHFkjWd8moLQk
DcQSsezdh/SKT3y5Piv1OMaUqIQFKjTNL6TFxweB20B7oxx9RkVVdwcYbSOxY+p7
3Jg8igpWBQDPWFqQyslHZkDzKmgATVdMxYCgnDpfhSyl9XrWS35KC+/kjf3ls7zf
moTUkwtqDEKsq6jXiwjCZQkrF2qX8EWh70xf5uAHtISEoCfFAkNOTnbDGPP/DPCh
iKRIkEG+zj9qFPlqxZy4xOAD2eOD8+L0YlriRTefLKMehlK24tMyWLPR9/HW0Odh
n2UrGNwlyL7+36ezx4+KYn+Bn6FGe9lXM/2VMHWpjZeEKW+Zigsxgwi81maG49VT
rFnJLwsXX087hvKgrBkXwPOB7rbWi05tWPmQNtFJDxlyZA+MCMRMO/wedR5W7wqr
zU+BZUBN0kLSd2FYGrVSJw1J7JZIWSz0LYjOxw3FZbzp/RPhfYA+jjtJQ1YCyQ4e
21cbcuAZ+PYWe61qbR/Xk+6JWhNhJ5JToC34QlGrmI+fQzVLTjLOCCedgwdfqoWB
MxeZgJGrnat7vYGSa7kd72N/bHSRoBbhS0AibVE3y1u4SxX2olcJly5R/fJYfdX6
4MY8NGVHSQUMzCNpT8vi03PIhDC5rCx5VyE0gOkQVACL6rpB9CeL/pnvCjSimKUd
bSyTNzueVaOzbKLwifJ72P9keq3g1HKUibBO6HCXK8QxB0aM7vewJK+/UMRikSMi
9L4xSVvcUOjP0WoxalQDieidCgpMHtvt3P9CHDHVkjQzkMK6rmq/ASjnqvnvGQcP
EDeuq7n68V8Y/Zk8lpHb6Rxlktn0c0MKwZj4cEw+z0UFqN4V0ns4MmnSmaGszcm3
yEvG6/CAw6LdAzSnMjAJmnFgYV/Ek3ZJEqdPfpqOhOeZBRgm/Lis1xna8v3V+sUE
GFCe1QKlo8Z7R/r1ZNw6F3SlwT/YTzq7LImInwdjq9sxoDysoJnpWjrR4yBgFGU3
UnhtQxnAQg2kn3DDtbyZUHJFYqqoa84cStrsiARVmzLcv8jLkvCMQQKFhBfn9BJm
IzyPvyosDgkUEsohmN58JBv2h3XQDBX2DvQSMFj7Ayuuw9HPL8hHXgdUCZLKf5W6
tH/W8gjFTMS2/GnFlf1fnQDz4E2RyHwndkCUNI8CboQVQr2ndbmIEstzWdHD+iHj
d3aVcucwc7lO78KtduU09YNLoEJrUfWX0Z+bx0JWGG6mAwFLHSnzaTLO0BXRLO0A
O7Cz+b+elWe7+vXrxFkH47f+OlKnuL5JOFMmbhBpfqgkL2zICi+Ut+42ukrYmGHP
s9csGp1QlN9Dgvu6RwrNYq+xRWZIcMa4NIC5sUJMogwNHW8p9mCjuzO6sUkgdbKN
CG03XXBmm44xJjagp9o+jfvP4+/QZIs65PB9MRoY9+v75dzaOoeitdSkNpiqc7pp
le+CkGkoa3kPQGhktQPBPm3ju3+UtbBZJIlq1+7cWbuAaNaH23Rq9r0Vdr3x8P+P
C4x5FTaan31LOp2w05Sl2mI6WGEQ3UNtQLeZYlKTGSdmTLwcFPrhHyC9wDfXh9h8
wzbJkIrfj3XKlFKl2fD5pvOEMcxJ8JGL3VZDry0sKViXIlmn5bDJEf872eiIJI6t
49oDO0z+Yt/FEyEdgDxIy7fMtYhFYJiJa2peCWgMT4L2Lr2wNoXXRbAGZmwC330+
3SvPmwVlddugTpq+IWymQNevm7eBzfDHqCaxOExktL+Vo89hxcHQBwdAO8WehDYw
xqijdaEpM8hDqS4uCJ2fdUcWCcYmIt0Hqmela0qer1rnQiM8MlcdVv1FGKxZs0sP
Armyzs1VbRll4fuIZdLlpx1hH/drqMwo3PJKJNaAVWqD4JSbg7Nw1KGTmgI9HXjz
nioVCLmRgVNN3ha8qHegNwqm7+oKD4dCWun34jngPHU1ivJKPVshm6YoS/MRqI+1
57fU9j62Ljn9euaBj3Y6SPleQgj22nqkEHzZgKov7CWlMdZrI57ZyUNylcSZjquD
9+zYwR9aZyqWMZ722kUhWCxrLV6EdQpzDLJHCwv6zxTU8wY37IfPZXvExyfMESki
IDD30CDj8FH1zCJ6IlM/2DUDqKlNwMs2xoSOFjhwDP8V1sLazriKMvD+/q665vmo
yO352TbrlQnnFMwYUhUUZhOvleYF678p6Ht1+U4EJV2pXpSkvdDQ5WHh3c0G3V0F
tnNaxEJZlOJx49KSYLDZzkUDeHQNqQdjY45XV19eSwk9Q14xEJ1NKm7u7O81ZSHy
NFDiMHmDxMdaYR/mdHP9ainD3DsfT0sOckRGQerHzjV7o4mqxxUaUh0e3Q6ExRDE
yuFZ0y1WVUnUAvng92SxsW3FzctBEMNmIlY0/ccGLkS3Q4W4k56nwa7A2/KpwUcg
rorPxNkYZ/o1oCFYu/tLcZ3dgRrFra9bV6BMQaZHPtFRdtkPX2T/gCU9AG5oTC26
pbJOKgeR9g3QlsiXehLyIax5Om1V51a9wUsMq50SlmWNMdUrmzhfIhfYPk0+Z2eZ
sMS4yQbSwhimiPXLGkegEPKU/PrErnQEsUz5l1QN2g3bUQ0rW80RBRDAKojxwe+v
riLdjEgqWjSYPZkf9Bxus+sOxc88NHR8g+CIDpBq5r4lZ8bMXhpIHAyUXw2tcYwb
5/tynbhspqj4fLCZDGpyUWNxL3LvYNrxdsmPoUmap3kwzMi56Ctz2BdWrMvQFvj1
3xp1PRU2CfmSSa3jNPbtq28ty16H8aBIecNIav4R5s5UTMnHx3jrCYULy71Nn5jz
/w37Pihdkp3K4QM6asQi0G/Uw1Gql1f1YEUJKT41du0qUB1PVtArhMwml0XeEWvm
uXFK1cTKfF3aDjmqx20SQ9VJGg6zjpFGhs0/nENn2TecqSkMHTHBoRdh9e4J7TRB
iv/EeQDwhE6gWUX2/k7TUmiW3E6DIYkEwAK/bJ9qZadbs/EIhe1nhvmVyDGH0Gb7
mGUZhuy/DIRKhvBPJR+3wrIAghcaDelrwhiKxmxwd3dJTzZtPdR+vIXzhEyOR5ff
ZVZSyOdAcQvhjhqd2wFp4Q0KxHcLh+4FyB2poN9M+ptbF/KQ8NPyTO1BqSEHoAU/
/AsfmCEkel+pFEX+ueij/JePCnSN1EL++5BGRFOaPjiHSZrOuXRbNTJUGIw9YQG4
Z53dMJrAtV9x44ReuTdo3mhSHJoj/OdORwGXn24xuxXpci0VyRa9S4BJQoCf2vEb
ySCrtQJCVCXHCj1jp4AQnx4Pdt5k4cAffxBiJJPZOkE6k5d0nt9fdSShuhd5c5/e
+3RigywbjaNCKf06P4iAC9q3wuBZI1ThErkcwU7xNbLSFOd2l1JNbiJOlPnOOp/9
Vm6jpXe0OnuFATOED68x+SDbtW2IZDmhrXOU+Si4CUSOgrgukhggcCtMQYOD0Rb6
vU+1I8ATtM12YRmtx1DILSqgOGbmtxX+2lJMWPWXLJWavvCA7f8o+sLSZRy0B864
eWnDcfKZJ9duSqwVzgRpPy6k96dhNYUO2J2i6XsWX03o1Q7T7OuWjoRhiNKlWdKZ
GPsYXAEMxNLqlfOexSSv77SvFXgC3g1jp9Cjmq2E/3EdTzBGFooNYPA/+x5qunQJ
q6zo/CwIbo0sPQxPhtNBvUbKnDDsvj+AQcOnACbHw5okDyXwkUEOH94O2fe8yekf
3cAHbsYSAAsRUdc9Jp+SKT1LmkHHwGFMOuKDLN4+SaUzuaEmTeFJGvCZn3g0k5Qi
X6ZqAKsUthfGcZfYbSP2TFPHfkXSmrdQVar/JL+2TZhx58zn6UEx+M+DVc/cCwBf
DnlBS5iP/10uW5GnwKxt6Az5hCKlXL4qID+/tkaG4z0BhL/pwji4T5o7IWkCwVeT
WVKXzxubYEulNyh1jRoScIr+PCBpGAeY+mPdEqwzfHgFR3mxfxzNe61DYLiDsS9C
706sjDO2pDLOU9JI8bUAmFMaZS0Y9m/0xV06s4jEX/uXUW8dCsPHm5kO7dTt+zeb
zeQvwlaAFFmwX1m8Y6OlWeHrXLwynSsgHjjQCF2z4OfkXeKF0SyijH4dB/B8FxwV
Npgubuh6+f3F2oQPfG5JC3BZPne9WrFdi8NhLIVL3x3ceU0kn3O3doZy0F2u5ibM
Cl7EShZI8Fglbdt31lZnqxSLb0nNKjAvfllqtLRiHk3v+1EZOdSvvlbxv5n1lh5N
JiMxwtv2/wXk6CcPeESyMZkrB1eKSnZWV8aR7gpW/Q4TjIPfFeA7gHgbFMskdtL+
EJ5EHvoZwUY0zVh9wWq92BvgOt9KoDph5LC5CWqceBhEA6uMnOF/ynWUq6Btq0Xj
lTFEb5RWQNvFZaSGGtckpPnK3zvlwYTSan4uyW5zjhuxUyZQeGCdt1pu54lT91gR
ge33LVCNDpj9mFE6KNiHqWSy1w2JAiJT/+1dEHPHDA4X4rrf7bKiWvy9ysFqlFaj
0OW9e9k7vIbt34FYhX8muybAvmNHXnfGosW+fOYz+7dtByKpYcX+ku0DphiumJhi
8RLH09DBxB+R+wmWO7rZNHGdBPrOJ/e99bQrc25xuXeZHjwjgorrLx0zqychsi2f
z/nyMFaK5MTzhimWBAgo75DYZUBQDy6IR5CeZv+G4T9R8ZejFLa2IflvdwEnECCk
oiwIGADPYnVZooLoQgJ8vnQXbu2mb66e35wZQmmZmMXgPwRHu5vKdhHep1GJ+lJV
KMvH0V6elhTdBpiBCFyjwBkkyInNMK3ttrxYryf4q3craJ9FRn9NPVzTNCpDa9go
+I8XaR9uM8H+Y2gDxHQAMqueWwBI+iSYWqlIKtF47ASj89Nn3uy6gxcY3pCYmmLw
5e124WqWDLJhkR9Tj10aobynqCOz6fd6/awXsy32Li+L7Ox5XWBp0fJLjiZlFQPB
kkeuF4xA8U1vl2JQCuJZnns5ARPgEW3iBIOtDO1x75es9Vc6TBZtmzvaoGVEiEda
ZJRW6jrg/lZ9792Dj4rcnv4YQz93VC1Dvja9K+Ud0nX/JYty4Ao0V1Vv4XUJCfTe
0O5yrhR1e3KvZF4svBWBhmw7FW7QzQWptdcgiWheeTGbbYBrxlaJlyLgNSauSGJh
6J47PhzHv2r2dkSco6+DU9V3/3azqlNoXFqJbwog4PxTkclUp/vvy4vy3g6n/RiE
qiJ+/0xzD1dtfVDj+YFGaIiUvmO+kSMNKwCOhJek0Y1VK4UnzNSSvHfoItTgn8Ab
ylnHRDkXGz46X/1K4E9cRbiGmynIKqqRQGJTbOQRSjuoXPwmxidKS7uiYil5Myaa
UW0TgOdlWGL//wYEuk3xuKZwq5XB0TdjlLEJK1bjHgkiepcZ9WXayjveIarSDxEa
7nj7v0UF7YIdzHp5h0pdHubbdCsnctg58BIYJiaompMiKnoGc5TMWIv//JX5aFRW
NStFsIVJDp4qS64U3QU1HceBq6Ha5ORPI4hMf0GQUludLnvpJrhovO7FNlPpgQdj
gjy6HzgFtxgD0xMIqmwpMEv0QraqSigmrnVu+vOPNy/B/r+CIPFe8bFIoYrdL1QR
Hx/JBInEXcna3e/loR8xCRDpP/zU6wuI25Ix4F8fBM0lMoVwcEtlfnL7sLcwnUns
3iK7WCiN0PEZpP8V+Kv6rTHsWRSeCJ+qNUiITOYmD99B5nkFQlkRmkOgccEx8a/d
0cRUngaWVc40loNchgIiIdH2xlSctpouaMHJbQT9pb0VTylyJ71zM1QaXrrWcb1O
4PlHTIWxExxpZqD3djbGt/x8Vt0Wbp597TJGPfaMGSuCTQ0VZmoknRSQuy2WPjQA
0jX3LDxLnO2fGyxNFt6ZuQPDDcIGkuGqh9qts8PdjrOKrs6AsWBYHQdgnfVg8wOT
FP7Yb3hdbDIeecVJEAzaF8R6z5QzNK8Eg0EMRXJIfXDGYTaWXyYOUWRd6sMa/InO
VygvitRer2VISKYD1sCWW2kjONOxudWDNyTGTV4IDrlJ0K7wcbZUT7Zb8MDCn2p7
NmVBzjwR1IQHz0wigYoGzUF97kNvVRIeu48P+On8sSiWuxxZ9p2AjS/aQvNiAcFg
8jXYtN5kh9Mmiflrdx5zgf0cGbuer3yLC5HUxao7fGxKWWFngwVcRBDbODJjyGIK
KWAoTvMH2vUjuJ1Drx5/0tDqpNhvL1P7PePbSq3Q5uZSmalLbrdrhkxFarNyivTB
mli9Q+4MtMq6kfxe0zjnCWe9zDUi5GswCmu/vUG9skF1FQH1Zlug8w9ByyH2LN2k
+/W9+MI90fpVAUrVcJZII+K3oMUpOpt+/5Jm6S755We4jFUyIG2/Cpg+yf/dBUKZ
l+CMzh4DOMW3bfFvUDRo8P8GYarNZ0Zxxk4W99yvjbUX6sGs5EB5ZKRmyusJ0Srd
gaYTJBeCY0+cYDGvtqwVBrUCyFwGIh5rB5CE+y4xfZ3UVM9Y9qKeIJOa8tgTTTuU
rE3+F7WozlP+/sPrktQM18rpN2bs6sK3KY9q+QgIk77XnRV9TzgNNlnZudVHeF27
v0o0CAMtNV+SttPa8Vbs6DBzT9ncx5ox57vEQaRfF10Dz3s4Zk8XkkdlfmtwjiPa
TGW/qXlDkN9D1hjl3zGURZ6ZEUZ5y4jLzsDSXZYOUMyh/+Bm/IjUPy28k5TbIKKB
FJuifZ0hoSD9s71aOxG85qDxo040JyO+wETgdwkC025edjK+axZgGsgM5LcmjCZa
xwsUQWxLJSJTVZv6/UbhCq3oOhp+xAnfHMAAprabYJ6YDjbeYcZWgmBCYYi+BGEz
3B8Fd1/YMWtJLdW8zNQO9q5zN40xuDw94FR33giJmSUw9NGFMzXy5KlNlTU7on8L
Tb6waSglPv0LRZpVvon684BrpHHTwp7Gv2dQeLPhfGfv+NSy6RnB0I7InpN1g/pY
Lvr5hpbDsKTXiRHTFCzCEVU8WZ0FBH44nGDXvooHHJ/o/s9AP0CtyYEnaMleI9mx
sP3hQd1+HAcrbypnTjUhrDh1XZ4SqqNcNsUulbAfKJSvRUUUWZ8KgqwoItLRoth1
XkyREJ+W/sUmLQiccgINIAVcRcc44YAGlKACQ0X7SGb1WCkZ2kMQs4qQIw8aXNVO
LFW2s71ctbnF+w13oO8kR9wVF7VLBnXtF84lM1rlAKIMNv6jBb6TGFX1h6ov1cyT
K/ioVzNzpfcDnSsYWYhQAsBrYYY0SSK6v3ccm+6UxF+mzu9Gx3OEcM2Gv4IyT6J8
xQM2/93/VhZa+uF4SPC6nYRAzG35QhADe8LN0amAliKbZYEG1H0blre84quD2NM/
j7rbN2Z8yoTQY2w1j8wNAOKEzoUeZOj2B3A9Sqgu9t0hKspKgY/DLv3XHXi0kUV4
LRuM60gklB1sXXP4aSCjJ4O60BzyZL7LBGytUY+n4XYaLk1zpfnS8yklwK4kNuKy
xuvCUXOptw8FK28o7OeAA7/YmmYAXqZgt0K+wW774jxI/+IAec9kmmqspXTZ8tlG
ULdIMqGFclAjpoJXZ6nvIViEcF3oaetBptQCAPsTOFpNuoznFcgiV4Rn1HCQKIer
epu9iohbfOLRflI6ZDEZLrA9sNeA7L5TnQm7555LjHT2KnORNKBcn9BGJ4IO3l+N
elcXKNUN9ihr/mvKXWj/RNgRg4dUjWaY7wm8KVyUquwg+nFyTaHIZEZ5Mb2GxFB9
3ECZuiJGUbIzejC2/wjXUdV+EeYsC2Uu6B8q0jihVJwgEcjmEjSAEI5k4jDfKaGm
mZurNtmuRX3sAIELYYAY3NFdB/Qi8jEKmGZyeBFTwUg8aJPNdCKvxwDDDY3Wbfvv
1D0TZOT9nhWYkgg+XAdOpOTgyDKpcTb0A/eGEC/94tRXmWdV/SY77V+cA7M+8n6W
idC/j23GOKX7Sf29tLa8LYeM7AYbnAkv517uOubPg+drOKqP1m3/Pe0tg20wdYdU
Lft3gsarWbHyz8QHw4v7D/Pbg88fEqDsvQH8mkHX4uUPyOO4+dQWPfKzovySzNtc
/qsxwBqSdK69YSNfe8foUuMOWXPpXurcXNvTk5qGdGhjowMwVfnORQtdYWWBSfCK
Lc55zXxyv25J+U3/LO/3IrXxMQ39KtLQiys9EiYjBiph9pEIjBQ/gx5PVI0GMTEN
KCl3QKQ8oKpvjCk9Poe3ZM92NGqPF/GAxXzmiArW+Dktn62/M/HHd8xjCxgc7TiV
2/e8hRSbtPOkjUBb4PuUC8PXjHmEHWNTHy7WXZtTkviaKuzOHcuPCCwoLrWibFPi
lYofW4xcp0/kn1NutRPmyjeYknFIkanIqZ31mY+KEJVkaDM/IqoVj0oUmWTrKKV6
GJkUa+G4HcMDmOhhC48T/pjFnibANjveZCsvctgX7X5/53jB5a4xsfRpH6xPoPiF
6CZfe3c9O7VHc/plsVEXiYu9V7T1Cu26Yjh15FtJNEQ92FlbfIRoUmuDOUMmXLwA
thffd9nk0QuWbcfXiH3XmKSp6x5D55Q+PDc8LofQisdvqHhJ6JynzShzkNf8OH5c
K7ZOCUgSF6Mb4ppmoPQRLvcbzCzInw3C6YFOSxrmla554ruEadSEdU/n/o9FIlpT
ihom1fqNpkcLp9S3z0bGMpfaRzQQufCWyvn4gFxk5GZHbt44gEqWZI5QcYVTBjYS
4khB8TldPoWpRdubFXPMa6copxQp+ntBTLIx9AQBOITcqrhgmRPHTi13g0iLYJTx
7pvS3iEYtEFDuj1WouHhXGUQRno4P7BJA3R/nF6ehQ62tHYcXRCIGjxUkpUD+Lu8
mtuzEAHJSBQNOEIupyCAP6+m9gR3cRbyNBmcEXE/H4lCcIRoqtYYoHH6YL44uMiX
/2GbZ+4MyE7YaTuhX7E/GNoj0yJ2TGMFN57ewZR1sGFcDW/MLPBJ2oLUnKO+Yb0l
hNCn/peuMucAJK/CgX20iFGFI30NRcVLZQ0+el3e2qwRmbhW8i77/HZqsxRtAv5E
yZQPLvh1KHOBBT2OogKDbSV62tXvvA6AOln4YDx1O/EFG8PUHdLxFWwLVZ82B7GW
ZjV+rmdE311P0zTnRelkJzTm9giuDtFFBZEL0EUQ95unhzZvzHKdTf0ZzUekRjec
wF6j9XtAvjcFncGSCjvIL3uz4Z2iKFWMIszXqLXR4PSxUN6nlQwGxAjITrn/ZlVv
VMETm7yPazgIBDFF5iPyc0n/qFxZe8TxtDgUtglgW0dxNPaZZG3sahc6R016slW+
4GM9XIYg7Rn8ln3aeRJctYwn04PQcJ+Oz7zJTaXhIWNclWgjHsmbtqa4axye8fqd
SjDJxgN+BI9z/YgspWi+t3QLmsv416JKXTp00tnq/PG08SrDr6E5WMlf0zJxx5mf
3Gqbo/94V9GOKma1x7raVRh5id5kCBjzRvG20+1vdywuHEWZIvUHZZaWsnY8o9XH
0glmbesVrGGWvC5RXFjGMmTo6oHmHoutvnUl4bs99G3WCWDPp5Bb9IwVI3wL7Odg
FdcyqSYvnMJdvI9Fzbpc6uABBBVoHNLYCHvbxJmPHjAtvtpfx7D7+YFgmFLV+gBZ
AGYLZ81wSNE2FFPdRVbefJw2KuBUUu0HJyDtHswYAkvxXoDoQeSg/IQJwnENfLPb
NKHvcwFBRHfQohBTUFGxUPI0nYmML/KkWGVtVZbyyhs4BfaZXqTu0/aOF+UrQv+z
ilPROtKHJvBaJT017zyZmkQ8v2LOYzqm5bgHB5fATSjJQET+Ht5F0c3vbjgWVckS
DYlePChb2PLNMslaUiUc/SB6WMXOgUajsCcQYqqXDNVPi3WZVE4DLLP8R22C5KPv
aB1MX1nFDWIiDGQTDkkdIcqoWpKd4yMv+4DY1FAMjT0N+GNxz35gWQwX0aUuRYGg
pXwUBOxg7dDxXFH9psdmn5SDZuKRe0wg0QVbKG94PSBtK7AwXI3OUfdHbq6aKoS6
Fmc4jLED3JpSoBqzapxIoIxmw2Pq7Jop9LUh1lLTPlxdzBpDDV7xj7Ek9n7iiA/V
wm/l2W+6haCBdo/WW6wBFKyk10WdT43YXJ4w234RAollpSGYewdOM0FQ4FLwWSHo
VCYCyvPw2zwhIDoLGhmFxmjRuaVTFlLMKrz8GfQFFJX9pIREXvkm77o7x1Xa5hX7
e8MOawcyAosnylWtHnMDVYPYXTswn9yK3qvyyd5JOW/1VXEm8FuLUPopVbk8UO/J
Ez9xu31KU1w4iPoUDsg1bP63/aFRL0BQoiWRB40eelf/BoRdH13vKVztlbHk0iIj
j4cSAyKkleprdSdrTwZyo0DeUDHtJla9k0ZUwk0ApD4YP/adgBokFH5TTO7u+L1T
UhKWF71TRfEbNMk59DiybYHvPA2m7L//X2xwOLWWZ9DnkdV3PpTduGDHJ+EnjXyG
q9wxG9MvX9rR8Ub/l7OJEjkSByl5rP8tp+ny1m51F34aYeDezlGU/v8EfDxo7RGB
c8fsiGjOgIh1foxVgW162PQ/QCJddtnLMmqRhL9kjDTn8cm83lbyvYOM9N0lA6zv
CVhwys692uMw6WO3rtCo20BefZ0QXe9AE33o0MAcMsiNBLBQUELmAZFuO5SVLXd+
hIJQBHxyWWQxe8lOg9l63pObvcxwiAgWVibSFhQaSxerv/2zZvTQdGX3tKdVsKSr
k7llUepwcj4OCpVZWlPbSAjvGYtpqdCJgRCM/CLjvarCKGrUjvGvzauYiJL6pV0N
Ixwa0Khi66QK0Y6oXhzsA6dTHNC/YX8IyMenhCDOzqwkOqH1RWWFcxZXyVd137QS
ZwpBv+wyBmeoUqkoSrKjhUtIIPNnuk2N+E9CkDS4Tp36PWQa8BD2J2Tz6dncVtR7
5OrqtTOCGXtrrFCApsr25vAQXTvQDe1JJ2gPmJFjp8Cv7V3nXFrtEKplmThvTz7v
B1OL0usD7WrF+7JbrmdsZGc88cqQlkdXw5JMviIpKdCXIAO5V+xsQSZkgMIr93AO
FnjNe+L1n099Eftg8Kmh40H28xzABlsrXh5eHMoK5yVLO8R8762f21TFKyJrbejT
sGCmFr9mU7gh7qhYJ8/DP5YCb7alyccjPKl2Gatwzp5sTEK2q6jlRFnZy1tb4QbP
iho1bAwpYoJcHs5fqy6H2R/WsLz1hX+LG6MmjedSLE4cb+k/KitLWCW6RCBKaq/2
iq6prQWYUzX6fxnl9oQLC4GJbj+zh9XvDq8Tab4dk+IQ5ryMca50HSypQF5StDxU
GvPAVSBz7f++FO3vOG4dimpCL5n9xjD4Xy5Nmc2AI2OFNQ1nXsbIcOx15RFyAb5g
uhrHxKSq9s1GTm8on4ZHhfAehz1IukzT7iwC6lqpSqxOdvhqOfPPUpwL5O8wZKRv
eTJUNjmvtKI6wK5vCEhSDeKi85nXiJScyNL7zNXRpowrzDPzU3ZfbDGDt/L5nHPj
9fVADDT/8p8k+GMSKPnIfmEy7ixZViYjyvfX5R4BLDBJxt/RcpooqlpiLb4EnK3l
aVyjL3sEgrkNGuYqLlnbWkK+fyfRAEdpr+vth0B3irftvxHsGJk7psO0nR2api9q
LPGtOzucGPXatJ7LEj0Qgp1HKagUVxWryQmWqkDtycdEuXExMxNvq+wvzVa0mDpb
KGpvS6xnOLcCqroN9jwUhYY+mf5mI3wZ0Ecu2shnWdKKJQ7DvYjFr7TcRdV4Xmzs
RlqWoGdr6JDv+8evDd7Of80Qq4aycPyUEGyQ3jlRd0NKQ2RN7k7EACHcxcmlGqHm
IREMMqv1nmhSiK9W52kAmF7XLpXQ28l9td/Tfesem3YyKbbYAkrxiM11vwC7Re/D
r+p0pbQdYl/O6xiuGx/HWW+MAH8K6WB2sFEIFBlcl8QJ8lm1OtlujtEoKyYQgPcJ
6+6UsQimdBp+/1PpTdgiIinWWaUWcRwe2X9cmkMeeme2legYr8Y9lXjLztHlzWSm
oitrXZ+d7pTbSuQDFtOr4lPxpbGYyYltPyVHGfMiXQld/TR1irdo8bfmhBCyAtLW
LE4xNfJ4bcfhgLAInNLgrSx0uY8MacQBs0yd7Vn9xIcapDBdM6eH6fxEIMe9AdXz
rIJNSM26EN8EnLSHtKmxGICdHUrtXSZJCjoGCeRIdLi9zaDAGWqSmk3kpfQWDnZk
MffnsyBPOXLh92ASbxV9ezcRDcqASptXhJpMQ9snWZDX7vaeLueTE5RNDyYMPAkI
hWX917umIxsdYSQ8LZz4olMXwhk871DJnBnY6hwQaDyKdM7on2esEcyx1IvLXHgC
wTmuS8cFeDFVZ1x3IEidAg/bnidG+xe0IyLg9Y5Tt+DSdGZ8mXcuJYgLcLGaMvwE
WVRHuWUiJX13/7UywVWaVRCYDXr3t1OjucWTRyIo2vqyL4Qe2eIKQb4NAmcKbQ/r
7ov5xBkl03NvUZNRHGElaFmlK1mFroDxeJQcuRNDqGez5irVBXAFgPS77SA597aE
92xlDQgd2k/kprb8+QrPytYC/Y8atgfY/0eOT/HJ3ACmfuUKs7FdRK8U4Qi/oVgr
xbY4yw9fp5I25d/jfZCPapv5noU0+z1Oz4O9flWBP9Wd7Hq37hMtDPnpZsndeoYX
nXSNTWvB1iJQJ+B1yhljEEXsnBL3sO6TR9vNDmhIpv62QcB8oXjxr4bmUj1IWBYD
I9NmSwXWB88B/7WtIu4zGofANEeMqIFXcHhYmR6D6FP3yv7ATywneJiHmU+V4M0F
JpNbl9khVk+f68X7b+7XBMEsQ0aBRbwHmoCUPDK1s2dxak8edVHk0ano10WzRz7A
22UhlvU5vhHQL4bJoHd5zEdWnluqUT0urnv4B2Fk+vyVak/+fFGQQewxUg3vFLf8
4dva47yUqGYue/PJY1U3O9NG/qmWjE1wn1Y4IHEh2nRuz1cx7Fv2TkNGj1JUbph8
/7VWF1iTjoSJfkun6xhNi3st1y82GIu/TuiqKo1fVurq03p++FXKyWONtPZlekdH
xnX6JBUP6XnJSMNSbkdkiT9jcYAHWohNuDY1Dm4w4OQzgofsB3sxLPLUvkp3+BNR
ujjHsBqr2SG25EXSyCWcibqHzSsc2E1DA+oowZmslTUT+jojCLL7+0PUhGBZK4Aj
6KNhgDs2LhPxaDlVhidGx3a9cW6XehKhv51sFsGuNddChxKkQB+/x3nzFquGCHWW
0OdH1jsG2JtZlDtYSN6opeGaYUuZjU1FEZXelNzveua7hi8zGtdR2Wbe74Wl9526
vW5ozmBmqJ3CscEJJThNvLdcL9OKBezZ2UIwNpfLkLws28pgkNwpkPWFwLo4GQ1J
NHXfxX/iALFo+iRNuQP+O4QVvE+BxHd6ciluRbcFwQweCNIaU4fwNkWke5dWxlbF
nlgiUYPOPpRY9xOw8IOlevJVAYXkhflxiExHTYKfKY+onEUadcaUps0QFFY1fPJq
/cVqFmnEGY0bHciOyFjBxEiBvr153Tjx3izFN4eR3szm8ip2s+miows7/wOMvRXI
TWOLwOI3CsyUOfHHyRkncvvhRSxgE3r2c2tjgp/GHHW+1JnxjA3oImjdQO0BwTZ+
rnBk7fyPCr5liZ/2xAYRQWkeA6jtVDeKO3/E3Jgl0dlRI3vGZ+Rttgdu/AqqaDQA
oiQAvZkYyUEsUPJI/7/Y9bi+GfidwHOKixWewa1kluYZJ3bWlwP/aWgqI7jvc1C3
nxhxzGkWd8YYesA1Ssb7n1LJEN8oTECXRbB5xL3uhIOWGXAQWzIlNiSTL++hw35E
vYC3bqi/6m3mk/XXfJuOneLlr6vWRKunKASi1XKBNRMKh/5X5KujnjJ+uwwn2DDP
cBu/Sh95nlTx8UrPmkEywM0RAWThuHIs+jE10y2DAsIN9fnpPNeyHUcX2a3l5hIE
Gkp6tx38BG/uI7MZ23K9xv2OwZUBhRYHVEmKDMwtSy0K8xr41sqhfIkr5LbFGhMM
vzkSl3stn6eSaPg5WPN3dBIVMr7t12P4V15ZV7vWEm8+QbCtj4zvAcY8YZXKtrUQ
A9OxgbxQejjkh+r3C66AurMFEbNUyyJ8peiCicBa15nA/pfPhASFzJNG1vTYNjJM
xBXYhh5ZuLCXOkliDIcyt8sVU/U1kgNJgTf2RUoygAedXW2zePsgfAjl/6KIdOFz
ZawxO7/JzC9Ag4SRcBPqE5kRG1uNHNyXt4k/rbslnCx0wn+nTRK1XFU4XdYosbkw
NMdkCc3wgElobcs4ieUzBfR0g5WzRjiEdWVlAas4kJTSpfdv1h9u9B9AD6vJTa2M
gd/k1iDioqKQUn5NlcNybjo907/+7hhqqERak4Xl0sZ2cAdDWeU6F1IowqpJ80Ge
7AbO/lel5DMtz57HvfgUYlvewBpyLCbaVYjdS/ThSxAQ1bcGdjMV+8YAjtgM+3Kx
DbmnvBXZUSYTJfWfu+odLM2DS8cOAd0dIVm9VZ/ENnqBkDMr2nyv3JvifPinBvrm
gQvq6tSEKqywDBMe3izUBFbhMAFSih5emSwjQyOL86fDGp4X+CO64WcC/POAffj8
GIqfkRk3dCe+RP+lN4dHMgUVHcJ76EvoTto37NhNww6jEgxs7LBKO+r36z7y6pWT
OrHjen3kn5MtJP6YC55yuuIKm1H2+nyjZdRfy1KV5JwcbI7Q4DjRF9QIda3NDBmz
Ow6hnz9V6Gb74aqohr9SeVRBR3WF1cDIlWCc/92QGwspWtyW/YPgt906GN82GkJB
OJs52fvy+hdFampu16ViQnQZsa4hfUGlfnPdMaLFa2B+ICn67YFDRYFNb/V31xH7
7vuwYLlBkcRfdFyuSrOubJ2Sq0t2B5iQcZdImGQpG3AleqeDXKJ5lCy2Uunpu2rT
A06uuHS2x76uumColXFEQL04jgSFfjd0SlnqeNHQAxI9XG+GaBJwJJbjRPVpJFH9
ikkEeMyGxnQ5WAyluUKp8LZMrW7GdQRNdIXdZDuEawnH34nqA00iuaoCyYY2Bud7
fhZhdkUEL1Lumptn46e/UwVZTdtRYmT6QQ7WL0rtDonIjCi7ZLMClSTULg3cZjm7
wPfpucXIn3OsFOr4VhsC5qaywmNzl+cP0GXJGmpVX5vAF3LgWpLPQqA5/np5SVL8
r/8avf0KDbmeW8Rcjm9RQhih7dOSxsofBeb0/h8BvH69e4kPPsWRVDrSRYn6kvGf
IC1hgpY1pnmH6xbX5v5xDDaQL/aAfafSx+ZVD/NorAZMbFbjD1gqAwhrEWb/KM0U
RkiZpqyF3Min71I0ugdAn8r1VXosz2WVkT0HqgH2XYiS7igZM/++gbAM0GGuJMid
Ua28Q8BJZrKJZRWmQWOc83xw+R/ln9iP8FBjvX12xEp8FL67QaPlCwWpz4zTg3hA
fQPByri3uJWCVPR9d7Fygp27E0W8UhKalt8D7X8v82gwqX+lFGEOmWGA9ONZq0Tn
8RoPoUKn0N+IoKZpXOKMG0lhy/12oUw1MH3Aukqi8SlC8YKZbjVQjvI7WhArKaW2
hnrRo+exI2WqhTopVg/BQddz7GZLAM4V8Lni+jPm4ZifGpsVwuVCjjxiCuNpi3yh
tvS9QxnXZv90CuCUWFT8mNRz5rL9SpWvXy9VFTQeSviCcloKnwYcx0DgvsMDQ/sT
Ub2o7xISTPOrflYywGH9Bu2Fp06x+Ja1fq7lW3M+tFPbyrxGXABRso7Xu6+bMuh7
5RUU/4ioFyEOVrOa+yTB7PgtBxfh4wI13qYJ/LyHZ43eUgEFfg/4SHEdpcwhU1p7
t2N1gm9hNpBm4f7Vvkht5wasz2RWHz2KYsSyxsyhkWWaQgjha+DDCTxI/HWKxlgo
MpXW3lyaNBn94gPo6V7rMWSO76CRImWTYyVU1Ju2YK4M9xlCyXDG3UnE9y2ZppSA
Che7NnwiZPY6mpLg0i/aEhxAUPxpBpUwAKPpZV9XJX240UaHtqv50y3Ym0+Q1bxn
F3J7YwDyYEGK2s3ZvGhq9M1JcCPw63HT/WgsV74SidMgzDiAxjN4yjItAQFZg7p/
eJzgaq1IfeZNsSbNmj9k/JktTAk+GiO92dMHwdEK80ePN3ZpQ2m4K/QZe/v1eFVN
AQ8sUZ05tFMkaM916b6DZqh0CPPgTpHN/poMu79nAfqufVojnEN59saTMdSnpWCI
U6bvm0vgmfIxrb0A/SCvoU7MNV0B9k6ac67fuFDlSQ79FBxi0PE7PyQ9fw/wyH54
VeVDlL58U+y4K6SXcOP3SejGGQuHwJ/9kF3T8mdGSzoyJ6WHx3vbWtmlbaOwDds7
BecRrmAsrsccrFerdaBDKajFZIrV9dto4zEuP6JFyYThVyqhzFpVutJ5tOy0vAr6
x771SQn2otyDXge6ipnk843s8Q7V0B2oUIt6/J3KsG7zRmnQSJyRXJN9u7NxNht2
9dBFsFhvAWsgu7KIpZKAK3isq4mfXnVP8RGGBaf4n8wY2fL+v6iFb6GZkrQaXxEU
GcpmNySndZQ4iQO6e2dLepUuib512Yk2Hk3ucxE5cJCF/50IWl6P0xGhjqvXDdil
xCtbeeg5MYb3VWp029yb3suB/67cW7mmHafaumD6KWB9OobZNBvlN8csWj6KhEsg
7yE7ZJ+5VKijdVdU4V4UU9sCNeEW3mdCStReP+cGlCOonNzPnTfkiQo3/mRNhkTW
MJ0nZS3wV7cBwgetJ1r6r49Tr7AUVmyuC5M8p1QC1WNo51IMMM19gFsJjVDeE34d
dmTESZ2l4xlX91YfhntnJ/+TLQiSyVcdKt2xw2pEvNbxt5Fyw6vxQUjV6bLqPnAk
B5TSFcqxYNovTlxNL9PPMQn/u0ZCqHl/62ocPULEHFaRqfK/u67HrKHEbaSKezCb
Klzby8Hlvmwms++jGThH6MLtLoqUY0fOFco0K46IXqjHaHrv/k5z7MXH7IqUTTwV
BGKlcROZWmAWu44RW0nXJjr78yVMQK+8jWoVIvzgS56jzN8awwhY6hTEmt52bA7d
v/OXkHetmzWcMntbFmgJoM2kkN+5BjeuyluGcV/1hweumNXdTwCzZyGRDHOIG3IH
mtcldtoyMmbm1q9yr0+c7v0GWki22nv5QrVXTrxMy4oL5UfeYxy6NTbWO6HCGQvT
rCwpT5D+HCLoN1ZdhUZu90Fjm22ZhMXNAjnSL/jinxUtGGn20BX52jLScbnlzVrE
0ARjpdL5DF4/IsAiiUJpeAkGGknVhMGHDq5cl9xC9tHFyHGFFEA9X+ruADDXcSTn
F/4eJKC7pJzUl5XbnZW1Dcn1UCbyZwaSnNyG9/l2V+MWWfJey82AAi61Hd4LErz9
22jTN/DOBVXcpW3jyREFn1Wa5jSKkq38XXeEUx2jSudPjvcL+D5Bbjrvz1PR6b+h
Q8wwWcHD0QSeYUJSbw9DFs/QqHKiEaYQNkcljHnN3+aytMcxJvqTfq3Hhz4Xp8U+
ERMBDwK3ex7+YWXC/jTp5oAMNchbLhLt9UbOsestROLPet1hIbDCxPF8LO76oTE4
Y/obqULMx1UYDglxQfQvTG+O5zign7L0fMq6Zv+BNoRGFaPfmJTCfTpD1bIg6R2+
Youadaa2sguPgptvFHmIGwYAbnIV9frf3bJf4hmB8egmTObnQQ82nr1x2bhht/ov
CHKJZnUZ/dIobqtui3wXNu1a9z8co/4N36yoyoUvMqcB9kJtKgqQg/sr5eb6U3qG
n9DbLNJ0MrfDPtxtyZsedr5pJFo+iYEnXoWWHl7ZC6HpxMbCg0i/oV9dMB3fW97j
vFwLIE/6wNAafgu5o0jrfdwxaNIRmLcFVQJuGshMlwtRH7LGgbW/tP7PVuEhhbUI
BGhbIhSdRXMfcD9QSmQDXPQMP+zMA7AwtNUakH5LZPc9qvMNOcsFP/MlGR6ZIPto
yD6TQ+cWDPyweAxVjI5la/NoG7l9xseyFNqI6vhsvz8rsRMybqfK205LSXI4gSpR
swsD05Im1RuqNfYBAD5Zdpbp/oEAJT5anFTE2cGMbqico8wyTiLBCtsqkIief0s6
Kkr2d02boPfxtcJGZHlemB9qWB1M89ECb84o7guGUcGlXRn5ZzLAyD5JWkl9Fmga
jRBbdgLWKHSkeYuIppfppfzS8kqH7UnYD9uIpoc699C8koN2893NQVWx3qk4ndjc
vDa/H1OZRtUfUyDYDaA3EUVL/3X89mvGBETqEkWrxv8TNQPHaB1T3Q0eO6HNllUC
vtAIPqhB7Un3ywZylfZKfX3UiPfGOpVpbuoU6oNnvUeVkM4wCmHRurfp5iNPC1Nj
KPFrYy44AZTh7E+TntbAjpiAj6duhQLC4UvNBIsXofLebVNo1zY39F+Y6EwA5vxI
UjbVVkvyzRrj4WMtNtjMKq8B+LeYxz2pYL82W34bqOFkrn1pORTvu/w3+BldoQCE
Y6TFUR+AACPH1nq9wT7EDSjFlxUMMMcYyey8jktrtAWr9MYDGU1tYYWDPPjwzyZR
Qda890nwMXpYLf1SEiZa5wZMtdK40ZKYMZlv/7mXNa5/H431LFUfSDIMJf4YmU49
n+XLOgG7x5mwJxGl/YCSMvl+cKEv/31HNt79abh4VOjBuLOaIK4u68InuNffHJkA
39ipZNrbjuWGBomogt1K3GxoLBw68NYbW/rdZ+fMMZA+PzmDIK5l+LF+FgaGPgcm
rc5UFdWWuWbZSgqkTstMB34KSRzivU6viD0v6NxGIzZ/VA+PI3zkCe0CnG13nRfO
Vn5v3bKf7Cw/CDFULNO989oLMHfjoH3mJxaTv2EB15Sb+qxmSa8j0DY5as6zwthP
DO9QgEJ3GGrtfbEMnduOseH7ViTx4fP0BQ1S+jYo76vwunGO51Vu5YTKIa4KYcyO
wBUkjXHfz0nwKWNWzfr29npkCU7I+MF6iPVUA1NS/YUw67ISPSxvvVCvqshTMXBp
f8HOmgfmm68zN+gdkJXnb39HDA1HeAz6GsHD8s6ursJEuuMPB+fBr/yJHtOByr4T
MzkWrM6FZIzD1fCy01A9h6kYQsKw9hf8HDc4tpBoxq3OzDpR77t6aDHM+IK1xI2W
kj1Z9A2qyBFFJ0FTd4bTlpGkVwqPXZF2xaQ0jgY2nzwSaPTWnPQqlB606jPX9pL+
OKdc5Db/XJzumGaUqgt74E5fhN6ntWFhyp/TopazH9Ssrj69pDAqBTz5pKkSUk9Q
IinDKJvVdk3NBnHjntUgUkpxmfQPRgGYpCsptzoFedzYpcAcn/tqeCumJ87IypgI
+gX6B6Mr5JW0tT4c9apBcl1XvpXVE8UkasN0X7x2LXKjY9oSBhswDyasp3kRQ3Nm
amcQHznoc9167bekXLtDubMg6/RjB+/iGVQ2iEr4+vf6beR/b62NpUD3DwRAy3Qr
5T5AYV/YguPCCn+SZtGck6hBMHVhd9ma/fQKt8H2v9OfQy53Zdfkik1Sltxtd4Fq
nWqaz5a9khemPDvbZugT6iMU97utOQzsWIipOodBJOBeWYxGiEsjiA/O/9IW9wxy
VULjpuw07/K342RGNpte4BQL+T2mEgJD+B+jbWT1sKBKrtbuq4hPKjCx0r0ck2yV
0Q+bRXFXHwQFNTSCbKp3BSiQ8x2enZ+Oa5IOvt23vgY2kiZj8490xvHj9MPqhDhw
THUoTMM56WRzAvwJ4FZ7F4HSklAnTjJZXIjpTcyIZCIbXCM5l+rLxnSoSXfi67fs
iiZM5RPhT94cfqm4KICJlPwmLLFz8lxHLd4eDPeRkgYUvdP/6EATTT1E+pofshsN
KEAeF0vjgv2Ns/xKKQFJv762DKBfo/jGkinRYZJK475mBY+GMRBZfftoqzG/iZjo
3qf4OjkYI02yYejnJxOUGDcRX8pK72rl/HdDmn9YnzLMtokYObPkTA7M/CGZI2QC
3XqX+CJQmDF8NMFndgW4wCgWj2MM9Bhl/wMqTQL9Hbkiqby7st+3NsUPvT55IR9J
WEWd0DdcUgikMB+8Ee9MiQu2i+cmf6JaTlyjWivLtP6OF7KXnlGvcBUHXAh/YI7Z
QHnmzBSSZ9jC8RDn4Osyqckm2ZYxB+kNfQk6gebcSuRzbZ8auTv58huGpTtUmuCq
dO7/fr2BPPDyBv06qnTd8IKXHtN5VxiCkgUoKzjf8wpudBjsyGrO5suh2rWv/N+D
BW0/i9wZ3+JtB9R+qc9u0yFMuhy8bdmfe5jPisYsDiUHkAFdRJ8eEQvV0tAcplaa
2TokPJgIcX0TEyoVf7hfr700nvKFCwuzbbP4WjC65TuSI8oCUdEqDQmRy3BnurWL
i2VwSEEZ0gw+q3j+hFZRgPZZFfrOLT6g4KpXB+PgrkvtEzXvCcSfC1Kcw6MFGus1
Y0vmPJ6sWSwvZa9iQL3tOZGSTdobagmh5VGeYVKDSjwKCIGQE/5YoadDxDOGXwle
EkonLMO02NVpK5A9mSfxXl0RMXGH+HRI6AWVXMEgDwk5CJDF/AKxkRu44iwX1eie
2ucbSLAkoMi8Mo4TX9Zl865QtjAwMCAMHmw64gx1MDBlHe3zwlj+NUh8G+RobAkG
6agZzy+QGenpBwZzNYe8+kMzMOh9d+hN67eANIjRxcpc7wcT6ACX0aJpVOBetlkt
C4UpfBufKuB13Ha9Xmf5HwMROiTqH8/LSNReFx9D7EEuZ3+w3V47gS+/1kF6nY+A
0k/JukHWCma1zUfKbnqIiWBFsYNkoKyyvo4bKKEUl9ETcHGTs5bbeF387Srbezlu
m0o/By0WZt7S6K2ONx/xxz9LLmW7yINB6a1YR1PpKFKjHLujtYFnUW61v6sG/TTo
ECw6IE33+ydfN3r1tcKrhcdJJ53AN+7ue5GCO0x+heN0SFh06Vf00nkxDH/+/5NQ
s2e7pEhm9zrCzpgq43tsw9WtaZ9n7L+zDXzpjB35VkGw4JXBA2CTyQwFky8YHsXA
Ok85khhEEtxzcKymRiadcmafvqeZvunURZweJi8OttwuQV3ZdfaoncLb1iVDJIHe
5tVyybEh+fK2s9M1qdY0qhPsFZYlNKm61fcP2NgkcxIhUWa0VXjh5G8tuADMWBHB
J3PMN2qyrdjKruezFbnFbnpsnKNhzC3uzFIROOD04eW1pMayp285ff2Vsa5Q6iMd
Wuo3kScjnbMGmaXnSeUFkwzF56s9MLDNaTghyCgboqfO+zVRUwl8p5XNZkhoNGYf
ykoB+QHr5EbxN5YV8IEnGOR97Ur6RzWIYQ8IPXze9wexaw3HYXcueJNxwxNeQDSR
Bv81byK9IkELowisWGM0Jb3UeusZ0RlHutkgv6VvSoaU1U1OsmbrxbhbVqyqWkxd
nsFUQAISHUi/MTme/TMJC6s4FpbFN6fpKuAjcjoHiMuGW8YsDZaFzplggeFli9XE
/Y+ktsuPjeS3oZY9PeKAontuUnwcGoPWTxrDa1szi1ftnsD4gcDGwONZwvNTJSM+
OC9LFfYlh6xP8vrTNaB0OUGvjusSXSnhSGYG3rO9BpZBWP6OWBfjSIFCZCeZmBKe
8Hdjqn2kcFagv7DKj6ec8LbnlyeQNt9DGdkmXAOE4yYk1pZ+5BpwOOq5dOM+a0Dl
8yGMdX319s5RhXZL+P9vZyP4vwMjJfk0VqZR7/QAdmXbGQVCeu9MJbvB1C5GdTIP
cE0CdwjEFs2sc9sksGz0l+xOnE0NtFcgELU5g4D6MNDENgr4cE8/iefy2a3Wb3NN
yKdVxHTjTqureJKHHRo7BNqNuxMahncGxCmJ6dkltNe5pN5GzC6zwzGJWCUICStz
qwO2wb+5TJ99pVSAMn0byDG/7TXYH34rh1Rmt0eGLvox+sUMRGR+F9XtkCJ+4b+c
/VYjvwLE9PyQG/+jqbuipEWj7XIBogepHoOvNIEy/e72ld8nNhWLC2cNzps3yYCE
rcckXoFZ8gccUD5pIm0JABEbyYuUB8Ex5S7bfAM6hq4XHMGWNZdfWPeG1nGjvbiJ
7ymHmiDh1M5AUgykjinzjg9wTblJjDT+h57YHl4BAuQ6G14n3V4n/EYgrgu8BQQ8
rDtG8IK7B3L1QB4p4MmGucSNFsHYREQbvzs6G7sMO+adnLl3VaFsrWBZT+g9zLlJ
vgZsYE3QjSWfBGyTb2bu5OAlKtvmErkeAOCMrA932homHRteYKooGMBoQ3RPC8bN
E0a9yM8I9xnIcXh/ByfRNWts2nRJ9AYtQkkl/xTk+WR4xxUNZ5PT0tFa0lO93z/6
VmDbW1ahy/mhCrJ2hgx5W77BpTwR2+1LrMrGdJ0DsXy7JZF8FrpnQFr6aDtw4I6w
bLwnfjhWv2l4XLeDW6kU1RBuLw19MqAWya0bX6/aIzIDyUmvdeETzmYg6tp22Vxy
tcsPGFDqHBnmnkmhZO7hJH8RxEaKt+jVvIsFTf9EwSGnVT+iY+Uu60lFM1yNDN4/
JdTmAOxamYoJKmdTnYKZ+0hq/FZUydX5Glk6iVjeQXWR8aexg8KcnYQ/KmogHTCg
iTG0K4DlGh6aEdaademFnaJX9DTpm1ITrBHS+8MSFATzpwSZp2t9pr5sn//SaSpY
m1T8Tf2oozD2HSwC4OgvWXB5oJdnDWbvUj1BBwQfTwjflnv6MqZFGSA3ZkP6zz0Z
jXHdxjVOBlBCZEYc1EjlYScJz3owqIsyWI3uPAnd+uuqIc9t/iXTg8b3tYzocQcE
GV+Sw7gdR0okV29uHgdwOCzSQJYvO3TfIuAOGwQaq1yipu7dndNXuLj6yvO+FIgJ
xvhqd2yrd12lq43CqfvqE6PbgiTJjpgrpn4LZcjMIadRN06vaIbL4qV6OfnVUftg
cWB7Kf1DM6VTH05V/NCoddIseMmwU86uiMpuGjGZsSpVE7Z16ZOC2GMgddL3aiCW
yXMx4TYxOCx9zwjNfsfNYSarTBspkTI1UJx9cH5tS3Vv8nolLTZwKQmrAgmGpA+b
djUOET+c6rB9AjDw52WsfplRAVM93DyUTH+29YBNLh44Bj1xhrBdZLas8MUToBaq
upgNi1+86abq3QliR7QJTHirXGb5/7Eg9EW6UaN8M9Xofqza6+5vRMHWNOB36YRn
HevV81XEqNpKmUTPZvqcj48BLAtY79YX7iN+YDc/6Eq+XPNsA8GoniP1IZWYCd98
3/dHNv5cuTUxvcc/rvJt4to4qtsJOox21HvE6dBTJzKfc45gL3+a5DZoDxnBRvCn
OqXYDSMLaAIbXI/3cMMPJDppU1NiKf+KjNp21AG7eQITcYckJiSXJ3a+9jzWOGpI
ysVR9Og44o/8hsfJXwDNJlfBeQQxYxXwZa8HAtwb+BLnprGUjBTH2GTWsVkTfW6e
sIgHZyJxm9/D+GartXyb1HDS/RIs32D6RNOsHZZAWHDsmvWcAKmMm/M5smAXUX2k
z4ALfWZny+FlNZkjO6EHVwAdGHoHVat+sIaBJ2zXR4SvazXSmHvhS3OfzhI0OIlq
A6/0tbSF1BlDnX7tpswSaxuHN3z4+KPDXbrmycpt9J+h3/YozNfhDm3jru0D7IwL
UH4H51WSsm/PmWwDFSi1aH15AP11g+VFTNL/plbizn3HpML+8lYGj82kZ3w3bkQG
10lv4Z3o+fxBL4RL1J9KtNh1d8Ip7zMVYhYoDEJmhgcm6o7Hbenkb8dmu2MrX2E/
mVIAL+aWtl8UaVoOiLLzirpTSf27y25eMolupYaGzwbqOxn7wUuXCITq9N2vMbmz
S2vlgYbgXr6nQ9yjkT70E7UCQ5U+KU/KbNiorYXnZWaGh3V9geCEkLUVmfZAoD+N
1QxTWjTikLNak/YsIvrAUTtJRgxBNxCckh/1Ik01ic1VFW6/7wPj/y5X2PTg3QlO
67naKCMa49OeK1ofma/LDTzsgb0fCnRI7UwKdj8lDloCdZEBvy9gigtmiORAb7di
FRXOx7CyxL3B91oZj6U9ebntgSdyJjTjAAJWLqwaZPLjfGKfltbVgTsg1yBr+bF2
f4DLboh3PT/Ko497r5eJiaSwIAosngo3Qwu6ikmxj02C8dzwqMseHzg02w46c76v
KeAr8+Po1MJIq3t+m32V1DZKhQqN8NdrgOLByZJMeVHqq9e8TAjy2yWgwHYf61Gv
7tsPP2NX+66L9d7UciSZixXURcO42OX2PLQtJO9Vv3LNmYVUgL/kjCm12xDr1bly
livcFQxgZ8zX3ATfy1sItCyafHblONF4Ol8gIUgqpol3GsMhrOE/jty2Z2saY5NN
UR7AomVe+t7A1gyMuP7WuRYemAGbpeHjmyrWHKlSJDyRv5Xm7FTmmSTvp+SSFPB4
MA6HqViUaHIInH0fNyG+ith/o8SGLoj2aJ2EIDQPbdAzkQ/WaqGW/y+KpOjTu6Uw
FQT97fhk1u5EnBtqKCwj5DUZSyddo0/aaZ1l3kt6htrIr6JFhMX/2EW0S+48hc8+
SXrGzLB5CBpMb5j24DcffUTjacC5mG0pQpDUbtMohWJ4sPox39Fj/COCAOPx4yAh
BRDo7bnO4LEa44y7upX6rRP/F1yQrWKzH4of8YYPFxDuGiSlWANB6+omXoQi5X1H
/AR5xei+Brqh0zmCxpEcYX1lHdv8s/B2Tuh5qoZWm107M/nai5LHOjcPAc86Ooy9
jYqz2nhEpFDuVRHZzFBpaaAXzKno+rcDFTkWSJMUgCh6gb4mhz7bkSQjJ+GIJYgP
q8nK7HKb73EkEi7zpDeIOVcCK6PIrs1maKzY0YYcPEJIbFod7acvgNUvr+Cn0OFg
RmvKt15oVVeUuLiS31T4/F58Gx8Xp7uIui+n3bkSLNUhfaXRJEMZa1nuu16pHgc3
Fu6dGsMad/bzSvehfXOaGVMFnLEsgpGanSMHypI78vjh3b0cVowTVnKc/EyPKOMH
jHa3y3AuX1oUrlzH78RVI3Pl2ZbUJ3KPpcC67NC9uB6c4m/GTk3akgh/nYmvPHpz
c2yRyCav909DWP2FxPy6mkowJ0r7MLhwR0PrYGXVuZX7c580aY+rlycoOPlNmZCN
ZDnK8UeEmKIEINuYQimpz6GIQa6op8wgz3f/zdtAOLhk54qYP3qRC4N7Lq+Hf0Fd
q51rqpqxmhi1oAGMe0TV18uA07gg9Z+ILeklj9GM3IkPjR8TLhmjjvP/XCvSUeEY
ZGIFrNAAWolvvHlWQMzU7bc0bJ5dZH4i+0sakwoOcLAeBurYw4lR14rBqqN0sgp+
540ta8ZmHMqqwd1k155EYVDN2pyA79xSW5V7WBcwl18adha0TzXT0Xh6ubWPv3YS
KIodEaMkLrlo/fjayO3E95KZZe3PhfAEBwoQO9gsKf8B6DTJQ6QJ7mgnxYzJzXNQ
Fjz0uAlu2Om1aGzyPOGpW4x5rtxq8xqqXQccB+CpldX/qAgWgzp6/sFH+b+IUkEL
NmQbsfDIfU4Aenl01CjTTBH6iV3Snnkp517ypRN5a4V/TUhu6IxkeA/l+Uh41JAj
Hg9HkI9sP+vc92Yvw8UdSWDQAF8AkeOEnJGEYaW6BmpBEwCqBwM8/ugNLoEy5N1l
x1ZMxmAeyuhjTHsROTnqmZtVVBDnXfO5upZVQ8v/UtXqbLn6WQOfy1/MOKZ7XKHb
NalExAVy4mF6d30YeM46u+APMlFKXXZ0gXSQ2/29C1u1lJUfX35en2D6Xv9ScWmH
TTLvLfQqeQbxwj+mrYp+G/U4c6bQ6b4SJHkrRlOcMycLeF7wUsh7+SKUSYA2IV89
eh9elfpieS+Byff3DiBQr3EiG75JaTcWjjMFhHIMvYkQvzUDMcBIjIYMTHafXbA7
MCfVH5j+CeJKgU1rB1hMKTxGx3XgYNEADEK5QaxFLrtShuMd1V9HubIeX0ljGMLF
fkjFjTiDA9PGlKrh/BroDQ9k/ZYpwYpwRzZYXaBGHYB1Js0Vi5/I9bWoX7tEsKz1
zc1VaSoq5jvZgbBHzoGOb3q8A7gq4nL0Nrm7GE2L5MKsgDS6DOMWrb5znGrzDxbJ
VINaqUL1SDQqvkPzAZbrRKEd6N1D/FrJRG2R1nJ/xsi9qj0ZKn7dkaX9fiNiYXPL
bW07y8jYrTJrc88IBDrK+jG7//4bCLQwojkR/3tOhFkcZHqc+uagHATTM95Z5B6O
xxzCz4n5vtAMyYcK7uerk7DJRCDwhwHIiGGJzieP486OsWO/1WTEL1mspJMGn9kt
vu11Rf7PQjv8219/AxSqWukZIU1SMyUHDj3WMZUqdJpPwxPeT2iYb3UQZzS5am4A
aopMuDImd9VmRRe7sUuF2jwf2Ugzr4dg8eW30LFv7nBI5ne5KAl/QGAx+LqSZ8Jy
azi9p4/RmjwB97q5zEj00FNa+f6R8ZiBY8yuRUHkwWfzQicKSIgf1hYoHYbpGKeM
ReZkxylBNPjbv1vAK9BNui5kmDa1c1DdozSFL+Puwdf6BD7OXnf1NIg8qtK/M1eD
/HFkc2MOxPDkpFJRogGQnKn60XVJ7vBFDzE0vqpztUkRc6Q5gTwy5YxKQrZsx/5e
tp4hQMBsJXT1E3GIuA6sanRd0xgsXf1UXXUbaelC7GZCkXVCeWprL+hE3Z4AYQs+
05piBwrvEGIfQ/LpVzSYOPz+Y5+AETbpB4kEXttCu3QtdWuKTBVK4AspSK6GMnsZ
SD2Gj9VpApDn9wJNGxJ1IHqAje0ejuYtlNF38zTvbNGwLF/C6iNLJHsMcRYhXmTZ
dFUGjXX9L0yQYPmGiFoEhPZQ6vHo7oEifK7wNDjKZEXMjIumnmTXN72vry/n4Tsw
922ZhmMPex9/3ZwJ2+4BAP5KCDAo8roLaOM4luFjuGVLRjZWRQSeiCbd1NU/OTin
dqi/tUeBn6P9c+DO8mixg+AyzNpf3CQfoFyl2kxgCeJSo0k8GwkkgTgtSZ9ZFCsz
C1fpRccJKqX3pVh1TXiludkLt7aPpwvbaDTqRXN7rZoVi4sU4DVCs3HbZzmPbFO1
0j3kxEtHfPPvrtiyO00PJz3fFMuIgXsRyzvYDiurUBw2Zpp9I3Ycp605dd/IItvI
sfuCSLcBn6gJo2mtHR9lEMoVF4IvigMbRzt3WDBkU8OJexjuWpL4a5rwvLwzYJMQ
eO+Nwb7td43AHrCbS4+6FIacPmuWYFvL8G4UY9vAaqowBD2Y4QowEOO1mXkjbjxk
kf6+f1DeO75tMu2M9AlUNBcypd1BO905hDGvi87CSIriF5Dhn5OwnVfY7M6W2R61
B7/cZg+Vv03B7vqSgDbD8121BepEFjx+2C9gT1kCZ/wXKZzjxAJVj+UhoIA6usyV
vW3WnA4UupgpoQjtUEykhRd0/7eXeXQp7Ktv7ARK1A5EZaZEF7n+ytoMMpn+TiYy
huZef3/q+waQUjbH7/9EwXEI5W2a61B/QKnAJvc7i9/k8S27pfNByLxx1sAhPJO0
XFBE2JXmmOjUtY0Ui+k+PSVs3ExmDxmH7uNT4pWEJfYRTlE2Xqu6CbNVamSDUZGq
z6nHCCoXQemDKEiNZHhS3a8/zytgNM1ajxlCvLWHOFGSs1gyj/K4S8j8E/1seegb
UpJpqW/PXQ8Rg7vGAs6OaxUMOC/CBQKugtqbBjIun0g5jAmJ1j+HrLCXy5Rp+QNe
qO9zLHJmE2g1zh30/42uneZuKdUKw/IMxw63zNIfF6YiH3qPa/II38TdmG9aAVx+
+slyx0tyUyxrOqQD31Bm1oJC4amxiXijMUIqjscjGw7wLfVpEYdBiH50tUjdSiGs
xEe3dQtVt6OFIGQIZXodqpSSz5LV4KDqdBy0iZMplOOD1LsgwKNeSwbjtndMirLT
QgKLUVoM6ltZitjGoqJq/xUDzL78GW+aDfSUV+vzWxGFh8Ci6JWyKuOdVHZk8fcs
Ec1W8jJgSQmYoKEdk4C+MzRHgnLaWNXSimbTD70M0BjxnMLo6QB2H6hc3t/nE4Kw
iyot5EGM1T/cYYpu+QoR74zGWaXfQoWqhByimRP95D2g7j8DB5K3bo061fSs9+yR
698A5pfbmAX2GWFZuo8KOWIMrC/MhHBBGYGf6cN81dHrGJ6Ritj3/IbMsj+Ho0Yx
kHpJ+yYJSoab0Znl0/63gPSwNsniWhLvGRGKOHw0AGS9i7EFP0rhM0iMMCcLoboB
FiNIypDLlPr7WWWGKgrBsV3ngL4bLpgmSN+zeg58GO83lwc12wwfY4mgO1hswFti
6ahRyIAvq/Kov0gV05w9qNO1NtKDEYN430i7sbrOjPm2A6BhrijJIdQKKV2iDD3R
tb1CmUbsPYGP3RekIcIJt+yYV7iy983q5BSvjaiy7l+51PorqqZnhY98ZmrGANSI
iNOeZKHoDltZ9zxGxLEpopD/VObE9NUO1/RubSNWiH2X6Ru0z+LEipWdL/IyNCfY
JJAg+PUKOUEwsox9kxuF/0m2fnTuwMMbvulsmMfWep7cJU5VfhZbO3M6XHFbM185
KMjUrSygvasoI4H3DvUBlRTsRDxV2KzwUl8faWQCT4A/nWasNpDculJAqo5ZT1eq
RQkjcOFwE4u86PUiWRMPztqiRORT2JvFp1OF+FLJYhg6ULNmsuoxEfO85AcSvlcc
SxeYplVVaGVxoFlRRO4xowKaFHqOZHbe6JxNETunGXDAETKoa2gMe3fg3TaqmEj0
RO6daheTwGrluFljQUm7wPfHZ4HaHyjKNSztkG2ycAeUvRN9MgjSLzBUxoeLja5o
iLV1fCIGRtNTsmfRF7AJ7rC3tjsNs4XQgLUqzZD6JY7+IiDYXEDBOgBAyIFCk3TW
Usimy7rtLw8cD0ea4LVjtBWNPqxaIbryZiPOybLmvGBvfeVf+cOh0RG7RLqMTYly
7e9yS8rwB+wZ8Vzi8mVIXHYkT+WRHXMrqVyLzhVPT/PomfLdCZwY2Bbe6nZkp0xk
K1sG3u/OkvxEN72mcOqDSfhFyXr/XZmK3I/HUoPP5uUyE6vLnT1Wl5TzMDX/iBbN
E2iNeHUE0PuHYMaXkZX+SZ5V3EMW34BZH01I8f/AFJNGRPfk61Bh4ROyYX/xf5Gl
QnxSLSooGdzKSshGd+cLLmereXftEIVdjs3pPlFiDWjTcxz+kBpKdyhXiG+hqSST
OBoXty+LcKAXaweKxuaf4qNScfXaIzevt6reAfjDrgavvIBp4VPKxINk2C/fdAwu
xl4KcNEOfk4U1G2qv5z8xvSuRhCLKXmZP687mYS5nkNx07MOfKuR3Ocy2B8KGcoB
BPbYNuefnT0Cqk6vz6/gJa4nOiHCUzKIktZxmrPg6Z/Jm2iFgSW7IiTP3RmZlEXL
mStAAU4K6U8gh7Xs3RLa5irykRg+IVU5CDWxmBq66Rz89XQWE0i70FPQtgNnpQDg
DKBbLhGWLgEQfcfuVTEQgDra/8P2o9BLmROLGV/ZwUMkNtNnbc+71+KztLeDX+PB
FXw73vGSdulMB7PrGvcfuvFHIgtKSO6TjzYRUTwBTlGeyP+1cFavfja/6f/5zA7e
dmba91z0bZvseQYJWUjNtIV1AnIMZAXJWCyQLieIazY+CgN970KufXEdbp3aDoZX
CcCTBRu12VtFHhO0mlbcHuHQ/23CoiNyvt7xYosd6lRE3U84CuJnWA9XVb7pt5NT
mIT9aNFR+D5PHrHmZ4NluAJWqp7LdtKYEKoovlPBnYdVPWx2n3gHdtWEOcL5gWyi
sh9sRX0GnmaN3F0QcqBXaq0/AsNQyMtPZnEROhPR+I1ZOdNiD5otpIQaFR+nefFE
uzhXv4EyVA+Wa3r4xIIciK8wfFbo/khoiaczrNEQkZ/GpLIQtz5eIkAKwY8u+eYy
n5Tt5lVdJawU87a/JIVjkvJ7euts9OFcHOWKmf547YpAm/9drahezfiPnPUAOfbk
qqnd8Sshbo7I/D4j8o2ZpRv3rKmcnzPAGUdp7y2S36hUD05dy2h8fWkfsw2ggtSu
t4dzLiayBRPT7ulPkmxkkAVz90WntYHMnJII5rhRBbOLFN1nBKZH6lDXJn5STa8l
qPluqFYaDU/XPL0Q12JuzsRt1PCj84jHe+ZwcPp0wjpsKxxElWmTWBrdQlAbHNAK
44JLSUsg+fO2MVfMSauQlS1MspyWFWWl9ycwuvaO4ezb5wOnld0i+NjfXiBPpzwY
fJrlf+a2r2ElkTVLUF8wcm4yljVAvtvcXOLO/KcOsEBlwlRHgIjH01BOYvJB4sPV
3WfVuBTqTF/jJkV5PGskvi5Ko9dJcTVScgEw1HycB/xW00zLBUnqH7poxf0McKKQ
p8u9qZb3jojhTW+s9TlvQctTUW3S73WCrljhgAqAP2wn18Lha6VZR+RFgXTBxx5/
koRo3I7hPHmpGGwkk6LaSbdXwNsfiRusSdXoY4AkviXI/eD5hrYLbsbNp9GBZxRZ
yidDy1HkDvjkQKnWz+GAqaJHNSz85PKDfnGp/rDMGzc78VvUg268/BQz3HBbM+tE
QpfrXqOkXG/4hXH+GImqnfILZ+iBLKUgp47WbqjxgILQjdIJp53p9siV8heUhvLy
IbHPshXKpHINBjrJ2/ckELeNVlcxyeidB2/7j7QozJAorSfzipborM578jLpazI9
zmjzwPlm2aSw6P9CH1qy1Mb5sGanlARhRPrh7ThY6Egnt5tdNCmyNRVaLPJmYtnm
MCYqbHm4nn2EYPpmMdjBDC2Lzzi6UmeFOiQZzciT2JIdRjqveVnWB6Lco2xC48P0
2JPdpErGMPjj5a9v6l+3l0uIMm+eD2ZNx5DJkIWDJqhj/9hUvPrGx2/W0ML0m32i
`protect END_PROTECTED
