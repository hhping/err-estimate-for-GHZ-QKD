`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCKWXeemntWR9Koqr0jngFBtuDOGaMs0K7ktRcqAXmTVfNIrJ6IOveqXZF7GVWNN
iL1TrmjJNaPXpIrAXzQdcfefOMU133lIBAl8ZFJpEB+6oThQuG/Jo58cpFgH7+zw
Gr6I/8vaAcfbClTpqu1L0oNZUtZb1LVlnB9LcOCAKOp0Hxurpz3j+C+sRJZFBXTk
BrBGnLr+bjh55uBgg6e8R66IU47vJY/GGyScnf9V29XCcT27VYVWf+ofX58jcj6t
+VZCDn+JlbVRmcd7teqYr0P4wVfi02ou9JXccZZNp6ZFdjcfepp/OH0s9gA4+ILb
LCz9efY1FPPd2RtZFGFheMGQuR01v0wpQlV9E25x8NWQOTAI5iSoccZhFkl/W05l
dw38S+hvJlEUtA6J5+7lQs+Di0qKSEXBJMOhTn+4/odG9h9QiAmN5DqpKRAGUI6a
Wh9ssPBH4i3guAR1MxetnJqo5+gruD2o4c/jiJv6m5TUa0jiC+umWKVjOa/rzIHU
1zJi0MOV10iHCS0IuIQA7+aXj/dw19vED2qQaWIxdsEXbBxuAkPJxdgv5/aWgci1
Ed/T6Ff5zrvBE3aXHyGW/BsPHe36xV+pTN9m8Nh4YXg3hcwU1v7FRVAfzQCaxOml
fm2EM2v4aGmx9f3k6LgUSsXaZx6y4h8zoXHn+T3DwcQL7Stpe75KDgexHyyJgdBA
4hK7F1RSCL6PgWQs0CVYP+b+glrpqpu6X47veqIgArpP3l87c6R9G56N634FiW02
MRdKQPHRRBs2fE9uOHAFXRL0hCXJekP98/Vxh6dx910=
`protect END_PROTECTED
