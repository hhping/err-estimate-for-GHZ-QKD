`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R7f7GrK9oX++S2S317UYVGULJ38ZQOEg4FGUOBvwc+v6OhGepF0CcHR+CH2SxELS
m8oKqo1PusyJnRo+Edv0K+7OE2SMbDnFE/rLntLl5yEVIekd4pfF9rveaHfwMDus
2XDbt8rpXbfM3Y8MGEC8zcuKlje2Hrpv35dfyKgNXNCR9c0RpS0kXKw9KZmj8FNJ
+7OFPeOtXnrRU2TKhlxXjj50pP6NaELh9sALN3A7eAT1d/nXIuZyHLxkGJSyZ3df
LnbzsDF1szoPg5DaRhFL83h9wn6thDxHxtlncbD/nSXrh+6VacyhqrYeCsUq+KrI
ghx1+HrN2R4VQ9GRthbUJuYC7Akam4uY0EP695ykG8GMHOBa3t+9+seFSg9T4pIJ
/bxZjazzyRSNeeoOcIutZvRvxm2wkKd+7wciWBU1U7gE/Y0SOqPp8MbuemXrpM2z
v0/nLhJyD/w/93YreKIbBjWUPIzOLUSjF2++qjEsI+UEIrQcjQPweisE17LIgtGt
GBTFbLu7OoqyiJ6UQPOoQYNqPqO9k9Wr5Pp2eRhhvLLJNCWNNWriK16kAE9hWxE7
M0xwqbDPgNEL03pMBILma5AM3iw6yLkdDUAepLOFkkL4kIQzCDfnGQcCISV37Gsf
BWoLsbYVHf7tHn5/MExyebXlZq0BPxWFuNiMUHeuQCTBxZ94F/KKR6ZSB1EQKhBY
XLJCOIYwt11T+sbbRd41zAuxhUaSpJpzBhskBgrr5ydAay4LmMJosQz9zUy2O47C
BYuaTgmDZly3JtroDLvHmAaFcMOt6wns/If2sLhqT9cxRDVEQ0Wg1k9aXWOX6w+F
qJ7gbITHAjf3cpmSeIcQZUtAdK3Fyp495G6KqSkBtyfkVe81lud11mP8OEcFDouZ
SKqXPcFbfI8IAdsCH6oE4ZGOD1TXjgm8U7uCucNGOdiwJ44rqSdsUL8oJi1Y3K7i
+u5LlEXvJW/HxHME46lcVBJlfYmaomlaqlK1kRtBU+1KX42GE9mi0XD2vgC8fipT
b7CKXlGp4sDERnJsMQaKH9VTwCTbPGsbWPIZ/vsMzYE6Tm0l5BPtIvVpTXANQHV+
cLgKYkLeCGUzpfldt8P2vGz2eASlj+Fbot+p0408i+hRCSdFtJFGHfHAZf1zCHKB
VoiVe4kq+1iLApcGKuaFU47bVoPAz8RShrSO9b6JdALNEZpvrHZfBr3orc/fjVPP
g6EV0rH+PY9k9C1aHsbxMQ8/KumyDaznyTqLtq7MlNovQQuqo5VNWpUSJCPkaD0s
YzO22PcESzhlxhA4+m5AWNI+xNwBkFLP1ggb0ZY66qvFZiFxapZAN3aEK1ik7aoL
PI3vj27XVi6gwsv2D0hSlIiF8ZCNbhEYGTG1tmNTyeb+gy2AlK5iLgYYJJVod+Ay
DAWR45ZE6Cg1wtj7Bo6zIX46Nzn2X9t8Kwg45ZMAArjlxBsQw/ReDixnOItGwR0F
ly2cW91t2eO1r1aQauBXzWSrYWtCGsIhdjPFRFu5k2JPDv4o79tgWGRBj38AiqIt
8Rr0b56HitT1D8wfThYe2NhKMocWTp9d+BpoSrgqZAhS2E2Zvv6se5WStdnkMXgn
36M1PboVTkZwY6yCCP1KV7gsCr6nup5tUhS2uIkTO6V/Kjwb22r9p56fjGICLRlx
uMPjDKV5dQxOvcCpKH3sl+zRcryQfOulOv8KwsKigvPWD1iMLGkDB/yZTJcXndMo
kaFqwFYL3KCaXRdl6MVqoATqCJ/uL+Tb6emSa30AR5qx28SBxUl2/BiGvD7gJHBk
EiRxQGmEY2TM+YxX0AH4lSdTpcVC4ULP8Yw2mgbMx666KyihbO4f5gFz/46tXtNJ
qQSyMyefDFVI3k+bhU7N/5NPgm3qk5PtmW0091WcLvGFudHbwzSvBe8dZPzGU9pb
o8J03z2zaz5RlpwQnVbcqKVpiSkd28ACJB73VQFdIUwrNxvxvHbkoP8c7MpJM88u
bwCeblosJvPfCl2tI9miaA==
`protect END_PROTECTED
