`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pyOt31vY95us2dPOvAlSae5n0d8aFf/bwyfjlcY0fqA/5Q/lqX9cmE4xR5Moyijm
xB5J8K1ez/JnhFDqKxUc9V+eBmniecMcs93MPG6nabBYnHxlRH11XcDMgdMJYm/7
sM1pMtxTjsQN6l8dccZpGdXPkh+HHIy/4EixJN2I6fx7QNceDWC2720kUR+FsST+
20GaU4a8w5LqgCMAo3gdG81RzJpPGSjm2y28kuPlJcKC4NWRaytUtntpAQBhZwXJ
3Xw8eyHBPdsT41ltwrIfKO8r/uAFd0BoTxxImciXPeHomNEtmv/mP6RkzGBLV/Zg
actumfdQudEqITNEl4QxronJyyDIw8PW7hFieI6hl+aqyU28kGKpJgLQbsJGPRcP
zCmymIGYEcIc3jrULUzUDAoDBVDWOkIZ9zPCWDpfil+YcprCr9WuiSzjFYIhD4hY
pUkgYM4TdI4PcuYUpTxAiLmpDOVEe6fPfW6aY751ROIbElN2TZcazLaBAcKM6Xwp
FegXsl/t4d7o3IRgcRRqJTT64Vek/sq/tvsR8eBry1YzZCsNdfy2/X8YlZDo2Mri
XnEDXVEd1NxCV2M9EkYsTTqDQRKpnYf2qaZVehWV6VMMFAsmHUKzjMpffqEu4SVX
9V2yLJuUQ6ghNqtVx5Zdt/jY/yFtBQm8/ZVgchxk7IvivAgfcOV0mSlwR5cLIlOp
/935RcAReMxNL24B5/EvgbKFm4EaEI1kqorwAPiU495Hui0RzbJbbItP3NWlYR+6
f392yCZCM3cKhFEy/DlI70acB+iAqOcptCdA4gMbybVA4D812fmagFtNfOE6jfsO
Rt+YCIp1sHNvkSHtHSFixLxOQlT96bhsgRp3tf2zYmxSIqi4kRh3l6Tdhpc4xaCS
j67WrVnh4FtG0B3dvY9xEMJEZrqMqUYmSelG4lgY+u75MW/MqY4mMT4sMZPXwX/R
`protect END_PROTECTED
