`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEehtH2tzYmnsI+pwCqRcfBNgpRsPR7LIdOz+akcody2qepVvhwiE4ZO/70g7Ev3
k09W5RrVjCpghrQ1fnzEtBN6cTXEjHI9/WVQgkJmy3VTRDHy3lLrU4c06HU2R87Q
2gkg36OEo456uk/Sk2aznS2+4IMNHpRwUT0lKeoG9tgNgJpaw7BUyEkNP4DnBu6r
eh4GlDyx7crRhR+0a6uza/zFXKPVmssaEXWLOJmdn0Eljy+PxtxFmewvNDoVqD9U
ZLXaEuMS4CNwn+CNt5L/Jw+JNIXs6Apm33cFP+5aM5PPDmg2ne0AzR1pA8mxHYA3
t6/VFi+ZCRCLQR+qwK8JFvHfuqyJrWy3nhC/muAowRhkpPavKHqxgGEqAhr3nGKI
`protect END_PROTECTED
