`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6cte4cR95QqrCDwQKcZtH4vJ3heNxwU+udcBoa4jttf7LZhX40k1yvJ2OG8EJA4S
biGkDVwMfkcPqEvjFp0N3OSWVhhsehzhL6bD+QDfiSJ6S6Nv3wwbvf9ZJpJbUZea
TGhgVrMwb25U+qYB5j/MlEoDbVRO46QRAJ6ETRL7hI1+gWkVCkw207Z9yFBZKS6T
6RC1+lgFBsV6FtW/qd8CuN+sQvdX9Pe8ALq0Mjn3i2sank5CqJlYbW025mnLOA0u
s8jV+Oo2kcSU1hOm+tgLKp5jxR5QeeYw9u2z8LnlCo/6vFGTYwm8mvkuXxoX175n
/LK5k2pZevz2vHzZ6VDyG6StkQqg27Eq3URWm1Kea16/Slqaom/Kch/Sc3UHZf8k
M56XBfWqW/Xm/OSOd85kdSMB69epXsGnfb7RoN5sUt1sEsX5rDjb77wW/p21RlpT
ttuxFx8GhOeLB06MTwmqhuPIBE37+so5QM54UuHP1jhmqGgTSNyJBtBR+yj7CnoK
nJTQClP0f4CABQxEcABY424s6NlbmXsBSaD0Z+KO8OgvA1efG6wZMiJEzrRmOPOW
3D3MeDVxMn1IQXkKx0rOaS7n49gC7O+mW8o1ZGuT0VOpijhN8l5sGTWj3Tq8ntfF
yPfazd4QHycPOjWh+BuNnqY5blW3YrbN1Q6mqIQGV15Z3lBiZzrte0zdAmZDvuzN
/tNY+U+FSzct3tIyPCK0O0fxZR9RVd031ydioQU4KO33VoNKWR9h3vx9VC1UZ38k
anya6rasDcxQWA7DMvfQ/ImGjm9AfUyB6uyPion+new=
`protect END_PROTECTED
