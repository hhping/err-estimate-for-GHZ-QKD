`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfehBdlTt8UhqJsHX9oiX6W1j/y7j1ZPNgXZhl8AkXjboCmWj/U3UQig+fGCtPmy
5ruF+P6F6LA9JuXbypRqy4ZhK4C8SN04RiPSO/yuJfWXgH5+JtM2pyG42Az9IC6x
QUJvizevwX5dbKELdmrMEooTud8A8PrzMqOeKl0NwpqxZ3kLWVRU9PYDToupXkVJ
bjfkGSiR0yN9UUgLiQVPa9/+/JQUyIAYZcVUMjnVltOCKfdSolNvD3R+9jq7I6Ju
GIYXSHjXTfFfdRurVoPI6Lt2WdyncnhczpW/bCk8zV9Wzb5GjS/dd98Oamnv8VWG
jRKZx1ykeypsqlo8RKws4gUpgkDS0dZg82PeLuXqiCA06tr8fOTj/iHThSnFcmgD
0Ihbn1u+AgkmR7Pjdl8imNPX8+MT/5ZNl9BdPcJgaegEX5n+lh3BznlZPF9HAMjF
Cm9NQ9/7MqBqK05fKs28XbWAXaC5lEsYVfLwwOL8zdKxSgUP0fsBR2Qi6Y32wkdP
PB8isWvsrMmQ7+j0/LUH99Ck+bTKLm/1cxxK6WcQrjopMJIqpfqoKEL9To53o8Xo
ou48MdELIoGP+lHq7v9xw41RaQYQPGGcr/DBtHtJv+wTRyYlE/emD7L8FB6Lw1Ze
CYUtunizUHg/RicFl89LDXoobTpEAATqnIhuin482SZ2l75Ixt69SYfajnumYWCr
0boXeWmsF0uYvjaFs9OiIC3qL9kGzuDzQs0RDsxjQ2evG+08V2HqVkvB+A0cm0Bt
TnhH7dJqxe7ATdkWY9M6PtlQYjU1DJHcxNmG+LQfMS8e7cvvKgRhq8zPy8RtAX8J
1Q15dV1r3Yqnn3hPAaVZAnVo4YhJSlBw0hnvr4vv0/1UKM1Q0ulhiRsRgyeRzvfV
nVrUFgTySIinZkpp1+u/yD42OQd0p2GeACfiurQpLn6iGJVvrj5k81H4bF8BlHZ3
yrpxrHFQ3rMRa8xEsEJ6jDW4fAZ1q/TR1DbeqEnSqfACXqoZvE8shjnEccswYKCW
9w0LqfV47Tf2JmGGF2zNH+9LLJlQqCHrqCmqQ0iMG35G2Wtv9FucNJolnDvthcU6
o4KBmzuXAqMTDkKW2t/nWSQFnN2n08++R7UYgQoufLiIYvVqQspH+h/B7ko819m1
DBYONdb29mesLcIKJ8NY46Cqk7AyCi4hJUeoiboiZ0y6LwzgHfZR9o3LWdEdoe70
8WkQAabTSxSTmlvQaxpcfl7nHkjQfM0xW+EZGyMNQ32f2yOlKwI/+1ELbsURIiZJ
2u19RRJFJTZnDAOgyJiwN0kPw/WFdUEaToudrAqsANf0jJtm7EDGazibmc2IQR9u
oXpT4AVE5OPnTq4FYDuG8d1gy347AlwJq/WD9ob1e64UKLC/L1Cdgw+pY33EvUtP
IPdo7cX2GSwbF46sA2hqLx3U4g4vLrFm3D+9SWR37tbmtJ/oxCnYmflvIUkfb9qr
7CJhzAnZxC0lxt2e09KcOdVBpsKZEmj4XlOfzZOii6E6E39JBQtA/ncj/AmA4jpj
g8DKWINXNHG0bIl+p4Hd3HnZPG22JMCsC7oJBObxeI5sZuVcK0Rjwwqeaz64wIAi
Yhf1pSsblKLAVRU19oFAnYlcLnjKDNe/h+7c+wwB3DXL/y/soPX9MiqQjId54G+f
EJZA/urc792KuGa+S28OwsPxAmfEP1wW/hJsumTY00ivJ2YyA3oIG8phEH0ytUEl
A0kS0iY6IAvsUJX6C5uHf2HxlCJt19c2mYp5owkQyirm5yO969OEh3t52p/wILRt
A3rNdL2J6Vm6p0wrpsC7jRGuImjvZyXLf56F2qPz7FbOs3C7y00gIg7Lshxa9PKP
XxHFJFsH5HAKulWwcEIJltpIhrEMAOXUH0JjjW95Whj7WKmQ93LClLn7ylUzfK59
2oWqOrx1VsvLTVX7wOhw0+r184FXv8w8SKU1779BJlIfkx+03XqgVTvXjvou6CZY
E7Uy4DHeGqkRrooXj5BTc+IAHUouJOCD/Xv05qBrjwKpggLTpX1ZuuMOOHnpwHpC
Yca9I9YL8bR52xjdTNDIHzNaYUvVbXmqaOuQaCbTIOrSkwQU0wI+4AqkVC8UKkw8
O2JvGD85IbHie2xPHrGX+avPWFW/VyIgNnDms+9C9KeOl5gd8aVpYU7zXpE/S38U
22/5kj0YGO5xiVoaWOgHm0mhsNYnAY69GdUBuzRKusWeDZpnfQlBbBZ49yF6RuQR
6d/RCLdwjiUKasWznRQnIjWcHcAz3a5ycGqUSpooo2PQxBJ3kAWbw2uZkQ9SbS4m
VfJsnQYqdLMIp1qgRIlyS8OFe88kmck5b+FwqiFIJyFB5EbsWMRoG0q7C43T7dSv
EaNeedojgdEwjXqfJl/f+5Dqep4LVWhurKVlubmLY8eSpIF9EueXpPEyrX+qMTne
QnbrWoliS/m7Af355HVu+VqE9+hO9DP+RzT+AXxffB4iyDdV3JUad2n9Of6WI/0y
hiUb0D7cZZdhQZ7vLzJpjtjJN6aN8V+zDlnJegzg37H+RSV5NJW/l4VxEJeEanrw
3iSHy1tLVozI00L/Dqjsthcv0lmi9cFWiEkpgPZKCJRwGAE/vIuKWD4td0+JBsfI
nPm7X1V31Sxy9RiI1K1qK74V6Fe8dzX5ED1m5WZlDDKjo/vrrYKZhdWPU57FYYkK
vyCofLFtUnc2S5slwiLgEqdsSGU3ftoR+1BJ1gzLEd7S3tBBkDwhM69PeihIH23N
yncPSEdIkLzq8SF1uWiBas5Lx9262hy5qHan+Y0wL7VlDrkj+4xfg3piJHPkz5kw
/n7puU+dNKS0tAaVcqZwK2pk1cwekXOvNKGdLmDB09vTpjIY2l2hF6Rma+ERdvto
VddTAr6y8kJ2zdmYzRJvaXz0huJ07J8r10ZxoFT5LbXpOGcvDqAxTGN5qqVPFPZf
k9gNpjAQPpujitibuLrrS31J5lwJjDagcUa+tBWiFnjdoeKSVrwozerfs/hravtv
v7yCMhJBca6lvM0EOjwyMg3kkc0myY3vVTzVYUrslizxHh1oh8EDlQmQs28XeMPE
ShZwdHMx4PGq+EHLmrvWtao/AGZaBvtNcwU0Uh/8QQNd8SWhYpdebAdprILEz2uo
eQMhDo931Ttmtz3FnyryMN3iLjQrAOjJkcv7LjLZjSNBz1OMlB5Eglx3qgKe97bk
sKHdWWrxkAUvfzwevaWl7jfOGgZYndHXqvjw9RENyVOHGU+7oOoErhD+/SQvDIb1
fZQhXRi1RYoz7ucTO7Pro/KebATJRXhykLh1ObB3kHjR9mhjLxntty8a3GO8oLq/
f10Gg3ltvOMSuq2ew7KjmirBsqIXgGhidkjZDxvA5Gjs40g9vXCw3zH/xGRYzKk4
pcJvmklM0nXaeWlIc/28SFM4x/Tz0OuGBewHimZlsHxPfmtn5LQwJnMfGo+ehoag
lRau/wKn5sZAGPH1jI7Lz3++SUMisg3MUPGhMDn+LJwUtIsw9VmFyKMwVXXMr8x9
GTvorsEHzjXYmZAGJrS/HwMRU8IrXBm1cmzOy3qQcPx7YVwhZDKlfmB93jc/zazE
3ax9E/Vsi/qL80tani9RuoXKaMu/D9w9WC2VenwMvPqJNkRZVhTcuyEP+F1W5ozn
yhXu4a5y1C4SaCHs4QnKdwW+dHGnnzWJGC+7EW+T+PWyIzwMsDdu3gmNrVZiMtcT
Usw4flb6SxmZmDJPqkaoV/kcWhnY/OKaUcAvVBbaSvmIypLv6bfmNyh91bLjS+T6
mMMtN6Z/ZBXLEdhDl4fGsAwJQmXPsg40ebjtSIxqFg/wg07iKHmbxjYLSPWUjTu6
KyA+rozrMIdH+/EETtjAlRURrRwIEKLqG+jUNBI/WWk3PJU5fCK/tLHMj1CC+t0Y
N/O6TGeMbOSO8UEhrRk1FMTZIWtKSdHxkJJte1Q2FuCt6d8lKidDpgX2azRoinyR
Ym7PW4MuhNRxAUTd8e/ZfTMFMXl9FgkzzAoWTgZdRZhzBwqhd5PJ/oNNYANlVlAv
dme9VuRKB0y9es9Z+KbL1NlIbqSbFYmDqqzDNx+YpvGm7JYcAqB0MsWbcnU109Yo
39sVTDLNbsVcPTi8ki0QUlOUT4ZMuXRELqxpkGbHRykpAYs71cXhxbRrMEvndFux
vEIVmWnX7PbnZ/KGdGE9hkQs+N1hQmGTv2/I0L5eR7bRwYl4ZqFXLWoPxN9ufsFy
sTC4P8CI+Iv8mL/17/HXYe+dIOXMfERd+TXcAl22XT+YhZcA+s+tB7I/O9KDzVM0
jBc6TpkLTVqFjVQviyqIRpmq4KFdvR7l5JohJc1NA+/cJh4aJUPqQ+rCDfeXdjSu
mTKDdvJnENiO0+2Z7xBAw6bNezA9TY4WnoSbWjYmY+Y97bd4f31LQpjXD6DGGobE
yv7BGfV17TVb/9pjnnSUDBCozSY2Y4jzFEhWPnXbRxfJTXH45/vBJvryUVPXfhoB
1/bBzpz4qCFEf9NpIwmDZFmdpSBzIXviuW1BqyKwf6KGvDZKsvvTEdEPmHvvfA6e
8fZbC2oOo5jROu8e5OxcVS5Z4khe2rytsDAuPGUPI1q13f6lbu1YLy+M7xOO6726
L0UJqLCoobUXJo83nqcNtRT+bSCMxq99j/E6QFBZ08Vurv+B1zrRvVQJ3ytR3NH6
Wr68eFsskJBBkr9ZIvDTVD/8Cx2NsqTaHlCrjnXdnxcc5fUl6Y+6afSeEb7Y5mWp
UZAKRwLiQ0u5EpIiO/XVd/fsYkHY/8KDtWG8AyF+QGK1t6d9E4+cK516wLfqUv7A
5NW/D8C7KGm58A2PasnGKAnXB4vPVrn6JpZap6HE/vn6PctPQiXWgZicsa6f2fJi
sSvFYdfUowZgG5/JuwcRpaICS1sFTUpdQC1mnrXzGGOuBXlNhQl1rFOfDTQRKdu6
o1NI3WZtHptC+33VpmZQu38qDcJ0xNapc2fcQx4h/6YC1u36azUsdq1QDQ9BidmI
0LLVVyUGMVNSmdAGaigWk0hq0d9ZETy0egXKM/xupmz93gX4xM8zXmc9Q5dfIcTF
hIjOAxIcXp1UXnmhgDrva0Sdck6uIXNXNdy4buZWqoTV0pJ+DDkGhToW1RtSmzoe
VNzH56SEuR0bV8aCK6QO17s7PK+Yc/7RkG1KulioKS/z+OlYnfG5jQrcVytK95Uk
bZOoeJk9ppwoP+SoEQ2/iLwNzFCGN4ZRcy8xUfBPePZkVaqWMamFSCwHLfIJpXid
OPGWkPPUIA/hBuk/MfFfWmeKYGgr3Mk9ssaZSPPGP3A8jH0vJs/sLoDqDDvrVIq6
YUdJFt99Xg3ld/ix2/lW2d7bJAXQR3M588foUPLgHtUJ11sqEfr3JYU8bkzbMvce
Zp0cz/tW3X4SNw+jF3dC6oDTN861/jSnb9QuBAlk0f7DzlV/dEiV4cl6r9XQnOUK
4FvjPE+x/RtyIiMhTzo2D32Zbe36QB3aur4teIX4VSZbifZPEy7n7tlncPuekkm8
dJ/06B7KGztZfReZlNVCZNYwn3C6Z8DzPZBbCSKAMV2igW8JacShDJppJZdw9WIO
JcOhncHTwx5sa/eIfAJWqRiw4cI+Eb9jlzjQpuD/ChGpIWHdRU2e5Nm8iCn3FNoM
Fo1yYXlB6/efcmc9VmNl6axx2SyY8wkQ2XP5GgZR4f/ZaRZb8WSQRTMEeMfgc3Bl
NpBHCJQD48Fbn+KFIbfHsZk4VyMFwvBKC4fRJJ4XdKh+2/GHbbXQ7KfqDG6AOM+3
JxrTZ/PB/zge5bdER8odMpJCJG1JXEpXEtrpZ+lZ3RaaQI2bNmdSCA/7QCcrR6W7
M2DDVAK6IG+1M+TnC1GHE/6xQZaDt8kxn2An2ekPovGTXo60wqtbf0WwL10T6BnN
hvqZxyO2c4TOHCSgFAZCDsJZZ/r54qA9fmAe/4q4WeULN4x0ofoKC8WZjhhPck7c
hi5kjdmVhEUpfRB635paF65DXjWS2pYMRplK2PyCbgnKWAm8T7fmGn5dl/geoy4E
VLnTqL6k3mIzO+dhDk3SiWwLW3y51eF19o6xzCOtPmfGdRHsdchH3fK0vqOCnudE
4kky12IChkY18dhxY/OAZ0yZc3Q+ik9fiexnrPVUelzcOuiT05sJvRpH/6cr9WWc
SAFFj8ZVZ0m9KUyIV0Rzih2Gm7bC9gr1YPgh/JTymJZ79xnena8to7ceIJCN3yzv
LrC0umeGxC6LDsGt1BwofD87ymt9cH+IQ37FZ0xkdLf7B/RBvUW8WO5C6R8oWhqn
mC7g268dPwhB5hSJbZCNO4LLjuIbIqsJIazegGMcFf8HDwc8h5/C2B2Y5z4rXO6Y
rC4zNyIb9vmKeh8JYD/Kq/teP3I+JeUlXKgRLXvhqFZMX7czQRrYPJo8cN8mCb4v
5/PMltb2nI64pdwy/48HCvPsT+ylygrI80yMZ8MtYWqY9yKccHZ9UjD6pPLE5hpd
VMdnViFsJgrARUfyKjwdYw==
`protect END_PROTECTED
