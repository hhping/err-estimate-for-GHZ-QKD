`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FybhPwpUZDcKu3vL6uTAF97rTqKUv+99UyUnf15VtLAx9w5funMU7W9sCUeA2hts
pOJ6+LudhEWCAi5gPVTUX7HMH/KRhuLSY3YQ5UMaJLSytpTorbLxp1wBMEe+oRh+
oYpJ0sAa4spC+CG36Wakf3QGLhNWCigiDcxIsOH855wlrmQKQnEx/RzV3EbBIGeB
Opta5+pA9IU/2GD+vLFlzvW9iOrVq7kfsmUbDpxE87OpI5urBNc+8x49taGhDnMo
LAJU0oEllW3gS7MAYTpOpJwTV2CVDtGq4Gkw9JbwZqKizTmQj6ARhwbeICGpklCd
PIyKe91t+zHVjydzwS6Vhe1hOOG0xkHPktRGSgFSrT08PqAw/d35BTm7psOOtmg0
bpWHC8aftIL5p8BEEfRxlZ6I4qcWvgzcXszwBKDWUAHBpG7vzjDrhe6vWCvnbgN1
lnlUxWzbNTtdhRycPtngJhdhak1KgydpVjBWundekQnpZCVzwLGiHoYeTAmBDWsN
jRhNd+eaE7x5bnrt72AUOM9DIk6edzoHNs7AmOSujBRA2wDGaI0rAS9wm10lFfha
G5mFPQAm7yK1xQiK4A53klwI4YWaBFEfywx+2ExLj6ywFQcIt2qNNgA2+3973mE8
GNKV3pEqaBCjFZ4jHemrsB2iNARJHHfrtHZlZTemInX7aHHI6hiR4YUk2Tx16dHZ
PsavJGg1pvu84WJdG68C0RB6DuWS0oAxyXEthWYpysFkT28tnMwUh0a81pkax6du
JjLprwtyyzHbZl7ud+x0pL8fmfONoaChaiwc5a5Am/LFMwkPcfo4+oqWr92+kbKm
cq4AQvNZuNvwICN43GagglcGBhwN54ozlB17rvwtr3ShqvNZNQpMFyqqew6mFHds
Ij9C/j6n13qiq5PlmeRf9QLV/z+NHiuc6PZNJIUYs2UQjthv9Xi0H/F6VV25k9ew
dSEGdCyC4wljK5nLVGNHy20EHeVaqvceD7xt4j31dWHlLIzCApZHd9NofJKG9L5I
G9/w9jY+nZIya45CdQOFsKJTnzNknqD/SdexjEqIdp6mm2XcSO6Gkg5xe+uhdERT
Bgy4n5XVCYldczcn2Nx21nA7AriFD5DtUiMvmKBeTZL3rjcoDC8QYoD2k8ifRXJN
wAImy/cSTMofGGK/8/LtQYP85w3UR1c/QLn2mdASDYVKpFtEPrcT60uA2WhaPZ8N
DTSxD6m3KRbJFZKJneSjnwiR/rjIMwgE4ve/OHMyYS1SfLLMtY2KHNbME3PFzakT
+muYwdG6NQLbhEZGuxEOjwufBUunwcZ1vcc/st0kSSJIxvZtdn0trU9zaEbj0qqK
tB4OrP0bZiqa8d9PVM0jmyeGE6UneGBHiM3nt/eByfUVsKi0mhqyLq01EbcfrgUR
dPlVmW/NVH+T+S4IUB3Xz7Y/lCSc+uvRwpr2eXaqIwnWW11C1SBKbEZu2d+CY2ta
jXjqYpZrlD25aB5+vau6a5aUNhUARdLRxyymnELMy0/1PgwTpZ2Xg98Qa6kkSzQK
W6Y5HyNEJDMMmGtlIrrhGMJ3meHPRa/ZgyWpfyR7vCST5eM67eT3OEfSXY7rnxFH
u3ShvWVMdKqsWGIb2Sd3LAg5Ajp8E6FjB7RDhQSvcyCtHFiWBr8LMI+U/xvZHZ0d
COBnZlpHVEY/zxi+zPHJJB6Nt42EEls86ly7+UepgWKU7BLMvxCfu6hWgboQ/KZl
lwzVgV9lf/ACH01Q6zm5dCXU9mKqVaU/I16PhwZsrVrml8r/FZeo03zZYnOCMgKB
A4V5ZXGs/V6Qw21NUVJlFrIroaoaCyM7ywGS7Vilnz8DobQo9c1jsZGD0+gPCKiC
0hMsc9xH6orRLEZ8wmzXqLS1VaGoL+JYIay6v5WlDS5SlghbWvHt9xKfTLncPUYv
PSHcOHWL+NwW6ySqH5YjiuLWcSsCjBXpRFT+hDXDej4lJJ4ND1cZawxgASjtPMBb
FadcIiKnSBt8XfTInTnsSOQwodezaAsSqWBV7VBnJl5jISVf2weEq833x4EQMYLd
yiBdq0pP4hb7eu5ew5dkbCdX2rVsq+o8xcT6U9iRcegiJpz+K83egOyXcIPsyuEw
5iA7Pwa6azRECQgr5TQIsm6CaHo4eBw1+RWTdH58jeISI+Cjc8gS8c/v/EKhFkKX
HsTpuLrddw7l9EAz6Qf5+LEKzVbP2gIMotSh4EArmrlGNQsHok3YwhORD3cK8Mix
8ZocVmk5UG9PSeLKoWSJCQ==
`protect END_PROTECTED
