`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mMzgiTPG3lDLNvkrc5qHcVSlOJzVgbpIIxyu86VYdHklX9oguYTI39WrrvnB9E+H
HEj9w5IjLsE4Qww4K+c9b1xhfFh7ih1ezLuLUYRKhCz/pgPdXIIBlyXZFPL8Xzf1
rS3kJi7OrGPOqEBmwxxe2JdrjlsAqcOrsj5/fnTjTBKtNEcpR0TS3soglIsS3TrH
6K2PuIEh2wfRtzowTTVupbyFvhh3lX1pD9ig1fUP9mSFuGSjiwuj27rZ9lGFcfWL
oSCH8PaJ0m0VqmxBhel9kbfNGmqYAGeT0SIMi4pBZeaSCWx/ThU6C9x5DlJ6F0wN
VO2Mje+MXAe7MnQc34Zu5km3OrU0zjlNooBpdK1b6mzCs9PvxNQCzzVoOG4x/I1k
`protect END_PROTECTED
