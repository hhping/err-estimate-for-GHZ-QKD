`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvHUIOeTmLNdEAf3VQy/jDyA7EobS0sE69IZzDjWfRdakDsv84TjD+MthZjjuU0z
RK5kKT78oa8RdEmGcTqdl1PSyYXIQo1tujKZoCdXzFQwQ7chGbKEOFjAbVrFoFmV
fIWpsPkCybtB9CrcayHJ4RTes/irlDpcVliipDG5VFM+qIy+LLF0fwTRKOW1DQ48
nTlWzQPyfPOMfV+G1NJ8LdH7zVATrGbIGdK79YTDm4WL09zCP1ntU14BuDdraZib
X29irzYGARikBGEj3BWX841aakEov3Yr9AxypqO4EbNszlhpKGTW8Fn5OcjmeZEI
7+PLWdeIkM9oWS5LNwJ2bMV9ctgVhfrBY+SoG53UYSSBI8Ufb58E8PdVM8JbwRkw
6auiFG+J2k2fjyA/mvNjYWCXTBqB1akQeYfXKEGbK6/ZxobeLzxP3KGGxHlRE+vS
mpImi1ABvjT3FX4SNo1lfJecDn+83S6v5gkR60oT6Yw/Sx6uOwpVdKq2l9Ou07T0
FzpYA3F0pDJgEAlLvUcrAGo//Nu9xplRRjSvBMLx7wZGCskyyejY20Vcr+82Z5XD
fC7rgxsCmBJcHnL97S31/CkUIkj+uBZ5yUegZGHj7vmWMlc9OsvpqeXGP+BqYocK
mj7jTz7VhFCu6dXJcw3taSKfOexoFsQvPCXhysC0x9XbRswHOoXcYcHv7mBrXz4d
OJ3TFxbW+hZ2c5jc2CCJLtj1HfooCfR36FM7EUrcNmacSbq+V+tsyOr2nMjkAacX
HWugHGurskfj8mKncRYRiMGdHZ16Ou8bA6o3uDu38pNA2AnN8exYIxXAF5DoStOa
Ib+4wA5JK8D1EI+4wNNuYdHj9Yle1La0TShx0m3cEKwdFR5LhuPw/XcAujjV48h5
NLautObGJIUHoby9cL9nYPO+pelnwnF9pE3hlqD4SBehuJYWAo1eqZhVdgwC8Ak5
YZ+W7WPDRfzbvOIrMxx5oWdC2pwtB5KkEjwcFkneBc2dKXp+MJ0Rhta/toAxUHaD
ee5hSnrjXKZjlMMr/8c1QMReb9DMN8tp7XbWyxAXVMHLLNjF80MHpsigMsbFvaAJ
COd5WXrMzk3iPb6WO2LeYFb2x/dGIoM7mt6Ugzdt8YpsOFpKoe7kjyMZW1elh3Zi
5rqofQuQqQ+mh35ATA83iOQLePJ3Vo8IVWJuuvbGDhpspTnpt6O/wzxBTjInvl/j
Ii7v0egatoJi3XWUbR+Kg8uhn8rx4Pr8zQGdIAd0F2Ri52GC4hWISD23JgPyhOB1
PMUJU4pLBHg0nhE3xp9o+6yvM7A0Z15FBRnMN6E1aBZk3LnWTAExknQcqtpsrbIP
V9/MTujqEZAYu7UlH3bO/pdDTqpGtDWUauHc2OUdwD/T59vlqa43QROBHKiRxzWL
KW/9fy2GFPbroXQDnbR3JyexHbHCFU9gMEjClxAS5y9HxhxtQ+yD2wAg86WvH8T4
r4ydKJEvdSc1qgD3EJ/Wn/tP/dg3RVuXkG542Tb6S97z1e2ZcPOyNMG0UXt8grxc
mxAI6JhtrRj5+HvRaZQwpkUny0/Tx4DY/jEzmBQmU7Wt80i4lU/p0eZzX5vfPt81
asRa1JIgHAyvoGPDtJv7dFD6q/MKGTfscGjB7lieti/YKJK8EaN8nhMuAiyu0gW4
8uoIuyz1wcIE9GE4LF0P8GNqYMoilsbF2blF9b/qzMyo94Ba9GTsdpeNQ/oHM/el
bp3TPihw0Kk+rjZh6dUEWfmvzgNiN75d2M7XbF6ysDPAGNDZ/lMRDvqIIXozJo6I
sli3++48Paw5WkiHStmxkjrEwU5tak2vufOAKwF1kbDlQoQEd/TgEAZ5LEoUvGmO
pRm/xuBQBz7dvhRhYx2vKds3afOnBbmzwc6O0I0ll93UybJsM/xRXQT3yX+AFKqC
xnMtXPqXPBIrfo97Ovp623kpZ/DWRAW+Z5siAa09/Ai8GXapP4YkpsshDf2/bNdD
1QXwwkIfI3LCqvP/hDmJIe0Mo9al1wfD1+Pl089khuBYljwlBOFoBFpBqVK/41Fs
0N5SDHm2Th9/4Uv1rAH00fx3lspC8YWelOpEprEBXivhkwWmt0Dj+ccCNh38XRSV
f9BZA9nD+i7b5AKucoOQe8/GdeXXK/zFeI7Zd2q+UEsqZbTpRAWTJEmuYku/tU1x
Du6Y4EXyGFkDHneHX+2GdgdyaE7ScF3wpmyJTsVvbdtSrbmNg1ZhCQJhrseFXntW
6GRsOnpasCH7JVmFd+S7SLXlDLymWVQG0BuE+pIh2kTkC5pDfgqKEj5vFWsPRtjw
moLuO6G+rEfo3lTklOupCrT0+NqW852T4xUiNcsIEs2vEcUU/F3KK+3sFGtFQ7d4
+vREytW+3qS5e9+wpqqrqmSCruJP5XuMfERRCyjUTRhQB8ltbGUqtJuVNmaxGqFx
vz1gZyWoOmifYfE7blk2TluvdYGzcDcaqFMnS0ZLRkodtTwnO/7VLaOrnrILLMkT
+F7eSUDlhDq2SSXz+2X4k7jYgaTwpbLJbekcvLh0WuNvPvZpny85/bdNYbQQlJb2
ukAaX0re77y/L8c//OJhklgnsLFkhOeIJLqUS8Zq6Go/EkKuHdvumUGbLU5BapTu
at5DZnown4du0FBJbpUhEzABGxiBTDFTpiGeLVYuFmX9HqIUxN76HCLAP3pDaJ2w
d/mawnZ3YYk9jELjB9W2tSQ7CPgAUoKWpYwjYc73GKWWi4hhFmXr9x9Aah9Cg5Sr
QV8gfLjyLgCMOB6QXFJnrnBCa3j2uOsQ9xekoRGAKU1QOwOIil7Qtnc1/28aIG5S
FenvO6J4fNzQEtUzg7AL2G9ELT4wPbHyUoSfqp0MTVlFyQAZ9TYvwEXvRgzXgvRc
6tj8t655arzscUL/JT0R2FtjEgWpGAOpy610HZzcKMwmfThEOUcKFVPQJvyCAmwn
83+32iV42cqgScTYaJFy/USZv59krIgwxrYw+qFUH7mqcWpzcSk6aMN0oGrvzk9T
688nf5vsswVxoDCblbiUIVcVz+fmw9gQRntnMX/ZKUgwKS73dtGC6WYWclLVLSCo
YklQAJCxnKuvyGYUNuWzKyOnJNQ8QTrvvhzWE5/RS+srKlL+2Uoj7iS6U9IwZIVs
s0+Du6cmo44THlseCemA7nQBPkRY4agY9dgiTfM9heoiEth8695z9DGt4V+2UEO5
lhO13X6r/X1wEljCG4bO2HYgaLq88q7dMnqMdcKAzp8TVfKT0Kynnyl7eEHX24s0
`protect END_PROTECTED
