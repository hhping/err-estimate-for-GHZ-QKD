`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rmqqSuM/eAh2cqBtVgsE+z2n4+aF8gToT7/yb/BWfMtA3jgOvcMxCkxkQ245IqoK
YhISbfTtT/ousVpDw/I0I/STIrjbl37dBN5GhqcAf7K70tHagaVylXEHgPLnVH6O
zxgiTKnkuOhZI5sE6kKSeiU+wuZAFYkryPs5DMq140Y5rlc22wpcqTmhb+3IjvZS
rNqJ1R1fei6YtPAA3YPGpnr/evChKwnbP36wt8NPlSP75iI2aXrFgAJNVWLO1XIk
9bHGS7b2eAeKadhPrhrncMEihJOMn/laUC8g8TKKLVKOLG5ih3I0Vv6yOP5DC/oS
geh/SV4JFLlvjPscV9ud9Dzzg8EnwldZA/dvOsI1TPOqB2oYc6UJsbqmgDfcuQUv
t2IYgFuGoSFFbNv4B0gsXzhkMKYQonMuI5VwteZXjKotHk/lmUtvkfPzgEPP28kQ
IDt5aRqCg3ghRcSabNVMZ3wwTzHM2bSsP8lAEGUIJox/vhbICAbY+8zCptCIKLjo
F6t1F3L0OK+oygvpfaxHHO0Rt9CwkpDJFaYjj6+lQXLqcP5BX4Kh2JzRvi3viEHa
kIGDRuediqOSo+3Sy+lab4+yQrxx8cKx/WVrpkdz1ID4768ydMTz5N0jrCM3X6wi
uFMv9OGivZsnIJXDYEDbkwaWmInDG52RzGZBnADQvlvtxugahw199K51nfSS0sPa
k4Odyrvuu90PZwjWc0f+HqC3mD2wS2tr27zCg4VQs0NihqvrkArScSQBR6DJyva6
2z+fRNkfYEaZBzcgx1BmhOQfuYYn3CQBLRI+uzKywlVmTNr5gOBYt2ye8Oqvut85
YjG/g9Hf88J2fa9RXlwxddKvkWKC6pm4hl9EKOHyUvB6wF82DO8x3K1kOLbcf35r
uxsH6BY0oq0sFLRudHfPXJPm40HWcXcT8e+FMUTq+cTxhd7jILbg4I9cTxx5/n5L
X8xzhXfd0qLHsikY+5eoXKXYm/DS74MgI3VMqgiGPZYcFva3OaHZ7ivEZGKu2fCC
O6iKXAgs+pWQbjxbLMAzdA==
`protect END_PROTECTED
