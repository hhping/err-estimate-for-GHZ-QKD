`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIMGZo25u6gpPkNsXVhhf8hJtIuLYXt/8piJ2cCIQIjGMTlIADiVe6iKtRZWLsVl
3WrWhIRjkh0RrGVeOyD2xOLP3xuHvMA28KT0X3epx4EoCThOmrPlZfw15xyeCluF
tq9OxKN8JS8Ka15G7HzaHNfgrLhHf/hoiwxiElHCGm90m+xaYZSR844KNxY3kVxE
zSQCm3SFR6LAqkPaZNYAq1HlD7Ft1/Xvc9tfV+zVSt1hVxn+z2UbBc5LQVHPuSD1
nNrhZ+lsynmnSHC8TeYPIqsLcypLuxIQ3RgkeRaRSCsBsHc5moJkjd+97U3/LmH8
LtToL5Lg8bgV0eHsdqi9rHaISIldJj7AAqoeHlIaCLi62CLDlKyIIu0T3jtkNkKL
dUZj4r7Unn+bO153iWtRC2xydkM9VIxmTOb2zOlXa3ci1d1MZS4sTVq7NwdgeCl3
1Pqppt08JVcINFxZNW9reEh4G8VmrZ4aAtGeY4UqOCqDh4831rvrdLPJdudNhRx/
DvRZIjh2hojm5hu3gIgRfq5AsgLk3DrLiIXXXUTgvOjMtGLuhHvVX1Zyax0Xxd8U
NtMOI3Wl+0DV13Y62WpOZbu3whx9AAzIaw72PFlxVx358mpTeWRopDNA8+qUPiKt
sL2xzeL/qBRyvxWHKirHrQErC5w23JiCkb38cnSmmDvQ/xj5Q3RleS//C3WSXUv3
MGp+p2w87wxSIdLKieBVNSNFNAL6n2t+5BMJRPl9f7hyGLfL46dIgfl7riChl5lF
tV191W/iXqHfvITA/AF5ho6ahBIK8TscFiWmmLhTu3kCK7oKPdFFU86k8vqjI1LP
hUlSs93keGjrFIt6X45r4MKzsog/2OjpzGvlmLgdCX8dS6Ifxgx6n3up86RHLQDE
h1MNI0shZybQslP9v+vC3lk6gBb3bho0gZcQGFePRIU8t5V4mfWiMwZ34tav72Ya
myHPN8cOD3lwAYnNeEZzQeKor+CIBjaW6rsZGwxT2/d1FXKSs26SlYvQvUY+Z59m
aILhxog+vMVAIzEv0enERzjK9ARWyzR39o6SAzxD40o=
`protect END_PROTECTED
