`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PyT2veafzQgyVUGYmMWC/5v0Wbf5qKJCtHd1USkMk+nT8VSNxCqIb+PQwVa/po8
kas1sW9AKsvy8uu24FBr5IMbvkcVBU+ulGru7tRhi+/oLgxWhNUKhOUnrVLxDuwY
NOBpEuCvcYODc2YlVTQPucSFcffw8H/6Nx7QAyVtlIQmYJIIXjSIcdF4rkelAtDE
xIvqtnzGrk3+Pqp8XGL+Z9fuB279SC1MEb2p3xymVrYpKSBgr/GfFr35JfYLYhA0
l+gh7nNPfmTuScoZ48q7Al66/RgFQt+XmfMDExMwcqrNvfw6IcnkDybQxIzpAU10
LwSFRm6z/nE5A7TwDdwJ+iLSZJVu5O3isKXu9k5fjsyKIh2drkuJ1zHxTk8AiFZm
Tru9d74hzazbML3jtU+T/MLdPalTjFyEoeITpsZdOR+LFA2oLq4xyilrucNmaZQ+
dGYPuYcTUmlneS3opTpCZxUulVevWCXR7RZC5x40SRlgth66tB1+2E2tpEDaoeUX
0uTKarujKw3Mrkg6IywlB5PDvLnbGYcJi5A6Op+6q46Yzs2XDurt/FrzOjrKD3ud
dNvHdTJoJpPSA8NeD8BLlM3hRC8w8xS3uLN+ltoG6DkkztYdV4wz05375nz05556
+yDz+qnLm/x/vVE7kwjJXSYvAnM80Zt/G8cb+aT7GrUtKuPdq1uYMkUizcWpCeUt
39U9RLDfgyravs6HJlWWST2VzcfTQIkm8zZxNzJ4sJEjPT/QE0FUQXjIwhNZNhij
OpdlsIRrfypVMRfG6D57w5IDRxV+DbQ8s6cRe/EBKxlPT1m3Kk8QXMB9zsbKW4cD
gOt2IR9jQ/WFCFvNbJz8B9dHXVg1ZDUkWZtVihIOpXVNKY1P7EOt1iMe1TuVwQcx
Zvug7q27AcTlUVrIVtD2Qi5fhGHXdY6AqKV4q6cdb0x9w3AEeVSbGpjZ2fYBw2E1
rwc4sdVGLn4iOgKDHl/IXmCFvQVSy3edYsNtIp/0NsN7OVFLZkx4TXp5vbZuz7g8
khgZYEKLgdDdvb6f8t7h241NpGkpD/TpLAol2keOM0X8QAaH02T//BI6Shg0/0gS
dFWDnifQC4xi2KkhNDyR9Qt4dLExpfLNM2CQKKGGXDdli42E7ycPCer/hfXoe1sF
B1jmWmJW5QOGYUKp7dpelPouhxA8D2zbFcJiNs5nM0HcSHFzVp57CluEpljU05pv
OBZBxRMglD4fZIki7obIkAplub8c9gOVPpnhIHQvxNfgzb3mcjuLj8CE7ow/Q74T
M5tHXwnmOQkObS05pWx+oSuPtnBo2eP2P22FbW9faMwiKjnWC5/tBaMDTKktksM5
/1HsnK71VlCX0XMRbJyzy4kdyctXWNviyDJK7k4K7FGy8Uh82SzSNy2cM6J1mMYg
/6bVSNoeK1swkTgYMfQ84MatGxSCxESQm95CU0T4x6QE+1CpLRdG5NNrEjPcoVED
HCG9evNPCdWzQjHrLbDr3tbolMIAldUGx56KU0qTM2f+MlAhePCDrCT41Qx7Fqs6
RSEgKTOl27sRf3d949x87PK8Z5jn9Mw9KvMOV6D7rth+jh91LT/D1JC2mYZObf91
NZ82tweJ9Az7beJTUgW1pQyJW7rrlo4gRCn/it8wFXi/ga3GjS1TeDJt9Fv3quML
htsZDqysPsGOIQ0ovMgAoyw1iEl/aUYIT9l3OFi+fgcwm5sDdGbZaQj4xDjVawFp
zqKMRJCmCbkxXhNi6GzxnIaLJLkInd+Tq70qyGBqswStMdyCmbKNhzkujZ8wxztf
EOt3zj6DiNHlwzkqQvkvcDITVvP/HYaGYheUjEHyNSpHj8dmNcYGqClOleSxSwCV
3bXXXnmge5kruEbn9IeYhA==
`protect END_PROTECTED
