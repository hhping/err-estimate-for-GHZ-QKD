`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/WWE3yesVQWdXDMh6/V+5L9f3Cu8Ek30/Agwe58l7v5gJCVO1ohAKzTm4imbY1Q
0rJTIbl9+JoygEGuTNu+CRI96+rcEqq//p3IDsuxxgS1EuMRSdSnIriX5M2D1rq1
NwICFjnZWqtpMG8mB+VGQT62hcsjJ1IMXaVbwf/5FmH8EB2eJtuZgO/hrOCHvC5I
+ZJ1gF6EYeFKfWFkoGL3mS7O1qfrJl7wTjhBZY7YBjmmvaiutUd0pGUqf4NXj2qY
U6I+X17J6g9gYbLSqSAc8Ok2iVdoIzItNmK9h6zgWC39Ja9j9mGN4ZLYEvwlK8vC
5i7568/LnIjxC5RAG3e7ltx9fb/ToMIG9ZH3MkAbnE0GsRKbiBTLiqet8gKDQo4c
PuKghldXYGSaESHwUaDeHP0NMOoxzOVIKA8ecjFXy9AJb1qrWFI6B+2dg/BvVd1A
KCRfwJAAi5C2owa2P5Xzqqifzxqa+Y0E3xmW67KWjUIT78pkUOxqGhqlg5by/02E
07fgJwGvUSsjZ3d4gJoDXXqhef9brYJs8SkBmKyc/jdwcJ/FfSrBr3p4QcSzADx0
+pFrWyKeq2ujDksXwFth4cd4EGYApOWs4U1hw90IVrr/zvuMuimevBbNOx38bG4/
gu7sOfJzZugycFVkjm/48dOOxk92QxS6RiaD3stFDa0nuTReup8pWl1tzJJwzQKW
eO7FyFgzRuApQP0ywBPoc+dgcxzmf7GrybsE3+ZFEWpHRALIk0xFeI6USnZOKHGw
4uXconi2ZWZpUJr/9pFw87S3R+WeLYMxDleDpD/vGFQj9mITV4w7I91Xc9iuI8fR
RkFkxVJ5pVJP4YOOCKYT7WSweoY45jefSTg6pq4JYACX0E3UgVeVwh4jumoYL8yo
KmhjMphfYn6bTWi5s9rIaFyKqvHqWbhnaQ/DrFlHvnDK+r7pqP+PE43ipoKw7ekV
evC5tBhMs53+2/2gkrb6WQO5uKuYsct/RH35ZmWjlevSyjOdbcHuVh9rzs1fCvbK
84r4TcJDQ7cpXon2VC7D+CIo+FqO2GPoIML1xxJDXvTW6Ik/mtFEDdMIYjaT4jQo
iK+VF/PoeWq72X4B51Ldb01oD0mnkFcLZ5Cn1kw8+AZVYWH/I3Z5HC77SLsd81ah
bZq2UfqXbZcaL6a5z1Q0kw==
`protect END_PROTECTED
