`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZt1O9Gz57FPXmRFvsXOR4iiHArB4bR2RDa5JuA3t3ozzRVBXgjdls46RF9UJj/q
D8JIo+Uk8mAKHYmfck/0qTns5Y2YXzSuF3T1nEDhnVDODQ0ytVO6GT9kJR6qNlf2
PIXq121Wbs3ilunS8JEuEeSggxdGngDUFBiHr1uzuZXTevbRUqizk77Qg+o6ha7v
pw31s4Bon0N698g/9ZaiWTnFlG9VaLCMu3Rpc4NfcPjGs4KK2W7wRVYPZKIvwHVR
MBFU5vvcGmRgi9WUxi+X737C5czvHNDsu11cFPSPwxT1gOuwp2YFhe8lKLvQ2yOD
m22io0Oj9oa2MosgSqD6VBNHIZzYOoRE3pjIBwEZBV9j2hE36XclDoFfcDcKVeqf
ZA5jXBwc3wQM4fFn7+2Sx0YAotC+n1YxWamw6Vr9yyWKX+IkTcsQ7hLDZcsKK0yW
Ph7F10sVtoqNMwWWb7MuuD05cna41dBFKbZROedbzRTboBd24uQcp53cA3dYVoRW
UGb1zHmQkPPhMD3O32WjEgN0a9oaimqVCcaPtCtHnbdb0thYp3nk4BE8NruTI0Yv
+1d5aufZvxTPcDrRaN6o52tn6ZM0DN8VqO7yZFvu2OOD/UdoKk/fk7kj1Lcotyfj
5rqe7C/Z4qRDdc4qEz9cYUrbwZtqi18sxPZGKXzZedKpLHrG+IpjRyJchKLs4vbe
qHAuPRj/9XTVIKQVFHZXQaNq+SgVRXslaeeWA1HduT6Zu/SJHly9jY4K9WCtlU/w
F7vF711xqP2leHsQK5Xof+puPkTp5pc+VPFltRUR/oLpsGDeweP2+J1Fh9ERuQeI
t02GIgvwcmE34CiJR2Xe11cSl62HFdfLn4slg9PQNjlMy6SLRq28R9UUBa7J0Rdw
Rr95zV/dTrCckCZU0tK5PxrWlgt3fwoMYu/bi5pa3wE=
`protect END_PROTECTED
