`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luLqa7NW80eQKlSaMAYgDxrtw6kh3th/UbEZorOBeVAU6gTv8lKkKBW/qi/X70no
ZBUH+PQ0ZRNXCGZP0YpbOeI8p3e6OrA31IcbDICletvh1hCty2uL1UoMinWrrsIa
7uUv8qmA6yNEsrKoprbuNE8GidcyZAXMvO6Wb6RGQbLFrae8ykTlA55pHkBePPpw
mPu+vtNrFegl1yL1IztmKGAfjTaUuHbljAVfo2Xf/wB0OYHcMH6nkl2+b+pYewao
HDORLEpjZ/SXwAOSPtLyxlIeR5AepvIhkSokVYfZQXfKFKAR41icA6/wFAJW/gIk
IB2yYIeQxzaE5MRy+GibK8TNZX/CmAsh1C+LN1OHudGKC4tEZoZBSZiwbaykDT8R
dyXLz7CcAMCDFNDXP6VKJN25AkQ49aEuDIp5+HDRk5NQKu9DWkjBXNpBUh/sv40K
pC5hBI4CD9FQXN0Qv03YGDYAuehQYwL0eaDapSAaldR/hgM/g8ObNkXf9lnIUz62
R8hc5BB0LE1yFl7/nfMfpbBOS9FzBa0Xb0ic7/v/mTviExNjSm5CXaF6AOcpBXFI
eRQqUWSFICTpwGh4ZtmOJ2XsQMA1ly7AazC1yeCt3Odbe1S9EuXdlmAXgwD60MnB
Jf8XSBOBB1Qd31mYbTOq5oLhgXo+dP5RtbF+0Apa3y4WgcVs+YpfEFTycUEqhZLC
mCTzvsw6k+z1QOvF8ej5sOc0SFIZ5gI1Y01xIYmq2rdcYYgY1Vw3Mbw5C/yoTPS6
JBH5+AqvhGyud5uWsW4u54iZ5WOlNYWsGpvU1EZUNYVMVyt5ZzdyEmXV5T07Gatu
oyVamfKWxYMOnQ3HhGydEJFPMLzRe/9R00hgT0+j4R1mQg5S0Ht/G/SN4uZGlWVS
dxA01i7pUUm2gU4+k/Bt1+Gu6Z7nDG+Ay3f3wSeUW1NYCN2kAlBMa3gJ2DFKnU0F
smNZv84aS2POtFigspD/4UUxvSJHtmT6hiaRpjZi9Y2T6zr90oBnBP+3wS3M2DwU
upctUTWtLLP0O2EG/i6/Riqque0spetN042TSpZiKZhCdVIymCRAfhLj3eO/5A//
ONoMawp+jUGifezlSwX2yQ5N0LvS3P9nAA/ik/r7utjZjcAuhULaSn4NoFGrxD2S
BIfqGMzS4bbzAms6f9VTqHgIv5RTMLWPYo2ZgA0qOsrEBS2mQdCvlka+DfEk4v1U
qR6LEBxVmDqzNtkluy/8viR9MO2BvIZlUuWc0gNczD1OOSXKKah+yOfh4a43Ri5c
SIF3BpMHHUrLpp0E18maS4baEJwER/8VEiEJJJQjt8Zj0UTqExp6r4DUMsqPo6Z2
lNjIfeCXbN7nEcDfE08Y3uQRVx0sB/0tjxwZKUlxW76c+2yrxfBaQBAA9QitRyl7
iXko+w0YXItcnO1umv3pUQpezg2HduHRgvCwc9sfZo3LKQKT5XoPFegrNduFbmB2
devtBwhsDm+mcQlYEmRYVabupa+lrIp7yZBTSEBdDOVR7HOnpCR/HvTmXC1GM1Q3
Yv0WZaa8pmEo+yKoxH4gNVatiMUSuOQdvZfDmdrZ8zemDTLbbMUWsuyOBP/S39ls
eNCBAP7XGO38hBILMQI6HByKF0CCoCQtDSiuBhYBv6L4lpwoCMxJGhkshztL1l8X
mMV6IChDRxI+LGwzoXJ65u0z9eEZtjQi5btMWv1NJ0P8i+wFNYyRLwq64BDqmGWX
e7ce3O5DkM7OZAHVylUg0O9mEMp1BZdv+waImbWWVEGtMpa8DS0WnkJklgtgd9xT
w6ytY0KQrRFcoKyBalHeeQ12f8UsqIsTxQVYC9h7AP3y48ts4qMwVDT7tV4aOI03
rnSDHo2K0jeeNRO+ykvm/T/GhHPu7ALIXhjyMPErimT0YfWQhc4NwRWZlru2gTPG
Hs2AB3hvLdHTo1jVX+IiYmeMadA5Waim/iQg3zt9ZWW6bcz4dQhHzQQjd/lkjFmp
H2X3v+NjE1k7nEJM7tHLzTPX3A6DLjubwGfsMXjH5cOaJRNVlwT1Orwh2+5o6dH7
sUbIw8cgt9yWHl/Nbn3zOGHY3QRsW0t/RVvx8c4fMARo2FQtQ4jEvF4MCe5ZpX/k
PC6E222DR5eSofTIuKivBewBIHfzYNumgsqyVqtekR+nNTFoiXb6810QibYVJmsh
uuQ1kdmc+N1svgBdw9ZqydIcsHonKieUC4v8wEhsm/88wqAiRshO30Dq3qcJ0pxN
M7xwXmG5U0i0TYdufRJQn6OL9/AH1M8agJ7vP7q4TymLPBZar/arsEt/+E2RVsEu
guR2NpHvhzeUibRkRXpcR7xHVPytkHXoMzMWd7n9JtE+oPTfC6AOFrbkjF099UgG
Kevx0zaRenLuxQfwmWIYIyQ78/BFUYlzEH5UX9OitjMBKW+UGr//gJPs74GbvctM
Shc7EItcrwbIQtvjXjaRwF4LhNC76l8iVqlaEMfY8oe+2tr/+xpWWEGAGPgMNmii
BK9HYiaFyFCeGvjUY8Df94fgcB9B03hVsfjllIvlx6VvhOlvWlSSvG5EmZDFmEnN
ZasZP0GOOYtaAmrW2GTV3xxt4tKLuG1kvJDxGvM2z0eKnO9ismj2kbkbVzr8TXQ7
imIPbNANMN20P15Fj9qrRD6ejpJfBmMxFc/1ozoJYYAESxTms0CIiaKqSi0MVGyK
daioPjCFnhohCr2sQZEVYq230ia8PTt9neDRCiOiZJUlacv+YvHby7/M+jIPQsB1
FC0xr/QhZB9lTBIgU/ICMC1SkU/7OBq9jb7+KJZ0PQbLvMBQzwJCOw4W6RHfiQny
YmyG38+ue1pJmw8BnrqGDsuyO2xJYT1rQpYOjkKg1GmKz30J5wk47SlRTh4Q5R98
fUCO1RIKdC5nyzBo61jlL7Qy5QFfsKYtFIm1u+ohw0UKUS7Me66IZ81YMJ0Kef7R
lli5nty1YCPVZqO0HuVoXJgcCtlE/wmuP+4deO6G4LhA1b+i/zlnCiKvHScnxMPu
RQW4UE70Bna3GMLyOF/+h9hkn441pAtBNVsVFaNmOvHhAU2ikw5qySEWVbG080DJ
J1B6y/f7aXMuODZyvS5QjTlcpkvwswwKOfaITMURBqXYjbrv2P5586dQWZ4cCWr7
slOH7cJmxFYWu3rMRKQcmlME4tWslSbcDnEJOpxyAdYRrb1JdPfkEVrxZQ2cTYGS
nJ0VfjSs1EIUcODwJLEdwH0GKG2DGufn+cW4nNu6PZYprD+ZLbxphu3GOmfDjp/6
lX7cZR8ltdxDESUQKDCqwtyCfAk/HVbzM1q4Ryo4jQPKPxx08+syxczxbQ6mLJGz
oRz+Z5QRaSQKP/kGxef8Rl1HHLR/lGqLA7+/qPdIasiTl6Z/Fe30iKxC0u+NRYlu
lxH2N7iNm6j9NynCLKm4imsQtTwTALr7RxicxbM0BXaUtQM0FnJadxDYe8lbv9vV
ZVD0JSZ2qmf/PL4OTSRXdpnY5qvw02JXy6KV5RAw81NDjP9JM5e1oRsf4j924P95
MxXk1hSDGEn+OSIolT7z8fHbYsKLoTQupy5UCerWLfJ8jvCbS+Kbv4d75EfMpHc+
kFdkAholQXk/D307yj4g+DvLra/dQNCoevLT4gOh303C6/iHTmWlRlh0E+p4h6w4
B6eXO1/q0bACHdDLNywMLtFzc6+n980rVwzvKEze6l1JRFL0hlYr8+m00uqskOeP
Y2vyyTF/+uFlXQdkiMAzaadsXMZa38naERuHA98Ntbbf2j4n6TaRSzhxgZ1xWOnf
a1M3h6Qh1g5ppMdoq1/v9CnXag+HHaTLKv4/pK9/GPoOI/hH5rtxQb5vXnvzO46e
zf0vuxg70ADes/318vYWL+NffqCU122hyCdIDzq5X+3F5PFSl9kp7JmUt3lkRo4e
5U6hsIUXs2U0QDCc+3PhLbeqtDMeyvcBwM5/qIpRn3/xAkG2dte/vBs9eVEQh2DF
ieW1n6fjv4veCDKxL6++HQFKKM88SiYM76S+cY+FyXXyob+uWvJjlpoEbhBN0OjD
fGYG+kCbduEzRgg5zpFvpnJdNxQpr7RLv6+LIiR5N5Z9or83q/xocP9062RlZV+Z
1+3HqGy7P+DhlHJGZvtVE/FpVPfsQLNHHI0FsfmNzPhhNfG4ngk/bUrNiOygARFv
g1uM9tu0o3Cyxzlak6Q47wvEavP0kdGt+0bMCwotRmUW8CpOi11TE/i/Mwb/HCVV
CgHAo7KRUHcvJ2odqKsybtG1U7w1vpSOm9b9//w0xaGHvYEXTeO0L/O0xWpApVBu
OujC0UeoIzcvFxLBqeRHfDZxo39MSe1cVJHz0WljZqGL0zFALgd3A6nv48AB67hi
w4rtk6yN2dBEomGn6PmDfKcIeCw1RKYD/tgjrs9IAGi/GfjTd7V5iguXOV/soEsR
QpYpPD18s5zvdtUmdK/Ps6l1V6Ih60tWHOvaqPkuxk3u/z0KJVic7sKkoan/2aBI
CLm1XRbYbvEWrX+Xu9rlKQag4+ed4Pv/3NhqxoKDxz7fqrGlXSz4xJ5rHeb5WjH3
ASrne4k2lTyj3+Gt+ZN2wxXPxVk5763DNpBcBz7cmoT6pj/zAh7lmEf+m5D325ZU
scir3DV2Y4n4uh7f+5YKK7DqcwqqV5AQYCPfffGCv/lt5H0F5UlBJz3ATL8N5krz
siIgwPg9crS/ddlPq/AVAfX+BvBkWGNHnWaNzp5bLmRIbpkfIMkn1L+hrMTqXFWC
UTldHhabNfx3Hqq/kTyQc1GbwrRdeQORQlEloQuIRXCNDFTKHVhTmmwXd9nHBFe7
aYiHwZbriuit/W4bgH1yqVfbf9lwZY6+USUTcsztqkojYtaLReNw6Wjno/WXgGFW
YCiWv7SotziwgmbfE3EqQAwYdO0EjJw7bLqAuB91j3ebzmDe+mj4iDNIGr/oX+cD
hiJ++cCsI9Uq1u2e9jJgOilZcbN5pF+VXcqBJxpCfntx6LjwzkvOd1i0fj4VQgyo
NEPR6z1A6RMnUb5D88d+DIwxU6v0wBSF50VDSEzAhbowuaaCRHZi3InpzscArxRI
tq17pZtYCGWxyYb+Ja9A3zDV40SZZjinlnqkSgEY7Dir3JG8qF0cTTh83h/JGzeN
kucqCRnZ4pN1/ctUom63m51aV0g/C2+Pv2cyXx6AqiWn9jM4q1T1sjXuKZ2h812+
rOShjlT4UXC4Cdk261ja8w6G3JNq/LYNqe+umHEbs34lRJBPzo+ZPOnn1enRLHpE
2MbFmBsL/d9MZkdVD7v0xRKW6h0Oal0p1OOmJTueYTizEkP4smenIG8TwAKyQYka
MBpE7hYPg9sEPTliyt6gMocz/w5XQkrRTkXIjYm8e+VWKml89QB/KR8BGP+9/X8E
5QsUW8YqgOH0dHMBYDG0A9jiIJxCkmauxk/clBQnG9YQqM9iDvwxi1OEEsUPg1Ca
i7s+Xdhpl/2VcyLDRRD2srV8Av4eTVDhzxoG0icMqAdJzCIJX05pH6Rt4vfKuoTt
K4XedGBBOfHG2miULngbQJ0eAnWcRnGbfH3RMgfyQ4fwdkjGYiS8NPYZxSk8kFGz
o1ZAP7fIq9T7+MlsyMiseA6YiKpUFmn9hKQA8koBzC0DpdO6Ak1okpYGoPhDcXKK
zVUKXF3/s2nv2V5fxMKLikQpW+fjWM3h0ohNvkYZmS1vyU7M3SZSvWjyxmYl34RH
TnTa7lgnqGBedT4eenPT7Klr7a0s+Ys53zBuYtApPINX1M6YGLzKBcfDLsapGxRD
aGVgTQ8VtOYbtQ/wbOFrYRU/VaVCH9OygQEO2osXJNuTIvqB6yiHZN1WZYs97Hvj
ukztw/HKcomIJVscjIqldXqOjttatnR+po4SortWwnxl8stl9i3vgh24cNXzivrj
7qxRnctUsEdvHhE+mLHurP6muJ1hFGcrsQP0dpcoZLsUhlxrCWgwyT2ATOS2duGT
rvtelgCdEY92HsNPvRK3JCXWnDN2JsJ5b/vILqGkTWD2O+tpgbsNXw5FYD0Hr9hN
THCR7XANhvBQ0M/GzkK6iZtTJPEhqtWAO2Z2C6bmsVgQdLZy5NTY/Pu1FK6ZGBOU
vEg55vXXDG4E2NkFKBv+QxqDkfVQEI/HwNc0TMyqP+NYkAHUANP5m6Excel8IelA
+h5M+5KfQDpzL2ynl3rxCm9365tqXgl8SjF9j5rAMAAlZvgw9unlT0XFmOS33CdB
zA1FlRoqc4AK9sJE3m5DnutALurD1lJjjXwIjMKKGlS1StCe1T9+OOaKopdothHF
kh68LCgCUFUX+cM0hrMiMOzQdhqVX13+1bQrXr5gg5DtsHO7G5ekUDu/RBPlYtMX
uFUe6Eqwtifb0tTAoYDQZc1DMyCgsY088KeBELoqw5feGftFtS1bGlXfkMTXeq+7
uzckmMKhGWyVwB9s/PbhNpG1gWkfGZdnrTrLd7vjnSGDLGT4/vWAAUmUAnUVAZzW
+SbYkfynr03xLL+nLlWAKLDrjl3grzDWMFPAlGJkgEzn1cvduWasutQYRsBXE5Eb
jNCb/cB1zP69yGln0Wy2w7abzSVhs7KfIAk9G+x0TUX2lNXb0W9vvoGD5p2fVPbM
0pFF8A2VYutt57qYqi0qCAEW0gBAJaHBa6dtojs0VgPF+8l3fqncs15gLk3EjN5g
HGt/XfI8oFmIujYHyBxDnFORnRf55AccsjPehogM8qJFKjzC+3BoaeCK++vGnWQb
+AMy9RkHBgrs0jZhnqmb0FHigvIbN9KyKQ5mP8ikiEJV3nRSU+ikisVri2eCGWQF
s1EiCFKK4vKUoJu+ogCWugNBEikuN4OJtnLweZKiY0JlnadSNsfHMXqeZ0NTvTxT
LkAfaMGUrDvmwq3k8RJOLq8SHR/FgGggU4cmoutDsngZZ4C0bk/S4LAS/DGpl2s0
bvrfx0BTnqe57YpcgOMoitYf9ZUq7eOxLNkV541Xjkbc0+30VvIcCpvkhhy4PWY8
lgiTABDhUnJwdfZcHqrdBlfT+963X6XrsUxmUs7sXeNbgs4wqhp60+9/wDEACO0x
hwfFVSiWXsbstmthSGCP9pAZjs4OJ0HVH3y7Gudc9Yrybrs2L9Lz1EPypoz/c58j
R3UHTmS49b17YX08r8fEVdZ9+xxqIZNzGXKLGrc7Qdu8dOYcwmJEbOBmvxFKy9Bh
T7XymgAwqU78RLOuzJT0F1DhfgIjVI6K3z/TNDqjE8Dd75dxE96t9StyxXLnBb7s
Cuz5uNXoH8NsthZHs9KiYYd+Nja3d6IhrOFigOcFHz4qqVAa4oQCwsrYTYYvFqB/
dcvbM2aJkl/CH1b7e7b+zEHhMBl66VXT2+dPIvIlmzowGKzqxAtadR8MYwTaiDF9
Qj+JPsxP3yR+Losez6bnZQ+xOm3WTgZtxaW320nq+aqz5icU/XQjNKjfNOdDo4gY
zn4W0D6EmLTe+RDmFB7Wl7I8E1DapQvHKGgUXlZM1hNwPPVTFVvNWpJ7WO/Ao+tO
NvcWhTCRDJikTTMGCrYH5kE21yXk3e/E6d5pEzAJ58w+ProdNOJU6EWKbCkI+0lu
4jTj5EpqForMsVIZLGE9PjyEvTxXhXbAyYwfKV0ksXikcpijjHl06rUgMGEAaKkS
QTOQeTZgaXQ9qBDD1nuVhqemwbVBM6546twcPLhylnS52gw1SYpr9sj0rpMK3rKK
Ehcl9QAvH8Cb8VVeJA7uqbaLc6g4CKjQvmNMaH7hRrX3/YkiNSfSgxAb0YpAgQs/
FUtjrfeZwupGngjCpfLnIuGrmhdtUbUW2LJrYc18/c22AeG7J70LKaAx+jljwppI
9ppU+WULWc6EuKO5EYjKHL/FjGLa0XwFgfkFM3BVUJ+mbF63EyLLXsi4jE524rDs
neRIPW0ETJR4qs1sea+3xuwQYxTRGy3+EVQBtopLh053VzPkZ7UM5D0XYf6GDvyu
tmBHbOzWyShO7R7off2XERwhvZ5meukw/UB6lbdGk1A/73Ba5pPLW940RLq3wNPq
a+AbFKb6zvk52Q+snCHSwoM30pg5jt5gLncRTLw8XVd9fNPUprk86rAziLaz9yLp
pOe+DJ5GZ7OvVLCDI2YDoP5kzX86xsjOst3a1GGvEeRdNMLBK0tcyqU7jbGb1U4m
J86i4dYDtfOeXbJkLWzypvoky7Gs0UD6l3nn7DOV92XNxXqZkWNwUlhLhqryuUD1
9Jv9ffWC9RbxCQAHNq41Yk7UGUbUb+2xtwngP/5+HK+YY25qtzEDrFPygZOXWW/L
tr40W7Q9J35S0vD9mg958PKSkodjvdTRfW4WBrrFxE2iylPSjM6Cnb8zuWaRMAHq
2m/BBhlQgMmqCipmqkQT4yfc5nAw23mz/GcNHfOZzxSqbxJGMZX+6xPQ/c//2s1v
uWhkRYVWxco88PhnudLZzn+uZowV7evWe3wkCfu1Pb7Vgdj/V1rXkv7J+UjvUhHZ
gIysF1Gk3QYOm5fWpCwqc8xkfbwp7wW5X3Pe4kYNuU93OW/TNlDX6PiRa9yLEOwm
cIBUEV8WAVlzHEWoC7Y+NtToEQFig6qXM3Du/atkhbh5HOhz05A2fgH/2u7eTUAI
2KeOdh92eRNvmnOvcV8isxH9FgKt726xaDDIScgq5WOd/7z4EVwCAOkA7sawQUm6
pNO7H+BZ8H494Y9AOTO1pADGmPW5o/G3qclhf+74lZoccZ/uC4xdxmiJPRf3G0k+
uBNNzzcoG1zCw5OyOv8g+5Cg5zzdR3YGuXefxEim9FABg7rQj8r4vnE2oqHEpjX3
xpNhVnTdlh/2yNn+PRALBuExvxXJMsYo/BogtkMEs/+ONk/40+ffIDmBBKHy0UNQ
GWeoOeSBjlbzqIqkneLlOL1eK+coET23mjMsTM0MystFP9d8VDJdNt8Xt7nA3lWK
s1T7RZpI+adlJy70sryx3idj9g3NSeT3VZ/uIJdt3BUEIGIT/qVZab4amtIbRqDE
jUfomehiWfleHC5/j+bvOQ1yjcrKoNQf6sAFNAruRcQl50HXLMs8mfK2oNUYQQrs
gyMZ5EHRegmy3usWibA0UmgeZDXQE4SYER+wQcl1g0ibpUAed+2Vy69MqW6T0ggQ
0puEfhW9/TAGotKGUSRK/24PRGKbuHmPmjJ2UijNlEoScQ7Lwb78UCRAo9NdrOGS
HIZ4B89t9Oby6kvPGGmsU71tMJfASPsWlPQ5VG66opfKfi5jE1FoPbnrxv4eFa/X
t6sOHTgPxh7VzJRJd3feKqZKcrtjiTHE4xy1y3v0+dDa9hK6KrvMjxDjpKrZAoEg
oiazzV1nzZzuFs4tmXVnI5rGdivE/ma32xvhg0BUg8LY/FHPsoHTuSTQJbUMhxSP
pz19xoqyGUHyIwyJCOrZ9GwJoWwA902DAKIPbAIyNWWYpKwAobL2B88Y3PziYVn+
VovO9vnCneoTW0z1KgrWd0Lr5FDtI5dbGgvy6OnQjt51aHo50lQwaOoy8OderEDf
sfR6CqpU7ykyuPYB1ig9XcR7AwNx7alVWZ0F7blDScoeln4330aithtzlyFYM4RB
y1wECU1tLYKVwTD6DiC9qxrTF6S4/27UP3CBG9Iw9chDJ95+vHkQzjGA2s67I7VV
trs4TwnKTM6EDfUPHUc8wq/X8KKzYDNCXmRHPen/LGyQi6SitwFxLwNeCCCqfpuu
LGBlQcg9K7zdjzmm2oqcU6VcxtNpavWjXaz70ZkvIOUwR4aZy/u7r15B/MTj1b8S
5z+ZOI2l7w2rbDb1763g5ZXLLK/VzAtqVQ5xixTCElYH3LzHzUaUIjoAXjlQmCwA
Vv4wwSq5IOm8pPERzCpW2MAtzCap+9vRT5ohwOKS/Nw8ZTlxLrPWgYtVCaPxPmrM
j8lNWA7JySz9TxcqnX6h2n7k2ZvE19u67hWjgSa1yqQ02Dam+ipEqGIcJMGbJPGe
ruRqbmXrLtrhB7lfM6h2DEhjREgHGNXQBNtXaEURMj/0XM59bLNIK1UyeaR7OBx7
AZc8Gqi70NkmEyD/ebVbY8q0n6BP45hn+Q6S+tT4bthMlXwB6sPuKlGBQCNOJ7xp
hcT7DSyUAxEs/62CFs7JwwVoDXEMyZfd/XLxZbpANBxy4IbP9+6TB8M0uKM3ATlv
01gVQ9A1PMSWfXI5IS00lGYMbXHU6OIaBoomUOs1xRxZKb3rjIy2VgQP6NoAhINh
jRzJzO6OyouGjPpgzIUfXt9cfK/IHB5vTgnvvodT01KtWLXWt9VBv/3h9Ip5E6Dy
zHQ2zUWohZgSXSMzPUjm9JVKhOwI0OfPL+e+yv2CrRJnrnO2gq+ZTnvcvvM0XCe+
V5aCYTGLvp+7rV6h/ZXLgAF4JeKuT6bY2/nTbiqtKKA5C2n+Mjo+EJcAH7+iwyg5
WSEBs53Rx2di3o+7J4kSFJPgq6rA/zw6jAuMpDFEmcdgBqjQHvilweVssLb24wvR
ZCyWi3eo17UD5+fjHSra8kB6+eU6Jg0CHjEad65pUZhdbogxo6ZZ3NnZ/fI+PqX8
7LzyOXm0jXi8f3QQNAiMyOGPjCN227TW1dIWS35/CiNQ0gyK5oz8F1UTxT9vORBm
hU3B5JFnav0Vc7HUv2hX5IMzf4UeMI9QEv3SWHLIQ1XjU4Fnfv/tG6p6YRsa11YF
oALw70UTnXvzxafM2GHRpBKyyXvHzgSdIMFVH7gMQGZ0+udLuiUXwqQUkSHUf5ce
PkYCuBpH5gWS8vc8rpxl7fbfsf59jlq4gndaVTBViWjozs99zubT/LFb5uXkdLXz
ooGi+2RkZLZk/y5PBNVCSXgOzs29KLsBS9L8S473YTlDqfvJ3G4fXpdd226tReqM
sY04ingmsEhHbFMiK4cQtQ1bWkwDV1mE8TXYU7TRZGPXVz42NXe8/4fmBU5SiBfh
YbaEgaTdlsxOaXFjpX1EXDDhTb7+equu5qBdrZ+lDpoxxlKdfJvJDnH+wahU+4l/
U8tUrLXQQevB4KKHV6bK7ThbbzRFEWc0mfJ3F/mf3ctIUSmjQqJbg4Wc1Ec9a80c
xKbZLhsnzz/BiDXp7TVccf6XXjpYnArs2PigjFb1G0UpRNrqaEZhRabguDjFqcfd
1q/FpX3dptcICOKhgE/vNKKVb8eh6Wyi2fgkyqW2cn0eLmFXB9BwnVf37/GhGoki
2Y9doEqW2Uco23ZKvyR0LFnLb2vTFQJadJmV+SSNTZjZM0PpILYBdglupz/aP970
ZAP9OYY+HrFCxc9HrZkF9smUQrU5BSSwVCYO3w4rk07jcOpQGnisOdv2bM//1D1f
RwrHlEJOGcs6iIeodAxPUfdtJ7gbS5mjHK4lUInWU/oLMvNa9jJMMWk9JK5Ve2kG
jdIf+PTeYh2VqaWWedP6IRFb1wlJM9d7/WuHzl8MBanFlOLtYdwP5iDcDP1PTe9b
FE74ejjyWd0VRVWhjHQkVwIipahSQ8j/pAdxJlgY+vBbZ8k4QZwGTQ364v8A2wSP
RDXxiAZM+8kWaifA5mqc9MSVz94x6n6mOGUncFRug0YCd/rLwiTeYfA9mBaPI0LD
b5rLPpEicVc07D18VUmrg1urOtoB4ZXaKpx3uVw2zFLYTkzO06e4dp0VJ1gEm2AN
BnAu6GnCuznZNQ6xySndQ8742tRP7htZM9MIQKTmQt4itZv9wUMZaZQTU3Jjx2xy
8FsCPd7lca3ljwEWTA22kAR2113GUKUQDoGe1mUcx3qGXBIW+/nUBafPyWH31vR2
qfDfS15AGeHmR6y8/nAAKqEs2Ae8ye8OdlzIdk/D4pWVuGFlUeMutCA7JYzvO5uG
pXtxeyp59bFWxuuA8FmJrZhtq1f/+upZ+Z3WzckliIkcsdhAOsnSXXxLgaHlTeX4
0OXjbNRgGpDF16jHMyUYfmJDevlZJEJdc9SyF05zFsJpFmcTDB9B1CAcxOU+zvIw
Z/cND/S3gwAUJdQOA0cIJl9jY81M8dndgVhjfvjun7Ln2Ca/XI4Juykqh69r6uif
HijCDfLuq6xyiLUScXBnbo78RYrGzo3cl3+5Y7/E6Qhgqj8Dxxa34ZeP+llAp79r
CtccNb4pnqXTSaJukEI3A2ZI6S7erPXJycYWjzIe81k6qbkLeZnNO8GQl1nMQj1Y
Gdh5wP9xs5yLsz88Yp65b83X3RIHQtEti+GuJ03n3DBwGCvlFikE375c0v/Wr5i5
qgj+QdJGVGmxZZiLtiR9hhqDqrwEZQCTRHaxEy4HjsfAxIGx/Av3WeWW5Uwk5gd0
J1KnZLL/iAhDEhiyIHdtON1Tcddf2ZNkYWFkoUmpVrBndETFDZHzqqhSpMudpHyO
cmrRfSuDNd93HTwLDxnTBmfGGytko1nT/aZifUawyiDICTBo+chaVivAE90MyieC
ZXnMDa/kgHpdMbPz6nhCYs/3OVK7ZVoVxMMCW1Q3c407lxsVsAPYKXITY9yiH7Iw
QeKdae6Plg5IwyrjZKCKzGdE7L+qW94iUKErpeQSRJOLUzTPRqjpgzoGH7DJZlqv
41B/xreh6sGPrh/xJIR8qzbVnfpkJqOU5Hpm6qd3Ev/pibtoFYQBjQPpLcIHd+/2
Ylql7g4SAm86fEzd7zTf8CR7b1+1KpEwDixEkQZoCkBxZouowJt2PGvDWqU7u6sL
LVyXRH0GuSPKtDdyHQwwsaOH35bTF/JxgLhGgURHSDdCzPt2s+Iuo+QlVrMk23t4
5+tGohdqroqz0BUFkOuZKckzG/AVKzOgbwC5MNBkEIJqyfcGbs1XlA9ePmTb0FQJ
O2Vq4IONyGmkRvQ7fpLwdqysEEJclAhrRqHkSc3jnieTmkZhZgmwOjF6TaCnmcJ1
k2pc+LgVMG2Ttpel9dYvolYbnDM6/No2Orj4+LoK2uaXtAOzwfAd+W1O4gk2HVwr
1Z/a8woEF+8Q8eA0SvxLxSjn9HgIYTPVBmIwfgtTviUycdM9kfnwPOm68Q8Uh9cC
AJKLF172TBxJfZF2TPIcpdWpBWfD4yFiU4fbfJ8Og2zmPHvxwkKUAxTbIBT3bF34
K4aIEeEsKBYOpOFastHBcZ8AJxoqcv6hTUfsS7lKNIxGM7gx5RFwQ/BwKSyi0OoO
V4chGAZkBO2oJJ1egviYfexg9xlr3jMYLlyNwedGTrGTwCmLquQYUZJK5tCFImbo
SWeQEI3WAnfCGN8V8fCXtxWBtSF7PvAKWOj0mU9tQqKPasnvREqTuoGW372W81eT
ztUOtdz5Xn8W2FOCxyxHcepih5/PrnFU1X65AbgEV0RoM6+AGnXX6vmw9+FAF5Px
2WSCUFoGmfOR9lwlivgGQjSfjH45hZgByKhNQQMenBkcRI9ZIpFPElYW4YkNY07j
/zEClEpVj60MbaykFrePlnPkFMB210MtC6DhwEf5vg4mh3Af4NY74it+b6rDngEz
`protect END_PROTECTED
