`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gdd7czahooKCk0MjuKTxGd6UY+KLuFB4dBjgyCE/FR3W6K0UbixdymsVOtt7U/A2
sr+ctKAmuSYBkngyqKHgZuOP+H/pXbgWJoqGdnuuw3JyQytNwSvCpZgb9puyH9BR
UFZAcEk1cAdVLcR3Tq45yvS9fIkuS8l2YZRXlKKrakJi+wffe8iix/2BcJcI3VIA
hTfOkzf2D+A/FkRqIhDjU48OdWV2ScSiVNwtL5EUX/tGCxRD0PLQIc2KSXAaeNiT
s4Fx3WScXcdtrZ5sHmfGCUZjuVkltPmppOpNZDAMnlvTXMDXTfjWLxn4GRedOTsu
xoGrHI9RijkMb+4JYMfysPa6BNo23BajUf6/K5ITLLiDD8xSBNezyanRxGU6/wOb
srvGCfBQBgFbkxCpevKhJ5NaXQ5Z5FOrvvxNtYEEvr5Ls3b5PEguY28EkwVaVXSe
UtEOOQA/CizzX6d3aGKOhOPuXp6cbQ8anS1yNR6h54E7RNAZGBRUEO2Zqi7/1Ffw
dDWH23vQfq2X8JCqbO8A2DoOFfvPDhjZa0rsx129umiQ3yHjMv0dDISbB49V9fDn
vncvW2HamTGD4SeW1DLlayqZNsS8fjJPVEzEY6+DeeENVeAfcvhF+4Ek1HFlfHYK
Q4d0FJ4rJc4UZ7jhvwCJLxSvp+WhvIEsFunCDvn93lwtFvsyblYWDGSWVUTZXZDl
7vMUVjkrtOLzpzMVPe9aZc6N7ONW0QNt/N+WCQAlpJC3A7VmsdiGkk1EeGxAlytP
IeRsTWTQxAvWk8ifrSC7Rg4ZmtSIpCmpJfCV3k7L8oOR6VA2taljIw48xApznAMm
2kHi2qLaJcl3x5eiP6dfa3IipZ9iuUpwF5xULwY+R1NTUJKtyuAA1MVQkINlI0Ax
QWpwIhvFlWLDdTgBB+TYqD6buE1NgQuMwcSYsrNVORb7JKHqLnOZl++qnf36HiDE
p//gPA23r8DcFdp+McPel5IVm/3/IHUkhpCmo6JaWrbgo4flzYQw+w1bgaftklQ1
/Zw0+1eO7KMDl3VLccvpYRYsv67A8IZIZiophKkIY/K2aZ8M5mgvtlzePepJY39I
m0b/z56tSF6uhkOrVY8+/6C1CdppyKpCB6tSrFNCQLR0Rmd9UPTzpt6RX3Xa39fV
CzOO6hoJi5mnfAU4jYC/lpaYQ0m3bG4RBAnbZsrURZ21aqmptJgdM3qY//TMys/y
eBR3KC3o6tuEApdcEn1yUhVcRxyGMo+Q/7dwKfASIO+u4sNMq2m1PeMStyuG6uPa
Qn3xI48nJXXq+RANFJPEWXvgfDnSTAwAhOTd5BD6saGJM0lP1VlpF4OMLVIXGBIZ
5gTs7He53mVZSYntIrFgVdAK6drMdDv3hzbS36qkxzH9mtLOCV8/VERJ7JoUU3nt
1RVggH8Gaw927FA+iGmxLCtb8fRBVD0dvQSzOFngLhlx/IC+LarhUB3rDiIBkAof
eggaSTfbSy2VRNHodPeFTflBshpLoZsxGwGLyXSC+dU924PRMyBEt6GZbGELWUY4
jyOOQmHMpK1V8QyY++v6df2rzWqassih7P3z70cwXlz2/9nhDQ9QoXHDmTqtFijc
XuPiu5eh/IzpPdUJ3NrIo5uO0lQENLncorcB6QkmsGNimxPaYeX7VaSs4Onw8PKy
GGftXyyR2q+An2NOiEBiR9Yh32aFZoi+D8FGAsHw3GuNV52a7AuZOEKAbrGjGi0v
J3OA6CE0BDORUE4Dc0Zmwgy+RDApGM0PFbKHzaNyTxDPCGObeplAaUqNYa7WeJ6M
RwGw4EsFvdfe+XQkNEkfV1qS10RAEafoqoZW8YVPW6QM3gMzFLX91ac+yd5+nGTN
JDDhmGVh2dV46K3RqkgP3JJwTje8BmYxAOP1VK++L3UsUeMpJ9KZm1zhjVodrGA/
nM+gYNss0Jxa4NaEsYGgRb5UCHNzsVZh5tmrQyjRWLvnXDN6iJXJb0droOlRA6cP
Hw5OZUPp2h69Cw2iZvBd9clIz0aLaIgtQggF8zgV71Gj7r8mW+StyhzMDvcOzqg/
SjMwzCy/+mQ4PO5mVtmv0MbY6Sj8ARKLvDIZjJpD3ynsOMqb8/asBjUZ6yt8551d
6M78t8ESrtwVtZ0O8Tu/643hZu8pHWwwKcCuQacDRpvJX+1uzqY/mrABFim8c1cU
QNolIs/sE329uVtGHuQf/waUvm+nDRogYcD0dsEx0ZZHoLqOVdY624Q3VMFGREqA
jCQngTVLstYfcc+p0Zvj1ic1CaBvBbeF8lZtFd5pvMt7Kc1JaYtnDpxS9KJvovU+
8iGQzFsI5Os847eGluhVtg4rNB+LZyIzZ1MEpjHe0o+3qu94Fbf3OBUaDzHIRVyX
5pgFldJXT5A+aBOa8yamtmF1RMggWNbuSyLApChVl6bzB+KRUTYTh9rITa5d7MV1
xzb+wx6lME2uIMHYUIKrMY5UDUDQFuV3RWf+rAHhEjwDxtnZ0XEnjSOB1HeKLF7g
fMv3m4FkoWrnMeWf/sWYjhW5pNV2l0mW7GL78AZSKUn9EU03yK063Jia39PeyJyB
FUNepACK4nDbJr192ShJ+N0KreUKXAdda7L/ALLp92cJgO/EWyKrsEkkHuimEjg6
ZutzPPn0jMMUftQ8GvBJtQ==
`protect END_PROTECTED
