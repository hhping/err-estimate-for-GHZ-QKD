`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmGhMH50mvMUKZI6rlbAqf3Wf0HIaRFqeuVxLur1s2lay6DvTp4Gl70K5ohtCQrk
DguDUZ9Hg2pzym0q2qUoVf4yf0sUqZIF5ZzmBNYww6AZdooA70lRovyXzxvmNoja
clCG1b0qHrFbViHL2XVLX9yQ70srulc9cGZor9rmlMkFyl34spSVgJ4tuV8YiZBx
uSV1Ej2DRw+XFkq3EAqquSWtdhMRW8Wdxfla0JswrP/cy7QgxwYNbG7/RS0wWZjK
Ly4sx15+rX25qnUVXb+SdgK+LZfaHFROPba/batRAgc3vQWTfle3GUQzzf8PJqKa
pwCuiJZmAkdmgXpe59LFA5etqm0Z/nAG0VRUvrE6Pc2O4Ucg1ILCG2A3E+b3mDIO
VJm7fEVlR8Mwe2OrkJA6WRLplvmGH9/eMVoOqh8/g4mDXkrhncMgyB+FYYvy8DEs
X+boRyDN18ROKTaaeK3FuG2jEQROxludRf7056cuSnwroRLi8JQnxCMZDBDsiSUA
SpfVMSSN2HRElEoAz7gugKXbgxI0uIjpWBpH7c0eJMIfFVlSfqAr5TpDZ4jIX6Q7
qfSjHjdzhGB3JDw8FQX43SHrPQje+ClnTOkLabEtflJWNIgrfTlPEUzp30xj1eaS
BF26BfgUVb7/Db69Fjb6Okar5LOAm6RX14qKBuzYzgJtQjXoZGyLKW3V+x0aNvlA
LxSBfVyhq5hvDf/+9sMi9xzXEjbZZ4NhkSTkv+hsK1JRYZIr+zJQEDfFkDjotZu/
VSYAr2FtIFWeqmWDPk1ym2cBPDWxrIC5nddSfC39T8Lgy7L7ryPK4ony5i0tJ7Pn
NNnhMbOmZ3IDdBM+xEmkJWtt2UpjgqaF5Koam1yvfFrv2d3IVtJx5ivFWAyMNOlT
qwyC7/o/KJQKDHPFR0iDC5mtl+NnCqt9JL33l+zdx27MIXlG8vSo8vt+tUmlfSKy
7TZQlKqE7oIp6wUjt1vxZslrVSiko6SfjHpVxfJVxbDk5sjWkQoJmrNDTqFBN2N2
ZetNOf+JBU3I9OuGI+3YfpQBEhiy4Fv3jtJwQrH3MuzTgHGVnX37s15RPMGUeJSe
HRZcNhmbfKysMgxvIeUfSIc3Htc4aIQQztBIEkkSFC5lMUj/C/zSDhyIm8J5Uw3K
TdgiCDnmf+xXeyfBbHToRWuxPXRwer/w4Hhe6mSsa/Hs/Ja/gKd1hcoaNIONyxS0
knS2tiTzvM2dSKDhCNzNFluvjG7RAoc5/qAnkHScBVYf/gXm5fpfftS6G/KD46rL
/nqE+apzY2fAQg0XfyqoddlN9On7VIWHju6CWONcnfWhHaUfxtrGJV6YKdo5o4GD
oMygp+LC/Q2QctpCItgsmKETdVVnu35xYC9lxp/L8AVdOTFDHW+XGnao6/avrc21
740H+l+Drm5Le2Syi3APUOXGgo5hsq/rbQjvRqDlugvyjQhOPzE8NO3U7o3Yr9VQ
KnbVjIJCewlSg6PoyR4cFb1m5ZeQ6DdQ/naHv/uult6HHQV0iH0K5fA5UadC97mT
mtGjA6OEXlv79MnG6+3bnNwANcwT0HZIlI9wycqPn8U3UWPiCOz4z+IXFswYpngp
0TXcKJMwS6Wusal+4sP8RHBejPpLaPC5MQD59Z7aD1r5SenFn//pe0jIJkJZcxat
pB5A6d7p4AmvYNvRhyGrkHuMMAYtOreJpU8KADE8YuWrwqrQBVSE9t/HgjgGBuDd
7UD0JeEt7y+K3Bu099ehRv3GJ5qhS5Uo1Axlk/WXszMB6jf9L6VUe1zd2vQ0wd5L
7xn3BAwA5IehanQqZ0SWyiawVyRVM4CoXzLg3kNcU9h0jrK1RhDWxxXqhvrAmFZx
9KtFPMs1KI0Xj70HqF5WMbYr58w8U+2PaGfVrkaADkG93TpuzMomdpCArQ7xC27e
QGUMe5aVMmU0ZVy+OXebfBg6cdxX9Y+ybRTpnbJg58TCDyI3qVfrmCO7aYcgMC+R
37Lx4V8MVHahUbZe0EM1WJ23Kt4xy+i0UGrQQpoVXGPX23EWRcQ2p2C+3XNGdXVk
/pTFnzMNOzBhdWDlqL0DReYAHBNhUEFTOJCdnvXqkRPoswG21xzogXd3k7pAx3yI
fCCmCe5W90DWF9tkCz0aA+OSKT1kiG61g1/mTWAej662wKBfSayq2zOnYrOGYsiq
V6uZmBaqE2kvmwJtNPF1ZUGYt7Xdq2cX1MgTcFVZ2BTpA27FlOjF/dsNyIN2yUDn
1Be6J5312vMBiXRT2CD7AKNmuPBHhmR8rTWs1F+skIZFck1Tl3od8ilLBaRnqIuE
W64woJzSlBn3UBG9vVsEro/DTVKHARzoKEG6D58VwkOHVwwDSBmz1id3aPOdt+bF
gQxa5n5TNns5rEm6dAoeqMGR0M1QV+s4P1bvoYhrcXdcYzBIHbTQy33U50AKSyhQ
InUgUax3Cy0grltcZ+RWb+RIUvu5rlaUyCrvuCKoi7ZwQnY/8U1wA3zYzm81+C6w
QQXThT0Yf+/jgCu+1rEYm2Tgtc9zkmE2LK43v9sE0kpkAxpM+GKN4quxchX9hjX0
yJd4BeVYGc+T/J2Fdq65vuZLTiIGu0I9Z7XoLDtr8xIWS5QkvOn8HZ+Ph7UhAsR5
emOXXAB5NPTRCou8+rRrRhGcPZKa9R4Ng0p1OMCKd0qY4GNIslVvZ4zi+edEOpa1
UBok4a9oi4jPdPi4ybgT5vMdTh0Z4uNBwfwcFQh7drq/i7R4YqIjR6KRmpTAT6tF
yJ9aYi0Y0XFTi0BifvsvRaCInQ5rhVdRhmAKO4SARXeQdv61gLxHhT0grL7Gnh7r
twE/lNUMBnUxuUYBcntI+9oS+Hqkyr47LJbPB92wPU+Uj7m/Pv0W5lVaHGI2FsYD
w46aldvA6vvZoAK1daP/Yw1KbF4rHMHCEA6Sx9c9uglbksB3alHbb9hQX6TeAKlY
DLeynIOwJ+RGQLdeyHI1Uc+sby38xr8faHzTYkSphzM80yjuUdb+9c+zKVYiGGZC
t6D+d3iKKbiKNVNZ4uzbSYvsfOR3Js18bDy8+X3Tffhc9YEkjIydlxnVNQPZVf3i
FZWfG9EBoOmkT8vpXU0NJo2B0vOOoJiVAxyIXgJY6jOtyTYgqEq+qP9v/E7RGcLf
4eGgEofA2O0fJaPKh1CIQhxo46fVpDvhLKNouVgU/wFbKwSOrAhrjpJNEKUum7ZJ
UQYZd65CqLU0swHyXvjJwa5zyalSD3EZQcxgcpINoc4I9vLgn7qf8uzqyOULvQyk
4GvgrmBPu8fGYIaSiaql5O+Tcd0JbIyTPYgF98AqzdhzLKBcQLtxyPtvLpU8cZpN
1PHiLN7Zm/jN+tyqBlrgTFh3njp3Abn8dF2M0KQypYbk0CA+/J/DGydG4Rha2CXQ
j7xhccCZEGipfxgsoGknpg+zR7a1w6E+2R5DMRiqBVt5oINxUAPoZIEBXmaUnKUc
QWC01dkuG+1K/ppNjIKQRR6+bBOTWTRhFSvJkT7xv7M4wXudWO6H5tys4LjPXVRZ
uGdT3EOy3hZrn4HKk3Tx5+me29z7KCRzi7uZLtp+lMSBSghyuzlJ1ua5Lrwi/Dyu
HhDgPtV0rN1YYcFQdEeZQ7aabJeahfZDzORxWBNRDzhBKeR7Y38irCUT5rFFL0Kr
zdVux6uttwE0CdNSFEFpnz3uN48ubTAZ7R/h1S7cTWSPOUWxWd51yddylGZbj78w
YYeCfem8paIWlytLTX1HBe9gx3vJiHQkpbKEKpMNK36G90ZmDqKVHlPMKqFGJp32
/iUXfHD+kChp1ig1afMJDY9gwJd2C1F0Y8KaZNbsrCM0duKSpp/yADme8jPSgAB1
+wSaELbEN6JH1SOQWwr6Qjyk+eisP/fxwnIgNu0P1/3CVplX7YEnKB43AJubuMQi
Z15f16ginc6Mq3ToWugQJFLsNRvXXm7WPlhE6gy0DIGz4biLE/S+kk5eV0WMzsP1
3D1PRM0W1/+b3guhkOBqb/4LOgodSFR2y7qdnVWBRAFSznRXRgbwXul270q5lVdy
Fm5BUenPih/SP1AJyv1bYzUmLreX/vwtuuKyI+XptUtl01cGOz5AdV/dHb18emzv
EeO456NzcLWvI1rs0uquZKbWb4YC/KbU5IIKtY35ctFIhVPuHIwD3bE0hO+87KTj
wIUI3v2kuMnsRTe7VOTaeburiVzj209tfg7B/BWnO3SkhPt8TslD7PN6AZO/V6N3
GolnTTRm+R8q646LXlrBwwRf9KNG3uXWP70i+1KqxraG7YtID+DVaCggLm4hk17Y
ycYvnEU9d0uuB5Dt7z8POs4W7aphWNqBs+Tm73rc9NZUTw69SbHmbEwOqsajl5ZQ
BwYdaG4CGM8EhSNdKoyskfLDpH0UYwdTU8s6lFLKKqXNJt49ipXtCQrqq1RADn8K
BQSi9Q0idLBTsvbQHqviH/QOhVMjn4CktqgaHpUA11a8jpSgKssmZaW7EBMk3dGW
M9mcpJD9Pyn7OZsi9uAQmuz+IDGITaPRprp+BUqBiTd27Wn3Hnd+W5lKsKcR7K9/
GT/IueGET4nDvdwLwZo+2J9GkZ/LeZ8mYEdI8Mw5gPHf0trYRexX3Ux9RauKfmNP
Xwnz1LkPlAtNvNXKoqMKn20zeMpV2p7JIItb8pXVUCiJHcNZBIistVSlHF33NG5U
`protect END_PROTECTED
