`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7DSV9eW3PlxD4PJNKUSu1taDFKv76jxnK9AS5NzjcCiXyse89WmXt0E2pq1eV31
afgjQ6jpJGgiD+F/9igf3Kh3zz6RCXWVezvoTAcKvB5CoG2aVIAgtddecphE6v+p
fb7ESFT9aPqSsdNVWVsU/qbETGEFPo4yIdupmJ+tkEgqq07ooMAUjvT9BubXtIcp
yIdz23LPIc3pt3/8kRCkCoClnPIngexn+mDyDha7jTIjZXmW+SqXSuVzbtea/kdU
1Dxd8sIlN/09LquTS7UhvofbMQGflreF3A1fg32ZDO/fAdW0eS45sr5wQKD65MDv
Q8j875QDciJ7Bg+pOwL7hySUN/ikgF4ehZ9UGPu2ZxKCIrY//VIELhClRj8nDIAr
ve7cV9HP7LZau2IW1U+qTZ6oWnDWlHXEWtR8/yhVHG1yhMLKFeMOSDHJ6GjPfOBH
rvw5YPsk7KMGTzgcT6Sc5HsOMz0Lkr9uwjRnu3nuLRKdn2T07Xgx+7/VKr7Q1pTw
BfLY3RFsa8CvnldSKRkQWXwaqS98P9e+YHCLWPa5AqzpZGHMQ4HlOV2Jw7Sqa3ul
f2rGQ7I/WSaGGEOYbsx5nn1AIrfBye5gQELP8iKyUWmio0QKXDwvFg6okOng3YOd
3aQxiwxUz474E2BwaQnm+2l6ERClIqIuCfBe60XFNe3z896FYA+E7emmHiX7jqA3
TyqCEoOmKOV41dt/qoC0cWjYGPIucijOHLe2uH6+t7QW0gAVFPHNAu3SFKyDvmvi
zY0hcWCv8zxpARVelAs0GJ378FVqzROiCag41eO0tRCiJ+6amGsrMG4AkD8Wec+/
/d38EMJA65cqXAL+yWb51zx79PxYDmWr7izuzl4wLdhZVhiC/s0Icxu2DXO6l9nq
aX/DSmKvUiwU7ne5fAw0929xLgBga9TlZErkxVio3zMCOstoZUI/yW0D1SkJvrmi
VezFdBpDXRWWYLPQpPIRTSoasMpAvXWxN1saSJ7QluMrdixJf6UKLAtHcwel95D1
FlSjR53I+ycyXAcTM4PrBsZJzxJvOKn8M/3CytGxcgKcMiW8fLKxRv/YI28r57m9
BMEjomfmmprpQlQd6dOfpisKF3zS9RoijnpQIvP94SPvlABFMuCiWJVjzj9EdO1c
gGOmKA1O/cKpUBXuKM9BbNiZiXxox5aTkcjYXxSPLcoUky6A+5vvCU9p/D86JOfP
aCUddTNjES/HcKZTK5DpdhNFZGS8HIap8bo6DQLKIWtlSDmp1tIvYtenNbvvEsgy
8gUunnwRrLRmNAmhLRz08U/3L/pekyXKMzqZpVcNOvHQd2mKSXOXqgF+T3BtrgeG
LRQ5Og2jUTVeqwhViiU6MfhFBBU2cnKDKPkvHwLMNODYgmAZlteS9qBoW+41wJJk
/fB4mFTA1CFWKMM7mehDTrdzUQCdck4E0wfwAHPk8VHUD6lpT79RMnA0FpSZBMvC
lBDcN9TWqSdanUHIGwrB3HUe9SHbL2A9MTWOERClxjmWy/c8EphQgBcb+0DhUD3u
XXBheTS7/fyEsNe8AMk7LFNfODr+K0egzBM2WpTNcocmgCGgcX8EBnvXbicQBCY0
9kjVvOxtksS1J/pudd+U1Vs4aCyi1N0F5WKbo0xxe2W9u1tCzZMgmFKb1rsJOwGg
jUNvHGWtkSaRSkmmKHUbr5sqLLJ/vlF5hbhUgBHfI8x/4mknw7q89rDhFMvINCwF
2iYR3+MoX2+iXLFZeVtVGHB9cbtwdkdbFM3lT7wJXbGS9m3hRUOXplhB2oNvReQH
IjIssyxm+KDfn0CVvi5dRf1vmxeGqvPWUt0NM5INCqANAniIxdbLro3vwovoDMI/
mzvqLmtU582ntOLn84X8ZhO3AEQOiNMJ3meGePgCVK/GOH6M+DgfcmVISHlHPWXU
g3gQ1iMRloHoVY3tTo+kPdoB3ne8jK9WurE5fMO/oOcpdBxnFalZs6Q8TD8GLIyc
91SUq2y+udDX7lSzZ0MOO7P/N+BxaZQEjuLCqKgreR54e6FeoFxtx5RMKkTuHqmj
bSyR51o8N3Uz8xA58vaAfVetDtGwHB1NgFYUkP5oQHoOi1fJGldNrWUHrK2V1brw
jYxd7oNfKSRCsJWTu/AD4VqMbF0IGNAtw6cS2OM/nAb7DOeIvUTmWeXELk+MDFQ2
bZGEYqld+Wdw63NiJ5+DiF/UFn5iERVYcFysqcNsNDCeamx8+uwNoXB5yYtZF6pU
GmO09jAPrPucd2ElGVDLCB2wotDmwmmev8HT7MyMx4HUEvUBT/qcZNcPT601cvl5
z+B/a7sGlHIj31Q1utLYO3Ml8hbqI4PvJvxCLmw+t25sFmFrnpZhu00XzkN6T8UL
lfUPbV1LKD7nVdVnkm6q+8S6K97ROSkLKHcD5O+gxxIsy532heagO4MS0a0VkG3j
wdeb+qVxJUPcDrsuf3ZZ+GbwjeqJRZuWhSpVUeoD7Qv3vS9os7rH5R8zwUT+NTpO
NtZbsASTQYbyy9zF9dflSAUZ+z8TW+N3rojOwagR910Qyqv3a0mn4SQw7pvYXEQ/
6nkRvhyvtbFcQTm1U7F2egqUxuugcrhGJlKqfmzNZFvu5JI4ckGPuh9EwgEij3Zp
wWReTlJmjkBU0Z4QX8Rw5ZmDhv1nNYLxnF6R9SVJxvgT2hjGfhFfi5QNsInBFxTb
Tz+VbJ+wgj9Q1gEvIVh9zQ==
`protect END_PROTECTED
