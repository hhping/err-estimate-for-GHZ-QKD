`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hpet8ZhG8zkZHbtzt07H47HlzAxRlUf4ImWGTwZV3YK8hcOhwxvQPc29rUmIWBBd
zrrBwZ09wzAEI1UL5PRaS/MXU8RR+y855UZMEjOU8GybVZyVnVVdaetAnBX92PuB
tZTClj2pTH/T9wr8n2EtneqzyAcnYFYXc7NU00xJNU6dlm3DfVZVFa78SUCbMuOO
NYW9cumCGVPgMUXDvSAHgF+T7ThwTVP5Y+df0heOzEkc2PoECXNqRhopNjagO0FO
pEkPGw/zODbFjqRERQ8aN9CHJUt0zwqE8H0iqd9P6q90KN/9IMEvS2XhBbKhNI/X
op+GYRXmoglVkWO+FAKxybfJ9s7yKDJ4F+1eJCItXj3IhXHVQ+WrfSMS+DtICivh
FF0QsDVLjU6waiuBnP0z7UKz7cs/rJmhtb0b3UtdlhwTYNJFdc+/bLOXuK20jlDa
+ectSWN+nY+mI6SZ4Q4JIw==
`protect END_PROTECTED
