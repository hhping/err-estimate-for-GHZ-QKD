`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aO+8dXg/c+KPyiYZsWcAfwKzJm1p+pDSswM2NmiTQyHjMReRv0OPH87vS0R3r+Al
WSYy1xJ9LDO67Cq/NlwW5sXepJf4BqnpIqDiDXui0ZMjsNqibF6PO3dCTsykKuC2
gfisGkkNXDFuQdXkCXrP52pstyDaAvT53Wcyi6c6KwT+kqG0zrFkcgy1boXounA9
OhLnb9X2WEBcG7E9jxGzqDSUz7YH+TgsbUtWJTvQvfQCuJNG6R+IWabALeA7jQOG
iko7a2LoDWp8PdvFmwZ/rDR2zCNzpXIkgV//RMXYNNwmQzoU/tP9GLAylnLAkK/k
SH6c3XIpGouZ4Jhw0e2uhp0FXZoCA9Y6tOtOlVpTxA6h5mPrbDoOiUWh8NL7YuhD
wrTfRQwE7Sc0u5HQUzWwJuoa5GlWdHyWlEtI6twcc1FS2O+rhwgLXB15xJcMDLJ9
+WzD9OjS634R0MzJlcDLrWk2sirXy6adqpUUjmhuO6DzP7WbLf/B0+bfREclS6ll
gKMQv6RneB/cpsVfKAB7pgFUkPQmqYTTCvzI29a3bhfIq1Y+sHoflsjHlpcQBm4u
yy1DwoN0u1biTSoyl4/pyLVCrr+lzds7MSapiskFl3RJcY1O/+tERsyPjWtF6IEX
bu+NW0rOIHvMNDV7FlhPZPxMAu8Xux4wO9yiZrHZWVxuQJI/ZtcUYP2qp5rBIRSf
EVN80piWr9uCyoGnTgaTuRcQ3mVL6def68OeaSN9piT2O93wg9IO/bRhxNyk1mIQ
K+i/BHeEY8OrRnndsykXjRjyzYqpLHQci2OSuwRNG3kp5pDC/NHdzdJrtAfBtFzR
wUqz57qqwYn2NVG7cNPffZJXSrXcSsd4Q5BZ5u5ggLo0IGS0N+PgT1UVeyXVdY5a
wT8F7jURt/cIn1J5rAnYEGUIWl/OyHaF09ZIV7wX2s3sT6MzNg8wa7rEzaTerpLn
mQEDaJKvhQ9q9+1EJxP3WXsEvmPr1lWgVLxbmGU/7IBgGPx6isOWdHU6w9tuzLT6
jpObdumkqx8jt+qu58NyIHOy/dSIknqnUmeFLvR4+2Mg+vJXlMDt9AUhxxjFKMTe
1Mzy++qqKhMHFl6e7fnMYGAWe3jlE0Jy4Kwx3WfLtbILv64gJ/dYF3Q+Fo5a/G3M
wtALAUPMo3rJ4xvasjVidlHmG0xcsjCVIAie4PFadq0s0nl2riNdM9ISBbmUf6BJ
neqOaF417HNqTAMbHNgT5dZv5hOyoV2DpJn488VSw2nzL/gVvc35qFAQbmXb+sXL
yFsLU+oQ9ObG417EGg6XABHEU4Q0QA26NmQbzpDRuzJ6ON9P1Lzrb6OnUVddVqNa
u0HPBmSKDRQmifoXcNs7OMtlgqI2MyeUU0f9nTmFXHBBUNhweFSZlbjWsootC59D
hB1GTaQWoNby0rS3bq4fLEQhgn0g6Q2QPBLTuD8jXG3SG02BpKK1va6YzCOCl8i6
XVwaI8JjeSDomNcE4vSskKNSPckmW5fSVFI3BlpSiChTWVvlO7HmnR4jS32OGbCp
m0dYJLy46pWc9PWUjIF+rtumiOsabvQ7EVqRkEWjec4T4mEIo2EruETYLaDtdaMM
KBWA9uPBkmuHnPrftJAPoDfU+oSmO2fej6u3ObwXtspZNf88Bh3Bo2hkZ8eR1csf
/Zz/ahEhQTTIdrFk0KMD/96GyCzD7J7uZLk3c3hYRe0Mq7ZSXxuN5TZAlJkUGIkc
F6lNWdMuek6vCKeHwMKHcUPLzF19yxuvQrVsnBORTRHcfN8UwIOqod8pxQP0I8vi
7+3kmQxV4enGSDTou04of56geI+yW4PzBclxn5bGQ3VHVlQLvQVvE3GrW73WYK2y
1M+bUtyt2ZdfMcCQwFOA9GkekIQi/DvEndFYyu+KjKtHe2OTTWjb+WcDn3Cny4Ws
JbqdfF+iA5qwh/HdKoMTYqo6nDc4Y0eFmJMA0efMSSFt8O8aHvl06XQ88xPvGKBx
ALCweJ6aTl4Ld+4upZxXpGzUQ7y78whACkInP5niL9jlEtY6yYUu86BcC43s4wJc
z6wOAPE0mXBSgk9ngO80YIpZ2WDICbcPnNDvUnuO/CKjmzZBVHsW8ZLSrtcdUTbq
bUSkKQ6HfcweLTDofO4TKtbVQZlfvbP9Fyj7NI5E1LwU+Pbl5Ip5m8mzkE+YPugD
+fA1wo8R8g7XtZOEoH3xt3g7qCFNdna4JFiduIowq490uF+3yb9ANLr21NBCUkYV
BAtKWxc+/ORXs8hDZwoSc6v6IrVogtn5oFxTth648Y5GZiP/2oHR04LUo9HcuncV
hci6NI1UoQGSo0oK30UD36CLY2gXzDhUY+6ogZ/JkHv2WjmsZfk05EtUtxoyka2O
PFrwyYofseMXiejFXRcvD1vn3oP6/L1Gpy7y6LsGLUmcvZdkHLnGOwAlHoui8sNG
decvZAHOf/qqJfHod04cZ8lu9w1HrGAPWo3LAG78cbmNFbxbtZgcISrRUWeLsREV
uJFOXbRSEATBs2D6TfI/Q7WisnBjJkgtN+tljOFhdfO21QppiOxcESFBD7hN8e7x
BB2o8EWs2AOBh4V5qmxSy6nT1I+lniWbnq7zVZi1fulvTe7CtLhxG986KS4MRa09
2n4Bb0Z49aKwfgBURSA1YrGf+3CzzSY6VmhVoafQ6BfSppIr4D4zvTsHeka4zT22
ewjJuaADZ0rfRVzuFlTSRsQvnZ3DnRRfFi38eQNXMvq+kApmR9PNX9APl5pPiR0N
MI5opKZrkNLSnEUzSmLwlNfdJvOMwZfiIOtYo1DC/LdxyYjiAId05mpJ5PoLoxki
0bvvdC6Xg/PvQ1Qoz0lSVcY32+RbDh6F369VDEdzNcvuve+C37CIYvtwI8zS0eVw
KdU+omz3DQoXDlji1HypC/dIRquHqwQyDp6Bfn9EjMxoctT5ekYG++VnbTTWz9Ay
LhUmBsrvtKvSK6Z4EtpINcbhccoiWIj9leJEcHEBtWzvTnDIZNH18QdCfmICA3YJ
oIKKZJKabEpsjns0bdGPbEEpx32g3WUxZ6rkCQDnXDLhJ14qFr0L4IogyiWkLlVE
0Cwl+aWI0rIbxnZ2lGGRC6viJNjIm5GRJJh5iBziTEPF4Duscz2BJFLBoChIeA6z
C46dMrU/+CwzXgoHtGNSky8MG3o9jsoR0mrNvcN9Q2mSZPPeruYk5dBAPaRisrfZ
F50nPJYviC2ZFIEWW93v4F8MGEz0j17R3HUcwuwz6p0ICiInLDSvpi7k3NGXlLNZ
EQ3qeg143nYHJnkTL0r/ixEENaxX+1BLt2h/5smoPzjwWzAaWYZW7479iAeoITNm
n0CnZ2e6wwXtWHv6JaBVGeTkislG5jIDTXVdAyjqxkKK7MPzHbCABbECgBkr/tJ1
uK0pNMjZPUInp8STlm4m5gZ64g3uVGCTd+kLjA598Gi0Zm6/gocsFyj94KLdDJ02
FghWUC29XbPemtUWtxLSnnbHPAlCiRYZMLNSsWIiBFXhUipf1rFcbhP/g9yNr7fb
Ff8StXJ0tTN/wYrAZ/QQ/SdhOkO/9FA2prxNQ1/hHqyl4rTTLhYaK9JYwqgNMZ2b
oaBNK3u6fXmzAE8pECpnV+Ych7WPlEar2z4EEczkIMX0bG2SnLkKTzsPcMXKuVAl
LphnSLAkKDlzOdHW8LGAJ1hTSFbCkayqftR+itm8Ltnru4RmwYK9Iqujjf7rFhSj
lm/Gul6ySgRAq5X5vqtwuVgz4ErvPfGsGLRYE+ZfEhJ+sGwSzElqkYPQboaSA9sC
GuvjvOZ6FsPS3T+/HGldkjIzWlk9sMJZUjTJ84td2xBE1Ih0Qx0G5/u0xKsTsCPu
uGn9MdJDjygtgXsRtngv/A2PzjsIV4vBNpBL8eSucapwk2oC2QYX7ymVLUPXf5Ln
x6lOBLEshn+g8VFiav/nFgbld4Fp7UCY10o+GY2u+bi0AJQ0wEf3pfMex+5dtMZ7
yfMpNFBh/PvzXjmjph1y/aI8u2phAnPGR7i7pCFIgGL2DeDZpBXWuA127HLUq/5N
FRGLRf84O6GPbd9yk03ULAbAsF2+dhD/WMiSf7+oJs+IFzCYo1YeiL0iRigbzXuc
Ddkq/Zi2TQ8LiwioWEDqf6CEDDkJ6e00Ucx2hlu3YG/ldnGxM2bARuzJIBiWk2tO
Of7NX8K0o0uEp55TFHvReb1gabJQv3HT+S8eka9Reg3kS+oeTynZBgmEaSFHrfaJ
cNY50GO3LRFZPrOwuo69KDHH/l27maDUAnBaaPAvc49DKhp9wRGmaV+iZZDjveNo
DL0dRKEdkh5VbzJA9Z9wPoZc6GW9y6APXdCEmol98YI=
`protect END_PROTECTED
