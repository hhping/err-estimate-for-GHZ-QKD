`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccJ9Sk0tmSvPdl81/hcXMSaXWC/rfIWa9rnSIowpE4+9QqOxaaW6NMzwsMPi+djz
118dO3SeKlED2gmDLafVrzdPlvCZqFPbmyLMAqdsClkrrNRk/j6qP2izvCS+6bVx
lDSR6jZHfn3o9xKRHfGgr28VCDQPKq7NakrJVnvSdVCUdjoQ4Ke+uEegdIXA1/Um
jSA/EEhT7iWGUBb3a6T/KB026+EsFxmxH99Z9oFirZ3iBHkTZvoJnBaBXR2S0EA2
TmkhbkDm+lV62TTVawPYE7YMHdO0Yn03/u3n8Jg5EQg4PcAA56LpmMlKZWE9Hk3N
kVxiK+MgnuKAer330atx6kMPG3tffA1eo6+mpst1Cwh9wrYIuG86iA7XjB75SirY
7UmhjPeguHSi/wL22Y0P8fzejmHa415YtbgJwfMz9jxHanuCuWAHhtyDS27KYwzx
BWz0fTPPi7SyQx/yasBbBnpKCVuSp7+tFvg1Jmp9co0fwxi+uDYGrw3lYhiIjEMD
S1GVPyMuRAiOKo5yHnzBW7TF8Eh6tncfLDvJeLfaOtnQl5dL7YBQUp4Xc5Wd61cI
FquziaJg5h0V0F0OmDHETVOyVd3FxuVp9P+HA1FBQa8MsOGgzEjIQThm2jlb5ROa
o3jQuhPSTJcFRXkw8scqfcwiWIq08bgrm1TUPygZzXJbBVpybKIC4eIDTMlyaXZp
sAkDV7ssTHxQ9KUJk8CmrToSxACRk6A6Esrprd50wnVjuBsst5juz3R+VW+FmCJP
bTZLYKoST+i8tykg52+ERhGuRRWiPLiciJnUVXtXZRCB9Lp8EaMzo1yk0U6ATI4y
tRV/gIloCaEUN3yQbbFfIW57wIMFBwvS0bl2j9/KBT0hfnIvUvny/DKKvGKEzZs+
QF8p5lOihLo6xXXNdNiJBZp5h40PDmSB86kFXeUlE4J1ym+UY2/U1QgPkRISCRuv
fzoLi8FMUru2Sefp+n3+rTQKFkEI4HlI1TXNNT8q7UPqx+1DWPhWj0k3M+qPrjNa
EUrGBE6Gu+BY2hgc2rn4ogzK24lwwFtSDFQLz2ZpwVt2wvITOzeDpDKrS4i3JrBC
mNV2AQE6KXS61sDeIJK1AOuLVVqr0YNKCanEdPjjIqVMSwPz3HMSVGWlKYgu7Nll
ctNvVByx7bHN3hkkiIOa+fl2uNPYKtAf9YyP0ZIL6dwbDz40MpMN4gEZbl6JcM3Z
EDRRSqokba6HrBS3dethbmUop5RKEhPBkB9H0bsPOrTjLXDUoRfmLFd+oRwqk8u3
Djk+1KF6pPVG4MjNEA6h5F6ymDqXv6L8y5qgU9GqXGiJ31R5c252AIcmKS2hsGPn
oqJ+8CWGa1aGGAhdT3/0BypDrAxI6RSQ3lP+MKXidMCNSiyqvXBK7tXG2WsJ1DP/
QER2vO0mbKR3EaHSuVgQhSeeGwAOre3ncBqoEp98+aQ8ecTohDBISX2NFgZhiUnB
rjJPqzFsgL+iApSiUWxEFTGMU5DBd1TlviFFoNvtnb0=
`protect END_PROTECTED
