`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7f5QYaK9INCyJmuwpQh3KYXbDTUmy1kXbsM5TMuUNOTwnGM0s3NtP4eqC5ks4YA
A1W8K4C6j606xW2C8STWYFkmaBaASWDQLPaMaXDhkGguDYT/rcMNggvDSy2x70bM
Gb2NoMRMW6wq6odAnRxh3zDzPxwmJS3HEaFlCxvo2GW4Z8eOObJBo8DqDiAgkIST
VcAFsp7k/NWBvlbxaKKHNxmKiCAclmnseI+VumCB60rcJrgDoDo5DH/wwF706wIp
X+a3ajN/pUsSwiS4JfdbNqnJ2BIPk9tXiWlQ0MGGuhkiKgvSSzvRCXphfd3nZjku
zSkft0of8a6WdrD1QppyF5aOTKkJ7iLBotclgjYq2Mjmzyg9cLrM1X6JOgiJXkad
nhEF3rwaeTJy4B+qZ35SIytKvjlZNG3aMTIyYcEUgdKfdsb0ynvaAS5cIp8ApBO4
gv/wGahhbjlQ3ZC7GzEFVvtVoWyjLeBzpj46TCXPzwdiAlWf/iJE6ld/LxrQr/Kn
W/iJH4e2AV/H5BGCS0vtaG5VqDqIghbR8boV7eQObXkS2Jw+UHZkY4Od1loeR+wp
TQaCoSzJuKfsawSe9ZNnWiyTFKb2L57GLbTyBt+69WmdOoyXUB6KV3wSNKQ5yVf+
I2M1Hggp2recIiEbG8gJgmuMIdmplfNlBHyqa8fGY/ZuCuKzi2Y1vhlxkC9lMg5O
lz4iKrS8bp6frC2lOdNc3ZB+zE24dpLVcj+qBgiVfmGjc4EP2OD1ZZC3Be1+RqKs
ptHcu7LKqQztPaghP57cBRtwBzCbho4M9zxBXID2Vjwzo6cn29PRhoAgCJsrcccP
qFc7rQbPrEbazxmLWonicLxrHb6hy2nlN28Zm6vEUv/NG6MvOty6chMpHSbAxefX
qPLRuAu+Ob/SaMpy8n+mwdkostS68wK7Ql6dUP2z10f1CRWGtWi0UQCiu13Cz28m
jTXc4gWHWPh5/RhffSPxTSgxcaGwFYlwqSYFfoP0R2qUqubxuC1Pa5oVS5hW+FKb
CFvDwKcWL48bDBXQFczVRe1TXZezY59XZHdFcT3Uv1xyqaqWRa/xIFHMVq7sAe2r
utYwzLfrzTmpQqOZJXp8NF8NiJtt+w3AEiowCUzwx1591xm+WPjh76muqegxexnW
rfa4+XHv1Fb/qQFH2r0Dm046bjkyijMfxJhXdkQwqM5p9PaPBijNt22Hz2scpVyy
SH5RXv1YgQpEEDej6taKuRRJCzxp8C8BR/adhKJ0voPfrpgmLXsHFK6nuIb1ehj+
SkKIEN0NREiuNY9gDdz75wxHM+Kq6llY50EAR2sXTkPIr5IaC54XraEI0wO7xYal
oGqwFIa9l86UNl9KXaScKthQnEkuVoFWNbzHvXQu2g0WsSZkcj5X5PJjSntOGswE
E+t7giS2Jh9SYm0rEwRUkLsZatXngbGRQAe/cSb8On3UY/Jlj/5FuGim1QmGd+OT
3hapbO6T6KVDjsmfyRPd8jnYZrVMkhjyt/WcmXiakcvdePeS/t6+oSmfamG+r01t
K3obAFFbbG9iHaR/xkDhhxlbg01TS7NMLiqNfPkpoqQUrXuBxyaNs89pXL1Waql3
NoSv1ekg3+nZ/qZpJAtY+1pbVmZlvXQBO55tJemzEYzrJbY2yi6XI4e/dzpqBDet
ytrtdiw3jE1g8eZkGtJTgt95Y9VU7i9zJ+EnPlRvQ+uRDEiAwrQ1gYAZAwM0AiEX
uhAGYY/K8nCiamkfXa2Otn+EE8ql+PNk+IxeI+SS8FWJ6VwPh+AKjqeP+hP/Fq0N
njRPo+HXZtfcTNJ2nXef22UXAmvNXWwXeEXxT9iuuQYji4LzszY3OJKgsDVIAYSd
7RJLaNKG2tIiYBfpUCV/L+oAKNuTos/1R9YzqRVl+h0MDRit3UpTv41i+kL6qoOA
5RgRzd1NvCun5gIMfku3qm3gHpg3ZZD7uBPz2nAZ9SQytmTccozsLuJCzdo/TNix
EsPKlpbZDNDqfv0Rjg/uq9QWrFDEP7ucBltfE1v8+IdwiAtr5imSDtoqzmg1qsfl
DajSqoR+QjJQ23btBU+YW5qHb2z3hW6UgtoYg6EFpOJtsvzMKM4dV3plfBPMLvlu
WXwW7rNMHRMexcZrhCYkEakkx91Io54g7kv8l6f+QwT2xL7bR+DlksGrunf4MhuM
4V0vLUU168yd5KK+8pYHsnVV1OglVOLMzoQiJjffekezbMOpPaszxfqnmaQ8Uppk
hIWf2nBJ6SpxUroWLlVnuKfu/PamKnGVzvLvZfK82UL9wLkEsbZeW/DYZ9SpydNt
3eXrjVn4wH7AEfmIGPp0AjFf2j7xdcbMej+4U7WoE+pq5KRY+H6u1okoFxzUU2he
u0Qx5uGeoCc2CZrSs1du5E/hEoIbDmw0xBHVh+q4j4F58YyArqaq8V7J19VMdW0s
JfkYg485FhurjyLPLENpDd+dx4VQI1OqIBxbWiZlZlxV/4b2H5sVvq7aidzo7f0w
VVMbY3xJo2K/mLlGqo9OC1vTTTYAwf15g3O7qT3ZIG6cZuS07jQYmCqjCJBqIZ5U
BSTiZBF/FFgj3iC6fYFALVkEDPgYyrIufJZpuITeXWc=
`protect END_PROTECTED
