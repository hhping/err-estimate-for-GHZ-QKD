`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G0ugj6rg28Z0VPWkEANct32nkFjnUPP3oWeSkm6+4lc3cpVxO7FEnAGZtiKOYDVY
xGsvTyHX4PaVQLtrIxJCGqfk0KCb5NBeP99+FMKh+5bEcva5+U5sko1FAptoLW4M
gqGIOlfJCgwB5TceeNHMnV6qmcjJKtLAMCXiyni4N6bXTaKsPlWqCPEqhPURgC1v
61mICiZ0vkIeC88Gxf8kWcX9wjrvorVlGhN7Ug5cXBPPfQygqjS7I1re6Yqa03Xu
LoH4aPohMepkOsewJJJsPV1nkSaEZvhs694HWgwqUJJ7cOQ6LztbT4FJ+59cdTd9
b6vEhu2vTGn+mJUzVD9VA3mSnErcKNHSXUTgUH1a7uCF7Ao9/epBGgyYtUurxy9e
pKDdh00OML+G64pQnbiCI40eoLeVkooUpXQSl+i+XIR/Hxp7V1vEqxiqrlG3uAwf
O4nokJhrWUxCB56WrVjYG1/J3JKSpB3fRh0RnrwSVzWeQCJ2KAKQvD3UL84OXByz
FqzTtqs4a4YRaGdR+CW+bydCPf6g2lrywdH0avnkZ5p9vY8/Di/GxLXCO34MHmJX
itpFT5s8i/Ee1v50Yiy8VKodcP+krofT4bL8ovX5fHKvNgwsZU5Wkc6w8WEPoEor
3w0aBPQMHl7jb2f1mMdV2ais5jdxvtMPBSepdk8d0YVlZ4PC/LW51ddsAcgjYYWG
38BVkyv/BIihD7DJTS8Ft5QTzMNm9/TqOJddVvTgFOr4kkwx4uUz0ZYOu2UsAh61
/jaBspLT6MhUkUCNp2q5poJchoFiK1B8YOTYxdBUIJLJ8IIS/t8KEvckd+YlOm6r
KYN6pAGBxVttlTaVMwk7o0HKidgBpiwiz2JuifvUEoTkoHIoBQQH7KAul/9Yt7ld
n6Pr/AXHAzpvILE+VvGkcVSDDhWa+YHUfp+0ZkyFp2RYXaiJDxwoCXLKpf6Ola+B
MoYTnWHRA/8LmbtVtXMqnqQ5RXyWfz+FpGTwyz/6XD3Yk/y8uM6HdNT6d3it+9c5
7KPXoetHuJm0w8cO8uemrZQS29+50UyYL6C94hnh6AJUix9TOKNoHszqt3iUGc3M
CQh4fcL4FLRVEBK8gDHyURLxlAJsXwqunYHH91Y8CNpBOwhNAsb/DCvGjQ0VHFz1
wlJk6P+CXzEAEd4PrabB+/2HtL9Vfm/PieKdzKiSV4EsMx+sN7ragi0jQufGYY1r
HzvX05LyrQrV+s8WUOIkmZwYq0+KIz2IiRqqEjFvUjL2/Qb+ttxF1E2YjNwrNySL
8D1iWIWSM+wN4LBfd0/ZYlmM3EHZS4VAAINzP0/oZn7pRABTCQnMH1trIhsAwn2p
VdOoZmQTVtCJczl8BGEoTGx9Sw4B5pA07neAzAhoyWcYlh3QA6TR+Vi9uzfHk0vG
7tHV25CUWJogwD/moBjXkGSwAb6HhJ0UA6lcKVQmDpzmiuLSmbdP4In5TGNY0w4D
GYanQWF9FFkJIqnCUlqq/Kjt0pbJ7zRleew6BoLV2dZoK6h5Dgao2wpmVv4ArvLW
C5vNxZL5wZr5j8INA7/X3nx22vpfiRvrQWA6E3+SQqHvkJkhNHKhVGgosLPiGmDO
ek/XnPH+grG8+fCjuvJ7/uGovP5pKuQFBhFl/58rrf0wXJ3+pBIhi/rEqqf1qEPf
RiGuNnIM+aTSsHR8A4Sbd4b66lwgRWNiBPB5DAeJPEas43BsS7u/q02iDrST/Dx5
wO3PFisJ9Buvv7IgIVPMsAX94Qxm0J3I8DKRz+9AOJLWkCvGXs1K84pVgybigB2q
2i2Qz8Q8W4fUvaBzBKb6Tr7nXo5vog7CWfbxE3u2opfz9fqaqh0L48VUnk/8O2fc
8BfQiXNESwaDDlJM7YclqLfdco6dmOvnxzjmES5IYhX/Wz8Ls0XpGNwNt0cwDXRR
XKO9axdW8IUbLtwsOOGqaT7F+G8aQ+fw4TG7PWaVQwvA1Flsz6H2GhMSW62alhWn
mnQAsTVbPflYiceC2/AhoBo5n7esaoElEeFdYdPLGss906dYrNWhmETyngaB8Vdt
r9IRwfiNzEBkHO7hrMDRvkHpx557K/R3NyyszQBCExabirobz9dMvJOYPhU6DgwD
B4DyAoyMx9muh4FUKYozRJj5jCvzehGEdHOh0CiqLexOP19/Kbpok1HyXYLxc/4+
6e3UNqjqQOXgRi4/Ig3tjJMjJZpRgeI7BGHot8WjRF8rhTobQjT+ZJIveqD+SqQF
QXNkRo7mvSD+heDrkRd5cLywhVWHXZsb3wbxz0bWiXLMK9G6+Zg1cZTMCm0cKEqP
WZb13UlJJM0OIQQ3OPzKOeoLWf2LH7USDf6F0G3jkYFmwy5tzjcFxQWSi5EAOQi8
cRphwuw6jPCRWoRWMNaX+OJA4Io10TjCTld2fN7c4/hA2c+ZfJPfssqeHBTEzdhU
TbkXzARTtBCPdBM6rDgcBg2G1zKOh5mqM6cN9K+rksNco0pV8GyVobYe3jUdxRj/
1hQnSLQqW9jZlIpNXHEF1YDY3a0otm5yVZUZtzga9NEqFwLcRmX5wgOjG3V/rSNq
rZ/rdyEf1LKRxDvx4Gkj5ulLnayXkWJxGQxVYQidkREj1N3bcvF088krmV6CvEVi
7Ww68VIlXvxMVvZJ2EIchkxDkn0mgvcs4U+Ka0jHEtYI7MWhqvlbc9Yp83eOW4dR
+S/eV1+6f1R5pFOvOWb1CDCzDZPQDfC5jGK8HVAFKX+9c1+wbbAG58j+uus4eF7D
EhAd6lrTG0nzaYAc+GwJhPbUh/ZDjgS1xaktK4yqTccRMpqvGi6PadBsyfTW1aEX
4seMdWzX+7/Bx8MnZK/fr9bMYcb3+DGHLsXTzGFuNYl+60Ur+3ckzvs/Wg1UymLU
QGmQG0xaOkNlhPzgGWOdyRK3XNsrsCTl1LsUUzBHIeaoUIyK8rxZZ1HB5zmQTUEQ
LDGNTlbXIwOWt0Grz9zGzLj+VPPdhhon70wgc87vH4mA2KdA5D12tFp8TYGzcmPY
r2uDKe1cpuHH7Pn4jRQSiG8U9TewUsVNWcsLpe0zxWdD63PSKncvMQRjXhpznTQH
3zA+42kQ1Mih1FvRLTHSKCPFRwCuxRfoWhl9YS4ZveHf6iyzwU37uojwzccbE/Al
yTbSqb6I8vyPe5XO+PPDjqKPC5E8aiIkCFAl3xwJwGanhKy0guS2Rj8A9oGna7Ys
IaO+97S3RbyQRKlE0Id/jKumnwnt9xtziOXcXfOfBmpoaVwyVEitryCmnuWqYyhI
vnOEiOahy5ht8dlAVV1VoaGrXd1BISbummOauRMX57685teMkibYSBMmrARgLfbD
wNJYkYvF8TIt2+x+qPeqmX93EnREsJHsKFkOqdm3kq0=
`protect END_PROTECTED
