`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6J6VJdzUYgInJEH+xu76tDOwvGTWKPBVErVY047zyvivfxxhIPIZa9G9lAiQ23hy
LSLO9TonT4Eoy5M55dvs3HixfQ8Xc5P9Otzhm768LYShZFy3X3EN7Yy/7y98mqNR
OFskLRXGt/FjT1UWufWNwyCROJIC0WevV+Xjg3OAlnJvGxnvQjQboF/RjOH8W1DZ
AkwZRbCLwtia40fxpJeOftfJytLgpumKDmuQaMV+b10uRh0BbTFyjJmpBI3iawdY
zV2dDVzsFZgZ0pT+51hECg8B6WFKIXiYJx7R4E3WVXlk8/Ill07fw3zAPSUdkLAK
OmpK7XSsktwG85Pnyk0A0QhcJe9CwqCeI68cT7MFul2/4GrzgTY494del/6lQXuQ
kqWBBLt5IvIdeB7M4wDBoBF8F8fj3ThAxT5C63W8ZwWy2bYawfiF+Ng9UbRs9vRc
hrevVB6Ed2l1Hng0hxiBhlWuQrqJxUPrM/bADMI097xEDvuuH+yAPsAXHx2Znvkq
o/LDIbfaDML0IkBZL2upy+F93zYjqDitKQXLijKvLcYo6Xk/2wikWVS6CRU9Bw7x
`protect END_PROTECTED
