`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNpqxw41qmeRcoKJwIq/aKNiNnsvTnnw6qlrW5Y6/gKSisnDY9d5aFpUdq3x90k/
/7pck97t5vN1hyAd1G2aCnj3vHBbf6nLvPbNX89i+iKh8LX3uKNYcVPu//4Kqt/+
4RthoSSH6v3CnBIs5qG3r4bmtT4rLowMoQ6NqNshhPAXusb51A5v3Tb3IysAUPzY
6fU/5qNDBHjTuoNfcLWIHy151qm7kCuaT6wfW5N7BGdZTkRgqBDyxOQmIxvwWcrw
3wAF1EYaRvVe8645SUzv+Cq7cb6+w6YXJyz6UTAwQJavNczwPB+vqzyr3El6T4Pj
I2GRjSLOUOnLnCe/gu068wbeymgViYuFNMUTAEJdH8XhocF1TBG4yBKHUSzZVYDf
+pRi/Dfibc3eUj+OLBsSZl1YUNC12501f/eaHpZaFIAGkKUh7bhWlchazrVYE2CV
y6uGweL1Zdu555m7mfMQGulAaU0WFl108et17AzNJNRFPhrM2xmFxlVK85zFmbHp
pyiVmnxsTUL2JJmXDOK7O0obBUWNSzEa71Iv7m0xPAic7gvtMYYbvYCfdzcAL4se
7V4KPRwJgGANkkddsC0DnTfzwaQYLjwFPM5A1PaL90Oq3hm1g+UF7BDsy9S5Vktp
0Uhq7Pq/2GNEuw0HhWbqKrC45697K7a+nmOHlDY+z0VwPyQMi+QaAoxBiL0o6+t1
OCr8PNRLN4iSPuRA8AA/FK+MXfrvrl0NaVtatA8vFMR1oWL0wU36ZX4G7q/whXu2
2fEJ5j7tuiC3d6lKND/LUdLZXnI4Th2+vYX/uzjHtf+7xtVofj7pLMTP4CQGErq7
iZHM7J4jRXx8ZyRDo6zodxu27uQjfaFbk5hhGdAi8rgsXwPSu8lwLqG5exR7sqlY
CG5wq/PLq31NHtuGb333kiNpFsfQ5bUjHCRmJjVqJ9gJQ3JgY7+EDw7vD8BLJEwH
/swYaBK4ApBJP4OmK3Y67n9iGrjYrq0dAfrB8qcJTew2zdLRoHoAqvvgqxeXhSyC
AtMUuLuZcfhTK+u7g/7CFSHpCmWkWnAlz3YDDzRc23AqRKsERIcGUoeKwz00wBFm
jFDmFjU+8BrnyIAgYLxoANlJNlwN2dj+5rKB7fNp940icJ41ndj9o1dEBXttA3mm
jWyyXWSReYObd/LATIu7g5QWvW0qOrG1Y34yxm+s6hoPkvRT65dgUdt0per+Hjbf
N3gbGqeZbdSQ/TEcL5YWg0DqQU4s86RKujDUj5IWvopbyf3yIHz0B5/YGtXfZqxy
o16XRW335MBTNE6Cnsa+jxAar93s1MgayT9XvDTXiUsBoolfCbmQN8n4OM5QDlj6
wKGErbvN6cNo6NPKJvInVYBELRJNZOTf2fEi7KL9/iyOwZCaplfQXtG3yT0j1yCh
a8H4H43BjE0OzAAOB7TsONsf7kqIafYgLg6yaxJcdR4a/5CVQVt/WF/LoXXTikm/
jnZV6QNSzRgiXb8Tvn+CoWZwsWpcJJO9dPFgd1NfKqb5d2/FL13lgvnppN4ykTDj
cLVxqDZxfsnkykqp9JWeaTrMxspKRMLzUS1YKfZshW/VAh2CA1fbOM+jkDS7YlE/
fS08uVWbHjYqXoguWeaVU7JM3PSsJL36BiUMYi3lcnzYGu5kLustd00eOcyo/O0c
JcJdIvckWbQvnV3JRo+XaLgM87yp7MjSes8G/9aOA46h1Kui2ZZ1DK4HMJcWUOIX
FLFqljqZp5H05F5y3RbPij6xv2eDm9HtW9nr1iWOxIgAjfWBPhwigcHiEBq32BZD
CxT2YJWg3HRYkOG9uKFxLRvZvWwB0/LEkXuMFjKNQ/Odvs9b9NuMZpDUGfZ7x7R0
Y5sM6sFHbwcRj2wGOgbed9xVAXXh0KUhQziLwoyRtwmwzUnOfUKavqP3ZGN/5nGa
hzG8bPnnpkyZEX4q8nWZN7shBc+Vas5sDMMCWhkigWwf0SNCskFy604AaZ+iS0cc
nrgIeahqVM//rNyVzU/Q5INtSgjsKbrJw0F3Y6DJA0+S96bBXf4XCokefRLetn0Q
GKFQ4faeq70jHXhX1c2eyeTG/RXsbPN2kSV+w11fckrcs4HcgqorWFSLc7k8omp/
G0iJh4bxg5vy47HGk8xJQQt0vUGJFa+C6V9olcMXV0BoEKsRo62ABiT08YAPdX2p
gblnRbrkUZWDs+NFLoe9O24AmLBousPjSyQf4cW1m+O1wueqEkh/0fF5DH+bjaUR
sXMALzt6qPuVRCZKRsWgD0T9cSfMQf2fy9wc6f73HBkW2Lyd9TXLe494LyYI0MDB
4Zoc6hCEXkJLtfynlFdH0efk7GbwefYUo8Zzcg+7R4KtUR2nVR3qg95SRv6LsPSi
Sa+QB8IspIZ2IF+rK6DOpWG3SbtnWd4dImAb4HM+RhSgkqeMAkiY1hyXuaBs8pun
NaSmcYuMNtHadod6IX/XDfhy85OEq15DpDJaEvpJEyfIPJyrmk+1+9ncyieRRc8v
+zcmIelWm5Y3kyGx2X0nzjYm/yRYFTwDBeZR2TVJ15pgSEJJtxMd0w9HTKpTeS9W
nGtWWFKlwAtmtKsJkxWhyGrmpGFxzFiSYhA7yFM9yOjHEIjEK1n6SMWNYjcAmnrH
xtL2Zc7ce/QzEmQUWEaJgQQBKujcaY4vEamKFr3lGSO1EyJXj6sR1YQfJb9CAbcb
kBQckZyM699hK8RgS4tAdn1LKiXfANJaBldNcoMUyeLXQhxJtEv/2OiZcFs7/Xro
QN5h017YEqoTqxitA6BJJTqX9k4hLIgf6qiOcyFNHnL4rKo+tkxLGyNbXR82iQAD
OG3tlFJMWEcAAAxrtjT5Qs/fE69SZJWwlTr7saN581cfI9sm6j+RysJQhHdAAvQ8
gsCi9Grb3IVXboM1azVZ+81XN2Ibm5Esi2uho1wlsv8VvXWVZOrrz6Q+g2PLq4MB
Wpjx+6v8BcCm/OGqiT+/SROsA0fPqW0sZu7pD3pxhaLaa0rH37Pczf7omfBIHss/
V6b/q/ebs2wVZwA9QvMoSBDmByfUBxIT6Sb3xTYcpXGm0/TCV4dawUBq4sD7Q7MN
2QoQBDFvgarGLftk0Cgc5J+XxBjjUqAPCdytTPhcGaXJ10zmFnh2ciHF4dPt5XSW
MZ235ANQWEMnYfPKYOPY8vgQdcArq/DaHEr0eAbz+GtdUIAanY83eP8fnfKkYqgs
6qrbDtEwldBVrSZ9+Q39fIh/HIvDLLjTZH+MBkeYRprKOMcV8mPNjOXBrUX7nSke
AVh/H+An0YUnLExwgA48LIfaElxhNr4hSTvoQxf7Zm9xXgq0zzsEhdHaVZN7Z+Ia
gzL0BCgyoCLvIaPfGDRO4WzMkTqomrp9fvYKhx+hVHZldMYYubZaNoRILNMK9hzz
2CbLca4Q2pYRwdTfImGHEay2zNpEdV5Kp/sncQrMVHwH7pYMcsXQ5fHU4pwBydI4
rA6CI+wt2EAxpYTUeAqa+QO1T1Nzl/8RZPtpmv5ZaDFc2BWXLHk28Wa0WFgfUbGK
n9ssaZVEyoYiP+DSbODzsGp629Ne0rb/yARo7v+IZB3mauj+utJ11rNJ52ehqP1w
wy8P2UQxNU885LYUNqvP7rGy2g56/qxyDKKTitzYcJCgyzoYEky7c4VjIcZ6XF9b
iQM6v6iT+YQ/XunKd2S/GZiDD7ldLhrTijaKgCXbRTwasEOvNO8xPS8dfnoMzV9k
05uCoA63kZug8sB/N8kT2LrmHzfTw0cA6V2bP1hHnbcj/CUzPbF50xbijudSVA/Q
gYJo0xFYwnX0Cpr+q41V0dIpYjzdaHDTaIUicp4F11JOvS6LoEjHRvD1yLeYRhK9
v2Ny8eOMzbsKJOdsQe8kWzpVR1o1OEVEjU0Zp9A1l7SJWd9L2lvYpf1IjftE+ndb
O6QHOjo4DDgnHQqWqCjFR90UX8oYwZ8D3hicth5rrRJL/XulJCtlHG9Bl+ooQxnh
wtkXyDZuovZlsd8B+c283xZC7FwFReFBuMxBYcFoGOW/LzrWpN+lddlHNOrNDK7c
pTi24b30MC1L8049Dv+Ar29ZKONuKQMT6rby04imcjI81xMfKfWawZCumcWj7vpZ
2j/EGE6X4u90wm1JsTASduzcAKCRpk+NfPAv3Wv8HrQ=
`protect END_PROTECTED
