`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9JtHMN6+SkIhSxFWTxE4uXq6SdnYHVpX7Kz+Gg2fOdIjNkak0TgxYBK3nGirWeJ
Wi5KhJ4ynpMu6DHgpFARu5I8K3TgcWMK+2Cn3w2k9ARhP3+f5IzCF1EBhaOdQ5QL
3rqjs52uw/JS3LjXGRqzpJ1jU3zZqtayeUFZhzYVTuXfLhFXLnombhLHzoDAiblY
/2TR6RrapEAKJMIfcC8tX+NAf7gFLwKcj3+czMbC14q3VxRCnLEHxyMa560HwejI
LZpGcPSWRaQ8taIRuvMBGNgpSVVO0Ix+njiZiyHvV/P0/AW1adAtOXey70qUaDr5
hdU5y8lYrJ0JfllBWxy8AdM3yVIMmqUmOFwOWVwkiRBotsGx+lG3yRO9uR7/0OSK
BGwsf3yK2CG/MmA0aib4AU0kMkgUe/B1UrophGKSfEDIUPdw9QJrgSuPTyh77X8/
ebCVn4JFX7HxRGyTFIuNO5iXieS3CM0aWA1NEc3ZAi+7Uf7DQ/jdd+j+j3Ofnvb2
A9LBDx41YzD3ETjZ+QFjO7BNwnLH3HRSaYpPJGTOio9lJeBryefQA37TaDgWQjVI
M1WUKahv6u69RLs0uEWJtOiuP5qwz3dE8OWlbdoM+wvb9SP5YVu+jmtcmEn5M+9m
/yNLrhKvxADx3jCsyCJDAm+ISyO9IEHj9r1wIRiytSN+7EL0mSL8Sfk/MueukYt/
TjN5ZR+w9eDL/AU8xFsGQp6yAjgmwrC+jDF34wPDrM/s90OUHFdYHI5X9F0NvKiW
ArOh8GUiYlynhYyOb/Cxvx9AA+zcvRhFULe6+x05MX85yz4YUzKO+rxoMbMOksne
BDb3FIMkOfzRDhqLBpKRblrPC4iM41WXU2UV+0+s/mIbC2fpiMD5T54LgLHYCg/4
2/GlkxKE72lxYcUzq+RJy7GE1bQDE6hLPGPSykSm9A5P3/dNzK4uagOQwkCEJUc/
B2G+GRU3WtvURz7Ee+TQk9fZxPbCOj2YeCWBYEpW6KGNJ4ky269u0nNh5VxW5NcI
`protect END_PROTECTED
