`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qwoQZn/E4Lhj9lUzyu2A+aIQhO77vqCrZmS3jxSvZMDQF1V8Q979Xq4AvQzNdqtI
5n80f6biYV92bwQPLxF9nDKIK6KkERYD+QM+2MFOp8i98DnCvVPXvTjWvfZ0cPmp
fudlF+0ofOt31ydOLlgplC02ItDMeeuW3We4KgBso4YKZmNUsGXyLjxRBhieOqIr
kROx3GxOD6RUG9xmQDieFL5U6StaQWNmZ74eSFmJrfzHrW9JQKdFuEy7XM00YTlN
FOEh5SyIr5BzRdSvNsVlOj0xHvDo3i4lACta8IopsArURGFn7rMcicYu6Yd8+bkQ
20pKBSBIyrhWq3y35rG0HNjvRBPTM5XkhyBaHLngiNs6PRCsVEIrm9pDhzHkHK+O
5mWKitAXfrSUYvGpRFcmPk7H6/g8ELbQ94U90TLvRWyq6EBJmBrQdrYeWjIk2Lza
w2EEUHPxfzGYtfAN5VdLpfo8R2O5TiXhyIBgo51MDLJcApGVpbeMkDsVJMH6wZYw
I5gq64T2CgZ8E2oRF6l+RLL+vPcWn8HjwEpMdV6lEQ5yLR3N0xRM8/YnbbdRg4kU
1V17bF7R4CukQ5rf0awOjpzMPaHLJY24TquiqGXhpsmfeh+FuAXrDmnD+YoyMOzh
YF7EjgvHL6AoFb8yIXRxF/XqWuM5t4eEwJPp0r0D2RJTy7HTTwlljRGw0hQtHqDR
xqu0S21WwnwdEkDlawtcynW4NHvsQ0Gg3nAykYijA73fupl5Luwxb3IRjyNWnRLc
KNRlWOrJIDH60yZz0wXiyLA54u+t/4XwTp60fY7bbdcDldmjJbO+IrRByE6ZbHnV
P9/L3oc+8jkdBEq2sIJxAmNk6d1AaW1xtFhenjwUmDi13vfhNaf6hWxY8enbrOId
eUJRl74mFACLZcWLnhvRM3tz0IHVPnkhAIjXdASUOkbcT2iyAiHSjVdVkYH6Xq/c
x2nGTqGxik+5EVIt/Wuhz4Ti45B2KPZn8pQIgKki0KQ7Ihk2EiBO3P1aJsD+AqRd
g7ygJEx/C90Ht0qgWRAq6RQmm848cJmRiRDcyVXWQguTCwvyFgtOezM0S1jFMaxi
6f7gNqttKgw7n6nUcvuiskMX4jCWoLvpsPX7Q4JxYEXie+7nr+IGjaKjwQJiLwNZ
ui6y2vSzyScrquXj92+gH6L86sEpaMeyS4yXu5RvMUU=
`protect END_PROTECTED
