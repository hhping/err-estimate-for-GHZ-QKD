`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gx+k9eGgXTTLzSBcW6lY2uBAiuf5lMp+LsPuWWspmeQDobH08zZ7TpRmR8GIjdk7
zEBsydKBc6GTn2U3l3ViC7cI1wN9++WycoiD2gqbOcQTDemuNyPZXz7UwDsfUv4A
8GLoSltAnt5+N0uM9WrTsS3v4mHIO1g3idFTGKKA0I+vKVjXNMga8OSkhlGZyLUW
X5xuitv5eRxBKDYRJ2SBtNcFKr4fTou16OXhILx4U3FC5aBh8XniG19zU6+aGBAC
nZa+Hf+mRjtzMUkp28MrJOgnoC8zt+QMdwFmZkuoapuf2/lRKW4xiRYWQOqz9HUn
t+3kd5b8LYgJ45Z3292UK0ml9Yo81wkwKkfxrFBZMU8Rp79LjSHEI3B1MS7dquQW
QIY9CVGUAO4MEvz4ixDbVPrJsIKoO6Sp1zsVh+rL5TBHVG+mOLb1ndhZ22L9hZiW
8M6NOlM8uIa8wTD9rMZ8VfYaFiLihMIKXzsQmbwnWoIvYM5kLq+PQYrBAmNEDq0/
bcFlvdMGZB6HhTNVO2cw6KT3umJrbneq3rFUcT6YunAw5+i2PEb9yM+v+6tA5DQK
SEG+fyJHpNeEazO/mmQimUvuZo6gszQ9DarqH2Oq0tqmcP1WpEUWGSTdoyJK3BF5
bqRSZOLfAleIu1IVproAG6Cb+txS4a0Cbvo5hWEflS7IpQwyEXllnhuxiHHPiJIn
7vqeeK09DKF3+K/NTPBe9oY+Dx5N/KXm3SJznTnVKI2zTsd3q+jbZHwAC9FMcTKn
ogIIT+GzT7UNhKU2SMFQ0yn/F1nvr5AXQ968pA9sRGaKe34cxHqzSiQGIltggCmZ
TxATbSEXueCUHynF26AGf9++Z4WO5LMd2duSHbY6qo+ERyKCNZAXpObzJRDcewnB
k2OKPa5XK9ahoMIUnBDO/WXwdFliDtCKd2NYPyL548ZI6fTYZe7Qkf67IZrz9K6e
wHC8o7FKEU4X7kwfajIBBHVSlfivFvX9CtRS+Zbtu0j261HRnN7Kkx9+ie2EM83F
ZGU4Kv2wjjs+jUx5n7PFiMnI7WGKnnBNM0Uvd86NzEjImhOiYqtWIPEqM0SYf8un
`protect END_PROTECTED
