`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VEUP9WJRdbW3vYghLJAIsa28hs1exf3542KTlh/P42n7pBpHvtGL+Xmgf6gN/C7Z
P3jLwreeY7G77DW+Pw/c+hVwofqKqNsjKlYgD1NO1b/TZyHOpvbDyDHURT6ESad6
dN6qFYFw5DC0oHzRrOSSoLcxjZMuKqD3io5+SOc9YnnDB+kdCvuxvOJP0Nh9gDCn
o6a+u+A+JivBVHsaDz+jUtOxIbi6SnCarW+CnmwJeKl/5SzOzcck1QMK1zUcK+dG
SkuP8jjrD3HwKhOL/HfFQMzc89uOSIDCKqD15/kqDuPLcM5GzYX+ZwKL58PqXpPE
OFWD0bufpmAWcgzsI0kxQSS1lFFSt6KLx+XPHn3jv0nPKarH77UFTZPWpGDQhok2
8Q7grYlj/lKzUixnD+f7rX1foSakTqJu/go049byOa7MGeNgr9Ree6xkQdLEWTOv
0cqIxmebqLr9cL0tn6/+d815iXlCVSDyH4WGxAJd2e0Uh5QxHdHWiz9nvOE67xY8
331LJudZWcihQXc4q8HQ2En9ZMsaaJ86mr28lgoQS26WtDlFkrqZrahT0ZJ1JH8D
tJb2gIUKdopvOf0G/q5sDRcjmx5NQCB+pL5/A49hc0veAMSTpU7OxKREd1mrUD3Q
CSTDtma9AvQuFpLCQl5CworSNAtlTw9AAVQYUTVzGADAXPY3Jjl7XjQmKwcrvY42
DIrHTrWN9Nn5ZkiIap8XnUqMkWNibqRuopY5gu3AhRyKbeVHjuaN5OfLgL+ekBHl
p7oYxL/jRSkE2o7zgg/5EPiKuKfQnFwZWcB9d4VvW+lHzajYzs8F1bi3FX1FQidj
2pHL0YzqlsQgtFwki1LUSMOJKyyvmJiaMLhrDJEVB864ViW9XxQ0nUnUd6sT31K0
CpQOKw2wPb25AdgYFCnv4nqwqCvwRngC6UaDT6B04RSIUmOLmHaVLkUT7Qce2ew6
cp4SWLnEGD1Yx0aGBaDTXYjp9iYeP+t7RLnuIh504XCA0Sh7xKuAJ1zb6j+KtGq3
ZlpP61/RLTRx2DjkvZ5WcbDhLql8yxuDt17ODYSt25OB2zhr/ubkt7/VMS4wLeAu
E7rRnRHHRQY0EZAB208b6L7F4KNCp1rNr7RYwDAXsSfvmVd7yglc2m5UaeLimZod
oCSNi8DYQl5lRzlxgtPjvS1SPokQXYPJ6Q0jvV1U5arREnaCu/4pL/KGUEFDB33T
4oUZBb4kBbUwJ8friXh3WCzfwxJe50qrOM5/FUVByALUGalNgstMQItGDedzAU2t
3qNsXb7J2Zsu8Fuf5HQ7dXVNlgtqFzwUoj9U/LpsCkbLNFA7CXXiQh6wq0UOaHg0
j2J9LmHTLo1hB2lufDUIN1JPoume5q8THFNsdCU/2ivRikXtN8PCUtDmj44K9TnA
ov4vju/C8lPIRzzzfH1Vorub2zeapVjO0lmrfjezwf2KBjezsXacIHQ+/74yedpQ
PykyOwV+zk2+3qVM2qMBHuQ/2t24meVFsirXYmBrSpYVi5rMdCURBRQOzbItG4J2
yBxgQzs1R0JSX9iZbsyIp6HYTBl1iYvGFlahP8v08kHzU8xGdyl2UpqJuPJtSo/p
PDNVG90CTYWsaRliPEyC2XfkMAGubZht8fETGQUHyoPYeWyrX/YlQ4wFtqU1kRi2
OEx6ohQIOR7GUzB2YUifS8zL8PFlrBcL/ynP9eQDyK5gNUMU9BMQOqiBrDz01lci
2HBihx75igQej2pxyhdChk899G3xUksLFOY4K208S7QFFp/cILV0OwqMCpX3NYr0
WGvbBVDVrpmh4FnwUqUdzwWJ+JomsPhkFqmjzkmIaBtoHxFz9nd/+cBTve0z+7X6
hXy6L7oUyUAjp8f73wGr7jWOSQjRBvHgMTnK2MKzUthoNNxPMHe16xVHmYM43qaE
p2bjbWmUGQZa5Rm6rp3L48yygqYqVlt0lBTI5QB+uDu49GadF5kLpyiFWlZoXTUj
eS5gZ8M+PTk710O4FyBFY1DYXnejDUrh89JJ3ca3cgQmQzR31II8aT6XWoOjcxHl
w1DCE2kqulXnKDUqKZr08rW2eD3KZ5E+lxP76lExlJTH+nc0u9kYqfJLwkTsVAv2
Y7nZh1wKNthUv2h4A3SofcutnFm9ZMVqCTrHTcV1/Lts8+sLrUvYvlRMQbILaEoq
7DGMXrhYk3lLVCxavticsb04qpx7gv5Zim0um8aSVlhosAsVuwYXxodl1pCou8WV
GZEoh7hxD58dIDaPxsw1NolIoh+YMb3VzoADzzeR1e27R5biFQZwEIb0wW5tMtPd
E9yil/x6jCwWbjTlWxm84rSNd+KcL63cEx1HDTMvYAPAx1JJ+tnQAI8k4i/14cp5
wx2A9UKmuvkrHdKdVoRRwwu+0uLDqZJVqNnPGe2C4Gg/JDv8FHCUk67GJyprWS8P
0+BPclGGRANR29oNTVx1haNyASEg+R/8KQuQqJMUb1ppY59uSnrz1rVFRNkzzo2u
js4ARAwR2Ljpk3hwsYJ0HESelxDKbL+88q94Xk6bjkl+QbQEtmai6P0JxkTFQ61S
GPLmNueOB8y/KnPfwz/rOS+O6cM+gN5z6SkNvyIVajHwXCXDPRcIPUViRbCGXNDf
A9Ig+zEq5CRPzEtevbdjUSObsRu540fD53PlTRwXUmJqx/075mGSj4HLwDHm0BJW
/xpkYp9X3N23KfHD24gznisQEkN2/zPWQwPovlL/MQWT7dXgKTHyVUUTPAEdZbBb
7+TYJUoger2BqatY9+fU2VvCNU03K/MLNa0/E/CwVyr4/Nux/yH+dSj+UQuLnZTu
muPfiZW1tiVCQ0uVB0YN6mWNWyIDMAb4oDksdhiA5jRMVZSZLd/3GFbL6a55bEyx
EgfPMiZfwuzjz6RI1NBHMAm1YjymuOXz0qILJKeSLf2YTEa38aEDlrXqtdlJdqkk
jz7goMmtpABd/ErN7TMRQcsVTRkHez9W93PK958VLWXxXSVy+BTitZEbNKqji+GD
mJngVazAoQqTkCxsAu4aCrFczsyA0IPhiCVeVDkpmwB060AsnZh7Nh77Ny/ANS5f
igE/jW+jdT0ZQSPt6mUy2tY5RaN0xd8oX6MwYRMri09CutGFHavWUMZXc8jXnmiV
G6QxN/Tq8vtc+EGXb59vY4557u94Rs7yp/88Z72LnOuVLOUkhQzIHksem/DMxYuR
fI3DXR6zFhFGUozPMm7uvKUntMXmpwIHkwQnYqHDcpDnlojzio8QNcoLBprpronN
Ki1BtB6G1VIqRCmj6h6h0fNgny2ZNcUUzsuI+/bPepb/dbPOiOW2HqScNNZrKdGN
sw8mQbpq8wEcbILVZ0WLa1CbOAcyU91hnMQHL9xbZXGq9hAdJ0dQhOjromtw0lRD
rCytk+bVmMDN14IQ6CjY4x2rb/v+a+/beGDDkObNZUrISwMODhzWzKlUzaMcb+LX
6q9xIoPqQMyf3d5iP+PIfF8GdpqESCGbYhaMtNRwZMqKNDTOfBCQIDNMzh+b6+li
15v3DefAPa/0tUJk+eesQkCTqUWs5gAh4ElTKW5WYXLXcTGMPWfClE9MbA8lF0Rq
RDWotSUKynIChX9qZbeExta0efp3yQbUFItAikqT1C4qASE4iYu5bN9+6makaPu/
+9ZcwVkHbPCdLuq+Wf6ZiZgEqN9W/SvdicXd2jwOuuqWlEDVah9GeWoEgBxShugq
AmpOY8eDCVB6/LDyOh6WVQc1IVw+sBcTm8eAj6eoGF6+9m/wpBuyBRhX924SqDbt
Dy3tzbWDXhJLoaRDowQdvK4GMy8/s05qnBhOVZA8X31AXI0yp6qQC5l3QOQ3KzCJ
59QwIcgzubxUde7copC972PBxs8g/hmWIbetJ4rOCPFFdgU3Di//O8OGxTwrwetL
fWGAhknG1JW4IhDjM8WEHL4cOsgzIzNGEjKf3b2eMp1uKjIOwNFrh2ytpeP6OFxZ
+gv9GSiV/dY7G2lJdxvDBogOM8bLqVPwAUUK9dz2Bx/TwIfCwAHHnxaOkpZst26c
cJyUYZzqLF+ikGyDAjk9WQsb49MC1JSzveWwokUrZhpPC3zmPBlIAPKzuF9fhUES
vihOrf30ROoAXhlwk4uIJ8VjSqa9BhyZGqACfSXjG0JOo0rFm8nvqYjXO8NNe+x/
qWxDH4H11m7ICflYs4lL4eLo9ghFCj5Sn9pM1Tgf9XcPc7XBiU508WjN+HWKBcNi
9grAJmp7lIMuA3+SGiMcQObdSV+KBhO+5R5cu7zjJBKED4KDt+kxM5ChFgV+iaRy
J48Ne/nnHizP+/N/r3XmkNMhCdKXOTMF9Tfh8KCBNMgi7ugHV0tsfPG4GpqszVqK
sZKzrJqPmujxHnFL8SRtXhCPqwEijsl0OFUFuLJ929O186a0CwruSOOt5RXnbFpe
8UHTiFN2cMXVupAePwjiWP/NSUOkUYbTjANMY9nsfdXdkye+J1BlDwsjt25vAQZ9
bt0PKkcdEgM3IHb6NIsk2Qc4iqKA16C5ZWGZsF8TImCYlEaTfQDat0kRfHy3m0GS
7qW35NdikPQUGYIgM80tvCPUSJLq4bQY7752Rn2SK+Kd1Fq4VR4OOVYkYjl6RKNY
ZpFKDKC8wvgthmw6P7Q//NmcyoYhSjcyCcfGSPCeG7ztmIb+X1jvRpzAPqsY/uNz
im1nMhqAaDBQRJ0bu7cl07vDbjGh9YoFk3g508t7ytq9INJGx7ZNO+dcLcw+JSMU
e02UnUIyx7q5UkQX+ULishn79hkh5U0uvp8ZbF4Slon5NqRjLcu+p3yHEYSY04yB
czSFdA5zRaI1cLpCmrExyI2kqDDtlRbVdpgRTyFopXbtzpQDB9tQCpUuJND+v2rI
B06Adfn86R8tb388VTci06jbSwkbjrQFL8TkHV/d5y8QTZm5+OBfOmrkrrqf2wu6
r/nLPG5gtwAjD33otEYhIZY5DRXESmYmYAfv2fPzqHqIIMCWqUaFsKGfctI+KGRE
/LMWEGN5kqvGgp74MKfaG10djYl38zmStOSb1Oqlf9RABU6Fa1WuSkhYvVVmGm8f
rbIQAijQBCR4VLdOOk47JGrn/Z+xzbbYqbGdGazwpG4pN46ltjEFx5cELlZ+oo7o
n7hlYEvL96JSEXuNhATZjk4Hy2Mk3J2FXad7Z7fM05gv0qWGIARXFSzm+zHMM1l5
KHUGS2i7IHr+ioWMMprkm1Vr5P8z4/YuaxzwzunxMSDK2DAWKzzk9xBsv08lMAkm
IJTWJEkhRWzjykJJWgTmiI6CYuhUXrxiOrwr80Fx8xPDxtVkdOwM55Yfr6Ce5PwX
jg1IPRs92A/eYw62I75WWVLfuPKROoRCMIWdG9K5ErD+77g47+1YEMdYTEmo3mv/
F0Kz37x/ojovkR1WlFxyXWwii+Df2Ff+43jKFvKOwTSNRUSV2rZ0406iMUKzIF1W
/sLyZvx+9c71MIZVRpdDGGukjS48bCMp5MEngE/OHD4wXt9iyO49PY0GfawjQZy3
G7dB+grMMz3suERO/7nWEdX9k+7yptCJxARZcuuxJf+BId6wXtrhooiYP4LZq8D9
d4suogY80b1EGB2REeCDa8JpykC3k0kHFRxa/cpgEmFMemLV34DoHpstBXT20VES
NJ1ElpMzounaGdrYupP/kW7Rpl/r6/GuT6aBjaj6EjkaNzsI5G+8KoDxnPTw2nz2
100uBaLLDzIAzfNpNJ2D6WCSOorS1rZsUCHD+UM2L9kY6HpMmMLFy1ByZXMF0eUB
lCJNbRGtYmU69AM3s39u67MAnf9hRIfeh701B9fmpLRscaRPAhismSwC70NTPs0E
1mGSZBDgjm/ooLyLuKmGUVIp4nncEXNKSuW0vBlAB6cu70YWaHBcLGTYjQ4E/TQj
Dk5Y2tqgM/exwNanAerw0PY+q1TZrZojUESsCeyTcZn48Hjd0ua9giCTcbziCRzI
j2YvmqcaD2g7mNZJFRuAeV+hDYgknO9ZDQSUmtmsM4WlhO5b5+aJTKfgd9pUAbA/
e3qXDaK7+LPTlBUsq9zG2QNzxqtvG84TAwDA8QAPbq7QlBLwBUct5hWMOZAegZYf
IryidmchhBa8dLWckfgJPDBp9AVyUetMRy07N+NGdZgD4Bn7fboDD4+yHdoLJjSA
sZcaQSH5dwKkxf/Ueu4NWD7lBnvHfkMIGejs5BVhAnKHmKTugi72ZhhMRGdHgRpI
zqlAG0DP0+f6n96LDqeSsrERfvHVCrXPVvJD6j9bcv8pmNx1j2m1qRz0+vq0FScg
hgHTRbIcbGRaQ5OAvELl8UMN8AFaw+4bEg/F+XvAP5z4PplHx14q7szHR96K4Ew4
H8TKXq8/UF2UAiegEPnXetdrMJCweAadTHJqfiw6VyT+8CX6S3BpEvCTt32sT9tS
DJgO4VF2X5QdaqfreKQeGMTI7eHTKJ89/ptDIw0byw3kAFIBznrJnVpfxIpDy7ao
6IcJLlXRwRHyfpSqyMcQbWJMihO8BLDVNwoHHlKlppzi/j4TjyZIbZ9Oz7AdR3jY
79vmjfTQfEAjurPPwP8/pEmpfeYYigWCpG7N014BFq8be4JNWBGmFB/9FVtUhlsl
W79pRU//a32mrHTvhBhAvoYcvaXKYC2aZNDDU5GJtEvz29uuCvqMZtlFiB7P9MEo
n8p5iqp3uVZMD0FF1x0Yg3bHe+WJ4ZD/tKI5lW+rvAxZlpuV/J5EqsWiryLT+4GN
UwSZXtzizcuN9f5DoWQHVSNx8nWOUWxk+An/jrAKEYdxSiMR09OOY1KlpdrEjVLJ
i4jfFxNBwk9hLCWGoEgUEwQsJODFZorr8n7OqGfvXs+x2DCuBHsOtSECoIyVcBws
wvxEHGQUisos5yTCKVB47EJQu2ph2P2rBSYzVJjup6oCS5lVUkJvmXJWDLn3Gcxd
a+VybZQCp9xFGTD8KX7xJnLHitC2So8+T12Y5dMJx2xseNPZTyrHavsoiUEZC1Ol
1lg9E6MXfgP79Sm1gBkwRt/X1uHSKec09Ng68x0Rzr7zKFK/jtiRY4wBuhdbSQHv
os+eY3GOV2Bq0aJscXazpnWoS1P3rYWZC+iNk2zp6/CIgLHtG6LjvpRee9b0hlKZ
g3hg5687G/4ndtszceRgw8wDXAl3wNXdqbtB0sgao5hBCM+iga8TXcU2NkbPkiar
0qwV9hf49X9qo5mCtGLr4Ge/ekuq16VgLOU9bq1raX5zvIRD/Wz3/sSCd+DU9Irv
7P6PM3UYixCYQ4jb0EIVBXRJSEc2MZM7+70pnLjPSCHgTD4pVoXRQ5XBsoi9aCaF
kEMa3Wdqnqu+Xh10oYpd/hpiLhy86L0Z+SiJR3Bv4epPITiTsjJdUlKFJXvukdLm
Ew1hrBI8dgkXFAMyzClO6iWMobFH4x6x3RT9dI2THElt2SHVT/BXpJJwOAYVCRuC
khT/tncsyBmg8nhoehwmzpLAJiObw7s6t8wfavbWzvw9vLDyBireBS1g2/EUmScz
eY1JUFOYnCh0+CurxHGP3ZBnsEHri9YR1SyMPkils8zU+0TpoIRSj+ClhFuamXu4
B3XNGvSkJonMLbbwEiLeKwJA/211jFsF29vRapkUt2HCc7x1GRjPaxGiDOvlxwKH
qAoxDHN5Yt3TiQbje5PyjR9i4ksbIV7LvYuIneIfnphQN6Uti6hE8/H91opGtiT4
vRmcXAy0RVKpb6GkAmPY5FoQoQ0MHbr0H3bWeHP9AkB1LtqsyLvcy+FXrv4qX4MA
vcYiMMlR4sxpnbeerg2+Lr7jCWXgrvYRFFAjZdeFtd8supUihbrSV/+AFBo7w7AC
DEjWWnTgOvp53NnoVh0Vz+qpkDbLE/Tw5sULjUIY3keHzEx2qi0AYBi87VNsW9zB
sHoQE7OGQmqRE6a2DettiyOmce1CpDDMufQg45b4p6XiuUU6Art3WDFCqtDwtJ55
kdVmEIBCBOdcRMxNr3wgAIN2r5amhB7vMDVlxHeLvn7YOEsGIaDUAGPO3DxTBhZU
0hrHTQtRgbe0X2eardlCUp7axy/9QvHkodYvTL4Y6c3cugjc5PiV1MXBMNUcxP6b
L26w7x4X9NZbP/viRl5tfRNTQ7RBErJo4+X3YClfT6N+vfU6zlcHlEOFYU6D6V0P
okktIapRIE53TaNrxvJ03ggN0X0unuL9ACO9STzRcMwbQ6ZD53iT6ua6SL5dYvGx
lK0UF/4yWMp/L7SIFDInGVeXvi1y9Ozz0spO4YOOTIPjHj8mveD5d7rSWq4vkPzs
zXIdPiC3BZDSJci9nSHVAdbe/xTdEjsDVEMN0Uj2fitxeCLAUcrI5ZJeMK0BjX9O
9VbmXX+lMqub8HFkj/kn0gQDGg8gd2dq4/EGgZhCD/pPz8+qN9Se1juxd8uZL04r
ITctbkKg6un5JzO7JxJEYfpGHJKNso0GsvM36jkik0z/A4mhT3YpSqwhXA86m/5t
hRY+r1RDL2JyMxzmqle8qxXMMWE6trgNe9D+I6oYnj5Bx5V9rAa7Ba0VMSj8oolP
ZJykqyhYofV9DrmUusGWfbmjbuS+O1/z61GtUg4Vc79KB8HO9RVfOcAGsm/eoEp9
vkCZsZdjnhcrIBY4BMWFxYtaiv2EmHlTKiAkLDcLAjSo0AcIu0Xs+AUDnc4ZEW2T
GrFWjf7suek5GU6dTfCMtcsFY/Am7PUGF6tZwi4/Rf+JtVzu+HR+bplOWNXaeNes
aaztqHQR+chYCk+hBRiyGRsS4HijeBDAl/xNFcRgYBJPFKUqC08sMPjWAMIIrWxU
g/6sRwQO80lKCQxiLE90LlIo8gLnOncHH93bx7AlTNvdqvH35N3HR67Ipe3fwQS/
9COAkSU30o4AddHnMzkEDSpanEL4uGk6HyCN7SRkc2DSAi0zJMdKGjNaKzjgw19k
tZvquAbeu/UhfA7swkzBCWW7TYh7TYvPEdQCAR+VX+4TTwaxDVBMxdZ7mYN7QSkt
tu9lmFyfBt8OG4voPPXxPHKhfVD0RC/+9PoYKTd0ultgzlUXiDfh2PtukY5wdK//
/9/5/IJNg/Cm4d+aSsLR7MALSw/ydfdt6sXpd53i4AiXGNV9I4uDBfT95juarZzc
fjAOW/U+6+1FL79UVt0p9tzbA2LiArhn/mYDbCO7LgTQqpI6hPvNPmLGXco7+lHF
AaRD9qOUjKGEsRfsQjNaJJd39KinRy0IvhMTqQbbFWe6yl53IkbxwmAyWH1N44kb
bihKztFSykQ5GOJrySe4nmxV0nnxL5aS3MJ5oywbETc/lsHDmv1De0MS46Fu7UDJ
gmrFj3SaDHd1mCNMaX0CVfSwjvQFABAi3U+zZR2VAn42zuAXiYOs21PwuQY/oYlx
dkar3g3TAFxCP5FaDVF77MkNi4Frjwl3y5tIhM7RgfNBLJOnCc+WckYSuT60Vp7g
14Fm/dAsbYjB+Cn+cZaosQ8oEc/xdTX96vSsvQocjBofNjm6h8KKqOJn/ik6kDJI
Cpdi5GFlidcK6lnqaOGnRxebcFODh8CNZoZ35rXfcHdP1xbAcxMGt9mXLi+Nt/Va
0LBYRtITXMvM/k5kFEMDHJZBPl+j/Ha36ZafOAEyGMYLxLNcdBYHyByuE/8opf0J
AC2Q33nDVy8e6hVuHqqGLEkgVXJtTmuqp0bBB0eBxTLP8ClVyolxyJ9P7DqtjJvz
nizfrQYDSEPhW8tOTmM+WC4JugDDPkWhCSaTwSuL4IsPqwfBzJ4k11EwoU7lP0q1
v2DeYTNHoTjwpgsBu6VS2NYymFkKC0hYehYAOGapKC0Q9ED3Dg1uxc4tzIK/J0oH
sjydw4GhXEnqqriC+SaKIDG/pPuyQMz4BqPol4+bXKTUUrtCrmwtv/BbJp+Y390F
8XdFWRsHGn4Xfm5nminCNTJOoa3Wv0DLuNLTuwcC5KMMlKIjemtlEdOCMGP6/VM/
PH97uB3ArJXbZIVcU9kjvTTqtAIMD8VwbXg1BDGKERoc/urda1cd2QrWInMdOUB6
1byqj1Vc5l55bsAbYIzXtJPaCl8o83RyWzktfJ30hcaGJCUh4aRBgpe6iupSsd7O
gBB+pHkjpjEjlLZSlrbexCfR6H9QBm/USucHUnOUuxmOu13Nkgh+62zUpBpDcVLV
tCFeTCHT6xbZEaKX2rwXhJeALHrxQ/P0LFk/UZwaJ/7qgikVgx0cgzgD8R3TGSU3
oRzeFXEtfSFJAfXzNRe3kKBhbtO+VThpBN7PQh1sldo5S0gXQ5elPhr8d+dY+hK3
9VbUmy1y0FwFL4ZbMQlCl3+sAMVJ1z+63tvTkb7uwfqfo7tV6XBzQ++iZXqM9Ftw
Rggg5bx1bpHRUoMztTE22yEASwzhoa2SKJKV3MHoSy98nXR14i4ewXWla1ULJiN0
u1xjjhzr4FU2k28K8V81wQnjjzofokARDyU3ozffaNGlp6eN14okMjDmZKCZmh0B
cd9vOd8xFIUkYhVJ+n9YyMsLeI61QFwsQ2uZcZLO1pAXce0VURtiq9KP3VDeyO5F
FJBmpHT/umZU21e1KhNiQtEWx+53Cjg2Y+kvSVz205+2uuEjEBIonbuZXLdEi9+t
k5wOUdkEgOpvkS+xdyaI7IAJD13tUtX4fS28LRnZKaPTxDHni/ZVC1HvbIsKcR2N
yRARH9Gf+mcw5IdFzhZlUy4FwoOy0zDQwebYx/n8btqL372+vf2MYCH6NmKxkGdU
1eVfcrFLK4mYXaQVMF4+kb3s4bx19Bf9FPP0PAGIxXbiQPn80gc/lIE0JZT4xEl3
i7xhqoE+un+fPRGIXfOt8O8Z6revxwSMVUv3cA+/gYlI0uxtnNmbIQNW6VDFe52c
yy/Yxg5ro7tiKviuTG5IRXYy+38xd4etAmDLOfD7x8UPb5k6d4prGRJ8RwqJLJyj
yFr1i5PZUyEQn1jlOlXrEJEdrhVU+OFf90iTCgZMSwFsJvHt3Z4h1JBk6frlYsq+
eUEB9pLwkauSyoPMu2VJOUIlcrXZKRv9UkUsDBXB8buBU/Q1tRa4Pvs1EufkDXH8
HufsvqNSKs5MqvA9vEkJViYUZk8HiKBr+jU+IAujnyaOlDhdIIF6IDK2U10eXDx0
+ELE5hZkvCIkN2+pKPVQZNmI6x0OFRyLZMvHDaSs7AJ3dBB1zi7COwXaRhezRA/e
lqr75o6edtpSFxIWzmLRO7BGlJuIo3muWnHRBTFXQ23My6GEHjV+qfbY8gRajOHM
supq80wK+/SXSxx5ExzESRDEfoEr5ubrZJEjrZ8Oc5WOIa/ikBW5VIyKyTqhfnQY
ydAi/JfYaKGnKtEYFxVn8ZmRl27w+OrChNjMJTHWarbe1UABux4hiLlaNQJe5p6d
NetC5PwPkNIvuPF1CYYpn+GvzBIL+5FlwJavLWXZH1zdblVyECLx17WypgUtLCdP
7G5GfBIY4zx/wMQ0J0pfZpShGvlLvnRRWGpTqV4tQQxtcCE+Crd82eCoA9ELcqEg
kcOFd5VEhKMEd0TzhhCa1Nv2f2DGBxcVM7iKtQZK4sFHhQuHBQCJmEneD/IaWu6f
m1NyQzr/nd4WN01+QpXnBvJSHJVh0yL04yFKzljFok7ow8Nwgd292luySl6nNFEV
S5xPzl0ouTLVtscVVnO8Ezr9Cj6/GzUreDI04sOjVRNnJwWnMKTQjwvGXex4Z2J1
B4DyFBpxLm2sHC+a8E14vgZHyt20Xfg2d30/E1DMvTTp/0uE6kQD7CsnR9VWuQ91
lbe1NPsMpNcTusUX2UKvgYr1FnoR+OmJCAIegrMXJW3C6mNCy5SyGdb4xWziQtxv
JuqXcQ/e9fNQKOm2kgZWqWZqdZnGFPyEdIOdMmBlNJF3DM8lOyWHFt63g3B8mNVi
wBpsOV5Ko6IPx9qNxFjVmQAxgoAIdZ94oCrRHgp41xWklFyEx159mL5h99iFzwr1
DQW6xAzigAYdimJ5xZxcjvOLKixNu6b9o/MWafX7X2Ii4iM8l85kre7ce6STTUvk
33urZneAvaZjDXcbyLJ94SE4KXvYp6JE+xz+arzLepHRaIUmqEvUglpez02vBb0x
Ijb3UuIVH1Pv1WF0pw/QkCVA9U/tx/j0MZmhG1PL8kMwBNrIzCoxMBTna894KmaO
Yw1J2QhmVwOVH6WROOItV7S2lmjRjD9+i+Eoq2GdDhHFQwSex4J7kOxQOo6anEq6
sRfdoQy3Bqhd6i2Jwlqh38JGh+Zj9NMfNFgnSfN9rxcOKOVn2HULOcKoU4YGy6Ob
dQFXUPlmkhH50uoMJGC7p+c778YvCiWX3FMTRLhPot/XJHFUCRJXSNyrB9MSjD3U
hvGdZGWyExRuZJ+hnT0lQS5KGKjR4M5WIXYyN8Z6A0RJDAssS9Wp57IUt0eJldeP
NB3uSDMRUNGwXPy6YH0gruQM5L0KWy/uC5zvnY6kvscEJfzHNLutJckk1K0WHpE/
XWAjr8hTw9qKM0FNbwG3QPGXZPVX2zdrGb70piZOTbdfUjbAARxe19yFErrtYyke
P5w11jj5XGD5XOD9AmP5iRYE9xt6VOT+uQ6NARCGnEATu5kIaQf2OEk/0Bes9jFa
yzE9CuOXpX1zxb7Z1pQFRd24MLyla9lHtUeq7hP/4BP+HccOAbk9XQw+oBe9hXZV
yNtsKYZAtk9qTXcEH5wWlK1mvJzQ3H0s20SAjIOPRIGq0pHiT/Sy2TA4IFn7vYdM
ALAVXOWP+wGm+2fTM+m3TUp2lgfZNpw0m5efgmZ691GMe2g9bKGIf2SmbxD2SKb5
E7u01uYSl2kSfu+pILb6MkKJoMlTPMIxQSsSoXKHCZZyOxrnZqhrP0JhE/gfdCMI
HEzn9ndhAZYQzP8xbGY02YPXOeT4uMe7ftpdFq5wvKTxnVsRQI/Y0AjWlTHrgO8G
du/WBVSwc2KGaJOty25aQvBFAOmP97QJRmCqHfx+g4kX5h+SCbk1Gbc2n2tK+/Pe
4osvCdfk2yePUk8ecgPSUO0ONYaIBekuJESlfOJ8P1tRH0ne76Gsl2zYju/7QQG/
axCy47FKYmxTaj9jxUU6Trg+LgrykCBce152ZCLzhe98V2v2y3zmnwkyjzHkGsWB
40x8bD2c5E0iZvTJU9mgxlDv3csPq6KqVO95OqRcronrhLft2L3VD7ZlTErng153
sMLJMu/IihBUyB7THxb4K0Yx/AFbUSM6ZL+kvIAOIg2MOipf8+lUgYSLin+7zOwF
ubLBsslmrIJNKIXyW6N14bptaSnVDoPmVFyPieD+YtVTvWOUazZmPpRfcSNVBLF+
yuOMZuA1Mo5pzIpyfr/5sKhxqtgYjnuj5vsOt4HDTkxEvHAp10pCeumc2OJ5yZER
ZBL699Wcu4ldU2rKIKz0vKZEpKAzvlNf/pthZ0lB06fJZNeR7byXeCRJW3fIHR0o
NRdN8PUhAI6Y5jDyihcAG8LRQB+rz5BQIYKs4VFhq/tvdV0su26b61xj9KV7LcIL
zpL2AjbYm58Zml4I9bublpYoMBvmTAlHkPeaqeLGK/qKKWqXrCXfvJB4VzEDIPJs
V7ja6bAjQRRowHOyJBmAqcm2mHD6DLcDrIvDoKwRFyPXz1+zigVO9H0mCRGvP+MF
hLomltqXdEWs73OmtohBIJZgmZ6Y2fszhY37/2sStyH8J6fcCTL/5qYpDWbywNVQ
rS9HBIWMNfOaV1ogXCYVIZrbjpUyb9YeOVI9DpEaT6ZA0PZYOSdIVjHSaCnxfeTC
nZlNBzZYfKUtzR7ZLFJlctRVFAXfErbSitgT+Bz/T7G6pbpmv1h5HxI8nskPrgqE
VQqFnLgOEwjdH6J+l/Cmj+uDGMDiG/ryKLZCT2xjWQq02Ps9zNu93mpzeDcsvupi
gEV+YRDfBogg7FByX9LQFMTMlKjof8KJkcZSiWnSUPZRjcXk4JTkLRKX/3fl0Quc
kcsj70MmtA2nOZ4B1YXXZ6PoCdUuEKPiFF3C6e4SdeqcOwNMAgLg2uu8w343uGkI
LiET4sB/dsXuuZZBzQGuzae0oL2Tk9WIOED8QThDGYvQBRvqbed1E6dN5VYcGSRX
s8kzumaVfcD/V2mQQlGGDBOY2r88EvHnwQCVMjspW58SNiTBZ6yMwLGuVFMmUM1e
gJlo4OJyFneCwXDtgpZNhEApuOESNpjisoeYwTS7kkAomW7HwAL/ryk2N8gPvUbw
a3e1edynnK8clWyqjboCYJM00yuyZVZr+touCgqMHkuml3d3fn75zLh8uhcPDCZH
Yjez9n6kBtEgI+qdtR5QR+Alt7YR6ihrd5DLGSQawvLbEeIDvprtjNGhb++SaHTe
kkCJl89XZVo/vtoz/y0yOzeDAgAdbpzmpKRwDnmuYbdT7oG31g5ZcDkp2lAUGAaq
chEPRr/vPFZDjV946PHDuWkjvktepehXgGeqgqGRnpqF0WAiz4YM75ChJHl0iveX
gurWr3afofPc2Qa/5IAzkXGJiLztsBBpzso+RZQy9asv376RsnpsgxmDBAPfV6TZ
nXaNJ03hoZ3nwnNCoIWPI+CBfIihQ5WCouCfywrTgXLpyHjWXtAmKZ/rB/HYPh68
i6cUJym6CLenOOuPvTDMlThntbko6LJdt+v0l83kHJp/eSbSqVZOqygFgmsLupiH
OG00A/A7n/PmEaV61tl12Val93mO3oHJ3W7SpvWrDxuLPtgc1YhTm8UeNt9W09Aw
pa+EpjjnolOHc4deRmTJ+N8QIPPoOm8oAOmF8gCGDYrjwHOVFREaYXiEb95WSEDT
2+xVnXokbSwws7UFmd2hq2KpUXK4U/7MZBwk/BOwIUt0gKxjjKWBfKhuW8664I0F
rpSMO0S4lGgwRSNdKeR8wpQuednLP8FmGIGD4VMZwCGbkLCrRRtpIGZ1Ow3q+e/E
tDXJaI443Q+95OvnhoIMaWUkhaxRHBbR9cQeqnizcyvIfkdPCap5ze7LIM7Pi3cG
ac658CE/3dg0j1USEAHCz9CxXLCwiSxi42ZoLrdBZQyLAA9epQ1NY2Y71nw6MYTn
PdTXRorIYBZsSNMHkjiulGaqjD/ET9BMB2cyJdDmCEVG2wtHLN1mGpTCbFvZ4wRy
xjQwg4mm1HEdRpaLyShOJCZlWDX5sqW3sbxrOslKy4DT4iYbIV8zroXLVobEdJWD
Kk/lqrNDa9/qXcZSVIV5I6M4iLkmRgLrH7SwO9sf1+MMKIJ5VIpvRJLDqh7AAXMF
saYLTYxIfR6Tt1tcYbnkm20z44hyZTV8P+dwdZZZ5JKZ0Ks4s7+ArlE/RdjKUkmF
FRKbKrh++YeTF2yZLqyuHquFvSUWUhGFa6TYj+vKJsjkmOdpcACRArXOa5l7Cn1r
uYGA9+tbx6DF9Lhjslx0dBaQVm+y0FhR1WrhPuE1BsVhroLcQenhJ6yjVPNsFfdj
O453n971BwfEPDwHIoPVB0SMKUk8lPOnzwpTovhSWzgK65GO2lAXcAeQWRDtmE/n
lh2f2CFxosme7T2ngLjMaYzlSStVCcv3AXmXNMVRciun2wSRPpIvxACoNzUXVOn6
/xDVEwcPUNVRVFRgCCUXV1h9xa4lKaMQfjI9qqDe0FgSbxp8Pwdv3ffFouMIgJcL
nUCyOb6y5GlQ8ho2EVN0m3zdzLKoMu0ckoRnGcjNt4McBXXs2r93ZbLAYj5CSIY8
pxxRWyhQNR9/Mkyoe6VGn5H2vCwsHyDbxadqzORD9SdjswfNhswJ8JWqw3tDHcfR
m2J83boDwljSKuJPfR4yeLjx2u0BgcYNx/Qkh4eJS8H72ZKigICi7lrxLv9HEqAA
gBUWmS+jrjeJ1c8N8BNfIPZyLvGI4/mxTDLk392q0upuKlcFes0O/JLgLgOutYq0
LGWC3+7itdW3cah7xA/jhNiAybqeM9lrLggS5vDoynB9i7SDEA8WwrVJZ2d4sEWt
BH0uARnCCjdpVBUzUfCo2XaXByxONK47mNItwQFEI6jinxAIsDC1K03aKlhcjmHY
kMNGvA2y/lW/B1emSs3GAMU8it0oBoJ/goaUd/Pjefsuhy423sprBvoIOQBTmO84
DUb9MyQlW61kFfTh9BgyO/MPZ7lFnhfrydRgZfzWN/oJXC4eyAHZ85e64iWnqDpY
lg0vSqniYt+OciiNl6Gh3QjstHrW9msmgwi+OWo3lOziTO559vTHeHolrMOkVvop
P1C5N/Dc+k3GDm8Ru2PIln64vkg9frFaMqZwlM/3Hat0/1CoXWEP9qjT3Z2Jxrd3
6h68TG2B6KgcQNbzg5UxCRO7+oaZ8V3Oxy1PnP4pbku9v/4wEIy5ZZncTa6xI3O6
tc1b01ho/R0YHqpLvFEv9L/rx/swvLraAOVH4fuD7seYCz/R/vDCQpQUcA3kRMxp
7C9iGG/n1bekbiylExykVfod55HxB5V0qr+5e6kWBkqBEzsAg2YbPjH2KBXYLd2U
I/ldV9CCuYeZ6vNPZnE7ey5ve+sbNxqk2SDbRuNGMUMbkxKFiSYoEwkKm7LLHXO2
4MAEVjJspa9vkl5CeTv9JA6QP3RPLclaCcWr1fzQ8R27iet0/KR+XP+p5voaOkGY
32kvq0hWwxac/f0TEAKpdi+AivV1csfN5Y/M324J6/uZ06cMuKgWOVNfOCb5+r3u
vz2hfSZCEy0lDdDHOpr3abrCK5/y4/WKvn3m6ZsNgQYLwfRePQRm10nx5j99zg3w
IlD+aeTIZr2cc+LEMTcBpwNFtA66WyHH05iTV5kp5iUAPepqMOFcg/PRUNMgdW41
4OwlXvN8D/6OSVJG3MlpFWvDPH1y3k04lF2TOn8taUtP+gGhKuVnJzibHOfxzV30
2rp7rULRvJuKwfioevBSVeIvoH7+naZgnLb5ODebYwV/hedgNoA+EuL/eXlZYgLY
ORKuug9SWEOgIcj7ng9fLVD8XQJSq8ymcGPcNSTwMVrDKhkGz4mLjglHnDWtVcRb
+TgzaW4c+Eg6OmheqpGVvJXV4Xf+xdQxTMP8Y2X8OLspi0b0+7Ki4cYo6X7dstBq
8yrvf7H50oVVkVfQqh6Noce83beBziuWxgrsTHrNl1UmHw2ivcXKWJ/oFHt1kMOH
EB6TfOkuwdCllNHZ91y4Qqeoq199ga/zMFunkGcIcyHBCFRqwMBqpxOHyijXQJp7
uOqztwQrfXozV4tdTDyAJmtnLyG/MKVNvYhySIGHOBeuuKD589EyS7tiQc8LN9Hs
v6pFPiI2acYMFZ7LwKVKfTa2N3kVX41c7liXqk7qKE191yGaVPn5zDt2vo+ZzwYO
TvpqDbNRCjC6W6itIyXIcScZdTBM9KB4qZSDvyyDGAxDqCCQsly2ss7XFyx4pj2a
8Lm9nUmjb96kXNrjLrkGQw31EOM3SQ9ofUrErz3Hjn+39bCgGpRLHAb7aQcDz4Yi
gXA4mN18XEWXSuITk5Z92K/9pokRGNYiBKsd5hzJdcPCQs0QUHxYmplxfWNyXjDN
l6iWtrmvQhsIjYfmrZlB7n/AWcWQD2UwiwooFqUkV6DTuzrN3p6FbAFkLvzSb/EH
ix5n7b4T2WXo5BpIV1/SNWDavJ9dYyRtBhLUW9MzaHYptfHqlb404WhYAd5IMXIs
pFrmmpjz3Dm8t1jEn4bBDxit4O3CR7RENIHULPgQGl5eTxSzuReciQHd6PLyQJrD
Y8v/1+Onj0ARQNNtx2snR2A+oILYMP51J4avAJtFeHvUJhrFiyzvc0z/+IlHpQPS
9gAMVDnOl4b1RAARpuLdeIBToZNqHXpCgxPxFprbohEkv0KaqmI9wj/vWKSIIOsg
Z4f6fxkAlMLl7zCu0cpiusFkDCSIJaQJJfzDj0pTlpMzIPqK7wdzwGGLWMrPPMza
5edyBG7ZhR5FFUmgxWSnKD4xDsCzgiGeRYx6j3d+BPVsHUKkJ7bdahHG4kBFrb0g
Ywk23utR6cJRoWjmyyNfR1sHfR8IAk6O8FUFOGSU7VI2q5PKt6ysY6yDw8KxmQpN
QlvVAXE0k0jmzGG8UM1O5tW/gmsOO1qEk9UVb1W5pfBqR5HZY98FQyxa/E436wmW
IFzmCdxY0Lc5DFWxZI+FE391M176Lv8MuPTzvwFchYKX3ycN/rklM6H45RP9aAuh
QNwsr+loS69IAwDTasRDacGRqLGEplSMZdiKPs+JI06tKyq7Z7eYhDrbKctoj6st
rbfDi43sd8otvA1UxN/akb0N0v2CCUQJdG+DWNq1HmlZvaMlN8+aeACaTc/RqnOc
yk3g9GYZQDmnE+RApwYHM3WAfB1dVVtn9HybrCC4etoE/DZYP2EZCSsCQ1gZnWAz
bvAobsQeIhRbD7Uq5IDre7KvM1GpaDPFs8opPbEoYIeIo3bgi/b70q2FHhxl2Rur
5hJmYkV2T2H5eWglfjN5tGvggMkBEfHb5cXgE9dTY7R7y6MUhhiS/j5rrexKtpE3
rVLwnIq0VYqt1Tsf0WtVqF27ozn5DujI2zrUVmqj0j2tpByjyEB7atKtCVvG9iQM
7VyRW7rb7FhPScwPtS64k5Vg5RJPmwu41E/gJmT+JYaJcg+/3TCUeZxHUKEfV1gP
CPY6lwxyCYlpMe7oJUTe0mmky76BFbfe4NVhFp0AG7RNtsUwACm1yohXStr1lyBu
26onmmlfabp3zdO5ISnfxiy7KeawjGCo1bSCye1nEXYD21ZFvNKs/8hAQ3rk8vVr
RzoQHJyGhIPHnze7sYKpKI/wheLbaa0qrGFH6/LkKJaMSrYzw6V7RbbOMXj0rGkv
ZZKMAuOgNbXBktxz+jHK5utfyOUzw2hzs/wOVxvxzLm6ub0/4UUdTRDa4QkqfH93
07ujuQHM8Uq7Y6E4mkGbRazH9k3uHQCssMbu/96WAVjaLaKoxV4AF0HIZj7/KXlt
UhDWUkE/FSD+yTqDBbfLTczjfjFCUCoqUeejelB3Bh48Qg0u7jtuIhiptHPaOeZ+
J2+5PV3ZCA1TSZ6GwDb1tW+KrwhBJF+O/ENMNoI6n+1Ukxe/x5k20yAgpVQnWcM+
OYXMRil/Jdvt1C44vWrH4Ab/ANkJokj5M6VChAtzbnIQFjacMvzYJHeTUY97bvOc
puPvTHn5WBO8jrAkUuvLX9/myVk5pzi0OyLvfgoDd0bMIRXkeyqvKa8q+IwKMaYS
r6/DTC00aAH6wCo4TLwpdcj5RPEdoKNlibM9DG02qSogSFezqECwRkK9MjtWCNvY
uwo3qSQ79RLPNX+y/Zx59nqgh0lMObjWxzI57MTRwexU3e0GQUQPwuRrOSI56p0B
27ZbvXCrWpkG70yTn8IsQIEWKAomvTvCJV4XuE+c6eLIPIHY983WmK44QBVoIhO2
ngkxCYBMFCT0qdWlYp+ZQuxYLJtesYliRkW7nX738RECNwxcsCjZVRvXqlZcB72t
ysYxkYqR5U7hXfF3Pj3L+gTZbriGT2Csccsobbzo6/3R3PSY9qtqjnFybUjEJ7BV
V7wLm3AKM5IK1aCk04znHAlPkOdS15jn0cRevzyHA1HCdHDXOkjVKYyMfn3RDuRa
uL97bHrwapMxn7Lz81dlwUCR34vZh+Dt+dEP/6/sQZ3HXYrp77NCyXw/xDQ1HjBy
xXbyc8zcctrpICma/oVIIst02zeBficU+sQh8NqNwx2myyhvoDuwerGwnhbQiPAZ
8QYEzHKJTITJ3zS9VAoTdERZZTAJKeV2lLGHVVhyJCeWbyivAK88DDY5QwAusREH
7ZgP2Jdb6Hj01JsrpsINgQwwKFKmZ8GDdAniXSU0N32sTofRLfUcGuDIMq534QFw
R4o1etvh+W4ERNnEFqhOc6gtV5U3Apjtt7Vo20cAta7IAwOjNKvL21Ew0lK6ytjR
EpGA5crLPEkXNENZywjZvuO6bREvMV1fOfNAhlt1v2ATiK9EYzfMwde0VI/u8492
bP0Jv2xNt1CfCtb2pQV9Xx+g4MCu6mxO8XqXzIMqnRWnhzScg5zPXotmN3JXFnHR
YOrI2yOEGUC6hz324J6XqxV7a7hn3Q+goCTXKvXrbh4eAQ0Z1K7ck5mNJPtcmk+W
kv6KRdAqQWfdj4FF2mZCPyVZomeRz+gjYIZqKK0xyRuVhb2Pxc7C9s80NisdTXw2
8mtnHndM/vMeTN1vBebDab2L2i107ZsGI3OIDmVzDNcVkRFKJeRSdkMbYrJltqIo
Lsi9kPzwtuuraWqSAbitITuBYAEjlXkbyj2GjgBPr1RHNY15igbxaptZXFZnR5vK
jWxoYqJBOrCW4CAE0B3d0gUtzMOx/yW1RJ0CF5Q91i3G1McZc/9Q3/nv606fYxve
u+IZamYISAm1y9akjxxw6+8behGQq42UZ7DNh3X3Nf3y5vPtxzSgalFvIE7AneCP
/FIoRDT7nVI4PDijQRpEy/90MQWvqhgpwnzoNUi6iZyszTxYa02dYbIz+fyTSDi4
Dnc70NkQygLddL5dz0tzrH8SO2wvFd+bCZDYReUWVIrkkbYjKTQthBLcZqp7prnB
A1Rbi3KJn4AODB5AZBsU5umzYzyvUJN6HrBxbfocu5wg7R38bHcbvmAljYVdXk2L
JxEOoda/REKpC8c9AQ6gCND3rAkt5DMzoxRwllgdw+rCwJ9VK+5d/zlkb/y8d88P
p8C2iIZyNS7qzOgWHxw0W/9WbuqUn3MAVcvQtTf+Tckwh5uBqUSvu+SVMzIQ0b2A
YpAenNaXNg3ahDE5KyRcWIouZrVV/2wLIcUY7pacyFBURxFO3pEUTLc1km15EpZr
hgvpYX4fruKZpcEbhYwlGstpvmULe6tSOZm8oKPnkxV3zBfgz1GqKF1iP+RFV5Kr
qoQNmW+aNGlJjiPYZL6P/8y1gTqekWKaumzY0+R9jdHkPpfDMYvcWb4EnRwWusGC
Mge+IVU5u005ATCNRgdDnYAYlSEGi8m1efgfpMhFQald9OEqIsWxDERw9S/4Y9HU
Ql0ie8b7rjRwlwhd/hgYdnQRMVk5AOqa76iSfNQUPsJrejsfGBI1+xb9js9d8r8q
pQC5++WH1DwclJTlo0pR2su4sXLUlTFWXAsWGNZT5+lLsps5gdsug56EknUvKQVT
hPAqsvK4B/GMpNawL0wPvlqFzaPHgoZRBc/se+QkvWDV40Th8yLSSFx2ue1Pkv1S
jegHTl2Ms70rQNYHmeb8G6uXCv6PnXiiSy3j/0/oV+8yxGKO+Gc1RI9zdd6Osdhr
i+4aewQbbbTwQtvTECGyn1uovlkovKWZ561Ks2QUSS29tonf7p796XXFX1Z4yac1
tA0yTfATDQvAAxrpZJ6vHeAQrhtwcQXXtidcG5OWvq/rwcnBYM7dYI+MNosEGMsM
VF2g3zu9O+Y/JM9bZyJmaCuaUdq/iFnkEvNmUsCZtCVnIftKkKbT8ob9AbfSAHw6
fz62FCyNkX16Op8U1BdMS35ZsperOXSpcSb2pwMzKX8b2mbOCUCfjsaSCLo/iv0D
DhNvrNnSrO9jdZSGRVKtwO3KjgpJ57NDoz6KGy+DB1J+lyVeMw4XzWgPDNHnTHhS
NsS3mSA4cJdk0FTD8A2ZK+9iiwbtQGBsKaJfFILX+1rulIVxdQMCLeFr0y10Ytel
Zhoe75eVHWbZ1bB1+sur2CKLSPggi2zyeoeecpjqRMFsvoKnOUeGR9Jimmvy14IW
dCr3scubv7HRDkjYrLA32Nb90S3z6smTC5+2bGjH2cM+nxMIb6/3CSb1ht+OsQMp
5HoayIGzwtFFgU7Uao2Zrc8xZGSp3CMJxKzJbn9T0EyngHBZzwRgRD5JzuEDoHdq
XOeGneWK0D3RWJMqMdiVhsV3jL7+iuw33d6hcXasnXYULcHIaraB2UoLXhIMb/LR
rpXkp223Cp6/9PjkDYu+5bK5vbFVlT3gjQTJTPIph4LNwiCyVqX5Utk9kX04+ai7
oiS1CS0BSMk49MmFJQsPwlercyc7WN9Ob/3qEF0axUtI5uBWaydfrTj0mTAk5ZfE
0v2LiA5Xg5qM8eALf1DhkRQLWHpd3/80E75vookOeJ3/U53olpgVEuaSrYyzBfgW
OAQC4cBQxt6KICmJKOtKo4yReV3EEKHD8ft08HqRPn3qcWvhKrVHMPYVil6Nmt5J
8qHNfNkvXD+0ROptzwjJy7EaY9ZwPDDAtQd6G8t6pUsb0WeCtEKedcFKW9I5E0s4
UC7GmfZTts9o4RX8wQURg8M0hfjT20Ntkn75tCVBmefft3v/6nBOE0RZHucwXcS2
R5mZNnyrEooIwWUf2mXcpCyxLvScgAgF8XjcDOakN6UAeRzyZrGJNgtpXRgYPQk+
ChjrDwetTjwdtzZn/lqcsq1RQtlP0dxpZC08+2xpkDidHvdM6i/VtRusg9sP07Lv
a0C1VRTrHwUWvSN0U4dDFs4wNlv6pCNyc/2LSdBJamJrMQTvxL0281KLO9JCNJ9n
ryDkdvcDFC3cRYTdY0TgKHX2mMul20JRpLjOcx3+eaJGKYg0y7dBBc6fxotT6Gqu
njvkBakvLqHlQfAwrbmOPHXfBcSWS2ppf7zIkGfB+9ViUxBOyPQYQ+bVMIrj80pc
lDyWhUSo32c6CCrjcwPhtn8CnI7T986CAS3MYn/yxRXzIP5zq450kz6U3b3eArNv
kkQpbTXzuo/mdOo7U/b6kHln5cEv/LFks6bSHFj/3+iuzKAWJESvMegdg8cjbJv1
WA45A0jOhoRRq5LUFCa2s3JLeMRfKKbEsp3slX8xaO842JoptTY9l0i9KAK5DKny
/8HPKQTPXYUdhAd4fjJDuBfm+rnDT8xzgD2bNzoRm+/b43bREwosz094ZV6FTI0q
TGzbe/53v+1Nk4RWMM0N07Ef89F2tECEBypOAMip6n3LzITVtBvohwx4M9K4W9bf
MVi/VjDv8pivhtFa57POZc64xynIth4aeH4ZtQiHuq+8YcopG4gyn74iAglzpsrJ
xGNrCACG8hJzZO3ktR05IjevD31eVt3ib3FFOj5jLTPTO7DUeBEaKck2wQXg8PZU
vyxuk5MFOE1nsYm0Vgg0pjEKOWeb2RttNyh4EWk5YkMmfxfMNGbQNpelo4lhJQTl
5jFlO4CgKbEvthXCr2cPBk6C3YusBAH/PLGxaDgtahYWeAVGm1JO1+4uw2Kjbrgn
rJHDB03/RQXNC8hjxh2/aEWBadwe3cs6cRTrfjzyRRYO58lVxeIwVjg7wrKcckZU
ULpSqe7dlag9wUq1wKtGqd28VrPKr0MlpV6qLx5ycVPRcY8rCg9DQRXWgNDCnb7S
YklfkgwFI2kmHxQQa35BuArCaPwaYCxo4Jc+IC5Pwxd8452DftjYh7BXN0guLcJr
ocVq/FzV3g4zy0RmMvYAR912Aic9qVZWuUNJ73S3i9CUcfewpteTb54GIDtBXwxj
7BZZrqoRJLKoLK05WXEa/ax5nt/vXQQ8Xt4wb+qpqlERxLS16xp5YCuds/dpJf64
EN4US3gJFL2EP10HaYhecqG0ba28k3CjRwfgG+QVMuWoFUiFKjcVxwOJAoWGX037
muXFXwNd4But25vuTk3z9AXVSJZTYqzgqCONHcgqIvhF8Ms3jt48R7P8b1F9644i
95nIwXv9851TOVNlwjavbh57a1eBsI5cok5K8FOqhPckExwWuaSVoo4JRJdbrqvC
CWJ+JPOfn0AQGLEM5Wd0O/Y/AEKsnlyWgbo7iR5RfpjlfUexonHImLvhchAesN8K
08bNEjTRofGloV2R1l2//8Xpuei2Qk106bn1ctqKCn+CM5ZPsmJWeiGEJFKU+ax8
mqzxVkk0Bm7fING0d07dY8PbW7fJ5y3+IzBdpCmtcbejGzKyrfSGl3P1tqwt+rQ/
5P6VOx41aUhT594YCOhgCLftZmHMXYIVpiGnnl4ZxW91xxBdb8FWn0/9c55NXwd9
Ho0RcU/6TQCynLVDxpCPdeNYxJreYbCS87xt3lMsGlch6HzqdBm8u39zdsQU/mae
hAmWBgEFoxPJTy3PVXMAv3yBwJ6YJURpv3p+VbaiyIyWzA9KkbC/3UIOk54WrLEr
4hoL0jmsM0t/PY0eI0uZBSJr2OFBXDViytHk0d9x0kqszEavyBf4MLJdE8Gle16F
oXXWyFGyVHvot+2X/iF0032fqhlZtku8V82R62bIrlUL33++xYNb3C6GbMhQHWqr
WQ5Sr57992NGwM9VOa9/W6MbMxEI067sWkThskmBs9XguMXfqx3vwoVopYmWRydo
dDAXnykwk+KdFhHsjHfO8MDpOnaxC3pgrK1grKMtZTHDiKYA6xxX20Wd9dlfsa85
GZlXk6Y91tKpQWuOUNL+1VLJbRQCffvjo9nw6/cKxsljsjFcX6l53eiBuOkSbKLh
u/fEOIWrgzSzmwSgMflWhtHThXdEYWtpjJwrQFw3p7Z3u4Kgb1s21Yo2zEhS4rGl
pUsanpQVljn3KXb35J8RRO+it0kKJxMllPkovxCnpwLtb/OPECwTfJfUZRKuj+bq
+Q42sUH/CLj0pr91gypAQduE+7gzgYHa64xBI9aGRZswH3UfYkfx8BNCURehza2Q
ted8/B4U38e0AZr6AudwIq9aKaVOqD8l6/nczgmMtAwE/f14yCOFU9dldSVIAhF3
YfU+mgo6xp3WjmWsHFf4bbTXj7moYvJ3iytlujVTNP4XCdeJtt2LCdYLxgt4p+b0
se28I2tbzkWkg65JvGK3mKdvK1A4Igb3Lk1tQnOLJ3FR8tXwRk4MdPTm/RTfvUSL
Z5nDxOLJMuTG9eJ+PwEfmGRme8e8GOzQWVZxg1BZzdbNd9dtKqVyi5/j5S/6mKS4
lVbPDfxVkKwNi/q4CSW8jA8GhjW/nfB1rB4Egjpyu99G7ts5zIlNoDfWkjkyd6S/
HSSqpuQIsXALzPcngqD8lCIO1YnzXXz0Dk7fkJCx3/2M9xrvLScfxOk1perVy9ve
7ExTFqezdJpd1IrZ6Ygpg6qAowrYaAzPOC3jVMkIeBdEp3FN2n/qB/kf05us9Vn6
WP8w6xqdJcaQGPkwY1o5HoM/9FXbBV2KwiTmf7cvssOkSY1nKoictr8KxrDjtLrs
XFXJVtv3Us2xyzFZZasZ2722AKWmIr4UQPWe+CtONd/WTOXLSQ6w12VSca1mywQ4
0AICcUZXNMnSxsvXhCsUS8Ue0B6qfBN/IXHBitbyS5TNVRztbO1cAP+F5WVw2MsJ
h8LiYmxWxGF7y5wNB8fADLuseXD89Ra23hjbFrAbPv/x9zM0Z2EPTfdrLckqA1Q+
RwPmdEDWYSKmSBA48Y96kPJnuPyT4HdDXv1xDLv0D6Ulp49ddLzb+Ay1saV7Wf7/
tA41uODEsHHJ5keQ3CffU+Szr4gNt32cQcLG2ZhJQvbHsPTh2Zp//lJeYccKA1a+
fIH/a+0PEGJ/OqEYUJHCpnfXJs5VeWCT12X6O+Kou8puAzueUP5HbcGkyFPAQV5Q
xk2SfVHnJtJFDnESl9BUBZezUR4S2iEtraR2JKkCeipomG6Dx/+R8rs8j5Jj/91Q
tzmr57O71szpWXyFl3S7pGQPA4DuEafF0/kbsJ7UaHu2A+g45cXorkkX4LaWUNrr
7BrpeBPPvq5UTqOhjw6X6UWEnFBBgv+DcVdTLAQ7tqEiASL7C6U2/HdNs3n2ViZ+
/USLBnnjNtWnphNfkB56DOZmpoNPrSUGhJpoIaUp/vCvS0TklScGcbdTPFNDX69X
y8OB+sesrq58uCBxSs9Cf4I5ZjnIK9rtGYtXbQk3arTbYpF1pQP29wcF1Hqdy2tM
sm/+c+9GTiYkLk5kZDTm/GS14zgtzgjsAQQDAae3syihM5fffhZ3h8xyVXhc0arY
keFl79ev/7Q1G8PCaPYo013GFJEff8qoGIUVlD3r9COWZ/0Lx4DvTJzp/llOeN2n
ceDVdDNJqTdw+4lxKX3S9XPvqv6NkuuJcegi5t3LUPAxVJP5yajrR1hXH0vvFNcG
oY23eA3A+opdZJo174DPiXH19nO8Silr37mE6xJl8ZwTL3FrC6NgY+BOhOpnDqko
JUWv9E5d31kegsC4A1j3NJB+bDm4ScsUKT1gLDMwjpI+RFPM4/rH0Ajel8O3RIdw
m7vB+ssEe83DTADxDsuDR8wV3Wfxp0Esku79IkW+Dw6hcFWjGeOUaQn4CcNRZgbM
alJZSuiTU+IV7OxJro7IOk6oK/Alt9dLEw/i3PWlPUO9fjFkE2DOmUVCP5Tg3bGC
cPYimLoYDN/FByF1z1GwVa+T0ln9F1VfGv60AEGEACPswGfziK+HN6juxINEwVqX
HKkiHdpGHOb3UrjZL0fjFX8M3h19XxUqn2zuN61RlvtBbxA6ftwUgyZpCsjDyAXE
zmCC2ekeo12XvAKwoDEWp7zD61VJ8f2unmizLY3DtvpDTImLBSaMdnlO102cK7rU
6GTb0YMBWC1L17cHaPB53+Semt8EdXh84EuU7KKdmpbIUqWom65cBMWHw36ZH5r6
KG46kgwvggIy+P2ed7CdSS+4dRSHK9I1OxKMaEtRAADO9aXbPt+kg6VuY0MZkwhv
X03KuGbJFcz0sfYGzSxg9/ufp/fsKvwD2QHf+vqkCcXxcTcz4VSWypO/NoLS6bs1
ctykeE83Osp3PN5fWfWfFtL9ci4NCBw+Z4XGQbeIt8GMwpXy3b8do9NmIlGl8gEQ
BpSKUeHXiiJCwguvS6VuLUSUbQp0IwdMmKP5ZWgVhxolNQM9fpLkdFEeGjgO3OKF
1rPXPDN3GcyWcYv2uImiVJF/2qkOILq/sHcmLTMNTHps5IXTHBEu/kBi+vX7i8Ee
+fdjxE2DHF0SssLDR+ZeS60rSqT1LH17CSkxJs1A4Y2K8cuFsBVcOKYPOsf2B6j7
wEFdL8dvhDKGuYvSt/mkoEsyRCe/1UhrN/cabYr9k9UUwZIySkEBRjio4A25pRO2
QbhGbEnLrEfb6fvT6pHsMkzPcH97hb54wlXzy2HjW8p/y+v09nuKSJpnh/FfHPUJ
nULzQaVMGhQVVaUfRKdbZB2Mr0W7WP0uG7iGhcBoiEVBuLvwJCPqmeye+1L9xEH/
c850PRTdstf0uoOUBr0KA3zdqJTtP5FFo4l2CTYSRjgI3Xzt+cflJxdWxUL0kn6m
+XYxDqvcZ8ESctJRLTi1LWFNrnQAZk98zagIlfM3vWIFNgO3YvaTJ7/euNkkHQmD
1HCmspju+uO+7ePwtnywdoIfHUFdQnemug100X8fK8JalmJkxc3YcUd13UA2iV24
V4MhBMLHf/UHxt4sumwH6OopR23CYeGUzTGTwmbAGGZpAG91V2ue49FzBSLAMMEH
XTfMH+5hLXVT0wxuxdtrcLxGoQYvbXXqS5ZwVSdxenRyzDBhFeXhxqWbWjdpc9fe
ZBHz7YyxxuJmQs+ZdIBhd5hDAmw3ThHeV6gk+sSoVn8BbMAp7g54kUoZ+7WsomqI
fy4zSduRe1F7aIVBUHs8j4Lb4iV+Qi+7QrI6yyWqrR3sezRyZ7uT7TxokfUXwFdk
qoXoJ/dLhByeh6zz4UUMEvM9/YnqKwazrEcsMlbtkLDKJrIOUAMosfL6QRPKSp6m
B+ZjxBxhaou1c9Qj4hhGmFtoSxKXMBghkQiU1TwQqdlZQi8zLXrX2jBN8ilNSc0t
IXSZz7y51o0/dHKFSEzcJDcfP6gy5BLRJlxKlc/6g1Ijpf58rGcuHShGVUXMYe2P
ntzXS1YZMTuqKeR54E0nO5rKTkAHSeD31uMpEzTMD9Yp2247sadYABj/l3lJBs8u
zkTQ4ecqGCUwSx+nATjRvSQwxsSONeD1ykFgZH0REbtpMxrXgZ5Jef0RFH3GW+VH
ezl1MSruJl2JZ1PAgs4ENB0Eeblj6W/o50g5GaIikh7bfRKDokZmpvqExTJZfoVt
FGS6uBZ72TBGI+9b9JuR5XXMF+1j15fykIgb+MvBifMwe+QQKAkXGZT4a9fWq2Z+
z7EmXT8+ETSyZsVGUy0i1/+zyFHENSajY3a5UG6M5NOmZIUzpJjaNJGG1DDClNAV
BaWcyVAX9beXawVldf6USAf6EmV+YjZXTeqg+dUUWfLbYEYxNDQRql5md/+qXTFO
5PxF4S6o0qHFSb33WuApBglvis1Rz98qD4pt0loGs3IUWkSRf4kTQq5zawgrsozZ
OSoGgabulBvL06NRqTr6R9U8p1RdmDVovXP/yFCRxsUFmva3xZx80gBFviscwdXt
O4nDR0oTTZPENmQUee4FH51XC6HVUEljxxhZvxiSDtHnHiIznnRFOCX8PureIoTR
EeSf8ofhl1bncLuyWMFu2WhpFebVmfcOkxaY4KUhbJMUdFzDNwKQktAFEUCz8jbU
ZNOpbM9opk4HvDx/mPNAfZaF6/+H6JGjsR7r55KIu5AQjQn9skRxPLaZuF1JztmS
sVKU14OHm3dI7edwiZbQmwczT6VMpNMteJy5pEniVJ7OFHkWQ50rRypkNu/9LXCq
EQqlLNMu6clWWEd7vgEcR+ZsHJnlMoKv14Tq5e6BpbhdN4hioamqpUAJchgN16wX
FQ0f3iRmus9vIPPu7HxL/QDwjmNq6nImQzqUc/EQa4QGZBa9AxUQHbl8kvGmQota
ZkQYr/RFViZXm6oL+8od+QO+hvw6tYpE0REjOl7Gbb5bjvHzDRZdgU3htLy9FOnz
XpMZfGGs7mKvowYII44eOzBd8QwznOKRhscZahWU0QI23wKhsfPuNymizEaDS/JC
TYAEYJZavm+pxWetuhfu2I0Ez3lfdrhc7jS4BUfqskl52hrjBx42uIpdL4C38DS6
xAoBCI7ysPeoWLYWxPjLKUuE8PpZhy5NejiwkD0jWDd6r33yQ9Pe4mChu5/Iaa/V
Z6R6NQUU07bqlXQ6n0TQ4fFKaaAf2IcxOQDyb/uEp8D4Xj7qauhIC7i16iQ3HSok
ydLaRBrog1/oTEX4k94Dh+I2kUvkuffUsph43bKHVeVGGGVV3KxhfxqEhhVbfVos
Z7m1iMVZ6f8baWZ4LTdvuSC7/jGSbMRDWxHO/CqqZIFAkSRhnDS1DWY3WLUSflv7
86MJIWfNgeYaOI7o3cqQ0+n3S02t668EZCfA30y5btjfMdFkNiJaQVQAqW3fpwyO
IeLHXfwVF6kHvWZuK3w6h274WBuPHB+2FO1mhoHIiaUaIqpSV66ZV8yRJIz7r9gj
L516Kin00pb8ih+qYoRR//SNKpPj6VqhobmxyStuXONgdAcnC6yObdHx4GTcuics
bB4cC11pyXDn3vKsNO4aW5LDtFQuiCjLN9I0rou8y0OCR3K3tMDgQfWQ9YKZfBDg
z5MNv7BdXckdds4GgnbwA9Z1WPHKFYtXsDrF6QB59FLfcy6Cy0ZJYuGuO9f/IScm
fJmTooDtUiC4Agvyv2I6kOEYHy0hPIqYVBLNZxSvOgr/tdfHjmF6sMBWn89OU/8N
YPh/NZLTZ/AmePVqi0ueBO/O/A/eCGcAP3Tpi6FnPiARpUMtAez0VWIhwGBKVu/k
MPYS6TxaCXofw+zKvPoiV/TNK5KqAHxKGhyuCg/zHrXqEf4XERdjvuF1ZquhLf/7
1e7hknM2F2ekfUgxrtZ/QKekmt+0PEfmBXBqoT++SHxKjCotCD5dXLY6YzGmN7yc
XdIxpM7ThP4PgJ7KbAZ0CHI9uB03MEphfJ0rcVaRT6A/g8ITGL5WTmo9dKF0cd1a
+snwXMLyQMEDuiEHRNk8PiUvYuXnqXQltFyvPoyL68JG5FrtPa8Glau0rv/dXBQ1
E1DSmYcDgId4h4uDbANv/gA04KWX58HDUrp1OScov64cPoCSoTGGVPbMVJpiJkmM
36A/V4jGy/MtKfE2IgD9uaxalM68Wgt3pR7Wi9/9EUBqo/oWoqXM7icUvxaIgYjs
ip7LncolMdDvltxYcv+ZLcRxDJ7HAnzWP82Pd5XHz+rC9R5tQqDp4Tw0O0MGY1iv
vkPlI6FBPeymYhpjT4E0/K2qYLZrRC/BTftJ6xKOT7OV3n++VMhK9F/oT+Yc8nmC
NO9iFTIBr0zGSJ1r1ugBCZCQPSW0Z9OIVWEvnbIwmAzXUnLKkc0A+rDTg9jrBMly
HKdJIqPDyGWAGAtHfUtMoonKIPK8fAUIhEDoe7M2SVwxBd39Lz9vJJIiGXuiVVh4
/d1kI8JD2o567b1uzfWZzOHejQdm2UG/m6nM1sxjGaWu9TsEd20nFND3j7VnUWKU
VuQ5/b1+jvDdhqQCc/yitz/3kSFG5ObpEEMTZZn9i+aTbAvd2yNzVR2WvMdNcJuq
fjBg5GorDwUBxCWtgvalakVMHEptzy5A2nPibQvUR1sIItfRGUz5H2HFyY9yY6WM
ROfJXNdabwxL8b0hwLp8PaN8RvWWiZoC7fajCBA36FAzH+cwMhOS0X/jZGdlI46K
HmQmr71+kOggUzk10k+XZCZSc+puB8Qj050dJ15vuKtfFk/kD+Mr5iUCWV1uWG1v
3wyGU6+C1qQyCUa1XETWY5Z5SGR4ATmcQ6XQ3KhggcWty+BoLOjQ8RpMQeqcHYOW
tWiFBo2sPH99t+8nHgbt0C4KnR+lK0Ehy0+gSIiz3tdg/+Bc74kK1uqJtbfH3UcW
IMobS+VSfLFaFhUswbCsuve3jZgXkxUbQ3GtYLJ41/yn6zlpm2dgx4EoZkDDothK
rouiicOSIPAUMGPfMMnTIAAekhcZqDERWNNDPTSgcQGQN/ZKXqVfB/cbrXkP84YX
QMxZVoQEBN+UwIMQBP2vYnfC0R5SVxHZ2iwDfY/5Lw1ZIHqZCWcl3Nq5JLE7ZVLo
mNpbyHk4DhI0rQZqdGelMPyQ7B2Bvyr1p8xe3+JwqVmBoJ4rMeakjN8b1H6SK9AH
d1a+OwxumokKZ8OnsNBp5oEgVZrdG0VOCtDKSmAyfLhZWC6bUtrjQD1v9MxgH/6p
8Se/I2dDYywYpXQQ9LAuP20DGZ2vxgqjMl83dfa15EMQ4O6E81ng7WfBn6jeaAlB
vvHmPsQ/2PAMu/0i5uiJlvcLcgqvpk9wi/4UFOyjlx5rrLO3ekg5/tXa3EqPbMKG
p/e0JZL1AdE734fL4QIMxAh29A4Vc0+s9iBxOSbWB1Ca9VL8dVqlGjgYuHzZS3FN
1vljnRMMeNH5f/Qc+I/8pn41kjJpM3RS0DnyQDJx0Pw4u7xg+yRuSRfWzPz9ZOXC
pc89jpwzIyBGNJxLhkriRyHDPQC/baV0Vj5LgLACgxYMmBWNtNbDddh8CTP1QXQQ
obFI0DwEv4tyqpA4kTqN8xAJIc5hGvBCtt6UyCctPrh1XjQpQwIOmL7Gd9/Mf1Cm
YiwOt8sxdAO5KRE54wwbTpKU7afX9DfKvgAJO4bEGpb5GniajHHry99pNzjCd4zn
DBNrjhA4ldUViOgY0L77wOK6zpgCEL+uO+pt92M3nSa+J/qKjG1PU+aPIotL3nGL
0sK9y1j4irqgRSSJgdzop+5y8YgcLSZEDj/NyA8fb6Fv8hkb7P6B5AcYHTrG7g54
z43srczU2pt/1WcxUSKHGis9z1GZeiIyKjc7qz+m8qiNRk2axER/gjFHu1jlvgDr
V6289HqnH+eV0dt0pnx1eS//Wu30DrvtvvyQIoJfRi76aITB7xxH2uF11SG4HwEo
InH01mxnxz8u+YHuGT5ahthqkfd/XoSvvv7sVrbbSEf0BkZxZkN8hy4Db9hueLEz
SEtMPLwqu0AdlL8c5wiSUlXviXKrXQuoJd3Yy7o/HR6peoCnR8vlgMgEEjN63L+d
gMR5HSli0rJQsZsPX/bGOEo1t4erPhhBtH8f7C2tpKIn6zU1CJfOifzjl+XnDaya
cbY+rIpJHRoWGrQEGWWLaooVeM6IR93UEWkn1mAOve2yVJFYkO4acakJJOOBmlfA
7VTbf3y2WH/7nTqEUitSVq1TxLbNLAX+LCCW6jE9jl1yKpWz9JP7jSWuAarHrXP8
TqesUcWnkCvpLRpQOFWe6B0OGeVx0zCj7yhIp1UsFepfXj/y1jjgdwFlGH2UpN5r
+sJgyhg/ur23H804HWRaPhd5O8OALoOQmgjHD5hg27VF5/GA6V88jMdW2eEEPR62
S5DEDvJ/ShJAbMKabUinNpR7pSZ2wImuB+vLsgOZHA8NT6ExtFYxod3F2hSKpujn
8m6X7rb2TGPgPtSHyoXnWNEm8IQTdzWvV5OpfMzxXGCX8mGVQuUS1/N4hxBH1ySI
5zh2lTLb+9zcxRsySkOzAPzGxEpo3y3Mpj0qMzkpRLhpXmvoEjbIzrA4CZMfICQQ
66F/rEgDLC4d4zumHoNKiVzxrWxDhY8BPUE0BpsGM9Jac9+dscCov41Ei9ubuTgt
6mYb2Kt6JLJkjUcg/dmIY1p/dlBGGk2g/qMEvvBeH1RPwutGpVSafVTKaQojVZeg
7/SiF8KvgCIMqTU2nnfYbQgpZoCzdNHpQC2dgvLthR1jwwIDNozOW8fiQNUv3CtA
PHTHNnj9UjgeCj76EAlD1pfdcack+jwncIOgmwEkUy4S4I+WSX4Gr4WjmnnHe/8c
UVB/VNXwpZRa5X/C0dauSmhNXj4RssouRwmgPO03BiXrcJ6mV6MekR+ARm2nQ/Az
OgVMytBrwMbjoUIF3gjDOJI3D2wtaX4F9qWpJkA5mi1BsKvTA8SrvR/K0oZUtD4M
InXY/MtugPZ8D+zGF7Da2Y6uuBlbvvZ/TPBtdAiAdrsM0LAYpFuUzc8wulFeeF7c
uXgJDx83F0pVL3ypncBB7D/MUDtV/9GbFMahVZ7lrEOKO9ouTi4UI4PNKBYRFGhf
EeqQs6VI4FLwTXnXO1uAMBv2xV4phh3tsj3U24RmRVw+d6m+ZrD5dJOReLF9VRU8
Y/W13KsiNLXIqbwadbt/TOrwMk1cBUGJqdktgHbe0hawrm88IQMFptioznIKY6cy
Q1pgrKiYONx6psEuwxQMEj8mioJDbBSK80eMVzZRA6ROQNfVz1tZIZkJbzE7s5cq
qF7x6GxLLPiTm0OmiZCb7IfNWQe4rXv/5Y5gzaMIKfVK7OAJYRK/h1XAP6T9MdyL
A9hJ7CVHYcnDTmPISMhPQyA/lEY0wrDPJMhb6m74m7MJ0iBLiECo35T7afw/3iOg
BmOhpx4QlIZKKdFO+Cs2m9wtF0X/2RoZtEJDeeJLsozDDgKvxlizGsE5vSBHHXYH
v9Kyn5TUrae6qSDDPzmVuiSmz9LvBeb98rzYPAuPvTEVDn60jPdi1r+5rYZirqYd
SBi1IO/UdIrdIy6l4hZkS83R+3C4CIPYoFLRy4pMiyQ2lrtIS49+bI24WNtN1zpr
lx/wSuukmTqJZ5Dqe2PMJKwve2bY7Kdrqv8araUEWNNgDWaTl+dF077U50dohtPR
76h7t4yC6YTrqa61T36GU2gAdG/MdEfnVn/CKU95AHQ1+x4uy92HBQHgHhR7XWcA
4lC6lyBIU8H6NRZGN3/5GVQmwbYCanzu/0J+K2I5PzFASWawV31X9ZFmfi5+VlbS
hrk4fdOfFlOIfQ8ogA3E0vb9RZufF+1S9P5LJ/N8H068RVSAkn00Ya1BDnSBuwHd
wVNCdNQIhPajVgUSTF7KczBZ6yV7ZuN56AUeALuO52YIxGVIcVRYwjmGZpOXVMVW
DTsWcCt5S58tgNXpxUR7VbIdy98MamGeoLDoCe3cxOrJ5u2UIauTk0zmIN0zbH2J
SKcr2Pl96i2qO0O9DX8IpcCTmHV8SiS0ekV6yTMQ3IYaFwUiceZn/x3uI7kNPD6T
zQu/WJndlpP+yubwCIFbH5BJrJmVRhj1ubDVnhAKVyZKzhhb8Cd8n8VSVohxDIJU
ECDRYqSxNYEyvfDG3mN6+Tm3xLq+3/YuqLVCZhg1+OKKVJ1AWpy5sy8LcufaW/tG
kGzjc1+UCMzMXZPoEE4BVYUsR2giX3WtzwtFx7hwH+f/2v9MSHSHTr29cXdZhn8T
AZ50jV7FL2hB/oB5PlV5XgMljD/mxuZDW2G5/ll6MAGYgoC2bgXvzkbm9hwc6S7N
qGJhOAaR7MimQ8m1N0h6exjbD96nBd8jD0GElyKW8M+CJ7xVQg8yl66QZkufDYEC
qcONgKrhYq0yKVG8hhLNdjE2QNUd0nO1IfUM14NKsofIsb0mY/bOenrcCTYNgfA/
Of2sghHf+Bvh1S/NWxeZADQ91HZJWBXmUObCSCc+mCH3SrzqjiXOFrY0+XXfYItl
Ryt7tFZaT0SAzrXAPCZNPq15JMO5SIuPTJPXmhyJu8ojoSYrlepJGRRBlAGwRNNH
Vc6Si6gZUI/whib+NjANo7H3bBmQg5+q8YWt8SMiZs1wyLquxBuy3uGDLzyA7Pkm
oDpK9kK1C7llMOHjoykOHE/C5VAKFG591ojkAjjMguwc4KJXiUlcMu6HDZwKIifn
8UBuKTLoY2SAhR9NYUc8XGW4U2qgi6I3klAivUkHEvnGMj3fpITiIQB+/lOtszy5
wfAXPVROdPBPpPWxlD7QdAAMKDzEimpZ1wHIEEvntQeKBA7+FEHcN+qaIM5EvJUx
Dywb3K/ufZWnCr49W0+yQGm/CmAHzeYsqKZSKRXHz2/i0zmSKjkyaz7Z1qbDVSzf
hw5+rGmvlW6Oxtng2QmQxn70uRReIGf5svijXtIDRKSYnJafvJIKaDH9X+PFeZim
6QmPpg+EdUWsrZ5VVmNJWwD+hlJdRe38IKY3AXtuOqI2BrsC/U5ShloeEVczlMSD
8SB9+7QFG7+RFhXZR2HddPYWP570884d4FhlECL03zv9MDitsNPkYjcaKXKyMDiO
wxzss58/85HBOpHjT55g2tlGtV1JTkt0q4PKmYqn2pdLa31E+UJSsOkrra78qZ5c
DjGQW118MCvLDcn2ciXFqjDpvCgyH66Rwg6DR1EmjsUGfZe+wHEA/UKM1Djj/+uj
dooBzLgHng/4YTH+nuwdWML/i7DAXzTfALIjMedpdw71JEUn3NXiBgDARZiVVQYq
pNrkkRGenh890DVSt9GSerzRcTWNlVfoaG8MaGdKNqbYOzJ2cmUd1a3ExyyksGgj
LvgPYO4Ut2Jw08YLsj/Ki/yRejDQeoqQF4xVqosVBhd0o3D14f98wpruYLd0y20K
RIJlKv93K7sYkW7XUHAWN2Um1/A4+UGfQdaY9Cd8fZs40lv+BRJLL83sy+XyUoxT
DRkgTdSHJ4d+mHhHypHsgWS3QL5UAafE8S/yqM0v6wca9Nl5u2/At5cNPv/Eyfh0
I3uDSjWF/NFyGptMw5XCzige0YDbsEwJyaz3jdg0oSjIYTrxHTE9yzRNg8mYu+Os
a9jlc0q3+VTvwynpRi4isrxPspVZlvG+4djHBgZFyfy5d8su/2bYbs3ea4vkgY/a
eszzK3ny/LjpSOiDF7ogR69D5RZe21J7B/wu02ugxp9Rc9KvSC7X+YCOCp+/0DdU
VqyrWpGsI9YTmdvu9oXtnmDE4IvAjPz7FTVb55dziPawO885qDiyfV7ZXdMZ8nwk
NXmJh7t5A3DEW0hNQOaPl4EG3sxbE3Tvs3ZRD5ntKHnqDPO1y1SBMaR/6eS2ozme
4s9p2UbxCWwOSSqZHaZhdbc9xgcZfyvMhBPUp4/uq4gQAvu6z8yEVsba9rN+Hwmz
+JVAK9feDM3GDYoZ4S/HthN2axumEitmhKRQ/lR26jKOEm6emqTyX4vwKbVKvpih
LE02LSOZXU8g3g0DJLwVJYQdPiYhnmWksjqhX+oYcUduOii0GbnPCG/CYC1A3wfJ
sL8WWp1Oc3TUOUOxScrNh3fAp/zuWJO4qC+HjwZ/IOGDBG1fpoc3RcoGjpAtldya
QdBemnx8i8AS1wuLClYqSiHegUjOMzxXHa6a5x2y32grX+aoQr16rWWkopImVSG4
Omxo5qgAJwm2c5zu3XD+gax0u5/pzudqvOJXiIQUl98p4WymqoHBQocAN039ynlH
npAgi4pAV7UPHJLKibiLhX56Z53pdXVfWTGvXhfCKFvqqkjly44WLy9Ylz3wxbOj
C6z4Y8BqkzXEmMG6BEm0HJj4F3UR50v9KBIM95Q1H7rOKIqwNLvLo9JeHmnIVwOT
wqFZbXInkXYS1n+MmwxjXgO2rcBjU9zlPzIOU6Sqs+t3RJR2Q6SAoqWQmDiiVatk
WPaXjFPhHQiW8AMn2e24ZMI58WxzruYFfyzsyps2cjCUbdUu5UfAKCN1KP6zz+Fo
KzQTVAZ58ObeKX2u/hkXcPX6RYBhefaw/Pp5gnhcTuKry46eTznNpMNXhjaSdayN
P5PSsTRdtknMjZAh3IB6EBcKa2yUT1zR2MyyWnoZgMDeMCUFDQl1VRjNYK/bTiMB
GZwy1g/nop9gUB8CMF6Ff7dj6hVH78YNyV4btrgR/tGlCW7I57EnLuwede3vBRY3
Y5TdJhiQLfS5xLJUu8r4qC7PuW1fq7mO8XDmrTZkvf3hbuPNnw3IkAX7GzSDqUl7
Japv9A0YfhybMLIg58/reikorErwiYslaXlqFDzsVtqhWaNktCm1sAijGnEU6hA5
SIhGC1UcIXy8eTwBBJyWIcLnz6YcFOrYEy1g6Yn032NIa/O336hl9t7ACxPih6s+
eE7sltZR4PHc+u+QWMCB6aInYt0o3+eb1rT5KVjbPfZceP9p8VyMwp2rxzslqoi5
ImgvDHrZVOgoPkh+D/NaZHJCYRx3oftfIaqGRfaWbOiaXHw3qnYtSS14XmUPgOF1
d0lPpoOSTrAjgewydBdpFhmTpAzaYXDPINEp+xf1LlluaZ5XBcUfiS619OzSj1Lw
MihDeYxB3JjBoD9IOylIYMguhcjUB3+nZ9uMkl1DjNhEVj1Vn5fsM64Dpkb3urGC
3H8T7ofOzdpE8aCI+3F43WIp7uFE+sd4gwlX3QAnzMteX8sl0R3dZ9ktgQ1/IyTd
gf/TnceT/kAwLMdNQ4ukx015HVQfke0cQMlObRyXpqfFa9kqK7o01gjkKl6yzQSM
6c8ZZZZQ/V+75vM1FvB8Ueb4mlOBcuLlMgZeQlo+74lBn9oVlQbyeAlCK6AmXYcd
tVSKWg3pT8DjOnWslkuYRZh9laVsDBFCQvTI/T3Ve8OlJFrBt7hmhTPZbaC/QgeR
CDyc5cWXerSLZXaN1gKweELgUImqFjM8wKsLX9HY4K15DSkw3Waa+EkI01NhIBA0
oWZBPvif4Ud8c236WEkWXUYE7CVMXQ/23Ln2WAy3lhodfKXAgwBL2hpx1ci1NVqM
cMo/6AiG/ul2zY1jDYYxgSfUhO9Wi/F/ctXbHos0Gsp4AXrIhqWBE48ryo4/CcB2
4zKckFZ6JAa9dI8iBYeKBJ/EmZ+i6203o/KrFq4K2xi4wWmM8mJoZVxQIWjER7Mf
C2WKkSfXj9aJwfK/IonNmBliVHR+s7HI0G1CK+rT5GqvYNc9ENnABOwnzSH5zRXa
wn9EPUnjsxjJ5m6dMyctSNyq40tDrTJLGiWarImFUwXWPHvKCSNY/xHWLM2NkIMi
0eYBmkD9Tuem/+QSeYFINo3y6ijdc+DsOdS0Ki20l0IbOzQyec0wbofTbWU1Gdmy
gyFDkA6F4FNic9OfFdsEQlt4tKFkqk7LN6WarCW3/iRkY/+U2aKrETQIGyAPebAP
JkXo7YaM5aHQLriSrsPaZ74+S0sOAsqMyiQXUodSgdKjrZBAQprY22/+tuuqpxQ4
krLVackZW9/3woCV+RE8RrPinw7ktCzlpf6lC3Qm7Duu6Qwo+c1ieBNrWLzjoHqe
Ngct5f0SYn8U2fmuKuxh1lPJbb5H7j1F3DXS5qCGHzaVlrN6wBZi/Z4c7qj9Id0A
GumevUicV1ZwpHVJKapUvq1ziZzJudOeL4oWxMelKlQtypL2j/0KK15ItsUk8qpD
azgf2q/hRgQA6Th7xWTQcQ0vd6Be+Yy4OJp7Mn2kq01C1/7z4DRozraPyWRXgJpM
nUpAvsjQPeSewe6M/Z4R0KpChXNAaCUboo3VPm7lhbYpfzf+3q/xy66slb1rY6Jd
ZFaYXmPNlsQESlnE+KsCi+JatLq+w1bm9Zo9i1bw4rxL71DBGPsWLEo8W+H9ybdg
1eB4kYvXLJI78++AOnvsSM74NOvtzkzWjOJgZlC5hZPFJ1B3nF/l8e0ca/d9myao
DYMsa1euOvvDCbOL+no34Dt2W5PB5NHCfMi6SVJykKH16eLv5Y7jvBGMdM7SawMW
wOxcFqIdJ2UH4OBvyDwUn6iOD3C+WXWmEMo8tmd1RNDGi2ila0jSNtBhYd9bYoNy
Sb/vbM3KIUjDYS7zn/ZaAXIQayHBYL95Aun9b4J5JabhCHPClX6Pf6fqFzSQ+ibH
nyDXirBlrKLVqynE+yNp2C7cSxI7lPgYV0hB2AYk3Vco3NEJZyJWg8hAh7zwhWxI
CMakaQBJ84lgUq4tCZyq4r3ObR+n4k3Bn5jmaIuubZfE30rrKqu61D+CW/TcpOil
8AW3KgrPVNtIhaKwnVzKFGUvN3PTN9XhbZxRehWVniqXCDa0jYbWB79QIpX2ehXl
naRgx2+wGkBl4ocFB0DMMpOHPQjym3TmX1q1mv9w6QJyXMh+U1hkk1BPVY+Z2+s5
SAbRH4BVo9Q9MaoVt29IT1G7DF+bwdbHdUjAgOAH1jz217TGtJIJjmf/vJhuV+4d
r+AkcjdCeITUVyrkk9dKoqIU9iyd9qGRfSOKrNEwHv9pqNTMljRulV0xhSIBf8nR
Z91N3EtljIKEFGh8qN0AYSobCwyYYm31QHNpLDm8eOoXQGnwpiyGbo5pq4JX7QYB
8NlbdNs05vU81OWCb3k7K239PF3Ef72XZ+Dx2kx1dLN5vgyH6DgaFYwUu4DO96pO
IULTNj+hDGYDs6zktgbsX62Z8niKy1weBcvB7iph1c0pCLAoQ9VBNIJM9w/snAk+
ydyK+qX2mg3MZYWi7NT2AQ0/ZV6m0tmf+VtrX/MXvfUe6OeA3ARJDJRMG8ePKRfs
16c6f8IqMh8bknnqUfN6hOmXkj4YNaldhAA2YmeZ3hLC2b27SNnyoksF2MPua4G4
S9iWN42NFR6RsSfZorqs5A5LQ1v6Un4wWiZA/0veS7oDZ/RA8VIiYW3uNLCrlitw
1msMu3nj0NZMqVCO10NlnXv6Qnex7GYxWREOqqjAeoIuDnrRGHXT7fx0wk5VRdyl
QsdR/eyBNI4lAx8xWD84qA9gOBQxBy3s55D/j09ae5W7qipVLbOlCtskkJvib/dQ
R2xlsBhMwDv9eLcsC0o/Zz907OhicbVd2dNH1T7mSII/fFICfPiQRVyFausKcgCi
9nX5Vx3OavAkZv9wQ1zcq3gPusSoEQU8yrEq2sv6AIR0h/ny0nPTNh6hjbgYo193
QtzhnvcYW23R+m3eG3dQAIY30908Mpw19xtoSmEUYRdGE+yr3Z4Lv9SxHEbMB5yn
TRass8RDupQz0zLP/6GQr/p27Gks+1TRFsYtRl5xOhAW9gr/WBUVMMHPqU+Pw9JL
6Q77nAMdIEsSJ/QFtUx/wfwlzNUTuP4TfRJWgqtywBJ/BEgksEAOcTN1Qtc0aBkz
5ZsBPmlkkNG4eoAwOIfhbCQC9HRk/h0jUiUkROCnQhd2fHJSvSbU/VWqjyKNKX4O
A7vI3dYpPx6khT2BcAI4FOwOu1pyrd+85/sEIjh7tx8CJrDynJEexRzGTqdsqeUY
y3Nrtvsmo2NMiO3q1IxtnSnz5ARkJc2Wj/lRvDWgOUEsibcd09LdI0XP0zj8WYHb
OpuYcfSHOvQlRuUtEvQI/UfXg9Pty2my/lfRRKn2r9mEIqNpmWos7eGvHQbLw/ej
h07x+B09eewwjl9OXnPYVEPvIHr5qJCJmbh9+oUdtdWJyi20HWO8vqnqK3zr/puv
ZzCBVm2s3i7xMWnydCqMlZ1Dc2s6SsAdVESmYCa7QSJaTMUtkWb111g2z+rtEygi
p3FeKvG1rfP7f2hXtWezm8+Zys2k1gbn5pHesTPHCntjgaaLxeWuE9HWVP+v6NdN
ty60QHCah//uB7jKWALzoDZ/lxgFtC7kRKjO3WEfgGIfjo9Var0XrS6ibTg8vY/d
fuMqcv/hZJrFyLTSHOjxRNdhSOArTFx7cGjnRgo26Xb3+j6+EDawbdGrXCAEIuSY
3q87DIGxVkpUzY8gf0BVhMOQG0Ao8qrORyEkSPjZo1CxUCmLq7mq2JX3dF8Op6v6
DIXflWXBLuMlJ23YokR9ykJ2kkvQUOx3hXs5qUxVlD6ifjm7tcWjfmQG/HZAeBHo
FzEZCR+BOamFwjNR205F04jX6bqsdeYpsH8A1CneZcxTXzqKy9mFnOEzAJyEmkHJ
LEKZB5LYPRGXaK+x4217Uyzj8cl9Nc2B2Gehp1Ewj0XxHahGlu4CILWZiYoGZ/jr
WegQs+UD7fv5Cu0xUw7qX4YbzvK2voJbZT+03lOToJ9Uf4+QoCLfUdNhkQIEL8fs
YdNMW5R6jctsOj3VFTPGuaIgPyxQBUw5kBge0s99+DNnYExjvRU7jKVhzJt4BHUW
oAd06E1BTHJUoMAkR/lneWewXsRRcgTqFfTUHXwoy2/62hzVGV57Oi5vuJwZQAS3
SQmhw1XrcynNyaYZA4ZNoN8R/5atkx+7rrxc9Pnrw6lIGSt6iFqRofu1v4oQf9hc
gedvyyWf8FzKqY3NCPgQtOxo0/M1McXWhHzilRRCJekFjx+Sbns9XVWE6Rvq3geW
h9q9pGBn7Q0mqKs+I7ImAfPLcxJ+/QgMSp1DbdiJ+a9EO0PVM0R/wuqgWgYtCCUD
FlLY1mxsgPsFqBjbgC3CXNsrLPbfS9xV7KN+++igsTMOYYKw3WYNagTirtJBiw7u
9HA4Je26SD6a968BcPEA37cUuNLKB6TE3blmqLuHeF6n+nO7k1hosc6mAR05mCXH
YhNgxO7Yi49uIKj5T/zkdyGom8LATRwlEKKuzkHw/3QtICWTcPhdNXmnFNF3GBPR
2lTCvIXMrmPR1FjASLTzjUdqXLfJjYQ9SD/Gv7Cn6CLigNdWS275gcxHDe1WwaBs
orkn7GrYeb2L4GBgCtydPQnsj3Qbsb2np1L1TM1hxsmiUK4aqAlqpPyIjmORaBsk
c1e7/WPDbkItwYeCjhymr7OQl+Bpj9v62rzQQXpgw74en1rCO+oK9fDBroRprKRx
J8qJ+ZikVkSn8jXNZ+wWzutKhCTtJnWfBrOGOMf8a4gKlDWdEgu88q6dKV5JxU7u
7I9WHAilnZbzDlQRBihY8fDZ8Wast96aulB+H0nIbrA44ONU6qS3vMfjKiqOwz9g
01nzycZ6Rz33gL7qNQJslmn/cPeKjA70yVmfB+O/AAYiY+vOkyRM7eD3FJFsy0id
+i/0Z0FgMV+8kQZRuoUhwFIdoSjM4Rv/X+bRIGVKNvh4Ws5PVNRLFf381jOekq3g
uUothZrL5og5MgZexrz+ShzZoeuWe1uqUiVVCoaY7nUzdgRFkJFaQdA2bSDUQ/9P
Z5s/WCIQU+fsjLa+eZ2Q2f1LUJPihEW3++jSOpWBbQuZlSyw9dlD8CBe9DsINIva
/WzxKuOHbSndTvcpgF9cSHBM6bsTvqI/vjXnyOpG1mOLcSdaQaME72FuLiIC19ic
ijxqhoR8iDMYsIiBKIZls7Jb5Fg1qsldbPyXXAUqkK637gDyLI0HiD5hEIR8Yzme
1yo/XuoutkToGY3ywlg/bVnR/+/ycpbehbzJIvV/0oyi8TDjtPtv10PzUXiUsvFh
vqG2j/xVKdnujgUeWMsEdrLUc6jJ4jPVla1i1gV+UERVsPFFCZtMokk/rc58t1BV
FMfipb2G9Wl7yxHypL5WKyUXY8l0vCOf3qUpU2sUC2agquaNFwZ2FI28frbi2qkf
vN4WHtzUcI5j3uNjuB+6tiYZYWqmmbglw93dLJIkJFpM5lRKuZAlgryNK/wnHc7A
+/K65/BKNBfblfQgL4Rk5MGgP2P0DJlfGg9LT8lDD5Iwve5qawaZSyI1j018n2ab
dKd/ZBrllZC/3fMgR09UrK9QmkfpfmsRREWKjc+zRMoYcjE3cO5K76U+XkyVZv7q
UlYbnDL/V55gUsYhFzQMO2KOqbprCsB37wc1Tes/FfYVarqnPJ/ODlKCsSc1TrqI
4+CtaxC0EP6K1RjbCszvL04ys/n5CCTslQc0nZO1RUM3PXR4mWSY0b+/92NKnRX1
ND0UPL8PkLD5sI8b6p/3GB5TZAc8kOJlDXQOs+GKXRSezbfrCFTK2XqY4yrh9VDo
myqylupYpcvCQpIEARhFxL21RlpmNQfFIMj7WWBq3UE+F+pFLWklNYX3o+JiS5aQ
iKsMUvNYc4r/nVz2+G2+ErvLhRWuy1ha/8ItiLaGcJT3VgRIpxqTq1bSZD1PmTjc
L85jvvrBOLyXQDv+KjNm96BxkjVM6QPk8t/2Ub3TMtcslWyO7PRnLYMJb9b1i61I
j5dJ2v9xPj2INPqJJ9ejJznoFavboUnR5EL9KPSg71kvKMiq04hc2u89b1BD/5m5
ULt/tdHL5JhQ//E6I5vTK+KOfq7qdlitok9ns9B/N/rO2SzOOTBgoa9uRpKq/6ZJ
zTQLxASLDiTbsuQWxvRsvhaAD/U0dF4FrGectVixxciYYUU7Y0oEMHnHIgOqCkCf
4MeuegGPhNTYCo/wJ34NJwCeQQTpLPxUzgHJpA5bhyqCp8YyJENzBXHodwPsq01Q
Xp+ot2nQqvKv18IP4J2ss2r50+Qc8ECetb/JmTq3fZxlAgmHQk7ee0PXQjrWXj2X
am4L11GNZHQFc4jmAndlvpF9bb356BSJfCfn6PPYyWsnqc4jm+EpN2EcgGl1lDmB
ni4AH4R7tsXREDYZM4f+xFqRRgfgKsH7S6de4qh+IWnxw8cNNKsiaOn/p38L7v40
c3JW0Js+pQ3d4uAIX2lup4eU9tvNnsJ60XATQTeNXNBjKTJeeXYv1bbpRMg/U6jl
qqVRmDIpFqVdjIzLqb7UpIgI/lvkTI+xxu+IwkYGUVNs2PZPG1E58vwV08ZaNTEX
Dxp6o0byY36VRwLPAM8UO7h4C8/D2ka7lWXJoGtofkbswdYGOpgeBEb2hcvi9sgp
wROPxrNdTW7u30s9XL7NDqVHt55X7uUSr3iAkTa86kDDrDCPy2BCwlblf7JxzBXT
a9V8cyrTFzJuJvpvFygtPj79XLIIQzRCMYSwu5nLH+o2Jw19TxUalqN/UU8LSNtw
CY7GqrCVaFbOIqC9SWXdAbJ1+aD5ZgfKIKTYJgRx7CO/z1LokGKYEbwrTc1dJ1y4
ladPRSxlGoeHEbaIEhnS/EfgFdmlw1jFNsPePLW1Yg5Ug0OnMoZG3Ppu6hLh5KPA
UW2eYf2K5ni/akmiaWqRmOYr+LPb9f64v2qvk2lvT9r3Xv8XGMMVw9Zx/GHc/XBU
dVs337yKpoUqC+5WcEY3a/QL6s7ToSzGhF7elOZ4SkXquL860jWJ7AoexLuXMg6c
VScnDGVG0EkeSSp2m662cDgDXGMOG+5pKKBvAA8SEUWPESvJ0mwCBUal0nrAhyCO
bQOdLCnl7orI1+h7n3+WpuqNtqF8QPjSulA1vsgUW+WJc4US49Uy5id2SIUGr/IC
05n6tZ4EY9pZPZTpqlywgdwI2gu6DDTp1IBgRQcAmZnqaG333qhhUnQIyMchi8DL
PbOeH5vjiZ8AQjlaLQydTuvQewzUvRgxIVGdilF+taqTD4f34ZA97y5Sq4wPTafc
5siA413HJGx/uya8N47kXtCAZVLSw0NV1qg3poUFt5X+EoM02VkCiX1Peb+mr1+/
rkF1NeqrB44BGuA6XT+R7qXs1CCJh4K8IZ6sNFSQLl9hWylk3qoxTlUQBstNDWbS
Ou27w5cy57WCu004D+Nf6Z+poVo3q1VpFLerzfHRSdKL1WYBMqF0qF1BXfJlmOPm
lmfDStkYENbEFf1Lpqy/VpQA6Wryn61W0q+pOb+bylQ4peDpip39NN1tB0eOCGqT
jOR05xR6osyYq6+DWFo50v6ItLBWMa8raobprw43Lg2CVeYl/9TpaPRQRwXoJP7J
WFz8GXDQDqKj9T4LFVLoGe+6wt89+otQ9kjBkUiHKtwEHWaQgPMHDsDLhgqUt3NQ
e/UfZLGF4Nq9RTztoQBbvm0id/uS8x8Jkc8OgJnaJj/ccQgNY2hCsqpUlxFRrBAm
8Mje5XIsbLRorFavip7psilwZmifrm2oQc49rpkqIANNCdVlYFsrZAaQw8j/vwQ5
54kOY2loELLaKO9cUoW1ZYHsRMHglbYhaZkIuy9M6KTqo3ctuPKRU9MIROKScfs9
ARQ+YQ11qB0MZkKr0o94XAN7YvNmgBGx5cR8Fex+MJGydJCg7HPpdzEDxzBQ6uZc
hf6XbvnDJ4FYkUvrj15AC6WuHhFxuxNOLt3gTHvYLQW6k+4ASDpy2CGXFvFFPVDM
Vrsiw1C1ZUlZOUL1G3l5hIGQp7Md1xD8b+BbsRugKuGG86Ad7tUqSOk2hG39EHxr
PeuqWfJZrqk2kHl4SUyF5ZqgR8xAy6DTNX/bT5PRgEJJZ7hGSfZwQjq7jy/1Iz4Z
3+8M/xieDYJr5sKkGJRjPl8M2zr+JgKa4eD5DGcysVq7P4pT9At4Pqlgu0VyaA+G
bTjnNOx5u3bfRYd7b4By2wYA64EbhUwIIygClPBX/LOG6djQ4+4EB7DBAo0P+FtM
yirxyxJzKNHucZCV9x+LWGfGUR85PPlAnW1Ql0Z5oxpprtk9uoF1XQ+doA5e+MT1
dejE/Xp2hUYqE+MfFN7DtG6kYxWoosVXAB92aeg4zdw6HbUvEZRpLWQfE4Ve+E6H
gj/3GFXpWfJ4IxBjE3uCDgAu9mcvTeSTonWl73o0MeWPWeBPkcliCIrm0RTDtXMf
x5jJTxle0yhTAqprLE4N6FXkAcNoWiPwMJnvEMnEJ7itX2UB+6A50sOwAvg/4W3j
vT4VBm2ks9vwjaT9/W0dfm0V0SBfDcYx0cNjRFQ2yv4gBUjPjUQQUztDhbtttDSz
0v5uJ+cWnz7MD21EzMMlXF6CkntTnohhbVxUdje8evW12bWS1LYlDSZK8PvaD2ry
r+9tKSbgeb9he2QDiO3ZtREJDMs1Wb/zRT7Kwn5rpJ/5LkKTdQPDxQEcsXKjEpGC
sagJp78c8M69XPilOpQ8zCyyvGn6E5paIaIhn09Si8MFcRcQp1/THuvWfiDNHCAm
fGrtxeJnMWemzvNhT1iVJcdp63mcgP8e0F9E1JS4PNP9WvmP9LKj+RbfRvRFxcU6
En+DzL57j/7AnZGXobqeW/C9MhBuHcfxB649SLLqlzUEjXS0wfgmpZRVPtjP1d3S
irhOwwN79cmDchDBPorJUIwHFgHVoe5jK/u5sfgpCb6AAV2CCmF9u/4LooAtwtpc
PJ4EUBdoSAOgzY2A9PHEeTKPk7Rmntb1Kd4kenLMfzWXvwBrt/TPCH0jQ4n0M60x
qyQ0Tjz4gL2Kw/taoEWF1jDmQpe4ocrwKOrG4vL+nIsNZZne+iSYd7LshRWDgJVq
NlDzFP5fz+gwGhwg2MDb38/CgCFl2f/i90RiPH52ChPu3PIRIq96a0kuTOfxEeOD
f5qjITASQGs278FIOXD2Bbx8HQJfTZ5WYrDXME+pwevHVjbTGQJrzWHdZnxi0VKO
uBQJ6I7yY95+t+R6FDnUNA/pXfYPL3uW9vyw1XK2wkrfieo/chVwAEu3H0KXOCmT
BHfMtdHLmY5jBh3F4eyP1I9eAgKL6yh9/sefv1/6rQ4CRH/o6lcSv1+yqPZsZc4+
FKB5te1mfBbYMcLZzScqvuRCaH1CZ2ahm4OOW8TjABqBpiqtgc9VL+M3p7kmvoFD
aRKe1pNjAdJp+OCmMwNslXs3QXGvpkZ7a3k7e8BdWF6Xn15IKWgN6tXtlPlnl71E
4zYdyb1p6EjSAXdAvZGnQZcXUxfOMAoVpSubdZpOuHP49BLKI4UOqJ1fm/3Vl2Su
34sHC1NyUWzPWmnINzx+dy8V3Y28hLHpqRikf+UwJ4htKZd2Rkba+h5iLLHfIlic
MtZNfOINrgddoaAFKsMzgQ077gCO+qlw9DQ6fTKLs0ifj0Wce+mfVjmK7c3FE14E
xxWOeaA+v0g1illYtO3AXizZlOfKf92157yyiOB0LstawnuohjfJ6gqBs/AFuvrH
G6MX4H4SbQ5EDY1YYH8hVjJ7xS7TofM372SeqPYJHx4+ZVkmEIRD6zrQbV4TVGok
b3GXTkgmXl+IuNyo2OaP7AdCFtfg9dQrydDRPK4bDFtXiTbXDXGjliqbsdam7T2S
OBaZ4RPC6FCxD9bakzu6ItQJucBGK0qqGCU7OjEhfNFmjOUD8DnJGl0TKkp6f/yP
uBkz6v2cF4PF5oHF56pC5X9uw0eDnliEfhPofFhK7VHLzJsNLiX1bokhAj/+rTyo
x4XYD44jyUm+1gGx5uA0ycC/JTPd7kxmSYV3LyVR6xoHbh38XsPDzlt+rBvBvr5n
dQCgR5SunppFIV1IN2wO5HFImSKVsGYV3gD1zmHiRapdOlhxwCe6LwiFn9JUrrhF
rh9qoEyDrw+Rubbx3oYG2UKcKuZHk6HL0gLvvFp0dCQpYAcw4W/XpEWyef94I2Uf
DuCOFy1cY/JEyRuuyhTbxoaXbe7+oKy0loYGpckYkm//MKggAjHEkmTgDtnhPqCK
zJR6Xnw2NvtkG81ZXjisNsRP2sYs/tiLxV2soR2WTsZfFxz4Okc7KNyohLdOBj1G
26GZR+A/hK7z1lay5oBNfelGSm3DohHkLmYeGjFJFkcuhxIF9Y2UxZDpt9H2Cu4V
q5WCIQCwbLBJpbzt7APfQotec7b9xQ9USkp2TlPx9hXHyeSIV7j3zEaalIydyDZJ
eDS8QGeDHxz2PxpiE9YXKuIuUNXYkK61KHi2KbSoYvidwuRB6b1sjUroMSXgTbEx
9u8SOFOEB34zlQQilTEiJ/7+Upf4Bu4RrUalxtjy/25y/t3aWVxZ3zRHQvRsIqLY
MjMknAq7rD+DIhd4sDrf1RnL2GE9WDdaJ5X8gJDe5E6/A1AQgb7+8cO1oz7aUGd8
EVvdlCejewwV2W/1O98XQ12JLowuR+2ikYZ4AY0mWrJcNVL+1hkYWEvd8jxDpqQ+
+hUkmKmrjM9rDoDLLv7YiJi55+HwbjuqxI5U51OLkm7+Vz3Y4uY4AqUPYr0Wn3sm
2aAINLKtb9aRVz9ckeFEGgznGl3+TOX5AVy3ztbiPXDPWRN0DeZIzLYhZkXismHG
gi6h7Q3vpdNXxmjK4eQKnw6z8L6F094Addi+RdR3pwbfqptOc9kqr46ASj3IKWgO
boIbe17n5eIsbHOxk1jr1Wsyzk9mdH6+MrEBo4PHYmshl+dG//+HjQbCDGWj/a8t
AhXgXtEEhbqrPB0/oHgh3G1obmy+vCc5FGlWQhaniEUMNIyp8z8ZiI23vcNdZBgs
BG3MUfIyZzIxk0WMIhjtpuajsOlNGPfD56Hs43jeth00eii8wg++eOZDhtabFnFF
SKif+4EwRyEuO9KcxjhU/k/iujYErRUrvMcKPevwGHyz6FI/PYJ5fQljmrIQ6/bd
U/W35984hNb/rxQ0l8JL25sYNX0rYSI0DSU7G5vNeN6oofHK1sybd/hXuKz1nAyT
h/YJS0KNv2WD6DLmp+mvYwsTUZCUFXLBf9O3Cg5s/bKbVMPwqm6Da4nLtu+PJJ0P
DUpGXRwEKQsfBCoXQRo7IZU4ddpr0Af3nhnPxQNyE54uZn2bYec7nZvWmEbnYl6u
wkyOSL7xLd30IBsx28mHc5rN3gfztwMWblEayfIkubIApu7jFbiDKgJNIbivHOij
gLkrjcfqXgOumOlt5RI9vqgyQDMTQTA1G/EOFgaCfSA6oyWcOEg2e6mp087Dxr9A
+B5iDorRgi6xUEk7HRuYKzKaKrEHlAZKWgaJmAH64Hu602datCUUVV4Krit+i7s+
ZzKZx4vGV2wzxrTU/UFNOr185zZ2oRi/dn7dMhp0lUhGOd5vw0fdcBbYzd8hI1wf
IJLxBwdIujw0b/sJXVG842f1S/OI1xm5Q3MKOgapFfQJcXpz4X/ovkeOuTKBRud0
l2AqghN69U1e11/F95VgGxIl5GnvXbT8WgkYuJt4kEvccHrPSOXnSlLFCiiwZCEB
sAoj+TSvMZ5HZo81Kb7SY4o1X/AnweFdmqa7g/EDETU9I9swy0/GxkoQnOC3nmcp
A9/+BbfHo3r9K3v1tqscH2XOUImbth+BTobGaG7I7CvYXBol+JZt/cUTjQPMubiX
AnxkJKqrbUC5uMS3R9ecINQUledyL1+7Moq+m1MI51mMEUSeN9ht37Nu0RnYXjsB
MR9b03k3hKforPWHS76BDjQpz3dTVsNsvKXvKmifFWgscVzOU6sP2lFyrNbZNoU5
0EeBzKP6WEAAgOpWZbOY6hCjVFF9kjBGV2pWJoaaWs//rXgFiTz5+qGzhf8DCPUw
hMw4rj1JNkXcmMNQeoFkkh9A9t83COOpgPPXBaOQDsS1mMMNgJGNqE3zylsqr4Ui
PEyCW9hNcj4FSuBB10swOBw+V/q9z7NC4pD+ZVTWsUau2Nt2xF7VHejGTidF3Ci/
1BcOKKXXdK55SqC6kS7U0+gfDpuvoAC+8RsJnmF8UcaA5nI7V990umAFU+NLGE9V
3D4furDtuSC7dfq85Nm69AJPHDE8b1RNBigjZBBL7Jm9cM8+6KjGmLIOL4I9So52
ixOOsLFkEyG19wkPMk/Uk7SM252izCYMPlV4btevHZup7ekiX8jN8Vq1qB+wuhfM
SDxeo030OpRBN7nIFp09fReldZtXEI1+irwigM8UyIGdbwUMDWb+1NSgnknQ7Tr/
DxFDn/hTof1mlRmZnIpMaGNRq2p0erXWpTIl6ixIC22KpiJsG07ttkM3fImMjX/l
5xSXbNw5oHl5NDi3mksUfsrUKNlrKp4DRKoxjorhwebMpuLVxScRTMNnXOx2v18Q
lMMqwsz0mLmP6UA7XO6/29vvGI71SraArGJKYbwuvB/sHllf7OQ4gILvMSEgaOnz
w4dkTdwwFlPINVlEyKFAMDDDTElYVjP+kPNggKAun+vDSx8pxEZq9mKzyEN8bO3o
CwPiy70Avw3aC4vAoDZN64zM/ugODB/T9WLsxrqMckyPtTr7Tp8+GKhEKCAfrjJM
2DjTmpYJgrX4CVuLM7+IXcfLt4md3HEI5NRmG+dYKnfdf1biGyttEoSZ6tlinthY
44dfOByEo+ZCY4D8aFlTixxG1ByMAfPv/9+O49GWGvCcuHMWErBf47g6aNYscALC
X9OLpPP7a91DE6oR+ftXmMVsqvxlkmerYLeGw8Uk7YeYuCFtf3SIvqvweC46fBqv
LepeHTE3Vj4xG4dTqWdFFUZD05SeEcBKn8Cyr0lxrr/PR9fo3iVWQx4CjkJstyEs
/l5Pfi1V57lTG9/QJriGrZzMPcQgHMqfTmNu+6Xdop+c1ECdUQcM7c/i7eDEV7uy
6NFXFmaoguhNjap7KJHJ/h+9U1RErIzGOQ29xgsQ/QwBQkhALlWnmqDVn/m+E6l5
scjLPPyxyx/ZYZMyKmH43r2weus8XM8RbQFig1ctW6/TcmeFmyDmtrhC5FPLYaXu
zLiPQe7N8jm1dIh+Oetc7MNSgI0dK79NaZgtEs9LnqvGmQxjsNX6Wc/gkbhBF948
KauE3+vAUzSEevYCJVAL/THDIkUVhc0ohcE8LxZqSIu+Fr3jH/9pwx3aZUGhAGge
FlCCBxSlvuQHlUFJjJIZjtZoh0u7aWXcgaVXNw7QAcKrSBkO77Ipn86XwuW0rhbz
WpuXDrU2pgeSeGx6tjRLE8unlmWR2yynbXoKNz9eQ1K8SscQtuwFIaBZ7Gz9Om6B
zkGl55aOWEBABxdeWutNJSuzsVRYY1M1aukZIqvaAhYiCAlfYGgXXWDKqEXy8DFp
VQ1did55QqEJD/NyPLFhUvR1gMcnGxiYdDLVV+DoKdUzWdLqhjfgJ9Ab6JAW07Yp
M666oQfAMZx4FeBxpimufNi51FObskFzqYa9WJ16DcMrCmd+g+7lsLRP7/n1h27Z
az8S4JsuFrNbQaKq9uY/iL+0dDoO7x+ElRAoeiflUgS3b/MBUZe5GJykN2ZmZRIF
+uJa8IzlZo7Hz5zL8Y7VklsZLx1dD5aNwlgez3qWNxfhzj6UknEs0pcwfW/pbQJJ
ww5G0eIvEuGIiSHXET/kInK5RCuPNBQ5anRsbsCy7JiY5pV2pQADD+kXq5rXxoID
0Gf7yO/SiC3D/J6YjwwFodDMJsfEH8xuJTavO3oefulzRluWCO1CoJyMO/LleC6k
fiPferoY55GIA3vv/zg4Ymsx5tSp768sPO2rAHPfHqjYuItlerVdtItxdETjkW9V
WdSamhD7sRRmPCKvKNHoYJ/AopVsJY8u5cJe0pZvwxeX67ipVkCjj45S3LtLa+qH
CcjaJMCvjVqjyW5YT8Erqumw1zbZ3jdoKaBIP76tm+5EbxvzZB+cAMXK1k+yUVhR
4mvz+5cwIpsf1qpiK4kSDukpjDrGcr13ZmS6GiPwwx2AmBNtY4FeSweAh631F2cs
7rTOXJQNdoRJL/e112X8Wq0f7upVdrSpTsX70Rqi3wzrNVgxzSCdift7uu7hpz3j
H635f/lI6y+5P6gJ9/TJWPb09iuB8mQTIaC71hSFYnNv56Z4o/JVT26Fw+tUBOAN
jGEJKvybGLyc88mrlW90tjQKkzmNh1JpRTozKbxZR+UmeHyyO44MCQpj/MvKcy4q
ndy6saYHreVmvN4LouFIeFqpW3tqSz93z5VVWJDx+teOW9faBvK3vAou3NckqB66
7AdN3FiteonGJ5DMnVcUnSV+JL/QbFZpUSjTK6WODjKiDYlq4YbVUGZrO33PlqDm
9iK7iiFXviiuaMAgw/tsKMhTftm2h+mhB9QoOA0Kv5kFgMyaX8xuKEPG5Kizmjii
/2q/5/J6KRfwSa1RTyCfmD0AJlIYwqQAZ5WHw+9OdO6JQ2TlxgPxHCgfwwpv1P21
iE0eFyw9qSCsM2SrLKUlJe8oSs8GrjaULVQqO+qPOazhtkphU6fj9ToEyMZqGEcV
7aPAc+P3D9M2yB3QTdvEEuXohT2CscRn91sZkvcrRZZQoWFk6UouLof3S/mWIACJ
xC/TtT7S9ymc8mgEYdeMF2s+0qEYfYzS4DEtl9NbBJ2QCh5KMLDhY3PP724Jtv5V
qPWkeGc1rIowui7a0APXPWOO96NJEWBo7Dv3+MB5kh7HS+iFANYpNjDxrU2XdjYQ
ZfIEWQBUI845bl2bUEaMw7e3d5IEjY5tk9LSSaoVYECqWnMQ2+2OOyGi2JJtqF+t
IbUy9MM9+B6l6X2iD4QZx5QfPlkpzaLAXNijZYOt4tRQU1Hfj6vXyP/uiLBqduBj
XyJuDl9dW1QXEFMXHQW60Ve6BNGdvzUVk+1akcNMZwkxSfaDqBp9CLVJi85y3Ej6
zmmW3mAPQfluzTu0q/Pa5sg0HT1DElUDyDRH3Dm3ztIOWM+8708I0+9pw64PdaGG
1sDr2yf+f4lMLpL5Ig2AmtNixw6qdxMwvgiCO3tt1YwPPVI4KgoPFk/CePcvUHjp
uUdcl08RtcEDixp9JVh8oq1C4DJs6OIa9iiBfmPCZxg5ztJMOycLGS5yksKnZ4Yy
JWZD2sSIX3w6r9RKVHn7VrjbFxTr69d1jWqCUlkkQmZWZ+3H8R29+iFXuyRFGOF0
Mg2qGvLLJ5vZYhZyBFasBr/xIavA9Gho4KkBL5ek2nyXeZPI3TDskr9C3JAANVtd
Bkpf3OLJ9HfmfBZYfaHgB5tN6VSTag/4pDq9y9evY/xUygUEkXymMOTIHqLjzUNI
8uc3SND6+Jjafdhsj1pdeXbokMds2Cl2qtQj927hgv5q1hRhBGaoV5j8+8vdGSHQ
TRpwzQokj1yIMu78F2ePa2PPOy52gRtlCqTCOAtBBi20vZdoH2XSAfu2zbpQ/l9R
uG48CkGbpqdiMTdr/i9bJSdFRJinYuee92YGhwLJH5Ddc2M41IeEzmIafWRUGaU/
TMPuATrPivig440tekLJEDJlAKsnKW0GKPTJFF2WWz84mB32L4zG7Iff3O7TU/4d
USkAYFD7pYhx1E4wrqk3uVkl0nrFNPEuv7JqoGbUlxKqtk7IPxTYp/wNUReiHISS
vYHWFRV0JJchJILflchY8WjVlN1n+wRkU20BksGyq5xP0dODiVyoHk5f8NZP7H67
muaGY4n39MQZVe7Ik0QA4a7q2vgR29RY9DCzIUCsshdkuDNwdSwcZC4bF9E0g/cf
0geycCaJj+xxZKlsYrNEccp0dMgsWPoQdqX27rVrYMWA4tclUCUYvVA8+phPIFTd
0uydkBkYav4kgFVpor+onnvS26sMYnja+Qg9HWz/O5NC33Jup8IVYV0DgqXexHwR
V22X9sU+lj0kXj4rGQ/vVWuVfDJrB5WDcRy4bd88tQt+pCtuP6ADOZDhzKmEh0vz
fTqoCF3sviiTo9xbPrXrtz0j2PcYFWbzqTHZRbXhwwBgy8DRx2OkPBlJTdD8wPzK
P6KN9A+DW+GdTKu6t8a2orPBalZXY3/MMBWABdfflPapXzy5p/Krm14SIxwEDEoU
HCjlLcS0E4Eto/NFv7OU7HtpB5Qp3ZLr7seibePl3LowWHTyyP2MDFG2lIQv9L32
5Apna9TPpMGocniH5LXh9huZwjP7tdtXaIxRZJ1AG7VUeVryjl0tPnqjKoL2VWWj
v//vYPcSz+4kxOIB67eQIUFmNVeVX0BteVVCxW8v49ficF6DmQyakrKs0XTmfkNa
J8E6IbZuQKOII5cnFFfDbNsneaDfSmMF/XLtysM4OyToIvKwINC1IcO3VloXxOHq
dIaz6khcw7wfC+bebGJeneY2TBguBhXno34znt6r17K7Y9+jpQzIGw3Nme0inblW
++jqjB2Dm8e26lfMyvrlaLNqdTqpvBlEIfvUJ8uh1+bze/Qie5qBRwwttZ0NQla8
qR7ds32zMdDHERBO+eSm53yVSbVSutSaMZ06DlIb9URx3WHkPpV47L6Vrxl7Qu4F
NDEikxAjHv0vWSUkCYOUoLCzln7ISO73nrm8aAyv7Y47eVaHoHGw0onaLMRDB9tk
ASpm8PVzEVq3U1Zk2RjDu9MqFjQGS0/aiiIDfzsogFY8eVkcDJOMOIpTi1NOlWML
YZcJjiOnPS2pPQVFOvu8bJEYmU7CGoPU7sc5LW6m+/tNeBqYj621REjkIBuLJwUv
Hgi13V0adkAEe8lHx1R6lXa/l281Ch9PIuKW53qvklBDN/v2xF5HMoJ85mL9kSya
u8348fVcfgHouVQYHEm6M8JdTbdxOlRRdMl3+TisXoXOw+7DkbgA6TplT3Ke7Ne0
dN5IAGgkfkxhCOMzltYhZH8Kp7CFXx40Ac/CXZgo9UaXttw8PZ9bxfCujEmBld7N
wHqsFllqgBdcphM+2RDA3lBOdBs5m0iivmVV7Aa1k1req5f1VrxQUAUp8XJFYbYa
NRd4SrfLk4qaz5b6KccCLkIGmvtPqujSarz+L3gk8Yx4oRD1+qXuameZ6zt7Q4rO
yxfvVIYDoil/G2CK6in0FPn+Appg86QTUeNQdyq+3ae2rwSDvKMzyMgUaSu5ZVZP
ddk3E3IHXfLVlqvSYBTNqe9I4Iw37OTYaQ+q0QI/kclYwmkX36ElJGzoeezvqHpd
6PJLlrSWCvoKpjuAlhr6uXOphk+mtp2a7P53bNPiaTejaEuuj1PJ4YL86aPsiycz
dt06Adio30wHyUYEAckVNNHUgpXoly2hsFoe0V7CVlb1NVVWK/wsODShTMoxi5JI
PZw8XngjCBohJBy7NUB8K6+xDU5UftqaFzMoZatRGBPFoJYjNNkMRbigKv+Zu4mP
J/9DSEdNVfHA+O2mra5+9xlkoYC5G0xY1E2rfPcsrjuDDcXI8AGBhc7cDunCSr7N
83/mdrLq7HYopus7kwPxRBAyFgBJvOQ4SGvj+ewKptC3iXQkQlgbLGnMRHLBitoq
qqyfteTrTFwMGNy6BLL+/HqboMcdStYc6QYLcSyvw1PkA7YxYU2X+0NhGWaAdGDg
3LsDoshWuy/YY4NYeX0vvod9k3kLzoJk+uKPf9XCMGBQN02c9+C69O0whBbbfP/e
HDihZOlVsVCLUKVIqkevhR9M4zKn6UAMmc9WLMcv81T0lL3nKkHBGRwuXkSk0jKx
jYQ7wXy0th68Az/1ndBB/M8+5gC4nAmWaqHsWukDIb3htcpOm7+kkNXqpVWq5mBr
rXCgvSnjVf5tRJqHLkBbHpZdjKNPkV+c/qnZkxZDQR0oiwwC08WejRStfWn2bV2D
3GcAu62Vz/GQ0ObprpxLMg4HVQvEixdLcR4qKebX8fI1zNX45r42d9/88qVvRWMU
LtBAwl7Z2BRWVYO9AKzoLUrAk4cefZf5Y8nG6dgDoj0D1meMxi/xrxUI8sXT8jWT
x2vhBsqp2NZ6N54J4hmK5LjGN3jcW0jzizVJWa3kh2YiZ4WPPwU3GqEcYQag3+Vt
vMgEiWPYXYxRWiLiPu6273IRt48l6PUxmSPCxt3Zrnsk8rkxcxvgiiZvBbnaiU5a
vRlyChlRXb0LA3/hTLLl4ALJqxUS96NUlW1iX4PqADdjpgZ6pamOXG4OwE/Ie5Pj
Gl6zrpFSLC9Nbgx+o3+W2z9tvevAxHUKhzwOBVZosZ0UNe2KbmeNx3KJFTBudqmW
+NIl/f44vU1uSIVo5ST582jGK4szBhN3QljYdV1GJd7X5iOdH9m2rofCr0Mtd+CH
aMYKXOxKg2nPccSXR00cMvDYjUXzNMs9BifaQAqAPytjqFSQN2gBeEXt+yXj0Vyh
SFkmTwEb+KAPMcXkbiQstK8S8GsudseA7CzUqCG8c421BVTEVv5uIDVPzmcopwX2
rQfcIvXBL+5TDPpgx7AlKw0+ghgm+GOyD/F6fHb70UWHqIaTB33vlLqMnC9LTFMy
Ybr1oEJ+BGD1N7ctsTNgwh9k7qsU59bsknWjPNW0aZ2vZvQ73na/xeDGrmSEVITW
d1AafB/L0AINWOYXOCARuKvMHyHttuVbpmx5SadyaL2Ajg7Jy2LuRaknr8DE+3Tq
hcSw4LGEsBr3EzFi1NALan/oSjTDgLKRPb2ls0o6G8QzSuUalYmenP41cY+CV7ta
QttxH3SN48Lmssj755wP+endMCPmRF4u4XBr2//8ChZyywfuFpMDU+HGCWqnNb5U
roMvW2JC4oI44JXjEi+oeQiDf/LbREGKHVd47+e/5KDHfcWipo7zbfFir2nC3Lvj
p2VFjacINOKWLnvJhoQ1H4Lh9Vg21pw1fjtdbhiqxFUFdD5LspHW3swyGdYS0Bv7
9Y9LvgmY4z+i2ohxDLZNytgdyCAMyRL7nr7HR7nVQK+SeGceIEhdM0ss/Z6lTXiE
/KaxhstrwtIIIq6Xfour76+ECOQkGN8RdhxNpfTger9gAJwKfxlOPWGjQdBBQvOU
uOwq8VF8w00sSF5dhvEa2zQvXW0ZfxuTo6WyxqqPTwu/vJzDX4oXH4V9OqcTZXyk
EVyTlHf4gtZNU7DIThbmdvquL+oP0GkEp4Q1VGJiKO5J2S1xZKuMI6t3nuL+V3yn
Q/Xpo/2qznz/xNzib65Rd5H+NsyH6r9Sq5WT44A7eMuHvbpa4r6GucsiZ3DAC5KN
MF3l7DL4Xol+j7UQwJwBMftZxhC0F6gW3AE4ux7K289H0gtGtSnOy2NkLaJTYiLa
qe2hf3W0AYDH8UNZ/lD0DukQRfcZuppHlwGBhFvA0akbLiKUtZv75q9CGDOy0Gd7
XyGcIlt9tyjbMntQbC96Y+YSwCPO+tRXTdTczqf3yU0xzw0un+QRlHt3CMn1Wpq/
Ir/ryS6qk8m0vMyr+tEU420pEo0pzJO2r/EWlffjciIKanm238+wYIMAxZz4DZbG
1xDKbq1bBGyimdqhFrQ2xDwIYkphNQityC7tTJeW31acQiQhhUbTX4TD5JleBZQ1
u/RvEqOYKOsCtN6SUrnD5B1LeTrJX8SzCf0XW0kr2saWx5iWpM9Y4hDXEuxZQLpF
IGvUmtTJLNyGiugV4vAbo3SvOGtolNdTJ15TeJR7jg8tj5AorPvzrca6MM7PJJ7M
29AmdtOwhzaV3DYdQ3tWMivsmqnLJdV5AFy3o1/RZanCqDmBX72yGmn0StKVTQpn
HGQGM1SfB0KIfRlGZiV91+5nmUb0eax0VsOp/BVCWoHmeYonHb59bjP0n5jEZ4nG
fpuyJkruR4kn38soBfAxC8UApD+yw3NvLIbyt+WIBV79/YoctBGgFoLcm+Bv10AF
n9bDs9Z3/ylotPo0viNTp8AQj0HYoUxlmiDE9evVBSmoSePPSVbtgAVsv1Ncqh22
gfbLnRw7fkf5nqty3LFhauuHK7EkPvnnSnQbYHNDvMjxakz8yFtJB6l7KEJQ27k0
gnMuInutzlFE5JgXGRJkfF46AQzO97/GzrATGcDK9nyb1XyH5cW7oWfmRyugzqs+
4Z8LvPBQOYfRCrBXu9a07eFy5URbKlo4EK5DLQaiG3m4WWOds9kFt/msxiQmv2Df
zAHd1mBjHybiz8o+xzIbNe1qMb6KrLsGvqrlTe1H+luJVfjEVQGfYlDQBjGO/j1N
GJHBhkqpnJRoPG9TQsZw1pi2iWix3VVWxEIq4Nb3cFrx64ODDyP4PC7BuYe0Strb
3+0c9IdltNqx664RP+bc6/SWBvK+HY5A3llo/s7joOUuuLzp/oilQ+RiadWJj6Rj
V+tMFFqUmoen8lRmudoDYtnNBxv4v8xl5Kaihy91/51HD6Vga/XSnmoqW5NOdVmx
hhuuWtnpZ3wVDWWtxH5x0vVbf/HmLXwqKN/Ot2JlPd1SNMX+juGUYzcUPpWa2S0z
vo+QY0TXnSKEC0APbImukoLz9TyseyWRf9X1/wv2kr57AelUbFo5cqEVqAMmF2wl
JDlYapEx3T8zFNpKkX/OZzU1X5LPfZhNjCrF3Cx/yARlxR547+M3St5jxzDTtto+
oKNprbbYBubOXr0nWPApjVH1JrjCvevbHRop4hHz+PwQP6+knFfaaf3+FPz/hLlN
hbMHeH1GtmFYJJS1k28mwEZ7GbAm4SBZJLJqouE8cPaYr3YjdPTRsPgQvrM4vUlR
2A9bxhadf+zzdbwgdiOcU55zkWcpHwyhSfC64f/jEt4sHNeTb4ZeCjFl9fMizUZV
BsbMY1a3TRyKVmdzVfiRdehTSPAZB/DmEqFLrNo3B9B1Y770bZJ1TXBWG1eYvGXF
gmL+gq5JidLhUj5GjkQ0OMqRsmGE4JsHcfwdDwst2DQfC4R6Sw/LcbxO407vifkc
Ksb6kst+UjwFfwaxCxXSwp+nKNOy0ZaD10mkTx90KO/c75vUzqs9J90ddJR2QcAM
H34nAg8DJjJufg1AvGjl6FxKd/63kS8QsaefyZIVAsUp62Fq+sMOAjXqFG8QfXfM
NYvYpV0en/R0m0SnhonhJRfuPTM/vdAWZSccxrrC1IfgSzRaatvy+OvLmcRAWWG8
UPNJcb0radHQbJ88fdE/2R9NQEJ61juHPFm5GfYDVKqWVLlMgtzuJUvHIS5W05qd
YjX+46Ix+X9uB1xv63TjTJI/dumzaLoMb/HeP/P9sQuV7mrsSFGPfuzCa7ju1tH2
ggrjD3iHZf58SuCiWxaIh9Dyb8ZLwBqSnuh10B2b89VXuim7XOVPbWbYEIXgjXQ3
Zmaeh+Md4APV6ydOYrDsRe9KN0YNmRAowW5jgdwc+OkXAPdt6C9nUe+/IRql9JM/
9FD+zAWYh4gfkaUdysPK7SVm206d6gLbxMPcKTa3uI1BaV7GeLPvLmLjvpdcXSEh
lLxzu0wVlvCwsgm2manMGba0KIB9DU4xha/I/swpu6o/CvpFjP8Ru5N/mfEtEAWS
qFphhTFlBDwimFSLpIdIp8h2rFhLFLF08eB67iUwji3xTzRWnHSCJogkynb9/pir
ru99MngVpBXAOhBa0zYus3rmdyT5bU9bXBjzW+VRRXE6GQ5RFp/5QeJ4mlRWMulY
IfVWxls5PKZcMRvpMsk2CCXxrpYWlzVdHDpkpMIHADst/NJvnZOoVXkPqBhdtdF7
U2HbZeUlMMYHcVOVer6L27ZEmtPoQq4/cCCDO3xHGYdD5zbxTFwJBbmt63QxZT3m
j+Qt40uaa1opDn17w688eTT0dXe8jkZC50qNaYV1GlDUMOnzz3G3KNAyd+BXQXGt
txO64fpGylzMqhdWo5Cr5O+gZUYmqT138eVHYqRLJ3kwDlOsmQD+ZxUo0tfOLLC2
/ZhpiRMN7FSA4bKgQaoK3U9EH5ug+L5bNA4ceRd+1BheoUstp1H5tK1POfWyy9Go
xiq5WNjuZjHLp+aShAHx+B/nPszcEqFzvIlA0X6KYGsLVKvbo2S5WSpa977fJA6U
yNbVoRqUBka3s4ykaFl/QxYZmNvdJh75joxiby9PlFO5g/U7agotgNlVzAVchg3O
4bPT1lUURJU9o+xYemqdUAnQBsTITL3jqrPSIseUEI3Oesi4Y8ukV/9dfWLo1NHD
uQvWGM7SuFKDh5WkIMua4x35pDCBtBDcFGdMTCHjYb9xIiWSuDUpkHvdjC1EQk3l
Pml83L2cD64C10x3EihUQ1DQLcZd8F+YLhSKYuKXC6kFe8b6Be3JrzSS8IPusu7F
0jmKFiBVZ+rLAunhUKeYC4omKcvRMhXY6wVVpr1P5c9bt0SOV6cFgJU5jxhvmn4+
IUrvcb5MKu7VKB/5n4LHEAVZKaJEGUL9L3/ehLl/y9ZxgIeqALowuUjuwhECklUF
6mO6wy/47OoLdMHJ9kk8JKtmT9us1ihbwhOFbCmgf87MLnjm/e41vMckVDZV4xmM
+vfSwVjtVuSsbDoxpS4Zx+Fzg+BLQJ3TgWmYWp8lWAaIl7UECkhOJFuGaZdSoHqP
Aya/oUprRE4zedfzMesrHuZ3yNYiUdtsdvYlC/zWJoMWNwEzPvUw98dnQqhNA1Gt
qlj31fA/udItm2bEFz/J1ryclYDKHOw6aBMFZE0YbIEJ2T6UlH84/q+d5z6Bs8v3
Hnv63xptkzecSHK9a8UKbR2GujGBLoGA7ZVqmBa3G0i6EdtJcxClOV8BUyRyjzwt
CyilrxvsmeX++2kUlXlkzgyV4NmJ4ssiO1oiHZsuyoOuGniXKi7+H2blUCwOlBZ4
5fNjR9y+6AtQPkM0jav4Q4nPzl43q/U4lnufLq1wR/W5MrI/oa10t3q0b/yM1lDR
BSB5rCL+eCORg5QONVcmnqsAoFJtJaUeRCcyqW2+J+uT58khc55P0ruynjIVNkRw
bKG8u9ap4XgJFHl6D6k7KxlTyczxGhvmFlxUqzuURirKsFVKbYZnCsHmT1hm06u2
TuvDOc/DdSwGnRErZFDm23Ech3Cx/+tAf5jmSHXhVBNpDctOxwRbG+DLg7Hlei7v
ac7NVKb8mvIF3XXlrVjSAAdEJsm+8VQFVPWNebppqSsuu61/eHFzLkIBq2GnNAD0
FT6ElLglpSBHsXMw7c9rjm67/YJ3xWeOYpl0hqOmDyncZDIe1/M7hBh5O4iPtYen
EGOoNLwoudzytlXPaio6umuRgaZYGnKMO2wvSqPOzvRTYvrk5eMeQmYUw/peL8Ii
8YfBDMup3/0itoV84PGCfZ8VyILz14qqKqC2XL6o/pZHYUN4i/Jq9DWfyK8kAG+p
zZaNNkYfFv3o9cNP+W2LPCwxi2FH+btl8FPfjbN0hnvxZJlx3v5KNTADYV/GPmV3
hbIDHHLt5JUYopgkaBWSjwmJ9SGnWMdl59UQJh+HfWMkOSRx7rPpBlXqfVoqNQYk
lWzKRE+qTPbWitfjfCrWaLm1oICH+F8DQ75m5swfsFhwIdfiqdByKI9I++OoLf35
YwMV4HdCpN77VGImbNtLwWlhpLhaE7j27gHReQVX0w82r9M1A9EkBCwD+Siav7wt
EGeEH//BCMKA69B5sZHCj5sYVXl1RHN3Mvcqos/Ns+fLTevB4EwPenfJbDY19zMs
gMPwnnmUJ8LyQlQptZbKEWSa3dQOmdLGLWeqHW/s5o0UPOx/Y/4+JRBsZ1Xoi2j3
mnHU94vYQSU25WtgaW24kn9xXxryovfzr+b4W7tESogzXCT+iaeCbavhkE7KFMyY
x/i9h0sGDApXWcHvmPIZbh4ovg94WYrmQsvk+ZS8yIhzbuABOeg2X38+YhPpPsq9
zisUlpVS4ejewhESblS/P2SSVOPVo3VgCDBeU/sYasLqyyBROj2FV3eLcebOAUtC
CstYFC7JSG6kY7TOkkYR7lKN204nELR9Y16C7i4Xj/E77KppmA54ccucPoE/gOlh
WazViOHqfMz4OL73rvdhEyWwkVmcX28F2HgIHHWkv4XqgEuf6aTfVo42zQAgVtNO
HQ566RKZfD7OAvucgfGlJDBE4bkckG5oZrRMRjFqbMfR2SQ3rLyHZ91V6PYxQDVS
EBgtEhDe3GvsOV7J4Qks+RjWF9awJSAgAW45Nm9vQ32kNqgtnGWAZA3wlOrCjrzI
YL7BXrZcokmqgAVOMvAvzP+glGn0POIy6E48W5p6HdoSKVhsj1s6QtnOD2CyC8qe
XwEIXlJNH4UB+pPaCQBp8XfUBKDjQQXjpI8HSVmQWmtCFQbWPemSHKaWvDW1N46S
+HFtzbdtIT/HmluoS2koCOazWtL8t/WorByOUuNS5ln2suCy/gMRxEZaFeX9uLvG
43LcMeBL2PKYYjgH/afm0eOeQ5jx45GWDTdZdrZYncbPadbuIjBEWoMOmjG+Ak4A
2CYIsNy6gVAyw9KSLpDgmVe88f1kBPYv5/DpbiRObqVE/dNae+HoxVyu/D3KWxbF
Fg6CxqYV6cXxwduYLdc/5ZQ7SgxhgObRZhHqs+Vr4JtY+uJAdsV6h68iqmbKBaTI
LnEKhHC6triMb7TLH76A9uVKaplBn3trmn2h6dkP2sXVc5u5isBY6NnyT+4SuJoJ
m+PImjXRKycgjKD8Ho1UvNvIVfJAhzYKSATgTpPrg3sKkZW4qM3vCx7FkWs12Eo+
ZEPrqQJG0sOY3lqfWXpigxuuK1J54WvFs33RufDtNA/hKl0Dm2HGJat2gCVQucG8
6iDjkApYujWo1BQbsvS78xvnNJMs/z7wrvMUUF+qHA9kBbAj1CfYtXubqvqgnKq/
xBKVzugHtDvWWYci9GFh1eT+T68lyI7AndIc48d4K5WtsK0B3IiO8cBC8H7wxOqg
HBqj4mG1HtSZjs81/KcNgFZFtH15FhzaHa2PcgEedf+sPnwx0J2SAq3HpE5LYWSX
pPs+g5zPbcYO6K+b3Bl7ONnuOe/3FF3HOFd3CQMWvqYvvCaXCxNRNwgMG+COQ4Ah
+E9FZqgrQ5S+YDEb6IZQTPX5oWWmhvcMLXQlKHHypCVTh+FZ7hziCm4IKB0Kg9fi
0/KGKEa4q1wD69EoUwvnN3HVMg6QdojwnDUR24OrfM6Z/nYxFD69fdCavMr+5lFR
VCkMBW4V22H2XsGlC5BAb/hgaFaCJHeubuH0f8wolpP5hDsjPd40vAAb9vQDL0YG
h3El9GvCy6LhjFv5XnEshdLrAfgQEl4Zp5siDUUSQT++1MknQSovEdmSBewub9FA
mwr89MDHVl53ZC5u4UFnue1dLMQNBpicESgCezO0B8xjhUi7eRejIXruNXWN3Nnj
25ZAN1mnFRzDceXM7JTA6WqN8JHMxvaN7sBZ1JnJlyihw8rtRFBSXX1kEmTqbA5i
WF7tWu1YB/AE0GqlKMDQvT8ZxoMWroKeknYB/RU2VDkkL5IDT/qVXGA6uXSx0mr4
exY72TSfpNj3azx8sZaUqN+KtJ+DwCWyuIMMHnK3MKWOINZ8FMnnijUskC9FiI7u
XCQcXmPNc2Cct2eyplxjcqwsMiCms9H2/qkfxIWj88jJjxO/Du65Nx+9BVel66lo
kwL5j7p8CCsIXQ1yFiIcLk7Yf6XMZxK23kTPwGCUjuLAAM2CJDoOWrSu6tSb9Dr7
7EmR5O2Rz+yjhu8UUOWDPvREni2eHS6QkXW427fYzGThqVmopZxjKscDa4yONMJc
xHY0WwmETooBFmY3yUO2TRnNHCtqJmZ3pVXGwcfLBM8l5i1tq08+sUNYuPFKb8hy
sb2NPtbfgM8lpVKNJgmKwmHkkf1yahB9op3J6h3pMbzIDLzWHDQ8N6MeHc67KCtg
wHYAwS7jkZs/WV1B6jhD7JWRyXKcDJdY/46hrfD1dj6X8Oxo2iY79DsMesVlAVHi
+jxmOReTcO3fkHUMII004B6dukrSKdz5/qoJpShpkyHiIiWS8duwihd2uBzA3Wmn
rQ8HmAH99tQh3CWN8NCFcInW6WpUMhm4ejVLlLy+YTVpW8KmS+gA4MuVfBbi338S
fyo0hAH0EOmPASxvp7F6QwdsIlUh4/49fHHZUygD6oHO9485ztLJJW88QFkrDD0i
2axnrNuRkaBeMD3SdTbRjbCGvlERLtiMlXaaN1qCf3AxwyoYMN5bqS8WmeByIAyW
JyihFTDas8jrusd/8rDi4TLTpOdCl4Fj62oaMEuWMdk3tZ5GSlw+Pi9/mk8JYhsQ
U5ejk7vOZpxmlQaIu/1qusLvaI1luDdh003oIAwQE9BvQUtiup8QwvkPnullMilG
ms4pr9fw+dzNxCzBSjaZfTAITZFMABgjwF4eamCeXvB3BCtVnH1Lemo2ggxVOvHi
2ebw6EdK9oU2sDo3xHVaVEj8+Xcq2Gpj1y886DHo5lKe69isjTfTW01/wp6ZDB6n
ttHd/TKgSq8fRvtP96SFwtUr+RIkaJBKS3avp8p6ytbdrxE2sIBZNGB3QViAvOaZ
1VIpz+xDngaV1odeTCInHI7muuVvv1gqkXdAItdYU0EdnHOIJXdp6QVzubViD9Q0
1ZUckW6T+7PNHSIoHi6EB5I06C84miQpkG2jGiucZHD5FAozr165XnUZcKSX5XWN
Yyd2pJutAz9sDOKBYjGGCI1A9W4O8Ihzp51Ym40WTOCIltQAhuQ3vcOqKvoTKlj+
eNKViTdtb6SaeS/cYLVgoGoI/NS8a8I6z/EqOYvhkMSFbCvvkQ53ZxprPS0Ra6u0
MnPRSEcX/YNzeOjrWDuR/o6sTc0a9PTXhZ4N38hCIB4f1Gp7WPHF5Jr4Wny3t3FX
ZTYMc0nvuPOWVaCiwrUSK6WxuifFl8bxBGh8nUupDuluR86dr1UYNbxMk7CrFZoh
b6nyMKw9NZGmirg6+PNhXvcmsOXUoyq4EqESMiADu49WtHfTMf0SZwrXqMKrbkk+
1/S8wORm6VTi59nmKQszyTuiPaqCBHrNSdrGSlzSl215myBXJz3bPypTJHHjcl5/
UPFWNU1WSh3yTz00EaBjIw3w2V+F7zzmdNO/F1LuvgM4OVyfmnU/tg/iWic46/40
feMcRnct15T/xbVSz6OBupMlcKbwBKahNvm1dYAeP32/zGMw8o+gSBZ/dL7Ne5DT
d5Omi4pN1M8XzvalQlUUO1QOiDxJJ9KZ5b33zbMZ1yxpkfNeDLmLHXKvM1xvktt+
EsfuUE6G6oP5aeWeWaZ/prblM1btMpzfXY9h5tGj3BrsOTZO7TQRG5BNiNN92WpU
XPEPCTCYv6t/at90riJnDzt1RvZuRfoFtVnikSsK4VEiaXPzdFzEubMmq39Qs9+V
cto3qjKU1AvRRFMU8KNpZxb5aIOw40VZ0gJ74z0qPfsA2hIX5Cx87jmgoaWaq89o
C6XedC16i37gfoIV+SsB7y/0wUiPK0ts/GlMQiIIOwC6AJtrs+vg/U3vLcfQ0RI1
TUw6j+wZ4Mjjy49tpiJNVx0xwtdbpKpH3OAzDRKWy43o2zmTUH59GbQi0Me92khV
Oh/h/r2YkzfGnm2hGCLoXAN2Dk/9WBl1XQckyXUYdXbzIqDVAEoAN4UP7QZC7H9F
4k7eCAfWVHpNRL3DbSoJfeBx6WFN9J9nlWsFsA6ZgTrjUZ6chnAnOpnB7CnK+w8A
MRehC3K+Crp9Z0WWs7bVr5o8y1LAP/T/KOSql1IH4GRJ9XY1Ex8IivrdlF7Xx8Cv
5ZK17YEjQOoexKU2O1E6CG97DIi8ckt0tI7XDceKC6qs4nJHeaR4D3vmTDLd3rRv
sq/ynBRqPxM2J2ZjlDQO/LSlGajo0+mN5GK1iB5N4oSHUdjWKpLNpPyGqRc748ue
xGM1k7YYhg7vD2vbDEbZJSfM/SzWOguZEkk9OauO0NXL/8rNTFVzPUjvHFNclFgC
z/niDt4piesg3Kd7tbh6XUvvH7dnYIe0EtTG24gIRHPco84kSfsF1Aes7VlEQSj7
WI1+uVpc4Ho8VRSUF3DHrgnhqOlIhzWwzuWuBqBwlCgx5HwVye1HPXVlem0/JxxD
FdwVh8pSHDuYq9P/jTmhLOge1K1N2/ddFfM9QmH6fy03XbQozjRAa3Cc72//JYuX
F5AP48YuFiTwfMDYTVNUSp+hyOJQyuQcoB+LaR0Rs7btvM29f6klWbKQNEvyD+jM
Py9Z3ZfkmK7tIJkRyJA+3t4E63uR4nQkpCAcdQRRbcM90MnWH6H68hBIOAWzqTk3
3u5bmH+JOCKTZWN5MVek/ShYvDCb1/GTli/1bTx2GabhsPgnzDYy1toBOts6dRta
WG0NzrssY9O3i0BAvXShEM+9ddeKygSsEUkgDb6QjOXcOKQGf7JhZ5dtBxBPm4rO
UNZ52VYhVFHzsJpMrQ+9eRhjrnafex3tiLzVyZuzaFxfntGwFS1dn9kXNkP4Pl2B
indBfZ2FthZceMZAEgE0Y95Fzd+ucOayOU7s2eMyuatDPn9kMModlJkUxaf5Qt6/
mqMW1uLfa0VqPBoakgLvitzhz9RCFTFtLiEsf39FSxNTpmYURi2ALHRiRhwDmUcL
O5RVCnp67K3meWl7/kdM2UV+KaOYVAfH9J/DRgAvBuq01EAikJgEFzWp1PjS9ygY
DyTPL+am3KELgpc3v7qn2rrHNbxOixigUuItJgkmqYtfs+fUEC4qrgF2qCL51nbt
q8GGod7mqj/YI1I+l8TuS2/HK+ipzXPYS/WM19vwSxS83irVyWuGCb2uotLL07tB
jU1NAA2q29Hu1i6xIrbBP8ZBATFRsQKi59dBPClxyeTQEmEqIiyHkIr9YvSccQQm
RrnqRNCaKs3j0qvqQ/yRczrkXXaiRWlJMQGzGDSI/zLZK+N0rZX1DP4E0TBl66Hj
0fM46C56iHLKKYObfRTgBMMeJDQVP6uzNpKdN7FflXDl3qMbR7JZJAHAGv4AI3pI
Scca40ZpPIL2VBQgvawnmMp9mSZ86VsiqMdQ5JwOCKvNY8blZ7Qr33FNnzks6M9Z
MpffTFvdemelD4sXCIclcbYrJ7VBkX+uSqACMkRud+6W+HzC1Ocur/6T16EqI5yj
xB9fcqvHRaPzPiMqCc6d2rzwICt0Kc93f/mtI6UP9otON1qhlx/JHYRFpaa438GD
OxdXlFyTE393ntq0xE+gUZwokevTCLTi82LUb+pK9CTJrE7LFiBfTIa3QNGQscB4
FJew/Vx8Cv67JIEpoSKhIp7HrYC+msCpqR6WRc802U9QfVy7n0lwNdbheKWauhcd
3VhtbRr24rYus7aQvpqqVaB79S7KhN4SH6KVgKEJRJajCtLZMKMJGyM62hkzSiql
k1QBXiAOCwbaFm2AVwrr+w1XC+fQle612UdpcITbVpBj0gNIVW3j0HvKXR6xMap3
XwTqvrpyDI4k4Rvyn/hB7dEYv7+HIzbJxxra4Pc2wHr6nKpX36IpR0vIOpPCnAUM
9WEUvE0MNv3uhAH8p/Jr+lB3/WC+xQ1ForDZVNl+k4D3QEEGsdlROFWBL7rIMx30
6lG54HRu8XZY/r5uXo3NEcFcXhChxqkPwP0ULI1i+BujxN8opQ3D1TA0fPGa0q2I
IN7CpRtS+HDjqMAnjf4+/Sr0PVWH2+TKWVuuDz4YgngGM2YSyMElQgeFK5yQgYB4
sZoBC+Cl92pl6N6z7vF9wqyuIupyg19Q0uM0VkQKFQ+qx7XDJbV8nBCB/WJMreQd
N31UbMW4ZB1H0r1ApQ1nr6zXJKLAbagJhrkek/ybt74ABRuPK25gV9Mq7ATigQch
SXUsvxW1jMNgk3RuV4aU0nSDoKP2BgM7FucK4pE9yI6B5EVrUqp8zq77Y4hraB+p
Q6oxbGv/wqAvyDKCDkv2Zk0KINEvC2NMWbHL5NhddSn1kY5EMV3au2Cx97l6ZBuS
6YlPbVtk2y2EkdonYJESXxZsMFx9GKHqRwGUEIQoCzUo80+vs40IkszfiGMlU0FB
7ZkRbJijJxgXwNgcTJ4L8ch197gL1qLef4B95XGk6xdfWhSlS7Pi/1okiL9oBxMl
msJfvDtIqmVSc53dvU/6LJL0CrLwQP99GLzcCNVAEELGYknkZvvoXaX55VL4PWze
TxGEJcdx9uqfEcHf2qSLOUVHYPHkDFopDZYhbXOgwSs1LSchFfsmdR6FQ/n4f8pg
S5lRowhP6feRsdUKAznm4Mhrm/EJNyNknrBrfraB1vUTb2b+DG8aUykGkKVEDtT/
jhykoW0lYIBkGNHYK4aRm0/hpBgBoQ+uMHy+UGoarwGH6B4rX02cGI+zeeSOUhmg
HIG+wTmCmJQqSC/bj0V34nY0hpQ/KnQVU4PoVMn1Ajgea+M+wCLY5Xr6sD3q9Xly
7dh54bbi79L0uWxWriVANIMenTQEAAa2dgbu9e0Gvfj0n7ha8PN68JPZ6AjKX7hg
wTiKjvk4cG/8f1z3fbWEzEzGzPfuCglI2YYRo8tqSAidlaM/FB9+6VPsMlUBKGK/
XXlpBWnDPMJoIZlTqol5UWmReiCTAJ+/F5U9WKplPBbQo+KnOzV7Ta1w05G9RCO3
6iQ6wronMIfnfYRuyCpV/0DwzifVqJEDo6nsmnAcv3t/220foN8utbE+MxBdMg3A
NPqi1MnXKxRIeno+RFvYx58miSo/1Xx8NT2p5T9g6i2Favb9hRMfSZTN+L1MEZ4R
eYmTi4kz6k4Te7LHGqAKUBkHvkgE5xGIPO2ggr5UxwK6l6J2WFRwrODLUaBvKWDS
QFZu6UkuHERD7lZ2AZu949pu4M7uVz2ftorng2QwVBq476fsjmqoda+M68fWEe3l
kzI/ZqizNfWvvZeKTrP6vzx/RNqQTy1uSEbdOVhC1D0Mqnr0D7S+k6OoHNELV7xv
hS0c2Ucunn0Uk+bZ7awTsODtVZYe37nmBSFGn2rnJyRLQAKButa+7yRAlEEjSjKw
nHuV3SFnbxjurgws6E6SUwazI+3ptN1HRXlfIGDXjbGEnOKfq+3yUjpF5Lfw114d
0zz4fvNrw77ywuVJ3SJs0gyEPwbYnBLd9ZTSj+ZH6yI+CSONW68jdDiLzY9EwzRK
8sGiWcIgqKAjM9hobuoNfAC5wo75wScxThBeIfgTpCfA5JyaPYor7lj1xp/92+u7
68yOMtEhgZHrITxBge4xnDkBwc3QKYQGyeS4lskYpWYRkr8x4I3KYJ2flSpXM64c
JrQ2G55+98DhkjR3wLaZ40Hac/jRpItY1u9CAJx9le82EFKgUmzRDIjMVNA9pNyB
AgwKc1Au7eoZHrZMhhXaY/X+sdQ5UPyT2T7BRd5X22lvxPJxn55pSkGj27cJZ2lA
mvPdhSBHe2Nigwo3aGXl34ARDNYGJ+Dut/K+7cwVmhXalW18bN7cvNwdQ0OPyieh
2/JXQjLXhaeqf1douu+WnES2P6Xwkv6k3mTvlAbcz+lXRw4c1QiPO/f8Vkkt4IFj
j58h2pzpbCHvnHSTJmlDWjtN1bU3xHCwM7AR4nB2xRk=
`protect END_PROTECTED
