`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CNlt1JUPnDfHQw6CDmoOBAEsTgR/aHy3T1TJMpTBEHcUgJP3jbqhayQUOEBmIMIF
a1hJmem16OGhfU9/KNB9UH2T5rTW5246aldQP9MO3haqB2ZHoKb9DSMfgfCam82r
mZywxfDneF6iK3jEAtY6RDelcApQZYIR1r3kEuYfe/UCA7xThNbFAV4Gh7Yx989y
Ry/oP5Us5iRPMt1N9Z1SUqlJG6NvySDIw6dHjGpt9qo3xF2EnqCoQHe1rpoW8yfZ
sYGhSlwztgS84cieyrSyDkXu3ZfSgDxrCnr0xRIFOgt/ziNep+mggOHTWcxXsxIR
j6/zpzvetidN0AKtRPeuI2IZHOX0vD6TFcKhI8tJyzfrwrgerN1o8PidX9hFN1Qn
kUDQeHHPFtyfIvzerEvWpdo3E9qkxJZSY0fH2REQIgW0ruCDBwdujr6tDP+Hgrkw
kQpnGIFrREA4p3yD0P/EQKM64an/o0F3gu2QTC/+3gJgEuYYHCwDUl/oDOR4l773
Ydor7R9NEeT6lKdY9H8l9UVQlO9zZQkXbfw0wp3FXJsty02YQnSCFiCLOnHFUw1l
rh+TfQ0kRNFcivFX1s7gYWTT3PnZA78osLG6pfsT249G0qyygFys7Ij/vGkxCwNM
WrV1lbXuQd3UifzCZRtPBlR7nMWsHRt28rrVV/MN7VFZE6xAWjdbhlqPGtMgOg7Q
Ez1tldFlGIhswgo5ETTCoL46/Gu+DgAFNUt6uok9qKLK84eKQd4vb2/w1pDxjyML
zD8jy/hJ13MpX7H1zyzTKAaVoabSOaLBgIxsW9vSURpVZ0eTUIUHZ6ZWgTVXs0Bz
179IvKywH2wcHhO7Jm+hTbcDC1EPQ5RL8AwA0HAnLaZ8laETNohjiDMxHmXkPYj4
DBR07zzX3wvFdmvn4mKX1eF8QtZuJ4SkZd31t9sqAlzKkAkzJHANVRj4OZB817h1
ydgWa37KrIt6B6ulMo66Go+/Fww9eIX8RML0RiPE4QTU7N/F/IczJuCXBnDH5qzo
BchE5snQxokcQuNMdzGB/6jRgsiy5rssX8gWAZcfJtuFu12hI0MhaqICHY4RTY3l
VM9yPx6GieGS3GwDlK6a5wHj3cuSCtQkx5C8BWrDNkj8OikD1pzVjTFDSPguVKkd
gHN+d75IoG5WPto73M7hZppeCNmOqZGQoopO1do4zpBgWxbvWVwQDRLlejQsW7S6
LVCFEh7XIWIrWqak1mcFWag+7KALdjLxSlC8L8hXeMDHPv3ceXMIJy++L7XKsuxc
xOK/gLteewpRL+OGorKG3mwzhQUmsXycwT9hgdbGOAyvso7ty95EFNzdhiGaxMb2
7N9jCWwvW1gWHAnNdQXmnO1IGSIdMnki/OOQbg4kha6x69IlpfDbbzTgUhf6WFa7
sYTqfv6tpN7oFPeT5m/H5lFyfnfij1Skg7fEsoau6U1u4sbdY5uyt+urjTx/yRhL
i+EUAzViFsDmdSmIavP29SZcfizyf5/qsCqu18jKejgI/phExI3hhde3fCufwxlm
OqWQuTMoxC6zo83jw34CmguIKqQKaxG7xzR5z3prvzUl1xE4EB5xGu4zuPmjQIMe
en0pPHyCamdTJBDGTXbeTGkVhqorNSBYJX0ieimUCBF/MuPxKMWV94bph712im4w
FUYRVmD848LnWdSdXt2s2FVzb0vaTXmg05RE1Q9SDNZgUOz4jXRTXJopaMYnXiSq
RJWD3A+WvA5uSYw5Z28BkJctx7yjcKbNle/OMflLrIjCirjL/HxnapAFt6NCGRKi
hOFxbjJsyM4LHSltdVXVD+Dai0A4bNf7Ii2O94ZDRUAV4tT2zLfaowG0wi1XRwoD
to0SbEUChlYVLXE+sud/DzYorwsZkr6eUF2TIM/8K5lx/TFmf1yRxwofAoiEg661
YgGFOh54s16qymK5vueuLEBoEKA305hLYLSFOGaHL6Twleu3au+cdxv0BAVKqJ0e
biIPBimuV0KvTufepYKwL9GINQbvfRuJ3knXVzmT59AyJVquiNo3llUh0s4KzZAI
wGU92giXBekatPoO2Gc1/Wkgtkw8UwL2+dYqbUbx2g1ukKEkwFO+lxqSoLpdSNVm
cxBSR47gpnjSW0CMkdPywcdE9uAQAWRN3P78MoJoE5I9PxBC8rJDJV+AEaoV7ebH
v1wc9qNscD3DbphCpk+HyjQfwFE3/UNGpBk5P+q7i3n/k0PYskq372uF1C6SNeQ9
24bgJiDUsoypjsepn+Rk4WvOWkG9cdtQu9WuelSB77kfOMX5tx6+FpdiUFcC3zcX
blgD2v1iQvQD6Z6KeTX5yTUM2LBS3vFAEste8xNm84Re6AWhLP5mEXtHUgkvG8Qo
B0N6eBu2aHCBUEz/WWmrzTQhB7+G4xfgrKjsv4PB1ULER/oIIQMxP8j4CgPMYuD2
Wk1reWfCHPPtqg/cE2MHf3+9p+ebpJciejIPdSEY+06CBGOG2XLAr+lJAt5jpbB+
HnnKi9ku0yO/EEhAywG3N+K0sy4Iag8rp6XxKEd8HfYw76jbKH7+VJKGvUYuM1SQ
JZjtogfI53N3sJhixdy1lx8KSPiSHExxdZ6FnROA3sfgoAbXAZeYE/Fyj+6ekKb9
90q0E7Oq+SKOEsYlM54jDfH7WuqwmrS2mXLV+jHh1xVUMKxRJTe4pWhLicHmDya9
Zs90uQFm0HEjmLyeOv48EoylOebehgtsjAa9QGl7i/Vi9JUX2+2/tnpXJ+kf3z6o
l7OhwpSt1/QuaGd3Pk9nXoudY6aCxDVzYOWpIaclM3GlFju/AOcbrpUSNdCTx/gR
urP/ZUAfb5d4nxm8N3hhMjAkZkqgnbVECto48Q4MDmg83OQjZW8RFxxJj2u3pxDW
Np2nYO44xR+9FMXlLMqlscb19v5beuqmgqZZIq/uveG/Hv/39Q8Qa9MIuLaFV2Qg
R0tP3vBGV56GUsfidezii1+pERB3RRCkiGTJvZU5P8vuUKbBW6zaif6YoF1XZdIa
zdueuNwYxKbGLgBPh+bGBIUVOLWZquZo34Xds/sNijsnSD5Rq+SQ/b8jiDwbMPjb
e72VnoadZ2/GbvKvYrxMqVIpHnFp7PcVfgozoIydwXvmpBMz1LdOmIvwkIynxKPZ
hL4o3cQ7KrZzsGo+w75SQASJr5X/qePBLcMI0kbfaM2k8Np39+OTsw7ISPKffN6v
WdNQrdHXBkjhXdNJlCjDw5U61oqLhv1RvaTNJ/TqQw6vLY4pcF04HrHwvssDWbJ7
ZrK1JsU2OZubexwsgb2lDa2WIcW7++vb8UaFHTJgoeZd+ArsYBCLyA7vIQumLYvP
5vP9XKM/m4eaI53g4et6ZCHrw4G5taimCb9x28hascKMVUlp7M8+b49vVY57GJCi
InANXba38yVs9TSQHjUq0r8RIsQeg/aqQKNzdNsqXap7AUuiPfug03CU1mgmNURf
lb8Wxdk7HXzpkBqtCs8L5V8/c+SEGHKxqDGl/jOtEk8YU+J0JU8zy9hWBpl4QO6z
mUyJYZPlqyZYMLvADGVYKvM5EALyQtR/bWqm97cjEnsDRfWcoA2mdjr4N/MpY6Ss
UL8ozdpRkqHV1xyK996ACkNF2w3wt/u6lROScuE/VyCfLeVjyY21nb9ubFHgB0NE
+2UfEc38JdZppG0O1B4ETlcD1c/yGL1Ea5D/8d/U5PiQaiva+vdJe9GzB5aKx0Pn
CpQPG7fc3vhnCetz3bLWgqm04s1CancS7/ooGUtzUpP0lsapmSFqcG4KVKzN40iU
+5ceoOlixG4D2TYRgV3TXmeGRWR0w8NtMj7X8v1NcsIVp7xJvtaNDjQ6VRakACDZ
83mdPw2Odu6YeLSDq94XbchY+us2KF+SHvcv8qrhEq69T3Fu9xjj7UJ8N5twBtCu
KkFGB0C1OadIZEQkDV4xOerc3wSdsR89RGq+7dciVYN4Is0uKM9nzu3aM5c7+p32
afr67JdCtX22En0+5KGLBYY4evqP4+xpBPX9EhmrvEX1CYyd/h1kGt8svvXplV5N
fSKJInWLJBunCFxl3H1OhGoCj6rN0aqY76gM6sR5/ypjHxc6RVRixP5tJPLcy4BM
rSOmTYq5R2QHqcVLiIIR4TlyaJ+Ana7WwbwgXItPOBbQhLDqVwQKSk8tT2Aq53mS
V2Rxhmd/79e6dAHk0zXCZHcDTYWWcr5KYCtDbxvROqFc46qOzvwWrhSplYt6WIMB
qJv9U85uFGB9pXgjzxtMtd7fg8+45O1VZwOC21H+RhhepxqstCs5W4daEKU5R0CI
VwjPXZzfx0nZa9o3PJ378oAoUPj0TrQQuGC6YEPnPmt9ytGT8LoHkm8eCW/Od/qQ
ytf0ZFO+7EG+RuCazJDITkjqghUYtOla+p2ISOVBaNaYgh/wWZjJEw53+w+iDTbo
FL6xj9vb3EpcAL0sSaHsaJXvq6Q2UmtqODGZnVE8EEvYVDd3xYuFfvv8QNrlmGm0
uos9Us71pxngFeRWxMxhoywcsjJKNnVF0tXae2qyB7CP9mVCGB8A2lDvG+tge+Ul
y21CTT5tzNEfBKnasSiYKaAulknZsAr1MCv4gfOZJHNJa9h6C6jOg7A2ZvX6g9tW
BclFSIB6EcQ3/hQhUsdLRQWYy4XWavNefhT4HGN+ogMG9x6h6BlICVMqv01RcQF3
AGJnvQMK84A7MnLUuhOfN/PKUVquB7O4qFJ/FfgTihSbgIyRmlXHJ98mxMVKemXU
lwaEl3grQbs9nvC715YYdmG8YEVzgqxtEmlU8MD6b+hmKHmrjJS2hbsaR98GHKVq
JEMOhVYqHzrOilIaqRh+GV6PQTGJoWgpRYJMMcnNLHhQvEgjKHJfc5wSX4jKfz1N
KFr7v/2FCIPvW4T/q52gPRc05Z59Uk2psUBGmRajbCGFw3ulh3VByru1VkDw0cE8
f9W/ODeuHrElV2WY799B2rWLQzgJ7LTXrOyf/1nwUKO+6Jn5T/U8VKfYaSYljt7r
YVbWmMKx4DQYWJ9ITqrlF1ig1DI3uUINepEqDGAomGPQBqknJxPPk9ViIbh0dATh
618qEcdxMcrg5gtBwuM4MmcLbps/i0S6KEcX2d3hJOGeJbw1UVeCvGY++2LgSez0
o5KwpE6syKRiP4bemT06aQOX08zHJC2kQKn9cNaAX9q16OTCsB2o+vl8zH8EDFyT
XMQoNPSML2oupCRKNTFEE7A+VFoGGUngO4Mg5XNeWkqZYX9gyz85gYMkJI78W8o5
CMdo3twVuNumf8PpGqLqdHv2d9t/sS5xPaYST6LxYG0/ejRWAB6zmChaZFQphgiI
mQJedPCfyp9i9kF+0lGquyA9fbUkhjkx0P0MO2ELPJxelxk2cqwoijNMhzniCF1t
TKXtVMs5HdOx9nY9kBHOaaEGGx5IHwxsnCpWbXsdPWkdg8LyoucQi1eT2hYMeP8T
9inPx+RnoxR8C8x/YAzr09laYpCO4E2maP2vRvYdz7S1Jg7FQzV5jCFR8TTcAtBR
37mQkzVt/ioIPfVIiQWdAhxauvxl6x/2O2ICeL+QtscxYz9Q8G8wpSDKPU/57CbV
QRaDE7hE7kt4lrRZO3WvcSvvKpSs9NZ+QjrcZsuaPze8EN694Odta8Vd+ns7NQ+i
xtZSAj3f+1Exbkkh+JHCSPQjX6pglKnsHMw4ADmbqT3gipNXtYnyPnXUR6JbvNMW
0LaIMITA/yWO9C1JijUr57vX+/FHJ5GkZO9ggM+dzh5r6tYkz/MVsZBNuCqA7alL
Il431b8zvaVQEHaJ3TwU/6mcramBRtvlbvCXTHN6RRFveJbwmeyrddRqD3rTwgRk
cxcLR2ehc8fPwAy/xmYxn6CbeqFQiHkdEEQ+rNwVE5JG2Jxs8LutwNB/43gNu/dL
ozk+WpCe+5tlnIU/h9XMyGR/utATzJYT3nuV61o3oa3hIi/6CUydiAvlSovfkjf8
CrxyCLAtJCAc7q2bzOTz+xlxSwkq6QL5nme9ZAThA1Xi+r64tHLGwpBMd7GKrCdI
8PkxTEf4f/5HllP3YWaierl6Flq45lc/pswdj/zgT8esHGwFSMXwlo9dOqMVy5pB
uAlHBHEhpQyDg+iEQ/yVdUCT4iiPlStbQQhbQdWErxQWb1l3dsqO7B7uNFyoUHWI
IE1F3Z/6AGTN6i32prRrDr9Hbi/b1+xVfPaZLDaV+f6Zui6J9HQG2MNjTbhqgI7b
scIesuStIGS5WYOSJ+64p9rL4dMXr35k0DhtkSyqhi/ZqORrWCdyRIvGtw1cgkKw
T93UXYg15SzDMBCFP41oGYTS8cj6bUOZIAJ+Yck5wZRJhNgS1CgwM1gfPYQqiNlp
fY5xI1Nyduhsc3Hc2h7fhe+/hcgDJqhK0Ov8A+GbiVs25yk5iEU0579OOaCn1p64
xnSGSkJjObcZgt1s5mSPocm/KfsIJTjt6X97mHi/KzWIr/dKzw9Q0ndGm4PT/Uxc
kA5tHJR80hhsH639MNJCxSFTok+Jnrmne1WyTIN5AfbmC8s05fzNOEtKlv7eK0MY
O0mQitViamMMrOLUmczKdGHxEW1u6/YfrfPdZDrrztXoKwzTCZTpmlWodt6/uvaT
0HYDwgyRXM9UbwlvvAyy1IeJTcFIgIEANZPjH3Ldw6t4r7BGMMBrWPNxtwNTdC4p
c/LMAZPhqRMuWapuDFWFb9sfsjL0LFeaBoPTsAUphnGRT3+wqgwlzgblipGJRQZf
lFcTJFQVqi0q8pO++aYdIvEQ2sD3eTxUHLrkqHiUX5iS8Z8iBPlSUd43zFx7HD7G
YQnCtOsaVPpkX+/90lFqWhtGtMBBkSdwIBUxen8FAyZ78FfnCZvMD0IRPtREv2+k
x0atHZMk9Rp6q1RAyhsVr/URyho/ybVGNrVuVYxzya3b7J2MKwIapqQJsnFk2io8
fo+iBuDV2vykcjfYXcex3qP6OrM9/XIycgPn1PctBEU14I1UHMflO4T21eoUpsxb
6SPkFNxVCPdE7/lZBtRLLwcMxnriZgAUV6My4j36+t53T9x6QAY+8FILmKQMa8Ig
ATzz/dNACAqAusot3Jk58Q0fEf0XSu6aJExrDeGri+ryejGzoLacUL3Z56IlAxY+
1ThwijmAPMY3Id9L9S2uxetep/2H+kl9+N3MSMkCRnxo9C2GdkLl+uzUiBDXYpa6
Vf1WWC5irjVMmr/jEDdeft3airpC/41Lg4xgWVp2aan62YHcPiE9qyIH2YzNqkdc
J72c3PD6r5UJyAfvPqOEaFC2/619SbAFUv17DuLCeR1VJbnl0jWxMkVEbIP8DX/T
Q9TkEu8T0DLIwCTg/MeJvWoLyOOAqMt7zZpAHJldN2/qs2sg5v/HSuSNDYbvvGvX
iY6KG7X3fNYtPch3B4uLL25MxENFnls0HDKQcR3Q43aaPm8MtJAuOarUbDnVkTLs
D/6J2/7lCwoFn11VZTe1pyCKEQlP76uWgU4rtHRZtSCz47irWqeWj8H24bf8SPuI
NP+TSQ/dWnsqI2NHwgzjH8CvxqI1dz/zc8KURGJOhnnaCpgTE/8f7VInpVgOQ6Xx
897cHx0p83qF0tpr9/JncUfy3/A2gFprlmhW9YkmaiHewJt0+TXNxtbGxfHoOMQM
RGA3poA3ZEUvyhiSWdlxR1Y3a6VvvuShqxhcPZowVzfuxJGiTBFN4RFeBFB8IaZL
L6P0+ODw0YIg/uXnjDHeW/AHiJLTxwilozp3o/o9Cr7wOOZ7G8GrEFygQmtDdhSr
dDROZeO5xiT6qfp53cL8wXrSViKUfQ4GXkb3zkohEG+QS4OEoQdPB07nYlbzBJ06
dUAtPMUfndNosW7O6S51pAHgbfARXbNDC84EcYexTpEfCQMZPWRcJw0/DKjcZIje
0eZZM7jusD1/G87TLdYqP0qir3yQ6z8mag1I99w8vlWQ+qsCtoHmXPuZ3CNOehDf
IC4E5rbrDA/ZSLGVOBXuYEmS2/AY5fhQkN+ZsvZnkMkMa9gvgwNQNrTT/NfGv6ar
MPWytLpC4a63KD1OdOCpNZVh+JB+Vls6FVFnihfbNWBH+mey6yTrENH7GdzABYie
EdoY6hV9vT5ZeGv/K3krN09tiZaucEAudS3W4kMmosOLuErQV6vj6bdfXmqRkyoW
0UWsJeCjyO5JEx06Y4s2WruaMYOlGmNabwS63MtUvEjEIl0WPBh83dTRgyu1dYhY
zWqFi4FAImRcbTYjd55TFmgbdHC7+0V0mS2khSYxY6+tIv2wMu6cvgc01ZNRCn/z
SNwnQPQ9Uo6aYx4WSJhwiGX4ZOB2odVMr8h6HtiwyQ6KVCFKxmwUCTjoDW0RLidr
/K15Dn4iVpi1lPa4c7YsHhoYhTqqu6YkWitfa7+G8ySV39TPvR7YpVVS0LU9xPMp
I8KSunxJxNkZ2b+ALgqI3yvi7jTKzWhfKTeM5H5inYYdGVqGgMy7Md6fXO5tP8Pc
xvHCzfc7eTSOcRMezViYI97zbswqymwsoP+gNJTQxXoFi/9STYxCAO0IgDrqLpW9
AjuOnasyCJ5gdi2dk1ePpa8hrNm1bUZdziHGzFgOTW0sddO0U6mH1QREsIaD4t/u
ota5puxcJVcISai8gjf1WC8tZm4d4qVhwiZyVlPgr2rR0MaP2p20pWUplLPwx4om
Xv570+5+pWso+7K2rCTImPu3Hs75c9od1QKkhwOLiJjkR3AkVqbAwhpOGtJP8q4i
ZJeY+OFtxSD8F1VdTai8EzGbCBeROFd0jwcnXJE1yl/M72gVDMclAeyszx1EiKH2
wcSPGv52PTaprL575dOI1IIADM4P1Ef4AH3UAGfGd3APn61Yw4vhMJRa/bz/sSxM
p2K/4jDmhXxsI9hIphaocUHQh3IXjvOVuxIQ/rK8Nd3/b30EpBXLBYQGN+2TqyYr
XJfsFIRBUZPQfM06aAueZ1Xk7CvpJorPO3+EqRQVG9Br57nYOywaXWJDlk4ZjR7s
nphOsckgNDNjGKTwkc8lBm/aiLM4BsRsCZfH6lAd6GiglntSQskGyJjQwKp4NwmZ
YDVR0XwzKoBOaG8mGYMIGnrWr0vDi/X0PeWBhf9H68bkZuP7jK+NZ0A+QHiWNDXb
5hWPdzDvpCYEvi3yUypgymBN3NH/cqjz9PHIB6Tmy8fTFNQv9nd+jBqIhCwRrkHa
PMVnespA/5PhlRahnWJj2g6YPxo7P9NfAuyeiF/6SkK9slc6V2eVu58XX3SdGWBk
+SEMhYVaZ217f3jtQBGPospog5333GiFyPj/APtuy3Hu0gtg24qQeUKuFu8Ye2lv
x1tLFrhMD5CAYrh7PoaEOObFtyx+KtVTS8QSYTowcLNQMXDLjIkFssedQHUJaYdA
aB3TWTVdMDLjZeCo3IjRgMsecn49n6RPVhYE2bdAXD12SPbCobKVnkjNyTqj6GFW
ldm/J+Ba191lx/oDVfRdKLAjfAxZ25OLDU6My3ZoWCj5U1gIyBr8Ee9Pc97p4m0e
tzaPSxzRb3AXh6ZdV2Img3uuuDY8xfqZ1XTYzj7LycZmsdix0zfoaLiGRKL8xHfl
IS8Rhsw6RbeGqQaLRj/bPieM8gB5OZD9cnWMWCKAbK1cbPMcswNo2fzrHycKb6ic
CK5eCNxEAgZCAEYHRM7vdjqvuqI5LfMMUxulJEIPIuRWRagqPSvVMbPseHcPfJZw
ijKu1Ax86P8tsN+oBHS9uqS1WAlX4YZuAwv8NGMNJ7xRucogZNR+qHEgJ/FDNdAx
AYSGImIJfyb1B/VtHAt6kzC1qPKk9Tzo5H6dPUdYkfZyqD3Fc1/1AOl2FF6ZsbpZ
eSLDEy/s48cZhSjG4vs5Re2k1j6IVP3zCcZh2xD3hVPpVph9LObD6mHEh/iNhFYX
htv3iTfaBWONrJj5SH0D/2cXdDrKW3qApKqwgMHhxElJtICslCqRIv93vCb+fem6
WAzMhBTxWTLOK9gtUV/JAeBvRrse0Q3wgdQXOhK2N7zRwKKvxLxB3QDKMEreMTai
kApiwd//a+dtZdF//gOF/OUEPCSI17/Ln4Zogeqv/7qWyND1qYClO/Ne/0YloRWy
S2NQ+44jqZh4pbTS7rmYElF6k8vkapvUZhbGndKrmvdzCiSnSr8THDBkKkemaGR3
PiznXapBXxKed/oBtMUFCqNL3G3E9sZkAXM8PQXhB9QG2I9FfvySrF73HG4akWMp
Eb3PPzcW1DiewchRsBGjFPzjVp0lxy29lOIxa6T+XQiEyGlSkvtGwfopxh66YNRP
m2/71ZTbAzUxDxGMOPLDusQRN3WroZpNwE6fGfEDBQUb4/pHyu4WqLKefxi8/dPI
nm4CWyimvsv5sCk9UAlSzZ44zLN70OupHybxpah/efL7oF1Ky/m0VLcxNFWO3Fly
qe4sTII73MRibjELBaKNiDhzd376mM6YNuscpg3IUWpJFAYAXnCMbbsJ+9fz1Mjj
qbWbkHKxkZCxJ+4P/MwRtvh+779ZfjrdeWsv4oKhsf1rQnYOGyP36RXeLwbCsYrZ
QfUQOssHJvFel9lqw6nqgdkIhlt8FVUM8iwh+yfydiKOd13rXHE5jfm0+J21/7y0
CgTLWLK2fqImfdWZhemiaEOKqNS9nJnEqEd9KtcIzQruGBl0O4MtBjC62RVQTH80
VKyMnxPNKR7TZEyIGTLnFUF6zZacizR0XzVDdFpCs6AlS9CsEDo2VkvZIrDZfNbD
ZxHsqPE+OnfYJF6E5L8V3t1PeV8OTVeoeNGk3dsnYZKdihb1dGIuHQwaVbEKFqPI
Tlf0O3xRdjwVOpTrFYwcdfpGspBRd5tz94C0qKI9KHGakQ0KmXTl2VufgTT6Vygy
ap81qFu/dy+tXbKD+BAqoAnXLEJZhUbhXwXImLbCb5AsCwBJJ8GUra1C9iCXgDkW
cukLi4DmMBtvGV/xhYEp43rcjpvdoLHdVKQf7lUKu+tPC05I8qAHxFPvBsRJKAgQ
W4jiCz+saSoM+Ill8dBhNpfhYM1WmK53p9Cjx80NymMVNsvmaNcScppD8Oz3oGW3
nqS8RkUxNcCBoXGD7eUSLBfz2zmdKTLrI8kHs3DrkyW62UmG7XPAsCNUsYSDByxj
TMJWZxkUyN04nyjqMQAeZkWUylJD/RQOjNqk2WXI3QH4TycTr8ZCdbIqiv+Kj5J3
F1+hUEEQqOFHg1tAV5W7UY7+1CVxNgKaTqgARfG7M+WczDWrq8yjqhLMcaO5ehKq
7mDOQqj5snwChbiUwd3kfOgjsL2fUccbuK1kEsmOfx3BJCcvG6+VLheCnHrEojmC
1DpmiPuyl7+wKe5veg3xPAMITs64WifXRQjQL0qFgSoJB1d1FWcnN9Ycm6y53fRh
ZF7G8HofLjGFwf+e5oPc6qB19PmWRRDXNhYVcV+8KKBEG35wUY0zIVuEjt7gDGEa
qtxqTcg8FqagkkqwKHukza8W4Ac4HYtRSj1Mzxrj0ekikwzFpTlIci6NWgEGx56A
v2ZWyZlI8FsALXRLl7OG90PAOmc4kraefPNOnRPslpw8g+kXJkP59QnSdER49npe
mxP2OXsn+Kp5KQAooT/HNewjR4UeJFEQ+9Zup2ETwiHs6zA2GqIljX39VU4loogn
mQQQ4zFKRWj/trxWGVCet8RD7nTTrBxeqm8OlEUh1/3jX7S9xfHuLQF6uw8aXJ/c
9Y+cFBW/r3eawJnp0qX8nmKMY3ysg0kEMN7zbMYwyzxkGZGdp75XRkJQKH94OAzi
rsHK3HDu2IppHyLU2KkgmaOBPAjxjYzar7Hg7qA8AYBvhBTSoWfBctbnLdCELUp3
qLao5rxiTt/hdRVp++GAhlgjPAFy9BzZuXEqVGDISC30tZHAoKQAy4oXszy4R09Q
v93QEaEoIgFrgOxP4uJhCmurX6AVVjWymcleugPiylncBYeW1XDsYGyo9IOIuGH3
jCccoBnh8xCb5+bTPJwJ2IooiXjbO+P1RWuatfL74+ud2/Zf5GYmY6bvwlB8F8Ok
Gkjyf3B748KEPCVG6iB5V/k+Dp7VFR7bSireVaywvHZx6Qx9PAahnAX36qrj9pwg
NElTisxn8BpF4xKBNUUwzPisxV14uiUSSLfpPes1j0mUh/O71ii6etyBFzV9Oiaj
Cqg8SGESai885dm4rMYxxllOx/wkX7D7YlZTS8u3WvoV/xhdeEsa6fIGvo3cYYA+
FhQILdggN0dei4//LWe7wslPOEFJ3tphPnRr2jwTBOwiPALuTHn+cpBy8+w3xQQV
9P+/cuK/bhBeyeJjHTaV9PR6pfBBl/9zxOvoSBe/MDyft820oNF1pWtzXCBecxQJ
IeNUN7Jh8B68MMjI7xkO3Uo0oUTTdlNRKmYPgbGbtmGVPliw0KJR+OzxgKgJbD7G
NMWyaG0TSz3I9TTe7d9tMu990rADPh0wv3Ite+jYA+a4+3fMKpUUK9BOI/yWU0u2
Xwkk8sMF0OSfGCmCKNteORYI868Z+IXomujXNC9vSzZGwPLMKgxOGRXXEruMHFaJ
cgiA8G97h7fLcfkrc40VvQeLpc8eYPfhdueME5i05ZlAb/JZOA4vbU8fqmZan5Q1
lU8HM3xylPOeEjn6T4UtBg9EFIbuZyzXqVT7xHXCieaSTEeWFayB7ZvfQLbFX5oG
fkrTM/QUXClyZhG/tSwShX1+wCDC0XtVlFisYmEjQ997RL8KFKUe3Bhgxq7FWsfX
kkbVTi5w4WMlbjwljLwSst1wa2zW2vZf0cTTIrBFtg20hAkvNU5a5EXE/8jJ4ZIG
ARyC5FiwXTYYF1Y52eTr49jcc5POwd81oNxFc9KB8k39GLOjAtagz5VAGIl1irby
wFJzz6rh1pIZov96db224Zp7x9hOotoxk4Qd6mSPW/En8Q3yHEvHr+2GdZNlYJ3I
K7y7Uc+aJ0fYcoYs7hhmP/h5g2BhGe7zpz5sXjbtZpWPoaWjzwUBk9dF+9F2xiEa
/4Xrx5JIxGkv6Kbyr+G+LM1caZep4QoAIGcGicesBwTYF3m8RdxwET1nI/SPAsbg
C0CyV1WHutAjZ90ZPdMIxCw0mUGz00aJEZjGk765/kW4dlhxP+PU+NoXGoI6oGk9
BuAiAeiSbXnvjCypoUGPqCcwHyKvJmn3pC87MdIPJIfhpez8coPPOfj3d1fRrdwf
N8pQoeEZOWWujtFXBTWva0Z8QRpIYo1x5S7t9uKQmjvkPOK1LN6i2S7JXPK4QfcG
PPqeTCozDr+sZHcwMDsDMtuYYvM3OKSh6O5dOQh2i4YnXfy1d30kdxWE9PKb39Fi
fwc+Fa3Cqbr/lEUILKN4C2SrS/W55l8cPoTxLsC1tZREnjkKGvWF51okHSHkXvVZ
dflsbZIuQtftPhG+9mmbVMMv28Rb4jjz9xCViDgXwLS6MraoJBda8F+P8JrS/I9f
RqQCDF7qlrbCM+eZoTswIUdgFgwz7Y2BKtQyz4AdzU8cuZvBzGokL37QwJaGzWYR
XLV4QV/z35uz+bqZtE22Xh85SV/OKpGHTW19936a3B775Op25bU3yX18z9hVhqdj
iZFGtjQlIYtIhlqvo/vrAmdkC4deaqS7vqbb+obm/a1VYO2SkM7ibkevBUrn0a3M
R2fC+hUBEebyf6zT6mdC+FWatAr31UypR2LbTyMgafyo7Tp+lBq3nOcUCjb10Qsk
Ko4zfC0KsRyLwl48pJ5iX902WnQAnGNazHJqzIJRRisZvFhoqquSneCQRdW1zH/u
jwGmeYXG4PgMQvV1UfZheVeLgwBzbgVI5QVjfFnmP7rpk3jFxBfymOJ6CYyNCPlQ
sjjdealfywjEe7pzBxxyrqedGvMgq8XGetzbxlN4JjYbSYvVtwLAwhjtwCcSmToO
PQAo8GERzkNS5lpmMOZIJvemldfTaVDDMsR2wnY/U/RXPQdj/DBwD7mLdopuDGf4
OEgBfaIFbMyayUK27m8giB3DNXOq5psD2hmGTjF8eROXcgC7GgZqcZVxVOE9ekn1
Fi38z9hHPtPedSiREuNqFAayg5vd0kZTteBvlpmtaSmcWDdYhyvYLlXWVJnHvdcr
uK00AQdU9tJwfRjeBNysIS062+eOSDXqPylzMRhFRXIJzmpqqqFDALCcpyKiAdu4
/nkddSJuXer9bO1pIYksjQAu0ME1a8Y9EEBrv1d08WOCUYD6eAZ5CD1cQuP8DZIh
I03aCzdDW2MtfaufNtK0T033DilTktDTOHU/IMEJ7gN/Zb20O3IahvfTnVJ6Q0Cf
ygp9G7Rt67iD+u0a+QfQUFbjWfiRqt0npqS4faW29xlWEotOxMQ/gD4+q4tF0eDK
OdRE6ATA2z2iykhnDli5E0F04nH3jLNJ5RdOUXP69I2aGRVfC+gxn91N77M/lPpZ
kV6Qqi+YFN6GdKV0rAmBePrJDGjWEOnIKT/95KD7xePqUYkFtwl0BSXMVnnNmGTT
702AllRT8TFQMbZIqaLiZBmeTkAfLJFQAovZ94/wVU+eSQryo2fQ53UfHact9Ovl
W5is8MRLz0UBxxe9Ec0I0aEwqc4ZDW2F+yDyo7I67N27HINGRpnzA5hpS3IO0VdM
XM+VAOunPtCzhL8YOmuZQsMpR7TLQfOuzK2Ipj7EZrec5hlhhjysdXZ56BMinpXP
Z5TXqBtZ5YUqX1BhQjF0ZfZhIFGv9W3GcNgB9/pmKsmgWbnDfiA3MtiBLW1DL/Wz
vL+AvdC3jXijqsh/0/yMD6cETzvhpvlMcZvPlgAf6FUDJ41IOlK53ItO66+NZKo0
hkNtZGneCnYa5YF/P8wguvngJ9+2yWl0sQMUOqT6A2FEkpQ03oOUK7E4VVLd8iaL
1Clq70mUy/XExJevvLZmCvTXMdc4yBx7Qj8EJ+9Um1gQ4YFQc/0rD0ricIfSY6D/
C7dPVR/w5XHSuwaHtD5vkBACf242VrbyRQhdF25KXdlq659yDBTwFHSTUmS2iCwe
9j7QUeNEm/yTFAKgKargGShn5zM0I3kUDUd0Qubid7e9j1Yu6g3oE/c/LbFCml9F
tmnEKY/ba6aVSqOhFMOfZQbcphMnCWtfZHcdyEfMjOfPIcFnIM1PhMBjwKvUH7KL
NzgJhKA12Rjkk6AsdlHi1uzwejqVU0soiFHMCrpOJlsmn4EZ6AOUmNgmNAAcolI3
fA7jZ/AVQlSrkG7I3ExHE/ut/Q+7LRe5YFUq+PjCuClvWX7WP5hQ1/sRB7c8L5s4
hx5GX3G+UnC0TqxiPve/yAoGRVN27hVGYO0RcVQgTSqS0i2cn39eZkMgoEti9+B7
88S9ZVyUMPbHNb0T4PrwSPhgWmEaAthhF7adJPEhrEJglNr/EfRMxNBh9ClKq+Sf
cT3XNPeAXKvc03NLrmHoB8jjIPs/YCyt5JpN7S7kCr/K6CSl10/GHUqOVM2utAX/
HvWPbBKA3ur08ZsWyj1c1FlsTZ0zUrPyzcA/6hTkc3ffU0E9VArBEtreM3abPqSd
uc6d0JPWdBIQ9xgrhPne3fQWJg2vzo+dUgGwfNVhZgh6ig9E+bKnSL9e77WLnXo/
KP5YoktStripJRBI2VPueteamfaat93HtMOuRAPdjhiQP5ATQjkw9gA60NkLvkJH
iAEQE3X/8RLFB7fcinL3rW8UTHepG0jHBuQPyjnQT2/pUqzLmZVd0ZQvCZCQxB3T
82nOOSi3hI++VkdhWfjfA7KFCQlgrv+g5CxjRNH7yB+cfGJ8ELLeCQqbbQ4ybMI0
chEC+WGH9N0OVRKlyvvi91COSSK5R47F05K7rM9XwSD2szEYUN2Dy7KHX+SX/GVy
rWM6fOFLP4L9TZH3WDD4xOVhw/R4bxm2A9HRn5z9KYOVDKuwOO13UqWE6h2waR1/
Ama6Lhf0SsGnUgQs7S4ZA9reSBI3Imlpv8Yme7Gf3kOfmAZ6nNNJHHXecjTXQkG4
YGbGXwETyI2X0ubtX0gSEDeFNvGaYXsB2sK1AGAGeCfSPmDi1+DjrrC2XAJ/bZ2R
Z5YMw4184JOFvJO2dQvlUNyVFkiFNe5LubvXbRg8F7G5zkHG6Iy6NscszTZPnTF/
WrF9m0c7LixH/tteq5tuGQpoD+IfSl9oUgnj1pYDnlBsc7kxyustwBZs4TH47G5R
DFxKB7ELtuB5G98Dp0SuhoLdtY630V+jm4bqzoVqCmiwz59sfNjW7aC9EgO3pFFS
bYWMWyrTfiYGPvPfE8F/ROt0pRzAbWd6XQzTFnrK7G1W0Bno9wq6miRoWRh64PGc
8ZOOZecWHPGBT1gser3wOT2+atLNpUc1ohrbLdh44zPrw12T+T8Gq3rSG+/4cA8O
Ov93Jf4572FVNFG2SDDcqWDGKWCldsnsF9AEXBq0ZW4JDxWW8OMENY0BnrlsafyI
E7vvLsAsPN/7pxo1vigSPmHTS4nn3WbZvtpnYNPtWfsMSzDUSevWgCET843gHExW
ZbkU9Ftc5B1D51JEuRTAQG+qS43SGEuTd2btYRp9OOjh24BWQ05PtjH/0TDV6SDS
XSrv6Wls8MnX9Ys2YWCgSSrbGEJWcVgfd4+Tyhh0YTh1C8fzaFxN0EWXz2l1C0Qr
8f1twu5yq+kIihPlKD7nAx92oh+Qkwmi7qz3og6VTCdSc+kjybYRUfnj5mv5a8Dd
aaxIl1l0MIAXKTPtQVt4Ux8+PAqIeQog5wP2DKTaDnPh1meZH/nhSTPONOC7mypE
E2s1+DJingjoelxWXUKE2ASPFQlkcaUplkT+G2AHKXjuwg26kVskmS10JdPdGzKX
0drPkCa3lsw2/gPhlNgjjffGcbfrzpYHdjWEhlaiplMG5IUw7aUSUvCHUZgRdqhz
wj4xD9p5phC/dSeqzWyutQz6LFo0eGD3urgVfCKgnIDL+qITdDQWq8VhhWwWK3Gu
57ysghYfvF6gkxa016y66G5juSq9I1mrHuxPZT7Bh2XkiZY7mnXUx2CO6hEAR5cQ
bgL9LhV5sZ5NMKtwn75pH3AfVJDD/CUvmcaMHKNzm7wk4PMRPebOYfM1l8CyljPO
FlqtBcl2rs68FDETJWj18R40snktdd66chRmNR4et77zFwOHRCbgxAW6DbyvngLk
rxeiAyk1oQXf6/2PV55zq5TuvXNywfjaVTHGfy2yQV6GEc1VVCwebJ1hBgddsOQ9
TQ1HBgoadna6Z+L36vCJhb7j60cYjb+YeVIzn5b4A0D0jB6++myVK0rjieIh1uPN
CmfXmetRMEPfml8Gbic88JoeIz4g9/9UVTUX35oLGRfzH4ho+j1jB1UawiAfXP3q
PjQ1Y9uH2U95Yn4GUtMU1xGVuYDtW1FngzdnO3qU2CZ7UIB/EM4F5iconni/4ieZ
pEc0c2HCoxMcqtyrYtOwCODhlhxX9dQCr0svm68tvCMsHf1t3dMwqrU4/3XbhutJ
saV/fsedf2/0s7lSvZIolqBMsGXq9GQpiC4IllDjXCmA5glrPwnH+3SG18G4roJJ
DgAq0/kH1qT5gqXWaQ13gYOefh4w6WfXzid+pKkpx95XdCTLCSS1tapmMXFl1M8D
zJOdQDrzIIUidnfW4fzOm9mGZGpend4v9MM0AMPUPd9eZnVfwg9wA/90E5Dzl9DB
Fn4GED7k97NT4BYvrCEpefDwooBGYJCeBdZrEdteBoqzmHe0v+TRVPiChEoOWDoj
g5wyiueZ5JP/9gi/n4XWnVwEiIpL456m6J2zA7Gq/b6DHK4TQgEwwg0EqFzbASTI
Cu7JyxNAr6e2xcpMuj7VCXYUip3aXWDXAkZG/MUiI+kZe1bNHSng/lavcDosm5he
9JzeO6uwWE3r9KOwC/Wr4E5vvld0LYSG4PHTr9bOouSYMvN5/Ps6aEJtL4nzCQi4
sNZI2eEoC8fuwgtHkEHG+Y9R9zhztRTjYm8gjGyfLdb4wwMDARx/+gcO8akh3FfW
yIhrb6OTZjD6v+lH27EV8Cqij/sMK3JJPbkhr3ttTfL7vzF7xM0d1NWgeTezOMv0
NxY6yX27zlnFzX2ruVdfP9W0oa7d+ZfJGPcOrcxUrZYozpGuGJZM8OdsVPslOxn1
m3HRG12Vny+TkBkKWX4DJXxyZ0KW4dZqi8/GPj3YghUI6VWyj2U4Z4ZI8IHrmklh
QGh0nL3joZbJPzg5786E7dgkwV9i2NarvrbOK4kJOxA1OqbCTtyIJQsl2QV6PD9m
UzIaNBcUh3dnFNiuUJVyQQAVJR5YSjo5Vt4EaH4n0eq4wKU4KWxx3C1vXJo2hEEf
mU8pSrIz5FO0AfFlCfEQH41abYC/eqaMHyiNJS4/Otz8lsqAoF4MHn8q8iLGvCs9
vSctp1u1ukuavlEo9UBNFBQxNrolaj32+bg3VKsHe70tMUgQCaw2Pgaxsg7VJ0yN
3qC0a7sgYtEzc1eXGq7VCf53ODYgw3R7/TjKYQdStVKJLCw0fJ+nYBm2skOvRYVC
5JpUkrVGquDNDMdwp3O0SPXORRJtjl26808bVxcrnfFOCmiBQFlbn1F1MJynajWT
QwMiNlPRR5A1Xzn+HYssaX6Gl0UZN86Nl7uTOHXgPCHZPK9qZBMoEnH9te7XhxaT
j+1voyIS2dZbq1AET1uztlICSv6gQEqrlwh11y4BA3zU3F4XviS1VJcd/4YMngj/
M2SaQdKwitKtW/Ylp70W7752nES+/BrG03t/iMAvXFK5Mkd7HdNFHtzP82pMmral
VvDu3rNsbNH5JzhH+xht+sh/q5sc/o+4TQehvouZmsQBLqPkiyEw1C4XfmwIHcBO
nl7MRI/bfjVU4i6Fj2Brnc/+Oz+OQjW2dos5L/Qyvi6X0+CYac5iLaF7B+tRWuU6
0uy/uEV9CzhRZxS20uhWXihEHBzhCL09gsAZJT00PuJlaxw4+8sUaU73RFEQ6cDy
ebMZnE/1raP6wVwTfs76Vc2TlRLUz/DRQyyS8Iou6kZ4qmAjBsVXpWlAQSSXP1sa
N7/M4JiRDSPNPIKieZ0RtJ6bWgK2zStrIhYhhZuNhxLl/yk4eZ0eJ5l0AQx8JWKX
1jb66Cc9nDROadBdrJMsqAGbjagpaVvmwoGFNPtADUVE3sjB5LdO/te8ZV1DGqna
RygNp1tK8wzdPyAXcY8aT2VzhSy4Fq+BVeFuydKzaecfCXj3YpjWDz8vrAzM4G5a
Rf87PIrddj1MjlCeanntzIHdWMr8UX9Q6biJDKb7qRQP+MAm4Dxl3O09efWvdxOQ
XPowX2zrLu6cDUxn8JuEYxo1mVcyzya/4Iqlp3vldFgYMhgv4VMp1oIpaMF3gEan
oc718aILrfgBFmC2TcLv/jjGyZ+2BkG+snVD+jCtcw6x9Tra/1sKplfXUQJrYh1F
czYC17xKA2i440RRJoSPIxZVxysfvs09d8AkC6B9C/qzM4Qp6yWYYHdd7vI6xy/p
F3nuaegNZVHb7Mk0jMK9VEe3rf4cdCiJBsMcpmYrMAJFlHJRt99fbUL9smwxORpc
PGgCXCJ4vb6mCcFky6bm4Tn5HqWYOcKa+8r6duQOv/Vo+nnmBijFHRNctKWfcYxR
1kcB778kIS2mNl+Lg9Q0lf/AK+vJimeAA0uQvMeQz25WoExOT13C2/nX5XEibMky
b8aw6aZRYTGfDEqCmqVAvrUyGRosotNzM5+bDEJi8G1vjdOZJR8BGnKOekARraWz
riNAK/huHqwM8hdDgVptUmkZ1RotmqcclEUC2mIFDoEbENQil8S79PCdwuoHCsiq
6wNyM1hJaWKm0MRUoMCXJYdgwJXEEYz+7zwbMg57hKgfCom8e6wQr2qPKub9zBMU
2lEcWIUAIhkZKfXoTq0wgxPc/RXBuUJpbff9gKkHkiqNEqqQ5Sq3Sz04es01pM7j
0321AOtJg2WxcawY2tk6kJuxNf1KcsjAbMFCj1qlpQt+R/9nGOvwMo4s8wAuQyZP
kKypxdTRqmxN+SM09AGTff12UOG+1j+J/DOumBrtCBzTEXQIBpsUu30woEeOWv6J
v/rNEcC14ZaSdzHjYCQ+HPBfLsfYIEG/peL8sbXxzpGyBpuiABnPoMwSxLm4uy+I
b+8EoymrH5abXJdhS+VWveumYIQ/L0gggUCItfRck0poyuv0Xwc5OdAM0M8WHLZe
qJGUgGIt4oNk5Bni+zG70183bAffFMqhFfDj1j+JnXAH/WrCeFvZWjocES0ztJGl
+C48ioxsR8t9YTvdr2Ll/ZSKQwcAeiHol1mcJDQcfPvOYEshscgqtcEsggmTo29J
tosjgBNpzBBwvyX/J6InO7Yi+2G19NTaUW10PkxxTyLTBaqEvaAcBLNIs/P5A7KE
8lTVU2cIaP40ru22YbLm+L13k2FhEspubpDQBtiTiTF8m65+pz99gmLhm/PQTsJr
rt2OZWDUJHXEW2Jr+n7bUJFZjbDxb28duotZv1c4nOR0nbD9aRSh005k6jJBFHRt
olK4qlzvsDQccuXF/crAWwNw3Qs0dH0tUIdfHU0TJHQyv5ATPGqmtKVJk0SeS0U/
4oQXfh0s6Gw1E1JYV8Xq8wu9mrPFRRU7yA64BYaZYqhmXDlDvys7NpDlYgKTFaz4
gUHa/6O5yIPemOt/OSs1Ik4qO09sfXd8MuQ45rYF8NqwRZlWX0eFX+xqYeH+cXZP
naMjtCi8N4UY6E4ePfo72ik5zed6eP0icqPUsnifuFi8VpUSdSy8CWODvrzxknSy
Up2Dn6j96gdNbp0K3n782ZXMwn2I1j1P5KSUw/Y+Y/q2bnD8JcLVkPKhOR0geh70
CYuUVfLT/tu6paL+fRm92W/4jrc1bEhYLuc4pW04xSjYCnnl4nV44dvg0KwkzQn3
Jh7HvPyUXL/XCocILNqnldhNwqOstetaV5mcDXu6N74ZiiyTu0u3kKML81P9iGHG
MKWL2ylAVDwPC3ZYlAtlm+sxbqk3TGKh4Zq8UP3mnOxEIw7FEVFb6bnGOq1wBXfk
UNmvZRaXXg3vOi6j0EzsBZDO7l+bkX4F+rRC9eVpPL5FCsSGQKUZr4Rj/hB2Cizw
M8hcz5799UO0VTBnkNzfdH1kkn64L5sP/LpOwOYUbZAyAZSZ4hMtAsvkgQFVTwqw
eH92YlNdwx3Av2ytA4SY1JcXzTA5+fdzRDEnwyUXUyq45JHNpAhtaqABgKNua/AG
ItH9n7GTy8h2Amswm7N/LoMtjJB6s4l7Ard7qkMX0eDYNIXwq2YxuxNjfCvtr1ac
WuXScKpbHIsHo1iQl9E5P8XN3ePQ9JGMsaVoZIa+k7zwsQj/lSFuuKLLxQzjU4F6
pZCST03ODr72uVBCqJHWlYDflW4UqgGGZ0+SgsmtlVrxB8hrmO7z2wgIPvdtHOUn
RKCXEYra1vGvPLOUmbPgmlUtjkY1Z8DOB+WTl1wPeIGZH9JCe1UZ7mbeLYwfHq82
LCi3EWMMRWJTIpl7XcrbU5cPeE5T+neMsgaTwXWelUj5YHY8YBlfBRw/Crg42aJ4
FRzGph5JZL+B9CVKM2zrI6E0Oqw2GHIwzn+KANn2SmA7so7u14sZNTjsT+zzjLuc
ifSuTqVxUzY/NHqaXi/OYv3Ijji79nWN/bCI1p1D2r1aSMe0rUtihgV/HTg87+7H
H6rsUh5YYGfpAclqIwBHMwEXv3seM4wSdKg6P7V/aCN4gUdnDErwyRiMoq/PpqKk
OaU4fLZVR/886rKS78lbSgOJkjvxJ8qMb2kdV7623hjDFWm99UBprOxPK2BZCahH
6fQ1kyZhUdmzQMshNYqNIG7/QGueW79m6Czn7BcPNvj+0AudZz+jT/ns13O35Mjz
32EmcFOfIcl91n19B1mBilg6l5OYmLKHzyXIJq0YTLsO5IJJDbsnw/iVO68veMLh
dA4BiN9wYxk6mO5MkWbdZoc3pZTaY7NOU+CE1KeuAZ/+bEq/sttrq0WsDLqlc1K4
K4LnDXcycodJiTEZq65aqtKQy5UcL20e9BqVizU21ezFO6HZDPJr15lJNAjk2VfK
A5iEDhVHknGw2KnzxAW2uEO4TYjFutoF5E/Tp9q5STx+wXb9osqLe+6H/0mBzXcU
qPiMscCHZzR5EF4Hbz8AdGWFdPd+gD0POwCKrI1FC8I8+hrONjfSt0xfy/qLNbQ0
J+wjekHK/4svOWJhIDILaTqEt/vY4CZfrS0z0+rNlSAYv84GvwqVDO0BZk5fCkIq
wxvisWkUbP9IX2jQkiDQm87Kua5UlvPwhGLt9stVcp0SpmZW8Zwxcd0ui/Z133qh
SFtI2FVUyJjILRoxXcVhTn0vC1DwzOFPwo/9BmB/K/yujsW3IS0QhUFrgEkNoEQI
VouMKUxaA55TS+OrbqUTM4OhwwWRqiT+5dDIIDSwOLv44wGGm+yTGW8Z/n+2HYXF
ZMxqUQEJC8fqT462j8T5yB4ERye2mnyunPIVeidFGDfSJTv4uBxM16wmUclvvShe
sr3eUBrv15MijUwgzL/qEX+rWsUStItKhc+JUDE9i2Ym1pq10PM41783Gg+hDg6I
KjqTjI/Oc+/0g8DhFfrm59gHGvdSDKaz5QvmJoUCKK8tDocJ4decfSKnH+qDs30Q
oyZRQkWhXhpB25VXxryU7Mydu6ddeKhrKHgE1X8FnrUbNXfSN1A7ZgDnYVOnmKIl
jRxVcYw7y9Ovm17LBtFgh1BIuLxAZUWVi5rB4HVZ9bvxECGqH7yptIdvv/cKkOjf
IDboZF+bjYZ8euk+bQDEM3mKGPz/S7aKoHMArLjFRS0eCmgwvElC6VSKA4d0x+lN
DgTYDmyz7FN2IMV0JebKbcnKa6USTbTKEh170Yw3dFHo/1uqPNYv/9DJw+wwiJlb
FKvEw4JExG0k1yy/EN/6JDo6cWaRUQobfjp5DXQXSViUStSQl0wX2vnHrHBAJPwg
euD3FYefhR5o+qAYrq0EShoXV/eAc0lLxY7hXmbj9DbLzt4rWKsRvkzrtZh5apR7
yk2JdTxXAdVIaYH0hfF5TJvnlQpy1jli4CZEwFagcP29F6NHMWzWjWZkI/vhY31Y
VRw8uh5h3gR5Bak+b2xoNPou+FPvdOyGAdOj05uHHS2k4GzDGCBDgvbIyhGb6gzO
l0vEcvJx+tk0DQUWWgY1JA2XHnSgyMAemdO0BBQH/dOmt08N5AXqDZcRBSj2w3DZ
/3ZdBLpwqkUqODhxgJ3daAJEKK2K3tbj+J+OrSaUWsGnjqbCB/QtjHNlSoDE4D5n
zREeLtWFeVnt/gryfPuY5m04140Nyc3U0r44ARz0isBsBpV5IeK7dZXqYLjlKG2C
HeInfHK47/GS5AZ48SivhKaIgWYYRXI+IxJ3MdVPAM/ZCvsYFAwo5kKrFgdciFBK
tRng83xPu9T5ymVtJUGawQJYYqyxU7sEsSmm0pOgK84AcrcCLgOORP3/xs06ktmO
EJ4KP6GZ1oh9VmauX21lG+tVhpHgzIy6TNUK8z3foq0gnR/HdZ08DsSFgSJmBG2T
tMK3ETUcTA8A/aAST83faIMyH+5XuBnepJVZ/FsS1qxwvu5JWRMvbUNQWga8uwcy
m5hAZ6stNQIpbWgzZJWBPrEqdZcgWfMp+LjQyH0oq8cVPAVyc1kRafe4ylommRw6
BgE2z8sE14QhEUiVR3JFuGmmuoFD6eIlbzIWKpIuxw3hT9uAqCS5AHAF9wtC+kE6
QRFa4z+JscwKz1FcWHiszA5l5EMl9lT5yDBGqaHL4gMOrCc2a7ZWj4D5r0D7w8SQ
TJ19lMUUFIntvtC1Z1ooZJ23lFm7bZukLyhWd8wD42s+DUDWg2fqFLMEPIIAzk3q
FL/DgxdglwsRZdwbkbnuG0UowW3hzPDoFRbyHytZzhKveAbN54Bex7bByzgtFzHP
q2xubdr8tHXYL23hdaeTtzam98v9bDnjhGPkhsfde2WbBSv/wTWsof/tkG7yJpgR
g/8DkvVzMhBxDgngD6YJFvv7RAy3h35RVb4vX7HgXDwfsqdUluiDuq2c+0D5eR8V
XcznqwedfoLA4+vuXINQXYqgk+OIAOB7d0vjvsDP8Lwx/xEU26TMrYU5ePGisJOf
1uXLK3DxoWIvJFDPFzPFfxbTLI2H3jZfqvEiI297GFKzwF2QRw7+7HRRdaaDqQNm
fJVFHQxPormKCT5EWHEWdrCTdAku7ZaEaVzWLp8W2cAoiuyCoXjGjcOtnrgYwo/+
JZc0U3CkaRevHj4AOm9nyRKEYyU7GCUQSRJWwiTEBGVQd1ZSKqfeBs4EUeO2h+Xu
eLr4hRVQ0gh9ln1p4UX2qWGTR4Ji4Ck8TkiTeI3UeUhZnCDIU/LLS+oa2S5RigOt
pCWPuEH6wznht/UFqEKAce1Rl7dKVO2jTE7CvrVICAzyBQHKM/SDtXQfasPI+k9q
TnR4JWqXn46vKogntbk5z91rhdxu/Oi82GsVU+lw7t/4+4AnUGKZw4QskPvLpM7V
ciS8kEN05ONvlUctqFQL06efq9vlRLEKpRs//2OyM8bSXuAtzGXLaZLeOBfdQVRV
SH/6mywp58Kf1zqsXiO8nTD6r9KjBLFOuQoKQXJMl6/E//PuU+/cYHZo7udX/X8h
HDDGMTaWpWEKWgY450OLN6Xgkt+Zak/rWiCVCSp827wOCWDFZSrqRX9mLKIjza1u
heSxdcUyHlAzWvlBIY+gd7Hq58zugJ5ef5CtwHiFi78t2DMaqh2+jhMTzmxvL8O5
aJ84odHZoFlNRa/UzQe40nEcHSHjK6zssPbjJFUWkVwe0X/H8RzrJDRqNkC4L5sQ
a6/CQwaL/vBSOctH1EG9/Vm80aZRXhxRMS0FmdMAX2oP9AQyXL3ZeP54v012PuKt
lltWq98q5uAlQjMIxSJgF73febdhmbzYJUJH595lx5eUOSvAlaJFlD2W16AcCYvo
FGeRsR/Mj4NdBuU5WBW4kFsOWxJ7W1dW+VCHtCAvQfTyhtzVxwQI9j85qM8DKZIa
1skeqmk9kCezh7VmhqdPASn+CJJSl+gHetYcnm43ZKqKVH6TbBKAjhXtC70fHTC7
x92NsyWvetbVIOgp5X2xHVx+3/y+2aFqPQ1GqGpcMbPHY7ckdsFBC97+ltNZhBAG
NfV0j8kpAadUIdu5EdtT16RVMtWNvljy5hRC+UXDPdS0F3d59VXpx01w21z11N7x
9JPL0QlcsMHleF2PJlfqBlktIOaW72KJpVPhR+crSmSYXR9r3sWT29x052YFLm0O
/1uL0Kgw3q+yv9aX+gxVjLT3iPFQ3M3anNoLDn4kb/af0uWpMaJmr9xl6JGePxNe
dCoxvuNbVTDQUyXuQFatpD/reE+V59c7PnRQu5q8tOCYGyQLwfAZzRwZJYBcs8NY
qYnQXDc6d5ak/vwu+bCTdxF3MF+rIctn+BekHAwfpvJ5AzyZocXPyz3ssfr4dYSw
Kb3tNvjEYcXbr7YFpiVCdKVbdRwx9Y6Z24wCbYWs3P4fOnMSB9muFHfXMRntJ5pd
hrZb/cnufE/hGplt+9BUvISRux4LYAxVAKHbVK+k0wSwkpQ0Fc9ZKoRqyx/Wdad3
Js6C3iWWi0YqzOFmJwRyc437tlfBHLPrkUslf7TBgfpBTHo2rhbJhzpe60//x0Pc
R88gfzhmUpWQ2lZWimngm9k0oeFzyp6qWnq0UMnzBt7sllXzzQmCAGJJIE1AFV/T
yx7nKtDOdlhbalYfM33PPHwhSLM53d81INh08KPdYDK7P+bJl8N5TohawQnIR5Pa
6+GV01bFIcEWRWrRODdzeATJg1uBmhptYL1IOklkTZwv6BSPpkEFjnOAdrbqb5O+
CKotP/ZUA12QeFHHEEPJKY6Vmx7gLNP70ZESWQEYuc2VlP0v5RTU9ifS/W/wQ0xQ
RHYTfOWDKVCwpkiWaw8EooS/YpJ9beet140K+NycDgWuVPfClOLh+7f/QUw9QjGH
7qst5YyRiHqmiaD8DwRKCwSpXdgjbbNptTOlvduIPaGWeJWLQW+EwMN/JFGdDYEt
3qifCCD1GLy8sxQrxkRLBE9fk39Pm2RCqPPRWptltnKKkO9eB47NPynbipIQJQ+Q
0IvWk8EUk7SQeMex5GdkpzvY5pmUQIrIWXl1W0UFwFRMzDVVL9n1W5fZQtiXJRKr
kFR4+WlCaJqXlQCXSmhn+kWz38JGNJBEDxkqbohl/8aHmDeQxMcgfoC4XYiPOE5N
r/w8dMtaOKGWOp0YmJkU20YDr/5EG3yk/SOXEoSWKX7W5bAXL9X0xUZuHtYns2KS
1+fCTBjppjl7zeEb8lCwaE2gX1l0VRbiHR++55Pz8XSjYGLfe3n1qsvespARC4Jl
3uNeDwP7FWuk6i5uQFpZ7RQ0QOIoe3a0k/3VhHDcgvP+l5G2EsCD99yhb8knwuqf
85k6mAW7hkJQpHqUn2rJceQ1GGqEwghLQVt7ehsCsFPQPl33U8zqK5gf7ytVkRnm
b6zR5t8MzwW++4yv4vzH36D+V94oDJI0WQZlbCN5BlLJ+HcQKSDfSoEzBmA9Vv4J
ewWZPys2ltc5WqOBltvNry+l0xFSR4LRlEesp+bPZn27ZxIwNl5xGLSMpeCv00RM
DagQHSSTfhrdaYNoO7QrPAEKkYPU9qII2rAx4QvisbfPrpOc9+OOMf4j7Tlw+0rc
asYC8yQrT5C+3LnO4wGcgLdUK8DMw/7h3Ox3/YAWFLmhkMhMcCxy6BFGCI9t0onv
YnC/WVgU+p+eeRhy/9CoGvyXRZCJdq77+ENksXoh3cK87iJxiVlfPbRRPO3UD/vo
kWAPoNJapnanI5RhWSj/sDn/JdmoTnkLGb8eY135rXbBdrwGESl4RAygvpVnZ7m8
j6eIjSzAE5UKb1YhWkVZf+SFrcwCAqbW6rO54QUYUopv55Gkr35rO0GH5LZBt3z7
2NMkUN+Uze69cF6T7tawRsUcqqg1cYRBLcW3yzjYgSVSh4vLoFFn3w4PIoSRhYjQ
u6CI0MpqaEtgTh26ymDHX3TT96e+47adNRob+ldhgDC6tEqwEcBvWYjGHVH8aNk0
1YA+U/F5TZ/29CO2sPy5i1j7ZI1+Gj7lHuB7S5QVHOirJKXtl3rVpkMjAFws0w3B
9ELbw1Xs6FX+lemDui8/cvEYd1rRwAylJ5pOSNovGegLQUp+qmn99H9fWR/0q/pW
bbN+eEQeYKkWG3qdGPG/nXxV1yK8CozFoWBwscO2hSFHYDUJ2CbPX6tcdfj16NWW
EoXJhF0eWCGwX0z0Pei3xCN98ZxG8DAcLRnQBbjrlv4HWqssuGd83y39KaDAbLx/
EVMGrMIg/F+pHthZb5r9JiFQLvI+KKEPqEKbdTVMqjuVLHUeqzZ1DucXZEFwr9eH
19frKbnddqSMBPwyAkB/X/WCDpCKICVC2MchOlApyij+Z/ObA+nZR2tJ8f3/iCCY
1rwNrO6EIIaDH72Y8RHN25GYAW5k2ncvGuY1Dsj8cG8wYkIJ93UCK0PkYAmxCQyp
89sNt4GojYZlvBVh7Sg991v/IQAoHFtmzKvdRm2Z8E4jR1/oWvhz+ETF2th2I3Nw
a4H6cmGJ/KyiZu5nqZRZoP5HNtES0lShv5IYQXGXrkme0A1ODeiyNvUfr25mwFDc
wcpRFxgviNW+LLHtN6/yQS2749QnG4V/OCoamKgnhCRVgO1Y4jOMEiUd8reOaobU
XYzzZJqiGX8kJ/C7mYJsEI6Y05XGY+lENCEpjGjXp5d0cnKAvXHDIjNI6OIwtxtT
/SvhUZcFpEnetvnoPLAkQr4ce2f1HN0FoRvHwigvYuVoT3+ZGNvaXZehhvLsejgP
CgZrurbPSV3upN3+ThqZ8qbsB1VAkTVN0xie+VVMEdZueg2xV1tMUs0w+jOq45NQ
lVWyk/x/LxyX4MQwNHb7zLNZR1crXRyvN/TBvCVw6YyPff8kM+JxsaVQfh/1eQ3o
qG6dx3v/RQ9fBawXGSc00J6JvGeT1uvk+cpiKMP48Ja+w7LsJJFTkGz405tm23cw
IP3wgaEcXrb94DHvW5ouooOCms3xuDgJbdOi5oIBEsVCVQ3igsmTLQ5/z53KZSB4
ITX+6Yo10WhLnHnQsi0lzpGSpWsWX9KWPPSE8oT2tbVDzVm/BXJMtj0IIk0T9uWE
1i3zG4sbyZkK3KHVfocDLeatfT0ArxHv2PW/fn4C1CXR9bZQmE6hhwRrRGtEDj1L
BYTqHaJJnS878X6Sl4vkictCXdB9p7cl2sJ2e3ZElv6I8+CNg7K977bzCrkPMdBQ
v5BgnvJwccTCmCnb1vzgu5USxFStQs2tZuLDr2sbCsDXWSR/L2l1g1m8p3RgnJNL
YHXWkB7nuxj2fnIrTxoGfmkBzsHwfmdKYu4iLGTvU3KNtue8nBNNd3dRhviND5qN
GYdOAfAKe051Camq9O/98psvwNTwQFi26TxfaCLVduTM0CVhenB2El5ZPOnYsV9m
mKZ+QTn1tdP+yLLLfx+C5gte4oZ7ZqZ20oZ+P6tDEFsI6EVxUjl53kTcxoVd9aPW
w2qAiyaFnikPYobc0+UwttGbsoE32v+pYqFal8F7eD5iDzyTzR+eYgPX6pzCPNm/
F8Rpg1geOubpaZ3wcwFK+1lyhvzM4krKUJNtEUR6E2VbLADHIZgAMeOGrwRX6232
iQh9bKU+S1g5N+dUVKMRyIDl7rEtKwe4MKiEUWi7wVlo5HY2Ad04uIor81eBckPk
+FVjc7pKWBKGV7rPwNnaHq6Z9io0ncivo0KQeo0B24K+Zqtjfh6PDVwHM6vCw7as
LvVTWoxfvu8faYs+ZskdUfF9H1hcHRwXEXlhyhTMk/dFLSE6Ddb4Z10mWahQBs2B
HuQXdRzR7xjJaeCWzMaUPsvFQBmqnF+36WmGpLvpZhNccbtwO3pmYpKU/Wzo1O+r
LZV7YST9DlCjm7cXQwQZlWBEr0/2Cz1eCbbOnZE05itcFtG6t/bEj4CQd/O23kb5
qoc9vvUkG7oPQKyqoD48lPzVAlbXhbiplWR/zk8J+q66LWjqauNGT3k+1HY1sluZ
/VtT5rFgP7byG6R46JtOBb/R7vHSe16aN7/3AeELsXg8kSScNftw6nw2YPBnUHis
M3nINMqj+ZASts2rdl0GWJoSfdu4VN6S27UZFJj5qiEIcyMohUGkIpsTwF5B8HP4
rgYUy2KzyP3CBUFvnaZLdQ4SSfswWJi2bx7JnbqmigshwVKxaWRapUfcTsRlOg22
UzLnZimNIidrjPG5Sy9vgUfDs5/p3Hgy4IhlW6gHIi6WZBRw3QNOwpdrCIFMPtQ7
FV8lj+DMu9tPE0cVbSDHg+wPkMIUvYSYlq26gCfxlTO4VqABQDNykYj6tzPBkvbk
QMoKFHFwdjgMCoQ1shRUoxHoFYYPDZWzZeG1va1XnFHHAhAgTFduxMeV98xgbCml
14NKnKWH9Bz3OYtPygrqlPKxWEGfzSLi4LONTsp3cxf0B6pR933FEm0s214z4dI2
4727ocPQOP1MGtpJsNlYZpWVbgR0KoWgAd0nRThHGTbvq+JZoWevUeOOEoAVR9Rn
r8riFknk6uIPoG2i18l6H+rB5aErOM/sOLcM51QkmGY9B0WH5YgSE7tRwMV4HOPt
yjhMmwx2WoZ/08MGCMezJLAOOEJAWbFCEjzCA3DN9hgmdgD21gj3cvYq03toZPfD
TOIidcJicGd+R9bik2h3z7Cj0/8We8qyNGrokWonI2cxznoI++3Wicx5LSKPOeGU
PuUh4SIwiqdGIHQ/ScHNdMCQb+qSybMu5Hm6evRjl44Q6ccnf5FkjGrBmqk16fqv
6O7gsO+hA6RfvvDqxY7vDA8JmPYCKln3FEYkw49+ocP1O4d2Z1TRUrpkD6QXRU1J
luJdcFUTPmsdak3vMj4MSO2QBeFzsVTq5ZzE2CyEX6Waof6dHpaeuVKfrruZGGhK
pdr/kqV8muRWN1emLlfP2cVzSFjYIjWLc7fEXsvHMyoZi4aBsS4OhqfHNW/yC3vi
8XoXQUggUMcbYE71J+SaGSxxjGjCbQcMSWVIN6ej0TRDLFfb1JPXsiWk885Po2qC
lOdVOhcUJ+TOcgt41MOnxfBfvGSx/xpV6yeI1cxTtWBTu6m/qhHOo69ewUT8OHOx
e9NxX6EAgshByI5K5whJxH13yCmiDCqnCFjY5QLKpT4/UCgcfozJFtS7fTQGHNAv
mBLbPEZh1UFcuMDNyjUUrQHhKWx7pol600DEzGKTVQuZmlhD9clKtcLhm6/dRtTG
9RjevhlzFsyx8AbKj2G/duy2h7vhYmMkhbzQt/wJBtSgh8tknORKRyy6gJFP96ox
dlannHVzGhDC91n1br/hiidK7XQOMFWx/8A8l7STNLrNCUC+fD+dPjqxVoLywGrc
4sJ3SKc30nuVcVgVpi33U7tcoT1Ei04/B4sd0LOMx4Mc9tInZotqvFb/p1OgMihN
IoBBSK6BVJZmrbCBfRfN5ACNvtEkRpUhIgvv6evHFKONqG9YZRSvFKLZcNZUbw09
1i/2BhCk0VFfH+f0/i8ATUlkCSi1VeOSq6WfCaLBQl5LRmGmmMT6LORdWYT+7qLZ
ulkDFYQlt/axT+mRZivn1c0eTCzlNEU98eUsu16qHtefzxbp1mrAfozU+Kkqw/cy
juQ3MkULKN2QY0nfTfVJfCAw7CnLQcTanytOLPUQQ4fz6IX/ndpo0IizBjSUgW/t
k6Q6UV+bNyaBGcLbogHdpt8+h5svsmuEwA9GdEd0VZppxU/EqpllipY+0QuJiGvr
EkGTAqexHIuZ7xX8uUTCBa0P72VaLyjT+dpegQECtfd0TdmzfHE60c9Oesx6jfg6
FtwHYuBHyi1mugxElw/dgOOg2AENgiAnWipTPl1AwHEsvq8fpUZTZoYLyshXWBVI
mo6jeU3XHoDwxiL/nWFxLFyJLgui6PIvNwabJkaZ8EMdW9SXYKfdRaPwQJrcOjve
l6zeamxr1oapZBHqOAxgyHauprnXeXwciOPNIdlaJW6aXvtWIXHo8VEug5Thc6Tz
1Z0A26A0tIjzbITEGJUUU1PqoD9R6r7bYvD8iV1uUxJNAFKzxoSWTErNIN3+TkO+
waBDgsheiHipuOD5F7edH/qLmNIr21zRcNVE/Dig6yTIZDAdG+5eDl5X5KG/JwRp
YCSy7HP528+Xru8nrGnSgt8Obj84z7vZlpny6YmeoGKkCRgunrMQ7Yk4IKeAScM7
OtNcY67wc10I58xcTAXdo61w8x02SKT3lzsAa/A1qDOQnzV0Wb34NPXP0sIqra0w
5o8XJvnsol+1p1+c8hBTZHeE92/sZf8cvtgFCyOjv0C9Ija+RmdUw1zp2FTILppz
3gp+4islPFOR+YRGex5x2GU3nDC/rWHI4lf5zA6AtBjKun4n+SS3rvj1POPHDSsp
FVLbX7k2ngYt7MxL5oZa0VRjcCc6MhXQu3qHP1J9lHTV3S3WtYBHFn46hsELP1dr
dQQhIdFHIApGBLSAdZBZ/oBNfmulOKjuxyjqNrq21rM8IAA0GC4VyydyLvDMcaYa
rBXqOf2IvGDW32g4Ie0macUB+PFFk+OUsIun/EVH0Dfr4ZgiquK6HMLtYLBQ/GkI
1xV8l0u3Bn0rWdVC1SYe6HmOe+GAK+p+0ZAlUFBl1vEwtNRjc4ajNaEgRvOlpceG
krY9mrQfJGLNX9rmBsQbkDSh69wlJxwB96SKzQcoSUlTUprYKpAugphfS9m/38CP
2d7ZNfTGgVkcWwe2bao6oXISwBzsMeUkrRETCZefqUUY/aZ3I1JMNb41j5o09k6Z
+c5hgZTLoOCP0l1wraQ7y8tTJQbaYtSez2vnNYMA7ZcqENh2JXWtJVuMdNUoHfwI
u0AY4Q3Fo6vZapEB+/1sPGg1r/3WLGEZJHhJPxUQHYGaXiEGuP+ez8wpW5buQinz
oWrhm3qEjrWvN0MoKlQvTil0572zq+VDI1fkqzj++22ribyeeL+5Cs5yUMzKGu7/
ZrJqi2cBOFd5bF+nL7IKEiYuRzk2vMedl9ae2nP9moIbCLfCvNm2TwrUgjhim2OV
TPkuHrBsWfUoogHk42jFgOYYTjwgTDy2rH4rocau33jCDb7N76x6UbtWCEq9ZUQI
QFJeiUsd30DScXZA7wCEi1+X9I8grX/pEA00tZtg2rrTC2uN9V2Qhv5OuaU61KUM
B+wEDu4F76ASXtQ+LggbgQ5K56t0/OygMEDhJTYjAvVizfBbVduifYs/0EIkHHhL
srSXZ21YW1iU6UkII0R6PDXuIl/eqeuGUSkZDR2Qn0qA+1JXj3ZPR1gAayXEiqus
GGfKWWYZy9MD3srCUMTxjSisxoFXe7/QcUiikfCm2bXhOswqYl6ZRNXP638kOSaw
SjYHAbqsHpS/LU/v7IWatEV1wRYAbNFK1RKKgig/q1kMyG7M10/2TZZVqDcY0XlW
fIyNOU62M3vqOOFp7LK78yURpHtU7dJWn47Yk9W9gPrQfW9njSZHbXgTIEhgx/p0
ePhQmJkMvC1A1xr9Asvp/meRVpV9AmNfmVEvbk4XOQfpCDet+fA8lFYdza9vu+oF
cREGxvoJxbr1lzP+JZpCQd2WVREAFqX67xWuB6YL8Fr7s3ZaaYQ2pu91QfdVyzXT
hkwygYEHt+ACFVRN/STbCCioNNPx+h9KOzk6pmlePykc7//qZS+JTC7S9sucZ+FG
x9cf/OLnsW4ItgpPFWowj4ot+uF38CjT3qUfO+jtVHtJdQNrQJbAuJATYOWrBBEO
1U6UJORlt7Am6F491u+QhmpEwiEpzmOw+b/s41KTBppHPsCaWrqI9Kk37vULylfk
X1IhTCb1Zc+TCKuXtOLQq4EGJ8B9rJ7AfMswWJQ8UqKAZqgBVGoHiruVkDtLJhPY
VI2E/Fl4X89EIVnm3hBltqyZR8otpLGXshAU1fCnqy9JtzjRpSMBNdZsdKX2iU0E
8LKcfSsh2MBr/uAGgtJ17ZFaGZteaoQvlcqP/HDo68bNdF36g+gEWiguiFxkU7mb
uE8Qq919b7OPtbT40OD4z3mWKTk7dFUu6Khv7LL9Uiu5wtS13yx9Bx+J9fybdrr1
fYyJgJZjTNW1p/TYX7cb6SCC+sRNZgWajsk074uUJiaCYmQnjMwPdDzQ7jqyJRFn
D7Kw2GaTbTx0aoSbNs8EssF7WpJcHd/BMA7NVpTmC6iuEm7cNd0LkC/MqMj846j4
Z6/WFT6fH3eeXC5HgwYZymDWE0iIZCbA1xTzEXOYtq9fKwgLq1V1hKaG3JjmUbDX
KBmzbY+pXFQRZvp2dXkN09gCB19LwTHoyy/n1PP/KH+IPqBrrRzk9lHvwZ5AmF7w
G9/cKu/CEISOscMV44JSMkha3z75TFC5GTIIfOImonfBJnmAwTPZMlmNI6Rp0jvy
SjmetwF9HRKn5tLlDLCcSo/NJAE81E1kRzZ6zQbQxcQINMIKlKS9pxA8eXLZ4tD/
jMxXAQMYdIJ7CpuN6ux3CFzfe4xz9GlcOZuTLJepyalVKkAGNaJ2KuQYBiVAFrVy
fSxfSfu3Mf+BFAKZPO8ZAh7Eb11o25Ufp58ag7h15UzuYWysHWazx5YKK+gmoYvK
UeiEoajQvSvTqtMbC1pHLBWJv3bIVlPEZ4o5IGZOynN/7j76eVw7fdxDlRMLuhW4
yNHqKuaX2NuSWcJ1SrkIYNsEAC4osCt8XmXAM/TTIp+QR8nNoRcGE4xCKrYdc1V9
ux0Nw7ebqmU6s66CZINb8Z/aQ+y7Fz4hufSRs+bLAu64F1ksxTwDXmaH/ogABykp
1byv8Gg0qBjfEn4YkPKqVIXX75m7Y7AsTaKdK159Wyrx87cjML9EvzuUfDSy3UV4
0Kqpl0nxEVXuVjLnWSNwYl8lkcHWK+hkpphyKlfslGmyTFWbZ8CfoDsbLUnsmvRF
gMM1PFuEanA+34dKfdzXlxfcDcNgmjUCDOhzME0wAsBHtc9lZyD3UeHUSqF8OrPf
5lbb6AgLv4ftmp1R2aoN110kbL1Z6w5VeAgasFW6yE9/dKqcHHLuPSct5IzSOyjp
RZK+m9x9WVY4i5Akzn418FHzUlTIj+zHweXd03Qf6TkJTMUUKo/vn5E+/pA7MH+O
VW71xWDS4ZS4c8d//FG61JSHVjKTGu2pP1gpuQ1x7YquafU7JlRT9KLu0Scs1DoH
rDF5H1P39m9kRbf+wbk2OlLgPvDu95BxUDlRlUgwb6Je9vWcY+NGhFp1EtpKenoy
ADt9AV+t1Jn9bv87ktrvbH0c9ykUgQwr5yIZNTVuXpMOAcvrrUxKI5z8zXYWtgpv
bcnCVI3Vw4hztkTxmGoUUrJMgDWdBDIvVr1xj3MF9T0DTNEhDmP4SZQ4QA5JuDhg
R7+COYH5wTkeAosX2Hba9+8xaE7aKLFIJEw1fQogcOKIi/ZusqBCaVtH/Uxttf5C
NuYo5pOnzVQQF7zDuUnW96ofMhZw6bx+iAmBoO1J+CuV/5esCbsrFeDR7wBaDJQH
nyk0aZy687IuyhcBbtAYagHgStv9KjC6EA29YEfZTz/A7iYU8S7kujUPlGxs8arL
ndwgbU1OsZ/yP+TGRUvsRqM+XlZnlRYvWj62kjBG3Nx2oS4QukiRq1FgoXamJ7Pn
PM7qMTYNbUdevX5MJIaSgETxek6Txr3i+n9VqeoSsxJOQWcLux/l+LQba360DxBP
x+BDdXRziTnJBoBwMxkoauTouih2H+vR4eGiIXS2Zote58PwA4rl2HobWRtNxlZJ
arGiytkw7vHfigJTtyGSVxQ9ABsSreQAXvn1CU9Vz+FDpakFPIo8qmYUcf/gQ8Xw
li1IFQLcZnihOfzop/wyQc2iYhU8X7AaFh2TxJmlzp2qFUpkvkkIdH0JPD/KI2bp
K4N/lQzeSo9cqMMur6ik8qvt3SqqUbO3Q8QJGlWeI35lFUI4bi05jiidBsf0RB6L
ge2soiXtlp8jByFa1qhq7rngZXoncU9F769mOVJpvAWOV7D4p2DUd6f4og8THOKC
Fcn3YHBDNF6IOZWG3gNmRIBh7saHCjCicACONuiVQoZr87AlZJGAQY0FZm/ttiya
hF/59Rs0N9/CEMYs5gk+NORzVtQeq9u+q+ee2xb8LSSGXzmamfxtNUDLLJ+hEbDo
QeJzkqC/wwTotZzGMP5ZndRsETgMHz1HeWv1aEI9H6X9NpcaH8uKdU7INwApD9AV
MMJCIlVX9uQHkLQtrTRpOtAce4vxeganFVUJaoLIym5nSxByVbrG3IyLhlxW+yDo
hFGdklM1X5Y8BOgiKXtzON8zn8OYWTPkXvLfKEkTBm17IYCTqG6EFXObMzpdA37Z
hVhJ1coJKZ1QbHb9Sv+9xq6yRRf8LSzvLsNkRZ5scj6OqjxCuTyWvUIbJ7rlQ0l5
0oGxVktdNeGQrwR4nYNnx68ebGZCAhhhAE3kbXaXHbQvwx7+MlHkmNWsBH8qG3b3
Bd22oc6C/9BXFxokrPZqU/WSH0tjQD8f0DCheydvBVZm+RyKufuerpIxm2XlsW1r
IB1da8uQ043eiVikUJHMOYqaw8Nuwg3GlTZelMm7Iqu05Y3IQTgmXxgrJBA35SNX
IHqW3AedvNxqLFL0uZl1PuUDbp8AGyyaOJuLgew8H+Hs5L+OBRLGjpfHQhmKkVqo
8SUf+4I1CSzVc6ZcN0kYf2ZId4BggyreyqP6z5viynng3ixB1GmvVrGSU9vQiav0
d+jpWijdAoR5OsrJZmbf80xJufjoay822PXgDj8jxLXGOLRN53nrGjOwAc0fauc0
hcmaZRknS8oLlDQrLH+XlGvBiaB60ackC5cOTxjISQjKed9fwoc1dflJVHXxhaDN
xj6RpT7EL4DrUVNCtrGk1zTguicBWrhvrnfQsE4UcKHoVPngJyfX+4GbEbIGduOa
7iEpzVuQV70L5xlzfn9w3PihWtlyYJEpzp36sjNYAroq2PadN2nmn7eOsCiKeeMp
7oIQQWDPbUqytb3DYAe858NjVsuwK8na8cn0mDZYsnWqwnHxLnlMm/17m9Z53drR
JxfOkHJqyN7EMjtyW0QyuG5nPHS0TB7Fwlg/mVcd3+0bFEEesUmPX3BpXCUV0dQi
L50QBg6MbRNT/3uz49LXpTDJB9p5PVm6AWvR/pStw2A4LU7+EOg1Fb/6z1pa9bdH
PbDiOjt97Af9dhU5cUvVrESjx0U577Lr4oISRp0KxDiapVjLU2w07SCi834vB8xb
3SUCQbvD+iV19H5y2Lq0HJEhEQrKP5rKSYZxtgS802TmYua5Zdl8RMMwS44fBjuY
IIkRIbSzaQTorRR3+NUHXt070NL2JdQXz9atyBpcWXsWrxmYnd189Fi3+BSInSnQ
nJ7hCX7f8oJteJK1iZWPhj8XTUqIWVbXfO9dXrTroD1bQ6jp127oymDe2FtQtVay
XBgSGTBnLpOl+eCmWV0lIffiVU5AFUXPuzd0YAWakkvsgaUxsB5yRCaZe+Pjvgbm
Ik4FBLpSbSHotB9esgxrHLtalyDB6iI/XBUBOSYmvAuB3+ZgYtei4A3LKCLFbtNC
KyWtRh9QBIduBAdiYZiRrmcceb3P0kRxVpD6bHSkzYRgFzwI6HRoGM1H2TycNYWA
Bhe0+78OzmxxKdhsg3CpJ4aKjRMUE4wxGY30ua9uoDVSvQapkUFjkG+p35L8LETa
XqfC1Tdu+IzPd5DAKdzJK30PaYQA/U9k1V0FTpB8JfWkzfPzatGyCwQhOxJBUMiC
gdfTOY5J6h6bfPaXiBwQpMqjV8vEi+oHJHW/LrGkJJang5D4FSc6zxv6zz2+H+ry
GioA/fHSRZPSq3+eZWKmeVcyJmEwwh2cnbRY/C0oNulak+QdLYuQGvhd7oEa3QRW
oAI2S7niJ1HwChRE91jIb4DKYRzlc2GEeLK9/BLtIuG6+hrqsIK0xXel+iJidanJ
gP5gDgee6Not461r73iwpkXScByXiYEAL4PMfifOZ215O22FrMPS+pl+bCL626ob
T3UDn73Ei/w/V2dBmim+C7wvMlm2Hrg+vIv1+klJuXHPM7EuoOIld+1S/NyN1cVb
3H6CTbb+TbYgXkX65OCBS+Iusxqajc5cZAF3B5I1wgmGLVEPtGNSMaaUCzh9LGhL
5KRm3dm1pawTGR67aEGU8Ynchh3qE7TMNBX4fcat7gTvzt46lDqmw/EsNs4UzMwo
RTTyAuGRJAiesr6MLU8WcKWrCSgQ8X2MiBRvs60bKiqayTT5PORhizfklmdn6iQp
llSVqZuSFWettof1jK6ejVLcYUvcUukzlT1NiL8ivq2EtaszkUsj3sxiuWXU9YRg
UuORZnzcQcpEcTi7xU9m7nmm9p4trNQOxBa0wPNNFH/uRPpqs9kQSXZFxB5R6VyG
72z4fIUjCNxFgwGOLunhiD5EzN52i8BJTZoRSsl08SXquJRRg8tUwF+jRTBice3M
7tmZ5DHFky8Vym6LDvw1gtTpwDdEGFFU+QyXlBMRofAmUmsf6xgVxt0Oqi/phqQM
uA0hmiSudDzCCY2QU0wynhelFBSiiPWqpVyv+7Td8LaBD22HN6siDNE5f1Nnjgg3
beJZst+EeQceq8I7mJTcqrmGHVWMqfJflAZdoy2h+pMLSpDtfCtm0pFFTXKhxfdI
xwkaRny9O2ltkweVcygRUZ0Zke0KQ5fmJmTo/b9DtLGgtgcRwPf3GcVrBkMQ0wif
/oysZZo6Wudwh7bCbo80herrmyj7GIFDkXukjFUsIfu+06VwK1YnMjodYKhweoiI
V03WXxaYSutAVDPoWo2frETaSrqF/aEvox876kD0AzYz9hi3uw/2Cr7WMkzDiHH8
dEzEmf/KmG7W08Zsa7VVy1zB+01x58QUey7SoWrLBC5S9YHA8oJ7SWB/t7XwoQnL
mTmBNlU8v1CSQXZlyxa/jvw+i/X4K1HrX/caPYxx2uGYUWlTJMItacJndkJzjVxA
zFJ78dayu/EsJmgLXCXyNrYW6BSAsDeBTaHkrx4nlit+z7dYSfQGu5PPlqSVKcDJ
kCROsVPn8m3NwWMAVFZSk1/sp98PrGHZMgWPHV+S8K0AoXzvxos+/MTPuVyXSOYv
hgHKLHk0gePRHXoTy9n3LW+b5o0lWxT+Ym5gHrpTf4qcWMdHBH0yYMWBa8y6CXfA
U91+7T1X5e70EBF0tJkbmY5y4RBwS4S+vXenhQTawtcbfGphwnf1y8FhqzScmwpo
m1hFnnJumKwBGgppLNYS2DIQVL/mNtM07hWd0gThovczGtxE6Zcc07hPowf84UGw
J/HX049QsRWJt28Nw77IGk+7CZRymYXk9HLegdKhMpUmcR5CrJ/zRJeQ5ONEZ4aQ
pObTLAQpOmWfBy2jZRMQk/syNxzIaKA9K7uJiOXdLbXf1QUQ9B1FcSfzsP9635ox
WjmNnQreBUd+x8/vDU8R1zaEUWnv/tNOoONMpFcqkBijb9DjM+CC3EFcD8UhLEFN
lQESz2nwob41N/deMK2hayhvVmkNgzvX7uO2iTNke6mNq3PIxpmudymBup8B9GVE
QPkAKHKRPrtJY7eXWLms9dF/GCXqTiOugMq2EO4TsgkaeRZVgGxiNT0e2dRkPlm5
L/g5bWjFop6SNhiuc9UUKpxv7VAyYRR3iVNRbpygQQFZTb4pJuqVc4FUlCCP527N
7Wlzyy2gEYvjm0DJfq7oAlWPFFaeNcnrDgc8T5WyM/DBDWOH5uRGyjJrrhh0UT7m
IJ0EINRZIeIJ8BHvFqrYYdbgR7YqnxII0PqfXp/QP+eWiMukKhJEp+L2OAf8R+yH
KSZiLPxSWGMF+qufZmj8SGO7ev3UvB8rL1/x6mjiwy5TaPwFdUWEKzW+zJcnOhAY
ntzrm4SGLFbpLN2zdcezkGQGMxRz3kBMMCu1stkfOdIAciGngxQKm/Y1/b0SQ1BN
hVBq4ogdw6yRlmhuFpzE/FYaiCPY0Y8dVIC+yyeU+AuvfcOgBqy6fNXIyvIReRgl
zKqmWjFgxnrXAST3yEelM9gQJTOKbHwtGHUejrdB4QfGPQpCktNqtaON5hX4FMSq
K/Mr0gmeEYFBBZxxZnPtwvvt+j0MgqmMrtL6z3ncIyJl/cwrZOctPI7BSYJYgFZt
6WAni+P7xShWLFBDcVhQiesnT8laMN2xG5CINcHJ39ynrVW3beyn6fSPjx0JttnD
Cw9tBuoB9x4ob8D2gPj0CgwRFH0N4zGBFFceKRBBRqIC8wXXvDkgU11AFr4bzYMp
zdIO/xdr08e8qUrrc9Ps4u5MmUuRKR0PoMBk2cESdwhAwE7pDGxGla6Y5E06FUTP
G22WACNa45mLa7lhsz8W4rjyPmz+Ua/AEm+zoednBJ0rr7s/jfBlU+rDjmNvZxK+
IP1ZJUMEh8srw2UV4FV67oz4Q0W05Yo1GFqkt29Q+b0+1kWIVOWrR7SD7uU+4FY+
g6OWnGmSaWSP8MDe/GoThr0iAv4AwHCAw3bNIA8nPbdo5ZgWZMgIbu/qwmNZvhK1
fJdTOiGHB/J8PTsEol/f98GuWIOkQm+95qVaXB3yXKq/xaOPYhSSM81AVjyYdEva
lIgY8IcoIwswBBi256sMJacL4y4Xm/fwsCjoovM2QIihdQPXf9ZufxlC+L+fHL8x
gBAJyhPeAvOkDC1HjjYId3WneFMB/oraLiRqi8YAVOtiXGVOsAY4OZlyYDcSffDM
iAzfFSXJc9f52n2KhsfK4L6u8jiL2YWI2+J8iqTJMP55mnXJTumF1j5mZxif2cKU
6wfki/lpnXtZmxF91c8HE6I+45aFy2hE0biQyXmDXlljOCAVAShALD7aRIEozRpW
IfxuMHnzsiWdJAHZ50WY10Q9tV7ptkluu8zwuhqz/hx/mPLt/l8KvXjUVVWP2VdP
WSPOg/0aovNojSam65tEduPyMDkyaHZ4ESwXyNfddZ6KfVL7e7y4QjMbeBm7lUdN
AuFUO2dn6VZU3nYMDWy6MTjBv+kUp8z262nmvtv6mdi9BvNP7Nt4L94QKiyE5ZUI
6sFoniN9+p6+SAgkz3rTad2Zoz194lfLLZUvvMbEShO9Zb14IQUTRQy5CN1XtpJt
80ZIrAwuiiZCz426WB4CpY+jWwBrsAY61j/W0UtEgQAliHBKriKbEmgJkGDx3lQH
SNPRSZOFMF0h1kiUdCwWt6ODQqik+xSJjX1Z7sxSEnSl8egHAhTSiQ4EsId34Tsk
265BNPfjGEkps9BA7Vz+j3ANtnb2TZUPqkBLlDJFo0eFdervcjPtAfKu4uAk55Hk
cPRJX72Bh5RGzAENG3Z4mGsSrOBe20SrDKtWRk43wHqrCFn8LkVPRzliPf7NYOdU
9QZcZ0LPiR/XGV9uLWW50cfcA2nkj6twPVDP5J/f5Oku2DJICWIwIoJj8aKTVB1m
J9zY0G39XEF/7s1LIrl5OlXQU7hKFGjSIW3emeK7WrEmjCFkMEhqiGigpHbY6Icf
do8qCjgI4wB7vLfz7x7bpTbh9GfDXsJTbUHR5JBiAknBYN5J6ZDW//w/LVATzZRc
EBGfKqwA1BAW7FHPB3tSrQjY90ACBrmA7R/gjn9XDpRolhZXOPy1y7w/9qM/rv3v
7PtXnBxTi3M+38qhCDUUw2hQCCg+lNTIzW2nvvE7fjrJ05bXQP8OOTa+gq23svaN
vGEWA4HJosBLmY4H+ClcAG/fxX0gt3gGzmeT9AS+66+ImnYwrJkNENPO3WqMwZPt
M1XmKBUw+fr0aEcUQOMlzBLQg/kS3kr79To8OJOmiOupKZM/PUWqA73PaoVjun4l
qMNrllkxynrpmmDkaBEs6sF/Qp7P9MmFZL3P+Scbrtv+2zy0KjiofRhqkCfhaWiN
HR4tdw4kUlMxI6wLCQj/KJDGKj2/K/CiyLwLKXXt99YRK6g+RacmaFDn0J7heX7t
MWwcZyu2tSFWU6osRuUPzTsoKhMQpITSNsEcRaJ06BQ9EsvSAZyHtoswMesq27RD
PhUE3xHJ/yFHwAsXhMTkCo3OXrswjsRxDIDe3rpPyJN/7gktgTrkBIAUSEHJUofg
Pbe1vonEmwT0HCWK6tf719/bTA5Wavw0QbEKXRlUhNV4hDK0kpLiQEb5z11DcWrK
tJgYdHIRdwjHehgsQWzxNu3BWZhlHx1bje0HQpV8/R3lsHZNytOyAIG+S5/h33LZ
qcRRo3PRd0ChzB163bCbJtibcKCaM02z8GjNYLCbEs6hg7PGS1VtKvUhL8OP0iL7
nFk6+xlZPQJPMStuv7Fx7Qb61nzwsupwEXdy3f9pqhn5E0cbmgspczORpdxbmJME
UckPJ3KdOM8NqoG7LLLnSxRrrWXvo3t/rELiF5WNKrIGehVdq6zRLMF2MWJT432c
NC6wdF+XNBYD9gg9okLaIZKAiTWt8OAnWNyQhPCeFertr8EmU6fniayzUKc1+s2a
bc0Ajcmz/1B2QfBFG0i317TOxJDmA+dLBrPi0NJBeOjxEYjlofPT+qmo7SsDlBi2
uj52jGHMgl4YW0w8kozqv4ORH2Hw8Gg3db4lxyjlWSZ4kupsof6awU2dWloKtxEY
RDWH5+yWX+Odsf5kFA81Cz4ABO6uWVhjDk+9q38TJsOPFZ9H58aLofoKHBjamtci
hzYmRDcAUrdjUWOeutMlIEccqXQHfJT9iZggSxRFN98F4igSFZBVThyduh7agNIp
Cz/9YaHjgWtCC5pYbCqIPJe8p8IX4HNJqC9mAhhXJMlAE5TJjNc93CGsmklmj7IY
9ffAXRCsgay7HhlCYfL1E4xvxoQ7E1OQitOlJ+s7bTSH1IOr9ZC0Zy6CSo+2epp8
JvcDeDK0sqIODSmz1OCUpWUneWShSwXia57CvBVNxEy6eohAlww5y86EBlKEldCI
Pzowkjxi5H1pNfl104y/b3Zm28T8A9ot8eC9J2ARx0YivdAj7K/ScwYylnzOOR3P
MTbOcavYWElq+/+2C6+UIYdzsuAMfQDlRAhdflBLFTN0Tcng43w+i0FExDiRo+XF
GlJdOMd31EcYfHzimSi+C/xpZRU6JEPOdbhxulacAiw8B1osG48ApgxllK4K1UOM
A7CsfWeS6V+gL9eWSP2pzP3SYgO/MfE2z0PrysiqqHrq+q3PTIEhzUwLcOVerC+L
c6C1BvgjDXpzOFM2u62U0VofTJy0jDei89QSlCGdV5P7JWiurboehxEEnzRMRpoz
mXiSrGm+CuQ2fau2udN+Pzf4QzkFnTki40asH0WlrL59qSoasqEPRwDgAj21Kptt
ln0WZxKHkBebWGKR1WYVFfDvGFUd+q+iqSyTQWFRgDgtP4mYHUQ/qeTIU5p2XgH2
yR7VdqqPj1e/9QZNtcCd7/FA8v82LRs3sLezkIXXgt0ZF5Cx6MryS3dYgzBNvtQi
AiviKMuIvo/ohuqzUnpbno8bxLea1+31FTZrAYwmMZUfsmD1XAkNxyzBAaWtWnq+
stSPc0Jo9xPjeEJoNMd7/pwzuODjwTWuL66r06isgGOwNuRsyi2QzW2nkDlewR0n
LiKrd6i1pXxEzCYKxskMI7FaBVyzSyj3x6k7fLI/5JPYoJtILNee1tBx6Iu9EeMc
pRkjhvgwOtHqH0rpTZ2KGzxq3TEGVLlDO3BFLfTmUApkMtaTeCKR0z72l886B15I
RM8pJXNuMNQCnMrlWcZfEb40x2KPQZNrfofOU+LYmi0ElOPplsIooQvvVX6UvhB6
iBlqmoulpdEOYaSKeI4uXlR2FN7OoiezwKK3wAtCJYPBGPn+xAtNvndFZs3sZ89j
nRiv87QvHp/xD9m/K7YvFQu/LEeCTIBSl7HZmTUooPOOD1gx486+nCo0wgPN806F
q7Njn33STSLncQ3sV7D+W4Izm5P4E3PpFA9CjBe21uPMl82aeIjXNQKaLu9JUN0B
2NEMECZ8jHjeJWWtgGC2Jxjdw51zZErU7sbx9hBpv1bPcyUuXHaX3Soal+ooMaHG
ydIjGJPUluQZJDZNzBS21SX0AfbPlUjN6xl3yhUumkWNnYXHkKVHqpD9Y2JeoRAE
PjoSr0MDYQjR4mY9GkC/UaEK5mkAtA3NFlqv+aoQWjlTofkzEw7tMWStyOcEOn2Y
mhGKjHiFBhDraXnj5f9Bpjw2Qa4pVppGkZdoWaki5vJv7Fbj3dUQpCkJZbi3VVaf
R420/GcjDzelm1/f6t0WYGMo1kolUH6aRrM4sp7UUVTLDrYIKFxde7vyJv/p6pYv
zaYlbDuzArwg73jnxFnvi9kSugnczqZVgQY/oKjE9cVuQdu5hEd7vTMdQTsXIUak
o6OkJFUiVt2pFm1ILz5RfHjG2KmGZotPOkGRxuufEIA3tYZTksg5QWenCyrC+a8/
INHcWmB0J5rYCO8xtQqzZhRaWnPwfovGlnq7ASpk2YGLckjab2CnkIBL0cS0EECM
TXWgUQk4OOa+3YSOJRq88FmouqnP4FimvIIrm1LhBAKoAiyWamdm0AAxmi/LFDxi
ajQr01ojBTq6M2d+45EQK3QryLqUMlUpPQetAMH8tS4P/K3GL5+qMGhTkvsrH5w/
WMmBS6nWCmqNq1B6s8q8u+AyrDbeHRhuCPyi5X6DmuIMdObg6JXoZiOBX3m5/Var
U1NguO1TGL89o6vRT/umQX+YbznMd3U0CyB2fdKHiFLTxmXY50bbuIDNkk9/+462
p3tQAxIqZX4E5HgFovBAmRcw6RryYgYtEPSaJAR1tsf6lKEVBmMyxKnTJjAa/Ftp
M91PXNF6sdWh8xv+O9APu+6oB/hvUrVcROYyctMBaL5NkrS8Hwody+WgqOm6knO0
T+pIg7eXbyFuWnyjG6fOIscqMOQE9kwixdCjHQeWVQAPIIutSHox4H5AlGmyh44S
8kHDHMbBBNTnFtc6J7dTLLsYQz6rKeoslbFZpFhNKrJyBA2iXr5XHQswMZ8YM8yp
Tn4yhdPs22FfrWiFTmkBpiJXefSDKYGR7yy0rwlYhpl+pNn/n7lRGQZ1kGbFG331
yUYp1lCvPKhVgrkQZEKIkSYryozHBgSbblIRbEUYTY7h0Fmi2zOrQpKAZPHF9ZKl
SslfODQqcLAKCEsiglbYpop/0wWVWqL+w/3gpfC95/PN3HJ7FVgcfm6SBT8J7ent
y3t8mwg6q6FjHDvFE4vjhwRqmFz3YMMMD5wqCtUt8DHLjwld/VDqLLasIF+nPgln
9Zh8/pvu/0CMAeCRLsMSMiUZ1OPvo8m2JCFCs3hvjAKDjHrNiTy8pTZAm4fh33bV
CZjFwtvUqDp3mp4qFyh1WBV/qQxyccC4UapKRmhXROvU+rlkAvGVLdjD43hmWEQr
zMhhkGeZNbYarC2esipdblOsLA87VgfIl2NAYMvsccJuD9fkNsRLPbnIDFg3mYde
7ECV+Oej7+wAdncfFOKvkFZQGFepFNTxsHwnDPjuZ+t3kmtUt7128dxw2DGFUFmQ
e3Fx8+6US6j2rAY6m9ai2CSfLLoxW26OO34XdyYhno421+up/tBxNhGYlou0UwVa
dUvPa/FV0AptCmk9QpuyazpUSDbHbu1csi8mKnIwZsNjsifFGnsFPlj11HSlH1Gi
DhlS7REz063CUi9PtXwJBR77omq+3WTtP1iQ4lvsSmBJ0lmHlq/BVRn7KqIj+DtA
XZq0rAI7Hv6/sL0vbjrjS7UH2esT0JT7kUny9YjuKMS3EpFqgOd8BGvnbsNFdmmA
GaNsRrdAv2AnxdTd4AeQ9pInarH7ttD+m1qV+qOyofWBFrvS+IG6b/OeJy85xNlo
FhSnGpO8BF2euCyCMzu0gKKUoXyl/j2Qb4rkZ0nkfXCd4hMeOiWwI6UR1qD76lic
nmLDPApqw7WiucI1uWkrRy2BpTyIrJddvdCZJY+NdIv0l/HIHlUctZ5IGk22kOM9
4Rohq1sdusmygl4CMhXy39kbfgWdB/SfbKOmbDZOZFhrcPkTI053DBdBCOk7eiah
nulp7YpnKiewxL7MZNKAP8L312AoedjG3Joi9VLTZGqwcVom7rgnxResLF1eYmAb
rTs06Le/Hdq2ukPRNeJR0N/sl0EbVsHG9uHre2WRJEtmVeP2oeIL4Do09UF8CVsK
E4fir2Ht5oeKhGOF/xSNlEv0JeKeIK6FbKxRPezrAe53m778qsjqO6EInkDeBNrq
jWm50YtxL1tqHqNxa07KE1oPi4KaRlUI48IiG0zj0fcIyB1nCb+RaeuuQagf/a/T
xvzqXs9Y1mb+TlCapws9MNVioGlQ0hDNDndQN+ESqbBctqp59YUUQhkGM7Pq+j9E
vJSds/HwHSiBHS0f/Zu1a6U841fl80sZ3vjrxXghR3DkcN/KyQ7vRVtQJTBcyjRL
as/FOLP0HfLmASURih3fCYg46PsFbCJbaVHwn5EeHIcX+KRdWe62IoqxV68qTkYe
vo0VryMRd9bAKQfnZk30HJ1gez+m4ge6mWYIsSOW5ItaNg+0/UrZMJ+4EsPQ0RjI
6AlMdVKJTM0Pz3ZFDjL7zvid0oEo9TtFlahRqCHZh4jXPygyJPQJgmJWPo/WyL43
poqGGVxpHHJvk42QVfW/kxNFzlp426p3UcK6zTU4EOcd/ZzqVB+t8i5dHozDl6WI
IUtrZkVQcnkbvgOXbxeXYvrtayVLkKeB9IszIMmTT9of/RFMYZ9ayCv/psXutbiF
qo+0Uhha6eKoyuMOssop1+XbqyKDkk5Xt8iOCarKQbKU7wstIqEbkXsvlOcPjql0
m0tpfe9rve59oVx1c0MsuJyMc+UNCnb7dSLHu70bIvdkS6sYsaTnyxXGoq8Yk0Ak
Ju7BfvxbU+AhFyBtfI3JU58C8VaHclEChibgDai+j8Mu/ohNc6k59F5s4lwxFJmQ
7qAAoFc8/ENSXEj041PVrHw7Vdh5jbd78Pvuj5Qvgl27/cwGqnUIMDbSWPiBVCyf
mYiaxX+LmgoR5LFoU2vmEz/ZAZiLZuY7ER5VnNzObX2FkXBW31vXNqCCBXzjYqNC
YvTl+y9gDPAJWyWlEB26EsUfct+DxxYF3INXIiF2LqUkXr7xtKzUxepWAGbXCc0h
j/t94iG2s9sstO1MEBpdDNeGzRtY8OLG9ZfXAVbfX1iYVWGISinjPzJbuCZLhqii
rKtzThCKve8Ftt0E/QjMb1Y19bv6CY4RIKjJrLdzL3jEcE2VqwBYFXGzUqrWIUWV
9pT6/qDAunlsLNC3imHe4+9OeN+ARaGkWQzIIXTFPuHtdSV7e+ePxexRctLmeHsp
ZFtVgRyq8xnmFFzzPKs24DVbhr/rW1YdWBqsUgJ+UPKNa99JC8oHSi8ah43AQz9L
dmvADg7lMpJXGLiDg9+r47R/mG0aHld5uWwWX6pHRlTtOGoLLQRqHhed21qty906
9jlzqSx2F5m7g2PB8h42cG6DQd/lu+2MzIdHTlbDLBTiG9oEGKgE+gztWFKDdunG
K086tfC8h3aMA01g4TkgbAguPhf/50AWXlsSy/ih3uj1SAeE4tlMTGJl94qftW1v
HOUwwkedl759OtX4/ZRYvZTV1IsrRKC8+iaLQcsjfik5KCLQKemhyP92kAnvyCuo
ysSY2abFi8XpxWR6yuNjE88+Vcm19zuS8R84QRgRQWkjTtfSQe/HJSFJUdtEA83g
XcezWq9fXaD74FiWtqeH+Uud8XlxXl/5UEvBaq+uBOFUN3nVSqhs0xP6TJF5DoRZ
QEGj2bWq6/30DI+YsFK7k0OqsmegmYsUvzxMsd1CIbUGRitAeuqWQyrefC5j9zPl
AdWtZzzKkzxC3ZfeMD7kEgoJLsLG3AZVnArmDJo9vWZ1cjUWeic8zZKFIygkArbW
zvnz/9T+dBVuBKUwD/2CZXeWjj/ZtxSG8hoeoz63g99Yi0/FLeW2kEFLNQPHe/rQ
mcfutfjXWEPfM4t2ArfC7DSZBSv2QZZWoY5+UTesqNU56qJozqm5Jtvf7pzyniGY
64N4/6XJAhq+iBccm0g9ZioRuevg2H8veQ7ELS2lLMJjv1x6Jm9vTg6pehRXZ5ft
dWnzSQ329c65VxjK/KXfFt4QRmbgAvSwik8cEfPwRI3Q1VBezlqJtaaoRFYknwJK
JenybD9mUFIbBydNZbZSTsYaubHwrorC1Dpljnq5u/UL5+cHTJtAG5hNBKvmUwYg
RUiETpSDJMkaoZYW3d2A2mNiYgTK/V6ktU9EUPhtbfbX16MnNWPLOAkVtmOgEulm
8gQ4TL/M0zRGxaiQshrlEL622dOaUtv1LEP8GiTW5L/8290yroUq/bMYb4bUyAws
09wOdD6UaBqK/X0ZU6k//rrlkgq6gcEwiVVwjfAla4XZZtTOf/Q2T3PzynAEvf/9
pwG/Lz5xlfjLKntW/h0VZgwbwWgwnAZfBiXE/eiycxDo05zRyH/uU6YBurTfRcok
5kZ5KBX6TXjUpiYoLc1gBCxcrDR213O9DAyCFz8j4cCSJVEo2u4kgKXOxNgIhTJH
W4fFGPFQvFxZZyF0koy4DCYIixp/rKQQaucmIjJqvozR9Pr4oKzwBzHk3GHIdsxi
t03MonfzVHg3wCzilvBN4DQrTON9B1IIaVbYyIforfUTDuv6BCZIoVETPhaMyNQM
sNP6qKou70b0bzxfdMtb77WbFFNQqFEBEvzWsY5k92tT1YEdNUmG9TxS1CViVvC0
AXHX+HCrebRPKrMIePdx5hW/Y87Ojg8i5mTFZb58PsO0DVDvHQ3onhb/ophxQEhG
6YV4CwSo/kiZJ20UBT/lRwWjCVGdN5E0WaWufMe0LthOShVh0IiYRoGQ+ffKT+Ru
qXe3JCdmS9HPBZ7LXpMK7/njJOccHpXFpdsS9XkHcagsw+bnwLIW+TCSnf5mbfS8
Spnk04LLIuF/Il5HHopDrm2hJWUO48IHIVLDR9thQzZSu9SUKDGQH2UCQD+RL7KW
qATAkTUiA93sOIJBsd866UpNnKnY5nLp5fTR/VhA7dosQRmMKl77X6fQYh7oorKt
7fzcLLG5sYaUq5+f3c618wdBCPFHg9qCpSchhyN2Gv8+3CntLKwDNIyTUF69smVt
mwShLiCPAVwjCNE14U6wVodBM1N5ILCI/DtZiCKb0GNNvkltujoFfOd5fvHNuYdD
Wp9t1NPcAWLu1mW4XQbUYZ2juKDy84x5Z5REkZFD5STEwNKDuzfSoisy0XES4rxm
fPec1lw+Y8Ul0+jUJBGTxWsL0QQlc1kJk/z8ZQAdbehll8vZUH+0b6ugJqUvMPbX
qDyF76WYqDzSkLEv0K/8pYfgD4VOj3gYTCqcNlbJZjNJGgzWwSsbpOYMcw+mXkko
pBteOSxWh1p/z/H/b3vFj+seNbGQaZ0/xY4LzeW2WMw68PUWrt1AcF6Y470YkfhF
o7iuLebnMW+nOkW4HVAqMpUCzM1dLZeUyKIRiXGM6BZptrGV8ut0GRs4ASevAEPe
iwOURgRU3NDFeDoqKOHTyct3yYFICdsB9/q8J1/oZrXhVbuaWTZp5MPmXu7M4Ijg
CEiTfGDL0b0YTFKS1jmw/r6Vt7Yfj6/c7rT5/wIVsAn7n/9Rq4FDw+k67PfqfSmy
9zCkRn6AEJ7Ro3DXgzycVxNjlrdnsqq8xkT1K3tYbgFHjjgbbev58NcD8H/UrRA4
J1JNZAdxTfafiyn1dLktdKVcG+KpkkRZxTqPBqUf7plr1PENGPkeiJMc4m3TT1CB
2g1G6ppY3o0L7I5ew/ylce9Zmyucn4sKBP62F6bRCe8JhobazBJaIE3TjDHKSyqg
UtzIItn+zfouzDUFv+HQ9MpBD/HG3EsClGZomVq24cd0NNPzYDny1BYnSiFc/pkW
UpW9Cg3+IwtgSNFO4D1uIH3/Z58BjPY2GS0JsBJica6h7WelE7h18to0tm7Oi48r
BdOafVIkrXT1qjX4c4rDuhZl6ykK+mY5RleUZBWxHggPosBF4XsMScBOJjhw8cxc
odYEsF8ut0tRm9R16qQVYsu4DHzor+vv/IdOoTUtYgegHyFNJgcD1l4QJG3GkGqi
D+KXOXYV4hVQ0xcZKXNlkJcW6YN4CRYbGZxeeGuon6DV6R7Z/P/qUAG29prh9T4N
K7fU8Q8xmx2HvEbrW9n07EBPvBgBXtOBbMgVojo6ON3r2q44cct2Gk76L1xpcpQ9
XQf9LgjQXlrzl1bvFhIWxQKcRWcSbI75nKzjoO7rEINBSut3lHGrh694ZN3m7/W5
gLxr/ETHClY5jOxMuY34lCDmCYNXerqCY3iC6ZX+B2JVIxd3QtctigugvDbe4lBW
XxbVwddyMxUTlTKSpBYE4Lux/MSscxh1+5a7sa8ZhgsKyp3ME8SLTtYQVnElbyMv
9Bw+mwIunV8b5NJMfh+/tjBu7TS8gLVn0c4PIY+gKEo38jtpNIgZ8Ar87RnDw4gw
OdAtN1SCzW8zkbaNGgMfQXj26FsSvD1BOsVVRDDgjgcqWF8YkjPxsMSMkHURh4Ue
DE4qNbeHCxNpBtRDJVSPbiQFdBcspKZxf02lIcSSQJZhSSzlVPIxUFdNvQW3MmI9
RTTuzuJS9VJq8PY0L4vEkzZwmu8xsQ74sw0d1pAUEpOvISvmGFcCCdrsW8VTAfAk
2cDgyNxEJjt1s3bs0a2c9Q/OnPHiI+pNQK4OQjkFFDUv0f0s5hDw1YUT36A1EtT7
vdRD9a+Dzs+gukvzy1AqBVSXUZaNhFRrrKoCxmaGfpdz/vsrRcHIYIs8OtKyuJq4
xpHGB1H5ymC1RUfOiJWM93gClWXGhGQ278EemyolGigVCvQsaW5hcJRFi8t7+FVg
8q94WlWGU0b8jyKoK5bz7jb8/NsUllIDLO65iHymn6cIzwt4b/KTRkimF6qP3AF4
tLJmF9Am8prqG31XgrwGrbUuYGyVX09ikW/SNwyDt874yR4K6KaXU4u7fNMOkOx/
oQePw+4JZRXj3TOVnEQVtgWowAUU+VNTG50beecDKzRqWiWlWUQnyyVfCQ1dl8og
5cjxo3LTwAVaMKTbq4oui/uqme5IEhzG4/l5YD0dPaNOUzBGlF6/pP/GbCWJetfo
FJjShFFntXDPbHTKWqydw0vv2hvFNnO1jM6T3ec/ORHeSF78c4jBFOp9bpTc69tR
UVR7PNdFRlqGn3X2NtsHx3IPMNESu5gUi0A3+krJDOns9g0QejK6GsJhafX9rnEj
k2U+cfV7glmi6ehSw4IO4gA1lbsT22PgsIcTG55m4ou0zCQonf1AktWLRpzNPUSo
J0IS/f0qww3D/Uxsv0lCW86QDFIO2V+CpoQi1K45Lom9+PcyO/T/405+Xfng6+/S
rugaDT4m5v9v9hAjFSkq4nU+QQ9nuLITFItg91QrQfgmsabxWbD3Re5DeIPl6YCl
pBLJxVdEBidvbhqE5YmyZULx/IgQlMzrTLGvoscexllzi3ey5TnbP1B/Kt+W5oNl
l4Bf7ntaNhu6BoL6FRhm41V/Cr/1s7QNPFAm3Y4fYWUjTdj17imQiDwCrahL4Idt
t1+kpq/KI1yo3keQhUcotPz7cYu+UuI4de/8pNRShkIEFaaCEs9pIhKLtP7Zqqyu
Vi4F+3yIKfNFeKyLuPig2E6CIUnTkwCoBLhGVgZtjotlMoFq+Cgk6sOT/XV5M3Lo
I47ovYxEwuDDvYrC6ilv6Z8MAsatu3XgdtDqeN0wTpt/rmYVm2xPvgp6KmWBAvnZ
iVymNomzF6E/4H1FBSI6M0VmhPgqR8ZAZGwJmGyg7DrItJHJR9Zi/zl2GDwMfeag
Iy9eddnPiL6fgvuMD9bJ7+Izth0MEG6V3YaYhARxT0Js5SEABwBz2ghARI6feVpE
KLGAKKUlfLxflJE/Bukq6XufTXqLUigIoJf9XA133bPj/FjIZdVRFuq9p8aqMBS3
wZoEarbtUwZG8rWCND0GLG9lG9W/WVdGGikzJiQnmjhxQb9CR2jGPSj/HHlBtfjr
eoNzBUKeKbOPJwK6jmvel2JMoDMuBtVk+4+tiOLuFQdvSMSWUYxBIoMLNMSmCHCw
Kd7qSgPb+mgsZg5k/i02I8zA0n4SfGaGpxdgCH0tiNZW8zDRxhHwk01YWvFptUnS
Ly/GKNptlzkotyU9B1jwa1ErWegYs1dOkox8R7vAS22RqTuFn2CSYNDjlRT+T6ec
ymes0BQ6PZPUpLElIbYNR41mtfxNhzxoU6vlxA+T3oeoOiHO76n6aZB0+kxTNgaf
OB1lF6AdMtBvVPf97/hyZr4OTBWUZCi6sy+QZIPDCBkMDlpii7a3kMaY7e2+2M9V
QRwY1xQFfVo07cabIn1sZaDN4WfWObejyEMfpmEiOsi9unhlhluizZmjqoCpaZdv
Ypocc7B0v6iu+F5PabqexULHaGUlIx8Aaj4HQETUfV3mG6759/e0xz59iYiWloyi
Rq690Yplus6rX87EK2fh7RNEzdK+TKeAxyWFJ2Lpb/hZ+wR2TFZUWgktvXODSWLx
ysF6SechDWRUYtzDhu0wK9lTz9WppG01d/eKxhA1dOpI7vGxFtNPQcLE6nMGlFyy
MNn6kzMNjf4pRpzs9E8l5jSwsQberwy/WcU0UX49RKCTzSTiN2rmtgzcQVD/4CHU
YpxBu5/I4k004v0nQE/NZAfeGgemhGFSE3aJ4dP5JPyPMVNtxCrjiQS2Agxs4n9N
FEu6aXWRaAcfpKu33uLbJjUVm/doeHww8/2zY+M5UmhKtIdsANkzK6IdixUjA0OB
nlxON6f/EDXd8aLg0J0ZOBWfV61lYgMjFbNxSjSf126+l60oOniTx4Y0exBAYv8+
fDj2FF9+sxhVybTxyRxCKq6Tf7/3gXoAl6NWwh8eUFS2Xz+Fa7hpiIotG36EfZci
xSXDLTIUvjCblT9iVxuTLHpHowL9f5PgP8jO9sQzF1whlT50G+ECHONv41XdjEpI
Ju6PdHIP2NvCLL8WF3LOmqzYE7RLk9z4DWDAmVhW62V/CD694ScFt0kJu0TxKK5j
/osollKvcjswQkY7goE3POSxG3M48NJ5hPf69WTGJJDqp57Wmlsxp/PTgzhZawGi
7OLxTI2WgvEO43u0xVUbexlEu2kpV75mY0DdOlzL32bD6OXw1BeWdOS/7d+jO1Uc
pVzxHpd1Rq2wOisSjwz0xbvNq935hzTeRh18pgsqdI/jAA1MCsNaldFeIKg1hBpl
Rl7lzWHfbjaX7j8+sFFFfRmDd0puNE4d+9tOgyJkaKAKF4Sza22QBVRwQ7rOS0j8
pR9BLFqYljXBgNN+4O05Kguxn8joIlf0cVlI+CkY/A4zAaYuC9mJa5zcwrHQPENd
dk864/BXSC4nCZF8nIclpjgLbzhWIU30sPjZMAs+1DTidFanxA4oNHTBNJA3ZN3w
RI+lSAPhdey4mF7AQaEMehXzblWIB2Xip/UcVHxIsKM/Q26n+eYsKjmdvv1vE/1m
0qkYSZ4Sgihgr+nUelgidFoKs6ZxVgiLdmn9QIspqu0NYfEF21qafwonH6cQ8nB0
l7ZsqrrhjFgu3Ww3+d9BW8a2w97pKa8qbj074eJWJIJ1Hr6rWop2VWnLcFBxQw8A
60nxbK+oviwxd4nzTaEUW8zuJEdNUip3PBF71DmqA2NLdSMCBeJFko6zihFnGaAW
GFAf7cyQsMLzqyt9fa7BbwIDYes5TGiO97jG/pCi5J0pNeaUGmUoKLt45xGH4wsM
p22oAJ/l9/tAIQ42JDjC3cbotMj2rVR4B2vqU0tc0mDl2DdLwNgvn9Zt+OE03POH
0M/U/HhuZjP71c9Aoy9cL8xbJStatTN88d1cpNHyY6jb4xFJd1w+xOMG4sub7SvR
+rerHUytAX1dMtXujZ2QyWQE2RAGRDMB10tPH390Mky6p2TV9b1nLIDGuBT4geh6
a1B4WXOddYMkYU2sQFoWTvUmDQivnPEpwhAuzUIu0sozDuVci5PoGcS+I3ZILX0U
pvF5H1Wa1gvrFmpPlhdj8hVzp74VuuCGSI/XmpLP/Og0YgTOBIqe5pqRzs+GdlAi
Iqghz2e+T5WW4w14aWuVlUxSIka87kd4TctnOAE8oq8X0oSpXlkcokfsFTQYsSO6
Z9KUmJslYq5M+2YgWC/GFH2fzrq7rxnRfkizCIP9l8rQiWgxYGNxnPilm4SgC6ls
rS4r9ITVSD3VW+3DNZQUgJJfoTg9tFojxuQhLL5fWCeNX6V9uY0YFXczkc5xsCQP
i7Ji7dYHDKuHxBlMdmJwLpr7kTYdLWY81TY7Iba+FrJ7fmep/Bf223dtHWFCarRD
2CHjlf+PLiLgDC2+wH4Qll+xsODZfExtmC5G4Om+p0lC76eDYRnklLQ6E26p0tU4
OVe9LgVp56H2nXdWw1r/vXKcrJrp7mwMyZRhVMuEAkbG5RYmlONMF7t8LMeKkHGh
H1pTFyUnqmGsjn229ZXNLZuLKbU1cV3Z1+CuTXPLaZX+i8AJi9IWwcLLV/0fTzOk
RbeZGo6e+RQr75uNByoQHNqBfnZ+LIojG9x4hBENgNNv2Or2bETzwbOJlv5EtC8O
HXdAt9ffk4+xz/lpUL+xSftdJ5p9Fm7qCPjL1je1BE4rs8deODQMAhJ0ZadMvUJt
R4tTwe+VKS8SibWAhTks9MjPJnrDv2N0865ZvRxiJD+5CfkDhqVSqNau+xjU7Tcf
FUMQTRY09iw15BfRirC3RBkr/iokFA69XZtJeQkuSss62OVgN10Q5j0y/SXiwUDZ
khKpfCYMAcp6S0h4sF7Hcgd3QSNR0iO0zw7ONwyZffCPmGMh4DjGfT7yqRESr+Ft
+Vsy+/Cxyg8S0+l+jXAbOv5SQ/Q98n/Ji/I3XBXmMJcBFBPOWgcUoRMjCHgXq4wL
aAubVDqRPGntD2Ck0Wp+1et6+sn3tmnk/Im+hM2FjSwfqOhltXB6xHesc/p/UsKu
GRqs/HfK3gzlNgutrrnEMpBGtMuNn8gnLSXY0o2XzRIkFjUEz3jAZdLCjz4bf6T7
Ua0Ye+NuA0/Ps8aoJVAMRdqBFBqf6yYagqmXLsz8UMDC41T6+dBbgREGh9ivU8a+
ukUqCQZv20vQQ0DlgvtEgnbRssoHOH2qrbPmwy4E3SYjonuWEMuOKrvG7bygDaX5
z7QBxLUebAas4CS/sqDgaExWuz3j3UeCPjV1esOR7lHTz5mqEMMF+9fl7y00hSro
LE/JF1T114k8k2FdmJiMwcNLYlqrMrJM2RlIxd5URaVhdqvXhxDWTKw8CrerNPW2
sjtc9lzlrW1FbJCm8OdrPPLnSTpXeqnQFjOmBP8u+D2Y9mJPvuQtoT4VU+bkZK40
0JqX2T5CAWZc8y2V8qeZLcpuZtaKovZfVcS1MJwRwkLLCX+iBZUwtbgYRNQj8Sty
PPjIWQ1zXG8qL8JtA83GZ2hxBMj/iMolgRe7Uur5um3vJw5u0exzWTRjMtEp2Mvl
m9QiE3SmAFt8zdFMVVyqdBUuJT03u1aRYWdlyKhKoV9PX4ncc4THpURGfwwHSnvD
kujBvdj8HiyvPpC5gJbz5/Zq5Hl7BSbJTpPzv39M/6Ib+Z0CBgZo6KHb9zJNWgBa
Xa6ro/Df6Dcpv5trLEzGvlqxAxuOpMeCfYojDl3IezW3dd4zSlk5C9ry7P1SO7wJ
IjWuVcC4bfMXGS9yUY0V5HCLo3bJnIxrsHV2CIL8wxvBZ5mlb40yBE/MRN2J+Oh3
8PZ6O0PkIe/70GKF4XpmwFChUmS1WnPbdx48aJahWN2vtaYycyL6KJ0X2gGDQOD5
VznseEqPU2Xf2zapj20FIHEiWhSUwwC+uhYJFji2njyW5SI/fNEMg7gvo61HlfBZ
Aw4ars54IPLo2kRzeNPPNIGhsT/NJxxwD1h28Wj9g4TVoc+kWOeY9BO+FgNV8dA7
yizk09Qaq+HlFx7+HM0Kwli7k0sE0eyOKCMLQ9LCdr3efP6aLweC73hsAlbM1yg1
Yat2shyuKi6DBsS2WSksKd4atB+tSKKSVleI7MCbiAiCwnMhL5vkfezS00wX2EE4
52xrA4E598qf4nldr/0Oiivc0/yhaXeIw+CqIz0duwn0uH2nbkq5pB/ABGBtqd3x
r5X+dRcRPh5679fXQrF0N4irwUr7GKCAJRJeSy4CMNonDGs6XsBpxKwIVC5PWK+s
lLUcATOL30PNd2jrB1d/98mXbNuItFrEx6E81Dfc1cbFY+x3xDF7OaouW6h0ERdY
uuka1NHlFHzk2xV2qYuoYePA14qrCCTQbjW3Hznsb4QTqa4cPpmc9aoZcDrnkUAa
LoLs9uYxiKADrQnRXNtd6JehM8JAo96YXcglhgitGzZefwf8OqbnPOrAKOGv/oKU
+E5rIRzM3BzQiFfHG+LnFtqO3hjK68VR8QeH1RTuLgzZDATg8ZXuOyXFMk4Q+bbm
/lg8RrtDD7QYuRfvqUUi1v17Qsjit8V6OoFwffk8+J5JaZ5hWCETFcofcYagI0E2
/ichpMcVU6qCHl31ETFmXL7IO9VB54doYyGORCgKVsCxnoxV4kQUYRd7FAXdtMQY
W5k3EiEx5NFt9v/bAzRvi4l7VeUsMf/bpC9+1/GOORG7F3KtPefr7VHbZHcQwMG0
kDKnAQgQoofObLSo7n4YZBB7RXZDmfGa5n4ittJZ2vC4Xl9bVrZMAXUxYIc6Fvij
Q2w2Ygpc1X9Ry0D+uapHT+XyrmI1ADrSctXmSf9M2QQJ2sctBzRNf5Si/ZepoFKh
hs4Y12j243X7LUuT0vdvoS/IyMf/ylsp0NWQxVV4Xxk06KtN5I3lsy1bFNDfc47K
1kC7oIO5LjAKhsigXWH0oXRDacV8QzrApTWJvyIEtJY7/9Lk3ptOrylsulCKHR3E
L5UJ6u20DrFF2JlmeDPwlMxsIKQnQyz/NSH6BwNg7cZjl8kK6A0YzTryfv7jXij3
ZYYOiNr1R02FpOyKOwBrnLS4EztGzjJ+rWTHtJVUKAvehXalh7QIZwNKAyvUxzml
X0nTps116ccmzWCxfkhQJPfDEJmpH112E5nlQtAKkwRcwxSHqq0kW4MrXEuioEGF
toB17Tioh/VNTPsq4DPXdcb2+M8FI8i7pUp5SY6nVlFXjsrBHJ4+3GjuiZQpa50+
Ggzo6MpcZlIBdrRXjG1QIUyTKyJBz1EF0aSFeouBY11i7J2irJ9q/KrmfxeuRvEl
N6EgtH84diDk8Enj3EjlNQOF8rnoB01no9e2TTgHl7teAmXfXoxBBT1UITHDM7Ow
fEWJXf+Rq+C3g+8ghHWX4BIWCe06wgoLmleecuO/8U2r5eJIAxvz60KSnzmU1wy2
RcHeP5OeN+foomWbR0CbxuREb653ZcWqAuMTmtCWSiPsqzmRDk8XysiveqdsAzl0
mQDxB4gWQpDugu3Gv1syMER1m4FgLmDBn+/dJtv2uPuXsTFIcqA0vGC84l0VIlXQ
g5/6ETWIr+wVCctxSTncWM7JRc8nVM2lS++94gjc7D3LA7sr5vqghjrte1OO2Dyi
3SrZL+axZGluVtn/HMGhyE4btmSf4l49zpBBSronPci2j4L2EKnSTdUkWpfxsLIz
WssnWBz9WJ2rJ3Od9t5BNj/FdG010mWmZRSJNFNoHQebGj4u2aE0vcOtKR1D0LJd
MFIki6Ya/OiFamOtVeqrRjZwKenUYTvZTSUXPt3pFW0KUcio/cEOt3q39W53DgWS
7hrhUyjudyYa4CT+ehIa7XqBrzGlIeTjRJ1kU41jgj8eWawtG0HaTYzFTGVe9xTI
uHKe7GgkHUjyGdiO1HRvmbL7W9UPv7plZuF1/Ywl7jgyM8VZlBvTUEWPuvAOifuu
Nl0Qnu3zHZn/CAGT7Lt2e6ooDtqf80oL7UDBBiS6Ig5QsxJQGtArgWMDPrnXMRdD
ncALD3y8AiW+/Jt/i+KGKC1MT/XAkHqDMahlIhGcAVzKRTZRuSRIuLaIbhKNKbrO
jzBZB0YieLVunGZfynCCeVfg9k5qwgiQGoX/KuKAl/3dYWkbN2Xc8tD7iLcNcNkR
Ho6zlKvwGCcd7iE7SUb4+tYjOQXA411DrOaEzhcmSBt/17k6lmtQYQWfu+KDCtJc
d5nXq7612jluwst45jmbZr/YHBYioonHXKJC5GsibESRnqIyCj2/IRaT6FVUjrKZ
VLIwlU6Y0f/X3jAqmPuZgXXXT+4vEYbrvXJPcdVriEwB88AHzZB/VW2kLyMWgdPi
WJbGkP8SlkJVD5Tf5FxzzEEjdlV4mpa2h9Q47b2PRDhO/oP7w2pUA+45p3kstnMt
7E82Xy/u8SNr0UiFjTzpVRp9BBto+/ZBMUcYaUL77Bd7/NlNUcN94i57QHP7IlON
qDiB9AjwEd/NkjFVb6Hbu2VXUzrvhnIKfstbFg1WBTb3IG/nrLyeZZCdIw5sdnLb
9WKptWxrAwHdxBEqGJgLQUvHRY0IaACrR41Jj1no5w4XbHYLVzdOqNHlRwHtDlJK
+JLbUMD33O3GcKMvMz0ggNs2wftPCJqCBFjJNQhNZpchjebBsitOPpoiYaIB65oT
yzeNrvrDMz5N4RGMQJZ2l0dB8pfrXAa/CQROIyl+csrKIdf8WffdOWk4/GhBHwwy
arRX27S2pPIBC+k8ah/TY1D9HhJ4aB+xLnp5SCYL2DKcOQ9a2IelcMOZJMW8SUg4
8vpxo8eLNU1750tS3Beyc548xQOEwoIAchMaqEvJGEcSQ11ZTXzvzWJlebqxtDzR
5UChHx31j+k0gmm++ds7Dm9BbGqIPVBVeyqQERIX6Xr1dCpTL1kYmKKESlgmlIU+
uvghoEUzz4pcSu802N786/FqFYlSDbx2eAX6nXY4XRc2n0fqoOegng2ZOVVyfosJ
FKlofEydfb4ip/v5huJMbBKsVhJ/fIHeoo5pZ5r3KC5SCCdqtA+T4yK1RQFW2Zxn
JgsKjY0ojnp29dxeJXp2mt4WoDxVFbXnHVQ8y70eEqF8vhjHALln/Aaawy+mxZno
wV6hmhi7q7ZjKSkogClMGHk4Lq8kUaYi3ZQ3ZmhyCFHtjFEwyNt9yZVMsJ9tfxEA
WNyKzkQgWvNlsZw/g060ohhHTjjFbEm9u/rESzKK3NAnxEN1UUMYguyUVpo4/Zp/
CN614buKRIPcnlPLP36scEb8lFXYgWCmSaQvotg4mgQPzBr220JBdkUr778bZZ6O
nZ/pFYkCD1oS4nmr3kc3aXrs/EbRfFIINnOJqT9Rdu4eKpy7VV4o0qmo4pBal/yA
xjJ1a3ZdP4P8dLYO7ZK23q8UleJi3vCpe8V0gdJiblhMhcmlvN2diS6/R7VsUTxM
WWWfKqVNsDF0ryPNJJbQp08CI/aeo66qG4kvhjZ3rsExbABscb+2p88oM4H4yHmU
0hhNOGf/9KZ8MFWUl8FtdiryP25Y4rlx4hvVVx7sNrV9/OSFAdc0enXxebYsb4RP
1TDaAWQsJ6QVjRf/NwhWwIadCLJ/OBgM9KNl87jECZ0JtdMS59BmmMoicQgxXiMt
V1MmIOBKVKZWKlu5p+T8r9RkZgJ/FTmKbsWJfNY/jWjjn2ur9uJeQOgy4xYYusLT
JMKV9GfsA9VhYIFclNlofJMscLhh3ouAiYzJoiYIsJ1GryZl+oznoY9tWogkDzpx
2ZiozxxBmXT9EZEp7XknPx0Y/a8pSQxYNTj0J623rL3peCd1/Tn1v8zJHNVS59V5
ijZ0jf5DIMBs4Rzfko95qDTVSLuy/VgRMX1h874f51vN+OaKilxsA01yehXN00Fb
tnUAv4DDVXsWViOwUhADG86JzN237wz1LtIjmq2ACQbRzBPouLZDDMKQ4mYsJLRM
S7qvvQcixpRepkXPtMJ7tQIY+rww/zKTm/rfQ0LYEWTqwu9i9ktYLtPcsbLMXtF3
FplsjOrr4umzaPILbe6it9EtfZ8Fqg4iDXjljloHvuTOTnRJ6uvRaeg6yR8jB+0B
IG+umJTScGkF0A4pO1mRqbosYn/sqri8Ef3oB4rGLnBLZr0V1BZqZ+gnc+6UsGhB
v9NFlLBM3p5867T4Ji+vHROADD0izjqEHRVWy9qn8dWVERAwHERgtLvlMVrJsl13
iMnpAAmx9wCqCvU17clqk9LTTgsZi4NNiXRcs3O7twbvsTCdSFhO9OtG3rd6DUuZ
I24SrZXxRqrv8xCDaD9BZlhS8Dfrnip4TaaAFRUHjmxJfRDaNwHR8jAoQWiYUy/3
pDq63YbC68P4J90B1+7Jb8qwzdla1T8LvR0foMqJfh8ayIkGgUSG/VPyeJB+XYWb
HuKxsgOWxrLG3gL1UJmIe8DrK5Mh9/iZOok45m1VAynsILC+RVogbbQ2EvtsLejQ
F/BzZGs7Udexmb1IVAmX3CsEtNhkhxDZZPo3cs1vqdkNCyVDZGUMM9AFfWMp2kbW
VrP4aOC4bN8TzgZIir596LoN/ltt1W3qqVUu2bwMFitMKbixyme5RSagvMsgrFhH
zKyFMCxCjZSu2FbelZmcok4Z/JTWcS4PsDb+9j4cZsYNSuLuxwq7fNbOkeNcubJd
UUbiq5DeWqx20BSQHKX5qbPPD0T9T9XnNyGeOQ/bJsY96Ml8hUjUmTwRDBixZI5a
aQYiqGYbmNLK5e0O+dcVvrLQleAn0fQrx4HEzzwt6EX5+hzu6h5NhzQFZM7gOkgB
mgXeOdpWUJ1DppAxcRyQynsSeSUHx0njcrvzNJLw8e7vfLiiY4vXrWijoocZUtqu
w5A5N68jbpgjrwJRt2PzsK6afQCe8TyhzUHW/N8TGCdjt8A8yNXgbKgliJV9ZdRq
HNuZCrzfUKPbAeWQrkKT5asj3acE47Y5lCFHiBH94fJuFJs5PVf7MwIjdrk7z/Ha
XBfDQjekQpR5Dn1EH/wCafihmLs8+uaFKkJp8UqeAZijjxfI3dT9xgahHjKdDAUE
lHm1B3RHGUf7MiOKxSk7wDwxQ61D9CoQeBVdiNjC3i2rmh4PbM1aivQhWZtAL8yr
iT0Wl9PEyep5ZtUOPNdZvuEQ/BhZoZq2RrruEhivJMak5YWw9c46QnHJVQVzPXZR
2jNuBwGV+JxaUJ551/Pui430ohciZnJVCtndOjKkKjBpTK9rZZnQcnokxLv9TzKX
tTpGt3WNdgyWUPmNNI5JdYQrjdDXsbrb4jlQb9+JCl48n5oU4p1u2f0IiHC/xMdo
00v2gZReJ+S0NuNfFqwujnhF1sA9L/gBIISaEFQPcerijhkiiAbPvnsIP7qpzhW+
3kN4dW0DbY+oVtJbQSICxjE4m1LabtDYzzVRanZQROheRmZmGK4NsGQksAOon6OZ
SCTf77C5mPWC0YE9c1dQNuWPQ+VefEWDxsm5M6HQQ1mB9sH03vQrCyZVc/97mh/p
S5lFQcw1+qtTkTVHRRJzu64s+5D+CLNCBHoay5L/pKcTpoitdtp8+GwUXM/NjaNy
EILfe4hPnCgj18dKQBOH54e+DqCgBN9D/uc1cH1cUMN363oPUj417FYAVuo9uDfn
otAdY2u326XOux8aa70u/Vp5lvWL9HPKIrhADN+vAVu3suad+eubcdASok6pFtBz
S74hw7Nn3X4G9lOI+QnD5Wlyyl4Hb+9nC8K9nmI6riCsjYmTUcUhsaVwKJMaKYR3
KhRSq8qYZ+aB3sCC5fp9ymL+eCQjXyI4shb1BW0buBMma9Hyt+t5rNNu956UqTng
7df8ypi2Otr5Dby9tLg++61/b4fk2/Y9+2+zT0ifZEeVL2sLPymQcyQvKB/bx2za
XSkpcZYWlIg7hYDx6o6/6lvGin8SbqhRPNzhV1pXHg4wKKGO3YIMQxk/dtKVgzNm
TuX2towgqQ+Q1VFbVKN+G3GiG4RHli2IxLG4I1P5RztnU4dmG1VSH1unjNQz7oxp
hrChbnmtETt58ks8RGLnmt5fy7PaSvaE9NOT8gH2rHp5XdfpwRM0p9rWhhSF5po1
ibypBTCx65HK+GmknWQphrBZKnxQOkk5fLaUQwxY2otL0gqA5ARrdAozsrNeRAgj
h4iG4sg202skKbD1Z+UHpcH+/HBItptdsGLsWUGZIOzX1heUSM1yLInur4C/y3FP
cvgra+61Owx3myOyIGTB1mFaDeIh+glPS7/wlcVQIggTQxrQrpGkIWwqka2ogV40
pTyG5MmHFI0bJ1/TwPKHx9tSQp/W4J1BqejpObXSfCOg9CLLkBZd4jJEXY+hrsQG
8v5N9+xX6VxZB67mkMIwKLCmSggZNswI8ZzyCmcLGD7keCkBdJZA6RaiSc6O1aqY
wNyNKGQEinjZj6X1bnyzlds7xalt5NtzXrTu2tXXF87c/ISJTJActxq7moLis5v/
u3finHMoG1B9AOxYLc9Yo9G2hNTwPmTJqxvaNwFoYyocI0989nyaWiHFjxTqvV6J
NZrj2gtTGHYmD27iGtQLmCVfBUHgwBTBq3e3k0yj5PkDL6cdcImnIiz5Gsoh4/Uw
Bf+DHL7Q9dL3WYAPTomtVGhMWZ/9s15yo6D1CaN17l6HRSqTUbKlfKO1lQ4UL/d4
q93XxrTBPpSYRXt5qCt0c3J0t5yHkAybCn0nFY2aExgeJ1z9h2mux7Q17lY35AyQ
qeXw4M0Hp9rZn6oSrJ6kF5U801S/1wq467066hP12nkRmD61FDlYw2zvn9wHlmyP
+4jVZZUjw7HOC2lN/6r8cvijZaPIh4wQwuNUdnw0DGdexcIm9XWx7dDr5pMNaGKa
UwbiOGxPQc8GF4V1IPrg2phvkHiZxr4eZ5P8fdTAiQV013gQnGM80ZzYh7XVACi7
RQEELYyoxhtqW0A3kNicGAanXVrxUtXicck/9IOAld0sWGHoQAtnv8R3+bOtrLBs
4taX71jlgeW6cIeA2TT36NQqMz6HwkxrX7+SJVD3W5krGfK0+xfNratAL1L2VYnG
sMXYJgEqAJz4RyqqDW0LH14lz7U3cTfpNGRpJ43lYiZ/GjyuwjShzw1fj3mDv3FR
Ptf9bYTEOVppRZQ1ZvcFGtyYw4dFNCoFtbIwDDHLc44MJ9nysgKa7T6omshymM7N
rpSs8CnMzkdWlsE0owYuBARj+xRYsL6csjoFk9obqzMNP/ntcWit7kel1079nhC6
nqboSH29ldFsYW0JDZtqqA==
`protect END_PROTECTED
