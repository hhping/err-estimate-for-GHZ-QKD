`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LM5pnWIxb/RXMjIEqg6L95uVjioHBhiuADbeDrLipLLa5cMSHZNVZfZmIVglbTfZ
rOlkhD/VMlAjfyrqPCLDcP8JH/F5xM+Qo5jLXJuz8rWPu8739/SJVWC1EoJVY9H/
KF+863f4uKpD99nUAgE0rz3ObIQ8xNIMTEcr0Ant4O4GjQybeEyjAMyYyuCPix37
rPaGk6pKC3SJmE8Z+P0zsJDXD5jtJUqiVED8kxjZOla2ng21Fbd1vhTXJMKiHOyj
6fMbZO2U/8lFiMGBWX9d2G4qowlbXyBE5PnhqLcgO46+WIU+4ROJE2B/p56/b3I3
i3GVJk5rEAjlA7YM3ceMmPZSmqRoZHhJFthcO2GGjBx8GTQZdnZ1gN2DY4PORdIj
C7iuW+0MqBuo85rVVstDNEphsXlTz2pd/NQYD0I0SqGH0Ju1EnrRawgGO+hn3idG
s3fZYCH6sfGHyHBhlheKeIpcbJCjw5JRxMUlwLwmlmzB5D/Ryi/AKuXkM8U/mZpm
84GVIYOWO+gJ6JsSNjxD73jSeft13GGstMxenyh5Kk5LW8e9O39ZzCYttD0+rIVQ
Gs/UoZamPX0zxUFTvqQWwu3jshy5l0nEvH2WCIiezdMJgSo02LQ3WXgBwCFUsP/W
2gPHU9pmtb0Tfi6xRc3041dSHsiBZ4WWp+/U1UD4PmB2ogEQCqWBKWi04P7pHFAS
QTx7gT0d0E3rtTO+f/HLbR+TGqMxE+KxHuRIueDpG+YwUsSWgcLQTNSzMEp1E+xQ
ffElHL0l3SeZmbnjD4pOCdtqlVJSZ/vO4NR+T0bKFOBClYszHonoXjTPNp02DLhP
/KbTILRTLvCrCzHJtNpt02ow3A2xB7SdtKcQT/AspZnZ/XzowmJeh+gDI4Do1bBu
AdqHPNHH+HuNkAN7FWwubLlQ3BnMP/3DJiQGYnRczzd7UbvE93JYQD2MjRPxk1yC
c/iu8BKnJgrALED+jhi92dadvcSgNQaeK2/Yx/p40R4MH03QKZAlvsj5fbGxXTT4
M1pLUizWKtQb9M8Iu4K570uQgnUwef9bfV4ri6hhxH4gMdajiyniVIKijNpwuco8
WyyIKgyz70HqRoEBSZyJ3m/C9eCUhvoVmLIOxtAWrqNb2ECDqshrkA7ixlJFuKHB
83eRbiUXYk2HVQXKB9e0eIqZukhGGNUUqypsq4OPEIy+Ibd+NXJFGkhl9vDjJwDo
mDnhElg5zNkZR2iVQhSKGBs2ae/E+uE6J/q+eTojEuV/ksfzD5gMV1m1kXTTkc3Q
bZQCAj15+JLj2neVBkftTEZ5vdsL+2MeMuwiXssCPNJSz9n4h+Bf2ImB8FyW/KPy
excV0IospqM10S8y6k/tAo0EU4AAd+DfqCe4gC3wFICmQHFIjoGBkf+kTxDut0aa
Qp6xpI4IUVtYdr1VZXrgzSqask20Kfx4Cm6rEqszhqnn2BWvhcf0MIqeSJk6Bi8k
Q8Iip40itPXxAYjdZIofibLHJIx0rY1/Z+TZ14YUZIbmZsaHowLm87TiWLmVz3Sz
qi9t1xz+4NlaMORQFhRSB7DZgPMSIzmwfbYDUdVIbONMGyzp82A92lpGSSzd1txt
GaBBEAA/cpirTP8ZQKHldrbQ7JIyH13T2edVZcwkQAc6iN51+G8PfHsDzzHudRCa
OEyVpGvJzZtIdR1phBTDmNhGI5vmb3ApEmWlcyZg1b3Kh0JwRcm6yGLq1MPYHovv
7OV8madlQ1PXP9/oe7KZjhTT0MKrsFvUQQ3bOCI6yb9oO3rIzsV258ogFyc1jB/D
p9tw6C6oKFhe5YFf8E+p8tGedS6KR3H8he7J3K+WC16PPvkxzki2kpgBRw6PfZrg
arjgKRW6zEe04edjfEZuUu7vCI9FKTUazuF2wa8mXHpKE7gn4driF9ZQLjGmTIPp
uUPfkEZq5CcSyXDskzPrvX0R2KQ+sDURr+5R1wWWa6GAISxDRZev0FFWBLuQbXrB
r8IWN7loR45FismlV2YK1/VYTfapGBkBAAAhVkBXoEY0OSLmSoBwuheTeIPgF91b
xwXpVL2kJ1SNwfin3aH0AaB4iFat2oDkn4GBJyIrk6Y6QHObD9rVykhJ7KNftMzl
TlAftLXrSLl8IWwj2d1R7/y9FiWlwA0PCfK3CwNZBRTbRAxwt6Oem0aqBMWr5mA4
EBIotrGGrAtBihpPgExso7p3fV905awget7cNmSh5D4RRrGW+FjM1wWr4z9dbk0Z
V6cl8Obd6YMFY9EmQwrYTVKBoum8TDlOeyCjeQk+0rjvGLrB0rdy4X2rDnF2Ropo
yM1Sm15H6ZwdLXyx0plBTdwIKYcjSWklPTRurxvjV4V2/0+Q4mtNioawruk9tqd3
LlOe/QJniiPChpqYsLML8tdvbT3CD+Gy9JVPPsKwhGUtFFlRuOuWDiAQ/D/scPfR
KOdfVQ5ko/i3yizShIUuAnrLMaGs2x5I7mPV0eXezzgIiCvq/hpaK1YbSS8Mkwmm
UPQWa62AO+X2lLlxIDoda1LC/2RyrlJ9Hdfk1H2u5ZH4dsqmGHJeSJkCjAuPhR8C
iGwrMQweF5dCUowA3tDSis2iR11G7d4h0U7fGku86X2lvgAigd3wR+3lcw1AAC0G
oxlx3LVzBCRAyYfcD3LjUnRo0MHQywTv6jEy9YaRNIrtWKGI90F7Fa3Zq9bg7UWP
df2r20ZDv64bxaBx9PhpPWW8Rt1i6jVtSqEflvLozIPXExeUvMcPRFrCBAWREumH
6W3qIb/z5G740tr65+aWSGIvkP7h4artJtCC0s8GdzXKSsb48ERx76pdG9nLaBMo
4/OJ1mWS+Z6I4jNEhcayGpGWyZ91Q/5qFzXErjr7r0+DlOetsBPXLikhvZe2i2Ky
cqWYQ3FKdeRu/4mXYSPLHDaAqHm500SL6u62YYtZfzYQGASBXAXYFgUMFYBSICOA
FEG4wJdKVj9/iKah9p7Xh4VWHpSW4LwHvGWIzz+Csv91ijSW09eDcwmmbcp7RRib
rBc9iH1C3BWyPwK9od+mcYXsu9QOQ12ngUS25oZPs4ACti21l+e1aETv6wrsdr07
vhEBAGgX1tHQyCgsP15H9FR27E5yc/olmiojd8dikrkG4lVDJorggBxJa7tRBS5s
UvUsZKzlCKwZNkggkMZFAsOunA+qvud5YzzXVjdlqFQcWdvfwCwM1JahIUQU9g5u
tcvZTRcEGDkfMlVShQSHffqehvzkYGgWzFwRohXkLzDCzl05gLZxyIW0Dg67Z6sK
muS/MCCbcubTBrLYqkYrxJiPd/Ik85pppgaW6fskKdiqCmXwJThq6bIMet+xmaZD
oP5b+7DhC/AuMWZraxwfdtpLPPTRZ1Z/QS6Og7Fb/I2tc+LPmS8gkeOcpC5GYgc3
zE44Y3bvsn5sndr+KfuN6RudlS4FESeCY1eWoUOnX3TONFdGOqqt2i+FJa4Z7hvC
bjbsQs54uocPVtG42PwHD56W3Gl4Uu3u87N/LIpl1+k1D75e8jkBs6RE6WOK1wKC
8p18OEuPOWeHZJacIM7yLOXsDDCDACd+3b/cE1BWCCFT+bjY5p0Vjyodu96GdneK
PUcyXWrQfsFvVTjB/j8F49COuKlrdYMBLZlY9s0GsqxPDU7mkDuhcUcrNWv3jLRZ
l6MnqhL8wF1aFwbrrP8QhserU5p7P7I4onV6MtJ1R86nRE/1JE7QGVCJjkWgxS/r
Ea8YTkrUPm4hm484xQ33AK6wmueFF2TznVEik5UaQy6xdNCgUI+GHzpojdYtrTwH
Ut0gTonVVt+JzsP0fT/p2svqDe2NNfgxM6Pl4QmyhsMzknOvd0iBHcyptWBpZIe9
oboBZMmkJkyfZ6P8boguC01AUvOllThvRPn27Rya5PfhcK+mypUWtd1xsrDdVztF
47P9jfvJCwjjtJDIM3Top2AfyA4gcVGLTNQ+rJWM+4Du4iCVhzjFDSHpsCO6u0KN
tio4sCSQ/L6yfF8R7ouQz5qagtvRPi//fVk4Nwv5tt6Injq1LdqIb5qj6Gkkmf8I
sgZbe64ffyDwsQb4FqNIaydk4869QkPF6SW1HA1OHYhrK4CccVXwDgtaHKa0jSX+
qMRaVn0g4xDgjIvUjNJxMXME+GXx64y7A7+M/r/DZzcMPEoF1W+eXlfkiVx2QwaA
roRZW77kNvBLHpV4HLnxk0D9f19+F2douEfxY5rkTM8Rps0MR18gyq5SmzaUvowK
hO4lnpFWQsJi1pOTGTQs2xHjeKaOu3hXJIYb38hBX2+eCdZJCmhIitvhf1IWSFCQ
QfIdld/vdify9q44AtvnKkEmPSeZzYnB8tUbYcPtzstcLJoMkSLNtpH7Z1EOflzM
kTtSOZa5LMuGVnrt5ERV7J6LiM5+KJaOs1wyseXZZ0hX+9PHTwCSxgR8oHZDZFsT
LParGTSZwh1R8mmkVKRN/nrUV2xS4eCt4yzvtN2pAoJiV+OmplRztt/JROM3XEiR
Sjsz5zM06rIfUI+W4IW6UI0SG4G66xEwu8cSEdl0Vxv15i3TgSlf8CMKJh2aGiv0
qxoc1pwj3yPCryykoI6xCKN3//7BppeGyhgyL3rUSYOm9e7GCEulLFA4w0U/ta08
8gXuoMQ9e75SYpIelJA/pvo0ZhUnnwBBse9EqwcUGWcpYN+5b+Lba2yx8MvjEsne
xM8WPaADA9oG1zOf5Z4EclRI6aGQGtBWjmjvj/UdctCRiToFD1YcU9MPFRpzLT0a
DcDPLoAJiZON/aZBP0kc31IgNMYWQ0kG1ohPvH/98h5aMLI+GLRLW3fcgGYZuKtr
l7X1XnHnAuFMWgAZ0CwrK7Url5JVvbOIv544exkAw1xADY6r0zRiUgpn6TNBOOPJ
K0+e7LDINdRvP4ADFqCaTmnEBCJD1Ey6svMNC0IIvnEPg1YlhpMDg+lMAS3d4jmu
AAQh6mobjwOvLz1+gEARCHY77BdRx9M+u3t7GbqR8vKDjVXEwzD+KAi5lQCOWZH9
NYjBncnnU6yliP5IwopQJOVvG2hgnlPl2S7QtXzNx1OHfqBnZKH6gYE1YdFZmVVC
vVwX89HNMeMMZdG/s9dhytPYaEPDLDPaTZn24j567YoWRwq4jqWnJqpE5jK/0qPm
sHm1o4rBJJzcCcn58817nvLSDuRHyIbFUf26VFN4NtWAfHTejVD4cor2LG9ZlyOq
eHpiduInV3Z4uoKkQw11F3bmFu7qxncap1YMFfeH2qLfIl3EJO6NoehI1tAAdXq9
FnP5psYotb1tPrv6grcwuStypxnXlMAnIe+JyS0tF/JG577VUZn7KaYwg61upimP
4YF7Jkmf+OKKz5vD362lNnEdooERcLubvcO7swUWsvwcnNipWaPlBhOzBZ5Ziht0
P/dhpW+P95TyD5QXXgWUqDgevDhi32/LxsLRPdxRlqSmVfDXAdEoRfv8LkQO9+JT
0hFiuee22j+cJxnciSM2LwhCghSV+gET01OVYrjAkGyjWrWBI+1tUq+/5Ajy9E3W
hl/jtFAKLdxGCwE9dj8e7l9rzlEbAYq89zdhtlUk+leXFjW/oUOpbTu93GRqzbpB
UWViwGFfmdUUauTQkqXtUjb2tXInTKd/1cPfB50PoW4rY9km1YiUhugeZg+OLdss
AeuNpuhOKAFCwHWKVlSmjtvoBzxiMaAZrtQEdl3p0r8/a6EzXV9hKUL7k1P+0Xro
8S6lCzi0NmZerlnunMgeNcd7kPQrRJA4vrEwLm9XKh5E9JhnoJR6LJIAhpA0H1TK
1znMtnhwOzhKwVoLkmpXu98N4ticnQvOgSAm0Ae00XBx2VrUda9ZYq2TNoNKWdc+
lQ5/7s1f02dpdd9C6AZ13eN6p7WuZu63wHf0NF4SZjbjPAOuIPxRB2ww5h5atPFb
5cQ9Sf8dm+OedFebu5Oi8MCgH9OSSrqoP5hiFE5GYLoy39hZbbgPk92DniRy3gam
SGI6uuumyDQEkp3uCmKYXZa3BAXlZJCQvBLETXsoALOy+Oq/zQ4ElWfN5m9hVkJw
nySgBGL4h+7Ey9c+S34pp2RYNR5CDSJmbe/QaGADTcfiGGaGOqvI5o6+QSJcDRpt
QjL5b9u2dujmad9WoDB1CYLDIOeQ4sLL8ajzEAJsy/8f29k5pifyeuJE2ZYtK8sk
do5fYICE/6aIfH0AuhNhwxnqqniGkE+XuDHOWOlTT8pB5ww7R+gy6nmF4snlQGtp
tD0Qfj7OmGvxeKNl99N/W0gY94WSqCtJDc+Syj+Tj7IytDL+3yLn3NS6LNeM4xMg
pYR9oReeX1dK+H2C9b4mp0vXZ0eXzRw6smLBnIdUB4OVZKGuCV0yErJnIQYM4O8j
OWFaHiQO/K6fZSJZ/nG5/Eootn+rCML65ZPcOVcfVdO5U2Kk7xsw9qGiYOFFv7el
9W6IkZAj8nEv464UGcHESpxdeIxm3G8GKFTZvccCLVqlfRZHs2o1WQlzk/CmWq4k
Z8GjaKYzS2MsN7v4YVOz4FzQMsayNfvu926gT2jtR7ew6JP1v5cpv3PN5AiWJH4J
hiek+s0ZWDNP6mPIP8GACCheXoZ762MGlNg9JCa9nGWUTpod9AaKeYWRh9FeLth1
r1XJc28gWWuNtmSq0/rPd+MXZ29Igoj1VY2YP57HbjCecnt2rsEPZORpogW5MwJM
n190lI4D37nL+50P6R+1s+rThX7jR9snF2vpjJs/dm0aEZXd9P364NOOTVkGvdiX
yjRlFSnoriB5w9IF00BEJ7asfhQA58oq3kPn5gUS8CiqxHekeGSPQ/FgmAJ8o4qq
6ldWw7QDKMu9wYJdNKk1d9jzWZ/8TwlqWPW4DwldN2fSjAQy+j1qV5wWBmN92vBa
GsBhcjiuj4Gcpb61FhsmB7nuhxJ8Nt9FZRFfjywAxhjk4eGklQmbn5xKjWOwmoIW
0366a3E1P/YpWNzAAg4EL/sYz6VzOW5+8zQe/uYwSH5rN8DxI42Nf6ngWUv2hTiY
HCstHKH0yYb2c+8+U9SmTALk8Rj81HLIK1xs9+RgshfehCb9gnhjggZdlIVRTfyb
2zRzIao+EkgR0vPw3yY6fU0nLzm+pVyfILABsO/s/luixrCiTrDq+/zfgdmCQ33y
v8UWnvcvjftRR8nKqnizUd7DTsmDjUErc58W7MMRJXKsNlbiD78dze1uF4U3YBRN
Inmxs6ZS/GLhZ+MMO2ZzS1W+GXVn6mu7EYlUqqra+FUhu9bfHLxdPoVxB1+3zQyc
inyw493rtwjLJKcWWUVr+ZsJ2t43cD9OiuJytt1nK2SrF8WbBygRwkEsdigW1kRf
wN+woVRIKGAyy3UD3fnhjIlhaBs6QLv0wyj4jpdmFdfmj2M1K+kiEYvtTvDGmAa5
798M6aYxwWee5OJtvyhvSJiPOBQB2s+oDv56iJqgL9E+Kd7xYwYx67iQ0GHdNNYh
xoBRQEloGyzs1u4DUL/F0ZsimdGGYLeSTjk6I2mrJkuTovBf27A2fteugXbSTzTv
nEuDIylXMzKsq56kpnexz++6tUuv9A/yDqVk4zSkox7lt20Cnx6UCoCrLBjV0J6y
g7tGkekJlwhWjaVeedjJQ35DyX0N906zHF7V/zaJaEruy1IjTEZgXZ2xTTam3K9/
kGfkxrpk74MMVjRHXOm8Nzj9Ex7e345bFGOi50ghPtyVuPCSL3lwfZjFiNfksL+3
z3T01PNtmVel5XP3efRJc5mtgX/yuA79svft8x4IdwerJjdUd9jIibqfMYB9wD8r
Niy5bFrA3mHMTl10zmi6rWHMulFkXuQC8fW30J+xP9MB/JBw56eZtgCJE8PUGkYN
thi0CiON4j/4AhfVO6M6ieJqTqxZAtOuCnKysJoNArxkOfKWnftIHJnhf7zF6oyR
kOm411TKmCINjMGqhf35EWhcq4NtmUnKF4jJjZibTtoz6Hbq9wn5jC+OBxI9ZHeb
IkbmFU3lOof9fwKJd2o3DweYnbMkNeL2wVMY6IEuib181/yK4se2emqZDdiysCPs
hxPT2D1FnZk0wt0vcN7n63T83jcCFJdKQ/T5e6CfNKdkyPweKe0Yz8DCxMvOU2Qa
m1vkHe+L1gPFf5rAEIgvkhX74s0fOI7MAQEnAg3Z4w0R+k/+GNrt5pQba42e73pR
qmTF1znh6rxqW+CqLn8xn1UBz+HW8buRXrLTHL/CiG9XdL3CHVL4F5RrFh1sh+HO
fVnxNx/UJmBBqZ/G/QeN5WzYKbkqqQN7me3pj88j/kkBVd7jBvnuYPdY71gUQ9OF
OKcIWNMv2U3FbF6Hf+XvicSloqNMKEiPp3thXXRuYzml4XByLQMNvUG6cNzUfIYn
+voOiMAJzPhED0ihEtj6Em0Gbdlk/+h59i3LgCoKZ2frlYKCm9SFlY1BYbuLztXp
wEnDiVHB/RuJ5NjRFXgyjvS8wpKmDyp2JYwRPg/UpUzh8S3bSEOnPdvsvl9I3ZOd
d4VS+WO89+uVj7Dy8sp1JiVTldMEH2GDluIGXBK6FG0BPN4cwz9jcjeWn4uZHsV8
TRCB1yUorBWvgio1rpmiJyfD1F9egzvMWxGLCU5aVA08VYm5GgRp3TmlJqi/pp4S
RCxOKlE18k1wza1rIhDcN7hAaRCK1b08R6Zzzf+fjAVQJsTPmwQmsR4Ooiwl/URp
j66sOkd3gQvF1TJUITapU6zFgMzfC/BbZkPZx0vN/NQ0Bw8a0cWibA/tqg8Wed8L
0VrFp5fz+q4gAelNm9ulTcYhjECXn8nwHskIul2Q76f9s9HVWBX43b1B3IDpaIDt
KesKgZBmSbCZtvu3ECmt+0T2uciyt7U1MPPiu+6RcHzPEsfVH7G+9ai4h4wRVTBo
64EHKDvXDGcNgF/D+JGKvsTxuV9jpkM9peHUvDGHj9KcrQaITolLf642I8IvxJRb
evvOh0SQ/Q88vlay+JozvZUkfaS/PLcwa/K7zbJgRfEr6IGRjrVYAdgerFG2X1Wn
hjt2NV/eerxS3yaFSTkOGMqyt5j3Py0ejBzVPDPZ/gG9K1p6TzU8IYEQCqomGueP
miCvAipc75vmAY0d9UWpN+Rmq9xUIaVrr1b5fujENCwhT5+tIuoZB+yhxeQj5cxl
UZfpjem4dOypOGOyNSo2wdhheqZOltylDVnTCo0+pEJp5xsGoXIt9hhGe2Md+KOk
T0UKaqlEEQGT+VnYkIzi3Yhg50J49OoocgD3nxtLRs0XUrQ3yQoAZfqu6+18hzhG
p0/IfQmKW+o3Oa0FeAzYwzasYYOPtYX4JSEzKlkBKEfJO9KJ3RRkOMm1s8Ce+RrP
3Schv23e6zvL4xgFEjMzrzpJTLct0wGjG+I2L7Go8GqBYAw0dIVzLjHfWaaU6t5W
asWp9ZPZrNK14ewo7TXm4Bcio3Y+7i4bp9wXiG5DuFJoFNftHS7fOsKRHb9HPdIl
57yh8IaYDtr9UMxpoz+tIFWSTWD4AWh64znomYROzMu4Tv6OXeT5CkFNWF6va2jv
15y6m6OYQIE5l0s6lr3BHrof03CX0m8KLMqbZIk0K5CDb9jzbxoC+Qw9YnLSBXyf
AZEZh5Drh+rLKQIam9Yb3L+jjWZn27aWY3TzCSGkOsQ7NlqTiLq7v+f/4m3rNFvY
3JR64lmVLjbrRHJi+1Krrb2g9qFrNLY74vQKaXlzSW9tXPwelKk7UBScD/PIHUlj
ef8IyES5ayMWFOMx8Kw1FCjJh7TOh4z3ToC9GCF9ZXCAGM5WUBlKoWTw9xb/dNyB
ifCKD/fzbk08H/MyJkOYPLwbfa818eLjcR6oHxJXw2d70eWWiRIAEet7i3QcbK6E
9w3RptQ/LevTZHql4W6gX5zRCIesWQvirAFHbxKJOmiH8zkmcayyq1RxCUUrgI0L
N5M80dZtwup2SK96MlJDsgbMJ8ypL5oBbMAuL1n8o1tZz87dISE2QPwFLptF/WgQ
d5oWc/FH5WRBCHFHnatV7TJjCPNBotrDWxXkPzvOTCcW3olaQ89UoTUk4tyha6Pu
AWyakCrS2Byum81GVaxpcLI8AQn7syJy2nQYfZ/tcq/g+4+b3PG9ptQJXRgXaZ2g
/3/Y2+vdnzrYhYdNVdDHkuXhVvtllp/FDmLtfJkfFWpWQGjbX2a3nq48B4v9uccp
P/r0U/Op1NsgeEqih6/3HjlWDIRrsOh36f4moQcc/0FUTlFMll6AVeSI3ih4xIvQ
PvZGaL89Wh0CnJVmCeED5ylVJfUD79CaSfyAhpvQ1nJrH+J1F0keXagCa4eRyrkS
5JIg+Jmj3fwcv08j8mrjrsc8e6cBcdBKo62LDO5ZOtNTtL894avczKwvKrJ0z9+W
Q28ikwjBgFxJ309oMRdibQ4wAR81xShVx3lfy4FrW5QtE2p3bRmr3LnKVUF8WUhm
BoAuA3YHHxZ7YVZyPlH16JBVBLvQ0LbcT814JhFq5345RHXDBhQOu6Na3xSuLEny
Y3psh8vPr3RSO/oN1FJ0dSJU1LNGKtJbpkhjZnU+iLjdkPBhYMKZzU0YuVphhVlB
XgwbJp/GcOcm9mfGf+VitlLKzvyFOZIqCyqP8v8wfG5mQMpa9RcE/hnhqj5twx9d
R9yP7sMQoG8Jzaw70JP2sggmt0+X+jtlhd8CYEyzoomG/7slrG+eVenK5NkCaKfO
pcrOUOTy7SHRUBmqs6ykSG8ZEDxiPhLd4RCBmLmr5OekT6Pq0Hqf2fbPpjlsGlJp
yl8XyAfu/M+pIYRY+1PaYBq3F87fBWJIWYfUWiKnbQrCJNmJ2r7fvHhU/u1PWQEP
kAl6x8tV8ROXW4VjHhHyVutSwXLv/n655GCr6tWockzSwHlQzRUr1q2OFkNhJGh+
du8+N/qEj7SAd8VuueHgA/z03Yc8glrlX8BbBkf3BROblnIGpgJMadOAnc4oxmPk
/py4YbsaP7Ylh58LgZAQ1wfEGkTnsAIthQ2gP/WupbiK0JOPEw8lXw+v6bYnr4Xa
zO4iskVlgp9AtHTOwoC1DqEvvw07m3bT5zo2mnNUAtR+ZCy3cAcfI/kpoXzGKuLy
Qu6fg3xL5XXdy+Pq6SG3ixehE/YbL16Bcb13xzDcUHfisIfn2GfdxsHzJcLwril1
k2Hog1FcqAJgKP52fZG6vMB6qBKZqNlDrFOClscyvuw2AB5pcxU1FuaNGXa2/Wcg
WP3NlNtXMe6cHtHId7Y+AS2Zwo1c684QCnzIiSD3uovGTL2uwyOBie5LJGHhnXHB
b1qTmz9ZqpQ6TZ2ouc5Cg5aIkXaxvfNVOhGRcTRrdmJlzHdMPuK4NdlG6bFpSWi0
3kRV04yNn0FQG3eE3CCxIPOCHv0L/eTUdAn6n/DJJr7dO4NMJtQ9HXjVMR4bBbSZ
q3aiM6mZ8YG4HRHgBaPqi4saoAXEqDpfNo4ZkrbdzSXEyohknAQW5tuZIcJU7tk0
+ESK1MSTNI6+WEUxqJHDb2c1FBBzy4LCgEZ7xXdrnlLt78aGvyK1F7+uTWORCLl0
goVUxca8Gbo88CoYW3DJUxYkTW1KAo7x98a8+k7qwD8XRkl1Ir0UqkgDVR5PZHgU
zsk7YDbhCOl1W+uEmTOVUiwIw788OeU0IlRFQxaelJJNQQkzwsnMRyraIvzCiXxx
SMvIt/dB9Chcn5sApl+25yGsL6nPULF7yjya73EtXZhPwcHb1bI3uUtCpCRXzgaD
C7hAF3O1jONkL2CUqxw3/gT4C2+PU+NhMqDdzwJvVvhtvl5mvJiBEqRyTqrBcOvl
RJNrVIcw+23QSirHELSMN6GV2OgZd/I3mDAq8KgeXWODqO3l9NwwUEtSkE+UXaup
QqVHVLXH1SrjwqgQlMLqa3u3leICa5bV4ilK78PK1TkLnrRrRS+TkjIkhKu0wDaa
5nKs3YcZ+C3IsPR9/El6XKw/HywxS/gYw651q/40BXukA+uGVUs5EbGtbtJ1tNLH
fqcMHbGmJZsXcral9fNd67f8LsbrJqUHGKTq8KKqeVaudiSzuY5Yguv2pKXPiA6e
35g7Q+1OP4Zyq6upJ9Tkr8mUgk8OEMkR6YUG2FsLq5yPGWH6fwcyHqqsr1rCyVmL
gAEzK5t0QfFMM7n8mPYCYacDuWVEh4WqLtXmg8YjpqC84AOEjHQD3bQee3IYdzrL
ZEROUK7XC51N+K+LOIywzm45hg+fSfv6veawIP4O5z/3OgfYUPadtPpXoLQtqTae
nycd/XqxBUKg175xpUu7H5q5MR6Zg6KBUdOJ36G5sFrRLjvIaO9h5TYxWZmTQXYQ
Y+9duHqiYN5TxhfNR3DB45NZQntMERDEzRg9Uh1uKboe6iw08I8kHmvawAT3jaWE
glHxeQLn0jP1cJOhqb4UhVF1W791O6MTjfLUaeHCgRb+/8gefK4qZNGKU1bC2GXK
MvIuE/Y59qqI/MzWsBKNy0yz9OW+Wmg5k2GF6JHBEv/b6DEHA2hfbIl9t69GqjJn
Azb4eO4fZW2DyAy1f5C0wwhSMWwf8d6ePStoASw/nJDvdQzgsyryc9wqYdTEmg61
+oohnTQkCdqdLISctDuiSu2eHVKSM50fZ7AvTaM8sXWfu5cHa32CoV4AVFWOHpLS
I+S3j0r6Z9sK/mFvwZSnpOerYsP+hyAEvOkOfIGYZcOTx0zSdwWUiBt0w1tA6jdB
9iaI8rWE2mbvgeTBBG1qP7SuSwBl+M2mr6gVQ1RQA4ARfpNazonZS8tqUgE/F2Lt
4W4nM6/Io8wwU/txDvfRQi5IjdVXz/RbF4hOSIogmf9JPVoRWefhqNJ9tRfLn8aK
6F4TYgJPFwLye48YVnCfmuYrTZv2Ao+tRLykb6SsDDifVUnd1zCQyC8wdqqPN4tr
RhwtyFCBCRVkDW0BQTQCoGiBU199b6USoijI7Eg4S6Gd5N2j5OqLtANoWf5yJee3
GGFC6ZzukEOKhT63qf6RYALA+nVZRHhrXRgKNbPVjRVGVf9bxgcPnJQFWSq6T8gm
yDpIhFjY1NqdoNtJVbVBW7Yqwx2cD1XJALUwT9Mi+QDrVQ2qajW2j83FvnMmx3LP
u75JLjZSYxDqBjwjP43vzarl2bFbDRKZjDB1AYTKDT3jyb0APPTTb+q2E7QayhCu
ojTKXL0SskpIX6F9kcSWZoxrQepBc/z9/CJYmRfSWirD4YZV6NR/zvWr2518mtSR
CRBR/yIgjdRfDvZs3gDxsCkk3lwEM2eBSwqo3n7vvs3sfsaMAWSmCEa+McNlgNA/
QTTyohAMnk2JNQN63+2vhhGoolhKYcT/AC51i1SfIbjbIjcO0Zi52f48ysVejeBO
zbo4NWcAi2WPv+jiz2xoXBoWfanpAEDSfkoa+0LtcSpuP3RkFTrd0W3xO7FzOLvm
pi0e3K5+wdVId9eLhUStPewH0QrglI60lWt3xxmV4ZZUvoP9APrsc8lOKH74PjIZ
I9/yKih+RwAha3aswltSDaYYyPyQnmLRnZm+ESapmtVEqoFpYBjlsh/YUOkTVu9A
pH/o4jSRZbuntk5kQAsUoLbHpqnh+YHHoLfcNikKTBhyFyLCAwdXnoN+P9FhwL6L
GGAAAJ7h6sQM9NFn8ImYhkYynyRHf38vPMctYKAzBGmGj2gNfiJaDhnNwZpA8LXK
yFE8IcawyKV5iofbi/M+WopRkaQOvpvaG8p2HR0LjO/MNQHvQaBHhu9Dy4quvsD1
aTz2nWsHG2vZlxxu3dBR5C2QVynfdBIfHP03BoP6uOrBM02vvABwcnvBRtZQ+zFR
fhAvOXyYxstrmr9AD7yRzmT+VsAjzbWX8ezlAAH4568iOoWoUk+M5YdvBjGS5ZAd
o8gT5dK21G25VFJIfdLlhVhyCbEu1giYTGmELlAeGWvnv9XF8n3jn8u+u7hPON/1
njpL+4zIZURFLp1uzTD+Yc2646G31NivEWK+GLtxo7wUEBLGwBXpWMJCHGHdyOMa
lSdO9EfmEn+W2rkOGYSOQZG4sxhDPJnE0zYbPv+Qf5+cVQ7y6ZSD52uUsI9/u5+I
siNMaGsbWPbUYOisGD+byf9kDf/rwhmNeOFag4DEwm+d4Y0/Jc+cSxe90ZWZFy98
HO67nPV/eL7xtO8Qgbo+TSFLxHU8coc+KOSstqjLXrnNpN9QfcolXKPWBFNPKxoi
8SS+7qxMg8R24PfINXXJlAjoL8dBUNDhja1iYAa4xMlUGeQbJ8yNxU7TWXiTMe1n
fKNpwl6eiBvFaPCeU3xt+V/8hr0ax07mjAVbmkPbJ5HBO69WDhAqElnOyShsI1gp
dNNtjdJHD7es1O+aeds0UfA/DwiI1lrjvZohUr8qeUhQiEYKMrNiwroEf+7zksD8
1EBLNnXiRO+Hk326oetP4Y2apYPFsYmuCcPcDuHvxArAPKgoyG6Y1cYAVvO/wW9N
4y2vrt8Gi9hsSiafKBbRQTNQgdydJ+lQG5sR/bzisJagqu7msjeS3KPABxjmzC6N
oKF/qCTsSP0UWuh6KNR9Xq6bYdCBs9FKunB4CM75vFcoVSe8JZ7ZYkLNGiej7QYP
qWtZO8f/TXobkCOBMcH+s7ZWq1O0G7k4O70T++WoKltmoGMKUZU2Ju7E7xwLwAUf
+8XTTUrt5W53wbnxH6SVBmKP7xiYFTv+Ll4hKZzeqXoxbvhVc0u/JnlbSI3LyYhN
YmO/8OncUWVew+59PdtuH9uRGFhQt8lIN6qVueLTyoEylTLyS/32hxLmCxl9rmVM
czM2AdM4zK0qw2ZoNU92OAV2bSeMswdjsOKy5PhG5YWgm8J1InzQOTkCVGu3AIid
+wj9mUjbuysDWWu3jvCBSMCMCljVg+tBdca9Jvspur2qSMfjEwh8TRXQ6wGCiLPc
k2gBNnr35rDMWe0SvUYgP4mt5rOdDaq8gLya3QxyZMqypKuoh6S63yfaxTTB7cIk
vj0gn3N8KU4shTvwn0I4m1+SkPSFiMM8tRcN1o8OBCI8AtJkloUQiNUWgTkij+IN
9KAfMawULG6uL3NrcQhYg/KK1HYwbqNYhgesJDaClQJuXkHYHUyibiJXous8v1Tq
R+cpfyGdaOCW587Gkx8r67HzkuKNT9xdOAruxjctgrfLTs9VqXrckFrTS3gEV8MI
hlS0/LWlpc2gfy2OCgPcks7GzyyUiNzDYJf0jz9/TVVetKf143YzRZzdlQQaBOEb
i+hfmorpCCK+DXwjk3cenIFFU4W80Mljdjv43enP7PI1KZGCOEehQZQBpc7b3ENB
wL5osOJHubZ9vsx9r4rc4t1lPY09DStlRmndeysBmJ777dOFU9m3f702b8XL6Nl1
VGURII+v0L26psXtqqY9LbgKR0bH0mi2l3rtG8EEk4joR3DMidIKTqnRNXbbM90v
8dTEvEZ9qIOYTno9VBW0G9L/1Zyxdv26R6lOTElhYYahdGdTdTrjF7HW83AFTkBD
BBz9sEY6M21xDm/cKscVHpvPECRVLXkNr5gXXVyAu/kKYlQjyb1PRyO8q6AE8Dyi
cpjruKGOVg284aX0FEAT6iVNoyqTuaqtj7bScSjR3omwZ4wWAkrrChaGXEOIjabP
f2mqd0b3JXzg7yDeThVP6qTIZ4LbJ+J3khKBuBriTbJTLcqNbH04ca/WZSEgGtFM
3bzWBIJugvxgBQjz5KPytZFt+n3hRQ48an+1j9k6it+C1RofcKQQcp+tODr4lym0
VZzXTu9Oq1A1GYiG83RQuqN9slk7vx6kRYAwjIOF6WRnA3MMGzYZiEktn8lA0n+p
UgpitKXFwjGKintAtv3IuLNC09xWVX0e3PTkl6ct8yqn2BY9yGbQ4XHTIUxRj7LQ
cU0VHaUNgLeqY59dhkEW4dWY2LuxJwP1rZzUTFI56Es2WR2q+komXmLI+m2cPRrU
d5T+vqmmiKhJdgylwMBXoI2qJYFqSoewj1TH0YgyOxpW2ArSNpFUgO3UWsERjjl0
WQ9hzlhMIejd13wOHF0xp/qvqAk0DFIDUFwtX0I74WWV8/WytdJuAJj2tU3ASsHc
VFCveOOWs3l1LznKxiXjEpKCHIASCqb7pcLlGsDVqDadESLfNKLWpy3zmM9mj/y9
S0+bGURDFPedPiXzBEOl74haoVnM5gR3e6Q6AFi7kNAV7Cunnc/qaPtmA5noPeVO
54jT4xsyEI7BUpozH9CyJ9RAg60rTO+yukUCxXXDEACbu+x68rqVjTeEBARlC2u5
PNTA3Epc025eguXB1tvXdUEpCMh7HAbS4vF1eLcpkXhWW50uO2j7A3fQubPym6SV
gxvjiHprM8mI5IXJRl3vPACB25fIQ4Mo1dKQdmLmx7nTemp1f0Bkyo2RdayS3UH0
lEFJA8wwDmKf3Dk1PYcX2O9kEQaJf5H0xpVOGwFUNptkD4aDSH4UQEh7oBwP4xwT
j+F5UduiYkuwYZKpFqPmTk5s0ry/wzVwwSMm1d75BrMciV2PvzP82BtS1rT9Y+AK
bAMzTs+JHLgX6Go5k76sk3g4j+17vKDSTUdlwyv398tzFBtxQYNsm21Lze8CRtBW
Z4HhhP+IevZjqqR4NsN6U2r9U+bOUiFMd/bd3SxskVD6kQfDnL1IanR/lo64Qn7s
VASVyrA4HBNkZwJf2dVkz92W2cyN/ty4dteCVs9aUGrNjZvBfPAHRMWOY4kVT08f
8eV3lH40KdixOEjEKi5fpeUWPAgvG3Kv8hhSK+fTSnPqZTmAnDruZz5VP2scyUNw
JPlE+AF4V/1x3I5qE/oCvvwm48VInVO5xdzN81tskYfDuYSSidjdEjprgQLUjIZt
Sp4LWcxycI8T902eCold9hmT761Qu0qfbOriS221c78XapSS/Pv5bto4+AST9+Km
uQVEQhC/OMTeA2+EvCRl+Frl2Xo4f+5bBM1vIFTsREGqIFhYhQdEuQbe6IClMrla
v5otl9MgRlERzEik9Xxf3Mrra9S4jQZ5YNT2wj4nK7+SokmVQUVIzDHlgbD7/QxV
PHb4rHja8WnShb7RA/kZszes8LRThRkWvgT3XQmXi5x47DTXYAPimoW85I7ZQWQ7
k/bYeKiQWqL0Q8Y9gPc3AwvZKa7ljQbR/WwOeYWPJK8qrIy9qJ4e1W9zZ/aJIPEA
wjPrsv6GdPg0DafHju5dCRuQd42e/pIScXbqajItdu1ac5NRM8Sc22a5FYjLLkp0
Jc3Y9LSzUCfgA6Y9j6HgJ6eZ4DeituUuPRdJkSCRCkde9Ha55XfHsN4lS1rwGKLm
n/EC3EOZvVV0yJqstiNDL/MUH9eYNj05vbvgxhJzoO9qVDBLzzsQD8K8ts6LtvHw
dATrcO6REfi4iToV1FbAOdnL75n9lqhgQQXCab5EdgqFJUgaCP0Zi/mdODZjGvtf
87DgCxeXXnjHyFiZvTuQGGrveL6SXEAa7dgUaycjLD62dmu4vJXreW0aDBYVuEyC
NbL0PQWJkl6Buy3QPgUi7Ty6qWCyADYF3M8IhuTfmOiMTKkuaXVs4TyhvRHyxvFK
SVFwpRxgdXQSDUqabs7fdwqhkcH89vISS18ZWopHoN8LE/2wcNDbg7r7WDwdDz12
+fuiNEliNKG6zU5A0e1hiCOgFVzv/Ry1RKXWpbGYBloNZpW4stmzl44bEUO5I1qS
HYH+2LBM9fRN9E/Qhp3muBzWAeosgh5Je1q5Pp9xGm0wRQixA5aa794IpIXv09Ig
75cq7BYxhKNQbYPe9BbYh1l5dfM1NnVnAnTEh9ZIUY64Pd4pPT7NzGouGTLHtuby
2fYlBDCK/hU+scpSoEn97WtfBJTSZUEfugrBv2bHLMQyVbFE2UfvGQsBmh8C7zHV
QpAtlWrSBzVZ0biii4LMdR4mz6CUS9WEqmXFyPPGnKT+9mIghTaOFqdQ9ols4fyc
OVGRtD53io4Djgv0CknTnJiywp7xpFSEyiloUqW0Ha+xdVXVMvPpRfF9XBFUkY+g
KxGK7ulUldDxuTNNKAGgriIugFke7L1in92xdsIzc+iOUJWJedM2TNcrgiArCEy2
O9BZr968N2zyabyGWC4ZIUQZ2djvLbJ81LdFEAE3pw2MllyOiggTvTWe2TbFnTVH
SrFR98SRYgCUr4y8QvwByqL3MuXEUhDOQNaWUsUs4VtIObTB4aiPLvkiwQlRSlsg
yNUrNh3CwqujyPXNhWE3sRnFHwhr7YkrdzFx28Jz3kImzPfGF/7Gihq3nzu/4EQu
TsgH272gl/hN0DNOt8Z4QkkFfyWzVTlf2UNOVuo51bDzF4MvNDqgSVpqsHAIa7wv
E2hcxLagZxWNxYKIwQ5l0mOyUgcvXp/2knexyjsJN4AU3kIfhyprkr0QypccCjIg
3YSwp8bJxV+zs6L2ShSgIi6iNYlf/GFlDdB8f14Gk0fdCElvhEflcEGIrJPCSduX
6i6ELJ5GuDIjupb/XpedEmUknlhbsAcDbQPlGX17XAk3lhhWCr2eU4MgDlNar3kK
+fIIhh5N7ShkBihuW46rnF1LWB8sjNPpNs/eBnnFkauDzgLD34u6EykznkvudHZS
exZx5FHz1ZDIzlO3XPMo9Y+amzhr4bG6QOVoPkJdGB+yTBxx6cEPzHG0RflKPBWY
aDXmfEs9TDCJ+6FPzONdb9FtQwtCNdo9xmWwzKeTr2MuA4U/0IucthoVwWqnchPd
P0hXMEcKP6QTkzmxav/UQ2fy28MjFm81qSKYUfPkhE62MAuNK7ANKW23SGHbS39g
0SLqofJaWM8bDIhp28kzEg/sYvHgQYNophE2WuHKjJK2fjo9RwqHMSvTa8OG/qIL
9c0pt7+94JPYlTVJxuk+gXw/uiHjmrTP85zOca08B7Fq3BLlPIb32jmbraLshJ58
S+/JxoS/b+uRefm5tWkqqCs20NR6lD9BYFAqoQLXCbJVJpcMMqMWnePeg84cMCw1
++LzQmVTSSOCsvGY9c+VtiMXOxeJ+BqfIhIXPeWTFv9d/xeJD77AHgk3HZRuDNHb
8MV1X8S4dSIP55TPt73YMZb+dvQo6yYrSYHjHMFjBDDBG2F1l7c6a1VC7PE5gp1p
R8q0wHU9Zgykwe/qPEwPo0WdD17LzQDn7G133EbbX10hCHoJb/CXbOJhX8FE78cV
ck1Bomsux1puyTUtvdEV7siPCWvcnRdpcpRqnrsfEKz0B4744U81PyzRUauQL1Ww
pVkNmkzN+6egIug8CL64twJseRf5I3XX01rX5Y0QcmQ2vKm+m7CH5QW0Nn4E50iw
+/5ivVsJKgTSghgo2LYjdN3F/62kVoDhkqIsyUy90aRGPdxnRFsy4O5JqHU9Uer8
2tQZc9hqZyGEKJiruEfbuvOSYS6eZ/A5gTIZIkbr+GHpOJhnkDAU4NzOaw9DcQc7
KI/jMDPeq5BSQJ+04cvyMQIAUrKkKfEiUZFoKkIlstszJ0pJ+vcISFjyqlVyn7Eq
DCFYvpO1GMosYIVPEl/KoHv5bc9hj8QiS7JvYUvoV+DZo0FvPTK4ENEsilyher+v
/Da0hLo8oyIXo6SJq290/qo4u6H7yCXHpNSOQoq/FWmwr3B+xm/+PIokZEODG4dI
u8+5Ddtu7tBwdNc8BmJKfgtY6dPm1aU7sEChobuZkr1ai2bD/R2qRsQtRHDRbeYw
FOCK21s94RFTgtwxmRSf7QVBPfGbAFZMccBjfsus+6+mEGxLF1O7nvuI+T0i3C45
0Sj7dqor+0YoXNjzY0ygZeKj0GUxaJ9U38xUI0IiIWlmANbmKsdhh9rgzm00Rnbl
Aq0fp0DW55T1pjWBX7ubReUXKgdfgxyueZrOpWMDm48QIdizeHBdspjmUgnVCg9k
cCG+6LO7FqMGdiOg9PFEvaX/3UwD1etgIhyYBj2mQiFFwkROxMVelrVe9XKulhzt
mDT0sxPExoSrx/AzkXNCDnbaDOtapWgMgVs31IFp7mD9WN4KMCEJuFNYqbCCZ21+
6Hki4ZdJGJ4ieKQ2SD5L2irck1qqn2bZpD6CQNYgbde82Y3cGy5u/cpHRTqrZd+w
Z2h4dreRnxRF+oHPgFsw5RCCcWc3ZweHNwfnL1mW89V+k9r950I5v3v7zN6h0VPx
NpsHmgeySJleJ4JX4PdebmRhRPNsBsTmqG8VAMBjvGreaQ6eO2CdzAC2cVbjMPVR
fI+hFYueBxCDalhngeflJB/9fZwlcabxgTSbi0DG7lsTI7zxpgNpqiH20beO/AB4
5zgsc3j+0b2n4Jrf53UW2mmCl2PS+cCgBfYWAKPX6ce3KWmnqhxFIVWdkIe6K+dY
DWG2cbN57oX4+xaO2hN57JXtEUmLfR6LQalD5Q9o8+Tseq4HrUx1yBxnYNDEBsSW
qtm27J+okzsCnzWXju4qqHu3RFGnIezuEaE+5QweOq1wnPrKeCKQEBWctf7dqJan
RbrLXjuPDTlrAAWb+HeiS9TgqKZscCbo2+Gy5gGNfjglt6F7imr6VCQeSjcZbMEX
J8TEuKkt4WqEezJXikhuxdjkpNJsWSSWDUJWk027EHK6+aJ0usIFMa0857FJdWob
ZID/7vvjXcE87lPU5za1RegvSiVtaebktOod8oQ+CA5bS5Ch5f+VHxpvNvDI7o9d
phD7iVFq4iBBN3qeFtHHZwn9I/BtbdY4Vgp3DWuU0sBuBsdVNqSwKsmPczTQlCmu
3XYDTExmHLm9singj7akcIvPQRV5zuxS0QKVZy+b/SFFu7mTz9v3RWrsghwDB6bz
jr596MIPhmYdVGLwgiykIVh4L4oxBvsB5dunWJ6HxnH8D3JCQpdBER6CFUfMCgoK
/vpB7n1gWKHhMlaGXN/ru7iC9RDoiT9u8CoSDLUlHGpFe8KQMgQE0m5+Ft2C+6Go
WU8Xleb0Iyol644Jm4ujipbQ6gEz3SGt9DHQdQuoGO85FbZOVpE0Q92OdlZixteQ
gN8PulUURSKpxbwAbqg5Uf2RY1s0k/cYjK/q6wG/3zxqBwW1HF+n214c+znPrXTy
rLVIa9aNI+c0+TUukhgKInaL7FCAahms8glAeB5Q5b+Yb2FW0JZo3Ni61lXxKMcd
g1Q2jgFcgxplcrF+Zv3ysvT6ewTZ1VFdP0a27V+hrKvfWbXHKEbb88ySmIt5c14h
UcGJAyvXqa7K79LsHIJNXFD0tEg18SEvOtQZ210GOZ5FZdy9wuoMvxYNfU8j9Kek
EwDxqnhS9Z8D5cvuZOVK5EfLSJS15OGVkiiiDOpipkF2ZR9A4WFPwC2aypr+YHmO
++xOn7yJwJKesoNs5SFWougGisqxbir3d5OrS69YTvoNfWxZNhnone+mgtXrAsDb
GuEkbqEwcuf7KV9+DQ/nd/3lyDbOtYSkSCMxTAO6zCBP/mbf/c+6zlJENrymQ0ow
EUkULuzUZxEXdiMgkPvUcKEMDqxNjxHWBZi4gZBSaf9z2hKfQDOGb1eEg1Ziutes
42sy9dEXtwC2d521FG9rpZmIo5Sa+WxaPCLuPmqUX895vBXy2x54ILIgaLqsKXi9
UAmlxQFf859z6+kuieJGXZXmx6YZEqVFsxCtu77ld/1G6IkNEL/g/G2vB9FNpfs1
+ZGpQmSgEI03zYOncjoagxf7ZcOEk+EuS2s9dhCS0/uvIb7paRex4S8zQ5jtkZNx
gG00M9sfsx9KNeLObgZo5zJLyVakZxMw737dlqTlp3UWsEO+WOnDzC97p/Je++kY
is9hYgCnrORXjOY/ai27xZX2B6PusXOrcCenP4JWJgCYhLa+yB5+1KyhjIzcO5OL
SWOTTk23vh8jqZxUIAZM7Su7+yYVLy+EkS3MGBsIsI/W7NGpYEHdQSvdP50vh/y2
pca/eql8f5BMNRSrOGrSItSJxxfF5K3j4xKiNZXclTl26ANgm+60Y6a8UcxkE471
5FZYV7AZc/LzuxDtjBEeoZYHHeyHzOr1MRWbAmBBZ1IBOTnauUSk55IqSwjOXO+0
XqCaXdbu3MN0UIMCcHYPNOWxzFmL/iJTTKsgSsh9zkfEnMVNM2G5DDdZ87iSkKlD
IIsPjsbCqoXyazw0gH7JAcrTBjfq8VOBZDsQIG4guq1EYqAu0MoXMBiNGZnfiyhP
4aO8QzKG6zIiyqxoabGUvkWx+y0T/0UMspGo0fFKnW7ncgbb4SfifykUEYeNo2fZ
4P2lIHxoUJqJj7ncwDeRl1vf7T2vmYgykfllFOBZwh+0SPg8f005HklpQ4F7qTtX
epcEOUP5TCqQe7oiM23YpieBbbY7EhK6GR7ez+sWKQUNtMXWJeVLb/6EedffwYnF
7Yr+ZyKSJ+3vPxxPWYSbPBRxq/IJ2HbYnpPf4E3bWji0lZQjdq2qUXkmpWacM5od
3b/l0qCx7BQxhaXKK/y50nJHxgHxLSakxQmFQxsiTB77dCeI9AJ5gcrXv44e2pNm
iK2dLP1ArpFXUJJlnboSuhSamdnBNqMMOrABS50Udm2XyueyY349hOxw0MvT2dYJ
W/bHvAFvaoHcpVKLJjkN1lLXUm7NPCLajNkK8BrAGNsGzVNc7ENi1VIgP3fXaw1k
xV38jKwQpeCaWn9ak0gc/5c/Vt46VEJ0QUR6x6nj/x1DjbplXIivN7O6nIN7T5NH
ugvUzEfz4AfLiBHm/Tato0MOc2r3CTdMsr+CZ8RIvDT7q53YcZrMwOR9SaK+4Rnf
8Se1h/nZvVCdZ+91dqbJh6a1NtmArJ1zKHZl9+7U0LJCYyeuqE+fwMpCQTFYnoVt
xYXaYom2FHWFul2pNewrEuyssRTZgkA1E0kX5803CQT/q4rdK7p1nmo+fP+ip1P7
5tjGOtzhUtC1iFtnQrZqLWpJoeATANGjruNbyHFAVv7WXagTzP1VMLgH3q1lKnpn
o98uBOeK63vf0CSk5lxTIrRHXnaGlUPDoPuQ4wNrx22Aoasqu13o4ikj24ZwlgTa
4A0HvnBYFrd7vMnY6c/mBHP8WRx+nFs26gMg0lYFyQrMfKdy2+s5JnoupZcPTG7P
FdcSSqTFx64F0i4Gfdp8sjgN5hwsCfeRZxpQCdulC2xqGDkhKO9uzk8zp+yZ87dm
jejhA1/XgoA/rm5reHyrR2jKJ09EgPxVokClMo6JKI0fxU8NnROVrURtk92d4YHA
Zn8JimwWqmBVYoLBuKC4+fWEhYcLiwlcl9uKVWuOzIKOlw0R8G0LVdWjuX0eGsZ8
DpTR5zRKzdnNbIfgzNcX84g92pFF1Yt4fhU7K4ek8TFTG1iH8qjwPdZBxU9m5v6b
W5FlyWkfgp3Rci1m2tdpJocp3O+LZt+xkw7jgR/4DI9EyimyUcz09PEUBWAOD2rG
GwEqk0JZvYGcmYgFV2/Y2nuURC9eEXOEKmPjKaaZ9uff1a+NrKDvGaJh826mrIkc
6qSAUhVVLQVPB6l7scdAVrDo4Ux1U1dRvytHJCccGu7ykEfcxcIxsMJ44d8SQ6fl
SUWNcRNC+gliYwazlOF2TvByE2sh47/HoCQq1pH75Eo4joYyx+hCtEgxofh7W8jM
drpeiap7USmIKPxg//BhqldA1+o5aRhWD8E+/cxK/uJ18Bi7Y+XDUdqtGs27gssV
PCZt9nNqyV1fhbuTG76hpSPMSJndZGY+BmWeODOjxDJAWwnNzb43E2tI/hB3OM3d
UobC4Ux69WFT5wGVJJawUuDvLocqvhVV/I19OZ5JgxF5uoFrdNPIMKfUAQ3UQaBW
r7LeTXRhSYL74uOWyG9b7QFzM9kTurD+IrYyzzGIS8iJCJuaWgB8U3NByS9gK5bN
OV1b+/Zkmi6drB+/Ornai9kDDoIsmcbqcJ/SAg3ObIya6CKs27DxdO703ey6gyNp
WZCJb5BTmQTSWRetr7ygJ84fRzToWKUXShiN+bQZyeZieRz7/jO5oagdWtW46LQW
JWrvd9MuUbeIdcY15es3QFuKvhWrMED5HK7Ixf3A8vG/r8rsqibDS5yA8i0uPLRV
lO5qosFMmStYtdgw1rl1nJUQvOr1jJfNSiaBkil27YwUtEvYO22nnHR3r+Gyjntt
eCqxnXr5V+JnJBOqH2cJlLaf4id4f/lY9PkweAEAFmbiQNYHT+g5pUgFQ2ZGh8dW
UbowEICUYZlnIZTVfqVGym3l71rqDvdNYfSV4tqpbQ18gDQq4A/kQZTzITt6q88M
38ZrF5mDghq8qF4F0h6F+LjdMPPBLOfkiuq1F8gYhmHQtxi9BYo6MyRfOQ0X7uNT
Q7c/N0GI3bw2zZXt51K+orEV+QWUpJFG5IPlCZo5OPHjb4I4OjjaVcXOR0N8qPai
K2rD3+3mx70y2jg5OSbqvqB/4gTJHVOTA+Zr2OIvz2UfvoB97NuXVxxkzT4kY956
V3dguSVQA5IDtTaTj+feN7Ufhk+41YpAy4pius4k8gQlvrX/Adiwn0OokKmfJzks
PAQu9c0sL9u3pnbbWk9HtuFZk753SVHBLDyUAVufYf+CMQBgriYO/kYWON6a8wZ/
tpGtFwXlOBCWoyLCmjF4YULfAD2+TotfHiyffIxMR832G17l6k6MHBdoqWxO8LwQ
ZasMIQr6Go9LUzHK9efW9fMMtPm5WDzbp4Z8CgNofPWFQhIGVHRYv2A85KYDdc6O
sKUz3bOMp+sJhbef8njtAppuX+bJ/yjeIGFdZyCgqTxC1s3ZK6vAQxefiFobpwJD
wcXS9Vu7slmNpizZRvqfHi0s6kS9kI+rH0rD/jZ7JS8BDLsmv8Tgdv8wY7F/MkrH
vAPpaqr60+w/juUsYd12e2q2J/Y+Xg8q5RyFLrjlOeownHKyfdiWaqVgTMkOULV7
MRPCgz8SbCNq4Zx8iIFqlY8sAkmnUk6+JJd0AVdbI+C9+gni7sAwT1V3O+Qr0lLK
5EXWoDbxv2xjBvGjg5KuDBxMDKMe7lD8J9w01i1jw4wlTh7ui4LxZsltXTIlPwye
flZ7DWg4YY15TmA50jvAe//voA2vkYrOGBdNMCAvdVyF0khqZaPSpDXwwRjHKJ5D
DAq+cfJFDnJwbX2aBRRcom1SzcFdjvzUq5pQRlBx/Z+DhesuHOea4lPedqKac0yS
9yKJlZ1opFf4Ed+V+Logq1cpoisRIkRddKTKqmi5X4hJSYyRHnZd62c/cFwLbpC2
NeK/yd+kl2cPFBoFkizIGT1KIbDOhED8qgcwo8HmA0E/Y+iEqMrQ7f8TbqiGHxhb
9gLw8PDEsts1/oeak4Rs8k/iY2G2GbK7QIcHvWe8rHnob0eDGt1fIXoYAVZbFYX1
ULeaKdOqvOL3iw3GnRcV34Iz2p81CkpPeZqP2HmsHFWxfc5fvL2XN78yAVlZM6o0
xuwlqz75TCUVaHQRTX6NYaODhTC0OYcpzHSOyWRO6FqWsoyOcdY7o8kjmmeb37oE
OEJtcuZ9EaIB1g19cevklPipyjpAWEafvE33Sxc2BhXjnJkxNWLyJWLiaK378Xhe
j6UkdIOt2t5Xk69hi6Z2WqSbCV3sFpTi0x4UmUaXetH7UtvYpflZCn+kO8VHHnFW
LGp7WJ8FhzBBBCf6DwFqFEcefXEnmtB/QNK2itAdxrfx/XyWUIjPDJue+cAVWlpb
dTX9etqAfJhzJht+GWjENHwk5o+nq+58MfZ/y/SEwrF7SYesSzOHYiNm+3sK1paS
odelBu7yhxd1gWNLAk8PeDyQfgQ1xNL7ln0D4hrchkJdiKp00MHzTd0F0bFONibs
iHnMCOOFvgy2vq/eFL7PLF/FeUmRis7lM7baFscgVHDrCVrM8djPejdznuoGWGR1
EFAVnDZV729vogeEOfF6eTixw1Tinso8plfos3Mzf6uQrlUJExAtiKoZwvYuia6V
aYQJh6NK14R3En/8Tdhs0Dc1rQXmN/8Ds7+AAv+nBM3Sw9AICzpUpQ462/xP3vxY
+LM6pmz+JzjbDuWcdzix01K7tG+LjyGXwnzDrAP+4v/82jxHBK/P00fvxEhpwJnG
s9NqXeAOozgPtvwnDIQR9xVG+P5ir7AR/sTxoeD3tb90tgJbijKNGcfwYJ77jAfD
torn1QqkTyCBLGLoTAEqVxyJKu+GNZEEtkS7FJ7dlUV9Ap3dzIatKDq3BY0ngzra
wZJTqcYPbb+8RwzP5qWjUbwFRssH8ZnL4wjtyjWtJWlnFDkDvR0qL6uhAJtinvEX
fGzZ3W+JDli3FfzyC9Mdu4jiKnRhqscr/gqswCDIlKfPZqjmhguel4rGI0YhpiZQ
psLOe5oG+gLb4iecpLXVFQJKrEdbEHcjlWBU/6E7UVKHcI2484DLrCa5L2qkVJoZ
9iK4ugTDiPotsZi+PuQ79i8QxVpTf//IzGyydj1u7bPNAYq8qSBLbKEsZFZSuDnv
Ya/1Gd2BbUk0yxuZ0k3WjAuyusrbNsA66bOmpFI/NfnDUwIART2jluMdn371rx7a
5+3mpimd1pMOm2H6c1xRw1eVtgnuU5rWPhmln9QbxHIs29oCmQK85HTR1doCW7gD
UUBNwzuG7ArUBk2dDvXyNfHiwzw95TzlUfzhdFUfMAOFyoAuj/2GItZ1bSjGdFrO
xxpN4WUbBSGMWUXIRMQjWA4UX5wLFEDKWSvEEE8LhYY4ZNOwjHkthhYnAW3NUF86
9+/akSZMACYAvxW6+XjekPddD/87d2GVXdobKZnyqmeljfXtLrRnICPbH2N2sGr8
fBLfZ1xMe8387DqhCXG0bQttxwXRbF9UyKpI5FlmJkRIgdOjtYIIM+9ThlWa0n3b
NqDQcmKSe9n1lSlvhvOQCCKXiCAFrEm1skYT3GihpEijeSymOtaek1Ps5qp6EJNJ
28WC9n9GOpp951QVZIAT/yF1r7I5AE+xkrdUGZYBnZW0pNNGKHtDs7r+RXDZXMbm
vTGe5dnKvGesrLN/8n+My1LZZAtj9BcPNpVHfIggrkuDqKLbu4vm7GZ3QZeY7psf
qtCZ6eRm8Bj5xtCeZ6IqWj1QOjQ2WxP/icvOloXqnnlr5fFICoIOGdGpbiBByxAy
pEYHaTy/T+DJqosRj4za2qJdU6DSGD0Yh7cUHrdROVM6s0a7OzBDOHs8jAm7+glv
5cYOyTCTdtr+EeFrj2p/M7MFrvhgrqNO/F3I9AbaO82FrGgSGwSNWzcixgU743V8
XaRAtIuEeKZ3vFbVhLXWICR+Yyf0NNpiHofWENpkoMaVew9/Bdksg1808Gjmcdax
XE2Q4BLLy8aXCwk2swlJd8g9VPS/dttID4WoRP1MzBqySdMNN1wmutTea75yD94x
+eZrWfHWgCk+Gth5H6Jg9Qk334wQjkMkBw/PLfcLikYuFohEqy296qFjR5mfEjiv
f0DKYHnBSOkAZrTIhfkSdsrXBZuPtx0vRioz34WGQBPP2qoUd8nFA1AihPwQXBUb
IbmTb00ClG73NnSntoxQyG8Z2CZPyKhclRL7jQeNrH46Vrbzm6rsgijIkOmvV1rU
DiEs1zMbgLb5AyIJiqz5XrCyOXW3kPlQTN7CdjK4D+ibbV8ZppZ4eB/705RKudJJ
8GV0Vc2Td77ufTWMm/+jr4AIXDB58j9fK55UFUTxWqzK0wzQ1wAJH/oD6MKxwrVQ
71jGN02w5tvPJMPx4H7e2B0ed9j/NxHXPvjLQPVEB5vfprUoB6wsPOFT0AJOwJfo
NYt87f1ZW2p8yrZvhR1Au4lz5nphBelSpdTvCyKE/iGYcFi0XoUjbJ//DCY1Fe8b
Ufd9pvpKPXur74eksl3uHR4KmoQxFPqLrPrysA+YZAg8FzHEbiQRByhk7iEDIr6M
wwjNPq6320RRJlCce+zK77Nj+HHUJW/TMwLbJjwQTWDzmokPNuY5vrlqjzeHD3ld
wMV4OHViDSEjaFGmVtV4+7Zf2aQbwpJkZoTa6/S56o+dxxNZCVVntQw7p/YorgwT
4TOq4MiIhv1jygu6RIuUigTt0SS/4t6D2xWbf133nuHFMUasvLJYE2lH2xoWTKNQ
x10m/14ZnhbpTrjgxGCsqL1hIYb/ApjQ3SvemKxL9yLuVInXhpfRe2N1UujNqnMd
gpI8QjnOUOHUyOuGJI1dEelf10MGOcNDnZJ7SiMj1iPhB5veKUSQkkc6lBdVM+EO
4/ITc6jlFijzLLxc+XbaOCg2/bAXDgG9PeuOKmYSjRqxcWIKkvsWO42iMMGRuQA6
HlLcgSnPofgxdtGBNJ2nayAr2eby3Yl4GG95Xxf0AlZQ8UJX6SBgMLLSKneLFdN3
zHBEESGFx27eyKEvOIRvvYMgj0eoJVxshKDIElFepILFIw56JXxOy6QlXW/fgK2D
j/HpWHAmNUa49GcENk5UPQ4fP+YH0GwRqhp2l1G2W9a+lw/NX4ebY9QZ03YzOTyk
jWyix7laZGg962NQM6y/AtaAfSB+8UUkmdJJWDgpJo9SpDn4a1emkfyIFeyHp3bb
hGXZL1/lgIVEo8y+5TMkbJA1+lDoZUexmURhbqv3/kKapuWpk5FMASeVFAxw4q5w
5Lwj8/YYurhEk1MUSiW30ymKaa3BM5X5pWwjSXw2MjmaLcEJaBBQGtO9EGO7hBoj
5nkfy2K+keb7NIIf+eU8vIL/Z6Bq+7SC6t3/ncifVt4D4qlrIXrGw6SBFHABuXL1
j8Th6q83JYyYwABSstXe3hoS2VcLhSm2zURWcpzVe6b82fgvTTP+nynOOuisYKCb
9t5fyRmf6754iISDv0k1OTWhcdUGy82zw8oG4khb0Fk8RD3ycPg0WbviSjPgwMtw
ghlcj0BqWCc2U0LWvF4C6/CZv3OEfqE56onQkg3TOr258oDi98A11cWuLVAB42R1
uF+bVx2f93gMIAYCsCdhAKHcvdmjqExrKVe0Qt1pfAYBki5FQWt7eQ5YYvdvYaB1
cbukhTX6PCNrxa+wZk6WUY4KP6yTrLXToV/wcl5I4/FVDAm8PNW0dJk9FSi8H8JY
rTq9+xDMUET3k2CKOuMB571qLEsL6KwHHHD+MOAUxsRkREOI0LSeBYUiB9q6BrF7
YyG+yEbnB4a62e95cqyMYJIlpH7mjtsRKCLTRzHk/MqlYGHVB3vkjYLY+wR/3kQ/
Ine1uaQYLJmHKN67jEfSr5JhaHi1tWcIGBG35QINZJkmqrVEKuKP6uhES/Guxj3v
095U7bPuG2ykacSZKqSJtv+16AKZvqdvBIYtDZlhKSATN5vbSBSYwIaEyI3d21kd
nTEJiCDB664yMrW+Y+mEmFWX0J1/OgUMU3BYD9pTMLlECdje1FejxwNSMNgMnMsi
5nWV7SAXNCSUqm9NdWj5Dt8ssCeC8/Qx9fAoy8jdoLAfAbRi0NZcxGh1fxwT6WzD
kMi4Rwx6E2Z6jlePnXoL5jRKgn2veSTysmYeT4eUcMyfEthT055wEBRIrYn9Yv2n
QgGOqI/AK/sR/7JGl3wHh8c7vVXA6djFLnKVqADQrQ33qlqbTc6Zrs0LzK9tK48L
O/pL99IXpNmeH2mRE4jQAsOCaOT9HjF9rWD6t4C4lxCnqpkdvn30ksz5Qa18P+2u
HhVK2U2Qqfll6SmDQwKc9MgpyD8nw8mo0in7+uczPcHXtUB3JBgI/2xDCVdtUx1Z
CmrhEEIxHlsEkNnpe7v+d5cty64IPqjKql8+oBnij6hbJ196J1EX4reOpJLAQoej
FQx1je7VtL+7ZjSIk1++rkXPgiIN7/o+RErb9OG/aeR6kVNszEyWhmhRaKFCB5l1
FaTSIcdLCrvI1gJTs5KeJy+en+oPly/i8DSSBUOFlDjlVAIsTQFyPxMdUfSf35NF
p4e+yuGCNbtao9UU13/huAEFPeFLh/e6DFjEHhKKBTyOKmxXj8mZW0JAyktHF3f0
F1gRFeAjHqIQBTJWCr+uewH19LlhFUyqUVRRPlN5ET5OSZkquhXlYIfNhsBIObvK
GRAuzyOpQCNR8WEp+5NDUgWTRmztB3lqkZqcd87pc0nrh6UEclCHJaHGxc0HnxJn
sHeNeNbETTL8bns4c6mkl4mQHcfee5dH4QGnQFJdt2Oago9bfVCxm9XUMjSvaOP6
4frjv5ui/Q9dICmvMdXo7vUobZsIrtad3aRWbj/0FMgKzJArA31HxKbEeCMkGJHv
YbrGHDq6SY7VodURAX6ZzIK8jCm2MI6dqT3sDBmB1MORc5W2o2ZkLZUpxMcZatBz
XtJaOo1ktT/PD57WdRUsjEZYksGS8IkZ7EvBPJKbs4BBs+rtR9YNNIn4mEAG/4/k
4NMXz0hjSVjsBcZtoNXQkhy286M6E0me3XvNsgQhZ7z32XWOxT2e66PDrshFRnjI
ony+RmCJQziv/l296UsMHli1JoPCrPldDC8zc8Gys1C7MApEUYPQ3O4I5QU/1gbC
9EHHCbPQjMcI0L3awPiqIGQeh32vSXhvYlxUttwLpWJhjVnjbcbkvD4N24d/6Yvo
oPYpMvYf31xuYDusypKNbz2IGNLvf8mjiSsP0C44hlh8fRCPwSFgqeoup8VV7m0j
0qobqBbw1cm0vZHjhnU/sXFMCgImVTbn/QW27zYv6GMMKevhMRLcg5990oGjn2Dy
vJ635OwY+TmhwJpDmni7tRlqIOuD5h9wbXl3jMbebZ9FQmLhAZyuKo6HjGFPkW2P
ZYpqUQbLruzvcqkAXEwSEGAcVwwqV/UypZLbyznH+/lQxIN34g+fh3pIZvvhKl9A
0fXf9dxW2OAYqw15acbXtqbw11lKQiRB10DWvM57N85Zw7CGW+lHIYxE8gFODHaw
qmhpZ+7OZS44+7qEres93nKU/+GiOxaWyZ5bNwfUR6ppQM8Mo+4iNSMb0CrL69Xn
cKyjoDVNFOTbn2+l/pY7ouQId4ikTZ7tje38u2zmQHbXptlb+gET5Dyq/K7m0fCP
HanXdaGg3dkQfQfoIUMrtr439yufq7LMMghS9+Dw/Zu09EqhflnM0nLK7U8LDkUC
ifrhj6amloGijKTc3aK39guX82D9cpFWXcisCmgDCQICFGoWiQNzogZHmjsVGryV
kMNkAZjgLM/heLn4QunPw+645TDJnfJnyFD/kPEXMnMDyEEwtPt/Fr0TjtiqiQuA
YQtk3Ujk7ilbJaAkrBekrvnevpmDEYsBCfjKG30geI8etRjSSJ+4VmnA/YW1AT9B
lB0XV7dF6o4oQtKUB0h3aZBsZY+4kqGHOh7KbBdEQImMpqX3JRYMobqUVsQCcHBP
TzZVPW1c9KWPzzu41vjM+KMrtR5P7MctPZ8al/6RUN9uUoS4yA+/tdbGbDktrF0W
flhfP0r9opJuiy1ISp+WZO5sZKwC0Eez3e/QizeIFRQ8UuCbOeH1fKWWte9hhGER
V+yUeDDAqU49MhlIzazmuBY6vTvqvVtFQKdFXAowJRXY0TZCOMLZClWl7r260Pul
bpnchNfPA/FozHeibtKmnD2ea1s1HDyJbWeQYlES25juKR49m/nx1hRxx5KZ9Rc3
bxR6bBq5AqRR6GBTi0tO+ALU5CwAiIjda7/qRxyABM76SExVhP+HdE2n/f2/qpdb
lwIoUgFrBo1BCcL8xVeu8OCcyU1qkG7IsaMC+wyB5Wn4Ud5mLkzr3E2EREceHYbC
fLx9pfM2A91xkyxVZ3awOc5N3Mne08b+3CmaOHav2hRCAzUa1vGE8eXgyHtNByBj
Dw/8oPSl/UD2EI5Cvf04neWvmwD5RmBEdGc+CAgkE2V+eDzDjLXBBM8VLzyGCzHI
7+KtM1vYts4NXlAHrtCn6HF4/qUNbnOnGF2ops2ASIHWFSncPKhHQJLlwnVpzEu1
h8DW++Vw2WE0QZBhKYldR5Y9BfU73+ujV/02Dka/IkvF+41ZFMGPYTk1pvU97R8g
mB8EEjInER6m4JdyetXPbAfAjzRUKe0j3xOOiRnWYn3VoZ07ZLbkTMqmQFQJxd5H
z661KgvxHFdMXEHU/PJ9L1qqwHUY6+jVnrKPNi7nhuC0+gJbtfjQ0ldoOgACKwqi
6GWH4tmI8DvS6AJEGm//n0379ac3YEZMMYwanOyxvMbpM16144uX7/wkknG47wLo
kEb9fTWos6KeNWS79Cfie7WmXrc5rsyKdHlbsQu1Kg2S8+qptwV3S9iT5WJtF3Ft
jlONcJQBiFXQcY/mIjD3/ggvaXKyfI+DxYM1zBYw6iw6T0uLPnD8HdTFHzy6BFdr
c8eVybz8iNlpla8tDrz+3Rw3T5MT0IkrTB5Hqql5x/HwvfWlVLz46UVUl2caIUtl
0zVPX+h4V/jOfSeDZIYqulB7TWDB1B32A1hTf7d50lRgqdQ0Bq8eOxG/Svm9FCt9
mXZNPALPKtxlTYvSxEfzYLGM+td3Nmvubwp9rp7VVvY+A2mk1p8wQFsVh9UctTbW
zokSg9s67NTXe5+vPwAfHIRApqbZkRfPrX3SSqBkGqdYjFr3d1poAJP4rdk2WCzr
t0tR778od1bpWoV7Lw7L2aIsyR+BD0rlhhMc75wB1g7zhHC1G8D8HGuzo6QMTWXQ
fQEwK+G8ClT41riFU8Y+ySbNhClL+FLOFIwmAgYvmbwxw0CGtYuf4hLuiK+m0gTU
PjxSq6nzcxsT73RD57rPJWIxExxdP6ZhzW2hv0zWSBApQpu6OzIxEgw7++fjGWEv
OQRnIHQbU5wWWRWSEdtfQSsMHKB2jnsLnhjwcaHJixrKIVfwGz4iYOS3bGX6crw7
YSE6Dj+NBP1orNz6L7Uk+0+GeOpiZoxGgr3o6sujZ5PpFxABYAgzMfbrkToScryw
cqU8yH3HsBb+RRSkiA/Bn5ycu7mUMOkhcvFHNBLI+/aupjOQPpshvzNjt1dYtfBD
Tkhn1Gq2S0xvtEYl3DDp4/ASL53kaidPDCTdXa330RZvY+I374NLkr8TKUpmQbsn
S1n9s4vDsYMWmALy0IT2ScJKrlPXfOmg76cdYuX5jSwmFUAHe/crmOHO9yBOli8H
F9DhJtoT77g7zOcupgARPG6/LYc4xIN1+KdxrPOaPvj/GTNjGoUMDeXmTkuw7yHw
g85LG3aVN1VnORLAA13jzmV1zwpNLJpPrXAqYtgctBU0urAUwAdAm2LtvABudKN2
b+tym8rMkaB1zYm8OpRNV4BGAgNc+rvHxq8xa2qW1z4grAiiTT1qRDGzq0D+tGIy
tGvd9nT59qHB0XWpw7EpkztqUbACDZ4Cxm6q5NRZZRYTBZ3si2230M2BP4t5INZi
EeH56PNMnBXbD+bIYCZlCr3siHpVuFxWJvi8Rh+6SDH45t26fXfqtjU1g3hLn+ef
YFfZ6yaVpaVukwX36KJsLYLdtRKpepkn0hoSV/epu33yeSHZdUtoiaD7LIdaBXp/
eJ0+vO7VWAPwIpq5tgLnNRmh5t6PV4jcTpHq3MncNJhSFiMg8QW/vTpyLua68nJL
etLB1XYNdJJHupM6MIodRK6A9s5ztwQVW6TiPeQAeihONJR6n5VJn3ujjZpAya5i
eaX84moLmvSes5yYEdXBh739wTyIiyIvlr7g34Hj+2siq949o3WADqE3hBUP4sO6
Mrh3Y5u8AB7mLC/JBxDn+dCbc9L4pRjj9nXWumM5EOX4gm2fmd3ASL5ehx5adT6N
wXZvLJAZtqwSoy33n7dSjEom5ds3C89ZITpD7pqGUstdyyt7nl7u5/l3wSZRtDP6
PteXgl55MSWChGshIV+YsslpLAPgM/vOVGeYAoKN0ugSLe+JBHcYUtdSOI1ddmbv
AOvt0WHj4iTI2xOj5u+dwFUJSE/2ph/ncqfB6Cw89dlxm/bdRE4jjBlRPUjPeylj
zqRz7uEnJXoghOBFKBwV6D/TzmsaqZAMfpSqcCYdVomGMAju4u3D164Y5z5L53i+
RBFP9HKzGbWcwUBoMlwS8Pwkd/ywsv7LbfoMiDevT8znZg651Pbb/JifRF21FHWr
JfaWm2QeBLnv1f/JBDO1LFhBCFZLTqJA6RzvY4skK3ByMsHT7jXm4jRj0evljsTU
Xhnbw9sD6Ei2zrf1z93Eqe6tTA1VA5gV7H018Mbld7gf403NFlDDyACkyIb3pirE
X2zE835oI+aKMuP6zldSM/kAVVWJylC5e91kNGP4U6pvW61H1NH8+AjL4eO2Ottq
JG3Nj6vGZW8ho7o/YIfuPEFSpTAs+PVKfcbxux9WgiqY4lYtgB3LVe6+lRjIkT0T
f6riaa6+BucdfPtiH+KFewqZNUF2fJXYnPg6XynVNGgVLA0qbfmJBKqM9/551g4J
cPirwiF4dk0D8ZpjDdLw/WHCaUBZWHyZwFMSfK31iUDflgw6ekFsVYdirfZUj70y
LfIYScj/dNvkCrnYydiOqxbUX4MJ5t1cmHGkxabc5HNl7mnM0CbfYGzY5l2diBxF
vj0HR0GMledMI9YpQFAn8EOYarlb/i9C8sAdZGAT2mrvbs7w7Kib+SAXO1sbBuos
yyxMTDU3rvhrspcZUTV9cx0aChGY9pplAh3BX2lmOPoHcpOPxruvySItBPk+o68Q
4zCcgdFSPH9SwNO8igY7Rf13nbUNw9X56L2tVXrDWWojpv771m/bi9kL3hA/pNY7
6vAYEgJiKcSQ72TlYXsz/9bdJOcV7B2d2v56dt1oBMva9rNW0okSdLiVWKlKaC8u
S66sA0BZF48zhjjvfxaCYPAZcVDFtekLQNzxefKPZ8CsPv4fkPYx6DXEBZgPdauH
SMXzH7SA2CW2NCEW0cWIGQ3evfjocJSFeMS4mCX2xiOULSsiMqrcbSJPOQPOHC0o
wJG0bS25eIXgw6/kARbU4jneCFgodI5PwOMj4JI2OB1GYHBZg7PKbH919hukNavf
z3lwBko+y9YA9enQg2n+bStIvy+ccC9uhDqth1g1Qx7ijD9kES9sA9UEcqWo6Waz
OYb50ZfoYnstLu/aTR84OtMv6RikcnxCFHIfxJv06fYabBnHVwsyYfmqN+oX/mtY
n+mbBMKW5/RtEqMfxjCPfQ8L/BchqzktiPyh7Z1ZbFF4Yi/z0lyl3Ji3I6ADxCbQ
rJcN7FkiHnu3dxJ4nlcvgmWBvMv2gKT9dqdPS+VuE9slrn0ozbiqYULewZeuZNqp
kXossyblyjGwZZNO3ZBMr0zlG9yeOGLybI/rH07ls1vr5sZnBAzjthBkMPffSThV
4SdnDWRVVdg4wlRkDqdCFazS9LQcV8aV4u73hUKP/XBE6C9VmSYHhWDCsCIAHXCS
vomq4JxMb8TdhDE0Y7W+qCSpSksACjvky4nxnk/wEE2pF4rzUs9oTDzecn4t1uwu
tr4gaKk0ac/CTEqBftPIPHaz8eXC9PE4zm9NcYeOwNmGZvTnIP4eCI8WPSVl2U3F
gYx4COVRv1EYBgQKJEItFiAmBeEnegt3N7j/QoOyuEllFzcp0Y/TamS6Lm1+0iEA
qQXzCJtZ/IpVd1T3heWxCWJAPUIXXcYV7CyrXgR39FA/eCT8aDXk9nCryt3LYCKJ
/3Zh7eaU8sQdfR+TSAvn5j5ZtJvAXefdbeDyjSQkH2UaShidyB8QAMuoA9sTG0Z6
O6+P+8GHUytp6XOM/wsHTyNS9cyA+Cyu/+zmNj46lMsxZxWc0DAQSdEOXxD7lj8C
TGWZ8aw1jnzmZblXseWMYlgMNqww6frJY9r8SPCzAYGqTEjLRo2NuEjeKBs95IKh
+2hc6QYz1qYWi9ciA0UuyyvvLRIigWgrll3uasnP7d81SAJvvzhsxOZ5ywdiJyGA
ZGXGTMDWjLFm4ZB9NpiqvRR1+Dq88nBUMM/ovAE7nBlq6ffxmmGv8t9NdRW9oPs9
0IxwCEHOPWWGlvZVStfEbsfbztsbb+uCiqYGJgx499zjYdnYaxA+k2vo7KZcdlaN
RI5A/c33ihVeodAcIFRuquNyBHI1D8T9hjcPMeV8DPRiog5CAD7cpw/W4QWLA5ho
LOUHBRHBbBSyWNAeWVYmX2O5iS0jhz4QacL43x/yqpSKkSNW68TCcJBZP4ah3Sl6
EboEjtj+dvf0sjkOuT6hFEBKKbtqtPyoT3lyefrPOm51QoN+cHqpAKc3YGLVQ67L
sNdvmyhXpUtD6cd7UdPi0E3R6XH9ZrYmD/QVXWshEEdn7wqT/X7/UjEVJEGu462a
O0EcBv+M/u+oI1dkM/Q+B3c26AesCL3xFAWt60w4Dd4S3Kamg/MKHkSr+cnN0kT3
AeahkqtiUbtaUi/CxIvm+75J5KucnXhnLhqlUPmZKoJzhhfXNYKrys3Yd3NbEv1B
1kaD+WvrXVp7RQU96sBaCfG1uN9q0ooGmBSTeCOxYRUteQKVmIjS4k38SH1aEtL2
mD/huJDJ9PS9Nn/dWeZAjIQ9/saT8ODsdkv4dzdmkUZOxLHvkKJSV5wIOAlwtOX3
0wJOX6cOGvsvoNIh6zJP8lqrMCFNNlRMF2zjb6sFp+0Zh3MtDhJbBH+/IB0UsD44
MV9lu0/fSHzuh++X0+xKfh8FU8oLJYDxY2h9GlbR9koK8bRqdfsIt4kHjbgXni+y
M9v4JOgMeWgdxt65aExhi1XKPbZ063B2hJh2v906XJ1LgRbU7C0giU+cqlHvyZqa
jF9zpJ2+kZBHRcXOLjqRTWN18bN9LUkbBFc1IvOfATIYuaJyViM6WtimoApBPiX3
b0hHrQ6yRhqUPGNr+O8gL9avC+ZEsdW4VuhN57a8enIpx+mIp/GbzdcBhwfx0PsA
aBbCQrhJZRmljPnMue6PP73GwSoQ+lW7Nay7bPDJYJz6gw7X7SbHPb8KUY4EXrXZ
kP77sBA5YDGR7hMKvqmKmQU9RRK7BFMSJHidprdIm+/ED06Vqx1+JIdZl76VZ3Aa
o1W+cKt1zSxv9sqIg51m0G7jyAwIS6UiZFdMExkGvzZd+/1FbapJeX5JaHlaD75J
ZcRiBis3dvdq4bELkZTYzdmk1ez4YItE2xL1J/DMA0k5RncI1MTs0CQqAV4XIJ7S
XDLCYNeqreH05VY7+P9sbFCCEygkyP/1RsP2bVF3uvIcPpvOLRwtDZnzhcY9wW1t
v9kIuwMivIVSrGy9hsUg/k2PLGJmLCyi6bXIHge679zV4yLayv2M0znXJIKqarIF
9QVvk4yGLj86oQhGxpiQ+HUYlwUP0Ces2S7WJ606V1Qzu5ZcaWheLMQH2xpmvxEM
MjzF6VUNKxTMG3B2Rrwf75/BEdAzMbBPr7EjSs1DvNWlXWOJQGvqLLdM0Axf6xRe
FdxhpV/iwc12adCx53vr4W+0iUT2KY1O3HL2dFkItVTu3gP9KdBJ4aSIl1sDJSFF
oYO3RGNo4yjHuW08ZBKD+p7fhRGGOy5wuAmom799QIiee9D/HsHksCzFrzs/8P2I
3naMENAkwRD48hqdCCDqM82c9c04DsjxREjQzT5w6hv9zqSu1R7WQqcUSFyS5H6e
N7CR2VhIxP8hCC4SIsoU+/9AJPY7QVz3SS5xUE6C3NiydSlnXuNUqj0OUHMI81fY
/Cw8NKAGMmp5Uz1USLfbjJhDRaluLmzxC43axOW5bsHyPDx2bim1xUzsKew9zjP/
9CV2zVJo1AH8Bv0cDm+PYNidD72AY5NLnmttz/TbggL8r0fG7rD4Y3XLW1NIv4JY
dSU4aqjRyxMK7ErbAKyys6G7q91cqyQaBRgN300VQ4O9WH3RDCAgnE7EklnJoeL8
umaCQVRXFUzOBYJYbfPwe9/PV8zQkJMX+5e6egg3N/tMYlMFKG7uO9lqTBf9jUct
F29a+qgptTxu6bOi7IjlJkeNGgIyEeO4u5WokzVBXPveEaUcL3nLJPt/RL3eF0Om
JJgzXjD0VTlGhgCPa74nNTkPli/AEOzYox86s49HhUoRPzt2bFby2QOn2PHLA1h+
2CnLJlfzqNN3Snul4O5rznCBPOQQIdnrfAjrOf5W+M3sGNRjWJE8Z8R60GkJbTsG
rC5FEYhuP21QDRCQxJUs+51OT2IKpHPd44Ew384CTg7pj3bsjoKKlOEDB8yYp+j9
vRdXaAAsg0nYPVTASJ7u1phrowGOwPKpyJkMtm6Hoi0lyLp1yVdqQABfpHPcUXEV
U5UW5CAjT0u/6q9mhcmX7T7eXl5OjZEjrgxNpR43iijQF78owqrb6TKTvbvJM438
glHn5pKxiZdJJv7MUiAVi1MOJJVVu31ETyPqxc/SJxq6Qg/s7jEKGgfqux3sbma4
83OHzUfyOGu4DkZBBLqdewCokNRWcAeCQXHNh1KVE1qE0hO9SxICJh7Efq9MWSdF
Y38VBdtBf9lEZDd3Z5cMHf3AyAIE3MDUhQh+jzSdhs8pro8ZRvQOyPafeb2DOf6E
0nn/2MAU0QhruenjCI14I0Ro5ZQzBzp9H9Y1w7fdR+fcWLqASv5pfJlcr86m8ccO
nQ+DoAUH1VUIMymS8suQt2rzt969Mgeg+XL5PF7S5C/MV8dUzxKYXUhwRJYAkLwa
RJAJB/l1Gcgwzh0fHlbfg+9UqyhBthIZk0tJpAm0w9cGuy+vbrFpHgPdCmRqPDBT
JP2tHktCtkJ1s0YiJfqxV2xyVjBURI/ghMluO3AlE+aN1u7wQSc3B8zj5FtUG02p
E2nFbV5IRyvfNHRcS1JrcNXzW2nngwpSw24tqminzP8wXZTl9C4+3dLJ9H5VdQy8
/SgAbnDu2KQV0o8SfNnbnhjpgtntBw+jTnlgUwtE4Gd1QwNF293y2Iz7q3tORPHP
pncc/lNDNPWe29czBtGWOHfiPzATOVjeePahqCkrmkiDlyrgu7ETPG2t4Y8dX6Fn
WoZwwKuiW4mjYhpPuXboc3UIyi/Bp/bSyzDHCP6V1GW4h3lA5um0MDuegJRktqMd
azHyDzX+IT5fP3qhv8MTjgPV+5BmRdBYkUIMF8P460rEcR+YdflDnW8dDHFNuFxj
fOD8xcgvhrdVsY8YSEzxXDwJWo7SIJ9LGbikk2a2wRCpomT9CTWIVsGN/hgN0xjg
w1ydxQU9sEFISQug0NQv07QWIcsjqzE7hs6nE9sCRYH6/NvW1iU/UgURsOnEf5G7
1VkyEtgi0LMU1X6TZxJAI0TAEn/3Nab6fPzOX/mAF06H4JIG7I8SF4EQZGjkeyNU
oA0q2pipx7+Ij0mxfr5LY+WfZtQBcbZ7aS10cxLyYYTLyG4jwFvdS+M+AdmA6THD
LuEAJMM/wLclIuCTaCWO2Z6OKScwGCpIwi7cLfLQwwGbOw8cTFrEHqby+0aktRE+
2F6LWAYg+YG0LwgRTqQ+WfXH89oCaYk8kaQzcg5RShQjgY8PSLg6ZbF3uxo0oRMK
T4GOCyRaIK4D/CPa1fwOnSzOuSZQQPdEuodvwhRAITUgV/LzRhoBuLivG6sucaTc
iV04sbrxfFgvFNKy48xcwT8LMIJ/JrBnhU2hmq7eQRZyc0oo7d8jff+F1aHisXi4
RpFrYeVmKPJxTxZa7H4f8N5o3uULhXimHQBYtaiWDptwyNwAKCJKMQbFFf1trHMs
jENzuWRjDRi//1ndvTpUe0JVTIUG2JV+jeMY97lm3C0W1MwAHmV52D1Z2qi7OlE6
8RdByHZwwHXlMGZeuk2wE8gluGjTArNB7r6NuS/Qwmc4S7LEWnEFul8uXG5JmR4f
6tu6ZrTgVP8+uaaBdXuQJlLlSle7hrfxOvK7dkMsgdNe2N7vwTEj1V6NiVu6XWMN
4QaREeWOf1u9kkEBzu+1MpHgtw2xpWA90Rd/bEbP5XQb5scJr5pvAyVrHQMw9a5G
MOwWcij1rftNfeBqM53B8oqzI3Getp6lJZBviXZ9aei6MnSM1g7TLhgzD7WA48I5
vjZ0VHJklSPAH9gLwJpDH+u1/H1CZBTLcoyq0c26ZuFWaLu7Dk8v7O0OuetR5tlw
HHdw97CltqbWdJ/Go+yk3dGc9EtFgoKJfPh3fS0atRTfHACHq/nx3tirxRk7XF+y
IecOKEpKYXb+8dLG6eXceuyBzKMnLHvuUEXM4i/iysW9YIL+Aon3MymPrhKL8yB4
zBm7ONZuneSyAf4UkHee3ZMOO5yh35oUI4vUDNqLc8gs3niT8fu79mAlwS0xEmeW
owu7FBOoSOfXcd7cnaQaAyeYXI7F/uBGoLtfWyZRbv968Qs8cLMQhYhhVHGEzu8l
34jRg0xGi9DJWj9+3hkol19XJB0SxCunoh7YMHAOKH9tJii2dYqcBd7sTRD/In72
H9jDVakNo6hu8jRN25eYtD4iXnpyf5wN+YsXq5E0kAp31NKtAcawHaMLi1R33mYB
5tdkvSL9Ekj31doeB2TPSG/xsW/EJO131jscwrd7o8EDxsKzshxkf/yUjBSQ+buk
wnsGEYeLcJAAIMD31ZgqvFG4qo3n/ZgiA+4Ctj93b5vo7mEz238TyCRItAheBc2N
XqzoNbnsyHfTQFGswlQ1hYIAtHt+1w5NPL4DjtWNtxrVELE56H/6XIllB49Qhu9V
DiBfWfIzY/dWvkQORyYdwyEpAaGHEjto3Qdz8gCqRcxdaMS9ukbsTOBafBqcVHfh
qG9crDQyK09vtKbXbQnDsGmD1idYjtP5lA//BsA9MZ8pK6fyx5UiZ2u8fJXKzjWS
HxTGmDrGVrfNEjd0+JUwKNEZKJ6U204a3rzHknHZlCQzKBgYmZyZyxeIz91BZEfS
Fp9qLVUvuGjNWIwIjbA5J/ZOgaIGfH03Oh3wRe9RMvtQxi8ChaP5C99gH1V9wcba
jbJz1mOYcyofaqLedfxYAIqQwYqN8UB1LmQyweCUjFOr6+Zd/qaQTkzZwKFmu/hU
TUyX3qrVu+vWflV/qHGihCRhCD7RbUfKjNPmEj0XQD2xKph0lvEXRmTsUnXxjSY3
/Xfklmffhe+gy6P0EjB7fq63TvnxEGdk4BgZGak/gRNIxkh4iYVg11pV7m4k+4a/
BRpdj3chCtbo+5KXSQZCh2R49Fge7MhOObcppHtJyJLb+VX6nZa5v4J0Taui9WuB
zrfKfxJIhBuyRLPB+xdOLtzNb2FjcgBn5v/3z0Ag176p963JB/Z/Xz3wYOe/LthR
tpQBhd3HFaLNhJ9AH/bb1IXoHvd6fda8CxOYWyGu+zdA8xskHSPMhjqSa0Lt41P6
7lgsBBkRRjCho2KfuZcafSuSq5sqlTkU2PInJUAk15YHkBSo7qgMz1dsJm1cHtuv
zMVwoONRtUmSPHkbWJzn0h+vQTsxund0zjstc9VKuMcfB0ASVLFtV10067guiMLl
M5YGXqIQHzCZM/gWP9MQsff+IUg520LFPQ/6QDV8KwWP/+76z3Tij8etw02jKbPI
6OE6Pr1iwwiKqCl5qTnExhBfs10BK6tCyficBi8axTiYHLoKJ7NEnB8zMyDCsJGT
cciWETsxEgYgdQoSYdT/Xy4yTYZ5WULyUq1N9yg2RqCOGi+1DpHAfB1UowU7zItr
J3QtP3BVujQXahz9EawqG86tTKbtcgor1KJkEuZUDbQvNpmeRWC1xBjwjmD6Ci7n
WEQoskCOg6L6+BuG/rRvTLXwdgHXe4CLDhWi53TRz0nosjzZfUvBSAeUDEhVgvIN
a5aDzwB+PivfylqPOsRsx+f59gODqm6lG9e3I8+LGWL/Mcrl4VmB1l+utkM86exK
tsMjO8zLvjdoICeNaxwp3QVKkZuRzVNkTNetlHZQatrKCvhPmtY3x+9pCLjLAimY
2kYRU54arPshxP6nwXs63dMGQqEPCOSPUfzNDbAPMVUoBrqa21ii2cj7ZbvQJe+z
y6InIopzBfrV8N7u+/KEbZsxhJq3oBQnKiKX7Q4ieMlQ5/hO3qmHAby8gSfomF7W
bKp/oEkr3CO0n44gvufpPKgGw2CO16mmMDTY0twGCTRXBTfdyTF2j/hHXMnfxfA6
yEg4Mn8t/Q10K0mVVqdf8EPaEfhNGpI9x/tjraXIEuT6XkZTckDZW11a13uHMm8z
sHIZmvjSGsSN4BYoxUoVODJDrpXWnxMr6vleqFhu9D+y4Az6LN25Qojf7S0EaNmD
1yQhSXkwHgidQD9xC/OKucNakZ2VSFWF1Kw01gkEnCBUhydZSgTtZG6pRSGEOCCQ
6gCbDGUQgDaqI6CRogmrsbBlRseEzX0PMCd5DWERyE8ylMYZDHK9O5hFS7UJQ3NN
wXoZ40pBETDX5j6FJ3w1n9t+h6yScRSRk1PXNyPuB6BbkLizxrxjJDhSdaTjBxqz
ps7EacmgfrAZGkPiv3vU0ffegl2ADviUkJvwPdfRkhyXxKOWt5pCArffnx7ERUm1
ij87cX8KYOmLs5Zc+HLaozueri4tOkEej/nvJ+ktelVuJZSqmT7F5th1YjsQOnwe
puWuLHTm3QYhP+mS/Tr3/HLgHMhSgH68a8B0JzRSJUqbvBb0HjNC3aG9fVD3ST3v
Jwiu1Ot7ziPgmrrhZhAe3NEXOFDd5s/Nt6KZYzjuYVzAWjRhtNPOXInXOiF29zt2
I9tvfIQ8lyFFWMBfifYrXND5G7vZcGYBISpA57PUOU6T1AENB0AvqEcVHbr7L75D
PdcPJDat31s82HQUMnecRfV4/XAsrNTQ5y5YE07H/KO2nK8Wnjge6B0l5A+kGj0J
oFzB0M6iSHsr5G+bvApJuJDyocRKaSqa1mbVeOrXBVcyn4nEhnk1N99c1uDsKg7J
RdKfsy6kCdrQ32OqK+no9J7gubg/oFF9BjK4yCCEAvtGm1lcg/hvobmoPWW7z1WU
e4qpMKgkbRGfV8YRFhTFetv2TRGr3lLmyAu3yowOxGVn6WDPHIaOL4unAl31TjJe
pKANyAazpUWHsj0UsJlzm/f9HUnybfw6pRWHXdoYuGmRjh1upPmVC9u0FGFCkw+0
GW+vP0rgEWUcLPwB2JuPQs/agPsuz9TxCOs+bHjoGymTuhTxvYKUpDpMELXZ3aUf
TxDcWEam/aMBWZNKeCLw/SzBx56Xgz15B40U6vKVlEk0zarP0YNQDDEzOToil7Iv
vrYw8a83E4ObFjxlybj418sorTCvZU1X+VbhcDOdGzoXDWQlp6Z1LF8mbieLkOfO
YnjoWxh1yJ8uMQTWvWR139minD7ZmB3aWFXLYl0CwPnBqOT0ms1VVYqOv1TV0TSR
3s3yodL0ybX6lWFs1gJgcHeRBEEIe9yVRYnRTkyXQX+Y22/2feAh+xOvBe/89PXb
zoIY02vCymBd70hZoFH0NOzp7Elhm+RUCxguBL/wi7ZSDVhdcd92yCL4i2FTcgU4
SglAHOWgFyNZpR5Ed+vG+RZ8BspltOK+zohhdxKobbKiLYrI6euHSQTwKnvG6i6W
dqieQs+ayX2Rqwh0+/F2hcR2r+3q2gQ+ovdUV8gN5JWEcOPbkZuN39hDgC19mKGp
mQimLNx1WpvlTOm1pB+EEM8bw8kFqdthcEycvhwSRtYkWDmbzkly1bMmL4ukFgcs
TBY4cWaQa2ual73flDv95JdSi8mYCz0tZnIaKJdWY9CdrxoMcsa+eu5yToTUwy3a
5Mv4PJU6DR3DQcOD4jBiHFCLjNqoNFm2IWK88dnhAA2h57Q6Mp8u9+KmxPEpbM5s
zdU1Yh5hmdOsFrQC9cYVk5pnn4MvCa+wqNgxT/gGOLnanBm67Ww5ImSBvH7wt40J
Bw7x5HpEeSMx+Q8y1h98E2DAiHsPm4mRTTEcDI9g0irYnmaGqhWnZtSOQEhDKasO
JTYTYWcxe+skVRU3XJkI2iUbYqL5a67LVF/KwQRHjqT0KHpE1hCfyEOu0S11109w
WnYSoeNtUnkrm0fNIqgvnG62xaQv741AveaK61OI9tHJniOmeFvwuw6/Qjq6NXRu
kp4DW/CPvb5D4O2Se3N7xU0QyG5E+1RSpDDLJBPmD0araffaTRlfbGnPLsK+tTA+
YSaC7cgsnyn0Z8TOH5X2e97Ru5pdMZ+l6KEC+9+4wjc7oU4hoPzNjUvXNgr1p327
n0oKfo8urHwNLjuz++li/kjGkSU6L0s+7pY+H0ZZtVx6ee9swcAuxRDi8l19bGFA
1gMdwTl2fC/9D0sAN9V1yIJpaVEUKRxSj4iaOL0FNWcHMBNRtmuC3C+w/HGhQlnz
li1qvnqT+QVhqaF1kwXRkGGKn9LDqmENk/nUyyrajenvUpdaO3Fe5Hr0XCDUWN6v
O4HF09UEpHGez6aC/LwAv8L5BpRVjtmJEg7ytAyqGpKNfTw0SBEJ6O/p5NhYg6xc
Ow2Qj4QhybPhTYbyMH/R+PL3Q5hzeTZ+2rq+rjcm2E4WYWZVbnBu7QDjsSc0KgYb
arI9y3lsWoz44zqyqrSy5FOBK5ZdiD2jyyvYf+l9JSJCv7Gz8o7GXvMkoyAp37sV
sS/sEo8BpY1WG4FezV57sZRX9aX+Ar5c3RFDgo44P6Z/Q2i2f2+tpT3lNH+xu9OE
A8OrrGIzktYo8uIKA1gmCSDvw2hsInozHtDsQ4XgYsjixLg9BJE3Il+BC9dPQhjf
IfjnKkSUdT7YoCbX3C9krmeqk6kPUgk2YHVb54twt57pc14zYUZl+UUcUtOFllmX
TwRlqpSHPhjYkC1omQHW2x4RiyMhwPZA1k4xOMqhQbviYICp8r27AzsWWXv0q1LG
0yMMWV05/G4L4lTd5iOOfzbFJGhGLdpDM8m7nYOTAmeSk2H4fKAMr5xBqRG7vnUD
rrG3nnG9q1iXusEdlqtiAEKI7evvbSOVjPXx/MS/NrBmUBFcbmf01I4dziYG83Hq
5qsbCep56FpIk9NJXoumqaJsY36gnDEowbm2Xef/oO3Ndw3o0f75Nl0xrYLQbgeK
okvOAcv7QdJaQTP/4FKdj8oQDHzWTpEm74Gy5EppHxqseDlT5tyBZlHzbK+m5lL2
7ond8PDZlfnwaI4JHKm0uNR+S7JwJaj1R52FL9CboqPmIRhkpAYepisxll+GoWvB
uVX9kMd/OaKRahQ4Sd7qdaB/bY9VTMb7hdo7sVmAjZJoccoz+AjM+pHr/p93TRQe
kt3ULgYzSZHXNE5Es7wVjdxMMFbCg4EhY2nLT3XGPuKBB0QZS7I5HpN6iyLmal82
ZWFXCTMamqlGiPbqai318l0KpjADlf0/24TdJo13JnneVYPb8TC+bGojvzP0BPlJ
6UcFnXXuomdOh6Zmf18Hyn13c27EnScszMNRWqnmdxdKEixovLBA4oLooAcWhWXw
m5s9O3tneXVBSXMHpNTsFgEyjSlJMAzT43JSr8RRjeZvF8c2Gt2Ff3yLufuHoXAl
hK+dcSr03KzFl2wm0uj0OCuPrxkh1k0MJ5jYEeEmNxhLh3XiLDQhhzvLzsDWdDH2
G6aN2K0KuosELOybbuf6KTnI09J4CFpEt4eYqoML6M4krP/o6spDxp2cwX7M0Uoy
jWeer/7gEwbu/MnNHMd7eaG/1eIgkzJK+KL+6+KWpSjhxopFBYiNn7IfMP1ZoewQ
vaWHzW/qnneifBsGoqVfRaPOZSWjKQl8lc8Yrpckp3FAHxucolUvTQdpb7Qh4eV8
9THfHJ7LWtLDg5tfxJxXnSTS4u33nmZ6+2w4BhMQ6wSNZOrN+Eof+b8RZ3GK+r3i
/AJQe06M4FGK6TpcUU9YYphIjynw1Smk4afIKAOItUI+9e+CjtYWqExOGO+Z3fwV
4U/htH548jEH0z3Ft0f+qeMVTag4PQ5/djpWwtU9HllbxbTKcThy86kITVjaJIFg
dS81yf8d2JjVl7mrV/Vr1DuXuZwbB1xRT88p5e+zOUoX004SXRw7497NJyXYyCnX
BgzTvVq2B3b6Hha+SM0g6TTSGVrUweo8scWrVS0HgYd7O1hCD+bH4ehYTE8tES8e
WUGuk6dyeXp6ny2SvWwKe7c6BP4EwPLs5EGhLvq71uHjEu+NRnoE4LFWZc7CC34i
ODJMDydYiMvdbOtEguMYPVb/ZneiCX7UqdB7nwa08RwN08z/rR3hksolE/XJBnz3
PMyCipmFZqYTUIhVZkKLOMPlCCkxZQP1OLu9utZpFpwURKn/GfGM2H6DRfmU8GJi
fYzkNyiOXcBziQy0HpcLTIMVRfJ42euZIyhLEo/cO6g0/B8mEB7iaj/DUyKnh7/w
5Y9K51v8nqbWXIWOG9z23K/+j4kHCsZF3jdxy3jTioEi9KsljXL7d/IbT3twS3jJ
1C4f3OCO/CEDnTbtvLjyf5ff3BQk5bMXduWhWeaUS35NPLhjckVtfpyHbbnMGb0B
EBW1kY0e3f3mr0PS9/YjK8r8CQldfmXy5x4cWJtUwXoXUZofgG6DhIuyxmtve5dY
mwqJFL0732WjE2LAaWsoDAeqy+vUexsocorrxDT9u4wg+QEnfIrpa0TMziqWeIus
GqhUuss362ZL5A9HbBq0yV77sJZV4hQ9a3u+Saq3IQXpei2NX64HJtuwxo80Fuhb
HzCegIHoSByGdZP5oJAHrSyR8j3eWO+/MGix0JEHu9ZJ4NtuaSOGfDGJVGbsWPN4
WNNKLO6xWlVFqbESu/vH1jvvHugOZCfKSjIRo3hh24Ru+C8MGnSeCzGusm9EHbwj
MedfacEUCh0J6b5S2UhUU+TWU5g3aVPYiR8I6p3IvThxLh8jsglKIUXdy4N/NV4I
mm+x/i60mBffwUSoqKaxzhQq3bxYbIFyDcq6V8xPwb+loqcU+BW1AthKa9axW8wJ
P7bHdelN4qozUIsyGfrMR2yWjW3zMkHpft4htbrr8RvF3t/Rba5OKC7SgvD7JwH9
hwKKqFFjhjwhkLopvUxKLMFxKzrjBUsyM7N8lWeR8FzwQpo/jGR3gfB9OBXla6Jh
PL0nfpJCaKppxNiilOv51Pz08cYqsVQtxFjdhb1hJHMGRjCvKAQ5gtA+MRkr2VF6
oh0X2ZA0nvA9dQWh7d6Ug32W/Firbp8nqYU11pwHa+FmtW59FBrQ7cNIND93dITP
arSffX/b0hsO9RkryL8t6F9BTbxNuDD4NaCTN7afS+xNVblKOqiWkQGvzPV41sER
BonHZ1w1TAhPApEjHsOXelqk3W4fiEAF/tIBC3S/QpoLdVUbx3i3/NaRsodHFfJv
2zd9pn+Gf7pFaS4ejEsq6WJ3eDNxTztrj9+HTuwQkwtepzl6QZ58NCZJNGBe8UwW
a3ZUd4O1fRRopFfzBTncfX7vbbi7AbXSXTfo2G2rjhxP/iUXdGoQKuVSlZUQ9fEt
tcnI67luuCA1PLN7NztYh9RNZ70Txl5XvnoHTMklsCZKI/PE9+Won3wuisr9/+58
z2QloC886t0ZuzxoiFoFkBILrAHJK4inHDInXbqE/QXoHM/tLjWtrvvT8Ap1Ymhi
atLSSW8w02Q25R+LyMU8lLOil9SAkwwIhYMGg2xhsxL8lOg21QR5X66nPmnWyXQL
v09g3xNn9RTvz0/FPMlySMSnkdXw7HuCIbLo7V56ebtbH35jjdbYIXMl6saqtEw0
iGSKgMBBVHWVmQOoiKmAdElQ7MQXW7WmUy8pF5EDn/kSX6JVFyEPa6GqJlUJ1B/n
Hzi+aB05ILBVZxwa8aPVa5Rz2p/1MbsNNI/TehSAaqFCMrjtvVOkA6Q3nco6jPeo
TUWmLjTKDJM43U9xWHHFP/9w1H4C6z8cl+lZ76wqNhhCTIUgv2F+OP8TdP4IVqph
scyohS5+tTZ/cH/FxIrWuFuyEOn5bjhfhMd1HbBST3gE2oiMfy/gENk3Y3CnRpR2
PAZ6E7nbayjwkasfUaJ4EK48TwscXftZ94+6er88BLO0eyqGW78/qz1mL/KSRUfm
hzNnzoTapwabODE/s6V2JvPsL0J5xm6xy8eYV9rDfSkyrfbDTd0FVaJZslZEBaha
Dkek394Ow+wzefuGucyTPrZjwUB0ZPP3ZaAbr/+bwZneMyg6KxTLIlTjqVEtpwwe
qmkPTykJ9f9vEMZIRjVNndMXgOJ2tvcEeUNPXPvsfJo5s1lUwi1LSwlCOmiJwS1P
bVkoO9ai+9xaHOaEktTy8IHXlVFDOuDr7pu+7R2ZNf8ByqFWM5cEHqlru3Utw0Pv
Ec9EpwDQONWIb8+0/SKPFYZPdofb+3nxtXGADge4cTxv4YDy1Z7WJEauBJy3rqUy
BKRFW+eAB+umMDEClDg0B5hhYIzozKSq/cetE68qOlZ0TgJ0LEwt7g6yQX8lDpxY
hQh+fVaVLnfBzUhB637zLDr2g2qc2KtDDKJzYTIk0wsU4guNEPBAq9GBa70NQFWB
rD5FYHrW9p84cVqD+aPH3kabzUj9d4NJPDzHG+YkdVonTCSPpOzJWLhLPUXlfHnG
JimR4A+Bles9oqcm7yNVWSDshVmDW2dTt3pzXO+R5csAcDgD1xDcwOTxqikY+bUs
qSlxImKChiU5DKbkcr/qBjjfBfdIysNxPyGJet2KmXjkzBHbUVT608bbOuHtZzQV
imxix43hhCyW+8iTBgsAbxKn6CqQniWvejnXjU+TWxnfzt79gtLgaK1tQsXCP7ZB
dQr9gJ2aasmei4meT0cfpnATRk462nWsh6Ag+wkWPd8v6TvTDyK6akRVGAKA8qNS
Xx5S6jo1hXzr3rmbi/aM/y2kbL6bI2WQaqjek9eXSa7M82RrKbi5iVhqr/RW2bEU
YX+AxiLXA8xFO1DubOp29Kt7GUZcVsELMGf18lq0PYgJozxtRD/vLNrdNWITsAfL
xef0IHitVWQYk9iVtUxUFcaQ8thP2h6Om2dG668pmTBzifzssUGNPZhcKit6wVwm
UMuTgTJOovmbUAG7xszuIK2EaPkF0DXGlUTNYVzIKNMTMvpXm9D0Lk3nSiQPoTsJ
phMFG8Zjx++Wk4seMCUSImfACEHBvR55rqMEZPREpKIpQiv/6wbX3/sC4LQwQWVq
LdoygAGvkyoumb0sPuuqIvcmnE6ojcRlSJxz476ynbofle73uwmx1gzBloWw+ZGg
x07VQabfTDGymKk01Q6k5hjiO6oGO6vrrmmgfnUh9OCTjFDkdA2XLkuY6DZjW8KD
4qShotmF1e/KNaB3JDjpR7nEfNhKdtxqiegS0Uuxm1qeoGLgu8MYFD/59cEt8iGD
Psjvw7sb+n/VXFQCBpUnvuHbrZ8Xdhr5yw/ANJV595PDuxesRbWyD83Kw1djuK0B
RUmjX8V47gNX9a3IlBSVg8J2e5b/QRcmisPuQnfwbLYYPfOZkj6fVXiWT+0Gp0aH
qbv+/iigh4MSCMabO5jeh2d9kQakR3MCIAjl0dakTqOsBza/Gl43fYK39FP76oy/
0OslJjbQkzeJrHTKohY0O+pqlvPZyQbnacoRaFM2FGoVHdwmvpIIFds06ctsozVm
W3DEmkq8q6XoTWx4osuP7CqhKy4NrkJZ6uUvSpXzqbCqSFaESDkAjPW9BrhM/F2s
i+MhZX70ijOHQXSqrQvS222pNnEiSG353GO7Yhyr7GOV01GODp8rRqCFkjpBqETf
Jk0/qBM5XmYyc3ppu31KvWkWIhVreX7XuVM+1czznmnik6yRGrTE97T1m+T3sRrE
4nyW3Uen9LkDNZrlW5Mxs7TRvCgFUTj7T9GY3Hpy+CPfmc4Pkq5XbrVuy6v7hQ20
qyoxhIky6MJ/vIzUM1Im6XTHqOUVO3etHGMRlMTVnrvHTfdZR6kDXKR7d7IMxqyc
UcwEgi7zAgka/RYsBuXfXv0gsLZNXD67j00KFAwXa2GKsigvbRTe5YY0sZHCZXBa
Kdd9GLccRgDxWDAXn18QC+W25+7K3Nx7BKTmOXVJQQkDQIzrbGSW9NolA4coOE7d
J/knhTnm6jpYCYwkw6ljAFJaXZt/R/gBRKRMXi3CIvF1AF2IiMgF36Jq3lOrOEOq
NFSBuQGCH8HJWmbd2TKLDN08QSrOVCDERnSIC0PwMjCot7cB3oQ6eh9Hd5fb/18Y
eFvLlWpg5j41I22fo54F0eOPfMCGcCTHus+gNJR6ng99S7KIpl0NQj8GYamIsXe6
AZnF+ZxnXoYj5yarKD8k7n7PVA2hBAdFlF4i2LWLIqRtH/fNeE2UjKVJ1KvLuPOA
LzmwgsIvt/EKcDKbeU95vmsa6yO769iFsrcn3Ox09WK8Q+3fz/fRpH3Eaxvv/44b
qZ74g5PJlWI72j5jRorXBfahGt76hxWs9/cIY3FqY/ey8AMQ8U6jDChs8H334HjJ
Js41w+GrrUPU8vz6KQvpbrDbRP1UD3Co2wnjC6PJ3CLBr/56twiKS9dkYy64pjMC
OJETis/llOUkVqlI570CjHOkfd5KS5WZkIgLLKaYrIvqC1BQohIXYjNz78L/Nibh
Tdj3wtI82Uf/7jcTkZd9zG/ahNQ6MiYLTfSIHjpTgm4Ad/7XAmoY7vPx1vY9NUYZ
z6Ro6PnhNt2OhFIvFEMuAUfEl8LW29cTehpN0MsxnNSuvpczZNo56dOhlXeDYmYH
Xj/q9hinbdFc9hejjYoaTFQq4XvShDrX2nQKqK8snDexFnmhU0pFXetijcaPe304
9T9Sy/RGfpDsN9N+tyyjVBvoUTvFkS2IyI1wkdszmwO4h7Uvbq+8rd2I9BoO7thc
Lp+rMqXdqr8zFwg8yPn3YG9eZeAdcQZW7qjjqdDqME875eck45wFK5gxgNv/JwVs
UaSzvYdDZE0rlEfK2ZtjP/oS+hes5q16QvQ94uz1wsubf5hVNzvfBEVor3V1XqU5
IUEHdL5WrBKWMzxozHG2TOsY0rxEDwCW0h/4Ri/dNeeJVe2Kc3Jyz0WM0r/Ji4eB
8KLB0uyJmLCSd4ySGRBaQHEcVfCPLob+HKpAdegxK+VWIv1ouCf7NKuYzg4342Cl
EN4sIGV/venwUoaLmsC9zTgdgL+IVCXYfsMZ5rxqp3QUE4j2BSK3vKkpn7b3JsSx
AmcMilfWDO21VLzNhC7D7V/dFYcsW1GZ7b2mzFIXDWbfi9S6SBMt7MBs8HUuBelx
WjRPWnqSBg20IREqdQ3hknYYxYi9AUJZF/9yeG/BMPvdIkxSv9NHXQcr+a3AiH5/
ZAFZokREDQg3dmQZU4AE/PkTzEunnsLUnPKxZWeaLS03tj0dDU4/wWaJlBJPHgO+
Vcqt/QXKmjv5G24QeKqMdKFlhVWIse0I111K4+sMofJftBxnzPSogVMgPxR2WxFG
X+ENcJ4LuZe9Cz1FEm3DyEwWcGyP9W9IsXad+hw861mknVrvcbM9reCOMz7maH3T
laJgBKIxGgPIpyTmYwE5E/2MWwOks+FfbgN5PNhfGXpYgxGe8ni4SodaycjoD5SH
MDrID7XGu+XrZ2dhpiw4vk8ZJuITVu83hKnFh1BJkondbWOZBVNR+LgXxUwhr5XI
emVM4QJTqLSjBrw0Ky1Fzc8Z039cokNZeoNc8C+ogq7hMHHcP0qH4xy6fDmOCi1d
waiyEKhjp2FEWqAagUIrdTDd/PfCsWDhPioliiZsrvBJSLTA+umDuR+EYFoj1CZ4
E2aZiXxm1D32Xd5V6RS/T+nvQdezDz9+yqA/SUhDlW8ygsHuTtII04Afvnq2B22U
m2l40vVHt1jC3kAQOH97GubOhd+vTIh862AC3qSSEmzfS9MMnyTuC4x8Umz2WlcR
fvmu7ypLIx5P8616f8O2Wc+nDwqUSYVNCnI4Q1Lbm/KFWcVTs/saM0gAq2q3ROgZ
HLsyKXEsdUz3J+FnYHyYZtAIkIIxmIN/ovJuoLLzQDw2VarJI//LoW28+PY/+Dtj
q1tKgfzw6dqynNjcn2+pSTqJltMaCYAA7kKklNG2XRh35ceSjJdVtboPN6O1KPvl
iTzOR6kJvErNXCqyMrHz0MZutfxnccBADv1dbd2OZkQyWcKUIPgGoF8O2/D2HtLc
8UUJlI9hoQORsYkiZhZPdaRnnywZOBUNSsc6n0jBk/tRGlt/0yJL6F5h+YmOrQt+
uAoH8JGkl6fYXPM2D66Ubco4qjLkWbQuaGV0Tzpnz0LZo2UXcW3D3S+TfcBroJm6
XU3WA0Wknln36L9KPxRbMOy5oOAsaq3kZcdMdGrM1aRwDBHU+n+HoRjnHDRX+JTZ
av7RtApJZIxZD0uXmvS1NpG7sk/pDBRNfToknMoJFm55Q95OE0NqEYcibTWjSXdA
veo4QzXrPQhr7/B8dt+bo2T+t1f69XhBhHVLoTyCxyeJ1QR4vmUcFXCa8KuerWOe
AtzsrMwyhNCvaCeuiBUmrD/jjdHXPHE9DrJvdWrl7zjI9lVGImTD1+9uo6TLvx7X
PxC8SKHKisBoalMCqbMIS8JJksJ9yntwZBGjDvQFkMJqCNC3uo4WvFyDpUw9GCRw
RTgLtN5PXfIsGlgIdvYylggdmGigBgZV1qy+gyXG1kCVm9ipQdwbz5CLkDhrQn6c
KcMQqBJkmU5rHlN4+hOZ/SofbjGxOJoAJcck8JBhq+6mWzaKsjUP5SMYRSwvfDjn
JrtLBxV3KGg38hx8BnIT62S55N/vg4F+LipTHNuHUWqrMiyx8lQD7qmxVLO7GruY
JbDyHtOxeoeKTbWxnBzpXAfRcruisLakxzt9um8/nGfGm7AQ/mH6sNkug+QGjIwJ
Pt/RG9fs8e/I2aO395A0FeNQ2g5GDX8IUwmLmhYEUmmBsTiKoMltaZUD4/+ns9iO
TD9u9i4ewPHuGiuM8p0GbzTSn632pZ9IMg9GVQnDlnyo9VS+2uDw1S4KgwGNXCjn
k1a+1ZqmBzzTCnG6koJ7GiCvg5Pvf9Kw8DAkx7vGv6K9LjRPcfGuXUvLkgpY9KwU
F+/RCfWRqOZkTVyyc097E6tdFdGuYzn4KM6dkL2sfWXYd7zDrqEB6uCIugF75rIc
L9Frkj5PQB7WhQKCwY9MRF/8qDQkK4xkIQMybNo8Rfeb55kkK18Ep8UzKZvmQXyW
7DTfWLGiIe8QvLnl49CRA4543pkFUM10AzjBGWP49MOD3j0VQqDDxLq4OqShUcr4
MMBBlcZSqEP+OUaXGXnpzARY1fWkQZSOXelMWuf4EGbQR6DcBAR6J5KM7hoMfnmN
1K+owEEWdN71eyBs4SDJUOzeA1cVzgSL0657CmHTB9yf9xP+HfU5oC1TORHdUZ8Y
uF8oxE/yF6pTu29dDXScYqddo8It8jJVVkx1vmGCG9/OFIb9q/+nR4k17DgtovwL
KKs5EffBAfAE5N+jcL84SMfGNYExJZiL7b509DgIMNBvo+lJblxeLKvb3ddHGt7P
Cy+ce2AtAEWSGnghPZ2KjzlFtLTU05BL8RkJ+4CEX4lPDLdr6O5z9R6VNq1u/aL8
/P45Uq29NCPLxPy+j2tjLqAanOW7tMFPHTDKbt2NubXZSBEXiHFpzwFVngPP+wCV
d+fTlJgH+pSNtKtHdW+4QumVcLh+t/5DrcBhkUs7VEBJ/179qoCtviSwSUPDGwZL
I8S9WhJVlWsfBmVPAyZ091yzcrbTYGp6dwfSOhyoBTjTPCPT/RgVmxXY3s88KHuT
Z/QgnmysTTPQUsm0s0LEhXQ3h6qVN8b4K617cadmCRAjzXOjDH0TItE7HlZdZzUN
7SA1BvHxJH56yd9E5oQjK2lRFQkAlng0bXrtXyjzj3cT7N/CafLpJy4KlD4VKHOO
Arb4cenciL/tUxo6Ht1EyW9FapoWJ6yIYtcO1GQ1GIEtpFzfKQzYUYBoVDYQlpYf
dL9wXoy5bwyN99iQCoj9JCvWERU1aZuaQikeOhCOGhWq3Z9muCNGtphtyc3pWB+h
VoERNXhEHIw6gbks1RHYe3YYx+o0CM/DSC26PYe8In5fEkPgR1b9NqsckDrXmLI5
PiAw+mmt4QCnRhzjRaUbujYQThxS7FMWdpds65YDGLMU7lXINh9ez60ik4HuEdRv
vlCTQUbjq6oPanNvvazr0oQwF7jwhsbWm+y2SL7bcUljnGIBjUAoZPXYAuto0qGn
ApUwwKIWbG5YgL6s9dGRQRXkoTRqfA3cCbpMQSMnHVNOHsaDx9IkHdSIuQ+OBolF
zxAhxz4d8BH7kqnBl4rKeCyzAyz49+4rpE9gKxZlG0oXnpLEOXqttzBzUso6jme7
LvyIumU8ZlKTzDahw3h5oeb69DgerzkeBVfaIvAOXzqrTXHsXcWV2xV2TQT0+FVq
6BE1dPT313OQ/yN3LdmZVRTmE/m4gyLmPztrzHlUz6ZdUC4BCA/v9C2pJ9IomV1b
Eme1Ew1T8InymCiilOejoDMB4GomJbG7UAy3/a7TxYbpcb8HBzBYKrQi3MLX5+x1
4aQanZeMMpZdtni07PtBK9IXT+sSs5Dx81HtErwRBKfuYjFhKR2+NEzyT0/BFa8k
YY3HaC0ad/8o60GNXYVW60BkZG9nR6fxHWttF7/mZbFy049QYt4dfEW/LAOlOM/4
WtvYtxWBYwzDou4JHZfmnClFKVneShZnueb1UIOI9HQBAmStV4Fl+a7j5QloKxJH
yKMB4rwmK8xnqgA3Qup5uvrxWhTMVSxBzY53/O+yswCalkr3VOFUCsf9DohQQHOo
h+fyhYnUQ7ih8Vsh6/Z1j94apWbEZWds1kc9e3iL8F37YqMo6/HFbkhBdPFh+bun
Tlf2PdLugKodmTIBf9DZUnwk6xLLM/fUkT3zg/GiaV69eDxqazyBvMnN+bDJI4hU
9MOjw60WEi1AMir1DwsgHMy8eDUdjNYn0m5F/AeYbuBMbNYpukeB9zLAPQIvd6KI
oNuC1JIOCcaCRb9bV3Oj8KfCvHkj3d0SgDvDkIMtIaVen8eGH5iR4hrNTHhvIoIP
hxoc69li1QxVsyErMUbIoHdWPSKHdqQyAmApvBh6fUmA4lXKZbsNOL00LDqPvTY6
TsQdgCKhcpmUGexmy5jJGlnreF7pa6oYmGsXOPGiyREMFaWE6oNhhEUQjJrVrJrW
yw+R5asegbafwIcPZo3e6n2UTPnXmCwPppJaWVnHggmzYRZkXUbNXandPJKDH9fy
GoIJs9o6IhHaqEIpjeC5D2IHRMKencs0u/tOuUr1aVQq7WS9ad9ROnAsXKQOy/Df
Z5cjot6XaWGosK0qhq2mFPVsHyvqFo370FYMyePhooK1Qbiyi976Vk037cATiqnI
EzCn1QUZZHEnEQ9qVuubptOE3OH/CjEAtJ9LhLywnWvQFenJRR5USGU8qYCjbWnS
LG7Hx6G2qTBNUeowbJpP2u7cilhHXj3qMEr5bzCrJfULPCdNSx37zlME8MskmnZj
lHHOvTD3DTY1av91G7Dw+l09FoJZt68Cr/2+Rb/l2acQ1aVcsOtcnLJpFLyGHksR
YFWPmEBRBpEIGdXuCaHzi7CONvcBZdGMOhNXQ6pC2D0UY4t1muA7DW1la8GPiLj8
rIPBd+PIeYPsmm1T60is46mq5QbASj0tfSfMsNv60N2Ih3aWP6nONqIpSoXYRmAA
wBJDdcs5euIaTydvsbTUD67sBB4pr96YlIMl0WlRlnK+IoKAI75hgbxSCLWmFrXO
DEOgjnIMdj8p3dN4kjFExJLzpGQkDUf7H/yz+iCV0GOv07IBNG5TPJjrOJvWUnan
KpMslbRPCuTUmy+Hlq2rzgjjgJ1RI3yvi523/Lv3Q9WrmZyGFNBHclEfWMrhfLi0
b2mgwJD69cytP0zHCh/NAA3MHBDcUE/7FqH5RtqPhULtSv1r8XmgUFIidg05mTXA
0xwScdZfX5NxH+RAmvXi81IiYU4HAq0sp84xioidPoW6x0bAXyC+AVGHeKS4GJOo
ABhJmzOt83B1OOa3+bTd+hcoglZ8D9vQjvpW6xOLHuHOCVg5MrJexWObPqb9Nma9
REyOTv2XtTAa8r2eG8xcDg6/JdBjhdBzOpqiDnPzomDGSAGGTLyxCQAImbozR9Mh
tXL1WU/ul1A4+5OPxBbz3wIFrC2M9ZmGNA+1Cbw0mqPcsGoT5owh3rAKsxRQTHbf
XON6EtrI6KPBzjMleyA+szfUI3N/q/P9VAc+QbhvGjJ9WvmVZnW8QEVYRmws2Sbj
4DtEwLckCE+FYGQChI5PS5kzqXYOYxlY500omXa7lRWBt1rg3TItwXzsYBUPGyBm
wxfDuxN5cjNVhNJ+/QWciz5ZviK2p9Q/m17+hUuBgorxuk4fJK7ZLQkknGvHgUIs
yr6NDxo6FrkUk7i959b/qANmB3joPgSx0XQ/KOV4kxTsmur3Kgc97F9VcYk8DWWX
6fcaP8KOTwdrs/bwuqCiVSEYxgyflgapGTm7UQnoecYdUtDAtgd9n4p7EppZ2s8L
vyxQuv3wIADhGEOZItq/eGKIcbIDhc0jg/BoeP7t+T7uFq5Yzha7L4UIlc1C50G+
mTc4VV5qp1RrkK7inuvlK2F4RRXs4DiA2z02zaH3olnXN5xiOuSDkmWAFyWIUaxv
nB9yo4VhAGi0d+SwVRgV1KlXMDPhd/kOxHsw9DZkFdUSuaMRBxu5VJykXBDJ6FG1
txsFkGkPhPjLtXJ16Xkm8Pwph/+E5nuswXanVDCq5FEvt8+JVnVjXBdHXrciHGLR
kdWGZknpSBOzhxtyDZrGoVoO6k41FQD9Ebb+fntbsbi+SpQXFzOAB1dn2Y1cRBVL
DrryORp+KZdbPxU7UaCVlic/QItMyRo20lerByckDYgdgto9zATh/MC5aFhlcE8U
LbseeOVzRZgheP3Hzhw0QCzpQTyUJ/C6DfH+3vk1bhXGLabkVfW5HUXJGnnRUdF8
oLcI/9RviBQnrTuRknhyyKirws9L5KTRwzFwK8JKF3+/0A0JZTFMXZLeqx3pW1Vj
w4xV5rp3m7XW8Z0+MjzIPX1ifd/hAi1mSC8/a/rQ7os1LjnyuNmjqGBT5GFzchkB
EWrRB9fHgBj92tjkPIdaQtZhaUXOCPUM4FqnXFzgazG8A61Q1SPpZ35ILmFGVDXr
cgFMn7+b/A7wZ2ri6HfCRYvfwQwDjQXL0P0oquBjJjcXncAURClaa4FK6QDlLodk
50qwpi2R9JswYoU7adQVjQKNc/FF1m8zcghUMA3/EkFZS28lvkpjfy7aKv3X1I4w
K7jRFzEnxnOqlBhaYbrowuezvY9xN/RGnVRY8c4JZNOLMbS6BteTRyDw41nGUSWS
OlZHN4gMI5ESZPEQVWdxnHA/zCKeNmgWZ+Tq5MCN1hS9klZUgqAK3Ul8vq8vw0Uk
OHif97qpcyBww7PCSIjH+tSTUyMt7nrF8Eetc/NPlXriz5cJPkzJXz7I3zghnVVt
x4R8KZ5WWu+dfrHJSTGlshp91tMc8opIUYsogs0nXV7VuSU8vIyC66K+0D5BvQIP
lgCQGYEi++1Go8AUB3fAR/gyRbQtA39Z0tsX75pfSCMsev4vu3I9PlVvxWOh5yJC
GS4czX2MAQsyED9lUt8GYaKVZ42PZ9OrztQsRoEhUDnSJ0rfm1Tz88HV1iPzVN69
ARu9jHeq/i1Cy2m2Jkk3lwiKpGnTcaBUmphKrLSqN5Q+93Ab0fIko415fVE67YK8
W/XKpQllTUPTUR/PnjRven9GRmJyVLRxlBjHggthG9PLGLoBBtXymccVKFwLo4ed
Z0r5rluFGCqiNRruj4RudPOSPfJ5H2Ylr1zXh28eFr10p6vprkmFJb0PhmhQAKsk
OI2yMt3coIuss3CCjjCNJ7dWIcEQgaN2rHlc/x9wNJlbAmicYU/BHr2AloP3QclV
RM3C1KoOn5UmAulcI6pTDY9oazyfMt52K+KJtacsln8848X9DqsHRO5dv9NHQhBJ
djw5GHcgYlDykDl2KbBNYG2UbIIZ0F6YT191DfFv1ES4L7K5iIiJuMyAoFZJSQXu
HfRAYjIook3rEJk8LR1AeRpWvOJW0DlmF21UgQHwwqe0AHCUJPzKO6SmTSt3UIBt
vbleLm4K1tAdYLu+D+Uh/BSui7+B7/NLOv+WZPlReCkEJdxSzL8UfAWwfn67cgOA
LQNQzCpat6yRnCKKXvcKGUlsbs2PqNrEq6igKIgDVSWLWie9JQyDTzqmCfdd9WF/
ueCZVvn6AZZjRnwKL2iXp1rH+VbSa50H5hiY0Svgl/d9SLOFKQfbfLoKoUmKaOTi
wSIxQI5FIcefvYp7CjWwZVky3Z6AR/gP5rCVvBhSIP4wl4V5gMH3lEBqcb+M9XrZ
wKwtaf5uhnXv49roD8niR5yCL1mwBh4pwhKWKrBigNTpiEatCAQyrLU4pjXqFWLH
Jy+59A0+ctLF3RAHpO8blTDDbfnSkh1+WmLLZGzlVXIoRkVf/KatYJt/VOIZnQwH
QRATmj7f0Z+/uTzjFnrJFJ7Rw9zzHJSPwDowXut+yOwRwoJ9iTjA6kk/TmkpQvRI
9vBqgrMY3Jwq5gCx/X7zCsWvl1LU0kaT9J0ZHiDCNHSPOV3Byg45huFiamYYptUa
Xns10UXsm/+d/62A78GsS2czbsbrdXrF6IOiZpmyh/yQGDkqra3qUm4er+tyb+et
NuAU6JhH1NdzXaEDq8664zL7OJMPUYL5PCa/mnzeLSJ8aE5aOqkOL0oxdauBu+R/
nB2uWzBp9dZIV8glmEwFTbOhxKneJkyB0KisuRWQ66OmZtskojMxpke9/4ryT3k1
f4VdMp1q3Nww9qaOrDZNDt9HqwAdvnxTvAMRI/vR4/TTyvLLhUqnjQD/hv9SF19i
X1vl01wIccdi3E/g1jEq0gZdiz7CDy5Rdi4VpgX3K7YiDm8kO/I/41RT7HWOh37o
1Kw3DnwBxmcGTcIhnsWvlwvmTSeRPRo1LIwbWHTJfD9F3G/Dsk0+DRZ635Yl32xy
P2sL6n7gVRVATmHOBMbyZ3zmZZyXOR6V3uYhgNwkgClSeT8+pnKqjJ3JCITOxfJG
fkM0mk6gkCJn9uWgLUzPOVm4T3eOxQ7jPm+ZNYLrhhj18xS2ePyDmb+qO2Gqylv7
Pn/7b412nwKDVxda+7eLkB5viwRjWMspEsZbp0LV+CC1Fnd7CBwRQDaT3+kcIg5p
HIYgBLlQgns/stsdduHwR6RV+4/PAIBf4tSf41qBUtiEt2DXlsX2lHog2tOof7Zm
H2UiJRqLWeKSI7BKdNaGwZQ9dyg6BN+Zh7GCfEOyt1v/kMtPXvEbQZKlIh0kqTyn
+DFTXn0WUskI31Fnps+wwQ025rXYMqa9YmJeXVSpIWRfE/hYEGM7omYjNK9qOeCI
KZIAiLJIM57fYZeh4UlzAC7ZRixTZq/1VVPYPrvYIi31jJp6cs0qSH7Kvl8MtRPJ
TlmXdhoCvTqzbDHco4hmMpF1VnXm7aVmovd0ycjnUd062D0nisHLgFRN5NfPZLTD
u3Ja2qD34VzQLC36j670U+16VO0pGNaiU/jATVx1zlk1cO073RltTo59ZN2A4kVL
jHFiX7zsl8ntMtLUEe92SLaCwNMmkwOC42WbxMlCPHaqBFtKx0PMV6GX8ngoAfA3
pDYMLEe7AcGdl+eGSORIxfGYA0CZrDPSq6JBtWd4JNzwZsao1b271hKb3v4fP9Hf
kh+xX6uKjHdyj6UXVeJc515pGIdGZxlKqCUOXuWpmaCi6QYZC97ECnyiE5ucqLgx
aO1hYfR8i8PeQUWyzFgx7NcYqfwNPWb6oZ4iLkInmZ5vJ6s99QdZeIUpPHuOYOCy
rcPITklcYNzriPHNScFcsKKZY5ZQVRxyDLyPq9wRpNs1ZsN122A8kVTGSeQruHSZ
kaJFr1sHDkzjzOiQYpDw/NHzyRMkZJ1+sTowWpP0EvY=
`protect END_PROTECTED
