`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcV35CYf9s3lbUbqdZQJ3V3QAaRZN4FRtld5lEQAkobNvk0du1VJGj81uAiTEI6M
ZUs37twr1Wo4DyFLniGsZQz+jmnrFx9ZsC6tMdn4oi4fOwM7dPYrifTVOaBeTnex
MuaV+qy/EbbI+sxzn02UcFuewFa+jLoJOWE14vbe/5psJOi+pauu17eaQsNJY5Vz
V8XiaThL6pUbdX+3jBww3C4Qd+7k8K10kx+UTInxpQ4ZXUg8kTzElJUtJbviZHtQ
JADKneZJO6bPS7b6zpBdjvv+zYnwZSh9DR1fh9V0YxMsryPeSNpEvI+bCwHJc9zZ
Y5AvoxLgv8s0Bbdthyw+8S4zRnb7RbgIkmM6X4Fe2vF/AJZxFuu7ijFAzhXkLyxL
mJwCf0FVaOXyCpi5J8Lty0BdjVh4zEdMRMO9l/TdhXxYdyS6bGd1oD1ENMlbnJDG
bj2fJK5hDfFXP0UWdqRMCWhIBbRu4ZK3IWkC6+LUXP4RnCylAPjnrPVF0CJfwCj/
yq4OyY6bwlmTAuKT9AO2JFkAE7HHqirQMLG/0rQt7NoeyE/r2GaBhd9GzyhAdIVR
pckZIoIzrrQOoyXWM2ouKdqQa0qy5OCMy90+OYgvSgcL8KfOZ7ai2PseSPFeR4St
+avA+sdPVCZOOhGU6ySID80b7Rj7zZb2v5kfTSx+2X4SyFg8XQjdD9mvJfPNr/79
VCh3If2ebcegL271U68AcMQHQyA1GxiyJ2mSefIAbjTBkhpS8fn1VEhFK355AtLW
2tPmVyafWJhDS7bgBia3384MkRvwK5uEvnS7l5QCcPbjFq2P5dCt6YdDwj4QENij
`protect END_PROTECTED
