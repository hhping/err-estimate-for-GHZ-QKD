`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kut2e60d2m+4nNxsXqxPJkxiNnKD+caciXHr4wSS/SG6ccya3gAalGbdaOaNJWuG
IgU5oNsQ6SyqFHGQAa15gdlDkUASq1lo5sHScwNJLqJIsX/vK1hfx+psnmRHY61S
EmfpqwWKEM+vwY8N6dl3HIKdzLstVCKDtJZrfqq1Ojj3lV0+nBVhR9Ss1CgWoywd
GfzlhAr8FGjX2MtT3oD75/unJlhyIpvwR1Rir989YNNXBWwazdlf9ZqoegBAgUfO
qLfkDJz+E25Ky0rdyLLuN8macukVyTeASDbGH0dBeMkElZRtHRRSguMJCwl02giK
7oyEVlL3vblM3M/mdZOqLZwWxYAwBXX5AWl3l+8SsdvwUlTlHGjtoSZfb27rqPF0
WpBufTdkfyUntf7XbYOXXqFk1/bK6mJLFNl0GL5h2m5lYSqxaI3fDsqd+J9pAbFh
GpUJmE1yj4Z68A2bVp8bCx6JbjrTkcgWyRyVWBoR67XNtkXz1qmcunom5vvyOSpz
5Dxt+X3VUvBA3uEZrLIlYVL7PrIDhp/MGD6jzfCbNg1rxn7Ih3d6SsbYmDjNuM4m
Bt4G1tsBhJSiEFihgS0mhxCup4tlfEVHEIrDYFhoBGhjEfLgRrKMk0KygfKFXrPI
fBu96qWjz0JimbSRTLbFQOi/+B0YpQHbs4PVslQit6cdTfQwBPTqy9Jt/q4BVeHR
vbwUQqTYc+7wHWYA7pyhO4ybPKNg2fkGAR+biZ4Oafr2SjcQXJmYWw6M0I02qqAN
vSH7uo/xHy8FZUDyiGHGcAmn3YlwnRD5Psgzk3a4+T44EV7U14ne6nR4Vu7JbAin
DYpfgV7q6sJpoJtFn8CijfEnqf0R11bVKGC+RWEMRWsbVZ5yFuovDwMiut//NAeq
jzTZTAbkPZAEw0TTZ6yDU0dXRXetyV+IEujS3Ly1BslcE3nhOGa8NbmwZMKXZ3+3
mHiLgLzu3nBClmMzDWdXiJRf6QxkEAG/OYWq6uKMGuGHU78F61aegcDj1owvvSqx
JYLlQsm2dxq/A0KuDPKpFvlQ+VdmXzDtUqk8lPDLJRU4LmuE2KWVBdCn+2wSQtmv
hqX0uutNxbutBeZwQ6BV1VIqRgCaRrjya1gyqIREo/9sc65M0Oi2HSIZIfAYQmuP
mChaB+i7YB8M8Q96fVjSZR0Qn8D20DWU+7Zs8dzWpGXoddkLREnzqRVcZKJIm7J9
UcvNGabK2ua1JdVFeBdhFdvNStjwDU/WtUAA32XPLPhjJ9AcB0vl+uW8VEF8KN9z
rlmR6aeEK0edVOXxJZ3BbIwdm+FL+EAnZW1TLf76PI7GbEZF0TSPSyM0+lgYFr4X
Eh+NEioNGEaS5F/XKFUOi57i8cUA8JqqmbSCoIk9OvyPXX8Frd70Zb2NGC8eoDsK
qhu4HgplbBa4FEkvGTWfLSf7nqWdyXwSs3wxgQ8Z/QFtBXUO1lXvsqtR0f8s1N9/
vd9J8BbBR8kvEhEQB4OOEyiCJ7pbEoaT5DDGFweFdWKMzbIu90V7eR2/nyIXL+yC
5xvSzkNq+yqHtSPlVhDtfLxvkh+WMlDDLmERb9GqNn9ss1K+XQjWnnHXIv1SMXHQ
mC2rj8eL56ETo/oRGcYsAHXwQolViGH9QeJpaNMg2cAbc+XpDIOoXvw4FvvIpHUA
rBwQHgxUogiE7oWebyR7/Cdt3k8bXcnJn2q8ZALyYuK/Xcy8U9tzDQPs8OI8Joy9
CprusnumDb7Osvo46qsy9XLG/Kg+YqRvHAPfBZvv/Smv3hB+/HJbDtWaS6KXZCML
YNnFI09kPY4RAiT8pw+26hKMSkXxJOiqXJvVvU/xykCgI1K4zV7O+t3mK+dJBvtD
SI4tl76phTMucQJ+ka+SYveVLf+aPPngdyt5VfVQndBe3iPT14BMga8xLesrzNZL
xLtsrJTJQvEc88LIFLkhZxcTuwHO43gwphAE49KD2Q3Jc0WdaarZ8GF3Fatc2aqt
lRAQKAb2B8ADJHOvck/0X9Lv9hE55F34pi6TLU2rP2HjCxGydYBU1DpP3wC0KeHr
3W1LfGhtcaO5tqIvSY6IxewyHo4toWXGbL+72fhhPz3JqEQpmnJpDfKfazPADwmQ
o5wYMYmloYc2VSSi3bkHjmd8crC6qK06EYch9awyHAGQlplwI0bRNRwaUfNtda3F
9jLOpeKUkBbo4nRvH+ia2CC3sxXgs9J+OQ5J43y5xSUo2sNVjEZvBwU42Gu1yRZ0
WpXYFmSam9p6+9FL/MC4ykEgzNFvfGtBoQAxTEdY4o7WO3nO7C5MDwT/qVLOsk38
GA8MtESL3JdFDsU/S2diY+U+3P8Qrl+NGFH9eBEqglrtILFIsTlKfBDQ2VSPTwLO
PJFdvBi0HnLY+qutTzz2gRdhjI8Z91eZUzQ3bzWYWRtWSq5RbnwqEKYr/PUu6EVp
2JswouqumjzaViycT76vlfMJz4rjvWQYBQ77uVLgcgvsjF7JiWtHmokzpf1RjiWO
BPCaVLk/SwNPUZwJVS7Y+U3S78XvPgmDkZz5TU8SObIMC445P255AoZbdmu2LIOM
RJCVKqTSnO2JICzDGQbFYk9aX3RChs0hH8PDjxM4EtLVqFMc27x9tk22QuNERI1x
VSikXliuOXz9ISOKDZrsWYUVcIrSAH/CDyaPutYNBPQvq05ZHjMZN/tMRhmjY49k
Fkk+P+m2DcuoE8qL5ktlUwn2zasRXzfM/iCkFAldgRLl7m1J/gkWRXc42Oz3oXnb
2X2ilqDYwPDayZo8+9nTRzrjjiP7G+0UgbXVpXFrde6M6aj6Zpbjdl/gR/KZVlk4
VTw1JIqhOxMJf7U874qNtEqekm5JEgsb54we7OvNF2kFLOtLHDIYykH6T/5U4F8Y
ZKdRN3xVytxDmiYR6NO6Z6ladzzv+upV/buX5lIJCZ7+XbZ3JnWZGaELSAbk/ujc
2yh2z7qelCUfbtO4n9ZBPDaSB4DESEDrLB8RA6Q3VlQ+w9APpsw8f3BVmpywtjff
PgUOG7wXPKxplstLvpnmvo04wg1+px3nxm09fHq//ncsFoFHSjol35hpiONQvB2Q
EAyAB/32urYpLs78k5SH2ilGYJOU7PtnhCaloZCoMXn2ptXjugmyS5VId5uFwNvu
ZWxVkJSMBfmsSvt9+lk82Tx/IUE22ixypjNH7r471hu1YY0/1926ZweQN+MOxVdN
iA+6qNvkiAKzpeoMQ8N50siSpZGXLfZBU5yfciiqAwpghAnBnCra27MT4zyzjaAy
FFTXmG5mWks8VHkdOluRzLsD2NFcdwNegt/+NqxxP0PkATmX7Go4v8hjk8VSy7Np
nM/KHjzfHMQr63Lai+N1/qiGKR3lQScZ3wCfK8YyEmKib/vNOhKdZxhPwbW27Sbt
xE/ZunxNH7stvnyeTPYRI2ubdwOs708bwKc7rU4ReKGfNJiTX3F15ghjMakAr2s2
kGDF8xD6mAKHmEQtu6oEezmiPSof16g7oOP5BUc3qa4cptESnfIvrNFYhojgwPWR
ASF3qrIGybllF+ScOXNKCxXntPO1UdwEDhjgnTdaXKbEYFV/dji4qsnObfCRv6cS
cssCVx8TTc8GgQSl4nBeOFXg+W0KxZKmcSDi04mVpuaw1gPonmxY8EWsWZlGQwNe
yRQga4WwrNcuYwQjtUXv2IjuJPtJtvdHImO1PlbuK0VjWjrehsN2nOrYjo8kSMZ4
YpytFl2P5VVogtTC6oqXXjWC3++RtcSNhKaq2PaB1We0GqCHJVFrfXnk3EwuJb1R
+zcGpC59o8qNg3DWZirSimdP8+C/JI2KdFteZodkRRWxXB0Jb+gXjHTmvdQC1tKG
IhHnfOc4rsoSlEJ9Bo33Gg==
`protect END_PROTECTED
