`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5q/boqO5OkUlKmCk4YdxDGV3ph9F75QjPG4vZbotnZmglZ5ahJ+36U+1232vJqka
K30TlCPoIWd72OTzra9G15Cxf9cdHXwdJcM7pYTZEbPdqtCBgcqFuyDNyreqQgf0
EQr4fctHRcgLOQML4NtTdQJzYhH6UHwnfvDgpav8/SBqK5BEF/pOk1bB07DiBMqv
ea6K53FZKs+wQWe0K4CyEXsbRhNj/PBHw70KY1Cs7L8Aw/Lc95Mc3tSpqoUQyQeF
ueo6WNB7ILjmdEwKsQnlxGexpAFplCaWbKQ9QvdVyTkpJBcNT/ANIemTp8kgHttx
KJ85UB6FtGnvhm14wtD30Et/gjK6MLyjLqOB8wegVuW7YCmhSxJy9fyB/n4slTQg
3bZTlLz7t4izE2t2Kpf/ABbVzeDR0554yRtLRC+kVdRx7IWi4ie7nbmGpncg+neA
jGZcA6MSavk+XhJgaleWEpfYSOAgtFLjigTkx59brRwKX8pe+Tqxlg5C+oAbVPXt
mBi3L6YKqbhp1ohqnVGF1uFdW51fXQcGoMLIcoMVEL4Rqg8KURuG8f1r9HRM1dQP
nsK2ChzpdgCi1K5UDUnObosx/wNbBdBUbvZSBev8IyprgeX1JPoN7lCea8HtQcLS
gRXLI5+HHBIclZ81Kg9JrCCbvONkiEKVL+NzCsCW+Hm19k/XfoDhxpVP8lPxXRO6
//v6B2WbvTjGJSnUV2O1rahU7OBtj/kyhBeyqa88MZhkaHnJEYzr6Aa9I6KtPHSn
vEqrluzgpDNuBYzAFuedNK6DwhqlMOGrnHlIU3JETsv5i/IbQpCkAVMzw8qhgmQp
v+8r/UjvPjlpsOJMlT2hKeHmulacsTBFLXwJAToNSR6p9UzrTYC0MuWInRmHm+G7
297goIKrOSrjqJgS2jBFSvgGatsaHJkV65BuLkm0p9lD5pJH9nPDX6kcpDmUTl2x
mfl6XB7p47x+CdyRUV2RR0sIQjexAye+Yw6BhFy0Qfw+AiGRTr02esq5Mc10LriH
YCSXU+N1q7bChFvPj88DXpUgEFbAPmcA+dFMY+F0+0E=
`protect END_PROTECTED
