`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iupo7Q7n9pF9Nx3u6dXsOWUU8rpGVN9cn1vbeIV99eDVdXiWIPzpO5zRgfzGwnbi
AVpBvYEUYXQARolKPaMWd3qPg2e/ChlLjohyF4uEnuYYsKBXAA5YW4PDan7wwfOy
74WMjlNIk4LeqTWNQ6Pl8muBxxipSv2bgU+8ScXojxB4H68/uQbJh+Mr7QJNQAOP
nDKtpxavxUMQLWKOnT77AYOmsCZ5Z4S1OJqAzqh019xhqDwlgAKVyhST7rm4cVVi
o4RKNYLlXqCBd9zPLUFFiFFsX3lzXFZuKqbKddbrq4tUNxY/AfD7E6Wy1EFBGWXF
7OKJ7md5/FAQQKQYTuL0M3sgCKgIPLVK9QFFFe2tAJiuPug22Q/TS24N0skkV1fi
VoBDJO54+TFX3DGs8XN8ELb3Py8R0MmEebnPFhWMUmfW8PtAi29tG0wzf1TKJcuB
OszDUililtlYktDSTkjuxflyNJgDi0kwFuLVCG94nQ5WOHCKaFl4ZlnZO4s/nWhf
f+IYZaf8jsA2nE71gOq3RiBmDkbiuE+obzf7ZcyQubtOePakSLUFu8j/mlkM7XCI
NV8RliUDdM+YETQIW1rosVMF8huDM/St3zihuN+S5oaLetkQs/ZPdo8lQ3+kysuR
xUl+KY+mJ0w5yRYMMoTUli6oAHGE4+CLy+SoNwS5B2b2KIxSyFz+7Fb8JmQDtIRX
6rZEwl0sxAYvHO2l9NBiLO0I/e6JHd3BTQ/OLkJAUTEpzOioEeUGAwaAti3OkAKi
VWo1sbx4Q9wn4u0O5lJXzlNpEIRkmWs+Ndj6OL7F3HDqDmg4k7OaKWOK3GdKnmjL
zfs0LzO9qhqfi/38+vql7BOOf/Gdjha4ApsMfNOzSyl4jyneHhDzauevUGhjn1hV
eABeoN1YSvfzjFqXb59KngvpJOXoqdzehcHWJMqbxVukrYNpEQo9qXyT/PkViHF3
IeMxPVhSb6+lBIodn6ThCvhArI09we/m0b/tb/rXrTocTvtgrsL7c2kiUQTWMoE1
XQytQHu0qrZLIFq6PFsntltZjay0PkK6xEP+wyUhljYr6waEYjGtSkOh//VLQZmx
Z9U7+AUE3PB5ezO6Z5cynYuG6FpECSUh+raJVavdKA8eUfziDzRjLTu8TpPkU5nR
Z2//mR9xzDA8GLVAEBpGRLVWdOsMGb6oqHatOgtivVplMLeLEEcJ3IXMkqnmlDPf
8QoJzm2B2KuFXSRxgxvowXw7iMAWtmuPuzQp3aXlCrA6HUyb3udVz+AhtCvbf3zX
YTaT/QJeVnGT340+1NkHog==
`protect END_PROTECTED
