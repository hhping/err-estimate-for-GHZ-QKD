`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcBmf+W6NOSLHRZueE1JTEFB6RU72eblxlpWO+q14yhmEzlfJwleKZGs067ZIEAx
KgmHHdEyU+gG56dV4E+i7HJbJ9zdMaodzwzxkXjk1rAXaCea32/om6jJRpiTwMwz
d6WrPNJpmOlxVt0O7vBuIbbx21Vh/IGabgiBGJ0177SIyTR2W2NQsdV+tjrym5q7
ogcKJsOUcWnWp/ERwFO063MOX7Z0SzrTJMe0TssmB7TCbHKKF9PL+CAvHblAiM6U
p120Ac7EeQ78/XkeILRQ5Dp1bSAmvWKa3xwBc5QU3viOx73W2/GE0F/gEJ0DCIp8
tGPvCaS5XqSbBwtCXpp4iRwpbyU8IRwhSwpQTxJv9bsVk1SlCkQRfNc0TcvG2yHX
4OBNlOWJJj8441Wg2bOal3eeQsv1oh49AtDw+zsDdAmdd4ruSZ0EantxC5MbqXhM
SVZu3d8kLslSkLHB1Pi+7VLeSxnPDRm2p6IIoozKZEWy6cuc3Rku7ZZrOYJFL1on
7cjnuI2DIGxwhHOBfCBvXK/Ae292X+wIVPovbmK8QsnWA3lB5hwSmlb3zbAbC8Ye
AuKeQ/nULwwmjMYzoEQZqg==
`protect END_PROTECTED
