`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNBObH5/ErpgdaB4XMaK6xJGneF+WncZyMxnLboGCWNU5DaLfKtK++ObUGady3Ma
nWNUga1FZaTpSnu/YmHdbUKR0XOPwHvoZg7HOltEYz2r31BEpXniepgzg1yrrJF5
Z3GU94KAvTDBq7TgyiIPu/lxx8NRS7joDh+EUC3upNU2oIt20KZe7LyiUHr8J7QI
p1YpVIq+hh2TimrzMKAzQSZf6XO0BzN688CLMMP2n4A/oe6Iun/fRpgn0cdCn1Gr
1R6Ky2hxdSAdj9daEyGY7YEIlRbqPBHe67qxetO/m0Wh2M52HQSkcoQcgXYLo26O
CIf38vMv5lMFedLypdNqchhReHIpoPcYKX2+5vclJLb17WVGKrspCgrXFUUiS4+7
JMmqwV3WE90cjQG/xbNsext4/ir/0cwc7tLUsl7lShadH/5rnkuBPDDFmhxPLeTR
DVYjfa0ZvhNOA3kwH052bYXtVbdxCxVXyiW2GjMUph8VrPFn9R4kWMMYZv/yr+6f
ekw1xSSadifVo7wZasJ4be017mF+GNx0efeLfVvYlxVqTinIdxE1vpLN2iXWiRFU
AO7RIaeWIPrXhjm+CvoPBFN4kSmktnhD+pTPrGs0sTy2RwTQeS+OeHca5VpYXODH
gZfPpEw+UM5PTnQb0cSfuH7nXLDC59DXYdW5sEqzwr36T5KTDpx5ShLCC8a3oNdj
4OdNdpfS7Ai20t1yfpBQku9f1Y3RaHrH4VfVtxYN6TRK8zJh4PEtqkuFo8a38ZKa
4epdtMj/X8jnD96un2rup5DOFebrwpuug7G0DpR54ts3QvIef81j6YK/wZ8ASg/A
mo5a9FKk4rAcTXlnNVFlT+KjlttSNSI0eAQYyJDL+PX44JaRqITO/y9k8kbXDPsa
rW81pTwhOseX8vlMmNDffzArH13ztlO10tuHzvrscb0eP3uE3v/ZTg6GmvEFEjpE
KDDL1i6VCVDGFgzi1VtNOgyOoBCmBbkJQdnVE3/30B2I7ZHR3RRRtG5D2gIRU+TI
QQRcagkyPhRmCWpWum6VOyiZwB2Oh6aDWatxoxzJEkHMWoQdH4lk3o7MhEKd95B7
vwMsT8kQJk/HQ8c+u+C1ZBOxbok6Ewzu1EGh5IptA9VBLfS9C+sRcleYRJl9Tdq2
tEUcs1g6fh/+yEVUoyV/CzhkvXQrgh+p6G/rZZrbT5DwlQ6AuudfVcuCV8KaCBe3
Am4aKTIyPzbNinacajZb9fj7ze500uE/t3pgFO3AW7+spNMKkYUVKnGLwdu5oGok
9yypLkgewTjSoEcXFyjzJjRrDVFrdFAI2PhNP8RoYd8xGnQmcjcNsOzJO+zpHEKA
guanyNg/JMfzasbxqR+yfbPpfd3kY5NpF50o/AZxBznxvp1KpvKrnsNEI5VqZb2Y
zxXQnCHw9zF6acy4/aax2pEWKc5HMtNPcwS0ttZanrVTiV74OSPwQAN1s2EmC258
9tNsopR/TiPYan/xOaY8jsXwVnPV4jtug7XQj6QfJKuD8tPy65+TYvTYXUBeFSy1
SWHwqDBWSTPndRYSK8s6pXEHkbyoLw6uwi8dJxaW/cAlcrvLY5F66hTEDe2rUnog
BEwfF7D5hIQbBYfBBSoVdfP3Q6VMm0odHS9NRXizIvAqsWCME7RIuRIjUWD8M6rC
U287MYoY50xyU3SXWHmvctNS8MfU7lT35S9n4BGvdcO9F0px5//e2YQPAX9XiIm6
g1nL7lDXVVJTcAqV+WORVpaGVwpAhKBkml0iTOK8UTJrEFRCnx3PeLwSQ1E90VIp
hBSjzoi+a17qZlu0Kt/W1Rs41no1y3fKnWD8b2bZQr4syKZbzxdk8uAvPPGB7We9
imjzV+8rOhFbeTxqNPtiHavFqSScHE2YP5r26y5FedGYmC/hWdU9SDUbYsL6vtNV
FBqaB9A0uzJc8geeNRJAD9WOc5WuJJVNtBKXJndG2ilMDe0FuvvtuosdUuIr5dQD
jh6oFdtAsKi/SLzEEUv/2z+vLPhmP0kRCi+EnJr29uV6rqnVgOt42vGDfhIT12WB
FVIrnZ6/BurIkkKrHYlLeXiKQ2Z8EFWUQkuHMuBZuPY2CCHg3MLWstqtH/o7xLnw
PK/B/nQeeRkvvO7QUaj0RR7WLQFX3mKz801GzYTbYxfLXQCNlvewmsBcye6o8xnO
MuyDUhQeiXQvwT0T+VKvyGAEZ6RnqgGwXtcdM2thVCgqxl9PcGwwf4q8X099Zwwg
ZnJg81lmDDdJ/uNLWgAaRXuC2ITWd1/l/6w7ITwGib65lHgvel80ck3eE+/OGePZ
a8w9P1TPGNXLNjSQb8AsxuH0dIXOODKZyqXOX/NHMlJgM97jIjcqe88PYyvm3r8q
oSuDSMkP0g2mSHvH+wsG5g==
`protect END_PROTECTED
