`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7Pre98MJGuLwoYv3MiHyEx+XpSh6Kwk0hvj1kTS8NfLcecxnGhSmc3Dcr5OjkgM
E1aHznxOu/Cux8PDBt1FEGWBhvG4eFDL2ARQqWRJ9J3zPN1QzuBurBEs6iw4KBag
qDQjZvSfkPqUbmHcVLQabYl/fJaPp00W1GLFydDnTt4EHECW1dLg0XyvfBEL6F0e
i2aNGerIVWJkdPj+pbQPTRbwLP2zOg8bDAyNjfvSP8YiV38RICoVbHPjAB1KeNxw
Q4PycxGWY6lwNAHsSlUUysbaxNlFmVFozSSxQL78haG6SVaYtceAtq6z9Y+GZxuq
rGSQPPmKiLVrAsszP5T3N2rno8Z+iQUTQIuFPIzrSzpm5hR/kx66LPwy0NgrqK0y
yjx4PJaI6a0LcxwgIW0yR2MN8/Y7XrygNTVjqIbJ+/AxDrqA3GqQFSKY1j+NYBrN
M+B573iwJL6l2hgmEQmfq9DilSx6vyFE10Ake+bh8aUfD3KLLh64YMJcabTVWJSj
IOxZUCZWKfs8AwxbcevecpTvU4nOzLBuUfXB6wbE7aCRKjkFZQi3nWyte0pCWdvn
oPmKU9QdBp3FElsFvqclCD3LbiJ/XIFItRGmSnDgExJp4OcZXbszEEIHnR9T8FKn
/qMhaBdCPFk+TlY+9a6q5LBzoMUZX0f2JbV0C6stSnjhAnE0kPVNdQ9euSp48lJs
IOr3LW4Kea5pG9yzBHw4CAycsdbgP79bN5QOsFOEc/DF6YvYW+TBVNzV1dd9AI4w
/bzIxARtOYtIzRtr31GboFR1h8hD8ZCXrbUWPJz0kQU+cSNymWGr347rT2IoRQSF
opBv+pKBawNSM8FhV7k5EMszsqDPdxjsPm+qEKrTQqJUmp7Rs3/Dtxr9ilIBew3a
SC5rqXwGkp5ty8OrQ8KVBB/C2qA7HiKBwOrNo40Apsr2USZxJQpdhgelxNJABLN6
XT41Nqd+ROV7XNzoPoZdaSqK2dZY/+M6RIR36rNdpVmG/mUA7GuLfDayeQi4spkr
qsBq8OVXWiqQEMiK0leeHPmjZulU/GfjH0Inukzyq12+UHRMrPkVg+sv6lj/uAQz
yAXXcWzoeJtagH3q07CcF5l8JKihfdCw0/TJWj+Wd/QmYpLEjtrSW9WqG/XgizyE
Dhvx/MA3ypV1O7GxoUnj9mQCF/CILAds/PYqtJFXXYPSqwpXfrTubiWgqCcEeRk8
Rbpqx2Zp3Miv9Xtla1XqK09jaU2KMlQO6Xcjao5Bf+n9LJqmL39OITqheQ9cpUwU
4TnsC8g1LcU4bN4WY9My/aO2X2wIhC73MBSR2YzBFnKD4f1++bbS9djIN382eY48
/1x2PimpnPccPE3+uyElF6oYkS7sA6Fja4MbFCFV4KI+FlaNHwJMk2rIipcCDgZc
cooDhg2lD/gHB6qXcUcEbgsuUqXq2UHxkahN/XGPt5khNVRxn5zgANF3D3pTtsD5
WIt1bSLw9uFOTjEo5lyH2iwk/QMgF0GPrE2R0LyGzHYumnY8umjzsiH2qXmBYclR
t1R18oqo5DjbkszcrFbCnZDKegQk2R11BMhN9FbjZNzKdkUHpNVvJIA7bZ+DndQs
Y0DVmvWf4N2i1SiXuU/mKqNIsn/oDeLTRfGpidRLr2Jy4L/SsDjZZszxe6VyhPmJ
YrtRsUp1KMS4S6OqreWHF7DDBhGtjYATNqGHK7E1Gxgo5rDRt8ngiNRfFaJsaTOk
v2Mq1j/Qa3aGS47g8dgvIN0RkbNObwD+xom44V7utokE8T1wbO+ln4diGoIAmyOH
QJmqUzKuMOJIilN3Ae1BBSAMA+/PIwulS2DCg5PNUjpY0fBdwSQev+3k32pwa3ql
atn8+qz5zGRp1Yy5lPE7FcFElADS6kXlzH3VqrqEQOnXtEduPtk/RIPbjp7mXo5q
R8EBsb3O4GY/wPiEdPI3vz/yyQIL4c4agljJHGG0irZyIg/k+kI77qVFCwUUBZzZ
Jbq5MqOCquzVASQkEHJirSPxgvmBQz+zG5A6yeOXsmevZ48mEtbipSWDatMi13fG
MhJhmmWwUsVQpWG5k4LWD23OBE1tPec6mpvp4DmFVmC6BGiZ+UJXywpJ/EJfNtke
CLjkWfYgz0P+R2mR9M14xBSj8aUicu0IuXDy0q7Q1gohxC0EewOGN5kewX/ydq+7
QMEnoiOQFCcbzSBilQCUMW9XmEPFQukL4GPzl5QbnBKS65p2rO7C+9OOu5OFrJpO
/MwJb9a6MeCz+WUrDvgAVJLbTEMOL0nIkhSkSTycIRjDWlHfbBj4MwGuqc8o4Y72
dKffuv+SXI9hOG/UMWkk41DPj96J1gilipGXtGG+qJ2OuTAbiPy1r/xfMq0Pzhho
DyPvocNreDCN35hAWLZSRrZUBIeKjxTqZ+sSHxz0h0nwlRlDbtk+I0eU1lOk02OX
hsJirrJQ9cFLzzkunhoKQRGZsMuHsUDbR+WK/00gG/qUWkvoV8PuImwJ4hxVCWE3
5iBX+4f6UsRk0iEUdbssuo+Mbrr4wcR4dPfEsGfEVxGX+4Fi/V6KicUCsH3O1u4v
gYKxCgJK/QybsY7OpyKYAlpz5eWMB3ZU6KhIvsu1Ej3TN2cYP2m8xu92pTCmYbRH
mXNuy0KbxqR2gDl8nuAeYzZ554b2IlyfKNUfYSi66dmjgSCuPFEA9mN4nFmBPP2c
`protect END_PROTECTED
