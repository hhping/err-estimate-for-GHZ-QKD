`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Idbw54eQzKztgSpsmlQBC1B8tvCFgIRQYb3t37IBFh5vU3hRPOHI4w791QLc1q+q
5mb2ZRbJHTd6L5MDgqIX3An5iK28gNt8CkOJvxarWVCZAMLp4lbLhCdbnL8iQMuU
L2HA2918kJIyPB8EMqiG/tEmrFeUQoPF7G7pYIGli2IieOFMZHf8RXGd7IXgT8PK
1+FzA3R/mHDUQTGfbk3dlfFRxAtbz38Lnlam/4VZVrbaU/2EvugHbbvlmIwHo4hc
SurHunVcHRNqPmS6WK6zK4WbIynCfkkePm8O2bIIf6FnAoQPLEPYR52jUShp3Xak
XxjZT6f9fCHc/5Bd7McMrJmW2QWAq2GgKW/gTjJ9ydRyqSwhsGK3rKer4XZG7R3q
OU6v+IubOp2nL5hQFYCCdQ==
`protect END_PROTECTED
