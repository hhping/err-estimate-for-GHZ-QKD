`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
771QAvhKLXDxR0R7bl3+Rwro4DEd3TgsE2KHv6Xrb//z93ziuhhJDgDj22scxhUj
e35JAOpAi5RhIf7eW/pTEFY6B4TAjIaBXl2KxwHYfi/hinOq9laOxqElp/OMXw36
JP3J91VgkdkNWNms+UCRjHRIZwYvtf0JCrk/4vrznza0Wj8a7Msz/m8wwn4hbjbJ
u8K1NP16QM4bnYByUZdzWOdxh+GIZQ3sK379W9/mvPgHP5mSBCoTE6/6SFqvbuCM
zHu8fz5hiP2UpZGQGJgB564QR/A2xomabdjAVG+ZLok7kTcyFxtlAjIWutok3lal
vvI0tTHMF5Y9nZpQuxZMRMAtL49VqDW5Do0wAWDTgDJ3+o6WG0uHD+5/ARuzJVF5
nF1L+59XWTBqo+UCi72aKlc8lFmMWY8JzlwzXTRExzniigpVnfHD4U0XdczSGb1C
lWtmccVxPhzpuIJRljM8ejTUgtZeHL+v1fcdU6FGp7KTfSeYPpXg3QCdZqbpYZxS
2/p83Zz0Z98F2c1KOVebLLTLueWviq/aFS9GSDwSmapiztta2MHErQOMawB9wSEH
`protect END_PROTECTED
