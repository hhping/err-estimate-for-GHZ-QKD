`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbNfbiQRv8zNdGxKRQgy8mtXnFD8xGdE1SmX29XUqx+wFnVfe46VI+Gx8bhvjoI9
XpfNlgEyG/PBG/KWc65DMdwf3oDD+bxnTY2IeK3cCAECDBqioI5lF+IYI7plepVM
kh/ilrFEKPCn9Ydj11f/aSffj4pzciTwiTJn6yG5cSLQcvP8ltQVKsQWr6YvTQ8S
eHd2oJXcDgA6aMB1r5zowbaRPct/L16A0lliw6DJTVMnFNqh+fr22FhVbo5ODP5w
YWr6MnkZ5OQcWgGY8ALF5kvWmo1tgaej4sncV6L+Kt4/JRrjzKLs2PvzgkPc+YMm
JqKpSeJWYMl8Mg1twiY9D5af3TLON3TGA34Vimusoz+4pQggLK2f8fAJZrTUmLsf
+bpg9NPTNgFuV9MjXh069HALEmS7i2sJ/g4TGPVsEWF307pDB97M1b5I4fCvnxZv
eHNB8tK3DScsjUImrue4PGcWW5KLC9D84v5us2BlnwfkzDocirkSYCldEaUNhW1X
aD+7d26Z7MKyzj2+dxDtbRZwT/ogkiJpgZ/CWv1C3qFpKeSw2m5dXSLR1WiI9ku3
H4XMgAfHt61cseDUzQcvp2XPnF8MA8OhVXkmDfCPzHmQki+rIGPSqlz8JKQjgFlO
EDSxJ8k4PYMaCM0+380nV++8a+gAAqAzMk/Q6jVM0G02TrHGs+aQBWuB2pOXQamF
6EM+RSfYbmGqq3hwpgz7uBkLm9WZQO4orQ0IgGiAej2bYbVXKzYdR6HqbVD0W3K3
zQNy424EmcX3S3fd+zppH1DY8BxvoxsTrMmqhaoTooYhmAAENpeMea09KRdbhFQP
aMr+N6DI01R0OSDOJr/3X+bP8aFVXl4LQrZuPpmc5+lZS0cqVAfQx3/hu5zWHxJ5
rq03cDPvZVWaAu78MfoLMH66ihdLU8JVsQXHorYhaj8=
`protect END_PROTECTED
