`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wk5ZRM8OlNRxmbGQAoOW4lxPrJVBWuHYRz9e3NCFYWc435uz1K692J8eDKbu3ZyB
yCRwBvTKkZOEor5Qc1ZxT5cIip67aqPgYA2SYXx8huRatO5g1YPMhfYjlFh5PuK9
Q/3EpOGA40Lv5T7gSOFCUS3R1aSHpwMp2osbNZG/GKx2fnKbZCgIS0hS1iORKFn8
NwmUBRkKuvpPSkcy/Hgg7sFF7xWn1aKdLaOEgS0GfOgYm09FgxusgCZnEFBp19pq
2odB81iXmUOpIdiosVkf9vtlQluenhmUWh25vVUXlijlYZRzHwsoo6osU73MWU3g
6LxbvVeP8XHv6NBRVpODy9eBw6xz8BRRHDctOWNUWhXQbVmWgxz8l1VUEVOkQrSC
XAuIoVgG8ybM5uTcbFfommh3m9WyYu9o/CPn2smpG6dsHfe0bHlZix3vdrymscfj
rn4X3vy3Dql3w0BGs8IJrA6ZIEQu+IdyKyqwl99IHD+VszMe9C9xDzBjnyPO0lTy
TJyHC9I62pOgWlavJS2ER8wsM/mdl54gx2ASJutEWgW80cNdNc8ibHYpsVHBRrvl
5ftWQIouzLvqVL5OWklSzo8cD2dj4E89ZIYFk7Rs8MJukRIy25oObIe3sB92VccP
s3dt/R4NFFrwsS5MNVvDB7ri9EzjBUW7o12ZstbKpA/1udytEjDEAuEsSGVCNfFg
/m3WI7T8ZTkiBBux+ER+7w==
`protect END_PROTECTED
