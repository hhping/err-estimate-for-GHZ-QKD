`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZMtN1EUX8MT/1Ys4vhWlmcBzLVZa4b3NCDaVUtzIMYE7fWf00n6iHjrzxmkrbdN
NLAQ7Dx3oPgkcAM9vjuE/39z+t3TXwB4f6Kuy9HHxUZr2iC9H7dEQaphUC3X/Cmp
WD4uOr4LdVZuGHzyC6Z6S7ZD97atB1cvmcEoZu2CjEBcvzUlfgAQhoK4187YO/8X
zF0oI6cAJroSF9f/cpqkWWLqYBP0ms2rZMOUoYBPDNPD0SqvAT+YyBpX2KJPJU5B
xjL3oAv3wcBedHoWlv65efFIt/0Wd58JD6fr6qHTUVo2grbb6jMAwAgb/m23BpzR
aROuP19z3rXTajSEyi8J8y22wRWr7IUE61a7AFn0sl9G/3a4IeLCaNHQAVSkl5KF
Kp2jpnpWI3kKq/NOX00cMHr1+PzD2fGqLT0nTWFZV/piLYNczB6ZrlaAwF2HWqZu
qK8a79y/at5JWtV5DXINZUQJrlT+vs/ceNg2Qs3NqHWoqeUHJrZO4ynwD4il/R3R
caU5GZJyLzTo9TmmPP+s6Z5VEFOlK3yclY1hse0gEftx/EWiu0VjLtLOURw8tnYu
YfWFwANxp1WPba6CJFxS5GX46PEadJnY6VmLfr6MvpwVemA9kYWEYu7lgttegvku
W6OmsFQzBVsEv4oRoX2wChbGPbg0L0VGIBn0qoosL/I=
`protect END_PROTECTED
