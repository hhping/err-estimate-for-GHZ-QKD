`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qqYnm1mksHiZbwt2eiz1ee8Z2C876mAtVAtUkaKYBxmHSJDiZpVSqP19ecMK5r4
RJDf2xhxFgxjaVszRESN6dqMZ40TVnwHL9SQZ0t5hyw8ucAh0uUF3jNMvvf7KQ+v
aWPm7IdG1267ZfDRpBkOYrJIhPkg2J7LmyG61C8oKlEXmtyLp3QK+WJr2n/2v7jY
+hqdCqmzaykPglyThrFWumtPNEBYsksXRAIsRyIgat2/kLgPpSGRat7zS+jZtZeD
iupxBpLq7dx9eb3ofB1zQW4vVX8lr3z5PlAGLhSsEYOcfN6FPTY2W32SpMgUgand
4zjgYnQPIe4GO7sPsMCnAi8oqGKTPp6vS5R6SeGTfQcfU+Ir/PPlXG9253FRUXV3
hyMxIusV6ywNXaV77IVRuo98ygeXMApVhU/xqDyXnQMF5KymAlKzesOFnCKAXA0Y
wf/fN62SAm7U7va4gS8/Gwph5cgGp0p6kF4Mod4lie85ZOqq8fA7mQ4jMtYsMVT0
qV6qCk22ojwCS+3FJ4dl094pRoa1AmJ32mmvmznhc98KdT4zlI4QYJd8emVMCO58
NVStTMCXKEGRpO14u7kLE2VPx1MLZPGsPgyy+6iHOH66/TmMxKn6eK8qj/C45NAb
FQ7NZW3jRvLKrE7v2HUWWPQ2YEHRW50AbbfrSSEz1Pm472AST0wi/hoHkIAvvpza
PL1zSta5wruJQtAdgv/imVRSHlGeBQrQXnqwBuQ4OVpRV6ebl6KVNCcLZhw2bUFh
wHJ9OE6bptlmXvGPQmD12cXxze9z98PiRCfkHz8/HQ5V5QngzXj+iD6N+oCSiwY6
4zFYuz7zfM2NX6aznBCM9k2QPoW4lUD4UZ2YRKr0eaKE1Yv6nfZs74gjlTss7glp
ick2lhUzvOyFfh6ionknBAVrADp07JPVc4gvLdAXc7mC3kTpMpJt9IQNh7Osz8G0
gP5mYXGIMeW28xyZeYbCUCFynuSOeFTGNUOFZrmUVjNevo3ie0Ie1WH5u+UwSOSy
WRaBVD5/cL8OsoIb2ooPe1LbmJCaoWnv0PI1gKdB/9vDXJ2swaM4REa/s9MYNzT4
oFHt92bYdBVBUpG1DWMC1x4tbGpEHAtZUudIeW6g9knyyKPqdwtaLsDUhsj4CHrv
TX2isCcpPXmmfPKG8DfbJ9xDKcG4QnrPuxXxjZQJoiTa598Rb3md7i0xtPkVLIxN
owvK3woiq78goVZXj1Q21tBnwq1O6+Ba2h83jGAG7SsQLx9TY8F4j4xWJox1IBgK
JgM9CRtiB4u6ywVOYbwm24hvjLRazIhBL6XKO6Hw6dnQn9zj1yKdIxzTX692v04C
cBYpwXG4iZYw22eIb+iTUaYzaQ4/BfmaUPpeoPmh7kJH3XhiZPNcV0vuV2RTYYg5
Mua6sJqt+50vDhKHwy2Fsxocf+8HdwexX6QQBTWJhno+dhkzlLP4lY8emEPoXeqL
0gSolgMZWVf26ebFj8JDONFpB/CLb0dRt8U95JtoPbHDhON/y3XsuN2WVG2n6o5g
WJRWTQO9pHcjHzAaMIaPs4dR7WPUCdY/4l4lxxcMHxPJSyn4beod9BRNUZQsBQKB
yL1MYURuezmAeGND0lgARF5sVfF2eBYGLmxQJ6K/Rz9t5sI7TXrsQi/qMlC8GB6j
3rbnRXTTYuR4vYjI4GcBhvyjoxhaoBOBsKuzzqiXRP0ib42KmXOvUdKVTcdMjzDS
4ExqSD5iWkuPu+ZQJXge7per0p+Qfrr37gp5akjhupAitTrr4b9rOdyW6VQ1zbPn
g5Mm3CNbSf34JWTXez06NYMMfzZGIcZ44A+7+4e/VCjogWeQCpGz5XrabwPE1Pve
DsnmAzA8yFjRuH6lh69UFxMmlj5l0vczaFn1LZZg33ZHyGtqAt6YcnA8Wpv6hEad
CisvAFcwoFtAyBWXXKO05sy44vqZRJ0k63CGJWo9YwqnOzzV26Hbo6JhQ25jf0S9
pFm8G3F4Hn6ALhMUK22fvJGk7HZU5mBuJqftGvtJjRFZN+77VqbyfozkUJpn7s/Z
+QRvYG5kAZZ2EaDOyiYUnyQl3ExVAXfy+4aerIgdtJnSGbFdTQfVUeaOFu/NCERt
gExnZd86RKtMHbTGcAoeZ0u/lg8CTGZ7KZkbuiS2jmpQuwOZc/81oFqReUXYrKYe
SGhH8OC4ONon1yl82iGLzA66qSg0XJ7vluNka5XGQIxnvxt0RtTiyjPNLJGIVw5D
NPLtigGImjcUNu2X2TvXQbwSfUlY4eh8GHSAtguAwEiZivA0ZU+iQigO+Z0Wo/U+
4gNrr7kj1WxSWXx+6ynWQ6vyb7LWMLC8cKAPiGB81a8PDbZ6/+YEUFBtbXJToiUN
OdUwtIdW2Rrp8eI3KxB+oTDFChH8crnmjpa4/oDkCrh7FSE44jA9FdbtHHwgvdoG
/As4pFAqK160IA1LIrFxU+91ow/C6B2Pr3Ar0MrGPKrnqG9/kS8xMSe/M1mfGvTh
A4EAKM2ilIDzUWy+gDOlFaeev0yt2fBDFjfdK62YjUfcqBmVstEMHdaSoy2k6Ilk
qn/WwMDjfSUVfO962R+n65oKycKFsZchYNpPcEvZ16kJPVKJ3PLaY1Lj3V98jF22
Jrtd8qXv7A1eiRhbz1WLTKDpxFwCA6646HpOVLH5gKMWVrX+wJyl3thoqVfcQTrf
ib18A0w+9Ppqd6BKhFbIpTOWFToxOEdP5QV+2lN6Z6mpvvAP8HX3u38AL4OgAh5J
wjlqTFLIysJfWnAdSESP91Dq6YDASwVsZ95CL2736x3uw5sShDtIl7VCWYgyupQ5
RY3Q/OjDRWq96Bp6icCbYVuEciJ3EgllPTLkGWVL30du1A6lpiBT2lXHXxEG20RR
7nL5+BClxJJ1G6B7xNGi5eUxnxH8O8WFmYytmgJzz3L5qnNtlQ0JbUypTWrnH+Bi
/ZXvpzVE5iSlwqxIDd9mPLPtfxB/R4BBIVpTWlYjTG1gCGbpKjbCp0lQr5TPLclH
D0GhJFA35ljJHQEQW5HCrd742KBBEmaoIsdBG5Iu0uX+xYFOKBD34CAJZpCJ/qci
40Qa/xeixpxU3zLLneqh/4lQJR/wwdgRssgTxXFu40VrA4YFGa61FKesLw90dLhP
7vJdW3GCt9D2OsMABCSJ/HCfMdPlawbkg+4lL06660rXuLO1T8rW2QrmxJfrTIYd
OOIBzCHwBdEd+D2Lwy8iWCrHRMaHhzQREKz7ldtPYayMT/MhRCfdPPkR1QukUHo0
Ec4IYoeBgD1sBti9qZTDv480BOvb7TOTJHItTY78N9pCK5Fk4L/tl5UyW0jMs8CU
a6BDX7m555eoyhLG4hjr8hPQdbR2fAQzhAK3cm/IRPoMo2BUfa5ECi2UW1n30wK1
RNAO36oDAAE5+L8zc/5NtMiPYbqTx3l2/k0+0e6TxzHLO355a6WdNcyR32hPwlVF
oOGPMhCyqsgxpbyHZUmPGcXvBNwCAYcnwvRG6yrMC6ZO185ffV966gFG6XbfRj63
pkGCTZxKaLm54FWUsjsWlVUiYpqi/K08HGOu2dWfjf9bUyzkOqxJqlhZqRt95Xyl
`protect END_PROTECTED
