`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5zZEssbyIPKonCZ9pHvxn9kqJXJ9j71t8t1q8LXNiOuMvc82XoRzvD7P8whk8W8
3hjS3fEU99eouoqpzFw9rNrh/NzJQGJm1DFQjEsgRPWFHmsq93Iv3CFag28dbzbj
Bmwui8Imi6Z+NyTlHOegVWmr2lba/Z3F6E+wrYHiYt8vGGXdWLnujYsfAntVb4TS
qHIQoKNomdKT96GT4/j1QppeE3Xid2ex5XNnRnhGaenxmGuJ1IKLLzGPIvvXI09S
Eifl99XSDHn0bf8Sml11TWqxnz9Ynr8uCVWqMVVURoOYFxmEd4L5N7gqTNlrgtvu
39PMCmV/xGz8EJa8YDsNhDreiAwMsGI1yPwIIsgo9exY5XuaAv8rQrMLSSUNgjDX
3RuXt+ElevxhxO+BJ0YPUyOypabpF7QjPcnhOCQoY7b1vyD4hLtsHtLDawfgcGCJ
ClN29QQwQmC1yM1GGfymzUz7rrduYZWou4+kk3y754j8c4xb8XtbAqMc7i8vd7mI
mdaWKnA7G2dKPHC6+YpEwoVB8iHpxTZyPmAQgoudZWABJwEV86lnPukAZRVsQiig
u0SAE2G6C9qHTqhUWRjofIo5+8kSICbDmXqhR1qdWQzhs1OK5VgRgxhNapD3Zwn3
5n9fnTH0+wByTAAKQ2knYUFSszklMm8Cfh0cxBXgerhyX01p0ZJeMB2MYHrr8z46
rRNEXYQ9aFSRjhja+n6pTy4cxMLOAppCk7kgzaz43zV3CiuCgtAeBUIWIu2fNzK1
pts02Qb91hYbSGzhJAc1Fl8HZ7WiUXq3yVCEkn+m9fLln9o+CCPo5Vmtc0wUqmi1
TYvaH5aPKJAYM/24VVS2lpLvttI3uEtrS64uvxRrEPYE1H1gU7W3LVDkVLoi1yvG
n0orsFbr64tPtk+IA7il0yrysUVNld+1LI2J8p1CkME3KZbxQ1JPjzSAhRaPYqCQ
UYtAphV3ErSC6dWSaYO3XLBaU4IItEqkrItHrg2I8g4Rq2JqzonjmeGwnnaoHwIo
Pqdw/LahE2UtO1KJHr+Ou1f3FIAQYFDT9kfa+773ao4xqY7IPvnGpNh+XF95IpCQ
GdLI5NO3zVkFfGBFtW6rkNXSdG2JH6Uo95iUHlHagSMGlL1KWg37w98GsqPtPtIZ
d2g4XH1HaRMAm8MLicPTdpEn2ZoW4WbCoiciLHqimK4WFzHPeDu0igYxZnwnMeYF
Xn9RewWii7G+Xsgb7tsgTy2ckrw30fjixVfhnqE5WjjUodXNvdVREyIkq4TXLDPy
LqCovOnARW4qFdwQBzWypZEM/MBHVVaRPZ2QOScRiS9xvjOVvYsY6XnGDIsoxI/k
XiUBFfoi2NlRjKPdpiaq97yxv0tr8JPM9zdhvYkAvXUpngbha9p7iO/DPrjsVglb
6TT92kTr627dnnVOGfQ43437dUSILmk4JOHTvttoFzrHNrz9YkFWDmQmpyTpeRLe
hSKeJ7u/ihoVMf/KW1LC+kYl+6iWGeXsGFFgtyb8CjqHtCAmjMdiQ4YoI5zO7sAh
msbt46PJxldftS6tkeeY6H4UWMgbqKyIqcu2GotKqh8E+7M9R4lVFFkgSQVy7gPA
TmM7qMEWPRwei+tnvfckjWFK/xKjePITTCypP6QlZeq/m69EYeoVrXucW3mjFXzQ
fYiv06uUjK3Ywg/+NDThMzaLD5hCy67AA6D6hhrlV8JiO3gNKbc7sglmxQNzaEJU
B2bYjmh86SkxCOMCtvP6h9YNHz6YH0jk73MOZ4aARKP2eH128PfhBwhJlUqnpMc9
+TmLA8rHCQkr3jk+leu7pelMEFcO4qQyLSDrGnQzGKA0HqOKKFWC1DUnXpdhb3cH
pNFr/I72x+BaypLChK45IRpEGd7ViTZXQJTI9vMwjvH63xwhkqxJrnw02owsGC8f
35dYu1y80PCcFxoGuLPgS6CPzAUgWuCeo2yb1D6tM1LnN8FrCuOAC9tZOpV2UQby
4EPMbddCCJU/TQkDJ1Wn5VOtd4fNyy1VgNmE1pCSS7bYF+cpT5XcMVKjbuIy6AUi
GSSeqhCRk56SMXJeDfL2sARvdruYrt72r77HhGFdc/9lS/Up09g3Gu7JS82vEeFs
`protect END_PROTECTED
