`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yElLc5lQi+CXgp3qGOpOlvBL7g/JHa21G/y08o9awWQ0+fUn6mGudrJoMKJSFF7y
N17vPBvtse4aX9TToCeVqhAQVOZb3CjHGEL71aW+Hrsc6JO3zwEMUf2GTxqlmuEv
OiFbQuzmtSSuCKsNx/nX00Z6hZ7hVGCtktvgQ8nic4hm6JTJi3FERPMe3whVtey6
ncddUPvbsG+WMdax75vpnMH5v+jv5sHFcMvi+3WclhVa+bIZLghuW/xi4cJFLVEp
H79Ybsp3LSub9ZOGLj2/+KkvIBfu+T5NKtAUfInKq2nVlYmefUkuQwHGwsTMHJUW
Fi6RsfpYOfCGQ2+pMMuoLaYCWY2Zna30goSaUtRzWFav2fi1ni9DPOluyXGgYGke
trW/aXBUClk9RNhYsU/zCUkuGR22uwS3S7oRA6V8uFEVCkYFV1IhKUqrxNffbgbI
2bsW8eTfMk/1usVmhXxTkn8NMHJYc+3m5YIc55Z4Bei/rTLq/0YmQv/+mZ9eEaGZ
HCmOEtNFm4e5TUC3NEMtMa1mzBySUHrlhmEL1OBjRVYi9vOsibHzFJrh7XZro+Yn
r3SJ2BnGOpKIOiAxlA1N6aac6yVHzRlIA1jjWZ5iw5DBzP8tPsN/gI7lmNI/WVw0
B/BSQOUXSRgqb1D/37QNB6pwRX0sguOUjehjIXeIWdvmyiUo4oEOcHEWnIEhWJYw
PMOGoFzPx9fPlSabq0tdt7aILCrwhNkpP8J9isSyj1TpHy9fSqTn9H3W+awu0HW7
2vWPIfQsScpbLTCeLLOCnP55HAh5ilhbGs47x32Tq1D7Ut9HslcSZOEitm3Mtgwl
FgVCbmOGbrjtnadcNvtz4lE9JdEj42jcq/Bx0U1CAulcqIgmb7D8Ud3lLtMrGb8S
O0B5u6LxKHYN6mtVyy/VOR2pzPEBDUGUKqFU0RqDlv4RhqDldVjgdN0xCo+S9Fgj
7RinWUDPQmgdAeYRZq9Ps5XeTDEfL07DRuAcw7NgX9RPV95s8kJPsZpsjj+U0Ns2
kZ2piTf45mNFeYE72YfSMA==
`protect END_PROTECTED
