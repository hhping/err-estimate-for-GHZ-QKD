`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSulHpSQ3VWNL/jqt045Thx3663pQd8P10K/W1OEcN4ZIyPJ0Ns0NUaRBkNPEYF4
DAjgkh63NTKA3oA1S2ZI40HYORxwd9vk+3Yw8kP2T17nUr2V+KdKpBJmCxe84cwX
tBI1hT4y0TuxSgfNQhvATzAbdVfdH9WL4XPwC8tx62LfZn98i/0y0KgAxJE4Ip63
iwLrTLrBfVgg2OPx0D7TALP4NcCdOs40972n63ESdvFaj6Pps/LSteN8iw4m+CHv
ah/jk20GumVLKLUl4fC6EN/D0p9BYhxd1gzzBkeVwSU5AjuHYMayPh5Hs/RH1Otm
5gi/qqD4StS3kScr8Tqrq9S+mlApUEIa5IjcilpKmOhZl0F3k7pExZhohMKhKSJt
SzDwTv/bwJ9PtgN3wt16jhM/nyYv+llj/8C/i+aMKTV7rLoakbJEKAfovQbYZeHE
mJf3CRY4cRcgMBOsbwSq4JHq6NYAhg3cxtrIwdQW9oz/r3eELH/WrRgle9Pb0U34
h1mgSkTjKZGLdq40AlxbyhAfIi0q48Bmv6xLd429pwEEHTA94LRKxrhyokVNZa6k
PhXuNM2nzdCbayXIvuusUMy5/DAfoRWzOWjYy05jRF1jU1WpJxW7ZzRceEAsLJSw
R12vcg/4trwwZNXmlP6y+OfEeSZjp5p2gbe0UB9vTyFLQa9YgBJl558YJNa9EFHy
5JL+o07R/PUv6bQLQDS/Ly5EnZxHc9fRg2UPK3bW5AYPS+b335RtRELMtsBTZicd
lfb6DtBHsXjgm2bmFkcvFM4KQYNRrF7Nbxtzonh12S/L6VpAFIduORdC2LcYjfKe
oSGWtg7fQFIBaN3cfGRCRg8WzNXxZpl5RoDDmRmAUIxPmixVtNXKhS5jgU0BXx0i
jtYHZYrI2LRzQAxNkT4T4Kjvd1y3Lpkn7Gdak1U/xdLuJhbAnCgpmFIBpVIqt8Qw
piy+1k33hbo3oZfb9c4trGYgVKN9VQWWdADrr5+sh0+iEDKPmjE7/LodZ5AZt2tW
Bt5BjicrVkiFhxYEQCaYkGTY+GFrnMcj2hOtVAgHrIyWw+IK3xU457iB++08IfFh
va65hYCHqS5YMIJ1W7bns8JW3GeDLxA0QA+ANoICWbXE6ZGQ0n9nusuf0RFUaiPd
9ANiK39+qKYHf9vZkVTdgIVndUGBiErDyQOj1Dtb4bKC8E5NQq9WuuIbDLyR1JUk
tvejOVkYW3L1olxcjBzPjrBuFTcq+43SSsBGwN83kWuKBc9XRN86ZjV2F3xYgbBI
rzp8nSvr0UfgPiv86692mQotm/hBVCW0b1znOwaxrNpgXsc5FmyPZqjnFz62RMkr
pQlQXUpkrAmu7NvyRuzXXoeDSmcJao68782Mgvcv6LgLgcn5F5U4KD0ZnjwK/4Lo
3YNxWmTuOmeZjqeACL7pSuF7hhVZpJZLmk1j4LNIGRN2h6S37Q9G/C3AbADRuVwT
+vXHhSE6Q2Fmm5/JMck+wvyNztE2Vk4U/hVoySDfdeJUUrt4fzhrHgHamtcNBj1k
Oy5Jqdpfpwzq1QMYLKlDkNYmAqyysSPEdQzfOOqIT5sbWFZzRKPKBewL406Ae/mx
`protect END_PROTECTED
