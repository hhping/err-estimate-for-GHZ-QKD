`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HC4uuUDq8PUVujCkyKeWGlRIeVwoHKTQSOsLnsBmMGmcpkjxA1MV8U26Bug4mPyg
5w+AXaSKb1fOEMlQrEWC0MpYNZNHs2YmDNh36h10j3Yz80gdfF1OcXMAOqDoKfbc
2xdlpNkvXYtXSKQLuIGjNM/JWT/4UBNq6p7fAkjp2L6K2r7AvYSc/Q1r725zpLzO
SfH87D9duOu1bwTbHmFjfSXygt8AV1Xy+aJEuhuuUsuy2NaJZYlfBvjOVSFkQgzU
c5NFPnSCRXoL6PUIIzXJBohUUecneimWNin57AGqhsalJTseI1iYfvZrJ+zut5i+
msghWGoZICrEiyxv6VQiq0DdG2lUBr9ZxvATJaCzKGUTfrH13QejJeiumK9c35dE
7XIhMq4m2vuN0MgllYxS2ZO7wR+x+K5UxZoXoNzQo9oTEh1+DKFUnuR8CZryqwCH
OeUuOm4OEvTCPKGehfGTQeUQqqE50zcvgetLXudLSwOqoOyMaJ4qnDk8cxV6E/6/
rodOxy4e0Hy37zdC0ml90vwJnxBNscLvYvgg3nDuSrnTaF9V74uLbKu0E/aNydlV
6xaslI7tWxzHRDtUyjfBW2j6gQ3v3wZ5yJ/GexHp4jzmdBWsXCv0RkDSY6POMPFy
HvHQbmIZaAT0W9wC9Qp4rwXpZ9J6agyMappDcx3K4WeSQ2v7gIgEuht8XfNnYzz/
cAWNu6LzkwrayK6UE2Z571/uwfr7shOpzBFT3z4XyPJDbmV6YRBU2uVoFievGNPq
KO1+UByL7qHOdCsLpaw1fHw+4i9ckgCB6JCaj8aUzux7ipzK1GYDC3t6r8+QW4Jp
UFE7nq5A/TiiIXdAu/KaBwVcrwtiuo+VX+4uSiRkZFp4uQIEYlwMo8OXmDSg/GJn
hIfi0KoHlvNDF1J/pDwKv99bICR8q1QNd/Y6u7RRnJy6NcjgxF5y4BQVU2kA2hoR
W/T+HSB5mlGi18z2sTqFiHNoteK3P2wNNgjxM3QqPh0fgazPmqjXUU6i3ZSZ5CJV
`protect END_PROTECTED
