`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zI3KQOMD6FrEvJuVmXZv9t/zFRJadDheEu/1zdeZYeafTZcfu24H7noUyZWqSBjE
thPYwhWsvoQrhEHleB6Ofa9mLE2kn+ugpObvmEumgn3TzbAUIbhOlQIJGu++jkMP
a12oFFW3YnuvNZPTFd/buZCLjP4RUMMxD0UulWG+RX/qjopaPEtijFDZFWVk35Ah
LtHNhBq+RAT64gXpRqvF23irvlv2HLnaZmJD+PMRV6rWWQWs7coXta213I7Z2i96
eMJdyiU3iG4DgBxVeZeFF70xcRloigNnmTtTCvNolFsnUYUJ1nEkkczN13z3um+c
m4xwKYfIHUi6xgz7FycVVwbGd5PxczLZmtHhPXOP7qqtg/DA8HlDEJw4ycsNymjv
jmoDoCLsXVmILvC71AUU+1wNS0glgG1eBV1us6a3pvfAWHIeHA5FtvA9yCxwShQz
E8LYwRyU2ixBRACBbPQY5iRshewQ2emVxgNdqd8CIoTyzZUzlZRPabMK3qjuvaQ9
9J3zeCOtKoLFeeNe28UXeGQu1KBL/nrUKDXuA7jphOzwxtddYokIvtyDQhm5qfxS
NwxuL2er+UzwthyaA/hrB8GlBxnp5jEO9iSBv/DR9F2ecP1DzV9Hu1YgUXw+uzig
wIbNyJwgzlydQiWL3H9bhmOqL7upv1r+OHH0P64PjhrN0x22BCX7scQTJ4K0j5o6
tZKrooehW9UGy/tDM9wRO8elcv3iA3iOP71zTcltVfFrz+nCvX3PhYvrSe8QQnld
nJDMJqzM2ljK0NTGS9Va05LHAMPQ7eaed1o6rD1Wm/2fh2qECdstn6Unmn9KKs11
sGFoDqeIhwBzfTwv0L8kv/FeIA9lkKb4EEAlGx7NljnBkAmxtH+5oC4oWIlztNyd
AC7mKPl3vyEM/B+OYCFIZamhT/DpJeVa38FtH31BfGGWgUznGKc1C75PbfXe0sJo
fwZWA6a+sWosBEoZC+D1nTsqLgiNECdIQpUdEdEkIWOJQRRDKh6SdsHTvJwgIdix
IyOdlN3eFIJpzmBnKTPehNmpfTEF1WDqgkyx8SKMXbaRobWH0eaEKMijHZCPXus+
oSbdAcH9ZbG+9sgA6MS4Z8DyZ9b2UJho7CmEyHO/LyiGWAmBcxO4mi9+YjKQ9gi1
2ubWHXeZNIUylS+VzPrxKjlze1hpe3Vu9B17jfVu5/XAPpd15IKK4wn9AZOxlH4y
gdH1/mCiGZx6ubq2iUDmj7RWqrcm5eRjwt38yQsnWfwGAY5Txgp9kmmjPcVPrF3Y
rrl867OZApTZydeLcSSasJLvd0aiFPez5s/oXciQHcFZMUwtdTZ63Ujei2TtEfmq
nCqW9+2JGA9xKtBLS4KY/0PysfZbD24SRt+oR8MsXu3LLP5liDSZzJKBon7BMJuw
6EQfewiuFQRgYTug40cpqSGavayInQud/RYIbVOeR9jJVBHkmFDoKvEprPvLBqhD
38NJgHEA+9affGaV0U1ckdNscT7tBxRbZRJYd2gRGxDYN0pUSRD+Mqm0ksuUts/E
ArOk80FyJqZB0NrlQBQrjJu0AWlaU1bSK1pp3wGwtO/MUN0jyXj1oqCqJVeUsAqS
gcmppbrU3m7jHqANFjhQEWMns/yUHVDZTojw+iXMR4mUkWROU3ouAivtGBsaU3Rn
kONIwRq++Sl2MoYxQrvYW9yCs/oRNGfb12YZLqwcXCkQjQH7EOELFzNIwKMqAZQg
9cAvDDARyHHTckhMw8wMlCB7gNWB/mxX68unFv2IW2h+COQDLvYoCQPCRVPor5mw
T5G4y/V8MVPyQWnhGtYMJAQKpJtmT93db27I6HRwcjw4pH1VVoh8EmlDsip1Rtu7
Ftpx7HmBjntQcOJNpDps/fE+WhZ6wDKtpHCsJEN2NW/6uTpU8hZc7jCJHEO9C/cO
NjQFkMZD3Vfm3cYY5TI7CO418H4a4VCDD7hvBkfGjlzeXan101jRUFeX1HlT/Gga
o8uRfUnuE0gPYG0+2HqbqfngH88I2PAh9tKDtd6RUsxGrq5qGJ8NtIzKsEVVRA4d
hbfPmI/3aBNyOLjj3xhqgQ==
`protect END_PROTECTED
