`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDOG5IArm3/AhYa7bYRP1OD2cy14g0Nc0ND/FLqkeo+Jbhxh2A51EmJEAXR7+CG4
0OKHFZDHJuWPrmb8KtEcLPMiwwzaCt9tOn/gnsyIJoZo45CG47XAk/ynKMqP2Y7Z
8h7imKG3JPKg6PUz7m0f+W8YjpSziRbejTPRAILs+zyzg/N6es/kkKR8upUw/hrP
REsOSHw9DZAJ3Bt/olZqNWWMQSCSDDdww+SAxd6aIVObF/Lsl2jGRo+hB40nyQie
yUDgqPQBekyFeOhFIsQvIfKfIfckegRPIfcChM2UgKNbShMhp/Uvv68/i8i2+KZz
B3TLLDevX7wSQr/0Z5eKDcPlIfuZdMimO2Cz2ltDQbapx6mV0dMAg1iViAZ3i3G0
Y+hLMA7XUSVUEkzt6dtNO2YgpMYv0dUXgn8tfb63eAKAKd9nda4qT9ucJcNx51O9
+4QjuKOWf7ihNyZIygjtPco/5n6GFvmip4oE9gm8Bm+emSK0W4097y7t2owaCASW
Ui3egsimvrQKIGLNKLvHu3Cq/wNhihmdUgaYctmXXlScZ2vRrXf/tprsxgpS2pq6
hf+f/3bDsnNSUlFFt54cPBqusuWuDzEAr26mMt849EXZxApH7/bgFER6IpzIo0m5
vJN0BSmGIDxu+42UvQk61GnFoEjNOQJHy2PTYJGXfnxwY0z/SyYdmHEGETpURFnN
T3wNG55KI8o1VX2m+ZYc1beMn6J9QcRe2N8p6ZuUoavQf+qWKJKsX7rjepVIKAnX
0zkxEr3ToZWsF/22tUC+GmZ9zyFpcgN0mzYoxh46MPcKAYp53x03pPfbB2zOh0v4
jUr68PRRKNiQer8nB7UYBrwqwznIy3ya4NHeRmcrSb3aVNIKPi+8xV5o+1Wmbp2a
HxOfzSZU+jfANV/hWJfu/0B1l8RnLt4HKfS6yhaCg/DFQhVOJ5VPZDt33P952MCc
3EJyDTQRjX6bmNMuTBs4PUCFft+fXr1CubOtZMZevSivAi/Eyqol7ANEOw64PUj1
T/tOS+nbKiJwK+pnr6zOoPVN5MCwh0N7834JlC273yFCQmXeYcr+66H5kHhnz1si
SsUImUTdEOiam63Aque2wp1gsWAIyO43xK51OtIcJrhSMh/4+39qvuwTgxxTaNek
cl9ymxDFKLmQO7OhSVuaib9Ne+Lolxld2nP1dMiMk8rKSwjcRX7lszMoaNCeGCFN
9MpQ6vuUugcPhxEkA8wr5zDCfTs3aAECzPoXOaRmTHqbF5tfvndxeNvZS38iEZgn
zE2f38nj4Yx6jEbr86hp6e5KA8aMiD4X5r54F+bg/mUkR4pLlM1tRxO/XoFcKj+7
voaCGFsYu1dh6FRjqM1X3dGMd+5JN1f0aVkUj0EO0O3+L37jqzNq2np+bFdEjVX4
zq/1oxobksDvEi9yS+5dirj//4PdWW6U2rdX/ckCD7LyOo6wgHjzQzy25pNDRavk
cPNbu+W7JE/oKqyuufMGqm67UDZj/3GdnI4RHSZLm4b9qTRTg/Ai1mXLplV4Of15
t0xqfHxEGuv7t2ncGXqmDTYSn/aIdUDoO5c21uLaS2xtE+/wGyadHY0NJXqITAUx
jzvJYpWKJ4PxfTjUPo07ugIeoA0SmBi7gqoJBS/Jy5eILqm4C2zCDr6rM5ADmDUo
8hcpKZRWGZyHuSqqs9XWOHeS/B/sb0oiSa2p4wZ7m57wA1SO+GenRQ704W6VeEeX
EuVz8oKlJj3gMRQHD9vmEqxIRFuF3+r/1n8VCPR+XSIC1rQP5jLMiGbywizN5Efp
`protect END_PROTECTED
