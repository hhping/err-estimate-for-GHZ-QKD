`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beCdCMZeRFb9pfDyL8rfehCb1PJucEOwpUG+DbYhC/3RNEr71TTOA90M4CjpBjxu
P/bNZe2VxiuAZjnHmO4TbNRAuBRovr+Aik9eyknssSTClDN8Uls91t1+v5jb2af/
bu2LL2Oc17vqEfX2NbphlZ2od851rBM23Uz1dfB6qLHYuC66JNpi3devoUYvxQWr
mz8PikOhBUUnqZugDhepQ9vPdDiQQgvZS8ZDkwoJQ8X6PwBroSOOhPNi4n2xYQyZ
rCaQSoT/wLvWNHmXaQcnPT/p6aEXIfHJEIlbBKhnkT1BmzGqN5MPtPpUam25907I
tAasdqbtChCWnkqfEotYFKz9V3yn4kGs2Q0/oTcAekWHRTNI1Gv/cbycdQLs7Iud
b+UJGbTYxZvdTugRPk8pKcwzgWELX4+mcyoKUKWyDySe7GIUY8xQtUPB3ecySXZF
`protect END_PROTECTED
