`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
niZ9vwlfLhXx9j4ez7oNnjcA9D1SfdduLon65f7EBwpu+h6A3lWH0YZ4KMZ3XvNk
gXe/87lb6CSwwycjQtZw/Ttzm+vx+be45qB5WaDOgM6xdjV5uStFhTMfs3KndD2i
sbopGcps5QKRqfP/W17IbgXCfS/hF+ROVXl58P7hlfy95bXYTwF975KyxnNcqpxT
xBAsGEU2QMhZVfPjC+0/fFczM07A/VLZ63L6FWxI9ZkFne2uiO9vgCA3Y+4GQS7+
bbFDJg22QbEMzMQV6fmlErAXoaMMDc6+ODFMZoyjCwU0rz++dj/56NDkzyaFe5QJ
7R+S8XuynbYBZV1eOy5Db1IlpbrE1rLy8rgPjIkkBiBRn+/ZcnLGMMO0619tccuw
kbTCq3uCglPdfm/m9Od1L09XyerFzHRJY/MWvoku0sb6uWVKXgf8JB9BgMfis3tc
TBMI3W05I/uvASF8z1++0RhP0Orsp7/hmOuY0mhYLg5JVjSAyv3JvG7f/tmO/VYO
mxVkp06yDAgLoG+0bis60CWM964U47YYeoksiy8f6pJP1x7qIrfsMmo00/nPE6B4
FlV+z39t9jyEvLKOB5RCObkUCtCQXsekQW6zyPraLFOTPHR8NDukwzBMc3gxglEl
JyHoD3yqDP1+sXzlTjjvv6zghgpeVeOfVsGprxCyzsHhSOeetpkd8dPCNgU0bTvR
BzpPg73i+UnrFQyLrIZ2AFhi1kL3gRwBtOTOb04BWIFpnLkt8ylyXV68iiyaE8lD
NItA/HVIDOErai53+GulGowDUmxzj0d2uM937rhbOedq/3R0+0+LlK4xJ5o3hK7v
6KDaJZULKtTY5HVTVEbTCOEu9BvORXBnKbHzv8ANFiKETUnwM1lL4/UF25YR/7E6
hLVopeD2itTTPHu/NKKuScHNJrO7A7F5WQnofMtPDRznfncwdh57EJkvJmBDnfwa
VYnVxHcOQJFuYXuQmYwMen7S+NGi8HzE3memqctwKXfuOwkIkEnf1pnK0+yc9BE5
4Y2Vvefds8kpnUPXZ0Zxj3voyFwo89aGUSLh76mQBF+lSKARzZzAG9a2DUT/3kC+
TSFqqMCg0rQeB9AZSdTV4OYUxNC9X/Nuias4sZpi4rLc5j0Hb6mL2xHoTfxt4i1q
kcRWuZEErd4Kv63XmYYfL/rVHCmndE3bdckgHRSRyFycVilm6IVq8ZI3caF+r8xe
pZAselsCe2MB1GFFg887n/4tlUFgIShomx+AF8rYnRp9cBnU3i1oKd/TUOfVRg0Z
J6uav9aTb945vO2YNfSQE6IJ21s9O1C8wuJ9if+Du+CsI7D9nX1WLEUjuLz0dfOQ
rTf1uZHSE9yYD0Mq1BR+ScIV0512Km0C1TmfqOpULotY1uP5e3xvyDqiPOmW9BWU
DUwXl/Q2RwHyHE4dknTNoyDVC6UaqzWub0AiGsuuZ6AwVb/UTv7fRMOdC9cnSEnz
p2ztERjW1OVyVY0n3BBjaDcNnQ7JJ0iMc02nxKoaSDYilUM6gxOhVarEtkhXBvL+
7hkGt6Nl5FY1Lxw+0x+6bxNv8b/o/r8/MDjwDTjA4ji4GNheKMRy1RLeFFRDhI+h
zim71snmkvcsJ7vL1QdkIAfGSx3f3O4JQD22aLG9MvRkOgIQrmmI7askevtu2Z97
hluIYhBPUGQ4YgnAckQjDYzk+hz9bJAIfnOa2iBgs0XF+TJwV2qdZNIkhR6W2M3R
UDtTv+T8PSeLGUGUZAI1owune5x4Ej8/4xB9fcHDUepY76GWdcIbDHnhun0qMo0m
6k/rNu/ZhxikeUOGJwRq5URBcNPU6Dk+pyuKahMv4Kiv0EwogxsRbgrE9aSPe1V/
Ms9woiH25PxFTj/FnkuLTrZhSjruWNbRbNULBAnCuinButsrQb+cxQFB2gTHHIEt
TJgp5kq6X5YT2uwxpw5Vi2af2432crPW1ZHlV6ydJrc2oMLwe7ucpEkHcS6tv8Um
/E6066fHxKEagE9J3j7DnZKTCxbvFr/v0L3k+CprRJ1/XspZWBd4PTfMGfzXkpJk
hA7sa5NHP3wp0FlEh4yUaKmwPSbGfXATYCdPxEZDLQMWz9CC44aN1hoeIJHRqMbc
`protect END_PROTECTED
