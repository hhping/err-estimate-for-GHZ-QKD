`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
co2tmt5axEc88L3c+zrwpgqnYnNoIy4DzVO+YbF9fxTKylTyOQZfgG3ghC6nb8kU
7tYvucqrsRCIXh0ocGed2kFHD4ZlLF/kI5UvFho7nahTBtwxABFjWxSbfLdeKBjl
GXHcG72S1Np8wURTcoz0SGVldD4EYHYr46sYLbJWS7+JmmGEHNQXWduiap2YWE5E
imM4SGDiDsXxfyR5jVMefMiVpp6x4K4SIn/7dIYIAK1xnYAWqsd1md1t5BYj5yLw
+tHXRbyv7r5TmP8TxrC7Z37zbPBezJ9nnI2J9D5Sz/v0Pqzne+upQM6LqX/gbrkC
lghcIWn0hE70BiIjJ9sPJd2atfFmxH5IFHS2Evd+Y6G4m6YSySgxNZqzi5hOAUWq
Xb42DDSH2f1l97MMl6pM7Jv/I51IhqMjjvZWWZ3FeBIbzNalJipSMoet6kGqAoqr
z0YAw7MGDf4StVFAqHhAzkCqHxvpu9ACZ/qMApTYtLBfueV/Fl0L3LO6Ceamdch1
aX7mI4tdqRd20E3y+38t/ch5a6kL7Pfob7j20RrVcYX645g7QfS37N2DpvZ8K7et
n/miSiugbteJ+2gyDLSrPyliJHRv63aVEYxfRitevMFfH+hmSLEsW5NLHdDc0Sch
H69o0KGY+vKYktgSYPcJInnWRFCBflCQcR1yYt3U52QrQK/9DEbkHnrbXki4A5Rx
vfes81ih3ql0XKsiXEFSKWcRHaUMjM5EFDZhEf+n+42pjgl5G/m9BDNuBx3qi404
9zNPKtg2zzWe60LCFVT//fjN9dxxgJCFTxBOORDgjq+9tCOJ+3WsFVz1HXVM5m3E
Nh02J1ovHRrnLTIK6e+Mg9W8skEdHWCdTk2z1zqwVJgao1Kqkb3hMn/hw1nw1iw7
9/ipWXb72fGjWP+oJ1YheCPJVsIPFCqT6xGlg4wsnPfuBkAL84bo5nf2hsQ1nGYq
EryzAGfrpKoqDE4plIeiSWc3lqzqjIekLUJ8JuQkt5MulGLCCawbKOrinS1fUECe
j8kqdRfyxlRA28yUG1cVcjCpG3PIkIyguY+sCka1ScHyxuJikd36Xw38DR+cx5LH
rG5sgffftX+bA9N2ogiG2edGCPUqbN/Jwj9rHyUaQH2UCPekj44RGkye4CcUaQVd
sGonckETfOlnXHY8nsi2V8Pq/ARBnu+D2U4Tszwwy+u5rIxzeF71wPwB8j9D7no1
R+VKdrGW/w056i1nHVmnr3n6gdZ3A9o3Lw7DSIzT0czJRCBPYFifnjaSlcF3lnap
QoKS2fcMSuPM3y4anpfukI92KyEuKFCvlcd8Tqnud5uvk5tqmd3vHh2QlifmLSOk
`protect END_PROTECTED
