`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3K2HilaYSyDha6K1CNnSFULJATW8PZOK6wTz0WnAJKMsGMMguB6G+qsrCRhl1f4C
KcgvqtbZD9DOfJZQAxNF4qeUKtrMahN6ASdw+29sTFpwBjyrJ96NXjmgFRwTDxbb
F+Wo0gmdwd8DiD2N9Oh1mSBTnoW8rRZ6RNBhEGBwSpvEhfWrqh+peb0KA0FUJC6J
9fN9cj8uiN0qSLk8JmDQVdH3ATEmEARIf+BA/oFXYkyrmMl1nl0mOTTFDDfYVaw7
e1Ak9ofKA/9VPdZDtDh7lRVvulZxWn0mj8rj7OoioJkC5vOmRSPGVjvQFLHHN/zF
5mGQpYGV/BYrPKLPMGc81CW0H73OhbUDkSbU02xn+n5dX1Mg0y/EtV/sWvt4iZ3G
f/ryW2UID4JdWbgL1dZBDUiMf5834LVQlREljM3BPb9Rh1OdXxPpBj2GLBZ3/xX7
vutWBphbZ5rASjXT9rs7/b06FJcxJnS4x6tVVc10EBZIMnLQ8aGJYBLH/nF7Mxs8
CdJieTnKFLTLYoUi9GgNRR98vUmV94as0hA403LbjvflfbdHMdzdAnXHJm1yScGn
hds9Wc6s6Te8GdCR3WkoqHzHiJ7bBbVMNUt53CuWv6Cb5UPiwTqR6rz8mRBiYk0p
ToToU5pLwQ2bSQmlsH+uXtX+RtP81SWw2MERfs0freNhA5huDWpetvPGoBPLTwAS
Djc9f7DEZul7dSTpK6tqBAY0sOGFOBis3Z71GlbgyXCJ0X/hz2CD5L7q03NlG4c+
mFrE0pyzSROfeFIyMBNlYvjM/S7DnwQRtP/jEIqyQBJhdF7l0JPEdC7p95azzQMi
2SXosy1kDLnG8XL3DV5N/FKfekcLnOFc4Fqvv2OkoQUrUvyh/cglzD6BfHhsiRpE
+ppTATCusvBHm0MxQgMbJSYp9kOb7dTESC2ykMok73IQce/UStAOcHpxKudsw3by
8ez7T+XGQkMyhldMNc6hBr1cBcMG03CaGRKSH2ssuWkdtwKLz+UpjfXbLVogsFXQ
1KQX4SsoQxGNKFkP6M3+PCToo60CcnwNYzU+8iJOQuaC3zan2PkLg+vIbrAz6KRV
zDwNjyX+dGQVSvH6heb8Tc1S2XcRh4olwWGrcUtQ72A+KdD2AgRt5c3HP+TMhDCY
wKDYsBKnnqothTlMmI5gcPMAKtdXqel1GdH7+QNjA0smGifBcq3NvGedBCsTYyuP
g5vYGUJiMuemnDWfte+djli6KgYziJ4mqUlAPK1buh4a1NNHgfi7k47oWqS4e8Qg
MJToqxCJgjwVfafWutbgAfnf5n2Xvp2o7xfE5tlh1GUdNeyNOhFDXpF0nRR+pTHJ
bSqYm1ofsDUJl0oto8rtjqHrrI6pzqiKve71GRbFSpXZQxV3Hjo2EoIFdgv7g2O/
i6VwVrckCuaoAZdUozF6Ov2g69Bczg3ElH0PnCLx7tYfp+DkUThgpPX/a+BHD6Za
JO+ZjfJWZVPIlsjAkek7VBBt40gmlhC+geIsNEqeSU3ov6oobZz1WHP1R3mqCFh1
tUHcSKKWvfzeDLq5lVUNjeRNbtOXrwwdRIUhuNb+236Uxa6edbIHMazE8cRrxYQW
uaF1kj/6HjQ/M2NsQRaUASTOZnpGnkGXNqFgCrRplpM4aYPkpMCWf4HNvag8hYYb
xlh+ruvPAgSUE1fE6h6XSQ0K8l4IBpnQSFM4isQlzNzDMA8Xq7m9TRCvwP7E3f1S
po6/Cc3EQ/mGZKqmVouLO1X3HhIxg6cdwqflJjTCaJ24nFiB1SFah4FlgtLPRxD4
XbN/XTDvbCitg7RFMykikRYAfeRBlholWvB4gwFdsxapJfY0g33BIuFhnTuOAtVu
B46eJFm9iiS4v/qwHxROXptEQ7fSM2jHf9UagvpcNDWFZNsKzisGDccgKvJykUko
/O80BdKNm1NaT7vJH3HEFLRgxGIDxvGHiqjIcGPCqoTqpJ2zV1kd8l1huYtBpFyC
frHNyc5KZw6Je7+U91oytFYIuN+gXvVho/VS63QbVZ45coG7UYUoRBG1t3+WDBqm
yMuLiXgchxkasFN7vDbroAG1TjIAVEZQ4DGKpwziYX4b9eHpGBT2xIsgD9EZ4HBu
CMYtmk4lCfllD6f49/ocid2dJFWLvVE3/qM4G4JIAa6o1SBRWW4dE9PvUTahdm/X
8FynM6HwneZQGgOnmbg5e8vJQxF3ONGPamQ9sjKccEVzn0eUAMAt4ZhHIOj0TWV0
OL/rM2YMZGrHNzUfUGBgCgicLaoI01biSCt+ChyJdiso26erQJtvTYuPoJM9lmmd
oRZAntO88v5CECj+YUnHLNfH+2AabdwUAQ6E7AgjZWoksBZeJp1HQx/fqKWDsUaG
9K/MFrbSED/oSSEFgJYheoxzPc5uW1eZ0q1wzqXmTVRT+YQ1sCsla4Ir2PMl88jD
MuIZxaNHhtuJmAf5DnZnaC5LOj18H5C9hKpii2Lb8jP+Y1sR2BM7XliDNSNzDg2c
5muRIv/WBGs/0VFa6UZ2f1CJGHdT0xadHgRheymPKQWRNcTb4tgixJwl4xwTIHqZ
vSOeQ0U5YBPyuylsU5tw+jSk5OYCXsaRbylNAVptAfGLHLJDJPkkMbhAONsG3hz2
jYrBxeqYKBJEvnxtAL3O3yyPajw/435wITzIsILt06yoEeO0XgOzhhcBrS5Nt00N
otU8rotADB63VTsCkviVG8baONd0bpqllYv4TIRRJX0+dkIeDWQdgQauJLc383h1
wftWRN6MIqbXRj9/9pIPnjvNaKImnwQWVQgmMGxWFK1nq0A/juhRwp1dEOMgJ5eH
whUJZpBKniwUXrjSbmOw3z73H/DQA3R657bAVL+ENMgMgGGMh7iPVkqh/AaOlRGE
I0rktxsx/kHKGEKHGgZ/+z1A6OsxPSrXDd8MtkR4KzAlVrGikX25WcoEStSXUV9w
`protect END_PROTECTED
