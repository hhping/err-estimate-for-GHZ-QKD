`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UF/3aAL4qxiaSn+tKqcF2lwHAkEDhnvMcoHAP96a6DC0bECpZ5jd1LMgdwqs3xtG
WQxMlFPARTCQ4qOakJaJitzCCRT1X3jUkGGQoXF5IhaT6y90ugJUa2sspn+3s3HP
Z2xBYFHgSrkJiDwrlEp/hURfKNYXx2zV5Ylx8WWmO4XBeN9pFeQI8yrz4M3uIYbZ
tsjzrjgNT8AIcRUnYZ4fEqbCGCxD4u0qcaOZhyhKzWTlmd1kGCM3NluU9sNamTZQ
9PlohcNWIo0w4WtPnWYlZ5v7OZMA4iaoD6gLFUsEB31lWTH9PkK8HdF7dkUUbOHG
CemOv4rDEV8b4v8uTScFhPoaj4rbrOsSWTYx1kw3/qRe9Zr95WvRMXXk27pFLDPP
bjS83w0GlIQJ8k8zaT+zP60YUlY5rZDBESOYlg4WKcykOjDKnmg087Z3zNuObAFK
/BJ2Wef16j9id71XKtnrod2HmqiHRfatPCRSCzbtu56VgygJgfk9ORVOVofnUnkd
KXshSCLIl+RbjePwZjNMQbxwrY5rFbqQ77Kafo3ifVbMcQP254Tw3EaDMaQckHsT
uqn0RD1Gz8LGziP73EcrgY3wphWpXv6qLi9YiLLevsMtrElFisc8nNmlv25n3wby
`protect END_PROTECTED
