`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3i/XoqiEePOpTIzfSG2WiCRyWYndfJtq4/0a/72TYDlBjAbWAt2OMesrac47t02w
GxuBWVGqaj4PZIihnU8rTo2JIf/g+FDQuKTUs/ZbYvalxx2m19K+7ELwBTSx1QM7
x3dDhevYeQjVz0G9pVJl/1fXz6VLnotGfoqMtfosLnWnknYUEf9680vOQHfzLuLF
bbmBZf4QrzRnVx8IPLnLasED18XjjyuEDJEQUnMf6//rit79yYxYYlEOqEpqbgxb
6ovNYDwmHhZAVBCuZE/ow9CRUoZ5dUkUQqoLedD7Q7+R0xcBRp8H3GHidDkENhAe
aAU62L/cr1obBLLpA1YamOaVfEGdHINo523T7boahLd0QlKe9dk2lUPIShxot6J2
gGukZEaFLu47eJYeAzb5D13Dh3p7Ltr4A5AWssJO7lcgrYRcMBynKZgoc30+bpKR
OEA+LHejjzLPu+GS8bmynchafxhDqf/czwn/3SLux22rc+3s62U24m2C8cY4EjeP
y8vX8VraDkAgjitSWGoxKoWr9zllXmMAOrJnspu1Yr5jt1WWzgokCWAhQag55JcZ
FweAJYdbYPATI9LQwwgIChudLl9QKhGWRhLCF/4bT9AIZ7l/DavBR1fkIz1a69Ni
k2Xdn8ciNg1Ffy2D1dc/ppF7PHou4gOyN4W/8dysyHa5A3bbjiZ44NsFa+X5qh1c
342/BtEiZC3DXfPtV4SvyQLVkvV7gy4w/8o9bujt++xHonHX/Lo/YZLpk8ZgCZQz
MH3Y6OnMvA71GzblLpBfpQbxZkcKs7r7hZcIl+EpqwjFENjNzLNoz2H+HekWuurR
QCLIpj+QMzr2wiAtRos3ZEh5p/937FZEZyNQNvya32Z65nIsbwbh+RLl5M/HHVWR
SRvFQETN7HmveUB08zSuwgvr1TGuUZqmPMPDqrH1+zfZzZFqATx44iSqWI+QJCaf
Kp5eAwPbhfnC8h9JQAWnp9Vv9zVhXvpLj7nTjJ4dkTonYRURUBL94XhMzl8kII70
Ompxpk2cms7muyEqcQPKXDKDsaVHfYnFsc/dFWaMYSMrXvflefICweqzdVIBx8Dj
07/yS2XPqLjKBjQ0wXCJDULATnHp+RJoryB9PQm23b+MNA1Y6nEH9XzcfMsRhdZF
nTVWn2iHIK8+z0QSsAS5vvwVvWCVVYg8OTnEiXyjSsaQc17Ar60xtKRHXHsxm9IS
7pEJecLlusZuf7MZZG+bHsynwMT4Uqm0PWijsqKEYOXozukT08QeejwHVS2Rk9Cv
hPP/YTBcKH3+ZQT0qcQRuRJ2xhw+qYgALPQmDx7niAn4+YDlvMJzpDIuwzy8zcoE
ATbKJul/FaBB2PefivrfH2B+jiUgJXJLaBwEYxcIynngk0ySkWyqE0QJPCOt/6pH
4QBU0v79r0Eq2inYjUM8hEnPvXFUYxouQ3Rpq7pvwPygxqSvsBS1B5FUHFIvs3j0
JKBB6vlrPT6uDC8/V1F5sIDNEqiqYzK/fsZeFlf+C3W1Xco38Fx4oP9B1E636sPr
lLUcxshlYsJoFGpJ0hrrxU8DGgOLb2RuLS/mJwq6ZruzoZUC7ddMlVhHSU0UtCKq
aX6fnIR9C/k40QTHaCiwNwI7Lfx7rOYqs8NilAc319tGnJZhTrcmbSLHlzhLgrle
/yfBHZ5mBX3ONKtU5IG6dCwhc33zi29Z2CN0dcoiDEKsWXhRK3+24VDWi+RbPphW
6mzx+yGn/3bmYmDLS8BAf/JkoAtDpDddO9L/CRkk+dlBZtp1mXeZ6R/R68YJ/u1w
k6xinuXLiwZjlB7tEMg+NHpj14+AiUQJf1PGiKvx865Xq5PME+/1zx5KvzWT0OQG
SN+tt+7CE4oRnXe6w6KtZ0eDRIZQFu3l0GqKXuRSPSF0kwROdGxeHIL/58O4uQDs
m4SFZQuxlsSXvkh0gAoxsQ39KQXdVpgqCckl4TQM2JpmGvPNe6aAu5z50+Fg2A1y
R6ruxAenEFhwiYs/FY01MklCbuP1NIBYDuYU+9xbqAyAwyZ+36HUskUWAcdzl+vu
S5c464uFVZ8AVw/2JXriPNjOJPfq056sgMQ+U38N2/6kdMi/0UKFdb7/nO/Pcyhw
`protect END_PROTECTED
