`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wsx5+baWlmKiVyd3EIKxAeQmmqyGQo77ohetv/vIMiRkDaRqhTzWcMHOdg8NFjfR
qhC79E6yu8fqGqiNqe8O5ze30rYRgMXYLrCrXZ1Wda+P1QqH4bKCuMJQiYSSLFNS
6RR7yt4pCxKOKuqXUr4d9SbyLLAt58YJQXSpR0qBt0pL7zs6Ud8cARWqmbUZ/GTe
W1LbpL/7SJ5ZiJunM2grZ0p/cBcAvhR7GGi/3KfhBhfDxUy8wsA59knwhQeIb3f3
ezakIoAMkvOv05rZnkYEqMOk1nbv/wk6nF+UyhJM+ShXT3Ty2IeKIMhxXmytpWrj
2OVwOqTj5A3xszS2E8g3h4nYsv8jewYxNczYLesSOSXLpWQ9o7HHonGR2I7g7XRo
XCo5zLn9a06gKkUIsEUyDjwha8lF2lGWm6D8LtQtVD2DUXSwM0EogFShr+FiaEag
cvP3Fmfvk0aY5uPhTV+IGv5vkhMy9oCUTKXy7kR4/6a/jhhW9unrnEhTVvpl5q9i
JRngemUJyDL2h/cqIMyK7Ud+fvCTzLCzmDebm8lrypeJ1toTNbAixTBBTc9px2L6
aZVeFcpEymdtOFM5Vx4IxLZ0weayN5/gmR4bTpGSBcQYkEaS2HzBAAz9vMBF5a5d
xHunkYILJHp5pBfyEpdkgQPmQawVrxhKmXGgq7kFCdvHg99RuoVS8/luwWEKcrRr
vy/9Ok8tA408Q7cvBjSFKoCoJRkd17x0IU2qYdFSS4hgav14uKq7pMzPr0186ARS
Na8JSuyyw/bJnraW2rYBr7wVADmYaxt65bYbTY7OockQok8xPU/I0zp2X4rfXHSD
QOQyvhQGRJ0OamSJjHVyk6hT5B3UtdEGXCf3bZonsAcQzJV9950tBFcKIi9ZSU++
9DhPeOSgSlMZQnRRUEsWsl1ixiJA2KPJdUI5TmL0dMIkm2cfVYlcWxzCyomoCntO
YzikZjr/aGCaqVSi9aZoNt929MoMbnXBEkbZxx+4sfBsyhOoMFxEriGtGAQc0YvP
6OxG76TqflQFcp+vfqAxHLS11pL28OpnIAKBzafSH9fQcZBrCYHM8Gl2pzd+AiYy
ErZOcXYmo/k/rG2BW0d9I1H73ixoZf54rjFcfvZ4HAf9ZX247vZFkjHVSfBr2uVF
wkl8AXSmAW53hYEU8BeG4vL45TNmOd2W/aENZfjusJKa109RkHOHkKd2vdZtWlL2
rFqDJ8QWq8cwfF/iF71eU5CVnitCB5noi2tqUL2qXBCvpjO5gzxXT6o6vMi78hH/
F/o2neBuUDnZGHQKgrYIVW319M6AMJhz0IyZ5Yas7l0CEJmSvrs7LZBQJ7wSZwnh
JS60i2qbf152ZBAuY283UQgPxd2WuoiYDOdSXs5e6+ueT28lJIbmjbI1VtiWh5Ts
b8uS6RsfP6kuLwtPk437hVkRy5DRPpSyQBRvzzqFUeQigJSp76jMgc86kL/G6ozj
hCPY8hNUFA2AFLePwYfCF6Ss8bZgJw9+VvZwTET2geUYHkW6wL7RXpAsLSm24XOf
MrzW+nHm0XQRIiFAuEIRt0hw89gz3jf7KYOsSeqAzK42QlkZ17DeDalYkp+JjeCK
7doaZl+A3ibFp7IqKN4JAxf6DgtkSNVZBGj75p9c4Y1sG1S5KLfXtUelGfSxecmC
1H/rJEaAXn5yaDmmCx2ZJFsQgCSvLniU7OqwVU+lR8e/nLPtaygSoKJoAH/RLGtt
sLBMruaeQJoca6zvEwZOwH5LqucGEulxoAVUHzKmTcM5+3D/CMPC4Pt4e7Y6f4ne
aeB4XcEY6vK4Qr2TnbGvDhxF/xivoKl1VZhFYRq+ULYq3eqm5kJVRyGloqQKm0Ez
DVpA1P59QWjasWGDRysITMIa9TCbq4o7+bB3fhWcEajxxhk6noanLOEiRtByPY0W
pnVq8rSPnNjJzxL09MjOOmD0B9EbopGIsWVQ8XKl7URHtF3UtsTnxBxsG0uhkN3E
/XERd/gjuzbW06GMGDyo849GZ18ttq4Dl5Z6p3VT9YXoKLdj1VtdbD5747UDNOwa
ZuiZR0QPScd+SgHmpxcyHSGnfJvwNjiQva2g98cBdGI8pqVWuf+q21HvWwyIA/0j
OTZSzCfe9MFMfBBNkiJXQ8MUp9uOnsEHjqDzGN8s+8P7qk4ISeAPyitIX+ce97s7
KnMUaqB7IOy+SmaVPk/GMsDVcQ4amse7tpLwDwOVAJzh/CgbpNn100ex7hZOuH/4
wYKO08GzC8QGTBGiCToIUjaiFTDTdNZ2UQwFYGyHQtWqpQiNJdm0qfUaeEkTXjIS
9LVfYnZrMBC0v/QnU6NuMSmsU9rWi7eBzLqmFBE66ZkxD8tgqHwFZLZ5EFefnhy6
AjEKfhzFz2vfGGGhW3HhPttQ5xzJxmpJfS+FJqancQ8nmZnTrrjsN8S4X57l8beX
/ZRiuf0lsH4gigz3QF9ilacbCVqUlrWE6nOsk+FC9iVtac62bsUWtD/DOCojuSwF
wre3KBlwKL5o7MElq8GuioWGlLeMA8T+8i3b8lkXGCm2ihFn2pMWZO9Rlqaa0rrb
mAueI00NF/C1tjYhSP2sQb2T4qeJG55mykvhqE3UrkSYVKDzDK5vjk2BiqwedAfk
c1DtdCTi43FsIL02rbCu8UJkOB7UpPBuhOWygxIx25EeX5tFtFzjyCAhNhroMsm+
vYSXPm0wtJt8qYGZhqW80Pemjk2dSti+gwyTADNv3jklSmKWGoIPC0JH1vqnQBL+
TiCbcSnrb2IW/x2efF7sG4Drng7ALJvkDVIgcIm8Z1MCx7ZydRVDVU8iM68WnH/X
ibdqC0UvltT2sr0aipLc9lFAxauKwLId7eWZQtmDcngmysamZNTO/cXlr20E4Qcg
jhcUBHRp6rjhHsbo+i+6HXy8dmsl82NYBWDXUsVeGAIlKLg+VeD5IbxJf6taAyQ5
7aTmE+YcLddulBHGSTcLher6UgMwYlpom6lvbHv9JPCUuSSyl4I6B2j9/GsGcaLh
POU0KL2zmXRj6LKOOZg9noLgNHDS+STeH0LiH0DuRfZb5vAlZtlGssBHTbpuN1z0
NOPbLLM2+A50w9Gz5a6gjj2y3sPvidkEOaa+3iYxp72M/HFsIB5TGMDPCw0lWWtI
48F4fm+/jKzRv9Ce75p7XbZpchhxPlBiwE028bZjljD8pYAk7I+l+uUFzEJ6SPRa
Nc1l3NN5I+vOIQ1KIxqgK7Hh72KUGww7XhtmkcLDj1HR/tlMSYafBEuAw2uiuUp7
rC/ef8V6VE059rMfmdbpQ2pRASt1fN0IcV2GEehNiG6F4BvhlicZKNfwc9OOtB9m
Vi5UK4uoHqPESzujmR6lV3WjMQmUJRNO0RaBvpUu+Wa6KMX//G5UQiz16UuGCmtB
fYnGLD3Vnhr2V2r3d/CZnp+zyt+X6OHkVoevL0/Cr8kAFXX2yYorvyv9oSw8+/Iw
vNfrfAfF6bVOXxPKALs3aSk7ntXwyb40R9Pj+SP/AdnyQM0t3s00nneAkhfVlqIj
nLnDQzlV/hqiyY8RyCS0zoezKGPdDWHB7epqdT9pGWGAoQKUEMszA9TCAhJFY17H
PyE1nR/ziUKXELFnev8ukHtHu2MTisz+YMDR5ht6HQZGNFfzJ0qxeNxcSnHgjyk+
00OS1GaRuCRpU0PybdLxnqLkfzdfaaZF1wTnhrBRywY2T/GmabgtSecED6FX+JkV
Bp9YHERiU+B55xzXjxoG4R616B+ijGE9J+8V/4GYl7P7bu0FbuHNBeNLJ12NUPkR
6oj+hZQTa/Tjeicos3vCjShZeVH5RS8Crz/aDcWvxZsTHO3nkyKhKLx839MRhRMa
nvmAqEmTRQ4tS7GTEFHKctM5GMbC/2yhDDJbAHXwgHnPRQM4o19ltOBHYQk86+5v
I5k/8GsSzLa886nDOR7owMSpkcOIK7rcbZmteCP8GhSZ4oPOO8HB7CQ9trqLRY0Y
E4xqTcMT/NWHTdZN3JRL//jUKUu2PI/o06SfkM1kaHshUHqk7k6b9TldORvCK8VY
hRjTV+GvsWZpqYc1CmZXSV04OGD3H4ssNQc9q8+BW4GsaHcLNkyplTCCH7m0lKk5
3vcrbBD3/TqiJno2FJiROOhG4VI2TUBZZGli3IaEpNxqx1Q+qbje5mYvTpz5ieWQ
P5BhhcwK/YxGT5k5WdynnANwjN5dUJc3hMLJnz7/86ONyfnwNYvkaT5e1dbUuI47
vu6wXcphFbtD61TX5EWmR91ygu2lUp+NTc4iFthwxkB1rjrgrs/I9p0F75g8Vebk
RpqBXKebbGAwN+XXZQ1G7wwtIMvzZWHkr1ZAvoVFceUZVjrEEgD571zsMw6TlMer
ibwW2WTiVYYV73CHkQ0zdT6Z6gAQ5Woiw1insodl50T4audiUOI4rXZMFz0tTdzJ
Fe4nNfCW2oeFtEud+I9+8I33QSbwQUwT/Ikmbzpeq/oOY/1OYdxMTyNi25Q3a1Rq
PRqEo/opCjLf73PExq16acqOzhdi+IMGNHH82bSr3xyutD45YRBTRH5I8dFaWoG3
dDH73W6ZbBJfZFENADwRTIHwDht4KFMlCka6HMawDwGwWXXe77CYbPW5guSxud0L
cGBaALgaV0N4emnl/4HD+jxc1i0L7yNvJ3fPDZhJwQgtXu/fMyXSsyfyJPaeFyZC
Eg/zhSn2I6KHZunWbmltelRp7O8JvgpBiB1Rx/7jrHmS/PEqyY/Dce+bABccqr9N
uUeKwJoNqgI8EAAm0m87GljqvvxZZdA2CtHNgOUMqMvzpr/4XROYvrLbSrp8gUM3
uZqHKFaPCOE8aM/t9/Sml4MJNTXEd3Yb2GqAUqn07lPuV6MKyaWLg2X9eHFN/y8K
9kcxSPkRPwFyhwpuiuXH+Uvfb4EvckPhEuFAAD2A9VpKp/7DZttPILurEmcoH5Bh
EWBNiFDOU7+in/s/h8QMupKZuCYhFPPLsZ40bcMWUxSuuqL5JP0HuJ4ZSaANXhli
xZ1tSsc+4/sBj1h00ado/sanqaScS7E1qxxKx4BS7R5IWfIHcG/3EziwCBfOBsOk
/cihVFnmeP4rlcXy1z+zxKxLS9SpfeMb6caxwvL6LWVtTvD8ojwiuL3wopKhyB2G
PWgPsGURCfAvyD/utRI1MugAULfMrc1bU5XdQz+NDkAsA5ITOPorSP4YNO4wrvSx
Ppfju2tQvOLbbSL5cQHuDw2NNgUVX9GRGhGQHPR69zhf2UUlOJ8fXmY74Y4cul7R
6GU/Gmz33mSLnZ+Gq/Of1W1nRRclcI1CbAwsA3ZItXO0ODhoDoqoSxLltxxa0Umx
XAIxQdJwNCdquM4Y3r0h7aOTXokbwmGirouLFcjYK7uRgIDW4wXFHMt6reVzMLP/
SLIFz83US/VLodCBQLjDbWerTwu7j4dVBAjoXloMTd2VE2OIO9ptam9+de8UR8vl
3fT6QrmrNBmeF5HYLQKD8oq6EcXh4YuQsSBLV3IfIFro/gURo01AnoiAiTweYmO6
/4yBqZ7Zp3VuNTxjXLy/hcRkSqaF9IC8efCteipn+jZ3GqCsEkYVZGz8BPxW6qFk
gNWcPgYPWXgU2m85hQ3aFia0oXUxp6WIXwyUMc6LGC2+CVVmVkmR28CId8amxbBM
ltHqDEpqZfMksCFW7fcIZdT/MXlxvP85j6jKlHkGVMBj2QZA1K7SwxP96+b7vlEA
Zckry0wOSNHEgc1OTuhZE/Mzw0xZvs2V9z+mHjhTMQf+/arAgAlVZHVodd82lA8N
DAH2WPH4KmRLkRMI42pFUuEP5pH9cOdGeQr7fKYXADCn0ZJ6kl2xwErKZgY8IB4a
qaT5XojczuV1bynX+cP1qtVSYGe/oyKpTDXpWvrtUS0vG8QpL8T145cJvJidaO2u
OtoV6a1ZWuVtfNhLV4s6Rf9QYxviz34LgdE7LciDXaNVOBhYAhL+m9EiPDjpyeWX
/MAllC+06INWNXs7/DTBbsdbPpDuQBLtnIE8Si9QfsGydfbK7zIvZ2dNh24RokJs
bHy9TyHDu4o8DhomkRKatviHW4jAhCnsMyceZyPccwFaNbxpd0GLaxqiVLTHKOok
5q23/YFnR/+yiCafHAtr4XOP/Uo3ljpvbS5XzYcd5c/P0ZZsUvCdu8KyAs1MOZcd
6UUDa5B08Z6pq5ueLWE58MnftH8vyXiowDmrXL0RWwDMSVny7RECSt1wl0f+CfF1
R+yPxAMezK2Rpl1Uhc3Lx2GtLFAgaM+wiuY8UBOVz7pzqkNFuaXTyzGG7grEwMtk
oo6rf/VIXFbV1WE7ZkElCF87CWMRTOz3+mxsxiEzdlFz61ooxAB7Qda6Pv8++U8C
jZFVMn0p1p3mo/BABC8m5BleWrfWSLvC69dHnds1ZFBoL32Y4ol8p8oOUP+sLJUb
SlBJdKJLymjczST/VaS80e9fKOC/GhHlWwfmdzfFQ7GqOa8rei1yvq2rod5nyBjw
l+YTOR+yMSj8KjDKJph97f1FQEoxmdGtBSmL7yS2vFVqyzr/rDS0SD9P3yJ7hXad
VRU0XPzXk7fmKcvMjk4/vZs4sFIGmv4MOexr824Pzv3OLrx65vSRCejQZAo55o1t
hS6hcqN6gBzvrz2JDjf/TFuzQ6tMzwqyTm4VyxypuxsQvw1NCh4atkqA6C5eP6dE
BDmkefH0uRxQm2Bk8O29FuJNWbSBtY4kC4uYn5/M4n+q91UhfkPSNNA9uwW3NeRk
Sh9gRLu5dxcVVV2AgRMXPnrz3h9Ah8vwSlRy4Esb/DS1VIA79TPz80Xa4c96h+1z
opYLJ4e2rft9bOOW01Ck9TdmMJloLq0VR9N/L1TqdCPRtUK3FLGPgbsqIaIQG32Q
+4+hd4m7P2khwC6/Nt7cs4hVjM62ej630z8HdsUsFB+yqCPa3uBXWqDq+dBFdiD6
OIYOigOuFae1shdglf/qUt6zApqXTRMdoOeZsDJU9kIo6jj2wImlQNPjQjkkQ1tR
bm6274BX4tbOL/fQYcmd72q+3jGgglA2YsXPHYEecevJhlb6ZIqixano4PCcalps
aBfq1z9cGtY0Jm531S+ypEmDhawsxRR70hYHNP26XOG3aCB1rtTz+DILpdVe9y+1
/xwdY4wteV6TeTzUMB6GEgC752TYE8xO+T28eLWeqStp0IZZNhugvgRYZd4PN9Gw
2gkBzuSAU9qh6X5uyQ5SUDO5FYv8inv7s96L28bDDTMs4StofbvDHZPs/31K/62h
rm5ALbnT+noS3gab8ZmzgASO8X8JLnJHnNz5IafZRKtv3CMUULvtXEypw/CcH78m
/ewcdGTE/eR5ATcjPlSP7EUVGFHw2ZGi/kofQkvuKREHKOqn5OPJ3h5J3f1UE7No
o8dTmj1fPjhxXns1l6f6ggX7cLfddjl9qoSSfluHGWUcjbIvtaSw4wUmXyyveAW9
pRANhVd9MD90N150T59OmDxVUOu63zeUIbk9tiy6A2Jpn7UOkabKEOmPXO46u0Et
uit6brvBpA9YVOaoCF4HZNgU6gLAJEMYyTIk/NjO8MqY3tXCNc7LrqT2U2WEAwJZ
VfQnW9cjuLRazb2kXPiJubB7ssI/WYIvPgZvtDWIsFU29P+9bJ4Y44eBZx+Q/MXL
l4JHtUstndUzx+0RZhZo1Oed+fwJEftrwrqSoGffqY9/z5UFhaXqYl+h61qJWVzU
5f/Nw3ix1HruRPIPG37w/BtijINKC7rOxkjoCOATXFiV7dWdp8cJvXdFBQyjvcBC
B1OYt9LRes+d1nfV/aUyr8FSg3dKnfhqbh3bfA2T4DUOv8plfZFSc7sx65SHEqjz
r+aAPQI4y2gfvLZ2k6AuIioNSECBglE++yf9zaBZ8QFbe7JokSJgAU1hU5OtWsMm
pPydzFcDcBSdXCjFTQwlG7qt9/+O9GTF/FsWh3OmF3UkX/xHyLrSZ3T44zmZ7mdi
Ew0fy9WgaHOIL7Ro33PbYMScSviVbCMAlbuayFM6OiHEvfab5gAE/UfabaqLk/AK
ZZwfsgEjbulBGj8Jx3890uwhbr92rjwk9NxMTbNUucuySrV5z16FA8WawZXrXjS7
TeyCekmcyODCc4bak6jISMpB9dsduOu3bJUJiv/GOSOZRDGHMV9b6SIEN+fbHUtI
8aqxPRY5dlZERUXUdqqnCTUm0EUizdz88VPdw/0SzOQYn/YqdcLUbA0hoJ2Lxzlk
YjxZj4xPGeiZWsgjO7dmflArKUstLzbTIHaDSoJhSt5yZeWnmVjwsYMQ3gpuR7e/
/5EXhAZIYKWdm6fIZzkylZ0edJmOfumQL+HXMacF0/ekYWLrpRWS5HJvTC6sXDgV
qr7pVsz77WfDuVmHHoEcdha04HKALQL0D9oWG6YCFEARiMaB4T+jmdtHMCo3nXlU
ininkA1PcwdCEA4EJsNj84xXpCZA5Vk/lYuiuTdt2iVu8oECeB/uHbNe56v49d8Y
RaaplAf7Mpo9M2VcUpJ5AC61ckr4hf/g4VFiISw1ExFRHFQ5AUDJ9C0+TcmqsJ3n
1Xy5AtgP7uEUd2r38ygO+RyOPnUmpQyFvk6v5EisKNoJ3f/Op4d4wECZwNa3tTV4
xlnLekFMcVF9rLGwYwAQesWNjKDw8CfXRbmO/l6km4t9KwUO4LKMlofIynOwGvHK
sXgWUagOp1kVx0lAXBvMXPlwkbJHa/tsy8TML/9jeya5WTNVuPgJOkFkPk9gEJD+
8MukwGh6EetTxFsXyhVu88oLMFYpEcjTqbUZ9t98k3sp2V6Orcc83ur41BzH6o1H
jRXA1+Hxozo1Us/PfczIV2p5IGKtoQpXm8O1OWE/U2h6AkXDDH1xDlV7lfwhqrRc
EJTiV08R3YFPU+kHYSAaHBHqC8t80xrvtkklTqA+d6YEGjYJQeCOm9s8FdENcWQF
RxZ7fma1+bQOpNuhjounZ5GsOv1wftPXcxccuBUONchNZgeCbXODNRinbxFwikoI
R/RIw0CcS8KI/vRsP3XMdR3s7w0WwCbwOz4sKuiy0lNmgyZ/pj6ABPjTy7LA2t0s
uqjq5L5vrQZokSu9yUMDuyve7eu0/YTeTSLX8R+n2Ur4STZqfZpvaNDuzq8zbGcn
2R/flZKXhlPRFwYWA6HVmdIVY10anPoIHi6h7x9saW1Wg6GerOKA7SvKJrWEHxsz
xjiCtbmj27p1gpRljOHLLUgkc+DBVu0TJkLQeXQsqx+XO09GvrseJycSDWuFF76M
H/UlAcqk1YYpXkGGa5QLT2EpZg3fGHXieU2gKouxGCGsVWHc+TGdBExF5ZnnTO1V
RiL1OgKxkA/Ehswn92dMqVI63+bDGwdEOxdhKj+nXoItC4j10uMWV2ceMOAAeo8z
Kf5B1Ag/kVOYDVwblNgXSqFmaMH584i3KfQ6KbduQWsO8cppk4jDjVX2Arh8teav
Uto4rBdMQ650bE9Xnzg26OJ3msmdLdDPp5AwH7hNdoDn8R0E/mQYbe0CP7Qmpxso
48fvvBV+OXzZxA1Wz9YKr2IRSLgPRLiPVOPrxWdZuWN2zYYCT07w31ztp+rhlPCE
WJ/MXpGkGC5qUv6C5uYVQMKM249Fd9USEqh+s64c0V+lZ9EjVYNm5iepjsghhW0r
R0U/eqFZCqolH340I8C+ZzGKAyc5ypG/V8eOXlIYyo24YJ0pLDyGxRlK2w3tEF5C
/Xmx0Pepa0tyYNx8Sjhk0VMToL5IKTMWM9gCj0SNWR1Crk2nr4Q6cuwndxDJx+XR
nMKmyQW3ZsCO3+8flR/941k1smsGR0qa4h9PST1+2/w6ONxlm5jaMv/Y3NbESJZN
TBOpdqijLINIn/nrvalTbJ+C2Gtb77GK7/TuOIOKJ2recW+2eozkGP0Qc3ED6Lw0
WL/TnTV4NrmQKKFMPqcAy0IYn7bTpe98zwntb3/cWYvfIn0THBXLAb5pqXxPl4Vb
spUc8YvPVlzALwQoslgKWWN4HhCNhgcEsRooVjpG4Snqm/wox6HruZIT/w7H6424
Nic6UOocp2fRw0o1u6KEKSwdr73LpZj8Syo+aKaikscFq+aLG56tuMQFfiS5rptH
OaRVY1t6eNxgrbbovSLtTt6Zca7wdELMrkMi21Ko7yioQvdCVHZ7vy+kS72kyzDg
GqNLRAiUJzIK7pMEru01L2GP4BfcCC1HbwdKKMyqJKdLNGn3RqnvuFXRGE9bG3xw
z61PA8S8/lJlUNXQrgsbTMYIsLMDXlCNvKVpsHlKFAjGCOczb+BBZvjKfJczYI93
x4LMw7GDbMMrfEStki+UXFjNPvr/9KliD6SqtxRwrDEvWTghPeLKgewqwYb9ZwLx
NxYUE3MmNUALRpM4zYtMItRMAI92h2RKfebRMPK4G8lG7FBZSPMfaLA+gAswmcph
ZxYRlRP1DOtoTzbqz+8+Mq0NYA+Ofuo91HIdTYWEd05PSrFTKQEpt0LHE6SfJ9TK
GckM7jZEkpzWxPcb79Ku5lw/UvsNS64q4jrgk551+WYC6S6YNMTgy787UMD6AytM
+2WbBeCiprDMwC4/gpIWZbZlWGYbVTrf1QuT+VfLdStLEhU/oEe8XPoKzDpvvseC
YogxPAEyKmqsr7fnUoAUkqPmVw0TeIF9zTkRwEW7UlVnabkjuAUXKZkFet/xNlaA
OP8Sz/vwY3dI4Ga8MK5gc7vCNqECZgeMfo2e0KXw5Fg/wF8GRQGSthX3+rATn7bK
0ADWfJQ7vUD+nMBuTgwl2sNDW7Xr1ufjLnYg25AO4UWWZAh+1XL1kCkzAHgVxCKA
XCpT797aCTHvCbUz89Uq/82/CNE6Q13xEBHoMMEgNmsQRQT5VoZ0yeFfPblxNdQD
iUiWYWN70N5P/cLK2+s1hN8I3H17liPCTukIYef4nS76PbwZymxnGqGdz6c3uCYV
WEeuW/9eWFP3vS+GucQ6M1+VsaX06Vx2T+iMfo/RShjNwal7T0dOiLnM1TdAJoOb
w+Sv3WPLgCmw04Wc07n2+sfKK1GtfqTkm5YRJm8Ba2nBQt7jY03tVUcUlgf06Ic9
pCqcYwI9VaSiwGAZV5+OnbFvrSZydBo40lx5zAInkYOwbppaCOzwlTYqfTh240GH
uQHbdyrpjPXysrjp1iyW4mJ9tt3otHipeYxQGWJXNXhHExaKselfyGGCMpzAhLgd
NuCLMulq9Bkk3cC8iah63+R6jn3bXrDPwib5HoolYmR9Y3eovj7ezS65SeN/MDMR
8yp7HLYifLT+MFzrINaSPMRd/UrUY5SB+SA9M+YSVbtLSK71yLaiiC6tpniVcyRV
ZLcT7fHamgWln7visRecNGu648G2+m34oLW92fsHLJ9fHYGJzdNtVXAzqWTyvY0q
jybBGc8vnHjcG+Z6SKfNg1x3O6T1pUOOiPGdhy7aFaYXiINx8JclNYZXWumu96E+
6apquifLxG1TzZW+cDqMy8Npl21EZPoOnbSujFnLwI2wOwntzEI2lazwh2OUBWzJ
Oc9zkN3/FtwlV69p7wWk6hkgKfLVtwKWGazkU3uJl2gCwBf4s+2mhv4K7rZe6LQH
2vaybI6qwZRtUsj9L+DOScIHsJhw6cg/5kz5h0wkrpZM+rLUEyksi0g8wFQvmICD
fn9PD9J0jLkR3nNcMenrE/SrFxTJNIxQpeohV5qRwb53hd8W9TOYVZNNYzqHePv2
3A6Z/p2YxulPZEpWBUCzAXFjb3jhRoVSltPVU8MfH7emrmfrBVcfMTsAYdccBphF
mkGwuPyNOIUU+0Wydb1H+KxyzjYCnQoLO6rOUCH5s2+OFmjktDMPz8heoleKjgpj
6dseXgG6HvPnzEBzIKnbdmaAiyulApF9iATzAqpZdoX3rlwIiuogH51TSGJQBWKN
jdXZV6YU6EpTWD+oIVicx2VHcfKucwNjKvRkiusOzzjEkPS04esSvud93S9R8esh
iTEn0cQ66drIB6k1/rpQbcjz4rF/oZ87ydrhBTSwaNyHr0n3Zju8F+DK5GZvRGqN
PHn7JXnNHr/iTVf0JO2RjNgg3AlI/w5iDpUg5+5sqZxyOValoYGcXFYfrEJHTuEu
okXnUF1qLEqsWwHZigMhNNstU2s3CjAe0lYGgsf6k0bEeH+NDF4kNLE9VTzxxvkR
kSo5cidEW1bIjzB35dZDf+cNlrQnEMJiol5SkMp7RcztNt8XtPoBwmZ7iSmz8CFx
pgSNNBH/hvflfQiFkjijIGnRvO0BPkZ7g5Ha6ksb4sUsQ9sAiTW5Om9sqW/WaqQD
rXCq/y1/nDEWJRknaVDM8pV+umTL6Tf/Gn996GDLWEEN0T7q4v8RojFDqOKldW0z
JdeDvm1pAk9ORxW6mJutLo2QvyAp1ceoVO9C0egL9O0v9Z2+9nS/0BM92CYwE+xM
Nz1/H8kzNyhUXM5ZvAg2RU+xm2Y0PJs5CtqR1wlPZE4tFAimLzz0dVheeXKKPP3m
YVvo4gRw6WtdEVq1spCHjTtib1Q3dw5/v0HnZh46bnFBfyTpsj5xIf8a9riguXl3
rH/8lwF511Xuz+sE88SCJe+kYjaJ5/iaNAQ01oEgMPJ/qa4q5ig5fM7QLDxFZQ0a
GBcUVkJ+8ftEjLqme0wrj4rs/rMcQuS97IQyMh2EGsh+oDtTvr45YxQzpnaDNh+p
NSs0h9xBvCe+sesKV0/VnZBletPZOP/r+izM5nUi0C1MEZn6hPshP+alusdURZ7b
pC1zDL4r6hwHKXaNwav/U5mgXM0SmU9Np1hVAWf8dXrN19oW4nQHu7oGzT0ald76
S6eMlskwXskfEc+ELqhxdmwq43dKmguxKnjWRCuMzZEGNzp+MXI2EaeET1hFCJKg
LLiiq6K9lDUV2sEAJ/acD4M0Ortr0FL3zzWXEZClZlTf5rKQ0dNPzw81sPDVLoCW
LyPeINPXfikJ9H5Pw3urAITvjCBqB7PHBym7miUJgVjC7WW1/UK/ozWmhGx2+svf
YNAh+InRYX3033aZI+hD1lfsTWOv9ebCcFtrzkMmXan3xWvUQE/GQsHq7pA1LCPJ
BX8hx6bix51wgO3jXr1zBjjMcSR2fIAhhcIqDnpAlvCBjabmrqp4pssWv+ANXJhf
vLASs0BGNJPUovdWjZCMO14ub7qGTneLXkIuoLGFTfwcTCd/3dqsqnysd9f74m1J
3KrCWZ6qUEQ+MUQEANwDjbjb7bOaFKNoFgmrLIGeh5s4Hj651cpEX9RS659bWxQh
adY99EIdfMkH4WKGoXbAN6+QPu7vsFRN1ixsbDr3eAGgob1MrnqggmAc+AY9CePt
azQCumUZC2HgGoUR1DTF9bAHvm5S9Db3MNf+yapPSfpxvGaoJWDrntKN/LQs0YWj
D8es0Iycwp3RX26kiAQ6CKpss05ZBuXh16mBUOgrahewMvB2n+TQK+Mq2J6ItGBh
kpOiwV0qx0D1zbm/EIDyjSg1iHKxPSrGrzD5Tzea1y1+Ye1rVvsrSaQLhzgtWK/F
ETwQT+f6vIqtuGtYp8bLCVgIeEWWmTd9BjD1e0oEb/u/Id5Uc3XOn4OLpUSo5rkS
9AfOINCJQEhyTtkTfsC5+IupCYUf5jILbWyqmEcxL0B2I8I/0Rnjpxng2rFjBMSp
h5j4gAbz9eHQpaHd77AaIjm33MZM6faftFoXEFYQJJ8Ac5FCZycl04v3jEtP5CBg
zFmzKgeH0CzN1Vy5ECfw3WYe/54SqkhJPK3QFJL1EB05L7s5eaJBewG3tdbFM3bh
nE+tOm8OSBLJkH+jutT6b5W4eyapzZI21aiXNnDB4bNEwoHxXl+Y6LTTvSEnAqQb
H9RlIIipvmD/MVfszMLaJ2VEF4s7RRwVmC7Tm0emFQtSjNafNxiNOuyDM0Fh/J/t
6WZKT8aQ9duD8o8s2GCEiMaOmnmsLVnsJSo12ojSZo/xFOAnZpOX0knEi4rIwLvS
Xnk3bH5+blT8ONO8xUh92mY9v6OXfVMStLnkRnH/cAkgqcrN/Y2zHIiFSFOwvQLp
DlR38R+crvWpNiLCNONGRY9+k+2oM66krHK7r8kCblx3HOl1H4n8syk8+waOxH03
/PToX04PbLr8c75Az4aV+fLopIroRRgCuA3dn2J1mUTioZngMAdAbHfJA1FT0mVh
BRmN7++skxBZt0OV9LXo1uFdr4f9G93Z62bxhcShW/qacLY3P3CgGR6A0zwD0wOM
UUd0wYk8DbZJDl50pkkv3LQKp8+1nd+mi5cA2vInNoEbKyeX25PU4SgdQLSB96dc
EuNO7p9LCJzj1yJvmESb5N8aP7+cuPxMTHOIddj0Hp9a7L/akc3QNUB3CkNm2XZz
2Yx11eij0kUNxT+J50tN1VIVtAC5IC3zsRDxJj8FQd4CGg4FRZUb+byKoKBNzdAk
fGU80rOE9fEmOJ1MZyLEWxPLlQyTa0+LCExqx9Eoix/cbsQ8dtrPCVZsHxpzxKfU
OiIP3fsC+vCgbVlieMnHs2GEWorEhgi8i/C3BjTtZAkX7Vreb8una/Xryv0BODkR
KvhfRyuz9l/In/OJLKTN5ono2Rqt+sNalc21HirCFpbtrGceTjtJAcug7BfaGsas
Mwe0+1Kjh+V8vow1r1RBslZtkyJBCCIREEmHWhNu85pDr28oXDjuOvMSVqCML903
BUJgNUeNenVWKIS/A0ojtYXmoulk1Y2HiRu9HT6Zp94GiYhqN6FNXpw3y4UKWilL
P5+/mBowbUW2hoGAxBkyACM+w/mlYCQsSgji5mBRp07N/4a4KVo3NeHlYHzASZSC
IiAFePM1eaoesAhz6BOrYaH1VovYbcBT8jdu8QqM+U9U9CGqXjRSAp5+bqDZQ22x
90WenZk752Q794ZnSRSOYRtHS7rXOFiXwQrpvmLzIPY5+ZoX2n9UwioBdp0SVb+0
q+G8Yci7hL+QgHNRhxVTfmtTc3EMZJEABApW7VuaV5AvHZnzCg1vuWFxh3Ebb8n3
1xuQV7n6FRqbIbPQbmv6if+O6Ujd5/sbEK/Mnx85kM6xcW3/ubXpgN4AS7F8gP62
bZD8ODrOR8VoGDvxGcaDrd3r2DFc47btTu+UJI/NMnMKUy0G42PBm9cNso8i/bS5
Qvy/9gbUmTNi3/u21twBMNkGNFn0xOOo/v/R24X6E/LYr7CqCF7NikxNykv5cSZn
1RSVnHhByOOOLt97KDnUmgcYAjN2gvdJ+dXom9xMW+tJSuoo5NRycbLWabxu3KcR
icWS9dhbk3xV87Pu3IKeFI53G6t0MJZq12vVLO9OUnffNB3bgXZC5mQ3BjOVjUFk
nJGKvDzZaz1aPoC4vLOzh1OmDcHLNP0fn0oRxPnIw5Vh2G+hV8bzxq6kZ8y157MY
WOgkJzifDXw5mERr3iUK89BhkhFszLYT+WSkt2jG/4omqRHIQ7IhmvpByPYAEjNq
rtRy5LV8NThJaJhgBdaVGHK4LqdrSYZSVd7bbnoeXoCYpMQxba9L/ez6SkCttP+9
+otX/kD2u1BuEBfr06nphhoyuMkvITsfqHvfinxDE2rEnhgU666m9ZHkKMljdyQz
J/qlq8bw7OpCTeZtybaCgpP4fYy0Qa7DKwshU5BIBAMJtkwFs5RPq6bcp649Fde2
Atgw0UoDqWGGUFY0c0A4hutuLqUgmSQtv8rGZvBItp1KwX0ENR/2QaAQjKISzBv1
QlHlb3ZhyUCB1BYWOdmVBF8AUZFvBns6YCgWcYKF2Cxoyp1MjLSfHbfz4OlWXLPd
3P6Y4jeE59S/9gFl/idrFLw/p8b6yUlrBmmNrH3sYZx2KAQYB1XN+e4gIlVgr9y0
HnMqCasI8+pWiJSr50Bjgi+60THchWKM9NhFb+j71TPsKnCcG0zOrtd2vn+XT3Qw
GRIJCrbz++Zoo/2BhBvh+yCr+cFz2P6YYvoM/b+16xjj1fsiBBpkCyUVJ6lGyrZc
qhvg0Ywsb0FIQ0ZCnA3vGpnPTeJ9eXzC6gzkHWTBTADsz5hW/WRJbLmOD4/8TgUM
v1EU4sX+Y0++OjIbhOtPWH5GNAMIL1bTyEkMGzWex11MCthNXlacWIRqscRpFSrj
V9HxpgvC0CajwhB0cK694rs23S0UybSPezJHEVpwSZUn0gJYGXVq4aJmeFLtXsre
DH9OKFeKZoNkeL4gOsvrU+v1PdyWD27kHeCZGvg2dD0tvz2qbLzduQ2qy1Nx8LDp
RkUilhbTIEHje3+M5s/OsMwCphrkqZzEOLIBjj2nriLZGXaaqoJ6U9jww3z4mmmK
itzGGMaAJZrRxWEE1q89RK7F48edSiAlklQRfv5M+MsoscugAKU/uURl2bHC9Qmf
3oyy1Ucu02hWBypLP6W8tWjJ9rL/3lBudWzANAS9fe4kVvbzqw+qEhbwohi7OMdI
918Wu/OIsqEk+MlyFNUmcF6TmNp+UNOpYVnHdMtQO/1MBycGqA7ZleQH3qoHJj1E
T4VZK48+H2wFi89eJiZG3psuG/O9j6bYgWRKS0Rx/FBcYOJd9BMGmK5denugE8Pe
l5nRw9xaOvk+FqllOKPTqYxKbA4LiBK/6Rk8XtiaqVNUC2WByu0ExTyuutfuGM2t
AAyol+V6YJbUlCozt6cB6vgtv34vyRqWjV33J+Xmxc4Nd07RFE647SsKT+UaMJ7M
hEJJWdiuOAR3iks2CVw4NVzMOn9RWl4N9Jelz0TY0R/fosd1YonP2o977uKy0+R/
fYsoGtTP/UZIaVUF75Oy05inWfc1QhUrpBHHjTxylRy0oK9HhvSo+8aZ1d6X/nQG
CKfBA/wdwZoVG29RxzoTlOnJ/Q3/Z2PJOzHnAZgSENVc1N2kJFqfx4J1fzu6wi7B
sTBS7uUWH4M4ND2AfJYx/dwxlSnb9yI5J6xCCpx9U7qYxGpiAnQBbrO1YRliTtvm
q/aCwldDTGe1HJr3FBMVsKAAezCEBc9yVssMvv1k2cyhG2ET8jtVZ94cinUIATwk
vV42YW9mrbMzcBQI1WO6Gku5/kuwgeFaW4vHZiVBFeLMkwJOjtaYRHwTLlLSO2+T
blc4ejq7iKAlQc/FzhC8g2E4mL/lfmYZEivUVy0eOfmtQDU2q94V/YYgQsGH5nyP
vKetXQZ3QwJVMD3tfneJPQaCS0HoAjb+3sDNpAjKXFUWyt+iWwdqwJ9QU8lp8BAJ
+uMZkPgaeFW8ffg54/rTFZnH+FSOWKqJlca8hBOyDCY/oiC9EjllrSJh3j0AoxLO
OvgQRUMddbxLw4InTQSe0v5jSWMKm3b7iWyNeqcnLymuDlZchB0tIvQrkqGDZvxG
7S0SWZtY08GpSMB1Q7j1Xrz04pKq8zjFEKklpk3nYVLooZPogqAvMlhGACFUtzsu
xdn12fEyu9rpWFEaRS55ENCkHx+aTrl50lde+B1SPl52gAv6s92D73O3IldIDCzs
UEp8bDmBLSBNrvrj4toj7YN1CUZsHrooLWEdl8O0HMG7QQ79LdILvczAyyDjjnUt
ppiMnb3cne7mWgE5hlJtdNPcb74OaM/V5fdpBWSup9wdra+1Mkjcr0cErR24hVP7
UVhUGlxJGFMffpBxV/2iebzmxpNdBN5qHZo7IvfZ6QNAgz4Lm8GgDmeFs5/T5yZw
1pbGpoPWbqx85sSkfVz1vkZreKASgLSRI2EpG2h0qNcuF8yD42yLyZRhLEE6dSdK
KUvgzLUdXFNuql7JD+BCbYuxJBYqGdawLmwKuivimZBgEv7cAzimrBlDLmAGUmBU
Pu1wLh652glqH+HwehCBONd/YdDv91YVI0N3l2y+y7GRBqIVpLMNo2w76dOOJkbo
p0fB0svZU/iAZBlG4d2ixCQiavwY+8RqvS1EQHUNDDxvCJjP9I/0OLLal1omZ0bh
Ccare95W+Alk6xyCcxxGPTLXYM9zhvnEJfAH88wYrdVmtNG83nEU+WpQ7Byul10H
WC7NI7eVhblcIUFfoKfGTJeAhmaJbRi6qN0ypFqR9pjNuB+QRKUI4NMDmzmIzavQ
oO8PJbmdJ5Q/+3IWHGFNPd4aa4j+pP+xkk3ER1+7LLBCqNiS74AfVQVk+fGKcsbK
iqaIwjKTY+zQa9pUd/C2s7kHdrEzdXyhKCtZ3jvuUkNzz5AF+Oh9R/eEtBBsunmB
bg/Xh2rZQ6VOtEG9N1Cu454Bx/Nsi7HlVtgm4JU30uOn5gVfCi2hR5es2aAG2IWo
ulPkC9nC068KClE8/+xalriQSggQeYRZWSGZy7JxwEMgP7MhPj3wEnhuCH7T7/cT
yGxt0KKP8LsEaN1qEsII0NUPe3HS33Wbf32woasll/ti7KlwxuRdjmAKzrLpY5eh
EmP69cfCDbaoebLrTdLZGzTaEv5vFFzr/13HRGrxmM3Q+2xIpN1Ysg5t80FsjdzS
i0OdmkatQGeZ4RMXWFi/tOzvvysXjpMTfGecu1Y53YDQz6G/7+YFiebZUlmaK+pn
5ORXgrELqxKvAuO8iooJrRYsb7KkMdWZe3X3f0Er2A3KHf71BVjFdIXu2pY0JLgw
2NKen1ulMHry37K+4jLuSp1tGEGX1pglcg+uoQYgbUot0DQ/amxoK7A1VBFMevwx
oIeLE9BsLuMOUZuYZHlkvhKODeCzFtprdBIMuocprRG/GO3FEwRgNiKIvGCoyRhL
c2g5kM5rjeMpZ8G65OUUlppJUPw+R7moBaSkhcJtwJmcBFX3eGUoA57fGkI6u4hy
/H6P3Fl33fxPIKQM7wZL6Iufq9D6V2uGnXHE3wFNkgYKrpqSf7rWAQpXs++rOBvQ
ZWxLUntuBn7ICSLoB1bzDsT4GOef5uzU771aMXM9fQaferRV835DklHG+RD+YYhE
oq0l9HYnFl7JI3JN53RFl1tAoHrR8SrPRNNLL/6djRIBtlP7R9HD8JUedXJ9PkpF
IliNzRkQvfmNgRJfbZw9A4Wuz7d4xeENASxV21oyezI6t90iUxbJCsZ+mTbDqIgR
ku81Hn9RV93A1H1rNLFfGBaRI4t3tWJRQL2f85V7gZqT/zLlF8kIYRMvWJxSXk3X
Xs3GqR25oqlkMUmTmQFGpM66iqlNDrXD9PZm0byU4F6NDXONHnqhQ4VsYJfa7ZqP
Hj6qAywpw9sx9GGCGI8NiPXQX72ZPImZg77c9UNRYEeNmchEbAlxGjkUhRy2rB19
sMN/LGs1uEiAoDpzU+KHo8tgOliqkibuQu1GlHIxGDyXPsG90HbBjKopOMbJByQI
bzxPjXE44OrZpZxjR7hiibZiK/RDnIb/oze07L52soeNIu7SfNz8E/EvLwgBEGwD
6wUs5PYi0V5DIxIoxU98WK/YOGXv9DVmUlCHwPxZ6Tq1al6tSOez2+zK2fKy+87C
WgpZcSPtN5Fys/9MFqKfI3bUwUn2Wc8jj5Pd/JE0BZ6Q5lTLKQ6Nj/U8ZVE4YPjT
k9gJyUKbouqeqSeImqt6cfeRVqQyOeJHdg3ap+OcRVNjgtK6mfYBHeG33kFfckTU
XIddCjYYejGaUMyEPLd17vjcc0wjyPP8hNydXwlpqYMmk8OiuloiIub2w7INLMvS
67dTCb53smyZvN43HSzNdCfn1F/+f6LyftpND0ykWpuYGFFy4Bw0AvEhpJtkBFuB
mgNq9CCk/3DIR99A1bajB1l1bdwV1dXNOAoXK3II8JE8jlF+xLX9NN3tRe0A0b6/
mlLmcQeCC/f/L44+E0g6NKCXDfErr+0mS1MpD0euZOS11uAnrlGxXSIt3HT1+CZJ
6nJjwpv2fs7kFrjYkHhf3MUXULM68Vzj6QFJynPZ43ipFg5gr4S1hxyL5cV1dS+d
WC+vnkqOAQ7UYrsgne1XcTQbZ4YOqHdOiCjENEhjmMM4QvPXXDsbwNADEX1r0XmV
isf+TH/t5XlGeF2adVfYBYWkIlbW+KYKQjm+mbX4dUveEp1/0rzLHGrKPkxmpzkE
RqUf0aVqWFEXCm5twBQaPoYySBKzoFSdFCWwkSzNHC3pgCb+moUp9KqJ1F6rWZRO
n2MTvcVQB85qL25rThIOisQTRWHJDKp/4EarOi9OUu+QuSUZU+EceB9yXiJT09NT
tv86d6G7hnAPhnqZ/j4b0fEQ4KjCRBMjkECq2kvbtTDftMAPJhD6ZfOtaZnINFXt
49N8lGH0sUOeR/l3zwhFXE4BfuUQ8gbl8xNKRgIwTtzlIEgN9C5FqT7NmXDmERWS
qjqrvv38SEWgy0zNWK6ri7FxWwvGe2IIADvUS+oet1N8gsRe9EGJkRVkBeiFQXLL
KEaz2WR1UkVyldvjejimK9KBwygnG6jVyW0GKUBlrB63pgdn223XPQ4i99vuHU6G
nwBVh2ZbyqKi6cGpvWENAK3H6sAFUDBQsnAXoHkck+d4XKgHQl+LgaiCaaHZ2SZZ
bOE0rU+xcNZu4i17D8zuFbS5R3tQ0Ucb7pGdeRHGBicqsqZpMkrsOAGrrHqYtdPk
/Xe4Jd+Fx7PNFJJPL2bXWNwvhQqsD6Hsb70L94eF/pwddzjiJK5kHgDFZG6+789m
tbRLdpeG1zJWW6UIOnF4Ecbl7nbKTmzdB54+QNmQ/kDVorzW7NTj6IRDhgofbFQq
D5YTbGKfSD/L93Wz+cf9d+0GnYWPanrFFOXKcmvPw+r6QqrdcvUqDoNUMgFMogj8
I+Po5tqXTFahwzIZub3xeckewgrHQZaq/7WjyY3Y6uKsKRYSdHQ72rqvEBJPcW0c
ldsk/FXy6OWVWzdgmMCLjowWzcwCnx3KP+bOjbayM80Dva1Ix0t6oOhURH5rWNnR
Jci4E9+AiaFuIEDk703r4vUjvvPFeOHhjlSJKNVLUMK9rIoEKMGxzRcijJRxC+w4
maxxjV+h1/3IQ72pEWaD6aMLp9mtHaV/uZmpIa97Kvrx9xeADLOz0mKZJz73DOVk
I31mwRzi5q1xeCbRV90A7vXiohXYqqOTDFHNT4aJ+a0DTtXLtBJDZMJfFC+Th7N+
pUuP/pYvTQSIU9rcroACuLYwBQtUV09TYpRMjA7Pmcf1041Y0y/5D91Pi2IFzvzj
YvRxNwp6RFLE8TIh6GhDI9WraE7l5EMcTjnintEXTaD3TGJwQ574UFat5b3ZMjqF
LgnjH6r0t7xCsbndKJzpGYXS1P+4y2C9X3ckIG4cKZyGb6HK4/bkvFvBrQrpGegJ
tHYAipn1P1A/C3Ekyy1nyftoVPXQvN3Kc0L+spqrVv3odwza1eMRJF4N6VcaiOPU
Iw5VQTS3mktqYYnOX93ci0G9c9ExOyArZBURseQ191fOD0slGo7KceeyXoP1ScXi
GXoQ+IEYrrXj1PZUvEHeel+IsJY6k3wrvyaFsKmwI10GnlTxxc7nj3zN2Pn7KzXZ
NP9ucwATPV/L9hJ/SyCQvq1tThA2kM33Y9mvzZejisJ2QCLVpv7zLlSsXYUjMKHD
A8LX/RWlT6+ztX/aEmwKglUk5ZpN5zk5DMs5hEfV0qdQ3cKFY0Wj88BLO168LXP0
3yDFacZeO2dsfth4HHKicx8eao3p3/YRhweToemWVkRG7oxyIuXf8Uuut0kcL5ev
6PRBlE7OpXGl2rL7/7ummAsF3K2iDXxjdHyoKcC0lr2aSt7cZxMC7c30HcretD8N
jf2AVu9Xaz1fGspureW2x41ZEWIVY1n73kGgRE43hB0VDrOIHJTuaUedyZHfA8Do
N+GKBEIq+tnckc3T5x+/wiYS6XaH8L9dZ8ikBVdjhqxN5zQDe9Uhk5ta/ZuBv4qq
8WVopsY06fi+v3sbm50hrZbqhBP9YsIrZDxLmspOj2H4EjQSPyUzeElZjY5dgPs4
s2xybbiD03dw0ReeeNyifHWpIc8cM+2qwqTrbM9ce0k6x0quuRtnFkXiqqhRMtYC
ChmCkYkZQjiHN7S7V/uwRdN/esA9rkDHsWei451C7d3VVvCREko/iW4Yo99BsQG/
YmyhrF/3Hg2hwmF4qU5hDQA4SjQvAhwavkscmx9YoG8uyFICHGH0aJiRNmAmCIE5
mWr9UZffWc7Gcr4tiZWkyYjvjsA6P/y0pVzif66ZrjQiUfy+eth+tkPpGK6xAlKF
F7ZdCxWXTqBk704URnd+QvqZ5AhIZUvEN7RYvtN9N9Af2SzSUv+DFqdlb57MC0Jf
X42eWzZgp49/hb/MqXPUI4KGYGJFeKh52BOUKfYGy6E/vxk+VrwswbnEjrpJ74Xr
exA3qpRI81EjGd8wd3DztpoTnr39lDj9KU6Ru+SxIJNEAnEE6rKpS486O17wnmoA
Vvz0u4mQm/3kt2DHi4LB4TdU4bnEpiZmelgI28PZa03aVfCXPvRZ5eRyRy+7yYB7
CVXzyoxqQOncEx1DjNNqJ8Lv4J6pdU3Ql0gtfcs1PinHxx3NNuytjcyzBUAZS3EV
q5gwJIIz8Nk7ASynOhy7JS8xZcnDfokETEza5vZM/YXfd99u3+rb+ZrL7aZoHnkt
8gLtFGyQFEMqOG13tedT/Uo/rzXlkGLuLnRTLA5PfkExMqSvEusl3lZ5cFHv2en4
Sm48nA9+Mftfk3c5wHDaVj6ZVnp+ao1qTgPH4MxSXRLgGqS3o3UzmQuLgVILdsZg
28BOZeK/ABlYgrfYPOGcTI4uRTNH22suIjdskp9l61Tm+BjQ6AVIr1LI1WUdezHu
fjW996jU4X8/mHQ7kd7gOQkWJi8dhvOwrNDCxhp/OtDNLURn4dbbGcLe+qsEnTYl
l8qUfQyRfqqK3HV58zPRBU7I/VRF6bSg/GJ2nGnwPtxABBWGXHNKOyIdrHB85yLw
apqtM06kJZ++CzO7QUXO9xg5Cxwz3KZXw1OyVeCit9RcBNlL9Ua6Tb88CbuN9t4Z
EQFHJngCW5NR5ygOMb1mgxh2jXMJzYO1CcmBCIvONHuJbB9gJeZCNIqdXuSJEPjD
JRJXa8niaSNPGbGWbjtuO0s1LWFN26HtPxGVy36I7tHLsJSxSWcIRABwoB9e1y2V
gCoN9SM2BSf76V57/L40bwUtQVbYFDR6Wvfp/9mhC2epgU4VKFLMaun8j/6ZJErL
Nkq+W4/l+IlC4oE1DdCZ/5S4sbJU1949eoZbWqUXzqku9AdJ+ndTgVQk/x/Z3HLP
jOgBcD9huXY2uG3eLpMNZZqfei4UpELyai9JNzOS426n6+I4mV4pHy8fQXlnZG4G
zUgSXEVz2QVSe5kwqIL7Ly+wCsL+0aPEfXSaDxsQQVplGLrHQOo+1b/e1AoSVJTX
6TjRbhy3pKoVWyNtqjNFjmxT09iO1nVCByLdQwUXMQkAi4akcfzP+tJNO0OYdvH1
mbY8y2eWKktu2tJNhhiTFyJFV6A5n0Bs2e7n3adZzjjHY81IwFNtP0+broGwbEqu
dSNMRB+3X0wdbjutyjN41NU7UwgkQmwtJ1h0LD9L3OK/eRVdmPExxiU4ivAqwF0t
oumHUXuC/J6+5lCNwKTmnHguOKGf4cVg3QnxxUcKjvM/vTyhVbFGdzsOFfKymVYY
mpFo5oElp3RzV3W8kdCQFpHnpKL3sDhANJlN0Lj1IcI7aBJApGoN87iMiiM64ddd
mUUuZru6Gwe4cdkkUhZ3VDSop4+m0ptGELbL8nJdRajUDOC/3xmTibiE9v7llKbb
5jmKdAHA4/KnAsaqXe0Fmtd+QMWluXwcuv1ZpDSgVg1ULivUMjoh6W4jGBKUmW37
LC0AEBm7wDMzf3CpsXYT14sYliXgTcDgTvwbUtpgn2Mn4nyILyXVjkmtyjl3pcuc
+QYpgadE4whNh7rOwsADMMB9xtI75uRjXIA5TlOKCp0edDo/52fPWgAMpB/pkmdU
LFll8cm2KjdnPskBWxX22ki4FjVWIbk/6ap7Dv9dQQIM5hT/F6QotP8b71tXzyCA
19pz/z6Aj53z13i5UWR90PfMPJMvcyBIU+Bi9AQnwJwgSd1VnloDG945YeWlUfqh
j3U55H8yXT4VpBBthHWKjZZgBbmbnLEn4L/+xZ52pZa45zP42LaGat1vTvOMP/7e
j39IrZilwwckAIkT0dl4UMK+0LGR6Wq0WsnSPRyJuv8RL2UYQTJ8ALd9N+QYhgMC
BfRxTBTpo1OHf5H7CPBg+Rcu0qykEwUOCkMEwvYGgKfcfH6sMRvyf9SE7aP4AzCc
RPT5au1t8cTaLj13VuF9JXLHsKme7mEeMblNJ4IaD7jFTUdQt5ag0B/Av53enNRI
EuURS9AczPHK6MUosR/B+CxLsuz1GgRj06+Bv3mHtDUFznVgCYAiAY1tY6qDf3Vw
wWpMhjCCX7RP4OflnNDwnYycquOGyTj2SO2K90i3Xnzy91YDgrcMOWs4wOV2gkh4
xsC559ymNCkBtW3jRN910w+sGsB9mFm2B7TeiFV5bkjTpTAzYKYOFhMKF9ZYy6bp
hiqy8W9TkbBHm/EDcLMR7IhHksJa7AYPuz2qd0PaRqcvE1P45+JVx1rjcRvPbTAN
SezBiivxMveqySLohISglfJ1fbmRaS4/HvGoXiJxaMdA87iTq+GY02qg7E4N4n2W
gj4CVvZA0bEAFyFhyBMFPNeKsmhq2YTx37qFLJ09zTcXiUnf0tebXXFdLZcf7kGf
Ol1gnsA/9LVBmzVZB+STAQvhjuq9pDCZkWay5rW8+wA5k2mZsUQSj4I/Fxt0XDQi
Vv0DXkILDG+0N9rt8KaTC7g1xw/bDcvfY+2kkUUi/PYTMnsvJbp1ZufMHV54ApUs
JdHZ3MlNCjEEY1gZdEFAWVh3iXWqzEUDzTBbLhHRpXKo8Lu1aobBSoKwba2+XkA4
xkierCD3q0BwpgrTIsGOQnKMyQk+FLaRWVH/ax2rJbnaE6uqTA+5jCunw8GP4SZt
SUuQSZ8w4uSUsEov4VB78/qwevK+WJhd1NJu6d6VvGCgq2xev9LJC//jCDuuBhqt
R05szZ4A7xiVrOcmrw6lUHP4n0z4lYJn4VYYp0Ro5lO1DXconlQ0OPzwkPPIboSc
NZ3/zkfBbRFa32WFQaeZobvZOvbxO/X0d0heD4OC1a3OujV6kEvkQOK/NjL0Gh0l
YsYWe9DfUke5m4UGvegaxCK1ZfPhZ6HaYvyrz9YTUBIwenQ35o/iXA4ZqHdvJTww
RbRt0aMuRc/KPOe3c7v1Ap7nCM7GiWkkwu3DZraaWti0J8O/UhGItIXVFrHsc45f
aSugOaP0CHa1Y1vy6SAl3yaGcfXjQsmAZ9LT3wIbV9kz9TI/YUU75S+Ducv63Xvt
oiG7KQmfwLks+jAUre9JH7kZ5cEicvnqiOT1eTMP5yLwnqZ1wOtN2O/1OcVuYPxB
up3PzgqWapwHseF7pjrGPiwWgB5wmBkBrqxll1kPHTkFylzYlPZ0/+JkcskBLYNk
ZXpcESyTgkqhMAsh94AD8jqwllzcpx2fLsHLj67iYZoMMeSVhefJFKaBW5wlB28U
4vunlNMQwKgzgIfhA1cX0aS2H34hYBfBn/aLakKTsa2yhZiPDR381luVuMoFBbJ4
quV70hvpHSyxFs5FaUWP6iEoqMvGktSz8QS4sQxpVTNNjOyUMUz6F+T++FHdVClj
qjWrMSDSpm+8mtxiwXdv+nXUbA14vQGsP+aK7B1PjP8U/+e1Cl9P7tQn5fmvN0nz
lc0RkI0sexcVFUd0V0XXly7MnJRAshxNXMoXxfaECbqFqC24gywzaIMjDQjXjuN4
jZNoGUKHTagTQKaBtwZLEprDlZPE3UyHy0M0zgOdxhWprOkDCf57gv0q1K/vGEnS
THU+NDKw+bdwKI9k8JshHTEJ20wo++PJpUxWcYbwk5XUcubOx57bAyUR6S4Q4nh5
N7rVppQOJOpeShrzbDWK7XaPpNaLr79uYJKHkOKTjWCgiUe8Fj6SyiyRKhs+lweR
m8eZCkMKvn8I769lPz8z0gwMfwk5Iiii1WsX/SDrPlKeSitVV9h6gmJOUSkogOz+
M8vfTOcJ+N5a2RfDl4iYV8tsWnv0R5Jgiv4nx5FVvJqOwEMYKCkROHexXEZO9NEV
BfNxhBgaQQWGXPuYb/Mm0mZ+lyjI9rsRzcj6zRTVQYHY5ebwYev8BuwsGLGSu43l
rVh9fcYjLIh6gMUMIh6cO0eQ3hcHAx/axo8Jep25Y/nMKj8R2w5pPA6b8DC8o+uo
DWUJrCqfmYk7ai2EBhctuPEGPwJQLTF4sCDJZ6mEewAXIw8dXsKtRPSlm7lPzelK
X4ExOYljQlvlqk/3Mly6qUU7Hz4WEXBFfHu/kl7YDe4dNl6aBkPi/j22Zc9CERpc
VH0NMXdFfk/szfeGm0OEb3Z8xtvKtsmNhTp1IBIMvIHzmOUKotMJTg16clFtKpXk
hhmWAI1iC5X8oPMHU7YrquuSm0PLLkfcExGKQvT11l2qTPbEECDi+Kxx3SKCBmkm
f3fQVDjGyDBjFWGEXrxdd2YjykwIUgEv+bwVZ1PZVOGkmc7XqrTczUzyTy2Ud7yD
UAtOmckSN4eQpCtB6MBB2bmYqRX9WG6W1ORQsohfZ5OfNecQ7c1YGpRW4QJYTfBm
IpII2Mr0PumsFR3du7/kcUeeYq6sxbMWAQEMUKjYEKOBAXnvefghnEJf2Ql0pFNp
13zyXAnfM2+A7i/uLmX/x8O0SCph+4ia2j6n/60/9eM2r2hrkySpiWj/VKFyMG86
rBA+D+pfQv/fl4hhtXCIwZ8blUGzr44+2bEVYZcXDfWF84TmE6LeLHeDgRWbX2OI
YyprfUGkJc1gp4xs9aStq683EGtq4y3tF4h0olS94dnbxZcrbfZCkhpExIOtJXTR
d5UdxpvFgxxGFhqYfAd8G4j2PYVHPfhGx1E9DIqyF5SSeAgxD4NDsUxcWWygCKkb
6/j28YiEPVZXfM0WvIliKpFFEZyP6K4EUaCwV25CcHfxnqHcQ4s1KGNIa6pZwrcP
0wQXVFOH+9ZK5gBrrx/kosreJAfNdtksFTyKMLrl8S3pnxrkOCHzE2GVG66V7jaP
FJijmTpVGEiTfIU2oMFCjAZLeJCtbHD73n6Ax8CdDCOTBdIt/N5qkudZxLvcIkG/
p8p4T3VUUtmCZ8gpxrrl+lw1EBgjwY2prWAtO7Aum1+CQKT7qdxFh1B1V00AI4Zg
UVPzXRABp69hEWF4v9DmS9hZG99/hZ16YXSkMrRiEKVNOrSnz/4Y0lNzWgat+eE4
CZk/U864AtgFBs9iI1+zFnVIJvUUz8tebAtrHO/myllOAyeRWi11qniK8EcyDM15
03pXsniF5ESUR6hZxOIr17+5lqAVCmrmwGV2Y8XFye7vV3JeZxrZN28l8lIdlSNc
N0RvrsdoUTpRG60WkMj6wDmVsR5MzDQ/asKdKv814IwhEIx6wFIonOdeITg/FdEz
yTuIEnGJ+r9Picxj1z40IfrTU7jE1g7XH5W9qoUlG9V4IWPPsBZ5pWz3xpDY+Q8+
FidX/xML9cTlgHyBLtm2RtNU8wWCnL79Q95CpiZxoS1JrGHtNfEPZCbHyJv0/w1x
eBZ+tD58M9UvGuKwoG78fULVwtpq/MULiOxKZHCRGklM1v2Z4WSA+69x9W3EHCQG
sifiGI//gjH4aZ7d5UVUDfDvsNaYbul0eMJq2An2iX6NtCQwk8u7ZB3aXKYi2QIs
4BXrKyy/5BeHuu53hwNTJ2n6pwwp9G6WtELx03f+l2g778Q3ZpIUE3yXruS4gGgt
4yKtGGu/dhO5EAEcTokRl96LTxPoRjGR04LOl/N1wB3RnDE5r1Jw0PYEY0VKUMhW
1+GBVUqV7MhisRrHUOfR8A1Txg/LkLVDtqEGdA0oqsy5MV5SJC4qCKwTj8iv9+7w
UOx8gPx5FZJGyVzVazlSSqSzIMnbxZl/PEZU9W0Ldn7MhJ2ygc07fVM8uKFlPKx3
crZZKr7IGUT7IE6SKSqiSrVl6S5ylUPb+xiaSh4k4Bk2vzcIu4O12EBYvARL6Abd
MnlQ2tIZk/tKkBt1ovXwpjMdGtZxcce75dSVA+3YtAmNucSc3nb1l4lb48GagUex
B1y74CndrgPRUcytD3QdGYxJFVStrAd3e7jlawVraaLnmtUVA5dQg2SiClkGhGeK
qUSEiE0UDs/YM9xQ6t1VT3ebdnGu+GFLxVu8ng1Ji1GWFurvm4PVDzUzXDSt9F6e
B31dNF6jW7QbLPqlKOQqLwuw1C35tBAuDzAfkYzHNdfu8bH7q7DemMoR2nbvGTyH
IZN0L9f2XzoTaBJOnw/9tPt5Xfyd0PPb+BCQzY3I14gjCXiZOS4W+uObWEz6r+BY
SXTE7GK67bY71FF2ZTh0IZHqnPnoReUZeoSn+JMbpM6HcVUQ7NMY1hzYpLjhxZJU
HGvSnvF5KEEM3a9riaMt6hZp+tgUPbDd3Ox5FZHq1ZS1UhEOJrfJ3rRp3cvkTo2n
5X3npjXnhFLB+6TYzOIUj1ek9RCQJJwO5J89KjJAzJuQCGB9y7+2lFsQ6kqf0nEq
QaBzFae5d5WC9nTFc+MeopS8HXBC1/zwa+iX+Pni8Z3Y/yWQrGF1DJbbBelalTqc
JW1NyAxQ5EMBNyQHFDcriuFIGiIHo4Q8gMtGjWRtSUWxXHqisbU5LIQl0vBgSbpX
jg6P5M5CQoSEkeE/NyrhgUWK4YCffikJGXT5MTfQy/7uTQQ0VeFgsMX5yd9yqWPs
1h8E40iSCsaJZr9EQtRfJGVQrgetN19+NmKZngVB2iSUTlM1hl7eWfNzMrb4/I3E
Ok10Xwsk/68ohdHqjfRGVBc6JCbHZr2ixjce3Ekm/o6gBs+AQ9ZqWIt1jD7cqdVE
wjtAWdPH2Wo/+rM8c+EnEABFjTf7d7lvRrXK5n9bmzCt3aoOPqeQC7sjzwU6MKSX
qAs5rFD0H/TRFiCEY+FXVvzRWUX0DRCRSQB601TP9QaftpTvb73gPn6FVrwtZ5xx
vdWC9yyK5l/JxDz0ebsubHoEYh1VeY0uvvQo5vgLgP7u5KEK/D+ReAe1Ets9z4Ly
BcNc93A1WSW2pFMdVU+u0m4MB8EAN7PBDYqWRykH5YMMHQI8u2KSxlHuUwPqgBER
hE7SQ+YJXbvqVLBThb3EYQXdgwTA3aLSygL+Js34y5xX043778LZLsZ01KxYCwdR
5pT86yP5ib6JUVaMlrwpnUTnu1+cMs6TdALFqqLBrANOXQ07olBjIw58i6KQWPWb
UUtjhUe5F/w2GNZd92DODqtVNodr2sWSv0c6hTQQzqnRu3AMivGdl53z4uEBzhY3
/fYcmvkq0oLtv4FeMw+kmEp9+TJ0UMp+F80oCRiEMQQxfxB1r0McsnrdIFCQb6Re
oC0J4gVgqnRG8bOxq6Gu5ygabkj54Wo1Fe03q8UNcvwAS9vfOpH5iKMN01ZMyOdj
VElEn5eG1YoNvqhIyjJ84J3YMZgKHApQkT8ZHsa9fvguaRNZoUmB7yWxddJHyzF3
WapXtcwhXG1M/AVNXCCzqoAUkPOhu3cN9NRwjb11sciD38bKO6X/y6DDy/6Di6YG
KEAuBf5U4JYl/Dnp42xC2ynDdjWcZB6fNjade4NWVCa70NP4qWu7yip8BIkc5THM
ujClWx8QinR+OFV9vwGrlV1gjkNZrDs7zEEd3Mess3uORZK4FRwje/NFKMDuKVwL
0Ug9z8Tx94nyfi4qFdmO84+/q/Yeg8nyNOxCg8WhnGvnpc9my1Dw/4RZ59tInms6
XxULcEJOYrxg0snlDCBa3o/96mB5FfqNqBJyPoKyIjyS6P36Z/GxAwHbxoEe4rn6
AQpvCYUpIEy2VRQJgkOnOQiLpfpCZ3eA2HxU94wx07aqX6oL2MAqveGox2Qof9X/
zPJmWUGvjh9uL6Pub5x0yNOdcVeNR9Uhc/6GRGZQt9u1/tTtCTvtUldbb0Bhyo0k
PqaI2aO1UFPqb9ZHfv0Vicemm/MCx7k3ndheAzwGnPhhDpRvRCGrXJMkX6jwEGl2
Z0XiEl/Xh6MSt1jyLNv5TavfSxef0jpod8cWY2ljz5Mukn4uAxCY/MB6NjLhT6Ba
ciyVHO39YJvz10v0sk6ZbwLsxwLPrdkZTLca7+54FkhKylWgkbosw9HMtxBr0YyO
3IK53EpRqgLhzjJg9eg7X7fURLR31iAp7gCOu6HahS6PfAfNLKADT7/BgOITZ3su
A1a2PAfyH2ssUnmv8UrCT6aSHMYYF5sgkw11D0+w92tHT5GCpwyQ0wWdHDoPFS12
ZskUqXP13E/SsmgzHQrM8aDVd3Ow8dOnhqO7mGFqMBzuGzUJvTTyvqmgQjJVBOfl
QJ7G9Xy4ec6r499KfNHhQuSerSVLDyWja4iDRaGByrXE8ihsYj3djwQifSmCyEby
6Xi+mQJXvSJv4/w1xQZtOnGnuKpZd+qxLsuLqbWejEaauf8gfth8l0O9BWzjjBVJ
LPCDj6EYgnF+8GM5+KlbcKsxhPWJFZ+h9eSQ5w7oRcKmeO8RxmmK1ZDlIOYF7O7x
fw6lXpL/HJkrXHutB+gjjlYdknztqXlrC55h7ZP4b4RkYEF2Vm1V0Sp9RjmhVao2
jZamFNFrzX8KLUaEVfF6BZSaNjqaS0GDUC73XB3yrsYnzhbpAzEqA/yu9+pVjmIj
hbwkhaSm8Ei071kuJ2HWkLBTGxu85wcoNDDs/R1A6f8+T3wtxBKYTUqUouXWkaSv
JCfMkdEQWXZk5htdTBjd/lj8mHBYBqhNy9IVm80lIVSoE/MbZs1T9yzkAmB0svaQ
7hnHVDTQ+iWfPV7RjfN7z4uCKT6cliEatxm7zSOgw09qF4nlA21+rc3sJQk/0mew
YKw/yyR2MiyTVSzaVANw3Kmhu5C0ptbi3nKgVHPfrqrFfPT+VDUNilmg93wm0LNc
SV9SGbMrJDgALYQEGcPzn5iscksPGThk7otALiJR0I3tvUZdZHWoYENAxER3q5ti
8lQU491R1PwAFwSmYIq8NdM4QqrrxFQzH30cLYkBuvxIFL2AG1fkDy/ELEDToDsC
uiS8L6M2eSEzQ6T9ECT4a1JkjxMFS09wUtKdHu3Zssp13zywV5gzBf1jLROfDR2P
IhyatLWxLdYaDbqFFaD/kqbOFr4i8wr7NFJ2vLdJY2LoWGhZ8XpYx0Lul0BB+7BM
4EEOWbiN9Llwjr1JUGz0VpS5mTa5nPDlF4OCxwHGSaTQ9kstFBc6ad+vHJ04gi6L
6jqzDz2cJMvFZffz9EQ5enwvqF8oHMfN9M//xSzC2HOT0kDRhcAtrrSaGxpj27Ae
aujp0qmU2oIRwXOZvyyPpfBZl2w5gI+dydD8nB52EzfmMYKoe3tvZDUVhPhJvd+p
LKXnHPwUUAV0zpBFcx8UhqrURApBof2mtAY4oUJ/HpYOknv7yZrMujh3cZB3y4Lz
jTWpcg1jYFD+UjK1p5ks99baT5ZSltRZD4ZyNkhs2ibH8b4Et0qjPNyRWvNTAArX
dnvg+/ksDL34hEnMIVirzi0jV6m2L3WBrISsxKLk7kJdgCpiXrU9wohHOU7m3Z0e
qJW2Ibl44sXzAtdtA+kZ05Z7tMVyG+dQJjd520rgRx3HNePQX29KeLLWSmMmzoQq
7e32CH7W2otPslQVw+7MSLB4PKBVGIC7Z30QQZGm57Z4gWwJoYuhj25EAFD0/a+v
rVXr8K1SyeveH9VepDc3BVJz7tZjFUMaXJTC7Z+7XdLb1oCVqQqVtXiETpnEVHzj
5dFmssrr6+Af8nHv65XRWSENn0pob/wyEe66WuBLR+gmkCu3CTetuXdCV62hHGCl
13yMjNqKzljw4jLrlsTDzWhdFX+xsU1ZtvSsg7NptLPEThGcgNJxUfc52e4JAjga
2ld+8Bnqg0eaEU5BTmd1HfqyzuB0+xRcAmNN6+nLqlLN7ad/pobkf3+BRd4d1kQI
P/aI7hQ3+9j0BUVdztnY79R4VAu7J5ZZnKSkkbtTBpyP8nbijvst8R7W9Nzjgb/H
9xmwPwYWeSlc+Fmq0ygnNGzcDUJorsLxBPuNnqLR0cJmgRMe6ide0Ys7nUs4WFVZ
5D90XSxacMLe5H6OivfekL3wnibKI9E3HOVYFVcYjgABYnERzEEApzrtrxMnSr7A
YXSOTOF8PvKYYZ1eofRavjyLgWCGxdaLZ7V0YRWYexttu1tpsv1jJMEhpva18XL7
xNM83RiRTVZP8scbMHmSrC50P/+WXEZ+tbNmdRJiMUXr/tJ1ZhQU0rBe3EfrzX0L
JMm9sLvb+esD7lEEXtihySW0lO+hy0YCMw/XVbldAIltS9nUp3cMkpqiW2Vvj7UL
61gWN83nphSorOy8jcQrh+ccf9ScX/ZLAGmF+IpYji4kQeA2sBfQxkEog8j0qQAU
DHUqKDwW641KSc1zEzx2dVT9qXyrhwHCTEvRXy8gm+Y81YSNrMOPwxLUZs41a4Xi
fv1xqUunfLjn4f1bz04KCKgRyIbrz1IVgVklaT+7TjNywm9CBY1/uM+QeZQyjTkK
KueqGV/uEPAcz8MEX18IgIV/KjcU6IQvmHmr5mvboLfSFyP90GXkmtLiIgk+1rzz
DEEc1HvYVL4evzxmnTmxmbhi3LxpHkHIK/RhCMgpLgEFMXDT4Nj4r3U0+eTr45ug
iroD1ryX4ozFv+AAPEDrJ0aJo17bRB+FXAqDpHsnBuH+yDztxIBr5kfzKYAussei
wVJyCrqnQP2pgRhztSYArAvtpkVgLRouwA8E0y+mFdNrsDmO0Zd/Bdu++Dr0UAaS
I/fulbPcc2pMo3pRHXeZlMm2nOUHVR/UEd7JcbiIX16lvsSeKguLbywQKNCYx45O
7anIda8OHwNmCGKR/jfVlVm0aEZZS7+njvPll5Z0UzyiFzYmZB/or0/dnFhf71X7
BJoUT/319w21FAV/W+23Cyp40AMplpvn+oEM89c5KuW2pghGxqgV5sTHf/oGr7Na
rF9d3G4OVoNlA9NtsNKT1fi+u9WLIhcNXrhTaNEQtO9TZ8X5+lkeM8vmXXB8rhr0
qAoFp2uamymU75hyeCMoiuHXwlQspPb1xuLQFh9FcNrCqSdlri12dvZPWG9CD8lc
NlM80YVbe35+9e5kS/kvOduDKAy875+ebpUfurZXuUccXBmcPWouLLT5OwcUy+r0
B27wxs4TIA/oVjziG3DRfGPwPvKkkzRcCRPo6bmG7Cjcp5v8Z6ebyD2LZPzOcZO8
7enpLQYzgccUBR2CXA9Y3b7zOZgq/z3soxVildNZhqe0OU6oKmz4TTIYjsDwm+jK
6l0ef1KBhFBHXr46XJkcay+FEaBL9Yn9hTqQmrJU3ixXZb2EuyQG991ttVk399vj
Tv+eaM/QpCS0aBygHRWfZT1cH4UYUhP1QwG1WowB2tTcS6gdR7JoUbN7E4N5N4dE
N2Bqp4P/1qznfNxl6Jwm0vNO+lMRQzlaHHm70TzrmhV5KJMuY3PaIj37HSwYws1o
3R4jzDzDVfpdYatFLTXNEmIV9IqWCQWgARtmalfLyLFTi/aMH9HUJM2vVP/1Km5W
yVqL9DbB/ygj3MezhH15frTkuBRMlyzGxsiuCn2G0tuduLxL6PemEyw6JuAR0VF+
hwIHaXh4Eak7XtihaQj3mNmnO1Nq21QHb/9ZHcaOYFDMKQQVETgEyITb9p3HoUvM
jdBphsTA8nVnfD6rwdszAhnOlyC68QiQo44bAESSfNIpuBsOv813CcYo2Au6UV/a
uUSWcSBEByFaX/7MTI2rXmosQxHZrrsnn/noCEeSeIQDnc53xgsVjGyVUez9+TGn
E6LsO3el+XYN8VkWHu6xtA49cIyaIEVBT0MRYC0PvW7mFM3htU2ym+Dd9NOldJFK
RSg/3f7tMZS7aOg1cmkJ2l7XcAQrTkbfKxTNk7jtG550bE2NUfQIOAolcMH3ov16
70K9QTlN2BpqkBuAeqYH0KeyOLI/Y03fokcmYSNRPgb3AwDMm4FWI3umXqnUj2fV
QsS8VCwwH2igTk3ISWU8eFzKmivBh6CTGytu9kdQB+eU/jiDqSOeFT/Rii9zcHFT
BjkRFMkYhtkSU9ILlkUdlWPVn4to9oJi+6hryc6yOsLKWGO0xCpxmx2GMSpIrHop
vGUBDwCydTWgsvbjpi6YYKroZvFOfMoMgKY0mDQJiz2jOWiItU9hrllSSr3w3Hvo
9kotpaBx+RgfFsnKqcFC+6rM9/3RCapq6L3DSEKMTQdmzPC3Vzoz3iUgS8Jm6otv
R/uRv5OMOQTyZp5FDKCyKa7p46vzZRhRb9xQeBMf+rOPszXpZ47syawgBcwuolzz
Nz6KNIgTSQ8AVMtDNB5pL+M2LTv64G0WeUhXN7fMUoS0YTMvRyl/b1K9armEpm3m
CjTdeUT4GPaiymZqMUclI2MBsB4Rgv0hiwZaVjgC0Saxa+RPDlA+YvHPpx8SslRq
jfNm/YtkzYDy2P+UhxnwQExs9/qTAL0yvdnrBPFSpNvsU9k8Fs4uhrEOpuGX2go7
nnSJpiKfgYYXK7gcbzDYGv0p+mdSiFJnZbEtkjbw0LjuLtelxQAEK0IRlBHpP6rx
bFaGcQbPFHosktQb3uqyHioRoT5KdVt6oLBmDZ6AzB0LMgDIVVfHQUFVeIWZuqfk
CagaQqqpZ6r49pT3TBulkktfeVQynDaJGtMRCwkD515wM4vIWIrf9Z3uVM6sVINm
aC/WGXue13ms/r2YbnhnmVUBjtHoE6gjTg7jDqwjWvqR7BuT0ZKZBMsnFCziR4Jm
M2bcZ5Wtxb5v9gOgsJ4uuRxTZTd5Z11Ps9iwGMDfjhyw7X1XPo4DTBEYhE8Ur5Xd
hy5nOhAGTj8UNEQeFu8O41Ytcf4I3ddPgITPrsUU/0VO47mbgN0l6R2971xiFoF8
1zM0Vifswc99Gub8M6JyYIjhU/muaUugZ00HRwIcr5xLhJ8AZ67AcsKTPYj9RLNE
EmKBmb4ISPoU/fvrc19ar7aNhkYL0T5BieBTn84iccDbTP8n1rQxxEYE7pF21Cpt
XCQni5vMzTGtoEppEhbDMmCc97yumKkmPipBRcXcnWdFUPyGDuFlpf2FQ8TNydp4
1CJz44gYtFwbmZd47QZ2ONV8qQBtDh+QXUclQloIYY8SCy3fNyUvdpUNj9gAoM4q
UPxcNoL0Jphehw6DEYIEL7z52uDGT0wbfrfpEs80EtVUOIfEVVLIU42oJOm9Q1r1
vVi/nZDUvM6Sx9kyDDXQnJU9sWgPX8FLj0vhXpHphSpYML8Pu6vZRubIpCSGg3mV
dXWSt6tpbVX/asOg9ypBjdTHwCZ+kpS2UKvj2zLVEPBvI8lbULi1mDFTQQcGCkJ6
7ovOwuYwVM7RBnUvoQ7OazibB1aAs1HzxLYNI1TKHMQgzE+vFNzmBNWjDSuJE0KI
Fpp+Kdm/yGsn4Q0kl8mKdtQXpnjHH9H0/f560TyMAOX3hcFOry9dwn2dPEnnxqMR
5F6X+tDNYosn7YVRyS69flrXhmjUSHm/qH1QSF30xlhb/+RrbsqvMK8jVY2NKiqH
vyDpPyTLpkEUKtj9/UizN3zV8xh6QQL9pWgrWKD7RfYfc+IvLx2CU8hcrHirHZji
xKZ9aXfxh7CwYah9oF8F0I6VUVwsu/0tttnhHpr/9CjF8rRPa5L5i0uUTNQSEXYg
DUgqhbx3dcVPrnIqD9z0i3VQ89QPubhrnaBSH0PQGxgbAZ2P64WCs24pBX5YenBl
YhoUuMTUqbNIPeghGBGLoLo+dmW45cZ9iCUvpBpc33KjSS0dR687qh3KPQ3J/n51
9KTR4w+ri3ZVEHssJCKgC+OkVP6QpzlI8dixjYW3IE1dyVIodxtN8R46vKkkhqB/
oS8TDrpBpU1vcW+EwFXDn1wKAqipKITJql32FL6eSf03j+CsP066gL5bwzN8sv9W
dVpnSZbVqUVKkZMfet6cZOYfp7b7aKcZ7He+JnQBjm9lylvSwqlB+X/JQKfqO8ae
/BcCMuEm20/Nuc6WDKKB+v8Xn6UnZoKVXiAQ3yz+YFLlKoJA02PdPf7wPWxyWdKI
vgUMtvsjZhbLSGqkL+E3/GYngEXjxPNiD09DtAjk+uwNM7h3/Lh1eAxODjLWoJ5r
HVw5OQ1kLm9zbEgwDaOdA4XeUK0R9NcpAKeq7gQfIWljcvbx2N6LWv+gQtwRUFUb
CGWKvBCdPL6n489A71nzF07cYFTLU4y56cXyhMYkhLid1dq0QSpl87BEvR9+n/Rv
tUEdd3V5x0xv/nHhL/SifRCF0wQTokkxiOVbqNbwlVeBDyHcXkP2wP2xCiW0wPvd
a+GMRdyxQXbKUW3tb1pJD/vUoZY0AP2ro7ghbHcAUTuf3kF+4p1e0gCCRAiwtKsl
fw9fyoRPYOcm4Ad8ZNYJKjWoDoJycAMyatzSU4MidcM9+mDqiBVNybKL3ZUIahqv
GvFQ/BHXZc1Mab44AltCwUx5JXcsU/sjVb1t6ZRb+f0WLLDVlvjHWZqjxVyOfqN2
XS7wIUML6mMhTD1s1RiqwQYscXKlAMEhh5yMcMv3AXJzvT03LwRCastI32rvEzUu
ZCwWxuSiXAHgCnEHAxPT1K8nlWKsFOTxY3XwKdtWjc6hOaRqiPkKIA7WZ3UOecSo
MZ6Y+W0xQ80jYe0XhX0jj63fpyRqcTPrRnaHL+37bUOVJjJOG0o7m3gLRiUfiyDZ
ms55TlPKDhPyLwNYbCDrLDtoIJUa8aYO0Jmv/cb52zaaGf7412LqNclnaim2Y2r3
wWYBwMlP4pmUwu3SeJnT9Ei3PKM2BcyumpH3ZZZh2G4ZGzTy7PBrkn2wU1nQkKiH
SMxnfwIgFd6mchySDFXFRJunlqKGd79UHXVJbsBMGQrCCv5t1AWWcMQnmuJpjVPy
9QC8WsCrKuhmptY06/ndu0RhmY+RQhBa3ZeTn/XTLFLifo62nnpmxG2dfMgAjkbE
kljxc5UBXWyFCDKXFfqvlrbR77CAzo41ae6J1OLnvKVKK9vyR6ATKM9IYnIbghrO
rLMAVGTYMUGOLK8avtyTAQ5jDqdVlFmAjrTOBH473XaUhflugriYdx2d6P+pLT6f
1jFUCRGtvxJMfV3Z3hBKMurs3hqANpbRuMNJgu26sSmZtm8Hi42uopQcI8aEtUUB
U3CfhDaGs0iAUe5v05pUP8i7nK0f1U0BmEpsC1AxGbq/MzU3JIQb7I6ZOnBr3k8P
TBhWSkHZPI3H2HlTnle6fuqmecmIJ7ArSU74dl5EcKjyaGy26KDr3Bah/HEkdDBP
lD0UkbJFlUVzdv0x2PSCguCCv0B+4Tl+BDGE3f+T5PcT0dio0+KGas1DD9ooC9Tp
WbDRGiqm3snXQG17xpzKXq5dhypL0xCeTfRJl4z9KkdbCEdMLTw0Mi0sFvhQFygR
6pVZe6J1qW4jdOoRYowz7bUr80Z03ucYNQuE/nmT6Vo1MaKWqoR7tC+1+AWNV4Hi
i0hHQs9GCg35GZ+HzYlpIGgjCsA0jCXQc1xebFZ7WGifiLQxTACjOcF+W4HOISrD
xVXymXqQWNf8AKzrifpkDolV1UL1u4AfSJ3CibtEV3sJ88mgim6Rkx8MR+60lKC9
tv6FqCKqCEpo7tcLuVo4f4rgMAnHzFmPXyV6QZWjMYZiTOVW7cWI2wbrHJ3bXiDV
m1tKafSanjELClxUFtNCg4rl1egui4cC/uw0fCw335V67MAXMXbmoGsFmakmrKyM
Emn/yoSsYXrYGBobDfRrA79APV/dUxFd6iAntJsdP8oHNfB81z+L3GyDOMsrMAze
D017j+wzkstK3FPXuArI54qqV+1iMUnZyw2w+A3mEgWt+xrSjXBZcboySVgnVNMz
A4Y13Ae/7Y9/7Nd5zFSuM7zei+fsNasgixrM8SoXdYXgp1nupoKATbg9z/C/rP1i
NbBGxhrUScVIrRRIeNdZbaoU2oHudDNTvVRhD7cc/okpZKHK4Xs2s4LFqKtDLYiT
xhP4YIYNwFEdBWdIywJRynMKNO02FrCphlbeNDVqNcm5pNOvRD7hRMsSI/WiDTwI
a2rMFtSN+PLt9TSflci+jFvKPaWG+BMl7Ae8WJpC7qpNSeCzuaQJTkQ5ISocdiiJ
ro6TC+ruLKGzvc7Ks4lJMh0L/wWOj9XZAmx0fkGhQagBKK789fWDuwx3fFCEt8hd
N63VWZCRW4B4iQcWrg1pWkp8wAwLNJ8s5ikX3o9cehTPmz+w7NoaXnSTJtKjWAQI
muY1liTlIjUYFeGE0nnrVeTZqDBTpXDLeC8rzhRj6Dbf7YV1aBJg+panmnTwMxlW
5yCHFOdTVXpdtKVhFx3J2wD3zLnsv5wEGJtchvR74tW6m6PDqBLwws9Lmt+f8P/y
668O+1qUWPTa9x/HwQE37pQaWMYUnlo5LDDOJhOrjyBfekf+1nmjiC8bA3c1WEAS
KPgx3hBB7DVOaEaouy4kviaqEY1f2+RrvJ+4R+4Up5B9izYHUh4iDmRCaNELqixm
HSKAQXUOdJAqCKKcXB+DYX9mygDPpbhncO+2UPDGfOPFZwDFbzSF8OCREcY+G3xN
oQxNbIH3m3Qp/ScF7MpP+d/ujKlOO6M0/GkX0cgp3TElY+ug37JIZlAKhPK6WViu
mpZLtfEgEevxxfSBs8dIZeZwX5fCuLyYEGAe2pZl4d2sU/jttxYHw2tgn2wcuF9w
oRBe29iXLzKmGTE+pQvDc3pmARV0o2XBtVS7AcMznYK+5r0m3q9ZH1AGFg6k2UUQ
zk9jYVOTTH5i6vUATiLJgPvgysr+5eNNABxHY5YoFIb649G8k4bqtOcx/Lobsd0p
XwdRWFugZ5eTvkreN6mLPrWY6vUmFA4cddRXe7VVlpqVaRzuWS4sjrhRAHHTFU8i
0+f1yubK2La2nlwLqV5NAYlKFOCEMV2Mo+trMQ1MV25zKX29nvPtGjRZdbMZpBwG
1pDGSp+bJseR0UvvI/qA/bWFjbWp4sxfASrWYUh9UUK/VI+e4WZ2izJCOi9xAGxg
btOT/oWwTh7fohOts/4g8i4v7l8hAV6VdDMv/equom7vDOrKz4PtldlhX5eNrgGz
8jXqrUPeGrjSzwZ92Pk0OHl46TgIHaP0fcNfpjxeLTzga7Hcka2PF4QaI/eBlYtE
PWw7LcHrfMZA/0L/0+gZrZ7QFvJBj1ojnUHDHRKBaN+GMlgzKp/T9YzA4t2WVRbb
Fx52cznAD9OfshDyulzkebsY30erXiYVYYbQ9NkmKbM0Zl7f1Km1TGVg8o/PuLGu
BpZhPZ3vdRzmRX5F9BjTrzy7KMm4YGo8PQVcU2E5U50Gz5BTdEGpFKMUERWXbEMz
JqjkFvwM7OMqhf2n2JNLKj+P7MCS46UkYi5DFopC37D8JMTsr2YTcoNFm2N3XWcZ
DdPeRohBhIzR64ceUvMvOv89BuZrPX7otasb78RwPLob7fau6AdwALGZ4iAZFk/f
yO72l9rGKc+VSU47sr1xrSQgUIpt2MBaQtxLbbQXiyywMZ3lm3OSKSgjkXTCaywR
P3AIMt/JlwzyxPoWYD1z4B5vO9AWrPAMPGQJZ1UFemSFr+HJ7zJqxoxNTnRGesOO
72zznPk/sx7V0ldB7MnJYIaxf2x84Nl+bLHggvKduEwT7YLbvWZT02FpMj4hKGGx
XRNViYLvtP/sGXfSaAWAbzqYxo2KtDv4xf6Ts4FgONZFOvgTXbjvA9ykm/0K8DnT
ghRwrYGdO25M2iwa4gIVoJa0/DUNZttZNz0VB5nsbzqExBeu67vtVmumiXg17Xpg
n1vBc+CYaH+ToXr44mwNwlSqcGtV5qOnaJvptFzjH/+2hrabVdWnxHkb1hzmVE33
g1Otordt9NN9nQUr+gqpCBaXtGMesis9ETMbQgXgsc4aCnFuYH8CdXfSSzW8WluE
txt5702q1Tuk/Il8gy0z6PrBFk5+r9d8c4fb6xwGzTGfPUfne41kJ8mg5emU8Vyv
iWCKNw+NfBOT2L8tCPxF3LALn/jJdnYBVLokFo9766FNYgYO95h5BWmNoloyb7tC
QarScnmWv7hEW260526HVdtZVELIqudDySqJLLXKlQRwGsegttbspOk0Ai9aRGgL
3wXI0yUTMGCpgAH9jo3mzUjLq+lk/OGrpjUHgA8Oc1mvBNIoIZAgF6cRZmhBuos4
82/3COwBkHWTjmSR9UdudU18Rp/KQMkPa0rDCJcxw29fTncSN/yoa7+0skJp4FEy
9QyUWRXNCAMhY/D42AwexnyQ3f4w1mbVqbFYIsJS+dqvgN8jObDKY3VvWL07M3o+
gT1X2DHEImmdSHMBIl4DBS4WuSD87dPthri5Qi/V7f0y4owQL2l4PBPW57nKh3kJ
5wRZ3DK9f7JWVUPHxnKib1mq7AY1uR/MQLqZW3W/vkXt+XhnCGyCLlMhcc12cBqm
6XFpRPYlSJCXEhJoSJx54DkSF3NLO4Ly+pghdPaOocBE+Az8dnGZfIWZ6wnu7Rs5
BoERczeyW3KEkukNyQjfUifT/BR7BSx7S2/uV50jz1Tk02KxHX2fgoAnRNFo9GLY
l24x2Yr8nMKTffeZ/Aqs1u5/UXi/8H9pI9kTCMSJ9xzThW1ajlGdEAYg1+txqox0
oJghTB+DFRn1XEIR58vexzOZO9rXWBK9YwuHoy9/7VLRQUpbsWR7HtdwuawOcCYE
UuGAqdf5IQTwKXp1HqdDs0mSxf0/wo4ACTRtzt0MO49v6OJKoVsjFp4NEcNgNLA1
AMF76blLqPjlredvJbgUr7likx8YRX+9OTOXjlfacEtBihH6k5Xq/SQYbuHOWFa8
POILRyNAtynfr7Dz8E8wa1e3ER3WS15/+Q6ywEAcrkjXIdTDvFI/epKzD+7o0RCr
gE+lfwuijlkqhhX88GsB7AB03/SGfddn3lfkQOQE9aRSj8B6+QXe1YGwUEFLlAsi
IcW1Qo5pb5oavbc4EQWYSaWKseal+cYtnTzACaa5w+wfnMvrC/h/5yCxIunp3MaW
F8XmofLX4+FXtlk0bpE/hefN5J11wKYR2JBqx8Il2bQrfTkgN+wgTfpkAGm5pu0m
O8uxLX6LHsg2xNN/GOP8CzRz93eQVRxicsvua7kTUvKCIcdC5EpjzyYfjDBWloWg
T1I4Xx+mwfOtSLDGYIVENNS/4Tjw3PZCl5d0Jih7w/TWHoPw+wvn6jZtfku6htjC
I0VCzI0EBHxQX0u07HYLi6VPT/H39XZAFaqd0RiGZlCbYYLPofGzf4Vj4xO1imdj
8hkqvKn16U9Hd0S5E2mQ8QD4v4xLwOBsfFx2nqMIXpogNF8AzQmxEd2xrqDrPF/n
u3EPJWDMyB64Ekvlc0LtNYj7mZkFq2OGLbn40/vUm6OyRNqZBP2pYYo8x3XkRHoM
0IhFuxVc9K8mm79Ul2qBg4CJCTyvW/AMIsacSi+7oBJHITdNwZnAbwBkTkzEF4YX
hYbD0O7+5XGyqJOZAl0ISmYQGv1ZcXvQF03XmSCQmKcwk3yD2tJcQ7WVJodXYtdH
rpj344hmVpkopqlCtHiv44/2OlVqpjIxkkGgvjH4gvo5zMDi0AHHaDgDjfKpedkg
CwyURiTBZqFkmBHD6FSQ5ZCm0YkwwCQy8ZN1fb3eJqKcMTysgp+V/TjbBeU67FzN
MCgBa74x0mZUUU9PJzTvvFTn+nRXF15+uGrls8NHcRac8tX7at6wEs8IviwrCLSz
GCaPvZJ8MnSOYeCB5ycvaxK1y70uKlHGSQMXpuBkCns1IPf6iYGOCE52LMohAtWD
k98SdHSSaLiXvzYNndFXNIo9TDCxA7PTkFjlEQQVpk92ZfhwKFF3Lzsbp5/a9KZ4
/kVtU/fjanbHHD9WArVGzVLUgBicp8TayuQSIDWcZHILOpz4JVMV5ycMZlrNZJ0k
EzJaHPokXiDqaCPPzspuNEBwoxIz2xCz4jcHALH2zdTs/LReWLiG3yzpytfX5aRk
5a3alBn82vso9mGKm1UeKDpkgFwjghqxhESDIlCnKIpRpZ40My/8YYx3DeRNNxc5
I0PyVrNW3mqIiuZwfUsx54hIQh+0igdPXs43wXDrNtK7AMtU/vgiPWaz5gls9SEJ
oixL6r1SkEBUXwwIbBqwNl+vClWR1Sfqes8T7Tn5z4CoGqq0mwlvF/P9xukEkmHL
TD+wbzU8CJD/AHgiXXr3/gKMq7pTyEadbTH9ES/GqBPfCRgjr6LANg7BHmvBBGNu
dd9FG08sEg9wU6omlFJqSvYvLlh3VaWmpV8W6+xU71gfW36bZfkp42Dq7sLbvLEC
fA4X1mPxXbJPZSj6lAvcKsBnL7sRjBIftjcMOe3zcwUyc0HFno6b6gi2J6dCYkU9
UwyYM9JzmjBmD9IqCyeRLDpCsVo8xNdfEz+7pMx0V9XIDol0NlPaP1/jTtCrlh4P
gPIe1JVQTvOIl2kxoh2j6HCmGkFbHhBxwoVS9B1eOEwc6tXnb37weT8G9C6dKZsx
bwuQM2Uf84Lo7ZlhPYdAjqmzLXVAGi++lyGjkJ+zkZYRkPWjgJf6t1O+CEdpSfRh
PvmmlHghgYpvVdzZfB6x5K+f6tVD2CRJwbglOqugP7kp7jn9CmtvL+Nqjdv3YfoI
apSEBdxIsBfIiy2wNPftCHnkMdTvNUPD5P0zWCdc2Q3VZLTj8E46JE2j/YNWVNUv
jHhCx80R0WOg7N+jPF1ssDhbDyS2VVbkTJwY3ed89B/cg9L+6SwKVIJs5oRHkqm4
VMwnkXNPV6tLfw7Y+7DBDBRh8akInjEiPZvaasTfY4q65c/CknmBvUyyDB4GbSJN
kjLcTHosUf4KzQvUmALdO3D/aMIFFQtZUmeXpseVWLsQI00ouwpnfpg7d+LU0uV8
5N0TJjkftLrLrnWEIv+4qxbSMZlMkEn69jrN/uI/7pOmf7jh2U8Crk/0g2QLvLWm
sQH5T5ciS9XN3LQjUcLJ5sXoJzUcDi5HmZeu0tZnKcjlNXQDp7ZwPpdoEQZJeSIR
7O5Bc0gd3Ufhzf0Z3S71e7udQLBRpmuhQgeXuXN6oBD8Fgd/jxM7dDvoz/4weqOL
nen56Fj6vcmk5RF6P3aH+v5XJ2Nev43hp+5/a+iWV6fx0SJtZYk0Z3kK+opTwscC
o+frSZDwIh488rh9nxXR/3mR9dEyh40na4uMPdfTSZ5fs0XQxlj7N5TiQuDpY7jY
EoWqwVIQuXz02+bpWVFSdsDbI7ik9VHBtPr71a/KL1i8RSI+z7lZ+khh9rFgptJ0
K6oMhbAv1CazZZPEmRr7OU262idjb8GDX/AQX8q70cAMT/vQX1Ja0zocrQNZ+TIK
2+qrSVePowA2Xlf2kczq7s/7x8tp6/kDGvGulgm3POSLFKxsWdg+N+MmyuitZTAU
9ETAY2vVPulyVb6rS+uN3l9+0wrNTCbDVPgwwqpvtv/5qh0JAQ91IywoM6D7DUrB
UQdvIt/aKJ0eybwXeCmKuItch5Yz38+8uIkvBu5Lu5BI6YVycrvbbY29C/AsCEvI
b5HRBbkV612dZe03Col+p/mDH+D+q1zPpFWFRDIzd55Q2b+Oq/56GK/SlFtSypEC
e7Gb2+1C0kZTY9CEXWsN5LevOBlGyfu+V2p/SXX7x+TBuGix4lRIaDR1pC4R9qVF
uVhtc3hJxNRp+nk8KRppxgxgpmr9oSDFiThfr+QrcSf53GXAYGmRaCOE15oEcTeI
HuoVL1zw+Cyj4ABrjoUGe1BXVRMdPZg+A9Rox26EkxXWk2j89m11yLCAL3vZOTEz
yW+OaQ7NHSXG310hA8LVZlo2Rqf22rOrHQOnRP6ZVTzd7QHIBEWKsa8Zfd1iXzj6
T4dt7vs6vGpppd9YOAfrvBsgHt5UkVuwm8wc2EN66+9AzwKjWlo/tDsQSdGd4soU
YsCdnsaDc1byjFukuoAV2DvBnT/HhsM2AucoZbne2cLHZFjq0NT9dZPOLQGL16e4
97DgHHNzEcM930n8IM7JG7ftIUmAZBbPIRJHrQgWXMqnr3w+CJF9gUC84GWpNX8S
pjOq5WV2KrEzAmk/jE/MnAqlkKrNGnzPmx3+SaExq9kErQ5WFoIkPJgPhLu7w1Og
UREOc1FR4+gOi/DXOclTL2TuVeT6gYYrKg5DuBx2sOkX4oSpXGATfXaAO5/KfDga
YK1cQoyklZ+gcuSf1v+PIriLjYoB9iGmJzb2q8ZRM0XXz7JD7t/zNtg08uuWnWHV
SpJfLr/8uZoL7U+gp9cqUQaUMw3slahqEZWq+pufrm/RrAaKz0P4/71BkuiT1LzV
Xu7x8moJBaubXzdOOGAiUiniS4LaRPMiIbjrSrR+MIOdxuvnMptm/hx3AukL1Mgw
iXmLPAkTXV+dHq8cKY0TmFhNtgNBb0EM2VYkF8gGaS8sdJZb3NEF8tiyWrgp5ZJt
MrqMBqR8TPb6TluHf97m9q6DMD6gvQoqbfdK9sF/6DoLSDoV7bXJOCKXM1+nheTz
f0ib2Lt1KI771kdO5cyxQzHvvUqxm58DXZ8lU516A2FMw+LT2Jj0OAF+PSlhOLpp
DLH2Vozg9Aszv87vu5RVUAeK8tAdrjA8RN4Uznukx5OXS0nWsaWTrdOgqakIXf3n
D46C+FsXU6AK8eim7UXjCL89c6Z4XzfkE+3c8fxZns+NyNFPOxXbcnjUet3EAH/t
QJ53zcrpQxDgqPuBsTm710mJMXpP7BENJrR6kG8ScG7lyLYkmkhH+IAsLjVXE4uU
kuEPNuD4ZJzY0XQrEXO0jK5lT5g4DI0jRUsjSUNwmCUKxHLCS8GcbZEtC8g7WUET
9uWODE1b9WARMQ95jMaHHMvwfzYUOoyour+3BdQL88ELLGTXRC2Qe67NBu6sxo1v
9ax2Gu6imSS63gfAkayjElZ2yzu0M8yE9mziABeevUgskoATgl7sB3gMz9iMJqyi
hITd3W+MCbFIeBeYcFXstJktgLfPVwSET5THq+WIT/o0Z8gCDMUfkQllbEOGIsma
cZwRfkBHIgYJ1dw9Z1Pqakm4064qwBIToBFzI+hGMkcXmVJ9FrNpwXATqUTjJLD0
Uw75NNZBJ5+Wq2Q2d3EP8hq1QR2O58PlTgAyJEtWpQGm0KaMP/BCak8s5prIfDIx
f9kwhmjg1XcrxP24SHbZjXYZxXRnczrtBMOZrqa6mKYJKexNL3T82izuzUmFh0Kp
HUunOvuh0r5pFn1gHn/znRquhb/546Wty50F6UA/tvRjQy7ErhKXqsohyWWs1KFv
98AcF6cZSN27VUnbWbpc3Y2S9uBUW/CvmLbf99Ch8FdwiN6qqFeBFfeyhXw/buZ5
GGl/yB7YdwtKE9GpfiKERQzBFv2TG9WuNjTaMhRRbwPrmhoRbXPGI8+tYexeDBxO
w0Lig1/5m+b3+kgwzibOzgnW0nOJ8zaDa/Jz0zCSfpgLU8pqHAXHRrijzxKIypB9
0KcVSnfthhrSQzL4vc1HgliKh6nnz5z6mQO4zZ+g2UguYxjyBqDK9iJ/vdfe3xh3
go5IvXevjcxUVxR7ZmUjH8AKw50u9S5goBATSFNzDe8A3L8uYCUUxW4dRCC0C9VP
yTs9M4Ji7LFrnIC+7GeLn2DvpAo2OmJ6XgI+JnILT9yH4zUy1l9l4fCcuin3Tgc5
xELcRTh97PHCjch8E5ePeW1sC8Fg9nBww/DOQxYZJO9JlDVlGFn94WjksS6+NOMx
qouaccmXoQwu7PHUmRPDFfC38TSsfo5qPDS8Xp2oqvvowIh70PBpjP1e4MGG9dbQ
J9FTji2EWilybJckKbWDPD9lIAbEmPCCXBKff5ji+n613gy0uspFFzDdUZD7D7aF
fCobLfQO5pjgv7Msc08A2vGvfKMFjqGFwwkijw6qPkPzKTdd6Kai5Sgda7oNE/vM
wPEyWDphULRHX8Y+YFKdkqLIc5oRKQ/BWbjiySpbqpBj54iXyZEwoB1WLb46h7wW
pQ9p5p6xz0N0nCSgLyyIC4j6CSrqxtSBKGrq332g8wYMTvREb9IuwpSK33AZidbz
UG+y59dbfK/zl5/QfUnJQMLvxodib6LUHrXQF/okHYK7xc7ZI+VpH57zvLQRQyWT
lyGlITniz+CiCDcO8tiy4wQdn+2iVQiAut77m5wM8s5cpyFkSSFvHqHsE1VejUkt
OHNB44iUe0GgZKA8CMTOOi6ZHm284Qy6Z7qZujIG6fzdCM8DV9BgnLSB1gbij90u
fV5etneZRWn0kw4XxpZ1LaaI4aXIHMu37XOvm28vjXyzFAN8M3Nur4tjfTogM1in
fJJBegqPaANfWnNbZoh/esqffxYgdum4rT5hO7kEl4nA0r5Kdb2p+mZHqNEOIdpX
jUmTFLxl2Gaauy/HSZOnxfT1bkKL2whHQwQTmYvUwnhLgZzLt4yLJ8zTHvUBOe9A
KHTpBRqQ/CDLbSmsB4p/DMy2eRzmKv7O4p2sw9UPWVRSxRSTgI9yFCbuaqyGqN1D
5GX9RXRL/0OgMoBiBjIOW8RaxxtBpvT4v3zL5bbdYhkD4gkvzYG9znrUeRu+j/R4
A7DnUmUrH7af2kDYfuDWaz1F4MgzfOQJ7hsYJyAm42DkwZ5d/6l3UDw2VD0Kx5jS
lkfB9SJT/snp4JJe11mJl2S2NXu5dheueDH16H64+MD79WvrubB8nfEah0FvlDVw
SMAbO7ZlK69cOy4T6Hf5B8Z2s7KxuzmSseKN+UzUlXVcl7JkYUeNfCKXr0fACZhd
7OZp1FrQkofqO0uYsMjwd8wBksq0XYU9lYr10IO6Zdbdw/XgpwCZZM24CKI24z9I
kfNeIWl+tC4L82tvCzPh09DwvzywhdxY7U5QOyFPUsGEsKR/vZrzCz+9JBLTbM75
a+b0EXZJo33pTUIDLLqw2/ackmP0Hrb3ArSKW+bPn0vaGMpIN8aqvgB2bluCuAHl
KV9V+AcsYj1UHrwf6NEaY/TZMFqKLpfnwmiSKPmh5MV/XuGSgvGdza/NreYetNBL
oaYGzNZ+P45//R0DmX0e2yQF7OKM2RBie4AtNH1VPfaqr6EYqMwbzRszCyRZ2I03
WC6bse85ugNH8LTMpcc86a2YNVmC4WKRD1rktbkK8wCh3k8DZ/3Kub/J3uf9OGjs
KP98us2xGMRXZrGu6q/BgZWWtIZ1YWhzFk4j9zwUAmoDPazSA6cVVs51X3LVtbAs
YWPSiV4jFKI3/WLN5Smjgkg4CQHrD6MWSqNc+7G/eRFAUV5yhp9P+5k76f5PNvS+
L6+vlTmk8N6inW30r12z2D2w4AxWlud0weVW4MVS2QghH6HfodDT9h5BUfi70r6N
sQZ9PFXbuQ6E0/Fl2oCVRHEtsICV6GfgIuWBBdAhnnR96/xGaTDW3Ii0xhbm9uvz
v+BLR9cvPdQhR1PPhKoBP4jJIAPucyXCdAbHA9masmCffH6LD9ZFBuLcXNxOA0bH
5RSdkTbDpUe7aJxxD0vYhnExTISiPqJHV2JY88e1u5AlOfMbBB9akpBsvynOcDGX
hk7PFn2hicXNyo3GALL7Fl59AgzMUQiv3W9/AwCAcWJ02IwMo3IGfzKWbIquhlWP
PMtGRvxvpoL1HmTP/WyNn3nVo/t5BIeqRH9zghtbm3KsRXg8Iu76Gu7e849CLcVV
yA/LHGx++zdb0dxXX6FQHQpVG8o1jcuuuBCnlc/iX3zViw8DJq4o7WROpxVazdGP
lzM9+xS4t10zpEHrBXUKjvZiYkxCttHKoPshWfXf02e+5pl9280/Z2Oup1kWxWAH
LU2Xqy9AVG3qFSbI3AhqB7mQV7xjVS7qGoiFHfU6ffZX8ZwXCAX9O4oAxsRemJlU
MK1xuSf4P5EmiKxyyWlfNJ3rMemqN24l3WavFMbSt/ESyJtfrggv24YcQhjQOkB6
Cct0Cp0gqk9YsWPtJDNA5TKPM7hm61OCqB/RHTEf/liFJjGzpTdzeLR0d/U6Lq9H
uvA4rPBhCkY3urkt/DqubL10ihb8jBJR3ZZpsDfPDgevRV7ApUaYqiAzROjBTGV0
Vvlgnhb6NHDnrnutjeeYXwh7vcItwdgrmSe3IMFsZPxh+Vt6zRkBi3Vb+sz+WvDR
siosSAg9yqZJwHGz8KjhPVySYdphnoEV/3xo/ElwVkFH9j34UMqCFBeCbJjNUJDx
v4j9Hm8NJTn83iMq7vXxJnq6vTijJXMq42a89yU7rUObjLs6YPI3lw1Bls5m/HD2
Do6INtL0NizCzPewqqR7Xx/yLN6TnzGtLI5slgrQq7JzRc4VooxO0Bp6ZjGggs/A
pgqAQghuZwF7dZwVo1brj5EiqMaiIUgEBsEmMbWhVMSVtz5F5L17QbXl+YkQsR1m
3XIjRZeBMfzvQKlvtXYN+hRs+4djpYmKShtdiLynGWvqlgx8XcTAgJG6W9ejTyiu
HNBVOsDaj02JY7kzTCIZFtHMjRxM2qow1Iwl+wJBRqnIGm2DPv+zsDSgR8YpqWxZ
drRVoAkchjPUSJBBpLZMnkjS1IcN6SANKRlNokO6ampMd/6yLuWoghhWRy34aUe3
CApmNngDnkxfJVY5gEg2HtSntV4114KMZa9DjB0amaQtAL903xXCepxX1D9WfI4Z
0hLTq6ZAIaWAG95ucFg1gezRnv4136wuMQodrMEKQ5rHLh1zM1JqWWK1XbVH9iOM
wxj9hYXVh/tL6DySq+9nZSftJq/o/ix9Ay1gnju1+7m+tHgO3UMc08ffJeKHuL3D
Sba5dtacaNMSoBgitZcShx/tTNyOWa29zES1CkdJQrVVcWfPSDswZm9tz5kuacMd
cWaLbNdnrEnZFXgpuA8MQAqwpqb6qpCFys7vtv/8TtZ8TdS6JxJhci2eXKe1Bbao
Egfsjnxr7AQGRIORaktYNzSL1G9Vqbsg8hy78SgElwvR1gjRKlPoyhAemmrSDczO
HwyQb+nUIjrHkvlOLj31RtDQHrfatyUmgTfwMRlIAT64WOsaYIJQ29i++EY0FT0L
Xlv2feIi2NypScRUZx7OjDOoBEIjY/GdRedG5f3hteL+OpZThHC7eH4BbQZ6DrKs
bJfcw9MGLKj8BcQf8jvTc9+PlKikDrHcP4vAP2/XLYKMwIBcf2MZ2FYhF48JY8F6
PqgbiQveXxLCnAqUR12HpmaXwjXqETVLBd26uW3gpVl/RaaKml7wT4dI/2DQmKHG
xfIbWqhXGWdqVEyG9MqHLWPFRzJljuqlcW4Ej7f5jWfwxFeO+GTFEy2pk9Cck4ua
CVfIJGNm8hXTqfeC9n+7+cWh/kaojpsGLCsv+z8PpZGHOsA3wfjIIEjVGEZ3/QDS
nPCFV3Ay7hgnvmznxFa/uB8EbcPYvYu7vF5P3zwjcKZGvbpA8jQ+hmC+nrs7vnAc
3ZqMsf8sKtYussv1EjaC4UBFZZNJXkVAKjzI7oVDMN6X9BYixuyw9kJZmrlCfeJa
QVudHTh+e7hio7cmfVwu9aX7s63bvSOm2roUw42pYGSyzViFviEZGJmk47Yr+fGM
YncFXstvKeYMGt4+9nwzk024ys/QUUDR+5bZE18z3LG8p/HVHLjPZiUQfa79aXG2
eneM7J9jUautcbPS8nsz70JW2nWYEidDhF05Y7pvc7bYD9vLR3uk/m+19lOJAiW1
56mP0Kj7NR188i4G4rkP+mq0WWj0FI82qgO8jsEUKj7dmM6vbQ9fpa1ZF9v5EOuT
P/Q5rfSulSTlslUg+LfbzB3+9gQo4O+JANBPHMYuXfAxlVLKdGjaUtCW1xYsmXwq
nLpGMreMnBd00qbJz5gjfSQFDK+VUeISys+0fw2SbFODRI15d1uv8GRzmlq24NhS
jpq2jNvKLt4Yx8k0YK2dOlOvlcnnJrhGco+o5XarBQEZqJGZfrgzTyABMB3Q/pWQ
kVOs7GJksF2vPjGhRVZiSy+G029HSesYS4z/IuCsHqkn3TC9ggaTZO0d/G4ARzYA
E96CdAYNVN2Z/Od2hsuFDfByWhrkOsSQWGslTy2AI85rpXhLnfdhnDnuSDWd8An3
jptp9STMmKdy0+G9/7P2UUbQ0gZmTd+1LEXJWYnbH1haLCV8QeWMsTUCoZRk+cI2
Dr8eu/iWClQK5bXe7SFl4kY49CJX2cWObS/ueWulq5GgHB6itK61zfEXoIpkaLjU
oCOHTYJsaRa2zWQWI5PbKTzBLHQ22UYmGVPnfVap+7In9HouwtmJW5fXwY3Yo3L6
DOUw4QNZTKZapy62ERiLgtS174xEeiV97+9Cl7ZJzKJTLSFyGYxQtivMeQDGWF28
gteKSykKF5M/ZwfM0D5w5AtScU7HXwnMOyATtbjDx8IrHY2CjIVe+oEhCZRmSnAS
yZWGhZ6T3BnXLfmMpKXQx23j5FWEZ6qD7mS1rmSzTJw7LReV+umXqgP5VgwZaoPY
8UW+rnXa2qVloBbpozNY/DUdfidOlrenZZZBxQbTLoLTLmdMm/JSrsI76qrk1k55
YnH14Bibh6XzT2T9sOGuLQ8kp1150bRMnxkY0KC/Sn45GwrNIIbrD6ehcWhhtdRp
2hES1J6V/ApIKbWIhTYrh3GXGYirxN27Hso8TbTGE0gD9Q+QRY2kwEpr2AVoAv8G
A25RY2XpA9YWP3JzBPHZWbnE5IGwaJglKjUFV1MRZtQwNZDhU+CIKwPv9lL1+JI5
EhbDvhJ0hHw+ABtwOkaoXj8N2O8BKMmlqSnD3W8hcb9GBiEJjFNEZ9ndEFce27wP
JOh6BrBRZ7M0LJflNCBdXpTHunT5ZvkMXm8hDafRRQ8NfLILFo5HfohjrS2qs6Kb
AU7HEEN3fQ6CyROunu9DIbwTusqw0HxvT6Ue7GlDWbgLoHaPhgCoYgiQGEaNY/BH
7HbGCgEfNmJXletY7/9pEX6NnyS8o0MCOROmI6llo2BZzKoFBfOs6aUmdraxrkjz
VwHN/kmyudE3QHYDvKusVe3GU2bTqiHKASyc3tbPgzbq44+sUTTWGXwmCEksdPmu
wm7aDCiLprR57lpTJiQJE1Ofks4XD64E6LCkZJ4x0w54PCNlyOVmMWf7mBdYAfFY
bo88oG6Y1FGSyNUfDz/0vRM2iDILSUVLXKxaBIIQhODX8R8IPmUW6Q0AF+bfQDr9
gteUzcOcQ/zDnXUfotsSXjAFczjz2C+62oNFot3AzA4x4WWfHgKvAhEmtzLiDTn0
43DDKlLZNfr9aoif2Ys1PlzN/ET6FkcKsQ91mWtFFIjk1HjMYWFuuqj4PDhSsqQl
jgpDdq6tZq3a10bSQy0vKx7NSSm6/CP1DaunZ6H+wMRRRTVkzUv/jEmLVafXh53b
17zi0LzaWR1KOyDkCbyvSZGhQN2d2WqtgS/bnGb2jthCr5GL6nzMI8RmAAIQYHBI
U35h8lGLridQtNu/FUMHiBKkr2ubRpkUFG33aQPRzuky1b2bkyfOYw+OhM78G9ih
iWBCIxh1VGaECJgUZNPPBEXOEpMphCy1MJu8He9ShDlhoG12KMkMPfwpnfz2aUAG
PWikOSW+v6D8fdvqh7dxU75G19PT63E7PposrBzkyg4VmVIz6KKssUd2J1mb5HaB
TwiSSCPVEMfFU1qp9WFhrUHd5reuYjwO0VSfH6mo0w375vFqBh2RZOH7tw1w7mBc
tmwfTfzNrejHXi3508JZ/Yq8i8vctP3ujT7UOM4NmJCTF/jyE5VOAGbEIkRb3F9N
u/5cHJh+tGG7QRZBZV/pRR6aGRq7QgMz7uOXSy7UV5bKU8R925uZA04yWSPcgbIN
aWDHWLHDbFKmRJjLqmsUzvnjIqWSuaz56ZrCNIrPVRE/vl2hWQMH95y8ZZL/Hgdf
yptdqcI+dpF7864C0YOAyDEwGL3VSjXJnC+F7yBFuehpSroQ4EjtFHRIY63CGVGn
K8vqwCkDiA7p79lXEjxCN4gTU2YyXPpyB0Q0gQ/aC/vLu8f1sqm5U17sU+s3I90/
Mc/rCDSdmeEEwy3NGg35pUbl43AGrVtDe9lnvSi96Iis61jj0E/ISou1G6KYVUXd
YGCE161IEloj6P5I1mAW2b120uPh11tgNeixNKyci5Y+Dsz60FG6+1qfcGpIDk87
BmGjSMjrIs/G9EWFAqmxGXiOliDh07KdUBEWt/chBzfv911Nb72iRJRFTxWvUqaw
2znJDoL1h2njOQlGgZrSG6CY0pw7ouNEBWF9h9Di4kcW28dmVHJP4GYbOZ3PYLA+
3PRI17RXWrghpUSCCAPsfbr/WANyscZiaxzIMfGHGX4nlklJMnMJkakDPMms8DEt
FZCDIZOC5SVQhxC9FObfOQkTXLCxkUo6VyelI0q+BrfseSLlm54Uyi1C9oTG99S0
GZRzjP5W6tWJw6xpU0LqJTlSFSANQJ8s8sIJLv+Rbr3YTpz2GNe4xrCoX+91zmlO
1qSUzmBkJXJIPK5zdQ4/C5ly9E8/vlar836VZhMDfJCviY+pSgDpkzgG/DT8ASKe
t4Jn2UzR8xujkrCcA972GPurNadZK1zQmZXrseQQ783Bigx+3h3fN6CxMpFqp43H
+DBQEyEDdeW/rKlDcSKbAhKR2LPi5kiRpWVSXQKFNnsZjWN/Y5WMrtCNGe78SPC6
mvsxcG0zR8sPOD6W3X+omGRSEyDe8gAaxrT1dvhGVc0Pw7uPlzp+ByTXjzmhxScH
TsruuOS9LGrIi5AyaigiX6ksInfBIBe+xjqAhaNU4I5xscPXtr5TyHjUxTK+5qf3
IJiT2U5D63Yadg8U4fDZ3b6/LrYO6bNVMwrn9BPUr7bOTB0QmXoyZMt8dB8FA0C9
k2nHjI4UTvHzw3vTq6XA05SRXUfSUx6cQenhWXGPUMaR3rbhF/FHnaAUS8Q8CHV1
hWWQpTaSUveEmbqHBZLYu7hou7TPHzL67ViHMQLdK96bOa86gcPPw1yYngpMCH+m
bs6clf6U/2ZtNpBnOt/g1aDEMw3g8f/3uf/FlePGky9snezAEgWnH6B7tQn/UYIJ
W6nuEJ5DYOfotKLFU19zfviTVlT+xeN57V7YA95NJCCvXwatI1fmQkCPCnzOFxma
VX57EsJYSn8vv6ifMWnhfnMUdX3+xQNKx1c62SQJbcPRpEzOBKG/rvbs8TuKK1fb
ny31anz72zzBdht8Zw+pIkDz5gXbIquNWUoxo417MesAQ2u3DsQiFdMr+7bVYxlq
01V3XpgdD3D673ovUL554UkkBPkUx4x/ELPbNtG5McQJYl+FSAb8QBSae7g4QIf0
aIir+0yxTETnLzWtxxg9GSNhsNwWaIo9l6J8xUjhysHHK+eXK7fR4or13CcLXtGt
TqccV5ze5tfneAmUk9GNva4b2xv6Q3yICWdZi6yLMy382c5aOzPGoGmlV0wWV9Sx
nVbeIZpVhhBoxg7KkyO4rxRxK21I7H4LrXpIjaVy51WpP2GAdzol+3dfSNDhVP88
cwJFvPZESnVjPNIOo8kPY3zl8Dn+b30rthfsjLfdrG6P57R9iCBXitDoxbQ5yyhK
MNdHC8UaYbt+ixj8f+7vX/jcxPlWkukuXEb1kN8p/Nriqh+ag551tlJgnv8JtlgJ
c/y1z4rI8HKzv3MrcHYqOAljg0LLNiukTTYZXSn129H4zy+S3cTjICCLocAfjJZD
8/pd9UuCJMQK/sqZCwjG5ggL/BT00qy1nfk06NNQi5Y8eUD7CJDVq/ZfgsyeFL1B
k74P0EtgkBOnMq3p5rA34MEltwgiB3ExyNsgA3sNykFcNvP9HPzsYS38+aNE7qlo
fhMCD05QOqC7M0F4D7g6wn4Z9uOcPbaMdDQDyxB/seTwGgpKS3Xe/admXoMD0Hj2
FXkMvWiQL1rfsHDIgo3E4a5I2qzAmfi0rQ69wEeScNxGS7QaryLryQWmexB/LQ8t
KRCZ9473zCY59+/10CyM8wMYdX5GNbQJYBOSYuupC/LnMVXDOyVh/hs63blnMgUJ
mLUzczc/5mEEorfzLq4QQodasHFjBSeB6Q1c69YtcOVZzYzMTRI+8v9VQm/wp2By
v6eDM3dQ6gWCplM8waQIk+R7/cMCaQ6CfWB9Uep/dryauxorP+XZLh+9UBKUL/+h
CdKD3JS9ixlEhY9H2VV2y79L2ED4KREG8ZHh+02Jzjau7Dg4BCUcKv2hog/7EtjY
M4xs0MGtQy79nfjdT8tXehhpBl+ZHUD4sW5hh+NiJiDrMR5imz9iyNmDj0kzroRw
l5aXaOwsTlqMdjTi34+/BsCzyDRmfLBNiNMdODP6wd3lxaIjU8w//UbKzxS05gOT
TuXaXTYuKXkmUTB6ZoLmKY1ljcG0MYqwxjQIZIXS2yPkKch38e5U+8nQMPZBgQpW
S7PMd6QgEtzY824oVXGYFzzIV0/KGUJWw4iOhJCB+NrPj1CDaPAO9uMobPlUtRav
VyzQ9S3R3rJFHlGvidWnxEXd85DPFY5K435Q/N0FUZ5lEalcznzzFgeMiMLWdGfd
pkRzFdcQuJPPUzptuBeM8vSU+KmmU8dzBvk1LHq5w+iUnXF+uSaMjymHacQ+pnKQ
kmjDkg3T/WZjfhtum44yL3PEvgywNrFnIvsRDd+zATvsOJ52atJ+3/e6WxrAw5yE
nk4ejVDVyV2aeZcgdJiIpHB2KAGrAeJ+OFdI9tf7CEQcGFn2Recvg5CG1w1siDzz
DaWG8JBvzaPQLF0IpGurYc4LVH7T7HXKdLSjehZ23sfS7Gf4wvHjwZ378SEk4uwt
cuzv/dALzvuIFy+TcgfeeMLxeeEZNe2rraYiDebO6o+2S6Ix/1lJtBnpnkZzuAuP
PDJjqQA0EH5GXnaIxqQUDq45SO8PYgaHIFNZux33vTFWJoNp8jfb6DbB/PTHpjb/
hYDdnXv9dcdge+i13RQhLp9iciOMdINpwn43rv0gs/sfiu2bzjwtA9sg4r/YEWU3
Vnl0HFTFmC/Nfytb6k1RCE0gozuUYmynlZ/ubdAhGq6eOC7dS4b8cMhOTJ8Lc6KB
VYkTo3Pyx2hCkN1E36P6g7hELBWc2sr171BAIvwdZDOeUn8PNxyOAbIFd05FaSXl
UKj+yud7/USoxr2OWZ7o5S5F7o9C0PLVCQffJhgc4bgexgTN3ioFSeOmlUJSz0HU
g9XVDnnerVRduuQnbu3I66deWbugANl9QNDH2imlDQqC9bexDuwT6LOwBrtkO/su
CtG6DfWlmxL7UaBw7t8oXj3Qj8EnUdnCFj474U5Tor7mW7nYo7DSiRtDybUiA4oZ
tFAn1SXWqnwmNbKKuKK5oLNZ81rAY90Tq49l1GgGgIPFxqI4DZpIs7eFh2ip7jKR
HArIPcSKTqOaGrnhSMYW7XUIStbwBP8vc+6ydbvgKWv34dIMrhqv5dRYjmcOdMbN
Wywzt2nyt1MUwTaT/wy34qc7ze+3I/ZFDinlNDiAP6JmM1Yws/9SaF0U71XogPW8
Rp9iwiLa+iIGgLp9qAIh6sgNpToGJbP0qUUkZOHTd73PApgglXrvch4lc1HD1OAd
O3gwGdcSErD8uD4zI93NfT8mKO5998kYMdMycMouX1vKFlsoEfV5+2GsSCBT0KIX
gognUtrTYKpJvDTMviufkGDkzK0ZenKjabCsiQP0a25U9YA3Wtvx5NQuO458DFEp
ClDA/1BPEJbQjVNarmVpV07D9vJKjVCtN+IC48zK1igk4XwBpppgE8Y0O5SpLE3o
/ekyrL/36VQOMeQLB+AQwDNlnImB6F0176f/FPsEavoGAB7s+1Xk7XRC+Ppfz5at
6tXY9jAdRBy4fKMATCnpahzQN+KcOYHbbepOgNua15RztH5GbudITtqEg6PU0DfC
ahjdIe314UPhffR1XWqyG8+5D1oRBeqlT2dPKw/Ik10sbTRAOxBhMlMYiqtrSXyY
riFydz2gu+iIDjata4LoX8YjPa2OlWDx+CeiU1H11lEMi/yz3bWdJrmtt4z0yc4L
KQfpXF1IiIE5u5Evg2kcjB5mKA1t30Vkgf4+FARDQ9CSCYk/78nX/ArqK89eYy/0
yX0Sy9Rk+Wpw9Ps0n4mVhElZfzWj8q4b4SxGC5+X/VUj/qWFfpkEjx59/kHHMdbi
JAPUCiVD+1jyHg/4KUd7YG55tyTkS9+bIrVhvbSJBVMgPAyRoEUKZPP5uSKiEdBA
5RgrJGhDAMG+pCaOjdV/vJ3J2wDsON9n2GFG3rK0DNXInCIAreuWAM0ymOPwR6HD
Bc2NIB8G8sXs/oYhVQ7tYX1yEOjiAQ/Jji4ZqcluLUVeuJW1dRS8tSLI9owkKkCP
q98UjbVAAS6BmS9dWODsEk8djbcgAXewmI+4FPZ0IXpdl4LaKJdNoilex9l/uLz5
NP56x2AF3hLQR3jPjaGCere/Nh6UqDiWldu3IvQ8WDkY1g+g2ZNYYBwZhDVm2A+k
+s5jMK+eBYDRp30uebmYs+XJ+09qQE7zPnIE/3knxN6JFKZhlNevg2uvJ4cr0pfN
IX8pkoAUeivPVIpN6vFOAQKkYB1oL4T1P5hZ7wiHb90J5x/F1QPRodJP4ZQpdC6N
PQXC3PqCexE4FYInqh/jyu0CvmTiOcmJc3onO37a3bywjl95UAB+eMSxmzgrpX1o
XQ+xRmG+ABdD0T6oWH6FZ/FHqnsfh7Njo+qU7ekPgI53xs+MFpDfwSOB5ohyuogv
omIHbZ64bj+xIReRckLxL7dO404iuTCSfIY2B+iMv6y43H/SjGzAvcFU2IQhxpAg
fplbpnOUBtg2V0DYa8RKBUjnCpqM5y9j6CVkknWJZti3yircVInoARseMpNfBy7Y
0MdL2m42LWMoXRGjOCyyPH3fKye+DyzAkU/+b49yqEhF7uWmAlD2QHNrlznWn5V9
+Lx9PlqBjwv13jQHeDeNf3z0yNeHAvrs7WewCvNdkFrF8elKwXUdFL/TgAZh5AU0
gJ4JEzxkIGUkju8lfrDAxESL1kbHnhMlGnPMefqlSvgo7CM/ah7p7ldOuPCgu4QG
7V5LByO5WLrr6xoUe5/6goyp6MwWXl5ioofYLUv2WRNHWk2+i8oEoOBNe73rwYHc
WA6J2rUXH4JdXgT0vixc5Vqm8XOujZFsBHdD5MOvqmdkB0+9ATMuawXSk+hiyKP/
ey2BT3mcOg0Lx+t4AWTgd1RHaN6IsmlrLZELRUC3m/OVWivN1BKBbAklEAVJD8BI
xmVeX2pvL/1ca0TMtq4oVzWa7vC/7gAhsxgzmCNdewVSRbKeNQoWxLdvThy8aobM
1RooI9f2VDqBE3z3mMoVU/v2pHgp8ZX3r7xVLoaIrM+Ktte5P0lj24BJjk0R9cHx
rdFsI4hm3/dKJWIokrFVdte2eeSmj9DeXp2DJRoGpBk/s/4RLlj8el9TLk5j7QFc
fkMZbWXmzRWNUAcB2Z88AOqGAOjavVnD5aGTQgbUMafFYyYiMy+GoMjbQofarx8k
kTsxb5CqOf3YhQs6gOHSSMItYLrX8CXINLuc2uOuTTtrAxeWgQKApwbnEnrt2Tzj
7M/capKoMdkCr3zUZX0XKQnuGYSC0HLeiOcnYV4AJQCW0Dam9b+ollnWK+5yuYyr
1WGb5/tJf69b+cqoSDfUxon/aOX0biU7SEJr3Lmc2yjcy3PzBA2pyPEc+MBHBRqQ
BUhKWdk8At4hT9L+nu7rrpAtibMTknE8j+aXOOEr4PnQjavzocRv8r/UtdO3S6xn
53kUVIHtd3nYDSwX/GhPvyElpRO4RVsKx1ohuQXdBWuBIGmaE3wipqO/5R5E4y1s
9WzB0xpOxhJFt7XFHR4T1SoDagRDCvjsIe02I1VgIp+dEeydLh3OXJnRcMKiRWI2
CdTeEfgFcpJdNXAS/UAclacnjsPITE2xBxCNnH6F6v0tNbU/L8LB4qyN15PEEUuw
g5tU7rCgR0ySGivcWqPt5uHYHAd8LjzLlCeLG/By4sW3g9Qgiir8PzNym7HV50zT
Grv2GHRea4nDirLpEkcnlWbEfYBrfacKVU8GriM2q4n+umZUUh1LzbLbRmGw+aPv
AKyTfrs6/KhHM9Mr3mKw6rgP5K+RrmJMlY6Y98xs/nNugcv44Q2XOYjXxh2qHaoc
O7sRwgoGYl7tfik8p4unO8wVy51nKEvqBEJnRC4EHGxwBu9tXmLbHCEFCSUhSoiL
md/AzN/YQ/6WRqJJjgCSxweAWl09N71aDPGt4ucLf27hU/hAMT1Dx1rUXQp52VTg
jP+42KrHQ8S/CyJad48TrXiILKzf9ZsrDOWy8DbM2XXj93SeAv5TRJw/+Yks24+I
v5Y7yzyB4c6kwT8oL5Qy2ojmfQB42Jf3Jte8Ba1Fahrbb8PGwbSRHLzkTXPtXdH6
Xqyj+WN8nSFkkOx7JJFM0dzi/FxXxfbOrM7uHjAL/cY+Sw2mDBUSjeSEDTD0Ycd8
r5+hJrsIcj23z3Bhk5xx5ZCC+IPO1rqw5GSvAC5dWIx0P7LpjrFirgbGp88VaFWx
iPptoo4wMwLUkF/S1DajTQpBSvdTfZlqCrPMRD+RaR36KWvoNvRFeuAihHmQjKuK
EV9JPkiAqWMwZz+1rzbIKYfeAWtTCAFpLVP9zUOKCl/0ndOiLOimN53dngJT9QTV
9UlQ8ZdPMgy70Ko2xV8HtoqKQ+ujRQ3z3COImx/ZSPOikGGSV9F4v1tEX4kCVhdK
KzRs79cot0SZhG5kplvtcfckkZD3raQPFx5KOxRV30voF7+Gqfzc7XAfMn5iESQj
7tPt+4yzIr/VrfwWEYdK08jHfLmObZprm+RCglFWQmxwIs7b+HuUeGCr6442JJQk
nUqh01h7zFHO/s+JKLSSPRd02RfgPqUQmetUnWDU7se8mc/oVax0St3m4/+6wT7p
xvAmVgJm1IsvMmG5r0xmm4mG+jN2tEGBs5PsVeGmrtiT8Aw+rRs+qTEOIFtzDx9U
MatL0HGDz7Uioc2zHTnEm/QNwZzSl2t/pqoWYLTJph+SnCp8TRhexe2B6T5xzZ+X
g+P31hXICYbg0JonK4NSYlO6oIZI6dn4AJzvOb3CfTUafZalt5bdhD8flmt23RVJ
Zo2nJ67eqIfWnu2/3hs71CysUc8XXp1sOayUU33DvB1IR+WdZkXLzHS/9Gp4o0zr
87Zomteb2ICOFAEwyCbf2JkQNQQFrybNWb16BENTELLSS2evKrPrCTGVgD2Cnvrf
GdCXZoBQC8Heh1/HcpWrYHalHPBRr97Hkp6wTFob8Jky/yguCTID2kcd46RyroOv
u/oHvwFIV80YbWpWMzZ4ES4JBk/xJ0YjCR7O3cdSKGc4PLF5CPG96Dd3E4An7ZRK
FPVS/5JH4+ZOxvpgvOYlxBSiVJPJcd1JGsyhp2KmyDUhg3CDKacakIrjuReyCOHi
Fe0wmK9iP2vlcr5uBS09Vf6UelcC3I2jb5BnnqG6kFcOYX9xnNRhLpcoO4d2bmzc
KBm6EixduUDyPNlC0/VVg6AhtfyEPv2euNCCDhH7gTikUqcIhbc5WhR3cQqWDreD
GNitz50xm6+ukQEfvi6J0qa7SdHupgvSVXy9NqJbrnZEPkE8/BVC9VRq47iNqS/8
ockC1HSXx9pmY7l9O6KMFBmSbSoxYqipSChNl0lK25xPQm5hkEV2X40TkjP5ydGA
`protect END_PROTECTED
