`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2OxW7qq6Fl1uKnePGH/JFlvmYHGOfo1Y2U0GvgoONBOiL0WPpY5iCXyfoFeQ67c
aroBiZr1B7mDPWvjCa8Sb45DCe5BDkKmYOQ0G1b9F2qgZ5GxAi9hQK9Aomicj13d
S9l0n3TWTw/sd2RSz+JZzKyJ3eMHVBZwW6P3R6pYCA1kC/KvMckuSn4m9wsoYZ5g
jLmk+FeX6V/rSbetegKIcJHbBfw2KEMN1emZxBnGXE+tyw6I3WQh6UviYWU5OnW0
yijx71qVngzMuVBqgHBxpVL+mjjHo9cE8mPSwjrZZW7CtCSg9QuKikP67buECRvB
36pA+7E7sYMCJs8DqvJgO7xZyjOgdBVAmW30Il9agOSkKWvPyjXQ85W1apA0NaXY
nIpX1k1AhpCAVLK27PTZJW3F2n92TOnvBE8m8ShLrv/pWUUpiOjNLQrq3TopcKYd
t+Mfq+DLpTJ9xHHJg14PpeRHnzWsGldW3i72Ng6AOCjfB2PpfkvBh60nTC8XjJWp
Ya56AsCIKu/HzQIftKC/oY9nsz03QqzBmokiqWCooY98zMPXNuegsDo5d+vKctD9
t0W5Oa20FShPJocrLsOZX6nCBNSPxgawqt8rMMVfAdG9dowZbq9vaA9YAdOh9XU9
4DLiVWzz0ttmC1JhhWPu9CfboJ3X1U6agBHeNxpNDAQKNnMrdhE+Rz+k8CpgN9hi
LBb2QEKeyj69iRB2wRFXJtwXu34S4LCmtUjRSom5dHBVChSS1nLXsAgrQyFJK5W4
p1QcORWPPJQ2MXVpzmXoIKQOzkTIpSJFfnzVKdrdRB2u6xrBWl93Qf0OZLspfQA4
5UtYG4HL9NzpfTxCNbhazpj6oz1TYPEzga111yeINiwmiGX9a5dkWT+c28YSgiem
wdEUCgot4M6QdybZXNnUfBzXX++k3dOoUhj8+AbvfKd0MEDyO/e7PSjU2zCrzi5q
trjyCnLP5+9QeARh8rOPzaHUl8+gZgqGhmdyQJEdtxaE+IiTtFMQg911+X1vxXFv
5mJCG4vt+UT//8zM4HF+Pnwt71VwVGIAKz9FFHCOK49lt6XALnCwUClbIS0M4paK
9SZpY8WY97grUXGIOGNHUajk1K7nj9GFNzX0mYhkIL195OwgEW4KC8hdN0XOSKI0
ehj4VbLQyD6bw/zRyDFyJ/Lr7uPr5EN8oDiN5lQA1RXaxwcSif9IuIYPNviTFjc2
VZxVkKBuzkzkfimMvS9bvdjvXvKgJvfaU+NFQPeMVVrof9y/9917RekeElO9lfXh
7W8VAKzP/TwKlTyTbnSyl6ElMCzSHyq35jtC8OvcXZBON3nMcMlHVJXYTUmjfATS
PIzgt73v1CFRZ9Qdt6WLjrmuLK3ktE1cP8UwtnhxJDd+J9iAT9AisdA0VYEe+qpk
Mbbaa7FWEQLSbYOo8DUx3VdzGpR2EAz5g7sunHg0JSJWulhxmhEL1LCom12staHZ
6LOqSWspy4wlOnYC9OMoUywco2tmR4/85JFewictVx0yHOLEmw0ss3MHFBpmDW5f
Fokg0BqLm76uKLJ4khY0BGzFwGBoDefz3SW70EVSiSIiGHxTln3Ujzxk0ZYo+5ft
pLx0Dk3R3h3gSpP00fvHZ2GGDeMgY4lxcOoprBAdRC+QGO6PufaNodH3HwuHo3pJ
CUgKUcSQrCk4aYE1nMnw9rNXXxrPqnlSgK9cYaVLKrpmtJXOm3SnN2OzMnRKlNKi
z6tRgvXBfSvELGjY8DixIR4LJjYSpIsZ6h08IMLemNYqDrG5SCRDcJaYrxnVgSbs
l79Ztk29SbPvdZfNS87/ucxdQCNLBlOnZRBySkN3oG5VRpMVqj784GHAxrd0YdQn
fsLZVOEWUZGDHquHv1MXuInLzDmrccbcbz3mx9WkuzbU1RcCL3bB1nCUBPFdgV86
+tRN6uPsUf/e643ziMMRTI6XD4m4z5eDZ632WeBcSbzlWv9l8vrI+0p7sTX2chrZ
z47fu9bcaq3rUKDLHXdvHeX34pIY867Wlb1J7+rd7+wSQh/sD/z7mNNx55FsAfVY
8s6/x/xDb9Ho8Ycz9CJvR+AovJlxhOi9evgnUa/MVr7r7vBgqGkZuAMz16ATfhhS
01uf5HLM/HjxMufB1b7rWg44aj5Um2ZUWgjKchzQdrQF3MbPUOUyonDMQlz+/31f
S2lynM8YMB7GqxaApjC0TYnDgto1+G+tDRpq5vORsXhG9T/I9NOsA6v5H32UWniW
mBpewqnMrBxtXelEv2MZp97SwFVHo6RAScAWXnFRo6YSvQM9CZLcrxRS1nbdK45b
080CnDYEG1tB6be3S7uKz9d1YOwXFTQy8l4g867cANx6XnAFVn2V0rdygizueWQY
khRaQQFD2lobdGpf0oPrY3JzdXhl79tYk1K1Hn3D6j+jcrKFeqNHJUS/7z87jPSq
vkk0lqcrHG0CYKIivPUzZlLzlqhOMRcVbl1D9Y/AerwX0Epo0OyfK4RIjcXyZAS1
Lal4/gTE9ojjXNxixw099ckSmHN9gIVGMxmDk1Tdmnx444W1zejJermTcUDSV5W5
9V4YD9ZCK4yf/FnLy4DW2PewLrF+RqFwq8TT6qvoT2PQkpnvJEwTvcgTehr7LsWg
5+Eb+0va5qBNqk5BhsocmMzBDCdiGKvAoir5e8rnegpZuJOpr/EKwCNmJRKTJDld
xZg01/C7bHJKJHCao8/CZP946HxLgB1BvmluvICOLEAjixuwJGLz379TePZOUi8u
XSQjWbsR9an/18iIr/ieKr0F2cnvtRKMkntb8UchVuqSlcv1I9gEvDqZSP/3CB4S
nToKV7R1MsFINxHQwzuAPdpqFmA2YxnOywan1jUD6TCN+yPGAnAt8oPLZ8HkwARl
b48ChkN8l8cvWdysSRFJoFoZYKpi1wpxFDgMh4Jak5idBL2YzQR1lN2Z0gvSEq8k
aO0ZCzHj+R3u6OY4W2HQFYely8zE2cdE4nTqt+9B6rJZB2o7inUynawgOGUXsQNM
naVqDTzpxYAoVbU1reF+ik/npboIV8kuW6m8XaJfeum5gKHrbCarZH8L91yleBsW
1VVk72eNEAYdmHJwhj1Isagih7tJSR0OFAMHf4jKuVFvy86riU7fAzqTGG42h+lB
hUi8ci8neZ8ZvioA3zHuvl+SIrWKB07YAgVjDmRBd0cSaCsKRYrFfmx3sjHU1fmv
5SCf5brZzldLwT6XOSQQWw1EhB7rYtArDtRUtPDw4Ck2hzo41wH41xIDzG6plKnc
b8YVzgpiVtdF5lebJRRCxx+g4se86UG9JXelklZP1FsEaijdTVGR1njo00EUn7LP
raeZPAgHBn6X7Xe3yR948p8JIFp2KeIvyvqEEH9LnfpzwpL4mbVrhGtJbF2V47Q2
N6m68A6yfpcpFDxJjAdPxARIeB8+QTn55CRM7/W789p7xOGjYhyzrTIxhK0MFCLa
6FvbifRpVtGLR6fjvrtzWwG4eoO3lLQpmKQzF24gz0RrCDSFmFOT6KsKv9V2QHTZ
8kht5MNTNpgJpOxS0ZQO1ZILKudxa7V/xI/qnGLVXkB5Lxl07L1eMGn3qginPs/d
NDpGOZw5IMlO5+ObEmB5SqReNThLa2HPQDUYG1yuMIlwG+ssHqomjydmDER/KqFo
GCpQnMLvZNNN9hxJDhb/Rmvg/73BglkRs64GGvHUF9c0aHupY5Ep1ikvpc1E29MR
znwc/AMDT6wGYj9/J0Hf6RK8HmvkmuL8X7mpeJKhj+5EOBLdPYtJ2n9cvTzXi+q9
Tj1ef8iRbfWGYqbfOtCOlZxHN5eIV+cvnRdQWV496hPEQaNCkBKg7ayhGwWd7e80
d/3eX5PMiONhghx7DZ/rI/hXZ8DYdvhPsV5H/XQnSRYs6vbKjryjdU4QIx7N9XFR
VLE4LbuR6Ix6e/1B5NIYWDoqnTa2wTOapjuhW5/KmfJMkppZTz53+0LIl4Gs/u9B
LQaS5eZeKmNhZDbpEA7UhtDrKcOyzsJHZh9IZAmpCk49KUYi0PzK2NK8LxkCENhN
Ghon+OoA3R+F09JJKMrINsgKb5WVEa1pSlUD5mO6dUKYPnXOr0iGNriWItUxjZbu
o90XSL9ShpzMj9DwP9LXF2W0XvO1aHU5nSBodSAYP+H+vsZ7HJxzR89kIvxSPjjv
nIeGcDQz62gtoIaaEdaDoHELdD22Mg9YUq0BMWnc5wL8jlHhjHpVovwt3dEOlPyh
31D2j2nFuntCrJT5MZ4juW3HZlVpGGji2cLwNbVszmXygnO6qq4+htj2LiNzK4ox
GuyFKiNo055HLs7QOavizgLRKprdost+LtBnay6aUvb68Z/NzT/ccMtD2nBMnmZi
mfFlk1bRXWne6+uwRqo365eQpNqmxoL2eAbYPhrXrcCzxCS0MOksSTqGXB6uMx9x
6OcgCzrOdgae/kBl94Me6TJYpBmWNI3QNLwoKfhh30ZvN9nzavqYZ5DIGviCtFo0
qWqiIK3HGr20rkf7IU68eyYev6dn9uMtTaJ4Aib0Q7d6Rgaov7L2kuzlisvZFNm2
MbOln7Lo3eH4pff86VJxQeHCSir0+DTF7dKmrCrzjYJqPh+b14mHchf3KC1EGiOC
bHSbUvJmHq7zY/PgV6kSc9xabif6n2RD54Ggdm/+JmI7Rib1ybyffx4pvIOAOKzD
Ge3Q5N/E6SefIOegOsIZ4AtoM6TM7W0ETw5Q09K6+HnAmW4QTvp+YV9171KGzPF/
bQU25fHyM+whYZWqaRVUIcm70CBWD1PqPkia+xg4prlci+OYmn4nTp3T3dhYmZ68
xctLnzKDpGoFD3DjwMm7jCZEKS+H8d0UOOwZDVUYu6SjOSGGl523vD4NKkLprSbs
blTG4VKdYuNlQoEhDJYSxA==
`protect END_PROTECTED
