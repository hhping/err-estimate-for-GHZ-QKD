`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzUnqB9sg8SXCc1blByRp6ktZTFyLO7DjnK+KLEiF3brl8lDoHQ0MFWQ/wh4x8f+
babP7xQtYYW3sw8kVXwBlc+pxt5TCxfuoGI3eHVyqRXmuX4/GCtx0nBMPiGcfkoF
Ftw7Ku0ZpW3MPbvWqP8QZxkGwnRFrYxOq+lm4SeEMPOxP62dslPHDXtc0Kzo6Zws
15RW4VTnqeEMHRACsA1i0QoJosMfk9jCM13bXkiqMY351k8IWfIUbf7J8lW59oT3
KkojZvQi+V+jvSfv9hoesdpoOFC3zl/CCpka0acOZKHvbq3ycKKY5gHIibZgb1+g
B8oEpyHwwtIGf5QAOrCeiCxA6RJ3TI3P60aSrh+C2Dj4Y5qpHoKfiogyV2DgqHqk
7kaCmQ3vNzC4ofWK9MHyVrRZx8jXfrcDr0wotBuUCHexpsHJ5utZ6/tYOqAoAW6l
EwAlNgQELE2o+WqGmDdENEXadJFxW4LuBNyQLnjUi2cxV/wDKzIyx5RKN5TfgyP6
zsR8KFdbeRhgPSq4k5k4GEflFom/zo3b08G6uui01xmhjVBO3Pz7yAhL5/P6gc/z
uiE32yfry4ElndnCv7QTrRb3pdrRAp22/F3a2DCbym3eOC70Mrr0nnjpv7s0knKS
P8xr+7mTvfvFBt+ccjQ4l3jrtOxVcFCOY1w22Wx6Ha3hYLucXbRYFXT3QleVf8O7
iLHx0s7V28De8I1l/EnvWmxpmjO/rJryhNsLzRhtBqUvNl6isWZbHI/cOPGllY6o
23KCxoz0gQTVQpPXYmsQlGSSqBqGr8fK+f4skLIPL8Dzy0b1i/uw85m+mIO670nt
QAZcDIiQwF3EliK7VSaoOPPxw3lt6agvVkkoStfLus8KFS6XXUzBlKltlvuf9dg3
ytteTwrh7O/WbbRPNTuye75eM4DlKb8hB7V+zcu2AsWYn7GcmrjcxD26ORabnXjH
A2O+QUzugx7/v/MaUOED5X+Jqon7Vn2y+N2X9shmnCafX2sdPt9rdL7X42hPDm8F
KecwvGDW185YKhJK5UB6uuc84Mj+xmJZS1+2GkZ+OxTThla/8f4i/jUsHL18YB2+
vYtKV6IPei3aflgUtbY4lYX7s87TrN/GxqYYj7VG33CvjoXbeIvLz4CKwAjbEQCI
BugQfQG52uDZ0ZiaT+jXE1NCgJn1C+F1IVSgRUSg/nFnRu9t/rXTUp3oLGZnZ6sN
5FEvx2AqTniyVhKgnijOP7lFnE8+7rAImghUvXRsUuQkWDCHJwyHo2aQpfpbZSSn
9Y0gBGgBVl+5dn3khBqRVNIsPvImaaPpLrtSau6sg6FB9u6KE0/nrmJSATqnUD4m
B1uVxaA6sQgZom4PzDqF0Tgw/xEX+XLaNhQOQuBn6wAlDqUreUc7fyIZkPinPkdb
YGLoszjOzckK2BuRcnGKic2nX0zqULDz9yGq8szClWuQev8IUjbQ+c5dEOwcpkNW
h8sG+7ewhSOluxiesu//SahNf5BVhcq8wLMIE3NZ6FApYachUJ5/o11558AyRXZq
ZRIiquRYcPzQW3GmDeK0Kh6ScEEdcVtIIQZa+6f+T647+HykxJYL05Clf2y595Bf
xMkK+cHoKD2ZvwKIsgRhQZM4xrggmBF+gFRzNI3iIzvukQcDUY+WrNtTMG5ZPRq5
mTM0bMGy0rfTBRHjw/CO+AIq7cYCGOs3t+Y5iivb+l+XIHw1JHInu2uGcqliBR5b
eKPxQcICNiskvhrcZwe4cTCiz6UGRv+paJiNBPfPQiADi00Qt7XTpkkajkKMbDRN
MyqPt/dwU3KNra02Sz6mR+PxYxCPhBOabpvUDbeK8com28Zpy8kGZrgUvW2kOfXo
4EGx5Ery7TMhEruwcS+gZ8A55O2awiezSP33vc5ZUpjIBEy/ft7lXAgvFzzXneus
FUjh0SuTcyuXbrx+2ek9USsOOXoMMEzJgsuSkPV+5lLYZOxBhbBwPClc+XpeNfyK
OcwCDjC4XRR5AB7QtKPx1ds3Ebx92ZbWyKHOGeGBtSVbs6e5tZ13CiVdVuOwPXIo
aquHgk8fzO3dIklPutFtuglAi4ZmhXNQuFIepEOu/O6v8LILJTl5qgaW+LMskVtf
/kZIjaDsHDhPNlvjK5LeisKXpF9CEzEvWovuz2ETuqb7E1ZpAWjde6Sv0KZ2t++Q
fS0jkpMSKlwubmdpqO3LfeKkTbh4X13Lm2uvFeGw4j7Md5UGRLpSMUw0tim5WVys
ZzPz3QRoFb0mNSBWJpepdDTTVFldaALHRE9sYc6BhwCyoiaFUkHHHgM4NlxipQ7A
ZNWEwAfSVSiqBhaL+a6AFRCfZjzlikPfcXHrgiDqfLO0Sm6FqG9eOh5BR0V/uSTk
FzYc0sEw6KqzKFqa3ldJkP3nwHrGGPWog+IWSRNMjEazziZNBm3A9/GssZ9tyf1T
0oDtz2VcSfdUwG2aaOtYaeJguHh7oBWxYoeE8WAgmxdUr0pEOOqUYVLo3CSvJZxo
55DZqQ3pdA/kGSilAtqD2vdLgB16EYQm1RGu88PHM1+c4vhrcWOxjA7YZ5Kh3WTe
jlTFnIM46sKBKnvZWjT5Ld6Tl+kgBOh/9Qly69Rn0lWrApMESUDB82Mwpoce6ixE
SxUYWRUv03WMqVItrvIR+fj59x0TvMV6sOL6p4sr/FhBrS2N+Z9pQKgnbh4g04/n
LaiM2oOapldkW7AIuhLe6W1JXWxkbXt9ZVFZF+/Z67BnMeZ2FsIkLgYlurM7QMqn
omYK2nejMzG6eTROBrgNRJPicGZaIgYy0vilKVa1VsuMcZ18TOoZL8vXbm6D8bJH
7H77bx8Q48yGmV5+6AETfIU6iPfc4HT5JeqBdRdZP7GmPZeqEJVSXo0j5sVsJDeq
YJd48r1EFZ3/zLUVXorQfbgja1a+OusaOPLlhsURVeT1vMK0MZgY73vinb2qAVJs
DlRFwNu26zzdzKKp1Z+8b7kXkNdqHQOV5dMjgdYWL4Z/7G4HQqqkz5OWaCIGXPli
T+/+o+bWQMOa5hT1sjQXqqRbu0SFo9gtSMxYPpou5/6NCYDb+Gk/CLMa+03c1Kzw
RZyVu4GQckPizchgF9xKEqt4jbt8P/k9PasOFw9DrhSiVnKGsQkfrOgbDhX90VBD
1LMyNYbhInxP6vXoxhxfKKFMvi1c2xA0GPPxkvkP3XL1365y0Nt9CZ20SmEenTXK
ryILjIUwRzhZfj4e8GNTRMhN22yDqid60uVTpEFU9BvBEOyDlGa20/CoDSVAtfLD
lleKaz+LVtLkt/QA8r5w5mfldiDgvOTqLNrcsfK6Qxt3z+5QWTfBXBFRRCekFqie
z5PvQSyCR4b9vbIMvaUucTOhKAkTtNLwx0Eq6FYzsJPMvxO/PawlzePoEj7s0SOv
dRw3leGEEoLMv+/YZYwvE0CgYOURM/pWDJlBuyCApnIZTaeqRBIXyK3sk9u3pDPp
WCxYEIM+Q9BwdMHofZWn6Y9iwqMsyRcz8f6dK0Sl/vKEFNYA8jSeQT5BRtsekQF2
UXxP+amM6nRO6/HP8XJwwwDYRlCsK9Eb8ioQLcNTXjjGd6gOKlARSpuFwwnyGoZ/
6ChsXHLlqdoG/tQyP5fV+2rKEg5ARMF3sW1dqz7cVfbsuoveIRgrs4jiRtnBo47f
lzomXihM887IwtgSGyMpUTU2JoRM1aDae8llJbK/Xs+s3A4KfHBtBEy9TTa01KnL
hhfa0WBRrHcTY5EsTtGoqiF92ACr8JWZuyfEsDA3vgl0L9nHdqWiQNlEGAAAnvdy
DBj3yA+s6S3usZkklJSWtyd3w+9bxrCaTgnhs5BJc+Jtzsudr06pZArvUdIdBUtu
Hmq7agAgXRBFV9QFVvRiHdNpKTfYh7QzsFnwdXk1Hk3KvRmUnFXzFz+7yLgXZHR3
lGz9KN7XRF4lkMjVpktdLQVMjXmXO0tyXjI0600fcwta/wcSZajlojQkUIf/+Ln+
xyJiNrCsGmgFHbLdnpYkUBr5EWE9JHV00nSFS507YXXMirIVodcfJpC6Xg9Z/HSj
5BL9x4u4X5gT1kGUfXtrAasd//4hP06hoeCY+gW43d5MgOciadQKldLLPLLG8EMR
+Z4ssvW90MYib/A0X/P8FjpfhnIqLMi9/VdA72odPV3VoE5m6uJGviJbkeYVZJ02
R7fMtChNkV0Aair08OhyvNzrcFpJ1HbkCpIVVTpsGjxqlwyHcWHbM12TuKC1RZJD
mNvmxjBQSWzjzIc73gEj0lITTRukNB6RkTV1qhSzvVEwqpQvkAwLwFQZ2DGmEzoS
zDdEPA1jPo23IiN71VjMAnWvAVioLXhf6LkWbpaNlLr7inPAd+DkM9xnwnriPrKy
VLC9phWV+UzzJ/9Ig+CA8jcbAoHFfYU4ZKvt7EHilRelzFuVpyyX+HY1G586ysYU
0i7DpVRS4Z5Q2XCZvzSBXwtcuG9h/erh20TTduExkoUGqk0vl8b858BJYOgLwPSb
aa2ExVR0KISP9TWyN+xHzSPuv91U9lF+YmfhP19R5bR27dDOo+ZrAChVbvoKQi3j
LN6FvNpnFqnh4i7RTCNEYanDuKGpzOVKQL+Rmyzyl1X7XtUYqg3Blp3DjrKxd00X
nKbcCE/cr2XdUGVk1XO63nVTEtdSa5cNDMem8ldOwVIFcP3/tD4UVy55c5khoEjH
fqtl0Z09wR1XcFzk/VKiQYgZdZ3KsHaFDbWWyVK363EPMGSD7arYYie7DOK+sQ2I
BvgLSmJvS7h6n0OBzbOegm3+tNwIaUVXzTs47o1uy9l4+dJ6zm6wiSBml7HHSJfO
RXW7b9zdWV8XAafL3c1SRttnMSTwv97fnWO9VX63ZfbOZNKt/hgCUiMIr7J/cf6T
l2yvBpC2p0nU4hQlZLJ/eqn+tUhjLxQdmNMhKA2ySjbwoK4oWg/c1/KpYa4OBH6W
+/RJtzz3AUs2ri9H/C10mGy/Ysmo3zyQN+YPHwYdeOWsR2Wsk/8UFympBSqfNf/L
hiGLG3f+WESG1KQFSUIa/WIBTCXONyFGYqAMgLyAxYAWjGlprR1pKP10qdTYJTGp
WQWt3682Zi0gt+poZPNuH9auQxAucnGmsLF5jXYyscWi10+xOn4xfSEosv6MA4Vo
U7iPHcXFhYmvmYoR1zOxSOmpX4pnNceBbXn1IZ/mD37+t+veDut7HMkMfpBkFtU8
suRewkA35e4kmVoRzhyrFFeu21yKxnapFXKwTh54gmJCmaQHAWTdQ6nudUEL+wR0
e82XIt3DpRTEp6Y3CfN4eXtoiIaj2kOmcBM0SzZc6QFayffZo7fDDNSvxTeX4uNE
/3l8zOqmKlP7pckNK94OF17jh38HmCIZQnCVqvg+WOhHnlxoC/aAHJJKiemE9MoC
F+cFfbdzLfpwbZmJq/iSpTK/BPs57tHkTT3adcRFdfxoYeTgYnnbC1eXLn7xPntr
ejQWaBo08S78WEM3k8TzAuSGIhNKxWaghIns1slTIVk+NliXkH86yWoLcrP3VUQS
PxnNRR+pPfVZAVPbezIaEC/k007GhU1Cq6TAVc51wUcAjC+2PH+F/9yAXdQ7GLz1
Ibr1uCxfH8UY2/AzfplMALLBw/OBFC5RDX9jzTPhUYg/FlDf3Es6NAF+msoJwCdl
SkQ2ynLA7FFseGxs2TtGgkBQeFn5U1V1AwshrtNTtHbHEKSkLstRS72fgy11Pf5B
8v3Rz8zIIBWupOO//bpy/5HiIHK96kauNJiiQeRJgGiUxHW8vXzAh3tqaE+6r9FE
hJA82tEt8uVmHrB2uHhM31UGeu8rabG8zEG1N9wuCT3u2ZebIqDD6LxeK1XvFVHb
2Z2Rd6D2vmJmoqG0P4qpnXNdj8sJ0wynKuAslIrDywjmrtK2opJa9T676vwzYNWH
WiZ5spH9CxvDMqWvwAQAfoLf05BlTgt6yvPSvMAXIQ2THv11ULILhbAc5po70JJm
4VpYwnY+wu4qZNKyTTxZAYrQ+ZKEOx+qqO0MVyW7vz+wJzcmaq4XvY2ziwNsLGiS
5yUmuqRGNpEexFjEXDCUKw5JMHuCkybqwRurxfLZDp9K3c1+YkbHjTy53aDDT/kH
s/SALMJcVWA1LHbGx2fKlRN3eiVnTWNL/zyUTz3Qq+aF+N5lItvQlDIfFfD0+/C4
iydxlsMI7oNtLgkbpsqPoI3wDH+7ndgH4w71SA1AaYk6I1OrAKVO6NsggQh8qufK
6PkhVpZ8fDdFimU1hGXs1Fzi24gS8UyXIOY9R8lxEI0DSJL+AbrRtObElXFc8XyA
qP11/rNahWReYdUE8OszA7ysxuiyByw3zGLQPToLihWQirMH/sea1GvpAU1MD8R/
J7nnwj4/PDnhPhtzX0Cd9Coet57BbaRsOEbr2jRz8E8ooHauqzZNLSsmMI6zsQ6z
QHMXLD69HxMYSeRMNnonjtDLSKOiJ4eRFYZLRugrE2LUZvOl0WOhFSk4WQFS+rfW
4okEus8o4rCf+i0F/Wd13AjNGJFfxsfmi/HWl7jBJOYvHZRbWvS4KoGVAn/RU1ND
LXVh7AQLxrmamLXJF2cpR2gzBk0ofO4qsETLbYBCja4zyW8Jg6pHZP6rj5ZqMYAN
0sgeK0Ozb6ASntSRYZV2Gr2fnQyIJnrMoFb0RTioGJWhiOBn5Gn1WR5PX6oRks4W
V714ybPHsEm03ENoG6CaN/yUnrBulwJH6OsoPOJZPLnFjK4PvsSdsJ3Pk4l1XwR/
rbh5ksq5ZencOlceDF8IMxA86ooTfTpA95PULdT/iIENd9zy+L9RQGhmswkshA94
nXnE8sK014yxKYGxAoPIdeI8o+LAqZ0aNzP+qNcOUaLe05CXmru63li+wes3iF35
k57psFMdQUQoj+Tw6iMHMCacoBIe9logPaPwdfWfJ0zpvJVqIdiB6+tZ/l/kIzOq
D5QZrMmeE2B9XN6bdtPRk3XO61cw0ZnMay7v/4UQfatw7b57juCTS4H1UHD8L8/T
4e3LGROctYqREv9ebzKXwUZ/CpMwCxpImbrN3VrijFZtpSsFZzaouq/6c4U7XenC
erk4A+2k+EMYY7gzNqan3HWBt69KlkSCztfV3LWYhOZR+ZoOVP21uqanGCpAuT0n
0Z+6D9Qh4qpIhYJBh/BFyHaTIpWLBuxrM1mrNlwi6sATp956OHTBK955ZuSMTron
U5kE2GoOFImVEXG5Sz/XNOp/NG/cqjB1cNdoJNsNUSOnQrXgdOVZWAzdvRrkuK2N
wQv1GNINMjJWCZa74URgHEDhNvIx19eqFZI04q6rifYKimRFbvw1ALCvoz7bsZFW
CPfXsmaYt9LpbRn4LFYpQeyL9vH4lGFuh4Y8CNDfLFry6D3IwKth+fmzD84g1Rqr
1+/fOEDFDdfe25PfyVVy1P+1bI9kElyyq59lDt1oT3rrVe++RjEjoSG2r3jBHbTJ
kcEuQqBbvACgoTLHIzJh1pr3lNZnHhYCv98BDewgKh7+ue+pHZvD/QO8lPPtTqm2
bzHq1ZOzcb+9ZPSs5D3XjGfcZ9prfAay/VynYfaimt3YbRMtaEatf5MSYjnsqtEu
2blUYXsDUW0lPqC9bK9ehiUlhQhsUzikB2KM2a+CVlyMF6VHapvD0N+85OkufXJk
JG95BVGCPhKeVGrMiGOlcOF+lUz83y0nBFC8gqrRhvrjeMOIGBW2E4dxy2/cdXC6
jXQ7Hz2yw1K5ccs36hzFbc/Azy9gdj81CBEpvRqfx+fYGgEyZt+B4O6veQw0RiYX
WhcPlf2Z5uxk2DF+Av9aJZvjqBK5BkeZ5FMW2bzsnd5afF7WrJzp2yOEnRnpx15K
zjVxEnxDhINe92KWF9TlRWxIKM8s/QNrVFxUrocKiXYZhdQ6bCLaQYTsPisNzvzC
3uJ0wtjDqlm7jWENANA3fV8c+czc5kU84gU6sQK9ElcXr8YYw1FOjPDca7TBTQU7
aLnsPGCXxVRlmMI15BWgJjc/63jLuSJn63zFs5PWJEYIj7q+df0ywItD9+X93stz
Y744FD5bsPpitzoMdx3fvKjew04ZTg/hMGv8FRaOi+KNBWyAm79hN66gj/Ue1b75
/QJfkWTDODcyFfAWurx5qGmy7cnRNwsw1RRIsuDgO6wiD6c0rUFAtoq9fz74sKh5
r4OLQr+wtLVduY+Mdh65dXOM5N3zPsh0JmeJXLCHQjmoQ9XCDS/4TGn7vQWMAFRQ
lD6gYW3kaV/FnupqFYOGIx2KZ62QV+uYK+XRwsKDKUOlWbOvSGRpmhijAlkoN9k6
XP4p+VvhOey/2HuX/Wq7f6GTG8Es12D2Rq0WVN6ov9Ao9o1y95DBtt60osUIOzeK
75fCx8tjHpr9IE0lv9zOLbNAVILmu315sRU0Oi3TbCrU3ZZFxpw2x1I7V+kKWa3l
mxRrCA/ein0h4HMLEO+OBAqLD9sj/+Pm7WNyamo5wbbR0T9avQpzXqxcWb8yez7H
ikOQDGKDDOkgdmiBRp1y5lXRunDNhVfld8SWl7i1GUYDdU8kprK5GH9vBHnNiRsE
TXLz4m4bt/xQJNBq9iGnDz3lYG8IcaOVzq/EcyK8sEW7/MuW01DW++CeUt40iOlQ
Nlv779Ja128zuOFE91WNaa5oTNyj6sdS+oVo4ivixpFvAcBMdE1vXtamd2XX5feg
o++lJCLxyfkz2FipnPrLyY2cfguxYX472uszQOtifD3LoE9ze9mfvvJ+D3YcTY4f
YDPqHIumVtDfUH1ULKWeJjkC/w1NCClDAa84kyluXX0w7QwwfiSkLkhjypQbifF2
M+mBvLmQRgHf7edteWMtvVh15JcCTQ1WZdsBApBrBzGYZH75y8GjEVuojsQFo+4F
G6agWu2Ah73VSb/aRJV9QPNyscumNXQw6xkECbrdwZuoAYnzgwy+MYfg5SGHeNX9
oukU6x+YBC4JDjekxvAd6e3/ukfdiBKzHiTM5Ts+vo3jC/idkgT9uGbcUFfPQjgW
XTd24EZMmnxFOxBeWX9SaAW+wBe3nfna0CM+r+Lh91LvDwcJE2MAs0xXuxIYN3nu
hvGI29zyqVSo5TkpLqdO2yxmFU5s5mVqncvnGfBiHoyzpBe9F7q7ioYYijbbofsb
0w2JyNb7o+Tq99FhHQXAdF1sKkanZ5fPKSkugKwogWq0vf5oTl2pI1EOU06ncIOQ
rPKe+DAvhJPWNWzeCqehi5u9VrXjYH7b0PVvEhiut6X+ZKKx8P3F1iGixY4k7HE8
PGiKXPaALfcPmEdgkn0uaah65rhpSN1BKtucKJ7oa3Mu+rg+Io0SWhvABU2/+ryI
as+Xalkgrb6tdfk/ZIOmnBEJk4iof2hP5XeRkEwUov3iCdgQuJmQIcl6/Cv1g6Iz
WLGXqQZFoZwcDfujPAPYlZAF8F0O0qhSKKF01uQd/ryernSZCxFFAvHRlHQL42aT
1aMuLULp3jOpVJ84L7mLHgPqIwZyn5fXVkEgF+QJR6Mlkxiqq8O6ffWnMcRdheCw
wdQO9gkAyip9tK92UoX5A0agHCQ54OTxKkxwXD153YSwzvAMGE2/bZq+CyWWGJhZ
gOZgDI7OavFqZNRUKAdUlDhE7MvaZZnQ+WDvmfiVVF2Th4KZ1zPOVvPhCEblpa2Z
8iR5imkNJIDAB4UOuzCKGsjheGR3cxVdZQquWsvCg0dsClvZWx0SuO2cO8Cyx0rE
ojHGdReJuYnLblNIL5giyKADdKXcn3GwsWzxQYNuxEw5dNi56Qn6sQvVPPlRXxAk
8dOg7AKDmHLD2b0IHs2OArR6xk+GDQ8uCS1WERb06cZp8XKA+nJ966bs5zAWQPqV
cwB/qT/k2eaiJkm1LxVFhpvft2Nal41fCN/5V0FpLIHFv+2mWuyU1K7SGBJjy4ie
0H8dKZqreAaRtpKM9XrMvM9IztY0TO11rrAvCl9XVooHrcHRKR7RjjCRzygPTie1
QmUf+xIQbqe/Z3rREsKAlWBorAvkD5n+qitT+zitY5/k43ytaXUjbTqXwiH55BnN
9N5dnmbb3pwTAHqD/8+NCw9mlosJ14oR5ZcGwfNzC9Xwlq2LPJg5z7b4usJrk+ow
/z0XMn5MemxleM3SecmLb/ykxL5ECnZRGyZR4mFtmm0FHY40xsla0Da1aj79Tthw
sDqEb1I1kNQcxNQpaUB8ljRIhf4hwVo6wjBTW4EAQwLIl6oQ1KkV+7GQz+gLUr5+
ipT9zS5IK0NQvOrilvuIolwmmb4IzHwaBQr58aoTt05zNIQGkfDG04ixTrNtLs03
fn0TXh8FEyhbJSxdnB+VbtYx4UDc0qv+rdBlfgp/uAcuFZRFPi8ntpT4RRLuzQt4
CsRHPA6qcAzosBLxrR2B9MzhiAfIhwlNz8QDf5bpC+P9imkm0VpePUBQeu0bjh43
sFdrrI+0c3C3P+h5g44leVbsfp1SRuAX7AQyFVmOyTb3v0xW2g+BwmMovo+Ai7v3
UCNLj6KETkFQog1XWvMWp3Dxfjh72Ndkp4O5nP6znqxPMqucJoZnXlK89URPfntC
U99kjDZr1ik/zYkApwKvrcahbWHS7FgZRX/eIc5le3yhwlU/F9trbVQKUGfG2OWz
vSOXhWFthWG/85/8ADwfy5ctecAmlS/81USNqufOLtA3TWEGwOSFRJJ9qoa0IGve
ZhlgLxkigf2geaswOavm1ObUsTv2Jdh7khPAg3vibYtfSOrNpt0D3fcCO6/0ep26
cbwa5kkK1+b7pNOWTwVnzuEKfgbELLxdqd67W0qMqOzE985sJ9m8eaxVyJaFhrdo
gtVF/pCSM9QEJ5S8aeEcmgoaZi0J2/4cSfFp6F+YqOljtnWKgB1eS+2oCFnVJlWp
qyAzoOe2XO1vQWp6C3RdOYNKz6R/0Jdb/7g0vRROROsERwmLHADC//ZNkkXAOdeH
b2+R6+JQapKwv6jVnsGc1p5qfnjSQa3VRZWlYwBnRPCvF1tOQzkFDm7/ofhHHYBT
KZO4UDDcdXCi7V1hp/HFoL4h1mfO1+zZyiY44clVI6N1UPyLmO+jKGr66PDUELeV
wd8Hxz/smwkc5PgPbIaIi20BekQvNsbgClD7ryusb/sHxpbSho84RmZ6iv6NKfWE
c+9SGrZT7tljSzo2YLdX/e4++P3xCHEYD4C/VvmaSLMt0SEQHbOO/oFMrh1Kh5t6
YcAjawPrXN3bvABXBqMRVhUIs1pHunCWrm/4BIejjtKA/ffu0GwYPWbsBOcHXzxd
gVU2n0kH8Llf8TG/RrKqCTYtTbv2i19Xub47gEM8Iq6u3ZcPAvf+M3hkTeUmXKOB
nRRTAwxO3E0HTHtBlpb/s0okM1q3Y6YN9b39egyirb/YsrGrdiFVI0YrTMZzh+/e
hLlRI3cCVm9YfIoqSWw03XG5ZKlaJGS6u5ggORt+zHEbWEPWIv09/8NHTKEb/r97
f2Cn1+qWvcV/lpDro3YFYcgFRKflKQW7gwiYQW/6oJrS+useL3WrkLdOupcTUgmF
VzojtlFv0qZ7Kc8xdFniuGUw2VZUYMY9t1HdGyStEMVv9sNbE89zRGj1PdAWbel5
DSkrVakDKrQHhwCyTjc1WmLObEzCZ1moeCuk9G7ao1nQfgx8CM1b3eJCcE4MF6hP
Nl0WuclUB8HgyAHOYTGtxuOX6vaLVHYaNcegHpc4zILTUoUkW7FefyZnI8vuUEN+
gyYacVoJ0IgxBJ6DbeNaltIDRWPiF7G0FWnevj2AaaB2wXLMMEk3ikvjzpV0RGw2
w3eM0ZKT3URoSG0f3UWFQV4giUrvg5qK9sjOqit0NF9MPjexBl8gAKp5XdRBeZCD
PfwTSZqEZCdQvwNU1G2n5wCmo/lU/pRsOi9pK2m1nDH3mb9ZWC5vNoJjkcoWS/Zm
Fe36+CfnN+TA0mFB3dvsbVgJYlqcMkiwDrV9yI+yGvJuWd2Ejl+M1S/HfSnWyVWu
aidy2eWWYhdbU0pUkMaqny2gkH1OFKs+y5J9/2KCZRwCpd9/TbzlP1SsAk4fGJrV
8IAs+VUPZbftSDg/fIQ1rXi7lA77ZRu+Lu8oOXluzhEndJBwLWS0o6/iom9tvWoR
j0Oo15tNt447HqJYqh7aokERbN2di4vnvZ4kn9rxbWSsZ32M7NW3v+hMOQ+RjGHT
Un64i9ZUkgmRNayTlsyBRWprDCAxeh1FW71+2fyjdfuac9lEzlIJVOCMLfEg0tIS
iSuDE4pu/aNj/H+Aq2YoLI1qfhCtxkHPI1Wtz3Z6cpPTlUEK7DKaGZ/uSsKsYUKj
3Ii9lUq7D/H3zMMQQcMwkAECDbVlU/NRaJauNrhoNU08AKJ9s2Z8/E5CXjE2p/JF
346oou6Crx7EjBEWuBnSbJ3o6xrz1cvsfUAInS8Gb/K5l7A5D6fMpYlFpwaGhl7L
zhR5WkuGcKSybEiA1vV2ar9sT2qgggsm14a0UpTU/PYVQZ3R9J+YM+pCXGNnj2fk
jONCXMv6Zj5zKY8L6tuT+lI7l65KZXz+3j6z+34dNWsuN9miitbsnzPor4Ulgf5W
WvYzVmCHHH4xax8mwxBKkQ25QcbyMgLeM284yBoZx+yCxINyxoaZwyy4yUXC41UE
hc0VyYWI2zcj9vFTPjRuF4kU2q9hrFGwemgb8eeQtcDOd1dH9pnoEt5EzWqLFzma
cRXrfAStmFhXujjfHl59EHXYnqE7wJHObVGmi0cyOa6mSVVfi/hLu7OuO/pf9xJD
WH5Z0cISlL1UksLny3NWRSOjwtwm8RryDA1E9l4A9onPIi3paXPj5iM/w5g5Iwfj
2VVY0Qywd8J+X8y5A/sO2ikBhcoKzyT0b5ohKdAFPm5VFjeuw4BZA8Y7QWf9pqsy
O/LVbKb4bC79yZ6ssbbJlam+m1iZxkoMzCN6fVYBddNktSIY7aY1keMQvoQ4fDJW
rU4rLpfOGJhYYBhg4CQzwAhDP2+oRG5cv/tlNn+I4UeuscqiqBdqi5oRg3CPFXgb
BGQ8moc5gmKUoLJ0C8OFjNDEnofqYprk6Qd+B1zM78NKypOJc379FdUDd1XI6RO/
BmxT5RyJ0ruHLWPppj1Q43GzhZZ7l25hT9hzTGFU9ModVp8sEpvPiy26+lUjIlJK
fIa/Bl88TW6Im35kxKdpPOKleO0/dp8A3CTDOMB+3endtBx6Lg5LDKd9GkAbEENN
M/27F2VP+mRE0fYRA7VrtFnCF83WdPsLYHeiB6ff9ybFyhg1ZxJp1xwUATBskWlv
gvqlYM2VTLumtIqI7XSCi77Kj/2MflpZCKno9VlHb2tLwhaPTbs9j9VNyTiqNFYm
9aOzxeZJR2ouREmS6Zy1BTn8fVt7GQXdcjsmDe/t01gH3obZ188CWFBcpr73hLQ2
A/pFvkijwQSgqpxYSzKrzip+6wA7h0C+r1uNgJqrIyQ7A7ZbkO3dzhGfhYf4PmjM
4/nxWIOTlXQoRVZI0i5YOFwxoMAhztel64Rq/E8fl0GaFHfvI3Wd+GPmb4eT78nw
RI9ao+VG6PnqPpg0COYqmHVjP1U2HSdw6+imqeDxutkdFcE+9vD4VlSNJEm8I/Rc
l1+CaowEoX7Hs2RYyEj8g1igbk5tqVbsmBsZlF5BUN+cVaNn1iJ83nJui/dmuiR9
LmYcuEEbxN5nAkZcCZ7rNovHtc9S/uly5WMj3T5C2JJ+dAB0jYz9+KpuHqZNwkSz
t9N0HsPIi/q9yRAG2dRFvcvLmNxojTl8WsrV+QPEsepsDLacnaWExChznuSQrvHF
ztSSLfNM9FjCY4l6CulatYXUOpKKU4SfjJUtfQEXkKMDXf/UHSjuKevB+wU90ftq
D0rjJMOmIhuoBIcfnuL8c0xvLD6Pf5MZBKtm9/+DFUYnxFWCC1o/VAj2XNS7u02l
iJrE/zDUL7/x7OzRGLd6UOV5REf+/I+N3Dkmv1CNwiwnF78HHNuoW2L/0RolMIO6
+vwgHzWMY7Gtzm0UDaqdd1FxzDIr8Jo+nvLC5R77iTOme5SYNwG/QcJ0QR5qTN7D
YiJd1v+HE9vjinTiPEzyxOXOc89RJg2iuMZCpTRG6p0GpohRFHbWN1bqsGgevIgr
cfmvF2dFsiX0+YACk7z0r8zu1CN/xOFBnuE1jFVqgt3Q9x80zaBIt0wZ4RrFrtAr
sR6Lozcr6lxCkB1cujQkw7HtImHhn+0WFsnofWTZCDiM8Pvtp//F8QIDhN73l/av
Z4H8hvtR0GMo0UtTD1IBJtE0+qXkY+Sbajy+zBXLFbnnAZJcQVfJMR6QPIP3Q6Ih
X93Z6VRVvgqeTzKn+Vur0swZpnPRvoQnU2zdxc823HPhAL/ZkCI5BOywZTW+KGPj
iQ9Sdz8N7ie8j1l88DCocRyd7b+Fr+a6jB4/rWUiOOKYlQ/9kVBsexfSSzOYUjmA
omUzJy5gg5+Badejv60bxN3rns0Q4v/Thg/lXoIDZngzTPliLPdk/w3z2Adk/Zqh
s181yGVrVkwihDnlwUzR56R8Pw+g36SPgYU0iqD50YyuNU99CRsH6ZRWrbH+NYYp
nrG7TbIhD5UUvwBzzoJvoGOh+squo7ufbRa5ibR18V+ciO4B2GfojE6hlYvobQuP
1j3wnW0H0x8UrbuDyY+Xdsibe+hp4exQcd9HrOja39/EYdeVylevb+KLAmdnTOx+
7R7stdIoUeytY/R3srix3yYkHLbd9K3VyGMuNpUXgXuEGIrh2MEZnwGLHEsVLyQY
RZc9QwItiBO64uwjcO84OMu5rJhTDM3zxhtY6y+Mu/SPQf7YrozrrHI6EotIt86Q
DZkBblutmEB/XxfYYv3na7LBaHgUws+wEh2f8QbdfSlDQ3wjAnbG4gEwaf6GvE/w
KZ+X2R5/0mxnahEd0pc+8PlyB5vBo61ytYmkAExUhHBGE6bTwEn7Qtxzh9yEvZJq
nZHgt7BqHZabQXJ5x38RKpCfz+wSCpOWog58c9Dz9k5RK2Ui/GruVPoPtshbLwbj
JEj+xVKusaX36fbVe99Xu9GZ9r4AFssc7c0N9Y2q0y1xWcKoq6pPF4OvugK7tPKg
lXnSBC3GuOeb/3b03zbZhWtbf2PUfsVASBaeoSQTfTuxfbgi/fj+vGNulgi0WHJS
TCgvFen/Yk4SEH0uLZaNxkgtiwTMoUyU2z8YMaLBsF5h8kSmS0hGwmjC/Dbt9fQ5
CRPUn91ZA4xdH/djw7NRk6UhzYIGpQvxrPHjLZ56uN02ZlN7B4eP/FAN79sVg5RM
bbzMSNbrRpktSQ2MePz6KAKjJJrvSF2D4Qab0DG6u6ZNqSbhyzzPgy8E1sFSwp1l
yZG+kRRuw/zEH586wYAQk5o8yxdPBBrIuUtlgtTe/ZFXNhnk3q9smyrWmyi6j9nU
7kFB3HFMQ4ovUUWcY+y4VoUSFO31NiiqKuwG2qiwatxeKh0i92mgvgWFCbBxQz7D
HdATLGqbyMlDiFwSNPMEjGxi/+J82SL5xkfGfhQ9s2fbnkTGiBt2scIuX0pCzdFO
maoWIUwccHlYh8GWE9nNpkofX5BYwpojHaoD5DR/2Ti8LAybO+j7iBIs0FZThDvA
5hM+RCYmrXGfJnvLTnYN/8NRAKfB40kcRzpsyzBy5Rsn2zJYXdOTgP3zxmvzB8ul
4P75DHLwXKjDNFcb0APHSWKyCsHGwopV3Q0F+DXo+djv6T1TyLLvPVhCU7qJJ+UR
FZLh2mhqNI/jew+1s4bEv2NantWjW1SQXjZmhV5m3ZtfQTSCNe/rN1zdcD0ve+lx
q/51MxidwgG8x4uqvsxfxdEXXYebuwrZjFLTtJ1+ECHyj8x0Kq8ze8wTeUzANuZW
fJejTtGfdCitHQNYdaAok8GCpGOLGouuECyPq55oyoCmc2UPNcdOmp41ao+9z5U9
Aagmi52WfCuXsae9vYfije12Q4q6d91VRAKLxVkhDlt25mT6FRUZ3FNWY2wIFPgI
2nIaeXKbGLlIpmvaEUMM3PfI2QvAribSBENJpT616U7C/3GtdU7oXKZaJYX9SepA
C009v59A4yNU7p5EEOJfZfG2CogyB2OaJfonmgte8rBxcqzXCZoqnZGEgrncABKz
MXmK3IjrCeVqWyKHixv/9+uifNq+falhpNKdegfRL71GZSxV6F7+Wpi/yD5aBfII
TI5jf1LYakc3ZclSQdEtXh6VXRmL1dGxRunMNPsGYbgholZ9vHZK7DbZldD2M/WU
c/LxebuZT68hPNwPVuKj9HqEpn4az+Z+klQGzZaFvbrtxG6Gq0oFUwC0aUA6/sfs
eDr2uF5ANyHpvyiWFzsI/ZkghHPMZB0gOiwV3n86iZvLxFpiO35K02/5rQO2gMVb
/BL/8+lnAQG3n9ArNts85lnbdq9pMcup266dGPHA6/b4NhhJv+1h5jbLzSi833ZD
gyapELwmkx4YukmAIDdPZofqjJ8emp0BBTMrf5WNofILJ7n1zhoFi1KoPhaV7cBN
7S3A79DJt4WGCaecR9yg5duZkaEf5T5QmoSQ/T5+w+QQkaTYBLhSzbDFvGyiUqE6
xGPDug6Z5cxHP4lksWjtM0pmyQi+TVlB1jxUr7NpkbNEkhwk6JHbG70LxIscneWD
l6eqd8jvNeooiANuhKc//2TNT0KUhYmJfMJ35WgnRHd05RPigtpgS0jjfTuoShep
RsC1txUEaqVDOME4go6Y8zMgfXb2RaRRt/Z/TNxHxp5DWRw9ZX2TprJIJXo3osh+
NqopQDQdafz4Gba0MLUAOfssmBU9y4y0f3DvqQwoNjW5GtJ/mwgGdyXCds7kUhAa
WsUnIwTIybEA0upqeGc07X4srOAsLYVobk6hDM6KUsZpGzdS5ag6V1Me799X4dOt
ZBNson8cbT/YShs7jbqI068WVyoW+S9ahZGjIOYsKW6xlLbvkvk/AeLlDNTMEpg0
tRWk/AtLqe3ujpDiTX5r2U/L2xKeTivV+AZ6e83xjITRCzvK6s00bBRujG+FVqBP
Yg14/ETLyI2Z/AkvDoqYURVtimpxO4XXArSaz2eivnvqqM0NVzcZg/EtC/pXhH5a
kpCymQPvhZoYH35F8mt6912rJYGNfuzk8bhZEsIrE7vjWrgo9T7JiUptQFby0yS3
Nysw+5plKEobG6BMv8EAC2N9t8sN5X+QpgBXUe1w5M2eIKUEc00DYbjdrQ41MYC2
dphcxu9w1656n5flVmFqjBvrbc8Ap4oWpSLMFg3S1cc5up8K45grhRKE7VnKBfPA
VNJ9HdX4DgliDj5GnEnkj+Eg42cPrD7vjEQrvcy9SfS/pItbJun7rtnZ6X5ygQYu
4qqru97Dt/AVkKzVEVbMPjNuSdwgAUSHt2N/JklNUkqXq4PusQKNdG3nA3ZBRlkV
pNg07RU/t0wQ9hsSpoFjGD7ShJEGmAoLumeyzcrawpJdXpgB32KBC33zCa/G5Pkk
IIdl5MYgEGlbXtKRmQl7xxD7HO5wsg+NZdpvU16YgnPoLVXvTP9lzKJC9ASb7Hm4
UZpN6/Wbhk5I2vA9GNNmnYnbXlakoSxagq8rrLxkQbg4C1CMjbpS9DfTI0/oOV2t
elhCWeWZvMz2nvHa1xh9g+qUXMCo/LCuNxIJZqLEVBU9lekcN99O3Kh4T1w5VS/G
CTtWxn4GsT/BK7CafuZvb4Ds53KHapSfLR31HheKI1h7MRsjtU/i+BzQBhyJwZGr
swF9/Uoz3i2kBTTOVVKH2MfuvKvmVf+YdEBuvq+LGa/wwKwvj2I4w4MJVrxnyrSf
WMPGOHX4FhbnvZwkDpBsLoZYTZxFYiIb+U7iB0gofr6qxoCOTPPMAc4CQMa6Fk8Z
IOmmwkIUBaSobjcKpv9auyZ3ArKip9wznBJcBXoIGcmZ/hyocs8oakDghU/JGF7S
Xkunar8jYrsLkapzw9Ba2Jl9MkYNn1GR3D8PQNC/IxZ1pZVlJJESAlrl7WL+eoMH
ep/CEZ55cWOqssg90rCrohP4sKWsOzvdN0RVuQSeKMuW6w5lKJ4/qQfnP4B3xqQN
CXxV/fN277X/BS3CyVvvBA+sqCZkbOnwshNmSyabwVx21EnQ5+R7mgeBChzMP9Mm
GFsWph2+aeLmE9s8B14qJrO4lvlOuyxmPkMlPuuolmXRtdIQuPfXzegPy7hEHqGY
Ld+IfBUnsst7P58widEOybt2eicR0wIuBaoo3l+YZTnHlIe2gfjEU+KFayWk6tGP
q+WBY9nkmzqORgXwy9ffRfL6tiHbmry7jjp0+3giHhaXmdKxkINJ61KXa2buDgEk
fKVN/PB3N4hY4pzPJbIVFwUZaeY3wI+qXy13L9RewVEfOF5dZZ1ojXFPIt6mAByK
6uZEu6VDT9ptuD4z3aBGQIo3dxNj9CQqZt8kWzeotLoSeVSjVHbFWIGkY0h+3UMt
9ldaKnxqK5gh1GJphoAbAiUKuBCqy+HUrOArp5CC7Llg6b27JRktLQwJP3JYUEME
H7q7G1HQZ073XsVFLfquukGoDWJg8Wm8Khljc4s8Eq/Pm4K2SEsBMqxRHgs4fmqG
NASa5bbqKNuhcyKuLb8hHcmqHNKt798mtOb+tFCnyV5N9+obhX+y8YebTb7H93Ah
ELYNpE7Jrv3UKFzQBOIC1BXLQusIAyaVSrSzJQF+T+SPrForBJT6XBy8WJeLTUCQ
3N/RlszCFF/koCnxUQo9vio7Bhe7wTS5BsfD9eGcuxsSfa5zfa9uNpF4YDlT61hC
520GoP5TBfyhluEk2qFjux+ghhpmOba1ltuqAB94jSGcGCHOkdKjDFIzCfkbrWkH
o8hgq0uwpds12uaxkkUWT3ulnIx67JFIRz7jU5syk7nvBaIGgq+c89Yun+n47DdF
6h+B7nC/+ZYf92X5mcGMyYEklt637qwddYgWj9KeiAVKd6eio1HcWeI4KnSP50dn
axNjsRDZ1jdUYrVVBWakwNrjj8IsEvdT5srz1HyP0kgrBdM4/AIlZfIGeV6F83gx
VcxJGZKd4llhtNTpLFuEMlScl+EXOEGCDOfK5QbX1Bl4hgXccTB5pOxkxGI6pNRn
4Kj5mjihqUVrw4p827xDWq6HeK5Kdm629XVqcR6TSkUW/vqHfF9KKaDqhVmqgPoz
+pjsFg68tz30jWy6CS5gqOpJLcD/HY4gk32Johe52R6qwz/1+2WasH7O7HqNrD4+
gemV/9UAKvI1b2gC5T9wIH/MND551P5KxPQtPVQzcfYpw5VDd+xmZH/dn3RMjdrU
y4tnHhDub0vfgXLtxfNhNoqSYFNns1MG0BhzeCPV7yU/Sl4fkMT6vlrIaDtGqUzi
bOc8F2Vnfc8TrwMpXQufHrIpRKZk797snv01FWQu6HEmNvQ6t+JLrkt6OM80oOBd
BJuQJp24LDzFXSsea+FONHt0T49eTOvJAqtAuRaUa/tyQ0UQAJ+MY5izLm/5tGJY
+6QVst6KkfvKUVfBtC9Bs0MMeIqhQatPYZWsDLzBF6AB00xd9J4yibRNNHLvtne6
gm1YDKIJGoOCck1SpGu4KxRb9HpxCdQ1TYWwVxkDaETXEGK29tC1tYGYac7rppXB
gvSOvwyrcdnKkm8BDs8Qdov08LqRP3VBDFWiNWuQJtdr5yC4dkPiuU2ytD9R3gSN
XkU8AuQ1/YB8M2e4ixUfVGAuAHKf5nJ9DPOUEYCjQfJg+a6lCQryzJWIbjDAjfRv
/43JNuc5bESE9TBvMOJJTHJd9ycuJbrRybnCqXri8Abweyl3OzWFVDHyAqMpp9Vf
umMSumZrGrYYS9xdq17+1jodI2mCdLn5rPhFtsGdnA7ixDJpdRG7m3ObVM9vkxIW
uwYlp4a+O17L6DgqonJCWultEnNojHBIVSs8DNHxfInsCbpzrLQsLnCIDQJMoJse
eWwmvZo6s4vP/QH4K5/AJOmwW6LSqH9FgdtcGSI7WnMq+Q5SJvoY+ne0uIxJRYr3
Km6DHR8YTaBLT7OhwDgI5V6SLpUMyMdFThR5fhGGNdJ+Rz6uwFou2tBBkdS55Rcy
RlgsBReI5ykIZf1gmalOwMJvWof+URWLFzYnq30nqcNLl2ke/RSCximYnyAx+EMj
xHcthAYeq9tCtg1lz33bdvFsGLQ0+4np9F+sLM7pUi0v0wU6BR3z+ETxwoQtl6ZQ
EX86s7Q/Ezl2ETRR7eMYuRFwUnNVxe+a1oMSQYX5cF+CCBAxxLOcmEOL2nN+0pAK
Q4oSVXk5PEJal/13I0krMa3YQSHwg32wfb83MCxWd+Ez0RGH2oL/8j0l72jdAOVf
pnhazSsY88jXQui709IIZXLLq60eEoieA3Pf2B2QJfKKOI5EW/je3WH6bGLrc0lg
tXAhYmSfm3Nj59W2DLhe38opnlHm3ZE36CjWHXclk0txMvBuP5uBe0VZbIgqlYTg
D0aGM/a9iuyMM08nOP5tQvEQDOqrlpS8Wv5DQ4ocJZWE9MuR7h03dTmhRcrgZK0I
0LKmk5/SvjpiJHGKPzlN+RkWwXNRlB0zF1fgF3hYUFylQviLXACkgoX9wUZI0DGC
z1+Cw8ufzHLnJ4/dS/pnrPtJ2c6U7k579BLugKXL6n7PGu9nfZMls24+hVW8th+Z
IgAFRbr+AuAVY7zJT7Mcbug1bX70WqB/x8y+eaHsAWUw4HQOLBOLpZkg+rZq6TjH
PO1M3usrzRzuU3zAzSrPxxp2vnGOfyFvvToSzxdxavurbm+j00iRhZrew1DESbO2
iNBgHBdjol5Nn/5SJ4GJ/TaTZr6ECiU2umtIheUXn/44ANejMPPFIswS2h7JA4gs
5PaUOxGgNMr8QazFbNtG19+eyHxVKSbBhstyqJ+g4DJLb/E8qqd4uoApwUciOqSG
56YVVGRecE5oFLCOXdvwCet7mo1RcWIynFM8LiJT9iS9lEGN257Qp0diBMmynyL9
K7Gy1J1MnkAODYG8F8fpoq4X7mn0NCuG5o+PgdGbc/nLC0pBhR7xXVR+tsTGN4mA
dmTixclarML7bHHEKx6nG2JtDhaRfr509VS46ESm2/B4Dk6aXhl5uCe2h8wjOrkf
pJ1RuOAkCFEKoq+vobRuVxkFwoq36/pKsVGINoHwplexSWYSRGZnqs+k2D+55mGX
0b7HvrgxXQ+ytafkx7IuGUQUb5BDvg9WffqAn1/QhUclqa8NEVpBVdC9s4IcNGLW
5K/LIY6/V+i5Z+Mr7vdp1+NEdtB1K+alXuTps/oMQ3A09ZA4fBL6Y9gvRnTsHvAd
1CzcVokZ8JXg7W8NjT+DShs7VTxNZ+ExvSYh07xghn8Nr1yJ+tsvPB4+PJsqjaBm
Slsus8E8cJRQ3c8eyIX2WcVDdn5wNXwuVAVJiCsjyCR9QkFgs71IZGo3mFwgww8A
PokPaJTzOyrOVxLu8Ihhpo+hTWGxCYDH18DCcNgjoDYCeSC+HMh48lsc0LpmFALX
QShjyElZUBnSUqLVeoTaR2qkCEYgNzjYXqCtcRmXnrFPRYP1swxr1Ade0W/SoZIC
Wa3RgYJHAN/tcKUIloDcDFiYXghv0VcMaAjKyoXMYMvyy4vFwwRSzfmI7JHIE5m3
dYG3UQ1Th8U6UO/ClwZAe3A6/nz9vf1l46Pi9X6LoCYRbg2OgCFnOQtpWNQXsja4
LFx2XxGg5HOqCrLCxgfXOueOHsKbazgXfGkKccPDFuynrarivbdU7cf+F0ShaHAJ
S8ve3/SPWDx42BB4n0fOwEQqSebWfuonzk4Oy8voxeTKJrLn09PnFApf8kCeRdUe
FH/GJkZe5jUv3kdsXRDUjstsS/5CEx3K+PZX4YTWlL54jNvESM79k6ENocBE4vWo
L3Nft43WqDuchgsFfHky5NkX4E58slky3wzj2N3zvoCTMr/4/0QjfHNbxq1YdFKj
Y4a/oEnr6i9Gv6TvtNAO66nhQLohhNK/ullAUPG6k1/fGJayomINOhcc2R4mnnyR
fvLghgtyyLtGtU9ypv2/fjzpLFNL7TbvROy+u8XxPOimgEPfVcNq/l6tAirmfsAB
9BGTlI+DceaqOx5fShKwG1iFxNbSxanifnrg92mhiQhwx5/bFpcOY1e9+vsfmvhV
TC4giNSfTaE99X0YxDdybqyS+5r8uQgBQ+86c7heDjeftkxmuKp9BT1jEGZv1viy
z+ChWOIxnAM2gu/KEQpe81YEDMdiB7JOD1u/dnJKvKi3htyZwd2/heHjX7829exx
B9dowLgwaCgVev8R9S8fjNeBEZZvWHz26vDDO1qF49GAujklUpfNRCrAnHZNGo6a
yXfp3tM29vpcPYUJ7NP70a/N33o1LwcrBXft+yzKLAiCelORVYV/EobRcjSZp3ZH
pon7FJVaFZLMPL4QggCLRlWyLYW+HT8fB3xfvEMAtnWyvTsw0psuoecIeTJXvJZ0
fVj4vSj/q4VNtMxCYzTPlBkqC0Q75vCXlOpLzMzomFSuYEKlranle/b4HOqwu/nU
jLvX++oj/N7qg7V7+eGSOs2/evPVQk/O7K3XFa8Ws+We5AWz9los0qzyyfXdkR72
xyGzIMIJhcyzM/T7EDMNWXRm45VCmwXvbf8nyWR3+KtrJaAbwd/fhhX/oJztAcSH
JNtKt0RY1o3zuCD/v9dqwbsP8c55zAapwWFqXGjX2LDcYIfy9uwBgL1meot0WcXX
DAoug5eAW5poaJ9K1L+YTKKWL67VLCVQTFpgQG1uUdU5O094Cmf+PwB/xjBCxUm3
+72rtClZheoSUdl9yrOxFc0Q08VvS3X/zmBMw3S2a1jjV16oZLmtOXMEuEfnAC2V
qXgoWM9AIHjhUsWOR8EvH9oZJ/3usOMSWbAw6ESvRYC1OGqdUEtLiluAMHeQLZgF
9eNBj17zAnVwB9iOF8lqjpBIpNCYniu47WeFAoehohvVlsQZTmlg4h5Bd5+FeYxv
AdJ0UnJI7NQsbtxQOYhEYLx9e4f8DKRYzrRxmnd9hU1a41GY9KQG7onzwLZkJgr/
AiGWZCboTtjxTWCqzXYhXh/pH/6ZawSiQ+g/LiQTIeSPHMV5aH7VxYB9ZHBKxjPW
C4t3RgvWBB+kCkWouJuzW+6x81SGPIV4F6/gjgSl+oc8sfFRpOQAW/wjG80kSJcm
9meLwoq0ciFjiDSfN7OAmQT63Zr+5IK2bgjIJzUlEi7VL1P6fJx1PQ7935YqrLgb
Sgc/EP6AM1Lo9KgpbjTAt0FSEGsH5lGm5EVnaPfCimm/vYdQC1b/wtDRW1AOrJAV
MepoYezbRUTxCV1RNfTZp/qReKpkT6Ffh4+yuWt8Q1egIokP/C/xU6k2aAVoRM2q
7jjT/1vy/2vQ9GHenACC/HIjegAVOXuYWiCsOGKIh1+S5MvFCsgVHnocp8cCIlF7
Ot8k8G3t9u1Kyp0ICVXOxCNafKDKDsy+/X1lISEEXlEcSp5SCnk6gXeewB9I1kPH
VHB5YxUKmvfeQbNjD5eKpGiol1Ix6vYbkrBGLMvlO9aoAfu51TEKryenSisTkJWN
31JvX8Vx5I2/OFAFgVHIcNuUcm4zbJ6ieSv6e3Cah1OfiFfAC75b/bdDiAjZNgDe
rlYtBHJaPjhpq0nL+InETNlUN58y+bhKsFuAherwIMKDBBm+XZtfmWpIhhFF7Yk0
8Re0oOcu76MHv/Y0tQimBBtGjK+cM842TbJOSKydpdmJ4DWv5KUPhc5SjAUUyzds
BHLhzR3xEMY2yJyq5g3CoMbRQgRiyTPUJ20PQlyFQi6twOsIZAg2P3L+5scsjwVG
Wrg794zKnYqdqF094Rw/Z6d0Ig9rB1JB/IRnysKjSVq1Ljfo9GL5LDVu28bE6Gxw
YlHC55N8NaNgd75frFezw7j5NaJB0nrjLwXy8+Nu728Foh2TAIVF1FJdMD05Gfkm
ScuRbsJYNkcVgCx6EkkY5aby/U/VGIozqH5slkh4Ikm+nT0ydsp6axdPpVmcUJlI
JdnILGL6/XVumL5VzMmFNLNwZzXtpexAowup4/73HUgGLNTgjEwsYC0HCTjHePbs
vH7CcRm9t58fo/mm1lmycyh50jjjXoK0RvLhT7iFPOAxeGAl9oaDNDdfDASTM+4K
lalS/gFghMjXXoTf9W0+50QZ2DnhbpGCXO9gN8y8U8px9UMKIaAaK8BuRvve2Bh7
sxDArrVrShJSmC4EjUFdGIkHvrgAMXlNNEsB54YhuCPnfqCH/Og1ZBM49ieqHjcf
B28YaPbeoFNJAHRt9cIQSjT8t296yCy0zEcOQ66vcJNRPGYw8sP3Gc9tRhNXHi+e
jA65XdRWlsCA0OwfbeKNn/yDV8LxfT3Uxn3X4313pXaKR7S6M1BIxhZ8NNEPTMih
cYON0dzFWu+g639kj8UcnR35CdbhOW2REtPEoP49dJV1Xfzb4TM1DuSyX0DVgmWD
cpoazgG/DpwWQM5ZIplEJ4EPXltXWtz8jye5KsSq4hYk2ti9BlAbWABVRWxpEhqz
DgunsBSswP7ULOupOXyg8xYfPVSIfGS470bqbWc+qoZR5MK9wYOl0odXL3dLbsSc
MDuywmoCn19CjJd88bPe9lz0j0xaVI3qTPCrh4Hte7uwEPS/MDhV+ERn4u5VRsNW
S60l0ePmQcE7mbqewi+QaDaslLXrsGASi9ke2dJEesi/qpbJMkWvG3EumAe9Izzd
qw+TQlYiDsv8DrEn/LHyhxE3SpJkAGsXyK33t4TOpY7dZiZb0enW1H5Z0dz4tUM8
hd6WhU/6TTCRqudlqULCE6qpwPZ3OydLpSXampxS/+HIgd9UzxoeJFHtrsiQc7e6
wVGU7eUPs8GgMw7O7QOlzbLdIjvywccvhJUw45xbRV1vZw4dNs7Zzkg+A9D/S6Sv
7wGWDnXHNIUXg4U2LKk3b9+hyy1a2dKa4g/nwG1Sh9E3HfabvqZ17FzzoJggHDwe
NNJuKFrFGpfCJBKJCv/kVDIgGhqgvsCsOvdp0QPHQ24OlUYY0g1PeI21NzWwV6X9
4Sdj2hddn8uP600+SRAY9uSS7YFVQ0g5D/uArbrt0itS2pnI+LtSpafW6V7PPqTP
SZ/oqt3U65DVCLL5b5ZaM3F2UsMK9rRSOv+aGoZZD/qRo+p95UVsLsvm4J9V1hcq
nNKJ2kpJ4EBf5b2h7cmwFneC5B44b0EK++dSANHoZughegJzQJjCjw13tP/3ulwL
UlnesArBdeEhjWa6I/sgvj6SP+A4Ef2MwyMUVt4Go3WbucDOnGMB84LuAJNqhV3J
D7wXf+5NZX1LbkkUU1TbWrAoDL96Z8kMs5usiAcsoZiORyYUQPhNrGAR50qcj8NK
mpi6zNk+2wvkZEniXuhT6e9ws3HW8Gx5WUrDFkrgWBWHu+RlCdA7VdNQ0ZBuKbc7
wBF9SU/7GqjY7M2GLxx/6h5peDIyRLwX6bHJbZhzQz9xyVRhA3e+64ZvQkuqPseY
cApZFppK1uELXBMRGH9Ll6DC5MHtelIkPsv23Mv10ivKqz2204kr1FW09lREozew
5UJmZf1HS6mQv2R+OH15FJhPofWn3fbi6tU6ecwaqXT2rRLLPyB8d2qlQpwEipx+
I52X2R/aOc2Rt/5UIqq+FDJ1bJ5vb7udZNf72yBcCk74fD1sJxIzgGa9EBXJhLrM
bVKcLz9jFITwcU7GYb5dEH1GHqUOzQSjbGhAUinIhAoZEhH9IibFq2iEXtjx8oY6
X+9ZSOQ+m0WJNOmfDh5vG528mrJC/eLf9UC7ESf2JEMcAAU+87i7bXHgO1pclpdz
HTq+gOV/DA0XHvzzzqwdn4HoqVKS8yf3jgEOaeIRTvPh6dExT1hs6I7YPlQ4Eaap
Iff6+3E6W82FxTIepJAyRrkplf6YCeiyfE/Pq2IM89xVzZuKCWUlK3PkYaFo80wB
1vpIPxqDWF5gIhX7I5MI4dAp0ROnSUNVYj/ExMB6XJpL4ChG9SV7WOIp23N/za/Q
atLAcdnHqV8ItUUmqgD3udwzq26uaSAF1PKoKjaNHyQrLrabYH3XCCHDYffjtUvh
Fmw5qg+0IeHuQ0NimWbOWIx2Llqvr+0fRpdjaZdlHx0eQkBkCPMKWULauxwR7ULp
HY7xUseuIy1mbfGeZjP1a/RMYG76a0u79OiNN/7Jt6Lm8+bmMBa8PbgZqAGISES4
dEumMaB9s1rbY8zyj8B6TgeyL0x3FM5TmF1tG2bOranmNj5luWFAuXqqGf9VG1cn
C6rD36ZbBwKVW/G640INU9zP43N2AsnTIqPQYhK1auB+beH8y2fPmFs1RyNQb6vu
KHHEaJpxJKJYP9RgskR4RXIaGsmUBnTL3C0XRRakG9p4vqeDxre/ZOi3crd5HEdW
hwJRDcoxrYwvavtmYfBg1WHm/QOWI3TYuMTusDTzreNevkMadlLe22hBACqf5zic
n2/OAX0LwivZ2EsrLNjRGhm88tOj4DNIaSL7ejcSQQ+3F6vbQ2LNwrvl4n4cpz6w
2zz3YhbwHF8QqEJvGHjNYFNKnxzyz3kCJ0GCQ2yCxiQzMxUcXCoAK9dl2HKz5Ioy
JQagbCmupP3OXzn9zPpcby6QA17UuivyFGbZe3d6DRRLAt2s41VpSUBYTp6XZdww
HaQlfNwrR3UnJoi7DVAuqQzvb8Q5a7Ie9xNkmYe0TAyNlGy3auPjWN+lLPJKvRkb
0eNyALx1/i0P7ozt5R5I0VHcJRXs9smwiZB6AifEjFfdlMo23gvwFlNLNxEeEslE
k/8LMngOK2+tLfoPfEryY7fGh8enCD0gQVqcZY00sbF2xWCMikgCjcmb39cqt0F+
1vbXLdllw9JZqAKRs7eD43g3J2+UIuOpTYMZcxmCLUKrKZTnCMZ9/0JhWo8oDKNF
OjOQIpqQoHMEPDC77eFUGhmWsWF9muCja1BqLgT/FaLcL3srwTZn8YWp28WdAD66
EpB9ruxBG1dAyo6OQiIXPbzJeZuEXty05yskYGPTsjvv+CmM6vK6psm44FvH7wWQ
vfUxZow0E+fbQNcm5FUF7d+N4vlk/tdt5JZcvMdvVOe9FVeUcXrKvDI1xgRQzcAA
xryeBCFbo8xfz9Uua9oQp5GDLXEHcmsp9zU+yyp7yKaUb6RnHgCV3+OsSfQklUR6
tG2p5NPFLZ+ctgfECiI5Ehamg+LAC6dwleE+9SPU85EJZKevSNJ0CkDB5zXkPMYf
v6i3Uft5ww1ghnID0qnme+aYq3StyJbA+xb4L4oi3JcMrfeckdJq+hHE1CU4JdYy
JH6KklG/tUE9fHJ8bc5w2wQLkdgR/e051J5XAQVj+RiWb3Vl8ddDjTTj1DqsqCQR
UvZIPx5PQw8uaSutIbinKucfCNZBleJXlmPc8ZNM/G9OSw089tkTedc/CdoXX9g/
bxjxUyW4dWpkAx+GhHfq1FimyIJ0Wr7QJyJ2ajZvfGastP1mLeDapVBp07+x5/xI
+ER36s/PrJFizA6+mjm74PRM+2+uA4tiNPXvYmfHIsu54ziSKO4mO9d+FMVSodMT
DSFlo1Qig6fjsgVQCCc5MTHplP7zLzYR/2YPQhkEUaRfKhAKIuJO42xlCisI7JOh
TBLPO65Exy+iuplJvtnU26M3SccDKcll/Pjco+nS/jrO0mr5bYatO/m7s+4EOYm7
xABzlLbSE7ouRDBNt1B+vKYFPzGVgpLS95TajU/h4fieXkflllauOHzcbhFOpaZP
66mE7s205C8ndcPDBT58nQkBseMr6UBT31NEG+P0aCvMUqmXx/0EnwOQ5FjQmsNG
muGROPMLU7J9wRYBOEjCQtGCG7mcQI0Q9oiENRJ+e4vTkg22x96rCNE3ihrAhCsX
qyv71wgFrOuTGLJGJRHH6KU4ljnNJ5y/HfaqOgtIChm1aIwYwh94XLz0/zK1Vh2h
E+fXroFWCgftf3e0Yn1IbXRWucDaPfr+OxJo9H/td3eTf0cxq/onIEjePw4SPVZP
zigm6SkQez0uxt0/lCEodUfviKE0humm5eGw5Aya2uyY/kQIDEKzyAVviZOm2RCh
hQZmbMuxhHmGEmFHJ0cO5rVsND6jE9nmMnclQflxe8vnoNgNSywXfUD8hoeajWzu
XJ+nCSE2H173kX7M1ZDBe+d4pOGI41EBHzOo+EMA6c0fpgkUSBw1LVLaMYnwUqyG
wEUaSxgjSHoG60M/Xp8oxKPWIT9ekCb+QjysYKyIpkgsdcjciLbrgu3NRvIyYlw0
TlChsad141hH6q/7Hc6gyHOz/KpGkr8jx//GHIA4sQ+9dPq5FM/BJe2+a9fQrdUL
35sd6lmX124wOUVGYUihq8OkPx+/3Fh8PKGKqaMxW7q/0CntMi/X3anED1TNwRHm
9tx6pRj6VzfPJT0KMNGEe99Yn3eX872ayROlls5IJmDT5FUZ7uQ5l/cI7oSAxURf
fas8d20q+Kv0wJ8Yu5L1Al8Ec514HAgsjolFxTu1DEXZ+Jh/ww//GOLKSUmAaQ4I
ulX6JEpcZMK94mxJ3FgpSbbhpGprTMtd7f8vHo6ONjNGQoFLX8nt+ktLaKPsEKPD
LvEvZFfcad3MLyEAcas4cNhEd8aiu1pWeIw2EZzl+h8vK/wbpBFeKc/t0YSTZEXc
QclENyS2MbopK/yvnXyP4o1pQyTxWQatUGN6u06OJnZp9MgQAXUigALhinJZOb7R
ZcV+QlISY8B6qd1WCWnJqfVjLu+GeEhcoUqOouqSsXkqOiA0CrBrWmbWd8afbi8O
kNMOwKGE533ILn+B8Vz7qHEa7TDWXTqBxjXTzrjEdXOj3nfBhARZlTkYGI6ggA+M
O3akdY1JaJP2N2NnET8M043AyFMiWpJTnvMowU99uaOapEVG1yJcKJzUj4GTncdb
VP/AItvb9yYuctY8NOeuHXuGeNj3cNjiykHLaAEGcVgK7Sz1HwuWuyL9CMKDonON
k4NFrW0U25C9/AFaEbRYR7gRNNbNPnFjziy/T05Dyt7MAWxqfu1ywJN9DuATJDfS
GGS0crIzSUzi2sErowLdynU6Vcif231zLMG3XEjQ//aqWfnT83v4laiEJ+fNff40
T+2HTFIloVbN4gyPXLkeJm9QJH0xHyTXi41nNm2xmM4GB9DMd61YeamJpGlAXDG/
RpiIEE6B48hrhf6iy/OQE+X8RVeC5P1xpXwqYL8UnVr5tQMwSjfAG9cXkaeeUQOI
mzgan5Pts8Vt+h6XFUQw0CrzRIrFhZEYrE+UODB/UTELbR7rffYuihb8ZDhmwMNO
bEcjGGN81sT8WJpEwvWSD1ZemecxW6A2iqsn67u/S5Fm4DycSSLqyKUrPrzd9Vos
2WAzWZRvkpdP+FtKt+04yML3wduF/xVY7eN8KGquTc4i3s5pgwiuc8T06TGBC65Z
tC+GL7YNJDuITu+JNSZpsRrtySZwe/SnTfLUyTE6cPDsCHEakZsQ4i7Y3Gh5s+rx
MNroqcGl6QgfCjm/x7vm2PdoFXw9nUAyYjYR9bHqLURReuf7PiChHFgskcNWdwZu
Bbrs9tu90/3LlxH4d6Zxixzzt03iy+soyoTGw5pPq+2pjF9o4I9yoFq2BjMnez/r
evTvy7LSwVpVOkiENhRjKxlOBofRfsr6KpMOT7y/Ww5T0L2TO9pXBRl08Lzvm2fr
7e99CAcL1459lzO1TYcRhCc8WnfSsh61cKpYqlYxQCm603QyTjXKdYvUKIRAsegx
2H2GOAPwC+TG1FjqMX3IoF+LeY9aHxg6b7gDR1Vh/NrF9BJdRlBBjRPo6i7JlVLh
p0exEZUJ6XoNewaL8pl4QvdGD5l1skiBOafwDvMkp4ujfYlTp4PwjoXXe49xd1B4
9sp4WPOytE0MpXHCU4XJpUDXRK8VimxssyvRyN9pVMjApt+fZqQW07BU13AjGlJD
XG92ZtRpoqFf8f9wI0Yc+i5oYZprZUEL9kApJ79ObqQIGEeh38zv5Dh5ZBtMTkb5
L/aEHGHkJUF6EOtlMsvUNFsFbhVdV8MZYr5rbWcb7hbJlNgexnlkuzqL9vtoK4Ng
isoeZF/9lbuMBNtJezmr4qrJ2+BNgO9D2ZC+wInAXtcP2uVn7BFyX6Y4QjstUJNj
hZotIqGpJ5yCSKZrOmBL+iicpExJXzvQWpn5nDcLflFzEEsp1oGlS9YA+XgksIQf
cS9cm306EqUojKo9MBBOpEKcrYJcOCNfmR0RKSmlGrluluhER+h437m97lTxGVvv
aq9N37u2a84ExI+E8tvKa5KKWp5WFFdc6bF5FzJwhermThlwQiNBBMG5YxLf2OfG
iszjrtgvuioSxUDYqHmjwrpr19lh4F+BTU6Lc+Id5OQut/yTULVVRpEzrrWPrGSg
/lBtxtBi2Zb1FCwyBbQXusw/vzQBVh39MdTKRHcsN5yUEbePtaONzZlICZ0lB1Ew
CZOgRW6qNdRXeAVEZxaPSG4CoK4kPqu5yTz9h8G5YUNrTCS1BpkLfamTuohA4v/E
rCmXDnYjN8Tj9fVUOwQmD3V2UeDCl2hUAYLlDZrjZeh3xozKdDxsBRu/dx0vy86B
FjGQeliVwFFUZMadn86qCvDUxAkzKgyazW0Byai6eUMYrtWlAOc19EgtqKau7NvC
t7TFKORfN8m1+8UoBboS5zHKCF9rIk2Sa7k1M5royxCHXQIJnDqltUUir6LXx/cE
X4s/RAdchoIv2GoCNsislV9jpFWMLyt+Rm2Lp5Q7hcUzT5QM+Rhr1bzmUI6TE86g
YpWC3cHrCnJIgOmZNH7iFe1LhX05pHrVSwy/s6cwo38UNz/kYHShgzgS34E9bS4v
0U3jyDiCwghD3O1kow6YUHsGEkwHPwsrCDUqN62lk9RAoor9v4dy410jJnNukGS6
GueM46c/INo69u1yLwX5MwMfBoz4PhbiSxmkKCu3qASCfHCGaIcEvBifus8eZF9i
uhExXT9UIYlBnmMYBieXZFwQVbKTTWyfzqesawIbV8RdtvMaUMoO3ptkowPQDscA
qfnLNcA3AWhC6oaGXrZCAU3wH+hP+60PCvJxdej8ZpPc4fQCPKngkydyKBvgnFwF
aWVxdpV5et264n6M1eMUx25ooHvthicZdp6iAPjcwVrW/RIRNKHWvApwj1mt8Tok
cQ0RV7nTYnDfrobgrMREXkYt2tt50EDY2ByKo2XqLYctv1/ZgqZfSCbI15Kk9zVE
OamLPRTMq7YURgd7Bq4xTNX7Du4Hq+cc5T9rRbSxCgmOM02EqVYjnJ1jwF6bJ0cf
qRAA72eJXSWgv7eFBW/v5uco7Lyum9uCAZld5n1ALcUKbTn5GetsYT/LfOnh2WsY
0GHkVf6n0i3RqY+gYXGvumzVG37JEKTMkE640ePjSnKHLqg2NP3w9zdqBXju3yP3
vEkDzi9Lm4iFx0GPU7oiCdBGuCGVrzWIxvzpgYEj/9wOjZ4ije7hzV2rUqdjVbiR
uCgUUYORUslaG9ujikP38Ws0yMpKAvXUgAYDOxl6pUKmDbXFCxDqlXvwcLYNMavA
eMUjaQ9rbwHOVh1KZgEGXARl97Y80ASAAyM9+tphzsuruJfeWXfcD9XexA+Hn6Dd
yTM61gFAnbCJyLAW1Q1vXpVgZBtmPeRq+nEuna6xKvKt7Qn/t9u9ColzY3llsaR+
kZzj2zykBOj4sbm10w5fBb543Ga3LVArRFONQmzinqKBQ/pI4TJUir00zyDaH6Mw
86tn0/63pIzHeWt1ITUjcTmItrjqhmwLG/MHIXp4uUrbq7p0jTtGUvdlykuBCE6h
HB0u32aQLwbFO4UaH03UaxwdWLjw91hc+hanuOLYI+DNgPCuMsP+UmZIDgxdAM47
qjbLOjzyTJh+95jOdripym5zQqpkcmK/ksTG6NClTkQn50zAd/9PM8ppRBirD7Xi
Y6QIG+sYN+UjedN1ND9QZB18XLEfhsurLBkgpKINf/hipQTAuY+7s6/+VW/Buuy1
j2pSmMF/Sa2feUXCDcoUX2HrZ4bSDw7RjUujqzYnMgXyoOfR3yRIUoMa4+2H+EvJ
Iq1MayWKZbXihcgybdaig4nuwbndmzVMcvi2sM1Zs2ly34iShkbJ4UCtCWEYA2Nk
GohAlPmyZOHNAdqg8ijeykiJ3Vb3GoCgSOe8rMeOaMBLa4djU8gMqDU4jJo+yNN9
g3HVrolQmJYrBYbJt7gL2htVUmMd+ym6cr6OVNn72rtSbt5lUfqy5unnUZFRVWJa
3czCsTWyMcLvHpxDs/s6juOXK2qf+WUq4cL+03b3QHoNICBXEKe16nEsa+UTh7fG
TsT30x1IKU7fVtUh5e0o70Ie8+WRDCwKq7hH2XsAeuAv5VVRF93vP02PBHvIKEdM
J3MLaO/pNL6IBWLW96/kvTSJ7kyeViPY5JgWYpiqwkGo1iuipn7Q7SnrQ9nHn4tl
WnNi7cQvEO8ym2gmW8bWlbjpmlJidQWUA7xQeaS3SXYMstea9k94+9+97K9zxnuu
8LmhP97IhrceRx9WBY87t/uIryrIfGhX+aZdFXbnLW7QDRI3wldq1YF+iD4JHEc+
ndhKdUN6HEHHxbRqbnhmInnZH53ZuQMqnC6mHgd0vGxrILnJCWRhbHd0qFh+7B4j
sXlxOKbHNEX0oisAT2d5nP8TqM1EtB3eJeTLhA7pvmMxbzvclAZDpaGWNmRrkSbg
kGR6dl84OelIYTbXjkvKRTrzoqQSFQwdAo5LeFuM3DRBxXG/x/sb1fBjtCRYDgfn
6XgWzkiRUeM5YIUYYpsca9ViNWY45YEpScChuVhfRXqUavNJSGt/nRqxhWJydGPO
Z21ezVLKMUGJDo12pEazYjlHgGkw2uiiPO0yREIKV+IFHJ7wP0gbnBTCazZXRMLO
MoQ2i69ELf/lLtDwUjlMmM7+DRDY2xeuXQ5ROmjPejy7VrUQCaHMyjkBM8xw+Dum
2jUzboxn+yknqsIlfqUUPDV+8Ptb43OfRd4J53iGggidLbLTm6pbAPLW35WicF0C
w62pHDkUagGvN9B/zcEna7aDITPPzAWNTIOAdyIbiebL6SWgG/Jz9ogbaquuOHEa
oh4tJ1zXxyLpexYqglvpXUOT2dM2/VAMKj1RO+oBtot8IcJx/aD7UzKmvuyQHgWM
pR2MLDZEmsgsVMxra/HTBoOlBMN7hzfLVYFvuEmrQ+bIpY7V9KeDEU7XR7q8y4Hn
644ASmbuX2VhNDbPafrCu6Za+Tw2k5HZfrA0Xfk3VpaMFgXzxWw10cRAnvqb5Et6
AV4qFv15ZHMVAsMmb019MVxTBiESCwXUqZMt2EWDZi+JJymx48c2Y0lAzE88xHFd
TMERryF0WziJ0GuNcIVSZVBLGt5g3WUMkpZg1WxtRzrDo4dOate9SLDGpUKkNgG/
myT2bppa0uqtESbFWZYeCsKjb0sExkhwJT15LOtxeWgfSlhIjsOd1L5cgTp7saBt
q15nUqUnxycxuDB1PyV1pMuy5+eP2LE4bk4j4sQ8WSOof9D2so/GynIadCfnk3EB
zkh5Q2hlDUvAauFIkadK93YvE/+UEZV2Azx4E0t3b6BPdr99dsGVPcp1a6FkvAYC
TK757YRN42iaZMXulsUascnt7dWZpUqXzG2QoQ8iloGtGm3RC4TiFYgmWkvJsswj
BlNqSfF1qnJLG9DOTewUqnLxQv8eenRhQs8hLydqhn06g+mzm7W56JUGHDXvsGmS
uSnGfcj9/nCpeC4FA4DgauoT4hodUdMBUtAFYiDusLizICwETf9YdFo745WfEKAT
/uz3AMgjGtDhpzNzuM9C44KscLANfufq95PmlRMtXJn+adPqG46wAyamb632tvci
XXwqFqr5kxxc0lq2w3t1uDGupOr1abrxwCLdYdELv6cvBXmLzlMzytNSY5jxc8Ax
9SgFULHHeVD9CDSmQ3TyoAkj+eAd0+u+jmL/MmQj1h3sMgF8+CGSQX1WEM+DbvHq
z9EiH3na1yYxT2sBjhldqGLoi5SUDUFJYdSL/lMEvU7KZNUEAROhwuF5PyWoaemo
FOUP3Yuc53KCy0u6HySimJJR4QbVsry5oYwI2rAB7gT1pZ0vvj3fNhfzLDIy4nL7
sTKKhbCbZlYHCw/Pi1nxr0iHp9WwaK+urnTeK82RlKqjacy19Xz2ymqBbZNRdUBj
SjJx6I3CqxaLpKEmQj7zeKOg31LCgEawhq1vVlUtZCuFOvQdaCgtgt55kn1kmj7t
b1rwiSZAb8AwiAXnKw51IyWEUf5Aj92DC6W/PGjKtMr/BW5uWPmwVhkbrVCwiSGg
8jK9svWH/S3TIr4fgjdPcfBaQSdPBShvya12OouAgoDcgQe37b99xFTHLe928oOs
Jv/NZ9LKPnxBj6N9fyFcJxM6HStXp7104vQiGTYbyPyhRNC9+ccaQSMQ/B8/ZObJ
JT0lyViqbs6Ycp5dNNPukGerfjTzy/vmkK0mcMunVvaaiSCfD7b9zOKxoV9wNP4n
F5IEQSytq6tYA6jtpYg2Q4LF0Cnisu0k6qy82k8NHEiMB1gLKEyxF79IRkLw90Cl
5kE9qQLyAQVlJLkSb2YnTy5mCaPDZw02LSxfZY5C44CoXZPbOxJ0e+aeKwpf1OEE
NLAl6LLC5HF9ZgavNmuXHBIydYPhnNY7IZLNPggcmWfg3oFMVbqwiZWPTSSts2o+
YGVyoL1JSrXhxDZ8g6BvF6jUTH0tmsSDV0X9tok7dDjiK47Zvmrmi4fLTShi9Fx8
WX1KtWwd2KS+AWcKSFlI7WkGmfMDtN9RoEMsNcMbt3MDqY1nRdv9NamlK8H065BE
lJGTFC8LJzD0xdPE2UM0DH/7Ag4xe0srfbuxkF9oBMBWtptxiaEiVWF0+n9jIZKC
Eo0VdDZ7enSVNs7NIrN1kRFhfQyT3T75ZdRfoQe3VijffkM2VyQ3gnCov4/7Wlh0
EcQ40t483R3mg12a8XZN2QO2es/kkvNAnACZUkFlBp4+w3B88UsUPTK3yytlpM8S
LayxBiix7ysyzggjHWiFtSDcLaCGZcWfr0w86VVTVGIMOWWgz9ZTzGefuMEb3HZj
rVvozuEKi4yIFaItMAfYkHeGtdjsxFwy3pu+3Ig9kUS8HO1tnEOR/VYUj6k6S13e
bRFrKofHrtdx/SUXbNz1esq2uDEjivt+yzkzTSaiUmA+LOs+6Le1Rs2W942hOYPn
4pue/Rn0SJsRfXnwNFrDkwwvB7BgsO19qr+hWNaueWWCWkUXvg9LpZdlO+ea9/bG
ZvrwggzY9OjYGabI0vEzHQHNVEksAYWL5DR1KCuLOOYUDbLmXiyVyEnDkPaK8zy8
exjqOBdyUdIIhyX84MgTDlA9KyjLFeHm+cDGi2gmljj/oNmbnkmbvAVHJlumOiYW
jwacjCjI5xxpIj0He0LwFnaqBL7x9UnalycmesVHZtlL+3uOZw1XEFOtcbSPzj1n
Fm1uBlHlIldQpyiTwsZIMbpxKDTPB4Q9U1r9PUsLY0x8URQXv4TvcZwJtwTZOqKW
4t16UulD0smPOuD+cVb46OPepUy2FFroq0LFGiJa3AKSrROVEdernpkM3VielMU0
5TvfKoGPj4H7sQmQqtXNZQy1Tsluw0opy2WRDHYi92B4yE3GEonnHWbtADqEFJsf
UAH6hevIsbz1gi4yMe1PAPbM62exh5tTrSN7mrW7eL3WL+UbJ+4GGwU3tWL7IyXQ
+0AL7UIELQc75PaV7f9iLHcWkgRdL/bFIlxgQP0cErx/oV11I1unCxwbNOj6kweM
MksFbBeYisvWM+v5xiUhTVcEbNKv7I10jRAofd8GYmmKNm4MnOTJ8uCc1HBlFSuK
JS2QbJ5RRY673eWbn6JL9Q+J2Xl4R0zOWr/GqMDBbqBCx8s+fe5nn7hqAwhviDMI
VsmWUsoh2VogP85+BeujwsNas+mPSuwr2ShPANvfPRbWESzAEQ3mW7Yuyx4JVva5
ou9+U2nwR8lYu3TxlOUinBWg5DMoj7EJnIKfR0seTD73TfLdjOWCn4SNnbo/grZI
z1uFCkmk8F9y0rLIz5Pkn5xvhKH4iUX3iIMtFtQBhMk6X4lBRYQFMCPlpA02xmwj
VpudN15tn6KfARzlsBeSHbzcWhxHm2xjofVYr5hxan5T7s8uD7UevH3oGBQS4PTA
Pv55nl7In0K2z6f8Mx9iPOmxV9f+k40IbDri/2R152wZ21wo48+ZHJAAu6n/p/yd
m5B/HLFuKl4HlP6O4gFzVgfX3IA00Wt/VTGOgFp6FjHy9wg3gAr+Cp0jvioHk3cv
05PUnjEngOcFiPQ0AVQ2ahs+gYgeM3VrAbk1sbYyMQ1fywXtLDQRaEodWpGnGXkU
h3Hm6mlbnUw7/BXu8iIAnQuMs2XnoMRJJv3mZrS7pLo9oOx0I3W+X1O6sZarrdOO
Pq6+bbe7rglTV2I1/ud+vRfIrdea837AhmVNI2K34OaxPdRtkiLiOH9SRM2BtSjl
IRODPHx6IhYfhWUh6D7lUmkOCL664lhYRssw88rqDtfPrTFCoklXeRV2N+ze+4AX
0fADg+/bdC28vDson5rJOUU0jIqTAUhkLRYwJ214e5aZ2S6WriGbkwJ0JBCLmcxP
q1tZxH4zzN4YaNTjR1imCikI1oE7NX8qk+VKmbMWq+burwjtCQ9le2syKi4vl7p4
JHOztAaWPF2oJVz3IjiNjzXaBVc7FhBfSt4ZxRXHOiSrYwjMXatTK0yBxhYcfp04
FEqwHrQVwZZU8ZMDyUCCJ6SLhi8qKuxTTAWNOZMbwqfgvS6Z32w7P8fJoi34c088
Rj89D46+vlXSdUHo4kxz5ybcGo+/IRnlCdhHSO4wEFrHy2AS2N7EKBfEi5JI/nbQ
Xinb8xNbWpfx3tmv0kJQgtkUf3rNLwEgv3WFEW6CnPekhfaXjcHZTOyyQ3iFDflI
sUtC7XsMRY1+Dy7TW8tFm8GQUbfOZAmhoVktMZ9RSMygkUpJVkxRmwgTpFJaoaGR
GN5s9xwOsnzpzbFYJcDuBG30DVrnyxKIYFxdK0kRvgpe1r3dyDPqON4881BHTesM
jiz0Lb82YU48VLimkaw1hAWzu14Ms8U0fYw9uLh2cIyBLfSszncJIW8a2umkDd7i
2ZjKkDQt2wtp2d4JrkaBPlikNBG9Zdjuk72FtYTO1cqqev4EY9B4OZUPOYDZjkul
QQoOEt8UJSAYGm37fIWtdP5HLZiP0lcnkN7/uaFLBAHLqKKpX6VG8poueg4qWEMP
+9/FATpPCAlM0UhvCX8zm/xIIPMGh6JX3AMcbjk7e/ZruWONKDDHo4XXO2WJ2lh3
5ZWjGwiYXvoefZaCg11UNgl7LKU5Yjzy2710pBzL8e7ZpbEJ18WBZ3JIbXhAE3Ju
OXCzXaKmBSQP27+quNewkYmL42mmgecdMsLN6VHTXJy05KEVEx3CjI08JOMRcZmZ
Js+OPt5fCPfgUljyPSlLzh0g63qSz3hsDeDiUgsyAyUlcBi5KMsVXISlvuAQynm+
faw4ureJntK+1jrjICjbdLgBhNZYV1DjOFHsCMi9GZjS0Hh1CgkOlllfbPPR58VC
IeZNwW0PHMD9L+n1JmDFYH4n0tQotEYiWbMrR5/ffX3D75H9qYzPKtN7LUSFt8V3
WEdO9WrEHsFkt/vVaSNKrc5c5iq4AeMBAvd1syjLRTFI/8m1fNlNQDRxJxwu2wpK
ReSp705v8oe37Xx9xXR4iboXpsXMAPMKfc5eNCAjOJIU/5x/AagtZY6P4ejBtW32
W+k4OnEcxxwKz9Ah9W1p7WaHER2nd+vADQjv1oDVGWi10yt/Bn+NBIzmN/fbIXCk
piVdPsX4lBxIRZ8YV6fa9uN8PMNw2J8KQEJlT607hYriYNwcOJjKAgakaXrdEjIX
9ytXuo7HivhqXTpi5FtNrUqB7B8zEP/rsImp5SyF6jmrg4Q2vspNq2/qSATqlXAC
u7jHaHWNNb3OXE8SApQFnZ/HNuB5uauSnwxwNNxcyn724gFCvesQGL1GOfJRCIe4
48kwqQ1jg89x9q7btGNE7VDiR0oS3tk3HCrmtL8eoxmjEnVYyZAopmtFgk6rIy9/
YMexBzWP0Nlio7yNpkI4Au0dnvI8AwvPdX8v5oz0W2UNef0ZmpiSPUp4CFipt4Ol
jkSJl31kmKnPcPDJSDGfhUFcXkTDWT5UjfGFvRlNm0kQ5gAD296xt5xr1I2XgsgV
Zf2FZ4Cx/8SH+TOfux8SfP6nrxL3WSOyxjunw/FJBfjX+59PuSpAP8GE+IEI14As
V5q+PuVvJxKvzxTzWnQ28Lwp+9OfUjTa9kOLQOHGWbIlPndZClB5uweNlNcAzl2/
ieZ8DKJW3SMxq2H9kO0/2DLJdt8gEqpETGuHaULP1/+2MPcfTPEeH0cl113XFs5s
to7DH+OvfO65h7fm7vGDjnFeQPbq5BTyXTAFkSSPvIN53sBPw2abKbBuzevZy2CQ
BB60EO84qNQ1u7OcQCvtkCYsUehm+vXUYX7Kf0wyY40toTmt+W2WeVNQY5w9LoYi
06VANwFRaXRkaiswqqS8nMnULm/wadk7STOfrTn3oEdD2D6sF/TW5cihyPgV4Pw4
raRz3XZvCJbJNVsOA6NKmhEWxMbACv0OXYwAHDAYdTWkoE8vVAy34Xqopr5Rpivh
LFuz9KtLcQ00Y30dwvkjXPMq+B8qrPXlbkz7z8cYz1WAjtccIz0zaIjbbNASAuiS
T/IRgg3WCZ3oFMDnQdbHR7Sh/28UlhQxdC1OxajUO4FqsWUv8suMJYL5jLCK2pqz
UITN+P9UPUhkx+T8+FiIcq7UCdSfbZd6Vxejq1KWmIsn+QOjMKbYgmknlbiIbCBE
qN6Jj4qBPP5+S3mebgteOCc3qnjWYIyhKrkQQ6kpbBt5RkUC8WDXNaypXwLxmX6S
7y4ZHanLftT3D0vOv0m6uhTNMHkfLXI3i4FJt39Rk48zJEvnmolW4PeqelEImzeZ
3IHFmig2+mUgbe25tGqe8Zh97CouCL4almta4JPG4OFX0o5g2lNFFkLKKCisp87M
WrHHRHklYB+k7oLeKekMIiqThZY2xVaQnfS8LCe93I8SbZ8g6Yn2nuMXWN9sSsE7
lEi9NtANmRq2x1kNI/MmKSRCzTevqI7VgArYk3YeBFZPjZxfj47MoLxQ5NYmMI2T
BzNQpr1c+erc9p8iXIDsmVlzvL4AHBTqPuQVQ4jjxxYCQqqEHSIB0oZlpPLadZnp
ML0cI3iq4kReNxPa1hbCdZEaL3q+1Kea1gPFU19DW/uJZdku6t/tbr9FeQLJfuV0
1eQpMVECzzvXnGkZ7ZDgv59Ddm+Lg4IJqVzQQNnlsBKmecxR4QeHffn+A6PAjPGt
dsRWwA9pwqsHPj0Eaia93vi48x4buoms8dEyG6BqHgxKGVuEnvO5us30n2fLz1Jc
AqQ5NP/C84I8B+t4TjDdwAY8zddbrNwoo9hMQkpLDK2rch4/2FOAomAwNutvsnZ8
nZ72eFN1FiQ9wiFrLLXNl6w4dpfJ/NwMSZlJdpj2i0ErXqySckhNhQi9n0cnb6s+
9LPDSRQRWC7CHN1pIOgfK1xtSjxFqAbtko/tiVYDQOvIk/jP6IXml11EhM2krDZV
MkXDQE4YwiGNI/WuXDbeo12DUMU6/oUNbEmrIQQezdKK4xE7TkVTA6imDztmpdtS
FsBgsrcUMOdU0+RlRNvfaD3vamFTjY24SKCfADSqyGoEFSD17TVHd/TZxPCUOJAk
WCUNFk0+sKqeLTwUXPsRaxAC630rErPzawve+MOVdpuBlTcVUk3JxG3NLnJWpEPU
9PmEh1CPZaIf5vA+moYwpXBJB2U42xBJh8Rydd+dlX/PgRTXOrex5e3/xzYeBl2C
SgJmi8UEGKjviEQru6kZxbL0r/fW3HAhCaAXrOX+QCJ3kXKphbsi6Y0CSlowic3h
XgDDYQ/d8nPbhgLGhPT/2Rk+te2cp6tcdyGjPAsaodLhp8Zkcoy+Nvuv07O5j6Yz
Ter3pfAo+zlj5QTXoYvxUy+wOoxRmZm2jhm3BJqWH87atAiGRGguR6CfKEmwA9BX
yrgrsEswm38amGcUGkL2tBqIFOQxJ+ScXf4STUKFSjCj1QtScuPUGqKNvXSEwHtW
TIXid5DULiV7LbwIT/mzGvZrm9C/XMsN9/zJehStFHIuxBVF03h2OuGlSzQSJdkg
u0akVuMVyfWzLTj/zJDCbm1JqKy0znQW8EWW0P5X8xhLISchnMOYYjsPD9TsHRXn
j2CviiRUsfydkIvKwX73rROtgE8kaAm2DSL1sHHnAehOt7yMdZtbj5hTzurBjNLZ
cVsKPKAXSjVwJaKcAPxKkiBXVxnycYxHDgDtx++Dcu6Sw3TfrgNKKdCU/rhYD7M1
SaUp0OJ9A96TQ4s2pGfqfJgcfgoOAKxEPF6rgyPZc2CKpUeuaeA9RZIX9/ORF8Od
edxZe8M3RCHIYQuulMmpQnvAvrkHvFLROR9mG3KHi0KGNyIaAC9Y1CAK66XLXeVv
IuImjW/ip+CtgTwIVTrwgV9d8IvH0v3icLi+rT2LYLWFoUssqjjs0kMRfo+kPK8f
NjwTKsyeHhioKamK/eOJheqSc9iTlAEXoWLVdPq0j9WdlmGo/EayyVVYttAo5O3t
tffaH0MVYbGYh/qL5OPGzyCo/RM0+cO7oNt3PMFNAJ1sPuCcHhZljWT4QDYFbSsi
Jw3mnWHbMA0tpIs/5EPRBjHlWenwxZ7AL/ojeT45vIuqoRpg1AMT+b9UMFyqgBKl
EAh46CYUybhXj/tBUljvJS84DE2I0VK8GnUiTINWzbIXq3ET7Yi9cXqWRYV1NMUW
XAbklBKx560YrbWAuVwuCFdGNqzMFEfqtuyvvmIpd45+TbPOl/E1ZlaNytNPu+Bk
pp0eeszRCvsnLZKIFsFFT4S5OUwnw9DuVSlVT/YOPqIJl5gI9FyRA7ByENFR37dQ
sVtCrXwlfv1O1LPTf5RMqH5jVHv49m67Px9zN3I2jXo+qV+IzpnGkotXEYctmHSX
7PP05c/rn1acoOvphtO44U264qFOEHJWJ6rs2XYBpVn5Y0t0tzDFnwGgYXVbg6UY
x85dNLeOvjcHeCgS1BlpIkzx5JgYjPvCdMv+oIHbYcPfJonMWMsil+0sevGp/rJy
oKMoXNrY44/z/k2PIphqJcvn5kQtzNxpYXakmeLJdym/DS7n0AIUOZRq8dYSo+3U
t1/7ne785OJ/3lD7Yp9JY02tCffI+AqYM7RgEMX1HM5uHUAn2tEsGiheQWYhI0Vi
VJ5nencVZ8b5vJntHA6v+ny0sTiTgYbO6EK99oei+NImVU8RTdeQNsd8Yad8+9DB
9zxHdgInF7t78tIGiK6tW4s6p9BTz7TpKI7N6i0LQdHvcveYfQtvpXbxhgOUL0rJ
0Oup0dy03DdLaEsxyr2r1TuFjIEM9nF4ex/M/TDXXfY6lGrRo30ESWKxLtDfLpqk
ucxG8j3bmKtm0c/BYBPITR+q3od21n2CES0zCDHqwhNoGA40w2xHM+rp9Uv+2iWL
CnR35UR3DtMKTTheO6bSUGSGq+HNl4dI+ibAEg709u8f1gAQ39tDkGJZXiczkMc4
IX1J+3tsJvo3MmKbreYxs1kA4u3THAtk1kITFUvK6LZWQsv3uXQE4vX8D2uz9MlD
o/cVlGxXrRE+3Z3kOXuj3Ear4JcX4j7S+6kTUU2/mnng+bH9ebvkCzqVqu9FemXj
REdpd7XHyZq9NsIEleD2Rk23qB1OAv88bzvipSl06EELcpkNMDZ4EgbtVy3w8tqx
47Oh7C3Avllab1v1NxPIbP2ArKmDEPqifKU8J8g7Zm1shqXTI3dmUk2p4DnWnGg2
eyTFG264zVtwuEsney5/pK8Mm2CuApKuhxZsGCI+vMNk0nFBe5vqNBSEJ1m4SSRM
+T0eeIA0VlgXDqJUdbcqaq7FRHcB454ktSOEdCp23+9OOGc+BByZ/AcbnazrCWbl
IVBjzadj84+OIArdhiGhGSWHcrhBMmhx2FKYz5+CqQQX0ZpzFs1mefN/u7W+59k2
TnoXxrz+xAGv8PA3N8o7zA2cfflo/72kt7Sg4mGlk/Rk8gLJrV57ZoSL6QWMEzcw
u2wVzvnXWS6YJvO22BwX5lG5t3XqmCs6jDAWpWHP5F9armgYLCj7UcsCcSdxFB/Y
zT0A9fwkcJdIzEwPWJdKNyrlEjvF3xFFomONFkFoDePtI4RcRHUe0n244rduMlbL
LHqEFwYPNLQmPXEpudAus+N5d5FdHjbvaEiLqkfFu+mE7VufV4p/ayPzRtooFioA
ja+mWkennHiYzCgAxaDopgDTtZB0ZcNKB9Ax025QAm2FNmXf/4XMbAqNti8km6kI
DEF1GYVKNx74G9l0blZeLvvJM21f0m+e76SzlUUf0g+1pezpCQOLJIYG8TY2MejK
g/cb5NfcPJrpBmQeqnN25lIrq4QbI1HZwmyPrCKhVtDofY8tQAM4tbxDAkk2lMKi
7udRKBwu1+Vcha+vYnJCc4X6Dkcv3p1saSH9ZG+grZxuTozpVDv1uzx239XTiZ5Z
LaA+kb9MgP3QEbrFW/S7ssFuif3FR1gTZ//1E7SZtOAa8lTE9BUuYaaalm0bUIrz
NrRmRlyi1gziI0y2+YYomF8ycaT+2ZbU652OsKuB83Iagx48F1aBoeXs6ji8Xnai
Q9H620iPVw97Hyz+4kz9ip6Q1i7PLh/7KY+quLTMSb8QSVJqF8EDwaEZRQ0l1Auu
SAY3V5JXgsXvkG0yPqsFM2Xxwx+oJqLUgIgFoXNlSHPbp8DBbmTWPBlRMFWOl2oF
tfgDGbB9An3D1T+rio7FgIvDIEGP3QgPp4+8E91MlP1B/0XF5cl+NfSQ9jmYihxP
ov8EXmlemT74bY4IrJJ3T41sM/RJ7HnZT4Kh5nQVLuFeM/UC2fDqbUpQSZFAHvWp
Mbu8TwHu/aiGA6fcwMUAyobjPUIfzi80RahBAc0FwJird81Mq6g3vMX8lLJC9LBC
Y17mXPx8qfv7TP2vE6kdbUsr4i09VduM6e7NmLuIEmEvKABYTukI1hc0HwUSDELt
v0aJVIiL70BYE6gk/ZiCn4CfH8g7KV5zLG/tcgca51bDnvDSqXIIxWsaLjatGOmd
g7YH5wqhXrsXjvpepmnQv/V/Q1Gbvy1wOEk/8S0UH4XukA1yBGQuyQ86M89CBZaW
8Le4dZYuGIGp+5D+OB4hBH6dd8T95eqpahskbpfQ0Tf3vGt7YvjUnNGfELMa0dOm
SIXV+I3lOrgrqfRT6IxN8X9sFSA0vCp4m6XWT0wKnPCVpybkNAiLU/qQgWzJFIpK
JYCbdNv31kiXJaz4PQpKDmncohTMcWM67fIDoP7gxEuTxIOPYCQj6V63k5FmeuWj
STXUdN80OIV6T7QtHwlIuqp+ZEOh7PU05rnUGj0UW8U8OM80c3hzXHJXqoxpf6w+
yyZ03zl5Fl5Blp8oovXLC4OBpnd8FEJCx2EmIwEqGZqOObnhor6Mb4M6LwZ+o6v3
h0MvdqSPhEPYS/GE5BTyBWn5z484xuQo9wwP6nEwN0XBOEaRBLwoV6cQRv+77rMk
UzBtqeWkxR+VsbDqLOMJ+P3HcRby1IQJFFmEQ8U5O/6HuMSuZPSbnFywOB257vH5
oazctm1o3sZfc0fbcbIHA2cfpHjfaRazeh9Z9neYx6mIhC6FH86Q2UwM3BSldZFo
dPgCVm7baJvIbf6FC0Fssz/bbnRJbKArb7hrMIRZvVbcFQlPEVnkotMEu8mxdyGA
SLkg9MIr48a3UgNOwxDrn+tvLRLiq6GI4XiSuzOj8PYScqPrsGSpUUilPl5ZhYGy
9RLiU7WEA35y72+QMQMHxiA3FKhFJZfRxXz3Q2SMGl62U9NQytZ6UFOzVi+uSl+R
wIW4O8eCPSWx2oxis/I4360mNJyp59AuKOW7wDYmHkaHOmVsLZ92uUK6JnCSgSI8
UeYZOIN/p6+SYf0yl2tDKeDsAG1iyt6VdbyXoIWqIFu1eeYtveJsOU8TGmvZFtry
2vIDhFDEVj4rQZ5SGK4Bmf1aPzh7/ARuwORo7qYr7ijpVdCza9dPm787KYHHmGDU
3/yNcRgaqToZh5ruyte89+3aaGWS9ieboHD9jNIlN8r9jvoX0zNSTdt2DivCToAx
lqBDI/+y1kHQiWBpVV3nkxB18a8VSj3eFQtNGla1tWDa+9p6tUcirDsY5dK2wHx3
izdcl46NySokoCw+odLCsZPNykGo4fcO2gmlzTB25oC2fpDk8ArkrFM+y8fCx+Ig
+SZBRq45xxGppyDIoBw2MfCeGw8irQKV9Eidl9gCcUKD4vTC1U7yZ/tcsIRa2VUr
jhUKYn9mXEGQ0LqoO18fkSyBUCQ2UygDtGvcUEIeAzpnfqjMFDPRx1L9sy1Eex7+
N0O4oMS3clZuTcnqbMef92eBCfys15zNVedO1c+ZY+jQqV1FYWrC2z0lazCZIWdk
LkiDAOg+OnNkt1IN4ZoXuAboYRS8MmHr+q8BiWplQX3lYQ0OReh4tYtRHDknuS01
GGENZ9Zr6ijx1zN5QXap1pAlGVMqZSA8xYqE8491Dv78sR8YhvzRKhURxuDKE/T2
AQmkfxru2LUbUnxQ+y8g+VCsgxOTkbjj7vE1PJMAp7TvlCdxoRgMFm9f1pBTknNK
UuN4TIOnAiR80dWmUgzxklRodP7eJ04JfpjU4UNCuCH4Hwf0Pm4+eDIIKDj58DJ3
Frz0IPlu9roYQ4SawNJOGk/tuBPruRc/S+Isvq3xa0Z0Ee9rP9okwCvuVOQxmPb9
B76xQ9/6ShGQGA7FkySGdr728iOK8NmSZsMYZvC4t8F1weIPhoAtCkKlBpiNMYtL
ltf46wKfFkVN//iDiJy/H7uqRXxIwnnxPpUsAu67CjE7ww0dq9KEoC/N0YSyXZeg
jFj2zhSZ6vjOhjbpnHM6/CUErmKAMmknNMq7OF0aoYOMunP4iY8C6aGuT1wlxQ5q
Hgxx4zGPEQUzKaUdz48sUorOG0isgV+SqKRG1tN5dicKQjdrkRa3ZM3DA4ng6CXv
DAvPTYz6o7lP55N0jzOfMqMWuMtRal076ROIj66/tNwcNuDqzT1B0FYJgNeZOFm9
cuYBSpZyevRTcLVmVyo8oz0s+vkyQ4h2i6hLXl5QtK3z33OSTpnyaDc8L4YLcVb4
/F0RL4RpWewxtr51Oq1XLHqiTjk0g/wiBK5PYa55J8agGXPy1JOKfYwhiXMpCsfT
5G79/J/5bj0P1uuFDWN4mIwMIL0IlC/tJA3j//EZeOe24rTpi5kJqQaxtBIG1GAC
tnac0ZEPaO3OkgsKsvECH8Ep/48nn+qnH2X86+JQVJGE8hRiVmBLfbUnW4ZpVjVO
hTi1ys8CBz5K9mvmwHyPVS2l98NBeTjki8/dNQn5qcIuVQRrAP1stOQqmcEuNV/C
Bw4LKtZNbh4HFCLQOrHAOFkzhN5LCA43y5y8LH+GA4X6u85pnBLDu9JC5cHDsJuJ
Hr5rzeD4vpQfZw+Ky3jS82hobrAs/h8Ta6FOTf7vQx2CvnmgOrchUlZHgHb/SiiJ
X4zm851N62WHVlUdOkWJHxIh4aOEg97LKvT8bK2/lcLVy/TDR5GnhK8zdLTQcAlK
HXBzN04xWgdd22MpMQ0afH8Nim22F7LZ7RzT9zqNEEo6jAXH6yjEaR1C/4DoQ300
kRu4S5TYiY6V2NyylLH8QPU72MoVJ56vX4RrwGME0HhyKjtmziT/hYKHidjQTalX
5dlGtCZDAmBlhKPZP6Vc/2rPX+8AQVK0oNPbagTA96xW+mILDgBXHO5qecis2iDk
vD68EMMJ9CJBzWmz63SPDqXCgR1XbTrSVDhVy6ze7PD2J+sKEUzjogd+4y6mH3Vi
4CN7fw3Clu/U9AupBCpeniZevflz64HsTKN1cfwkKCl+5mLcSFNfn2R8a+4IML6z
FvTJTF9gUzVZGg6/ebb5O1dKYCjlTQLugJof2t2disTemPqpMxNzCUjRfMEnwV+K
1SiFdIJ5GFUSlBtN1FifGhfPb5rirhT7yXPg0/kla/Wv3DpNzmGYBmubW8HxH0JV
vtpmo12tPb/2+GYepHxNh454kgwN4/ZK+h0nn98juxNLGdUMw++4DKKznJLTB5oN
SwFNVqb9eJYBY/RGTgUfUyMoUpwbvYDescGpMHiTga1OZaiOnt6a5aPLeX/L02Ey
Fy9aJLvFl+fISAi66+iGWxTL41CbCIBAO2HKcLYfapyp0+ePCw/TgjY5xoYLwMq6
Vtva5yIHTQygp6xMT6ftBcdTJmtSePztzov/HsElqEt8qJ/8biFuUgT4gWEu8Qbj
ZJmYq1Sfd0vvVdNB+FuGYQ19Fe334dKgP62WX6rlLLhFcjPduO2Esu52DIjWxpzR
Fc6KFIkMnFL0LnoCV0RKNAghh7FiXMVxy+g6p8EMK/m1wzyJXQOdnt6YB3IPpGKi
AgK7WLSkkhBq9ShWnNp3VommE6Jbb2+FIDDuhX/6RxbxTgwvcAVInNTvTidD0NYm
t3rJLoH1QfbpiFwni9EQItU4jPDKu5qenBCaVWu7yqTIlkzygUgCZuIB+5oVLTev
Ep3JqZBY5hSJcVbW4MZvSi7e6mf+Ks46Y1Wj78zPgGAcmKzVEOK3iUfDfF5PGnMY
Hps5p1M2yz8uD67ruX0b3/rH5VhQDIfOgLHqB1tj+nEISLKnkKkt6ME/nc5O1G6i
X83Mkjtq+bNok1k6DUAgCwHy9wu2M+PcnnI5gp6KC7vk9OKVDAc7ApIjrg6WBl1/
lo3c5WWX6ie+THXqqgi5mIjLgGFOt+Ap0sKHRx0+7mGd9+7fsoHlFg3IIg2aoF52
PNIUWTtFJrVE/qZAL/hYsCouz6xD1XES9KmJUdUiD/C32MxEltPNHf3aaNbQJEmA
aDBZK7Yq2E4xyagtxUSsfN36ZqEsXK3SL1F9h5Sxk15SCcAPFs7YM8OaGlfk4Cly
wzRXFEkCVy7WsIuz58Fo8SfRd+qFklP71o117XeS2+g/VGW4Y+LCrDvv+3JLpoX7
Yo61p0SIo0O53EM/kLrN3RVHOFfVgiDtHUcfsj6Qozyn9fXrFKJ0ktV0qQE5ZLqg
0GtOG5/e+mAmkb40ZpN2yBPLsn9PP6CiPXqVNHNTYGUfRJXYXYFZWYRBy/E2db/L
E/0gV8+2RBDOIlm7K68BaQJdfGGp34T+NfYPOJs0gKVuwiuGJgT42xMmnan+X7m2
0VfaP9PdSCEcdkKxmI0vF/bhmN4kuM25ZyC/c+COKpgaoSL/QXaZyDabaXPHXEpb
+jYfqeDrqviF/pFAmekMF+IIQnytG5/QpuPPVxMcHmgf6FQNOJaeo5x8YoetA+S0
ED+k5lAjzuHqDYQkUFI2EM0OLDjc8cUZx/CN7jqrC43ceue0pXzxscNpAIxHAR5y
qU0vaXiWRKz425lLAuuk2p2F+AktH3HixM+OZq0wwFmISj31Xp1Xrt2OgTo3xVdZ
zP4cPZHH45SJpCMEixEWK5nq9rHdm9NLBERbDhgDjlCgNudt84+/77ski0ijQNut
1sQaHpdQrVFGOujYH8J7GkuaAlpKYjSEU/zs9JFk/CLnQ4N1iFPt2XaEfxmT5xQ3
0EERd23n9xaImHoQffW0r7w1OCNrNC6aoDJfKQESaDP8sECnQEEdn5ALecP2+Vq7
WHikIMp4OK/DNb4q6Vv056eVOdhirIyNwlrcbdvNOdy1zFK3z55ubyOL4hWWWKXC
M4v4huj57zowg0hTu9Vqqsy+whCBUfI7iEwCTvmtBI+4i1LDQoms5b1WxsLtzSeD
JUYt4suOuNMwoor1bEaWvUeitwwaq2yjQTMueFCb/7r2Hbv1PHa6ET0VugOZMLid
g3ELJZG7IWuGBiP4U4OX/D9TpwEMzCbY3IQauF3FllcX8PE3IY94haPJmb8nGiDH
iI5Loso1muL9oIYgtwqNXRXNVjSPYVbfA7VqB5TtyW58s049iaJDEZg4dYfkAHLp
hXMLSof/UomHzTbBlj9tU9RS6XEqAFARsFekQXN9oZF0t4y27xFFouy6sNJnuaog
d3V3RHiZmWRaCGIEN9m1EVtNCdoHxNZWHLfnPCli95C2qf3APgg68Ctak1Jzljfj
7O17G+KHVMUNPMZp9mUDxhmOmqyiGlagXByvCtd5BeZkXaOfTtWui+RSTwdkS0bP
f7+5wYMQ4OgMID05cIE+oIr86DaWYX2RpHD/6pUFf2EyQivHlu8B8ztM+f2DTawe
XM3atf4MDvsr+cWKCWu2EJst/47peHnB0RH5o0XT2Ka3+M1VLX+IroqTM7EQHjJT
4zczoi5n3gjr291Ar8m2+n5ydRsqxjJMHu1OTqcAnuVNoONflW/sMiI1XQWThPYo
Zl8nsuVF/uJmj0wmgvZZUNghMnB+ky2+TSb3Ykrw8T1BBNa9eyjYXjahWI/WtweM
psXk8KJjaczwIHfRouJsusZtDMaOhcFiAwfVq/ol4gaVa8k/pL/VGdVqwXffW9s+
3god01Cif2nJOTQeeHeFR96ofr3ojyZJ5Km/5mJejqkfFfqNcqi2IGcHPSzs5CYI
lv1/YGeb64t3jUox4Qb5qiXdI4xQ7mHX7MYlojFGDfnS3WOrOVzbIJ6fSNooEeJv
8/GaZ06dMaCuQZ31NAnmwmkRWJXJUYTrUJ68DkrpRrBn181DhO0MFD91K9BSu2V1
SpSR1jlJ161KVE6QGPlEtx8zfNlcxsZ22dAYCv3rYZ0B6SSRLYrdTVzl0nqEcN0p
PQawfJsXwXjo2pgHxg2nAr1enSnrXCQ861wk9KeSK4mNiHfbsAPc1iAhyFtdSt5S
bfs46Ycf+dJsScLjVxVTnQqZOjqT2+FoXCiVkeTtXuBT5u2fz3LB8oSiEaVixtSv
jkz6IA93uLQaNeRCc0Rm0PeDVrJIFD6mefP6j56583DZPSXiXshuKcMt+G1t/st6
xDhj8VoSPtWthhDi3LuilWPUXM5Jf8WoWzS+UauFi5bwEoqEhhWods1nsP6he6xN
hRLHeQw0h2RMaxEUzVk4N4xbnyGdb/7Zct34jUKocShZc78jhvvcxy0Zs+D325WK
G2y0iPFtUuzOeBDQ2z3DD1W3l+xllKAQ9lHKRPnPXekSzSkJ5P5zB8QUk/7LMilI
lATT3zFAJHS1A5oZU/sm/ge4N/4ZrVAzJ2hq6IjMe0/qrOmhlNgHAecXUngqHNmI
hGhMdss52zNzI4m3evuctpolM1RQ1tvj+qtyPW15YCGUZCedd6H2Tcr46w3rQoWn
ars6aU/ACggcrg6fF8AzPwAjfAjd5OVpqSCEkbRuttKcrGbD27n8MGJONKLf8Q7s
qb75/Z0RnVbYnAvrnsruIhwOgiYHHQdWu/jA0oznckYFAmEevl2T4rQ900zzbGog
t6mv6+yu5AbBXMcd3lWg/qw1d8xhlKghYvvdUoyuMMDotylRUy/bV/J3Rr/YmL+E
6Ui2cDln+K0CeATcFLG+Y4nNaPEFyxglV/UzONHsteVipKdGbO3H2MbyrMaiLfMP
UwNnpj+FZo3TTDI5LDyKJ7Zwyd5hs2rqxNe5YMFXkBdBQQeNAqQDFNL3+Rg5afP/
dpc0cbnIKmlJh+I9rccH+V0DfY3chPp4FSyZEnoveYoOQWA5+TuvnHHk+vzDLl5p
CQHJRrs95dmvrwqi/x1C1GE3gIi3S/q0JsKnNaLpsEAwkLgLCYfjk5U/pKDXDvYw
q8bMKb+g3aDeCRAH2duj557xdlaDFz25KGcEz8d2+pJ+cl6Hs8pPdS+LVx2VhCna
6I7bo2wRxlUxydVCUl3mv69nZaR25G1P3IRVgTwJ/6MvDijGmj7UDgr5qC8W9QHo
dLCiPuX1ChT9yb9O/rkujr15rsN91CyVOIifbXYqV8Vu/7+WZFxwzSnXRqB8Agqd
X0brFVGP4rZhXJ2BU40EUtLHlc/PDHHuFOlrU7TeOAzbeyL0D3c1j4CU/zGCUw+T
2SVTz7Pl3lGwSXL+NItu351XI6wT8s5RlEpIEeQszQX6beDO3d8HaGv+pCuYt0+9
W8DfPrxrSXxWl4hEa5r76N1lfkXT7KYxpI2pQ+oIDNX/GPbK0PQ26/DNIV2bIPHV
TLrWqlDSRYiLwLpN7Rl0fXcAwsskmfZrqSmNE7XDuWrnfh8jtPH4jyLhb7KbHpJJ
xX+WUr2UhlxvyVQ4Vbs/7498OaIjTZ8bxk5iKR98AGXUV0kwlmCNNlvl0WJwR8of
zA6zE1Wfok78pBiy4PCMjhTnUGoeXIO8rEnVbu5SmQaSDMq2UN4MVfRqT28m+PB+
sqZxdukzSZzFtZCmfTpc6lsW79TmeQIrHEmY6dql7TKJleX9902KELscq3P3Sk4S
Nh9O9M0dcWPHhJFdprduhpFxQyAGxkvUBtjSB1rFAkNiFzKO0rcHATES7GySDOnz
6aTrGcGbkrozOjVApnEJDOAFsf3b2jxOs9DI4mLI7AMVRxwBmNDbjJIhQfDwFIFO
smZ4P/zgrij49WvGafUtpe6dHN0xEiQdCMbC8s0TyfattZYSwzSccSdZLLIVBSIM
z4LJEoh9A7D+I6oTaPcoRcCcFnufcfqKmy8PNn1xnv+3qk5D4pNgRDjcbkm/B7hS
BdxlEYDiBLW1M70KBL2xrKFE95Q4rcgM0Do117nRDsMNnmPtIkewWRakII5TiZa2
Oxb3HOo5aCKuRs+XnDrmCfIKyX1OSWe3bRVUBPE694mYD64Awk06F/rjs2G6n7Ak
iyVPTh0wfK8O5ViMYHUwVcwhr1V8rV6DC6u7Xb+Wvta1fp2FuAdCo1RRSVfy30bZ
ozJzXHj92R1qULUMOwJPCldGbl2JFbS9hVAynhvAjOay6Tv4KD6XbIUHcIjLswzS
D7OvB6FjLGqW63rFqey7nz2ghLWigehhG3XSOZGFe2LDfDzNyMNcor7iMhPw5biu
phyTXJUDyGqhExH5CRu9fO4ApkBDFcAoNRM90Mn+tiRtfdN4kId7hA4tMnSxGOif
tkLcD1s5lPcB0qtEd71GqVYsziWBugXNsSjrcbuv75Wqc03MD7RsdMilBUZfrYAK
4BGZlOZvnIMrM9H5sPaWlvnIrr29O/nBDu6nSYMVKzpjBWsiQMRPZ01JzOksbX3K
xHOFvoccRy7QjMPUZmwhnxhJw0auVWgA6+igzQ1gwomgnD1AIuIwzwliuOQ5D6XY
Tng8mAXr3PGiELgSKg3k1uBgYvRRrTF4esUQbNU+vr0AWpEgRKDQ7DU4ifcwQPfr
ilZvIDzWYoW+GYQzO2RthtArRK+h91Y/9NEE0dkn3xy5nuVXFCx4LEPG+zqDk43t
RFeXaLIv62kb+Oy97L7OD75LDYNnQ1F8ggpwWsIyZA3P2oGpU4UzpLIhPCDqcXek
zvO1KqtKa9bzEYpGeREZhP8LRxVXhd/ba02QpCVxEej648G+7CGHBMV/ZrJIwzcy
kCc9DYQB7hvXzCJingaQqEO7Ku2cr8M3YdPBKvVfZO8zsK9qxTIW7a9lJNumm9Va
p8YhA25oILeKy/ayCifiEOJTOm35qo/2TOrrqa9I58k72zcSDhVDr34El0AknLiD
7i5NCeTc67vgo+LGEug2PCXGTA1xjN+BnFNrIf97ViIY5THzv/SwE/oCl+Dz2Rf0
dtfJzmtReYYZm1wXSKni8OImjx2igftrpwrDB1RCaYb4J1RQogpEJ3giRQAA4IIp
aw7Xo3altimIUbCtUVyDuiC38g7mu3XAM8yh9VXj+qyRD1l+44Tya7lMbjI/JN8L
hmdtRx/sUWOpDtNNXVB+YsM/UK6D99Yp2yLawdvKSbTNbhPFlZLde+hSNBuK0mgs
SUjU/RF7DPpjOLp3WBqPFj9z3KK6eW5Hdyb5F8DiSLVVBSIwFDPX9Xwuhk7Oby2m
e8tju5ky0O6FV7weMLpMi/bhWVKYppeVxgkE0A7V1TZ1BU4GhGKuCUMctd5Xk0xO
3yfO65R8lxPXdEVZpoYuyJ/A1Nv6/z+D5mHkxYeLwjlh1p9cemUf5FdZPcXcH1L+
BYG0HIvGN6mjo//bbeDphEvHHMSm5ob4zF9AJlZQJ0jpWlU79ruRw5NusbCBYWtU
SSZHLzIFHqrCKlLZTk/9istPXmyweUngmCfH7tWpNhJLhQ9miM9DfkjujdSnnoyR
J/GyiyUH+lOhfFNLt5ae/+JZKik6AmL4wuaoBvbgaT6tQdAZWzzhsygTAkm+XK01
7C7Fu2km42TuWKWxuvxHAUxY88+wiy31B86bWvjuY7b8CcD91t2gcbTSz9cdMTw9
yXOECo12sOSJNxXapJ6YHbSnqCjd+6UlXp0Wn2jrrK9zqJ5OdDCbeO4ItBrdhtVu
NVAONZ3ohYLS04N9lqJJti/H1z9OECgUHevTAwiqx7U3jTJmWt/JjMS59eQdE++l
HBNDubmmp+RD9/omPzH+XBJ6AfIOBVbgxNwMoJDrYC3Ano7g6uBmCkGT8rRUG/zs
PpuwiDpGWwj6GY8mVCwvMMiKm3dv0UA1PYBlVeL3GmvYoaxoPaIt2Zjrjtk7UbzN
2YV79IKWElZT9xdzYkzXOodNyQi0avUhRQmMu9c6a0lA17Qqdx2o9s6oXq45NwoK
U5w3Mmz3BBl+Ql0cc2ZsTGFVDlcsMoW/h3IaKl5dx7vzzvDyPN1vI8ZltTTlNW0A
4CbtYwNc42son0sUpMZ0Jbbf2lCz65JHUD9SqfIei0zQbp8Vh1aeiklxEJ0VIN6H
xijeE6s7X47mb/7GZmGcy4pWuvbp0sX3StGmf+H04yHyZ08HN00EAGwSt+Im9rul
ZUgmury21kcKEKvwMWdEllwRLe2h4J/jpZ+YNPugsLEQDh5OpWGeh/32IodAQ9+p
Hrb1CtV9IyY/qVjPSMqMuvsJKqvyA4h+TuncNkz7OwH2KV701PTXzxTx5pvbj4yO
yTfgxRExxDtBHT80qF+XKZIQ/dfUqQ/6skRxuYeONDnE+zSF+W89Xwmu59Q0kw3N
2srW0PS16fkEmz+5djKsUVKTCnvm4NPikcszKje41TCio7BJ+ZmKqEJNcrLvjQnP
MDD72mu3RPKXJrL1epKgP8ydF3yvmbS+DAoX7DwbOR4t23v/L1EHYOOzPZ1oPPut
g1/tDn6UggRHMM060VY68ICGgEIXEiBM/2ez5H2O/7QvKogyrx2fdP5NvnPJcDD1
DEBFxwZ/f/2ks57gXTGwIZ/62PiXuX0hJ4BBJElY6ljJYedcESCRdrO3axXqJ/jp
GcDS/SIRqG8qH83H4zqtd3FIZTFV6HxcPxMKCBwmBpRUsx13vzVmeisxEj9Cfuvf
S3OZz926CubhhZvBokMhlcDSK1geMgbyMj7dsDLsZx5BPGEehlNhEMmyR7Q8bl5f
hyk+JRnKeJsm4NIdQkHmEESTEhTX/RWSTaXTpYLfMH6TegMEPFHxLAT44zndCumd
R0z8jC86bisCbjXM/7/mGJiGMenahAibP49p1jiI4wpoKB5Fq49ioQ+8Qz2vJcMb
dusebm1t9h5VnjKPdhTJ8/QhdHhwTtzcf6W57dEFRGzNqj4anOask3H6qhri/8Y3
bUamFyuKzTnZDLnNMwlN6GLiYkDY/L6GysPSxibYJebHpLFnWYN3By7GDK0xKYeP
x3hmP88TCAguEmHWm1MY3LR5GhZjvlfu9DuB4f3uSnnOvfKDqqrw9Ozenqga/g4G
SJ46jHEmb2KbBeIrufqwCRpzh8qpFE8BG5qkIfQeVumODu768/m0JPQqZhDm15Rd
v9ly6HqCyui6oKWKLaDsTMuUiXUPF9dytuxRNzDL1kp/9cD1D9QPjOtYMxxshM2d
uXck1Y/zHtxczHHu2kb7VaSnIhyQTD8Amq3IGdcaqwm4qEp8gwHY7mbWOEeRRpBk
l0sO/GFm1Oe552h/DHXp6+dM4nxwY+bRDTdMBt9dHHPq+lZgiTFaYkkxfbjdcwO3
0Fo2c2NvkqGPRKPj0RSAWeI7/zcUgbmsfNYGXUjFIvKHXC4AvG+rMPQRt2fi5f4j
5TX2Ed+jznPFge1ioq2Y/5W36PMd4K/Txnuo7HjGzpETCs9Xsk//GiRYQye4kztw
0IfV8es96b52gRsA0l39Yx/85TewHFlFPTpH4iil2ebHSl3WSWClp1FikVx1o/uh
v7TjGXIkj9JtvCd96WKp1ZgBI58DgYl/1RCPx7wtJTwEO4kVa5xFuo64IOp6lCee
HSXuqhWEycy/YEqY2koBQ/agT7A+uYKY6QcaxCQ2/od4aydmcifuuhgeKi2UChrH
2zn6J9bt3cuyFCuZDiTvWsiUxyke7TO96+6YVCN1dUC+6gWbaosHQ7MsYKn+5rfj
BH46Mu0cZtAv+KmFmmwV6t2xwcvRHv3QIet9aicHLPEhBFCTsLZgkiq4PmsuXfpR
ARlGgAx7wCflTLBAOzC4EYfNB/vwZRvx5WMTeSsWlM6sJDZOVo0+23lXCn4xEpj+
kbubHP+65mrSdgUDtqsoCL9UHcfbjfsJdzh/B/VTsv1fDUitg9uXIyVmlNQ0XWB5
GjMXXbJjSgjg4oIO0RyL/KNXe7I4BJlDovViVV9rFsRAd9fMKSib1dSZvHD/DqEL
bimqfAlTKlRCgpDuQKG2j6dSGcdJK07p1YE0LUQIgNH3n4zZHMvNgYlG/h20qNFH
JtgKLiHbOZWBZxTSv1legW1nsm3/R7HW8m5SKGQAUX0kR+OoaSf3+omjI9R9dZzx
nO/t2Fg2+MwYxZs4oEgFozGDk00FYK/IBqzGAfuMb0mdYOTsB3KGSUb62iUhUhFD
s6ot8OsYXjbI9ubOOymLBBQ35II9XfnQ7wnDPJJsS6CkGDKjzMP9H3fDkbCsU/Cs
Ayx9SYf5BEaWfM6QUtFW3zX1VnIC65qXyXXEHLlcWGYmfspRp2ElyNdS8LgtmjrN
yaP89pL8pMMGhfzXIDYcPcLkfDWEVcyTrV48VY5AwEYzOKrToYqt3/TiNFBcYC+n
HhZzMv2LnPE8m0qiAVtYp3QRy4cWUV/IB7BAvWa6Bk1QVKqoA/5ejh4MNDzhn+/G
5am5ikPA8X+EZqkE4YYG4WJ05cSC3edhg1zTNgOwtn8LFldL8jLIJEorO6WxbT+2
jlLn70LTKzlD/wfe1SRd5yvRe8iD3IwpDC1MS5QFLZaIrFr9Mj5zOZY4qfZc51Vj
fxqoqwBZgTwItzKhCfkoe4ddD10TDeXWh4Ja9Ch8CZPvz4kk9dpmgJWB49T+TBdU
c3OkPJvVMOUfU6IHaQ7gmA/NLXO3NLLhC0NpXt2i/I/b02WJWs5yAzNdqVaX3az6
EWAxxmNxVjAhb288iNdF4ntJuhiVg0wU2hfFc8UjfnccBO7m2MZMBb0/poXpGQ37
el3VKv4QdrQ1Tlo1a2mqWuTyMXyip3zbC/lasNg9F8ezFJolg4LlvqzKlX8nNr3H
IRSkk5LKV8ITcPZUcplUVBIcz8558MzoMD5/ErV0Sm57BmBzgiI2AdC2QMXEQwj2
R1McdtsFAu6zmWaF5EfaM+Q2tXJQ2qvW8pQ0r1B5S9aTNwC3KQ5Iuo7/XNvpBB4h
80OMlP59zYr3axtBF77FQ7iYzxPly2JjnQJZ98UlcTcF1zbUSnJNSn/VNNQFQygG
1z4kEXoF2jG6ZjIfYpXhEqkKfZTamr8ZYrM8LXYhEPtACT44+Cl/7Ah0DPnf8kMW
xcyGCSjPkk6S1/wQ9cj8M3oMzFl6s5uxYF0dEcem55M3zjFgAeKzXpUE3wAtjjgM
dL7zUDVlbaKkDHjZLRDITaFMFa/bzghPuQbmHFg+R5VBN+Sq1h6PAVj0L9642Axi
mR37N6A/DSuQTCMgla1R+unUlMyICHy0tk7srBXOPI2ZrSJ+lhNVae4XKE035WL0
eG6JL2EQ/+LguK0yav+QjyT1nkthbDmLh0nHFUInlk95kHveLa8jjxehHOiiXSv5
nBGsyLhtKhnK9+zrYDO0q4WZL38mkgN1VnHr1prwzLjnNbH4UXXl8hnHYLJioOst
hdNrcJrk6FLoze+X2toaibh411l46oSGxCTbqrpYk/0KzRMB8HTcBjTodEtZqinV
YmHIAXsCSQKmCwaYtML8EPcEWsIokMwIZXwArWiTdsi8cSYa2PXKhB/YZrEIuvfS
m90uDJp0F85RYEiYnZEt5ZUnqltpAfySQuzdVWB7eSbPzC2q1H5GyKOZk8bpo345
ZwRaSg7XSXvpBJU5FSu+Ds1sReUmnB8G0P3BkLGqVIaHKWfIdrlC/JtrYhgtH/U7
cpj3Fbp/Hb0/lLu1funVXbTuaM4CoOGM3PFuvPBPo2HC7oOUt/yHjmahKLe7cj4q
1HQxyZdOhvuSV6N90/lOpb9IoDzPP9olMUIuegK1patE4Ut74yP7dzQgZH71u+TX
4G0lyRzLX4eMgdLDnu3O1EmvF9EharEYIbHTH+NN2+uvz1fwDX43WN9M65VQ15Dq
L91mn83JZxirAFXDoseST5LFMg72+S02WXgM4IGZ7yjnFP7Ah6MQPsr5sgvs5fbn
5XMoOKa20BclvCuhcuYV3dZ+0zPT7iv/V0hILYv32vspzetWKiGe8r/thFXjW2fq
LNPr9z8czJlpoROCqAL5k6epclMG3EAx6rzuz2uQuOYt3mPdKvnlMIsk0J7Dez10
Kc6MC6GCxIZFLFGS4vfWXlOluJWvSNWWMlaQ8OUceMBlxD0ITRFeufxJrjPI2cex
Fcg8kJ8Q5yX+Y83Z4Yey7AdVqAyLfa4nrHy6VttEvNoAe/XnRvwHMknsVJiqUNaD
gN0FHvaE6Ssdlfq30WudoZeK9F4BWSUJ9fLfumrvnC4XW3zn4Vv0pIKiup1agjYv
myC/PwGrbgHSTI/uWBhF3Q1FeczhUXyug17dyj5OCpH7lEuBrZ7Lq4AH90LytN05
5R0heyyw8AmkuWwBmDknmXqjXUFUSHyknxrdTDoG4lnR8kDolOXE8bOaNNOPk0yS
rhzc/vbk9/CvEGsHEI7dpSA0qy0oxUfqdPbvRmU5fz0mdre1Z3Q0P6ozC0yV7edT
afG1dNDhEZYD7ZLM1rxjoNyP69/EGjpDyO7h0I4r5StCftV8nKOJ8aPEV8ChbzrK
CKRKFBL20Bhm2OV7w29WGlQYidMDGMEoQAHaaEe35jOzqlKNNkPE5yLSv5HikbsB
3ni6qWufdUlF4JeWNu/d61zwFQ/4z0+H7U8n49DdqOIMd+SzXlKdod4BSUnDHVhV
5t5Kq/7RSS1zaJlC8drt7PHp7pjp89GUGSOwaO4j+I5FpqeI2UCXfgt6FSygFayx
aJf1qASgFqJ9OJ2e6P8yFk3GGa7Xnqis7zLl0v/PsTzsvVwvigDgbG3uXykLlhc9
vrN+/X+Mfzn5IY8OvUmPwKmBMafqT/VZu5JQocNieTg1ZM4XPGieED0U2Lr3BaqV
AgLKVVz856cmuhUOC2KHnN2oX1IId6BSiExsY30UkG2SCFmC5YCGE2SlUp5+CbOR
79aY13kM+iMtv3CCY4A9rtXtQONknT/JeGxSOz7TZi5uWtdH0h33B+INFGoBmcGO
w+iZBNOtp2EAPf5/d2NcLQ==
`protect END_PROTECTED
