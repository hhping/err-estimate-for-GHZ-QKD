`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u2YtHoyejkQ791LXZCx6nOudCIBbP2OMrxiP52oUnvNTP0isyX6L/c2QzxVElHlg
F4dWj6K6uhSZA1TOrpMsaYSBKap58WYANlsDHWnbX2iPxZSUvi9c4mMkLlNPlqkh
/VuGTBPuOXHHraKhRoNF8+/VIBRX1AnKGqy4MfrRBbOyrfT1BGWtyY6Jdk55FH00
i49Fg7tOe+LNB21YOAvNamjQD2RakYTJ5bHzBO01/5pKpJl+kResq+0iiafEzYu7
8UtaBpq7Jpi6bPIs/rtpuhQtfQg82uaep+0pyoDQx3sD4KFv8il7Ihf/pzGHBrC8
ZUpzh9um1GC6OOjdkvs0YpCM3qY2Z7IKIDdI7lYbTDiL2IgiA+yLeNYM5ko5zlrP
wwEbkxKL/YCvIw4hdgQbEZCIjqw7//ro4hPvV88KTABvwUS9d9DA//HcZTAIHbRg
BhLVywrO2/GmuO+dnrSKD3RbeLsJB5GD9QVcfvjk1W9Xda19FUXeYe/sgDQngPJ8
0fNw5HFtWwMJlaLowc1lo+M/UtBMgCLWVzHriAigbt3zlajqK+AQp7FFhwAG4qgf
5w18aD+7O34KgS3++Auib7iKd9q6ZaAG5CbPH/xN8wyhszMcX813c9VuJxm6Xnaq
RE/H6/07TLW4evwCMa/m+q/kbOt+Wp650hpbW0+LQChQ56LMKIjbaNvJ+x9bBOem
OGtYbXvYnrnyJavG1eJyC5u55iYCBC0GM/wsuJ3qozexA//NWTMqzdSPdIUDMRJv
klhUubM0v+GAmhWwZ0TZlK7rDQRQCLvmFnUT+d5M0zSDK6dIKGMAMAKzliDJ7tuN
fpOEvcE2FRF7UNpUE/K3vW4IsJPNjYxuC9m3Pg2/KlwGey3AgaBtA+1rdMUBIrkY
naemPNZ0GzdK97nem68/oZCls94U6K9J9JlIRw6Eb0YXot9122hF/VznnwnbVO0P
ZwzQ/tVZcJJj/2uogMNYZrqnRs5A4Pop+d0YrfXuX+yTiZdCxlYpTKjALxYv7gZd
1NZCYqwj5m7YrFL0uoaCX6GXWZZ7s19lpTwIySaqFELJDRYLdtPwTsCtI4EBJaoW
`protect END_PROTECTED
