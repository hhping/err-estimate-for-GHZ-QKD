`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J56aW4aZmuaJK7rbJUyiJFGjrEOe0i1Yj9dEkTbYjghl59u20ilnTcs49XkV8o7h
7XO0Ap0TxlhfNoz1YXXLpRi9N3hZlOY92X28446OWQUq1Lugn4DeAO6T/qO2DKhF
oXgZnHFFHkIx06yCaw1cj8XgPll5l5ixQMHAIcIPwvB2fWXIipHph+ZaBs03MDiM
nwLgT7dDGQ77Jp8a4oakTb1SdLWwcLlPkYmkhrAbJK4oVKaEQANBJJ6tUbnAdIQa
sVegktMw6jlO0V/C22o7ob8mELe2UasVC4UUWQVw9/zF5H2dWVEPQNCGXP9NjQUK
7Y+FO1k5/ct5sTiUVL+mK6POPj5XC/sMrF6+duk4dXI6X8+XCN+Wa9cvSNgpp4OL
mVDUI9s1TfIa/isE+Dz4qn+pWNTWaYdttTLk8D3/BNkFKYO+8Txk6ih7c40XecWZ
Hpod8yVqwLNRlt3AuX3IUsq+nnN+JG4QM0R4oB336hmFbBKHDXOwWHAG7N2hCaSj
socae9Zikvohla+ROd/Y4+eidAv/GVeoFuMrFXUfxQdIGfbq+o0/DCfhjbf3k1m+
mj5Bd+zl1kiJWmqjyta5/SkF4G8uYOmZTUx7UCyQYSQHt7/+SpvmbWm/9EHgWcyb
qOSuQ7XbUGBGXjW4C51XSwP+oh25bia54t84ZQUr/m/HNQQo8/No1B+x/MmO2EY/
tr+ZHKGzFVzKEw3rDQqx1YxijWDDrirup2b0+8DSSS84wezbV51L6W6g8rzExUWM
oErrC1G+McpDHQ6wvm7bKynjdBi0z2aKaMPOSC94Y99daSdwK130unnhMoweM4y+
n9EFTjPuYi0VGUDSIEOuMl8D+Sj7JsAnlsVw2GdTnl28xkGpKTjpb4INLgvq1v79
8951j2SAalzlaLUZ/AweJ04sbW5HCV91/G4iXuCdqMlv0FTWm35MZGL2oHjNYT2g
r+W+9PcQugk+E1l4Ueox36SbjQjQAOEOfITc9lmPX9uAg8Hpo6N/28e9iqs/DCs8
JrMcbWElb3Gq8p3xwUh899JNJGsqGU7bamLdNA+XUh4892JTx4PkZ0lJhqLdsb68
D6Hzdyof0LmUqTsM7l0Drt5BdP582GXzN2s8dSzkd4ivpLHorT1oF7qpFtW5Sca4
F2vZwEe8lXh+ptanFDTqor0aWnX2FzgGjrryNW115Yu7Z4tE2hcdSEWNOBSwCylU
kWDs3tfJgRgfaWSOoKJxFrtLSETpiDio5mJUcJ9TQ9ugdh45wbAXSBpYGMrZ7YSF
M10MlWLZB/ShQPigpNA/9Re4nNx4HubrsqsHhyfdzpPrPIayWwuyItsD45uSGusc
vSFaN+fISPHZHx/bEnsOw4snJBmYDZweJN07XphLocuZ2yEgU0OOVIzQpav/Rn5h
SHrjaRG4jih29IUFEdbukLqm/q9UBTCUQn1IPFEu/e2USG4O4DETm9OyJ6fLav9b
p7SohpHjk15h8XAKwbzR1YY6nXplaI7Rga6B8x9xhKEHG2jlhmisKt3t6/8MgL3K
rgeZx5n1+iAw4s4g+MpgUXzQ7cPF7Km376OCOz69CJLwNTinlxIc1khB51Sn/LSD
RloMZfLJJpCHgGi8mpPnthlVmORYbTmeyzhz3abyEuYGlTpQXRLlvWxPYupAZXRf
RcMVTZderm2Eb2LiDfyjC7lVyOrGva7sgVt/x0/BBvnZVg5OQb5ANNFnWeYD9hMd
5CeYPehzpT+38PLSx/mGBE6Aog9A1F9ucyLA4tqwF/31hp8rl9llemo7ic8QMovV
UwcWCNDvw90cw4ZXOywkgspJsXMmxWaSIQF0hqGoD2Ao6YCAWziaXmKHj5nwxCeC
yHe3viO2sCRoXu1em2x+Jz+tuov9KtWyQ1U+Uc4MmOA559mHkTN5uBfla3ZLovBW
bTpVYZyz9DtM8VwOPnkplh7F5BG/p+052TgoaWqRwiDIZ6XSWXKLvJuTvodRLVtq
8vHVMKOizo3nZgR5R1dDuHx/7WB5LLKnBu6by0AOOL+lGXjtJW1dM46BxFRWhn33
ZdtRGT6piLTY8w5wWPfR0luUnbIGx8tOka2V4ygEKUYN98hnsrH3/0dBXGr0+2ty
+lwFLPfedV8Uo0K7oNJN8cb/rvWk7xj+tJ8HVdM/HoVijOpF/PiGbtTzlG3O7TQT
8syybKeq6A3SU7JXvvmNUiCVaKsK0PSzPANuTeuykQKjl2NBvz9Frhg/tQv+6IyE
F1AvTvKg26zR220jZo2xsqvUIGhqcDgyEx706OnrV+22dKFqSyY0AFLWadF6ZmnY
HJjourW2ej5JH7RVsC4Qc4CcPwoIWK/zxJnBIGAwbTceGD+ESMA0XKtTSG9QuQg/
8xXaP9buvUGDGdjrJCO1X3YQC9UZ0xHXKsILci195yxgeDZ7/zwQlAc68SmiWzFW
YTPvEg5dxNWKC4boY495JNv7nOqrUgocN5YDuWiS6W4c4A480URnbNVpEtzxi7WY
o+RdrchR0dsNnp08+Fouqg0q2kvllyNF5medyI+Na1xu9n4o2waePIo/DPPTPdVW
X6p5HtpE9dxxccr6FajaShy5puUg5zifmOXIN5WXODdYUtdPS/Hp90lxEfSYS4qY
ihodgPM2qt7F9NSzBUOz5CWbaYRvrSTsM4+g/CDipulztuenQhafGCx0LuUXnSTW
4P3dDSpKjiegHps5dL4ax6PsfvSpH7KjivtyO71jZRb1ijGhodL/20WTgocQAsPZ
VKGp/3ONPepjZ1iJkG33e/Mi8ckNzEU5hUDwuM7bPjL2iAqkrOlE8nCFek7g4+Yj
LRVFKcovdHh5ygEWUpSB6a27ajd0sNnbAFn1ubbANpAnpstivqZMmi8qMq4X/Prm
M7M8YsZ4nxPdOnKeoXX1Dm+VHfSBUJHmsfjwXi239JcWCUjf3KnJ0qygLK+GSHR3
ZolmL+Px/3kyP8CVSbasiFDt7PWfXSlgbvh/Keoex5WFb3usUOL3/a6gXQdYNW/G
xGwVfhwXx2YPGmWRC5DuAxebcJNLRx0dIspFeTzLveCcEPb6SPhYThOOCaptG+NG
6R8oyswKb0NFHNKkOseokro0LCruuiZMXX+AoeO0OFfvx2R3XogiBhOG3GC2kfTf
g+JfI5F6dXruTeVPooSEWiW6yb3sJxzELqSZrXjpIHNwqiWZL+pSw45+uSj0jRDX
EI+SLUlPJhTEYTNEP5xarpsh62D6tLS9qiEHULXFhHE6gwLeCKsGIafUaHavRMV4
Yj0ozd/+oBFkbtPwETenxqeQctrLGWTxomL8M3oIlui7OffGEzjdpJHgVzWuu+gW
2zfZHZaWwed3GBSrmeMnENCHJlUFsfWhojnFM5c5IoLsWH23SqfpMlXGkPLTkjOr
Em/xWvyZ5VE1RO6y2Hrow0x4xVJSfilCdInBPeltbdvxLRTbT6w2j3EGhxihEnrO
ynzjQJ7au2OsuKAmpy68euAyceiWMwcL66a48vCfYP4iCXL6FFgvIYVO67cJMrhF
xm3uBLaMP5lXs8bWaWrUzvxVjTFUpl8rDu7BX9dA+u9V/dt1pY6D684q7DJVRnfb
HTYvzilj8/j50F/sY8lKWEeTjTW8dzddn9UBCZls+WFXr9Xq91d4PzYJRE1Sx8l8
vybUKQ5aSSHmSablxqcOKUAqJxhtjKqBczW0tPIZDkcg8s7ucqIU1T6gprxXI7NF
r2ik/75SEJhlwUaNF2TOywgKVRCIemq7rL26Zl61lQGHsH1VrYhKnForIy1amFi+
/yRLOOqE8OZ/oLsFpXi39Ou71T4hELyTC0LQld5kQK59aDqvTD8ssHY3HAQ4chJc
iiKds3erTGR9r41d779gz55Bf0W7wY48g5AzfyqCcUsBBqH/TE1myTjtFjakOUXI
LREb2NdknKyeCzDJ1N0aYf7mPZjhaWHa2xAmgrrvpgdTuliZpj0VDs6X2QGBr2P3
H09+3uEgcPY/zWXpPGN2pb/snIhEmh4bCCYwckeMnTnMe7Yaustc4kCyw825lqoD
dC1N67OvE6GmddR/xFF/ddyMI3lHKdEEA4rM5J5jD2hyI9PtO74FcZSNNNObB6/G
kqDP1xaVz67Fr0whqKzXvXBqOPql3ThYB312ev5gicNvBpxRH/l5W7yLwJysBF9J
u/zJtyOr0nxtRlGJWvwYXdPiVyJD4YibavxGq8fEEMDFbl+UGzbJPaH+p1waOAV4
OBq2FiPwKeEwaGlvzkrIbDBqT2w9Ipt6KwpK9Fdrm5VczYkNi8RHAE6s/T23vpyl
0b1okv31gouMURAVCy/vCX8OAnOD3lS1r9bJ1kbW+GZEOcyzkMcpeqmqO93PVdyM
TdVZx3p+aeasBiN2ZzFbqpJc3kPO1J3Sy5CbG+uuqC8czCTjRlXl5Ss12jOKOGJM
4SmOqkFrNm90XQM7HNhhz1ejfvzTP2+Mzrdmv9U2Pamu8CtEaxPC68XwzYxJv0mk
qoJHvTAZQGgYUkW9/nhaDusc/754pMm7WZ1Zg2fPjJ77yz5T5XBdJxJYoG0hCfp8
8Ncq5VTLnEPRqFFZoX3vKic+rhX8Nv6f50nd0Axhh8cZYWwLatbXBoHAvCICygyK
vOCOXEZjf7MyeTKZdy7QcbzExhuMD6Gd0YS7dPG+Xa1AKeI+Ez7R8QjKUm4k+K8G
RIpGHlEuED1ErsXvAtCSJKJ3WDmROxfwcYiG+g/WOT7h5lzTprW0p+TU1FH9VvCD
pQRmtnAzR5/WAUy+hG/nq83BrLCZP4jjgKMQfp1JL9l4WudeZ+3KAFk2sIg24lfv
LLih04HYVRu6WWjFLnrAF2xXvF0YBHn0cVIveQ7FfgcXXl33f+CYfyMjN9Y5+/E8
CezQZA7icDFa4GqnA31XS1qlpbkfmdTOiHcAZB5j9ilqNyiu9882LpGNaTzImExu
W3YZGQDxatKIrmHR/lT26Cp/gOXEfJEQe/iNUDQfJ/pWQQvFus8u1uL3YmJy4HtO
/wsNe/bRPPr179uY4lcFjrB2mTIAS9KLNEBLh482pSsC+VyoKMKabKn4hD1JwZNf
G6ZwHo50m6a4sjsjOzKBYowLCQ/cIXUE5H2uWsmBalcpROenC3KDwYmuEGrtRQu5
02+P5e+dXIUElKiKou1zhdY1PCZWcwzi66jtMXHz8yoCJmQ2Ah3TnEmVuBURNdZ+
pZv68+y4cKONZhodnKlEv13ANsTNtQqnTZ44wet9JSVz+K1ZY7kX68MFK3ionpom
q/FUevrxjtsJPSxrRwoHQPFJdnOzGTchWAZcaMKxUSnGRy+aQfJk3f6ydLT/XY6G
9XlEtnb/T5z4WQYjjGGxXyZE2jZ6bbvHDKLaZMAajQEPlRTLnx/UPnZ/lxOO/n+O
DSaSvG/B6HefRG5Q8PUGbCpAxVygdZj0zufsNHX2Us/StV9zAxFm6uCT7vHCS9zG
LnBT5W3EBzA+XqrnA+OkcJzs/PtZ7R4kVVdV32JVheTWkN4Iyp1mveBOLr8uj1va
ECQxLpLMTd6d5m5KurGcm2ZvaC8X2L95tty8LuMS0XkP5zI7bVB/MRVSRyzGNLXH
CbxusgH2UHlV1IUVp2qbLWCTdhL6Rt7v8CfSidjycpK2jbmT+0x8nK1ddZ8Og11y
dpivHhzNmbfqSKhWSfJXY3S8h/WWJiTUoRZVv0HG3qPwz3NQnOYXNHY5leCQ4yJD
ImzBu/WiuL2x1OBoWMBVJKy+cSGYfv7QrEFPWuCwRUsO2vR+ivbGVSM/9KbDL2fu
SFYYPwyeKOnmgMOASfiRhOzsQasvJveUX1d4uq5V/mLZ9UX2ber9v0aZ0pxZW/h8
236zF6I5LTp3M3Jx+J/5PkbLO0uK5/xURdPy7NGOzWVDfd3M3TXxsd1cydxq4P0M
V7QalCdfx0XaJJNeemKHubMIJGByEp7Hg+lTaOYHjDGPmukjCk7g7EBobObU8PlK
2U0LwaGwUKihKt2a6YbDo1vFJEFTUvScMuz/hCiQnN1ItW9ZQarzFZBG7X4Fpv+W
Ct1ToIEQqh8lXJAZY1l6I9+u9vPcknl9+2YCFU5NmRTvnh3TQ5ubbRvTEVLw/HCp
iYAl6s2YQvOYUdUHwuaWEMq5udiLIaCatq5NZeWWcG7Ipp8PfA0L8WofNUkHDIpS
uQsu2DXx81IalYIS/oZF3oGPbUBwJCUflv2U8Xucuj+qQkDvvdqooIohFmvMl1hl
xt1cJYivPR9a2lBh3fi5z5F1Mfzs0mLrw7aAsw+WYY6TG//JU+ky7YFqy9PmJJ7b
N2pHbW9N8yshA8HsvIbTu68GbAN9LgG8TLzjyZ1LDjtcXFT57mK0tww/vw8TC4U0
V903FgsFIxf/8eEv6xxLe3X80v8+xMzzp/GEqM518Kug5HM9CDPnYLIMnlFOLYel
0L6+jNIcCZxxbFb7nhPnhrZt0FmQ/Q/jJy7Tm/oyj+7bAAtqmKPT/IJZ7+5ZwOuU
NBH430pBSSinuyVV6e+xvw6nUJiST6Jsj5lXuL8qCzMGsphsboIYMfOLQJYciv4m
2ptvUJSDUbm4Thw5ARn12uPqcTeowM4yGN8EFNsqA9GzfZKzqkE+Ia9iPdp6OiDM
QBtQ0t4eXaiue9CliDaWQmIV/UgAYLRbmGsGSt/etLo0dTndWFQHCTH4uOYgRGma
rGxdPXG/n6ttwAl2QRAp8W2niIu6kIvfsbLo0N5/F5s7DjgMZNl4pntOhjqSG8iv
vUpDoCJjHew7YBuaPPzv7jp12hxyN+NGObZ5Lvokbd/8lMZR94V79VWdLcfOFyeY
+9WRM0qluJWIwHZmVJGbUcqGewhNRkp5+CvBkaLSrxezidHf4fJxhs19LYQxCOWd
i/WIVWSQJ4075iwQKtmc7oYxjUl3FAAnClzVG4+bU1+kXW5w20qv6qFa0u8Q00I9
QowVZJbvtEdCHDIONhceKJ+C8NF8bhLXhv6M5r9ZV9PgvnOpqZTyX+265Djd2IkY
2R7XOprtzpQNc8c5j+TK269gv+d7S+PmuUT2whdXPytOn1sY3TBAbYTh9lpZZky0
kX3t0eeOnLDqb8tXyjdPmml4B0/am73VcO/zPfmV46sJS2YeZl0InFcv2uF8PYZt
`protect END_PROTECTED
