`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQir7XEXwIikxLfU2dqwVsLLPO1lj311Q1DVRcRix+L60zigMAinuZA8N/KnhbQv
ZHuty7znv+BuYkXGYOQdb9pobBUeanBZWWtdfFakhbzGvvTgDXjOT/PMqfLA3Tk0
ATdqWwVhVGYwvWRglenJJ2tpahvehGI9RKofGE+pPCnm00C8P40kEM9XcP4A1l85
Q/qvFTN6ZFsisPKuKoovCUbNS9r3SCiqgbE53UyQVQXxUp3IImx3jBjfRXUtuuZq
tfDueY0PVEkCqIYIp5aDj1jOawgCfeaoTS7rL/AuEM42BL5c/KEAF9cSgldDRmkX
b3Ywa4JE9f5u8fknOlemYNlX/zf/0ENwI94y82ZNinKVjQBYZ3nwS5HRDpuMOc9K
43I4y+jCka3PWPhgdojw7g3aN8rNtHuDdMhoB+utmA5IW1a78YIZ5ZKXAbSYB5Ac
MYzRvPDbwqLHURhdR5fPzrNMbhg7YDeYowkXUu1V61s0a9Q83ZpxQWala5wysXE4
ETr7QBKZzCBCRIMSTRZsmhiiXhCwDsq+fbYOo4ve62a/SPKYbc7wVijZVUWiz6Ro
0kAmb3jpqGvdUIXiudlgIrqx68KKgKhO1j0+iFPnk9qB+jh0j2fdjxc0JEMVl1se
DN9z9SqVvizJXhq5DRvN+4ZyiIqRhov9x8MGm5Y3H3t96USwo/2nFHZVYScbn+ue
fmbp+QwVSnJH8XGekVHG3hpqJpQuCLndsEeOio3FHCeiUMkIacFz0W3JPYTGkTJH
KSg2xC/4m5/S64nisEmEh2czi3bxxdslYhLkuABGsGHaC08TvkYPGbWPyZw7G9dw
y6aqLb6p5WkBhJTB6/iXpXgXg5ZaHwnmXLSh/pyyvzdmCIqgOG8J8rBpuG1BD1jN
U7pQIR6QuSSnTbidxWMBkciBIjsKQxKK5OcFxBEMB0gs4QSwjbSBDOWhCRlXsc77
8g+CnfnCPaSUSqcZoxpP+egyhtm/ygAoKqBLYkJlgVRxyPuO4k0emAdMdxP2bQA+
XxORRpmHHRk2tDS15txeoj7f2nDkw2luvNRRTK0c0xPVN0yKU+ois4q4ngoezNKW
jVUePz5/WSQ9jLNT6SITVRpw4x7ODOAhUP8bJQRkbhiLn85WWG/sL79gsJqeEK00
puDwaBBgFolFyhxwllCN8LbxXoCQEYu2quRjVGoj7NLI9UQTjRLZg9Cwzhwkh/a0
F26QHIaCcugoREofrYDXLAEnZYQxxaieUsYgHOsllRo/8Hn6caJPbBgJNp8md2jy
lwTvD1h1EOy6YConuUT0f+/Bceo6ITHSREXnBfxRE/CHLrs+k3wfXOLb0Rwcl/3x
pF/U7FCPfT8jTquY7NoxQT55+tIqtmVcKwBHGQTrvcqlxLZOczc0B/E7OcNCg7U5
agzHUhCzCSduzbbfsieNRt03R9oaH+Qt5Q1SMZtqGfTOHD5ld3rdxL2/YT1FMlXx
UbqJY6RNJCvCVqxtMT5Big==
`protect END_PROTECTED
