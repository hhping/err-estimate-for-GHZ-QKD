`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLNZfu0kQJNA+4h/BDqvrF2LtxWEJNrJ/Fxb8Hjks81IXTiZdlgRXz01K6U/Jw/Y
eWTx7oNywl2GIUEabGoZdmYLnEChF5nO/rT6Li6uU4CeWXy3PmzqyUy7sRI99H0j
c9n4qUhDtmFKsFlXX/UzbK807wFy+/stVG0B6HVgNTT4j7ErfxE+GZe5rwEAbVDY
FZxoMNEMqEFjUqJke99PD4D3PGgkiRTJuYUt9pAirB3qOgAe4snZcpnlPSOfRiXr
iFl29QvSR5xZo1Wk3zB9aSwo4322YfFb5kevsrW0ZCy9NtzQCAVU0+F8Sc8Tm09A
Auj8tFmeH2tWwCgtEVWdMQq5U3nZ6JKLWM7H+g4b/b09wj0vbTY/VO3e2DkMVTy+
04mVt2fBB/nBJrsC+zgRI2xMdwW+YgVQIWt7Y9cEKcXOis1OqwyARn334cObkGP8
ipWcNhYbQRgjt9vjYPut/xryZdgkatQshQX1Peb8VatMQ8JSsCweawEEVl6Q91X5
bG4cpwGdc2Wy/zlJH0UxNoHy0m9p4bA9oCdCVNZZujP5F8aktOukhhzk9GUh64SV
64Pv3XpsVQ/0pktdtWZgtED8qyCyNNara9VP28Ld+X1OZf8v6j0prybw6ty8G/nH
NOItghAL0MnH1a8/jLUA8EY1giSGsVsEYby3KuhgjBU01rLiiv8Qa9/45qeb0ID6
lHD5tM8l4gLIqOWuZdAXy2HDXBE2CmcRBgo99XFhqua7RPfXTH3idx2f/hUOX30u
VQn17Xly6fJ33tMF/wvqRqJx0e0WC1qvb+DIpwdAi589p62ZwEUofFXrXw6Q1o10
E93p/0wuUj6CgYG25A8StQ==
`protect END_PROTECTED
