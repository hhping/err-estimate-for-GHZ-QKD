`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOtLn90nD2sTvRCMpFBpYjhjYyKYPLZB6EOsPgpWQvN09lsEInku7tFCseKzIvV1
hgUIVLsnLEZSV3UdngPaXegXcI+kTzbYtvX1CrlacrtDSOhb3wczg+3cpZdNXbnu
QM6AaMrb5xQ4Tlt5ItaO/eJ+j1q9vKupLEseE4uQfzo72LEBmDCleUg3yOY8e6f6
qxgDpCkee096ZBQaeN/t3Ds0NVxs36c3BPoXnHe+6l38FpC74c0PjXr5ynL7zDp2
u/Vvp12o9JFUPWYhNoEtYQuOiqSgRsH7843x0kanWXRxebCyXXaCG+i8nD9x4KyO
KoNrOMll0UaDSoD5i+rcQRn7Qq3cahVzInyZ4i+qqinLSRItvmZ4BVdlsVY6H+2W
5isj6mrdbn3O99frPNtznCSCPDrdtyvL6+ZT1+scl+qpnzE+uZg+0zaHDJs8eR6Y
rhYUr0d4KuW1taHyTp5kgIygLiqHR9VXq7V60QBv6VyZZjzluLk2p8qn8BAqtNfd
oSedr85X6w5sXf/1Mp+SbN69osWLZgdhP9H4DpNgt7eXJbrSzyih7XyxMZiSOW+/
AzW7hM+0xjLnbHH/GclTE7wtXSkApO5zj2DCMGjuVv22xyCJvIfNdFNWKxy2kKC1
mseSlVZ4gnjCVqetedqiJ+SgKf1YGds70bUiD3yh/MM8S2x+3vgf7ywilQrcJYHp
0JoCmqZIW5pUCyKjJ2U7OjgYCy7YEcU+9NwPmnmMf1sz+DthNGQ1Bj1ASKoQjTgC
fUdUgDfNFOk7TOKY+w0K0lE1LqGjIbxCs/pqFdT5+ANv/VxTSttg5+oHcm8c5UMp
ee1ZEHWebzbv2RSf+yJ/L9Daan7CbV2mfbpYq7gSXi8n4oAjljRKt0pVGqvWe/3o
uKObdngw+PyZUxnqMEl4bEXxKXo6Q/LHr8oC+33eTVnZUO2iUdl5R7ngeM8Ieymh
CUyHEmM0M2E5/Qk3n1xcW2GebVOv6ZOvKmwxJt781ZVC3RHMZowi2dnotZGjwmKW
vMhHPB/o6r8onYebgv6n+vZEUBCh6W2wl8ZORQlZOt1HKKBPCC3N4lFhTxR7N/Wc
Vt9rPUXHnqXsWjUsXZl+jOsdZiNEdUDxDQIZTRNOykXISpWCBKu/y4/cgZ9f5G0E
yQ/7zHi+pRYTWBgw21xLXjIdtNA9zT2DIhe7SmUpGa1YsTBAaXjcHL6/+K9P5h+r
qYx+uO+w+dffzhDEC7IMV4i+qdzPhTStKf5/PdSJjuvT+7nPdrJxLUK0ar5NNRQF
rVhnKgNlKQWFmzJ28UiIKLP/E+XrvnUr6QpYYgD27VxvuC67EzrchzQKaAWbZkra
xfqG99wV5GQhTzXLdElrKr1R5YLsZqUB25ckOOqrAEAn2YSP977ktU7cnXThpxTz
dQrtpvHKdVv/RASqjizGKj115lDDMrBbqkNtkGDDK9F2CMDZ+mm2ov7+orRb48tQ
+EPVQE8a8P9CBSq/fhFQ8e+fYnoIGd1Bhblwg4D6oRhIOzch5t2+Jgfncwfd6s88
OxV15qTbfSkcb7wWG/M8yOWy6BCq2JlZ7bKaXbIGfBf/ImCJphi3OMAF12LZntXL
DHjGKgU3EJ3mS0vHMUMtcCM4BOR/Nacha2LXGHRMazyP7KbzMdt7eW8jzgZFe1at
YA3aLZy9qSob+1DDVUYj6CMVXBKwFZQ0r0JsTCUlg8JggeAVYYCzm8YC1bXOZKLz
i6lRVrMn4FHpl324IgMpZq0GA5ZyV8P+U6fqCd2ClmpDrEqtWFw2yhqbLbI93Ibd
PW3nOO/9OTrjG1A2lEUEu2RN4jE9hGO6mAftprCMaD8Ux+4Dv93uEEsmMWLqk/pH
z01oyLsTK+sbxqHlag0p5eLlm3lTe/LmNGLWu+dDD6d6PhvIlXLt24cVwTc6w0EU
qyH3kIVnsVcKpmx0tlx8YBIMmfAxjBROhm0YRndUAftpGNy/uuMzmo717hxlHaVt
H5O+2K9fNy+3ag/l4T3knG49Z9WiRUC72wJbXXFZra+MQ/v34ChAER9krdlDOqSx
O9Ho74Xd96Oi0xD30C/pJHTOfW45HoDnLpTd8QpTR0P0ymahemW6Lln81IEvii+R
lvHUMjDJ3PcU+Ls3IVRIaDMZsoly0LgJPtPCDiTEe45iCXiUZ4dV3ZxfKPlJYrd0
DcTieVRK0B4FwcX+CeM57kjt3arA+LcpVn2e4F5DCSaYHu3feDWutD/hAcYU2Zd4
3AgdeliRc2YMOWQV3uYVTYTVZHSZndlCzQGipGLyvAGwVWXYxeex8FOn0qN4q4VE
sMyxJX/a3tdRx5dfRTkQ67WDxcGILstnS3baORnOmRRL2WXj1uo23eHo9fakWDh5
8gQSK7EhDyIA2h1qgC5VUvGUkyN64JHX2zL/DH72qJ9J7BoiNeA0JYRvRZL4slT/
WYwr9iKP9BdYpC9TRRetJ6bHf5Hy1z7Twgf1hayp76gY/wSatnGuPzk/9sbUsJFg
waH+I8jRQl+nBVYNb/jRCCWnY++N8aJfi+Z3pTw0dksjd4bHysK1XyLr7VGdW/Pp
zplyvC9I5Oh41a6wyHC5lmQke5pblCFMBwmco4lxwdGLSbEEjOdd46JKtHE5HNPD
RsKg6S5kVzuCBEohaV8/SiRquSXvkIiCX+9aCxUDdurq7+oNhHdKAfo2oRb65rKn
aaXTs0xteL4TMoZqW42lg8WQ+1GAb0NAvDvDcV7IrWT46m1FuYfBH7B5B4nrVafu
X/d9Dt68IIwn0lbYXnjqxjqussGBLT/pZnQR5bzygg4sv4enUSQgNCX2r+xFEigj
NoWYttz2dW1NfMjeGuSqyXMc62kksuYSwNBzHFob0XmdkSSmuTyP3cEz3NI9Ze+o
yKwQexl9w2/CrjZ48wZcYtx58CyceMAypiax/225r3ZP3MNhn36hbq9ViwvLD6u+
HnQ5Wj0rK5wfZQGTA5+0C3hETKC9+ZSjLtgu44nBvq1ZMssEYDwZUVFfVLAdsi5R
37alb8AyMYZzoUBhDnWaixE2M8R13SAo2WrIMp8IJw70Ei23ubE862luexhxHBdT
zMRpq5H9uQnQnV2nHWHHLc+BWWiPup8JC3Z5QC84TEAOfQujs9xQ3G/W4UlC3nDG
qECRoxT6hwHhdCdrUfc54kzhquMhKXDiSRobzaafFECbhVNe77Ucomg0D6LZBjBi
KmxoZIwRZKKcHmJ6kay/RJ9odG6nkLhZYw+bAEGM7Vo1098ILxQsBdxNVZxnjZGX
wxrgGwhqOU/I3GhCDMz/cXkM1P1/EQ0Z73Tz3Hy0VhnRRh4cJ9+k8h0PdjCzpUCJ
DKIMThRYqlMnh5JJi1jQWaCMlZiosZaNDrD5eXx6Ebkc6i6rI+w+QaHCp63bNZXh
mJsv6nATVZtzm4m1c/q1wAKj2r0mk3zpzLlCctUZymqUHuCN9ivkbuBCIZlASBM4
YMlqp7Herw1v9ppjMHD9F5/IkzFl2n/DV7i8gZm/nobJkFU59tQUxhJ+OfPc2ZQX
q1FDI951kOUBpVytcDYZcs+dKjwW0Kn2Anm/Y363yrCdTWMJ5rAJPGXUtKRRXsLT
VjQS7NM5Jwgk4oeud8bU8/GCRaCuGCRcUJK+yS6MuhjXgTrsa4YBeSDsAZibLNTJ
NekXq6KcFeJ1NUeL/Qg1hJI8FxhKgNtdOlTJJPnk9Z8VcO9EzmrUwP078KoS67wO
gj0reOfx1HBMcokH1XaDZQifsC19XkY1t23Yso01oaGo8dWXW5dxOkXz4+vygDpv
TpAAEZVYhwnSa4ZZQlpkxdzUEbJYdClYCfs5950+8oQWlqIRST5bhpGKa9E842Ux
v/C8WfD84sgRqieakkneP750tu6i6aQwPnpOh3oM7Az57gqLEYjcuE8Lgq7sD8rF
IjluMJU1g4KUj0hM5tyGaJ5XEtF1Unhkd5jTScbDQ/6gzK/f9EpKy0qsOHY2gOO2
zD3mMiRZivq34dmSZd0AGEDah5pgWoEUKRXcRl+TI8+H/p44VkC/iL6pGyAA1EhX
tnNAy44vYc/eiJrx7wi1us+80s3JsGVZ91uS9gmAi9N7gPYpH9zYM5FKF/+CoiCn
suQ9LuuTCrhniz7E8bCyx+Jw7FMB5Lm+iOiNt/U2E97iIxNCuEM+vZ/mSkq8Vx4d
p58iRsiCp/gRONEGFcT1ONUEeBPppRg9T8+TtEDkh6OrzrAAbqEbf3PjVZWDBNXa
KL7DXCwFvrASzNVMkJHxKI6CnaLVka+c3a2MPk2lAdKxnmYrDEcn3XiKcaGziCJH
PuTGKyhsA98Y5bQjtqaetoT8XOVQJmH8C4/KHxL1GqQ8d/XQqdIIgK0aNQ/1SuKM
nvOeEGYdqQD8qNF50db3yokoPyqVmYYlNblZD1KaLTFsmULzcS0DWPUPA/QeyE+u
AbQ/YmEvm+nSGN+Wvasyoh+cvrkKzmG7j91XADEyIeDyLJ0+Sk5y1b45PEItkJjt
JKLDylk3iwUt2BhVVaLrZBswiCXoc+VvTqKcQVIgOIjw76cTvpDJLUisNp5YGfSf
G6pg8WSHMrhrk0gUzjRAA5PE/NG7m3Pk1Mdso0g4CVf6bMUnUsIdMWSzb1ff0tm2
Pn5U8gSxH6RvxDt9eN0q/ERSVpsjscdtAwXOriBkEU+VL3A+fCqTjd0f6yVeZQ85
rFh/XVuPXbl3HGmYhRZMJni4eHHJwUQB+DrzO+IdWfbGpBFQrj+LjLrXv6LF1RKJ
xhW7wT+qu6M66PWyItvr/HmffmoA2+hn7fa9/5wlHRlOHVO9ZxhN5Avm1UdbHWZa
UgoawY8f9KGh+Z2e1x+qKFp/eKpcMWW6iNkFPj547ZHvPK0Gxk2NVzci5vGNrN7R
pbhrNP58GxOKQltExh02ThbsSed7Jr+vz6NDeTY+uh3SZG41VRVKzy8PncLZ3GnE
gpV+cS6Pxoo/DAmyL0aerWDmI9rcVsKHr8LkxCX8rnOqCgyOlAcxquWLhFAhwq3R
p8mt2XYlqloMxTbG1gRXRTCtfRs+nMaSOmxwFFb6RGsGrBJoC+JvNPkBYjC6N1Gl
VroeXerycfwnQziHdx9aYzYeZaTxtlh4o3W+M92ku1ohqEkXTLFEfRRM/GU6dtyw
ilckffXmoFXLk4sMImLDcqNlkOAmJ0Lb6FRbTS8eflmZgYNfaLKwfuZ3OQAUcVUv
WCPEzlf5PzdPUL8v6XWXB25L/4sBiK9IeIguYVk0erQQsHneDmdUsQhtieh8JnI0
iMBVwHZNdj34ciT7nUgMSaVlcwB8HKk5vnN03CFS8l8a+bxGTQKe4V0UpNby1upl
LPL6MgdDIb/RbFAOqwhZlN7fybaBKhzuxXYBA88rczGrqw0LTFsM0EMzv/cJHHQV
z+xlmaV7pcF1dGbIHt/fT9GV8J3BK5bsGOmJR8zbF4z0f+M4dTBRmx9tTieMyvi8
m+BBPsB+gBIWLc4MVFBdrwByNy0QOP2WVD2hVFbsS3GEtxCcM8zm0O+tkaFU+Pn8
6l2oJRaNwZo3bhXiJFagLVvo8xo2efjqjVO2gZOKn2+pRY6a4JKoYpZ+TrRhRHRe
vlLi0+x80cZMpGTIPu1Mb/ubOdNdK7/+ltmmH2MWu2f+Imq8p0zlEWB7hCeAs/8E
2VwRlcbo7TihiXZhVCgnDu/SA3CTdicfLXoICwhiNf5w/dsh2gNVh2iHbWPjaLjC
8V/u5tr89mS2qDpvhdluBgPRB14UekSgCCWyK1ThFQtUs3bTue77ntU7XmdoSXeM
BjyXrhy8gzP+yy6dTjVGT698WqCU/Wi/DpecVDzpd4jkrDZwHd/zA70KHBOKuN9W
30a5gs+Y7hvLf+Ahsy6mIEGDbegAdiTraoviekXt4U2OpoGHRkElGV/OPL3sJH9a
zdGAEDEHBU8z8DmZNr/jfjaXBXSbVbPYM9H31vlhZ2dyTOPRKWukHIqXbfVj9u1e
v0JXLN2RjdSuHlgnYAnO+MfqkEQyB+p+9M9CG6ZDwHz5Hm3aVwFWlOmWRbsdoVaK
M1vHChYrV3celVPYusEpPPSfSQvEiwVgrfeBw7I8oyB9fl5xd0jDqClNhgac+jYi
Y2TQQtyJ0cp21pZ5C8gLz/Cyg2QMuMQYxRJ+7kIs89oTW/XwvcfL8ZSqUNzhMke7
C3dshipGzozrtd1jYsu3sV34PFXZGqKiZlxGBQajn/kb7Sfw0h0BuNwbq/+4/IIH
/b0Q8HGg3iMhtuBwtGkddFxz6lKOzhl0ji9fgdmeU4qK6KzyRnSTGuOQpFNQqwXG
/vt5jOsqhHjbJFP5OM4q4chkMd2FbGmNNGXGtZY5od086bRBhz6i7HHjkT+7RGYQ
nsEmY8LxbwiITmpov1M+oyX0Fcvr6ptsK14bR6nDX37SVc09WYfJeavFyAUaDG30
89LbR08HAcTj76ZeqDZKSzZeOekXExLlSZvBs0Nb+8BlisVqClTJt2rEUBBzt2g2
ukFbBKlix2TNuXEajoL6BHez9WNL3cU+ZI6Sc26GZhFIlic4YTQnRZVx/IqPW4f0
if5Lhbn/u/oul0/YPb11a7dJXKuC9NnjT89NQ/IvX1Ibs70lcJejbGoRY48FHJHG
cKquURMiEfc2bti+iGs/ntmOeZRTACT+NV7wF2wcWIlk/FZWCOwfvqS8iTYOGScQ
/WhKbzebnwpwDDNA0gL+ZtqcabbPn+6asMEjGd7p/AAJWgEDjU+aeoDawGPD2mTz
eleiObbXDknZKrqaNuceqjvbvOYzpOFu1jJvQZK9dyz9zkZvHqghzp3kWrJ/wVNR
S5836k/IqIcv+ie1hqyWGtVd2YAHFPm1CJ1PL6wuENRoI+qpqCW9mxgOQzQ1XAyq
99IJtSFI1iCPg2ohHVxSDzoOTGJyIzjuNet/xYA7AoG818M2tD0qVX8Rv0HzJeH/
sSM4tuB27ivhL0jBoWQ+ECT6KI88Dt4w+LSPpjOvEkMI6OgpYKDm9/OdpZHP8zbW
EzW5KqMJniincZRFrM1hmnHXg5PdPX/LgUiNcoSJx+VQg2SbNGUdtl0Zk/IH3y54
4uBBrsInOdsiWzeb5ja2YNTxLy5WDrwLayfE9WjgLDYdKslD+3AFvYt+OggkJtFb
8u1OsYxPzbQ/nudwfXzC3GnxUwdLyoSH5reWwGrXnBE/4uX2MyqNAJjBeAvjLwGH
eeXcnBPxjDXUzKfMRJ5B6mMqiaA+n/T6C3tdkAQxOR4rufIEHKFgAsrNYaH+9XNy
WmBw90E0glOOp+YLzwvS8a9Jscfc3RbnUh8GzTRx5+8sdQRz7FrvkX4YDo2BkOYb
4oPbYC9Wc2fVrZ5DFrdH4hX1VN1WgcNDpWT/aJ/V7eHSbKm8VgW2Y4daoKXpMPfV
Jp1FSQOm2Dmk60gM3PvrYqhxaftmhIXDH5M+GiIKdovyytTi4kRN6dL0csAkCY1a
uCh4WvHyiR9Mi5EOSnjfxntGlALk2KgksZGTEpnFyFLxWTExz0ig6gHjqqX1q3Vg
8EC0MbX4YNoqZ1bFkdYS6eMKP5yyvSVAZIreOUgJBvobjUUcKnSy8RvWVp9BzB80
YddQyboDc1vW3Pp8rYZxu8XrkX2JE/E4iv78TuEf4dYU0o31QFjMDpfzS+I18FvU
YS0eJBY9W6kcYBXeo8HUIUlS4+rosGigSZYGiVO8DEmXT8B6ar6xmbtVL2gSxt4F
NJK2nGg3zLGYkgU0CQdad4eo15upWt+uWSg16fPD2nspCrkuLF3MZ9I66ukdSWld
V73iggQvoVm3FItcecS2hC520aIODLccKHbt/kXKOmyGKoNCOuAVGUZnzgQSTdck
NzphKbqwLJhghJEDiH5s2lkYT9HuJ0XTHB0laAoKsNb+1KxnMTwdvuO0X6e+pGEX
8r+Hmrp+Lcl0D1MtJ0wgIP2ha4StVpTv2t+tjXMGU78ikjjTABnB6ncvruMOhTrf
d7M2disrIF3rXBqsy7YcJr7MHpwaAtkGBD1pXp1wP+17mUTunpXPZVfwk5b0O9Ex
OP1ylLKINl6RspxMaR1hMlBQXmPdmKTzKBy7ZUu9BBdKVVO2/b55GEbjPk6Vptot
akZ6rRk4ZIlQdAQLiWIlRvtYEdVpOiFkTb5yd0BmI5gpyT3q13YCD69Uzabw/+UE
nql2Bi5sjmtGfrguNmO8NmjhgCHrkqPqjrV0d3n1/XCB+Gj6UT3vPtWDAs38Sl7s
oQvODbm+rCNMVb6GtbpwGLQ1lT3rBf6k3NXYeiMk0Dwlra0dALnGlTBCfsZJ6E3p
EVlJD/k+O26kXBTnz7apej4y4ADZB3IZjI+8X2Fj07IzVO79ZT5QDwlyyp2oXCNo
ae/9QPROfHgd+k7pG9zOVwdyfe2pC6el37RX+X5BJuAhXyoii9wxLUvJycdqJLcD
GiAU+xTy9BTaW4qoXL+YgjtQq0H3HZIP+7wck+i74MCwEpzMHXFEwJpvRSgRuObh
KuhfH5u2dbiAcSi01SaKFO4rV+2K/FL6kcgPP1IF31f9djziFuEA7Bm1xqEYi227
kheilVwF6yQ4cemuqM5cBcAIaqDEq6b4UGjiOs3X7RzUuIbNLqkV4Pw7G/bQW5c0
/NNLplPmosfrHhbSzCVj2DQDMcUu1auQnupITdo1I1LVD/DE3SIsHThgdtpPr/OE
7YH9hCceXGri4MGtDrm4INlYbGKinY7IsMtnS5P3plpO5GGWpgPUxZ7beE69xdHg
vRBi1wgCcTY6FW5rUGyv/Uu2327HWplvlo78fXYqujrEABzVwZpUUp7CXYKmft5Q
MHOf0ZO713zWFpemxfPkCmct2JgAmtyWrHWrQJmfGtGVu7DjrPvt05FS4RKayH7D
xw1hfdNHRT8tkeOf1gJC/+3B1wYZGP+Q4UzazjXUKLhYWRFZsKXNq/3azs2db7kI
qM3QyTngh2Nvr8ayXTym2ckRd86WsKvFbZb6XplYXJPfGZNoXOjDsWkOB8jLP57I
GOhnRObCIg9lk0ctrWpF+rxvTHVpJvgvVgxTLVUaT2+aFgW3jIrNwZju/cVP6ar2
KBazG52qEyh298DIUgAtQziZZwZQsX6Br3fmBjN52m07bSvNOkqK8HkZip8VW3ro
ROOKwes6Y4y0cIpGLIvaBbZCGVHXc4outsGg96wnbsc5GNFdxnQ4JINQN7iBbJqp
IGpQUW8XjzIsdO2y7bqbZzx4y5hOpqRIWKaFIONPcC01OXrDvAzb1kYrQYAdZduX
FO6zvn+BWcv3VxF+yFoY64IuvGwnF3f4Wae1AlTPjsvWyXmawibJD1A8qP9nNAW5
USBWZlrVR3wb4RATOuKEzPrWM9p9SVPJCAPyfcLnUebAdXqmU14eGmrjD17woNfu
puDEC9t9HFqiHdZ/nwAqDsAF0mTiByyveiWsRQpGee5XjnjAVRZlJHbAz4rJGGKs
e9U+R05AAT8TBIBRPkEkPUqdsU8D6+xQtc6S/FJirZPljgGxgbiPWdxSd9Oc+UmG
X0geq54ddcwejeBrYjiqSlBId1Yhmz+gGuVYMXVqBIp0mdTrqF+/jYMDI3Ow1fdt
0X6T6SfYgWZ3mRv5LBsyL2ktnUP5Ka9meRlM/tk9btm0iOSczWurOlaSo2zp5Emu
yFpb2U2lfLQMWNBZMuvK0VihAqqc/y4EYQIO/zqmfIXM99H6EM/Kx5X0rUXDMeJz
XmWTEvA8ms+tohomizPVzPTI9PXi09+kamIYyYnN0sxUARLmkZPJ6BIRc1By6ICn
2Po8DClVOfZWl7bARV5NSYRYe/xrKxGT0RSnpWqF0sDb13CggqEAZHGulKK/iBUd
YvVtp8T+XmhY1PLFw8TYD96uwi4OPDTejrRQRNg//xQ4wWGxqPoEBr8wBCMjtdwe
5xL3UBOadIB4nEagcO+VWHns1vknt3GUGlbXdDGbg4Wo8+udmGWpMeDAY7TImrIT
KEnz27ya8hQnC/qIEjihQ1Xw9mJz6bxBvP5Uq+bum8CevmRZExUP7PIRpCpS14NE
lW7nDXl+eoHT2PWfgmKVCi5XPHM3qTdX4MFQ5tJeuOgN2DZWv2o7cdtl+Z8gZ7w4
MF+IZgAJao33p2DEy+IV1FIgsZauWGOMu5M8LrdKr1BdsJbOXACI2KbSYiIS6Mze
PsaERNceScnS3L1A83eC46ZUlJevXiHr9aRw8kGapqejkm/264e4otEs7Rm8Ev8l
rMl9V0LxaOgQWdnEI5J7poTR/Mi1IHBR3sINu3cvLsKLhyP0M0PKocXl5qHU1VVt
wXJZk3A+tfT0Ss/RZO/MFuU1QHM1zevmdn3UvK/VKwWn7b3YjkjTeBYPFR1qp0D7
wQNaSUZ073KaVD+c3cWLWaaP7iBIhxFlmB3IVbGyQuS+ZG3XmoExHqRAv3m1LhAN
bUOKWdvfZJTAqnuuSHlcjMvDwmZQ/HdywjnVGnIGSVg/csoPY063CITdTOzS1Wbc
vBuLaYjZsc0aVR52434Osfj6Tw/dIYa9tFMioY77igijmoeztjCYcR3wG4lJwV9c
cc6gOL2I9obXmq71jKfq7TqGDN0bkHnfMumbhgWqVU2N0YlzI0CvFkDo9u0n/3IM
ADbe/SVOEaOYmFlMtUv6gD13fByXfgIH+hJ5gD1DDizXuJlQJvrU/glGN5giYeBw
rrz0cGB/3xMjsD7Kg19JbM3YkjSgAbYH+Bhxy/YZeH36ZMp9v+phgkT/RAvS9jJq
3xoZrnO4mbU0XC8DO1cpMh0mHPLgqhh1owDQRVq5fS057P2nu6ya4ExI54kvP9at
4Xy3g14YDECDR84Ies+TVkSJszbK3ZGOPYXqkrJD1GHIOWDYYhAILx6sM+8j7afX
vZ6uzEe2QPUrOfPRxeF82hSfUwHgkdFGtARgetHaYPKuKRwP7c82WFkkKUgK3SOX
p0RvM8b0hBwTfc9QCsN2NxFpgf3wDQVyQD/AQPYI9tFi1HHcFbz8dvnoQg98gtoV
wGSf7rYKvK3EazDxxx0iWgh0p/JDldd3JG2bgx/7A7qY4109sOVHmAnbDxOoHzD0
mEp4TnQyi2si1zXDFKt0VaFNVpaNZ9YmPwdsEwmq5wN75K4x7x1EHtqe7oewrICK
+1r+Dbml3KG1a5l7SiQd+g/ZOHSSjgLBNgeLWvppvz8pNs+mn/a26+sHdekhD6wB
r3mdnViKb04VsViSqfmpbAXysYSKuokY+xnbsvUMr/0YCDegHPc2XZjXoaGfJJsN
W5+NMnXaY+fcUmfKh3MTv7EUyJhiYhfM4Q5AJyS+zbpse8dNJeG4ddpPFtD1N6OY
mRmxaXOvbR2XXsoSgWhDByaG05dZha3+PuGUSU766C5su6m8JPrHCY5fn61lXxUN
u8aUfafmdkiILu+W5GMCq19obK77qpf9OCrSBsL8GoH6YDpgFuyIbVShErKQKty+
2QTUlwY1ajnYvq5uYqJbmWX30tjMCOzJjkuhpxNRfNcp/fl6czDLSbyV2+yDGfFw
XSxbxBkXXm1XVMg5xDWF0esIWW1f2BgLqlwM3kzqa3xqMbhVSpkNkAMG6m6BZ7iu
YX4K0uG08baPiAfV00hbEJiXi1SofgwY+q+6GQnrY6t3AakWmhbah9ZrGgsICmUN
QIwThBsYqHqQSZrU0IVUArsFb1gbBMrEJaes6NdaDhKaTvoi6ALI1j7nqZ1CazqQ
adMH4XWVxecp5jAgtHimboo4jw4Hi/w2htq2anixEnKvRVXhqtlmn0JTibpRAnxs
sJswIoe6hJqMdILVXYLfLT+GvbJ9wiojwpDjcsqwqEs8YrpiZd1/pLdULmITPEdy
EM/Vgt4EYAXLE9dyjPIEwMqxMwpRoxolq3yaz/7FZD/Etlr0TcOobIDVczAzTSv8
UJCeyuUnqx4o9yCB1XEjSgjvlb8VR7reViBAl0UzHFO//LYriLvmUGb50iwWCQ53
Vi92NuqJMNV6t2nomy9lpLzp9/MnXgWFMSaakhF2RQKwlS48xG87CtAR6oaqAIlM
xbMSM7/2lUV+U1i1knXGNPMQOBw3UxY2/FEoPYHzB+XOqgunyQY/WYi3YLjlNcoH
dHhl1F2t/exywnvC+S0QpRwEOtRUk3qQuc0KHY88A+mELgA+Z6KI0M9TbBAL/aek
GRjwYpWyPZrCp6vHsrj1YYSVRACLTgImQqHBMnSWqA7HdaY5nTubvQSMtUl5kG4S
K5fLgPjJZa7QKAJrrjtttOMtHrtnJOpYdpJ9bI4329sGI2Pi+Fwtbh0cUozWLSqI
QJAYUn3Xai/1K3yJyi4RFfubCcgkClctv6Bw5x8Za7oUeFGCmcU0j35GTfRRYkjv
NsXY+LEmruKQ3u2oRORcchzpenPTTjLm/AKvJKnFJpx8nmBgssK28XvLkC4rkbZr
bh0RN3hLUctgckv4xHAxJ1CgQYsePe1jECq/HohqlKQdLCsBi31qzP/QOMBqKbcw
x/2p/XNGsb4THgNSbeQjAPnKp6X2I3XXEneWGW/pxUzejljnFbGpJ+IrTQ0+j+KS
+0WxNldiajot74gXRwNB0uSe018bePoc8UPymDNzY/dpZbp9YwNwGdN7DHgFKx4p
q4ty+OcB+XZN9lHXNY0HBmkGLhqMUGiJegvEBKHDA5FkwZktOPMb36zsgz3tWNty
c9uYA8NNASLvSO80AQxYACGXzwtYoJdWGSWQwST5VFsTf7meEJ69Vv+EvZ4AEZpF
R16yK5TMwTg3+tcClV5E2Snqtttf15H1xXhVnghOau2nLd0/FrhlowrmpMzfko7l
rY0Pp6Q/V6y49030uaeRafCn41kgDP5drK96TF3TnOrfYyEEtiIyyoJx1LcvatYW
aJcxUqm2cRMbOjBHqgZ3fdbgS1Js0Rs9iUupILxaiZz+qxz2+vUOpJPBeJtBm5Eh
Z5R2hmwbh8KlxSJX4qstXTlSmKIJB9BICD7RGZkKoJwBU+5UdopVuZD2EQFrNCfK
TNOqGzO4P7cvcREj0a44eAQgHUxGu4u91a1lxbSf/RSRfa+jXfiobMtCdnYEsIx0
9dHM6SxH4KnhE+syv28GVrTt5UzWvfa6BFvu4EnrNy2MuyUL3j9N0G1DoQ7kd3AQ
rwyyMTPrmXIpGpriKjfsDVIyLWCIkSJIsItrE1mRb2m8qWY1YAv3NXbPH8w8rIyY
VCc/vJGSH2U/itPQGb2QaaPyaHFvojSzj+phMsFN1EOrS9uZlLxe5C4+4aVcX7gE
rop+GKNeTK0iG43copaBzBk+JogyQQy3XcoPb77tzPfYbFLcr4K/ARcwTthjJlZT
pHSuA73nKQL3EFZcktGlddeunXsL8LAO6HQ74WNFqY/z7HO9YRA0DF6Q4dXJskoQ
c5X7KnCl0dv9qZl0OxDlQCc9u/RlFEHBx8cEYLn4NN8fz7TN9mfGwYHy7Nnb2/8d
uX5O2Z75l9qPCalZWG4l7vbICmeEF8KXObeICDctbYjrUEam/xe9HVJ08UUENoht
y+bohfg/PBaB86YfUsHWr0RK5fykilV8WkmXD7uxVZk2v1P4PT+YZRXE/u3t5F5r
Sh5wtFbFOI3GyXS4aKP5Sk1dxCcbwF4+GH/KmB+RrdHl3A3bSjt0PwFhntQUznyU
mpEjTEuo48AxfiXHNLCFSOpqDWqnFhgiZVwHloFKlKHE1QcZzNtMUL0cbmhC6/dn
H5sAuza2pCWC4t8AbC2l6IxiwtYgavNKBYxADMCwYzv8sLolVZU4QNsBST9dsJZ9
cjFDNsOVUakXPtAVpml1SMWXW1xeABU9z8gSSJKfHNR4/Wqv/RXjLJHcQBkQ6oBW
mcb7uKg5R8p1xWIONS8aqfn2AI+ghRsotogKh5N3hfOabplXKX3xUUfjOQJrN8LN
igDiZ1RfJGEmCOZIjpAG93J+Kesh2Z0UsKAvo+qGujfN0+6rRQjNuMgwE+RyCIJA
MxG95tN+R4LmE83rKjf5+ugwUN3wExrmfn/jP65vKUwHVzaursrV5TO41dwIQ1WS
Il7w+mqvq49wXdyDAC20t0L2LI37GqQ4OQcUpYtX1Gg73whj2zsJYpPkk4rBpkIM
mwuaWNTqDPnsk2pNCgPK1kENOjf3eMctvUg/7MvlTkSebHhf2N9yEbdsw2G3ln/0
qYX8hNM5EKsnekbO1Zl6j0I8T9vVJEyoP4Lp52C4oxBqoCKZqid4CjPtigudpYHJ
osCLG9ZHy5E55kyTaE7rRQbfkZNuI/600ORqUpO1AVGzo2F26mqTtM3QJJKVOlBH
fCXOFhcJnHPqMx8hgkkTGCGyHaGiAuUNDVsTC/2O2mzR+aRcD3z6F3poMKpbrBND
BmrWlIFwdzVwmGMThm8q96nSQNbEvl5Hy/HnAHrfHwRhAmjajyFnR4uHvFdConPj
Ij/KX/HMcdVze2OF2O3Cny4q4B1RS25at1jqWcdsOPWAmr6Eh26dve68hgdlvD3I
6IJ1uDGbwBs8Wsf1Xrynv3h1lSJuqiE0mrNvZBNvgwtqL6vbH9w8tfykO15LCjGD
xMdVbHkSc5fst1E/cXQui9b15O47h51xSyvEz7UcssqwyoCCzkMJQ54RGrLU7uLj
BcU+4ILamJgj1qwbVRMQg1X+/rJ0vea7QtQiZqmh0+c98oVRPjmAg25MVcJFoMR1
hc93QvbdG6tdkhbJifkNXTEDR2tAYl/jvF8CMhXfkGgb//haqzZ2F7+/b8E2zCVQ
vVSapDS5F5Vu2ADldQsfbZko9DCip3rPXq0u8BYxmpJpZmnK2El/g3Lxfk1oA/AV
lPprRHc+anPvaQUScAIrtVH8jg3QttkiqyYRZaa8c4vuMWUbYfES4RyUsfyeMhnG
LYkn4RP7f4mVyjX1Vsj+9h7G8VD64XlhwEQrnxD8WG0JSxSqLB5Rk1sj+l6QnO1S
QXE/7N3bCYUSJpgnRmQ0oRubjucEPmCBcYe6/fOa1GsQ1hX7aHHyI0BDfqLYRw8J
MsCKQL21G2mZe0shVgjtOBnGfqERaG5kYiiS/q8xULi89Z8R6lNqqhYKRg9FRJeP
+MPaanKKh5fyEBj5IgE/AmH6enk5v7V0G0MraUddXtSBAg198wrMcPl+46xr79ua
eOR6Tjy55pFynwMPuln6zC3qKPSvtP/qPKUQ5OCqQn+k0UTh0Y9ZfSTjEhJ0do1S
jPz17xKRSDG+T8GicBYdhm4G9HvKstsyhNGB3HvJvRljg/62/htzi7iEG3+Kr8xp
htruWlhZaJzddCQnGqvBevQr8OZmVQL5rWge6y9AOnUC8fiqo6NRS45bWtDauGOr
ufNlMZcpfBo4pCHZuiGl2PDZhdMtJ/+FvUgrjeHQ1NvlYB2hobmvYi6+25S+keKQ
0UN47+7ww/YWb4tC1U3Ttkz8ZlBe7Ddyj8VoVaa7zxpEXsE9qHgrDDBLjBT1MCsx
0Z5WvsQIn1ujkMsPRvwRgWc27iJ/yy6Kp1wXpwMFOui2YicoNoQZAt96uqvrFJl0
YG0SFdCZybhpQVVAk+j1Sa7uXDTwgZREsw0HYalLBpEN78wJ8XVwLx/Iq2AUQQuy
WM9j37fzIRVCCxSsHVKYhxDYdwweG8tIgSmkRjHTEEGpRDkr9yKhvCDwaWR6gp4+
xprr78doqQibk+XfNxij6D9XTgbEX2eMkQWiOr4RWOdxb/LL5pndvii6qk30Kk8f
oR7XO0VnGmgNM8a8MUorfMJHwLv/4j/B/+I+CbOX8OKPTlKBYw1OEdgkKFXA9ypX
DLh2rCNmQiCd1OD9Imq/Rvnqh1Uhbku7Q+XsgpWKGHgm3AHIOq1X0oPJwNRtZvR3
9q5K+d8x2EVgUOU7IJpX5HYdWx0hfwzlhT7OaoHernKB20kEkSRMKmWps51vtiMM
WkmAPlmiV8TwaXZ/1Q/eeQ+c7yAnmBaPXaMDSTAzKpyXJNB0bnVPBDaa4ObYc+Pj
ZGMSTk2OR4UwlfF2lZO1zTpau8RnHrw5EyZSVCOLYOMGJbpVoyxOwhKEv/k5CPYc
okJcA1k6fi9RQp1dQHZ9uhu/3AbSUBQf9mP8OwpOTJBkC6d1vAommtLQ54YFxXlU
z/u0976e3y3Y2GFLlBDqUqvieZT1TBBqevRvXmnUFLBfYsOQhif5mr8b9kVAsRei
qoBmffDVnaP/eEgPMpILBrHgwreZ4rlDatUK5FB+1ygNYfnIuHNItNYmcvTaa9P2
A2SAqW0/PkqQnSLFEHB/BnI3aHFTOIrzUAoqmgk/PPT0BR2xTsRbfbQ3WYxBBkhu
m+BjJDb2xQuF8eLf6nOqcaNaoNmBUCja98z8iHSwd+E80A23xxeKnYKQwJSTFCxR
k7TX0M2jSGR4SIKnx7EsWP1Yh7AOq9VQJQl7PaCKSZtFTiZ/blNXjWD0ZsVz3aKX
Y5HrVrE3GuEPGWmP7xfQRz1ZO34YxSC/yZFaD3H5y4NElEzdWw2LICgTVh3n3wty
srX7t3G32H8Ypiepx0EYVs+eqrhL304k4ttGhr7PFdxguvCfkL9PVODew290bwdi
WKAD2WkzlhCRuU6CXbsOq8ZxyIf82MOEc6iYJqLolvPjmQLLRyLwvXh6EUfBNgnW
zxSX6GYswhnfgOi21dhzHJstaMx14QU3ImFxZg3OnNnmrGeRmUvzsiBUgXdEQLXR
8VkdRjteI+kxkj7bqu7/PfS2InhOvGTzlPFWsXoJ5EOUV2Vhb5oAgX+0MPFMTsGH
NrpvsBcHR9/AXPUPJAmpMCvBS7nEjqCqoV8TSdL9GReGos2Q3Lfaivlxhzq+Tcz3
Vh2JeXId/GkdvSlOxObgFwu19nsTupqWcu+BwNktbMA3bta/g7dxlwRVU9O0V6Nv
AMVdt5jKoEbPk+ay/kdzj8ZgYLY3x6mhvkgKogptlY51YAmFf0mqkbf7Oc6ux7Yp
+00LO4dqMBMZ9kf6vwWfkcN5hq3CWCSTZHfcr/4DBB3pyTftiz3xBrtkQxEM9GE9
14LjbUMyzEnxenGIEEdO9wpXGVKN/JQGSBI8Yp4adAfUZWxUZDpI2sC/Rk0oi6HU
GmNjXyvp04Gh4hs5AOE6eX6Jg2YMc9OB3FOTjF+NFumUWLiFjmMIAGK5jqbINYdM
itLDsc9M3iP+6q7RmlWYdoaraK70cvaSPlP2M2aZPo4ifFke5rzqlfNysO3c9zcj
7dKc8Cmh627/+XxPTZ9hRV2kJJg0+nhe6wBhI2fgmy4GZ4sJN5/hMbn7dc/D9Vbw
+/6es90EWF7UN5u5Gj4Fm5lhIZ8tsWWzdX/2LR0sMOCoz83BYhFZMuCtmOZ+BFRn
fW6lQxzbV+3EEOJF6NRnBv3DLGJ2zvkIs4cwegVqqQMQw5byyQyLLjgI+YgCXwBd
JKUV5NCBYp2bjD8CUAz/xnz99UN+RViUTz7R8mah1ROyLJeb/lV3C0U61/9/DWtX
2odAvwypylsQwG2m9znbi0dmO8i3S3yToq2WC9HkBXLeZkvh5HJOY+e7Z0LykWZ5
v084+B0+ZBuFd+32tT1Vh4JMNGAM9DHeKXoZlvwEEZJmQ0z8/CndQuxvD4Iw0e9Z
2LzAsuqaxtkY3M6++eUBJIphknSPdKwO/iIe0xCHLKHnP1Ho7WyHD+bweTDSbmw0
4I35yAG09gnZcvHH6fqIj4eAF/od6gN0QNkqxiiF9DeE+UxG/b2aRUtFWpUNiRu+
GxEo8omQrcuf7qSWLFhWi3xyxdyoGo3+Gh0d49cFtbyZAEZ0IRTbTVA14OlWjiT2
moUWlWNaNIQZsItblKHTFLPqfxlZEVaGhVVEFc7/IeH5Znksj0AG7uVVdnvPe4aF
ZP7NIpo8hMMTBTkSChGbVu6/O9zdhJ3t07SRxOtIJ7BN8mX/uaIgLeJcGi8Ez6ug
GLw4ThIH47xtuje1K7aLCujVaQDvsPPT4v+5BhynswTofrJaElv8t1JPAXjFa2jU
ZLtIN8ACxqWs4sY+uv2XhmzxGiXWUMs56VVZLQ3IaTMKAeBdT2nen6WlsJG8hGM7
hbwD3CfdOdlU9rQpuEKMVTKK3a/dxHemPZRPl/2duKBEduFEKMv9i4O1EjxqBUzV
bJVsVIAybC4THBMLYlUujxrtPRYzNx2v107NmdsmtDhHj8SRIuR/qaBxfB8KPXjy
v9osjS+YWiHsX2c7m8jsXxyn57wrcqmWG3U52qASnjQqwa+GBjoKzt02fP+7sKk/
hCpnVPM5CnxekQDFNxYuyJwJXR+Z7YPVaR73gh2usG2U0KycuT6FCFVPG74xZHj2
+MnYgDR+RAFvykMCjuCyGzJcKDvJl33vEs5uMvXAga6PNDzq/qds51P5dIX/ph4t
l7y4piYqmtP9GZSq8cKWcGq51N2io0LkpQLCrA1+MEimUPXeAFtrMfooRrUGGWX5
qT7yfZYoN9xPfnhQX4NrbBTOg5Dnc2aQLUOxUol/BHbd4zC4QtLMQQ+SvMFlrz/y
A5ZPSeZhSyP/CY6ymbTytzOrMyybmZQWHRLOYVCZwq47daClGqFmhgBjYLKYxdpF
8v3FvV7Pr2WSVtcfIeB7RR2PN4IclL/30GFarCVQMOV8ulU0CIb1u0oIXFEC7eza
r+xjRQJc70A7Jkdsso7sJnIkpsHN8bO9X/1uvVJM1mUC9uwvjfUqmlRaP1YL8USN
1WBGt98XFxE6tvcIJ2jysvznW6AKJA27s6eLQ1R1l7FCMUJOKXiiKfPnk39mycKg
uUcHSVLPCIt1Or6pXu0p+KAKZMtOs/V3sir3IAoRXUOLwLECGsltrPXsDzSNHdvb
MuoklxQ6sop25kVcQ83PRClPto1NyrbPtEygtvTbwb0E5xYPfZYxzFo4uWDXzUL3
Mp1nccuDeK5jjRfQmhchnYw34y0VGqILvrs3BgmCCL4+Hb48ugRg6VsolevQBR75
P1txUPsNBoPtzoj1GnFfyjNFAqbJcaYlqvvWw1LobO25uiwe5irLcHaKkKcet0tR
zWg4KgcnEHZ0Avvi71smwV56bOcymui7h9yoowJMAYVHCKE+RKvHGycKi3o1x2WD
D80NmQkjQb1lXDg1XydnLSBM8GmLBR8AKGKRI7f6rXJV2827DfW97JCl3lTwDLGB
6/D6vzXlL13ZkjTNjdIbJtONsov7e7hFUw9UOblm2C2XFkbD/ciRh2Z6aFeVevJn
AsgCiX79JVMvyBXon9Geo8I8A9+7DfpX3T61EVh/dWRFFBVENZOX4bBkKA0Z3Br0
J+P+ETanzDpPGaFLtSYdr4ufhNANg4zpJ4iY1lNMX/RnWo0ANm98gl7N1dKn7fk4
zfSXE0yBKckU5yBykul8zOV3g0dkf34PddYmwtwrNmTfyhv0qpCRLNAJyugU4Oc5
wVzNFO9MAyYdZ2G6ycrygUsfYo2PhxdZqpZAygubyKFKcGMjqUmAS9Z73olU0Ggp
8IFW+ssljbkXdbfV3/uMm/7gyc7fLjhogoRS0UWzXN06bo/s0KMSi2ds0gFVuS13
bDJ2ctvCyh8j3fcTN2iY4YJwecn/7lrFMxhpH5M8Jmeisw5pweA2V/qgQrFSxOTH
s1oUPrk3UnXQeYr9bZxPXVqLUCp7aXsDEQr/0pA4GNsYxG3Ee/iQ2HeLZSQYFlL4
n6lWBoZyINPt0eOKz0lPZYw4/xzZnAXD4qkb/nbgEOEnTXyqFYieeQ/EQ7bqJX6w
NGeS7j17Xn5fhze/8r691QhPzTiOAYEejRr+Kx76EulhbR6F1ElQpKD+Igo28u9b
XUhPJlkicgmQKXUQftE6UpvyiKpXKSIddEoiVLxX64mde6UzcVL4+1ldWBO1apT9
jjqHt4R025MhobHMvfIiHn0C+hiIFHxJaZfJqPYomidjJXrrAlkXOvYKeT5eIP7f
rLgrNUWkeczq6D0NzzdU/wQhqEtfBedypxPBtI5QhHjoGIc6JVIvZhxsgxZV5I22
KKukVUAl9LncFghMxR6fnduQsoM3l0Lm32ARdg0NOsPLY+sjhnY0T9I4DRcmKfmW
rsUsnfv8Z7RhHttOH7YKi+4ML8rVRWWg03B6Utct5Thn3xhhQOnnqX/poiJnfM+1
76jLnLOKUB8TW5njKsAdx99bz9Kr6d4rndwdCeSpBoBezCYn2VLrKT7pf2lqnq5P
QUud2iGQrdEcM1qrAS/iks+MRnR249iW4G6eUsutZ65TA+wXxB1POjGS3JKtVSHS
PhEc1j/+CDemUagEzhNvQoVTp2ou8lgwDDJxoZLwWrlSvkpb40GWe0iSMRxvCUM0
F+FOqD2BF0qkvOC2QnfM/zRE88UQ0Gbh/WbroAyl1KtajJSOEhy7zK0qOz2gc4zC
KWVf1YBn4XcXOQ+R/uUWHoJOxUS6sHlOk/W1P1Dn899QuZDZ2fr9af88tAeDVolv
3QzYS4pOnw5nIEzBVrQ0QNwgEOq4NgCjym4sHcdvidgPbxu77Sh7fWAmmc1JLP2N
3WaH9ggvIpLmeKrf3pwDuApy5IxJhQNxsaA1PeKFaRql3BzzMO0QeTM+BD8l1hNa
phiIUKEfITB9NLxaNiuQjSCD0BgwXfoR3bBuZ0lehTvuQSiUMKcm6j7rp58baiYN
o5B1nUg8RSX0B6Nfh9FSfU4ZY6epjfby5KY5nx20NleOov3P6CCSRNS1DKiTPOMQ
G7oY4ssHV/RxtdHdNFaKBIGBz3ELR5kNM1k2gjlzMllhTgEHP0LZtIgd8MxCD6RS
QwnS5Qiadn9PieDvDi6S4pkVXXLwa1G52kz1mV2TvytpzvT0iL8xJjUGJ/uEiuZ6
hdoA01ddphaRzZeWkmwmD3JN6TzbGvCN4H8saYCe66swRpOzUL/AkhU1h02aDr08
OK77CnQbTMpBkptl3Qeu4miwwM/5BcM4crM8S8hVfrCVAj7zB/wQ6UkzFoCH885m
u5sUWLZx4XgUgyGINDSMQdQT47OE9Bks10YSghSYiZHNoWPSr6YrM73NA1+hC+GH
Tqk9rpSxCZhh59nqs5SGmqARMDqokVJNu7sSfxdvMKyWbCIS/c8K3zLdN/MznIgi
Gt+eqBdT2asBsRy2YYXs9SRcs8SujaJL9khlt8XuNKTLfHIC0JqSYeFRNOpmg1Fp
Eu6WB2RysZxsxNy78/2oqtA8EQdy2ClUOce6js/BQBHnLnQz9w+c41UUK1DW63ZX
Z3maBjlCQTyymkEXYwR8eqmWgFVX5ho58Hr7lOOsRPkoRMoSFa6Yf//GvhH/7dMI
vCllq+WT33vlxJu3ns5w78jBCqVtkc1ZxbLOcBOJwjBKyrZJfZ7qNAGZA+VjRHfG
feeiTxy+m82C5eybElX6pH0m59nlnbKtoX3bj7XdkHlhc2wiI4qcjdEmaD6xOmyW
iV3QhjQI1OWMT4ZKX1vgoc19wolP5XpiSdnjANQ+Jfwvb2uk9rAJ7g+7qeGXLs6q
K7Hq9hETUEkZIcLF2v9PRaV+ibnCZqSjw89pcxXV2HCLCoRbab4/2l4EEgqtOBvL
sk+2St1fT5sxUS6kdhb3xYqhagUsJ/LfUcxD6tl1yZDARTnVyy3gHERSEmgTiCUz
PbDXVupgfd2sooivg8VzUz5oQXzHq5ZuK14kkKpCeRS0JnP4AbXOzQ2W23cHG7rI
fpdSqm1tur7BgTqw/XiavA/bxPXQrLdEsVqX6KBriRJUxqplrMtk6ighSxdc98gV
rYE75UsWcVxxLT9sG5rYuNch1ciKNiBM62vg6aFpFUgry9qn94/oXSeNqpVXEZSi
lGztYFddfvjFqYOkOuuUqDVpZak1Cvk10XiM6GOrBHJFSKdZJJNccQWf+IUBXDbM
Q+TbWTBP1w3y3iTuBXf1Jlh0vFGPQvjR3CPPD3sKOOQiKaiAtmUO+ajY8Yys6Azt
ZCBWK2JVxYf6IAup9WN5kHzKUDteOD8yB2v2GAAdubMQuzNuxwpLAoGIQUW3OBq7
VFJC+giLkQGB0sgT3kHnm8zix2bmRgrKqC67aPHgfWJJlt3+oxXoTya8TEIaYVgC
zsEGbLnGK53ioaRm3DNraOq1xbZaMdO4SPvfngS2oC5xt+7iH5ypI/mGrn1TdLCd
bvm7w4aWqyYNOoY76VS7LJMmz/fXjd/s5FwmxLaXT2ntRMFhCoDAO4mJbA3tOOnQ
b8OGgOKV83mSlhO1DGeYuP0VplXXCCt21k/WVplqJxeAZ6WhCRg3NE1Ukb3eurPj
Nd+OlophyRJ7qoA+wMXXz1aFveWPQyq08IL6FpLb9eMVMO13T1kdmrtkNX9SxTLv
WBd0PS0bc3dXWRYQIK416CAslNciInb2Z9yAnvxAFsfKnve24i8k57gtMZy+jx+/
nTFFXqmj97/YnVD7++bCYLcB4/kPLypGBC0IN1NDi3OUHUyrAMzyuLUNyuC+yheM
3MttMVdgFNflxs2L3fSXPrPX8cSudTODSfrHRgZjMpRktrvJx1aXWLRBUKH2/R1i
l7+SEM37OiizSOKXCa1EBR51XZizKPBJNbrWDjqW5AuUQPdjuJvlWQYefLoCOpbM
DOUU4bAjA2bm1lEU+5pk4YQPEri7PhIrucoauIH6R5zsupVsoK1m1mA62X1Zix4F
yfBz3P9ubrMElIcxm2DsGaga+1o0DaF8j8ceqJL9LvPYtOsCEdfcxupBrmo8vFe1
QeHrbPmuRz7QWlDdYXP4A32dbvIGpqaUA2sus+09Wzg7zaGzZexmm+YN/7qH2SWz
Md0T2uDJ95ObVkwOQ2UQ1Aw2RxBSCx4Qp6mkiKmCSMuW7O4XT8j0oUG9gKN/ipbk
nGZLiWqj5cF2xiAhKJyNR4/Z59G7Z0Jmo9O1G6CJ9wISfCYivjszDlNAnIYZEqpz
oCj4Oo/eH/2zO9uFmtNJDuKdz2EdxNyq/yk+vU+nj27wY2DqImx2A/IqdKRWdJc0
2Pjt8Py7YJufPlaB/6VKMdNsgpW0YLzAkZrlLQk/Xem4AkeerqaWV0g44Cp+ToWa
fIu7NHk5I2hS1V4LIkgHzys5GVsHHH5q8EEK6XcHe6Q0oie+kr5krfIbQygLSaal
92DIgCCg8i+UyZ6bygr2Lk4mq4nV7RzsdZtnsPBTRxM5JBe5B3SSA9Ikt/0Yg9l3
tN6RU8itwxXL289KO86oMYmOhwwXCTXIbhywBQ0uhC63AoFp9rM8or8JIX3PlZm4
TcRNsB7BQV6CmaxvSLVgyVLNcbUHOH+sYt9wLdFvxcsX4bRm/E6Hz7Cip+43jDPu
UIhlDVo7k8yz2gkxLwcu71dBqNVRXm0UGFv6EyYhlHQSHN+Q79nlnCqNhsgYt7aK
9aq9VDR9dyot6n9x5URvHjAgYXxHNn8PWanV1/nBEhfk7BCILM22nKaaLFbSuTmf
onbAnaia0rMRoq9W7ZiL/iXph3ua0KYiWmwn4E6nsTA+DSHQd8pcPgo7VTHybgB7
2fS6YZ/3NPfdn8G5vx0ftBWv4UGtCb7K54GPtTpRKfjL4nhEbjnYSmJXhYjwjyp3
4bMa7mGrAAZm+FTQM0LZM4jsic7xsIFDbB9Yl8JlJQDzB59a3xdwv+0S46OMvhX8
kskiDMQ70ciBRX+08yMpWPi2eVKlQ/wLi1K6uQ7GhPOTu2RGS+1NCjC0yYJS7PB5
t37MsmGvyhtvMOnCA1lo0neyRQmNFj/I3eGagqpBtpMWjfHxb7x9Jds+McWfcrFu
YMjzpti1Fx22DKXMOaxcTRpAdioCMW0RwgLiJvnME77CPUH0+Kp8K1uGj7/Pu+ZP
nJKPXs9AewZ2xxuTX0Twxh+PHp2SDDazXEOcfbOh9HEKtcvFHo2PN3fe0U4lGhMy
UnpFrnVaUvKLozbW7fz1orYy7x6YIsZyhTL9oKDHUSqQZn7y7gK0RKZP67OLn7nm
QapPXIx6PMMM0XC9JltjnlI5lVR10X8bsJyGGIFrqpl6U17McpIwcMqXInwdXExf
OKk24yvOcQpXt44EgpDIy1E7c4duNDbQbf5swEELqvaw79TBks0iFp0WidKWgDhu
diXRR68PIQ7ivOmMi3gzwRwsOtFJUUUzYMS+bC8cgG8Ybm2otgOZve0LqbHBk6K9
d1QoHAFfAUUsHnA02eCQOB7HV0PAT6H/OMKb4qQSxc2OTw/xKdkP4b/1IJZJwc3c
YIy/hRvwZbbj+MAPtIuiYzFFWhGY/yBVPVuh/Np34nR3ggUADupzYEiJiJGBUnJj
fnw5GiR4dJcFZgayquenBKm7YDbOCxPI9JyRC8s++3RRw1UyDEuwn1iquBrAfpqM
VNsKmRJ+2drJD55o1MRXEDw0oucrsXE20k+0zonvuHrdKjiKHNgFG5at+3mOc7Kk
/4Q3Q3+cFYieSuMvfi5Saa9nbPHVCYJcMRZ7xc0Sug8PjCOeRGaYO7qAUDJ2P/Kh
4tPrUpd6NpnFGeWt+fsVG7+qoLjvAacLbuNeNhll+OWE3HZ7ruxVXdmm10dOVHCv
0xqs3g2RacTepVuBV5nly2mXHEuJl8bYBBrjsexQ8QLMnQ33yBbDur5pkTfw07Gk
mudTnGCufAzrbBMh2e1RCG268893GdKQnM4IVda0EF1v/Wy4oYIMdTwgXWkzNVLH
AQZb0UlGupYquiesdg+Xl5wSclsXTRCbcmodWQ3ASVHZTUxyyWaXkZNiEm+7WzHT
EW5LhuyDaLEaJpVRQkZI5vg4rMDIRgjkL+FST8WoJsxJ0H0OAyxQySsqhQ5TK9Qr
CkYDzT8wHYdcIbvn0G1OKfPicPuDCI96kBXkGurN6nqMbvEvVmKcX15YHEU/n1a9
BuCjOJraeuHi9aZwACfg8RfJs2u31kFn6C87kXfrPREC0f+8/FJF1hxLWunz7LeK
SQuvbVM26KDJgTkW0dmaq48tI2uHsRV5+LtL+aqhTZ4Yoe81cOWWEQLCr+JgPrPL
8oBUVQhq1V3LCdmGy2KLCZPdQLSMnyA5yn0CT0G4HU7SCQC1SBdkfgc5zJihgUAK
Bbo8Hem6hKflqVjz6xYPIbRsRdYqzf8l9sjt6lAN8FXL3Ui90gAYK4YKZm+UqnyX
jV4YiHI206UoocKn8iEcb6M/NMk4fyqleAVwM45Sevqi3aZHikDThGdho0DBgN+6
gGQp07bRHgE5X8P292magFvkTYclJ4cOdRZcPegoSR3mkTf0WV+OmsubEr7CD/5u
ZZmCWICPb8Y67M8vXCb1yfcEIg1EIBAc4DjstycGJD17dtSZwBhiA56tqO5oDqE+
30DBHPgp7eOTnaDDVhNSUuAAacHUcTefG2V9iv9T8oKUbqwigioy6PeIJJNQUfac
AjyGoYbaEN0pgsNVfxY11sMQwme/2kGa2rI/IGKL1jyyKJJZSP7rG4qcM4xX5eV6
aLm19t2rb98IIrheCf5+1W2K4oQPZLVv6/XnVOJuo2knvWAAgzRsbPQg0SZWNWm4
bA7Ak1szNJqkpEwve3kcDeNzycBsnVYrV5lbMbP2DbqFfgKG+Wgaw2NNd7tXIJEC
c4awaj5o3zYkvTgXTUTVCDejbwK+kKsEf7kojB6vjMzJTeISC6XxfcOJP2Sd3jcG
wsecCyt/qDGe28Egzf9qX+fjyG+ipq5rm1vs/2f4/hxrLkBb31/8z7FYK9iyg790
Cq1wYcQluS0eVQQZ3Vk4OgyZJQg+5Xv16e7+hkXorQpmEA/6GDfY4veHH7JBS6CS
4t64bl+G8veiNZj5nIQK22D50/PGpFEgiOjgKu1uOOtDSzzKHK1xQSp16V3TVA2K
vrM09bVY6g8U/A5UbXyD2v3nd036lv332dHS95MyUByMx76Vi02t1JZ/6WoXDBSx
NxWKC24Y4U20Emk+QPWTiAuZS6mH1F2S2AvVz7iULnooDeGZR87hLvZUKzxf1m0+
x3gqvdr1PXmuuOyxDaNpbI2N89ZDncm5+hEaMT3W6kGPGO6QkOLWQRNARDbIWwqY
eF0tquKR7Y6XP6RE3j2LBA/TxDcxvWUyzfOencIPq/W2Dp6HRdpOkMKnUI/UwXo5
Ev6EfSCjwplzbd/QnI/lDbyVNzJM7MCK439wDQqefIv+Kq63/RAwoNENsvrdxNyK
ar4UM2kky5iL/1rBNlI4m+vu3FspSCdMllvQFEr/CyaDjdfISaXt9kAnn/4roWWD
iPkvKxmetH/JheIMviS2Cl3FZAt3DEHRo7HdhiwUw+e4Q+fcWGpbl2C7Q0aUmB6O
UvM3Nu6qOGCet/wWXNyq00LyUsjfNm3LRtQgShV/FVSr61htq2FXjKBMLOQsP5yY
0c1CgK9JOArRK6zGq+VzfEEfyZ1ZYLmDxyV8wjo37UT6HkgheP9xX+st57sHKLRL
hRArqo5ipP2hbJuuO5tAhNfRCxDLcJUezuLPFfQ1GkeOKMd2ul4NdgeyrOGdpKfY
eX4UmV9EWdg59KbT0ZHdx1cAY6CZkdsGk8heG8LixTsyFLTVBC9PBUAhDvCeExRh
SZXCr2n8ovqg5TnaCHuTwsj90lMa+u0DbrirtlzgJEkM44M3OT3kODWXO6b/kOOI
7bgo5nhXDy2DrbLM6/Ke9/jjkn8PpWKglEjvCO6SwNEVrw+2rSs3G1xkP/lzq5ma
VWzbmTirwOOt1tlnYL0fULymM1Ch7+MROzRBhJFUClv6ahdlrovWId3LIFwZZev2
7HSnXPZqovzbQz/O/vShKdNWLo6tfEqKVC0EyNzAsFs6ASy4xCkDD00JLLhjRLCf
CLcqxOnLvxz9EFdL3D5BN2xqyfEQN5GJFCLyZ9e+ss0XJ+o4Nu3LBH9A2tstRBFN
X+tngPqntkET3kP8PdH+F/9dBElg/DS/evkll1PZxmVCLxDQkvnLF+yo6lPZAzbj
HcbDwIwaysy6u7D2XJoUrWhQJBG9rNVG4UTG33ZUefvuMM3Icu57vPGHobqMMtJe
mSaI1zvzWvJwAnyMBnR3SelKHySe+e0+mdIpR1dwVkSD/mbtWMafm1EGxqpIyG9V
PwbBJxlAUohbscsNd18VcAaXGeVOWAAIqHsxSPv1IX4kP06RfoBPX5L7cVGwYgvf
IsJetuZrQY/yraI6jY2oYYX2drUWUffhlFoYv5ITibfxleQYUqLLZdv2xoOHstX/
zfTxSmJec4OUFjTMBnvC86Sxd6o4h9+LXoDH2ZNo2FwPsiTQMyDazmKMNJDBT3Kz
V5lSYICFLNXwgmCQuTIM2yw/xBJT5HQJ53JMhqDpy8X/7rKZc8BSF9QBm6k+IP6H
NOHWo0pMHoUkMylmuat5KO/eyMAwQyKw0OSUuWtjWHSoAioD3QbsYwVJ6XrWSyZ+
z71SpGHJ1rDd5rNSG+dLR5Sjh/jOapCvJ336XbOY4macbe3kH6edcoBZWTwdHU9v
kENUGkrgCIQgdGOFKAp6KP+3vfxtQ41ijC+InPGMeuVkI7W3aaWWxwO+d6uu8qjb
RcGkyWXZYAucygu1q8nzqIGdytFGu4WBdgSXqBuVVZsww7QiXhcuf+T3acNvRgo+
tFSUsmyQT7iB5MW4P+NiLp+ugVqSra0nu7wkFwh9+uH9g0NW2zMJTQ2gaUB3cTTH
huA0gu7hyyZr61AqkFHgnlXqHN56oGLe22b6XseupNNLasPCSjmLCt7HbaD5cCDm
Xo5F1FGWMs++tjRiXLPPRl8MUUqI6LJw2DTBk1K8Z7+Aipi0WvndSpjMs7oATk5s
N9ITd/nPNK0Fix++l/c4z8mj4xdknKBNgov7nOogJ/ys+/1uRUaKFqLAMW6Nwosf
huhfxHh5r/6CmKWN8uq4kf4O25DoSlVj9nL3XDDvuvW/igqYBGb377nBa5vMBBcW
HoSZJJ7EKT5Fnx0H8Y6YZDLSpInqPvMzV9DKOP4oZg06uaVX88NM+MZ74hSJcJon
P/dNH8MVHq+poUDOBk+txSzNZnCelc3RblrvFaL28IIzLFU4ucj/o9a1GryCxeqt
iAw3CbohiDruGJmTi4kZqKXmmy7TmW7C3AuL4tCHULk24IlHlwG9m+6u0y3g7i96
TAI9qLx4T7+niIqaP3xi1uC8zb3E8mtyMvJ3bpzBCbQMZ0o9yfzlbiyeH8dr1ZqR
1a/sA87kD5dTSfHYh9TxkTGcRAs5CUtmPTxKeEvpr8DayRhMcQGYeGMdAAPeDIa5
dz7Cse46U7JjCdsAIn4HX+TU6+a1n25OG2lPJ9x/OZeAqC+uqrs9BB8f/+Mcr5v9
PHYQbPX/xFW51kIC5nmzxQMynD2vwC/a4HQAR258ymsIOIq958Kva8JXUrMujnuz
kG6pbfV0Q/jFS870NLvdJPCMc3jHTJkFsT3/ph9MKCCUl0d3YsMAP8ZHBqX26Rxt
jK4zmI3hz6JiazMnQyAlqsSJNxHGIKN8BmODYSpgbWAfWHINSNri1fDIFrd/TBeS
EVHDfgVUbJLLdu1JAxPzNZEntC68qWxnlKXlWUD7tGYYpOPxz3z/jdAb3+zA9Sm5
5NQyls1U/KW4HUjmKnmnb7+njpZVVLFO+evW+MGcdmE36oaJeSRCDiNG6D84ESH2
RiYX4Q7WQqWRcpVI+mTTh9LfmKYXG/rprCrCQtdhYcLiQMFZW8PEB4p2gv9SaDlX
d/dlcHGd6b0PZA53Z7Klaj2zHt8+NGewHn5u4TFFQy76ZZyC3A6fpL66R5AfGzPn
lUkPRuYkWxnqWv4pVZrZlFoXglhLvQgyzddR9wuAKzIqAr644bGFWRZ6sBjc/h68
L2s6j0Tia3I0lEUQZnrSr9WhNpVV7L1z4qfoy5XnPEJ6E6p0v3fLWFJRp88lAqVi
CDASoKQiL3OV4/HjImaKx1iNqxHYN0J5Ok7s3qzjIXDO/5yG71zAts7HLLouCb9a
kaGU+yQo/wUs2Vj8QsaTkioDnYxbuAONJdvY9hovwQZgJvjnXSJ1u6HH5YHTFASR
8Qp5eb7DCc/YhCeNTpua7zESUdhuYGTNNlvn9+R9VWn9x6o/Nm0z3WJfggxqFwRL
Hr8nA7Y2hpUpLxEjpLC/LApG9bjAFERxFDfNEt9+eL2s3AYTRF/30BB2XXdWArzO
LW/oaCUhERkKcmLQ91z1t+EbXGkjduXfsI1tI8bP6r9jApYobUkJeAu0ZFsia6NE
oYrP+WkiRiEELY9WpigyHjCMhdp7Uy7IGxoGzsJLDyhrfq+ZK7sTnKPRdv8CSDiV
R7uzYMZbgSTWTV8OjwnnF3uOV9Y8G2KvM6mkB8Jq0vPZbOnFcOqnjWQ33nvA8xLt
WKYrgqBL5T00P2b60dfE+48HqSNiNlGR4n19aBhhIWwRs21r/SFuWvVNMpZz6ZR/
Bv+KJ+ktVEfH/+ffPT6AeaWhyAWPEyf4qSXLLs0VusLA0q+GNkQGTiuf+bVwFED2
xueSg1EDSP/k9SX8JHnHqA9gYCfnIxiwlMNsw7AHtIUBKMCLLVlVY+7YC+nrSB1H
jlDN8eCVT3MWvLHRbSaRp4NVswecXxRA2O8+p2F1JZAhrM+8HKriNLmkQB4gYkSI
rMTD43crAmnEGtDOQKZlWL9/7QI3wIYJ7pFo7IgiQCwUEDFl8Kms8wQD7Ljbf+uO
nRJhw2g62UyQsHSKxlIKsMNyV8XsDdXP3rXeSKjrG8nUkKAn2gXj045oFtFeDHl0
bDHZ6v+OaP71bKBIk/stAbAjLqYMVngvBnHzrWvsxHfRwKZ4ptfz9qYR3YUHTdTc
FhWcG+AUTYN3YkKmLXcB6zY1L9wuXu5vlqhNnKCVG6xTeuN45TWNoScf92+o5rOn
e++uXKe9+zp9/Hr2RsfjfB79xMayThgVq75KghTih05Mn5FmZSHBCnjPpRmgKMEP
b9LHcZfzUBxAHU8wimtgb+1lUsbVIl8Oem4cVE8xIgte6TwNLlaG13oVGQ9LldCJ
0EFUVxfS4fKOVXudrFoyiXPr6r7BMSkbFJBwNrGGl8kQ9/E03ocZcW+omBxpnaIk
dOyoXx0odyIYcpWCjGpFXTPsD79MrQGUqVgl9bIR16EYj8oLbpw9/GOfegob4kfR
XDPCHHdV6fCWvXtFI+SXq8/8YQ7l5RSlMCU6zwf+mmCG/Qa7UNYxmqXRlXWKZyHR
ilywexatZMjthz2epEd/AcT4VesBHqVPqk9L4MXo3L8LQ3tbwFgRPSjFnnAjQEQ8
xRSecGEShHfKtbER3kw7eI2Ae7A4DVMtij6MuXeD1JcISnAtt6zltJLezAabf6Jk
tkr53LUSVuIp65V6clOYL06oY8ra2X8dWmuB6Kl8GJ0Mos/32MVankUblMwvDNcc
MwMmy84FNZ+HF6niUpfzJAks4DRXPY0829LViD/Pg0aspZ7EDs1rIUkz1b1uUNB4
7cygOcNEoEArlfyDDy77rpaH+SjtDqA8nOEeIVyaey1ZCE0YfDqmJ1X7GyD0cphn
QVU4w0dmsOxkgyFAf5kfI/O0InBluMRRBeTGmu4RZWO2d3dGY0Il0jt0npUfSPV1
yaDKAoov7QMmDBbCnRtdtDjc926ylUWlpJbYLb15hnXr6/smNkQ7hA2sIJjEwInj
/AMftWBoouReyeak4OUt0OdpdY1nSO+ei/wASFy99RhNH/duplbNOjjr2zoSSi0N
RvHag4DaIxk9tJioNMFDBngojHt/0Qj7Pd8CaJN5lEOz+rlsW478UUJWXtwPJAll
3urGCl/CIwiqHdtkdRsZ0i81crzh4BRHfJAeht9/PWSS7EhlBq+Ho+roADD47k0A
VBaEZDdWbHRjO2ydTWpmXHRCmoc5LDp2oY2JPUQoagB1/GEGV88tcGtQtE359P+Z
exYOBm/b8NQR1ntvSPxZceIWvG0fOEPc/vf5uLozc/XzvT4bwv7+xTHA2JqyaXLP
aOOR/EbhbdFAuIRSPxoRm9HTnloXSIl/LpGtq8quk6hv7P8JGCePcjGsBoNErKvt
J0do+ZVItvd2cCpJQvIorDWF7yu2eR90uyxCSrlwqOKO3i9WdtaqisOu4sp6237k
APfRCTlp5SUpI6LgzZK9Rf8isybTAWzGHCKzj3MBjJ1zT1izhzF43X1SUDVmI7zm
XeXIwiuc5AF+/fGbFyeRWb+sfNTTPYdKYtXT+AoP1UJ2BjrwAxEDp4WIqa4Y1nNo
bqeEQvUImNsqtfBG0B2bvkO7FvspmuNmDYOt8B9apzrC9zD4qm5hzjdU+/041nvg
fhKPgz2JqO2J2YNTKPQ2rjLtrbOw7eRIm9gEiEIloASA4tYJhHo25a4Q83RVz99V
o+QWp0X6A8gKNJR5xSngej7iDgx0bxOo2c5Ql9kf0Nox41ogT61gzObD4v1HI5YI
ddRLfKMt1wFbEXYKUoIV6fFgLATPGAG3tVUBYFMl8dkD/f0V+36YU26WLFsrCaSJ
d8ZITIGTDk2/hz3InnhQo/EmoRSjkNA95MawCpv/JBWTw1cTrU0ScsZy3p7UYFkM
VXJKbh1lQvs0MgsO8zPtGvPSaLcQNak29Tsn8KtwDhRv+zA/29aRbWwggxuwtg2M
VISEzCdWS9P0+knSdKGFTLmt4PY5KYw6yJWiqurz6lpXOa2Y5VQB+aADAhwcvl4j
Qr2i7jWwQtxoE4TlwKzqrfCxcmf7u28voW6AWm/AeDcnyQQnrBndATV9C7WWrM5+
f1okR5Ho+vtX4Mu0Vw0qZGUgkzcMZ4mu5y7D+qzRj0AA3pN4H9TfkLPvhutaWtbc
AJwQvh1nbwfjxYY1GWyxKVDf8YAOqZfxRjk0WzSB2iZqdptBt9yEjGDF19IHImV0
4XKtZjLOct38bDyamZD/sNLlZimuncsP60yItqxbhPZ9axZi0mRw+IR0X5xChYwE
K1COIscDhYxFSS7sFdWdw+K9AcKmK/M/MmKfOTsSAAXdHvAXdHV0Bt9RwIwYozb/
j2XX2h3TLnD35+Vs2+eT81RLXyNPh+nfFiD7MNcjZDIqS5kFmqUhg29MQhZLwdpo
WpbQEId5vPUelQ4t4NdNS82LQ8kG3msao5wujHMJG4czxRfL6vdaWxx6x7W77i6i
H6FwxLX5reor2kZqoe/7/e7Nii3wHBrVuF6lW/YsD+bABwWeC7iCmJrMI+A9hr+g
U0zt+XB/w1n1cE/aW2dMPflS8kpdcxBirse8oDUN+l0Q2OXNQI/diYS89t8cuIl1
zwnpNoM22Py4+yKnEpB/h4b7IP1wTO+4l4rCwBHkPyPTevheIMvrBcx5gGdPFZM1
6ljOlRKOJ2cgeVKK+Ec2urN1W0zx8NIYCOmBOWLPiKR/eFOc4nq4FnyG7AWjr6e8
Qj8gdvhnnqxptsxOsuRO9zk74TiZ0VhlAurGzLcIg72VVEdXgwul6GSfcl84tRJb
ODPQEW2FlxRr9W2OgwMzvxndwkmo2s9YxfIMVvzNW/I+My+TVJsE34mj1K2OEtJJ
Dow6OVfH/9Zp8yC3T4ZCfRzpsnmFZ144YPCeCXxeBEkrB8in3f86r/WhMqjgs8ng
W48Po7Yl7C3tkkhptG8mXnyQi9UPQF+j8OQ8LdtZ/nwrTJmeAoMZRFHOee2viYGS
Wzpx6V74QdqckkCtqDX1FjdsnU1KNJAB4BjW5jnJOahjV8dj32yC/WvEZ2qsQ4t1
sF8ToSA2KjxEVietOHlJj0xb8miWvcLLUl8AL5nHhYTQP6gBglX+EIQbxhC0nl9V
u02qW9M/86/09DJq/cJ8jZMdHyLo7tK/veHSpkK2CzddbzLIbu49/3ekmhJl+umL
gvlWLHFcMZe6lichW4kzdYpVhbtYrYvlDo3qSWr/0rzj6joTXoKbp1vaHvNu1d5P
/0CfDYy4PbARsIYNNneZvvpMJ2jIBOusfi870uACbk6HjNlhGVlVpKNzlZcbOSl9
+kbqXGxQQfp9x4IketiREfmhX1HiKU1IM2MZIc+VE5ph7e6K+Tdm67FIaHb/+z7a
m0RWdyNPS4lWO/nQJw5Ml+GBEO1IZv4R+ij7VhzZ4/alt/GiyZhkQ61q+Dy6fuxd
+keoe5ZaDXW7xDIW7gNRwFJgWsLwSpBIZ0/AKV8Gksucj4l2gBZuMjnyz3j4/PZl
pDANiYTq0ieOmD+LBABruh6y3gfHhtjsMMQS+5yyad/isYqKCorrUk8ATE4nU2zp
ZF93p9eZxEcRSKrl7qCRskEstZfpWGMemDlhEdYFAT77XEROcYrcnYbR/RR0+PrU
53H8nTAMGlcHC/lh6sIeueGxv7OBH7eK8L2+CMSzlO0o4ObUYgEQWDezvJBTiJ16
zeEoLeDtcxSN0UAgY2LocVmdnnpnDlW74GgM6RZRKsPbJ2hb6P/xGRTROsCbvg8a
23Ca7y8MpqhW6Hw+O8wo8ugsSmaViEpdi68xKuMs6R60G9y/xglm56bW04cBWqlp
QDRp+jYLpFSBr6GZe3bDbg5H48BTevRCfk7NNjQyotX7eKAjU5XMGlwesicLm3MK
5N0AqF5GvbMWDMGwwmLaasUJWKunfncF4K4sEHijCqHiSOOyGJQNqcY2tDpabVTH
Ny50nThFE4RDNXY0ajIJN9lsY6LkB4L3GjRHXVI/YdxHIVhPCxG5okL8fevB2ZXV
DtXvf7uPYMNViKnbD3TgTLYvv9Gj05fz8Od75fQ5664V1m/xo3/YMKMKRAzhzpT7
JANdme0dzy8p5B0yEk3oHBbQ0XEqUy2FrxaxKU6mudjnasKCA/k/1rcsmGF+L3Fy
k22LeU1gzNrCt8CJw11wX4rZbh9iH022ubTpSL4LWsJwMrxfwABroyq9uL1fKVw7
RE++aE1looCE8fGo8fanv1kRcKWkF8CDHFqDdNYkkDEWj3vtjLYWaH0/uYgKog8Q
0nMwq0a09AoQL4fqHXpOejG0Hfhys6DRuZ66yAODdO2zrc/AdbzPiOW1wWE3YvIr
y+Nou8ixf2R5D2eyNu3PSnghnHcyIpMzm3EiKBvroSj/IuMNYVgIJqi1af3KvV1J
d12Xe8gBmb8bo4zWTs6xj6nF3TKUBzkbXw5GXCGN85/VWFGmB0nmRCDJvYQMXmV4
wMZxUoASP8foHpL5n+up5AyNZXekKeGZ1V0k0pE+JlmecHqiVwRKrZHIDE6VXpcR
bp7Npqme086U53VXeR2OLt40Jef/OgvHF/4xqiWkyUDQlm5VweRJm5wOSXk+KDln
dOWxPPmyXkAV91nVhG3uc4SpBhs1/+kJoa5gTdOkdrddNonG7INzZWk6RG+julrM
jo86mxYr0jZ6omnJQ8SOGokgTylOqEVWEuicKhKUETxD7wsK81uCMPa1ZLxTSsm/
rrd/6tBnOpTXOIMOMp0BIFYalV7D/5b6ix588Wwk2W1YuHTFIPBfj4AWSt1Qgntt
aa/oq4XxuYlnKc49lQG1vMSByNIdSA1ypJgpL976vKx0wArXmRX2Jn/JMvcLeZwz
4zOtDCg6ygdoT+ZLctrP1HhGBS+Nzt/fk0AXWMk5nVp+GBcRbfZF0yGuy2o6HlP2
pDETq1+5BFdUcfvgLQQaSwGX3ASJ6ypE4U/jReiZ4oQwAd6C7jjsvUfnYHM5MzJs
qMYJz9WAt0IsMG0+FhEqIVF6ofqvtR9qKQz9gQfo3HYpzq5DUzbIryY7KtFCDyzj
psbIohnjmUBADyQiSAp1nfJNkPrZLvI5d0JDVrhiJUvJwNTnOpfwj4EMojyLBIa0
I9AhXSuhhsHpWdI7T4rZNB/HrRq/fyC6s9y9pCzyOi+uYIWfLxE53VdjD25/yD2l
qtW0M/CJDXocF+x+wjKClZJcxRh0aG1FCMob0OaD1MuhsjO3ZS1b3JHNLh1WtJEK
xtKVdFI5I6l9y4j5pIimiKRILZrJKX1Hn15pzF6XbUyuJksgXM/aLuQaSpgN3hn3
FxJwPnGUOXI5UNVRIhl0/68D+v3AY82OkYKY7JAtZOfc0MOEVLeuZfk51KjFLWXi
ORwf9wu49IDefqYuJ2EJnB2Y/ncTBPkBpRKfO2X63lXra0R5rKvav73MZPWv0yEN
QyJ1l0vhCnMxeEBaSIpha2taRKmNAg6T1nG5PB5xtQgF506RI7hW645ApCx8dDTF
r8A5clSgTZsoto4BBqJ/csF0twmYx2uNQKsECj1/7tqcEauW5Yu3gaG2EY3EnK9t
jZGvWw3rC9Th4O5hPBk+qhQltvDQ7DilNTaqU+dAojpl7b2OOif6i5Y0fb2Bqfkr
eZMtzhuLnjcdVTU9yLLVh0iqBQD+AbeAy7vUGx/tP6cfhQCSMkZWjjV1yZzbcBnN
62JOVk3wxnwhxdx9HPf4YtepH+5aKXYDUP/1dAoRExFC6SfAzq9+1ihVsH+HFpjY
CWeT1jlooi9W+cZ6l2vPQ7/xPTMSCIi/5BlfEcVxSrqIICrRa20veAGUaK8fikqF
K/+Vxi325VwlX+keQ74QFhHLF0vqJhj1EBCYLB28BUIbA4DYoy1V8pFJnvBsz3t2
4/L4WxSpGGixIMvBbldQdaLpTcgzW5izU+794j4UihrJ4Dd3qIADsx+cubHvugF9
tl0RQw4M73t5vuok0iRvHgCk6hVfDP20KOlDMh1CtALNkllN5ZPDpqnVvy1HFYIL
C3LyjOiW+UTmQCxm+YPHyPJKTL05Pgh1muYnBLYCxhJIkKXDu6+KOt2znKRgwbb3
kYpATKsf1HG6FZ6FPflnoZBiGbOQz0kf27bVIpzIXOKbGFW2lSbJU3JXdZLbCC1b
Rdt85yPT6e2/BmIpqe/r+/dQo6NQCJyYV3QrGlm7l7v1+g6eBw/Hdyba4azSTQ9m
RoywU0F3Xm3uhdfZWZU837HOQbZYSnLW/Xp1YCmVpPAgqaErFk6aW7i4omLKEHPe
8Qqqsq/AO9QN42IGeCplx+qBesP5IkTfOsQllAMi/W9ujV1qQXHBfvPMWxsW16D8
Gm2Fyz595rtfwSEOgX8JACDxcr+7j+v9o7VlfQN8h322PtrZCx848CZBtCcjron7
looXwTS6luOqyssBPVuf8wUVWeAjAq8Ep5KEvbjIG5qCtutEaGlQo4LWplOyUMOa
hSO7EpGcPE+L+rPyHQrerOFUCfBT5aNctlCSdmOEaBcH5HhqqsF6x9IFxEM5jG9d
I7jziOi5zUyeW0YOCPHHJoV3FJARmG4j2+5T2+xxyZUDlgo9PXjwG3JLAeE2q8fy
QW4pqYEzRoBm0fS5BVfG5RQH4HH/yXdDqDNszYQBMPI0g6Se1OfWyDyq8lKy8xm1
qDqQCyhC/Jex/G0yClvnVpWOFoVkMlCrCAGM5MAXudGHs8ZF/ZQI9SCBd2m2IdUd
3jgNOhPaEVS2lC//M7qjcUXTMGQLmQco3cFfTucB5ykbL/QMCGsbs0+bh9P6CDji
4DDiP56lAXvzoJEB0K3rTFEi1Ccd8J4VRHXj4i9w9ENJkP1F9VhQ7EPqH0PEWyMz
K5kzbd+3HhdH+v0A4UmKZ8I7S2WXSPV9xeRItVwqQWdWorq+4tQf3BHtMfHTx23p
RyJC8OC20Q1gOuVOGB/YpqbhE+IinZXJNOhEn/E3jF9uVP5E4CmvClPTAchZsO4g
Sd6pxoW71DB/ysCAk7/1eiEBLLCzd7Laf2QO25YL1BdF5w+fFolnUwnfYk8AE0hR
0GgV1mEIfhGpf0fszJr5MxE56KMmJNCeo3OPqfxIFy3XK1x6GGJa+VmSDCe55DSX
pB0h/RysJS0qFMdmxVqfN60M0UHu45SvTN+F/TMRizlHPF5AVmmMQ8u+5jgVEZbV
67nU4ipZsdFS2pxuzDrTNjcqgOcb9M428xigu/1vYCcrw0NNAKBqUEtf1IeY1wbc
mVU319rHeINJy9gX+JxSWyehkTp1xp2dKmQcE55bIV2Ye114dMCGXtIdlkIuRN6G
WThy5jBZlu5qsikEX5QDoX9JuSXIOZ9JdY0IOu3fGna0QaNnyraxt/m6pTrhxJzP
r40PM57FrOXduck1gmVHLQ3gs+oYLKwzd/PdOWaoCzrMfVVZFqCZqZcgy2bUmIm5
GzhBHdj/0QZsVYedB7DOP0pjdvvy/hB2c3o1EZHrdZ/EK0HUQwyoukgim31hPwji
O/RPMIXKj8I3nOmAGdUStqIxvobeiPuyO3cmzKYd8nGD3ZQP6uM3ict4PlDRfdi2
Cv0bUxvsV35tDGamz+Vp7Z7FGu8XpTNw1TjZ0NNxRK4punEb82gM7KWeE4HyeQ2y
9sK5iYo5vX7Vo9MDHitkaZdlR6BHmbKhLvFL9kBd+5uWlBB7G3iBriMQxPW8PBRt
zzSC5XAJmvbPzrI0IL8Q8DdxRXJg7qCpZIRg8oLR6A/SeuQI9W7ucEZOhpKzaunb
X0cy9FpdRPrtTz0bqaC18fB2T98wVvIEfcMbwQNUYpKfcDLIHBQzJpEo7GZIyEcu
vi/mUXFeSMzT/WknrCvq7tl0V1JoOwCQ5arTBoOYP1nn8eG7seHJXiKYACj9Ew8X
AinLY87OLRr4z5er6By6wvND50J4KPYvRBP7c1BUn8CEpK/okJbTzRlhvs51GOSQ
eXPlsprhDHvrkTw5pthxhL/4qMn2V3RKRWWOwa75QNzersqIFGM8zTk+R8EUAVIp
F8NZIW1ilhwDpFl7fdsJX0vSedByz8vs2wV5xXoyDZfcNYuXIedj3A8cc9Mbua4+
LgyM6dBSYnFgje/QE/HPlFfy34Cbgu48/ca1LNPzTtp9maw7nY7DaKVHUoKctaEF
ifszmHTnDpsF65EyzmLbVL5ddV/EnWrN/kjKh8obLLA2KNLZQ60S5ll231yGzMQZ
HwfSdJTxz0w7IPLpeHgAFK5KWvXweMxYZmRaIo5OxhT+wZrRGpgGoIfmGw48JkPa
u8XXOdrqXMyX9+tkZTjIeuZvXjaOoBwdnElHLPgW7RgVfXZiX0oA/tHuWIBRqe7C
RvTEhGEDE7U9MISQqgdfP6XWrSas2bKRJtdfhqZcCdRLuY91fuOIS6f7Rdj6zZ+J
t47uA2JvgI0GW5v+TSywjtLD+HALghKydsE9w7R3XNGxC/NCmr8OnW3RxyUFGFZk
kRkqc0GvWJSxS0irlASctOY3uaqgJ4dw+RMJzdGrfhm50ms4UN1mAfq/Bvmu8qOV
mrGeMu2byJBRoO0TKinvtFtHWOTplGXpjP9/G9EcMt4NrwVXtZNMF0TQkSGzcYJv
lZyiRXPZcO094hNN9kV6H/XLVSKb38MWihtjtLPBNgHgha8wI4joC5CGUg9tPgs2
dxZJLe6EoxmzQb+ZSRPBLvyucpfMHflRHSbPIhUrQmDbDE77KOt9oAgP/m8shl8V
KD8sgSosqBD3gPuUY97xd2gN6BKr60kKVQvswA2YlbF4nvfopOAihXXTXy3tUfDG
Rj7h+sCyPWDLfqZF4wJfYTprdvqYVWRR+5YJ47vhaxN8WOUyWNlPEy2oG5842cFZ
MNtGwuSVXx5KaKGKqpWVxiJs0Zws9Uf5PXzQcHwgngm4tCnnsdsVHn+TAuM96YaN
MH612ZyqBlL/Ic4+FvclD2wYg170K0/ILbVlX3+L3D+PsWtZCnDjc/4A/vPMO6y3
6/2mzLraVwlGovhBflc6yWn+/OOIiU8R6Z6mMN0MkuTkJ8itQa7gPXQEkqOPZDdU
vxf99H+bUlIH9ukBwrY4lQ8ck6HTKNoTJWkwc/9zRU6a39ZemiBHSxXfhVWUqAYY
xcC3c19j6tLt53Ab3nG/F7fuT6gYBjLKnjz0G7QD30R4qhzdbJnNA7Q35I3aeCw2
1E9sxfsF2jrLf3SFdTnbqDs4aQE2DWUVTe7i85oUEuQzVBt42E05ihcqIdAWNTvl
xM+q7TLrouAzlJ6tETg3wmFgPVCxKmxymCeZYKqELizGBMBumKENWQgm78kGA7Vn
i+4MNWoxqwkrdXSOFfabJpiYZ1OanGZOEnFDmlknu0oK8MknCe4KvdlMUTMagJLy
vk1sU7oVlEPxctICznwAyO6MN/DMkrnEK1zeLxIVBZeFcJgPl9wMgqN+HlBxIXyw
uciSNa98Hg8hJfuNV2+S9HPPWFsF03JKh2/Ux4zAduSOi8KkRshrR6ecerlSFkYU
VatoHDwDLcpivW1TALEyKaGtez7BMNUdqAjYsHZcVQdNvhpeg3/bvEXoMq590bFk
ZRY3o9dWS266PK5fpo2UCmOLTUv6Rsnjt+5cwCM+8jfeKItKA2UYghj+V/ea+Jff
fS3D2+V3YXcB2BwfebFJG4RR1c2JBbqn6cOUGtbG5qFkq7FhgBDLf+He4ysWs2no
YRwxCuTR147LSPCH+djBu+DAuaMEPOry7q6Fvgum8ZStFexnU2YhCWLFfbOGFYDe
FqhJiS8nm5Cz7QG2tVUNr31ff3/ivKCm0Ir1DPSpZMoE+SnZf4miXNk4/9yDFMtW
DDr6n+bB3uzUOwvyzDBpsDkl0BCdo+8B9xDFWZ9sqO9Rivfz0CAaLf92PvEo+PF6
rMeVTyxSbc6nhRUZcyBVSrSwVl+9xBkSTdDOm9+C9C4iUm5uHD8aO3ucOAO49YMq
9xHjOasecQmNmsLIxIDMWk6IIqdQlbE/9nlSO6rrk/zU3lmPovjW+VevAAKDuayh
QJ7X2Ndz8p3mF8xMJvnQYmeWbmQfAJb3g8/Ca/FyM9x8nveEZPVEikfOKMQxIg/9
oxANf2VzE82Edgm2QkgPr8lX5yE0Q3Yzi5+H2SueaCFLm0ta0WjSbaLi2N2bfL+V
fzrfRoYyHM/tka4HiFGz+k15m+p0JdUKMFM7qS1rWu5J/+3maMTcCMzgzn0cmUhZ
VBKNK9OlByLtM+vq2JgiOCH012cF/YBAPcs4mlLPAeM1H9a2RUvWGUF+oA0lQFGs
6apagq/ahmuq8gsmTmBykGdUzs+QNJI5fyQhFjDjD5eVoVrPiafVzyHMYfIIWSzr
psSSlIRzpyFqj8Vt61DQhBwQRzDyCCL0zKuBa+MvU8FytESUc3AJsISSr+kekhMz
fo5xCa6HtRgQIhl/fZE1c/sdggUGoNrvCxj5iWs2c7RXPXSekTYWJDmbFzanlG8q
WQ0OzsIaZZpD3MdkPngAIwMWPCByK6nB5p8VEQDEzz0OHl6wG7c/gyCswgN9BqnR
0EPof4LnwgoEVrHyglzdlZ7D5WLRv0a45RbMMvy65bkuSEftr1sABnMoKekv/Txd
SS3guyINSylgDe9jqRoUfnWn/CY52lz1hToEbed5+ayVMrc0Kjw1/+51qzsb/VeH
U8bYZJdB32tYkRxXZwQoRkxTTuama7X7iOj38OLmCUdlPws+wvPoizH+iw3bRtZe
RFD+B50HoWbwJ6k+IMDXp8Bk/JVQWFdC2IPnK87V/WGug8cltc7o15bbNwfIoj6/
jWhOeSOP//C6ca1H0Zu18eAuuv9uM3A9hT1hb3OtOIWHs4x3HVMGopC8qWb6W1o4
ywIORaDdfMGCj8HJe4VJamWo24TFdlQGOSoatW3h7gcQQG59ISrwwcnx3f/TfGno
XN/ck1ET/3JWJcXlSyaWis471HwcONpQB13h8v5NiEsA3AKP21pj/pj/nx8WbMiW
LsqVttWqkLd7Bl64DIjos+49En17mT3B+MCu1JOPVV8LR9tHUuVkuo5BsnwXDtyW
fIB5xl2ZjKi9ebAJCSAW7wDFNfUPCyivIT2JduX4bCQAnTCX4+GkCRlFqFPisy6t
DRjrzSNS/FLiHrCtfNHx5aht6AhoQtWTIZdd76WEx8sVJ8FvJGV//J7Oi5DHF67X
YSQj+C9P5z5QgcD50ulspgaN/tpLSBqHzJK0G333P9PuT/k5bYvFbDLHvDwN1j8X
c2dswqbycN8aes4jc30r81DFThhlW1d0zXcewjdM6UvenZgPgZOevue8XQI1IZ1Q
gb3X4LAiVmN0AI7LGyeGchrOk2fxlAwYr2KiWK4NPVveuATamomhEWUfGe7FY8sS
OvljqpQPFYOX4FG+slStEq82HeEpGDUIAC6wRPYcf6ZlyBpMyeo/l7p1X0F/PSSW
bwj7Qz2LwX3SNzp0jzZnl4lpJZOZIXJ5065tObAkXnAFr32rBasQ2wxihn8mmKJC
rtCg1QIXS1v3bieF/d7+2LR6iL6IdQvgA8hMVYOAAeqKaruwxRqHtER4G2qFZ9Vc
WmXiYXBBu1pm9IpXEr7C72plALohn/dV0II8nF7oWDrS2jStovdGpq+4Fw6EWY1i
FsEcmC7vTYSdTj3ZpN8lxODnzg2z84tOvcmlIUCXRQNkMcXsccj5vn+Or3sOxi09
SBuEudnsWTS0y88B4hjjN6avqNWGZ8kY3z4vWxIawcss+BpA2uAjwwUS1w2ofWXv
cIc/v45njBTREccMJeTd2+er/xMaplcHB2jsg/V5RVD1hRLWv+SuW/ONc72kZaE6
F6hVfIusVY32As3FnT5goKD7I7QbNQV4oiQG9gk8k9tNzuENhGoAv85+xuvhHVTh
meRVA04uC053NGcCzNBL4vltnMAaI6ib+c5IsEpkQri40u8EZK0Rf1yyxwbpYQv9
PyDIB60suxFekXVKj722ftk7BJcRD2Qiuac61uxwGo1R3BbHBxET0XdY6BDpezGj
SqBodUGu5vl17EdaMkMI+inPq33k3GFtFgXk7AgDnxPQApDtEYwcifqzgdQT8LQ3
8rDH+DKSmvyoap55YS8s0d13UkyCTOa2WXFSRKAOZzpnZufTVSotKeJ7xGZcfaxG
tfSwtjyv3wGbaKLJxx333JvJjs5J/YtckgJZfM32/YU26lZcFK6H8dpoIDzoelSC
O4bWqB7eruUipw/J317YF7AO7wxsiC69zq3uMfJOq2nEIv6p7svuv28EyqrOh/Yp
iX2QGPLvNdD1y2+WaKrodM27sKgDVRxIRZ1/VKdW/YWLIoNhDaDIheeYADrBiWy0
dxuZ5dktrU0h4KYGFNF7D08JYNrU1opIn7gktjGMvXIZqj9HnWoD/XcaeDB1kN/E
nsO8LMQ7hhfo2A56asmgUOhYWW/HbRMHnK1OwZXr0Qgx8FeFlJ86hc1u1yd7G8V1
ccnc/Epm3SeHGD1Ze347Umt74LwYj2Lj1MKaXmM5t36nbZ7M89UnCiKzA1vn+H5R
OZkFUqp7Hmqw9nvu6FP8AFkLAXxiV+YOfiQGWHD7w5It1HvQO3w+2hCnm6DUvil7
igM7ZPR6d1/Gpzu1EX1S9z2ySwYA8e8661MtvBNna4W1XE9Jh3s39Exu/GGCfPya
e3zqe8D5s6AzsY1VBBC+1IlzUM5PlytjKRpcGOLSxg9LODuNmBXHG/D/Ljn1Apzg
r6a7yV5fY1BUbsfNSqgdDne/RO0JBOl7UTfkwKuSzEB6pMdH8uAe2c/P9a6kkbp6
27HP9N4yHTISBEogz0pdpXdPtH/nHNkNuURgwNA9SJFJiRxCdNMIMGLJ+gqhdOup
N5o8dXMWxaYaQzWYOP1RPEozM5zI6V6eutObjIBubzfvwx1M0xBKe8UDAIE74k5u
hS73fRqOV42TnejFH7aIfA0zFJM4s9dCDdVmlAN0+HPlH1RFp36DxGz8WlTPNXz7
1M5Obso6BXCRLXRIDlXzuLYrf1uvzz+d4TsLifwNL5t3lwG/U88kXPQ4KGsVjCDO
ZSX9s5U+5O/bEjEkyIqkVxDCr9CILYr2T+qu1pl4LpGciVl8ZtfbCuNrTZEU83gV
xIe2m/xHHpujvTWeRxjcTkH1DhcvszJ1dEIecR/ZTHdVvGGJBmbOos0qChYXd5Iz
PO8rOLlcfw1k2KecO4AinrbolLIQP9gmDdH24OTVWAoaGP7AUn/IUZC5w4RbefyY
NIwydCwmUJK3S1SnHHVo/Ty67qwsrXrqzQ2cs3FKhTeWRvqDX8wq/xSXHjwl8Ztr
PZBZ/5rWi4c2uUx0Uz6nKpdwyGHQL85GAjdCoFJXGoXvUd3aq+mpRD4F94kWScp3
iuU6k7c0NjJHitO9Nf2ziTK+LHCEj4UKN6ZIDyuiB29vb3Mde6uDcJZp/UDeCTk7
4St7AIqCdYsa6w8yqHGZ79Pa70QV522OIvd8fnWAJuEwI13v7mX//+wAT9Ht1+HG
1w31tg/Ij8ux55arUoXMBeEuFQpuQXfgcgiIYgqHHLH35gCAb6wbx8gcGt8Kpnwg
wChnolr/DQkygbsYQeG41NiQ7Dq1p7LGgG9ZwHsPojLNMAZtBF2dIptEr6F0mQZV
LrWGVWm0QNwYcXRcSleKnv7GU/i4q8lQFGxeYR4nYU94vZXo4u65LYoXmxVAABhz
0h4Vio0Q6xVX0Ma815p55oNqbyZsGH3xrUAQhzAIJn0RJ3mGkIO/CCOQBICwPkxm
/UFQuWqqu96e0Xg0V+Bbwblutr2i2wBxWXJto5Vko4XiWiiOY38z1jmvSg1r5k8W
Xsint554QzrefFUpBf1npqIydieF5on3XkGvX7/4tpaECxNbhGjWocuiy55gLsts
wL62MpGR+lnHao9DajnQXcg8dxdG44YiCnlDP4gWd3TXBcsq+t9GRGAcC6vaL/qR
wEfDeJ+rzzHwoC72+/efQ9vcIblZSH52fIQIK9dm1oS0fdIhxJuCiPf0QDsGNCNj
953WMkelttNnbEFOzoZKY+rSLoJJsgcVGJljyuE9ciCQY5e7kaNIvcJpSy/VjgLa
OimNZVySXnDIIJVQiZ9mO/pkOFINXx9R4ggz/FTqrLzXGabs6x+/0NknP5No5ZQ/
VExOuxy2F8qt66g14Nxn3juDvTroAj0l8liw7tdqAtNqdHc+Djr+9GWcshFBXVFj
OhadR0g5TLuMVaReiCF2jv3jShY2ZXvU/F/i4/Lo3sWH919qjLzzgmJxaBd8OTeK
8/Y9CWUMdqcMbcEZ4zYAnWqjyE7EhJ4db4ClXEApoagTmQ8Nj7utxf+MLDoSfiQd
WLWlMXkaherPVI+GCL+ABDAY1hr2BEA3KuhEwADPrHz5yrTRqLakX2Yoo0BbaX6s
jMmJ/wZ0T5BsiEdOnRnlQsW8N+irXnmIV5fNKgID2QpPUETwsZW/NRWylflTAQMg
BorvptYGMBXBaEePkgSulc9ogLqy5JYH5mLQ/HOKmOKOAlicdGg91gUQe3CpU4r8
F3zwcIcXB/Jd22JBTRyVBylMjbUK6t2grlespevIG9yVyg2X8sS/oTSm6cxLX1Ma
kA1AF8iX2EhGDiNBlh4TxstznUVXmk+jKbxsIvn44bR8KTOaK3JOLnvicMvqmY0c
p7RFAdSMuncoivL0kkQZiDJoHefFO1owYWvfkYZO4EW5QjXDGZr/KmwAxESHlGt8
x0Nv7avSIrPUWJBgV79MRLTqgmDz0jzqKC8giXyBUxMoQSU01i+uYK1Xnf7aMLSl
KSktpEdBx7Yr9r0DDDUYLwygOWXa0sDZFyyYElxm/NfYfWEhHobpLde1w6uer+aL
C2GWFgxv10xwPCe+Zrpv+fk2s/uE5rlObbOj8PF0vkinz+GvAM2U51s7UgfcPBlM
v/mY5hS7Oo+CA85t1byQR98FvH2B/dQsF4seF28l1bmNbmsseWBx7AxdVCpyBt/k
/nBXHwEZuDJs+uIOcDncqevEk6xDCU3ykveLR+Vw2z0TEt8j+x0UsOsIau8wkXKW
tDsZ1tgLlKMGuyL1AgsH1T38NgG8gkAFN8MXo3eCS2m+gkYXDsm8EDBpZnIfo3i9
RkqtF6ooIL1R+S9LoXI+l+phZYtlSri7Ya6xB3SBON9gZq09OSDFnMWr47Aim28C
bJOM7Gx2Lqed18tVEDSdvuE/KlWRK9MHP2ZJ5yYZ0QVR6tMjIBk0liShv+O4eTN5
DvNqaFuXJBp7IaivaLg0nZ40SVCgQQL87eu+u4lTIpDlRJHVpZCld6npUWKerzG1
mRIKro/MOFvwHVY2isRg4M2nggyNxcfCs+Yt61Y5qfngm0VypMDMl7TpHKzWeuQh
RoqQBd4ZqxyTjr3cCD/VDE44franGxomak4VkuOKD+/rTLnhOz+Is0IQo8XLpACa
aFAWdZ9q/95jwc3uNwtoC8RhCyxn4Fv4dhYU7K31+TzgVMaKav0/+t2/clcSW1Xr
OQDIvOsACvUYHA7mUHskYrCnwDsxxX/eD8cOMponBrFBa3p8wflLRbrco/EOUfTI
peqJp1A0DqnCxY0frdGa5fUehgWCD9rPP9DJwwDfD2n5UuyChWFgifqTAdttGKOs
R88BEpxnh/ah6LXb8deCOSBOQQoPDdTNtvSdLctz0LtWo2AYJCMzZFMVpaoi7bJV
TvKiuzrhjVYZcylJ0h1y6VLnU6KGpJkBLw6lNk+YOF9pHdsbZeMt49UeyZg9iAJd
2juwPb8Kb1Cbu1Nc6GwrzIb3wr9cxFL6iHEuhakNFvHbdvKE68ULURmcYY1Cl+wE
EvJi/hQr43dLmwPlQYEMamUa+q4/gjTyBdD6h1GWJkXqwjcHq6IM3vrw11bFPzl+
9Gtz+tS0/4OVLETiB05nIo61z8WP2usxgkw8+ymVa/YclA4Rv2xtX7ga7vSIODJu
dw1E9ADe3+k+RuqUTe27p4qYfrlAa+2vhvHeJ/sPf13e9xJr/dbAiRPqB30WBAjD
cw0l7Jde/nm33jjyzzTIrccNgDv20cyE8IG3Ces8WvTOJp7VrQ5QgHQBLDYDFwP4
m6yoOy6TQ51UHh3xMNLBhHePD8vsTaGHzZDAXBqN6lMemF2QYiMvyPJiRyLR8TXc
utVoM5wT0wY44oUMSv/6px6iqXy38em2oBomzsHiiiH6wT9jrnMrGG79sdrGt17N
3MeOxKsXH3PT4bfZkamUM0iXjz0o4hf9jak02sI0FYB7cRK8ZEKK0/21twINDYW1
EDIZJxTubv9liwvFGfa5X8WpAuKy7V2yuOW+JNSiO3M4dCqj3huL+x4ji0EpBpOp
QHpt0NPisZhx9DfhmCdmaFwgmgdRPhVXOD/UqnTk5ued3JSvhZh++EkUtsLDfMYM
MRE2yY+/cB7FT33u/RLBji/JV2Y7cUxqpeGjIcu7wcQ3zcqRgZHZfwqYofnVC2RY
AZIBPhjc5JS1pKoqAzdyuKeIxonJUZVlxPj3SfqhDIZM0+MosCS7JgygVtpSCJTX
0pGGilujBsNajScOWzVyUVAU/kdSc+0HJ//2TRHxK9hLpImwCSS0nGvJPs82BD06
lk+XoW55kSHok6n6j+DSsri8pHzLrmcupHnmtqjmyHxpHoMV2QJF07MgoZMRFqVD
TrYmuuuWizgdlNoH7oGNo1+tV9U8QxmCYpfp1LVVrD5S/k0pkU8OBAdbR7CTxb4X
PzTzuJe0UB07RppI/WunSU6wTHWRs+9nUDCx3doBlzfM0WTIXaVGR9xq1gJIt1OR
4KS+mOo7CcGU0ElJAKDQ5ljDiQlE8pFEswebNoCFrKmYzFTJyP3B8H3Ob9LLa+ls
P1Kz1bMZOW6urCTUInel+k87EZO4lpnW4gXcn8CoyfBBl7bL5twRehZsZgMmLYCZ
jkiNmnVGPY+Cyp+pqyD2z5KoBWtiFkiKLmXA9bhyGGypTNKJrHrzlyIxy9y7Gc5L
8iUr1gJtBQq6Xqo84bdT0fxK6mfbcwgRmZ4heGhy5qfiWSY2yMtrFhmG3sMbRj4+
g3acwOepQ+s6ub2HnkDdfPJhmztSaHPE3Oc6ZCJM3i2/va8tvvfdEzEBTdWFhs7G
rFTcCFrj2UjeTCdsMmXDDTbgGIzH1v7tbZerjOwLdmKBsAiZTXhSX2uhbTlteMOe
4pQZr5kYPMNmMrUVhOdPAuFFYg7yNgxGHjWgIH+jIhfTyk5PQkXvZOTWK67IScix
jVKJONTpkOE35p99FDkYpvmqZwg0KLHTMZ+nruuU4gl0BVtCCaGLdmdFXZDQrKdo
KqbWxOtgBKTbU0IOpAHnyIN3G6d/QsfXsstnWbT+oxegcWNgz+uETmksblB2JnyH
eNKr1R4ltFnHQ9hxudH/J1EbIuFIS81QupA30gXMNZ1Yh8BfvOK86WhMpu0fdw1a
GDM3xHqQCaxZXfC3ByUzOoCMHInA792gzfwKTJqDLn+AT9ducFYFAZQigFmZYEk2
jQvtzWbY7DqcXYTX4J2W/xIhqa8fPq52UU3Ol3QKUSB65OjeR639WovSOXUCx08P
h7nslGe9yXIhpr54qTx4O4UllxoN8WokSaELDvWFwzKm+mp37t9n6eDYsvDKeAbS
UceXe5QO1Qar4cAHxV8EtDsoJ4Oh3B2yhIx6PjwebRnnskNf79OX4aR07q/3a/8G
RCI2WFiyL3iKT8QMXzLRDiyPyCYOM2tZ267pP1Monsx6FcnpU2LvlvhNb81khuK5
TWwf/d3yZo7F9o3UJX2Wx+szm2b8iO4c2w3j1Z5vTdxuCfDDo2Gdg5DvS0PGWgUQ
hbNzkxDXFgAoQFSs7BQyS1eCGx7xvgDtoF3vtBtByL172p+BLxgtIQCbykQp8rPm
6Q3Z3c3TaQzWTrX6Rz62DojA+Zc7cgM1kN+iNzSF956F4y/cGL5qzT5D0ZZB7Xag
eiyu/0HJXmzoUtxyarwPqU+RiX3cFGCoW1EvrkiTBHdoWmP1BudOIsJ04Qu3ug6C
/NJuImBZqlU7peNHPUAyVCHAhXbq2ydMeOwsTV6MOFJb1599dJUVkLl75Hned18a
sIXBnb3EDsXfr1P1Q+7MQ8LyjFWtrm4OZNO8YuZma22OyT8s1lEnII0hAVRz1E7N
SadurGvk7dN+qFeGO96JtwkWleMQooCO/BVEGbadGM+c0tcgf6I0YZLTwXTxwQLT
IJXmJaiZeQpF4K+pNXYNNR8AJVLZ+o3OUw1IfVv8hth7WZ/8btCfpu8wpXHqM/S+
Y+b4d0LswpDisD7v+8FmqXtAHa907xi3dHp3iyGwJ0tNLMx+0FHh5D1pO9Kw1y75
ngM+6AhDrquSFyU0MwdhyqW5fm5p0uxaV+Q93robKXCfXv1NWNNZQ+2Yfz/T1DJa
LZ7X1rd11FgcRs3MFRAU2p4f5Aw8XuGhOTRdG1xZZ0XjRL78FlwQSTU85jNMvYOn
zsLB+itzxRLuz+IwXUPPB8PAHmsaWmqxVY+mJ1rh5i0QVfcrnXSO+RK5T64W7udI
Q3F08IMKxp07yw2bXdVUuq4yPFowS0Whmka8vPnuYbKOUXb7kB29yDDG+1TpAwg5
+TMiK9PkzJldVmovntRtdkiXAUcmysauOSctnBzBYhmwM82MByGtYTC1oJtMQrZf
teGBzoPchZnyHuKJEZ2Ca2v/hQ7QtiNlviENCmPiEyUGZIiezk7ya7/Th1H7uvIB
gXM/w1HDLj5TU3zv9QXquTOaFQ0y5n1e7eA9hIL2Z1160yPRaeR+YDm09DqAp3O5
E0cJIclEEFDVd25tfm2YV3k2nhXUW/F6BxqfVWX54HMVdPDryqzaMBa9fSg+btXq
fm800R8SHHPWrG5Ldoi5sk7tMTR7QeCxhLnvQ4/6UwWq4ZvdgiznkUr6ZCPzRSCY
ygCY0u/oU8U5RvXaT1i2UIHLtgG3k+PIZ7wL9Oizkaw2TLucxVtHnbfTWk6HlFWS
DZH2mr2iCMNwg2bkiegGtlSTTW/FGx3XUZrv9isB2gsvCxYZk01xzkvbQ69EQ9jn
O95kQzz1pS/mvGjkgngLJNbArnFLVyQqG6yCOPR2dI/2K7DHyBMTXgCCPn8Ivu4N
8w4zhRCmp5CeRBHN6lZZAUs+TQa9k0Wrq72a8RslHL+5dKaXZYWs8tEvQDkzAi0H
kxjqGzFnjPss8BdDO2TrLkUXM9VL8uUK/OL9OEYeXAyzxlBFTqHajaPKAVGxBkLM
LbTiNZtN/1hOQqltg9Sg+YevTm6JjQwOVFCo4Vwr58uLw6kvSsQfSdXb6zsJTXtg
802GK9bAA7VFatnsIhG17xAZ1nacnxp5/ufzA4EE1U/pKk8p7tjjZMln3sx5NTsz
c6xm+o2r/GH03JBl3VU72LlX6dSbVvmGf1dQ/R4oNBYgRXMZLdYt5CZXR2RPKh+O
Pw3bcUqdfYEAMnEpbBTBBBXwdxekJrumMSCxan1ul+ufUIR6F9vEnTlmE7660gY+
M2hXgeEf8iA2MjHv1unnmu12XiBu/q2pmjnPURqGoZR4OGeVfw8EiUhdnnXnz+nf
w2XsKP6Ou1NH8BpX4sN88AXAgW9fQeNoeHKQN6W7hWC85UuJ6SXwugKF8TlEYhhg
RHihK3QU43W23IC0PxGzlFM2PZHF3ihWG19Mal9TSimmpi11VagG29w/PQDdWUgc
oXffnJVI21RSCL8Qvzpd+JyYKLuxZ//g4vXS6J84fRVCjOnY2OL/kidkERwaKIoe
f5c6Gw75nGNoK0U9jx/+6kbuXOeFeISzLUJkgj+pPaI7Hy0Jtvwti0D5uGULJ/Zm
crO/vnuWhWbL9aQatfJYGgrvMGDaV6XgkIZ4/DqfDt1Zjjq+HIY5Gf6uj0tQ8++j
DWfwXdhbgx5w99DhMEnMxWgrTk0I4S5qwpo/QaByRsNSclJVBfP2QbS4hObTL4l3
Wm3KWjXtcmMyRaZMoUh1U3DCP7D+iqs6f+e138l0CISY0r8S6nv38dozuzEejlIJ
bnH0g0DonG7dINk108nuXHsSVm+Iye95DHtZt1EyePstGiQFen9C1JSR8KarcQej
V2l5xuBEfkci991xJgfvuqgsgeA1tCWXBAC6XX1wWLwhbjSweqz2t1TW85Kraa3a
vdJ/0BbckqROK/ADfP1ZCRe75+MPniZX/G4uKmTVWDICQ3neByqTdTth8OlA9c49
uEOufl8vQMc6hqmjdpOgWjVyu0BlxO7DtKk9HGkFUy/ZMiaLvoFKFcA4I4uTbRco
2I2X7ngD8L6mg8ehmlb1txFr7/aud+wQVxDo224NK5ifYC09jLz07Cx4n1IHzg9G
r5Vqmub0XoE7BaTJAiUbWHmgpdyn2y3/xcP0FU8jBAtdDflgZW3bPJ0NdPGTeq8Z
YsYgnzPzZztQsyq5WJ1e2gNt+MzdSURlMGZViDp1h38MhvUyQME39TR82A0J8HrS
63ssbpEOCe7a+TqDPbHJUvHHUjCdwgoeooO/W/73RiZvyuvkcj8YeVC+RxaXIVsW
B/2QbjW5W3z2pEJnGQUQIeeqWy6Pe+iWFkQVvvmeRZrpI2HNvT0tDafWvTD0Du3Z
dcA6IyetKdZIWIYbIyC7SVX9Ot4LDgbTifmGTeOOBbECYAsYG8UT8zrx2ofGucu6
UO3llnV4/5qRl1m+ZBSXHTvawViwmJj9nqaF27tTJLR8kPk6cXi7yvU64HjSEFgS
xC0DHw2+5Da2PWpwh/gjaYFHD+0mQCb2plmemaTa2tlERrQ+mUPbHE+Z9eHaHm/Z
ntkfnmcCS+oObkziqervi4WsmPDmfS5V2Oa7VzQX8MqBDZ3Y45ht0tDA3cm+J8oq
LCtsFHLJyYNF1/VxhXknNmvAg54y5VKFnrRmvfvFzFHM1u/fbPp36FY1qOpkbg1P
0L6DWRcWij2917b2YahI9ENjK6F1LvNuQ/QpnPuDN16f9/Y37RyxaN6LYSwtmzxy
feVyHCGp6eYBi01N3/iGxaj0egwKeh2q7sw+3WjjlwypleYjGjQv+KpSONv93cJR
3bhCQ477IWb0SlJHLkbLQ2pQL23an7Rloam6BcurIuEWD2L+Z+TJry67tO46JtY1
2rC3MH2y5n5pDAjAeE6WXwArfYn9CTOSuFtLPXu4+B0vU+KM00TQbK8Q8UHti0nE
jmOzBJN5HFFepE8ZJVSIxuo3NUa0NZE8sUEnTwGpr+VqZyTF4b1vD6WYTywwMJ1R
i/s1A35zZZA6GUdsuewwKCVhzfXHEWv+H9bvnXQsu2cV2XjfRUMNE8oht6QLPpYQ
yQd6Hjxj9YnkXAOScZErHIw10KnOUunyWvNE6QlhEvS87X87mm6ubY0YeHW13y/k
cZor5vj/tSXRsk+6zL/hcxMAF9Mjcx5/kUzuDM9OyagAQ2q99jG0WAemmAMwDLsw
JuKQvvdYXlg31m9EqEzFDl8Za4lFTYZ6g5+EapjsS5uutI6xUXxF4uw6QaoOme7p
bXxs+8s9GgjGEVX5hy9+S/wC48WxwDUYOd1TutVdbU+5ySS+YFh64jpkHn2ldt5a
20en/HShWulbLF8QtaJjXwvTZGbAbisa3Vd0FnaROneQJ4g+8NdlFlQQLtRS/p+n
nev9j3YzIif7k8a5J3brX+R4joz1CdYYZe6/HiMcH43ytCmJk4DBSXc66p2itzf7
gmPj/TU4pkSOe5XSvgYgHhkQqWKnE6+QrbePLGiBnwcSU7JgQWvOCTbOyGdP4J1d
tLq8QbyO0KAZ0d9Egqcj/SKcipFsIUXoy43T6S/SycORhmiC1r4D7QVkA5G1Itzr
IMiWSG0g/l8f5XRS2pEfyzu3Vnu6NHIVipoyQHyyyiEt08XqqTxYQ1c3JbvO3RVt
Bee+mr6Hr49HgrYkq/Jrqn/UuBx1lhotMFNvbGcndBJNjvrbVlI8tpDGyeC2Qp2P
Cq3VktaV6c516lL3edCmdKnDlZOFrXXKcDHNeBCRrI36qOdjdLy+Dv9epy19exRR
MD4NVHoWHGbpiTn+zDamvqzIYKl/m/rM6yz8EE3nqmy5sAUR1sZIE9sf5/up7gJl
+axOS56fpkzPucKxtfm0FOUJRZlw5lr04MMgqB+/YV25iK0eBhVehpd9cr8ccZ7B
Bi/C62AutnP9TAPxjiglXyO+AfRMuY9skcMR0Xdz3HJAh1YIFq6X7LfXxPr+AOWW
kLQgQYT8Yz+wBM/wCO+qyMtJrpi88hn5CbfSeLz3IAReAmTY966JJFuE5fXHZ2XL
f3EuvDzPcSzBi8khdG6zlEPQOp1NR5M6A/ubtt71alQ6gWlPzEHevUXZXZYfiBDO
aTF/UuW7PL/TbWysPRvzI0L6O31Y5erhUtpJbj1oHPR46MKskqb3uiuit6O0tlh7
604JiyX2H5XsWugy52XSMDAe7xdse52vTilgPHG2cUp9hoqL2KK+dpfPTFIprkZO
dIl4XNOq5Kdhw4ZR094bmHbr9qI5ygqmJ/xIOrOV1cL4URyXtFCZWmnFWmPLVYYN
l1JFDQTVhNXCNgR6/PYiQFICziCU6ocIGkNoqdzwAK1rRrzo12sn0uyVL5iCWTb5
sPyq3Jpm2bxCsn9/r/AU+Tp0HWRSO3paNcd+KA3OcI/hmuPWpDSJxku59BjRO6Y+
1eCKF3VDOBewfMJZXuPw1xm0HUXk76KIApew1L9f431CiGqvMHWCtof1kRKiSBlm
jEgitgBugp8Lk8YobpqqUD3q0HMMC7nydQdgoU6fUZSBcPmGHXn6KkmLrhoRghN0
O8tTyIJ5asflpr0XalyC3LbCqaUot8tXQzCoFvXTJ4zQPA1FNq0JDQ+i/FpSQZ6F
7lxSGY+ADnBlfn8k0tNB9NRcplsIcaQfji4y+zdCuY/Bi4j6qxG0PmW7Z9fp76mF
sgzlYeTPlSFaY9pX5G7GXICrCQ/zHXL3g4sJVH1V0/aX7PeQNxDTEUQKdL9Qped2
MFziT8eiQb4V3wWt3vGElrP8ogAJvG777PGRrUQh5FwGx6PGSxCMzztt4XsIJuMc
shwrtlInqVzTGI1rtVpWIw78zzqrgF2rrCGdJUP+nRSkRnQCqsBMI2mq5kwX6s6c
KHmPnwmcpDbcnvOD/yinxv4/ad7FlRQUyCwApBRpHuueHtCH1irtP0EV8gmjsS5h
+55wR3dVarXtWfUxxMHuu9X6Skh5m4Cecz6nU8JCAQWv1mnniYwS96ux76jGjHKZ
vBfb4xWxenGYw3evfDzn+Gw9b6/UG6rOWDbfV7MUAnHEjIDQvs4NV6oC17Xrm0Vp
q+UFZF7LSkN1t5DzDN3+uRE1u/6codSOSXq0hWB/C4wJBfUvRf/LW3D0ln3Q3ecW
I/M5KEeQuslT3kj0Hj/I83w+FxpfKgJhyN+zV1XcL3QiOQV2EH5yg+uF3e4zsz3y
kMhgylp5Xapx9NwY8c/KMK1gBeqB14PDt+4tcSeqmD53VQxVzdeEesOMn7MoHH8Q
97KBSFIaC4777RTnjobIT4TFDCTIzYN8Z4keVl4xyjYATgHHTKgyMl34rD7dTCYV
sgaZtqn5AXqVZZeEgq1cb7dQh/RlQXC1YY1sVpCSUcTL4c3OvsNjOMw2v2CO/BBn
hUfs3/vqNoL9O5YH31HOkSnXS9qMGLk5CRVKZ5y3IQZyhH/l+XklfYur1oXKSPm/
4PzlCpd2KlHd7zQWuevKiRzLRUpBeb1VOJH7v1v3YkZVMElL6AmnxHitulv0qtK1
/jfUrxM1NnlMhKiMfIcXmPAtX43OiNuEvzfxk8XUjFAxvprNRjCvkXN0Y5xkQazV
LmkXPDvfRGzlucdOq0ns04pZT/esno0bFaMzOpzRZ6eZDBS+JA+PWx7/RrvN3QYk
N4SlhxkR8M+o5RMf1/CIjDMLmdFaDWjfT/q2xj5jc/j2EarWjLW4XdOZdu1jMmJs
Lr/nMBF5aNvf2NVL32WE3XSlmGVV63mW+4DYO5JAFf+Tg2NiFdKoZqtmMqVNBzOy
dkUDnDt3xVKtQxyWihAR3DqxYtmyhttMFLnsud8xVTo9fOe5PgNqdQVlliV8XCJN
gompxk6WD5EN0W962O25qdmTqTGaYcbAu2fMcHb+N8rShx0NRuP4Sv3Jo4jyxIkq
x3MUnipWiFSV5NGux4bu0mLT/KIOnpol29Z2Z6Ra0/68iA548rowaRZ7BI+VCZOo
ebXFYXnbHrjpbL1LMgmVOKSZVDu14FWffcpH5KIY72eRn8sF5fC9YzKM0F8b/3F8
hkQpSz9ok6zzGaNYvH+9BNBgmtjV2gSkfIOdRTpL+iu4bqGdzbVgd6SmOFukFi6K
w99ffRyycMDziIhcLhAspRDjwjK6guKWHstlbvw2HuHQB6e0CBLBm66ZdMsQ+UV+
pr8TLU74lnDFNPFN1axfeSTri82+/1/Mp74LF7uy5pFV2jl+0MVnWczDzCrw+jIL
6JMhIFWnWWRjjF8PVtGL4Qjz9rMGgxSquuoM7chjraQwTB0uMcys2AfAg8ocr+0i
ENz9JGwZodRSfSkQiSDxiSwaUY0y1uBIObg3E9rBy+OsNe+W94gLtT+zQPVibi+A
0GKcUO/njWIQun1xDdQDcgm0VYX6m3MT7jFeAqC4w+W5wiXwANrgsllOAFLpeYzI
LBWQDVTrzFMVDgi1gIZWF3Rxe5uZtZ+E/xnQGFqqhhg6nrPVbBzBsRq4lA1onkxx
YiAwfdztPk8q9Vm9SPeJacdu/KM0MRC7z4Xi5aj8G0nCskxhW11gAnW/jibV9JBj
FF6oBEvINnAka+rRnpYcjbLT457zivbK1Jae8z2BCobcWoL7LH4WoqGBTr0MQJ9V
HulJVOXYqe+TRnoZ3YFqt2WiPxaRix3tt7WueSlhmwsiVrpnOjSvEuew1oxHoKo2
DweUNLhdl2sVVvIi2/98iX0Cfq+ZQkhzMFiPUIZKpJ46rDx76VjU1DhlTkKEjmeC
XqzoU8hCTp2+f5GE4PpLqJYjN5HAbpT6QR+8rIBUTt5G/W/8MFPf63h9OrAi3m8P
vRfbGBSFl4nX5q1xlSQ4nTrUQwqcs7PtxreFVLuYxAts1ijU7sSPhHJJ2bZZINZi
4GMcRt8eIMeYPQPk7TPJRfrURmA+VAz5zanqDuRur7kxKqhhAsBi69WXz0tzIm27
9tXLlW3R4tK36rPGFh0Ka3XT6cmxHSXy2ajMDPtEv0PCw8c3iJeUm3EtHg6gze1H
ZrsUke3yRCTbBNdYYAaeWBli9MwIg72HMJggqRzbvNPACzeyB91PLmgR3qOhNjQ1
SCHOoBxGgFJyV7hGbti/6RNnkrJ/s5MmF/aMRCCtxmLA2PkztRxPFPS5YjjAso+v
0Hjm2rlVhQ5P+/4rX6O5RHJZEFHqtyJmlJmcgObnc1Qg/C+gRwolvReelrYygrpr
zjcXrUDKdGUD5Gc0U5r1jBcU6ucnWVFK8+3qX7DwavtugS0QwPXadNlKw211ZvJ6
yeeSt05+jNEsrk7KyZaES0uRMgiNFPRNjQgNzQiQjqECmH/wdeBymSgS6qo2R6uK
Q76N4Gov0i7slzaDpWrsiDYjkVxepXBSU1YdZOa4PUNgPuKp2tkjVvkHn4ZJHtS0
+mbFA6NTK93F+dXqTRWEvorobLVYdO+IH6VRa5tQx+PoCTCV2P5VgBHW/PICLDm0
qcIqaUxKGqxBKDz51v9Y6Hi8X8ibMH65ASfafiYjvrWgZ5fmaJQPoG5BCE5zDvpd
BsduvPbFIjsMGHstYdK7ezST1VzBsuSW2A9sqOrSL0rFVCJTYNZC3ggd4hE7gwoG
VF9O30Ofq72TP93VGxff/piv8t/WkP/yXDE/SUgHyG6b39cL/DZyRKiCiAFSzzx9
70/W8e67lvvEoZQKbvHA/8VtvBvJSJeCjunvWq7Br0fRWUIu3w+mBBYy6KNHZDXN
QlwTFwHH1D/RKNgWw9ouRrj7yfYMsytIXIt6csgmhJesh2D9l3hYqeAqaXkcqfUT
gEuMOSK4DrxYrsPlqnK2mGVMsLUWBuaQvsZcxEyzna9O2RNWGW4F3QSRgTPmyPOG
dKCKWOxeaWFwGQdU1IQBXP2xCYHyvuR7Ej5+idxzK1SIIc2QGhqUdLnq8TfAlkke
LGkVnazc4YTT4R1Zv07XDpif6F7OsN0h6ZRYWB4QbYe2y0DObWoyT2FXjfg+N4HM
tGF1SWcKEgucLqLGtAcomF1A7YJp2UU4IcdTNcVlrCn6pjDsuKo2qKMO+ry5qaa6
HILdsnEidx40OTAcpwAJyWEbtfWjmao9lZKIp1UygcrofHgUEynXLKGYMV1IO2ND
ruSx2yBTLxOlaa8uhpsOTEXGf9JC1Pqtz+U17ADAT23GGH/K0n13ZrkUdgs6lRc0
yY3RrmAB9EHwnD3XXv/lvUTd5KCRsBMqr7L7K2lpUhUbqm8A6DGrhovSamvhA8lo
5W8ukzbBR+Df4mLGGeYWd8o7/P0QeB919Ma/c63gwt1u/8ORrUKFPYIrzygVo6gC
78XJ1wnuS5JPXYlWJM9mD3sdiuiCOUskcTMFryxpbEKw1TcvdJ1fHbAaD/byKgvS
PMxFuemrULd26RQSLiDFfSfQTo/D/7VFdqX0x/m4xo7DO4MHiGG+luuGmqUW3OBo
WZQuJ1sLuliFpJioDlHNDpcdZA3pnnTAWB6W9K8t6glDnJzE+RtBfJLaNgjUSmmG
FBUNMVJAX69xTC2QBoGOVS2Arzz4n3cyBf2Bgtrs3YDWJxeapWaC/gZ6tbqpp9pF
4Zh3Pib9B6PjNHZ9+4znLKjamamn7zuZWnIH7wo/gxBuI4QYy1B5xATZ+1kGxF5l
BtKWdDPpdxV/Ns4bVhf14VcigVnLSRUiPPnG3XRk+VTMVVLzb2Iu57CpKjdanB6z
WRETs5egVD1J5VTaLA1h2bmvbDM9Pa8AXCFpXF8pqOVET+NCjA516UHi+9qoRxcp
pADvcnU0d2iV8f1i6wC2vWKBFJTY9UC3b15PNrHsMrddF5+uLamPQtR4B42yc1tX
qH0U+C9a800r3Xr4xdVMXD4GR4Bxc6rKwOoAByJDwCB4KghZXteaVLL3tssQ3Cat
5LWWCZiUZblj+F9ohgMeZysC0zueVhtuojFC8nYrvDJWhbg2XOaH1E9Ndi0G5m5j
i4WGQLzUC2nPJFQGvYZomvXXhN+JpSLKaWm8Lpwfgo73SQeApiNXigaZxkeMEhuD
xLky0Mggs1V/CN2J0z/TmNvFZ0KCVFafETqqpOAmv2KPrzfqhvfeGkDE7+gwO/Mz
8iCcNRVm2U1UsO9jX5szba5c8AlMMSt4RXBX9sEnTvhu4cBTaKoA5XQLu76EkqZ7
wEjP1e6UJ8keYMDBSQ6jSJ0U8uf6t6JS81l2Yr/g0H7iFty/20D0l13QY+/YDKXA
KVgetYqEtv/lJwFYCG6jgu2gQEcIGhb3YxcWWCAtdyWvXE7AL2dTiJv5UV+/3SFq
WJloF3gBFKUDSvrGmwjtO2UZX+KtYVM57cNoK0BUyHZ0KMMR/rz9H5UHEhsaYW2E
wrD+MlMCdFvX2+dGyTzsAii/FPrLfXdxSEgxQCTQ7r/GUFmhq1JpXcPVmGzX6Lvo
QFvApjMsWa8OeGvB7KGuFqSDeT1G2w+MP4LWm8DzTZ+sOxzMvkB0hyMY2PeDjt7r
qDwVvR9IRz0dQW3BFy2kkfbJz3CHLncKfzyA24df+DyRUNAA7pvEu4V5SYk/vnOL
jNKWiQoUAERGwLFNffH0fvQ/Kwivo7NC/gMbk0HCVF1dTxw7n05rQ0eTu/o4SXPL
/V88ZzdmOWmlUVvIrNZHQ/sY2C1PJMwbozuE86o64FSogqIWEQCKQSMzykMRqkKG
DDLR9FGzsNpPYX9x+O+VFSaTMefwzBBI9xajx766zXH1pLmNMOluKB9+t9b+ICJO
ExmTACo8VsgbvmwDin6GK0zzf6Gpbj53/+q1JRz4Ce+aNuExCbi5Mmq1RaYp8/oE
2BGpUugWDUa3U4pbfpDTurts2fy0G8CD41plVf5CWuQlTfnd0d1OEUpf8pTUPWMy
DeXhNkbp8PL/9B+gWrYnSzfccq8Adh17EsxPU7Iew+9U7Q8B5w+taeqRvwcDT52g
ZAOv214pfqef21kFrPtuZf+wv5u8ZZVYOnxgkcDaqHiqz4Qef2ZkDs+LbTlxFBf6
OM9fJPhs+UUZO8ZHHol0kKyoLlrAsAiv3uX/o5AGC/KmkRS1Hghn0qPnom3VfhEC
I1OycWFpXLqhTF1W39z3qTIC4QQ6dHThhtgFH+G46JvcUWlx0fwFSEtXJ3HR2Gq6
R/MFVqqhjmZpLwMXjkJ7i0BOP+tSeb7CPZvSYX1Cimic6+Nn0Pk0rSrVBVUklDf2
INHC1ijlkNOAlNPTjN8sMAf4TKVELdYK5iX12jV0KHWJlfFxvmW5YlPUJp7dbrGM
bPAUoLK5o3+ZAwOvqgkyErSuvUtRjrqQF+zv9g6NO1UFmT+aMwrHMA3/LGLhdqgy
2pq0IV7U7a9tfVcoKxwahpNF3V0qfnaig/EeQJrlYlKDnWIzH4+RunKZf8jBzW0v
AlKtT3TG9u1EG8P37vkMX2nbVyrMap+aK2+QMvD1PQJ4wRnr+eTS3aP+rI1K2rN9
j7ROcjJyoS8VxvZEO3KZibG1WPbYftJC0AE5zD4+hjBOWzJ28G9pe0HLIlR4wthW
CwtL0feKfyjIDKOWPZLwxtUsMlyVUiay/038ywOOtnbvSILIhncLq0U4gTCh3T14
ErWhMJhrcbYUtsKEyeWwVywVMLcxWyqhWEv+mB2dOLuNSUZhWyTcYPgdDos85poM
VKD91DIoNcVcpIl5kTzms3EwCakv1kl8gF1pcjrPTaCZdRZfSyS3XgvEOCPiQCjE
HxBMjj/tFp7JlRJD12b6FutXyBZcxjCvC5QznUawxpRTOKpO6CfsPxnztNPycJi/
Zfxb0fMhRJ7MzPaZn2PwAPRPwXgpzFcn/DTh0lhAdSmjj/Vn/9NJaz7O38zQM2/d
7FaoJ0qqyeEK+cSgyNMKL5RZud4YyVRnT18PdjERc+RIaEg51z5A01e3gwR6krKb
LID9OONSdpl7KVMKpFxyexbYsxeJSGd/6YgE2QPoCCXGeZPY/qMRa+WKz+A6BQz6
6WBwv5cbUUCPWn7tIacDUwtHVk7gvzkdbx1YCLflyZ9StyoxsWm0qrWUhYDC6oQp
hdE4HSM2baz+KLnDdhENjz9KzuX5RdkFZOnrmp7ve2nMkMhcdRjR+54rYeXGrPeZ
AMQbHA0qsaskAqJiM0Aqsb0R8b868lKLF7uoKi80ACS+VvCmjPS6BWLDP0YVCjBu
NCB3RAX+bHTJN45ZrVEkMG9xfRJWrzW/FabokJut2PU//+yjpCKiSf+e+rjC/5LP
2OvDKKVqTemlCNwPUN8ErUYCidHwYgeXVkoST45pTHYmUhsHepXl8z2YG8eUDLIn
+lg8yPJkqeXt+uKHC6SLLuTQGMu5CrbN+ueicFTVaADkujQkqlljH6WEIMohSHCn
xrEk8ixnsqUQ7fp3MIvcM8Qe9FLluwcJ66F0RStIRo/qUqD35TqDeg7b0JqFDza/
KLnQxLP0Gx3ZI/rZpKVBCeyGPVwPszewTL6Njw/4J0bsUcgcWZrWVznRCCmfdLbd
eYOuw/h2oZulGHTPMG/7uwfYvBHABG1mDunTFE4w75mW9cgH1lFqAqa4jD75GwYx
t0DiOY5OL8ym/ofyZgX6G33wgq2H56/6FpHu1yT02Snm8/Myjm6WAYpCsmKbPeT5
ibB/rFc4fI7AZJEfUyAE5QeKQzb6tjbUA2SEGpVjj2mxmcJgbXuWnGLhYuEDXLr+
/RIfwo1QUDoa5aPmC1MUJi5/9GTt9I6UdC5q5QeOH0mYCZVGDlE+NTBNezIMT+m5
HzEApawH83Era4AUn+mMS5Us0bRCwD9OepJRhESmSWS9Uc2xg0LXOgz00dtV80i6
9SSpavHhy5Q63UOubPPtvhohovA/70zocYRLA/ouBMNpt8FTs7nwpIDW3UGWt8/5
ZV4+eoFuupwxQcqY5VVmPrqD5N8OKoZ5uZCw703UJSolDVHMwOz+BNpYhV9lNYlX
BT+gkn/V2TiY1C6KFbZhKobFnNMchZ9KWhieuzIJNEkjrKBkQHENZT2ZQOMKr+4h
YMLyPmtxSyK/nAMKmvcz78/QufaktIVBYPSKjGL0ayUP2WgGh4OSJK41RUjRwQwF
hprvmGYjAFqrO1USWWfjeewO0mVGxyl5pNQWKJOqslORDQ84kh3bDAW8NmTAJ9Fb
IWFgLp5c7Y1Pf2eo16l3/xnlVgDxlJ/rl1rkeBU/3S2xJnMZeRlgDx9d9gGnrrNU
oqGxjJ04nUJyBkERoqB3ANrnHg/t00IvcUZy/pm+z4Jd6cMhvv5iHaOwqUI0uf8a
1Kip77JQucUAen4RTtLjb/xYhgzhOSQ4sLkcPh/HZVrCExEekuKHlia31b5sEDvc
0vzSSP95ZfkJy//FYemP6m31foL1IVNgkcR/yq0DVVo1bpD+MPk9ihQtNn05bshc
/k5FvBgaXB+CtHBP7g6YlZ5BMY0TXIXguSCUk3YmsCS0R4DSOJW4cX1BPD8uxHPe
Vt7hSXhpvjwRSfDF4AmRNMKRKJQpch7KGDyKEJyRbI+pVT7g23jzaxbjcvGrrYr1
TCFy6sXzKQ0uOGnCw9gIRb9444GLF9AHKHX7v5vlCsmtAcHqQ6pHhTAQHLdBnViQ
Y+5lzdEWny7CeFCw6OEAA/VTRABf2N+OfZUT7sa1/tSVYs5ai2CkLaLKAA+izLA2
ajv9emAdKbnbCyB4XwswF3wcfjScNuw2bWJLpI2HqnJ6h5i/ElQ+C2Ewf4zsoopa
QEETctetDUdqGOh+aap6xPEdA4gWSImxpC89zpAe+v1Yz0iXwOwz4i9OTTithNP5
BvNLhFQVWUakH4xigBacohHISj6GTVL4QmzpDCHgni/4oQYHkRDw+fKp88FTJgzz
XosTK+eA8tk7eDb8/uQ7jQFSakbZp4t5ndGwu0tbzgtG2Se9PE8WEGhQYSKwmulf
Kjm+DPMjoCcEiorITCquvzQlAWSd4xnAek72AzgSvBOAJhvb4oTuvCRjRi5DErkr
hmPAvjwF4Ee0bCIvE+aJ4z7RkK6fHAlLd3av3x1Rbx6/QY/pIobaRWf1JOKacVng
8qRJ2ri12o/1DrZVBW+SJeRS6q2aIb/ZRPyqps7TazbgRRMzauCTUYSyeous47kQ
FAlJZFN7W/42Z9GiRZmPwnkCjvPqTorcSVGbI5wOW3gJUfoD8fk6YrVReF2N1DxB
9LAqwcb1zspEl6k9JxVO0XIPlfR+wePOeTeiR0ErulTrjB2wWeo1pNakdv9IXfHf
6wVuA22neYI2d64YxNWa/rtcKCTXfp5NnOK4pw9GeKJa1x2wU3agBy7yZKugmnfU
JB003cu4c5L67y7X7NiBAsqK/BmC2FgIEs21IfNNqrQk5UgSgPoMz8smCK8K5Qwr
W+IoP4ilW95dXplpNDZTABmWHh0iIItfu9/PluXUAf2dfKai6kxVKWgthJwvHn6J
`protect END_PROTECTED
