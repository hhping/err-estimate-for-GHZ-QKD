`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ja6riBLy77Q1Gb2duQoas/isfAHNKz6/hV/Tsc/s2m/1Ak95J1dOK55UP/txCiTo
tJO6wasiU4VlPpvfJ5c+AumMKzflk1BGz9UBrDta1KL/jUE6mxxErza7Ks8X2/8z
Rv3BRWgmFTGxawrylbkq1vHAEt8BMUVbG4VDTFsKZyoI7oU5ObXa6Q7DBXmyfDfY
xz9NIjgdlB27mKGX9CQg1OSbm5LtUZkrRyAod3KfIt2EHIBkIVQ3/grjFJD5cidt
R2qOKkPTy4lXEzrbAyzmamMSX6bexWIIDIQ3+UavLVi+qfUjOXKrv6z3zAOkhE4z
xWkJaKuX8Ol12uDHSIdmsdEy1lYX0sKoV8EZmalVUmxe26PVv30J/6u6r2DdNJsE
3KJOzvdHzloI3Eu6pKBHxmggnHwBrvTMwMztFo7rpAjTfNvVf6TpfkDTXcOIOqln
vbkus5m8Az2NKxP0g75K04MWfxTNkKubLWL851eyoCQQbS9dz0ZlzX1mRQz1F+xE
ng8UqrieywOSlqHbjUva3NvhziDiNpRQuj6nSn9+bxY+0iLU6tobAb4pnn73AF7d
5JyIsp0LzEU6a7H/nRkI1R4+VdFtB6KEL06HZm4C4x7E82GJGs0KKzOEn1Xu29aT
NreQJd22/J0y41YV1S1LaJWqJgZlVHpJt4aWbs56UdAdtRM9indH8q4gtEYbza3K
UUunXF+gx0DdPNzG1H2kBOUXJ5PsrcCUDu9g1D5it4OA+hh3l7+SLLOKI0qm62S7
ogSlAtULqZ82EX9Z0p608H4+dLtCWjRROywiVLA2Z17kDFGUqQvYvfHVm0e1nEr2
yZs9VS8WaOOZNk4OXNrLC9ozl8NUce8XMBu3GZyGzIaYQltC8IaHKmRwsjHJl1xg
A00cuU1OqBMsXPUL2ehUEOQ9ZNr7N9MkLX6xJ3efA7zGmrV4wr6i5Wb30jP2pC6n
np5tq3q4no+47LSgZeMd8zIWWe+kHPodHn35ax2qfaeJ4TyvgRguQ184SaE7f0Iy
M1SNh7tTUBTH5+IdLAivbSieicLvCGRHySBMrUXzS863waT87c2y4XjkxtENxOJ7
bxV6XkNciw5sASZ0VE/DK+8P8l+8AAga8v/QeURCn+cBFXXCzDFmzpQ9soM+C7Ix
QmzPEE9pHMKFka7QyXGEPAqkrxJABHHaKeSgRTLo65Yd2odM3ZnO6ap3W90TUaeD
DzA3zHNo3xQkvYxybkNgHCnLAR95xusy7nzjJHQgCvc7ZclVdxJv0QfXWCaEHRpU
lsc2wDvGZfxTjeT+FaeREgYcvlgTPS2OfKowrmnPrIvXKWYXgxA8HPnjT21Qrh2G
BpSeuvCVxDPhwftfeDxqHuE4K24zKwec/1zWbTwrc0XCEhYX/ED1b8jJmUKnLute
FElMr9dtcLZtLSw713c9+Q==
`protect END_PROTECTED
