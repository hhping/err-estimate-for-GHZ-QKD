`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8DQ/YpthHHpCz8Su+wpWf9vE0XtjnHW0WcBFRl6qp9UkAmgQmAfy/BmZO0IA2tO
wt0/zz73rzfp39Ww3xC9DKqgAgYz1dRiT/q2VEuIQrlqH+FqEDnohYC4MiQXXeX8
KoiF/fQL1lNiM8uyEXTK4dPDuG3miCezrHbPxjY9o+ZJTxzPPLkWCVkiWnvreJmW
I5QyjVJr/BQ5ccGaXczbbFsxRaw4xHb2rFfgqPdP6ufMkNiI0Yc+KsAzF3cmsAOk
VEghDQY9OVFx5TKmXrP4X+JsSIiMgJHbIkT2Fr69JA/7qI7idsX+/Wx2tZUhXzlB
m8VoUqeoEt+gNVnyp7x7RkAbSAcbWkVtPEft4UAlSGjYJPK176vM1xcBYbBwog2T
XbQpF0CgApyNcMDL9a+ml8J/GsTco61QeaF2PP75zbtBvb53PTE2j+nSPZRLTqV+
GjDBaFj4XsQtBDVXV3ZrsXLVoiX2WJjC2ln+0EnAn6c91P0IZpN2o2K7L3rj22dm
ODcnjY0RSKge/SjSzouRNFxZ0lsbndiBkHkOZ+h68xBG7ed/+bSqWewXoOvj+3sR
Eq/Hw3DOIlJFq9i/P8lceuWSVfPGGq31elkm+CfAknzuOamIJQ8ftrrmg6I75eQN
xXZtDtck8mXAj7PruRNHyleSQeqdndvPxUqZuMbKwlPwabrk0wXX11ROVyrqUlUX
+BtUoYgjjxvcmaQQnSq1a0kqjlRDWGZDTvFf/4p8b+AiP8MexX5/hUfHBVT29Wbw
5u42udstZjs97XDMIeeUUpIx9C+bXTp4+5dOPm7y8LXym5mlugFoDtqAyrFebIbc
jNxjmJ1r1cLBGtqUWaiCA9QWEgBFD78y+Sk5fEZy/fm8+dB8R2JJpAuR4USdhOEi
F/5IYvpKFe6j4HoXD/FbL8QqsCg/9YCwLBXmhJgmF2EzRPH0I4TsSJPpQpZA1u6U
MpRQVibsjMxQ6HZGd6irh9eMzWVvXMgHWV66JYtDdiGa/H++1qN4LRY54jSZ1kNP
GNir7+YcsqF9c2u2xkc6r6TPnQV1x1UZTYiBUj2zCrr5SDNDjxs0z7/tbxt7Vfd1
7tn3zJyxq0Yw2/8nLz8/YsMjKVsmcNFDFZHu5AkkiiYp0IHsTFQpUmQk10WeOYnB
rk0rjYtWhuYdnBhGXaPAvG6juVKaMI9ur0qniJM7mK/B250ZpSnTmy/uAdyKQDS4
9+ZfTSG8PliNRH2lfjxe+dDay6rznzrjWvyVXm4b5jP+TnpwftCy9y0ygWKuwutu
`protect END_PROTECTED
