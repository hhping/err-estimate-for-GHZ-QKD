`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6Q1vW3WeoesweUYWVAOi6ukxoOc/p83TawXP6umejBu/ZqFIIHOWHyXXMbfeyFU
oPb0JkVd42mr7S48d6h9q4VAPIXoyUBRsGKJCr0IT3TpU3OvSJp/uLD9Z4/9uqV4
Xp60Ng35Zaojpjao5cOR597R8b1zF69m1WHGhO7+/kWJq5KwKc0rSOQ9TBfywJ38
iKW+6xw1GdaRT8jaO47Mh25RpwXL/T8YxqUoBmA8zKrhhNbHshRCTPQEjJIP55YR
AUOfPZFeRMXOaHz+p8ZGbEltRjdLdU/bb6aWStO6dMF0Z2YP/2wIoDWnc/3+Ru6L
JU74qZzMyCi8jjkhWHf1eG1o/SVrk1FITZzah9YFkFBz6CApxUD2prQalX48LWe0
Den5RxfH661sqNUSmcHtaQ==
`protect END_PROTECTED
