`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RB5FuB4R3otgFi6RV4WiaawvtYJ+IQYM9pECE9hDdyOMMg5RdSvY8F+Y2Vh7pCs4
gSBWZmWyI+Mbcd7y+R6aJH5Ir4LC4AcdB7xGvqc3tVJAqhjr53k+HbReHelBSGci
5gP4yHdJq9OJLLGXdXop+cUfTeC2ypkcj0JgF0aTM86qnuY6XcvI6H+pyPuqGz9d
HWF4mnlwbSGF2IwO7kbPz6RxgrEZea0r8wjEYuGaFivFs2N2SmSEo8s36sH8xKEq
cuDC6uAAp7ZMYX8VZ2hkcizPSJzNzLLBLYSJKbzD6lDQG1Nl+rgRr/DjgJBsF660
Isy+WlOmsc1lQINJilFNJtUZIqXCIihV8HnyNYTHzAtlFsDxbghL+yWbuT8Lx/56
BDopNF/xe1qkXHGz5gfDCNrks+P6MixDzLsrMqbod5wli+k5z1skvfwaqlkS/TLI
ew1hYSbLrPKLcemorkZf0u9pZtVzmrv4sVRp5Gi3JzBQuorD7PMXMXq59t98FiVS
s9ytizCmZAp0Y4eTU/g7VK/MGhQaCjp9R9KsVJ5CfBd8OZeUVly19FldVh9/74Sz
mljoVFRbO7u9dt+1FRTw1U+SdhBvRURh0rL11gL0KDdrvh93DsTKb2EDi70tw5f5
EIvI2ewl93v46/1EyqzEOj+ppVLFPAR1l8+aGOFoQxA27Q73dX6vQzNvwLXAaxVT
08N4lLSNEG6RLfGj1a9OYgtIjDqxyx04zWdg5VqCPst/3fX3A5jHHy0SdB7VGTrS
CrJcCuJvDAenIv1l4dYGm9+w/AHwTOkYllivJDsmL/ZkR6XcQHyMqy20JJyF0zIX
N7AK+yQ7I47YVIoEfvB3gwdRzy+IdZPmdO5hmuec2O5SJ2fBKhOiJeDF4gYOdjnc
6L6DC3P8DmcfbcwEOvIZC6+7YMgffEZpCm82o1JFQcHEdWSJUOnz2JmVtF0YDSKE
2qjQfzj+N8eVDElU6r/t3XeWqNGqmgbDz9BJQrMdogc5SkCZTC50vNDA5anwSU7s
SRzeOVUY71KYbRrZgAk2KgekOJ9pk7Vl1++s1e9MpI1FlggsVBjfrx+vFoA+PPvk
vfDvu6A7iAyPclCbAINRaSfmx3XcYgxLuFjy0qwX7r3zz1CANv8UXwYCrWpPFR/D
g/Wdcl7EXUa9mnS6pzuPLBfJtZ302TcvH7W6oGpzelizDEbpTL6t0Fsc+1jl45VL
`protect END_PROTECTED
