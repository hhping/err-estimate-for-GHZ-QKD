`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kf7ztXOdtjoSQtxvDaDRBu0BWTjVmXImKfxZbejX376MjdOYRvw+0zrvO2O5P3Z
S1Dt0h8Bj7rmlCVNtTVnpz3XlsgEWMg7F9tyx8MEfue8bfzGZmAIAihjcQFE2LxI
XTzKq9mhXjyOy2HBaiMg8RNqwoSlzypjuVK81c2BvrBLVzD57N444I//Juq7AhsW
LgLfCtLb/wir9YKgefv/oiBiuYDjr8rpDJgGgwxtyuFdsfgn/mvnTaXrSlS1w88R
BkFt7dmPPaZMx0KIFS/HvCXu6MIpTnr7n7P8+bTk5XtgPS1J+e9Nv9PZj488+Y06
aY0lKxD/UBGv1NljDirl9+wEgImjC+zz625DVeo73M9qScC7fajS+vZNjHTKUnE7
L55YfqY9G2zemJCNDx0ZCVZKWzLBCB8CHqcm5BN7ObJyNux5ZyDpwVgOwnIFcMW9
TsL5BeQ0h1vops21GWWgNKO0+zyKHALs8N0J+zkhmJ80p5hIea+3fUSvh+PhSoMV
Onodp4sz/9xdfga7gXXiHaxReugFDK6a4QRU6ldioiq3vE/xPrrc6ta92+hWFQ19
jDPFVHpZhlbFz5EB/0/EqXYpOVzLJELYZWI9E7jDnvtXEZYRa+2f6lQO7EUEkkBi
XpCUUWaAQpDNHr1NcySVTJkipkJIii3TU42SWyqDNHNNG7PVhZRZ66s/o76WR7b+
busyuDlkHQullax6DweZ6FbLUnj/pjLIbc6zyMiyCgZxgpqhkgnVN1rDhAHV196W
qhiksg7QzjJzuRMFCksTTrLcXdefo6P+rCGvG9S8CYaQyZRDSjJLTVZSlubginZd
Yigx2iX0UibvJ7RivBFgV5zMocmmZpVYlDBvOSGR1FbsO8L3JtKsk3HTJAWNN2UL
R2H5g1kVH1mO5DUysCaOZx4+mvWr/IE6k9hA95aiKtVAEsl/SSOLFunDUNfDigCn
tLWav84CBP+of4MobSFPJtEh098It0MhLdfCVreJHj3eW4JdsYWbPQf5elAWPtjs
7bJsjt9cHN5nQRQFbFs7F7yO0gGY8gFsF8VEnnbND98MEu7NN80NEALjnmMojxsR
EAcLlRtGe5BAcmy+LL4gt/ieWVBeEKu019WuPmL8tyx1dqVmtgQDuHPwc+zXHUeu
8X8NeYXSfJ2SwL8UWY69CDMVenE7/LofIJW2as+5ISq2fIbfZyZx+f3pEp2zeEzF
mlwJ2UIpMNuKGc0QxeI+6O9wPxpyYpxSzWG49UeuCkLmWmRNahl2VBSU6zTCcSIc
M4adANt6xw4aNdXEB1U4wK+GEPZ9qVmXbAe9jLFCEflSSh10gwKW5C6QbxYQTOf5
a16mu0hIfGK4fKBFTyNx5qkN7BUIYtpWgirdO0EoimbNMe14XuMT/BTRgso14VPL
MAuqz6cvxOHBM1oUs9ciWo1g0NwDp0zk5s3eVWWAGEwF9ap46i0ISR85XHNrRw9D
yWUaG5H4NH62voA7i5GHBhmEH8AGDEPhJHulRp9sTeafYmqZbAPM6WhElPZmoajf
SK5T+dMG0simYy+BpCGU5eDK0IlSr4Gsw2r2IpoF2YHggLxiy13ibWkiTUtfFHVw
o7VGx5bO17/cmiZZ9jxmDKj82n0bOrqYu7OYioKSkd1PIM0eKPPeewkK6n87Hcvn
rCWrbXD99UF7JPIy3ra6Lr9jy86cmvbAlWX5Wc/+tNfCtyfn48clnNvbO+sTsLmT
PWRJ0YX6lR2Jd48vv9z0GPqzimDRPc0uZcNNF8RvCeS516QcJC5fFcsedY1IZ0XQ
DN47tXp8+YImDnEYIol4/V2t6eqWXskvnxzF2uU8QB8LJ0HsKBwv+V3LT3uUjlLk
dQwSB+XQWxQju9w6xqiqQ3vIyVTuDSzkUoN8p2ugNhsU/hKOlj3esdDSZs0FiKRL
0kL/tdewZBLZal3MWRHM2h2rWjWa5dzB+qVhCPCGKiWplzACuThOLT8jIzFno+Am
OlGVpT/4oAQeuwSI89XVTpx8BhreL2ln58cl0iYdnyhcrrFaYUAbZ7xc8XE6YW9j
FRvRP77ofFpsk8h7/UgGVWxneWO13X4nPkcAmTaWca90v/A2pIvEWaat4V86izdg
qX/2HUR5I96QLwj0vCl5RrF2NDj6aS7aFR8eYR+50aLOtsdxk15mBhxGIObD8WC4
WKK+D0B4N7/Uwrp+yv8aGl7rwN/9fzUD25cJPxMkN7ucDuXWIdJIv8PO8lu0gADd
Qvorrh3qazTmg146xxZzXwNrldwxeaGWd6AeObDDBsrr06mq/zWDkSMuKTIOCFKs
7WBknu34yjxhks8WsDoFEdxyU3+ginEAi16bjU07ICQtAUtVeSGnj6XRdwT0eJJ5
BMpvsprs/U3ltGYCo3mDgFCKisf+QNiyrcXSuxvJgSeUyy2gM3aHCNzkeBUlxAlP
nseaOqyp8UELEFMIHmzi29VgEA98qT6Quxv8j896DKt7Gg+OraaMcKNOQ8JJg0ps
diTOgWyZh5Vn/Utq1/JcAA9rgrBv8NS9+6ReGWm7SXnmaCC1H5ZhbUNqccRunk2u
DmBO/I+FmGPSDac5HdYFvmVVuNOcsAAnjUzsp6k+SuH4N8tidMJ16W+q0RDwbKL8
p9yOSnaRSui+EOde5GnwGMrzwGuxT6W4DlZtjL9PZO5sdPGdxoKRdDgVMo5I9sM4
bdOTNzM0CIVPpqspVVD9qTu9I8HjhFPXz9fl79GCI08FKpOY+n+RJHnqn0U429VC
N+cKUCU0Tbe3xNL79IoQBWQzgfeA1dLY28HYdE/CeVMdTRZYrcTdoMQzv2c5MtVG
A8h6aNxYc7ZPk0ukwIOpQSQMH/QXI4tLa4mpOLv+1rrlMz7/n11g1J05BizvTE5R
BweW15TXjwh4JVdyaYjkTH0cXAw44Ofk3nT2yXuOGpT0RtcD0o+PUDABzSvCG09Y
hOrOZGagMBxpuVx3EM6pNUPq7nhL0zzwKmI7BCAI+vPCE8qXoOqlT81AyqcvGj6Y
lFvefhUpBByWN1E4R9zEbSh176GuMYNJ7sC8/mtgNQhsiljLSrD88uH8ZIVQ30mV
dxo7FIkbesGCQS/aNxB9eC62bRdJXX7yDDMDWyBOt5poom0HT6cUQj2KE+eYn/o5
Uf5brQOXm9oTHvIU1D3scFYdkmXW9VWU9CzLco8d07dvTmCy8JaEtqwVhdKCqHmq
oezI8ry4xEiGtTye1CYjXRG4eWPctO2HK1bw+g5HBb3jyoadlEeLaungjHWQjZZ5
N6IzFdAXiJcJ5WuNBHvr/5ig52brvBJo57rDJfRslAecmSTDCdFozWUFHxCb6yzp
w/dZY0K1edm0Xv/W30aZzcu9/4+KpFHYBw0hFbSWAuStk9bEmmPqU+4GgTZWLGLF
RJ/sR/rqGuES7wgA6K4t2kAx97iZqrgoFz2wkMZR1VoK4X8w2n9hgCZgNtZmMxXR
h76HF2rvbAjwD91TDUvuZy3IXYNne5x+2NRX2tBYW0Gmh1chiJkDAoG4+N934Qqe
MiDH2BaFalT4RJ3cB7gICiAJlFGjztAkp4l0k0GeX4hRefKMfu5QfZKATRteZRiO
G+W2rqQNJVV9sKaxoMPU1I16YSLQ4mnvbHbgpnJoFuRGdwLysanOK9tMokfBhoby
2ObrRqwqTYahFPQ4EVbwOTTZLA+cpGV7FjxXOU4J/Ksq3ofBXkjeXosTg9Ac/LLg
7wGtR2j4DL14ftl09Hu+bKDacvulV7kfg4nDBJ3Z9bHEV9aQjopXB3deC5I3jj/x
7Lj6vwxKQP3ZcDwgykFVMgnAmx/xyEdZE69ys9jd+Al6NzLx4bAwGCLuqw+juEv+
6VkyL3xlUChJJ0Z5OuMNtsaQtIJ+8zAQHzP6lxCt1+rYA//FQPQ22RGomqgdYq7v
X66hajDTz3I+BWef2NcG8Wy7Co1AyCPPJLbJzy10+h72NcPpp3erd7xJ49OzcJ+4
0j5SVznD7yrbgomrDq9fROFC+PpRtJNVkTUs/Xl8yW0+06k5aXzsYOHC/mnLHorw
MNPwKDmp6Ua0JbL0t2MxCgMEm6Q2HD+dbr2mF0BlfdHG58a7eGiyOK/GCHkuO2xB
6VlgvYhLU1kGUsOG/U40XHLkcZj+L4Ny2/NVmr65MmO1W8Omr1fVqkfyS26HNXg3
lrLudhEF6hjYDq6FecEdd/Ds9WpmiXMgbx1wC3/USa/dMPWkowDpqO65/XVwcQBD
kOPfpnvUk+5Y7QzahONyGuyU64lYSoX+gQazG6wSJ6A2WCGMq7EUskvhwPiAUIw+
hkhH3u8ZcIfyihxbeUJT93OEp7gFtLn9PcrnGGU+7e/PC4bPgZwN750gmYoyEcLQ
j0Ity3KiBttCKt8n0XdjmysYg7iRGv2l9BkmQCwLCz7edEqzLomYtLO7g1gYw13A
v2T1SRw6sFSvsHGwoByDTEtOJRSQFUlcKnaJLIeJB3IIaHIjE9R8WAlBTILIZr9O
6O4CoXKwlw2IEvZwFXyXOweX49CVImoNvx0UwwvuRRIsMib6sfcsJf2f2in9bOUH
780wUInES67C4LvX6mdRqlmduFNdWl94cRKmab6yWAGn+RABMebFhvDc3Yu1jufK
1Yzyv6cdiuCM2Itju8F1PAKbedewqLo3k3h1xqmDgiHSCYpCuJb/uPem/hIJKu6G
IW7/phfHofQEQ9L6x8whbK0UwzKJrIepbC8RmVn23/AhGFMHXl2xA8fAHoGha5tr
/nQtro6YbiAkUEXtp8rPQC1l+3qQ1wUjU9Bv704FLNhDnzPZYkWKm9fcUPC/E2jE
9FxZMDqBbfJkXYs6nXMMI4hDEyvaeDbpGv0JAxwUTEnfRnUoFWww4tcGyEQQ3998
x8tqF3YZ4JOKFo05pCiJ5SzhqbEOo4drecFG5pNJZ9hBNauEhucxB03qtY8GCAbl
n9yBpe/f4eGZ3Yw0oiHzEWnZLpqmqWoocXir1lI2zUQZWqUwtLK84oyTAe3R84fl
1he0Mptp/K5sxPoraCHIAN+ycW3+03SFSax1JwaSPIhxXRy2LvCXQ79EQATtvjDh
Ko/DeeECdM7L0bi10ssjfEq5P36hxMplu7DzI7wp+fkpFZUhnJKmn0jTX1m2yxZ8
e6FeOCuQQFD8kNt5+lTZ1THRHFPZ2zJ+evyXTA96QR2jwN3eLQ0PqxHXWxTMHeeR
k4Aay7Dn1A/280pmQhRFePylboLVpZibXhvRfBT9KKpAp98xYoLgG86V6HEKdwni
rvLUBuG5uprYOnbL4BXJdMijkrGoCl+/7JejZpU//tmSAu2xvn8e2NP3quON+dIz
Pj6dsXbz77sNwOcFDVbEyBhytQC4svEDLREwbMiQOJscbRX1XvhJK7oLkVp1CZfp
MlQeOM5vFO1jwqY41aCo4kvvKX6undWYy0ECBV8zM9igTcMUohs3J1QXTGYRyoWg
1qiZnQRveRowMNmCmVbPzE8rMf/pqRnXbiUWcSL5iMr7VVwUpH/pSGbqrziZAfHa
QhlI/+IwgbvRUMcQRbbJo+BXq3tDegWohG19mI6v5DqAP6eKaBPPaiNWGFHYwiBZ
2MY/7pS4uVQATgS7c22K9nAAEcTgq62BBt3d1JwMQl6FOXO8TOqU06oq7CqOZ3dO
wrD5sNhIMH81bjWkctPBeGcXldtsw/0Nu+fVRm2GItqwn6op2S2+ER9vVyR2BR7S
g9mNRYEL11cMMQs+Jmf4OZEKCyu47uPq5tPoUj9HBbhcljKfPRHdEs193osWnR44
+jpyzmeBx4sYGHVmDpWh1YYFHEyDTHiL0DmWuAJMcX01ys/MbfQLiPpUUwsqz6Hh
6YSsmbgUv73Q/7xE8BLotTfCh34Ae+VCw86Mq0i168GJ4Z/LpZWfTBLqQYl4zvEm
wA00GtiPdh42hFohjNc3Z9ps0DEUx53OrcbAqOmZnY9iqzMlLpany4i7kSnT7BwJ
go87YnAFoSFEzlwwcAr040tkNZPPD05uRmhJ8RR67JaZkg83n+owJbhEpS7WiXrI
kDlwI9GIH6KBglg0Ot+NzMFoeBIdXMXiVdaQ10hiLT/WYoVvuBojFj+iYWLLZ2o2
RTyrwOW5/isjj2i680liGmn0PkhKzyxXbO1EJbitN2evKUwPfCczPp3ViiYS4iyE
2EGmScYV9PMwYePXB0zxrO4u6YVJYRGyz+ds4Geo0fizQx/dr4UmduKoIMTztah0
hqE/wPWS6EySiVgObBFrf5y0QmOXGoVv906ZW3iyOAlogVFq5kstMavs37n2uqLs
pmbtkoWCE60e1VI8RXbc4qzK5noOBqRLYPBXaF5B8VX+uykm9qcI3IKu7GHdrJp4
JYiuNnuN3t0V7ibQCcDYnVvxsDSfuKXqZk0j6mAOuBs1ChMrd0dDBc3fOSqbiTAi
FpgShqJY73mOvTzKVLNIdmHxDEImoWnZBWHV//Po3im5ndoEqqveaTUtuvMq/tbc
LV66KHvELW3wy/CXdiAgHOGO7e0afJqRRc8h9m16OYdMryLUDSkZ4QzRSenTbl3a
p51ljMNw4Odpw1HIMi1qeZw613YS7/BiRS/cVguDLfurMVZqTDot67dnwJlhJ7Pu
adJhBPmyppzzbnHw6CxswSujhZ0AAfxomMNtnjLSdBYFfWDWTF9AVWSuLPhgw9oN
C5KrGhuy2zLQYcRodDqVEefO+JFPzWwFn4BjRhJAHI9/KvnpiHXx8C/arIcBa8kK
4Eq5ULCICfctjTd+dAx3D9WAwLvvQXCry/MBLRAQXzaXvSzp5CObWFmtykeNFRz5
QBzglhwijIjJZYi+NHJipogMeO0oUMNTZWpX5Q0albwRBCoj1YeqeOW5i+1FM4y+
dcHMEpGDU+X068nUe+zxM9oGl4cYyMGjY8ANNkcFpDoCgx3TEv+eJletHIWi0OF9
eni1dkZcrqHkaut7+biANZgvTk6et4+LKfeaB+yGxW6qj6Rk0kdt8ZVEj/5lGxPT
GTrsRfPlKNtcqvhpLeSkYa9+tMSe88JuInARVwHx9ot7ohgwm4ZRKYcJan+rBx3V
jk8fhblrki7NJTZa7eTcG5u7JhyXt1E41pkBqxIRykYPXp9zqjOFFzq9Ulak1PQE
+tZ/MkQLi+KTwp5elgX+ESRAUrwwpa5Yq3oxGbhZq+pzPYDDK9jjVgMATBzSE4gy
k58cgBu3FjZUzhloh0tOap3hcWUbF4zfUcIrfL8KDpZrY17vcm1OZG9cOGeIFnWU
0tcI8olHGopsWbq6Af4D6+hBab7pnQ9htuZET9XPupm4DJcHDfxgj2QK08G/Sbzy
YH8llikjz/qlvFqHn7zdPDEwPD6CVcwCbYjezgw9CEuzK49NOxvSd83OHvLRw0vD
31eHrudFCYazpny+F4zEzljVsb8/3TglSEZezFMwypjbC2rkoYb18d2+Z9BfxjHg
k63R3eWUDSqbiAXnT6wAD4lvOdGaX4Myi/Nwawr6lpeT9Ycs9PFiSDFwdcPoNtib
anxT6IWKle3+niK6SETwQVdNeES7xXZSB/MoCCUfk0d13rH+ZzfMnvcqz+q5j0PB
sn4dK93hSIjpe+QxpZzqrxSnjycof/SJbEcT6RcI2fv5y5LqiqtArWFI6ug8Zp35
8tnE00ICM5DyQaHh/5X1PV1xXQNzqkvL7374qERhxUp6vOGKAQdPIZtYZKFw/fEd
79Edpwaoefkl9RZLiVA5mQhymzD0mJzA6yOG1y9tCSEOTangnCU3kYpSLSAsRI5G
7DpycJCTWaCXbWoDHRvrZgjNavJiKJt6Q53Zt3AZw+SBDz55LwU8GJQw3bVIEAO7
a5VPatwuPeyWqlS2kMvnOEbHcHNwfyjk+ZYxEQXPT/PPangsFo+UMWWmMEFEem85
JHoEA+EVVLYv7tLMBSFHtUu+C+swYkF5vpnKqfKz2FMMjPI4UiTeWKxVFGAUP4/r
1C+KVd00sEpPhQg9KmQuq4JG8h50Q/PFyxKg/rTGhiL/Qm/tVvLnwWCed9attMs3
sals2/jze7AnS9VchAbQv0iFLpPrlfAhZ8sJmYVS/lyuI1Y+h0kzps5yqeBZKv0+
PK8/tFkHpws/7sgXF5XpCNtN/e8xtnuL+IkQ5UmPqCkxChlHAocLMLLVINpRYVEr
9X96tih+wu6JKI37olJZUclFu9ROEI7rh2ml+rQQ0eBcFVJRbxfaDiwioDF+WWF6
B9MsN8jSyOnt7ZoUCYJUpHXMmp2H+eHXsCeuT90HbH8piQ5gFnAKVK4gq2HhYxAq
5mFK4VcNCgUldnDmNCyrRaZCX1Qn1JFyoyuNSq8XiuFDRJJNBbBIqgE9c4uIW5Sr
R4lhNgT9CyWOTmTI5o8fIod3PhmRFjwRpZ1RTYQ5rOIH1/e1d5fUl+NjwfRUC5bV
ZuTtUxQ5YsP5Kcl00+ase6iK+YHjkAcjhDeBWsO8LG9POWwzXaK95ECiq9T5SAi+
/eSpbzciMVB1UrlZWiL+HqDHvBJGVeDN8M1fUYE8sCvvUm+6wYA8y8Mv2vdYILPx
K7Wx3uks8/+QGlnCyndGzqq/HSYWGunEllY2V5JYIlQnh6E8Diz5p7MmfaODuyu2
kEP7mX2xb16jfwDh1kJwTAW/5Sdteitey2EvZXAAM8SmHmBlrdTRzpmcJCJyFDrZ
n1S2DDjqdzik46nZ1i0EQ5XRzlR70HmVIjx5kQuyXbzpwNDrRObrMupACaHyx5dx
uHvU7cj/xTy+P5p98qPlbBmP72HvLktDqqSo68IrjpmTZYLqXRojxkVq61FGIMmH
npyyhFKfsE9AWwiXcebdd9UZWU7eH6eLaVIAVvKlqy7hlsu/WRZ70TxrZygLwhpj
OEmkop9qafLwrxXlId6unStU67p0YYlefhmUMe22oehHv/wtOfcC8INat1VFM2To
vAgCSHHPfc3iIapi8SMH70fPjpA1iaxQH7sOkj/uBkNDvd0ljHrZfqBDz7t0dPfh
b8/lMpaqyXz5eazkzWga5x2Bs/fY28lzhYVLB281bRddp8apTLU3rQ7mSGTIrBFq
2nHvAEaKIpEKsebGu6aBn4KhQTpg9T6sP7UUruozUUtdKarCQiEVtngmFka4oUC+
+h9wGw6vZiUKo7+ZTVlhsXUTDC2CkrIybBA4UqIuyqSYKkX3xb/MpdrY70vg/d/h
uzsbHZeMUmHlZrKToP6wTNaWYZ8OSGKgtvPAkLiJY2XaLN9NVk/SBe53kpKJm0aX
pwflanxBFcUHqieGd0b/PWQ4xdoEZs4wZ9I5fmGerijmuVHYVDi2NMM4pljSlVQh
EWXqKF0hGYsd6sRlZFF1KDF3s74gCr07vdMG6ASsZi/ih/8XyXaMwaroheReFZMx
qR7OdJc/oWlqKvvlXRLK4C354fxST31r/JLuhGTx4fl623bxkgJX2jBRXnJHvg2z
4gSOxO8ci3f0oA4v7BGbwqyAnIuyxdXsAgllI2A0s0Wt0UT8cNwU1tra6AMr3yEo
DXegRyBDuCGDAP1N1x9aBw3rXAqEwZVQRGshUmfxbwCWK4v2NkD4uroQZBPwIcWX
s7LDqcpdWhyuIkGxTkdc3VQBG/QSSIGSao3GlxYHKpf8I4bINRoISq6atsxuhUcp
ddiPsSfuduaAPXQq/+eUao+UllBiMqXKLJbloyu5tTDMzWt+C5a+I/jMBTRj6DqO
UQbsc9/gM3PyYm+V9LtmQ9y63VJFvrzvFJHGLoXZz9ZVtWU2QGJ4PFZbnP8oM7AH
Cd6yiIkYf6UBypN3bUEh66aiZXnncG9SO+R7Tva8NShIyCIpgjdtc4tqWC/Q5g4w
hp5Ax8yqEkrKUsdoK+4i+qVogYjYd/FN2KRiCmnZ+9WsuRASGNkz6mzH9Q8108wJ
2oC+YvVR4ygnNAiJsnjwU67HNHxo37mcsgFzXpRBohtw/h1/d6Z1k1ocY+INNaiB
eLDiuu1q5ZPmPuG5TSiT0zY2kLjdggd+pQE8CYqe+WeTQ24GIwjM400toZGm5idw
iB0vtrRnYI1qykTAJ2gyLy49axA8OJPYkfXMStrEYlfNnbdzigkRd1/MPPao1K+J
B2ojwNm4my3RHJKY9Sk6byW26wq7A1ndFN1QjTLVwtIP4AGHl8SDtNCz7H2dbI5U
8l8UwWC4PwCczaAnOLlVMA40V5bqoWyiqyB5jqPzKofdG4RCWMYMYrUJuzNLMA3f
E879gPKdsUrB5L0y16dhRErMG3SOAGTFQteBowATGVWnHzVJBp5So+Y2e5BkiYDj
/panspUE1ilNyI5iyqi/Ki+c7cRQIWU1j0E8fCaPyAoBgwfhGov8fiS4+IcJiuXI
TB3npcoZIcWHDJEOTxuiJpPAE89EDJcQIbFtj2dtzlJAqjA5FoAJSXztmZdEkBjc
+YrbWvylQYstCmREnumekoHE02Cv32RGA77b4MJ+73vqmxfkhLOcZDmvSSAWaleq
D2hFL6oMVKwufFgsFvpos32B0+Cgbtuo7nHO75WCjVyqptcJYawFPiXPfkBmsdwJ
gQlaUeXSzX+PKe3eb4wfoV8SYdV+/yoF5M7UAmKo3LdaT6DHV033MxjSyzWjN+Ik
3nIAmRD5S+HG8vwEv56vH1zOlXEG2lhQr2F8B1e75W5+KxLp6lNyXYNsr5DHK+hb
ue5zqNPNWhQh9q/0b4KAmHe3eTDEGjIRP9t+0KQ0CZsTnd7UaW5s/2c7+8uEXNMm
qxMnHVUfnIIQoI2YK3R4Qfg9zmKF4qs8V84S4/ZSk/S9x/GisGf7doJmeEAWDJsJ
mT93R4cq0CNCtQ6OPnEoePTN7JYzttlcSQO94e5ISQiD78zx1ItoCcU86+YPDzU0
C6eIH6C/2fXCoxeQCmvTPFphUBvve5tDplPb69H/WZd7phnjMaFRqhnpf1oNcT9l
oSk9QoYtrGaqjUjfnYjFBHFbw3iAQs+/Gnrz6qo/VcYCsjbmRUbtDlvSK8CdCZyJ
gNpLa1Um1r8XSKBWX3LuP01D2XAQoH82InwUDQOnbvaveLrT/zxEX7aKayyExQei
UFOI0U+GPt5CQvX78QvfUYmxlid2zwCpiDoCGhwTQYl5CFCK41mILqdQmDCxqGFy
onyq9CcVaBrOn+rs0KRNdIDhShYqqq5R54XN1HRUG93HLw4NUxK/pZwDMw4pBUUl
RNXk/0LxR0/8UJo4TwL/ArFHYjtew2OpZ9cujGuk9YTMcHcFvR0CiqLJsjEyYKde
+grkKyZgcPEMHE7VAASJ1ZTskigwFQjI/hwHD2K9DDSOC5VadAlT2TbB2ThkPN/J
jvIn4A6Ain1UUpR8yqJxR0q7BbYSfvbQI/1f/cyym9tdwjUpk6UgvHNSKoBwhG5i
Lw1Wl5FUAcwYCsrCI2eBgZphgN7+QCDb+uLlVLrPagmiBuxZ5hDC/iXWeN/HMZM8
9x1gHI/yO7/GfwnFxwvZ9v3KiGUrkuZAtx9d/WcFsYvIEqusgX8Cr1pRDDSw6Pp9
IUsPSjO4tyzS5cimaZmAoZWcTZ0nEVpXGUiMLQQV//cOq8WR5SOt1QTNgcZtdqjr
YcfWWlyJY9dfG99oWH9lSyl44TM8WW6ZdV3ENTVE9YquvlGQumD6hQLe0qAoEQX4
WHxapx/+9P4SbH07JpTL5WFFyAjh7hc4Ju48fEfF5NpuZfUlsIkjnr8pbz5pHpJA
FDpQASsyY9PeIuL0jpQzYLlRB+Zc+NvfRBrwjwFdRaxWv8XK7/EbrTvXpsOYO4Ea
G1dkh2fEkqhkal9fvPqa3li8bmDc9FTRkxWtH4eFU5TDmlv0OoPnkPfEP34LtlLH
Oxe8/sgemO/R9YdTPHLc6TbJSVHZkjYtVlRHEu4zCF9wOdCvXBdp1o1+Gzf2hvOP
WqDpNDD5pRyfuQIdXNWLCOraJYCU6sxkaCv8V7BmOo1E1LPpv8wmsqaBvHqJ3luq
gugV0qTE/js861BDre235EdUPr4nkmooPMlMyddEHbFTY7oEaecY6aeVWcvza8aw
v28mfDcl9QqJZEAySvkm9U05NWdSCg78HIipPTlc1bAmfwo9nQFDlZYJ/Dw00uAa
W2shKlLrXTaAvlEO4K8oFSa1AtZekNzpKtweGrEpct3hDvjEzXq2dIs3DqJytQ+A
MJSudqoUnfbzFeQ0Pw+zTCldkl2tvr6i7Gr7y7+TUjgxVXKTnL+Xt9QxPbzH+eK9
FtQ5WPAAmMr47sRA9nb6DAHx0fe/cEcTkH8s3O73wh4zX6kxt8+ZjEZj9gcF3nd2
pk7cTl+QHQWo6XOEI4zcLUp1Al9pbAqMrkwRheVpmdlQpO+RPQOqdHwl57hiQe9r
Nos0BuKQWkHUlApm7Wm8Q1I8tjVzS/4Z7tifZusf7dRgJXisIdCLsoknaA1B3vYx
PzBPmx3x31hjcHQplFfFL3K4yR3PTFT+IVamaVcZ7p6vbBAhTOI7RJE7t8VNS8aG
PyQYmFJigUDtr+dmPsO17OsVmolgYelTgGdMq/YLZAGb2pyUR+yUnUm/w/k1eG4j
8RDaAaHNDnsg8A7LR0gkm4En8ZhVjo01IWvktGgKCu4M/32rmbQa+R4NCUvUThkk
BfB+BRnHON+YEbJzvjlcayvzMZ2PSSHNkerN1S55K1/1qopQoHRE2bxjQRWBZfLZ
zo3BRzK62oT9ndJH4WcEVvLG8vkJVGUdq6u8uMXQPrwiutcgGR4E1mIAiIIQdmYp
6qqZHZAP5gwI0B24jyUwcw==
`protect END_PROTECTED
