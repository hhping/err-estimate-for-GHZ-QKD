`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yywor3JpyAQG0Ze3qqmuLEb7CgY2Qac2q8V0pN1LbFjg3SbguBk8r95cSpnN8TLG
gkDeWO5dmb8VbZNuP/3TA/KltpyHjb3obEWApn0XvFqOGG9Ki/kzM3qSEw8Hcd9f
5OnoJuHYraLSwp/rSFA5hY19Gwb9BCZSffttfCfqCZxSj5LUqs6jIpaXpNrpXY1E
EIgdtnINT6h6STXveEdVJvB0bBGWLqVlJmtNCGZUCE1+iQeSmoaKZWJK5BMCuIrs
IX1nI/PclvCBsvXXtE2yYSFs61Weafn1Kn9/TB5q0Iq0shjIKTqZRtqlO6RUcgfV
8l11QEnG1z7wiaPahuXhoXbTB9NZgSCbPDE8F1kOp9Ok7+Y2tjfkJVPMBVSM94Pb
yy1dqooNkO9XhY1c9adTERU0EgQ4zyqWaAtBV+bHx/Z04rcUaxwiIzATXeEmB3sw
cKftwoH3ttJDCdQCjzG7hrqKRfVfDVI3s5B85EzOS7dGjkK6WyeyjGOzcRNLnNNb
C15JBcDSWrbiz3U5x7eR5VEmzwvGrzxd9p9EOZSf/yIndtJi6z3cK0Ax3ZKCaw8b
XNCaFVXYheUdMRdkC2IOyFihiGIXlhv7AXSiwOMLiExxb2dWJhs1uqey4X2BQacN
/CkW5vlugAe1shYY39xvHboCDnoKudjUl318AvLtuuZ7XlGguSBRTmOqpYmm3Cul
ozTfF9hatE1bp0cUhNUcb3UL7slBIsqs6Pox+dGycQ4J73CdFhwjKFxTdVfE29im
ejktbQnLafCpDWLimsIyE6LpOepIrt8Qbl7hMRQz9Uo5BP/o9Zwi96CR6ZmPtwyQ
Notf5ddpm5BSBHcmmO1bdfyTVLTqF/W759DTOMhF32htuWWRIrnqHuMh7w6r/Ak7
8dDhxFIWHcelu3QApcnx/i3HfkS8NuKXINQlFssnC83OEOX2wuDu08IkTQji22Cd
jbJIeV9tMXJuQfqdKJCYPnUmske2koEDpjV4OAL8Zt5jPuVrf2bKDHgKP2whQFk3
fNBuLoGbhs4+BleRHiaceRPcr1dEeQTP+3wvKJ6sg/TJtOGFOuvOI3aPXWEbPLdd
zVnvMySMjxzCyXEueimt26d900A8fduEEb8/K4kNBJ+SEBfNEc19ZW0P3cbjprix
8gPyRGDwBBtrrX7utC+VsgK4T9nzvY4lnJSI4nbEhZ46TRQh7e70pgYndiwBvBtN
tlQp+neByLLAhXYzXC16VKaL2ae/1o40DW3gMPiSD3UD7cDSje9C6ILCUEeIKQz0
TL4YZ8xzZPIe8spmYqwiWU2vY0sPOLFszMIj2J4gd1Jx8ldx5hJM5FEfo1Siwcs3
r4OarIrtWA7k09KRbVKtVbb8IF47ieN7CRTQNCF9pPWS9gWjBkH1ZrRYtNWp/iOV
myabcyuMIvYwokGQEvZ/zTnHpGuj99zDBWSbXLJzXEtGmk4ODCCeTlncSqxWte+H
nXVuT69UuOwvznWOWha6sMsAMv/4nDvjgsE2aY+xjPu/pmntBxtGRVjaipe1dfCM
kIV8RhGshC5IgbMaqOTTLdAhwJnbiwcNzJtFlGGtpCmIj2Kyipi6xlFiA66HVtJC
ePGh46abqmrGGS2emHMh8WgQLb0/1L+5CGEdTzZTsAgZhcn+18XO0UryXJeXfnhn
JP3uVu5foqHpVmZEKydayGwyGcBrI7FzT9AufJB6ZhY/lZXB9Ep3DBhdy3qmjO0W
ux4yFCgpDJDrh4ukTkffB+hbCtS3YMr1mfzQP3K4MLzKHGiH7JxBVdULUts4vs1S
H/ZCAJgczKdhdWgGY+wesG6O0tHAC4R/RicQUO8ln8nGGsGi7FsDfzpKxE+Gjghz
9e4gBLn9ddEr5GuWhBz1+yYfqPsnKYIjriidBOS2SoyRNtk0ju1Zkuh0LMem28mJ
6Ani7hforxZjxTVjFwozWDsf2B6jjqSe8sVNNsu1G4TDgzcpz79pU/dX4bkxgJJj
uqUJUaCBNijVtSh320BVquLZshQd2L6sWqwpqpdrVp4OEpQeb4MlSJuEe8sn75gg
aaVoBbY4iQblZS7kYWQNgg==
`protect END_PROTECTED
