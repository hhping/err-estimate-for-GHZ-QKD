`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IkmD5zvtBjpCqe6+NJUo82PiAfN6K512Q4z7IJpctDIQlPUZzGfTiCYdzCONJOSk
7OV7Ljf1DkgkH9ihfUzgzWw87xbME0hOarFjVMAD/24+f8JFa2CNq8/A3f6FhHtz
rt+puR2vpHyW1HbmuZ3T9pDEaBZmB9iHUuwAkMM5XLGHH4WE/DiLypVXeGLynwCf
M/R3595VNUnT4L26nVRJQ4ir6OMrMli6JICsyb3hMxCJf7ILyF2ffWhlpIF8rDJQ
jvE4tdjvoW4mNlQ6HNhr7BB9d87CJB/A1Jr245Tukk7BIA7nXhaz7wdC1qzbAMc+
EbGkG6/UfHtv+50ZYMQZJJfriWnRFP0rvuSw5KnfWl315WhzDjhaEldNlH7b+li6
VwvKeqXN7z/aJqBod4tdO/OjTtRNprxqkH39FpI9tg8J9IFtYoRlA4Wje7qosbbr
FGi+XbREeYDe+2AnduA3FYHmNd7s1hAJ0pphNctgK/+4aVAkM31ebF2m0HHZv8LG
K7v9GFdah2CKSlGa0+hJ1eJ5ODPsNfyGdrNMGxf+zMn9RjT252wMmrU6hh/j+DR8
`protect END_PROTECTED
