`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3CBgrjsOyQLeIS+miKRkOD9CL6nyr5F2q2WeUqRmINBridcgugNJTjdxIrtWXEa
5WLxlqJfQmKYuGDJBt8XzBOWThjJ2PpqNJUo9gSHGU4ZqoNWwak9M0h12v3ULqdl
znxqPDv3n2io7qh55yzvzaARe/2dtVQxHCwN4ACwkHq+d9Nm3qJT5WXpAoene8xX
cqHu1jZuYMsurLvtJ/1xfKxltVI2VSR3LgEZytW5QwaefO84Dc2XI8Gy3dxrEAJn
/Xyzs4Z9HKFAtg0FvELs276S9h57ZtHrXLZdv/8J39ETL/YGG1DS/5LuXscke45X
dC/uiGfdTK3VqDEGfccidMMV77Eoa2nRP75K0deJx1hS2KHorpKubhF1D9l6rg/j
EaII6vwWFkN7trna7HhlsU5ugR+sVv2eiYvhcqTwNLovJFgNRr0h4dj0h7036laY
z+h5ITJPS66TMpbrTBtwI+WQDV2qYgLuX+t8c1g5aOR2tfpwMtASyyoh/0ipzlrq
Bm4edKs58eFIMJeMpX8fyB4Pei3NDRLgFzKf7dMIXyevD2bqzMLt+Gczxnre/XZJ
LacWmajPCFpAWgqypVRLY9tmBw9KdTVgvQc3U6gGzhueLsUzlVmgaPFrLsfbiQ1i
KYgKpZdV3pa2cRrf/hVWtaF9MUau6vUMxui6waRUbMB4k19DNHVwIqXQgAAc5Zdk
g/px9rzMxKRxwIj6JJDbZOOJJQ9ixxFvagZjrfuC//ZTIBuWQEKR1lnd4+Jr9t+H
h4d2TOOCgz7yVGMS9Qx5XjfP+aZM0NruZ/hQx6dxUnZUwEVnEK1jv3mCNbFp7a9S
l9xQ17Q2HYj+PUquDMvwDq6Pd4V8diNeEKjTVEBtGYt0+J9zdXvA5UxP0VDVY5Si
beGKM+KsijR+4VZhPW6bgo2morF2efmAb9aBlZ0LTU8ntuJcvsAdPDsJa/E7QFW4
mw5+7i1/qB3iZawVXNGazvY6f12DFYWzR/tv2XbCaYz/SaSLhCJSymIEyMdDCjkF
fA4Pv4zaEhwVLxMTdj3cKSRQ3aSrvBv8wbqU/wN/3US9fgPjr1ibrqrFsMNQdA29
`protect END_PROTECTED
