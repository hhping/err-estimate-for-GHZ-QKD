`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JAanNYWGfJTH8+l6Ng5AFGAHfx5wN+++pd9DcrDUM56k2sXYfeL85oh0jRVvDN3
nAUjoutI0sSFCLbyBSf0xmLQ0MYvhQJufW7+6meLa9zwAkKjM4UNTrnyaW8U+us2
0qSfwstoTLKRlcuo3b5PdUJx/gLORq90Cwyrc9yuwqizRkAn9yVTGSRmC2GXx6d0
Hu+kE+e8urwECTjbsNszdeDFpOlUPGI/2I1rhIbdgnY3TQIMa3HWZxL83zvri4Fc
CG9XMjRcD8EDkUiPIplB8akSPrqg6DIRJso6TsX7rzJCUwnn1mOxUPMeK4b/pIFj
/z+CplugEL0o2cD0kdq94vEDdKqtANm4O4dORNx44edb9x0yoPHlxjN2DRLUyHbU
E/2axYxPiKwTI/A0zroBhRLT9Ry2ZSUueCzz66FX8AOp6xwoj74/T277J5H4kQ/S
hXEhWDN710/8EihDvyzHyIf6blY0xDTcL2tOIzXAg/feMOQPAzpZto0U/LLG01LZ
iIdMXj10dj1GWWp3fdwRkRHuPC8X3ZaLIt9z49pw+qo=
`protect END_PROTECTED
