`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrVSMkrM0oTWxprifl2T2dK68dIptVDDbZYT/l2/l0ARTX2z04+sReTwPPbcti38
eONKOT2dBlzNnQ5enMGwsSvp0PIbWsN0bVpHCJn6fcdsqgjpmKEcSpB6Sx8j48Xt
aLZjHGoIDEQKEiohQwe6uCsoT0UAnp5Y3wYP6/4NAGDWj3S6q+CTE22E+iC3zHPa
CEoEGDQKlrEdc5fnzKJPst1g13ls5M79+DTKLR6sU8wYOX/xZEawZPbB4BH56D1K
W5WnCi6ChtaitvYR1wq6/YFzc1xSHfvNd8M0T+loCjHHojVdgfmEavEpxzVTvPWK
+ZAz4ndiE+XRI8b0nyyM7NoPiFQXsoXX/ZhjXkgR28uBJU012b6muuHxCAkl321P
F8yEWiQARB39cictfs8cRi3iWjKK92kM3DN2yXn9hxa102iqzarhu0S9uRWczRKb
nokoKO5nG8E+4sbFD9KqgVvaQILhV5yHcD4tvZPazfaLe5r5jYYZr9zNEAANN3ZI
yXyWEaVgeD/mnwwXuUB1pLk8597Iv06i2dcUHXSjLwuk0Gs4qiImsB3PL077k+RS
OufoUIA0IQ9wRLLm8Ua585lfQ1XtCvz7MLqIlGD/tXagIrFVvQIpaRNPdiPUj3zk
0JO5/Gv8E7qRazWiYjGDvbeoJO9k1iC4SQJl+/4fGooZdZIuhm1j6Vp1EL7dVBtX
k6jC3vvjSA77R/NAjUtuzDHn9gAheQCeq7P7BEVORwwLOCDpm9TkhdQHlxU1oorI
G/osC0IInI0/Fy0LBzuVMY4MZQkPvCYVUbL/2oqv6CAB9MoCQBE7HyVbNtxe/mOI
Km2bYuX5LPJc8fHXirYxazHOAKmNoT64LG/4VEVijRkCZN+J/k4fwOf93bBBdKXg
DAknbps9oUMq5EG7/YattJRnCWOXxy7Tvf55ku8Pk5xnrfXxtowef3oCdI/A+AXa
4fzhtwxMldblvB7J4oBdZVNxlcF7+yZbzjIna/S2qZI+wIIsNm8UsfmZA3KnC7ky
ed9YzQfZ9XjAR4VRJQSNTlHdsxv3yHVgnqWxADcn/bEyw/ir10WtlxXdNCbgVmXp
9FWPgdEiUgeG5sWNxMT/odEl6LywDb5nGoYIYC5hEfWpjCd+HzZCc9cWuuqkAioT
ySXkdPWKtXqx4ICquXFWtkOvlYcSDrlKvQ2fDq+cVf6q0LTKmdRhCbJIC9Ye8sdX
TsWCULYd43CO8wOeAxWZ+eLSUuAiUQKSo6GD5a2HQ+Vkfa1Hzqv5mnYk3fOTY7vv
KsMidh2h+aAjBsmGp6KzydBsycCwDt26ttq28nQYEW0Dv2XMqD9aEUjS/aZN6DGW
GO4ImqzvE2Phd7WvCmNKKliNkp7IrWiYbYKE8Fu6pwFyXGCLCJXBM8TSF/DWPM/h
cvKLhZ8tRrVr8NE/VLGl/MmOex50vC6RW+Lepav8K2ycUJZOCDfBl5jbJFDx5Lqh
Fijk0NeNi86M/LSe/fhP/w==
`protect END_PROTECTED
