`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxAS6MeDzUUdHTsykdgf1khUJ7rFno+ziaoHwUuq/nHKq4K/0qQfnefGnta+E33M
XTOCnLchFZ22N+5nlMb8pGn017T3kPXFR0Z7w7IM0Qak/EvJRKCISTNRoINe/MPH
HvPu1OSdkPUwGc4xcLOAkG05EhkHOCCLd85ZCHe6OYwj8qmR5PWMgDmW4tH/+/jY
aRhqo4M/ybSKO93t6KjZTcd2bmjDFricpEEqtunBiFgqJsXdmbd3N9AJ/5e76Zmd
81WN9FaJ20AC0xCKFAcqxBQ3DhuBduOSGpuIjlY5IhCpgvaGCfftPCdUwezN5ATx
imnhHgLKqHqyvtpKYfb7ZAAOqywkIavIMxwUFWMeAofpiFGxuUWV14/77zMMN2de
CdUBbxHwwBjjIuOklQs3iElhHAl8kW1k2kjZrMle7U+LlU0wp7OakGY9eLupRugV
Nm1HumCZR5DN+juUrcyBclXQ6ipzFjdYwYfEUTklfJ/KhVs7qdLr8qXmR8Hzy984
osyg7y934agjD66EAAXOFz1DCXFV/yneN8u55AUOwiil5FZetnWKSeTx3Mw3WX/8
p7CWXNZct7dLXgcDA5fhhSgVQvbSYg01gJzOEMcso1smpvN0URRKI7it95W8YlZq
Oi1/tcnbt3Q/C2FxVzlw2xsUvF1eWc5dNAIa+bFr5c4sn0Z3LajP1PjCI0EU7GJS
qLsTjsCM950NNS11+FzcLMHknvIv/Icd6pGWDKmpPuAnPaHyTCyCp/jLB/l7mgbZ
8RCYwkjRvF4lTACYei9IUu0WoYJ7Ksh5ArexzDFo4gDlAnZoMjmIWw4ZPyG1cBGw
UuDk4gWx7PSJLmNhLi4KjGD6fBkSijEUQMvYKpcfNibkRJLrHB1eNi5Jx+x+RmtE
n0+IBrG8oQCOVYjvFj/O7F+xqmnJCunSH3Q+rhRqLJMXf58EXB+KM5BSnko5k/0Q
/0gRSvJaoBkhzblkmvb4RUwovuc1YyQibL7xth0uM+CRv10NHyeKXaJvMJXh2DG3
6N9hXyMzgTS0wTkc4SgI/ChaVUAnksybGvD7WqdXQN8Wyi41FPlcN/+vRLpYAvp7
GvgVm/wDbBjp2AB2c2d+Ik15DiFRp+U8BRgMPDo1415hrE8o9bXl+ApXSNTdm3W2
592XYI1znvmK6iARlv+CBxErRBJM1OOLa8LFearNYOBh2MjoYE7zUc98DsPogMcn
x2vFgR448HqLGIZpHrpLnLI2+p/ZuRJuJKqUtQQkxplh7rZQ2WafYfr49auY+kqo
VwNuaSCREHBmTOTWYH2wx4K5r+4Y4Z8D+nAZjyt0anuVWCtoZd8igKcdK6sbmbmr
5f5uJCRrYoeKNEPYQnpmmCihgjxlheC2XeT6BTvb87LjDt0W87iiV3t0lqb+JZkB
3eu9iw7AHVKvpirWq9EZnS1lK1Hnxu0xEp/tY6W6w/vKjqTWychdK6O2iuO6Pnp2
34qR4nEmFphh3eM6Y5VWvYHQJLhrzgRtSJXICTdBW58ijEF7Fdmo4rQ95PYrEL60
MNJVjEXuTBKrb3vV7bPLYFkhdsrvuNXVEXEzA6LnL6akploNw68YIo1oZyz0vmBr
Y3Ma4SIQClB87GCtVxzc2yu6R3WslpP8VSwiWhy6OfLgtY615zJkKKJtS1aS/UH/
VECFm5YuTjAjSxjHllHriin/jtY2GJUu/svdhR1rqNEIDo3X9KazSLLh2eRDeDSM
sZOLCpbpkwHnln+vOpHoduxFBuuxXg0DI4x2b8EZ7fnCXFadfAXM5jLC7x/xbnBZ
g21Zm1LsE78yAThJh0ZOY2w2GA8vEm90YoQ7GhU7IbxM2DKOX8xFOEQibD8tmyw5
sIm4hGtib4dqQiG+fRqZQUR11rD3FqFRgAmSdmQqDiGovs9+lisLdZEraGiotzGk
DWikgPQtYY4zpbb8Mw0Mt4U0Jw/Ur+B7m24or7orBp7PHDtViuElfrTKOL7P3xOv
+UDeu6cn18euCZnquLTJ/wUVGUAlnn2/QY8Da+0Hsl3F7CxiFLfRUwA2YAx3L2jE
1c/s/0KhqbjszgX5FpOmhq0x00VqvLnvKemS69Scp10yQQytGBpSx9k6ItXI4OJf
72AabmwoONs0AmyX+FyxIw==
`protect END_PROTECTED
