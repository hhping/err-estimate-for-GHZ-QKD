`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBQf5efiZnTPumSklaSkLrod9N0Jx64Hej8+qv2DO68MIiCSdmhv0BY6JVzcesl7
dshAIrfTOiFPlER9V1zjl4St8ZK6uDuRWpWKP2WUNBzu9q2AkW/MN9vYga15K9UA
Yjmo3ZHq9Ww0Z68xBNqBg+N5KocXD9maaLsrHFsZ8HppKJEQvs/TWahJroGH9o7u
OI0xzFI8r0/9TTQg1YCT9NqI7BK6xHPk8Vd7OjIfbn8uHiRvr+zCTUHA4aCS6VJX
IFete3EH+B4A9p6cgiH0c0r64zA+0W83qIuveYKpNJp3zMKGurC0IwHabuAClbyX
cBwjLeaW6fvWdRawN8qgJfurAf7H6N/AIbESRWf4AQlGEZyGE7s/dyRxeLxSdn/j
SPuN6He4No9TfXwG1F5DZMMwSRTeBmavJ/Xu+c3vlH1b5e/KxxCnvxnwOGnHMsow
uSOmPrIp0iiNv3KbNogHPnoUApJLCQmFOg4ZE1s0UzsQx679whXGpU9kZ7s72/zH
JDhoCGpmdsQqjD69esGVdY1fUQ3iOrP8duKmJGzsSS3GtnW45reOK4yIvEClG1Ri
HIZhJNF6aPlFbMR1zHyfjG6jqmo9yuIjwXV8ymgLCei6jLW79dJ/1MiBMydcGbH3
3YjcdQ6ZkAlPLz6psBFjPQNhdoaQAL7y3qRASUT5vr/7ra0dXUm8oYtBJfrjYDJM
FaRU8FXOQyFd9uAUXhQfgUBqmcQU9CcZQc4Uz4MYxW0RHuLVJOg4zi4Gn/x80ggz
/ROjq+tCj81RdvY8gMH6JkF7Iu+RTg+uL2qLURxvHID0UCfo3LtVWsGpmoBSt22+
hpp8gYOYKWEMpY6WD8hC0d+Px1UgHkeiR7+Lvxmr/PQvgmmOmjzWLF7EPvjtB5ue
6PVdR4fHApDmyGg//rDn14gnnlSdSZyWr7qThAx5QUhmnSQWBZ/SYzcpXGiAJrph
+lC9fOF0RdkH1uLoD2wRXla7VkHulDvf5NaKaqrYovi2HwUkUj7lodNRdzz5DCUm
369BPdakOYK9vKrZRXFfigYvhuuNXm9dmZqwIXO5nsZbzaPwjlnHbHJnBSUvrNGe
HpmpYZyYULBuNiS17isJkR5SPI8H4N1y1M0xceHJ01AVIq+1Ruy0bWeiO4sq1W5K
VUjYlZWMktDmkUVRf+Wzij6a2eyLW920CcACq9p5doX2QNeQHlbUXxKWEYrt2kEf
CXCQr2JcZhDFruWJWYfa4DWPOq7w3UlUd/3/sEOQ7g1RKcRsOSDxT0iJCcOd3vhG
TfNs/ODNJWoftS+n4/gKP+PTXmwS99Vx05rdfapDdyL8iXKOCf7//vI5CODiWzHH
`protect END_PROTECTED
