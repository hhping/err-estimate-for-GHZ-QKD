`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YH5gpL11PxjxFbavz3qg7ilgUAJgXrjMMyhP+cQsfEXAYICBULcdu1rnhrls5jYD
dZuXQArHHkhNEq6I2x6FczaAwqanGP1IiTWmE6dK+tEALDyHT2SH+bIXcO83L2p3
rSsuHAk9B7nzvbXpcuW6p+qge2hMMDHNoRQOX9Ya69K5y+Nswwr7Tme+VxRK7B+Z
st+paAkkuHm5vt00OXmgbTwJ1gzdGhaegroV+HligJvBcmnLyWXtpRsx/Pw2xrob
ZPRzkAmyBvLobmv9M8Ez73EDwkorrMHvYqUOkXHR/QS7ttnB599JyK9EqqTRh75R
30Qbg9vU+rwhTNyIglYPPa+wg5ra9S4bVqL+n3TUOfM+p+9OuFROZc9xFiAEMBSX
Q5jRvddczOzIfkFd43NDrGe7oTm0Tt1/8/d55DeFdNtt2aizuz0omWa+eDSe4PNq
qr2pVjfbu5maSDGly8Q+5+Zg2x5p/+wwO0wZi/cjWO/DsPdi8xC3eAsQoeafUSA6
CGiDpt5i834YW86UCNpTGj0OCASGP3TdgWjZZW2OaHEz0Rt1hjaQiSWQ+QOF341I
kM6/0Y3DPJyHttZbo1GIHBARoz2cdBSOBV2uhrDS/aFbZg+cLKExZaGn8OdNjbgs
gw3j0JMyCMH5/ad4UGRFmGbCmMqbITK2q4z0w1194RxqUdQTOYlTLEZr52yrlKq8
ZLh59rc3JCPLmI9oh1NYHQ==
`protect END_PROTECTED
