`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1CHQf+oNQijVOEGaTye7XiSfHjo5DIdjL1xAXRW3rqDNyvgeZA808JX5fwrFTFY
qRTQz/biDg3LVQ2+fL3tUCk+YWvqfPaJTdOHfCl8rBoRgcsI3j6rMTc0+3RCKnGA
w98QgtXw+gH94GCmK+ObEjGSHrZs4YkUHiBfr0N5WK5IK4EKd57ULLH17R0y7K3I
Viian/FxRouqgUwUfmPmA3KPfkaXmV5lkoU3DRHuzv/TI+eIm2ul/pwe5izeZ07r
SkGAcEamhqTwYKSeXX/7oLDfrzw2fIsthYuqEvMub4cRv0Sxr2wc7YuZ9Jc5k6dN
S0G+ZAmYQ/CSHRGmevzwLmplJtjn+2HvMgpcWjdY8BEC9Xa7aExQSX4AaCSX4ibj
mYu85F8mBziK8xXHysIhThCoeNTFKukdBWmEE760qCflnMkedGchQDTWp86Rdw8t
dSFCNAgKPFTQE+WUUoxwqqoaTxZ7/Oy+gkST6+M0e4DF72Nv11x/DpSZqKGwJPP8
gDPTbHIrJJKfA0sZrBFT65mj57B7lAFOPRI2mUiDcldrhPPzB9MQTUpoQLOaf7rM
0Gc4CpOOIYmXON5fj+injyDfsanBFWC9vLeXF6ncI397uWFI+3ugn1izIfTkERwS
2rmwArRvP2tyL9BhiebrBZLXEdOavsenOecV9mjatT1Lm1yQSLvuW7pNSygT3eQ5
T0IROjREZSoVP6Ci0nJEuQmAKnFnZ16VeySpMDmZvBxoAd/5dRKJNw4yfjghtols
hJddre3cIhpGpAQRC11wKXgqGN+Zh4U1/aCaUiWRJYmfDQOr6CEQEQHWoM3Amcxt
sMFHBsmGtW24JPNEokQAJSUH53GP3YGxz7AtY9jQ00EimOqR5zCrmHBr4e7ohnzV
3x2ibi1rjwzzr7QKA1n/u1TJUOo7W4HmimdDX2e06A3RabQd4ZIYRNYm3yxEoDZW
z51Jh1/TWBnJ8sxJ+9B4GA==
`protect END_PROTECTED
