`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNLu/iARtIAu6COIkBmQIX+ar/S9HI17iQUHN9yvBn/y8pSg7+pH/NjNe6ybQVXx
0J0Vu37Y/zxAUdBK28BV7mVi7ngdzNs+OH7Cvb7Nfesqm3Z4iP33QwCPFfm+Qr0l
8eLV1Uqm33ADNojlDfdF/o3yWeLfhbeVWttPKDlNVDXHeH3TBMS/k+jlm7So6gGd
E7WbY9v40roVMvm6iYEFiUMIXEZBWut4fGJhoXScpZwgJLEGqlWtQ3fg93V18nht
ODnRIRrAtmWY47uWxj3W310XPzsizDrNhomguouca+Xl1byaPMUJCqrqJI6XESwz
cuDGsrGnZigUmm9O5iENhNb0GbY69fTTHDfFGec9XfTDuOBa/P56UpY+/dN3xMi/
L0ZJzNp334CZg5lx/4i0nC76jwHPF5aUGzYlgzjnCPHN9Pp6xWORsAXclm7F7NCP
d2/8THcg+Lm4tvnzvr+MnQ66PLVCv/u6QpOjqRUeuIyQ6AbKwDLxsCHqi9sBfeeP
fMkIXqGJaf7VTHOm2L4QsOiJphcfGbLwiv1SHjyMlvmFhc06hKQQai0SPf4SCAqc
Z55JT9suJJU5CWRr79zAYk6OP+BM3CD5295VKDcXWbMPz0MMXx8UuIc6AsjnSqdS
+nTX0uSFWGLlIbQddfCs0v9Kb308b0AMceELIA/Rr7JXBcTxLx3MEx7e8o/F6K3G
L5hXgk2Mr2EcqyaEe58PbgHwij5rHe42Y2Ba4JXObIFzoOnbVKu1tCDHZ5A58XM9
jCl2P+k98e32iXnXvQ1rOdl6pVxPvv1sLYZea76T6FrNxkQOuBjOzZ+5+vXnvERr
NQFkpGoqQlPbVhHUQzDRV1mGIGuimuNxDbk86fG84XzssJwm0Q14jPHah63mXW0/
kFkLJlDPgWkUzsNnaUbvQjCQ2O6bPshsQWDqJlU7wtxne9bLqeKue55k55T1VLUG
L55fHNHTiIlvElFfbdBzHA==
`protect END_PROTECTED
