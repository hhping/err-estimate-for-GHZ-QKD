`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1tI5cuG6co32nk12/R1/ntskZ+AZHr53v2bWjbPfdcFxmKQSzyaHQMmst198gTv
xnFASyOphoZQXBZ5PHP1BumgtyOfVHh0ZoXIS/hN8RuqLRiaGdbO6Ul+C3816x22
17iXR2UGUFJP3A2DEpd2AcHk8kAf6Dp+aWAe4Gkxo+Khw1OUPx/ap9lHufCxnyNZ
8nNkdWVkywlzt3VitZLBJcAE+152y2KGTXABB2criv52+4FJLHrBApqj/UgXjpt/
/6PZOAqRd5+8pmOhCE78dSXTRht/h31Gu2McbfXr3boqrZ91NDAq0s0WSZLPFCid
NJ9a3eZntmnPZDQVPpU75zasDrpi8DLbRMBqAV3jzVT8OF4R4aRA6fcF1mTHoDHW
miAF5hBduzDEw0RFcN+n6TGGBgO10kBFwuHsQUGd5mD1o4ypZKOV0OEx68ws9zkx
HP1luBS4ocuM1gR6COw8wnlJyk9T73qU18N5HIqbVYuDR9LLCA0T2aPHU5nFGK0A
kf4Es+lniDHIVhSvi6dKt2fqZHBpOWf9hRwW5oIzcr1Vie+2ozBGydzPdC6rxzNk
1PGRkMWofHEDDHiwluwxJWQNCMletvlNCZa6WSbDr4UEu20sm7Gb5aFxiSBZUhm8
ioewk0jndSxsyYLaA1prJ+gGYhKrhSB9ehBv6xEFrOuhA1Q72SPiOFsNEUYYMPcm
BHSgcCUM61BbXk0CTuW7PK7sWPX8UBQpLN9RN89iKSTUNFOexIGmmPwndNquYFYR
qoSKFrz9Sq9ftxGIvOLT4fFTY7s5EAYLNPRUy6jIsgx1TiXhCwG5JdnjT9Eja2Ts
+YEHvxk6j/Slp7WRvJC2ZwkfOS7RCZXCCIGfkdSs6wTeeltfml1a/qXmrigoyF4B
eDi3TuL6nfMPxUDBLq/sFlUZAn8gPMFryvHOedkXsM+XGr7RZzhhhnoCnGd8oCun
RQj9d42ptSaEu7DzHEc37Fm63S2Ghx3QnC9GTnJ49AhDIcxshwI657mkNrmKK6rh
3JWvELmDJWKgmMXerSzoDq0OHjVpn2yo5RX89MX531d55UWHHjLsnOePXdK55F/c
arHieiSe/qwetibDTc5hNj7e0PQsltkyErG+LVJ37rtrsAW53zjgMel4kvOVtZ7S
ag5bgbRurmLXxCJU/w74ETiGGenxWFelpUZYSvf1TDCwMUq4dzpxHTB1YwPfPvPp
fnLtDUWlpSKXpxZZmUx9hg==
`protect END_PROTECTED
