`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQ/rNh+UA2lxMmTSt/11V0lwM+3DNwvBOiD9SGKjQD+/ywOpti/memeENfoyk1I/
EOqXQYGC95mbuZk6uLAILpYyJrTCUeRFloMrVNULjuPrPHnbR5dRwsRcTwiMXKoj
rIfNPxRj5Q0EWciilh12jXuGqo3jq4DlATqKmrA77B6QMefbhQADWuTA0ZiIidGe
qBuPFqDf9yf0SInPOfo+8kL28ulDvWwabR6P33ykPzO5oap3RZuWtqqaXaI4SQ2H
QP+fx8HcYuf2ZlEIeIhqQRFCVlvy1HAO7OJhTEG7xXmvFUAMB4KcuMNdoGn9RKgP
oBlsHaVCfJmCYJtaRnD0xmoti5YV89mhGwzIfxlv3nzP5x9wTjy8pdrd1V7/dpic
2gia7IlgoEaL5BeDp/xfTw==
`protect END_PROTECTED
