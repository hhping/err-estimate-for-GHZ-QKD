`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GodLwS+6uLolQkfaHdfBCZV56uPaLKenov/CWCqpaEJO7iBKYe2j6nXw+6XdWi5j
A+kVxzmxcMn+UeR+bT5/jL/SvaBiWRWCEOpKgg6Cq/Xs0dwBHH47qH1rrJSTsWlW
tkfGZI3YswOeOAEHUmzOrb5xjFdtOX6pfD5i3ctHXd6KTjnY80UQ/wxCqFzKI8yq
6WGPNPhZl90Na2ZqoLN8J4Q5Z6i18QxLkDemr5l7degghgbmkdSsEGRSYXmUTKX/
GisTFi9/URy+zGG1CneMbHq65d7uFAgCR+t7mFNnC5XhVaFIpWEUJXVE5DUlD3CY
U19VdpueEVHaQQzJHbTBlOQn5Se/p2Ta6DmK1RRhEC7IgXgWXfYmUgaETNuAW+uH
q1502/s7Fcpqi61/LRvICZx4Yq9OBUcIsxAh6jbT9+GJw0NrqdTTQ5MpZL41P6VR
vn1jq817xVljZrLjyhaH5rmf/D4vMjrLJBqAGjVEcK/uZhH0kB0k0nlUlOgokKen
CI6VLJK1qA2IUujOtL3RO9psuBinK/fUd2lNIt3ze43rMezjzUTVNlM6eJ76eML5
U4tCRBCXgIhXhopvovUzzIdGdy5zp2Wg6oi3JqOXNmPzAGGUzuOPhsAz0k0P1VvH
JNet1eyY44dwQj4U7E8Q1aMzzF6tXwleqlj6HaK5KkVXkQMaUsCwYAn6/c+EilUp
WL8k03E38f0xetzT7wGDBU+7N+Qj4PL18SfkgTV4enydCoyxk7RlZMqVF3SVpszC
m+RIxuD42c4ErbuaZ/rFv8rADwfYQKM+VyvZY2QjSRPThZSCckl8c+2iLR70r8S9
C4brgEexkrDRkd5AWjc5brgcUn/8sAEw4q+fyI6TITkdhMBZGsBFKJAqDU7f4Xqp
1dwk5hRrU/UkbvGVJa0za2BXhhmFVJAwfJGvJfApEAmptbl8ZHZhzZdXtDv70noH
sd1HMlDQdulK5dBVg8qYFl/PclwbD3CzYoh7LF+DXCLpk0tVwxEjUlwmwClxVomO
7jMTSq1b1nOswM8OxF+N7QScN8WQwoCkh/7yE5zsXKJZTUEhgS+2XHdNSa0mDx/K
xRFLVmurHHyjgXUKGPjV5pEkBB0OQVQwuuk3fc0oDttcJJij1hkuctRs4yRoWipJ
RHoQDMTAZGdjVn5h1/CNf29xVLKEgsNl9njFub/E5pECS4nmnO3Q58C3Bax2Jx1u
MrgXA4CO2W0wNlzKP4CDikG3NGXrodhlmABv21cXlz/jvxPJdtAiaGPCtDjGRNao
fhLkEWCFN5QQwZe3Hrx7j6ZmdBOjl/GbbBEnYGQyiuFnKr5oHxS37JaEg4PKJ7Pa
D+wmJ25pFJizqTZVsy4hP1Z115yMkNHZ7XyOq7civlQqlObwCzMY+cce9fyYA23l
Y0ZXrlVWeNRFgg6n3YBBOHJs7vqAJBKQN6XmCH1agg62O4HwvDpxPtLy/qxcFS+S
ss9/7OZ4iFdD+weOu/RB75699JdrjNoz6FC48whFd5BpuhphLxLRZ6SqNz9S5fuB
BKvthsVFuZUvxbD5EF+Rd9NGQNy7KE17vMi6Dna1dV90nuSXBXjOsTCY8CcYCcop
WkV3bqlZDdVKvuzvKuLxQOlY3Oz9BY79IGCEWOovvInveZ88v5/4wKEC/tkUiGxj
BEjqAiGCHTn3iXK8ivTfOF6mRMIqvvPiXnS1hnb1s60uOJ7TehCysT37EklZKVc+
Hl9F+VZ1+/oG+MuaLStfpA/prUQ2k+vVgusdaQtv4Psl4ESLr36xHAmn4DBwoZF7
4VPsczqaZoo4Ee+IvmS5+z/sL0lo5B6d5dEDTqaBamOqCvIMa+IGzkbK8vxbMPwF
SmjnTV8FEUOJglF/DzAaLs8oSGGGMIKUTf3lw84iH5rJDjac/xkM4gx3hDng7N71
IxlJvA78aGTusHzmCYRRkmNmrYZe/DTFKvbVu7VPTLKp421YSrkVo4n6fcpGCY63
iolG7e6uqWbLBux2MLqRl44ST6Tb8gzxfSAV/ar9bz3lsgWJbIIIiRdaEMiFA/iX
NBXAYZRg9iivPSa+EOKxiQS14da2NYt10tdqK0QNBcXVEKcFMosCUPspdoEUauJR
FvV3bEGyccIxGXB3KZY6E8c6qtNSZ9vdup8bLTryvd2ZvbLZ3rLyWxXAwpniL8Wb
0OrdfuqaGF7QgSZAVByGCcIOdak9PtTM58+jQqrHa0Bi7dWDxKB4pVoLwc40hYNQ
eZxpNFNruGdR0HlsTAgQEXnL6LKQ071Av2g5wD4N8pttDh3Ys6l2TvtTJ/KOs6aD
KKKXD0suJGMj6dxg6tGcnrs4h5cRHWPks00B1/hMsZ3MMoTtNlO75ClQntWQtOwh
7ig62Yat3R40MBnZqiWejQqXguxxDc3z6XbMpayFQU9+ntCFXelT24SZVat7Iyro
9GxhzMueFl93Bs/BqYoRZzGgOEF7NX7d9K5BgCpbvagD2RjTghzutDUaS/Wu5AvZ
aycdxwKHs6159IvlrcRX0AdemP0y+is1ro6NjvspTu46K60aZIczWSetxHu6EJb7
O5SOIvlxySC+iEmZtoVXsMUPbI6fuwJqRTljtVtDxA6+Gfhg4THiL9h0GaV3HtK8
/dkqbCvxR8DsYjGzcTWdtiamQVKpilv5vawV92V62NuTx6kD5OVaqyiH31z1zivg
j0szK6EiGR6Q4vacxrB9tmKGhSQK9UcQN9d/8rZ6plgs0YoBtSxlGY8KOY/EDWX+
udjlaswCwf04IXLDcpMXNw46h5XJA9cpF5UEKHFm0SS2hK2uj2Kxk2ust2GZgQKB
L05Vzpttv5xxgdgRrC+getBMFI/8o+UOWKrSdY+Gzu+52DmuxrPwqPu9DzQEbGF9
zCNz4kOn+2VadmI6jb7fRRT074+CjYY+lc5ncepsDSXb7rJ7yA7Fm0RGVDau2yHT
D5uDTRbMvnKucx+Fu85LCCqddtmAoVDBMgwM+3dAJxU1YhIMw7uuC/Qx5/WmxwFA
gJFkIEJToDbtzjzeyrYhNUNJwSvaR7DTiT8QneFsUwEOSJWF4bgsHGqgsoLsrYJ3
nnzKHpuxltuO4FHgU6EakMfboMHg6NIBOsM+9wb/7VIu1GEloaeXeQF0rcKH1484
AX5pn/ANgNFaZw2FMavl8rwv1tqZmAuUPsKkoyacLFqEWjlWN2MTHlRpriz4n4bk
sTpecvQ9rg7qf6TuyeqmAiJdgUWvCmIMioLQo2hzkUmmnjDu4umHdVnwjqwNI28k
VEIkPG7FtGSAsEJOxFcpF3pS/QdSyQLEU8AxN2UwvNWBpi5ji56HMhqvfpbz6+7J
w4m4otZHaO3T2BUYecej6SobjdCJRdtQC+U/dyEoyh1YS3zVNgRIliYAP/Oaazj7
8+m1ZgMa0EvXcgAkprfsULPqe6/mz0nbjXrhF3gDWHqqfJ5/qN24yi8/54elfKE3
SI50mj0KURmZkkSu8Q/X5c2L5GWYfnXKGMjC3etilkhdsZEsEdKUyBgx7bp393AX
BRuIxyj54a96/ntvY+Ws5COxnBwSPNyTk8wrDG8sSR70aONdxOoSy1qpBq+fKyBP
eKKJfNHKn0HVlColQvXa7eQ8feZyQMqCdatgc9H8osNt7TdoFNMAL0ArqQLFd7Ow
JLCMTpSWhogP048K86bpkfwKLxxbVkreWF/V7g3int+YeAjn/hZ8yRJzaILsRnCN
ETbRSNvRaJV3kVgQ+qLQu6BdsWyAn6cezBY8dF+xRPFcYRWmP+5iEBCsJ33cEMER
mFQNsRmkdi3EjJZZkkfTrsOBEfoxZmjHcXJJzq7n0eDLl4RbQ5nAapqcLvcW7d+W
09ilUkFaAjd7qZnMv2dZLI4PIxrW0O/ZhNNLIt6sS/VSmpzDxtsjZHetRgRldqV/
AQgiCS7hAcVqGNtFD0ywDRIwOjNsio6UoIgoGNhbnRdPJE/eCHN1rqlqCB7qBOk0
pbrP3oujh8TdkZqycf3rCsA1bc9qnrw1fa4P8ikwgWjfCdFxtmr7JEqqOaZMNyaH
dTCwfwDb+urR6thHWvzlF0Z0XeSH1RKk3yp5qONp6HqMuCtBmBsH6Q9NFHvVLhKr
/zDo/16+M5v0RrGuSB6jaI8iU6XlHeGC4cr/VRWozD6bn6kNhKu2eH3MMXEjPpfa
awLi6wg1fL9ZC3LIr5tF8dN0uSmmp1oE1F6F6D5Z+2fTD+byWM+0KbbH+yURyv1U
E6IZKTQ8+D10duHHqBzZNGtju0Q4eOvSej8llTS7ua+0xizwAwDx5DMbKd40z9tm
IAnEX2wi8284tOWcWHDgsbo601hzANsFHrq3O0RzTc8yPwJd0aVM356Wf1q3LS7r
zgGnsFjKE4FIdsBFCy8/DbGNfRi1xKDh+SgjytOcv7l792KVz8Ki/pK13qkcOD2o
BtyEx6IO6Fw02QhJC+ywNDanjMzzxX4wmgTVGtXPGLZnBgUE6pFT3anD8LDO3Eyq
1N6uJcIcJrDK7vc/Wuc16fZ531kpZHHH74IL94F9A8F/JcTjNtZpbMeMfsbLa/5+
oX3y3pSIroHnI3s1c2WL3/zArnM+UiPtgaoGveOmeQiXQmV3SOGkUyUSsSsk7/8Q
yoIWA45SFsyBeMFEnrznFcZ8ypH9E4QkFOxa9NItlXE+YTI4/tDOK/pCo0yp3HNr
7TWSpRh/LljPWg5nwm7wkmDs7lKLI1Cf31s4X5DFK+Ql9f5BYkYM6XlC/FUlTfNd
HdUIqPa5bHDfuUrTdTmUMfYxxkmA/Tf590/FlU4UYc1tOjFTvAv+ynwEpi5Ri90Z
Yisvh2sC+aCDlIiHtWyJYEZlaulHsfNZfAiarpIw6Iuo5FYB47EGsCq5Pvj4irsu
Yj/BlH+x9ckYZZwUqqXTB8Ypb0foUZiPxBf7QJFjOdsczsPTy7BFIyE2DCK+Nez3
o5nEjvD3L95pHrTmRBVfTUlmYaFr+2vxx3iaoVzP3uDem4Q4QwbxIQnd5TZg0kLu
2pF3XrKalpDciIbaEZUKKW+B8bwyKNMhWl6lc1tGIPKz8PBexNUB/LWWoM16TruL
W7YGDHFQ/Cu5ds4rEMw5WUigKbfYUF6fBWozPhU0qDsDEehCwvVx11pUB3MIyFYR
hZt4M887urnh6mK4QDHuLr44UAxu75z5861Zmn6dWqYPalHjQEafX8KJ68n6z7JQ
AaEvvv+SxG8ZmiPVbFqWxaGDcIJYO68L60zmEcXs3E34stPUMqsLbmlhkrzdXC8i
OqlNj9kIJt+nxWrwVU1WFK/E00HdiSFVXSxVJUrHo5y95P/esuGsJrn7wK6N4FOW
99DM82oObV6BwVYX2yCtHLdJiMt1COxl2yE6Y4+YWkH7Lgs5FmEKp+AYfcJaIQIG
iEqAFa2pjqMToS6FCQ6sVsaCu4tafx5GGZTxBN9qrKSbpFBN1Y46mxUsD0awIGyz
lUm22yDX64IlW//Q/uiaoZS6K5tAJ9ndkYEE8pm0Au2oXYD36krWxk6ZHyQPMqA5
XxQcZLp++fTd8dJ4BaLH9Di6cbke7/sbWPooB+lH2eJmz7rrFFvm0eLilGlYKa0o
gGxZTPGcEItSoyxbzUpanjjdcJpW1kwpx7IIodIPyVq7a82QffysHjYKmyKJOFDI
Z8iiN31UXvmxBReBlLxvpM9MpUhEYxUicEO9vQZEhsAIW3sT+gSTkQAUuqXLSob2
7wg+fu9Q6WlZ9dk2nnD+fnsAUPqau1Jip3X4G/W0aTTQkmGPubcqTrRuwMnjYJkc
ypxs6JfFhn8OwyrxGYC+PZPb63bAXkjMhVJ6kvTF+Ir4kPYxxY2Pp+d0pYIg9NJc
zEN5kn9yHBeecU+C5NekaCZTsYA+2UUNJJMEkTvZmPnLTDNPTv3w1GnfuvQgbPhw
uTAK2M4pztXDpR3K2DOSElkng1M/V/2W66kCBFu7bTepT0ZGRk0nDwrt5brJKKRv
dgbkZiFH8yoB3kpWoWao+MLnFk8ZGlpQ86dHeeAPfdFBmvF4XjoFqoEE3Fm2mhdq
ceelmPjS7o8eLLlDnhjm8hz5nYthRQrlCQiZfPC8OqsgzgzgHCWQgmeb6sSQs7b/
ay7qpET8oZLTA/aZaRbqEGOPeIzKlTnmPoDXbqDKhA/Jz3rKHZueBbG84AfujqOw
B+pertkwFHf9Xx7GbE0ikuraTv5c/7E/J4ww8U2vz8HYieDEcF2q/hpzYIkvs8QJ
iqsHM8grrqpqpG2r1Tp1ycxtzkKc7bd8BAGmeVGQu9HPPN6ysQTqOcyMSGg4dbX6
C+YdtLEJUPUmk+W/ViY9lHFF4n5OmYKh8rQzWAYE70sMbaXxePjlz1K/FdsuexuW
jw9R7ULsJSKsTzP4d+PuyF6Hjef/3nyicVulOIsJbAaHiaL6aqmOY+RiiBbpjFpu
zu5UKUKd1f8s7AiwmLDIxrplj4+A9RPQBxYapR8qID6XvKhvXoymoHiOwYcbWMO0
zMo/4HZg+wMNGTUHcYVJ1o/64QJ+6f7ntJQkDcIJzce7dCzacH0Acklz8jCoGc58
UTeEhse9CWm4MOrzZTzJVaiWc7aRl4p4wKLwlT/RTaV+h6e81jVr3pFO1v5odYBB
pYbv2W5f5ijkieigTjngCI4ctfXWOJWDy2EDLyxnPeO81dCd6/Wv9rfxHDcBxxMB
UCC+sejUThgHbM3ZnZ6F0umnLMizbwDRi21/gffZ7TQCOx8ERK1GuRt/HILVmwF/
72sft5Dpsoc5SD0yQPIrXT+/Y6hpm3KEll8I+Okhr0jBOMIfj/m69FiyR9xxcC+c
EUGKElyxf2OvZNSdawINHnATZfz0d+a6+lK/Lu86+nREqlGNB1bLlzjU2HxgYyd2
rCjVzek2ps3LPM68VAtVl24KeIMDRyVLgrhNRRWXAaQFVzOnqQx2ZZMz9w/xf9Hp
g05EVOhhMxMRZKqYfTTBQ/PZXR1SN1T5OE/ostgSRpUhTMn6jlF8Sq3n22sYzHFs
3NnEbfuucKrg4NoDKTaoSx7CRmL5HjpHoMB7WCOsnDs50FVV0v65F2F57sQ+VsOT
RZZVnNnVMU4vD1UHH4iqdU9OcSjA1z0FJinFH2BjhhkGsIciRAxPyYMw0uWrzhK6
1jjDHIiMo8flW8rnRvQSnoeDDWmB7z5gLdBGmmMUNyk+ydiTsya8XoricJ+WII9S
ZVueExGBiarSiTqx1OpvdH2scyX8BqGPtGMK43Y9LnhHpTgY4dUatgEgRcu74O/f
WkuChqFGyW59XQeAWzADzAyC8KzsELttGSqtH3n58QP8VsX0BQdPJuJ7nAujPb9b
reNSPaWqjd5XNKdP5MvS7Tf9GYGrPPFJRAvPJISleDghO57dFtM0az/6kwLLQokO
9n0Jnf+Nv1WWDSGVl8hQhttmHvtLYLZpd2Y9yYikLQCKew0XgtLxi9KHIwTpBnnB
jERNO1Ut04g6dXUK3VqVIK5ZDKgb6xQgsR+PakhuovpeOAwtDJeSnIxj09a45o5n
DVFgNN5eL81ypwn0KwxOa9oLsTNdjyYAy9GJMjnIxJZ7QhqirlQv4x2v1jZb3yqZ
539qoEXE5yIsk9yY3OeEMN5qEwcEmiGWkEcNAMLLp1CX4psDEn4/UXqUJOrXQe0C
FOVCKCU0Tf0KJWT9WZU6Q1RwaMKDBcmNzkyL1St5P5G7+yQWUptnhbDu7Gk+Ocms
YZ85q4ky2KDIp3+ZG7hyuhcJ8qUDnrMryLtIsxKU384S0Sh4ZFAF4RUo1Ct1Yd35
8JB9i+FNXx1ENHXXIRPoV/gvElG/X+yAIxlm8J6ffjfMPGCM/lbm5BgD9UlEp2sm
C9R92f4Af+tFREgcUjnWwltBSZk/mFiP1eH7zTZyQ3gxmXbzZreg8vBfFhsKJlFQ
Gafd+GW6rhnmUQt3QtSgxijXbGEiu6lHM53CqqneNXckCywZ1kcnlos2WdWi9DW5
JMXIZsU2tamgarkoLAb8iWB5eBFxDiKfeQKk7zmB/vUOSKR3303RxRK7YN2DxRLZ
ZuaHDa7987c5KAj+9SFhHoGHJcOyExi+wahxqZjXAeOSh+vALb7B/Fcm9vyC4mtU
qoh+9CYHLhGq04aoslKUiajdQ9Kgwqvwp4TfScxCrs5n4cEScL6tsDxlkFiV35ji
BFwrH45vCEKhE/7kCoTgG9OASzc3bb6UmnYusDzPKejIOyxqRB/uDgx3sc8hCS3V
M0e8xJW+ZeFr67sNifo4cafBWS7RqUmRVJ3HMVNMqJ2rpq4FEbrB4Zt7LMsZWmsI
sedOtflxD2/fP9ayJ9h/z6EE/XOP1w9Wx2FkpnJI8L0xsQ0MDmHq2S2QuQQP2Kn3
//9ucmzFfVIDorBOdG2UxWLPxWMmdgxLPya5OU7CjDxbQ/HGFQ+2w+PdRJlH6TQV
3BaeT22qm34O6QJiEZQ50hhQqOM/4bxeWnt/ivi9BMWTIEEjFbYERw+GZoFsz9YM
bXsXbiADXoi6ap5iDMXes8t0MSpDRx03pnfDvgye1Lp39UWvWoSnlaYtf6n82TdG
mj4n3TL8qLWaR55jlpMNplYz7iJ0ZZJnYWsrp5k6rGM6oCmBK5eiGVvfiJh9AKjZ
bKbsCPraMIHudq68R9rKTG9oNAcnyneU+8t3VOnyfX2Ez3YmsoyQiDFLN7ak7s4h
jf4GpgQbPJTCcUjiRrc/TeM00BqlWDllcfp93F5MPdxWJDIHE7pak02ng8iTMBPa
1J0OG5NaXcE7MbIQpjrWx6HCjXuMeJDvB5d0Xh1g8NPVNF04vl7iKqe1aJ5FrKmg
x7WvgbqvDAFAHY3HcpeE+VtIHJI0hYZZ9wMYl8F2ir4q5ma2eLOq2A61WsUVpP6I
/7b7mO5D9d0iR92LowLWydmc2FE/DMkAzuB12V3VgxTH/QigwE6Z1n/QA786KoMV
CWPtwAOKAWQWY0gz2Rt2DtfPZp7UUduPJ3iZMf8oZvKI/yAubaJ43ffhNDfLkYEG
eUEPZtHTPIJit3km2Ky7P0/7BZsZl5wHf6zVUF6B6mIApsxpKJcqJsZt3rJvzoF1
aAqH2viXpvzB81wPxlk9sLlbK5D8sGG9ATyRCoIynqu6HI7gvGIcLle6FHPBVMq2
ejamTsCrV3DUvK0Xznsy/MYSUsBqAFSm8Zhz+jjdZ5x7EdLHyhYE+go/gBcMDEN7
1Ahldp3Dprx5zd+0FiRFHGWhpc3XpB0Sy+xzmv0VdL8Wzt+Pk5n0X9VyEa+eQnGt
S65DEnLQDnhRM+sgluqL1mc6c1ifGBf/46ssLUSpTI5aRzHNh2K8PIKkgcP9qSGO
GGZq55tEe7jRKIeFq5DHieWOhAmVUzqHXUmdu3la0dxg3SOotwFR/uZX3PPlD9Pe
56xNthGpuGVFxcQyQP7WDJOahC8nU6E4a2K1HTu6J2IIqfX/2EXn7FwjHZiL+a7b
Pt7CzSSwiQEdxQmXs5wB42JoSa8xA0w3durzrFbBOqIyEVRfzwZQQVryiAQVOgLk
kPZ4s54KJdzoTaEw16jGRzLoEf6/mUgwyDODphXFnOFJZXLEqbHzS+eb2p6qNn/A
MHzzAlCwzNkm807OzyAG0eA015CI/ATKI9J3nmQCThpJp3hqcnHhDzxXljbiFaQe
esFAnxTzgGvxp73M1M9wkXSHqughKFCDv6TXXU/rROynh4JrPcW6dOQen8g8ZdcO
/NIIvLyMroxzBgpMJV+F0hlcRjdrnr6QH8PFgJQJpwofDV8apOe/zt4oFke/0cif
YHoPzF9/wLUrMSvF9nh1eHghO0Sf+03FxJIde4KEq4dC1oIHK5uZ49uYzg/GaA6x
uMeWpgFCybCzcaPfumBq+sdtt+QDicRF3xZurm33Mb6jdI9FC3jdgUyUoQPcVEcU
lpN26MvRCaqvc54M36EFKNxYtTyokzOyLAA5JgeA8SyOT0dBo69gwqeugPRwqvtc
dGx05IUyzKXj6KWTY/27f49KOUgeybSlqtOspOumN5GlW04kT3x8E+e6ngbT9qbE
+fwtjHyT8p203MJhkBYxtLriunZ/6MNeA+teG92+ijw5lmWfora+KW053iFfUTZ0
DmT8YmhsTVE3OX/tfrZHiJ9aMP4EoW6JMUgnuEQ20m7YgJ3qRjQ/t9+ubMfNsUsP
0Ii+8yNjzhq0e+FazM57Cp/8AWn0s71lr8JdvSDXRmNCjK5PgbhhMEQWQfJ8Hs38
SuyxwArtyuzkrRRYIKunat7tiFzxtA395NujOOcTnTWYscU44rJ8O1aiFH0gDL7W
bwLobDRNHu65+JjJp1fyJwP6uKm4FIhELt+/3LWdfdB6VdSp6NVs2SmS5aciI351
Z25m2IpQQLmzSo+j+B2uloq9SeBb4F6kCQscmRyLfk0lQ1eY6OBIA6+mqMzJkE7S
ayl/VNTVZhkRKx/Z7EEfzATGizVEt1m5GbxXe7YVwLZ1U30a2htvSvVWIRKJ9kyK
qc1Pj4Wt3cp81ku6oJiqAaiE8KJtmEB588K3PMek89Dc0utVOfEJNKzkWqY2POKc
a88zfYbnxT/06t4vbCAbuPlbLxNPG4VYxWGziPdJHHyDh8nVqouCq/ebA0mcs/bC
9YSmHAnqsfwBNOHvwKDMQX/+2fZiMn0ZvIlUNdYdnSZqw7MPo/nAdg8Oj2oM7fKr
b1yyuB2mo4X/lZPIgXcBrjUIzJ/U66qeCROeOzIbSr448EJHPkQ4okl1r2VhjyVJ
cx1SPlSe1v3EZ3X4KigrIO1lhpyu3EuwGa7nKq6KviyP2Roz/vIlhcgv8dGUYOLb
206AI7Nqjv2y839UOqLHsnOut5ivyXZPJ2RErmkwHXq8nclpTmGz1Yp3iOuXZeC/
gtsUjrSwSRDLXO/ARrnrVNd+yx2I7BeY69k3UlcHJguAUTvxNvtSDRF1fIdyoliV
VMRWbCoSQF8Jcoe4FvchjIocZ+Nwlh5n11tGqNhe53LRvKjebPDfjZF0CzMg0IR6
2bhlOcBcDWk2p2bbTbYleyEIk/7wSbdHlr+quPfFcYhtI76HO96Otwedfss7LvDw
xG4uh8NPyz/vZ13dzWOGT2sKP4E6kWOg0iqhVyteV63dM3gXTcfEFD5M7HUUiL4D
NKFKkepOMgZJFSmzbHXX7iYLhS0/RxQdVRFOT0lLTEa6NDaUl1Nh2BaU9hMaa43Y
dBEhEhta05hJxV7XIpp4oQN0YDHJk/rsS39CPjHJD4Js/5EqIawv0TC55nZFwtUG
bBL2M7ANIXAxqq/FNGfWSN8TmX4IHaRi8EMfLZx9YMt9VAdyGdeyq+ufgdEfc2Ap
1qRookUo3atJtDIsj4A3/AQaJ7A90DNqEmuyVRTXBw9rnGOLWLv23SC5IRw6cbMh
BDixoUi23befzFg3oiojyUBZyU4uo5pw0EtdNby6GuqjypeuGHhs0w0qAjDIzKfF
kgqufjA9bwidevG5TFi1VkJOn/mvnGogQKdz3a0j6PBjI5Num2NaiuDsoEAFvVbV
99ufuBgc4/3iDct7VdH3hIMxWkH7DrbcBZRonwzXwkzA5Ugk/GPnhpz2QN/SPhIY
py5lD7WbXpn1wyz6CK9t4l7VCS4dBwySoOdscVNrUUbCJlSvD+UgdZEoskIQTSbE
gPMHGJpQLtKvrVKCmlWL7xiKdw01ZFcFsng/mN9nNW2M3GMRPFv7Ffd0PRpoz5dt
sDbqlAeeJb+EcRIjXHBI4jUFnoNiBCZaDKNM+eLUHud0MVt0zqLcRAKVIdf58N92
xhD6VjMLbG1K0AtpenUwtxAAUNoAT4L8TqA59FRLuXZrG26SWIblDdtf2Dj/0cV2
adZXOgUKRcwYrdmR5tXM5ul4ujUjfWcEuwhWB6NMasNw7VXLIyR3OspWRl5B14eK
171nk7Ny8TMdi89Qo0cYcPkgIYPDAbYpSDXAtFRWFmrENV9qYhdgHcHBeGmxMWlK
HGuu60+8c4DhNFPMMH5ro5gPISQlsvdvTHyHQaU78tOsNLvjmhmk77FxV4elFpcb
PZPC3xjmwS71ClFxwiZjFfgGn7B0km3koPmCJbpqfteKlY2GYCexD93oDYx+jIs3
ZtEG8TWva8jLMSYfw2ayCdfnED/m5goJTTgdVig2ydbEJ7VeS//l18jYXmw39OM7
jgT6HgEnPsImaUD90YJOhod7depLIPQz3zkh618r6UGEqR6O4g2SucdwZkSY9so4
GZA/QL5sjNBSy334pRMCK/Y1MMponm43y2FDu61Czmlyup674Na+KanXUDp6tV0U
wM5OB04ZOwWGHPqlmW6/SC46NHM3+dgI/yPHB7Ol+RFzbd9aMGwAjL+pneUDtn8N
FtqT31CPSj7IhAMlQFEYRbx89RO2emIKkXivsUim7gztuPi/4qXkQNM8ccAk+jDV
TzMIEKA54Wc1GIIJS9DLSFeVZpXT6x6XIlf95p1BMqDHs0a8j0z67a4YqONXGNfv
B4E7IHPSGklMtOwadfc6CVKJrBpWlnMfnN+f/9Rg1oDRfpJ/zz5FjiDFXBRyJRzX
vXrnULj9nGmLrdlZxujkguNafs69VKQhlPSaeDdmoiUfYZgXg/isF0uqAnB9Droe
pRxZ7yrQ2MG9wGt2rhY216VWymhP8lSIiUQAAGJ0Ytx3X7oUdtUD3ZDghn3S3pe1
a9tWCZuPIhG1CED7TNpwKFgUEnRZUgZW/PqGqLxy/+E7705AVzRltN2/29t10FwJ
PPJT4etuL4Co3qshywKNQPRuCF4OxyZ1yihs3OCP+TpP3mtnWRm7AwF6Pp/VBDk8
iH46aMRHVLaTCixYLSKRjYv8DCgV74Mobzi6X/9Vc7TEnnKoswYgTjuMhD5TI7pe
jLgr1mu2pQAigzCUvouNjRoN9oPbz6OTar1tTR08Esr49A/7C8EOQeVcxa3Uq/4A
fK9YS0G+rRH9lb9ETWKp+QXSAh8dsrIHF4CcpDnpalXtaMyeGEKxcr7juyF/yqOo
FxDXVxUDGOs0195bbNcJBQovkAtk7u7e2XJK6xjfBKs2iw8A7lidD17GrDG/SY/i
gpFvRyIBN1QH+MmnZGd/pJ8ztzJXPJtUYRKb0bBC5craZzX8+YpkuzDq+/GxRCHS
eSQtyj+0g5wF24TxjTBQeANJSAbFDUiXstasVwm2f7/LshUtagH4xookP8zhm/gD
CUuNu30iP5yoSgtZuDd5tc2VHo61OTGDsPDzCBvGXdG08WJ23cPhRVUlAthCSTQs
hsv6MgkR/VGMzL2UaoA2KHyMuMYlMj+tP5DVPIxE4ynHKh3PXWRNux4BQuWHUROk
aRBQqsPTGGOrgcuGmg0jJdnucXbKfQz0OcomkCpOCiKX2P/t4qWedu2/WdGzDNyG
RKvkRQBfhwOM+xrnzZEeGasfJdhUF7deweN8NWJMedkdWqMWnCK31LxGg0EXjBug
d2z3zdkF/WePqOLNFg90zO2zJdKjgpxz+NTNZ6NLJuuCAtjJknj7pERogdxvY98C
96wLDaKz+uzsWYmDx0OIqtRehDwMRIEKQSPfiwucmm7B+9RQvEYlBCtZUZdHK4iN
LGGqT/De56QHdovXg8d0XH3FdAw8QUBBESLsZ/CHsAHMLcx/pe0WKfI/mMGRv5ed
9VApMGghQVOxbORmteZtAvyqy9nLxHBJfWakbRvgKK2siKFRbbeFuKNY4LXqGgCO
bDDM9TnoVdgD5HIo513BY5abpJMn5DzN3spSL75YqMKqL+wHVKM6wkqRg5vHR7zf
P1CykbHdOeFoGjqO2CO4Chg6WsT5Nv/FsLxjJfI6w6VCpWlT5+7o/XKVlKnVXrTH
2nehQd9NDJdC1nfukV1XJUcFCS266srCBYjkHfRS6FCJlv6JzkYpzKbgiq6hHMMp
NUFZBeGeeTBdD6D6rUuF5Ex06Wd8AnUhau4o4n8SR6YOsSIBGxRGrGh9IfYiN3LI
VrL/XtRSvmrBwJAB1sHd27zlXhkLVG07PFdh7T2KAjZbrC+EP6ikHNB1RQNrJB0e
rmsObcEPravFx2B2cOadNJVFD/xzusIG8IKVOiXn+PZoLd0CO7sgYVYTGbBeeoL5
GQA7gR7cHCdWff4z5l/cRpxAdHY4zGf3cVrr7EyqgY1wf3f2/WjUDhqfkJiBJ8aB
/d99xBx6wCPTwfL4aa4IGpM3kN2lj8Q+UDEXc4zP+Cym5yNPNtDXzhOZaPLrhH3o
cmAqEmpqjKZx4L3w2DnfkH6OVKHqXArFON7ZZSZAlAr4lI+5t3k+FIj4J7Fp2nHG
N7olFQ4MAep9wC0Sis496MFSwAnNxEWOpJwChHgSxowxVIt+L3Yei/grdj+oY7Zg
Arx38oy8RHDxhYQ1R6zwGcgqH4OprG5QA60zABxmaG6ax/u3IbDs4jrU86zRS2n9
9RfiK2Jcyo0Jb7MQ2jjIreLFo7zUCGfdxMY3er8CJeJj+xpYnWTTOfKCDKEV60+1
0mrl6n1YXKbG2BG5XAnF58Ts2ZoT0Hn5oTaCA5VMmYhMpMIt38USPM4oH0McKCxo
ttz/vXorFfQGTiFmVzwNPYTvtx+0qDDP4UveQovLWxGRxgQHDPESCVeB/WNsJ1sH
7s/J2qKUEZRmu2Hrt0/VgONlUv69CoaxTIKXFVJZOvqNNfGbWPco/SqxeTHCSvWx
tDzfSFUf/K7WjGSznKt8o0hnvL+l8jgC9WevEuqntcM6t8aUvxfjuiCdSAXaAPib
NkAWCi9SasMOQeONImFruHq9k8/91XyundW51i3ZEPow4BXXJTF2oGzz+X2WHFa8
j4r0pQQ/sjWYx3w0DdG8XMR09nZZqsigOuVr6B0zZaeIGroBZeZQ5s3diAM4N1FB
k6jUqVqWRUdRMGW3nWAbBRKxBiaoDRzyAtq8EWuZAaSx1HXBYTxoknqRpz+qhy5s
rsaXIRlnf80+yX8uKbt6Mmh/tBsiISY/ti6cT2kKN1jgRvMZkvHdT+Dwq1uHvlG8
Gx9so5xZHPqEhQPmpvRxsAPeM5+THfS40Br5abbPSyOwebl/u3b5XhXD/mDYGGpH
UGkVm6UbTt6fYzNUdTamP0Tv1phUDLBrtO7e3yqGUVGGVGzW4LXrjGdomimVXKF5
73/pZQ/i0E7t+Y9OZYI7AuQ1ZQ4tKy6ephr3HYMvdhtJaBiPfSHYq9nsxB3yPkgm
F85uGMPZEBiKcB9ldTrmK8u94prsbvG/Smf9dvgoeSfZTpdwQIqi82HDjkaDLucQ
OkQQ0+vlq4xS1G0pJnGvuAzJ2r/iNaDKeBuNT5/HHFyYUFSDfaaUQIZc7i/k8Gzb
tqiJd9YqF39D8u3jKLPBKbXpT/hUoFZznAIPmmzNa1q1zgub7hIstlxwk5l9Glt0
7j7lulCofPSyMWaDspmhSL0LCHV0Mmm4XYc7NBW89dpajBfPjKvJ7S8NWw2DkcS4
59hZUAxMTb2GuI/ZGHo/IBSUBC33gIu3M2+z5+YW9+42+qb976cUV8pRVl5dY7qM
rCRLmhkQFwNxDGrja/FNb/oYUMYTqPuUBwgZ00E6h/FJXotwhqGW8SUowOKD+2M6
lTmW0ufVK2PkGO3oLQjPirG4lG5Jl74BJo9A3lnVyYr9saO1YEAAUbndn3NPTw78
BANU3FUWEmtwfXtbTh5XqY3iDP5t4i4b87dawlx2iIHVDZu364k7E2WGpOh4YDEq
cI0/KKLQBkeGyzDJQCbaVXVHiuaQEVNhnuIaG/yCeooyp0ZR+6o8ZL2Td5UZNhQs
ZGYITsaHbt/aS90zPoo89ThZ9PyqhCZ8JKW7ufktc9e5u0pIb4qyAMtVTEeV7iiY
MPpizGymDZVanJVggK0zFd/DlU7n85uFA2ecUrjFiwy7TrALgKhAV82mUnFLO1Aq
1KM5tssKVlEONc0CPai1pv9yVk7iERXmTf1ulngy4ydYLpapRdsvV8PO3Ium9N0z
UsllPl+IkA4OONjJESF95gWVhpAEVyKzz8Ru+NV26z7UXVjQyzXU0jH1EJk5106K
ntY+PtfEnndlJf1dYmCW128WhqcK2wJCaPFMOgVKu3//V97ypDc5vuDYP7LEa2Ao
owHajjpeD5ikHqmogS3fRVLCw0HoWG9bSanNUcziI5u6IErH9n+TUfPD6Ldfx36K
9mbyF4Ec/OkNrcdxBzfZKPNyIV813uNBUd3ACtEsZ7/nVlxKse2hvNugkXTAMKaN
dgPvk9CMrqYok3DN91l36OMS1DnaTS/7WKw1SWwLZKNVgE3Q2S/pOy0RNW99bYLf
ICSMVb0Tn2nDFgqYA7lT7V/LMCAlOOuw6l/yqbOpixz0vYRVzsdkHsfCLt+abXNf
jk15jLu/bhYT6+TPNG2P7eIdqowoO06s+LlmZPuFyG1l9vwbHOTlC2kGThROhvZZ
CRoBSrXObxFtevDsR/M2NW+7oGxBUw0zxczpCq+ZXlNco560RTYTqNW/aca5sdAB
Ta/fR0YkYhNJW3GbML7dqRt2LSa1uNFbrKnX9nEF5zNmVY1rCU4aWqX1FNNQtaJ8
Kd4wmdFhqza39g9PoNRK0/71Kf1V1nmFz3Jp+wAQEHVpFs35xNVXyk0mwJNsX0Mp
JhjKYJUw5eXIqmJEtpQZ1eF7uIcD7jgCfuMMMs9+Rn+48Y/DQPiD/tSqOCuVOlOM
Z5bV2XUYCI+BSXqAGQh/Crtlh1+xgfCxxM30zYnVWV6xx4bgz4DUp4qAsR8VYMvJ
5mRLvTcbAk0OqxtUEp2kOQvkiuJfggqcbSWxBR3rCcJswxBTGGpXyhQd3tKOrn75
bGRpXhZj0+eVGKMQBGjVIeXsDWovL+THBoJRHFJB+mJUf+ojkawycEOyBuXOCLa6
r41dWAG4N9CuCKFO6Lsd3j+O5XOdwa9nJ09Z3GA6rAeLJl8T6NkQ7EenftHlq0pC
DAxHJ0jSS95CVoenfY5jPGUdtKIYrHeVFUGt2Z1zNN2IXUrtNJ0tg79gbbhqyIVZ
z2jS63LeLTn0rruy96PMEfPf3HsYrDd+sG4Thxo1m/ta9gbdFfTA9bQ3YIGGgBrB
wABvunCTzLsDDQ9K/PO5CVQcjwiER7DxUo5alQWKBx2/bR69KFHD7VzmczrFfd12
8j9fZ8r7t4hlF3t2QnsoqEdHC35tzwlmkEqQOxWecSn8QnQjOyJw+A4xjzWngXQC
mCwLEgDJMYzoyW73kPfy1wLB4Y2S4bxZwjfWLPXdEM6quI8ZsWPW+5/gl+KAIuIn
R7qgNpb53Y8e8aNlMkXgY/XLLrcQ+o838sTjL/Y6GY0bVCwKS5n9KGzZ5QmgEL88
MnfsOFSUHiZHypi/MjYexD0z72oG6+NR0ebHeNLcPInnA8KmN7r73a66ewXn2m7R
Jo/YcAOTJe7enASj49wBTULIEdjEP9fpAENx/Lll3fhnWEfFl+cwhXO1l5bwIqkc
/4K77/tnjPxKA4BO20U59st0Q0jRKYAYTIk65UL+AaRqaNa8vp4d2DPOapqJXnMc
xIgu9hEdIKNJJ6t2vi+f7GWMZQkmbIu6EFQMXMj7UBOkMd/3anlyidexau+nBfj+
z/c1sboIm8NJpczlpz8lUk1zi3Gj1OT9xIg5IXPoiRfGd9KU62NMO783pD+oICnZ
tk9uFxyEilQ07M9tj/JImvy3Pn0oSdD5hMQ86R5ZZxVJtE1spReWhz8X3cs1aMKk
NhSjv10EjPYF8ArXyf03OUHqGt9qpDOqIwuYerCViKHphFh8LY0NSychFQ6r5vwC
y9lV2oF+9W3PGIed9k+B4+CuOxPLO6rRRdHFFSDujto4Qq7r9iEbruFBvzG9pM+K
En7QybXqJjdTC6RMwbGNeVlqQL/rgvemBLBLiEpqQT0lgvhLYfE70q9UMek/1Ms5
R0fBMK3c6YTDdyh2UnZchA/cKBaFjPJS6kq5ZPXAGi9G7gw56NRIXvDWSV8+S4SQ
pInOl5LUh9NLd43z9v4BzkmnvlOH05va7S9xPStEN+7376+BL/gQLHvjUQ1siLYj
RUSLfF9WNkhddX75kE4V97Nazt5v14z1reAmSDwO6/p3CV+Tnmm0emzVJ+4en5HU
SIN5wa3P2oA5OPuS/RKYofC7qO6WCYLNUunUmZRLmcKMo+wmir8xYEGUTsfrJqi6
EfUitAJz0Hq6lXcWeiur+KDoUcfDgw+IQMr92NsGkEmIFVWpSLttONp0Cp3dP/sb
P7/HJJPaw800iBA5uquo+e9ouwms2EuqllOFc56wMpeBdmTu3lEDXrA2np7GyO43
ZTGvWlkQ5KzWbTZ3lqKO/Q5ZfHO+f+FDm+Gqvt/sihMS2w/LNyVUcRsiAd7iN5qJ
yovYj4taRd+rAt/U+PdjEaPtWE1oUlBfRi50YUs/0U7k5F+vCU2QnT4VZGeaELEu
cfgaU55ji4rVVaVReCMIeyz622T8mfrob+DdyjgKhz9xLBkXzwzHEbYOaGYL1mqL
YDEBi0gjXtLlJgQ9xF3bjveEH3jIE9kfdzWwaKn0R5VmB3AYvM6PvE5ONK0uSvYg
3oT6g0DVt5p39lNJNg8SEmD9yJpS9q8G2C201gRo/qM6wk+/wK7obwg51nTXL93M
oruYeJO+EEp4s4LmoVlXqjyLmcn3hFqH6uDcOu9Ye/b7SFnUt3iJt6nVryvmGxq8
UtZ52moOlGB9CHQCwHh+TD63j4zoCfjjlUAmhD0LofBZA6lccxkYa4yFonsoP3Lz
lK6kyDqcO5VThgHID8WnSDvV0mQQgslkabgXR0kpoa+4gWu3/y1/DfrSVJQrELa9
sfb4PxXa4vsPPhfjmqq3j612KcI10StaaJTNxEKHPH1vuajWgrpoufsrvOYK2zb/
+fgJcHVApOMCa2wyTXyzfFjrAsgTVG7CikFcpdPFb28qw+2P1giMY+Wa1qGrxKVW
VgSTIKY9iZq4xfiQ2LDkkSJphvpONNbJ/hBgWC1o7xnczKtzK5yuSnCI/b07wfa9
dR/bs/+oQlFoSLANDX/TtLoaaFqah6sp4cXfKAX5zM54fiIz7YFGfPEBVnEj6dne
pdcs1XLOsONZmnEoHOsQjTPUQhmeTadLm7oMrSfpc7s59ty5J72tdtSJRLkI3ye8
SGP+ORi3ySIPvUUon9v0hJjFT3Jn5BXAq2NvpxGKk3+i1qrqYwPiHAWiovsVSvUl
PX8RvxwI9TSoN5jBC217+hXKqyubgNKGQlUPUlCv4b8sY4Kkg2rlTJvl8O34UfAU
OYX0mPfEtyrFvktnFCq4Bml34EjvgE8Nv6Mm+gxhagW0U1lLMjDtUmaiQQTDDR+7
lA/whf/V2VJ+EWuUPGP1YAgiRonShKgrHj7VMIEepG+k/8hrss5BkAveQFywwiI1
t6cKm8LOjjGV40IEpARGXmCjfDLxsjUxTH35Qui7HNmDakMRqHIaMFJuheLXObem
Mfayu+Fmd0PQ2N77G2hjxOGtbPaIx3Eyv4k1X+la0APgBKvSZY3VRlx0HPgyI5XJ
H/vg2eTlYNmEsYEy0edmEI11BO66/QHzmdLRYV+nqEadaBpJtztsPbmnwdOHYr7a
P882TIfViz/WVX9b5RNXfV3g1yaiKvx2dxc9o8+AZ4PcNVYWS2LHk/E23dHHWsEY
2ojjIaJsF6nuQSuuTRxnC4U/7a6ZEZKrgTvv4W+FhWBSbVtGw6oea+iBr8DsOWXo
v+Uk+GjnjO/klD+PukbApwunyXO3gG/05oWzmebZIi8buJx1g3SQ26UF0BrOVMZd
9mAQjnjcA7zHROmSw3dC7WNi7dzLPMzKLq6MehIi0+tcdcKtT08r6ukQtAXXI/KX
rjPAS4TuzICyn4mgv3oHxb1YS2oihjn1s2VXOfNtR4kZYScwZ0Nb+6UkDMTox7jM
bdIrj882buq1BMVWXM8DRAlnGumTFgcz21leOuyUNhS2XXi1lGWG06zphvzL+RwH
/AhmsYZb+2WLjuA7lAQ5k5U4DcQS6Sx/5pYiREp5Iny3AEfJJC36JqbAmKovfGSm
Ja9r9/nbe0t0ZXShTMBXzoiysC29rS+bpwpX+DWHSYaSq2KSCqvUxAoxQPO5Y8FY
EGYQQRoUTm579rULmi4BDoMm1bFyW6b/ZJlCN0BVwsDQNBIoAJTj2C90LrdnJAE8
zyxb/zWZAkjBZQf+VNPfPIeiDDWOJJSg79w4TGnwkGujnjoU0l0LjbwH/tewtOVd
gm/fIBMZZXwxWimkAR6XZSIOOioMzS2bJlaZ0RLS6qyCUQ/iAK8cC09JRQK376yU
nSeo2PP7DOdNgcGdEQgOaDGZvYU+R39wh9J7w0Pk6mnOuVWUG5zI+mG2U3KPR2Jb
c2FV+QVtp06e0FkJlyG0FjlVTP8NZzIu7YHwoPNJr25+UIDmbA/FF2D2qBJOzWxD
LG0iVr3txqMeZSZ9IWyn+x6PrBGbp7liMQqyPs572pTnoWesdSMbGrATwLMpu4tX
xEIapLhu9rQKfFxNc9Au0l4meTt2iYN5KToIm4dra+M6m6ZQnDJxOqWhko44A9su
nYTSPSzvY8oIWJWoALgtDdBYKYJnKUJnykmYyfk+gnxGmXERHh2SiwGW+1UJTWmb
o/7mcXBzJNf1j9mVtL/9/fVzvtutuJ1JHTkCMFnXAat1nHBE4M0RBCSjQRRfK5Fl
u+wFL8ZjPDPowfxLqcDhFTVICajhW/9rbgf1xtTk7nqd0bXcCqx3iJ6U2yjNh+3t
sk2improRwAsWLxVK9jrXm8IM8y5aSZEcsjn4ivVvyu+sn5hpDT48mRAxXJR1zn9
g1tv0aO9sowB5OZMK2L8rJ1CkqTgdnf8yjY42h+H3XcTTb+A6OmreEy2aJNWQjQK
1Cqyhv6338RIDxRbse33tV6oh3063e4OfXm4R9pVLo5gEWqE+k2cedzEnrBWM1+C
Ebs3ANJ3ntXVP7oEdGJraz18i8wykmO0EoNpFKJJaZWmdYqXrmSu6YcuBkMjnNHH
c6GtZCtprBlfVCDUAL8iwJte6W7hbZr8UWQ7hKMrNU8gTLYqhMWlesAPaaR+FjN/
mPWzVviJ5vKChFxXZZITrCNdJG0NDnJoHlw8EZEua2qBDXW9kd6FO2ggmiBcEpM9
YM1mLz1K1LyEMKwGDmbpHAHoDW00IpTE9aA4zPhF0e8dMkMNu8IW+NFqT49SNGi7
g36A97umViCXTR4eVaM3RRCtmrCAk2F7I0U2nPYZmSkBkw2ADiV9HmxP2dkqwIMl
mkssBvO6Q3+1XUSg/PRF7kT4qGGeTw2HYviV9HsK5kK9jDCpeVPCXclMLouMNPp0
g6pSRFYxsBwz1zsoSAB1zIufOu02WbO2gMDUBVi2VTUtW9HOcjc3Vyx7N8lmnN0D
JmraK7EEIOB9OQXFGrBc4ASVtKc0ueuBghICNTVKcbhNIyHCz9QSrBDECyqijdUw
1hzH82RXn+e5Z2dDPkISDzg24N9ct/ptmjfE6oS2+KWcQ7wloW61OcHXxMo9PFr3
zQJWcgky8xuKVKQGMTYuZSkfhTuYYXs6TTN22bX+Li+L7JQ2B0rAMZZYj24XJh1n
6WZmDpWauo63znCt3Q8F/6dEB/ksZhwKzm35IJ7c4T9h2U8A4lFKcNgbPLHLl+gP
Oxru5g+AZ92xMoprfjcjTkQmx18aZ2ZLK8V1DeAjRQnxWI97jxPgjIZH1IXD0HV6
LnVDlMQdfzqlaBZ6zpGuCUQ0Z/yLehhMRZ6uIhK+AdcdkPH7jaBHEWb6mqCflb0e
j3CPA0y8Vv4pCtuBjuyGfPx1qozeesaW0OgrOTmXOhHPbyorwJUPg2E9lpSxmWdY
DfAn1Gr4BWyYZAFU8LHYKqjS9ErEHhl79sowKVK0dxZwVackbXXpeMuQVay9pePr
u57bUr8b+a5/7qxDzeXriXgvAOTmVchKOvVx4R7QmFJMWfyCAP7XxbfqTB0tPIiv
tJ4NePbmTTDJeHos+W2iZZMlYU40rP6PTCblxa8fCJ49Ogmm55xf04uTx9xgZvJV
UNH7JHOeYb4tK/24ctau3eeWomZrktYXTfyisf4idk8OU/+K9kmyBKsZ2W2RbU0g
cR6iN93SdXKmRphHAztn1f7tMElwS8vd75LgZ+9kB6uyGaluvjqxQxFwe00xmHga
IOT2iS37BzrlsYGboTuUlkwfAW/AHeJcuX9dJFOD8xp9QkcxNF9wvSf6f3gesLYW
oEjYKs4uc3VoCTcCVjlwQEvUhi3OxgwwJ0tAL5z4OcYdrPVRvKVPF6Gt7hOLm7mF
QE4dI7hX/Im++DtsE1zftWkClip8RuSBJ9PoTuNC9lhWp5BDkfLMkTazmwPArVQx
hr/lk9QLslVq2U/sUQFEP368Cl3EaoyvV0rZmGpkXQtHYI9zehpOIKZoHctPhi++
Q+heSKsIduczYvUGOZjBUtkp60Z5bsSMMThmLD5lsQKMpptmiS68hpt4yxO5jaGr
FTZqhTpb76dYtlU+z4+ebzPT6YzSMqoavj4ANMnnRfGQAs/i22I2FSsUBMHAoOPp
ql9wOfknRcegj6pC59CkVjxeE9937/Z2OioCDs5lneRkWtF8/HEe+SAc7yJ6Uumu
hQqCz/KSNJEnOrAYijZ9GCC0Dm3WCypcOYwQoeCTwlHDoZe1GLzbLIlZNOoPNDmX
3jMUWuxIyfgC+neXN5rDkelwp1ouXg4DLwZbIAPCbalxV9/7InQHG+FmUgbeWM1r
NO74trcyDWBUH1liHm7Lj5GmuiwdBYccP0fbmRs+gkPnIMaYvhGv8gEJN29G+jSr
RA8cHhSxf5j/lUJw1z2swPMwTulwhYggKlH1/DkoxL551KUN2LZXXR7IVjrsgjUz
3+tOjC3F3IL18llxo+3yBwfvZpWSzEiP5JetY1koXak6BnMH33O7Yvj+p3lTjOCv
f1bedo6s0V2NvQ8L4uiwGMGt56oD56bOThSzTC2jyV4puiJ7c0GGv+yudaKDFgPq
4puivxWL+T5VXh4CcEpNAz8fLwiLqLq9rM5KTmllTD6Re3hFLhyJcmIHKyFm9cml
p88Hvjuzpx+KVGeWoxqCfxLaUgXS+TJHRAui4fiUgR9Xoh2zTvc10CQmWYeOQTDy
hdV1UKzqHTu4oqKqb2pYGKt4ov332vy6j5fIoxU+xpTUy8o1HzIXJpa9eBVjxSaH
kA4ZGVeSfMIgaqnEIo22crFGu/IxmnSynU1QmdWjIKpQ2QUBZOD7t811CuFOlt2v
UgVv3Azov17LKB/6M2mHa92VG6brak+b65vpFjaXJ7tw6SHJtcj2eZI9/55m9jSN
ASGJr6iy7S8G/hJNTkmqy7S+vE6C+s0Altqo+9gnZqiX7MSGoq5wbMxd1gAuM47F
TaZQlX9lUd5mm2L33OPCb4vJT0nIj/Kf5dINSYZ8fGXbG+pEa+CLERDcOgJqDi7J
Zzqtn4kGs1TP+PEno89sQUBiJKgOVvnKXovBzP1Lxt1U6Dhv/2YDEKUkougpkrtd
3VW00ploV6rNr85OEA6DAE6LWoezTonnqYtJBIHg9Ynp+ZL3nK/hsBb8QgBAP8K5
/p1Xy2GptsOySm/QA47vUzyrMo6rUHVwZWmwk28BAjq1gd5oLHkYyC0O+zhrbfPo
rAiw5nz6ZQROvobr6D4rmDHiKrxGjOHFGtuDqbp69FOmoXMSBZ6cKo7AeFN1uBLw
WGvVw1CcF3oqwZ8OpfIJLLQInw4iZfEd2wF69vXQ5JaZOVybvMgRIs/oHNTdWZZX
CfsQgDF6wAjwUlBT47CHh6NfR5GyiQdgXOOqe4mm0O1nsC4otPF7OMm6SGn2kFhJ
Uy2b6w0VlbPmhpjDw8+hEe3OScu6uwSNauzWxkXX71O+u0iRngK2SZfVhA4Pu8JP
qAs6yr/yA16PLkt+8MNaZqOcM1Uk/XJWynW1kJyeh42wffdoJda6ulxNf6zidBzE
dB38uLve3JT6830VV1WYB+FKWx1RTyCOllcmes9AA1qr7nWhXwWXfcTbdb2azHo6
7BSDYzuzgdUamr7KGRiT5SqGkV6ZTNetb3J3b0CMGv6bOeJ+lStZOLgAEmRMRxL+
KB3tUTEz0Ywdi4qA1kuD05JN4DHPEOZtZgdgdslstWBEgJbnMNsGkf+y/5TUD/NN
Hqv2pjkqsyd5Cj9brmOthvzLE+QGxToBasgHiMdYIvJaxTajZh/0szM7xrYzVlF2
j7B66a5Et9oU/iwEp8y6R/r79YzOONnZKDdYFsOlCsz689jAj3ImZZb1IQm8Er3C
shlonLEyTF97eSCeIlXLWmlxhG541yPE2hc1GBEGjfpfiIaLTHAXmA2y5cvZNPw9
C1h4oPp0vj43IOUMO9WDcTljxbyiBPphy7OTSEbg+0YirLQ2rh94BqFJ1BpPB7cp
2dy8aM4eWtNB86zuYIBiONqz7sa2VokFeL6owTskpc4CVfikuv4uwmTi8TKI5fNX
NF2AcN36ClhCXms2J4dx6Uo30P5M12F1RVSQATeLfrtnLmOCkM8v87LaRmkmsGNr
xSF4E+5fuXczcLnTFwD3zBO/kRyETw3sinGYTL+SV/k8Gm3GAoW7oNChW6Ej6M3B
TspYViAmKvugBA2x3PhBvjDqhfbiZAR8le+ufpxAS4O1FSLjZn9np/QjOZUd6Jmu
5797RVE+hrlQczKdDK5c+dLyk+3JrxEwuTudsgvvo+OMwcmrLCO0lHSp6deohKeV
c/GnB+BOGlJOd2k7htqBzmYACYMJpKBh27/O0jHk/d/AhE1OdJSoujYEp328oqsK
dfEgiOeUjRoIT0XIXJCpXcXqvg/iFvwD2gu8vE0imu6deXrrrnIR1cGSRS77Tvhv
WFXWfs0HUw5TEuazRVvP2GwMBh1uuTAOBX0ELgx+4UWLJgFC10VQ8Qj3sPNSbZ6k
WfBtw6PQJEmV9otrdgN6c7IZUyRFBIlL3PyYxOvV7rhQ9l/S1DrFOCpvn7UVAD5Q
6iCvKsu0yNFydFIAP6ELW853KJBBKa7gXHFbv1up5/Wep0jpWyUXJihH6jZEmE+j
fpp6IVIIqr8/g0fTYYx2MP6KIHtsWnKbF58Tr2qeLS0acT76JtCLvV05uNS9Omk3
fO3OX1OLCR83Qoa/tzC++C/H3a5D8D4ut6t5r/3JbJQPfrGsMIDkWg3DZZKOOqB4
vGr/+bx6LByeGWw3YzPTVfPVNeSFGDUonavZc7BTlgQcif1Cfgm2DTzHtDHIAD25
9xd2Ff1yLztabmAAkhnfnyufQ6rvMSsF7X2cz6PfBOHIaHL06KuKiclOhcAncLmk
Ov03OJe49RD8h3H1GP3bHEIMKIShiuUq4FNLS8rw6fIbDdTUCqCY/mUYPXNKG+DJ
G5DJ9MCv3WWR5c7PVE2w5ojysSUCd3riqZdgHRPksHb+/UCDKxll0si7smpM586x
NSn1INlq5bvk8aWiv9H2WgDGYm6x38rSKPoi2VHPTBsAOq7Yik4qtdnFTWK/BskC
vF0YeDK9Jv9DyX1HHLRfnhZXSMPLrVdgAeN/TS46oqMut/GWXL1krlaKmBho3mUN
Rm1mMc1fAhQ1IHpH6qKLyzCg38mHetmSTYP7e4uvlD30eJ8Gd4AYPiTQzSB7ZDxl
GIMAcfc5dzNIEJkh6pqIQ6YM5YxYrArBDB0l6ayFhutJoNtimnmgayp7Gybj+t/K
hk80yvdDfmRo49mp7qkC6yiXBhqRxPvRc6BnWvEGxtJNMRAKV8UG+Khl//5HOqzp
Pb9eVcAf9RoUkWiyOixVLn0lVeH/W3soLtAw9k3zQXMwB3Aj4NjUNFFmY0TRh1yY
zf5VaUec0hTpJgOBlZF+N04tsfYS6iQGXUbT3hdsirg/cbgFz+3oiuQx6i1R9ybD
aQ7PFvenzeA8H4/NoUkUmxk7RfxOPR3yrRGYn6iTPtH5TXcJ3n/1zw1XTlgtS+3P
YZbzbuR5vJzICSoAX7jXT+Z06d2xMcUsEIbJrGfGzxC5NhkVxsD7Rl+atwhlvYdR
4EIbVCyzb+JLNT3bgljihEFkWX1hvxQXEQ1H23DQ0U+lFhCLkWDyVjD/LFRsaMkk
o6/+LCwGIiykxBGppH6fM+z1Ill3xyo2ySJd9I/2bt4QurNcGurhmU6I810+E2XG
B4CQaCy8oV/rfMjnNL1zGIcqXqYzwojLd9tcu0/S3bDjldOS8Gc2/NlE4b+2tDMf
B7UUaOelbn9anDRAOMNPNN4tDPuJdXVP38npDAYkLdi7LohAhAaFeEl4CX09CP8n
JWkptA884NSMVXKHpkL/602wvAHgEygGLjE9+slMUJpFLhqJEY/e6qf4rXd/CExv
Po8YBAnVHwA/KwOTujW8AMGnIwmIbF7E06rIEFtYb+WQY8zol3aZfz2LbfoseM85
uUQKD8tC2X62RyfOAKO5KUdawE0SgR78AszMbgBQXFv/HwOvTEdS3Qvl2yio60Li
8fS0P+S5R9fSQNWI8dWXzUs5DnbSM9IjIPimh0wkrDO1JsX8xp1cIZbLiGz50FoN
zGiVXa9UkYu1bd1IQHCbjG89NvcyPCt7vFCjEiLgRl3bSgx6H74ckoL+X7G0XUVB
/fPIj1Cb+VEvT+UywYHrO9FgRPX5sRlJu7z3PJL+wAOUnVdQbeKkaMJZuaWQmSgD
E72nybZJdDUo7VA7XLCWp4yhT4iGORlcnBN9xBNGYwAEjyTh4NB7Gg2SxYpzqhVv
T3sEDj4DI8TJTaBcUqZFWKupoDlWQd3lATl9P0cbyYoTcjWxWEzhUJ23VG42E0m+
Keb1gX6f51YxmsWSrSbduTFlf4tK6B6+NhfwPrJKvnXDZa/El0MROOJlIEyL5AfM
UeYSOJRjEWil+FPChmViTMcRtXYj2w/vXRbrzCsj4cKzUbhNF8tM/Ey8EzYoVikw
oijMnn39PxFv54/WJfdPJfrkr4koiPALM1PTEKcMQBko0WxpxVbaihYpTLmdBsM2
FJ4qSsyo0c3TKSWPGPJw7EspUm0yCxf7ot7vSGLJl6lVqTFBM1Kd2YOCEnweXOjw
pJL3nkN4BhdXY9jRk7dvhNlZtmFxYugzuLWuFSUWXxoKf8xPhP5AeBhWmWH/PcLC
lmcQpXumYXPrZrf70YGU4quP9P4IpDhrp+fG1imaYMlI44wVFJdBZW12ropfPByP
e2MkXf5emOW2olWSmDJCT3+X4IAcjvKOcDIyxgfjm1lzEDHhihFZUQO3I5Uv7Ncj
aIRGdrKCABjpJ1TpxZFdqQyAw8JPe/dlo997raGOzx30wcfheHF44HsqOf9UTI3i
EAYJ/na5L/hjmT/JpN7woa6S74R8NwKxI/n0qxhJmN5JIVY3JkAiz3editDrM522
1WL6hVhLV5g4blVht+IAfiTDDp4mSVdIq/gXEXVY/UX+Ao9md4hTdBugS0bF8MBO
kgik6vL18N2ZgEQp/JSI0zzbApuXHuPZemfkQl2ERHq/3OEr5NDA61agprOPdeAQ
MXjRrE1nCOag79oPOj27gODe+BpZzM9RfAL8fkzOVcdBF/swZSBaqqCskmBdR3cQ
a1kpI3TwS+IHT/S1uov9m+js2a1UU0tCB+mmPBzG7oIWgPtjMiL0qhmg55ldkiNo
eZA+2sNZO6py5zg+0QlQxNlDiMCfPxZ54Ga9c2S39WXae3uBt5Hle+yYfaBMFONo
5zHvfCy10xpna9raJXjU1hIs+JB+50yg0AEAGE4yBHjQKzF/qz+ANUSXArFlHKvb
dexUBpApx1IvPqHJQlQrQVH/01n50O+0YF051sCwbSUzaymYapU03RWMlupWnfjY
qDRYFyobMnMUxRFe6xv1UKl/bGDpdCx4twBAdOR7kMNtzcYhpxCnna+IOvTmRwgT
MGQRELaOp3yUnJ3ZejA5W92OJlf0zv1RrmcBSG1eo/Jf5BtVQ0k4IAgeqGHxWP5g
tsER+/65QhGqr4Vqrp3gi3QxeSR0E9kkRSNPPyOfQm9nfK7YterMzLpTWocpoa9G
kKKJCpzyMLbC9YUlQyzR72w3KyIYUgxlukHfEbKiztvjxAKeP6Rj61J8+/ex3rtX
XpQbsZwfRagVhScvmhuUGYC+3fIwL6O0dlvwWknuI2mgQQ35qirIsrHdrWPMikGM
UFRkxvfhWLlnaJFjiiMz/GGFZzdz6dGmlO9Z/ap6zKEpHexjRA6Np/N4/4scNtLb
74a7oH5VLsWWHizEArUaMVvP2lQHiyhL2Pa3WxzxEJcc1flrAHayIVTiGg1cXNhY
Pq8Er/51ujr7iFN5PkPWlXHCcmVtyQNyXIvVd4/vJ6MVO6UbLWhMmdsl/JIDvMM2
xc7zlllvP7Xa77z7PkMLRaEF11nh/ZsynZlzRVQqT60bkJBPm07xKAKnwFO+vocp
b6SC0Q6Hky3i8xfNHS2ubJPQl9W4Xc+GWjYJCmoGzTUHepz0h3hTLX3aRKeYA1i5
gGko/EdOQJAWgy44alULurZxUrubDMktQE8g5L6t1zu7WV6kwP9UFbAUHKO0rFO0
eHNTQDft6ev/ZF1oemXyINXWl3Ds2l3A6u+PXStt+wn8kZ/FMZ0osKAiwiRfgEtQ
In6n+HPs1RuqPYg1OfLPW87LvjJYJ1lAhtbIWgGNKH0HihVEDPXsXVBmG0f9uXMN
xejBjQhAj9I8ORQRNbyceaqcGh6Fm5FpTLTHAMibIUDpi/fT7+8axA/vQR08X87b
nQYIbNMbohqBymCoLMPuD3ZqnGzHzIVPm4yoisMC7zNI6gFNs5s7PsKiGdRgV4LB
XWb3vhXkI3HFHIVotOI+qxCfJea8k/rigazCUNIKArr5RUIKMewuf9QtK0+wmwOd
HO4yj/URnpT57QdOfDG2O6ElwuyF0EDP+tXPPoeJN2CbQ3JH6kSOoY54TVm1aGIy
CeON+JPLN1WCA/Hpjvoj5Ma/M5cUSjQX4AHgB/LQT6gSzZ3lhi3Lfl3/B1stX5J3
kMXJHVj0/kxJjN9N60sexqDX6gExnDAMP1kwLFyRsQpZJQJFbQfS+TgWu2Oil6ED
aT0ukBVWUCY4zUm+oiGWi/4kwhtDNiAPnXZQ69RqVCY4toDr68+eL93SudRIGbKV
+/bxWQ/FNl4krurAO5vYX6VJB+aAG4ieQwS2wOe/1qbaTUuWbenCXsujgRdbYW1j
ML6oxWL1wY/MKEAgE5OKWABkTDxCxv+zNgNQ8u6t6Jzhlkf5c6svEfus2F9ilFwj
c7JjTe1aWHAGxgc5OCYuuz8Ry83gplSB2Mry8ugzwzyBNKcVb1H8lY0Jxi6jRvHS
SgBP7owgnRBoEjp5mXAD6ZeMRU04rdgC9nCxi0ddBcINW1WVeUJONB0glgcTDAh1
SHhbMJYDVoRyyxYD8wNvDb8yi1JnFWrwp0NIgCgQF75pwqjfrD/+TRtfhFeePdtJ
kp2yz+ZU1YOT/6DIQCsRHnrqcVLCxVhOyrbYvzigs017Y7/dUau/ePMXEyNLY/og
sagSH+gRkFl96XE1eSTJ+5ZqkJs6BBFgFvpjsy3veQ97fpEbZ9y1whVLvdbeuqZH
aOSkoOh4gFPzd8uLP8Z+hWWJpw9gHhAVaYRtIL+33hdXwKbSSssgR2KlN/3yP1Xl
w6HKa3j48L8rjMjY7lg5Tue31UTbjcLp7tCDz+cNvQyg8gozfkEgfiNcd+yNJwo9
US3fZ3BWwf39cCregaUcsJpGqInBvKAe1xJzmSIiqKSOqbj+IUSfletqNY7f73JP
sTuYXoo1iKxvP2Dce8SEYWboQrfm0mAL+cQoRGceBC0gDJgUh5yXhJpngjyGSKW5
//uDX7OuhCIlHmUi+a7BWc2sKnwbblz5yX22RgMmYKJlGFl0snRIdgF91p4dARSE
oAEcDE0E1TAhqQtrsJMTUXqtpEib9KDP+ekYSkpICEgRaPWGiAzQ0cp0xpKRHIwA
imRQIBbJsVQgqKB/poJpuw8f+P9EK96iaorRijSsbtXHXet43MUgUA/St/ki8f5V
C+9a6fDPyzqRCmB2t8nhlIK5nAK2tvq3ouGmHNYF5SnhtQZSSoYAG6wyjqbaoohn
rajtylYuYrhvHN8OOMxYqTJ42jTTVYBrG2GlrDYke35SirgHrDLOUHTKZ3/S6bnj
HhdLPsOvB5wgQdKdG90R/UkHWrrHIspgARM3pceWXwL3RvvxyKK8vTuZRkVCw9qL
D8OnjYFcN6vsH7M2MPDIlhiuW9EkWSgCLIFacOo44NDduVumKftOKOWsZ7wdCO0O
n3Lhu0+XbgDwyso1Wb5CSOuRoeB9QutsJzrLcuDBV9hNSy0vtq9fceENJJFOEZ86
dsZCR4NQT5qLwL4KpOhfi1GKSR4pgSAi1iZpP+4nuLBrKLpck9f+ZCDeHDva+a+u
GrWEcde850i5g08+J0XgfPq96rjrEgVyPmuw67rtT8KuqASB0d9kEk4HUhkx/g+t
F85y+Dd5nV2Vveufj0tcGjRTtKYmj7LzBziHVN0OyWPOQFmaUQpKtJTwPtI7KdKX
WRF5PDY3+E5T0g04qu3g3ZL2LX1VSK/x2SJIn+0ky+cyrosAlsKuQMm7kf349HqL
fXPkJsnmu0KXNuGcHPzuFGhRX8HYVSjdut5MR+p6Cn7paFSudWRRXnQlpHEgX71W
NqDQxJeKaZcurivfnbZroyzCZVzZ+zfP7F1gN14PvAuf7JINZQRHCVX2YC6qaIra
HhTcdCp6vOj2IvpP8kl7nNrwKSiLmcD2zf2R3g30hmxAwjYQoZO0mbrKb9U1+gFV
7Wit+60uVlOoIocUJM6Tc63JfjVGd1cyjAMj6UsvxSbVdYllUaPgD63CNK2VEQGc
zEIfRbACQu/MrSVt3Ec3cntOWS2VFxtZQb9O626gyojnNQxPyNk/M8zX50zPDyCN
lI7f/rjbbksWFOrJNQKRetISuGweVpkGO6pbr1rHok7yUEfuI3o0eYAN1+uMq45/
kNZR1wqVksOp/gENbBHdbq5nblhg7lNO5LQXnKF0I4irP8hD8NHP1y3vivkovWAk
bqvKVOVN4l3GkKrB4+rsZrMcPPxvUctUH9M2DAlUL/Niivhy3fA4/70aJXZ9sNeP
B0VE//wuJ82oTEKSyRKkvzea+B65rdVoUdH+B/iebEC9SHTpyv6basKmmtITCMSt
Vd3jnpsNQQ6eWSB5Xm42sveFXn33N+NrnYdsVYI5K9vyEtHQeR5GbUwpLoGK7Iok
7QopnpdRh5DnfTEn1hhXRGv5f9H75B+2Uuj2K01x1gV9qQ5B+eKksKFJdnsrXnuh
90DEPIsgX0+Vxcz6a4BQruChiOnWIu7egkvs0fiIFa2MxIjk6ZH5KuivCvTAVz98
cFEK9x3RwegxNN4AopSCOETB8eh7h3v347Aq4v226DUZevxRy5epM3L9xXBgdZdQ
wFLXBnfOcjX9jcX2EIApZICjOeWeDv2PuqTcPeTibwD08xB417AYpFiEUIQ1BoBD
Kv2p5rj8ek80+Yz8qF7/XoSiqhmMfdjNcERs0kTjpe4kNFq6sc/GOpDiya5383UM
C7DXff0nl+8ldFUmrOfwd/u1RYnYpQrBQkT+mWM3L6/xSPhur8GBq44SQ02LzDqx
MZmGwFYpdorpfcbtPt1mhANrg1GqeE19X3aFFeYjNXMAt3GpXwq00hYowxXAsyFv
Ev+4+aQhYHCyUB5ILNpshwqWWu6hl9ab5QRk/K8EoZBHxIej6+jLDzcNTjlOr4n3
EAFIdOkcLNuA61glR9scW7pTFBDAzGRTedembXwhjHhL1re5h6IXQvZKKxX1AQUc
oX0X9Geh4mlotBMhP/lxXnXkkh2/JKTARm/ouTM8Bkv+QS6qfsh+4022e0D5NCts
uOUlo5wU5lxYFbc6FW8CfQgIl3l70jR4zgL7WUT+9jrCss6p85tcTxZlyVUzKE/z
Q2wn4AWmrwm3Fl+qAcbqD+QJc2A4lQeVZXVkS8DojEvCNuD8vO9AXnRhdVCiILvc
EN1+zb8gWZ4UzghTUjQR1fJ4Ywau8J+zwxBS5D35OnYKReJYvaN8uJ5YK+wEUAqa
xub6rF1VwgcpXA8fckD6sCUPaEPfD5CJ2uVip0+ge6VidQSxrxxCFYKkFKK8XJFz
IDb+tTOCU5HX1zTRj+wq675dpa+T3cu0iH2R5WUjTnh3b8Z5jDg7XD2w5YMWJMOm
gHBJwq9+pshcGwkdKI1nbOHzB7XhbYKYUtrMf093OddNOvMUBjDIOsVykyrM8khV
2xXh2R66QgIoN2CUVW+EtXFUR+1gbtGn2fDCEQGX4wIAoebR4UhKFIu4HNm8LdWz
rhugY1zx83gOXsftL3IhunfyLQwet2RbXWNx1dlrk5iGJGthFSDpgltXPxtNLlOS
Dbb6npxEq1ZNf8mEREqDAK4FlcRHbj3IamgsBF/sSjGEmYVKurECPtiw4UnE1O3S
L/k5JJkBqDk/lNLVw70aX6e3ggiNiq54Mf+JoZhXMZ9otv9pcLT2kokK1QfQn09x
PRmDC/iGhYfYdiDKuq0JtZb7CmN5G9TYvXv4q4taowSnfIAuhvs7CRHBi5N/0bWX
+JsgIzTSSBWKOIQVl7kvC82lbQ7lSykzxJY1Js4h1nFeXOvOxdcbz6wDet5DPRlq
tLvfe2qD1UZ/yrrE6cMa6xlUuwovmdV2IM6PQZiSV94wVlyHnhVoB9v5rfWomPGS
cl0xOSckkny9Teq5CVfPWPYS/1RH1HSKPVF6JVP9LPfzNw4btcmiQaoJa1AWgckN
O4p1ajsWRJZTZnlZkq8hkQDTuQFJ+peg8mQNYi1fVy6//3dloOutszqK52Vr9fhE
bCjZBX8iD5NKsUZeZerWyFes69eLHZ1l2IACKdk0aPgulpjIHB//h2ADMzgGGjR0
7DeYQ0XNaK1Abv1+JBvbOxdL/+57f+Yuo43oux6uDMgYS9ZnNzuZHItFa3LWJfQw
ifZJ8dCJtqf6newGgOP3tWa0WJi0OOkcFlIAVch4rAnKff2z+bFW+sCThOKsp+ma
rGKurGeZrKCoZLcwiUay4gIpFU61PID9F9X0XoO0IcPcDzEDajCbQ4kSha9j5TDs
n0lXrvc9ye3Oqr+D34u9kCC1yiyFYXwMWlSMG0c7e90WJxx4urjWiKdTFVPE7tOX
5nL4iC1NLRvFS/70HGwFF1vxWmd8xquHqos72I1NSjRuBonyli4mywh9LBx8kjCx
785K1DkN709K5aCEEQGvKZg3tocd41e/NnWA0obJreVsEe92j0NyLM7xGgXNR7Jp
ZnmqMr4f2aqUl560SSHTt0+qGKOIx74isOGEGD0TTuIjcPXceE17YL8CxeEelQwt
HdXt5Qwm1AhEHkH8Gct1AU/SR4xnLg4YJbQUE4X0Wz2uUawgcPd305tqCAJpJoe3
Rsyt1FMfBEtN3Jsr922Xhp/5JOlKC+7Ea/SegBung0n9eNJ2dioiyA+yeZb8O0pd
XaGLAhmoc4XxqPNrPxUDxPnPPixZICNKh9VHYx3uVpHxcnqrBPzNG33bqdeWxWWM
paOX5qidGzoE509Vag+Ae0DqZHpzyg0kLUoBK2mxogdBMyQ8zq0GQ9DestmpC1XO
KMWraMgxutqBD1uS/Vw5hS53Z1kAHW044TZbF6+lBQFtxtXthZMYW9pOVd3nJNnN
vsInXHLMq/1n187bJZ+UPcPzoKzOG/IRN+8E3nq7Pj9/yCtl8Ay7DrRqNfgOtZ7y
8GOYYBys4tZIXt7sRc/iO24MEzu47hhSCnHLdeH4uwwOmWyhlvu8QbLIGn8XFopz
RjyIzavOypVRvWTFJi9Zd173l6WWYM8RVzUxklIqginMm8Nf5ObL3mvlA7AE6L9O
ktzWChcEZ+JxX2WGjhJU0hOsCy5SMk/fbWDzqmffRYFWR0hcae+xqOmdoYfTAeAV
oI6HdM/WLu1uCT5Ja7BIuor/U52NiP41jKJ5rWdjXbXzNYg1vdRNxXhL3hkZLOcK
jZRDAWcLyu8DHw6Y1KKrYdJdrpwAl9gdVQ5RUxzxBSYNdAPTVzEEFw04J8M7c1IR
06OH6xRdKWuH2ddkAH9P/Z9pRQ/o2aAwWzx8im/L/iwAnDXRtdI2M6+5RGbgVc8x
tMlnhoIEowc1XPWUkrN42N4H7+jvtzkTppkrsolBgSYKLpWtItuvuutF4DafdH8u
fMCaYFGOnqHZsf1bF9htB4qRJwhtVtVAOF4skFyGOCCCaeFY3siqIvxowdIM99+h
cjYUL+eJoqtKyixZHakw1VfK5eLgAJnOWis2oCQju/v6g+FaMFcGWDFSgsq0u7qv
LaEXStc2CWXL1m3w+IXQF/53zse5LO6CYbEYOtTO29CB1CgQ0G/0DSoh1jY+dno2
dFVINUH9P+toZFFUxrKHkI+GXQa1XWDkxfZh/IYzzAiigG9H//LGc8oEi3JEz99m
3XSe7fKWT/A4b+9ETMLLN9M7E6eqim/Rfnnm76ILfXtTkJtChVY5BAE1LAjNUDNw
yQbuY7ap6hYp0kWu0XA2e+7sSIVy6hgGmLP6o9xoMjYg1s6fIq1/+N6c6d3ZkIWr
tt+4GJiQvMnYQMT5DQBI4Z5BB6cYnDnY3zFQZzbw4vi5UutnrRthMWc21ItUaZrg
OB7PILfgnNqYKEkyxlDmNtbhUEPvTViA2YSvPV2P0QdDYTTsj80tMrrHuT0Xbbrz
QIZatUuNY8I/TsI9u2XNLsA2PQUXiyAR077R+sdXLJaYg5/wJ+e9Q1ptxBTmp7MN
mOcdnexuEjhKni52o11KFlGCS12SfQt1Z07A1TyYzqHIlqDjQJfvK2HUmFi0qyOg
f50BBCzm4apNX5cyBh/Suz5Ti/LVV/2xdWs1VeCdhsOSBSQ1so5zz+37COdahvE3
Y6o4uC4V50hI2aSDPT4A4gI5/9V3j0x+WpYUyKEDZRHtv/NvhxHf0Z0U2JIUsuST
SvJln7ij7hogSxzNJS11sEQjYqGhK/9Ub4U8IhAvXZC1ZRJajEL1UKTJx7Ioag+j
GxUOJyZerDunzr0ssZjHvtUhGAOu9wnPIUYwn8USgyxnOIbVo0z8ThDHabyx3IWS
QNkhuRBH+MX6qlqNGmD171/pMhqctBJf+Zwspup6SGNhvF37YZslYtK7De4dePHE
5IPRMMH9I7V6iFY/bCm8gWat7ZW05u3yV6Ga3dWg7SGNya2f1aECUDENRETch7UT
w7ajsd3wBhG9qX0dTmkGiEnoUMU0ULjRkF1rfPbtzX4W5Z0NDbGz82j2hpu/u9Yf
JMgpX9K7HqSWwoDn79th+W6CAPOh+yPIoTnqzEZNq7j5/9SqtUPsT3nRV2ZpK7yX
WFc+k0mV2PFCGVeEn626cFcNP/fZuryF6H61FQzVdtOj+h4GuaHZFJQptlApSCom
mBUcxWVY/B5IuEvoPKlIwKdHlrKN/00yeH0C33YnNpyiXIf+FKQQ4y3tzOrRoi7S
4UcclWt+HiV/tzgzUPpyVN3BWO70qeoY2X9NT5eCafP4KZGsSrN0Zzgk9fqsCT9d
Q9gE9eKK7oXyInbdWvZO910h7R/rqUzT7LbgFUPefY/UW667UTCDNlJhvVQnYMYr
kbvuDBcMV562jvMAid5TkHZYRXLQgkgiZULKa4BSF6ZsEjETPUNliDoUIB+EYMrK
wiv3rpcFFTgy9jK6IcMp3kpElkwbNHegFbyykmeUNp5OfXJHK6mgNl1Ba6krjec8
vJ362AoNCkyntuVp0A2YBMMB4lRMcI8grdlACBzb1i1iUuQaVYa5LvvG2AcK84Fm
QgQguwN3itIdzm7xOetQt+clBHPWGlAF3WHUclQX4dg+mTy5mv/h6ZbZgKCj6+WM
4s/6kehhhQXOno+vLr8KLDPxPAMPAFYI20ZBbRfRcRezDx5S7+SgK54qR55xbZ9F
usDgvZ/vWWGLJ+2G/SaHm2GJfe0TBnVkhpHczStZSQ+rz0JAXlW4nH53Qn3d2QkE
nnkOynoY8Pke0P0TNnA3EA0PvkAdDuoeTT7rSHtlSaR3uFnobw9a15YvEw/DZ7Q9
ey9EDcXjO6DwKL0PUltiqT1U5BXh25Gn8w6+tf+ph/q3En1tgNb3M/cvNc7dBKtK
JSCGZxOpovZEMNUp+RzyhR1qFXpGtXCxrnLUW7srUg+OOZYF810OE1HuSQQ/Ml8l
iblPaZnioRYpZoWIkE/PHyte361dAwiicO5h49vkPOTIaPPpmwS4nYJtYYv2l5uv
++K9Ip73bGNb8f1rHeHcvTTvGzcPmpiuXiyULKD51HFm2rZC8R2KVXXL7XVhdN6J
TrvZ9WEfqqidz2hUTCDicJq/NI7kR9nJRCYTNLuqwOMrTxzRQsKOTP+wm/Rhe5DV
eB3zWXI59he49o+x8TU7NC3lyyNwzBBWbE57E2JYmvzDxIOakJcHLm8vlCAgHBxx
K3nXPis4ABT/9/Ve32XpsmfnYdXwUwiginZUL9nm9gmcC0RfEjZQ8BuDO2l3JTr/
GkF8TzsDQm3o9sbRR94tJQGHrCGhTnRN3ru9sWCKNy4JIyNCe8DhClPeVx0iE3Tx
mY2Y3Kt1aESTFaqGZsQOjSugezicspWLcI4tlMnE2SqRbrjnNq3nXYCBkg2Rxi5z
KhycVLBKECzVN1VdHtWuJscxkeGHkOLjr5gubZq/YsMEgFQu18cQIjHKAiHE1UFu
LcZzb+CRWicaWJTK5uyW+Zm9k2Edv9yMPCSvE+lEcQpTLz925XnJkv/GcQEt5GTd
LslYtYMW/oDvvtAaEkblc7EX+isGjQRKVdIi0MQf+HAl8f0/T7AaJitfIRkp6xR3
SAajTCUIrSbuPMZS0g/c76Iw9fDgYI8+sHdPKoqobDWi2sDFadWEJpdLPSH95rgd
P2HmGrgmt85Ii1KHl4I7TEiWTXPGiTTrizqgIYQkykHtie1OebM9ipOKoA3pMWMg
SJxdUe5Ue0vG4z6kL/TX0nIJqaGkrQQCmhXyYFwNIsO20+dgJOSLbdh4mY76bK6+
VVM0eTeVBou5PUes8Qokr62+2aH/fTmM0mcpVdvS6bts2Dse4I/yV8A6E0zxyKDZ
e3/mVr4jQD9bhptqjvp4aR0Pzs5155yNcvLyY+rJu+3Y/Sl8wh9Z21HqG9REOQh4
sPuUpHOb6NAzMBo05pTYU3eauDSrxp4yQbdaxsccVjn3PG1G03DkJ7rrB+egU+yy
IBHEb4SFy48ULyaLMpMHG4a9fjNp9cwtGoLAbzl9JCgFUMPs50hGK9VwiB6UYqqt
5E5oUOXgfTjbYg8dDs+JDTfR0Ej+A7Ou+lpXF4tRTY65h7kxH/JgZO5uCXFAfj9K
ZFidCCw0ykUi9OBoqlknwyeNMIwZlkCNpw+oY30hw/WnWtWUXLs3ZFYP50tQUjlY
uGmAZLoe7DccE7lMk4OWUqJkPQFS9EeUlFv+UugZlJIuwRRF+QskrJq8tIvH3O0w
tom6jfddMaQeKsDnDoWXJoUyKedb7TT2YNl8JdwcYZSPe1bUHQdtQ9VXCJzcQ2W3
qnQQl2vfYqN5ZBsEF20pVE17Vl3B4O1557l4YOAguzPjCvrdGsYsvXQw17t/L/gv
CGF309hIXlK0YfRrXS3qeyzqh1xWuXUgom01V1qjg3PRupkYZnxkfwGOzIauM1AE
7qGRiMFhapVLafQS6Y5xrxOY1vIPpIjMnrDC4JXI4ydwQIj9cUMWcrz6Kx073Zpj
lbQmut6/b19+rY3TBpdgH1MIEUI/4+qcREA69NqxlSY4CydUfpFANeDMSarADoHx
FuUJ5BIVxtwBgW4+38OwecCYrjLehc5lb+xQv9ZG9AOjEL+v9dXlEh/mkLVPXuTH
pZ0Amph6sx46P6atfMgU7nNmPnSRk40PZtRAV3yJmSMbkICoseZoWCwnKB1SoapO
CgRRs7ZjbxWJvXusKdOjtHRrgj35ckAHbSI3h8C9dBpfoSJgxYJD0NGlpomvs/aF
oABPfcJ6f33QSTa3BYYxJT+eK4QnaFmDwVIu2998DR/vFTHxE2ooy0OpzLgnKngQ
nTVwj3W0P5wuimM5VKqmH7hxSgnQtjfk1SBXehjCOgnEkpNKAl9zNqff7s9p9LD8
6GzZ7h6rsI7UVz14g+OYYKFh7KLvTrAb1j0MRh+HcNYPeuPU+xDbZ2hY+5E/oAMa
IdMpwqGpFEXL9YNpQzZCwN/a+PgiBw3lj+aANLn4k3P5t3Mt2eJO7LuGwZL7dUgu
NqX/WzH4bCxP2AjuAkCnm8MUcpBxJ+iZ+qE27qfhMqP0Zr2Y8pbqP/YkgFW5MCcE
EUTSY+/mJJpJ8skeXO3CGiJcX0lNIi8OgC2Km7ZAuLjBnmWu+62Sa8Wmk0tpzl7+
t2aqu03hUo0UJ50IsGqt65wpxUERhHtJFVLFnzdFqmc0XWKCcjGbVjF2DMpyM7vq
5ousE1+LxSk0PUYfhg1K97Bvn/oicZytKBT+4nQRRh5GKepIGvkqZal6ML7tnyRb
lsw6gbGqN3tT1fbEFRCWaMF/3vEhjcT74+ilOfxLKnZbDxXcw5Rz0hYdkAlAIWMY
5+HC8OHqXc0TEuboBwqbDgSCBz5IbJN833O6AkxyPvnRITMETPm2w/bsGRPSXY9o
mu0CIFmSvlrpZjhS6tO4HyNM6lNgSbpF2dCiW7H/ntgaPLJexj+i3JjzeX8pGs+c
Y3GudeD8pUcVP4v3VXKZl1PTcHQqsbevRHLv418//sSa7a0jrW6ttzzpsNciT0Oa
IXocqcnhE4298D124Q/BROdhrUJP7WyhOUT97nRHoUhwipRfcWPgWm8SZBwoc2ZE
rCT0QG49bUsUGGF3n11mQ59ozHuPTz86QbrzuODVXmxd2UbWu9xA74dezU+4V6NW
iwv9Xhc8NHu01JC/UtT1XRHzhSNb9MiivivWkWRy4tDC7DYKQFxp0LnE6YU+eyMG
H1w/9T+kuyN4KOHxvjmMEVfltEv9L13dTti9YItWZnPi+1GUxcisOUXXpVaRy1Ko
ByMDGZnxbtvk0RoH7WzBcjpDVVFBqqdi5LeZMX3bbDLkrM1laX71E1S86VWnxeSC
VKdjAMNZ5LS/RDXCX5aHCGtnZ6Jyt5/ginGyAgt4qa1Awopyb0VHIyISYU+wO4J2
3aYY94PTAiSuGZuSP+n98Y+tFzAnX7ZF6zCBbQK9W8rfFMFn12dFlK0P+npGI0xF
1yPYqitAFF9puqSQKkVCa6chMk1si6XPLVT589INWy6QEVxMSCU4wvmTqOIqbNkF
Vgjg9eKsw0QSVuDkumQpmtiYdzoD1N849JBr5+4Ptfuw8WqCoaBCMuhLV9ucORy2
BqA35bhOGH/bhSPR6YOt0O03bKydEW+1fZ8AkVOhTaLpLLrsYOw6JbeAeURDDlW+
llHmjzgNxOVl2+b9F00yDyjRMKuBl87pa+CgW/bvu6U9DOD5llZ7h1woEGd/T7EZ
n5jMU9INRCiAyCGdnfa+OcDKDPnYQs/j098Qh6HwQQSRiKFoNHlST06bAdXEmyeN
QLDFek/FLSYDyIQg2qiIvh4sut+SiRnoPAkV0detW/Na6deffzCzYBjp6e42c9Yd
f0Qm6LTdK+0tAsCom0zhSzcKzAzlXYEyFFLTCc/CTtg7MYsSFcCNZ7MUFfLWHehC
fCfdkC5le9l8miF98NiFZ7+ZoDBVQZlxwnZHwSnV70iIkpJXuZPTiQxOu0+NZKvT
XpTfWGIaPJZx57x0WSnpt8CwJ6W+OqTNmJ3/YgmJ1nod4HmiuosITJbzH6K7zXkR
4kTXgXl2GdmEaNI1myfF8rpcysu//zN2l6jgh+X/7oO5IJ/QJVdOGiYpyfj5T56Z
PTGQt+yRkrp8IXuqtVwbLdj6feEEayQiUuwtZtrc2kZMjQg4v9n+LRkzNmyr0wX+
Y0Vju1X9XH1JNt/1++QvsEQAZNnx7ApAO+PFuuMgfwOy8kzhpiJ4qdr3YTKsL0DT
hKDV0ZNgT9o3X/YRQgUNwRFBwkAwYwzvGFhZhcUVrHIm1sNOulPo7NXpx775nsYF
kYeY0HRvLQsHGMsCKOH/Dj5Oe7adPP/byusLUJL/gFGp3x/9jDeRuBW9I3Nn6h2n
LXqsC7Ju/u3gxpbwo8xttlzW/lKCJ31d4N3QfcUyyuBA7+v7wgp5WlbHCIRLPvB/
BKoD1ESkNvqzJlzrmSpVTSysraivkVry75nIs7GsfAEHSYAxf+oDn3jz90vPT2fz
aRyXb4/K5uMpiS/3i8rq072pAm6cfJ7n+WAitSiQtWSLZ14gG9tm0A6NosiCkYBs
MWiFmy2QacXbJTkYLhDVBrg19qHSYc/qHtevtXiopjKzFLTw3lDTN/9hMC7kgI7i
HNrKlyJv7ZCrlXXN4/veZrVGMueBW3yBz1JbUfn+yGwIunWozTm6ucRuY+ATzTj6
yzioA4Io/9UbQCF1kqiapnfJkdN+D6NEy9I38qzxdbGy2M1F8xTk+lIePH5WXqVx
vcCPEz28ayVKfF2u+7BTsCbUGwHMpM6QNuNzwN3SkjP6raMVFxYY15DfJzS8o5ow
u/sNhPa6R6i3g4CGnwhU2edb9YlpJSJuN7opCrVzO+8SF09cljAxGm9ccpLrm4lj
e5I9jBiIKDhACTB9jgQXbOuaMFxHmvm+JvZTqUZRioQtduTARtjM1lAJhbXcqtWa
K4lXV53/dOShB/yJfIR034p8cRe03KtL9cXgG1Ru/uNMiwZH5dj+xApHNur3fxZK
8tFoinUOjDWpeJccoy7BmrwMluDwEzp9BJLYQdA1O2DPhmyJIn4qwuFG/e6DYcjq
wq0NDzHiUwIClGPvBIv6e9KQy9HoXwLbl9Ug0ksJxolI1W/1kkJpw9Uefaf0h0uH
HGQmUdKKFglaLXpETPcgYign3IxvGEQ5A9Dp35d7TxtiEKvaEGLlZkOQLvwHHOhW
tVtypIxB6QtYegVubhw5DfPVOvCq6Hl5laIdUqw/eOX1flWRuZse4uGBu5jnY9G0
YXhzbryLze0j9OZewIBmWGKn0z+3P5MUgzob2OiYNRLy8Bqzon8C1hDw+1TrUwKF
ZHT0dxy+wJmOQZfNeexQFaVSutOwIq/rjhXGNAtAHrNM9MzKnJt4mW41LpyxtoCz
yKz6HxhXYyffArM56jSVMxv/HU+HhPt7976qmF37YHYJtmkELTU7w+Wc65yXoj2b
U7XOX+Zka0fOBfPPx33DFyZmX4k04wV/9WyMFOC9FlMsnt2nfHOoKHWI/EJXWHn6
OTSlZApcbUoMbFgoKWLgkKQhbvihybgp29jCyix+fwO1nKpf/5zQ5AIHs6vFSKUy
ZIJu8deggUqexa7dzWMMNX6CikQ0oKW0sTU/EsenPZWGOXydmA1QwHQEPpMtOchR
1fLv8Db203Yl1tw6md3mwnLnesODnzvQtJO18nfdHpxK4TQ3h9ROBkkEX3uRzfOt
QzsRkTE/A9G9+l+0Sk+cAeJCTXjtosx5ckvhqTPAPXU5UXNhvlcZT4a3jgULDdOk
MgsM0pOWYdmq9mtoYI0H0CvJcFJBlefl5rtrqO5SiUK/H5+AcCQR5GFZGIN7hrNG
lyPSjGQALjeX6jMItNVn/kcXCNnMP+bDQXA45AwfFIQi2Dm/h3fuY1kRcdyZvuJn
6u/zkJ+4wKXtqF2wA1YPHNbwOpCqp+l4w3Ic3Ek5hvqSCgPWhXabTjfAEcYM2DeB
d4onhg1T5SetTYgec17mVe65vX98g8Y5gdwGDVgPYCvtZMrbORVM66mTmkreAlF9
2Vji5KKeCAR5iBfEl2WsHMeNucBzs2971dmg+wqpJMcBNW3UZsvEywxunfTIZV/q
I91IBROsYNk2qmTY0R+qWlwsqOIG65ZTHXFu4q+7X4D/hRdGkcPTf/V8kSg92c59
/qlJLWVs2Aa6OjFGhzAEl9gpClk/aoJ2bb2iHwLTt4iWjQsas07TyTQDNPwwJyfh
wrHyr5v4tbBl1iPspArTFYzAGWY9ajEwd/4zgIf96Mbd8t/zMvkoc/FVT/LsSvgQ
VQ4+6IXaCv5zQr/LX4y8grEUyjvOXY7B/GvNpbqb57xkwIIOAXP/o4weXF6TQav9
Zay5UYoSLPmWRuKOx5uKD0mpkTRTNyDp6UDWRNXMa9LnPTBv8yXG3O9r40oNeckP
b6cTCsNrEuVhGlpRedZX51jsFZaSAw9vgi5DLjAZ72cHf87MuEpbbf4g1qZOJKKq
5/FVRu3nkZb+s3g2WA2kd67lGfGVGCAoXvWtJaLhf8DB2lFEai4ecCHxIousAcA2
7yedm0SLORSJKYtyEFq523Npayf/WZX/yOgsUwNJ1ClS8V7+2ES7GjzTdiylIcrS
Fr61wO7XUVNC3JBwN4v5mKmg+sGqYQqf0K+BN84qEY+WRnabqprhPrACktCyEc/Y
HhPH6oi+lBazIpJRngPSQo56UGqSlONiGk//DArhXwIfIWhzPCyJPmhbPcY9C+al
x/EVuEbuKTxT9TZ7MxYLKAe6B/m9fPpwKWWDH6WSI2+78Rd8fjKAOnQlX1RMub/b
aair47Gfjn9ClJHlezVVr/vwJxTAmZtA5HzzCXtWkEO9MFi1+8HHQrt8IE10YfTQ
/4szhi3dofCFaSPEwepdrNorpSdYU1QU2JubwQQYctXOOlaq6vDfDj5bre3x3UUt
JjqF7F1Tc5TK+x0v3JBwphNg2HyuMu7CWfps+Pu9J6pL0lE4iMmYHxhgd2i4wZVX
8AxGSgXy5aAy+duI50z34bN+xEFjeQNiCuBsPngXrC0SbyTany6JwtxQcT8Tyq3+
JPcUHxxt4pTiAgFSAgT3RfyS3IBy20YW5dvXUl7JnxCR0EDqtJS/sn9KWskusSdd
K5a8GpRb8UhacqR5D6O3sA4tPpG0jLMHP18WWm6l/MGxI4BcIHEzLJHtycS9apKW
Js50k/7Z4BsG7nxsVQfpM9HSkrRUrmas6NtUO1AUdGbtoD7AZjyBaJcx/yPbJ93f
lFaAZK4ExMhYNETPm/AiZidv1UwYYUdfI01LzoxXAzdeBTMMixM33PDeGv56bT2x
ZtG6pp6U8WOIBnilRtrG5Tsup2/+q4aY9ImXwVrGBzNmGR206w7xx7gVEQVy+Myt
pPABmVMAIlo3LAwWoUKuWCEWmmiPdfXCO/2dby9NCnOuFEGuoGVluTH5aNTL9vQI
fK93Mw5ORxHlPhwtXWfYPK9GWt+fY/y/5wP1SH1y7neNayGxlCE9T6sG923iwjty
sDdqMznrpcdVbgnenQZ8ZWoP2FvMa7zXtJ470nrqNmao/X1zJuh/Dfj75Wn8v8Bd
7zvNWusW/Wm1LBYi29iPjC/I8OlbOpiiz5JsiGQ6XQHTK7l3pumn+mDb5S4GSqHe
FMetawK5LS5jx08Eha7ud04/C7enBsUE5d/D27SfoLeq4hFznUHXK+4cUmnGrHo+
pps8+fmkFP4nF07wvE+mY5v6uQZzEFetIcOpnHkAs21pSw2LxO3D1R73+BTBWSu8
nmTPK8PZdgza4sm/MUIUyqi65LIjsAfs6au+hD/aA9emOmZy3PQkVpUqyXdqe4yY
079Q4WYtqRTRPmT2p1wtxd1gzGla3FC/0rcmAXfKtQtUbDQLfcdvG+vcGE8PWSxv
HH9C3eLeDxs/PE15fl0Y3kNQxJyv7InIrJgmaaUOf+nUFLUpkrwlT3+xxkkhI4PX
5+t8SxctSvD9AXQamkzrAJX1My/ARBYv7mHaOb5Opa7w3HEAbFEtp/EShzPcmnQY
EnesNkzXT9SK3kvlYhsQ/LlfxDufeABvDC9MlHNFz87jXZ07J0foU1555jboKQ8b
yo2rsWXeoP6dey8pJTngt+yRdekTo3PU6QsLhXLaZYuxk7ymNQk8DyaSie+ieolM
hfGTqvwZqJcSKDiwgMHbEhkZhmk95PA8KLsOuyIAzmr9n/xyXquGLjJmz1k2vmFx
f94C+UZoMuGu6hTvhEjGxqfI3UsDUreRj8lo8g616rQTH1favBlizxPSFAkgugHY
8iuNOrxTFkefBS2mFes5CC3luw2xjUW+zslK7EHDgRbitgNIgVhL646AhbXaHC0Z
Ph+QkY2j4BMjIfIzEHno44B7PvEJYutMh8SxtPSULXNSJzqa+DCHcuELrDZwp/xA
hA3buNtqiC1bAuqqY2GWPPEWFSfuoojZK0u4KLg1CHCJPfVF33n4HSnZkafjVYQB
dhLO4yOxeWDsYVdOmlQVHZGFKB9W00b2I7ToOzUxBqUbfE/NyeeVZFniEGP8c9VT
FDsWpfd0PfrinEyB0AM8Sa6yVpZjd/dRTBKanucsgiKnRgbsZDk/UivLkARWcZ/0
shRevKFm6aKocv5s+xmEd2bmOjNSeZQcB0AYfzdfmOsZ4GxSVfK3KCpK8ek4y+/7
H+LFeGJsMpCcZ3xR29JrjgngSpuO8dw+2wskkiENOf0Bjx1EHq/mzFczD6IU5Idl
HlMgOQy5gfUpOBelU2YCv9uhXdVWpmCX17Swa9a/H9VpwvxeiSu2uyvoKeA8zR1L
8+kqygMZw1K2Hsk5zLSWLGZvNyks9Cw+1oEBcU90JRS/3Xr3tEModwazMEhs+hPD
mudJKL1dk5hMA3V6ZkxfLMBNFBe9mp8cZVf5Z9RzCcF5fhq+3WWz4/L9rlVaarRd
8FzcowWqT4DkMXq/0qRviWDkH3nQYw1/EIfLQTOFoJtYvXt683WevEjvnHxAvyDX
S5Pz4rA3/+gqTsVLfaWpOmgMmDwT9WL1EQXJliHK/duAcycS3Evx9iaIWHvrVNVm
UtVtm3rHsVIlJn9vtwaCubQ2CwzQoStenU0k4Dn/0z6lR6/SmNDs02rSfjV7GP9K
EsTCGZDMvCX0XmIB9jRwgelFAEB4f+pdWf4e3rSGO2weudEzXeSCiarA33C0NLm6
5+L+l78z4PhXhPTdr77Fp7ygIcQrE0BTpU59qOR/Gfwg8AjY/zmDuDu+5X7VsNAU
tuqrTvXC1LGV8FC6vxYxHMUIGkZKKpnvYG/dV6tlO8zrHo2LKk7RIZLcKti+OvO1
n1E2zqTrdFyDE+JpWOTSDYOFHEMp3oDe+IyUySwIaPiQsn7//rRfs58LqNIMev5r
y+8mG9oNI+yT+P8vNOJlAOsog3IAhW22yuIiEhVBBx/i9t4c7YzNYKqtay+orOe+
H+R6/Bn09PKYmS5TbEqsD5Xvh7C2TcqpaGb7zqtw+pRgjCwsREDOmeSgax74ZSIU
xSpbX6WOrlvfNzpno9GX//8usUdq0dGGgM/ycCy8rww8RUTsVgmWPSQWjxz1f9kP
n1hk0+fDNMb/PT4t4fycsFN5IzOByFrcAlNIDCqoQd2OtTJARV4hIGyDbFCXylrK
/lPS/F4EsIHtll2UhilrSE38GPXp+jAS+UaZaNa4x6HspBgW8qF5igMfEtLC4Aoz
4aTiisI9gNXc+CiA33y6AD5zxbXFaej3nrGMgzGcE91+BPI7IoTGOx81qbPW7iL8
7UeiUst3sFIfWXlW8XIQ0MjnG9RYQ7BY1MQHWpIzDCOMu+5fu0pxLHxIeqr0C/r7
QSIvp09Epfs7OjR5lM7WAJrZHBzGmXtOBei3NYVwJnZe0ddU/pSeujrwEAAg3OQv
EIsgCSZEoTa0SNO5zenKAVlwmFWXeYYbNeXK96JOr4LRbABb0hBVpzuVrGbOTyZa
xQLKgpENBs7bg0c327wN2sNj0TUt0Buc7TA6n3i8xWYLe1UmawXj7YQQLw+G8dWz
TGMzzL/SdLSriXH+uPGbxeUs0DKZaHeMUSxiXN8G+kUtsjxyZnKFfB47cvu1BE25
PaDuF3fK0yVTJAitvK15bUYnOlcUsQzLS2D2r3t/AkI0vtYrLB97cIDPPTTEMhap
sAGKdj2OBZelRapZ+UjGKm9WPbWtggQgKuhFIfx4ZO/R166Q+oXvzUQtys9Vplbd
RDC/3ubVmY4iSb79Fae1WkWlkweFkX02LJY96GAZQqUs0i/RE5QW0YHrhFvOKSLe
mOo07e9g+63uEzZDDBV0dj5U6EPoCo3KyoE/SwXDqOdybvOOl0B62zti5MS2J5+Z
zMOliI6sTW3ugzlVn6+H/UICtZO1TcfMeBOxDZ4iPaiZkg874jKvuQJeAb2cQTyg
1xDv2MEAZ5kmUN1kJPSws/b4cBmCw0Q8njQv/plCLUs7irjWukK/RMbNdie+UkFc
T4+NE86WKm3YslnvpeMYDRCicbVIh9SNuNTclGbfaermFlxF7yGmSDylJDiG+xYB
DCgDWRVguGtrW6eyKpgeQ5uUAOiI+sIpYnpsZgJdJbwfL0lCwxKOMMcVMg86c9ql
6iwqa84VZG731spf8ocBMw6ZETw2VAxfO7E5639W8C1ArraDCGhBIv6IAzt4G2WI
W9TNAPtyYMxSbgGT5TZSAJSW0FrTnQa6o1hBULlI4mVANjqY53F+pfKsQ8zzaHoJ
bbUJSnjmMHdSNiaU8dKBbpi8M9Vovoi15bEPgPkoB3ff0LRPZpRUV/f8EquVLKkf
zWmVE6hmKFubLv34DYzHWLTyyq/M4dpxISBUj1wjzdC31eeFwSfDLLD+wsG4mBjj
HA/f5KIn+ZrKLfJ75jdkxoH+1CGwsQpWub28mnUu/fydEEZBSkB7UOeiNQb5eFhB
pAIM9Km6CtEEnRgiFpyFB5uSdFvDe1zvc4Ki45m5WHKNKF2vL6aTtLsHlO+1ZJwD
cAJ7P8+nJXeujJMC+RIX9LY4TdmOdiUhyzszWxxtBuKVScSH1BaFGTGZcqf142yK
h23X8F4mIewf1tekLjqTWs3Sz238qlyAFYhfBzD9OpPa5VpWreoYGJz7sTeJoeWn
v2Ybyk+zjQepScKOiYOdMUkyhVbwDcn7v0H3XIlP+5dMEvd0NzsX+TNBN1MKP7GV
D+XWio1rXdPmA580MKHoZT3wUP1c+ycfwyz0ReswPF2Z6kLVEiZo2LjnEYb0lLGh
ZbiK7nH7vur1SwHihbM3j0XkaklRpIgiV1xZFEP2akEuHpZWp8vC6cQPGTpmPpbK
aDkqqELaaUEy9mGIIEUQJXiMvCxOeUopYDyUwVFXtt8YmSdrRLdDzAU9SKo+ab6y
vrjSnt6P8wZV1GnEbb3kfJbqgjNiIK0vy3bURuPLN1JqA0Z3jt+mPjauuU00sg2E
GQdBSMDeL0bq49EdofeCZlT978pXLjX4pkzDY/pEOvw6XhRRL/Y719qbd84p46eo
wn0nCieZLXRtkyZ52VPTn7O4lOfBE+umsZpiX71R9+wKtGyq/JHbqUKBk0zA7XZG
Vkh/EcJA3uI8khFc9wM9iZyhfYVXh/wfY7Hf01jfA5gLC2ciKUxu8zCTnYEuwkcs
HhZGxYORuWqQ1fhHHcgER/4nNe0w20RAFM9R+OGrNEXJFO7RDClX4enNbOq5cvuZ
+ePY0E05XAXY7aAwK0zMUF03gZLZi1ZrH5B5l8WeYHYKlpKJSENynZ51X4gIj1Z6
LJloZHmfivRltxs7lgJ5BMcLfNu5+YNWD7/4KVng91rTZkI9A5VTQvc3R2PlZF6i
J4spm09xIPIv7Ng3vix0ufiQKmNtjBUGYVBAwuVfAdGBTaiDwPqE5Wx0MHULgrbX
ADi7T7nKmVgDs3sLsy/09S/TzvkQvOiWx16NEDfbQ4k0BWXQN2ny/Yko55aWIFld
keXB0mvo7VKjWrYDX5K6o0fWv6ZTbSLrZbbdpzr3FvzzM/d3fFA2lG5wuGvSlFbp
3Hqk5onijXlu9NzCNkfdExwMm05gJ0iJODh1LPFrVJTNIJJ+NbcHvaEuWHbvYNBT
T0mVcx6NVmqlldN/Ih6vOMSEyCes1DO5ZZNOLwXaN1lqE0XLzTrzHTXhZ3fMbk9W
BIbyx98UDUhPg4fV81DYoA2SfGwTU148QjYrcz8A/P2DV1wr+Alg7andk3WNWv6v
Hjt0awEXr5vgeLtepmeZQ8i6B41Ywlf9gwDKh8/4r2gNkqWpltVaLBVf5RzohKn9
7vt9KsTljbvCRxFvNNNZLHlRKIaBgz7Y52aIojL5L9ut1fPzpTKHFaAwiF2UCDxD
hvo+ZJiN6K6VsVPQXzJKBPtxxfui64TmoMzwkWb9nVjF2hF/uYl2e9pC2iUZYCH/
NPfxGlXAhsoe16RKiP9aZoA8aXO0Yv2LniGRLlJh/LZjZoEEDlSxUhP5YJQEwB+f
OqRofjlgKr99cz3y8AiAIg7m6jtjEJ9YwbyCYlSg6s1CPavGW7Ry3dd9K2wNFCGw
Vsl8kefZ5mkbk5G1U5BI+SQ0sP+xUaDasqnwmelu27nMSQhUANrKYM+kW3jMt+HL
OmL+Ycwm3d64T58R6VR0Zb8OlxsmeC8spxOi7ItfX75Fepxf0WzJ63P5IBVfYJ4x
VhTQn9W+uZ1TywtKTYCRzA4YeB4j7QnagSrg9kZJdbOuAtyGDzfoEIsSjM4JU/Mk
2fv/wtAv3dEYcSRXhftvhblHPTVjudGvhU90ssn3RmWvfVZWA6d1R3a19AVdpc/m
trJo79jXR2cQwrtCdqbkcBx6t3dxBBA/aoLU8rB/JzDABxBXVsVDO6S2V4u1G5dN
5lDvOMmD7zDWwu4jTVNKEZyryk8oLivOUCxgg9HrqQ7JTLktKr48kNLgkDjR1Wrn
3ZGQ9KWwbFE5ZnVYGYwDfUaC137yVWgtTIwCozQruFBNCHtvUdAKVtzCf6gWLuL7
cXuB+MqXuYCP+thPWVjwcqp/xGVT6R5bs1NCFVKyLrmorJ7Qcj7As74T6M/M2c91
syghxs2fU2sCyze0ttJ8r83FLlVkHCvmLrZU2uxDLaFjtIi+aX13JDj22sPiE38y
fRvcIOn6uXOanYW8/TRQuAOMwf2oIyQ1j0C6DH/IfR1qPs1E843NDqChynpRGwJf
rqRSCS126B3syc84p5GKmVGlrSFJyrYAmV616WPdqCI87HBYtn536OOJK3ageEd9
cZC8p8BShvJbuml6uls8Ht6L/gPvIkD4SQ/H18Q0ASp3rs/g3+5v2pXUlZ0s3/4u
mRTEwnzmERtKvl9m7wkDpZPS1KfLsSE54FTrYzWPD6LOacFsT8zZ3JmfKOGJhr+P
2mUPWdxXJHbUvY3xjp2NQ84Y/uNEhDvbCCUMc7uRmV/KMTMxR0sG/FpO7O3ecVdx
FlYBwos38V7jwGNVEMurc+X2Df+SQtAWD5I6FpP3mNihi3yy4pjU4f/A3+hkrRmH
noye1LldkJdTAUmwbLi3K0B0gZVWST2BJAIEnf+VoxkMK90ocdk1ctUgRfwkVUj7
Wxqob65huoDA+SqldjU5iX6Mxp4ccHt7Bej3out7CaXFm74SDPltdOZ8t4HXhx0m
7zJxK4vJEQS6JnSCubFvytEYdj4gFeso/E7QDbzrMgR8wMkec026lL/w2k4g6MG7
5pXTrimriIu9pSlNlTOakUAnme5dxc8gaNOxNhUMK7CECY5ctj2LVPumJSDrc6L4
0+Zad1tWiOrnqkLUXHS+YgjWx1tpK6wpOijinkyauT/cdA6ZzLFmUaTsyAYvRudk
rMz9ilhgLWk3JpT9rsiiBYoy4xfN+Y/KJbRfcKHhvY94pxSUgl2Ye25zGZCsPaQI
hfkErHyBs2HpT4Tc6k46pJFN+w6MYyxmLO1OvjyrdSg+IkqTZwui0M1qLMAb5RmJ
4WVZG+WCPbKIKjlBV/+N4iTiL7I8Q7nmuhfQmmOhThRkGE0RCgBQW393zw2wpNwX
KlLoTKd/xkKtT8xBt16Gcelso5J5MUv91/8A+UbU+leR8TKFXsOBOtUfOv/Jt0T7
1Ucuyx0zS01wT+YYr+eYwywT+SM3VZvwNwlDnxulhHBOfxCFoJ4QQZkZMSexmVfD
r86Y/EmmGNtBDHQp904U6CyTAXh/YGa3x9pvrR5lygOgPOgnulNp2IhI/OubOAJu
efoEDYU2k11fZZbQlZgA8WPGqFeAWNp3yg4IUhBZfoBTl2R1/0AURqQ7/DZEvyfs
rA4KIt9nlDLqfcCJzBo+IcXlh1WZB8ZBQOsTMaM9nZv4AcUqbBrnwNnCrnF4XQgZ
+VetCipIqjxgjXMTLZwfhHzo1E6zV2yLm7+NbzGQd5ZWcslfvDUQKZE/ECR4t+u9
tb/2Lqc4aTIstF4s5LsOG5vTtfgJaeSxWJG2iSIDwqR0WqSo/JLvMqU2vwbVCQRT
pYUKLKw7cF5bOcCDIVyvtYIJsv5NmNRt8VqZB5SeZ4j8xD1oHCwAX/S2KJKE1l0H
m3UtoZYDF2/dDRwWrAYHQbpwlbidBH6StPnpk2C8NDHbFrpw+wqT3BKfP5QFG0MI
/rKARv0tT+wVs2XEY0LdHzgkFZM/5ZwBav1lPPUP29lVI3KF3Xg6GSq08lirgbur
Mh1ETfVdZi+b8WzuNzJAiCb6PCQCJy59oo+7pc72rRBPzlxeQJw7TVfkNuszudGB
TGMra0yuPz1lt1Q5aH4cxG8GGIqppVElnzojWLapUFsXBYRJHNixpOIL4+PeULHZ
iGQtwYpsgdgpjF+iW0XwR4uD1Y6v/01PIlm3aOePqM8TM0QQvuzLliOwqSs0GH4K
MHIJ6dE2PfcsdlL8Wr2IaXbHRMr5LqiQKmVhQgBNgDBIJor5lH5Ga8OcUVGKm3Cf
ku3qeD5j3UNLb62RNAcyyUT8bQnySO/Wb4OJQwXfORZqguadsuwQPrultwjKOdSb
xtdi3A7yCI55+gWNnjUKG68jagKuCsTgKeLt1CuYS5zfX16rrNTmxSUipodsJGoH
VAMZ1OrwA28es1wHMmBiCgGwKtsUfOg8Y2aRqZHPEiwCbdZ4gSTVLtQ5nj3RVE20
aXYaflXYstzAf4aFukNcVDWoJHSn9MP0nkczrkuNNajr0WtijCGxvQZEbMCrFRZL
gg0wGZArE7R73AHRIj3jDESTJVc4fPbcvS3p1m6gFN6yEIEEuC4DqJzchoOmq9gc
bvjcyv30c0YrojQ4/rIKQ0d/+Obfc6DO+2kljExdJodRD8TQ42JyEnmKbOGhKl+q
XEjb7wNJCfqmzaN+jml4xFR2y9R+XCKiHbtasgIS8WohQ6rf+/1ufWKaqLM2YPBO
tvlmjwfxNzczyieSFftk9sOTwL5N1qhZZfsRiVyyhzzgACe4/9guce7Gch8004FB
45wvprlhxXNoe3waKpl6QxUT7QgPUP29Bp/cEs/TEddeE9Gyws6jVtoPy1Nv5osL
Zk+0OXwj1A9CAMMB9KH9mpNP568xwh0eQuJSU14iADsPXHK/3SjhMXsgozcJVIMj
uOpRToK8evMxdQi79BtKABaRn8TTAmbn8O8CdF3ll1e1J/aVi04iBBpjFC5f9+Vg
AQiBM2X/kS0qLlXl5UXEVRh5qZQwlQ8bAZBRi0cOLbuZ46TsBnOQ8uq1iWCAzoqL
wb5hfb4xbwNV1a/Y3WKruEHvnGl3DRz4SrEDrKxwLtgEXqmU16QkKdh5nmWxqvup
xcG3AI8JAzxeTm0UxjUqYFQCVPsMBTD9YL9y/ORBN7XLEEAbbBFGwzMuUwrbcO0h
LGH2Dd6lvkBj5JKsIOsXU59nszQBXfsrwlakHAwYc6fxNJrxakrtLL3DklmBfhSo
bRGwvcheiIZUAt6eJjDAw2nKl92gGGGkWuWlaEtFs4eVIxC00xiGpcFYcbj/FXUF
//Y9WF4wD64aug7paERo53xoVF0nz2kkDytlhgVqfHhj3lmgUhRXEM0+PGVzbkIH
+xl9/PGz5uRy0HPJXQVDQy9LbtepG3QLcQxQU3cvruFOptUjUOEd28bM0tcVRGL5
KZ4pHRTIb6QYh5lqXovN3d90RdyRyqUkv9OQWP/Npk1szNoG/Wu85e0cydhmL7qq
CHLBh7/bjOQ/3crm+Mt+wQTt3wNYC1RjgKuQw7GNHloU084FPpBJKUUPg+hyTOSM
xPLMilgUeTiOs7Fh1yIYEIBoAc0Ndyb28hclFMEGpFiLExx5JIs+V2r+rln31Utz
N+q2FYzAKwalITPINfiZWv3Wp93IHWTkYDp/G9N9ix8MfzgblKz1euIubVBgltwS
ywGHUHdLFvoGlle2fnVx09fpzXC6s9Flam/9WlU0bYnmdyueaHrn6SxUilJNgGaa
K78yf21lrT5Aan/MDoye/mXE3JFB3FmFNbmJcW4J11KVkrCE/8Dpbrny3a2jZPfL
GR2LsFbilt7vJmLNNyVAlatQhxzy95UwXdp+LOIjIbBL/x51og+2uAY7uRyoiSah
C3KKzYJCn4fYcdT6+Vmp0MJMeL4knTnIu9nyDQQ5mvRdsCNFTvo3vB40wbr7jvrI
iqCLKdCXQuKAYsMIyFmUjg/3kKj1GGlTB+8zIqPalDbuXqL+0pdkfQ4MP/Kpzg4I
K7rBtO8EWk+ojRwJSb9EnVzliU25741/cEUE5Pd1cP3WumKD9aHloHAr1YbAXgLp
XX/iS/38wjmtfWiud4NqrWw7bdpMuz2CKPGdsN+Kj6PxHA6U4waH2gwbvVy95xTs
oPgszai4PHC2qIYTgq/IZTBfHWute4ZEex3d6DULOVWQXPnSN1ZdB3tuAf3JFXqE
SptmBou5uJAkywC8NDfofesyKx523OM5b2PZAwqUS9u/DMcbeCG2G7b7ZHNSiaD1
CtGLQEHRm1rxx7qnIPxopmICS2ojjTFK4bc4C757sKR83otMnAFzRuDtzLzGE1/Z
biEMs7C2GO4SQ0GY476A0ynR9Z6n0DdUCjH2s8XH4VDPA9blOzC7nd5fIJe+rzLH
QNrbDpxLr6OG2n9vLQvERyXBEGNUvjtCCukH7U86HHNwqjicRo3hu2vIFeDlG3RC
PiAe8lOEmKtrXqu66o5OZuZqrHNO7mR3TnVo7go8f4BPIKphuR3sa6VVKgXNlUle
4bGJ/8O7xt5pAegbTIndz/IsE9GFD3BoIfnAmZBT3+h9SNtkRUy63KPGLAx1wOpJ
BRjrsDJitXsD+GZCUjVGzxiRCdvyFAUsFbQXuqdcbu6/WPCYP/8rx9bhuPUGsLIz
QIKh2YS/+wcSxbqtj3C5C4bxwNJxy5sg6DloNWJgrnANONHkYFEuFdV+Dt6LAqPQ
radjccxDdbzBk0I8AgUxwuFC9EjKxhk0/NFvlfwT4GJEkmwun2TB9sQPcf//6L7c
vpY7lerDD6MTkTo/3AclDGKD5iYXVel5oewUXEqaMbQUeZdjTH6Nu8zQF55ToBtX
Iyq77R6ANIna4YOyTj0tjQayDkWfnU33yTT4hY1h9G4BTpNykV4nPdOdIQblnvtc
6Srk0W7ZkPNIIuzwccLs2q8Imi3omlIQCt4hi80ft+Gxtwix/ypm/192hNfnp8aK
MxgfI5nPUiM0VbejQ0LmkZ/DAXgRbKMRnrFKfZ2ztD9BmiyyMWTG0C2j3JYxfBNz
4zLlxt64cLmy3Vb1M3dAQUqSpDMgwN9MC+aU7X6J5+bmI/m9QC/yXtvipBxnMmX6
VGRSD7PrLzjS4z89e8OT54piZ+bP13eUCgMGWPqD1wUBdTfyXa9PPVfc+TmPjdih
SoI7tAXPec9NNfw6mG5123LYH/Z002P0CHuVhE992o3pL7Oag8RZ1v5QDq8l4Q1j
WU5/Nm1pIwXh1oYH7sG1gP2SXkeOdS+uBEpTWwSuJlk7WiDo5JWx3eTx2g834Tiz
7Yj9UTiGftT6NL8N8n6uPZVZTX4gBaklcKLpnIpfR1h8AGxPSXe0bcE7xgHsJPOQ
7CY4uTHH9m7dCF1cgmRKq23YNAnX0XktnWs7Jtbnsgp/k8a0aAcpcAuvprWBMVVR
VjmwlLS6CMlepyRMmuDzuAoXShAjQvXgPvruY41TdwNrXtWan4zhn4NhmAtE3hYh
aYv734C9IFNsj7bJRcWfl2PAdHzGNm5isEOEqUeQ2y9HKm6BGzv4vRUorxDjEgh0
zPZfXuNp3UrT2195PKeN6vPFpO8EH/wP2eK+QKfaRUWzCzjI0RA10JvpD+xEkR71
D16jk+mSh2xdo5+8K+Zc0AT309LoHz/+1yLqVb3nbe6E84z52vgZSP4xzXZr0zPr
A7WI971rQ6YMLCzhDWCwUUFgmAnpGm8bDRWIivZ+2Z1JGfrLlNhfDy/FaFwz6793
NBv7qjd6aB+jEaOLM4ojLesOYZXVruYbEK7zFNWhOmTtcWycCMMSlea+0/WIlmN3
5dlAWUXd1mxXdier/57vRf8SHTpl8mFdEKq97PqHMKaMkTgKtjPDl9DTNZxceTL9
9cZOxTzPrPKvsqMNV8TV0j0N/McSljnHZTvbKoHEMyEN7xgEYfuD5eZBkVVnv82Z
tRUXzcs4wsOedsDX6qFlwrZc9T5B7ILZGJZNfxK1m4zWtlxLhKXaBtnWuXgw2LRa
d59FKA1oXLNMsf9hNIaRe/sF4+ZNXwKC1INKWkZYbbPtZGtohaQMTx/fNkWT+3Si
vWRcT128ybn/TdvuUSEtsk6oymXYzumzFxpeE9tUuk22zI3EZKHF050WaSdMF87e
qqYKdAklEGtE9nJG/mX/9qbPAqGN5+ScIdRDqqu/HXWaUDhWAbeGw6weElyV0vuK
fqdhJYms7ZgBpA3jCqFgSCvd37lJkd6rO3i97WNGy9GMxIHMIhnqRyQHpE/UWPwC
KOUaePGe7tHTiNV/8gTpuiNJfljS+TZwMDmNGYDQUEkP+aXv2O4RCOQxAsZHOVw7
HZtDjALnrlGHNkVFOvm99bQ8LcC1CUgQtX4agq6Dn6CfSEaSIXQp1GnO720IZU+j
/M6UeowGPQJPGGYT8A9BxUIqoalcuGdPiIWT876wVY/ZkEhJUQvG0gCWwt5Y4wgC
8qNxaAfAxnMcbDEnLwSX7vNu7l1+k+15wDOpxokAlQzSQeW318YhrLLBg2E2FS2X
R7evNNnYmT1rQOCwZN2ngkk8wKJnMVO0afHK74fqgeDV9evkrU0dwITqscdZMN81
EN/eKsI9hOHnELh89YZk946tJCC5VfSpEbleKqrHzg3v0l+S9T9S3GCsL8fvB1rL
vBQS+pB6KAazYDu/iA9K3XlxRnUWipgL6bCCHxOVy6iRq4Le+c+ktgNclKsc5E7J
DKHcIhHw+PH38OSULcED7TyLnMP0aukr/I20ZPjSo8YIhCcIgqWaZDqvtZbvFXH0
S+6/xoHcyq4X70uIMieqqEPxAlUHCVkaer1RM/83epBV4HKJZfrcm2z3/Da0rron
JB/Pe+RfItl0mzac+eaxuF2CCWd6nIMVipbJcc3whADeRCacqgEf+t+CBCQhc5TM
JyE8+C1RRHc5X1OUvTaBgFo09/2lnzoitkdzW8+GgMG256MYOcP3hurx0Npy3msE
kbOCT/dqSlNS5fr8D1IzY7z7OYY5bswdw9OHPqk6Maa2KFYjAIz/krFNYMVELaF3
5MSE/qMCYsKCrIeUwMeqdL+tw9Ycsksq3FVGE+UCS6u+Bhuw0otzse8hn9lN6rvQ
d8jqanEeL0+Jixxlm8JMp8qqS+nApEFSbiHIE80HPt+jvFMUwemq1G8IfCP+LsdL
VNMuuZez8t/kAFbBdmGhANMLODp+TMO3Rwz7ocftkPVoPVsdnttu2d2K4kF0TCBi
/KSNj+XvBBPWMrgpTlN+iNq1QNDWbi77yZ+jzbcKtYj228eu8UFc3CvAcNgySP5/
r34VKB6sSLkFeaW/G9BD213IjDFrrq/iboMVlLO5jM5DdjtZeB8D91DcK6QlUCCI
vIXMY32BrQZYZKj5DWYTtGBord3XEmakQUly8+NjynS5I/NvEkgSWulNhqSBW+pb
yYlsac0sQeGh1ntalvcqNVqBCpswqJEDWAsNNNUZAvG6Z3qyMRlX1f3BRUg6eOxs
mCXw3EGegyDqDrW0CvpSv9KLl0LcxRkEqy3Lak90/J//9UFT9+gInsgV6woK35Ez
hktIs9PyfebPjviMObbSdD3jSzshtsFfbx4kdtsQBxA1zbWMhXpyYIkomdWIi6tu
BUY6MRxStSZgI0yL0DlM1gtIz/BoakRe/HupyVglmMzW6g0ZPGtFOp79fhrQHGBy
7PDQnsFgXsH2C1oQfkiJh6ZAWLHdk8VAXG2jFGfxCswYT/or94xtZft7V93j2OtU
6e/+tD7EsSwuQHBoTQm2tZ4/e5yRDw7j7rrRp2gMAZjrw4aodEGQ069hLMWeFFmi
QISqIvv/PWNIFmXhlFTGtd5q/eRY8Siu7ibpTVbsiT4VdVvnQAQF21OOraz7pbZB
16vL2VCfTokS8fN2soHt87s0HXXufZ4uXVLzLdIGIucCkWk5s+pN7Ur3aVhvsn+x
W0Iqbq2Ci8hL2Le5n+ZvyephRtts6Qc27/B8vClPInWtbBIUNdRIfa857OxClWdm
I3JJ1wX9zpPhCTsEhoQwz3/WZXnEGk6mREL6aGD5ditqe95w7isgMFyg4YYTUBGQ
sEGEg4Tb9nGFAE2kx4hSo/P9GHCtkS3xJt49NdUwnwcqFd/dOdP0tWQM5HWvwq0a
3772yMt1ScqUugZUgKEfR0NFuKKnuLFP3Wq27QmrfkxLPAuPJbkUujlN6Kt5Y0xa
B9R8IqQqVUG6UolVNvClmjce9vA1an/iQdF5yNby3sGIKduktHZMlcEB/aFq40fO
v83n4ahis3E1zbgWSQgjWzrFot5a2M8WrKbiB09N2RfuP0nS7nZwEOH93Wc7CMZU
JDv51764uGcCjUPRqWUCT9/Fpc+3ntUcmIzMKDZIaYruNbq9XLomFhwI8fWd30dY
IMbvME1beY51KoiaVy7KVkjPuu2Yky3vGyYtfEbSCO26R2LhP6BEvjOB4kB6BC4W
buQrRWV/nCcZdvLrXeWokGR4XRH8h4QK4epjRJg3yQWuYDTtea7spoGUryfxFrgt
GdHddzszH3+Avks2kSuNiagyn4jpcRzrKW74ZVu4ae69gwee2dXoOnU6QKnbHbjp
4fBVdIJe73IE8i2jVmMjhW0gFCVzI+yYjrroEoo/gjZAqzJMFL5XS6zu5rqvMqAk
wxVH8JFCt8rtfn9AsO0VBD1al4XgSrPPqhtZUIRp4vog+YCjdaFg/EURXoTWwaqa
mLErmOGUP4YsurdG6J1hZiKhEQjtLGpXjRqNzQCDxb7b5Z9693c4IFMMKMCzzVQQ
4UdlqVZ4e462r9vGTNrA8KPdGgYqAFtQs4SPLjsIwd2iZAC2KDyEF74tK187ytj8
8+u/41H5ZW9t82MWqcMEnNCwtFLfdxYMHzVOqKbvbEQ1D8nwu4y1wH0rxvgxuk12
e30TdPtS4qlUL27crUTAfyEA9ILYU5mX0R4ZI5K0o1poY6ztpQdj5dsi4Qk9u4Ro
lfYuwHKXIlUG3tcJpkzhIRKWq8z+j/48I6sApEDqQPsWbh6K3D7yoPoQUJupRn6v
AVcfnzG0KLiiY239UEVvDBZVM9W3cYDaLtCph5kJ6yo93aKWeQo1ax2lXawVcF2Z
fjlpVzuLmWLrz+cmQm/83JSu9PA1MfZ8DCkVt7VAXC7qunFmI6U2BYgpPBNj5pjU
vQ7LoM4OPdMkUTOnDDx+cncRXPZ0+ioM09Boax+B5tkGrKTsqf9iVFflRznXYCua
1Iu6MLzZc6iV2Qrhdih70awMRFz9oY7TCENgomOw/rYnZamk5vC/6aWhk8bQICN4
qoSNWdeT4gKsdl0ASaBQtWjE8WOWFx+W1ulBy4VbuzJRvGJ0TL8Q5d5i+rm6FUAi
0Bvr+SS308HcU8zPIw1ETZv2kmaAb0ViL6zc0/x+rd3pNhvODWSDav0cTwYQtac5
W1lvOR5a440q1xVZss6K2760xw0BB1vbvOyK3STsWM1LaKstxY5bxxg/3jNA8Nio
rM8swnJREQPzEmDsyPkOnSZbCrOCMSdEwWHcQNCWVGeIIX3BSQ1XldIcnNPz2BZT
MpZSokV/T/A4GThatgBTuEMOz5IYJCWReUqeUX81F1t6phhCqGuquJN7uR2eW0On
u09MJifFdKo54xv1+PNevxcMayJwt7srCyhFgPhvd8OpxCuHDdYH9bkS83Rbb6vk
BcjB23F1teV5gOXiaUKk1UABsC860q9LUHKUpA42IjcBrkCOaAlFjey9bzEfX3pR
8sFmaTMold8PkbWjtS7SjGIXqAZMC1Fjqrkh8PHQWubFWn8j9kevo2kIgK7p9uhh
vvxuMVrvViFtH8wDolAMENADAD9a+5j76YOXFmaIcabw1zAfBv3rrnwD4q3R90fz
B8My2X9omswFSO6B22sW+n1qOQ6gyVTId7tf4bboB6mY2Bb0IadZClAC8j++z7Ph
NZo/5Buvr6+0DApz8/0X5I92wGCrmbTQPwBCwujj86PZjcd1Jya7kaxIcfmx7nkU
2+bk1Kna6dhr4eJ7D5NlPkyQ2ODHx2pLx9NjtXULJSW97TNkiiz7UrcE4I4Zbtul
5srHDDqUCsoZT7CyPu0v6gZDfff8B5l9FRYv+cyWciuL6TE7RPPfLPjAENTh21bC
MiUDpHmfd+AW0fn4IsTP2wo01kk+ZJGUDTrTGrRBDMi5yVTAqV5Vjl9VfgJ+8obU
8Z+//3Bk5ARZaReydkaZd3nFjxe7Nm+XqkW3aoX4tn5sP4HdfraMEtVDvd/ijcbc
m6OaFc0F0upIi2QdpPUqsRbf/WhX8vsjSSG4k6Tyc7KC5IdoZDyxQ7A/ocB4IynG
lROieeveeYpf6ftiIEO2fHUjP636Eoe66VpPcXIFk009J3KkhHoVEHPtSVwKJM0S
kFZZD0VeeyDEUdyJ0AOKZs0g+89nYbHKs2Ad8RYL5DnAEzSsE92dXQHG0cR/AVh6
QGr/0b1TQoCV19moEN05Fy72YrwJIDBTyMZAYiNoDLu6DSv1ZnbunGJ8Sg2qIh0U
l/EacY6ELaZk9QtEs7wALfcJ2S779SU9phpasRjuXI8ej5pMVJONJBFzjr0sIbQV
A/gtxUbRy6b71XN51GBVDzUOOnybJRRxIUfL6UjlRjCBguvLAc50eVpF37pjUbdE
xvbE6YYsif22c6U1rh/ZuQRxGqiD2ttj9b5GZHpu/JoMS+BToKrFGKx0xRezCNj5
7R4TQFyppnl4nSs/w2L205MqKzbBHf1jX1eaTXebY/PzIueDc7bvgoKp/QJpAeC5
d1fwZRymGgPwsYQplrMS44b3xstE7UKypBoJYfADNYq1YD0mA+j7vkKhNjYD4h63
+2+xt7akTEvgPH8evpULkkTe9v0vhnXLXTM3178xlwq7d/SgCvYks5h0wnP48kT1
BN/owijoK0EINEJHk+MKeFGtRaUTmJBOttcrA0lC6Ic7mxNjvbH7lWLeFiutoCqd
5ttiW2l+RyvzI3k0sPEblfvhvPu3jCM4HH7228KfYa+Z+NPP2fc0v+R42R5dZmXs
t3Cgm5Nw+d3Mi7u5TiP75IZdro8JDTYuuzXUPXBUZOehtDtfkISoIr5gkf1PFAPK
CQ+Np5YLoZ1K6NXWj8r376OTyXbIAXAS9sau6mDqOwY=
`protect END_PROTECTED
