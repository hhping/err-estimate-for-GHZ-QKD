`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgydY2WDVZKdthtO34dn16dSUPxHlbq7Hv7pO3oe4nh12+Kk9Y8H9CBNto25hC+t
C92xk1DFfkT16ZsDFQYOduQ2PSsv8OtZLP17rDk6ES240Y5TBOBmOUDfRVvTPhBu
2ihDnGl46wOVkGZj/55e7TpevSP6yfjdUd3hd/eqD+e51+A7SNEMlUvew9ob0pd4
HRVCJ4Cnxqw1ky6wI1im/EguRnc75zJzlVN/LORdYA2DtMQRKRJrgK0CDNcxX2xF
+oaFIrpgqmgQhW/pg7AqXOTCG+JJRTbulvf4KsCpKmAXfQeI7csVLMtK82bqgZK/
8KiAflWTwGDIZC+LKFyP93G8T/U3sKOvF5C3bXuBqDF7wkyL+ZGjb06/r0irKReX
sM9wCZME1N50B/z6QzutzDOFPrGYluA14R7aoFFpAxprfCcX6516GQUCJAiXIehZ
5V1vjY5VEDoMvyAowNRWI3Ab2jv7ypxnXeOWOqttETZM11nHiubU7vn0MLCmM8Lf
PIQRCcSOGXV5MnuU4J4hN/En8noMjTwVR1dX5fU4QYD3E43lAybhJvg2MU34ZT47
pBuEy/n/cE7DfthhGDx/DIi3bTNNyJhlkxKWyF4GCYKyLNLLp6AsyQpnYAfZTdBp
MRpOf3Wzxfuh4vA2MUARAQhwQ5SFhP6+SqyDPAVAAMxt/xo2SmHoXxQlBPS2dXHI
JRehXfyijptKW+TIuwpXBjeHKGFgYLPERFzNLFItJQJ1gglkTggQqaZydN786tja
pPV28h42BFBc43BhauEXzg8KNWctZTDlXCejL6V1W0mY4GGWkveG0OHHBmgsCzVf
CjHDA8wdorDF8hbfQNdDDij2fitBrgvmiwln1hHXQgBLlIhhdB9ezJaOmk+bT3Bf
VoYeYHY+50AH6n5uZaTv5rzVhuclbVu7bk6MTxl8LI1yOjUhHbGkrROHJU+YxD/s
I0jaG7zu5ZZxXh5ZvrLvF1uUOhlOkpSWIygzTAPgBicCxWtaIkH+XHkP6iawWQs+
gY/r8yzOYo51nI8vbsYBwC8YPHwBTAKiPvOMykX+ZC1w+MtoBzaGuWvzwa7yiz7a
0M6/DvEH6hKWa+HAbu/naLaI3Qcgjjy0bwB1DnsxKSNO1ZmYTgkzZAsBItrbDcJ3
vAAKKs2jz2Ihmo1LQkYhdpKDPQkyp9Xm+VOQFALrD80waABYd/8CluLkqUbU80oP
gOSJo2r4t0qp34eRriNMr0fcCBPeUe1yIpAAugoA9Z3cNhb1h6bF8W8qQjyzwsoc
kcEuMay3XZls+ki5HWnKVMs5CkyNDtabGU/7wKgONI1DMlfptVQ+K/VTJD7vzxHb
qR8sAOooQEnrOdJ29deypnJCiHmE3ZoliMt6cvopPb0F/JpACPImpoQFtN06DHR+
M4DgqsUzQXOkWx54kZ58wLjSqGC9IQxfKUSDV0pTnWhjzem+ff97bXf59d8Yx7nv
lHaXbTdhYZqB1yQk8/Puxi+Jwyh4XFrl1+QQkGfcb1yXqSLzScd77zmj9ObvcLaq
3bfBkPrC9Y4zeolrRcc+5adpeXu9tCqfv+NF/+3Lao3TjQTFdmmr8sAqY0XiqTQi
kjCGZbGCH+eLAOZMI3mVJ4R4YrIneHr4Mg6xQhv/+ZBObL3offN+le7/JRBQ5rq8
mG0+afgjOKlpOA4aTJ7kQKiDGHvDnjGmo015vR+N/xzN1ElNSIogLSnaM8lvzSAK
26uCsAW9s1c40rymy+Ah9oiiued/Lw+OioY3AAnXgU//qm+2/fERJGZXjXyTkmSD
ZV9HZe6Hmg9AnYPrNFlAqxafew8h4f5VbzGdK1zTo9vlyhh8WqcSJlAIXN6nbGgY
y9hj3Ela8Y9yrOuQrSzmyVGznle2GpIDr/nkBujmjh9tz7sBF7//rzGcAtZ3T9pq
UaEEG9wbRIrMpl8XTiz6fX3KRRIekYapLoOh9MhkUW7BIMwJpLwtAH9h9L81RfqH
`protect END_PROTECTED
