`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0YWmo1eurgdSuOg0TesWYi0yvc8N4JfqLsv9U/G0qsxukzdK0MXC8wk7JjlTa7cC
AnNrL0T0jjQ8aNP6EAf+F2wtYKtY87QzSbQ/BkKuJGwlZobTdDtmxkIQb0Pikt7a
hpoYrSM2N2gcyz21laSOc64BGCZqGB72TNT8LTVVY6gPjmCc3OUmpOuKMpn6C2jQ
DcG9JNkYFPtxpbMZTzrLru2Nr8xIkod7beYqNxJxUcXxNy8eT6Qz7/BJQAnQbwBG
AMeJgpt+RQuNS1CJbPBgh6ev/VNVWQ0Ha2YUM+q5MbWaADnXb5sGSuz2M5iMZWqX
B6Yx52DytbprzPQuvcLQULe/NnPrYHTSYd2PhOrwl5QP7UbMI/gp4u7kOaVzfIxP
G/AE2dHtQUWUOKKko5PtTyHfKJSHvXsXKE2wbDTR2XVhzDd5trfRGrKASb2xfyfM
b6LkGU4Hom7atqK4ACY0Fg0YUR+fViCJ5sPmapbSR7j9fI+MIbMD645TBn/pn/YS
NtKZzGDzrfdszwsdYuJlzSCAjhHAapo/XltTA420qMhmbHaEoVmSdohxbNYdS4Xo
rb34eZe8fmGPZ7Y9KDM8SqLZdYhVJQUdgdjPdxJsjpTYyAQ6mkheIyKJworeM145
k66K+hjn61vuXkMljb7EIuxE14jpe6lmCBM/Fy79CorgXQwFUIMK3CFACR+H5mEw
YJRqLBLtmCgDA/HH3wVqvt1UlOs3JmVujzkdJlfiXX4=
`protect END_PROTECTED
