`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Pt58cil2KKU/wbC4EV4i0mt7LJhIHf/nY+00ephbGW4ojrt/ii1jcuQHFk5WF9t
EClmdhmmJkrGfE0vvahRWpUzbrqrqItPEaCDssfvFWdneYqM/JhqvvChcZ3wWOF7
dlJI2sadd9pht8CF/LiFbF1wALXsFeZ6uUDk6OlizkheVx8JJICUjLiF58GSyE4C
rBlH1ksRjR65ZgDlzEyd4aNfgLICPeMFJRWEkZdyIfwVq64x8nGbFTDQdykaDNQe
QK++Sj2hnEMh7RvlJuM2CF9w+rnnyzo7GWoRtt1tdEmLBpz/+HmooeJQjTPkT98R
LRxirVenHO9WKLbBcI0Nj+hGeYNANxuQi93ik2Jp/hZkUgDrCIXLxn44HM94Cdp+
9rglPUwSsZ7W3tXwnPZiqIDyrImB5M9JCvB8SmXrMQ3Fo5e73AzTawTd/vvVkVHB
vbMAuzN+aIc8DhpdBwLRitmCAiAw+S96fTvdw/wrMmWZaUeo/SgKp04Rg4qEY183
9e99Xgmknql+yHV/lAyqNWUjA4SbxXlsK3mJSqwgZyEaXEbU0oPca8eIQhj3NraR
+Uvma1f5QCUYYv7gFsBLmzBLPvGXwFpYlHR2VjeCLrABTuwVeuV3dvRlv/9J/eMl
076DuKpNDFqHsy08X9AMLjw8dPfmMA1i/rNbx9D/hLNzQEpcUh4B8jIANFQd+Bii
OM2nuPTgvmda8hDOUcrf+HHSsL1348GnCdrWfU/lj1n7fFWCzLS6IwuoOEIf9RBf
3BTbGe0kg9Xuc4hgSWHiDsPFET5s2LxKihJ+d9OdRHrfEBYEJz6GxILXKzX7FhVs
nLsOERiHWpL3tbum7sTbOCvfWloQ7ODP2aJOSY/dYEYOQxZf2KstfF3TNdCoKjA1
0lMRH64b2O1qqqQLH5BXPPz2vEUkVQkvILcjn5TiQZhxPnkLjo2oje8z2KkliWvZ
Pa78UtUk1y322WbC2ffYs4O87ajXl+vFuLtpMKMWdjJqZsm3R9ihck44JZIJhc5s
b31FJXnM6s04Z7J+fxIC3yyAWEy+jL3DHJfs2OcMJeoEvno2vUeJNT8XXx+EWC6T
UKcfwyvAsYwujz/C+iub/Aolbw0K6IQv2aaVJtbHJV2sT3jRG2hrKoMJtfV//AQL
sWxii6tlRsdWY3h8TLPG7bCjzMK1g9N6czqA9YfVAt9JB4O4A+PXN+i9iHc1xGNm
haoaH6UbmvvgruJe28jS/41T2L/Zo7OUDM7Ni7uVhvDQXUl07wK7fvAJ2fU7zMjc
KtIFb3KTjmVTs8s70I/h0VMHvgEU+Uz+Mly32qGgCwSJ/A3DzmgiF1xNoas66eTo
cH3A+BeuGEP71axuSGm4er/wclRleOSzxbBlqyHRuoedLBvTJVUBtdAsOPDe8WIy
WzZ6nLKLVrE5uRwtH9FLGpxsukMVKol9HxP7W+em/WWuWs8C5XRbjDoro533Fc2s
r696vJ471Zc5U0/wYY/yDe360qXmS4opZIHsMI9h0i9sE2H84TBx3yLY+kc2Mr+L
SgRABizVVCoJKWKudxDTW18/pT/TbdZinZfajFzdKf/I8FmYw0/gY2u5i65GWuGz
YSGSkxIhSUorwjGjpIIIvms1oXtsQdj/ca8gZNNutxRz4D3hTr+H8pZTVc64fHFx
XyZbsKTPxTdw9X2irDxuMb/GWuBH5XvTV8wJ5QqXY8EpUHnYe4TOWu+ExPrRaUMr
gAtDDaViof1ns0rsjKlrXy1iXpkcz8+6Bebsc+VXkpUgBpGmkoAHR0pQbWEmGkHb
oV6yKiJyheZ/DmwzwaBVhFYRMPbr836QTghkycx33fuqdL+rj2JL4LfzfR2zV8Vc
GtFDRy2AWn8AAiPnaKy4oVhTYi+2JBob1vv7KEuITzis+p/8LRxNFPgO77AAKS97
hucgYYqkoMxl7Xj4AsmiZOilIgs3mVapQp1IRM3cWcTqJlg2D6z2nLCEr6+HEQdl
jZXq0UDne4BId0FBPl4O1zdHH8lg/nvTFtwrJDCtIyKlkuo6DW7wmteQBn22/mdd
ga50+7jzE4pEIvpFFKbWQW4kqrGgqazVlklZ12BQqZGkPZ9M2+aRRi9Nyp3lDxfC
1PpMO71MlNWUk6cGNda/Vxa7r8M2xPgZk3Dg2CfSoGkg7slrQvUCzi101yuPQ2Wr
Ax59alOV+KYh+yQfKJvNoHW/vNZkeeD6J59f3uQZ+mi1y6hVcwuX0XJ4dAo45VPb
o3+XGnKipN6txrztK4W/MqLwto57iAvdTAMSfeXgZj+QEp6BqTcIE5hclbM+SCZ3
5On9aNpyK34h4QvIu5mUERNmIzIsJ+oR2qrRSZSXblU73IQxxWJJkTFf8xCCRU+T
hqJRKXJeNk2uYd1vJWpyS3VUIgTCHx4uDe6QSQx2fUqJtGPahBicMqX1RVHR8Vdv
xhTzKv4AEkywqV6VoPT7oeSB2c+8JPPcrSySCOS0CrGUIJL6wwB64dmA4RlDWjYK
Ukrfku9+fBKw3L0qS7wh2CKsaRZAUohsMcpOh/umbUDyofwADFZSZ2sgVJ4JI2d3
YH6ZAXJrYtZQ9REWRzGJUzpH3s0pPfNlR8G8E6oK2wtIdrWhKlSrbzJ5bSHfZr+c
ZHiNDzcvGQZPeu6kvsTY+4VMIYycbUMiRhYiUs/O/4Dzcrg9ijN6ZBsNzc5BmWGy
WJmIH8wiSvCGGmUvVejkH/xyghSKxEuoimzS1cJxz77AVtzle+RKbu9UwfciJhx7
H3w77nDRYa84KasGkF9lSSVWqgh468oHpBqA0MVfytHsFHXrP5X1GGcG9fpFv8WK
/foRN04wcs3sG0/GB5UqeVaPb9YX8ZfMu31FYh1A++QuiQmq7FeP9y30MrZ1i7/l
6qZZWHck3j8bMO21BsOXglfkHqw4plRFzz96qPDQi/iDvtE6CBVcdw5rQAxybRYM
Vd58eqii05XE+j+mPfMRbE129ur4+YOmuzKxR71SKSVUy2l/evYXlA/V6xtHXdQC
Q71vgQ75SVucivvCdV8ZaNjAUjhx1To/MKROO2fsPzhGCBSCZshnv/EWBW5u1Px9
eGXQlRVAHvPL6Gamd0D/AdNBsPaF3GAb/H+RrGfGHDLW7wW+XV1hmFxh1B7lv5NP
Acr/+57wXMfvWp2TJ7ru34wkCbng4Rd+jMURG64CIpBrrbqA8v94GPRy1OULQ2kt
zrwitVSMSgQkZBh56hZ6cK+o/Ju9pXyY0qhhDKn52WVnXUaj9t1FbAsNWkDjvuMX
wRs4mWbDW+gl+tFDP1PkRO77rxM3a+wP/sskXGOACS3T80whxibNGlJSNsPugaku
XSV3NI2+OjGHff21+OEfz+kCwoLgbikJYOZWt+SSynVrP8ZDoJ2bVppfDsAdTm1+
bEC5jitkwQksKpRH/rcI4w8PlvKdL/J2LBQC1SdkToCw0xD1gCONkJH+WzK9Ip+E
FG1eyJ/uC3nlUhvxLj8JME6VfFhzeXCiC3djpeRqrErYJBn5pNSZjRxxr591Z3UV
/6x5k9ZjghNPrgD0mMI7lxVtZKeXzKS5lW8dVSLwUVM=
`protect END_PROTECTED
