`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axNL3YxVlPkQ08HLaPYk6RGrq8DFXKGkcrZUm/HAy82gvlLgqKnZNnlXpUpR9H/u
BrmvTFxTzgqR9huk5ATNWKR0aRcO9xs6k0P4SMeO02nuePmKCYYjETEcyOfIMHLl
dan4LGRQu9yOdkb8a0Y+w1Za9kIHvnQYXNcAaDR2Ws9UOwfgpKPEM+jkXfqBKRNM
/JZpnmzC7svl4sPodB6xOXzwzAntFgta7+Gra4jkF4iFDfcpyG3Gz8nOnHuimQD6
252vz2B2zZrI8+QnbZSDRO6f0ENkwk0jXAEHDkWOnrYJGQr5s9b5njYaCOEf5tKq
J1G8gKsJo7kRiPutaP7Mxzm/ZxeBLj3WakVlOCLuufMOZFxTkyIbl4OkvqMTYWDz
KsdPzEyHWi7+Q8TSo+8lmOv7lJwrOyY5d8MVb+VaCaQU/91rYLAsZg6oLqLTuscg
sMsM8SVVnUYGHjqVnW/juf5D24vsuL7cnARr8aLh0N+IRMQu4IU7pvv6Oi2jo/FW
DepFWl24rJmo+Sgsh2lJvczMnc43UnNj48E88jY/rUeRgYy5iIzfXkMHNos51sg6
Vb7wnWPk1wr0FkS1f0SFQf9u1ayn4LxVzoXWPT4gzbBTWYwhtxZ2TtewrkpK45bT
Sac4WNfMD4UTkzLAVpmnh4G651SY1p600UMNtMXCv50=
`protect END_PROTECTED
