`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFxc51K8kTUSm4Tz/moosIGDcLH0ckSm0tt+Gn7h/b7AqMESAUCsQ3ze25PPlA/P
eNPZ8G/OIRpvuQBIL7oU6C9bOzbBF4DwF4kVGcgRRCyYnFNcH7457ZvokRLZhgUZ
jZfaNFabpA6yKpqK6ujXWzcRS8oSHl4yIgCY3Foyw+jWAtyiUI4n/v2TOxsmxghC
4Fz0rj+wDCfy5iV5eKjSvh0cMwakSwkopO7GbJv4TFowKY3fiPS4HWm5ffEonP8l
JPcQ9nQE84JuPsUWgNUdg8HxHTKHzd0Iqt3XCbZXrCYLlTNPbYCyNmn4DC368PqD
G7sNFNvKAdhkyl+AI2F3fFQ6RXH6XZlc16pjdcMuqDqPkFwAUEcMpPzjp6kry957
eUgea3OcncpaN5IHKxDpm08PtZqP04PYR7zq5pjf2YC/0ryy3OPFPLHFzs+gw2wR
e0HU0or2Cn4sPjpmR03st+ehP2V8lGUyE9mYSJ4cyyTRFELX3Bmi/j4u/Anx0h4H
DnXw8eUVEfZKLNZPlzw677PIz52Udd4ZXsugaHsBUoXLh30a3YsIVNO8CZYKsooN
KihZu+WoYWjwlOWeL/4fzc6M+AaZ9vGjlikNE/OwBnIb2V7UO9UE8fAzrOpK39xP
lM98o14MdEFl+YPGz/SJ3IIMtfv88JenyEPDM1QJPsZxp9YLslaAZspukjmu6UUs
wA4/lgpvPPbxxijbsnvjGZ/JcqEMqtuwl54O2LlFJlxBcQVXYLqtWMguYixRfeiV
PKl5/PG3pJW5tBIwHV8BCaZfrNVPD86rGSsbgkIn2kOGvTxkj9I+WPq22UVZ8nix
a9HMjKYXvhblUp7dpSlHjH03Rq7e6P1bFC4HIeShz4a3FAOwV/T/i9ESPcc2t5jM
or2ecsBMquRjl4UENG7611Y3W756ZPDAKe1Nm1hky+I=
`protect END_PROTECTED
