`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNmRI3XRS46S34Z7oRQJdoKbDQPTtP4vj2CBmIHE5Z2Uy62FeSWnzzET/aAhTcgX
S4W6uawspR3J8IGl9pM91hybMSQQvgnjP2Y0Oc6kHp4gU25z9kuqMeMpfFtQnk0Z
rHVSI09rvSe8ZE2Hpp0eVF53ayrFDUiK9RV98wCs4X17GpYrxaMJqhjzDRjRI8Fr
zZ0Okwg8AVsf8tyS3kPto4PCu8csCaZMdTrpXKGXvDNCTg/gq7sxuiDin1rF9xXS
wmhh7NkqVHv1YaAs8fBkg+WR5GZwrAaFsiBgPGUNtEGGULocOpJBVA5Pp6uvQrw5
6RjNZgN6jKoNY5nvrF8+PW5eOHXRu7EBgkGtcUxulf7oWHLy8HiuyoTHJfMVn+Pr
10EwdBhMFtS+0pjtVjW7PdnILir3GdcuqRpq+HJHiuDZHIg1gi1TYEsrOBSXeFTQ
W9G5zps1bmr6zbwBj2WalUUUz2104//x9uEJglAlQImkCk+YULUjWVve8GnIdoAx
vKn8madpmPKkr8QeXgc3RqXfbbKw1LbkN7zcufDqwbznAN6GvhwluzTZ9HzUHNDj
Jr59AD3JOIaom+Cq8PZDkks8ovkInllQdsyhMJoBZRuIkfDaIES5ZmMeYmtU7FPS
eepMZHYVJKeNzPABzfVKfg==
`protect END_PROTECTED
