`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ewf/GiWNmEHUCTy4LydAE8CHiZM0EnQYIMuPA8yZY5Nh1p6kavjmkbHP7CDicONb
VcvOHOV6esNwIVzliOa2RHWf/geGhd8rCFQQRCTzLp0GqB2Fazrbiaw10dQPY06a
Etiq1ufe8pjH2wSgrQZbQdWBep2gAB5d8bB+NR2NgMvXt1bz91hxLlLhZbstK6Gt
LEiOU7Bfn6UwkDjxdF6yJItSb3zTB5VHjd4dieG3PQ8/i0OrQq/FgGQaWtkEbMOg
FbJMI6Sy63m5vB74w0dop81mALmDnRwsvf53rza+5OIX/LXJIQmd+cAraQo4Ssv9
lcdiB2DjWlkLwUUcLpe41pGzCuU43x++Wv3Zf3GN0d7FZmBVvy0YjoGqUa1hTVJD
J/AiZpScByA+43hYagK1OO98R8j2PnL/dctIkOssYpiogiTMrUWmsOFIDK8AZ+hR
l1+t0ftU7tqu5kahVf4HtVpwzgZyoo3ETyJullFHattC0x3p9F1Mkr5ynBZYuDzF
D2Py3+dY66enkKbixuJL//FkabW8bZtRTlChTpha0V+Mslipg8FvVSZicqISHpQP
r6k/DR9ckr7g0Ko4bq25SnrUub4gdgBNOmcH+mRY3HVRTlzfSPeDVa/hzUJprA2d
+ybxb9pCmqp5KnEi+AITpBK5/JZoa2tq7oKQPGf4+czEim2INNFLbvQyYHiuk09S
zE+lvoheSh8bTFhkW/RE+7mdrSyuN/5p7H/X/w9vatYcLzQgyVqqW0qch+5ckr3w
0nd6ZhnGe9aMat+ItNRtD6lys6J5Z2B1Mfnc6ge1ntt43Z5zwWR4pwFYI9eaNgQN
K7lUPwAOLiEiNwOJKWJx2gT9RwG2K6IAHn2RTVdtZ3TBpQS4ERjMulgp+iBIZ+fk
zrVNI1wD6n98o9vw64Qcx3GhXOUxlZdfVbjvAr9jndE=
`protect END_PROTECTED
