`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFOCJK4DbcbG1R/tJCBbbwEl9Wp/vLyIs+wMvl+Voj952nGQocSNZBPIKJFevdHG
1Y3ECeZYk7buRwV/63i5SmsM/DZKsl73SwNohxzlhBzw4BgKMaFLJzRkewfNypaN
pBmC/Qrq+iemZnIYWR2ORYJMCI16H0+FJ6QxKtdJTAADX+hGAoFLxSIQDIXKEYzt
3sgIvfDqVMTdlK799jpMqmEIKAHbmufC+duQmMZkx2WUhu1jK/fKIFAk52fOB0xp
u16OExgPH6xZVEmtOJD8HA/nXz7o+MWf6IDjzaHAlB5mAXqdaZPJC9GFNwY78fIA
64vAGHGqzkIQW9VQTwqOZyhUAVR5WQ8x3SlNt0XDIwmyt67Vmv8rbuCYUGosZzwd
buVPfJfnrq7v9A4i9us0jJrvQXCsyOKhnnk1Jq+XDymUy2KByKruYo5OehrLma3o
djl0x1RrjKUmq1cL2NFHyP5d/DET4ngY6ejZxfgNT6JMlF6c7YyP/WyOn2qIqtW+
KLW1B9vfy612CJd7VAyB5QMPU4yUWYWf7OeZ2x3Z0j6/TnDEl3q/cDS9eutGFmj8
YOON43UnsVUDYpJ0X77UIqooZcTmnysLy5R12tozWbGyI7EA0u6gwsy6UalEe+Pm
WmbQx4I/utKlwvXnq58QuP0JcrAlENeKGThwqHuZSLRzQCIHtpIjbnsBjmfq02Sd
cmWsTGA0RgitYgqpQnRkbfHXHf3YMMIGe9k42zY4NpVFfmAyqZ1mTmjmkIkB4Yc+
UtiCR3467zOAN3HGKuqTFYlprJjwI1OHSUn9oxNgtDOwjOUA796MGxpVqhlhAKQn
xP0TnO9Jema5tpAeB7DgZtjR9dYV6j6R23/jylYcYG2LLPXnDvjZQUwHPvQ6G5qL
7E/O3+vYSy2XTogSWJ21IkLFM4fpNc65NhCHoTZRmcwfmWblOdLxpHwJuAgEkP7w
JHcXM7xLnpeKEC2J+mW1x6qZX0wSGIxLuDJRI+TotNgN7T2uta40DE++Wlibr4Go
Eo+NEbZTH4ZY5usy0dP1qx/WJeEaX6HyYayR7yIZjX9zVc+yQTUZuev0aUeh9wQA
327/fh0c/c1JszwPi/Jt0MET0V6ZJr0UoFIG9z5VlM9OyPtMLLJuldzuOUuj9HrM
5BM6YqC7iTyz21iVbHtBCHV1a7jifh6T8MvhpKiuWfq6PF/8K6fdL0boZ4sUOtRp
g/LGJpVMEGwAlI6XcL9l9/zZGzUtpJL4WySIEUWWN2xJMPDCpkMrWPHtobbFNclo
WO1iOcpu/qTc6Zlb9F8mQxRh2VsC/G2+nXu5xJ3NMDqZ4KaWr0x3ffX1wEJfWXvN
60MJoOqSTsFGCjgEY6ulLFokhMdsQGjksid/GyExzrbuHUYRFkn+eX9IsXJqnGm/
ex3rLafwiwrMfi723VuhwG/7gQRoGg8pX8WR0Nn+xQAquBvGpSkfiwvIbhJ+oSzw
LseB1mYhYEJ0XVI5eaQVXaXNWb6nFbxKdN9mkvYrdIs=
`protect END_PROTECTED
