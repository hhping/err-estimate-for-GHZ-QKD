`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9ovqZTGCJ3W4jYI14eDgERmiX4k1spi5cOWul+nljI4XDdCrhmS1vz6B/CZw+aX
cFUCxkNAOgBp+gBUbDQNp0tvr3LWHS3yfhWmIQXD0tR0CEIFNwtd/7UkFVclYdWV
IUyaUi3V9slnROCqksgIWRS531nM0M+3NmJ4o8eVvVfeko1osLQwN2APdDopOSPu
DM+mfopo0/GYdN3NiLG2jLeZT7NpXJHWQa/ZNhTE4vyKIOpxhnYKpUhUFmGHNh8L
zg1i9SgAtwqy5EulObxA6g5IPWvm3/siUSG8wi2JCuVViADiEw55GzD0MYDFIDag
BzdJGM97R+XQQrI9ch/sBqK+oDDhhMROviDghiI5gOPyS1QAK39SHoMtcfCPc19G
3mgoyH/4DaZnZa7xTJbG76JCRWysWMS1hocWIJVq2y+cqt7FJ6PF5P68ehfR9JnD
/gNllqFmvCv7ZUXZg7o3uyfSmCbF51oqRrkuIaADM3y6Y+fnl5dGxc4AfcymZgdm
02cFLubl6lcbTq1/tKwAzHduoAfK3NHVgQIC580abLdL+fTLF01dOO5TCx+wwH9R
7duyPOo//bed18kYlpuOIYFAscTRen+/dTXBLX2s9LZ/YnDxkMP4ebhTdVrs3kpj
Vb0VVGLGv+bJLf9WSJ3TXkKsVDstilBvMWBImTjQWqVLlN5GUsZNAvuaPOfQoT4M
EZ+bwkBX5yAF0nh6asdLYCNTGnSY40t3pwCqpdtJ7kgpzPh/FL+gk4HC14l1zJmk
EJEZ2Tgi6iUvI4zV4r5FSEqTh5Kme3EccmuQOGzNOOXsqJdfh90zn8mhw2aISZqF
E9zDtqltkqcQkwN0n7qV/KsI6bmvfXHFbiiETPSIS0FirUddSRkG9353Twf6YlqH
Fmge/MUiBXjTDxP7I6wWbdaZNz3upoLNL/ew492sjzdSWpzcooL1/FseSB+x2f4P
gBoy7ZMYlpuAgc8npmd2o7KvmzONmn9yelJmkg38bEhHxrtfFRZJhZwwC7nw64bB
r7XY0UYINczgpZx554guoWNQf8M/pvNsDvKBSfc10aGGL7rMfUwyZjFMVQ0M9HMH
1xyiYfaWRcaNcPjc3j/lanOqo5p14f0dpXJJqoQ9b0X7Ju+aRtSfiM1fxMJbLYUa
/XtqvyXlHWolnWl50d/Y2i4cu58vwnCOySIUp9+HxQBs7LRjlQPqWlnSWcVTpOIt
/FWC36WTQP5pvOKqRAP3iSIToTP523BMsxPj0aiXBBGGSamI/8vObW+ncNAsKbFl
ZXZ39bHAn9nwcbD7et+iqBd/BDXLKDcx+xbKz61QvV8PX6mqTTr83YSCqSCMRQpz
BijFoEnne/ZuUpRrEaiS0SPPXVQTb4iU3t2iFI/i7vWUc79zxr6ZM/XTC4XR5FnC
93ChmI2DQzvu7aA8Gv0LK37Teq0F4Vsh+S3HuXwROLR8G13xgaKCEobsY+fZ3ALK
dykIS6F8TAaPELAVyvTV7/GFqyvuxw5oFBA06nZv1qz+TglvKah97eXtmzdt3bT3
cQXTHqGnklCgjmSfjDLD5wU4iRs+fTqa5U722rEjoHSnoyBbrpMJjrfcewJ1lHlL
KYauVV7OmwmeiG+VS2hc7gvC0r1pmJ6UKXJFzrncEnpbb1tksa8PtVooPTRPW47H
mOtnDbjIl8NgxQkZQ0eZAIvSJsiPmVc21u9zRW/YejsDl3S8pzPD53qz5ThXMgSf
ZO1L/FBymu+4TEqW/zIUFTXkWkr7wiR7nsVXdU6FcwqIPAMfIH/r4UxTDX1zLeo6
hZDmg2Xn2hgTavQX4QS24FeMrti8usvuDqaXegwmOodwKW+NVZ+I771oYOIokt3A
qlPQJr51np3LH16RhNtYjPkJZBv4ahXcKwQrNhde2gHuEUBUQ/Bv1MWGSasewSQv
103mhGhyR+3j1VaXKqwoMdxYX1zoBhYTyx2xfylarLHiD1pxYJadUZbGTCubl5B8
WT1y6h26JGys0r//IUa7YayWA8xYyoPy/D4pCek+loq0CeyGriFE8UkmDsr8tOhe
c/UmMrjIZ4ydpcs9lIlqIiTL6snrttugE3Tnx4sTIqwdzWtNIPh41pNjvnyqwZBa
`protect END_PROTECTED
