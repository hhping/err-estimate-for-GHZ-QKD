`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pevZULXULL9abpV5PWLYGta3iY09MVrfoPl4ADkDR26huuYEu+BfgDY7VCYLOAqK
0Gd8MdvAsdFdI8h4SVeUyAN2BZuh9X1HTPVyPsLNA6QnVRhsc4iSERrLJuIvx+fy
i8cG4wZSHRlNOqrjWzimDEllBpshhvBc/g4yHtTef9Q2UmTGa4VcBdIKeTH8/5os
rQIh2GpLaONkBe9FrSbdQ/lEggFLVN/Vbx7ehv5zcreuBAcxWGOs53wTzRl6mFky
as81QxGvXKK2z4/pS1i3cVVvvnPASUBEaSzRoaa+5ZgGtVK8FIW9mJmPEzNgLkqX
S2Kzyb2nxVQlKWa21JadNXyRIuTPuUfU+9DgXuBfDi9S5jM9GYvOlKWAPjgVTUVg
Hxvt4ZjK3QmvnzvYF45Ark6yHLKIaww2rd+xEGPz1ncB0Zh6a2xPcQPFIATgB7ut
eYSog0T3NGM71XRQv+6s0PPHbvmvuNrnlU4Uz+HcnnYSHd4S5FEG1cf8JPee6vJo
fsc1ISs8s6AvbraYdE5DCAt0s8Ytvlhwh6UsZsPdi0j0778h/1oZn6KRGedkKFrx
bOv0SlfPbqz6u3Ycf4rRFFVvcqXMXqaaXHKlj8GWtxAVYFn2vCaIopikehOUtDyn
OrJBIJH033azUVPkq8i28pT3+kOljKZMrLIxut3C17UIkvHBA3R96jdqPrOnvLI3
h+fUqQ5yPFaevDQ+faoAVo1pG//GyT1cIE2XdIG44yw1h2BcPtel7X4CUS5MGY+r
gWngHvxZRBSMKE66l6jDDGFcfEsT6NnmXNNxZ04ogGYVjAgZ0olf/GD8rQNDGkwq
HmXxiVV94BVcwmHrxZj4fOriqJXLGtYj1faWxwrU4gsQJWJ+eTH64Av96166BNd8
LkQ7h586TrYNv63c7Vtin3HAXshw+x69bHlexLNwVzZ9AXP9gfnxyE6z2t5705iw
YZQ8SlU4ydIxBzZvcVWwGwK4kXQX6UPN5CwBM82J2xCeBuRSR8asmSdLZRySByEh
Tbj0mhBHDWxfQj1wLbVH3htxDnqejCM5kI7/Z8hycHKA00N/QxYioB12oHr8ANVO
gDxcAZN0qML2EmH3f2rZ7X7k/3pjyxeu6A1XmqflooCcCYIs9MmUwoXKkgiXAEi8
+3CHERhofkMmSzzqMM/X5AUM/tf7JOpI3lWHIM4lWWDqG2dmpg8HPdYLxbA1I5Va
Ef1SnpSh2rDN1OEHlBjO9sK+cv1lvBzAgf72kMU3ufI=
`protect END_PROTECTED
