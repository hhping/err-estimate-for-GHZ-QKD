`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kDk6di3ps4fsymaIBru0fg9Cs1lZ8leFlYRPfHoBkzZ7j/FZNWGj9CRSznnngbNg
3CkMG7xUIUryJoMwRHXypBvP/JtJ+6UM+aphc0YGaUPJVteRanVFqZLzJiNW3zbQ
SpOxWtmCQB3Wdfhu2FB9Ds63kuTdd425L3FlI8dgVQYjZR2x78Cwz4HLx1DNeoid
1qipIvplXgUVk4Xfc3W8QwbjvWRvSOVeiQ7Bdi1SvHMr+vrqGMqWfh6wu9GmYG2N
WIscGPL8gl9XuRyE67eSFUMnCdyfEIFwZhtV2RdufTBWeeahwV3Xo11KVraAVttq
DU4cEqkn+ArqNpnolp7XvVO9U8uNr1WSqh8CFSJS37Habc0DKuWCmAXSY97Aj/rJ
kRunAF4CzeVtpvOqLUmABk445AwwwH+VJGUE/Nq04dnvwXtKP1WPmlQ8FsbmZJn7
QGKg6KiXqTpQm9Bz3c2NuOwYPiffQTFZWpMtNSiBxV46CDcGkEvks3scqVlUu4mn
K4TIwmV5mf7YPq31lBqFAodgdNq7sVUB0APZMyfcAG460cJSzwREy890yH9PIqPJ
Mqh8RWCxQamxKV0oNhPcvMdNQtZg6aVHxneYXclE+pcscmEtwayWFo00zNmagHnG
IXF/pNRtRmniPccfF+l/cynlbJNj0HTkiDG8Rv/Tw+vwtqWAGjIsIuGp2uhIsgHg
PWSUWY89XMEj+Ml1DkkvbSLCyTFacYSGbcJ0+DFC3rwmD/oHq/MMlC0BQ51ZInot
cmuvML6qQuLQ8K5AZXLSDvB3bkZfeEXlp6AqdrZsd5gHyfPbc0FpyMXS5WixYs2w
q+DXJGKTW4k7Rmnol3okPtd1TJEUuxZG0xK2ZaJnt+khb9rLJ+ffiaA5nggF8DdS
CSkSzOa4l/pSmGXXSt4LVeQ/oj0LdunFrKce/tWJv0RDAAElPzIKlbgGtz3xoyuo
ZkBrt3svfv+TO/JCRDxs9E2XWGrVEsuDTeWRpL+a6hcc8aiWS8rEcEWkk7ztXWMr
By52YPb1aZhOiPhrP8rUDTBh7myBflSUiLcReeaV7i3xyygejykqi/ENCuV4WEJS
rzBUIapISwFEdMpQjsgdG9EB7GUMx8f1hBwGidnPW5PxK9I6s4vLq6KAYaQfqn8J
7ZEKpjZYMwL+gRFS5p15VEfeQX7MIoLeh0KZVBLfgjuvu5Y611iky+6ndyCanMeX
9dloYBNNH9Z75okCtFewNHz3ZKLCfO9W6GilvwYhV8O+bXw0JXfRwboTw6gvKwsb
MbYfsahmj1f+TVVh8TGB2+F0QVOaLP1WKxBVQRmseLMu2+6rzR+GApjGc7naE+wo
W1HA9bIWfIGbjzOZ2gVJmrl0/SHujCu2e2mdpG11yakG4Zoq8iz/1rMAkB7EVLoi
NmpWkT8cW7zMstdU0ULLVcjxB/99Ppi3lyrdzyhTwbbYAUqhWxyDiivYkiuHn9D2
63iUAaNrksf4VVzHlt/u3gBLmibf/i37PUQTobXJ94wsRvROfSZLgvUvZ2M3ut/l
JH8dPWVfyB70IOuMWtx/5OaCiDGHJoXh71+IJfIYfl+eRkl8ECPBZmyzWxOSyvxD
ZL4XJ3bLCqhwBip4wuibrzv0NGeo90V1HUae/DnP9U44TJ1uiKX5Z+YBCl3y9crV
FZjPyw4yzJFFveNfeWr1/Z5z3ISkWhkp2K0AcDcUb1K3Fx4f/UC2cfD5oJWk+SEM
X6FrTCQUN1xI7rBIrbDWFeYUZ8zWL/PDvd1aqKVc+hRINQaGX0CIqiW6A4xx3WbL
Z7wLJfl+0SxDbIaOViM55b9J/VVq2iXVCVkXsYqae2ah4znQwdyEfHvql40G55jA
i7pkA61M/yYoMzlfGUF+4wzeU09Jh1iNRsbgXdwc29+0fywPVaC9H8qVJJZMbpGt
BPkM1a++fX8V5HC1RiCqyb3m10SSvnFIIML6KL5z0W8dMtRN1o46CAF8jYvxFPtR
CGtav5BLhJcsgBbQtcgbjEVkTsgkdnJXc8ZQUn4/4/jrx9Rrn2Y9m0HSql9L7wJq
U9mzoi+Fz8ss6hmG+OGN3UG8KbK2B6SNEYK79CNq/QSdWrsrx0uSHfUmRIZATa8Q
62JJhSJUuaj1PllGrp06Mwl0SNB0kvD/rxmMTVNCIWRxQRkaxJu8F8dS8t0dhklB
erEAlruJnCyq58t2GJD8qNU/Ho6RhgcYJDRmy9LXlYX4PCQ/oEyoU6WcSYfiNdqS
PqxL8jZGHhfNaz1b/yCJ51pDH1vsRdWLLmiR+lnZsfOBi4nwU1wAM9KoirGIQ0oa
iFPW4WylWfCIZXZ5LZglgikA7inKXLRFV9rBZ8vUNGjXsRtgWZWmgybcoaLKsPXY
NJFRHpK4td8oWgqGlCgfW61Ir75JjLyWWvcOrsF2rCSeo3YRX3YkRxTskiv+Hw/+
BKJSbB8wNP45IqZwWEz9AwzRLMIv2VGyp58TmXVQmKGQIrHf6ZQyXkVjx/Oy8Sph
IZkyn5fKig4I4jTbgFcnHrk/5u7DTIhIh1zN10BOaFi79+GXyeG1CC3V62oKRneT
16WS99foTFfT7IkE+SknNqaKDVKlvfm1NqHTUy2rVDQ5YmLDugh0/fN7WqB90vPB
qQlKqYCT+r565NKMqIfQT2EpBGTVp42/o/t5le0zweg3VZ5ZBv4+vyEJECHHOhty
aHFhrNVNzcNhlKScyItq6Mmx8HheC3c59ZJYOdr9NN7nsMd6ub2//gFYY7chI79A
AA3q6tRTigndU3xfr8mCVCTCPzvOartfILlOEMKIhk8Kw4P1//RKupkhhDA7K9YV
G/vljpoLofkQ13f8gn9zkNYhgVEx5svXcXpaFkgRbs7xwq2c2NAAQ0XAdJFZrbwU
kveXfzTGGGcNfzYQ4txOcM3rlQ7ujUZwPgFBtHQJk0t7TNwEOokkiYPyNAZFLxUI
bkZwu2GIypCGSmJ8bLgNrJkGGyj7pe27S0hWS51D0EmcUHzqB2OfXp932TJOsuEm
70yHD8v3x5UezY4sse+3+d0N7kSTk7qLw2xhfbhCV0RipIbmPHmg2vDvjij/jxu2
uBMBHUFirDU7aA3TxNMYXOSOhFehKrBp7DRocNX1Ciz0lHBUMr7hXoFX/HhVNiLc
IXIinXVQIWGmFxX84zI//cFQxOm2rtHd6IgGgKaVC1xyDVJP+bg0Rqv/7BAT0vQD
VoKwNZHZS49SeGgWT9milT5HXIDKGt89c+18rH+8GCHDMkAyvR83k0Pd4ld8R6Fp
Y5cb1Awez0TkR52aOFzXMEE12ZUzI7VSliUg8xC8hJ4y6+y1SIDTIIh/l09xP8vQ
D4qmCNeUEmuLEgu1Rz2aMl1TiQZ8CL0FS06chDWv0jdtcUyK/DL2mQJIAlbSnhKv
ghJ9/XBClMdH2jlEPXSFC8GHYToSJoAIbYfw1hhmu1D7AR2dxSQzUoz+ujGK8wMD
YkA0pQAQP9aJCP4oa5sAB0+deK4gG/CgMxZGL5yhxreRh5DONpVrgJimKdV8+sDS
+pdfgdUPbCO8ZZNmH3A1GPy/TF+iFXznI7nLUvIyuEqa7QVCQp1rSPSJyBmQo8wI
yf3kQgo8ENduK30Hl4kdljwwN34COKiGADL/ZUSUipG30V+XfBwDw13D1hrUMvHa
HMICMNjOHs/77EApVmDGlCWzel50PUQgzGXmSvndHTiOQT7siXiK2s1eQ6LbNi1H
VQO+daO2BfdP6pV3RZX84BJix4Ikx7yThJAxd5ZlBaY4pnkbvnNIo5Kwpd64UlVW
Z/vVIQBQdcy0You+jDGwHi7pXSpXrm4uupxIvbaWLH9an+Ytn2QouFMCH4/TYfmq
Q4st/qvbNv66Q06wuS2eKq5PExP0CbNCgzqTbjR5G7TmhZcOCsgqbcFw8bUbW6IE
xR/TP5/Y1Tca0AQ9pAw8oF2Cnq1ctonG6nat8NuBgYE7ZFZHR66TAY6VmdK5qCVc
0Gu827Z7cMh0lOPsK54tC3NDdNAzBC7nbgxRpv2HzdiFKrt2BFplHDwFsYGldWRR
ZzDBHuZ+Vyk8wPOQzvy/t2TpBo1mVKAcwNhPKBvVnvM7aHvD6QPt7Guoq7IdxRmw
7H6gu/i/qMdZ8KEzVwy+7yvjtd13eU8HGokwOyxQ6axEJTGaZvmrKKJuG0+58SGQ
NjNsccTofgYINXe+9CStq1G2TU3nRlUpRiMjQODpCDV1FpGeJcxd9RJhh3GCVatD
v3MDpfJmm0bkawQku31xATYVY9idUWjtTtcdnsTAYU+Facb5ygbF0LIj1QPvNmjM
8eD3IzdgvtL5+KQ+51HF3xmljU9VFo+1ua4SQ+KTcxkQM665EENwJ+0x+QcyZ+MP
4PcHS8OqktEonqztfSv+pj/Tv9tuFYwMfI0RRG3XijWdbX4OTMqyTXw2p8sS/P9P
V8yh+11kSYVCNHX3LBWZBOoKgQ37Gj1nioLtLTKwLVvrnkr6jUvVL0P/Ze5yIA9H
DBqChoI54acPLfj1CnKsDzPycBt5GSsydjxbQ30Lu4TfRVNZ6KVUNSnvZKVM46GL
XRxvi4aKTdKCDHesZ3Fw+1FkzD6iKtwwxMg6kyXouE0/JcKo4VzGn7QR3P+ag4zK
LL79TAVSc98Tvfe42D0v9RR66e3Yvon1H3ekyYbjeHWklY4Upy1XakezLrtTYzte
PPjsOnG2ZEEIZMA4zA3SivmxMtMTtaCg3XXHrWILjwP/I0UoYyVAhKFkhqSMloJ/
qPCVsQZ0wbNx60DXf/7dvtItwTLCyliRtZPUeWRbeRXTz6vJPqYqaXYsux0a6Y2k
ztNgmfHq7dMnXtRoQr3NrRs1jTyytHoAU+385zUpqZl6MkbYGXKAGg2PeWKFT4Cn
7lE+weF8RudJJc7rC1QSbC5/CV3s5y0WC3uORlvyYblC3yemqAth/68/cZgm1rDH
Y88Tad9YdJJEeqF5fW2o6aIowlpa35ocMwJsanM/cznysLEAIT7BQ52riVSIWYvl
/jIb4gQPpICGH/wu38ZShf6JXnZzxG99yZHMY55qTIA4ucGuT3vm2zRsc5L2Fmkk
UxfNQlptOFvTRtFopkKaYIhzSD8CDbmqBgkoPp06EnOK4IJTuvzgi8ivYZ7PAwLD
E9wqYB3p9xQrAgmutnaemtZ5V4oPBDu1iah/LxxdrS+yPWlR5yddtej7+3kCSopx
6Px8vycsj2Gd+ss3mWPiRYstsDKzL88HBk+3zFcSSzBtZ1Otzvo0eQ4z5REMzbK6
ihenCiu2E1uv/QrZUmzSGtaZpMV09GEfCZ3ssU8nV53GReUaEQjiwHe7FnWIDjy7
9uxhFI7TawkC/Y7OVjHN7YFTRwdldmaP3TXqEX5myBqy5Z57tWPWQ0xbW2vE6rlS
4hhe50pdQq1TacjZQkxKBx3vRY7JxD5C8m4k+RumARUf/ERDoGOMgs9epuOH5rfs
MqlS+h3VDJ6KxJh5xj5L+V3TC6/1dW2mSzh2i5grCKniysoiBILvwxYmTJmwq7Pp
BaaZY9aROHSfD8yYEvPVZqxMG4BDAsshueHOWT7OurNFb4qdBXN3jfFIomzGzpH+
IQbgaZlFdtUChtOCGJyvTI2GSe/+U6fkT6qbMsmpn/f6QU28SiV9yfV7h2Q4AsHp
fc7QrVypQ2AIA9UW762/22DeZHIbWyo7ozrxS7veKUr67qs9CndX2S6ek0ki76Pw
K1PWZcc3rJlBOuvxQBTJb9MLytHstEugJCiOu5Ei2eF+jDRop5L/aWAJuvNQ9EsX
eHwCV8A7qmLuottuyX+PRj8S6Tirc2g3inlF1bvYEcB0YthmRfql2M5PKCOZvrqQ
EcYOOQF3Sso8c7h9DWp4Wlvmm/rXEi1z2NcIlIbYlB1AcgoW8nTrPSaT7W4uSLj9
AvbZ2XmyC9q2wHurWfpu6cOcl5batZ470bclc3Tp9qxlUw8xgdMF4JSe628jvt76
VqUdoguPKwE0lHKCU2Hz3gtqLSJdmX2GjBzgKCPUagMoQFM8V8NZNZrvmEkshKct
Ox4OZp6Ge0MvSCeto7llVNfSmud528yvGnrt5iRE7N1RDZ5xqT7YHmhum3i8s+QK
1LCF+kuvqjw3eL6nOEyOBk+4VWore1Ur119o8kf6/qtGTlKhXWhXtKqa+lUfx7an
LqIK78APIoQlswZY56hYLIL4sottl7YLBYIjPE1YuBlPXFLXoXrQDe/sh9Nhw9uI
0mdnbrB3hOVi/G3f4BGuuMobihSaIxqt8f73erDKlmE9mdCtgzPnVxS5Lp8K6LGv
S7e66Bg4ffQRT+9Y6IC9SvEhQ48jWy5bmEoov4alY43WItIU98t89u9xXz0XWoIG
FuAJIvZBHEns1t/bS2ZY2cx1OUosBsiy8KekwCtPOP5+n8AFoK2O2vjWohOH79S/
x1ejPhxdTaemLWyeXkp8v4J05UvxFiWvIwHqdXE52wzPubIBo8WMN3DikTgP2HEJ
cgz8EOZt7VlZ9AbNZEhiPq9ZTi6WW8Z1/x4I7gnTOqUtZLce38cP3qr4iA473Hay
NrSdDMaihu9A1uhW7MR6KIFaAdoMc0Y8rsgkQKNWFtubTpsLha4NYmttfOPYOdfz
mmrqYDFIRd7QEnYAvtuiVaQp4P2HvnmRVAhU0PLlmsuzZneJjzUWegrQJhG96F0g
6/9lX2H5236+NvVti0bmQ12Q7kBD9FuT6cZ/vA4YbBONWw4jOLOoLFUFgA/YU4pU
bg9I2n64BeiHtaLS1Ory6N3IiZwnbrxWr46f6kxlg2gy9nnDBTyPfy42slML5m/c
Dq6YRZAzbkSH38+CVNnsglwI7DnYHE+OsnMVJ51+vhxFuEPCO4fkp+hRtHuBDEa6
U3WyBhGPZuZLEKwS1ASX+vKj9UctsEkczFl3OJtDOYl3tkSjcrG7dgv3wGjbZPrx
R811KD9BHBzLOeenKBi406oEIWNiBP1nAep/ZTAI+jiIRX50K5kDzcFURiy6HpmN
jwiPEhCJhnr6oIFefrJccyht8GBElTEbf8k2t548huEmTbNfmrqjTZor4GeScaeq
f7CaHfl9Xq99z0DJM2jk/6YIh6JeQW/Ety1c3Spw5YkYs1kGpQoJd9Qu0tlyoLP5
dyMPhztt2hCzfbszESPXLqKiminsr4FV7URZRtrK53S3OTG5yvucC9+aA82Qjswd
vG1mhwUAr14MTX5XhDmxPQuM2jTsXtMG03o+KwsqxAaxOXyns4Ej9nXEPJ0z9dBl
DryhXs4EIEvhJihPe8O1Doy7IdoWz4eqt8oQEB37N6O/uMf40gkoxTE6sRrTwuPP
EWgWaLfemccvGCZPJW5yPz+VfWZQvYpiKBAP/Ba3yxp+kVovLaKgyY61GOGnblZS
SxqiC+DEhmx2io+856mO9Qo+2d3wW1XoPMOIS3YvHu3NZc4UZL6k2rNYHKhyVagk
VNhQYOpfm/luNLmNnZfw1w/wbwdM/bWCKfyU11mrSV+FFkV6jUG04lPaDDLbVLd8
/8gS7XcVx35l2mMOP/uNe3L37FX8/Yfva9XeWLRxkza1OrJAahUHg5byQOUT5hcA
gHt6JYaiCrS/487kXQejSIfjjaxZDEQsUrr7mKc4q6DisioSe7yz8PcTaDigC/F6
YJ9s/FXTRIRb3ghVaXAVHtlqQacAaawEThflzKUGb6+5mfFGHKD049JDwnnd0DYs
3VJBTr1Q1DH96k+trBzxpOadSPiy5xpSuXfg74EnwsfwcpcKHJZN0piipqqCFwPd
3zYCyCZKOYRzbp91dXp22e4eCl6TQNYoX+m2z0hzxrdyVUXKE5i9qn8yF8X1T4PT
4W1EjqGgNZ6gjqiGReSo3u7mr0NOgoL+qugPek2q16eSjbJ/09OcQFa+9tITdBR1
5bDxASMDeH7EQIJJRbCNvqaH9sxDKREB04Q2LK+SCCSe1Y34oabFt2J9tZKvl+Hd
PBf5q8/fbtOL1QaJsZ0zeTDCBtTnDwtWE1fw9NxCsKcbipq980MpywMuuSNWaIk/
CydWXXQgB4m77wQpXoC6C1/hQIHzNz0diqAofAm4MqiE2h8nKvt3YqxFuvWwSQxM
e6t9QHG+iHq3XsPHXsBtdE3itPmvgG04SiOsKoDfUtKhPPfUS8TsJEFj+5hhkh0U
zOlFY1Xwx8iH6b+9FaM5zJ0Ikf8KrpDhKCEzSUOO2xnE7tsGmQ0SPZJPQpaQrX4b
RHMicOuer6ElG+qZ171yPtBwDcUxGEZJML+cEdMeG6/i4EoiPm/WtaeDQg3bNtMI
YIJ9hDifqw2+92GyvwfqJP6ADZH+dyVbq1IpRo5so63PN8B9dHBYeWpSmbDtTp2S
fg9e+mJnsJhxEMekQES7+fuzaZ+Ndl4yw5DI8Yar7K+UpXxvTYAYH8uXHUgpZYax
aLudnNR14Fl6LDMEze0LtfMLVoeQF7WJknZNbv1cs9Em/fgsQCGU896Rzn0iQ7NO
DK59FSfuQKhJV2DXL/kFO07taTNgb8YE4eZlEF2YX5Jox2RCYLb8967LwaQTu2iD
22I3AavBxsckgaE1+7w9IyRqVNgSWT68Ez/OZ1wrIOSa88mNEvEDxswkdMOsduDW
Bx5UBZ6FjC1zXMpcGqC5oeb4s5qgQfPoKhhyFbi7eupg/Y9xtURZrKxMHMX/1Qe7
RFFI0phW1MYFeSI1lRFKXG1cFykE8C/9P9gjTjn7jKygt1lNdaFFSFYBvu1dh4mU
oqEG/paqARznsjRE28TNpPq/KCSONBiYTFYj1zn2bprEKVZx1P5yDkUMEAJWGoEE
zOg9PsTY+L9njAMT6XKDMf+soUYqTeelCpwprhOIwt3lmLHSCA07stv3rtiKCPpV
O5SHl+Ax5wvo3HEI9dKkBuuum/OHDOMXF3JpUzT6XRKdEgI+4PLXv2e08vBF4Uj6
6Lwayd3vY+dK1w+3pAxX8gYp//vc799Od0bvw3SiZUZJs/yU7cAV9RzqyarRtLRf
Km70Vr5h26Ag8y+ZndkNBPrPAonikFf3B456zbh+oWwN6yjEp4vAlmZbHJi8ejiU
cycsWo9jVUa03uI3nAuve3DIsPOHyGQRCIi3aXGx8zc44CywbFVJBRCXCNjGNwcs
oVfGI8nSrsedg+ZF6Ze937Rg7420Dtp/69NN36h/8LdXVU/vaBSXpIhpq2G7agvf
LIVGrw55bSxKZUHJICj0WGR4D9LQJiA8IJmieTT2fxkHcMPjZdoTebXqbJljxy/Q
SCdIBVcVGLVM3CGXVoY3K38/eHyawO5vOKbJfyWTK64fImPaPgyeaCfyDPcc2c6v
C/rxqaPJVAEB9o6pyc5ww9SHYiRX6FvIMRt9LlE8X0dI64CONHQc2E4jErsP47R0
BYDDEHs/tDyZfkgDb/VpSzFguNKPIR+kK7iKPMTZWcMo2lPl3H2WyAvynTWa1B3r
bUjCHg134hTS2jfP1oj2mDSR/eSHZDOl1V/iypXIBuYcboQnDauHSMn7NNIow+4Q
1Rlui84qFoQi9geFBAXGgXI1tNXXPbU0YZGy6dc4OXnHhyao0L9v/rSgFI0MBnsE
7xeAXcLTMiA33zxaAeguORaYrtM1EHxRJPBDFQbvB69Hsz3+dnu/EW2tnSHUXP4g
tAK897HnsCoWhhbLhIqd8jocwdl1aFzVUBN61on1ezL6qYi0ZVGFxrxjm39OfnI1
wAJgDbyVYrBWs6zYvy7JGf+UP9d2jAZsuHRn3xkkokgjj7hMlfSqvdCQK+Xad7nE
xxHQo/PPYpb5lITEoceHqjpmU72twTp1shbED6MFw1vKT9y5Z/a6ktOWGVqk3nuv
GQ3qw3JUKnmi/29PzjgJop/l9As6zb+lyFDU60tmpTKuz9U/mbSMiTVojvDNxtit
YhbtjJ2TgXMtJWCHCQLHdTkABhDVLZV8mNWlpO+Impz1cAkXGBPgbej750fO5tpH
Cc6YPel38snorhGmJfzsSWCmSdKGcTZh9Cf/AbvsOYLBk5gUC5nca4CJ5hgrM8md
vMTwpnXC4ef+10IsZrt0rQRtj4aXbinTjx3H+TLcjdwl4zOTTVOWAxvwAneJIAxc
oLUMnv+e2gOQTBdC7iXr7ETLIS8V38JGdsCP3HYJMuMIGay/IN5+FDDozMJKvhdO
5vPhpKrETkRjJNXgTwHvzx0Df+5kvj8+qUAUP+k2vMak1RKqZKRdWf9Ub2MrLi7V
jz5xQ9RHFC5Fermwo84t56Wk9nadWdX2rCTNQm93mRlmpcF3Kwfgxrg9ZD/6cOiC
oOmo5WZEFZ0feuh3kcv7gdIv69OMw/CltCt9jmdSOBNwDfJHDyWKGOy0XoQvIbOf
ZojDAeaXSDVDYFrxoaKtsWqjA1Pctddg559RPejHOjMu9sJLzZSWuYJFYNEWju/l
uaumyM+SQsLQZENKMtefKHmaqdau0Or/ze5ys/yInTdxssYxgZn+ApztIlB/rawJ
Ng5WISoygFvEB/nhdWQV5PdbeI/ONZc3Q2Ac3urlRNsH+qz0QlHvUIUyON7PA5Q5
kT+c0phizkpEx9jIiEv86MWKFkv6xsACHY4cqQ2jJct+xYNl98Kz1RQKzJGmgmrx
35icrSCOOLJVlp2l+NWIhDE0cOQ/nov0AudAC3HbnHzslhn8FsKmsCXaV9GlCgh/
aqe7+74FIs2jcfEv9yxfZQ0vt9DcMnl7W/65mWJiNbTRNEt7PubCMl4hEp3fl9b3
jS5Caku2vTVGoHpP1RF9bx531P1aApvBRjY7sWZVEr372ZZjxumsAK3mfrv79PQp
TC1xa3/lVqDfWFjfyVCRIweDpwecLl/2bdIuEP1LeiZzwIv1aUM/Cw8t+6O6+jQY
5eJDit3OBl7KF/dBkiyTwnmQXm3jtJ27MJWXBF9dMOb1N2IHdmJVTaqiwG2E6btz
u45y8r89CQzyMnDBxrMBFLkZ+1pPMaXMy5i7+zB4EealhM9p0tMMxTKJVPQAdBwC
iT1OyYwBYj6QZf5Igx949HURGj+tHbKIMG3q2V70xdTGQTs0aiHi8uMEdKBmDwq3
YAQshzlZc2H+0TXF6u82yElMy/18aQvacC5dTOCoQVNhuFO9CIFW5jn/l+9SJRGH
K3/ECcxVaJoC0x86wXyJjFOJmro1lM2CrhVFjewV3HY4cRpnUmPtFufrXaRU9NCh
yps8pdKcz28y4cntOhxYc0bm/x/wZg4kPjslp/i+0y6+hIdGoKakJahXIJBZUg4P
u9P7VCC2uPzodcPwp8oVebP/hLVQpKli0DBPrnCvqRkEjcgBk+1ohV+lt+RyvqqD
kAXurTBZSy9q0+7IHmbZ8jaYrZym0TBFda12lWhhC12vJJ5lkXB2+0jxBLCdSDg7
7NSB9AZaJpIVMxIj3awu8mQ3CfnD6gbC4ZsCDwLieqtzYZ0cYIjv0eiSPxld9BDQ
QKm0EmbLLhtPdTDKLLKrha0r8dNlzJcTPINXm31lOKfYPb2V7cD2B5OOZQbQ45A4
NaNQvhX6bQy2JHZaOyElB7KVJEyUAMJIpMDrQDyDTQfNuDcXQPhAdwb6F2MkYLPw
QQXOC0GzBvPx+EPZcXCvtoroSHCvT7NriDBgB11ZX3orcuO3A2ZFJ9JToxQykrGC
71fazX05bJ/JKPXkWLzPUYiIzmCQLfcgH8jt/uWYdEn9j6+8boEZ7H60vu7Waw1I
tR4cQvCc/Wp3RsSNzD6mpJfYSP4g8wPPvsYFk8sXIFy1pzhRvyb8Mqd6Tqm+gMmK
2wF/mIWVtuiFmvfGaU4TfBWAr9IjlTIOrZpkVdb2UmOxtXqDcZEooc3r/i4Hxxp6
tVOgvdiI0VbuPXt69MCoC0CAYYlxTIZ6fnOXgOuXBfSCP/mW46Y1PanxoE9JyRJN
Mw6nw/OPq4gmHMIcDXNgC5HN509wYXv025YDNcwtgwcR88RI2UEZIuikpFTgwzcF
NYJ4VuoKreEgCkoW9bYTxjxGlOWKYjIo0n47XIGxkBz+A5k7eyYFvaBUV9RxXM5s
DIALKkBhSUv3On9zvHtJeJyPvIpG2ePwXiw3q+UQUhRi8wqlXUTO46jHZkj4c/Nw
5a6i4q3a9XRXJRqhrMegtqA4AFtZ83YCQVbWFFeVj3xEF8zeW/TwjZQqH2NGw8c+
HPO/sBUQmECsdueRzM4kJKpPLie7ZbPADyiAN0p+VLH/+c6JYoypnkjmZdpXY3oG
mrdgY3f2tsXcBxyozYk+dMSSNuRLmcQ7IaezQ9EjT+MqNGAK2wCO9ixx66bHRaBL
Ogn1lMpP4v27QWSB34p6H5iGg4Pd52gYsiOP5H9MVtkRbDX6kWRkvVZJXfYg/7Ck
9Qwl/Xtkxu7bigTvDHcqNZf10mU4MSnREkpukvFhHy9y4w+hiVQmOP5CcoGP+ckG
yQEfOcRIEZwIYbI6dfrYaSygb5fiaJmB3Jh0cbfWuyleNgQFIaxC/6/iE7WII14B
MwGhuCfyUYhYaQ5KpXiFjWevIrYnDQGMTNB8AvLd9VJndumFypNc6j4N2lTCRJGD
yTQ/8XfXzduhn8z9AQeICp7XEaqxnPI5HJIPW3hnveCIPC0WdymEJS1i6aLbUjL7
Y3jcwTq9oYKgEHwmdhK1+WKVbfTL4eaD7Gy3t4sHn/mTe3bnVyuhNN2rJnJuP00g
Wk3s+O+PB5ZOn8Qn5kAIiZA/hh3gRo7AxQwwpGZ7C2xoi47aJNb6zWLDU7myisWU
p5eWC1aXZ1o5SoWBzoVp/EX/2ffa2dfzt0xWd3qHRuH3EjGqYiJsdIgeTzEZwB1p
U/MezzNVhAbLXNpPg2asJ1txLNggQ+vcPwZ29ViBUnw62LB2bl2FcZ8fYWMjx3Tq
g/UU5X69HZFhvazqlWw/wUgAVD2RbjvUX7bY0WIH7AbHqFAdZxzyPLbU/WvmUtNg
uobOJ8wDm2AfxXfmAUEAVWM+IGEwvQni28KS9SLuBH66JH7GmF40OYyOdsd0gXuf
WzNWQygeuEEwT5WN7lZ208F5sbArgMXvxborxaG5cDL9Sssvr70C9hDoLnFt5NjE
2fjq4JTp5w3XN80BwsauwaggWb9BIvyXwLZyTG4OMbFdU54XF6axAf2qtjmWKokG
LgJ+bokPd1A+OK+i3Q/2CY/yEXVSKUBFNTzGLE98pDdqQ1xKdEAQ7BBQYaO3c+XD
8hG+2SZCNqjXny3QL9SxGEJHHCJ5cyNhRF1mCFT2126xzZOTem4jRVpaLqSsxP7C
7zS2kU60idA465qW/r/sDVzI5BazoscNCBMOxmr5OWVICWp/sVinlRfjin8tB7vQ
QrD32onxcHgWYgYwC1poTOjUcf/CXsL06s/L3CwYFDK+glUgQp1Ibu5aCJ71SzdL
5KxsON6EQLgiX03ATUhVbX/+s1VvC175a2pn6zYay64LsfyAy6rM15LE546JHd5t
9/7PScXCT0MkNtJ5mw3YNOKsF+9KH26i4SCmoP00IyPCNmkf9r/8nRnZ7cr/pB2d
U8Vm9EMxpe3bZ7//oWlzQI1zis2neeQVcEHB3ULxgxe3N58vR+65Agq9yqIfdQJr
2Kdu0ydMWobWK0iybGxuMXvY2eFNKUE1nH8lIhJbXZWAkYToYnm82vxiSp4IT2Wp
D1jlV4B/ufIkCqEEFh9aakY87y08sN1/ghKueotGENisBXTljJoLD+7o4ga4JshW
y+LX4p3hhKBWJZkP0Le+pi6stgMhcPIUGIFGjwpNxIRlmsdNUBiITtGc/smZz1ZM
x3AR0eovjXqR08a/uJIafoFWceVhLokZ8dt/wl+j7/f0tLOSQKS+OxD7hEYWIcnE
aAH6GSoS4WRp6StAY8gHK+54Vvn/TbyJ8caHi0F9rcM05TI/N6nXMOLwZkw9JRtG
GQV+pTwMEyvkZVaYw0FiZHlGyhHHoXyNJgj65gUW5p5oEYsmDyy6wff4s/Sdqa31
G7aylwYc86LKvLgse8mjKnEzLBUJAexEuQW8jWVWBUmpk59zKvQm82Bw0UkxOz85
MlpWuOW1XCiqwhntTiMSczJXNH4my+RG5bXU9wDBaEz4C/3wtGR9Xl71OVvu5UiK
7fOc2ciDzZfmfRnYtCNqZmfsPjVXIIynjLpC3Wd6qr/7bieLj6Qh9PHH+11OFrYM
E8xYWQ27M4Zrtul1fSKU+mX601WGpIuOjj4zR5PaVLvH/sJNQ/KPBi0MQPJoZZiT
m+UrUfFYFKBo2M8bE2pOc05GtVwQUl6g5qVwra1DMp80dxrJnCNYLHgwj3NsWKuo
JutkQzNGdP3hVq2Nsos68MKrfVSsyOGtefm0k5q3CeqP4ueUJ9V9HVR2bjNsJD/N
KjFaV3NJuFRr2s+S6Sa+SVoB+aZxzGookrT+x4uEcQ4mowRpFx8iXXsi2JOozQU3
6/RFyqbmZbiQmLGJtcdnsMGVhb09OweebeeYlajHB2LJZ79WQnpH1+zWPvCSvqPy
3mOgqQ2ntvwhbvz6r0kDbw+ReQkbNXUVnjM9Z90JgJ4s2dg2ujirBKEX8Tduc1vn
g4GOpBxa4ooYM7/69Y+sQQPAugdn2JXNMJOTJoLJRFuLRXKor7Smtauwr+JNIttv
Cy1LU5qiw3l9C8USGg55s/QPb3UKax3Ri2bpkJpxYy0kOu51reOa77PJWYvZKt2X
4Cr9ZKZFdccknMqKlP0k9Tfb3SYpTPZ9udnJa25gSFy0aY+jGYXcigTiU0Q83VzZ
3nkhTwlvgzbzjMlKnI+vhmhG7VYg/jQcKDDZ45wGjjxPmPxnX1MgJ3+Jq3w+FGhh
TVq8b1SWcPj9kn0kAgpKtYTfqf2nmudBMxRQ3/NGLszc4Fk1e6zlS1CBAiF40h5C
Q0/2g+WNYTcSO/2WBDEh++3FRlZoOELr7iKqdi4IKyxFQI3/DTpX477nuP4b+5i4
dIRS/gQsFR85q9kRDbfLY+uPTWXLj07WRr4YWKsXRfftK3r3MHLrZ8dbdpUhZuR1
nCUJzCU6bVXWsNz6LJNU0WJevxAvPWZDp3wo7JUMEFJwMEjXYdDwmkZpBu0o+V31
WAQ0Pq1D57yNQ5bOILSRujvgsmiBg4F3z849OHNzpqeOyjp5MBd4ahTjj4yg3hXp
pT9LYNc0d8s7vdUUs6JIwS+5Vlq9Gb0XEdQgSZFcMQGbLyABA1PI9mEuv2ChhK7P
z5gEIfrKo3G3czLe7uZBwB6qbdKZf6gJMZ4BNvOkOKes9LKBpyEPTMSa2BkIZv1s
dCDV9xAnL8HoWhJb1jTYaMHTG7ejSYSthzVsCXj7TBmdL6Zy8xEn+Rsd64dzsSAc
RGkqg68H7ZWVAINPEd48N69FMFzmd7SwBfssBX07ZxgElt2XQHtbxepjN23eGR0q
vWk+FiIb7nPEQhQTiiEIPG7oxDkSVJ5Tt58q4F2k59cdiwWNl0/Sgpl6u7vAAX+a
yt/KBGuPncksRdwqZgiw3W1rFnHQImPnwaBPh30CoiOobRyAV052fJCr20FX/joB
dQXFPHuCJyc+81ehG4dwTGHTgSweNC13UhaPjY1XRcyoKfH+0OVUWnzeEaemhw9w
G0QExw5LvI6QOzGfsvip9ixBIhyMLlXQFeybvHNdwXVyotdTFXrfNZ0687k24Zdh
9stsgaCAxSJsVrNkt/ysy1Y28qoKvKB9is065BN48ZKE23y/hi4nyyB5OY6lHttb
gKxCazsXv1b78g4zyZuDdzJa7WUK3Br16kgQoN020vnp/zsSsoQj7iKuKlCgW3N3
TaPVYCAFdPkBsDcUwsMJOgYFrntksv+Ybw8uE0/wEvhj5+U6a+5cSqErBwTaKnJK
9bClJLOldS1+xP/KNZ1IyMPSCXyEBGxt1HFzQYcjcm5nKdxnSvyA0YkJ0lSwzam6
XjWAPg4PRuf1WnOprrtITotxUG/KW67XOMNF4ORJ0HFxQ/vFRcgC01aUqHW4FAtf
zT4fOQCcPHdUbBFaLayElyUMvN66wYrXCGXFQbTmPc3gjEfjsuaoJuPHfihVtwQz
5ES8okfsTI8e152kDlbQqQbNQxGNvXtqjJWvDOEKsjgYTJczvbCFJlioPXNAaRBq
gu5dt6BsBI/12RoiF7rS55Ogqi+641BHJ24kj/y6yZkeilDCBRpWjCCzodyIoQYw
l16oV0zDrrpJexcAeZI7eWhSkNTS+8ZqUyLB6GL7vaayfwbPRxiWF1bimWLkjvbz
pVbM3T1dMbRByHtM2Ws4PMz/Nl1zWkjv4bmh13HN0AKSrTqRUZhHMEMNjTaZP5NV
QheedTVDkjKAUP9Tq1qDeFGE2fee6fqbt4B0ooxZfcIaxDa0IE26CQ5ZHInv4v+d
Qw7+AzABmoy4IEIMQ6CumsiEMHiXkW5HyfJWC8NUt+Ftre0QT8fzPCoOmBIuZLVx
2eciYS6hO2+fzZnrK3rDVOi5olEH1PMtVnfVBgb4fbYf+ljUSVxpmgZgVnnUgrCo
V2v1GPDvmpp2NhOGRGT53eziPK0yXLPln/jH709g86/4i2cfl7ms134xFTjXHD/4
JMm56K2Jb0QoBM5LYPsgMwEEfo3ftTbnVJRGcXL56Of/xqLBo5YY8hEbtXfETk0W
7fqFIBST0uFOcFqG9JA58nHjZ20cuB62bUoRTqZPRa6fZmd0lz7atwjx4TX++n3F
xWdNGiIDtXWOLk4eclN6CGbqsM+SwHl7KLV+j0Je6DXmQOk+AJpW5ZepMeto0/Ca
pWZ73BA81yInrAR0UecbZbWIk3MvcAxRqifAc7b4TQiQe2DI/pU421cwUASLYGFu
v4HyN6p3y2MhD+lnmfyjuu+10Oc68rGZPkqzMK+npDoGkPwzlGkjjN3fgA9iVOGq
g4VvEckXwUUPUtuPSVOpploqBaR8N2zUAS/5TZRBBuP3PN8gPYmQmSvMayDllSxq
kw7D3Mm2xYT8Zy9b3LpunFHCD4LBV5IHEMLpJqZZvGNyduUExNtJ7eVWhHrabruY
NQTxlAgch77d9x/QXhdW4/WxhBbqfqgRKMIywObo7MiRuBcJg9Fl0wiRfUCJeRul
7TMvlUtq5SGvDHonEqJwwj0MYHy2Pl46YSSBnZOYYeXUbcI1Y2P4B5OZYWqfddxk
2V5JpUKyI2Ae7vN8siO6UtzcJ5qhaxEje2j1SRcFkocWCvEZ90l9PUEsOzWjdxbN
IEHghBKiOjA2sN5O54AEb6CKL7qMidnjQb3QORBmysDOT28Iaqi2Jrtv3jybzBaw
EqP+cgchBEjgeMJOdI4rBzoTaJcwbfhEPFGapE/L4Whuy9hbP1I2ook0jnk9nUiX
KBK5T0dRb8ldaU89eAQmmqOPHtui5PKCYrfeI1+HFqwYYGijx6RkqXrXLoutMZ4F
P85gE4i9lTz/btKOeiZzr2MALMoywCKdaDs/D/oUrfLB00HrkOQEEZUGz0c23OfY
iYy4EnpTmvD2Y9oNM9P/EUOJhTcgxsJHOf1INYL7Ng8TA55oXyyWG1T21F3F+bXX
ima4xb9qtk1yXjHzDbwCMJU9v6E/l0NIbhLoEJXn6lsVCWStL6YHScK+k23df+Fg
OxvPyhR4nDOL43MGq46cUFGN64ga68i7I/wlmzNTmHlzMC6vVephQxbtzsv+pwdh
Jibh+maurnFKpqlqTXCEwRWGzZXz4rnO++qO5TVOphAQ+yHt7cbE1W5Fjo84bOuN
zOTX8URtrBSJQgLw9oeSldJZ3tj/0xd8bZqkDciPdQ94RrubsqOB71Z/M0s82hY/
ZTy6UzBYN2ecKmSvMqwRXG3p0GfMEqRB4ff+7tB29yedZsuJ1oV9Y87y+/P3lbnV
9nkDnmQK4CuPZ4ojJhNkfLRMIpF4PCrr9Px5zdJ3YKq/hrEzUTKzXIFeYZJdjCVJ
W7GhsSiRem32sV0c8EvOiBur7AC7pGtWBRzeVXeiRFX58UCAjQ1qC3lNPhJRdJ8f
NPeRp08fBW+XgUHHAoRjTWYjpMNLNO3hLrgFF2slBtMo/wmYpDHRzc0u/6G/BW69
O/qogZO01cLwi7icj4DvThtAWfCTNJdYSwegX2cyZuYxIrTBONcyS+KqluuH24/5
5evbAIoOpReqa7qZJZuZZqnTkF+j0AvRF/O6PLwHjti0PYRJyrwQzVQe8g3UXEyu
D4DWcL6ViFMIXJgbNKNPCKwWT920oyRvME5hfXDTh5Lt60W5YqExOaVOSlUjWn5r
+Ibf3trBXUZOKW+77t3EmzZk/IkBYoMP8FjqKvQ+o+fxmqeKn8XmW60xiYtAsKEC
OGd91FKx3Jb0n5QZQlL2MIveP3iZI1+oits6tJU3y2Fut/sSnSNjP81F0/YnzlDz
euYxO2xvE26lj8Uyw+52fT4Wvk+9bWNa6B9VO495BFZFOTwatZ81Emu2PLIic7p2
azKScy/wsfqzmv3dq5Q9ns1vfHomLQziuzBftA5Zp9NWJIrTYO9y1LJQ8HIA8GyV
uCrS/pZVIR51+t3Xd5d85X2oRFsZQnocR8ZYIibHCs3+h/TVB5GCmqSbAlTE/2lr
aBaLF5V2Nr1sVCovC9jTWtQJRSDlprsAUQd4N9NMecrGr8i0bO7Eh154P0x3yikJ
QMYahRSTxutiK0eXubNePOcc4V9+KIMl7fSHoi7v5O1nywvIhLc6R1yf2VOoLYI6
Q4SVYxHm1B7+JfVr/vcRqXZPibE1FOyN5pIxM1pN3d7YuTsXZkj9dzSVP0QbohZ/
TnPK/GWUcVfMXrtZBAh36MBULVmqVbIqjAVpr53GShBQA/wEYtJAEp7BoKPxH8GS
3d+PLUZi7Fj/bqqdl74ko38ilvbp2L2BBUArCz+cNl82ZbXuAT60FUa3Zmzhtigc
7kVSuEX2QRHO+Mdg106PdxPjpnpuUjCr931hd1jKPJSxxGPL5/Mo3SglTXFozuVY
+PUp4gbQmR/He4n1GuG/HWRl2fSVvUI95Pdizc+HWrjCNBPGwGbVuyNALeG3crQ3
zcklvSf7qECXMkoR/WMqV7Pb0RcJ6uDsdCLW5aHTk51Fciq1p25C2p37r4XVH2us
nEYr2kJo6ZmKC3yr3UufGcJe94f8v/RNUbJKhvn0aWLvhLnVP+assAsb+zse127P
s+xb7an/hq3slCmNYVlbZdxLd6Z0W6QBvI7W5QOFjpr/HPbOBigIEBpHL9BmFqsP
6qdcub64l+aisi+QANUHIvLyOG5ckNNatYF+1MPOfKyni+nwFmxXeusgjrmO+dfd
fgRwHwkeYU2iQEeGgMUJx/NSCEmAiq5CTo+aVZ7Z0zjw837gWQA0URQ5aZkaZYgF
oRzx0hjOkBQAjEKNKBSpBuX86PtOWrLL0qVrsEIjXgpSbtMs/JmpuZPL2wqqblVJ
ZOe1WWxkMULPthMdHb6lfCezEhREGZCpaq6LosZaLfWr3TIa7woS1RbF1EQEYvOn
T8z0CPhuqb0qAiqyeSAqNr0M6M/Nxso6EC4pbuLGwJSEJcjkk8RnqVNwU9UGUGME
vGqux1nnXPuJdwcofJ3fs6o9Tkw1QQzj0SYpYayfzRxeiUJuh4JY6GnWgkJJhIQj
tjvt4snX4JpVxq1z4RPgtqqRDTbFqtrMb7rfUBkx07Vp8wvzAEenOSH5w4oVfuO/
AVan0SVYxSfNofXH8/mu8nXwWOrPF/tiQLccUf9RW+kQNai76dEIFSlIQfbmpY9g
5B6mu2+FcQv+FCbC4H2ngJNyRHrXhCdjGaLk1LZueoYm93/jNsne/4ZrmxjBqzDM
SvJAZCLF93Ln8/pg2VCCdE6PJeQDZeS7iTnI6Z6MJl4etYHcWgeUysKmSLLzGovC
rogInp+QaniVheDE3oDZWzzNUewl/6aN+0wMKcrM5YxLVABVU6sc148/gvXRMSMt
dmsSTLQI36k6sjnjwwI9k/2o4i2u1PB1t1HYJKOUczLtxCY5nscsibIXDOTvuKko
60CUZykJjj5AzDv3H14NFfMccRvV0lmyPUF3VJcq2JZwmcZCcW9BSU3AqgadtDnO
s5JCSsQW2SNlpuLcvm4uYcbkH3ericOBxu3QFpLGp3d3g5/8FsO912WTYKJ9KLEZ
gkm6hDCovHMKNBvbUsZaCHgBVnMDfad53RE2NPyGl7LBi2O17MP9MJJygkuIbr3G
b8EvZX47FRYl4XVC/pr2U82P4VS0r3vNoc/6kORMw6MWw5ijpGJgPNVqNynEkzqj
HqT6Af0oQQpIzj7B4pQnhonPw66KQgXWuobOqFfELRoW0bKBmoVErK2oXw9nqKS4
DtwXd2uo/G0rWMuJRID7+M1EC+3bukHG42DUHAFLCZnQZqNpFwTNJ98FcESUD6cx
Z2AcbEPbm+DSjn1DlBWNakBL0Ai0YJ1Nd+z2ub1Aer+Dsa84D+E5CsVr0XMFULp5
MwwxkkA8YeCvkO9HCvmMY0Q8S/5ZdduhXKBXq2TbU8Ukz7NWXYNyAE0qhXGOqgy+
Zb0dhxMQghOvRU5diadrXMGwmvfsmfbaWNfk3qdSQbGHlqAZ9qGU1Yw3qCHC3GPt
M8ou0g2k7ZDe1ibFLWnFIJJRF3XNiiklK9q84DeU+2pdrB/RgYGyz+dT2u5v1P6+
8RQ8d1fQzshf4VPQj+JXoN/fwcKMC7hjEP1JXE9bVsv7RqOm0AG1r8tRQ8hs9Dqp
f7/sTpmOm4np5X5UFRiQ1K8rGDbDFMRALHxXDS20RSiIi0YCNYWU0Y9uGdu6ROvH
hKxk6XtjQG9FKZl7rUYYJ85/P17UJIAG7LI3+lxpp3k9hKElXxN45lXADQvyKkDl
kmyesJapAsiSMSw5YZlFazwL6q0XjHZJAngIFD4XZOIQf+LRxLmoAceiOZoZE3f7
39ONtQhm2brzeZZk4l274R9yNLhM4/XyO2yq3NiAv0KP2GPlkc+DhhbIseN8EfcF
qUtBxP7BfgllIuLwzY84CLD38mTH239wNvLd7MY+vRQqJhz24QfDNGidamh2goWn
7glIZJAuacYtDaWHeTP7A3AVF7jaJ+T8QZuUoyqmQZEaDXWjmWDzYyv4Z3UO582O
NAhnBaGoM8VJH5TOt5ZChVFr9+yP4LHdiVgHulp6GTa2NnVDdbge/dgWvGK0y9Oh
am0VQbi7HLW2CR7CSGXaqPeVa7z8s0sp2duhLsJKbQFqEURpSTte3kzn+NTHyqpB
3tUNEWBLEdeRbc2tE3mJCET/pTP/lUEES/ewmZXucQGx35pd4OK18vW61NCpt2ju
DOuza6N2zQpSH5TBDdkIkfDwqvZvM7Ynj7eKIu2+xq1jZPYmQGf3toF1uz4TlIB6
lPXeJYNjL3GqWmIdPgaM3RTmUslk1XNBdAyEhj3awNZHRrPG7LkPxT9/9hJ5rvRj
3K/4AoFJ5it92eGfHwVZlAyjfZDYJNSeHSfdercpKECNOzZpaf7PBAwx+ayRG4c1
vI6PlBaLmO6ZcpetfaRRgbUVbeZStfudc7AkEUbDX8BpxO499smkL/byBi4ShYj+
vZB9gjxMqxOJacjgkVoGemS/2S1fTXhRzKIZ/EtxJRsz81HFMZKRhpBMGI8Q3PFt
eF4mh3L5ZjF0r5m8Y5aSj+n3Zs+Z+aTfeVLkqM92iTUC4FyfjlJzNdw3THM0O1ao
qg3kkzfIVKkWSh/5DMIZGhQ3pbVBGITK3lM6V88rMF9sc5mKAIaKXBvS+RZZcgNE
7NwCrGLGXKcn39YvTQiBZu6BB7nOCdOrk3cIykuhggwLoMHFFbHfKBo06GWex+pG
YEYvmC4APRwa9JlDYUYGVutIdBXlxTOEZZUk3PJt0R223eLR44MQTyN0HeuXUfE0
r+8qSvTRiK3pTeYkwKPBrrL4DckpnZtqbQYxOCOPu9jUjTgf58QLBGIvuEGUdPPf
pw/H9u8loJ7Q3WvFdOYuDE0e5BuWLoRnpnPAlw/+5Ak619pys0D8H8ewFJOnEabL
pxkfoYi54Xtt879cbtOR0BkwkSzYSKClCNOmx/vn9/QhW8TbFdq3n6IPiBzPfNah
z3RV8QI2qNoxWm9lY+8sLNOkdrT9b782NG4mw0SjlzSYY0l2IVTyivxqAso1OhN8
vs4ekGNl2Mc1j8dmllVtQPtRJI7uy5+dMWRaC+VkMhKml3qXd4MINlObuIeOpIN0
KEOeQW0H78cC5KX6hlfpQrAezhgaoKRoFsJLmEVil8cOeR7oVIJWdTWvTQAv39hF
VrQmcWhaw0wBFIwUps9O71pyCzMH6UZrPX4Zn2lXgEdupjocWgHY2p9XxiVHEanF
G+A8F8D0SO0bbI6JU/YfhKPWLnDuV1m2GuKcJj5GmFyvyaFdfQ1USFZx3Rri/3Wn
7vQx4UWCv1Nnd+oz7LJBn7nGBXDAxvBdeu1vD8t6kNsptziZN1kc0iqPLhHDaZSd
v9+XFgVaH6+pPd+Hjw+Hd8JXJODg9d6232CtUCDFex4pGpdPUF+HdCdCf6quEICN
8cLa8HbJz5CmiaUeeZxO1JOE9jPQsTyvpCfdBnzkilHJXHkvZgJ4n5jGKe83u5L9
KeLh3hOoIf/j1jPpN1p2YLbVeq6RStAXAgS66428Txgof60aRqIToVwEC4Luqach
DXwsIskl+6uYVQyeeGnoFO0N6safLmPS0UkSKfFZtLbPSuG7O8OeRIQiXJRxCcV/
Fov2RjmogkwKoyZegDcmLCdEFwQupOYeM3t7hlobYFfxM/GRTZw4fI627dRCxzA6
K+8HCWbuFyMTucMaGP7wxLfb4gzEhdXJDatRL5OF70TvV0bogxD0n/vyKPAVfUKH
bdBPvRHlLdhIZHuT8/2dK2RxglYAIz43YMQ9+9KjlvlVtFQLtRzZ8H0XIirihByo
2I7zGl5SJv7IJYPJZiUs7NfDH8uuwWj/97yiLEnoYTLcQ1thU2n8wbLiiGOpCe5t
PU+xPm9vPkdm5gjlc5Scb0MwyQz6pY92CCULkspCYe2lLL8m2fCWtf2OOpg4X2y+
4USqquult+Y4tvB7/rbL1yUryljXfxU0c09kd+AzIdVrEyjbPrc1YT7YZN4b1cSw
J6IhgxDnU5V+TDYscCtLtHCGI/wiyGPzLYCqMOWDx5UNJVvXGaQnPefh+uoVd8SM
625sQ15vahbDgeAFeSXu/x+wO8S/KS90Xow/uyfhVAmNrEXWULvyJFgoCiT/AV36
uaZtS4LVlfZS1TrBrdmsXBQUzzNXgBO9JvprgvSbApv6abaSfmKgFfQXtQORGu1i
oSCN8OrICZe5ORBxyOv7i9jtQDxyF65yuvoCVRVlJJ9wFdH6VzBmRv2ldxa1lpOL
p2dOQ0q4GxpTVprfttpby21MAU2mnBht+y4R4S36agoV9EalaPklngA/otXsAjls
mxYxSFpzos7sRRZ4/4OP251MgWn3hp61qpjkBQcf+aACRyz12RX4jDI6g9aGtZI8
Gh4BZlpKharhRvTV5Fpx3N1qJfjd+wF8UxWXjikCmmQimljdiYVA3i7AZkA8kbmt
NSr3kHNc+kOsnBSqc4Cql+uqKAYiNqXKcSTiPNdpVNseZB9KzVOeE0aZGqMIKn4V
ttk4TD9qd2DyDpD4VDd24cpOxO4RHlPyxhSrbBg7hhuNv7/iXoHVNzv6GRvRuQoa
eulA/96SWza7LsJ/RdQs2pjzFtXnGmqRAH8wjFHUVWykniE2MDiveMML3EYNEFDv
6yTmX3hxpqap2YHehd6GGsf1n/qgKpfC7nEazurgbgVioXgVA72ZZJisTBGrJ2vn
F5ma0l3Qhx28//sBEQiRtE92gkbX7ZoIuvGDn2XfCq2ojUnq0OxvjXYmOvEDaKGE
ONWO6YVZZZgYRuf1gjz5tSQhTXm2QybAoM8XubTO6AIXQIyGQt2+iiZeXtJYzOj7
V7QmBZAkXAggKGiQ+r28ZLz1Wojc0DSM63NCPxR47wPmyZzxiOyF7E3Z0h4Tar6Z
xwNyDyNdVHPV96+70RLJXCgvD3sJp2WJa6wusUp9Bq0wDYZFxw9ZtrtMC/nkfyrQ
WLq9A2J5+1o1YRkFmg91SfguIYFLSGed1odhnJOhhXQoYTOYlxvq1p7v0Dws58f2
2qgf2sqhVYk7U5Y/CTtGzeVB8sQsij2/pxl8tDSjQuesb4O2Z+piUxHK+i75Q/kc
C94L7o1PmapL9QiJT596tgPyLXskqoZ8tRjKX7d/UQPVeHXVws0+umE/KAsjRQWU
W7UmaQDZ6yJDZNj+YaqomZgCuUw3QhBr/klXy4M9kiLgPzVKDaLsB+a7HHcVetrZ
k+nYc9U76lq5Cpo7H/Vj2ZlofMhNebIGOb41LHh3iq6m2nQkAWWRGrW0m914siJQ
OSx4z4BrhmER1v+8CpniN1KXaSEBZOn0Vou+K4WbbKhzqSF0nUczdosz6P6uuEeN
H9fsYQpJ8TkqnqhtUduATsqxBm3T5MXbV4Nlf+gJfo5mNU/nFnPvKsN6T4A2+WAQ
JRjmRRweYhXzTNEluMOBwAYHMtHb0XhSBhvUk5KxFMc7jLcAqVwcDTIsM/P8qpmD
u+Jdrc3PB55N+5rKt3p7ezzc3AfO+D13xzsC39KzlEc/tfyNDlpcDRZTrhtr53Eo
PUm8NQS/5NpU+jq/LTByXetVAE6z/+XHdxGYoOLHecd0czk1Cggrjh0D9KClQlPv
RdVw//iLbVe1GlxCXcqPNQAHwCWDdyWECkWpdHsuxUJog8gJSyMfRPWMIjRJ/tf4
sd35xaZSW4oDZNal90tbJbN/k5PZIoFXKUrWBV54Bj/HspIJtaSvY0ia2B+EcyUd
oIyM5wfA3zqepBMo/0UrBnloAU0f74y19LJVh7QdHlROh+3gpU+wDk1k7MNgrLxz
140yZiAb4XoEXkampcGh0sCJ5rjU+rS7Q8E6hp6LPcTaG3I1cNaZzIoEV1RhLQXr
c0UAnT8gterEPgEz1YLZQ9GplUTSQJH1ZVgw6oL+ZVlUPz60CWt73kQioLHf4ea9
AurR8l/7H6u7RYiKc8hREHCSwzqO2Xo0u6siGFLes0remYbN8Z3g5rslF12+WnbH
oyqvd7Lp+RsLxDl1A3lBRbTprtWzjAXUQBXt7jaxhmAu7FH9zmBlE6xK9DqbrePJ
wOC9RvqftS0VN/wxmNZ33j4NM3G3VEnba9sDwOfw8Sa/ehJrymfF7IkVCykvR70I
uSGmDFh5TJqIu1w0UnU2AIGug5cHi8oMG0D9RFxDzuOP81m1y0ct4JttzzB/kqH4
nRcFYvR8IxyG3BA6RX12UwEPiNAxNVL5sfyV8e27HUHxGwSLgG9GaUbtvMMDk1MF
OGL+YhbACU262Yw+WVjCzlm2bNEuhlDA0km7+YWUvUkwBEbe+VDTr4+Wr74ed2em
53WlpB1S5FXHyhFAQSDzu+G0+heKsywuEYYIPalFbmVyCZJje1rU/JyhS1BH96Fv
T6yO/yTyMPpbkH5BjYYUF7pVLRs+7RsY1plHGOxz2ZOIQQO6MPX19qa8IWYq3Vpk
yM5zmq6JRthYGcVH0Y7qBF65LFtXE7aJGYV+AFeOzd4vGPmOmpaibi1SeeDnQ9o8
UQyzoDonNPvjeFhSc1QDBN575PZ/yuZzVNOqgP0Yt1jT21V4pM2jk5xX0SDAIiK/
FtNYvZVlwkoa+fuvSoQWQYDJRWi3fhzDWeryWjVj1C/QIEaQUZq0m6tN2eVB7UCQ
+MRdh5/gW4OzHf0i8akFv7YBs1nGjcv5cAxHChpSgDD5mKvk6ohlDdTIW/nK6VLn
tU41WkyCK785iJbBpZd+oJyLgfXtfLmGqyMlN3SW4rMLvYL9ym2I+5ysRv74lqzf
cTMSe2JRjDnrEkduGELdxAHBZWsFCmu4tAs2t4ByYpDygAD554/odh5EKWWzd/z4
AY/R4WwNuuHcXopWPKsabuWW4sxojnExmpIJTNPcujEUh3aaSr4lBPku/FJE2XfI
/GbgRP4DXyx6y2W+4dEU9a/wNf6/i2xcuF24i7tdeHe2yaPSBUAYli/cOuFejfwm
H093UsjofOWb/4ipQnFF7H3wRFgqM3SIOi0l3S1l7gMjl2sW2F7O0TwTG4GRTObK
VeXdUrdqnnCCSeR+KW1MamJzgDpd5n30dvKt2FslM2s0tt04FEivG4/CWIM+jLob
PwKDvAGLCaxiilkvNCVAKG9Z+bGxx+D8W+p0QtdbnmJ3JNNviy5mc1oS2fee/hpO
3ufknzazuj2S4w0c5RWYljkgmdre9u8OrKPb1UDYvtpL/iGszcqA56v14zGFzmIV
m+1mrKhGuHRFuRX/aSxjJIFZ+RRjTICkOhFvGxT1GVKor/nXE0n0Shd2lcHh3FtJ
QrAXtYIzPfuQu8gzgiETnR2mxUnqb7p80e+5rqSgBey0ZNS73nE4GNrrOpbtMOf8
27r/97xUtC8whUWue/I3D7rD+dmWfIrKRCdALf2aDg3ry/sXSzG6Li8PQVSy1f84
d56lJxJsNcqLWRJs366LE6DyvGaRxFyJta/kHJ7/5pyp4VIig/GL9PG+ZhTG/4Lw
oMD8GLn4FXbYXdDyX4aeXf2Hy17u5T9TbHcdZbwSD5mqsm8AdGUSsW5cNW/reRsX
ByPaRKOnPZTqasSKkK5JJVGH2jLP1cQxh2PRqmyf0zlJ0FPeV62LI/C4YJLjrzZP
mZZOa6vxYhl5Up5Yit4HXuB+yeHr0uSNdIbxBcIuJpS/2Tg9AZDEAPP/ItDT4TsY
B6u1NVqs2U2xmW60iNflhDsAvtBX34DB0HqN2OwlcdLyT3g/8dV/yZBlEGcPMuR7
Ueoz8wCKCJxysCDsf/bymMpSbwZMewmijE9hOEvBjW/a0jeOAfF3qQRPL36BjfI9
nAcc1nloA4skFJsO1oV7u5Uqyh+SPiRx2YK3js30HMFwZifG3BHqLu1/HSFbJqX8
JTPu0uWU/7+r1RMDu4jgkCFsE+6wIYjEbVmtR9rc1sH3IdOi6jN7NsiUU/bh4Oe0
tAWzdpgwKZldHhB1cnbGKWsaV/08BAeyioF6NTaZ+Mk3jlSczX+eyuJMB8cDp1G3
0j10LTMTJrf0LUlXBw0Mtwe64+PzlRkjF+XMUl0E2/HPbIPDRnXPmsaIY5eYkPRs
ITZR9tYmRMZj5OG9Rn4IYO/Dujz41qsXpC0zuBgdHAoAD1QVClmrSZzzSymfsGIN
3HVVh2KGD6lQVftH0acfiDF6PlZp0y1ZXKOpUO+y0knscEnEYS3BKGz7RP5TWAsQ
y3PoaRdvKorY01Its2U8qoI5cVTXW2Ovctnvmq5LvI7HvrYAZ1b8sutujZ3N2pgy
XZEx6ZwvaTs8aWe427dXlS8OrWh1ume4ZFoYKe9RYXHY24uFM5scwb9baB4+pjGa
R/Egv9qSBzOkl+OIyVYT3pRdLwbnbUR4aNpZ6Junrk2u1zXsaYSRku6ZR26n3LDG
ZhSsiPAJ4mQ3ICKTJAXndREYLGXHEV9P0vgIJqUFvdFXTinpCfE9njO9CAQnN/oz
jcY5KFofYsgfXKoCi1TzMqhhZwMZTLANlPkIRk26IgRMsqSYxjwfpYH9AEjNPuU+
R1ahUazxCmcVwfQsKriy22mRPTjYNyyYRSWSEV5kYmJ6Jw+lfh9yPU/3GInL+VU+
MmsLO0Xa9ZCWqXbsZv8fKjJK93+zUStL8QIhk8AJK+XcEd5u4IwoHuCawpetoOtu
gZ2mPRI/dlfq+bVJGOluz/uB6tEMxB+LPzv474jLGAaK6jMRXJA+I5UQy2B/7FoO
7U4MXd1MjGYvJcuIw8NtoG6/qSGILgcRs/m6pczSFM78tBhZ3xn2Zslvj7kq2cNT
bhVxaYmZDYRMRA4Gc3h7l176LSXPOZS5jVZiZlMYg75Sp/GB8lOFjyLuC3PXn69R
w0NG6nYSMSAgVbHjMtlXcN3//eJ9uH5u9/Th6E+BVmy7Q92Fh6EwpxYcS+5M9kXj
j4dpYYL0IEahAyAjIErbqe+yhEUKPvjIJOEnSL5PSHRx/BH4nCfc1aqzuk1lvQ6I
HqJxJ23ZWYQ112Y7ZmkJ2lQffrIQBeS2MO9BXwfl63AtSzRcuQnwHfg5Lsii1BMm
jtt0UCi+9sTCLyprzcYJHsrTsB7PVyk9BjVLQOQB2fyd84xZ6Og4a1GbQNJPMIic
oMsIVR2ApM7oaE2qgL94VUBYvalKuaypW8BMwtEwVtZrtBbnqRERAQm4c7nCh+Hh
KIjRuUwUgJpyLsXmhvRIlk2RqBLrLmIjggpQ+HDyYkkOHkJiUT+OV3eBnSdgEcau
uTWVIn53Zbp32nzqvEqYj7ujmc+ap/rodcb5hfnM5Dn8GCCg2k++8MPQcZbqgPh7
pivxRBVtLcl9s8TEzCj6/FwBY6AY/Xd+i7Ov1AoYZytL8/eVcIgGJ8wUpHAQ92QV
pNoU6iwJUJuwFv3e/lqMuhznoB0tRnoRMDO3CPwSLDTggYTaivL1U00oZgzPXwbk
DQ0qug1mWzM+reHl35VGHYb2AXt0TN+/GzVvTns73PvnBLYfNBnVZxkITuL7+xVS
BZc675EZ5XN4e9VAyQXYclQPvUENoByih06rOIuE0hKnFPdTBM8M1peUAcNx3+HV
ydry0ff7yk6n5U7Fl5b4JgrAe0NwC84BXvXEo5p3mVw6PxT9+CHg/Bg0jpARaTcm
up5NVQEIkj24bTlp0RA1mkqsVtpReNHYn4xHpzpj7MLWZiJNrxG2DjbJm0+PTVLp
z+MY4i/ZP4/+bljLPfBJBQ51uuymUzciJKnGxptCHZDWbvh8up11RzefLm9+yDun
q60C7kUhjWemwJ4EVf5hqDTzwwfzMyMMt1A9EOEcPN0Bps/EWyFLk521Miu5S+zD
D9aoObaOA3ynSVCp9TA3nz1IHa3tkfrfDgZMl8u2hYn3uRYx/bBZ4Im4tCch1Ral
1rMngEt81ott/+TAQ2lTxtuEIeg492un9PG5sfdRNqGEXBMg+gjjcUQMeV2EhDmf
qSIrXERvrrFZuM1vWwGCAhqlA1nV4QLy18YxH0TpKnMckDzFJQnvg+IvJ/Yb+wbf
HwOTuxT9qbKw/6pNa47jxWqSTc4Vhf9hql2FGe1ZRV5LU7Rl4n2rQXJcLMel4oP/
bOXxMb9PaJjuO1ZCOWJdq5HIQCOXp6ukQC0pDiaB09Zn50GwTgG+5VlLzLy3+N65
9uz7H6aRNA2IPc+BafOOjo6BIfpSrhO8JnrF/ld5rSYYj/puwKpYdsCXvqBHB+cw
864AnrcquO4++2yvNv+cGxrQjfc65K8RyK73vNPaL2DTZ0RRzMGst6ctxQjHsn5F
4rcliiV3L/RyHhr8rWs5EYktiXtj/JZJhC/9IEgzDA0LluPEIIXguAv/CENTg6dC
OEew1Rply3meMlmzmHD1Ty1HgDi7SXzNHTzJ+j2YQvc7n0540SVVHxX6xgoSgo2S
3fanU8iP5hRmoya2YGUz1MteqBCCpguGFTjeaCrN0+T5y+HNvfyJDphs8o9bybQ/
tlOkiZdgEwTExQZ/FkYyvB2qRPR3WYzav+EFgyf7iE+rxZJE9xAH9/4zlaZ42W+e
L6y16oBo1KOt12MXAuse0bcmeUf7ypEwX6gPqcEuJQEdSRJcxw3fl+LkY/O6HgK6
iazc7xJqebXYEpBJ5wysVkxoTIz0B3fEB4S9nMYfhEjgSxxbs+HlL4u21BywWRoR
YzZBC7ygu26uRa4k7HETdr1j1HZ30PDoPP4PX6SEAUmVQrFN6Zfnm4fe/k2K4bbJ
j4KtUYBY5DQ90HXUFz7AK87/VmniC4GN0lyo+AUiyl2eAjxByYR9PgZULNcXvNgG
lkoQwYutPzbLcC26fZo5f6XfHRPSHFr3UuD/iXAEizDmJzK3sloNsj+7V66XP+ey
+4+S4apfBKu1zGMl19BujY0AEP4bMrQ2WZoJs5ylX1GdaLUkfJfdxoAiktYCUQ2G
Bshy6gQhJqyt5ORclncQU/TW5KAbzPo7fCy5gfcmuzuTrqitzp26YNGgPAreMyk/
NB4BwPGdyJU0s6XGfTUKClpEHpTKLa1WNublaVzsvz9l1kEJh7Lp2O1UKnJFDm9L
Jfi7LBrhuhAARN8u0H624X37DtzV/HhaPmWPeJg0sT1IWx5A59KjjOLkyAmP3QuB
W3mC7Ssqe8IkngK9ehARCDthkNE1BwhOLrNcujg1ojQfsnNkeBrR7d6RxhxTJzSg
mE067XZJNPQIPdi9MK45oQJxODgxj4Xj96WvXzsMmKobVrLlDTvBmt1eVF4dbP6Z
mO1OtSjvu0qZZxp8ukfQ8KSDPJhKroujly3UmVR3Ctf2/vEtJhDh/BujpDzWvlBo
Dfos+8ka7paJPUQ/9Zpd6iM8i1lzfDxsMObBl9kA2HnDeMIDQkNFKQ36inhx5lXq
5/YLfIhY7qkb6Gq4t8Mzix3/42yvU8pgFGIEKg27HcGunwSnyT8SqOw9RKNYR8QU
HVut2mtedIerRzkmFAkPurJP/PR6uTUk6lNUlaiYXoJpn5vr3LaItb99X+VEoLUA
11CWdaQgUAxoBy/w27XjolPnLOT0C8nlZLPMG1XoxBGCjVURZAp6Cdc5DscBHj0J
q2IeoeVkG2KKHJz3YyMmu/Wx+hbaVCJzOUS6G0FjzSY98quWANvHFeKjZEfjRsA3
BDsv0xTAQjI3PS8hyag/djEVWuUnPcxX8llpsCd2ZT/ZL9gWbjnwX411uckq/w9p
wDAI5+Ny6uQ9E/1hZ0BKx03I9st4xsav+g7/JYxiEgLi9aw4YV0M7uerWbgmL25Y
o6yTA5h495MkiFNGVp/8q705G/IC+RFvqx4r9w4FHu8AeBiXbzOIY2NcLCC0h+pw
/+skze8o4dydu6nqLrplsb4XB0lfmTItZUSlx9KguONYp6WP9W+os+GiwpKzxSOI
3ahBKRWeNA9cvDZdXUtxtMAzTF7TAk1sa71zk5JFrAyZ1pU19f8oUdkVsvwbPTe6
CMMPVh7e/EvwEK8paBnMZr8rpt/aqN5JNzB6QWgcG3hw76QUpZqn552F8dheIIdr
WchlZRJLJyAN3sMWn4PawxceSbMEG7+X5k1AyrENMJ76acZeeRxeTJhuZVakC+bo
qAzrW6I34abVhVlV3G4p7DLd8ISawQginKf/NvPshiMtdwR+7l0lIxpEov6WR8ZZ
rHJP0/SJBrJCg1AaV4ezvIu7YSjnDQdmz++5gDaR2Gffw5RX+ofas3Qr2ClmCS09
FBHjo8SSL6BBNVjEuJFI02AoUy8RM1Qrnn3BdDi8eivP9ZfcaxhMfIv3G/IvrR8r
C2XnP6szXPdgY6kKm2nHGRJMUBtpkunGQ7dlS1RTDjR/kDNvdsE4ZR3V01p7TVZG
2A3w2NqYX5zM7KdCgnrbfFfLnX2BvJbhBTuyJzPfEb4kgERoWUQMzp40VCHeWo59
QMG9vCO5B2tb9iusr2CcJ+MWLEX1IPV104pkaInvTOUXwzcGH7lEcJNs1bw481JB
SaPVu63bMY8u+hvkAkyIvjqy5TFvwfduAz8ZfFJfpoIgnVTB2bV+BDwE7olhRK5Q
VfxmfbjHHB8GlCSdykTRs3RYJ6S6t1MrBpeR4ESu7N96EEN2e+ZaSw0iljAZABAt
DKzopY4u1r4qx/gVUAiQLrlQZQ4CefQkTYLPg25JUMt1jsYXIbwhttt4ueFBNHMC
7oMjpSX81o6+hMNQrV61QnjgbBySZ6OM8k9qyWnTezDl3FUtva7+V3BHz1G0zbcd
CfFDCcCrqAm/3vlsnZ9kQVPgE5jPLaOlviS4nGpAfow4Xm27pIdv4t5WWgZq0Ebg
jAkeuEda49MOAHARRycubBp6W4MNEAYA8pJmadoRFFMoukRJta4Vt943QXGI1ACd
XfMkBo0nFWzCGYSKgiAERxEEKo0En/bbukbTsiSwAI/Te/ClpVlwLb9zqDBHuh8O
JIct1QH+lU00yFvsSm1ra7XmqYvPCxmoV256M+fTjipPi+ftBLP5uGkrEoG+bA8p
4/e2MpX2VkXQ22h33z36bO8EktbD2PcPX4WMc9ehZHWwdM+iBAGjpSfDDX8kAudt
kFPtKYRAv4SYLxjVfk91VDFg2LW4YwfHk23DIfKEaobnBk3BAEn5pmwlZ0BeGt9U
YFh6BHQKl52NS+NGHjMy9thuhbInL5l5cGxA4ChNlQgPNVvdaycexaBwxrTAIY+T
eRQeQNCOA1J4snjwByNgoibMfG9NHIQ3NbUkWEuxYBS0SVLAljIeiINNF5g/C9Xb
lJrkeVg/rsoFVHsiiBi37J7MU2JT5zfQisPFnEV1HNcUTmZOYoDrDUD9tl6ggX77
vvaJCd7oNFnc+Kk7DvNH2tYrJLj4vHZ+gtHm2JzgVQipNTRz++lrK+cBxzsgy7xA
U3Wvqzb54TnjIwX6r6jJZXShd7ap9tGReJ8GFlI9o1StjSftjYv9prvEd/VHWzxv
KcXpADpub1EgM93PTvaKlkx0QGgAfWeptkTFl5JrH+kdh5cSlBOwIQobJcVGZQtp
44Ugb6pujmCPWCOd5RLjVnEcXccVibn9NpvoV2S7280/RagLYOLglpLuMgLvxJa0
qGxeIx4YKlF0TVVY/o8c79mLpU20W8scTbtq4u/XXtWTbP/bCe/dZ1htDgesZUGJ
Y2lf9qT93/IDax8irk5KjP9EobRHnImfP6O7JVIL5N2OTv2LBWGALV7HfsT6l1Nk
RhA1nXNhQV4r1jKP60UnLqEY2SYqrCB+rk4mVk226CuBjDH+UlzsVI5b6hMZqQnS
dzbvQpitZfv6KYDjdu/hzSqy0Ws2ag0FXDe993GZGLG0mm9C9WnPJLV5BDCb2F54
/jxx7Pc9QPPKPxz+wJnd6QLytdjtoGSwYPhRHbAziD+vZrzUIPeAsZqwKflIY/Tt
eiy6ORs6IYlpXi8ddP3NosccL7x749wJFR/eYd8z7VtDfDMicVc8v3f26YE0Dyws
JLqn6oX0gaaf0mLaxHHAojh1OJCigICipZBe/3TVQDRPSB6uDdq3Ua8Xc1sCFVmv
+JBb7pCpsNQThcyhP6HiXh9JLP8TkCsLgVgubqU9Zb2LavLdV/+tAOaUgYCwdyQt
fhitYD7i4ZfUB5K1yTdh/TH8InO9Fzw6h5x5iv77k8JQOr8jl5NA5HC2pL+V+aP1
tWrrckzkipktKOYfjjRpFm6tbLWEKLXF2ZaBObnDM9TWgjFG01SDQ2Lf+FE3s0yR
YYWjJ8dxXabScHBJgilbeFaYcfhEl6+Z/AuUpcyXpxYJb4CyMJ3ghK2v4zBcdi6e
9UUwCJegreEyjsLjj1t61Lhxt1jG0mJwMIClYRhlfb4JE0RKQxc3wmacZIJBfsxs
P84+q5027wmgNQFvACl/nDNV9WBoFSy+3CkWZw6934RIBZvLw+sxaQpDNyoiJfVz
38Z2ylmOW3avTzjGFcDPs7TiVTCS3vCXlCDUDbLwrbfFkyw+x+hljEsVqQVz1piO
eEvOOqCncxdnThklmnN+e4qoEhNmdijRbbDnVwsB/QAPZF3At4WUDx7RNn8A42ye
hkj90re8DCfbvHjiQWiIZUGZXv7a2RMMlQRFGlT2aIhR6MXBz9LSfY63rrXzAIMi
TMkL61Na2o8yO1rMQRIbXx2Hy/iFlfSXsJvL/57A6cFSYWwc20h8oFwR6nI39vxB
OxRye83mPeVtw3lbja5xZUWWs89/xTE5lRXRUxLeVRSsqrdkde24naZNXHAtaPWC
kn6jiFVmnQk6lK+8U5Kz2dnf098q0Gwq29ILnrDXUhCYQkEX9VZTekqAumlyGRLn
LVx1WM//Z6FDrKisACJi1li0sKai/7FvoOlXvuzClb3paDpjqUtzzxz5ZLHdTLdX
RQg/OiBSEnCR/7eTm/C3RpI9PeD1rPLXJcjrjhuo9MUBy0fqczULQWGWXzUFlKfs
PDpZjYRdo3bZyNyAMUY6mfO8SZoxThzt0Y8DkLqYBMeCfEVz7EyTYlQNyOxRiO/E
LhvoGAlwUIucuN9X626CWIsr0CsGSqhplOo3XDDcP2DtieyaSr5Y3y3aEkj58E4x
wS++AQrVtCIWpaBrcCJmfX+CucG823q8ytQB9tCL7HBZOjsFpZVAszCX2DoBuCHU
GvajjRCE/tqxiehG93xSzWFYIjT1xCxHBLAy9Vl231yObmvrGnZiq5uVHlbqXzGF
R3v4/upeUOXSehu2XUIPPWh75ihbV0+OmFoAt29z3S+WJIyTpbXfrzKd3GTN2HDV
l8wM9C/bspsDpklFATalpgRXs5/B10CaOn+UEXv1Q9I2ZieUYVTbKBMqUMol1uBx
iivvEpkXHBMJ71ymgLwRi/s+9sYQ2p+Vg93MsElOHjGNjNcEPp/m1rLtPZeZErFU
VVCy1TZp6H+3yvGRLHumS/6nRLp4c/8SPdyZhtK/CptXoUgcJX+4G8Z5HlZMW5Xk
BotRVvGC8NQoUk8AVcyHdii9HDc44zstwOsAO3ysmlYJlra8lzm2q1jbMnjS32y1
PE6RVLPFPY3I9GN0z/CXfH6PpYMQBlxuHvXp1hJ6gYDHWWE3BJDLNPwtjZQFOjWx
sQqbJ9y1yqrQLOqq90pPIc6YxkdzbcF+WtBKFUofZzfW19Heuio29yx4YORST454
xUb0jYW+NP/amNGGV0zEMI/0SRzs1QahpzSqdNV9CZMxFFI7fuNACuNokzRqhdl2
1ZPQ5Sa87h8RCx9MEWg052ruBMO0+13eRc7nTJok0kir1YwPnpaoOf8inKKmHv3S
o69bzQOYMsOP56h8PZgLFJIMGB+WsgcbLepA1CRvuv9UDm4Ims1RNhB43Th5nOQf
FqTmfg0rVa7THKyFJ4CP6ZYVW2YCEN8vn/DzmQ+4gpcMnHR+4aHR8el9+R2jFPJw
/uBIJCi0ZLqQeU9cSh89gocgO6NAKen3dEHP+LgYSA19KddGzKKTvbPH2AcEfyUQ
XY62QqK2fBCH6lKsPI+f31AaJektZnfTYldQpXKO1P7AscVMDBWLiQaHN49y7Oo6
LRYlVBTiDnDVovOnadeNxF0sZTVRyLnzvJWku6IH95ClUowBaSrhqsGrbLa/7HBr
B+TrlVMh9lnB/T2D3bj4nL6jipkm6NWnwZmZ6adxpB1h7CVA2PGnKjHvNSQOyjXr
mllUmy7ydeiRQbBEiDxl9utBxfsQ9lwGF58k5q+ScFS2KC41ABa5eUasMtb+JYSF
yKgpVEKvirEotLv2rJTcGjOsR4vzATw6Dath1bFf3tpVdAPyjkVJBAuekAUzJDDW
sPS0eo/2oGQx61ND0sqma+qejgiBi4HMP3ZTS+0bsnWwP7OPUcVv9nV9v839ae0N
SySV7k1lc47wjygc5LX7gif6kUnI93sa56Fk+HYU6MvwxzVfOcW4k52gPJHKkwUr
FKi+CvDsYyWHWTDJrdSuxlGveoIjDw5IsfYj0T6qc9DYFLWh0ls2cwoMMCoF9IGe
oXRuFuYqMHx8AolfJCNFg6gByBaL/h9+gw735vyOY2OdCR1ph9Wij24wkwSoU+SX
WbX3QmRzptnGGnTNM2m3erqbZSMiyrKH8CTGvu9+jjF0PW9hZpQm7yBQjRcMSCp7
ed5/nS56kwQpHE2Xgf2qYqoU+y1CTUvJYqAh4Dkysq97rMKfi39S9O8XDfGnQ4Jw
j9yarC3KoD2awOmOvmtvo46wXc3BGOinOmZPFdHZo/zN/gekFfK2qBcJJH72TVf7
GNBJ0pJfJSYgfrbCCPDguJeH7Jll3Wktt8v/+wpmwdDbeGYsuxchw9bHfTzxUed7
abXyOgQRL911kC30pMiIz9JcaFfJbh+LTsGX4ncnhchArRCH3jnF7e4UdRMvY2Vu
xVnS4n5ZuBgREqXVCfSyBAbXiVeXxT37qEvKgOtlbuD6pVB/Aar78YxyM2oIUJPC
+//a0aeWawvjm8HaA/ZUGWeQdqAK5V1NjkfnDzKTCvzy4AxN47yuMxinMHl23jaj
mQvQx5Y7sCiPou7OOIhM9y5y1wkZ1+g1dPU5gBC7sdXfgfit1sh3cqm+Z7KCJRVn
jbwWLjoegG/ENvPN9V77+I8RCz3DVBUBivNQhSHbKqFqJ7DNDic5hK2CzV45V+cb
21t1zfeIz8jG9BVJCYlySa9nGtXi/9nLdH4+gKvWZJKZYKR+dIdWekVVOHcAjUlX
Cn/vREQuqD1LELrtREyEHyrRRkluddVo8lV3FFJMT8OdMHhXow1CLXD9RUJseTDY
2msrqN9NNo4sXDQo/B/9V6FS5BXCQnzmTsxngLBNLcItHPFY2T9MCRK7vEm9WUxo
ACnhMy14XVwre88rJtOZMo6Cp2Ohab/9bXPWYD0BtX5SnNEAhGU+akRd2NLS3Pgg
f92QmaaXWz6lLQjXZi4D7oedyeuzytSk5Z31kpx25n4LtGZT9eFtPBgB68V5UBbU
z5q/X/3ZLL/MJDhaDzYRfdrVqO/aiG/4HdWnLAPZNgOt2zZrwbswnef0umt1VxGy
+s93o4nvwU+rUVlKvS7hW2RmhErrLHmoKcDEs8Z5PqRwfrYOiMzFs5VgWOBubQr3
XWjSyz+lt7X7w99KOhtzLlWEPZz3c4Kf+N6IDeJiSLOAGnAWYKhF7BHzgGo2+ca5
MDFhiT/s7EYt/Es/0nH9rDP7vHCnhwza2vcldOaUtEoewUUi6Q1m+zcsROGgQuXY
gkiKHBz+2tByq880AEpGM85kNrVb2TGeFEBgRNOhMv/rRuva5BRVU98m6G/hwadU
jMh6WzVdf1NQOC5RxyGCOv95RPH84YrGQdHfnCQDHE1vm/swzbJmc6hcQ298Hr/c
sS+4c3nJeLy1jKofyhPs+AhXn9YFqO4g87bgEFaqHVSOH7cYHQqpGwVb2b7ccWay
I4YgjtnVf6AE+XWtfUKzAKPO/CJZlTPDiXGC59CCgUnXhAaSjwwifNPGXN6GGQqP
HPHrqld6xJxwTYhdTbaTToVE4ySlYZg+s0m+fU3FjTRFg2tloO+Rgy5dGk0Zn5gt
oXJx0NUMGaHbw7i8K84XRnIvLA4L/ijRdA4RkMSdKqc5Jhd6EEy1kc5gQvuH6u9u
kMuakLlz/fpxzW6H5QTceg4T+9SGscM2qDH5qF/fhNOSzm3gNEGdvUnzrwrXAnh0
U5FFA4/yqjcS1QzpMaxX6ayPS578yJ6qCOdui60wNGeif4ei7EhPZwEpj4/eAVxF
cYfZvTgVQf2n7dLWIuvjF6qZSlO9uRwNyTU5o0gOi8iJ970CtM0o+H3FcI7ddf4H
vq5cLxh5noFVoQ0M6QJ06ZacEW2vbNOPnt6lj8C10kjqaPoSIHhjBDtfzaf04aNc
Iy2Tj8A6Quy5pQmmac/IYckujSsSpRlXUuGe4SyQedvfrmEgnf9sMbOjQ4+r7etE
J2vUlW5CzUxSunPfzQeZ/RZDFHlFiymv+q4bT5ttbBuulbrN3qYcJLoOzwVkuoF4
qePAEFggn6ow0onP4waMaLp/rBRrPoHW1FZtdyJJqrcKKR8McNut+9oGbFiFiAMK
xo6dJBJ0TLWNV8wof8jnxmm1XDBdjDayl2ZRBk4KkCCR/xwMUGOWiMxw9QGvatoM
vmr/nvIHySC9vEDcCQ+15Tvx3/X5AUVG3KlmImoEWUnctL5kZWSupsw+vC+iGdZZ
uq72xNatHaClygJgtPjVeOpAbbpFgCuHfUyp7/tqLbUuVhGVJCeHJBGsJ2gV30+X
FuI/R2HI0/ha3kuiK+fUA9Sk45AKVLGUPrSJjFWh20SLtupWf7YtAgjY6chHvLpG
euJYIvmMRNMTXVf1XjCTJVjw1f2V0+nuwy9SKPslURrzWvCyHjPopaEZQQoxt36I
wp9uRFkO+f59zpzi7ccTmRQ7e6qzgL0rvBrVkzkX7wOh5pW7Llwox9vK/dLRMj6h
0d/aK6frBu9t6pP+ppgw6EX8HCVkjVl+maV36SUAaMeJxMj5qcGTBfLU+JM7MEbK
Eqy87/PbouvMRmLncy+BwxvGLOQUX7aZSnYQMwFENAoNcNlyS9f+M/4Xznn+JVyP
2ZkIcGSCC5U9Jb8E5Zx+HSnkVSQrfsf5uPiPGXjhXHOdmrS1uLwFETYBSzHV1yvZ
mIrdxKWYKewxA8C9OxRbV7N7RdV4R4aHbNHGWgYUcEyJryeXRxY7jgMYGTn4B1e3
N9ZqgUTSm4jOHjl/LRiuVef4PO5jgSph6FIufIUyotxXeJiUfd7uCF5dBMR7SkxF
KnyQdeRSjsqWNMFvvwjtUJIn1yQbFTVyrbDNrOKgXsQLIlbHwiAteqNZl0j3GC1i
8ywXw+zfpBuomRyBaVzbvEO4dat3kk3X65F4fN+6KsaKHsDopAD/BzD/lqR6KZ85
Qo9AvDcCJvO+5zw0H8t/jPpb4Op4luB0ARfYSHam25YrNEDuy1ARxKNEG9RsynCD
THjPE7jvr+2/KMcEvwcHVxEOV0bdYX181Z6PFDWd4vPgQozNQKKMSFLgVETS12Pi
SVRr3v5IYssnOBUizMoN2Q9Op3iZfE+vfLKU9EY+xvE0pNfknIr/WUXJQlfvVqOP
Fa5YHA/TpKYZRhyAs8CyRSLKzDYbEjcjWxBsllOT6XL77dyvC9bac6GAN0olbgdO
2KrUa6DtY4+tqT8VXsk/dEIdkoTyucTPAHXsL7gjGE9QRMPAiGvAYXwFbFVDwSMR
LfG77l5ijre/f8bbSJejpov3aYEjB839j4PE/lgnnwcY9cJPY7sjh1p09W1BpNzZ
NFX03t6Up0SvzC/tHmDBszJp2j9AZsjI7FrvoiSQxSzvY29JJz3X81RoYNj+GYtX
UwlIcq5V8xHLKM5bG2p+w92baOZ5WpD7P79U4OK/kfAGuGCrABZU4khw+npyjMt1
F4a1f3Nj05glF+4x/DSElv6c3jmkFCbHAeVoVjBAAKGbTHSl+/dBrQdE0VMgPOgq
Ulmhr1brXsLBMD8XI1e1Cs5d7RDdKSMsOlC+uOZOmixqK3ljjUUnyHN9m66zA4DT
uQE9Qtc/8I1JK9CLnbVyBAej1gTqgpxmRho+APJqSib+NYe2ewLEdru4wbiW5J2S
4wnqclOw9rN8422UDNs+RTCJXcegQC1dHjB3PJ0xgVrBvnz3pBKTfSK3fa6/Gprh
eEWQ3gZQDt/46L5mGTsOHKEUG4x+9nSvs1kSIGWgyzxKMQQHtkF6nEjdtuG3vay0
D++KIZZ13IYr25D6sHaVU38DcLzm1/S30XOblZh07pT3YzIZsWRAgbv/NkpPdOWl
r8FXcesbvo6YK6S/mCV0nseFcDOuonljlKWGS5VIa2q54PAIk9DK4iWOUM5XbzZO
QntGPaaZ6K66755I8aZ3GmIk29vU2Gc+w9zX9z8yYYvadl5vtwWwVj6xTt3BTOAE
zhRcmGUA+hAQ+2UBFpA5YVLKFZHYcWJlECEvgE0MGzB/HUw4r8untpf/+jabzh2I
o9oYKu0ORBSHRRRQRo+G8np3eVtCAIoMADYe/GLB57hWzgsNAabUbxyYxaSb2ASg
4Z3aDJBWpkjstzVqdz90bUyONuCq1QwNVMLpl9OYM6z2ZGcAit1mM4H1i/7EEeca
/rZ+cIGjT8ZXhqFD9awWYp3vfkSR8B+8jI9pLCKMWuiC4UkRpMLZ3msf7hj0HVay
PlWcbKhfDBKIoqyBn6jgnOuB+CbyqLzVKnG++tOAfAtt1RyMd7tBT/hqESwAbR9p
WZ+cGhiJcpgm/YfyrBA2auV/Sn9vt9VqEItOPRYGqOpIIn/Q8vXlR8Zfv1kJ/xLA
PiN9TrJDRzs0/1jp80racbB7id78+jH+EDol9BynXeye+X73+vTAt1Z/V/5abV+n
0zUU1QwCGwZuMJsW2mMehUuM62sg6XjAbuw6dH+buWn3wqcKBtRCN5MJgE8++vN6
7zDf+EcToCnr97c7iFFMlmBeeq/DARfCCfybC2/RN8cjebnuRmQk5H3TihFv/uHd
vALYI0td50A1CIT4LleWjeP9ifLEbXXeq0m6Trit3XuJx55PuKabypwMtCewoTQj
U5e67Run6IEGrRRSTDVk7QjkG6KQEb+YJFotaWc3mgdW2oH2TWR9H1k4K6vXUsXM
EfNGF8DXpX/KRn07V4msxaFdCc83lDNGhAtJE1ZT9KX9N90ApPirRghp1QxtNykU
PSrTVGnbWp/pF7sBfDTUGP4ctElPuRaUV8KWGgt+xW4yqAhP19Yy62i9MX9593pJ
8MoRLP4FkE+VM63/m+6zjsA909MoyVK05UpqrdPdgu16UNGXdkXfj70JQIk7i8y+
CGwwXRWxqD0iULEwEOVoFPAcpDvj+ULtMAshjaD0oHe5MgPKnEf7AmIjLmB1pxkX
rkp2urLZuU5mda/i3LPYbgslkLQ6JhBo0caVE1VFzMAnAGSr/OzbXlX8FuHwgUly
ncmmWZOzgUA1YDIn/xHigsTJLRRb7avDA0w8d2BBcaCey7Kqo6atZ7RV1rJV7hF/
q5waoNC56a2RS4b9K9pejiKYNQ8mCgQ90hYt6It35QWLh55BJkTArS80xycDR6+i
xCERc1vgXIBVSnS8BtEaqY94REU/70cqhy24IFoMsRfaE1rB6y3vB4xegXfpVrW9
Sauw/MNQLKPPDHGlQYzt08j8NNeiUYQOndftGMSATHLHao/nUr9/nMO0ZGxUjAlk
W39Ac+XbpFOtF6B/wq4J8B8cUaS2daAbmR0S8CJBso6/gq4TlK4RyN/FKCdh6VCi
j+74lMSHV7M8UE/Zcelie/1yG1sXz5mGstgsqbNK4Jh/xgyZ1HFfxxEhaWfRinHX
QbmjYLKLuQ566waWT+EGKNqnJsJwfUyHYYVIZjDM/SXKulF/cgAZW24L4ROTNLE8
LFKqYviU6KKsIhldZxQFJNDFQr2tQ/uBLndCgfopOEz+7BfBJEy8uKXEHl1T3+ji
lrUpwYI3AmWzXovzUSoZwdrMQgIlBz8bkO3lxUEXBbFWpRCO46kSE9/bkDv6Xuma
Xv8DJKDVmXsQQ1x3ehYIoZiJxjnJuAA3KOy75ZumXzQGzErRrtECDkLASkCIgOGc
kn+2gz2/w9qoLeelhujFfzuWM2knmFKTXAHDHiQr3Enb9OoDLSLoYFZ1iaX6km9H
+rswfF6CFHDAHdcLRnj/1Xd0Y6TXYNKQEN8kh4Uh9JE7cCDSrrZ+LHcE6vEKumz6
ieOEN4ZuGD4NzwpAU7J6T4XxlrvuQMrihz66ZFrMkITDzYZHTICbCRpgdVDU/AhF
rYuvc2t4xOjJzwQtuWtdZU0KxRn3sX3NvzfB0ILa3QBOdiCv9XeI4cHy8NjGrACI
G+HTKkpong3WXwIQ2JG4pqXNW0jkGenGavjafigBZkklopHMI/lS7OF58Bk/UjYb
EC28OlhtqcBHx9lc7E+IczfAHTGBRHH+mgfS/aNScom9Oyk+g20cED0CbR9Qtv9O
Q60GKu/3V0U/OBK4Mcs9A+Lg4+0ff0ylwBlCbIBktlL428x3oj5vZM2GJtyncxD1
gtcWs1Me/OKipj8eoWyFXJzMTVwhWEx7dx1vmfjXfC8Tm0Rwmc1wubm1w0mDQCdc
AvcCjcaw74G9AUXFGNAG7EtYcQ3E4a6W5sW2OKA+yMBFZ2xGpkEXUZDkuYu3R/Z1
jMKicaSfwJT5lwuvy1/FqD8ibdt9WVOVIStyvyfTul7fkaAkNSTpFpPFuwKZrO3u
1XrjvMCFJxBoWgmQ7smrn6NGfomP79HyRWpzymh5JH4spMy2Bcp3gGihgZnwxs01
G63CT6QxbrXrzvvV86N9W8aAuC5Rg30CvAn/sgqxc0w1nXW5l5mLSWhYa697slI3
Io3fk0cawXwaNMcMHKjLAcaPMA0C7+hJ1/FfS5TywXXerDTob5o2W4cA0xz3OuYB
lOSg23l2S2/l4eEtLPS0Gr5dyZqhSUia6MCMMHx8Or3/0HpPOxnh4TWhTigiMa5Q
QEWWMc35FGOR7Sp3TUBURV02rUhZl6JR9ROYjClOJNsk+Tu+RaCp6jFACXEAGC9Y
I4Q/tWB4Gv0WwArqVgh3hD0hxpK7OGeSGYpFNwzbkpawY9wcvarHMiHdQW1htXva
OZUG3mJIP2qHGdCXm8Halhi8NYrB6Ns7VkfMu89muZHXotkUirwm0bs3t4zBW8/d
R7fkUhQBQKtLD8dL8vxX2lCTm7gCP2M+lu8lFMkyesxMpMSRMV656xlqB1ZB7njy
xjfbFwVQHM41oOFwuc89MaQIYd/iPULQBQ8nlRp6tyXj1QAd8rXH2iwTBV6lZo6P
aJrLT+TwpPjB/m6tq2Z4q/7VvkRBreOvqKmJfOelcGMCrjvaUkFMS6Rh09dMwtPQ
W6k5s+/ywT3dMeXCk/8ZDsZDtcoGbSKHJBh1i6ki5D2FMgBSmmYYVsfPHukQFWYk
b69PN6dBnMyGf9eYQG+kFoLazU6END7Ud+Ih8dovKZpMjfnwjELCynePcKuPpfwj
yqkxRFxZcE5Qlja7xhRRbTqawADCmfN8ocRt5blkb3ScogN6I33M40kFCQQspl+H
wQ496jRe48hCQC8DTGHA0bhcuGyZ7uIXAYhBQhBdtmFYNtKtpRKrXCs4rVuIfCiO
TKzwOZkOiUgBd68AYROTV84gd5G1y6Pnm2nmip6EFCsBmijjrTnbhaz8AFtCPKSw
OaRGsq6dcuJ1eeT3Tfa5YMLwVnBIuBdL7/0ImZTmFhUwRHTCRTGsmt5j8UBMbYQZ
etI6dta/7Q/ul3S8ghD7mkP16BdxqDLGbXuU6hQjdsdt96sLb7W+NNxGZkjAJ4ct
vHmRO2yjxk89NyKmp6+jwDtl1Ui6T+8DklDa+qxqu0+5xpxf6wZQWkWvCFH3sVuL
IY0mvP/8UpZ6uKf7qatMN2bDcbvoNSDbx98Q8HX32F2xI9Nq7yK+tXM8QaT3TNu6
e565Z3WUKBmOq9X3+tUzjsiqU5G4ZzmA5Jrgi3eKcpCQwWU9gh3lvY9WhwVjfC3j
xRhu+ocn6/GsATI1MJQJOw0N7BiVsRoTjGRrYWNMXqlBkrfTEBOUgamtyoWrSLUo
gIRmUnQsid9COcCDYfypwiXfltXdkIgorZWrMEKZpE0xCukTWrgd4nQF+b0rPC0N
a+JQ8DLnO7BRxjcvfjTo1ml5GJMzTc+x/5nhJlHDgQUjebahlsw/l2Y663S0dA/U
LLv+eifBJgtk6kqrXNCl7Vlqhrpln3TxXDEcAZ8xAus18PyMSE9tSa8tKiet9pxA
mH3pc+wchBqss0NCtZQnGmHYchqY2/0f8NDHorKdgGb1qpZJx+EuD23Hq9dO6A4h
FdQrUFw6jWO5MVxUobTSlvts8+bsSuV0ltqYzSi8vgnXteyMyAgztoBgZIp1XZtx
9FBlxEspyIV5Z+dt7eo00Tn6pmoiIftzm5L3zbSvGtiAO8zYZaNSX1PgzbuKi98W
wIi8wrvsQZuRxFxfSW8skigtDX1SGGc7IIs5fN9k2T1xhKUR50YQHC+cxRKkkcjD
QNT6NhgCnZk74tAHv/oK4WNrpr9+X+tWjSR7w28Za/XZImVXAHMxVLLP2CPssdLD
EEhqu2zX2ltxnXcpu7PQtJH8QgC6PDdEagFMbdgkb3Ib1ZqbQQE6Bz44ocakLq7t
7ClKDhFFKdyM2FGIeyMcWupuP/VJ+Iwx/JvElI4O0Yz+1DUZqY09ackuOf4+SwSC
rpALVfn2rhYFNqF4sXG/DxXncHBnd8Omco1BjNWYHiMYzFEIFCSw5pRqm+hJQ1Cy
M2n0IvwDqr9UmUimD71gscPKJK8WyMFrnCpxAC4s7rvGiryVNM6s/5JyLASuIYd3
72F3L+sl6lLn98qXbgvMgucXMi4OAYBjnL7Hw7YAF80kwJ4lAm67aRR8PluFNAaD
qeev2LcP0/960obeTM4u6ibRjaAiRtt6B0PzmWwKxymFB+oKG5oOqIvOqvJ2XV83
5qcgKiPRS+IZKef5QEssTpeZvaIhmeWzH/4JjyibOsD1/TpLzUWsDjTDe7k/VeMi
zwUJyMvFPaTJ85GAtSFzOyN0YlyiqVdc516gFeoM3D54r0X2ZT9dZnRBqsWeCyer
CCqfJyhKgQDIoHvwHFwOTY8f+tHwF113Ea5M6L1n6xogDWayHcOPFH8k8T1+ojuY
pSyWTxQrSsfAdoXtPupKR2C4/tSFaW07XNSF6+XdshpPHf4ruYtJ5ViEfTvAHh0b
XLrE/MYL4SwiHUFMTwm7WzIb8vPASXXeR6vxpMZ7powJ5a6Ld6ZLLTc2MeIAEhB9
DN4OlkqxIUcSHYtYs9ukcP8iKxIH3M4lG3MTZczhVGLhzC1d1fkDPBFpD8w1I5Y2
PSJ7x6fMLsU4PRqC5mJqYns8tog4wtwddtuoNCnWtVCIVJM0nuTAyLcBqrEwmT4k
6DoZBGIKG9JqDbnsBu8RQ25MmCJ2eVrJkwKRbK12hbWgmyWaXpFobowtCLSKRvGQ
zN8GhEy50rrelicn6bw0FhXUQVuwwUiLjfAeoEmRiJ8xw7o2FdklwDjeLYh2xcnI
LYCBbGsSGDUejupTDFx7KQeqONDu34pfrZeGKBC9+mD6lLJ7F1c5g8yKmSu6iFHf
byIOO/Sr++Agn7CTaR5R5KBo+Oo6xjbyNiXX+iwFCRfdT+2Lcta8OO7sxyfV2XTz
U/0psUNBsUvD9xAUah1e93aAGl384wvhXwLVlHplNtgbz7T+7AJbm1olZ8BuqP1m
gCaMmjtX5AiAAIUqYrawwfK2T9963UrmqaHmAFqHiNouvb8ivyPk37xnKmMhDZKT
FShI0w6332djCAoHtVCRDbAiWWYjJKKsxUWKmN22Q/r6XULfEqaxZoRKgHqB43MM
pPeIZ+DSdMWSB0BNOdPv8GRuyX8F6qz3ToLKmlNpb6+XV30bybfvO52aujwFrMbN
3XIVQlwJr5XUMrH9m66mNWzLu1trUeD4SFTWaFZl0Xz092aZJkh1qgL9XYuLkD9o
Ad77DHTtROMz0sDkA38P7A6utU5tMr/mqdlvRZ7ulYGzu5sxlyWYixX9GI0cGJAA
oKem/qIuOGXf6xuRBMoATKwCiZgDrHZKjB5Fq/GaCMg7yAAv6kNI7oih1KGjtSQw
2MYYb00yoDJCdrpcWv5Jk6bBTwNC76Rn6bMVnVVLz+mEL7ZXq0wHNzW0eeeCagBO
pjHvDNXV/MPkMAzzQkzqc0hTaHAUmcJeM0LM/xpegZ2ambp+SZ/IrgXUiojw2Som
awF0j1ZpKAHgvchueyzbbreQ9o4LUkgKC66J6iZARcmXQBSZDPmFnuAnQHQt6Tp9
ivKyODcvLF72cBdahHbxWEVLm67kF7CePlYpYUctoHRT56Kqkzn/RVs+d6DufvaM
7TT4LG9G6TUFCxX1qYVRjPZoxXwrHeRiL0H9HuQr2lCzzctOc9Eky0OwI4btIYgY
qCD2rk9JBcuudhw0pAZLOltmenAUvS/FanIUs9fxVCYxI+rE5Wbvwq56wPtcmk0n
shsNzTZZTXxl7gGdk8BCRAecAJ7Jk3nB29lnDi51en/2W797YI5z86v5fI7IDrgC
HTeUVNoQe8MqWPCR4czIOkLH4PE2BRgOoEH0p3RVO3p+qr3y0vq8yNTer3+/nGVf
iHketmyGQ0k/t7yFstyVNdZes2cyZGuY0TYkFBbJGNLWEMAMEyh4N2wtL02QoBtK
STJ4YkwXQN6hCTLuAnx6FvIRJiH9//eEwMZWx9IuLHcbCm5ejxS8iCHrJHyWRBdP
fL4JXde4wRism++zGaTdDJmY54br6FFYqXvXZ51Q4rhkx3Bmar00T2PLsq2F9WkJ
1dz9ayfMy9CioiCkyBPnyLNq4WMHpaOoBf9XbVrIIfHPNsqASDF61XTklBQMr1AS
fhmfQJ1seJcREEnYPq/kLH4FqlNowU1mVqj0quIct1tfKcxXWBsfrYn/QHySxJXa
xxxNWK/h/kcB9tWtjsD+dfe9OsALu/H0u3GDDuT52FSJSpj3Yh+7ZRtrU0lHjGfA
e9wwru7hamGSRqGaylMR4+9tdULZMigei7JAlOEcEyKzLWoLplpxqWQbT0N41Nw7
xthnV3g0zQ7LUqqsGnoPg4KYOcTsxai5WJ3BwpPNZl2cRmvQ97qVQyIjN4Oy4kl9
bDJuu7308v9r219V7LoI8StAaqUrUpcFPFtN/DYdEBSfxfO5iEJIEhI1l9nwTBU1
MFn5L0w4Y0cFss7pLEIxZHOAVVupyt5Bd2kH0Az2c9TT19qCXpWCme3sB6rtJZ/l
keQil8JGyb7euHh5gI/RNrxDJHr6baZ2wKnG1ySl0CwgueuADlMUjP0ws/1diQnb
mtB4vWom62IrZsf39yxQBy07iF9X99WlYxaMb4lRbx7ixUE9OSwqEHwolu7xrX7w
wR+VQx/xBfkvoSPfQXHTBKfJoMbX65cu8NsawdIiWo6BxS2QNHxlBol9hzvZEAAz
7oH/LDH5h/cwy4Xnu89QvgLY3rvwvpUyUG8Nfcia82F0xwYaDriZAiJxR5GTWD+/
QtJtljvsWEGN1ThXdXChE9EHsE527gDRLqkFCm8shdF9RoTHpgaE/Ay1y/TJPUha
EaorsriNWji1AWOv8Q3cg72vyDE8mnfpyvI+iEZSj88Roadj5vOxPZrAIGnTqW1Y
7o6ZSsOvP6sO/c++J3+nOmsNn3chkduRtunrzjm/06Ll/ljkdS6ELTmh8m9l7VAQ
uBHB12VUo8cZ0UsXC8SyXPt/9S1wMA/tX1WB7qGDEaE+85aPhy+d6NfKaqs2+NNB
dEAlk4sNew6B7ZOSYD/GVObMzOOOR/4zyR5CiTxD1JySH7WhjvBcb2xB1HW2OBla
D5FiBG9i0XTE8dGVoK8SkPmdsd7fL3/PcahGw+Wvjc4TDcTxUHeL/C3/5vniWCtz
b+L/2OxeTUYGWnaoOxTSHzz8EZg4WSPVIs0BA8DDGSSsYboM2S+dYHTSzqOLWcge
lzLrsvoS37mNq1HGnQJxnw12gAC1h8xibdrkIwkz+PRfzm6IfNpBVRSEw2gy4lun
JFHbtVUEXALJK+WT9KVciDQldL7JqUJ/aOheSbcW4IrOGu4sUig2QXfIUzd3zVPp
msyTvpbzOGmu2kGowreNvKKcRua2iq0qFydv/7OWbkgwAF1C7aNRlrGypYS99h3Z
g6MMQ7tXLHGr0uURV39bc/t3VcNHg8dRhCuTbQ1rVipR6H70f6ZCbPU8uYyoprJ/
ECsBS9GpVUsUPlPi+rctZ9JATCsNGEHx/Bcsx5GBIybe1t4yPkX8IS3TgcxBxK0S
doIXAN9weiuwIf1lHi9JxxpcyflWKmt4X7u0oclxoJiGXsFGwvhyvOsQDDlDDIDb
N35ir4Y4svkDtv6GNmR2UIrCC0rrZ2NyfUi9JicBtr5e/xdO1Mai3NQ+vD4Q5uD0
ONylvwRE3Rggwtf4Vmnz0yM29daf1r3l85O4/ujDImAXLF2arzISOer4iRjBO+pS
Z9OmEv2KdvIN5qtJN2G4L4uMRbXM9mx4dKXL2me5SNjv1mTRw+AdWx0KLiB/FFl4
NKgfL8jpeCvtrASkzrZxRxZ4JOUbKXyqIYve5s5pEZ7MieEPFbkUksDTzjNzombK
sxDe+0Myw39jSxXa/xeWI9BN4ESQ6MtDqA7qdPqH6pWsXCsG8TADff/edGhnTIh+
K+2W3yjdiZFOD8TzShRhMq7In3lXVjaWbWrtY5nfxKNbMSZqxZMbJIK7mnApP4qe
I6XcNytUbQ8Z5Sxw06v5SK5idj9mRDHaHCgBMI+2JznFwLuXO9TP1b3RgEEhOXLC
pA7H0zwkVMLALepK5SR1TR9rEjawcWvSQNy45SDpH89cZbkJ/i9L9Yf/ubOpoho9
2x/zmmEBYJMPG6eaURl8NsxEz3bT1R3VDkE6KeCp0baQVopVpvjtKOFFPR2hCyQz
6H8LfRXsOjFyvd3bmvWTEwwKwjCmuHl/UI3lOXKlhS5e7LNaw3Q1h6Ff3pgWBNl1
XraWUl7NWw1OAzTvsI7rGuwkMhsziVbbyGnU7osZtNIFDldpHMNF8Yrk1lpre6ht
YzAEYlZ4TKyHaX7rewo7J48ZT+urVllkuOms9mQewI118nByrg4bZVIethNjxaxD
Ta1/n6aeiMILhEpJExiFwtmT+EXXyxah8ZqQzDrUoypAbbfpttamGR//91moOzUM
St60SzZ3XjcUdxTDpI0wwwsP8VWETE3abUH8Q7bNV9BD4gX0OaLL0DXFA0b1ZxkT
voW5AafvWzZoIN1/T2GEYAAaQfbLPHmHbpRhkU9xmllgb3uWm2H4ECo4FXHi+CB4
gexfxq1YbE7tsBGEpAX6aapISMpgdGFHNtP9SvzpMzm3EajZcmHyrLp3hsEnuZHB
waKMdrgLEdWF0jkE0eysgi6CCPC/LIOZGAqGxYCikZF3as34m9Z/PLC0/jATmjeP
beSRg6MOjra65yZb3cMgDz/VOHK2TVwJSNaoUApvz3tDyDB1YWJk0y2dC4zEPSUa
+jXpA6HezDqGS761qu0Qcn6MEZ2Uv+tRYx/WG7w3yL48vnQ6nCYeHc6TzGa4bqza
ROZ0SywDM8VUm8lufj/vsLcHkwA0GqE5Bl9RH0wSpO3V5l2kByyAgldzU/qGlNPp
nNbzHhZCJB5giY/aACPPpp9Vhjbnkt4MBAMVwYZkK9Z2EfKq9KwYvsNH1LPTwdKi
OhMuumLiUMZECfiouhbAVlxG9CsN56nbPavzCdW0GaCqWSRn9P6kY+7R7fB+wIPz
Yqve3jVCntJvLp/rUjI9xDoYgPuoZhJp/DKbCSDi3Tl/aUjHOTtKjbDa83UG/Yny
DoInUVwgfIF4tVgp48dKO8WGvDI6aBDYtTPAzNqjXlzFO3YApSrBC4q8WILdSQEf
SxJ2hw63Yojscm2hYk5+ZYV0Tz6UT1i8I9jPOb6i+ZZyATBM64mBRdXIdkL/ZE/Y
8FzeooprJDk2roR0MHBDTXPMlY6ajP5A7/p4wBcHuHr/lAz+XiLsxS/VqFz5r7yj
nP995lzmpyGT3zQD1pIojwTxL3rcgJzhDiq8zFlIPqTIev4wHfO/1mbh6GUlvxYT
AA2Sh1g3m/iacT9AYAatsLhcMkgNAFBKYdiUraHuELXxiIyW+vvNCA6+X1+Kuniy
fc0UoV8Luu/YveiY/cZ8R6DizOh5DXu/pFd8GwLqbJrZeAbVUAmWIyjpTJjMLVbC
NETLL7i84pDBDpyupl+/ChRbrfpEV4BTF2AtCPj37RcXS+86t1aUPEvZZeW9nB3p
Pk5hcZoo1Qt4eBG+nGovYdYJlrqUtiaHzsJKumoMnzxT57t40368lGPWLF6WwRL6
pKnx1jGfnV2eUYJnH3sBXzG23Cma72Ff1PMBytpUi4NrFwGJnNx/ffo15ZljGlEe
UA+OqykZGwZvoO+96oOj+zTOKFx7KWngSOfVz53RkjcnMGl/ouUimbakLzfpDCoX
XUMPTzmajds7ZQD6oUv8dtfYPeCMK6nvION7nhaK+S4m2QUmlA45xZgNpCl2/nbg
qjtO5eIo2hLxT8hYInLwDlqX0eVZowYL1j/HrPCljza2+nMSjgB1f1fj0tIHf1eK
hd5c+L5EEYJJF7/L+qvxg1xyF4l2dysiVp30K8F0wDtYgpQYBcInhRJaZq0u18FH
wbnZh8I8LXI2Y+LiRDSniHZAU3T5XBHVl5WXR9RHThVXBdW0me5o84h2j3NehXTz
hZ1GIzpZzIvJqXJtfBCE6ERzm1zjN8HsNP2vklPFeUrq3H8rpbkmGS5eTm8Catuf
tMXbuAoAFUQHc4GtpJnwzMWW9+b5MemcD5VIkKlZXRY0sBtT6QWEIz/fpra9PMvR
iRXMOXMgSEM3aOyH7J4Bat4BHkqwOZ17WOnocI8z9h+N8KUNhn2E/6XrUSjfhK6M
03sIlqs2ybACxguPGOxJn7nSs/kRywjkaDkKcOf8UmRceDdfpCUbF2xEWUpyBAzv
JcwRj228CAeA/EthOoRFkrtU7RZnOhxiFODrDn7GXpvDh3R24r4mEC58eW+dg0w0
hbGnNqsjzBIBB1F+0WJ9SAAmtsyC4bcxHHLtAs3+BQNI6asb3VVxsTsvHEh20ucK
OVPKEog6Drn5EWKAGddr2ke96xvsQa7hPOlWiLMe7VhOG9sCZT5RQMuJHaryyWXn
0x2P7XtoiZ+VwaS/B81SNCT1ifccFtGLDbxtvQswUzyoyaetgabuh9PrTxMpGiqL
UaTxvXuLEkN4EOUlRV/zCCvweIep5nOVyrIuyWCw6mp8p6kRyBS0PFCEI2tEk4HI
amC6YC2o56QjYbrk6lPo78fN/EAbS4gXgx5rCJOxne+bPFfVshL0oLci+E3BgztC
QurQT/SoA/minU6I03waBb9r9l/Igh1vgsv4ZMd52627h1zMu7XbYCGdmVPgSCbu
9nfFmJEV/t1XSNTK54Nswd76Ra/wf7yxUn8m3FJUYfMcWbgF2mHk3gTupgeZM7n/
WeYKn6MMe6v+RZR97m99QUrlzuUBja1XMKij6NjPcSNCFo277oGgKROPRNbGrBGH
Zd/pykliq+LacHPI5mOmTDK5arZDVBtaEOeEB/iNQE52U/RREgMRxJfqk6OSECba
nEdi8iZ4nPEA7hNWcIDWkyp8E4jeto/Nh6UBOmAggjb2zECRLgsvesAmxTfu34ZB
rej/GyJ/O0sYRup+HnZ5O1QF9t/bdL8kJypKkzKcbWufh1kKM2rBKUdPOimYl4hn
2V11L+5UgH3F0ss3/aRSjL4VlG16xF/liMZikJFLs9KhxhWuaV6dQxukK39bSYaa
+7qKJQ9mop8gxNdaAZMaTMEgs++tXMHOrHbcD6bOXWgA0PcVXq9dt6Ovd9DZLsK8
VKKFEUdnI5zSayBpRmP8ZPAwRdb3Jk3rm4I4Ett6gFtNHHsryrkYlw2Gh+y6Y5dR
gqpkZXDeTB+yCptsDxTow175ZlL1prhmwToqeaWFAxWEICrdDG/ePFEqvJ+Pbdnr
Ur3kZyUhdwXkcHCoGTQC+bUr5hCrpfEgbMeqq5qQQK8Iqvj0yzKzhYTkqxwi6yBi
Nph2V3i8WvB+jhkjJ4NRQxIWILy2Vms59WR84M+FzVgJlpOI0K8UwmfD1CSZhQ3G
wmrdhLYNbPsgoTMth7nUqdfJs2gVnasocdf/JmLfy4bkNoHTT6JH4PjLAgoBKcgh
p2NfwtcE23ozt0GG3v13ihSjgBBIDuDBjjHK8bBG5WfucqZwwqNR9Qm9X9asdnuj
i0AvGNkd3TSO4GsNZv9WDkW1moYNpKXPHyE94N63pTD7pAWrAUU1kwblvtmviKiH
o62A+vKzQspVK+V27WfQw9YKBMxUsdwUQr4gkBvY+lf4AnfWibDaGkI6RDck8mSI
ev7mX6LFaUDpF5OOEyUYkdSM31ZiTtANNPOGqFdmOTVyr9hDAP9Tye4wVHOl9LOk
ubbdVh8dKZqRuTQ17sjxG9pOrKUTz56XRhVzrmNAYeK168m6I9fXq0UOgxRhKwGH
TCIBczYBzqkX4xKFP47hh3WhmZBrIrw3PFbvDUy6lmxSnX2e8X8xtNkGH+0vby7G
VJAw4JF66ie9RQeZSwxCpY0RnTMVZUmqhUa+95+bcQQfC7Jcx3UeBizbTSjjNgrG
Ri7nxgJ48uWc6wn00jHbfFM0n84BwsAS/JmpA/DiYcEprSo9NOnVnyJrRbHHgYFl
/jP/mc45+DYEsl8oSZTTzFItqj95t9wq7pQrx+LYTXEYhIWK9yWhyfvn8+1vwoS7
1OQmN1M9hTBNMiR/RIs59D3+PeQo5O4lUy7eimifT899/ktO045KE/C7CUAxO9TJ
TnAWAcFDHa3ciDvjz7Qwe+26jXI7v4t6mUFas6+2LgUy8rfuUuG4if4tuQVbg47G
fGLWp3IoVz9ChE+M+FI0V12dA0Qb+Kluz0Z9ufX7caNa6KVH117T4GaPRKHi7VTn
j3vUHvz4EzS51EqBgCy8XRkEgAsETpTdNbK4kBNHSBNw4VIQQfJJUZK3LjNezCe4
37/cqNZYfg5BDCaC43hUgTbEk5i8xSjHQwvmSL9ul6Yp5PuzEEmEGE3Nb4TZpZNj
xrSjWvBaO7YykZn7GzQVgpOo6mODgH7UcdK9UgDzaJLoPNrLOpFvzusW0pM+vQ/i
Aapxgq1VRtJ/xfNwBKpVy4/z0IgBE5L/q7XA2nCB4M8munFPy+rzMZU3X6eWF90q
S4Z/nm0cgyW7TKp95PG+9JKtPdculGRpwe89DuisxWhQ/UGPUMex96Q2nQlIX03z
7qxnc62kc84EXdU/r+moBy9sIByg7kZuy5dtxt5Wp4Y+ioPADAl4lRbgCIylI+Hu
Y1I6t/PyNjsjj2KMAOcaRcL5XhUMTWcJzOzrD9xB3hokgBljeh01N/2F3HKNAAJS
K/pd6kTJge3K4nB0dJ8zhK7N4sAGyhZeAspTNHWrGUmzqp+uKHYHhoJbfwhGRTuF
gLryDeiXr1vO+e/2PWLhhPEllSmqbK9EnGpVD0/iGvzYbGuXEhuZT3kpBCzcqHlX
fPbP2UyyI2Jm/RlyMQ0FGsFElU2kHQgGadUkl7Az6JWbbGeNL+ureBa0r7jGSk1O
1SxNRyGiXQsOCYUKS3GYhMZ+ThIabx77GvXmZI6n+nSoJGtEkfWZ9OlGm468SW8I
uWmLObtVclD+WoN/gUwFilqv262M0kQFY8y1eS18t4WIb+YIOnoP6EqhK/68SSS9
DLE05j+hSBx/S5kkKWpTuicLq6BGJ2Viqfwe/yl+Y2sRwpWdoitxwopWQKJ6ZYIe
JpkFvaxo4qSVWWldZBQS7S6mjJ136vjyTp/+vqLPkzIPIweZvVCkxEsmlg8smtxO
vq1x26QpCCV+oyFlGLzqjNG9CLt4KVHn02ZbCqRPEOVd3YbfMNMZsOcVmwczMx4S
jReDvfwknCiQ4g+A69QFtrIiL6mWqwRQKtCCkliHRIq6mcoIYZNaLO819dhBYup7
NdHk2e4nB91kQ+qN3YaHxY/SBW+UiadfQifKoGJYetycOHmyQD735F5bF1/9szvi
H76DLfGWO5TytIPNoknnSR5uc+LCyxnVpo2ev495U4jid0WpWKqZ77PjS2YwbL8Y
ZTYq9SnybXLoJKto9GXl5b/OUioI44es1RqMcbmSaRuswlxzxILKGrW7ngJV1KtE
stpJclS3RuSYQGqXm41wucCgnNQctfWc6C6VRkfwmsRjWYr06ojj2QNG7yjPUOxM
gGmgh3EgqvNmS0veRggR7t5f1egMPVcj/STxgCvRCUCBIalFz2jLvD1R0ZTTC50A
kzLdp3N6uZMWKNsWTd5464wghoCoPwYsUgeHITnkQZYFFds+9zqKiqLOe7E0zgyM
RK7BPs6Z0pIlfz+g3qYa5sfeqVH83ayxTbvbM8bBBNE7dhGqFiYfx1Uamf+UzuJW
5JUspZtC2KCbo5GO2080slX2VwxA1lWf8XhxyZh6Y/DQgDHam8HsRrttVLRG8va3
vAMNGiY9h5iVRXjl016nyT9LVPfsAlZF/KBDBhXG8gr9MbjNjzl66+5A5O/rzfUk
YMq1Ck8WGKS1eUjOOj0atDekB2NJb0Bo+Gxdng9OCDkCiuynzqUA9q7t7qXJUStA
BmThChZAwGF5+ZANyt9xnlAOp9TfzFeQlKAdrFa71WAMTV0vofzc84yAlrF5dE9A
9ttLgIF2eTZi0ud4iObaz3XXx3uAIzntmYzcNBOtOKbUHHPK4vc2/CWlJFoCctOQ
w2ZNqP2+vDYbOhBUdGOvKGy2jCyp9Hp4MQ9nwHuvAiNjFOZRtzQWxNNg/2oVBFda
pCXMtvk6XGOT7R52zx9wpHURe7zZgLnpTzGMZsxjaK25xiFv6nRQ9I+T9TS7Wd2Y
dTwQs1eUNbpC/LQlfR8sid88I4xMRrhyZypA8daxjTqEOf//Fk5AtvdvFukkMsGG
3uFXxyUrkkUhvnJaJA3BPu86416UAULFRcDPDMjo46DlLZ089l76+6X4oT5CADwK
TSDo7PhG+6jzkPCR7B/73HwFG0fld+kQkO3/j3U892VsJP2DPOfxdlcUXKQHZtpJ
6i0ze2px/LHNLku5C9YRzVKl3pJ+x1BYpBcdVr0MFBZK7eQLSo26M+VOIc0TQuwN
4r/O5XaMaKovq0yH/c+0ohlhGq62WUHi8kkiMHVxp7A6ptlmwMPbrDL1ZG9Lp2fe
pTLLCKnquOdHbf8gQX3AKICwCGidG77LTF2zs5bsHl90k+tUZWb53KocoeGfeSiK
Qqe5PzD60sXeJ78faUzIb6uW3UjT/6+OEM9DvsEdip9whU1/FhJ1UZ4wveSomgGV
136YuEiJLoDNoljp3nKbAv059+Vr0CXquoe0Coylq8W+FyQC2KsRCZYQoFbJsO78
l5X/f1K7xqK9ABiUflD+tlsoDkk7tRl/+gHTbO2JDb4W6ifvAFxgVckOEktvINtZ
qFDaplB2KsalMZjXw67ixMBX86FfS6DcJS6xzxykQrI0FzjBsLVgEy4Fp4yQCxhq
B824NT4ntb3Vw+cLjVRMIOC7qTdyB4J9tULQWASH5Bjy5uhdHrW+RyapEn8N4sgp
DRxraXGaR5UPVs+h4s1G4g+aI0OR53cDWHWHui8ZgRpHpX7h9ql+lS8UDn1t8jRk
a7UL/Tt5jNdHixcn1ztx3Z9cJSOFxNhovdzQFnqcRcZZwwX2iM3B7R8dBN3Dx2kX
NnXlRdp2HRO5rWdOeynBsJaGNN+Goc/RtUZXzy84KN3XGMbOO/216oIdZmOwj6Gq
reI3QNwKjfSg2p3loCxUVkZhFguWv5z4PlGAaDs+lbZLrxhJUya6EWapyJidqmr+
2GeoXfWqLDF2qDD6WT0t0DF+4KOYQ0TruGfJl7bChchVlnT3QgZd/0vI9IeAroli
o2gS9+7H+povBs2Lyn7NyL98x5hK6kndC8TcZ+vXIOYs0BGbknNqcA9cQri1Ywcq
WiCXsSEXQR72+hc+rtZltmLlMv951aeyDQYciXC5lS4SYjCLBA1cXNzaLmmPPbTO
nb0lHUtAQrpgm/lQ6lLWUwnmfV89BsJf4DNefE8W/tsAOPABhaK2TxRdAdBXaqV4
aViwFUat+3GLDPkFjkPIiWg4R1e2fiCJwrIQIgz36L50Hg/tBJ/j1UviEt8UbvB3
WQQ6sVMirUekECzVd5faw7jMP3lid2oGeg7BiJPYba2UWw5h3PLACQ79EGEUTmhl
kwBzlCMjFtJD2+4WsLoE4XQuK35Q+pGdND8Gcv1zc2MTkXKlWoWPJAuJxaM3diyy
n7Q5hCrVF36ZlllrmxkPbPFqOpg2PkrJNYuJK2+rtm4h+WMhoPdmJ+rAbAvardzD
xmTvrCti/bFGrFGGAtlhXE3r+r/PpdXpmDv9GxpbXusbwRgesXNShDx720kO2kO7
Ti0yY5+UCvZW4dVuGVXSKa+dRHVHK8xX36ui46RcrpOw18wRb2Q6HhXjYT4MmTMx
07ZjwrDCOWvV/S6/2Ir6Qavbk4bQG/GMeGzitIOELX5/2x/J+QrW/iqUGc/nDGW7
hY4RDr8hCUInFecmHBgn9W0qHZoyYoaJauELGNOiOBkf8RtZVASsh3P7CEw4RqbK
qYaLHW+ae6ps1f99R/IIj+WtE9KnIeYQyDE+apnymXbNt1SkooNTNhiN91/aT+Td
UyG+BkaIUCTgjktqaB2cuy5M7ZmAqZwzhBauxr3GB3MffDFQhYs8QdbBWmb9VYyu
k10aEv0MVWkG7PDw0oREHAdcblgBs39eqI1DtPisuhgjpOqg3KfLbFeM3QVC/1sl
Ut3VSlFP63e0AeKObPUO0LrGq3AVTYAkBZ7pFqeQKCmGtror1P2jcP8Cflg796zi
U7VLfoIe4O7JVnPDMxN4HNyrSknnKttd7JBkhJsfA/lvxN8lI90G7twhfrJn8FHx
sp5C4XJ1cFemkYIDbxt+4NWkPLfOCFmmoXo10yaJNQZYWZjvJYR9WgHX193/Db1P
DAnupfQJ2VtPL7TvAN7Z03GGK+YMp306bWzc2YXCFHygsVuzMM57s0gFELEEyZEu
aHcWZH0eRPtdB20odhGQo+eJc0m3W8GDBeZ4NcQwrTX5BQVkZpl29oNdY9BWcY9P
aiBu7nWBSgSqDErmQ0IuWL9OZt5MYmq96NPGD+6oDMiRstbHWar1eMEKMNYuOeHe
MMO5OUOvNW/NZFDpWF9yJZp3sH5uzR622efwSMcbq2sajogi9XIxrwcdSimLlSu0
h6rFIphfEFwdGtGWgpT9X3E1MIrkMe8yfzp6Vi/xbn82MKVkP4ljsaCL86kn8NcG
nQaIhnlPYQWNrIWVgXY9TKTZ5bzrwHJrFzZxRBSUireHhS7OOa9q58kdgodjUwiJ
u6xeIMLEA9ChLgsUJD4Ec8siU5US3QclDWBxCuQkK2ySfmwNNyIecggPQtgj09yz
P0KUOxsMxPhdCLqgmwwIQgj3BatzKR3q9w1TLK8fDP98JV7rhWbslY4V593hNTdG
7x9PeH35h8a4sGil1HRSiIJ9m6/aTgVBsdoJamv59wslUdDKTTEW0XituXFPANrd
HpCkn3kBS6LkI6NkADmwSFxNmC3MaHtA4omo7FEASznV+aklPiSKEjfeJP+wYttE
M5B0VL3efQ2GcMbF+Fj6Z/TFHvLKTLWWb+eqaffzJUihxvo249SoBj979SymqfTB
3JxGoO0+PgqG0xwdz5JL5KCCHXR6AKrpslr8WpILu2f38leQdq8jGcyE6bQwibUh
OJarccpDCXm72Q/OWU0jz0yDWkbG8b/UTzcP7DjZU/Hs6N7LoXihF2fUqaq8CulH
haCx8l7/0fMkzo2qo2xQzlCpHkZ8oLU7Fqo+4PP7W/rXntQoteZkDTqdl4GTk8/i
3kHHi7SiBstw/1tpC+ouaOoYiyal45tdMtkioAtlGr9gF2yzIqyy5kL4t+GQ+pRQ
N3tF4AfQgoc1ambDT9/ripxsZViRyiHM5dt/0PaY6fwB5SbDc6dcwDRB3D/c3Osm
mIy8xtafblqJesgqPIR+z8jrDq7j3zsbbVvn6CnkgyWzlcmWhF9id1EbPp0q04PX
JLRq9JKQa2rtVwVXgC9g6y5jey+JcuHIgHHcD2lkHpyueO34qMG2wN53z2ncPLD9
hazWL5Y96zYWlG76O6YQ4glHbF9dDfs5LaMzvErpWsJ6KA/fEFF0BIZLj0gUTCDD
LDwOuUwgVhK5XwMrcceT/rvjIs5f29IB6ZZreW/8F1d32ApDcalHWcfDF72ZX7JE
JWdbG1Ph5ax+9UKn8Phom+tnoJ3SL9BrgGWc5vQxWCWaBmCBvDNDbTodgbs5uRy7
OQ3xwiq/teZFzRpC2mvPKva6oEqEfy+q6BmI9F/3b0HJz7o69H+cx0uXNdR1+MzU
fJbn0cRyMITtCwWt+iIMFcul0FHYeRbEzPppU1nvg7tG7UlUtQADQnPOZb9DwG12
PRNF4loQhlbaeSl506np+0pGZYupsVj4R6ScaPSQ5kBaPebDN2tOAQOqMcZ3T24k
XrjSie/CIPzbrMvPp2Jvawzg95/6CCtd+xxpCUEkDGrJYaFwdcRkwQlHOMsWcF/q
a6+kOC330VCS6YMRghFanyFtPUrw3ALITyspbsmLSHzATulqLjrGZPQHfhd9yut+
408IZdYLH6IaGYyNPWGhSn+7TI1XYaHw/OeiVPuivBhvwwV942jGmooj/l9uqfqc
WBeMXh9fCk03TIdWtE1bxr61F6gThQkgkCJs4jORgmfhiBC83ZjS8zsIjOhHp2Zm
VAsJ2O4aR5SrdS9/0+h3026xH8hsXbtf9dfud6cZo5J9pvSdrUd/sbSwYKZZ2g4m
J0FIrGg+jJtzu8qFq1GLCX+eZ0drc1mPjOPr9rbV0XtbkhZY402mIrnIrtbgYiW4
mmG/trZHcTtGoDo6KbfViOJqRX/WpoBKf0Zp48Xkew2atuvt5Wc636RUbrxnNM4V
LjCs/kNFDhqIn9AUosnMzFlO/b6ZHKEJ8XFOEX7jkHYsqfRPGGiXidjYRDpmfQkX
wJLKL/RMr1ybfEiE98ArZcA75vyulcmFNQrsuKF58j+6raz45COZh9KJ8LCjsbIX
m98BSD9ak9bFQ9PhNGNef2qPus5GMhp0jWtBoGLU46qCvFb7VXarPLN7TUuJB9I5
+Vtp6XQ/Anr1zA8AVg6uzUFhmce9/bC0lNqM8evJQR/o2XqyMtWQNEvsWl3dW5/o
6T6b8H4UAeriMRbIzkLSfEUXtbtPCHJLXzDM6QHlWjfxYVKz3B7cD3ukWQPTIuNP
gbx7c3Nj7n/Ncj4UysKQKx9N0N9c8FMRJ3wKTsw4s4wtewPN/pap5ubdMolwXtuD
d10uGkfyQMj0sLxZphQl6u3Voa2kc2bE6kWJxjtA1H9npu3GkZ/f2W4pP1DmKwEA
N1YTDyfw9xD+SM1J1C0VaXT0Oa++Bpq+Cnu38z4EdrW7sDd5Tytmh0H0riqbq+cX
4Z/ZWo/dTpgXqdyLPwMyvS8IyVwhxeBO8XbK6a5T6TTBeP2VjLFqnkjbFkvQPbLN
j/FvT1Tba0GaH2Gtkl3DXiXZdKJlzlNarkmu+DAnNSUIn+0KkgPvvJVGI8BgEKVQ
e2Vrzvx5weNQJkSO/LEDQBleohot+HApU8ifZ8W3NIhX0Xw4Q4mFYUmllrPzoPkq
/04AIv9XK8VlQjud+mDkgrEMIF4Iej1PYHdMrhioUnRntNwEE9nVcw2r00BdUePe
VYoTArhcB1F+yyluNNzIzgqc7m10+KPCstSNfnzIxc0SmZbWXo844dO4kcQCtk5/
svhzXE4HPu9wOzKJcIeLjGBfhrg5rB181NXoRRAYESSY+C3qCHwCMh1kCXQl85Yo
FbH0JKnMwhTYpx8blMFheaaorzCZpPxQu7WDOTnAPA9LsnbP2STYKDMhBXUAJOgB
o/1s8qqsA34dZTmQ0bCFkl7ug/ftunnKjiZ5WMOmANfQFZWkLf/Ab8AKNC8z3E6J
m6KgmwI/v3RY8TUI2ZLHbHsilO2+aqXsUwWlperSrFra0Lm0yPSJszaaYVll6Ggu
XD7d1Yz+mmFAhbXtgdTrKKptR4jS9XbfBx+S7DC10GA+rUSVxIvsCZ7cGI5fkQV9
4rmxXTGxbRBUhbb9RyFxVaRFxAo2rmK7Dol4rPPMXtSoq/TSGWUv37pPwjxUFP03
LncASCd7zWZnJaaMOk7+Qx8y8xYZpOoaDg54ZIHsb4cy5zxVkG/9eBttFD+W6xjz
3B1NjUSPP9SyisWSvkjMYkk6jQS0WqG50Z93TCZvmY30l3+6VaDwToqZKXr07k2x
l0xB6iAupkcLepQY2182SX3mpPaPqXxWfqExNnFZUDBDld2AycjZ72f89Ukwee7V
sB9b1GbbKWI6anB03Dmmu8QwkWAQjp5gSP2lZ+aGJdpgRngE55Xf6c0SA313AgOP
LIfKRMDcgsJEYlLBwSf3V5o5yYJb8p44tDVKt79CcHnTjwgfGVcB/6Wx8Ca92u1X
FHwGVHkAuH34I814NcYEsdvTQ8yLo5WINjMm3fMDysp7HG/cRqyeHozuHfJmOIxY
M6ayizykryN/LsTfSGC/LzXbV2HdCer/r1Yzih+M6bI916Gsp9wV2G8GkDjbglZ+
6yrgqTQXWZAiMvggOz3oq9tgVhQ5bHa4Y5d+kv2klmWJ3P/kiNzC38bhqocZRFEW
lv3ed+A6PNSl0u10Jt3xWL2SND2x7U+9brbZXnBUsL/mJiZQR+bR72w/PUNT+KIY
yYCLPy5EGp5JUHVfeFUf0490bTXB0SmkQSbK6grErbTRuIIxqv4AhJ/2fhh/KLJl
XHx9C52bcrbDaUbmVj6WDfg+zdrufJ9achcWkI7I6+FPH3rVrWkSFyo9msko0229
0pe64bzgyO6qWLFFiJyQV13UljtVjjB5vCaH1v8UsS024zmrdRfumPJr+pz4J54G
XaJ7UTVLn3M41P0mTTxHhg30a/0FqqsGEBCIIfDXm+c8xnd+p0HKu8MnZZy6/v1v
lnCcEQh1v4Gk6jFBJIwE3a4vd3J5Xar8K5kVjwO4NGAIudKWg0np6LTtKwvxwemx
VUL/O8/SixpvlX7bZFqzk1sag/4yCYZb515G505ZKdi+5DH9J0zd1Y4bk0/VHYHy
3xS6csC/Wgq8wlcuemafCGjKBDwV1PGsKpeaPYEIcX7KwExuB5FHKCOcnixvDQN1
Fqgm6ny1R0p2d0DJTHFa37fqWUnJnaFwdC/HjcIcodpFcEDuaqcKc2nNm2CBmCZv
RdRbF/gClXKymOsHKYZtOsWBSbAewkHJAavy+FlzYd9dbN3Wm090USBr9A8PaG3a
BvYSAP5nMl7J5h9RNz6m4Z6pV2gm6gepYaoX3zbUaB8dj23puBK4d9Wk0kp7El8L
DLvkA+rQpN2xGdCAc09beSTHZKZ+v4by5NJ6KyuFNLpVViCON0LB9KdQEEhpd59J
5wYUM6UdGxYYAB93YMxuGnqz1q5uHZR1uQVRTNgIIoD0HCvny8kkfwNaTCPKk5Ql
x5oXyNZnA79S1tvRf55dbEdtHHhZZeI+LzQTHxOcTeDk/ayLjjWJQJtJTRwXcoqJ
+ijhGQnHuszRNde5/YfiBw0gqN9zxGA9hAm6Wu1dIig7I+6jfGJ+t/8dU9VqSWMN
BKVY/zcnLgTpyxpgGvxpKn+usYr0PzGBaVhEjaIT4v7mJru+ctSX8/CEoccpFEz1
NG8PPAqWiwzhfkkrec6COgSVkvIFdNlUat4avmPNaLUJZ9HsM09U6+Asx0wPHeaj
BH2PU3F+gjwKiNuMGulF0q13fHHzPWs5kFhhfO0cWUErm80FaEYTVsLK1bDUOFoP
J6bAg+RKh09F/g34Y+0Da2Q9mlVyeg5nDezjT7DswIii6Zng3CzeM/PEBZABemPl
X9+WE6rn2ipa0WZbspDOxmYiFqBbBxO5/S+KLcSxy6hpaqnyafqSra0iX1nKDYX1
gT+xC9e4BlauaGP7g90SJk9YvsVCCpO7TQQKJYMEprkeO9vTY7ebKuAv7iPNJR/c
RxAQixhcLwIbHz9bRvemNteN46e/ExCxpa7HDeh33Ajy12LQBwFiXeKP4/dtQbOd
eBcD926N53jbKqGfQQ9gquTKaPdZAsOEeVTiJEK7A4bE4juRYukFGXTEQexB18sN
RFhszY3K8wzm5oMjpqBiZigH1mo0iWb82k9bwwgRu1TPa84lQbSJSTBbwUQV48qV
qujqaL323osyeA2MFEq2eG0bTMe97S0YLjg/m87iNZAdxp4sMl0DvCbT8N0nDROn
FKeyE33dCGlN+7pcTEg1wdKkn1FbqRpNNVcG3S7lHdU8rtkKCoq3wRD+K7Qce1O9
ciQ5Je5QYEmyLzKEex8eNcGmk5N4cJUMN6NI69sMnFdn8xv+ExVraujNAuLMmjuM
qPULQpMrHmB04Eio6VXjHjw0EGYzEseXa+ZwmRo/uvrW3Ou70RnG2GeJPbHeiwTn
YifiLiU9w1tuFobdX/H16cYthjDHzOxlFEylov41ZlIFVPQRzqJoeDeAEYtaGx8x
Pid2Yym9/VUJkK8A28hVSKJ7COJ/eKfwAMD+vXIKnJxCwlL3/5MrJ1nDO7uvmzdM
8eg3gJ/5JMTymMDiuku5eXvCJcsbzKYZY7DjnITz9sIrKHcBjBQYFkTDwK9svHil
K4OC3yihuQTbFugZ7yMY5VrGJuHear22wdIFZtywm81lodve+U2esAmewyWiEBhL
R21HkgQRWNXOANpAPvw5RIO/+t4kASZviFLtmkuO9Z8kh3O1qFPMynfF3wIXhfLe
ReXKxtmUA/TVOoBl6b4ssr6mRL8NdtCewWbe58UgK0wcttDtJsXAW/RyC4t9tl1P
kAuBG4CSu1lU3+U2iGSUj9guyNb+iCMKotJZoZxrWn0rqajVp0xmH25Qqe2j7X/x
iVySDpos0MhhRVzr/FYje2DfvLaEogU6Ek+uc8WMD+sZJyUjGHc3tiMpnvhJXUX+
hIuZMD64lFiuCKwHyWdVZCMAmMDKEMbUxX+Kgu9mFoLm3pdIbVqtEHZ2J20FpkmM
Dnz/ED2Mx9ybK/83F2xgSaURfjj8takzYaO2aMCqPRx5pwW0laVUwjKuEfTm8Gdg
+JR+kHMSZS1fuKOOkF3DCbH4WtHzjKhC/I4CzWXtDxQ98kKmFYJ2uYJEl6SAhWAm
MXSXCDzFa0gOAw+O6x6KrIOgoolZjWGT0XQQMp4RYyYop6c6CVa6cdreCHy+/zqg
MgrnS96+UXYkgIzWH7SwPzbEEHy8603/9mn4/JgMNXIOkjs6JXkdH5rK82tB6GxE
WWgPXW9EHy2ePQYMao4Ph0T11oF0XHU61w4kQ9hEtwbvoLBAkftASgQWHAJeZr3h
8yZcvvmBbIvAdqcm9pw3X7OFlLHlOLblJe/waMlyDBZnmVptCVQr/AQCnI6MgWH8
0BkO80K3PGEKwp1yCmcTMO1UXWgerVt2HvGrzMk0Hd9w3oz9/B4aoRnhfBxIDMFY
qDp9txBa0oawJ0LmlFyvaZcjd+/qAzYG7DwkJ2VC5VkRRk8fKKy5i1ojE2m4Y2lH
drlUcM5pdoIk01Ek2xA3lckRuccpUYdrdh8ROdxrXK35Wa9PfMbF4WFlkBXB3Hgy
kh/NNQk6nHKKKLI6lCPfUSlISYIwx9BSVDH1/r30hJlq35MwSeqbEq/5HlUpQDOs
RQR4uwh4COHYDuv/aNIZwW2jYCN0GuVUdsR/OzjFaXO2nRW81FD8maBfMQO+iNKG
fSGS0T2v90cgZMu/QhhmSUR3DUlnRPMFOCMUQDxtcP/1ylj1Y1RQ31PPESmmOYrj
509+JGCjHsE+lcoZ714S7vGoP0WLOnBvFRoKcOyUUD2TECncrSBdASDDwxN5pMXD
Zc9v4LvbI8oJqjwcPTN9QcMNsAep2G/lts7i60KtwonFmslNPmH3tNQzjT7fQa7D
E0RUbSiqF3qcGaZKcSWX4SR+VHpaY8lS8SVLYeEqWbwueaWaf6ORg1d4egwVAm1C
K3PVu04ijYF74kmB+l4nDAjlUbJ9Vm/H6yl4GfnUrDifxBSCsSj1O05Tztvtop2Y
/M4KeHBQDA6w+xdSe9kEVRjKUPMmsZw7l36vWozmBj76tF64oIhtPMafhGH6Qwec
CmoVeur5MALUbYphFoUT58yhWDpMyIDtsWor1j2Ag29bKvDxHuZ4PHiSPIHIHNAs
tl4O1EsBaRWvy6LMqLnMVVULTvMeMpzCrSZBHiPWIHS/NzgedBgtU9ZhTYZApotl
tqSpVW0HrZhjkXuWNOu6EQNjRSASh4RhJrFQlG43AO7zUfIkyXSaOqdS5B02LQ3b
7FLCMlsQ4ZNTyGp7/9LnuG6l1ykdz/VqX2qFIw3frtaOOcAqx7lbdCEAaHsXkOtr
FhmkSD8iOh+XxmmMpZZSOEBHUNXVzivxDJyaQbdCn1qRmsAml7PB0TfuLk2FBqtK
NzBKJdz283ZUI1nr2+OWfqa4dN2WEHSig4KvSeY4Emy+M7mB69YilUSSTBBBv+1u
wy7MOJPN0rVx/YltA235gQCip8J1yOL75lNnKzAnLZJg1zwPa8uhoPKtrOWICSDL
lIeKOkrs9IN9zZOmjh+nm7b8IMBxH0akr80p1VCYlEeTyIHd12qrNdsZnTdrXKMT
MGx/djrmL5RiBLdEOnZkH31vYPq9ksaJkpxJ9mIZl5qMLcA3Cv2U2dWCtjWTdPVC
dzeNqdKTcofsrIe66Gm+OKfq4L3Uff4gNR0KQtBuM34IEsRJOQtm7vjBYcBXLtrl
qC7yeNhYgZjxDFcMrG5GdfSodsWPORKwl1xpNpQ/38klieGHiecqrLjRGqxXWyT8
j0RJsAhh3VrJ1L4Ns04yLjLPheMWwsJ9ayjcTj9yRp9jqhceYCjoV8uQd2TGOzv8
LBZIik4/Ah4PA8r9xcc41dlTDPaFMV01pVKf/Jq98MRGH8xF2Fz/Gel5uaQqmgPg
11TLEDsKIJ9QuPPrkvH96HK2FpUXUQq1qB2QF4A4xuSHaX5RNQHDEHr9Xsrtcsum
1evZzd2xCkPZ+Slud5HoIDgwZbIzBgnYESdtWC61OMRoDx995U8FvoLbDwPO9xu/
y4pfNamHq9w2KToEu9PQ2n6QpUFDeAjNANuNGrsJE8WoXNQMwcp2EnGm4+8zxljS
9hDznYsceOLy58pJp6YyCcOR1UdUtnHEVNPu4b5cqgVGeypMvwklGZbiRoOqBHQA
pK7rMiEvFIFq6RQ6ZEqL3/OjsHE026qDWzkxv90cU5cLATBbwIKLnA4UlxjEjwoK
3pk00Rr9RrZ2YMWIBj6kQXBLK1urcohWj8Ve+zCpaMES3YeK5HAhk8FxEuxyFec/
8CsB3XvqylNO3oF9JhgnElWIPFejmKxEw2BXAnM31S0Dy5SZoL7GT8TYVWM0jq/c
MZW2KNl7wW++LuypWIjMpYr87QEjkteDYdEvNUsXEqbC6ANWbUp8FrvfYKupVopt
p6AhvY1tFpgT6gTY54UMt/n4iyd6Ii+zp8NdsufTz/WlIv/IDgfzf5lP7WS9rvie
dF798oY5LFGVqDfvlw0GSyaynJtXZZyVb8/Ft0grYgzqSnJI14pwE2vvE2VaJbmf
H2Acn6iNAg0Rrc9W5Ukzj/Yc/HQgIiUYcOAwwRxrLljPP6bgRkWF2H4flM/w66uX
SkwTFTJpe6uwz9HZhNc7tZV+WgLHDsiX2Gn1z3PCMVaJ8XPxvwHjWWbncrv/lBjB
oapRlnY2rLhibqRFT3d6FFJDxl5LqQaJPnOzHheNu+dZ1W+1AicQUKXa6wxo3BJd
0WkwBsM/vk6Q95NuVJ80jFRlA36IjRy38abLWGGlwcrZxEJnCACMgSbUueaY0Lh9
pMm9fK6+xKUzfzI6wjxFgYJS05lrR55MNJbC0u+Ot1KB/KOKwwA36DIy2TlsbQXJ
3EpSgOIb8lxy65Je5lgM8xmtyfPaE/Hqopbkh1kksFLyydifVPbz+j5hTv7LxDR2
RWpsKibMnvdcVzR+8PFt3rye2f9DR1gLsyvADZZMA3n5jCbbIRj8GJqVu9W1mWx2
buaKNm4H5jN/Gzo0Bmb9ve1S13QtA/hGrmIjOs1fWHYOfOf9hFqCZloOxbDx0z1V
HKvpLo3ktxPKxo+R2mC1zxKwMUKyBQa4HvXAkMHaakjxwI4nG4uV2q2F41UOwhsU
h8mVf8R2DN0xrmAm22bxHOtyiu5xl6Laik6UMYKMvH4nZtH2xxkeg+omGbGnjpuJ
StRktnyXPtSoQoP8fL5ftRB5AcrO7H4PfWnUpKM90YcY9h/OGD3G6SNs9JERrLCj
OCtuXWpAeeeHE/RmlFhJxlxR3asBXvlnGatomJiUz0LDshEmJ15Hor7q4tdWGTcn
3vnNHXjfy/xseXocmzhtNn8+Xu/+EliwKh2iwh7WAvHzCiZWTja7dcTJ/lIgVOfn
Qqcr+rZ1orBZT1AKjdKAvF0ZsPtxc3ycFbS/BBxLMYdbQM0JCXH8qDm9mN7j5tEe
TpatoIqKGWysKqaw7vJ50iENR+g/r1DdGr/nD92Jrksx86E+vN8DDqdn7lPms9pZ
L0DBYCFiMsoyvMv5LEayCA6aUooe5lIiiBuJxJQKwJGYQoZ2QWFjJMHU1S7inIGu
wrIq+CqmRZYZ607Ow0Ga2xQix4ccn7eOnMRUVD+QqjkuWgzArWTHCl3kczz7Po3p
WownNmOMKi8LjsoHZF/OC1gb6mZCcD6e2xu7ZqcdB+fNT6oBkOMqiIk/tkIONUZg
Gk26rqIgiPxbGxetGZAvr39v0LD9YvYH1NmFywWc0PRnCuPSKPQoov6WKfLAYDiR
SAzDet7th4caLZNNbm4+62iJ/EQlFCLcHKZcWvJl14XbAZR/Ac14b6K/zuHdbEBH
VRhneb+r3sUo7DGENCbqci+o89tfzuKLMnTeboq/nGDmxrD/Xf2skxgPZHB2Uz9Y
oRQbCAUI+4SSzQf3/xlap821KlxSrdUfVxjEh7ObZr584Z+6PLHJzgxJyjQKsyQh
Y2ODogCaL+91GIU8ww7mu8/iMyUT0NaI4icuSwHU2B4oF0LYgAqcTOJWclC5hcqg
2mUCweKMjHRW4+Prs/Hyqnvc289w1Meko2VvWPU+lEP4RGkQUf7cwoHsT4c9+KiB
nY7+7ZfQ05bQDqynIDxI1dq/I6jQGOR7cWhZguG7zLNwjXC1sKyBIkwqenfYXNju
qonA7fcE4jNZ4osKB1icpQOV5D9mmQmYBTUQ2UWSQKcx3aVe0YDnPqrjOAezmKqy
QRQwhvvf+ko1vFqEQ8dXrIRmjH7x6q2ZVSJM4k6kFv5jDXHuIqcjD3Z8r5pqXNpL
Hokm1NjJ1U6cJ+KK9oKSomhr1wv92DMH0x37v6C+e5KvTG0cLNaoj5wJFShrFIwg
8NRsHxra7Vxl0NcUaEqem0hZXZpn09gPYGMAv8dokoxaoS0W8nKqfCRvaUQsgJol
4nk3LnC2tFGArLlpP7+Uqg4StSeJRr1l8VLytOHT8haALWN4eBEOzM3aognYXudV
7I/I5Z75iTB+JQIWgQs6yw3E9Qs2UEFPfXHQLVd09h3v5PXy74YpYVdhyCQvJFB8
cs7erMXVERIQffE9mQ9/5cQQ2sNOTFN65UXUlT3HSXmaBvl4HgHKrqiYIdRZpZqB
3epFO+ALAzyQuvg2qdtQ8OlpJxIrYdfCfJk64cZdt8hfqsU1BOOSZ+j3JV4ammmA
vYfAyzkGBnVWkfZs1AWwK0vAoe5pdvcZVzgT14rPJ7ZRxrMTWGWHcswsycXAliLL
/buvHcAJ2pr7I2l8TdL5HYGbsnbtiYHvypk5GhyWMSxcystZxPJA8xRXJFTfj3da
wveRd3/RmJJIJmZozUbBx1yWRded27O8sCZw+fmgr9GXkERaxLGXa37y/rTNGbGC
Y6StR619ZUcrwl4q+n5rijfCSYznWapyPEBdmfxbFoaQ8k49n3Jak5n6U/C0Q6SZ
wZ9lGbyziLIe+pSxIRAG7NESDioDs7FRklWgUoGSDeBmTP5JG5qw12aObTyGJuLQ
bkV5KeJNu9MT2ZzTjYzH0j3f3jiYCbAd7gHZO7EIUjPsPkFkVoV0LL5OQcTuIsm6
hxfNUD1WUqRIAYFVBhi4igdt3dXfmkMTdP6GU2A+blt3LqZ+Ei5DKPF7DGBpMe4O
Ld4nxJBGYWsTU8CQaQyatXdasnDGt0ctX1zG4NGuIL4ydwOfvSUXLRrXO0YIlsKD
PJmV4ixhSi3Dnnue5nMo06XLFz1FZtIguFE1VquaSbS4/eJRspU0Qm6tr6lOBrUH
vqb8x13/gxcX6KMDekF53qBFIAhUWUWd8c4k/rsrAZwai4vGSI6jUqduNXoL1MbX
35y+OUnHFozFfg537OWQjLUq5Vh4rfyVi8J324NlcctOhgjUknq2tUPfS5OOffMv
x/QAcReGGClG5l/Zx+Mjk2fRXFVA6WlCcIwXckz8QFQHLgeMyArO1e2xzyzMQhrH
MfOwwpIE5SbdibWlcCSo4IH83iWSXChZmLn2RtmxZnxIzukwVMWLIQc9PrwDiReu
9Bt1cNHil48A/rne0lJ1YtrbXkeUk3gMAZn5sWY0RWRcfo51AkkKdo0RjC5AeZNu
uMWQeCU3GBlOTRVzICCPT/eDOT6aRc6w4XoH2c+o1sDNBQ0TqsV1oB3SqqvtBCAR
uzVTAYAlAHn1h+olMYun8/eno63xg1S69e1s8YkxOyuzIHFPwx+PXFnbT5EIF5mZ
ohrSHw49q8gY1phNWcfopTK3BEgrzsHoGNXNIMNRVHUb9TEwj/t6ntwHcqu3jEQp
cqgL2v8oSiNWvQdaX8zBNFe+oDN0eu38di180I19PxsFYyhk80doP3lhFSaMiKYS
hOHYrTZ8ZyEkRQP1o0sYKUaPT4w7o86DlfKQynN6ZWXbwXieJSNZJZ58BHLxomSN
ygLIiat8oFAaDLsgqPJMxMpbIYxzfSbdMQziSeqq2kDzSxWC/+8VL6z3z9Jt/9+X
fLhbeOntmkAAKkBwqQie5/golSid/tnAR5Yq+es5sk7r9R3ltNC4dxHcoCJYTRbN
IMxzwYFeI4rcLrlb3JCJ7VkIE9H7KZVPjuRP0tW0LIptNHLNEzrsJ/UAjqTODcQb
DVSi1KC6x71h71MQlgc4YJ5UVqKa4XW8v8djhADHGJRlqEXCBBdLcVH9qCos5gpk
ir3eQXlrtIoqr7h/faRyMV+BkG8CfepcEiBvh/XlADUS3QqC4tYC/VJ8unNAmtoU
2i/cS2QHbIobMYqRzHhWfv7M6Uex70I0oj6j0SopMgbdjvYe/c23/wAHttCbPzzs
j+WA4TmsNtAFaCMApQaX6d5QvUDLHkxtvacd2u8Snt4alAaQgoHYwj2LiTRsDIuI
KLWVkrGBuRHVGvyeral3aQExCMhYrmq9SPa94GHpq9/iTJs+FeHuo+vbf/G72B5v
YVTbDtsZ2XQ5Y+xrVR6OPpUXC4/y2e/wM/fkAEUsLh0jN+7SUsR2zalazFpJaink
HKvKP+j6kmFak1zI76GLRM5T3g7C7HfdiMQgIi6nES0=
`protect END_PROTECTED
