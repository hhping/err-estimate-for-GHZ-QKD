`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wq5vFeQTUFJDfMjVxLf67myKjbJixEN895FiSjBWsia0cp7VIRwPxCcNbEIuxsz0
8xN9WcjdY7Oj5nYOYw0YL4ZOm/TWKeaaADARYbFaB/MOpPz7UH2npojxR0bZf0a6
3YeXuXV3PCg1qomzUIMBOJddLNAUUfEWtCEfkycoIU9yhqnv6bqFY/HJNDV+4GmI
pCMzE/EGSoe36OMDu4w7eBzt6i82li3e3mic9MhQ7JaB2vMRza9BqrWDHp9/okOu
Ph8iR0zHRjCGgGn3EV9WV/G00dr8M1EOhwZ9sXk/iOg/LJsC43h7wuo7b7pP+T2u
d1sccrtXubzdiHF7R1NCpImKMH9l3/SEqo8b8VKsM4yt6r8wt3BpSj8BlxDvZnqJ
Pu+PnbzcOFBtHg++dU7T8q44r3R2xYnIYWYofNzQpibQB9rMyxPXh9GMQNt248Lx
3DcERp9o7AVR1r7wTHXDp/XL7dXDF2zI1FswZlW10WwxpHgS+xa/g7hSJ7z52sc2
nl3b++hu16SANXbW+y9R4POCF7WhE5ozXopNygA+6I6Q+eVxd9k+WfTQf++z8Szj
iMkNyprulCcCCZ1fNHDYJ7HyEfZcvr4YdYdPBsxm15aySunrch3tnqB7x3ENB2X0
AeI4CBuMeDsDzj7A0MHJxXqRUPA1RAueFwLJuSwPDNjVrlNHr4hVSQYzcg1bLEHk
SAIGXb6IdxntLMEIF1oM3dJ4mManA9wYMMFWwCAYKVuYgMya4KZ2t3ZCIU4LHMA0
p7iB2HlyrNcG9JanH/mqw44CVKf11baQGN6Ve0VbKxDgxr8dY6oLXPEWz7e++stP
RzLqgG+8YGkQ7Kj42lAcP4BH3sll+16K3qmHQf4QvxfZqEq/feFv8r/RUUDeihrD
5p7e2cYE08eC+IRvGaBAtXVsCnGElAUtWJogT212/vnnnIEzjBC6OeGuzF1LuaFy
NS8DHl6WRMGyREe/Lb8ahSU9lBJDPOhVqhKh1Df2cIT/Sg/hQ1x5z2/qqtUMPB3g
KSaml+xv01mW+aP82ZVVy8qfmRgH71uE1Xyv6UresVVBW3yLavp93T0NVnJgdeTl
xGa9eLwN//LDibFrpzwv64iJGkBbv4wLkqKp2eErXDl6lf/3yHTPJSQUCBDzzIp7
lXEB1ruBxW4r1nA9dJZV5eh35Ka193hrcZekgyHUm3APWwU2D1CHd9MGoeis+NLi
jUggDgSqajcfa0lSo5N4NdzWryhyvobn7yjUSZXa9nDILQHnYeKfMNwfUs5BY1i0
TsjP5PeisgvhV8ypRQmk8EYQhc+x2nDxwlM5WPhL80w=
`protect END_PROTECTED
