`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfeYV2ASxKByZ/5C8BBPP/Oi2RksB8Ua7wSHFGmkZZwwz12tTbsqKk4toq1krDQe
/fV9rFzJyF5Z9uv8ldDBjjPuTpnkm4bphZ6OOaTN+OYa+c0UEOLEkXmqaA8WpGFe
2WgH9cdACVd4tScCUp7hMnbbJUWtjU+ef7vsEpPP1UAjZSdkHCZp8Nz2tb37yY5b
HcqvB+AHtLeLwbWtPZzemKkYKU9wsXdqyWWXAvKL72gi7GsMryahSkJC/do63ATO
D8AHSc/Lw5dg+plH47NeJH6hhXhIqmMj3aZjCHURBs0hVHYStnatO3NWQUBQwWzh
4v7knmW7H4o4p2zFy3EkLw45P+xYrPUGyZIyEN0XUxZ7DwAQQQLm1W1oTImqkbSF
gYukRhApdBgIRU3qMfGjcodg3iOBfmMojF0y8uyIWTwQ3tatgfvdEvK7oDYKssbq
3kjiNKMrAT8dqOAFJDy4ILrof7TxHXOwCRdWJHTlFJ/mjFEBDW/AAtcRiHwFLjvC
WkR7Hs0zyuD2vRJ5bXE4Z/Z1w2SrT9fpun2pN9dt2iPwZimNhAlBUDDi8QB/uXyi
cxw4ytmyYjmk3o1knPIm1PW3RVEbviV0uqCjoQJ+MEy8/2TgNcPYVBXoJAvlF+yr
rrqgdryv0dxoNZOQ9uzZewG1XG4UVgF/tiW3+qnPkEH5xc0ym6JK7qK/zSKr4MiI
OU5igw2rLZ7l1B5fCcl6+W60r0ymwJYaRqF8qBiOloxljUA/FXTFm07BodPswIPj
pYkQbaPBN4ZCjF+j4LzBlnlWy6aws7g2PVj8UeEx5EGmsn6vDapW1D00Y2oCe2EA
G8qJhloi5TJ8/E3pTDoJnyc1Pu/YbsmwJelxU9H+ZvJHOPpuFzqyN6f7u9aaconL
SZqs+tTZvB3cJ6ZLtYSDnfR+sNsCmo8neeC+kBeJLybz1WVb20ObFiU+CQAEdoh0
5pssxwMNjRNtywoNT+adHM7sGPYe8x5xLHjqDEFNqC/uPpMRVGu7MchUmx/pDtUw
3fLb9eY1aoIlMJdtlCPCzyPJcpol/OlPt/Sz+a1XrNO+Wuh+yCULNei0FA+V3T7p
irkuLp8FQ4TffrhqCVhFEBxo8U0mupkQth3ceBICwJsXZi32VDmMF4f2i3N1j7a7
XKN8lJ7matqhFjk3QSlmwLmraLvm6UZXQl0G0MzsD8uOsXHKeQOgXILPnMWXicgJ
JBCagYMVZTS8SdnYZXVIMdmD38JlwZitT2CpKpEMskU=
`protect END_PROTECTED
