`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1I8dF6E2xMI4GQDW97D1wWQjxMf+WPDCAT8Bf1QWToLyWfOtOEkyjFYIzpI0f5h
nsLylN+gMkzI1YsweQj4hATDaEbD35LtH/vK9fGbOIr+wc9YZsN9k+yfl/OMgpYM
Gm6fL7B0j6N2nsAhsufzuJg3hvOYGt8lArL577qGeHGjlaHm+bsoIZuq6Rxn260e
PI4hX9gDvDm+iAdka8qk4TYZGv6CAscBYC/2+WW3QXWJVG1v3SG2GiKcNhoLFTiL
YYdi9LzUS7awfI3HXpRUO4gApUjReB7dj9hEY0WSNiUub9kECsBJlcRy6MIv2g5n
/ePJIHDypOkErurTuPUHi2I1WSVQe1/SQ2Lniu/2h2Rzkis0VSyx/ulqL7vDAP7a
F3i/tsUT4uRciNzmQq6YSTH5ajpixl/XRT5z9e12Z/TN7xcrsatkQtCDHLgJlhqh
C20Y1IQqHhSCv/COBp0+TknA0mdfOHmek+rF1om/K7zgjDhUY+yZqdUcN57BkC+/
gdB/2IfACg6CusZy4Owh4C8IR48wlkgg0HcnkXholJaMSLFK7yJf5xqjW0aNHLqe
hhHUJohSvTSKurovx5eddDKJjb3NbkHw0wZIYpwulydX56Q1sMPIrFv0hCJrWBZq
GPTvYrlaYMMDrCiJynnvstFabhWSin1TPbYbUkUC+E+ndZ0kh+oSpm9WZESDkZAC
2K1bL+t6TMcWXlsmawVZVz7l4rhrjkDkH5SFfIxybviojNtvLzEwD5cqKVpx5Ipu
JlstpaDMr1BTgMhPmmzW4Ew/7QisE/+UZtELcIimrTef6YXJYcQ3kkh9IvX5DrDx
DR9fwbwpYuVETvcyn5be8L5ysD6DTRjOU9g2e2exf6g+eQDRe47qdKcuv9jLTnOT
xmDAS41bIZUEK/IPjK451+1/dKnR8Avaz6eUc/Q2ad80Ju3P1Gs3KQu43/2qkRx4
r0r7SqY12XJSD3OVR30KmJIk3uTzcn0GiIRiMDiuIYvN56Hub/uRl1TF8+rRUz+M
qiODIIS0VTcsB0bbDfOwOLsSX6GqjpfEP8QyAwmqa8MqDE5HF/Fwb93cxQY3EJ31
GfqGMBlzL3P9/PzNZR9yPuB4hoKHVh7JDj9wwnQJmSsATdiZSpAmHaTqmL+pARep
fiWZ9+xzaeshU79vhzmAXd6HJSyEM0Qb3MaP86xEmGceQxb0Y5P6gp6uGsFtq0+T
N1fdweZosxlxZKkTbHud3unt3YEIPcXDr8sGnKA4n1idaW/xaWZ6UY9MKVeYQukM
XEN/Hj7tZIiyCrEO6TqJ0EpCK59L05cB4gp0squT74BghiZL2JLmHoh6qj9b65gL
rrroah1ROCrQ+pnD8/FhnTXj2PM0RBPoi8hP9a12/qfi4uxHmu7mMJy/yl5dW5wi
AhO++tALHVHGO+1wN88DIrP5fYyRHxNxVVyDycaPTjAfjlEebef0B5kX3y6sun74
nOTOI4Xy64Wj5MpIZek6UL8vhIshvrckgS1IKjFLxYcWdVtz8DFxYCsq3rsMtO1d
qyTiEehrzyC2TmV7eP3sTTIkyZmOCxXmUeakKXlplZpzVA6m5dfXvuUly0f2zUQG
gEUgbybLaAXEXvsFJEo1CcxYsxV0zRtB/5vwJ+47jHw7T/Is8osz0pGOFq5IYDb+
O/OjunWN71l8Pc47FYjDmqItYWgWC8kqEUMXTGmC9w0qDKeYbiwUNKk4AX3FTk2u
yxcwTAnmrv2c4OVlyItsOOutyDJ6K/FT5vYCmM4yCNB8virIjXIu3Gs/G6Kw5EQ6
OoMxZ8Der9iz17YFtXuOeDV8dGnum7SOzOUIMSeKINuiVJfVpdwZwPAFm6NuHx2j
jQpqFBXl2zisRZIxLwJTwa6LK9b9oFtzFQtwWwsCMKsaqgi7mwIZZ3Pirgrponcx
lrnX1Jeb/By5F7QSdH6NfM2OU+zdRjWtVJAzkcFryW/NxtVfwWp5V75w66K/0eEr
dK2EhwZAdUgP1QEJsTk1ZQAbkVFlklX97EHzF2yYu3nuVnNQee3eObECBQl+cEZj
r/kUvY6zJwqzTcAhrhegVd4jL9nnzDtSRrAHcxDnWZ4QKrzpPe4VhqJj9LFJams9
69SpGrGs1S56qEBPa2GPaGGVe4Xb0WjhHLpWzmLONCukfQDZOdNWlD9ev5VuEeww
vf7JlecS7+Tgso0+LNgUSzqcDHcLh2czvq90MQjA3s3W8uHZJMcX0ZPxHz6BHg48
mClHqmK8G7j2N7jHAxPjCL7aaHthEv9WA+iSGMDqqvK5M+JlchCbrCKGaQWXaw3X
afqwj0pQ7gNT3jbGSOfDi2UsT7lgB+Bm4X12Zdg7eYOC2Q/hUimanJdRsuFsLfN1
QkmoBY5FK0vGzcX/3A+16olCfUN9adn+PJnSpuOwaiixbtzVof9VMXBVOuvHiMhw
eVmSo52+L2eWA2DYMHrXlWdytJ1c6gAWytbtqXa60wzFmvb6LURQVlXAM1khPk2s
O5LBxgpeP5FFBxR9v+P4q11sISPZo6B781xXAfX18O7j++hIdipGQB0+MZkvXNX2
GwqLuWzhfGcJZ6SGxzaiqqKb2ebBQCYVjzIWs9Zi0SvXaiFd3QLQqo1JS/3G2u6b
ccfDiJHFoYFUYu/RewdnNLr5enP7LWUGPfN4y/024iE4xqPVia+lQ+RnoIE5fP1d
7xCwEWvQTI2j2Xj1E8Q0sEthXoVBJy5ISXB+8S+HFMTbA0Kwh5H/ZvD74P9Fm2fP
2JCmmp0AWQLzFuO8O674iS9wmOt0BCMIEZdkBLFLfpJaIo9uho9Hw2REbOaMWHqu
gCz21aJlaNFHNE3iU6749X5aapmVO6YOFg5bd5SoixKIW8MYMtpv/wcyTmFnLzZv
ih+0fWDWawhRZDzdhpKYw/J3qRwi4Lp+SVnOK6pzhL6rlBI6g9h+FAHe7fR29bzX
SYACJmkJESERhMHFWqsAO4d8wyaX3slCj7vnvpC9o8eA0WdvrWyKFeJ6g87kpScx
63hjtSLo5LwaTuhPKld2kq0KiqKvKIskLomgEhpOkryCliDs8Cn1dl4nGc0Ytuex
KcL3Bsjwid2zA8gO6vVUVkdwQL9yYW8mo1//TFh3Seia8xDpzmfCrgtTGKx4qxVR
DP46BsqaRgb0SErlZVUo4sTmP5j5wDdsKI42395465K3a0qBMqnz3cFmS0ISZ9cQ
dqtbymVOomOPaJFi2O1Kyd0FEb+2J48Ddi0hKwO59FuCJZz3xtOvnbMbMrDsr5Rm
Tu2SBHnRSr63Syw7TUEx+OlGFjyyf1HGDwupcXW05xaUu5Y/+HIbbJA/82WfV+mW
apcZm4J4Y49H0O513gBt2zLR9oHiNTl2LUZRrUP0puVMWVY/6wS+0fUS7tDYLac3
ld9MsEFJIuM61r+58/ew9Bq0As3rLZ3d8+YxBlHTr2w2O8FCDzTEYwWOIRfpx6da
+VGHWkPRUe+xo5h7iCHroucfAv+ChZZzFrSR6F272x+hheaEWJtVVxkZPee/n/6W
Sv0lRQnTp/5VBeGA6UAB+2TOiIHX8YLSJSOVjwmBJzHXgFi31/uecFMxqfiix9xl
k/nXn+NzlqD0gCNcQIcQifbmPiqIBJKJCisfOm4+R+zMUfRIQppr+L+Eujt3yorF
zFT4HnPFTT0Y0KQkCosDVMH5mFTwcdm809351vtBUXW6xPqWivpN9u7OiuB+9dEv
zB4ftpXd4j9MgBQ2R+5F8iaSsgQf9xOo6/dVcp2DlikmGoF+eC6PNjy82ELdjmVu
tlFSpT1i6gP1aqiEvxxOz5sOC/fwQfWFNMcifydbBPu7hU8qior2asEEFu3JUwXi
eXC95md3pJ+57AF5CiEABXaFxo+W94/XWs9f+/qLUiaat67HndjjBJwTDptJXLmJ
YN4bbhXiR26TaNC86My52CfV/faB5ecB1iQi00wY9cR6PUMJ8UiBD1aWkqX+UKgh
EYm9/rsIUFCjljKUdQ0/mzD8eUp35xpf7UqxbTrJqN9wNnIA7Sz6YgzSVPk7H9v+
f9PtVZu+bJUJ+d/t1D0ltvXjsgWXrtg11ALie7X1OcDKcQUPMS+pnAEQ1Wk223o7
ijRPLfLRjAvAepMckjkNajNtVjXaOGXPAcZwyP4vNnU/I/HL6d+rBc/Qr2VKlS58
w7xIMxDhWhpNhkwYnsz1HqfuyZ0frAtu3TRycJjljb6d4Fo9IKTPGZCy2tdn0DMz
JPgxF2vHdYw/y7Qtzkzn43+tuLC97wCsnap7Mva6u99/dHFwiYShrShZcz6WOl6/
5xng+Et/XKmyDfWByyKSK/MI3ugRCUWItyHTB5qIAVoomdGP4kFSLCbYWYf1WqQa
VduIDcFsUJ7NucaEu1u/wm/KGRKXXTdgK21DPyFIHzxfn2qPM0hasODJtg4lsb5a
`protect END_PROTECTED
