`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yiiazAMH1OaEsPYZqDUGr37cqz+Ccrh9EdUs4hv8rWxjVLyo5P8gCqelsgkjU0kJ
sOjaS/pjnLzrr+ZcrDPdsKdtxx7QdaAbgXsW4rRQYpmHLlTCgUCYWGaVMuWFruHN
Ut1jXCiYpiWCXETMZd3lbIl2Up+taRh5bGRTk/pYcqm8EjfehOXjgljSSiBVe+Xk
`protect END_PROTECTED
