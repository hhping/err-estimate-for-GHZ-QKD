`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ndl04kmyje4esUaTgCI3yUJhqD1FCLe0gu4pO422IK2Q9pjHj6qVGxHp67Zpxn4Y
nMtqc+fbHtPJ56UmOy0phJhO+AVEpMu7JriUtm/KLVEz1i97VlUUIANBgw+s+xge
wzo3jbtJBZCDrg5KHXBCs3gbrJMFAQ9Oy++Jdn1lvamnfcilWRIbDAYwdSQOW8Kj
llcFEPrIySkZM22dP2c4+iEBHbnccjpC5yawtAiIAkGCWch4n2uJnlaKXVIAuRj+
5dMNyYgmv2Jz7nEyZuruSd2JNZQiVhgxTUX2QtmKqnMcZ3sG7MgrF/fhwhU9RB7Y
dw1szV2zCk6kou3RTKuXV5QkH49SgqoMFSH2kZZ+oLiM6jYgS3Hxomn8uVGzZ1PB
nIPvJ77ssL/A/Tzx9zffTjKHvd5Cg/trzzBp9nBvtVe+h9m4xCa+Mrcd9xyoxK30
8W0y6xDgAbL/FZv8EQdf+7YaUwihPwaxblfDWPCbUjNLdYMBULCVEYMO0pIaGnhu
`protect END_PROTECTED
