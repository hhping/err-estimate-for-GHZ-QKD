`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVOYvd2aICXPrjFPiXjQHe0c+sxALezrSFaZG+oV0oIXgdPoSHE4hGZRdLSPe2h3
XOiaMH6nhuvJthrL4brVmbVGGj850fu7lPTSLOo0r3zji+dT9CZOPCOtoCVf1NQK
o8Di0XxCf/jnv4c/Hm9hWfK2lgMp4iBJFUB4zaKRkA+IO9wildgREf0uTAEcAtbx
f913+XrYBqJj/Z0cm14hVY/q8zi2qVBs+bn7hBfqHEvU81kGw6ySK/S5JLo0axjr
dE+LhW027WpHlu27/WMIqGaSGzO8iUZDUJr+E6SeuPtVYykSVO/gCU6/yIDzeBxx
Idm2gO6nxVy9rXyqI4Y2c1lYUWgxlcgsL7+Sks5F5mGm9kc1qViMx9kVa9kT35iR
rmXUDVyqabp+v4eirtTjZWVM8oVQDQ8aWCwXl1Y3N7zUAAfk5CS+J3xTU4nr+Yys
xwUJZDE0Vr+nJfieDxO+j1dh6haZQPnJFNFDnRtSw6LJaiaGpfw1OTwEyF1heLYD
z8oEl10slLLJE1aGD2JBQF7hXqxv1JdTGY4jRQgTxBY4RAokQGewhPy3Vh84WY9Z
xbN2fczwr2kbV5WuWyv9k9yccAeXmzRCbHAENe8wA82YlBkHu0rFqvha+BnlvvQy
KEOSMEkcINWdFyK4rjODpVB7t7NBxzwxD9dWpE/52KYbOZlUZJAc3nbxE5OUwI16
`protect END_PROTECTED
