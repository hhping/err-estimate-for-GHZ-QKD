`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYaDxPd43gLWA04ot5Hhy6kGcMlI0iTovieF4Fzk1iA8wS2fA1Ec/SpOpcWrGdQh
O2eWEN9rpPi7pDJi3l3dYwkyXS5Ywfc6BIwcp3rG0VuD4XYD0TmW3rz3KD7O7U55
Rros799aTo6l+iPVWe1HSyjmNEOSxBphlKgxQ/sa23L27KHZKGIM2EGw2wbZ4xLT
VO8pTT3rLYBbJU9XDPP8/STcf+tTdQ/GqNzMgRCHiDFb3LUliHW0StqbzFBYYvWX
KmWCkkpnCu5/fK82HAbPCiZwssD57LShz35y6dyfWhCe+ufsEm4G5sEOB3q7eBO/
Y22qRg+63AykdJDqiigD0QAWW/wiGUCy1XIg85pvMtF5gwEtIDN4ER9babH2x4TG
tKoSjUVjv6Op73v+0hzDKWtAG5P2qMb4Kv1dFidu9fQGdRzDQeIaxyxwPuu3pA1P
lXifxNCEs+mOJk6kcH+rwAyEhNyzsXeesJ2BkxQptvS2MF7/ylymjDMOWQcCqVon
mWFj1XZ/5s2JqSdEA/hTyg7VayxcbWv6S7s4XLnn2ybC7Eow1ACt+MYbE/V/kR2O
G2b6MZtj7FqIbtwdNoPxrNLVDHmcT4sZoiOqHLnzjy8Wb+k2oVNcZUnMuLWIohkN
KguumYu/gSgYSzuKATMBBf98nKyFcNC7sjRb8IncbNvxVwtD2KNCSO+QAjeZCSVN
6lmnlnUt8GK+yPOqHjoPl2qFUaUwzWYXTeQD42EHP8N8UyEdmYX6aQU+BjTe2qEF
mXVe5G3cKULrJ5CfXhkvief80BJKTEogdUphiMvWKxaxu5vhE4fD1SApqWZ30Jug
3fWIxHpiJl/2YHYQ8iO4dvFYPziQvlvoY1Rxfzmy9DeONnBFBPrVAPa/buSmDuqw
U3LKq07M0MvjWK7dG+Vfn3T0yiFYYSuLewIAYqaL8yDhNFgq07J1Dx7WErZJJhqG
OiGHD0KPOShA2MuqUGzECM3MoDPCXmFpN/RbUDCbYE2oBEM7fBbKDJ2pxVgMK2Yh
Sw4J7zARz/qwdvI9pzV26lmNyRU97cpfZi5z1R+GbwUbLiYGu/VVVEWZg0T6BpFc
9rRu7s+oh1WwcizThbu1SWl4FNa5J+Z71o5PdQkJDnFvCxOT02JlkSjMO2BKfmFk
/2ZeTdaL2jZB04ZInoc7IuNXx+9A/SCQRajMnpz9ThiA1zqmfwiUIYIpfDlff0k6
ih1n8POrRoOYVwapGSUdJHQ4UBUOcNIL3vAnyxzaHU5DpIolmV8rSPauoJNsZga2
4HKL4hDb3Vh+kcbg7up4KqRuTJUqFpMHLkARQj0RyNcfsmXFnYdeEu0Ow8GyEjyN
jbAffx1cdjhTpwmFpTxtG+uoRWEDPL/J23GaONhp5S5yWmlWMHVgEDfep38ntdtt
HU/05CgPB2UCx4L+KMmsNOz77E/Ed+psQydsaIP7M/pOKrPsVxZR/E7KvJCbC+Np
yHyak0RFuOxibsssN9cAJlLjxPCIhzGpvd46x3gPcP1dq3W+gy5h2n7O2RJoDU3t
HO3mJ4yi70ngMxcROe2V2//SYdhYUiwsr6j7/TVwA6l6T7mTijt8qoB2efG11CZT
e7uNkn7LKqHRQ/aL5ODfcPUwh3tEmIyRVRbfNS27KvLQvnXwxXxKSx/vPFMJYSEJ
4H1nJsqpl5ZnCGEWVZZdJPiBKt7TDhlNTH9X0CRyojUnPRup43RlakjNw8AL7pyd
zBXNs+ytGdK0F5GXnkc+TLhtbMxBtvd54O/FRP6ZoLNGVNH2k5B3qdqAVTMG+srH
arHOSqwMZtBOI0OQFy6BtRqhqngO+Rq2RGQovqADY9H95z0/7klP6ermAKc8BG1N
fMtWp0jFq0n34vx9RrFBqWTh4EbRKAZ+kiSJRYYJgkN2Hn8xok0YaQIxVVJkJHWL
G0utoOMKuGEayS0In/qnT6k1KKznGv94Bnm5lzDUTCG1um0jZV06WgPa67Ng6Q4y
JeDot4Mw76DVbmREP7h5+avTdjbBHTkXprOncm9BbpQFfr2JQ76Mx4ggA8Ei5AWz
CZsLq8AXV9VmjGFA3CHIrXChz+7g9bl+Uc4T4CGp80rQgxcjysDTXk+i7aS8/OkQ
6uOfAhzeMg4yU+CaITqaGwdc+aJe2BfoxKCJSTCeQ+9FbT2tdkvm2s5ElBk1ef7x
fmIQ3TxhZ9uyq08HFav0edSCn3kIkgqfTLGITfakrdkUAsdo0f75/jKHBJcSJiaQ
e3qKnFEYVLo5zLKadjaV6TJYhEqH1i1vL18V6akNTO37UbtwiadEdVIXlgU/YXST
0BulfDk8hXaZVqYtq2UfJvcO0Gn78CaASbT7mLSjqWjL0zpbW1a1eukcLk4FtoZ9
83ZBVFHC2OLQ1XenAdhRCUWof7cS7EwTBT92AwAxbO/aaUvJXJ/7uFmExXx7fy27
tl0H+o0/LPLSmn+3HrVsqIhXfRAgSSAEfdvX6avGpbYv7dsshA/QSwBXpLnot7fW
g/AihC02JfRvI5TN8NPOFRCM6ml3bPiXhnr8ylVYAVkaYhn/xKnggINPCImLh2/q
BfYxFONI/QCWk2LmO5Q5uy0XntiRe5ulRNqt4aBwF/yUnY2QLwv8evs8x0ukMpyj
WzzhY82HKNie7TOWtVdu/X4yyD5pbj+ljzIXJmTo17eRuXYQqd0LWQN/LQucfWN2
M/9ofLpA0j0IXCV7BtYXXeIPvnN6hnpbiHF4MVQPZe/iSeFm/XLXR+05HCnZF15i
eteSyryB6tu2w0t11XYaBMT+0/3QRjjpCaKuKvemDoGEPl1hxXDJzRywP6Re/BnO
IL+HPnCIFj31UyyQ5r4wPv/vsLn1vBDpKPqxOGo4CB3RPXfkeSThdOvlVJ9u+/T2
EgzJer/auKPFB2i7WgVYAJC0A/hWzPcZeA7Q8lK7D2bXOKtWDYbzU99JUSs9t61B
X0ToTVLaDySPkM3BkggMOg7kJJ6R+bP+SzvOxYjPB5ivUbmXKnA+jUzaZAFDrG9e
wq4g13tZSYhYIw9cRFWl8uYp0R4IFKueIgswCpN8gMIHXfiLnt9TJr/kHtMH1yw5
8ZsulNALTLrftdGyaJhyXCdjphjlWNPzwwjh5lPZYWIzv3S5oWiFlAVRvjh6GZAU
gKDqYBqPcwwANr1FQ+8TeDOEWXWvi3TAc6GG9/ayr37Pwae3YB8Om5kilxGlGp65
xV9LgJ9q8QKAVBqDvo6Bsg+8OYNC4QzaLs35mXZkMrw0k2YYOviUlM3UNleLCxmv
8WPg3g2PKyLPrdnfuwGiN3h72TPmlzAE3pdOULfx2r1DOP9AYZqVwBSOOBYQYt3W
Y+EVK0vLl8daJHi0bXkIH+5pHZTf8MoOez8dbQ684luvBoxYkSWCKO0HaPxzvTz3
JTeqI2uXJDLOLxtMA+7fHLxiEepkXM4xjyKqkqCAhgYpd2Jbsk2s4ohyDc+sSjuN
az2tvTLmgo/o+hh6zJErLZG9h3MqJGy6xLyNqDhy7Lm3hulLY+FBiX2cCu0/2X9i
xr2KdXs/1dqbEzOZMuqCKB9q/OC0DYoNzlC+adUAU3tkGse0F/En+3eeRQQFNep6
Wwd6fE6RShN48J3tDh++GJ2SZGBz3LhN3axSMjV77gW7HuJPzCYeLC0gTJEG405m
S8EZCl/g/GuuuBiy2K0Foj9JoVO7jvPQEt4E9xWoy/K0ZWUar7Vvpm/7ytCvb059
LfXCQO8dQfjdnbcXY98RYFQ32BVrZdDEvYmxr4RaZGK/QiOFdcHAArJMNMGX1PTE
HlAg3N/V/XCeNYnbO63//4HIa6khM7ikwQaamg5sZTXQQDQl7Z1kqZ+DWhX/L22+
NvKCG86jgZts527RwlImmLi69BhWRbIw8YrfPcr1urAbMDD0LxfKiIw88SkYcGzR
ApSbmMlke0UKjzCay8hgmmB6bg7jM6wYVLQc4VbrNy9CJaX3epgHeU1811wlk0Bs
e2qcjBm56JsyzVkPII1Fxtz1pMhVAjuuCtcoM9548EmzSE20NcYJ/BWYIEP72TBB
vCyQO/+ZC4s7LUCXey9WBHraibb109iYq9cxyUFBh5y1WslHV5A2jWI2QM1ftTo5
85JSZ+Xa7INPsJjVp91sv075oj24cLXrYyrEIuuh5ZAqBvNU2A7dE2JI6AqmLv/P
jYYcgI7EWU+7+LsPpQvtKM38uvdLuTGv5RG/WK2g6JA7v7SkwTMkhY2GT7kcTmeI
eJ1zd0LeN6nui75+jYZXSb4oe9hINS/wbylmxDkiHhANCIKUkQVnjjJAdubO+uxs
1HZStKtjWdDGagoW2LIzhPenda3JlOuAquBQM5x6bQABQlGJN1Aey1z6witQFb4a
lqJFJ4OEepTg00u3eKlu8CIjOgrfGHozWhLdECUWenq3i7DceVNSVPuj2+ABaN4D
wD2pxCebcM04jjMM/oeKUGlkV+G/As6diKNZIHIXRQbqbkUs2U+Uuw9OJtOG2mOz
vlkFoyKJAZ1Muatc9iMcDDGfaDVnaorVFpMDi83mkup6fMvy/nL76zXTKPVtuLE0
9ksj9EqW47PG0Dm9Ck1J1QtR6t+QGxb5g2+MTyQjXyRtsIS0krqXXtVh+nKmFAOX
5zJzm2Vceutp4mcgBGUU8Dzk362huafPJWNKThECv/BdEWVBelDadT03YQh4S8kz
G5gUQZxWLM+A1OW/ibgrY/BlOqP9+E0WBfC5SevlJEyLiGgN7ZD3e90JAiXQwelm
opqqGCKyR/703KsciJA/hW0pXUYuljkYX8j00cIXyoeJClyPN/FF7r7eJ8ptt5CY
pNFYm2vwI6B+ZQpwcGoyGeD4l2w2bOLYXCkTyaj7J6CruZ2iTAdgeXSNrMeg7cIa
C82q2dse9LuRrX+agAyujL/FchzIm336p0bAb0O2otwG2Hp7CqMTZ6BKT5NYOQkZ
0OOGGE4QiK3TfLRT0+IjJDxThLREEQeeGTWyhUik0OCRmcg7UOuTVwoY5plhcom+
rFu0TxJfJ/ArLoLhsEQt+qSK4h9ssMtTveUDXh/0uidAHSBFeRL3rc7ULOuGaZ5O
rOna0djow40+fKHhHhW0ZtcnCEBVPafmISeG8Jm7TxbHy86SMv/eS0GQdED+NhAn
KXQhNa73lChPBAkrsryKYcSHQpZXvYkW2INhqJXk41n0id3N/CLqE2fWKR1FVubT
AnMD5kvW2GcjyHp1NeSAp2zkBjctydJfc+EqwQGQhaevSZUKQUkt/Hcg4kBZaFDo
PpQV69dSTuU/5Fk441I8IePOd9vOYfSXg5INMyIrgZQa2aQQaU3OHsA5evM1iY0z
12gMK4YPIdYhHxbmsgFBav2OExETKsPeK3/al/RWM9k71f1/gSwppxP4J/K5b+/A
eeGruaMqoReejFgcemtHn7O2p349vfwYEFaOPduEKI8oCHYJ4E3kgdPDdkoI29Nv
JhKilWkdbbBuHXXmdhfsx8PU0xKBsXjDbzpRHdogwQEmTtSnhRzTLt3WuR65cTrY
01CPGD813ydXjzRIfiAU2VgWTKnKcsMbjEafSfgqyvzjNPHpuBTsxXf3poeWh9MH
9WdoGeIvCq2X+LN93/wWdQlMVPLRa2C7LHKcalfJx0vBa8G85DttyWwoeMHi8jlz
x8CWQ3LIu1Pl8PdIJYiOamEfv2/ppzvasEw8ARIT27KDjCj++b52Y/0gvt4/x/S+
zKPkz/O0Xs5qrGhU+fVNBPY3xVdzqTDZ2l8qzy1XYuHyIGkOANTMAgiep6+P+0mO
uEGV5XanYHZJv0E3G6LhrN315yOOeYvr8hZBgJftfL9ZGuQiLGUyzZOlQUls9QVV
PvaT2WkBGimvwuZdOlFZ4EVJYuC1vCfMOwzGqwZ3V4VBVQ5zu1dEY3mZYsXVEcjU
7WA6FzvQiU69aTDOhtfkyzvPObccpWJCKqP0+iljW5MzPDEJi9n4I8vKbOc6/XX2
pJFltuSvP6/4bzIzHRvOAqwxIMmnET386bS31fgv7uvKpYDyAiFL0PZkegTNXiRY
V9NNInbeVNUpoba+DvDYIMiiXFGof6zx+RLMuzXbpCynTPAuDl6ebXrxEjFx2KLM
xMryVG2MOq0fi62ygPplmxqOwi0xF1Ik9gilKbpZAGf62JXoyCJI6a7MzsqJuk12
dLmC/OBsbwzfybjp3WCSjBae4TTbRc4f3ZIgtXo1UanJvOaFhN5WST8VAzoMoEG5
aIjKZ2G0PFcZ3CGQNC01PdaZA+K1L093fWip1AR2oJfHfwoKfEEWMqUeWrAbXMmU
tfJral3/Og3cpRBY9wTak1zgw6QQvTckytTZw4758PG1bCk98jWcuWZ6xgoHT0dy
5sYqB3ShTwbTFUOtQhZzILAvHKFujnQyWwLU/w2axoTaG3g3qKAqhsLvXV6Uf/mF
drFgHtJVEGJS03zvZbJLMBz3kZEUVwbDcDHt8FB1JEpPNZB4FbZg0RtXAn1PBIao
XCS52CwVP8i14GSPKZ24rca1QGdLBzjy+kfQD3i/HntsHG6sbEMWkSLF5ZqEnJRh
8y8eF8W4IbFggWQOAVGm6a8uF7YC3FWGnr0RBROYiEX4jP3isCUhk/h0y+4ojEVG
88BTdWKBC++9qWu8e47AwSQMj/yIJvjG/jzEnZofkmkRjFYTNGg93NH+bCKFS6wn
1tWssMS/xfCvjZd6PaeiY/delUCI88TGqt/JsTPFPMEp5xU76HlFfmVe847f8Szd
h9wyGV5NQWnW1abBCnpfU6hX7Xs4FRDlMB7x8yy4a2yyxFcLFRc29GtW1j0UhWo2
h/kmp9RTfAF2QuZCxiz4xyj9fkTNg+OGdGnC5Nh9n9SDtpPuYy+8atMX70Mh+Wz5
JW9C9nbnKifAZaFYZRZvGT38hThsP8wbSnLpkIG8Tyfc/NqpFalUrvFKFDN6QLu7
VnlZCrAXynQj98wA1WG/HIKwBud8Z0RnEoDXV3cOzZorK0THMJcvDZEVGz4VyqV9
OrQ17/UTLGWPVhcBXh8ez4wyrqiQRApGvxcyjrwPuvYvnCEQNDBeTdbgV3O6qzXI
MdC3BOhB/YCOGz82ZPm5VmgBOPel6iY0T643pOGPoZVjjQXZG4AAsinWrQmM3mBB
CC4gqVaghzPlcwLCQ2qa9w4ZJwVMsJpQLAwEOvm7XgbiOWsRaoeufwnjOhxobBxY
hhtXm6SS9w1BpJZ5gjSgBDroZQEhCKTqXzFiz3ZifYFm+fbVt3WDRdkQyOmI9qqz
pQdtFB3EowHVKKc5yfd5DdwyaTFg2OGvSmLM0SjN/yX9H/d9zmt5j0OUUIKyqVUb
ycER/JEo+gH9bBfctnYGdS6wgqqIVAalGUhKMOyAJdVKUgY9RsdsSrBxdOd8G/yg
SCK7Ju1zBqROeFEhPCVHiMqFtJs9Zv8MWd0lPbNCFJcA3/Yw7C+AQBuLj0HY6fot
UpGc2wPyFwbyP+Ec5y8L+B8Tb9+AuQ9fx0eYnSo4EplKFyI6hNgZQX9G1bifAvXO
D3QpUkbKRIsCmf7VEiqGtb15RWRA/yb0kq3ndVsAbAhWvaAtzy+IiDIzNAMRHz5r
JYZIS7JP85wihh8XoniJ8bR4dhvBlG3WTIrHdANLXQKPyfjAsfLLbXXjIfghfjMt
nV7pOQ8mUYGhTIOQhWhg4efsk24tJ7XJrmFy3PZEpvYCKUyfTfDMV8GxtkcS2h05
oBsK2ACJ2uGJ4IruD5X+lye2ZQIyScYx3Tj2Mcdw4Vm2FqKzFkehjLxbqsGj9jL0
t0yecb+AiyOv0EEnhKtdVULRKM1mdQz5PYOo0yW8w3khRCd1QcHISIaLaKJkI42J
BG98cWpjzTtk/CAI8aVMNdkep8s0OS3FP47dikg9sjfhpDRpCff6wo2mr/k/88xC
Ruk50QJ78buFWOrWFidEfEPOuI/PzraUHKo/ExzrcHhTdzdQ8dbfpFQ9GKDZ6WEO
wkcuNc91ELyLQoXXnsQvt/3Ya/ahB5dvYIMX3ur2X4LL66HDsnU9MYIaIs/Bnqbv
sNWILmhdx1d85Sv3vpbthrYRKLi5E6Ul+m8WVnfthLHylSMKcdEbRIJT/IhSJ/pf
oyPcLRA2ksoXsTwsrMgkyJTIj7ePnz8xoAPdhDPLntOrow7rx/txM/MS8nLrvKsA
1w06Xuy9yFVakacwImmblPZ4ObWcuJXzR21+i858g7+Q/cN+xgc5DxLVZBY66Fla
biTU6mdCLEQSsmPJScdhgLh4qdxmSg7mdxYXBDJCdLRuzxat3gnp1dcIuGBhDIku
WaDnniE5p1C0FEQ5e6EYQcB9nL9lVmp2Lwg12QVo2KQx+S4bT/AcgJ5Q/3DifSup
j/MSpvxi0dgHiqizFmzOsq8/PYZUjw94eJnUgyyz2+jxXLWnUuBx4UFuyUIMX3bS
OChkpKf/eZ3JpeEqbJpgFMCWa1mUwGy6xh91vlkof/Moln/FxALolJJFKb4aCyzT
eysggBo8S81zMjqnL4isKLlVnw/UirriVUGhj/bpfTZOfjUbhc5VF7NXs7tMtQRe
2AekmVzxlQAedPEKSAyJYPvme52mmuRBpuzKxsrc5b+SrafncWsXwnurV8sT2Qv5
aeQFZNvAP24vr0h/bKCT6lygcNpeIkQexi4NIlz1qEpcivM2kx9I0uelLGhZdByo
1LTCt71ic2KVk7gicwJKDI5ktk5GDB3HhwWrGPPZTkLpbREkBILFdMLGjD41DeV/
ZO1dhP6xpu0PSxJ58LknlROdEwABjUfPr6WnZcypmNEexZlVinNmIbT46sF0TyFV
ZQ6NT6GvigHhGeM0ph9GIKplXv9zcM1UtLucJE+OOBcMjHyGw8eNjnoooOlsxMEx
icRuJNJ4RW3ITurJ8KIdWPzEnISh+kbSS3LbWkNVEulrbLYhXlAI9ZE6cf9aXKFD
YgKDxsbgzw55JPz7199NoUSCX++kydqNQdoxmvPejL/J44saosbHT4CPMMyIsU5N
leP2P3sL0GafQSGIphSpQfV5YOufPBMw2TYFqkR+EMBo+PbuoEFPrnBkzkf8FDXq
Av144kir/5DRLDPs8dPnXN6r5NGgHwDcF/eeV5hqR9qz/UtBbo71RJjYPXy6q7kH
rJqinlRG/F+cJH7ONsqGGcXcTAox0nXj62uOY45bIxkxk3WyLDJwwoTHBxmrSKqC
QFEADOrLaiMQaXWDZzzDJePRomc4MiR0q7WoDlzMFFLKlK/GXP7efIIDwF1/kpyf
hgwnNwIYcr6HJMueNacSuaEj117RN3kCJflX0T89eKHHP6U9HU9IDtRISVQVcw8z
JBLZW682haWDI250fl9P13opcF+rOFSYyznCbqjTr2DDlmoVvJ/34hvd3MBsimrc
JnmWJTgpQ5/ImU8gUyV8fsXZfL8tg5GF51gFMKZYwpMHwgNSIiUmuUAaJUmfUwwr
8X4qXm4aSbJG0/Ox7kB7iIN455bhMxWfm4QoLW5n1Cx8DYxCkMVrCQqPKTKqY2iq
2iV4rInl/kfo70leTFnndU2ZBvw5z6+3ivwZxgzVeQobkZs4hw4uLBUVGMcW0H8F
U13BHHeUn6sPfrM37uWMiXT57QJKfyzzV2FvxaLzuWCtXZhKuzkbWZsSvmOb8UUh
9owLCyqSOVynJ29EivBhJkr2+dzVlRdkYIXkKxGOWOCXJkGXBAvarJmzPYI0EU4/
RgneWyufEbzWzYctBRNNtRbWMwXkXg8fDbBI7HSn6fg8gauoIYSX/axFUASZV6w2
bJVbeH5O4ij4ijz9rRklT2guX/PpALo9zbTowG1ebIJgS/PlR1VFdOgLzfHJxELd
Lxp3wqYeigtNAcriqc43Rl14w9NTgsiGVPfcGjBe0CMP/+fFDCQoxv68Gsm/FJLq
GW8XWkTsoz0B4Zt92f+dFt2EO2BDbUEfoRhwuwy4JJkOtJ/tZrmmx+EiZ7Yo0WAY
X2R1muYYzN/+Dh/dt0YnL50ZjlkgQH18Ye3seuJSb2Dr2i2qSZJJyseEbmrt5+gp
/9Ps0pATHWpGnzTIPpfikzJuzlHp+hShxq9Pl6GRpvoJ0Oihg9yyIbbVYAZCB2tg
gpmPGSUaMlZzFEl5ZG/sNR5vvnOT/ejCgh4ixqD/44NRq6HUfyuCFfkx5qFk5owt
fR0uL9b/HQgI6xJNoOM82FlcwQrj5nP/57wofisHy9eP5G+LjLTTClUEUcSucFV7
Eg0FAhu29kmTL86FcMGCZyShBEHgr/V9FTTgxCvlU+84aNXENToqY6XW0s+/ZTCB
LxxFZb3B15kC0A1eofp4W6FW5VB9Sg1jswHhZrq7HTBeoB/GEPJGs8VRcOfqEm3n
7UMpouf41vo/P7fSPbylcWbI49kY3qBctDhgHfmplHoRmm1u7KK7IFpdeIsqoTtX
1q30RsIwGQBHBPfUAkryCQm3WD7Zmj0j4pJRrKVFa/5hLftQp8YTYUyyc48VdG35
eG/5L1FWldNwlxufwgLhkzq+ddvH2Z+0HYTHcB+f7PW62U6zY2BC4Yy9CWY48HCB
xaWhKNFBO5TFeT0ShZuxVm5uQ2pOLqJJN6RjofYXpGNIk2V6SuYFgbDhUlW+JalZ
cjmTvtc0ocIhrbeU5wIP+DJBkH+DYQTC+BlJa2FuewUWebeK0wQCx0IurEqM5Vue
p1SrPgpNk8F1sWCWTm2QU+NTy2Jl88c9qSA8QN5jzrZGpmGAe3SYwc+xQtBsRAfU
XFlPEoaGfn7O0lUjzTKkBD34w5bESrVO63Ha1fLdHFVIhj6s6dzUaHMgJIWMAlwr
BiJUvtwDYEUmA4vuBQp0/oev39XglNSmZgm5ObpVxXqB6yKu3RZvCwiIr83gUhiB
gFsVYa89WbofRPcRU5JM/GncGn+5PQD2RinmJi0IwWk5BgOKVT2dSGzDPqwwlZTo
ZiLd1k9Ydq5WQ0YcLVfli6SHf+B2kEmXWYIQ0pJIklDAOTG72LRRNJB8GbXG+dt1
fa9UP/wGoIF5waNfqAwcDK3ElxeTE0kqXZxE5WgvE0YEloaq1jBSFFtW5/aP9nGQ
Ppp+P65yiRJk7nJdRdy5cENWWkVSYageoCTpsu42QH70dxRiarjX6y2DGhU1ohpF
MFCryRNKWfcIKwSM40umcRF5n5CKjaFHLhYuQwii/KOhnnWaS2PfPmkIpUu+RVox
NSbLSbumngG+22Br7xvvZSXSv+vBSTb3Di6Yil5LkFV+wNpDQL7hKa6jWPe1EexL
yIE7NUIrfof6qhfgYk9hhIxcAQi/Nki5QM43Fk0tEx0BE8Z4lED5QVkZCPjBFF6E
3TiuYR3W1yfxIGt1NHUNwRmuuwG1Fnm2rf2rhRgMXj6/b0VO5eGf0hCENCzVKMrq
je9MXpBjnfcaAt36mMmIT9tjd4U8DrJN7Dwzq9jeYLIt/lxpy6AmmZ89LwsTStrf
qb//giXu71lJgnzS6ZynxrUgmbyrz2W03vnIiIB/Vqfg41vJV+Ir2h7cOkz7oOID
z/oU57syVGJlCEwBdx9TL475Qtp5UU0jiZQ6VsbUxZ08nxtKeS3wdVm7RYpkkuQm
VDeZKDQPLKEqlg4CwFF0LXMQ5NV6u8XewXdBlRB2NnsniXPJ88IPKZBISnb78Kou
1dKNGgtX7xEz4EPOAyw7WxevEAEaKYJRqJDqITLA0yAEHlr1daKbQDmLpjXyb9Jl
q/kHZBkzANp1v2muFiss1qmhyN7/rmVLVb0jR1eL7Mi4gc+g0OtDkwxUJFz+NqMI
OHAQqaZpnmoieKeoNrXJ154TdqYTyfWk/9AVy1zrKNgb0dVFmI+UAmmcIXuJnL+/
7AFLUn8LdBC+kbOu5k/V3BVHMNu1Sp/V3h95OnRvE8UE8dRd262iZ7F4ZSwyL6cA
xv19e8QbUtkTAgJBiJEEAyF9S5pa59O3oDdV9jtZG8ZZrryRC4hH9p/DPgytuWoV
ldSx15FyBF2qshzSstBAxISOAU69EaQBs5ATNl9dgicO7WxEBqKpotgE4rKcFQX4
GAd5JUaWX8rIj3m+SoBq2tYohcAz7NKFjiiX/rcgTSlClt6761vbhDgt9BN8+2+z
oyz7gBQVeS9C/aOehaOm4Q+9q9NdzMpSeUJbLKDwpTZ2X8O6y5vf8qzHLQGvYxms
AbQf9cE6cb0qXtIr0LLZEkIEkeFsCjcSabWdhRikMK9ds4YvOBNOaR6X/N35lti2
EiP2lX5YIIHFpap44O2pcJYbMupiWmc6L02ROMg0M4YCLsc0ehIdQ689HeW+5CK4
7eSB2o+xMOXAnH7roaXPqLVHJJxqZuZXLUknPczmULzjhucWmTlonfMBv/NlEein
Oo8O3jl7J6Ks80XfIvoCIK02WtXMWFYJ76nyQG/7v85w6HjU+FpK+lRsogRfm/Rj
sjH3rKDFjzGWGDNM5JkJ6Hkybxygwa2jcrSq6bIV+ZWAmTvBR3RpmdHQzLxvrSC6
V6ekqGyI+s4lObY6wImS07HATa2siCEp4H/zz2zSUN42yS2kQhMmcoKNL1ByIYKb
FjsNFSTlS+dK8j6yL3jrxtAZS+n/UtImcSPNKWreJLvnTviLEb79ktvfoDiixNY+
Pa8knH+nNxXGkLrDnRLLehvGlgoSIE+jDYu/wH3mQ0kruyyCqesxxfitmTftfBxY
SLvBuIzaC5t8X5PwlArLoWfzk9xDZZTSrsqEzy24Ngon1ty+OWmumWLIegzpT9yD
HgDp/7tpO/bMuSdR15GZ6D/Abgdt/C4OXMdb0UVih9vHt7YIIlBtJKPj3Hiw4937
R4uG8AdCpgSiT65KIHHGr+oLiUYOSmt/0hPpxpytP15F3Gz2I8eGqXbCFYXnL9J0
OT6Po9A0BZt8nLfsck9YF2bg2WjpcG42eHpc/OyOGvOZDBXvkfWrE56qvMOZyt5K
tcEIrATcPbG7h1A4wlLYFp2g12HJFr+4+I4+vxyXYnRe+XbXQc4Sv9mvUhYNMwey
S70bv8kaaqJrDj5xcD/AswkaxTZwM84/S0qv6kbxG4CzqM2UoRPxOCeHJ2QGkjb8
AsbMJYoJwoCmKctoLHBuVmaLPyrZP37tFbEBlAeLHMJs5V/H4MLxh4Kzgz/jET2s
lnc7L69S8JipT2lQrRpPsw0aVWcoYmiYciUXbCgyr1byB+8MqRnKC7mIs4JW2R/m
ygXeKKtAjy2HXeWO2CB0g0c2BDL3V6NxpY7RMq7fFPDzVlJlC2qI6kMUL2sTbuQY
7QrabFxykK/KvYv9G5ynNTExTUdM7JbvnNRYTnrLPBA0kyTLUHnKTrNuBzrSPEtA
XMcVImKnO5xcIGNwjMITog45R0U7ehd16OARsZDM7G7dg99cy0YKk01H4JUu09lk
bCFgQJoHlb02kV7x315BWRMHB548hA0QXGAY8Zl2PaK8U0pgWEqMnzO38+GJrMbo
zOt2KhWdigzW4dTXVBTY7f1fDbFHLbyOii1YBaFwww5MRA/cjPmOOInUiV6EzgaD
PJ5Mq0rWhn9fP63pOkF9U/LCTURE2Ey7uWzBRbr4/capqPY9JODVebDOlD7SG2Fm
59deZATHzpgxEFEIVx5l3DB+Zord4yl5TnmKNzzd5vn4/Mus/NKH70bJZc0o8nMk
Sghg5ap0j5xgosecs7qQfAPzvWoMgLLi+ZLwvP53NHuwG8w9muxX//CQzxWptqcp
mG70wjcx8GLMgS5a1g48iqyXk4Kr4+ZEmU+fhHYIVwV3eUu7iugOozWZNfi0apWX
cWh+22or+m/8jRJYjS5mVEwk2ikSqwI+URjU0Zv9daQD8PlqESBhD8q2ZdbRv0RT
VqLbCqS0Gea5ETX2QeNfHQQNq2pYMYGTe9PFdqV2a/R44mclY4tX3FkGH83S1gVG
pzXv+VYo0M2A3x6WxzX8Fn6pLkl+c9samshGTp2GdjYH+WJhUkKer03a/w9HEz3b
yQDBnKWv6q3wrEXjeBrLDoMB8wBKYn60zJxAOQgh9URi0iAZbNQEMQWkPZVvrHgf
6B8rtr8hy5vpi73C+/IF5z94rCFfR6VIr1YTMTdrrimPKI/NdQ8xhK87yP1d/zCY
gH9k8/uLGHwqmkypW+54T3R0y8w2JB4l2jKCFGA58LD5+voS2gHX/o4PiesVo/e9
2N9qAPaGvCB89N/4ByNzuf9+pMELl+x2uqgUg6AfKstOKffql8aO4k9jke3Tx3pJ
s5dDO1muX0QECtIAnxwcfls8l94n2xecqBiIP8V/Tm6hbpsWEQCJGL3BJoKgM0xB
+Wvf9Rb1URhhs9aM+eh0QIqsYS9mqnuBD09UWeMlKG07isuQTpX3+H5b4r7jEjbM
yldLXQdQwyt/sCTEtEwlTFXbYNVkc8/tKvWrg1NhIl7k1Bu8ETXCy98VYJkzb1Cr
RSe61c6PxQuwljL8/VUn6GscT1kdgL3D0nd6rhEWFuvY+aT49V+FiUkgryxIU/lJ
eh6vrxVIpYWxt/Aq0fd77bSK/Q7uccMEDSttzAfy9sHhO7eNpQLK09h0H9r9JW6k
e8Z67xPMCKX3QOJeTuGJlCDpwrUMwivzkWIzhLuPgbNJdgw0+L8nHWLVOU12qYLg
trxa9gnetWsS8FLBOrrA+ZQJfy/vP1q2GmN2IiGtkZapaju4yYm7KI0hlTmQfWSK
Zb5xnxrx1Ka1vY37V/UYu4XJk1n/0uNSMijbPB+I1zSi+dIOtv8LM5o3R0GqIn0i
9FPeLH5gJSoB7pqlJC9UncWt7dLRmCDyviZ7yNr5MFtJokNxKcGl3MawhBonDAZi
0bV4GQUlkxw8u7DtMSNVqyRkxk4igC0SXbOsrmp64VfKMV0Z6PTQ3Mi1abciPWLk
wSq5muMETBh/Zjf4L9heoZbAqu2AmtHAmPBb7/g0aUFpMMLuNLg9LKg6B3NwczjL
kDZc7ArxvMH41OC8eGBkBxEWRS2+pJg7xWsBYuCo3PfU8VpVD4Vxt9nDwRWtJWxr
ebr0PB/g7U8fUcgTpifhUvbF3Pdfolw7m5CcdtQFE82xHFG73rXeUVR/0J3w8vqF
AMDyT2/7vRW9CMMtwtbVLxv9ZzCg8a5IZ347YpqvYldk6p4qVA3Yg5YVinnGYFfM
tucajarsFGNqt2w4rSYLzNI+pWxufnY6jdLelzKrr1tzrTe+wzw17rTsVjjzo5Oh
0n/1IbW4zxyFRRbkdH0KI3/bhtb/qUQpapQRVppSgadVz3AXAQp8/NN9EtAhAlJZ
me5kYrCD5T6o8luiyaBhamkssOYSR7OfMhAHUyUTxMg9UWFEavrz7y0aoeU18sWT
zSqTMh+21Zwli+OhdAs9IBMgJt90arlAVby8bOLUpEzEV4MDDyQ4GU9pqQOw1DSM
ZheXEmERJKSpPnA3ivuR0d6p4rOL07bLFSAnnLtaXGuP9qj3FCfrV7tA3y/bSmQt
zkoM/l+PUysq8iyKfTHxcctdTZMSwVwV82xqvfNZGbp5CmjKcRJQkPrFECcErlxg
kvHg96vhY1YiK6fRSQDY+kiWGyEmZyrumLI7VzFq+dT6f299Ddbqp33xMfzRYn4m
x3xwo9Lm1pupWCntpAGQTEJjvbkhYxqei//izTsRq0WzukBhqePiCorMT2DMe+l+
SB44krR2KVX9o9Ni3829BtpZ4gKqDlbWZ9mmOJy8H2+UAlxGvz15cSxxH2E1iZI9
8UM29W5aBzCKuFjXRQqYUsXw+rua/Jsuf2jtiorQhsjHJVdRDk14/QFg6Z7VMkh+
nQqHOb7ey2FW3mJndcvwiqXJXZo7Nxfj68qYz0KMzRRlGjCx8Z8Xz3dqcnYUAZug
gTMTsJQVqOdQuL5njWGZm8VXxpOejangqpvSTymSDvXpX10kmJM8ZWXs4+k0qveK
W/ZZASe1xABsan9oueAqPk66NfBroZ5zCvgtUnM6hLnBZo7Kvbk4spVnb5BQtHzW
QqMFD+LIKffJwsdwM3sdv6EUYMeD2bjqcRII47Sq8VucBY2ByGrStrHkxifN0IT0
swC9nvezEJfGuEP42a12v3TLNDPYV5TyyQQjNfbOr9okLIWWJrlwmAFB8E20IK/k
fNvyoo5FUD2ldXab0m8So4WHu1e3moBz1QAxqA/kzecnDh/ufjBU+R/kEA5hPT3O
e2e/rkj2tafsRX9rm2gq4xR6RKBHPKyOKOzTxWEpLtkbnQXV6q5D14XUm1EOC0Le
xdFQhyayWvuBHl8Gz7AGYROuX0bZW5pROQEho2CQFfl1bQinJtlA9cGKQHs3QJj7
hlZsM837OEbCm2+5Actbi1Jx7QhHkkou5IQEtyaf3WQidUyCvezDa5YeIUx2CVQD
CSZKfJC0Cez7gRWEa1MDXrBNPrEUOnfYITdVFh8u6dPfAsifCdqEE2tjXwmo+zLp
gNhCpy7XTwMfopWx3jsDGaxrFlT+LFfS7wRQ1JEr+UxYrNUd6RwneHOEiehIuJYf
im7+fF1HQ2qXAGOAGH97x1aaEdDYNS2Y/Aqml2wJvu1NCwG4D5BM1i+JcN81ZhTj
og28n20jnNBJkLggcxumkR3RbIOtJLVdT3Ym0Xqs5rey2wZsWKTw67EGmlMkM2v0
wN5YGvIaDjiWeXSDNIm7X/7AJ+TPZLllrVQjaj/NfDuS/7bKFvlmfD+WHjRHp2vk
vATVKw8uvYX5s8JwKoSZNJLmqkEiCGIEcp5Vf1c63mH1rhQ3Pee9/GOCWtNnbLJ8
jFBrQXRSYXkkvcVWUvSbpKgpyF+biDkZuAnY0xPJSbkHrSKd8NVYqriJOcyk8LIl
asVulFLjc1cf5+b6yaUcknmv+o1txUcgJFBYpODpJxF0LbA3VQwr1R6XMaBrGvMZ
/t3oAnKivk6RVZhXoBOoPUoms9OR4qK1Shdc7cTmWItQC01T9xGqNGK2jcF48PBh
xh6xIvWdFoc9i6moERH2ezPqnuCDstB1EIUcli+TEFYg+KzlFSeAko6VEQkQZTFR
Z/tqpC7+EZKk3SALLm4ZiHXp8c45MP6e3bJXeYX9tMZJF4EZRD2tm6UNHOnGPmWi
NlyE1P+uDJtrXuR70ggbVXHCKO5Qar/Cv388FXCO6O9VJ1atQr+E5xEhSPJ2qAqa
UwS9WYtWTtoj1/SFdm9rPuv8AG1DtOaNl9IZjNGbNq+DQlONOfn8TKTtcAszAsLn
o11boEYvKMSg4ooIBw8wVPh5Nc7rG+OIufHn80wDne7Fczi93ylP8rJuyjwyYMD1
HXf0YiQxKiI0lKfKjEmp+Tr3GARlElyPv3JanNT/FzBfa0w/9EXgFX+Zn2PS2KcK
fSNO2DnDFi4Wtktp/w7FntesKGk8LrF/0lQOtwfDuFM4YcSD6iZJ7AbMrm9FSNyU
k07X1dXZOEyKfZHDwXTkHYK1Cb0Ogk3pIWGqNEbdwUTdQ8BxeI69Ua5GcG6cLw01
+rdNoosvPr5rmFq5khSddYtoA4pukdFQJcgE7zQhfcRYZIJqFiQUbWDWaPp/ntW3
ufDtDcURXZcEhTalULO2yQj9oEvc39SDwF450sq2TY8W2/NNUhWmPQKoKusrArMW
LhLaoClsTGDjrq53XEHd6SXNce+njrMgz3UNv9RDGAobMFxMHJnG41ytQjs5R62A
rNVT2ddpiX6VKlxd1ceqOyUUIhZRVS5OpyKZTxrPHAd/T9FTEhlqFi2q+hNsA3bO
zDBeiPnz51e2OO9BfrA4RzrcXkW743aPRTk26O1VrUwQNtuOwhHSq2UNBwi4wXvk
3bbYr2VXZZdGrGZVJneT83arrgmWW7VD3wcnnTe3LUnVU5PIr5rzBLoMR8B2LXbV
+3y1FCDEQqMjtSSJVGEQCTqxDIwm+nPqZOGkgSWdSCFJ4IdHNEMc4i1qvpjS5Gj1
Tfa/ka5nXbpanW/OnLUaDZoRf0Y3+u12Vq0HkpJ2akaSoGk4ZVHyzcl0jbH2yYYM
25JbeNIb1dc+ZWRQs0jJggPxDvqsADK5tQbu3rT6bo0j8zdtlWV4y3N+LP3wttr3
JpVU9u7ar8j5l34xDU3CCdw58SnTlYjKlxRvNkiztIVBgWLLssgieCTJRdx3k74T
C66cmsdbD7m67rGRj9RxyKMI2S+dB0CPA6YWa/dHwsFD/TZ62YPH0t7h0FwYOdtN
qRWMk44uty5eMQzMkFMVUgBPI4EqwZyLX0cQr7CY4nJBaGHVwm1yV2jRgAGxVwDf
8o8Fyqdblc0IHZ2wJ5/+vveosyMoZrIGXMHY3ZKTURQl7Onpnlwh6wVxKu+4NiHx
WKNtyhSg+LdCL70u2isU4dxr+20O6mGKwmi7XGekfr6EVrp5ySheZlgNffgrR6z8
PluK07CzcVgxt1IsMxAI7T82R4aEQtSK41h8/QMVzrPsGuyt/9eIBhh8J65XVb00
Ao+CagBQXUsKIEf1iJJG617oeF9Z9l9JDAu0hJxCUJmeBv+GinWKS7vnCzhc/DNU
TU3VN5tNdyqjOqUz0jp9qUokVKfO1rvFRyP8daMN8FWdzm5kZuqHg+EdBKXs/ig1
uMyUEnenkZhPS87vdINbHyqDfkhkQRviPKo0DBx7wvqHhACAeaX25DSp0bu+YLLb
B5rz+5GI+NGv9A82rPde5P2g+IhPqRi+V5cfSGcVarry7D4KW6+XWY6WRajNh4cN
p9rZp3r+jx7bk3t3qgP1ekOfZtikqer7iYsu5Ks9DluDI0cr7ILkALIpESyfXmG6
XL2tWNcr1Qp7IITdJ+5qKpjfgwVorPQSImqsCTGNcK1dgQu1/Q+3semZtpMcR3kj
yaZ4fE2WUWIitdX/ie1kGKiPEiTIYjjZo5qj/PKRTHXaHNhSCBBuuuQ59PnZ1UAS
aXY82Mk5tXq0OM2p9q7GQliTBgfJ08tr6KOODRpT7+IGIEJ8QAuDtnd+jECq2GRR
V/TjLgZcr2cHQPzMydRehdY76p375tTA8fX3eEYBtm+9Ujl+AFzBrd14NvZCMsCw
70PeCBnzfKmZVMG/JyJF96wq/TLdtgPx0C6yEOqI1O+Zl8zvpX9gok0/1Ee7AFXJ
++xndVIPC+pYdghHYODIfRpaUfhVmcyXyGxs6ERw3NI3jxWI6MhL+PZm1/mhYL/z
ET4yr6UfIDdXg7xPdWu34BeSCzy+sGc0cbvlsx8hGwiSgz9TvMyr7HB5N/81lB6O
dr33/YE5kpD1qxSR/WrUSkVzuPtVB3t6CmWjCbaSI7I7PFfcjHWPYVDjenp+5w6Y
B0k7CICLIui0sP6/yeIsTtEHmZwEaIjeQXsrsNPZUgetIR3+9jCyYYFVqIj7RLzP
4oQX12GSoRCjbXrYo3BYBzIOSAdng6aNZqV+/eIPt0mofmmQsP4KWpeNxhQs5pNZ
Sx59LFUgA8fbPUg6AdvCseQiEsHBRDLF7xGfC93vW/6SaSOi+c+SG5qHwXfKwKg4
HXLsrIqxKMcbqcspHLTNSU3YKrHBPBKjIh+NQZThh5WJApOXRdNVgRQmjrYjPHcY
p6vxvhlUduxng1BIsIwe9EJiE1UE0B53LGe+DXjM0ua7o9DbYFjIpcSWdmasbhzJ
NuJaF6g3uIJg+n08SRvoF74gS7iwtlDFgz2Mhf+y55ITJ17HnqXkBoDLpdBTMayp
OhIlk0pOkGnVD5XrcI/YDYEbaEfj6m2Op0F/M/x6aTcGKJFDu9LWnOqueSwFf9r2
Sxk2qtHURSpjElIZ6zxVshuPGiIEW20ajGgU+VSk9Dn9r70etbCBERMOoQH7cZy8
F6R8gA+aWev0PFk9Yu/59xHLCw1GkkAcgniaXNJONeeOWyGAaLWIbZezbJhxZKmR
k1vJMSpmCCACemKW/PeuGtSv961KmWYjBcAxWBT+oIcrGazabW4C/gLkW+7bX4dY
3HvueR6ud97yh2CIadcnQguLH3F48UhVpAUks4pnBA0Sr6hqkwkCGasDj8JzaPJl
rQilIS1m8YgA/9QIRUcrJwS0Awj9zjARd+rxN0VJqxFk+lc9fmZnY34SnfaIf3Ri
LDCuOCCkwk10wtcL3axqSQHZkh7qlugSO56KQjioed4lQ7n0eYnsALRlsOhaiU0x
Y1X7OF+gxXIvUdlMROaKBIxVrlv5AhkYWhGLouu/BcKPQ2iNd9c5G9qtOzMdMl5f
1lf7//gCzPKPtOJoe4kKeR0PlW2xzYw/JP4PKzS64BtuwsFadLrh6Z9ZDPi1wfKQ
gkgekkzriAtNP2M/SxUs9f4QVYziLqvjMo2QvRqK5qwEz3WI3JWIyHnlY+IfNcSE
chj8gspK2TMrI38c5zrBe2C2iP9pBKkrSo5ATJ4kswxvInN5DXxnsnDlgMkF9m0t
bAmyzND9BDDIxSozJfdoDaH2RTQ/jOi5XEMCjFGDJWOh1z6lLyueO318mn/onzGO
hLdESynd9gO3ICfGPGui4tGAtHGivCIzFmEZNJE2CV1f2EWZYRjntnpDYlK3w0Ml
ZkDJVAtRxqpv8ktjL204F/y4pp4RrSMZ4vv8qpy5Pig4f8lvzwuEAsIhhGLjISSj
5X9j3iU1KzVvyzKHlTQmemPuWwnqE3pxroq/t4we2ofAEM3LbyOexJn4pdHg7Cay
MECrZzzYmljyDxDc0KdN7WLmxcRq7jPHh3uZEydRw68j85ek/+LYZ66q/o827YJs
n6AIU4aKpmilvK80KcsfY/Ub1sWa5RdDCiWMdjHfSSHv1rN/f78DImScSCgESAwS
2aoQBb3IdW/apEYKetu5oXN4z96iw2x4KC4T31ELHHiyN4TASLkYbWfM0Mj2DWlk
cBK6gEgRX8VJ2rNfpezra9XhpNwdAnh4ymr/9M8A9pXkRyU44d5y8btWsGQ0iOSy
fH+2Jh6Eossj2m2xagQJvI1+Qz/FruLh4Hm+FC9fMRhu+i82MEjJs0elI9tAVVqr
CvBegAnYXu80xpKZgFpGCDnshzjlVvoQSntDvm2cZD+/4Qv5c3iRhxI7nMqDI4NH
LvoDITDpaYU7+17D0xflunXPZos68cLRbFcM0oosh/OmY0yr5Nj5ukwAt7LH5n35
Ocm7yPiM0jOnhuNcgaV3nqcAvhXcdykPMkXfuQRIO2mzrrpEBdsDhPxhYFZf9C2T
ALrrPiL0jPb5YAa7dP4G3V4gC89IDHhFJACBXgMVWcPCBhOxEQyYh2YIrsq6KMME
G+bmUmUywZduPKVvemc+VlgXC9SL2V0B192tZn9Yjl5vUPOo522qk2SuMtgJM/k9
Ol5NCFG/oVXmtF9rM7FNSfkgpzl4Won0skFSo1aBCZ0m0Z/LCY4qCjwq9z4EwoCd
2Wdr5CTxjbWuaxj/3VCZQN/WDlA0SfA8RRE1+V0ePPHVH0sO68673g0EYy8zJ13r
O+aVsifDgzkQ9dSHGxvg7pC8aDL+VcvG5hGaiWgv5aAQrs2TYNzuOYxP9Y60DKmZ
oIQzqNcOk6T9lTF5zCAahBVWn87lMwy6ji4WzQOwNrnE5jAnLlb7ydeds9hQoE4J
Isfk8x7e6WMoCQPfronhGk5/nP1AqUX83psS/SQg1iAyBS6LqpWd8E/UtBREK49m
PqyZdJiD8tp63V9dquB7owv8okKjebKqBjYtmVgqfjrebwT68iwKig7zTQNtTZNv
CvSLZx26aPAL99F6XHJY6myHBTC4QzrRUAtBYsN1pMT3TXtpXqRZFq2LsBT6IOVM
QFOoK9L0Q7qC0bTOWCMTDDCx15Ksi6Jcn07bPPeXGAWfkYGg9fCkfIc24Qg/u6fl
FIahZX4KZPh6HPqTHzn8VVNXgz1ivm+Cu6AeqbN5nDAWmmHWeJXTBDIrKaVOt42V
a4t+gZPiwGQlGj1ymxKhV4SP7fxiUTj0qTumLTlUAYPmbjnCbfe7SSNbnZGKMdPm
fZ4HU4/7I0lYEoqMY8COjcfavMj3Py7p2v8dwVkds7TJBsvvwlVDFTrvT3oGW3x3
1ANxjD3GcYMkKLaza5IhQav+ueqthr123N4YS+NmnBNkWwWukbpFPrNbPMCB1DEQ
jRLNKnSifEl4W/u1ui2WAqhQyn9sx58xJ2ZRwDNAvpbBS112TkyN2KpiyIJ3c7CR
HONzbAO0dVWCzQ3DJxhSEYpy0uyByVofjX3DtpN5yDGekS7ZZW4LRAM6XV6TOnE2
3V4sz4fqS/F83E/hfQxjZsGr3hUG3B79rl9tVVgoOuUfh16PlXQRUkskjvH68YSH
AqlCdo93ykpSAzUEe0Y0VG992Cm1N6g2q2KATeMgPe1JVp5OsW2bg+erjCbBQ8WN
L+NbB9RzJQLj4fJQExdkEahpX75vcE1VDdpvoEOxgioqczvCwAReBjkX1YpbI8HB
LsSe/3wSfqodiHZbvklkrn29lh+oa6lx07DqrVrUxcijKMd6lRHdsK+WRF0A8eTb
V7pcHZpEo91YOa8cARhcr91y7FFBS0JVZrsz67r1wOMlGDHQw6qtxWzQLVYZx0lg
rkY8EzrOYNRIswNfkg9LQpzEjbHZONLwkNFtcqWubo0NIICN99+op2i5iVUyI3N2
SYjOhdMxM7xpL4OEYJifygvwpEl1lzu+w/MjShbx6CX2ty3GZJpPMmFWbvlUU9K9
APDMpSABlkF4pDd7AHg2jzUDz6UyBli0m7DHUr+Q1qBVmPMvCZDIeVb2kYJ2oN1L
Fcj0uwszx6cOJud9+WxOz+j29cVMehhJameKwYQsN/dy4JDrBT6lGSGW3y1kTcF4
BA8RfIcQZIdlb2M6vyF3366UABGxp3a3Ka8+YSMet68YiyCR0RPZdJUin7JWT5zg
3t607ifMsKc9rcvsUYn8kG0DwyBkGN4/DVNeF7MCTsJ4+6g4FKmebowXthD5eWby
26NJihK3VUNoE1qrBH7vle+eBYwiFgrwKPF3s0GDkxDBvuvzxGvd9yoDXY3xSnjG
VHzkutT+mrtcGvHiABSF4J++KRWLhXF8x+iGIaG7pDUQE5IiRjCbTmLWXakHZGPF
Quc8a3vMP98GcNBrm3+dmvCN+OhNF5BWi+hurtt8YRyXsdGZKTHRyH8iuHzG+Cb/
Sx2HCH6/eN+G1048DQ2PLP6kXZGnrQcJDr1bwuX2FaqwtCIS1m12I6K8CDxUcO9i
17MirKX521hrkMJmw2frSceihGIa08lgdtERcnGUvSHFuABwl/SAryKHdl5x0VDq
Hp5wOeUSPYeRQ5ODA3tr/ZtW5wHJQ8qi7WvDJDTQ0V2re4+hthcDVfhDw4TpeCoe
ml6qVLr/h5rWHl7VLZN9bIlNNLM/ULKh+knx4TKjdvnOuwBK/PaY9biBjXV049it
H8SCg0AORc9J3FLw7cPPQtqP3EVPIaWGdKIxKI+a//OHNCn13y5RzfZYCPJcQo7E
waOADUAmS6bkuzb5XqUjZbvV+3p851YaGoqbrJg1xL2VZ3Ei8S1bacTkKh7aNY0o
0by+YUxp46vL6bcO+ABMeXhBVPWLGggXf6CHZzopXO0OwWXI1TVXDVSvFvxhGBGy
tbhZjAg2zFoi4TaDEvek2fbbaOKbV0UY1JFD7cpyU61lfmdfp57/mcyhPR3X65bS
8SpessLEKfhE2kRhbwdWmSS8FZIqu+KkzGxCz24KQOUPmivgQE56CfCdAg7F/fjZ
CqC+JJVx6g48FqU77VxSUNLekSaq5kGIUcgT7dwyof0REoq6AD1jd8Op4HjgXObO
mW9g5stGOtt/X2Kwq2+mrGbn0pYmB9b3Xi6yV3RHoXgwpQh4FYTDLLakhOoW1A0X
sL6ibx/WIMUz2LvuHyJR68VdH8y98tLpSSDbcj6zA1mtGV3OtiGy6vAYxnV82sbq
bhcSk76bCYd0FYkZECFC3YFmig266dTQJG7Cax2j+QX1fgvn4GjRFW1wGJyRmstU
72ch45Fxm0Cbb4RiT+57X5ihHJQ/WL27G25X4yMrsC2zHk5HMHCXnuyENcy66cn8
rZcgbRWsFzq/UTis2ABAmd9dZ8/8plhPpoWTBswLszsIWUiBptQMhOzE5oNTIqYh
5vA1M+kIg8n84lqYTiTZ7DwHokqqH4zfH/uF1oRlnjjXDnTYeJTMB+Q3JzP81a8M
VwsD6rRJ5zz6SfYr5vHTz3x6X71kBVOlcCLWek1D4ZLRU+9LxOM3/OdHYplr1qj0
sj8GT9jEHxmOM9CBnHyixBuQImUXTKjSuKQGzSxTKtHqlP12k+uQAW+i7gQ/CE3c
qfq8XeDlyKRE7wn0DsFFrrUUNEguKiHdspLM2AsjwkrDLJFkhvfHnjqKsDdZVTWy
3WEiw/PVngFMhKCBvxRgmq9TK1BsYpnIkeFwGiqGYf7EMSZ1GPSZMTwvUq/xlB2q
+j5wcz88wMmviT0iibzQGlsNS1BDWvb7ormPoq7/bweccvxIIANpaEVRS3Ggi6nV
qQvxDiqTxRi/J6P8B2ZZqUk3pdx+0/tLOYtxEWPeB7x9VyN2PULY/zEL9R2SFLCs
3Wz+Dyfz6jeBel79Ncdpp8yBSnLvfh9UkeGbPPXh/m8fCKZO3VP2HQIwSWJHtgL0
sYSoUoelVOCgLz1pVqDzXWavGb/RkheJ32K7CUMlQwsEAA9E18J8Wn1vIFtTB99i
VDobkskGOYfbD1XgZvYA8GP67OJlGT9jBmjsOaCgFqybvDlkkC7ZGIJoVN2ZGfXq
7rWUOaaVPdFQi15mmK7HrtxiJ4H2kOy5QBUuU6rwgGAb9dNe/KmkZeMtdLKiM29H
LE7p/v2yO/Ywf+JQwXr5AS9r4vsDSwqhZ4rhwSF9ef614qOflAaglB94AokzYvx1
QoUV4/yMix8CgIIU2VhLGT4fjH81qRvW0ex2PXMSZmJqawe6BjQHaPFgZfVqR4g0
5xKbHL1/PTfJInXE9t577RkpnUYSI6og2IOdz8WizQ68nNfh+RzQk65bjNsjp6RF
7OLlNJ56satilm3yvYEV9nQ/PeIVcvVtzdp4q8q400MuL/4ATNo/ReXhF8gzKsJp
OAxtE7YK5JfKy0buo+1in/esxUL7Q9OkU1bjIdlnfH+oGBVR3yVJrP8KMNaW8mA8
/zuDA3Up29StplsZrnEWvzZyEvLUBfcWYzoRI4ql4Ob/leFkKKQpNXdMbX3jiAx3
nUsO8hPEs2qZouuyvPdiO6tg8cR56P69nZai+5Hx1lnqi+iF1ol3S3TsIWrkvtYW
el8lAKj1XpCGiNkHms4k6H2mbhsnhg8wVmp28SZSZhoEOQdLFCf16ieLUT7KzJOu
mIrSoFjwDBmb1p/b/c0l2HxUsxBSrnf5U+Rw4eZmN23JolZxq+sOkgW1zHIQlAO3
uYgW/qjMlUNNsMevWDEXszSzBNRybDR65x6Rw8sjj2hCxSZ3jiUbpik+pvKiLCwP
OZ2F6O/HhLvYCLevps5VT7m3qovP/NUF7mOHNM0V5DZhnFbh5urcXyTlo16m84Gg
AeENi+suG78jlC1skjJMaRKQpv3bKpEuI8dqsU/o9jXMw7fcSNnZt/fzELDyh3Jr
VkqztGHlG/unN5R9pS2d6nFCCeoPvmJhVdevDTfCE/u6AUeOtLbe9dfo0f0JrDtt
u320cfYYwQvTkgDABACc3X7Fp29eG7/RXQTb9zf2tkBkkDtp7UN7mrbCuqGuAgvV
7SbOEhlOz2Q+5DL6XTf0B9MTXpvsXWsleAFb/h5RDdulcZWKJSkUfviVbh6UvxHJ
PyU+cZKuDlcwkkcETF8CfJeTcZhg2/ueLdDywEzsT4hwm2t7NMLIToR25hX/jsxe
jmXK/wIJ1tiSFcvGXRxB1zkgVIsFYAg10pNePXwyWn2tYYTRSGbUbP1qJqha4bIF
FCkcnMTh6CpDBHox0FwJTgZPCuLlelOsL67ylQ9l4k/nmUWtCKwt6cZAt56ieD7d
+ZQQvUFxykHlej+XDq/zaaH1vdR2yY3kotsTusrQ1Z/vNFZ8u0Y3s5HDMWEsUpjZ
7J4FPUyVb/WRzUoQ8gj499nsxyg97gWYeIq1otHPLFYva/qBLJh9hcCC1n4moaS8
kl01YUQMtwQ5YuRDZIYbi4kQHRModyZa7FfwAfqQuveQjnHpxL9XJEr1orLjiEs9
GgXlVnMTUsEd6D1c0GL8JhisBrsOS6xYuECNpDqdm6KO820enISZsTHwSqL4eF/G
JQc28k87FiVjltEZhWdDABRQPvQXfAmwYiGxM/Co7nj3+geYgl3AcyPmh8uuQSSf
lO0iEG62duX4frVZI4ol0j2UnT84UBmMyRYvtIxjqkxbDidE5LlUHotlqjdbXz+3
Fq4zSwdy5X0Z/l9efJVJjdqBX8karRrV6Ex0ov+/gEDwupUcC6iEZ2AdUv7m4fV+
iHrujskRu6k5bZuW64vHTeIbu6yHwuAcFCJW8jmSw1RO2CXuxwqvstb8r+czY3FM
kZQzWHfl/m/1Mko2uY1M29JFP+PxQOqpNKKfzUANN2dxqrCjJ2QpM6GE8MTzRw+g
8u44TByoJcUHV+RTy0zHTKzzGhwV8eUNcgyPGuERY/hMS5ruOBenFuUNkr6NbN8m
eU45BS3pjJBjZTx9o1aIcsGnE1F/h+ZjTrweG1faewsQN4jjAY8Hyfxv/F8kEOJ4
EQFAaELN2Tg4OUyFNsWy7GYV5O+lgLuB2bkvrBOe8GQibE2kBU5JcNZcOT/cpeWF
rYKcfdeYUjHhTYZ1fl84M0nQrSp2wbrY1LCRHmVsdVTF8JKiT+8vBc1ucLDlev+E
mdrvOGICm43pBkk/icSTjbC5d1ALysXLArBUBZ/Rjx+OA4JjzKcno0lt9GJwd4Jw
zvUuLOJIkSpXRizwAWox1SCF+/XWcVkydzCxRqMEa3SWCl2FOxZl4VU972oexA6s
tNuL+kibaZaMnr9CRZj6MDcrNCtFGZmHZg6O2sRmq3RpV+Y+CZBa66CrBhOY11Lm
UW5FPdt2XabWcsbY7E3YhFVlntoCoEEtmSmIthf6slhKs/kP4cdKSHkpwYA8ZPdM
zNEfnrSKWRZKgq3+279PXmL/8DL/aWUiOLTKUQCOexaw+oUGgek5zwV32LqjaN4D
o0n6wsKYUhIakuqvVxWdXNNzUExDAcux9wBZVnlfj0dVF8BuXzoNcBY15ReVQysR
S2DmfacuWYXwYJExJBFyxOhlR3z52+3SxTNthGWK0hLLu7OgIsxlcXcbf3wZcCM9
dNHfSRo8WUYGD9SKWN3kisLeL9lYdOkizPTTNyd1e33mX81w+d1q4z5ehAK28xlO
lLeU7VusN3HkIthv1ujWc9OefNp7kO9i+8Q5EQM0dG7BXQlqRJkNKGWu2qhJAhlF
eDNOSFEWLDbXyeUEctJceapEGkNRwSNzwgPdtCIOXycxWfxKCDMHPKiBOaYEktBG
AOid9aZfRYRIK9l1MTZPVmWIa6H8i7vVrueDiKjN4dFTnR2rf9P8awYBPBtVXkFY
YPcrCqMR1LqLOoqraCh4fJSbZ50TEhWtpIJV6hjAz0xtGZsChHS4oG/wKeT0R+nc
GBbDPc+3tn5dkNNE5oqnZV8cJVUUSWxEqNJyiE3tByKwb1NviOrkjSrx2yhBPKXT
STVIoKPmAXvJGBpy9bdB679BCBUYctFFb0ckOg742DXKIf08u6sjz0MTfempiMEF
o+mAHIjaLzmrTAbB130Zz1dsRKb2oKwRpm2yNUY/GGM85TGIpCVt3ovCMiwts0My
rzHFWCKE3JpCTDpO14s4TsdhGFS3yv4uMV2+oImRDpuEFEP3T7g4805uDUarxGjF
C3UAID6VDtbdIOO3+7KuAoUrlSKYXB8kpXqoAlvngsjt4Bs2YL4dWj6UCns5ovyd
QtkH2Hgobl3uG4OJrvpFfd9L4MqpIPz+T8LspOEyg21lzyVWS36Cf/QESxWTdfR3
MDWI9F9Efvu3KbyIbmg8wlBRh9yYZAQ67eGF6oGEBqYQ74hcpVLIpW7p1ho1a3Tw
46SU2Pcv29xPMelhked1nhvNQorR7mKZD5trI0KfCdWGFw43sii9XT83MC89C/l+
uNzVh1AtPjYcknb6Lh3UILYoIVGUlgiWfXhOGAyQyw4W186I2yJHIWfN/msg9tyz
lJcTRX/oO0UZQHh4LSCAEZRhlTORKK8ULDXn6to15nKC30ACefygPXpWq2r7iiSg
SHmwBzzvSTyTe+bu+2rWx5jpZXJzTYx4kArTy7cT+ejr90kkxUQG5wahNBMXupkf
OJmPBxQdwalnP/0TRidQTON7w3F1Nh7JO/UndkfdY4NYjkDeUZDumISj/P0h/atx
/P4XwFuzGAoK68qVgNPTMMopPKnrafQLBiYdMiDmCRWd+Su32cUkg/0xGJ1unyZQ
yNlkUBKrWUsKBpgrTHGIZ5WPEQ4oLrvWFww1Qxfy2Bb82Z0SmPQAaqcfKDSUkAGt
HTivBFCe8Jhf3mcYp05zCO1H69xpq/jU2h7N9AcbiyHuZC4oQfcUeHMuYGAW+uqH
MJmwAzRecgPyceu+OvwDyOpyXqjPlrxpODVy6gB7/qbWU2Coo3rpVTVAmithjFt/
mmoMLt4sNIQpeev6p4PeZsrDveviJppUTAkaO1EbB4T0BtIPkZrdErsDFCUvaeRk
RUjSuF76QoWluZfpkLaA1Da9uZGkhPibsfDaRei5YiU0ofJZg7FTVRcwLdKYKH9B
sFDq85F95C6Rrd8osuq+SIknHt8pTXo95WQ8kkZnIl8vaswxPqMVSXhhTL52FThn
dIKKm/rctX9EcNF04AjwZVoH+9Xv4RVHWPAI5eydDRxI/I2SBD3frYKXQj+MMJiP
ePs9H/N0aV+17BkaRrc0usDs460ScBS5ajPOpwz3W82o48kmIEs7F3f8ax2S13Yc
4m2crHjqtapg+7+G3el8q/ECPQu3NMSnZH/HJMnJvKhmh5XR4LY+rEv4Xqfku8Mb
KuYjl/qkw7UoaSIK944U1duBZATtazheItTn5D3mqnhv2LHz6Pkq2LxKdJEo7amI
pSKfhgZqP1b8AkqI95RcrbuGH1/5K6QXkQ6FoPMs5UAgoLtznvmUkjZYo50WyAC0
3f8fE2l8Ge1zpspIKA9/dkOKf41A+hku/kdC3y0c120yoF8OuBk6SjS2wQO1RGmY
8licyIdEHZgjT+iXm/ihNuyTyfrblAobUfcPUwjWcsoj9CGLxVFP2QuBcH7XBcSJ
tfxs+Obp8wMBlDx1OeidTs88YL/V+KNB/CHm+ZdBGQ+0Bo/6W8cgdIdVIjnE+MaP
BIn6TwxiHjjQczvzLSocBl5K+m0dCNpvlYyimvLu+iNy3O9asJdWvETm7fCFk1S+
NBY4SUp+yu52YQ9PXjwPtVXPsMr/Q1gNF0lnbgqNpOvu+h+ytIwZdqk1gTd5K5RN
T/rkIz7CvzON2lNXs8y93gAvlTAVgrIA1UIRDU7q11JFpPyYAv8H8gYCh9d1mERZ
7hcipwwNEB5DTu1jx+hLcPDyzSeDxkjOQpcRCdQHqzZzw4NLLRpwtEAGv4sU5jJH
Jv1IJWePNXTr61aj/EunbnjBZe26OCAib9sWskp8VXTu0WLY6P5vWqB2HZHXcJLJ
Qj0OkF1sC3FBbtdwMxXQ13mnpxV8vm3Ib82wErueknhGByCCp52GBfMVBLqKzZuZ
J8Q5E9Dhmh4Y4+6H0oaTYnCrasGe8aCs/Z4dlTT1Dqxvdz1AmaWsI5EB6fYWzvlQ
EH+SzvgvX/OuHwpNy9is2DLL0wr9pcaetLO15NE+D895MYnS0SYrKAkJVcj1hpjh
GM0mQFvS+pA1XIf08u3Grylt3Pnr8IOMP6+N29kxlTTIC+z1HtFDa6+0Foj8ZJGi
LuX3MtfiVqo4F43v0EsZDkGOZ1Bgf8Lp5q+DwP6BcAxj27w38Ou8QZmLtpZIGlQD
B0pVOLWMoVTe9WLYYWviEzzdZeUQCXaNaRmSOHy+JJnHWQwPbgDH7n0+r4MbpSuk
NR8se84vMgtucP9nbF6d5XBWnm7gWAR/tf0aF3FQMC56hrhGkX2HEOpSkNnQzUvb
0355j5V1qKJzfTbHH8OQOK0zs7KgcWWFk+9hfFQD7t+XS3izPXxV1afzqjewd09q
esHuRP3muBY7BOOTJAnwKXtMJWtWYjnwOGciHGIxqZQuSHXrj2eveJ4sUmIvlt1Z
n08muV6Z3358pS1haXl8v5QeAywyyjC+EeE1QpW83HQ0hgr4fprqld1mjslbjyK0
Jgj3AaWIQMFDScxWFoKvewH1GkRslM37vg8saUYBZU2mZJmquRuOtjSbpWLnBPIZ
HW5Pn8/P+df21hyYWKvV5idQ2GjVOUc/Ir5y6zwIoa9yvzjbua81Wo2hQY6mwM/G
NJSU0IzT6C4K2KsNmfgnWM900w18s5P2ecYBf1h7/SQYSGKloxlyQTfkFL33gC1U
Qka+4LVwkSM9CzkH/GNPieCizc0rlyhI4IxUzRQBov1eeBIy6Ohx98cXTfvnnw9k
CAMiWOo8k+eg3+lL/W6lXond00odLjWE32g2lPdp5gGL6xgE7/Lep9eBB5X2qzO1
Wp7NUOGwXGGTk4RMSOEQrSt4PHhdmZeEvYzco0zvg+hDLsW7FGQjSkZBF0dy4nBS
I2ThjX+D26tCNxDfHvR3Wbjdga4wCzL7nF7KXIPC1+93vlubatRwyIFgINnn6a4Y
57/+7plmd2gogawu4pQohUFH/xVfyk3z223q0xZVj2kHzMOsjbeZ3T4e2BIkNhvQ
y3pWvFTSJTZ6OV+/EdFgJtWEB9Dvyb9iL6JV1OgBwp8jITGirmOACZugcSWYsIat
1mKFqK05McUrR8+TQ9pCm10/Bj+eUnKnFsG5zGYlqJyCoN2o9hTPKVJDR3pgMXl3
9KzkxbcuRRBU7amaC1PUfn3iUQaYG3cdecrShDZWeIn3wL7ARpJTDNvCn7X1RBN3
W+QzGoqMOUdl1iczaj48uG9VIjaHuK5frAcqFUu7vD82PlsiU+EqJg1JT2YQHui2
UtcTRpdvdpeFkTRGNA9cS/m0GaADV8339IhgZzUBE4chnVbBna5W1QXgL88ewFFH
N6hsULdyukGRKEa8obkYiQE4ULmxenOouXV7oOS+NbCAYUY49Uz7U69hCu4HTUvQ
J7t0ZtBQkLfnhqOn2BlHfX0rWeNEikwdNFX5RZsIrIaJygI0u39bnTmzvvNyFqlt
ahOyknNmVgHZe1T/GT8mr/BpWS/f8c8VqeYz7mTUO2zkXl+61bI9FYTZw43fLkKV
RIAVWE4TipOVoc45G6MULoRrqsBIQpNT1u2sX3fY8xVV9rqdGatj3udMTPVbbOog
20Oi6SxQ2QSMZQPyzq76yHHbk87LYhnVzqgUDY1ZbJag/38jeyyzEmnRyRF9Qrsc
Ngec9WcLbz49ExY72qPhtPtdqy2lOJGtsWKoVPTmOMerZ6eYulo1SpVKnDKDsBgL
MEiEfI+LGe8tRxNX+J+MP/UWN8bDBF7c5pO582n+046TK/jZL0ZITYatb58FXxP1
QzZESb66wPDRFDs790rwMQ81EsStiqxN/My37aRatu5PJ4LgXZAiX+FqKkRLp0io
ozDAaqbLVV85ndRrJExuQEeymISVoR7t6z/1ibjedxD0oAsOhuEKgf6qpX0riJUt
NP8K0mLJ9iPKHEBghCBD6VtfMh9wxlIi+OeUIPuX+OTZNqA7wMlz22y5Ugsjw8LZ
aMc4yatbediGDWc8RLgerHqYnn09mH08fliN+0P0LnML3CqoIV2PR3Ih8WVtAxcS
bzaRjeITWOOP1iHrgL4Q5Gy8eTKffzddz9+pjVzwRLFlN40MB6fPCtBWqbFghYv9
altU4lkJIFPwes1SwRfs46ngYPB7Rq5CNjQaU0uSaSRVfcainKKHZqY8SchWKBd1
RJz4uc2UhAE1sd5oA0r4vKW7WSv8rHgLYlrOeoT6VhY2U6uCVy5BE7wkCXu8FNZI
v93fESNLBTI2ObCanMj2ireULnxjlvQ4BWKkuoFJO8VCbIMboBmmrQ/xN6eZ44Li
9k/XxTyfBf/pDIB8LsFZwdqvV7LBjD+Dy89EdzDU/M3Ekb90Nj42bLt77ZxNkldI
u5GYarszdxE1yHQkYxx8kFWDbOKytMSbQIqHPlz3g9qDjzRDoLPKQqsSmcYMYXS3
bgjVic1Zi1tVB8xhWxHcO8tqmhzwSYiwXnNsm/AUuKkLK1oika0RrLq03IYAh2bw
PYnZSmgn/q1rjf//DSQP6hUKf7xRgOAwlx2gazIOsH7mUG6czidhTyJCp2fT3kQv
OrZli5kATOf5ERy/5NeBcjK50Hs6679v7g/f7hz5V6iwiQDixCqWy6CxCH/8X0MT
+zDi2ElbroACxlaCJ/pXeVqqXhBUJ5ho5puGt85tTVHj09O7GqhLT8CoplEIRCV5
ya8Gph2gAGkurVlZDK7/G1JQrAwpg4JS3IRSZOOGWBOvHyKW6bfu4qDdiFLyZZio
fjfxvpDgSSNAD0sHd4KI3LeMZFeXvyYNMPW99X3+W9P5HklyrtPbnWx+wmk4jugy
9M6yUGi6DESB3x5aUQ7TkW5g4b3pXHh0GDX4/dhX+E60QlRJszrbVgqe2OBLP8xg
hZq85uQDjvNNnSU2gF9bQXE9b6+5pSZfRwcwDcAlOfn5nvp61IimfoYHnz5CzIMR
NWYikOtFfa6hmKGN5AytTcNddSXc1Xqa35kIPnfSmonbmXCfPXLiJYy60uknFHtY
RRci3zG8tEuXfDe5Bbp8iIzUyfr0b/i6eRaiP5jtatltzo/sFnic5yrQ16ZpyiV0
9Vwv65TUE3Ah5fGZaAg8UzgkF50gU9C0XUXAbgn5udNYUu+E9kxct4QvzH9T6Lo0
JD4rCtRzTab9V+LyoV8IeOGzc/6vEmDEcUmcB4hqaHxJ7MOCvYAp+r9joh42GaPh
4nLNI5AGAmDW06yPbmOKl4TrJINRd4Ygetg/qz/AXvSIM8uqK/uBO8yF5duCYKet
OKTWJJm09mF66+9RkLjxw6j1mu8mdptlqNDiCqj3CBdXuvOF0nDzS7zickLYaiYs
EU8QAAfqKdZotdZ+SejtwjnspGkecolPMPcsJRkT8NpYpTZVv8Jo8b6sZHvj6RK0
VXgtlKcKr7+xpNYkmzMFXsLczlgCfdO1AavRWPAz8hIW9slwpLH8m3RKhdt74/7y
V+Kt3e3MVHOJ7ZQ0Up/eUwgg5gCJv2TJw0ZK7OQMHaHuYJ8727c8t0CnsRtl50HO
fXueq0wYAdSeljnPBX8JsvnK7OT54btIfg5c3pu8kBl6LRxVfYnr7L66GKkMecDl
41fK+Ob3no87RpLN0lQpU0IkzMCczBZGTt7+UuW5y8KR33tTsu4Gmk5FXnqIAAYu
Eoq9anNxSC+cycmdIJnInpOTm5CrWt/B53kuoisOYR61P7P5M8Jrnnjt1S01mqB4
icVIQLLAkZ72MFfXwEm2bUJywYnEt294udCsH1mPVKnIfmJ7ToeJoY4wvWmK7bJo
KQdz1jm5MImvRWq9YpozudAFyiclo5071O+YwF7FwOmjs9F4Hz6muw/AhFHwMj+8
b0U1U7MjVBxjjpZglPsxHDIAV+EEBqjAf/ouoezQgi4ovkDna0E6oSV8zKfcz8Qi
V4usf9MRfVmhU7R5UEzttFlCS2p2egWsNbLzldYk2BhHgX4mpVxs2Enj3CJ4eoef
D4O5IlRmcVDoa0YjssjWnnXEW7bl7cmbZKlizrPoMbWT5Cebo+nDuvkfwWXXltxZ
v+llJKt+zbzeB0GdGDF7hh7EiSumq52N9zawebXsbSClIfAzR3VIJi06AuR4lLzZ
DDFNz6Gofk5YZC4NwJlWWNXSZpHxGykoBGSfSS4JJlcV6xcrB8UUGKN/SMtTcV8+
6VJtt6/LYxhvzp1fzA35mApMeZlXaMx/GCXj/OY+7K6STsdnj7Tt8S0SiIHEqyjX
yB7eMSHHuD5Fg0GRqD3T3qMPUvBdphJfgE86dg3ltv1bzWEq1E00KvTQdH3irtpf
ms7VZvYjRJTaqCrOcFiKl/r9yUvvsyFYnfsJ+e+8oRHXeVcanW3U4X7fwPkIgIUe
5ycjwlkp5gL+nlJLqOT5k86MWZE9T/0SAXjkkC1PkqxbEqRuP5BGUmt4a8CJxkOs
DbZbfaqovTszMngtOagEcuL9sOAhm559RZzhi0kKdtvmqL2D3gGNmPFBDQj3XOKZ
TfawmweO75Dgrqe7ZCmHrtRjiwZ8ugBLeSonRI/3xM5a+TjQy+rKac07fW3yTkLB
7n0BXWque6b3pSk4C5YhnTC6ePT60LjSpF56qOiHC9oglEMVPIgE73Bvgo/m0One
rByV6iXqakb7RlHa8dWceUsCEmEI5pk8oADzmjEtFrY1OQ2zo6sLyOLNcikOituk
zNkbTXjZf35VzXzCxpO+7RhYAlFCKOYcpHU62QV7gV+C/NzUC0xab/FIBmhzTcBS
b38O12y2iq6lEG2FaUI9kjJb79UX45OrYwHQwfDNmuqDtWF13gPd749ytIGoCscz
54msWLIYQOtC0Xfi31Ggfi0ZG6jlKQ3L3XCcOG4SXsz/RHY3CkOVxnTaL3PXPXcQ
u5Vm7Q80/gLDmbaWSbureC1pPtc9SKICRo8q5AuSzUY5a4KvYK1+Wub/RyNnVyfR
ldFrTPDIcjfDjaC4RSZN5wRZMQjWBLlKnmkp08P8CMoWbc5B2LBlN4jyKbtsWkXo
3qEu2PGQW3OU5ZVJKCk7gIKhT65oqtRWWILF3Hl/YNa1P9NW5Ak2Mokdu65l4RPh
jjkfnMBU06KseRl6qXHKTLoyEIXHeXEkueoB7YKZ3/pKaMEaNcqs50Fm++neJJgf
uT76ZK4BHJZPbbnyutKFWu+X3jgqRvm1R/7OY0/Xthua6I7oZn6ae0qkE9zvxT+j
6sCVq6bkddv92uoSFBgiGibVy2ZvWqQeT6FzBLRZVOH7eR8QdrYs97NpDuswttnx
yrWiq2CVLQKm2ZXejfEUqbmA6o2SYlVTZbRFVQawfbMOra+4uAYSXMqS8sv7Pwtn
nHbTl6xC4uDEcpjqQ12uv4QiBUFQ1AW4zyHzPX/AXGFjYZMQEUJhUYzRNEZR5P1c
eHFGzz7Zww09ga60WqPXJjrgMHTuAOTZ6aKxfPqGvQ3Frtfg8s0/IbTs4TJ+GR46
b+pN1aNiKw8USTeE+6clHJ5EAj00RkpcszCMbWC0hwGnmOJ2q4grNWmP8FDogxAO
84XvGqilZz6spLZVCVtsfQeApoEa9V2tlLmFfqv7aRhlmXSBKK3pNxacAFIGAEJ6
36ihLxVrRqqsJV5QDq9BVVO4hKuaSlVBgn6KQf1rBS7OLShzpCdKB19lqWJgGiH3
roc83rsM8OwxnzrJoPTSsDM1QZodkYopy7x4/bQdB/WlkiQn7hLAEtnBJFKwLytJ
IpqG2F+UvuFFBneuUlamSxIuqf0T1XSfFnHbwHjpapsySV+wQ2ZwKIsncNwym5nF
CBx9fycUo54EBhOele16BnCTSbpuJfjLGUAdFsdsjV3mUP7o9uSqTdwzly1ggxy7
KyXEHU712zrnWDwliOD+k4DzR0qh0dg8Z1TWpZxDS5Dx0wxUto6YHWCNxqYodCiI
GX9XFgKMKRokcf/kghRb31Lo+ETx9oBmUyn7dL8s/qwvWGEq9wIMAe7T7SJ/xiaJ
pfIsefUi9jpr81EYz7lWhPeKnaEZ3v/m+IaCXiw2b6gZAmVj7HYOMROm3o3v8b8u
2meh8yVR8my7MSs52mAHkrgjR8CZArHkN0cKNBIo147/kmJHASXnfsri3Tto56KM
Hy1kS1NR2uRDDIHfhMN0yAOwHcGCr+x/pui+R5mcAms/rs/0ErYV9jf8ve8KsZPd
9VOt3Hz+B9+U4JMviRXoC03nSsqHy+Dqiikr6zxRMhWFb50gzRxYurrvbqmxHe8x
GFmjAQbKzB9AokhjCMFy0uyfbdPzfEdl4mrZr/4y+7ZKhvvs+azlSYTSw23+e/mb
P1UGumPOEyXn81LPxAu0qVVbp62pL4RupvLkUUvVX/xAJS7Q5wB7mFFR7ff6ipb+
pPk1poLQn3pvfiFq03ySaQJZnSHwX4pFytsqfSaKAtppi/w+7iqMLv2HN4YIRCMb
GFJxqpRj3E3wSriG5l9VNP6PU1VCU1QPcaO+tUlOT/FvW3AJqLvpUD5qYaE03ros
GUOuVRYYVX8ZQKRANF9YkcYmxa1IzX/DX91DLaceQ+UAbDSc/cg2CU+iBScBrdMx
4acuBQtecGf6pqRoRIfsohRnrCFOMcMh44On5AvipCgFKs8/L7N6UZgAUkOPfAVF
VmL09e6B+eUUN+K1Ev3/e/sWMBw16LpWyZ92+y/UG8Xda2ndeLvnc6sr6Vgr7ty1
0TG3TJR82FciZ2ycT4+bvhGIIgUpY8wRrvWb76Ie1aKTGYtYOPNdQ+nk0OjNktVh
8CjfBKtOfN6hbbKK4Uvvnqh9sFGZeNp5g8s0s/ivphU7mwnuxmwbmd6Pxk+OS5mH
1B1EuxyyLhWKx6CJxl+s9r1rPU54d3Ean7ugARpU/6Af1Oj65WWDJly9wHbXz/bz
1KKCauMrSuCEAiUQE+YgTsukcKMeIbfKB9/C3slxjW37Ni9gtTcxADHGJAuOMqZ5
P3O1bSWd3tsKkAXYA+8v6b3rpKOD9VaQJoq3Pn/wIGxLm/Tg9ZRgR+tCjaU+sUpz
hQWTr0VmHurF1zf0RnYnuRejXGhEih6GQRHAzUNgpPrnGbO+HxjLWrcLM3zf3RVW
b0butZtET6M7UQ+A4Tz+4SwuMTRyHx/2vIpgwpVGNKOvBs8xqg3RxFi44x0khbRJ
WV/BCtYKfidcHi/nNXG/TmhU5PdgZg277L49O81LbwbKpAUPN2PhBPBgnZPlhUZP
oIH+qYW/kTAbfWnhS2anNnkOBOiWGzP+zPIGHmbUfLIG8eZczPaMMyzcIdkp9wgS
Ss1JEe+jV7b34j/hPQoREhyy9QPenxj/NQTLIDvj9Wg8hUN/neOW2GT4eiRmJPLr
6jeR2utvjq2xCD20KTnYvRIPtwOEqKfSkXHgmvWmRxIMYzjDn5aJevQ7gzvfbPjL
00RiYgRZGyjQ52ENAjpZXVKtLNCWs1M0z3iYVCqc++vZBVqvSx2QQjC2hWvjcOmb
KL9rLQ1vcfBfZiJTGDvKKoFxCE0tc5cIYcvog+UulJq5k8E89Yg1NlNpFbkHLC0x
Lc1xDzj2thmK/vDdeFlFzQIxktvL4f+1v4JoksMseYVF1x8oEQfmIEZ08vi6haMJ
kiHUYjmKvQalRdnFc1KhfpMATRH4wbNgMXN4Lfw8CPvRI91eCh5u1ILZmms/qFJa
/+zJeBeR1jXu2TshEDbjb9b7XSNY2f0CYHnICsYiZjG3eRwG871EGWAfIkota9AN
ickt6WWRJdbQ8mA1knN6pnXwOM0BI2lM5BO7CqyxZU3eBEYPvh2Lddg6zt5jbulk
tkuQsmxJh0ID5GMufzAGZvprvw7X7XeMMnSr6CkgC4fCX+/d9KVnw9PgzIigun/s
UP6WBlqx9FALrNYoMZ1dnF6e1gO1kbLR16CawM5lXQwGlVk13DGRKiHzNge4Vv8y
+UhxlPSNxYZFZ4OXQR8mOyJPo29ScqT/z+lEkgk9QoJ2ZDJPKCsR3/chZXsW8gNQ
J2uNHO+Y4NVpxfAaE9wVZUIMUZKv6uMgeknNu5hNlw44V1ssLzJnwh5AJVEqih9J
RJ5QMZhGzoTUzdxjgBPc7Usn/Z6g8nQkKdnKYuSXs3bI5oJ6dsDHU2bHNimGfbF4
oxMugIAtJE/64OclNsHWvIoxzp6N0fOzRqChgQX+lk3K1qCp/fdAN07uEtOv7XFc
kaCkxwn/3WZHgWVd4/qf/82SwRUVMhleVq2vrMLbCI6mzDp2uvbrC7Hl39ad903r
xwgn2F44xPcby5zfh/CuD/2zmSxSU3FbiuwhrxSgC9FpRYO2ei+5VPE2TFU1Y/6u
hn97a+MlLNxZ0zkUFFofUBzrkkUPec6rBggWxM0xJIkwniARevBAXgpWjOqAfMwV
JmokQRjXLJmqYPknyCJSsWq0+lio+yg1U9gRJFlBQjp8kdRp8DT9bdPN9knMdvY0
+vRYFhAH2ZXFo+U3SIYs5+koHPbCB41/yeK2cwSlz4wYnjmIT1eLadWPXKHM5MVN
sp1MrJtuteYXIudpQX8TbQkHCAuKJ2mUqqfiVLwXHIMXjGjpUdSVv9WgAh6MKw45
1GnSilCz3BHy5Z+IrQMxNEmCBKAxkXSar5w+zgKn+yPW6HaomMS2pIEdzd3Kw0BP
i8vt5598SoYF7AmfVCuyC+VllJogInX2ehANnknUd6O4qL+S0S/6A8LyJiZmEomj
9RubkolwBnzaOa/rMEHIC9yTaZiarxxDljs3MxuE1T6GGfkZEd0A7UEUMdthyXwz
NV3g+y4DvrcOldq6jUK+xY38KAlU/Lc0vCAtxrFL+L1qxHe+qXFKkvm6FyJNvNy4
kAtQAvKklIc/ej3ZBtE/tyfTLkEw/wIjkJIWvVasXFQlvRboqra9YuU3k+tweRpx
UOVggYiRQPlDf1swFkq67K3afMCVNuERQkpCFvopNrLAGSgMn70mwdHWwLATq3ox
O8C5GZZ4R5CgBnTfRgGAhLRyHEaWu2XAZv6R+qaAt3U1mukrgWGJL7fanv8D4Zpp
osd/At5p/8UttS5VHMrcJ+OAFrjN1M5O5pRYvplUiUkY+C2F9LFYb7t/CJsEaLKM
uuoFv8LtEwE0JvTtyHIJIr9kJ+44tABP27oTf/4E/uDxFuC6qYPLXq5kzYf82C14
KPMmnFIMy9xd+x8tcFv1/u+VxV5xtjO3tNZOyOosFtvspBS+bXtmZBo9caxvsOpG
rBtTz/lSXje5ezt3pgs2WLris1Ypk4lxAUTr1MhIWVsccTuZZQw8ElcW11+x453I
NzKRRIY5NaCSD3exzgga8UCUFXaQizieTtqblIh85/9wSLOPNslqQs6h2IAYe+uM
DVlt5TwSmum5trfjw4R65Zq6pZt0DcB8m3iKrUF9esaufZaqCQJx+iklp2SmtDkG
t+KgQFBqd+nyoC18Iez9VA4a4qbtXzJhyIAHxDilrBe019CMrQ2Ptvf9b60B82H+
uqf079bYWHosQ49KuZiGhywbvYgngxBRFdjuLO4EFm0ijeV4hUhzwiZHCoQXRuNq
whWWA+jAWYPMKpOtX0veF96PDrxwnRAm9wS2sqJcR3GaywYFptMja9Zr/SsXYNwH
tuR4TIMn1+tUAEGizlIqjomUBINEnSji86JEwTRCA5yI+XVO7zy5wHuXvv/8jnnf
1f4fFW1SB4ce+IolY98qttDA3jTn34YTsGf/Mf8IgymC/RAjyGl61bnmBAOUuNew
EiMiljUgHHdBj1lhqs2YP8rS5D39IasOOYFS6HCJ9885jY3W9LUe8WtbbHetS0V5
ld/J8BQgYrhxlbVp6+b0QIV2BqqrS2bL7deIiexK0HDyGfIOXhPVET6S9pLwhq8C
DT98hX2oZ9Qx09bGeyRzcBjSNW4de3gnyDEV7ZzPD9NpNYY8kWc00mJZycdN+0rG
ewtX/YWMmPV8PgqvvHu2rDAJYpnBEx/kbKMWnEetcPQgOcoc+B4qhK1eV3nq0J7B
fsvwXsLJ/3Mbq5LgpaIeDZZT4JSGx+/HTwyqYXqY5TKWtSm43v9BKyxWQua8/4jH
iz2vL8Gtaj5SWcZrWthmNXZ6MGfeujh7Rpj45nbw3GPaSr5nQ3C6rqqDRXtn3tLm
i9ZiKZzlrvIOYVOYXmm0ZIqydGVHVE3MeeeypnsaESUK5UnCtbFiZtfwIDIZvMED
heemGUGojsmjgowFj5KbgRtuRcQnTJrs6WOR9EsZREsKKsNPoaYCPzFuf6AIf14g
YEBVPynvX+TOGRxCiXJsEaVDg3/1r6oLw3uB0B3Syy+gAo4jzuOHSK9/g5/qqF11
4HSAMc0gV1bouE3khgTaNDpOsYD7a63rSzaLxY67UIema0+dz91VIcK1HD35q+jg
xyRF+kZIIqw91/f9X0F56/amawNLlFu7ibtaQWH8V2LQXHEn+8fAUH4IY9Sgz4/I
oPniOr2KNic/BTDtzjK/697iwQRcd++Eh1TKbHf3AVL6AchCcmvxZfybMAsW1K59
4nb95jNoR8stLwpdlPhoP7PuAm/KL8qNjmosg6lfmnkmnffDk2SKkUBBgIcD6oce
7fxIaTWeQxliafAcS3vtjSMtwCN6pZII5/PjlWlg/Mt3zyCgZlpMpDHkCTUrkrjx
yxn6/w1z10SOE173elzOQs8oLUXdtQm81CjqPgNDa8YzgGpFZhI458uGwnYPyjEl
gjt3W6um20hxLnMp+p/HQdFR3rAg3//bWUf4EfXfFSrlOZdHUmJOZTp+gjYJz6c0
dbmkyVqHY3DnN03flN0xQYoG0t0V4Kt1RAlL+apsYzQXntmwbEKV4dKmDal1impj
8pbWpB5Rlf+1jpfaA6VqrPiakWXtWhVfrLCmr6Ftsiu2FINcKGR8BBq1ZAsEfw19
/h7VVU9kSR9Q+YXKyQVp148B21fV9f90ptenSG+Z3B9yWSmjh6MnNnfOmg8yKLj9
99Yg+XyISonm6OiWXU1N/o2gbVUrzPxuRjYB4xxQqt4i4L/z+GXpTOvjaq+Kn4Mc
kfrjLibTdL1Fnzarp5aqEIFTS5gQbQ9Ir8xUmmS/BbWbsUJCfw4D+8l9EF8PgzlV
QASEVEmRng+o+9fqmaZJXYatGoDq4aHvRoWGmeKhT7Gxl7qHWAWKZXB7wdH3k5M0
I3XYCyCm1C0i1tu/z1mfhZZaraaa7Ya97/+x+3EYdEfs28hQAyxs4YUEAVSSyiT/
9SAQXmrjWTerb1/Xaq+wHt211F/NQgmIBhIqqUtV1ux6JtsacKwNYsnJbwXDZrDQ
6Mf3/VXi7GXfl8GKEytUvcxE9k5Ro+Z36RgsbmjcV8o341yj+giLXrJppTxTIzqT
zKChTEtRiZOpJHlmHOE1DZtXQs4URBSYvPQAZRB/yKlO4ej43RdGWKjpL62qclA6
+A0+v+Sr9dr073Vt2tcZRkoEqpJl1b2k6YjND5Y6veFtXhPv7dgX2GX6tW0ksg6/
xPnwlaIpJk4eR8dL53Jeqe1BUw1acUOSxUFahmSmzfm6QZnmvkvwyWtGurKydDz+
XNcbfsLoFj2Pf8CJcq7lVk+5CvCRe1NzHRIi8Tn3VKL8PqEWdURH2H7MwWgTNoHv
DmOh56CoGoKXCijPAdTgxvc4czPbG7Za/8hirNZDDmR/E5JPNwFRun0tVPivVcgY
nmUVEV3o4bcRS7l4mON3S52YPp4oaK6SW7HMrM17REewCWY5YUDHqi62byne4RXw
soHGxkdnJmkrmg8foD/Dzr9Fp6yer44/p482y9UgekmZxrLmjo4ay0yEzhLkCnnT
aLu3FLu+M/M+Ad/r0UOSlKgktnFX/TCJYmlxHqIfEHuKVCgyu/HEMHsxLjqdFDu/
kUJN128BqAqs/ZpUtopQ0TdEgk0LJzIBkB61lX6KhFSM6aO2Yez1DSalX+X/mING
Su7AmQZzIlRANOHPaRkoBpAmBdwu8i4YbJ1MHiUKsHVe/y9jo7KSnr+X0LRdzNdK
Wdfe2HhGSTrJpHYsgB5WwY8Q/ONdrHWJiholldiDxlAZYqXkFaIV2Sq1mvkIozr8
/JBg48rK6zf9ynuUKwun7Wz/SuWqxEKo9nEx6aEn7zLNqXdcJVyiDiDol4K4ARKq
hBG81H/iSGuzszuG21+Q/hAWJxseH+ItZth6u+6hxQ+645w4XJykcGuHpMf5V8x4
nn18F261MbJR7hZUcQCYT6UTlwHG212soGD8GRYYshXCCatALID1pauEV6grI4KM
IRo+PVvsgVio2LTnC9BK7NZsQXgrQzGyAcBOJEszAi//1vQobvMC6L39PG1/2zRa
NHEPbPcW2UQzu+V96ZbEs+aP0lCdzvrqWDtm3yV/lx0OibTSRQ4WCQP6Px9H7AGo
wkYAUYO9p7mT1QRky/eqLKnuKXXAyqqinzoHUKAGJWZHDCBlhWZ+YfQmBIJIeuGA
J6hBuP+4TXxC8uyUYBBPQo9pQK+dKklNyQEkngJJv6DSkxBS3tNtqLUgk+xtzOZ4
fSrCMxWLssCWDRaGOaGYUv9ybQkygN1xHfvFAxs+Ua6lcQubOj0IBJEl1Js5+0KP
JIAbP9VQ4GI8zPUojCbMn1VET903kQTkXJHvnD/WqyG0bNcshijlsP1wulp2bT/D
FWPrlyw+pkNo3ObGssRhe/HUtXaRqlJu4qmH7SSAeWDE/dLBJ4ddP8EqwQpAX8VZ
y0i8C5/2P4cHCTFIJCCjxs3sb1HO6zqSfMJH/wTjfwGJ/w+tlshs53NN23EiEIb1
KoMtabF0JoTxbX0mLADb6NQdKoOLuk3FvCxkVzjyzOHfe8kmBI/s5xsEJ7cRXo0e
w9Wa8iCLJyFfcPUmank/KP1SF8ArkmsixJuV2+2hm5ffFQcP0LMTIzAYbfcNRqfp
pqXS7Hz4xeDKZ2fD3wpVa6I4taWNVYYtIFGJiZROvqEwYky8iVlaav3quk9MYbDn
vH4hBAr+1e6iZF8ABwIljSIgjbNYuf5L9O2GmkMYvoJ/6g1bUSDyL4tb3Pr1TZvI
UPeZAiNt0Q2dEILS4h1ZW0nzWprQ7Lm7/Yv7e72OBVH2NvZW6+ivpvM7a18a7QdR
iX/L9Uj9jUrZzjQmy1BH+3bDxbqke7WHqs7ZyT7GdmJnR8cr+kcAn+/w/BETshbz
8r8AGDr6H4GuzxnHTYdaWokXvIfeE4kny/WosJIyyZcTa+Szv/GfcVCm0TOd55Wq
OapJIoBlRJE3b6aM9QZMNBDVn56/RcddTR7nIYud8AeZWohNYzej1Iu2IFXEtE8t
mu9E7386KaG/ZqcMuhYugM/qTtF622bYjyZM2QzaziD3g0R2SzvS2pyMkzu3eZEI
rrqLB1gBL4xNKqW2txKDSbXNvKp3btkp/teGOqb7fCW21VDXrL5Rm763PucHD+Hh
9lN37FYSm6hoT9XC2DNGnUz6gy6VAzKlCQFzW+6jEAFt2P1pzIAaH0WTn7lahLTZ
V9tWty++7nw6kZH4rHmuvvecytg/BMHL0bcH8zXxJ3fpTBVr7vlrPXskfbrFDqPA
tAKS9KsWb8Lxcqq3UIN5fxDwekg7rugkga7o/gNeiHpTe3PVosbYRnXfmKmejvd8
nuNTUXeWvO40g2YdkWnZ7i8OvwpjPXgGRWS6wb1JWVgIH25ng56cvUqyFZ98hQDd
QL0rYc+5qQ81iW48MwL4XIyvy51ikFqpo4e3k5pMMfQOrmblO0OY+zcWa8EpoqhS
8Lhs2cv4aUBMf1r9rNhqrNHTHy8WOTWpu5OhniVQDVGb+JBq2xhlGKSkl/Rap++0
K1bKojgYGokcvVVAHDUPYJC5drfQoIRICks3dR1wmNa2+7Cqej5vd5ExC5nnqTpe
jT4BveNEBlTCDpdDLq9xs2z/ANFDihQJEkb1x5Rf9USNgwmUNtVnLBj+5Yqs9qHn
UX0/Nd4SGXZhqzgufkRLCcZgOkzljMg+c4oM2HGZenkxNZjKVQyURlWT2SUGWN7e
uBwjy1DlX8DXEoUPFcQOIfCdH3m5fMTc1pO++NCMbGrL71XeJUhxSwfeaUQYNrat
irvwu7unp4dPiQNHTu/TllOgpYU7AoBcRQZHjPklRbwD8NFFS0adCpbInualjsVu
8W1qDhVHLMm8fheWhfIp3CAGGepOvYnnIz3ak+KQNBpFQPN/fV+7mLVbXfYUikEN
aVXEy0O8CVhD7HZk8rdHmSVFdFMRGccQ3snEs/QfwonI1XRYJNnwBR9GCAXLe+ZG
5SFu7tnrnuGTpQNQ+oMNgqlv8br+6fQ1j4OvAd4eLRLpZEa1nb2LuFtmOWvtkmdF
ehQI4EDI4gUFAiG0+eqrMbg4gbVUcN2NIKBenllQjWWz5hmg4SmSIV7q51tRI8/f
VVIXPdFbcWoRMP5y5BbtVqop56hJnDApt4qd+8x4+w4R2DcMYu2KeX5Sh5hHCqWc
bTPRAKKwrpKqr5kUhmMrxLC9HPq5jNHEF/roJ5LxCj6kanKeuOlCkuKq4ioJGADS
o36T+glTC2iBSC6WNq0vLPVPKYL9jRdc7jnGqMvb1TwgogXXU0FM3jdB5I0XgYs8
Uq2zZZsi8pq0QUgvqIrK0qgetiQm/FJTUhCmw26O9l0PWq1S1a8AyTlT/lTNhcef
79FT9mkRQVUN57byJskPju4HkBrhQG70ACxHM70Uv9MPpMZ1FK8Lrq78DEWdz9Im
zXqUsmhRK4ZhFM/yPbFskw/kuFcpkTEyxk8KipRdKaPgNbsYSCi0G46Koad+UY1E
YWKLWhsA+1N9uB7BP2R23ONG48mDTJAPQIb0eIhMWdrrfFs//ak5WDPAnR8nTRgW
iXaGxm5Jk0/Im5Jl8aSx4dhfHa2VbULR0EdxiqMSVb2+7xcL8O6MjVGDN7sXYpID
/9acVCBdpKicEM1hPBiPMCh5ExKegKulwYxz9UwLbXRQ8kkdH+UUVyn3xbRarp/2
kHdxJoW2JsmP+/7fW+B1XGBNZF1H2HGsJwu43lBSXW94M5WxslDvEnvr2KYux3DK
IQ1W4E0ZEAAwFlriSmmDH9NUT1c8ZEdhZE1E7v8qT8fve5iKaMvSSBEs4bmHXyEZ
L5oLoTzVkEvDHd/BcHjTr7ATI4cLmmmIh/K192L/9zjDBE3DxCBImjyiiCvsO13+
7kLCnvE+qtK8quMXHj+3XFqXtJ7EROYe49pbToKTKHf1Q+YRDDF5cpKmtQ2KG61z
kcoDd5nn63/fjBH2HnKpqxNsFMGLmhdd2Yn6BbtXJfy+ARvUUsuUmEzDB77iTICZ
j38Nqo6W/pYvA0VwP8Y+tjQR0oIsha/RIhkE+t+SmYTdlisdYtGoUiPhfUGjL2mQ
EFHKwFjhMr9jjb/XWUlHwuanSCrn/XjdnmlvMUDheLEQGY5+QNa2PYCgLKeqfk7n
qCJD0QcZ0s6lWiSnD8vSeKL0YCeqQL1qDzGCYkVeJYlr8dJBjLDrscnB0iDyzB1y
xOKUnE+w09S8iyFk/YiYt5R9iI0Lzf1K6rByh7vD8Y9+iRB+IG8wsJ5kjCaqe+j8
vWsf9HlPPgIq9MJRI8/kPTUMGvkrNKKATT+Z7qqLGf7d2tC+44tAsNKcRPms/uqP
EZHNlvlgdGuyqYgmNm4sTG734XQhD2TPZslNx3ZvWHj0q9b/ZHBb8EYMl/XrIpIf
9SXd5ltt1eiNrCTKaD0IpEOAgG+kGKZrRNvT1vDCyWpSoyvoB1jY/N6SD4cEhhe+
6gblRB1QOUeH8SzGRTWyR7JlSzxSiSgTZVibtAtTw5EY7h/mQOS4ljW8JlYbbQTl
fjw7wZIZY4C0z3yelCBToIU9xIoi9WqfOuh4BD/ySGNRr5l8TgyCsnr4O/qB8G2r
J9C+hNkbuMgx6SUnlO8LWlJNxXyyicopGIzgSvnur05qVr4lD6ie7LcGzjH6oZXg
J0LkHgFBaciYKULukA8iCGyI9vmuVLvGlo1113N6grxXR0lOUumAQi7NKxbSl+9O
47TuP1h/R0HvMywRSK0BEhznZQYWe0ibAc46UhWQygvK7woq/msd3/Eoo6QjvlGM
3837SnDydGWZEHxMEBbrbxm62OCfG5pserLxzQiHSEbfXyOPf6ZzjFx2LjMosOVE
8Qqq2x2yYc1BullbPX7d288ruWyG/5UcI8W7PXtiS6/d3SK/bkDCSRA3KDE9pIU7
lMfZ4ZvP7Qq0+PwnICLtzx23ObspEOdWuI9xPGjxwlojfPBprAU0f3KuA+wKm++u
EG9PWaT3T83/Fhix9Hq3xTwZM9AR1dGhBXUtzY8xhqRVw2fEmUS+fOCgXjAMpZPz
tLjuSEYCvC3xIdNdCSRz+WWTMJYM3AOOEu3fhTbE0bwH7B5/4oPDWapfWffDhISL
alyYwiPDhVKgKZmoN9or1CFiaMYJd3uY28yy9hIExc4G9B6ug+3Am3llWIYVuicp
lM8fJbuSukV5UN1BKZIZvjQxBwbI4t5tC9Q5HWzeUcl9bUt+lSNIZ33YKOnxq10V
ZmdPH2BYQff6wZg+f8fGDFQ0Y4V82opehmhmycw9YpMMOV9BuABm6aJ4I5EkP7Rq
3/cxDxuR9ErkTdQQ4USEs3OZbN2jNqEAdE59GTQNjXA8u2goxvyShC4Ct5d7rOLq
WeyCwXYxqQ/aMLbuj4OKp/H1KZZ3bO2nBPbEwPB9pgrCOX+8+qiRi2e0OSN3CN8w
SmHqttHZvDjDfIpT7H5HCYrzN+mMCBO0S3m37U+qIuVKVkj3umsgN/eQ7Zd9V6eT
JaWoDrPvnJeP7/IrMgVOdJKcZN6WGhG/1BNwtY9bVaV5ZKO7DA6FTujAAx8Q06Ax
NoEPqBFU/2VvcSxC/YD3q5Fdc4wwKF3posS5EpfYB+Qttdjpy31ZWYw1ZL//6nkg
CZh3f8oM3XQoquWa2NVCYYWpo6BHFsA+LdxbWjA+0pe38d/f1PHLPI7qt2BH56cO
j80jPhJAsPBkWnUMFlkCm5Qjzy/QDeW2diHNkWbA77lNqPH6S1ze1KFKFwBrBLHt
ZUoa2FWJdnTffCI+269mIlLQdMEcobEPWFFOkZ4YcOI+sfjt01MululFxT9Ehk8V
NvIeawryVpIfTaacXUAZFcPXKyQ2C8PRZQ43al8H829ROJdUqobzuBh+u6CoU2h9
qVmM2wx4PR8HZSGw0eNUcvxnpvth/uKNqHT5ZhGl4Zrr5VY4lw/QbwYW7yi4sYuo
cKE49q70qAZOOLHxORH8Oz/tDCy7kHy0oUahQshiLsaNnNEs0Gy2Th62p5JXxaHP
XB5n1XB3cnfs6YtOzDc7l9kJ882/TeTPWBN9dCEmWo2BBnKrY+9eVO/qIDGd2u+q
wgRd1drW+19dHRHvPLBAvO4QHSnRfbjjdAOLHxciRrq4/AViWNjpVWyUSZsqSpa9
pwsz1sdHbQcjAW3gIBCv9/C+06PPM+XCx1WcvtZXXweN6Y7KUY4EBxblWh9mtWps
oH8AQF/g0hsW3zFOxOBf5FC02x8ZQETQ6QAMOPz6qb5LP0y+gqCjvsrUW556IvRR
lpZympo7aFvJqbcrVOYRosAJpNEuBvPP7axeEDaKG1KYHPKmEfNXaiPYncGSJLTr
yLuN8FzjrlR/r3ZDvvoRz1wKRItlAH2J8tsCYe+/v2uRWNPFLWMcckYS7kMVszz0
ovVvFMWml6s/Qh+X9dZR4RpM0Uz7FOutN7qej3VumNDB9QMw5/hlC2RuofhLKp6I
YeXg9f5ine1FllsbjUbXr5MVvL8gaSRxQ4brHCI7JwXNbf9jvP7+gjGx2BS5uib6
Mntq2rRbV+yaF612YOdCEPVLnlVzpYOmcQxGuiwF6kV7TAtfTZ6QnoItsRUcTfIe
R1sVYs7hZi7D8OY/WAZQM4dIOmAJSrGV2Ceqlpk1tRJY02aKz4yTb+0VmrlGbJT7
kXdUw8a+QsOgVdC1TLHqNxgg7GpgNb1jl7uusWuhFQwWPT7p31sKPI0LR9zupH0h
G0zumTRWznqTUkODAiV6tNhIJktivGR5+JzZWi0QuA5wxLM6jw9wcUrQzCpJTXaQ
pTcWE/1YQ3AAqhJxjAbrRMMs/mrydUszm9kbvBwhBbsI4BbxCrJzDYg7ZBHYdJpo
Jcgx7BtvUvgVDHq7UAMv5dmSUHe1o7m+7KX6aRsxf95TunryvKLPcXrCRT5V4t5x
9zgtOaxIYsLsBpWyAH/B2qe8yQWScTX+41dW4Z2Ci83Zrwf/8fyOQVNgxqiv/oEy
uV35Ls3QIM0f7s7ccHFHYYeRHiBWvp0go6sEtHv5Z1qZL8Qk4z8/B2647aOpap1o
Rv+JAr6fvLnijH+GwrleA20SV/3ywWcJ2E2r+AYP1v8FZYQFnwrsMdxVxGGmrbxL
DgJIy+JcgSYheaRmCY203+gqd3320orzReuhUFHhLSDHSQRVuNnRxHH1iwYvbw6A
G+9227eN5vMyVd9ddXQWankMlRjNxTcbucEsL2WezxE5hxg19kCFAFGy2FKDyLFT
ZHaV7OUzrek68g3NqipVZuTqM9MNWgzIL7LqPzj6GU9shOU41Fi8QYS1q/6XmJ0K
rJ7bBWvBjmpI3sEgfRgwzLv3AqZUy3TXupb2dcdmBQNL3PQiziXodh6H4IsV06Wt
ODmbr26RGZ3qmLjZMkfcngeeg05zUmHQjEEqFzLuDJ5yOs5rZ71GzP2bbKryT7IO
ESUFOgKj70IJCOHlt1PJu7jnGVSTpmuyEm8u9CZqM5PpFXLUUrnn5HF8mpdE2E3L
s6NpOTCO4SUQ2tRb6if31910BVIoudfJin0bQnwmxjd/1wL2u8tsMXvdqjfaYhh/
ABsmYLB89e9g5A+1G9kuWXlmLiRGFsSAPpsfmriwy+tBe1sKGztnhAFwMEKk+DFR
+dfkNDh4hpQb9h1+xsjAwbxt6DhjMhYZJZKS2TzPRvrGMCHyfooWvMRIX3qvr53G
iVWTaLvX4w4ZEV7ZNqZGAbXnLHPFY4+CdLi2Ff4vdHanOgNeNFE9H3rrY9rVwirq
yoZQ5tclvahqAW5VxUqc24KamREQHqvgjxzizQ/2M9YmqbzIglSPsT7BV63N+7mg
1h9PTzu3zl1zBKmCCIKdFqXZtHZLVzryWd54Gp8CpOKjcn5M1VynPaqKAe9+V9ao
whq+PCtfaCG9T/kUzVqz5IJQ6+xRK33QqNEZVISnesIyCWUoBI7j6RA57QLcszfQ
Mfe8P+bjTmQ8lfLTIVuRVnW++Ww890OFdQvquBbSeEkG/7KaIQMv7nPJrYfPc+We
N+dM7B1b+FMf92iYFUigEmCEeqm2FiXDXZCbbSTfCceJZB/tu9xIvROY4QGRzl1T
PvsW3Tty1RCAnz2weUW3oHNYkYN5A0te7pbiXhiVU1GRb4xSV8tFiA3mZ/25zJXR
M25aUV7YnFlOlAOjsJtZSqmLK/L8tfEfhnJudrmkZsUZhdM2+yRSNOFJl8RSZhYC
f+G8vxsZb6U02cToTW6riJcjpc7MqML5PKtt1//xbXEJzijutFMwHNWlG3858q3d
ljwS2jwxGmMIENyCb5US8lla+QJ+XhbRXme8EsnNvCa6TkkJ1XL1ApEeNJV0w3wK
YAIcSlj7+e6+GYVxapRowRZQd8Pa/0THnzpdDFXqY6XWK7Z20IUgLx+s2X/A7dOk
yT78PY3zM4ftXw6vgrdkjCEd3rpP35ZT8IHMNO87rcpX+Hx/fUiwNiV7XPBgHjC3
ZOZKRG1MWD0v5r3IRPpuGo5yfIZJmdyKY9pC8IsjGZz1I8uVEWD+y/ku7bRqmq2T
25dOEGlYEM3/GUTMPOWL7/k4+G/nGNKYcpdhgjQzlJirWUmdQSM6fhtk5O4kjDHN
OoRjUKMo3xQHK/NRieMkQ7+4Wr0EkZ8IcL5iLVPwLqfGJBeTFOQss/4GUzwDzP1Z
zxRHojMdmT4UiuuSnGz/6boJiIa2wkVwVpOeL0Ts2pVUaM3XvoUEaMZTO04Q6bFM
N7LjAzRkH5m6gWyBFPUUpNqyNnfFEaZXuFgus+yT9P45oPZA7ei3avHc4yloNwSi
4Jabhu+LFuvillhJ+o5rQqnF3GjeoauNiKG6n01wF/iK5VUMNLpMpZEmYKAXI0CW
LuqMJbZeQpF+fLVasjZLn0nttdB6b/rI+f9muwMZ+vbgXdL2KIx0MrJidofJ42RW
dQnsfvhVqqDEXzSTqKhzxGKSGslaYl9q6ll3GMgWd0S02eg/FwA8I9Ucr4xRluJv
SbbzhQB9or0wsQ4iGUjad4kxOKGq1HRlXy9JrtWsk5Q0Z/eruuzPXtlYJxvK279X
GBQeQIxA3c/6cI5/kaMUD6Qe8xxpl9zx/q76XdbMPaD7yp0xLf2cDJ5248vfYUz3
pTFwT4gmTvFF0jZ/Hd9umkFzErOPVrgE3dUC0VTPefpG+rtHWLSqcYYbqFJzMawB
M+O5iF6kpSnWxgHI2JOF5RBp0/67kMeDLQS4b/S6a6Aw1QRCOW7YI+P0tRNWbWmL
NO+3RaGJtkhmbb6sgKwxcZKKjjkt7UDUUairgVs2ktCQ7bslkjHNTMVlit8GGwUi
ij1cH2AEfLIaqbYmOBAoF9dmK9JYI8g4xhf+AeRDoijopwMo0lbZZsTKG342lA6g
gHNyS/c3Y6yJuVU41czCnWeEqs9B4Gq0slixCzsfzsZ/uD0UvS69zN5OvDfsKnL+
yg/GTBGnWWBZfAP2ls0UFyY9+GD1OvGLvsuFswDLvk8LJBufRMhV261YgEiC0HZs
SnpaIRbaDDmJR+1WU1tIF/t98ErJ28cNGS7UPVceO1j+bqOMpgN/Q0Eed8NKfW87
ogn8kZx0KiofO2c6cJH0evzA8MH7Pm/S5unY+/YjFYh8p1uX7Ji8OFJtNoDODu01
epDjJUM98oUoREhe2rMDHIPsD4mv8/9XiYfEMT90hgNMsDqOJXUhqR8MxpJEM16C
RzDlDHtx2Sywk+y1csXCDnAtnkHNYjF9XDW1gJ1BdcjIzUJCp8sO1T0dfDC8hc43
KxkmMe7uA2LvrYkNzkg1nIBDQV6H8nzWEZBI6x1BMG5siPP+K4MKWYnkaubyFJqq
zRFZyJBXnfT8Fcx/Ufo1KJRe1bN5cQ9yAoiyO8qr/oemSkVdoIvKA0qsJH/Q/oDJ
rpYpwngJWAdMqeJyGnkzzqkq/Cp+hB31zElYzZ09vt73ZIQGFsdC0uEY8vLOaIaD
uX7kSR774TMUsmj+js/rZKE/A0piZBwsjA6jYBYDhdqhq5txAud0ENSBasvYFm2Z
vX28+ZEbTyBzj14R4Yind/RbH7Io1QZmV5fVlxUq9Zzbt6gQQJjlOiinXaiYN4R2
0glgPdQvnoxIjBdaGuGFBRDCZZcEZU5mtfo6a32i86u8IbQJ/8CMOxOjp2ZRfugV
it+p5WU+BRjOMUgkwIYCcHC6vQ6BjoQ3IWXektjI9fvlxX6JWUfvhTuBEv8sssmN
gnqqfOwhEt9LA5ecVUUGgvflU9AF/cXE29KwvoDGsiASTSCZMUwj+vvv9hlRpGVq
9GrGt+/bJgRu4lUUyDyCkV4+y8DZPA+c5vUQ+tMVDQ3IQXQs0N2N+l1pug6uOtS4
KlGb4U7E6+sSwORmNGuG34EpO047J5LTYmb4dJmDrSPsG+nVmnybKsA9jNeODRSd
sTBVwTiRBqT/5ldOSMaXXH+8A1q/SFlkXw+SMYjjPH2lxcw44lRR2d+GT9W9CqXL
AabY93j5tGbZqq7ovouu/T7pavrd/RS9SM+1vIN/U/rCtuMcpCDAsJDwJomhjfdo
N6sEw2kTblQ6KapVRQDY4pKGx3xCuqHIjsKgP9Le8+qF38tD8oLDZU/OQOqdqMTl
Gb8IYh5XExdyMJEqpXh6IhKZagYIGEsfb4ZILdDeYTzjmjVlBwrAaUxO8gKlCMXw
qp5LcI5cnowec3kthiOatb1vjnvgZNK9ck8MnuEVj4ATjXrR0kACEWDXswAFgl3s
sI7iXO1kWGoKijBBuf37fMn2zjihwVxQVr17/rXOnJSqLDKZwuFJSe3Q+i/ml3RM
+dqd60Xo6yhAOLpIRVNc7C3eKhSjiK6N7Tv3cuoRHF6joYd+UGWO/GCskZimaGNa
PVEF6CLVXMc+NNdaxViLuRuHwzgr1CB40UZ8l7VdVlMUuJAkLVuURQ+sBJqhtOug
JtZW4PJiXb6A6/LzE1vzARP560ANBu1o/TMUCSUlatnwNjDsq1AOeIKZ9m8HsmmZ
15v5ylHC21AFtCwWQ6PxNza7fivTlRt9wr8J5R12NO7cH3XHt2nmcpEeIoh3UUkL
aRI38QlLkSjBM1vu6UPvE4hPPCRfi0cXBLvyYX+4Qv6htCqI/LjcRCBK9aZ/nOMk
WdhvQFPfNJ+NfhfUu9AH1r6xe+bF4LP9hV5r8eIQWMM83BnJl5PaDtXrGNMsETiF
WqRFrfh2BL6CCD8ILvJlk8kynDQZ8M0lEEq7TYERdLaeDw7SXb3Bu1w998zz5RFP
PBD/rFSaILKRTambxzkqCQm7bBbGczbW+H14U+SqxuCIDUij0eCs0nwDBnm0vJz9
KbXNseljOhUWtStOqHJnuHyFjtaut7e5a3VRAymX5QZF5AG+785rg2f96QWO/1Tf
l3Sr5CL4E8Ig9psmLNmzKh8/cURFqSW1KWPKpW1y7dkjG8Vj5VzozXrkYDxXeYz0
b7RT7LnONQYRgDXA+dVY/GDi9DY+Tf0rYqx3bkT7rgbRnMpQ610uBnq7tqJRoQDs
mrhphq8dazDh76F3mtx2gephVZq5b2sR+wr73ATDsZ8M49sh7PjlHaUMZn4EB2JP
qiuSyy8e2wFvQw3roLYLBRhCGZ4xHzvz1WqUK7uvnsT55e6Zh8ebECWsM5+axC05
ukLRvMQno9YZoQmmXU+Cix9t2MNYA8lDvfmubJpyec+mdB6JMuXDjFU/2FcRddhC
BOP/sWZuE4e+w67P0syDBohwWjQZFGsGn8ZT3kM9UBzovPmFFvfd4bcnWRQu9gww
JjCti/vmvybHmpu4oB1No8K7RXn3JGoV+msHS66PRZfK3jv9CNEIjGhVqdgtmzo2
j9vFYYcscfWY7CHqu04D7NmhykTBHmMcqWJACvwpJVO+6CwINinE1cS8abi5txWC
8RlFVo7pVkCNgYTndiu96JQz3s5kUdbnuWvXEO3VBhLIEG8mq2eZcXJeLV3EcDoU
dYnqdsv/6UNpUQPLhOBhxNftTxuGqz64QUXMwmTIVgloRhoCR1hjGLInKBx8HvHO
mZqJUdkf/G2vcdmpD8VSRjbo++s7EecJ5+Lq5wbaCoeRGclGSzFgOMUQ/0L6NUWy
ykgowvaTzvf1QOHCVWXwBhAvKUC1v5ynI1A+LdSrkFHYnEjDH9n7ItTO6GB3uivp
Y7+KGTa2KfqHeLyicSzRv8JGVVASaS1dzpc1gygakq7BWGG9SI2/djymIwhdv7zN
76MpZlCgGXHdfKyrlxpUBArgOL79c96n4cHGRhWOcoZVm8V0HZt0nWdfNXfK7nkR
y5SAaM8QhFleq2/GTx0sN+ujZjr4MLebIvQ7b9E0TT6VcGcLXwjqxhNxE5DVgKeE
09APTQkvaGgsUVc861asce8GlApxTISeJQu5ZTe4ohkq+1nKYa6wC/xa5ypC5HvT
BlXnXEsrgAajwpuCwApKS9D2xk6xeUbhH/j6xVDtEyd6A4aGb8207XguNXQfmiyR
QnKBzTjiB51I7Wj1Eem8GwIO+/IhY5ivzMOr0iV/qDup9VAtNvzsArhNKEBe79a6
zBXt6r58lpFQGFzPoxKH9mr7I0E+RYIaTrf9IuwBmE4kA/3DewIlJPqdPkentf3W
JySAMqqRQKdi7fLyY5/B6shcs2q+Cic5omZQwLjgNt6k0+qLVcUzwowjbeaGUZoX
NPyVVE056PRlTPsq82umUXQuTiJOJQbVqGrBGiuJm8GrBiusZryYIgDBnW/qDMMa
VG35TtIW/Kcz067+b7ejJQe2P2v6g27VAMwcSmUhpKyjVXU3SdU8OuEpDt9XT3YH
Zk2+tsN5sNueYBgErJlD6DKFqbn0/yRkAeXQ7ppSY76JsZnUQp3oqmttj0Ywe5XZ
oB4iCcMLfftpvsCX4JbZk/QyHCaxBTKC6BY/SoXSyyy2H8NMZukNaYgtB0VR3Ou5
WGAZz8Z+XHLY5fnRpoLsvDJdgmB7Pum+WgW77Pu4LjNWc581a0Bfft7bdxDZ1iuy
0Nh04Dn8JihZuuO118o5mvCYi8OVjbfJi9gCUAWTiOrVe5avJKmKV14Ro3OsBjx7
jGk3lOpDlyIO1r69CHrsurPsuT5dGMMApJ9Uzoq4+Ne7LC5CjRLUj3VF8T2eI6RV
waNuj1Zhj0wk2JiWSQCO+npbMbi5ZCzP3MKjOJ7/nYbmNSjEMXsYYj5QpV9MwtL3
OPX2HO2c5kkgYbgtaEkhVy0hZIxa/LqvzXyqhVpqHWWlV1RG6f7qh0ryPKvdoRFU
E0BA3alwoJBindJnYkE0HFtNWd2uDJqrC6toEYkWUKqo+LsuGssDPjgbfVNfVftd
vkkMeXyBpLb2e4z1t/H+u7E1FIftfCnlTIy8rGfQ59ytHl0E0UKIzP8u37BpIBoT
RvjryUoykYi68M2feIIdWB/+K3924zASZWAyxX5KVdESz2AHyMaOnqTJmf5i/b8a
fh/RjNsSTOH06Xy1RgQNb0mCDfKjAX2sjqjIiH/szBRVx24Cwq87AH6kdJLVl7bg
ar8ol1AfRoxhSSF5DMbUZNRGIrlxRRg3+DmuZEz3Ec3yFGN62NOrYfpdr95GgS9F
ZSaG4UOxk2XahxeYdCvncE6SeWDOgPsRznIO0pb8PBJ1QSX5JCR/yXeETCg080Nj
gCCH9z5K/SD8oYT+Hjvp18R9YJjG7Hb6p4SEU/XDD3SZP3bkarUj3VtbduLyT+5Y
OTKlYRZzFei6X35DO9BVPzcWB29CQN3SG0f/9/4GT4aPs1H+MwdI9G7afNripLMB
gFI9S9tEdH18LiRrSJXNv56Ks4urm0KziTjH2fKy4NNF1bYzheKw6M0C1vficZ0w
LRbFuY8nFPcEHS99QX5Z0FPqXp+VlChD0YirzDPpdphKb2J95shzdGyeyCsPJ5ss
U7xiUYjtvW/2CqgFbX+OroZcBHiejE0eTUY+gfrNBlFxXCZSqKeJJPGbZ5uQRW4C
/CL6S7mob4A5HynHjWAf4ZN8f4dXjJNHhDbtD24lXYsUktCk5Kxk6ZNEirEgTVA3
gAVoT9EtHJpBLRh37p+NSO/L/Xt3zAD33+413aSXAwyXL5OIaxIy9zMrvvOmdA3Z
7vXEi/j5ArDQmZ/oKCkuNiw6tNG+mzeinwL2KhYGINbeCfChQHMLB4GnGHmzx5gS
HBiBvhCk94YuNcT3VlnrrDTaYafMy55dCD49u4s/CgFI8zBgriw05dDSWUVc9zDs
R0cZMkT9onTTqPjslnwfIWrhUk7bymHUNuWFcjBOFnHyp+urSZx9EABet9X+D7wQ
nqzYguokpbCUj0yX5P4RrAztM0js/YY5nCOe6i7lTKAUNiAVT4sE6Y1E6ynp8rDM
ic3wrwqA1I11n/rYulXr/9pqZ7JTIoxkOZw1cuO6XYRxh7aWig5WRLJchhlprrNP
YyRaeqwhdOeIsAZ0ME+YOmfhxxOZLlVgVuaSDVOkA+e0r9+MXb7wOahZuSOESDIa
QcImRAkespfUnpduWGVAbQZ7q/Bn61bhchcY1XM51YrjMzQYx8UY3NRKdtSoMYdj
6dmJmIGSNz9r7IpPj/GFrVGx0351GkKkXLGJ6N9SX+r7JxQcI8BsVO7p0YR/7nWx
TTmRrXgHTOidEJT90AkeBHyXJ9iXO5P7dfOwaGaUCZhUkWyJc3UgyM1LxbKUIny1
ELMH6R19OzuYoIxW6T5pGKSdrdBFJuTpZUaRj4zktR7uW7O8JeyVyb9Jl0PM5bYq
GayeAkV/thaSl8YnLWtutNU7UsMjGePPaZ2H/HtFGgx2XWcTU4HEUFRtiwZ22B/O
UDniWxU3p497fxS4hkpFP/9b7Rv0GBKsknvCIfVDXH1qA4E1RJj7f2pc8LNpxCym
C4nJ/Wp2SNcWynHgtmYlxeQBqupCntv8rxHLBO4zp7RoAqLGk8tX29LSWbZwNbik
KXtE7IVgmjJEqAWMB/syPAIomWrvouVzrAoWckhZ6Nizj+e7MsSgedosmmUwUn3H
v9NTAMfpx4YfzmQbWQCR4cnm41TL1lsaFEgFcighlhDa8Sep+N2wNI9dfc6W+cIP
NlLWpzQ05OY7zpXV4AgPkdrkxebSrUJYbj3R6ChNE6JLHdXiIhxPln7fnJqglSk0
zNeVqAXfdRon0JYAWJjM6ubKByM0le133KuIfwKoXkOAdXgnpHlhNo9JrCKfpqS5
avo5QRdIrIKVqocjyTdWUIwdermX5FkgTZsRWJxG5/qmMXEZvpUaBZobqpaL/xMf
4DXyH1+WE5eiaDTYqrZKEZRqYnKJzFw9bpe7z1CepYU54amMr1m07IqglFRjiHu5
gYBGyWOt9tqF+BKsPlJ6ZD8sBfsMaO91Eo7hl6B2Qff7keA16Xoqq04oOqfp4NdW
AZp19svrZ2Ywkt66riNZTngnDEga7ACwuBcARKZQFKsAhPE5BMHeWA0LvIzgZjLZ
13x4jMXNlmzP8yW+1BbJ1kTd3/SDJupk26EfbpHrriEFYofMoQov5c2+Ni4qADfr
CKGFa3u/hwUFLGLBU/abD5ZVEJtp+AzI1VQ/IBTT0ImZjEv7K1fHnb9+mh63hXqT
ng+yyKcCyUedn+kgbU45AithzM/jE3WxhNgFmO6o/5lYR4XKVo4l09URvZZyHXeh
WTu7b41J1Po+TCfAapBGDLbdgSvKIolJEZaquW3//i+yLDp+mGr7JkRE4L5qvWNO
7v6jInz3oE+T20ubxRIbIrvSmNSbnKinehDoqIGJ5yt+PiEYvh4a0NGcDlDSQPxL
Qu2JyhAq4IfpQNjo/KJkGr2DdfTCk28NxiLy7s3bHV9HFWsNnU+o3VgFKS99Act7
KhON6/hmk/uIvahpiMVAQRJANtM1NDn2BTG6jUhN+2hawkNAwVpaedvTd8zUVi7P
YIPsMAXezVjY8CSiTpLvfD4yBE+hbhtjnMkso+8u0Z9B3PmXwwua/HlhyKdiBKYE
qNoxilFQGfyIXTgeOuCYTj1FhD68rwZuSD815IXtSprb1O/LW8R5Mno4Leh8RkAZ
7TVPMpGexXZ8GvwiBLXlUpEkvfBjrotloEHjPT/hBCJn4mbhKgLXeM5IDToPNwIw
G8GPlIu8+DyJQ3CnFEFxShIIpIk4/oFqspXCLrU0yG7S1j8LKbyJbp9uaIDYGjgO
7ASAh4Qh4j3zxXdqOEl3sQsaVHLYCPb1BZj9BxF3+6R7S4zVIaEJ4zAMLvWB6QvN
bH3OUNgAfznoYBhzYCY60JR8swyJ32aqS0/k2waT85/YazBMQx5KA0s3OhxqCqgN
aJTr9zy01eTwQixWaw1KDO49sisdAavKexXVDlHoId8nznup+paL7rhDuSP2k7U6
tikZac4SF3abSXHpIbDs+nW+rqjDDjIQpadDBhtLfE8YCDaTgohjv25TOcp5BnIb
uHStBjd7zdu0PUVwrN3iuSRMuZBz/PZRSxta/E1zdYKi52xkEQCQPpw/KNWsjIMb
lrxFq3IQA0EK0GXn6ty1RHlV3NE8TcwoTLERN7Vdat/Ydz3F1E92siZjd8K8gw4t
eulMG9V2Y8mGU9i5aaYE/0Zh/pS6hecXtEdm1RsEnODmMO1dsygNFy3kyF7Vmd5i
Es6AZxgD1JJ99aNWTDdQTimsRWjLXSmAl1PBjboQQLRdyn4DOug19Mgy0cq7IZjc
CCwJlb4dHySEGfNAIl+a+92Qs1u9UYUFEPaetzel98Dg5F0a37oNrdqduFNRZ+La
MHiOFEBmG1DsgBZXFSdgorqksYvJLD7HgpMqvC6f6j0DyiM86IuddfYSJdXiwNmv
zvOTn95YM06Gy325NmVbzM395s4RxkGpCmkXJ7ZkTZDsj8IHK6xP2ayE+pXiCu4s
M7/6oofiMErRWvb2YLifMVPGyCCj3+44dNe/pYWfzRYCNnIqYBWE/4WHCTZGB+ku
DsqIi17w/R2x6XWnbRyaZVIBF9PFu0OCxcw2dtWEvKsjuZutxt/LETRU+sfLHq3A
PAfrWO4M05DX99T2fzc7SKH2CxoFPNYQhDnETyMIouLB7iwUNQFErwHG6e1nk5RW
lTyzll66mVBz7obyUiFVdj+fOiB0FRfyJTVxKZmhjcONAwN5+aL0a91YOpr9A8WD
oVE7i0vg6/hSApT2+g2QNAZspKaK77XIbPgMn9pdGgiZAs2wsOhEBlp5PxzuTJ00
itLIIG1tLLbnO3Q7DXLlaWUu7DoQpkPDkIMpOr3Fz4F59Qg9yB6U4qd979dW78MX
5odZ+ay8rTNDDN9b2LWEVej9NRN8oWc0676oS9Vm6zh2Dx8RUGlrYda9rbg/RHzd
z04IrHO/KmDJw3fO6xzfSD7WrgHTxVcu6u+oviLPBy7qQbVyuGSrA8n98x/mSl83
4O6W7nNL5StFjOJYvrbyKYCI2R67mP6KVpjlxCboN6VGWfyVkiocEFcGXYi2PqGV
d70tGBKko/NlZ4DIH0lLQ/pskr/SqaKHIAC4pH5ErEEEIIsZCWGZUoqkhB69xVVk
2FfUFrXi6yP/G8flvNNKjekEI85xJKnPqcdAKfWi5ait/95PhGqkTBmKdt4yjsnG
fn9nw6KnxFcwQf/ywZ3higF3tjAacB2zsITTEvFDrTGXg0Lc/kaAiXw16j4Ga7FU
CiFmrpOl3OqC6Ea4QPb2+KTC0V9oGudiysV2suh94n6NsJMcWKGa3MFh/5Zy0RXG
qeTNi72R5hVxEwn8sFi/yGe3/cKAn0zUJzVROBtxrqSkP7cdaM/3vjMgFRqJ5QRI
cXMSa9+DKSXC5IiidpXZIh6z7N8L+c8CSr7dcl0yNcT0isYyuwS+vp2fOJKon7Hl
uMze2dh8fsamdfBC+NejFTXRXj7yIgFiRFywuxKypW4mCuToun0tLdLMISuF07nv
gmSfBmpQOhj7kW6pFri3PBbsEXWMdXaQXX3C4pMbpaF2vuzjBObMXVkD3av6WNNd
r6GKQRN6IiF03dpgym2KH310ImPDfIIQ+PI3lJzQqUc82iXqhDbgaDvLYq0yifPP
kYq2HQKOsooj4oa4qm43Fw==
`protect END_PROTECTED
