`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqwwxSM7SJZXcMJ9yaAwOWUGzpoXIL45cZqP+Vb41e5z+xDsUnj2ZC3roX6IwugG
bAk6M/inRvVynHnUAMEVmRpjhX/ZDbaiCR8Zcq/jS4TT9f7Kk1j/Mcj+UV04Uc7H
HrTAhkMPgWQ8p0U31mvdaRtzUS/Yv2F+1bKWr0gIkS6dYlkCY9ndKn5W6ihabh2Y
aWwBIOzSEFzBzHa/iQS9QfObbZ+hlC3g39j3h60J4At0hW8QrXBaRGE9ninccSWS
Z7Xml6Pupj9OkH40Aw2Qq6vyCxaH1WmZbya6bOWV+pogTocu3dWEpVlJlWE4IugV
qyPK+FBNhDklWunfSV+nwfK4s4ThWLuHXBhYZI7hYIOp5Y1L05+n4N5YPQw/g3iD
PL8sDBFWRdj8n8xZVfQW4EYWiSjwa3wPYuXW7GSrANBm1o3sNN7SOGn2BIDF3fFp
CdgDPPZ5Y9jAqtxtpVPaqfCjI6bi9L7tWb4JiP5At0XyuVApmbo2rGSenN5QLI4+
KBbf3kNgDMomX7nLrafPnqNHv5RiaYFYppe5uIXLrDqV9lfTJ93e/tCkba57DpjK
YGqYlMLgChSqoAkVkpUZAynm+xeXMqN3XXMezGzhnrfLiKC39cQyFMUpvoF30cFJ
eINT77wXA19sHJpYdyxHhwsH25npkqWFJZAgoKGsHUqKXQI+4nA7cCpUvwC8gtSF
opYB6VzKbGLnQreFDfp9RqZ1wbocbBEf/v+KgRFW6eftYnCucfi0ncZgtm+85N8W
vZ3HOPKQBv10diTrOOf8EhWGSyAM2tpsqJhKWdO8dwbauwfRO6DGDXuoXs734syT
lj/x9PKgar/Uc8v8bpjIRf5eOlnh5WLIvmcg70RBZGneIhOCSKJQqZQLUymgGGTB
9sK/ofeXTycf5UqQdDfJPOkfGLMPsjPUXfZQQlUuFgCGS8eBJL+DjyuYgbqKRT2w
p+HnADS4oR/YOlttinLcuy7pvlR4DVhS2cDILd48IfXEkDOJ72MUufpTnKLeQvqM
WobhhDI0nlu0lXzI63YEgeQqm490IhpEyWwNbX3N8kQQkE8bVnb5xE4RPgn5K3fe
FRwZEFZ8Jlsr3vP/XPiuhSJnO6dBKkoRfQOTHCbCkEk1ZPsfFYeTO02S7r4t778n
dcIrEq27ff2HQzeNz2wSO2rE2W6rZ1fTI1cHBEfwSYtVu7OlEGJhA85XkYL7clK2
lKShlnCKD51Zs9T7hXnuFw6dOlvS7on6acpv0og+dtc8v7JRToDV7U12dq0rHO54
1oIiAa5Yl7oEdcZ+3mvZ46/WAb6OXuSZ2BGskG4Wl6sxvVLNFa4ynp+ZAqGFz337
PizNZ3e4sI6eApNeU7WJbH2FEQpftNuuIOxGPO34ktSpZz9SJ6UA6C1cfuH3JIdx
/fN7ziK6sA5tBMhWkWLOr7gY3tJ9Xsu06JdtlYaA/yFdfup7DOuBfCqXiMZIjSXJ
ukWqwdSrUz/8ngtkfo209SJrYEFZZHptYELmcHSnS2UyiAZSaEt9JTVfJr9nm0tB
tyT1VvuM9PyvhT2Im+OUr+8wYbw2vZj703BQPae11VnvpPTt1ecBQTj0QBoyAwv6
WdwNNd6zSFRuBbSleBcCUfHKwsSS67Gzdrg89d5w/3Z+VolrO1hA60A5AZ4TeXvW
jxFrbBnTPja1QuGF9FtkGBcaMM8oZ5hHXYYd6qW2C4DNgX6g0mbZW0RJYWyBo0/f
zgQlVWNrConsRHNI9SYFTQ==
`protect END_PROTECTED
