`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogOQWrcuXk0oHTRr4HukXJ0/HPnHyN/R92B79WapDZgMqBsdsOvxdlDTsYJFcTpI
CHvosxE1wiZai+TOpZ+y+YiAl2CxhrtCurMibeXddLg2wj5N+LnZm2SDHqV3Z6ob
wx77AfJJ9DxvZCk/n4clXPvTVVd9pNb3idKtB/ZVoMShQPqOzFgxs3uVSf3LFjYl
7EpqjiQChsSq4++Obu4vsRF7CnAKm3jMQokLEWnuENCcZsZ8MUjukUAFb3E94/dA
aswE1mnFE+fMLpYPC438inEC1Le3t2gR15tmtahwJOR2nZwdk5IN97sdWvplrzIg
+HwX/U9yQ62ZknCWploPSeLZGhydCsU1VgKLHjZZaERJ5R7Fb+jX4JsMdBmqlcDV
sbMciJTRL41flqTsvHxRm58xWzHJ7OcltRgWqNsH8UQGZCd+6ehxjgnaHx6S4y5t
PoBm4QCWTzoHWxuw4caD6MGVvIxKiMMeTL7p+lPyOp6vbKySbztYLkrMtSyZNUbw
H1OmB9YEYsxeyatr9Z5AG6XF+4ITQ2CILR0I/K0QH0D3gPrdex76gIu0EzesUKf+
PUH54qi6z9u0cuoMPJF8k58p0z+oozySkzRHKDMKOe9NlqPYsxjZv2POnrGFGBPz
Frd5ET48j89N4ZqEfKpOxIhYpb+pMWo75nN4m/68co8=
`protect END_PROTECTED
