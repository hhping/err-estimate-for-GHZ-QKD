`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39XZVLnBOKHI4cwm2eDXTjZkevGaitIr1vJ4LrMvWzd9Ohg5b4SYycjqKTk9IUGc
kcyq5/4rpvdwpBqyQ1sZmePIfopnTOUIZtlRz5NuGn5NIcJ6jiehDYehFpc3WV6W
khlS8TcJgjs3f2zEVFijyvwECXPJrMkpP3U3S2PfNwIfYm00gz8HXsfWwzQwGh58
EXJ1eD2KW3hkPR4rzRgFhZEJW2YodOPASkxwUYa1GqDtzNHtHL5UAHSKytuXRtAn
BxPaEhI+Q6zb8GsIQ3G0ilQCgoHW20osMadDWHMEOM9YDYx1z1zSB0n8ECIwBypy
ELTn+QzoG6qstj7CstoIzJHPEo95uSKJgFI4LZRLlr/L+saBeCKM57/hFHjp5pVh
v0HefRls6ExKKktmn7XYrxCtyohSkhdkp3zhheKyWksewL0U0BcBnTXx6dE896js
qWM7iyxzURQ2sVN8UDNZnK3/osDbFpCT0GlWT643JX3GTC2xt+2QQj6JAJ3S+tx/
sJd7P5imHvUH/3p/Kl4mUf719iIrI/B7wkCUZV2Ppev+lT/pCOf1RkKy3bzST+Yo
AjpzISnBZ/Ofg7oB+4OyVFpltffcZALb4z6S5XH04WRNwkhZAvepeXRKygxOq4Wl
O+QDSGpUZedowYz4hAHfGLBVVGqYdeZX9ShbigXxpi5laAUj+yC+l8TOJ5JP2az8
+oViUh1lT8rFhnkniB85wUFRoq+1tpGEeclRmvzK3sBAzBnRHuSoQawsw2shGw3x
KYqmYwmLqV082+LLuvFDaw8WW8UwF7bSVPImXN7LbD0OUaze8etgBMF+tfGRboa9
2q5txpoMMYh/CwT995I7MH7tSRfmd3InKM3cbDu+La8TfNG7JG74hyeyAEqJ7Hvq
Gzi8mN8r2MuxjU7HnSrxUmsQwsigJgRlEgWVNkRTQTHv5yU1cDB/FecgH849IzKD
ZIFqbtmVDB8ObNSFe5LXdNstVu/kspWfuhh9yiQi9mi9N7uzIuLOAiWdsBpFXSok
MVri6OD1KD13y3hu5zMMD0OpJu0hAOypVjigaWOQczBDgALMTJC/6Oo5AGhx9fve
PwOjiK/ec5lu3H1sFzYKEudnI/dzoUA8huiyufthTQfrgLWc7pwmLOLNfO6zb/xx
s5Wc7nofYvAF8ZIIOKIRrOeudwFXDTq3IETDzPp1LTVFlghpzpn3y3yr7G8+S5kM
bdzqCsh4lO9pDbCm0Zfms3ThIhZHDraCG0Czpeu20/xyRGAjptf9Anp9bLrQEiBV
MhOWzAG6uVCIfOjh5DxA8o2yyYzibUtgQKs3Bpy2A54K4tRbFfKxq/ZC9Jn7567O
PiYGo2f9baB3VVdBgyA4nXdoA+GfU4i7BsMUo8oSvg8vmGAQJpYR2jKRCoos9hfx
VwJvxJf1vBP/TfJKkxA58rGroQUb31rojr9qOpxfaMUlnz7Bro4cM/5ywUXlBkhR
1vpGoiLFqxkCZ69rEJ2E/E3HsMDqVRpDCPs9g4xd2XbSft2fQi6bQ1ReQAUS8ogP
bagBVUvQJFQGt4j3CNbgn+uCAuzelOJK2kturWhv9vkCppzM+mcjT4p8IACWGOvD
sJgzOF892IO9yf/MzrpcAYyBx5hR12HAp7bP1JdZq8k6UoBJhMHZDN1IHJiolILK
Ai+dLRQisIPv1GIma7Sj+Pw8LrI+EG3bUXdw2PU1i/g5viDh1hQTkIaeZ960n+82
FKi75nc228OFlOgNW0EwMpBaE3E1UY89AuapCri44D/KhJbo8QSv0hVhyf8V17Zw
rmlk2T/c1vgP8zXINoBmCpO0kSh0EbmulJO1zsHLGLurnSoqkiFE9sGkLeAn4TsP
mxAB8whb4oHTpkFT52RwsrdlB+jppHekbMFl+oD7u/KbXczyQvfftd1zz73CEUZ8
`protect END_PROTECTED
