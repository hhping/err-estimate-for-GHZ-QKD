`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1ub0/+gWn+HhcOnZx2zACvYPpyVQux8sYii6ZtnhxB5+8JakkoXXm4gnIcoIcCH
WBXnVeD/hbnjTEFw+1H0jqlZRVlBskdtQF5p+fzFT8pVYQAPWwbMlZuk835d79ub
48baiGMkEmZjxT8HuItn7sREUuXQtz9kcHXUsFqgxkPBZE7ngCDa6Hkl4x7xFcwQ
iNDaNycQ4Ib16paoWIB5GY4vCO0jxMTAHBgr0U2TMx8q/0LQDj8/P+46Otj5BM2G
r6VRzySNMSMpu/jEJdjK9n7+H3r2510lObv7xv16fwCrLYAuH08p4Gjd9irYqOne
/dwmiO+Es5Zz0HxjytfAj5UShhHHjO3ncYYXpGUiJH6jNpJUXn9KxKlb2ezTpCbL
WMGJlP+gEiSkLtKJj4Umq3nWwFBvmMFh0Gz6n4OogJnhbn8GMy7g0WhaKpW1Al64
vlt2VAu5x9zEkgh9EC9+r2DYB0iNQ55DbKwpCxGaihRe+2qQHO7e9gkQXgN7L0G1
uHQk0FLJnpztiWXdb7fLBkPb06z/20NW/C1jB0r68/7d4pCcBmciQQ8+1luFqwje
ovrv92WE6sXeny+F5AWJXbn7NNNEo0PpBlpaJCLcKIP//NUGeOrTOXD9IwdHGJyb
wBKwXj5XtP8eIEr9CqBnetrsK6xBTdOgFxuS5I/jpJxoNCx9Pv4d3tSTN/4PcQig
2J3qCjlrXTvlVqvs5uXIKjRVpfoMtAZeGV+7/4ADRLlt7voMS88+5uPmWh21Uz7h
ID7jAsbO2KZk83PJ0clPsgA7wFxkXcKxp442BNAC8kZ0DTsdl0qmSPEdXCo5EeiH
Zk5pmdntDR/vMGngDAnZ3wgB3cHngEGOBMt24kZDuEHdXhTXw2nhxbqeDVLPH2kU
ekrS5YgcQXw/RZebAhIWdJsNGpIlKQhQYqdAskyJHEU=
`protect END_PROTECTED
