`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTaSGJfHsquS9ADzqBZ/lxzHRVgnK4VuDFK3EtKrfm/JNOYNha+sq1Tuh5tcSOxB
FKhWP67pMgC9pSIexjKTzu+a94fDsDAvpHGP0ATBIvlAGrfdonGuc2TkrZs2LnWI
Xd+31W6Kd8g2d5ffnII49JB8rQKUFwl4cwG5ahXXeW2gljXU5DJoZoPZLk2EuCbv
Rby/0ckCKjrEiJcoaOUwo1CGkYO5PLX0VKM+DpSJCrOHIV/D3l4MnEQcjTLJzXnT
dVVbx/c59tltEWl37ymabH4TY+ftXeWlBbA+lk0lipeNsVVaW4f6CAYc+ZpH4PkY
NsX07CkiiamI/WFoLnKTzih/dKRz+vfmthRk66Rzq8OGSHV6ZdaqF5N5vE+eM5wS
PRt16CNnLsfH99cpNh4ZWW/P/s13lULfjUbVbWQDgl0LLMD+aa0F/q7VApjgk+IP
e5NTvsFRUSTWR1udyHA/OHJSmvu07Z1zb8PnaURx3HEND5a1Cs2ivQ8R6t5rq2qv
yO+vHB6oNvE4/fX19Zh5HjWgQmDiHJbAFJuuCzAdB2KUJI+806+kXaK0J3+DQvRz
TQuwlHg2m6BeigMHy+W24D/RvK0zVBTZY1cr9Ci1zOzDiFWPsWawUQEtffoA0Zlc
TJ9bu8y8PMHTm2Yxeq8POBZxJxsEOjzF21c3UX9K5JNLHn0YyIBHKU21m0t6URxV
fjuqMUxrT8HaefAC2b9KulREKZlxa+4HIUDX10yMwQIHAQbvhVvVf7+E38ZGDUT0
Ckg5xAiSNVcSoyXxkUBpSMUdbUHXYpPxJYO+Otc36TlbsucOD8TlR8pe8ep89kzf
rmouRU4SVY0VreUheKI3zSABCyoG2ED4OpriwoWCKu2bz01WgrnjbtJEijs9vl3b
lQ1WEu8gu4R+V3A8WsqgHKUKZzDOCFDMh39waDauT2lCgOb45QR4RnaV0HWeJMVv
cMeTO9XgC/Z47D8r7oGxVXQcE0V29B5RFv4edb07FN++jPScpYf/8DEyfIXpp55s
5lN8X+yHSWPuGOwORD07Zb76qBODK6bsP+uKmFd1W0HhsQ+4+Ic33AuSakvS5tiG
i8Ms93j0ENse1AmYGiUAMKKlnI87g4vecFrv6O5RpDdmK+DPm8e/6xconRCAYpmu
WfDqOl3v30PLRboJ5U4N8841Xapzbjkdsazb/ZyfZXaSTuDtrOVxK8kjaOeZlizq
utqIshR5KXydZ7KdmKbCngD4qi6//7VKYCrEDLxAld0gnKhIfOfU+zl5QhmKpqYm
EyHSSDDkHh6S9SxibOqswGVaoDyQRBO5GmBTzWZZd2iyJAr98P4uRf7qcZTAjyRi
8kjyIsftEZyhh0lq4CaLd6cFw8gegXXt01cGEKxn2dgCyyDPu60E0MUrEXHQkMyz
zN9ixhUsN1cglXHcwebLF2m1IeAzlv+zB//wZsHBv9jGioffwAEO69DkTFqbKmCe
F0Se36zcUPqWOd3F3BgSMA876B1WHFlP7Ea7iza30wfGo2C0r69vhdkdNABp4ZtY
DVAGBgzg79T6gqo091/FWc3Hr4Gqc+0zzbxIathBZGhoo8mwpzN5vieXM89huvMW
mOZ2ZoJe3JFFaQQX1s6MPsD81Gm1zeV1U0DMeJxhVscd1Mfejue0va7TNQrnNCpx
SKyKONJ91hy9NmzU8r+HzYxIghIrJVELim+4/Gi7QxGHFKDHLUWjO5U6VzPEnkU0
U8LAR1yxb1/N8x2oyx3xlx3Bx+cotfbhOmAkmy2TrCVPEcb4docE7dA3i9Prcwm1
Exro5+ieHBDWGd/fYmsULl0KeoH68VTJIq5fzxF6v+Y=
`protect END_PROTECTED
