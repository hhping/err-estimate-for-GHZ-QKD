`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eob//D2ygvvlJGNios+OTHSCmDqW6x/T1PqHdpkFH6oWBIiV6ytTKWQbuQJaFmBS
EkV6QpN+/ra+j8wBJ1oKY3AT7QIYloCyJ90/7t+D4Hs3h+J/qfmnkcAcN3aA9pZa
uEXtB/m1KDd2O52CTJktOcxOqa3MfNRQKgYbEh4tRiHr9s0YdJoy3QgmftEDy7Ns
f6oDcx2Vc9+bhefm8uavCfDYM00SlWQ0GUb66z8qvugiCpZauMwsFzhmgxHbptJV
Ly0XVAEETNwFdbSiJFbAlK2XEuXlxkzmI1JzhQButHEACHT0fVq9qvD5YSEoSjxd
DMF1raYb/n7KEZJ96wtijLvmABPlJ3ajEzVqVFHoznTNO4w+thNnfXQKXtPZGGQI
Cdr737EJwwUHj9mwbrXPO/VuXcAFMvDugo790MFWWAl6GDcZ7V2aQ75DoqQvJt+h
HukYxVwJETAHsbk3wGrIA/TleL8FL8q34epjaCNu0cGIsD87Z4Nusb/1axYZm7Sm
1kQZTPtOoZREPTDm0XsywpfSXVunOqQimC66v9PiAlykFj2R4gc+YR2kGT8k1E4D
5SvZEpvxprUalGJV9Ic1DXit2zDu3KNAsPXtGUKBTqLlE1t6EQ6O5VlSQ8sj3aa5
VDfICjvGxtHxmZlYUQfWjEJucwTZv9V9we1q/96YWqiAv2w2/qvSoZcxKR/LyWcR
QpYpowWmjq5HzWMIiVg4ufXPhUyggeFay8tx0tDnfD325+qV1hZ+p4cYfacENlx2
3yb5wNcuUj8xhVONXVszhPIoGRfY03pJRNkoG/5AKm1lOboQs2Ad4xkohe70snoC
tmZHaweG+HHgeQigXD+0Xn+yDl81/PuvKOAetY6il70zYiHorV94rDAtnWVTqRtg
HloiYvnw/3b+27ZCpy88M51XhwDnTUK76hISMrNTzd6Ghq2MMlq6I872Rx55KP1i
89U5T3e8/bXod/YAI3qm8Pfo7cWEa92G8uzQWmHeDMXad217el6YNvioq2yKE6Ym
mKigdQFPmJ219RQBcnEcuBYVnyikDYYhOnbabLxPJ6GLkRDr+Io9+annb6rUEnyV
zND3OCPI+HxKu/fAdUi9bbZ7wmpwQ7+4Uz8WA04UAVOJDMZcMY1uwPPUrOU80fZw
4vvZJfUV/yI46QQBnGqnxFsBIbWJuXMaMrr2PrzJ6VZ8T4HPvOl472NylNKMNSaJ
KiRtWGXvgMpOmtDBmw3c08Qs0Yu05scIsYDQjAdJTR2W/SJw53+39Y7TqiPfXxX+
ZzuGQSgCuBTx/4IMmeRfgNIxBk84TBgqw8m8GA4Nbgpx00phGGxsftet/kL5svCi
0E0fbwNNlxBrkKQ1pRksFYcfeR2c0QUkHno31D5pIXuhj/WHqvcCA54NEoUDN2nD
aNdscNRYAHtw5Hqt+PCkf2aHPNTiY2B2DLOjrqUar5hscQ906KDr3SwXoHtEt+DL
a5KVTCQan0jaDyXbZIuRoQApXui8ROoMfPmYLZ8MoKpAKY3zCm4vVn8rs2c8s4L0
HIkDRHv3ZvfxlgRKo930epQo3jum6nHeSH4/AmzinXhbDlssrtw75t/ea9Wkpz8g
hvJSNVY50JT9RARh0IWhXAwKP3ssRA8vIiRzWnYqDyIIBkhFysmxSDUCr/h1pgXq
RRLQSyu7zAJPwOLLM492AX8vIxVVX4lZezz2XmXV1wY9ozyjeXYp3s77PoGnmLfp
nJZAAlBYrHzXPaWikcbZsGorYMH8dDk/qOBU6/OI9p+3QWJ5pWi/TNts7JrLwd3m
AznlD+VEkhtMp7hsSPsjsqJyOS/pbesUiP3eYjpnnTP332jqjPKcy5f2AiC+Fc5x
c4J9ipB0wWNIpwxZ5rsSmvRS+S2XztraOktavLeJ5awo77ADLRwuogR/oBWjLa9D
jXq1aVFjwnY7ZBaK7lvoH+O8K0eWGnIP3a8/3rcUBNwz3gcztKNuBHhcyCLKd3GZ
64/huTldjwwWa3OEzS2zxdwbIfOeB5u+iZFXyUKYMCVfUFST5pm2eaybppi/olSy
jpvG/hxEBuLHl/NxnjHbRj5pLUnb+5/jUBtW1ETSHW6dsmbuVrX2IvcPbmW9ptZ9
z/fWXqCwhULVmGKJnYfAjkxZs3hsnersSX08Xd4xZFs6T9DQVwMwSBKJRFZnO5Xe
2WUNXUcy5i7bzFVAwtPdnYInTwkfpZPaZT3A543Ek3A+5KchVFFg2hNaleMV2yrC
Bx8tE57uI9RLFLhjAPS36pFahCOnFHZwrvIuJmEL8K7igaXgGRlpEgiA0kx2XLtm
t40Dvfn+zIuhjQgJRLYxpMq2Qv1ozkBIuhjxdJ70HKcDgsQ29A0dGLyAHQ19RYM2
7jZwye8mNRL+lIeOpTfEHmBGAplea4eH6sguH4n98lnJ3egR+Z+9sylybv1d3aVI
5CqOqteeZ4zqRcFCl8VGOKQHtGgf7KdtkWkfzUSBFPdLGSQm/Fi07IhtnIhmpvb9
Rg7W2joZALIVzkytUaEfjxVmmusIqseCTr3tClBaO54LhpkcvGv/1fWsdg/eoHnf
2s7y5CbXz7ahBJTGkM7qTCvfB+p14Yf2OLZd662895B9oxD48ecjGG1zONZnCxd/
rj1KEuUL8/hXxKhMmg+COE/0+MxdvVlem0CvrOHBCFrtcdVQq2M8gueKIWUUeCiP
kDnGDGYUXRgSzA34GtqsdrFV7Oj1beRfGzN0j9xFVFGvrPmUyrb4/v5V2NzVzYrh
hoCTXbW0UpSs9pAND3KyTD8mJ5AgPWv137e4uc6N3Rk3GLfTo65STzIuvev46Dby
k0vC23zTs6QXWoAJgsWmuuDVKJqYeu/O1RZKwp86jKl9XxpYUDELB2Gmz2iHmyzH
l/2pjxkzyP84okmgSzQUng/YIreeBeNIZBgrfw/Pbvb+n8Wznp04Bct89gwfBEhg
udGIAjbAdrWGgrpLJGQTM75sTKY6xP/3FyWGlXLdUaNEPbHWIX3Qz1rVslWhMcq/
sDMMPx3Usc6uoYnhh5mm8B2gQ9SlBfx5QVKwiLYaMx+i0Wnt8SFeBJ+QHUuW62lr
VtnDmRKgyUP4PnFNLU+dzchif4VJiu8AI63sAJLaXfmbk7xNH0gsR7Dag3dsWlYR
UyhHzL+CcJc76ph769X8u8LksdHsH3rH+4medVYrIbRW0johBp20tD4Hgpf5DJPj
qxZUZbXnAS+euybd9v9D2xisvJobI62/gbWg4CfXXlrMLmo6YOGH1/i6uqdqrxgn
mUULaaTaBbXf5s63FL10dFYolUBouy5Nzf14RZVisY8BZwn1C1jpLKrDi5+CNqtb
0PHogkiP57gDGnsv3Nn8lMkVoTAg+4KSOctiScRqiAyJ+U9b5qaukI3KfjWd4nng
CCRcUEW16lyi/UhnJKz1zdBcxy0bhpV4QBjE4PzJs9/vddy1/wuXUc6tyZhIWglV
DemL3+fvO80FSHn76rY0+ashIvNpVqNnEDJdDQZ9QL5CGMj/k24SZcjEGjPAw7UU
kmF4SCzVCFsgJuVuQrWONOjyT8yL6Xv3eeZWsfmMPpTO5lvPIBq8RjlGX77dv9wq
ku5nqt5S1CXG1mWHbhZXuKoGdA6btWmYF0EcL1bOWiXjw0kUGn03hjHqCawZfLGp
PzqZWSKaAyhg4mO4Py9/70hyRLNTrhyroemo9L5o4NnObSLAPw86qQ9dWzOlmAvh
9bf3ewOGI6quCbMKeb6sgGcuF9zvuympm1ycBG3CbY1j9eA0ScHiDl1JNMUpu5fN
Z9Xg4eGGotCihrNJg18aux8sF1zTUW19PFImESoXJxV7RwVjrb1SHhgkWbQwHH7s
`protect END_PROTECTED
