`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0omyMLankmHO6fY+ftRd6i4WSeK5+swFAsv1oZx0W6MdP2U8JNXHFMvfihX2Rin
wj4e2+9sBqM2aASQsf8xC68zvR38SpoiSyN83S7qIs5Oco3mXY1RUzoWH2tDtn2P
IbAvrhviF2FWKIOs3jOVKDwfjWBc6FTSz3ipa6d66W/5z9RbHqti+MMJCMJ6r15T
hYqtAc3VShtVXCkfM1Ste6zf4BcFmvh17jRqCOY4aPMjC3LDIS7CGcYuekOTx7Rm
Wcm9Hthx8vxBibpd8BuWj27QNwMxl3dHLV9T/qFVAhiuLVSNCZKjG/521+A3t3A7
p95pFb2LLD5+6z9ZTrXUC5u6HRVu5Npx0ulivgi4mbTZZaeeDZ8qK2mw7FMIqbLx
9dP85t2bt4Rw8poEI8F2KOGxUO+yP5MAa+/+CxHBV2cTJllT82S5lBPY78Xmt23Y
Uf4mIoS+6M/M6oy95p7Wm/PJbW9phMNKSqyXuRfEJfpHJpeXIBfRGQqypENt57NR
gzq7Wl9xaJhEJAe9QMipGvgPcKoh1zBalDHy4LLpxW+Tfr+h8Y3CC5P44hHgvv8/
BmF/+uHF3OlLt7fjJTDyMo2l9Y0rXvf5ZcRdEo5sHa6d3if4m+VGGJI2599zD5zc
L7VwNIy5QDeMhHxpaFMTi+pW6rRYh7vm9jBqHAQGHQSP9bUJuKLZmUjvekUL/PUa
LjUzaGph8T2zaj/W2oyRFxBaEX1WpfiqEEdGg4aQjeFrQkKtp42j4MX9/YxwdPMk
L8OktCw4cIpK7O41Q2PN2U17oDc4dPuHlz5pX3TMhYTgsyOcSKhW+fmrdcL0YdVu
Xwpkk8k3aRBK95vVw8FYSXfLvgNtNHNP9quiXjt9HVFhhxS7OGxyEu81aDwD1ze1
wwKlez7BLqtzPE4h1IGrIxWqj4Awg3Mb8P/IzjkEA0aCRPBet66EcB5ZMvZx53mP
1uMgYKcadqey/4SOed2uKEqymkpNz8AnXZmVXwQMqMWByKReqGzzl3ro3gKqTCJs
TyTVo+sBmfLcVMq0bJbdyZNqWlZhk0wTmBup1PmRh4Wwzn5svFLtkgJeB3oBjoTj
tqzhk65/dCt81+GOHoMjVfzzwaji2X4pRS4SPB2A9PW19H7lzVlVKbnPxyDMDXgY
yyY9GR85VNqHmUxavQyNuGNGUVpl0GY71+ljTTpmwkVqQz19F6adsk/oNJqbOLtA
9HlVsMf5Fb6Ze7TDDO29o8eEW0yMx7HusNesrXhpGwaKjcV+lCxLReEk4tNf0syC
K6aFR2Ig+rRteqCzSX3ua2lC+Kyxsj/M28S1YsaZSAK0wGu/vKhWK+mIFvhiwTkB
7JoSOmuN70kX9c2lTvU28ZPi5lEPTTnCMVPAXBZzTpldGkVh1iJWf2EbfuWdEQeS
ikdz06zMeaKOMM91pxfynPJf60DySDyjCsXOxhQI/VZx1jxifFdz70EJrhMS43zb
kJ576ZWayE5QO+MDZ5YJAskc2ILafyVkk0RWa5HjoG1p3OYpcy/yMqFKaiMrCOr4
MSPt1Tsd+t7nKH4bc27EbREKd1qS4vSj3OcJWk2POZuXGk1Jzl9SppowuKD5EocW
Ba6N01/KMa+N0fZAExYbGCtJN8ufU48VN+0hn38PH+4OZp3No8VHDc4gGy++4e/6
DAgEs5IfoF5VCk6p7X6sBSMqPS5LOxPdQ0JdzxYOLarb6yw4yOAAV02GuVXAcjPK
2itKhlhEblDdGky/6A2RBmtRKCG2qYmKUCFt14RVEK5Gn7m4lAIw8++0Gw0jQJaR
VRAiiGLt/iVPGSMokKpJnsr/VaWY0i9rVIYGgMdsD9iMHfc0b2cGc79kyD54kg8l
SN/h90+PREmJn96IyDJZFob3oEvmkpweBTj5mULdqHVjk2nAa/PgC783MD0PLJzW
z1ZOQQy0Fjk7jIKTv7DsXNmKAAJWOVr9PJveOQSJpnMcyxCZYpt9i9iUH81Yn3pU
TbuoY2P0RYR3DZLOWVrzJM/cEES8SgImZIKDXPA6WV5DdBAtWEF1AUX2eYCfluhM
NDM9nx1lnnuu/aVWlDeI3C94/+yTumEsAJ03hi9pviVN6M6n/QmZ1TrxAomyu9ks
FR40WiIDx7JCd0T4MPgtOq9Nw5jMA8yVnXbJRecnch+34Wl4mS9ZhjX/BF2aGjye
vMhPE2M0m3eS6sg8dtC+uLRP8WNOp6MVeMy9sHYI2S2OHPXtDJ3OdIrNU/5+RYZI
FptI0FPtMyfDrI1zGD/SnUgvwVliI6On1bRrk3n1xwBiKUgVB5y1S8k9ZSPXe9kf
M12zIN9CwUyC7kbrOu7wz2iHKtA3gOq68xsdgDQsBW3Ez5cDvPVRX/kX8XML0ESa
3duwjCwx5mzzmFLY8UxBr6lNZUnYJcYCFLrnEEeMmT6HB1hpE8S10eMbFL7my6t/
Mb+pr6jUA3p1Jrl+iJ82q6CsDaxIGfaFIz0uOPcAAgmUwc0MJ3eLmntAxQ2ECEbQ
0lW+kr063h9P8ElB1YuTPgO6lnNY6GeSiojahusyJUHHhtQzx7/CXVEDaT6tmYTP
Fvy7jTjTfYuT0g7+tghn9taEI6O9CQPeYsunW43OTLU6YsYcVgQdllkAckN0TV4n
Xs6tpMr6Gc9/yFbXp3+5k1RLBOHSUbYOvbKdR53rtxYV8G4x7RvYn5bPxQNZ5w9O
P/Xyo3iUsIYOazFmzPcD69j0RftyAgaj2wWlpD5mj+CMtIQPmi3hT4ZBgluv5UpZ
/7WNIC0hrzNpK68wV6jC9lyYgsCw6tfco19EegyNJliuUPa5/e3a3bHQ9AQClzNB
z4l1kOgettnhpu8RNTB3b+F3s5rfJRpC786xBzKypWKp07h4d5/Z15jnByzl/k7r
ixg9/MrVrT3OuePZ+PM/pPShKV4QwobLbpPxibgj/1cG+83PECzUgFUP3YD9MqB4
HcQ/5FO04ArWFyk9XS3nvYT8JRhEbkaMuwi0OW8R/p1CyEh5u1vP7gvDfiuvvQWr
UrkI0ylBL11rSSUyyc6aIITzBi6fn62P1LLKV1o2D4CXIFnCq9uIrre/eeW3m5MQ
IuOm0zBiTFabZRZczbeVHLlxhbCjoIcZfxl2JIVp+N+GLGndATQQJ6OeiIRFuKp6
/8H3UZnx9UdaGrtob5MOCdktLjs0Hk3oUdPd6WGFf7vONF4cCUzgnJZx0XQ5fRDL
2ueR9CSvQDfgIRChhI8nnVqvLbUIc34D8NJ5QuVlXosalP8vszYOCMRV3RIFKfab
xDGDCTQK3D2JXBxCZ+9pm/u5Mb5iCPcdGm/XlmGWeQ/FEqBYKUOodrbnVeJPOHo1
c266m3+LXOsxaClTLpBHoMLXiPtz9Yu3mIFMPt83dLPwnnictIHnANPPxIXc5zJ+
S4UoeOu8oacM+7TLd4Of2ZjLY1WvaEuPDck3ojOYe+W0bHqxy9RtJem6ydnUQ8Ip
aZI+4ZDYXGq4TAdFOmbBFQD3n5N/bh+YiufLSjxDME7RRxKtnoXFxOc7N2h/KB24
72bruGTxY+Gt2abfWsfP5qtGsc3Rux9KCavIZF+6FumgSOd065x8Dzw02c0S7fSp
NEkiKlFEIcGQ7JWWyeQ+IBNd3u+iXfU2QBR9jtL9iR50d/WQIXY6yIdN0rcAwhh+
INrxD55MYU4RR7DXe7LZNUqhPpLGDXlQ91CYn/KWMQ1EQuc9Q9Ja6iqotoq2w6OW
ijbMHRnkppoGoaE2QDGTuCnEkMsmJl+uZx042Wk5Sb7p4F5XTUio/juZ/HiO/rGF
nUere0M26LWdVW82yjCASEGup2nHGoEtW00MWmvanb5HpbyOLxxlUUAj/mmmtfva
SONkB1UXNL91IsFjSleW9p8ElHxKHSIu+9vStF1qv6rVPhwK7qSkT8c2Ydtn07nZ
qkYVswikZcxlYUEmz8gRwwGCR89ciBmShFQtrOqrrq3/vZy/Lp6QbnsjqRzWrcWM
VKbH8nRtOiblIF9igdg9/ApWM339reJB5K4Kk1ILaTGDtT9kyBt0ELIjuWvb9WN5
FJwfCidfxRcReu6Xy83bNNLD0ETMU0eWAfRTfClGar6deyMJ9yuodyqYEDP1E/M2
PBjaSvu26AB5I32piLVLNKnJ4qnrusLJ75ggSln0tYpSAKOVcL2ZvzvT0JsytMFc
BYGYlvfUI+rCZn8OnT5m5w3xrjr4aPGKzeH57H8dDYtmfsNpV3iTFw43704GmV1v
Ri7h2nsxYM+ejfWwFtoHmQP1A5PRox2DsiCIveP6zUPDIRJCYt8qL7MZ180QqBwW
saElI6wBvX3TFvd+k/R8e7qH11nTQ1Mdcd6PohVUJCfF3qairNygFJ/LsvV3SGrt
NQa6ZoJDIcqDUQi6e6AowWNEWfpDYgDYb3I5QDLz8sLXkuK/fFcZJrpuFVYMo3yI
RHUKb5COzoX6ByFQa+w+456gYvMRjhZaJ/8KMjcwlHhBVuN0LmSNLIG0l+pHw7Xd
O0UUT4GTbq6CXgkKcMyNI4bYARr66EcwPuZRjW5WhZKl6ZczacQ5S2bkalfEvM3v
jos2TYuN5bDva+U+p38codMBeU5YSm/Wsp5bRW2+Tm/45KCPVvLpBc6zNXmS1g6s
bhv+aq9hkrfzczoIgXc8cwj2qsTpLXCxr5CjrE5NWFz4Tsv8u6JacnEFSdPUKyRa
8GnumEynG7Y9BjUJ7ERVcdqxhh6VdYs9BAP2+KPaDwxEUTss7y/ZH339MtfrEgFG
CBKO+gs8TrFz/KiCBqhe4U01UM32JBorQij8mzr3C1naexCdioV2biTvG8HPGoLV
umC36ki4qE7uyqnAgVPyl57u0e+oXilKHSpV0XI9mzbyQvV9X8RdFyuYci41I2D+
SCrCC7arjFIeeZw8yTo7NialdGkx/ysqicAl55wkss69nSIMjx4zyuLwWrn45rJS
CvSUlCKDH2FqOdVCzwEHSxJCwDmwFxaV8zfop8a6w3aY3dXmUArB0gcMfSWjNrDD
YbP+ME6edsw2/3qAzX+ks6JE2+Fzo9Czaw0H7AwR9725ikDsJzkDh7f5EFXUG40e
WkfZ8oAFpMEGUot2Wvja00vGVHHr2Mi7e2o7NmOsXszvqqZIhH2aILhWOCZ2oooi
dZ2ssc4E3xsTkk03a6DfbSNPv3ocFL2AyA6kqL4AQTKXOfZbcvVMKkKPVMb73CAD
3OZL10DjXguPmm7d+u2jryMckYajEWPTvGT6+B0qeIZZUcE1BuT13L193AaFcvLl
7aA4DMEqg2+7P4ENYl5etTm2Z5aqpCNOP/kUsEcpDxE82/YRlEg/NH/aKcltE+2R
EqX7JPFMcpDNkuGnkmIF5C6XyDff+BxMaGofGBF69k/Vb3z6RBFpmaWXwEcEJrIW
AmBMLHe37qKP4LWfp0tjdf19SGfvCByzdqWPa3EO4sC6q8V4P2Q1gOKW4IniCW7n
Bbj3AhIW3DL2VAYbHsWd1mGFPuRtuNA/rmSjGBq+DTeg/eaKl3ssIcdcny+uH8Pg
iNsrhNIo4eZ7Er/ZmiwNNIx8+445mu4UTthOUXH7V4ZYoyF35808LVl8i5LkkFKD
NYjRydo/f81NvDsMC7mkvipyZfiUggCAXWhT8+fOgXavR0oM0iN6qb5vGy/POY5y
A4WP3DYxLKa/SHZdx/4TCbvZGg+TEAB++783LUlE0Cd0MbHaw6j6YEAK0zTR/fGK
4V+7NPnAazKOJh7qhJ86eQ2zTY4d+w3kqG/kRaV8g4Z0S3CVm1nzu/4XRi0XQ584
QnWLTTOsmYU0vuC5IJYxw1f/BpjHyVci3ut9+h0PCcrJTU9UGi2rTOQKg2QFnU7b
hwRXNwbWldGnNJ2bw0at/Zegti4f5VyjPckZNnFdZfQc5SyEe7j1KMjE7N+teQ66
gN2JioXgva+ae8UW6pnC8Ax96TeF+MHDuF38gumTrUSUdrAs6znEaT7f8S08n8GY
4j5wDRFvHBYgSEO7QsgKc/n/LJ8rTQIFw8WqcIK5gp674GQKOfvXnxtN2wVcbEPd
h683rm5ug9hi/1AwLoFzR7X5E6G+zbZfi3JEiQJqPU0FX/0Zsw2bgK9iWpVB/yll
0UzDa/y6aGsaGhvwdPT2F2hNOGcQrTEbP48ml4Lvk1jdXv9xO38Ioc5YAIOv3VJE
kZsYtA4jfZYpRPRYm8KrZDSDuH53RtPA3b/6k9q0yeWlIwGHZQub5UCq8kmwtlk7
CHh7sxytHERCJH1Kc+f2g0Vadg5mumD29AyFUNT/fU1YxA4x7kpsfIFqK5QD4NUR
JjU1KzZyadAR/J85rX5qBFkhd2ze7syUkDchKW6fl0HvS0Kbw5D+Zv6n5OcYZfHO
pCTkWVBZ2xWA36awC1qMiz1NC5K7ZY5tk7RrM29JagJiyIRSlcETNBTU6dbWVl5S
cg9HZn2WdWOmfBv7Mz4bBFHmL7mkDKu8SdURXx8IBzP7yZBIustDbocPXw9L1N81
PPwFeTr75k74skwTUpZHVkhnN2wL8Z3QlSIYhBeHhR5i40eOj6Kg3o7wPZqwGWqz
PpyjH07eJV6s1uJPkXObqraNoG7ml2K6U+rjMK5qkaVimzSVRoSAAG7y22Eu8PWo
qmckg9bgb5ztopvz51QExq4kwQ6hzA/AvmZW5ma+3gLoiM3FtNM4jKx5yLmMixt7
tRQxbEpO3YXpwjynL4qUlU547q57N4lMZWFKZvxUSj2qThdyq+TZUwmiVWmQHBHc
xKNFIk9F4y//ZFr8w0zowLvcXxVN2R0pL1cxyiMWytJTOH8Cir1ksPTS64wvi4QS
QbFcvq6nSM0EiYNy6MU9eI0+s53CUVdVOdwoc2w+7j1UtU7EiiTC0qDfh2Psv42/
rfTgb921zdRf2zlI+tQ+6TXH4h5gFTxsFzVvfvpdH9Xa71kVBewbEXQXzbrsczNY
bSob5wpW6SUca5LnNdEJ2TTBBNI7iX22m2Nehi3f7nketQEx7+8d/tAJmdFMf2CV
xzPWVXU7oIb3sHwY2fjr12+KFtmzxCflKHnFQucxFnSdaIOUfUAgHMnSMf5VhmBY
laSNSCqjKzmoShPdRtBgD45g5dqrXSrbnrPLsMKyp89wS0c8y7zzM68hsAFmBPmk
HgBE8nzzaQfdwB/RE2l6994HHDeN98laf7P/VT+sF+fe6WuQo78ZuPvgoGIFvwDS
9K3/7xGW4s/NHNySuOrx7wogL7g1pTkvEZ5tbydhN1rUCDXevo/FAQg3wjEL63Va
JI6VKAbo9v4OnfWPQadsY23zeGpfEmAG2n3R+EdBSEGmFclVgf42Rdg1VW9P4V8Y
ljqOkTTRxfgA+gktYvZgf33yt0DpsWHxnUdZ3wpTg3Up1i8H5WOmkZ/LC4whlSx2
5WLD1jtLhhoJvO60Q6pfr6+pESBhPRZzoRUJrGMsN/qdwgLHhTNbeSMQJdx9wF0g
SykcO5NoFt8PfMTq9/AFLnUNhBLK8dIrDJMiuzdkuNSs1LkcSg2SUoIw2k4ff+t9
pVkDtvDZc/whcbADo1k8JhPvtqmpuZrcpMa+sbB9TerDKooghdq7H4M7uYu5vV/s
e52yrlhff5i9V2w+GCgy/gIZ8cOO2r6o+0pyc2HALq/UMD/jysU1G8G+I7rcnAvw
PDBWXyPbggw5IYvwEf4PywGYO9bBqB54i2w9bykVxwWT2MhyqlMk3FbA4veG+BAE
91JKHInUFF4RgK6amKBs9280KIExN+oLWGsVAE7G1dvdNjSI6BvA0ng+Jy+JjnQH
n/iZLaRqvz6ysYAdNuZv+waOOfda0++3ziZA9+5x0C+DL4eA1vAIhTc6utCo8qi5
0i90gTnMXcJyB5m9A0wTwDoOThY3tIMAdJRnG6H6XAWZVETpPJXqBGQURUl1y6Nl
i8tt+dD940e9cjHAOMoIT9HfrykCspPzg6/zXVHKMWsPAedchS4Wf3EggyVaA5ZG
6hgeI/JfYeD93si262mlalBGvkKlrtSLGxpyMiPGRvBqjhlPUpfqA+ZZ2yO6/2Vu
JK+gt05qnEONw1Pn1qxJcsYgMBJZZ8+jkSMFpWDw9MKw+4xiReJdF7vzS9jcZMOX
3GCKpmQ5tBUrPd5tr7b28MpbUkMgnLArBF/QBP7zhyBp1jaqwVa/g8e9VqTbZ9hK
Gy2h75Fd2Hhz8DLY4gENx/VRj3pvyyuh4iO2U96vvwjT6tHiLrhbhUaz+7XGAa/z
HYoBDZOdrP+jo18RIBmp4wCKeA5Wmuqcf6NE79Ed6+JSvj2eZ5TaYGgZxbW+X1CJ
B1FaKCFGafLZKYF3q8qojsefL5BUwqqULLAuPE+/QYcHB/NT3bz6aA+RjT+yNE9B
tgrLoGfqg26mTynTDlD+xEU6M1GwEpfjJGM6IqCHkyqEVcqLervovzXEPqPusNf6
8qAjX13XtUWO7ZqtMJu+t5WL472BSjODbqSwRUvevftSE3FnELRm8DbbcXyN8Hn9
SSBSviLwPnz71ppGN8eoz1WiQukrOiL+21O+J56kpTTpMEg1Dyv3LqIgpXO8qOiQ
Uao8FqDdvbIDgMwokRmWTCVIK7x4+nDtUauKCTVpysVGMSh9I7sG3QWVlcTpEayU
Zaj13kExsNiozpG8xqtJzDeoMwakAZJJPWm+VWE8skAvr9tiDfT+qJtaV6QE9M0C
GXnkDTqGjRns05K7OGaZWW9fjzF1IqA+alrrHKhMnFoMzVWt4g3+Zp01SMVNIDmw
/EI3hrHUf2j3TwBZOGs6PDHgb9OFXSmiB/yne+ddH/1BAE2CvYeUZsLNZERA3rlw
RlvQsg5ovAopPkI1Jd/udEV9h8bd6MBsjNITclB8gIHmZmk0ODs6wCL1ZOqWnn63
i0XBNi2x8MXiqI0c+r/dyTVrgh9+VjA2s7mb71jjM2wW8on1jJoCU1mHoptb3/qf
4OAbxudSjzVoE1jcb8KLsxX3T0V8Lc2eS4QOEUTelCtxrIO93AVOgCn0B6xhZcEu
gioMSn2DCJe44vPtR2B4S92FNovjCuFkBr6vq4wr4/3hUteGtVJg8uSubWKrADwK
2pa/J3I5/QswV+72p2JdZ5ieXwlvUFvyb6tamJ0U2tcqj0Frord7F/N6khyu+nqb
QG+8/J7fAKTdA1l9la/lYQsaojOJOjtOjcX9mjSqhgG8MfiTHvx1Tw5+aBRpJe5B
3rCxH1kc5Vz60G6ZiDUC8leNmgrZ6jebt5z1B6fK4MMk9HC8yN8PdLklXM+NfdQE
P7hvfv0nh7Fl9mylQtKGXyITMBg6MPmKP5yZZ85XUxmZEB0hOIPg7EBmE7G3VMBp
SnNnjgQORYsQq2REhWBAc5ECVAmEHxqy9RfLjUhP5aAJizs7gPWjQ5rhLV+MoPCG
WRuXudpyB6Pe5t8lUsejAb7qV/KuYn3I+iq3Es4Y+MiotNswFVNU37dqxUyreOQ6
F8ZqKzMXgSmhCFbXsSjHcj658vvtj2LmI9zDBzCBm4pPNajUIPg8IzYKq93r2mTV
md5DZucNjOMzw8yXyBqJXPPiOH0zwQ/XOxstDzPt6Izigd0o9uMbPhdvDGmyJWhB
+ZWNCJ//rdwcQq9DV2o6fTFuyheRn1Qe7jhm7wkZRloQQpTo2X1jjuNx9JAwfI9+
fFCkOdie/S0exI7EgFeaNPTg2dfhpUEm3qTSsujKiJvfplBBNtDmKyTveMUe2bFU
uhEZQCwTIOs15/eaKqxJGBxeNB94s7SAI7mfpITpUQXCjdmyZ1ZeMCj7kjR1Wpmo
z3CEsZ9Hcx8G6LfCdtrZmFplsd7celAYF0jHMt3GFun4xWeCPelKtYjqR4/3HlyA
anj+rUYmcrN9U7pFIMaYXfbvgi/SCeM2khW3fILtPhrj6DVpto/uYKGPBDsMu/dN
xratW9qKEyjikgkoujPvxiboKvDXnaW8NyuawIhEtsYxKVd4uNfDJ3rlDhxXvZl0
Hqb0nwdBT5JwpN1fPCpGfVPTGnJ147f/6XJyD5eU9earyM6VDLBmt4OxN4PGLGx9
ffXAl9hDvBcV7VgKIfbooZn/UznnhAKE/CPDTMD8QDewtkHlEgrZTPMBT+SuoJvL
LHIKQDbNUa8VgrBjGvXJmus6AZJAEvhsIruWhHQ/Pp0NwVachdR9attF9AZklyVe
1FY5haRPuq3aNvEF9EI/39VbcNkVWFNsvI4LOpn+J04CGOMgwhhOB3iG1y/8VYun
SD7TZ8j64JxyM2SzlG6Z4g9zmtwhCktrIUK9sR66zt13hmDiSzWhF2G/bEx6xc1y
dGXuykqA9bS/kDvs2TJHaG+ueBOkCz0bpzY3m0GZLVI9JtxFTucNXPvjqd2YWgFS
D0umSn/jSYs5cEpkhJ3e0RE1Kd9lGpwp+jOzFHCuVgoLWrNwoHCJevvbnUxBQWcp
HOKFgElvToc7u4gV2CmZKVQNDFBgIXvOmogvkIkf+rK4TIqTOx+ymtlPwtSITq5t
rdQvBcx81uRqxYJySgoCuBfWfApRjBI8WI2bNGl4BVHlMTrz/CuhczCtWHC/wC7B
NiehC9FVSEjJDuWsRFGvuAAlfv7BvHbEC59qEWPGFraxLprOLHDRxzFzUCWVMkAA
viwUdnyQMxXlezB1nboGTJJPlDKuljY+PBKVTKyXp2IIT23PnX5sfPSoovYW6luY
URnjY/GwvIwayefgG0NZThR1rDo6xpj6oJdODL6p1d8uqV6fjAbx7Gt2v2+CJ9Mx
Lh/ZNVLfXr+Elb8oF+4EbvFaR+zretVkzbysUioVq9ZW08jtC2zWnjfpkldOUEhq
ddpM8yhYsSADq6fstIHaiUkl1A5JgA7Jncp11Wc+nusUyReU7BX4KBFkkxefJp/6
ZrGYn4wOwGgK93iW3O0EpUdEpe/UScVTKlqg/Jbd8fg00Shu4mXj++JePbzJ126U
vF2raC0dgW6l4DLzr1Sz1UVb1awdlie0i5lgbDbM05ab0xk0YpDtnEJNth6BWz2p
uTKTFxx3nhbSXWQ68BCrogknd+M94wX9P3MKDmQDP83hAzVL6xGJEBPxl2xTNGGc
8l+yc/m1FazyEDaP7ez5Ub+wU6LcuxFojCrqo80p5sddAnLQqq4oVBYrPCGXS2Ed
O6JgC++XbeEvbapy5c/AJPTvqK3GDtY0duIacXzeno0mCKG0YmThOwII+aBolcNc
TRFUUWLyOjZvxmweCJgXwTOxaKmOJxwZNO+FDWSDeMZ/8/yuIzqYfpQJd+uxh57G
Xb5b+tCD3vkKviwQCPjDyZTk7Kmtzy+eYpZbuqVudBp4x192OAO3p3Sam01S7LVG
OlK6OQItFec7PsmRmTnEiMKXO4il0cQkCIYYHzUVIxj2s4Unuy2w6Xeq8bcEc8X3
J+ky5PneBzCy1yWcEB5ZLcpWsci2xYcaOPWaxmrEOS/4kYDzVHfviWLUucbWLurs
3+uHLDUdytrim8VN8RR9/tD/a6VchwDVC3Y0NwcmcTmnf7/AoDRoR7fqIpTRc+Ga
lZcaZBJpmtI3/FvOdaoUatzECDMv7959BTUSh6L7L5Zf7FwhCQfBxrQSSa6xsQFr
695PDtDAFLZQCiu1pnbdaqGQrOz+vyLo92cSUuOMuwpKA9pQU1CxIzZTZHk+obpz
+ajPFMrh8pt3KkKYO46PZy6HeAUTeAriyVh2m52TTnas1CSacWMfn3ZOBWZRI3SG
4IeUHbwKQA7qWde71sWCvof8gmzbAH6sEmohWcGYb0oSuKeaDtmx3iIAWQIeA+HO
JTOhLzLY95IOvNHsiONZlAhkwPbBSXkLscVIG1Z2Js+tJ4LFPYoyRxZYRlfTGtdD
Iukm/skHGCpQNNMQQuc9QWtGGr/P7jxqhJjjbvI2He08rJn7Jg9WT06UsQLB6+44
7RrmrifwQrqOLsreBdYFVIoxVZi3rmcUGW/sd6r+8vy+iMQvfWxYiCWngSQVQoCL
TSaDBZUdJdO9CZBrw9yM+yho7NJtmniOgj3wuEnXdiqzyPxa82ErQb4mcqgjbcKI
BK9N+FkHuiYsMS6FHs2cistg6E97O/vCDy5S5LR7BuBvSiFX/hZwmXcgiTE77GSo
/lz4WG5AXVFTcPlI9AJB4GnBRe6mKZwF1kWM6IOjJkd77Py53URr2rQx6LuXEdS1
J3ZIk4nhkCDnSh8P+gjzZRAWvkALJi1sp1rmBOYcqfJ8dwpH9V+MZFxw7pxNenj7
Kx/0XwK2Ir+3ZvVw7VbW5wCKWW2z9Axrz7anK+bFVBqWPhhjHfRQOI2PvvdxuUhX
M/5a31CPVDGaEb4m9anqy+zpqAXVYXDm4jaYqvZIIjc=
`protect END_PROTECTED
