`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62mGAZn5UivvyfYHS4ouTSpB0WAi4Nf+tMoC6XTQvcDYCl5l/E5HpTZX6nGfoL1Q
/eQ66qmXvcKdOwcMPS58yybdma3L80vv5tN0xtRySrBjsz8pFe5iOPIK7MIvnE6Q
kXpWmmuHXPY6a8TAH1wLbqOnauwhcYRt+5K8pXcbjkivC6Ub7JYVcmfqEvG9LS9T
gs7MQB21IGpK3Dl+C1wczGogsAOGodC1MZpJD08zowfFQGbVKCTOGYuHRyhZdkpR
oXq12cEk3rqMNWnfITMuebQ4LcvOEGYwt7dF2YXgBTHseQfqtbGlPXC2DdoHNIqv
6g2P5V4LQ7YrY7BBtCNtrsEf8IjinziS05GrLrT8ZDrvf5O5PNIhIkdakc3Qj8Me
ID/vFrOtViPKAyYTJOQmJCKtUwdzwjr0i5gez+wckCrLx3wmT7y2WEEVsKhIVqPH
ct7PnwtM9A52lYyowyd9kdPuZhf3EhYBr1pyTaQ2hYbJFmiovp1UJ3/5IA0EzkKL
A7Xfzx79GKxxgxwKi4Imp6KaBshAuuhLRn3Zp4q2Gt7jORN/SNVpZlHJ+dE76mY0
RTO2NVQejUx7oC8Lv6to5S9Ur8IILweypHP8Y3WtHEC1crDJvnweoDaczAPy67Y/
K40+XM0JAknVQ2TmWdp5Ska6/Uy9U69vnOe4saOFkU7akoO4aPu+04Sh5eZya8tM
1h8ZkfHyYm5yRizjCkjeEqpODn0jMyJn/mMfWij7YCQA/gwr6+qhUWG2vvcKjZGh
D/URgAW/wSwO6tdGr0+yD7lAvNZfiY4iT2YoYH97wE1pD+kYWCHsn5guY9sf+y/Z
b/a76RjDSpLGTrNzSmieRGYxH93Q0DQ5sPk9kUeD8+wzVFVMvWLvSzaDxEAK6sJt
11uk6CM9ixHzXoF/J22UcOopE8E1r3L4DyFxaKRXFO8EhyhJVV+tQVu1QfydmBQB
wSGfpfLASuCpn8Mv6Z5ipzEacJvb3ifAp1OKdLVNfroeT5zvqvR2a3mwd3TaTgPU
XRU7mR2Bw3GkP0HIyfWa1NaO07nkRptRfVN1HCe1dTJ46bi++UPBvn64YNGH9W+Z
Sz8OWbYhEYILLvr4FtzWS9rCmB4xNulkm2X9S5LoXdWHIl6SU9XPKio3czMH2HrD
bjnH6WkRkialS6Y/061EZBdNk/g/Wx4WdR2DL34Ln9gqN8vtAoGtIWdIKLTpqFIp
3TTWMT7VSxCHRMqkwBqDMKFw0hwX0A1PInX+mKf9uHRBGY2+/xf49dfH6ZLm4zi1
qDFb1OYIVMrv29gmof7IaY08vJB/8lfnT6KaUvegpSQzglL7wEvQfhAuf+lpun5S
u46ComBvINOT4g558bXHiGJMe9BwfvaQYhV7HNHf3MXRWXXF7FC2Doz4dJhGO9PQ
qIt4lq23KWt9QH3xeZ2HRtkPGe4lqK6STPm6TwLpKLnyWToROpd7E3h4xF9tf3S6
UwCUA50+3yWir++c0Hx83xrwf9uv4XllgV3KDbwuN7XAF036BuLnyr8CCTOHRLXn
vCGuzViTHx7qf5tjnpxES9B0Re4i9fUrrY1Gx1mVSFBtWYO7n9kjaQ1u3PStk62o
nlHWeUECSrXcuxJmjB2EoshC9qaMTTFplotxDZciTVFrMriHcFZr6s6N/DYsYKE4
/Qjtx1EvGjpBNoVsjEvq6tHS/kf4uw6jt7wrZxtLCbrIXcxJVp0GMTV7O3eua08P
225PEFmXp2XrX/YkIHAZ4PqXaMPpRkY6+UNi+M9+bhK9RdP3XxvVA/ApHNB/A0iW
y3Q/Ztvb3MsSDr4yxk2pAJwA6NwyLI2mC8uPxBVLRc6Mrdf0MG5NwDg7AVb113iz
Q40qamqMaiNTHuieU1M8uynS0lOpycaUs7X0fbl2Svu8LrJm9jsprvQszAa4b2ww
rc34uIJ1B0HZSwxa/twNQt7M5kVu8jNm8szJyWUBSosg/jsHSjt0lrxnBv3hbXzH
Ns2kjbu+dinaWbI5z+s1iu6/qBztWZKQji4Z2TfOGJ9LzDDmAno/22XwtblRMyPV
3kxSbIyInQSvzFiQP+kIsbuv2UwJ4a0gh6joiAo/13EvEiQEISxm8rAPOB0TO+Dj
a0xN74bueYQ65abfm0wPjb/OEtasExi5fkyaekcFddGst7IyX9rqsVlnezI8a2AH
92RiPoX38nQcaUV1CRQOZ85L2V1nwcU/EU1D9I/pva0LM6Q3704OvXyVbuv7A1JG
B2g+PfTIx9xm+5lj5ysB2+3Ber6AbQYsife4iBu5iT09hI8vI9AMeeMzGtNKBsXu
kvFfTA3oS+Jna9de+LsQynzIvbfIRr357Brzw9E1adwHiUbxH1jKLsv5Kn+oXYHl
OXumAVzOpmN1K8l/zu70AKNiI5yajKlWygO0Yyoaqr/bzzHPo8xlT1w9ypG76Zp6
6o16y+SaxTp5rPmUxY3h3fe3bdEi8Q8vfS6fTZyDlsdReYnH2O+dUyBCiMpfIQu7
VX7rP3/6V54bs9yNArJ5snLK7G3/KEgv+b5wKij35c/NOZmNpt/rUxMqrVqGI909
ag08LQ08RhLC5DOkAVLuoMOV5z2kECWKyU+BptPyohyefRHM6ICAY2V9UECIsdMN
xN2BWsd8b7mmddHehMBBck5KU/Yb0E/ucUOLnKkDtpN8BsoWzja4ax/8cAHSmMFl
E5Nzv9zdPDHeOn9hnbyZG+6E5bHsQQx5QyElR88oNptGa7/mTVlcntTUMzpppmxH
t4BZcw5zam3y+UojjGU4z5UtL0xxjiqdVrN3j6Ml/hdFtsJG+Utjx4vkPp//DkeE
6K31HiVI4UiegtYuzJkrLkOcFoQwKFx7dcB9SvuWKU1nosDP+57wGzeq13W4ozP0
3P0lSmd2zeqtmf0OAwd1zo2M2jrMTQp0mLriaOjV0saXTBXCudPlQTrdPgdfG+pB
3nU+ID57LKo4E09xkkrPbmqmuYMbuYpGFmDIgUm4ZEd2WFAd7chd+xDdpZU4+FQD
kbp987ZZifq7DOjRAgW3OEioV89adLMRKpsUuUu9utqmmR9ebE4qbzzaJ3vyg5hN
7m1o7LSqPBEYZbJJQZ3TIoxwdwogt/GaSWZq72meRpgegYyUFhtAH2/0gKs4oWXZ
URhlstSjeKF6oTAuf3rhCBFRSs7howG9CN44d83ZkpgppEzYuDGRNV8wXTaerH2m
XwBSG81F7GUlihQ7jPFR2Qc9k2iL/nQ2im9fCV8TcvLo8H93Z3ovh8DQfeVcGVRv
4d5MyJOAN/a4mkTOp/WILy+IXFJ/ywr9g9jAic3hwUnZI+v4LD8xTFxCVxOlNHI/
Li3pAvMrg5U6CUJyVA3hPQoNzWQEbsLajelz2OgH9R6WzXymGMONspHYe+L4y4yV
DRvOH2YDqRQoFFEn5j7tmROtQ4kvCiu56pRBZa8ETs7NCBavEvs3qjturoE+edCk
Qnwb2LSzKuxUupw9Zvf3Pb4sAQIBx31V78JZR+d1R0E6jFTNQotUqdw+uM+bypz7
BeO3vsvBkUgpdlDahBEtJE2z8y71VK2aVZx2odllpWi8VUid5YtB66vGMGp8egN1
9Gtgvm4O3de/QeBSGTAffavJASSIc1gdBTrd4EIBp6FXyTu2niPERAbpa/i8RSDg
1u8RdX+C81Z9QFGvdVgU1MAl3WDzRiy55MBbxbD0QYA3Kb+72Y8gR1r1AWSHtlNj
yBfx2YbApZwtPKyNOvga6oSW/C8dU36S0y/WGCdE1gnO8wujBm8+q/41Uqjw6EEI
gdEIE+CTXxRkRngylaeeyklaZB/oHH84KtcDDrJ9gCgPPVwOl6iVsjtL6QkbpweU
W0uejxZZl7eF3QF9sHLOnLqc6xoAE1PkdLewKWtP6DdmilOldfddTtVxxAuPHfh4
y8/Da3+ZeZIkaXY1+oa3SJZvrgWdeXUKPPhhDmJYP8M5XZEpc1Lxl1eSIlM8MIYT
S72F7BwyuCV4BSn4+kZmjvq416U/pcYQGnKEaQbHP04IXMy2YZ7ylUz06WHfd+Tj
urcq7Xxg1u2UFEw1Ckdm3K5rVS0DLki7PgTTnFRaBVB15DapgsSAOb4RETnpgx9z
2TucjjAdaLvKXTLlzrN0bzVM6GwkVs5LUgSymqJkt9siCuP3lySt0BtVdfd67DOb
xZ7uK9rc9Bf6QF7vxXibwn5Z/lqTk6bxoGMXnnusTRCxGBGIs8Z0m8zSPvPKcszS
rELxaPIh6p1V62A9bH52YykUldD+qWaWNep+RdXuuA8ZZCqA0T/2fzybd6UEpFAw
M0gRkEZE+7ZFklJZeTe5lwXHCar3jHrCxrIF8RoeqJYZqVLfqGCEx8OJ31J2GL6e
CIwl9ddlcMICNSoREHzk5dPqf7i3jpy7JeOQ0jVpo/pULeaPUEVaLA7wiPexIFMC
d/woRt8qeCGeA9H1aXSpS6KYPJYV6W3a3t1dCcAesMxdJ3By+/zvwPUIXotMIblt
ds0beHl6iFA+lqbq+SOr671s/Q/Wkrh/l+dM2aKe18xLdAfAhKd2Ce0IY+X9DZzc
CxI0yYXm351+4RUEwiAkryfozLqMeD/Ftth2NwkpmkxSP6Ug+JhXznrYr8poOTW7
`protect END_PROTECTED
