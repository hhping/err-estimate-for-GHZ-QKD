`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOWCyBEY++DkIF/0frPTrD9HoFALyxX10EvjqJskiKyirh97pnkRsb3U71Ap20YH
FpAv2Ai0CLukGyJC3TpScdGWgtkv7JQ+CQdc6XMUauoTTQt25JaV6qC1sA5BsCA4
cqzkpe8HU+m58UI2z9F0qCQ28ANx7Gjp5wZMejpUiQi5JDq0/jtKo22EaHEltcDS
/1fqfigg3PP5Z7xJ6CKoSRjUPyXFZMzy+wmWIlfxt/v6EmgrqfjXipZg4t14EKMY
8ywLJUZhSOPEdXex9cO3WpcM1X0MTM3B8wN/OH0U2wfxsoOwPQeK4qZ36bdpz9iv
3uwhftPnOULYZSRlfsHhgbdXlM1Ez82n2zKZqL5g6VXxKAIISxltZ0EI62feoYoC
Fs3ueEWxFy3EPmtrQPJGx+9p9lLd0tpO+fMVjER/H3CYavFkFxMDjzT6S8NSqsVV
1Yo6Pjh4uIgjPzphnvbIc0/uqfNJ+OmE73g3E3BHK3MHs1XDTZkGQSEnxBOtV069
lEO3JB0X725I1PT4pRLszmyadtTleOh6y8jYNr28S2xn/ONbFcippS3r6zBW7Ui6
GWGuYJ+iNvq7lGfIf/pktx/moJUk9wGOujHJbtk74WXJFE5Y8nW8s/u1gIqf48zt
g3TbjFqm18SjWhoJZQ56QeKxTSoetSDo1tmrE2DKgbGqASleKyiTtTa+PwEPw+Io
7u4fH1Cm8r323vAD6LFPU75KjZoxQDCz2XsARf2f0McB1lAMqqGSXyutT4EYEYZi
NItgGeGBC94GsQxejfxUgnSzBkJMleujimwx+pRFp0YQ6tosvsdK/j7YRdkZiym4
hj4ywbyFTDkFAdpX69YYL3K/ZW+RCHYV8YZW4l8M97lRsjy2Y0MyOSqdkH02xqnW
5BrPO1VzNydI3w8KwDeZWn6lx8R87JbFTnM+24HhCV0k0EKdDpH9bYZ+aGFDzt0b
tL0l8imz8z2Nt2nIU4Rp1/X+4YjsSjybsEFNgev/PCgTGjkNRvsiBlGixZk4g07b
d4s0mT/n5g07xHRbtzW9AD6kgXv9DH/qY0WwrDC7ISjasGJ4ZwoKdYu2BE9H0+Az
ru1uJg7e9CEXVZopj1YzQPg8jZYX+CFOQdnAW2QxZMWZiCB9ZzHFDKg2liw3nhCf
cBY1Pg8whdSMykV5XbX0G2hE3UNUAmnF3+zQA0TzOIrBXQP8TQu7BCBqDIyQHj9Z
U/7unjWdvD24EHuNNBlWJPP7u153+22Z8pVW/Fr7f33GhUb6//Mbk4wZxxsvH3l4
bCweCZ7KK8aL78MRJvwL5u2e7DoE4GiJzNukMFVjzOxefBcUb/ftNqudKhhofXtB
lIxvyqrL9tHE8yrmmBEekCGIbngI7Gs0Pdn0oVehLZeiQdLBSuVYWPOyPL32xh1q
3A/NUMiIbwAoVNYMvYGpfeYsk7GjdUr/V5LoJzTfisOJvP5UnJCrf4iHFa+BGYuh
3RcerY7leBWzvmTDWi5gSGn+rMCGerQe5qSMYyYh/Nvkj13vm2cJVf8lAI68Zobd
n3czHJEz2L+ZSUurcVjzYxMuJZRH9udJSdCyzDwBq2go/7JgH+SFn9CoDfCQ81wJ
BtBdf6q8zjTkU9ufvH6wOJ1hIYp8/z1KBP0wxT+OfFjb3ppdrX5K6RjzaU24kToJ
71acueQa0wdcPYK0SF1lYOXOJPIKuA4QfIWTfql4LaXh+GbTYQgDCOt/tmE2W+dT
0dBCKgIQbkCtrFLzBHMgOChzKayXzFwxsvX2fqW/tF1NcAOgprHYz/QCTGft6JE5
UCXjXGIuJHAncHJ7f4ebGOBLsrMY4nQ4LwLAJBwrtmRf17TO9fqtFvXmE4HII5QM
19l+bpoFDDNAvAAwslcg2tTBDEIrT+1YWNXJ+KzP/GLPZ99b7lBiABft0zeSsrof
IFeuY6okff8iYbOpw0ONZi7OKm42feKaDN7tXv/vGbu4S6nlS0rRCyWPo33FHlnr
oQPhGGPiBfClIqBG+NM4EqXNcXDHGt5Ajxzsy5/bziR/tGCAp+wghX4QEXBEgyIW
rD6T3+pdHZkdiXkWSzcGk79Gp23MmBB0HgEvCaJnudnFQtAyJ7/whbgXHZzKkVOv
bGnnFoxU1U7EgKlbFAy68aAoM0o1CVQIxf25R2tNBib4Hc8Lftnrs7tCyhHQQ7IH
unOyFlxG+713U0dJ1jhNL5I+P1SDsJbTEb8aY4ul9Bk3i7lAYqS9qGY/t3hgoav1
l6lmKfUYBdnRCVu4FYNpJvoFGC4JmlrOiwS185Tb5S/bRjsftZJ6dCRB1sdARN7U
SJCBcWXl9BPjf0NHjW/dj03UjW8n76VZgdgjVjuVoNofFvTtu4l8ih6vqF/pXfUh
oMpLbwdez54i5Fytxwt9ZwW5Sh2LjlwhPPU9DzEBh+sLyFrOk3KpPsXEBs1lR8uV
xK5dUdvwefYBS1l59Lm7+PM81/FL4hpnD0Ph4DImOhoiRN1KDVIwTrPAmEGRQE1e
AkS6FYkCJHHtz/Ovs3915bU/qytXMGOEx5MG4IneHIuJkoVQh/p7BaBEwKg/3WSA
Rcw5s9Ev3LmjR1F9YSiBTsCwnvZeS6aa7PIXeeA0NSY3Ey6E84ejSQCS2YFAoVK1
OGOVi5YQIBZUdbEF/O5zjXYuQsxFMU6Cv/Hs7D/IUDmB6nlw4cDQZLlogMwoiDYu
7NIJSEbCOb+I3/LW7d+sfL+FSy9PTZ4G5vpsXV1thlVQ/vUpqmeStMIdR3FpmehE
hfh7reETBnM7RiLjPBq8o3vThoHm1z104nuUat0ro+N7xsoOKZwU5xEpggKBRRx0
GW1q2Jwo8+dKe02z9EpH4yf0pgYYhG4hvKdcEeumV/j/Tfpyw3Lbkmh6I78abt32
6eFeZgKQ/Di+/eQPm1OHmfwcZs873/bHXqHoy9UWSXb9DGD0agSMlP6lpD6yl3Sw
SThNtqaU2PfxkZgruGQaS7CrS5GZTjvSED8Zk78yaHDowRGJWyMvkumoo9TUh3H0
rCCG817SSfiIgKvgicryXETpru8iWuHrDIpY78K6CBthoRNx+RJcOiQV2s/Qbjs0
e5cOdEsqorb+//gbDXX75pmUlWIupfdPgCwNszKQyBKOZBUJ4QuWh9L1/SeV+9A2
s9Q/afxAQsw4vAIOSV92bfDNF6xZWbzUbySafkJAMflcsClJpzIe8a5NuKDkESAc
ZirA1CZ1vJzz9CDbvCJDvDkHeQBy9vBoJ6/wcG/vLbzswqUo6mvi6BJoHrr5E757
iR2enGpmamEoAlL5Nngjkbnnw9TFdPDW8VbIeEoz7Nl8EO1O5R5UuYcyGAfxP+16
5bDaS+UL1FVfnciW84R6YVZo8TXbbbSiL3847tD5iutvhrG/gnpCfipSwts75PxT
urFqVUOD2CK0OWE2iEytQr1hc99zUZeCwjO8ha8OSSWK74DbJgvkoZNd0xCFPaaG
rKjYcrunxnsdUduEwmMKVfR4TOXcRJ2zfzeRMPc4ewzu2v1PsiGe58WaK0H6lLWU
48E7me4tOZQT+EiQ4gJfY7lWS69I9up1tsCMSC24QaYwAV6F/4S5IyXYMn56I7fV
S9VcEvhYL76gLfIzUXN9yTos/C+ykjafhYS6Ho0NqOZ0xNCRTD22TtBsaR2hzyeb
j7OJ4IOS32OtY8IHh4CG0aTxpg2mM6EaiNEJcrWQsGXB6xTJDIDzlXg76fj8OqK8
q8DaK4hrT8UryBzX4EbSP23zpCLxEioDtgY4U+LlNXv6mWtStI4q06OgWoTdIu6d
DBaZn7i9vgaQWYGiYpRIpRPA9UHYtP0B08/KJslrRnYGzK2Tw9KGXUWnEQ3MK/q0
xkjiDrCeyQXnOtKkL9tJnghB/Ld2tsr3NgBf+Sl3OoiogxwlpvK2NR3WGyJSpwiM
gKl7uUr/ImfLSkvqT9k7mD76PvL/yOlSFk3OSMxUC8Pyd12rEfawdh8d/oOOFmca
lB+GV8mW9nctAP0c8N0h8c8rNc8XMvG1J5DLuX3YtP/CrSiZCnA2QHAB76rdGXaV
7Y44akKbDDKPjByr9HHlWp/+RIGBx7qyDYyxahSvrA8G2MiUO8xZsPmOCkZwjAHk
jFlbDFX0Z+DOrmlKFhqJ3gjGHS0heY1B5jmx1NZkNZtr51gjCBnHIFtQHRU1KmOK
Q6rgmR1CtJmEsiPVtL3KL836GP7Lgtu6FuLlPrhi52fbf9W+K3d+O0kJeM/y4Bbo
PAbVXRM0Mtfs13QD2HlD8pktbLQl2Pf3Wx1OiXQF3ssAExErh2Z0WIy3m3DVAiOh
iBxEnn6K2VEZfs3xEqwqF6NTe5D3TBTKoVwksZ+ek61Du2TP/W755FCIyI7FB0e8
ylPwauYGu3NKzaGknJUlP6XFys9i5oghSpwoY9pXXe9Q4grx3vP6ihhJa2h0nc7R
l/ZtrKxPwNirsl5HgF1i1+MVTZnDVvwitKTV86L0TUYh2NnzRiuWE4b15pTMZWuz
9YoRRqmK4h7GczdxonB6GgtxWhWyLw3UjUzlPmUX7Fvd0HCQ/DjPSanAKgT3LLn2
Ev6sBG0124UXmj/9TJNWqoyaUkBb/E+xDyyy1/D8dPBfLG6dY9PBW8MhMaQ+75EF
nOK7GvD5dVvR55FslpcH4Vn5ooz4nGlI/nxXTlTDlr2IV4BdT2NW8S7GE8lr71S0
VMw6cvG8OQUs4/gg74yDj8ccOxw7nAyulTzpuFlTU1A+Ff/w1ryGYReJWrrDb3ES
kC1DD7yy2HGKqAqAa415bsxB2BwgxRdYg73CLtu5uBbg1rdIKHErgzjLHMpNaRqk
l9Kdn0r55679icWQFDVP8X5nC5LqmYwLcsypUxhK0c4HkZd+aJQBNZ4OkUX6UxRN
zUVateDCNeG8xzL1yGO4UYUEfazUI+MexA1jylEMYjfEOB5xDWzVtlIlQcMyLU0P
7pbuQX6ZIr7SD3nd53pl3bR2zBzn+vJ3UhlGzMzuuwApVh0kYb5sqDzTjM3kwn78
h4EijTIrSq8ksJ8/Vg6uSpbxaP4rHsSIgengNzGRYu26nw6O8FaekClxy1TwrhHr
Tl1WrKOP2zEM8HdHL9V5ZQJnJVJqP1v8Xs7EonVF/KoM3ltXXyjmpaFYuZ2w3bO8
cNumFYAr9nJeAkMjA30goH5sv745Aj4SyscRLiFP+ioQzuRci5Di2V2FdCZS0OGJ
zGPgKAOfqMxUQo7oDQbbV5+8iQuLuZtP7zX1GLPGpaviJdVGGykLvwEn538iIQBr
y+xfZ8/IxaSOM7BEMvvsk9W/lGxpGpO/TTccV+3/zYEyDgPzOwTmX/3fy6aWr0o3
JkWrHKGQngJ4gLrLs8YZ13dS3yFApk/rStovgOeDiQZ+kT8TILIlabTG240XQDAV
51NBGxbbEPSQuo9WNH6ve2Ht/ZZmwcjMgZRr7MoZNZxKuKNpJK6wVj/edyMMJH6l
KhjEJoBjjBa8xm5MRVAqTOmP1d3XL7XaVi8c9uYW/qUDASHiSxcJPeVj4j1dIyHP
ELVL2KxlbacXazM/xsm0EGRcCy+9vw6YqU/sDuqM8TusEn9w3Dk4C8ubvJePasI4
PxFlfuEyDiM8qllNDnWWDx75QIwOmfL0YFdZ8kvNKvEYZudl9XnuaLw1AeOJDzFt
xtmSeKetK2+V4P4dqB7SeYuGpJY7Oju9ohXTHPRD11PcPvy1HB62OfIzimEzCSCC
wR0NywA4+IEEF2EmtuX5oYS/K9SJPgwyc2R7TNPFs3kWSnBaVnZOkPWIOzLWvf6e
mYYr3/WftngVPqu6qvUXjD4+HoIU1kRwR28iVUPCmqEvczS9pAMMq4GlraMjxi0c
t5Ug2WnY40T1L1qa2PhyEMlM3ihoEL+0y3kbqY/pjNKXyaApd393/e9pTu5d1yvF
32maLINgLAgN3hNb+gjCXwz7q5pGKmZ9cX33fYu7wfE0E8ZjB0VanQfCBY4gqpvB
evnXbFfcDK3CDYSog4dL6WrCT5stLPgLhsFZ8VAwe2/9K6PtHip/AYWBnOdYLnqx
rBgbJCaS5Bm8cjpZd2CHTUhPLM21uGgQlg1eicciOH/RQwRlM8wizQJsTcS2Z4Vj
hSHUgc1q6q5gzQErgqht1qt0/Mpx/MVA4Xt1FX/tTXxSNu04JOmQLaU7mx4Wloxw
mHyoNX9p8w5ae4NyEhzhFjKpBy3ZU0VWhnAxHNe+7cvtSFr+64v2UeSUDoNN73HD
qfMuisQsdvxox8cIiJQsz53tbs+lw4tu4l1M/cP8nY0AdeDDGYooqCtimdA0+VYM
Ma2NHbEYHz/+cH/uMhWm36nPdI6A9Lgp0JoWZLJB1MjfFFmpIXAkgh0pxXEqfBza
BkZaslxhmCzGz6v3QXDvLawI6EZsrIetsjEKMTDBbmnTN53x8jwDQ9NbaZqB9wvf
/zv8tIFSnXVpaK0zwm4laOShGNQ1ZD9e4alXxJbNbzTTYgh90qvHjif30ox3KSXb
GTIbkOKYRPy4ciE0Dm/5O9Yuu8blOWAcgKmv+Zcq7pERTYgt33DIT2h42+Q+xv3W
/uX2403FuWzW5HYGDiDc7CbclFxmk+a+7LUawKqWB9vkaU93375+912Ep4tvhfaf
yvZ0+DcTjwlDAb4NIxSVAA6GGiiml/arojN4d1fGhoEcHBaM94pUzwiUez6FhbJ3
Zij3rkxW4j1Dp7hkzLYAYjRT+wpceksPmHScl5800hGiedG2eHjXJ3rd4DOm2W4Z
wrl5c+vRnC879nBPgurC6o2ImpbXuMjQ48M0KjLWCgXjDZtE3/M2mD3HizWIDNBl
hDO1MvPXm/a+Cjk7KVkJKcI4Y1EpgFuO5L84fYkezOHGQOBeU88DTmmfKLJdHqpd
HRoT5z+4P+QbMClfQ++WCtpQtbCFHLNFJ2qlnL5V8BsAIHTtfIzBg/U8JmityvUg
Dm8RL9rfX8hRN1DJGeCpocjmiRFawrb96oM3JQKy2il82REpvbn2CGSQQkKLSFKT
+EnFkmcjM7vH+/ro0ORkhSOBi1pkI5IR8FHsKdscgIFP5xIPBdIHvt6abvsHyVgp
ZPzs5P6MlfN4QnoZ84MWW5IhjU670Z5iotvqli5XBEUnFMa4RhpqMWVUfuNlFz5j
ALxkjVRAGBOnP5A2oYuKW8vXpWO8DPIAcX+yd92Z4e35Gim/J2snlNV0BC/oK3xg
K0KQkVV2o5xEvAuMp2d7cW6nNRyt87KU6tESxbW6XK0dmencGrIk6bOO+Mf8cHAP
+NgUnqmd3ZUiwJayXdkE5Nnun/hikUqMGR5na9WXEN1g8A7uGGIhl4yJZ9NvEIfO
2FSahzsqlzHZGJYnhni3f9mJBd2kw5xzvRC+6uZDxHFZB9hBLpRjtcwvl+spWsco
GfeFp4qetpht6asOX6auRXCdI6qm+unayf6834KM6oHZQA7FLTvG8gL8TTM9HZvY
/WSFuHZK+206beFZnECJUSFLt1j5bc41reFOdazVaUpzOGRIT7eN7aaPdK+7rvDa
R8ciAWzcA53Kkuxeh1zk9y5Bla0zhUZnEx3d3bTY8VxVoeJ6zx2Dpe3HpjoKq13v
keQ6ZREu/iRHznqIJJROLEiS6pGZugbF8gCHs+4fIJQZIpVWj41LP9eZxV7PWLSl
uppRAAHNr3wXk0Pg3D74Dwp2cON+imHHtcVcQZLJpTVfBEjBXpL4JAxC096uoNOm
tmg1jdc/332b0TBWXfg19KOSdCCjx41uEi4jWnqxH01HGblHXESAa+CHkbew+Rw8
dVX6n3jFbYKVvtXYLUWGiUDTkQwkuAlMR9OtKYDNuKOHLN4qnBjuwocH8ILO3P+w
le1EdQPk9Ag9xWWa3R2L6jrsuyJL7CPEddkBs6/E0rYtzU8z5qhbOlNb4be4Pr0x
Vr5XPp0AjYyzWlQY0VaKKBtlTx3K/adC81WddStuRXuyS4gHOj0TopxB9wGq4PLq
l9r9+Y8smMX16w/r8ceMu5mKDI8R0ZS7I7ysoDpgAuwD2bdsJsS8J3XGyiQi+TKF
+29W75f8bQpnQagGvOuZlpyKgnldbfhzuUqIKGh9SsSmCaehuxoSZCA5ZVthnX5/
o+1wjXnH87xke1jRatYlrkSS0+YWUtwfZHhoTXBpjD6LYwFdguXICj2PhL11tGwz
xbgk2BJf5x/z3Q7bKpLcIZ+IZwI2xpybjXQIg3xagOWHeVFqn8wniUuKUwy9eWNV
ffgI/Wu/BjSqfO8Ts+nDxZuREwq0jQLrE8Vjn6+uvIUsWC+d3ci2B+bJhOGX8qIe
CxB2scY2za16vuYY7axrtDrzt+ve5LZ4nb2GzE4taIMDFKvCpgbLP5rcYiAuZBbf
NuqXyy0Dx11uUwXw67dBgCyWYIneLNtVtK4Si1tSCH4URFF6LuqgExlhJlBF9xcY
RJkKcz58QzvaFOjytv0cprV47x9PFrvQ4iAyNZo8xs6GmcAPXCWmkYhMfMgFSFDR
FTK0x6+V/fg2ub+phsA6tc9IuQ/S3ksXeCYmF1CU65ylfuIe2Xhgl03ta+QJdfTb
2TgQHX/fJAeUqlZS6zEZSn/tQOFMzNSyD+UrAvwPJOg7bVJUHnFa70bySn704HRP
lJaZMyy7wWb1osXjjktkGcNr1Mz/jaoEa3YoMKPAXDwUYDXxsoT51xIUrfAIFZJg
fkptPzwUXJYL1uRBINRzrGMbO+N8BMZYr5k85mU7dNuPBO3Qr2BDDEnOEfHhE7uj
EXGl7IE1BwVTG6kiduf/d3HbNu6jazbcsXDsc1L0v4WaqCcJ7IkynbtasKZr7QZg
CSDucUoJMgJPMkOpMOyGovR9YhsUIlNqD7JgxiK8CqKmySlSc5w22isP1brJvCgY
rqY4A4EVlXYcFdKrFkWxCO69zU+cJmXndm8URPeGJM97PimiXBMH+9O4QEtijB1b
VUTfPEr4Z/TWu3JrmNs+FA7dPQjoEjyt2vGWAIblknMyS3tmt5i/Jw8uunE/s/ky
3HkOBroz4V36ftpAqfLOWScgaPvI5qe8O9s6df2djPe+zngSZlzQzURxvxz/G/Dz
0zuyLtGKjKiKl37dViB8yYjHt5PvPj9GQLzqFIMw0nkMGQOOHru203l4pptics+N
2uk4hE37q+HNBI8Y7ZSGNdw/nQcBK6+pyRqr4YPu4Vqc31n/tAtp+BJM6egAlme4
F5/cFeHGAD3vdBvRsh4IK5bz+GrlF3ePAdJeyyg4+fDxc6yp5TpXUYEFWji4Dtg0
4/FVy1mNqgTqVuDvsYIrJsyG8VvfDESWlDxGMFSV2T8LiEvlv+Vpt/D1xyMrLUCi
6ErofiC2g+y8wJwk33gZZdCF2JG5A5upJ3AWb8VvSKXZ4Q/F8AzJBRg8gk0RbHcX
9gsAo6hJW2fFTSu+6fgbM6IYaWq15UR4XM/dmL3qHyHIrt5161Rtlo62LWgtXNlN
7z6yUgdgoidIiBxsIk0xOM4IvjT7WDx3Flf5l47Ld9sjX8FkIHEKVMRcd6CQJfpF
QPSvXvzPvFYBrJVPaslspJY9b6Dx858gn4p1zHjcStmTd2THO6NfhUzHYpk3Zf6l
ds0+rFWGS++9a1ikSlR5s+882KAiv3xWkUGtVAbQBe3Exh6tiZRLHfleEyDnhje4
IMKo087tOH9DLWQGgPDOWqlLPCwDmbHKj/gmvLGWFAOV1aGtowjlmH3lVmJit3cz
hxXjARY7XLmf2bqLyuGl6j47U0r2rSpPplKJUncHX7MmOUrzmZ0Op3A0hD1MTl/4
OOCjcj1dDioVhwUXQo0fmENDkuJWtnLb1nEgICwLQgd5Mf3YABzzj2CwumXKYRKg
Fu0Y46MOlyD7YOlmi1E9u9Qb1cdz66Q9XXw7jE9QSylK+BVOtqdQCR6vW3K2Y2ex
NL9Skd5zkIhXD2DDeeKe+e4ehzqunUshQUXi3mOWKH37z5kBcBMASzM4SITrgVb5
abgkEizL9awefsidkN0Ze8FBcq8dann3E5vb9V8RXOYGkFN/8mpeUOn9Q5m7YrY1
6Hze8wZwvYnmjyt1ec7rNdIgB/74MyDZ9oyaAVn7J5Yyu3W3cqKhz1Gu1+ElwW/G
Y9qd44hvNM219BrewwucgJ+TNoXFK+vwYPz0egm+zourhDGODh6Ni4hPcfBFc/jX
7ysgQj/ghYYv6xm7jtHV/dQYEkfEntQ4OX8nOFh+QOPHWf3OckIMsufb8ig1SBDt
p1rSWqqMlenwvOuxl/CTxpPdJGi4BOr1u14+BO0z0Q2+FPG07hgQr+1ZAmMKhMSD
pc3RO097/Za9xArCOmaP78uoN5a8ABDiJYnqaxMgmJc6IRA6E++PECPuc4cj3w/P
dm9hkuMxLjHzD5PEsG/HyvwhueLEaKgAFw8UT/GSTCC1ozSarCm8VzacPc+BhPa1
O9RM8vbkoRFIgr/duEitoD46IRftPuFPSnsd4qnxvjw7Nma1cLc/KOG5g9rxJgzT
eT6bgpTkki4VrYs/Y7g8IyvO13Ys1k08AQzs7xfl86wws//VlXuQiHM6x9puewFj
tKiPEj/43f+hKLygpsiezjPGhAxin+LepgzVcVBg+ZFNKo+SewpOxdnR2cUGUIdf
Gm9hgklbEnCmBFeBDAqsdKWtnczbZfno/BYtmBvbq8okNuivPEIQ7jz5H8oD/cKj
19nOm0PHh0ky7wqV/364EO9ydlUdihzBdAhkYsmuYkIDNLmVRiJXhyPbI1741rU8
eeGVa76AC4DWPtwsFcWEVk/TnFarKjMnDkoQlODw8xc/mJKJSPzb9GYy4zrtXSTU
dH+IIveCnWx3PMUBHmDpRc+tiv6CNYs6YRV/d1mk1pMrlmiVw3WlylfI8uBhf/7o
S2sNQYRCGhoe/refoUlPQEznfRsem5HrAUd3zqDjz1HC5QCF35dDSZQRINoEUtwY
THuG2cs1iHv/yuEw/FSU4JlbNV830dQGKa0Ay/BRfAfrVar2rGol/EfS9Ll4DvvW
Bpj7twQz/1ZGzHznOjPQXxldWPuXoyGljr7dDApNrcwL0FjSkR7buJL1rN9pXKWf
UA6527T996Pl/hUaY+MrGsfjyD5jORfH7RdHhHK0OwftKz/nIwzRONNJ4gJ8BgqK
LulQ5TjZH1aADS8PDHKt468frewyWutChYn3t8KFWFy0My0TEaft1B1Ou0BsqQzs
W0mFi219BPwKNoVRCxQ9+LYb176IE6YPmnVlvmXrdTxiLKKzleOX5HR3ubDgS9Eh
rI0i9u9XC66+sNOveFLXwgV7YmkH9WnHirexXA3P6nY1jH/YJRkXf3swa/1ER1wm
HmQPjg+69JVd1iaXuDWl3NAtHg9ho27RGRRi7zasvoyaF6IJq/bTYs2nL28YZsad
3B90EfG3KcGNVe6dsZ/P499CFlhk9CLKajz77wJybr8iAqKcF603xhCvhSJCMAeG
nY+UY4+hdkcNzAkk/lpqXNGRw4lWDVMF+lPc8WWylgONN9OcfRd71anTLgwVKi4L
y2YSXMp4qWOpuLmzcztwoKTzP2g33dSzrC37IcGOmLbjzRckm4x83iT2sTKUxALJ
45ifiDKQ+wHw0pqFCSR9FinHcdK02rT/oKf2PWBbwsPjTOZPDwMdN0NQRRGVHiye
loPRmXKnpu5R+mq+pfmqtTMWsUDIK2gZV8SGJy3PAJWuGOfYcOb1yUSC/R6peXI4
loPgnUFrMizrFxn8RM5QJB2x/DBE5fRbJ9uOSCgoZ1/dMkDxk7mYqZziSx+XXCeV
QSTmJh4K30n+KCVucpT03wwum73tU/04qPTFDzbRy21likwVJ0iDiCLGpS9T16NU
eMn0ECHuV0c+uwVplaGegWgoHUWL+t26W+QpDBHDdZX0+GvRL7nfHM9qWHqOHR7O
TwBY0RC3K7h3DHIUr0KGIn3EqJypg/ZJZapBJNFYLU4Oaaiy2OdKC60EmgRvq97i
l5RzjmlFT+0mhmvO3eqQGf3hvCsa0Mven0FuUFa67dxsrstk03sXusFsa0MaBYMn
NWfz8NBgXayKaUs+wCB3vGuzyQyhSJSX9tE33hPH4yt/kckpo6b0x/4NqaohzGMH
iXRQIrzocfBcg/waDP2Ci0Xf8cfxxOzApG9GcJzre3NU+Qi4w0WS2Zo0KWMXdaww
NxqNo5nKwwQNLH8g+GR2mKA6XL1/myJVv8xsMIw0fCmmH8L4uM7hEDSstfMZh5ZV
FQqC+5O0hDf+M5Vy7rYkNtZdulcNXDTrripD3rOf9mbqC5dU9mdAkqn+4YSgqczb
EbFHS9VesNFnQ+lG7CO9m03bXtgMyrf4dDC4n28rsLgvUtwLGD6hkz6HM1m63n6C
IJqeNrM8q/t7eNv8nOE2JTzyBsykLnZCNgamKgS5wjhTmD4zuqD/ffnoQ8F5x4mY
wvb/qZKEdDFQmTv1fWIikSN8C6GCWxW2z/UScsozmErxjE1VeSdZvibf+WqM1ZBY
SMwOYhBquwsuSDbGec1vjP99RgqUK12HjRdT/kb1rz2PEHx1IplT6sfsu64HzEMT
/kglBQlUE5PtLN5xSfH6EPjvouin+zeozgwt36o/u75uhxqZIy9S0xxYL6MNZoT9
qVN0IbRjxn7HLhuMKN80P53+pshIR4f5RwQK3yfEXzGWvrfWHZU91af9EKWetlrZ
H//fAADNURZdkAj2Uvowa9jCtkvovn5lrFc6VAHwUuYSirRwYr8J0iNVqQRWc0k5
6z5yrQ4rEBizv80oLVTNdv1L84nu6BK8VZAThczmQ6YoAowY1WdMfhL41UmkVzK6
l+Yuf5Zj9mepfcJqTPsVDvRFYQ8tCDXQ9aziIGYvcCKB/bd5TsBpPaYA97lkbsd4
+bgTlFN+MASmvx9v556DmEI2q8J2//Why2KS02mwgmoic88hKgq+s6K/tE3eB8XS
keolV0qUVmlgm0E9Dodtpioe0DkAVnw12j/rFa3NMtqn0X31kxY+RMlNd9pvnTMa
FdDQ8qYc8nMy0jxEtLm/SGh4nnj32TC+xhADWW2KYEv74Vk1fBdYR18JTWrHc/wS
tTL+BeOCswxNDZGbJIUuqrN/Pfnqbd3wYPZYMiVbGsQ0TcWmPljrbwdyXa/qCLYE
OfUOiEVQaaCOe4bBGYeDjDKMa7xhlmn4ptaitNN7nOWFdamJhgOl/UlJpfXPD6r8
xTYM5T5xlsyRKM67R0HLlSWtO2gLKPk/KXdINZLKLSaQtF61P9u6PA0gWaET/ZGq
23B7PTfKca91tXZy5AzaYcccWCZGcadaLD+5Q3IvyGfPVRrnB9q39Vh5RmAPWJYC
Gow9II0WzqxqV9F8ifJzZ18mzLWvZhx8bFIvWacNEKtk5zyGNnJoEmCYDzYry3cx
kG+DK1b0YfQwUAeGt4xSQ/aljpwOvNwiRqcHXN91huXOkJw3iWAf+akwInF7mQQa
4Glx0Jc6p7ymUSLZTrNFlRLIm0MccZciOeqg41eGaoG/TgdeO+7glsylxXAeaPMD
VTYXSsQiQIIA4T2LTgVNn2xZODA7qwA2NJxFaD00HbenW6KLlfOJwygKziFrVVVr
n6z+GYZhYD0cFMd7xMTsrXVPNMjrR43JMU/8M4zrY1vxeFylXnoO5clZJKWkCl/b
lnkx9LvBL5YJ8lV0xK7Nf5Rgza0so1gpzDihkaLXK1zD5lPWlaAwqBsza7U4lAkc
zPgyd0/W78m0xUjVkbaQs/gjfMOiAavediB1+XHdi9i9VqCvRVoXc5A7q/Lrks4T
hBKpSrZ6pFOtXWLxG2eDjNSldCY4H3PY1Jl9kCFE5DZWryPG75C4VfDxnfV7Ew+B
j/xIIoPcZ6UAHywoH/732mSW+2lgkd1UuzTL4rLq7C+gxBPA4XaOV9wi3n1znI7p
/wbaotRSW2MznxdwD2dbrxB3BVQl3piy4xTTgb5wbGJzbn8iZXlY2I3EP6Bt9GtK
20KzwQDZR02W/GDKZCBj6OcJjmh0Mz9Ze0VTE56cDeWkMJqfpUfdzeXuKIGLDljY
mffo9sUOJpSnQdAhlSnJmo8xh38BJ0vmj4Sgd2eQx9f+KsIaSQ+UWrhciTDZIYLr
1+KdfYaiHMV8912QcWTotrzONZsiqHYxGCYVCxUX+x4wcRm7ZYJKPE1gZViZDM/9
LmKmKdW6iH0Gmi1y+dJlgnqjkF81vIK2kY+9+iwWB/xF/zNn+LWMsFMKYSupwzzY
387OYbsF8P6PDtvIQoKVo+mnvKh09Bww7YxNdBxsY7/vtrevwygFnANAKveKR2Jt
FvxXbBWiLE1y3qFRNLhooKhFSppxT68gpRLIpVKC+7jX7inNuxlAwcg6OCL5mI52
0nAjEE9f082+djDqoErH3jLfk6eifu4uNV3ScZ/3CwSv3wjr0wgE/bt0knBNGAzP
fsP/QD1fcx20azDCkpZW9KOcVyt0ls4CwY2J3tD14/HfVHvSRzZzUwj1IhRweejU
Au8v8SOhDYzFinDDg1livjlJLGIKu6FMkis8Zm571zIyXwEm9ipq7m5DhveiVKuQ
MpjmJMUwLly2jfaeIKVuwpW2KJNY+9UEcMxQF/TuVcfNoW36sVtRTYtdlvd6IIcu
vj9MiAn+YiLzZNyUkRu4GL6s9YtHxpK/t9QlXai9CIHyrkicTGnX7R2azol5sfxu
qT0uSoDJl53BXU0gJa8IoyxVDs07loNekqb1GzvCAjOuV9DaUxKtud8FypQGTpNa
PlTzee5cqXD0WsXwiwdfB8LJYzNlOY37ss1WZUp4dNp/Dqe+eDeSHTaftP7mj6dZ
6N7ZJ1YHy79oJ1pUstEJ/P9oRfjM41Wm5y3ajxlXLfStBrM6zVuge/+ipsFo7aqR
KaXes9gLr8y+4c99i1taspdDDmqU7jfc2K1b2Ac33SCOhszRX5kwzYXOwX8D1eKY
ah8M0qfV2pXhae6cZJsiNw47Gr3/72aGGXWVKe5GY/L4i5UxuxsoO13OHyPWnRk9
2F7ALCRN4jzn3iapBBbtU0YbYA3APkzER4UYhODYq1cQ/QXLOINZxsDnJS+W+Dc7
XkXfrQ0911PFE6CQLs4/lKOsNBWo6CBE6/kxSWlCBR2edyJXQcSDyYH5UrDwGm8v
eEcTu/uRbj9RvlVePJ2qZJNulaUC2jgjx0SR1yeEW0dZqg6vBiZ7H64Kv6zsfCI3
DmUQGx5bdRCtnuZlMrkB/u7IgMcAFk4QMgo/bfWG33GYVGuT52jPS263UAwCZjvZ
BkunkgsfSsDtntWP3IH1Us2Csy6yWK7DsZBfNCwB7Fh6tvTeQlhZ2+tohGmRchRe
vRb4/1RWJhhDYNfwlpl/zw22g1cEzKpWAle8+iLTOgcRcAQ3lNC69WW1fCvts6p7
zXEbRIRwuLTgJru+8e8tllukX0iEFOEYW/piajIvMvs/XO75tXzB9CAFQ5JftCW9
8U808BCPxCpQPqyZZ8TTF6hE+NJykdDgyZ8LdCg8n+nGDzyQbVpP5EEcklr8Cqge
XCIJNghJ/zzk0guD0xD73mGejNeBm2QausT5Ez0hUaJpkUUamzhXYMPL8wme8A+c
SUdgfaNgNDUGfE8mge55k87gQsZi6zRFZwWtDDi4O/5IbvWof8sz7jPVHIheHTHY
SUcd3mmFSSbpB6Mkl5IMez2aIhMk2JCe2vV7hkui9NUdOJXG8L9aiHF632ZtJo1U
7VmRUqXxQbEYOkUnT9fne7B4toGwdQ/udzPCwKhCj9UAbeJuzCP/3CvS7Migqway
iDF2PWAynQgYkG0AoWg6yWF8olqQSYyta4iMz6Ei7rYhygYykFiqB7fPnBgUU3GC
J+M2ADkyG7O/G/EfR5FDtXqXdVcXEr3wZTyHV0hLxfK3Vf9EegjfkrrbexBACJb4
WdcpseZFXNtIZ12n+AIkEaqTubditlTEu+gkHjX+xn1mq2bGK8zggkdaZTQTx8ra
8M/l3EekD3ypJocZgWfNQ5l+HqDenyq2F2nGAdaIyqMrQY03cjyCFB43A0ThEqVM
mMxUiKpD9IWqAFyjzYum0W4YA0cL+GYgT5X1Ko+4bEHUsIHVlaVHYVNrxxFlZ9fd
HSgvJWelVveacuYqrNc4S/qUNf/0fZv+Msj7h9AJ5ab9B1mia0QqNuLpJSl3O7M2
pqjaXdl7/wkzszwOAc8fOs9Q60Mek/wQ8Lby6l6q09AMFRF1fEX++PnNe7ouQOcg
l0ll33b3C9VvJgKFdkqjdymKmmZD51uHJVpYYqXjcQM7gdqVp8JeEkyz8Vo6IF8u
MR46gsfRhZ7+kGHt6z0/6mKNv1+LJN/yd2VMBxuwsv3cwV1x6LA6k+RfMGAvZg+Z
8Yg7CHLBnvb9YoG2+auiysyKoilmuhwbvu7vCkoqDrJ0JsDgaalHumYbxtF/2r4D
Wg2gmpqXKxKMGUszHRLOIVTWWX80adVX5svhlgkjx9/oXtI9pW19r7g8SvW5G5yf
OL4TOXYX6Fg3ohSwxgzLmUnaTq1ILDlUiHxOR3irewdjvJw0Nt47GuDXnX+HEOZB
b61ad8s4SJ8UhiN5FIP5qKJR53ejRIdathg4+NbWCbFzp7ZC8i2Bd5MxHPFEyNjV
JIUzRWe1xVbb/F15gr3kfHA7wH8JgFC1AW92Lhgw8FstTTuXpZu7SSvWizH4Y1Of
QwvugJ7eQzSz+UNQBPmkso8/0ojkRBsfGyML/jHBIZWoVChTWNB8F/B0PdvITjn0
88z1rcW855ui12NxSfsjjtL2zRm9WcsR+Qy0GyiBk9JsfQfbg+mmEwYnbexK4mUE
KYMKlqcSHP1bsKFcL+ZySwiwQcZEG5A3UsfkEalkK+vWJd18TYH2oNV89bDLNDtL
Ao82j4p579lQRKS02ierCV6P6N4siwl5qRofi2b+mNgfCNZfiWNWipcMJh0hbtZX
n+tJAl+oR6iRcGy5qw5jM0AiUvwKf2/9qP12+bPYCeTbawu8XzSvgn26T7UCEUEJ
C/4hjiuiVOmPIZeu1kN/n/A2n4ARv+vX2TGSt7jHkS+8ibrOhvDxZFUSs8Ku/sl/
jto3XmVI2ydsL8oRPy5ZnXRv2Bm6ebDQvj8bLm9cBLp8LG1smHHhxM5tEmJ/VEfd
3/qKsDp0a+/ytIFlo/NpBbfjsqdMEvHsOV9RC9QFUrhzU38OfO4P9vpEcV1D2/To
tDBRR78Y5IQFWzlg+V59ESZ9cj+/5adSsk7mYACuDhJAAnOrIhTGLeIqLcCcPjVR
52jzwfXiA/YMo/W5VYwSnBku0DPsp/rINAcc5Yn/7PCDcP0j9qb11vnk6quephc8
/D8X5VBdPHx2d4lW4HuWoUSnokteRezLcOWNr/+kojttXoAc5yXcuNSxR1NadYDV
lfVckjeKubGrIG+MwKMxMWe3ijHrlyIqIeb3hxAbIrpjjYO03mqmOf2HSHbvpjF+
qQKpsdsMsZdf/8kXaJDIbkLY0KaSFv3FYasMzxAT+V14VKQrpv6VgygtE6MWOZgj
3vNBRhsHnBQD60n0vwyeBpz9pn7tq1FNLZBJ+MY8UU4wbsCvgxllH2sWeJ10COAL
ugVEWOoNzFoqMi1+mjUbd+qzc7wVj8FTK4m9JFwqA4XbJyoBBegyGhv6NXpAb3j5
bYQ5fSAWcMCbxp5cchPyCq520AOSn01o2LgCOr3Dfob7Pt6PI+bRlkVRW7SIOyz+
Jpm4ynUrpyH6joryfGfO4OZc7uDHykCoajK/+puSBJvuaD7VA6OBXT5WmythNjeO
0zKh8PiQEoA/RJLxv9JNB3DSIhAjVDFACBu1FmxtH3J1/LpTpvurE6pdzI0A/kNz
SLT0w33U4Lfz53XoasyVp4XMA6A1LMh9eAZDpC0L9z4AKCd03D4POp/KUPY5sTzN
rCwIESj1b+WCm2CpI61bEVXEpbzZC9/MmqrljuhjcipXBcaoTAtiO65RVs1+xnX3
b2IUsuU8dSWvzVns3Y0763LuHfLExTIdCohTaDDx4q3T8qIq55p/HF+2q5OoFAgN
FDRnUmmMm5pmyggm7sxUSt8xzUlAl2dGzmFv3LrTLUgWMUwr0GNeq2IatbGzLhAf
vxxy0lpf+v0tR9w2VEy7mNYuxVyrZ88j9PwzCi8Riv+unW7+BwtzSiOMRDgm5D4y
OUQvC2fFq0e/u3/OH3esFqW5XEqQBn69PgNTH3l4tzV6cdSCJEhpDirKBxh80607
3eijB+xbYjTxRwo7wAObqV5LTGwpKm+alw5n6SDleaXHH0stMb2aSo5nYIZSzkag
3OIZl8RCGEH0U3WbRqDoe/tvUosR6XOJTh3yzIeq+LKAzNErWJ1+bpvDuf98ZGcR
Um6ZfBbZKBSxQj3jJz76jCwWY7gZC36hqZhEHG60BBvZ20V3WR+CsfRiCiJk+Gc0
HvNupec3fAXwUqJ++Ey9TZcsH3rtnwdJ50RNDnzCqSrZJwwC2OikAlENSnj5k2hq
EuDYAgiuGlvRPvQRdU1cEAD9ttZUQHgPaiAVtwbKWzB0k8mQPfAkL9wD59NsnypG
jzlO2sSa/yRHCDghYflGDd+mruO9fcdDaNSPCRVnnzjIlw+eNd+DITUyFDH3Hx+P
9aaQDXbWTLqLmw3csxt/H2dsxCYbIw4TSBXyOGmoeGmwSAovbBj/FV7//klQOFbG
FKGtWnviD5fmbm24r17c7cBjxvRNr3z+DgRd2gHAq9GPUyDfqMhPhEPipZ65W2lS
aDjYgvxW13rQrivfKAYyiWcNl43j1yE+TAHzA8g71iZ1Y2nTPovFi9EtDhtd9nwO
AmNtQ9ozdTXraCej5CxHybNlqrnD8UnS/QKeA16t8vKRH8bVE6n7JYioQ4VLRWd3
2tTqnZnUflHMmoI8IBk2aSWt244WX0ImXFBe8tP9ZlHnrmk0ht+Qcpc3wRYkKDc/
ioBySiW8JUDnSSHKisiMePF2nfUKnCyjzgjgXenzhmAQjnUQ1Z0AvCZp4cryekkZ
D3Dg9uSZe2vg2iQsIQ24BGNhqxzo4yWct9pQCLh4n06vBdWCocklAwU0sJgIim4q
CvLYYqfz8YIELvFMfSDAhOlTv14z43B6KXun5/V/DcgFIQTj9ZjuoUWVTkQ4IT53
1smHGghrrVnJSzT+pu/pjTPXnTv6+Nc+1m9oDW3FWmBOwLxp85pE4DGksVB9kIZm
hYP/dv3i/jPjEzaQmyci1Hb6sAU4vaXy7tOHsaHokwi/jqW8Q3M35UEMOZcWKdRS
5eT6IHQtxaqoiPjlzQfZegDO2Mm8DUd0JYiJBQBKwquzUI18FSEJRN2JapeflNWT
VyMYInh2tfcXs/DpePHHmDb18orBBADFLvIkLOlxOZk+6zAwPaWpIBEis9pTyTe3
PbrocM1DNc7GLcOEM47Vy8RBgvV2ilbZoKbcloag+eIqlrEOa4bAiW4ijds+boTf
4dmVJOUZS7ov/WO6JhkzbfMGtoeYum32L6c/bGNnh/6KBRY3+Y3qfxL0PmEzdka1
oKW0FmaG/lFURVKn+SKT14egeK3cLb47meARP8lpNwixbvuRC1XgUcHAPK93B2J/
X5ODbBLPkXKBZFsIh65AP2j/kBPGjX5QmTDdXWjheqTsJNVK0MD2bUS+Q483TXnx
GvpE2Ty3d5JAzjjonvriJIbvMDYsBerREuaFo2krbgPVqvRDJDq50sYfko5e5qI+
2ridMXSKJjDMPuPPXOFuWM/veJLuEjz7URAp1tOt9l+nhH626HI0Eez8Dw4Vbhur
89k/ChvvnM8shuie3DebdkSwLW/f1okYTq3TvV3RYvz4vjanxZZizYwXh7h8oBXF
UdQ/r1BtLQDhg7aTgoRlZyT/THaShI7ZkcmJiufU7Q6Bp+7I26s9oHsecQutEqC2
Wz2F9QWbQvl5ogZdyiXC0MlUzR5MESEmd/fbSzhoj5c+Aw5Wb3Ado8W8KYlT8EuE
bTGjjtBB7UWq9Jv1PY6WjXCwazavSjDNIhWy+fEOPl7XdildpCsZiHJXO0nn93hu
6HxRbEZiIv528RHiossrX08/pdE+jK4CA1J/bOmjcxATMhj0aSc0tm6q0wLvEHPT
a6m4tNKXr43wBS2LCg9JtX5N+a2X4c9Z98YKupiRiw6bjLuRLLk8fem6cpyPptDj
C3VcJyXLhplJ4meEphrvOjeVOJ0on4S7YpCyttaeBhZrVR/B0zY+lVUEeJpkshCX
uIJMJcL6aQmGOVTfnzibhuh4eprn6xWErL2+SWDlHXuAWFpe6RlANKELqYq1aTBi
PaiXaPYxbm5AISkhvnT8o8nCXnofSZrtH0h5h/6wSHzIHdiYqsl6nd8/jPmERPm6
FyG8Nank/1Ts3ELEEMNT+zZIs+8VUxU1jlN1l9Kbko9sRxxiBEmSDnqosqnWrdGK
uEEs9ycudwQm+Kcy/AVYfH948xsjRHG6pZsQvgAgQA25KoXT4j+ROUu614YsZ/ss
SEAz1xIucGCKGFizyG+Gxan7q38bZfa4lQv76yOmQtFfpPcd2GX6J3W8Pp+wPCiQ
ZRh0L08A7Z/inUmt+xcP7Rg9NyTYi77WGE2ZitnU8MhFcmKjiHiIV9Tkd5CwG1DQ
kPZ8uIAS8Yrny4EkXJdi8MtNTAoLu1+r5oaqm8rMrJfjXg1ENUuDBWoP2zVEzC07
InHv2a6YBZdxQU6fmCSjtkggoepv8TwkXEwM0IaH4HatMQAl+bJE4/e8MKyM5NPv
wOhA+bn/rEqifnWbywhO5cVt+kp1i2P+DDcQYwqIveEaQYzhHL95Zywy/btd3pF7
H+pn3CTI1yJbaoOQHU1TzQwjZiDiF0LyQYpRc52O8PC0rllcMZoyJ9j1I5220Jrm
RsY5NKpb0qo/2M2no2jkWefxTB4WZzXt/WLNVKADHsMdtVDjxnSYQ0lGg51bdj19
QvjjKHx26UyJbWbc0raXDH7xKJ1by74Uud57BWo/TR+AWy0hT7Mi21e92ZkcaYT1
wBffJ1IFhypV2Xopb1mhxXN5pmR8lhWVKWi6LxMxwj8peJKznDitnf5VGrxkbU2q
yaRQRsknegG4JCrcIMKtQY92zxVnX95wZO4JeRGQc5ATUkzbvkOWGG9l3M5Hj9j9
7/Q8R2HPRHmIf3ECze9/Z3Lwtksu2BbY1ECvXHvOUCGbqT5+cNX20k3dXnC9FeRQ
9YDawfMGemFBa7TfVwgy1WucOfTvsZT/KWemPvptoDiUUkW1RKTCCdQM4Ohy1N6w
rNOJMh7s/9zJ/UJXBlbtL6hxSDlkEjbx6tAWxZ9+opb1eGSf7TNnuwP/T1NJiLuW
3vcJ/Rj1gHCQj/88hAvqRopIMQQLvB+nkhSg1aZia/2ySbFEhPDRxOZp00bHOjkm
8Brz/AOKki3gBUqFSXz87i0raU74jDfSa1d58wsyHFgIgbZqc6DHfjXh5FlOQR6b
4ila2yPGvr9IhufHTbVNajyyGu8HANZsgeaVldy+3XEJN1KHB+xBCu7VOsQehUFw
0ljk665RKFXSFEtqhlJovdVt115eTYZ1629otLquqh8sJCIWuoSy69hexXDonpNX
fm6RRDQSdVGB33uhbk36EOoJ3ZdBBGf0UMgh/JsNOHgXtuagtaLyjVCTKK2kTXJL
Ajxvqe0nVumRjEc3F/PimxfgGuF1EN0gsexTvkN0lts9Efq+unZX22qxpyExQbRM
Bb5rLJgPa5s+f4AfOB0v2ugpJJv+dBhfmIQ4l70Qz/855mhYqJhTUCDN9iAMxHsY
kCsqCMQi236nL+mrNNDn3mTLdTvN+0Y6WPVbrf5RTdSfk7C7759WfVSFBuG83uJN
GjZtxOpmxo77A7+/cDAoSKh5NEw6Mn/OZU9QRI6NP0nfsC8l/Fw9EyJnTKJNxIYV
AtWOe2eutRiQxv+bh3jbaT1SmHCz28jJKqEbW7dcwLvv+td9DBB5JXNKioENeS/P
VxAYvKZ692Odu5uHN3J4q9Ae6lZldYV1aVy+F8yla4uBQQ9Mju1KT+R0UYWoGywA
nYxWl56+HoDnVMd7Rv47mX4QDjbIsD/RTs4xSO2oAZWUWKQbLjoTv81orF8hEIC/
MkoTWnUp3KDsqzLrkYAHhvMQICnvWGvbS7W90rAZ+ZbPa9kHm30j+/PJtLU2NZRP
J+kb0zuRsePQantQ+Z7b+IYnM/pd3m9UCdOMUPkX84o/fGFpJ0IiyN/bGL6cmrQX
Un3u8zxFbGHhCHyGPNaXnflCoZMwaijZDJHy9F+u8XcKAXbJLD+hsIU1WOJokIdG
XvM3+XgRZqixUEn2AjB4u6LQGZUjV0SsOwT5d6uT1RCJyN7r/GiI6rk+oTaFa0E5
GJ8Fa0EtaOsyhVLI7Q9fR/JJonzs9nS+FO8syQ0cew9s5TEihgc2oRnArp3E8QKQ
g67VM4euv1c1pMuEI1EpcpRKk/jnKVHOIK1CbClHt8Ra/IZaDNKuXHw+tcbnCU/Z
uvaHb1L/Y8kI07t9FrBcFFi+HY3EQzREUEMppFtoLJQDpQrvW7ozLF9lq8FKSpff
TMAgITZtos1aUqCG88k0ON/s7ExoRTA/ySuPukSc/W+DTZwtLkkfU3ffahd2UMOm
khvvsN/p8EqjRJ04pAN3deuS413nwgE1jz5mQn8XsbdYogdl1gW2oWy1tadZhEWg
4GuytGQJtwmnnEI8qOm7lXImMA9Q1jjRvNeEWneiczdyPKd1/s69QcQGNkUyIGXl
SCmZH4FgkdoobA4TTfvZpN50eVCz8U2M0SBz0cX7sZuxNPNL//OeGzj6IO64FAj7
pQlHZrqOoRXeWNRdp0deolTDBkqgc65SKWIvTqpuIcPZs6I+v9Yl+h6lm7Gk6ifY
hgaSwaRGiQ1WD5Lh/RqJgSF5PfrXmrClgXjO/re4QREYLeTnczzu3wAq+ZEyB/h0
xDuVtTsdXMXBFuN2n+u1UbaeBTwhTESk/891gWiSuTv8Wt/+oK9AafJ9K2mL3tEb
EquN6Vj421OGNDg9dClKRA7sWPWh3k2mBQEmGZhU2dy4H+ua0OB6AS55BZamSPeQ
Ar+Csz8iHzadPr4A5wSD5XMMFYFrCA/fZW3+W24Uxkb+bvxrr1/c9nTqnqbOGfeF
oiLDI6Wweh+1ygwbrGdNc0s5V2KnTvc6fXosMAoOfRAQBlX0zTXz0XqHgBEoUiYs
suzb8WGCP5FjsuNsqlk2IiqA5vMrTAjQD4KoRx3VOZ/Q3Et/YL9ht3sm2OqK7hn7
MX/otOenRn0VVzdtwEBB5ahEza0j/06OtRSLgnNt3Fq5tzW/HNwEbW8gxGNX71Ue
xs9vSwx8QZIOnQZ/igHdiq9VtHLt5m6s3NDK8KR/P7OQqQ+Nzxi/JYsFEKy69Idz
Epwv1mV2oUts/5B6M1jQaXcE+Kc2Y0XpuAoKvsOwTS77I+i8kUtxpjpLs+nPvrAG
SIuJh46kgv+EdHWzczxtYn6DR8ispftt4kDtYDSFZm7VqfoIlcqe+ZmfTs0hGPkR
5CXoRwsTfCZ9Xm2M127CR7hFadqe4/t0wNbM7zKbc9gmfzWazaq9KnA9U5CnI6HR
5QsGxmGDcn2E5Gsg851bBI+6dNBH73TjfHzdRhOppZ8sNZ7yDJAIwvA7oo9yKAFa
EG86q8R9S/FVKjqVms0jyZR43qGV2hnOAmFbV9wl0JLaQMu8v5g1oOn2rVM0dpkK
BGgHVWAehIXimA/0cC4tYQf1fIO+9xc8SPgERbTCXH8+EDtmhNm6W0Apt713qXku
C1bI6OQd1AhwPgz9enSr9RnRd+hv9b4I1brGC/xeCb0zKi2+5zndISgE9xzjqdW7
Jm46tY6AHPRyd6rqldk5Ed2KqQN778ucrMP8rI8OL1ULjhSOOiD8+q289sZMkbZO
2iKa9STeMCTt7+PtHEHre2/BvVD2gOIW+mvZhMjY3PAR4KoU0LlRrN3Am5x6EG7V
zrzH0h3iLm352ABuIssDxqkv6iq42DEF3t0rkbqqnGcmFs/eKPzrJH3P/Bcq1ydv
vJQ1CQ82ySOmtRsuZCEBicp9yfnzrwgD6eHnMXBVPDyYj4Y4Qsf1lsTQsxu2ZABT
uFu/RZR9CeheUug+zMSoW4KFf/bKINrwkrcreqCegJV276EvABK+5koAp5hn3ZGR
vopYLPXfVFua91cdXeFRgkUss+nV8IA8GEbDSJ/fUKtthVVJdWlvAEkvnSfVqelL
bOBbMRbBcT1xpmJM4to5kaDG5u7Y3OWB1Xl4FTyYi28k17mLtkSc+Bf8uOR8eqrm
Y9ZUFEnOzjtfjCaBuj2OP7+7eZtlxLv6qyl+pl5OovjOCb9Nb85QTRHkWg5KjbNv
RUg5H0Dsh5XoHj7MVgb6WBqKIqO8+UZltDD7im1Q6ZE+y5NS9UhjyHHRy7PAnERw
eG6RJU+yorWL20ETIapOZCA60J6nh5ZeoumuaudVt9qDvk2/FXXsJXa9Ves0OJDy
7oWgbpORet7NhXh9qYTsP+MpQ9F9BA0TSA4ZI5/dWOMe66FG5y23GsEpQS2/Lf6X
qh+S8GGwhQty8KAGeZNBuUcj8pnR4b1bYpsrjqiTjUQh0AYhlf/I2v+u8qKSrdXT
Iemf+K/LnKM1cO992z+wBxoqibj2LCdJ5SsRx4l/b9knVjOlZ5flHEHdnqBp9cUG
sdVOKxvIlEm3sech40Inca0H3LiqcqBlJorK/5RQyyr7SOf1U5JIEh47NP+Hpb0z
NFwlyD5sE75ONx0tP08sZipPXgqRpGF9KJ285wUYx286Wchzv5p2Qt/hXoG6qHrK
smW0OUr2GQGwZJc4c8EmkfIzULMowKzQpX93peRMfAobMf5jModT9CC3fUJumT9A
cL4pnGe8kGPlwoqKEhoYOnxJmojPbjmVXut87Gln+T+a7kHX61FBWAZHrQVvxknr
jZIGHf+k2y6Of0Ivvs909JD1XiuUTIdu9r60aJvbBdxBoRkVe0QRUIg056ail1EX
aUWkOZ49UjgsPfAe1Azkhz+9iRCdMuSeyMSRhfF1TqXLuFoCPKWPDujxRzNTvHaZ
c6gAjwyPiypsVu/msypbd9DZjhKuau5eCBy9eKfLap74CueIDhGzvku80yDTOu17
qAbt3+p/8FRKq/gDUN9gMTCyNAweVE6EWAkZ/PcMZQhpb1shgwoFCI6mAcE+nY4t
W+6JXxl4sWptxAdNUV6z7akqrVb6sWcdX5cDJOj//6RaBK3D5G0URKN27Q34MKqk
qb3V6PD4QmDLwDBRxlRPEtPgT8NZqIs4AA4rLyJStQK/ZhTZrhQba5yxZSegHjhB
x9XbHX3awDIvQ3Hy1Gomg1sFTsKNo5q0QihGYpx7A5Rsgyx2+NL7pwR5xBy+bgQs
XnF9piitDUKpSCS6oyjJVPlEHmlj6RwlJ+d2SAA4TffeThFTpeLDJMhB8oeEfaOR
Pf8wnyAFOEjEoIF/C13z76GRmz4ZE7+dF6+f8dO9qdGd+Ch7vWV6wBR3wWMEi6a1
4MYIC7IjdEdwuX89k3adCew3Z3LZdXZVcAPG6LbNk+E8OKy0+UsFWf/syNsxkN6D
9bP/ba4WiMhvI4Ve/fOYXwoEfbvutQgC3Dd2yArVnJk5Feb28J18a8f8PX+7p/aU
6WmIIKXAkwKosS+yN2WW/JTGQFay2tNCDuUeqsYI1VMW/B4x5oRhxKYekcxtv0b8
cpP42SPWuA0HlPV7yHn6c0VZuDm8xoiwtz70qcq9OnQ0fsN3LjEQZxi00HHwk2Aq
bqZoIEkKbvdn95Pe/Qq3CThUT8vA/Py91QGddiK2aHcewWEVdOlpVL2yaDmX/n/g
TQDIEo4UfogbnJjzagihsj3EXP4XoEvGagePV3jaSri9JA0fhXjctah49fgCjOSC
mAcZUc0vFrCrOs6UCSHTsBgYvwodmmS0f6Vqqb6fKo2tQ5yMY+RPDRkesJstCHyG
bjJ9S6ttvd30mpf5OU0Z3BaSEj6ugQ6EaMIQg4pBUiCqngvMlWTmi5SEjUrPZi6F
eB5T6Bs/bLgXBTIwCi5O9pk6MSlTwaZcB2r3hBneiI3Udj/oa9YL8u/j1QStREab
1baq9Ax3Zmc7T1VSUYMmFzuTvA0gRMNI+7LcF7dzaIUFu4Twa+vNZ9z7CYjYtsTT
E48jC/O8WMsE+z1ru+hqUnDOkyuPuCIdxH2aBKbwHbjb0q2gwtRkMRnGNaoXaicf
EK5dctmYC/IjVPRiaZaKfQ10texTTiPvb3Flg+uSMDaUiD+Oapr+EZu7I4C0qr76
oma2/Ksmo5s592M6DxLnJ+3R5mXqudqduKerrf2UQ6XEoPmIhkjrTFmbHCDVO0ox
8rOuojV30QQl+rRoooTYcU9qGoOoertEEz9VkGuYO24rvXGiqUQOGWfdVB7y0k5K
9ss6loY+n+CdNk5GFkCrmMk3PAnf9eAU9tCWAQdBnQNyzJwBqMI69rDlubaVCuy6
Yd0KC7WkDCV9ivcQH1hmG7qLQM1gvBHuGXgohEXCVinHiLeo6Y2kPydZaw6Ttyom
Tmkzl2dAjzPu/qBQ+wekDutvYb4ISwBVDPWRFOY7lIepPrhAAS3ZhKioT8jZB4lB
SyFrRtaMjTgJIl11xYKlhkvGP3HJ0S03lnWb4Zv9p6R2ZHOEtRaE9sEct1KrpWpK
TvmHTS4xrKAdcTpalyrde/hc85Okqs1AL/IcBA2O4QYhrrFxQNOvjMoud4TeL88m
zDuxVuCK7lU7CoWj6zkIR60bw4dfxOy+T19/6UAA6cjvJNzgpBHYeg2XsYL9e6QV
sJRahl5GW4XuuILFRV8WIIRrHOl/WrOQ8mhqazthBq97TuFoZhwejhpofVi0MnWK
kppAbVXPXPkyWpNr4js1PQVOvC9oWIHGKbCnKaySgyYw20AUngWRd1g3aCzZfkPX
yigVG7LoBuTgDgvKq0SQRcJSSlI5YXyaASP00VaixgCE7//HsRkIoNhUItdiuR8t
jJAO7dYB5wyDB3XbBMo/m19IxKsHjqKVjSp7mYvBGgbppO93n9DKa1gohBkSLo4t
3p60cP08M5wTjVbuKvLkn72SsGFj54gSg60oQfc3G8oBMzfZ91Mfhx5Mx3VYZYF5
EPKEe7pJo5l6cIWBKpO5NoznwroB+gb53EtI3ty2STRGV1a6jczw/HkhpaR04Vb7
0HCWWKYQHaztymDv5vz31y6NPeq41rd4K80wZLFf7WinYTPfy1niU24kzyOrpbjp
R1UfIIFvBZGlO2enbf7r50JgF/zxcxkh9nWEHY8qLp0e4hG+Q9WYgw/8r4wgIzzE
vGxWenZak0SXFD6UW8qAPxYBPYRAHNrhnzQ9qceipEHc3reSFXw2D9Kp8SoQGrDz
gJrYvGuhzEB4JeQe7ayBwY9N2JUixCHPo+3G1YLojuRR/62Se+lUtmhE3At0qAFY
2nYcawEwnnqOJW1BHr/O2iVCbFr6n+l3VyAGO5Hbw6+KK3uoqG/nq4F8bcDOThN4
b0lGc7soDV5qhCLaNm+nfNmN7Owmxsp0JjKnfsstt3n9YwtVf1FQow36221Ncrgi
yBFG6UfmCKPDhvQk58Wlw+Ytz0DVDj+eCltGfX4lDaixdap7j5FVFhpdFSieGCsP
UQexa4i9gOKmKcRmephu3E9J+mKCq5m39EaPXHtEFv21DLtTO9QZBmapWL2t9aDp
sr04V3FKwCUzaEvmTrUyADZ9SKFRkz7NypORPlJDNVVME0GLo52MIoEY5QtdM3S3
FgD4pEF7DDRTpG2ZFqISYR7LLt/yM195X+oltxi7Q/1sOOX85AjTwONrnPAuIcBI
icaAwHAkCRXa+Ai+IbRtm+sTQ9qyOnSGJXkPTm1PCbZMSXczDC/1TABw4UNTj1v0
xrvvVYrFfvYJpQswJB3fq4WMBt4sd2nlBgvlHgd+EHy7ibeunfFsVar5F/UMwO+A
kyi267sK8aujLytwxNUX1edkwCYY3YMfnyrzZx23hIVTNLJsESXJovsiOP61dHUA
j19F41jfTwV1t5GoG9Sq6GLKf5Crm8ytXy0C8L+xGzEAl4RL1cJGFw5y/PtRYtSI
S+haSXbI9ErIB2YO+Sdsrag/AzVL/fwHVYVnlx1tqJrSjB+lotMLqUp4xdKOOTYu
5hP4uWcTKYgjLg3AEicvHImmol+to5eLfpzhZNbr9VrD9k3EMv7tznJlr0j4RdT/
Ww+t43tmF7hiPkS4X988EkDcot94y518c24NFDSlR1dhfDes/PhSWR3+69YKOrzS
ocpd/rTdiILSyQB1F5v/morrwWi4EnzZpD0NxUi842HMuYy/LzMsA8ulnk31TH0t
PSonY0sTDqy8ZNCa71lWNviLm81I8sc4j8/vUpRxmIEK6EvLvtVs2ELQC45o/Mxx
B7Fi1ZMb6zEDs5MKVZII1pGvqBpc6tzC2gTxoOochq/BHbHzZCZ6Nb8CJJWmsUW/
pRrCVfM39XYU2qnG9byO4e0fgM9b3KiK99obyA4YxyJ4fS7R3U1ZQwAWw7HpH9hz
1GamoNz5wEU6386/TRvOqC5ZWplqufykxmHfiS86EzToNIKw2t8xmtUFMBj177dn
CFMTdra91e/MrteeI2ybyYTcBic5M1QzEtpHa/+ra9xUMzvCEn/tdypwQhx91Twu
4CZbjhc7CxAQh2+VzuXjc/IHiexMex6N3q+rlKY2X8wwPP2PrZ43b0sYrtMJnDDQ
xV7cDlQjewIKHbe+d9k05T9xFb0e7H4Szfq8kx4VHaPOZYfuIHaXPVf9tBx3foQC
tR5PWt37N6TpvKGg4HsysFx3J/DQi0AffMn3nvBBUQlYONK49BcCu1jJxgHuTfMz
Q24yPwWdIWH6R1LGp37APXjcJZb7wBAKBkVEvuCOEZzpBavyDjr+6fjGrW++JFqD
d+Ugd8Z8RaJIHQr1RQo7Wu56IQ+vPk6RTWeDUTSunjdzOHSSLBQ2lW4OPOdrsih6
NhZrVKA3aax7ORNhjrQk7iT1+56+Cd+YnHIXxuLDkwNrOxwZJo97eCYud21VWxog
9yqhJBF1Bgj6K1dW2rQnH9hmeinkSKz1AUucoa0Jl9IbiQ6iJ1i6HNs+TAJX5Y8E
hO/Bk7Wi60BO359OyD9wMFfEIUFLCeaAqLMsjFk29KuYbBTbse2Mf1GLZinoZKlY
43iydrnMrmpdiaKQdAxTUfGkE0PfNsO0EGQuAfPvQnRswRaswiD3vPGnafL8Y60I
VQDMnWCsJuCWvMppg0pJMWmCULTNN0n326WBBmPYFeuAHlnhGUZ0feHpqE8LHi0A
wCAyF8WpvO2BWmynSe1NImXIo5kt2+5q5Z64qKF/o2wkEm0O+YVTJ4CpgW2k682y
VRmRMiHPow9YE7UunRQOnROGG9lS5PDfvSuUOBwM5gqbWksmEspdSuBWzfSMLjiZ
QAfBY/sh97xic3FYlWZUyr6ky6j1zkcYWl2roq4UTZkqLnsV9ZoIGuVAZYpG1X5C
0+Y2egD00daTeh7JNI0kHxB4wz/iQnT8GuHYOVxOUFtSML7xAOfhjI2SEl6qj8rP
XwVe+5dzxdEQlBg5vqDidcdiriz2ZHtznpqYBVMU45ZM4POYFnuRd7oslDlc2534
oS0KIruGi/goyFlY8SBzi2vftLNMcjtvhTDYOwnz0PiLCBoZ9p3kVAThWm2f63lg
SiFPbDQu40CsxWngRJrG54vSkzd3jhY82KsxSVK6KdlNxS5yV1rn09lzB40M9woY
R1aEuzvD1hYi42bAf4SDE949MFH0wZ8jtcM1j8pRhj0b3xF5IiqYH3evawgDl9Nj
OQVs4sdW5h2JxOAVb4f5892l4nahuvDeGACS+QopJxF+Mc1ByEtaSNInZgtzBbcu
x0FPabRmTjgs4MEAnoe2/KhINynxwGt5+8UHtitf3z5Fjhwi4v3wt/IGZQ1r4L+z
rgcidf2muOy+WwlV9pZRSaq/Js8wj+HSp+ldvl625H2UyJPCXq2NMWmbOOWCj2Ul
BluKCiOW6LetnYqtriIwGILQy09VvnAgDvYujviQ5KYRRyuhcbcwjmXoh3j3fkkM
wYd3aIf/uAion62winX7leF+/U6Vr4gliWd5oMzKDv71/75KLdXYm6dUu43ckHaD
gcBbJvTsxNX9P9phbfGsWq+MDtSYn57L0TD0CRic+ESGrCZBNMsgL+cfAy2D3z2+
E2w9iKmsHy2p6vIINbZth2M5ykYH7+yHI71QclQrqAdb15mduaAR6xT9TInhCUum
zECQvyvXjwa6ZOnQhDahhuIv1B7TQ/aZvl0niyhQoIlG/2p6WWj/I+zo9ivNI/I/
CSi6eX4XuqatPD5Rc/hcY1lVPXehSnzz6/xpcaw1kQ23aqoOLV6ErQECDD6+86wP
LYAEgG9Dj6oMfjeCzBpZGPQHD/MOVS3IjrgOemK1U/h6e+Cbhuga6JochafdE2+0
FYs6EtgDnUopxSnZemfrQi8oNT02u+RPzjO/T3lscqVoEcx/Sw2ObasjBqcf5ZoW
BRCutpMl0e8AM3JKRCfVpKKCH45ZoFX+Qf45ZTfyxyxDI+cFfINX/pLq62QHJKk/
Dfy5j1oFuQ0nUv8u/2MXgSFLTw/0IwoeRsxNrpSmbcypxXTTuhvSszIdhESzFJzS
XAFpD61evySDkpM1U4V8izdojhmIEtmHelpc+oxTAVodvrZ8AcfVQ3YI3YalqFYe
WD69IgPzWHXzyAjFn5hD37Ed4NPwZuvZxGwZAJpsle1ejZ8N4ZGhDT385eoFU3+R
2+GJq6GLsNCOUauz1s1PGlPXtgj1NtG/3L3lihhhaxrkTbfbZ5N5JGh9FqmlML6h
BTLp8unKajVfRJUtoFENFAngA7Y82eD8mM+7BEt7tSjvz/EKDbk3KCtq4nIBZ8Bs
iYzXhwzzQ3jz1Rt4NWo0p11XkZNy83H+tQDiU7GWUak4/oh0Iweacu0tAVJ9QxyD
LeqAEQ5iqIvti0FPIvCqbqvXNaRy0yuUKfRWmc1QmmZxIGbeUwKcoChHo7Qnks7Q
e1syWPg3Ut0YIYsqpahvaiBAYI5zNcl7pCgQaEV0eswC38Lg/Ula1Q60AauIOv3v
CJCAWHIYVJs4xNb3tyC36WlTrAqVN90RfNtfWU8vv+9beU8E8soO1k7JSkz8LeP/
5AYcEAKy8NDY5ZjwtiuWApPR4bLUWgtXmM2pMRV09KUvfbAVYjguJE+/t0htsmiE
8AmTTFY0dc/NOoJXGZMaUo9mbGGebwxP3NQjQq3HucpmT+q1blJe+lI5fOygA9az
pe1bZ32QYmeJa60I7QsrASiLWjrkSFRlCC7FHNoXfDZiuvcyHvnHmV371Cyj8Jj/
60AIwpB1PaC4Vc9KVUgo1wv8QXfXomfPJ+1g9w3CvzNyx/6nAsmLDY4A8w6P4VyP
5Quze5HbI2elfp4+h0aaZXh1nCqTCTjPw3pKHX8si+HRifl02TQAIBJP/XjhMkHm
gy11HkZA+CkOjjH5CJ4jPmMrm851wvVvdYTzqHr6aL1iWhb6ltve9T9OEHXbXNS4
ey4KGPNQ6/HINznxWAUOznNxz6g2oDK23/DWG1I6+zPgmUtWo5gmYoyzI1wb3oke
gvgmnwA2qmmh+PY1GeFL1c6IRdv7gygEwEV2s/+OMxFhkE/bfmumLuV4EpbxMw9d
QG1Ixevu2m3F7AAaiuwFXOVc67h7UCVAqr3Z9J6re0PjgatwruDVBoo3hSFpdNkg
FkDzxU6NUqJvDFgIXrtCHehPcad5WQeSA7w0JDWVIgR2FeFD/CI+C/EeQ6Eo3En3
OCG/+kbIeE9Ai72VBs+TJGuoZ0m0tBkGwnZPVxTjpc2ELy+Dy32FwPjNL7FoYKRK
CcTNVVJOCI44zVgUgu2XZs56dv7WKJZa/XP3gL81vQ1SQYcs175q9rq+d8a3Gq8q
G2hOkMGFKPguVpu6EGggZUT73AuEs3KjSl4sK7p+wgbH+mozSeszNNBWS2dZYG7Q
3EhjiqAdx/CZUg7ukZ4stKNa+fPAI9MxirUnXWDc//Mav4Ttpz2JceNq5CE8rRLU
YPjBamk+EH7dapPhBr5moeowAjejQ3LaoFZEW37ec1oc1g2d0ip2INmZPwCr9nL1
nR5LovCSnic770o/iA3TFwK+UMIZLEbXtlZRPNDor/612tFPm/7IVvmaaQz02Ro5
6Hzcm3Oux69Jo6+k/evTp6xZi9uejYS1w39DjJTYVrKgQyqfgkTDgy1MSxtHTcKc
QMJRmeYNT2v8flWlslTGHijolVSHCCx7PUoq98FGCU3QngjBbg3zQuEcvrwiQPJ8
fYCraxWN7Zwwcbc5HNCpffLRu9sthyi5uqbppnGbukge8r3z5NnBMvliKlkX+y8o
kYnY0ytsOGCGahA/uAnx5O5vFqbLxx23CL2qZCXCBXYPmmfATPvjFTgO9HAQBh3p
fyx8xfcxRIUgONgeS1IC/xgK0sle7P6zJPVqGWCCPheZxDOCTzZsQMC2meNIoABO
Q36qkEiTTbI4CRbRma5EhY3yINQdqwcDpebllYvrL9kKJXBoecL9+M5r9LybZir0
Pl0SVh9+pVoQGTdz5rjEicKw0nO8eMv7loM57/03yrCNQOl75p/5fMaStMhiKipV
WKeNDxya6zLtLXTqvECzgLCGkImUoONWbxzeqeLIxKNq31OFEYLKuQBHi/OIeYuf
RMexeM8PnAqM63+zsMtj3mz9hQcOAJepdV5bmn94PuT8ZE5ivytcy9IUP702bvVy
okUM/x3l2/kPkhaR6dQCqyq6q8sfnY6xd4nTpiWXbR565MkMuyepY86Hr5wFb6sK
GBMEJuw2cyssld8PIZ0wH6g7xIyCbFvrgXpLC+0MlPrp8JgH8rZZWQDQCGwX8bMq
e5Nmj3rHTiemMceNfQTXd2RFKzYJii/ps14JVToJy4zfoyWoJk0xRaqNxj4uKCzo
U7TEWAJ89BQjZ2GI1bmX+7xKeykmdmZvaB4zMZ3HU0F8QaDtt4B6faGrRx6ZBenu
WWMBsK1FOYmBHUp+zm92jfzQUg8adQHzB/5r0F5gmWv7kS500YNIlaZnZ+13JF33
iBzF+D+74+cTglsr2d293ur0D6P/8kfJaZ4rpxZv/i70aJA8NuIJ5FSYA+Cka+T+
5AzZK3cD/XbQ0qB38A4RsQ7q3EnVOnhFItKWXEmXLTGNgey86ur6MOamZ1nxkkRI
fPtSO1aIKnu/RifBKf4r2sOE85Uxv/pO59Ip02CBNgYKJSLd037zGPRRaH3EzCNI
wCpCKbzLybjuLrJXK4ElwAyU6xIopfV7BTeB+yy9d+h4GzSknewiiRKxVykcGz1d
vCzsJFukAsWkpRcYsVLPFcRuQESlclq/c/XRKKHW1/UqBFIKQMk24NZZDcgWBEkJ
B8nMfl0WlyD4mUsCxsfgVizof7XyzMDMRaF/j1NLxWROS3/nrlsiFycSNMpdnQU4
MOKPTollcvm/QBC8vs1xakBZ0TGTHrT3Tka3Thujt37Beo4rgHnSod6vqcTF681f
NivQcPyIZI20jcScWyhMRCXUxvu53dXA5nzUnNTM6KBROJQatvKBqTlWJnl44sbg
X55dsA9r0WLhuY5++UadupARu1bpua2hboY2/IefQJ4rfoN70imhYJyeoKs+TQtt
VK3wkRmg9PkRPREtGTyvdOOgOpdS823ZSblbKwOlXLe1ixfVcOuKnS8CltHn+pSg
c15N6i7z6laAmr9RvIGRUtQSIE5v8uKo9zJppFy/JdYzjMxweSP0kFk3JMV+PcaX
tKr2wFwtVD2GvYEg+1QbsFZozOrDyKl+FnfKQtF+9i2U7J1aLiL1tbTu4kyoIo4z
Lzice5gowtHNIkbk+wROZ2Fwh3Nblt1+/hnePJtroXUCnMFqr3pBuMoFDjGQXk7u
aEn5eipUGIcbOIPHAzRmSdxCrItZdjGHRtboE7r/o4ZF62Ibb4qLujNerRasi5dc
5CPxkKGn+jmvbUmj4e8/2WwdvpT5eB/sA7vhjQF5dazmK8hzUa2jH5LZft+xx/m9
CEmzz2JFQ8ayaQGUxnIoEGXFB7jf/p9SsTNGqA7QG0JiKISkMevhsTNUML442b7G
dmOzp2zxbJ8qJ7zdtB2SPIEifJSxs5aCvqIEmFnbYvQRDEGxQTeEumx58qneBFPh
VtOMRqEsueZ9QQLV7ZAwJwC4eqQ8S4t6J9Y5ZVYZlqF8tXOnk/6cBn/SV5aLPSDS
bz/Ode2CcgjHDjauyxcjf11oE3vv5dsED1wasJHkhS0Or5ORs4cTNS5pELr0y62z
U3QMKMgS4N0TFYpQxZ4L4fSHqATefcEha4yvhR68XxzHJqTDvuRg6epxmCPWStBv
clwFlevh8rrmUtmFkcNi6WzZCun4dmsdYynvD927v5ay43j0Cvqzhm+5qJVezWl4
51KrQbVeEGAKv5CZ1vWquUdGizutc4ywXHfW+1gW209vdpiMqE+pJVhEDWy3Tsvv
ZuJZ7WrM6wBvgmOte/maqJmgoZwBkGKypytHXtIr4XvzOfLbzBW7cBWUM+B3r19D
BgUBYCnJnHe0jBxc4hgfqbuWKLxlA3FEUtzxj06COAvEey5YMlD77yp/UWYY6YJc
KJzmB2VRG8C3yUFLPY0Y5ln0PZG2l0RnAMNXSYEXzouxLAaTvvMRrcqhu+r787lG
V6uaDsmG8+qLvNTI85XI5PFN88G7SFrAqgxRYxHc/vfSn2/wq6LvIjhLapwfb3id
7wJb8q/N2eoLjOY+ezd7Kbb/pLsuwT5HZku8JOgj/bWhuRN8VUyzdhLltiTdwzVq
7Gca8q1KGbaNMg99NrfISC7mwKm8KK4ecA40Z5FcNhi3/bLXi0kYQ3tj8m1kiFY2
6FhKp0ASLF6tIBk4o/SVI04wtUfND4duk+ywS+pUrNV/5Nd+c6jr6JtF36WC+oyx
56N2Tmn4KShy3/QwaRUqBhpJKqy0pQq2PRDwqlqIfgZpaIyIyKFtA4Er7sWjduwu
dvgm77fUJQ6TrkMfiJkZajwJ1P5isVLLSJ7LxKPdGn35j1NMvXuYUMqTwPKxDQ4y
jFu44eIQEyX9maHsx13V71OowitnzhzFqaBWVxEPgKyP3NRqA9KSf22ck5oewoUN
4un0m6nJoJRJj8PO2tiyICIifWAmImMR/a0rBEH34g1Rs8YF0yj/J94mq5UBSkxZ
9cIZfzJ0L/tMoX5rvKFqKQYvTUHb/VxPIz1lAxY3pO7XRF1GZQymcYw6kFLc4NzP
/WCUREKqx2wguHRX8MeRHgWFozl1dKtRdCfYynzruLT6YZhbuIaDblZ+2URzyiAh
sGFmy0r/6wFmPc8BSQZkK3WD4PMXuviDtod48W2SAptdCI8bF6eO2PbAzlO9o2Qo
nSd0BYegU0aC81/sifFBtpZxfNb8ciDDAemggKuQHI15lrmEKWjH58d7P4kjp6DL
m9ZyR8JSj0mUoJDF1hnwzys+lIcpfpRtHlQyUVDGH2V/MhnxS0mIPjkLgOVkYXvL
nrsMJo2CHy45M5qnLOibruEdyp5QhD8Uq0rY9DfjWHmb17EhMjxW95534X87PLLS
PY/le8D7MEYIgCaIerXhxDb4tcqnU10pAv2Akl2E5g0y24MnQTUG8Hb90cOYPZKE
+TeaxEV7CZV5tRhCHN0hhRrYVpZldbcbV7f7/QtybW7p2USMHaBRfHim23w56fU9
cHjFLTpgjcFx1lmojbuUrDcHqmbIsJYaG56pTgKBs+aG8PAK+n6JLQpX1RFElAx3
jppFjNMFyfKy4ZEYRbDMZBnB24TAzU0mBeCFJ6bTwBjwisLH1t/xismDzx+D4iZl
+ZJPfqhKb267G5zkdXiZzMkY/Z3xbJf6k7BY43AbF7nVhfJjgB6Z5LuPCpbcVobw
W5RPHb5U2Rh6yu1XklsDeVhtGYr6dZpnVbcQlmv70GX3NzxiVGwUt/OGwIGVPE1L
YMUztHnCs3P38tS1xvEUQs6q9gCR4YGwnWnNdgaDvaSjrdAecPgT94AvDYkuqxMz
xma+AWkdlrxUoex9DD/lWVGWcYHQH4afl6xAp7NjtPo8ObWo2DocB6UfOWESmoVf
p5FgIcrDge9oyqmvWgmQ+wCF7x8KIU5NX1sXvuDeDUZOdDpE5MSpfSoQSwvraC2e
Zy/HYZ29mL70mMK8jy9Ula9QiED1xrCm0i5WJONVV4dyVv6bstD4XoSjcfhOEQUz
USwMNTiQRyLtFMLr/XpVrTzxY9zL4656AFuDEKLbl+j6GsBIUys3g9O9mUIKQG//
PeSNKVZ2pd2QBv5a1yjs4bW7rnuGaGbe6WPKIIK7EKgQUScS+Jzf/wVkdHmivn2k
mfIJnjrY+1VtBJ3a6Pv9HLJ5xD/wlJPjn6LGzEaneDJmaFkqRpIr2YtJ4mMLUoct
gx8rXOpDBszt27vAZWxhmKPSPyCC1VxvjL14l5UwpmX2tu/4JFWipB2KRLA2O11J
C8Moz/f5+86dApyMxi+HyL4bYeQjMjfC1HRAqw4K83d1yxVz3H8om0pcSpvmS4jR
SQzNfqzQji0sSh7v4LyTEz97b938KZpZdfP4es/cDvhu5p7SyeEbkcHvpFezX1XT
KSNIMNbBSBuB1kbOwIB+8P8u8ulQ/5Q30HNR84OK2AK4Zznkem9d93flSgHsoTjy
oVEJpUyLkrPR2icLvsvQS8QYMRL8vGxgM6S8pwdVF35RfcK02rVe78OI39RKYFun
1IMCzlIQgLjENDWEFNJI/mBFXP269y7u8Ovzap+1lD+8GML6Dcpa2tD2azR8FcMT
qZ8toJIXlNJz77AxSW56fWAa0eIorY4sGgrcX5AkcNbAh5Aerx+2SWyEHb3uv1ea
eSSPFjBRY9rkrjqM8qMbQjnGB3jH2TatOHWEHQcezXoOZduVy2mSCGrO+9DRakBf
ZMD0QjYpT+URpwNUafWkFxS/yCjLcjYvkFbPAFwLPMH6JYJQz+ewwCafk635y87s
OFncTwRlC0YoAgakYDxqblQSVLOhjnq/O1iLS2SANvO/c3HWOdtrY8NEAipLuBQ4
cTEJyIQQP9zHJX1ePlyNB0CeICXDX6ZaIX+iehtUxgrW0gLrDbOk7sQFI8GKV0zB
8ptyf8oKQmRi9F02coOrAb/ssKKHyNc0UemAldhDbO05TPfZByCiZ/CigUML8bVR
d6hvR9eCd/8inc8LHf23kDAyPexIuWp0R5ehO8xMBWFAs0+d9uu1oMRJqziJwsK6
DLTqF4cBaa30onRxnKVVjj/9WUQdpYelV9npucaLasT2MxQ3vL32TqH/nMNje9Rt
p5jnEjmf1MaMQHzGSqFoQaKmc4OC8Gh6lfNBBBo87ljpz0c6nok+RRO3EE38LjUy
/PTGHjXFA76UFAoWnAUE1OtNdejHtadc1bU2P/CjMWjjVsa838LEYoU1sxoVbdml
9uoYMyhxTPiFBSibYlfBOpMCEXEUz5SyKZUWAALuamEHSRHIhISLjK/hk+N9inQJ
98MYXkoj8xh3rT6DEv9HVqowJWKU1WwtN4IaP1KSGrlXqarNRNJXF4/yURwsdVfM
gQ7A+SIV2zjXTQjuJ9Pe6yrJc+sCKwWLmFS5QniJbu9tmBHRngOsdcecTZYviBPX
whyxUD+FAkyLrFosdhb019bIVoYL6gNp6hucby0juxTbCg0lrM9zS6iYVZBC5cxb
5VJ75dc2FBGUalf/N242GOEBQOiXzWgxYZ2hdklCcNoM1j6D8e6+xVXj99JgICun
f1SsOe/CzFiXJrO8fZGbp5pE7bkQC0qUCgENCUXiF371/EV0rszcBk3OWDr1FNS5
wk4fWCSeGkD348U0KoJSzZdaZVa+q4e88QDDU7vNYR2GgexfFCdYA+8B1NU0/MqO
WqhVC5mUF6yHQtSh5xgqu8oM2y6dR34qA0O0xpJWPL848ScJFoUma2K4Fp4d23fa
S6Pb3XsLZ93F0XgrScq7Z/Kf7HIb6550uV1HvtVcPbncsqiR+QwLNbnhoWmChFh9
qVdBBd0AjrTZ5ewBPlin//sCwFi/j5laBX95LbAYaD/ASx9u5hSy3TjnMs8ZagG9
eMGdQQrjCIjn0+Ophg6SVcZUlGb1vsHKFe8bKztxyW7DtXENTdgJay39RZ6XNIxc
mO7j3jqstvXrETDyKaAV02gAqR+uvhX7yDmNAUCHUszFBkmum8Wu3YtBkJ0U6iZf
NGPprhwexL6lT8DGek1WPQcqtlcOkyBqs+eX5WEtN/4T+hOzuZ+i2mEYmx1CREqN
q+A17TGWTGpz72deJQZrqNwGsjQSydtBZPv/9l7ojWIh7uxAM0WSJauQa+CqPOfY
B+Bn0xrqdWHgXJu9Ro8CAtO9U4+cBPo07+RkutHSz9WtdpkQHjWjPWd5mTrLIT+8
ZNJPZqMSJdSTlpBQeKNPMbAn0CmteW1oMRNX1tZbfjDOqVKfzLjqFnd/z9hG9XGl
JblUrDOjdOEnM/OQoEsYjwUnzoI1KqBXc60vAkxNhor99m+AP4OM5tilwWEMU05S
kGj+Qo7FrOpth/2bsK+GMn6yl+a6N6GotpNKVhhKqamM/krzcZL9YWJoua1YXEk+
5BddNhT8cVUADwQ07hGVZNxyevjcbOLtMR9jTeLRoEkGcVRd12zDNVFoyR1w/30c
0vu7ceP9JYdTU+R6Xka4+Uo0wZLXgi5FlvRbb5zuWEoL44T4EaCGVA4xx6BxskAX
skx49OYuRBplA/Bz89+lVlEUN3ggp8tGFzTREBbBWMRvTNF0osV7MGCC6CcRY5ha
qcxtu7+wSWNni+ES+bxps5jMypPtTwNJLKvSPLABDS2PJ6Mr9NuVFd3Wb9hrdcJB
Kxt+CB/iD9jel84YSoooez1xDk8jT3bNk49cW4wWizWCA9DbAtMEz2WcAAa1Csx0
JkiWMK09VYLaZnMlVZ6HTYaAVbB5t9I1wCYhsrBDP0+6DFmmG0fkpYRIZorGwOVt
I4OaUb/ooelSurmv4T9dfT2qvTUUIv5g+KRYFMe4724obTgMg+4bVwa2EyDSSgqq
XAx6jeQKW5NvZs/57oHFak4rwpeNdAFCGfWmtjhC5KAv78c9a2NrFr8OI+q2y/7m
qPdNs3zNWc2KFPcu7kEip5t4F1MKSC7lDoxGP/4cXfIN1rTKgVNB5NBWxP0GhsEL
v6H9jYPFuvZfGcdf12W1d/0pvRUzl2EdY51WkfyRoMf2ForfqQYXwfudvfiKeMBz
gtj06I2400Zk+sMwuHDv3dW9OvtHzai5fBveXeXhu4dxfXQHGsSkFd8OXlCLjtRL
UOWoJFA7okJUCj7YO18PJ/g7YS7POy+JwL+KLTjz+P2eJZzPQunUpGBQJ9bFGB0A
XOzsA7Blat862pKuNsqKAJSEjv2gcu7JzJhEWeaF4WvxnlxQ1Ex5gX8GvQIlFq8o
WhUC8yrBcFrD7kf9U9iAU7aV4QHzSqUUopFRU2ASzW4wEhf+/fKJcPXscu3GGmzC
ZdtrLtZ3xMrVr/ASpI0K4zcO/mrdb9h0dAmWpYwKu15bIxkN1K+1MiuYQa0PyezJ
JTX981uhNghTIP8HB3rqImAUYw6D8MK2nhcgdwKAw/pnfo0C7Bgto8LNaphvCaJx
8Fe56/pApmaQMp+KPUWu/4vIz7NJumanFKUglB705mwpOeQFWnWncF22joNxOjCo
Wk3Jop3YJ6s0RATOjzrz9KGS7NMGH3MQuRSlls2/McNMTV8FNFmiPzg9XbHPPh4e
UPuFxT/oqvFYsHEx4Xj+N7azdO8eVj+keKjB3wxW7TSplxFrmK/rR+IQvwSV7n+z
Bx0utZIXEuYjArFEGWWSZ5fIr1G0AGDTcTTOCqzIPUY0xOSDxZRMNHbX0Ew7b2Fh
KXcm9DOAw4M5xI03q2T+DnTC/VEfCZ4VGLubJDPOcj2O5DkXl6JfN4/EQFlnkpLt
OLmTlwVO+JUCUUVA9H7WdMKz5bJv46tFxEFOcpJzknLoX3kBa473RCXDy93AjTp0
nbbNjJKRc2uiSgUEQYC4YKXp9fQIGf20kPH0X0kNKUx+cR7wqMi9v+rYYC4L1cfl
51R91d91bV/nl83XNUcbnPyZiaXR7UWJ+XagZbUBrmCgZ+rtpaYBwIgULnRGq3X9
cSgHgh1TaZuFo+2RhaJ5qHgMy0mAR1wSFkTqjhijg2p7LBkK2vPsOzFESdBdo0TO
Ot+/TytMEQY5ysUKB8As+shJUyhtwJq0BK/mgs/jKctBGZ/fGa7hHP/LtaRVBwEM
F7UKdjVrhf0QgJBJ51bVXBFm/3RugT9xhZi7+9XmAFdVTFrUmgTwpl+eRttZzbHM
37XtJ2to1gBhLg1yem8qanrV/Fo7eRe5rqMp5bGYbZbVT6nxYDpkvevUEPWZSpNs
vp+gnS5awwFlCbANrmERsL9dCwkDK4Joic2KAaD+bZB88KDctEvmr/u8hG+3T7U8
PARSM8b2ooAiUclFIUHvcoO4EJcfN4u94uQa9I1GvOf3TJ9lTBZe/SxKM+3H4mDk
zyzl2ki5Q6dTmmtEDjJ4afe2E1P/OEGF6tqgR7Cz6Y7Qyt9JdabjZnF7h1qw00co
1UeJmP0cEN6pXmQN0XfBsObpOpa6ijUNDDK6i3WkWpcDsdPL5YIorL67uC5FztoN
Uw1wp34QhlowiLXpUkjV5f9FqVFmpKZepxDVGuzyVH0lIqT2CiqcgxTpJsaxZmgy
PBwX5csIsBxy0DhB35ztBYeG9rxHpd6aviIOYJ7KDgr5v7FElzbSCk9QM5JtozID
SAzCVYaZ2iyZYD33uw/EyH+lEpSLCIucF2j2UH9aXQYJyv7/MCu1V/NzW9H3SCKg
LhcEzMh3lfYyPv8cTrMfdF4l9jTBVsCNV8aiVSFi889M8LLhIQNN3BoPq7AiN5p+
UsWc0JwFX5jogKnUTSucDs8bh7O9lXL1V80/OY2VH1Y7hyCWGSwSdUzjdtwb1lt+
PcCrIsup0IPH7UEw3PnDy3lZBn6OIpGO0PU0zSSZmXvrT8I+oiHq6aM+PJVNMnej
PtM8oopvamMstzmwIRQPAXCYre0q0RP1Wxo8Eb/s8/8KdIJOMfB2061BptTFk262
PR4WXdlmwENkDycill6/pOY8vla5GKNj7q+ouxC+uwN3FLInL5cnG4RwGhOkc4vP
4CBaTcHQGe75vNdTzvThcB31jxY5tw0rhhxGVmv7Y/hFSBExr1pQ/z3yoF6N9RLs
t2xbRQzeZMjWwP/Obh2zHVwvmGg5a42OuRc/FipJMs3v8+PzKZnx3F9WgOIJnVYO
gNk9ZxiShufcVOkNLlWk9PnAGfy4mqMl8APn/SsCU1IWTAyrCD93f6wMgpyYf3H4
74iARNQwvaoomSk2pkDJnEHpaa22EXglKfndSj5iYRS+YmhPt39ztmNdBYR/dfyx
o2XbJwv/yq1NqrLw16Q1b1BWl/JwOUHqQC8Mk7lobqMmpEO4llWdUf3juNFGlhI+
7b2mtKIaJLSAzFOtxAYhh19t1L5WdSNBK2wO3MrBWhrb+FxM5yjOtbBMK0d5cats
7NRJK1olGGmwzZzlLK3W1+KJtLWw/XxP4VkzkklsAK2X/ZRNGrjrjEfk8csrSJdZ
zNcwliR0bivCOcvjfXRl+hj18Rh6PXOLWWu1kIw82pvEaWQjo07V5JXKWTZSiukz
NHS6jxZ8EgrnJLBwWEmRkJWx/hEJiVwiBDIjwEm/aRbflrPKw22D+mhfnnsYnMIG
K9VwkeuGleZrNXNzvpVAKvh+GDDL5u7UWMV7HWczNjkQKpUDQnv0mbCtf9htcIek
MefxmC4tpjJP+9ekgPZ0dpPhCe1udeRJ5TbZKrihB+hJYYyC90RFc1L3fdG+NiRq
A/05FaV65ZCMYn+IuYfbMDgNQdwfq3oGvHaDCx6ql38LBvTG3He3jdtcn5jdDNFl
s3jc42WXaLtybQZGCjNFHfkXtoExm55G18cST7CDarSMom+241NFoTaz16mhVE0i
ND/CnFgmFDuCiVlB3jiS+yFh0CtjccaB6zRxV0BHflHFGU/oCRpHnUiIHmdaDlv2
q6lQvrBhf7r4dmxx8ULBFKivGN4IDunwx8rocUrORQgqHiyEtgYvdEFLQNqFCRvM
gFMTwHJnrLcqZg4gfygv76o8f4vk0+2eDnETkDB5NgekTJ7p+BbA7bHQFhutWduY
LnklfCqBKODAw69vXA+tvsd19alKrC/u6cRZeuc7tvnwwLThQAg0DxZVUsOWDymg
CJa+zTPgIrdTrvLoRWERlemsABnDRG4G0OmQou9JD8GbJSgkW7F7xC7OkUk3eYeY
bEvYdd2g81NTLCgp4Xnd8nrLP7qBmiETESvFUb2k1Ujuw/BvUxH5Z70YrGbzVBUt
tqtSrZzrHCIxGvH8Y6LNwxUkWbEz35JZVJF6yKOqElR8yWCBpz49yQyRQxrPrr4n
13pzRHm3TQQ5LAnR1n121BoRfP78uTdA5Sn04w6mr2ztXOE670w4nWPe6efZ2W2K
DQ8CpnFyN8Ptwmx2EZ3/csEniWTf67bWCPWDaZckjSTuU+YGBjJ5sf1mILP8NXVb
Mz6kWUZtsXmGFlPCk08yPqg79d3K85ZhYQmUIBPsZpu9ULIpWBEOAnpVgO9e7Nm6
4+3uFvF3BI57hLrp17Ha1VMLN4B2aERB+q23sIu6ZyF1OovnQvSdw5N72x6nI5cn
S+81lQ4/BZxGkuuf/NE9zzzf4UpTCUjibHnu2d46fOXnoIGfPmPy0wmiWdXxVK3t
4T9WdTs2YI73bsZ1WdmbVhFrPATK9YLYAtw0CbRjtJ4p3bg29GgRRz+sQTFnabMH
y9vPO28edqVpwX7S980KScrBXrRZ4ue77y2E5//85aKTdQDb4jo6PlnIYETQoQkk
FJMhIGy4wWNEfOYzvssX4LdUpFLmQxvr2gGNr6PmT2Ahx+VrFqEazWjlHtKbsJFS
X1RX9HTznyONH3zzmAuNbfQQ6WjUvvKw0n6tTVZtwBU1xp5d+qRNK99iXAmSoKVe
xu+YP2y80nft5jfQfDu0cMFyO+O14miqu9ylvhlMfEuBfwPCemO02JeXzYLOqt7q
n6nNljeNwYdShxuKG9iZejcD7WKY8fr9bvNNgOSiO1mPMdUOvooTJlYrX/SXpCrn
YJAuYtvOnR2Rwr1Z9p1jJyDVDqWsZ2+Q3S0bSjNyMiV91tRs9WyPDYAHMw3NLzy3
e3G3Zt1xfxxJ8vlFg0VIY7xL6R6zzkrtLvASCuiOzluxP+m7PjicjjWn4NsrMXPx
HXhfPiWEmPunI6dI9y9+DrJZk5w6nmxA21Clf6I4jO0QCsqmg8qHipJVWQ+04hf7
pK3j/FcEpCHdEgQ4OTwmmZH2VelZTS1elgeUSM/M1XN+OKIasHZ3yk0kje3XgDKP
nRAz/igvU555Rv0+rH9/S/Q7V6J6y2eqbXGXKrOX06aoXsWvNiSSjpCPaz12bUTe
vGt1j5jkaFBUEEEPDniI8OUEvdgJnpVPppCMgaE4DbHW5wgAPPldmVQVGGchiVvV
fKtH4GWAEbqMe+ix5QHzIx4Pk5bKmmKt6GhbAYw7qjZIzpWqsFnVSD3/VuPq4f7Z
Tt3vZby73UvA20j4rUJdLd1qpINQbzmp/7Y3f9suPdNUGooRA8RhwootnR1AAPrc
vVxpclWBdVgZkGnRiHr4XHDBQ4ENv5jDKS44BXjSb8VjzBvTmxB+eFKEbkljkHnP
GJAQgQcRW8juY+rCVsz4ajHQ/n5ABPLpXyWipKOL1C3eK3WOULEIFqYRAoFfuDj5
nfmUa7c8Eqo+dH3MZOP2SlK7Wf8a2OEbkwaOykWr0J22KSQyJ4OdoSDYH1JTwa3P
QjgpQpu2pD84xWdor5Y3QGOspsMt6bys1HuMYCLqcIYi4sYHz9TQ9unitNaC4p0l
ByTQYRwctps7ymb9KKOazCNAgmwnbimtS9adi1ku3NQsba8RpUHythP4Bmt3t6ON
O7Nc+kuLqFKqJlZMbr9hirpjmorWHbZ+3fACKVzymp3zj6pwF6PTragMo8c84vei
GpJ5kIP65whZiaNVqbBwjxUnyU5lR71lCkX05O48n5EhBue123iRQG9XQNRzN3So
24Ym7suY99bUzY1ycDDBDxysqj9G1TH4S3sVA72tVbSiiFseClYGTXnwJUfPSYHr
ZK03F6E9jf3j4Cb/2oDMYgmDccHouPqCmhEJCJCUy8yemzLwqXDW8xW6YabNhNB7
SC4NAq5QFAPv0PM9zyQSc7xuxTJ3cPrU8rYo+czsPLBm2gDQVJ3mcjrAewSapcj2
MQ3/kg2Mbqve1Da7X1tjj7eNlU94Zm0jfYiKNQsUtJmNbaL/XQHHJNnUguykyk4+
1GbgPzv5Iu7/xdGB2DhKEbMY5gTVrd14v1oXRGiBorveKHnsomYWeqv6LjhJApMM
xYLqwES0XfjdeSBSvcFiEIRxXOuU4jODbrqaRdA9rF+4GyEsZFl/AB/UJgHi6mIN
7uZGcnCGwaU+DhnY1CPyZ7rslJBUikA9BBX96zbETRWdIFr7bzYnP3ebVWUK+wUF
y9piqKpmXnckBAoVPB0Hy6fp9ZKiGDARkYSrRZulxOns5lLgugIhKruJlRGX+BA1
cRlUf5wTs2CAK4ilS4YBfJCYJMm0AHrEmM6lx1+5b3GXMVPz4De+MEzLGiF/Y0EA
cG0WUwGEHwL3IVrpJLcJ3CkjX6BWzRRif0ACZC2UcbwppWbgBlaadJwlQ/OUcYs7
pggV5V9fzW+L2U5JWGsDWJ1Vt/xQBtFjgTo00ZR8myLVrvTWvyenM3OliMlNLOXL
H8t0REUFcA7fTXnYDCN2Yn54+XTRPLAOo/8fdor2QYU5VL3gF5mBKj8hd5AZsAOS
Tsu3B+1fnFiC+gRaAfIkviFx3CtjiRbHnSNvDL8QZkaMiBpT66d89Q/lbrW0p0jM
V4l7r/gsf1Ubd5kObC8cXMrqQrgsEfZ6Zvcq6qJMnMYR8rGAo+URJl7MWZ/tTiOr
guBMFNmTQihU49kmt8RYDtABjhbrU4MYrJe3djKkEvSoOVgLztrXzeTOVUk8mWCO
cOp38oCih22NWaLxKZPbJGopFmrTgeP3u9SbphZqXKDxlHW58q2nnjx/U0O4l/eF
h4iHXGvwlkfx0nLm3Ky74Na/5A08b84fQtwGL1tm8ZtVMY6sXTrg0y5y3T6N/93J
jemsaIfA/k5w/CR7T3PMRAr3/+OqsvoZd7w0DQhPaKoMSeXxP5DjcCl0HKK9w4OG
22BkHPG2jW5mE19TNbEtsXodZMRuGywOJLAGTNNSonVN1rpMT3BVm5w9NDInUenw
IEOdm7bPJAulbgttM7GmTykvyi/LOzaLVeqNjxly4kiQSp/wkfBkCxOQTLOuILi3
mtBBLt6l7i1IEgxhDGRsRvex3mGkfsLg3KZ/ZMPo2QqEeDnJ0eiMAqA1hRGxs9uU
hVUkZYpmRpO7rm0/Sb41tMBKZbYoSr2fvMYx628DjJFYL8x2WM6orPcFXeKdEUCF
UTGj5JUqJiUI+4RptWfu6cIVIDzg7Aa/Rz897VIAbadlnTaEX7y0ipjz+SdOQGR6
sBLQGi34HnvN2e24tI3RHskFd6aXnO+22QNl8QECj80lTsnAUto03DsSzH8bcqFx
QcabMjT/B5lfjckDuAyTOOE4LuXvtW8wm1D8Js4+8tNXE2bfJhT1R//1CQccbEdt
HsqcxfuJM8Ue6d6tDp3UQe9Y9j50g0GmiaIdOvOYJ60rZYra9QpRreyT460A0lM0
DkEJ5u723w3LabaQGAx7qkTr9oErzmlUMeZivgfCsh0r9ZdT9aFXGPCAp81KF79S
GlJZA2cSYzC/bZfQLW6L66zBQfxxgRXPZDvwYvkCV1TFkWfDycPYH5eHXoUj3Tzn
qm3vlAZfCfZE04WMEbpMyHLCXa67RpPdhhCJZNvVypbAUv45r6Nae4jLrN2wraRz
bmLnGsew1odI6OKSzfagr2phxZiRvoz9jHahl/+51EjMkB1Kalvva4hZTQTRlfsX
ahq2RxHGLbwXzKM8Sd9z2G/DfLtEs0Y+RAu7WM4jfclzYFkVgCohk90mUzejMd5f
i6fFZv+vqeWHGJRodHPpr8y4SyYp15pRNtqZVSp8cH0MP+hp2Cj+9xPxCGyNhtw2
wOl1IGnFHFQ/DiDP1W8I5IG5187gBNE3jlOrWLR3NFjHJYMmWtZ8JrPNZrhTu75G
dMD+3xNG1jygAdICB+ovsohNYAlP5VC33dJ52l9cIYgexyi7teIZ5I6bhgJjZ3WM
XMwqBQFd1oHAlkce8o1kF8+jfAGbwjRCoiNGlQdh9+NABSAvLy4JT64yry0Zc1CJ
v7Ttg9AQqPuvdJO1huKU4xKh15i+J0NHWLIMokIbhdokCS7sXymR9HGg0m6l88Xs
+KGDGy3hgRjgWg84/kJGC6CRnvGVfbDkzY72HrMvs5N2uv4k66h12KBlnEOj7i0b
6gLFB3yD8eE3tCYC8767BfoqBZCeNdtgsffmLKmgnUULRQkabvbGdSGAor03VvU1
VdKPiXW4lL6PW8dpB9FueojzycVdfbonNtm7z4KmP6WOebpN8uGLnVWK4MbxsMrU
O0TEQRyoZx+OkwOCty3SOawXr+HY2NG4o3u8NDEamvNE4pHlBiKT3eVcMoyerx+e
6l+pHOrIFdY1ZfC46oKZYxCL4Iu/cHgs7YMW17mRc9TESVji5dzcMdsT8PWk9ZmH
EEQGe2Lc1aTsfUyTypW6FHQJec//mwAwgPCpANw+RxyfzkGaXbNP+9+tT86Hlvj/
0jLPIoghmPVNZU2tIZkSolwOm+gbl7BbNwMhKsWJ+fh+i8fJV67qsnTiRky6z/kj
Gm3500RYQz5KM3OJ41WCA7h3INPJXb9uwkMmS3hMBpTAsAiB43G30baWmpVBpbcm
9nPm1G6d4vCeYZK/LcVNkK0+InJDA8hZoHZcJHkrSCprzD6EmG2KZJLYVbM4U0K3
Bu6Wz790nfaIoqN2BfEhfIaMySyJ+uAguCCOD9/E1vY6VSqR3cxu5LBLXjrxYQ2v
ObxDyWYMyf+dgUdCVXCtu+RPiJBflDSAg2yvbTK7eUo/2rP9IKcbv9mUXyvNWipr
oloBfLs4bOjnLlBIAY8aefSZnGHvXP2CZ7VRCT6r3aEx/BSg1/mzzEDM3rpI/w1k
s+UfaFcVN22bFi8vfRio9QvhTh31ZGx2p27P2PkAMaTqipRRg9OnYLCa36DeXxRj
qKJVy0g53j2GVkgbqMvuXrUzjqwbfu79Qu94zGR8MpuQjDVYjeS7uVDwq1r0trUA
WF4Uu+yWQlyuh/zFJklYkZZwKXPUyENlYxmvpOmlo1frSPq6QFgSvwE7qxwQxYYP
0Q3rbA8dPaz3BINIGb/rCRhMXKlZcrq5VHVkIohMq48OZrB+IO3V6xIJOezyQi5R
jPOwwURozeZ5LbYYV9X4jGVQQcBhuCZr5+Jg+aRtM6kLzrpw+pWITurifgEI7/o+
fLUL816eQZXZHfYPj/bD/lnhygpn/7L4be/sWLEX3eFLUqGjvT4sgxYyRi59cb+M
Xfd1dDBAQC4t8j8NRVfGxV6zgziDrYV9oQyKItRJldc4VD79WJdYaETSftT9bBGT
XI6d6OdukFdiVONLAt/Y54di8HdMivKxAdXvm/R25fWylY6vXljgfFDrydFN574r
uz+1T2+H6IfiqKT7UJp/GjHcQkwJ5VoeSvD7o8pLbjiAMuXJ7/a+l9m/HYzy78Td
EXcPGKIW7cK6RzQ+jCwtpO1E0PCzwgkU2IhEXehHU1e+wx1WU2AHxXulfwL9Ew6c
wTZMG3UmZ2A3Us22F44uiGqx0aN8UpbGGRx4/gVInvhAWxO75Y40aOhJS8D7prmH
KYbWI2V3v3kLOFAA+dCa3zrpNS1Ky/mXfSnzCk80yub7ySF0DyPOT0KP5GAyrLk0
e3op2jYjHzTIjGOhZLVqsUk9WeM+jh3JDF2GO5eqsnsOfjpHwIyei38erCMHnz1T
WDn4pzjJztSoZE1l+9k014WMfUNuyBqZH8imWynJoMnbj02LdAhAcbfl09aIHmWX
ecwbn4ojosKfuTfAg0GMFHFx/EpNqy/0ChLAWWqO1ZCCB14C3XdIE0V06UwpHL+z
qu8rgRj/HZ35iFRgVYGVYsJ09DSMqSiCQ9AgeLuIfbxKA0C3nUt4hc7Bb86YfQr+
PCHIi5RQldVtH/jdu9vC/wWxsGomyrDtK+zPgIB1J2ABtPkWek1kesj4vC30yrXy
Yw5SHEK30Nzd8UJ38P45G7BvoonnR0Zu0bsMXnQSmNSaIJOZJ3NKnI+I5rZYjtSU
nV4qdXJTFBaweS8UZHBfzekaYWOKi0LOpFqyrtHqJLrOYE8wMnRoXLnDWLgCfyaO
HJkD+erIbAJAvq+vE9C/MDFQytaEjtAVDBX+P3R6w6cOE8ucwUX/hy7Ftki3ew0a
hzx2CvxHgCWtm4agkQi1zCiH1JQ4iaNiGRvhq+pAdGEeCMUmRv0WQOkSyctW9jgD
Sf3esCuBeNF9XVr0HnMHqS4Glu5Hvdbgi5pagyl2AH9PBGjU/jbEm07OgSJtgEYd
2Mto5T2FlRDAM6bRLMt4MXB89maButgxOXufqOSqkJPACLxyA56Y+IG3YR2HjDaY
jGwa0ElfSHR4MoK9Qt9zQxFbA2dF+kPb3jxBnSqM+6VA2s/eefLYHWID+ZVCi/MC
UNd+G+eOmb99W826ESFaxrY2Rq9nYNaLVW0cTTzp0Qql0VF9vZnGOsX4+QF5j/VB
hWxouU7rC9pCFmuzMvJCaccO5UEB3br17lSipaa9PU/bzch2FHykNYlZQsIFitcH
aV2D3bHq8fahMCySgHrQg3RnXhF9yIQIOS4pbwZcLzrxYq7UBg+tImL3vY61JLvy
15TxAytnp3cLaNUeAexlHTcsWR8qKfVR6boURTjPMseGK1h67myZfsDzGOLM+CoD
HY8n0yHobwJ5c7HdjMP9+d7aaAaesnPo709kWnuFH19BfVW7f6/pWQnZCQxrXYMm
uu+q9XtH3qTIq34Y5BdDwKszYxKSaRRZH8QD+a0KRmZINZdu+KEIxdvZAcAcepLI
VpF9jPU4icgnaqW71mURyYm3J8y9B+y9gqn5zV7+buZau6cHW/M6UrjxW5ES1MI2
sE/2nowiQGUrpDdDs9FB5SDnmDH6hhQcSKk7DaKCuAywE6Yco2eoGcAefIZkR0//
Bz5Sh4+1TU6Cp/GFt9Mh/IQ4QmglQyCHxQ4Y9HroU+2i2gQkSA+v1e8NLVIQqyIE
kVlmG9tEmEAyz4PI9h3JP9QRQWRcASE4c6YkstdV3jsPTAgvHIITTEWubChVKmkd
Q7wywNSw27HzmlgeGScoKeXrHEEBeXFdhGRok+hVw223OmJWdRrRyZ7KCbDqYd2T
TI3RxEqcA/gjlvHdbeZK1reIpETVWgVMlFYgWBqzDevy1f0bhnMn0ausvCxtm+Ao
gWRbxb8QZU1wsUidMlt20x/dpFEt6Nvmr+8R2huBuJMxjskVk1QgCHFNKPN8mMMJ
a/P88S5O8hbPTaKC9kmfWmXI2M4ZK5webD8t+aG8r6SXCE8XSLeVIqSaiZHRJBnp
YsLdhL5j86AW08mtndDLh2+8fG206pOLbzze/GJfvf6njWQxr2R7h/XKgAS/viD6
TfOcleVQ1dPa+wX8uBlfO+GYfFHdjxM8P5ZtziPJhvQ0TX5+O7S5w8jJ19+8SXlb
NYdYL5ZSIsUQVLT6ACVJcJMvdAHVNDWrjjFm2Htojx9iM+HJSLPO0LAGnjtma4T3
bz2nFQ5M53YgxZ4LZofwdgCfYXHRA77tdlbJZG+Ps7dkZACZzwzltZ0vqjTpJAdU
2IjYKuNUAVGGA6gj1b3nfFkEOQMaLdwTePqXz1GWbqfAHTXh2eSqGtCFYHD6M63U
E/BO3YrXDx+3DXHF8Wt/4nH4iziydmrDuLHsg2wrmqrmvSJNgjHwHoF+vLF/pimT
Mg44RtnSegbydP7SU3cMqvkJXECbcHHBPDu0ObxWPCJKit8jj1N4vsvryIC6Q3DP
0coiGQvs3dd3VDtiOOsWxGLXd7bD3OQxzADpOj0/ntsQXt/4Aq8Is7H2Xcz/LfDh
OrOC4/bRXAsq0+8gSZwUv4M97pAi1PgnFv0GZYMCAgX+LSiBzW2Eht+XEIVIce8H
FHF15VNGciY+8EtTt1d/0h99FNrh28jyvzuxTAydK1njv21m1RSvbHU3K9y2o2fz
8pk7HWjp+UcWdcyTa55dzzppVWwYC4m/eFiXxa8KCTWMkXetrmpFovrzVFTTeVqf
V6qX8FU+gLnE1Wrqp++a70h+OP2tQxQyUlKFQDdURCAise7cCSWj9AUxhokLZt6W
NzRBIf6G1wwKmGTZs9SNfRIKNhUKK34luM/8iKElNPs537A25OJ60Lkow1P7DmKD
omyC/tBlMzdyB4d1PcwrCIZSqE9KGP0U+kK+gBDZY/9AGzYDp7RYmYJGB4I9R1Al
FLj178w2qbQq1hYSi0I0EIEX8EUbq1nBaox8uA6rdzyTSRAgwbqihoAnOcTWTC4j
PmTnaajP8UqKpR5uFw2JO7RIdTeOY1Lp+uO3x+qnzbGUFuewpPkxScVsdPIJxRRQ
AQB/x4n5tCtArwInYIu9pwUXa8clHBK7TaWTPjHOfWJQbEqq3hI5kWIhKEwPqJ3l
KS6ZkFzsHmUc/g7J97lhvzZaHNDcX4MFU9QG0omKAmd3JUOBSDJio/H6V4gfIAli
TEF6qUARI/uKjEy+UQNlI+NNpUkdIaD8wqHmQVTyhrxOi3LAaHx0oPhZOA3nW8ms
mU3M/vPlyK25m1nhKpLLjTo2szGHmsalBiCjU5JbmD+xsOnp8YECltbdD0sqHotv
+gUUlHNIt/ud8E+wPifLU8YbkBbxXmzbdOFqgQnYRiykgOCMGCEMLLcDVgLbHq2h
dhg4Tlc7FAEx3P48JFIUQ+WXAtZqGYt+6jN+MdwdQHK+fHiAdIveV/8ycYN+flmK
iSva0bHGv9Y9QLXZKYQuGot2odS7YQG7i844K7tC/a7KLT2hyJ85RxlLlfvpjMb7
TjIUoxPYVCcWDa08qB0nybKrkFvKjQNzKJHKpKgT9vklmkgPnkpS2T1InB6KfX0F
/U4tViUIRlPxxNnQOQ8Ptbq0ndn+RJt5PFiaY/MQZglkFtxj3hsIl4F9Imi+9Mr1
SOutbWHFz6qWGCqNmNOFldqVg4wxFzZ6xwEerQqjb5cR8YijTehv+Jt3lbd7rQRs
rKICxsSEZdkVyGMieDfK90GciFRAWwrdVwtLd8Ty6NznW58X1/5RNZ48OgcgAByO
R3ylAcriOXav2j+5tL0ikg2uvfhITDYhXN9sJjwPGXf1nP8v93RyZtQo6rPwujkT
+zS5HPhn0vv8yNdnZAAqgVPllEGF/Svy6umY4Cn03qAQyLIyDG7o3nwqJ+WmZwjm
3iZPJEzOJw9OjrDx7CJY9X/UHliVwlcjyyR1/qVOFVUrFgiyL8AYUSiwKylWHHWI
e8CplY/t50F2tx0kteEZjCS3zvec8ECRoBnqmtD1wfh6TaSvQu4u8/EyOchc/ICj
CvDDVpMtXtxVzmsviZ+eJ3vng5iGGkg/gUb3I7EvVBuXzgZZBxNtJjV2bam7iUyG
SLx9JLaLj7tEN8xONNWsl56lqaMw3xmQdZ8flCTDs5TTlAc2U+prMPkAq6pSR2Rs
QXV74FLMmnAkKP9/qLpZ0jotz76kDAIWgM9H6gkNZZiC+bCdix2SuTZkwzdvUgf9
F6t5gg8FNLmghN5LJPYs4vPcwWt404p4XDtt3XgFYrTUzoWEhvPxgmfvLhe5manN
Tgjo4XnvbwKGVn2xShExT8q0EB2bd7aObJF87TG3SjxYunFCL6dyT98Jy9hwEkim
+jFlSaBsl1fGsXYN5GnL52Dhcchf1m8t41LL6KcUOqws7JSK2IXLxaUclhOx7TP4
Fq86F+hy046QPMNm92+rf9xnlGMqYDfYX0JW7YsvDf5lHUEtSSkM1Z2eFCFY8Hrx
peMDyN8acU7YknqpccD5uiqNI0oMSWREbcnAyr6Og/q6aG7UOEtc5z80DSHmaiyy
V+jg2yWEvSgThoy8PPHnfpgbeU5Y+QnTfXY1YrFw4AvsKeix0yESfyR1vj21YLeV
NmbeVnAOyXnU5g6JkG9uYkTFrQa0maQKfMxZ49e18FF4sFV1WWaP3Wn/IwmTaU+V
lraxX2rormEpKNrdxTrV0nyOs2y71B9qWil0U8e21arstLEG8FFvH0Mmx4Jw2Ajr
JptQIWGwMNN4Cf6yxTTc7pSVnpwKrr5Hou8jdoq8u6WKlHUZA/hxYH4pXWm0Upnx
wJl+CykugYGcbo0wYqOm5x9P+lPYTxDxmQJ1cMXRcf8beQXuUKk+Fz22G/zdsRf+
Pioo4ieC1REj+dC8b0/GBfEgyQ4G8GfuQRNbiMhk8zmGkfCh1cntXHnJlXYB61Nv
QBQahRYdKGUyg84GkBW/XaFCoOA1gKnvW9QIeZCDasu0Yj+9IyYp1yxdcpiG4yHS
ldH7haW60zVgw6KcYUyq6I+2o5eUBw0j7iwJRfRxPk0MPNZd6LHhOSrIjF9UzJpu
3GPNboEK5hYfgorNYaF2pbVUR7z5fqhMx5MWokzftKTMYhRrOoZNlkcljayLIva1
g5r4iGxhfLbRPrzSK2eldRS9HdNsoB7Uj6UoIseP8xajc0bVwbCZzZ/EFTu4xAE+
QkV460hpXYbPDI8hct8BT0hAkx4IXgGdf78HxR6tj3vsv4IeHMdsO1vo4gyBwXGX
vO+x0/y69elmoTon+MT1SVRSdh4PHSEU/HRDE9lW3KA9DbScdyi/tGy28IensIUO
fVlAUhySQQ0F3J7NNCp6+Gnc+NLguuPmpR/QhypWOqZSQwDcBfUUbarJamfnwwJm
mdwSOhZhJhccTFeqDctpYLvD0Lf1BAzqCVfO0GyixGa4fukGN7hrn6ZraNG8HJOT
CgxMHEioK4wLHyRNWCbJP3o6rn7YRTSQryffKfEqDe9y+S0K7JKwtB8EEY37sIuI
MvZ1fYXzkHahrakbLsFcnx0X6vmT6iRKMvt7t/yRyPQspveeiaEEW84P/eg6qDfi
pdl7SGylB9Iq3Mknjg6Ahc0Cox6iPLBxrj5ncf/QvWycgmm/YG0ORXooRZLy6c02
dHX3HD3tgpP5AoTj5gN2wXaz1AqEND1+hviEAsg84wM+M5incxPtiPPhAs6zBukI
/ZcumoxtR9Pj/ZiCjh1VRT42noHSmpIPo/Fdo6ZX9AbjsC3JMogQp3UdpZoLN0nD
/aOlBa1FFWStZqjrdx4vXIsPNyPZ+8L/VLFKAAZKmFTNCd+ybYxi/xoFemjo09dE
AScbm8fus7EkjB/a5AihMi8xaARRBCNzvVYWTRq8CuzXmYiiK/1IEbUApH506G9J
Q9Gz+cZeK6cTixyGaIM9U0sVih4/MeHP+XQod703L7v7LMlaBCp84ytsWu1WGkki
uoxiumamCqSyK6tWvmlspwoGLOQWjX4eui05MsB8Z1UShtmuAkxVPBPpp0Sua3By
qNwJcVCG0Iznq73pyVzQAaqrU3fttLOBVgoP8mpvwgguVaUGj/dobkIfABjtIa/g
axVM2Ung35oheANAN2vmkhm2fUgaB6R9/K9KXofgUK0X7/903Eq20i6/p6k1f4er
H3E3iVhN/ZBCjvW4083xXkLAeU43yTCuFSJFU+XM+TF/EgssQ0/mIKDgIBrffIlL
+ejC1qbc+rx7xlati9kRAc8DxUwWqgAjkWagT/ZivMAiQsYfDcCn609a4plDM0iB
LjrefOQIHI1PFjJ4YYkuxONzFY2f3Yh5GgYvDMzGDNnsY8cI/LTQw4PhWXH6CfUj
PUO/r5v66nqaL6OvOe9HdA4/9IEKQURq83EM+pqqQlSQ7nsYjcxPFEBlKMMsmdcL
OCZS+QfAsBaMUqCsvyzl1R8PguqTshgWc8DwAxwdbo2VewfEYK7dA1U6U1Z3dwxz
eKsIsLS9jC1ajkTpbfUxmnA6Olbg77kgDQU9/ctgr7eB/gvwD3F4mVi/skKmu29K
rDU53Ep3IIR7MUBUXLsGWBvmsE2TurIylV34Bm073xunASKjKizdonS2NR6VfTF0
X4t4JQuxg82NcCO2NrHChxXVE04nGM6DQk7MuWcGZLlr8+a0YC/e/H8SK7ksZaJ8
AHXy4iNDE3N4/7eSCl4MAsaKGTjKDjrORIvJ7LS0YGpXTam19CqS51mHI0B3ozjt
WtvRn5fzM5qG+tripq8S689qaciSKmyMeA3egNlXJRrqjrmpqogEIrCA5etRhFyY
QxjC37gXUa+R5t5fEtB6Kvy2bN6ihDer+kLZT7TC/hejzWbs/lMgafi/tvrYtN4+
R9sNtEi0OE/T1QhsGyzlVIguzLPpiK+dBkwTsUbCC/5ezXdCSZiBnBebf0cjxxT3
doC3BXiGEjstGqbzURdxaLMlIknYWymzOxPj3dftxpOqyLpxdopNglpN/c7Fpqy3
ZGSia1x4WJCfFRNdW32bBgN8k+TYz0F4ti+O/AMXKo2ny0luZSfYM7ASFYtwIAym
ohb2UmnEvSplxGKCXfuaV/c38qtSfq5ijYXj/5ifN5sgT0MF2qDvj2i0kUlVu9eJ
6jTmfCLVrhIfAFnR8pWTPlnXtQmMHgc2bXQzEnSA3sQKz7R4po1WO9QAf1zF9jti
b5bSYzjWR/RFvIuJK3zQAbuxjEsz0Krp5/iwkbpCMaw5PnshAkf33UlG/TuGjxmx
9DR6PE4FI7chFHadnPKwsvqvLi7iO3NmjIWjoVY7Ej60UT3AvENlD2GfUHNLyHX4
Qklgv/RtvJb7Nbah7dYyi6nn+PlcJ0Wfyw5OwdVNQ2u0irP4kwuli4eM44CcdEaO
mWc6SBhVY64DpJbg3gAp+BEi1bM2kz9v57hTZcWtj6/qSXTDSU/dfk8pHUQVbD9v
cZEjLWm+B9pQw3kgyKC/NFXzyVck5/DC5F+g2bELf6rQQ0NaFowqCK0YQ6H/IUzX
io8VF7TzStHydB1hFmQ8dYriLPi+vzhgcvjNugi89jo/wFLLxvfVbo+ty04z4YVY
OdWbun0nKomPxVI3mMS08KLJT4r3xDa/XMT8YukJ6/x3lG1L9XnAA8U51rV1Bj79
yLcRz90IzmfDiOAPHIf2sf0OK2PmjRly9OI31tToEMPgPWQZH7IgsjIxBMLuF1/m
3QqCPr8Km8772q7XZGczocLUhMEM6L52iX/K0TUN9Pigos8RMoFPJhSG4/EqVMoL
DH7Rr8k+21kOkg/HdGQ/oSHlJLdlty2mzelVQDBl3MIvG/cPBcYGcCpNmHFJnne9
Rt+fp4qlSCYo2ZNgSf93l4DBKpzE1qVd1kwX4eJwqsSZ8N6vZvvCWwA/uIkTL2MC
5yEB4p7Lf9wULDJqqGYPVU7kPVxEnNpGPhforC4kBdgYmCGS2RvS2dFi/dz7VNew
F8yIiajpfjJYipy6ckiyyxZZ9MYIHvt2xFmYpyNaPEKoyRxVst+IC4wkqlfQUvmj
mU0pwogrqyRvcTX3gXEryA9l8GNHU23NlBlSiypyCEbci6Bmafa12QQy+Zf8hoLo
kRYdELykxqIgnKLhSRe+eIpNHqTtjD4CR0lq5TVlaPGscb9eH+RKtPOvozr8q4Hb
C+RNw0K8FLo9CqIV4nzgDxSHJXqqJH7mZGdMxjoCEKWsWPUomPXTthJzOeWITi93
+wwlEqytSY9oOxWnkYHMwsGaHPvnU8L7xB1Efog/ANDkkzZ8S8vKYIEf1nDFdriW
jxpukNE9f8YVGGmcS/HAjvhB1jmmPHMR5xbcx5g2lhDP+s8AzjSzGp8gc3/4l79G
4NlixvhDLZQD8DDJDfsKFoALXAZ7ANj0vF/ooie3jcf9hBlAdTmd+S3AsdIF56au
NeROtVHZ/E6SDi/qp3cQ6ISK2DGpLVHoqt+dX7iXl/XkagOoWXbSjGGoaymryysx
7Xbx2AyNIKeHOkxTdY3bdqq8BBfTNBhAvaw0i90cN/JwBkgXdaZ3KE9Ou7urlRfz
ApNp53K6gbyUl++wFXwtrWZbhoaWnSqdcFlKevEXJcyBXM8Zdqgw5bdFqWlSvKsm
cKb7laUhDzPU4mn740CFSQmHOOuj7Pke3r+EQfXyIV7jDKKXhsrSL4PO6tk5eSuX
3IhsVMnAcnAaWnLUrTxnkWExhraT3eWrLiAXkuVEeIyOMvukDKefVwoTxehzAhKd
9Mcv4zYNmvD8cQSIMijj4FpAou4m/uTijzs8Sw2TYMrYvPfRI60EykWYykpgWna5
S31BBpJhoM6oxsQxtX02hf9n5Es8jlb8qljHS3J29zqC3mRzOptXWAFUMnzj+Gpl
oCKoqFpotQGcqANq6T275gbs12y+AdBbF2ltrDSUtBOi1UOH5c1JOfBd2jBlKXcx
UhoSyZaT2uBOT0Ao3Bj/StPyUfgcjCmfZLa+As51sxlS2h6XB9POjl5MtIT28Zb9
QPWFbIjwDAntYNpWnRf9KhPnJ63sirmgY2x2WQ3lKkCnObLMjfL/CkEzG/PeCFlr
DRKy21E3ZYYQWfj8BHDDrh1AHVH9g9ZOIm/mjXHYjkc5KV03AdyaJKFWqCE8FHO/
8W8TU9eNRgVAV/Gtzt7qzovUlsBOgffSbdTMq/dGQdNoAWHW69fXY7OyqPUmMysD
wNgAUgy5S6R1cnyW7O2fXwVsuUZscWwBkfbfFKz2mEm2yAYYcs19cMcppKrkWV4u
UUlGGkqXDtyYxGwDlgqZD6FkhosyXRkoQq6ApTsetRMiyw7GyURgq48fpro5Wh0l
REcs3WceJ7eNL/oVJpR1byJAmuFvhDwrogofPmeNoAqCipkKaIrpepa+w8ALEKuW
P5kR7KOgV4StbhqZwNaXJfgOantU0JYKGSYtH7kn6FPfwvGQwXXkapV85N53iNoR
Q3FelE45HPtsFRkxW6HfdCbjuIdGs8y+MDTleUlHRHUe2D7ptC5mtW/3O5FiKyvD
fFxbdc3T4jVaej6N9Nrvu8oHNcYg/ImM32Uze0DhbCR4jt652WedV9um0B35/DQg
p2hlItVfYSjAQUAL6TG249Ti1SrS4ARgkYaf2PqaKrappcWwvBoDLAf9/wGpoDN2
nzW65kEB03Sok5H2OkL9JUQ0ifowXr9eZZpmTZoU4kLsTR7Qbf8cJiGe73dVt41j
ikX+Y5GOwp5tSSoj1SPzRj+9Kkv4+Aq+m9SiT6mXtJXNqXWcMK6wfRRfsfgk9qyP
rlXE1nMKNEPmB+ryAyt3ZjtcUSSQSVRV/+90WwVDrvpGIAw29ILM4O50mpBOt2DP
urhkN32iM5GJ1Xz9pjDzEJUZoIYTZUUi9S8Fze9MM3QUY4CR0T5qW7DFLS8MJZ2W
DqOrPhKGQFhg4bTQNpP3EJiBdonSdkl8Odd34J5StzKNF6K8GLLueml/6h/9rU4J
ijZeKlHDsI9BVdW62Mi+1KD5APMvLfe6P/Zxei3/SogGMYY46FWtonM/Jjt9zrk8
oH7puT4E4HoXb/RQlD9XvrU8vJBrD5SearxrF44Vi56A6AF4PrQ9uMtgXo6n6I4s
aMTMM8iKN5hzwaxiPXM300xArAaFqprBidHiolMiwZUUB9SfmfQTxp/Wyrk+0Ib6
WKIpmf6OgYla7l4Oa/Yiai3cP7PAsrwf3nv1QVEJjDyiPqnpqYo7vrSg51MoPb0W
z5g8bYZshefO1Gmg24tNCqcNNg/4F74MaDotEm78LENzXuz3C8JIllsAZ9+jwaa5
HF98E4JkR1aMYHQt4yUC3Pmrx8ulDiitoiV/+lXy1H/+EDSQD0vdxlf97Y675CVB
8olonPUs5ZXUx8ftIh1+QUVng//y1v+u/FRLmdGYlBYPvCVpYbD3JLxNP7olUA+i
EdahpYgnx744GyArswAZhy9aPpw961uOCTqsoZjyplzZ8r476uHsqFemUIjZmKbY
MB5ZEPYNH3UCg6RtK0Y8/qxF0UknotR592sF3D173bPHVQqxdxMiW/kdyjsQgwbu
V51DCBFkEAhAZycC6DgKzYZcL8x/mdqfUC7pR+K5QgR9qQpHHMZTzQorLEDtFw0G
lQ1QlDmNZtyYaERfJizChQ4KgNPxFYYoXjypeRPRKvZ1cyyMZbBaSj6Nvqw6WlUX
togupY1pmfB0D6u+DiundPKtkHx1t8Nz9jqlVjpFqjdQq091sY7eDrx18AxCo05N
P+chwS5nMWcv1NkT8OMG2U/6WJ8rmlzXIp5rn4RO09PwVKat8K1HLNSoWvsGROcz
NC5rHxOjwEZJdJ5N1n3xNJKKSYs91jcpmGpeTDY5XPTyLFRrPW1n7rL1xZ3Ft3fS
5ApbsE0AFv2QRCDVPOnSG6oCTvVl4uyB14b+fyuVWxg4RYw0lKwbtH6OJOZj3ZpR
CJvbi90B1ZNHOMP1+lYAKFv9vFBIgTyVrG2jEIdZrz2r2XyZq6014i6ML43JtQJ3
DqmDNfzz8192IDM1kC5OdopVms+uE8zC+ufyfK/6AaR1gL5AClunbSTRAnFHYuPO
DxindTn6kLyn1mNsWYSFBDfo7NBXKHIqNkpLtBOKzY5ky9VlP4myJjmOW+YEn3Z4
+fcozxW7akdlNxaAACh6GyBiFFjPwmTmesAemdDQ66YT2TfUhDKn3NAMnrPdT/hU
4brPXh14xvcqffGhoVad687Uab2Y4uXZzcpurJXgC4vd45GT6+22H6jRYo5xMCCd
K7mHMmj3wp/n2/7bQRJGLb1cIq8ZJNLv2glIBwMRPhDD1YKTxTyHAln+avD8BhyH
eUVESyitmBlaux167JHS5qbzeTBZQzexVOR2FkxqN0iS+G5w0sbf4wg6xSTm3ShN
KxFxEoeVZ7DDix2TaQsYwM+3EEWsZAqqiFiB8fhJu5lmfJsuD6DRpiV88zuIoJPt
9u4+yCegHl5+AThXGXPH6VPkBl4dP54dSDp8gRJ4txAmqw5k0NPnuG39lTckWL5N
2R+970zrWXfV+5tnP+1HoHuyY5ubgPQ2lIddyRXUQOTpJZo/ZhaCT5R+w9QHRfpG
ToFaSJbKjsgLQq/TP46QKtRaaVZX+In8de1ve+ZmCzOMOaDVzpMNsIDJbz16bwzn
sClc/NJvP09U6gwjrT7pwWzxzuz7sKjxgrBaVYnh65FkCEdPP+K2VzP5o1UMExjp
llix2QPPRuCjbzcgnYGMsIU+qklFGp3lKN7Fgp++7F2gK4nYd4BP485uR8e3RMb8
7S4eNqLSRp+zVVCBKvJb0YjzUhdNY9q3nylHi/xMHNCS3VuK/0B2Zky9o53JkQi/
ImpIfJt8W9V8+Y+1OR7iwK+/xSrMQ75FtFXYwXz1upa+5r5pmwMX5W7jUA2ATkvS
e8epuq9N09LUe1dxUspbRGnET/MmsupAnHDh4dY874WT5fNK4BZf8udpyA8LQbaU
BtvU1YPgdNgzGjp+CMkU3F88vbavxOYcytu4YAepb4g/YKjTJuPzykT49cYTyKw5
TxwgfL4Cv9rhED/RVkkJLN3BCYuIpC/xusf02D7yr2iJcfrnJq67BMBqHDb5j4IA
c5UBEUZfdQbDtDpMO4+eul0V25EnEbyp1kZtDcfaEFPPBdIwR2NWcC3lCgo2jSJn
IpPiBqW+1/ezbwZWPJ1nMcaYt/KO4dYFh4n/6kU/bp7HDFB3Lp7hsMVe8m9EzHzy
wmMc3M8nubc01ztA25FeErvNz5wY2Kh7/HHET0guyaAu7XHagtF03vPY0xtoutaz
JRBXLunK8AH2q8/w16co06UnvC+YktUniBsGThq5e49k5WSBEmYiU0CAttvluRXT
1BI5ofIBCoEAe9rwOQahu6ACzQy+bVH45SGdfdFvprgQtgrOO8y/cYELeU/p0btX
064fLnVWdzi3X+q42EWphtHelxfJLAi7bBQbxbCgGxAUiNqVmaqX/KTjlR/ccFjQ
Yripn3g91Q/U6Axqyt5bqOpONuV6TCubuZ9yoWpFakCIR84zSzVJ8Bpwj+GdNHdG
DO1CkoAbxawCFC3aSZY6hHDjjvajM3XVjEtoOnc1YpliO4BQdciAGAZ5kCxKcnm/
S2jgWmWHk3vYe5Be1e/rGUkPtk41HONng4+8svK+lHkcIJdAdb6L2QPzNzBVK1Ub
Nub07aGqyBIBjIef8MVCHzDD7s7jbIA8frQLUNTlVrFhokP9drEIE5wZ7tn2tl94
jQch3ZFjj2G7GdrSuXEf55+ys86lTOHb43ACAAjhEcSQC3HGR1qEBiKZl9O+hOEO
k7D7SGRfQi6Ot0C/hxi+F81eQmSYFI3rbN7vrYMAdjbL61soGp4vtJd2Pwkb/IoE
WJ8T0Hghjq8HT5gcFs58w4mcKw+QL5ieTxelZpws02L0S/hgCmL+oMeKcXBYXj9u
bc87ZwC9JGOD+Vm94QUd6ltt4S0wSH47NRSwl0qEr7nLhH05xWURODQw3m28TsrZ
naIV0WkncWxRxs481+6CFSGZq/AkRLCLHjkHTMmRdkxL/cdW1bmTLLinkm6ClG7U
28m3LeG0tZFxYCQxh7UMm0DrPG9ETlDN3+WomL8EiX5HVmJ99RXP9t8YafZ1sGdG
vw9b03q/GAE61siIsbZP6c2tRXbGRzGhbTBGxLXvqabkLVuXrqptzld1UqXixkY4
e3oIkcENPDP9P3ZJ3OGs1uTJEBPxDbejJ6ROlEN8HB4HnwiJA6GE2xCKR4SFjRfL
jE0VnSZ1QB+o3e9j93x70oVe7oAra+73dB8XHXeYzWFK5PGA2zJBKmiu3Cu2+H7t
v+0X/9e/xZQg8T9Dn/HuQCejfmmWhsH21Phj26mx0sOEb7wIZRKJH8k1iyAtFvNL
4Sefx4ZfuIuplcmdqi+SZfQyL6+rLOLCGNRrIofscnOJoahKxY8txLYJ5VMqn/zv
FrYBxVhTedgtYDfGAwWECnDj17+puNbiB3Ee/9CzslUiQkVrGRLkT0Aa5J1XcauY
xBYBKPhJBPPmFR3EfhWECPenFdOTFpXHgdOTdK8uzTm9tmuiS02X8WOjebC1/b/P
yK7gmhF0B6G/UGHnVpQWEhUNAE1kpndPojcSs8TP1Rr/ZaB5K6pmOBATvWrZJc+J
Xyvijq1fUQeTadIhsMlLHV8QI+YbZGVHRWuNaFsNIguXr1fERhYG1JAeNLJe3Fz6
WngLLcU13hDfVJDkVrBNxOs1BT9+EPCzAakP1k9ulXUvlDUZXL7Exiekw6R7qqMg
gIgvkeiGtu7GWsBayv99D3fyIRiNO5P+jLnzQdMqq+9mBH93qgwp0qkRVTsVMU8q
gE/UEVf0RCSAK5g10YoFRbTricySfWdDgvlmJooyCRn366+mfDKcJJmvbyhgzhof
+iXmRVa+ZR77LnyHF2Nrg6TO3J6VpIcZyFM+sozF6ypQsVpQIeSeVJOVZeaDOVMW
Sa7W/cVDN26239f3gp1rsPtIRIj2ODUi2RDEEnJ9CTcStidETlz+RIWHnVWmY60u
cEqb/kaBSi1aWii5R4EuJfAROk+1L/L7Kxl+9vel3GKBU+XYizqBKyOjVkALYuCI
l/hygdjroqXgX3HMRWkNvj94ty1uzVyiPvMo7rlkCJF5Q7f2teVbvGMT2jDVB69L
cpX2gQFSxKf2MwMRR9FRMrUbBKsklNIyheinMQcKELUoDjjpmbeyrYHzt7yTPDYC
+KifC4atN3bBZzEvFIDBmtB389t+Ep7UD5jNbrvAAZ3ufKmRmUHaf/g4UD2ELdry
xH0a94lKAAp0/xi/DDyeNgW3KTxciOU6xs2EnEU1mB/y1PC19wROpXxqaEji2aWn
3H584RjvHQjOGuI0RzWXrJdgieSHXK6uHysZuPdCUdfMwkmVKk2mGoDaRNXpTZQl
viJ0WMUvLYPDBeItvAcQxbuDfd4vetZucl6Y2mQEjGeulxRSkFn7HqyeZ+ZRR4w+
OUGDKqukXEgre8DP53P7bQWYE6cLi7FufeySOigJyoLtX33JBsr3UHcz0l+LuB47
NPS5KnHquUOAkdGHN/NbQx9kmmHIf01AG9xoasgtM+AuIHY/55zZ9DIb1Dc0bmaC
QitJIWH9OVCa1CwDMhJ5fJ5iALHYRMGuTzdi5NzVce0BZStszUONTjxBRuUx3/W7
/kE+r3EFsBIk5BpoIdev4ZSc8B7ggtH9Lsx5Jkm8QCU4LUxmbt0MryrV/KrNDkpI
GE24odVW/Tup4lr/Ldj/z3PamfhfudCtNt748boBZLtD7a15YE42GwBVj0XBeK9I
Vc2w6u3biRRJ6Sc7uZJilNKmTtw/k85+CEB1CoRZhV6EV67/WrBYWLA5MsuBAJEu
O7mNoA+oup2DfcNowrEzpVX7/JnvQBiECuWiUgCrJ5I5+IT7Bz+FFgrbTM1vzMmQ
VE/UR+xNNKEUenHgJObhhQQplYCKfXJvrxJuEFEmsuBweYDdWHyGAqTkXsN6NxRh
g6JWSvHGxGoR+CgF+BgOkpI4jp/V0lvlQ9Fr5MHGrcEKoCjRjhOR5M5fvKnFqodK
NK72EVXMUM2Gp1CbceeaIzoLrI4s477QmuGSU8eMmC6N4m/AQzqjKMjwoZRU+nv1
xOoXFlcUDfYZCbAVw2b+4LTAljQedk/ae0JBbQMjYMqSSMoZN0NQ1IS6SzvXIwwa
d0mQVo36SOEwTbH4HKcWoKlaeKe8XNQg+EPPF6Eun4EEJ2ZQ8lIQ5wEilzAKeZ4V
A0KjBPq2/HMXD5sXUo8AVutWn+xtNd+HvFUGOu4z7zZkN3h+bh3s1RzAzNk2MNPm
yddXRS3sOqrxVErK7vxZ0aRWckQHBtJWaKgNpHOreDN2AG4XHN0FYNfhEv5nnq0q
ynLxz4Klu99r8eX3ehOLXhR5pjtIw0xDmLCbZlBzc4PWMsXe0eK5W/Ssu2cKbzkm
y/5d5N7hupIcNejVjGhQAbteAH5CUnjLKt0wK1DWdN8nE65MRSBINmmfyysCH1zr
bXBPdfxuLlRs2VPQkDnnSX1aD0DUC6YoYaCZtt13rSlVZnMvJMzRGdgQLsi4xQ4+
Er+05YrS/0kjY2hbYuScTcXIIhe2GYWGUSXOFyP1mFpSaWzSCGL9Ic7Bg+mvQAec
Jx2X5awFM8sd185sQ53aMDg4WwIGtFKDQQx7xhVnLImnQVdKdf/EzmBy2BorFhVo
L3dI6MJrUmafoFOEjs8dpFELSZjyPojBxQCbXg7LrYPn8U0HiAtNZRn8XTCQIbj3
NX9Z3WjoAk6qtgA4GSUYuK0+s+KHkH9IYzyBHLp2fkQEkm5OkZYbl8S3ZFMoUaMB
Epyh/uOwQFkROXOiS6HlTlzKNWWUOtIIkMbyLQAL0gXYtOzB3vrJwFSnLCoLDZ85
bM5DwnLJeRLhVTumONcqUeEhqrQrdzhcgVcnvY6SIBF64qt7T91/Q0ZWiM749IW6
VNi9cOsbqy8XPIBR2ENxMJGLtSplFgeQAaE5ItMwvYdCGlNkPPOTyydnGdE5Cpv+
ycqqpo6itL5+GWKpeG0zODcwCNQR9cTGaGordf+AUD+b25XZKxGxh4CyM5XxJxng
yFgfxYxcesOoJOSmVZ4Mf0IgYctriRR6P2hlEBRFr3vS13S+fumqMu74fjlrPnic
v22UzYiHSXzq3E3zeIUW9hI73diwP1904MG9+ZFv4/UhaVAjxc6vvXnDfJTAjepg
/jMPJ8yXty9rSdpIj8k/2P5QY8BU35788dxTIU6+IihNvoiJJq0rxGqK/O9QPxhK
DTgYUiNDD71k+uYNTB/KmHrTedGJutfj1zgc/XsUDf9lYM8tGj+cdVcfxjg2u3iG
cmF48qHNC51Q3quImeppvZjQB55yXKJoFnkQIoyh4h5wDKXoMKcGf3cxV9WvBrFl
Jm9cVtmyF+8XzJo3/XQL78TAloXedpdCIeJlBe0MMcWAOXptThO1Cxhrj6H7A1yY
WKxsUOsspPjIvpAbvvi3t6DqFSIqC5UkGtE2GUUi2Ol3FP6ipspdR9DfMXMaBVlT
iuVqsbuisEDAyQzDvXFKuY9w53ZYSqzpJCVvgzZ6M1RB/XQpIILW0O8LEpIcYyhx
aL2u1b2FOdfFbfTpKsm6dvjUeyC9fc5kidsuxMdheFyOhT+uLNY+pZPqjDyEs+Dh
/+h9kbyNe2suyQbibjYI98elrMtMui0WlzfLOHms47LqXGfDXdWr/lLT/MO1DBVE
4/X3FUxBfsWXY+gHO3dwoFID8FHke5+YT9vsU5os8bnu+kIFdX/qUHHXhT32Zknv
NaF6uCPAf/C9f1QEtqltqLNa7fsVjBLqxf1rQpdIViOFw7I1k/YRSDA0LNrDjcoM
RrhXjQSEKyiCi9rpLHUAR7AK3xmB2gRMCSFaY7X+1b3wruFC0A9RJX7RJFEtF22M
iRRt3jBIvgRnFuxgnrzP0ahlrT3Q0tvkR5ToEyMif3yc4laWrHgzOpQNflV3BYnH
s6fY7YnaOFLdIeJb4hLlq2bqrKIaFIyoXqWoXigPkO+rDrGkwLLLJcoCu81NMVYx
DjgNZoMLxMFqEIF5DnZeywZmGasCmKBs3Y0aqaPgL7iztK3Jn5AzQh6PwPpJ9k5L
d8Ew1jDfpyJJyIMobkO8QBZQu9VJy7rLzfgNmyx71rI/K2CrvbCjq8qjy+YWd6vL
jOuFmM/n+NFZ3ARQARk0lbUwtKWehGmCslvqXcbFTtLZd/qx4oleb+67Fj2RG7Pa
YDRXXT0ZVRjVWiAo/ZGbqK6Wj4UwLln0ZnQXnnJVxT3s7VA5tNZrNXZnOvf8wohz
UeO44mElcQyvHoSQG2y1T3/3GmTsA6fYcSvrTg8CPPui5JFUVz3emMA0VcDIqQ6A
5aY/92GC04OHAv474sFzvIGnjulUJtzUqeIJL81S6BNEticEhNbIW/TXo/tVIGuw
zfFPLyqxafhLnM25q1w3f33fekwsMhSujvc3POxijBG8bvvRQVtLwSStjiZIEH9d
XxgLjaa5PfTe91qjTiBnXQN6Oe6nJjVYJXxg8zxqAyD3JVHoAI2O34wqiTDgnwjr
WLe5nt709XhAXJA3XSxS1ue40LJMS0vS1e08sT8iT6D0pD/JMbk3lYVNPXRJaGIf
pgNqp3PluhJn2iM8s5Za2il8NapYrKvagVz8CjwygTVrY6iQSYZX52EioBisnahW
6aXR9IHEPIi4inUPizUTH8JF9hWnBuFTNsBF/za9vU7+5h5gXx1b2Rie8CNZ9g31
B+75yAcUAImrIh1lyStQZazhY3PoYh2m4Eaq3J20LMTTztn8QFVZpCEsUdXoaV31
I7a46GeEkm0LyW2BaEAsDPQcMkXjzmS/AvSoWqXWywY9DeNsusLPFFdMI0l4iEKt
mT+U1RWfM4s7TiqbQT9vtdpiFQSx+/GtlTEFvNY+4Gx/L4CriP2OLwcwnsM+aiBU
AdKusvxDTMbqKd0PW+qOQe/BL+u0CqlZc1u7xuXQXECKjffIiBsHZyfENRzsCQO8
HSae7S93KsXOVBJlShJ59AAhM1FdDfaQWJnhV5FO6/W76StTvOWCDy/SrYOFNadg
ml9087k/Z1keJPvPpB9Fl43w2ZW9h3GV+8eSvOGCwB2Y9E9ePnZbdiryQgw3Tm+/
+RTpFtEtAooRUjlh8NXcQBJVCupA21e24kX4ug7DqUvisoMj0T0lT3WGT5XK9H8+
9HaYbl1T0x/L+9rXWJ71Eko7ED69cn2xOGLaXiQean+kssL2i3layjJkUTl67ZBM
tjsqaaFPwUqQA15nfRZ1kGDu25gXnccboCoBn3kIg7bq30CFFOgfeZ/19thZMllj
Es6Qon5c/gWzAn7tZbu6x+FceLr1O7KwHydDLEjj+SDJgEPGT+aNgLxxPWCn9llg
YuJ5nOJAp4dqZ9kAM2cZcM4uVQBb4+M16f41MI/PO6a6cLJoezRSFRX6FNMJnAvc
FwasdsQ3vhTHvB44szzfcYBNMDJb84czlizQ/59X5KL85L6Ryrt5mk5Fcyxe9Vo4
EcqVrWA3Uqf9oDhpgoPcN7gsQpFMYZe70QhxQVQo7MAaeTSGfMg0gcPixL6Neipv
7/zz86PKN8LcOPAyP6zVYGySmGU01MQOyfQIaB5wDwmxoN/minqcVxrrM21CRI7u
Z6eZDveV1HWpaL/gYf7FH2FRvXjo7IXMrtWFxY89FZEFkGyHQvIEqIPl8j3QoHDf
/+lk8n6KInqB6N6eXnoaEceLORCVTt2s9SanOXvi6xktJrZHaQ7tgz299PjHNGmi
tYMD3yFKEZhke9JB7Ehh3JLKn+1M0fY8L8q2nREtRuEjnxSceiy1KSp1kRWSQFDp
LgqQ5Nnrky0kCcM7/432S4s5iemRG1wfUx+otbSP769l++mvXiPhMDc7OXYaK0Ns
oqrnSWl4uwE//BwZHI+XecBZ/ySkL6YgaY+Q4/U6JWmF+Q2Eivx+LkLqJvDbO/0D
e5OcLNbWI4QpYY1yN8t7DdqVstshTa5aadJswliK+U+m9wi+31Y2WEj0yeXTENLa
KSedN480V2HthT0kY0WHkvkPdTxp3hpXyn+y2awOhxMNaElQ7rc17HU3DVn++rXt
gT30K/f/0KdDLEYFKloqh3Fdq1zGc8PZUZbEURRAw4sJeYdvbt5oqmeq95lQEa6z
scrUFMo6QZGQLmwx2C3+/hlz68B/AXpAdDLtWyV3BYOUsJJqW9SqmyjgA00Sz71e
XiCUh4Q9sHyWRUQRRQMZBNkHHNKSfYsmIRsQ7D1HaGIOeKlqUNVyM+LdGp8fnBu0
Q+ZjpVym4INDicR3JDAjhc0LhbgNTpSlKh1Njd5aAt7C3a1rY4JFNg1+bfxGgMIc
wcjQurnP55YNNDwqQS47LpfT95wgQNG17MiGe6lOwyg4rTDYyYlDy5u3WF2HCPYI
ot2CUwadLIcAZThuwKykfZBlyS7upQCvzvJay0KwulmQjQcACOB+/9WKS8vC6USW
+okgMAjJF7lsoshkpJhma3HTi6wEolkoETLpgZpE9i3FSosGNF2xV9zK64mfo9uA
jX+61fdz7nQdfpnhj25uOu/qq2wGF+GiXGa2jeenTgvOuAPauqSBP85PnoaCk+ph
U+pBBoQsly2quzO1GDBeVSmpW1AW0IhHg8aMFGXmBAdRQrpgaFYH7xHVEE9oKQgM
3sOxF1ZDLvx52I9HwKOJnlR3kQjBmBSBwBiCse9/tOdfGDt/vslDadAEOF7FHGbA
d6jCYm+cWNXwk28kTxvpDKj62/p4eMKnSPfxvv5CAwJVlqhRtZTwLXrdXeeNvfME
CUT6PxetzJmIi+g4/6ilDdeIJMqKSfIi5U19IKUOn9rSmfeVwBgpV1drOHFueHfG
kIrEM5o76CtBzyOpFEWL+LcNbj1hojCCzB8S0ucjDZ1xLrl2+VBmYZ8X8UDsg+ax
PNPNhwC/3JD27l1MPsctllzNhDudypa83jlo3+gENoqkC39cIIynEyKB/yPRHefr
8z+O8UiPxN6oB6Zai9EgwOwz2s/KwCcdWHAMsmy8smQBDav8zbu43118mXBGTwbr
FIgjLaWgW4tp9095V+rH4JDKQaJjlu1vwVJ7Ob9xwl0fUmtSfBH9yw5Be6ESqjLD
xf7aOt7DulWHO4Ye0zbzF8OZPPx1eE+s0uo+1NoYuh+YYasxypl5QvhmKt1uwCNn
5LbEVcHMkj5y3NLCdGedBayYxoLyPuolKs5e8GMPGry6cFZO3JQvlljF3K8fMbpj
o6t8/DwD9OXrMvHvciDr4qFTjgp+vKz5fV4HC0O3YsVi/tq/immsEFY1I8mPrl+Q
3vtF3LhdOSqnWKopNZA+DxjCgp8Jp90mmYUdwQfSKZQgIDfwLrjdmtGSh3zFWPRF
Ag2y5MVMqnJ+BhTPgy4yVpVTA2yNM3ZaToDVmwnp2qJxHsrF6ORh6yVMQkj5yIan
OGRxctDAp/EHU2h/wZ17zwYvAvSceTXBazn4GMoWwuINx92+CCFHKNhtMqEdUY5+
Hh9YdsA/kZnR7FGr6j6d1O9Kbna98loTg2/CFPg0/sBQIl4+c+mxAECOgZr/CEZX
htDRjm1pOOhd386Gvy/f57nf6sSCQdgOQh/DcDbbn5uvigadu6/ZVSqv+QfgWD5/
8Tnk11ukJ9j2kLeuPqgBxoF55Afk7wzPk5Di+gDfUV+KJZeJ6kodsqHqitd0v466
YAZ3amOUd8zU29qKYp6vyjxwEb09kJeh376ame3fFERxk0LHtyoL4doToTcUb1Dy
d1/zHGDQ+AK0DRRZI5OjsP3ZYkPrrNuS3U0Wq2iFlWcpJ0qcr/vag3s0322BlSEc
/m8QR/SUEAVtHmNJtfUqMEcaIebGZINd3TwU78/hymv4xKoKThsEjsKEKPhUBbRF
UJtI27sPpIl3P45O5fhDvoNNcHK7lPZkcOHAy4CfUcXxDFsg1sb9tyEiTMe6IyfA
/7QNCciV7FVZNPI8pH6weGa9oUOztc2/djeHKaZ1TW+2JvhcMAt53GwxLNIIX6R2
yoPlfssuRMR7p4tu1CWRYZr3kbpQnhfhePbcMmHJIPnHF74ql4EtgEa/htvMKuNo
FSmrZnrx30x6cpdFpib0bfZeNTo+GOfyrP6Io/71iWNe3bWWelLEpB2r+BCm6dvh
gl+j17c1VhBIiWqbkX48kzdainqMhRU87KaBenV5TwqZ62IoCcu1ab5MAGG46XKU
v/Rq6hXU+YHn5sVN4EpUpEmMSUYV84ZIa10ckaST2fOANREkBr6WjBN+VFskpEQi
QrsDzNPYPDK7G0XOfLvM0stWr2Rm0xuRipFmORSgm73ZRfgsuOxa5sv03nn+tAb1
L83KwpCBhus9eFuVMsyro9VN8QtObq9kBbE3T+MCEcd/I7JCqYoRAszVlMlnCcoO
rFK1sqyrGrR2c7flsewbly0ldIfte1JQkSxaJnI4Qnfg5p+52kb12WKSZv3uRaMR
u7sUFYsAjYCyTVMgO00f1QwmQGmft67O3ExuvjKp8Qs0BsomvHgKF+HlItpGdrAs
jkMHTmovbmnFrFbgdRPmy1XPYdVOEWOMSr2Y2vS1qf6CgeSPeJn3AM1b9JKM9OkA
RIBjywSMv9Ha7NTotOUWryWrhTrAP/SZ4OqIUisr7bYg85Nn0Acnh6SnqbaJne2n
QVPeWEDn4QhviN9iWlzZeYvu9/lIgs0HjYgVW7xk+8/MUGVpZqiVpd/E6luDV2PB
Z+tQVDN2doNkn0zoN+bPw3XfMIghKR+P66dmqIRS3skJbk41ez0MRh+v/jrsAL2N
ypFwrIp6Qn3Nk8D0NwMUiXnUKnFNaoI+vjxJkjndWW8u3up4PdpoQmYwoUaxLGQK
rRlyU09Qy3+QfzJVs4rd1Z0LkU4jzWsIdWBRLwlIZWMmfgOgvhNB2OefKqv4CNNi
nbCo8eGbSjPwdKP+f72vCLyQVZqDvXx7dnumdI3CJknW5aUfv6a2rqOybNM+bHop
BZLQUnwpkAttX5XznUiTVDYk+Lq966IhVZDWAU27ALF8bU5DdS4pVTAUkOR07SEN
Hoda9P6wXeD82hM3CJgYvBjBX9zRWUSV2yHulZJgfAxr/zUK/rtrd0/WV2U4/ZnG
f+9fRmzm0/Ysarhe9k+kVpqz4q7AyhRVtywiGEK579MGGUhF1i8x1yrhZVhsvhF/
jyzqxSzcAjSpsJCS+Al9bd+hFz7g8OPhf0oDO4+bOwK7w4dvVr7865OH0Ov3GZ0x
f+a7pLckhNg6b3700NUhCkfNHqnyz1ynfZzRKhz+jP7Pv/2dTHxfCMnHQnKfKtx0
hITS4i5xvX+8v2PqDGJk2hYqjClGs+JlHbxYCkqJGg3rDoTNmZ41peRevfVPsoiI
UJ5Iqq1qfYee809RykpkpeJfP6F7fDAuiA5C09p+ICHmdO/yYZ/S5wUKbDn8pPY3
sNNKStSTGBhsQtiJNUTD7013gAlyrQdoxGR4nf35YdcmrHar7Fi3QFkK7LEUpy2y
XBPQGFCeDEsUsNEU1fuciFj3R4t3dcbRI8jiuVEdFVeVWfGImadpZclO21bUtZ5L
VGH96JzTC2X2J/S7wL5zNnBll0lzGvI2NSRDufQxX7mLgQI4RUNgpSA4boleD3pI
lYRFqGIiodDASxTxBsl3I5Sx+3KDTPxJfuFJt923/lvcfurJ7axIU95vILs3ikFf
B6Gl9gETGQn5rGj631k+Kti+Nz6QGesnt9EKA3tWb0GBDnO8Uz8AUzv9J09GshQx
wvc6oyqq5jGtNx+ZYDX5BmaXwnM6vkw7MAbW5SqAbNiC4li7pnsSyLPcOFQ25Xvn
6j2tD1IfidD+LqnkLSmfC7rFRG0Uk2SClq0AZMEjnngTS0qjvUoX2Hu+WPfLK9jD
6i6soGbmgJCIV5EcmN3wre03lvKyKPeLCf9zZq31MhN2xC9esj4pM9uO4lNCfOPB
2rdVwMBWJo/Dy9XrrwKq6nTxjTWsx50YyLmlnBDbpF2xa4k0WBwUg6YeCMGMTDsi
CYlYpugSSU4oOdsgbTxYw5ogmgfeobftvNH9JFKy7w/dFMFUTF3VVNnehpBXkHGI
0TXzgBU39MsKH4O7wcdyiX3/48vT5jmyB76vKJDCYS+ywt5L/8q4P5LRzwHixVUr
EBUNlhcRIkvcGpi/wYnxqM05EanqOIYz76oxsIxjycR0l8nlvbsDZjcCynB5cWlu
zTMwPS0eyqlDgGdA4gqfXo40LMIyvsqY0XIAhVg6TGdlAoJnmxKU8WaK6NFi6neI
4+kG8n3tvoEv7Gy2RJvnjZcPqbqQOLYUj5/4yLj9iTl9BDheu1g1HMw2/aG2zUio
hRM58t3Lq9fR+WyhCy2jBoYTmBvvZMQtGvGXWqL+I81P/x3v6mx1DUyCAcqc64D3
r+iQ/zMsU/2WTmlrKwKVRvKwaSVrqIE8Ojy2C8JOhOpD5q6/GAzut3oVNOEtNUb2
L9o5mfcQEXaYQdH1k470WQcqF2pZ33YUKBOsH/92dLufyTducDs5QDNVoU1IMdpw
9tjhh56BzezuYFDN2EiSiPg+lSoy1+ryAzjuCh5Nx3Lr2oVwEzRfQgj6MC+GOM28
D3GLW1w3iIQc/vm42Gjw+vispDxgDcrg82BHiKHxqNDx6NHR1QKCmXiZpAEYxiBX
6FIyPE4UB71EtogzGXumS3y++OY/myjzs8ibm9RazUEOzB/U1v5SlAW4YuVl7D6E
x8mWHLzSAXz1RAZtlT3BOAKqdowAEL/J24E4gWgZQOMYkSjnQGnMdmE4dohGqm+b
+3w4AIfRdGR3BYbMxh2+2wMIKA/0or+pZdorpighwJY7eU9MiQbr3hGK4k1t+S3a
k0jFnXO9VF5JH5Cp3gO1FeIPE9ZxDKx1e3TvMVuTsAFeJOZ+qHR+OiXW9J5eSgpe
qAiiJ1a5KLgygmQ/pYu99PuYp6vBpOgkBebrLpqoOuEM+qResHuVgks4r+vvn5M7
3IsB3IbdmIVKSAdvR+cF+pUwtROKrgid/Pc5n1+n6cRkpWHB649+SCXB+Pwm9RRU
ycwPJef51TvppdGoYx2lCI2wxw6R7YZPkwbv9ZKm/POroph+xB54Bh+KuQ3NAR6W
8kik8zPTLnDBxT7C/t1B+0UjRmycEeAwmgKeE7Dxwrcgc+mU6393vYFbKabg5fnw
guLLGImM1h2hy9WlXfB6doVw0QYFI4C+BsdC6koYlNaRkR64aSdtyjDILMfkihj8
pPPCTbmc3Qy2RX91VzYibBrU3jz95nNTHxr+Kg5EU/i+CQwlczJ6YLNODJjt6uBE
zRj4Pre35Tflfpeua28M4wFPSSjrYofbVb3p+sPduessaaP39pDtwd+0n+3zsONO
asx6v/4xwb8Bi350jd7zGebt2hdA8lBEI45ntYPYAMtCqVWo8edfNYJ56QIROtiR
B9sH13CUYsDUmbAd0iQfDozxJMNC+CmArmtTnOGFaW3oGBW2/WbH11PaJP+UqTmn
2yj146wr3LqjP642DaodiDJraej0wretoGN7ii0E+olgRQM2aqZRiUCmTVXiEuu1
OGnrA8wAelxPK6Uht0CSv/iifD2WWLxaHVdzV68fBMq2aZimdlG8BEOUKgig7abN
5BcWbPgjp7wNBV3Lze+ECpEBPlGzvdB4GF+JaHO49dMXP5+3OMTaeFmvYyAo5L7u
R70L38MntJcgBgKkaCidUXfYOrBB81/YPfg0GDfRHBqO7WWL6BUqlnKnxKve4Q8m
zTR41V7ZSjcLo28kfbxolwZl7PLs3l1uytjbbvwKUKpUvOp5HXel75Dr8uqyHv0b
RPGiDu0KdXr6u1KUvfuJW+IgvFTKKYYv1ARTE8tLIBDbQ+gCFV2mCobkGA2W/y/T
SAx/SfNgCde9CedjEK8ITPyvm5ePJ1GlYsHOuzZId8+6J1Op4ky+QSpnaSawMlkF
Q2K8ud68yGYkz9jOOIoG2t9wxhbOatQRG212GhGe9z6UicaZuXPEdvbuWhUu536A
rPvsJAHY3VRimFRr7TL4U6LXUyC8khisDJyA6ik6yvAxnFFfdzUlUqABSvCsrn1A
ocD03durQTCavwUOd9AzSOXTgP84jIi+rLHUCd/J6v0Cagcl+5VpUmoh/c8jbXR+
9hdUFQnD2tf1qomh2Ab13bYxiQbmz5LCyskgD/DNRKhHmFV86ElfRrldm6owaEEy
nWId8ZQphF257LwO1+IbjHupKrk0f2RYGuge3QyaEXO8yMVgVBTj1A46F213XhFq
o5eljyk6SG8EfcAlQPpQN/3QCdbJEdJIm/m5BcQhIekX4zaxB2URM0dXljAwaa+c
1pA533Yv95+U6w5YFRvy8RJF7bdUUDpT6tEBQ6+DWLLrzNzrXi4t91/CneXMPEsf
ouEQL2v8u0Er8VmES8BtuqYZU6Rv2OMQCSm40NMj+e0+kMt8sb/71iHgpBaA6cFq
plueLPL1kSL0ueLXITKePmznjUC836Jd1+g5BpC5Pk8U9e7uI0ZrmcmWoslqWuMZ
O/zDmGjXzEwAOSXciFSXQ/fqBhINFGAmlpPqGmRkMIAQqDthG6ylLr6/0T4+0YCf
cKfTnbuwGxA7BysMO9trGGs2TTQ8iF1Q3nu/kF5yQBuOHTRNcPi+MHIwo1TryyS8
27tklgX4iOGsYEqhJMiLZ6D78IP7lMZG9TbSjMSO4JlvAR/TYUBDoVlaG2GwKEyM
pecmBf1KIrLuGfeYBa10Xx/fVFxBKSNpgsCatDhjREZDbus5Y2EZLZ3AoHyDiF2f
yq6fZhuHAwajOqIZPyihm6+sxs4iQuTBhaMm2UMhSq+IXCx3Lbkw8mUxhmtLZGlC
bfesftn9tWOFnM0cNZL4/Eb96wbCsb9R/VXkIbRW1B243HwZrilyBDvl7XqD3npx
BQirgvNPA497z6TiKciY8LPztInOakuWgFB4c4oJJ/0jc1MievEiuhMBHQRYIeKu
kzwoRXLSzc3RQTm42RhsYtLwI29rx+M4tq7daBLfK5BiJxVEZZRF+d4k/rT20u0d
RnF640+Yqt038XfE2UCOfr7fM6y+KwwY9K7Eb1LtF8+oDyEGNehsvijwaYgE6BTH
ILmPGRoll9468cgnxAZq782S6kwkGvAIs98nVkOCRtAoacNLyHFyGCKyXaNPacUe
2Adqmhxvk0zoYxgBcw3/Mp+4tEvaeIvVQAYUfTTzf3CA6nbLORz6Qb9Jw34iOxim
j9EakgvjlNEbfU0NvRESgOwJt9Qe7utkIuUD4VwEg2s=
`protect END_PROTECTED
