`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gch+tocmt6UBnYhxSPomx6eHQdaSCDJB5psRTB9zLDVCEklomtpUV1QxQv2UEIv
2OK2v+X12NkC8jPK/Rn13l9pOdX+KTA8hcfqrZm2BhiMG9ju0VZYMR3wueG2lyUL
l7qbfxp6CIlap3Lio5x9TyLl7siJNX4xtHWhrPvtuvIJ3/QyqeI/N3zGI0K74dTz
syFw8Bx1dwZ31fX30BZVN+QJTbeRiXqZ2Qckd8FN1KSW1ECxD3Mqm2XmuiHwBvDy
v3IN48MDVNFQ9mG+77YnuBLhD+V4ukGoNqzc/6/7lrIopYjIKpK4tfs5yBIIWfOE
1jN1pGbbYoI606bBQNFEcI/yJ0Mc0nUNuljCDz81f6wntHu1kDZDdQFHchIJ3paK
7hk9xdHoYZ4L0s7xkGHWSXnbQ1c586cSDwnceGNFgbrdWG9S68XqCjkgBenfSNym
ycHQOLV4ZrMTDqQDmPQQQOO+EWxl/nGK1n2RzLxLHfm5BGvOMTX+WLdXeOjlECU+
MO7tU8nK+XVTtRDlPDcEt87T2fk1Jg/unaeT1eE8PQC8SLtzl9Mxuly43nWf7e7t
N7kj3ozJeC8sBYguDTyDo8mpaDAFxeJYzfNHpSgUgs8vHT1RS1afGtLwsiNH9mD1
/1c1KCxMyoGCpZP0ocYws66xmOwkfHX/bpgiQv0S0PA+gYjBHYLVxCIjWLb4Coq3
rzVQrc2ME0R6fN33LksU37J4nAFlX2RAEHGpctUmYRMK/8E7YJMsngzTMXKLF6/J
VPQVQheXxkxkkv/GarCGCzsn9QcNRHq7QlJN0OTPMoY=
`protect END_PROTECTED
