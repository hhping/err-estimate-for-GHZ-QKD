`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgZQZMLnTKMYrREbn2KmxdI/fMETw7rkwkjY8sZtuh1rj1SooP4DEt2nMPunyCOC
VGmTkp3q9UC2e4gWjiS1jGImXZXaMqo7Uh+BV0MH/p0vuquJkcXC1NIuR9ji3tNI
I2ISW7iwSDgZ6CuwHs1ixbdBOWTkMaQrrqWX/Yb5QbTf+6QcAiOwXvJdIY3Rg9sM
duDEQOtPT0NKtNSzBaBzR42pc4rzowYKQ7sfuydosQvqKezDqCw8qh9vVf1OI583
mU2jtQtHfPvhgiVYLPtlc1HDqMO87PbkADbeO10je5vwlyrRaNHZJS0NC0AfqXn5
vNDOlYi7q25nCRmL59KkdXhAmJpNElwuSaIFiM92z8v8jnndIzTNxNxDGuMuGxw8
wLTTClq2h1aaNvUzpMMy1WzE8N+bMSdpxzvjCAZ2NEDgqGmPzoYWIOaX/cxAriDZ
/2u80kErQ0AOtFKaKvyoMS8uI8IbYExb808SssExSpaarcbhBY0b/pTT4XgmGM3E
CC0buD4gmmWUylhMTP9yca9FsaI5mmqHetzPkLlo85FckXiBSdBuvx0OXxeM3xef
8n+wp6KQNIVS8VYccSa5dD5pzij808l18PiIxKVDuCrec1EmAcQIOSaNm1qMoPe7
/l9EZOejur4vHASwDdSoDlx3qpUYpurE26MdGoC/EAxNt9KU19FFryTNOo+2PMJv
gvqI3Q5FCxseVsE3A5sf8/V79OVK2OGIy57olUweMa93joQkP1uryV6tEGu8NlEO
rBTligrjRf0NhAj2jVdSHd/oAFEdScLlcnnfK3uZ2MBPSDFKRU+7952L2OyN4ikk
1BWZgROLT95uhOwDBZuGy20bmoZBWdL/rv+JVImaoUlrxEjS/z6KkPZjdHT8B4Ek
MGNVnkQh+5XFcV/SW04ITXd8MVlKS091ZWeZ/mnZ3ItGVb4QNJkH12nurf7AGsOE
TeBb3CwoPtfti6J6MASEMkAfTJaLwAAliHGSDhbzlvCHsDGNwYMkBDnoDbylVw70
sa8xVto8Otc62OsP6KY1L56Skvtm44Nk+BvdlmoXRqWGKu1wZsYnDbvOK4RH0LI1
0XCGNmckUtYJT2/McQ++Aqnp7h+l15mHJMOup/Q8VYTTaQkQFNd6sDyw/G6wQr7o
grv9U8rV/EGnWjQz0f8OxJYoRkSKyTChfIy9EzHU6YfC9eaZ8Nhd+oYfLkh6yrhW
Dwm3LOF60VP1fwtbTqaoOg9sDlBRpLtfqxZ0m8ybV085cYTyD2M9bxm/eNhExZBg
aVP04KR1zgLXxtweVE5DPIpgfnFX2XFWT7xvuFN7AR3UAyeG0BmsTfiiLYypkd0c
`protect END_PROTECTED
