`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T7Ivk7xXvpLAfMm86b+5xvQxX0EEZWonQW+ZhMys3d8ItZIkkNhfR4qyY2zXOuKa
llD+QQ6sEZR9RSYeKYrLbzRr22aJ55wr38gDV0TynTTvGDPcBcMeDGkEAgkULbw6
hjajqwmJfbfPG/aBebim9SsfEuZIXgq075kkLdI33i/DQ4uMeThoWY0Y501yZpn3
MM6EH9nT7wfEFuKitJNO6taGT+7ttS0skVkMe+KxAwBOQdBVb9T+jQnetl/uDpkE
V/PyASfH16g2WutuSlillCyj61+G7yxp665VsvbwI0g6m6IWiWxQdeBMENi8bAk5
loeaTrqHVcp37Nihxy6M1qJ0Vl2Ezf3hILz6R6HUtYnGnbKOPqksFngH2vslxr54
yHCEmJ+7iadnFR3H3Ls5D89YNcF2CFcDe0eNCImcabmpqc4JuCqogPocdxOSJ/wl
pUi+J0Mr+2kvXBtdANXz46X4gfxkyqhRb1ixTs+UYojpb9D7tHyPo5h5ZKDP035e
GQeAua+ihN8jFWdZRcDQX354G0nYVEcIkG67HT4mqvZPTW7f541gzXgInPVyiBn9
rJfrXW6E2dtNOtPk7MBZvQ==
`protect END_PROTECTED
