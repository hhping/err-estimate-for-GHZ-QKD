`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYsdeLKhciupdARfDsDiUnOavR4pAiBNly8n//Tkwus6ai+SsHDf1JnV407TwG9w
elSy9b1Wti+z6s0UQk1020RmiCgmFbAhr9AhNOTOe48TR/lLBZ0+P0h93u8qRSuz
Kt4n2ZXuTV8RoAiw29k5gzo1YW9EHjDI2SbcIUL3YXQJWitMDOuohvqz+Kde1gL1
+2k/fBvIHzneOZfKr8vc7RYNovlQX6vhraBuww46WqXb+d+XsssMgP39BxeKHmTk
n0mYgbKiucSo/FbQQw9dpkLuHRAh7/fDbZWPNubdJGXOyFNVX0IqBc2HH4GO0m0G
fHMRprVxUN6Xw6uz53FfbVZo4hY9TZ2gVQFDTuuH9PLLDX38QD/hcXZ9AnvinKXQ
TDTGrvIgr8fgfYJ7ZZWFOQ5mRWJYT4q09KuuKd4y7zvryCt412QOVZHHdQSm8T7W
n5tSJbuZ28D/FwugMaI0tUCx5aMc3Vm8wi7tHzUkWT9cSHl1wVrp74PM3huSVWNo
oZdMjsLIaC4iis6N1xWcF9knrs7pQcNOK/WGlh8QNIs+x1LFfpkmIbMWTsipFY1K
73Pg9vSk8PDcu6AY2jxSSgNfHxttTxdeEp7yoagdgFwAf8GvE2JTI6clMrGOrViu
4fOgpUETSrzXD2vREvGlHXiAko0G7wh9Ux6l0kf8xg/EapF5wtgPxAK+NTxi/qyT
FJpGlFH8YV45yqT7g8D+q6whIsr3sS+KYxep6/hbBAxRii5+vjgkxjLQHNj97/h8
OrPeQ+TmNtwZudNrrD8QDrm+G2K/ru5yvoEeAsFtsFen/xTxXTzG3bgmlsE1ciS0
3R5uCtBTEm1ZBpAp8KxlVJeJCoBdk/xpbF9csmBtDsecRx6445IkEzSmYINmqqdR
kJ8NaZEyM/gnPCPtNPoyMIeC4V5sMGHbnf+6LVYt8GoTTHWi6z9FJtWOaQCUahjw
R53VD5CyFzVGUrtZh0+v4bddMJkoA7k1pXyk12nA4D+9j3qFZ9LWAd4ywJhikT7a
KBX79Jn5iYosEfiO36+JdSREkD/oGua96iNpE6k98pcpJKLPZtMZsGeR7yFwu+HN
NssTyyyTJrG5Jb6xtPy2FNDCu/hDCoR6y6Q4ZO8w5s4P+hye/oiBYIdVNFgzgc8G
lXVlr0HFC6H7qzt6elntCh0GPOQkSFy9rbFyOPTO+2hpP8Ti7pu4AhtS2uZ33c9X
jrzfGWll8kMK0HAQbnxg6knZfRcW8mINTjnIDWsN93eCDu8JvFNB2p37bvyre2AZ
DqnOqv2HEhdPiVWpUjlCR5nMpu9AJmp2TsOqIwNk02KNyNaO0/adG0WjrN17Dol/
zdDt6ph7k+o2/kQy1cr+MgWzfZLMpNF8MGVgzSBTs+vulrzymwYwPpvNGw0jr1PB
BRNQXaKfYUwtfi6sjLF8zXOMBGXHBGWCTQQJSSuWeIKHDnnLpZ9zGGX97vm0WzXr
khJ9YLwqUapAD8g7gxe8P1zz0i6VGNIHaiCX7QNopkyKdCyuxw/S6vhMVzIpsMhr
iHPibdYwr4kukcz4JFnUkHALBtSgWINgQ/7Cvbm9KGpDQJZDHzet+jBRfaHiXHtM
QaJJGvsozzPDl14CLz5EMu0SIEBRr3S1NQSc7pP5DALcUKs2DwFeZTsA3awCXFYG
YRIzgqBcHoTUPkCRXn/r8HGMdtfVBJmQmZv2i09iKV4=
`protect END_PROTECTED
