`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqZc+9BcZtuuxyQclslwJMIUGlzBi9YT1JfbkDVtgy0BSwq5L2S51ysfbLWU1uXE
WDRlEFCahCKOAqTxoWylSXnjwr3DY1IYcCx/DOjPc0eVUSRbo0AMjcrLTEIw3juL
MKLsaJnuH/gODsqqjFxLGTlblRV1TQaK40Sq/x+C752LgaTvtxA0ocJ8/tgxcOIl
mcY22mte5u7tfQKG0Ru3vWm+G0abfERfRw8ZR1k38Mdb18F9s0VyLiurobjeMMIk
mgTT/JXtuJvEtHmmBhDkSj5vtdD84QpgacVvHdJJHdcrtdsVwaF4x7wx4ouawM60
t1F7f+xoLSpsT8dS3CGUcXht58Eqac8xkruLKybZB2K2xsjZqPEvaYS4wRzY2t0B
jqKk/7JU+OQjUCsP3GJPt6kXXQsRyktICwhFjP7tPc8esWTJU/cMxkfO+nnuZQjf
djjxczAiw1v5WAt9d/6mbgRmvju01UCaGg1Jb+xDZGOJ3OGIBhiIUcemZoPVmc3y
T8mym9A4zej8MJ1KHTsXu5V4YVCY9PpMix/u7DGN0y5dd/jh3lhaKSWGEBI6hdxY
kR2YoxMUGUL5uXzw49na/84ieOLeXJF9q8qU/dvJ0zlhLZJEczdgsZ9zj2kEEBrP
ml1EKx3hpQlyFL93H3eKvxprHIW+7E4ZjIiu+qD1HI1AN7ijgEBh6Z3rCQQDeI3x
PQi7PfZywkgO5grdAfwUaMn+/6PiPMsQPKfevsv/AiQ0YQshjhfjUEfA4nnFNt8w
wgiCjBfkp8KOxP14J1EQkZ55ZXqTy3N4W6gGtQthaQQDUcnES/7YEk30bWAYO/tq
VfVOATD8hol+Mxia4ScQ4ytkHdD8nz5iJ0/8vDDOHo7GqGUv4+GYwhJYUafPvEFT
R+rbCSrLnp/lFZIJG2tz5D6iS+ovf1xj0BYrcnAGB1rPjmXbERI2O53fRUvSMNbm
pbATHg08wKof5JwcNckZsxTxrLZbqbzljHA+CXzpGtZjfHRRgVlUdQP9K9HV1SQ/
`protect END_PROTECTED
