`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qo6vMlNN/LeSRQHsPWyHwQsaRtuW/+/7SdE4fYWT/YqmbpnNcx8fzFED24cdjts1
O827pjb+gqF4Mbt7pCmpYKmdWF6kAGiz7bcOQ3/Nt8y/GfqrMEmDYbW8ORYuh44n
TCh3Py4l4miE9Gv62yIwOz7DpINLUAuw073hgkGfvsJJEBXJVyk2EN7duIlAB1kc
GtUzgXCJ3V7syM6umQELixONQ6/VwPsLdgF5e709UNVlO5KSScd9M5E/4zhMnEqs
ullEF8dAUoBgkDJysGBbFqRRKELxZvBw2lsj1EvKMqz/xfElrpZavFW4nmN3xY1K
ePgDoB2Ej0ETNsiFehJ0flVz5Gf/BB+WeVs+pQkriB+3vgSPQb0Puf/am98HNMr/
Q/hIMv8NNCTLGjIx3m7YdFAQ5eiRNQktWDJP/fKYjKRVwkrgCV3aLZnRG0qatoWZ
g5rbkjsNB7eoobutnDj/os2qHmbSOGmZuO5LBppBxfeAigvhpRmzc00Dx7aBi8GS
lDu7UapZUz9qWur7HLUzUqX7sC/kWN3URvrAQD4e91KY2ZpeDlokb8V0Yh78otZ+
KggsLBjM7CUYwmlI/I6zMi0uwiitRfXlLbezSlWMWt6+/rbTz0fKwjU26rYvi9CO
dYuzoDWTxiJH7gG2dUfqfUoC4VVTB+TX8q8NA4D1kLbXO2LlR/rMCLnHB34L2yaZ
jyvzZEkb+C42Alugl+MI1IvqpOi+mA0zmwL4NlFCXsagyyCXlOr6J26wpyWWz1lx
coZcOoRDU2c8mLGKsLzuayA8Wyz6fdd1t+QeFcYFzSA7DGC6nyfuYNSmfXRswAQg
m796m300uFz7AAZDX95SFRK/ZoMYQpoKv19U8WWSMslApoAXGQeOeBtDjHNJzg1J
cJ3gqKGmFmJ3LvvzCXCYjft4cratCAzLTB7ryZptVS5DTZfC5koic/SJv2tTjHRg
abzPRNFxNmAY9G/qprB885j/oCxC2hsPKVyq+V+wYbCKc9qY7Xyy0t1yVTt4PU8X
48WXt+nhG2V6X5NOBJaHxDGHmydMwkXC93b5d4B1T/JJAixgvAkG7FuLuzswgehI
tMTAWt4rIgtzSkUnxbLTfYDMKOCo7LcYGFU5B/GLbUhFCqyeu7hAolI8SGWft8xV
YpU6rexdQF+81H5rhaM1kw==
`protect END_PROTECTED
