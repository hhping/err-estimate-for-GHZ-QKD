`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSROgSiXbZ/bsUoEC4dmlcSrNW6Am5usVUV20TWrMWpq9TYJvXcxvNgyTMeiw2jR
/TBdaQTG2IrUiyHZcIg49WsOiAt0SvpI0gu5Q0JBygzbzd3acWtleX1kNAEg3OvT
0ZKdd+mtXR9EEIJEkLlVFM8/i1sYqBNHOjvnOqtsPlVOAlKdORSm77y9bPmo4W1I
p0aZQDhlz4eUCt3GLSQYrlONKjSEp7c55kPSrl1nguJwsiR0xw+PCVHeTrBdsPCr
I4A3eQco95qsCnDeA42pp0ipWmB9MLNeA3vvnmdv/Kz84NEJBfB0ETBjxWeYb1uV
3eaaEqDjFXp1IrheUbX0E0iucUeKwWE7Qh3xv9rKWDCc1VKyIJpMcI673PIKtSjW
aqyW5koIAgw/KEVEIMgjKIkcw/1zsLP72IxSTBRydSJOaqd4FIfQzlmklUxAz6P6
wv2/+IPKsb0an90xzhBMJz8XUO9b0idQdop6uDwbgssUAgDakrYsFoZptd3L9aTz
JRZxjJnaeapHIEQOKpvzDM/pbYxzAikugrOMRfTcpDmbFBin+Nm/D0OrE0DwtLur
IFgTXABA2JYZe29g9YxqVADk1bJkeFNPzB5IEp6H0YR/Ji5GmJZK5WGRaYemHQDY
lD7jSKuMtfy8I3pcUpyK8MhVj5i8v5x5KKt3UYCHw3bANZbr5QzHzIvr4wlSj5ak
RFfJGvLtrDqAUplRJ4aZ7r1grOPyOqsStSsMB8CnHnc=
`protect END_PROTECTED
