`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4wh84vhe2zr3Y5knOnA0FnPZ+s/4VDoApfgoFcscBa1Sj+Q1XddRDGxBLrDRigp
qO65Y+gUOXlHi9rNd7gl0fpAhtJbtoNWpRm9NlGJCPrI7bmBP9mew4hL0qBoVmt8
lxr3HcecuhR+USBXoYdrcaGZF2pOoSTOf6kIKcRKTNOfch45qM5Iy+1o8MScN1lG
KxltPrrNQ7aTctf8AyjvYzct6BQMtEOLYy6Tgl4cHMq0dchD6RJToc+S0/ghX/oY
aYw3GIgX0mDVl1V95T17nce/7aQ6gPe7OGtfWK5wav06wV9bSk2XCljB31vzScke
su5ZsFqLeU4WMoHtTR+tNAWQx4Om0m7UBT2HOCloaVq+lytG7jvYXked0ajoxEf1
SQRBCXQ00V09xxEN7mMr+GW3Y9pfCKKUJ4+3k2Q603+Z4asqtDzElenf0TPHJHss
fLu3C6Q+Xxt/B19UZ5GHLE/1Mk4VQwkr/rEQOV8IAx3ET3K4IAfgm49Ob8bvrxSC
`protect END_PROTECTED
