`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQwRNrvkxhPPxoZa0PFIqityeNJZixAxh5KGZklrVWEt3gmeeqI57uAgZJAgEgtI
0AfBmTAFO1UxGKECm/ekZvq/D24gLLFz03yuLEby/ulvItFGcdfTCWHWiknEbCRI
4+rv2Z8PwwWuG6ky0UsiY8bHV73awndUcTHdi4Tg4JFlDQDG77T/HZ90tQ0NWLA3
vYVl1Wu0PXRxiB8L1I4RCQFSzRx1WUeogX9r9vHYvhCcG0InH1cA+INJewUcuk/f
Hb9YRFn3aSAZn/AaRtzz5Z7KK2jbi2ebml4A4QC5MiZ5+X8hThUa8ujQio0jsIAg
tNj1tc9PmxTjtXaHg1k3Nmicxf4NLbydpXb87u7VRfZn+fKUPV6TE/CndY3x8hb1
ZzRYddoU38roNiDjrv/r3xy5WDoU9E3rdnU3jikqEdYJ6fUVRr+EZtryg9TfUwvB
JxoY4dwk6mSSo+aDiXYBcxyzgzK4a94i4tSIisy2hFuz+yiF/s/rXjBq2d3jb0S+
VvXJdEbwliVgHAzHLG9oS1OAjjo3I2zADEZfdPKddFVMqfzTuFIKwbhoM2D5y+GV
2+j7NyXxJbT8gyAEIaeta+8tqsflq52GgquWSuFCs77Iq9etzWbeENHgr22k2t4p
UirwgI02z6ZtzRIlFC0cmbB1J5ImJyWPZrigbB2LmmRFewPGo7V32saNynT2EQig
f1RalQ5VKrroPXEuDO3BAiuQvLNng9JLIrSxgLvhmcBk37CLqcL7WHgTliZpIoT/
US9te6emAzshy5e5kwDB7s89NH8Vfk0S5D5KMF2O6fB4bbXXj4KXBCmrco32Ohsy
4oRZeVLwn648v+NkreE1Ma8OAduWA7R8G9H29iQAX+zPhx/tiFsLU8oB0rV9Rw4p
cqHcGqSFxIsnmCMt0uLmMKgm8X336JY5QYnSilFPmvj7zGd5LORnG6nfQrceAmki
GnbqKAlT1S1RfssRMOUs84Xfs3lfl4++Ala4J0atAnADDxWCuTfVq9uHTDKC/xGK
pP9sI778qQroNyY59OmHCvNgKrYtuTindQXLgEYuWXvnhieOblC44oJiS8T0RFbG
t8slA4GoXZ3QNHfkP2R3vjofxuOj+Qq2oYyTxrVtYPYpFJPu1kzIpNErzqZ9gxcn
+Zk1usFZf+hDIE+JIymzZfzS2ZD15f2z/b9mbxprW5+DM3KE1YxkJ6ORsGWQJlqu
SwtZLRvYLGbP7Y3QBepKCqa9vSYV3Fz1tQZZ3I+REQ1CdfLHWcZEGmwTZmHfIOEf
5oFMNN9I8/5E7ClEIfYerl0OYdCZNgmI3TN4Qp7i6xgEKi466CSJdpfzKQ1SQYzH
zmjCuqf31aW9HaEupQANIGnKAvCyndvLHgB87gmQOnmPu/fE8+Qaf5jdyfmtFqKt
LhZjbqJcpbn3z2xxpXH9NLqkdi0aeIZde9ZBLmzajKrJ1eN8t8L8Fmrbw0gpLO/c
+lY/tVqG0O4cUYZkwtAwwrhcUeRbFhXSkUekaLJjGlhortexADdzAHX8/nS8glLE
WoSMhE6AGi7Fs3rXVM1Oh57txAKoPOGKMiXtRIDOKAvFXHztmHKezdhu3eoYDDUv
59OrNYVuz/uwW51o+HZ/xiZGfr2t9cwSJ0zrW6G0kUd/tp6UcWTUfNIXeREEvg5R
AOur9taTO2w9qL25KDIdZ0Yh+Pu8EKH6mNFlZqC07U7xePSqbytajauaA8XuWqEC
MYnRedx7uheso7jKESInrCjcKCZPflVIbGB9UfEP/+eXxW7VUvY33+O30AycgSX7
K5hL7NT90ZiI7oUHH1+Xsu8cqwjqQ++NG3D+iah3d6t1rzdjkvwgn3L13Z/86xs+
iuFshXFFm9A3lfKnZTrL8TuVPaQvOcG4cmbRWUUfjT5jv+KdYMZ83L5obzrC1Bw7
CFdF/LokQdlU1eHFpIaB4kROtxRMGBd6NU47Wz7F4GA4fj3OopdUfLnQd4QZ4yAD
0bhE0qNlRhmwp9BEqsm7vuyufItwYpHDEAIBbo5jSit3Hr0FIbqj70pWGBAMZ9yC
u5jA46bk/Zv2t2vTiywWeC3SKBjw/RZtoeuOVBZzyWjjkGmD76FdnE96qIvTh8ZM
KVbBTgoWM16ltdJDzS7E2jx5Bnw4hA9pI1n1xodu1wABc0ZJOEewUa6/wEC/3+PW
Tw8yqFRp5cLcL0eik92Bx7W3iGNjW2Wm9x2lcQO3vIlY2c/faeCIEFvLbfgbR46O
n7wEriHfevNcppxDNg4US/VNAJMLTISe3TRXrFrLBqE/Smwyrc1ebuiUtroCODrK
NTUkdjw8hJ0SUFArmTsG1pWdAUaePFiDZLASaT8QDIaftwryIiAIQwlGArCjol8d
LgwCBaPgUBndzbiKh+pqCSEOde+TPmn7iL7e2UPeY72K3knTyvsmcgMs03VWohX6
bY6Ju3RmpBv3KQpgch0p5+LGmuRR5qoxqEmnfrXYLbZh/sLZtXp7ZLg+tjuIb+vp
GmDqJXIzr6ub4bh+LYuJVnnkI2btGX1abdw8BVM2T7ZqZGEqLMjZV7cqjwK/+bhl
p2meADjsu9I4QpmRLceXKEiMa3A4AcZwO+mJn3WQKk5S/Ifkye3eDiagdHtd0KxH
p8FgifAnn+e73u2UH76VxheOUanVuQjNwxJvd+3XOacGxw2n02DZquJlwgUW28zO
v68HL1fy7kDfd2vMr9gdiFpfSLfutdrLzdN/7z07jtuzJBEVMtSxh9sA64VPNAMp
7sOTYsL1B7i0qnFDc1FTZ7/p4mImAH/AGKUksEAhEMiQOunrcyqpVcfS0KZMjNcs
Obh/2hjIxvrglgqiDRFGe2KEDLrmU/l+IkfZ1t4WgB1k5lNkWtUTgxauibYzNRWN
Mq0nKvDki6EZRpjXprujEp1QvGlIyQVyWAIBnZpxrnJ9fCg/zAP95rhNsfX9nmQA
KVNWAjNAax43gYGNSBlal9SHtVwzVrl8NKlwb81221iMb3KQ8tx7454So+Rd1/3Q
yLw5ezTHgAabsoBTbvKTkAuXJ98Q6gY1kSgxZFv7jmRl9FqB83P6rwEnuDm03eh9
oeMgeVu0TwHytwyh5Vq1o6FK8VvOHftugF5TPzUExFDsSV3IMeVRF5Le8F6BCZFn
Zsk8pwzboZGd2ntCDO3GmEuvf8BArGa7v08KlTBGByUBNq6ca5HWi9YUDCsKiE9D
sLszlqk7pQ367xJ3MwT9kWQ5U+NhXmWKxdy1nS+F8jwAeazBJR2TkKNVXPHH7CKR
loi5AI22aAQdrKEb/Z978FwhyMITPjs3i94YP6099RDgXPReZFBxOoX6E2ux0fyf
cCjPpMpOyd5SW7t+T8YneCruuzU+FFYp9xuO5kOvh2H9Y4mS8Jdy7eQUX3hZF5vR
jlYJlxGTUe7JAesfgDXHKri7BymPYv2NI4KMMrtyhP0ZZrFx2buu0Wc93M5I5RiP
njApfTQdxktIAvd4GFE9PwTNNMSqnjo8j3hS72axlANnsycHDO8a/i6s2BRiAKeA
L1OzsW7yXgNdccWm6hwex64Ty/B/m+TG9WxcDSKQY5OLvZ5dtks8CJ2sH8xVHd0l
0rBdinKl/TLMIijad1+oFCXE2LyW34uLTGh7ATbeXhitqw66oa82THzospKvWgtq
Oe6mBQ2bYxmwiOwbrUI7evsFhNRDAkJixMGoCy0smC3k5SYUAWAYX6+tyEth2Xe0
m8vfcPC/pvyQ6OqXWvgVskffYF/csG9OYo3zXoI2KO3zuJRF7/FSnhRPOCGL5Xxs
PCuDBSd5eXlMi3zwqMwdJibpld1RQK/YH81FY0Z7BSewiR4KFAeIO+RnNPoxGpHp
y6F2ASd0k7/mhKXxbILwKjfUBD+t47MH/eBDoROC6wIqm0q6LKLRExRMNvLI5i12
dYhV4HapBGVglmbKCGcHj1y/cXS7y/4bT8YS8AHH8BQEM3gh+YWhVlaYVcSbxq2x
3RH4Y1NCSQENkZRABuj9jMw3rwJ4wnA5FYmoWDNW4Rn6OBimoY9N+nh+x24jT1vb
JSU+wVpJ6zza7SqPK42D2hFjUT4gQ9tbFdryYhbDyQaErDqWllGpP312NPCcuF+Q
KNzeZ8TOfnnevGLENc7SHxpGB9P5rwloFC+7oJ3EQNj6BveqjuKnsEuzcCcZdzpB
bm3KCuvV7aKYG5zYNs3BMM8Xga5oucxIbCOsa9gnWrqe6lrcyW2U9mMSgU2+pXuZ
xVFOSL+eGd8pntkrEtlUEuJehczyWWVSa371FqPY8pfMiFm1PLLQaOch2kFkDmey
M7+/FGYcDbJXxZfbUNKzk+jnAaHmR+eyVesGPOJo/nFopUiEvSV/vwl182Vs1d39
iOvEnKiz+nZPoXAGutRC4cRkoKL/U2Qztl9QRx/N2ULz+Gy4G30WtBIbw41lGGH/
2c6cEUPHMu1e+yLecpEsrMoZO10vmocoQ/zQBFaYfWdm+leQiq/uEXO6ENC9p+w6
+DFWt7Jf4BNgP1Zju/GQEYy7EnPm/1tA04zRXJLAlj0nvwHQiMkqPsx5nTAFTciM
eli5jIIUZjvQSyBa39W73PrKqJwwpWGGYM8C5qph9pySkTnQy/XmNgUJit9nB5wa
0rwFSJ/4NTsBn1MfELH3wNsqzbAISjL8UNM9J0rmvxi0ieTKvK23X3IoN2uDe5tq
HC+eiRiL0obq5wot0sXsfBUMNdKSSDvb373aFPwA7bYTs1oJBC1W/PQ7K7v3XgF8
3pmmOVAEFlitT99zZIZ8gcqPpIxCl/NwpEMoKf0z/fZ0PIAqTU9engGp5h53+Bnp
mZPXrXKz3qaxVedMM59nJVwR3rDdMpSUYOeQCeqhGGMYmTWF5+CBxJWdbPqWHnaU
bnvMxyg42R2kHSHagyyC2gVF49KOzy8/Draw0eBx/49XEJKjakZwMDU6UzlHh9N3
HrLIR5UDvpy2+pN+CCPl6U73zLhGKmjZsgVXomOr2QKpl8ptNxcQJGdCdxOgNfUn
v8J7Q6zXzQnGrzyYOFam97AZPRZ6BeDYPPvGc4fkGUyUYtdtVQaa4jUxUyEKmAXf
baza0jWUGpCNC84wempKiwNxmMCTQ3diT1oGXzAsj0T4iTyz0NbgbPxUucoQSSzJ
KCgVwGmCaREvchO3qQJxGZy1IqXjFQYMnvUtrV1xpAAOHYTNVBrKH6sNrNAuczBS
5HwvluSOrulD1enoGrHYyJfqd0z0vKGFbphOVvprUQ6ZLUVxMLkanG1T+ZYC2+X7
nNTAez506DqtpTlP+jYXGT+nvl5ryz9al3Ytdt4mkIiEztFTyG7oTiwEHGD8Hixy
dhIeIr3l6FcASM+pOE3WLN2ai57YG7czAXjw8EYRoOpmzeccueVS2Gd4+/mbeTxR
jh7kNwuSJnf3Xwz60yvp0IwAmWB66JbrpuQbjBKIqC3VrQzpZMgnFJ4eV5IILP/Z
N5Q1P3Lpbp60PpgnYrkQuuzzjJ3ZkZW+sGm+3OpbigekTlPQbg8Dm9tL5zRQ/fex
Klcrr57tgdOoU5JMsPIsZy0JVKfEiISE9QRBVhAqa7Fx0hVEdkHsjroPUZtrW0im
Eeq2i9nMXxs1+V3wysH/thTdDZxjJgUFyfTAc1y10Bm9J9egZ1IxID7jQxcsyu/G
dRbIOosVfFLmIQJmbNLS44K398f/ejwA+FxyJEctOt1T3fwR+PtLLi2HDW8lCR2i
g7FgpNtSZU+8OuA5UbYskQ5JYUhEvGwdtP1fE9EbHTjdRX2SzIzE9ObfrRyL2N4B
DQCegCGITCLFX+9fUYmX9nzlYO//9zsgupe4GCB2GatsUK77R+M7WN6FySELur6E
GJjKfLP/kJfpRPQeKaCq33R0Cyg6GYxK2MQBnYS9sDJhEs6Ee9tvM2dKkV/3NMuI
lzC/uGEXFqWaH93GuufyNPQoEdpF3Y0JTaW25fNpjlBM8Xq9mRH+H3wz10gBwXmK
DdL2oE4/zLe6r07ovze2BkUyinQiZR3c731ILQnwYuXiIiJUvJYV+vYQq4IdSemU
khlqI2LYzZku2rZzO/jbnWqP0WTI17SZdcPxHyJXwZzims52CT1BdEL8aO1cfp6y
sD4+loKmjJWFi/vqI/OmRuP8wwQ8s5gq4HmqUg3y5JapdmaCawTx5S48SJGAitUn
q2/kEju1+g8PyJ8/bsuPsnDgJDDo8mfdhnzN1hLIdhRsY4EHjiGaLER6rpbV0bCy
csW9w+7UBzSiBDLkd20RMhpAVcb/8kA7EWlLLaF2Sa6Dl2Qd6N8f0K5hJ/WhlmhR
WWcDkOL9NPT26efA2vDuQ6ZrizpVqUWq/z6te/x05wtat2F+TUq8yODtEVwU6giP
rxgjj5fATZdddedBtmJeLKlDf2RLg8mxnek9BD/fGVnrI/D/eM3/Trr+wqkNYZJQ
wBPvp7eKyP8VYOneCyZypp0QSBBpqCz4xZPjsafZ+rxnNcPZFE1BWya3eMNtukAz
TzJIKUEFFNkaS9mimaUnsJla1KIaf1ncW+1KdN42B9kRrEBkvGcM0N7ydnqHo93+
rJEHBDhomDrh1Fwiay/UubdI4C/xeD4veqSRxVyT1pC8DwKRJHrQd3RcndkFmKz5
UJY7/SnRiX+fMXLghu+joGCIx+uflFRuXqtas2izKKSf+Dc2xpyh1xTY/esoW9Xc
7wT8A2QQCChZvS83IGBBzGiYm5JGA4sJO+CXsxwdoyvFCu3UHJVpi6HUa8248vqm
qyhAseCXSXL6tZoduxd5P2hgptPMWhBXIc9r7FEIz9N+lYfDojtjZ5iqGx4UhHM0
aLvLQwnCPlKMUOzE8+I4HyCN+VQSjbIK+PYvEbSuDzzcnEP1UalwSQAKT/0SJE+N
qvwl2LvFzIe8K2wAcVFaoRo0IABVo3EnSXAx3AcNNQuik9jtGkpE2pCjslQohASX
Qmd4xOKujBT6EKuAjPSF+eTEL6b04uG6su3UDCWDrmd2rF7LELTOr1GNONnCiMHp
2CsO8AN+OrfX01DQSNWr0VcABoWAWMxNFe0OifwGnBkanWZ729iXZy4fK2jgk5D6
ZzYKqrEn80PW9FKzqj9wALqeDLhXjLdFfuKVbrnTAv8tOXPheBFpjRIW5sghJihl
9PrQND7Pdca4eDRB8O0DyURP1IhlKlpk8pdpWssEtQvpeKp/czgPS1vtzRu9yesg
QDrf33fxO+yn+s2H3fTElwZjU3rWNMF8qDZ71NFacfQqODtUUxHlQkAMSLQeHgjX
Vk9iiVaAQbAoVh/oAgtEVm5QVt1FUmntdjArY5ABxf8YEbDq3ntNpcmzBEuwSNY3
0ICr5eVzz94SHhF6lN9hA8f0p/vI9b5nZQiir4eo+NwJISRu3LLJ/8FVSlMvbBr0
RTEDsKw5QbsbdLRJhpw65qU5KQwBz81LTwYEBnwmBRV6+BoRR13RDXgS27vRD4HV
xBmoBcV/fnUJy833zAC503mWhn+UIdmviMiJiJ7Te2xnhyx9Tq7OgvzsnBYutGPG
ha3moa9+F92LL1btsA2TrmnE9ot9hEx3tu2aHtfvaG5OO774fB8PO5QhaDbiMUGJ
XiP+VYvE3QBxx0fGBX6H30/Zy9QyQ+TdKTv2D949W4GCYkzrkl/nxE+UsuzBf5mG
sTho7XBjOUBpEEQuwE/xLZGIi/C28ioMN4i2Cs4WUru6joNLpSYmx4dcctHVlAJP
hWwld+zQwOf/T+FY5upngxHwPGkW11xhMfXkDbRv3jaX7mpiCeu/OfCLaryVyi6Z
JmgCYP97N2FVRjGVT6ZaYOAWhcj2LiEKFMDosQ+ioVEHyhjJIlauYNhQv66Rq8Tv
JntHbQ59Lvwu0qVRDWrOWq7BpcKZ963wxAOdoxpmSWB4HHs8R0EHtHHK4ZXxjxww
3zB63aUMw5zeTRWE/rMso9JL5VaML5CQQssF0Qiotl7yfLTW3b4KMY5VNC91cdVN
mye+4p8JhWA/O8Yj/hvIxHm6XbSTeLvAGai+tVb3QXYp2R8KBomJCyefmQz7Q68z
Q2gOYI1en8kIdrek2l2vqkrFL2DXXsRsHuUjt8cyF/GxAa71wcfXyMgXNJhH+6bl
kTXRebwWMVCAHq/00xfAhFm+1EowTybeqCftRjDztXBipWtDqrEYJLFaYs+KFiko
w+Rwuz191MEW4j9QzqRdLZBbbnY8eeNUdz3pJWpZJQ2729QD8HRVGFPyELHx1+q3
/RX056Ez7B37QAqrmNFyrRH0F6ycJP1FyP2SfNTc5k9kMfMjaTHHl3Le6hAxYG/I
VXJ1MJ7qKDuHqaNHTcrYpHd5VLASX7i8jbGP6SKRoMgYhMxLSVyfYxsa8IbZb4/8
lngJbrFiK4uCtsSOsfA7ULrbc9eFXOvwY7wACe41jtX9hEiUw77u9mAYyzJx7nob
Vbkoh+W9Hxty+aHVKup4TkbblsbZhwz3NrXFjIwb7YFs+L0qQG532uRbsogO3XUn
LlhawDHv9cQqOseIDzLrm980DmlK4ZeEWG8iKDiOVWuOJKM0dK1t+nEAunMenFa7
KXhO/1EYWlav7z7krpR/tcgWG/TUWNkwN55h7RxxwUulLRg79hjRGI5jDaeD9sxM
/3NL3HgINfeUreIp1inNFSDZlWfLMXcnjK+4Qfot70scYs5ApGMziaMinLZVeDjt
lBTchDT5PpI/XL+DusqLPm/KmX8jnmnXR3JfveSeI3GD9l/3hH9CN5y/kEzq7CkU
Zqu+Zor+gCkh5psWz3WTZWBctjNGUVSw7ze66SdPvakm+MpCEYRWoJZCadisLWYN
te3phcMdRDXAX47tUjjhahCtENr4DcVJJPYW0kGXhKDtpSfAlZRnSA6FZD8AK/Wa
34umBqAUbjZ1/h+WznuVWAebbaxtmEqmq5mBIZ8zaDVFfqAm22ITMxExCuipIakX
GLUVFPWPQ7ytHQGUtRql25teHJqkEwXv/m7OHO8UYKTyRMFsAUqMxjZe74IccMXC
tROC8CFnUU8ORZLiMGq8kJ9CciPooIDp81MySMo5bPzRtAae4IhL/XdSX+MUrE1T
Dzpb1mqyfIpK/LX4eUh2tr958ypsI8Hiefx6pOfeB8kJuF2uv8IXINxlxpygWtj+
NwoEoPcbKAbCUqhxMrMeSOS4nmHFD3/MZDFpgGYryEBwZnbwWzJl1FxlqvLXh5JX
dhoeyF5AgCOUweVWdqnToyBPqR5c/a6PiSpXo7XJq+by4goexY/kftSfUMUAWDbY
cXlqLQALaadVsAq0hD0rGV6JAci2Leot3WeVEsE9SGUgnUriDes3fprjze1JUSTC
1Z21LBGkj+eDHiYUECMh4nwZdB/k0dIVWNJUtUwMtP1/wQdcsf+sgFzqEHWI1EnY
pOBJnkC1L8EwPyR8JyUll018SU8T+hmrZPWwjiseR47LPRQbs8qkmpsamT4nDSA1
+EwhXfgMU3IbcZ2JB6qegeFmX6iXFWg7uRbAIvCqyESIW0Sl7rYX1eQ16QhHMUoA
Cu3nLep4AQ/6w3/4VJd3dQOUyIinMY33/39sgo+N/sJC9WFZx8QQtAo5+ZZEKFtR
OKss6Krk+dUNhjXZqHeuUWCci1vbPTatL1B4avzAAPN90mIhQpjAw5KCfbuQH8oy
e21QSf4ANXCi7fSQ0CL6x/NsCRr7f+5Hdc4Oo8C9egjEvogf2cOeeUWYktyMiV7k
R5mhmZyxqtqSyztj3NyTb8ySfdZ4USUxtH6FuZtzpaJ/AvJMC4vnvyA1Bp8bSt+2
SwOstr8rhVwjVJkbyZVDaIHBVJ0mt/TfFCgF07IM3DqnmMG4CbV/xJBDcdhIduAS
vT9UKhq7cFutu48EuDRwiXqgyIl+4Q0jnihNFNBn8J6RI5gdy90Cx1/F7FWn08+M
OKN0rimw3A9GriwS7yLVvUFeDCJZJLr6m2ogNV8tmAJPPLin6GHyU+JBoGF4VPZU
/uzX9h5l8FgwbH8CqC7VDLlvxz3FNx33lPidK3dKGCrSpyQQOYC/wxcMylGzrxEB
I2BOOXzGz2Gq+MnLVHogWvSHgxB/CuuaWECQotcO3Xrq2/WndDb7jdu+vyvyJnxP
o40jPpJwLE4usP6gKNF6v8tt1ivfYz238U8O8qZ7pILubpOvsQhL+ED9wdR3lju2
t+Wm6DA7C9blot8IG3RnKTTd0p/KXWTYYIFtETF4LQYEhfzEMLZN2u8Twet7FirI
L8Dhq67rF6CDrEQW7jXgFsi1VW1fIFzNJYOfK7zHQ89ikkhEvrwwFzg38ybBUhNH
8/HBosgsWAjNbMJbHAZchWWNfMTek/3lXccryLxeQTIG3WwrEiuFOmdKbauDeQsc
6KsSm9vM/s1v/DhE8rZXsah/jb2Nt/1EBVKM3MpLcd0Zv18nwCZdpnWJoRT9GLyN
Q7b7C3+iWNrp5YKkskwzyZecF0A+tllJgZQx9RrpO7lHfBfdqFpzzzysspZAveQG
PmG6FpjEqxsRK78VHxYJ6w2YI98R6wXCgdnZMmifI9DnaJfx+/TZbj9vtjiR/u/g
NtUjH39yd0eiaaPLi0Khp3VVldT0nIFUUmWGC3eMfwYT8KH09UfsDrUARaFC65eD
HRvUfRQ6IhQe1NBtE8lBxIaa78nCucZvE/NgGFLYL0ZUH1PtR8kB6LamexLyoPz/
M7xGvMHtN+AfQDSXeqLyI5SqshpqOaNQux4z5H3H26LqfTBxoQgnWQRvnea9f1J1
RMrtLy3EK39/Z9PwtOWXuKd/Kiy5E+4AeE/FlY+nBraP3UjKv7JSHt41Hr7UJeAE
e4bDPoUIEP7iMWOitsW7lb0V5QpdWh6BwnaprymWP1Q2mEFdk4jET8wba+SQnYdW
WkMrCEoYUj9dZs/z1b+QJLjil6D7WntRhaqyPn3b2Yno3+l4GxHnT9CDw5ArAEfo
2fYMj5zHILZ+GBmbG632RRMuGB15NJ6uzga90C63VdHwF8+m0fCUfLg4Uv7Jcckj
CHIxjJSbOfXLXNwyT2WhlmTA3RL85phsx1Tn4sbbq7+cKZSFOKlIvKxyZLtrN8lM
xq6a2bAdDrmbHhSsnljNWWszLmry9/7UoIFvD2AlmxYW73jr5puiOr0yvS0/XN/D
HB1zs/YEKJwAcychujM9BWj9PBaACgLjGH1pY6aA4TdlXHJ3ZQz2H+cJuOKnkyv4
rZh0rXuATTJkGeJvrRF5EwnjgWdYvGVouCMRGpsUKCUCMbu2hxSBwNd7pHofyL0h
yFtwMm32GTdkWlcA1xpy4QCHkeQ0as4nzFQDO02Bgo9gC+mQ0evugG1qqeueGqDE
LGsYOYD4B9jpa6YthvokeMvfsQCnrqjHCKCtwHEvX5zNEIjCl5wvE2yrJ4Y5SFe7
`protect END_PROTECTED
