`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lHa2EzEwyYDv46oWszby2V3HzXkhMYJMcip4Ch4Yz/sImWTQvubyF8P7BuPMzbVq
7Fo+PBhJ0YQikpjEDltbZsGA2S27G65vEpqtu6aj49PWukBbdxqz8sSCb737w9Ng
FhrWZIeNSK/qBTumgnDMGpXiPKc3DcYVPT1rmF08GKGY3KjXIyL5x/NFWnfYtYCy
8RPL4v6GxnnQXQ/64mqSgTTfv5g2pnFrqyrwrjTDqrhL9fRxbldWAEafHgEtqpH8
mA80TfSKFraZXvz3FAetrJNvHOAltOxnKB1FVi5uUwFeTiD4bbEzYqtXjGPcS8LK
YTfOQ398P1BnGO8bTMktUjXXiFAlBP3dol4mI/7aqVaHqxxayanP0YygpTRoiNkR
`protect END_PROTECTED
