`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DwsSdv+l3qNq35mUJCD6Xc5Z+8zwC+zOhYphG29JpARx9nzFP36FMHAn3EBXJ8gb
fqBCGWXQvNzKRsBSXcGztyZZVm8CFQ8K/f1iqees2j7ccQ2YwKI4rESr9DmBsT4W
pCGNLSjYy1u8BTtQYrZe5DiCthGeP15/WDEPaEBchJlL3jOn6eGkdgQf0g+QVbvj
fFqoB+oNKbe/4U87X3kPFQkkhadkFePLM+9C6Jv3HdavZ9qIFwyVR7OV5O9DLtoK
40N2APau6CrYuTrdrzfVkBwIQpVg7EyUbbpnW24qCG5emXQXi8XdI00k8KKORJA9
RitTXmcO9zFPoApWYQNb/S18hq5ZMgS8glxpopDSZfAwjJ2MrlQ8qrlPHCAX+E6V
EJkEWAphHGRxWU6lrI1e2BBOhUGEnb4MNeF3tRYC3QWzNNtVPgRNXgiLk913Wkkd
ax49B3koAdNGAEgRvW5vLRD8XkbDIwblC13s2AXwANkqxekA65GCzspEM67fy2cS
tb4Vw4TqgKkydQyAFrqIR6yvau38VQO5Ase/aEaBVSaCGwVpWC9FNWGy+6FOlWv+
NmgzbolTRgRkVFVrd4GnkKP2kShSdr50yipqW45HV0FYlAuCViZIJbxfsM6M6iUi
8LPCP8KlnwSu4MXIDapJbU9Sbc8kLKVa6ShMfO0KvcwOqvYC68ZMWMsXuoz7ha6N
+0E3wLmxd1WKX+Um8+abIcfUQUEVodfFqCkejcqxqPpdHIUxOUuEmUYIl5F2eocL
dYJfBzpVH9JC1Xull9w1m9u6Vg9noW7Qi15BSyucH6I2e4HVl47IRPGyhaQuJfOU
weO6tDRB1jMh688Fwgz8gT6cbcZfovVvWD7unrNIu0EYRRmdC7DKq3U83HAv0DF2
ZE66fba4HrVIvXb3sLq4C5GsvXKgN7wG0QxEVrywGWv1EP1QUKTJ4rqtPiP/cGyE
C4no3Dy96YZbPgVsekNmepKMvY5HDrMm8bmDG8V4kxxUphHgqIdpxu2x0waflp9s
VANMCIQikUMXv3Ju2cxTUJ0yOcqIGvZus/Al8z6ikYjZQvMIgUxx8FSHhCPsXxQa
aBvryHfA+8FXsKJdBqO1o/ESBvjWTAk4AsMYf5Ymiev7UUCpKdNXAPiVh2OX/zq9
LDULCasVTYqCf6ORQI/05EZ3QCSXYSb1ksuDH78F9jgmDxVYmiU6CIlPb7zLYsJi
t44VT0yXFPMlzoDi9JxZr9fncvslDgkQddSt7d3MNLhhZsDL0GFfPx7XAbL1TgEZ
k/qkhOHmyr4TQ+mlKO+G41CrlJyVC1HTVJIwxRAb12rjikr5OIWUQSJ5uNuwvCNM
leE273GdNYv8wPsuGsVd/88vGl1eEnbdFtFAvFN+Kj8N8Nkee/8Z7QnABM3EW91Z
RCAWiRYebQX8mqoNgmkGOkZtk455zykFwQBBTwy64Guc4YxYE0rBd5l7HUyBpqEY
QrV4NAz1opF2bNq/3800jxMsXZ0pSRX52fTv1uWI0+BAJaCrIJczWhC1fO3FmSU7
AMU5hlY7S1hNNyWipzx0vXiixIJdKuu9/SglRQ7vE9RtEvbBcgReAA4ZigrbNmzM
mqRoCknQ1PV7XFMeU23c6VLrGH4aeO+QdLgAr1lVRVhJW1ywXaQvUH8S0t0ifDL3
16AWR0SzZJxu2CKNNSIbXQNEmKzcbD4SPVkdnGtRREzGGQPLhw2nOYYrD6tywqOE
ZyBLap51wnMeakYf6GFrtgbQccbH/m/ptRLZSqirm841fSh+l6nEWAsqrlIBMrnE
RMq+Vhwek9w9MlWL/oNXWPY0e4MG2G9XqiG6cPNL4kXc04jCmcNtYImuipT31yjX
LTj2mw0JoR5xeeBo0ulkeOpBOwL4DkE1vqCIo9RSHvfA8Ef6H18TdIegf3x9mESv
693kgpEOoPUkDVkEdYmKpPfy34C/yFhdMpXezQHl6Hwy1Bx27fanF3Rz1eQFEaS7
hlSBJWNH9JMWwuciVRGuGjIdSIL6ox30A/eQ8QpZ/847QXlUdtxo1RGoPucZFi2x
KHjzLO1E8o5GsfzKRyQYTZlDZyVpEuk+k6FMHJTNto1xDzrr7r+6vi9ZS6U/kV+F
x9yug6VXMLrMmvTQKNAzCm0K+vrp1sl/7VY2fcxZ75A=
`protect END_PROTECTED
