`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5qkM2KtQ8dk1xljrsK/lDjaonBNx/3HcZpttkc7s861nyv/LNmXXlMwS3mFdUFM
6Hq33oqzYnkXL1YSQxy2xJQNz3v80zJ+YxQc8yjmgQK30YYVWD2AkdpUY/N1HIuI
5VIXK8EfQFKfv3v/zcuUELgvxnVjNu6+BzGPBPmz0goc6OvX6P2GYoaqOZG9aVrU
9vms9kaKAo7LSkTMW8Kf0sj321XjZrW3q1yU4NE5E612q+l2Mlota+od7HS7MTA/
2Q3K80l0CQoisKh7CoKtTXITTXP9VNzF+96ELL0Jmg7oC0RHtd6ZAruywjp7e6O0
ZzQkWSix8dr6qBQjinBLYnLbdFNg16ENp3VfG0brbzVio6d0olSS9F/6H1CrSHx8
HrKQupvMFFN9BKpzNtBAF8YNW6RGQcIXWK3CsuHsgTYTHTe3cm9rNLIRkBYs5WV8
TQR6/ESUcRa+72KrY1a924vUBKJ6yWjpurvifXOoae0gyR0+FGowv4E1Y4wawRHp
JKC1CpJsxElUYFh6F+lp2/ubRkbpUJvRE8Ic+jryZIHugpA73JspM1rIOuMd8W9i
NCnh7qMzIZPTZIxisTNR8hWODS7rR5L0nkW1GzNUIMicqkrP9aEQ0saDJ78qG6sA
RMsjdlsM7HycvK1iTvv74vQVG1nEdELGhAVREZ+sGWKb6Qme0/D/6ztsl1UY8pqh
OCfcz9AbcyGDJ2eWK86CamqV9AgYFzDNG20yHbq+0t6NaZK4gALE9T7e2V7MBkaZ
tW4SBL6Hv/XfSWfO766grFg2ctNPNxJtsO3dn1H45K5gjlC541f7Z/vIP+3YuCYR
4UhMHWhxIQ4jAXjHGggtMGlB96iWMxBA6wR36BJ28D1AAbXo1dNktcLB8kYUOppl
6DNpQU4fh8bbWaBO1hfI0XOdGU23h0FCL3k+nmKVx6PZvtjJVLmbN1qF38ZsxMbx
xyC4utQni1uKt1ZbIuSpGQ==
`protect END_PROTECTED
