`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NaKUdOsQhGtiItCA9OWFOD1yAKvknT34Vq8brHj7dMXTV1+TbGkiGBvDOQ/ASgED
rIWOiMaw5o7J7O/j00K0M0lQBTBpTxfHm55ALjQ38CGXWiJFsvVbeYRHx+pj3ykk
9efjn/Ty42nIYfMvVaqCaNhM6+uV6bMusRVe1jrCCGn6CaWMh0qJTP7OuW0JZAwx
mNab0KzGL4nMF14q3VAIv81XjGo6ZruU7udr1qMeGPprDntxVFNPyb3KaiUUOovU
Pu/MUqmo2ioULRfpx2kVtZKocvm4yyOhPddfrAI7yZoNc2Re1iVMfEL0Q4GGTZba
lzQguzFK/75NwAANNPCS4C45TzOcHXKt3gs6hhZrrKH4EDNlyq50GT2WtQCB+V3/
jr8wffsE2FlFUXa56Y+b/FbUWOYQuolEqU/H1wUXwl6o36g/Gi1int8YW1xN6xjd
WFUDrw5R9Eeg52y3ygotMQ==
`protect END_PROTECTED
