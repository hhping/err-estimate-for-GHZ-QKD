`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4krXn4iLwsvNDJ70hVZdoWV2s9HMxfoiO1eYw9UthsRIqHhk0YnmyfXKhUU592p
ZImKleHilqZycp6XGPVnq9JRLCxZtTLDJzl6y+8XG7BHkl0pch0/JwyR2ipFp+Ae
FESaFAJ2w0GAmnfUOctW4kVBHrk8JNlsib/SPLZZFG4aa/XJzrugqKS28I4bnNxg
0Mmu1hIgOgGy+Vy+omPQ4qMR2gkpBYxjl3voiBGCmH7kXTUa0uAnDWH65grDBR55
o9lD2Bd3jIX/IOD2Sv/ZSzngJUjUsPJpHW4ylqfhaBCvS+Lom4vOSQ3/dl8u+0ye
jQxH7QoCcWyxNFifJphYmX5qaBphUdN1mMiJCuLDmfuqRw67TVdGr9BqDt4C8ao6
tJWrgRg5isDsIRpMvggMKyl+WWnKLnO3S9uUCkhJ5o7c0672AjPRkTfQNfyeGZAv
7rivXf0kErOLo0Y6p+ClU2EMgar4Do3tmM5QJ2WN4YNZNL0Lw3nre37qWHnkxl3P
pZ0eFijKWXd/zwVP2uhKuzi6Lo+KJ48oiB7fnRCChPplNMEFq6fUMel2mUIukLSP
7dGjU3e1pxaQtztRTKcpxhv2dQGSYjgtVLIJaa5d17xkQpNVegWWxpMOHhng/+4n
Yo2kGVogWcNGmTKx1cx9yau/xz+B4SO0A0osGT14RrL6U8VZInhEQ+EQ4kIoY6cG
argrLXOO+RGGbb1OrG1/7cxLdQY/LkHdhLbOM75r++74psyQVna3dpWHt24HTT5a
Ugjo/40JV5mSox7E6cLJgRpGXEqMWJZq/40GGtmmi/AziefhzJpbmhsjSPMDlc0f
0LHcrrgmh6qEhV3rO/IDjZzfM631ijv3p4s3NjfJnyPwSenpcpkJ5fAx35cKbX2v
9+j8ywAiJv8QmPaZBItb4xg1J1P7YsnEcDRT7y2YAk/b+XrH32krywaGkbJ7gUDF
fwDIt82lQl4kGoMvfIijGw==
`protect END_PROTECTED
