`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHWuERqmy8s34KJzhIFX390XRsXIcsPYDFMyCICBNV1VDMSmN6Ty2qQk0o69OavL
fwnQrmB06x474R0SugQbWQGMQn+xIhQxBne2d7NjC46KwpDDgH20uhpi4DsWRvW/
m1hNp//Qu1V0ajYkFlx1gi2yvMtsosVp2+VIDaDqqzGqgt8i5A2pOJAqQkQFIVSU
YBn8FF2gEtvpOpR5556uZZRoibjVCxs8xIlw4p4VRxXqSg+KXqXvVxpyNSrnWjSI
8RclVkc2Up+wD5f+kgERajeg/iERur3Vd7V40v+QtlzWv0I5aY3uYFpF8nZBC/9t
SEWahW31X+EqPIO+NKxOVT/oFTMEzgelsxp9yq+/jQicjy7dDbTqe1GP8HTsudI2
FladwCwn7HbW5pFD/lKu+fHRg/ToigvIN677zPnA2Dao32hzcECAX7MerRNesa3K
cmAwRbgU4Z7e9YFovRH/Pqt5TGn+lurua2F7cgY+wKq6KTZRmfaJriSbV/0nx/Ic
nnDp3LgyYKJsbN+w6qD9uRZOTk1sTQrTyyYrle2WpUE/B7i/8Wk4TMX6bQy+bE/h
O0ADO0ryQgj/Df5ULaAfENUJW3T8zpMWm10aYLthPGSuDRlOuavyaUjebP9BhOsD
U8sb56M+o9fvhb2QE6JqhRtQ6yJvDKCF5KMcMPO5RcxKdkkpT+r3OfxDSMTsxP5G
1tprtgrqZKRYxwTvBGEU3gVDC8DEPPupLMss+O+1UhrE/RyLDtpY9SfcIoZo7Y+L
oQlCXgfCpOVedYxOaW63EixTNl75kZ+evCPQcCA2wQFlMThtIECcb0c9xURqtn8k
9lCmG/zcaL7mf9uy8t6DMR158xmXhut4dVX0CW61s02FyhqOSZx0rc29bGVWTUw5
ou2w2KG/ZOmUiqKSQ5Fp9oWiuEpmX1TZy2L6oqyR6GVLVhIE3CsD1SZyc4wrQi+J
3OjAL4Sj8Fc1HXayw1XPhzR0QxusAP3fbwq71Rr1f/0iT+a5oIeLvxr6aSS/tO4P
moK+CCtKHWV1cqMqLfr9lUxu/eFyEOuLW8zQNYhkV6IT7j06DMwAQlSFPpvOzEtt
pyA1nodc5INbOJXcIZlBJ0zMKucnrCD3+3j/NH/IdEt1sfJ9833TScsMn5hnBpqS
37aQ3rSscd8HMIBK6AkopBE3qhvAoSo6vSfP2C9vmNPZg4GyKKZXeEkHGXuxB8Qm
1B1swvQorLhbCwpg4NBxki/zBhEgHdZxVkhnrg6Uia6gQbHCjPJscNbV+m/1lBTp
mB/M+RDDQna0YwD68NvZPc6d4V9K0fnb48Dabmiiikf3kn3xhjssikM7c8hTkoeD
QGRPyiaEJU94t+UOjZHvwXXwfXrbEAs8FkavObx33ahqIJl1MPcRJtQ66MPxqxsm
lDpggF/D1XyZTx+g3BF6CqLnlh39Ar3aC9JuIYCWx8tGj/Xtm7OgbSXnDUnDVWyR
udtI2pgcAEhY921DAbwwyhBCw1CZSJ7SU0cl+QcC6seOYUNtzVJJslRUcL9BufjD
A3i9wVMIBbeGmJtBcGAAT0yXWAZVzAnIVfTMNCTxxeDOgOm42lfcGeWOpA6Nwg6K
cX+AZCBxLGz3ReBaelY5uob31h1qnaz73aWqCRm65STHLZvdK7Tz8XckGERhksQT
C4cwg4bjpd85dDwfxl2LzShU42SG99BzUc8EO9XEmgt1jcwfRh5XlUJ5wB0o8eoC
vvTfYysfYr6Y44uGUFdaRZsWARPWLE/hqa2NUR0C3ja5DoGNvexMMi57jMs0kg6Q
4MDpkWFy5VIR1gyDb1qhLotN7zmLCpnt42AMxFcif+XEuLjWuOEN39udfz2rpo7P
4VyA9hH4DJDzGQu5QTAHhOK/YFOaMO8xhgqLuJg8gXGqFp7P4ARNF+F+HQRa79FU
`protect END_PROTECTED
