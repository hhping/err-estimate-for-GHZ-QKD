`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1RVenLVF4RAYRuBNFwHE66mHkqmzPobxVLLqKrJnrDCj+bPskgESdfTXpV5WI4T
JIpkkWOVX8hCWbzKyF0WJnsGH75ikby0bXtEKWoU4IkDOtQ2xFLUN8sjmui1dr+5
hkez6h67MFZgIGSL06RAzw8IuhWBPSpsDL6bGyFl2BP7N4S6FJ6DzwjCeCmPpjrS
sgYdohIBGVNDM8guR6/bhT9TOSA0LyCqfen13uWzjfvk5sDRqAUpp42m7W6FK1fC
CcoJ5a0KH/vyEMm0JBDsm9JBzc2XvuS8xaO0fG9KnTF17lgH0gKQoAaTCrZ5sgWL
mpZmTZAI3DWjQ8Yr2bUAMh8ROs7B3zEcKksucPcoTDR/pJJ5x23HxLxMYmqDmJ3U
GReuNOjRUkKHlFnkqPrM+BJR04WBZuVkR1pbG9HEdThmvEe68aWgSxCAmrlSQoB6
mqhEVdgmfMhDmLSar8JXCR806Ql1ix6JyMVLNYq7DWXJTF2kKivMhG3Kei1C4ct1
tlqqlVjAljvkvke8tIfPliWClLNzYp6K9m4K9dD7IjrX9D9fIu3egmcxD4AkN5hC
Y/nR0BYOhGE5HnlUgeAy3dqWSv5yRGcqMFbj03cQ5Z8OjQ7fxRwLpyljPofspuRP
T0knLvj1s10rg8vOk54ZZqGFo/k2qCLmA30yzn0PEZOsp5ooLmiQ7f+9jJMe6iLr
08KeHJDhtw8QuBnBQRb4FUmsX6uh8uvVUtcOTdAIfFkvEVwN5EP4Z19frXLMxciN
hXVYMlOyltpoxg2UXED8o+OS3DjKpZvdGq2AcgLCLsGMH58RMQgit0DurhWX+jsU
PILtmqEVTYBJHHh9hJbpuhNEoRotabCwKEVe3zs9+Ik3c7XJGFoTTTpJ4ChXCKsb
V+ItcwtopJ72gRZvD9GcuZRLRQFLSnK9fzoUwgcCDbNe6u7H0ly8SSCpAtGuRYrD
tUvDv0XDqg+e+m50Ed2tF9zIgws+8Mjj54EePzEcfSk6t8wVx5B9L9cEkW8K9XgH
bKtwEeIApnqYfpquUooLfVGxXZX3JMU/87FH+fmadj+e+7BWUmv5zF40TRwZddfZ
dbzanu72CX/hdIyMmX7oYyBbfw5wRUnTz/3rjd4zyclGELFvPxHRcAaiftikkmtM
xgsFzh8t581vKnEJrlkYT0/ocXWjuPsB01Q0CVBbVs2InWeAhohNDRi/A64/ZQmw
k8S+doA4z+2KdiAJWM89EJe6dwTuwSsLl7MSSgu/JD/i81/yey4Hw6jZU0r+JXgW
GujtSSIte5rWmLWBMiqcSAv+G7LyFfjSsrDyZfwxpibGbuFskv3C5RO2iogbLvqS
t+gExODx31iw1AukXN/quFD+byVvL7INla+ANdl8ZMNhNz/q/uCptONyftJrDkDo
78GpXuUVCgDUKFpVBilL2m5/bfZxpcOIgy4A+Ja5al/hFE50sNqA0a/f0jnpk7eH
oTcNvb0MJw9jvyTWvhim5LwrYFQmdWeu4RsD5aB1gxfQTHd860fSVNBmkTT+I2gY
dteC8QBdNIU9TykW7HKmY71HaJFqh2nX+L376XeyzrKsEm/FSB9npPjxxUWkv4eJ
HLj5JXXarKaEGRDKe8xNcpE7yKFF07pbO0cXAq/4jVS7+3uvTN/Ypt5biwFQsrlF
wh2r4FfAlPAVOXYsxrKC2u8L0Se485JAyFAj/dvQtvDaA38guVhmASYTrjgahhzn
1NZwAm64u2MpWVBIKDVK2e7JpUNcvr1vOl+/aolO98wMzZw1gMD+NoWKg96d4UUp
kuZO3QmO4tpMhvwjSyYBlTbwjwPCcflSrHk22ciBgttpUi/hxm892BcsEqzE9v2l
9K9r1JeBofcqe+Y81AdK07ggemlZ6j6jArJrPOZdZ35T55TJ6G07dEBDAmb0krq0
P9Ah+SGQtwxm+nH6zyoQIIHfAeT/vZdrnS41VKRUvnD4Au8IYhG4puQ5g8xeCqhk
zIny+CKw6Y1eOr8YQJ8RTYCy5U+HzETzMueyJUbCVfpWl+zLnUeH6L0RuhlWr1+8
B/U/IdqHFitpAi+Fh5EX1PfYDDy4AyKs1ixx/F8ZCfOnNuCzfgU4BnFXTck1Fom+
C+SIweRwpjgS4qOwxvvAFKkSRVvwI8L4yTP926scXnSCvwBSX4scPOjiOB+dWzsc
6dUi2lW6jJq1fz3c6YaG0cCtiKHQt4q3Hwek/PqhbA5jVQVT84qfq2s6Uvh39hWh
bSAMFvxSauJmIMIT7b2JhOyCo/K7vNTfofM7j14rKtuzkHc4LpmH6dZj2ZRK1IlL
AxfxX51ZLeHoEkqgwdXZpKNxea2pevwebDCr3sFsUE6lnhAjaapyuMi3fLYort/8
uWo7lerGd/TB66g8xIo7EbLvxZvMXZh6Azvgtv9oIDBHJkPw6p+Oo0DP78RqeUTV
eB2p7K7vWrPTh73xvtWjt2jp17yOvLtQRVk6p7RjLGsxGXueHELnCZLIrMl8ns5x
eQm4o8SgVprY7e0W5StLI4iUPgBv7pUCOpypmSgTT8RAYu27SFCKxwpty0Ia8RDk
8q/uBb0UKqA3EjuVg/w1OvyC55K4ZfWp6oATUW5j5d/ncP4tYSDSbYNlAoZL3Z9O
7vR82ZZePDB4QY9YQuHCR3zifYOdmNeKia/3s7RP6NaWGnucvzkiM4rVEQQ0g3Pb
Nf5olhfFHZzQEOTMgpxnVybQGh6JQOvZ2/UFFy0TABrXg4KCwHJVZxa2z4wHs3Ud
8SmybnmOyFI8o1OkdGnFAN57Bh6wd0NGfjFnyJa+1zDBD9cgyG4hf6A7Qr1nUGcc
gxVqmg87NPd8bLDr8g5MbvpdKzCVErYoqiCuqYZC53vODMr9JD3juq6/hlSo0N03
Xmha3AvMquPxa6giXx7iMEDNi+knl3bGqE0E+LRJ7p7OGUmEPzZwDCPh9J9QMmI0
9iPU3uVd6lAq0K7W3JfRoJsc6Z2RP7mwJJQOUhVP2nrQgqGyU8BCr8d8Dp8VLbY1
wuaBfNV3kSRRdq5tqmcTV1PPMc3uDLp6x/WowwDwCa4xP392vUN1LHLpwch2vHb0
3LAzy1pWa1NuBw3QcxGjP1L1wBveqFBk16UhLaixPYQb60lj8n43LY5W6NSWumeU
idVHRLZELPfEoP8LElxil11YcF6Wbd+qzWlrcrJQi4pMNY6M+INjfbVFnmablYJi
42+fk9STsxA3h1+s8F9gsAV52w+HrFeNjSmvVrt5L6HwyMv/v47gB9sx7iR8uswP
KIkpj/5wobDsHmRC2yR5rl5IaQODUqInhYLyGu6vbRKsquhZjDiy/REAyBXe29n7
ZbLJYfAGcKaLWz9bpMyph1+yoK5Y5XlGInO+Xm5L1KF/zrN+w6mWzi2UXVix7Mzw
4mF0EYtzike7L31P8Njm5ml1CUZYSXDv9U1qlDLpLKhZ7BXRR5/GNqLplLgcbgnY
e2iFhDw9cmv3ThTC8sGOjLCM2OIH726ZkDflq11brgdm5yLF0lolL+B8x9/wdEAn
f1ncd4AB+8ZZ313xurcrPDjXqNoD+8soMH7d+Fhm1kk1P3KPOtEfj5eMRAftI+ah
oMMkjKAmPJqg2PZmbATglKwTqJjd9dKOVBKD3gdjgNMuyn44vqkfy+NUHVGE0lCm
Qko4uQ1OB0iqGXmxwkApCKFwfp//E5gMsUpUywappCUrZo4D8d0UuHJl2IzXU2zu
7HrYC/HmW+/JLAgrqmvrsvUWhey/DDco5g8muH7AB4qpAStCB8zn39tU20su94RL
cMc01RztsgX68ZesnRkkOxQQ3QEx+1zDe0Rde3FWkJZYn5EmyhGbMBAFSEvVzzQO
5o7nTE6MueX1G4sQsIBR8N2IlyfzAz1x2h0YguNMogC87zf2iWgD42NKmmv0KjMX
4pCT9cNgMPkLcc/SSD1k9RAAdaRmjG16i8X/E9lISxZIoB+xia1GxCkbJYAZv2bU
/wq2bAmF8kltiu9wXffwibbSnsboAniK7YWWsiTYB20IeeA0r/1JTXDkBeO8DIO2
/C6UfR3erxr6zRaLnHN/XscoRcB/dmdMSnmfA98Kk/EUzSr5h7kXL0wI4V7SKVO4
uwSQlrE0Ke9pDxLG+OAVmYzfr7NbtsVH1L3hxNX4haEHrntFbimgJAFgZ8uPgnwx
xQKFxDNVOHARhRYQ5ImSycSfcgwHZChPAYxDi5UCulR7d/X/EiCjDI84OKNc6QFL
8IXjFREw3j70K5KRwEQyJaOGnEuTmngjlAmZo/aqAz7DVSHl0AjbGnuDIHxEpL/4
fDiNcnl9Q4n4jrMlsl/3qnpDVg5ATL3C/focdQs3WyWSJ/ds3tb4G5UTDX6wU8//
gjODy6mYLgv20f9PphIDVDWy++mlGSb3UndwCWNkuCp4iLBo4H3a0MGcOn4W8FGx
MgEgxBefivAlYBn+8Ganfp9Zae38FCYbih47JqVLxL4qwflKFht31IYOlbPYS8wH
sTIAuV9zhhgX7WkJZvh8FZwm3JpbR7EgKKurrh8/6oJCdoQXGCaoN4e9PzRSad+P
DQVkpZ413uY/gqrKYlQQsq6Nlgfcz1SM1ksgORrZHcGr6EnnfNQ4WlWY4z8JRNre
EpDrF0oRSPv1SqXkG2nVPlEHgGhT+p8MGdSjMT7aVCeBVyFfX4u+tsMGZvvHql9s
74GVZYayF+66OqHhmGBdyY7lfoHdH3fzQOxsRd5kOpluGoEhLrKxSFwqg5rci+A6
bxd3m5tVNqUrT2j+Ql6hFBEk/fJcLoDWLkhgP4+J1T4=
`protect END_PROTECTED
