`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24NdvATTI0iWj2HrjXvLwyNSSmx1f79xiNunSKjNcx1H+4Sv61FTco1xhbaWzKLR
KRH5MLe09T2fEl69JtiZfMHfFt80X6vlzTjCLZyABFgrLv0BpKfpGY/algAwCxEf
kJkCum3rKiwk/ItvlYHWLE64Dh6hN4cqVRvc32L/S3FtQ1F2gRW9qPmjN8yyITR0
/tvChajlboXhiMa7Vw3ui/y11fj/Ym/Aw9vgd4nny84gAJIYusVw1+qgsovJkiuC
moeaDrYGVJrFVrNofjL/aMFPMGg6xxsS8p1VpXlLW2f/AeUu6R2/AC34oa6++mvb
SJQd7bmlmMnim/cbD6EOfBg2G6H2RFKhEv+El9s7NXyVBevsUpJE8+AaS95TL4zU
liyy4/ddK+KnIFbJlcIlgoeRe/9ej1w6qRxrVbZEMDCJi2eI2BuEuKKxU1pG1hck
iiCF7V9Uoqs1oRMlpAeB99CvImMLKi9LeJzrEMeeW/fxBgPCMkv05W/viCeQ9wlr
JTiCayf3FKWcewRZIz3ey9NnxnO5JZUhW5YMTtM7gfxN7HicKPou6/hFdoaK6p4X
fpfkH2teFDyoaywkdMRU0whi6KWLJrxyEm5gyb8Se2/qgKKAQcySwXM4sxt6zTgb
WtjrK1D2WEn3qZKnPTI/SjXZV0F/yOvGMD71xxtbWG1UFlbOgztKvH+o9JX+pSoh
8Y9mlxpoeU5wSJOkGlW3Ito44x7AKwlSxWMx4+nlVX/T8+KKd1wSLMD3brtymdpO
cyiq3F8WqPnYOUVlYf2IusvQYb5eQxYxihOUdTdXXk9oFsz3Gv9v0MLKeOd8vxvQ
RZ80jQrZ6oUYlRoTcGv17YOtoyjN6EnhCva96ua92GNDIQIfgNiOzFvKiYZh+xGp
hp00vzFo0B9PCGbqxqHk5rnzqLWtREs6dy9UU55Uw9Ua7AI39j6aSx0OYBk5POc5
1suOKacwTP4PYfYv+FiS2GPA8P02ryhIKrz0MbmHx+yimm0UKTBxPD+V6RASzdjf
2oSpReaJZrrjbkfiE7Ah5zAU1QRVMeisVqLKJ2ouiUnel82zndX+BvKJOf9HqlvE
G+3CUDNlcE+4Ml+FGTeC4BnwQSwtrhaU408hKOzn6dZz+zbDOEZG9G+W+pYRM2lT
PYA13hddPBJm1UxiyhqCzuRYx06iY88eaP0fYBL4R4fMS8TzaAblLShAOqv6Vtyj
PiaU33ihpmSRhve6eHvlG2YXDLtqMqvwI+6LXrjhsi/KqmQUBeSXmSr2lLqEZHIa
urIDXILI7JJV/WJwd/OI/Q==
`protect END_PROTECTED
