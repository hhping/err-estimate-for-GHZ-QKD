`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkscFU11fsW22gK98yKXDdzeWcmhgOLs2JBQsO2xsvtYiy/fcKYZJcQ0OLsQZ/Ee
b/9JCXJ2WaCqBz+r5k8I7lvWhK25X1HQG5NY6r+7IVGDxw4sDMvwtEyOBhSwppYO
uNDO/+3QeMg/stXexjmReMrc5+8j8lJ4/dxCbeDsiXU4wL6MqKwWbQ0Ch9iHzrPH
Mkh+Qsub0Of3uYNlAjtQzoT95v2a8T5Y82PRqoBEnCnzv3oOfuPRRkTyGsvuul3U
yU7hKvJB56/Xo5tpdl86BkoOlDe5vBz0o05ptHAcWeMVs99q4NE2NHnlEp5NVaL7
ytM0AgrZTZIkuyGYQr6RoDeT02UG6Yo7kZFJuvIr4yuxB7lSPlpavem89QEGXMiQ
p6848eOwWx23BKLYxFnlA/HPDmmd26XqJLg9G8riJuvfYMRI/jI608tH96GpIpxj
5jyEK89O1NQPlwIjQZNe4ZUX3iezPpZamZIGbCuvgdOgCxeHXIQD4aqIzKeZPu4L
znokH/vmXre/3hGK+ALC5DFply41xKplTwnAMzDzhbkjOCa5jm7peFIFpOrKfc/f
71fE5HkuYA5XjadgkpSySxVfQ3Bi6atkx72ueKTn9y/lN+xnXtxFJU1Dzke8QtuW
hPppb85UPz1khq10ymnNqsx1WkhdYZxMi0dXGBLtmseNH9xtKyyhNV30baAWM8Q2
Tphswpa2igM+Vd6AgwbbyUtDkW3Rmd3EJfRvbmF3sBJAx/gChNyIxmYVpYF41OTW
E3ePJvioiW3nttM7XZqF5c8qTDEKhu0nZiU8xWAA1C7IMG3V5x2f8d66qk7Y/Kvt
eipyHtILcfCldSN+PFPiVRL9zEY0mEgUd6Rp44NISjfOioqp+FfBSWkw7lEM4icf
XZNEKAbuKGiRfVKM8iTyYN5fMGNw1YA2FiLQcoY0QmnbwDj8XTYJjCHOupB5vxCc
MW67XbJ0P8BKY+r3nqiW03d4haNr04Mc6mZjR0hgq6fLb6VlonEzQV2hDNpamf9V
pBymhCb1+iijOz3OPlqMmuuUv34OLhSIXllmtaTK4t8CyYfKSMEXwYhAl/l1ND14
+3Cwrt0cpjmaWwi7IRWYpNHnmUqn4poeo8YAJAHJjq95eLXE4pVIsL6YyC8g4IVd
Zx9Ho58mmaM/syQfhN4ajGV+MICWFJyWTJjR3Mip6EhEqFrc6prqBWywtAPKNB9+
icU5HNBsVSy46Ocz6wmvT40EXI0DoDQ99xcG4EeoSJOYWoZYVlfE4Bb/g6EEgQy2
e2ktC+KIc8+X7C4krpssLA==
`protect END_PROTECTED
