`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SR/hSTyW3JF3E/s8Nzo+80IvlpZDei2MFlKQTtBUkfk1a9jOAgMj0byeEZb09+yB
+TVJ8th2x0LKbtcYIRMgW6BpH62ckNIv/Bh3NH6EYbzqVOTKqdGvdKW1Vky5AShB
SSnwPcLGoIANZ5OvT10OyU/bh4MXqS9J1JdSPkmNCzemTTgoVqlZYdqtwWG/7V2a
NJPHSPWM+N4NqwJB6zUqPvOqkpI2P3uNBYzx+EqwcXMucuFaO54Hl5XRKMp+gsNc
k/WJkL0B9htnMYEa87Z4Ze9u3hnrjkuXlNpB65QwtIrg1M1ENge6UvoMN39eoBbh
rH9Z7NB9JHbi8omQun/Z3o3iiYmCcGaUXdcF5TNT19SlsxLVOiKptggQrwDtQMpG
El1Qp3nzSVN73yMXys8ToxXldqE/Hh2NtmWgyFnpNO657Fvsy4apX+vCsWqqoLYy
JQmpONcViK/aOTBU2lCj1CHSyJHIBSNzpyzO8SDrPZ73qXSPy5pCeo49pVVkTnR8
/krbwVt6MfI+pYDEykKEAUNGTJupKi6VCRaSLeQnd5QfIur4zR9ZqjFJKUj3TUwy
4bA6NQ8yUNfER0M9dPflQBzef67gB1PnZmUYtb2CtQMVpQd1xFrYiGFwznVq0y4G
`protect END_PROTECTED
