`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCL6raSBrm72mavFPn+5+WbwK4WxdcwVrWK005RvxjHc5iI83B7SOH57POSWwGg9
pa9TrmGOHr1qgV2RJubvbxYz2tshyg4nX4hxPxJUTP7DRMVOvxggPGCIXe+rcaHx
dr4I0flaxaQOIXhknc2OVKkC0Y2D3fp4LhP5BF34SP3Za/4FhNNyFgEHrdMlQ96T
vnasnb60gdd6SA4mAD2dIkaWODayw8BYdyeobHGbsRlTNi0UBkIZ5YCMMeZZ5Zne
9WrXTwoZZ5Gs8BOQwAEd5+gF9A6VBvp0ZVk5H/50JXKgrI4TlXtMsL+E+hzCV6Mt
MFqKYJBW9NRDrLwyo4eTElAT9jAoKYIcruUo2tplSsSQIuICa2N9DwRckbV0p/66
X6O3+iSID8zxA99/tk+d4AgawtWjMRHEFYPWigukC8cM5kjbfFgRsAAKgKZizapy
BJ2CrX3xOTCO/DHKis3ptWzQx/wORRnFpy35V+atyIi+800S5itdfOCak/KuGY+J
aLOJjOSGR3XyBb+eGsyQ3mZhvSUuw9tlE6ggA1XUbeQkDyILiNgQxGeHNR5m2MIC
eylVJmxOgsiLt2ZZbZq0Nsj1ddz6lVxZ6W5/q8ySoNpuJ8aDJ+CemPAyrUV0+LkD
6zgPGnUfk/fIcTT0R8BvVesjvFYPUbdqQ8yYFHt5GJ4DkYj5xuXhoXJ5FvZRInk2
nv5vOLK9CIBVU50sEIA2SSewm2FvvgRZyScqiTAeaBtK9dXAbqSlM6ZxCSA1kLPL
/MyGi5JCQxCw4UpLK4I60Tg1Gbqab9SnROCeBVoyy0Wqxz2j6Db9asHGrwWkHi+C
FTlnv5zDMry9RVcYlUJsUUqBImeo4SpT975060iFonrlt3YHl5yDj59de7y8WotE
9pUC3Qo3YynBv7oKqWJFKuZ0eppan/fsVH94UoqUh3Z/WZ6RVHLxrGmL9KFWILhn
idTIjZ+YySUWghIH9gM5JADbTFZAxfrAQ6DixH2NvzTF0wTI/e2EofsP8i3fVIrk
tnN3aVfiVP9qkkP/dE8uEl4fyEoPS6IRsGSZjmJzjX/S1cPR6P54GrVJKqH3r6Sc
jda7vyy6dlw1/XmAQVM4KcCXdFGrnHnutdj4r913KXxUvPPSAH9C1YcDXkD0tRBh
eXm4Qxan5yItwYx6b220B0tYiE2bT/NlaMptX/rg3EgbRvCi3w141eZHLyTm6fjq
rcDRYn1XrbV04HA4693gpGkU7hPbYzzE4rW5xTVfAp7cr0yOPqf8pJxlTmwiVaAa
hy6iepMBfm9Emi8yN5tAqtk9hjQGLNI/jYUN+QTgmDAT83VU+XcXV4JsRER4+SVa
10U7n+RQC6CoyGfXi8rqXWE5Lpn+U8HX0aSpDkSLwYGCJQ1h38y9zmlIB5LQLMPn
JUrc+WHy93F6T2HXMyCfNpjPZRmmJM12alvsg8kQo0VSn08gk6EJVjUer4oizEjR
frlBLmxVVD/DkFVH3mUuDcGzBbJjpngwaX3o+aiqttBlLcbIjexhLcxbxPfc0ZeN
9xJcZZPll9/5NoTEHYH+RYk9hCahqgcy+vIcP1lTI/GFkPrUvR7fMjsb8MVwqSbV
JCR8ZrEkZpLTzcolYSOuH810Cvh9h12KmkeZNkQ+CjF+S9pJFl04SsEjKJIEb9xU
BVMxBopy3jl3nm330705ORma9MLViRWuewrFSQVEYQul736t7CsWxV17txmHtb+c
ifKAIb6r+U97ZcbEBjGY4w==
`protect END_PROTECTED
