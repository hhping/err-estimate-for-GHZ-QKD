`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3KbGdN7AyADaWU7wXWon/mreHvfq8S7XCfoYY9OudLopb2j81WyOwQYBtywgjAo
cATn1rcvOrFrEK1lQWNIgTRZprK/hBBSThn+pktk1LhgaXjOlGU81oZcKeGWrOCW
/JAlm3eqUGk5pbIOMEx2IZGKGHHP3ZNReibMhopZdEEq+8OLfrBg2GiUhYLLQQGX
zaCGD+JWPtuaYmTVAlD3TvVdQYjGr6rm1JWITySwDrJzjMeoOyaEe1Te0nJdv5UX
aQZLvJ+ZMaOydEQIJP3bTjpAmq8HEYcXzkB8/KBdWvpBiYqwgDc7lL/bur7x3Qo5
3b56UHlCiclMnI+8kKUwrdL9n2LXMvt5g322cPegDRKe0dhbJz5nTzG2AUilPzzE
KyUZPc9xsGo7UsSjlThQATVF2WZlrDI2ZdC8KlOJcHqhTWl+rTEZvLI3jDca9387
cGnvzep9nbRKJOL3r4+C0699b5GMZIJyqc/U20rOvO5NUzOgPGDBfjd1vxmOlpZm
OysJt9I0fmFcHngWkO8CMvlS1P/HVlSr29qCnGLc5C7xAWIAgVTiOMZfyR6zTN/l
eOhRz5mSm+BGxRwO6cVA8CZUEDiGJIwtPBSdiQ/T+khW2Vu0dIygId5GXDsv6b8a
SBLd0m5UxQJGHvaSk4pliyzTxuQpqeMY1V6/dDNOR9SddccSbTZpZswG/mVCyI9x
18KNTTttzba0gkv79mIpitINBK7ZlNDuQMHB8CPCw4kOGpFH6KlCejQ0Cs/+dxIZ
IgsJO1HbFmUsbvuEypmwzUcKB9alyBiobFikdP+fntdTZ2HjTnOVaC5grXdu9Y6t
ZDYiow5RhzH4R+6PjHRVwLW/Fgd8M8aJNxbe/nPyM9Sbpt0teMxgmKdaSzGY7NQP
YSeG/ezQksvY4UI2e84y0Gpk4pDbX6zjMDK7k2z1N0Jm979o8qjVZe8N5sgGPxxY
FVS8hVFIoW54EE8eQxtbzK6vx9iYK2wlXCcTi8oA2kwG6Ihzw3CU5GlXX1//1qxC
xZKHCdNK5ONAdtCeCOJzcVTway6BZYZIVDBaTJTF92e9zLucmlbYj2KdfyD4Ci45
xzAG4mIxa6Jnhpft5V9MR5bNqmqjCnavy9+ArI6iXCMOv6YnWHMMUSG4zY5ha8nU
/bxmI1Va4G1AY4WAHXbwl72oY+U4nlEnWIKQvUMqW78UlLzR6Y5KMMfh/vFIlQSH
2uhaitJz1d01dYtRx8oVWbiCbha1ImKaLmzO6EvhGbrySKA/KbpQSV5pXC+J/FIP
eKgxfj8YuNvyyX8JmZe52ssUXx/kymrNj2eZRRYRIIRzHmKoQySrPcB5SL9Xx63e
0b3fSk10Hmk+aDZP50Xx81eyWieW3AMx+DLv9CgEYp/PWvMRKFKYL9hxHaHb1J75
bGTrJZAfOFAZlGO3wlFq1dWH3GJ+aYIDlQb25JUbrtwMCaGl49F7Vfv0NvEKV4FP
PJJMxYBdJzDS8qbRgAF3XHEDaGXx5z7vnsSShBsRTXBF/6H84yr1VgHWCo86hDFK
TPN+SDmV2+7+Phuogy+hfu76ny4dVJW4GAsc50/gFa5GC4HovRjUQPTTd14k+o+M
sITDV4isFHtZ12emsdzZprpC7EhPDJHhGak61KPYWPygVMFbWVZ+pi7edFFVo669
xgPkhWADLgySG4foK+HVVeS/5geDRYomqRoz+omjCBBtH1jc8vkr0qeQSiDRqRvG
HOsOUln/BbxWi0J+Wn/9/P2CeWkuR6mTHIPKC+WEFesFD/7zse0LO7LdS7XVVIdx
l17gn5njXfGliAWPuv+ARbrnEypXrMeigNkdVgPPnCRYejHaRieZT93WmTTH1pcs
EQ8sp6SN+1cu16es112yBGyI34r85cTiuwLzcElG1IBDcotg0B9mW1q/gpkcm1FJ
ksdHXcUcZT6vVKc9WwPobaam+WAvnGfwGCWBNhHLJIsA8G5gDu16StoZWPObc4Po
sP4QxP2OrDKf8licNASv98BvTy3so+ty3eQyqwktHGPQKKVNposTvnMJNdfMKoMT
i8aJf8Wc4reK3msTmh++Xqn1aam1r2FUJMo5gxhIAb9uX2eoFy+K+vDLVPeuiR5s
usJRBlPyq4x/lyJ+MmehvQW4/sOdR1vhm3QViFm94ncwm0nujDU9Qn5b/uCeSqYi
IeJznWk/uATmw+qYMGD/3WcFENlax6brH/QakJEDn/CcGOwzWTCp2v/HqsyGZbyK
xIAO0HqIP4C6YsinpcD5OsPtEPJNWDP+ViMJO1OuBSJ//ibAxoZu7tXAMTx1XQ/D
SHwMvKPfaMqgRHkmlPimBQcykbRns5o9TrDWz2UuxYoQxsIluNrw70Tz1QRUTAWW
2Rk44FaiXvWEIRwmjgFNMTOZgjIC5kiw/vTqPoLfGhjRS47cnKwtmuCHPAY2iFhV
zrzDOllV8iT9yvybCFPTMFJv4NoZqfi5gvBElNlfWwj+Mt7YEF5g8mxBhXvsj+Rq
vAh6LironEJC7OkYtwf5fJC6lBTAd/FoBHJe2BYYGKbVk3FpNgjHEnVipez84wbH
v0mdnOW/TS6MY3NFMseEqWsQ1W/On1fCxrzsR43NO0lKgiYq3ZryzAI/CUh7S9tf
m8emfXAX7tSM2aIcDYoAB6kD97YnYSA2hrFzmilE4PxeyNaANbT5eyY+FQ/qhYnb
jzHMYzaJuKO3iSOsmBQIto7B2gFh4jKs+7aqyKpY2UBxU7+PIQOjHb9StzA5a1OU
BDfCeGmsoUQ2ewnFcrxE5gmiQ/upoFh/fBkDvdzLF426Wtk86H4xB/lIfJDWVJN1
KiAW1sfy7QFkSfnr+cSikJAYSGUm/FpTtIxOSIcHhY9Exe+UDJ9ruJ5cXcMd0m4B
nY+pVgDw6KFwLhcsXXEYhrraihpFKb0KTPzEB2IuP+CQBc+oDKcq7rG/FTN3+n8U
ZHbaa1M05OlSTkCHNUGx/kqII4eTCm0Rf3Q/f9wYLvlVrWAjauI+2EmAmNqCFSao
CrPYZmno0JaDfzT8TfWzgc+5ZXfRh7ovM+3rjXfdPEaafuJyXOik6u93DKSMQluU
vfJB/gZyDT6rtagcBMuxQn6jmwO6Vsh/IRDONx9/2Z4VxRifiEfnc9yJJkf3bLdQ
LAIWWNpdEAbU1JMAiWsPTvDFg8d4+qcVdpRGOCYDWCNFqaRT6KPtJgbimV85ClV+
bjEIhW7QjX2gfJ2cvmrwUlHnpyiFlReA3kS0vZnsYK9HKneyie6iwgRxUtJ+QZZn
LwIh8TyralVAQSvpX5K2eeE438P3IbRI2xLZDrsu37UUoFNaqOWuSXRId8nlIdk4
u33CBHeVVc2ualhqRkaYqyGs4E770pzBb5bzelaW+/Kvk3NoRkjoDzlWGcvS90Gi
cRjrxTaKHg86egsNrWsSKuy1RQBvaxNrbTp0t9NHH7annl7XqlZYXyaSqJuAq7AX
iTfKMgviZMlcv9UMkTOohs/Hll0b+6XSm2NSvS1CPEFylGyHlQELTyNGatLY1b1O
zLl5HcXxLrQRFP57+teyLrPoG1DXhrH+Aq4Oxt6TWiGVYp2Mbyzht7YLlZ69hKo6
VzNISKHdntmtRVEFcMa8FvVAeRUSOz+k1NQFtmy58eaOhtmqfI6gUfL8Sf6NkhIA
f9q+JUVrYSmcMWTfvvFrpM6JNXSc+EXTnEoB5G82iiNlCaZPUEcHUoSXC1Csy8a2
ddGfoBoddyDJ1Onl8hJ9gRkGg0r/89t/DTheoZkfBtEBgawexncI8YoPG4T1DEPX
C9LYS6QGJ7RD5gHA94HRtowI+AR2Nf7TApox1pgtoQVT0DfJJEt2FiwxLZkclYU7
ZnWK+mt6DB7QMNMe9mVBbzZmn1TO981GjvGic9m38OZO3zNOBSQFRp7JQwI/z7Qn
2BZBLHsFsd4zp9/BOj2uTZF3E3RZFqsmdbqTKqdNy1tRNXpPZtCycp3XRSn6b/eO
IqR6gKEiAh3RQPvJYx7kLkrrIs18HCBpLR3mPLrXBYZO/8Z4ioz1knKwCJAEXdTA
z7Udw0xvgPxFNy0N6ViDkaTACyNBU+07nDuASxu+V02XRiXKhPkzRMsmGfVbSjvv
mG+emUJytj9cB1DGYIc0s2e/lkefF516J7hYJx73rMXFGD1+ThdPwziMzNm+lgEK
jX4cFUfVjTQZecZdkEG3b5ns6SlTUDRfVY6vOuDITsK0D8wxA8C4873TyYIOQfFD
QbFjWpkZ3brFXLrj20V9wMCqIrRVMh3F0n0DLnj6Q+3EPQz1+hCTTLP6Np7of2T+
eXUUP6OA9Lg7h0iAr9B/FfFPP3a9/KmPyT0SgJnSDJnkNwi6WgvSYfljp/s8iikd
cqrhz07WPBP7awMoNtsHdWYNRBZ1SfwiVDxwCobM+kZ8KjlH1cgZXKINRiOhBoxf
Izn5OPC5JafFBmlt6SVqvbCB4qEa3P9vumofr55r1V5dOtozzJfHPkwqABJBnm/S
3bcNw4ecN8vzCq3FkJ/X4xrkqFVPXthH3vgE6kDEhMu+UUGuoTDDYG6WH3lqeH86
CkbGyTU6Qdll98W7mt1vUc1xMZr5t7zxfFAS/YJ6hvVd/KNTTTNGvcZC559rbCDW
QCFwBzf23DSQTQtzCHwSyBpGWscSWbzxmkr1GImW+JYv7/0oobXwsJ5GuEMePIXl
zurWHOrNdlrkRxJ4jPNnf+sfF1pefjGCm+G7ImBy8FUHfFrzKodnOEDOifw4Cwnh
PmB48JbX6VZk1bRTfENQzOjimDxPsGdhn3PoHS96EpqQG633TS8IhiGq6atk7h39
BboGFVIBZTgXFnIYuS0CayHR8tk4hECtbLl2gJX4kT8DRvYZhDovWdIFT6s7HuM4
oFG3GKYqVepAYvUD9fPsoNJYLGmjha6OYEWTi181V8EEwHGH0Yk5YjcbNu+xUNgH
+c/RL/BhIHuLRrRKkzjCkVLwbLNCrHj6Q+I0YD+Uh0tho49AVmVUfMWvpMVlOTZm
D7yfWkLEktJNL2pKoz7RXqNKqQj53XycsqSl4yh3vDNNYVuYzK0Ke3uA8waKS3wA
17Q+qD3JD06zBCMsSv4mAirXwsmz2cbvWb/bPBh03Fkt8fKg8QMxkhykoqB4L2RL
1EIuhknNjvmDY5dnwLt6OUatKwGznWN91ep5qoNIsUrd0OCAPosCwNT5bKj81Ei4
0Ea2UDmK5mFIMsJ8lHu/L2zLzkEQF7UHQYdkULWbOIRia/YBcr1D9Z5V+Yfv/h8r
VTtQmsIQH8PxBQyMqyoqBrvSeR4CxNnJYgKfXbLMnJvvB+2Y9Pda5ppywI/vtFHw
Xlj0lCulrkrYOKhCUWiNk/7+7xsKUCR31KiVUB2MDDl6454ekc6fDPd2fpQi1nii
70ATRyeLoBAa6t1mCnlQqGNb/3eNS/w//MGz4px8iOlPw6vmwDXSyNapNgpMJrKs
2eTTmGcHBVV9AKNjoXwlWKnvsWiuqvaPyQUNQRZbEET3oRO0WG/qhLerjK45AF2V
5Um0eM8u834XoB12lzCLaKYo9nRHUkICdnbmbvv6pa6mnyoCaW21h8GgAEz3Q4I2
35Eb5Zx+FMqf5yToIX/6NCtdL5Y9N/nmaW+0YG5FXDinnr7SBy6DpTjJoM7YHCBy
n/qjrAJpjhxTR+XvAB7FSD32+3Qug6omagvSjxGLHbD+lj2cqwloB4GQYu+5Z8Nt
DGbyWAqCqn0UxSN/OXZSWz7IoORtw7C9XoYfY9pjm7mLxvfCUenZs4jec0m9G+YI
T/gWfYRHmkSdinLqFu7uOIfG21qrVID/yvWJzrSOZWAf9dCAOurtAhqXetrwNgRG
+G84mrFd2oppCU9YXkQciZjP4OKEwr7b4n3vA1qFNhzkr0psKN3TFHHO0oMiMo86
fUqzDlHbQ+qp2vqiHUILdTAod9TlUQZlYLxi+9/EOQxG/C+S2t5bedZEoxmBp99g
+Sc4vvgWpu91P8aDiEjAYJL21wC7NS8oKDUls9dKGzla3yfZlI2E+isWuMHnyp/G
1904EqnmMrqK2AsIMonxxkGqKHNFjYZkQoZd7So8wCzudgMlBqjOyrypNFI5h8OS
N3MN73EN3R/h4Vc0kohfkM1vpKyNEz2WDXIkQVqvK38lsxwqvvwL8/Q5Cgb1eDaE
TfzfP9+TRsQpvpORW8lTJV98RbbqbfgFEBHajcT3cNo9hj3VnuehulF1xjY3A2Fi
S3SIHOkEv9j+y5TpC4rn4+7pNSWwZkUSyKBf4jmAGv+kDsNmoXEmREGaik7EJw8t
wy80nsvo4oThgO4U589QBAgSImvwVHiITcwIPuP/FroIj5t0n505P/luHqcs5K9J
B167eC02eOsUFvCcychXD5o65MErFvgHrIh8yWodZZnTEDs4d0gI/Pwl9+nrUYf8
M6JpO0Mo0gOIvPViVoSLua0i07OasTx+tK/cGrOrBpC2IPRq3/lYt+mNJsIqWzFp
RT56JrM+2GqFXDLjKo9f53goBV2BeB+3BFmhFtJk5WN/Oy7mxYa/GJG/zL7RKgcz
yOg797cWrEwAw0H5G8Hx1UK/6PfTr/7BLWig3zNECRoFCEL6Kx13FnzATKvJ/Wsr
qhVSe0to+QcTZIFMEeqJMcXO2hzucvqE/Fp3UZNNftfnI+7wfXARv3luYdFOPCd/
bR2XvewmHMVT8ZXUC1S9UrHElm4S3CjjnMu/5hJXqINbFvKZzP9T3a4JAP4Ls5Xl
ERnu8ASDHoxuGndR8i/557NtLbnhxbNnp81GmykS3PosM35mWXDVbEGeNL114SMW
sEjt4ljV48bupU2d8m+7P2FSGIV1EygLlk7insLD9hKCyO97/tc4JP1Qms1BN5pa
6v7ta33ppjLHTPq1sxZqIjNIUYcQ4DIZazS2h5mcMJn8PEEnJzn8qz+CKDfRiW5e
tY75i1yyEJPRykzpg0UT1l80+t2skzcPhHl2VupjdOwvuUInwNEzy5Q3V4CHUDQu
U5sXmCxadj9Ap36j601lZOLGNrPiFryZhYDtQTdr9Cn6SHu7CKlpgvrjE3GR24LT
qWZRTO3Iw+BYRkpKPdFbID5TNObabbXJsx9yZKnyAFp1WL4REV0hcUFJjcVQJbk4
IM0pxGvhS2x0L6QFHfy0Xi3PgQ5NHtofO8cI54IAle7TSV+9fOR8uUXtd23Sw/uc
xfeAlzIgTU0jJw9e8YN/HIlLx/7fmX1TKstc3iiSgsHyNyPMEX4Z6sfz7fpP/Dqa
H+qEmJ1BBnKARdGFgjJq8xYH/Tsldy6Uq8w0NSvxr5WSqEEGXgEbKglnyXkLDkXk
rKcHzpITEubiTF+IXXfFn5y2ORqB3N5BclJwHVAQkqcwsVMwM5XCI98lHfzilE4v
m6VqyNzTCukEH4OGENTsFgbLRx8N7R/GXQhT6H65NflyZfGfk/29afOboUPzS/q1
3AXnEyviWkwMkqEjtUYl4zUcDBsU+D/0rzXQeq5kysQynQe5GaT17RoWGCBnDdqv
AfcHnrc8oTOp0i55U25TGQ7y4pnNQI9ZFH2bluKawNAMHETTI/E6bW9cPmtjnpvV
YT0Syk9F3uv0sz6KyRpbaHO+vqA4p2j/9rxp/vsBDevGWsqPP7LzE6xxkEGSRfVC
nfG2TrErgMKVwksT+2OJeZ910ElbI5iwVRCqN9Xhw43RevuPRqkwqjQRNEx+ZU1X
Z6xUvO3JbiQnp5FkJv6ujq6nfCrJ1qK223pro9VirzgIUj1Xpr0U3BsDQsUWoVG0
rM8+nr8Y+XeZ/NFGk0+/+US6IBZtvxLVzmB6odgGLa9gD+GM6wXNUu/MPDnIuh3P
O4lEojUdrjnlucjyPqmqlv1E0G3vUHbnjWClflCneVdMF5UN8psvIiQHqnZcAAtH
4xEDhs9nwliCNRw3+riJorrYBcTx/CL9n6l6nc5HFK/evH5CJHr684pFQ/qlfTLQ
fMhF/neeza90mAz6QwsnFXuM/fV/NAKXeBCYExpr3IPFUJ6JObJ1B7s3ADMLgzJf
RNrJHRczlvYY+1intdw2Qkl+8Ju9p2YctlKbuXoxSeqs3Qg/yXxoB5qMHIMx2TUb
8bKeWFwgYx/0g7Vc2OcYP6qu0a7MZLAPeFmbUv6iDgw6yoh0S5uSOuDzzDr4Vjim
bQTTnQDzrIxe7G05AdvPMvCrHk8b8Bt0G3hLFyxKCUlGPU1gs4Sy68fQO6q8L1hk
Sje4vXVbIxhavUaOO4gK72drf7xcpCJnR6uzLoTexe8UibZzkAagsSYKT+nSenEQ
D3cEF9rEyp5rX8SNNG36mExgE5/0AqkkRVcuHzJKe5q7xwSYF5qU5TmqpuNqTnEX
H2/W+L5INOMqGk1ju0BtIjySnK+4bpmqyq7kKFWRoh6VSMusJA8IX7U5hH9mNl7O
K8AAV4omzFZrD+Tyo8iIf2nGqTJbo6w+sAA8QO6feeUA6AXi1ADzyOYxLCj8Il6q
cFiA630+j7fssG/rQsECPxRYVuktBJhUQVkTutxgWKaSN/xUgJk9/Amj0ZXCveuN
BjVaiI4IHu+rMtCoSVyu/m0V8guQZnF+8v5WgbYo2prHtpK+bStq7n/dMtn+wmou
h688jPvCRtfd+3beHC/HuZyZ4sPbPJ5uV5D+/um+39yS2EXzQkvhZBtGymn1wKas
fd59IZ7MSBIr4IDGqbCXZcUN7HsZbHzN0RrzjGVeaVdrKzjnbjEy2LfhVd6qruSy
F7ijJSxKh6mqu2SeFgIRcIU1YjwRQIrMgKz8gRWjUwjdML0pDuV1A5NJ/8fOfADv
4vakOy7pvtmwguYZuD1LmDA2eh3hKbyPtKH3pwwEjtqzpAxfY2NbKu3ErK04A6lN
+HVigQ5Q7IKo+wzRkQCucach3h1oHQtU91qEA/QJHmVfQm4yk+qqWbWaU809DlFi
BlK0r88wxvBbw04ee5BRGUPABCUQlIAdFe94YKMr8j2VxUAP+uXrCg9DcD1anKGn
DezEKnHb/pVCT4NRZszwUw==
`protect END_PROTECTED
