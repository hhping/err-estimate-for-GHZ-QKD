`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6otXCNLriHqf6OAyKQUf+vKk0y5Hpoh31phaIB2j5K0effoUSFJqzvgSyIf0AnR6
hA/fKHAVS/yJiqGZb0PA2iJH1JZQpvwWEs2YZOtMgxng4kRbVBPUXVcW635+Atti
DtpB8t+gFI4flbstyvoBJCA0ozE1axS5DvegjR7uPlXA0T+ikCClNJDrX3gNJiCz
CG0llko6YkOfRiptPDF1GymudrWYHla8llUYOaiFkc29/WweX8GVY72+xS7R+ehP
4RRg0gVFuUlOZUR368xk0TxDRb+77/2J0RWp9YDi8UOKV5QBmRpiO7/6WSpqUBow
1BlL8n1YIdr6NbqPWdsoiPNOFEC/sbNSHlOHkPivszBfPPpP2p9CIycPEv219CyT
KMoPYUqaB74UKCzuuuVLOPFBnrOwf6uuZnUj6IVE8SxUzXm5zmRyo9z8FQTulu7H
tnQxcaoEem2bZaiFsckzJEwm51tpTmajYjAkciTVVtFu6WXBFGDF901EILrgBIwn
PhScvAT/6U//J3loDZXGgcMIcmEL0y4uTypLmWni801DdB5M6Fyd2epD4QGqOH4J
4oAiqvyxiRHC4WWpz4Dr0SFiy11P2VrIznCFxFebrLCwcFRGwBA+nBoh/8ymSwto
1OFIGjG5N3IKNdUxRSQHddWuGLcxp+b1VLVLKrtZIOQ+gjzxkPYJBxeZLc5VoJkT
N5jPEnSnXD0Y9wbHI3MVVFn+iVa3a6jlbUGwhcy4du1Xry+SFvHsASJIojAPn7Zz
ed4H3+3qQCmkkvqO8/uXsFisIK8iujkRuS4ydmJFfb8UGQySkzkmVEjXWzLjV/Fe
h0Dl9KOa36stMsQHbPLetQ==
`protect END_PROTECTED
