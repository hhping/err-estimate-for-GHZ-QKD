`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cPL+xJ/Y7VNdrvpzpmr2s1ToqAnr8MgspDv4o3YS5oPGzMunI21qLs1X58j+QmR
SnlXPt+aiwV5YkvXWDjH7VjTNod5AWid2tLhBLw9cPuvxXaj6cUUaP6ASWNrvMUG
FNoOvTGl47tuvJmiCml94y2Gvt1vfnKY8eFVKY42GApv61ZbnYlVL9HlHJbTnJDM
fcXENiDVWqjx7ji5HEc00p7QvIcmpDY5S3QbjEzXR9jWoBUVZG9PeTPXK7trGQLV
xko5Pl8mEKQsbFAPVnmSF6zWbhfQ5Zch1gmCdIHzWsnjnB8cPH38XlYDormMPyt+
m6YSYxlTonPAPLrc1RvwWtwZvcfxh9Lbfh1QIWyYe/1H1JOYYviUh2NtVfbQmM4m
WqOQX4BMWkTif+IeA/S32+qIMMoJoC1mYBD2Li+79qp51Hapfn0p5bxNb10K2oqL
J38o22nhn9EEUqJgqpsx+FUN6BLF60jTVL+lZd27wBSZmq9UwWSKg0lzO45maJ5Z
Gccsrfra5Y3n+k16JmtRlWup5APgyNhgUDMI+xrDDFDXpbPYaNVZDMQu7D5I+gX9
lyOFDSLveVcChsxZjQlNHXc60lem+uPWbS69A1XcqhhRjFaj4ym2UqLSvbf6YVtf
5mK/OmkArD3Duwad4WtkgznqtuLAWcGu3Mx7rhJpOQphvjLC82x9laioWKIzlKN2
X5q1kE/vy7BhztVvjjsD46frlE7XKWkxHTMZ54faG3peS60pPI89o/tp7kMIe8Q3
82z5DXHm/klaUyvQlVI3CxgXm5bSlpPUWdR+pBpbLrDCX/49tsQCXKeBbOc6qwfT
HvrX/kkGAh/zGiD8UlxI4TzkBLNG+5N+gx38OBLxui10XH8mKNE8rDk/vcVH988Q
b2x9AmAZgKPSfxJ2RubTsXnNyR5pdPKNSCV/M/noiHWArdw9Aji5vyogehYalKOr
4P6CS1TtX9Nxc5b8E5eRADfAMrq9p/z+VHm9u8yeaQo5VSEZ/uIgh7KN0xdHR06w
ZfzCS0XTF8kiuPfgS2MmNvblDsDQbDpUBxu/i4Qgldlnc4Ep/i4/m3qYayYw3PqU
vBOibBY/aEmqHGIqk/BVY15fgct9Ntb1QdlrWFBJzQ67QMAuCm2E5sxKhtlJRO9R
UtIiPmsy5old0mL4JHoU33ghCmjQBaTK/M7IT8ibGK0/mWMXK5rTAUepb73r7cLT
3HkIWriuO0X4QcrlRE+9EA==
`protect END_PROTECTED
