`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yorRqk/FNzUB+5w3H1FZWcTx3EMQ6+SZL0ZJs8L0rWNwvXsZqc7pn7rI8sVsKkGs
UAYvokQ5h1plPsHuLIJgyuL9PoriWh3E5+TIXoPwzWgwgwC8SVcHGQ+0CvveDNex
J/CV8WrA6tmtGRtQYHCSkSHWwFuWGPtMz2KqV5vP2xK92aYaGT1meqXXNAwzGUmu
u0f7sRAFLW1FISUAOLfhNXeuOYq/7ABKckRWgTz8/IXqlOIZAkqYrwX+AQQqCA3Q
3TdsBwMlI5VNjnfJiBnlaZFvbft2oa6sLkvelXBxb1FBf1HRv41CeZ2i/XThRKQo
v7kdRfMVFlJtxHz2H2aMVnmh4dAUwc0CCRmHPjPynYudbbrfi3aF2ZAA/FeG/734
tltNgj/6CnYH5l+5n1y2jwfV/XzwCFuq6vYHYb+8rAH2tFGdzxS48/Ne0V+/4Rzt
7qZdCuio8oKRUW9pdrEj7b87NNqtWt+0K5LENpElMSnfVrLiUFgXeR4bsHvpUq8t
4eHfQx23HmQB6yvaqeCR0rMoZVUkDuKRWIWp1bAU/bY/cSuskt+/gEGX1M9IC9Ux
`protect END_PROTECTED
