`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lBSECVkV0ZkvurN6Tf0jNhNGIvLYmcqV9GJS78Ajo/kE1yF4wTj1CUjimRLEGuwh
Lu9Ee08uKN9OcGbxELMGegtUoM3WhSyhjoMBy1N271J5CBrUU/LpGXyG7D0qJTqW
2la+P3jz4S12tLwGIu9GBMUoYXZg1KUC90WsBshUcTCDOC377jKQmIrbAMt3yO4n
fgZFJbiiokInlOjGlaDDhDx+962V0zCjfoXPOPliQXG5rHyO3O+4ptJu7bXOYbp7
WXU63MvAr/0RcjZ7qwHbIYtTZSj8pC3T3MBfK/BDGIbT1/zrA8OrpE5PhZ/Olica
qa2Rb0VTjEnFmcJ1eMmlWymne5hJQokivhy61Pvp7RQW+i6VWlmdYxxsllInU6Ke
jb6zY8gGyv17x9eEaHGUMxk/BtQrgGSBnHHPgygUvcI9yhKRnTGGrTTqmjbbp1zg
iMsAchgpjrpvSfAK72X2Ncy0sOwjpPg3QNiEowzk7/8p3Ku1AzN1INlcmwjICc+n
XsizPukfSDGEf7SbX0uMs3o9ZvnLyLo05FqlaG+B6ec0RfqOQ2sLynB96Cd0XKzc
ocmlWJC4yENeu5J5W0ggWQCc6FwkpeWA3TctIChFJl04KVbPLiBewuGzJDD5I3W8
LhpBRiHfjaJUyKNPuUntTwu32fIFy36qLTADOQEPD4b1yu7qDoJJMRhhfml77QJn
qYzLWcNBrLNq+89vJN/U9ET12GFSNoCGSh8dFf7tPeQkN83gOLPF07eUGgplrHIG
wpXFKQIz/eZimbfyu8uSAVRSoDXVoeMMttM+ccWL3yBSrrtJ9vc5TBLH4XMB3HAD
4ZyXw9YdRrl1nHI6trvSfkV0NaSUHg2mMhlNXQtT9hdAasD1Xfg0qfMIfOD4YlGk
JiKZVFT+aGfAECbYAIkGRocSEit7PyWL2SK7ahteewUYvrlMTreTrn9x1GF046Jy
RGyhJYMuvRq0McP9nUETVyJcn3dIMYPOVnrLwhTkqz2TIwiUVxnAJ9dWK4ALj62g
jdtoRO+hrtvgCyyPLDy+6FPfN9NcoQFHV9h6ExM9WJT9KnTMjg/PAILDJBxn192S
GE9fH6e1G4t9g8/AAJiQKbgZvgFyiXKV+VVDmC8MblAg8MDtoHRHnKjoeyMQxDjQ
F52/cK9mj4hdHxduLfdCpcD+hfao7g55MA4+Cqxw3wodXNsiEJNKn7y+6xAOy3Gj
eUOIqnqH1m93Js1xGts9x1rR+XjCNR3dHfnJDmJ811SWfOR+C7RXsOzqE7rDiu2y
zk/+MwKCn3317YEcQUzM/fstQxSlPjKiahDPhfIB1gY1Zd4YG9/q5XCcqpr9PkfS
OPq7vNb8fpawPkDbFQ986awiP+ED3YlyhpAj10vwtJCSVkDpeScz0fB4B4vBqK97
bVPDJJ1e1APh0MhgnaXZb6tGkDZV6Ssy9u5GUII/g4qF0W60IAxns5gOP2NPOck/
sZ06PZDS5kh861yjuT4RNY3SNNUoACGJA8QOL/tC+tHS5QqgxqtarYAC6WMtHb/j
2Kcr6B38tMhpb8ezC7nDo50kh+nbRGlOs5TFXNNrl2W4ty3maN1np1+PBTQDXRln
nBkku9lGIXDsuQ252VwrF/QQbfqs1T/44ftDDVsz/HB4W3xwk1xq4eVUia2TH8X3
Xh5C2+pHgvi3eBMxjSnybIPCL7dgDFKmbkcD0liBmvZO88KZ494SfF/teNzmajqu
XJCO/rEkYMKxNpfGjnnyIAoxYXpeD2vD9vf5n+XOdlfWClpVcHVLoFSWA76DwSuc
AhPYrxsqFhhwfjd/EjFHKctUjjuTASxa9C+MsjL6tw8vmVPFkQ4onQD2+3JfGivl
b6DcEiVzbkitzjImfVE46yOkX9AlkMdkN8vrzHScswb8cHFko38Dui8fjtrbGmGz
VWESM2NWmSvZRU010soZAWNmTboBdb3+8LLUTrlXqkta6BNKQ1O5xIsdBMzdM/Km
DekHAUn+pPlcKexbHFZKgozCFqvaoJcq7z14nOXImYy3cxDY9Y67ox+nBWHmB0YE
yiWjtdtk3Uq8Ghd9J88wN9xnrbtN5QRLPPnWa/FxVeyCSTUbkVijvHt87bdyPOT+
wMxpJCDT5wunMmJ+LD39ZxX074JGDBrxmRzBBbUNZvp6k6O3bDcwDugSFGRUSAHl
rQXdYoKaPBOO9GKUDi0a/VL5zbU+Lgf37uR0uNbW19SlaH2wxa2N/qyE89t493M1
DOAvcRtt849Gtv/L/fwfpCFv9C/USQzb3+AHl/wyPMWoJSIEhHF4XS8tBFFfSTLO
uM2uhaSdmQSfwXGxR7tKzmy4fCg95wSt1Y0Bx5aeiIExsTD+FrqfIpXnc9lGESk3
kiZnP5abURRuM4TFcpJyrCs+e+PphjZnVcLU04Ybq7pcihClEB+KRR2j2xywvG+B
mHHt1lL/bCGhoaQiI8MQ+soUFi/Npib8yXD2zibO9YVVO25lke0jftQb6OSOw+So
YH/GDjEr3r4rQjkxHT7d7l0EPuPFCV/9fvui/MgrUMnWf+H8kPqk4AUduk/wfYxq
VUpXg3vBhHmUhSPGubgDmptgwaGHPOIAc7dDJ2aAiY3jqY9lzbIMKNKPpO0nO4DU
3lqyf6Ysv9jZ5qVLJiXRYUJmdqaTyJneApJ8341QPj76DdyDDkc12toWXT0Yv3DQ
72VCGGjr9lG+Q3/N1OX5NQVys64KkV7FD2Y1l+MEVEpL9+PXrhB4ON5AfPyQgBB1
G2+nlKL+fET1rAQjzusBZniQq46opm4fupQn9RNBMcgfHWUAcFLo+gxEvrXD4yVl
lG0N/ImBJ7I6YhA6quoqoME9oxPL4GLvReGmwZVzaXdqZcvUh83GYVUXw6+OASP8
X36F+4ZUvbyO0aePYRFYoplGhmpla2WKLN7fWz+HfzZwN5ol/CYTfgE0J/AbFJ16
Doj/i/qSH13cDI8lJtu9kd4jN3WqVjy1J2mp0SLEQCG7MrwaqwRzJRT9hSGxt2ud
WqGUVKq7gcW60F98JGrwpPqni1B0nnyPzJoyrsYie31ISwrqSOwdvuY0fEg9dRK0
pokotD/nafWslWbvgRAoFO0CJsj2+zO7VhbsAJLknFno072GstvCWkvTymE6LlM0
Lg8V+Gypd+uZak//gANa2Q7bPl5AnwOFEpjjexu/53tmUgTzgJIrdZNHMjf0jAme
JxkNndvrPE8GuwdPQr6E0FdDyUA2Dz1AUVp9iCpZSr6gvADwc/yJZWXgoCkwD6x2
qysEq3eNcThAEbHeMGBiG44dLWpv/0zolClsDr2oH4UA8m2n/bx2droLzWcU9CQu
IG9Ox5I77zA8sTMKhLOj4s/rUeX9VKpoArKpcnfzoKRd/GgcFmC4XSEuGXBwKJEt
pRlwbQqVfERRjWJsbIOTahLan2fv2ffwW3SReJlHNk8V2RK6RU6wLFaXfwYtvtnC
BXqPFXjtiGO1fEShEuRJPOZAEXPhYIDd22SLaqkvrekV1GhgpvOe65SeuspB5O9u
VmCzcwiaH23SxrKgu3v8OZuyDZnYKYV32Ay9+wzWeFGkgar4/lqRZP7nHOxcREeJ
gFR5kNWsyC8kh72Z2lnpsFztonzahfanWlUlREsXlBD9N1TkhTAZfRAnO4gJTqan
0m3fc8eS5uX14RZq6QIl7AzT0UFrV1liKeq3g15myPHAr4d2ymHVRQgZV5mDET0Y
lfhYxdEZj2+93Ns6mUShti6q8tge59VFFs0ata9iW/fUkVIxrxc9s7sypp7MmkuG
IbRqXL5K/wG12c6x2oj3rWYc4/i4sCX6NCBVzP/y8In3mhiK3mOpz0oQ77LnZhbX
XfIbp8trVNq5brOjzjZXooi4SYDZiyYSwULGlJtZDZMN/zHFBpZN8pDzkK0m1sFs
SiTlbrHqqSqS7lCMH4dKywk166XVWvzWWCYvmey9H3oSLacfzeWsuqerDtnvAmFm
jgC2M3MFeDphF+/AbSsFgbPKLXYVaTDn0YUSvdV/Cv+TFZdAeTrqJxNO1gOd+dk7
X7NIg7LGWKP9YLVUI5yvWBDXvi2V+bMBMtZS8jfmr4ILN3PurArL31XDaoPMM/3s
xQf1QjjYEK3UszuWtGICaMOdTFAjC7rpWxJNYKV/TUs/wV6WoMxREhLXUdx2ZTKd
VI1GYxuLk10gsdavSVQOp//ShH/Ey0yhSyU4zas0ZGUpUAKuOLQlpeio27XxwMH4
MjUUHXiK8Vs4Y1pkGvEzPw5mwzeCQrIjTJlYiqYEoeFMQOd72CbGfldWmBS9kROn
zGV4WuCpMHGqxky77NyjeVM8/6UxljLY3YtRduvOPzCUhLqDDuQPFTJzBKzyhsNH
3X1VFTVYK5zYNmv5uFJa+qP9w5Uggj/G9v8c1FJD3Aha4gT7jkTBUvEf8qddlPeo
lb378t488AKM6mThGFRRS0ohCa3z/zYfHgNWLaYsZdSB1H4P1yJQn+h57Qg5bPE6
b7lqG80bZ4Hp0hvr1oaQ+1AIspDETgJjUGDVmAr4z4X/vm5l6V8dVkIMWQNNAib9
jl7mpMcEx5ALUTaQVhAEHRope+evy3H3daLof51erG+LWECpln5RyXH1vgM8OBSf
rbhn+5/VomOlt1pnbGohWLPcalNTorJaWJUpOhPsl/hx2uI68i9QuQkceXkAg3ql
UG/M9Ygo1TynBVqSrP4ZfY4IrL0r4sV6byNyB/QkNpOonE/u532n40uu+Qyliq9r
NuL9oz92KlN3f11DZ4A07rQmwn5O5TtEehRoWRSjOvSinMiBsph+Ytd6wBIyQKvG
phQh3SGORfB9B7EHwDPFE59c/DKh/eNnDiVnYsa2IiussPjuBnthHGWxowlEfCdO
8rWy+gGGsrNMIzFWPSTSoJ+77GJewUN/PtbtjdKb/94yIc1wK5oYEoCk9e3lwha5
J0QrzcqlA3OtuYaK10CrlU52wdfrl9yYYqJuqr7Egwr8W2z/pKC7Tdmr1he45/md
nu+jEma1aOPBdTVsk8Ez07djBgzRwG4WfGnoT1YIeoFVnKS4Mqh8Df6g33FIm/a4
gzrJ8Pp2PsGZWlVURZ1Lt/+G172vPZzxUW0e9TmGj0YdRNjAdy3ddcDmwEXcrjn5
hYfjpE7s4tx5if3/cGWWqyWHdUH7cTPT6m57itawEks8JOD9bSFitBnWUm/esP3q
NxV2SU243bcZSDXoRGq92X7j5sgcSepe4kxdPNQjRAo/OhS7PCsXJ+yM8n2vzT0Q
mV9KO1spNkTBsmh00g2ezb51SMFFMKQL70Dq8ocxGVHs1gp+t/BmVC0cb//PtaeP
xhyZBzHUhahbvVx9jAXhPwq+7HOTgAvmz9dDMezf+3Yhh+B4HAdMCOHZ5dfNOd+p
aDfD3l8E+T2o5AbmKYwJDBRvbommmLMUyVYLrrBcFpmr4Hg8xig0JQWcASDh97M2
iDKSOLR06OcH7qNlrItSwjoNfWkRSFRK90XCdWr0rYBiPquUc4fjjNq0LqvINnA9
HIicBuz90NSM+kXs9pCQ5oFq6qe/F8a1qbFo5c6xe6GxZE2vQAyjEaINwZ7VpE40
X2jxw6mAjbSFHwwxCp/NEPZeOej7M+yoXCiRYIXMd+8ykOVfDjsFQ8yHYbs8ER7g
dfhEx7eq/xfEIzpeqKVbgKHkQLiA9X2zLUkJ3pPlnrKcrMa/rGqkFRLW27WCAiAU
FM4bKeAMxw5YBppye9gUdnPv4yFdkxCOdjw+ddFLijDscdnX9lTJUAuALuAVjFCm
ksg3+CgBx3V26ZJvwIPEzJeeixQE6l/U8gtuYKlmY/3tuX0Loc5t1SFTK9m8KxYN
OP+VC3tXyB/tkO62kgtg7p15J0RWHiY6EnbJxDtUC7X4eFt7Ep+I/euS+4Scft1C
klbegiFpJ+9xjow3MGZb47pKf+GfUf/rCAVhctusrIgAUaO2xT3KPLRsao7jtvBl
FlOyuMzQzpVuWOwEDnh5XKfD44r5SXfDVqIoCJzCd/iA5jDp4VbwdHYs2SmIZyvP
B0N5mBNyzWUt1QZzMZAtOFbwLzXYEmLx070ZUxNdwRlZJr5jilPzCDrZ75T9jU+k
FWzfm0Vi31zM4xq1aVneDm95CkXsJsdWnOZn+XQmoSBbjrfAKy1Gs/YI1nkKe6WE
01kp/ixlCqNt28tEG+Z7mlLdF4S/xtPJrqtza7YvtUw8U6zLzVWrBpuYX3iHu0S8
8SODyZaxU6do7LYnIXPd4YWy6cQxt9Zfg0+IWHBIRTWtFfMTyNqrWHHnXAQCiE7B
B/TI454LYJtHeWBUpIeuJoDEij+T/jY8XHZlXuA7tm6IXxoKAVZEn0nlgVM7jw0I
CgthWUNasvamaQJcmKnl4et/tkn980BeQ9gu2I45mYjLrAQVDDBvv5AzcbWRVAsv
ZfGULK8N2KmTssKalz5ufhxyMWARJlZusHJ2K3zB/DeOCUHLqamb50WegBWrd5er
z0P4jIzg/7wcTTRU9VDj33XjW8kKQIqi43aWTTSYYlW6vRAAwkJr1hgBCzSyi7fm
ZSno3e82YyyY3XaNPmpg1zGGen15aQ4eIe30FkPfkn1UGXaaWiIGqWpqZ0/O6mlq
4Co7PvOWHjh2m7CH4u9X6h0p3FEKDbEFq8M28WgtTKLspQheTMEG4EHAf9uhTHUE
qozoR0PL4XD05DjwfP3Z340Nm3IFBTngKkvaYk2Tt5vgTMazjO318RA0RiTc9tqe
dr7POFEvuRdhz5/yf0u/prY+Gn3PdGL4sk6OvvJuKju9NvSM2iZxvqpp60tHpP0M
e+mjMXrAEW+SB9V21Q45GR5bKOp9MGzkGBJmfTQJSPe6P89C/r5ngg5FR1HtIa1C
1R7qsICqtPZjREdKo53uEcaruGFnFh2Vg5bfg9dy5dSLiIptigxmJwcPZzZRS5s3
HhK0T16IKucu0FH6RPgSRce3KpRv+9WsZXlQsoJyyAe3OugP3uuEqWzcGrv0Oa/Z
zn3xgF/hx4WB5hYHciOi5pSTnBtGrJX/mitsp+7TPdf2WWTMwC7HOpc8+n08N3bU
LWB4OupIfK/eqhoLW6KUJfP47Ur70xN8x8qCdRvGpdlL9HRAcWEMYx14ekAtoveP
rCFTm/qv9JchhqZaSjUtvOigJhCYuq7G3fyU6KleB203H7KB5i2RFLgooQ2Rg8tq
BEU+QKwjKc1sjnGArfx4ixy6FIIesfb/xfknQS4XxuUUKM147SQMpkTE/m6iPBM9
wC+2N0M1BL3OL0PEBYM05v44aoTsNc5RQWf4h5W+oQRq+Nvg+8f3ZP8bZMslHUua
qrpHvxKg3NEsF/F6WAtlbzxQ/Xw4VV6orppRK4yje9mdGZTK9Zse+Ukg0Qf6ykg+
KaaL7srIj+xtTDLujNh/kvcpXGuEb1C2V+6M+9JSAporzsEf+nkLUTvjDuq8iEFi
eCRq8j3mkmnhExLkrpSOifpehX361B2eY+Z+SepcVMyft0+D3d2t+1LBKl/GkxQ8
GKLCjzdJP3RcaFqjqIVcq5Gf5BoiffOA2ecVqEB7vZQfacxOPcm38gF7QMGIFXWy
OAP3LcqGx9D0FMAGPASL/Jd7wP9INKLHLyHWt6L/9t1ob2XXzssM3KEnp1P0jKf+
W8mG+J8Hm6gQAH/c+cK29b7F1PeI/lFPRw7YeJqqfoF8X8rmKIkTuqzyn6qBWSzp
rXrvInycvjQHVZLh62cEIUKmNgxt3CxId9Cy+jnWMEeBkbcC6Lb32hriwY+rNfv2
S+rtsGzc+29E2Bm4p7KnXwQbF2HqnAA6/TOoHNyVWE0hs7bta4KiWUCIUjnXF2A/
0wPXi0clpgtrZSbWOZd6IXiVYPWkBvyUfPutXxw0tzHDYYZJsS/WvCEdN2T+VJ5R
mdigueezPYuujS7AXtqXb5SHtP2S1s/olwkfe25cQG09kczDTGSJSygbhdiRi6bD
QAMYHiF3Oj+4ObQHW8sVFzJGBVv+Vw5Vzu3ciTRJnsUmMQwGUcTGOMzVb9ekx2/L
dKN4t/WzCeminOFEfIc2K6NdR/0DAVQsC8FeAt0KYcJZI45sg75+MuzIn9rBTSl3
ZzQFIreSA1kaMo4w92h4Qm4b2Tf6uIdKNLeEpHlQY/Uabynug7ja5dAbyAtH52cb
zpPMa2rTYgDU7TZteeLf6VleX66KTQNEVjNyFIc9vPONbWSNuu/WITtDpqD6NyL2
MW0Jw6azEOlrAR2j2YV/Dz6bj8n9H7Sv10vLvg7EtVxcbWMTsj6euMjnzbw1PQIH
axv9nsFUhy10Pdai/9K6eu0niqCwzH2/2N+7e/3JYWwzg3LNwlQF3RJQXC/kMxDi
TpjYaFn41FLlQ58864ao4qidSUsr2UqJt19Wwzc/RAj9uq8OpcSGbMCvUNIL/2zg
iI2py0Yn9DBmuxUErZ8reX1uhivDXy0WG0UBkiYqetUWTfY2+muQe/s21z5lOxFC
vL51byH1tvhfFPWeEwjaYQDiU1B4sYWZMaJhJCgktzu1q+PP9dq/f/+qVYQbeOv1
FuO1pkbRG94W737C15TiQCyX5VO2cDx+YnBaEXUcMnHSWxtbb2bIhUDm7fKfYRrm
zeFqfi6D7/7y2iD201Xk6TbVmKq5q+e38hgbPcrWI/9gHjdVkTrvfjhXB8EWCMVT
KhdF3qdkTK95bOWBsChN/n0vlKt/YVE0PJYlKeOX0OIk1rB1RgHU5cPX2ZOJyhoq
mDpvGiONxtYRAJNPhxhyNrTXvdK/mLq0NL7L0+qRSV9FRwLM1kOIhDV38qTbnSaa
tTgIdZa73MM7BbMF0pwKOwRn+WIS9NchurvglAIYy/TpYokTgZFkzvW2eMGOn8TD
wan0ZimmZnSRlbtVXnzLcLroa94emZsEj2rUYfwm3K9Mk7Sb5cS6FfDw9+T7iqji
95KK2ns7wDKohzu0zAUQG6mbPYri4ubGNuzH572weedyOHv4RnD0uOwYSD7zVO00
c8eGNj9FgiDxwz627L8BKu1TTALSho5pkQDoEOSVX1FBj0c2gefJWa9KiMRl1pSO
bzpzfwi2k1kBlRhMDWer1VfxWP4Cra/2Zj9wlNHd8ZPnMcid4Kx9hGLg5gIfrEbA
2vneZixJJYpYLDJRULfADCh4wkqPEG9jTDL3iQ0mxV9vYGoge/EqPX8B/VWGAK7/
j8gJZTIQdquKhVb2FYuSeH/tKvYHg7Fzq4fApuc+lJZTM1RjJHTLfkLgspBvbtvs
yqlUK967L4ILwvuWihd1FjH6sn+9FG/dVgknCafbnkNCfAVVCSjnoKAtUFlwF2mI
pPZ9AZGVBpmjmNM/9+5nC2axXSBIneX8wK16T8IZF0RZQdbaLKyZsqlN0QVlBNsq
nTXhEVixM2y1+wMzeP2iScQyLtQAY/1rEnM46HIuIuh2AE06ATSf/fONcgybiC+x
GsZMqu/BkG5i019/KS87MpWDkrLlGvfrfIf4enD8/QZOzSrhfRnwAykE7r2IKG0X
P6v4+r8wgahYnhkTTJD0A3/qRrUiS2/Blmjkxp7tRd7adLJO68LPGJvk0er3nGXS
bgZWXDUK0Ia0aknuDL2mjloTRKa/bUd5odSbSbiJ/l9GdwDnvzmWNrLyYFHoYiSD
Q7b9VKxruf8WLwGdT1k0LqQGR+mfoYpgHF1zcG0ydsruGI2NQCtjxfhENl3lMTRi
qA/6m2U6OJcmDK9qGvh/e0j5I3cH8gBjOJI0HJZVwntOo5dd7Cb//rFtMclVeVMc
b4gANkcX9zuctQLHQtouVOnFGkClq1mQOe1Fsou6YQLWXgXHzg2aq/pi4068op92
y0rx903YsrlVwgs/VDrif+WkDVqRwVKkacZzIY/FKAmttVI4buG3EJ6G5UvQb+sm
Yg5fN6mB7UwTeHZnWD1fUcpxG5MY9Xq0S1qD67M6wmPbYqQZtwU0hhpBv1IvuSRN
gkWT8UkeS963PzofC0CnkvOGQClRihWlaXmLfeoApawKtCOEStwqcIKoI71RQBjG
sPa0IzBJSE3QbWu8ovERZNAEjLk6f+As5vWGoPoDX4EXGuNgwY03AbQxv1ujKKsA
juFHrfXt/hR4tJVbSIIZTzWOjEDZLEpAYoj2v/U78oLnR1u8LdOM/Q2otMTvrmCS
thjHqKMAmhI8z8jo3du0cx/4V+8iCPYgX+ZaNqlI7m2Pr3vvv8WG9Vdd1eQ5jPDM
SYtroX6XuRulwU5G7AfyfcqFJmu3Y4CM4lnQyQKG5+mLM8vP0pzf2hFY2pohj9na
v+fPavDay7Z8w7XRWr8R4xFS1SIOHEIvLwN4MxdIV+kQ+YkTQ2sg2que0Sx3Zm8E
cBNn4AMydt3/aJ/HKdAyrQx81rSRf2WjXMVwxCOkfdAJU1oJTxP8hnqSTARvEett
e3PXViWZDRPkdjr9wdh95uorPozOfTUgdoHleYIJNjcJvZdntyaoFRK3yZULdV2J
QSQ2FFZ8NT18cJ1Wo1onYjwq66dWO3jInh73CF22SBGfZ4Exe61QHt8F3VKmhvyc
aQbvPb+CMJDeT581uiI8detwfjrOyhN4fG7PDIvQOFZWhUQkge3Nw3GAvrpReEZJ
k9w/S6gqncNiQA4D4UaHU/ZPlFkBJib1pcWuSiLg2hJCVTqTp7a86kt1y6oGb8jz
VXSkay9fxGAvHvRj2PKPoj+c05Kb28vhkCsrNx934RkErJs8wbx9d45LutNeL27I
C7HXH7CB5U4LIACv6mGbaNF5MPags9Tl6r3So2CXZ0KhiOPlzxd9FXpHIcE3T08T
8rsH4DcLdymMrhmHi+TD3KHoPQQas/7X1tn6O9dwmF1avXLVN9zePs4gwAHx2HTA
qGPdyK/eNCzWBgfXisxvAYU1QHoz7xLFTBVH/eE7sK90gPlAqZEyuN9QQItOeUkV
eeh367Ax0Xs4Hks6mIWIk7V9tuli6WoMoOivjQ2PCLDZ1TmNxA6tnYUf50W+5/KI
yV17X/Sz2q3k1r1KM1AmCv1Js6Y/1lYBRmJK7hSjaXjCXgjn2jq9hi+iBk/8HhEW
XTQvoZWGBQJLuMsjfLCeTpfs2Hbdmjqxyd8A6xB78v5KOm091Owcv/vVaAEmACQh
TLMHXIckaNoaCfVGT3/czC8aKcLQK4fhXNO2/ceXgjnktmWLEPNJk4+Pe/gAp0xX
NyJ4qV6+avRPRVwLZc6kIFK8ujBh1nd2x1+96ckjqa53BcdV8NG/Za8klzYnZCLQ
Fc5DfZEqMKxrga371FPVsBRQw7ZVydD2MHnUGra+0tWtl/93BgPHCZZXHBg9/rQe
YKhZahGYiGJJ7SUHjTkat6L2LWHcsbYS/jTdCI5uMufDpqTApyYigONzByV+r143
HPxD5JGkgKLFYXbx7vFvh5Nbda6ZM5Y8hibS7NSczNMBD9zMSFaEZaNsjE0d2zOi
oUuwVkq/XVKqwl+h30Jt25EMi0XHtG9pgSb84SvhSDCPYKU8qKOAU+iejxRFefrx
SCMyvCI5LaQU4Rn0izAuaCVWwWJ0p8/BmENYWUROl19s+kPn2KcEfAlHFUGQLzdQ
irqe+ieMvInp00P3H7jwuQTJbXFH3PXY0WM6ehal3Ktgd2r09XwW6OBjfXtZ0Bf6
rUmRgPqcGm/QGzBBbR53jJLK1G07C1FQ7Ro9QN0YmL93oZ1oaCsdmqOtA5UcFUEm
u3q5SmkN6orRB7d+SikIIsbNRIVI32e6lNqusMH7PoDJ95T9+Q8p97K7LHC/tm06
rgNhfHhyVxsqShv4tgrs/BuR5S6OXucu8S3OLBov8rqC6PT7wgjqz93hUDBdN48V
jjPq+q51QtAyLE7Qab7ChdsxBgtQvu51F4HKsjzRLlB70FqSc20aF+5PfnF+UHpO
yCessyJ2YtllvVuy3ViViUYIVd8IFKfiW67EBhp1BK72xz9yP6ZqA7i/iRqqWUVz
EjvB5LKiFWjX+Nt9NWhVL3GIFhy6jJDABQe5qNJUghOO34XSYYOowPZ7YLUigXYY
gQ6n9IOeogPpzU6Q9ykkdiRc27kUCtEYQKpNUDuOQJCGLW/Ws78Dosr5QoWBlDyg
E2HUs0JuXFjI88RJGJenj1U1QWTPJWCtmkuO1qRu/4WlbJKO2/bQfbIu/61a6x2f
YwLPs1vHEf5H9L/Re4tspPxGl5QS0ipX+o+pocN+wBL9wzHu0419IzABwecUwLH0
H7/r+HK467eq9avuXyLznf61sXI3q4lv0hfK/JovQ3O9iY36uy3vpCZpLWWhHF33
2PU13oK+B/lIbA7LniZCtASfL968JC5InhpXmgYzw4jYG0ZGor0NCFG8pOd/YxNc
bDEHQAphzFbq3VaoD+i36IVEiMKNFciZ1iQrQIkus1E0V26SsFmTmcrQCQIneW0Y
z/vgf6b9OauGOeCii2BSe/vaFnJf4zO/JRDL98UAXhnJ2es18p7R/EN+ljmcgZ/L
2A61Q6LXJQYzcbKI6tdGXrAA+ixkkzzco0VjB7iHSA+PaS+5xIC7D05bpLwH08DG
dApoFnfANYSsUMzfJBRu9k8O+1OcpnKrOvxOCQXNadzEdUZoy7Cbag42J5RReC8l
W3HjlJqq5yRun/ymK/SLJWydt8Wliq6z6HDkd5MvtC/o00hZC8GkgbfWsi4wfi7p
VAx6/lV11pus0N7FTtKl6ScBkr7JFcJezlOBTWeNfMI8cFpPXsYlPyR/YlG/dexG
d8dIkdR98TLnKL8G9FDytqqYBUcPHDSDXRdquH8VTxhuuAeyhbN/sJSEagQESJp/
qAkG228WufuGLun40nIbJvVMNlqn62/h/ORCusS/7STV6Cnwo/PESpLPOlmGY9Sd
/ChJC0iqyylqTEZDJN+2o6GjzuG1IBZb2XFzsssh8hXN58MjEG14zmbmEHqDYmrO
RzUqWBqMydb70hzvXFapFBw9HOeCx03uhPj3SoaJY+vYwTf4DYaulHG9WvZUNs/y
yWtl4Y9nF+5UqeJNmT7PgT1ifnHk7iCDF3Xo7kiI0dvf4Ybr5XUTlXXnDytrrMMO
XcDda5Qwr5yN08xrFUkqhPDVYZLd8wBxj2k0cWrrkin9rTYLcsIydg+w4a/Q/j1r
bxDb7kdttA7sKuxu+ZItfRglrjoF0KONeQbdtXdwaDtOWGPAkq1JjfL+xk7jNhYv
QuDuPqg3oDqvFNrO1TD4I4CXNQ+degEoFUKHQDrYMelvRi3U24Qr+kMD16ipmopa
XS9EYIMKW++ZiIWfVnZVB7IgITXfOXzn29xeL/kl/59SchFOeg/GsN0lBWKWoNWk
jc6YmARqJklgWujq+FIaJhk11p2C6hxAoDqRUl0wN7tZeSZ0i04osoTyRNcZ86+/
Yg62XGXOew7z0knwKkogyk92UhWVPlFcTxrUnfLEHXEBAXF/3yxUbiU1Wu0DUS1i
nsxHyO2GJud2WhJ5aDWVlHBnSpG9Ovxc7M6wUIdGX5FAnKlIUNkjAPEp/43ZwPxI
ldN7fZzMrggjkBlfC7X7x/fKFn8GE0ySLBrCKvIv3CuGgfZJ16eyCOCJKjZEOt4e
jJz7umxpCNU92J4Yt3yVUmEEDTc+72S5b8dQ6p3O83/Zn1ByAVJNAYaoVDYDb0tW
QEdn2HXba1baE7MZgi48Ox33MK9lbT+HwU3jrouRrxKS6Njc+I4ZSbSHpKZAFJFM
p8IGod07BASDWcF1IC5crIJ1VaQr98A4n4UgsKp/8WAzEpEQ8lQfVwpxSD0FifpB
GlRsgyVsU/pMOjiW8wAuY29sp2xQLJUCYVBNt5fMmRbRGzWp2ESTp6oFLtf1tbR5
ZfPkWS/7vZ2ewJCju4dV1fpgOGYAomxbrvXDUwgTsvhRxJMN3I1rDTQ7KKoJaAiY
TQURYVQvoDKzK09ZOg1dWTzH1hiKRggdiME00K0MEU7IAyIEPcP80TTQKDLoLG65
1JFicpZgixrlTF9g1oAbhb5Rd/xVOpin1EUTTKDmLvoF3RSETq/+YASjiaii3fD0
eclUwpzLEr8C3nG3Z+HXcx+/U0ABgzvhvFZmr6tTfiHj3/U+/v0YSpkrkuXvR5OW
jxfBOuQPPOCCSUHnU3iHIQ66S5CgNrZKcUyGl2pStGca1RnabbABmFcYdCBL4VT5
GpEahzfLLVd5vv+0SKQD941PZcvmu+Dd6NCSStLtIC78ZyfR1YZaUnhI1kTFaeRD
PoCSLXh4xppzGR/Ad7xkO9Gnf3KKjc6fTVLCsu4XTV5FS4vvJjlpJPHz1xd+g5a8
NK80bU5SdC0Sqp+ATs4eQ7aH99yZ143P8PC9VJsQ6h61U/p6JoTxRXrx52Rz85NU
Pr9rAWGDcYtVGkzuK6ZBeIJiZlCA/TNDkh/hY7LCgmBKMiLcZyExAYkswYu/dlA2
Yq7IxO4NjRtXDW3RBkBO3vLnLHPemWLJNmrToUzLm8nnBlI5QsgAguY5+5gNhuWd
z5549CJkSf5We0qkZECP/d5TzN3a7oJgPuNCcFpc2rGOIi8chnGDXRMqUZ3sqTMl
24XpbSni34ammUrls6wyzSXDOfFKC06/W3tk6x8vmfeKwBexoolvvfSWNqj9pzl9
mO2v2ix2Zs2uILRMLebY03L1wAecgUFBx4l/sCWCZCx0Cpe9uEGC777VcvC5Ae0e
DPTorDFb9O7mQghxFKD42tGIa0zkGZ3R2nnYC2a/+ydwb+znrj3kFiGMfH92SVoZ
B+RcTsSKkzid1W7kmAmIxYnLZa9EEiXfsr8DfMOXcnrjkPryqnE6FyrCibEWtYh0
oSDHVhrdfgd4bmRpcdqlgI7/PMSx5JBvCGlYBBPBdZ39qyK3mqLVtDCWlNin/TMD
KHuKTKzwKPSbn2kguy8xVwyBi4Eze+a24DCyOMilf60ASMjSGaps/uBMwqVtQycM
LS5XV/mLfwDPZRUWT4B4eICEznQMrRc3babfufAq4ig9oJ3F1iWrIDHl/EZn29+Q
yCjlcUNREHYNWv5Wz4fvB7IBb6Msvn0H+MSLvoRbnscyq1ZImJpGS5bxSyKDNDp1
f29632JAzddSBmfqvO+/g7l6m4iExTMWROWJmkpfaTA40P2gFKNze4Ce9/oQRwQs
Cy05GqTpuOeIRkCFd+KzomtkAIHC3dWi1kXwFMpkPAwPeiE6fK8ycKz4hxYddoE3
hRU3xXLzS/dOpGDR3WEEo49pFgpe6E4Pgh/joS7EAjI8+68mHHeAxzsUOXnHaR/U
yEVgGBwRHk54+zxtc3UWIDYWitBQ+b/PNLuln36E7EZDchAUJNj4/foBDoLPofnI
+wP9IxYocsb6mAaIvQRr81pD+4xsUqIikDICfs6tsCcML0MGHiaZ9wM62pAgqtAf
fac29lBh+ApEEk7yavjJTGWNlNIJlMiK4Z3jxplBHGOeaiS8DH3+FGPOHqutPPlQ
SAzTZp5EWKU/JzYlbc85bNaP96uAJBrgEA7E5L2iVHN8o23XQdMHWEwIkUlfWE/U
QdCvfPEkF7tAPLTVmEzRrmCGyz0PMFEQgjZQ68fnXJ8Y1CMoALR+2J3qpjYIuV/V
mYINSNMBVkLQko2BdcMfy85G46a82tzT3qf09L9hdg3l8YPbnS5KG+WyWDEQhSZW
0ALMSb06MHF9fkKTEGj/JEw4QL2WgEFwIu9ZU+vlldkOfDMWVQfxuYBSs3dRNBAH
iy5tIcUU3ZwY63MZA1pWuXwRnnz9uMI/Kk7PhByGZm+K1E6bHXXv4tyBR0oOMoKR
NFJMmUAGj93zxVBJDfCke5a0sIgyARZD2BdcZ/AdHyjLAc4zwIHeeox7iEQ08qpI
c+ALvKpwvLX/sY2ArVDB+F7yFGqAp/abGUL1qVxHYgpE2J8Oy8R38riBc0MFFUir
ZtTZeyu0WjHPjhJ3UsNM8nZQNT40GmXesL28tmAty+7IpoOX691xbSxMjTM3Wm8i
086aBHKNHP3uqr8ke0ZGehUceneRmCG9tjN6CdHKcZ48YRCwnY5mO1gQfNEYwqh3
/Tkm6MCExGKgpmvB4Jy6fHCZeki6j5vEMrHOAPe48YnmzlT8I6OqoVvykx+idzdv
2hpwn6q33cyjcwncdXzL2HpHzoqOmcmGPwamlwQshp74JclpFQALWa0++d+Pe67E
k+9jD68F5idQoOONqBxPRxj1V0K78kZv29Nz3QO+iD/TRuhNjqI3Capc9u1Juwd+
krx4Npor+bp+XdKfmfLVCV8ZBu4FmtObur/FA4FpjXFawZYXIZ4sAwltNsv8xK6J
6k5MfVkPAGq7ipvRgN/PzsjG2Trh8EL8RRX+8Vp3V6eXZQPE6FvkEhbEOE/DFwMV
yhA7qeHUHTcA/1fjpCRFrcZvgAsVUQLe0iD3pyUGDZh7chJKzbwLLKSS1MnAv82R
NY4U4iJTdwvWmjLr5feBAaEjupXosaVOElIavw2Q0HgJvbHEffXyEVpbGOQPwIyP
xy4MLylxfrVGJwSq8RgMBnvSWFpZIIJ/B820cjlzJZ1/VXgWG+lfSJGFzj+tx56/
uVKf5L7j/2AfYm3Ym+GHf058BHdWqnvalXIsIC9Q7M2Rax5Q/+WIXZoWLq/Ey+pw
QlonJKioqjYXXcA6OqVjB7QKG9K6ks/RTvCpnGpysiR4b69i7Q7PYtIROpWSJ4F8
9dHfa+3sqXxlOKWaEqI2GZqYEtV6ybT5YorSKWXuouKTWki0uD13qnfuKqPA70dY
zsNJUL6hse0Mlo2/z5krvSaEBkSAHxhH6uNRQBcd4cAgMd4xUAkyvX/0dBFdKd6o
HFklQIF5MmsNfnnWPt6RlIgM+MRRDfByFksz658OTrEoQ3UJ8cFRDq/bGZy7V5tX
gjhwrmhwdhC8yZHo56lBtmIblpa6AzaOmg7Mnk2Fxe9yALwNAeMCaf54t9ebT9pT
1f16Orpt6ztm/rvQkM6zJETRCvGUgBGiUUh7wR4BMGUWJn/I3/yn/D61whQK+H6s
UKUOcdgoMe/kOytuBPkOjw5p2v+et1HgEOnsSSyqOzJGVBPzTpOQ7cHj/HNhu+++
j8nNKZ/Hr9yxBIIHvdzwafgMpxd8wemmYIURNtZ5RZoo2OljPdCgAOO9NBhcbi9W
Qyklf0sV4GoG4hv1bWJGG8TVWx1aM2nWB5Yyxf/K6qM606UaYa0KV9zJhwZ2D07h
RZNxfMufAuHSJCqVJgcUXHBi/Whtc4z2m4UecuU5EghHSeny5mjR3HCfixf1uqRs
/47WgFGYP9VHZNEdHbamE+HH20Bf3VYd1oW7n90Lc3JPoXcENNORwbQ7+vrzlSH6
dqaH6zkC7IHOlnFoz5G8e/LVpnEYyEIN4eYpjeqfQvoDDQkTSaBoP0nFbHcYSRRN
23E33btgv9LF4bYBWvLm29FRon+1WNOURITOE53YawLkrQVfqQvCuL6mldQaIMWm
KJi1A+uXtFOkYpULMvwybqfM4LRNnWb3+n2BCCiKBLQqieAzD2SLrYWZjvaP4xxq
uMmRCVlDRSewBvesdzKSmT913ic1YMHzOqTGxmDYHT2EVR95u6593rfDYhLF+b4e
di12tzrBoqBhm6jCEAGtqN6VAJZhMgaZW9Ls/kdEryPDfWADbN+aFM2cS880aYoE
lflrnVGBllqDkLcUw2J/xTjyICWTQQvwV9zXQgYUj97ZcejQGPY1NwI8tdevqYCY
c4Ufu0aBegjU/UhzcA+6y5CQIFnHbdxy4twsvAq36vFhYgCLn42hF08dPRc598uM
/GA3//+pVtVfW627aXUF+fBK2f/vi/23JHcA1dTXDAJvwXOL/rrkBgc6/WUMJLor
u8sy1aJtXzYvXm5lEFDUIFt2pXxPDutC7l2/SeMj/WyLfOdkwu7/WAaQa7dP59cP
rDagil8uNofaSlogJxW3n2vYUbUF2Z6P2EB9U2q2mVFv8ZKeANwH4Eg+DtXSRyOp
l7J/C2LWF2mRjh63neAcqMZR/7XuZ7tRrsORoC9YNVVKsRxG1udMZN+WR46/RZ6o
izICgDvhIiK90HduJLm6ZQZNABHHq5uPF9mv9BBlOondLzwvL/HDqXbXcUK6860B
S2uoZexFuIUzt1iZUGezjonkXMMtbe6Xolw3kHYMTih3q17xrgIcmLkphl0Y6XlP
FBwurR5Gm2TnCemC4NyMjIQYvaABAe4gObTkXK6YDD+ga4OiD8q5VYlRYBqWN8zg
4z7iHLZrAF/DDgG4pkJHKYkVDVfqQQMl7TqCa1sYzjLEbXrgPOFuIU4hi4wSub3N
6AD/OX35I5TOjkrBPgSDcrXhYFqpfe9mbXWcoUjr66AU3tQUld9AXVfkFXyZC+BD
UjWRznq9xLusXwV2KpDyGVYyqO5HqEYd2sBPpCkgi9YS54uG/djbvGkAWS/HbVTt
YUBxaXpvLm3SoQe6unlnypoUw8h3UJwOaKohdvN53lIQGiL2QoiOv5z5PHZJt6uP
jsPU/tyd4GBYrd7+bv+sfwHB6DcRF8w+ZvGSEjvOAwYtB9xMMMw2PLDluShA9TcW
AQYOv3j/cBs72MaT+dzq1/3WzeQ4YvPGoIDruTs4awHS7A7cwdwUJ3fAN5GiMHU5
+jVH+x3NI5mY8yoygGUtmOnE3N9mpD+kCTE0kFBU9ZBToqqcpidRyEoIPEDx+Qk/
ZxPs2NKLW3S5m/86RQgzUCUWYhPyT1CNHHdtEzLW4lsgWwmjQdKm2s8tKtfNYW06
JIofvnvf8Wwa5Dlvqcw40sWp47Y7A750ac35KZlmZQ63VuG72u94/pUNAbysdBoB
52/4bWotJPMsmYHfFF7eMbKAh+4AHJdDoSFXhoIH696Dm7d4XiCu+W04/S2qO0cc
uQpAQmgbZHZ+VBAJASnjRb83lfsJVgj1oq5b4Nd/Q4rjeitbOKcXA88E/C0q9805
wW7ezaCr//61sobDBzBJ8pCctHNEpERIL6kc6UScZ7oZWtiOUdrAqNeglf/lePx8
aB1CoFD6Y6ldpsLtw5Mag0UxCjO+ekENRJVkMTfctps8fp5ywI97sU4MzlI4uaHh
xq+sWhtUpIyTqIe1nrUN4YPsp9HyEO6r8faY+8chKETesjYfWOdbU2qKAX08e/AE
aX3PqC6eFjqVhREj36F64CC81a7Dmg7EtTvPJ276w5QLPINMkqJo1oFANy9H8WzL
3PsouWUiizESwSNHcbSB2K4hHItY6GnQiZNlcEC8wYOya5KB5ltSpjpf5QygX/bf
FFcB116xLl6oy1hc4atE0fTAjoZ6C6Ii39WaUUOSCI7OvPQmG0nWL6p5ku/Vuqag
uxH0kLnUeRb0WKHDP/JP2poQ2fVRAdxLk8Q7QPs/SHDJID7aE+ZSaH3/VMcVrJs7
SK3oMlgUeKDxUClboN4xy7QjCOlDU4Tkh14c8KQvxFonp0aR2+2W/Ll5i4KMkZlq
NV8kSopRS1yz1jM5GrbJ22Izifvju7oZw/nGowztZJzd9V7B/6P0YnUmkRUJS0xk
qkH6K5odYk0s2aX9Iv2fPHF6DYTROTtBeLvIbuyN+3YfXHsGA43Hragq+izv5Hi3
Fy1A+83QS0lm+QCmvSZv6diwDjKzqfTcXMRdi5sCWOCfqdWMr+CU92zLtVjm8nxF
X0CiQJcidBlDMB8Is2vCUm2p5X/25Z+xhPqY79mc3+wx4ngxtV7d/SBMIAsDBBAt
rsZ1np+OCM+63LELS00ySPMN2kuc250E18yYd+wevj5/lSrlfBmBfMsKFMIImA0n
eVfS54y6vC5jsMHKwlsTOIdnrSBRCUDsNAfRNUU84bauTROYwNo/gbBZkVmlp7UN
YzI9wxtDIgUcQCM8G7Xa9cbsW/twrmHYWOS2p/2qZE06Wt3ZWWOmtYYO39oH2aQH
ZokeOCSzwJCZSjHH3rvmaROvv3NCwrIMCo9ySb4Yg0hSKdchkY1X8yU1NYzZLBlo
4+QHfGEjelHLTASlgd3R20lpxuSqHhc8YP5suq2iEzmoizN5MHoAggHGEyXgTQ+2
pIlwlmfD3eIMdpFQsGeJmMoIgWAGFXULjBEq46Skv/k4ldXYUu6QYTq1bjpIfGL0
tkhLIEUwpyIMXfjvztVTidt9VV6RMlzNqkhSX16kvdlS0CrqK3P4P8bSLX/2RWMd
35ZcR0R1jTeDDr0EavzZPv/P0FcNNeh0LKbb7UYSSKYFErr6jJq1AwrW+FIW2UBQ
kLnoZkCgEoArnhYFUkvZac3IKtmVwk8+HRSb7bKvBFjmUrPK5JO+KL5IVPmZHVBT
L+TNv9bB3VzoThZ/uKK7FGN59x7XJH4IZz2OMKB+NqiNu5iCynrdYpikCx9q/+1I
IGWPo4DsVDTJua7v547sZzuRr0JTU6m0Izi9oTwS+qCZpNJEbZgI6LuA9FCYjzVn
pOzQYvN68AIuIE/RgiX3ehliHYC+kN9Cnf/utKaFSIRcZ0agaVZg0xb9I6Yc1BIl
Esji+hdLBc1DXSM7ZLjFmBNdsfBIrrsEXpY+we3IjsZZo+d5KwpYOcqVrqjAz+lC
RVf+e5CDSzWu3bxS38lDwEXFXTcNVEabmYpUdKORZxrgGW/O1FAhvDZsdXQOjsXr
MJI+luauaC/wj36bLc6convrafq8zxmXJfh/LNdl//3CWJIun/z0sBEGUxNQIeQ/
99E/trxR27NvXtB0eIyLOEnu0zWP9ZVmFqGNCeXozhR9FW/y6XtrSjVGIcTUPxLj
X8u4XZyJHgoIw3Wuzhg+SJRD5grj5ZeG1rMYMCgiOA6GUk/XuqaRillRUnhPEwI0
lkTBLI/ieTYAUuNzjUwrOMZiBGZ5zoU0iC+4hftRNHILJhWt5WX3cGdfaN+ZjcOL
27VL7l1ZKYsq9qkzPU4juACkv3TL1rfeNc/pQQnEI7FwsUeI0HwOhKccKtq8Tb4Z
N3EMrpjc3qXSU/QrrZnmcEI60r3WIOPLSv6JtGoOm1aAMD6DjkOg+bORpMb4855S
17PYSUKwBgNkVKr9LF5aJDsvARkvYP7OKoG1zjK52zZoSG8LlKd9ntySw0qZmUtb
NrZ9c2FfImL5VQ20Kr2Y6J1d163h6qAoRJXRgCzPPlKfL7iXkN/HD7TnlITE6yQL
i5yg7KkehhAzRbR6jtRRdDxrBNQUa4OhENkA5FgiaJx5tlcjUVDPNl+2TH0OFjEX
tmSMr80GeT7gf2FxIJE2pa6ykPKTn/vzcZhEga2K1iFy/KyKfl6Bq6zlyXT5zHb4
h8/mCgSNUfmUx5BeRRt1r66lF5+hFosikJijW6J4BnRV4Ys828ueRzexMtyWmfFy
OhLmtD6ELa2DMDoWf+UjkwaOONzsVwNXFrYrmR7yOEAvRvHCbc+3zyqOeUcnT1zA
eR6KK1ZslU9j2USj7y/NbMOuKzRpRNJF0z/BVRAf3Teo4HF6qg4i1cHhZDiW+8NA
wTlVCI//DAyGQMK3pT+wNmZSndIS2fOfTBQAwJON9sZTmfQTBm9hVqjgLwHqdH1r
CRGjTNXVObuQhIY/Nd1pVXrZza6aJmcRa6qc+2IwGKvyu9y5/KM8qU+Q3c1YZ+d7
EdgX5KfLBbRmn0E0ljnLHlWTQFm6+I6iffXfdSm1TUy6EL2LW8n8HWj0zuU+kUHs
INvpT4r+NsmBypTDqcwsxgBrnO+8He7Pztun2C6SV/nl9ORyqsAL6qGViY0NWaNf
w5rZxvEzzOF5BmYTmYDqJPUAK80Hl8VG1CpHEPHy0aBjpUDpMSZee9MJtYQ2XT94
XPRYOlMx4oAJQenVXsynZnxmeThusxzvjNYOMT51tbnX5DZQiFdtBYV52xliGYnk
OtDdOjL2rBi59sBCL7uI9z8qKlbM8tmXvuWV2NnDEdltKSDe011PDPiG3Fa32SX6
qxgajRY8Ub/Prje/rUsxZ2gm0D83KnNX5IsblGvk9ACNlEkd+sTcenGx92TuJQ3h
wqENF89Swb54UVxyqRLOvVmK6jQNnZQ/M29i9G6dXQH5kMTJ6ClOOqX2D8R0g3Q6
otwB/yYJkWPnv17G60RV4Et3ImTLm/bKrv0BpX2RoW62g82KMlgtNeIo9/3XP1Kc
vPZE9dNQ+BdTKXHv07o0l93bV7B+7E6pcRupx5XeG2n86vWh3upNPmKjx+Tgxjst
csAE1aywyA1qlsKaILOSSJLD0imI6qcNM9o3S1IgAY5hBfYO46Ai5BwqiR6b7fK5
oY+FL15jGiSklllBI4uT+Xn3Ln/vb95TMbzSeMhS0NMOItIZvZqNYBpSJk+SqG8i
yH9v4QSKMmVpaB8ROz00KMrs5pW1BmaQRmLRGXCMbjLaycnFnQvkUoLqW9bomoSz
jSlWZdxsMvZ/zRg0ljfufPGeSiwtpP09iFn5JKrPpHAD8whcBQXJxUsQ0cGxc7qu
K86lo4GnT6dKu7yGKP65ae6klWt1N6t4HNFcb3PgZcMRLMSgdArHNbaxf7FjuhgZ
cOYgA69ywzNFbnxpiz2elZeD9Z0TcAJeGwCW4F0nNEd3tSfCCQmOCrwhrPhVhvr5
ltkVVKwpKpDOnfc4G3aoT+vKAqQvzbHQl4RPE/ZdPs8BBxphuB27lPoKEL/UlKKH
sMCFwaBo9UGmsYpw6WsNuREtQnKqGYmi1L/DgSN/gOr6TpOD/Yn1Ngi9PqOSStL5
j2mfrg7nwTYoEAB7ZjHHDxpVU1tZk5Qer61wBWeHBgLQlp3R2Qzv0yZoiroL/JPV
CmrCg3pWyJzRH/O2jVZ/clMrtE+2hAuJHLgX0sdPPcOinMWOIUDR+8s5nFy/+kC4
t2SR0ZV00+47pPop3RxNqRsZK/GoyUhAQfEIefH/prg3dsyzeumyUZXk0bm4bPlN
1cEphWrjKV07aPAUgmyWLwMBzDP9AoznfqdSfBDPURnjHhX98EuGRyaZ0v1y5d+R
qvIa2+AQL3rsSIe9oR6AbzbflsogTmuzO1+b8U9lXpn0pQJVcfkF0Y23Xg7mKP+B
ZP+024L9TX9J26/QMqoGRs3LQJNu1iog2zndJGMaQLfjpxFg6VHBUvxMCkHM0uOk
8kesMeiUknedPVGVs9S6cE1RNoCL3qecABLGE83DY5t8ZYIVHZXLvtu7ikJmRycz
DvnlekgZhVZBhQJ93i/zXM2VdVpBePqorTjH2/kYcucw7qtb6wEJeBfHKvNUE+Fx
Ao9Xk6Ybd9CGTIUKRUxy+qxES88mul9x9U9GQD8+t+YGjufMfLsleqUqAAIbLCbU
ylJjCqDm1Nr1ZbPSq6DSQVSL2aeYm8mgLk6EHunQUlsjhKqwUzSGdzMoycDmAMo2
KoiYjVGKuzxAWdCZnOVK+V18oiwtCODDz/wBbWAcHcHiEruf5sFSVuCB3pIqVSIz
RgzRokbKXB6yCim/+vl+omvqiolTTZX+FsHJN1BraVmrHJ9LCetNVaHWxSAIwMLf
QFrDInGrxfrgeK7dEyjgbodQ2et3WRBzsMkIYl4SmRIPaioyoHFdWB3O2P17c5oH
Q1md5WDtQSGoI7TaDxtVeksjy1MLN0YWSMUiZpjLRmxGljgnqJJB9821Zb6YF/60
/d/6wpXp3lQOdhbxLNCcoSHZKWEs4r6gtWFKLQA8gnnfdILT8ry0Lz34kIZrcFpc
rJZG9ZioH9g3AHzjzLpDhLjRZugyOS6BKF7C1G1YXZfNpvYxT2mJHCgxKp/N/NqN
SPJ3xeLzHljkqJK5eqgmaAxRLV0v/QcbXopCVHhaZdYu4wPxNRqyZdb2MEJEOy82
GB0uqfrkqW80csH/J7GLrSIpQG4xAVen9RxxkDR/tPhqWtxjGi37JWx0m28+KILq
7fO5hILF6YCG4nEEOySRsbmokUabiauqAWM0bwalunikXgLQWVsKOCzfZyD8DcW/
bVbwBS/rfcl7XoHWrDmygfuyfATUUAhqe0c8zeOE8uaDqEMisrQ7sMkV5xy/pV76
hDlBZAQWjqg6brM1sF6z+ERDWmtBcUmgrT4DXBWMTYS669ZdENHJ9rdDbMPyAxeA
C+goKNngi89EG9OnTBXLS41BDkzPYEKQsJwPHJ6QBZxvTQUjhL7d6Sb7rrn9d3Uh
cA805TWXfPw46SePA13WfDujcr60UzMgmW8Mvy9T6cII1SdtOweboUc2eJ2Sbvi4
+/HFcXo+LOgklUxwi24ab4VwAc+7ayiNTIQxoYZWqFYr+Pt/BFM/NmVH+z1E6V3/
1MMIJfMvOkdWz6QcDQMecWW5uVRZPlRHk9DES+dPjpUmfaEE4sMMrP6euWfP0bBR
8OTCtoTXvlaaTNsQ/m1EheceQ3xyNRbeCbYHSF9XXxSBNfK4WZLkWCldkqpZM3Fy
1Y+LOTW/ymYYF3VPNsPguStyiPxEv2tXj9A+PWkG6Z7/Jk+h0WXBPH+4LPxsDpE+
DtdH0SKaISn/QGkrThRp8FYRl7OBEgA0+8YjXnMKQJ/tR3HJyBlGGuTPi8nYroth
tw47qHwDANfQXqeR3Z36gqs8z78VBzs9hMc0FkAJgdDkWO5PX7w9ZC3FHkSDuKc9
MUXwQDKHvn2KBzdmbtg9W4TSKh4//lo8xNbT0khe8i9xPOWOubq1EkoSq+EWXb9l
JIYZlI3Ef+xVgQhuEwZ77Tdoc0tlnYGCG3nmXeQMDilozmrAShVpyLRw2yeGGvSd
UhPLuyYzLrEZvme44EZMX0/lqZq2v0G0ffhQHkvVnFfKF4Yaz98/i7Xtkl0UXF91
5/OzzNv0v6PGZB5h6JhpZJ5XGnnSzBSqg6bq5auQo16YN+wHhyjfk15zA8M5gcGW
tnDt2jlGYW8ZraWKImSpErL2n0Vugi3AxJP7k6FHY6s9cFyTP5AVFyIXl3qSI1gD
AdgdhVshonokemUysrWvbSIa8TYvRf1UeHil6WNvaWYASi519bDzlOGV43YECCng
p8I2HPePHNFBPEHbyQ+K+azNY5Y9JjwC7XzNz6x6WLfnQabZl2jxjSEF7xSIwKHX
7B8ka9FLkQSd2IiX/6r0wVYIZ+Cyupu3b4E1G9pfPBJ0o/LzSYIrWrc1ysyC8d9E
nWGFd2N0bJEummwMcWpBdB30MdIft62BHkbZZ3F9xuT/nM7wRzPlLgVj4Zb2NYIg
7inGDp7/g6UAGpdf/KJYGRj1HEtPhAevvkbm6MWkmTgqzN4qO37dt+jMPCWl4lDd
ymSulNkhknb2g308toNOKviXrYQHu3mHS2CW2RHh+oDMHazvD6gQXs5PoSmop18p
AhBbi97yPueUGK0BnObDi3nxAE8VWVFRuKaiHrr8R2DsQ/kW+tkdOVqfyDwL5JSQ
NK1OSoK2RsseE5ztJbb8ssIPBFvVRKHC99aBmelovLvPWDgEAY7c+2fQzjDVZwEM
9fWgKVdLlyGlHCLCsHyS8W3oqciB48XHVmzFrcaGVPSiNLjsJFQ8BUr9pCVDh+Ek
C0ZpQSLi0M6Gv/gW5BjQxKcSoVilfqxWgaHUN37Uq5KexijXAGcnDBDpCd4L8Jbw
y5GfwnqTNCpEJ3embjXHGThttS6VqBvgBJkBNEEs7vaC+oG+h8o3QAM6uW8Zai1y
6j45SLyRQVidG6gIVGGCu7Dzb8pHdy7WdIofokXJWEQCdNigiSJNatpBX/ZHRuqY
87K+yHZJTByUtmuq1GvuuXX8HoWWwi6Yj3VInF5UZsRfZLR0wRxivJcCQWIWdk+e
vFuvfeFBa22d/Gk/aS6j2HezzV+yT0GI/tVKyrfJzTPTwfwkdlA6pgNqZflCIyhQ
qZSiKB3apkdWO/7b5zF10lJzBMNWsjULKGGHofU4n5f+vFNv9qHXv4nYgVsw925N
7vIqRSCueh8NcgZGMbbUD1/WJrArm6tl9Zz6W6KU4jFFKiSGzQCisRSwALZxe+EH
T4z+Rk/opeeta0H+eglecSQ/CKqXhGcmrOFmq2YocD/C2WX+2/zYvUBhpVfFkpJL
re/KJh42VcI8Yp8Zztf3O8FvSvhc45+g6ZhUo5mQqCJAarwuQqsystPNwcAQITGl
I0vg0Dmf3W4v1zXLCQD2LqiNjtdiuMyvtQwUcBvSJbAcu0DMYiXgWjnAIycDuGcq
IjZExN+f1TBxtuZ2o2sUOBesed8A0q8HHCRL57Zlv8sngAARFONIjKjLBiLqwPOU
NM+7ky0eouHtT7TYebLpWihMI/HFDnpPPSIrysyZ1JA+CQx/jdzR44gi5F462i+k
CxuxP8ahNIyRSBscbz9YAy8EiQKD78/kkirZm2vsDvsU12+xRDofP1CABKhexHGU
mqdIQHO7mVZnxENjia7MQ8vE8wtt3+ElCcHPhUTfQOCtkp6rqeEe2+Wm7k7inUse
g/f+kYwJR5jBYwdbyKpacQuAj+5s9L7x8fjafz/wf66zGVGLAou2C3Uv+6xSCVkI
cyu5Qwrv2W+CgXi5rCyjeLu+svRBmk9UC2fQ40eRdB0+RsqbSBJUgiFYptn+scX3
gkKkZLcPik8q5oKtWWB34VnHHKlRl8D6xACSC+prIDlfrsI1BYwj3HQulI+y6m27
HgXaYAtIDmSdzpUeGw16BNV+fNxWGUSaola5ANXgEHhZBtS1M6PU5VFGfEF2Dd6Y
FUJeD3g8h+I766bhnh0nouLaDcVH1BbTEflVEkYxC6r5fs9lic+7h47635WMiH61
O1V6XnezQQkJ4rP0r3pMxiozBDzJ0b5TCmGviCIuI/dvHe8IvQNrzID9ldh6ZOWj
46PBUG0I92rYGfX9SgT+M3fnVBAA9KK5lWPVifwvGNIxrjHea9SUO5chlzV5GNez
Vv4+JLrsT4k+934jQN2jnJzv82cdgPq9aQzjZ/wr566lflhz+xP+r65VPO34cemJ
CP+4E1ETX4vaIr8meUNrqVEp1Spe5xNkCNS20/I5DTHa1lBk8qfFp23kY4DlLTAU
rbF09e7LfYYJTSuWKl/n3EhzPm6QG5OhB+ZesbgXK8ZU3UNc/IjCMCrvakJgdkig
V0yTD0tSBstiGhM8EnlBasAv8DDmgJmzO23vZVFkER5v4zkSB+2FtnQS92rG3JWH
Yq2kCm5Fi5y9XCLcwa5WzBOiUndZQG52Y9BlGigweperaNaaOBAS2keXpZmBuLnB
DR7b74I+/T3AZtF92X2Yo6h8cpIv0xl9kmZykxVMfqntp8Mq2qSQyuTZ9XcF59Ho
15UqhTQ0K35018L6YDUe/VgVCVaa0BK9ZIO5fXqztzMkba1aEaKPPUHo0oQ7KWjz
/GdoFhnxgfbtme6K5bg35OQpfQikDxLmRZ5O1odjNOwymCGXbd7ERyL39/cviPwf
UpLVBbkdx7aeej+hGB3Md0JdCv0pDukjjKkWOXQt/qukTfLsRpR7R6UzplmE9uOL
ZbvqVpgDqDXqKLLNkZgShdmQfuAvllrqmDHGubhF7vQ1ME4ELfwPy+OOksnQQ724
u1u2s05Fjv98gc7cxaMxfDOKhtp6sZNJqi9Vk3LwvOtSy21EBeWWgF8JM8tsw6pr
VjnPaeZogSFi3nLU67bqrCQQ124ZXUd15D1Mwzz4NrINYHr+hrMsy6UrJ8k036uv
P491DvvzemoEJuDHFLzjlB9t3F/ZniNsOVOYhkb2P643Vt+9pZrngPjQ3cctpSG7
K7/p9dMOy1C3Zw5WV14hDsmndG1gzme/cT8mHntgFlFspMuhjOW8t34ejf8+hKsb
TVhQ35RMuG0jwARpCItpJu0p2DvhGYhLEsnZx8VlRXYzaO81JTUiOGwD1vObJq7N
A3+QFiAGKT9PhYgDxCr6kXMBBNjPFz3dLZiI4+WBWSXKCnJ6fQV+usm8hU+TvNG/
El1WXc0iqEasFgVaIzksYXR7TR0jjWkILYxRczE4eP1tbFlXZOBhKqDZNyCPKYn7
TBjeNpogluwXUoszYqrF0RpT+eA6zdcCSmFXsrb8TaQ6dmAkdR1feTE3Tp+15yIH
v8kFJk47++mS+E9uQXKq7SGvXX8/7ljqWxKzBemoMSkTKcgSRrllRHJFS3OVRMgF
HNrRwETypvbPgXoB1YA+Bj4Ccsu2cwuVTgR/CmON70eXwUmTduOL4jb6c9JxEfcy
JFKDGASjRJgbl0eEF3Ow4CYqLuOFwlF48iRLRHdqFPXyro600H551IXCFO/ZQlEd
M5Jmh9E8EG56DgUX3Ua/R4qvyGcQs5pUWlGd9kVsEf4rioMsDwcSMrx8XV0hW+zS
7/KfPt+Sa5WBGsFkMxO3mIKudEXm5W/2A97/6ptRuihtn1rE76GeAf3WGh6Uospx
FVLjA1q3a6MFMOBUOBGvayzlSl6yyRcX4iswYy7LnGD/Ajmnd2oyflEsc70k6TA1
pESrkcLHJtLQ3JUZryGf3Xi44GYNCAOjB8csw/HVkkCIeI3lKrISD04VbKUhAsvl
n6PWighObFyUyu9lr4Shm5ePMDmG7dcKTe9Am0uvDCFh6PXVaUTpToxztoa5+Hzf
yetOIGRFPH8gFuD8vqujKPHzxJcW1AhMO+wjuYtdi8qpologqwXqzy9XKfIYFPDg
0ip0bOmulqFW80F7EDZoF0snM45zzlu3xYgAhRMpDkpae1ZjnTWN0HONWKjgqIw4
ghGI6vaQolIaGtnKzYeDchj66jN4PMgVGiWJlsKO4SeCUCV27uXy9ZwLnjqYIJFh
davq52Q/C1j7NjkZEFJBT2MrCHqa5T0to8Ko23vwkVu5DemPkTRAJUwRDAv3P9GT
f5sAKiYBuNQs9deOpgIlSe5cNpRkNGdSJtk/eREs+qCknM0lZ2AdLfHnDFdY2Ngx
qC8C8zgnaQaw+qdNPYF8mhv/Q4nScTAsoOOHNVUJef7C0vE1OSKISGJRxA13498x
uhHmWLwmF5gywmfKxZwlfQBgoRC22TSamgbl7aFc/L5Lz1KRXzvDt5KJnkHYTvxK
zhpzZBeeFdcOKm2BACzsiB480mUnmMfC2wSFE6Lm1ROcnvNhpOq+GTqLYMxFvykU
ks308nkfPYU6a0bMRM7jlsIxVvtRpapbUfY4QcMfqz6y1ZoyROqNgS2vuVgh5c+y
RE0EhoCftMOOIREVYhbdjGR00JMelTprqKuOmhCQmaVc6f0Ff7eKj0bXgUHK/bsp
s1Q+PpbpizCCBYmsqoyG63sA+QnKJMsQCt6eNHBktC6xBt9Xi7SkuAFmRlQvHhMc
vprSvEMvDTS8fL7jPNHg54Ia/YxA+9AkZnSlflZjmwvclPkyttYa3dWtE5N/l59C
m4EIaZQk22YMGcpDFDPEVPa0UACamrRwFUZpB90EvzlFWdTgFiq7kRX+vJASWXHH
zme/RWUGxlriCpJkjlOY5RiWINfq0Eu7qDDA7vJbdAPolhEjy4D9IhWZ19s4BLFh
bXJfS25w7WhzEzjV4w7hSkZdtvRgOgYSM8uKZoLplBevBSEAtZ+oUe/XbiJyZqTH
820onQHORStU5N2e44af5rtQEgItmPiLN8eFHREsU0iTO3VMoy7hBZLe0lNUBohp
296gHCWwiBVamxh/yqKIbE8etzmbdqI/DX77PNvngP98kQSm19F9151urXQ4E0oh
N3wNZrwzLX4LBAE8rFAFyls9bFurUFN0B7rC1LkUutRf4tZt08j/4YqNbRY6sHJp
OHe5mnkhNpJSeE317eUGbNK6jfq++F2O0GTxCLrNfV8rkSxReHhGMdD349V53Pdo
HmF76z/NODPDu3Ww+fbsZ6eNdOu1ZuDbfmoIhOKckHY2pgdWiyWV4TZLXtLHEnAU
pMcABgA/oHFSihUJngF5qqMRuDMqGK4kMssdJM3PZoLsgWfKZZNWjhjmF4j/riPS
Jc5VyzbEQ7v9UmUqCKsz+5DNA6zBA8LpnU+glEnmJT9XWT5Hw+oHrB3lePtm8wjl
buztkjd5yte61zlsuaQt6sMJy5YUM7uu7Rb29gecgwfmqLRbH/TQmZhBfT6JcMFd
z90BZXBg1tZYXGzzmp12C3tC8xRr1pfg+CgDfl6PQutKM3LUvd52uxqXx9bGcRUP
h8NMQBrLSZ2jRASlGxhz2Cj9+49pmoexxlylxegLuBO+Jf/0jhImATvBIm+yPYnd
UXZPOO3H/IH+afukddXCZ9Hu7Dp4e/Pa7SzbGbgsJ7wgUn8Qmn1lO6RDDDHdCD5z
qNaGdlqs87hKMthQQgAEwCtO+ErN6LVM+ur/o7C1hyD7Fxrwe3p2I1sSd8UsbbFJ
kjDHTEnDolx3KKCFRi98mAKYHLuIjuuuiA4xFR4BB1vMOerDE3kEa+dMebJVlnL2
k0EeHauGyDAUYJBh3lY2HQ+zitOBLTbg1/JgV1nH1G8qJWmupJ+WiiIK8E9ZKbz8
CrqK5IycVnbCD1YCWmEQ+hYgTW3ADPYNdoQJfMLt8od4Ib77Jm6fuPDecjVufv7H
e7G60yjKb/ImGuBv701SZ1wlg6AvDJH8488u4AdCfoWV9yqHMsqaWMSfurJN2S3p
I0mJTT4Xu5QigrH1n39jmYorTgBg9k7DSETcLkmjO6GHLLtYWkntwMogPy/1LcbK
77YeFJRIYkDm41NmYuagNjcDVD+Z8FMpZYj9n2tneUP4qa5G/ewlORdKIvZf9wsO
dmNuOp3skkVgomXcEotFOOH6PqZFmlVbAWht7ot4cy9IPIVH/AVhreXg/+aM1PbF
A9me6vX1swZ08fr1ArtAzC7lCIP5H8Cf0VC+bCq2RYzTFM8e9EcDYPWgt/8NXBNH
cpxiBN83TZhc4QiAExkb8OMD2lppYMYsDzI1H5mAO88v98iXxI4HvSaA0URFje5x
DamC/U67WK7mzNH7QQ31A1s0zgns6UNQ4nZHJNIQ2hdQP+l6mWLZw61cjkh0SPu/
Rs+gNxpPvMKmJrAcz1HpIfBDBd893oFCWWEpCjUF5ITB/wUc/RN1q2wXL2Aqf2mJ
sTVHOGFY+2B4mkkjV4q3yij5ZKq420gbxNn6SHHiwFxlkt6B7YERklYlNDP7dwz5
R8OkhM6tDt+ttrvI1yhGYNJ2SzjgtIQfr2ykEjzlw+JTaNjPiwKQeuCUBQ9+pUqc
7jXAsyqeYhtFPXFjAVlYIoAaWL1I6Gke6kfTYebHfsNpezo7WngGt9aua4YwfNMY
moWegAtGucu3MDKSDs0HKGu/0Tp4Jss3Ao9nxBRy87GRMfsaJSer3rhHigj0HdRR
EnpUzeYwMzAxi9TO2LqbQn37a5aYU4VJ3L5yYA19sltbM7+lkSb+Hca1GNAwyQoS
ITFFWOg34HFA+zhWP3Gzq0dL7T14eNZ/Nkj3X9RgE4btzJ6lBrYUGNt7bpSBLEzK
iiCazoFTuA/Zu5LTlXJs1AFuDKlM56A47gMCLdixMeLUIIM9dO8r8aRJgwyzoH0u
bJuGYOYWV3LYPcjKP0+vGjFEl9w6lsk6Bdm9/n57bbG7VW9G9WdiG/m7Rocb4qCs
qLC0fpyZlk4PynFTFWjlLbvbpl4caLBFcj8O3XrpIYwlF8bYEyZXmzFcimMOgYWq
N33GdOv2seYQadVzv/IoIiakxUJ3938KzE3cguBXthnJWqOmnTyV7nMjRr47d5AD
K7wR/1/e26g+dZjX1se2CBesUn66utzxen4Gn+gu7PqNWX0hR8Q4PEVZzT+TpTgk
dw2FtYhvAwj+Yb7g75bT1trwJLvT/LP3DZE+CnCo26ppx2ITQaXv7Qc9HZ6Mi8sO
+tzRF9rRl2Ctgfu7S9xjg5VIWr7dYqv1Ey0jds+UUSB/fkvZptKqKrspfsiHQUE3
sVdgFikBc5Clu7lK/2fOMLhRcaCAoeD8D/yt85G0UYN30DxCREnirBAKgj00tyN3
wVHJCtdGZPeWlNXUL5Zl22Mq/+NYWRxMD5TeBIr9LD7/aG+LCe+r0uQlrespj/Tc
eseABPDBCaLxnRl4qtBv+C35djPsbQ9s+CPpxjn3I9WEWYfnmRCOpCn94RXlET/4
gHk6AA3Pd7BGR96lNR72/uPbC8WnqoSHfuMzUgWLohN47ee8qd5bPFBx+LnQW4gq
RCxyrQRFvEYRGfHzK2qx4tc6G2KospmB6oz7CeMyiiHw0+lhmEXDZllxA0MGPapK
PFjgAku+L2O9wIepXFWrL1Y6+O+s90vLd5szh8eczqb+U/7SnT/YiqYFI0YH9OdM
JftNnQWZwEAmtGmB+a+3VY+QOUW/vaAJO/SJKpXXmFHMHQVeEWwmHHdKVDyV5Tc9
lsxprkRdQ3X+ryArZIr7SxXKyKmxzFSvUKusw+Kxktj/Ph4j1aXoLn6z8hj0gNv6
d5a7lBPxFR8u8VUbXly36oZ24WtSAqbRRabJO+tGZ35wB2uJ1uwvWL27kZfwpqlH
cDWbC5jRCg+m7JyHL0/Qzc+y+EVYwwA+gB9UzFLvUTqNdMMhq8ohJPOULodBKMYO
Kon5u53lqS5w49nrut5UQFrkJhlaVbasXUs5xBxlcvWTDZsjgaD4hZwo7LrXN862
gFLPDq3BC0pWVJ4qAgSxC9mqLyW3emBBN9nbdYktmOMpAyckt1fSEvOtY2K0S/3v
0OxoYU6l68B6h3/mVWm4V74fNHL3966wDB6x3T1fxoAplh1n/QPgsrvJGGk5SaP8
sVTAv/Z6Abp1gjJyprOGqqyz+Xj67o3br3tglRltDfCoePh8igsjMmokgo/J9cy4
oP2apeF3aLDSqtXjM+ZzzMTOJNKD4fnx0ZwHtbiGQl+SY0W4er/8uoqkA5eOFV/z
DI0j66qpe2JxiR6wn3/7CvqISLtm2xdpfsOJPljTc1LfoXmsXC81rzzvn10NRFiD
4kjqj12UMZjI47hyAAz7+Jk2MJGf+joN7LmFt1mlvF9JIMqZswYtoxaJRIHv3FBH
5931TCSM728LP9tIlfUeCgcnCHy9cVUyTTv46tTA5nUglk5KzB/KLR5C+jhW1ebX
ocxFh8SQsn3uIvV9XggoXp5mD+2GsDKtaQ2T/qSCcRisMAcrAbaXvuPpJrYeRLzi
0B4VSf0JegIZvUlrqC/tBynmXbg/xnRRn9Vxptlw1gLYhgT1RjTkGJoKNT6GuFoS
iOmUKnu0v3DEUrC/BSnXWN4z7DzQUsQLxk/g7HDmqAawhr4GX0Y/C3igmtPdw9Pd
weuvlHLIcV+v7dp4PiLKkCXVTlOfVGFzR9JFwMrZe6RP+gi8wGBVOwZInnP0ehib
xOyb+c3opp/Ac0ANpXhmobKA+DvZddvok0SOiYIoV+SUEXVEoe5xXTBORnCc2/K8
Aac2uMuGVfz/FNGgSLHActmWcZp+7BjnpCrOPHE4GxDtSrx276wQ/nVem5qcZPd/
fZoMoNUNLdagH6QqjppW4W+Ohp6hEblPbxkZb0JXQE79jo5QxhuVpCuo66Y4AG/g
maz0U88W4KaqIRaxZDp8UsgjYpPAruWCzs4G2XhoZWfXjw9oZCfNMAvVzBDSteV7
OV5k+b1mO5Ud3phCTk2pIuOYhH8EpV9muA5ICdltjqtTLUOVbb52tUkAEADDpOAx
OcYnELOPk1XdHKfA5QMMDUfAS0Tyh+mvbNtFStyjV7TXFU345R/3JL3K9jNM6OnV
xhSvGnVwre4dPe0P/iDh0sFPPTdyx12vv9/Ti5yZJ7w/ZK8k0v4R5jh3WHUu4vBr
eSMIs5Qsc/tuzaz0Mp0vJ5huf6cWZH1x2laWonwjtG+tnJ5Jr9s/4da/80AWMho8
oIKruVW3mp+Y/DLoEQEXXPGdqyt3zX8oDZBhDq9+iyvnnmYJX99DfGBK6Y19Asvr
hbiQqWs9YNToiEnYSX5kqPMKwXeL9Uo82eOQPewF885btZ0gn31VQg9Kp6dmRg6h
xYhso8AJK4I4kHxZqpUlaNUu/8qiDPJwtXMft5GPUjk3/9oTVl0RNeTfdQ5IxpPH
R6wgzcBRSjr/QnmtXQQ8emsByjktUD9kTq4kUCg62eBtErozlVLIux7UVJXMxGlg
Tv6V9A8o41Y+4CdZr9bdMsVYIX7FSXXt3SzlCGsSJfH9PojbPL38V9qfarJcDFoM
m2qrjKqYTxAcL1ooCAj8LJcuKSFpV3jKXXX194LrcgyOo8c9UGhMtFHMzJVFu0KJ
jrpwjo7r4SHRzN72WmXbNbHIlKskk1yXUeb9h03vfGVwgQGUAj4T/JGBG5q5wktU
8yaFTMuCDrRUfhCF9kOx+aHWjH0Tc6ctk1j4EFE2iJxzzuavLc+YN5P7SxbI8p22
c2dlXGo1wwXoM3VemJwsVYSfteGaOj75LwYDfTXJoy6zu83uxt78etyXTssWwm8V
2A8UcVxp7KHSFqsz3rYv7B8kMv4ORxVoFtHFY53Gte+E1o34R8iRCRKfLzyaigwM
LgivH8CjWGTV+pC4STcZlFm7TePqojDJPzScmfbKUgsoqkoahFjzzSzN+80x8P+w
16AJSpXNeXA0pgR2hwQuOouZDNsAy6HCj5nVXrQiNh7ekjdjtE2Q8EJC9ESSYh6R
QimvgJ9iNhGsPgtHvJdWECuM5CqMCxLLzCgMsb1tBq3afRgOo9Fh511dKBvXKuko
Xz8CEaDdU26Npg2Cyn6NRJ0o9oPfNHLzPcHTBf1tjj3AAYU0diMTQ71yWC8gL4Yz
mbu4lv/whFE+O0odCscpPKea4L4MQY0ah/e4NFWZL/TcrFlUYzdvq8qvMVXaonlb
7KmIAyIGieqgOE69TapMdcDl9TM1dVKHmrhZGn04UK7ol4YOjKiqZ0JEZ9H2yIrU
DS9DwV79iCV/DDS8jBP00duccBzksoXLqTvlz1o6QooecTKwX0NYs7tgMf7OpJcN
EoZVN5igaOMGTlFqr8ppJh+mbukDfiFFp/sgnxpLPcdF4xJ2Lev5b9qQzd+meb73
A1uU2VR8666/m/GOkz3NcG/q4evD3uAYO5ObXr4YHHjS7QXYL55mZ9i/r5CempQx
HFS720HQjQeN3ZUCHT96rtfU2TreS29B4ERXyEoiHqk1souqXUcU0DQVdbIV6l2b
qvud9wcljliBlJKJ+f81J83ugWnkkuRN4I8gcVfPr1zC/hH01XBTHZ0x8kAEN+GC
z7E6mdHVL8U+uxHnDnUL9qwOPIBeIdOr4/Z4BAr3wpPnN/LahjzEhEFRPT1M3K4E
xJ+1l+n5gT12/MrElp3EykTJmsoK2pSWqmWIkkdHz5J0JdWano3M4cRh2fwtloI5
o2qL3OpUCt8uzATEHgWFAKn67pr8QEbiaxGqLhNgT9h2FqknwIawfeQAdOqLoD8S
nhOa/z6fwP+OY7r/z1w8kPyppY2DhIcgdTbmC1SM0BSHDfMEDiCeU3SCucbhz56a
0ql+qWiHCAh6ZG7zfQJ9ebLIbp9ccunC1qLosElHL52fz93zs7WoBBowGuMMFWCP
nZ3o06Q/0X5b/5BhD2JCG8fn+h8myfrs02Bsjx02S0ygIZ/NND2WbQMdPeJqjnLi
7UQ3wFoQViRuohKj9GsJVZqIxMXOD1mHlpChvSB78DOoA7qFYl52iN/nNBhueM73
3dXcWZSxS2loTHoCPZfub3uwby5KTmXG5J6G04YbXxp8ggtnKM9uGYwK5iliOuSZ
UAVP32EA3nfJUmgaX7H975WoYFMc2uTM95DFKtcecdH6c86ptaP5BV9YDySDqFub
vQ5PiaMMKgJPm3lA8nlSyxRZKkDgMBoEcw+jUpHDWjc0MPWmHYszbidR69/p9zgH
mGR0fpgxI/0OuAcnco/W5uCwJTZM+yOPPq3zf9FaaDTUl97L6HqaJBlJAVSv73MY
iiSHh+sOtBXxsr1O3zEGu6m9ICMr+kO7Cc15iD9Z9gA+A8SRzyQ8H1LGcLJM22Hv
r8XGxQZ6Dj5tlMgSOpUo0qRQodvkGz2Prh+RtL/mlhcJayjiq+XMfg7GfZw7i3Mo
9Rd4BFxD8AihJnponCbr8xHxqFCAgBMnoDCLV8iiC3BUHSqXGTw1BuheDN0IeLJM
h6YzOgBzwVIDZLjeRf0If+cOAbTlD4QNBJ/aUHjBJHgA70eM8nmXV/oWABWI/wL0
2C7Wh4Sn6dQP2XKKmKQkCd9+5xoNDX6dvODGCj+Qa3Qf9i2yzy5D1zAPT3r4jOcI
bg8IZojPZhQOK/WwVry46TIC3D5/UGcQcgHPkfCSO0VT1RCQ6zSdyRfKdDLDnDUT
Y4UIq1cvVG2CSR1YSmYCBOimzbB6VASs0/o6jrveTUXU6flw19ouh5L6uT+CSb8a
kYJKMXJmobtyzJcY7A4WN05/bi2dF1iYUV0aQ5+nnDPRYFf5vHHCzl2VLZsdpZIU
F/NX1T8ACsmwzcVfHupi252cA1pXgYX1ANQhG7gDCkZ7gPdQJV6b5f+KQrOKzbdw
ZSZB0WTe8N6O3hgfHSWw33FCJOtJalFOASdaacywar2FIa8V7pRoMbN737TIzkM9
mHoe1Wl6tJo5JSCvUqZIHaavHxEzLHC2xG24KHBOFQ+YBh7Reg9SWJxoE0fVx81+
/xySFgJ37g7TDMdYn4nFsqxi/I2396urB8flrwv/zXoiAhe5iKXWbC8rmu0/BK7N
m+P2z5trMt8Q6FlwccJ57fVC3YaHGBksbXpuMnIUcduOsE78/WBmNORD2rVA7Vpv
u5kTeL58lzj70kc/zAiIG1oFKiYxnGmXLb4eHDWxBmYFiSQOH+EELUky2vAYRzQE
Wml5gxIDRYd6Jc1BEaZMjvlkKJnhPswCsbEnnNyPPNoqmTxhVwZb3DVteLnxFqSc
29S20Gv87wnZds7XYs83I3+LrQ8RrEGgp5gG6b8f62/PZoLS3982/pAX6GFZR5OT
UbV3Fk4vrABItdhtlFpP4BKf4cnUDmH+6t87HBSUIHntreIBdsqhmORCXHQcT7Jf
e0gLPNeIK9G+7HamSSTJ0a2ofyHctqOCFD2PWu6lQLabD4IKiJKVyqE+QwKXjr1U
wPsUghZm4eNfjlEkWAKuQVlSc3L0VukMTmfwYVdq9E64pkRJFrRj9KzGDxMhUetQ
EKYkyppjR+S/tsLb3qUg7Bwbh+LlaEFohNpAcMcZs3WFXi5WcNpbf4wxccBt3Lw1
bAsikpQcZK5KvVzQaSm0SBY17b/TDw12oG5H9mf31ADHbwKWXgjwjCimn5XQja1d
2lbWx1j4ph1M9DuhhH81D0StC4nAx3QEFR6STHosdOF8Y0rooJFgLxGP39KRRZGq
AY7r3B2lRopPfPyw0GzGVtZ7/evI8qOFoJGgq/8/1B86XYU6KLjbyv2FyNnpZrjh
ixxjfn2nnCY9fQ5LQeUQCs8+nkWvfg5qMUBpx9LPJswVImlo8L81cjbQxrxaiuLl
Ym83XRo7Rh+L0ZkOuc1SjP/PEC5JcJaxrQGr/QEBOS40kElqb3P0LdI51cVxeitZ
gJ1MWeSEwxdeWVCCoNdSrxUEUy0mIs1NPAGL1a7imJNTfkT4VddJWvhUnDbTj6KX
1Ufirk7GuBwoNFYcj/t0CxwRmZq4Fln+4JmNlzaq4J2Su7wD8L4omRXvPFqZwk68
Mf6snGh+4tjdecyFU6GZf1nIAr4BePdFzZZShpZ4Kzygx3Qjw7T3OV/U4lZua47D
s5Q6QfoqPkHPDNLKo2UeV4+6uvIy2nb41XcbPSeZCuH9Pm38jE3DJ/1pNLKzM5+g
s9uv6v8K5TWFB+rhhBalDUBGYG4ips5F5t6lJLDi/FdjYpHkxujQbNjun0LdhpVK
gI9zRS0B24D4/ir7S0EYAcBzUIENYbB8XJ2AkMbJILfbkEdy9OIR6hT0FTMLh0HO
ZDopdLiw/Ga6P/wvdGP3S/eOEKCDlvoLOtFVMj9ZeOyGotwLoxGD9d9LRcRNpE7J
Eon+9CM6T0+cADvSAKROgczXx5NCDSWS2IGa/OeDfg/9UBb4uv0ZU169y5ZxKUE0
uOuZY7a/4tFMvpyzIcTmLE56dMppby38CK4RVbtLaZTy4Oe7bmMeIRU4kMJXhb1t
kROd6cgJKR4tD9TrIcCJMzeb1Rr435XAhSr9lokpp08dTz6UMUEQZLH4VzvXTDhH
gLT4SaiQMTIaH1SU53UeAKL0ZKVQ592a/SBU1WMtSTUJH8EBqF2rmO85XZ9T88Wc
N78VY7eTaE8rBh7KqzDXJkrC7o4QfnS12X7AaBqWbhhTNTL64nLwp4vVY/cZtsX2
OqmhfVFD2LrbBQ+bO3geOMo6JUvFWwhQPoatKs0ptxOWau7Dv1Z9ZgdbmHCiPyFJ
3ClnxRoiXLhAlO9JNSpDjGnfWOaKvVN4wjc2Y+ni134Bd2e78m+rYiMY6uQNKh4t
jcrDoTYknBSL02TZPCF6dtiPHjQ/da1oTquQ/EZobXlZSafVJxZRlTS329FtPa7h
ypVOFHhX171MzQ9iCoYtscJLCrMk53hKOcHZnGQmZtdlZFpPuyQtu4D84n+Lq8OK
jHrM3dvjoK7tW7P4AqRqYklvC55OkP3fPXEWH4+OS4zj1oPScck7PkOxaGvPMJUW
gLxUKd25DrNusDVTEGGk99WYoCMdgQuvPjQ7MCRLQ1asj9yI0Cen4A/SL64OasQE
deJ/F113L+5AFwKBqZSJJ+6tg3pjlGjs2YISDc0GWWgGYREVAu2V2TTBiuLzp6Av
LtJZhSBYpYVYmw7B0tYqG3igZdOmct2tLqchvFTo1d81eujLnH/S1/QNX7Y874JU
YUUfQt1nz8Ojpohk/cSXAI5UxDNrOUKqnBdtdj6cgGZdqwaZgTKGC+VPr8g6WlM4
72WzjXqz0NMYvFywjSVdCO8EvdPIgo5zGhFdlb7ZDYmnY/RSHK8cQXfiZtpY6Yje
QtFZT7Vdc0zgr0QY3b+rzMA+grjF+DguLImO9KRWjTIwd3a7xERyiGlLMpnUilni
p8KnzyJIGLIM6gXs0HIlJpx3nCg5JhCwlmP62iw3Kj8rC4MQF0gsm6HLq9lULqAz
FssoXzDFrtU0AB2Id39ODe7XeMZC+990rj6qFd7ipxCirAO5B0FR7CKWVw5ezoKk
Yp+qYpFVW4CAsDRGKnUnm5V8c2/YUKHk/Yet+zHAUHnz59ZbKkQJgbbBEB8WxRWX
jH5+wMPM3aMyApymmnQEpXzwbq2x8qyjL5vGDZuKbfar1+JRNESQO3z2xUxw1KY2
qGzsAMEHGZceWh2v8PkAVbXdbWQpZ7Wsh2mzRltTEcuzevCPt/a6rIbI110DbIVH
8g4JZPfHHbQSkGz8pbSIdvhWie4UdpuAW5SC/6Kj50ICGnH5OB6ZanV/dCfA3sCX
WBgheLe+eEXYrrxlIRL5YPUwpSWr6Tlb9iS6Is0uw/YlG1VEDRNodD6kPyunsMWI
qLx+F+yroe5UwzUEd8QHP7cXkCd4R8s3fIs6q/nGpgmho/ELDTwYbczRKcebkWcz
Se43tpCT5oW9dGsxRwRAMcK5Zb8A8pj9xwbBbDOwk/DHBkmTl8DuFAa+sKihq+h7
qhUDrDI+HUnMuQOCyc8xybtsOuEto5lPaa2z2sI0ZrDB6Bo9LiaJoMb0/QLeddnj
TFbC2UdjMWiBf4Ri1lUqoSo0opg/+l0XYjKJQwjx7S3d1gHiqp/AnFEd8KyqAeAu
HqZSj/OmD7sQX/mLsJM550lEY4bGwqPEHHCDEUGtPieXIYhKd2NzXJNaYctC3QWN
SRuhYh+5s7LJgGpekPNo5s8VjMQkNXVD2awksLcuaUCq1DucrRWuT6arDEq6ytPg
e3jFW6nrYIWYnKdKkyAiLGtN/vvbonuU8dCrXQMMx1IDbo+sKqDZzYlc8xDxk2Ow
p74UOw1mYud3k3OOq54bv8+8xJTgsnhERtyufGPiOiCd3o4Xn76ymWkhZ+2Hn3mm
Of6hWuT50eFxJQXuTh48UYCYYre9awmAJe4GxMpIZRzolCFSWt6i5M8qTzQEVeJp
DmSQPP57m8fqoYpLFQWuhpljVoPkFCme7Ix4J/mUXAFpy4XhgN1YTWnHgZBlDOkI
n31O1qo+5JqVE54y7gw1AgTtvC+sSIxUy0HMbb+Sfk9e3g813O1nJLSGHEoYVWtn
qCOyJJgy5WzNzDutIwhOYOgaMle84DgZkv04TlHZaL25ub4zcvlAWncDNiFv4V70
4JJQrx/pM66AsDrxLIP20aF8v/28QBf2FdLp124tW9aOplCWXv9jXx0ErrYoYus7
knh6bi7w0fNS56H0xeJyUNYcJwXj8CU7U4rb8nrNUoCSa7UTjevxL4abYem5N3pV
n4YhHbbkF0CYi/lOmANQB7z0Fnky6jcU+IrZ5AtxWz7P3G4WH6p+Vb9yIN9l6Y7Y
NkHMB8FIKf2JJlR6SI8Q66o/iddtFaQNAyF4PAOsURrtqyyxpLp/4z58symewIu3
Yj+nbIsCHvpc5Wj6R8cQSRDQfkRMmruszWApYpXyGzGa1jY4Y2x2VBaqG7h9aNWj
h5fYRIiWLpXYKCZEGI+SNipF4CVy9d/EyDCyKcFHJJWp8/NOa1A3N1WZoPZ1B7us
0A/yv0GJeFrpDE3nUg1l7t0z90pX6D1PaQwD9ezBj7kvOhhhdu/a93zmSaASCKDT
cAPPkFfqlgT6+9LJcVRWcJUg6sOBONUKgZegKDVTdcItFKBmCgGx5PnDzM4nmgFc
wwMLoMck/PrZzTZN4rEcn9+kYnsJLMcd7eAgNu4m4Qwqt9I8E3/dVeXfDt3hYN+b
Qfu3kuUr8vd8d3A2FRAFlmuXU8kFnPbBbjUgh6T/YXQOy9xPbrxEoIYGWzEjWn5A
GO7WD6FHrfNBg0Nz/rwk9XFWZxh2JK+FNmugUEDz2yJUoOdCzVx2zhTQm+K4L9mi
pqiveSZ2yWyZ7gkUaJV2yolEZD9p4aoNGj7j00+kTE9EJiiOLYNLk5MNs9EXlPJV
FUGAIjQEEz5e0E9YHK9LRnw+OnlpoG+yq2KuuxItTisfps36ybT6ztmc/TCgFTNX
Fq7ZRflC0TqCIu7UO0JqreJHhHANoe8blzhLa8UvuwQnIher/4ZE1lSB14tCZS2g
sUbNJT3b0RRAtbUnakgFPUuNaXq2xgcwD5vuWRcgb9T7w+IKwWuWwM9G6kEGWhwo
uHDsMfmnwgcFt8w4+RUerPFrwolAuxUKs9KSsdYqU5HoPmbIKwK9y+T1QAD+HHpF
Q36HQ8j7mXmJdEYgiYVdh8shAFgy9nlITOgsEgT70mAws8ikLhJHpgtHu1mZ5gEB
7sh3i+9M23M2sQWsMMINsPTay+br5XUIEm/HCheRjsaL9TokxQSDe9C0xCDHWAkF
nMqYz1Rj6uSwbsz1rDGJBGnhMCuHACmRIcpIWOaePnv4m3pArv2OAyRMd1RmoGS8
TJTmCkCXKnozna0Mofro30ed6ZzjlAXWodn1ZsMMi9wQgC5dr4RQtVGw9+0RL9yl
BrnYUt9CfnLrNeQa88qQcpsdCKI1h1d+PMlaVndD7zTwU0z1TgHEmFQg/xQ/mLFb
fYeZ/RAz8kaBT8e+Di8wKGo/X3h0c+bkTeoNplRgLlIUc2/alhRApZmq8KpxwYkY
vUsOVmJYH7Z/n7Txit8SpvFOmaN68biw/cTvTKQ8eDG+6Ap5/awgukm0Fx9cBcne
E1ucGCBpiJougFKAJa5jVicZYH9Y1u1kVRYO6Os2yVWM7cnCsFm546RO5Y9rSGsi
TJXpExPkwVUa7ha8BNrZaLc8704WXq0hk2EnEjDVq+J3jM6PgBfOmH8B+E8ye3Su
0WFbCLCMlfGyaDoQTIORWjTTxGt9WffqEkIZUK4DcinKna3296TlVv3P962fjerB
CSK+Rfr/WFNtfR5cVhztO5qFkvcIldVAYO7fMekJhJQ/FKJHAM8OvRhPHYCj+bDc
UU3EcdQAjJ9BGMjYH9VL8Aa8NSCQ1rwXkNn1KqWOpEALOEy73ivVvjm9Z6zIzlCA
gTJFySd5WjeymI9kBLvndxGRrTR0CFsqblKWdwV9ddkQUJefnus8LqsgLD5B27OM
9t87+ztmdSZnfMyAY3kvfzmxYGDYCcXrrKCBq8rjqh+iOYYZjYX0xNRLPodD2Xy6
YZhTWrIocF4GXsmiCV3o99BDYQ+rRk/5HZ8pethO8z1WFXZzHmFyot6pKJw1g6PU
jRf5BqPQXrmZVae8JOqbYzyQNsy5HfZNZCDdMM74FmCc8spNhnJVHwVT6egyEQew
p6y7CVruu/YVeO5w9wOXrFiEy3s4oZI8TU8FEyduAx7EzB/t8vosgMmpq0FNNIZX
uSR7d73PQogu+aJsAqViMW351dDsqETNW0t6uGzSBmZNHdGMdjgn5VvHWIJ/T7yL
RTrlIBQHAPIOYJNpK1p2kl1lcyNH6pr4ZvJnSyX83FBtjFaQvEYdJi9042w0wCjW
7LLGPG2FuUKCLg058ZBZjOXYPpAA58D2sT9luNCe2WUvA1AoJPYu1aVys+oAqFTn
4Nj3g3PgWtLwdLoVKF97ZNMc0iFa0stPTPuRNA/iUr5Y7gX5hX0jXRRMWUAkjWc9
nvZoqC4zYrW/exTe7ODe2J81Xo3+ZNz26XMfG0mUZdM6eET7Km89FnDFfB+aTVkl
2Cg2YbK2qCYEruemo5e/pd7MHsqQyZOIfXSggNkqwXbkLj1fcTwP2SwDZfdr2I3k
/tafPPqsY6UOfIvmDZmnP8ru1MEzis4X+TFAnFrjx+XYDtZ1nViSrmkqhq70C6u+
P7rRYEQZc7PH7gCpK67mFy8cCiuQeJqz6xlx0wDpHv/aquA0Sl3eL3frTJkQH21S
2XmJIf/DmVhlrw0sSmOehGeysdV1drDOH1dt1JrwBSD8bOgwW5lb3yYhDab/7VrA
NnCpGgZUys9Hc8nZGcRoaxXrlDhGj++4E7N386K/vWpswFH+Z+3yZ1Fw9P9GqOpu
/8w4tPyn5Io/GogrfC95le3EkjiIMltukMHUcyIEqSOYe5brTCivQU5fPKfYiwkP
KGVCiXhVuLzC1gf+l8HiwFr2frM4Iyo3+OSap+nWXZsBwXHRXZq7I4Rm+U1fexOn
eoED3v8b/LUbdl1z9346YZQUuXTGDod4WuAbeLuHrBVmr1ClbsCsKBUSmrF3tAhP
hbGtelK8Hkc1qUSCqPkX4GgS2ONG9/zrO/ZgzFYwo0iIG2eBwxdXFM5GXFurUi3m
Z6jZ53daYL8FVugdFaKceX9XiFiPGF7NMKMDMpQkv65n/afwqkHxwpEQ83DZyXYp
O8cZL4UtGZQrhc10K1S/qBlqzWTKPO+6Us65G5FnwBLk7GyHi+4QwBitAUDl5wie
OaY3P+wv582ZLViVOGtJIPBw+Ag2CJEf0MUo18aPQ2XQmB7IGED3cXo1Gi6WRgQk
UZD1DtMOVuBrrEvAzzUtkN/Cn+rzcD8nDf8Mae8alAT/cy1ZgPW5RCdqN6Jd0dQN
NYlOdFPg5AgP8jobMfJBquaTImr2xRnRrL0mJ+fVuQSVZYnwLQqWjoePTgKq2hoW
BPfhbyfTcuh6VKHHr/0UlfysHZt+Ez5dWBT8OgqSl8opweBdaKInSqxGXOxdCeQR
T6C+pUjD6oWgVDJjcpN5SdpzJWvNFX0+Br4RT+QzQcCZ5yTMqD744wwarSB+ih4K
S4qGk8vd+h/NsdUYfBb4jZrpJCAipyHZ3j6vJRN7q3a9bVLsrGvGuFVzEj7LCrra
PSF1KcQS1s5VDMl+DJ+8XV0dbKJWtdODZoC/X+ybym+4hP+J3N9oevCpk0CWi2tr
ZHLfmESCJgkqBG4hWOEtVQjR+7n5JFqWTKH1mePsCJbMAwL0bue+FoRxdpe6wBEi
8aRhl240jvJpGHp0AOMzhQ/4S0YDek/pcsgU49QRaNU2k56etipVQOvkHlOrRC7H
8yInrKxa6esKuafph5k56fqCvtfuS29bklsaQbLGXX9nQNH2+d/VZfkUMOT3dGRg
y3SqUj9/S3LSaFd4GiLoyHUXzdu5i8BSf1BefcxaHzaaHwIWsbrQxLxwpieXM7GS
6rrO8B09gw+opuYjNCd7UdacK1oQoim+xc3I7OOH5HBpSFicrFKR7gS8ZEphqy/y
XW7zf9grwptjawxMiOOr9Q8eXlZO0a/46fnNc5OaxOr3wf0EY2ktELcd4FRcqMVC
9hKtHevg/tmCBqUkdUUe75k/sb8+4iPX1TdCZl3/zsb4r85nH9abp3YeMPqr+ATj
7TgaQsgIfcjoQtUGA9xAyJpO8GlbgYj8IOI+TAj9JQqoMwW3cJaCVrdbzBxf40tc
edIspNgIrjG6pioc5EtEa10WyhaC62eRILtf4T5nI9LAvw0GBJUpt5O/B/WvHHUO
TTXCXf/VSyalv5SRiDkgwqzf5yvbdFcUrVuI67PplIYZuVRoAAaGvTk12zR3W5Ue
lY9IYIxXtGy7B0xkVlOsg4wUeXDy+dKnJ8wRSEcHLQE9qkyoTHE0lB8kwhzQ7xaz
buDJU+OKX19BTjK9RjpW3itAxXPqYTCJ9EBmYM5AUZ47AqW+skQ46gIbUJpAJG9w
kV5HdQWLKlf88Fg19kAvBpcKs2C0m+TOUZtz80BYSvnEtVcf9ygWgbyprdHJjOhA
UabZX/zlBt1Y2qoHP/mfRLm8f6BEsgsJS9o57mFjb6CbW134t6EM4at43/x7j+a+
5bTo+cyCdSLnWL0EQAb4BYI9Lz7pnMacFsDTNwzIxOU2AU/lW6OTS9KyYPFZteDl
z9sTnG3Sv9LcFZdGHDrLZcRDcrdjWnRNPnILyXyhM2XywAizQWS+X/xPFXFrLfCe
I35jINOU9Q5LM+z/irQcenYvlaK2Gv9xPka7+3Plv/Gz/tKxgWjCe1ZlGRaxODvq
6agSwCSNeyKBKyT+j79Nz3+MFB/x4POCKPJc1vPX166dHUQZMMMOmXRu9AHa2HN/
UOBq8utnuxyzfIekQASkddIufXEfqI7H3mAtoZtdLaEdoo0dSDkSHxhNNupuOW9S
Z5xCJ/LFBbDY7pW2YysSfaQjcTuuu6WIDOtl7BcUavAh34E5Ht0/U3i0zD3/YHs1
O+B3vMcQvpteMdkh4yc3DM8Xqs7HlZh0lp3e9nXr++8DH0UCHvhw0PtTUALMjC1u
6PKZIULFJmuedA3ydRqPGd4T1OAmkh8l2i2tB+KsY7tunvwDZ3vi9OicQhwTskQv
HhvEPB8J9WmojquFrsnVrLJd29Z7EbmgfzA2QMhgjBwmKFoaBF4TwodeKeB5CI7b
9CxueBaRYeJ0XH8Clr7pQbO5fPn47fXx3tZNyPECWIN/Q4ARBx+A0cB3forKhMb6
8Gr/G3SXldUSzYKngfa7yOoAZ2yn0X8kdu8lQfw5Xxh7GACEaa2oMWaA92yvGtLC
QJrIFzENLQyFvIWtaSsA1IAGGfd1lfgp4dAf8fvxngYCkrrDC7vye3ZabFtZ+GjD
GZTuD6SluMrcr6h7tvkytCZR8tdEWubZgNrcyV7NyvqlbFDsfRMP0Fy2qLD8O5Nx
Yaw7yaEJA6a8PUzz/X4L3D6A5Lpwkf17p44bs/PQ9ILBWBMeexLFfhSvTdt+wRCf
y2qE/maI0gQ5QUWFc91lzfPq1sZYK/podzmACc5owjxuLfUHKecr325U3WXjI/y7
gH4bcr8VwKh+kybpdDBiuzpp3VKyZcno/vW+6kQ4Le4e1LW8pD5y83wjhwmYdx8d
4tsGGlSnWu+J3ABrbr6N2W6YtNM9x7MkWwPHv2c9m5UGjq6aNVEaMhUuMC55iVEP
4ROw4tNGByis8yB7kI6MusMiXwLPtvNkxki/5B4IriU8N0HicM7bZ6qplRAcIf9t
Cg7P2Gx76rvYd44YkXGtFNKQoOX1RkUGn8wE+t//lNggU9HW2QbjN0oc4MlWtIvq
96M1685W1TYoL8QvBFfMTAb2+6K+sWFhpuSfSQW/h509vNvoGdFLmVEryaUnzGBG
CNaxhuZx/OOPi9Fz09bnBZGLgH/8m72/i9+bL+uREAR/hZmPDZomv1VGKP/OH6fE
/rvU90WUgf9yhKoUYvk1uN1YnWeprA/WeGFFZRf/GgaSpI+CixH/cmTvJvr1cpab
0yiSObwyg8WLrRd+IpyC0xctE4eH9WXowGBuyoLDLwyK5g8uqjdVg6t6RhEPI3aU
o3PJq6gB0OSpWAtNpF4lPVNSCpA/MqLqXDr77e2wGf+DJbWhflU4azz2xRQx/XCr
CDbFvfZR7j3A6Q2a7LdLZwOMBlDy8f9yMmvr+Ms3CrpdAJte0z1OewzAdvkCbOyd
RJJl+XNU2y0UiRCtFyvoqdRKcRO892kEhxp55EGKCf1wK2pL0Z/kzc1LuShedsVa
+9EHB8a801Ox8Lnqw+YILXdmsgr6tvlrDl7WV5893oa37pbbCCI/oIc7D1ClaQCN
bp6O+uDjWKuWwU1AFDUiOzLlTE1i3hIzbHeX51tvU8XletNxX2PvTNCO7e5Rzs+u
OOv6LrV33njjLSoLufPkP47/tzp/asfvsmOMO2glBPV5KJX6wOH5v/S1NLKpi1fp
Im9KOGeZQD0ZgIcNWhJy1/JOJq6lJJQrRKIVkP0z/zsSuS+lR7e/uV7OLpRlX7Ot
OGijtyonds+eo8nkDRaGHFZdVhN3AJVQ921ntG2rla9TuOjD+JW0zI26iLkzJcHQ
SZnf9weBAdDvMeKBUZUy0lScR04EKEx+IilRaqJ33rpoekXVyI+jb3RiuRv4Kjge
2Lf9Lp1Wtj+ojxtZwW7OEkXi3pncm/et+kgQq4DJNGjOWTQ7CjV2tJMFZw2EMSON
UFXMyyXvzwehN72mAXrtt25PfoomNUptsX+lnmsV12LMig6YXpdJCARUyoLf+lpS
LXRFE9F5k/yARcED3ubkljLNxQTFBhGf+3hNTL7E1q623c9JfBoTc7mHE6Q+vZFE
qrS0qr1ECUgC5q0JSGNR5h24f6u8aopLfg2DNnLRFQ8mAJKqym3a+WNS9kbMFfOg
6i5fUnpvTEnnX6I5azVpB2biTkjZT4zzbfHE//RcedOsw9vtBEQjmEAzx6k42B++
H5xkW4Dlwzj+5V5MGtduQZqVhjQM6Iw7WsW/O3FtUx4r0u0Bq+sB/BnbiVyS9tGr
ZrmJ9DCynmNutiQFTz859bct1q2n01vTa1KoNuCTDcBTGk4jUtIUkqjUCAMPKCqX
QD0wdUyb99ztN2qhx/yFYeRKYLOf9YQyJMIB/ttOyuAukUcLrgNCrX7IaELWxycL
+5w2WgFqHphkk998RoJE9DTL5y7lWxVyfdlNNgt4GkNMtbuliFIuOjN02897AVC2
hoH4SulMtXRcXZI8G1C9OvHyMG1N1LSaAgdadMBqD3PIRDTJ8TAPAkz+zAAm3auZ
qk/eGMj+2deylRvW8fCn3xrfeO+o0TeRKfb/wpzDuiBww+ONTGnSBwfwGIpbDWhw
Yq4K7woRHiRwlT6MGneNKvMvrxEJ3Ev0V9b/KYbblxt5VZ+K7XZZU8dvdC2zyf0I
ip09nlzwYCms7a9tCMnu234yEXhPy6tvbxm4GHj/8IT7DWoOU/76oaiDZMmhkPTV
Ey7c9ZZoGxNOhNiaWQz/JtHaFw9dW+fG4SeltIlE8WFncr7T+aRPK5BjQWVFyKWb
5vVegzIq2IM3rpgIFC8z3OgDTq5DYMtMzNV2xFNCXDGwvJpjaHCjg8k5H5YYop3K
jmmxW2XSB2tqRVeYyuNJBZaucrh6xvxMgwodA+njQmJRov26+nPzj9g/J5jLWOJE
zCuyzsJzUPqPoSOY8kYiqixFq98YfTXYgUUwwpDcboDFvF2LBp2gZAjm6cvzU68C
pnf19naTTZuKW4r6kzMgbd6Q9mFuVc21SPuF9hosU+saY00Fwr6kCHwLG9DXwBSE
dacRdXiiJ6wxjR6s0e/jtP223ayYOqP4shvXpTV3nc7iiJNAZ4e3wxhVBPFfUrFk
SzlkDKpo8dnHNVgKQzUK2xQ8GbeDmG0BlF/T0SwsGrYmvyHhzrSUN5R+iyVZRHyc
WjnND+ZmpIhIZkGNhJQUisr09ZLQXh5AHRSz2DlKqaeFU2AQ9+Yaa7vY8XoJq5yZ
DZI2d7eJ6fJ8NN2CSFJjCIQZce+NsfKWMcQ4RjHeLVFtQgFPfkVqdHFLj6uxHVIa
aq107rVumwTI0/oZntB7tLOjYczQGK5CB/3WDAd7RWETIHICohxiX8HpSQvsTSPb
SePWiJ2PArCHlZwN+8/yxLftrTIDWA/2H3S9iC3a/Iq9kGaNoCuvflJIdPmfCPWN
0kyNaaGQjjes5erKbV+VaLTQhajwCwIuXdUnYC/bIcTvyxg5etZEq/Qt3yTJof+z
HBqzCsxe0/hBY1y0R2YECoTKEYu3RF0gW6FOzmrXBypCiMRE931goOuhJoT6Wb2s
w+3rAXiFU7bZCxij3o2CeWW2hACwGpWBi8UIGb1heWDoRDMqh4QPpOr4loc6gZG5
ILmYHbLryC39IwGSncxcQqiPFY3X60KKk5f2FPFXsQAvvpJuRytdU2bdikF+NLrX
XAAek3cMTpJOPpQYlYxn6/dmgBkG2A92uKh1AUstdRryIIeNLKtMpYUXwwNF1RNO
Bz6g3fRWYboYi0iO9j2Khe2Y4F1rGnuxdUE/ESGsQur/XnrtyPuWk0CKQjFlQGrp
8aOyVpT8Csr7j11QD8IqQxWyktB6WPfERIoJQfmTQkIoU/fO8TlQoE6ySR4rWcyN
qDk7ufLiBdZw5KmbH/ZSNlAe84Pf7Uf0NxdSbtrlnOrHePGlHL8pYl9LkeIPAmlo
3/jhTkBJfLT5y6uBlkDwVS9AqxMSAnDD2EFPp4Vxbm4iLDRdHrey8NV3bKPYSCRC
va/13aMPd+WmukJiEqSalfLN5g9WQFcDYWoOAqmRzVxjhhy51AwkgSZnbqxBjBWg
Z20ErQP4vCdPjZ/4VE9304jQF7wVx7kRVsCbS0FADdlM5gwiZ5Kt8wtiZthB5JpX
SlW1ik2RnrnP5SXuB37PfUqOnwXUZkLvOOh3eNnYFuzuYh3npSnuhcm9oY3Kj+yc
/9ygQ+dtlYs6miOfI4j3ircvdOtQJsePQBEag8HTDCSuLRLP0ZDGty+Pb1IQSXPi
ZnY+Y+MYilCKT+xG3ET/uCClIi4lsxfnzh5djcZW3W+tQFquM0iCzPuDy8pB47LR
9F0XCHti+EfzpLJCEQ3t08mdN6KeqgobExBoZzsLn9RbHKjlbhtrR13I7MxPMW2q
0U5h08Q0h3fZ0xMXeiGc2/EdnYlKvsi/hJPel4ayKDu6ZLwEs4h7MrC+O1bICPxt
pj83x7ecoaLpfRiz2wpbjDOrmz/UBqX4Cs7x0LCR1mo44kfh0AghPusAsqGPzzBp
Os+E6+10bsu/Ln0Md/43Vn7ZjMIJCokBjc9FCMqdJC/6RAxDZYW4BSDK+FTyiuiN
isyG34CB7rJ3qfb4SJTiJQSJu/9Yb3YD1ZgWj7zQaHftPe9O/j9K7i66K4AsVywM
juKUiMaKSVc/YHcCNWT8Flt/pMsdXvO91Y0WY5TsKdy8k4Cwb4n9kfxx+IZGjjiS
K/e1R8Gvn8RzUCL6vLy4FhARXKMa+Mv7In6TMzJ2AmpO9eEWaIjOHYYKonecdkxK
FpuCoBixDJmCnZzWuVL7AtI5It/VIPgyu2e2QZ2NUQPfMFsJ5Bxs9805FGnibvx4
GuI0yxvD6EAmlYjysqlDK6DgSar20No67Sf6+7c5HG618ir3f53S3f3YWylahLH5
GyeR2E9GfrsxlMLe0iU/koMWGDfKzx46ef8n8uMl2SXA0h8rlNdqXMSm8bz8L+ES
G3p/A5Lw/7omB4owAq7PjZ4ZdZyJLHVbfM21LLEaSaYyUG7LHuPuYIAysthe46xZ
wnRCaz8o1VGjslrnuuD3fvvKnySY9QeIIHgkztOET7wdV8fjGBw2T5Em5xeM3CC1
HnzfOfdfoBun63tPpacQvzbIjFEc//I9mS9ITxo6JN6xSeteSWAOldjWQRrW02BU
9hhnqu0O/fv8bVSK/mnSfQ0hxzMLWWWKJ0q+YinCgU6STZQuF0IK41X6afwX7eeG
ekgosFz+ALFL5tTXdCoIDNkILw1SoZ1MPTJZW5FODXwRIG/P5+mySeyxpg3egTiA
CkTgTFDVb+iQLAo9X9mh8Tc9WO242URXIsWtkPU2uX4BG3WlHhFTNwzcIVtxM8J+
ftNIIg4OqtDGSzM6R5yKLSTVnR73cP0xpamYkfk+KQXyBv1fwkN88foq2y6ZwANH
YvXKbUaWeee5FPBZF4zSJb8OvxamSDtnnKFY2BjS+wtJJjt5iu9GbnF/1KlYtPFB
xW7sSt9wA/+yFrDl5jM4aVeQW1Zz6rVKPUsU1TychAwI4A9zcmthHQ3Iu/Nsainn
VEoB2zUmUmsI5vx8hGcsXEpnVYLAiOaiYryJH4LaD2l4c7hapHoq65WEC4J1WFyD
KihmHLsTE0jm7FAxuSurV4OgWR4qTYUzo5aX489BukXWBJ38Hzj3+tnjg4bis9BI
8RoraflChZpwHqo8xIcA0N4k9e6jJHOjwImi0gRgqqPUqTMwi4jv1BsNLj3sIpVc
TB0T4XdngBSEEBJa6JaYY9mJetOrI8praEhJolxtn9Jk8rFl+pcAAtdVpcaOpVM5
Q6ZmuUD31uzLwuGxjM7ESKFpiqtJoSWuXIu8c0bfLLrj2gkqbDt+9vQ9lRNA4Mo2
T5nqqd5jyWITBb+DD+RS5K0mXEtsCjCNSa003ld99S/HIZaciOSSTr+8wNgfi6t2
ZNJfna6QZXBLIvu5fL2xJC5ElKNDZvgsNqeytb6jRmrWySrY6Iz9UvW7uVV7b2dL
sKNjGHH0Mst3Vist3J2KppV6sxIz9+/gqKycyTm4kn6H0hZ3nxftbGHPiXli8CNI
EHfoSggrjmcHmhWmXAyQaRZ8wvjtAIafMZmfy7pdUoEDVY8eo9MUzaH90PTgI8A3
f2jUuiDOoxp+b+NqBVYGtVALgZb5ZZg7Cxou3JNK1C57XH3z1ZOXRXhNlqH3oTsC
KMsXXo5NW+YgNiSEfxlUyakpG4e1hhiIzr4Ox/zYhMpZwxA1+yh+co8hv5wok0Ha
Flm4OYHnYmUrjAFr6VOQ/H0lMUl4TITmNwPghHjoypPYOpofSTNs/ER4B708kfoW
GXj8DkAawLFI8aSCfrMBp21mEbYGSFY2YH1MTlt5gaUMFfCSPs3SRcYQkWxacXig
CSJJU1tptSUopsqgZxu+GdBVF/X83EwaAsKCHUDcda08Xmhjeacl87zTP1Jw81N5
tbD/jTfPMAofBaqzVj5tlc8bJb/wVLmhl7+eDC4lmeIjhhVfVwClGWJM3nQZEs8t
VqIF336+V/te0OpgX+JQBuqH66wcQmi7ialBBJV4z/ZOPu4JBWIv4pQsex4hsAHv
JU9DPyuP0LJdW3wPr1m0oZnVkEz8Gxysr1uJQWy0PnOAJegZLjB55b08y3qHB3oz
w7TafKE+mY3UnC6F7AyxmrfrF2cv6Rh7OYRw0PF01tExi3c7WGuPceRCLr8joIL+
EIYUoFU7bN+BLBKOp77qdopApA3N6i0rI8I0E7MP2D+HJCjbOeiFem2Y2e7NRbiG
ZawQU7q9/POvAfoFBuyMKxFmx+eS6pQCIeB9O76jcOzoGYhx6EHAUH7MFIySlc3I
2g/Iv1bU0LctUHsk6Va/NlbDCiy48bVbUrYpLbTO6n5F65zD0QHtPcMj3bbvbZk6
ITOYOXC+03heMYx5WdJPZrxXpu0nSSLXPsXVbr0yfc4bmDI41+Nd0JIRrAuavCl/
RQuioWVVaizmHesCmhLkvmphKYKb8kSgB0nLXrEj96g346024QmhMT+z8evGTUVR
cB2Ou7czrpLn806rLJivvKQRgkuGPw1/CRyU3WeadJF4XxvlfdMsHLaVAv48RvMI
JiPsj2Y/OKX0VdWxPBIabYUviruIus/+D8jkHnmVwg1gAlPtJp7+brZj5HlkA14N
rElbRVKg+bkRRajyXtPDgH4jSYNjIEPxn77zCGRaM8kjE2kE5n4XI4Q4cIm+o0M0
0Zps9qaoNBjbvjgSbRYoSnW5r+B+xh+cBqJw4O+qzS6bmSTtU3vI8TLMcNXuU1sC
Rl4cSR1YagnC8q9jwb2kikkGyxhHy0HKzanuHg8LcqI++hn8d354R/BmA8YKRWKV
j76hghGzRc+ZAj8/kBUmnTy3aoqKSbeHLXPYubMim7Nji8818x6ueFW7o2gyaQ7t
MKYSMzvic4JCBRRVeUWij0e4SS+9tBA0Z+1pEieRD3a9lEF65Nh2Ze+xMvKl78dH
sTw+A6iUh/yKomH3v7fijqrS/Jrv++xRZLeL+LUNPYOjaFUy9Il6vMybuDJoo8UJ
XSsjZAUXRSkKuxUhkPN0fEt3yk49wJGs/v3ZRLGtIh4DR43mEJt6xWYpydoiTMZE
5z8EhwUH/FRznVJcdH7y+io6bs1VRE9DCJLEnmW7TVZtHg5unCtMKARoF1iNKRBQ
NFPJWI9eEx7jXu75AXEIfMSVa/AsavtGZHGF9VV8bgibPK5yntiCx9uH4eHwEhB1
6YWyZNs4OqUEMrZsRqd84Hg/bj9SOuitfp0Kp/iVSFz26UfkiZGLLko4WhWeogM+
ul+1weF5mNKHKvm4oroFGYb3SVRtpJdUjzvltMtZ5VwOBQIuW5hScBhdz2fTNZkB
riA8hLmdWE4AyD/b4a8jAX+f2vD4HAwzQhJdxErsVA54S8ZsykWhHA261oyxRtuY
g1Lv0hz4ZNM8rZ+SvnE/5I77Zqx3AjPie1I/fzK++LAcPcfxwzU8EFsx86uC/KMP
SHFaOst2lXumRbZr8x2DzF7BmxZN2Tf4MpvfnntuGxlrW5VYNxGj9hTcml6dhGqr
HrcstIADZ+d4D5McOvmkROPXBiS1RMsnq6RiRExrsVDYePz/IL8xQBWQcbER4dik
nAOJbfTFQoosgkN5aCgM/ewFVP6v4T+WMYOn4zP8yPZjzMOZUUQ5XMXwvW0kQona
QvIBGuR6oUc1PH2MHX3xa+mBL6Fig+FEek7laYfUQP8hA1nvE+Hr/619/EZKjPeM
SbCZbWutPYYQQSPISVY40pGosWxojwftflyZFysg6DieL6sPau7KXMosB+BJXGhJ
PXEpf4lEm/Wb2Dg5jql7RC/jHJN1+iXPSobg+4r7kW8vFpRRV5olG6iwtcRErrtz
PXs/hYPWdSVqZfubvA3AUffqhbCdtu3AYBpFTBZNBbFvYJ4wR8BFgN9hbf+5U6k/
x5BlB6JS/qSSwyzB4hSY06jLDKcH/G1JFLcC1uWJlBsQHiKnyYic33PBC1b3GSAa
4xs55Z5rCOzH0d3t74c6WkVWC6EjW1fSL0u8OOzIszbxkTNghEMNOzuLcbgyEami
SPs6Htvh26HBkCYMHg6Bga0UpmcYHI4333Mbjuu8eKaA8NdqAYM5M0Odr7d994DO
BirSpcWukkz4CwKi/kJdR4wARLevSUg4rQwZGiMgaM1MkLvKwk3zgnyEPEqwdiaH
Y3OTiEdvjvyFz+RI2Bgn6VFW6gAReiLZaZ8qjQD61zQCYukEJDTOnZEvg9wYZuir
K7qqpqD4zXQeEsPBJeU9Sh0dI6Yw3tiWul0jqmAKkXCq1JcAzo1SSqJHsGQzhiB3
f+x1abzqLf8Qz3PMrZyMODV8rpojIn6U/rY1kLeq0EWw/zDSZ31xvXoUI3zxezRl
7NEbBuenVTPwzL73MJTw6vzoEZ+QlucNdLIkwxNrQWBelvin5Ky4KZomvehDQboU
HU5EayNBKUK2NyWHrvVpkE9oUvkqwTMBT1ibgDuA0Cf5rS82AayeCmNcZOEOTL6X
pxdiHk7+n9i0R0+6xN2eBk1ZFqAjb3sLRssWxc/UhpbPYPqrZmWIyiREY/1As9xk
ID24fDBYPtsGVFFzOBZfhrx+sMOicijLuurS21pHtyaMD8WH/C5nrq6mU6ckHvW2
UKn+hGvo966jiQRZ+dewCCojNpn9vtNQ5e1qfsQqdUSVgToPON3NtFdy7FMYNHWB
nk+iDUI6gozCKrXLMl7wcxUa7QrIBJrvLoeD2bA13v1SsVeudEitCmwlfIo5j1EA
uEgkvht76z5AJyYf0O3UnRAFHtDPSzDtBDKALSwsRNuOiu1cJXYfO0I2ZBCaPswd
Hds77Zk9DCaiF1ocLO0GS0+TxLHJAaiZeFhBKTxTQWpnZclNJKU58Qqdzd//lvYm
zIbYO0n1rBF33i1Rct+ksP3fol2AahuUt19ZpdO1sqLG1vNB59RH/HHHlqN4BGot
cXhUORSj45ZWwSiVhyR90NVw/9J6R7/wdmiDPmrLcD1NT1ros7KbkrFyquWdyVqm
uewp+Qavj0f0M9sEjtEinWdTbiD2jSTiKYf5jbFJWNvMk2sdcVj0C+CM1nMuH3CS
1LQpbmgFjNZsL/437GkKVZivLtyAxCPGR3XBKBVYpAJ/b38VeMGhamJ4oNPW33h1
gpETEx3GVAoervXUJ7RqeeELDV6zMlN/8FXaFOx/pREDu2euxMqmdT1iI6JjFx3M
IYXlXercsuVNpepQFmnIZYmeQacxWSO++B8u6r3rQLs1qOBMFHYCXTdcUdtdX1PS
al1LfC+lt8p0VNB1TIaPnIUSdJfg/reIR3ZzDJaOemWk0Uym6zLMD46lDLzW7Tvv
VMS41mDiZNm92Rbi62r1ALka/QGmzea9hBOBs3/75UNJYe0vyYAdkGeBFkV6u7NI
GQLK5dphrCkqyYmDp0mEu9Jnf2O9c69KmF6Sa9wao2QIkVbllqWnaaXGs/UleZ8p
37uLmpzfMbW5eL16pwe+4/g2dK6j/SSylVr8q8/OPe+llq+DOr8DWvqKYWSYOwLe
kPfs8IUdRNj509oL0VHee6e1bGCy9ww9vwtIVQa2c9JNAgMEdakzDQ3N0CrM4q2h
psQVMqkbfsvi4SBlKymDS2yyDC6f7Sjkcsip6euReQry21gilBKWQ5iwfkYubupW
V4eS3ZNdHODnlVQSNGWstOwURr3ylwx1CV+9A2uE3f7CW+78YBsJgpMNg5C3l6QE
4KLS9egFPSMxJ1HtFYinLbMabPA7Oo3zZiB0oHr890KkvoH0NzGD1kWFGUGyJ0H3
fFR3RFu0GKyC5yXufnmySaYkP8H6pifLqggRIHpgIWOmGvMnYvOzt/f72gNJyGa4
f+GbtlPQYxCPsKOeNjR6S2h1DOhWzMfE/HmwDSjc04uhSD185RC8nOoBOnG3wShQ
8Tg61vmGF1/fnb9hOENf702VEHYU3/EVXR95/AP2GoxE61SZAWPmiemLhJ6n/krM
1Yz9/QEnE0ldKtvZEXy9ETYPYA543seBgVyYsiYpvdGCintD+LrGggy1LZ31b00t
6uW2R9XGZKb586kw4SpGQgdoELzS5ecAqHm5D31DNGO9Aqn3jFlhWSTsi+I17vDu
DxLhUOgx6RY8RUqTnZGoUT6k+A2mtHTz9mOvR+9F6Gix+uWLcJu2cF+Zl6s73MR2
JjjGZNFnSP3qDJPwx/am8JQKnyf4EGPOmq06HQgN7zRJEf1o/IyzJlgzdnbi9ewm
/Ak9ScutmuQ3J2yV0UMMjtqfi0czzOm08iExsyCwC6KkmAWzUCVIMDBCO3/PRC3b
eXAO0ZKQq0Jpq8Ypx8f0KMV0EPfhfrqUmVtgpfiVCRNHzghp6ttLVgVB+2fC44LK
bc/QQIKv76nsJOA2dxwPxVt0jiq9m/qIGgU/cEbMEoHzCVtaIOVUptt9GqBc1fIM
fo+3kVI1TNYJIPbtxtfhav7AcFJM8pnXAYGiAQ1PZ5aCsxQLzDlsRolj8o16HxIA
Bam0MG8rbBzclLwDebR/rDshVxG6ClcgSdmYkR44qZ03UYo0TgBdCOK5fjnV8L8A
dSDMS5B7kqpiz33NNkOqhpwpg1G6aPQl03V67415nu7ZUqM13CU1JuwDUSwdhaiC
/mcnwjAtVMaLOGoQW/7oJ4PJPugNP3ZgwmFJuzbzYHJO/GnuNMjfXvWt02JLxtN+
wYfIOIgrpj/1j4gCJDxXHXSyRY7fdbGB/PRwwwl+g8giJcpq4ESZ6WJU4RmuDMVQ
hinx/Ze/1uoKLi8dXTRylxcwwKiOgW8jMHIZlBjdDpvPnV/Vn9RoONRMYgogWpEC
aSoMoCjtsGvI7BdHA3eb8B7OA1S5dx3sXIRQ7AJek1zvFy132lEMSe5KeV8f16wz
GCvLbJ1FkaEJoFAKAQh4T2mR5O4X/6oNOe9+zVyScwXYZMPQbBm88rp8DFhisc1m
w6nmR1IoGkAJPoy2PNtjXqc5bX/M++r/7EMtO3JJs9ScBFvuhtdL06T+jYMcCgyj
cPr1HAR1mRho2jn0zsJOEVFUhmdcBm1pv/A+3D9MgnWKmn8k6AcMiZF4zXQ7i/mk
t1zSyBHI4DkEAfnuSk5L+u0UeUX+K4RVlII8q5dF+M8QQB5SANiDVt9M+ymh4Pta
DooEJ3npuQWQs6WyzJdUKCB0Qgeo5cJovfk4VKwcRa013Tcw4k0kxQM6FNOXyvf8
v2QeSIYHXmwbeKsjnxO6swHTzbLt7tYbXyo0CI5nqvzeLM7ipSNY4mwckaQkrM5i
gBLP9MBIC/Hnp3nTehN5aJ54VZmu5MqEeJ8jamD0yxnO2yjsiKLmLby6DL63Rjgt
/TNB9yTawjHGRsMkuc92uiy7X/bbZoy32QYkPAuRTK3FsUpJcZGqvRBJDEqfGWa3
kNh2sybQAH+SsA4Ic8B0xr0BKGJefbK40qwKWqEedLm+h/pagw1gv5NDVuvTUggA
SXExZh/84QaDSMxd1JKb4xWOmKpN19lq4HVq1QPvQi/xNi3ct4eqJOuEHKClr4af
cflGlDGoB/tjvo3veFp6GEUkPz87SZh/lVdkrlGNBuq3Ui7wZx7R4WYD8audBqIu
ay1ZeCxRzzg6qmE5pOloMtpy3mZViP+CahU3nFXLXlVIi8K+3QftKHYOtYrh584q
NuF8R6gQ1tRu1LDldLyhrKy1kjJOWj/TQGZdBuZQQQtEwfhVALaPJ656BlJk8A4e
46U088Cr59yv/mO0JdnBNETln6ik4d/X2RfWNFyt+33zDHirjP2Fjtl3B6M70qC9
L41cOAM4T+ZVJkKXl+wOd5BU7WW/2AOj+YxaTvLAXUlI+H8cSxJ1zfsNntxJSblR
JUQ+iSBBrUrmoVqjE8qJ6d9Pz8LoduT5SJI5r9dfgHh95w88RuHGKLRTts2FQoFI
sRmFm9n2XOM4SpnbDaQDBLFC7SN5jke+P1IPhEkveoeF9JEU6HD3gRv0Z8Yt/skI
Hyyb5xgUfN6gT/GSO2KopDC3l/eEnMSqK4xExuT7Mmuy0LuZdy99flg2WP7JuGYR
`protect END_PROTECTED
