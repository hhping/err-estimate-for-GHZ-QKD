`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bmtg/OojXMovmbXSTFAiTIAvQkQB/31BGBTHJh/TZeSn+2fSyR6XExMMSHb8onhh
tlm3c5nVBghKvkjpsFIIk2ywE0X4tdfPGbPix2vXjJfM3k9n3IhhrLKywrhFKwXm
+IHkBuwD/usEUfh1H4n863KdPVdBRBc9pyUeuFBX4nJSBSoiEJLqJGS7o+mH1LK9
IRws8SNj3g4t0ZKvJDBYlNS8FQcej6GiFCZI+51zSRGeH0lMRWYG6D8Ixqbc/qzR
OU5VemsCkfdfCkEhzcZFzVkePXOP+EV0zP5Eu9t/z1XMV2/fz6Ij/M8f2Tlqa6td
FKvIOZleT7oHLndHmtKDGDcJrhubxUy/fpHd/q213QD93MIY2wruBHt06xPMYgn2
voa4Wigjrv0j+w2gj4DGBKX6aoSANyvp0439+XdS9fAyGFpcZmAxgUdIU/Zb5XSx
NOI4gvI/w6RNV2YHHMtWbPffIB+Xbfh5fkqaE7tWjLoJkpbGJoCoVbe+opQZ21C+
9OU6mR2AdbaYJTRkjb8MQ07BWnYhu6Lq6w2enllyHMIhca6R+czzPSFUucnuJXGz
0Gha5Itooa1vszODq2dIB7mNrUYTzS5Hk5UdhqmwtUSnPebEP0G4q7YnlM518+xV
UKqsJ2vV1yhvAzRteNRa1SGj6ASdoPShb9h81WgU0PYw3Kbzo6L2ZIWvKA1dWK9v
Dr3s6bBuGdSba6eXTXXKBLYx+1dhYaDEe2499IbP79Cbl5TGtJIa/JhgfRNEiL5G
WHW+KYrRL+HWdZHg4q7OrMImLli3oWRsZb1o/+Dq/reZ6ybijokiJJ5QJGVCBixX
Uonh//8CvCrSobQdO64zNvjiOfv7vFCDxiyDmRKsbiRzN2eS7zyYq0s9WtiGMY0+
hd9pLdH3HQICXXnNCkL4PrbxMWDXrFkz3XzaPByzU9l7/F4gJ8xPDNRDHxa9XW0z
j5MAjc+reAjKhRaKW7fRW20OaQamZOldpxI6oLmqJT3ZT3iyEGuKB7PNyAvpR+9T
ShxPnfWc9Q2xDgv/i7XeJUFWNwC7kM9QrK5Z11lqpsM8F3Nq++y1vBbrZNqN7LlF
FQaifKP+OjE9lDN2na1N0BuuYc8MKVdV0ZMpxK+D74SUiUO5o0q1z+DlUz9Umusw
a/YpOJTo9Z9cj+ICt1WD/WZNqpBAqHVPupQCIVrzu45E9rJ68KrSB0/FcSNxK3BY
z9lUgjkFVEbyUmrQ6tjfklXsluTFkkIsHDbBNYTjZ4PWI8jRh1EBVTFLhQdwS12p
x4Un3Bo3UHXKzJiCUMMYyS7rR1/hMTB41XaHHpvoQOUN7BNzPls2fcCrKpWohsI2
EG/C2CAFJwD/Ho7pBY/eFgWOn+vTcIl7EqLFsj8rNAYZfsayyu6vPB00LJ1fJ3mS
Gud2wihXQBGwOhK1THdJ5uEgeYR7TkQYgs6UluDnqBH7sDdzaZzeiiL2hQrulV2g
S/r/cm0jnmM/Q4fQmOisD8EgSAfywZWfihhwO+RDzToVaYb+0W5cFeVNVrM52qnY
VDnAkEl4+tYrkHLf9Y/xuETy/Gy13EcY8gIrQYoM9NEARgM4uqgjPR3PbK4tNTPY
IKqm9F+8exYggdTIoe8YVtEUVfmwK2M50+efR3r1sFwaGs66KQGKqXofFfRgnbFx
CdyiwTrkvWQUUrtiNx3zkaOEPQnaSycvNZV1u7NwychCwJJbQQ8l/WDtHMKsSkCM
nP05GmfaXjjL4cgvbNH07lv0RSvVuy2G20smyIKJK/TmgYaBVZEVP0MKCRP5Rf7o
u0QSajPIP+eVu8W4F4P+sNjO7cXcIXu+u76TsgSArR7CNSBskMf5Q8HFK+P47CoA
JbNhI6mhFqEKnc1XisRF78/IHWKxx0JrKyVkwpZKyk+Ro65f+zvD2dobmtVeKR7D
Md1dd3483fLS8btjo4Jls720sW0OkmQmAMxd/fd7P1mmNzhhnAInA4jGhW3BRuux
bs4Lhm9GsHjWwQg2fVJvS4xlg4Vc1n/CH6qo1gBDMRsz0Oj1LHFmSSR3zYfJnDMb
bow8xvQja47iDWUxQsakzN1vnKPDbjMcaOqcSQLCeLa1qbGbVbK4NZUe4n0veCRZ
l/lCUa7ALpv9ThcLF5gwh5tYiatM5+mOMgeEpFKBLtOPuxJGqijW8JlNmq2bdw/M
2lcmd4b9wpoGlM97w71ZLzGxF3HmIARO8s6Hc9nnulwXhyb3rsFdPE2MhsaLxRe+
2BKgb+KvlsM8NhhP1IL/oZ1LV2yD6RIt26nBnUUQgudqGfZZGZEMn2jZygEitetb
BaqutKjmVwivaMfShfkike5Ce131L/7rkcrXg2kJXSbGgmAsiYtS/E+OLED65BtA
R4IQz+7mhHu2/pWhdFjh7g==
`protect END_PROTECTED
