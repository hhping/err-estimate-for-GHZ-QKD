`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+o7KrH4Kwwe98Cx5bxwCKxtNM7E8p8rOZ8oH/YlwILb+YI1tdLbukBGvODy1/Gq
+6WBTlb9T2A8gX7wXBb9heD6V0V7oNSTq4dnu7+OpfY1/gJQ3NqR89jO3/ceisaV
KNaLSSL6VNj8AVHRGRXCl0apz1RpM3IAq4MUgSVkjHKwrnvzUiR5hrZf2Bc3xeFr
TWHDsf88j0zrQFRXX7d4WebmFDxGgt+kAFPpNUREe8rGWHmd06fADjLBxtIwBXr4
c4Vcud0A3IoTIK34s/iquU+EVELy3HntJJXRP4N4VNKwTdAZqqgpaMTALwqJsyf5
+Z3Px776JLu+DgjDNujTK9gIjIc2coxyMM5E0NgQELzhRinXpZQ2X7gCsbh85qGb
5CT58UCJPuWmvYAnn7lOAIB5LCR3MIGgdZCe1nB56FUknbocBiAANLe9+5dmHmbp
VXqk67ECEC8S5EmDRlie574adTsZVKfvUWWszwC3GXcDrojLduf9JuXwBNXhs7te
0PkiVPppCX2Zth7nNQn8VEbFmFXBh1fWVtp8qqnbdGXhvruwo6va6/yTEkBpe5bm
lLzR5t7PoCrlb97SnJS4RAcJuhQQQE8XaF7SShHO4VNoGREOJTThS7+KcfGA7vAf
1f76D68A/6F1zu9d9gQLQA==
`protect END_PROTECTED
