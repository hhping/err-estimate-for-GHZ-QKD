`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79Rky4b+1QrcLgRJ+7lA0YNPgINPPKfcZQjPB0jbtd69q3htDWnRC0aOd3mJsuRi
lqsRkihW1/X+gEluohY9swQy349AWFMpsHJksG/kmN03udyOIjmmUvj93RkQ4ufI
WnKGMZPSHacu7XYCv3OVtjeWDdQNWdXY3r8snyyWmnKK62GTi7a3j4LJewIZoHCY
5XaDQ21z7CUew1RqlbVpJMMjbgfeSS2tpz8H2BHId+sm0iqTG09wmXLiGx5TUsOc
JVw8y8TOZcxVThvOnxBPh50MsigLepV8bjCaOUMvUh2nsxCkqNFsi/NEW2BWPgEj
dUVqDYDFdgArGY1NvlC4WT3Z40WP7YgBOI2J67XYIPL8wYhuswqq9SkkBtIMoqRd
`protect END_PROTECTED
