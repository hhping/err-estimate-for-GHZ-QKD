`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RvMpEDQ3Yk8s2g0HIqQay4h0n5swoqMoDKvi9G9P4GSH2VwdzuzinOu95KqdOzSb
V3st9tH9Z6IOsek0kuGKyudY1bZls7t0XZl9v5ZvB4bJigCogJvO/gGx5ptd7key
qnV5XheYDPTH+ld1z/atZsqg1HmsrgYJy/fYxiYFaV9DPnoidAyxB4z6bqeDsTLA
72CjGaPdghk7T0OCIIrXon5PXAp+9QkiicDTzxScINfQB1knqyCRq24u8Bvp3dtb
VOUpUCyQermQIJ26Tx1/kZ7iisroI2VsWQTNuB8H/EawgjUfMem+I128T0juOLqU
75z7u/VygIot4e1alOfGKFwc3X7QEs0cjIKy8a3DlqeQw3irbPXaDIsl5uGKS+La
eLK5vKAt39mJu6fGS+OBIvgr9HjEdjoygIqNitpw14B1nvnOufHiszYA9EfSohTi
iRL8J/jeoMlMCUAUoDFKAnOWp4FyYp9a5d3AzP+aM07X/7PCP6hdYxNljxdkazTf
i5DyhnSB1V4NQ89NnRewA7l/L3ByiPJwSJtqdG4HWApw5LSBnWeaGi0XK4u41MdG
S6ULcFc8/zx6d1MH+XMLBg==
`protect END_PROTECTED
