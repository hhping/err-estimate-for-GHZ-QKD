`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVfLBM6ophNGgg2GnckJGVAPTl/0gsi7O9gAKLZCyCczIaPpaqWjkY4mp2xdeieO
PXLplI8qG69WdkJJO+Qk/ow29gfUGRKVtqlrSVtRJwhUKIbJ9To+buagUW98Oer5
1zJHeQM+SbRNXhefDvl2gEzD79HJBz7oR/HvyAQBwrM9NY07zYBfhbrKg8U9KShU
MKONJSsSIyTTTzTG7uyTWlgFKaQ4+BtLdFcILhJP9m1vTtBLsu9oiiv0FojMgJ9l
4Esc8eR1KDF9eedm0iWZ/Mk5n9/0agcLGvKl31BmH8jiSxuRZR22EDoeH+44aJjw
9jqd14LjPz+lkbo3NgOkvhcTU6uHdyg99P8u1y5+vWhqbCATj8qqKkK3OSEYmSeY
VcnyF5iOP4aoycdBHjCtMLxbRI4C2Q4ir8362WuluiWtSmLBFsxHJDhRQ9DFK9kr
o/eG0nzluwIvQ0eUDsVMYYRMRp9PxAcwSQiOby7NlrizV+QWHx98RsoyZh4nhSYR
emfWeMtK1z5uTDNkoIiwt53HQqYyNN3OUA1+xfO7Ww0tkM3Dn4RNtGqOxxTwTem2
KBUnOKl6XT1USsimb5i28mc2Nnsl+f8/Pxywva62wjHTacX2pBzkTmV9OfcWfZgg
cqNNLiNKhUZLlB9PrYizme8rhT04LLGaVrskT+MfxdU6KAqOu4B2Goii9+FIZVIw
WZPyZupPSCagC5NgTwIgx4Gv0MR9o+WkGwKrDXT/zEkxB59khH19vgQCsTgsxaAJ
E39ciHrneNa+gN+7tuUlI/+q3titZ9aLHpkDrKHnsmWvrt6C6lSv++5IJcri7o/u
hjQxshhZrAYXSQfk2PUfHIT+5/llaXfyhiEjOhIEfBGS/coJ3gKtzXoHoR9axusl
Vgs0DmEVqt4LPa5cIU5t3fZkggiLz+hJb5jLvXo9uMRcYbXWeigVf6YpmUStaEk9
VVsrxTCeV8wlcx2lEf7cME8OOk0BxCwlusUqh/++IkjV1wihzKgVorVZgfOitjIJ
5csP/aVxrq8cfOZtNZZoWxLTvPqzIX/ZwG3kkcTtKRyaeQ5d1knS0B04L1lqRvz7
NLk+agXH3GCAXeidc7egY37cTVSQS+zBxkKQh/UJ2XJVbxsopE06g1Ft5mhDEsdH
opih4Qc01JPgO3dAim/QWDXXADOQpM1DnUcgZk90fgP1z5oUrq7S00CUEdCBaRcP
2lqZRs1VahkAuqNuWDvA1vKwKNXZgm05r3h64p05rgkaqPZnrYdTfIwCejlO3uNC
glSsu9lZSFdWRguQ9Uh6SzExza2z9z3QAWDxQ8kedk/rw6WyP7ox6XWl2TnNu4cI
GxZvoi95d9+ilcvhpDGp5bFPbU7hd+11lqU+bwIKSX5EsPDa/5ML7qypDwu6WsdE
Y3RSPpyleJAnJ3plbxuNrSPv9THEc6eLaqNcUArStutMArmK42T9ESvwBCDROAIW
P0+aZ2Jm4k0OYYoP2qcvfm3OUvVOaUNTN3N1asVlbLWF2CGYULCxmubLpmVs3tYO
BQPKNjEkWdaAS6rOXotcWOi/gUg/vgsz7ytEv6Y4C+YHLqlFBeZamkLadgXbgiyY
az7Putvl3pxUEPHYJnsyDRd2Nf+TJkv+m/zFw9mDISn3UDGtXX9QK1Yp9cMRrO91
Kv8b9FlY2FuEfTrZo9H+DpGAR8FqP406eQD8KRXkeSzva182zFRED5J4p7zypyxF
oRbFKrs49oxs3PFGHOcqy8LB4c45Y3Io9/cJYYMvXWAdoir7BNoE+UUYk3HwSpup
teCnnyC8JfOguuKWQdtkGlmOYMjE4dz1Pg6ry7yd/UQyvl+bSSOW/+BbdMqWQhLw
X+RuezZm/4Ct/IUtcBFwAhhaQKxFtxYgxzTsf5Ea0f0ePBN8IHB2jSQB/dsGMnmn
9stLBh9p7esPGc6DCI3fgcMOQtjmDtOjsKxZ9QvWGC3vBFCauMxbCx1oGtFTDnls
vPxputrFOdTfjFdxzK1S9a5jOFhAB0+hRL0rttyVqyPVc6d+YADmpTn511Sl8iFa
OOSJ4JwXTeBrvRErldcJcr5ihnSdQrwukiY1K1p5+GFA6b60q+tmCZARPa1KUkJb
4XOrWRAXSHDbUNKdll2VpTHHNut6xrcVDQUqp8TukrDOP5o289ZbwFdOknPPWS1X
LwoaT3C6kimkNiDrRWjR6JO+BJ6PMZKDV5YJvrkptl9fNYmsE44dESIJxcAVsTra
iNNH0QjxpToaf11ZXp719cmdCqOIyR2Uzb0iIicywspJNOyP6EFy3Yx/yWhGpByN
XYKUb9wpXwHtDJsUx5mOYAbTJ7Sdl1M89n5b/M4oUVHrhgc8s0UF981zEtIDEg+c
bEpFgVDsduTye9kLwR2I8f8EfMyBKNE45LTonmpuGTribB2mDL52D1YLy2INxoQc
2pww3G6u981obhmuzsEjnTtZcjpEXE+Vs0iR0MgWeOd85NcBIInlQa6zDx0QsxY1
9J99NvHo1dGeK6vkIdlPRR37EPRcH02WHT2iaK1sp5jK2myw97F5rx6JsFEaEOwW
m9hiZJAwHgCb80qs8k9SvE36je+Ggty1M+sxrxJns0qCsQIKUf/9I20ufliQxTYs
X1gtm6wCWmZZMEn1DFMcxstR+T6bU1FVsDgMgPQAqOEzpCPQJdDWcC1+Flpjgnh3
r3s+x9WNsGvgRkYc+i6NhwvCcEFubikNBPRG2vVIBL4Ccf/BqFUPg57zD7HUUKtr
S4kHt/99eZM2/+xI6rVSoKKYDca8+PBI/s9UDrVMH6BfqS3LbAGXnvXG9WbrGn8V
BiZ4BoH2ZOUOEJqM/YeFDXhZfkgtDxXzStu7i8/Umzi7mFlQokWoOX7YjxnVQlxY
Vc7uyBXOxocDvm0GeZBq/KFTYETEuTwj3IgdqdGkVMLrjNTOSJTrkIRQBewXnUin
/MSsClmjD1ioy09lhmldxQaCcc03vw8Qa1Up8vIiNe4FRKHyuDQ643RO6H/MWCuC
U6FtcEfQJVtuF22DlgFWLEBdDMHeYkp1IJ1/IzHP2Fen0XRDRfPOf7vdInbHwfOj
PYp0cKsz+RI+mWNzQfr28YOCxp2BGDr5xlPM5y8N72zxBqVuERp+wI/IBL2KvgOU
ojqZgDzBu4sauHQE6GT9l/dpqHNaPwcuHVAVwSbZKmPtsD9PKA0dveEtK0B97IQI
PQkPKbqS/y5U3bK6gIw8LYPmAI831+0L/K+0UnA6QXjW77UlNiOl8O7ngcwqMzZ2
nwlkiWDZpHANnQCD8s1cV4W9KByq27jn88/JDy2A4kWBhWdjANYCYBDAfXIPWiGt
UMCqLO+aZ489luxC2qcS1Ag5WM+wBPiuUpQinuouO96UvZlcpLnS6E+EUbGZndgz
TXnjLYbnOa0h6wi6Fjv3522xgR9bmlLz2Yp8lHOXoyM7MYTJMOoZyRshQOMUh3Qg
dMBHn0kCaGBUR2CsydDWDs1IeFUmbi0XLxor6WmB1qqDO5YzTLPdR+vaTfamUzAh
M+oNnby/j5kqBFV49VKaA2RLIZ6bpy0LAXkT8cjG2lhxf0zuLY8avSQnYT3n87Zh
a+lY6+d3B/9EXLbpEnon5ksO9M62CtjWFs674fSCWQJvn8B3H9k4t2BI86iha+/f
8J1WqWUYwocaAk+Jywy/hWWWwtO5ioFSSaPV6P0gX6C5a1jIIswwX96B2vXiNrTu
VwfbQ3VJhqlpS8SxuFkzUb48UPOoNkFMc9sw6LBXqCR2gmWic3fWUwcjIbcQh2rG
NfgC4ZjZ6w5A53SqWlKNmVWbPXOpV1kB/6MdW9o59F/VV2pQUs8YjsZstHgBkoN3
+mbgV05rJgOE4D1rIrMwbZhJdSRR3dJ2ZKUn6MevUWo63BFfUvcvkprasAheTPfW
rrsO+w4PHvM+vYDMH0iAhy96182GRKgiXXaT8qqNsXShMZMnlxVjt9ZgGsVpghf0
kEv+1QFgrSb8JrdRl+IhR0yFRXsevYrJCkgGodZ4v81nix2+aaiYLWerJXUpiTQD
o2o2gav4V1iXp9h9zuSJvrXZAQht9TvhVRdI+2N04VPPPsTD3NjUqspJnMzXfyXJ
0Qurq4NO+/1Z6EXSAm68chI5z3KdNSbXoGXA/8y12ksGGXxTfmIGnDD5YaZ3Frj5
Mscclx1N0kUcZaY/gZrYT0kbp6NtPu2GKGYU9LjKP0f4G1P0zANbCc0HT2EilrhC
68rHo7anUijzxvx5bXEUZmxyfaFLmbXCLdUtThWw/GAoCKNICFIfRgZKrn5Ffnx8
kqeaMqrJBZQo10im+g5roNWeMlBc0R3HKXe3q2N/L1idmyPfPZNngOfQnOzYZmau
CnZ1/+5SnjFSWkOZ9ynJHyFLVYfgOboQrWg8EPt/GF/nRnDPAetXzjLADNLZY8Yz
ZK6fnjRtiPtZhJTP7SecFnAxVHhx25SbjoQQ8qrOaIEych+u0PIR6utgpzaXG3wL
hdbzwbUPaWz0r3VNCoFgDTLDi7mGVl/l6kVM1bv2wwO3+Z8bUfvZ5yeraRlh5Fek
jnAjSd6qOkXnzcdg1T8U8cSsM3azcurVsoqDErMbLaidrD63HV4zRahBBfN5KMbV
lPQsJZnymkFdORkDam/rrfr3EDmB58217XUT+U72rl1fVSEy2xuFN167yo6yTSOE
lFEFftLnpk8pUEDjDMF5vcrifSQrnYIexD8O3u8Z3BM4E+H9r76qtCJ71uhkaCmo
/fpvE+NegJLCfvwSCdfy3Zz18x9/oz3wFTGz7QNfFGlBnP86voF4jXkBpbKEwwif
y1e2gAgfMI2h3y+Kjm90JbQelMcUreZ60sKmfmOCxDNRtAlw70F6tu2ZpUvledlA
9K86ZjTkY7c3HMY5gf2dCu34F6YZz5nB6M+JoWeo+EIe2okJlrhDFrg9m4/+NzvO
yTuPbf4+x4v3cig0Wsdyu/aIREo2SWWq00dlFKsOFW8ttGut5Y2xBKKfXkpKEEzr
uGi/VTVa4EVfxk12XWrsjsHp+gjp2A2s3Z+U4kAXPuVPuZjNsm/ZgEQFOapj2iVJ
A93amdwnBEirh3HML5Q9dH0eyOY3fvdhfmjmpZ2YBjfl8Qk5pq8YWdOrolgEj97d
6/BCJeVXr4Jg8WSBn3ydSPudcigiecrvgSlbjeDXlIF0HLk14KjWx0zw8+NBv+IH
usB+5P4Q6jK/nUvRqkcp2IdhqUttJkkQoS/H2QMlTUst8M2bg6lctorn8WORToWO
nXRpiyJNbK7d6wgTNqhIniwSCQIaeBQNnR4GZacymG2Cd73C+qphqFEvl4ZzkAAb
gDGjm507sery2fBicr4NrYL6XXDkcm97bw98Y8mXZcCeiqwJjrJNewCq36idVRxu
qSjbtjm6Y4xW5jbu5UJmtWW//6G8p75Z1q54zLpZx7LwtPYUMSKmZqK0lQyNQSEg
x5it95nYFwhLIpGQ1Y/WS9ecnSIsmJZ60fDnn161fwhnvXc9BMI/STjRmptw/mM4
RPhKPZ6qWxu/0TPzd74QVYx/dSYOSq2/BfXdvIMfdL9+u7Xf/sDHi108Jvd604Nn
oRS6S9qMDUYuY3fUeRUuhH+lgCIdPD9xL5xS/xM3KP+8bJexBYsTVcxGVQ/6mgHM
7yxE3bMX803NSp9TMd32kST9QTdauFKzd4I7Q0cPM0A/Md9oSa7QQZqcY5kuylb0
K6oSSKcRyODsKDsnTxXT7luhO9XyhXTRzYak1mL9+JTxlOcYmxPYriptGP0XMUJI
VULZTv2G3KbxhHawvqhTSy1maPU8dufjuegBTg3XyHIETuJsBkzumP/RnRGwZJl8
ZEzENMxy0egMqxVDx+Jef5Tco9W5CrnsspGbXNAGk6GhNZ3clmUUFYsu7E2nA+hP
lxGwbPZ/72WMVFmOq3EHXt2YrBaZ9UD9mur3925XEbrCHQCwIYqkW/qLKikEz42U
YlBucqOcZj/XZiz/WkFBCZDvdY7ML0aOHtwnY45OhAdcKIeL88Rvph3M6gLC3/g4
IK3bBKP8KhWwcihOCaWF5vXr/rDrimbN3Ksypg7+oSbve65BVMpB+CcvxHF9xSvp
fDrU4iXKtKOuOZ/sJLYM9kxISrtSFF7oZNfY0Vn7K5a2BCnD6vBlLbs54BtpIKbY
l2JEnaMAuiyTcKM/51WGqxZ5k6RgIVMDtPXSs6X16vIOJbPvqB461ERgmuyGK5TP
TLVDYKfEkvSh0MotkCDixbkqsnJa3NutiOfmTT3ua8taa/9P29Yy4A23k2nz3AqL
FKxpXXrerpMwWkEZSswptyKWNhK9OIZo6nhroyKNn9/e+dw8W56Ps43Ffl9vt4zw
TGQBgZupnq+GbktePIL3RjRnoKpil+Icvw48vxAPlUx5P0xGWfMuSPMceeJtyudw
eBu+zltF8yfNKE9PYLeeFIKOvtfrVocDzpX85K8Hh9vgibrxwBvGA4/8R87R9Xez
s0UaFgt6o7bzXvMGLg3S9jBVJyhNTuyCHDLFH8f++Oif99YtI0+ByLzTrEYWrn4B
5GEGr2A+hKkybutIxhLIqvEYcP0NPX0vcvMQskTLvGmhUVBQBvE0R3ID8wJnYuO9
YJ7kUFPI5/dXyCoqPg+2uJk9TbrpMa650zqZaatJMAWmN7uZVbVuBzQzn/d3sa6Z
abW9bT/95KMm4u5JXjv5kdkN5Og2qJa8CDX5YoNyLR6CUX/m9ZbDQcs6dBjglZo4
Qu3Rrx07XgRyetIFyytLSMIflTmOLve5huW+McNxvkfbP7aVLxyuH/eIC+PXx2FX
B2J+4W+jkaiW3D6gj8cBnB4bgx73JfwIycPaLGUgIokAEYMJAnTnFqhMO6L9ycHt
WwnnXcrDsxD+EIGav4oP3w3seL1Hlo8ACTM9tC1cPFm6mJMOUzBI1LtGJii6+h1/
OA/KUDAC/XZhvC6O8koVqfitUkGM1hln33319ROZuREgqPsQvA0m7SbpPmAWiHBZ
OP7Z0YrawkSj7K7i/Z/RfJhwCP8/gi1wSO9obC3Mn0OuS6wtcOrmlKfHt3hR9jO4
W0yqSYM35MFJhFCdcAan4stcxnwWxmbpBOoZmOtvORcGEd66w3rTxge6jXZAKATs
5NQNot5YLEbpwfIUAV7bMMGBR9VSZ+ExtgJNYD/vYwz6m6McnvjnOTzjb3+/2kVO
e5vP3DIfRDF7/3CI7eGPiwex6Phj31OUR8JIq2PLAmMvnu371916mAWnJbYr+gaS
qid4PuUx//E4vKulfcNDosipRH7cKN/JOqaSCjrFwrE/wXDcmnDzUZskYW5hYlmv
jUnoLUKefgX27dYb6ffNfuHEpnLFceBdh4t3cqCRC9fUXw5LXfl+wzrUbfgQAYzj
+90/QTHyqZ53VFq1GtqPGj7fJ6mQJMP2RU4sDVRKcZOzzprMV3GH7UxZdO1SJJsW
PqU9JGWF7fB46W3SxY2eRvsB8jOz36mstFOqj2qPFN7TwFTfqRK7AfJ4t5Eduoxv
zjSx1fg7pLDrPJLUK7brOgXCkHaEzKeFfEB3oMAwJHcASpTB1U8bzK5Mzg0lZ2n8
T+wdrvme8eIAQAk6TXRdjc3LFD5SC3CPg5iRBN3vQyZ89BhvrwdCEVrGA/qUVVUP
OoeLgH0thhIW0JDHuehZ4Y0j0Ra30yYG/tN4cJ+j6w8dsUko5owTIdeXSvGRn4YL
i0dt97eLgfMBn+lGuH8wEyJLpYaP5Md+HwGHVjTVbutMpqDl7axxGyD3I+Nvz4PI
UuVct8sPv1ntrgeh1BnyyU6wplieLBTmVhhsdSn9L+yH4XZOmnAqG8p4L0Wgcg+X
twcduJSYeP/kwBA8eJi0EHKy9b+MMtwUymDQuDlVFipLfBssrKny4lglSfzsi7w2
q2nT86yRjjOLfsnUvVhMi5vEteIwQuxMKSVE3GXdl2OKSrL0rNOYgxtmVTxwPgDt
oJm9NZCs660kVBB/zw0vTK8ZmnV0TlrxV0Lzd3gA/q5UVDFGrhzP0pDuemb7orCC
uJ5gLUEi1GKK+461acawDSwQ7+dWh+wq+AOcYp6UrzF0VmsI0KX2VOoNMc77eX3C
EGP9LA7YOB1Qc6FqTW4UkMwZbuy7P5frnUdfi6ZZm9vUPplLU98I6HDufocTNx5q
QR01SlG3Dyxg1ryBb9ILfjkfQmaoBXxXA3/B3cvBZcYNh0gj+13m89Bhb0b1FPD8
quLy6vA76Md7YNb/+dRR048ahtxVGcAJQumePE1paOBO0b0krJ7Pptc2DPmmd+Ht
x9QMjfS3FbaVtyxyeI1gaPDDi3+jH0SH6HBZVewvNZC+YZh1dRvJqatBLRSiRVkd
exXLJ8Dqk/fmOu6nEKS1soacMz/0uSZYcRsLrCQq7czLQHq/4S4cOvJVO+UF9vDW
/W61ArNlN7lA6LGZIC8BR7Vq/hUEbzube7Z/Tv7pLMCDkFZmpxRaAd2wbjYYUKfV
AGo50ietBRQXJjGrrgRJFjHgRMNPJKIFoTSv2AYuypKzi363bxLnCEXHfmB1ASij
74tlO854JsSc05I5J+CKUZi4a7P+uso780MWFjeJKIS80EJUnYczR9o9iQM8y3g6
GAYIziIIVrKVs66vzPwC4g/wbkRfOdrVTmIiQixCEpVdOF1R894wxDwIKs1/ahfd
CO4X9PGIb47sCiAiU94p61otwTSZ95GqePa6D2Jg7soNLSr0ZLKE2E7kNObfCuRN
iiHuns+lN1JXMIn+DmVMd7OiP/nYLYvtkAQSTgizXInQLqT2xBZ6CaHXNs6qbuRb
hmqF8fXeW0MG9812xz9AqvFpCjFJiZMphbPutEX2hNi2Fahx72JU+zwHyImC1Yqm
LAfZmz1WhmuCmsj6ViyZXelB+gvH2bSOqDX4zjjshNqb2uillutRtzTPgw2o/eBp
rhXg4yc+fXrMID9SDtxhhhwBTEy8P0IxnAGZTLPy3rxlvlhDNXqiaUFhq2eM2a42
+UlfGZXHzBGIptNhHhxazxWcgmnr7OWIzPHecvbgopfYVhfdwIGu4YFnhq6Fuw2G
5Q5h4fR/kzr/IAkBsBLKmfasfFZWFkQsUxVsTgYR4P2cDsKus4AcMoOf7FFSkFPb
8a+qTcC4MbaqboSzvAzi7tY6gO5GFvxBS3kKz7zN6LL6/hhQbNzrizAJvaxvdDL7
caQa2dI3K2HSPRMFk91jMN4ArEmO9F8dHOOO+8FpycE94mZiLLEq+sge7qpr2t7w
BtYRh+2QrTV1PUxZDk8x66jtJCF1q8hbr+K9C/pFA2MgpDdFXjLq61uuan+5fUry
s7+FVzm3XwQSd33aeY2QMD5caGHDCv9C07WKUWFcTM2sIKgJw1SZU2QrnwEs4lTB
vZ2sIJpTzqQcpvJ81js2xM/J2cQAC8L+aVYhJQIXOop8jEjDiG/LMz6CFWWJfHUc
+GtWOAWTJ12GzruivNDcgqk5FMv+tvj6VOyMy0t8F2VkZUdhbuoMrI5AV2IA+1yT
MPzuE33BvY9WtAQlY1nFeVdnr0ht+bJmEXVutqHv4G2l+HRtY38J53SsmGQjMfPQ
WljtwJlejVUD0/ojx2j1Z+rScPtm+od/GOR8nrfIHfHquZaMKWcdgwY7ZCh8g6qH
qdRoEW2AO5J5ZwwbM9z4cylwVcBEy+4fVn/ZeXTElU+LNgSL6MucfldyFZkD9ouQ
+gpWEQchp6PBDL18mNxFQT0e8fFOXXiWw1It7IOnzHLlLnoCIp6CfVO2OqPYmYwK
TisHeHF291ctRWp9ZFVK34wudb48T59yP4KEdoZdtwcc7xMWK5t4xFzvBgCtp/hh
atpT3KBWEfGJmAgyBukweTFfZrOnP0E5lxTEyGoCv1bfS9ntb+os0GR9FzvqPV4K
kZ13mJwxvfx2GVDjj2Xhz/TlqKh8niSoWKpiWNrM3+uOByyAJysxl459lERuCDQR
zOeD6bk91V9hXsXO7cfonLdGtuUOtQOLXn00roJxUV+r8jPZ24rbTfrkXyDC9tkG
qlmoGqyFS2X7DiKcD8pRpI0mJRb95a9PN29VZR8HXIIxt0rmol93ud0Tb7crIVe+
Md/n4MO6UWOXdL2m5JI7hXL1/PsQkNnYTHuMsm57uRkiI5eJ64Xvf/hNvuriY3ev
gFMj0bA0rGd/fhg/nRtZsPz7zQtVTr4r1kmtO/iuezk/5uRQ+9kVLoNZbF+TWCYq
rmaMBP6lcBECrtX1xakIfZN84S+hUuW+YJPGBactaMeHzoIc6PyAmebC017rzS6+
lUCIKVYBhsdpWZtBKIvbySXjY16cOnnmbCm3/bGWuTlVBMqQjZvnO6GyqEX3ojcR
9w34rzHGrGA6pJMh9Cexck21VbvEgiafz0IE/KHKWhFn2AAVl1hRyZ0clHpGXU0w
keMrn2t2sv4WICIBcwE3fY6TQiDPISALGqk/rPluJwMkAGyFpQUudZE27+VVbgdA
L9Vwxg690Nhg3q7eYiompkermWPLyleQtCu0W5kei/zTMIX7jDRX3/aUbl2xk1cQ
xiSThr5tfzBdq0TabPQaUep4mqDlweijJoVY2MYgSWfYFEQtDA7UtW5eR1t0fjxK
vvcb91XcrO1K07lgwW0X11YJCYQsJUYkCxBR0gSGVWy1F3FwjLQQ5t5tC9dgxAJm
axBJbicVBzdNTRRtYzZVe+ehiBmtSbY0uPws9rdMDiruggXPnc/EWQr5XpkU6AA2
sq1bnTWTgaKllNRFoylQvBcQiTQGinMXi9SEOzvU+pDL9VScMQ10W83JHW+EXUKf
zB/9v+MpsTQOr0riAD3pFqcjOjlZhRC+UMJmdjnpkHhbrisw3Pr+Vbi6/orD4Gw1
GAmEJnCwU4NUvJxl3XAkPXxYIeP65O0WMbUn+Sesc2POVGioVHqKhXcNmVt63bFH
2KR7QdxBHccMvXzB5n1vpXMYwE+7CexIIcv4vnxGJyEO5swyCN7LWLHCABUARqB7
OsQUZcLmRhiVvoiilycIIUIB3wet5rcp6Wcha4dbbNp2yr2JkdQnE5Td39sLPd7y
Ya8rneZj1tMl/xdGFmwZgvJAVWkhGf4WsPUWhp5NoCmR5cnN/ViHqtlxyxuWWl/i
BdDbf7OoHQ5LpCpjLVux1GvkvxCH9YkgoUjGPq8Q4IOyn5vmO+DR6frI65If3Izj
BCE+IoRwxir2lXheyjBCX6HAtEBO5nmuNCjeRNvOyIZgzutYAsoPXaTaqAMhJcLs
3fofrA5gIvvEX7ZpInF28CiQmqjkmXmgGQmDUpk+WU+TpVhCF1Qm/4ukUsOZ8YGg
Ryh4bXyyOBZ2bPCTjsOeY2NPmTcjaLQlRLvte+4WyFkMueLE18ItGhpWP4rE2gCF
Nm+bVkdBj3BdGF8wykjfkpvZ7auPYfN1RC7lSUNnh8qEJfUMN0vFpBKrlFWmxKKJ
Xuj0mqZkqwXnW4MX9SOMx0NoO9DxT74WNPNQ+uYa9ME6lbiTkEQBwDfNsTw5NFA+
Eli4YPA4uYXjsDsqKjsHn+qGm5AzN9m/HkNXckmv2trzCLedNlVy3VRSLRB11kda
z2hMEt3QIMHW5S8XDtg+P+BLfBPPV3q/L08lQnpZQFumTLoei7ZCyJGz3/4Bt/b5
cFC7nhrr3EEofDCuY/dIfgzyPNaUTuqCzDvab63o+vU3bmKFjszG3Zwl9Zz7rNUa
+pw7dGigj8iddwfPcua8+BW+53yiWtUWqmojhiFD51PvBTRuLt5ZzC0s4QMfx4rv
bXZbl19MFZfpm/yPPhw9E2D7ZMDavA1pctK9jRR57tji5Uw01EUStVy60Gg1Cwbt
hkRIWLI2MW5cB/0I8nof5SLeNiD+TckxM+nhK529tNMaXeQTP69OxwWUh32Wv/dB
FhlB/5LBEhe86KYxY5heTpUSg6j0gCXV1fK7Lv8xwb3W5dne6Hmo1RBjDRJss9fE
gb8zE7aKsqXGKR3bo47tCnK/NZrB8pTB2GVSRqW59guQ5qDvJuMQmz/gzn2j5nTo
x2fNsbhJKcxV69y/rmTijAkfiQVtv3DT3CO2KcgCaLfP+SNzD5ns8zd/3Oz9qDQZ
os6g5ek+ICohO+xgN+1thvm+VlVrwm1Ip6sIf6jOBLudvtRao+pxjsSFGUf89MGu
DMUYR5OgnBcNFQ98Ct73nYZrwqIwY61Xt7QW6oKgUQaqA4GbRJx7x59Wstk/7nqq
919wogPyQvCGMPOZMbFMJWJPrFj2HXktrcU+gh7WL6/JEZIg3nlhdDviqHSWzAWh
Dk9tj2oMxXWMxI9tsVnyNleezCIai4bX4YVqNNgJumFRqzUMPYHmnh9lpob1Qlgm
K5I7cVO9/Js1/U01NJDDvJBE2gi0r09+PUPTIHGejHDJ7CLFsoXIe7RFgcGR13CJ
X/bC37xKc8dIFmOIIuw8p7RwPGKl9vdz2lx61HuRL9+2i6TxYCaJb6QVG36CCRf3
w9/EitRMcc66ZVxESeCb58Q8G1smUHPj3fKV1RLuYlxvEtrXis377JVmqV7SVXrX
E0Co2MSpsd3+odg337fL0C/YfXsucP1cxTYhPk038sKAgTVg44gAKYsbALjuwKSP
fUDBEoWsIAde4iSsQeklE7w1CqgK35UgECF749G4X5grckiuAXwM6SXN+RInDteF
qHBzkDiMztuIjJpGXWk/gXPAVLMlWhJxS1JYioqbzeqJoWSw9i0e8GZaqCKihS6i
45M/x2bJEGNqMlCv+NjHLAOclUtIU+84cj87RgCfKkrfn4csp8MWuAfflQtqzRVF
uihDKsfpUjT+WSW3zbKRZ24h1wAcpUIPFAOXQMWsuqdPGaEnYVx5/obE/CNShajm
vq3ZSMbyZsa5z1uJ7sBVjdrZxLXExw7GkaYGUE4QmjYFD70R72yAXxtRtaaN4L9Y
1cMNMXmudpjQ5nje/Ux5COIiHmfxQqdvzB1Cb9Tvzm+bl5t/8peryYQGE0rg0HzP
iSZanDHf0RKvfuJELtQyq2/DN1aK3EgQ1mivMcYYhGsVc2LaRzWQ7wsGnja790AI
XDP4aKLbM7Mprb/U2+2m/tWIj57gcL6j1cdQ1LGN10lb0RVjgVIKZF3sYZerwBg2
lrZJDqASbzdOgK70aBa9AP+sgu9nzqxl0fsrKYPLyyY98RyNhAZLU2Bg0XoUBpIw
UBWgd74kjD+//5TYVXokdrkeKjwSdVAtYG/lhy4tTanmG632zFBP/lvPXSsvPq4Q
4EZvjGlxe2Q3j5T9iPhImtnhXVRTPyrkqHWfHLaGaMJDnMqde6bEpZZUAQus6F6z
jhq9kHYXma2hMvmEd4k8TufegkXEN2xo05aRSQeOseCiqU5Y4ynyAvObPvIwe0X+
sl+8kAQxYHInLAA2qQkVV4GIylOQ5YtLn7PBrV8AOFYWs6rmMoRrSCqt0po7HzRF
6hhcHejEzHVHtkIBWEecTjeb+IgzqOAcfL/Y7fK2wMAredyjsWWafyJpCgXOAErG
mEI6IzQVlApheGbJSyJym2YmkZiMy2JfXl4X6lP4RrmVM0j9y/zn+CNcmAI7VVOs
KDgpSvV2DFRje2xWRk559EBxhlh4ETQUOeryjyLYEi9DHkiLwGdp6/xGwMru6n/r
13aCc2Xdqut9ba7Wx4OLxBge2i7dxHsAULusOhuXMR/LAGBwIgOfPUqgIPifaWMt
SZuUgGoVvF3BPdSd0xkhB0lmjH3JOSLG99bcX20KjCQ0CxOL0jZXTVzpltAeSlI7
t1EPrDQiUMaqTQqtdl4rNPoc5tcoi7qUSFUe2UwIbDXT8IdEQfS+CaeoyFTCNBCA
0EeRP5o+CPL/kgS2FSlhkH9862UDK1wLlJ8ISRH9jmATK0x6uYIleuYyr8/VyWEj
4rFJsSjtZVxnzzZA2TvuWEkvV4R4xJnD5fXOhG8mSRVtIv6hor0gRnXDvhm9tDPs
5IcdYvJGRFiOid+J7cWPJRbJmM3RwdHbZe1nKzbSC4JIdPGdyqGyvbfq6ZjjVCWj
irWyBNIO5jR1hoki8xvo+S5d0gyUKihsaPS/HbgTjXTVoYsAWKjoZAlOEaHy/4i3
2I+ZT1T3LlLXFv55zI/3GKE3CLHlfUNGL0J7fe6iLKZgo64ik1O1sv2bDOAvMd2a
OiCdjfYjTY7V6ihWlkj6NfVKL1ILrWQe3bzAevgJMOvgy4bE0xavbHngdznm+bcP
JRXLBO6QXI1dinu6IQ8Rf+ohlmz2xuM6zNgTYHFZuUwwZPiRZURKaHbz8OEBIFj+
QGMJNl84/aDa89boi7fTwqP81TwnyaxjSGlYzxxPejj12Yq1HM832Vv39I5gp0PT
h7jzTE7fsH5/lQZnS8729+OrAHTNtnv8homXKlO/87rkDSzORd9o3QLfu7/6olP0
ULZDNzdoELqACvgJGyJI/D47qv6GHLUqYMnYFKEfHF548a3HbohmqIGZWtLPw+h5
KQGS5+YJKvQXM1ZL2mct6P/OgT6MrJyr4bBRAAE98VTDLswpAxgpxmLAQJivFS6k
SZObuS6jU/8NHFLnh+ProoIGa3tDovtmGoy4Sz/deQWex4Delze4aNeE6xbAKTiA
1xj8cmDB0V+f+tq+tQCTwrNBpVIng4aoxclOPB4On+iTc+XMHy1nnrMyMHZ3v8Ku
RuDnr4mY8TCmG99UBEVOZ8yd7ZPEIiH5UfPkwP0+7CArLE9RHMJWXWQaiIsypoZv
pEflhTiUgBqsKfTMCOyhMrtPyxMYW0NTBqkVJwk2i2VqL0InMZFsSgK6Lx9ruKwQ
S+l5k0kvK8vIsOnwZONlOZUqLGM5Lj99EJIJMbGltsCF6A0LcN8OKRlCEsRPZQ77
Lr9vxLOTD3MMmrlbwZP5F/R44Ycn5D4aqHmoNjZ6r1PV/ulw960GoZgTOBfyzavC
XAC2bqK4mc4uN9HMbwjybDi9Uj2J6YpOHsHlF8udmhrvvUxQI9YwRG6Lq0aAsk8X
UnIKzTaI/TPOxwFcPFOeiVTh3yf+zKRCoCT/5f5yxRfnrADvO4MRIc0Od9vtGeKO
4BMibtMn4Mzb5VRJsIbOtOPk/kAWdWfulH8hTF20Hou2EIDpXVeRE6vkvjgkNWPr
8DjPAD5wORu/Y3LpEtRP55yLsD73gs03ju+qC4RBNWjFXGwKIUKsvIaSRgH0Z8gQ
ixygkx9/lsaUbtpZTGiD3coBUSvSqMDFcroYLg3G3ykajqKEBrp1X81PGpXNYTye
Kqcs9Os7TucZfxd5k88+qCQUD64FX9MEd6u8uezHHj9LU+a+u0akYB686eUYqzNP
CgDuCb77JEq/K+fl5fIYu43CoGuLuV99jzstMaznyL31EN+OeTjGzUpt44EBRdF6
KRVv7VisIayhvBDEGcADFGLjehqaLD8kgeHOMwcLUVxsqW/vqjIlhQPLNjoSTKkV
3woTmCLhqXgjOj5+twmHsn8Mo7GUfW+ojgJwx4/frfOd+lyPzHf1XkQt//HsxRe/
EVuH+HqOzMCcpDnTwubxaI9Tppbbl7P6+ppPS82mvN6BQ+x3I83oKHyWQ534OY5W
E5KfkejGy3sIk3HEBqqYK9mpdvVrlzglwBB6e44Rf2RPtdWRXouafo8TFhTads4q
aFYl/U26yqD3RlhDAZBgsh9Ifn3udIsmCBOXoeGJ5vcF7YoL2xIoc4c+er+oL06J
yfOn5D2U7eFKCVqEx2xIKaEap5v7sjopV7V2TziB9bMt2pSeuzuVWavrj22Jm81H
jgx5yZTBXygJH6yaW5S6ydPQu810YHVgaYH8XS8OWYfFk7K2X0NjLUVxvIfuyuOc
wR8ungnh9Kab4+wFp8EEArim3Tne77njF/O+pST1biLemH5NA8u+H84TuBXSPYzE
toni+Gvxvpt5nEtfWQc9XeTjpFkbqo35C74GriZQ3z5AT3imKX7C4h6Gdu2sfVYi
RUVPhgYZNTMhM1Izn464zedE+77nfGUdcVM3TC7wgrQ83r6LOK1sCsYCmYRT3MhB
4ZZGmHSC0nTotT9d0Jn2UcrJks9ygnF7S+VQ7FSwqbygmJNBe+hG/QyjMoDsbUpm
cUrkQePrGv2oIWnjYJuJ/Fid08j0TX28pspSkl9vOFS48OunXS1hJp/1zT/2eizn
Ah/LOoAc0XPhQa2ifXKeyXgjVOOartL9ApkoApQNDHhmQpC0BiLHV+Z5wUz/+nAg
BzqHyPWu61DUePAytLii/3ZGiobxfx4ozW8kHjFUY0NpIsmrvWKvyCZ7afF/y7kF
GMOGPqzP57HpbdJyLvS5IiujE5pv7XdZYSTbDpw4QEjEgixy+hJDBDk9WdmEFivQ
XMyttNXMLsKznx10BGL4HJHwG/oLPBUJjntMEYGNuCuZkWLyrkJblE7J/998ubix
v4LLYtqKtjVT2+sCF7tPO+xRY5gZovTOk5Tkn3g+9St4ezdy+ak2XwoBoh8XCBW/
q6o7VQGO3sCkvso+g7qfZcm2bfDKjPFPCP9cPYc/kKBu32GI/Zy3I4Rp07A5dWXR
TCYt21kFwTEwTfOgBhqq46BdLRaWQL/xu17NDSSPxHZ+adbEey/juL7oFb6Meoi0
OXVERxYfGlsMIDn0GOeNy8LgLfpd+s0dLrvC0kQ9U7BXyjXh55Z/R6ACyrvVDaXu
u4DwoF2hUgDVbTo363k6v0UZhvDWiCczAB5J6jURAfZcL+BD2wWCTKPwTkeJC/2f
Fk016UxYvUI/gAw2I1SGcON/gLJVsmSu/HytzaA3tCm7zsPuaY7O2wzDkHGBS5oR
nRKjEVxVJrA2kJIGRj33hg1dgIFDUnx67cx/W8XM/NVriIR1/bj/luNTuFyOLj7r
fdvTAFn/G2G8Ilqumqzxtmi68Dc71CdYw7MI34LdcPM8xcMJSdCEwwi+pRMlPb3y
2CJkjydwUZDn6ZCCCM6ZhgXle2gUXUZddyg46rBa9J24xmfFSWUCObeyrGh63BaF
e89ha03I0+OomjT6SSyfODqwEI1VDgO1V01ONmzkUB8X+sr0VnxSKKJ+HNdahcz0
DtzU+G/RqlpaHeIQUaoeSwFVfxyKH2/zyYlsU0+mlHt7JwaPJMQZXcWt+qB79/Qd
PfexIIj0gpWyRfrS1VbmECUUKmGrJm5sP/OcAZpLbE6owb/pPY/0Zjdzi3a3dKgX
0ekai15EyGtiZOtc9WPDrtRMqHqd1D3yoUfEbfcaYUbV0YD3MeRfZa1Mzm7H1ZSn
VKYiNrDENMY8XcRqCOSLpVISEaufOx7zxv7hNy7sEJI6KsAYWSt38XpK7swthrXz
DWXdXCqZ3g5Nq+V2ChkDexzqgP+1NHwP6yBz6n6Lcenl+TdhYFhJOMSr4z2kt/cm
5C5JwworNzgoJes0V1pKBC/IebucMowIluD+jk2aEzTtoxOeBysBg18L4A6Mk7tf
JJ7FUlpmdRAmgHZ4j1IKc396Uv2tHL7hSh0mImXOggfok6g1qPHHO8jJypSDPoxB
Z5eYqrp9U97Xg9pWF2n8AkY0D80JSvYFaOTzYiJ6SIPAuXA2DgzgxIE0RWHgT76O
tJrWUy91NNNf93kQL0d7i/PkJq8FYrxv4jYnswuNA2MFM0G5yLr4JfeaUwJH7KSC
lMfy091Q7bjQeMNizz1fhmU3bBBM7OM1lPSRVLw+s7ogZ1hRq49kXss0rYOG4FrS
iA6QuK0bIytBPcdwbAyZbU/XzvF8Idy4Y9uYM5UsmJFN54AhMCWo6EMU7daJ65qD
mXhZcVWDqJL2iUiByhTiyMkGcP6ECZNlRuiLSrc5l6k6rLtC1WAB1fxPN5YJnY4K
qraW2x4IThq+liCxXZfF0s6QCo/ugKtMNznnEcyKyGesJa8XUAZhLW5b1VNemSmW
paOcm6m2uWT5+yu94EmWlIShdMH0RxxMd7D+Jlut2j815qswtk9/9tHIHTD2+mRJ
NaDesZcWb1NrGbA7lD+EzJHTjPckZHWUv2EKgqu5Vnelb6oJJ6wlRk0S78UsO0St
hiqC66bVKk2PcRXAMjz8Bprd/SNOVRBoEvQ9AMDoVgFJzPML/3FDxlFnMW/4Obze
OzWUxWgI3iS2VJ6ttuktChKfumd57ZaQnejm12WtUSRihEyvF4Q1zBbudcV55RAw
+zHp98/2jf3cubVN/LwHceb1Ioth5dx0oTnqq+bi136LNfZIZbXsBzhdvrRfUhIv
NRksrCqjwRIzxn1h74WC9Asl4sPtFAdp5JVATBB5NTuzrhJp0ME9w2rsy6rB7xwS
7hRNJsDl+iTxORHz3ix/StobVKFF6S3vXpNpaJO8Emq2eGlPNVgB5YZC8Mv3lQXD
/cnr9EnMR0MdUPm6fg9ca6GPsD+DOPlVUPt6b5luwrZAXdgUhI2MuqPD2RryFyML
FT38AjNa+2oKx0BhWdzKKmLkuhHTd6PBi1e7ja6Dps1aC5vH/6UkBQIT/YLhP+pU
txo4O8RYxnJs5ys/vM8DGuNcwSJuXoHrD4xArdVe/vX42cJFzEQ2F9ApI61HoIxP
LnvHOAi3RHVnya0wPISg8sudW7pIArVzX98b8J+JVLyytLkcI2PeekwlScko19WS
JP4seHP5hCOjF0Xpsl7WQPVqZjudceKUniVserBvEsD67IOBEnLCPFpiHQfI4uWa
k3EFPOWlTZCXm1f/coTWQY8EwD7y13SJf3VFp4fNVMMaXxxNiF9Y+J0T0fKW/QKR
RuipzA5sJYP9TdgLIhNGEXnyMwT4QhbTe/m/pFcMa3CX4Gz/Z1GkZ3YR8SusZYyf
wj7Q672qsHnvKBJuLDVghea65JKHT2Sw5zltqb2v3j6BCn4XhQtdDkVAVub0dZnl
Y8YAmOl3UYQKrjAS7vTFZTt27bb/CmkhmXvfTzgMLZiYpf4dGksCsbh8UWipcu5l
GD+Vji3FQIKRuVghyLD9olPqyfEX46nSTzKW7/W7v933fAUz9Ol5wR5rQpYEHMSb
Mo13SmZaQyTEHwUWYMfgFMBdDxhvBB9WS0lpg6HyHCuXbDth5yYuZ0m/Pew45Qw7
nZBaDNNCNypbVqLsl2zJxSfU144RwY1uDdkC9855COJg8W3t9PLHaymOLN9jaj7f
AbYzMsoSnVPmXxwLM/3L/6/oL+uVukojopGRzqd90LG6wAIMm6wxX03sSRhgbt0t
YL2DErseFV7+DTMj5Tpt8ntAJ3nA6dWXY/+vmwMC7Vuvjr/tkBMX1UPeZupFyvdD
/wqMQgbH9OjOV7aRhTuElMXpXCpvdchGxAW+1AJxnV2t53/eN2tJ17RvpWCtbAfa
4kdW3/2axteJtbTLF0b6bunmuqH8SIicHSsbwDkiXdmF1V/rZnvYQv+KveKAztQd
O09caY2ApyBtZUPZtvDgfvzLkHghUcwusN4VJS5jotlq5s3lZw9P79ZloJ8TO00C
X0+bdn143UWTwPDZOTnfbrafO2bs3RUuAvwWgCp783MoU+Phs6MJ3SRXNvvUOBZD
Q+iuywRo/AU5ZX6qxErXNcuug8HzPHnZPxBFXbfA2pwXfzpg8ErrLVAGemUWkdIR
I+MCNZAMM80LJ+14pdJYEXdS7sbyPonR6e/dg+g8SU8bRsOcO/XAXpLEDnh6eLKk
xnEmYrF1rzNPr5BpcfyPm4qCaCpWqlGNgPLuNYsLxk/pl3axHph/8eEvN8mNv0UQ
UxqZcvq6aQUsy2LR+kd3nR4CLfCRFwzqWv8P5c6Obfw+nBK0uBUn1Ssxa/+eI9sO
vgod2gd/EK3/HqgIfd1TEJpOtBs8ODhYM47ctQffgBQ5jL+/nL+FWOgryoWyfbOh
ghiB6o6MOMEtmujVZ9Fd8lVo3CF0UQf//U0J2nHBsxufm9now9I2nrko1lm/axkS
E2LGPI9nB7rRivQHUPQF3awPgjii8E7SXix9luCtAwLAa7OWBj26MWd9UbfRRNdU
xrD3HocEfTEov7hmPiA72sIDrt8lL8nJEH1fTyuhIyFBWsegNDP6NW0rIozgbs65
uwgEK2S4GQhKpeiL3Q4aylUEgAZRmEGICoB/DsC65BavlYHhtMuUrBI0jfU3LOIb
aV4Ir7ghNMRu/kuQbsy+F04xXGycKAP1uCDN9ryawo97zzFMUdGorRE8aTjNQ8yD
VlnoBhScq+LSt10S3ScOzrw38NaP16pzjgtmvRoe8hgJadIg+BlOaRuvrceDPSeK
hhxSaTLksPsAccqv9cjZI24Vz1ZMqiZF2UM6dwKjTwtt/i7g26YcqCui3fmLq7Qz
xd66WQ0E5iPDcTeJn8poFCS+7fj+YOGk91yU6niddq3iM3OJsZWtfCnqhFv2AIMW
yEoB6TcFsqa+2GK6U2QZM8d1WtrbA315uF8or2+inZyGigbHWqN5G44HfhGAsnYE
07T2++U1oKeFvHM/d/elQAI4nssds9z8ycxiSD8sW6N7SxQ1WiAUNXuhd8cHx/KG
ufO0q5MJHptY14XrIvvUDkm0lnp3AHsHt8ByT7652s4ycCqMJU6q70qFCikTe8Pb
W20aalOA+jnpcOl+5h304UxzdlQUSR6hD0WKPCavDbEpwZqB5AYeJnoQPd968GTM
yEoIxKhiG6zE7q49+tVzbuOtZEoWF68gUb8An8GkCKJ42g6aFKQMqF9mwxPzK9Y0
7B/gTHB6jDqiI5YBsS1ZLRwEJizJKkgsMyWZu570USoc+I9GBFMygnvjO6LbqAcx
OhNS7m4+tkiGyTo5VbJUp16Psv7K3QLJJzVK/LrrZYCdzKs2WEegyj4Yi3oL9p2s
Vd/gtKY823eIvUb2Po12QBrAB2we/i/MIpn0A+WWYy8ZMijgom8cLdVgJ6c/EgNu
tJHjzCghPmZKdN/q+2irMedyMBzvYMsaFy1wDu8DXiOkBVqmL5qFE8PGtkqcEbIs
U1/F2cgdRdotRkuoWyFuZ1f2/c7Vr7yIyBC8+GC4zbKQ0niFCdXF6B6WsWqyEeLw
LFMq2co6H92ulBywFpBjMXThOzJtGe8g4aGzhoRgn7V9xM5hCnJENKFMkH7dhHZg
2ruXxVA2YlUAHkGyICPH4cat50yKM4XmN/bSUfl5Ltfh9VUuk51qCGJbWmr8eAxV
O/0c2iGyRUzbrP49EMInpDqmgxL0bI/S76V0eaW8CFfjQaOz9iKsxM1KRYAf0pf/
dJacCySvFkJ9qKnqY2m2Y7gpK1U1CVrDVdHVaZBJZXgTHnVSbZkTbyXI7BklsEs7
xDJ1QSEJSAx+bb6PR+YF0MtQ82kXGnyrQjDBNj3bgXXpAWd4LIrsH2FneESbO18b
uaUMbm1wzOUPJ5NqMRwSSOGNgH3bWTm4cUFDCZAGtO/9ioZBUaEGU3XWqUiqO2J/
eS83bYW0zyA8AS1fPB2ODikZqhBoLGaoe+eysghB/wLfp6i/mO/oQYm8t3Z+fWx0
Yqj1Cmpe6pAdMGLcvYmBd4bYAXGrAcvUwS1Gv7D4LEV0T9yXa+RFuu0as5LO4/GM
SAGWxe2QeR0hrsZLjhcSpbMCHxnkq+qTHAnnQ0MsUXNvrzydtUyPZAqW3cuY76/C
dI61ARMv4t6O2d4Cqr93J+XgbYKyZ9cDdvfh8CYmW85waTRZ0NtAjR1FnkFUizPY
O/luHKBl0IdemL6WMbsk84VAJOr1AHCaDB44I3odAIOPVf/B6d56gC5v6m3/du0J
mYxkkjFxcvXswvFTHUYrzXYaR+pXDGFp4aQ5iT4YJLkWa+/x25ggRHQm0qTlJ3kC
0v8VKdVOvnBu5FCl3UYHKwp+A9qczlQrevJr913j/K45IXxwK+H6UsCSDl12URG+
ZMspOe8BjbhgGzlQPks2w6fkb6fK/7C5z6Gt4xcMjdoqv8CDg0XLPPAZJsfHbsJB
fLjeyHJn7n5UiPdECAZBXJ3xhFANdIW3hH7BNlgHZTU+MwbqlB46ZO2+7UE9O6K1
dT1yeAO3ZGdOwiUH1qsnzQ0X3ThWn28m8Fd4fIcCZSH8XUaYGrJ68JDZEKgB1MfH
ZLq5NMoxACudJoQfkbjzDMsGWBf4oshe9ppQvAVi1KApQeapHfyf+na38ewin02Y
H9PTpcQmDCwjX5upI8lGd3b94WwAZulu5hpZy+c224sKWDBxzr4hMKujRKjkHeyg
XaFPDPY50BjOBwXHmolyC2zRWhUhGFxLonf22zZ+VtiHZZJo9sQjqixDdPChJh4K
f0S6pCrVO+d+hkIp29K+mwclP6lMSqVfPsNC4NA91zWrgWTiMPrOLac+XRjbdPz2
a9csoXxMDiAPDxJNMwii7NPuNIEfl7Zqu6VAHKGr+24kOmG0ZxXOixeQ5gNlGJbB
sqHd4TRUC/76DM6HKGhADY3fLrR0Q28d8ffR3lTScDgh3gjoxSCjZggxwLB8VlNV
cvs1i8u+eM/qEKUMiIz/upqdd6BhtzRggmg5xAZkXOPwNuhBM+UcAIxgC+kS/Kur
Ejvs4n4G1jpHis5EH8/e8js1ENZbfnDxdQo+OWnLNi8v4ZHijRBL7ryW4EuxaGYR
0iFeJKuG/JA8kcnmJn1+Yr0DWCwLQdlqxEYYPaPcJ9R+FlBb+6OpCmWbaSC9F16q
TS384Oa5m9K9fxOMRKHRmvfUaxz9lD8IXVwUEGM7J9kWpQJtfrMscsl9fRaohReX
L5e6nFRcbgK5p6P50laFQbnNu38njx73aUw1yLUTo6ggr8sGpXjlJsF5PS3RTV16
+ZB4ar0S/gpVix+yB2DKum5L5d9eqZVtN1EBg85LsFKN4HDDQkmKW8D3XdY7tkdQ
phDas+YQmmN5rjCeBL6NSUP4zGVSMem0xjL/qDHwubY9eymajN23MQlqZNolo6Gy
zRaEtttoGd+zcRIY5dNWDqun5KSb46ungAeZPSc1MVzSEB4kM5dkrjbZQ7shJY8o
rnk1rR6A6i957eQUgobTL5/2O1OfjY1fAZEj3VRzN5xvK7qnOg5L+S/j2dI7GAmX
xYiYnVms3kcK0Dok8WLPMOgcMW5FbiS1xZMyy1qzxtj5I5gloHci7HNP3W4o0ooW
7UYAfdL/qi4B7MSELuUjE2nhiONkoR/JBLl1t1ZMzkamgM8oC3DZKKF55Z9tyRQb
U3iO5xY1StcvNdEqlX7a0KnoEqZqqNnqNfvrJSsJH3L4LUDzXxskv6oSP667YlFe
JwiqYtEv78QizyTphfEkRGVkl0ZZ5nbJ2kVIiNdeI9g/l4ogiLSUfGf1n5/vklef
/Jc/IqcOP7n/vtnw1QCMq+ZA/8eaREmz5GQCiSWiz4uJB3+289YFEjSgjFqrE4oq
IdHXoMLV3buWkpeYpgd/74RJY3EMk7PbeQw0v3MZLRFUMj1CmrAMLxLj7ceI9gze
nd9oLkAOf6/y/TE9PGqRZlbkvNlbqm0Y85ZCfeJKsjSvK4L3XjgWaBlzGQ0NwwZd
pi8Rc3nH7J+jHf91FyiVedjeYUHb2IT547+EZJZX4oT6iFWJ3/uShXENENVmCIk4
mzaqm/os8/qUHzpLIVliwr/y8/sgYdg9jTwPE/1GKN1M5CaM38p4Vc4VbdQzR5do
Vgc/8JYV/c7exwzxi2Rl9a6F48yw5MYNtmgUJO6Dxr84JnbWxZRyjgbRfmMCfaqj
ijvzgAG2vsD+8g26x5iu/L9DuKK0eyVe7kDXeLE96owbS1FzFclO+rhqojGtMtqR
ukdcC7kBDoSwKRGDFQZKVf5EmIMITPpvn2r83ZcuTDwSwLYRezcevuH99RTjeQDQ
FzjZY421ZK0AqrLVQe5wR9S2R7ZKzJeqtDu18cWKvVi8iMB7nOuUkD8CipIXAKAY
QOF8nDiWBNMwnyfusyA8FY26U2L/pOZ/IstTCFc/F3Uc5CH09GvmRiMsjo34Lun1
XKoesrGpcqe8rPv94RKa3VlGqcS33eZC4zYAqs0p0b/hd85dLtzRRXBRbt90ANUf
YXyBKv0HVOrXTw1UsNnKL/pEjuL1Rg1v/7XKthc1FwpluA4YEBrhmbHckg3pen/D
POELcIsJsd0rChECV4EdKOeYfv6U91//vzfpx3/4cVdyw/SNOJuD2iSkAV8vp7iP
KSyI6Qfl3PLYKrgMqCRha1CPhEqMxJpPs+t6XmtngoN31HucHU94N7XVfzX/6/nt
GKJGAwfwThwm8AjZsGbTovK7JK1MNb88a4ABKoxI5RBG6/CI9cYlrC7S89niAVms
YZ5W+rEIxMWwzg5OKLJuroTDxEDPmFEUiaKEQvrNI1jzEnlIoQXWkCw5l6OrbQtY
Lye7k2D2xaA7X0aThULkBreNmfIUX6STJ7Qbk5w+/PrfRdygrTUbnjtsU3TcdDOZ
5NNrAibJR1OmtJNldowEVDVD1czZMnZYok34xtUS9KGrtSgNIlpP4T1tdt8b0Gwc
vHDwaEmtDBT1ZNDAdD9zgeSg5BdkODoQ8qhvbD23eE6Ocj8qoTYHz8iNzVGdeiIt
M5S3S0n+zXq/2iiu2S/bv/Y6JBcqVv8ILd+67Xl3xL8SmFwWu+/T9WPTm7MEnCWQ
BUthGQngScn3Az1Hkl6pupaMk+yHhNaMzCJX4hW+TNVg59csXGVqLKCa/h9Q3UYg
vyvcH2rgaLd/peXE764P6hPuJwHWGiB2l3VjFGhuTyztRh7PS/iEFCv5SfURUEk9
pd729Y3l9PkIoSz1Xrgw9Rd4baAK6hkFqmJbgPQqoe8MWL2cZ8CNNfpROplhV5yY
Jr8nqaaO+wyBOvnOBa7H6kg1hWtoTtN5X0IS0ikZdbNABWOMOFpolDIDxA60xj46
AmzBOmnTZu5Ndkj+AA0VcpwvvBUehFMnyGn5UwUcrOXcbcqgoQuY68Kxe33byghH
Z6bPnc9F9siFxORSZ6jDE0NtNqeukxvd7YBB29qTzaM/RgzXI6uN63ABFXW4xzhe
OqvdX3Lcl2UK4V5vxe1at8hXNsVb0NdaNo74F/dDRpMSsawxzn1WIxXuJ21lzThu
HQrSHqQXx4YHIsnzEbQ5ieCKvsEadmA3IVbUK8I7+yXGE1lJbN+g7iRwfZWizejQ
G4qbpeQ5yZTzOyVP7ypGSN0UHdcEcAldgmMYcdVJs/DkhI+fZC3+hV/Rxink7LtX
3PG+pVLmthHPrKUL9y0YL0VO/xUlb8HGyXemEnQnkWhlTA8Aa+IqMi/irePdKOor
/GTq0E09imK4dJt5EOQ2OtjDNoxB1QeGY88mQ3mfKXgTKxepjSM5PoLarU85GMQj
Wul+sMDwvmYcyyEl7KwS8FVJG6PktgzIIusXMnCao4WmAzma66lUxLMt6T1+20GL
EBQbUDyYMcvcJv9MeO/Dh25nxfLvkwec1obkM3uuZslJyreJ+yo8VpVaWu1L7ldB
J29133DHjp4sgsFwKhPES1CiIvIgUfUmy3z4f5VI5nBqGYSfxZ2RzxI8xXjOO1EE
7j9416zmJFOMRVtjVk8z1mMKQSnm9/94i8Ga8kLI4TZUMJts59ZAIuhKBVSqxIJ8
rbY8PMbx82spWlPu8abtZBH1noBVgxMN9JyaZf2DPSCK9wBrfyssSxhf0PY507mG
4+cEGJLDYhA0EuwDBpPJkF5fjmagPgpZ8AJkV3rkuFj2fUwjVSAjePuQH5GSzxRA
zMSPsUQSROz9nowe05T2HWv60Pd/If3xp0xmH0KBLLPbm6C0ydZzgTJd2Stcygsl
HXWn4yDXkp7U/2JMojvS8c8Q5zAaH3gELD+d7fG2w4PD+nKDmB6SqxkumOWSkXYd
j4eVs6Yzb25ljZCBvlLVvUoxEjm4yuR5wEjyAX0x67SohvaExgR/HPOMGl6DlZz1
PnGqbA+r0U4jWMdUs5H3oxfKJZu/zhUXgd3JZRb8E4hXjAfczYjUEneEN9Yt6ZEG
HzqjwNe3+C8Kp0Bml5eAIwxNsZ3LRWOiTaGpoVBDd7vafMu8SRgQcAlm6CwsR8P6
1uORg7h9gHMvALX+lFzMGaN5J/QETU5xM9HhWBukW6EzR43Q7Eu7PdARvkcmhpQj
en9M4m5S345I3YKmC/GA2XdVPZNEDFGngr4yxGR7/UdpUxc65znHv4Snb7hQhFJi
g8vPgabUF+zKvFi4BNs1X0+iwF9JEF8d95PnLhfyJJiYFU2oRMVDUT4WPgmeh3Gk
GIzybPq3oJbs+kdgTQopgNf23GQgqvMCwaIgTP6JlSKR5hsiVJACls5N1xvX9F4f
p/UpkMDR2qWy8OYj72mLpEHT4G8JbvFyD/kfih2FzO8ZQ6IunJL2WSJD/FuxQnhu
kfQT50xid300DA87fQA9/Vv+ggy8zN41AtojuTADyLpqUNGxjICtCD6Qpb5/kvqL
s+ooMZ3dhyCHQtr3df1U2qOksrH1EMVXUhCIru6QC5bOrEdPZ4ndQHL+G9bByNPj
2ABWb1QSIw+XMfFjY1HQGOU8WaZYtoFsPEqTTcQBhBdMKbxEJ3aoIcqiyLW6I+ik
zQBnm/63BQCYeQBm2ehSGAPYLNvJIC6axx2NLQC3zXHzzgkm/Gq1J0rk3tINR/zF
fv31JYgyX76TYb858y5+rphUJoDN0TbRH39j+zDtLwIhpuznABRcDq8cNL9nkyPO
BEkP7OP91aRmyc4GFub5HipykCgNeDv9BY5ezcE93D2HHeyiu9Fh1SepKSaH01Qt
LIe+q0a7LbER22lOoc3aK3yfcQq2JUGzwLtE/6oES+8gLigAGtOuwqhb8cAPMgsy
2PEuxVPODKh7pmVvb2ZItvBXFI43Xjk4r867TbLy5LCpmAkUXjeu6L85srpLV609
w4jpRtRi1lrYNx9jKYepBXg8kkvzbkZAXXsYp+peNfnSYU/1sdHfLa81+rzIUxUe
MtAMdGxcTCKu3DnLpV5/IIhEtEBYFROv70H/aBq0zge4q1YPjzn0piqTpvbBh4kY
m8tWLT3hppT84kWMYZ6vBoF3jECqNQGUNcQllZv2VIGIORrNwYMbF6jSokRrTed1
HoG/U6wZ9JF3lC6jvseYX2ZsqskrhRk2MoP2TblIFw8I3f7ytHmNCsB/fTRfSCJd
4YZJtjJnL9g7NbwJ9Kvjg2LAuj3eKJDIbAzDNKlnDG/nQ4IFBpDP33vvBgLNdHDM
0KjC0WX9buvjoei9TiFFDpYky0c++Cq0M6KdEHORHB8aLGqZe8gh/cSWVpk3CHVo
wvkTjviwWTy1PN4NrVjYG9gsATZ5zQHxh2lNK2sW1LX0LcE9rJEl4HptUxFpOjRN
yqjr+KjxRdxe9PBIxEVHe7SPRYcJO5GCvUyLDLG40DZzXvEClHXkbPmT7QgGs3MG
7PxsiZ5LIbplt+wbGmigbDgWpaRGFCfd1CgJGR2P5EffqSKGXQ7ebF/61kL9C7jh
BHPFJPg/E4RWi8sQp4AgxnCi2J+qNauC9rJ6l0ILcAlWIOhrtfZvwifzAv/vooJs
0Pad2ts2T5lCLK0dMBzYVkLsjrac/UnzwR5teeejWPA/vps5XY/6NlrYhqNgvY5q
hjV3WuWjqfo/uUJlUu2PFF7reFc0jL8YJ7MY29hrzfZI8tvpTEU4KVemK2rCP8fL
htLH2WGpeoEzgwelpEc4Kk2cMbJliP5VmHILidnKDA0zHOicaBZDSaSDqIafTrie
H8YWGQuakAT8jsJXJ7wfUEjP8f02ARahDp1pBBamKj4mv05OU4qfW6LIl99c1Jcj
OGICo/W5EyO89ntNPzKGZfnt5/BgpTPVaIC7gv9VonGn1S+PQM/ZlNyxFc4c00na
WG0HUnY/MS5GCLXr7QEe64iXzYO/PPSBDINNkNq61XlZDfgY1qTGTwlGxftSQNry
S6T8l1CDw9DgdmGWoiTJYeP+vBBE9e0kDUsyo9hK/63eqTFXgeL0kyQykj6cOyr/
BYnt7Xl380OL6GDh5uHCPFMnPaps9MNxZTGrNs3u86NcpiiYeIAWiQ0SkdsLAW8W
xiVXSdiGnggaIXGJU+Hj8e5Tehb2fCZPkeskfkl+AxGwi3Qqu62x21Z5ufAsi2rO
SdeK5CsI+dKzuUiVcGjYhHMVHiFLCcPDDN20jSAGYQge+dxoWw1+BBQOWGZXiKze
I3lsB8TGFbt6GVs79I4SqxJBwrP+Tju66PPlXySN5F5hiGu/j5Y9OQkMZWB06kFl
KV3Z+T/TaE5hymtF1eLrJhGbf5Ogb3bPypAps9rkhhVNlNzgNB3PujU73I2M7/2d
1jRLgBJdDh4DKbccaXxZgwdh8P8klLW53GbiaLV2gowYTrsagVi5liJFubbYj+hH
ZdTZJNnt9rsRFJ2aIb5YiokqCQZFjeu0WegaMefro3zy5lzKHL301gZLSWFwe9kZ
0PvdU6YK/piVMccHTOq0fg+LtmskG4x/4p1NcXHMnZ57xUQAE8VMQNyEw/fthNbo
Xzp3pjJF5n8amm3f5rZlnZYG3ZVv+33N/jC1gajmqOu3d4bnIgfPUCDrqbL/dERx
eGr5QvXpSGAXihEWSUM9cwddikNmfcxzAD+k+m5yhbzaw1q3s1aOxdOAQkRSnIPv
iFwrUODj4Ws1AqimMzpvODd/UNwq/sFVTeu3+EpbGjVn33nbJSvGoHp9oOPXyKmh
DFdXzCZgtffWAS+eW45caQsWIPCszqIucHOGbE7mCwPLkSDbjlMwusmBsebOBPda
rJWMmI1FoJtekcVUdMdBEptkcrUe7K8JUO3B50R7FLwU9IMUetStwfvGvHXIoHK+
61BR7JjIkpfSYmtn2SeQd8i12TbgJapG82le/NeMCxXZxTkP9QvYuHmegwPOhuUb
c8bz7G//GpUOQax/KzNZmbW9n+egHPF/LlpthiqNbdejVMI2pGYM+4xzhx5EX9qi
zopJ0aOAbLlRaMebAuatN3m+yuVT8DLdSKuVOOUPLsVg+w4pwwbDWRw4nwrEJV+/
56Rw6zLt06KLWlWzyjW+bA4Y1e/vU4wITK/lXp//ogLtoCly8qHu3Wh/Xwnoe12I
jwzRE24/WDJssSwh8OnCxjlCTeRSq8iCUNpERhswtoLwxyidTfQFViUZajmuNYjW
Bzb9AkPYex6lbTWHPab7sY8DpyoTNOSdc8Gifyx2dXewIOXodVJ0Z6LDXs+6Yo4H
PTRCvDTm1sHXRSHESzMg4yofzthIkNrzm5KLKkzf+/NX2glM+HAuCwkfzqhD1og7
e9PhgKFFnk7i6RvkVsA5SEw78p3sEQsZQM/GSjZpFV+pG7Zo8CSORcZNwLoOtxuF
RBjSJzYaPCch0DfolrkytJmxB0W8Hk61BcZmT0tRs0IgsmVhqb7VkIb6/bYqEcay
7A7Xrjrnuvy0oeUX2EDYSGNDWOz5J2CDTuNUxvbw2VOKxPZRwL/uPcJjWr8tAnN4
dsDgrUZnXxcpKbQDnWS1SgHbu+jI1IMfX39lXMUM22Ph0MbLiPFLHOffMUzhFF4X
Paw3QbHXBV7DjCzthmJxFeJ9wzX9Ep8+HmESY5bTVRGqM7XX6aWhwNVtmlY1mk1K
jJRwBJlJNLS+WY+Z//fzzd935rhg5TspnEAyM5BcUm6Ih3rr7RhtO3BoNn5+eThf
RosVp4/jvNMl0pd/2lRXiYi9n20EIUXGsPq68pe2GlJRaM8/HRgHEc22J53if8Fm
xKWWkMP3a2EMNkrvp/G2Z6wxRhyjXlPpXlzg9PYKKZHnziG9G6D+ACao181xiYQF
KZryWbR57TrTguXA4+vB5O5gIRisYtWCkWjDJI/vZmFEz+d539vs9Konvq2G/VgC
krXiS3M8rp/FLm9raCFDJqELbRW4TcQjrw1FIQy1x9ECNazqigUmROrMWzEMliAP
uYi/QF7Io9HakE4ZsGhxSnYjjLIOhlgdr9nT14JijAPcYcBy9CfSJ8Y903m6DYla
dvXEbh+76GL4PQHaKsCeRBSUKqglavvky16aJA4vBoaD08X786sOGLe2xVGA80Zo
IuGYNnHY2n3Fo3viz8WRLieAQppCjgXm+pIKxZKDZuWvGHIfyI0bcH9WMV8DhIAq
/2GjfPB1grUw1+VZDMSmQw4cJURO3X0CHyjj3gZ2uQXuXe0DJ+JwrCjnvmEq0GVc
WsDneM72HyZn4cU+wdfLy1PtnNmkazuqddTyoI2ZDUzy5WIXsLI3mmG11IvQ058J
9dSoMGbz+JIYefXf5QF4Wz0TyWB31jW3knkb9FmXy0djTJwGS1psKRpdwXf4xoN/
O3CvMi1hA9UZaqe8lE6qhkFFejh4DxCGtyodrLhsncR/EH4k8JJsz7GhNEHvI8kc
lvd9czbaPg30xHj3Hmh/48HoW324eCLic/PE8CQdvKmF+4nP91Cv2qfgSW6DYXQs
WS1gHr40D6PH6IPtOA/1D9b4WrtpF/1KLDb/V5tLt9KbHzm/a9ghYfIT0hVlwrdX
xFFrG2uilOlMfo74qiwkFQ2eQmsHexygpEQI/R0DmtQPrT7fcAXUGM6s+PvqhYv0
EYTd/XQPFAEFwga7mo7eTswXtJarFwaNlns4Om46hVzcSGMXxd0VulQYvdh0hIWE
IC4fOxR/wkREdeZh7LyN/0ZomCUHioUxTF1a/hz1FjTZTLtcnXZ4AoSjTXa5uNu9
egEe50NxmiWTJlyzC0+59jzCTdLaKdCAzCwl7FNaKQo9PwmULj6GHyvnSLDezshI
lE1K+KCkNXmEPtUJQBq9s+sGv8iy9TDlFAYXnbt3vMevp2QB9ldPP0XNRSDWdsl7
UvAzURcx1W3/rxOA/pew9TQYncGs4Ukz5gxei+iRR95dzxXSSW5jmpZT1epbXtSj
nVI7f+8KbNJ3DyO1W5J7+FFWsDQjrxtT+2gb0wmmMbLAwysDLS1B+bU8zoEmzhiE
aqSWa0fxU6toFm7bezUQDWsuA5z+EpTOIykR3graqqIywBEWiKB02JFWKbmblp2u
6gGTDPfH57Ubq6m5Ar8QoZIntIErIQaQRaEJ+Wwv2ubqB4heIXek/vNroJ1cZuPu
nZevTeQgsYDgOY+F011nOaeJ4XycU9mRESk02drn5HGm9DGmcMaWIpfwIEpmV/OJ
fwHQPlA8e+ZRryVH5qthrxqMBqWYuz+8y0j+aO4wSqA2ioqquMDCaZ9JCIPyKtLl
Zi8b3u7gvO4r1p+Yw/SQ+y0pv+42cewovtQTs3RnJek0q0H3O/u3vAcqGd9Jdf7P
jGJRt8sesDT2iEPJWXXxip3VIP+PLPHLvrK5VaQapIwr2sDdumSedc9HGFEsDkxe
e2HeCXnFlzIf7kCs0kcklvQ7GPTfgda586I6cnssPix2o36xixSrM2X+XQRXNm1P
LL+b9frcispR3Mhz5ZLTXCpRdM2J1QPobTn/QTz2xKIF8F/j0U+qJed/XS/40Jja
iALiko+4xBE2kCewMMSKZEWOnewYoxOyWvXDEO4zvZOH8nmwX2no1Uiuwx/PWZm7
+lCXmqyx2iMrHXIMO95p8v/Rtdurfo6GIl/5FcEDu0YBnzeCxbFdxVdz/laRg0dz
kptmupSYK5vs38CSKlqfvP25DZXX7gqHwLkZYcdZx8V483KmBfF+NfHs4aepHCge
/vH8u0dkzmPJXL1I77xf6kTXngU7QZvJiwyFHLBQhOMx+ODE8f7XdojUerdK02h6
RIzzpJb1Xu0YNZCcXegDhc/5TInLJTffVR8hzLF9Fwi+LqE7y1DRGPw6vdy7+a2j
eks4SFE7Q95Y22Xx/UPra93ICEmGuU1rv6s1G51W7QEBHjkJiv3iob1wqlu/OvCB
S7qaOnO/5cxjZW25pS1h/TTK75sRkL4CbH+8kW/2uEQJbdNYAmFl/ZLxj3cfwTEo
uI++WomHJg+/CP/2wjdNqR1SYEKe4e6aBqPVhcFMlt0JmVa2TWPp99RY+mmBPPpW
f97Vi64oTeg+Hk7Smxevceg5k1PqQnP3eaROzuI7bN666dIVQtq6YeMl2+h3jdq1
jJil4yDN8FMLv24R8oIUeqIV6o2KxjDS+KFD7a10kaDBK+7piFV1+gFK7Slr9mkY
9iIE+ovWm2gDVopFiRWrqvmwYuBHQshGFPF6PgXC768eErnQS4CQEL8mRLDjAHbm
wVnfS8UjUJ8dht8J82a4qLyT++6VuFjKJfjo8RPAv5O1oAaz0ZmEowPdbLpFnIg8
0y4MnFyrd4gADq/qKSJeXvCrjjYQkZopxgxY/zIRo3UJ6xOSyT8tMW/yqKQyLCX2
XRRw+CR8rIAWun7m1a2Z58WZX6GXDsEH2TW24EZz8IfFGTVmC2ZaCmP6enj8jQYO
BsA1hGYEE/OSjlfi8tarM2xnxTojE2QTUO1KU3Ql81sCvaHlbseU+QewP3IklPqI
RT3mBeIxh3MrZMcV7e728gs3TiwISGoLjXW0F3QYO/QYr1tLbU7oiE2Cme+TgMaM
eJm612uKC6D8BMxF0PceMtEkLn+XCTAHHKVJFZDiE1N6j8vc86ULNg+78atuE3lw
CRxsvTQhiwh0NbQtMJLkhwaxw2aKU9ZuDj+Y0Wq/iF+TD7I+r7c+99EyVE7Iiohi
ziBN6JoT2XSaQ0jkfy1h9KnYL2MPC6aokIlYsH4D+O2yZWt//S3eGBM4aEu28JJX
njLlTQs3x4o4Df17ieSABXVOyIjqKFRPSJx0OrfOsY9hIofgDh8KiXvsGFIdnRIc
gAP5VrjUi04xbUsbgAYwB+UbPHcbfTjjdTbIF0fY+C6PADmrEXeeZgJvoPyfezT6
cpQNqeevljjv2tiE6DDqh0MMmSVNIwEDoxGHz1xB+B6V68NJcteOTS95ve37475y
inxhnyp3LwAOt5UCW2MkJLPW/ok4DTiYTXNTvo1QyKFod0jw6rmAD3SEp5n9EuZ5
NyAQdeCscWvCimTpe/qJ2V2gaot0pTNA1cRjo9xQMlpui73BZyOC+Mp/Sl4O9JD4
sB6S1Eg6j8/SZQuqiyZXXgvDGTF56UwEoUv9uov3Gj4OeTeiEP/hM8IQwJDb4abX
dQN5XWZs1vTJI/YYPWX29m5KZ8PvYT7EvR+Jne0J2tN2U6CJvYC9FsVBRT16E9dB
fbzk+BzJvY/sE+kKA7JLO2/RYm6HTnqoPIyAC2C6e8OAfz6sSJ/tWpEpPSP/nSdz
THIQ8lZ6SpFyokXtNBRFHIE8Rt7OU8dLY4O++A0yC9XqXTZV1HPR83ZXEvSGhBjd
vNCEBfE8uudNWkqh9+Duf2NVOniA3NXRklRFsSY/EmYYjM0zPHuHtj/Punb22wyd
v+ZuxOdsZbxCIrMp8W/jWfXjohGSlmBUa78icYsfzwyBkwZWZGGZN9TsvGyyxGyR
gmasZa/8KVN7+N6yc0DqHl9MmBGCD/gbVcekyiQk9meXjQp7z2GfPfblCf9iygVn
XPbB9JNFOgmi0QHIZmxurP4UO4bMvf4x9319W7TkyWQHig6noOIMRJE7R9X0k/k0
QcvlvGu4s6OGd23rTY7BWtgyHukcsjJL0dW6sJuaEyxwF8mycUYlMoh8R/QEAwyv
FxbE1U8GWR0Dvja2LQLvq4Pa/beW5gHhod+kWElh62afiA0EjApwvMBqkTaG5s12
tomsi48PfdUZI2QQyHv1f5rmDuBn2Gkw0bORkQcMWF+l95JWdsoo9nws7N+GFDBs
YTXzvoqRF8Bjh5nsdyglrlnNIe3cj1QYlipwIqyu/Oaxx8fPQWRMLWe5FA91zifI
FWTbRH5vjIljy3MTVnKsRtJO0RuMjhSOZL0A3nnSwyZVd60GaDXf4VY5rNITd9vK
S1SEvIrwjgGzH73yVpc3RZyUbruikHixmd3nRTfDpiuyLjrA81pc68x7LXUs8az0
3QmJqcOOuQfeh36S6TIZI5wFQ4ed6+xykZd+UhIF8Z736JrMMhxxf3T4psVZx1Sh
zTCRNstZ5OjJsfiWe+JFcXnwsK4nU3ZGBhAFM0MqdKEFkGDRLI6zLh0gM4PV89LZ
S+oJmSvsANvd66vOr/fvRUzAcdn7HGLFx7vAVfMQty8LyG6Uk0tE4axpoey7pH7W
j5huLcTxOC9BntoUNJfVMCu+iIxjZGZ+rBJ2LTXuJFnlUG8mtTk0fcmkHEAjhUWn
LXsOV3ORtaHZAm1hjBpyh1goqXVtEwf6nhdW48PNmmZ+BkT/UVfWWeN1DNk8Sh5B
ZJSk41Te/+M6VemJJWpDbhLzcpnq/m3idHWO0YX4ocqXMgRECYTiKeRockST74/j
J71gNGF8Gjjf9OXq78jTYwCr1rVl33R2NJuupvFI7rUxQDSUqTDzDPs1tKkRtJD4
bZvyKwRvsYPw7b+e4hSZYm9BnGJvb1hVb+l1gNRbreiG5lmWuqjSVgyz9Zs/etWM
gzpgQAxowR3jIRWdqZJzX9Jav+j2ub+sdteYKWbnnjzANt+NytNekK45pIuTeuAs
NXWVKW/FXPh6AtahUc/7YMkAeq8tC0JL/VCq6m9+cthdEYG/M/IIzhFuIY8RVpaq
HuRUmBEBZSRnQLHXOTI8Hx9GN6Pq+XuXtXL+4zU+EeoUg1DADZVkYSkfE1PlknmL
t6YG4GlPMPuymiXBWN8WWuSSCUleF8djvKlwpwdFlfTlRx0rMDq1sOXLGo8ozgrx
lDjn/Xh0c/WWK9XeU38Xg/rH29OU5EFOWDLOEoR+d/8Q+KZMw6/1QjUiSjAiFAWd
9NruFJZl9I+mCc2gbocQbyVDS3GCcOkSPk7h3aTDxux0vBEjRhMOu4qfQ2JJDKHn
eISFICRXCdPGO+EzZkHzBT5vrh2MMAvyVjKdZ5u6yWYS19Yn5BwemeJHLSW0Dww2
YiJ7XebVrAS0TsPovunmIKaXUeyNaI+CaEAfhMPtaust/2kff87rloyzjwMh3O8C
I7GgSNm1EsIJ8D1stK6JYm1ESLIrpgDBdEUcbXiMzFJRrBGnRi3+BCvKhuqRWgaa
2vtkVOQlRy1KyFxgImxm8mueArqckbRNZjBQOH1yIeYDIPe4KsFG8drPuRUlJpHf
AxQkpgjpgJk5cOP7/88Qu6qFUH4iBOmrnr5KGFc0MVsoQappkzERwPEYxPFLe9pg
8x2ouBzZEjiTjvYHONYJGy3TINLHT6AeKVj9H/wILCA7jOsdKNWWmaniYs3WgNwt
X+7xVeZUUxud25VBg5WLiHhXyFXI9lh5bIhkYtyrn+4HKuk1lNYb97AN35GT9QfG
/RQiwZ3nS5mEvtlBadp2sO2dlEzHWrHymMtVDnp7ZPHB79JtfbbQ7QGh8TXGhl50
3NuvjrSWT1285cM727ZxcXwM6ArwskAKovGPJS7P34/tt8C9oCCl1AXaqAzM4K9O
TxvnqVkZBGFYllmF8horwwk38S+Bc7MSc+4h8dz0H36NvzVSDknBBHQIdFOsvERD
64NmNbhvSDqMJXOmngtw3f2D849/bZiGhH6wUr+OhN2WZ164j9UBpJNOgX95nvem
8XqzsHOTCqE/HyFzJhJteE/cybLlazFVGj7UUvgIu0j1vouczLtlKRfIzd3/IMd/
pGW9rKMV6a423z9uLosCDQ6+pEOkKz4IHWybRlELNGPihFm8N3F0oEufEt4jKo0m
H8K4P/5clksycTl0sn4k+4ZRZIwBPsMTOz28ae3tOvwzzA9HbV/F8Q7LqPfcL/IY
8WfWdy0A+QP2sE8RRwflDK6V4KtmzMfjj0lDgcJQZMz2kZSUdBJeZLJFOPi8Tbgj
PXBk+Q4pvEvsTDh5LCkBAHU1UoVdVM5wEXoman28kS1006zUHfYLF2bfr/PfjbB3
DceR43CI5dfkhqvmUrMqyosetV1qGXYNj9i+OAFUV8u97o2NIrkjzhWJGiNimnfr
9Z0GUK+qeHiPSyRNyP8Tg5471d12eZ2l+A7z18ZZtG5BD0n4drSwJvozgTf7s7jg
Pm7A4L/ZEIaw85kyXI6EMbw7ir94q4/BorASX9xr03pJ6FGFj1fOFy5QnCGOkBHl
DpUX1f9DcBRIA4jTiyVIzuHtR8jpxyrNBfJzxXPbRlsuEi7ZPN7opc1xQbtg26nr
5bM0z76zft6bH+FLu6pb19t9NjxJGtS8kmU1hwbHfQPjQwlejZU9zZNCB/KmNjl0
3X5A9jwtWqCR4MFy3x0DDsgZoO4TWBM4+jVDzWmDYD1auuM31xtOZzj9OjWkZDUO
pbMKGR3I2P744tMDG51TvyoRsBpJYxdAP8UkA2h0UGby0fhKV8pk2F2fRCS3sqEq
Y2JfzXWiV/xOZCEBJSS4pO0+06E3BCdM1BFnyT++en2WoXsOXP+GWfzVsQbCqMz6
zR7SO7PndZ64bha+8/agvFirWteeLy7U5awqjIPgKSpX5+smX1onTSy61YMlgjKn
rcJwD/UyGhqeR2htuaFX3vtv7X4/mrTOMBCnPPoSjH5pPQAO8utszLAn5ZPOzjVs
8hpAZmerzlEkbeCi6/HOBtO+8D789PrwCCM8cHCsXEWitbwmxcrj+MXlYMuLjjw0
tXkVmW6nINW1zvJJ3nVgb8Nm7dJlHvQ/w+prWbYzPr8iU6pRs26pwld0oVSgbGeo
Th6CJj2FrPF4bgqwEFIGcOGejGMI9ipRHDs5BUuARwmI776yfChMOj/CDDE/LyJs
hPaJ81bMRXhjdTfTZW/SPIamcwiQBT9E6vIGu48/mybPSxq5zNIDxMgkuDgoQN6v
mpmh6Xd9LrMU5QFUCZYeCzP7fa8Z/3EG519NCRE0i56r6sy+l7ARlR/hbyLMw7ru
BmG7ZrAZmzPu8YD6RqsBc7CtXTf6RyOiIlA2WMupeseu8g/s2boKSYKnnhNi3EKs
2BX/oSA9+V/dMahJaexPheniT5RuEYph9BginXE0tmqVWNXtosYWJUYuLpZ7Fwkr
QwpShiKVMiHEUt6nSUQ6is6yxnYNjuj3PH7Jf4ng7/MZn3Tbm7e6fQtzhLSMFx5c
bSRf9y7RNXk3Gkr7NanfcCUIlgkB0XD6jhK3XVGiyhg5PJH3tZMoBpdL0grJsMTK
R81kN6f1ONSh/xZDpb8tdXSC+BDiGv+s+vnT+xkGJi+tryUQ+3Fem9xXPiD1PnT+
DD5rVll3y1oVd5xl8WpiWOxHwQk1Dn7y+42m3TyFT1cd+YmjQoN/1NxE680n20OY
hl+21tyJ1VvsQG13uofK6CZslSAECa5GqQWc0vU+ZfzCM8sp2+9GrYReNjEl2swS
oP8EH1AyELLzbTjRv+NzxP06xCwI8pNA0+/wCMviLSfRHgyyqKV0JZ6e3t7WKyIP
kW7fGGWQXB8hM1ylVbiqJha96enX6W47lvI+kvmzds9ZdLS9rrKB6YSYBifpqlEE
nYmlIEshS6EfkS1PgHT2WdHSB+rgfvkedMvAs6uQfzxELRl92tKcm//cg7uASHn2
zflL0sqnhX3mdXQ8BNrIlWjiVRl4mqUIqvHfx2XwfSlj0Ol+txlYDb4zBMs4O6Oj
eoqS5y+Ywlg/9QYpF4Xr+zx28MSlc60eKfmQMnxHX7uSh5RCncKQ7PWVaBQKcIS0
OpsXFO6OgSDsQiFD3giVSAJKlNoDsAb6SKYp+58sEqToOxLCGbsthazXK8yC58Gb
0+MYuo5o0sKeLufbAjKM1crFPy9mRG9G+SNytgPsZIJL+dOrlJDpU9jf0EkFmV7e
tW7tgU8Iz2l2YAu/67KfaoHB5wAOX/TguUHnFUL5i0ArGNxPma4tU6/HQAnfaqSQ
fYjRiTewFsR4IiP+yAkakdGaIa2J8V6QgK7/PSSjuYSx6T+xF6ACha/xOVMvYarW
Gypa2StIcYUCcqnerRu+XmqqMQFJ8ukoTWHOyezj0s7d1usZg/amEN4+mdftRigZ
bW3mOWF3xLQ7s5BQW1p2i5otE5DG1AGoLf3WvIiXhR1cdic0QAZxMcpBLV0ctob6
xiJOkSmY7mpBhqghmDVmHUHQJzWYH33zuv/IYosqQKjCzfUgzyBOd9hOkFMCeq0J
cSV2UQZHVHGqDcmNVJDI2X9yOiTxDnDorcsaD6772PK2hZglR0mxFtpRYOZdzZhy
YmYMqSpSyCRmFLSZF+cyG0YIawOHnSCeODG/S08FyahtrMqhcN4wt8dDNVzmHvUd
dq6qGnbQiAuBIqX8DRfFtyoI6MTCzGOexGuekvbl/hbsbxwL0jRhEg3ttVvjLXgb
+4soo8rcwXyd8UwfnXYLXo7Ayn6UCM7U8GelGzKram3yUfKDzrtqY9t8QxTPmTsy
uI+45JGoeBtjyF4Ue1aTm6Vyn2m0nu7sso/0wAsdxLu9YAExVtuEsHSxrZKPVgoI
ilt/ohD0ibvv2mQ41PtV+5TrHIyskntgk2Lp55o1dDrpgbRFt/OGky3L9/hWJiJD
u8iNYafUmxT3RjcfIAElUNoJN3XyeU4ruQCYELvtDFrqcoCkLWa/1RWkMOhtVCyB
QktL2y8OgT8MmN2+Tb9/MXgMVtDBinw3AMCob6gK4Z/7vQLxHA4NIyFWVV3ZKopo
FZT6JskqYiduqvUfnPzCB8I7O0boIjZZY9ESSYhAladk8EkZj3GPnoV5NBtCNGPd
GACPAP28GbWssUePGvURVbeS2KlGyvM1sF8fBpJqz5br2+otqxtwWZmlxZBUJmqF
9bK+rbX+RYA8lLf3HwD1/ZW6+1fPCSmxP3ywA1U4ub7uCEywqMggay+2+zT9RD8S
XLqqCtTfJjbS+ijw4zTg1HYg8C0PlQXanEhOAXpV1aWMEr3mO/c/4AjhhVAkF9hM
OVuMQGjFSGdtYTHocExfMf4d1rDpXZqHs5HDiXAs80kLq3sJMllLGnl+eD8MXS0o
plGW/zF5cGzl4plZr24wJnuWjxdUJYXUW9Fk944eiuakk85p/6rsCrFb58vhT7N/
iNUfdX6/wAp7suDxi4XRNzFsoMfBeEAJU6//n84IcDtSdTVGeuI3vV/aHPsVdiad
OCK6h3eJm7W4IOYR6mTso4NtOKf0amXw+wwukku7spXsWYl1Ivi/WVshGFe6cZGQ
VnpvAQ/h7rKo3e4O8ZQNA2GSTAllsoxQnrdyAI5kskpqA5NcTWKLJCfvq5LpSWWQ
jmX+2slqztAL0DkzflAGJNdeI7PM5dg4BZp406qXUVI30BlMn8gytTRa6UMl5ayt
riVuWza4XaFV/mdw7EPBh7xKHfw5brgOvlirPDuOsxPJHAGIUB84YvSWQByZoQMn
qRFOEOdVv+QWNQuOT8AOjYEsnZI91F3d/JWazQ665JNh5F0r571JojE5nq8kpC5y
vehctaKuB3gClOMioVlhsNuDajTRz3bXv+dNB+XUnurnPd4jPtWGjxGgxU6qa1jH
K4RpZih+XdcGbTPinV9lqqA9YUQ2HfSmJKehs288fjqCa5bv1kh5wxkcBa4ulKYF
IULMQjMjX3Jn+fhGUWDU0JmLNXmLGxef7BieFd+avSOqldEUVh6X/IvX6piylYCR
P46H1luakR4i+EONg+lq9O8BZHZY4fubIk673dgqn61vWfkuFH7F3y71MFSDjaDZ
uQ5JaOK0annJylpGr7c9L97nUPNcPXYGYdDChNVXMNN8dxfnaCsX5bofGICxWybY
8kbtA+IIAGSg2juT4f2ng8NU5ST888dMc5iw7c6RZMfrImFS/fC3jsnYqlJB3TRc
YKg0EntrJgLkXji1XWtKzAA5dhkkxFVIhwOo6NRDwFytfNa/Hthu6uyCMKGGgtTM
rEk273LbAcQLfKEIitS7dL1PweRhK1eBLWX7nF/Vd4BpsA7wFHYAgLwX3cCqY6mH
QAf9LwRc3FiO9dmQcsT7VfEsdGpjpTxLcpomFVBoefiRfeQqNFYLDU610x/a13Uo
V1TbO0D3R8lJlJ5pKdSKXNFzOCHGTDnwW+c+Sql5s6riXd/x9OnZ6EvbqFNGPVBV
tatAkNkUiWo42vt5qAEC2xzZK9sU4GTdvNBuVi2iqHUeW28vyMJ6YsOnxMZiCNRM
iaVBF9KGFWCUbB3mBrmqb+xMi/C/aXH0B6icruSTVMXiAbxovHwgMgTSs/iQt8S2
sYu95d1zwY3SV013nXWqp+3GJ4JD7USJYMQd4HW3xTrTJgpqk8Yf19C1wW9DqPGJ
oTperufoDoOaArZx/5VQhO7Lbt3KQO3sI6dZxiymLfcCYkyu+uV94YJgTV76Ngrp
jQS/VntIJ49ckDxkDgMh53+EJDZHZNScSX+SJHGPeSI7qt836hLycBKyzAVP88/6
7Hth2eLzC1O4JFGpHy8ZsWyXZSUTwj+b/kIscBXzzANdNZh1uWGBNcxuXulJr9o4
+RIOY2Q5GPXF+baILqIXQa4zd3hbb5EIw9IUbgI4XPJMyKBcbsVyUW+jQXSXIHLG
8+kXcRhgYOVEkSxwUy2+p8NZ4f2Azr5kEh/SE2Fh9lpsygjklNltFSIhkzSlv6Hr
ZGvz5lCY4cXF5mIdU0FXsy/HwMZpVYYckEYqRHv537DXsDRDx026I/HpGvEN55bV
RTqoZEMn4SG22eQSGBWJJHfSxr1Mjr+9zVPIW4U85NVhhzH9MLqNNgZRzu3Kyq1j
9UBeBGybrXBdGcCflizt8F1t7xnVOqEYcIJQZIjoW65SAHyV31U8Wu0I+ov3KXk0
GZp0HIbFKNR2TMO7Yf0Ies5v3IcIQsEuizUOkEOJQ2QtyTbjV+rgV5s6KcaHxo82
4kzuB3up+X1m/LdC7sowqEgdrBz+MR9NzqL3N1Gum6/aTk6aims5v02Tsikcovx7
SOCeqYFyQfTtGOZXjbf3NDiWr3zgCpahavEr5tiUjb4IS4+hzi0G1I+9ZxTpv5/q
t21JRcDBDNpbvV2WQX8DHncKlkKSs4YNzP+IB4uxlplzO9ODBT6ia+3kDmckq+ZW
jDV2vot5dlmJJQeFs0Fuxds/JlbhH7wU7139t/xxAqMG2B/BNAcVlmKC29PZgxFi
jYxlRyRX9xtcvFl+HpUO7wM9M4Epp8E6LXE9fh5iNvRkTQAlP7K2Aj7maBZMiIym
RdV6BObdw86MdHEGdxUVE1OtH2khBXXolFTT6RTeFekEHaokFqvFwwB2fo9fyZ7O
ijotbuIKDjki3gfAzcPulFQtGgQvgjl5lPPHJVmhWaE2RgQb//rt0xY2U/mAR6v4
AeZI0DcjDAdtC+vJ9BFmmIxUvDv8DvZMftgJOZ4+vebcWgWl242kXI9EV7CRITHP
UQ5ONTfHKqQajXjx9qFSU5Hr3Lb1fCxIrI3M/uNZHqEb1aFrztqf+sU7VykY3Q+c
9MWKdIObORZZi56ebm5Z/9dNhwejyzQinOkX4m0bng5HxdWrC2SFUPWgjgn39OiP
lgWg/ZSsEZJYhjjnkN7akm0hTGjckngtrxCGBVuT3LWef2g8OwSr4n0GnHf01a0/
ElMm9b5e1nEKHTmBfwAxRvkR5d0gk3ekAgC8AoHhFfTdzJf5su43vPuMXbfYeiVO
H5ijMNz/sRqLk+oo4f8kn9dJlkgtyQnWGtHXmwy8Qp97CyWRBqIPqErx3H7P+E58
Iute9dxOv2XPecmxRULGpBf1ZYLUctTwgWp0yqzfkpF1nFgT6gF5YNIgTfjbcQgn
Ehvn40V0XvIkOO+gd1HahRJXgVd3WxikF5cFn0/g+i2nnAF5phXrvZHuTG8Z+8eX
Z3gsnpT+/NHeEMpfQ4okSdkf/4cmfoMDHBrQuDvpGSBuO/WZMNu1cAisBiitPwKv
QxSllbIYXiftorEJGtiF+L8MF4Qa7UiYI1f0Dtpdx3mEcBGThG33VBmg96U57WNY
XDeoxyyi06RwCLk7uu/kzuXPkxgYi1vIZJnXXr+dUcUSvMcSj/CZor+4IWSK/CtX
jgRgfQR9993K+RmiiAfHDWCFkULQ5TofhCHRX43E1B/aadWtxk3AW+CKsrzZ4Qk8
4T7II1SV8fcwdou8tCZ3kw3Xr1OfIbw0pP6noCEW4DDBYkRDdlGfRAQWf4pD0K6Z
jJ5juU7Fzhc4Ozxen0ebQjW970XJV/0iTeVnNGRYW9pFwrUn5H1gBTxZOveRr38Z
hzJ4HZp72LVSzDNTdyN9YiPDZocL9yb1Fr7NdqGTE+pWDV5kJFzPtXNVGEfanUkq
KSgSrCZdK26AYqEQs5yC8WicvZtk8lwKPZ1nW2mzjUlaeI9uHjYEerAYOL0bqSzL
hsYAxSMgi+gA5YTTuSVZ4KjPBF5/TDCy5+N2G8bx1MsuIHgfWAIuk3f1tWyTh5HZ
/wdqFD6en7yry7ZD7nEHBvb0X2DyucFY4FDR6jzlR4Hr8lE/nnT9rZ6hRv85JNvk
QIM12j/KcnKbBsi1ADrzVyy0/1qHH1OeaGphGa5bWzJU38VP1HhucP7/Obzo0djb
c/4kU5adDP7ZXtDGMZrritVVkwx7euUPXZh9AnDbQkbkI1a4GZUHBYNpKaHslt1W
T3uUboUedOc28t0uNaxBXhaS30zWn45yyAEe8yZfkvJ45O7tL4IzgZoN0sIJzbG9
PA75/tw1yqcQgVSG5knUKkaZE5cRF3umwuD9Hu0ynkCFswQD6TxxGTqysmDMCBPu
K/lEjl/XnHLOMye7N97knVZiqV+NzMT2XnN1JAysHMqkngWU4atHKZEtZ/cDY2+M
C6rNow+3h97/E6BZ6Tb4joRffRknYTKuQ3M3VpFcVbTmVrEgLJ5NWj2TuwoSHA+D
j6Jvuy34Ue/NTNXBYSJqOdi8mpJ+KkZ9f/3vhxyz9TEvejlFwwEwZP/JM4OCobIq
/pErB40iBxI2pL/vfTrG6DP3KHiV0zIM4r2Yv3tO+HO0UIBLvsQrhV4VJ6dhTn7x
vuE2MWyvVYcM/J8vSgJz6n/jIb/VRRZ1upbysahtjL/hTTmtKG1BD4PSOevrCt0o
m0o4iQ8Gk/HK8QamI/6t/R/fhKXKO+VH2fNEYVxsbfmN5oV+3rrkBcmUkrsc4DZi
amxvN9wClDtNw3eBztdFm48LFcFDcdDoUqh54KNEmx2G3iZ3kKbYfOMDHbr3ky0h
n9yfQLv+DXYDt8Sn7V7Cxf+Ih6ffHCizY1mJqRo3ZBULXjG2oKxOB4uUE3wrTo+N
KceJjsqlcSohxqYQtN8FUbOueTKZYsrP1VcP5p01Hn9w+MwHjUQBZwfKy/8XH5oU
41B5Bxvx07TRcweV7pM3Ng2QrigoaFA7+bNB8TgU+51uweNKdIsqgqukhJ4/LuNZ
XwmukVpzxzbXDjxAyAyN2tpb+Hwp0iG44gfsizOqpunjsIGNA3xCsIA7DOufdXio
ADJJdtSoXW+MbVBE8gOcJMkNhY2r1Z3ALJsLzGu/tbxTVfQz88DeKrSmYjyJ9Q9H
2UEeaNX79Z0VWGIvGRWofkFOzGXQNqMzlEe7ErJPzBrjoX0uOzZc/lS0xdDzr/r0
uaY5UCScgFppXLvO4F9DjvWaLjdLxjdN1lfOGONdmnM5iKJ5faDe/m+KTIH2xn3p
mqHfQ05498ODZsHE/L7034gm4mbXaruuh1s7J+KrqkQYTfh9W0dm5eXKsi48ELJi
WWpeJJNzQwkh+zzxThL+yDq09pSq33Yg9kmOKfps4kEO6RXFJ0GyIcN9RJAmPo/+
B5ikH6PurvY+xTzCHE5rFMadqqxNVap2qTLeBSqoczm9sY48SnDtCltX8Z5tlcw2
g7LTvFpEF9UJ7ouyjfTqFJ8T6RHsCIWO/bPs88Ov+j3z9pFgVdWhMIxKvg74Yjpo
7yVNk3Uto7rCi9aYE1e4LMFFmHS5pGFQstk3cjNGJqtl3T8I6Fkyx2nxh30R7k8m
Cz53CplqlPm0a2HSNyvtU3tnYgbTbp4tHtkBQ4rN8aSSlFdfAmpFXqd6gvOEW3W2
/QzITOwhfgrOqVN7M9jqeYPm44heTBi5ZBIZi+cJRGfR2pglOJ0gOMEx0LH+k8o3
MSsN/eFWfClhAVieeLGpuKE7e1jHH9xIlo4scfo/EOdNH7CBOhx8Td6IUWxwd7Tb
N4NJOxBiowvQ5sbSxWIyTBIwgeB4V21Rf2hWGunTPEih61KuuDdQ/F3BPErhAGkX
Bz/rd6EoNUBuEQdpsNRlwJ5xP02MORSwoKVGi+JAIfpgsjY6iMNWx5mlDI3lkDfv
EnTaZBnUi9RKg2yroBYsph721YQT33c8o99T1ZvLVTtT+8V4fzabpuR6yIqaqVX4
t3jQn9hbDOynqKKG32tp5Q1idi7/y/gGymJ6s3OshyQRmTvrKcJI0e20L9of44he
WNzqmt+FbO6csXBoIA5NYdaWKqaud3064JjF7TlBewhzJcM/L7QDHux9Wx/Z3jif
bhNISJs7iQO04VkoHkEHZsIzbIR5rTYveNyTrf/uY2I/2hvExj7jwr0qU9Al/d6V
o1wlXYlNYqbB1BBTBas48Q3Wr1FctBl34/KFe8Q0fWZv3sHtTOf2IlMU1yoNcHMt
eq37LKOsTYiyzce8PAXOZhaH2kPuC3fdrmsL3OWm0jyHpPF83jH7rmKJKaTScYFQ
hMFWA/rECz/uTLJBj4fuX8ATdL0zR6rvz7rtsP9LMzOhPTTIrr3aUAzJAynd+/0x
0hitsoQRQEK7gII1DzcFmwZa7oZ9RG82SIimqdi57fcb8voNugQMVIViN7gajBGm
fdEbBz38KRXgUHb4ZBjnolSinGgCDbBtLu5RraxEEndtQQ0zp38RLleWaH10rAMk
yLbHkO7Hp9EW8SwxzppdW3FPKzH3/ysxI3flanDYLdUIMF4TapIfCixLkS8WRgCz
ZjntNTNXjcT150k7AIduPkMLD+628DDhlIXAlMTdvfMudo2XJkt++T5qAEtPFfVI
3w2Bx9YI9NP67797LSfZLhRdC4vPDhdthmxtEzz8rvFNrgKtW7WqCXVhFwboFqWH
uT6xm27MOGIDseGVrBQHfmHW2BeQIpZCPeU9EJ6hf/anPww3l5sFQ6kD4dslHJ4M
dsDfa55oyY5MYQkSuFErn9pij4DgwctB1cU3WluNKYFG1tNUSnOhDGbl1YxWplWG
i/TcHJySEykPDD78kR7oV5WdUoSKvbwUtWttdh49qfBEDAVPr+JR26ftlrjNN+xB
NkUd2WyMN46i9StWWQvoqDxsRPfZhSksEUVwE/Qn+QA6iifk2KoXtu2qSbsR5cYO
Jx7lm5AsPmmWHX6ZgXLX3ijjo7Px9LM/Ao6G4wmf+EHfLBvMtAk9021uIuHE4oxJ
RfxRwefbQQgI9wY731HL+OuT0ZHiCeI6jKxOiKdBeRAHHLWTD5ICz2f15+aSEUDA
dRDoak3nalNAoAFu44fayqrf6Wbc417nFDnGIgpoPslSviUJ8DhWnynvEAVoCv76
af9ajkNrBRbkW4BTRtDRVVGVQJHWOdacqOUQESTCXJyoL0sarEPcK19UmFqFXuZu
m+B4MUWyAycI8vRUnHeEoUXOpR0g05Dy+Nl0wvICivZ7A4fVWYJRzfyWnM/L4iGZ
hkFs+/jm1bHxZrD5+nypUh8AYWkpb966QxOWKRMxMpxrK87Ooi2OUuxy54QYaj7g
MCk7GxZoSc1LNZl1eGJMCRd4FyzOKLy3VUT1utuqZ5XOup8w6eX+bSeWqMJn8abC
RNtxNxmb+5JRa4SowSYVEMHW6fBO1ZHVYXbzETHAI5SGb+kCnb65OjqUd9CfO3/k
u4ngbAIL6IQhdJPuucsubXRDu55dxIb3PEz6Jqjx4w+qVvkxdO7rURCZ7lgMS9Nf
UpOQOCIp/WDkP08ZeQ6bONr6uoPkHHdFmEc5PCjUkLP7blCIAOPt98PukF4CWIf0
3jKbMo6XGFnFk/ObvuKeeJdAV0zAr7ew7L6at7YDcfPWrBTtkFnO8GoEpOcb8HwR
Qnz6GjO6dkmHPOf8mcVysaE863+uLUk1iZrmHDZwFTV6CKoGjmr7p67lkTF+em36
SYP3gVzmtCqSVylBaqzdo/7la7b1VP4NZH/ykv4lPUPIR4fIYuW2TzcqtKywrhwI
nvbVGLev6oPqaEvxZL1neyE2dqe/J9tDOHqHqWH/bPtwCGuq6hO+ZaoK0njoUYqE
nw+cvTiW4Rw9vX7DTS11F29vcsUxo+Pg8hADPpGx5m22gtFBDdi0i5q9jrEgQ63e
y7Mof0ffEEGxOchGpEWQURkhHLLRj9fCIeJfy1hV8noE1R6LXC7xdTSeNM9JDcPZ
tt3OWIME0h0zK6gk24S65dpf19lyrwDWh17x7hFs/QbU7HnyYZYdw0/lfOP/XW3l
waBa2XUzktvowiJX224C4biiX7Wu39AJeq803RYHrvpLcmnyBkv0DO63du9UvQz4
JaRczmcAfGlA9ZwCg0o9yx50ymCw+6JuTeYOxmPt4iyBDy/H8BFT0ya1j/oHFTjV
puSpHvYZ9rr+bkpK+ZSXP1FyIN0CYdb8Iwba213P7wjAfxaX7ual7RC89igJlNYt
/kUtwamelJeqweMYQm2gna92+bLv5/YkvcBvbDFOxLSCDZe5w3DF9ixro0FoGWhz
7k0CzvfNH3D91dqMZ28c8mdeJLrEV69Z3Uz/VtnSMNM0EA40zkJleCKaAbv8ZwMD
84qGQ5xe5nclbFLMtGI3SqLPFfMcok7+4gqqv0A3pJH/wRqGoO3mqWVYqf32YzVJ
prPB95JSU9qpo3J+3YpyWPP30HfSbsXMmshul8KHZ8Z+kvr8gfk2C5uCLmituuUy
+4rjt93IbgZVTJxrYXsV0JQm2aT5lrk0dZf7Vy02CJIUgauf+JUtjib2UkQ4U25q
kojZCCb2zgeLyb0Oo6dlJnNrOVL4HP1WmCUaeTYLS78woSRruMmasUAsM0TvEq5V
ETatFuaVXahTbYq+M0AGUiM9kRii5guNNqYLFe9esGcr1BFzwnMUQx62v1ySemCu
FFPkiuu9jvoysCiZCSIp+HIicNjY6Qo2tNgJQG0k+Cm5thZNI0xSpxsfsWcuZXEK
+wa9Wki2rLmWFImB+4UTgQ2kDchdMm1f2lo94pZThscHPpjTc9/kmQGb114ymmdC
K9gmmID6KCaRQFx6drsLIUyjJQvN+ygkuYt9Uxoj1Jt445t++3ejTDivSQf32TRT
joAwoH8v2eCoKxUVO6xghzoqoZ00IIiYUAEd+OSu9DaCoIXhjXznz3xLUR4nYrFo
UGJI+G6dRNhPAdLBdyPAbLIWElsDOGUrStfus83FBBGhlrs298TEmJNaxZhzAPIZ
Y/dPDbM1880G174uFWIvJ+hjrd4JQkQntMAwv/mXq+0apOS9U9ZaRw3Dpd0NET7L
/jEJzm7utcRsXwQzKm88GzqP39ThjArkmcavzFLBZJ9alpA8fQac6pZftLf71M5h
dUY/xGgW34kYh2+Jc7rLcacIhXNjYcBKa7voTbT04SQrgAdxxDpNGGhW7CL7lQP1
apJluzxK9KDRigq337Lp0IzsR1u4gF1XchDpeKWocNvts/tJf1YoCbaJspOTOKIS
/A2HkkXVMO/Bd2kqbynTzg8TOmg1q5U5zmTrZFv1fILtRYu6X8povYn3UD4b7hkD
hnPkT/zmGAsBYt7BAgQfcKi0+Lji3XRBcsVbBhmGRyRGmG6EAb64bBxO7rFRPtJg
L0OKsNwW8sOZZLDTu4Sw5RYMz+KDfAQ3T1D/GM5xokJF6dC6VnG6evb/uuBCl3G+
6WDNiYtDVgvfo4zn6fIhcwVQu6jFxp3dfms7TWMcws+WsNxZLVMRVNE4LudKg9O7
joi+EpYBMxJXxT5HRKoHgh7TWHptV9NMqXyYG0xdrqWLigoH5+YZZikpYGDsx5vn
kHFE6c3+yMZKvXr472r0VVhTCik5+4F87Dm++Ke+KpMt22gCxzEGy0ymuVQfYWCu
vzOPQl9hFih/U2gVwPmdYRWVlIT4NXmPfFuI0YsEWICwjZBA6tQQp+Xf8qfWcMnL
aTa0lGGAbNAKKZTHEtBz4+zmrcOED+cKvvr/X9ezSfFcE+k7ey6cJZ2t6ky2DYun
a4rlNTOI0p5XnXx0TEi7sv0p66Vl2CRAJ3iD1FOXLCHvUfSjj5AQ0OwUECCsl4aL
B22lm3j8/4idD/pjCvZRD1xag2Ws5rxxpH5RmOpanswozZQMAU4hXoOlKykcBhn/
Br3gMBVVZL3AD2+lWPxKLS57Z+ea5QjythUQTXfe33DVbNxHF4icK8nGyLnZ3dN8
SweOdKAHkHB1bPUuHjansD8w/FBfXF0ygsHD27KohKS0J8O4fDSOhnX8J31FIqd4
uAGRakIQTxe0Asz2iUZpnn1BNDqRiK2QA294KliR9axg4OYZjpHKvSKwCcEAW/LU
2+HweuSjLnO8rPcqzktsTz7yjdhDkdvFdV7Og2AgqftEam9tKCNeZ+sJKNCoNf0M
BPEkqrk3nQMgXQj8SEHRVq7GE2nNVKoNO2NjNUNNAU1Up52vzZxNjXMrAmC87d8Q
33SbBlYexrgAxiGjN9hOC+9HYrsh7LbMgdUOsODwRGr/XvxshX7Wr6+XCSXbKxXQ
9+1BQ2+v6HPkwXjrIPfbZZ60PsL9FYlEvO4rkqXz5d1YUfVLRsWYVjNTuRMDVSUV
D12xOkYJ6fz+TDRQ8h1BVGv7Hz3jCgd5za269H5mVtWi03s3qgE2W1Rh5wCalpui
RiiIQcYC+j7SIuquzWR8iVmr+1SD8E4htiO0HhchHf04+zShDj0hA2J9fQYLtC/w
ICvC1mVm2KJDOYfe4bBgYU08B+4xEbY3peaoBvDAIc4rMBSFVO4yRh8PZ9RxCNWu
7gTbgCtwgCx/h2/nSBsn+oh1ZFQI5bek12ehxUGaIusJEmta4R0TyCzD/M/90e2a
OA8gXWAtQbpChC3DvJ/AJTMW5hA2AWEoQD120d3BSR17t5+lEjk+Fh++D4NiNR57
Ig6327F+XoH/2A8yyt7rZHu61tfxsqynHqVQoKmvKEtuPBEHZ4yEgjl3ifvA9lB/
GePEf7z9ZMCcDk1F7ApVBdvwdw4yNFwfNvVBTbFoLABk8gJgpp45azZeCwpNpvIt
CJRm9GFhfgAtMpP97k88fIM6au9DUFXAf1pAjAVgCDkDTAxAtQ2hyhNKOJsMGu4x
OiahC2aEitWZJc3q8ll13a29eg3Cv0EyiVPlYH0mvgfRyumdJGbUSoiC920U7wj6
K3sfWL1fotvrdd48L8JI01hDa8YzOGczez097C3HrjBeklSsigcm5RuKNFH3EiRD
KqxJtYtcnxDVPdNy9JZLDiTigz6W7qM+jBrv5DzbdzN1nMTWI0bU1sB/yZFacd04
fNQ9IAT+grYDq49Gxi8Iz7qqKUO8Z99uC+D1ffc9SV/s5Tavh7abraMRcH5WTTSx
QBo6GMlG7CuS6mX4xzT3Ne7i8Yk2y8I2OIKnDcAn+tVftXgL6ULThGBx5Hf5JjCu
vnNjCD+nRYWZPPK6KpAAGUBQXP9hl4HiI0A520VADYWINTQSUmRk9lK+wPVO5ENy
BMTRpg9CCH8VGmSUhbFImpDrJnAm3DUrK8lo1Yc/XwK6aOZcgkXGAYMM/y+r9iVV
65uKP16BrjxnWvzO9xu63hlqOSxJpY5IrST+VChlWrlH913e0Thq2GQ+5k+hyAvD
HUfwPSMWaSOsqgfKm0qHsf4tYcnE/IwkmK0LTNHdDKIrMjrznSSqCuKi8g6WXEMi
+Owdg90uLdg7uj830zsGDc34e3tqSDyA4FkMH7g05KZaPk5vxb5ySF5px3A6X/9G
u4QlJtYCe5A9dVY8bMIbGR8THK8E+fN7/0I8Z0QFCggieEsRwI0BUO0Sw6KrmIDN
EviN4R/pDRljVxLWyaFznONmPPkEtqzlZqciTGucV7J2N39y4xJaC2lRB73FtTzO
DTWTMnYSaVLITlmj8SQq6mqn0QXedLspCX7WbgWEe6bt1FGETsfJ7Fu0gEIMRG/Z
BgL9BMB5+hCzztyP2mRaulHoM8mlz3ufC7JZofACVRp9B++NS5hme8bJb6yUqlDk
ouUS2wQT3K6m+2G6hj4x9FM+9qOyZ7mj4cD+vRTroQnV6harwRSVsDUeJfF/4CPF
sPKYTLAsdRhZ5rIAjseOneiPgA4K3AT6iLzBbDZS3yDAsxvoPhBIHnmYaMn1j8BY
2utNi4xJuxD4IWV5lvOBlP/e+/xc2HjowV7acZJZT/Jue+qN8XyqmYYsga8kZEKA
dedIW62MKwuMRdipvcYfMBw/Z5jRcFCWKBUYw0M8Mc2kQP/CeC7BoNiJfGipBTja
TWZhLE/F5YgqymlqcZ8L35iMpMmO5+OOEwkXIEZfxNKbVMbJ4rNm++5rZLbA/g9z
pcugGcownVIjCQBP6mOlDSjJ4A5MirCAoZdG/ZrSHItKvap5uDFvrDj7fwwTR0aw
FTEOu1fwSHDYyrCeF9KphxkQQKl6zYU9LSQbM2te6mBjlmPgO1nX26tHwe0XkLi9
QrY/uckthGDFHCwPJDZEkTLl6/WW2MNOD8yOTWNl6Xx0tnVZnO6WY19HplGwf1kZ
WFLEMltbrH8xZcYQwHhh8MijG0HXnmBGIyfM9SlBH8Rzx+Zl3g6pmTGtEhOmT2ye
fvVskUmSDs2fAVjf5PmhuJwkI/b2+49RVgKK8x4E8+kSJMZLJ2l+RmvR2rl6GTIU
fQ9ZOcYtf1lC5HDSO1ezszcNJjqdIcln/K3VZwmNuVcP0NGBz8hFlPSsB7DKDmO+
OCGJaPG6jnL7mk1IUMUIAkZQ0CshtSdc7zKD+B1iYSsk4fsuBaKbJUB05zqidgRV
XrofgcSEmHpFPXo98saaVm96K0e+uiE88j+8sRiVCdB9lrqGtu4ixhE8SN91m7z5
bAO26ZCN3NBpFOaygAEdtw3TEJR6NCCBThy5lpqe6tyIpp9liVbqHHfwFFOBU3Rf
kXmq3TFaBaWlMPv7JI8s2FyY94msN1B/RKWu7nirji/ZJUgXa0ZWhCmobfKhDMsX
Pkx60EZ48k9nOZ8+e0Vz1HbsfjSHDfpONF1NJM9BRDTWH5mpl8lHgfrdA0QECUOS
+bljmE4wcq/DmAF6e30aZX8Q6iqplFHbiUJyBGF8bRNWTnY5+roxsG8KFm9anj/3
bwpSqzXllmT26TCTGZbQ1WDUP9jHe6fwsh1BrxevtkCHQ3yZRVJ6M9mqoMANJxP/
j39oYwEdPXGMAgs6nIWK9PCN/x55YyU11BsbH5DqDniOYtM+igjqY/qTEI81hlDJ
nqeprgJ47pIpqfMxjs6sRjQoVsEeFBN9T083IJTqzPB6H9ut5eAOzFPh/+iuN1a6
0PkR6K20C1mBT0dT7XLiGZUbop5j7v/WX2BJWYJx2CPCc9Y1JwGhwJ0uSz9M62XY
DeIjeooLRk6VC9Xh4vRzmvjuunKBvM3gvp20RGPBrIZ28QwRuSfJwXCNXkYaXucn
9jJAALil0Z6o5qrPEJXz+b7ZP8qGav/KAz8M/esRLu4YOg/PWG73pqVuvk+8id6l
vcbVuTXZkuLXAI5IjsEkAYw5W6NL46/2nILTLCSjNMTfAOx0b0wz4uva36jza9W7
DJxWVFmHseNJTTKxx5KOlhudB4UwLFY7JOPkd0CrAeprDvKz6538CRwmWYQ3Y70a
2wiKGwjb/hgoOwEuwoXuSXBgIKCRdoKuiB2M1+AG96tTjU1UOPSFnJ1Gg7jyu2ab
Yi0pu7AGEH0weTKPaqvI4JfHKm4XzRiULgSnx+4lTXGZmV8qDHnBMyVw7hLPz+Hj
YFuQ48BEJU46H1uukXERWmW9rCBHLHDqdvJd431H3W78nq7PAVPatgG2Qv1jcljh
I3sACBxyZL6+aXwWWoUYxoM+cLCjHotlREusA8CdOiXjZapzEnybn1ZBga2nYA4L
ydy3G2qSk8JK2osuDDtjkOXBUbEdDdeYrMOp7bOdALhVxWfs/4vzrDP5wjgWXxy4
7mMfr9xVfGe9b2X4+WWFPD81EfttObgLvNlyjotS68z7oHODV0/GDRfCqRX5Z/lC
2MvV4yvXzdSsH8eysrfI+/hBMgMBoHV7ZkzpqJBUi3eCagu6UAQqs42X5dOYH9aQ
SAh6OAjkedkj8QpksVYl5lJIGEgjwiFxrnIZV1Trnm3oTp1rJSRxSP9jCsQNudrl
qq1CS2m4AF4/edOVQz2GhL1Nj4ciEC3Ao/8kEVD9vDF4JPk6tbAAime5v0BDzjwi
8Q3L9JYhR9vxWLeJsBC8AHTacU3wsKzcV0u/VWN22vytjbO5FJLknMZTEH8a3H56
aA9zDmuHWLr0xni5sQHJ89ODEzHFMh/X2mD0di5WfL2rvfORDzpng3Ugrdw4qHu5
wmgfA8NDVMGbXjWKZv0PjwgG5QnpycgSxGLu0J6s1pQAl7Wmja2iMWRXtgmjJkCq
OROHXgtFrrjuuo42u1+1MY5Vq62Tuqddq0F+rT5k6flAED3uQikMUJdMQiz//3yi
Q2rk2mofrqqTYT1i7lUAnyTR+ghkZRTq68TiFrGXEivbIU53vVwFKERxgPcwVOVs
/yWDUKuHX6R/el4XnMGRLmFrcJJdh+gNRrcG6kbAIczPpJxe88xDz0MdusBBFj9c
f55qHPfSjGcgr75lNimmVGiZ77+Sf5tvvTWHTDbxB3wgQG9ed3TQdrF/nZI5uV2y
7g0W/hPZ7jqF63QuFUKxKHus54ocsiUr8Zqhx5drpxFFJUwbRZB45LPcnwGQrAG1
JhgZ/QXCoB57caNo9e63VHmbchv3KwjQ5vEcoOngT/GTXbjRV/K8qTdvsKDpz2j3
4f4ZeWYwbcpoCcfgbiLjClG2aI7RJXFPZAIr52u8PkfuOUHO0I5F09CttNzxoEaA
CTP2FXgCp5QmoZB2N0S2OLnQrSqPTfS47CbowzxZ6NJxEtRmMreUeKg+wt6y0M/h
EajXVRX1L7pF9uucoF6Ouv7BRJOhpEYlx/8Rz4ae38kftL2DIOux4bAzIWJJmi7H
bsllkv9KDtzk7Ms1Vcdlk4s9TEKfuHsJbTz1kmDP5K8+A3LgGxOnh2AR9QvAL/ns
RXWqLUVhf8fzTsjziL3H7hXTTHEgzu9NOpy8866FP8gPDnATemaspwGOS95+CSWA
hDKvHzSaIzhWyiCDaQzpiXrhRyfb3xetya8dnR6VL4yXroeb5gVqwK/fFxgRgqNa
Axx5auihmeFLplCt6cdsVuDTXmpuTuMY2UeX7BxlSCZ2N8HgbOcVz5oren5qxJOh
bPCEzKMsAHF6ME/Tld1YXSxq65mBc57QK3NDdLpn05vtDElw2j7YaPlgigsV95sA
rY/Jd7Fx9ZYpNAry5ALsgl5kgvlnLc1dpVLgQnf9eifRAMd/RBBhnM0csDQO5H7l
H/eSWkn5PFnAS343NJQnNlCKYGSXWwF/DrH2/zEOzOqaNvDhwYMx/+C+HJQMOVHc
bnikkJIIGPf6PPQHVEd4mCQ/o++Mb4CmHNXHpIajD81r0mTvnPBdsv8J0Sr2tYwV
HVJtxiNQnyBUmoF0mjU3kQ+BZjImoPFG5uihUsY2B8aJzlHz7ZvrAyidslU8pwvX
li58xH4BgnAml4gTCOvtEAwf91RMl7TCs75BHxNiG3r2eWjjs3FqsOLLbmjyeO2N
bGpCDO84iil3WtKTfFmxF2kT4tFqnm3Q6cBibYAmcHL+SWk2ppMJA+6oPtuzOBjs
Ln7z+uuxeuiQCcOFr7iKnH3jWCOY2eXWX0xpk0/icYJjLkvykgQwBCzohHezU9nv
RkNsIKe1GLx8W8hIUn7BR401SMaE2tHDLNUOjzI/RJ+BmCeps01VxAH0OJ0jDeXR
x1H4JELk5EuPlwIh5pjrp6cCBrWLYbxwEDOrrPOAolo3/C7GKWksAvsG2DSVHHOH
vlmWiAL97hzcedeiQZM+mHePyKSfJLuDind9zX5mabdr3HC4xVp8j7jV8QG+PB15
XZ2qv+GBB+gE/ESdDLLW9UHYy+JBUIqQGvDgADCjcWjW9BS5rOTmOz2x7noPhYrt
3wKxxg1d1HrTQ6tKQ/xbzTeAEpPczdyEAujBPEM6U97VcT9rjNJcUyxuizVh8BwW
kjB0pCToS5xM1f9nkvyXTRdgSeqgdE6/WfK4MHN5WzicmXgaKY6xMYr2wjNCZ0oh
wIy3cmWRg/yG1JQcHuBBEp85SoPsBKqgiN6al+XOfy3WPh3N0lP57wC2lyH2+Bhp
OtvrkJ6R3R5HXN6E55s1kgq/KnNvb2JW9dyM0OSlAiW2mmMrcC1JvcnnUsIIe6Sl
Pjz57oU1tXaOJ0fo29spkfmP3iHdyoXG+tkDeCw2Uo1b66NOkGApoZqo8ycJRcOh
oj693jTXDU5V5X1ZMC0xNdKwkAm5YiFk58mrbqiA7VoVKKqnXNbWV1FT8Z9MgtU1
PuK3D5D9nwR6+4f7XR6TXQWSJlAEkXd2xt3U5A3TeK5zOnRh4Eo1H10TCctw/pv/
GtZcG88+NpfwVVXJaLqvlc4gcJdr91MnqD/NyEzyvmTgf2TzzkiXKq4U1nLnOC8k
8ujRlwyiHvn9Gqr1RAe7I3NhAkOfIrxcnXQxTa6EVg0IQgr92XyAUJ+qxO9j8moj
dwM2wu8oTXCHh+IeIOqwIs1cAXVwAxAhRAs5WYbsg5exzOGVfBDm81fiotjQTGDs
N1ZzuzAYjY4RZneWpLLqBEeh5eePWecmhlCyrmeHfSURYP0x9eXa2mfgIdzSV2Aw
/Nc80a+nhV1tDymLlQbEld+ZqGVlBfN0emhC7Jlh79Kli8L2uhCNxwdL1b1p7eq5
hJ3vNRQH7NBP0Pv47rBJQOXtMGG02GNlpggECNW1oabBkvpzCrvdF35Lj2nHuGjS
+agbYhMAlDbfSlyO2gPi0uS5I2MNgaYMbX580KAHhEZO91WF4KOQgnNku5Tm1bR3
9m9NnzKSoqyoYvQYnDebZteaJCCXtzP4SZg63Pveii8Slk3OFWZNSspdQ4zuRO8L
oGT8TEW6FipzaYXiq58AiwZyIfpp4BnJatsJuSAGLm5KAzb5tUEwawAqxvpxUfzt
vFWROPfOv5aMY0kb07t8eu9uPtmZWHrzg8/34wsth4454msuGLRZY7OesN9QEyd4
69hGZdguGsCcB1lieUHLhqlK5eO7mJG8cskKhagw6D7peIU2es+i2JTNOCHD8IhU
ilINESsHtOK0Q3poHYEhxY9z6jFQDviKrK6HMfiv60kXGOYTzgnFqv16TtztNvXG
hA/DpNl/x7W8SQdD6Rpqj1alCUx9ppKvdP4aRucXKJSoo46GNd0UmJQt5+9GsdjD
xFExDd8gv2dk7lk01khkYR3LdSaQhCiOyP1RV2OcG8OEeuMvwQReLrQEa6FdGQCH
tQtCTe79CRYa0gbx6bwaNz4RWf+lqKcFjC0mpsLMWP2z7xoMKy/rpP6a0/J1kNnA
YME0X+he+kE1PWo0UbyJR7TtlZwwkZYYwM68pq+9vnGiMxTWBAL3MgrkbNUfUGYQ
FaUT0gowSu8vnmzb3QItD1ORsLUfLFnaDvlNTiYLetjiT+LvAH1MUrIuwmLGuzCM
Tujg0tEAjcFML4wmQdm8+4E8tlZGs3xlIYjRbWNNw0qpBYNTyfpfT0lIlcjgvgiN
9bUBp6hrR5mjaYugYL67zpuTjy0DptTPpEHgFhBn2j2EhgkUEt7fOErJUIpeDqCT
k52h+uLu0Vp9gieSwMb6TYgH3rN8GCOPgNGbMTVP345+5LZZ+5Jqjret1exOzQRj
ky+w6yWuJEnJNpA66tuztoS+nB+loqj0lzVJlUVoiUoKcYkEyJ4wNzMAppfDszrn
qxIJsPOTxztUKmu9PepH4KIDwUpgiOOkUrjUcg0LRp7anXC/M9YiDjz+bU2pnA06
bFpObSumhYeEzg9o2zkdBdchUxtC9l1ZVUpZ5mqAJX63HUgAniirRoq/cl1EhKmW
NqLQAJRwc/GTlvdEZHYOE121ia+zDjuyQHItB0vIEl5VMUqneU9Nu/VH+DE2o+/G
Viz1Va54vxUt2qj4J8Rnb579FAeea0l0KBh3TN6bu9gkV3LAoTY6s6TJckOG5YmP
tHdamXL2Ya+YajA+Qh0l3lBPus2mdvt1uGyqCLqWPE9h8q9CiPBvlRhL3p6SZrq4
aW2arosyLqRy8vH9EpxIuMNtXurQW3iSRNcTL3QSn4zkJ3pMT6ULza9RkJp/aHiL
oIV0KNZN/dpKEls9ULSKLDLL0jTZCt6wIok+YiwBQwOZwQYgbX/62KH8FyNp9WP4
EREhHFIMRsyqJoGK297e7ppe2FvTkcfOb6PD/osGTs3OD21SkkWLBao7bpyeLNBQ
PakJU0BVFtaC5+Z480HdYr4u9qlz9EeJ5AwrQLot1qsAiLEMp8McMTCGZ3CkWtzV
sCK/s+s5BAIH7x90RoQCLW7OnnfIo1CYoUEOdYyqgZEyBJQlMWJFQeDjE1C5xSGF
+uQAHrg92KJo2SoqUwAPMry3yTv0rhOy8OY46zWuV6wvS+3KKdJvjQhrhNjmQ8gU
qA1LcXPfd97ELbBkva/p0nzsC7Ch+c43UUzynwr24GJYJcY76YwUFpyz2dLzN3Pe
Fnhm9zcMktAuVLufEEFZXtHVMSMZM5LhqVt/ZGDf9aYKQrvfy7inWGG1n0XON8gB
3qjjHbLn0qu+zB62gbkSg8KJQp+XgARmVoJLTW/T7+QWZ3c8xlC34vxjoEBCk09z
jgwntF6QTVY1iALFkujXlkauZP5BwxBEfCmi2g3WLUuea8HLwAFB+crr00FLCE7G
tdi8XG/uS2MhYeX09uxPpBJmhfWS3e++XoInHTuTk3xh78Ecnvjs52RzjgnZgtvG
C/wilrn+SC/92s9R6Yn1KEkKuTLjoWx6Nll5z1ygMBpqkB+mRJf610f3XcEKIT2r
6PCtIr9sdXF+lbHh0agYSYCepieQpsWvgEcTeajzTuq7MUtd5WAtOamaPcI+ZtIc
ULvtC7CRsLMoiZsg2d/uuzQ3WJI+QGb3eMNhgIoWIn5JxNaRmdk7MJa0YNtyv7ic
DZ+5Wqfjrngno5g8Nyk5N1GnN4y0sG0RTviC6s2CJ6aB1M4VbsCz6Od73zjLJgbv
uSnmeJo32mgBbyG5cbBtMDh+MoGiw0qlMpcCfqlV1uRmn7awi6N2AdGSB9b/wMKk
bcXHOnkIVS4O/MlpanD6d4WliBsOrmDUw+FrF56yHVzZo0lKeg+Nz6I+HJ6AkjhD
2IN+ubNn8BgAj+E9BvZCwQHY3v9DBYsSV65v9S/n4AzP93gOB8ROcblwtmxfbWPd
ojdKaTkbo4Cs63SHfkMfTU4GDIhvi3KL86tcWnVPJK/2uqYbHkgRPDLIZaOWu6wQ
DWBERSxRl1xSN5shBFohxhIo9OyPEX5xoKnYC7rCD/C5+/6YDqOfY6b6uAh6ypgX
dMXJhyLJwN6/+tBSSuVFqw3VhLyU9luxsd6/ALrtOiSNvXsZzT5tPPleISyBMOte
69/grYPAxTU06Caju2uwCVS64L20IgoiJ7qXsi/uEalLPgDWLCsyjS1NiZiGnCR+
j+jB/muNMOOQssLBqqs72XNqgrFwoAVBPKhvj2fN85fnIjb0iZoB2LVSnjC2YDtz
zjrxWc9q6pX1j8wKRrT3ZZWwlfZC/ZHOysH5lm7A8I4bNFRfLEroZw5o+H0n6sEb
pVSU94eG48fNU0YaLmmilwrG5gqIPmqrfVUQHRJIxlX/9sgggmo/dRT/kuoeURQo
PRWZuY6W3bqveAEaV7JVKtk3uqlBZMC/fdGFCdHs2sco9tppGDhhTEqM21FQpcC1
Lh5OS+TXyItnxS196K9ruCVwSKoIt0sEDNmjerY1++pxBSZB0MXryibSq6y8CXAh
RHhQd4iL+kQnWOCNdFfM4CjvT+sRB8Lhp/4Z8nsHvY63WsDrEAZwjfufI72qf3OZ
8M0gNVjuAoas9y/3UnUIWrHw6wZEdHhIuMwcXYVRiqGE4rYxYdsOxHTTilVKwxiC
c6SwfBfEfTRq+Hth+gVjV9Zzj6WLQJgJs76L8l6xsilASNj9yod60nFdEMSvnHv2
aKokSk9fPpLcpnHdzOtRIcp/VQi/BICG1yAgPejjVs60XAz3fSd8CglSJg7epMJv
Hb05vJLqFN2KZrdDqhf7WIESdlY89xe4k8psyqWlpCu37oY5hp1VCCovR2M0OdY1
6fzg9WGAu2VDZ4HyJ9ETVxo1bQPcyt3TzB3+eVWPRBN4IPPXFYOyQ2TShfye6WbU
jIWzb+QYniJVF927BfiqulwkFRGuvx3Nw0pcLFd+I6D5azAcEDNlytbPX8/Ch/uE
G6NDQX4KDWUIVnDH4vJrwKIoDn/0KOq7SFFheuPAHCgsN/S6n5ozJjAQi6TZfsJ5
k+FJyy5De/jGYxUsRz/XiOJ8oB4rbLrgkwTMYIE/R/aTcb/mYbH/KUItR7a1wdI9
YbRwrXhYEb3gVgJDu9KWElpDcZXM5kqH4uuA5RVu7BT6JgFlFzF+iWs/cksBfSZ7
KIhVX21QfSR0WCcts4sq6aehG8FFu+12HxWmqMp0LjlhAGo16xNb1JyK20osMtA1
Zwth+MexLEe4V2i6ytdiRDmN00jcoo3krNqNWQRX6JYKJXmxafcCMRj9ruqCbEBt
EoXtweSX3vEqi0A9woHttvKUwIAyKdYS8/daVtl+tSvHQppP5MwA0lV7FEpseNis
Xk9hKELJ02hJkPrbo9cuAJcuP45HYacMRlie8XQjcK/HtcOjltQVpsDroDOK2xiG
RnhX8Q7ef+uFIqfUdP99Zg3d1tpkeKRq054u379WDTmHe4uHEKqobTGXq8O20amC
kAIWewxopptsXaTekco8UEwK3yH70Z6s+PzbPrc/q1oOpqF/JcZgxpMcR6UDbNLl
YTIAP2Z/EyOZNW0TTs05UvgITbhIwU5wDUFj69eRcpGYkpdjnSUTryizIf/aXAvB
yo+/SNs+Mqns/PYwzRsUGst+++xJXubC1uAGX/hjlF0t/AVk9dbRHcj7N5jbDim7
azEgxPsjHyigLuYbr4yd0TPmp4aVroaBt/uDYZAIcjsU5hbv8e/WUjZux67RT4ym
EJPz9P2nu0jEDqyevl4y0T7mqnuSaPtQ4qFcPVHC9VhnURaP7ZK3cGcxGA+bHVUU
sxs397BdQlfFR0xpBjzodJ32tYX6hcl88CK4N4284IHrAXVg7KYhJjmL9N+rBWdM
WKT3IP8lbp7mApLfGMErRXzmucLDHXmEUWp0O1sh8XFnRV6bIdK1dlZSpLkPsPpv
UV3dpopX6VCT9YAPAxvpT324SyY7ImveHbTO8/dUE+i7FYvgKGY1cZ3t3WrVOl6G
kjtG6obeaYCnnbNWE7yXxA7etVeuwlGDeTeIlQL3d3xdCvr6NSuaGVB4U7ebeUMe
vKfWjnCyqh1xCCEnw+HkjVCf2OXhmAgpjEUBu1ROxQ+bV+QBvynl6uF1hAPWOk4z
FFkvGG5whspeI8QzbSKTfnBvUyHp22YmMr4P3T0pzHNA3p0z5grB3yQmP+vfFgg1
JWm9eXX3ZGSJPRd/vg4Ppz2w0u87ndp3y/gzkOg6IKXfYXZBjOQUes2ToC9eYjKI
m0Ew2vwomygRIrIwueFwVkfp8IvjQuGCD+5kcySk1emwrvhymFGYymO3KP1jrdCW
KY2oltV5uD0OsbtTHn71yOyaU/u4HjODxHjXwhXtAmxpKLJ+CODGE3tVPgKBtECU
h3UTQsXIG9v7nhE2zvv+Kc6mvPVHTB18nsEQ0kWt5soKgUxK+YCXg1LtP3mTvzr3
i1OCIptbkMu3wOdzwSYSr/MlWWiAmuk57PWE2suuObBmfO3SWLjBcoJkhnOwI6n4
GDjtUztFTBVF+Rp874EuOtEqZxBmGZAjkhedtzmo1894Al2D4S2/UpIToeYXF8PD
JoHYWuzp0rtH61Sz3SXsH0bDL9+vpXabiwVeWzyMQ4gxuHDRJwNv9WWwoDEgAwBd
7OPN01CJZIZNxtIXfAFFLmZl39a2Jc7aptW8rYVO4uXRq1ifodMhYWafz3p0R/0Q
+KeAse5SpQp+sDw/ro1FeEQHDLce1UU2scf6k7ryY6Xi9aUPat3eOtEY4zD0VTqF
0Y/kCtWkRW9PSIgtSXYl9TOwHbkI81FzUgRP4o8fzV1ZEkTOA5ETzz61niHFZWz3
zvk2OcbnYCDsh4T2suNTdDySNouId7iwDsgq0gjtd7KXzSOG4vUkUMe0h9eNWyEU
M7W5shc1M+WCmfd4y/YZkOLzflYfBcsvbsrTTgwU61nrjJ0+TPpCLvonzkWdAob0
q7rwuaXpvLnIqoeMJd/5UrLkTnFj7X5QdzP4x18e2l4cOeYk8BeuxhrmVRQN/bIq
Mm1Ix34uyfixLMKjyw7Mml2LW9dH+SdTyY4Gpk7UM6H0S/2QlV4E50fd+tdTaCb8
A7A7E9TxYkF63XgX0WybTwnBJLyEH4n6+7G18SFlR3/nahGnDW8TuGft3ubkO542
ZVyGXg/VM9ssKNQGOQSo9CxBQG/o9GA8+NcPwDbJBJ4EWPrANEsYyD1jMAbnIoiF
Aj1HqtmmT/E1GvgTTSGrLR499scqPfFp/ABbDAaQqtMPSRALAoUjWe3KRVZmOqmh
1lNG8LQntWs38CqHvGloPfmp7Hcb4z1SN1kphiLUxLsNSIktJ44GhH8T0LbRb9t0
KpcP7AnYcYVECaMWk8rRKSDykRxwnJaJPQAxat5oePCp4YE+MnlDkGlWd0jffGlR
5jtQOy0PXMbNdqfnW0Ud1Wdvd675V4PM+dhB83+gykzAHbzlP4MwzwcMWEHMJdXX
OZ6LPqrtUlvLW2DKfxlPuxRyhFvXT2JJqPK9O/7JWUEMUNpf0xvu76SVpzt6FG2K
+W/k3ijW0G0GuPseL4hbCsfjUCB6vCLSgSnXhLkjUbIoy7h6VxLkQycOda5PSd/h
q75fLzIaicDo1c0h6LJeHrPOgBrgJ6iFp0umLz/9vKfRn0CB+EnsO238GZJBwzYz
e3zXLqKTt96uO66Rv1GTAKTPKanwvH7CQx2eIIydXHpIVNiB9hCL5px/y4AjZnEj
Tc6czYLoqYtbM3mKeOB+Ypi0JX5DHTF66QiH+9lfhyP4//1r8wbDRStJ+XfqtoLp
UqD71Zdu0pT/eIqgFW9KrWzj5GCkrKBcTlW9LZD0N8JNmvn9ysBgGuUZpdiNqXqu
ehOHBfxQPzQNncAQQ/cEcVTKszGfBygQ+N62JVPZsayT1xQVqTe5rIlzrCAB0tt/
QaQwH6o2PYCHsNEzfpb8dMmZGLdtAKvMNamSIdjQg22OFLCp6IcjsXPvroINBe0e
Zn6DuH2V0wUEuxohcXA37KKRKqZB6sdGGE9rBtqbWekHgRkwQSWZmXR4Ry3SNaZD
edKiZo+lK8NocAY7t2iS8g7TY+U5891qfBEhk7ccGsRwIkXeIoOD/Sr9XA+Vz4k/
9ToOLnop2QCYSDIGjHnNMmwm1YquxPBurRa6NDx9pOdC2iNPOSKpiW5lAOvPfhU8
XUnKHoYR2MfsAPNRldqh1cGHQXWZAAj6g7xEgpzcHLYNp/IwjKJvkb+zo2smmsLc
v/h1eLz73cVwVZCmA86XYSbzWNCGs/qffSxUShk7Mda0t1tmPNQkdqutlwMVLMIN
97kqeARcZL9SYJv6El9pdnNhtoLTaE16tNgmQBa4SWEkN+xCXM1KA3V9uHvIDZ0T
4ly8icwJevsmYQw/HNkr8e9WSBmeCSVW9JjKBzUYjexGX8kRWoXvdz4g3MEs0WBn
t4Nl32HUMUuhhP9iZbHJqnShFUFnsorIgAdZzQ0qDJGEey8SFZdM/t/lAt+Ac+hn
cN9oofgFmrr+NTS/QYVDDtyh5Ke4Du/amRu16GFcTE3/O0AGVeywFpJhBEWzNGhT
m0MBWll4x6BT17+Umny2+ykt9IKwCINhxPnOlN6Hne382Bf1TKGfPpowgFx9zUoy
ag5VgUw6C8zTey6PyvQ/u+soweNlxLduZWtCngLqQdyzNQ7Yn+GAmGVI3OfxfY14
5xOP5fYeituAHsyx9hC42v1NguAEElagE35/rDHm2RhR0Q5zU76urACYOeqPNq6I
GrQ8NTRW0Gj1y2dzQ8+LM7NSNpinR6KDLtr9jeeWj2hgXEoz0+mD3iLCmYGxVKtl
l1CrcdMl9Mu29BD4i5H9oP6u1/UHCqtm2uyTtOJvhFGm9nE5gWisYR2ECU3HgLZT
yQXJ6kxL8b6yjdN0RCmWvZX5U+YG/FxYQTR4F5zPShPkAwyp3FnmGk9QR6Yv3RJM
Sn1FYfJg8wrfnMGkPAEVU4a6e/Jt1WnOwR7s0FBAU+qaTLzXjAtEMgQqvep/sDFp
erSYT89mQSa2oSkoLH3Fj9zNaDNVJhZKMpbnySC+wWW8XxDAjY4bmA87NmkeoOR9
RZ7wp7YS0EDMmQ+s87zxUexcwwjLbPGcC0KaPv1GnGPtkbXHXacAuLQSqWn1S31S
4lu7p2vQrb3vewb5L5hOocnyZTXo9taO/o2zEnspPVbptFWUOK62TVygRNYBYBUs
XeV1MvAmy5KZzSkmWNGFf8c4jdjJx5TqkrvPSMzyZrukL0fxvVBCoXMbxDe4bSwG
5lleFzLZgeB5Cr8M2I1xPmio6knuot0krpqpB8lSPGbFiY1QFw3C1+ceevrRj/tW
8HMIuISkwO7zXeAzUM3pxO+PX3wdlICLeTwJJlbGQwGXRzXUPXmzUvqvnbsF6Csr
`protect END_PROTECTED
