`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/oPrVr2fF8q5ZUrnNc2R1wnH88MovRyAQZOYRDT7oIylx9AO2hx/8EGKPHtk1oxh
ynoo3YF3CL3j++JhhsEWcCWVlHYK4V256oJIT2dRVSLpRQ+9KeIy4aI34YUEB4ss
H0jotqtaanxVMTJcTKTvtW8ZyqfUp6DYvyQgn/Qu7OfRCwLvd+314amdm9tFeygT
Ejo7Kc0pFOVKcLWhQq/WJ+U2yqYd6tVWp9F/YqNcPtH+by59oQN+t/56688a6p6F
ciZbHgQnc1I7nnDavtlJmoDx+VBiYarZF9bthbiwvbK/aGieztZo+lWXy7rEPZCx
woQwxCAswQ8XEG8ZoEKozEKohuDgk/ska0xroBZDTr918Tomwj+OP5W76jKuh4BS
DSlKWHjZj1or0/FwTZg/qG/2SPXzWfx5uMn5pTO6a23eorzyD3GMjaSGPMRQBvCO
mC5r7mk/7CGk+MJmpWEObSUNkI7m/hu4UEOkt06KX8f7g3X9wkXdT/3/u6ZiPzz8
d6jePoz3jitFvFeQS++8mRAc0UiiuLyUAe+r+vsDpnozDtLaTkC9cnyEQIeQqK69
0loYgmZyfNvrQvbyYetGhkRDqj6983S3Kjohf78Zh2hecIosGxYMXrj8DvL8yurk
pzYiOCpdcjSyeuDQ9cmehwn4JdRRl/XF2Jl/phyUcUoCNTxC6uwMQMGxsfWMrgVq
zqjVHCrIPLYkfqMkc47w0MPPDCDQZTRPu6pop/YdLTtNNWLmt171KawyFooCBrf/
1WJ6e4/kiYH+H8qLd5MbfyFAakWmPhef2P2fGCRWnogap+dGb2Wwzd6sqIGYgMyi
IZu8WDB0yfVlSlYszW+uRe6nFpKM3ld1m4nippoucuUnp2xwhwZ6H8DOyFYUIFM7
5hQxvsCpDr0l+pCGVQS0RlVeAQcq8QXGhSyyiPghTspyIpoGoUXGaB0HNJ1xdQmQ
pJkq5mhBN5mgrWwMe5XpFmF/qlFc9ldqJe9xhQzOnFixUcMJ2rxnIZWmYROvLJo/
CYC866Z7WD8Xm65NNSt8ereI7+ko07KWzX1ZV3RQq6G0ikpqtumugJUio8EnGc9j
Y5Xp6g19bSlcvrVNHrhqV861X1GnOZL5jpnIyuSPTmF+og3U4XxTmNNRpcbWomog
HltZsTM0cXu4IUAKNtAAXq+xkmUVpwfVe9thUXM/3U4jftkaVlQ3KWvcfprKPcQr
//uKknmz+APp+bWvfppAsAArVfhgTt8Kq/Jz7Vep4AE=
`protect END_PROTECTED
