`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6Th/jMxlC746AfgduDfEQYZoyqcX4rtCgchRL2X97wrx3kbIHeHgog31dzX1x00
2ThdVXUP60vRSzPcO2Kf/gX1aX7SPTrKC5Fz4mCDeva7TBuGK1yD5d9n9p4BB0s/
mmVUUe8OOxVfIrrxayg76n1nt8sNuvYCENjADLcqXy/sJcpd3t7G1qP7yaIietou
Rrz+ehQGCeg86glxhFFwqE50EW6Lt0y0HGKjfj/pPIitjd8K0FeFMInTnLlCb9OH
t9JTy2tkpyhg+9Pasun/RKf2de77wZvwjI3Cvq3j2h1dpV3VL20ODtRc35YZtz5a
Ler8A02U1Rq9lDHqpQEejC8tJUeYSwhqRREUbMml1zKfHEU/3IpxetUm8m45yPmz
p42vqDe2GD/+QcJvbAd8ZOJfRxs9uz5T3Ovyyj3DKljV6h9KxwbkGHeOGgNyjjE1
xe0Be7WjYqfQXokTEOoG86vBdslMx4TSs1YU/M/mX4wh9/zS9j0xtBeWW+FLIAxM
IiqoRASpBM3jCklWjYUmUnf5P+3oT57oUYNFbNyg/Mtxxc9PViVyjPtnngnHTlsp
3f5bpxpDz1qwqQa2INQc4w==
`protect END_PROTECTED
