`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QikZdV9tAOEeRGyET7fSfzj17Kp16pKrMWwKpunk9rHRX0ehWHPasK7h+wZpzEuz
Oh66t4mjWo/A9dnUqutly7k1Oft75KRVzDtjRwp0rEBe7EZxvPpY2iisDZtZKtAA
hOBwOeOkcDg7Mvypov7ACGp5pHRg3y96B7n3EejyBFckSIkPP7Oh1aGSoLFbSJQv
///GBNV2zqP3g/Zn3XtKCwL6Y6/qF8IV5ZqMLEyah3lY2L7RMKbvbEEYgLxkUBvY
PoiDDvhcOY+CJM40LmB+47O5n8btYMLIG4Tt2mzLMZP00iR245c12JISUln+c4tE
5bnL3svvteAvsJ3Z7Hld8VyhfSvSk5PEjzpn5CjBSFJzvElQCvUBLM/2GcqXIQXh
HkNGblZluIgej0jfR3ZYWmhhuV1+OR8Ae4WIxWPTZlmqg4eINtfVDj9eos9l4Mqi
XreZWHvOsRQxruDroptUHeYBSBitDVnJTuWrxYQDqFScCzOKlOaPlX5FTnF1ME8d
fNDSyYu8KpgxP7YLQ9myYcd374KZw0l1vkb645YLFZeqbKj/mZksPOHxgpXHh/tw
PYcOrgGhLOGXBiJvbDmMTDXmTNGW27sJ1M40Ikr1yNczP5IkeEllpxh5VKebS3Xt
TMV5pn3aopOcbriF0AMXOHWRDvSBePGPY36g+83ajfw=
`protect END_PROTECTED
