library verilog;
use verilog.vl_types.all;
entity twentynm_io_aux is
    generic(
        interface_id    : integer := 0;
        verbose_ioaux   : string  := "false";
        sys_clk_source  : string  := "int_osc_clk";
        sys_clk_div     : integer := 2;
        cal_clk_div     : integer := 6;
        config_hps      : string  := "false";
        config_io_aux_bypass: string  := "false";
        config_power_down: string  := "false";
        config_ram      : vl_logic_vector(37 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        config_spare    : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        nios_code_hex_file: string  := "";
        nios_break_vector_word_addr: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        nios_exception_vector_word_addr: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        nios_reset_vector_word_addr: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        parameter_table_hex_file: string  := "";
        simulation_osc_freq_mhz: real    := 800.000000;
        silicon_rev     : string  := "20nm5es";
        mem_contents    : string  := "";
        mem_contents_valid: string  := "false";
        mem_contents_updated: string  := "false"
    );
    port(
        core_clk        : in     vl_logic;
        core_usr_reset_n: in     vl_logic;
        debug_clk       : in     vl_logic;
        debug_select    : in     vl_logic_vector(3 downto 0);
        mcu_en          : in     vl_logic;
        mode            : in     vl_logic;
        soft_nios_addr  : in     vl_logic_vector(27 downto 0);
        soft_nios_burstcount: in     vl_logic;
        soft_nios_byteenable: in     vl_logic_vector(3 downto 0);
        soft_nios_clk   : in     vl_logic;
        soft_nios_read  : in     vl_logic;
        soft_nios_reset_n: in     vl_logic;
        soft_nios_write : in     vl_logic;
        soft_nios_write_data: in     vl_logic_vector(31 downto 0);
        soft_ram_clk    : in     vl_logic;
        soft_ram_reset_n: in     vl_logic;
        soft_ram_read_data: in     vl_logic_vector(31 downto 0);
        soft_ram_rdata_valid: in     vl_logic;
        soft_ram_waitrequest: in     vl_logic;
        uc_read_data    : in     vl_logic_vector(31 downto 0);
        usrmode         : in     vl_logic;
        vji_cdr_to_the_hard_nios: in     vl_logic;
        vji_ir_in_to_the_hard_nios: in     vl_logic_vector(1 downto 0);
        vji_rti_to_the_hard_nios: in     vl_logic;
        vji_sdr_to_the_hard_nios: in     vl_logic;
        vji_tck_to_the_hard_nios: in     vl_logic;
        vji_tdi_to_the_hard_nios: in     vl_logic;
        vji_udr_to_the_hard_nios: in     vl_logic;
        vji_uir_to_the_hard_nios: in     vl_logic;
        debug_out       : out    vl_logic_vector(21 downto 0);
        soft_nios_read_data: out    vl_logic_vector(31 downto 0);
        soft_nios_read_data_valid: out    vl_logic;
        soft_nios_waitrequest: out    vl_logic;
        soft_ram_addr   : out    vl_logic_vector(15 downto 0);
        soft_ram_burstcount: out    vl_logic;
        soft_ram_byteenable: out    vl_logic_vector(3 downto 0);
        soft_ram_debugaccess: out    vl_logic;
        soft_ram_read   : out    vl_logic;
        soft_ram_rst_n  : out    vl_logic;
        soft_ram_write  : out    vl_logic;
        soft_ram_write_data: out    vl_logic_vector(31 downto 0);
        uc_address      : out    vl_logic_vector(19 downto 0);
        uc_av_bus_clk   : out    vl_logic;
        uc_read         : out    vl_logic;
        uc_write        : out    vl_logic;
        uc_write_data   : out    vl_logic_vector(31 downto 0);
        vji_ir_out_from_the_hard_nios: out    vl_logic_vector(1 downto 0);
        vji_tdo_from_the_hard_nios: out    vl_logic;
        pio_in          : in     vl_logic_vector(7 downto 0);
        pio_out         : out    vl_logic_vector(7 downto 0);
        soft_nios_out_addr: out    vl_logic_vector(27 downto 0);
        soft_nios_out_burstcount: out    vl_logic;
        soft_nios_out_byteenable: out    vl_logic_vector(3 downto 0);
        soft_nios_out_clk: out    vl_logic;
        soft_nios_out_read: out    vl_logic;
        soft_nios_out_reset_n: out    vl_logic;
        soft_nios_out_write: out    vl_logic;
        soft_nios_out_write_data: out    vl_logic_vector(31 downto 0);
        soft_nios_out_read_data: in     vl_logic_vector(31 downto 0);
        soft_nios_out_read_data_valid: in     vl_logic;
        soft_nios_out_waitrequest: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of interface_id : constant is 1;
    attribute mti_svvh_generic_type of verbose_ioaux : constant is 1;
    attribute mti_svvh_generic_type of sys_clk_source : constant is 1;
    attribute mti_svvh_generic_type of sys_clk_div : constant is 1;
    attribute mti_svvh_generic_type of cal_clk_div : constant is 1;
    attribute mti_svvh_generic_type of config_hps : constant is 1;
    attribute mti_svvh_generic_type of config_io_aux_bypass : constant is 1;
    attribute mti_svvh_generic_type of config_power_down : constant is 1;
    attribute mti_svvh_generic_type of config_ram : constant is 2;
    attribute mti_svvh_generic_type of config_spare : constant is 1;
    attribute mti_svvh_generic_type of nios_code_hex_file : constant is 1;
    attribute mti_svvh_generic_type of nios_break_vector_word_addr : constant is 1;
    attribute mti_svvh_generic_type of nios_exception_vector_word_addr : constant is 1;
    attribute mti_svvh_generic_type of nios_reset_vector_word_addr : constant is 1;
    attribute mti_svvh_generic_type of parameter_table_hex_file : constant is 1;
    attribute mti_svvh_generic_type of simulation_osc_freq_mhz : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of mem_contents : constant is 1;
    attribute mti_svvh_generic_type of mem_contents_valid : constant is 1;
    attribute mti_svvh_generic_type of mem_contents_updated : constant is 1;
end twentynm_io_aux;
