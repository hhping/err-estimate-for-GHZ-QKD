`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2Kb0FHSabPQKoYRGtaVGa46mDTo2ppbPDJTjFMPdIrrECOEUQnqG8eTOa6aN3/Q
WNf1Sac3o5/grHsdYxhZBIQcs1Qjp47+w72x9CtbYced36GKHyvBGAMa/yXvyHMI
Go8KqURptjmB796iZff1PDmJ9cr+AbfgA0afHECNmCnV/xOmXDCcwZV+oWSfhvMP
RsHnDiPrgMK1mgPLJC6qE6Fmrdcrmgb4Y0rjrd7NRwXACOO5qnNkKhDr4sU/2bXn
UpuwWAoXlFEeIREqoJch6vJSnkOOFJe8XPCag9hJj682H44AzZWDYDpDY45mB/MF
JbUT4IuhOhg+mgXhLt4zhGDEOgwn7Q0UzQTZeswGW9v0fNUmWXa2JW15h+E4UzVm
SjKX1Zq40OpbLU+pzJKcfDsgaoA6+S7nhr61bREv62qjnlS8UMpRHvVQ/O61OP9q
ZCcFB/Hwd1jUilmca7xD0+WNK33yczt7adn26oZ/DX1cRGVHvcY+31AxwahDSg/z
4G/DsI8j4t4lwdIdmMnETJUrDJebMuUttFgQbOnPzYxENPU2kYrTvroFYcw3KFlD
WqyQ5x0gcuPlEHz3WpYDxMceJPCCWLOugs/tytPLvdtWF65/rsK9GyfCKimvN2yr
l7Ms697eY9b2dzceVuXR7ymbzm5gXkvT2AVIGiOxIaUeoESmGYuLT6bCO7AgK3iV
seF8GOIylvdyu+6fQrgQso3dN+jTgVdY/VDd6gEGirkwOfot22dJcAIaei2zFvdZ
f8RjMR3846Edn+MV+QM7BcXS17vSHgkT0sjiPr69IJeTDazLD3Zlwj+s1QvjTgBK
1zzMWEook5ir+m05o5wfF17JDDOlo/aoCmVuD+/wF8TTB596rwFY+ng+LLeV0ye5
OggKO0FoMq9DOFTZ0UD26yemypbLId6Bb7X0pNLK5YCXYbYI9RXXM8w0ZWT1hq7O
qcWtRcePtHaJHqbsW71961/jqsLPQevwsxUlBEuju57SE9NTYeSsQaEineRZ9wMs
nXVtFkGAEMac7sdylSV4MteZrgPpqx6ywAgWbroSUbcdAqkTvtv785c50NPQyh64
tLOgbfK7tFMBwa14NFgAYh6IMR8EpQV/9ierrqdFsBCQZSRrxUPLE2fk1wQzCO7w
PsRuInuSJCcyGxuoylspdTW+rNBFyny3+GbfwRmYS9/q9sBrbYZVtqnHyU3hXV7p
Ie0pfxdxVwbqkzDPx70BUSOkbqN0pBA1cwZSW+hnNbq0w8YuESER9fpD91Gyo7qu
sE1p5GMn/O8PCLXilM+QQSxQMcIolCddizc/LjhGULvEOI6K2M8RG5UOPYjzkGHD
yCcrqWdQFArefwuKKAWpaLsa48JD35hPHIhrf4GMyLVHQLdoz1UR+1b2r+Oux82P
orNuBx+ytzmfZxkYMkDA+Irkpo8UhO+R7Whwg4p5MKMcXD1feDb54XgwlaUJ8cOR
q63II+qM+vXAK3zG2lE5IZB6W+yH7VlFwab4wWwkoeUnuriNIZoCcDEJrkRH1m2d
v9lm57lUSH74O0vy+Zn9ltO5kAsfQjy5cYZb3Pb4ks5BARTCQyMo11nAYzPg8czv
SDC/U/y42x1vQOPJWeLDNn5OVjOYMzAc2sYWJz8RgX9idO3LbeioEQk6KggziRlg
qJXoiz9O9gLmSXmUDwkrj4EGgCud6ioLDzjtUTemrQRPB4pscy1D330hR6VUUf15
rEZ9D9clpygZ/acg5NKdO4QhvauHmB3hpuFagCdxr2zAwWYXdTEmezxeNtaa9Wb7
svGam6PY0UkuAMZPXPjOhOZGYrSUek+4u1gz+9Umi6i4aXpAxUDgDHMFzrCwzhbI
gWIvVWsk6W9wkJcP2xtO12cnkL12s5vK9oUG4goG+s9UdNeugH7XaS8B9smpXxxc
`protect END_PROTECTED
