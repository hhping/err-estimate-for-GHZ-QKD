`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvebPWonhRKD3XELG8jX0egaPmKvf7UfuuxWP3vW/UGEzMt2j4oFUBEw1s290EUd
W1ipW1lUqggHTfTxTZwVyLnJGiSSGJKw1kNYHqNrWb58HVYxkE4m1/7LntLUvgWh
3dF52ZR+giJERx7jR7fUYE33RXGqAzhL+gC2RgkWtz6VSX81PXoVBsZURls5lIqT
XCVh+2PCq2akZiD6E/Lf9FfYu01miU9ZrO1IsBwMBFss4VZer70R8uG2edt4v3ui
3jLzq2BpUdeJMNvbtHqWm6OeJ8Bgrs6k/EjogbaHNH93MmM+2q+RjnNg1mNbV6vQ
wkkoXuzPHNL4cBwQYtqj3N4hbg/w3coshFL5DNxZMiBO5eDW2nSowHSpnUOcNNGI
I4fetyIH9xKInLQR25eyyLaOKcTmhcENfNAGcm2x2bLKQdNEF2rLlApKa67k4IR9
V5BrJ3y22YMiVbQPqjMC434lyqkV8D7QTI/8oMfPbtWxP6xsrJlNOIAG1RFYw+Ol
XsaZ/nOl0eycCW8hG+kSFGLlmqAslMfoTC5QanM8KsIJuR5bsqCuDI5VUbns9xHU
TooHqQoPA2CZyhQXhQ1jCATXz9sD9iFSNyAj59zc4YSCrZc4HUkvmXXCVnX+Wu3/
u8nvdlwbgrAtnbbAPsMw15Dk9SWubyWxqfAF6B96QwEPqzhFPMSjASWtjHLhynkT
fb2zCXRZ0qlS34wexd0xraTI7A3vY2owqjzV83cIAvstdKDEZ2TqA73U6qwU8Tvt
1Kl1Ct8YpCan81VJgd1TXYENVZNJFjZYge2qiDFV5guD+SYUuDpb8MYWAB/8XKPE
aPuH9J5mFBV2rCJ9otFh+HHx+/30qjjMYOSXOM8VJjUxGPcKstZIM8JiO72+Vibj
uXvkPVm+oKS+vndovZdPYIL6d+mQxR1oEeswK24VqeF7hvdshqT/xgkoJ394Y3+R
9mXG+O237iWeeBgV+IHriudAEV8pDC91E0e/Tm9Dda1WO4aEWLQBrh4toG1VeNUy
h02A5+jKNYoE2a2T9ISvG88ECQTs9oClhfanDkMMrtdnnDMnk4gsR2fDOxcvpB3V
`protect END_PROTECTED
