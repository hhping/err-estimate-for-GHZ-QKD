`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqGIc9cgRbNWYyBeTVYAKAB6Q8fep0Yxkqg1oqYruP6+NW/wcUkwyqoTbdGGx5gm
lbTTLNm3hhejlOeR4oGSI+s18GsQN9vAofuuNEZiB7LOCwe3jkafgCFRP+wR9QLI
4Gae7I80d/xgkeuSyQZGmUVFJNCAdvVHot0EnQZ2qHtZP903valZAUOBv0pTztTv
v8ECiU21XsUZbkca5EapcRuRwSSGhARiy1yn98wBvSVaslFOYqFlKACfregnbPR6
dbhJDsMgcEZZGqDouwCk75rn7WU/wbdmv5wehQ2Nq/Od/rVBO1tz1JFniMmdFT+V
3vStLSwbFP3GiVsNU2zXOeFHO86ps7o/VupV9kEQ5QFpZkXldNO9LM/lAPvEjxqg
2eRkJo4oQCDhZt6n1NWsF2v1c7ZtEZKKz+j2AK5WwK5XG1MmDeiIYFfMRHM2tSQ2
RoIswV4LqSN+67F8KwOsIsa1evT1OC2w9kiDLFXoWOc23VZtL63CVp1KiT5lQhPb
vsjrNkiaUy4IYV5GKs5m2lfuU8uIhjmL0uZI+5EL11D7Sqh1/7+LGVKMVMXhFmK2
qOVSZ6clwaOiqrymtZkgx0xbDVud21+MMkKRQFJFo22qtRDKcapjUCx00SuZoLki
+TPY7ZMV6cVBLiiDsF8/cnB55sNgKxR/6g/JBLeG4FW8cS9zU2MTb5QbJKp8HgK+
yDHTzinV6kpxD9IbJ+UwR1tyi7nMjuiAQZWJ3VOlMALKiUV9L9zzAGRNOnFuMEm2
0eHRDgwgu86J+5MJYrcG4pBMIZz9F6zjkYezVWINHmMONP0S81MhvJSmAbDHOCuh
wtJePUS4MHnVpOG26rpFLdPRTMcK8Pe+4A6E3AqPqZhkcGMGz5QtXiIy1eT8gzz4
pO5oHUN3LYiqPesgmBqlBC1MHveOKWHeUl6tiLIORSWuTXTVZIlfHzh6Hli/WhMI
hzUvjGuiPeuWLNv2N+rHnZffEblMe7Iew2iI0AtSRjRGNZnuXoWD1kHXstLdlnwn
+5H+GWrfZUlc5lH5WPkuEn02/P+eQHNq8V69e6mJUDzghUMpQODWjYOhFOeQL0FR
ClNJJ2fV6V9CXLjvi/EpaqNihmIko8jycLI9hkhXh9tY7hUJpPiyPL7/BtfC2xI+
fl8qiQ8ORbECvw91HdWf7MAob9EHBeFoQ3hGLTZ3HL7fEbbM5JNhgB9l0wbt3x+j
`protect END_PROTECTED
