`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
STuacn0osMq85KRfrDOzhq6s9ktP+MUOiCj0JY7J1YSzP8ZVxpvumthD92hKkP5J
GGgXSZb4BwZq/E+VuhpAKq2hJ0/XFEWmQBgp/cuDODcsu1FrBX9EB+ifV+RwBbeI
Di2lFrl8BYWlJiyu8envh2rPrhFrGGn/2J8I3mxqxlc2qFaMaLPK4fTWS5Tc5l/R
OCMXGIcySNsGbw8btula889ALk0JIjDUP6gli/9h1G1CJY8fvxtp+4nTWmyRnIOu
OUS/X/z49uUzNLTrkYk3pu4KurIVwVU5RgpA1Mc6kc/BOrbs7ndeJMe8m1G5wvXp
z03WSrLa5wZJpzQUElJ0NWbFdXrAGd9/CbPVb+lHRQ68Dq4cbl3gimJ9wxZ4j/po
IasUrTDjFWgtNSkbKmSKPJWnEOgiu0lDwr8p43RJ7aUMtY/aFTnxN3FhItNbfUWC
`protect END_PROTECTED
