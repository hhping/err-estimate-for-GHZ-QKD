`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQ7Kmh74lAzBpiWNjcRkwg9HJt4WtdTP+8urLllX4FK/ryZSpxbmmejpUel+cdEB
wFDXuQ2n62gZH1jtnk3MD6NP8Z18PGT2q2OdGS3FXcNvn8GfxYiO8Du2VW+j52bG
q3YTAz0ix/oRV4wi1Fa9z2ZZggDcpbPOH9gejXVYPRqmNNXglutqfbRC2AOtxJTx
HwR1Mwxojorv/OiHZU9ukriAfti/SHCb9XyIRg6r+QB5nGSIvNeTALyyLHi+lYC6
lhYhCTA3FmpMkT7XrA7z6OZs4x7YqTmTJ/R+rpdL0sNv5kqe++kyWyeuMUrGRRlU
Brcyyov3EqKdvdspETIyVohiVmY3J4zv0nVtRHuLAi8rWrm+KerOcqMBuvZ/oQia
Wgg7+532umHmCU+L0oL0pbOCRJ49XADYOLCHNSKnvEUgewfWJxQ4vh1APcB/tB+H
Y4JB7nap0gy+iqVaUwq42GhQXleajiXcQV38tLFGG4NrwgptpKfA8UujnmrIl+D7
Fh4C3xxQLQiQIG5pZ09cOFQqvZXVj8EQXa+2rME56r9VKZv5c492mdMyICrPA4Bz
evj4WRI9AKYtT1zk17JmqsXIXB2V0lJZrY2WzdXX1UAbOFg5+KYEgfJJS3TNBjJH
86s2SyQHfJLfOle/30c84SyTvr2GdIo2n3bEQr4LGTxeFhMHm1ZpyZjfMWTGQdSe
XLVvRaUJaUMCszOqHX9zhurIVVaGYshxC7eO2AEq2KEw3BF4Ih3m1nfDQsoL9pNP
h7PhIfYK5qknVff0CrKbEHzZ40O30fB0c4B1GI3D8CL/gO9OreJzy6oA3OZ7y25G
oiKvKsG5xLYSCnf4Ts3PYmIElPymDUWVWM3Z3wRZfOAGRFNkMOjt2GaC4NuVoBgV
xmkVj6I88jZmiU1vZdpeaz3vaLX0iaJQNgw5jsV/qTEHDhOlLHc7yUgIvF66uLbv
g+hvY9pV1N6fyX/45IMkCdQYK0VgOgrO7lDQjVUcXG58IvHsgi/zL+ifnhxvOwEV
DZjoznDBO/h9+hCrrN53PCbaeIbJLlepf00/XR0GQRVW2KjTO4hHHfp7uRMD2oyN
qY1Y3ICcuZtl2pR5dij4eSDlX12sqWut3sYhF+URaQsNLYb+9Kcfc3k1U64dJ7Iz
PD5SA3sj4HVTCqJoEbLFb8YPcl7ITaDjz6XBZJExmZ4GKKnTqyq1oZP+RoT7X5EY
ZOIQgEJw95DCnt2jjlwQSDRF+0orHPSA7j3FNAIxoYI8vGJnpwgZd9e51ooCaDng
/rh1vvZ8BSVQlLAfMcM9AY6eL4GEfZ4xYatKaJiKI3IVdk7Y3XFs3eK3TLOy/Q6K
3YsIxRlTXXmIaqiWfVVoL9Uhc4RZxHqf4aDTCTf6UXAX7thmioWzbJHUk54NmSjF
02LL/FJpQtga/MatjbyoGzTkyYwV65Xo6rHrmBEYOAEEENji6CGan7LzwBc16WJs
wRpyTkzuiNfk3vURtrm3nO7nVUPpEZMTAN7tH8g3ylPO9n50OearGCULeIIGg9ft
nLRMuzZwblXnEHoNTzMkUYH0aQsQrvOLoRQ2S7+ZEDBH7u4v92gnl38TnDMTnMaG
yfaHNPBu1n3eNtsKQiqh8HDJy/9uXPLAsO0wDC75FnVBh3N+OLDF6/lq1nbfvmcK
ykOkB/4zfs2N5pKxx/MH1T4TQjqhzWajj8U2Xz9c1YWiLI5+nruto+KWRdW+ufmn
IEdaGHZOKYE8tOB/tqQphpZ+yS9/V3g9W4+CZ6XqQVF4518Ec13rF5LXk3fUKbnk
Qbi7Uhq9Pu+QPjw8Sp8BXVezJTT+nNPpLylRHgEqbs3gb0Q8Q1lcA2zYKghL2RkV
8xLk7B1fBCoQu8u8fHGfHxpY1JIbEGYbqStG4B6MblS16F6SlcBP/cBByTWB5zKt
UfSiUuNpJWHelP/DpJbum850+rewttjhhv6sd6BrPPuXn43KiALCtbBrZmbDjnoR
Fq25iAmwRIHz387xg8Rs8PrnUxgHx3sASmxcOK3Fw+jlakPFeTaEZ4hesJIqsMXk
w3ZNvxYB+ZGog9NmiVQFcQyFZdmt6OTGzkXJqUBW1TiAmNTYBHba1vsReV8Dd5Qq
bOBX/UrD4LfEh6KEspdVDgbbxMQnzpxk8Oc/fjOao4ogShFausa9b1MNk/Jcf65I
nGUSHe4pTRZwBS3xQgMGXPGrBFEoR61wugiukmahiLLcobtHK2+jwHMKn8SfBfIA
uhnhZ0gVO+mwYNQPH7Fe5ZaqTAq19S19w7GImACMsIEnJCGHHcPtCa3QZb5Ie7+1
OLJS9LjrVR0IGXH20vx8rSa85BPNBSqdQsFj4CFZZtrvpfp5gfhcJ/AamG+kYGlZ
2bI08YznTjpLwXwN46yesddbRvePn/NcAuJZH7JIcSjpTLF6qEAb4zk0kzZ8wCat
q9aY5yRlUUBv7eFUY4GeTJdVGsALfUCI1Qr9YrHe+if43nSsUuO7jB/wYkXdFse0
3P9dAdhR4DEpL0eNHhV6wCpCFMuLxvjSgyv4TJWQj2d0wG8wu7k4M5mbKGqxL73F
kba0gFOH+R+VDY0DObnCPcpd02sVOrqCVjSr9XrAUEyI80tmqtUiOj0CXzwb3rYc
rmxpO76WrycN3upoXh+8cFa/b+MZevfmOtCPOg46Vb3ZfwsTFykHCM1gJg5Fdcu9
5RsqcWeX08zX9pnogr6P9KaWrnCsuWLhAdKz1XmKb9F6u2FUuCiTBnyDzjpyE149
69RPZYTixEtJNMJkjdW0xTJvn03TCGsbn1U7JESUILoBWM7XQeAzlSTie/dnzO/m
2JuM/LNEz0O/NN6ZYesR27rsMS5QckJVH5D4qwMbdhtH/m2G/JL4bWZfUnvI2LIt
TjZWLvIODOK6FPXfvllfQ8xxubrQJjKwmc88iiUndMMsg/Hhy6Nf71+3e4JYayRT
5ZXntzqrOIXNxVp3WGXgQiq2NPeUGe55HI6Y6WayU8GxKrMokobzI6AchsQcKKLv
tK6Fk4+dneUxjb7K5TGct876dBOd3S33bsMNq+h/t4900wTihu5x0egy1QmCAL7N
CFd8FUyk2zG5jc5eaefCs0Jya0+ZQgCavGDvPMCw3WBUZQfvMc4jXf2kSZ4ALdpW
mcAhk+JDZDLmuI7fZcODKVu7+wsuL8sah46csT5RZRlwzjEPZCDHqOoP2GSB2Pnd
988bqsngV0GXgGEPWe8c9Mld8yjuUfIVKSpf+EAziu3TWdkrUki5p8qHJC0w5yAF
CXUeWAC9IuV+f2pnk/yrKtotwJ2P20flcDT0b5gE04YpZlTeC8qrZ+CED3F1hBWN
+KZMY70DMKCtwfTBRGKSwg7CXDiUK4OBEuJxfMfbiuqXt6g2l0jHt2nAg7I9L1D9
KAb8dmjzo/8nzZQed7/6adbdY+YRfd0I87bSLR0xNPylfQaArtLcZhFcPk6wR5z+
lXLvDa8aGbtCkolmiK0DYLI0YUwg6KBNZOVjTPXfxPqtQlMG7A3o34zqW906q3X1
1wl67GtM/t+eL4bsth93Fj6nIuBSwBDA1GyELBrTpyLESjBCUonh1Vwpp7vUMxUW
90NIL/OD7jI/pZ0JbjzyIau/FuLpufC78CHxXFMWINR0UB5uBIvgEzKo+lsjhQ/h
DfRQyE5ESWYdtd/dq9wxQ5HX2Ushpbjhc9YWLrwxzkpj0d2AZsh2E5NKd3gp/5iK
2VuIswfdiUcw3vg7z/tjJNJ8zHK+scudjACOBBvBw3qdH/HqeljRU62IL0lGeHgv
UwZnqqLm/YJteunojqfJerqdwJZrHGx0PKQxnLJoJ9jCX17jFlQ099O/l4zbfNmG
rdLlmLcGVrbkhlFXk5fDTHXrFxVqRmKpaBVzTpoNFhZZq0Qjt0hHZ9hjhc79ekQI
PzgR/TcovUuxRg83FIbmvxjBZbRK6c7HidgeOWNRKlSUwCkcgFbxOy6DXIA+ml+2
rYYEg8MDCbqKWG4TVLtRqoC//eHp3ETzYtFYsBaY8ueqfeOU/Oh2LMnn5BluAfSU
QZZ1Ycp+lIkfssz5xfDQGE3+tQ8qrJ+jfvSgeee2/Vl9akjGhlOeuOncCKpZx6Tv
UXu86er6dhgj2POytVA6b9pZmjqLSBpVDNUwl08e0ggM9hXpmcHnWvewhb224Ft5
JwJwFxJE0OnjvqjJsx8t3Kbm8WJgEdOAM5/+Xv33XcWtP/4YZ+mf3UXHLtZUJ0pz
bCsQSWwZeuQ06mURpcVs4RSYoo1YFdO6QvNS7RkY6IdWhYnFjHxMy/mTMcBM2OBU
WnCoj5dXN6a5Mm514t6cM8yl6h2gYreb1cN+vYtBvj5I3XgI6SKm2IqS05GUIqvz
+mSR0FwsoeuIt8W2PPaeZJbRTQ25dEO6BwUh17WGKkMVPvW7zA5iV2jOU1uVLx+D
i/kE1RUc/s/WR+k0OsKhh0Lr5F0rba7RkcnzpXMyAFOGYQnMMXhgfDI/ftEkGjwg
j5WvRk0CUPWSJtQKK7o0zRwvyIOyEwRlD8I1/JhG3QpSphqe4BrUaqLQqy9mo3KU
zXeMi1CQ8mgUQb6/XLUhSBt1r5R6Szja0g2yvZvqUskuVBBsyaOvQ24lpZcYnkJa
GNBY8V/guMHPSc5Yed112LNGVhW0qoAbaDtOxY0ysE5g9A08PyyySDnyDQVGpo4K
YcVxO2eBiBaBDCJgmSFmzfAJwoxo+4QDv+REKB/wpL5v6ac4LFbA61LsGgtoB3/B
fA91DRS3z9Pt/18y4C+9cJk8fWzDD3g/iEAllxTi4Uf2bM8xJZWcaxm8uIQb1c8k
4WvINKhhuTvv1R/5t9NwynXSwkuz7Zr3nmkKmUkj7y1fGJsrTViBEXdO9yTEKAwY
GReqOmmumem/e+HKPSkx9OYYkl/MsBoQy0JLmIW+kHiYkSGWRCzj7f9CuOc59s0Y
V69OPSGX6LAEytYh6CODCyKmNPMUYBKxZ1lv3oG1AGN3rMs0ICS1FAonK+Rc9XJs
LAjYQUoAJoNtTEIysCo55PR3Tsdi+146JdH+fULJ7oO/7g78SAgk6NcwVsQ/qJdU
5sHVj5YdkpdIxRwWM9JnxYaeV1ZcbQP/XXZdPr/Jyh4/AbEmFz6UkquaD0BVKKop
8nd3/Bg6EJipjX7DwLMGdfWsit+Qzh3CApo6UKSE8rFXSWO5uOVReEOQ9eWVaaYu
roCD5fgLvHwXc9nBUTGYtp1EsTQH0xm79jzvjQ9g9ILoYyVr8X785BZPaBV3Xpnc
VmpB/4B6896dRJZUP/BD5urK2+Z2/gtjMEcChS2hBdti3K0ouCapfT+krhG7p+dK
mBQBWEet7O9pqiRChKWyOdKv6AhanVgYMSV8C5TGJG6Q774+TAQL+saHFMPFiRjn
V1ngtWLpBuPdYBjJ+STTHHjGcfYWlmEWMEiAUN32XtcdzUhHWfYNIkb+jd2Opt4C
40aOyshFEnd5dLVYlUHesrzxfxAqy9+e+6gG1oAszUh2ysI1ihEndowXHUsB+gug
dbDZDqqVXV/NyOx6/EF6r0d9y3XaCJeL5vvK2fKl4n5K5dM3QCOcP6d9EFdKqgt4
h/AhZ+t8sQ82MbCaaQidHkRarSdEOdLbVpyYx49YD4TWK8D20ICB4vciYZ5tQVmZ
MFE6NqrKP/18vH5phH0HjDEM5oFVH4M9q4VaCt6MZLdF2FpZ/FIlI6ANfNLxfy8v
izinkNRaM68FPOA1VV+OYDBd6aAEovBiOTc7ZsWb5VEFfpF9+qtSPhrdyDJcx3OI
4T0N9+BfFAjXdcum++8EhL9Nybr7Mw/mxr20DYwukpdfhcq0vOOUj3psZZjJsewW
kpjSY1ZtR3d1Pmzh6JNFaX6jhz2cjtHM+HFYX+oJdKMfj89TO/zYhvRyn/8wqcmM
mA/P4zCLiqXFeGG/IrUCYR2JgafVz2JIjOpAkJZqWonO9b17+XvFGyN6Sd3m8Nfw
AHRiQi7tnfmzNctmFZP5eDi6vB+CPMTQO3ig6wxK4Zkma6qmuWXoVhWI4IduwrX9
8t83NOhaM6l0fOqrxXhJFExntIA9LdmGYmx2tIJ4rD0gRfHtus0nkH7cgH/Tp8ad
nl1Vps78eqskP48mAAE/YFKfzQcc0A3+qjMCt7qFyXON0dwnSSEsr1tCZqPHWepq
MMBUfIZ0EsnugEc6yOJpUezGeOs2rrUV24iQv5CZPcIfuncgwdQXF6QPG1oATWee
iwyL95J2IJRwzl0/Gj4MYYClyfgSn6/LnD+iRFIqOwAZU2Vj8PuTdLjkaswlQsf4
nf0ByMPV0YiapHIeqDAwvq0LclankxnPPlvNEZupAi3AjW6/RcQzgm0G3T4oWk6F
3AjhTfMg05sVCnD7L0c6NKuVgzSnYUD5lwD+2Xx6RGMXXqxI49Cjhmf61QvjY3A1
grzXfXOv/JiFPvUcwP8P4jEFOHrxYVthwDaTQeejOADRii/Jl4pEfWPszPQy9Cnr
ZKd5Ai6gNSGrLhYnm7RaVwLnmgeiNh4joMk++ZenxhALYHGv+pHrbegPZTmnFAnG
GFYvcylIvbyQn6kBBkgMR+rW7V+My6C8Fj2cTGvucUFs6Fuia8avyH+xn3kagHpr
HAKqe2qec70L7sABaVXVPqeJD3e6cLUi4zkZDiGtBe0W5G17vmd8grNvHnRXnqXG
7CC18uGoAriPvtE8UKq+84Xatyb2Fw3rtuXPUGTePJ1aaklwIQ9BkIuAa/zkZaxV
KSJX7pV9aUywvTb7B+j9NCG6+nGKpSwaZBzB1kCXZe63a/SZNKavGYbnNmWCPe5q
FRe8WlWtScQVxvlCoeKowX8RcGNBrB9Bp8FLe52y61FaeIwu/SU1xQiJHK1udqkQ
sFmWrfvRt6zJNFLvfl43KaiV5jcabQPhr4XT3m+4RW/EIdceA0K94T0euUZN8Oei
MgAU+akkyrrkj/YSju/Vimz3nMcBSFf3pbp2MK9xJDo3zEu0IzdMdYqG/00zRvG3
D4G5ioJDxj2VBIc0A1M10WfItMyQLZrP4+YeJPTw8rCw5Xp9Wi3GDx/hGu/t5QFo
7Ztor1vu45FCzTvTkKDnMFNtnBGuXkd4a7S/fFhTR5zPYJzqvWN1XJ/65HHuggiq
wKeuWyN0Z5psTbXXtTvDAbD6g4yVL7bXoRaNuN8YvUWnLO4RRi2W0ajxn8BCXdkB
kKvzyPFNRdmju6ZpzgWiLwvruujNTjRGKsG0MJSc3VEmPxYy5zWgafQ0AVu6XSZw
Svk63Xkac0+XqwGV8GVrBVW6HikDQAYnDy3zc7gGw2qIprY3b91wzaPpfL7ZZJwV
UHBXkdbkTzgvnO9bv531wKD3LgTXfLMrLmaPKsJTDQwHoe63jkMKlHYoZEaM1yly
JAs32FsdX8tfXkNp7ED1UWZJ5WKWKKXOr/HJDqAxVufn0wK77AEsIcG0b4qIq8Hw
WstBRZjXShF+wujIAFIqm7W9cYW4EkcGYxE7UYR57E/Ir8s/aSZJFnrLvqVksar7
jYzwrb2XhJhuS/b6RRVTm1XAAS0WhAs5ICCOeko4r/NfU71i3j6ogqW202vTiaUl
i/NZSEMJ/TpAKqWJGaRf7QLqeAKdwfNhoQuG4wZHRr4Mr/daprW7hwxwBJGGO1X6
dbebyUOGKqyHT/R9idtsKvQodDMK6zmS1N4HDNleVHVtLi3xq9K/91fHiPfmMOXb
c2wg60yuDecOFYlF9NTr42gThaedH7fqoud+xm87mIzARGaZjbaRw/rw5Upo/9dT
445hy/8rf4MfTTyRhN5W4Bf+Vhi6hsV4M3kfS48N4hEyOB5VOj87+byXnlUrC6qu
f2pfudiWyqHEu+2FncGh5VEFJKeeJS2W5bh+0y1Kg2zKATV3b1Ed9zVZieIJosx4
ApgKM1N1JpIGWL/lIU4p/ZJmxeitRVJGZp7uDrYgqTD4xOsu+/BecsuJsuPRv1Zz
0+Pj1FMRjU7Ru40wY4MQ6+BLpSHhIa0kz18m8nfU/YsoO7z1df/osPcEHctaxhGu
WGVyK9RKxeRXrVsoBacxEHigjHGCzSTA3gVGDdfe6xho5tx8JunWEy6kXv0+SfN3
XVT/GdkgzVSxV0G4nE/GojdMxsKNDJaIHBzw49nSG0L36JYWZR9NEYo4NfZIREKg
VdgIKFEoYrNTXrJMcewAfq2a8TJ0PzgCpTLEVVcfcD++YWQrbmGrOsrSDTupYGYm
axpCFYwaToOv8DuJlHWf/K8ja0hZWV59IMf8kWt4NwR3CJE+n5ayWQyMgwre3Fpr
3NBi7+3XQ6JKbII6MZIIUoh24cMXmplWWeE7XTfbPuNhq6KMDS2cpux5UfX5R7ZK
fBlF/+L2FIpiK8e254u7Xtpas9QbilH7CsQHyLIN/QQ3SoQUaWUOVzwL23P6VOJb
QiQTn0IErmwGgAP/RVdxpX0ceQqUh9SG2Fb/blQhpvC44e6nKQ6NWDdwxrluzE2N
IlmbvnsvCL+dXmX1sOfhYdjemnz4Br5vVEyz8DheNhvebxW5tewCIQLsARlCRAJo
vheqA7nq5kA7xOL/SLRKFZffoBXVsy0tV35sor380GQjprdJV3zgsdJodbjsRRhB
Fs5ej2rx0DMUU/h6KfGFnHuMwfZNvULwC8zvCvILU7aIkAofrHVArnZSA7KUSoEe
VovdBAAjmspHfQfPlnPGAlSwYIbtQJwGX3fjkXlMRh/7VUm39Clga0llRcxNMbaD
RDwC771XIF0AW+tW5PFlWxgbW/Q0e/GxhSSfFJ5eYEW7Vzae7LOuuMWesczrQIPT
1OG+RqFHrQa7v92y7AGseL2oUBZ70R/uNtMtkFUfNvYWwbHgwvFnxETA1HdwnsGS
KUVnqvZ8w5kOZGd6aOISyCC9gaIczrZb9DVnseS+mtm05SqVY9m2Wx85b5QpAtql
cQwpTvOd354SXYqXV/4X4kRZO4x2N4De/7OxoHKB9FALFlvbU1qPKfZEM1kYOn+R
rpy6Ql1hK5zCzCkj4LP1mrct4xAPs9OFI9ChdkrNjdPoXG6095C9K5nMFC0RfgxP
hQQDG/oTQXcqnV4M9CFi0VL40yeVryUDw5pCY6ePeXwl5TkMGzIMRNsbuRn08nKG
8LqB4r8cc4Ik+s6AzqE9nE/tdmJO+jEpLJOV0exVKksJbRflE6YVndkoSlhntX6s
6LI2CyRhBd6YkL7st2n8D6x4ay77clm7SuRJWC+MlMZl+PdfDzRTbxAe0JVKl5a6
vo5X0bTweOA5VMIRq1K2o1gXL6bVzbvTiTUF3HfkN0U7RxyceymTRGJrmaGEsjXd
ADM2N90uwjNHFE0/k21tRq8FaCTz2ief09ybsykd1Y0TG9EPSflG+HR4ucK43mYr
119b3mEK2esbreGd/cuxpMwR5nJREV8pN6FcXD9TNLvVP/H+SScKD2+pz7m4vtw2
xRV1bJ0PLJkYCCNcmB8/Yp7jP06GiH1RtDJIj5k8L608hiS6XUy+XAb84eLY28oZ
AIsmSeaoL2dhakLH0VZo6EwDazTUnbXHRd+vnfAxDZs3d3RBumwHpoGGKzy8P9zz
cRtjMBgYEET/PcjcKDQRRr5KNL0tbB/XNk3ArpYnoBAFmnJMzMMCVnRi/IhnEvZ5
T6QrfBauHB9z9b2NxRjnGHcyNqGrZPvv2l/u5Ot/0KiajF6+9kTSByk09/ZoWzft
pK/MVTLT7aA+1Rj2Omm1P68dilAbsvMBBsPnrbrHvmzQr5Y0dQieRuMy5Gql9Ne+
Gt8Xq9qRUWQUju7xyBBjhQerTyNfac4KJ78Ra/t8AqHNDHFRM8D1Pnbx+LOxwI1Q
UH3oMNSrtl0MgEKh2b3l/E2fTt3Bdh52QwS5IuCuLwsyGK39jSWwm1/inlaxNPSQ
hBBk2Tg6EY99TfNv3u5KRi56p8AVzxysABwZh0OvGTFI0Y/Nd2ZdiWPTsFmuQwn3
PqteXmYWQ1GA4ExV/np0isj7NeyAcC/CaD/30AYM9AEjHVIBNe7LXq4dIk3J4e+o
S3NnMGRrqBGuFK48nylEAOEmtqvfI6zEasgJdliDAvxHw8SPLsaTS39s2kO6jwWr
zNxCySgrFhz+iM7UWt/ddC3BTwBCT+1GMTK7oTzatl7xR/GXMae6w4Od3EoEppI7
btCnykFU9fRoF06aE7ko2pERZf7TDFtK8Yd8qndOdk3XQU4poEt7Woi+lG3rcKei
ynzvW1fyCBaczC2jyAtzm5eGaBgmYtoDuDGgFpz8Zg+ewF7sDbLAO7Wi1v+eWYOe
6oP4b3OIKGlzpoCF2YYhq2SA0ITrKNPGjbGopuFfumIaHhCaod+FG7eJFkhNxmU9
d95xyhjNMU+3h7JIMxOXrW5Bacg7pxfz75LUG1qfsZIvt6U/Z8vONK0FfVpBa5Hm
Ca1WCUoWm24FukrhuSVGfxZlvzcZEMsG4Zuk8TQ4ZkQYzs2fW9Vsk86zW4S0W/mD
L51Mhfv5J3c0XO/Zx3xBXsPfA+elUDwQy8zxY0Lq1spmbChW1gtt1D6GAmML3K8a
k5HeCvNrtZxoJOlJ3CUWau45uwf0pBSty9MbXc845wamrP+20TUhhOnP5HpLfEHs
X7xAI0xzli0U+KWsYZ5SAxCBODOkOPL5AZE1BWlZUq1YcTh3CXv8b/C3DVUcT3wq
9C9d9/L51B0j1U6yz60FEk1UPtJXiTTFWwHwkjYHmqqfxE/oM/Kut+r0MbgMQ0D7
DFLjJyGaNDjf9sRvQJj8gqZR/G5DvMoAlVac3Jig+W9tSUt111MtEDJjGjuLc8AF
tDpDF5VaP3z5aUppeqYXtLysnhRfCygrTPfhVOC2qGUkw04Bp04kHDODvdlTQovs
UUBHTf8q8jnudJyiyHOHoiW2mnIJZgg9xH9/csWNarnBReEbwYmaj+Vk3yWM1TIT
LS43VVPA0sqpOoc4vk++tEW2vvDqn5Wsl3kkQCK47ZLq0LOixmhJ7cLnl2u6hbOg
zb0VKG2pgLE8G9ZaTtw5rMltVHINuxPzANXemKDF8prORxlp1biBOjoyvoQ3MhHM
QuH4azQg8m5b+k/HUXVDIBBfstuXP2OThe+f6/y/as1CD2iSutDZs0z3j8uA2HEv
Q8ouzR2/JyjLMoFuuvsrB1g6hE4GmHO6kH/NmzXynjIoLVyKrZ+o5UPS3J5hoofb
Fg9pSrx4l0UAzIdDqiCpDKDC98w1LuW4QGg6pcw6E/Z+CxP8FTcao2aXkLugHTYQ
ymAXB4wQi8J2k98wFFSXgHg8i2IPOdGBl8VHBYLiZyDY2Dxy8uO5ddZTEuML8YGk
ghjGKPuNXy/uvSWcTHOSqG3Ii7SZqE6jVEI9ciO0KBq/jmVlH9PF563yAESbuE6T
uvW08VUzCZKM5Uxth9hyevV5jSkexaJD/AU+Gz054hTrcZ+5VoeN3BtRQaUAKogP
HpbaEfSbC3X31Oh4ylbvyMXBviiCUzSSOmkF4zB4ulsQ7+9cMuTF6QILqi4lOsY+
SZF/EXoH0nbW0Mh7RcHwg5yf+u4c9aOQCdWJXWY/akg0QhRKDIW73qCvih+Ou/h0
z3bEq6DWtGj3LBxsZLlBGKmIOF92vWd4vLanYCqt6q+92+ONQS8x25pOTBo7knHq
RvdyDudrMwcGxM06J7X4AHjF6zcPv4VdCgHQgbjVJnRbzwtS502boWVLaBsrWWTv
hN25LWlp/M54Xt8JG4eCu6d5XyZw6IXRTPenlauG/0Ys4kLRgF/Cq36u5U5K+BTB
U6FCW0woOZ8XZu7B3/Oy7+rhupzZl5ml9rXNcmWkyEAmW/P7vZhaZjgnFED3v8lJ
M0RxR38hi2qdJRFgYlveZ//a2Js6PR9C94z+ZruSuvqsx10msTctdTUMlSw/MXDs
53p/zl1kvzeQAMkAKrU+XHFRayFCgClWXL3/locWTcOfVNSUlrUNRTA4FwnOH+/M
lbO90R3bSTGlHfKh1/QU2D555T53AO/nvZVmP2ij594hi1Ic816UpwnI09N2AYeT
CR5CVMbbo+GdnOZWrrcQ6SXi52KBMa/BH3ooxMowxD3rM3LBUTSlvBMA50/HcSta
ry1ijE4dSvkvj56Zt1sWu1q1fGMFM5edroZ8aRVBnNEge98jQN7l2arQy6K6tnl8
TTQAhnoqOWdBoR5NFrvhX5T9a8oHMxg0+uvjI97A1jKxo4eGg1lsH3n4hPFJUCUr
rkOtetnt0dtueWT/8yVuOt0rIeGGR4/3YYd6Pc5oO5W2JQIJtuRTOfQzgVkXw/Q7
1nbD6+d0TvoaB3I6LMch6UxAXrjjbvoZR2loPoUq59uBwlKfPAdMrZ/W3Kj/3IxX
P8LtDH+sYBrMfvQLfGSyTgA3deiH1C6zrnoiwjLTImBde0rKP0SSM6B8WgxNvy1M
KateTSsWrRfZTMd0yJ7fCUWFXdiKZdfrkiuhJV0VbfKblVZHv/l/2jePzU1Ro/7+
F6NLmAYhDlKZORIsOIaQil+s7ff537Ww4DsMEPue8dvmMKJxWh+gPQJ2U0Tly/k/
y5M29MIDtQtLFUEWPr54ac4R2Sqa7LKU2FF5IVD/OI7TK0/g8w2xpXRf08vm5bN6
Kg1FzWWdmJdyg+QViSlGtP5oYK+zcbQR8JE2o9R+l/LFT+5eTllPMtzJAP0smdfI
vUQiOi7TxiITyovYPbNRu8QCD9WdtcLokxVakZntVpc+ngZrK1uhlm7RXNcHjgXa
/69xHFTwB6Y75Eb9Yt4HfupF6HZuQaD1FsGmSxOcQiZZZm+XVnYfHHW+2gnF42Te
1SkZ8jjEFPwoVLVS8JnyPvjclu2r5Z7Dkq1iGAoWqAZcoketBedJwGdUOHGFoOgH
aJlX3XC9qPtgYIaAkfw4YTq4nxNZ0lqs7AeBN7JhUqgLi5Rb1Uf4OMIySp6hKCMC
LDp2rnfVkN5EGRbxbsmNmxddKJtkP+lOjRIp2cIixxqxBRWE2x5ALlK3VxWF9ydw
XvynmRHzR6Hqh+e29f7/6chaiknjlZEO62QOrjALaP3jAPCkc8Q4ndDTU/5CASZG
fqXLvMY37wlZzXDzk/y8u2w+WsrM8GqOk5xtCBlfG2nDhNQRPKO2UryY1IU/0bSz
h/dUohcmhpDy+cqCDUkJVmE1DZka87ZPABike6vrYUSzx+3Y/3Y9YD4AO2L5Eyo9
4DXNBm0M0+uJZv5UQp/KduXBHKFz0eY4gv950CgsxHCepiYBTBWvlQ3BGxYzRAAD
ndgogtxun4EzsdPG8w8WcsBnk3AJLal1PUz/O74JRHxJQfuweB1PANlaT7SPrFuL
AYmPdsT5WHlI1IaIWYslh+cT3Veg8JFIz0xubY6TvZ4fohuyoDPEOz5dOYs8Ht1b
LULE8u+rVb/E5XgeSK9F3p3wVVsR5UYYxqMwzFHtADtHymid350XOzGZaMrjozjA
OlQo+Lvd++OD+4+AhqSscIUZvQ67sp6r+o3rLUOvojaZAl6Bs6377cDu+RZJDFyt
VCyeCop3es/Mghcupiqdtlk9QVUD9eTj9y0LNPk6FrkO2R/mQq6W8Y0k5mQtCyWB
ovXYtqut3rObpQiaYKczFiRssQo1f8/f+MKRaOcegldM2AXsz59PaljMu0HvOPIZ
kfm+O/FYfZvtYZXpsQr2DOEsKOwCN8nrPjg6UnIv4Fl/axPA9EWm731iRl/wFTBQ
2qcFp097d7Ad4j/FjmlRVTc/3R/dz/2aokWBYwU6rpmgSK7RF/6V9RqpiOhkoPfO
n0JZBHhiHss7TmSzFE/2FwCGc6MawzIVZyoahaL66L1ihWtCSqj2aGItqafhwscP
nR8svI6xCIyW42kzVW7EJLgcBhYtRFJOQBx5J9+AqEiMpjiWWGVjmu7JXxOHbEiO
KSibmbKefN507bwjOJsvkAUbgMyGhuuRMr4xm67RHUJOUFdp2Qn42okAuNlM60of
19HGqlcBlKpxeyhdlKEh42x4bJaTD80h8iPLe+7IUJh9XGip+ObdjtvHGY/Pfbaj
szAyP4BAofuEphMh+F+EGiMk8kF152vYud4zH58FBSXGYNQ+SxyUZzlSU0yqU1yq
IxNDSB3V5mm4YFGkILdTdNQ1rfjPbQyObmxifYy4/YjG3/O/uG1t8sD2Iacz3xXi
UIdE93RCxOz6K9WliYQaAHN3MH5h3YwXLOE1m9EUoLW2ehOolJ46ODZ3/JTaF4J2
exuxcpL4Ihzh05uR3E+T7qpsTceIp1l+G7lvKFcj5BGVUH7I0sj3qCgEtgoY1T95
BVCCGmz9b10JjMhdPkRCzUvNQ27RVUrm32UBHsEmUvuI/7wWvJL1mLc5+SMM6yQw
mC3DukJYWptzrFlDuXi0XryPfwqUozgsafQcsEoowTeCTpdQql7Uoio2O2EQEjgm
FUPJ35owxFtlqfe0I3BE8lZ/SaybMK/L4Kwjo0UOUusWYFsrP9oMOqrI4EnYfP+T
QKvFX8uBZhAPvLdXBA7EY0huAbOZYjElHH8sze5IjglQUna3NaLmPluYbbdl4K4/
VmsChL4gjuJ9F3sRNf4DB+z0sJ0bCunRtxRD/Kf8rxoor4kVM08ugdp0oC6n772i
ez9QRCI+F/QXxIwlbA15VsQZm5TCoyhwQKJfogKWlVeCLWaDwtQKvcOu0YnFn5tC
d/7spjoE5D7nual6IZgfMhKvIhzZQiibEgWX3a/BU2bEyz4Wfw8Oydrk9b+SIijY
n9yTX1bexVI53aL149md9kzYfSuUd20PwQzbbQclyyEHLZ9CCBUN7uGdHx0aFpVq
QRS6VicZBjHDZTJb5grujxdjk6PZviFwQP4Dz+mWypXdJUlTf3TG7kiYvu8zaUvm
Fnb2gABmG6klWBBheea+LWxV8QoZydbg4WCS6zg6q57t1yxHdDhtdySSdFTj2F3a
jqQquJ1clXuJgxmy9E9bGYt2qiMOqnOGJoP7ZQ7ZIBWjdqO8lgq5ozSVlv521K2s
7MRieoK4qsAsQKqiWkmv5EtXnDFgXdh0zpyGKUwvFqIK2+Xa/Jjj0IbUhoD15Jnj
NdARsn1usfDdwhga3DzXLh/AdGH5+I/sPcvp0Cm4TX8b62wZ2kCxIztPDpygSzdK
IdlspwXZoPI2Ajdgoqb2EOxLuW5nY6b18KbFyG0giirF9bK4WIXWXJCrs2mqDDIU
svzCOI0Pb5NjQ0gx1v+vkM7tIogk2CUAtl/yHygmsQ9NZySPnfmy1Jb6NmWU0J2B
2WMcD4MunSXjaDuYI0eNhoq/2qw+PbA13wumE1QpFrPIx8gHyxNl0KTeILQgjfir
XeWJGkyuRRwzUtIN/ff4tTbbgPO+qe99nmWjDKJS4wO+2xLaIt0DVn1kcxMRTpVK
65ATJbC9k079lj67Lb7DSrMjNdewMAtBN0LkPS9KIEHVoiIcCvcsRXiy+YNZC5Hb
u/cQQ3lFY9vVyub1p+rXuOmYHXKnijDNKhoqmjNwtHkZYbxrKX0JWGj8Nst5jmxF
B+t1LwIcczUYOzQ3pT5yahSOnIGBE7d1Lynxb8x/FGGK9nitmS/dxIbHk5kiAHjK
L+XCqSeVJD0TFERCkEN2syMwd2YRAq97yXJCet4bppEA5J7nhhcsVGTLZmdL/oqC
iuKdbacKF8IwB/Vrd3BcgwX2H+f0A2rBZ3hHs2ntgb7EhGh52oajpKGQOVQaOWzO
elLQIzzP368MA3Qj7pHQqU6otTagPrZp8YuF9v6wutMWb/WwNstEs/m77qlEWZcN
3w71AbMb3k/zcTG0bN3T+92V6QrQ3C14UAsoBsbDfmI0kMMuyHen4faCsNB+IySh
VpIghnfCZpc4pHxklVM/icws5+RWSbmqoZqf/TnDDqJcbEKZ+cWYjIQ05/GaukGe
J4tHyTD8LZAuqpyNI2IJPKd/z9XcdiS+N/cWOatDd1sDtlSk23tMUsEcq11/DKVV
YeY8takr8JuQFmS1pxp68Nc5zvt5PXj/MQWY6WTRcmnryTt8F418XMHhrBqYAQwp
iEuymd7FZfKSVWNfC8rG6WpZdkFk+jET0U71YMA0l+z6C0JsqyW3SYZ6RsAIwmVX
ak/6H3rUZsEjdL67T9zsK+uyW5ArjKFDGRYKGmTeCTyaesWN7IPTBYl2v1YqyXnu
adJXciaVd5mFxRN1KDM94O+wx6bYpnb/8Xqn6G2xWW1NhdQ2jg1xFnIT0AOFSbYW
dco+xL+oSTPVLQCT0W7AzrGy+JoQ2NSjiohgB/c7qmYpvgovkrTHOWyrO2bgM6Uu
aU3KYyVr24pVCIfP/G8OWmNcXWgg8ewHKnX7lVQnnwPrABUMs7/M0y9zpswxen3S
04xtwhjmmF3DucU7/aebUOYBgMXnj3ax9+XKol54d+TjD1x9mEx9oQ0dQqodGhtA
a3OjhamkzMOFr3SuRjIdlL9m1Wm3DGZtACm2ClzUu1XRKydLFzinQodlSegQkYNL
TF9JMa9goHyd9ZXS0qInAEItJEhnh/kT+/vv+NTrkmIa9NPaZBjNtfHgNFL9WYMj
4lO4UewZaotZ0NDUsvgHT5wVoitiDmWZFuQAdtnhUygwJ6BzdPiWhMo+gtrhG6SU
pbY0nhOwp0Xz8nIL877nm5vnm/cUlEATxFVGtFkJoV+PLVYGNuSWDLRa/ivHEd8p
97xEOLt0Vzkv9o9r3WOPe+a6TeuE/J3tJdX/ky846J61E48KTT/UHzLNvxfB9H04
u7olXR4dWEwptKK0Z66Vf+2qBavQc6YUud4GjpS+l0Yedf2elO7nyT6FSBalKnS2
EpoWnD3oFtRsL7aihlUoTkjdxiSkaHOyCdt6EOWBNlhiaSpK1Ehhmah63Tr2bmwk
je0x2Zk8oHQHAkB46EOHs7NqIij6Y7660oX7r+rI0zX+54HddfFDfQ+nEHc8wfis
2/Q2177BUNcs2YaFO5s1J5OK0ucW15M10RBEAKQwfMB0ef+NVhJY34cyCGU8ap5o
GN3aUXfkiT+0sxvmrnEsb05Npx6WUqTMFj+wNHFThTWH6566Bfp9dhW7dMSUHLzN
EpPxJSQs47Rg2XBeHFjeLRoosA50+uvbIx2BIUYysIJJUxkL+z6aMopptUCeh4F6
wlScoFygPiQ3EBogmgmydmN+SFq7kwXFjdPzqmAkA7tYfVrqSWM6plQ2CmNX7dcO
x250a2CMS/zOOosu/W53Rgd0bkPIKl3rroHeUv1NOiC9etSaiDPF9Rgui8tTpMi9
cV9srr1SSccd9mqL3XQY++UUMRd8iGKeGruzZ4j8jk0GSkDfDqZUNYtGhrXri70e
t0OY6cZ9Ul5uREHTwyPLqtmWSvPXyHJjqg7Ltc1YNX2cNka8aHGXDk3zt870Fdcc
HsO4LFjkvUL+2pIFstyzD8aGH1vXuDAv8p9wiu2TxPtUhCv7pxI/McOc82QGeRCX
K2sDVQamiKpdW5MXA1IkH7rFhX+CggXzv4Gg0gNZzTduG08+Qx2vzmwHfOZoKnPf
KrEGRr5WODa/PKQ03lr7jRqwaurzAVcsEQygM5cKZfUnylgap4ijMgVOXfdfWgeR
yNxmY7zVTQzJz9KzDALW1Q5SUy0Nz+4aV6x1dvWi3AMvGqyClb5nWbGxfAXSMSZs
Ru/dDLrXzP+ck+1iiXMKnM1O/TgEvYXPsnbTqOPmutqRCVycK4kHjA+M3i/O3OOC
XqJ/7TGwyh5f4qICqaZXPX3Mzd5/2bMFPmPzM0LKkaM0cCoVOgWSZiasAYgdY0FT
csWtqpR10V/P38CGpGFJIBZhtKwWxnW4JN5QSDh9OsJ9WovvtTyy7LiFjIR6ZjsZ
ceonpFcHx31o15mUfG928RD4cMCpsX3B1paTp4BBV8q4/rlNR+rklXW1q8iM0lfl
TkS51hgL5GIPsgcqJ3uE3qsI3+h3nW2vMhq54gpspVoMAwOBiEsa54tJ0VjkKDe3
2PEK/aj3KJ0X55wTBazuFjAtFj9Mz+2Tt+vXjenD0lukbSSL+BUuxo9LDNgPUJa5
IRSK5XyCOHBeTHpFmnvTgj/k88P/fLXpSrKGFAuYN4fJebntfU5k86TfQJjomZJH
U/sy62OVWQin8k/jX4VqiRPg8gORj/uAbUobyTSNnsFm/Yva3j5TTkOTSRdCmPve
Rt26DJ6unTBqwjxddLmrU59ZLeXWAR2LUA9K8iPS9XWOPqEzjysOyjmyS6bo4Wfn
0qh2pzcPRjvbDaBuDytZ7jB2D0ezgdBdQ9LGSUrX9AqtDP94haDYwvv1wHvK5q8x
hn9KKKjDN2DiACalPTI2bltfq0+B25v3VOkRAYwWy6OXJpHMXRjxuNtElkPUa5P4
pZ/88m0B2ZA7FDTxqkg4hod5PQ9hU7OUKlzmunUN+5z8TL3UgG5RPl7+20v0SOM/
ek2mH+fxlxFngcOzYzYeSYZganyWDj9oNHI6RnxxWgswwydqlda0c8TzXh6Ca0Xf
X5vfjxXbDk/ppKLPmsUdGhXuXzF8K+TdtbINUmUnE9b4cGhRxHg7ysnbHBo+Ulev
yFoIdhs13asn/9UqUkUAbGO8o0X9Rm7TpjrmY+O7zzxU8RXc0W0hpGRd0zEgFQdl
2P+4a9f2bMe3woiF/yDQPWwDbvsHOUGxTCDTT+7TJC+QnDhW5CW8Gyaos/l6+Hoe
LKP48GaTXXNERKZwTVOgkDfkQr5qVG4AP85+UAq0WYrtQ0gmFK+FUykXA+h75D8z
02VXeNCTi6Gu5O3ZjeWB9KFCF6TXm9t/GgPk4Y2vRIi8gD9jpNO21daGhJlrZaRP
/7HWooF6z6h+5XjmOchlrF6z61oyHmJHJsHPYKtxyGmJBHsc6ckhsM6XVhf6JPSg
q5bKwybEdGG5+6WzeHnATYypAwEUpLvSjRyTB0PK193TTfr/zLV8YzT70wIF78I6
miKXxFmEPHYHxC32gxCeH3keShD7L4KDLqbvhP6Y6Xd6wyRmmo1CDjk8zIAV3dd5
R8NAHZvYGg80cpSfO3Wa1Ah4kzrIqXk90rBAfcrRF2OVbRYy/KeqXiQl31+8fHxr
hcqph3JnL4L2OmDgaioS+Si7gwZbV/goNQPWT5ZnXura4uGlCqg6oI+LBFR8sndf
9ElMi+TblySKQXq0VgDk97b263gVBQh4OSNBErBPyWlwe9FAE9TYBNGtcMt1XhP1
QfcgraWI4wuoh87WyrLoSJHfAjvV0qZw25vmvkqOT7ZAA6p6v0etc6P95e9Figxi
2Rv3dSZMYdxX7qPMzFoBMKjBaYTwHwTTLVBE1cnIoeIsqtpvZAUhwHbhmn1B1XfD
UMIgezBG1zfo6syZR1awGiIhr0sw0FndICApBq052yVMX4mswy/fm1qpV60cPoEG
i7uyHNWmiTFZNtnY2YWkGlA+7VY9Pzzv8qaVy5luDNTd4ZqdbM9afHbz9cdBgq8R
x02ZWQTm/E4Gu0/arZDWdOGFrdlE7bymE4lpaiIWvILhUcEQFFX29Pw0WF148vlW
Mzjlnvh2SLC/66id2Uh1WN/r1cc2kvSXpx5jY4J/4xg9m5xGg1GIxcFU7fXCRXPU
4o6Sra3s8nEo773kN74YBjme67Aco60EoI+avxGsxRi7LVPLdi6z5E6ELZzbrtK5
TwxtjI/ZnSRZk5D7tQjCxmPnNpzILjBXW7XJLouRp/gj4JuxncbeUfZ70tvbBCQ0
hg8oTYFDnoWRVpruy4i6iLiJFlEt3SvTdRGEnpUF1TT4bOuajUwHwhkFA3j0zVYi
JtPU9wCq8rODeh8Dm49K7WcU2HUnja0ARtwUDlwfcLXRuVi/lMlGd8M1pXWsAw+i
M+xOmDWH3Pt5NlrFGqZD3mFUFJ0QmPxfzw1o+RIbWu9ZmLkp56+AkAjMGXGOkRhL
VJJiNFgwLLPLZNgL01gReXF9WZ4AgoTuANjb7yHp+6tdg8pVy0/n8+JcAq5OXhxd
adpE1dMeZNuk8+Pq4815kC4ErPxo3kb1J94WAzNaFCvtVFaJFqYM/4VyEdtZDI4L
hzSL+6ML3r2YOoqRa8ykHvBIeWgwmEH45zVANdSrsu1gvlnCQaj/K8tUbDmT7t74
tIhmRFwyNT6tJfBTtAatdc7gflkcCQqn33MtSmuocWtJ8tnzeSB+2y44XoLw++5I
d05zrccZ8P1zbJUqm5huqwYvVF576sMBy7PyHWUx/pidAU+INKHz9Pa9Kzco4rgX
et3iwWC+aYOeXVA8oeuQ7IjJrSfis14zWK1tmyP0NQ7DX6IgXT3/Rsj1OIAHLXiW
ENIhA9cc6FCM8YV/xV15AC10yHm3GL7TjmwEtlhfA3gMM1oy3GZds3eKFVKXx7v+
G2crURYVcPJRwzRb0qVjAeFHBjszmDRnzbmCqUUas3TjS6SCi3UA/EEu5iHJeWhq
ICtpqsy+7/JEdfyBodpX8a+xkqurxePbyakCthDjBbEuOkD0z1f0lscU2xyhAg4Q
RNX5LMQJ4GkP6ZoGwjVbkKJ5MF15qzA/UYRLcgQfqEgj3QBZx23MEszMYreBiw1P
Wx7afl7YLzK8aQi8FHsYLt0/kZ4VQoSvJwKOI10mnwTpiyY8fU23MSXh3g7RQ8Vx
bNI4G2AI7ZRFhPDyvNayg7WJsaDntI/lqJkxxeD6UhizCdqplilvUxU3gUey+zLF
s3jwp7kia0sYYhmQN8TvpbKXhBzOxB5DVjOjYL3XNoSB+/cJGN8FJhwgbHdL8O21
qY3C6TrbO7OKsR1m8rQ776NiSdKzlZeIPgu6uVPpiGc8ipcm1tcpXXwJx+Izt5GP
jdHe7bH+H1jk8AfYoojAqk7Xk5CHiPoygv3OdtR78fEGwjyB6ngoChgimnKkMv97
qLSf9tva77H8dWd+JYk4OYP7Qr+unzPI1nyrrcvlm0bIks5rt5BLTtwB/lHfpbtL
Vnbg02p0XR7jjN6lPOWcHTckDNrmJBododS9FOvtoFRKeWkEHgYuII7l2juAS7Cu
sWNL1oPzlqwmAbgXR9z3EUnJna/oXHBQ6KKusdLkWAAtlQ7CVTznd3zfZBDBvYtC
EL2InUFfqV2r+BuTuWd3pZsCwbPH6/zOp3QZkEsywGBe041F2NK/GBKfe6cHKcm+
NsG3QXK/fqlB9kw22k0J9756XLdx8OvVJeGOvf3xVXxAOyLJ5uniDNAAeNCLMtYA
L1RzNRAsA3S80Cvcb4J2BS0fQ5MocY6d8QYGKUIQHncK6fSrxliusyIT0hpGBSm2
Lt/gaecK5sAJFSozwGY4pXFvNSbZL2mrQXIc3krInuniT/UtZNdBsrC7UWfhrelE
1WKPw7HlzsFmOAPePGH0Ois/XPeCS9uT6Ozd4NujNdfsVsun/4jhKpG7EefQjSR/
gD51LZL7PfJsDpZ8+AzSYrOzwwQgMm976+HmwLY0c3rwEnQxfQ5sJIe+cijU3uL/
lxx8inTr8OcC+jh2QeSRgLpbWn8EI8IgA4jB2XqNdJu6+9EwEpL9ZdhDQyh6IniU
iW+dnbrHlaVh19dTgYZ8vvj5qlFTPnhyam2TfmEG9xBO7gKObV2QRzdQkAQwuZL8
VDX0M4LhJKWer0pjQSsHmeALj4XJj0ciyLkE26Q5j0rh6duXStmjp2sPDtqw30+3
sPlaJK2urzJprqGjUAI38BG8BwPoSMS0FPGy0C9J7LfWieqmDJbnp0ZqgLSqC5gj
J03Cp3jHqdCmGBUfpleRkioSVZETwwiiyJyaNem8cfehCyIeOuBae9dKSlMlawiD
QLCtrNp2zIGifbexFD6qfvb7tTNag/8BJr++2AM3xUXjVPcRBWwANjwErD9W+x0t
mgDqQBgmKElGQL22kBh/kOQPUf0nPnhHWMXKzpbgmuxACARZX2pYeeuDiLDVPvz6
uCAYAr+rgCy2hC08wdELWD0FdZURcCkDIt6XSuWBdnVL/WJ1s8NTWq5CfXSloXnR
joqFMsXzEyonZFQGBupoBPtLmHKVeUkJWxG73zA84bDyCycji7Bg8ztw4TiFxVEs
+qYnX7iC2+e69p2gJl5hjWtzrk8Zf07wWzQJP9VsTa62dLhaoenSqf78+1M2+Qj5
pyVM0O6q1ZsmYDLoGWGott5rM6EBYo2zUVs2UA99KHcjDoH8w+OMwuI43U0tr8v2
j0wY4ws2fHejEDKWMKqeQnJPDVHx9ahdvmImA5TTtLlH4zBToVrkvRFuxW3kUtxE
raBkRqcG+MopNorsP44o1UrWYeAYEJl3kRaRdloS2Zbmg8iZTj5f+qqf5glwMU2J
Sr7eXxY0WjLDV2qcy4qisESIl7lVFlTbKYsAjbSqHXc+Ir+jcx4o8OFiGcFApwb5
7k5PjwAV4wuY1XYbqAoRkJB3G8e+fzS4D254mBanoahYtZgT94e6jguMKgzYC2pP
9tdnHqZSY/FKL5eFqSAKf92/OWtMfinUj/zrW8Pj5IuGkpSDzssWsH2fQtc6rw4j
K3PFG1M4QpRa+HG/L8GhAs0tsgTWQZkA0S1tKCbYMKOzrkFnDjYk9izkw06+5Zw0
W84HfUf/65vJyQhcbuawaW+9llxXZhCJU29yYHTvp5D8Pq3Jbn5T2Tdm993OvjVa
A3GuoskjvLkln3JY9io+PD48R+g5b2oZIbUIO8nSZHW/trbiyjJUUP62h3kTa4l5
8kUq7jAiE/LfBCu50GjDIYN9FCBYXaYACdbmMy84fvQxzPDbypwOHszXCvRGqGrU
D5LDSUX0nGXwuM0Nfq35rdmC789nc7LKpv0GM3ZhCTRqW2RoScfnfz4eMoZsok4n
qwUDtC3byXgxcgHbfzGun/ku+O+lOZcRCLMT7VTXTjXljNL6NChJd/zSrX0bdDwT
wj7Vlhgkb1QOBqFrR8AFF/SkIks8AFZsBymtuhz1gXkbxS8l4pE5GgFwb43tO6hw
0XtKbL1FHGP7OUqIf6X22e5PiA0M7YCaugUpkduvg1oZsJyCNN6o4oC2ZPZiQ/2t
1C/aBsMKF6ie/FTXnoCdZmnJhuYoTdTtE9qdCLxWKVBp+0QnxXnugmWgR8C+Vq+8
Mc+iBYrzLIETbuKw5d/4jzrXLwdqHd6LU7aO2gAGVvXrMioNWcuZp2Nw2e4f1N3o
TqddtXLiQ/IO7UYeFy47rxMVDieFDSfvHyzlVTRG9IizlbETLZuCO6iTkBlATJdl
KC1qt9/i9CNJJAEfd0X7Uz4WaLfE+AQObM5pI1W36fvW+7PRZ7ZrcotpmKViAyVw
OWdLLZig3h018QzHSe2Xx6jW7T0XKAWvsH3lzwDM2Iyj0uiTdOWBFDTM213E8gjm
FGDr8Je2R3u02GKq6x6hegWt3aJcI4vm68+LwhKCn+cFh/ARhRSuCKHD7IwmaYKN
jXz1ZJEM0BIOjFofAyBVNsjfl7jkGxNR+0fPbgE5BGbSgPRviOQLEmzOClsc06iq
PsBiJt3MmPVaYtgAe2dG3Nfvi5hNIrIyP0x+GpGUHgE6S9PVTEjt/ETtpd2od6oK
2XpZW7wTzpVS+MpIHV1ESxLNknwhfgRiZpUWbCJ6ce6n/rPwvQwgQryxTEYKH+ed
knowqoyiOFirWwN8W8ru7deph5sdYBla6AX6UQpOgocRfhxTB+EEyZ5IYvWzXADi
zbanGYq7i8aKFAR6D7PHuom9pPUdkOvBEo6f4/PO8c9k2HQmBEj3cZ9qwRg3Dc+Z
UF5oueYEIXUQx36KJhIus8OWx65e7Y4ldos0NaAG63I7UC2gTd8+YiMKfISuUIcN
79CvrohK2oI5gIYxUpeVh2bt0xUCJ3c3o1wUU/gnRToVBb/sfB+89tnvnM1dxok6
o6a/BfbETHH5+i+V8JTprl/k2Jp169zwom7YYJHvV/7pNkSW7of0t0kT1qlo/eRs
iHweph1Iw5vg5OWW8HNfMzhLJIeG1ggmwScYP19Z09JAUjWQsJp1v8xuTQW8KOSw
C8GvYFPsTJGeN2kzZhJ71yAuaq+5Bz0bu4sXzaxPaPZQ1bRGqxXvpcdEDyv1MojM
oSQxqYptjoatNn80aLrVcziq2U6QW/gfyupQOwDj27xVWbY3EAwRXPoyA0Lt2UrC
uxntwG+sSBj4zvfyFrSAOBq+7drQX4zhW0TwSUer89uI1MA1j7OJXBUmnUWOG0JL
v5cL0jFICf8sdCai9yfkvlvPbSuNbuT/YSkIGV5r/0Qe514KbQ/7bWSOn9nYlp/p
4JX9jdJ9UwmylM14xTiYiK/OK8WEkLZjGckdZZaQpIdhY2auCDrFr1av+g0GJ4Ki
8Srd6VeT72NM7ukZr6OKZLdFN1VOWAmRrmPte4fRd505sF1zMHSN6DFYQPptNlp5
FKih/+cfQ4jACSzmQUSB/M2U/9OlbX/kYlGFwpEpoldT/xZ9eZVD0jQurZEOwoNy
Olm6NtPdvzChHC+sPvAMKdJlhUClMNpPlVb450vEdoQOTw+db5c8mhneKQSUarrm
ziv/VADSiEz+8oBCr+r3S2MV/gVP8nT/1ZR3xnGDltPq6IUY0UH9tCkMTjcjXHoh
l/jalFTSmNcM07hE7wUhOAuHSs+inKQorf5AMy6td2DAH0JzgLI+s1jn1GUppyCr
nRZdQtXXSPqXpu7rPVUot7CbqRPuh8y3qJwa3Axk1yxa8/JnYbUw/AVQifOmxHp+
KhYM37di3c7lKsbbqn414Qu09A/XKKIqmMmPuXT6DMaQPPMlHJBVOfe0a3zX3Tg2
aOjjty5gGbCwUjPg8BBzMkiTWUsEGVzwFKnoiEHgWCkkpm4IgrRbAXzmSVUPKovb
naHq19oFpzT3zNvn/E6dO2xRfEzzw1BURW6gscKgBXM32znFem3LJ+E2Z4WhWuay
Iu7G1GXG6brFj5w8Au9b3ucdLmuvSUbF9V/JggwC70qRGeBWqWShDZBQQNNSwaLv
6uDUqe3ODTzkMXu8JBWeb+bPqEBYNUYdmiH7ql1cIc90+OsmikRe6QTXCG3ZTOdr
4FUSRBGKIUJcm0tFwcPJlQGsObyJzw/qS0RjXy23kZFc0R1VqkowskjTs+0PVR7J
d7NUwOyD5p+VAngNUUyVh40F6VHf9p8nBCUEQ468Fj5sq0GiGYQRWsIzqLG2SdRp
rhYlUr0PhvL1nazRVRAIbi7T9flL0/rs5F1AC8evC4H0isSA+gqUowJrZETBvRsJ
O66aOIXf4hwZH/L7hBaHBZJl9bcU4YirQVCLn9f7J4hErpnzRPBiwtdl81ayYwGx
r0oWLI9o6gZYKJ1eLNuFhQ+Z9RDfzi5v84lXhRyXYj0X8wW0/KsBdvf+IAHsdaA2
3q4mDg80cL7PnM+0DBrx730+OvgcgBUreGspD4CaTVKXPTKzpxaHMjOVkdwoYGiN
Oa0G7y+B2Ork4ps9EdVeah0aewu310O3CBcM8csGgryG/Eb4JGJQA2DjIt/ZhNaM
G84hDLWlY84/hvpVz8Wjy6VAApgidqRG47tSDIJCDifFhlk50WakH1ooNz8XUvoh
CR6xP2bsAMomWeQ+ZW4asw1OD7UbJKyIuy4qtF9amay6NkKvxMC9Cbjf1E4RPWBI
jM9hjuC1w3os5sTzk1Sff+44rrKAGFDn+ayFOSQ2e3r0p2QQUgbfYydmBiq3GBxP
JUJ/hrU3TH4fDFSUpMlZeHz9dmlDGFG+Xnna4cg2xncixGQhbpazsvOdC9MN7Hmd
RFX+eW6HvqSAeOD/N7Yp95mKaA0ap/ucs7rNa+EJ5d6SU35ynjBwnZK7AQZSgJKP
fFwJofbQS82mczmfGUxd5WPPoZQnR2MYRMC9/Ir27OdFFtxX1AESCDNg5IOfUWwW
DwtacWch3dP7OIpgsOveEAuY4b+myBBdMNy3B4evN6ALOpaeV2leD9SaHGwoHDDZ
e3hOPX+ZoafvEzcS7ezAmfkxQ3f9XtLkh5UbzmpvFr23wAoL94lB/Pf0D1rglUX0
67Es7menphKoM+l0VfKhO6gacxVrJ8EAVOEeq+zFOwh44KIyyhs7c3jsrzJyzbdd
7aJK7ZavMSZfc4Kf1ic1D2Un90KtKXZXYlHRDMkdGp7qsvnS6hMw3L7dGKa+e7Xl
1nLVN5Tt+NwhnT3eu2LvIMyrgDikn4ChJJBjPE+9KaPlvu5KxFy5qWWaPEKyGTnC
Nb4pkldj7tv+C2rn+0n4/xJmUur/mJILF3ehy1H0mAWRw4FxNCyeSQvgjtgR9q/V
2IWgq3+VAtUql58KyrgV6pifEq6weFKgfa7Nh72V2UfRBQo9/DngJODrcljzX395
cXHKAk7kTSghTTXa8PesmF8pwbRFGxNqjcKDJpq5oJUZZFOtOBgztwEf7w6jKHU6
8mTQ+e4vTJC3NeyUGVA75TM5zbWP7byQD/eA57t3p3tPcrR+NGIFNeJ1/lcZ0P9b
f+te02IPDZfViED/x1lLUJDz7stahm6zrobCzjC64eB3PrgyeBmWKplH/9aElpxv
bbZFdFFWuU/w9lkEVplKehm5AX7cuTf2gzuYMNDwKOKrwN89orlstuLrvTKUlfe+
wvM4yFTAFOVWirR4BZBfxUhCGtEZxlsECRKMLFo+B67UTT2aq2dNXhdqQScyx7E/
uwHNVColy7hjxhaCsvk/1Pg5qOWZu/v87X3co9C/LRXCD1xPSZrp5OWTlQ8q2TOL
VHfz5dKLhHuYyKp9DRytoCBJ/u22BYUYxCerSHPRh+xxPntRqnGueADsgqPP+mFL
K/nn7aNQ0tCkD/lMf7Blik0j+jVpapneU7QTM8g+bAhZXTqoXUykYQMwDkJHMIdT
gFY9LwS+14fp5i3Li7+bpvckLqSVLYIgNrg3Rx0wRLwYBUbjNqPaaD0pEYkA1SYD
zLq+cy/xFW7+dt2v5Hwbfo1hork6VD8bPGR/uD7qi1MQH1RyvlR2cbnjjvctQwXT
NJA9v7L3ue/Q1SimNhNypaHHCI1PIPz7zJT9+mQNpfhDWPSmgkzPJUHdQkiaan7v
30TFHnQSTUC9ZvPQ7gctQaGSUWowdIj0TrLC4mX9rEVxk+hmL2VkAAKP2zSyEEAb
06w0Xcv+GNTFeh5XOtU4XuLAbaTJ1TSvpyLw1URmaZf0+1dY0p3ZCw4N5GkgByS3
H6a4Yf3w76cL5oTGQfEzSR/TURv2/pYBiPIt5+oEd7Q6t4GPgysSGXdCmT0iMNEH
lVERtBAS47UBwYIuyNmXGs96/+hIwt/oUPXUPvI52lShdz+LpmU36ZABCy+uO7eu
ZPJCczOF98KMmPo/rKlAaYBAAJktpixdWQlMdJ9eQqmzGV+8KYNQ30A8UBVWAv1f
rjkQRAcYxcLRH+OnlbAqFcvmSPSXKJMiiAa0/OiBgjoVL211i6Fytiz14Fmzer0F
NaCqcnG+biojXTO+5cxEe1Ygn1o9tHV0rRMG0wdrBbzhXPwwhUqrkPXFHghXlv1c
LlMMVn4YWBLwGvRgEkQJw2ARk5x7PCdAVmgaWB0ODAZ3Wobf1TyauOZ8PBCrm34J
y7yiM/TpkgLHvLA3Pd3H34orRr5jvCcwZyRyP/jOh5/uTrvtIFTo7wFVoLrGqH9L
cN4SyabDsf/m7KSO6MpLKqUMDHBclF7fCr4hAU13fBSbPcAAy5HAXk1YgGZn1Con
GLwO6xNanYLwd8SArPUgfAj2zSnub4bGsoNmyLMZumdhcsJqOW4YvPViggQghcRt
LLdWipPabrkewpTF8+B7iQ067SJBujbAx8akw5omdVfI6V00fM1pxC2TkXRDPfDe
9+0zyKidtm7nXcqQwMwM92mIKhq1fo5ZrGj8/7OlBmn7FkK1zbeAKTjQ2KS6q8vu
6Er7j0P3wWFUtvz0koqmJEqcSuTcU//8ORcPIf7ro3ekSAPWthh2GijBkeIUe8TG
WvJuEdnCeaXrhHZ4V46+ZZyP8+xZP2RioMz3dNpQ9cfO0CMQhkKwfUIQ9m1APN2G
sEzqKfuzHHF2gEfgGopkLrO+91VnY1LkthoM6mgL9xcc0mOhXLGxugDmzpwcribX
GHpXp7/zpH9WtFMhwtfdMBmlnqQ9KxXU1Kdwn1oIBG8P0oGJgozd7Cjw7Ma00a7y
/dOZTvO9u2kb2RFaKz4Lc3sUu1AL2Z9TgcqXnI9zG6IAi+tm9Y1ea969kde2Mxgg
lYX4LqgrboFlZ/fGpOZdJrf68Gr6tBO7L727+fd10tG+Sn1Qej1U1snaM7rXmsz/
rlxbLUHxMllFXqx9LJT8nazrdXdWhPgpO2QDq9/FwIWdjbz6aQxUqP31m3SuoxxM
+G+FsVaN90QcvL0PEstlAZ1Hb/5+tMI2YXPsvVgnghyJJH+2qzONE+ledLmkj7n3
v6BlGhxrmCf/1Z+L90Ul8ejW84lOkIugWe5vd3koahN8wUhlkQZ7OifKXf1UdKgq
mHitlQQoLrYpw4nL918e3w==
`protect END_PROTECTED
