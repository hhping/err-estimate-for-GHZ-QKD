`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jWBwunvzOsqGrwt/xaswGC6A+ldmZRcL2ArHj7G5z/RUQ7fDZQH0Csr/3SyB1XP
dWGqxCdvTotIQPrCbnwrxfJKX3iP2xK7vHeGZvWCHMjOpJbCYsXB1wgLsedYx2XI
GpntTYNlFUh/JaQWJ26j35cC7XJmsNzpT/Ep43SqVdJ+LFJnSdT9OU7yiv2BTITN
/GOrkLlbzQGlmh+ASGa8yhOEnnRw8EXZZCz/Thx35J9Xz/Ag+8e68zu67taMrX+k
cpNZv77cidUp4uyl6cMuHO3WGcA3Wym+k/vLV+T02qbliqACsXB155wEy18hYQ7F
IuUcIj2UAxX8xuD920hm4yoGEPN9hLkVCkHGq9L3QU+a/SmilRij3JwfgItX7Elx
KBeTCCnQGTypS3Dr8ekgHFUIoJI4JcQxRXsjNurEYJK19ubp5LMgCLsSItoASQ98
CM0+GnAOnZtw1jQBjzhX3r6W8ebn3pbZYIoCOQySxETNk2ADQGP4x/lrwideg1zC
bHXp3t89dki1HuG0yaPw2QYX/bw54osIUioT7TkmoX1dFJ5PG7N8PJPRqOvVikiI
HcJu62jroocjm3Ma0RYI9Wot6nHTRz5DMIJsBAZ4EC9w72wRg9ilk5WkvGRaJbVG
dHsLMPHYdIoIeollEGvrcIjSO1T/U/cwSs+pNBspNdplq4/1kOI3aXrEjyjiqkUJ
OpwM+YP3jKIAG8sfngY/4CFzbliOGapDKClmoTAqgKW/G8CqWlLuJIVCQE9zP77j
YmiElpx4bBtn3QGXU6qNIbBfkXOSaSGbVRodWF5uOO9eqo2VlRP7u/LC9WE5I57V
4pafxrYNDnPLFD4M+uFqq2SlibCMjzZw9aeKZGW2KjJPiXNhGcuAXc1klRNZy38D
nqQ1HLjQfVOsyOSV6roXw2t7a2oGCfkNHnnUT7IsoCc=
`protect END_PROTECTED
