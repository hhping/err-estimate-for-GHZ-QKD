`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tk8lqS0bfWgnGrCCVKbxgDoD60M4og6JvIX2QpGMi/AapMySRVbwi5RYqWNknLXU
8Eb5G9iIcgX63If5mUdCQG2LX3biCIWcH8Z6rFAsmElZL6D/8yXpwxJ1DuxIHpLR
uBrzAyA26Y8RqEUr1N1Yb/KkOQhWGR0iGwLgQZJWuUuJ6/+xn2X/Ui/uIxSMLb10
iqjmSqn643PScLgWnzAm7epkphqLGX2cH8ePsYmbUEO8e8wRBgtGjchWx6VGZhU3
AvC0Sh1s1flXupZybacWxdba0KF2iZJpmbee+3iKEEJM2uRaeJdLe13zsABvJyKH
CxHYVGRVH5cspsVTnWsxpHjxPEPR17gUjl4nfJhmR8Ge3f28jbRfX/T1nY8/pcOg
lwpBCpKLZJ6xgvbfBji3aVxiFm1RurlFxBggHPfA7T7sP68QZeVp37vDdHTayXBJ
u/ja3bHZd9lQQvoFxicQ/w==
`protect END_PROTECTED
