`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
liOmXg0SdL8cJHUvJ9+vPDk+GbNh2puj7mFgxbSPtXxV4tz4pdK+Lt9E7jGPGNzB
ZvBHBqmm1+yMKOAUiEDzQTXA27BY3Xwn689gYPtZQmnblMV0iOC70RqVvthwVlG0
JhS7JMHKGpXcL6MboMJGsIBgOpmmOONdbC3J1+fRO1bXd6uWR3WgkkyrqF5FXDWc
VvggpRjmUlpGZDgnDh3vsSslADiEWohDX+OUY0n/IQTYn1H+NRjH3+cHaFMLUCYj
NS+Yq0V3LDFdx2W7x7pVgfcxSCkW8v7HOjkoMQgsd+A6jtDkWKhursYeUKsEJTmZ
wzLRcgwXQttW83jOHh7ka8ZBYZ336nw2J9wzoRLDIIITiwgI8kA1jH3kY1eKhLUN
qltACxrkVD+ZDXdZOoLx5gRo5PIFA9f9sPUbI42vclWOFleV9Aq7uDa6jKZrh4C5
CJu8tLHw//xJWzSHF3WSsAvrolVJfsCiDn7GiyRaYpiISHwEGvCX3bvrokBa96Ke
h9yHJs70j5Kpjpy1S9U7+ALOM9Mf1C16cb7Jvj7+N4SZ9yn/2dMDIhYrI8vuM6HM
rvH5AfyCfGZm4cMETXk/5K8G+Wvli+h41daOG4vy1xpZG13fwP9L+o+z9TAKVNrm
AzAOc5gVyIyFnwZTTzdzzK1pEBOYcO8EnvdaOi8NTZxpvo4s9+AUM8ZrvdvRZGO5
2YfqreMbHpcJl3GcmEoVGeYB3P+gK+FyCqkv0qRxh+rDiI32PZuXyssljKK9Hhz5
eRjlzSsWeLsbiBFuQHHikXT3qvfKz1JYfyfxClRPj9NZa7/ity5Db2G1bFL1QspZ
Eh1kjOTXlvk1h/vVK7CtImUs4ZnGLdpZ3DCjBygLr5LJeG37eQ4GqxzbH3nzSiSX
FrRpzchGhO5YSScgLGZ62IAr8PKNzPQzus8NrjVmSPzXD5+KPEJx6EcFtZNKPcmN
WlsEDvEfUtap6k6GlzhMCCVLpBMVwLvvjhfuNoJXQCo+eSz6hiA92GEuiu1wLELc
quWmlgoHYTz3ruHUZ+EH63Ea642aV/7SIWahYkDyKY6+Ni6Sd7uQFbEnFejzyXZa
Vn8H1Q2/EnlLaq+nYTCZ3fo08oEj05JUw6XY9V+Ub07cYvs+sVK+wjU/ei+tWzOC
fND7BcVvGJvY+BB4R8PvThXOvEfMf4rmR63GTaSae5CX8IZ4IjKOK+6pksUFDLIB
MfVchvU0XvO3i8Jk+X9LNT7/+rXDInZOB8m7DsG+l/fmT915i3Yp3v8gOpCSVpH7
EUpqDYamUZzacKDXB4IgdJvf/aglQGfoCyfP1snvwJfRkzB4/yIRGg6WgU6OK7mU
tF1OGXZBgSM0aoQbBaDNpDD7viFzZxkR7Y287DHnwnmSHjMNUNk9dDwvwlDXHzOS
wdDVy70qBUIvqdyazSrxKqBWWMxnHr3G2RjfvyXWnWKAolCHlwwnLjnGCzVdTMdG
+p1Ce6tHUQkbZiR93HxvzN1kFOwKP/yX3InBR/YpUnWV6RoilNG19EeuMp6nr6J/
vgYFFPIe8oVIt0i0QTgu8fcDUhxwyhnS3cw08t2LlsK5vin1gPK3MnjzG0SQdQhO
ib5QCtHcm3130sYsHzOXIvH0Vq1YOkj10xIPfIgeY+453L1kwNfgf06z/wli3AwI
c7ZX6YiYt98cv1mnVut5RfHwTKD1UnvhDeuAEV7BUUXk3LYaZro3pH5p/1ZpYJEE
XrSBZ0WbDLl56saxAVevkZHi9V8Ckdzi5EWyQx8Rl89IaJNOyybVnPYY03nmRsF+
U8jcKFbG6HO9i6EphLTXi8pNSr5qzo822vydmjlwDhq5mgNToJ5rp8+coMwPrPCO
FZs8017frSlQL/DGDytQ6E6Qm4IQlTTcbAey5mSeXvZZlrCeUJzSNFwcMOdDoosD
EI4Zu2zd+7Ipx469tmSqhaSAxjI0mJxVQMkKuwYn84GfQL414uyZqrHJ5H9Rwboc
spg+WT9mRqVNhIf9xHHRUvDLy794I7WgBmFDfN32uTVo4bOLyjaENd+Awgx2hdtn
vNmOfVVpohkd0oj+81iHKzmLDSb4dd8gk0QvsTnngBezaLEqYfS3trpQugxcj9K8
a5lkyksLdvWTbZFRLky2bR9W0JBWwakJS5GYb2+UTnO7vJ8MnTIf62iPedxwK/G2
b3S4Cyb2nR+ZlnOKGuedAjUu08EctnOeg8o3RYsLxltC00OgV/SQy19AqwpR3hNO
7ce+UyWylSH4FYsWZQ0XVTavvFavntu3pvS8c8qBg+ymopFfaTWkXg/zVDtu+DT+
WzkHernAsdyG/SCNiHzPKbvwI9aKpK+Utabg2n5LP9+roYUazNQUqY16w/ZCtWj+
t606YAvIl3741AXoV+AnJR3zBsZVrg1qsmtnMceXf3bJ+oz3mfidvPUux6mF8nDY
ww6HRbAGcjC2QtR1PW74K0OuEqARVQsaqwGxVu3gLwghrIdxDcAYPpnS/fKFwKoq
X604nl2nOX/JlYjmy9SN+w==
`protect END_PROTECTED
