`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zh2uNFCg2EeOXtpI6H51GKZ4EaVxTDCSESvyOlrOzQ0NfrR2YrkyJo/e90WtK3km
Om2mbWydK76UsCjist5uPu3Kt9sY30o43Sttj3/7gjxKcZvxb6v8G3O3g/JrWAoi
r4D/SQXyI7wisFh5+GN/rGOteTbjA5GgBReGHhIjNfEp8UGZ+WUQeaJigxb8lmRy
4VMcfa++9Ppj0v6C+iJAjdinHsQboL37nOdsAc2Q3PLlcI1grqSf9KGtHzzUvK/u
OkVaStiee5vCeEgQSjw5dy23ZiQ7EEXnytF1rm0RStOieuyPgdra3msltIiqMQpa
RDzd87P5DvN9FgGHsegsBKYCxS2HrQxZCfROSXM2MjoBYcoQdVaBooGgzNOtbPKD
5mHz/F0rPZDq5wHYg6GTmoY8LP0+KmQY4J4t+gTtmYvfhIF73HQSHP58oeR8UAqu
1BJ6H4Qrc9rnnr2M6mFNLX2i4qEMQetYKLxWHlsfXBeNOxqj1U5adQ68Pk6KRiuL
UGQSIdnIHFaCculu3FX70tLILqyRtlhbRzof9xRpKhQgaqDmq9/FcLeYVszz7geL
BHdqH0PMNHZozGoLWwqaujGvSSAsMwKcS8fJZ/7GKvwM8F8742C0rgxbTRKLz4ZT
qGPSko+IwyRGwpaCIMeQJxFHDjcu3D+iaykGBptBsDJdvyKuUttxBCHdZ5CGDyry
676IERTe61GeqnO4jjwBaHjuCN9xLTekXQESFTtAAuH318tJW8VUbsmhqfrgjQ/z
7/MMfDU0ChVqoKJog6dSGe3KVulqz6vBZpalA1xOHNYTyV+ovK1B4ArKJ27s9Kzs
1S3fjRslns7MfbneTi+wIHDJEvhdDQwZ5fTSWMS7/ySyXJ57KylYm0KKwq3+WZIP
IO4WQDluA7UKgFZfE9I1B/Jcw32myKY4ipH2YBLI2pr8x1zNvuIllkR6XVFWqf84
FyKD2LQx4xFY6jqDRL8yF0Uo+8AkoKvPRT+6MXw7lLc8mooIBk9lK2DLUKi3XIxi
FATW+cRiP74arGal1RyTxtGAh0Pds0h9GxqSvSyNVb5p44Jj6mO0UVPcK3VBxPes
7cEQWOoB4yDDWwg6TTHd6zT2E2Gtr+lrNEf4fz1XL6sUuFXqA98uEesU0Ke9FIOG
`protect END_PROTECTED
