`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jdYvVAKlIVPQXQkwCv89MChQIymF6ELbsawOge6AUOts298FUvBBUaBr79jhCBgT
4uPtn4LwMfcO4wv1+1LfukDAJqCZn84s4hvps54tyUIwUX2arTENz9skGpFJCL13
3G/0wlPEmTLoCUID1t3I9Voshx/d1frbrZMK/GEBP4BZmAm731IL4UTzhzw/Za3f
qny1uGOsF1Y+j4HM1tLGNRxJvM3xG2i7qEB+Z2rsWr5MgxnJGRiRpTStZANwcz5s
8fpIL3uKZWi5iqdsnXYexQY/N2fH0vLLgJb9EcEu6sOD0xAw8rUldSPlbkrzlDSI
3Mgtsjz0GUxLqaPwzO/VIzms6cF3dHyTT/BYs0mOcODzF4eKQwQh9uvcCVisZdRo
kq7vhv6gEXxpYbhTauvdiMo9x7kUVt27dyRDE4bTT/eed7g6bKB14IGPeThpD+eH
`protect END_PROTECTED
