`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z27akRZl2yp89V7IFSsUQFZWWlnvY+kjiXy1lf4n1MrwteJnNxi+jcoTUifHJW/r
3UV/TB8WJis03fbqbU/nK3UGVv5g5Th3u43NXQ0q5w4X9Jtim4GGINhhpHTXADco
pjrQTUNxPP9iQMseLjoR2QRz9R4ukEVTkfUHlPoMWhKZKyg5+QK24U82DecdLp/9
3uSwFVPJ2QjPLmlfOJqZ5dHgcj645OhPoTLLQ8PLq98+VPC4yFM99lJrZGOwRAqk
jxmh6+Zwxthcahrx2uu/rduTQEV3cL7B1i8A+zKMSZRIu1xdHSItDnx1kjGuG6BM
bmNAK/qZjTmXJV3igaI3vpBl4KfMjD+OpbK93ds0z9sHGWu6lEo3Ch5d0PSRcuOr
LWKFry267GUwIiGMc5MohcHeYeE0oUzWrGQEvEbleM8nbWA9yvTUR4eaUX9/B1gt
6x9ht9BtKwQdsw81fuqbyQafXCmhXWVYKn+WNoRLVXP5BHSfv/s+wg3p+TO8ZmGw
J9KsYXv4MzQ2U24xTw/rk4VuikksVwJy92PHzdZqimyAT1f1Qtrd8w6LaxjrypyB
WkeFD5WoKqVKBMKGb9gNdtfSo3FVOQkhbdI981RuJ3Pp4ulnkSKUCI/Wc+CvEXKz
/frsHi/GyLIMqa5fXTzTnKu6QuwK2rKo+7xTqF8LSSlqYCDkBMokVhVjeMwOfrqb
YN8nwFXqgwLWf7KSOAEdtLgEx26zaq1vxxZfUpeG5ywzbeTBUvUIsK4iiuVj0cod
oCVDxzckkwmHjc3PpojNvLgSZXvYTj33qcOXtIlTrUnJxkJW6oWP51ldcfZRZE39
rDMZpOGh0a9QBhPhZWH1uTwycSscIKwmLD6Xd/z+FWV0RkPl3S2yGM7bPKdAblnV
QbnzxBwTIFIcxHomnQDUXxZb5s+O2R2iyPQKJERAbi+6UEs2bvQuDsdp7Ju+drpf
gJW+3meGNCKs7W5TM6EkRMfojKoikJMIeTsaApp3ip5PhdFxRVOmHxClaXjpDooZ
mlBbmuKA3VRzsZFO61yIQzsU2sWWUs64djPa3+PG6ORrOc88skvt5JwbSRiEZeLo
2Idexwyhqhd3xA4fWVw6jR2L7WcvhPj3b4ZEQJJKuo1eijUHBpXaIEY0c67OtoNT
ly0QYcGIzWckKnHrIU+Rx3nmHJh21O50EGeGBACF6k3/uVE4/JGozD3DxOMpJ6aR
J6RTGc3IYqfbA2+OYBk+v1NR9yy9ghEgYeM6qAWLWDqWftQtiLnmagOj/VVD3gRZ
CFUs3oInI3O04+ctISMUv1vQNCF0ay10lFsrnVgH34WxWpebkdL452W5HrnyuKiR
QTr7e4rncEanSrjInL4Y5SvS1TkWzxcx+A92U5Iuczb3FkRjHmG6NHr/CwOKNqlN
q5tDTHWZPguQnDOMq5vmYGMkbvrfNvjwZNTaCkLGL++iZ4WqUcVqqEKIaS6eN8JZ
yX6MqtRBtz12ki3KY420nENgI+g0dJEis6+LH7FF2jmoV+jk2IdH2OQO2AV1gAyH
JUbQHTAgIOb+3caEllYOCSWOIjt6RxbDebtsv8qCTU2ekLZ3uNrj2XxVo690MMtw
+9NylG+B2lpz4ToKHVNyFjJ+lKeMxRPcd4XBLfiRCqWmKtVVjuKQpde5AwdUFUNs
Ht+y8c3LIJ05yUBxKG56eKlgx1RMz/I7oqSDyw4OmI0QvHl8ty3Sl0qAUyyLPuY3
ixzseIFqWFjFF+vGKVmMChR1UxFOxCBbqBIWb9F2BB87AARFwdUncttFRUNB7SxL
/IP21ahtvdEF3GCNqR7ee3VM3LFopOeotEYEJEXURcg24Z6hTf1/bWNbni4XYtnz
op3OhCYEvtEuzEmcXlSMtatjj0PxgW6kCNmD15bk6tJtECAElRNIrTTt0+QAuJg1
K+AzcR4Vpqcc/fQIZHcg5JAQAZlU2bo56FubU6g4jyQHXSuhdvvXLqi5iHhN9y7H
CwAsGQmorSUlbm8nqXA0Yi3n//cknTElIlZC+EIV6ftBcUpFyL6bEu3pERBEhzN7
47BOK5cTygruTwsYoN9nSJ8HHGR76CYSUxvQRTReTHyUA0dntoK4rCvg/i8iMVGo
lE5TLx4ZYJX/PSeCL9+fuPhYzlY7il1qMND6e4cPiQhE8bsdrucdz3UZopUew4bX
4qSmwN4oECVOFgH9NnpyG+bl3b8Yf3yd6f0QJ5gYQOkq34v6qczRVYzkRVHxQYya
W/RN58vKKsDGQiE+AUh7ELcUNiAwS43ojujk6+ML2/znftiXyoUYDtUrdc1/zooD
GccnM8Wqm/y56akFGBjG7P8A8SiFYwxgcf2tfz7HJBC7RX6MKNLMLgDC0IXGm4jf
4gyZ2FLjhpviQFSrJ1I8ivwIfCZMzy2rMnA008OrDYXINty1wGC6KKk6pHSRfdwb
mGzDWS4WLLBmJuSGaOdCnkLnAspbawFByYq2pLszjEFU20lZimJ0U+NTQ6+2QEGE
MTBV82NHmiU5lLP7N+zII95y6i8MCkS77nsDpTYtqE0BcU6Rg7ETQQ1e/Mk5qHZ9
SowriKwqK0zyvZ0hs0qZ9jmMfVBsTiwCsPrEypfmZAsKUYQ3WqWHcgwne3hm/sBt
XdYq3IX9oKhXz9HnuhQQmFyrcmOGgcEKFHcRK1Xecm1AuGl7QGW94vTi0jKtTs4n
j9SwxRfZuNCfBlMosCqz/69rx3v+2zJM+vfs0B7NX3KdtSsmYFdju4yp7gt8YsZK
P/6IuTkSxoViFtEK52Fp0SPhuxzljCNxZhK7iDP9oZ+He2nLiJjcb1EVW2QwsKfx
Inu7jXKt/rUgo+HKGkIb0zN0mK3QPbwZxBF8wff0xYlYaoHdochJNbQRDNBgwkVh
NN/OxSp2TNdCnIyTuqj8NJElautKkvNRTOBgIM17r+DOrREf6rP0OqVs2VIYIrwS
oBCjJnMa5vrTyxu1WpNiP/bk5KufifLiUIgyxMBWsWPJFl4ZtaYfVHpLK9JB1gjM
DBRsxYVykFq36yA+8TdGCLL7TryKW9BKeKgWKmFzKMcdfERrsC+o6QyPr4NJnwuN
euPHyxgZIi3cQuxg7nvaIx1pu1zRIylqsJv4Mn6V9qF3GIlWXvH0Kn2PjuQTre18
MTdj+mCSp2/S+BZrI0vgCJTvlBMz/wHYmjl53m4Vx+VucerZ/Qe2VqEiuhSaQFaF
MVHwQlNmp/XWSjJIN4mogcpWuUlIyIP2b8Y+1kXi/EtYHLPZILt5H6eWaCbD7iOg
caMSQUDYWRzzkq2/7Akj+w0fRTHQ4IoDzGM9eECoxAAtSZTSnnezGTqeYlzSo18Q
KgX4DR53rAKJqFs/0IQKkG4akCgcofmvujTs8MnKyby0rzl+NdmbF9UCdXz+WXhY
+k9PWqv2Acl5jJBkOgFSscg0qSoPbXCbHZ7zIWupypTjBJ5tS5l5pbm3JYlNk91Z
NcyWwVaN3hXZSihNjdsLW2yGLcUbU9vyN0JsFOzZF7dJDvB7UGUQF42OJfvYjNal
4PqO0cwXxKaVNfYUfWt9qmStSm7423HnoThUYehMGamHDnKMWuhmxfJ8hhVYBl2P
1OEwBXLunSaoM1s8SXtj3n1v9TG0gVVuBoKoJXlrFD6/acyLfZjv/SPoMfejEPTY
G2ty/JXEaZx29+e16kbZ01T9eCTU+xHxM2dcEd0+YzeOOXhQ6HfrzVtJtb9Y3C8P
rohTthuobrfFZpeX/YlMhiSmSYuEfuLkrX4jwv0XSC1gLuD2gXFEOpBQ2tbSfGad
Poh9qcoEZyDp5ljd7JGwEW15w1rfZPVBl1a8YTyd4DeqUXl+/5NDbkDHUeKKhOOd
mQVfUMo4t5Bbe+sEzXFlbyZNtLyEW1jMd6VFQo2vvQzlXrhKrUw1+ruXudJI9IPs
vpHm1PTKmfr9z5UGfs25hY+xUjS76LoG8OzBaQSQQ5bAmEZ/cL7YM0zzoDf4HAVM
CorORFhvVUufqG7VXcQRSHgUvnk9jv33vsXExqyAG/GM53/Gmnkn5okvckL26lCj
CHCxEOoXf3g9a6s7j+YNeTzHNaxgFS4aMqmZ4oib80i46NuF44D92j3LW0nK/xzP
O1G6rtE3nvcDUwA0s93/S+wi7iNQ1V5wxCJZIkK7zX7xDgXYA+1qUNbXLGkvDF8p
G6Z2rK68TeFLTcEURYogndrz4YgCxJVSeP0USkSYxI7dD47Qw977/Yss3CrA6r+q
hVo4pYLyEQheHawwq8SufhNFtiUKW6yYp/LhMgrF8zYISo16qPpahdBqviVQ9KPf
kKLLXfX4/evTCaLsHhKQjJo5656TRpTb/iy96rwgVz2pLwq1yKQCChihaCbMLKdv
nZkAoYAOjrvAS9zQAV2mt2Qc+5au9A8c9IhIutQEAVFV5+HEFtG93lkRFeVzm9ZU
DDcht52ePxHReWoFJES9/mLBAyYInURReD7WlIE9te2OzdfWKhItvGyDK+/sNbSY
HnaH3jnzj7nIKNByhpiyShsC/rHFRgDCEzmEbfkxSi+UxT9LPLOsfAGQ6wOOd8nZ
aHOkZvJ8Tvc2oa69QY31dQDkdNV6PpyGrulPsHDZzIxMzCv0x/DXr3mzMjSP8nSo
S4WUa+h3fB+SbxnLzpS0kIg7Lfa6v0n8iFfIG9tdY/zowzWRJq9y6hdutjuh3anp
nVnRWlBcsY2EuRyfNhZmGaiCuicVmdWs3766WOETjk41jnRR6oq2PuDaun/bhM3K
g3qwHS7COUyOn7N40CF/XuUakLVBXGjVno4oQzcYIaT4Qp/7oZTUzlor1QV2/R8P
ICfj8mBqM6N/uqNXHapiO3fSYTWF8JJvPjrw+uPrKkOXB6MDyuwmbP60lnXzh66W
LqtaHbXccqgDSldFx51/bDqqOcSX+GLaHyQitQy+ZRm8gA6Ak5MvI/fSZt4pwVRp
0YkJlR59K6eKCC7mukKiFMuATpB4t/7uJwf7IWLWVwuuaqFERKkLqBMcRDge2q4+
AebzmHeSmWvPy2blV1iL7Ns0Sbp8Hv2ok7GQ93gb+yuyGZGAveKQ6sU1+gj7LTnq
rLBgVPCl8/tfySiLVca3hesCuO8tD+BKXOafFuTk3WgpwOS3nP4TYGpLfqUUtFLG
jSt0Fg8zRSyJ9qXvhgsmsUPumGCi0hhUyNP8+rE3fvoDpMAd4G2qvVUbR+H7RN7y
INIeSpHBibJh+RfELcyLvaT8Z+gRyq510dd0JmK9kIbpPvulFaNyiVtzct16yDNn
zWn0aXE6sl5+xvbrbib3V0DUZCur9kpJbbTJaSXGZ24dEB37ol/Xmy2a0CZAP4sx
hZH8uV2HyJF+Yq3cviZVTEMtNToVCsbJNHyx/Rx9hLryH+x7Krqhgr2i1fBE0UCG
w/ur+j81UqcYSIlLebFfziP2sQqNA8NE+9nfFTGEXUZNPE8kLF1Z/LKjRDUl25nZ
/GCCHHwyrxFqRvPy40UvgE0TrH+epXk3MSEZB97buzBiTVicp20Cp+omJTGNA3au
AlFuJRF+QxGmPjYS8LqmMmHytVtEGv5quhlrL5l0+fHAuIYkxnBQsTkliKd6vAUF
sjyHKfWY3ypVETHDgabI8KCg1eG1Bvr+48PpXy658IbqDT3vUKNLOqJ+9m/o2y8b
+DoEu9gnOIcSmxW/DlujJ/vVGLpCcTPUoTh7RvrG+kY0VE+oVVVmf5Oqn6u29Anp
ljpwuaepz0wzwQDYfiu0wG9DSldLQ7YpG5tOBresJkEKs24JELxldzHZDAY/J7TI
sG/dkKfepxZjyQX2gBOTVW8qtViIQtqoC0x8Y4/bX62qnXtVcfjrunU5aC3Q/NTF
1FMZXUgkFujOL7loz27XxUiUc/4YzICzsHb7zqkk9p6NTv5IxZ648nU/pLhryEwV
aDAq6XbMIFHKah3NUxvOVuUDRCKKbhwBEYoC1gOeSedloxrR7pQi3YeTEJ8xbaDh
IAkRLN1Mdr6isOI5a5pLCNTRxe4OzaF3+nO+i3rzkiJdQJqoJ1+4E7twXiAowkZL
Ta+6grYJvNpQFlNe7rJJGauejytv4UYrknAqq3kZAhiQKL8VGHMujSH7OIVX92PM
6lBAYOSGiicXzAeNSZauUuYfYHKRL07a/4THzqCXjRNVRPyOFiOHbyelujUWbr25
Yv5Amq/gP1BjMs5DMTxyVzCzQVg9pZ22a67FgK6mW0+Bl0/n+1JCtT0/haCBRxR/
OsPlxtPgKo0ft1TwSZWLFiDIzTZ9v/mT2EZLektHeDFbEze9P8kSTweEcyikIYS3
faVK/M+678scWskxm5rq62AtYjSv8bTJw+J+G9N2u+UtDpxZFKmdaTFnZLiKEcWS
jftK3QkZ1cDUnqUZNB2cqfVxlqBvI3Fqbvv5ikmyZ1r5B+8LUpDgPCPk5L4uH/sa
lB8mFITWhrG7ek30xkGn9ODwya6coYFKVhYmCb0RS+Mh6h2DoSbhMfJbK5dM1oBL
lAax1TMblmQmCRtF4jYBbLNLA7SKr4ZBROo+LHDggxX2TbAmYT8NmFw1fUl54E9y
ZuUYlv/YL4+DbBmi5w5fWLJ5qILzf5qcMbKQitruS9vBDv7RzmsXXl/lIEPJ/wwW
Mj+VA9piZ8EgpdzhysIDkNT0vmob3VUFPQlB3TSXgw0yPtvT0K4rBjRKk/h18b5Q
CUB6SQZBHrlvaeP1NjQVegldjkOCAjbyzJrXfvKKc+oq4wvmwGSOxkHmO7Gy2yoZ
K9/RX57T7eLCXH9IZCDm1SzgjMVWYV6Nb7EPg1ix7lBkpVCaJ7XMYUrnMb0dcqS/
d7f8y2h4MeVRircvO0b7oqL0g8Qd7s4WbKfuot4CI9q5RllvV21N+Oqvwpm4kV50
EZkSUu6nlAgbLaV7c+7YtaO7ZNwIbL7D72fHVeiaOijNSRHiSzb6x6jV7PjWkcF2
c/wSz5zubvmjDUCjsyyYO0ADGMezIGQCnVhyXVSCx7O4fyiQdkMufCJ2YyIKVwdj
BDy28aManQHWdld90Z10dZw+T7E6cTx82HfcO2+EJ9qR5d6m1hDIF5ieYv+gxd0y
fh4oH2IAywaD7nrW05LOrgg+YA3JDQDCJQ7XWUrLOqdpLk87swh9N6sb13uX7qX+
TkKB1zxRvJZtBthOTQOjDSWUtXgM/GoJJD9aa32FUNgGeI65iRIpi9TOCGxQ9i2G
7MB9R6ChdblV+tGOCcEjg8WEskHrvNv8i0hjpRZFDQCAX9dBZLr9QplzQ0RPaL6f
CjyHjHMiYJAgj9Ad0AaiQs5zfhIzEX8U6a1yC1wQcPB8TrzInCGNUwkhkE8rIFSK
0iluDctnX9lGX5io37/XQPR89LqASIXfHNpmtcnLktPjx4wkarK7nkQ3n6qwz5Jp
lXSLOScw2QJMnGYJHE0JLOqrj3JzyzCy/Jn668aHvYdN9rzwFCUeZHOMg3KC10Ii
xL1txBZlgRtHdZxSzp7Q4oyN3x469gaCkApQQ789rs7+rppiSEggcmcVnpfROF2+
6MxgPxOhENvIhdHLlyiZWmQNZHylxzKjAIDP2UJEfTn7gHmTL4aXbCFQowhMfLcA
Xratki4xcs7ejXFY0lnp9hpyiF8jRDY5vwv/7R3hwchylD5ooRHtuUTokpY7XbV9
Luh0s0tmwORPsTYO22tO9sBnkSbdmFBNH3qVFdsCZy2SI2mi2JnJo8a81nAJ/yDN
bLVB8TtM4qYaKNU/j3cs1+01J4h0KSDNdUDAub+lNQZjMyBbSOvQZiPNKt8rQmh1
dArMjsi02kOPV1EvLhbk1bKrnVjCKhefK8V9eHlDEpy41yAcCDe6gLDE7DqclDgg
Ojdr4vDXwd08HKlxMSH2cFa6Oay7h0OajgqQR0pq+1KLnDbl9DUTZXu9viK8jBsm
nK9Ps+nUHPxuso5ms1jVxzHk3wovhy01ZHAZIOywyc57JOjttjRALyOLekEPATCJ
5CWo+NHwauIE9lUEA5udvg/hsAw0W7H45jUCRf8N+Wu4vpkxbnUClpG6Jrf5pNoW
5EYsPlFBzR84nwIpjPMiP4owWExlQQfdaTmvtexJzWZqwHlU7kDvk1u68waXCJNC
lEo0lM1RWplZGa0d/cxUr234DfCxSivbhfkDbzI/KJItqL5XK/ezL8dah+ATtDVc
Yd2o64QMgMDqWX8aRtQyxS0VpcLD88rDAcJbb/jW7zpptzZBYaruKV6JxT1iKC7Q
HqLPWVfMoPFKGkPg8zeLfGjI+PVZGvf0/DOM4pVeAPAGl+U4MoVRmrIgFcDUDon8
LTybyZSeY7DproTYZOY6F9VM9drIxqnRLcGgjMSj2ANmaI5RF7FW1QEPBf9liuZ2
YgR6EXjEVcMF5nWAJX0A7JFmmY9tm/htr8vslJfaXSA5qk7W/lI8DyDhlLYq0j/2
WhG1hMjkeYPvPn7KYXelnG7cmo7GH1ZQnuANWUY/MLre9FdViCrt+8GWS0HcLnZk
WHB6i3rpHMlkprP+ft/ZfdghvKufgWnGGgUk93NhYNgW8LQApmXsAp68JP8xB7W7
a27FwL0zarinbRuELtuatUDEaIfcrT2eINU6MyAPdBWKJtxFjNX9v6vKxUVDa5rL
WHh5zDQ2gufugfSg+CQu3inRFrdHtHrTkw53qjtnpx3QdYmhGuhJLTeS5GxpJvBs
xwRYhEzOvsBZwZ/oVIO7Um6QdzOyAzON3srP0FZKqtQurtuDv5EP7Lf7BIHcQxe1
Uj+X3tMxJaHJkR3Ilweh5aHqHv13r3qmN9N2mel6ggcfmzdE5J7o+EXBFNdZXIS7
2a1Yoa6Rl1MLM4R4a+FlYpqmVvSn5/NdqoxImsgrT8KeuoCQBJvrjiC5JS34wLE8
+7jYEE2Vr07BEHmhDeJZdC7pKxB3X/CH0uwxp0BfJmfgIZ7OznV2Lh2a4fqK9VKZ
UV2aylafvHOHK4A0AP55z9FTDVMftT+QDtbWDgeQdo/ih9y6EUDfGUz9YVY0rAcv
yHlOOULrV2dRXSwP18/FD6MuIKgq7ytS9HAWllS8C/oYEzg9dGUXg6RnWnSaT8cQ
pQ6qAmKfAhK5JjxcisKzBBFunSQAyML1y4nFNAFaMAbNUjdCVJd6y/KZkkqZuR8N
QhEgTyslV4li1QVaEOwoiW3nuiueedxNuX6t7hinMcoAAmCgDYKwlkljKh0btsIk
QrDIM76Ae0HHHbDxk2Lgd4xcgxjtsKxhqZUH5ksJbeL2OhEmKN62bCgVA9dR9ocF
vW+lKVX1UxghWNyj/NXfOsTLjIoyrtF3NAxFvrPwqgLsfsIn+n7NeAcbxr6eEnRf
9yyjyGeofuFhmoteEbZi7bxFECYywcgt+wm4F4yYW4PvxjAGUSP7aeizvOZTc2nt
lTniar501tjoxrdk9/R0Vgib9D7KVDmyQ6YsYkBD8sbCPQ/+WXC/TrzLQBxSjkba
vKVyohZqo6yMvdElr+S/Y/usRfA2jhbBWZwzDft326GP09lCxigtpFmiCn/jdAos
ZUS6qZoH2jt9n3EgPcc/jWIR1mYL47jb39m9f54QDe7MY/2sH1l8M17CL8yiqqmU
O+gaIZvDvgyuBDwdiJCc885lpoWlZTTNzd0WmO+sYJ7QNMZZi6Dmm0ySAg9ER9tp
5Albg8V10q5PE5XfOJFWWQIrDLRibVVfyVgPkhdZiX9wYI8CW1u370aMAzLH6MVT
uMuTqFHvcYTQjWceICNkudJgdizIcg+JPxtVcGEs3uzjRDz/xdb1m4Y8g0Oc9Qh2
TKmx9kcC/S1AS9mHw70ibq3Bro6tWJ3RdVG5IMP0pqpkDCDeAjyKi3hNhULMUAnG
uEMdS2WbIefwx2+Ynm4XvnER/unOvF76drYsTBTNzT4QufWxfUwI6FCRJW+KtTNv
BQ1KGHWtgaS/ULVwgo+zOtDM3IjwKg2R1SxDA+hHxSNlFIKfVkoEBqu0Vja6RWdt
/5d/qwBrU3ggEvs/PGEgH0eksktaB+Hpb585TabI1qLY+m4TDw4UMoB7nsHK8SZv
BgFnj3lsD/uOLSi9kcbnHIUGrsLG7yb9P84B5FqhD/tNfX6aTgrjvn0eMvyoU6rc
cKb9u/+574Bt7T2dej38EzwB74M7yxb+nYOh1C0f2j/9rTO8hXG4YwQaCkwMKvK3
wEnjxH2Qo0bBfoOLZcKK47allviJmgKhDzCXFXfBDYC6ZfzYFPiT1yJZlUEsO8Aq
n+qCAyEcOPJkinPRWhXrVKyCnULXP+Sz8R0HDJBkVFgNsl4TlVZ/tZepGtnKR3zA
HVsIm8SnILN4FN2ibhWw5iGGjUgJ8q/+EYXLcajgiORSo42b0fUioSJC5vKfo9JM
s1ctZxRCbCT0StLqk1xnthErpFDA1XwDHNF6Fzltw8/AigGbogNdVlbdXSfsuIki
EW8tGg9mNMw5pk+tIE49She2WDYp9QhmbveJNjRQLRNeuGhy8ocInQao22Gf/s+Q
CuxBavl6kmDWd9hp6GTCF2yW0uCS9U5k1HNN/NI1d89Sxah4sCeod8Ig/Fs5SdPN
6bsu2wwYT/pkP+H7RmMf6rUdu998UiQXd/NwaAjgjpKEKddSEi9Wl+aALdKwWlii
wId/ueNQfYHrlO5GJqPST9wf3UIaL0D6eKTPbjvzNAoDb2fwXz412nrCIsKpyR93
I/mnPNN2atz3IW+qAuxqVPpr4vaOpK6re/vK+p5Hwtr89WReoB5i7kPnzNI/tNOj
ffPjGwAptE0mmI7aZ4lmqopwa0BBlAVZWCDsv9duXj2GD5b1bl5jhEZeB4AUzm/y
gvoGSBwnzrG7CyS9t0D6U/4J+SkjdVFWln/+V1F6VfCdu+YV424oMZG+pxbNvJmd
aRaOcbMhU8pzOIwEobm3X7PvLUwpeM8SbltA5hfgmcQBs34yqFxdrBXAafX95EQb
TUGW6njsUypvqEcuLEmV/UxdeeoFYm33PBZWlcv7HBHoK/Wvgn1S1j2eI4mTvr5a
hIu1HskVkDwbOcAdTJn3Kk6sxSdta0R7gmS+1Bu1HxLMiFX+5tqiTRHCMhbTFFC5
InRaY2ICAd+fVYAX44j27Nz2cDOvqMezdv6mqf8LD7zhuDoTqeMFT90N8oct8s+j
wnCesaBDJgDrEkXkLR1L9TdMrAJd1FCIVenB1Uw33i4f63ZgV7eu+MJz0cA1Wrlq
Dl6G/4eTLudj4KQ7M2iOYSEIUgcApbpZsP4q13CjmOVZTuwIsF4xNAM31g1UvYhq
Z6Jo5Fi1IdR0sB1Ji7s+g6mwzAb1yqf76hplkCRVHpVQuWhlriN0DPD3x5MJsuLX
wM+jGRbAweM6nNjCFdf9obSGD3ikZErrBckaN0rQhxT9jjo9+Kb488ZfsHxg3RAi
fTgxMlxh6Bn4ZjcY+lmqkmXzK/+x2tfom2DPjTVSRUfr0UbdK7jEPQdMfnHjywLI
rp9KEfYihF6EiQ1cfkNAxmyQBrDayoEANB/gSF0YREHQR1dhkXzfKR09045F7Gx4
1EQpo5NsOZ9XQLEQXp5pEOOAH81tIiZuaDTzvIl0ET5VR84MpeVk7M/G5QoKH+Du
A6UqRWz99RoAaixb4/5PxQypoie8kgeNUbw/CfqF+UQ6dHQyGISLwqiVTF18tft4
NBcTjisvwhz8xjDMFExzA0cWO+36w0UCda6ZTpv1TGBvt8eicC67Ha5tvu9JFMeQ
RHO+jbnEaFSEauvEJpmZjDNmNclI/ifO4WYrhK88AUxzGawkxkLNgf44YzBkIbU/
ZMR2RnjN3whO4hCIhCmGUAtGbn3UExZZiMQ43GZjV7fXEfprqVHlg9EZhqwIs2MP
S4DBZIiWsVtR6YDx85e2KM9Rc1jkvCDcJPdx4GabPph9FrDV51Olgc2rKuWF6frN
4oaMERHdONtqdvYqjNYI8BFbG4Q7bbCyHKv6ZTKlAYJSJZAjArThC2TUCSpJl/ac
fhydRxv9QEVA5EmMopm++So8NHjaDOVXf+na3RRHidSFsdHJT5gS9JG7zdXdRzFC
/Bvuch9rEA83Yn9I+E0f8vz1C44DRjuJpf1fDfgDt8Hvv5FZLI7DVswZewzS5y5Y
WPE/Q+gqyWIcMbPwOF10gOIyeszYcc/iTc1cdYG8g8YyqwDzxPFii3cyuVafJ2eF
2HQ72rC02YNGVlQHjzOusV7KppNGgbUBfDbCWA6ZOX2RRJK2Ve2KUM3fL8J9+aQx
eT9i8FQCpqS102ylcz62E0JF6RkuaoduN6i5FuG1Xx1+AwvMIh986eR/n24DbPGX
54NvYiKlCGrfUfFQ5PhnQuq6zkkupAwRxPBg3XOpVfEXdXcOuMfwgzNB4XBWulU9
S/m6hgeB3HvfjGw33PiFpYDaNfWp43IgR+M1Dty9DYlzVHSMc/5TKPDCe0EsPFHL
hbYpzH55b0D7Si9yTbp3djEOk5wktJxIcncSgbN0x6dhct0vz7YGR6vB1NUMyR2J
PVzjXDnSPDSelBXAP8OqrRDu0p90NASVAcc7QTWks6b7QmE/LM+LVQCOvV+Y8Sv2
3nUF5BoRvLOOmxta9NHsFK2l8aJm4zDpkY5dOI3MYcHsEkskpVdv7cQwp4NgH0o3
SiBA9/vfA+oXhUJtQLey5ElZoSJ4TOKMyYoVSJZEzK2tNFSQd8aXRA2jKyskHPFt
aRldKDGSv7QgQusRY1mT3KxpU+bCk4/QeSNXrP3XIHnxMfaGl/DPi5kGHl1Tveud
GI5t7Lj65EKucB3/0pmPSwsfLWqfVPSP8ptpY/9j+bfER2ekQfNSBqgMta8Lh0uv
bzEMjm1RcXV0S5z9xIhLJpT0+eDIhIM5KCjkrET+Q3U88vZr/0eFKDa10WbXK2qa
q+adnUAi+c5BfuCa1P9DJPnL7tRglA4OAILCfPaYL5g0Jb+DMpbzJlQPvPxl5LOy
HGIQHzxyMdjhs41QZ9AEUisbHph5tibUC2KgLPeA6bIBNcCPV7QoVhE8QLdCw1bY
9M2G/70h6fdBvz1seceePY7VixVbtd93Yu+r9tXJjq7cI1ZmubSK/0hRE2j8m9VX
DsoiGfE13PLheq0XNnqsWEEYVB68F9L11ErG32pw9bW7ikvd8PN7NF8DVGlrIEU+
g+7tzr97Lx1uu4QQaLRYieU1FXgcpDKxKkm5ya6kBuHfQJMKzLeX5h2k1b5g/KX1
ZXfwo24sJxA4N0u18OkK4nUkWGHFrksF8Mq8G5B+3Dx0f1aTbe7U8J0e0kX6X2Oy
PX167XH6ezov2FhH+fPPBBxclgKZXFXftfZs5u+obkxO9yBP9wwDD/o3q+Nkvnv+
sb/hz2UqRvVuCG4a4wxQdw2FRYnquWrbW71HOnjJKtUID3JYpdCLgvJOyj2Kaevj
VL+V9ataERTH1YXUaRBuOmsZb+JdWNXj6ZlyLXLsgKk65dPBcEyOXQQtHg4kBkYq
nrxz+0N37ozT+9rDgQ7u9my551xbVp5LYVS4bFnYvvmdIgQmld2ClSAdY1e5+2ra
l2dx2EZjHO990BbI9CGpBEm0u2YHmGC6IXsbZ+EqWKPETCGjEHCTyMGPdkdnnUau
rJ5o07XD8fGmScwN2JUIYzdKjHp9Sl1MErm81Sxs7dfb1uXJbNRVKAIkg3VIa+Vp
YrIsX+RNT6XixUQz9bGS8zqv5bex3ArRzk1fYzeiA0uAUpQy1SDs/Bu6CVl7P96P
r4fn3HOL4fl9LhihdMZvm8677Jf37g5PR6S/WL48cWZWaoZc+FGYLmR0+CWNpcEA
XBwd8ygQTUlExUrTo75n5HJwMJtTdlJBBcpnBd8IVlCvbrUFUG5Kw5KNAqrQaHv+
YmTaN8jcMDIrRhg9oi9JAl8shm1pElBuidTc7p8YpCBI3IBfF5uxUiXpsQtLc6Op
LQ2mEQ62bggTaFhcxXCNntRMH2bB+8GZ9LUMZmkVrZn249QycakBxih19KTyiP+f
JukdH2VHiFAckD1vLUW67sdzUrYqmg6Bx2vFLHu7CQbrLMcGOIrqb+jQlpDqRABX
aQHj9xddIORpA992OdkNqBegSvZ0o8SiMQYT9UTEGwg3mer5qBBbJ9FK9uQF4aRm
mHp0QYe2vK+qlZbZFxQuHzn4z7pVt9IjWKEm+ZD6CkKa/v5U/9JUoyODNklNzrsf
HM0lRlq8ZDouRLL1og7lAfHdYb2+w+1IS7FuT3Q9dUTmCuouoAsa3LkizBgPxBgf
HrU64EbQMgJT0HiLJqxxMwL2IctcnuX7pvGRuZ9K5pzUzCM0o4gULAUptwHmQ+W1
DT5iD+ZqgYQy1JGbfeMbpAy5w7/9s/qlekccdS2O2/OmPtdx6yll39W1bD75GvEd
8RC6K4Cfj2wApSy4teaSw66McouMWgW0iin6C9QsFdy3xt3ykBcaS4ZwK9TMavG9
ce4EwZdKct/LV4UqS7xfjuZAKUFX1QpRpD5si9KrhIwaAuW1WNqfFDropV5xS5XQ
rbGwizIx1Jd9XjBq8vJQSnIumv5bSHelFJISaHJ0aJsIdZXt569NEOAvdpmPEfbZ
V5QbX1Y3Z1yZczXlOtDAD9dadniiCWpb7SAamCvQ/3ITgokur03aMLVw6EllA4Rx
la1M6PmYQ7Ia6dvIEdKZ1n++3FLKNfdlghIn10+Aho1sS0jhuel8PxBea/u05pUA
hbjXKSebexNJweiXORhA9BJ9DCmPhLuHt9ShqdqSCzad3NJfGQ697kGcmncJzsRg
Ayvoa5I/XOQGu7Kkzaj1kE7G0ZhUtBwGGLnYdfm0XtnZzjZwNeNguxCseUAKXzd+
WRQBLXHF7j+Krrrzs0KFEAtzl2wT8N2c3iyIspZC7CCRJH7GE80ZLlPtfcDsk7SQ
JME3WQvdRb12MVxWEQYui08pvkg0wNUV5JW+UbFpLQMSM52bQyZHJ8ou+ppTo2xB
WNJgWpCj1PB4D4K4EZzJ/30qajklbEe3x0Q4/Cbi2tz8bCSwSHM2k9JnVSExjk03
6zKZr2fICeNPSoFwXxAm7Ix+fHHC8gEh6TSzdMlrklVAloUuydzXJBpUDYSR4MAY
tmshyXIrNlgEU9HRPDlmG8cWIqJj0kZYZovyQWuQJHGpSDhhGOOvJs8kF6mqOATW
eemIAKaeHFuUJc4Tp3M802dUieJRgKb3xRiFsQna2Lbl3klM2wS/KaEC48a4JY6a
Md+Pr9WHsZ2w28/1gf4JlBrhJV6ElEKQfDWObSzVAA/eTAmwFO/+juLolBezpMsK
5KtKPlZ6gMOGZ1l9tCmTY9vkbqaVsOQtfsD9kuap5DVMO9IDU2VkBzniseIwVasw
1vtL5x767v7GxtrhEsyoKPAuURdhcZ9H/CMIF+swbD5tFqujkhb7jbgy4lh3T+iS
12g61vF4XFfVc31RZpNqHvJoXqbOjQe8PltkH1HZvP10NP0gRWWsNELq3rusJv+s
CrWCcvZ6pXGq7wD97zGRAPWB2zyG3eDXyDy4U51EdWz0HRh4fEmD0BOP/xMhhbYu
A9j2q2aRZDBa29H6LoPF6+TZaG+dXflSgUca06nnWROQXaTHzT6LqLfwmYz90wfE
ftm/kGkTMKZxyXUR/+PYb/EZsUdPmK9AwBn5W3eUhjXoNkFT9BYn3n4/DKbRCE0R
oecd9JJOJ4PWrswWXIs9BSwaYgevvPtiG6Bpn2c2g0owjIavRJaPEcLKTTD2hL38
gj9Gl9oxodW1BA1+o1Umi43PRNBBHI/KuIQSJo/Gg8H4jkFPeQ9PZS1ZwC2IL+3O
AH+3oknfmXIiMCzSMfHXDcm1gAJO+pSHkYrVxzjbohmiG7IiC85if+jKU05oxiYX
dBKkLvIAjDmTLlbJR38zXF0Ywzt7pZJdHW0bjfMmlzYT95XVXQ0+EcomOduFfcEb
56ln1FPz3Pd5rw3ijzzOMvqDM5RtwGJlJo0/AYpUjetpEGZyk8d0aUm4Cq2+tCL1
nAhB6l/2uuoo79XFsO49mzK0wdIdquKAVelOAOiZyRZI2DXHeXMLMvile5dpYqhV
6jkww8t0DUXLf7FJY+L9jWpEmy1PekZAehAUH6mqKtyAdywBHRmDaiuQHvCpdQLN
mRqrbEf0WSM90urDqwXTxeK63s+KzFNNf6ZWueoNyaAyYHVdVonDxr1rdsXG2lz9
YPtZzpheauTb0PO6ED9B43+ZUSNg0DQzNdLv43tTH7eyN1wFuS0uoBh8tQVYAyI/
jSr8THDZwNRwRw8Z+uX0R1Dwit1//Vxn1Lm4nUTHxjuvxny19sxyUlH2Rtag33bB
XKe9DTh4KzHcHyjtEOvpv8l+D7Sgq1gYMYN1WR0qU6hg9C4rAm6ZGcnGhPnWmmqO
o2HDcTH18AJH4NHLd8uWQCxHbdrCqVhgO13UaUiZz6TIPGP/7wmK03UnI8moYAPc
Jx2Ns8q0otQSQtJf81jY0i4QFC36Yrxxext0uOsDk0Zf4gmESIdgUZBcGeJ7JmdI
47iJFqlxHtYy0ZBKKYHxollcnRk8B+EXHYCdYeYsoeuFX/AZ7QL2N53KmGzN6mbi
RwJXiHUsFafJDZzHWj/flPFGrF8JZ57qXmFDT8Q4rMZqrP2uVf7/8RaIYzHuX+mO
j5ywTxXKzwYPCq3w+Qtx/pkPS1dyCMJcPHaK4cdrP9Bfkqq2X7o91CB7/L84b71Q
19c4xwYsAmfzZmDSkoezWf0E0hNuC1F+vNzXBFnsNq5hY3bFChSTK5SHklaHbDvn
kZdjT9ozby0dDCFEXh8cV8gCfKPV5kqCPbZ65+4WNrp9PwZSREESuztI9zrlH1QW
/NI9PNXU3tXB/RbqnRz3/FfNQy2IQqIRKlGcus918qJAV4lEklNfKhnRm4gGpc8N
2ruYZCJaRM0MsFo+DOe6g0Hd2t0m68BgJKcStfklBijk6T96DuH+NOXEfqCwUR7w
HlHvXprjGPnHdLbgmcf1BJKKE7HOY/ElzH+J9Cb4Miw6Q0R8TAvcDjYdLzZN/qYn
essJQFkS99sa0I+w4j2mh+vIxM4dM4F88dn7z53juXN6UfGjfoyw9v+pfX0Nlgae
Wu7ufrbCnjNRzEOHlNL1lJbNlHuaSkemQACadeFEFPXxnlyFEUU8ZdDMFLCGd9id
szsXBht3lrbWTg+/O1asXDzp7AL4n8XVD5EtGarsicnIydD0nuRn968A94cPsVZJ
VXG96k5uYU4NDNYYtDxKc4cpEo+cii8t80HoOTSPYBh6hrpqSEIgYOdyWwbcnIJO
O/ipYZaonVBEY0A9odNjiJQHYldkDvcHFntayT4gZsMFJfuSkVXEo+cvqZqS7wOH
svvzvka3Pavklccnsao9cKxSCzh7LfQZIvDCPhWRRwEYUhGGfkMcznQUIQd03OPa
HzgLQMJ0LHPTd3fDWORirknT3U/EAHxD76yun7gP8dcLczLZNsjBTQsmuTDxGROv
pugcygsQNKUoe5mCzQ+1YLGLp8UTe52Gg7G/lkGkW3CUOPEWVMNsMbWv9RIgqrqC
iay7w/4zw5rJNxNl2x+HzimE+sIX31n0ikIraj167EA2+4iNuxkiYr9quMTnbUgb
+zDoySga0KzkOlhn/KlXMT0OiKCSFfQZd3vKqJJd+zqBkCsT7mn6t5tnadBKLFVI
mfxIxj1gdw/1t/Px9Bv7d/JrjqhuA8F5Q1OAli9HRDIeyv90MwGqn8ctHNjs7fP1
hMUmyLy405xLJKFzY+nBzS0Lw7evLr79ccUnXX6KkhGDsGQNhZTHAS73CRomdiMr
JV76rI6P81jeu/l7o9no1e6rZgVJ+ZBSoXRXC03vUmdDHbPctiL+V9q1TpfAI6Wy
Z476t9wkJ87CQ5oScgplzv/Is7WQ7Yi0aHou1RbJYnhCVccDgy6LrG2UpT6KRB4Q
Vnipf/2CiNmVqVZAN2I0mAZoXpiaUgtrXSUkMGir+o4KJgME+OBuKAAauF13LTWf
Slkms9Jbs4Dq9XfRafmDwPBQN1jiktS9xFyETphSyUYyhrR3olBHHbYT6QOJWd0G
K5n7rVAwqKz9VvMkTsMXv67uM0hWA7sxuCr5IBMzpnrFbbAalGP/gwWXN5mhNZXg
V9Sdu+StSl90c3fVnNn4YQHP/N3/WG5lzXPGQbCZQvbNnerKVHLZg+JBZS6lwC5c
/otYaBbam3DMlA44XakK+ae3QtcuavIwKVnasJHc7JagOYG8EELB4jGnF8eL2dd8
JnAulv9n5TYLDJ+59mExyaGjRr4pbcXEXBFMJLsx5f1ljEocUWsE55YookEYtBjB
/re+CO+wBqwMN1c15j3oxx13uXEd+7xz+yn36tqnTg3UXotJzSuvFv4XZZ4oSSQo
Ns7o6k0EQ5KL5ohqCRJqqLVwOUpgnJlC3rnnZtK2hYffsuyELfY1pXFjTehBqRrw
DqXyCtfHxRJw25iTSqODL1EN/D8Cvbk1mbSx/VWmuqHrMmhdqKIwvgzYMhAJMgrE
KQsk4p3BoND7SCSJrr0mtvuKKpulJW287ezZayzBKiaKDjYGqfsIIxbqQdZLOavW
tayZNQk/UevxW5xL4GacSGxraIFP3oukRuc2opb61qnT5kXzcxbOEWBP2Ocjzrjw
UqCQlWEetf9Ble4SqFrT0vLWLrV36RT87RaElcI/+0K0BPebAU95bFouEYwp0iDC
PYcfW4C2tp2QZLfXyOMonp4KjBLsukus+HROp9SR1Xzqj1DpcUyCyDKlHyKwCb+K
VAp9MgiURRjsu6LluE/us3DWSDAoUkto5qh1svih3vGRhhTSlA1HUP0HkEDy/cvZ
feJnj5TxvE88gPgmp9PhRRT2bYim4SOqtDvI1FRvZjTBhdDuIpI9xwyYNO8YprSF
CNE4wLklSDYdlVAhT5gTV8wP8yRiviVcTp8S4h1F7ZQVgNQm329Bvb92ce+3JA/P
WG+Wuw/KHtLh+dA0YPQv1AyYSOBG14AoCvE9Sn23oi51c6mXsUZvTf1izStnyLzf
rOjE0tIdWNDTaqoFgBUYtkQtADHWR26+feSqzbac6DmhwWJneWfHJLpY/IoLxQYh
qW+GTCMIVlmFpbfDLWh/3K4VFQO8yYrxGFPYY6ObA8kPvstvk01B6TOPLhnj7Q7A
PS4DvNVw0hKXIzmVfT5khwpcMi/AWB/j03ZO7ANmrNElKEahwyfUget7MY/VUcJm
zqZAKgnZ9rY2gxWfiE4iBvlgLGvo+GaxDWtgxOROwWnb3caPgN1wQZ/SreS3M9nj
Eu0d3d5UVCEJscH5OS0/rPgBeJHrZ33FXEvhS1eYGHvSnIZLaApz7MiRX/TwnI4Y
SVtkVoTrkC7fyZ6Xf0k2YgrnsxHZ61iLO0yRoNYlWrtFPJd8towgUy+NIX4YctaE
ppZkilYM1j3piF/XSPjgSDjoebd9j9kWC5csrK5BlUi1Sr1IJuPcOV4uqLq8+bpE
HHzRQG5gub/Hq5RG049i5sY/8snCHdVPzoTk7V1Zs9xmZUNb7t778Er7Y6kigzgF
r8tds0ZZOScjBgaklb3xZzwraGP6EA4MlI1pWHGNtRaQu1NS8AmYer3tv9/DR8Nt
ZIAozE1i1dMbdGhm54pHZCEBHnlGtWiCKhiSjReX+UEu1v1fqAf5H1Dlbm1J0j+l
jape1jNpsA5RIGc0eeiERvwIEodhrn3WAFRdm1jvUZOl1Fpef7M4DbDndR7QtOtx
9Z3WLDP+qCpF3F67HC+306tO5WoZEnChFquGY2mvXNrTVnjzzZ7DoOremxiW6h1y
btzsatp2Niui/6gHbmDF2a9E/28Jtq5p7zFmuFDEiBB+YH59KhaQO/kHJYG5NSGZ
qCjDTG19OktF37tsglE5Fvd2Sas9voMTdy7Mv6QwZR50TY+O8jkfcBBwykxy1nk3
5T0tUzAmYj825ar1yGTrcrRibclKKJh1uyPsMVr0brogCcrfCXK9F+rAmzkk+v0j
R1WDYvpnu4hrtfzl3j8BfoWQ3UD/bY4H5/oIR893Ym1fpzGKJt8EvVevOlR4Bad0
/DuUwKOzjWQliUn3bRoZLay5VGB4B3kVw77jLvaciXuNxASswMsioecrlCWBngk8
o16WvDpUTe1Jyc2ylU4UQTSNUPCpH3IrAkbJAPk9ZVPevCNeZODT570+mUyTI4II
qlh83txrAhuYU65qQoTTSToW4FpB9zlAE4x9v6nTBQBGtMYjLli55vLNlq3215Ot
HNuEkTgNwZ1PobBGhVoc5o3FewZChuO0L7eKLdZ4q/P9AMOCcS1qVQsFif9dtdDe
qe0jhpWEQ8Kp9GjsG+zb5x9FAsHWPujh7ACgcSoAQ6l/whbDMUMWOYOXt7YKpIia
7eoPb+RFs5uaF7DhWeUheQdCJoizrdyFvoLjeNCm3lJ8RY/vS7MOnEYDp6Hnx0EK
jgYgK/eai1ESnRtcGQHCcyPUx83BajUfBa7WjFvBtAd6QushnQgcfmJqKzr62Nbm
0/QTg2S5TiwyHui+xB6t9HqhWUGdsothDSdKFVY6E6fllLyD642o4YRYjJcSigdF
kBm4P+SJqD4qtOVLJ/9k8CwrinIW7MNlR7irgv6Ws3lZ+fcIfUx+fpuA1+Ew1Nmz
+mUwWEN0ltfhK/I975PKD5OtXJX8m8V47B7RDZMKBERT8gKFwF/Uxa2IzuVvH+wZ
LnCEcX03ZDMsgAgPtSW3sZH1vKq7wC4WMYcsdeonTkfIQ9/c960cohMpqEsoh88w
h02UMzKCZPpBQGbf3Q6Z97u5u/uF7fMCdl2qTF+3DzI4HTWw78LGOO/QHNiyiCF0
gl1REihT1JehqkRbYaHVpuKRiRi8gdvrwCDv/zDChn+hEjIpvPV98sztldtomNLZ
FGWSEjk9XEr/m9kuTSqJQjnOwvPE73RItUlIqRb0oQPcP8IFXC52k3K6e15axNFA
hSomls+o+7u93P+FYUtPFD4XZVdeMHYq9ASQs6CjbWUQljK554X3XjTz930/oh/e
KkoXvK5Tw7v2TZPpxajigSH0JN732fACZ/OT0ugLAbC50Zgmkl6oVzY6jHadvtXJ
tKsGvpfEJVnsBa+VpjuueGJaDrZ0M4Pny34JvnHdKmxVWQP86C8GUrBNams/Pss9
KImZ/Ei1F2gXsIbOUp8QaMX6ZSsO+4Z8vvDWEJso0d70Zh/JCEQFn4wJ3EAGa9vu
4CegTLgY5NeAbQnFsjVA9s5coWvwi5AEwxcdBGdj2DDDqtf3NYSLGrmjys6f23f2
CTfPK3eq7zcWMjIa8Tn4tQUFCJbel8wToncwZUa48ztRGzgoil9OD84DiHPxg20K
M9PIbhtqcIemvPev10LlyfaAYZRhPdwksk5ukIakmQfTH4Cb9Xf1bbMAJzA72IF+
rDWHbFEQxnyP/9raa7GTMaChDwE7sVMWA3D4K/YJHXDbLk/AtNzKUWrDWEfu1PKl
rBydkJKsNAQiFxyp8t6gW8Flp97E3aoB2OXosvfgDISoAs47DV7/bUFYRH9qj6DC
ngEO4ruXivheS7qg7l1lzNUMWTNpaytB4j7CIOo/+qPtQ+nY+x5VIjkfGeYVuMMy
XBxj08QAIieDuB5nxSp30W1eoviH1AKdBm33BtK6wT2xL2BkY2zZV2e+C7Gz0Ox7
vByVAzjeF90b+dcdiGSXXpR5BfHarpE7xXU9SADOaRYRHrr2gixI3R7oGRR9avbV
j6KdM7Utl+UnGVMJvbl4aXj3PQPWTo4FyanuSzqtSysTb6mjE2QHgIbfLHNhjlVN
pqt+5RbDflE4NpNL92NpK47aV0nYp6r8F7hZnaYG1BH2lY2a4m7OLBkadON43C5l
+49e5L64LU/xEqW4tH/yGZB1UlSFhBF+/iXg1C1/rzJqC7CHuCvocYsIwmhbMD81
22v17lCln5Kikh2OKxd0PiKn/XtsFT4h3GmmIEucw/EYTO/FqOjLUve+G4zSacL1
gfEL/MhDiNra9b9JY9ZYNlXQjyNputrJD40+Mp32BUr/crQHOGiR9hxbCRzACS7x
BfVpDK8ixTi9rCFtSEShyHX4n9nsE4Y296SZ8ReOp/dWoahAulK1Z8hj4Sv7V4da
DpmUwroOEzamCP+01zs1Lv4zL4/9gJNI/1d1QeAjr997CbNrPj/txRjfx6Q9Clze
C1BbBm2iDyjJ3xpQFQiowgkOamqDcN5dLPFrJ4KqXBm7NuXoilmsk9vuW0r0i9LP
pHbHkdKQpRwkywWkinZbUQwBAfAPqYOBvf+RsKszdKyyvjQDl2tbkwAB8keMho2Y
pOepDsyedPxBCJ4AX3prcTBA7+XOn4XByXjRUDcccupoL4E569jD/DceT5t3f9RW
dOMS8kdq6mkO7xCchMX/vUmJA0fHWFGDx+/SR+xMmkMwGekM/+j8s+wAtmXJxv11
UQfg1RLxPuMhw6FxUWknaavtTLlg4DYO0r9ekHEnYQdhJc/On7kSZQ0oNiHYmvKZ
324Rnc6ZHyK8DcKcIes7nqlfOzgVaPn+zmSCHEvZJQWKxtxphcSalO5xUPDP3+XF
ufeCRCeSnP/aNVwMzmV7CdNZ/CDzSkMZFb97i8nQ7BSK73kJW0CRbI19mV1elE/D
TSknEc4A3Rr9oS1R8O5/Ofrubhpo5g66IBWukGuOISuuDlJaYqL6LxnNUWceBq6m
Sb355kYQxBjE6BQGiwb5aQ1eJ1bSUSbBkxHuDn2OJvBNgrk6CLuIOE7bj4xS2doA
XjiV8JRZYKG76Ygs/qZColnTUI9R99g1ZGtOuZBQ+bk9vBmc3m+i7008IdnoWm8r
zM7hZtu6DQ3mc47MVIcmZUEX6esEhmSaGzIFFO2xSt48iLdmip1Yvb1Vg75eQJkl
o/MkcvIrVLC1DuCbqNqV99ITcMqA2QB8uWTQRPflFAfatngO2Ko9JRv9SqBicF4U
3roZGyADy/BuZ3t6pU5vea3xkjTYgdF7OqXQm84ePc7DzKdJ47oJadXN/bvLiImO
JZoh5vUGf04knrKshm7K0BiprUfyXsNiyu6cPPNsV4eCIl2urhQjALGAvlneg00+
lhLCLG1wNUbN86wx14ASqQ43AmMDDszjcJjTk1Jm3XsrAhLSbf61TCRn2eOyf9yh
1P7LkwMjBZEbpN9SnmLBP0IGrLe2bB79q9JX+eAVLAvHikGKgCo/2oZ5fodGoAiM
FW+VQjt0uxcHYI9c+Mx6SmsFK10aqJLtmsnrLjUAFhJ9fw0ojjW2Hp2Rsywn/Zgz
BZLa3dtweG+4jultCV+kxEgIiHqoF58/AHWvc+TgqK8GsOEFPkoqsmOv8wi8+2cy
l9D5PWSpQYD5KXIi0DiQ912JyveVnVKjT4HzbF/EURKBPdUgOXCOm6WoGVlzbXq7
38vltYxl0L2VDeeIM9ItsvValGPEwyl3hWwdWhdEhf2mtqDkI9tikP7pHxCdEGpr
andwYt3PtLFBp2E/uS7RfilgMtA4G6GU7SJYN8BOTqV64I+KioL1GIOCLT5XaNGa
UWMx5hZj00Yx9eJzyGiUUAf/UsPl5kfrh9PfmgTIs+gfXrAj4fYMVgfK2sWfnBah
EJxWLbQI+KLwQBM818dZz41NJullUVtAZ+5yxKd7vN792oR3w4Jolupx8NtinOBe
zpnjrzTILxY2P8bC4EYMvGWmeN2CagVZwCRBxnqo6mkhvbz88tsMFsil9ma28qTo
bvkZjPgVKoKXVH4Q7Py/oEizKthJnwoaEdGN/dBHm5e4gDrGdnmRh0mw8SLTG0yD
ljPPNOlpnsIUxVvIl+jTluV0lOSFIMDdcaudCdnX/3gUEHLaeSxOBlsirYVcgLvB
RpCnn+l/DBb3Qq3lvN9Bh+zR8mGZore2yMecJe5kBa1Y5EyW5fidCdHRlsgfdbUw
GdWC8uv63WdSMV9oiaEuniFSLBMqjosKfDRhhnU3SLGwSTI8l84UsvHIhAMnsgpP
Wu5Ew+ZKyWOl1Q75qSR99LPfbPAFZ06CG9+o6CB6WLnECHg0H1c3cf00ErBRr13P
86k4UncfebpNyyB06MXSJVCeo+mECb4rAXY56+jcBTsQW9LLmsP3RaQuVxsrL4+Q
WxisTIyr7Nl1t48SeAZNTt4OvWU5sNPoKMEKmVSq4deQrtV6O2u1flr/Tg+5/iyj
hZqlhMmSSp3ut8PfZ1s8lqH4YnKlvJg/efK0iv6mShbW3cqK3kFdYqNQmDowdVYJ
GKvycv8ns067u620pmuajdTyIK1+8ZCgMRwDPUBQgfXJTIZo9HdRhXRh1snKWSRa
h5/RAFKSTKWomWk41Aj3aJ6DsSXvrPk1Mx4GpY52KXHrgXkQxyl9e7CO/ywAgKU0
arQYeBsHMP/QTuiODS+uWAarrQA3FBIgjHl7uCzxZVRSoah0PPeoJAw9WBgWDTC/
z0kPi6flGq700OliG5HdFPAO9hSpKTImxUi/Dm3gPIou5W29gvbgOCab7pBUuS8g
h+hsz2ZU8ECMiYborUBkUBFOcAypvcTdphOvQ/QEnaRxv4ZJ2sw3C+EPecpZ9X3j
/+n3vjQaBsqBbnAtGyrK/i0NjeOiIZccS9JJR1DJps56s3HTuA7YcfY1fh1tyhAI
hI8+qyVOpAsG89nW8663gek/KwGAERFu46NnC+BjctvwU2TqneW8T2tABQf2ddIl
e03XZJgBu1KljAjs+/6Rq25elqS+PWs8N7WAt3K1i2d7uDGxeJL1ezA3ykW+Xi3f
2bbfdjUn/GixnV9SjkZn9pUgckrPCtY6fw6rFUfhAkNDxwkpUW/DPmq9q0ej2vnH
dxuWIwW4HwCruWIth3BJwKHZqE+aSW0Twwk4BpoENfcZ4bQ5FBv8c6NYF/zdyXC3
WHeJxlzS3mSQpUVQogDmafcYQQ6IBSrtw+8+SUBNcQyScWHAb+4AaF2hR/zEnGii
jx55SxEqJfxfnoVlTzsWDqfhHNsi43a9mE2mSfgI9dg+a8jUNujxYR7lKvUTgkbZ
qP1QLuPSu29fJoSLJaZ9zfZLvednVc8BPvCnXlL+Z8r/1yB9ghKigu8VWxzW9OPa
wua6qwihwP9vE014BC36m+i+70ZneiEQ8nGJIn7xluecwLcXu4LrqC35LwLJFqwe
i/LFTRLbk0niWRrqRAKSczsgwie8BPPW/UoGmJMYGEXg7ajfHqwJs7+9+cRzAUpC
g4HbCKQrcXBDfxp6b1uck3pZip6yt85d1b5aVuRvKpcI7AcRf/t2cgOwh6qXGHbP
SnEEyyjo1LMhzpn+QfHyYrUthVSWzHTMEt7wpZrnsHQka0f5jQMrdUc5nHtID1kN
KYiU8ugV134SS3FXyQr5bjXQDEwAmL4fOv1XWWR/nPVhOxS4LegPEC8I0iK0cky0
4gY6fhxWRrovURR8lkXfqzBI7s/vorAVHh4ajIjnh+kqSfhsY9T6NPG1v4WHIsdL
vHFbylBHvqPwmfc5w0vQp+QH+aG5FIjI+lDb4LPNFq0lHun8iMNXawB02cHd8fWh
P0Uv311bXy7ezpYzTH4h7anTuYwdZpUik6BgYgPYVQsRwly4cCngYkJl73S++NPG
biBn64Wa9BfatvXJpR72DVwIm5KxD1TV0enzTYAEHqrQooFyH/eLuY1Fnmfplf3j
IBr4szp0LEF0KNUybjDp01vkNGDM6GfonF8DHbtOMfzdlqsGZvQPLhNebS55RA3F
1sDOTGtgFuhguGFIkdwFX1NjOzuLQCq4zdS2wzVRc34EMg4XBXioVue8cTnKBloM
EfS91dLgYmWq9QtYE7vKsLqaBTUBE2xF2Z6E2H/gptsNPGpslSE4+f+X17Hdt1Vq
uPm99OlC926VZ5Y+zRVHnYcYEq9dv0cJIw9EMpi4xtnJm1nZuduv/DHKVuU06kDM
JY6HnYY/c+zSBifZCAlZl3+I5ce9tPsbMdE5SOmNr4lh+yekwcvxZwPmB43l392+
tKibXGEtmbWift8JWQukzMT8lfMGSLFcmoLQgC2/r9OSJqx3Utj7MVA8EHV1uJrs
ii4ZK93Bge9kIpSyGk5NlEfigjQ+c2zml0J0LQkxhd1tNFloWgph++f+uSAFDozd
A6EPat6ms/zKL3A3Y+xlOh+JsdmuxT/BVFqobIsZjTHta1eRkPNiYqfPpBEAmexn
R7+y4f+Ykr9FlO7NhOto9DsSDT86VOk3P0ZEy91Y/v4E6AEJTNMMQOIrLKWPv7pF
ROnYX36cheNDt1EceyzzGbOTuBGlt8GAs0tYKQehYHqXKiEhkumGXGfBzJ2gk758
c/MRalcb5yZVywzIHXDNa8EXlCsSa907dDWU8BAyMo4ztHtATmmX8oRF6uZzRUro
WgWZLAllG0o9Nby8jNVwqZ3/SkAG9Orvw8wS5U9A8aL1MeyU9wAjCOO5Zo2vVxTo
SVPhBxKXk6zjqWKBqhz7KlUoAx/UsJKUnS3SvAICwLdIcCrfc+FZjWiLyBSI76Yl
LUWb06tvSQ6XkbqSAd1IMoBhg/kOHTRS3IoWl3F4raGOcImZ0Bd1KIj0NOgteHTC
Mc1JQ7sw9q8Zc+bKTDJkM/us86r3tDdQgQXlTEc7+lQPrl4RwVLJWX4nZjxnWPVU
6at7mJoGChenl8FVN3u8nd2BbrZI1Jsxx2DKwr8at0t/UAwyCB2U9da1ulOgWmaG
oKrIoipglRsPGlIcbBET30VNDGCxi1clr/m09ab4ZGkEDgBJdL8G8xDA0SNFM8zL
9C5I8rlNohnduM+Ye5BCuFaVi4cLFpx3ap/joV9ChUlNBvLD0Htt9sBY7rYPJPhM
OpF0Rjf3bKfc31VWBQ8QtxPFtyYe6VMLuQUQTIiT7JDmG3RzatFHvkEdnT3b7p9j
/NAah6fM85kAEi86qJDu/trQ5M2aBQj8L4aDvv5PTIYwVnAbphokxuyex0Tzobn6
UMUlggvQGyQno0X2nG9HD7r8GXimieC8htImCen8jGm+nFcEvCD10dvnjkwvsaA7
EOZLtSV/Qk15pS7J1En8H18LzcFUq9AsLBygCUUz2kREwK23R0r3FrNmGSTbVyEk
C68ZwMmsr/nCTiftP1gFPFgWYK2QzYpQYXNEzA6LpSfI70Y2Vh2cTuCFh36Jfrlm
B/UVr/zNvosuoGp0IfSEbysGAhvx1pDXzQdsCkJIKOyihaDbAlie9BoJWRUOCtFS
eLHJR8AGx2+GzDuMUBcynFabDkLaqZZDZO5TZRvJ0SxU6JzHcKF6nYnSPuDjbDLz
i+mXEFgsYW711LDdZq32vegVv/n4OvDpWLTk5f8TNYeAO98SN+j7fM8ab7miOoc2
bmNSA8YvV2Hf4VU7L2KaIzGbcbFu9MidyN1mPvfkqYUHeOonc7yvyCuPjcALzcSe
W5BsWRqmnds8mNkmhbBeyOUhTrqcZiDMIZK1TWMeTmQQ9MAH93tjNU/VdwjuOyBi
rv0TOpFbYti5sTPgcMldFNmLJPuoFtXNeC7wbgHp1YAOquO2Gxthx1OeEBvqlauc
ryphGPEhqGODFpqMTwIshK7ixhRjtH6tMK2CAERAgQj1ZSgdkHXrVFpnmknr1O+a
nWAgsDmg3sbstCFrD3UuSSF85r8Ym7nyRhcCI9Q+wJL4MYuMehtYkNgck+jBu5yH
VKcHy2rbq5r0aK6VxrBESmZunAJEhcESPbPFzifzGrKF3jusV+tbsBehyVvX+vXH
eY3VfOWej+5gyN12pmfcbP3teFbMNyu9Dhz/HXK0RF5XsLq7hH/yM0ZywttSdoXN
EaeMcEkq4+b64T9nUj1D1usj6jZgw08h/nkcCs2O74Ly00zE4iWQLbJkTaP4DBqd
YRtkeRta+MJPAUaXi9KQLJg1fSJcKxIBCXyAqCxAjJ22U4KLA38Di1S+jPrux0QP
mfKp8o1JZCUaNsd3P6Se9RlO5VaGncI1o4+mEBytz6oWVrGLmKycUPL7jzCuLDya
afQBhZWGMegTcPGqHRD8kcJ+zhHnbKsjga+tdQDBWmjYwzAotNKEQ0PQME3ozseQ
AER/YrY1w77FRaTc5b/FxgIF2Axgw8ZDhMJ4BQT9v6QeXlmVJBjYk10ptcm7q1Vr
bfSStx9p51LPCRMZbmJd6VW3J4t6GGIBrLuzlpAcsTexkdQNLvNakNHQ+7E/pMiG
XMpLniDUfLfT0IKhKXzX4Mk8bcH+inwnFo3DdpnDQ6D7gjW5/n7QZ7iqxvrMuoVD
od+arr0gLjq/o+88LsJLxmucHVkTF2CsPaybJRZjVZNdhxaIIP9F3+YDldyy8b1M
nna9YFNOi/CkqyKT7osEW6BEttvj409REYqeXrJ7aHhou9FadvPc2eIitrJh51oT
Sg100FRXXsD4pRGI2GrDxQIqZzdO5EtFc9qJya+iowv9U1e2K8mliooIAsrlUrZO
iRh+ZdIOQ28ShN+WKuMzq+37jsLluglhYm1VFOANQ/M2rbUz80LEAv8+E2D83UFg
auBLgWetnzJ1w7OKrujSrDX9Gs3LWVu876TP3QDT/6VXNX/iQx8y03pEMBcohebc
mkc7bLz788skVFdP1sALmgMp8IopOBRvyJT+SxyGJrly2bK7dIrY5SDF1QWX5tmG
GTT953sCpIZq9sN4pIL254hGsGbsbb5+CL22fZsiR1s0qIeL8bRTbbfeIP+pNJ8G
StjFP3NxRrEUkldtB34Y2PNPusdhz5ieURes5cMT9JFrY449OyIOCdgTWep2D/wb
otFq1ikOTaa6plr5VPPbcXOGOqJLH1fg0a4W8MEGzIeF9QougMi9csjVPyBZ0T38
U7Hf/NLqjfL38qjZfJYevCzzNodfp6TcRJpHZ7fgKxLbX1m5gjTuvG3RJjsS6aJS
MHz3/oU9JkSNGi5juKKpYGmwXV5js2WQ1hPjgAA25pDG/ZKnUrq2pGZX4pMH4c9C
vajKlIZOujPMa4c25H97dm5tXRlJESYjuvxGv/2loGVvMkaRTD96X2sUkwKx+fWv
5B1IcAI3BzIo78QMvL3m15WKyUkd1LX8nC13rpzlgFXGGpR/lnVm652J9jxZMbAB
hCGq/LjEBVNCCo+yHc6afjx6NZ6LoAB8/i17ipFmof9dXpR0iPreSGF0U6HkxVk9
+SPHEWDlrEk54P+/c/TbGks7ft4cHpej9d6+Tzsr3FwBCB2JeEfr8zoh8EfSNI4L
6AZ/NlLMpEKSk8yggljQMlG+t+pucFT4vkWPf20JCj+vOefzUo+8TgVgO6q3Qdag
EsyZWMqnHt6wRlpGBDbr3+0kIewfb8yDH5EKBqLpwbjGWpIvtMBnYnokCSZjuJaD
YA11Om4vIEmKB8oPKWGLjQ+nKa5niNlJOexvJoZcwSQn5cIKIn4RHDLzopjyDKUF
dX530Lxoo55IOqsV1DAUYodL4T6H1qPUIvIb2b6ygPm1nD4XnfhIK9YwUtO0HaH2
819WvRfC5+jv2tqXtCTKYKOU89IBYxBO2hD0izW76SEJx95toG8wYuPm6xWlN3aj
WFggTO/J6+0t3Jj+E9dKgVYdT0t0z7dPjiYcNJPrnqED0Om0nxcq7yoL/DoX1Us7
v3QRYgqpksUhecilpuqfBdam2p2P4HjI9bqKraDgWOFriiQ4OwszLkgtJMr/E1S6
tz2yEJ2QNliW6OmfHxjzbNA2w2g9OTqn5ThXDyT7efdsk0LoUPHjJbGZmKmAFaGy
2b6USD2pE69Lr+W09YL7QrZazVmXOamAf6pIPV78Fs4nFMHd70DFADM99ft7Z8li
SQxqwE7rklw9TSBiqGW+ty0FLsC5I3eqQho1J63yhfWOqhdPECjsv4/SkKxJ+gXe
DmzNhQi2aC68XnWzxgVptkopTP8Cb8UwXfPN6IQn+Sn8OdwHpr3AiRQmJkQzNygr
Au7GA61HpI6I/2RApjvDm9OXU2hbkjAjSmM8lKudrrhlFTGKC6eJXcpCbdE0Paef
EDvpZ4PXPaz7q49b86Ya8G/kyGOwuAKncqzj2pRpI0Mhfl1gobJ+Sa5t7WCr2W1B
iA2dZo41816R0XR4c7/odgQBHCqnxVLIWRmPee+c/42En1QMoBtb4Axm+KuQp9aH
0ndbXUzVvVVC0gb/aCZg56AyCzCGt0jcMV1aZOneNrbYqAA4jDUQ49DZqvypsqGj
3wvsSjEosK9WJSfGrf0aUa0xxubDpOmCTB2UXF2N2K1XlnLZGQGSZxZc766M8JYd
ubKaZLBKbBSYe+ArgSjjZp8UbQfcJu8dlrUCBAadrvbZphdiLWG7Ly7PNKYPYo0Y
UgVpmnedS84MA7rBFCJz81MsQUBV7q+9ZTmc7S/2jKL1ApeXq+XSaGBl1LXSsbjF
BOcscgTP/j2ABSsnDn+tzpRqEqAdy7PGPbHZ6YWQnJN3vtuv5SOxBr7MynGToRB5
2NAMllKnxdNLkYQBz4XXpINgueGtK8fkCS07m4yEHivc0pe+uj+4eoxj0McFE0M8
7oZTlXpX0QjICrvnj2foBQ4WF8PTBilSXgwbx6HP9mkEUE7ctiL2fbfIM8QoFevK
i3TXDjoPkglySntyR9Ez/eLkOZ3BIFmNqxV5tqVNpb+2Jo09k5fEeabfTQxshtUK
bWh3oTwIYi5EjQjahFiN9gV5R6Il+vqPEULGef2p5yZuSV2Tyfxrx7v8yAAVEIC6
zCDhEK4rymhMdzZb9mwpqPQeSYMi33vwqogYxJ+nKGL7v6AIqjSQVkBKpWnvZSdp
7WM+IC1s+Vrq2xmCEPtoTEEfBSisBcDArGwVhvpKvlIHg1G0P1TB7yeW5j7EqcmM
+hvtV2SiaZw3n55d+3nag9a6Kp0HbfYc2UirRWSCaweh1dnJunLXXM6GJvYxCpzO
QliuyexD4Cl4gkoaCTpE5GsGgTfoW3yHq7bWimRDfCeInlY1t1eC9/QxZhgGY4i0
uQ0H9AfA5h/gRcH+FXx8ywZHOWC+S8+sWGkCBfpvEAepwPIyZOSSoeyn3GOv7AlC
1FVrDD2V+kB2H611NZsZ3UNSTOLUKlUB73yH0N1rK8i2FXW9wtuwVkYbG2/1J4V/
HfSa7L32rEHxYe6wbQ9TGtVt70Twt2HSQ49kxxGzqz9xU7zxyrWC3+NF+IsHZMl0
fbBNNZGevTk0gOzf7o/YKciSmHhsNGdLetH+/OD0Kn42BveC5hYjtUdgaE3N6lli
1+SrsyRyFXy7KyH071yFnqxrBFjSR0Eav43in/22t9iesO+BBVndJZYdOVGfxpJ5
QdNIBboJA1oCDB08Al2IFo2QGth5obNFhw3HaktNVU5vHym2RvLPSoF2SraJmoOa
bEAdhTn0kTx+nyPkDw1LmDl4/Ii7PFzIrE2ZxIIZWJhidkjzOBRjiLHG8Dg5h1iL
hyoWzq39lc5cBAc6TIZnbf+kxHY5m48EZFQl0iCJDTDrhx+DcNK3OYGbxBF9K/sH
cPBoRErFo2a/eDokMBW44+VCCKj2sMnI4qLu8hJ3pAa2SZ0x1frNgL3rDF3GTqiB
V23WNu7WoI6gq/U5a6rRyxs4nGG/4S91Ov0d89Kr86fhOaisr9VfUSz+Bf+Akfph
Kk4cKXSYSfixZ9fzsdkiicTjtDeZN3IwT7hYtjxUXyw0ZBvigDSo6qT5fGZ5iFuS
EeFpBwL6NF88dZQinz59zv0Zw43O650J+vIQIcpzVAopzNCcA84xg4Ne+QnGGxut
Xl9eAQZqo5cnsMTnp8/0dCinE5O2hZrjgjF52UJ8bNb4+fZj5FoX+7HPgE987I8S
TjqDOuj9CAUoA97/4UNXRz7Z7GI88zrJwfE4xu0MKKYpembwwxgYbQEJdgHiAplt
X7Zs172ZsS9wZXxGuSDY0gnqHiwmUj5pLvLy0KPvNTdpRU/RqDGu+TYuU2giPpEt
LII2PizVptRvQgumsgQ5/faEGQRroPOBbmq6oJqVu8IdJ/sOprMd0jlDUIBbRFxR
v0vcghlt5EjnqVsacUTXkjco0UQvdana/9BNJy7kwmFM6O+5evolNDhnd6Z0p31T
zLx8+YCfT9PWOnrk4pDGxl5H5ZHg3rEfeC08JwN8cif98wzIA6ZAEcNooknNURXn
O1PpTZnCkJGFFMufr26PwKBBDhf/8Zm9KgFAjTEeVDYKOcJfkzvcJMc1ZxhHqufk
2hWch1GxzZ6aXWEoWCE4VHFWMkiXa2utLNDeRUndXUnuecX6GCcs4UItFFmGu/n4
iwhQ3f0wBzpjs+3NkfFwIEZ5muCh9WKxPaRgcY2PiRurFqeU0amIgWrfGUYuPqEo
1FVpm6PQA8pBauOJfUAqU+C2T7BruLJxd826IpLVA07Umqxi62GyD1suu90jeYwc
WJFKy5XMQixatZsdr4LUUl2LLFU8upJjc+2i8XNHqz2CNDjM/BDphp+0Yl/XxSAj
GGZ5MgSm84AmjdyJGkA3nGHjtM4jjxCWZtWNeLpqjXvXX+qsS9FGozmuK10dnxRj
CjIMzP7W857uCBfVKlkGf0G1bie8f7UIaIDlPIgbUzZ+6dZnn7cKqneuLr95xEBI
+t4F7xGR8JMxLsluBkJsilxFuixQmwaY0y4DCmoUkSnGY0B0R6fRTMez0U8FJaqi
YdegitHxQWFLpENHpRG2P52gik/c1/ZBLzSG9lWMCJLRuBYnNv1B/BKJc7ELJBEv
7AqRkA/Eqo4VHhSsVf4mI8ouGrkE4HUiJMsLy3b16h290kddMETzOByX85cFH4UX
a0RVy/xajU4nwXXN2D9cDbjUdjyHubCGOROfgtwbYCDwU/g0qfUhlMNaubYbYWet
wdBfOp/rFaTX3R3HexE5qGp7rqxszPqR5GANll2+nPDy9JA/BW1rJp6J3dpqOqWP
l5CoWeMiIw0KPJVRl/7Cmsj+lW8wvVNdveEGZkXl8Y/UEbS+O4G1mD0vhPC+9ZDm
BVH0GJvuGXpUjcMLMJ++Z/XCEiIzRexwFzlj2MXl/oz9KFV1R494I3vDoWm4jR7T
K/iuYxM5lyN9ooups1e937HsBkDca+rdY7CAChJNgQCpKP3L62aWZh8eAq8LvV1W
UtEs6Pt74CTd8HnANZYWp8zHgzGKeniGX8ZcoXCcGNtY2yOLvYbLoMwi3NodTYxz
k4BpulapSTdChvVwMKHjbcEp/qTYzyP/hTfWh2sBEkikQRhhEFeRlF3C7J/qmCwI
8F30LP0DHtuBm9ZdEdJQsm8lkfroIEfrMPOzURPWQFzJuv6Tn5zDZyRDDKbZJ4Hw
qvuB+ZtCUvFRRnFIAZvnzSPS4rRsfYweNUA5Pgu2tsbd+E+6E1tjlZWOZqKh4KHa
XIq/gkbSM9aQf5STwgAeJqNRBYHeZIfkybvX2X2HmKtvw/r2dOr2DFg8dhnS4qjg
qkrXzEWx57kbhj7d/WBgJ/8FoGACv6hDFK4kv3LlfAG9LM1j+6fVU6ch9nrpiF3I
iefygHjnWtLDnXe4L+uFJpqr/qbZqVlcfVL8TSYtnMUJ6YUX/Y2LpVCctJqwhPol
fvQizf7U6tQPIRmTKmmKDO98t826dfuLLqxYvUCL73WO8wSffRSc/qGsomgihtpI
sGjgZJBr89CKLhLcVz2lrjzUM1ER7Y7f/dngFEHMb8Fa15DGjQvHKCcolfijh3Qq
wK6aF1RM5hFLE1ElmEQ8RCaUbwCxQ90ZOahLU7K0aJ5FoenYwhFhOaEge5jhXXXR
BoiUj2Wc2FwRL+AT7JccrtqYleJ9QsfCR0g8eFDPw6U3a8QICzD6ApOEd57h74JV
UaojMB1LY8a1pYNfcM6LWTBSIOwfAUFzbPKeuuf2Rz3j11II7AdnBDYuasJrVn8l
bRi/PI/rwIm5DFwke489sQthjCqNwrAcnzoTq2t1ebnLeWrxt32FhxNRV4reFp4M
2Rnv9mor13NNHI7i/p2xQAhg/eZ42d8p0eQ98n6Oa6byNsNsU7UirckSQS5bIDjt
gBPd978erBj5Kfan0KaF09qSw+34lCjfwq7z6+gUFnWQooDRFsxqIY//VGyx4bCN
AbcZWddIVtdfwTylMC/H2K1ebRucAfxMlPHekSBqcGemEamORek1PeQkGP/48b+h
m+JMzBwVj2QkbjuE/vw+BVq+nHOAFcUlx9jfoK/YMMcdMMWDLymFYnPRhoivbX07
zDCBkmuSSf3PKQB3hBy8mrPbqyAxtM0AHWB0ymJ3T9atIWO6j9huepGzKQieHoMj
MMmdmPmAifexLh25Ptp/aZ89tKEdLfNyKyegE+K4khdW16MvYI/XloVRyjCMhzUD
Z5dXxKmoTVLTWKKKOCd9X3zmKWQTxKR++bRpZ9YBOcR3pVN9YQpaIsvnP2T5UNLo
K3Wg+nSYIAXePD4NAIlymWFt6KxgN+eD8Z0qA43UK+NYrRWiBwY1qD2SKHF67fl1
+tsOgraRneIHGXez8KiPJXvI8dyirvj92rSRvupNwipDpeHeKPWkxJMuCmyvvDiV
9qBEo+aEpjDPQIOPxtaqD+L0F5NpkbH040OIDeal3d6EYWVm0QsFfWtuIm+M1wcE
yf/E2KhMmjqSSfcUxHMqEKVDgSvCbW3gar1GSqhmw4sQxr3JXyX532UvxFrIII76
8DN0ychNbb+T6kE/ef7Aoxu3IRToDhRw714+iaX9v/ih4RvMiAB77/eCLUY1Kpkv
grxsubBWBP+sDK/730VuJeeH6/OQtM2goRPkNmBfACr5/xyNKwhuTqu9JArqwujD
GyZTcM1KihAp4K7q/WpveJsmhA9kJyZwGwWzp+1oqExNcp94Ah4PgKhEiDlNQWPb
TIjgWdJrdF1Zo1ID1mVGIkmpfGTgDPsz/6NhvPw+fsRmWPJkiQcK9e318wZPI4Tr
MeNlQCHmZfLvOHBdQeH4okFAEf+yxjzW1Xgu0kjB8VPq44Y/EOf28pF+m5ZtL2cz
a2D3RD82b7btrZUthytgbY8nYVXNuAeEek5QMQYi3gGP48TPPZxneloZilIDImQ1
PL74CRJeflCs6Y6YnS6JGJaeXiwBQBSMLOZZHM0mUjvd4s8T2SkV8yu1jiaKWGHG
M2oiSkId3rIXMEzTzXqPiHGI5RnnHJm9K4ciFjYs5nYbgadH02PGLnUAXpkJ3YvK
CaILA8B9boPHOTvmJSqFOvqzcCCTCM8y1nRuN3ZR2RcHl87+jbCLcK/75giO7Mrf
XEeGE6hgxTsqMkVy3VnJpdKD3U0dl/u33oQnpxq33dlVBHmkBYoBbuu0pyQPGHl1
Ksrrd5DETD0MD/T1FWGBh0CJW0gkvrnkGxFtaby24+HGuiwXvQzFPkS/ZDvezAC+
erofZ2YJehe+ba6mo/ugYDf932ZO9jEuVzBOVTrGLFyzmH4Nmn9kPI8rH9iV1acs
d48DHQJ30OdhxBbHxFgr+hpgpnNNNsT+kHl9lcYVVLZwY0rfP7Rg3C/ftLnNLYiK
nW/siiTC4iNdE8l3+5X87lRImp3NlcadCbv0NBOtNk1LJQnGoSxfFgFziDsIzBiu
7lEh0rd/iiBM2CGgCQqLluyg1lMNwD1JMJ3GWUXrbXiF5Q4PjKKWTuuTOooGpW13
PPy9dEU1SWi6SFQ4GtcEDA79IgCwji+Dwxbiq2TvNoPMqfM+nY6Txyb4uA1hEkIu
TbDVJJc6YNu2TgaL+hxX4YYE+nzCqZqB/Xm9iuLYM6d0BZLfIlgsiBC7tUVfQrQA
aIEmfRiEqriPtSUfpzp2+rrZMxybsCEVoaFrtGq8+4NeQyFS9yMSANnoV8YimIeo
7AeyBp8qG490eH1WyEUczEAnynj6cf/dplMV6y3ZlUTJaIs0ZLRiwDmboTTahbrm
zT+7ovSjIqrYCt7eW9WHs/bpyiBP4uk07jfvBMMFQtvy72gtxKwGMPRWu4uvGUpp
8RaYwBvWl5Nb92Na6freQbfLDC0vi3mniI0fn2OIprQG6bU2V0kVVNupJNoh35Jg
zwoRjE4hMqQQkzXSF75Brj749frGjPIE0Op+FUfQaZE9n1UcVmujbT2JCe6+Rpsn
zQ/Gl2RGC8cDVIH4z+fPJhRSom0g87TdVVS716I8KzyVdDl/lhcyjV64oz17eHfn
wZNJ5amNnJBJHY+sPxXBTPzZ/KlzGyyHae3Q9zUHXvCt2X0Mj/7lt+OsFefIhq18
AHUZfW66IAAO8swSoG2lQKZSaUTusHwZtSQ+M7yf85GN2apMFv4oEjDgDrN4mK87
H70iPxa3MrmOtrUpz5oNEqenN0iUxmDEj5fT9U+cMh61wLdGUPWhu8/k20a7eOjP
r2Sra8sAAfRfxsYlb0X7dY5LWT4AXerJfg5uDWi31JKzTVpR16KpIqZfstInIgmh
rbBisouoj4jTYrrocapycR4iwewX39hmmMMzMJCTd/bcPMFwpnYxZ40eWtJFU32E
acYiUqI+8rdj5llw+QFxshQSagFIKeuvbCYGb+AbqNa9Sgo35YgmRUH5ccRwJZ6c
OFSXJS+xEWj1WSm///rs9/tSIdxTKw5iBWlBV3MumZSwI1houyVTye6IxgLzBh35
p1ydqh35G6cQdxL1ZzB4jyeEaZFymx2Sp5XKAQrNx6hEXDtSDUYT1bNdw7quA4wD
mItKVRsKOH9HvsWBvN26KQKhMwovMERlfgghOM7LCqasyVLFEUdVDzec6AxrTVMq
yLqzWVdXNIKCmip1sOiKMxGtx1gsoMbShMtTgII83d5ugy/HgYS271PFf1GKqDAa
Bc95+MA/ruStowupN4876L/b/wK4+bLGwJZ5PobmsEiD8/KmSOR+nBPXSrp4iuuN
Veil7IqhscuhU+/PJOdFlSDSdRM46xkGL5XkXmlNaAiX8UmFvZKV6OA1NxpJ2EhP
7MyZ9TQtaw4J9fGFkutpiloTZTwyjKr8s0fiCZvmpsGYau6RGkF+r2kV8+diQpNb
Z4Kg9cHOcRuiYcmyn1Tkl8g7TfPXSsi7gx5Z8R6uiDR3hopBNeCFELamyZ+nwxlb
mc448aNdj0u5EaThx3Gtc330VBxO2cHTvX1bQpHehcNQnH7Rem1xKM5NRmUZqO0o
1i/ngQwPB3Ipvh4fqxkjJP3OFNRieY3NYFmf/AIS4oAF3l+qKHs4I5EkPQk0XWxy
xSJQLqL1gYqIF0SilFPdTuVy9aXVQVxG1yx9x9mUlVOB0Crq/GVl9F0Ro/K6Y3UH
lVrm/taprpRiX/vwrfKtx2FWkDlI9uD3SIi4H9NlAfz+b4P574/usT7I0nspgY+x
p5AFDK15M85T/tKXlGAktMRmsJ7PSZBCjgfhLDrQCxJvQ6WofPJx2b/z2GhadgFP
tCFM1oyCHwReGXoFC2UM0EFuyYeLBIrC6mYltbZrswXkU3e2viEfvlC5cZwTU0Qc
J1nRJBzFMigqnt6cuaqUTI4tF4cb4xFYbPckO3NjAkf8lCk0nWQeFZWHeIvBCj5Q
9sGSaZe4COTo7zTIF6S96rPDpp1jRfbjhJvvoQxABBUYFymxEYNJgw6ljMDKyqVc
au9Bftz9EIcKNacYhfYlitch4I0CrhCKkM9ndONqzaDIqEIxy4eydPEww3vlSyVO
NesE4KcbfqpgrYTzTs+TieOwNjGmhYXEk81cKKn0xeJRR6ijrrGpVZbMElzPQKSo
gqV/bcccF/QS8brioax4nmyqbOvlHxdJCZU8ZfEStH6liG0bKzK+9XErQ7fY7CFD
dxuOv1x34DomhsYSop7dK94bspT2DQEIXI/fTvsfkxJQTvBaBl/fitokCUn0HuFr
OF/QeadohDXXD9VSPo9GRrlWafAiolg7Ks3DDSJMFq1MMMg4b079CL0T5SfJlTcs
Wy0w2bYF92YXigNL/CivYRor2pvftMB7O3EaUuU1dEI8mpoYN7A7oICp7s0XbNcU
bp9/QhtYU6SsGsXVfyQycoiLvN2v42NCQP4Cp3v31wFW38g5qC1Nc30yopt0VPQ7
H3t/YA4OpGCaQYbSs1NXH6cjjR37ihblm9tRlskxb1ZhAa02eWZZOVK9kgDXh+iL
zHE/0+ibzeKXeVJtLk7END38JqtfM6CO6w+xgCQI3c4yeTXU0QYPg3bR0eYVBBsN
LGxuJt1X7wupmEFbjypOQNcugMM5okXAgz5LE7BPbKE4crtfkzuHYMHb/lqcF3CB
ns3rYdB3XrOZfeGe4JNosYu1e0JjleWXlUlMwpFzrx08lOrupof+Fnjz5DQdkX9I
M2rI+hJsh3DS45bvZ6t5rnzf3uWHWooR4woxKEapLziOxtQTduUf9xZ7ZYYn2UCw
3iGU4yz0duEYKyAUvgnR/I1TPV5pflHO5sVhXUSRrdWDgmWpWt/HviyeBKPiQA97
zyqkxzkalOCcsRb0VsLt0rGNIG5FxNpPx4nf7ptWgDiCXY3T1BpMFIizzme9KnUk
Hpzc8dUnSVmUSdTHNab6oqi+lv7x7I/RTzLpZVvRSuR7eOY3aryZJn+svlDXoKC7
csVuJf38Sfpe0kQiLpCHx2of7K7FeNXZy2ElO5nXv8iApMMwu+irTt2Dnx2h/bP/
DPCm8zIBbotsbhOVzS1uaB4KrQMXCzRwbYQIzW9xhAFTpogj+eck0OEtqRccJht1
10Q76dgnAE3JLaRGR1an5AuldGz/ZhiPiO72+snoDYZlY1zv4tt5kqSgOfoEjXCR
a4e9Y1Hxa5cFKk1JaKeDC9TgfuqxndOKXKJhuUxtR4srA+krZU3Mh7+kH7fW9OKP
QltALaIlS7QYi1ni/eKSYvq+W6CqowTEliIBIMTseOsku2uQvEqglqUUamwpODNa
3u4LHb3H/k04+X7UuU1A0IziPtMbPD+lpG/i6GRiKTO/esiJqtLGrgeP4agHsWbd
eGwrqYhP8BueRNqwu7XB2AwtCTZomdOroV1IVYX6Jt7rAr5Rm5mA66L05uEC99Vh
GvH71X9xQtv6OeMK7Qqy/9mlUjrm0nF+ZPSdozgLN7jkBhHA1LxTFBbZfAf5yUXF
dgwGRe8CC3ANgrEJtsVCyjah9ucQoRjtv6UmpbBIe2ftmHflKfG3quaMIRWYsHPI
GQl6GFBg1TW31GEUByFQXo1U0Weo9vb4+bbcYlxB85Up1ubCAcbq+alyBIo8utYo
TazR3GXSoTUz61Fnt2rohQzpgBScxLIuDPeYkZvdLvhSwVXd4rI/wpsrtJQpbu44
UDo4ENcaedO8FMDeEWTL6ot6wHL1+O9aLGWzGFbNSbnFiGBK8uqvqMp6ucwauEnP
ZC6UX6IUxso9o/4d6rW+t7A71QcCqna83wtwVsmWCxuOFGF32UB3O0/DQ4AoXNgB
5+P02x2zFeAI+4xvzQJQJvMWf6l1qcixtf+Ln5awPRHOZsVjxpcdv7/ZPVfTwvU4
vtFQmEA9IhsNQiwKzwHaJMKVdBRPXotBjJy3Z8Giu9MdLPva6+8yeZoQysDmhuts
Xf8chCl4quoE8TOdssh0ia3l0QjXNVdgYSDUAaLWyqY3cfaW7PQjUYH3HNlHuCGF
hEhbajn9MfHzfm/hRAodyQCDJVLtnlamqlnyFbnSoAVTa3BM/nsc8PwnK+cWY/Oi
OFiiiV3AX76Y+16AZLZClOmbn/OG0axGPVJB+SF8LLzsSvqbyHbwMkRy1J2Sz3nX
mJA8PM9BndjWIZV6o8zeYVEb+HzqLVFTrmIY3EdVe2fWODBlvDNNP4a985Ww7z/W
NvJo9vgFqrmYJzug9K7VE2aVdCXu017iWahBmC+Ib21J/J70XEgFurZM6IEu+EzR
LBT/dwSZZgnq9v3xuq+XFOfZYIxT1fKV761SvgNEoQBwyEJSioT6JehhrcPCabdj
aP2kXV68bK2Dh/oT4bKkME/8q6s7vC9d7k3uPwIkqzzmq1e4lp3/71Xv5IBfUdmx
Fz7ZE/LTU1b5VbOv7aiP+D5TaEhSTI9n3/qdlD3SqjysEwgIsldOr7gHdMpDF6iC
GV64u9Fc8ZjVxF+Sp3tYIECp7hhkRE2QtzJ3Sy6d4v7Cnv4zo2oJshW8ARa904gS
+Ko12aFQJn+PDVrDOkW0gyuR7dOIMq/MBhXFKy93ongHNkSn+5QCmVn7zMt06tUt
d81lH77m1PIT4IocX4pEbPbD4DoaK/6es5AlEjbnU0ZW01U57nyTuG2jRV9HiZ59
zw4hD5YdMX6wv+hsHM9Ewo4Xrtoji4Wq0kfWD83E0vQOipvxSdrtDCvKP7pTzNqz
mFtAoSFIpu1vQQlQLS7aEvM4wA824xruY2AQx1yLbbHvLH7LQibgHuIG0ZZtqBt3
U/GgQ3UIxwhOo0pXKFF06thHX8+RECxeH17ixZsqp4dgikujBmU4/70MnCKaMXFN
0XqpVEaevgMcDm7s20P9XixyDtyLW9k5DqJv8z8Qr6Od6aHAt/pwUPoxyavglMah
HVHH6HvPVpLfoh9wlH30ugyYZHkD3C4wIBURZHD8w5PapINI1KLj6PHT/j0UySYV
UV/GDfamKQq25ZS42oxbVfJnn6givxji0/vcM/7xNVOhiurkraMBS1BwXL30J7PW
84FbeWvmCbJdVhJz5qrMEJLqYUaU4TOpggfJ92M2Ca8enbdhcQXwAn70uslnJ2Sl
QKpADmWwKmUsVzk3GZwTvLhAExEPiCNvvwxuw+Bbd0sCioEXh51iHIrdtSzH8oWE
vCbwouGR/UgD7Ez3VpfVh1PuH+vNsMXoR6ltkAwrqqT826Sbd6oJOHK1wlKfNktl
BMgm3oOK02bB++aGoF1djq/t4zUfjMpgrNwxwIL3iMOZLA4UadExCchJ6PGwGq6n
qmejZceHZIbY38dpBmznwV18lArV/5gOL1KNenUDWhWss9OcWF4yEAkYCprT5cE7
M9DoIKmYX62iMwuxMSVfkk76gcdTo29sDvZlgtm3ah8dtySzaRXvdk9vOV8EYwBV
5OKfFafejTfDXJiRiT09bXLalL2H3PaPmT7RPTFHcR0j+dSYpeuRpbPZNxf9M/2M
/0u/D0I83knLrzVdRGF0HnWGaDtYTJcAVU3aq2MltafVJe9venc60c21u2sdD6QY
LuQd5Hk9Q5NU2TnU7oHXkj7cbmIV5ZVYBu6VMQRn2YXJsbfoDTGXhhU4a5CUNBDB
m+HE0XCubblTLFNmaR5iPRDPl1itINxYLsFCdciMmACL9z8r+CBq4LBi+vWKI0+W
QMeVWNl2xuMbJ68OzvYrzjt2I9SeONtJhdzgn5LhBVgtJHMXBQTZfPxLrKtpVLiP
dWMJtayvmvUAbCbty/8uC/ZKoyY2S/wMjqUqh91Y4AytD824xgdRZKuTXNd0t3I5
izmySzJbfVMoBHTgM+qDzbTeQ5LHF+gPpN+zLPrq+Di35j9eD+eQtJKubiH1tIjJ
Ty4nPatiHVIlX3hmOueg1TFx0AhD6eoSLcibwEt7kEombbUGZFUqrQfwHHfCX8QO
EmbmIRD2vMIfqQd/RjEPr8Rw5zAML0Eh/52tpER8/ZyF1DP7KYUc1agnXH2HzcUo
Fk9OmYihHTzUvmOqevpyNI1FbFh2f15EuB0UG3dTF2J5eSIfOh/xb3fYnzXHxIKZ
PkTJ4d/XV6tHu1cTTfUEpx232QKyK48mM4klgGZDfVrelZiqonyeDXUhCtQU4J9O
HxUbIiWPir3XeLomksM1FmYi1iAJR5fzPVQne/qOYbOqeclIG5gu+5YJGgqE2+oY
vLfm9SknMhI2Iio1GOBasT/kRsGdEZfV4qaNY/8mXuICk8B3+IOwoNEFhG6lyZdU
lYA142mdO1SQfqZg+9y3qGdGEcHOHGvub//RNKif1yHRXEOD6pCCj26y11vanhDN
NHrMcgoJj2jw2Xu9UJMY79yNIHhIkyHhCdb8gldPhYLS1UlZV63f37yWlNEHFJkh
sGKb2xClR40AzdLJavk1cRvphj+bRqu08XCBFYP/5Ss2fc32Qu1l/kCnldjou7ei
NM8y1CJvCINcgPUg1UaJqRmUu71YwHg7OxdXvU2X0OAYFFdhVkgrteJURAJBi0c0
qj4muciuF/+8/iCb0OAM0r2o9sKTj9Sco8+uXjNS3fmTRDqhOZDUBkdyYw9q0wBe
db2aeR0Gs0pyb7BHgZ3Y7MRM/AufJryTn1moCdb+KYLAtCIoCf7f2Q6nhOHsY+Jn
VUlenaWChvhvUd7K7bBEmYxU1VoHwixzhQ+U5J10d5gJOjBHsGWfX2qXrfkSVlWD
gwFq3DGIrptW7oDCCUMWvTcq+5xdHO7bjFt3dSNJ9uN0rMcgC0gM5aQeKuzL7g3H
QkfZ+IezQ1j4Wt19/9mVMEu5pOMSGmHfjY7SNDUsVQxT367s+MMFmhZmwQbEYLhV
rNVvD0WCYrYeUBkMDY5K3Qo1DGV8g7a/7GumooKPg97RdBmk0oMUdKTP2m+eHuZZ
nVcIVYIwegZ/flV3D/O+0q1Cx5BcGJHxKVZPPVcWvYiGfCAcaO0QnglHcziiSsVU
TfgNqqPL8e/E53w7qa6Joi4lFIMva6Qb2fObiTDs0j8bcY0N2GAnIu83I2Gvtg+2
FjLwk4YPbuGvU4zuHxeBSEO/3+G1fHQpzyftm/jDhnn4wFr6D25IOT1XAsNvfSCr
kJwSd7p3UshfswDiSl8l61pI2nWoc6X/S9FyuwqyrdTzBHOXUNmW308ico4ACzEt
h6juiFzkXR7vk7aE+1/IigkMPNIpLlNnXCYu5gP1E3dzXgFAwjzchcQbg3OBDrON
ZaOEUMSjufVD8wPC6mdWNRAMbeJSP9CrjAOijoE/FsiSBKrHBrll9GJV6EueSBB6
y5uNa/wiztF45Kjk7KPdSEj5UQM4ie6ydwZJqPtlBg5hZZitgeNQpl+eiBOw3m+n
1AEDVJ+mTZwYgZ6H/TEAPYAN8seGAZ1ybUaOPTvGY/VorYmWFMiWWRXH5VvqoQU+
yyHfQBDqbtIBQTUGTGwLxudICVEfGtDZTZ6fCOoFiwJFHlsH1abcfikEylyhGDv+
o49eF0Eum3t9blADzzhr3LNxoavj8rl8bhFHMne6iyZgKR5wjRSA5k3OCpeO50Ua
3PpaVTe5rPFFaxZ9N3gVeEc+ewM/jUq4viqikZdwbkTr918SEETSHjECAXOiHPn6
aSuZBfmqF6QbgL0NPKxGGftd78jY/URDqba7gC1qxfXwIkkAUvDTe4Zsc9CcRLUL
PHm206quPPCFCOEi4wEJ979k/Bi1EaW/1Nw93zwuEDoC137IwSiYSC3TDGDnH9ea
LcHNFWymy+xrSMssIjjgnocZPM1O9v+wPQc21NtOW3YFsLIXYi9lyRxYGQn4zsN2
9p2XdRKa+zjEf9kAUnGzDCGAh6CIQME2yvHekfklOnYMt+I4dgKP3ZD4CreP8K3K
iQWxw2NC8Y55LxvRq+DRnIDN9As9256R5twiAZiuJfQ/jhkCxEfHGsEFYHQ9P4ek
qNrxZx8+6Pg6w2i/8zVdh6+vg3Wc4qtoYzwF35bCltZg3DgUpAcTxJyk8JIyZZz6
9FDLLgGQ2UCW8pwM5a4t+fJr0dIYLW8T6F8dyf4GBYR/zn4uhVrzQdAhByCQWc3Y
96PLhOWQ0h2821CwVHoyIpDw1IdDghgYRh+CBN//fhUa8SAyDbL2KsNpYXZJpVzF
S15smo+EbCvepXrxa45S+e0xuJED96G1E4+w5op+ExuJ30zRsVglu1NlerW6GYxb
omWpNExs84SGnLnTGaeZQoOIjlsOC5qB4Ngwqs0Es4IGKhWpAsnplx5mA9cT52uH
ETuT15N3jus73KTF81kM304e4Xtb+MtwTB0enNuugkyWI7Bl1lbQYh7Cs2a/U4pl
bQsWwDpwGrEXdmV72Vsdo9r+C+mqnJacQL+QNn5zIA/d08D5JtMovYX4pqdFVQ8F
D3vdQmnOmDUVJzqaOokMsg0HC1Rp0r7oGhvzyq3V1mbrVJYmhJfSuy1MWX8vx7Ii
eJ2mrx1KHoQ+AqfUDSy14k261wapJQWuVo7x432SKnaNHzJ1ph55FjK5AD4I7O7X
0/rZl5U/x/YDEvHV9s+PEy3vJeAmq4Qz2P3RsanTc+7HmkT407QC60fVVaA2+TFA
LrFajKjmgLgIHA7BE6pfMZjQAlkmoL9Hyo3U4/jAWZ2eo3x69rdzn/IUQQVXrXk6
j+q9H4ucOoVAdKu27lLRyuJUnUDJypr4oaBmMaYFD2rp6sROf/GW7Wu3I7LNw5NF
nmDPfHinxHPf+o3JL4zKJJo6V3VdXy3f9gVoAz9FA8NOqZzIPIv6QHjL5b9vNkIN
mK0KqrfxXs9gmnG5fP5Tcr7ty9Vmeq5i56XzNTHRjCRHwiPNwFNj2ov2WQ0nu+6r
vhVdqnEfUUPLP73CeSI2v4Y8Dnj2ZP36xmaPK5ktZ/rtufiNo9ZyE2Tyio6AfCR6
+JwAXHF+FR3EBKYlraDQRhyuxM8ZcG3cVrIHpH6YU1ia8tBzJmFIFCB0pAenpD2U
sc75mJogefweO+Z4na6t6mxcFL5O25VIBfkUNYXAtpJSOQxM47S01HM1/Rnm7v0u
q3Zfkftyk+xiidlYQ1p8ZEqmqJU4Rz3z+rnA6tjx8fATSknb1fxOIYRvlQr4/6No
jiA0hy8IBoTbfoY76R+6tUu3qrP2YCU0VI09bY15CgVZbgokdg/lUUnxC38smIvm
qCd35FZsIjKX8rbMjQDEvfux8PZGjY6yTbq9wjUZfnVv3Gz9t0imXWEGsaIuh6/9
tJG4I8LcbOP3XJjX4MPOYcAskfjR3KQxCjXhnrtmVPkh39lLo51/qgqMfPpEGCV2
MyaEFgQeOAutYu2hAAUsDQNpclXBZl3hXAFXtM4Q5PxD7kGk9DtQsUMB6umBDhYB
YdcB1ObZA7We70Q9tFeBqmBWTdvHiC9e6BISdsEveTbl/a9gfZ2cVNOgWHmZNLk5
KiKgELU3P4LGneYd3Pk6h6b3+pdi1qsOEGkRMUGxi1GZ5X3xcIO+Q6o7dnHMAR5O
FpzeOHwi/5yE20ND7vPJeMd5ELZcqfooCGeRQUtI8kicoEyCPfQvpPxoFpq6HdTv
KNv//+khkFQVnlLfTH49Xav95JCXyV2aKKYgFKTkkv06oMNHTRC1xVCXaOjoINuG
eNvOXMCZjPhrpEai17vZZtYasLPv+IIyVXyB1hOvihCOJiFTyzdSwrP0xm5gweaS
msal/zmVbMPruQz9g2Emfutykstcr5Ys3SBrOlJ/aaVDdJwxU/cFq4RIot4lr/au
bThZ+26v4RzA+eREHLtv+5GWAdywTcSEFs9uJunbtrEbbLatS03ik421eEPUgyEi
WAR5u8RXplBgbJZasxf3Kzy+otGhjHwoY9inIcDwipQUqkRBZBaZdSzoUDHR5pgf
isASjkmkz0rbMVuREOjCcSRLCLARPyizhI+DU7Bx8G7swcyjTwa2LnxSBTAQCN+W
sR06yE0uq7Jtc32e2ebo8Bgn1D++fpnw4d9OQwzeONdj4JcgnSn99jes5a8xmVOJ
YEn5O0CuTajYKItGSlzhJFUu1aYCNLeepMY4Ez09gRsWoyFsu/YR8l0h9ojzfnSw
rxBt846cX0CIPPI+QYgwcM9VPWJ65WCTwkdChJSaJXQz/Apkx7UZ2m3FDSkjsKNt
JSieShzfNVsj4FdJpnO7/I1V/zbjQhW3L8/AjGZqwwZjlDdY8Cl95zQQ02jjilcc
+Lr16i12vLKg/zB11dv7TRpIs3nozsRqpkDsb3s+oNbXvH5lRktY7rGWsn9PpFSe
ksUgfgC6p7i3BYS/icBtJhgT3rN8wmkZ9iiUuQkrtVmJpK6LSwDgmIoKtjQtVaNF
4zvcaJkLGphDHF+Qwp8m9mFzdrqDDL+xA5m4dX1dOiVCp8xsRXSxjdc6fiRkAeKr
w9B9Pk38Ze24F2hUXCut0oV1eSOpLeO+nKXL0P6+/+LCO6oIAVwdGkjNeyG5beT2
jApid/ZOISkL/Vq8X4UUhpN97XeG/Qnd/Z+Gnlr6I5Oc+lA4izMT+pfWXzXc4Lo8
QLTuRfcyo6CEVN7iM7xFWzUwy1WVu9X9Wl3yQKgUa6ErAoSYtlFAe404+GCOSf1t
7SecGH86kwqrCcMXMGU2n1XZU2Qqc/tt7PxDUv3Qc0cLR4K0FdDNzHuIA0Z/GeK4
fgdDHRidj+4w2TlrxUMDAAZuXkQr9sllm4BMsvFZVFauCYH5NdiDunB+Hid/UqQN
zwZvHqUmUVTBc4+xfheNPAHt8jyvmqAFai6mDa5Nxf1KpuxBxh2PFegDRx7L4yB0
QtA2w10i8CZ3CuH5MyeVeo7FW1bck1WRPpP53wZERWwf8NKsGzRMdhjWdptUvnoX
V8VMcWnyS9XTuche2fWGzguy5aCzN9RTPi4LrBlBzO510HmnUuz7DKBKYDig6qiG
2lcUU2C99lfVAdA45YT4rZgfYr+Lsk7iDZM3R7ZPDYAWGDaSE7GxZqrz+bkXBNGq
9/ZNZnOb+LUtwZD6k+G3fM9w+6PSL8sgg+N7g5C5HgEN80spyv2ljscg/wHluurp
SZFQUAbTjkNysTf3YD/i0K/3x3c2cahLu7z6uzlsTbe16b0NrIALvLnYlOe/1U1z
i3mNOwuWRoily0aEFR4zgIXZ41YwfIvneLQ9ntD9qSCQ37BMWKbOHbhL7h/M4U2T
dfEdp/Qs5nsmkqHkajFTVHYhSUR23APODSJQovP3eNdOqZGg66/hGIcjmVmrQRSE
KN1a00jUcmV+MOtfm0N+ORt1Tt9zItlrv+/6riAAi3D0iZbyZFTogqNsjbJFXt/r
ZRafye+KZ6sasNyBI3I1HiXwPslZU/zVDYOMUcsY22KoRMMDo018kfwODbO1M31c
rCuKSLnMby5vrIQz6cSgv5rjtbUXtIL+LWGF3fRYqWgkVYJzqq9YffGnoC+z1Ab4
8lsAzwFX/ugy3nK7cZlqn49IlYW/IiLDqLax4w4ahrm6uetJ+mBJP5mGYZSrC4d7
H9kxUnhSiFC7pdPIiujTZmyFJTQ3yWv3yf6hlyJQMjrHTt9foxikHdbFXXiaIwac
jzR96td2oVfJBX2rZkwiF6ijVD2fZdkrkA6qTkVQVaS4JdMVPTJ0MuxU7ArVun18
+b5FqoKmzxzR5YZsPFaoue58267+nBjQemp7rVfHRviwCUCD1DML+8vHJ1nVM1X/
s1ENd50XEqN+7LqMIXcvmN6g3rajVYg6JL0VsUlZN3FfU4KUxBqM5SxlVMXwaxhx
2vk69CPqpUd3O+i1587m5m4eFmYQM3gMOLZ4VkpNv+Y+ToBVTohLXk0o1Z3xlEU8
cUXKp3+rCPXpVxrUnLCJexyt81ndIY7S0CQX++0zXWeuY8Z6tR8Fo7JoNJxx+7GW
lKW+1yGoEjgOw7qtn36UzX+VSGg0B19SLOGof+cRWhxlY5e7/uwTsdXjkXo388EM
T5y3gAy9J7gDocomX3pXF5U3/cdVRSvS7tIresAurl+WDPTphDjzQXygvlLowXtj
2vu9oZ4DrvZ7I0lVFA9+PT2k6T02HPe9I/S1VhYuTXxNOztHkbhcqTyc8qcbvfLN
H4DK4t34i/VFV3hJuKkk+rEtwir9qwO//To3DnjkFGpr+k8LDbLotmBMTBzLCxUp
uoaDTmYz7w4HaTF5ka7a54WrRjkmFCWPhrUiWylQzMicnAPs9VDIUOIJTXyTHB6y
yMy1j0osVAGRR/wmusqN9b3g8+EpBPbNQoYFqbs5WxAutwkxNQuf7wjHPZKsXTqb
Key7/rMw1LbBrA158nDNT4eJUrx60I8xUcRe2MWAhV7ZOAbb6ZYjJ9z0usUpqQfM
CspULZxpzIkoAR2WVOcIViQAxgPunzDo5TVdjcobpIIlAe2QXs61Wy4n+F/5x39S
OOIeh0iTzJ12znsfYM1pP++f1QyOyh1JRRoFFWF/eopI9MB7i8THzYxi0ja40Kd4
j+qr1gSxPoXbnb3K8RPO3/7bpqf7EGueteyYnh/o6e4S0xb4HbDkDRrbu8UZxKa3
DJG58LVpbnGWN/av+6zorW1ql2R0RGG8k45Uj72HpWPmcUCJs6yh12IP+0n6uHDS
ol9ovfHij0J7vFf0610EMFgX5WBXK6t+6JqVHoBoyqESwn+Jt9vM7oxVONDLkDqe
hYNTn9jpWWBHpJWAZ/JRaM1pHKuFZ/aU0M71epiAEfNVq5pJb1leuoE0cYtyoPU8
6f9kkYcK2rgY6kN9aW/Lmm9XiRALmij0whFRemSTuxJNo6sIhJF2oZ3uqjGY2ap9
PUJmfJQ3Vzqt1OhBTKcLxptdhF3jPi3Bc6bSxqvCxQKyojQvQYeNdQhh/6ilGD1o
3kS44/Eu5NQQqN6zClbMUJHhBwy0IsV8C+fU2Q7UrMytFRtzwxZLeFyfuVfNhFmD
ZmXmdsENE4S0EfYDNUA0RTh0EXxcQsWIHUBj+tHoNoZjQywnzg9wgNUV+TkQLJT5
BdV/mRKQOJXIhilZ+WOzzNEMc1WOUJAbMnb6MHpE/3wXE4CQgB6yH/1sLbzPXsp9
cdbiR6jkN3u86QwOQGet6R6yoTqphppDN2+lvPBvxG2+louWaaG6kz2JbiQZXhZU
zcYZaHFkRX+bTR8nS+cIVQwxCfte5VFDfFN5Jz8C3vqOyjjA35NqTb3fnx1l6K+c
ibc+nZQiByKyVXplEga6dd+RtgQuDQLR5mpSDZVp9sz56NrYNf4RsLXbEIjrnm09
4U0PzX2geIKsGR1+D3YtXI0F+xNy7B9YoDTENj4HB9opVRIbfvrntq424sQ6biBn
Jl4LjPu/diNAJgjBIjHbtto/pdjavpKodzlne5qHrqdtplda13ld33gWgF6mD3xR
KZBSk8w9c5ordoOEX+VlFbFqHctpFrcJaqaFs7U8oMgEDW5mLViPVkX+aRetODsm
nLTgyOgvKqct4qc2gc8iQIHmfTiNG5ckmIirAEg2TW22UKioTS8ccMKV54zDAeBQ
BpyjevCEkVars8PBH2kkOVCvfyBY/FFGfOU6JfnpAT31pGv/gOrvOoD3R8soA/Pp
Z+jWO3O+ww+6xdRiarm6VV3o3jIxNcobT5sbF7yj6TeVpWCZnq1MnwttLqvt/i9a
Jr8wnVtPRfkUDVM1DYcnLR9i3QXKv2tcjUrbsZZDhNW7XzVMwLX4vMxpvN7plxCn
Amg2YtIIZCYZ42RIoM3COFMmgBpuMEGm/hM3wWdM3twQcarPDm1gzInxHUuo4iJf
xBlSpPK7/d3A6p0T09QHk+GN00lZcs4/CpLXF0usz6snQ187ddyAsiJKH1pAISVm
h9D3vQ5wa2CfQgGBAZWa6gP0Gn4ro6fTVMPLLJxkGGlTzGPeZc6m80wvrV4gzQTn
eytqkkvuuA1LkrucrWUHzq5fsvp6oLnp2lPZ1l+n6seeeYj9v9cZAXPuU5uq5nYk
XB9CdTth0klnvIL8on8eEM147+k1a79Pea2nnV5Bd1RVIrSTSbhpGMbld8KwFK+j
J89bk0X+s1pS2gwrcFf3MqUoKwTFBasxOvdxBlVmmmQRgPYwnhQb3WU4HzaPAVSw
c00ZqV1Qkv57t/4OueFmWci9OirzvbtSuAJXJ2wAjZ5SVgtW467VJJp5H9pstbGs
PhaTpTr2RcAubz4lwffozi3L/+DhL9nLCB2qeGRLR8wTfIYuf84mbl7/CpnrymFj
JcNPBrF20ZCx+WJ8CI9S5E64Wk0REXvgLQl4zIaiw8ynefh3lBmu7cwyZkkWkBoK
OFBVvj8rtdY+/w4A5E6QGMAUme8jr06yUbWuhKfDlV1q/90+h/70rpSSlcnP9NXh
DipTWTbcHVfm/Se47gHxLDjG4CnbD//k8Hs1j6b57lrRA3SJZTS3ViRgHGk1BzMe
OsA3AYGVB4BT2T125tyjO06llLb82JEVzClKj/I+8byZ8ry4+6bv34jQyXE1FPaE
pyNg3SAuT664G43qH1bnWkp8tAbOscz390fy7ZWOALvxlVmaeznGEzWOxmtLgK1p
Gi62WZ+9cGzi35LgqHoNmqm+DkWFBIQOnnkh0v82/GXjwwbLo9dSyAd0gcM2ciO3
cpGOTMg2d8VfsSaRJe5O3ee/QJXJm3FZx889xL9YOuhGe8ysDhkyh9BDPaHvawVT
qlp/quZ04Uw3X6FWa8dtBRFw6REXMKPwcZozNxcSQRIym47092xx1jllfAlvCuPO
mbSzI6QW6UYG2fyX506S5ozncsb8Bsh73XskpW77zEekwaVH+xyHq3RTktkObY3O
T+BiI5hCdjg1wFVtsKfoCf6Fy1IIs7Xda7g5qXfTum9hlmM2v774WprKCUu/2V48
GO9spJNyjp42PFmN9IdwTJYd7LRpgJmnmuxsODWopcpyTdz1lv708XEuINlI1q/U
JJPDURUUu1JAbrw2gSIJ52yPK4bsLM3j8rUg2FtqpXYtSmsADinKlNJPMbNQ4Ajz
iYD5xrc2eq3UooVeVYh3jlwmvCnZdMk8ygdxvLK0l+xhcOL8C6MRb+H40b/rA7bc
4r/l2KVf0HYD8pvqG9lE4zNrur4keZDVULEVhdHSM6GZRxdsI0XVuGsI3u7ULxnN
ewpI6xYM2maHC0+knEcZFfC5A4z52/njAsog++mM3xt1XXs01hxm2g6ZsCmyc/YN
/r6iRaurPkAPGmO1i8SfYPYgCrYN4Diiw27SPLmzBq1G6w3qeFkrce/+ovUgDzJ7
50omhyVx4GAsHhCbwXuRAwGefYsROzWA/FUgmU0jpBre0BOBz2nFdjz2rPTwRT0B
sVb3ssKRQUCgVLh3a1hUGmxMY/4v87wDkKbA6c4anqYPLUj5SHaep/A5HRkdObBi
9HYr3RVu77MDc9ki3JSljcnkYct/rsvPUBfWookR/tVb/WZecfqrXFWhN1ficZCL
HxxhPBRKxjekK6O0a9oLKdF2YBtKo42/yW5Y/X2IAKi7sdpi8vB7nvWbRxzolVbo
YKexklmKoe+W1BF3l6MIcpOJ9ChGM4v/xMTE4iUKgAWHoS6M5UAjLDSW5w4y73Aq
dO5EygKN7NNXlsIF7oXryczmx5LRWWmegor3DvywEcxNXaq67lL1cCsy40Yo+X7J
Mdh/g0Ltx1mJ65j7dtYd2y6x/mZogoR1ZZYGoFUV6oayNE6HxXQPSNbJT/G7kw2m
jwaxMvn9/lLvqHe8Qtn7lx6pQD7SETnN1b3NX1XlJuTqwtTIoBEi6zglQW6axfmn
wPvdfS1EKqnvjzgKg+cFoBwaJWdrkLML0pRLq7jxhiclnkLea1pRy1MlT+NqzUfD
XREmECJrEaj8VGxsCQzocSz/Bxv7z3DVTuVe4/JlWYW0tTonDrGlIW7FdBZO1+WE
N8EdS3IDNbgiyHZ5VFM3CxkVJIDmJrnc2vyq6aBKUh0SQXtDLCl22yXGyg582iNE
e8S+eYQrZQXxePnXh/wGaq4KVmBzpQktxAYQtnsFH5Q5SdfD3/16IcerppVnHlPn
GIv2f83XaqPK7hVtik/FShOBSgKJjXzdSecPeCl0iKHTPTpv7n9XoBaDZiP7DXlF
Zuqp5pTGHHt92YkykVyUlsdV8dJyJmKnIs590Gf3OdJpnMjry2FIvQS8fdsBsQXn
pitvVq/ULTrO0aboHZfSbXJiz02lwoDBklYj4HW77D5pqPWqouQhCQmEJ3cFeF5M
povd4UgKrBO/dHBbqHrj/SYgQd2yrxl+Z16w9gP2nZcI2agPdEG1tQVdH5g0Mk7Z
SydBVkItjsOb41cUurzc04+KyFMqnC3wnv9oDPodonq0I/UlAWjyFnXQVdgs1gJQ
n+BKQ7wLQ3XU8R3Vt/pyIlmRw4N8xFwmkwsLXYGT0K8oYFlHihMq+hbAgkhH4wfw
9h+2umCXOF+xLWAtOaFOyrIiEcL3GiUDFyl6bvFRuOGKCbf2F0sGDmWsOz3MXXhn
Fy2rXcKN0cdoSVfxi2p/L4B3dmYlxIwiLaV9jVOfikMprpjTpGcQniO+PscBfsmW
JxF0AHjva2tNTryCyr1uM7PxzKU/5fXZBqpn0JIkXiOCz1oA55MKQnVzonKaDrW+
4Lj5kzwkR32ynF1R0IeGFpQrhcOKV1fFHrAwfJoR/JqlbYRRPtAjfdwRy5clipQT
2rQ67C/nFIU1u4jixyUGn7QHsvwSFl6A+it2eOx4MaQ1CIuAVDYwwgD6A1tFMxZq
ob/7djiy6dpP/BEvkkhDoFFRQQg522XBXBWu82QYuCfZqJAImMMta5WQM2q2yI5p
AQdL2wQk6bSetH20zk2x+iFZoShAIROMx24xAW6Znt/S/DbHpgm5sM33CCg1hri9
152GpO571CMRaLDzhp3EiMHRwRTk/gL0Fn24mB+zGu7q50p04Ax/AANQc+r7wsHA
A/LUgCmfzNSS8e4m8aAmGOn+VYnI78bVfun6BnHePNO3Ho7Z9QW8XefBSPcD7SXt
5TFfsF4aFNe+RTBsREHuGIR/Ye0NZWKv6uYammcndoC4YY4i4u5hGeVbo+ZoLJO9
qQeaO3eplCWCV5xP3Wjk8xPpjEvdzlv4OaWuD2BHC1/9AjHrhde93ojDDyQTjA6S
AjsBrfaYbinWde/I8L0EbhMRAh8IQvO1Q19WrtDCVYw6kSx7mWCqbIL1ldKfkyXc
EdXk8Tc6VltIrA56e7DNuLfkZMe/wCAT9wWcMeOgTOfT1kOK8uMtQHWOvC6nESWM
a71dtNuS1avlyjp/mBL5GRRM9xRBJme0w1uM/xfYyxwzGqD5VvExbHMpGre5NT92
+C0dRl5TRZlHCgqi8hliFvGwCTrMPFHbC7r3/t2b1E5dD6tixQWcb5w9e0T3OZQn
NS5b4LrgJcfs8tJOCSS9blXe2Sm74/e6EaeneMwe/gM75f+3woq22jvLYd2Kjnda
s65WcphI6L8UuC2NeKqSlhcxmKOx8m0XkjqfB5O3vtTNzrL+SW+q+PnySmi6kP01
jiQHJVioBcw/aZGLiQJVCbsAo6/XtRHt2zKucEzg2S2Kcb8lM3y64YC1lp1h0p1+
bDcbCrP77T5SZo0z9h7LClfL4XomZTlarYXAzK1g0Z1wJzxxc7YZtRZ4YUDo2JUj
1/4apYDAZ4XQHcm1v5lkCydV8WallFkqPjNdv01DVCK1BXeBSVcbfSjowXCfmrVF
NBVtBESIAvOK4PgcsyhjK0zOm3JkplNNuDzyS+mqCNiJSUw7LdAy4RNK2XYpBDCh
qx5krRv2sDeJRiPMMNw+RJuYWZoM2xK2jq2tnQtKapWWMq6FG5sqstSOcCXDZZlB
BsUZJEYhzpMt6bBqNYnlDnzuoZlHDz42Zmj0OpNLF8hBFSzcoTx90f9HItzj9Rls
UoBdOxqh7zsgbBC3x/SyzO0Pjgi9KXqOOw7InncuY+ivGNlEkcqZpYWHC4JrRkWn
PJmCGmYUDQzfbnpHYgbAAmN8OyXmfCVWj+AmEHOMsT8lwOUIGw9/lTVmhRzOUaT+
STuc481bLWEy+zVO89LwpH5Czn9cVX6P4W9HVO5pqpHsVMX4DgkFIbGgUcGcnlmQ
mXVE1RdOsISdi3CfPr27hj7BTn19S0UMJVTAHCTCnm3bVH40R7doZqQByjZ8r5cD
r6frDs5oNrkxVGajQYV7m0TxkrCo2oKWEGntoXXnjf6igINU+2OBWIzcsg/q7Ywv
/KVmos/ETNXizQpE33iIGpVgbgYU+40oXBEcws8czR1rFk8CJkSAC7ktkMzaM3kw
JJnOjMtwlzgcWoDy8V16MBnY6VyzhGrETDT1ywjjZS2/Hg6Cxv3aupNUGp9JOdqc
RxNu85m7q6EqLQt0l6eELH2x7EfIDSD740TX+0RG5Bwp9NHYP7XpU8u8pZhnt8L0
fs65kSR1BdkAwuMfcoHtWAimzUqdLIZb8KAeIovBWi/NbZfvp8jhPRICPvRd8tfo
Ksd1r9jPwQlgN7isbzeeNyOowCVoEDOBZc7w81TFXCQ//QnjwA0TbPIjng6fCKNB
ix/pHUYc8J1vhkIB6/75aNnXgyt1972ZrpgNYfXknoak3zMRH90HdOa5rkHA1r/2
l4adLo56oiyUAIfAeiM9syN14955qt1PtNxwC4yaYLAz1RQUtFou0sN8PrPtX5+k
LkstoZF26dTzanKAFlCfP6H4YUCz7Z3ZGpi116ukNPFJCcilnHIZ2qv6a7Lo67b2
xL3bwaHd7mJR47MyxFi50E1IyWgSwx6Egk35WnaaNH71IHCq/sfZIqD6g/UNvO/Z
WQ0bBEaFo2Od9dj+18F364BkALu2+ivre73pBy5TKCYIwn4Bwndhy0pO0D9duzuN
MwJu0tlyU+92txBYqn+YgqozWgShWTIes6TR5xoDK7h6cPwKWO7KIo/rgc8K/nfD
J0g+k0nxGMmJFHgXXkfj3oDCgpPja7YeDoWI0JYVKUfaA6EFQqhAxjzGVq3J4Cru
eec3/YueWq0K8khZy3UhknHaicAC88JIcDDoBXujbxxls8XurgvdVISxsjj/fFTQ
IHRS/1OFTok44T/IpIHY66cn4ZqVx5qA09F5SLrtyWvUifXfqjUnWR2eRBKzoXyT
OQJG7BOk7Sek37iJrfKHPB6Y9sxlclniQNumwK/JvCuB9+FwgJxV/vy5QgYfgHke
Wv9e4u6HDhJAs9tgDCzuRU+eUBlh9bkP36BgzXGuclr029n40WH+aL/VAbV2JAVF
RBOgh2vydtGV6K5Wu4ZnAY4JlA4aaqxveJ2s0SnSZuz3iU149sSkQaVBNYN+l7Aj
4FO7udYWf5SpoHFRaV+j4i1ahga4HkcersxeAZP12715inYl4VxaIpbK1G2VKexG
MWmNpbr8Y+x863IQXpaQryOCx6frCfnlMhxYdtqCV9XsyOZ8u5GNa6YwIGBoIqh6
+ajhqeBCT8199tXnlcn/hiE+bt6sPNI21J+LQnm2pnf5lga/FDtPSYKuyTf4fRlV
oIXD4THNzPlxg2Op92FKV551nQrjBotZ8dFEWR59ONFuLc12hI6dT877sqdNxL52
eZ3veiUU7F2vQEDDHUXtQZBpib3SASY0Uh38M+vVhbtmNxgBBskRLX08jScwjniW
mmMszZOVnkGL213LNlvP6na88/xLh13le1gqqjD7TOAbPSRhn5q8aLjEX9m/wnnX
BA47YcuqQzdVNpU9MQ0ynWJGwcx10NiEfi4f3mOXGG0GoYd9ccrJUrZ1cW5u+BEL
6T4bp2+VdGV8/q02+vZcdVCAlNb0uD6jxTOHSoYGQXhuWE9vfNUTEeHTJujlLTS8
XmtrFOEXDAyKYGrQWbPwvCDcxVyCqLqUn/JmkyGZxJHJyZBlcdfT4SUsmDCs+ZvX
QeySv6WIPZiGbXqN/MVXEbCVISbhJYmre9CqXTbGlPImTUfsSI3Tb8dHmscU7MMb
yd4JfHto6wiNqfXJX+1VoxXq88m3TwBWSV+Nz9V8bE+G03h77E8N9YCuAsSbNkL4
kc3ApHs231U5g9X/frgSzTYpJKEOYQ/zdKdgVLRLgVQX1vZ6CS6IZx7NWt5zMRoj
j0oion7+SE16JvEI8YfAE8k61o9JjqZvO3rgmMCvwHe0Tsi5M2eopLWsrDD8P5hy
gzyz2vD728w8bODIDbcK8svuyAL602433mdS9FGmcBWQEVqJL8Wewo/ggMQIiFdE
QA2F5W5XmgylJngQpYhg6S+0l/qBS+ZJ3l1veXEhnEf/xfcr3Tf3FxTa9REJee2D
cJMg6uWyVsOCchPmViYXjZ8/Uu6tMKeF5n1RFUbXHGE9gYmg05Mi042EUNDrusrS
aGbrCgpR/dujDU6Jg3TBUbgQPzwkgoFWcjcBS9RqUNq+DpiEIKQgcWSAwWD8+egj
lf/VdFN94eg6yw2Yn33njTa8lCE/eWypwX7LofstR4kCvQVEvNMq8sT0zQRoRaCY
cAiBU1UYDGC30eO15SjZujQtNgv3LJcR8R0BHwh8jSspb/Ftd2AqaHsicQ2R8/T6
tLKaSMzYvV5GmUH4fCM5N2zguiZJ2IwDWl6jg6ppoZiiGI9dexsHR1Yg0/hntOTm
lp/2kDfk7QLogdPyVDigIpNDSUjG2p79QfDwNehHAoQxfgcpl0Zvn/fTmuRWBAxQ
FumuuXjKeY+kd45Epld09A9kQDtcD233Wxde5WGtwjSl4kINJzS9o5knbtww4p99
KffgWYjKKZgy5YvmG0NC0tExMbq2eSm8idkTAk1h/ByH8xgU83BRhek09aVfAFYQ
YEEg5u2u/oY7P+T9ffX/fFnGz1bHN2OUVFbSAaj+JMnmIa8URyjdLODy5RbvVwiD
DAp36QpEkoUg3MvLGeU13Hat5Um2QghF63eSCAoPsNDv80rzK/FfZ+3TDmlTNI7r
59idrMXvEJKXqS1ZbDRkOuB5blW3dnBY8HPx+t2yaBnypvYYPMjl7yxJlVypioGO
4/Qf1Yy2cHCleq4kA8pG1M4L/dm5d3AzLwFKTH5Mw1Zuhv+V0q5BmCYbdOSG/gGU
p1pQH4ZquRA5pi2c8bkyuLuCrwdetKTU6roiKYrS72JAkr1UCQKXitWuwP1nWxIz
B5vOLd+NeSsbkNsNDtM8hosFfiDYXK8s3a5KbDWELTTYw3iI350T67bGFKYbj0jP
DX5+lG7leLr426HzsHxrRWHcseeFWqdNkLE5sx4oZVIbwzXsESNXM5D4KFvs0FK0
srKAopjoZokxbDaUBW5Ua8oAW/RDYWjz4jW+7iNg6WiWtphdexTX9l7AjtcjxePn
EbuvqHuIHqWkhQ6cXF49sPr3+iMQ3BEmByZU0mCYlXdrQiBqFA8w4ER0DJpiTAEY
8GQAVGxhOwuHEPIxvf3fd1FIMs72I9bm0DO83VJgm87Tx1SBOnyhcwaPr4zACAs5
QqsUBP8+vqlmgPfM4F8UcMLD8OvTf0odiQT/zMaqQspvoV50goS/6hrQEBYiuLpp
QwCeH5jk2sZE0TY7bb3/zJW1U4YQP46uxmr/t3L2oulebchX5qDqHYi2UIzsbFo1
qxWDKW2O/cUZYAjjpdJCn/OvK8bAMQiqAN5ZF8fTQj0s+jQvlsXIu2tZvB4mNldv
EYA87hfmdCXcG7NQZ0wim04KSw01EXgnnZX/agxIbyp+PnRGdPTf4wgu8sJOC/1t
7+j6GeJnAQr0qifvsVvAH/FlPKEqZIIwAsDHJWES/93fd7MfQMrYJHigJQBTYNNH
McPHc9C8jI+gWfWsbc4fac+Lia5uOpcXXfgLxHu8XdEYmQwp2ncobYczp5dInQYP
odrHiXK72ksU7lEr1HhUzXnrHv9oXA68BiyOwwvmeXd3TnzWSZrdkXEibewmIeRR
knHXzXhsXdALrqAYs8VNnz3qguh3FWNjqzsmv2EpQjg4We9wXcZawDP0l7PUCGHS
ElMZwGJ6WF2ytZXYnhvKX36PMBzuj1Hk/YFJb8NF+KbWfhxy6xRdUxv4bYf/YFpn
C9T1OgTYj07v2m7a8YYo5DU63EwXaoHmcjCoa8Lfg7DM9/To9aoC5bsvrZ8ikBcU
HK0pRjMl7M1JWw6kvgAXY1lf7IGZQCXeLmy7lk5sOmCJriOidRF82v/mt4tRQ1vJ
vhAFMCPsxL0PQcChBEA7vO4VLcIdeMRT63nSoOMr0acrqvA4/Pd3znvKNNgLfALs
OQcJ9gdPh+ATtX+mCzx5WztDY0g71faMR86+ia1CUGmkWn0z75X4OulsJhPTHDGP
nNgr2+esf5KdLkzWQZJSa6zNW0owXR8xRjozANY6CI1j8TVE2K7EaI7HyRnmBmd6
nrhZHaD8oamXV7VP1iFduG4QSXH+Ao7isCReNV3bPrF4BZqwTTaQybyh77tGLXk5
lrkpjjMnSUtdhrpyrq2N0WLFr0IfXhCU3MWFJX4Kup+C6hxBCpsd77T/6b4mME3q
W8fx7S6hZxVXU1UP6sW1X4W9d488Cu2Zm1cxUWCpD76A74TwYCQz3ZSkwiKc1Dt/
`protect END_PROTECTED
