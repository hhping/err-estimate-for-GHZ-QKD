`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjyGNAFSmrhWPisKZX2JHb5/iEn8PQz+eVbIBPdxY9judb1P6G2r7sSWG1UEWuEn
LHLMlEumks5QoLF5hBmy5HJzyjy82maGcTDROUusi83XEv+kGD94JpYTawXni9NC
uHMAJKNUS8JtmbPnoKi49w8lRpXXVPFop7SaAms0bjcxlLAZqnndZImQd7GzetVj
hgodsijB2DYWFxUTKyBzsMcLi/MXnI37Agso2owUjrLBgRGBqj/pk+rxg1coaklE
b3XK7+Y+4cVNBrfW/uT6c/MeleTQqhVKh6EGtQaSpwGT2vfd89ozCnbk8a0r7cCz
aIGe6C9Y7gV5l+EQ9ivwUaBSAZlXYXnMCdPhPo82Wilh9QVB0XZOKJ1SM2y0Xej+
EuwwfLowk3Gsdp1u8BNN7NmCp/fDcbEySqHZMoHHqC4=
`protect END_PROTECTED
