`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X57FRRLSWsXg1UYrv/F0eAn/C14epjDm7MHmnNyEQV5ToEBNKAvjDQWYOK1VG7zd
8OVYfAnqLC6FvbARmIfGjfPmgqQsNireJr+RoUb3HLkl7wHWBWc6jnc24RHFDj/1
5mxJnT6cCuw18MMEHBqKHY/tdtRjAJQe3/RJuP2LWbC9WufRIuSrAk7SDL0v4VuS
TZUUCjY/Dkk7A5wCTd3uTN8VJkTSIo8EuGRbIeI5NXbll+V2rlI5l83W8d4Xk9IO
lEl9AdpeiSY7Cie5RyYrYoG3k/i/+HlkzXH+xV+pgtQ9hjBQfCgCKk+KOe+aNzpW
iLelG0gHdZDdj65P9OlSfiNFdYlGuJv7+/VTQ9su5IKL7ZYQGq8zy0946XbkyC19
ViQBk87eK+K4kzqVTjZs1cvZaNxkuwsQ7J//Hoc70F95Nu6Wlhw3H9xavkB68Pm3
mGk9MWDHZIjfvqh+r8QIdSWUNo3MgxxH3zrVLUkUzIu1z4W9XVBTNc6NkjESA7/4
5t6XswGcEhIgiHzLHgRDnk0Q6Hz6xzjp/Yb3AVbwsb/wMqZepE5dcGsbkxLK/t4y
+6c9ZIZthmUeHCkSJ6+WcWyAQdW1Shmm75kJtgCFAzEsoyAgH6892rmEbXgTToRj
WLmWzEgq7JJw7DwzliWXDQr5sdBIe/AoLJtiH1yqqIDaNVFsqNWgO5nG9OzUz5gt
9xYq3DXlJfVyH8mCqzZ03lE78snO54vS6GROxB+ZT+QfuOJkuR2QMPUp+nApdSup
4FiJ08+Dp7P06pREeUH9hAwoesO86JzHgQ2sP3S8t3NKwoAD6QyIUGELzFM4f0V8
buHFqZUT//U5C536fMv+7IzATfDoCcQqRyz8EFygIvF33Hxtx2/iCjB5YZoaloC+
sem4sZB+xPVfCzgDY3EAjgADXtN6PrNDDjDbVkk6BFTCDCBpRTApf6prMi25H2oC
Vh6Q3KzflnC+prfz7IQLE7ipXcjt8W4JqO6YWFiKAg9Tr8Ua9NTItt0TCv0+4AE2
wYcssWykBarNcthzvpRPAIFzfocH9o2fUGFZw14/N0MbrZMx3ntJhx2aZ+jjccsT
+4ey3eF7CJcw5F8Oswyag4F5pwmTpaTRF5k6hpQSgFeVtyHl3Q1Dg2n8WX8VliAM
eybmSSxxNJCLvmwkEXaph/la7SvbzeS7O4OZZbLpWDzSoItH7Dy+wi4RkbL2d/PU
n50xRG2sY75xhlzuL7zns6dN7MS3bQVckxE+XJlabzXS+M4vDfy4npOnEL2YwVco
H3yTIV9IiGWCCutvs/yVb4ZjXuzNwdk/BwrAOfmx0dGJn9kucxTtFYK8uePMAARl
mL3lsKKX1+ipqM7yiKNEANG7f3RmMCFRzizxTn84gL4b4qFpQjQbfvuBQYPeDWve
a/UGodQoYv5yI8/JaYV57+gSwz01JGLbz/87Gh2UqCi6iLRuvlymv04PMs/wJYPh
skKAYqhyDv+CLvlL6xx/IwmILe1eN9kjPWYXutz7K0p7oW037iqqerLqDEO2Ss6r
W0pTOQWj2sdY3WBos27eCQFYLmp9lYcM48vg8hjgBqbkNxN7IcvThzlG5PnJH7CN
HkXsdWaeDF1vCYsTEGpa8TBOPFOB//CkVggptE3OTwkKorC4MGeQMHROAcovvcE0
rtVR3291CEv7v850Kms1H5b3ka4z3pV/4qv68k9uPWNZ9SnTZFY2ccl7SEHjNa2P
XdFAv5/F2oNfMk2wkaZKog==
`protect END_PROTECTED
