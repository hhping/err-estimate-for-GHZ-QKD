`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c+sorTypWYsgdN1Y3coOViy4DSn1LN6Q2UX1O8uYhgWugL777383yGd7Hgtip6kg
QObfbwSZ9kb97LKzcwOgOPvoqXtuCQYnF6bmfSurL5vwY1dN5Cl88hUB60suTSu8
4SkdnLYR1FiZVfsBzzeY6b/JxwvZPjERj2IEZz69RPAcBdrVOLpx/x67Fgut5R7j
vfPWY9kouDEh4nx5F7IQ8wVlGE3+0OFi9Yz/8DDfK8whguKxjEeGBXVgdKQAeL/C
3tzFDgS4dw2oMcfSqdRrf2jFVom4ihWNW176M29Rw1eur0EoIeVjJ2oxTNRA4AEU
wyyiZGZiHwFSeXRVKaaRBDKKo4kOs5nH/g8IbDDKHuLV4BHFmhzkjTeBJ4/sNXg8
eLoGywPBdZ5MQtitBRfPM4/SE2OB3FtUarswGpG29DutUOZz5mFFn8juT3eFgdZK
hTh6OpIiZrU/BE+HYlkicsXYB3SiZlXul6KznQiGlpDgXMwQhGKWSUaU53KXzPMx
ve57GFaipe3yzlbQWeUuxif2mVJfSCOcBmv7k7b048f9L6wYwKAqcxrt/mVSMrJM
J8WrQ35YZ/1joW7QI9R4K0NfI+q4w/UHKdRczx2B1SKvEovvT4dLhpPkWz7XeUym
Q7kag0EgsloWKUkeddI7g0chd1C4A57W3Rpiwld7JhFnuXo06ezy+Ws0AjYy4gQy
OWSaGpF4c+w2bL9CKrmEx7bdVZI9jr6PJVANAxEzEIofHVrlYu6Rg7lHzll39O9G
1APEDMZBUC0Cjv1v6ZWn+k01scUkSCoCgV0KTwSl37Cs6yOzWXOqvxJlsnJRAHHW
lxGS8wXIw8j57vktKU3c6bY0/xWnBf09XidunOvCvetxJhXzliMU0rf0LOa9lydK
yBEI/L9P9bKKseELB5S6gMTc58ZVnzelNaf+w5oqlQ5ro4Ih6/wudj3B2E1HPepR
y4gKd6kmHQlDBYDfeyTpZnW2Rk9oP6L5NVjEUshJvVczoK/Y9aSlLhajFKJmPBAQ
dGWy/NYdbrkn8reWTedm6/1GHL7dT8h/QQlSVK4MmcySJhAn0p/7zvc9my5E0l5l
`protect END_PROTECTED
