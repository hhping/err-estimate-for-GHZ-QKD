`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uPiJ826aC/mbR0zY3IXX4qtLruFgzctW9YyMsOy6BOhtrbY3gYU79VMKH22S2Zj
luksW46o65TCJNvLskGN/DIZ1KJB71Mj3b5o30ufVhmRklWwDlL+pd+ITCjpxVIo
kFDcmDa0Nq9fSlbdx0wepWTXhzPo2ZDB7xdhLRTxO938mmbQ70EYkGha2kNxbGcf
ZRLvcnkl71gP+oNGNA1uLD1+tORjy8PWsE312xsgcWfvXkX/BC/Uzq0/SoOJnP5N
4PHvnsdG9Q437HBPzgTUGrP/G64iJP81+jd22NSnMgcVfUmAk5EVALee7rQ8eFyq
u7bO/ClYaEYcke9K4xghvqQadzVe2mJCmSEnPOqrTXLA4euSS1F7ifr+kfFf2wBR
7LMDrIbzrc1AE2CVKyJnDzOUy727katdLNJCJgBNUoiwyv8oCnUznVfDxUZcG2SS
C+FHfRHVrjUfbYuPw7ckgIr/fvIOiz8u1Kb4W8hmBiKSfOgmht1x9neVjPcZ0EEg
Vk/Rdq+QVGRioP5W6LD8li8tiLERFHx7fZ5DohGB63xVOd9uZtxjRQiX8AZCZ3Qj
7nsPx+WlBpOPhcYlcYCrPQ==
`protect END_PROTECTED
