`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCRdVl/5K9cBbj7bW2q8Owp1PfcDtNDChySkP7ntlKCr6ouBuni/uAdUvy0GztUY
emlKVMShVXu30IKXI/wp8XUBcwQLwopd5wFBaUKEdDe7+TCCd/ISzuJ3nltD/Qk1
FLMkZa2u6NwbSlf7+dUBOgp+LH317NDNjRzx8jvisHP2PsDbw4+4JeHndxzXnDX0
e67DHri2V0W4+dl2HcL9PE6YpsrliQJK2t4+BfoAfkHSzuCWPc4jh/pmtU0tTQq2
33jrQN1YJxo3OrrDaUK4L/MbpR0RR4brmxCJPREnJfSf/LjZI513p8WuZ0kwD8Dz
bpTCtk0KFA+xCs8cEotdbIXfGnVSd38CDXmMVxS3y6RcboYlLarFTe4coaWPWn3H
kWF1ey3l6tG/eikXXgUNKZ5WYvih3PodXVhPPMUEJ1pePxei/V39FEoUv132iTUV
RwlLbRJs/gBxRsLs0ak06OSlFbdDDe2uRwgetfZ0zgBox96WtGk9B9uYFFbYbDK4
aqyJiW40P1wq7yvixPWgCUg/qmr3S4zyDsTrzNa3SBtUGdwQDa6L4a42daNENzZT
dJSbU+1TIRUhSsfyUNma54vdVIGnA/7Qduur0oLz1FLvkWKtDT7F5WLtdRS1UGK0
5gT1sKLamQC998GnXDuQguCA5iufieWlupEMmE6mtZZ5Z5d2eCUdR73Mtde5jnM/
wn1CAmcZbsQPZ4Ml4DasyM0DlsLXT/kd35bOjL57vxUUNRWwKc0HxWI0qYA9AA+R
Op7fOpLyUpjIrN2xEaxvLLHDzV4PZeU4XniBPJRrtBOogoqP2Q6qLXYDUj4LCT5x
GQNs9jmgljo3REzZTEgblHQuTy6yWdt/q0wIX7OTzoKd4/cM73Mu9X7EYTqtRPs0
s1xx4L9s0XToNLgkQNpHszugTHos4V/9HrzKaXPAYwHaKs61fJsWDz6vsNAz7WZh
8WO1PHSU5+34JKbxulSgI84guIiQ8rX3JesuZ7d+m2sl1iqjp+vL4/qjHwn0fRh9
zajF60/kDE5y9rQG01/DUFLfwJ2FI8szGvbPaXu/riww839pnOe03Vsq8PetGwjo
`protect END_PROTECTED
