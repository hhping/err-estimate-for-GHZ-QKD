`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JraMCnJzJYWHmGJ1rYGPrk6+imasRtgH//cm75Zfmir+S1X4jqDdRyl2i5Yg3QiY
yW4D6M6JlQT6L15eGH37raFFm/OUslZf9NG3wikYV0cgRod2DR63q1xCWIoUrZoo
SPavwqY8B2+GeCro8/6xvnTJ8wSyUEiS6DHg3bj/AfnHAUuZjaI3ZV4NwrBvckoj
cfl3G3pgWZjVweNT1xOoMnOEiPPRTs8oe41qFTkSUCWWqzqyczIPbhR87ED70GUH
BVNkdP1y8wOEvec/ArX0j6H2ek3DGNz9z95JOdOSrFerV+D50lR2noTQkUtRg0PD
uf0MeawrnCSQQCc2eDPQObSZMYWd5RsWyEVf/ifnaN2k3Kr/ZSrPbCUrrh3UG4sf
KCdkKebGcgjbTJP1psgbG8Il4BHwjhbWlkb4OKAVQXubUSDIUTeQ/bTa5FEvqdoU
fYR4lnijWhuyhZPBpKz8IOpZWDK1YOpIIy3W5te22sStYD2MFvNUBn9IoHDzkYph
j7JUARQBB88/dnzxwjth9YlgvwBNVe9Sn8RVEit+LX35+kfKLehKjb7WHMRTf+jJ
18xzB7TkNn98R8RwTv+n9VhPjHeDDLaq9VAs/OvovDA=
`protect END_PROTECTED
