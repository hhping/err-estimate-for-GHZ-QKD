`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wLSg7BoUxK2yKSwej8e5TMznVs82kVEqIUoiXhBtAuMHHhyxVOlppcBZ1dzgbI+C
tcmhH9nUR13QXjb8XYJ2Ge4wXGGrxiuZpQ2RWxnx0RJHTmWBTHZ17Wrb391rsCD5
NqYINqgmDOjwVjRt6+4cxbjFf2l6aQihsLEHhnNJf47Erx0Bfy9VVCMeNfRJPXNw
rBAiQzxmxo7sS7rbe6LFwfWzfsSmS8qZzVTxzf+/cd0ptVn91IBLZ9YhWf/MSrWT
jdNLY5Hl3qJ5NOkg2N5oKNVKr7rI9hmqSPZ7FQQK/AeqDHWiFg/ZwrYOEQeEV9e5
waFxYIOviJ/STz29rbw026rsWLQNoj5LQFQJVE6TEcKH538OS4Ij/ImJk49Evrde
eQaILSyIPcKGorxSQ1AmIKZcFTuIyTYgnmKyrIwNM5v9I9AITiAP1Tt5w2olvePR
UsLdQtaYz6OOYNCVb8btQKOVrIKmZ9YWOqOKsE6xF9A=
`protect END_PROTECTED
