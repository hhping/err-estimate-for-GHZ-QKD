`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5BepWv+YmvKuwcVxSic4u9CTZ+bgSkkWrb5FbPaLaE3X0+HR5HTo9Bsc+hNyl4XP
Q27AyMeh19hN0hAiqgG8GRTNN219PgyRAnPfhkbAJhgZqtol2S+nKVla1anjbq9q
Q1WjEvHx4lTd+dSXD3IL+GbzKXxcvLnvoxgqC0PJlxBzNSmGMzVx7cqshnC2PdzR
nL7AX+paZcjz1KohYW0A2ApDQ/w1CNcJxLfTmXjO/BmGIF2e9QN1TJ2QAUwhqPgA
/Sr4G9lZqaTupMw11irtU6FB8gzIeJr4P3GRa03tgoJpaFOX+4BqjylG4AtUEZcX
uBw/X314lQ7W/xHusjALfQ==
`protect END_PROTECTED
