`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsnJ9D5C6wdGb0HO1FgiG9IB766EIJ4mWKHfWkA3pMZTodemL/FJW0MHCNEaqgfv
XYHUBZ2loiP6TGuiY3DxeDOBpen4kBr80N6OoCI/g3Ayppsd2NGFGvG/Gq1iyRbw
90OZ45ga6pojeaDaV49Ari9+PY+EojgJ27tXnd43nSdgnps6cipjyCo3Fda2JuFT
w+1kRTtiBZp/Qre1uOxJz8U6/nERC3K6lDcTtBeiQX0/K5xsW+yqGALPAOMTTShM
EHH5+Olzz6VeZigGYuzLjIeHLKvfMzDji1jehCqKd6oY9TjGNDJLzoBKSEpqOvH/
u98cYQnwI6RzUR3+gHbyVO9//eabZtEJy/LA6qyNr+M5EuJJSDLrBkFTPJZKFCSE
GtFyU2yQGEINrNVsz9VHmnnQUnLQwK3U7l/I4jQv1TT+gcsKpKyUMd6kXptLgEfY
CNM4/evif8cCCsn6h5TGnlxk/deT+tcv9jraIv1CA8R2jtiyvGbZTkFpGgvhTtS3
HKiR58sEauX31AIANi+35apm2ZeeRZj2LK3J2/5GBZGo9jCP5EpydJCIswPIUFB3
ho4ruY1Ygveavxws7kd9LDq8QAwAPT8HAQysH0iKXl9DsAAN3KGAvW0wsvQylAQr
KPJy9/vkGoOxFnZ01vnE/w==
`protect END_PROTECTED
