`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVOGtC92qMqIh+fRu8740ZhwB00PWvIVIxVjS3jvTK+Oczni0acBWjFz4ETS25xZ
nWsHxfui9mQ50VHkVVyyy3G9cWIF/satMSGmg1ONyuXAZP9JAkp0OWmEY83Gk4w2
zBrsb/21b9+D0erqtWdS5fHzwPKmVLHdov2bKKyCTOWkXjc7obhVBP+3ju4WtlNv
6Ug1dL9WSOACF7K+jEHcfndi6g9YW6TILTnlGmhCxbaw7K+vZCMNGqbLtwGLwjt0
pFsrDvciLs8fVrV1asIjuRzG7Ar2HVkl3TcvWn/Jbiaga/zBKBW3Yo5RpGUnzgtU
6xeGcC5EZ77vSnIA76H3YZjCcShY7jgukqvfrts1AWFZMfc5wdDmU/xgeLHLngNc
ZF4j4ZpmP+9SwvCu+yKt2WKuazfWaT8vD36niN3/mg28u1JdQsiD2b9qwYn7bSeq
rtgVVc0akmiIcmufds8WcCi7txSl09lT9BIYzDgiqCgvuocgGvIULd7M0cxSBs6a
ZgF2bcU3Mumu+hPjJUQwcLEK3yYqRb0ukRCCiHaX9KQLEAdAlnpfSrBUHZD49d3K
6dMph24TNw4ZGJduUgJdPm2NepCdNFek0n09wmoZ7mnEv+3GZvmpYxtvLQImlyLz
+ZnrixAtAlO0DHOlX1GVNDDZ4c/RriIz1EtN3jLsQkPKN2Zp1GKDhdEGZnU4TdBx
NLQOfKYbdAysMvGQ/itn+kDKo+3Ko9MOgRBrYx+NiTRiMESI4ZI9ya9/q9jc9q7B
LoahyL4l2Cp4ErEAcO1L3joWRwMObNLeyT/p/8gFEQuzXTzo9xx2FuPZZDBK7cIu
LvjyW2V09JQ9dn62CxG6sAalvKFZQy/yXGd7btAGWK5MrGQkJ6bEtVwcnOG+tLY9
B/8/xd0/k2DwkAyb3hz+tCsQ9M/am3hVlRmdF0TS7BFyKPLw+gNxVQ5bQm2MmAy0
iBlmbV2e4H2+bMKwQB5EkjgPaTskVgu+zMbatCKjIJ4ObmSir+0uTdZ3M4CyF58x
6kvAZGLqnkUqyWplEKE5kNiy8HoonJUBNIR318SbFzGNBB9diXtR6ina6GrmSHzO
0SENrYZ2KJopbg8d6qvl3uQPd6lXBLmnjjpQA1Ujm0LYNmpXyQwHWvsici1YPzXt
7w9NOsm0j80dv0Lec5z8WzdlUo9D+5jxEi8+pUlA0jxXTi5MCjaULnj6FkWzqqK4
30x6Qa2ldW6+8IF20Q/r/Oq1wSn64PBYSn8GKIo8ESPadxDFDwc4fRM+mvqjV2eA
pS17RKtne9hvLyaRqkZPd4CD5jKLQ5FtZYUUFdtWbVFYPsOGIK6j1NIFivVf4lUd
4Kn+EhViGbYOjms9s+HfunfsNAgIp2kISiIrPkB6FE289OmvFLMzwY9EAGZ5dAsq
`protect END_PROTECTED
