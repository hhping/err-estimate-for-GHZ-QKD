`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G68p0qTH5Kdnbn00UFc61C+NhXp6NMuINsmHBCjkiQOilI1ugSEH1P6WmYSOSOyQ
V4nbS+B4OZINztC+XcZZAhhP/cDES4gxE3cB9NOSEkGgop4kFWcy86T23voPmimd
Pi/zIiwcY6mN2C0adeFXFXFmlPJgodeF1vx/LaGQlfhtNA6S4vzICpuMtlqVDDrl
0CLxV652PjwK5XyaE96EOQ1ew620rDqf7tDFh1+7Nl7YrOrBKvFR34ba2LZFp0jd
dNCUhx+03WfQ5UaO5IRjE6czR+b0o6UN6o5Ig8SHw4qkSzQJCQkj31dCG90Jm6Cz
vU3WZojO6k0rYw4nwd1ZSeVp1f/wm5UjKjELYqE8sQZslN/iUWCsyfIbwxaFpeXP
1NFbiTTdMtxCETzROCX+k6EWG1nmEaE+pMJ5/m8vifjLiIe1Lp+PLGt1xotB4k/p
DD9mDg9wzChdgGjYOLenyjqy3fTshjnjEF7QefBO9mK4T/oPy5yOMiaop5crxrLM
UeVxRcrr0xQoznZ/vcPb71tdo/Xkyidw2C9HgZIKHifb1DNb/aBYk35eK/CHvV8A
GKg3O5Q253hGG0x3AGeCs3iakICKsO6NmlK+WuDY8pvy/CuGYvJn5GDWQTA86nOk
k/0DlMvCe21gYza4GmC41OlDqRrhXChYKRAJ4VwDqLicdHf6y7cDOGAvPfEvk5e7
L4YLX1CRHTMJlL/5A77UKO8ax4Hic8asq5tnraTZbUilwnng0ZgMObVsMNj1NUPr
g+aYMhwB7TR5Epuhy6Ql2HNeJSLCjphCCeWV7zFhxqrbc40PhhCmz47wdL/8isZf
V0uAYHbuof9ci7Uy4fH45vAT0s6B1LgVFLVGdmz4GzEhDETB8kp4bLOmy28moedq
+ZkC0MX1BYLvgEZzBzubZvqXmaJ4RjIpzq0kVVdlT8jljtoTc7YNt28ey7OOAey1
122Td7XxZ33CU22LtBLw5bKn/UCq3IxaACt/I2ekROlAtI9YXPytZzzxkhsuFrdb
Nme1AThyJYGIY5ZLj3PT7rg3WzPi8YiMG1XvCn/hp1aHPrcx+2cJpSGonLrU+c/W
vUMezdVQlBzkctkgtPocxpYC7yePBMGiNY5uy3F89D7QOVI4dVSUZNMsZqxuLHo+
4HSKDtfEZlwJWty2jLdQR2IKdCXFim3IgpUqNKXRJ5rZzjl0hGIFADPaiYUjzVkm
AZUVYFb41Ov8xt7tFIoeJwWWaVeDD6rcc0xUWCrJ63OIBQmJxIxU+NVob2Lf66WF
7Jdk+C9V5K2I6kzwqerjXmBt8jdoQ281pQpW3GNTpX3XX7nZowzMjGI3ZLs6fGRM
wYWE6dCi12t7ELLxz5boRocEtw2/84m2FRfxJdbRKUIpdgZLkvjC20kfjZxrqf8A
Z4oNTBhLBzsN4v3a0UnAr5zAdNl+9iYGFYGdrSk7rjQO2wpFEe1epN4ePIt2pCEN
MXPMdjP2BvPdefUUa6T8M3PYRKdoLvZbndN4QGCOdlXf+qc1JNgCW/8qngfgkhjb
QSPUAXEGF/KDRGK3RT+O9TGqPSIelYIdQFu3pLZLxR6uRlqxW3xCuzyxAlRX2+vZ
yWJ+MfGr/tSgyAdVvjGB0wvxu3e4p4shukEKf6YpTq5rUql8WS0Ww8GJInfra6rr
EYsujwW1SfO/8Tf3J7vnmqR/4vBPgkJZ5FuehCB6U+m6CZj0/rR1nBoyW/zJwEtC
EOpC1gVUZ0YPUmwoAIa8fHzehS/LjFKRL/qTAC8F+UQ3DbU0WehGlGaLLxjl0DU3
9O+1beSL3Qr2xLnOMKXKNfIXJ4P6P03CMatKnL/yScLfsWKcNw9mwWC4Nb6iWlA2
y6T6OCQHFUTKNGtNilLj1yV/EDSWjcmKdMY2tCp/vbS62FLF+D+Nvnfsf8Fwq4Pl
OKxwE+9HV4Ia6SNtUZqcOsLU0ODQ0fwOdoAVt1jEevgwxP7HlPslDt1fb68VMOUj
hDR4TIdm9uHtT8CHngVYC0fV5cfM1Qy4JGm1bZYGpxLh5IQSbYpWMpe1GBkgk1Oj
82xfGzKh98thv9OAOqU/UsNuwnfC3kxBB2Qx98cX7DwTjgIX4SjtZuK7xlfmBeQk
hgmjyYAzHLr+OJdg+NpTc1x7kT/4vKzdLG9JzwbXgOCyPYqZkdoNd0LrV8o4WB0Y
DDNXqAitSn00rDMF24XrCu+yAbzkL0MZgrSgSPFZ2Mi781Kwlnv6vAbByaVgg7dA
n96zAOLKaJfjMtir4+pAuEWYWywm1JNoLZwLh9CjTORzOifJBJnqiPm6QM68Vv4g
UN/vvpkIdRYUSioM4ca4/iNLnpPtuNiyKr8kmhnVvdZo14k4rSgfbUzDb5o/8aXr
z8S7JAbje87T2eSm4/yoc56V9tAh7u29gow6J5y/CTUph5tuitxwPqgjX0OWi8SZ
kuZToGCu5Y5UjebVyAasOO+bbj5qvs8FOa3nFxsFhknhUZsEKtJvEgznxoh1fFNj
JelFP3GNjcwY831d9uK4n5Mf0WeasD3joI68BqcGxZGzmgNWV0IRvxkxDsjgO0d8
W2y/zOnUgEuw9J2Va8KbdWgXBwmCNlZddzZ3P1Bjrzwz5EgSwO/inpffsinXG8mp
/lrHOzFaDpYQLz2bWhgcYbCrqycrfFLvp7mP4cNEIv5oh8Vw/wYyX2oSdy1ABeBY
kOS/sv48O3t3nVxpy6nhvNKDFRsT8VSjyh48haZrkXfZ8IEws50x8fdYXqOJzglr
m6SNCQQrejwbo66eSfndkn5g7xJwry4/OKnyxhbJy1fHpxaffh0bLkcKbO2ib2DV
WhL4NBoFkm83qasFUe8/35ATYo4tUVX2YgHBQ+SLIfegL+JRhe5FY/xWbmmOlIVY
CnNJzh9VXh0HJHYFrpr9xfn+uUp+fhtqluX4CQdWYm2b9XBn7bCmyNZkrHGisLxh
3Bh9iCpv8f/bFE9Xt3jMHXFcFcZi1pivpJL2ePiSAFGEtQRxwjDqmt5/zPo7CADp
ZR8PwCjPipTTWTRaL4hMwpjkft2c0c6opICrgLk23T6Sdy+3cHsNE7zQDwd17aSB
MDzePFpttGP5e6WnAbYg8B3ylwG3dMPkmMzODp9e6ZKWfea1+XW6YJTPFKS6cA/r
tQykG+OH/nvdMYXms3T14vQt0OFSatuHK5haR/JkSfNgVLFg8Q6h0e+D7GwR5D/P
1ehu+uP5doSTXhRyLwwVXzAPoAyELALAWpE0BRhsHbXkcS/xkTcY/dSeXrjH2k32
hWKAxTVe/ZSfpD0/Tvpr7JV+VDtUUy3NEkUtMLeg/50rYjSiGy+YQ0HCCjOY49hS
QAIxMHT5sS5tddV7mKY3KGqGIP3ldCmlA2Yka79nRreMZUWE8VrGA8yKdDjMpKlj
4JDxyqWw7ot6NdXnhjsYfN1Ieu2l7aEClpk4mO2cOznHWQB0OXiMxKEU6UOcAcQy
cAz3Qc/d9AfyaYghn/8WoRtxO8+QjsrfXKtth0RUCPa2BaYu9iNfvXoE722+5275
tm7ebw46mTHipKvURwEX25JkxdkopEbspucurnFv9LU0yyOX5HEiQD0/AjsefZ3c
6xwpYREGp+iC608u8qdXa3UGrM9ShM2GHysvOBIskmR/cICMBSc/i7H6gqtOSYPk
T/5q3UoN67e59HN8zB4zZ5M51b2MVMsM3TanjdFzCUJL8Vd81Kd+QbQ7rLzQtUrU
IWdASUt4reysnJ6RRa8DMPx54Rb+VmgCTZusDIjjBqN1N2KZQG610QnFVr+D7RK2
MVu0VJHrd3E5SZGK8cjoe3mSZPqQqd7wrxijtNs0WbljjaYduZAM3eG65zmhUOYS
pyo2NYSYpf11BmvWqWUaa+ZtFgkKvVQRpphOz+d0mveyK8wizzcGoy8ENDL/OUrM
tTtRpyPWPYABoJUsO33k5LG1uESDnZd8JY4/gAdCtD7jIWLGZg+x1vXHK4S5E/yq
V0OgSJLWvAyOf8beYrYFIyuoY+cwIzeDHxu0MAELsbgR/3cs9aJvf60XM5DyQ7u6
9sxt/0Vl3EmqLUFZlaE5A9ghwKU+r8EPrrjSOe9fC9FtjOfZJVu50u+mF+PXC3zG
CUC+prwwJJMgtyKTTz2GnoSY//Qks6vjo3oTZBZ6G9LmKuhcERSBChUOyNSIPdSc
NmU5s6CwQAPJsHm0d+bo4O1Rq/vqbQk01qMSlACvQP0bIxr0AGBzp9NRaBQF2Rlj
HCHhZ9sZ7a00fumMvrewECfU6WZQIDXCzfodPYxqRYOQKvJkD+ue45uF7AoihgeE
8rk2+8cj2LXiYJHi8lUUoPE8Iu3lZa7hv3cb9g6KiI4ntbBD7IzO0EPQqt5oYcFx
hZXjTm30F1jczZ/elPzsQH48qVVbBcYQJwccMlZje1/HGTZjKy6veKk6hiHC9z77
/f7A1B+gtZrEutEyIDb1GvfVjhII0QAvU8y2kL3ynnSDaWT+fHi19S4Ch2tZe/XQ
SHELYBpJ5bA4qTRsmRnoQz1aH9IoNMl9oic9Th3MFulKonSUHYjBxmIpu+is1aYB
yMseqyBKVb+4o9XTcppZWhOYt46660/mJH7z6AbeHizsnNyghLFO+hQ1IUn3/vJK
bj1Q18SxfjwIdQPMhUkQZr6x25KwxgJST+GOOjnl06sba+HOBM6WYTfAkiskG0Lx
leth8lPb+6jYnT7FdktlmfnFztDmVhWyOUy1+2g3EGdLTZC6whB50M1HJSx5GrBT
vSyClYCsglgcMVN2snjjzcV1HA5erFQYsaDCknkMIKKkDBzTGg/RCuaTE6+jUjte
2vIHYaQ3X9kSwz2LB0LQNG9KUTO9IWhMiwoundy+CtfKX8yO/BG2XMPcHk7hGlb8
JI7XHhuJB3Qtuh0wSb8a5F2b1i1yp5QOxNQwqJwaDXPa5OzYnw/aX4Ngzrt31GBH
rnfpZ3njLJ0bNgCRnKo9XdEsK+UgG9njTNbJ6y6eBsvV4+m5wRP0W6YbTFj79gf5
/s9VPQBJaPf7sg7YmX/i+pM2zz8JXya89QgivxNkVzyuMJSrbh2k3w6p/99Fzo7l
Y/itlP49JBcROBI78SqGD7nITTQE5J2cAI68/oOTmjXck0EI4Iad0x+dk39vNFmm
AM9h0U4GoD1eK5OgFNSFlkTIvmJIafss8eksjXch7aaAQIcVhRJnpyZU0di4/aHo
0jUbZYOIGjVkSyydgp09NavStcTutf0FX61faNI8zEbXCcCZnytv5QJf3yQ/R6T6
eoJO6faCt5AraTdnKbCOQvav2m2npkcZl526xeBUPxsdetM269dlzBavZ89V1d/0
+rBl88RvmtzpzcO14LyR1ScMErtSBsg3scnh9pNHSE5bUzGfjtUEidWf26WrjQmg
ovaqavUKIndT3jzZQ1TDtKhQnj/SNmy5qF7FKrB7Yw3U7TJ1WjVbHKQ0vCQ+XZoU
DniR1v+i7i6jdILae7HmL6ciZljejRUvYAUqtzkOHZSmH1u7mbvdDdANO/VzZdx2
UeQ32sTL/q1LWqWQ32t9+leN7da0ODxa6ygBSl/Eh/mRZ4NNn5Halja+cd6ccBph
McdPX7ZAXqvwJvAma7tcpJ4js53xlSBptfOGOy6fB4a4JAgdehS133ACIVRPunRZ
tEgRJ8oF8PGVIGWR0eKobi60N3kclhbn5OXm3DRyyeg=
`protect END_PROTECTED
