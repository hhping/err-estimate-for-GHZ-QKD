`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2bLRwzr0kBib9rPRxDvbWbQAXDzLltYhQm/jLZ3erYMiYoLF/dyO2whGloDUdvo+
TuujE0cIA9mJjfXfar9n/l8sn15c7yxG6Ep/tOpwMbRhI1QqzbnKgbyDKr6Z9Cz/
XwnlPq2/AXR2+BvZvvd66OWiJEJXthX6vTPMPHoItM7jMz/iD0ggBUu6yo1XQHsT
6ygGKpTHUk5kezmQ3rhk5UBAYef2iRoPAfvf3mhUvdotjTQIS+IYNtQfCZwN7yOD
e/4T5gLEzdJ46Epfmc8hnf/AgBAOAbZ3PTPe8JK3W1nEqy+T4+Cd0tHB/ZMNe/ae
oOEfw0M/uRcLj7gSN97NtyhtUNzqsrzWKZUPCj9CZ80EWY18dqXg3Ogc7ACkpQEn
A+6EdR1ddsCB9HLTt29t2prTSvsGXIQt5WuTsmmlerY=
`protect END_PROTECTED
