`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wwqcc7ov32nogxgw/CZGeG2JmTrzLDQvHAoivUL/htk2Bhufx6oI1qfM4tz4wcis
Rzg3UdbBzt/SWTmmuPViYp/gEtHBVDRI7346eubcmnrSJexz4CYpap1TxsrmrHvN
zFBu3VLbBUtEtAbUer9tnXJlZzug4M44yKI7aZn9vGyIepS1bV/oI9Dwq3uFhaPo
wPv4FmJjQaxJVO8PnU+iHt50FJu63Hl/I+BgHuI3GuMAdlPsC9o9Dc3LLFVinCs5
ZETlTf5jGaib3PuoRE1N/Cpvz3T6Xw5aIYJb/LcCPwuNvdvw4T0W3EOb5XrOYr8Z
koivp9ZPeMyCOu19bZX3vF6DDyHjCZinr1etnURUYs30B8Q1MSr0MT9RRO7ZMPt6
fghXHYu8PpRXBkTek0G6dXsrBx+CYG7vBI5sEm+Cr1vZ4f3v/B5qhoOTWO8RkBIT
33PICTaaaIVAOfhIO4ZmU0NSfge/3Jw/roER14U2XkAAjdluv23Pl3ZwHeTqDRic
V5D6xN1mfMehPY3EelpP+OQ4CIvkuJgTgHaEKngZmQZmZpKu+BQaOjg5yeiAFIDa
QfVDrbFsRRtJd4cuUtVvYhULrmKwiwkhjyh3UUrEUvEIIS3v0hq5Fe+jmdQqgkaY
LU0UzvlkX9aQfxaR8J8zhfh68xNWLL63sytNTdkkKVnEu7p06FbN/BcxM3XmlSRD
RTBxAwhepITe1dQmrIWkmz5NGh8hOS1WV6ChHJBDHo4akvLWgF7ET7/LmZJGiUnl
Pz6G0Cdh1ayrwpU45VBLOLfDgmR+o5rILhCuR3qrMTT8pOwrXRluj6MQlqunLEG2
PtVCFMrsDXFR+UvX0ItboYuNeHSJZHW4jJcrnkM9JN7zJAlTDd3IPJ/y7TnEnRxz
YRufiGGCeCJl8RRBlFzmfGaLV7lanGcwSbadWPz9F+NfRUh6Z2kv+A9MtLOg+STX
SBOzHQB8dW2pw65WQ6r9h/IScipYiwz6ZxMnl623V1NUDMAqDKLBrYrf6XMukGYg
tu/tf/og2ehxCTJo73rfOP1NOhBs/qEC20EIRMKbv/J5iQnt2uwX3ZWOyMGK9sy0
WHD/bGumfQMw6TbzuH4nECbmi5u+EFUgLGuqtAz9HxLjMqSCeN9uhtIuOmKJPWeh
rN3Wgsi9ubqZQBEWR37c0r1HVcQALCuTdJ9fhJ1jW0XLCdMG2dDYABtAcgP7v5sc
E7DT4ZbYWMznrhraK9LBGiCuSWQnn0xwUuXSIv6SantVZbTkz4Ftr0HfOMtL+Vcs
lAbQCPTBwr0Hl4zj5Fix9bEYe8eozNmOzLWm2/eR6JXFKAm+SVTqG7pcLeoyA8Jq
NTC/G6UNKZC4gPCmmL8kWHYhu+dKZ8qdSkBjONohtHbTlRDaLtLAGCt9CT4X+Trb
Hkc4qIXOiI3AwKNP7eHzsBmuhyo8XA+cmq20+fzqOZQ=
`protect END_PROTECTED
