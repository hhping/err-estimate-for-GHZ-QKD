`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJWU4d/fRAq60ieWRpvSiJVAlkugs3Xbn7+0D1nmU5LWVylEMRqaS8qkiRgye3eg
1JwqkfhX0WNTphCudK7UoAdYgBIrOXoqYgJcwJ3946/M8iIQpPVgEqwYVGtXgEDv
gMLwEtKc5vGm7klEkUKffkwfbOU4/SPmMrq80bMJ7VHG3vljJrx4wElIONpJ0eYi
7p+7YKpHDm11L2wDc4+Lg9/bJAKi8rcGrCag1NIQ1y4tLxDpaPIfU4FtPMnksd1J
IewxYK4jwhu6B2NNUXs1FzMSoAeBpq5wVoozHb4GqAKyBVjFLTSoeXi1IXlDv0tl
jF7RA/KQmKtu3nYSrInCga1fxDcVKwRXwBOM+sUuhqHIxTBHUUwuYMn2WOayMZG4
Rgx/7+Cu1T6aHVT+tKgzlF+40enBzYsFpR3tAON1sYqTjA0VboFwWVbQdCg33W4x
K+NLyB6Isp8pt6hsRm91lu75wbXkMScbBCvXjqo/IrpejAo7STxqOK87u1xaTm/4
1yYf++pHrLCZxw5MguebCaKMrZ0Rb3SbSRHenTYO2RQ7+DbLj20H5sP5AfANAVA3
XenWdeLqhGEMaLi10DHehHBrtv7Hl9AIPg0mwun7cF6+tqx4aA75JejO8zA3iLf6
6PFObfAbIW/RmFBLZQ5+xB3ABiKcesUR0dVZOjC85lXi4HO5HP1/x3n8QATYhRR5
4kw8HCUklvAWPgypXgyrzm47s6Y/krTmZo9jahrhGk+U/sa3+aVNW/JwjGVr6L41
dsq9RXER68pKjzKwJom4fCNDPqny7NXw5gjYk6Kdw/IwFakOdqNB6DEPLtt6JQRp
DLtOQLyi8yBT9dT/+vZ1QtZpr9426IRsX5iRFG/UgbuCVvPRJrjuG1zfiNvRgstz
nZkxBoC/nu5atVStR/Gjb5ul0+VxQ3p0Snn3GaJHbq0mXK08yEZtP5Jemi0ki8Zb
uFwkd66TUxRH+dfYq795mfcGzyGQ7ywtJToDX9BnVoWznQIam8j4FzZWW3y5vIN/
hJYhkVGdD8nyQq/FGzmCkUQMtOj6fhR0p0BF5GGsFlyZySMDo8tywerBBzrB/VGZ
BV2MHmQOEzRy6xFF+vIObFwPGwIgegvOisRtvSwaPW51j62++CZd2nDc5pwzTESX
FNN7A4v0/deFRlxjGh1nyI2Vpv7CiVOMM7ZZyvbcxL0CW+7oZynUgjwt873Y9qEz
TbI+W87ualfnTlYuX2285cgx9nO95q8kg91Ly5mWHDOOK1CsN1Wb06wzRr5DLIc9
cYoT3UC7UjFRbO79nPj0IdyhkvkCtK+6PnUhy+mhOu3Xd5mPo3n0XHEtbtLzKXyk
JlpvYxuiuJeeGHCvMn3lNZ+EpTRO1ZS613yTsUW1LrDAXTaIqyF3eYItGQIWaJ1g
kBlAjJ3BtfbJs2f3YzSIqLCt+43tUB6FuqCCjB75iaaiPjZoGBhe672p2iH7WfcJ
SxAH0EmFgfbd0suSl3xHLsoSFMerx5u3iiCs0KQtCwctAy6qa1lDMXLQzvuTR3kK
Ux2/vZlT5ky1aBNkQOtVyrjUa1shzzkQ/k2sFH5yIdsx9YY5CY6UtixLATZZR9j/
zNKCgGaf6hHDh0GCDfkNt9jvNlEECmh9AeyC4ax10t4M3u4zW5EbIZEM+/ZHqR6s
yhtjhCaAn76t+sfc1eZIX0ihLC8p0dUsZLeg5WJPnaN8a00zfBsrbsI39jmF9pK2
ETrnJVb5xDtHDVO+hn5pqBKsrBPX5UgUP4jCCt8IwtiOOvTQ/rVgAF74oWdIixnC
amApj1eIHdmGz/r7/9qq/9TzJSHjb16CqWfWyujH/7xkM2ZcZGnzXV+7XVP6UClb
ip8bRRUp7qP0GJL9fcUjKReR4Bgn6bbZOK/hwJBwk9OpeEAYrwTs3U3DaEmbh7Ra
YFiQsCYe1bx0uX7mWRhTbzUqk9gIjwzjVDUzCv5HoB7FOH8peVRz4qetQk75Z8DD
mr1Ksld05zjhz8NrhjynoOe0I6gUOBf8rQW9ubCMUCh9z22tP3RqEAAWTJXhricO
cLwpiCXFLRsKqB0yqZOOyeZMKH7AxSz2xt4WQwO7bUf8mGVNlJkBs56EZLfl4IH5
+yoTfy+nhJfHZShgl9Q1KRJVxxDYjZQPMBilOqbUIqYQSwbyoTMp8KVsrxJxNh8L
xsKxNJwKnvV+Nt72GPB0t9sYpcMCxf2ut8qw/8A4pg5oghTPDLfQTKoTUafR3A+d
KzGsvmBhpxgkxVykcByceTOSoub1jccW8rUTI4w8CLapJQjc3NDei5Vs5P0CX7vM
G0EM7bjiR62/c2o4p59l3L90bej2pXVLKW4aEROrI5PA1/BuU/wy9ONMrmj4bOX/
yICJlAwVaCiTseqdi9PNsG6bvWD05AgUjo89dYtihqPIYUjJG/rVwMJuIfobjGLy
T2sw94bkQOQGU4lJkAGyg7YSxZ96fWu3rrh/bNnACHtxGmjxNGwXnTqGDkibNN53
7sIuwXLMSARlxOpte7f5yGKxupltVrnAzuKY2k6nrKxqMXXud8/S7TVYC24wp+js
xX1ZPklEZvpDUCeJlOQsk0EREfpWFX7zVpl/sVr+GoQYaTeWe7DofxK0B6hSPg/e
fnYAZQwyr0Zm+UJ/AZKb2mPTrQH0EK9rJHxTgFtqXAia5Xz6PLlYyHdSdiCViIv7
Tt0qny8Jbvob7q7sXc/vNzbTUZVd5xO1WIfDnUmlLPadcmdlguIcV+gYKazNDa1W
nY/AzIPGs1YhTMYImWuwoCfKz4fdLeq4sE8hsXE6j5KLFoOjAU/oWQkXqTdfeyb6
+BOp5QDFAX0igzjgkbU9UoFm/riWCQr18VEdRYktPImNrKxICLuJvNvpx4o10ie9
MIcEXKimgQ9C2Sf+t/vRDrGL9NyFTVkD/oRjPUYDF7C+s3SlCjBfIYE9zeQwL4tb
a0bCEoaOa3u0DGunycZDqbrG+2+ilnI4jWhqxj1ss+5zwnIbwvKzQZnbxy64QFHK
rl9ULn2CN1gCqdK0Ar5PKq9CVWTrp/zXT9wQfwSfxrR2i+1GspsroGqu9WUvtI1j
K+8lwSmN+vLsyc1ec3+yDIO0Xb8yMcG7aidzb/Vlg10NnI5cnMiALQTe9ag9c5Rh
eYhQmvFMq1Vd7suoXXNqhOby8+XlxdK71RRnNDqt3TrOsysKR2oz1wormx/xSIfj
wiWVtzodXm8DNbxY9XPWBmJdIOOnGdH+LLmMXUiMOeTs0pyqPAx0UpQk6efDLHqV
uxkov9Gcv43jIR98l4aaSFNHma3P6qTBRjY9Clo3vWLHOPGqpMJz7ifphK521yf8
z8rPGugU9ocIHmXp1aikQqn87jY5M0dBNdxOK+hGtcFC4rI1APrRN5nM+3cHedAC
F6k64KtkBu+wkH4Dxf7r+7kaApE3Y/0nhmldjHebRBrqpQHxKqatCVRAtJhKxS8E
ismWkt6zuNSg/jbpXdAb1iM3sOqa0yGy6PP6UQvJ7+rcZKVeqykKbNrFcQHgIQKd
wF3HxAHZZu6IzmtEqspqonlNrCLCFaHANfiDtsgSyfyqYNbCVsXf1Qmfi1zBWWce
vVlOmkdYtMdF3fRx05mWuHWCw7UPTzZfPVtsntFIe0Rh5l5sDuGXf3vC2YFPRKIq
Doy72+khABLwAiUjLVD+DmnABG2ejRN/6oakHIgzWA7t0qco670IPLucStYiERtW
ZjnXUKdK2mupV5qFnGb+2gXkIBl29LCFavWpfWGVHg4UK2gm7+yMQZ+H8JKYpKOD
Bb/hS9cRvxGzWZVrAXIY4vL4OMT3TFFu1BEmyPCKsdL0wtNbEesR6k/LLysmEMRD
K61J8WgTNFzb1XaE9kizsDv12BgQeqC/5EPRy4ZgSM7ofsYhKTdGjgEeGyXaeyBk
FcB4SmfNn1sYSrXB0Z2MQhqoiyqzN0q4YcN90OL1VbNtWmERSHBblxe6SQPIW90H
kqiuMsvgNnu6MgZ4ZqUdf/rEEJqrNm3mwh1wiAb12tCNiNVp2nDwBEwHjXhYNJeA
nfEdtA4F8uYXGFLjj/tRjF6LlWHCBJ648fM+qC0vV/AHRcm6Ze5C2FV7EixCt0SY
MuSEmGudviuclD35lKmhNkQN2fqUsNrCRiL/udnXBTEOtTl3kNDR2DO+MZNhwDPp
ybsLevEqIIB85XnNmkUlSo6Xo/dUNdT1kWoVIiKiKy6rI07NjaseJ84/PDU+ZWD2
V2ygW1hwazORR5nbwl35Pc5Z6SiRXDhB6ksWqNkRZiCcuE8RZEvsfG+/1G69oRA1
2g3eJtQM2EBCdpCVZPVIuXJvJqeSIgMoGlUixh7Wd/ojdKwqrWAcL99sqap9H/o7
I6p9fnb2UDOgmm/GZK4aqQWSYAxbVb0LZ9vbfJa58VjXl6cXS/at96hU6H5yTN0Y
mOwpaWoD3aZZNtvmFge60033H7hkG2fqioElJBGwbvaOBTdHBkF3mG4QRf2W5yXK
tTuO/oRytulY2HFqOaTQlI69Zth/GHsLWgqTEOFLLFKWc4IJW841VWqRJgj//3dH
bqwfFUf++f4xft6OyzDW/J6wBTh61UmWvDIKm8h4GYYQCL+KSphmVdEi01RF/z9B
ofKPfouHBRI3LUFZQF017WsV+a5RgPZrVYnbB1mNMrsqeeSJV2nsYxI5P1LSksVz
nqBpNN7SQ/pRnJ6PQsrDCJBJUmuEb9uiFN0vabAXotxVwWenzJhT81o++aIG6IBm
1JP5XxQWVdb435gFiBNezSZefrNh8dsOOcs+6dCXJqTScUtPMzfEBxMu16gbPP6d
7Wmrsp1Z/Aefx5CIyiYEyoSEsXhfg2ZPJIqrV8RiwtioH3tsLq+CfxaOIek/FT1e
MEXyYv681YftwOWDIPEpK9ErXnEA0xERwcF+vyMu02r9rgEXQQW+366ylpk3grG2
c/zKYmRUoIOCaBdWqnsfPeBP0Lt7ETa0QKPlQHJSCXO0I33LGh8+MyuYdiJDigrE
p9UYfClwyxr6XK1GvRz3yELibnHbFSqReLCswK0tjdPzO13wMA1wCpqC5Z/m0f4K
eYRmOgzbYa41FuSTK/FJwTLFP/WAEdrrVirlGVJDE3ruajpOIxenDJYgU6H33NYu
blAhVRe0r9sRN5CyvFZaZGiBTaTDW3U23lGlMBpWGSmssKucTHcyKmOzcAictwyj
XI27lJjXLWdSwIuCaNoLePOlsbLplgIRN4o/fGWMgOfNEWM9EY5Ry4zzeaMq1aUY
I/v8sq/wcNj8ILAIalCxcvyuxbF24eBUopYm4Jrsj7Bh3oJzmiPDi90B9HKc90uD
ehvF2Po1iFckU1I9MSViJLaq8FNmLBlVN4oTPcvsOlRGNve6k9NYdORrGfbKxdXk
5CEW5XP54SMDTF7bhHHdIsjDcSltREkJLSDSnOVusaYVsBaPnTP230KgTh4y7DQc
eQZ7/AyY9J6KIRx8Me/rbmQIyqumsiCqaa+hra9h/3awsuWirfyvEoHjhITFpsK9
9oZYtlavZk06QJ3vP/QECItw7ckmhzmMYABAT2orOf9BeW82+Q75/a3sLvxRLqWJ
eEqDOhz21TrUAeDdhgdoIBWeP1PLR1PQgMYaURTGS7yqp0UIztBIFzo8KLuFWpY6
oVTx5cOTrWNismFdXI+/eozc5ZhiL0WDllJS4WPAfyZs+5ZZOOO5g8FApymaGbij
SPQwTm385MEI2P/hEo3C5Cfw0DMYcoILL1bzsigxu0eE9b6MBSlH08aIJD7tnhvZ
Gu+R5MkNRyu0GLi1klqogyvLOPM3WF7ayrcL/22T8N+gYz/yYFcV8T5vOauN0gsl
ghFAUU59Wrw5WVXG5XaxzcZ6r68Gx3xlIrrIYr3vbH/m09d25RfqKYsX7+9XobFL
mC+YlA/pb6JhHc2hyFJ6fGh/xIpSaR4gBtGOCgi7EM7uKjvDjJUIMJ1ygWWLitwn
AL1QpSTGf0UeH7sWcIjMZ58Lf7/1gPpMB07dqHRF866D9PJKVOwIgNUflr+sbQoo
16bV/DJ5w+23tW7Y31ZvhD1AhzP3CH5bK7aE4xSnGsEqa7q0hGhkOvHyR+q8fk3W
mFGn6YznQjFt5iKd6+WdzQhvtUW2G76lajvHjAk0JBQavyFmjr6F7a3vBURYDi+W
s/akjtm21GPG9XXNyI+eIJ37koFS/noR1D1LJtUQjs7Nry5vtxdm6txESmLQH2GP
U4KR5AMunhVkOM54gqvpm/9RT/OxLnGxPbUq6JIZK6whP6M+/wU5pbbl5hFM8LKI
s4bdhBSFS9yTXAJRL5BfjP1MrBEnTVViveaU1TXRUuch0bLp/rOFYTLTjFfg5/gO
1a8znSvX5ShhXE6rj+I/L6fMzbSIFMcabnrKoh9Em3gC+dpIWr8akLpTefKNoNaa
sZPF+Eywl/vXQKt1XKg9aCb2BTk8ADwVcyfTplbLXDvlbuDKQJVNC4Ku3jtmLPAu
2qeNklo57wV5fb1JzTCo1NyIeuv3JYilFxjn+P7r6ThC+XTiVKtF5E/mW4eQ9dFb
1c5+gbMi+4L2QuMNIrPN1lQfJqO5zgKvb+kJKzQ/qc+c50qqRosqfcNzg/jPXBo2
2vB1cszPXaOswxBURPU4DwuX8Qk4P59xieIpQKs46e+n0pwF3Yl79l5MM02PWutu
vzsIo9ZUtX1b0pHp34Vjj7KZUZCBctpuRGWrD9aAt/mbHBGInF0fbr8BbNpQ9QHH
IwOlEwsBlSZdmliXAQx+OmTkWXFb+ylwOcslWVwXoIik9yW1C0q/wsau6GFuzPOm
l2PKU/LqgCoUK+y/LIBeYWZwTNEOxYCJu3tSn4xTDK9/DrleRlQiTFLk1E+PwOah
ijsPYGoKrtrLqoMh8PawhYjIZyxGeBOq32zbuRlEzDm3u8hPe4eU3DkEb9g2VLhQ
lznblZDtKpWSU5IDrlCa45iYJNtV+o1jIArK8+mogNF027mWD/K6X+W5AVtEPNAz
3+kiPAiFL749KLycmM0xtY3ty1/KttkHn8pnUuFefEzuUYpvSnP5yfL4ziYufn1f
LFqbNSuxuDNaB7UwJdJxSC+1Wu9Wz0MBa+nu+1Dat++5N0d9nti83OradLNeCofN
pNdxv7I+TGid8sGLsZn5QecvG1wxn2eOM6EcuOv82367hnnvVGo8845vtT6e1Uyr
ZOcfL4bJSnUJ0h7PMRp6ud1IG2nO+Wz/pzkDQB3yuCkm7sfnSq+X5xfJgjs0gyyy
A0edUfIP1REgA7P+L+o30BesbeqQnT8UI8p9fmyVv1sTjYGLkIUCloi6ru3g3LUb
dK9qPbSzWfFN7Duned09LjGgYIcy7NAfvYn64P/jub2V6Dw4+Lnk0/lmhVINEpso
VDfZ7NKf2CeI3w9vin7lppM1qr5gWz4FRcy3CKQxsSz8WJHKxyy5UTpu91TPDAaK
VOehMlUhxhXLJa2/UxsS8h3eSTPFBvGm5yRlLUZIFK28IxSJloua1xIXl2RrLsoT
Q/Vb63BmIL5qukD+OCPGWrL9Vl2AZb2jMIm2t8N96mCwNgtvoRlp20sBEz1PjxDU
aQE96IZIOn35Cj5FK49zhmu2Yu5FhwvhVnJt+fZ6uP4coeLVMGUN+uE8EIv1hbPQ
Lj1xdW1HIOCAu/SHmD2ZwrCoB8t645LoNMQI+rpycCvCFYp0Yf8x0JDGWHZWfm5w
xx3RbWmWIygtBtw3FmVwQH+anLmyfbe0Q3PDlCY57P6oMOZhY/9qREIbfrt2svEr
mqNyXu76G4ZUrOS4XlC4Eo/b0y9ZEzd0KLniITLpfqgNjvrblpaOEoYHir3VVL3d
6YYd8dZa40nK6lXcPytZKnhvj0XeZUoe0L8gDtDckg+00wFO9Z+cdmjFbi2fAnq+
MCosyXHV55O4XCmRNk1w7McceFSe5dbnNjMwmU/c2RzPtrYg107P9eNdbP/Si7gj
bEY/945OsdinkilKqJrmX+ItBR4GPgdV4k+uwTAc/f/V3OVWIuLJ3i1pK6qvGaAx
wky1oVA1/LckVDxU1IVdM4vMFfz4AVrFjr+VaXF1RHDnRwPPOacovKSGRJeE1NrA
Nn8hkILXUF/MkXwfSypx5sbc/S3BF16ywd3L2bcWLh1j4fcVtNEtRC1Jju3WXZEB
Vm9mX4hgyHRNUOdTpJP/vLMBXBtMwEu71PHaNfwn9mWNWuUQY9np+R+vxRlrt1iX
LYQw6OCGOVowe4uAnNMCyPMTeZ4XqIY3q7hGIMFAjEnGhRxGFw4xA6Jxwu3c90LK
mZjK8TXQ5EcmNZKXneo4CeYJTGLQMEn8QUyTvcpEzwc41zrgFP6h15JIWHVJzESr
F2QgXQu2uULeiZVkkBUcpDl71pzALmQD2eUS/NhF9gtqXg+XXA7IZiMVzsj0WJjd
PSG0kF20IeUGoKb2fNOQszwDhKDIdflbn2XBi+cRFbnUeCpMQ5PGcHa0XNg8YCdh
2/lEFxDwH4JKyTK5UaNmcSPTZGyMQuXIyRONIMEbSOP2LUOlgTTGqegpR/q7q+qm
4kcE6CZ/tGVcYUZnuzFEOnqa6QlZH+POqq55254KbUgnUg7EDKeJAxDpzBVyrFUj
d7ZIbHVTU9O6f4oFpQKD421x8NQNmyrqp67gJ82Xc68I7fCobx72vsbuitVbvC4T
MtS7hLZQLkGNBxHVkJwA735aHqZ/NrdyEsRNqvZhVUGiBCmEc0L9WiApwJT8HLUS
s5IfMfKyaF6jGVMHF2Jc2wcbnMAqfCKEAJTxm0YFUm7+FuEf8KWG+DNlyBw7n0bd
XSUYCJTNhUxTa2t9Aft8aCpoatIaACyKQhs+6Op0Xgno/3+b2EFNlj6dbyekUCfe
r2lBM1vhZIbji4b7lahdk/nBY+cE5BgLt2dFH0ilAuo95+L6mSDiZW1PtqRAG0nf
glLGUW8nLFoIcnzVRM1+ypr5I+h5rjEYu6O39TYqYjnsZgXMKB7kRw0EG8GA0bB8
KSyq2X9ozghLeD+a9cf7y/q3Kyl0tjCG+UEd2bB2ootQaW2ztIkRIOODhwYOHsjk
Be5u2m1zhevLL6CEFbSiDQJouIkm4IH7rJ5fhDCRpNSokz/O88z+yLx4e/yOtGgd
UZDSqQD5HmG2MpxIOJ/jeVdyaXbs210lu7nKXlAPfEO8YGqKvYEG48h6VgREyYJk
KzgTvmG7BvCojb12U02WUnRhpiV/TiabWZqnwRnBPIgg6hddasgN4tBDDzSdfoq3
ZfXicKctjMkaYW4FA7Sh+lzJduFkSjxpvN4dpE5awecqvqKn3IYoRhQeT9Qgro5L
nnq4j5SSa1OpUTnPcE8ZQYZPAF7XPo9YZ9B5ko5SbbvM5lB58IbATgTm6c7G+vjJ
DiPOnrzvbXweEMEfg3rGrfeGBTq82EIJbKq49W5/BajIxakjOM97kGkd3vAyjw4v
JsUfyWtULSYGevnLtAqsswzall68ku3MwC4/oELvlqRFc15oqB1d6uxIOkQvKSn1
l0piVwoKZO0F1x0OffQqVXUXDgM28DoRKaE614nCSBZJCRQBm9cgS80b0EbObBYp
Dk7wPI6IyFR5BYuoMszEg9ST4GwbF81VfxEYo3ojFAKqEYXjDy+bzadrm/dCSi8v
RRZUyhHTzwd2vhDgOBLj4s48PqWOFto9MQzu6pVPJZGyjZVBMZYj52liECaNg6eY
Nau/OFlEiYGwtTXP65RsNA==
`protect END_PROTECTED
