`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3L4Oi5ShMLABcZWNlZzj/LXbFaxy33Cv1uo7ZTwj0TjfNGjQDxKJ8u4FbM/swmgV
cGzcAv6KNzwmyX9QghshFpkatXay+9rIz9fZZMaKXsB83/yaPUlwxBAQwteEaswe
pQUpXgzLRwEiX54iePxkI8GJwPYnJEvH/AxBu/sbLLs9pHuXIdWydvL3kimKAMss
yVONN58Hfd363n3XSnZxBT7ipDiAL2NL7dRC/+/BZQUpu/3BKY/hEFamSxKZO17E
kqHowGVl5ELviK4BUCUoggUaPETUHVTjcjGVZbopr+1KG+3B81w5NRFpQG4O7GdA
5qG2zlMmf+SXULP6Oxr2GVb8MTcngWswU+Eu30wF8QfX0lcKJzPDeA8Pi8b3FYZM
bogiGxxh6GbdqI5DcmswGoICz1yl/QKlshkbARKXkt58vKSnRrWeXcr/MKIEjtmG
byCOV0fnlCC70OHwL6S1D8Oi7R4IrtxVZrbUDWmDotM440OgfvJss4AKwRX+cyob
4CHXl2VNRIiEiVpp0EOzO9qW2e4YDuRQ3+MfFF3R9Mv97+fl2/u44hUeqaepVO1M
da6bjgdQsFT8ACCjomL4b86b46QzayQQIqQyBy/sD0QAEea4Lv1nkKmtJKiCYAw5
`protect END_PROTECTED
