`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZe4gUscB1tYrFKv77/SFLHZ3oEjRlBP2+fVnN7nhxxlIbzVe4ByB3pShJjZZgye
Y7gYkTUmRQdgp5Il1hDgULCeMc5kT7PvIL1nGLTAkpWHGqYs5PfWMhdFe5gXcHxE
+6cqbh2nJaWOUu8xr8Q0pZt+BjKrml3QqmyBVPRLiB3QkwrpM62ODg+z8It6nBlC
5DFUSbEN7oPgxCm/m6kiWobWYHw0MclbsnL8J8Kz5uMAEbOmrXMv/F8IaZ4UELwa
OsxiX40HHq4VbFdQrPZrq/1tavSgyFPGTKO9kuVqdLB010rcL7flxIJvdFKPg8TV
irFHFxfoMUvWKZxYDshFow0oZIjFtiJDXB+pmNFx17lQ14OtJxwHkuna+rX8CLqk
QC6DiAH0n00JaWaEFPO2OjwVR2Z/vOCj8dq3a0NKRjqQZAHcipIIBMpGUwCiOohu
2LBBq1f0DzvCNvdfaij+Pg==
`protect END_PROTECTED
