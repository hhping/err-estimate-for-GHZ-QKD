`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CtOuqngXC0IJtg2Q4zoW1VyBar/9xX2NLWdsrj/Sqwpc4ed3t7lzqmrUmXibRvX
PkqzzrRvBaW6fayIMZOCVIK1s1fIUYLl2W5VmfQbXrjopxY8xlGaDGlcXS/Fgzz0
xKxlEzrtMmSpEQWy7avT3MBA0eMYe1VYde2a/AQIGp5WCAD7yCNOnUZDjlFE1qF/
HX+M/IthRyF0oDFLkT0ov7nQUobjeUQSWsbDiCf8jSE2arGWUhI8BhQwUB/vtbHO
5FDvc+uh9TJNkgav4cCYblNZxMq41AVib8W1iHpCRI2eBTJgpYsdsAsjNh0KBQ2K
kGGJZGavVAdqNkRVGcf6BL7Qpn4Ns6FVMFH0q3Jyu6cHkUjuaVqv/qxObTWcTtoD
SeOq/ZW6rnWpC1+R6OeVTnrTNXmVuXYgw1Bj+/l9urtjQJHdhEaRqjb8LZT1r68P
/ZzTYyd+ZsPSKskLSKFqzq4JDwnyQsCiW/AuVVM3aK4eWDaLuZPkFNcMkgN2ivMk
qTaCxR9XP3U3LsqHZ754FuqkknAdCXxQjMZVW1azVknRbs4lMvCr0Se/6IgjbAz0
atE7MfndkV4Lxv9jtf0HovaQQKQnvZFnh154jtyU9hi8hlnplYWwRaPruLcvgnKa
bt8rL++8AcuwAOzw/3FDf0BZQ/5I/QwSLj2xAVrBwhhcDEBoozK0M0ZFSClh/9DP
shbfZlG71BcJSkoImBuD90qzVDq3AigfadNjLvraE9gZ8EtTn+ThmEhFSq8Qmnyh
QzzPPYcxK5w/zMfSbCU6iQy5HTz2fZG+VYenFkvEvNAlHmxQStEM6O29AQnWRyS/
QZk8QKX20ut+dEysa2CMY+59by3+V5XoiyuwQWc7yM+P36iUiOIEsYkihwuZbwG4
D2D03VUmmDc83fXw6wdqRlE7EuhArQFRIbeIVdVva5FzMT9Ts2wUKlQg49uAO9Mu
WsA68l11r5/DXbaW5WM8y+2DGgM7wEDBj9gQ/cwKlCKFCaomAeUdIZHbk6cYYeNd
SB7PKGXFVQrdcgmpMt0otij1BHdne8RxoutO19sCcJtv7TcyOYRNMOUlEXkug0b0
aztsbVpbTzlCEevXFNHr8H1vLF2/viB1dAvfltNRTEox+6l5JbRJy+Cotl4cs/bk
wK0/V+CKFjEK5ziS9OEKsuhWx8wRT8kPiS7FovikrwSQGJIQcG3x5TF1TOmPl1Fj
FEUC/22eAcmaFThRmMyhVqZLuu8VkXoS0PT/5PjZipIXB2S7LA6kN5IIn049S4Mb
Dj08Sh2tgccA/CMPsmcidK1P+D4ztL1cCw+v30oIDEcnEAzdc86lW0VMol57dHm8
JYbcWzS43Sl2iLxLA7K4g8rrmIX7Fxvj/fX8DrvOk3Nd7NUS9UfZ04xoW/8HeH7K
TJZYsnb8gm6pJxSRufZCPtJuziqLyDKX7QlqFZTw9kC/wXeHA3EJpoM+ljKmi7ws
jOQPXCMnD6CS/Sa8coHeRHmQvU7iDnHQFAX1yNhrlD5bievolWBYKjqfcqYDUYyJ
HI6EjgnPDHFFrrEwcwuvSN8gtKH8ppCzI8Sfp0/F+G+2Jrmzsbc02cPSaF4EBniG
qM3FjkFLAiMkaiaduOtgWMOULbPc+4n6TMYkXb/5Gi1i4r1WJJ3NOwMr/3LCKw1A
BNa4a1ug9GLF07H5A8lC3h8OCOts5ZF0jH9sQ9YqbYYTnRn6OMAKW0p/FFjSMa/M
Wi/GTzpsn2W2fCppAKoIfAaABpJYiFxWz3oiGWCyM9iBJvE3orgt6lhR2hCBE8XU
G+pLf4OB4kY/2HU8mFZo0CY2ND5pVDF3qNrCPth6WM7HfqFRzImlKGhkm+KJDTaX
ch7l26eC9JppNO8qKPQii6uELEtxOgCriTvlyx9fzNl3RSod01M6V/KzwVzgmuBV
MXDrCGVnjAf3HI7yV99T4m+daB4PLW1x9UFPiFAKXt+w+RIlUC4KFrQ9CZs1+4/G
K+TZsjE6/Aa5vGrKWf6Y3FP1YD0V+NxGtQSSSX3OkAd9uc9EtCNFhubqHcP8mR6j
LET3vzTE2s3/abVzESIrr3ufpt0LXUzeioKsvHCmRYOfn/CflkR05QObMMOoc/GG
KvYKvmMJCrEfVh48PHjhObVVk+uxdIoCT4aGc4v0WuLItVSZHpaF0PixljTyszrl
KvYM92V5DFMmkcbftWu+OIp1HXbcFtZWsRGM4N4KPjD6dVPUPpRnCTZN+B4mcMlo
0gxh9zHUffL0xoL+BZtO1Zby0++mvj6l0u04o/UlyQEDnIur3PYtvcUJTZQhy5UA
sUqCwgp8edKy08sOr/TPgv5LyGSKwfrrP+1D/5qxDX0fGZiE4znlKQTiEdyPkqMN
Ten3+UHByNihhSyc16Ak1ut/zG+UscGzYq8O3Jd+4moGWEwZyhvjFZLG7l5ikkSE
TabOCYmcbDjgW6VYKefC7a3Gn4xVd9ahgqXiKgLNGsZnEEOcDHfmkicxHNCyx9qi
eZvCFfKcOSAxoBSIdn/w8LdzI25fdnvgILPsAblSUbKVyHR3vzgXaoz1nSk/++VR
8mGINXTQbOSm8e00K0gxUmBIuJUlqVZ84AneUWZ+fcbBWN4R7DQ1aTyCxOmYzcqV
FdTmDoicM9+mPRdihflssBdZD3PjOzgqBE1gA6bQBG9ujJ93q7MzChjNpa2qLfQ5
M6r8uRdG18ytSDizeZdNG7UN0ibDe5nqMG/ILgPiSSbqaBGTvidIT2VehomwSpW8
g3nqhw0PTyFlZj9dx4AyvbnQg0TIzwECIp0P5IHou/y3Z7VptkhcnNV9nHeCeXg6
EDE0pS/hDzeu49bz+Oc2SSOCSWjb1RSsV4glG6xlCg9RVpmKfmvt2F7HwUXSh+NH
iQSJqBINoEwFS5OGZFP29tfHhS1zH99pjH/Vmi1g5Rw8ctZbepI2B6GF201anGDl
RQOVkU1OlMKyAK3q6k7BQT4o8Z76aae10gckXkgwrQT2pzrFsjEuWF6UmsaohtKs
RqbKTEsHFh7MP8NR4p1fNxGda55hmwLuArUvQVqGsJBmxZ97bzuulzPV03FNbCjr
H3WAuws8fGyDHIMR1oYNbaZjoZ+TCcNnSpry2ZZB36z5bheHoUOiuLnihhY4dPch
syJgJxEDKa/5p/V+ynMrqw2NoVHnuJ8YmKQnVQ0Rd3psHojJ8T+QhmLL36KkIiG4
stvmyZabYLvBBJwoyrcT9BEUT5qhUEjIQx5LJFz1Nky1resFK9aHdYjR5z4W7qdt
AYBE6M129KM4vw60oU6JfknUURgHJHxK1SsQ2HJkereT62gVTase1f2bI+h9rui4
9GMXMdXESGcMLjiZm9ruxGgOaKdKAkGbMzXNBGmZZU81+1JeIIhmNqj7Kr8URpIf
2Bjt55XWgIR8LvFKEslSZfZDzeuPzmac7izpODlG+f+kf97V/U5x8FS0GNf3MkxB
fG2i8XHaMtn/B+48fy23cldlIu27ghpmMXX7Za/9QtsVS1swJTl5NL553AeGjWIK
WSqGBJa4ggN+4oihQ6eXn6bcZtyX3uMdBig2FTxfRu00plTF9Iis9XxlURwhYa9Q
7T1VlZ987ndXwr+it2NVBbtXRMFbglc9h6s6bAhUt8/bluOxqb7KFKIzbo7mCQan
VEGzy3HO+qKgBNLLN2u/G3HaSkwTUWlJksYTy3Oj93+S+VxjyJqLjE9fIXnpzhmv
uffttNr6SRenNieWR125BZO8RE8/OPlk5hv3OYX89MklTVYe550zoUtsMs560xj6
SZSXTKFMbXijbLdjYAn7CUiI3duwdZz137df+vp9cpq0iFNQZcLNPKxWY4Jn0/2x
BEiCCsMJaqFR05RRxCGUahAXb/FgEkV9UFaiBk5O2YXe4u1CezLIprvSFr6VY1MU
9PSooScphOuz1wyvZ4vT8EtNqgc8LbmOrEypZMpcvVUqjCi+RgxWp6+8zYx5Ob+T
hXxCYH7o/Mzx8kmJb2nKvCsWGROEoGCKldICUL0owe3nrz0t88AKtcLF4sywN0ws
VwMpxd6rZqPSzrwEtDWGO4NbNsrKH3JfpbPJO076RRXJpRJdT4v5IpW8xYVbTie+
bfaxxodmGcF3MC1fBjjklYE2zOUt2ekQxZNgyR1P/adjjF7NgpzLjKDlgn+lkCHf
jju31hTtUgKnAoQAusGMPRtPRc1H8wZb8uiqp7NkiUPcgXAtNqZzMsvb87QrHcO+
x6r8tUXzTpDg8wVuJVkx622nKZw1mBPMplwCE6boTx0a0TTBkh9uthlmLkQbi8Sp
dWNZGxm+FLPDy0UljFLfymizKBIAaheMaEtMl1Es01OSpUE3RBilw4CxZkK/n0rh
m9D9J2T62O+xnzhG7zbwiMlPRTxBAdsyLcaz8WhKsnc7wvUqj0wH/a8NRDQc/SJm
Tdi3t9KZndW/ZO/JhX4k2gJ7F0t8DQjAaXR0Xj/TbtnGlZN8H7R7iw3P/TaMkb2H
Z+6qeyPwotTu6cH/olqcrvpBrYSbf/a3YGpjA6r95aV84MKSI3LgaoNpn6Zgwl14
YYEuuzSQuGCrYWla23/cCnTWw7BnOVgqdYPmnExrd8WdTThFHWFpfiaFqUdtGa26
aG25t7QqLoQ10xQsJDyrk8eOwgwtuUU4rsK9/drd2lJUG3xpcHXVZafyk8jmLniK
KSTvzQ4aeOWKsGyBxSkvjlv4kwQVqzctMRuo+QnqVCrutOXgP6a32g4/njuZqLpk
CjAmiH7rPazO+IaOYNF45Jwf8BAlmRAoc0TIXLgebOAI2DTGOtv9T2Q6DYz51brs
PrYoy7woKnm7+EiDEKw4c/XXf82uJn60D9kzclUl3azOZ+I4BxfxC+G3bm6HhJ9w
O//+IWHLbTl38qJkwzxR4qswukg9iwxd4Vbclfzfq9PbeoRgUsLQhsVJzJQGBp3f
Uoyk6bj1wmeN89T9BelkGzXuqfXFrx+CcSEs60xr9pl9eZG0KYzyStnrXP5dCAVo
I4ZYBYosrvPB0QYOUIFocm1PT69mONo2WCNfY7qbffHsnmC++1gKDpJF+eiUv+1e
ci+JYCQpZYo5JYVRGm1eQNHZqsTikAHMYaJNzIBE8PVs1JRipvNhhx3x6TKmuS+8
PMrBYkcCX0yNnI6Czkr/6dElq4g6lypPiTByaMWMW9E8vUmh2GmQbAQexHZzFriO
Pkpt28tXjOE3PuRn+H/x00NPoTyhJn2T9V7rtZFn8LJU/EWURdk0iQJRsc0kP7dP
F1m+1tjT4+P7I/2xeL2+SlBT4p1lr6R7ZPYF7HqnPz59K6LRwj3cSYuLznv1dS1Q
Ruo3seJqXKOQUEaGXrWe08x7vMbVypq5wSGQNub4N8wcsC1OF6uY5TAyuMTtNsho
LV95yRtZAoaCb8jqVtw0gNi4uGsqqYg4/ThYtTBFnk7JBXv4e2npSvOxKPLbhoOV
8su+Dev94HpnNTIHWm8XKTulC5YccknBRH7BiYhQIWVuNon5tZyqUGlRTQjDbMOQ
wnj+gq9VOtzGgKS1xRSKrpWcp9JkZUjuXH9hOhsa9iqaxIVkljoC+0fEfIjBC6pg
1NelRJ8oBi80COKGd4mRm1tES4NOhJ/ArPRZy7pX11u32Qr2AMihOZ6/uyjINI1i
0D6bUBrvEu38s8QkULso0XgLt/tTyAWbK42X2wUq7EGUnM4jLZwFugcSZZrRCNR2
IWHJKx+zSl4iiV68mLnTg86Du+mfMRsC9ocVHYAsGUGTj9HY7PiN1EeaXgYxtA1E
PaAldplX7XBLFHzAq2rPyQix07cJpk0neA9aXkGDtzn29ovUtB2njbJtP5jkHj9s
BLk92Tf5AdXGBn54eur8tX6EFCxWKfmQMdZqO2hlIpHR0r7ml6lXS3i6JWHqvcB5
D2k0Zebn2uzuZClzYhh8nVe4PGmHsVVyDdfyDl+nTzL06rcEtQ8SBP2t5YvjyWCg
ZjSycybvuHuOTHtLia9vMq5BP/j25da4iZXSDBHyvNX6f+BjN0HzPX/qo89IAONA
4d/e9VgC9RJ+8TjPWFH7Qw/8mI1bvAzZocD/15Hf4nOB4C/xOIuCQxCOg48el4pi
9f4mc0RAUOrWAhh0VFths3ezsTNzB3rYuVmbT2zfdXMNvD0u4YqQ9WagPChgYqyR
Zhj+lgkMKEiDM4Wf0VhOHkwXXx66nrF/71RSphXoZdEQzgRsStwgO+uSwnYAiaS4
NCx7PsSymQf0UkviRufb7cNIeGdRrZDwXw7WSQU0HpI/Ndul4MjYzvR2jfytc+f8
4TFCEe7dEieXkmLkE3XX+m3o+LW59DCaspu0BnZ5joscphQ6M/zDNO2QCvoiLjlv
QDVPUMLcUIMKV6OWnrTEB+LCL8MhCRpjSQvp+Waq8/CcUTeoYc0QT9FYqEtqQeaD
RdGBcue7ppW6qw50PmOlp+Ds6PEf+Mc2Wxgdz3lkfj4mSePtCXTS++0EBQLWNXvW
XTE7lbGH76yVjP2ldrevO0f3xP30UkORwDXDTQf85bM3vFglR6gPM46cP8z2txVP
I41fjjPsBp+muIE9CR26Tgj1JkQ0WCkgYKE1HV3Y6QkwxebhloYwB3G38RWnTM8e
OCdiUuvY4sLR7s/t9nGVD4u0tlTvnbkwMgtyfGw63HTYRxN9qnRBxtcpGnLlYLaW
L8QE132VTm4dqqVjaP9fvG0tw9j7sTPihvd3pdsnPCZYU+5eaXDF33AiZr0SSMvM
DORM8dVWO7QQn/hWNT7tO/IIVLX7tPSEETd5k9vyqU4Acjf/q1eIYu2Tk+kXckg0
MSDPpSF13eE8xMScN8qi6SI1UudDvAb407Uan+0hRiB+2yRYWwBsqaUzNYzD+GTF
SsW8rNF8kJiyUuPA0trN0plJ3FsDmq8/Te/IQAq/8dJHOsKi1XxZVM3pmmHZScAG
DPWlUdlU0yxtE7JV+1QL/VqHpMqR6Q49H4u7LyQLnXkCeHRy0cE5DSkXK4kB9yfk
b4EKqUFcLroVoeMLcvaeLwnblDfyjslW2hBHarbe75uF0aWWiIPsthZzpbhfVZfs
I6TcZieVfhW4tDm3IN8uAOWP4xaLB1c3lExXXHqpAKkTb9Wwa/6CI/sYaUSIpW0J
ZVeFMI5Z/XSMnfluZlz51y3QAAWEbFlmPlOQtncRbIHvVCiLNus6C9uGojh4IBv/
uPtUZB0m0fxt7Al677kgG/0IwxSih1tv2bVQxN8hnH/WcVj/SM+Oxyw+b8x0xoBZ
ePHusDGIgNRpL8uGyAYjp9iiGKwqNOy4ZrS1tdFLAevVzipcBja8stgBP25rvfMT
5XJ1K9kgFvMmw8qNpZWpxt46lVlg5bD8bVi288EuTDrA3l4+pdtDbsN94uGq+kOg
YlYOo0qKCGjLkjZKLTcfQI2KooRphN2UFiBEcuiO6tdZ08jbay5K/5vfyZ+ThdZi
6nko2QU3y7rZHSMLT7bqCWlCWjdIk40H1jWraC/suj4nCSjr0w9Qan5ED/J/a+Wi
cPO8YRF/g5qk9t6x0j7ucuAFUis1cUWA1JnIovTsyAERjphOwxSS+lLbk9BRl3w2
pkDi4Qcblf4ZsoPrqJ0Ou73jTJMq9CNo1jzxmv9Hgd7wVsWwBiiEbKM8BysLR5kW
NzzzCfjn+I/UyaSZs7Kwj01d2yd7TPHOnn4qIwZxtsrpy8Z/hnolwr/EKEwzt7Yl
9Brl4qcpfCzBmgLmBabJCIpTBah9vE60ztQb4Ma4M3ZPAg7Xxs7PKQGNTW6I1UJ1
ogLdq/poUi1zApZ75BlR0lqkut6lA3Fx6lkSwXlucQjKLYWeuCDrRZ1OZEUySdBG
wvZKwE4NOLL6jTB9sQGqw7nyqp2olHo+qil9n7YUTt7B9YdhSGB3+Lw4h8P0q7en
O6BJ8lXidvEdKHQPN2HRKETRnchN1maT6tBmksk1Wsw2xpwwZq5FpOGxyjtJlo/n
Fbp5AMf/L7JI/lKaR0A6nGevQYjr4QwjbmgHcyarPnC5hJ69EmNxpS4MD5XMIJcc
J9nCJ2+4xGvJecT49kFkiZ5gKEjdBu7ghP8DAdn7tnjMo7UKNKhXMGjJtQMIL0xm
iDp17vT2Ufd9tMkXlarqzWrCnlwWbDek/RHVWbjMndaHTta9ilDOhSX72JJavKwq
u8rT/9tAoOFcIKO9kF2zaH737g1AdWOXNyQC4/aYSprRbGaIeGwbWsbQe7d08Eru
s8VAw1hrTMxWTd6P7iO7wL9w2L1Lv/qSnWNvSd3D6XKtUvkMxmtAhR3YYv3Pcp+E
HmbNsWCfsyRvUGkpj9VzqiwWY2ngsp+LDvn/Ve/1OMV5MbLryqI7zm2Z8+pkjFzK
jDfOdd6mSyjRYzsSc9OtF/kJ1NL4LXjyhJfzPyKYGimlX8DOMPNUlh0Nzk2PJKBm
ETaWSo4fkHb3+wTmlZy8OVGug52FefB3K5jKj/QOgC6+G/sVMuEpsCjMeCmE4xNS
Fs0gkcKW6hropS0RNjnVf1kAAKX1i0wE/lwVub1tQQy+kvTz0m0/+A71SZ93l5Qn
SS6toHTS06263xhqpAxhPGkzpAL3z3F/LHWNd2CyzVvbXwkTtVC0/AVe0Df+s3wk
xCOTPFoM/bSlHcuD1zrhMUOaYDwHtmunaUovSDUc7IPYVwkxCaRMzrUb/F8B9H08
na20ffKZRo3oYNA+DV7OppircdBnjLB03ca9qahViYWUoDHpwqtsKjMUgxWIyf/5
IUM1p4EjYSUiBLMwiCZxc1sjWvFRmJVp5s2SskvC8orTPWNXRzEek2zVa2T0FmzV
AeRnGOLA04o+97MouRyHvrEvGvD63eCtQcdXycatvqg417BcQ6DLGVErrcp4Wfnf
rNmy/GbYbBIovEdxpkdRj8IDJNCp0tKLytkNAo1VfG2Ae0kcHc4BlAaayPLCmtqK
RjdNkJ9qeEz2B0KGfJ/2W/jMKXMKe1EzdpWegaMe1RnjPU5FgGNfqpjOXJBGwfTg
BX5Ce1owklwQNg25mGTR4tJyiQG87xqVc4f0T4VtLCPWuL3mRD5oPsbOyIER7FIu
agRXiPKQpzD3hOywhYyXne9E257OgdgvFwjZxslf/yqCZMuSUysHyAIk2u5brcA0
RqARCWqn2tGzj5TfNAGiTu8Wu0bWJ0bUTO9yFarHH0kt1rH1nraZJ7CTbObkY5Y5
WNPOi5X/W47ESyF25kZRJCHSA+xONWHMU0L7wliI5pL83LHPaEbAmHB7Z/THWFnY
qe1uNBoeLt+DgRL05nVAbNbPq0rFX5Ili/uGHGy2zS6OiWYS5dbWJjbcSPjmkhgM
z21EjtDBPZneJs3DI7+2IktNFuK3T76wWvtFWZV5GSPlJthLXR+sQg5qw3t2g8k+
9D/pCKXJxBNaiXH/qsLtL2qfNqFnrxjMk+naA7+dbh+3npFbvKVZF3LMiqHq6yv9
OXZ79jhgpSl/QyQiqLSg0h1TMCEfyR2HzCR5djUBnRN3LKw4qR/k94ebHwEeGDOx
egzb84GRxiPGEgmFncFEPxbZViMPpoPrluBPxHjdBoX4MjpnDlFP8AzfmYJzzig8
dAylwDJNVWFtsmbZlz8z5G3tGdN90aEVmhrMdfX3c4a5Ep5TIvlrxT+G7873pDNm
U25/D+oaPUKECaNJL1lvM9QdFX1qmXAw4UUK6AuzbW5M8J9U3E6VWilwW4mcUvTI
rbFF+W1ZQ1rI0h0+QIDuLRAlTXo2QM2RWTH8uBJnllV7rez43/dKDrWDyyVhAfXD
xf8KKeGlHZWrZBzRQNn5eAVeTzfFAB3S1a5ZuspQh+ANs9/8WFPr9zY6A/0Tu3r2
5XYnQWR63YzCjOC+UZaDF8R2vcktbgLHwf+vGYzb6/v1WZO/n9YTBMu1CkJHV3FZ
X7NU5dLxmHErkiB4oRfPM1vUuKNEULGxPnRqjDV5L9FObD449rMNKLuBez1eQRWh
MwKF+cqLzFMW0TZ79BMQP8QbeC4Fd8P234yr82euR/tPi7ULV6C7YU9QSmDnaIhp
XKRw4wdmkh8tPygJm+YpvrNO/Zdfxu9MN0RS8kqbpJxWMtVW+1WFVjXzoUh/r7N4
aPYLwraN3td84TtyH+NTN1i4iW8HkWWSdhrs/Knqg5JNe44X5KfP9ZVrm/KIUFH+
J6Gpl5JZdGrN+5NbxGsbOj9EdXMuYlNugl+j/h+CxxLvUg2JNaNg/5elfmAUz0Om
fIyMlZRy3YrNg2zNp1W9NfVWen3F+B6BtW0JTL6cqtBNQh4h7SOeSDk2y9bfg3uP
HqOBH7sMzqTNFIfUxuorX0oduVL+lLd0JZY2OA6q5yJYxvFmqcuT7d8q94FjJT5/
q+71whtFPus0SsMd1xQXjeBLK7KTgT8ZwwKwfP5ZvNj6ZhOomh1JD9f8AL6GSPsB
Ge19csSTpmEQxEWGJrqOtlc+6kyke5M2dH+JbHXuHvAQzSdPUhPFjqPV5nmMDjDz
Nqm2CPWpgeyAikdgXwEaWlIw1gHJ1RJfQWzHjYnA8FryumaSeK6WritupOEjLw0v
oNvAVl8jjGu5AViuQqfCMPImiqqpZH54udy7n7O1ePTIVnpJtQ9FLa5LMh49o/xw
ZOlMBMNzdxmbyV6hOQ4s0RV7BuZPKmKP0g+8dj+H1yfVXG6c4yMKWtsV/QFzqmdi
bj1C4CeUgYhkwkuF2Co+ccr4859ejsHM6qcmymXv16EH1CG9JIxrOvImZYsXbMmn
XbvH9PibW2S09fRlZ+w7W9b8x3QUibFZt94B1YPvv1fXPFPzPyUbo8zef7WlPLWn
1AvGcI38RUJXolZeIDZ3lpNm74xoNSzCY6s+XrgnfELCokbbzD+E2CNYB0xo+YBc
NpXelLsLVC0C5JySwYa1oCBZwBHM0pxs1ckhMMy/nyP4DbgE4jtMrw+bM/LIECDa
iAK64adpGQi4wCHQ2+tzQsyBuBsy6eMmgrcoUDBTMTBJ/LuWkPuWzWMf0zztbm2W
u+aRpwt0jd+b8jnyLEQidr77Uf8hw+MmASxoOAiJdseyEupC05RDpzOOI6lzX0te
Kxxue7JUq/MoizpBTpZSjTmXliNicof2p5JSLLo5mpCWWKQV2rlKUY/ezdnnquPs
DLr7hbNgUxNWifkULXb5OMuu6zWra5KbkPwtvOcHmJpKvgtJTxQ6DvAti0A67dFg
FW1aCRXqzf9VSmZsFqtZFjPNJGrpRIt2p+OfNnztJRL0SGhIhAWIT8VKwAh1wPSe
C1Jy2bkoEwGiXk14MU/9ld/5vqKz4hj49+jgcWcK7k9efaQFJJ1n99SiDxLQOQ/v
qJMlT82G1V6R0roGFZQHYXxaodjgtXmVZvxDCf5ieI7ssyV5PNnwuWan6vUCXzov
JKWzpgkCAPQUKQw5pg1XgzQlNeKGjXrVDgNl/gSy1ZA7ZTJnFXh5LvcRxJBQCi7f
/oODfEJO/Jd6YziwVXgJx6dtNiUfm+t7oaZmVmpYBWysIXLhqHuLYEoj1I3Jvd9z
VPj2LqvSbqbiHC4CoHNOG36+DZFZ5b2tBbgvAQ57kL2Az1e96qtnXtPghrgeIXP3
ho26mFUwHoY9mjK6gwIzWAKISPbjzgcNG94zCCvPAa2hiOxNzVAYyFjXitIriCaL
+/cWOxrn+UlbViYJywGMO0EKHXho+j/s6AcGE+egL7E7Az12ZrafKpALboQU5xbl
GylUoc7UsOqQxNiXYoAnT3VC4ennii4VSw3SmsnXAvUkvvenf1hB4SUqJ+bMQ2tB
gZfyZfyVTL9hzN0dw1UhrDKZvDDu9QAaNe0r5OzL42PFJeDh8LeqxKUbnWkYAsrj
zrFSd1LH1nm5dYZYt+U8zfHeTSSrDxZ/n8PbSTGggg/jH7hn1ua452ddSbKRp9GC
9xYF+Pi1GfMyclqAQxAJvk8cgSEbRc6GK/rh4I2pZa47FyEwCvgz58hxtr0q7KJs
5B3/NtC0pIwinxK5VVtLP1J08fIntUsD+Qu6NCgMcTyYTy3B/ttQGXLqK4aGvM4U
ZKNjT8rAK6iaOq7/YUqi2MQUBN2APVap2IIdLD0FIjYHo0Oo6HhrJkeIE64Q4hnY
AnZK4tgv5Ay768CaSTaCqrNKHQiLWxzV8TubJcgmsdCb/Art+w8dmGdZs3iwPzjZ
D7a2muMNj0LEVI/TCKORm12MnOkjPr9q27IPY4rHxf/GpWILeD8YfvT6XajQElfP
mwBRX3XmF1mfA92ZMMOqNr2sgKDALyB2xVehqYDI6snoJRiZt6nmgUiOQShwyfeF
8U2/Sks2q7LDTSAmlSsc9wnm9Mkv9z7ACjIl5T5A7jQDYX5/MyDBEcQ8KfpfjDrT
Yibc6pKEVb+cIzaTEVJP+8224l2kNbpfkfqutePNDCS4xQ6A5sqS1u9hwAkUPij3
zurmmpwQDU5qmsSzuTJ5whbqPR4PbwdsX0XwY9vrSiAPS2AsZlrWY3e2ow4LnYHd
4vVxqAscvDLxpAt0JX158nFUugYpBjJc/CmwSOWAs+30LdyslT5yOFY+d4uZHo2X
lslPaSciiA6bie6L1kE0G0WlP7zPhEzZrEGRg03LfXEVjXtUIt4oUUlIZoGo96kq
Ssrl9Hb6Emy5ICQ3ElZ4K+/z2OF9MPLYanHnF1fTT0KcXPG1t5EfclkTDYYsmNjl
ZGBrH/Er/gyOprUZ4Q4ZwGcyMe4mzZpGBfkDf+EXx1trtw6O0t0Mf2YkLyZTQdMf
n04w41mSCImuvo6bNcL32rIkovyKtVJfGggdXW+1mtyd08jA5nQD9giCkf6qAl3S
5H/hP5ZJpHhIt+pmtOEhZwUtjhQ4Ijv0K5eKNujNZY/t1zjGYga8A/DKQaDd4lqe
cO38R0r9TUg5o1Gi7MTdod+7b3cy6H9wYMuPXhVH7Kam8eBQAsLZH1S6IHIMQFpn
sPEtV9CtAZcPcRWgArD5x/X0rZAsYcQ206BJFD+s169VviFUlU7BeZKMGAKFnm8/
HA6+QnEp08JgaYm15qN+Bc4DG5MxPUHdJH2cElPrPuaKwgbpFSRH7Foj9tq+30IL
8op+dWkI9Tg/Nc8liQsI60qQz7NYgVwUGAG0wf3+2oAVwRhcQXA7Q0c0iyfcvT9k
2x3qcz7H1qbSjD5mydajXPvb3SYQCYsl+FAuFEKYmsTWYEifF8KPdj4CltT+6Imq
uT3xYOox83OAJrAH9ZZhqV++1JpoQvuOzxrxAANCU0RtBra4iqqhvepyJZ26XXt4
g6XcdUFbPNL/pHBYSUNjDLDrmtPSLPurbj4kRMiKe71kSaxBs6dglfOjfOGT1qRS
Sn7/4Rlwg3LhHU2WmnEbmX6x8w8gYHRpmxPR/Vil9k/MgzHdJ+Q2PpJw3vlrJxni
FTIZOCF9gLPxCH7xYL0O6hrv4ToQw2NLM6tUwbqQjMBYaNrmRnQNkcaQvJuCZ+7m
9tFCxBkjMQ9KHJpY3NrojFSM0eF834qSS0f6hTPO+1UDCQpqdNJNbC5UKs59p3gU
h4qQrBNkhbhcrP22JJaaK1fgEAdVRrOlAjWik/Zn8i7qcoZsJ/2M5zWPwWmEpDPw
3Oi+9IaewyqhGjfVMNwp9LKWDwJ3aGtWkJrFos/9AcTVYIIyq+v8YEFhMCb6nHVk
JDPGo7PdjxlbgM/Dw5RSGvQDfkI5A+V5lbf2qjmy4RHOoRtpLfYdzK8T549oZ3cv
EAqsccv8KA0VYANf4c/wOSzNTPxEbj0zjVzSoSIBdP9HW3mzk41M10K2wRYPHRBz
fnI4q6GQReKibTSC1kDVNYY8IFlcdI0RUnbeqGLci0dqQxNmCFYjnQh3M0Les2No
V3IlHFDSrHvnlSM0Gahg3w7QBRlyYlsEo5dpZbDOVTljCFNKwrG7NylYfpJXahXo
7uMbK88xWwQy4Uw5pf064EgTEcaRdg2N0J+3PK/ghD397LFfsd1OAqMmhr+ixlJF
psApjY8g5aHdciXVRuEoWTdODAjRMRoYURlHBfvJveqkI8qZRaPSPd92YPdY1zMR
qiwm6PBitwtF1DDzuXtMCoLza8SI49zYL1FaKMba/oy1lS6dktw919RYuMXsCIyI
33bw15QhtEMUZ/EWQs/QWqRkr2BHa7Beino3zXrhuUG0vp6v1v2qXUY6sCN63uqF
P5Aqllwl1U3SVKA3cOd4D9X3JMPOIAHib08XHApNrQp1vh+Jsol1iVZZ4AUn9POh
hORFoW9ydocwizGjvfNUs8F9mrbr5LX9q89hX1VdpfcDEqwuaSilXmDt+KpVvLpl
bwWwzLj7Se+22amArQNJH8tmvifdLlrtZMJejWzgs8pffS+76o4bVtpjEgBsTAYi
y+p7vn4OP7l8katF1O5eNyKQMSFgblpyWLxB6Qq/NHQhVEQyYoZYBSboDh7UqCBh
eN3D5A0xNa4O45+KK5bQr1bE3YloMXqOt34s4t/Efw5/V6SA9Mj4v+NyJANaL2tI
7FZHVcMq8AffkuemtK+prNl9288l++owRm7+fztrPBkngg0jgzHkIs0ihlQtw5ZR
H7UTHIv1HJoGc3Dp2tRhKmjdOit5ndgGrecMuvUvlCe5B0bCFSLiUYnEFVFB8llL
MX4Qa7u57I3jMtasWl3EsUT5djp8df3T62ol+iYAOUluzAAV6NI9hf6Q8NgC1LAu
FT6+FlEroURp0fnJF20S/xHXLLR5DPnJsaDQG6feMtMJQt88LIduyLP3FiijWd0F
IndhETLXIOYAKO+OaeXT9wkKDghv1qWAo4oX5MlSon4Z7AtHVhLnIhCGnV5E8Kps
3+FokXn7at8bG4PBpXdEqErjQtFKLuP5BmTA79oyKLb0SdQW6Wr55tAwyWRI3j7G
wdbsB2fRyJu8hkHnbw1K6P2dr/ubtGtxk83YEs3CvnBNzKwNgp2+qJy0MyYmNQa0
5RuHMLewF2/gom4sJt72+VmcoDtqNd7C+ONpfflz8o6SbAw1kWy2wprFdUdUu4CD
XRb9f5WLF6ZlNNpI4VBt+yMlILSG4+vNzGpse2Nia0/dy2n5WMwj2CbJkwm8OmjM
RRvFkD8zWM54Gf46LI1JhVrB6XjOMEosuO50wM26zyYbqLH799uw56grr2Z4lZDS
LC8RYgjeu+dTymRZxwGB1z5IV0IBNzzeAYKiqKJKCkecMl/dvGGfxOJsXXTnY2rU
G7Gn92owedDdNmk2Z+Y+3BL6RdCryfCornwUgFobcoEwWK2xW3ZmFgrrw00C4A1Q
Pl2MqH2ogR+nA78E5xEthVBG6GdnI5NS1RwSz1Y3rz3QDIhmE7C05aHcz2UbE8vZ
5vvyVjO5zDGSBFMeFVUDa4YDW2eZFXQvFSjsPguw+PlJ4R48YL4AJCGKs5261rNk
dVCQIuutVfD+yzzLVjVqVvdZjqw5hjPvaeHoFidRt9UkqX/NhXIdzJmZmSoC7MCc
bmvWIAlYBEuq0hC+p+H5daaE/4v4EMgUiQeDVO3gdbT2vynfnswTOUVdN3alBsVf
PA+wMK/X0w2jBKquLrK5+FM0V8bdXNrDg04fTUjMbZzRpJWIX0F7EnOr3t//sQaB
6KtJzFy+5/hrludDzAZG4v+3m4XdSM0GKCvOGvFG31GAOZedWA36yMtIqzsh1rlO
Z4pFj/EVrEjOr9HmuJVReEUAsN+U+4YR4G0X/eILxCeNF/HUH/rJf6RbocmUaqvi
qK/wRMb3Kprob4FNrt4HTtvxFDeLl1Mbe1sVK+6vwK7kk7LVHZaAUDbw7tj/D9Mj
BV6InGu9uxypZXLWVNaltNsfwMNNJAbhIq08F2e4I2aU9PUI70S3PwXsL7jQpqVj
kkx80/s4Z31d1hovgzOH3RqVmYovpATcNB5/3JaxBvcRyBBuzHeqr9RXHotKy8VP
F7QbpdeJ8PgNomH0ryLGeMoujSTbTQE2V12+v4OuiAeHQuqciRnORjfLU/6b09sr
+FHkHuW6HZrJxNmzPjUMyHsp2+bp87LD8uMQWxPBZJx3yV5a47cXBOvTHLIevz0+
OZfBvZkScyAgQBJFt5W2vzQbHs5azikZaIlVSLGKmEDSJ7MdAVzubXjSRR31cIWe
0TbUeTtf4IJkee+sxVMg0vNbz4GBVIyflnvd7uRrmtECZOp4Q36AfHkKBCg6oULS
DGFjEIU6HG3z9tLyjouSaGiv1VI6hHlqQhXja783k7dwuWLyo5obOA6KNpnZc8io
LMaWUjMoBJXXgconlU4ptOWmATZflWXb93nErdMKPWUsQlRUHARtCSLJou5BdgEu
+qrkWwaTdYSVgE+K9hhlAmMOSUkR4lUIck1ZDoOpa4+oWr4jyD+xyatZz3sfckEG
vWvozDoTAHRqzLnJvfHNpiQfepnn/3VFKhLqq98dWEVQu9dQmldqTGpnkDIdOJIX
0UcHJo6aaMhThJ9ZdhBGHcN9rwb7qgImM9uwSxFtibgXaoxisbNjyfZ8qv35WJHL
ZUOLkheIjaVbc6Fb8jrhR36Wld4Qw+aPr8JViCZ320DbvXABYm7ZHHQ0JLM5F6sa
d2TzbqZ9ft3HPHV6/QslYXhV3yh7EiYfQ3J+z6qMHL7GZJh9cKmliBBhD8CpUy2F
AccugIR9Fkj/g6XmSuysGliJGRcyxWyYPQDKCTzIIJ4jw66XoR7qsveG8k/9AzJN
MWq14/FGZqh4vHu3Yv2sQmGdAs4BsCAjw2BK6zjgPU0c0wKfoIw88i6bsMvkVyRE
uBJtAnsxo65Ldf+Od342LZUusLbC12bAsAloBiiV/xGF/+GnzsIcYwU5rgDlI7Ex
g0CmQYl8RcLhZtaR113+GmaAN2c1pUu40+vcRCMb5De/0EA3wmtlyEfyFQ11fKDi
fDfQ6ZXkiBQPrM4MtkJ5KDAu0UfiUhl0hc6UchsToRW9udbvy6/0RPWp3P4rdZoj
6BJ0OiIMxHwHNO2xXeEqb5ovDgDQV1/K6uUBaWGiwrtKLGkSsEdOOwyIGgRspVv+
yXFdOrSHGKyup3dT65JBWDWYPk4++XCq+ZS7CHWaxEg89Lb2DxArY6p2KKzPIk1W
h2F8tGKYUDWS563G3EAuR/hIaYN/UG4fTdhugmvHH5MezHZM/KgjAGD8Gq5s5Nv/
C9mR7tnzFtArLLWVRUl8kPk3UTQYgDEKV7n0XNLHSX4aqa9hHKbJvz6V8IWgub7+
nqsxuRCRqb77ctWCIEfjc7OnLVzxUEGwKmrIySHRIQVbCvfk0cqlXKWT1QmrYMbQ
MijYBBRmudkPS6cqrG13uRJOrGFkCYa8aAohYu33ltsxGQ5kALJqTm6QvstpWBJh
Z2rPnzRNyX2zsN9tCuOQqqjxb4OVxEukfOFtpgV8D9kBAMbT72i3I3sZz5Fx65Nv
KOFVLVCUBLXmVBLKhzXnPTc7slh5X8ZQGXiY30TH5uhZ38bd4twr25jmXatB0QdN
8/FL/PB9ggZdvZGcFsf3yJXs0eW9aZ+A3ng1txZeENyzgYkbxD1Cy+P9+ht1o3yU
yiS78Z5Q+geUW94Dl/mvxpnWWOkknLMFzH2ZqcUmm7Go7bdGC83VD6g08Fn3Lsc5
HMNYZgMRQ/o3I0nr3UvZxe6M/zz5hQ3BjZtHC1a/iYaEzR+YvQl3uLYyW/Rcrnpw
NHEtf1ymb2NBHAAXVFm8S8/lQre8mugpTFJj3YAe85U+oY0a4umc+gcbl2mysZtL
QHgvd/z316jXOWVQmrt+D65lZexg39BUDBP9wxWi8IWLzF8KKBcv9634Ta4nHKqZ
pHtX2/w3ys1QGmFdre9RhK4NLgoEZPPkve4rt3kBx19siSh8je/VIW+y3YjKQmAQ
1C2hGNOA6jrZOB1zj+YznwL7A2FFEPtJX2R5WPMrLi8GB2F0gQX6IV/L7ynMBpy4
zj2mLx5N/78c8qTd7phd/ryv4zmG36YM9QPrElA+BAy6CQYwlnw2kK8cdYzzdu3T
QaMRehjuj6T0/drc8musSfdkih8/V74uszaK5gip+n5sqCYF60IxDPGZe4h8hhyS
82ufU4LEBGyWzLy50v/AGwJu7FiNARkmj9RVRIr6oadipvKf4VBWAa8gmDKyGjZv
FGuBYBTHxRyGUtnM0ItwBJIozOzrQls6b0k8ya++2uJzsQThJKmI/wNTx8b+kn/T
O4Oy6ZiedJN4/Cyvx1/0+cYMiIY8aruS4O3Sb+iun5k3glE/7kLnYkpKQVxgN/dg
smx6wBMp4X3KSqkCF2EkZZSj4XqdOteR3kwacAubqOYmsMZuAU4AgCxZJYLzo4Fh
UE991RXLq2fXADp+7b26jIfuMBl1TPBKYhQLocanFN+2R9Ol7PPG/5f2RuKXPiCn
dYU9BYYg5P8ZaDT7Yov7g6B8x5Cnz5lLl95Djl+JpADaXCu2j1MskPeL9QXINt0c
7Lot5IM+2mGhq+Ohf3MUvhJ0B3W15cA/WVfBLIVAZBIFRPHFZPsiVfGdLEcrqjUc
GlMXxJNzJsznRuhgY7Zgui8X411JHiTR1fyNQAa9eZN7zmB/upjMcY5FHHpjOm0b
5sPmhl2Qx7RLF8xliUHXt4gal3xBtm/18+SQ3900/tlb189CmUBAJe2yTeFiqyks
MpV5gzRoEqPb1yS3G2m18mn2B8ODb5VvNoyjsh2N4VkPS9Sjmc/gT0Sq9GmoeQRe
42nYLB7d2Hw10AEvUVre2rEUDABhaeaazPhrmUfI2H6iqct2RGQR4j/RLsTbcFZ4
CyXlp1Z0OZIGUJkMAFjLH6NnSwHZhUShZDKVPwU+wmHMRd8u0bY8a4fUumzHHwC9
r5ILFizizLOUdan8hcGGWdj0J0gGFkpEV9m4nATtwoKERscGWhT6fP1aImkNJrK+
gJEQohduIFGS1ZCEimSikO7pSE5NsYWSUGXH2BoZGFQqKL9IKv4ZsV6or7DprDFv
hSzMDwexhYeKa+KnqtGUZK+dniqbqV9T/wsmgHVHBqGoroEmelBp+IbvCQHlyR2O
QdXLVBuYsaOkh1riDGE6uzRPMGewQzUvAcFq+acSufGFuA2TWzbDgGiXoElXuFi9
AUWFHKDgWMZytmmxHfs/afWIW1dpoaV7Gg/s8qm4IaIVKbylJzkZPQ09chItAx1R
mbMCDuVf3zniVpohRZS/xrUXaq4xXbfK3EHm4imPNhAN+X1tgD22hfX9Z36edvoJ
cBXerhTUv3xtYzAqnVn7H3kQ79oJ/p5SOAAHa1B2A2F32Bt4y7yaHVCgJolT9lg6
zTRZxwQRb6Qkey1gkiX8Aobms1TyJ/QyqLYg/PFy8yCO023Xck8y3ULrh6xGnQcv
hE1pcljoGSD7f3ocROkei0J3POG/SvBW4eFqupHGs7ojtloh+lSe8uuaWR2M2vrD
qqAAqcr2TGv2eg6TMJ78sb3dZi/ow0XrG35dEL8aGdawYM1QhA1dyTueZgIVJW7v
B4SqfznF7HzPqoRZ7AyKwdKO58O5tbV15OQRuunPbbOaK6F9OUgrYH4B6IuymDqv
8VfQPON9v4xbQN4JoHOrc1DQXOnREbDSBFyw7HnAkGMMYr8VNrRycWOse1rNR65X
yk+KohINcxJIP4P5GCzWTM1rbOtVbqx3ofCGoqAyDhj7b40aQRs6lgmGp9l4Qzj9
c1merW0l/Ha7wJsL9KPhWfjOSX6zjTFjDZ/MH/kQyBZ6btLmlQzwa9FIn/PnPvlk
PFqRiokU1pWRraJ1o5X7tsJJ1UnE7HT58LUFOBtJFs+c5/66+qGjDRRZBebVePhp
qMdj9oNJZu/YqNhQ6BFTDcVXtpLeZYtjDlk4F3e5MFVvgWk4kAt33fe6vACxezkz
wFKZTblCR3G4JNM5LrxL81e0pF2K0iecz/z1wDXoxefBY0zNCQCEgCqrzfnonV5A
stmGk2K+vXdf2RJ51YvdO3Q7KH2pd2FMd6lnl7EtxBae8peC3n46xaxvRBY1pDmc
cidPsvAjAij4tswnqmOvua4xajk6zE4QCs2Ko2mRIEF+5DZT6K+CAQiH15SoMG6u
aeiw2JaMJklPopwnnkLGK+EAKhkguhGfhGTX7I6hAaSoBuTGmBtUE2g4NJsnwWZ3
1fggyP+ptKSXzFoKVjNgZU97z9abLCsU30scSiwxdTchEacmssw7tbzG3375In0S
JS6Esh5AWShbIIFcXmHn29CrHcJmH1XiY5owsEiJTqVHhF5KiT8J7lUnDTdsmWNs
3H92qCZElVCesV5lfFGEZKYj4NvgQLiu2Upao/hQBduYh3gkMbJEjjL05KwxZCrS
9d6IXdPERJXEeBHg+x1e3bxvbkAuBe1NBgsutCLBnOTSzkyAr+IBEWpu0jefb5p2
FHzp8Yaq5xetg881eVpM8rXWiMOWGgOM00q+fq9VVl+LISEXUWrXpA4I8fmfbFgx
3QmMZmXqFURSmyp+4pDznw0ivcHOK1HDIdJwMLY/f7unn0vypG8mIzChHokyrbAX
jFATHR3hOhmNjOmT/tbVA0onQhrFXT2umy6phFkYErQXXlP6eL5aFmrwRxeGmgxI
JdIb/nCdjr5Jn4jw5o6v10hUBM1TGOpEdpbDJ4tVclDtOwMFUAHABStHSKPOYKUE
h2TJYNeEGwq2rSkVtZW2WALZlb38Fc8qrzAgj9s2cv0AIc0UshGiPOwj1FN6fiJI
Ta57DhAgQAJALpcKB3vNE/mCXMdvOT2mUNzayF59tyIUoXJCvP+uJABat9v2z3Hk
Wph2/5AtqrCuGpp42kODY9rWGpERI2E9+yA6itHRS3wgXkZs84k6ZMuQUqhIahxK
NWUXmFU8XOmK32dIJtT0Hf8VsA0gicNm6JUEnZzQ2DkAo/Y8MMsqi4WOLiqtWuIs
x5WKIyL6WYZ/DvZq3EgDsNFeq1TLX8vcOgtT4YWoyAm544P/aWEy8+MziNTgFzr/
Lb1hokbkaI9L7k42ak8PNBitlntE0NBf7N3dMf+I7DFdxnK74FnPZXjGmG37/B/o
QS+FFfGeexSluv+EDxzmyxrHtE+eVwScDlQs7TGaYlWcsG7K1/BmEwwLwnv18hAJ
HB1fFP2ZPZ7hBiKBvC2cH0La583HsbvUvX4eAvUgZvNWAYKQ0bdNoikAUnwWvbh5
la3JEoEjNQyWaeVYc8//w9qiZsxnFq35gl3PZqaCkO8F0sXFigOyHSk8aSTZ/us3
565VuV54CHZGHIw06kBGjF4jK4HXkSmcM/lu5tY+Cr9ilIJ7bCiKV9BdhoWsRiP/
u1bGmXcVx8dJrKoHA3sZdvjohipLHcjUPXXyFqtqUXxAWioVDzU2HHpQcbaYiAKj
slaAGjb28VqrTQnZ4d071V9ODhYvDPeq4x8ovQ8NPb7z+hBHIMTZvrcuFr1664mF
IRNvYLa9OpBPU80TmPX0ngDnAJz+1I/iS2EDRagDyi84xF20KY1mzz8BqyjeFgFP
9sSfM1v1p3AELKc5JoD8uXsRscV5IpeNHHY0+SPp0WTDp/I/R/ftthUdey2rD3Ql
CuICivx5i4p8d8bOULLwIVx2Q7Hm4XkVZ8iEmGdIt4UHgMClARa6qdLgKcFXGTFL
ohPKk5TPoB2yRrwStwngUTb3h7VQgjAzJ17CH3OTFMKnHiuwap2GEXzkFOULwgGm
w08Mh3p2KA5WMh4GuOmyKK9jUzRXp4a9dk0YgadhYt8+6+y/QO2F+FDkLg3XG9Bf
ZfZW4RgoC7DKuMbsxVwndOksiLAqZw8adtDcr8bKuq0b2Iy/1ZiDKwbWJLRVTsSH
Vka+OkxskhIEQiFwMZE+HR6u4V+lDeFxtGHsUCE0+7VrSdSo+grIhvmVK+SOKqVU
RLYM4V/rkHUdCA7OZ0QzTDMJmc7Kw9l7WaOC9SkF1x9Udct1tGQmckAYx5KZfaTB
y8FC2O0/k+ORmO7UDOt5o/HgyJkdAWapNZ+qRyqKx5iIA+/wAFOC536kOqJM5Ger
oPARl7aQ0GGKXKwDWJ+55E2EBrjt6PFXPdk3/btplrAvRIFnNL35N0TKCl38+Zpz
VdU+Lks9qITNpGXp40Hz+yhS8kvXMkE/EVQGhpkhUfaIBOlCm8FnLfQ/GkTmCIZu
n69UqoBG7WPtYy4g0DbYIWXvPehWEWCDJ4+3ONtGJvOQ9fZDKQGGHvkf5erySc/b
YlZkIdxdVLbRi5pxkRra7Jb5s1VmbClmtjAziTzcnv1c98hbX81SJFkqaBGDXNQQ
3MFlaUbp5b70iaN+dhItrhHZ/KX2IrEHxqh1gXEL1ST3XlXhvgvKLscPA4sxgfZr
spLF4v5/d5LcTx5A81ZFXDMzI2Au9GZ234RZZQzU7kf4TUyzn4UABUrQwCctWlFK
iZheep8QrGSd22GyjGMFaTicnE3uotd6DJL8r73zDFh2Smj8+a4lIk9ld4/kab2/
cSvPlV0aDkPrbkMzwdl+ELXULKqE5Zux7rvPhzTIMb+cx5FtuECgbgTBiDL9Ci06
1kMnRezhjld0j6jAeJRc/yqa1QNpZrAOdFKiSq/s85xvSwiD8t3OUaAssguoLsKl
XuQvqiRRnir1afmITSIq2sLiTktebA9MEqKBw9Egfu3DuCgT5TT/8qVQT7FCKl0N
4ixXUETJTP11yvMm2rTUdxSBYwPrY0N7rQXbx95e2FgBGt6li9ZaDhTQ4DRvoJJA
mb6bH7dUCkN+xJS1hdrqNMqXzfBWOT5tIdrB+Ir9i9B4Sk6YH+YUAOjU5flS+x0c
wNKIZ4NWIQ/7fLjGAoC8W+kI6vvmuvKlZ0EHyyUfPxcd1FzV+j+mcQpeKHGvjzgm
brZ7y42dSKskV9uVDyFS5O5/VD8sbVi0inDaryKQAciZGRq3ZveL2NnOGvKzy1nX
pvWxAsxhTQ7gcEn3m/8aSARXhu6jtB9FMQ9H595iqYadty2j+8mGCwDfHXrMcCso
ARmBy1uS5Xd6Rszzu95QQbmIhPeOlkbcdoKibRdwgTKR6i2lI6czaVSMTOop+vM4
J/5HAEl9YL5+nvV7h8NpsJjkPYpim24znpMn63ic6fOgaGMB7CnVc65GWHkIgQTr
+rvgzqqjl6gNLSQP33c0LZC4CHY0H8CDG3OruwvPD4Lq3csZ5hPM+HbgTJNZs36i
e1f20IFo9CvcAWyhWHZX+wYBldz40wOVnYP0h5PKaLVTES2Fu9nAZl9JUs3BFbmF
1LhJP3gZgMG1vXVFInP0zyKGoECXlRszyvG85Oefci+WSKiSqF52gEpqPZQNSbDp
N3XWWjEtb3KfXnUKHuSaKdYSKG8sqGPW5ObUxWEpWkpKYlT5GcyMF8azTYaiV2e2
MGf7UyFhzW2Z9fZnbNRUwJNlZ7p+xZOiLGoPBwdKysUjvVn5EkzgYid7B/3VaiKu
8V4UYZk/YeGsM3Oyck/ti/grzvgsEqoNcgO5aCY9lwSFJf9HdT39HBjSFFKb3uv+
G8CoNUIIhydhWrJs8MCyBqBAkinOOq8RfKZNhxGdMYb7ecBixqQhq5hwFbB3QoQo
i9/IfvPiGeOBKnR/2JxpGtg1u8UVz41GP5cJA29j+mdZoq+Ff4+d/b442XKMxvH6
VASoCwodO00xRHN4RjESGOEXVDyyqUE21kJxchfpNN6sxpZMRBbaXiFDl7BnkWHQ
3sDwF3H8Uf0aNiFwQuxLLb4z5/1G2b34i8U7umZM15EfF8K7XS63r9+jasRRySOt
S3lPzJxrJRGizGmld8zHGa2vgLqHKDFPC1iWBHVizUgJxXDiECSqTC7URjNIU+YT
QE7XFdXC3PykJ08j330Kn3ckUVNAVGTG93BSA+7GSnm0n42BUw2gg0n7iZJ4mgdX
UgTtwZP2eRvHaVksrhSRLAyIX9pdKLs/Vr9lWT4Y0WMq0fHjNfHmsVbkKO1Rst4b
0/NkNaHO3EBuuUpW0XEy8mVIjCSA5abGI/AT4E7ujHLr7zuVlYB2ubyNqp9CnTqn
WkiVBhVqaIv8KD/hBCVbj2X/K/MphMlf1RamsKa5EOTMrI3snmFQcQSn1c2H4vnO
W+bIE69TX8Fj2QqZJcyA2ufCwwLNFgaOETpAZ6oRgHMKy5B2li0aG7wYFiXi7/Cd
6ApkpYZcRLGqG7oiBwhbzoOI7KYNnPYleY2UjLjJMLZ3YDOtr3BFeQQRM8/xGUwh
E8es+Q/8efwJHT9jk+Sa2wgUIKY7IWuU+vGxw3/Iolpege8cc0e2GZ1NY4t0eOmy
7RqA6NejRAjFeA9Zcq3xRuCn/d0YHY7mst6ia3nTTKu8Fq9rlNb7HP7j/CCnYqdJ
bAtUPfDFeNEl3drfTsKO2vPI3PifxPmtPt0olfZvnr5bMOwrigIbgGInBJxUjaDa
O/BhUd6YLazE8fMqfhJTb2OegpR5RHhY6cvP1NRPPi2nJFJdY1yvaiZPfRVV/55s
KeNw/wpnnv+TygMcBg7E1IjNJuLdbaMdSB0NWytf+H/rutABR4jge+hHQOxn61/G
IV+AMEvAukIKgenFVmD4xf73pcrNMLcbZPNR+MyhY6PwpZ+wiTwxBElsT8MHv7qj
Jq3wyz9KS2tP/Ay3Kej/FaKKYaNh9hR3ZODitifNLtDElOIv0tx+cpxhHfjZgX1w
iUffzwW1vrdWj2aejb2krq33MdTRHA22BHbAjPb8gqlTyNeoYz6ilAadyBENYmq4
4wzVr6GIm+rMbSqOZJJdDCtMgAyBbW3lgmTYKhShLyWkvU3wP9zetl/dZtxRHH3e
owDYkoOZXdm9MlImOre7v+2fNpXGWOoOAmeu+K/TJbla4peDnQ4g75oYGk0wkzDj
E71+LHHwVw/quijxa7i5l1Cvwc1h+r3Q3hDEXBN4QSEXd/kDG7hC+6dF480F3Kji
np8f22Lx9MXBHX6nw6NAldaSpjjMIqjFHArUqvQ4AOxG4ap6S6H4QudwytCg4isC
aTWHmqgBsqUBSwR3vCBhepA55WptEt1emhU6ZUl5FcfIGQnF1Zs9o/39AGMjsbaJ
3U6PCd2Zqf0dIYaz0RKFp4N+ASUwCbqojHzpNSppjm8NKBLD7k20BGlenFxeyMKv
0Yyfv1T9R3VD2nMCTst7HfK286/0SmtcK0/Tl6n0A6PPj+s4uK3VT0iEG9XJOGYd
miZCETLOpF7sxT+9kVeOYqqjItfi1elkPJJarga03uh1nkGgUrceNgagNmZoJZRA
EN/OA57lFUq7I+hN+uG7oYx3kLiCGj3UOsuoK4/qKGIMKPxF2Y70ffcveBxrbp87
/VYLaRPGPY2ta1MhcOsMJP6OJFzNGd1IZWopTjTwlaqEbR+i6ihHG7d5+Vwf0YVh
Oz/dz6OxjEzGKNiTgWgPH55EJCaMyIeJRfjbLMvRDhluAtmYS5Pr0i68Yv6cbfCn
nP69btFY1ODInDuuPwokIvUU5rM9wRlPRGCEE+lQoewDNhQ9l5RpyfaH4GvY44Ya
muYEu47xt3mezsSZgYTLpoS3YzJoFNMGgr9o3rhH7CINd5lhM3oj8//nrVs8oaNm
6lf4Mt/qZljDlTEryCAgPGdYgqaANpdF8jRlBK0E57V+boDmkw7rGd5HXB1fhAfW
7rMv0fHktUA7gxZogUX6GTx1qe/hXBoOM/SJJU9CFyojFfCHzSNWvV5RmZGISnTH
z7qAI/3v074UDMQUPghylbeSeBY1ClC3CODxap35hzQ5XZzGxwXwzoPSvwrFWwSA
0sJ2UcyLRU2ywLG3vVHP5N+xu5E1pGvr+HFu1b8fLzK5s9SZuu6zj/CyIcJH1udN
gnVD5t6uxAskFMqn+HKZjvIRRNruVBz12tzgRshUULrukL0Rvy2hGHTMiKFGXlUy
A4GZAvjSZmFWVlC6DfEDsCpg9DLJJoPvEBgA0CdUqRb2iQRLFEdkjJE9jAsQ9jLF
2vBqAAlh2qmwXifkyRRslgnllEr4BLm4QVMsv5csOALczHdGozTAUUXQnY1sTlgL
m5yUefp1y/v1OQKkt2UJkMNLEyVWxlwM3VjctOv+ql8d1dBnu4SDDMOGLTb5X3ce
ggmiydWsY6n/QDWK/JK2/HaqGBVZPppYPWqcWS91ftPXMJS7EjaAN+vrtGnnlCz7
EFUGhFiII2XSzigUwfipGs0uJnmq4A5aYoDAQSUNIkVIgip1IgLN40bqCdPD2ON/
6V5VAiWfCoOa4CrSg6jdMbHDMZuyQV3ml6yZB7/BxpRBOw24t42P19fMCJmXC+pd
gAsiOipUDAkBHsLZvRRViqYHtQL5c0gKQAYMfrbhaNN1Z3gY85JUcjVWWXvMRrTW
1YBtiTAfRFHDAq4V2qg8+dFoYXBuygN276god3puFwc8VU6fkbSQmUTKjkVcwBnQ
MdWHeuIsbKhgMi/pMZwx/iKHhA5/gssRfMiPV0JvCvyYyANRL/big0RH2qwNW+8W
034iLr4wIFq/ssyHNeKLWK00EUFW8WToYbWTZ0MPue2A4QDiLeJdjgWl9vYds/Zd
cH4Uoc0/zv1dFxI3mAJ3RaCEmZbx2qYOraO35ACVDwIh/xW4KwlSfe+ygR4RRIW4
LIA4gj408Kv9Eh9QqpiyJmPHKDl7Ok08VPdv8XxezLHG2uYXDlq0x3JKUh6MMnx8
qFI7U/5itOv5bobNotiX8f3hnCnmbuypbK+mpVALoJjBu0v4kWP6nMzVS9Rv6VKP
Lb1x3M4a3Lsl41/R92QZWZE1N3Wg2yjQMSp/I/LR+aD26pfMG3OEndudBXAzs8Zi
fpkv/5MHYHKDSF9uCNi1vuiWFbk11nikrQrqR/w2uCc0q6tBsT4TGwK+exf5euC6
TiV43MM9wWm1Kl0LNf4rZvrSYjuNHFfMjmK4yCyW/j7KEdvuKHGiG3VdGH0d1L1/
+uvf7ZKVJZjPddr91nLv1wcYZ1KrnD78EY8hL1WDxqoY1hW24P4JKQCwHAzTjvcg
HtBGCFxfyMbJqBZR5X7/ZhOt6Ye6tA6jErmzOfkjKaZgdIo7ZE4DZwD0/T47V0pm
lJ+Rk5v1cspbwdljgqpLysYt8RgSmECZMZpFZhQM0HsVkZDC6gbNqJPeftdh+K58
SYsfN6tJyYyzIunlh65JDfArI3w3clEq8p+4w/TFavWHZuGmaTovQQUJSBWqDK7i
hLogSvS/CJkaWzVyfQNZU8CUYiqBHCxKKbLWiOg42bClvyNFW/CIxfRmMAW2ECSJ
sPnCeXvcTLG0I5oQ9C7+Cxn9y1WdVlEEa6dpdNs3Bu7Bqmzt7GYCpZOM+Da5JkdG
TZBDQYaJJLMmAPLly1qZkrNU+1AsFT+P3lTTpO2k47w33M/PABtXBTIfsXnf3W4i
S9aA0sMRLJqQIe72FOXe/RAO+DbkKPDXoijkTpNOkwDGlkJKRR3BSWvb+Wf0zspt
4Dyee00v9PqyMU2NytRE/oIbeBkJwzE+/lUU1N3y9XHWVLh/wXeXsRX8Ib3QtuzC
zl51Yq2E58TlOPKKHNcDLTs+ZE0XfxhzUHNumVkaUXBi9pDLTCVnVQWOFuIuU9nS
l+9RX7lLbU+eD4xbi9/rtsVOV8VmZF8kkE2zyrHFMZlfGjCwYM41NT4aRoRW2ah8
wzKrUB4j/UvD9OqR/A3h+c5jWDHoScDlUaBc0dcbtUvxXfOlPqsohPISKvO75WYJ
17LG+N3u8cBKvr081e2mMz/2Gm1HkAcuA3fAZ6FZFD4yF+yaF2nPFA75LitTnre5
h+pa93Wsy+xmj8S2uFh334Bnt2IJzrWBAOHPcgfaAr+ddh7mx+0woAYLFtv0v/v7
ru+1mOrDHCcJBy/eS7kt9Hk+cCb0v8l8b9WxcmOO2rjmbT35O86W/beFI6hTWCyz
kllnNN2RF9fu4cqR8uz1CH27M+84xrBrdrH0xKCiy9SR+kKSkPtPWeVLFNIn8my+
05Btr2uQkqtsx0VFOGnfaISz4CXf5EOrVQeUi67f2HsD7Xi0OHk9pf+vZjjJQzFL
SxmOcxzt2+yHHQRXAJUhem2aDDowLHQujbCRazbReTsX6WCTqxCueyP//tSxRNIo
T6doE9UuXR8z6qOBD64gS1RFJ6VgdCtJJMAidIdt0QvAFgDIrhq0dJQdNYbQ34Xm
RS/PsO3lKu/E16qfUfHQ3wsvhXBquzTC/OYn0B1Qq/DkWMcfygfBYxXqWHeTkAob
R3b5knQ52mX/7HhnVvJAiaMGZKLwEZUbTpCkTszkq/lj5U19mfk39z9SvmQjEI9Q
DI8hWGLxZXDiLNFfAtjoIUgesZCks7jOagjj77YLUiUqaS5U2nPBnpwV5WtToyvE
zrYuKFnpaRcR2tY4dmiuxDT4Ls+G/BBHyRocuZLNUGV5mBw6MSlkyYd1pAnoaM7g
JilCsWpZlU9AQeMPhYRI/scP3K7ujsZGPHjTDLhOEmnGV16ARQc5SbN+HET/Gb+l
6mLJx8HQzCFyUF52+EK+vU5+Ys/Y/gQJjLiqOdJyR3Eh77LqWCoummfc7BfvToO+
slfkspcfooNj6xURCZVzTEvuRYD40l3P7x5ADKK8Wj1gAwaf3EJa+Fz9mXEPs2LU
NysDc4Fb+09MmODWZNhWs5j2b0L/YKUnyFAOe4bryFarNkWZoiUUrYiMwonIDLEk
wduW1jVuMs7ytjraoY6WyQD2KRNg+Jd812NSuBxaMaOgvq+SxAnPhTBjDcogO2Xr
AcPZiyGAXHIYZ0QMr0GaGe8gN509euBVri8Y4aZf8Y/p9U0t/IUlEup74lq9M9Rr
2gjGnk8W/7jbyIH2EnqgTvj3Izj2omNtUGq3sRfswVvHYwH1dmwDbnzZc1Iwdq0K
/sFFbjQCm/uNFTF6gnv/w2k51RoB6Xz1wG6IKHc8WVV3XGZdZCpL9l1RkBeqVTag
8Pn47NAdfEB416Rq2GpxD7nEEuOFjLRuRRiFWa8QZXVdJ5VfsGybVqxZkM5FoaF7
o+llqPb77osJatg3GDoO7sgXehWo+xTyi11HPZSUguAdRRlhVEKs1QfOHBMjf52U
O6VrJuxkp3ljfY45sDZy6pEXkNhD35jD6P1tmbcJqS8Cs/l8FNhi5A3IZWN6YgSg
Pc/Qaf2/sGzuo7+ekKa18tGWI7cVOFZZvd0FgeduSJlmT+s2upO3lKZoIPB1AZdj
9C1p1fJgYmMD12bYu91beXh9ph4/jPFkx+WEYsRKqUmIzlyIm0zxMO2BLI+slNC0
FZmiBAnWJ3ImvLW55cSskIuZWGiyQd7kdy85bQZSalOKatM+WQNbqA4nC53KnOKT
Dzb+XB5TQ2Kf4uC0JFpLqc0PVN2pmITN+LtRv6lIeei8I2CJ5gVdC971h8+Mwf4t
zwOBryJraW2S1Itn0h+5AxTPAP63kyBJiqBkyHNCHSa9GbryzsIAZ6jVgjTdDBTl
ENup5FSMPm1lcyqOzOlWLg+gFkXiuz6DWm02PMOhMjZSXZAoLykhsrXrF9ymaNEA
mgj3iCgZtYhKi+yBE+VV/2PM4XYcdyvNd53OHzBtGM0nBf1lpA4Oxupo64cZ4eIR
a0ijOQEN2cRNUyKD2YxTjKFOqkEeDHs97KSCybBXPRNmBaiWAoK1Dp3YnG7nVdyB
BmMA//mtfocB7q2a7/CBdyU/2mVCdCtZ+TRzS9qWFevVU9m7lA+0Un8kBqJQ3Rc8
auJh8rp+jY5d30j9AF0pUKI7MV882GIcyYX9D6dkIUw6I68MGdc/cGdH0LnaOOPd
H7CQL+/uh7CXWT83WPJeNa4CIp8zJz2BrE/PmmVXW9UC1IxuxPoliQVv7lng1kjH
XWDoMt+mJSwZImuXRoV5UsuCI1RoKhnGZQ9Of+HmK8C/8KccEmNE0R3ZsWdH62zz
jRUhSBwL/5TGNm6Kcxk+eL8qJ8YEOJANPeAPBxM7vWPa/zdGQprbODvR94etaDxi
w1JSlBkvbr95eGm8jqRPe5sNeOFdNrcDFl8tb4bn/BFpvtefa4KlcNTDmKxNkbFM
4mdojr00qc5cBr0iJcfjOdn0Gcd8UHWU8QEF1bune3+WFcBzEPjpa1P2a9iQ8zWm
rMTNEguyIgJve2I7K/0YHDivd1ki9QZibuTJOocoVXHx5wiD0GAI8s1TPk+5ftKN
T74mm+zD9EL2ex8xryohJnQxrmaolo8ZQsQPs7bETHnFv7CTfOd+46NWOCIll5DA
RCw9TrOsMe42jt9vZiptsDtVDrtJD91jJe3ng7mInk6y9XnXmJFexgdRceLXHCv8
sCxM6o/4XQPGFZf8U3X+kjpjAwhpx5feehNq3Pkeg4C0KIF4i7PG9fAqDuPRDRfs
dmML7n9nEwbELje74FUMr/8qWr87dMWlvDuLrInkI75uroaTFCMn8CLpZ4+DhcNy
lUHVnMUe3tY3PJ4PVCMRGzI59Ei7jcRk36SR1YzMt80yAZJhwdJVPQ/o0KTf3DdD
XP0r4BwPZym0AWV2b29cRvWQwCbjCfbfYi5r6fh/duXcp1Tw066Vj0pPHvkv3LqM
JEVla4Vts3EdngZwJkqh3L+CmDXQXdXeMsEoSr49kZDUdCnpCMHrZAXvOV+eysll
cqKj4S6hG6+Q2zOQlSPt2Ve4eIcvvAqtboAQ4kbHkBZE4RN91HpbrW+aKUQaCv5B
8CjO1vAk/amhGNotDSA6k4fezhi5gJwhc1PsGZOZ7aq2vX1yvwaQkt0WmGiZRrEy
Mw5xpBbMQp1jKYV7wC98bAAXzg4iWhIoA5B18vmQ9CIxiG34pJAyKI04T5s79R1B
u84thC30kel+2jJgvzehVbMNcHHMss0HcPDk/AafgjbznZpj+lK/AEET6fe5I1+F
kJA+EOXGbJz+OrJXkrbWvDVx84XGTUgstDDisZdYaA96uSFW3UMI2vfS31NMI0PI
sd3vK35mSafckyrGoRdmxkudj5on1QTl0DDGkcinZ3zvB2XMPcHQyLIC1uoCnXuu
CkoHVTDsdklRQIjUNMztUJ+LG5NZj008u98NndGixEL4n/DbmUMVkesb/ci1HhgX
xGMiV7mnDo1SoAEVEdK8Q0xHPxFNP03ANBbrxPvnqC4w2IH9JO4cOgI47JVCPTp2
uID796oNtzyPzhfJ0hmkygYYEvxbdNFFpvtiXCBN3DPMqqkwkhAHts30eMUZKrI7
zTAA6qNIMBTIwEZ78jnuPbviQHy0rNf9GN/BuDVCobQf1eAwzftxR4GsQlrmkhSI
SIwqx9J0obGPt9/WkMXCaofPnLAAwzp96tVtqAEB/Zb/GfX6Yn6uzIwNKjk5q7RD
iM8W3h5Dyr+Djq1zvNdEeadhCt6OZtXYIQMgOUq160fgIgXCQtZC487V579JlPBh
XyjjD4gVzoPh5cfgGT0Z1YYIUuDJvedd19GyqMHxmLl93y6pncCAq0B6698JluJW
rzD/g/zVrZFOR85AOqmdk+7TnauOmvAWFWHNahFOe0MFgmYY1Qik5qZ3vbL2PZhD
W4hDR8ZiMdjCRuSMwTAtGAP0jxLD0vNUk+ZbR38GNhNdAFkcE11BXd1zFkCJkhqx
hukDwHTPDfic2gk2Ndxm3HyctNdxLP6BeEjV0UPolNayT2kK1PgorxvV4Xd6hoJe
8gVCA53hhe0AQKnH34rBfadOEDRSGAR6R7ZUCXlzJ0LJ27dR12yiFltYi8xLpwEi
J/MYXNty5k0z1epJRuJuj48rAk+w35zJxicTXm0eDqlPZgGxcz6QmBZvoVjVE8aK
FKuvMcBGpGPoBUQyHz1yZ72oZymYWGcsH73PyaCFY7r12CyyT2w21Og4nOTyRgwq
23dLYUK0fOrS/RstaGGNyywfUumTVzLFcGb6bNp5vrEa9vsRwT2ray2Uu3Om1KE4
wLWGlCIcJjioXdH40xpzdinfkad2YyUZoCcBX02dAJpZAluVz8/M0ukbfvoujKRM
fC1HkoGIrcNWMtkCMAvA3vDI144/tsq95okDqKjxooPw1YfXNjqQdkzn2jnYvzR9
CThcB0P7cOd53GLvRZql9P/bZ1PRn1uM1s0N65zibtxFGHrhIopqgE1Bnq6XSkmy
bBLjEw7A4Wi9GhzM0s83ZGGggrSXBbsAYKpmMr/2vg+RSDWcTXG7KnqH4/o4LjYa
J9VOWEBp8PkvtpM9W7YSzlfXKRqdFf0OERFibLUUuCzLqRJQudor1VNvNac6hFRH
sTE0crLU1XlvBrgD3Q+GvfY/2KeijAQ8twwKyiFav0oRyIoF72ucsiZVO99DA0Bt
O4l+aDgpHEJjIY/syAt8qs+E1dgULPa2kzAcU4nY8Ij8m3Amf6kci9L/dav6vAi9
I60zqWwUhQjuHUifG0Xs4WKod8FTdrkW+6YlsbUT2vAJ+AJuSIalxnJRl6uwOYDP
WmWwSMb6rV3sQFa2uLOOvAkjEYMt5fFPTHR2h/nDB5cpj8OywrNWG9oAvo47AaPO
7jUx1pJtrUEiVwccG6WJOoGEY/M8f6B4e+2imCCZPGupzqCI81z+EDwo1tZaJVB8
0bBoX0XX40NMulnVQR3J08kDUhP8GM0+zUCSgdGXYE4qMSmwN7GWycaDF6wqN1q2
SiyVSmFE/6dNoNfxn0y49Zq2WXmw8nm5Pq9LpzqTMEA1ok5VBp/VMwmC/Br6AfLU
rSip0bFZwCTPQnh/IWOE/2JVMXb1VJZPeEZuwJeqgLiTyTUz/5Fs0HpkwCrs65kv
sbZsFcU9t/p2WJm71g2eD5N0718APZcDN4dAk6QgWYCYrmXAkzchobVjo/fI1dEH
UFcx6OHmg/wVr6EW1vJx91QOX54ZPweWB8wq8Me5xDtR/XtGGb5cFKO5IvMZnRpR
ZSvf+fRuJ/o7qqsUCYaRXlpHPE5+4d/RQ6kwzq0z5DGMNxsz7kD9fnn6ZoLRa3Xs
55nZ+he14N7u+61omarcJe48GUkxsZt6ufSw30pJBHCxzhPlfry7nLPB2CXBP/Na
uNXFYaZFL0d3cPH+l+oRJjLFgAcEJH/TX39FSvRqMbIuOYHuRnCnukvhtHYupjNi
+pJzIlgBT+8+Dud9jVz5GErhJOOi/uDufdmY0MObA8QTFoV1S2NosREzPDDKOFvy
RU90mI1XrAJUImcLUzrDIOsblioyogXYGjtrnlEF3SJ1hcPwFWiISeQsLjmyrnzB
JIYTd0cxPinifYp4M5wmNg8JUeTujWqQ+IID0KNNAdEOBfpeoXCxIQ7hAQuV9607
bVyH7HQN8p9fskuu8fgZ1CjR6K3IPyiYAbh6rgayA9bCVzyn/HEOWXRBQjYEhwji
tjLrFeM0/zbR2OVzEWDV4yHuK97o3qxbz9bvJnJWnIfiwDQzGcq2uEejtcVl98wh
iXpfk42uzSaKRUVTED3Wodb533t75Lmorj3subcJTrWewypMkkfcvap0/7k6eo9j
j+d/9gapbM+dsr0a9ONz+m19sJhlL2iItCR3bDkppcXa3wH6Q5koYa4tZzRvF9gE
SAxWFj0bAmMuu/hs0t+oH8B9ep3Jxia+Jx9JGcqswUEkknolybM3uYPKgEh7PS8j
2TbgfXugj8soOL14swMPVgFsZqCfpAHfJqxHDbFUqiLeqZjJBgwZwe1e9Zik1jX4
+ehSMEhxyGy14eBeiTBwXhg55eN/QNS2QpTyCTnByTn6tP3mJHfhmRvmfLJtpmg4
nrfUyg+4iDq7/7cvBPbHDn21VEuQ+yXrP6cLNFcakFrdxkuGVQs85aDZKOthBQGk
T6hcX8LaIR3ybyAiOrDa7rovSAe5L0MY92VUa2xAlUFZqlnLzqzMaCDtmBSzX62e
ZuyNPfSa8/v2Hb7iRWPSDTAIVDuXbhQmlZv8r8l4doRNPzxLy9Rn/M1DoN6S6O7Y
qfzcVb1UJ1IrKdAGsPRgs0/Zekq5gS2UkbSas8GvPkWNAibnxsn37V5kuzgywbR8
TGbKKIcvVGEHCTMt8/jrl0V6rycyy2VBMtlOezmfNRv5eWWtvaIRJzlF6M4EiZLf
qXmr9baPKfK2VDQrIy3HiMvOhY5zVq3PMe1BNxU6yJgdnyBw+PN/wihwaYFyJnps
SlvrOw4xRyJ2IbXTWQMUlQPf/pcPh2il7H2C6/3L/AyF8MpJ7sQIT7Z98kE0OXcY
+zl4LL7PBPDENQTCQfN26mSaOQyuyThQcsF+7cUpr2iKCPb6TaWWx8ixBHQ6PW1a
NEqStha+xKrRkJ2Tz5IehzWblyB8g39CmMcebvV3ypU0eyTd+iztw1WG5GtAtTXG
5rANKwUwCGUiITDtLIIFyKv4pHNZJvNDhlslcQr8hbK0sWePz8qxpzOrtSnjvGMz
Cq4dt4Y9GOW8FWI35ocwmQDIG1965UD4RTf9YJdAa1NU9QhySRSq5ur7THW/Klt4
0icfrXBFrG6iDIhosDQJJcfZZY8fSH2tF54muVkB3S9DVPECJyl+8s+mRrBM8G85
nkSYAh72HXcwmL9Tm1anyPzeFN5i0vHmQydmM97x2KK1gDP2VawzJbpRPBoE3Rif
terI6SjZO7UFSDTGB+PuU33vF4ht+O40NOPtitIZj2VOzrMjSaPaZPLqMHMJisyb
Tk/ONUMzPGVEBrnICIK3y1O8V85M5eANlAAM0Qli/WfwmrYcBgiTulAEo40EBvw5
/d7Ra5Yt9fMphwkn5YW5BbN0vsfyBgdJcQUQXRi2yedxfYegWXaDwHgPxsh3sdKo
eaAmvy1NoEOnQF3MSR6NXb3xsF5peZIU16FB9yyps0rwqpLRK/b8esJncC+DXlDr
svl9Jrv4ttImPxuZquTrSscQz40F3Y6jCpmYWPiO5Z82kNmkVkAwJJUEYKEoj7Ha
aHnatcGpb65xE4IFciDOWnYCdlmIgU0hJFSMDwJBafmYGYj0yhB1ATr1NUC4+ozF
Z4W7ofnijvewgkb6QAAdDtlwHa3VcrR1SskuFrfuJtIBHcAtaY6M+cUy8lu05FOj
fkoG7ctP26pFVGcFda8CWXynQYFJI8QeYGoJk0hzrVa5af7aNhTkkhOxau2shsMK
2DoDVViShFDhXsscXrK3OFfYfWxSIvU232e34SKRB0MWQ146AOWEw4WKV5SP/o8H
So23DWzmyZJHRqyihfUN3eL8g4uGppBRRjr0YyySFgyIZjHgIs1KOsOWrcGf5Ng+
KgJXbwgffNFk9hlPof8oK7/9U1j1iNaEz8HLJ1owZXXlSNhJbQnkoQM3O2RvGmlL
B238m4KFEEgI+8YAglzE7KwFOYzBfLGaYsJmD3ZcTsR9x3lmShCdnJe1BOO/AqaA
+Bm6bt8dw6/AVVmVem7DbjCrZeflVKNddFlAS3GtOMK5qQj3DIoeA7Ez6inQyZD2
hbLOewclmFvXYIcMta0mJ1lsWpcvgNv+WL1hJHJGGklJC/FJzbINoMGjM7U6Mu8S
HghJm6xqXzSbXA7C8T59fQFl48GUIM2tFgh8o5Pb3JYF9t2xvP3rtjEIMcPSaQJp
15Is09zPCpodNBneUKrtzKA6f6Dzc0LpNZFWRTuTX26V0YPoQnG7SXVHYgHVkHJl
sxAHenlHvJH2M3y6TSJhzEpb8Nu1uYj4RT0LS9VXgTNOo0W80HayedOSQ+BwVWiG
P3TJxlihNeO0Tb+24td6MZAfe4kxHd2t/yu3YQnsijjBeA82Qtnk+suB99PpzFdX
AB+J4NfhnMA853CPR+osGAw5dXSwzeToJaGMUlg3uMFwkg1xgSC0nEh1j8sMBcYE
EHbD1tfvK59QN4JxIPLono8TK9G1wK0dWFd1tPXWNQND2fwTWV8GdisXHNBPHOta
wkV1GqBv39mlE9OcLEooaoP8zuefiI4i1eKmNjAmwAtF2EB5mCG2tdQUzZGMFnI2
apGSwbNfmhj76RvU19q4nI93CQlNoAU+Bqo+k5m+KMtdpQWwYbRRsnaTX9cFxRCH
GVR0093tZrYUZEC15459u0XVmiY+6oDkjnE1jCaofs24qKvOnPuWUFNHowVNFJ1l
9rkBcAQ1QM0Al5LV8yuhYT2vhzXDKcBR5I7T/CIFlNbZxwaECzwDKOsZe37dOFYB
NB11QF2KNAREITn2WzMd5j5aNWltqXbLa41KtbxLUNxZLD5vLAjoaVsnf2En2j6/
UiIh380CT5USefaX5jFwY/Kdw4awolkmw95lQfRYfdZA2OHbPTQC1u3hYZeEDqHl
5Ip1nW03JOCVWC4ZdHjpAYNmHscxUqfYG+eLs/Aa4p4iZl9XeQWvfkhPwmV3ZvdW
IdJb+pV3mVVMnQsSjwMif2YtcFHjdtZ+5t+jxiWIw9SoQcFCWu5M4O3ZBuhMQJEv
itsS4TQ/vULvdYq+ZJfhAB1rZovgk7ji4P6aXXz9dXGSNhCPazeXHxI4u2IT+Y0r
hoi7y+piDC5lgQLZgMLbRKdZZqle4CosfKxdvF5V+FujvtTF1HHATcn6IS4HtnSv
djG9Wa9lgMXOAg1E95dui/RdcopwgTFFsXDVIvWWnw+yoTO+LKr62YNmcgUz2Ksm
CHDNX1bENNeHfnQIBiK1W7y8YKV5qRlPnWtzwsLk4F+hKbU5gNUfr5zMio9h8QOs
qpwXuNWb6fZ5nnYZ4Yv0VQINgeS8IkTPGB18bi/3c4SaTO6LY89zvzQknyqwvE/Z
KgPYLAUPqsjbGd+IF4Ns/2VdM0Ngy3LGdckgilwJ6IeUFqKMNpaua23ToCbOKY3t
N2CtaNxzWFpfINI0+ccY3a59Aq3BbAyKbOMfexr2lid2zkCk3Q+K9K8Q1i/d33tx
otkkXHmfiIdvn4L6QtOH1wuZsGOSz1ycPprHT4xXyxuh9nleF78pHWGZH2XJ9E7G
LfjXOt8YnGY7WWPpn/vAN/XrwxmEWRayF4CIIxebaKJWXPP+gPiancLvMCkaZ3a7
Bkdz0PfHLwXSf5fa0ZGG8RAItbf80qKFyPeJv5U1fGdjzraiGMg5DNOHQJ6L4xOU
rJedCaNDAtbqrWJ51ON+/hsJJklnn99xZDEdsjdq8SBL5PQVUgrJ4hpdtbKjCYSp
BRbtCtfYtHJsKsaBwxN+eJqsTaNdHDPez78uJBMJVsZ8qu91HbusMose55UXkmlH
mpy6CcQAqdL7Q0QyOHeFIw+0fZyqgUGG6MpDY/hD/yku+AdeT1hfnUc6wueu9687
mWMMtw1QPxOASVjZ3XkSA5IYmokLZ+XeOk2n4UC0pj58HJa0RZJbNkPbPlhACV50
+iiOcjcJTxXFl9pakO4E14sWKOsE9MT6MtehdMPXbOmQdNyQ6SbRdlSp+rh+LoGT
vYmurPxU2E6agLQO/B1J7yQcRl/QPrPN3XwfKdYewIQLZPV5U+S2VAuPUE7YZSr6
ruN4fIbZYv+XUIisQxLw+z1agih9kGScfOBs1zgC6cdVFRmnaJnFfPi8RuncVgb5
8Ja6KWk4PggfiU/O/NVBwBfGpXPvh2q9bjFitGguvRADqZXqDncLNxrSwREJ2sAB
mZLjjyfUYAoTw3yM8qXxfIXdu4am8zlDtqT8ENMxMbHRqrZEjDk+qdsxPiU/2UcF
lQT06qp5jBVXX+DfjuRsBrJeVAgW87qIgq560LB0MoaLXNIKteXrarQTEWgI4xir
02ENezlDGgbD6RkOmDzOx15+kEQ9eEIYpiZF8NjIz8jACkTfn9CUs+/cJeaIDnz0
6PiqIS7kNJ6wcT2ckhDIIw3YV0oIio6LUtRZ+HVwwVOxMoPpiHDnwh/KICrT1BB0
Z/hETXLktg82Q9y5Wk03h24v7o2JKzNYWJLs+uYJy9I1kfUMMVdHsDfbIAFrAJj1
TABp5l5lKJE8VR9CKhl5uXC7CGwj4HDXfpJdJcBkRa9abwOmln0JYTQuUjXNmIVP
BBlGWm4mxeUAVsPFhsNVuNeq9cYUJM12kXGyByarD9Vq1S6Nk7UkB6En18sd0axK
i3UzfcO6VDnfktYQ22j/mu0+Kl4OW0U4h913YH23LlHxC2ZExqZWDP8NFIn0+8gn
5YRxmeN+KD7+/oVxFlWLT1zQwrv0LavHer27bPOQtDGOUPf+92QcJ1qFddtTBbHm
8g5AoRPjtP3kjckScOsCNOIkGIYAaDfXBcRHpl6M7kpYadyOweUcvO1X0G+8CtXu
1OyYADqBKd/4PvhYr9eFwyKTOld3atbbDE9NeuJPI/LaUno9MO13W5IVoNSslUhr
anF2ewdhl+maWcPDDvwwbiKvXvVgIssDXGlazk4XBe34ADrE2K5lvaGonHxJktE9
h56kWE89gI0rDbXuPsygLLwo9KXpYRYy2vjSWf0kaEcZTY+MOiqxJuIB2nn/rpKF
hkmJTnBFfMwwWKgejuAixyahYRZBebw59mF+lSarF/+64awrG9XuFmBUhOAm1BYv
cNXPdD9YZUqnssRcu3Koreb3EGjBeTBZh5Vm6PwEpPHEvWMIZhBcF6rhktr+579/
mLQ8fVdF00oWiQbVTKyGv7Us3m4EQE/jD4LCGlEXm4GRE9ZbZtI18YB8O7Kcd1sG
bO5sGEOe2R2C1Hn9LCoQ5FECDSWVdt7BhBs20xafMhIDctv3W40u9NIyttrZQkGN
LSxkvigawVXDyLW2bBMaL4/pKz46BcJ/XgB4P6t3FM8jk9D/pNItNG1phvaf+rlt
VCgeMNl7oXqTTXjVJiVHt3iAXAqaesoYvn5GLgo0kD6fh5PiEK3GSdIiGDSYAZvW
kv8kYs8Mfyf85rXZ9BcW9igmoror54ltKGcWTwBuuiRfVZtqZjcFtO8my+Hegm1Z
rGHuyA3xk9ZgpqamCxBjTFKn/Nqox2Lni5XgYzfLhzyKYdDw7UV2BrozFF7OM7Je
nD/rBR8+CjSZPp73f+wphCFIglb/X6GqFe4YqdvMIIPYP/bc9TP9LbYk+wm0iLp/
afsTIeti2nm++nSV/+qVK+x/kAYO19Jw/HC2elb1PWUL0CnejvBnI38c1hMJcNHh
971p7aF1Crj4tyvlsUOGvwiqANLeCW62jSKdom9PtLN+W+mtMoPGG/GWIIUw3Gvr
ierNMLbu4lCr/Oy+rGFG8uCZ5dDXiCrQE+hTTS70Mbs9zJtgM8MlFzZsEDe1HADp
A08w49NHKRFirn7HXIZM/yMFgyJOX6+gKggSwo35RxDLD7MJYRFtQL4ozPaZL/2y
4gboWYfbSVlOW//MrQS/z6/V9VqDVTVgYky0SIBXwDtuIGOaI7GjHOv9b511giXv
MTmC7gDpOIfS3Vx7QEEgTUw7SjlmLkQ7k7ObF6cy4rnfc4uBU8yk+qI4gxksFpQP
d2S8v1QixPQLC9rynSWBAKBFzGU9QPFFbTZuJr670S29ktkEcidSrKyzMhDC+Saj
thKWbieILRacovpEDr0r2IXmWSbqku+RxpNTrx1IjgzdXZxbr9Q/zOz7JR2DeExE
zWMazhKnDEVgbgam7FuizpJ+t4RDcEaexi/dUdNBdFVAE6JDbzVU2s2Q6R0p2xTt
8KiJNKdnXnqdlxdXi9wOqY9wCDppuvIMclTkMtJPsAwSeq61ayRnDys2TlEkskT+
mHFUzJdPs8tqzumM97nwUdeYaKqTQOeVVLl4+kLmkfUCIumEBpJBWNVbe/mxb4sU
YpkRV+SJrQT0gqTmpq73D2mXN2SAGA9Qc42SSztqRKuUMboyTjcHiI+oG4Zi0Zml
FT+o1K5IHyC/LPZE0rPWBva0SdR2EXGGg7RysJnxiMK/frOb402eOTAEVrmiyNKq
cl8D9IkYu3feQ2Gv0eqTr5kH7uy2O0SR4VnIkCGSzuAciVkl4raCmSy3IgENhTUJ
lDJX+ETrH2b6Q0BTUNB/wq1UbwaLFW5SfZr/54+ezTsKANSxS9WkFb6AuEv69d0J
5kIZ04RZmuMAe6BfN3TfdR8EZU8pGqoIGTRhpfDGCLkTqNBx0hr28My15l4TvJ87
Y/G9WLDOxFf3C2yEBD3IBh7KVBxgVHGTA7MFHtjP2GiLCzie7XdD7j3guk812/j9
OVUbfkKlHi1ECEcTeCkwXPK1PhHj17aOgpa8dpeShObLmZKGLlM0+SM/a4M1vr49
q1V/ZynP8YHqV2KH2crA7UJE3ojEd+isaVSLDFbK1O55T/JUW5ruc1xCRf2HVJB4
syjdznI2iaDg8EV2ugRGjSCq9QYDrH/JPeh4QprYC7DoFAGYwiRu8tsY8H0BPZp1
JrdPakgH9o+1+e7repUXbUHkjkb2CYW/UygPQIPaUIaCI/R20Hf3pPCt+aBCuk74
zZh8yc4TDNMwnij/GmqUTaEYCSSyP56S1IkfIpGzXkhK62IsFox9qo6cXmgb1V0U
P36YyFS2b6s1hIGlnKnN6SsJF4HH5JLJp7fA/NHixr9Ue87LZ3g1a9BXQKX22+mC
gekJ3BRX7Mg8lPUhEOhCppNzPcr4WytC4M+xS2MM4XUhTRy+whFiTTN+Ax38EQPd
D5jGBC9PXaex588hxYzVmswYacZmys8VihsS9KDB0liT/1Sl9Ce3m5gxohB0T2V/
LnLAjfrhSKUzbJ953YKf5GmitC5RdnG/s/Yn7F2F+1en5PO/gPmAn/iK8Ze/kMql
OsPcicIAtFJHRdEi8IHSHotIxzRpcpiUko/LeHEete9iK+WMneZVXhySFxowf+WH
ukRtnJ6jpyVsJFzAfK4QGzRDLpTpgm2uNz6wthISpeBqgdycmSKvLtv6V8FDN1VH
aKjA1awcHD9r1PIb6s54WuQNxTx6reSuGuAYEQiHA9NFJPTQxzYjcsNlZnKsmE8L
CMVQezOS/noG9G/d6n0sPf8nOzdPTGigKmW+/FeOpbyi+b/yfF/azjYOLiJHN/ok
251RCBmZgRwaPpaVHuTatwtbX4jRAItW8i/ShzxgE3qbZlG/gVA5QpMuj29Y4Cfm
qMLbNDA5afVjXiB80hDDWNM/9ruk/LaFcBeFp3T3La1WbZZZeOhoAjXdUV6JSRTM
Xawyt8pwPSydS/q/KYsO2w2KIKRjIuOP0bnwFN7foOni034ZCwSMhONiFAOsYCV+
FRa2/eqCCWjOMBwV2MckeZjaEH5mFRUMJ5LzSokrIT4KwW9piW6oio8o5n6hTKzH
0S46kLwLOD7WPOxdDLJQSs8+cKiHOlOccDCSJKkJsmV2TgMFhI1Ulz5cmAz25O+U
T8KZpRvs8X/wE7/USEblGFkQgMf3aAPTQVgnroee7DpC9Ky8DXSqq7sT9pVW9kD8
mXGdRrQyOm14OT1G8PF1tr5UeCfNrWj7EJ78Y1SQyvS+FdiCo/ISL326Vq6cR0Zv
RV0jpSD87OWQbrZeN1ehD0Ev1oV/twxj1/KDfWWQdPzpqMgDJTr0wZz3Qx62m2/A
bDPQ2uNdC6aUx329rIyoMrwSx9b/OaSqL8W3XVK96gsqcoyNIT+BJ5qLJUXBhIaP
A2AjvXyhGX5AvXACVABnouPk/YRBMaJunF7AbXqLJq5gcrWUTel4Ux5AkukKG/J1
imzZVRK3HnhwV6GNwcePsA/cxm7UZFF228kn51JTyy7NWnWcNolrgPzpH2ahz83L
9IkPqF9vYkE1iU+LGB425z9xw8fZTLJXHrq/bXKngSApy4bzRpf/8IhqDhoTyq6D
/218JR5Ol7CX1qZRdMOYi75jDZDkXlTpBaokapKk3p7r19RuKueCX0PG73WmrS3u
2nWZk81tSuRInp9FKbeYBqtCUCkYpw0EYcZKvqG+CnmQEuA2zh5hILMsYbipu07V
BVKSCqT2rKUwgpbzMutM+70YguyNrh6u0vSSG2LCb3Kd9Pix8WOZ8izAIfLJpycE
nBzK1GXxeerJkU5Kg553hv+mciCslsVEpq+Mczdlh7Q7HnC3iepKBAJaaDf2iozg
UQMcSUaLyp1TTwiXURPXqiB82l5wJc9G8ly2d6iz4h7mUpRJFQMzA9Cl4MaL4OEI
eG5ScNvPk5aodIRqY5AzY67mVSD7iHay8bLtqgS9ngjrHdgC7D/cIklNLOOIxM3c
NZjhv6v+WFx77Wu/Pfv4pvWuUOfoa1Gl+h2CTNWz3rTcK5yWRGWdtUnUO6E/Ssyn
jvGhC6gtcBIbQGN0mW5Ab9gPXxRapsKCAGJtxXxUXd9M8GLy1Vs15/g1efudHn71
EngQXal8WfzORbemaHnbLsprLyC54YKujmFW1GridCiEimnsZ9h11UxNHMZ3yt88
GyTzhN5yrWkLDmm9DdLgKRrGa1Q6OCuSGBQqirpO8rokhw5h5SXlt3oAkUeEiD0h
2RslLky3Ll8YCDH/47A5EaDLREO3hRRq08FtcnA0N6/3LmtlRky68uPAOA5Tjsia
oc4vOO7EXkbvFYitlIToO/lGHg5kF/Ji7DQsJ962ZJAiCCndv5+jbDh59GWonF/r
IjjPx9Rv0UFEHQC+00rxOOU2geG5x337fc7nFzU46vxb+h1BVTkW1girdps4WPJ2
tQf03JGRGzGqooGPEGXwsPfywe5E3Sh+Ni/DN24gcnU5lw2Fncb3B4a2oRmg3xm5
UxXmdZVXz8ZjegiYuQeQoWlruRcOBesngkwFs1fQ/k/pplcfDYUx3le6bcRAmRC7
V6qRsSv9Dan7+TXlBqyxbpOxFnQc8acj/KEHMqgZCy3pK2gI0m/ai4poIgBnZH2B
1deOJa1xz1xUe6R+R8SVDsyXjRpjlazq7UCSnX+WU63VAfCw/dZNTsuqAWVPt14m
IZ5bPfcvH+geUHL9ed0809ndvZCAreJ/nju/UtFqeUVqY0gomow7JplbEOnl+Hu8
0ElucJA7679yWNkayGnppxo6GB0pgomXjp0sul+AbJuz3akPJZG4E/LyQJphCUv/
ktphC3eymguUnM0arxMB+6JE2IjsPkR/DaahG0OPzCJy4xwEMGZj9bda+j6QCxRo
O4+VF6E+Jq/kqrWZoyDRiXsZ/9HYkTt0+V938JOzpZ6bBICJplPw2dYX+0sHQzxv
jV3jjRsMRrg8Yz9YoJSt9RaZ5eNtvAYnWiCq9fcQCSVZVUXsPBCElxZqAPB1KvY9
8gq7taBJNsy4/Zcc3tGTJcbT1cH/X/yFyVqHp5HoJYN/adIqxs57oeuGcKWXVkvC
7Fqv0phDPn+rId8m5tNs8pE7OTv+04Om1ADb4O8QCbf1agwMIDB/xbHpSg1w/YQK
EHz4ME7IyKnTgrdDFZuq0uFKqN6oSQGyrvsEEHW2VhkbqmJBtXagf0FtTlUg9DuG
5LCAIin9ega7iR6NzdRWWuwPaEFfJGckEip3scLtUtfHAVCcZV46lWo792ztfHlv
WvnpZd1AdD1NOcEysn87rjZCgGSuGv9t9LhO19fZSJMPVJaO87MXlhQKmkbx7HNs
H4vGpxby7ZktuzRr1ltrq/+IM05AoNmGvNmB7+A4Q9MteS7JeZcHUHIYWgo6kGOm
0F//zbdvsUmmGQJ1A3aLwViv110G1XOMS4kSrlksn2Wuntj4wE69JqdZbEI+0tC9
blMV+SD8gZtyvCcQwa5WPblXqjjpTNxzb0xgCyNb2ciCMhKBQJYQDwRr6ovpTVzW
8UZRZId534UjINiqngYgLs9JXPbvJ53wZEFvYsaThlPYNmkm2BqRlHtBzVJ49+E1
txqOVGnzbGU5n+/do8ln0sHZX9SKQMqSzpe/VhKfRTCvPnt1yUz7VtwLloemh2Vl
uhtnqhGpyvDjqG0GI3qw5iDmeQo6w1vjoSBgRAbtFRpoXj04GehfbjGd/9BUC9/Z
f6RvH/ln3m0ASE2Vq+dkJp+FJh1JWrIeb2I0IYEHphYT7aYi+K0RCMFZsCQsKIAg
do+nqWPyb1wh9pDd8DH+QL/moDbSYu13ImwgCnqraQPEWQAN5gc3ZdEOlziw/6aD
DgHQ8rCu7xhmhAtWXMQrxTE+Oku3noUDHJY1crMNVNH2llb9vjdeNIdXMSS+RCJ5
yNnKA058bzlLSOOeUSXryOAfYxHWiOsiY0L+5w37PKWnFYrRyM76xnpzLsge7P0G
f69O8ylDlkd39vvxXSy00dDiCRxPTTFpRJX7L1gtelAxmeSIgB4zPlI/LoMQTqW0
khhcISitd2k0+PYIpWnJUZ/CnA9ZLt1H1mU7xvwToxkAHJMVr6A2XbLcnjzbrmY5
GLBercqxfHw4lPQtkODXPXxlTFveK1jd8H4smkn9ldI+wf01lHPJdbJ4DRRBJv8C
d2lrIED9KSx2XEC9HwwmpkE2xuuzt4uLoAWqjtvSVsxHm6k0toYA29jCaxTJL1/6
fFyxon53REoGYpHlwJ4p9FFvXtcVRdHjunO+GLDDHCEKf045HEg4mpjQqQ6B5vPa
QacQxMqPHgZZSj6KWx2CLOZqRkDENwW9131WUvb4Mg9cRwZkq8/iO9plvP+z6HZ0
PY/kUGG7EV9oz9YPpYPazPQxB3ULIquSNUZ9bIzVaN5SG14OAdarFbVFutkVQPk5
72JWjtxw++QFys1yDq3oLgGaQtU9SeM2sxcBB1QVzD03LkXdwiH/wYK2XQD6/cK9
s0/XSfKQg5UyXAF+i+rx43iEZbPQViTSBOfQExNZTttvXW+UH7OLEms7z0FdoebD
sBOmFoRGzPiFhPzCsKpYsk+WgIDhl20lfrBIuP1yt/ZetCzPczsbtVFawht2RoBF
PDe8c26Vw3R9nY5ac3tOcL7MIqHKfCUlhnIMHPaY/PllWRXlnHh3r6TAspN00Gu6
/Qf5K6LNuyB3TVP4sxiQBdfxSyXn/BQ6OMIu8xmVNBP3pBbK/Boplm9s22kGVsQe
wz52M1kZISpQss91rCcuy9LLzEyDHxEzDQo0+nd8AR/3rxllGuloxhvytEG+E7Og
Z5xaMSN2yYW0+qpvXH8SLgQLM9LnjAXNXJG9NY4caqhsAluip2SUiOHuaNC1prtw
7ESf6IIMT9SMsgaPTTqtUOuNRVBUht+Fcm28NLdQUAdtv30ZLFfKmZSXjUdyv+Sg
1Qf6QaOwOxXNUxW4eUqdyaPATreoHTIbzF8Ha7D3JiAnJVFJCmSCrHkAQHbO0JMZ
KFpUOinLiyNOUqg1AXifFSLjU11an8aHPw6Kf61qHhfcajzQS7dj0O4bqdnKdOBA
QdiUpCNA/fPxTGNZzk/c6qnv6YoOX58FtOt+Twl1t3evnpF+Y9uVXGu1Dsq/OkpU
BLD/3cN/j1Zs88BOQ8HTj09ghKxKV9o61i5RXjkblhe/g0QB14lJ2AZuP2U6uJTz
8BHuNInxK7hfC9dGjoGMzuuU9PtgD+1G6epgvx0f5wYIWkpSLHLtMjW06OZu7oZS
ChPpYtYnkZuRRGaQR1VF0WCb1hzCebXX1TvrIdjWP+rNq52tyrsmskx+aH12aHQd
uQfgucI/tPcHNRTd0+4lcRF8kOtHeUmJjeYmAmMlUc5rTfHXPxMZPzmbmVEPDg3J
H9p5fmrLyrT77DPAA86tmONrUupsf8pzTSIcgibWclz2offfGCIe0TKT0BQQYKn+
Znev+cEzxzN6EedcCx04c/0/40pjOgLMYnGQB8k3+sHcMfjPopLXpU3qXbN8iYLC
2E1VJw4/VrOkJoV3QSBqVQhrfBKrSP3Hm9Fd5Zg45pF3jqDosC3fDotIf9m2k0SE
8t+I3cdbtTwVcfqvddn9WlMGFtCeyO0njob6pvDMUmAhlIyS2xBKGHlfeZMrr/fQ
9ShSj44byl5OGNBO05rYzfPfea1CsI8KytPVzikw9PrLJhcfHMkxyAna3DwbXkTE
ijy4S3ubedzVD69B37rrfsHX4rv9Cq6gTV1Ca8znYf4wEQ7b3uGsPVAcw0UWjdSZ
jo23zmOtz+YxoSUenV86azkH23q2rs9cfPCt5SNfqSLTcOsatuNVzllzB2qBFmz7
5vjBR/XqDGc2V1czLU/c15Y23NT8GS2K7bSHk82zFSuBJqd0aHjxHuLKi6AQzxxn
eV6/SLQc6/SOv/hGIsxVAZgPeBdrJR0jfhsSbJhnM7OV4ovNdjS7AtJP+v4pXcTp
O+vmMiC6dkwShRZAOokUEcjyDBc4mA54FwAiXya16FI+uEruruM2I0RdGc1P6Jxq
GwmrwdB83SsX+I+XqR3ewJta43j7bnqkvoR8Hm2JX4jVV8N8movqQL7DsCJ8Q0iC
OPCrd0tRJ/8agHt/WLSrsHzxoti9gwXCm80zHmj+qRAMHkYri42ReqkLAOId1nHk
Q9zG311zY5+kHmZ2ZEz3seWX3nrWth5DCYqYd+yrTUlrFRVIBsQa5rkBZC+fHR5G
EPg1Ke45bN+sBgMtfQ4kPESHGMA6zJCnDYQiPtjkZ5CrhF+6GWm5QVzfWoRwXr2Z
IprAgQnSir+hvGksTEFWFe3ObKR5OzzqejJj77yDzvvkAZYmJVTY5jxmjARZy+VZ
sAbOJokrgZI76OHQ+kel22b55IKQVjs3WlgTY/bgt2pmlAsViVC4yIRVl0Q9jFAY
rWXPoFOr5IgzJGmS8xTCu3d2P/PbLTGRi4oHdrGOtslM7cpff//haQQ+SBfsh24f
7oZl4I/WczW2mQUatuWsSv6G53Dgu1AGXGHofztfTXF6uYnaC5BVDNBBDRUCYhZM
NMj0UphjnHmJmhvGyGu9HJEPoLCTnW4niNkECofgvKIn7Yqjs2xeKJpjenhzWfIH
3+BvwT9lTDfP33wPMCtB/Fs6rSi9LRxqRLumoT+AhDa1YRjIR97/3QlB2AjiQNJI
ZEIutrYgbnX6yojDYzhLgQvfP6X9pOOmMwZ4a9DsezRUsKi/VvUNJgb9Y39v5SSD
e2B8SmvKjHlAutRygBAKU9n3ofvjXqFLxn0gsgS1l+DPIlUF8F56tWLNIHCQdVWc
6sSXwGJZg20JtUSQdvTut/KtbdlUdMDoRioqv5UvpN9JpaZYsJwFM2d4wu+nEFIe
jO6j1s35XPwplyX136HBp3PxtfgwhkO2r9VtpQZbfHPHp0WMa3twb6e2LBMN1+cO
14EeocfngDGGWtsn2HMP5yspW3QW2C1tdb6kDBBz56yos2H43STkbVfOkSHXsATu
GNRh7gxE4TeECIOBjL9Rg7aB28ph7OGbsQPQ8W3+X/HLSpOMtCAIIBlq3+F5bSRu
LK7YCjC+NlzhpwmLo933lD/boJpL7oFie+JrYIFPg4dAmMHzDL2cU8h6+XeliaXF
BRB3Rhvsr1vEXqR8EjC+iu2Hng0FYErX0VpaO5ArdSr8eoa5hjiiI91RoKVeYTjO
8Om5k9imuRAEDfDohsLOCLCK3qgjX/IfjMARvW8L0y43PSaE8iVq3Cykw97USHXY
6Ux164+GK34atClMxtTltsbPgi7ix8wSKI3mS/2XXzxXBZeiovsLz5wnNsFAOy5Q
cVhX2eALLApuPmwZpkJr0omTvsCKwleQbTyfaLxp6tfrAedeRiBRAKPdAWn6+jvD
ST7P1pVK7uGxi1c2OzFeLLGAAh+GS29rRXSZkEHdC11iJ4xJQyVJvVR00siQ5pV8
xRRwXqd1rLJPLQHDALVc/5MFIQLaEZFBhVIEnIg3QmbyXPIOUr1daIP1xEd24HL9
5QIO8ebnygaoeGDMQngnJpa5Y757mnvLU2F2sjA4sxYbOikRrSgvNx/Zm61CZTDR
/bByWmchsCQUQPPoX6NE3+yltWHL8OA0ACWdid2VlWSoM9O2bBV63jr2kUGnctki
RxXM2J3+e/fdqv+P7T+NfHpwJrVzUcTo4rpIfeSU5iGjH2419WtzRrlUV5MhN/Bk
3pEWHMIRTM4bZgr8E4aaQiw9Q3aosayeqMueCUtwUYWdX3hA+SJZ8kPR1Nxqwly+
r2+S6ecVpYQL2RN0e6HjIVLse9sQh8xpqMwIo2B3aK39jOI+K+BMzlMsone5LfMP
FQFgnEuLmEf0Z7E5hmaofLzCpzA42kdStZxZ5EHNWJNxvEIs1rgpmXR7GKnK1K8y
LVo6nOHw17i+mdL4Pd8W4knccuQpOamnPhx6Om6NWOG5xNBB/QVYGG4ESxFMDTLJ
AdGxXg75fU24+jhqsV0mCBaZs0ct/srpEaM5MNgmD4OkbDFMLTi98mklyzs+T4qp
aankK3ArBc0cuRVnuGvh2EzBv1AddLvQ4kwP40kKFstNUJXSaN5jhk2bTHE8bevS
XLi+J7qnGpW17nLYB/mKiwyoGwdiLkykKcRpu7xLslmXtMQC/WnZD1xc0NkunfVU
WNFqTO82T99nGWyg7Dv0LmaMc85jBopr6Fatgm1gwR5Yh7HewMnAzfzahSO4u0kB
v2q4i33MzQD35+lrwkZ3vatxI1f1Pc78JXHHCpjn1OpleJZvvzxNoFlHCMj6qA2c
te1YUeMGAZnDO1/2pYZo8Kb595uZ6oHvKhSjzhSHGxE24Gyfm4CxDgAPkeKnVb5m
U8u8DIIIBc2+PHEwJodL5SJ3WszCdeIjgoCBxZ4X+P+jvCpp1wbXI6vmztlZGiMz
f5ochBIrxZgRKEC1APmaAhrGJ8Zv/2FkZIxM1WrN17Rl5TGsnHBjSE5y6hZjnmd8
mzsdEPJdj8bbQ3PHG3zguS9woEXtQw7NeDXFjtXvoRxwml/UXfJGTQGbLkuOmVqw
6BwCzCVucSL1zylXanMnpqZ7ed1fm6r9uyQMzVWnuFcY5qW+oacTmVz4qKfGS8mD
myllzb9QGuzp4j+EfTkgNXOHUbv6cdveW16g2IM8MCyCjzrCiMs9QK3jFcgW4lZo
0BJ2GpufEWiq1YdchCTTqyX+n7LZVWaTqDD0mijxMH9vbpkFYSJJNdSaWdP2iuyu
Aa4xtaayQbfInh0dIwWJLKgnPxQ14WdZnuMbV7YjEsqyDjE6UClrvvy9mo8Wqla0
ciM/WISd/S9QLM7uTUWfk/SnUW+KzcOVKf7cY3r+uibr2XhRLPyc+6ivRWaB4uuH
Rxc7X5CDzhXKH9vUoO2NVYtU5DxzYdfmog3mD+dqi0twjauhjP3SVDFkJI9IJiLd
rLQkTA6m8JQew8KE2dJ9HX58gnHI+13zr2OAQCcZ7n+7+PN7EL7DnsjhtGIKZfrq
jIlHm/hCMUxfqEj9DyB0YyvkPqOqJshOvFwcTwW5UvoIKwpGqPcO0zE3TPrKh8t2
i+dKziPx/11SX+9RwhmqpooIyqBxeKcBMGpYpT4yxdWia7oVh1EeZOIek6PFNQh+
eIsij3nN/eFGB42yY7+oY2LF+akdhUTyX5DqL3t5STkvKT5ie7htgvDau+8J6phQ
H5xNDKBD76KCuEuKpBECLvjn2FMPPuDpfrXUSYq0pKOAMd0yBQPTW9MSi4yAlI5q
ptOyaqBiGTpKgk9EQL8scuqldvOEzgX9rupyiapDXTGGMlcO0XhjgjejKwMfeRpv
ho/fRrrOk3GNEct5rK7U7UTQFNa3FJRZsNH1fvfUjSfkqvDsMuRChU7pGTwm9QSu
0sp5s/HiUgK/vG+MyKTNgjaR2X5mWPLkFMjCYHcuSl/a8cKdPhs0qUy5gxF9/D5H
m5NAcifqBdgmLWWkHHFcrXIljyvReRuDB8waWnZLDiLjvLPDjaAewoe3ebgAjW3r
IaFHIe2FepcTN8n6vhKk7s2LRloj0ZHSCpZig5WIWDFyO/ak8CiHCrw46Mc/gcSA
BIAlj1/Ycg8uUKS8FxD5hxpX4Sc7MzUkk/u2HIVsBoFeiBc9E66STVbixDZiUkbc
XV4FghlScN/OQjuoFXYDGPf7YGQT7PiSPYwL47fwZcYzwcDNKDV6T1OOj7Ocbaw+
ebVT9tR0cMKs+qQvVcq5YAAcC+ao+KNV0H6fT2N6kKIAC4ubYf1f1CtrRiVvlb3X
k3MnlLOBXfhD9KJtlnEeGVJgQnawiOfUADEvf4MOqbIJtE4TP/UxkSU+eHVrmBei
o5FjJHTrjNIxiHUedHYMs0Mk4pWSAn2cZSzAgiVPTivUhUCrR1Dl+TCmKd/tULAX
Fh4JA9tbLHq2NWPZS3QfMYjptbpWaCFK4PFP21bvElyV7PD/aTmvLjWlLPdLDr/0
Yv2NZN6aFKil8RkbduHYE3YrEeVC6PdHnUj96EJJpv6be9lXyPnW6U9LxiK64Pv9
EsPAiHaPM8uOVZJ/VI63IFLKkyPvdeijCxnKHpo/SQiID/51ljUtvO5qiIFlnZo/
ahzx1bKGpegtDCLKZ20D/wNQuAQeAiG6GoThmkFiQTtnsX7m/I6kuByKZL21MbC9
ampfcQxa0gntZ8yPMBZXN3Mv0obdB4sHbwENP/87hhNl/VKmgt7OzHXkawYDLiuH
3ytQU//9AVAYhuKe2fbRupZdyTm4Y2P8mFn74f+5WAqOO3Zd5u6/b2UAZ5+roZ5j
SigTiz8AXqX51R4lx8hCe6kzJnr04VkbzH/VpiRpRmJRUB95FOyA9VLIXNnv7IQ0
kOGKPiOkkUDY9GnxF/lGwDdxO7vTrL0JS8eCEQDIDGaT7y1KQdJ7t+ku0tT0XsOT
JtfId3dWaSLqDNPXc+r3Tt8pVp59n5auLkivd2Kuc5nmUgSO54NUeAMaXKs02FF/
YPjKzeNp/y6DixaEfhxbtRFFbumbULbjx2UWq6dOBgDU1JJbFUDd5DATTCDIffcP
xGo2C5m8jt7uHj6YD1jQ5W6Hpqk2J/wKlBiuUAZBmHqxNKV7BVCx5munQzdJKndi
UPCqVg0xvpuKku5k3YBoo21Ju5buM+ssCeZ0GSDTXC3+KRTKkcc6H2JrULL3Wbv6
kuyBgKhCOIW37RNG7wIG2d2Yo4o0GqN/0PgNfc+R3EvpxJzKmv5vbZ0bLoRC0P11
D23homOT/sbTKiXv2QkurxJomYtRacWpxGInFQzfIpv/sYTM2uSN9BrvodGg0WZd
YnTvavZNIiJOtoyVvSPN+7p4FsfIGG+ZvB6FMg3xyzqh610bYO8zBrD1YsN7VjpX
66wvUuLeTHUUhXTOc5c56UJmTvO1K7irkZGaniDXiLusN3/QEL/Mqg4WgRrxvDEU
va+mFr76CpS5KUPTHXfiKQPNIv5LH+t/MF9LEFxplzq4L60YuJ05rbHSJ3rgfZt7
ukkA6ZnErGz6ICjidNxqPeE4U9yomeifr06OaPzF6vHaphflUeTp1UfzFOIf5nzd
UGrEgJYEDETzrJICkGuZ95SqDbpN0VJd2wfaytX9Lp6yAKd4JUXISbva02bSk8MA
oJXnqZknZxurVZCDwPT2tXCbR4sxeQGN+2nR6n88P2BNHPEXLot0xk9qr/2Vqdsg
GJUZ2IgrV6vxCuhNg34rSGwY+XfAdc30HYAfG7WTQDf7Kh8d+vYFOw4/vt+DlkMK
FBzesleP0PB78JcbWVcwHuKQEw6Rr9fS8zMR2hyVXUZhrCiGlH8Xf7R8Aifpb+xJ
NIt0cPZaiyqDzh0IFDPP8G+1Q3W85gD9Zzx7UFkEelaE1+9NyBqUiORodg5DI2MC
gx0qNILNIxA23Gp5G1BRs+7uQN73JNkREkS7MRDkpREl1yw3Eov0LQEmYa87DuZr
2wQrFKyeYkBc1Jec3O2X6FAl30zb/aCkMn3azfj51HsaDpkso6bxSmRXv7ARxEWg
dvoHMF2yr8pxU3fstyQWAWwFxZMP+FdpUi9PlWPtFwQ28q5G3jlZxK/MM+GoGoFs
hcjoFCAOKPk+TYov4oS6Ll2gMFRuo/bRjKKGFAiIPWd1IvQoB2hOz5qyl4iQe7Gz
2d31qAeyymcUDYIg0Rwvj1DXDWnFur7fusaA0Mro4WZFZMKLfbwqsNg9rOTBkrb5
NdEp12Oj5ys9txR/wpLBYO1sS19ACiimtrbFOAkUpxgEeGoZCqIxw2EdzsqE6VTj
Ri5GGDgtyV3G/AoUP0V1ZP7ZZqKvtLNPgVB3YOHUCCdLk0whrWv5pG59q49xqbU6
BZxv6562B+dpoMbvPS/vDdWIMymLRDPTVQEV75tl9X2m9Ws1Hb41ZL3uPKXCnIeD
Pz7zUc0Yl9u0MkRgFnuTxuy9MGZs6p2UMm+oM30aTTw93lLnvA3B4WOsfU652eiP
cbaLOKX+ISIGhIo4TEd5TEM0BXR0kpS+wF5C2zAQmXfsVMUEERafVIM4UNRQx+wN
D35Dv5lbEWdt/kMZGZmbcDtrmOCozGkypLfDArXJgQCj1kARy9N/cndSwEQQKaTc
xVwVnnkF6cT7BMM9Gzbrs89cpE3d8mw2g1FQeCTeDdktcYxFvOGbUyJWP7DO3Dld
CmXYZ3WA/CEjd5Z4jQ5rhHMQzPNmkOryp+7/OpQ9mwuJJ0IzfDwW+H/uy3+y8rAx
6p7k4KASoGQkKw97D+ltBlFhOn9oFsQQDjVy6pyOE+AVDyMv1Xak4+grEBSFEcqy
Hj9vTetI/gZ12fB2cPUI1+lRxTQqWdQ7t+YVVJ1Q6cA+KVvB6jMmPGz0Ov60Tkw4
SMOe6qeyWe1lMW73C0UnR7yx5lzq4f16Al++kIkwZyqU962sdNFKvFqf4M2AKUXm
ScxAfmmutbBQwFvlBsJlyqbYZBPtNJUkuglII2NnNiZ0sU4EYorIE0ggKvwg3Afo
q4nplFyAlb8b7pT8BQrZhEyido+cf9xfLZalClQRFGbcM8lNvN6dKtBdSIal6Ckq
ogmOpKQ4ldb8Tfse+jt0YmA/LsQULUh5JFouQ2ZWERTEXM+8eS1aGu19AFLOQIOR
gIZBANb4wUtlPVrYs4DUidU0kdO+GFsLrG9zehGgKYPVin6rfUlDTBT+7lHpFL0B
4bzGEnoGspwPCwgJ0yeq/TBUexrZn6GdmpMTO/W4Rx/8LkWM8IK6Gokt3NicpgCq
E/4h1mLmk34MZykoARseJBN6nvHksx57Y6txdMZDwA4qxq/TiQHZEf1OxlHcCXdm
1nYNDvzi2pFTj0qYAeY/xxSio/yJ9eTCHtZd+ablpOZQRnxSzz5p9LGLu7pzRdsW
vtKaAwdXkcL3ihY2OdCSOG/NawykabCecYpAoxPlIfxUYSEdiaoEhZrBtuRZqGLL
1YxFcC11Ti1vRqGjAwHP+bN1KsYJi6xOsFk/I49UcptLcWwzbTyZ0/1ovwaPlGID
Y1W2vAw1b8+7noAINC+l5A+/TTCm1Cwc7ajDPi3f1c0+PwTMjpBa+LN+HDFixNWL
Ii7GEQgz6H+LrdX+vvkQSTHUF0XH+tCHTPl99p1gbEJt/nVaKptgWruhYDtEocwc
f0kjm/6x+VqECWFOiY2mxJAUf30amjIMgDrs7BgfdrkGyZZ9Dt0nJVsQBlb2YgsT
kGnEi67ZH0qliPziFmBAjwbH5v6D/MxiNN2DULsnVI+rPo+pSstvW9rXxDeYwdjD
5hClyYbRDNzpd+/VDQ5vt5z/obXMVBKSHg2QuHW7+MDh5fOyjkzDjZ1DCCpy2wt1
ynwBECBQquFCrw5PnliZ2AV3SX0m/gKluNozaLRBAr1qi5AM5H55ILJqi7Sc/Ou5
bTOZivohbaS1Sm8Q6qKFXMFvWAvTXMM3nk5BswhUc7OifYPOmeqiTRTzV4kBGLhj
QslYnGMhkPjrt2935ha3G0knK2ieNBS0ezfaS6CImTemNdaLkHieJK0SuQokNNdA
gUMgMK8SyR4KQRBnf0j00UNZT0a9Gi/DBk9nGrVOR+UXUKEJ4UPpp1KzCuz2o7wU
eNkXewJ309Sv6vYDba+VzfRMKfg850YzrHPBGQVSPLbBwB2QIkGTuXaxeNhascow
HnK+Hdo/8eX04EKVPKhFKKVUEgfKf4raybDndi8SMMKFjui5vy0I17dUhpSRj1EZ
khT8I2QC19lOLCgq6VU3fNPqL0DicN58kz899OFLa15YZQU9Ylso/ix2ebZSyxgH
RuAqZYrZ1Il7LawI6tEPloVwHXffvCbWPy0KmKrFzN7PqHpkhdhTJAbJIU0Ru7Y4
7ZbEkEsGsCLtE7J++/3J58FcxhXHY/4LIF4jEmaiggqw0LyVcUgwy0m9wCVWb3Z+
J9Y4BiAQm45Wv+81KHofPVV2aSQG+cXeSF3Sq5NUJgm8Db+zHFC0/BTDqUMbQXF0
72i5SJo4WYtPoU45HEpAb5icd1X2oqy72KVrxFhI1Rt0OMdbP7AIDFoldqqt305n
Op77BLeIesG+yWBvhSXiIFSOcb7KlwITpOB0zUB+gPKwnvJBC2qXeRZGcfyNRBKz
Se+e/9h+V8XkZZOFJuNWKXLe4uujjgByvQuPZiNXUXXeRdT7FQRv38aIivpCw5vn
xIQhJyc9mZPSz1JpPUtR+DLPvkkZzFBkxvwjWNDe1oiaF0rDnrhlYPpWsTIP+3wm
xiuvYJ8Rf1z6qz0+j1zWf8zFufUNTtPb5sCf8xE5AkXkyXcdjaWfSP2KAvHdKbuc
UZle9RsO5QCb9RkcSDG1XRPapRW3tDbu/tYJY9zkCc9ZxpLb9Vf6UQfpfT8lHB4A
z/HIfWoUez/1fiPGFDDwPQMd6ZHvN67qYGkB+Jt5/YpTxLy/SbkAeVqUPyNlWHBW
z1MCrSmfgXEgQdzs1lGkfEbP7r/LHvwINHCE+bMkdqwKkkhCW3eLfqxhBjn7vYR1
Qyi1gTUEgI/dRsh8zcr55P8ukUbjTHRCYM/sTqSYqgjsAJEBs5jkv8GMsLVzi0/p
d+csEq/bZgc8tyuJ/bdCi8LhcmAgQ1EjB/tLJFkIusU9qgoxlBu63LyrzFs4frrY
e+VlHfgDjftwDzJ2q0E2VzrPFrZEjGoofd8ciKKMSmEPbTLrDp+GxchAyi1nbYN7
RfVCdl7F5T0Wj9CPF/mqmpD6IE2jzVWjbXnMkaz+gcWgt90gIU71gXqJRMqkWDek
NJTKPVBwv/pe4Pnq4xMWtHZMRrX+9kHg3iq3f5EeqQwrqhn90zgeXL7o24OirNAf
bbowi5qxsfkUXYNCR1vvAbydMw3eSbqMd2tzZS/ThB9i/oS87St1Fv0rVCTDb9c8
Bpvx3xFEzyWmlnI2QSYmdJUxV4IFK7BSaaJ7lUrqZRAxOrTNxwW69Wk4Z6lOKHMJ
xpEttITRFG8YsZ3BRv4vWuX+zZtUAXHZnZH69OX9z5W0B1q1HGl1ZhQv579Lj632
EQnr3Ctbuh+5FKgg9rBg0toHux8IiXyafs96ayx34EC1wEB2DLdNEn+GiukDdFCl
E5ix8Y2fS+yuRm+VhPQJ5jvbYrej0HSoDviL2hq1jfGtVozk8mmh6MgdxJNLwr14
OEdHw3SCr35+GAemGA48P8akjBCJ5Vjv7Pe197p3n1+XMY5RPVrw9MF+OLJxeL1Q
4qD1QPipyNczY2WXTUG9lBtO6jcKJnwDS9uM8N04ldQJ6ZmuIAvvOmiDTgisiDUe
QXq/Z78hzRBIkT5OSS4TTcbj+LXhfvcGZCraiutJG2eCHmQbFqJdliT1U2N6BBdt
Fr8Nobbhv0pSyc03+HmZwP91DoG91YGnD72hF1ULJeTR3FTvTB04YwetlDNnBpKo
ZMZXxNthiIYRVJV7paLCf4E+Yx4gSMkzOAWSIP12Aq/u7ZH4ajUxRgsbLFyftVzu
+hFIMebbyr97BG4BC1JdH0P0omncZXUfrDpoLdaSyil5PXaJhDhJhEHBmXXzt6mI
tQv/Q3ZiCWadFRHr6ADWGGwxsZ6U8ZMqm8uAFpqPFpBP7vsEuxSnF1lo+vHMW/HD
s/WMX0G2+jdbkkDlNkYzN/pVwuH1MLC5d5NhQmrzpU95JVW4IucRpMC6G+KUBGO1
rFuHCh3e2NFJtnugqSxL9hMWT2eOivHX6ScBAhfz4PAuqiM1Ewu17vdU5DNpDyDN
X81cGryY+64vQ/zCOmDXD/Ch4Etb27mJhA1j2LU5Za/EE5sA4bf2uddePwzAxHpc
CdH4CALI7iIO8l8xBkw4r6pN0K7kJkFMhk4gIGymOr+DT5R8Y/P4zh0cxekRJcV3
Nlv2E2O5gj8tm0Mi2YivRqTw1oJVz5F/S7Ll2wpk/fynwMt1A1GDfL83X60lr6sQ
IuOevbmS9wJ3Y7RJHyClwzHxn1l3IDUzwuyW+5ULnvVj6a4sLKd/c2iT2GfTWgYb
O+bAstwRjIfiRhXalIjvUvJaXNwr/HDzpu6IHBywwnUv5LM8bha8HYBIw4LFdFgT
azkaY81k+vz6m5E5yZcXWr5LFQquiUhqtko2zjlNDpdT7oe8Zxi7E3bg/sBacb0V
NKyFbpl22NmjzbDGEmi2085PCGGdrSc608wo6TZHFeuA/Rnv6b7JCOnxIdr39t/R
4vrDGnE04z9mSYbGkGs5uqKk8v0W834/2xTt9SWSsZuAdP9HhX2fbWC9oRorbH2H
+CRdexrRlijNqw+0PA+A9kZFhRR1PXVjxGQ4L71qHoY8k/HQpEXFWH9n66L0ISjp
H8ECGJPXpOy+A3jd/0SzWGXJKOP4M6UD6OANCXfcK0zvidZRIfUhbfSv7g/erJJk
ufQR1EY5tpyari2hUITgu1xRzcHyxbAaDB6JZX85S3ClxfJQZeU8MZSHKVv/UOfK
pUM9b1MSMRVjFcYszvMiCLnhtd8KcDAdYfD96T+l2wuUgygHMwkcLxbMAN65pbLg
J395Bi9hui5GPBDMgqn69l75h/cxyVMUwWAnK8dyluixJiF73gtMzVQTyPawMz6H
VEQVN/0TeLcF/MUCTY2oGm9yFYW/3W4NTw47wBTzEDIX2CVzXf/fAVLURCCKySvw
FvzZ4l8VOfc2bYnDyxCwo2LSBFB+ue635StQDqhdb7hi1iSzDl5yUxGD3g4HhBn5
77hYFYyu8XNoJc74Ix9G4X5dpHNpf/QCH9gH30hJm2pOrlCcPgLuW0MksAp63Iya
5eDc+C5xX1OdekI/tPLd7PqPrdN5NnAsKplkxL/6RQs9aCAmIAwP/HxyIy5GtbSB
ByY5X32ubzAOhGI0Na8nI+pIrOR4CJfxHbpyzIRQwz+IsxKE3GxR0Dz4ZM+iqOqz
ehtNbvPWDtw0SQ/LSmaAbpq5rxXUDgAQmW2PbFys0xPKSnJIj2AXvdsOyvX7xM4y
d9JIIofXhJcDuqMLdA4ogo6mE1iSMIpb3g0HdIPv+Bn5e/pVj0L5e7o/lroE819m
LLJJhPfM0Cqn1lujEdg2HBeJW683qdSyvuG7gnpieO9Tt75HUNZxeof6jzZbbtYD
Faqyd9yJ5ETDpqsCuYncbLT8nxaUp3PY9MiDc0rurTF+qT5UgE55eONk2T2Ffq2d
1iWj89QUZrT/fJs10aDKclc2cQDxZErUJfKjDuF0Mwca5dlO0/Dx4mezK9HmHxST
dcwzEhxZIy7ezmYXnA1OPD327jlblzVLX6pz8/15bndqj1VAMk5c2SfEAWTaB4Y1
TA3YrwIiLRW1yMUR9V25h6uWSmWNWGEGC2tB2p4Us6rL8h8pQsmM9xUBWXGkzprv
xfwoOk/bJbNw9iGXki4y4BmU1ODSXSWeA8QhErJLZYs1DX2hieVRBYn3BjE0QWH6
Vt700AOE6by+SSaw9XfT7c2BQfp1+7x2wV8/Fl4PWE+02fj8mSGu6wnAhmLT3xF5
QqWS5WzG6cUNE3RnPhqmxL3/RywVvafNpVgU8rIIlfiYEdL64wCtH9hW7N5ahITq
iIM3J0erfS2Pd5PXQJYR38Ik5pELaIeeqa7nezv2XFKcA+Hiztb4RSTuAkm1zfIA
uHxghJbGsrDdlG6/e14jodJX8pJ9M81Xs5s+D6vHHFiNJL1yN0sTouIzqfk8FqL7
VBvwp6d1A+Ps1P8tt267ZYmXfph+QdvqHD7W5EXKL7MlHmTypLf3TqNZQE825VSG
lxlniCnXOGXYPSA+jQEYLtbSCYnBsKYyUeDMvlXYoj1376KTwk4sFNf292Jh/wgq
zZ81bM38qgeFIkWdxwT3N5MLuNINXaxHQaRlN2ERmg47+JNsBgpQFs+Wk1ETbJjk
xU8BQkPWWN/1nuWOTEocpaoRTVUncYbOJ315qTeXRfgr+EEYM7HmnQEDGjsgO5SK
vIH3mko/SJQwHGG/dvp0PmWlZvGA4+JLTp28y8IkgS3/IRcP0KNTLTlaGWJcyUrC
z18+Nt5W6QYzXJ/faM4GW1mKtMmVTkJiF0uvDMkGvg45dr7WeBR4XAQ8HDk0xJuU
Pkh8CufZqnMy37CyBxGJm5ULHmgWcRKM3aVKUKs9ykjrNoyRBcZU0HINgVvcyj6U
s8bv5Pk9kmPeKpEmkQWzAOtNqF2koOf79DDEDbmAnHMXtPkXXXVz0qY39IMBXcn/
Eiqaau/PNv2NKEDP7ZyyR3QHVCtdfNdHQtKBFAMOm8rCj+poReZbajZyw46Ocisq
jAZmO+LmTQ5hHKastM5+lP2J7xmA8JczS6IM4kCilrtviuxMTTf5YSEiM3WVUSRw
xeq0xGFGVs50GVMt5wqA2qbdn7lM1HUfnCnL2znk062Em1HScGc/kTQbO/EklBWo
Ka7djupjKbzUBRiuhNb3f1aLFz/o7q3SpLZsvnjHYTAb8K8EFhGNnR0exyOxo/Xj
KvL/JEyWi9wiSj2rnnuAG4qLoT+JVOSu0npgUACxNGZruXG9qGNzzT0Wd63gEuYt
R+xy2PVXfgmn/tRxQKb1Uq1sqNYfLvfGkwCQW1MsGYn2pa0Mc+Gkheep06bNmjiz
sFhSILnKhOuHfyODcEB6CGCvciIhe6DmxAE57MUnvmEP3CroKFjzSNoc185r9L3R
4VRu4xRxmBWCd1EOydMJqFNK1mOf+6tEafEb6Uvoq89/XTbQwzfM+zkas0bXgEKc
YizpXC1rRErXHP0fesG1KO1TEu/8j+v3En6O6v2AjjqQgHHSLLiqeNs4KTyK1QKW
Xmt4Rw35iSwFqYFwn9AOB/1LszITVkM1EC0TLOCkmSNI4ah34rZ9rvKCPbhf5c5v
gw1P3mWvT8UBbiu0zzZ3VWdoac+PMHxbiljUvKUiGJz0XNf6IDX0iVfFQKRO2T9k
ozrumsYyf4lMW18p8IFHwIc3JoOg79AF2u6e0/IP8pTXT4+us/+F8zB0hcymKtVb
K92gKzEy8fqgsV8G28x7QaTlOxiEcz/L4Kxac2In/IXStEvW4T5vpuYTg7Pl6toW
YuiCkjVYz2lBtLU13ePZSCo8aiZLOH60Mg13/CJa50r58oylw0VPFCpilwRlPoar
Qb3pxG2xf0U2WOY37eXDWnCT0YohgZBkBUO3N2dl+KvyhQZL35FosEiwN++G56NE
+Vs/ExdsuOtPc4HFyG18W70PgG2HHpCocK/cT+n2yoztKU6npRgieyeNR7L9SOyK
ApI+FxoWCB1fGb0Rf8vlxyBXpjEDOgX7NboHV8K8D8KkNNyAcPDFaKfV3H7G8jH/
lwVEqqUWb7J9K+4qaqXhk6XGpLv6Dt3rKVEoRp1xxldke3wmy8P+ppurMA4rYi7X
uRN4qSDb4Ca67ath/LsO8py7BODUlRkU7qDFDVH4wmX4OZOjAWK66Mm9gxwYgWsQ
gffdNXvqQoM37043Xt70HGXPjCecbtk0z0jjY2D6Y2QB/G33bhWhxc3dzY//bTRN
uDMQx2559FCJzDQk1mpjVUN3NSzCOLV1p6gh+DRzLbK1GbJk+3p6Z/vJXNQE6fGe
8+1r0mUqmoqGvDYbpKA06fkL5irCFVS6Ph+OYC1L8eXrdERl38gBuwzV1omI+DH8
y/XrPdoMhx9OqoymS9dnjGuVQJaGPaLBFjL2svVLXDb0FKxD6D0DNGpeVRoOjN9z
GD0F1IyN1gtfYh+TkumeVoGqxGXhMJpByVsIFNSMtoEooZ71lE0feiqu4VbDibZq
2gMxv6x8QtZ2ucwsAUOzLs7EeVuRsLGslWiUq8M64xoee0j5F7TajystupcmB2Uk
7qBvoa1Itl7kdorXtbLp8oE51x2nKtHWrSRij2tRuiXqVn+JBkyW1aCJKZ2D6z2v
5yEuD9Jl06Ci4uCoxvGg/tpRJFAXkpBRNK1+FX7x5+A05LWnssxDyP5J1RBnUfnw
LxLIFuVlxtN/aIwGAFXv3uwqAfW5s6GGJrquZc6QzBaaBfLf0GJQPbvFpY1gmKBW
okA9Ebf6Ju8XzfX/qAWumCSebKxDG0GYiYSnX1IQFFspHSTgKDPepYKVAX/qX4hV
Fk7dGwdZ7pfEwcRr7ZvW5A+ROE1cylisp6AGvmZusof5i4PDzwZgr7BKLA/56PTW
9qRB8BP7tihTHoOsJeaNGdoKOrEClRYTsyfv/1I3BdTynFkpHXEByU4dF9+PhH/X
TfMhCIuZfkvoaCIEpU1+5Qy4HwtJqG7KovRqe6KTBz51FeSdnNcs6WGuFPqBiohy
E2vO1iT1IqmJhJOtqKRbApa8lfm8iX73016QQdK3L2rUBNB7Onjv6eQTEREezV1Q
Ca7OZVIDYXeyZJNp8Ws2HrdZCXFUvZf7W2U+GvMeaecHaceiTSb91DgeK6Z7nKyE
z+PGIZagoBOvkIIve/E8cdhcvD2VDcEO8f13RN8SHbDYoRkAaiCB2ezKsPRcF27X
CKU8BDkx86hsqbmI9o0kGzEsICxRy8udaacOnPaP+ekuSvd/JtX4owbieIIqVCNf
geCoqSpWQ8zVXMNEf2Wyqbfl21S3fkKr4JuQWeAjGrDyLgQx48UdmV8zV+Q+7CzF
lQx+W/Ty3cBxZukCuMf0iq1aQFU76n3DFq8HdWc6PWIJdz7nSIAvl93rQFZTFu/E
l/yxJHW1T0Evm0EDwjo7jrOOMlVOzCWNkGQI32WN3LEw3Aj0vNvueS8XxQ9WlWVo
7NZQy2HwTkYNnVhHwtln1GNL2E6yXy8pN58mjo4AajOfyeuJEvGdT8HHaR4EU9zf
ehCW/7QF1P63GFAnAT4U4JG7fsm0yzbyDNFzk2RHyikq661h9iqVepPgeZ8LOTUz
YGAmKegqNn6P5KVsb4tnDFfWiNe6q0dyIBg9DYjOgZ07Po3z/x9fyxIpjPQFzHth
biEsn52Ra9ra8eVjm2SVbGBsJqvit3B5npvPDjWiMakxt1aEbFh/lbuKz6P5gyac
LFccsGYr6FjXI3vwwjMat9Jk5TjGq3YIhSr1dBfZAoEaca+PgZ0K7Syp9DrTTgOo
siwD43PHIohSyZuzhIUJ+h4KigE2jNaSf2EvAWc69e0TkoiOV5kTEKEOCV15wvkK
af8EVG5wnmIKniAFWp4DhtxbSOD5WuJ366JGpcGbKWCGXhRiZRwHeqt7jg28DPr7
7t/B+YteY6/UFGYLPqhbcSpi9UVht7oJ7BxinRC7Bpg=
`protect END_PROTECTED
