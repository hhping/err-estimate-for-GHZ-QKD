`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zj4dgwup37EBpUuFJiAkMMoQ4N/lfY+xPwUxCaTDY/15fV85TBdL8DAqVhkMtK+D
O7C9WIB1Off5/e4aNr28i7wD94KvE8mZYhf6wG7dHXMzhnNLtMiqZ7zyLOoFd9Yn
RmNR4RqBHzYNFi3O0mhvBje7UxRUkzGaHfOx3+ClWAZlTL3ItEuDqvYl2qtCxgZ2
TQFxLIj+7DnYrd2yQY2TCjChgoqf+PJ3HVXmUZqzdIMZZDXQ/Kx574d+8Wz/ezGT
emwjMwdPZCjHJUlEyX1v0DIBMJCzg36pVlwWxyE7JnDQp38LO5zi4tejNfnAvZpN
OaJS/VSYhpknw/rAdSHF7AWPGozzs10aWwynxoqlyCG61mYp2Bb1SVRpsm39JhWV
0mQ2moUbwFi7pq8fVu0wsfmymp+K/pul2u8gxYbwIZeTkb8mooArZlPb/cYgzufs
Jv7ca7HWv9TDISa12AmvVy37O+mUZML4LEjEfrhABG8nX+dUZWlRRSSfKSTZZGNI
iFIzKvBTSEfHXPMIZUMoyGLZSbro5Tpm22EZpfsRgEde3rKAQwb0oHOocgzgwUDe
bSQqQvg39aO9sGGc7RdRrvv/nzJ2WeGAndNHW+1EVCkVm0f5TLf+3EThTDA1ADRs
iLU1C5x+5LWBhQnJ1wsX6eWsDPy5MvKBE7+/gIaF1n/WGLEYv7yPYuhbxYI8O90M
GLoQ9a5JapdIE80IDR8k7Spft8zM2aUvly/BDjfi63J4B36x2/HQ4IKZszP9roL5
yZwDwfs+qva9vfNBwDum5CIDuSwytM8XxNBjZuU6ZzPbDKOd0UqyF+ow5bIqfVOM
xwJQ45C87xMEPCzxkOkE1EvCHgsAo/diCDxJJGZOTbHsrW6onAlmFwWpOrO2CsgQ
2iQJwP0OpTD01CrV25qXlxfm2EmQ2XkBlV1opnP0vtxBCEwbL4ySfWd0IO/Ge+dO
Tua5O68dUtwnUXIR618ik8tk6kgnGRGlnYgZ2n26ooMXPgxLFJLMVIfWNyHtJACF
woGuqaj5m/yktrigwlBQJk9dz0i7YZ+s4tbxMgdb6LHbXtbfBlkfGSuU2UI2Sv1j
ZHV2IC3+7jBakE21HvaKYJ0r+F6v+Kw+9iNYl+YEpytBjEuWiefisqznUUHVPz9o
UFWnbFqbtkVaMKHvuCxYdhGtLb+dei73THaidYRsODNTxAWxRPA03oPxDHMpv3yG
MIwzbdZqK4a8xx+BJECQcekXy314+8TR7FbeKCPO81JpXq1awbMipFwvT19auRXe
PRIdLsY4RFp5enT0B6NxLIbKEcdLi380itbApaAU4ZidSDMtdI40avWoDkYb5kDE
hX7ZyyE2BjPK8pxVRw/1/89Ko05F7V7WxhnO2b2/+ru9eU6330iL084jtpfPDWA8
SkCNnLYe6l7B1IXe852AbBSJdyS/nHWxDVAM9zKo3wW+5G2ELHSttnNonxIBI0dt
qCqubWVVQTVAafAF7mq88NGg+46vyI8wXZUTgPi8N5Zc3bpY/0roB1d/q2jHLt2r
gvaefHV4HYYMly1mD/UYM+Pybai/paxCeGvMLCSF7dFrZYAWVrueOu+37Ogo633d
os0FiwdgEOadXJuYfTwn8+t49n41joty3+8XaPphpWxYZeIN7IbTtnVwkBZN6919
Zp5Mu04pSLzT8Ae+nhwhYSihG+qFJhVnNKqIfbFv2+PwmrE+eWOnbM37aOh0RVI4
EgVu1FN0qyD73Dc0dgW0yHgWnVW9KuHGy7dluw/dDJNk8VNJuUoJCKZMjEnbZxwY
fFsaa6bUgrv8DpyQJI0XSE9rfXkvcToCnyfzqBytR1GPzWnEetNMyS2WJJ4x0PFZ
AbZ9CvyIeFQ2nXBVK7eEdZ+SwwbfDvxZxjSoKqql0Bh7eMva36DF6/QM1jKXjB/P
bElAwTPcSseoLn1OXYgqeekwHtSHiOl3tcfLKC9lI5eIAL5doOI5phWBSxbmQNRR
/HUsSioXVGRqH/HAVyRoouNBWoHdd6jwNx1XwKgGg/5qpVIv/kFVOVdwNc8nvjaJ
u30RJVG3zPZJmQV+vhH7P9nsMp4VyT8I1cAdh+LXQhMKpebyGWsF0hSfbMbKSOwk
e1gxX+5whC+ShyKXi1YUCIcADsqOHkti4P3k0Zk/DECYcAq4YP8auYpqoOL9UjQk
Ml1L+s64CjvgU/MyTAB7HvDhXQ6CDjA0skwYBdx0TK5hLMPDETYr2bTu1/2LZ2S6
FOseyrOTCm6M1CFRMMK4EveEkXHsAgbOJYrQuUZDpEA72BSAQgqQqB63Cq+MUJ1H
A0vpHTEbrogOpvNUJrQcTJX6S7njz79SlFBHHBTK6wC2jqIjsbV3jfxAHmrEk8aX
R3hNPJyOg5kdBmGQrS+lQiGVTVrdW8K0H9VnW6Uxe4cQT5ridR8Y521SH98RIs/i
j8/9Q2aeOBOoi9bsJclJbzz/bS70ECgkKPx1fkeHwOOzKKzGRFJkohH5lhljmYcf
TJ7c94oKZo6XhHn4DxBsiARi3Iubwd4brkpNfD+05Gh7qT7w6fWjJkjEU2EhfDBY
xm2rVWvCChohpzVilQ2pXPQfErVnWdkQfYaFjv/wOKjnke3j/EkJoz0kwnOjusN7
PM73n+lvSIH3Nh6Lzz9YdMZnr3+/eDpvQxAnq3asK5H7IxZObuHl1iHHKCt8tFXA
77S5/ufXiuDKKWK6Z/ZrhLXHZmBe48tGwVBfVj3jSEyIn0BMw1I6EXrTpEZdp7vi
pnM3PVuEHAUhNQzAnqtDC5X8smq3vUlHwZEUa+IeehpzHtL8ccBrg12zs1dqIESD
4gdJMEiD3jjB9PaeRZp+2kT0tOqhm0+KMLqPCnC+zhfyI/Oig6NhsODpnlQ7EVcG
HGR0ublnLXe4hcfOwe6XVvQhThE/vc6eBsBkZqVxLFDEe13Jg/I2jYjiBueq3gBM
GEX02HtMRvg6Tmu0iTYKvUZSqURMmrSpii5mjPokwYQXkhNrLdgwF5VLedNgoshr
bNKIS5UC09XGnMMf+j0Y4nO2IPN2ZSTAWtXAuZwIQW+s5aGcYqU6nC8ZBmRuA57D
h3aSzza96I+b5KrOOLedFIPyMqceepegZ4N5AVg7JYclvoSpdxLzYNHLRGmtN+yb
cGauEB3Q8HX+ZvdFzCrSh9ZKtE6lN7BDp/4wl0ZXPtuPuiyQ4OaM/jHte8/NGeab
8eqMcBzwegL7pw2CgLRSI7urzmje8usudXwqlni1W7jY9S8jbOmeJR4zw6g8mfDW
F5YXc/A3Dqs+V5vAG23aQL/ENMyz5GF2bKOjUIm5EfFYRU5cK+8vFdpW5AQKMsUE
XXbaNGV0lTq9hMpV8Mu1EcAmUQe1KGzHWkgf8L/dZOoqKEoWHICzX4T+MaVp+Tvz
fqxRyVuGa75ZWBG63oyEQnqaAeFpldnPvCGmy33VG6mt1FTJq7dD4rKle2oUViV0
hlVdfxnPZceBnZyZdDRGlo5yLB93j9Pj+Iczm7TNa8W3fFC1OeXy6ot8bBw+tyxI
ZaVWNccuu4MvX6JRoSEeFHJ0vMAE+WOrfiK3p4CVXPuw/H8aniRDHxPWepkxA1+e
rgWcoWuaClW+hs/J8nTGQzg8Uplix1ZLjJv3Pb/X8393kqQSiA6MC/8FhvZQJ5Yp
KVHnVumc20OGa3qusDqCYJXreuIhzwX++GK+pa5NXB6udj/DZT7ldYAmo/jXws34
asAKYx7dMRVcIMRpfaLNJR2j6BV04FiINKucfUVWugHW+XiWgBBn60Jh7+oMg7pk
/lr/0ICoBDs/nGs0hJPeBS58tOebB1fzzJvgJ/m8KbWCtu+H21TBNmqbCFbiy2DI
jE/A3hnJhHPsKyRIZ3B6OUe4mC4rE8/CHtc+MseV1ziZh9yIJANHSVCvjjzu6/MG
AA4QGapRSUbcm3aeSJMIWR5N3UTDu5EBTPZN+4DYachgQK+UqPLpisPmsL6a59yF
8usF9qCs35xGiPSNw2HuxHrJq8LVGaZCtBU1snw490vd7gmORDyTSKV8Ngd2JuFM
VS/DXtfKUgPjKSvZ/BBfhxI2dimEYNq9oMEUeM/wClwvSioRe7GQ674zVm2lncuX
eICgiAk78ry1yFn3WJGt6scL3xDIgVVWkJ4uwodzQIe0mUPUOECAZ6VJFzKCqIfA
Gl7PtSKGtXJbqs85Kiv/8KQBrGXg9Qjklr/bhk5kSDnbwkUKJ0PGlUdCtDsVCKzR
JwaXXmaEPFGDHiHYiVc/VL4FQQz1g7A6LYX502I+ilj9SN2dpmMl4pHrIsbURv2z
t5+9gFvm2qr1BksFOK8hlORhZnbnt4OAP7oa/5NetaoreG2MLp/peXHVey3mF5Th
9sp2CkW3soLZp2XCcbQF3ekvkpjQDUqdrcRnhOR4UPduL/kF59HscWu+f3Fi465A
LPbQc/2XHKz1DfiFIidCcgqez6tirxn61H4fj27iT3oB7hcbrrCzt2rvRgPKmnv/
yfxaOM6UjJmCiIAjj6W7Fc9zW60W4ak7C8h7llWvXyz/c9BUz09LtWMvsL7PByxK
OjGEDQnXPrYE/ebYN3ZZ5Arc1U/3ncN0HFbbBwicXXj28v+cZui7ThPBjQDNSXXb
HCHICeAwVXwoi88/V419KqPlJXRQH+QejaEnfR9bD43JmV+7dvrDPpPSvfJkFYVj
jbvAtL/7sukBXgW+fWHNhbRfFRr3AUzPeNba+KInp0Gc/iLwSMkmAnRfPVfTxFv7
Z8HjBQvkxw3Hc2HJsVHWHQaZZyekHll0bnDvZdHBFCDCDKaEoMLQlabl+92HvewH
x9FsRfonpjW3ugSF3iW2upmrY2u5CXYLNahaFRy2vU1khLanztV3hNXQVV4xwbbR
QJnzrIHNIyTc/VW6Wg6jHPGa7Q9VKRMjWVFaluzmCaXn0CjMMu2oyz0qPH1HajbT
+XC3DR8QAS5umZ31FzvkV8OOZst1Pk9U6ZUAzv8IoNQQaQgjrfW82F4NmrZmcx0B
F8IdkrinClxU9x3KX4UFDI4QzNVIbw1WDxkV+Ba6AAvttCgbC//V3I+ymeOur7+3
kdzXrMwOD3jEtxJr8KJwseNP7SDjgleGtnGuv6pyR/KILYxevnXtk6BDfIH4AHTa
0Vc5bonzPMwN+K8gFLbuUh7kLNJHkzeesSE3rbOYXo/OeWzhhOek3QYdHoeYp8bA
BqFfwdC/kI3eOcUOMEY+LUrQ5KxUdAjTT0lC3ZM7YIfXuC5LJHbmkt38w62Vv+9U
g+uirnvVEldHhbWDbnnfL7FyWLgsYFyUKFNtJHUNXmu46zZhCQ1pq3JHq/jyBvPp
KY75eHTbTh8yeV2oU1qlZpyZyUa4eiSfybiCwwNcqZur3aiRy2bYflif8C5z/GsB
IY9NsI6gB/3k93o/Wfaq5jWD0hB+2V4VjK9OLGExFknEbKHBNGHNegl6IoivkhMW
FL0ZGV5RqHTtQzquOR2NMbPpsd+ec6nFeXEse5lj0uU6tEPX+4nBbAeX65ImZBTA
wiOF+wv00+/NkXvIcm168WozHFwuIyQmBzYGm4W85/whZmTf2hTqRL7uLvBpd/gW
/BUvpmC+euj3osU4AyWnTqmGCIdyf6duJFFZUZ6W0h4RuXM/l7v4GkeJcsncXL84
HZXMHWKoPDTEWNY/CBgP4fm+MHYgSPJBAssudw4wnjKOrTdxJYWBGTZXiIKR4Q/X
AhMW78oqu6hJxAC0OawwCbq3yKgTXzFgIEKPd2XFeVmz9zucsL7Qt3cTTq0sEIev
0ogqtyGqmms7HiRL68ZiHZMcJJwL0cIIX+gSsDvISOH3sW7X9IbaiJBvQvscpKAl
xyxugwLRsWCyBeU1EWzpmw6QRQ9rpEDX594Xd3TfbbPTG7mkgHmAIdZM8yrodUoG
0rP5pkTuFl6wLkfTE8WExLN/0Wk2FZbAd8IJsrJHgf3gj2+i3ZHStAS8eCa/Yvpl
0icXjuZ7IF+3jye7/Wb8FIvbWkbVXbuitIflJmJNKrBCcowyYbYJqv3crc1f2mVD
H18Ep+4KIqHa9wnsTxMo4EbF4wRJS89TlRepWYU0CR2+iEB23/pPWI+iUEA7UCM5
1uLOmn4wnppksp+yrHrHjQvP+b0LRIuGuiIkaiY/6SAQ3cq2JX5+PKW+LPm3EPmJ
IGLBek2RxNwz/VyJn4WPKNinsQCJo6JqFieu/RmeMhIQnlw0bfR1cVkE8C/wDEfu
QAQp0zEdDwFvi7fhm5MDENweGGnBVUyF4wh5PpS819hN9yCFcFbD7ItbjL5zfi+q
iZRBa8SFIrTzGmNHKjO/NyHfYLp7PIVhAx15/ygnuGmxhYXI18yHL9o1Cw55/4yG
EEH15gFZ/kPu/arLvX7UfrmrggqIf0twWIT4IeklGtHIZYUTAK9vniCcxMVd3tUx
ViVlLc/rC2rLw90yE3BWvy5iretP7vMPn6e+mul6FxCQ59Yg/BJqvrdfxzbF6BPG
HCbHZceCRWqh81j+y663bsr1FiaNlh9ppQXXPPFBvDhFr3MgkXWAJ/COQizYguNv
KB6C5uDbXz5Bg3Xtk6CZh7tN6eqC+3IjDgYB+jULUFZPhZgxJ4jyFA59TMVYHcHa
sd0tBEyaMaqOv1A4GNqtkRQHsyTK1xhAxuP80L4jnXOm5jNEtANZOrnOmvmW0tBN
umqbCfrV5o5dqjER+IFBdXcrf0O6l6MNoKtaBcbdMITYyVA/faU62Zp1oIa7i5oY
yorZHDvyH63e2casYcFl3nKuXLavMJ51hv3A7e9ZGWTAlci/r6sK9QNWCzRf2sxs
Q6Y2d01tI1GPaWvkVaLZNZqxhqv2HMw0LoALESDU2hj3aTJc/mqY9hGrBPYlUwKc
u+v+UQUHNJfZ7ElTSlxklGXXCPJPyQH9dje3gz5bkbEnL09R/EzW8qGSdsoUfFCJ
9ODJxXRYmA9DGIedmDmi+tuZ58zdazkBvvPDHsglSG1TTMI9q9o3YgTZpL+JVl12
0OXsyUg+ADoOUoiW3pIeHfcKuLozlniSHIUwYbDDTHkVvnuqYErHd1w0zA/kxGc9
1NC8DFPdbvNTDqpawPKCj66JOalMMrC+pV6FXEnjLDIqgZxSXTrb3+iCizSzeGuo
j3ONlJkZGCncoVTxHPHYryY/iy7mhE1gidi+T+7h6zkfBaWpExellkpm+ekjwnSu
XePkwpH4H/x1VjEwIzQcREsLJbTmQ2JHkPaMG55YnE+t83wdPHbjOAtobunlVjkc
MnpjpeAbq1CtO41EUgX4xl7WvCr+1kcMSuDECJ8HKAUOFevU6A8IFo7D7NKhK4OT
4ENKOx3TJo6WlmxO/jMpnfHghIzh+BkjWOFuFm29/1FdW20ovDdgVtxdvABYcIT2
GVM4ChEzPbtCpepKFL8lVw88Ty2OuxzyMLa1CnQ1UTKGJ5xs/lSkbFmg/T+2n+7W
8lnDeuz+aDOv755kkknGUVubmyXN0KHMg5TS8NmcY+Sz9JtRP6B8lOi6Ivv4S1R4
A29FhzctsAr0UB/0R062rq8FPdHzXkcoA/MeB0hNJOyTTMagapASpcSd+FU8X47p
ldYKuUkOPJR+xhprIwEVej3ySbET4N65pypnQCOPN4Yj7cnbSIerUAVbdrHOpPIy
iCo9EvtWJkwJC4x/RzG4w9Al4hsZBXIk2DvgePxXtt3jsLcDmHReYAEBC61tu7Md
4DMCqy2MsBU+d3ahtViKp1BBFIa+zlq2K6QRFbR3stJhSAe/eIxyxvHcp3BR4j02
Uh98R8cK++OwXK6DIP1217Rg7YB+0tmpwt6Ifaky/V/4Cmz541A9RF/OWIfQEcqb
8J7JKKoOecSyhy3gLDlNoJkziZy9A7VcAl/kFjJ+43unt+iafpIdVCJDu/Btnszz
YVkfzltt1H50xlnyHRb29W0t0u5dNV5AzJlZNNH2+k2R7Aypob8IJoc6X6Z0Kpcg
O6KIGtLoIEbCFBODK7CDSnPsSWaAuCyQd/uRjjGfrp2k7IIduId77rqxvk7S6bgP
ORIcYaRSqVcyXqHG5cwzPPTANgW2VIL1CWn7XJYC35rVweBcmS5LMEZWxz5RjdwZ
A0NxizzCQjClJeUzxDg9SvaFAkaJ3qTl+/UU5Dv7SCBdPnCRhk+lm98OOmZS/OaA
fvuejzg1Yfx+U91WbzezITqo6dX+WoOTTzFyAavm/9Chuefovy1EPrsn//hh7Sxt
1zIkbCUsNTms2ZhblymYhGC/5jTRoUwobSKSFUDrK/cbYcmLrrAfbT2LzyN8emX8
YVbxNkah0zovCNQn2WZhg+6Ydx1WrdvGgnka7hN3NMpnpXAporrnTDN5nEEDnOdU
`protect END_PROTECTED
