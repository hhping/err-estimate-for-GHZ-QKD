`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2hVeAfk6nX77txbqiH0QYsZBam4vVFZuc+y5fMv+9tRP7WAo10XdVFn7lXRvn5L
fuCTC1JK5dz0wGQaVMHFc8eb7M/fV4/5+qSiqPNL8/1Tr9GSYNNZ5FJ6GjM4+RWX
IIqhCmAJrZYfiyLy6KNbXPCfBDIdpzbgm9L7d8OqvKPEfLLREDmU6PATiR4ilewt
BhYFnZetm6St8//E/6IdKMwI4xg+G88wbkBFpvbfWcEwMsNmoW60RIQSduu3DtRC
O8RDdlouOEd5FTuwS6wnLk4bt6vWInK0hqnPBLRB5YqybHCGeVttrlLm/bplJSh9
miRIXh4pf66RB1Vp4jujPbE6sy94vEKnp5yO3l6+6eRbcPgs9MZYmMK0D7Fpvy7n
+TSM0KpEzNRtTMzvaoJiLt8C6y6t0fYcsTFV8hLGc3Y1cNuDRgxDU4c/DwNAqpw9
505E7ItPZJjLvQ2mE4OD02245UKy6k5buuHfa4dA0J7KAlpsRglRwMOkCBluYa8V
qqJ8H4n6UXDx7pOH8BvOaYxpm4gwvZYPlIHRyGZkNGignKfIbaDCby0w5sIWeX1z
qdg81KLku4HzXcnF5Ir6MdVJ/4lpnKLGQ0mTuznPPQi2o191HJ7hqYHznZrqbzI3
`protect END_PROTECTED
