`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJLnK6wthc/1CH3jJ29TTTMPeKLxJLHwX7Suc0HEJLJ/Q4pkWhByCebAvkxzcr2g
0asmdm5qjT7hof7Gpnf7GdXh3U7OT9y2mwzTRTRx6KuRYq6tUv+K8xVZVkkaQVxt
9m7QBAwj3cHNQoNLGswqdqEjBK7+Km03cZV1eqWC+MXWu2aOMeY/DSAkti262Dkw
IdAbFeASazGZwvOaGPBz8HFjeiRuALGIPGY0MDfnD9czeIejNGPqfG0t0wah3xWQ
BIlejxZmH++/r2OUgSqjy0M39188blXNl0lZSwT6TzAYsx1YtrY3D9BQxb0e8yEg
FOgD6CYRKsNhxGXqgd4tU48tXFQmuesCqc2CJEa9NxnbqqesRYpFdtKP7ybwInmS
ZdPIh5XoN83kwWmts6lexvoqV7sPvDP7GwE6d6u+nFI6u/iOpFI4RudzaZEon59Q
2cQFFGoSHHxdOZG4dYU4MwfpFW8kF0/ZVFmgP7AZ5j08h3O5mRsEqVgCRru2o0LJ
YiDSowWpLniPa/y9va1mB6rNT1ZAe82moHFFTBOfiv962lJ4StZTWSpE9mhG5Mj4
H0pPLXLl+Ob0sr+LTQ2FJuqlSBTawQqsGdjW8tRn+TRTWTu4BqoeltqFt7Lw8ovw
Y3pZX/b2W7WcyRFnVYye2OWw4wnCB2Vj6xl+lNGsotFrAq4KpCebM+PW6zfGbhcW
ysOQyrGFuOa5OqhFRSo13By+AMPm79XUYsqZ9/gDFJu+v9njUjsK95Wp080DW7QV
JqTR1CVJWEqDYHxiqwXfSvYIQ/qHT0sBib2YItu5saFzYVUlcuDiMNQMdvuAgwOw
2DtvijqHYD867BzAt3STsP7dOlg6I4ELMJJ7ZZBRmduX181/8zBxN7pm9dp6kvbq
6lI0Savt3Bnu2ywy2yFWoXd3gUILFIc2yejTS3xMaq0S0QzBOW6v5YzAtpNZ4jJ2
zDFIRQmOTQNbaan9MzA+n/Ot7k7fAM1L6gDD7rzPt4B53NzxGh4gSA76PyTEj03l
tHfO9apBFpopfhZtYZB1cujZFrMTPjeb9Qnl7e5FUk+/kuUmjWzVirY5YCU+D6Lh
lAeTnN/Pk3RfqQkptH4JgRJoQRp2mJYCh7bbCtjwaqQJK6k+974aPznSLblUVOcN
nr36wXZcSrwyNDWJ7UZB8C81tTmf1YY4aL2RKbDizrXMejNt2XZm75noYzfAtdEJ
`protect END_PROTECTED
