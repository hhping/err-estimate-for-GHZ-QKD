`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EzfCHhytzAPNDk2L87Pbm/eJS//DJqLzUc4odi1bBLHn6B+Z0L/w7yABlaMOHuhx
LhtEMpW3DgLaYc9Uuh+nN1YARZoPMzHfLx6KBmX2aLuIG4jFynAZSz+jgbYlTHgK
VR36j8shw1QvuXI7rIKC0XjFa00v6HeqEIzzh8SHL+RnnJ8Al59nTOrSF0lxGtUF
UyWW4WA3/SnYKsy5Iy4rORhKrQ0RpcEMpOtxiy3YSes0aSD8aayY5AjK3DMIjL1/
JgyM/Tn2mBDwpsh+RO/B1Va7yUC9/m6mOdI6cxLd8pRjLPlyU22dUZD7YAd2mSLt
n5x+mFS9C2v8LwK/Xo2NZL1PlYpPnNKbWRxxCY9A2RZuSZZGQ+P112rN1NeQoTd7
pRkBY1qrAeE6BqCK08lYA+g37E2JBVUO4IGhsEh87xEzujeMk3k+dw2ZMrU5OBPu
rShL0JBar4F+7zNOZYeBSyrKVvtOWFxyZbTQaSqlHDD1gzt0WdvmB52jkYsz4QGl
H1dawXtauGGN9h6nzoW5HrQk6eD+PRcCG+iQFJtGmuF2L5Z2/l5Zv+k5cbhfyVE8
`protect END_PROTECTED
