`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQSAfFJtpuLwfDbJtXjvFNLJ+E8c/osRfuakOinH3vsu1JiLDkkEpO/u0i2qk9rx
CWCWjGWCUKUaOS8o1hwMRxKeLqf8axImVtzFz4F3HYYjYB+SIL58ake6XJI3w85E
HAmXxjYxOdtk01ftuvwUZJ3DKQvKNL3F1ypEIKRYcF/FKnAy+t7fS1cEcIr9ZMS1
IqdR5aDuJjLwFkMM7tYm2tgx2lOH44xcF+MmCcnFPemMKVf+ScLQu6dckg9Un81U
+Zr55synthHkFXkc2rUGJ12lALzuhyOns1BtV7HdeeuU/h8LKni9wOwF2EbXLNLQ
V4kcGMVz73NMm1eMtoW0c+bPyaDZSiGY1oQ85hGk+TueDo7Azffofghv6xxUJRY7
q0aUiYonEhsTG5pYIL+j56uQ6K1eeW3rSVL2QyyVz5M24Ncur3lvaA3/hgDKSIUU
Pmqyv5cQBznmvRriPjTYmSeZ2DE0hSExvxjiY7IoCbeCQHzsaXzwu/RCMJAM/sV3
EvIlscqdPINXVwJS/9fwJlaUFNk5iHyi9GqEhUhkN7cuUM4b0odZ172wmzEqvcCq
moEdDkpYkfn4se5yN2BSSqWiGLJdFQZ6MFlwRgQKPKaN85gnAKQgYTPxXo7pwxgd
Yr58ZAG2I4kgWicJPgPo596RN9AZwglVEw/DlDxy6fbo0htuXIdQk9sVnq2psOYp
cCzvzVskdsmoZDOInCX2ixYPQrWEH9kbgIGLzAmvTBINSlBtU9RxnX3rddrE4CUz
UVlUDRl+ai6BlutrigdPhrXuUo2LPfnHiRaMNopwi0nsnXYL2gweZN5htZpPJQ6W
3a/QTdLjPH+op829RVQmgjjG/tnTxzJSSTOgh71wfB1vNJKbHJMElKNdaWsoQFGg
JsHdcaly3wcWbZ1upZ18CL4LZTi4bhHFBl6aXgwbf665Ly5GgJMCee3vXR5VroX9
gX7OV1E5i74MwO0dl0fqzSsTtB7VxUTtULyGF8mqqWxsJcqsDhnUuWaqhJpa1u6D
nzRrUe4jynn3RELxLGXV/uwuU6Vh7MMKzprX5e3jn3KVwrkZyGyPyWRAY5geLpVp
7lPJ9dxfUmlYcCywuhhlqrv0zYn4+KYM/YCgfgXkc1LuQjrKwwZk/jloJrXxcVVn
K33BWS4Coy9rVjxCzVSbmrOlJSCe5BMkobR96pOmtJDYv3biJOUQobCcnDxcXpOy
62gKzGlBU4C112WE2i6+6l9o9ab1qdzx2qXl4DgBYzNhtwBt2hybXjPDQ5EJBZe4
tBMBFlL05BRt7ek5+Iv790g7/TSbEAqSQq64/qYLNDCz5fzGpJ5p2AwdEacm9isH
xN7M0HHYUa4BuXec3Iq+H+TqlMBcNHVn543MiTquss8Xjb32OL1G/xr5OJCx539Z
3NFT98kYDkUaEuuDOvfittlf3X31qZ/0aGoSqPcerRzp90Ck+SjtIltHarFi7bh5
sXmDXBXlt/OhC4Cqyl2Fx72LGLDwbshz+8h/RV36c5VmdvKSejSlMkUIgvzUDHx/
trr01D2wjwDqWO+vafLTP2ESHz02pVWj61lVmJmLqJemWVamkdDxpGRTeeXnC/cc
cnmNyKazPb5GoFPVpPMfN5eLkEFspF13R9iAChKnMdLoMIdPQzSzemBpjeOKnbtz
90pWLhcgv0w4hGjI3cOPQG6yiNXAroFN312bB7bfGi+QkkgRLA0OjuWFeMEx59mE
fexHihOK8OBKKTLbIGjUDNRIAcLO8qF+S1wTrFlkfxLSoRHRylinczzReiMyhBuI
7twzpY4Srp7uvVPKNVGVvlwqJf/zDndNz/uJ4zrXwdyqD45L5Sial051A9y0r+au
OrgGmlpwgrKk/x6d9jqXaaDF4pjvctlguY2YJzGTUQJvj1wEdyrRQ7NKGf/80X/S
TTIARXvRB8prqMWqrSSdcF6pGYqpgEuPkX/opAuWM/mJG/+Olt+C0kIi4YIVElTg
jIoRuDx+2ZuuIPlLfjxK8mCApD8wS/qk0vrufMxEEeboqVZ6o0H9zPiRWWmE4ClU
Ck2ZvxiF+duUN6BBonAuxUSCLxUwm6IHAhqq9+ajg7Gm3hkf3adUDt1q6bG/fXMo
1194aVzPBsWpwlin2UDVm8tM3CNSJYuuNH2WAvTpjIW9HgMKjtJYWcuL+Tbj+ZEG
sQFxpr3sRQjZ6avBzvF1asHK0PuTQ+o6EyfwBHIOnxSzmbMRcvZVirVa4X9RN4gQ
MspDqIIqcTxB8IQtcyzAOW9ZVjVMEmYLhO6MYwGjZUTUkq+gOyx1gyF81zMrSkZP
goxM28t1bbGLNkWLQqsitA==
`protect END_PROTECTED
