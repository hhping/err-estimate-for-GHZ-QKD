`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15i7sG8xJ3ACbLOg0vDePblWx0dK0E/61gvmde7YTLTSOTwtlFvvjAEKT4Z/4k2+
b/UxChIl9Za4iRkVTq6cQ52F1kTIllwVRfnVEyaHGeSreSpF+S/+8CC/FfuBImfj
XLRZ34df628RYjmL2IjERblTB+jZcdFu4QAdVH9e4aHsfTVTHjs5I+AJjmiAXZoD
TWUJnjLvudTAPTDRIYt5TBTYlbtpwhdfvBwODXMgb7iSw9sHOKDk4BB7IsY6ZRvD
jedB7Byt0Z4bIwmDK+06ZdHWJcTynHwU57lVLTz7rryxbyegI8i1YmyT8Csa8sI5
50xddq1DUxB4qosOs6pJgt0XhOsNGvOZ6pVfuV8W2VHs6KuNLLSzYaBi3mgSYlk9
MeNW5WBAlfwKfSr7XuAjFU2/Mrk3UYofmNqeG3sHr0QFLlQickfEWN/ruzZvXqMl
m+O84N2aQ433LkKzu5c9LP/d7Hfn3TVMu8H7ApZjaJ32RvUixX36kYwWX8my1q4s
1QjaRlaAI3K8QZhdLSFDlwVxqPCSrl+SGnzgmenJKwZ4qzovvRslibS0pDHxBXik
cM4rTDV1g2XuFwQAg5yppXCVTwl/YSZEN+XuDJdZZY3d2tOpmRqh/fSlMctAILEs
ylBWTLhn5Ilr90FBWqPecsxh5CRI7y3zmure2upGyHxUO6riqhe9+JZJfGdATOXT
cLAbd/2Ud+hhM2zLZ/td2G7T53ik5ug+6pqMwgmTwKi6u2kGRqwbq1AWturzRJYQ
vxMhCPwOsdESDpvgTecHNpfFG+2QAv8ypbBLnZ2GyTzZzPZtoSPk0Gk6ZoaKQtG0
3YkI74pXL0AxyzvhEVhQVHX2xopGbQ4VMN/lsl5YfVNyuW0a33aYMuiWPnIk6Myx
1rSOCggmK2jVeXmXkFjqvjFSR3D936To0bVfYSemjdyei51AOztcBXyygxJBxkJ2
8q9BRM/aVmXigFIWS/2ufndNIa0Qcdjx3q+YVz5sSv6zNkQMxfojvA1Ajw9iggW+
lP/ajZJQ9YVucvHwHqp+7tEYVRwJEIihoPLLjKYV/HDKP81OPY9lcG35HyZIZU1d
AU/L/Izo+GAMj7sX5Zd7B6XM3RtuKZK8sJGWm1Yv1AipykKCukKarb5rgqo9mrSV
4Y2y2StKa+uCviE0ScYMjrltVMrFdpYwgYDutJyENRqJPal6codSMwQyJsifRLyH
SN/hIn+9UFhtKZY+yWj/TyZkBFEUnhmdVQU2fqUYmSk65JTuPfHH2q/IL2E93XRX
D2Wd17SQPgve8/qvBmAB1U//FlwcZqH6+8OaYwTTgSNsadmnYHyvgiceOlGganat
U1oKNHsX+mp5VEjiCFPqP457fjZ2qIr3ZoqV6Rt3NM/hjc8UgzrreRaIYVclC58f
XJLRo3ZgAOeYqIdFJLGdQH/gLcEq76XdMH+3Vdxhnrulu3sFIIzjJzBTrcxck/Em
YM9u7WOxjFlH4UKj1qb2gzFJnkpMjKA+4ZJaCOYsb2GL2fRvT84Lqnpp6sq69Ocr
H2/nl06pbKYuEhkeHOlljektL8cbeRDogjfTpJXGoAS+8RE/6ADnDh6rtteI4JXy
uOkZAEKtBJU4gNs2f9Hglq2nkvJiulmWENyoX6lxZhIH8cEhxhq/voHXLNAE0UBf
nKbmORZlnSsl2PUtGpnKA/tjLpM0w1g0SZlq//tMyaX5PDfUtC2wE4nvkIlt7CON
DW5vl0EW95S/Jmvw3TbZ8vsIpWDCXhQIIl5gKDwkAE0hSucLjRTo18ls3FfW9FK+
cA0wHrgHh+e2zThFnMFJpRgbkpvQBi2T25Nm/9VA7sqCebG1Hmo/B0GdeX5UE8Ex
cvdoVCDSxIOJCsIzt9OkNkh4LOEzthYLFVHMmhZajZSAEyqjJttYgfYZY3g5dICl
e51qr9VCyo9as4EOvqbezKij9G9Vdfqkme1L9U8THVH1G9HSJtJw5ovMb9CsdQXk
hXj+ceBiyxt+aNgI6Z56T5HkKlkp5ojLUYjPoOZkPoJOpOXDmSs4G9TPxGj8+E53
V+AnjLI6UlwuIKnWvxACv9+Nqui79FsbQ2+7HGRk6AkK6lJVT2/6E+nLlr4Ek17i
c4LE89Pe9Kf2RFL0x4sZ9xTjkd6jVHtScYsCnBVHm3fQ/cHDpWZi9Zv36ckJVLUg
tX2yQZ/OR0wHgBSDIjXTlSZ1MiJUGSBXi+K1IoKZoCFC7QTQ/VjCJIB4GODK4dEg
yJtvgDXSAaiZ8sFxhB0wpmE0T5OX6KXM8QcFxFQZHhOUjxs0KXTa92+tX3p3dzhw
ecgc0IzUPb+OfPYQMroRb7jQ8N0Y2mp8y3AyM/c6jsg=
`protect END_PROTECTED
