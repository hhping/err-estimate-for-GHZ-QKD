`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0fQ88vyQfw87NyW1qTKWrqln/r2iadqDcPbeZ6gvOv0hsW8hEEE5cOg578oX/bA
4tMX8AybMNLPvxoC2AoyLa2zJwfNYHKBwmWLwYuNkCWVFY0ghkxSpsOa2Xaci3lG
6NnXiOmUVt+qdkuja6MDqGaJgrCSRQ18+7FuB5QqeArgByLYfQYltJNmVASJ+ubL
Cb4Ya6kDkCEiA0XeloKJ6mHYKsBnqqaV2IKCCPIvlFDpRLS0dXPkRP0TpHgSP2WB
NCCruTXZvFHn2xkhqCKPKOncnRokmmdiYdYeIXVIxiEFIgmhoKde0gbcFmSH26Fh
6XMQNygEO+L1nmGhwPyaxJUyDwnX4qzK49Mbg4xwLPpFpqP2wHHc6iYXNz31Pp3m
`protect END_PROTECTED
