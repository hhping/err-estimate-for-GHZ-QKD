`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/HY48hPbssT4HZRUkidYNBnK+KD6PL+3AcBROY3NJoagND6isn9+dI/HdvOR+XAs
Hb5YHaIpVDfC9qQLWI0oRUJcZBF44pjn7Rbkpe85bsh1cGptkQJxcseU8sX2k7xR
tH8BlxluMRZnQKrDnupzKWfsvcOWt9H5v/MbWJErukgsNYJy1dLS2el27aGiLclB
JCXSBS7j+1CR60PrOQxJVWIBnvBB3I2HW362Wi8KWrQj55GHINk4WTN37Thx9F2o
I7lSsZ5ZOIii3Prx6W/FMauX1gXL95XoBMI74M+0SdnN3plPsCJT9lUHfEIru4y0
9UDi85daEWneWrSn9eAASPrRiysc8qJVQlP91w1RGI++/zUix2LFWWafazBkhn2R
X5Mu4umoZ3a8Ir8T+tDGXv/iRLZedmvPWEMXQbD1G/RDw4JrtxIw5BprE6X5YFLg
evkZBmj8LK38XTGvpT55BBd+p14CzDY7SVasRESwQpF76d+iFxCJkGf+8u+lrJRi
eR4F71KLmeKG9Kj1wcb3jltpEEHRRvXVTSQU8dcdka7KUutsng+SNCrNgo1f1pJJ
5bZt+swS9oEuZTHcxZTPej9HzU9HT7o/LeLC8tdCt+0=
`protect END_PROTECTED
