`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfyEqd3ufj15OE7QVAqP29n81hnCutjs7MY9btor6AthI5NZZVTvoFvsGAhmzPMI
BCLuNuRdyZyUp+uzoDODiq5tpxCaTxJB3X0zBF2J9GUN/SCyvombiVyv+GeCBeHE
UmZrumN7oCl/laxb4t8VnJQgB3lxgdbv9rwPVLzPCNliDEA/by1V6KtVpBPyBQLW
b7uAF0SoYkv/bQRO/+XZY9tHERL5bN8h+0Z96UwhUp03EOv2Fs9Z6WBqSxUDsQLb
n/TW5Vaz2vrFThv39/1wVbS2Ky6jp7znLBQzAqZqSQibDez6Z+T5VvmDG2axiUxz
VXlvyremGuuRlfKtW98KEdrueMDOs6d1hJNugx7MTOAq2lGzkjs+Goro00Zw0iac
J12TbNdGHd+bXXDaKa+UUDadFli9ibH4zZrfYDLCVD+Dxk+qKbU68QsGQwHQ9vsG
bEbTWEPraimT/e+W/5c05XukDprRQGVZtkHWpiU5zrwjVwMguj2L6n2Kl5ydgWpJ
UYRChMNGwaVdykJoKf2ViVq5rc8G15BEIB6tYr6AS0Psg/2LQwG4zZljyyfP/v4y
hFGt3wG6PB3EQCfKFmC/UHkYle79CczQ+jwJIaUiiDkoN+wsoJgRtjI7gFFvSLm1
UV3x6UJ/nEfLSOL7r79hz5hnVYMU4tWXg5SYW+IhblGUCSSuJA5MmB4ubvyf+H+n
xx9kDujOS6tzX1VLXpzFLgbvTbc1As5Bj2hP2/iH8ItviM3lv7eG2bfQxsC8ewBe
3ql5N3Qv/lkwnCZl/8K8FCcAv4TMdT8ZauZJ3CbaLETUamCOH0ydUcWwHnCtR9K8
6pNzUPoSjOFUkcleYieJyWKsHUI2n8PtksLORs4aHU9QsuM1xbTK+fsXmBjkBlny
LhgxStKJOzVDO3pGigOOtG8cmUJ6VfREkPjY20VWCZhtvSH5fLbSSor0Pp/tahJM
3GD5owdg0tEMftcWs2pMRn1/BwTnF698jGcJzD9u0b6cn4byYj2+OBar5opLr2Cz
I8XaTlOb/b1SN5ICo/NaV+LZgoWqJzvchLc2U7r5Qzsm2IkcOpMTQM4NBrnWvwA9
amXxFfVXyaT9sT4yw90IGG1hwqDCsw40b0ekDstoyagbBJvORdePSl/Sj8j1+MZd
FR+u3QVzqn2TpCoG9pfa/XHyguyXceMfE6moY6Ofdsbhu4v+obieebSpceqS18v5
4wLziqMpeuuFyBW+oR2Wxkj3KtpKOujMojUGxi5kv6IZsSlmU5Ak9TIKv3bKuXrw
lyqvKmLuTEuMaK9CQHj98jLW+lHdhGte5mquqbOpB+7NoJs5hCZ0N5uS9ErodtEj
bIjs9tV/rXk0khzNOuqgkplhEUROzMuyR4rdntYrYqXgdsULiRGxoCuW50PFrs+C
e4GBFdToy+M1SPXVnf69VyK1ZfQElnYJ3uD274g2JDPZLAFp5/33Z7h0+gQuMFct
QXWI/8cazWaAL7IMaYZao923M1YkSTDhk5lTAbTw3Ims759CCjnRXVP7KP75eTUP
72WaNe2fE+aUVVeFuqG4fr6qxpdqAAgiqP8JKLdBydNv7kNq66D2Jaq6ua3NuL7T
CnTkSSh0AUH3KLxNq1sxIvNq/zkjsJpWXS12fgT2A/z1DrRNaqjXNGy54/W0vleB
IhFug/pFGWB1NjIn1REfg36uWpi6xkGGvt7qFik0KWV9ratu0fSqyjkWyuIMOu4D
nFunwdpf/Ic9Ld+C/nSPSZ9XEqaRTKvYSZTreXmjNzYbTyDwIkgs9ma9fCiA9vDI
I1AeokpDdKGSYkVYV88S6dDooAqJFrnjyppndwfE+b4AYbYWWL8smhmF/KXFShF5
qQ6RfENMjK1kiIbc3hgp+yMgcrBBLy8zHCJDRbnVcl/l8maODQD7nVoDeCd/hWRT
XGP9QyhH+96A5VCzow+Cs7wdfDG/WKbarUeMAPhtYSF+o3HgxDFaUwiuQhG0Tule
Hj5JnXsJvp5SDrgigGZ/yGhg7ljcHgk17Mx/DymECKc4rHYMTucK6wOyEfSfpneg
gTF3/W+ZZZoyiN/GsPZlN4ZC5omiWO+e6V1TRuHg4Oj35ne+F5w64Ie97XTchvt/
7YOJ7U/2v+MtnEHD7pzb7xGX2GqMW+8I+dljL9P1sfwsRcqqfvFzLaGSwqlz2Xjr
7LRVeCbo9naq5ZdiD8Qk3XSCbg2Ba9SJd6gpIKcW87OX6A0M/ie7ZhipMLAx7I5Y
j9mJKRotwASJdPWERCOnR4Mwqdr5cUcm3/zTwGpJxVt5m2Agm0uvOLxIWtw7TEiS
bTy8HqYmbJ4vANILBVW1RvIuh0tCvO4x1PTSeqaZ2gTnUjYLaGeSYIRl0J9lrCnO
COVIMvfa3y2Ak10Hg7gr/GRtQIvgRKxp47Xh56yFVEr89qPNt5ApZcy4wq9yzNb8
cgM4szN0drgPCKq0Zr6tfI8kuPPVIWVzNkZzh6QIGCXg9gGGEmLr+qqioIeHSO+Y
TEbwEKT6Qar22vxDohiDSIbULdGcF5v6VpwbRcgIe0zz+HKHjdrIKS0scVjchxnc
+s//rlULAR2mSkoE2oKyCBbJ6ZTMCzQrdvSKUFasPYPKQgUtuyQcJ27AoToJ0GAp
h68BR4UBL9InXJWCc9chyBEklDeCX8+CUk5mU678GH5qoYdhPVief+hpYELRqxGM
Yxlaoe2sxpaGFvYpmG9TmSj3PU6HWg8yYpeykq++IhENKNP4loOgpOelKOBsH48Y
5kU3tU3yAIya9qpBtzWjXf0xfY8mzfpRuT834OZBXAyVYB+fyk+qYMLUQ/54M+pY
u3su4GJpjFrTFytWDRzvm8y9uMi1t2GBorHBc1eXQTOaNdlVhM+O/1MQGhdXw8uk
fMzwFcoQw1wBU7y2Dqt9qQ==
`protect END_PROTECTED
