`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovHs37n2tvTir8C3HOa9nvZ30CH1CdurVE166Vzj36tuwSpLtn+n1TeqhlkDPwas
J6aDJIYXqMlDDbK5jaNcLDt2i+E6OLou/m0A+uMry5nCUIBR01IanOeo4ER7qw9t
1Fnll9YpCPi5ylv1jThjrrXYpmn5b7928CdehEtA5Sb164OaFFybO/FmDksmOl4f
QOGjNiLp5u0oSVBsd+7RiTsAdfyHLIzp01RPOFKaW9Q=
`protect END_PROTECTED
