`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHoYURRGZf6RPAi7tU2iiEblOveB426GGuHBvfL+5iYK7q3+ikRIx6+019KTrqht
9yTRkSlJdtalXp6T/sroooGNcal+u1Yb+QUgNjhPw1MmS+TgXwFwVM5vA18Rlj0c
aItBwbj9nPgXKr8VZ9oAoJqXSOybKluMK+3HV+/QK94iFDP8vXrkHRBv09sByDW1
wFQIvR+6shbvNFqDBZSMSHDLEk02U8tQywLDiRfGpns3HNpZdBC8AfhRgVklWzc5
jVq0RQghc+NaBkeZJI8Nc3kxLFhB4m9u+6vOYc+attfKCnckPN7YUssFsecG05gr
qOuoc6IlGqRd3aITBcqYYKbI14g+JDnfV7UX9Bp3g8xjZi4jogWUV4jyiTggc04O
gGHWqaCc8jfAuzDSXdYZ5qlPy8tP5zRbAZ6mUVTZQaXICa/N6fSVTacDsjOO0ytV
LOML4GIPcEr1Fzs2JQKmK7N28XIfTTd/9czc/txLqdSGBvTNYV1TTsgJt81+Dlcy
AR/Y846y2V08Swahw4tH4yV/P6x7l7o7zMYisQHUaMLVcwFYOtrqM2h0KYjyVpXY
I821QrtL8GFr6DzEsbu5/rHgRhlfqm3K0qEwcvluPQ1JTedIF1ItPQTpAn/UnU4G
mWkmrj3chgzR82wVr+kBW2x44IdlhI6NYbK3Td0GSL66eF63StbxHFOPNNGr8q1k
wCNar0dc75C2uUigQZ955xAPPw2mVuwpERAIKYr7gkCobPj6pVJ+umydVT/DDlAL
5/llrN/vqohXUPfwv+TQs8Mt4M3k0Kv+AI6sMhqs1SGoU2g75tX/NyS+eMjbbmPJ
tMPD9em8u6epEHKtCcmDs9byOTmHHRjP4YcDsT5eVLDGhekeis1v+W7HApb9jSiN
JEFWnoi8UsUlWJiDoA5T7hDsgATn5dt2N0dZdIoe/x1vQMG+xjrOq3KSMHt7erC9
wYGqnExsdRLz25pb5K/aCzPUSacSzy8clmpQ/R41srH2zR1VvbAExcc2iKeqgwfT
wuvSNdE3Tx0DIqLl0kVj41kajvQLjCru6tmnzMo34Ws05JHQ20flIc2IBOeQJUtL
iKoHdNdsw85XUetqxOfI81wcysm3OIzuhS0QFRJhyCcS3v96CYYqFyImLIOlhVxz
SpZukeCuTeDntLxAP6jWYEL8D8zxCEfuA+6UqFLbVQGddNHmEjivFAGNbwhhuYOy
8/CowSMDsb2hkQUt/KSLdhgnsBmAB8DqtDGS2rXxiE/uHBZ1kR/gMRGN5//jA3bc
caUUMc7vFiKVElJmvhWStlgaprFYmcQkm668+P1VLtHpZOnVodjTwotKL0AkUJHU
FNuV2GRvjSiFEGTvPnq0OYwbjBL8C0HsRnBlLp2pLw2ERXjVQ6GRfQrqCDdQUMMi
y5TmArb6Itg8DwEElTK0opwBQK7NnsGHs6b2+4L2l6TdDDBe+k2XHe0SBV6ED7o5
XOh1kxwcQAzfZJrh79d45Rcj9Ttx81iA270SHDHwrET8VAtBHqsLUBzxWugJl1z3
K+H0izydfjuGqLIhLz6FFK9p4hGFe8l+ZbAEpLgXnEb4fx4PZboAM7BJ+53Dkns+
3irevLH9Ggil6IKaK9d8KFgk8h8msfBQ8O3++58TZmfNMNQOlWgUdG88hGrmPFoB
9ngt5DzJeHep0VBgCZgdUCD0h6vybKYU5GD0lsnGXzcfpBnmM6SMNw+i2NxkoguO
ZApAn2Y4SdSd3bkrw10mznGPDDPOqCJp2PuS7rMALLdy7+vg3IlWA5FDjJm75ks8
EDH83gODpHxL2GQDNBgPe/7zbNizStD79EhhDxAdQYO9264BBxmoGe1YCGX5620m
tP2XYlELElsRHI+2CwxVLwcivzdH8Rd56x8T/BKZV8ucbMJyFiGipDQBmPs9xXJ3
A4tFStkqqDVK8/ni1czVXc5HmxajCs+lzHrihPr0Goq3zQZbqzPmMRwdvFivV8Sk
lEQ4OFSg69zLW0oLt6ibwYj/VvCEzjbi9W8Tb8K9wQq6ydbIoLRwn2Kkr7C75mOt
eXMStLrW9/Lpbz8Ik0oruE6+iiMHH53rccQnUUsLjSceEVYVlc1SPjhNhYRoNMJK
XcLEbYSqEFLZLiBUhQXBw6IK+QKdA9EDzB69hBzswl/8L05fgCQDq80J6LenE9b3
ZMt4bog4ZWjQeR6VE42Lu12ZWw+Q1DEJT10VzJMAhM680loI3/haPjVFnM/FE9p0
eM+apj7mdJVX3l7oG6RG2HOSUWixgYBqz5PNdWyw62dLqwkoYhkUfcvsanCi98zs
H+Ee85PPFbbzDxCOsJfauw0Ft4k11pX0IsNDUjijjgXBiOOvl0Ntq+i2d9DbnzhF
R5LFGQFmRoih5gThtAkmnlRSQsw/OJVHgZNcsDyFywFv1KydYKbluPw8pyChd7MW
wQkVcZUYsfjNW4qbb/xtCuUvrhToOigNZ2IHkNg2Uw3eC0aDjQHfL1nlo7es5R17
k+FsFYx8Jc1N0ymfZmmt0NtWpAIaw0C7pyuNOQQWX+TtPYG27Qp1BrkPjcb8Edho
E9+HvyU5sayBW1PaxekdGli52kcWRBs1VlAfpEZuoyhesQ8HzwOOMz9dBFtUzVx9
olhaD7Czkk+qwylFYqu4rtBDxA16tgDhUbc4aiHBy8aJDix+Akh5Je2daSPvLKKu
gk1vcgFuHsT4Euy77wAq9OxpGqEgxNDMjaH4qQn7l98L2Ju4fMpUgh/GaOmIAW9m
iw3abCC8YouaMSP3Gm/P6j4V8oV1j+62YwMwc5M42hKbIe+C7Egbi8y5zCG+N9CL
ytVSBFMebnxHQNNeG2YoduihxoXGyH5BXmUtBplM0xDzBcI8ssYoNWxtmBMMXrmY
C530Ja1eTvMoH1t4AisUosFG+rNgdXAKAR+ruJ6W+ynmDZtobY7qtwTlMjZ/B/Cz
uQTTpKlLIUhUnPh5GSId+uX+zfbj7a5Y8BP37EOEVn2YXRC43yt2aBx8HTF9Z4O0
rlFHf+bilqUAdrkm6wv9U6mQDkSWYEGI9gOwC54fbxqJ7iHDzGMHnxXAd9Z2eMFV
3B8Q6yYLL9jqKjPLTkpSAxO4bPY0HNbLD3LrJ+WDmPBFREaSuPG4oH+Jc/7Eugvu
3dXh2EwA8qOM7YdJosyQdsqcWsiI0t/pqIl7f1IpYoh+gutwTbyo3NXUqtxvvOB+
MrL4ptXiFGli2oMZFVjic4GWcpiOKYVXtCg51yEMIBoT1lFcUZTxK9Xvh9qI4KYU
SINE5w6Dc2xrospnmDTLoZ2jdWImShF7Q5KhMCpJuUJxEZ/evGK34ERkV8ESiZXi
L5uB2a292ZDOnjvcoxqAG+16DzSItX8j5rZLO+YKd0aiOpHDI3XWsHl/BY++sDU4
QB4Bhr9NjqIsUslL65FbCQ==
`protect END_PROTECTED
