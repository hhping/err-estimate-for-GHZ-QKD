`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogZtbVx6DxzYpb2z+RPFJQEDDPA7U3IrRRNkmrpG5z7XVLtpiuLt3je7k+14wpns
eEOAkgt47IN5EncSMq8SVcAn2t+4BQxJNHPa8TNdV9kGunif50xdKps95Z5rj+Tr
SY+nx25KXnGqO/FK18BY9M+crs75BUFsKtfFyKZaL3bVkH74i+oFvFFA8GhNwgwB
vcWw3kyGja+s7gNMeQ5/v2AKFMpWJaIA8nGLwZesTX+Jlkd4R3IyUYzbEDSu+zcD
/qpLij6VQphTWVW38orX68/A85Yu5cdbL/F2bso++LoWwBf6KsAG3u6Jfpg2zHPP
tYb5booOPEygmDqrFkwbXTdFEB/PJEg07HPCjj69TLJ+jK+cduJha41+7JenA0rY
jKRC6rsha8Vupy7BSGD52gV+YOBn7eDySsdQD8IqG/BbhX2ZPeqMWmDI4fqivvgh
xo3TwHP1W/UHOn3Bdznjgu3ZOBcxqYgp14m/94ImU320VUOic9qO7vT0j12zOX3/
syuFtpoqz66sZ2pPWVSK3t6eKYWZ474X5gIxH1gVUJg78ymyphpY/Mw5/ytowax3
2igkmLwI+rpAAFuuprtpNpR4E5IQE9SQx1zEbyjGEefp+v5pYlezs826gUTIXfC3
4HNxKMYU9JRRxQqW01u6eJe8fuljMYcAgUhBGABYNskOpiDkylGQB3PXIQVlb5bI
qhzk66gsob3whoYNHk1hzw98uoorXhQXP38aLqndVWKosXgqeNs+8/np6QN8xOs3
IcXYMJyKRE5zWqyv7rEvHvefIvcy9WZ8hd5Cy/tVyj97OOc/6j1vidn5w6IcTszf
mpBiPKKfzGPJ0N8hsry5mg==
`protect END_PROTECTED
