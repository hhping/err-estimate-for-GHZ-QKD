`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hnxzBxZddjh8TEKpQdZ4cf9ovtsaghE++TbH72rjQQhk7Ae66XKPUDmrLbEvF/r8
VpG+6n2p5Vj16eaAOgG5X6KObpZXM5ZV2Yrk2ziA6ny0b4hC+ueU+CoUZJMPS+a8
+ftLt0uXbNlbMb/Xh2HC4hel1aZYkugXpVTI5RDp37XqkMf/ZzIKo+4qXVoFIvOh
TL0HOaIcX80RX+QqPQ+xKMxWZSivvVhFeo/lIZ+ewykhSQZUWJp9nH+U68fa/tJ/
NMaJkT1VgRtu6F+wiRjIGsLJnfwZvjCkgEq6QcDogHT2CTZ0xAEW0vv2hVS0Rgrp
+BlL9DJNO2zOUWl5IaRsKOaHfoBBP7GONG3JaqJp5ryzNZVUCea727Itydq9JSiJ
sBpJiU8j2+gev851ZG4pXyNUvI+D95olgfBdhpFxMaRkg7XGYKGS/KauKmwNlnON
ewWBhXWQNqLF6nn19E1HuC3tlBuSgHMaE7VeLnpXSuOZ8lPQKkODVkpj5eaR5FLP
Xlv5dPvNF49yvTaj6HVh5HN3hH/R/qxeY89xD1nAgi2QEi8I/SuCA1axRMetvJYo
8QaT9WrYga572u74GcX43PN3CEGAFWJFMDNvTfvHVfdW2z7Mb7yjiKVzczV7gQLi
eTqx4+La3NnIx44QjLRSQDbQgSflHptXBFPn9gJtVWkOqoKuPpvYhtb5xXk+lVWs
gK/N+DSVa33cioftKrhzzd0rkaL1H44poNgzmorajrJx982Ea8W9YcPv+U6KOvwM
Qq1euaQsFXNTu6Hhe7DDy/ICIE0EfhUUH4fTN3BqvJPgspVVfAHaMvEqb/Yol6TO
133rRmBRNp7a5mQ9CL1M9HTx/4ZnseErKJMe9arod0QB1uPU7XO3vNHN0oT2KgTb
Tk8WRxOctxYNH+78CnCcb8q4ba6OV4lxwCJp1N/FnnNy8bw0VdlCQTKEp4Ot7nf9
GitY85jTOJqahCAvbpc4ggJi6leIBTwACp36gFC+Z2QXvOP1PdUDi1HF8jbWQHlF
CqfUYEqYEqpCUML7UYbloAwYZASZazznYEyyRJ+6o7HXbogQKLtQK28MHDh6hX0I
iFLo4sOFglXkvae1yEGC1jguU8LTfMNkkJfc+jZ0lyF+68aUtf5As/asR8ciSmzr
SpY8uxzkqcWjRX2NXZPF+UKsSMFmK7lLnnGhjjPCicQLwhzWDVH6ZC9XSvqb29zD
hsUqn9Yre9EWaSSN3Nc97T0RA4+S6h6IcG19CPP0pflV5yQ5koBvvy3vJzzp+PFX
bGc17C/3HXuiqlPPyGeHEujqNrJ6uBIXcUUIjKsjjNd86dIix09s3ToDZzcUSCjq
P7dxuEoAB72eG+I6jfTJbFyaK5bL9htwTH9/+p4esk0aXGgAoNaZH9/XVD8LlQkn
Z9ihDHgaEt9lvDCpdUYw2jHeGyMbG+rAsQkEHJjEi4wAHY9ikJnGucaKVjCr7T6b
VKPc2uupLH6coOCxSPbfFJkrCflA4l3dPoVafmn4YJ6v8YG/n+u9NPb+Lya2dmTW
9ZSllsrvEp3U74zaGbNjXAzNM9NEuEsaewW/tQPPSSv4A+1u13kCu3UpAUlmyo5k
Wo9l+HfDNIBvSrQOTMZaaKzlDepKUaSxTHteAx8L7DatKZa8DPzCm+XneLghUgKc
JcCkYGK1elfPp/046X/rYjXYCDJxXBwaqhDa8Q6zTkFdYXldduir2ktW+1OSLNSc
W55QEK1NrxYMriDjLnLpGKcLVEcsmnU/IqjrU/nLzZUnUDZahqheLnOwJW8mkiit
QA1G6DAb7bwT/lfDssQTezKymTdrRhMDSf40Gf1h69NOcB9GPiO5sLWwig5li0yu
W2KtFq1H6inf2m+bycPTDKHYs5bLjKXQIucffeVqL2mNu36AUsHE3RkTNwKAt67D
XJM1MM5GdyrwgK8wN89ROqqhePXqyQNGYxDtBglTujT37P/FVcidpYWFFuZRVw8R
yRw28CPOR1oERu/pJOCMSIsVNiGh05fup4DnbnNyZZdQ5fphs/2UsevKTfPUy0Kz
a901GAV/+811s/ted9zOoQ==
`protect END_PROTECTED
