`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pnYGHdwv4+7byEx3D6i351XAe1hLOkV6etP+BeZihdvG7wcJarAokk+SQUQMJEFR
CIIYNnFEYmo9TQTZJEQXptx9inCBSsuhZbSDHYNRHVDCPK5gZI8cPVVjjTHiwIVF
uhm6yzrMtndCTle/F9y3oef6ly40upTrNrREwVv10gDtGc2mzbR0M7AvBaX8TFEu
n15e0R2bi6kQxR9bR+ArjqbApSxmBBeVlQmw+QzH5cA5tEt3J80s4CwQki2KuuTd
V+MAb8EnAbioYc3wMVRWtUmzUP7wWcZN58xvYKo5zd1KooDhPnpu91B2cANFJ/qR
AyzlBQnGpTxOUg6tG7BY58NSSCmJyV6cYAVR1dGaXPDbcXtbICVpXxnXyqIwMmF+
pS1aln+84ypVpqiOn+GPZTyVIPiNkaSLdPOkyAbBVXqpbqEtq7kMWGHsvOuK4RQb
3ZWfhNF0pPAVjbVWWXZ53cjYCZOaTOiCvstKU7J5illyKtY44xSrMEmt/CunPebT
AlEylk0a/yJYsURCbzu138Pg/NueepGQGQ9+qWJg170s6earMhFAN1i8CcJB/kIu
Pkmk/tXBCHeEUWs25kq18wRChsZqqU1R3wd1dq0nJszjjm8v2HzqImN/1h8ZpVJc
H8/EppAif7RsgELjmzJiy0bHbbtNulAym3XZwe4vv0OMuXSfLG4rvnBK13eNk1oc
RSr9on7GeSoO4aIQ+CIj4U5LOCnDmOjiK53kN7LQznmWMMGSYr0V2c7R+24uQerY
M14XfTRdisHEGFeUaKDDGZOB0gAqINk9eOF/ilTKHv1H8qriwHyJV3jO37AYAiV4
2YoYuGL2JJW5PDAXPWVUj9r5Eh2tHjgBssXLyS8nG7lK8nGljuH0GOb8WJtqG2tD
kkRAjkJJmcsoPBDg+vMsnpJ6TY0Kz/WCIZyiFJixGKqTuI5yWgp55b7+nt5HZvx9
CTdUCBAlT6hWCfDYU3pplGk6yiwSKUJbOnz1ag5dRssQEZ0BaCQ33hpcAW5VhDBY
p5rLjRJsh5Ya2aoNqWLSTcfHqTW7hYxaBP3pvRyn7HYcBhdK0OksAndjJ7kF3v2t
SB7ULV7gEfHtEO5PYzdDxI3oqmlObqXnxQbQtSyyWfMv049Tz9LtR+IMI6ktz9gT
2pFY8XIDGpIPw/SBY0YSHQ==
`protect END_PROTECTED
