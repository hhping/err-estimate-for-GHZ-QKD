`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEK0jl/3UOC0+F6GzSmGHjrtchjOCVxniRLrGETeqB23wMNYVZCfhDqMIICIS8dS
fV9JqRtx/2HshZovbK/fv64Uuv3eGH3TYON5J430UIRjOHXLhGKE9+MjKHMmw/BO
5V1IjWuoTn6kyidiXWCnuOoFnp3mLyOLTBLUnp7J4CDAr5BET8Yyr8I25jqREESN
djRTDhTW4ja8HnVi2+Pf7xbubaAq/dC2eSmLc+srJ2mXeUV03G8DA9LxIqQQ71VP
Wb6znRXzUQfXdtuU9XgSKITod9CU6kf2zIqmivJwdIUSqvT/aUwDkOhioor4M8Jw
8AuKqfEy/BMvQC+6HZfDLDYbpJYnqBSs0wjNcz948WYWijfcLZwuLwj5/bt4Jqwy
wnLAxtQEeP9yOEgncihdZBj/JaxCYUIFkB6fUH0lha98MmvYWMS0VXlcP3VaKHVb
c2OqbMfe1YShjLx8KbMZyEAdS36eW5LRBlIp8x5QZELaj/6+lt0uKu5jdCpKdTWh
r+fH7Rb9+iLSMblRz95cUweRduAyBNIqG5RIA++x9HH4Sr2YZtwAs8cDMFz6d0l1
kMWDg5YcTSyiKuQkTLT0D9UeVDCuknaLXSuniXe0zyq6Tx963dXoF1dcpOSfTk+D
0ZWI6LHOlL9z5785gTwpjBCC0uJjYVVzWVvFR8K2zopI3Y5ck/uqwzi6lCvS2Gje
IF7YvqixHCP5iz8tO8vTzu2IDFcYlW7Umv9GGZ5AEv8wI+Ahdd95ybJ3lN14YOf+
SUJoziPFIusd6dVZPDgGfi2be3CMfMXtb+opOFvsmfLioOFG8Ekxvup/sH+pVr+5
3pKjVuO9EBIMfHxeZfqKZyfjhvLPOVYlUEbq+NPPXdkk66oKLNnE7WR6iyO36LkT
eUWYSiqUm05xK6aHpbOWyHlPoqkrELyx/OgR4MUzH3qBh2IY/e58CuijLWjrykT7
3vqEmQsYc+32I300vVel7w==
`protect END_PROTECTED
