`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AbzTgUaTDN8dWVCBon+bZjwqNWbwNzd5hPXsblMvvv5CmWdKYdpPl5ZMnCVEs0KK
P6O5iVPouf4ukFCV0NEE2UE3Dz/jC9JZt49n1NZryVfvqIYUrtz26zrOD8NFjnnQ
1H+TWKVJddK+lKVzjobNgcRWt4xOVl06mT6ynk9FK3NQL08F/LY2pES1uPdkERSm
CRLXUSrourGpZtbh2ye1abFPdHohlF171R9H6rkFx2UdMKud8lXXhNwNV3qIg5vO
ns0D9MPX81khK6WdJI3ir0n09ftUAFMyfSmawR85d5i9PeWFQWjVmyfLhKn4AQfI
u45ly5lES5NYaACOuYNuZJ8dWdbS3DTRwmtYcr35iehfHh9dlRzLgQ2vrup32Ctu
pUvrOYAMTnrxZ6BS1+SX6ZcENU7Q7cDQkc1ItVY+PS+JZ65EpnhW7upe5XS+23h/
HmcKOrfdELRJRAUgwWHtr2RMKbJ8aiIKor/4vJwEJkZwRup2d+GXv6K0MRTPx4Bz
O+6SkxWm5aKFZ4s+318+27XjorgHkN9O3cKU6WuOqRcrhYFcviMMWznSF3tGAgP5
BtgnuhT4349VNYcTiN//w7JUbtdlBRYe+VvJCP024LqSd/J2T0rKVJ3nhd7pRtNq
t8xZ/l4luQ0zxLomtCe6EUR8jq91VXoIZ8D3ABAnIwgAPpmB/sQ/PTFOx7IGYP/E
RLuHAjoK4SlSXrsQALA92dU/BnipOsTUMDUQ9GnfrPs=
`protect END_PROTECTED
