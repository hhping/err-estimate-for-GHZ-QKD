`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9+CAiKXNvGTFz6PxDEBfYimgwbEKzZwERV/KVWydb+YCpWGqVBDGKhoJac+5/RZ
31qCEgkfxevANCVOub7o3Wngos5VMsndTQp1KYy/Y1v37vEPYejQdVztZZaqs4nE
FgwiIX85Tgh/fsOUM4crTI8mae8dOru32CLyL+9Yd802+GdZ5/rviP25sIl/Yrnt
LEfuuv8ajuj10YoCNxA+V7fXRMY5+P53aOEUkv6Gf5C3aD3FccuP0kUgKDxNJ7Nv
W9MfGXD3eoA+2E4vVKuqtXj7MYgI8Pb1Pu4r7Yw4+bp5AFy4QXyJ1GM7yN/4Vl9v
JTugtsT2otqfE/5xLkPvCY0MJuxsPmjdFTiDJkjIb6b2ejWEhqmTgDfgbAfbOWwx
blVCjSBOU8pT2MFx7AJYcw==
`protect END_PROTECTED
