`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dfM2rISOOASNyJVqRqx/UmZRhCyt/GUTb6IdHNoAQNcmaHCT0jjo50/yZUrBjvXh
8uv8qD/3P46mcK9YMhD+UuzRowpqBCQsmDyESlvNW8/dgZCTp/63xxqaq7FJU7rn
dOKKhTHpC8PF5ta6lSoQD7Ydr2Z06RU54/rMYeWsM0HjN7Yc3Cza9Uqu9pp6WwaD
918dLU+oq85Ew2cxuXjK+7O1HgK6U4bzt+yKSQujuGfkypCDVi6aK2K44ShVrLS3
MSsTI2L/N06OUlZyN9z31zkaybrj0DSTL0wCihQIYut/DVLmWbQSlm3zT1xVVF2M
4cs/ZsxqzpJCFtK0ZuKVDWc3QHUnnWjau6NCLZfuDzbVJXDLjkbsPZhkpsxivew5
QJUpS/u7+sFknqp3++HksEPqHsPc2fyyZMtJ4erCW00F+dnqN6KWQE8lDxaMcCEy
nR1m0kaJP2TuTel0rq81WBQ1CpTkXzo3PQrfvRKuB+d9dyiXj5rjdO87nxYXfwYl
G8AvcNHtbOBgzKqdhCq24A7uKbbCcECwj92moPEvNpXrLiDbzbFQY7TITMPD5hNR
GLuvq+3UwlK3CcOLbgxVdYZTuRM2IRUQReL+mFzWhxBtj9uPm7Kb3KwnSTcsEF7m
sbkw2U5u3xQujjMTh4DSynvFyUrOaiVr6SOrRoR13hZLHsso+fFSiLsruDumhMB6
3tvxRZN6O77PY2Ed8YDLVFOnr9VHJeq7LJob572eet3FrfXlRlmLdfbneCq6xwWh
euL2Xofn4th2QfNJ1wld5SS3qGAftTtZYMMuk+z+lQWrhzHd5UFajsSf2LnJ3SLe
51e2lT8NOngFAJATehmX4sQCyUv5VHio5zXJqcNL+87rrykc05jvH8trbcfyl+fR
cF+o+184eBJT5MrbU5Vv7zEmPHeGp/c6hV5oYqmbLiOrK1bsAJS/JC+8d572xX54
FZPCH9FVyFZtGRaXLpLxTLsiC3bB/JV43eSRr8p+kNw8Niz4B0avLrXDuo0VpppT
jFjkSpVW0tnJk65HJEyOQLq5px+PpzWbFP/QtyVt3/IAawchyY/e+FGt2gWXuoyH
wqoBXJFd56VB2s4jexOiYTyWiBABtGbtyhR4p3w3yUucPXttE6YfSOUJ7UzDq2+b
LGYifk9af56OHOZsMCu0xxFXHKA9PD/q1cgrbmU1+AI/UQwWtiofvVTEjpsrmMug
4PWYaTOLArvH3aXguSKJ8JVbxU+w+A8ZejX8zXxnN8TKWBXXN4Nh6mk4I8QUXI1f
cq1RDHpWZdlgbZuTDaNHtyTMEdJE2pEVfEPKAbgDpmArg7opmNHRLB9zvMdzHCWY
gTcPScv51zv8oz5VLNjPohep9oUHE2OqbyoD6gSZNg2sAQOhC1EkR2H+bOgGAYaX
antxIoWv+m6c+9a7aIN62IDUPKZrUki3uxJw8Hz15+m1EQmm7JwES0Z0k6TNQPNN
HbixKIxss8csP0HffEam2xkOnnJa6PsR9lJrWEohn4gbOLIAWMjHI5PqIvFhE2CX
RLg4xA302TuSznJc2SvKAnUOy41YMJwGW87IrZ5TAYwGSY7iiEd7+FpEb2VUhMrB
76Fa5KAonuuPHlelNzeg8stxiblJ7m+xL+HsobrBdhOP47ID9+bs5XrxrVlmsidO
2C+gSiwOPfakRAnQ/XvfMJ+DlAs1VOJ4KfIwwh9Tdc/6JIRtcaPyI14g5LPJiMcq
QsqHfRHVnd/fcX8dXycBt/VZSyChcieviGx3NIUdwYo6VK13AEwPS0xQZQyBLN5b
Ou13KpSZW/vqkULVyAQGRualNhc8GVES9lKlT530Idv+JsSvS9zgnE90t57XgMam
wQ8x53OTw363m/3OMRXMrmupmKK447RvPLCiLcCH1aF4ZMqf14q2RsySzdWd9SFo
b9WuyJecJCTyeYVoCnpGPeBFlySG8tjnCve3nh6Uwr4eBVyGugxWvfeN42aSuXsS
AJqT8VGfQjDJlGx32OMPyx4OWJx0oXW+pBM10ATjogYj+Og0Ws4jjrubYIez7Gx9
r6EWmsD4VtWg9vwh6NScJX3cDJFNQFPCaN9/BZHZk0JNSItgksRLOeF/L8i4/QVs
Iq9Ew7Y5beh4Ejr6/NueouA00VGnR4GuxVzG6CufkYhvu/BxUEt5LzWDOEY0Efxk
AC/3E8WmXxeOUh+MPkD6XtXP0fanJ7TSb5XZhXtBTSF+xH4zH2zwytFLnD7FbyEs
0wD9fqLPqDw5t507NDUYwrha+YCXjkplily5fID7fAEfmSlI/dbWguoyYjwf4jHI
fuFC87qRS1AxxJZBznKrbXiouJ1+1RqevAANjqkr5B/9Hfq8o7g3DUExmV5IDDoS
S76sXiOPltQ64/WEHlo3X7hzMIY9XyRLZkqhsDmul1yrhpPwnaBNsdsb6EmTi3w5
Yg560bBM41yhdZ869icR9wNnZDsHo3SxyGF7q02yiALZ6mCBvFi7n3LyUgdF+HMT
kLFNw86hfMNmAGSUW/VbkRrZ9zDc62RuPCKedwPJ/LacKVopfM5WYTwq5k6CVDTg
DXbWqpdNv2oXUfXoJHPru6zCtDpTvuEnBv9sbZCvxruuwheOV4zs9yJ6Z++8m7S5
aH+0VMJeS+SZjXj/g/LCARBcHDKMNJBkY06WgVg1Ayd0ygTu+dRMDqw1qjLD4UGC
jb74MXqC2hkCvNch0brmlmY0eHklI0V9otD4C9vyN246r7g/lpNtt2Au3olh76Jv
NBnuKbd+nvk7iFpCFU1zIGBN086BsSEo3FVNlHGxpV1iNRiil7hAp8uVDKIlgxjp
oWsQNWsmTVnpqAwe4sGaAR+utJOA2p7TuwkxbHXgxtgddafBRudi9LdfJCNRNKUw
u+2USAKWTsjCSWIbeI0r8vb75CIy69J+4UyCTNinJCZnUP4q6s1uz1KVorwCVSsn
o7HFrxGoh83tGg4XLyF6/wp1ned1wtaYBzSwNxC6GEg4XC0w7jTD7f3QQcArF/+Q
jVw5kOocVld75vNLiVOv8GltnJep+cePmtX9zkBUiOWFqYfOANVvWVt2FIE6gAvS
IXtyJ0EuH6XjrRzIVN3EkIU33ykw57650zx/FY5kWkfZb0j8c2YAJvu3OrivzGmz
JkVZxm7vfKuhRo3QB0VgM7+sLScifPk6d1gRQLoymOSbXcrjLkGFPrYBIMkMcfDO
3x3JQqoys8RerSuzRSmm3e+Rw1tB8JB/B9ip3HJ98yz5jNQCx4dw+fMHgWKqifWT
ktijuDfaJQNUjw7CXuQasZ9R3M7inHniP+fQvq7UWyGNjCoJ+rZ1ROp6qF0RH9g/
X+WVq3uTaVc5tOOalwCHmMhN06v7EdgvABv5uTHo99xN/uVM8WX8AGVe87BJIjLi
jzzfXcCgCHMIKZUEiXYc2jZTUNQRRLzpIAOtVHmDNykJ1LuiBgU8VRre3af2CNPd
mO5cws/4Qq3nC+d2P4hu/7H9WaegPmUmJG/I2xlV78thfRbcYSkIIL0joASFIBPl
dRfILqwYtBkvbMydizhJeMUDlcI/GbLk8g1QO1TnAoJMw+1901fsHQD5w8T8eov/
DbgHaWcT87yFD2R5YioiWktjHRv7phTKGkeJzAsdoqotxgRtTHGV1w2c80Vpu3zH
n5TF89Y6D2l/HMquDRJk1E/BRBuoAZtI7MXpxCsvyxqiK4YcRv+Q3MLxhTxmJUiz
nQdqG+C1Ydhn2mYyjiKS7myVR6LgkNEdF+ZdrhJSeB3MpyD0J5m700VvhL/CX3L4
QUm6GiJbqqLahjlMYEXreK84qp2pqKHZ733+xBsQg8Z0lIpSwCPQ0co6BQG/QWRo
GMKRGzs59PD8/5JDs+Gc5+Xr3/R0UhV/oSkGYCFXGPeoofshYSaKbEuTGCAH/M95
64vABUY0cImWIY8h9HRduw0YzU3wIUNQ8IxxHefmV7ZKstJn4Q+svkL6OavX5LQ9
dJ8dvaiPG7vddvfuYXNMn5R66wsUHDb75gA3uxvinthvYZ6NnD+9bB568HiftNOu
/gdM7kbomOs0ejhFwVmQDz77/ePBY1j/hLNS/Mjbds6y8DOiltTCT/9oS/3BieAQ
xOnttf3jjeHe69FcOkCLGPcbtp5GKgPA5xEEj1MMPCr5S7S9K+SCe0bMG+iiOsjf
imEQcaMeONcPx/UUPTuKuWHh6tozPn2DaMo2FV5h+fL2x9/zTaN2zmFJ1OBCpUWT
e2FYpOg8SLSC1/iZFs8DTnYfKGN8RFwuSc1wohMl0tuQrUygzRXAX9Xhd5p5u3Wf
lDYzlVUQ4arK18AuSx51ZgZerttUeJQkeZWz+POj0OXRrfqFInoQulH/W4k4F1F0
8PQkl2J0oVag3WkwLH1X6Hm8/gSuSApxgSqIVIHCMawms6SuSrttL6aba7Q/gjCr
Cp9AHRNzWP8H583YfGC4XAMq6tf/ukN1DFDcWErHzyTptK4RqA4aeAnMtFMoTqDf
R+EYWf3KIdLI7GSnsRh9jCCHE2seo7pZuCChv6slcNTBZ5cVwHtTcbUqKFaucgkP
t2kAqeSGUNH/f1z/z473BcfUEZEdLqKuY2cZuLAOtvFanYZpHef7lVOD9TEL99Xk
jxvrjtEb6XGC/yXyB0v8I7EEGi7nDdHGE9LyUMryVCvKoL76TvRLHTUTljOQ9rxt
yfK8w0mBJ/hDZEgbVlhDklC+Okwc8QiUVNixAdMG1+FL79sDxPYkU5uKewJsnF4Q
gxfLxLWbcFKy9UDw+HCY0d8ZlXe5Iz6LSJaNyHJqdCHD6BA0O/oTvCrNukLWRkxj
K4FOmusmkBfO5Hjmku1f/iUHAh0GsaNxYE6IfVYTV6ETqCbYxb4Xnd79LwZ3ypCr
1BqXXgNX7ufmLB1pTp3f02B5NzaxH2X1KlWtBX2uV1ZidRCn53mZhHgPmL2T5CQx
qw9MPhivpAm9FvHVzDJUa5d8qhMYKUcGtUjt8OFPw4YH0fSETIRed/2AAVOunElF
rbYwh7NxWVsstspf+tolR0kUKZFHd+58HfOfn6uTIWicKzn+wj8eO7CsMIwIwubb
GAKcdR1OejFKww2gJQH3g4RyEtb2kC7aR07ba/mrUKabBFfDp/9n1OuWUYqs7n8Y
d5Jb/NzpSHzsxSc9eF8jePYMMkRM7RGVkfn1r882ana/uycMz5DwiGnZo7yOdT4d
XoEg+f+1sr3jsRAmAXox7IFEfhgYNLtg6ALy+pkehpofVahsM8CWJh+QUa3XDxom
YWgLwbytn/5/MdhrRyg3n1Iu6hDEys9U7u06C8fa+WV6U8vSUmP/sHLuO4nstUeA
G3gU0RjYOSw2wk49LHapz6DMTm/hdKOwGWch7M3ctwWYZ6WeNZh6/SG5TejJ6OrS
gUIMi5m52QnPwcbKmgPege/jM6HohVyjGpj47L9Dt5FtU7h4TKLCqwfYzpMXpmJR
2dslM3ecLf7zJf9rVJ6zm3V4RmRvBk81qINQrvpLgb7KvaRqwGf7Znjb79tl34zA
tBEnz2Yy/KGw7vY7tiOtz4jiEyia2BPIG1EBT446pU9wep9jY1rlQo79j7bVDfT1
ns7eH664cPpl/btZyjJ6lizHyUdRC+butEP8W6VOJkOFhvTj8ke4Qq5KAo0d3gyp
O3KF864re5gYWWQsv+6N+vdJQxavt+iKDcbCh3yQ61Ule89qKXl0vl2rvtxjDGhE
S7ddptaQoP231aiSvhShIrTdgB2pgjWJDTw7AGfVTzzHWtejT9cThD+r27AOyKBQ
ImDKP+kr4zXGqpPexXgw60xpQ2hrwqY+nKSTnXGwE2BCJ3+ePZgBouxuKA7AA+12
fB7RYuIVl6e4xUjvlATXEtFAtNdBtKHSIiutTWPAROszSwZQG7a17nAQ+KvahmV3
Fve5ErsF1LriZF+5gmFb5UJSlGyqg5F61p/Q9aRnwTZt87lKu5qHU/5pVlA4fJ41
u0bzwWtm6oMDujxk/Hs2/AnB9185xKqmjRYuiDgFffRHNIhfLiwJjXTe4WTF1c4l
mQdiGftHgkO7lrQgzOl6Z0bk+SZ4yvb00rsjSIDdCtIsbaQgOhT/n72DMnoJBU8/
Xoo4W34HUH85BodyU3ampZMoirM4aGZrjcZkamvX1TkFin2dyBy+kR+bYKj1GWN9
HtrG3Rx/t2qL4KGRpcFf/kOfhZcqEp5a3+5pdBcJLWTqlbDQORDzhPM9t3TFEl9G
hpid9aB/ibiuyzncNuMvdiID5SLZlvbAjiaKYnccKPeKWbLAPjEmPUDrvp0/7vHx
VCW/oxW9DxcvYU+s/RntGxToDG4Qvcn2v44AW0iBRmHlcfROaNUaOhTLJtr65L/e
h5JXI6aBxye3ULIJZ+ZF/l1RCSt/FDXLFnbOdFuYcnRP7bV/HtGtxWxhMYz+VUd0
tif1ldRA2NgIstBPi/feN6ULgvUk1JXMLajN/d8RpCY6Bg6IKK4DDow/vD+5V/1a
jVrnv0EzxLo/kaKMeYP2Y0I89owEwRzfguwWX9uOQVCtsPaSqaR4wY15DjsczUfp
hU5SonPmskvGcLPpe7ibsJ7BRLeNm8KGCYfqL/svUkkVdjbxu0U3SbhLxFbPCQvu
tAOprcTnd7ehFGKVvuAHNIDRUfZqOPJdcXXJLERunfJFQpNYOk9c5+9bOsyf3Cgf
M7c2f3s3jopbljZdQPH8ZIf1ggYObGk9dT53ASn2flG9+aaOUfc1RiEBg1xJC5Lm
qSgae8OUOMH0MOZ3j9qtI6jQtYVPJuMHnJIksMsgZ1m+nALp/x+d/5KPuWaBC5n0
A8mTArg1XIXZGoK1zwJd5liEkA4BmhO8+95/XjNXFK8B395TQDsVhvXLUUXLMUt0
Hq84ezEYQ9l3jCkniizQMMKd2ScZIiK2NKlgg2QCdZUQWR/R1DAbm2/tBO7HePxX
lLfqMnzUwMIKiONLLIZE2UnDvHa1cEaGOBUCm5Ns5ZuuJRccoXW/j8ZSpNrOZAPE
tNdeXWdXuCPqSdgHOrLl9p3Y1N7Emw1lRJg25fwoaPJWTC+x74rLUI/c3kid+gr+
JR8opZ7m+cSoR7uPf68ed0cExbdZg2Hzd4TM5VPv+U6+6OFcszHem1AR084LT+2z
gJZcEiiqS2UZNU/ixGZ0itwyPqsAxjgrPppSwPdaiSjhm/KQ0HjawaSQOKckGZsF
xj5L2PLTsc+lFexG4+Cx3ImuOcV4a+/IpGKxwIpwK2/DqtGH3aulQPlSz+hEh84Y
x184ZlNVeeXe7l8AVRuXw39zI3ksbu7V2OIOL8ntumBf59qgD5f2N7YYubdhPtk9
jI/Mvz0Bo0A4roSyOdFu3yLrLLEOq4YzAWtqahu11zfgjfp+8FG0dCMO6Fo2818W
RGknmCe+e2r248IrEdxT2f2mW+TLBrIc6v4kLZwfIYMcmny3uY3sVDS5HsnDGopx
Dh+5e4AktAbIO2Q2+BF10JLWUkZ0tmY+IVN7Dyvs+0otCeGBfg7Q2IqAmsN7xnOO
dt1UXyjSGt6lJXTc9qUtE9jZjK2J3uIahgHT07J9rF9ODJgiTS6cG3O2LeSydLyU
VkKLHCGEv15tVojSE+r3pZjHnODhbNxwiSYi1Uq9P2Ij45I5ke9MbH2d+dxDQKO0
Soe4aYqW7Z0mk5ALe6OqnHb4HilNTBeQst6/9TjwKRdkzEAB54ddOX1/a8Z/neYT
UmeNErDbtn1CE3ddmXdI14EIufw1jyGPaWxs3FdueaTunQG97svLJv0dPkemibn3
WHKXGtEOeifjJvNaZ9JcwQUgotYrWhc7EWFfFAgpDt7p820vGtfmJGXQxvrURvCz
Y1ZH65oE+xHfT29yBFtSoFregOuo1JhwTPgQTqZTAT5lfiR2Fce5DxL/F54CAYL8
Y2kxM7/vxDrMz/IPBQ8N2DbPKI/avP5nIcLWLUTJmHY/8gL2OP6jko01sFvgoPWO
onwWp5CttdCXF7R4nv0wm04NezWanKZ+G2aAOq16KsDBMl7Iy12CzEMpHI8GnFJz
g2LaZ/6pdxt5dtkqxVtmgcauOn9MvviHiPjfaDUJYJX0fdKe6Vm56yR5xAcBidEE
lqs1X3zO+TcQG2cGO+nGtlc1EAQA22wgcwRii9gyGuQM/o/7yBg++3BfsgLiL9ma
wk45LeQgvki8Nr4BXzeYCqDiBjZP3bSGLf+mfMtLBLRpMDin8y0sAfULJZKG9oSH
qF6T1Q8KyT4HXNf/zlbnxBNYL7S2PHJWTykS5jdFqY4btbAFVcqToslTNvOs7oNI
3jaFXob/idC/8u6uBoTNsMbSQqQco58Q5Q0E0bb8M0pk2hrnCTCzeba/8dINjM9Z
gijJcMtTP4FD3B998FdFYh/C+ohejhR+ndX4CpBWoYT3k7K34u1i+WYNHtyTWQGz
+FpDxP72fZDwxP7vCSQg49Ka5pPVF5qBLc3WyOKOXxxGOjXRql1Z6DdJnE8qCECJ
LOQd8vn5hYlPsWlO2qj3lV9BC92h7CNMJaHYacguCRIH3P1ccHdPv1oAjSc+twtd
2IzjDr2R+CaLJ7sCLlyRE+VI+6lBU+57Z0WaBq5Aib0Nzivv7SCoRNo0qZk/q8s0
/Nw7s6Hpx6jq5f/rpj3gI2N2dcRiYowVljDSFZjnmzbalSNDeBqhYW9590B+jbVf
6SdeF6qZ1E+BPki2x4dP3q9WXFFGYtgkGFxgaS9zPgpQJQN+MvR+LjjBzmJuY4GP
EyqCRx7L1LqrO2UQaOLqzCqyhUGaDDmXY9WPP2wMHaKw2TLZb1qYPhK+ikyA1cWD
x75hgewQJtJGTWf4JTt4zwv4ksF/v1BMC76tQ6ht7Akkk4scLZJ+gNQQKjlGS4oN
sZHJM6Eaw1PdGtLWBgEpKBtthQt4nAvCUVBYNALXthpClIreSJE6uNs8Uyd9Wo1d
OLBFGoxosnR2UUdWG/F9KcByn6/b3MvrhOJWfS2G1nvtXVEQQFG7bz4F3zlRqF5u
2MoG/5ZS+SG++Jq6sGsfxLsyAIyK8bcw/EMyyJ1iP1U3Ibr4aeVNOZFKODhwQ+Pk
TZfgUz0yzQcGnqTFXoF5y5d0YgwJH1MuV2e4cu7kYi+Hz1kWroBFcapdXRYN3qlu
vvNwPoUUjxnzDs1LgS/6aaOFHUTA8RvxGOQ4RPE1KrTajHaKDP/99QBrXYQ1UL60
CDo4BYIN/NSJcZiW9o2ObRl8VNL2jD42/eClaUGEyxJkCBMIRFoRvzjDAyDF+Ks5
sJllb44losoUzVSdsYO8LXUifAftJsT7KhDDgsPSoUgawZgxBASyUgnJKe5MrH8s
cT4R74r+7svmod78zElOtzNaUrRwLHCDgATxan3jfx4R8YD5fbl+2yld4v+Xaxwi
1G2GnxeNhSX3RxN+jhgcCC00eSwxqw3Rp4jPmOGcBBs83h1B+dDqW6IM58DboMc0
degHaNAy2awLtG9beFWyKSUx6F1nbcFX/u9QOecOTyeSmKiInD7YUVg3d/Pj90MS
4+k6rjACjy2bt3jTLeXE3LxE0SMOui4uSULXvHofMlgib8OPVbTwzlw0w/T5U6ZK
7JfXSBHjNviezAEii4pYDC88L2UBpKqjULLPNs0UmWzsiCXuSnIbqOlqPwqsPGQr
C/Qvcp8b/u9TRAwdC6DFFwUdR6bAdiEZO+h000Oik8S8kWXvQerkBdyRyDq8I8VE
gPJ+uHZ0vpqu8kpP4uJTkYIeVArmQqt5rY8R19VX49A4fWOsrEicuZReXVqS1eZs
GggTnOtk5E5Iqk0do1mFQicFZWBBbmnfxK6PvbFvoloNfrCo2oBYk53JlOGBx0Lj
azupPzwmg/7uQ3lazvvS43P6bLhnQdr8BMDRTqJSDcKYj18HnOAmCdnnT9R4HgG5
Cvqt0UH85QhyVTc2tIijhIrH56XffQztHd8rdtYdcK/wsmQWdTvO0J9BO5oV0plp
u9Sjkk9oK853xPmeWwA7XdXxZtUR9xuOrAH17XO5k6Yh9uJouENbuC+fR6eS6b2+
MIvFlpvTQRr/uBxwxi9GZB9zqgnRYWCzDd3ji4I0MP0jcMbiffTliS01zJeXhPn+
V5jDWF6Xw1+HBRIoOw4Lcvq+VO3kEu3L2+COWIjCEc1DAt3++2A3mgoEdwADzuwz
cu3mfUouuThzW9oyY9qT2A2/B1xGBjJoCpIeO4evaxL0KGsEs3CUNtFxVoPjXVy5
44vpkvD8ars9JIa82YA5AbF1nWKb/VOLd6aD4v5YkfFSuyWKE+FHKvjcOgdm7H7F
rPNx75P/0M8oM/hHXY+JcLJHDjKsInLB5g214dZiRuUvzblK8y0SsPVeW3XyxGiJ
tITSeKcTDmYM5cEFt/17Xa1FgX8FcUHdJ0S8zRGUlhpLZe2LDHT0Xdc8SD98RViC
kHId7vKlbwS15+OOfZp1FFJP44frzdP08+t8B6mxfQHzABmXLMp87f14JOWjk/3d
zbW/kKddmq6xkFCy75S6N7MJgB7lAX+nkT8mD6HNdnkMFsyRTuHvRhV4CCR6GE67
RB0u+liWSoQFNWUWa+wyU70La1yii9YTOKFuV5wGaaYXDgJBihg2bUslud1L/RlS
Vxnl+azACPT8VN5DeEuo49IqdeCeAbs70VZ8yMa2oukuZ3cGqjiHmCEfqadT2ZTD
KU+9kxTUoERfcRVGCH6lrwb6a2H3bMwj0lFbUG8k1KTeV1+Qu3o3/F6Wh/fc7/td
19QIOThAJIdjx+zpNvz9udgvC/Pn5KuTqQ3F7qzFMYCQIKnDV/w7bH4H+cxDX1JS
uIyoLtSzFEPc/O13hhz0MSVWjFQYTdnZKOgPvdVC9MYnkSkABczUj7s6Ic04VsbZ
jpOv+lUr/kDDx0Bm0aK0QCAKbjiXrbqIsh2/R5QVfymmLnSUe12HjqyXao0idVKT
GCFvTdfugrWJkUSUnhm13zWA77JVdgxkrVzgNsonAqoOzxdmnAHnalyBPWetoqna
Zx4WuslS+62FKTHx+ZILOLqSM2Mb8FZ+FbD+/FUYvz8zumC+x3O8U3rAgNb4ryaf
QaZF28oRCQlX2fgKs2KV0cgHJm+T8eE94X84yxyOUFq9XsvHx0Juz3M1bEr855bS
1SqAhVZ8ek/VJgKO4Wj53PZnNTxWBRxs2wbNjGMv78oz9/LAEaSmW4gSOfDOF5ew
FRaE+3CXoVisoe/PEdpAbXJjL+Z3FhbKOI9jFfUq/SzPE0qjdVNnIoy95M7PDSDT
Atl5kIR5p+yt67Sp8Fod/bqWK4NSTFkCs/VjC29TDjC4DutiN5zAWV929GUYANNd
LQGfhRAcPmAOSRGuMolTEBer9dTheASIxmtoXNgQXgjkfxmrgy1NNJm5e868DsJf
w9zLHpLpAAQf0gNSxDJ5pVy5hx4qPNM/X0xnvc8I980eNYufnzUfkoGyb+Itzoz1
GQ98esmYGdM4FwBtzFGr4Sj9vljzvRNSiZVbo8LLOJ156CFTsu5CsnQqj7Eucyww
NXIdpB5jVBvJ6T2rnIqmmRdSy75HeDZMVq99o3qM30I8WNuOxQ+C9ktlS98Ok0m7
1ToaDWSI5vLoNg4BLdcOO3F0cuYFxsEWCUJoA0OW3ou28HvsFcxsIvCXofGsooIG
QV1H4/a3ZQUClesfN0hvBz1MRYk/uH8JXZtgficBAre0v5QNLYMGMrd8g8uAR6AC
ZREHYMXfyC/QuWZJApODUZPISQ/L94gIQx1wyXiXJC/SnBe1qxgUMOCCA7OZtUuG
5nFLDpmPSPiwhF7qYeH4qyHyltsURE8xRVmkpj15asPnsALBKAiiCU0U3mO8NRRR
SvcRcrw67JeHaswjYdEC0Sj246H5NeZ8qnDFId7lDu6h7g9aZXz+gso78dnuulCj
0FG9S3Xp2q/pfMuFGACbD/bbb3qZ196b7DLCmbRppvEK8BL4Hd6YC5tuj+k+Fgsn
HORXYxVQxG4uAGX5Ktw1B0+osSyzZGHrSBCUQywHonib2YOc4yuHmpVhxYNxAskZ
3f/Ce43oTbHmh669+5d/efj2jhmqiNzXHmEHeY7wIiRhGIIx6xOOHQ1qISYEib2K
XjfjFBsp+VI+T+qpVH8BibbFfF03OvosEkRcRHzBtoWki7gCFheHQEOe/gJ72mVT
59LwcbpNYjHAoDYnoKfXpotiDUb6/WRiHw8qkx/6i+I=
`protect END_PROTECTED
