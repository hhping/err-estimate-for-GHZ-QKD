`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9K/Boe58umOrs/m6uZFGNnegS8lgvsKYdxp92M0WQTXh1xae+ZEXZl0ku6+M8My
OoKJQxHRhEr47D6bRvNTUH7jMc1KilgFd8jnZOfVRvmQ+LlkIXIlyjTyyy5ahW49
FH17y8GgI2nEu7LzoDo6axpbcmvZvnTvOjl4P8ix0tdKOY/2GAGiWpT/3Y63T1lI
U8EiB+eNk1MeTPw59Va2JTGqeN2Vrfxm3pCPwrSCDOTFKzjZdE05SlsAHoIiO8Z2
/GjClXdTqp8gEUz4AyHDNHoAjOlQ7ywRSroSoSWJka4kSL3EGfMBLTOJAjgJ5Ie3
DmW9ltFYjk2049LWZar0j1hJac3BlZRyduxqiM5kDZ9scvHcpdLOssEjc0CYEXbl
Z1TLy8g76KhSNUpGAVKByPq/U4+OtB/stViaz2q+2p3zRQ375rH9BXqr4sTj+eii
Gj5jkr7SIHSYpwzCAGwRVp3GNTxqY18BDyGpp80hS/J9HpFEBNZwFqaMu312TXBY
cHlB9WqBN0lgw3c+v51Eg32+6ZyR27LKiObUQMX0MPhNVgLPumrT3B3pm/v9V5Z3
ic94jSlcdtbbWl/L7HeALagr/x3YAqkrK1mKhenW6kv/VP+OKOb/9G+S6iiy8OBb
rp6yM0Ejk4hQOex4OGcRS48CNYio2eGKjBC5L0HpcV3chxWyzBDdjRV32E7rCJ70
AruKElj7hHZw9yNyqJYKLaR0W+BK/R4nXiBoY/VaLjXj45MY2Yqa0Qc8UVnWwh9r
egMqoititpU3bDgzO8ymoiiqRtOlIQlTqGOwiNiBzV3mJiX5tuCTwhonaz1zMBEY
kAWcPj6XI0J+fjE0StCcDzTn0g4dLJ4PY/0hcs0amv50WXL8uw5iIglMUi+ftw3u
hf3akVNHMv0qIFwROTaa9R8WFY1fQ5Qhytz8KNZmK8mbgq1/HQ085qghgXYkJKkQ
Hfjlq5ILOnlsWgKefRxM4jnfSGLB1cAYMAEEMajNc9X/ZXOsj0bZLc+hPwYcSvgX
Tv+GjlVqiH8SuZ6QeboyoT3qGvShdujBILTt1LYYg+jEPoEO2+t63Cbw/pNdx2RF
9MlkyKq1EhhtYSleRR3wYrPzYSh2vJ+tvCLhIeto2irIdkD2ZqQ9+oz9yN5jhXp0
sJDp6NUJM1uGZUyH7HOYN0YsDejZJbRH3ud6etdhGpBvVsZxqolTIh+7tgqHlF2R
DtB+JLtuWLWl6vbF6KAXud1AiD3xq5xl7obJJKNl7rOsatpAAMr8b5JsEATctVng
4yEUToUk/Cv/tVUAp2HZ9tEfnihhSwtGneXZkLDUQmPz0ZksCsPWJ82QITM7kMI1
4y3IDEIEgDTf8lmHyKSzqseuuR9aRKqu3UVmV8hhahPeEU5X3VXetjStKkAcSoyw
75g88ua9lzFKbftmkXWhPO6ZDhsHfjtT6W11tE6p0uXIJwh+3Y82LKek5eucs7+X
n9pcgOCbx+XFyz88/miceLjoHzaUua+JqIb6Y49DaMJef4gNoXD1YHmscUzntuHd
9M3BVJTyQd2RIpjNg6eHvxDLEbwrqtCVIppA6nx9k48XcjD669vMBCKEZZdZ8+wF
s9VZwHBVVglpXBmavM282Zy1O4+GMlXbk9fVD/khFuJcEedq/DR+4K4NOpfo3lcF
mXKnErwBezjOOSskvSEpL/5DyTUyfmHxQmn8qlVJhOUk/pPvAkdg9w6pi6WiDaDz
3HuCKrrUKueK/8ns73CciVYdOK91oX9+YEcF8s+fD5XfjplBg7C7LRW/l0GNZ/T7
KwY3djs2Z3aYs8UtvKX2B5L7K4X1k753zQc6TmsQc0YWyEhKk+F+eJq6mvzQtFo7
8cImIHAvoeIvYuUnzfWX0iKWf2QYK2qtelEiWQ/exTY6ivhZqXveW03goMgDzSyy
01B710NNEV9+JKUGwlbD+40iFrHJcGzPDSxHbrCXA3mxYCdHJ2QNj07AmBWfiaF5
LSWc8mg2CK2M86hOsD9BkVXM2Ibevd1X60TONFQ6Zqz+jRBpa1IHr5syX58Nt2GS
hjIizn9Fb7Rw22seGbOrS2uYmUxQjWhtRsGwQ7DRI2BfBa9f0eH95/LG8roQ1/iu
Jvrf6I0EoSKDvGCWLb3SfIbVx2akbdYSfLlH7AMxE2rbUBwVXsdK19gQtlh7gXne
wWE90OUSLv7lEahMNyNUKkQvPrIl2Evp2r3ewAngL8TawV00eX3G1LlXJ24nuATr
5NG5QJ95cqdn0301saG0kIhcrZ0a2Wh83RETmFNVeeuk2kQrcUdl/tzyBP/eQwOH
l6UO4ww6euh8EqwvUGL5Zeu4DjzcuZt8zSWUaIgQj3byBbqtxWR+vqY8ynyNRqEZ
0gd6xTSavO3BdvWCrhXoVKPP7ewTdImmRPHvOkcXoofo69ZZmdRG7LHjz8GGOziC
u+kA0i1uOaTvSyslEH00SvSYeIgYqLD/7pDdYA3DDCmXLt2hJkp1qx3bvtBg0m/y
BPrrrH1qlmhPaekbKeGgZOymsqmgIsDnXlMF+ElhWMlbSR8WI/yuoVG2xFluDdc2
WcBYaaRj2lnjd5TeCuqRcZUIrOvGaaY4xdAn4tTGtfRr+fnBJ6DiIAOwNImx4wG8
FKmVb82KDu2Zw+VqLBV3EGt6WS+74B/16qY4dZGyzx6HkU1lcClIwpOdnRJkEIo/
V4PQFg+12XGSASmGllZnX+57MPfILO1jf99DRk9+vGsxiCKKT8WzeaS0S/x/YKvq
Em+eTz9M+9Me29lTjuCCsZhgJ9qAsbCeWDXAfivpWG2bMEFqoIw/2NZjNOp+Z5SU
c267EEZhScN8dh3XWAZ9ZMradi89tfZ0Ct+1Xusim966UoDdGQyBscCDENOhAtIa
KjC9hlnPBN7ZfKLAos3j0qMOuBvHjf1JnRjCj9/MsLvqb326qNwcfuYCnOROF11W
RySRuG0utM5MQROAmFirQg==
`protect END_PROTECTED
