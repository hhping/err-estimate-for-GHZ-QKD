`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+NRh59m1ROWgwRPKGsrUh+tJUNUeX4vxCFs57GaqIJ+qhNMVeD2v7NuWIBe94S1
wUFlODXH+hzgeEgxnCy2jHbKa98y71j0SgiYWR2Ryb1PFj5prJT5yc3Wjhp/Z6q2
iMmBSyjNnPZRrTtb6A01U3a5wgZjhAwETLdBinG6XSayUu+ixRyObbQ6Kat8YcqZ
yfvHei0nyQ15uAblRPNc6EkCY/L8pkJf1xiNKEvZ3GphYP0pYHrJV5LU2G1/yNzf
6UWK5RLnabS9QXh27vxEmZGpcX3L8/lal35bMzzfXogpYgID+5To4R5p3404b+Ti
2er14wLCbekzyKTFcH6Qde8nyYkmO2OrhwLjsi6nnIngxIeaKyGLFeJe8Z0HmZOt
4zXEjAw4M+H/NFdMokMJpggtlDHwO8Tcq8sMKQPEIhAcEk7/qGesEiZTjxrMd6KM
Pw+UuJxTB57hC4+so0pmqbtcze3ADvD0eUGHgl7o9w6v/8vBXLZNaoqMpX/3u1tR
wegOKEAPei5ZX9T6soSZ/WpKf9OTzOMo9Hrn+PyDoHY=
`protect END_PROTECTED
