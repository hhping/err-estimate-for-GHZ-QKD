`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WkAFh0TH2z0fj70USdvHL8eRP15NCN9SNjxFujwjuZ2CG36euH1hiivzAzt9Px0/
R2ObEHB3gD7RgITk0drJ6Pz8ze++4i86OxfHLCtBg/dZDo7rdrHyHQg8rbnRenMQ
eX+wsiha5yuEhRCdzuMf7/lrCJIDNpTDkw+8JB28ducEb6GWkZ3MESiCqVgRKlxY
PoTa8xGI82qXX5g1Us9QAmGm7yIDH0eA7WJxhITBganSdYzdYkB9jHzV/Jn/Ez9o
rh+ARjn72CMJLGqY1eyBJIH6gLcVCRyued8tjUto6fz1y0PPtw9WE2Dh1bQZfAL6
cWkbtaHWm/mC3z9P3+je3ZMJIdkQ8sExhg83dThBdVeLyI8WivIYPbt5fRE37IyW
HhiVjryT9Lg1eQf/iHmQBXkW7hmxKWITIJBcBSi5l4YuiCtgaVFnHoXOXkWFHnaj
cp8QKTrlTUT4/Z9woNVMBlNTHdwMB3udoSzBIMRnafYpWeEgILYxRr50FhE2ip3x
fe6TuBbRg8lQAuUBYvhQsKnZ0lCUX/6L7JDLZPAddGI=
`protect END_PROTECTED
