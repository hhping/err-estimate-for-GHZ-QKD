`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWftGdlHBykO1WnbSPFMGv0na/g/ZVI6f/5DcsA/XwihGzqBB5StAQdJc9xLztlg
yqDnXEUn7pUn6QdAsEnPH+qZdzfCALfnb5LGXZzC83ZUJySkIha6n9r13xympu3t
a5vvsX2Jan2AlNiWnipf0BAlr9I/UzvQonyvcfMhOILRp/Dl56/ukni3OydxUnl1
j0FnfKp1OY+D2gOgohQ+mkPR1SJciD/F1+PnabvSTU4HdAGhKuMiYr87RQUa6ExQ
79HqabAJNR+LY2loXjnOc5G+WTjpLPigi8F9ZWnZEOHbxllWuJmRfays3OToJ4ys
Oz8QT1l+NFiiiQY47vLecqkRO8GamBRr9j8O7vMc/YKgA33Rn0x8F774gBcI6vr5
CYe5pjQCuGtC8l2+cwBxgpyMxxjQZkRKaNQGM8tqmb9rw23MvxmZCyensjZwO6+E
mBBNhE1qgHzaWXlA4z95aIgoAvBUgGztXlTzeGnjW+1g8oas7BQjDUL2iFofvSJE
f8pQ1nvSYxwreIBEOtt9h/+nfTL8cRUMdQQldaOWSTWN/dqptgwffJZH72M+UZSF
ssnAhm5L0h0Ckf6EulaP/+vGPM2K9yNKXGZMlIbnMaSAbmjn+MopfOdNQ9z6BIKH
SUIM7J02j4CHIbhpoLD+/YazEIhMKUdikvrIjxoOQrxU8lOdfIr2GQRKIT1K8kly
BzeHHhSY7MQ3BET+M8JDAns3QrnLVxqEuRTyARicantE+q7VMcwbak6vS5FwBLDV
`protect END_PROTECTED
