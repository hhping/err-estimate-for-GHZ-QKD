`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p3HwokpXaVvmtYczITuVP/1pNpv2JUdBb9IVcL8D7m4DEHvbRBAQ3o3c1lGlrJnu
xUT4hjQoNGgHw0c/Dpoqoy4xAC3ub+uMerjUYQFI5P8kuHQ00mvtK2ou1k1UdUTl
ay+ebGnlNJWSXLDUAHx17ShTGriO7oXAx7+69fpbr2P43yp5ujbzuM2W/R29Yngc
7VU4vQx88BF1bCM0xDiBaAU+2BJ5MqRSuV1njKICHd2s4RK5U3I6EIvGRAt00iIF
il6YoeV9bUK1xPWf2ganY7ZNMnnfzPPI7uTMLoRZrMRtQoOHuARgojPYWhfADyz6
PvDCfu6e1qhCJKUIVA3RT1cOJzAyXbpmK667SVHi1MgP12ymPcKQWZ02CrQTG/1b
l9JO5khD2DoMHSL4eqOhOO8EeN/MYEoHF1DiCxv0pxLrNNOBguf6+hsiP/VqUPKB
W2nDWkRituq9w6oValdV9nX/sys+3JqoOJnuuP5dwbpdXJC45Zlqdsq+ieNIpr+4
NesDKWP/LZJ8OWZwvvSh0neaGcjD9iRMR1kJ3OTf4kE++jBqJJv3P8Q/U9VzwbPy
LQvjVT/rudRGv9g4CcRQsdUMPvVzBI/X6kIkULdGPVBIb481cbEaOfEfmz4YuWZb
iwH/weRSaUddLxGoEOfxOs/t4yFSnKB//q/gw5KhRiwJDU1nO0I3I6gotNG7Z4eC
lQC4Gr4gwXZHavCVm56bE65jD24Bt3XG0AW28RbpwvyUNgqgdeI8VXD2oD+aBT2j
S4lGx4I/BaL5SI9L6JYLwJrGpn2Rmu9f1nQZfOFHiynJ5GgIeiBsMZAMpcsuitod
g/GxxESXYSch9XQWdhYKGB2jVA550VJlbPtnohPRs2xd8OKKaMndkK3BmagSz6sM
DXEKHDgK+9YwlR2r13dTVF3IAamMvRusCpTq/iIeyEDoh7AjmYUuFQyw2cdM290i
7DbsTdUyXsSib4+qREEBhsT711n8ZxYu5DSALOnfZpXzLRSxd097q+h/2ZUdh+8Q
R1UdTDVlOVPbCs30Ap8A6FvSz8rLzYv1yAAlXaKxVWw+FwQJrA6PKRz9jl+hZ6y2
0YsAbgn0vqsNv1ksSbLG4kmAs+i69cIKNRCrWkd6OEbX2rbMWHtpCk8/qvfu5Wxf
8HruZ40qmPPLFXZY6eJ2n0cD70so5lwaVdK10hxqILQ9LTijpATplMp2SlXi6AjK
14yuMkLc0F27HhDxeHr4uYMfnjvbcUmr79YEHoymb6122SykOnhD/orsQtO6yqN4
O90PKfKlrNvrTOYy7q/3as+F8ZYmkM5iuE4TSsR85UwuPXuHz3MIu1XcyX3fsfBq
c6nv7iTZmLyb+Xeuij84/g6TqQGO83+jskuHkIRT0CkJ+R4uLunkWIYkCv/Tz5Zf
CXY9KOqKEa+hE73ntJT8zhhsJFaeh9dxckd+g4XyiTWNUGtbnLJCT6zLWMJrpJ6Y
SuNWG5KTnpSWycuX5t3O9xU6J7GAT+U/KPopzspOe7pbaaiFfVnrsHzPyaeKI2U4
OOpLp8ul6G/TqU4rUzDxF0D+NS7OsFIoLTXpUaa+iXvBbFLCOktbKZYOTKEJ2iSM
t9emYTAP3GjxnluWqGkZGOs0bWUUy+Jh03xYloBT9L8YtDjuYUSjTRyEIqZTAfRy
n8vfQcnC/D0STptjmGKkrtTnVVd/yOdg0sX1ZiaqaU7aFm+96smjkbESRYbVmQ3p
6usAqS8BBUOUi5/Yj3VWDfDm0VpeAcal8ylSt9F+h0k=
`protect END_PROTECTED
