`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8/gmTBnt7etVjDRu9A+iOGAXKZTlw4VC7opLDnEy8TAtdAwSwNzALGyy02sC9nr
qm87Dkb8XENG9ltPTEyXkLMUz9XRPmbKk3y74K5d8EyBZySYAw5iGPvRkekegcDs
PJr8ohQgv+RMPb975CW8250fzWqUPpp4wjeIgndYVWTDMHQAIRRgIukczYN8kuc/
s5dZWDxNz6YTLdRAccSm+VcupTuI0zUjVfXpjw+VXAlNQ/e77Q8rkzgDUN5/U2qm
5uhixG5wacLgeTmwpfSdMpf2JCKuDk/XE+9Vyf6wa/B+Bs7UHs/uyT6Xiek2WMQ4
4syc95sPDCQbs/hyhIWwTJQtwpnorLgd+1pdsGl1yQVazQQLPXl1FZv4ZdI6tAXP
1a5QuC7pitHNSCNxtRaq6p2h13SUtkqW9/J/NDfFIiFiC0vGds2g6WRvWpNg8gXt
dqx32edbqX9dx280edqNugJ4rQvuXFX0GU2Whg2Ss0ihkjyx1hxDL/tf4lWwTe2p
G15T/eh7ggnRJ0a+2MvE+JcRZR5sJDWN5PQfTxpUd5L8+uJrF94+AnM+cV4XusjB
b3LDylHoSAjJhpxlQidM4xTw6ZIjIGwKUfZmi76zCcvCNh7pTgd4gb03/RMMSaR6
Bfb7CAdeEHKR52o6VIYN/WuSlqhWxzvnIrK0CMaxbE89CztRhfvQvTpmeVoKjnli
dveoIreUox05Dz6IJMArz/o/pUL5bOvPew9vqgRZ66srh5PK1YgULGa2C5l8fjpr
3SKAEkVS1YMo1hanB+FMAzrx58O7uICLrvfGZbDQ5EXqxOUc5+otZcPhMboJciwD
vnPGSmyuI04eTIFekyaShiriaBycz1uoHAx1rjNaYTN5vjmh+uN8f9eTJBZhX43r
/2a8X0aWM6z1K3IFxfApoKuDoR8/jEUih2FOe8bFlT9hUxhbheHEgV3faBF9X1B4
6vFybG1G7SYLjV11Ubjvs23oZCM03zk7qPwL9H9w6QePaJo6nzIoJOKiKJx/PuE9
BndnOEbjuIqRNB976oEAQ0cushzj2nULST6nWj2jPEUT6jf1jql39DEgVt4EIXcH
IucwEW12jC8oP9wKopJZqmZaRb26mBFwSdQHcwlVBASbaNHLutVgWVv8nE11R8VP
lNchf3v1HMWU8EtGuhCqZsWGtI7e8+IVaWKZ65pnZZvr5BWiGQR1dBT/Y+NY+kQj
FsajRCv4KgIVtGx8kszVsoP0DDS0xaYIJ8i8aZU/qc6CC0uWFq4na+nI9erZevQX
Gu8TVRJFcBqo7vKW3xo9N4yr4EtZWgJYHOucqYytSSqPIYMZdKrPUN0qeTDPVPhl
gIJF/pWEBfU/KCIhcMgQgTccLThDgaAqIn+vXbHIMSnUSAWK8xOYzRgJAYLl/I4B
FYVgukk4IXK6gJ3SDH2KEyJcPfxdMEvpSqFKczTH4HfBjdZlheq+HQbYx45gnPA7
HZak3kGljmLmsuXNAA2ZXDqwcgiW+HZsX/kE+rU0/E3ugYAEvlkhaOnUF1vqMPwr
xSt/QVZzUQ1lEfpv1/hoMWArCeDItOQuqMeS5A5ENNfMe4pMYM5ywjPOhE0i3pJJ
WKE1k8XtYY5RYnzYknKt0G8bEZaHDrnv98VRCRbWhfOzsxu4aLedTvRUgrIjTKvj
C1nblwRTxBVp3q8cOFLnYxr9TrLdouvtrRz2GBmz33HGm13AtSLQjoI5leeTiMKU
BEjyGfGmaVIeFScV3rnbXcIwk0xaAmz+rkMbW1NAti6lcrzIDHezv4Iag8G4xmi0
bWhnkX0KaU3YfobC3kKRb0yzcbfYKmOHBcr+oa5p3ToTPFbKs5NwRuUxN1suTqMm
6sUNcv/VN1EEjH/pRVrAgp3+ea+8hj/nuhufWZItLzr4YlEWH5N4yQZyRr1P75zT
NjGdKbBbk9TOAG04KKu/Ac2lgDYLaib3uwqnTyVaFXOrOMDGl8iBx6OhP518h2va
I/d/WIiLamx/54drqgOrxquNOLIewtGrCnnG/6YwXVg15pY6q9W8FWbVJ+RJtTi8
pDSCTBetbAcWR4ia4gVWN92dkHa3XEgCsjTudJughOp1QVYVQSvpP5Q9SWt0PPVx
4V8yDGDmRceKyowwDuRakMzLb4ziDeStiNMyaQmjTUqabIbWkMZjd043piPZXt9c
VX/M8ric6kZAlYvp9mrHm9yx1Ed3eGmGPpUB10KVmseDYf3D3ufdXvY1B2VfDqSO
WSaOEdc2XZXiGje7VozrZxEHos0D+s9fUgDnLpYoGcSAiDji8QzZznATtfWUhp6E
Bp7Bc670gJZy49Zzf9bnMpNTMEV7eOGK9CSOUQUVYTKRPfb/y5TgR4LNRIlcOtCO
5uWdZmEy3VQFjlQq8rkMIXJQN3ByDXEJWb3lU/Jv2d/mTIsd9RmUE5I0uMj4i/Dj
d5YH5PTbOaQxHhw+2/Tr49p3pIe6E58oPTiF8bRH8/Qw8NgXTSrZ1gh1udIqdfoM
MHZGzi0E4N7zHAJy+X2YtDN5WkIe2ioEWnegWeLNaOcPmaUIpun9xakNRCrbvhje
QtGxMksG5Mkz352oiCy8m2yAG2Jjojssl+j+eP9JxnR3lbSZZlHyqIBiunYfNyCh
AVTMv3Mta3R4/FjXkQgS7eCCvOImElL9SE/hyzHDnqa1v88iomR0M7v+GvH8hF/d
g85QGA6QgSIOVteltbs5nWPA9SFIQb4jH3OdRG6mhVZPRvX5oSOHg5i1On8RNleP
TrZGXzjYEsYKVC74WUoaHY0n4f5ZUEgXIctHYFrHT8h8MycL6hRg7BrWqD4hfxbE
z7wbdPQkbXfH4wX+u2UGwwStpEJGl83LN3jdZwEiKo4li139bxuLaEKNcnz48CAe
n/Jc2ECcSMQum0lql1KbisKk/kl/QA+edoZwDwxSRNiaZF/FuXF2lk3nTQhrWW0W
xfRxA2t/fNuYy9ag6meMXyxaiVbiAM9VA1atyagANm63sx0B/kZEBC/jomEVy6vF
eW1ENrkZAJCBIMaj9TO/wZUMWcnA2AiFlTCAG4V8BjIpOGCxVZysDRO8sG6Z1H2f
ANQUVtNW6VS9ztaZlCv544JzdjopNvmTwm0ORvRvAb2CGNq2sGKnnZedHKO4F7R7
qh0NpqQni8eLZ7SfkfT64OT2paTPyaGvhg+g1LqVfN4rmNM34oU3bwYIj8wIREuF
lYtrCMOOQbr+2aNuD0s3WLY9zUDm52G/y6SdZcW1ZMx+qx/1UA59Kg3c1VX4TUQK
opizZmSrPABmwnXigKYp7By89hQFlbzT1Z5OwXlfTqy/bMmFAPJ1sjYslTLmuAo4
25rTAvrvzE/VV4MwfysqYVqeympOIdztObJLtVZDR8KfqteuiFHenBqCXjJkqg5Z
5/tID4/TIhGG7FrnPluxuqXt20p8767CmQAWnNbQm2tEaT70kKXwfkdnrIWGTZGQ
gNWAEah99Df3cUlCs2jCYZkJseOHWAMuCzYVYFv4kRZet6DJO2kNszLmP4vuciXM
udTq1skGvs+JDeoFDgQrjb+qAMZ6OKRZ9LbmwD1p/Ik/N5TJQz2iRk3lL8BaTQwD
4N2a53aq1IOm13996xBDsb8Fgx30c6EZcRLnHEHqCD0+mG5QXmtI+i+LGBHrbsMG
B3b5KDRAGsBQTJOwHKYgokX0g8ZoqXQCA/VZBgr7rzR+zTPAlv0fSI1K/hEga5yj
IPUNQ0S3kdd2V/euXTld47pDpWtFsi3SB83HGSYt4ClQU48zwu3K4JaPgjxxCyAP
mJJd5IInRni/BpgtmCNHrzW+sZuyOM9ZOq44DyBjq0bHcMzFnmB38IOCWOkNH/LB
NNrtFZC10jpuXIjA6ug6cMArvVQu7fMGRidFFN7jj2Yb0PEIP3oYWPDfF1YXSgvN
3i8covpJXXAwzYuXrOb2dAZUPVvpziJHxvS3v+BUZVjvfjsn2BtLsiVf4zfwwOyl
uZ8/l6DmTp6l4H2+OpLJCyE/nLrD3nP4gtwqp5CFU6koWFDrGvrOcxqx3L5TaBjg
ia43fwKuq/dz1ADkdb23H3U81n/NqbfT0T2gKswn75wqzCLTYhFybzTgGG6wHLAA
g05Zq1HcU2MjMlZJnPgSUTObcHYLQOwLj0wCA/T0uSlP9iDzEE9pWucU3D3GX3o8
UEepbWW9Wry9TijrKvTnLCCyrscNKkbibodcbtCpYdKOYxqVLzG2BiW6SHRka2HR
1RQ+PiTCAxJegDMHyFIE3uivhxWj073qnSZNgZcZso5ArVSZaaitxyQdYi8IZVr5
W+vRqhBbu0Xp/k34uux80Xh+v4Gr09mACPL4Cq6CxDsye36FzVxSwHNbbRXbqDuq
c5/3WScIHPOyciSujukpA0qKLub9uS0/hUC4RW5AEu1c+KrFkRMDusWMOKyY6dqG
r4lW1dPJFFI9Md91C0QZbon5kOE9HC+AGL6mv6tC8RwRE10MEWxG1IYcMhEYSjY7
kKvr8EzpHo87yD3QIIyHzn0gZukrNxq+Z27+9UZrajA=
`protect END_PROTECTED
