`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9YNVa2ReiwIgE+0UZDRe33fSejfg0cxzxQXLY45qwmbnaSoZws4ReK5cyRzpjNLr
VNttU2r0jrZY+nOhisoWz7y6HU/PCC3pEPatz+fSGImSz8Ml2vNRwrsEwKnmdUOh
87GVvmgnWDez9EJ8iriUqkXRzcX9//p8yDRz4hhhTgphdZZr/mQFEOfGGIQRseH+
ZH1rHTpYYsibnp7QeeUFM/lRsuMS5W7Morl6OwcjjZmJrb1224vzoyIHk8BstOJF
Tu3hzKGXC/gdCXGoqEKO7gcXMG1EVnRPGKiUjOBUfgmKBA6OD7xQE9h+Od2YZzv+
F7/hPzLIQeqEGId0ztKOWDamLS2gLX9Q6CZOXpD4zGidquyYCuCzQ1gA3Y04wuwm
Jvo8y6Rf1W88VkbnDcA7cfhp1sKrHbYJuznHYxWRMWWt4SX61D1crGGGUzsTV/aX
ZCHuc2y9oxZlm3II44zWiAegImi609bExdxPaoS+yfqiWKArkIH+y8Xwr1vsDS/w
ybYsG7niR3MewpQGRw06GFUGjVwYgUFyPvTDwrOJTvKFNenaCSVpkGDvybHPety8
FKQotKPLaVUtw4PYFpFcZL1foO4vnWAq/oyiCHjMYw+UjN929bJDrCGyeFSu2hP7
oNoNtwp0+2FDTnpFaEM8SoQ7kaeAOQko4R/SOWwHsypiaW1M9/T0N7/Xz6uRjAmK
PpkpEBJTNokc6fR4zMbCJTD2QnBIjRU0CCfL8Ui1jA2xTUeAe7hw/xskQ/PCHYby
FlCPR9pv8fDJ4NQTADAfB3l5axHoHaqgVizOroz4X/pv8JLek361/Q7geFtXEMhn
4xJXH3Nc4lk0ua+hle7VO55hQ188fq7pmsdSibdPjEG68u0Hjs9vBSsmiDUrPeRe
`protect END_PROTECTED
