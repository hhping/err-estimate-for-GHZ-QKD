`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDzOYQ6RCOK49lWKggSNDYgOS+vEPV2cTFW3K+mXZ2uz8bUESCJ+yc94yJbdMP11
Uv3jxKitMBK8Ojjg1qyMaoVhBFiRHEaX/cGPbDQJD7yb3tJtsYiUvuM901qyoZyD
/md0yOsrNCyGntphFIm29ysFpzbEvD2Mcg4ckZlXDdVVmy7sM/U6UoHcCIw1g1TX
MnKyJOH/Oq9e8MQKzb7ql8r1NoKqUABjuBaS7R3ckYVtvfx5PkinAZEOaiXE9cL2
fehbXSjRlydKdUVMlsaRuPhopUpUPsqOekR7NrdkUj3E//ORKKrV22x83BReWceb
Uxj/JMLPMN5ZdZ0M9XNBQUQisCITF2yHzrdBaZX+sO9i1vZaHgZeMCeBzf0dCx7t
xfcNRsacjSYU8Cz/rV171cFCVBFBID7gvwt1aVE5AJqHJTR7IkAgUsD09/lLZmLc
rwPYRw/GFFNBigV2iBMeZaIJMYMPJSk+umDmHvLBUszvKlca08jRfOLlTDVujsTN
MPtOz5GXd4RLlDPMVxZ9W4USwc3JmxjYY/ydHV8vH7FRBIBSv5b8hcckAd3R4xl4
4nSngeOya9lH90Thu6rap4h6iuNV2PU1BFyTaOXlrnx6UxI9X7PqpdT2iG6QlwVG
FfDe5aan2o2jJSvXy0sESk6LmdWvfMxws+zzUKxIlm72546I1AU9NSdezilgFPBp
UbEemv1/15qKcwj/U2HmHwduS4tRHckS7+ZESnt9k5Ar5rnfAAUApjEyicQ1FDKo
TTyDx4UvaBNOwSV/2mVuQOGdTiVRgHwgkEHBqRebPKICcRNE6o9GNDFquwV2t+Hw
PCrLX+2wqaHjmwUf+u0Z0ASou7WVCk30fH2pn8ML8IWWgnuDcd9C89nlcqWcwS69
DSezWO83Gl6C5K03d5mBhOCrL+qlkHrZSnchrmK/+lcXYgIY5WkLruCpj6yb5nrN
qaAXjtGRhaMr4ojFCv53kv2SyrGKgNHUmEgDJlDB7l/+wBCiSDZsUb2pi3i4r1iK
5A2lAeexoB09+gQZ+RHVWiGQa9y5epbwT9IcJXQUZxryTOOMVyk0gZPzcA5/oYBQ
BeOC8SYODDzBKFD6LHZOzb3ra95u5pTPPjRRq0mkyPAcZ3KKyCHc0YmPggPlfe4S
OhopzxvXF2hOm42JlOaDFxtuRarIrahoUHl78b3nf6whK1KGXksbk3AicCwnZw1M
g0ryeA217+tyomwgOb1tsiQKc+ti79KrjEFJZCH8IBVCjDTvzaY1j/H/u2XmgqVf
YB/tQoSHmT5+hK/K36/7wHuGnXd9MZwYVZT3O7d+E7wMZlden8Cid28gYGmFWqBL
sJzvrig7NGBonLb/SOI/R1o1lerbu6n9+ZzqJs2zyWg=
`protect END_PROTECTED
