`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNnjNWXPSS9TNGL7sB+T3aiawg10GS5KbM/OkOe4CF4vwE9FhDxO7Kk2LN9W7KQ2
eWTqfh42NjuPBELPaXH4RYBgxV2eKUy31+m6QOJ4HMkjZFEWDF2lnFIEsooZezFD
Klf3s2tFvtm8l0aNfZU8aBZ79aygnAZ9oz865ni0kmQHlqlNBR41clNk5TF3mJF5
dJMBPi5FUvzNruEcMfyxnBYKefJkQNLYWCokBBmqsm0x3agh/Y43V0VaZ1qdbxPp
tajYwVEoEtzX6iezHznKEB0Kq/MKySJgbsGmqQPLi1G8CnhUyTOA4S5+2NY8HW+e
Ig4/XoW5YvhNcFec5nsa3cLjWkNGafSqbAyoncM5YxfHkA0QW9oEy1f+ggjfjXkp
AKRJemxUm5eYf/h1Sm6NtzCADDOV2FalKHVs4sdrKXr3BZdhzb3Vh+LWXBelpVsc
ZF47H8hwjRWqCc88ncoXP4hxWCcSGd6CbNZzsCq0uBsaFwPvsl8vsl68wxCKuyPi
vkshzfa6z9g8mPKrEEmYthYjd8s2xp7Twu4W6qfdwW8pwMMAfVAvOvDhMIhC6H9m
tBV074AC9k9rgcquTWm2DPEV9LHwgBzsa+Nz6bbzw2ssvUrP3mSXqzv0nuuz5aS8
bUmIW5Kqp6wopup1UdEkoZt9rdDIs5UZLz1DPjsBNXbWWmHEdnRSSPbdJgw+q7Q7
bXcRfC/oaWAxPcTGtIfirwerA9SiW/JGXzd/uYAMl+dWZAiZq6JftX6yh5y0yh1V
V4kKbBSg7UiKNaU38BuzBdPBJtiw5gZ5K+Xd/nGZb62veVpoQ9Hxjq+93yfo2zwP
+eKOU/+sprqNR3AkO2FC5gJjLIAX2E4tAnxxRiyw1VWB8Sd/nyM2Yggg2I9PNABg
BWst1aXnknz0Ovyvh9LF0O++gS5rsYceOA0o4jzfay3ENzpcN6aYb68Fbvlh3G4B
5YcUI51jfEg+F2WvmNrrfmGUQP9e+78Zda3hT2htIc+n/YJAaH6dHq9nuKiEflrB
m/EPPGR58/fbxU+BdGCPxJHp9d+8yIxmQuW3LkOG2YHCo1g1xzKPdtyWeR0Orque
U2GagnqNqqja7fCPSMEowHxTTqAW4AEPEN6uSBH4IVJKxV7AwNUUQ1lrfb1/+7/a
1pwcN+1wHPpPC342zN9BrSQCNcZNOUXSrUE/ujzimklQzDBdc9rRkF6v8sIGVMAp
G2az8f3SDsdDCXSZemBknywMB/soHtHNeYEUpEHvRXk0XhQJlpzj9CsLr0IVOXWw
CV4XE888WKJVC8UWPnd1sEA0IPszgA+I07MFoy7d2l3qJO9dhWJ1qsM7KAsmZYEQ
O0iCkoM0pJjgzt+G9SrWPt6bIq+39TOpUakdbsIfnAoVGC+0eKNuS95jF/KiX8G8
HiANQhOxXleewVRSctSaanKG2JUkPR2SUQioegeqJWFBsbbREv1XB5Zn+eoOnTSk
1XNSwegZmWy8kE3Vr9f06EHelU27wf/fuqbIDBmMuRsz9n6ElT7aVafmzHn6IXQa
EzRFHTBHvQMObGM64fdhbBidXdEYkteUa9faJ1p8flec7nHOdCKXGYawh42sCjDT
CqKBAP/JSS12k+CJY/mRyZQHBPlAlAB7fjVKm2DNOlW/lPwrssQ8HeyhkT3iFVot
Jrx8T4fzOweeGLWO2LGstnr9y0tsPKal3D9EQBy8d3kdNz3+U3jcEQYN51ph3ijq
2Vfi2xyTTN/BpxdBY1g0NBVdKzYsGctIhmaq8mXTkRotJXwqACDH8GGdwsVSxV1e
YltDoE9CF21nDA4pEl04HcbhVHW7vZ8dDVFoCXep5/piBfueq+Hu5Gr5sWBAHIBw
/b4PDpHjYykae421Z2s3XG0hmo8aHnAtvQAFZiaHOFjYwo/kHYXb/Y8qwftTyDZP
3Uiuspl/SpodjMbaNZychkFQEn/ra+590wXjj9kU2jWx8fGEwKs/I9cQKA1he/1+
E3gBP7tfDnIApPaqlRuPLARvcANDu4/nxdBkWPDX1LAN3h+T7WD+IutnE2K4jPVb
jmgPaGkG5pprI0Y2saJ4X8Wd2E56uuQdssii5BQgWjHgbGXahebPWgXbwxQfhHPX
bW8rv18TIcz1mfZk2RtrgZrQ1RbnSvgIi8pSLhpybMtph26aergKJEQXLYn2q0GJ
W5I8SN78hYHATr8G0Eu9LmRDb2Gel/btVnA3KhBFIcg03SGBuIVKE127To8UvJZx
madIkWPFAgItBf6NzMZRUcoAcHXFYbeLwxXZdBtdSTvr+lha5qPwyXgUn3HQnb7O
a+IptDfn5E+x19X0GSzAxzx67MG3QSNrIA5LX5RloYfDYIJE6aXxLMh8O8zMRgQr
kUm4Sd2ZNp1rgY+XANO87CcOBw4xos3cUIyhIHRPqBgbOSoxUKUAwep/rcmRJTgZ
rICgZ8fvyarxlDY1oG9WheOgHHhgK3GGi5NXRgu9UdRr9heHMh1oIMJaT2MMayZR
l3OpKHYn+Ict5dxIjcljXb8VeYHuibwBYzQWPE5xgMyvrgKtSUb2X7NdymLy9nUM
a2mXUI9jYY28Qi296zBQdGCOsd7woSSkpWQ1+J9nr+ciC8Hxx92YnyHy0qoUYY7N
O2losEmjCJQliptTXfS4WYml/bY95MzbDU4BVZS6gbDXSnMvFHKhEifJoy3o0fDX
ahEEklkf0YIF9RYebEXVoE7RiGlBLVmeodLmsBDR10RGBWe4+xVM2laYnIS8hhrC
b3FV62TPEmiYWzj8VMhhB3Xt1b7L1k6qKR0GZeztiDV4dB6dCCuXHTBNtE6XsD5N
tultWEs0vbGitx6WmO2pGJYeIdZChJvBNVRsUGAh91whRBnRjk6B6C+29ipLbGYW
McxAu3loXAkBkJCYdPkW+dwMhhzhUKM6gad3nIKzJyL7TkUQ2ssN5WuOEFo/00nb
8WizPb8QzKTDsf7WZ5r1D7ATp7p/b8vPlYwxcuNrv/TnQOWFHzEu+tnxLhvuVtpO
d0IDR6GcObs++UOLqEGrTlZ61/U5AsVGecDtpuYdZjpTymeT7UoZl/HsTR+xFNH2
4YaFiM78/WbeomonvkKuh16wVSerabFtWlaLnRJYLi52lMxKdALdqB0Yut05LGIu
98yTLfcVVf+DBOL9IhCTQB/mB5KEsTClXg1TCh8Ksqnk+F9RSsgAEuOVR9bt994S
YfX7YkpNqQ2+rk+zEJpFiP60ENstzgXNwzlnGhkIIG/sB2u0PqYn+Ps63VJwHsmk
DBgMmzylcLynFOKeB5Emx830/YK1d/MOwjb+4BaRxSprCdR6bYJcQcyF6capupFi
8R33K0qhHm60oNubt0/tnQXB49ceD6UFqyFmvn+Fds8dYK7mCGich0Xx8xEzDcRF
/AVbrdG9MkjPDNR0hMVQgNp8Rx/5U+HTrR0bbMtNzcwbDkDO7u4usS6IhWezrOxj
mtU1C6oy9p0U5zvqw/ESyEyCutJQH/rUb6HGVtLYLyqtbQl05sLjEcXgnt3YUq2q
/78UvpAPD1PCSFAMCyO3Za6saSPmQG3QJ6T0X9uR2nlNnD2NeeNG0vdfG7BCHdOt
zlFb1ekUiS4VyZjzswVvy5iK2U2wAtoXMJuZFWU5qSiR0OMaCQQgYRxoxWOrSSuU
AZ8GODlQacRa+J8UPhROgdahsuA/OFIk/Fidgnv4tsDzt8w+64UU09k0qie++kvg
EWQZQxE0fwoYPCJZFy340C1/w1EU6L1Pslhc1rmp9LvvWZvecxgXLADYICsX19ef
iVUbmy5l/pq0xsr7KhrKz8gX5OYw4L7dGTweTMoT0uqh44QUiUWJBe7LFG6X04AD
c6xL/VqGsCQn4AJbXq3EEnKtnY0dBlEdi7JABJzmN0ZAEoMIFDZLfgbcMjz9/B82
`protect END_PROTECTED
