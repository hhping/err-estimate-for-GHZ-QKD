`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjOlJsXWunFPIbjKtqiI44t+gONzLWjUll3mQ94L/b7d+V7QHu2XMKDksn9MK2Gz
zu56zD/Juno+f3ebi1gw9kkVP+GIFszY1A0AZrET4kAe+56/GhcrrNdYLj9W/X6b
Ydwy4c0NgQqXXLZ5K2f67BTwV3+XafO6+xe/dIpO5pjX2G0IApZgmIVuEpow4fGU
a+d0IaLoJkwblGFWxpUbkffSwVR+Bw/vBcjBt8b+0cznpjvcPXbvYiPzZXz79Oxy
5M2ZnW3xVxPILrIK/SObuTZD9srQ3QXFX6uPYW/UMRn/7ib00g0q+FSm2uhXX32I
LCHzg/PvV7EXQaXD5Lin8c3LeGuapgo+XbCf1eMG2kqrRcBBIg21DbiIvQY8Pw+B
WW1znKBovED5fonFtU7Gu+om8P11rdiBLHtoeqxVsq92uIiY7FaQC1gTTDA6zpzL
1MVL6NNKvrcd4tegpYbOTG632UU1uxnSlBCDxzQbudEE/tYUDh0Qu4DJ8SkIxCcS
PliqRh2CXK/qL2oy42MP3wja6pbot2vHKnlCyuY9Nfo1+TqCbsFjGEid8l13rWGO
CJCqh7EAcqUS+2Udvs5si63IoBVAh/NFd3lobtjm2puBiH1uNjpPEP8MCDg5ohF6
wgf/nkErXmch85W97ERCL7ffl952L53eeRbZ+B6yeT1yxVR9iRYaFe+8STSTDSOW
lKxJpBUshtxp8mnP9pyU4YosciStTgE3kokMxp6yyfq3Kx6uPGBHWM+6PZcE0I/r
VIfwt0Qihv2B9cGpIn9A4MBj6WC3jLyhHFLhP8rm/G9vSJPxUOjXH8mx/oDu0jFF
JKHSKmXiFhjEMSIU4os7w/jlmzhp1jSCHSBt2cDvHSV9zQYofXvFB1vd+lWD95Ue
dJN4wvkx1Ni4BT/t84j+H1pVJbMySkY4WKOH0/k1crgcUunIBgLm5eysmoHBROof
giFaOidwAHRxZox5MY0jGToiH1d1z3GbJMnuPbvaXN0h4UUKZWS5BYzWGcmAhjPR
gRuVhhvKXpgPMnmKrN0VnjA9lC0bjDmmqkYKtQ+G75E89ttKm/UumijrF8xt3I0P
`protect END_PROTECTED
