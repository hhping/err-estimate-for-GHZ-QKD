`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFrzda5Tom4NGK+z+vdDzQ49bevw5KSIkH3323dRT+7B/a/dYTBy+IDXQCeJ1MDg
ItoHrF21J3/9ff9uXpjInXlfPrVIFzSt9bzakPdnrVdw5X2kOQkv2+ZE/3sU0WVr
A92VZqTo+9ofX/ABNopAdcrT8OAcTAKPb7I1aq2sj7FAnufbJ3ChIgidovZ68Hbm
JveezpsC33HRl10Q0yhOFs3cyNy2tQxOqS2wmP5FeiJQ4RArZVLLP7clunobwAaG
0vMUNVZ4HIGavh01BiKH5kwDdLVQ6AEBComp4NhBK6pfcOj35mMQrtKJeMgVCV6A
+he/zC56NjVunSLRxcRn3XxXK61tSWLJlMnv9bs1GnaS7XXAJf+l4Znao8Vc+4Ks
zApyEu617x/mKJO8l5kVS2zb/MkYeMVxMPBUfJY0bG+IZ7EfFSzGfThTPD3WCkgd
jNuVRtM7HNUDmuTh62dwYcceZVDuBR/wwUio/GIrb7mKFaRbjuEZLdzxuqlLzbSC
STnrPukDSrFjck/fi0Wj0u0AIG1SXhgB2QXfssiborakEMCTs5C4QzyBYkCnm1vM
KG7w5BccYg9SmPmRVt98x5Ogrk7+RJp4lNiSTrflLnjvny7yAQahxAx1hCyxdLes
85wZUUDChXXUfnITp1uFESyM1KMrnw+WeDc/u3g2VF1RAKMgBzjOqAZ96iNU2pxj
`protect END_PROTECTED
