`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxZ4dHXr7oPuQ8fu9/Vl7sKeU2GnajXxRI3nT90QJWfLj7YIHBDDH0+sfyPcnCvZ
4SAbUepsEh6LquX8RVemdfFRucnDeimgrqLxMv3/ER5MWZOtCRIQi8g/rrZce28H
F4BpP47ntL2bdv3JATUQzr0QeWI42Wd2h5UPimStWhpSggn613tnRTSN/84DhqtA
uGuJ9qBX+VEUGEnbdJjy5pwG/QFzZz2blKNZ6i6D2Zuy5ads8cqzogHq+7innmVu
oPS7kB0Z6QfLS3YHYVYB98vxn3VK8MYOZB2LY+z/6Qlrdget3Qo64Z5MNE6kGL5Q
H19ZnrTke7zNOevNm3CUFZztYiUQOYjfIHywKZ6zJGGc5vbuUZ/PyEiH0LvMuMdD
goF6nNfAl82RQY7nZ6RIZyqHL6iNDnys82CBWLWT0YGn1132f4YM4baPwstkojJc
/zTmh5Ozea0B6Ai7Ho9owGvyyvvwfmZLT+Tttf68Y8Qb4IcFx84IFoTMrroqsgWy
XrMd6X2nI1wjEqJiXlcED0pKgU6NB+BvMPHfMJ/fj9cEFtlnrAeIAl6QzfBWsY8H
UaRme4vLVDMIj+AuoPzehpwPVhyGpi0gr5JzxRKdxleAwYDtHjb+cu5TeSNbgqgE
diKtG3PiOVZxL6UMirKvgXvTMunJZtYwbUZEeMQysnbjlkpULLc+tGFdXV3q6qkF
g+dY5XNws/AYFcpT3bYim+/Gnfv8meN90l7j0wpy6TzzL1OV2yuS1671mopnzzdu
BY10rZDeDHX8ikHTco8IF/JbKSrssl0Uwa7LSOLYjUklnEq6h7hHC0C2u1MKi8O2
tFVgLtWdum7yFZGvzctd1e98/fyVlfmMgZWFbF/oIHVRQFbO9zESvfxmw9t2RB6r
RZk254qwqwIOsV6p4zHoe69K90xUEPzi4odqSW8caGtXR3rsrT/gL9rzF8dstXpw
IbxyXhHVtzZXLAguqqVG3yHHA8W1fTeD2xUvpvtHDXoIvRwegmRt66dWRjlwfG5N
wU3QB4ZOvAo+ukk9z5/GKYymXkgYG0x5XB8Fkl1iH3kiKibaN9CHuNbQ1e4FHLeY
BDfFCaW3lH1CeWmBFDSIyME0JA455ZaO2Xxa9ctgEh4BCKtY2RVrcYZDMEjUDO4p
BPhwKELgox9VyAExW38z++rS/7MudacQ4ZzlIm1tudkFboTzQxRcnSg7FuOayjvq
yQNgXDw06xaHLD0gep7CO3kRECDYRWl/Exp1iaLq+ja7BhEWec6k0cUZj7dNuSdB
4n3ZSPUCcNOorsPc10IqpVhepnDSVF7MNz61yfsIRnUo9oEgDx+TJrFNvl73o4OA
BjiEZejVQAjdcjsri43+h60EFwlyePAzkZk+nBAAgtf5YI35onK+rhk7ubDWOrVl
svQk8m0R303S9ju4Yxp+ZwjmltszFYAcjH7BIQqsB1T9QDWZZiP8Y9ya0thy8FEo
ufzD0rOS5IclQkgbLSfs+CgkMstVx3R8oceI+g45QUYKoLh/5ktUn8NoO9Xbf9xO
/ZX30Em9wBexjw1i9VwVQryIzS0ohILp4L/rt8GvwLU=
`protect END_PROTECTED
