`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2RsKZqfPrK4jFxYT1cXwYHtAIbkSRzNzia+HU+kzr67kmpheOiRkGMiMjjC7ScMc
tlvLTfzmOHNpOwhN7SticRcVjapas3tzE/YFV1QkkZMO3yvxbMU33FgF9Othh9k4
CZ6LU6aYgRipZqnyvHvzBOZXtrfHBZVBIswXXWxQm+obt5lwAziyABzNFoD8Hazh
1X7PnIxddRzAwf0mn6ig5mYyV8Vjht9byWYNaL2sAAnhLIBaaC79dahvt0PryHzM
sFCcaw6tCmBShwxXGe78W7X9s7qUpbju+AieJAxwHpn25EKYMO3nG2WI+pdzyjOa
xtqJuVsKkIGmDzL50PSghfPMkU4VX2Zr6yRzzCnri1EIOk2y5tNoCXSfgJNFW0I7
abhCS0KOEaij7vjtX1+bzXucFSECRPZWbdKvmDR2Rijz2sb9kiFJ0oGLJ0+8lptT
uyH8di5DphOAq+o1xmny7AGc2MeFQMPTXQEeCuXkTDb1M0qBV3WqmYTInRlb7D2o
`protect END_PROTECTED
