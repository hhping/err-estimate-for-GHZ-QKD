`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iHmbPEVJGa20+mjvfx4/AATgDk1otVT/0L+X+mrNlmdBsEkxch8KlxihZdmieK3Q
iy7DPmnq1APB6V8+WbtAGAXih3tWYuCejoS9RYSRx+pTkjc+NrpXWShxmn+DqUi2
/eAp+zSVP8XsWaz2OhE2qL4hG2ft/K2X7Y0+AstqmUPkVMHIMk9HKp/qKcakDaeE
cV4vhWeLi34uktiMu6lvIbY3EeeVSU49K0O2tiRRgBEYbtLWju1bsjRqZDAL/PYx
djfUoQOFn+GTxudZLBKrBpsKW5tIx0/rVMWk5fhIpTWRZVEdL2wqaLeKpLn006yQ
nv0T95Z4JJYZe90+DbYRw8sl4Bil8mSks1N2nCuFqpV+PYvjI6cepASVZgryqROF
tEn9SU9/PCreawMPI7+q94IHmeknpOK39l5HAa8BguXTee9BETZJ9ziIViKyaxyh
M41fjCS5MhjJC7R/xmoXN7XI9FP7dBELPNINygqacB49qqEcvrs862VnLbY5giWF
f7Br+e6FItFnB9UH0uEswFI7oal1w6INMrOlfZwUYcijS6qBPmEgsadL6cvdEzcO
ky1xNm+m6zplFNP97/0Anz1oge7HQAAOmptEPFxLpuYaV0qG6xKrI0SmC/NzZ6xI
UfYrmmQoKZRzIvjGmcmkypLLWnjc2OcxY676YmbIG7TJHc3mKu6MVYb+BjDLAaf0
kjcZw1r39hVd1jhn89Jci0rZEyDRiNfXMcAwtRvKKAPBPTI56G96RoTXUXFHu/xa
1QvjDjHTmXFa0zXOPWSotdZdsxchjJCZ80uaUcCOlv4bgMghMT5KI0DfaoBqAmKp
Us8pc53s3ZWIN35qmLa30r+1094TqCKl5fH0PBObaqZt0uwZl3RKRCPzmcYkCyGg
F0VrjpGme8bpN6cbmxJ9Z6z1qRvJ//PxpBWjfyhQ/GxhylLmL8QaoR8LKvVN3Day
3hd16038oEr+m8JQjWLYvKLT0s+rJkuIm+j9ZCz94ses1sDqguvES95+bPfmsbrI
gHvPA82c80erW+15bdkLh7E6jt4hr+TmXQAaHU4+UwUYfTfKAH5vpYBiBsb0MKJG
NFRTI0Rd+sH1iUYFLgyp0fSiwdZ2nY0RBu6cPMttiO7c/9Xc4qmbKQcxg1DK3s41
zUYO/0w0X9UVlss+Mnrzs0LK28AnVndI1qUraOcH/Dx0/EbG3K10JIAt4hxcDqws
E3VjrbJef1rpDsd1TD9eFB5u1/iVfPfSiDacBDzZ13EB85ffisJp/e6iKygYmVk7
MI3+A5qYIxyBSQ+8xxvjTdGDjoxE5sT3PF/3jf6dd7yUzJ43839SIa99NHBS7XI6
uChHVOZ3sllIAJOzsmsLB2/pOC31Xn2Q3BKdOKEXWKkjph+9OoXDaL/32+2nFYkN
UQL0TkNlaOrmNUJVvfUPZAmttKwRmOD/UNhyXxoshHnGihqWfXQXaAjc14328B4G
MpTNe+0PtufWKv1Z3VwVXl3swhehNWqoKRxPIyN/s0mmiupQ2GgCnlWXQjwDx2oN
AYwO8VFXY+IDG+CfdqHuyrn5hA9RK6zd07NaA1Q5n9+bt99A8z2/cq93YCJkbecG
JKjW+RKxdJ52pF1ygnRB+dFfdJuJrsnM5T8TOrHmrXMk9vTKmwrXqY4GM0hSrgRG
`protect END_PROTECTED
