`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rWpNsQdh5DiLAW6Q25wlZ00pwA5qkyLQKrKMkEtPlLZFcadGvqksS2yDlA43mLTT
myclqTRjmW7+xp3R/a+u+Gan240+kHzt6xAQcvsFG1nV+TLUPhyQwQaYItUrbQIQ
DCcSGroSVRnRazURebQdOzQ0ISuAF5oJekd+T0442FGL6mg/KjU1BogDrDlYxYfz
9BUm9x9aEinTXGhg5Cmpl0myXuR8Zea/YC9JxvaFK0ptVO8mAtlwh1G7AEgCaxsT
kAqVjI4vwGlj4+hkoR8dxyYTeJVrHlhBKLniLY667vRY0XmTIaCpLQGWWmTMkVZ6
hJvTtq9pLUyvl9GnbbD4Z6tHfNHOuum7zagMV1lLR8fh1P374OEMFFmu1b9eHN3O
BK7/AYhZ4EGRXGickx6se/p7HhLTFgIVUr7ZqY8nh3w1vWiGmAq/5Vie1ULBGXdK
YlTbGc8P46NGObJvfaVvqZxcQlSGDMwLV9oBmWtifRVqeHEhR5jVO/gI6YJ1AmfV
ESiz1+sOw98qLB+3Lv/DnHHWevMRejgDr+OAB37xKEYg6B1tl/hJb2QniMpg9ex1
DIUKzkwLttAFck/qn7saFmu1z8UQ3ps2b6fkpclZQBITxGKhMW1pIHgFouZI7GZU
s4N7GuHxa2tagqqLO5H3c8Yf8KzRn9rCaHM4eWTG5so=
`protect END_PROTECTED
