`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nKdTf0pC6JpfdujwsYTmbXW2VSlarLGM+9y5sPjKziOVNQwXN3fcTVjdlIZHTMp
/L6wEzzmfsLT+9KUPQgW5WA281xTYZF64wqHH9NPENWVz/4cGKa27U3AP2qsyZqA
FFwDoaxnwjRIsVffDOEzLGWPgL9i9cb8zhMN7KBOY1QR6GY2LOlfRCmvDXoSCN7k
iMhXzIuNL9yQKpIVssbhvu1iHtyzwV/zc/7tdHtJUKQDZ4G2GP1mQPYv6z7r5scP
9h75A0IiBLbn/IJKPAyHTjFBKssnqih7nCFpE3hQqBdtseKbWtO9rnpFI39CjZi+
KtyKZ08kAbkn2gZ3ll0dj8lv3lFQ0tuludzypDQO3zzWF0E2q98PFufPg2bn/oA6
1+aPoGeX0+TJgSXyLzpg/1hUV3CFAnuhURcJsrvkzvmlNsj5jgypsU3VLYdCOhFm
kZBQCiDVWw8Orn7sw+2PxXC5uo3Kpx3jvxMwr9mz9TVq+SANm77yrZJGULn+VRWS
UuUEd8YSq1dbBWkdJF1wNTCTEFWiLVEOYUGaI9m2/avBLdsvnoqkOCRq7DXvTsYP
BTjZtYTdYMfaEh/3opmoCcDwLJiPX/6z3RneMnqAygGzbsEFKQ3EIg88XFLiKmix
up5NIHXZuz2AUZRoL+DBkymiYQQe+sKkHcUqJkxHjKBOpyt43mTB8pCRuNxSEj77
DHvpgEKpGULJZ9Y5HhMV6FS/O6mdyfiqWdbSlJ1PMhak5U+YItpvgTYrARRF4aHK
4TAYlAZX0j1GILYXDzvkK5qvedvjZXYUzbKHX0Ou/s+d6CCwtFRdM4hYnqOWic9X
OTmoRLYzgow6rbUwnJsmy8x2uaXCH9LSXEr3HXQdFVPtlgyghWuQz+Beehex+yrQ
T9UfSCwUBE/mnl/qS/6f0nnUQ72GhSKjK+hzpfFMsLfjWuiGDzQDw+IfpjRc1ftW
R0ZzU2C+ZGd/ZdX1ackcZlVjvHi7cBDBh0RbHyEJodCO9sNa6aCDiuErqFQDj6tq
RF8DNTaE9DIG84dhjCqH0mAOXwdNvkQh8RknfOUXnx80T3FsztYKvdbcyFIiIMVo
a1PYpKQXBa0KcI44BHS5iYi+dxfC6mHmeXog7DjPRxFu1GzGDRkMLQVrzLZdJxDG
o+RY2t10/BRpBV2y1fbMERGfuG002B7yzaCBB4UEVLlXLD9cNRvHi929Xq3cWcEY
Hj7mAJSpFsnMSkv6xvsGpXa03W7RGKEgRSnfyS2VhpyKJpOy6UD32Z1pzVM+NTru
mpsu6kS1wt7OnfdIXGqkjWrbSkcDP0rypP8B7e2kyI/Pjo3BArw5eTvbk4Gm+0bR
Y1SpVt8F5Gw+EvVG892Mf5pLA2TRZvVXrvu3RuNsQJHQsQzJbQxVTic8fu253cuu
Jr9aXrVRx+jZfpDbaT39U1B5yLvVR5nIseb+jZ+6aBKFogTJ0RSzFxG0Nc7K9cgO
K4+JXSJzYuBqRXTdVYRxZD/5pPRz2xSUCMPOenKKhnk7MnWONOFO2H7u5NUySLb8
WmeQlatnHabxZt8quIXpZ6Vsi83KCB+VM5/7pGcDsJxnZ/QG/+1MA8O9psTwg4m9
PhmMnBGJ4pqBUbZ5ATXF5FQg+ikhpHXPyAIYVlCu7p4U7wkD4oI0rNilxA69YIWa
Q3Ul15xlr9Mc1EWTRsjVWVop3WRobi9c7FH7BPd2C4Bkrgu8IZQ1owggI7aPY/I1
2NI8KDPByi1kX8CgSf4sjtagmqdUtBSrKEp/iMc2kFOtbR1y7+DOGz0M1G0VwPfH
r/ZbMMpdIgwNPb1puNhj71RzWXJuAx+XkytVnkQ7gfmDWChmPl4Z+CNYWK0gxwlF
kqFDW0K8EUe7M692bpqkS5WHtBLbjieAIHnmDWuAG2BFTs77p5ANxUSwnocGpWPZ
EFaK72VpMXjVQiQwz8bmUyfYdWHT3USnb56Fc909sNlWbuI1f3UQT72sLLd1S3rg
vLnfEgx8kAw9oMhNw15y3FrLDuNeUFzWSE1SNaCCU3o3hYvBdqSmPBaMTRJKBF/h
oCUoe83qU6SKk087BVXe3jJ4hKoRC19uaDGZq8XRQ0e9EcmxR35ru20AVYYrCIP/
YRfQQrHFwHYb7Q0Ih7bvMEnSQnBGQ1Q/nzeJbqAQqMFrYc8xTarhqCaFE7KWTlMl
8KmimZfEMs6NX9CndAjyZlKUZWit+W+PZTH+kSCZxDAIaX6Z3Q5NHhCPoQTWUBdE
rWvxWWUM/AGCwnqR2qIM+u7anMX0EK2IsAcGBqnMa87VPwtpkHaeJ/RGyJBGjJ7H
NQi1NI/QO+xsom77hpaFmYcvb+LuJpxwaLfO3yh39N0=
`protect END_PROTECTED
