`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QN0Jh5E3lQALlJXacFLpjly01GZoQeqiBKbo7ZpvX+z998tVPW8YOQo+dH301Skk
rFQDMmwV86JT5jk5bANhgv6mq4+D19u1HGZ1x0BWwLOARd9+OQGmP8u+f+iMR0mW
VYVsfyIu4Wv+6uafClcs7BMYNqwdTzN2ktGd3LA6J4thHn+0Ygw5caIoxgBjrygQ
soZWxC42vGKNGkYBFRwBxex7JRB3Y/k2ZXmLra6DjNd+fM0PLaKZE1nPWa+6nMq5
mhlDoqZqxG46BQJe6clw2f0vtz9gRySCwcYgFmiU6wZxuw+CBP2YKAknR6pONmhJ
ttBAcYHi43wQ8BAz8RJxBMfJ6bMiidk+CdRSWWiQclleOfbnOW5rKJOR2qG3YP34
MlozfNCxvaK4GhJpheH2gK3tTcPaqw+VPeqPQKPv77DjNfC2UsYjbxeMtpe18hlq
crLPcgItgalkqxoZP2Shz8nMWeRycHvQ1+elGUXxWL3TECm4DgyyxhhTkxlv1olQ
YFrvZE79OwkxhwQjESKF4MfRwzwAx37XKH/Ur2xM94ZJLnafkvZXK+jX+MNCpz6h
khLXG5/hO9WVdAGOs33Jpg/Nu3xAlU/8owMyVF0DXhs3NH6sk3SkWxiWfshow7Tz
vMmlrm+MhNxQGFMV2C/FUCF9nHa7+byFVkolLT4OCN9XBELOguS5a6pRL1WCOnfK
sSMy4pLmHIEDo7X4jp/qMQBHFYdXMX19TKOJbXlN2+ud87gB3Y9nBX35/Tme65TM
CrtIoruIwSyzwhOMlC/4yCXlQcluhp+E7pA2psLVctxG+OKc+LDPuSVLcFR/O49+
HsiOzZ1g8dQqoyPiFueTB4A1cYnm5G+wffc+xJKrZCNvwW89wqsuFxeiTxaGvU6L
t3bg21+HF/oqHIP5YQ8vD8rX1EiXNj1SJRIGqgMUGXCp/aSfnVkn7shni5ayZfA7
pUyBZym84GPyg4axrFiJg9nEcrO6s7GvcESZUQI+XZ8Flg6bbCBIGobQdPIOtDFL
L3PYeKCD3Vj753Xsx4BrEVwT2BGpmHuZ8C1oT4jDUxP6URQwa3xkFfeX+DeK5jrT
OItII1EaF58OMKy8KEHnWWg/zir91/JUJOVwdNKA7BVJH0/DfxZVM7VQz1DXP/Pc
H89VQvp67Il2V6FzaIaKwjZCM6Qqmb432d3XZMFAeqsHeDPbYSTvtpykOj+kC9F4
EpJK76VanrgjQZ52easvdzpVdVNP36Dlf2EC2w3vQilU3P3wQpyWt796cDJtRFfw
lEk3Q1Bag3GhnsVMnbGQMkmgzzgAYk1TbOthLpwRIiHZY7309kXn3Bxls2oW0txT
HNPs3hO1nYBikg+2ylPiGS+Wz3J06uDdk670A/Ny+Q7yj92SnDr68aBJ9D/fAc9w
llWZ7iKhfoyldMiXKEFmPT+xOrNJ9jxVM6dltYV3IWf+wB3yCuq/E9IoWxe5DkuJ
XNgjhGITNYjPad19ALpadWD5sutOUjeTx0QXwE/T9dR7XupsEbkAqcomEBXVY1Cm
AfFU0UKdux9ywxEm9s+to1YnmKWI9cKCOi/arzuAXZGbiBqEC+2w1BG8+U1WfDuR
+U6ntsb880t0AwIFElrv8ZKFmwvgPz+UP+LtV7FPXc31r6im1YrVKPGJZY9RVgyy
/OT4BNMqP15AhhDSuJlbq0Rms7FGEArEqEqod7MFIeHYMjf0HzeNfJallh9xBOXy
56O4WXVCX0nEYsPfSdVgEGTdSUPhP2h5WQbXSP7lJRRqlstIow03Kqpb+/hZn3zk
/8durTDVf1ksAIaViZjwmCTASQwa6jGOkuYpL4D/DgsHFnY7Tzld1622qn1JRAcy
cSP74Qu4/NOLzQqT9cCEqxQ3wNOyzKj5EUE7OSzDq30GnKXl7XeYAIx3glO7sQAu
DVrPUdqbozrRftoK3iNU/8LVxLaqN+H4CvXFx2JIjx99xeiAHwdHG5WSmCvUtT4B
`protect END_PROTECTED
