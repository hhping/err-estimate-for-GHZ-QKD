`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BPOcwR/GgzkTGBEbKDM8SNpPNWidXqwTLxT5SSn0J/NtdGGEyuQeO0Eo/W3kpYFo
y1/RJKUX/PxFK4AdzAPs9S8uCH7n4hFeScVqkskNJ6ZqTBi7JHrAoq7LV6Zy0aG4
HiYIkDjaDnGt9o79Hiiv4q8iu30H5D6hJ27yUSGHi6gtA1OJ+eQTpkzSgn1H0WR2
X03nD1J+ed7Qrq/sLG3G2Vsc43xxLB3diSt+6C1MYmmq5NGnP3lUfG/52Ch0qHMI
hbcvsKVBNZ3p8XNF2VCoAZVZMIrW4mWxLK46TQbeDjvQIPvDjLDP2xXrIH4qHwI9
B6ZnydwaxmSnsaEfWxUA+9XQPp5E0nfiMR/x8gKXbP2XRAuvbb9/nFNAvwPoMjVP
0P16FNWvI6ZJp9iOVs/GsZQil1x0Lqvq+yIOfanUlCmhx7T6IHPX+oaNO/Hvak8g
JQAP5OQjg5wR2NChzrQjVLIRkaMbbnXLiOlVY0lJyrf9EvZiVC5AkNMxpx/dLKhy
IMKosnLrC8CbeBWlIeTtPMHCYg1eL1DuSDVA5ecQpPtNXE65TVFxCOu1GUUaDwCb
elRVZiYMxddtq9yrWmHoxOOaRuQJOjZxBNufsNy4o0UJWXAIT+RCB4nTVKWodU86
c9eeYli2mIpYZ/FekezgqN3ocZYU8lclDfCd9LFctw0etYUiwiF0uHwMoT1NqvMk
NcuV9nTzyfIxUCWVtgfLB82hkcAYPbWFMq6ElWVoUDBoXIS0nTOLKUd9/YvXp8Ik
pVAsTDkOhNXId71lCT5vEysodjAEjF7HScvRBdrwWG1E+Nvdpj0VHcES9ULxwxnI
PIyrYQiYjRoS6UjsRbql3WHdeerijbMzxIKTUCeiUWn9FnVPMZYUFCZc9OyjE7OG
0NL9NmlbpQkWWFtWeedgr6OfX/gcvQkLyadEvWFI61+olY/9O5Of9agG/ZXiwh3r
Q9nJIrvtRj9ck3aQHY1keoFnJgZ3MTuQ1z7hfO5ErKMBuehWXoET1xaKGcp4z3KS
iIQbg98xYSm5JFo4Wb9g0ZbYyZ79gK6hbkigahf5Lg8xwr3MvUHN/qa7cjj3F1/+
VWBHgNtoOro6P4XMXJ5EavhuzeMSvYXhl2E0NCp8JblMd367qiTIJIUSQ7u4o9cf
dKMsDOVBt6V+W6XfwElmlt452+/vBCkbIg6e9gRaL0cX6qzbG7txJa+8DuvAnldu
GLNjDeYI2AuGGEHxPBJhpnBgcRa5IoICqlr+7TbkGBILeznbtRnQLNDcTeA3TUmE
KZqw7OMrR3eWfwN0WbtBmzthjGAutxgiqPWZT/9zwQd/B0rEUfDHYTsoT+yCa2wM
ck/AY6lghQEP2CiSqAbnI3mLrMP4lrhQ+wohUhqvuudvJ1W/Vgf0lVhHsj2AuSka
IjtOH74tdHVHHq4ARQB33857N7Kf5EwUu7y0+4WJaENgIlIZ0wTzny6Kf6MG81S2
sNVRUpYOVtqXFXcuTZeVUyhF29Brs8nz6WAN3CGdNQp1UZ/tKoe0mUJh+DLv79dC
nrew6D1oKoRh+wwB5Gc41zfCBgCkm98RSF+CN37CxoN6ru99sSUaBwVl7g+qzcRi
PWY1nNL4dGtpfkIOa7d61SaajqWwnASVTf8WBEkjL5gm+SQUbveTYyOSq3qh/Bu/
P6zDEp5dd3VLGYyk0zR0Ijyhn3UPnglQnt7jXg7/jjyikyXwvvnBNs+P/fPJX3Fg
3rlpy+kSCuLrSU4kQMzUJI8xmbJBwRGdOKFrdSh9zeFgxgp2Zh9gMQMS0owZlegE
JC8KL2UzV+W+EvDgN6FFohPoS1COnKzqG1fLOajw3PCjozZqfPSXEClehqr7OfVB
QzfHDtPwjYls6/wZCEK277putNV6C4PqgDHph5RBhsdMq7fBYFevLx5yTzLjzxGx
0QF5zIPxQ/4fIZd9FWuphxrW4qYOgyA9/+XWDUktgDd7u6tQc11CjRBU9GWT37K4
TRaqprxVQh4s/HggBWvJQiBFLpB5u6I3p/BYv2o+sf1XW+Iw7WQwmcKz+ke4hfta
a2UD6GHV/dHyv9gdRvKToURSifnOgPxxqRiczobPCTXXaSM7i9rCSKebeKzF5ZJu
UuNvlGpyjoirW4iB0S3dd0qV8N9jwEq5BD7pcCtDtE/msuf93EfzToedJOC43w6A
VMbl8pPgWabAJwRniH8ItJ5/BndMwDL6bASTeio44HllsoYRLVQJMZvCn6u9DFUZ
bslDF/sSW0HwXwHGVtt2AuU0jVNTo1D8epv9lAhCwZf2GZKLZJCRmt6mwJzwUvKJ
AFkWzb8vf/NAw0Pnzwkxl4N7ue+babac2L1pKbQIAHVOY48WrAEhPYMR4AXvdilT
AVHnMHcesyrG6FY4g2wwkA3+S5OheJh/JKiMOEx3+cjaLdkxSzEEsy5no7nCwicG
JW8BWc0vxnp5rfEVHxr+eYg7+92Pd2igVbVKFFmY6yxG8PWh0xUC241YYoi9YDpa
4rcqKj9jKflB5C4pLFf07NS5ug96nSiiDNHwJzxDs+JSSPYeZQRWKWBdXgAiO2yh
gQrKeWiseXmJFeM49EBw0MqyuTHoMD1f8eEdlWY0X+vTkW/RfGLsWxgV8nlzINlt
t/F7QWYBe0aA8+iTxVo4cJD08i3eCHr/RCUAw75tN1wRnv6fOAygHxhfO9sCZmIn
X5EZL6pLHe+4BJu7+K7XFxomRQXVav1Dkr/0fmhPdbk+4XUPlpbUoZQ4IccYVre5
13N+r9fzvyRJzGpdyWnGzGDl6PIPWZNUioyiueY8aFLD8u5ybGwc1ggw2X4RsWG+
wutXfC8AYI1z4GPc47XiyV2uI6IyxX2UiN1vQ1xIriiv7B+yGc62+r5uHnkftWR2
X9CBQjqYW/de3jDI5KEF0tAo0cEydqorHlUfgjIfMWrG6ZWpV8D1ELqT0SXNWDLT
CMAaTHlcvOMdfnKRLh3Pwb8NvYyWiSlThBxtX1xuDrbkzdSBJjnY2Qf9VLUKIqcm
UDiO+gMdmOWFOvXAi8kS7fMKDLqNlnI+4lY7Ozd8ZSZPQQ4N2YLh7hua9+zAIvma
TYn/cGM4ZYUkCPJaV56qjwhqRhEASGPUvRCjMXNF1iBrUUqw4k9sxSs1qw/qS7Kx
d+k+OW5O/YRWejYSJz8TNixzqnW83Iak7Ek71X/cufKD/pRLzIMA95eZ8JGz8JnK
YDrZZVlnvkYzKAqGmIu0dN4kFrWDeIAjnArGiwIJr9DF6BCAT0owrzvfmnj2qkFb
I6t2U115pFl59vxXSmnu0VBJN1xPRf2NOG6VsutZtHEgPw4iXuQF6V43sxB0LTPX
ej1ajmXFsAFkO2nr+qK0ugrlmbEF1Ocxuxc9lWIpaoi8IP0qRdkF2EX6nZw2ueKX
rDpLiUevml0aobBAagrF011dC4RjJqSvyUNcauI94PNr/dIvZ/eGfqLPxccIx+g6
gLdm60FXlccjuQxgUne2AbmWqa65xsepR8lDYngpSAfJAaQLV9Tl+2OheX2eREBy
JvBxiVVzLZ6nQlmtUSwoYyiJzBuBcc26QDn9hb4DriE+LGNJ1S97MPMLuZAM+brt
ufxoXt3rSAQ6P1yCKO/YUQm6fKKH0ZR3xkT0SBgvjwM9E3Kx2jQLFHnmhwAgxQYp
/FkIgCB0VN7Zpx1GWIkHqznwqsV1BRCW5NZ3XMDdjoSTaGfuIjzzOkNqRe0FY3JR
/GuhAY7OMdZui18mMf3Bn04C6nKpFaaAhbPsFCsisO00MBqcgUypu1Cr2RXotdON
Yqh383Lm9+7t5fjNcOF8HMmOAywIH8BYyJRBKyS4Nw2h3bRnLCQaDk6HbGdPkYBZ
E9/75ySaRh7HOdQpioWLX+CxjUavZv3LfnWqHXt1VtYzQhao0Me3TxyTX9rLP0eQ
VSr9YtD5w9j17dSaxC5tQgfJBs1FptT6SUD4TQOqp5l9IKWHpHaUTgwfOAxPHxUi
TCGGGbSukVxiSQgCGG4dr5H+/LBmOsOtB6Olb+c+bSjL7+EXHBvi5Zy6yi5u5id+
50r/ebbg1DlnLBv8bEV0elnH1+09bV5EA6SlNNgz2Hz5jevrj51JoNFKPq3Gg6Tp
q6HUol2NlU8Oeses46WtIJgNrhjsBYRDbZiaHfr5rWpASwx4k34Upv7W/s2eVY6s
GoI9Yn/EjE2c7Xp4fkhCgq8NkRlus8myVGpyzj1nLTZuMjyWFlTQGulL3Zmn7Rdu
CzYUHi+fQg4eW2KoPStQZiQNExFc58jTI9vbGAqez/vYue+9kP/o8qKKJXqKlx/y
u/NZwk1h6g20UteyXe64rII+/iyLRPMmV8vRbijmSqXUdtcCba+fGAqBCvSSyFDr
OE5CG1au7JHv5+BmFEUhC6DpFYs0NqSHC1s2Bztv1kIPYTSSrLIBj/+Xp1w9Nvom
RcAllfKXRGLa9bXPwAhvmEoYpal22nmfp8EWl3wsX2/dKb+dtW/W8aSQ7yQrF+S7
IkTXzv5UP+vfO4OQoRRoaOtNNweWAGAGpdCa/62V3atcmW6+FuOwaSIOY0gnIKqG
1bg1Vlz1mpkI8jLSdutQVasrP1TiiOXGjuz5Vijl616wBX7JoMN9gie52AQ/ZYea
Aka9xCHnXUHfLIXA+Nhg9tIRLQ1xsRhwRu9bmsVDmR+Nk7XKCVZmYm7hwjjo4jlu
0AlCHboa9NYIyAokFwb1bc5mHKVK8QJc/Y+fiPX8+Yw1ZqdZ03ph3Tl+fGd4Jmxi
hNy2LLXUkRMXGQsvnsrtX3FAxsH1PwE5aoFVLulKCyHqQTwd8T0yGuiSjhck09Zn
ZEyIPFNcHsAV2pRT82VUZ6vmCwOdWjQX10tmeKUOiwvjqyEKDofDHUyrNeMCT2Pz
540gmnXgkz+VY/Y/+ncoU4ZkdXExZNq/o3zlBlHN9+EnEejjh8xDpbUFEEhG0bmX
CHHGcAW2ql4W5m4oGyerCwduD9y9E+C4rXJMinIO1TVGiMCPSQei20kyHxNxo1+d
gpuh5xfOPgWv6WYg44wAHUElLl+zSlX0N5usAEt3wAx+YdOTQkZ2VvMYwi3+OXzK
BKI0nE4aLHK3WT1d2LqkHpJSGobftdNwyo+uHzOSwgKEMrmvcdHJIYtdaFRQBoEA
7u1wMKYnOMV+blS5g9Qu1W4Omm8AANTqunQvEM47uq6upYY2ep0aXDQGK+RPxWEZ
35SDSCqouFJ2aHhS8t05lF25045S8tlhpplgUex1/TpVMqXEb52GarcndX+2SSVV
AKj1LvdzIfxwpO4jb4ZJFVrKN3FEvBbwApdWXv2zQJoq+vMz4g37l+oxmskNLUcp
5PQAc8hClm3g7rUgMIi8co66jfoh7+WP1Su+IKXoKSCxSA/w6MINxH2Y8iq3plDq
nfZ/ordemDExgzoqCCefPdERTDA1ef816Srv86Sl95Uwox/ryFMlUDfSS39Vxp50
O7rkh5Ue7oBRC46WuMFn0kK9B7QZt/fDhK7je6DzZndw8HAaHB3siFKZJ8hvKIUA
ZADrboK5UsyRIJMAcR1j+vF6cZOLPxbbEQbBbZGi/IiBD+FXv4mxvU8vmMT1Xc5i
qJ/5oSZGSId49VcGbFb4iBaOV0MXMKftSZwZuoHjWVBtHWNxza+NN/KvpPkdia+T
IQGKzdAcICRhQKkYJju+4pYxmQYQun3lQNxi7TE3r4oMFTZaWs6TtQVQOO0D/TvZ
ibmiLQK9JaolH8rXDlmSlWNW6VE64DGZJ0Kn2EeFq7he97eqWDV0sJC6kqGkrFwt
TF4kmkJiqqLkBMGUjpzDV4FanVO57ppEGrTooy1Sq/4Cvd0qM2eHDRMYZJzHl1sJ
KMcv1CmjBZSVdhzCuqzf0yFA8AmW4DOjhNI5jCxoxPKhMtpF6M2ZQip53mbPdvmb
LUXE2pwgc2DS7dSkN6yBa2pJNMmlW3tqEi4xhiAbQvUPX9I3/rF3scXJg/o7C+kc
FA4unCvLWjxIk/G8CwxPEgiCG62JR2LTvrhEVRolb69dteCVFgY8FoC2jn5mT8U3
sVo+QV23AHcMvltP623WAXGqZpE0Nh0eZ68Bjzeeq3RhdGs234379J4dcVsNhsC9
sWm2y+B915urd5syUOAyR2waRHrK9+5MnPAl9vHzzlNavKOrA79TwedPZ0AUDi30
owvkuihO+F+vpM8rEnRovMaHVIg3UY3CUAqxd8sJcdURHsFjWdF284vxLfIj4+A5
le8HhTuUFahCn1gfnKg/sp987rKAeQj8xepTA66uGleD3edScukiK49jl9OkonBl
PZJujzb/BtqlxpdDEnPZFme5zZsFTDtqhbamkkaUriEfuy04t7zihDjKNJqsibjC
s7OrSVXKFd2DjvhCZ9zj/TFZzYBjEJKEkpAreBMA7wmLtLcKd3OlR61y5oBWums4
M7hseZiJAUNv914PR4kOBF5MbkIsOaMcuyR7VMl2Gdn8Im8difJ1U+bnyeIxvClJ
bNMBWZmh7ExeB6NVfWJ9bW0c8DHMWSHCrBxy6kwzIH+PbhbQKJO3BpRKk1FjaYbl
yhyuQKW53jlpvfEcTzCUvjmjgxpRbORPUIR3PqCMg3gkG1OpnHEZOz8qJbHEg7hC
iBy1MJGPBaSspnPBwLihTEly8JpfxDjRjb/rGz+1OPh6xgys87KQ2hSCGd2Iq1dF
p9pRLWaW/pecWps8bjjgxBcE1/7WddGN/ZNO7SiM8bKrrG14BLLZayP3IuUe701n
63i+EKH2YgIEUYZTh0gnXte4zxgM3qzdZKl6JVhTOH8bJ3ljyRGwLOrhh2JhSIyF
uKSRUFXa4tlGcYHypPNzZaZAqcDh7NnjD7zXk57ZA7o4EfPigjPXDSEXToz3FNye
8ycxwtbKQF3o6Wbc2WfbBjDfe+N7RH/NuLmXmGxI+N+hTqIg/Dj3buT/PDstIhAe
MMuwQbAgnUzOcQEBVQbDOTUPC76pkZeNcogvkzJz5Y+vR/oMuf9IwyCZA1xXIayk
Ot1d/9mdmXg/CUpXzS2hG58MUmWtEc6lPAkmnkk3elhYk26CHKa6mlb9vsTiLTq1
LoO8ei3jHZmzio2Vx2j+W1hBNndalDKuPmT32SSz9Abe6Huhn3S7zGukLs4Bb/aI
kHwV4QPLjSpBAjks/ecjvASeYBoI1ZiN6nPK7OO6916AoF9RdVprcI8CAumVIiQx
hpbwAUXYKvKaLoysbYZ5g3qfOPKocX2UMRHg39cD9gYR1Jh9VuFjHV6IFqaoppYE
qcGN967Zh8CACZjjC8830i50EpNLD5uPGFV+TSZD5ScBTo1zv65Va8uEhMLRxVcp
JNTmz+hQ4JpOWkB++8Pl0Z6kPmpRWaCQ9AZgQ6ZLFth8kGSkcMtdYIgKxkI/9PkW
aCBexgRF+OsygIZbct+xc0E0VitEDXUGqvgtFufYr6I6QQDFYmZPVFVb0fLlBc7b
bBs2ofMWn1MSxd/90djp30P6vK8CAgU8TVEJI6i7KWiq34f9Y5UWcTOYgn3XJfqI
2fDaeMNIP7m4TC+Sq3NEUA28CSWD9QgemNHxZFBtfLGBGVy0OK3bDcfygjVJ9hpW
PTUx0tgpjnpzLAU7+EgcDQDS4ugTod1obI8Ff+Ofud+cFLJLUWTdq8xM8hbjS5kh
3WqWdpMfUCItvo32GGaQipQnXqhxqtNQY+EbhFN9YHezJtCklF1Ni8IRC39EoYlP
2gOdj4vaawiW+P8ysgFCzLA029mEDZXbhuwS52ao7M0KobJlkQyjQi3ywWjDEKoH
J3t7OEIeBvMhhdGO/tbbSHEWsoCBJRvo4JWGp0PJTTkMkY6jQdRr70x98lJ7yWzh
q9aTeJsWp13ZyfVHGvtYqgmN10CaDPJc1lv87si9NUpuJ/Gdaeq3h7sRckwJAJth
/FzU1nG8e75Nn7VUIOzB64q9gjTN1e19g9LXGNNKetdsxLYR1sk9+IoA9WNRWMLO
2b2ugCBhYWqI/XWv0mLcq5gBoEwiF1zBx5IcqJlq+YdMt9RQAGAG/vR+3OKkzcOh
vb4MBl6zYsSy8/l175muDfy2MkNhoNIVTSfB2avZSfSGfjP8H0G6iI1y4pgwbZS7
jA21nXgbW+Ltg2yyOdJwpUBaW5JgzW4wPKFi0fJko16cGWuloAz7qQp4s15bHoTm
m7nHQuYQnY8hvfdCkCEHZ9w3hZIoxBIyd1aK+oRdGPfbaC5sAmjAZ+TcmaLdkm9X
JOVGG/46NqjsD2yq7BluzcUxY0qpESbLCrSDUyCSO1+lilaxRbhvSxlpyBzWX31D
mTmKT03noloYLhr7AJK/qbUGawkkCKJjQcwTsb903fim9QdHW6oCgrEyPSS4JbaB
15P+VvOi84MU0lcKToQ7FStrxqXJKTr2MfVPydyn0bM5DyGAG0SRv1RCf8rXoufe
pV2P+sVbMdtRnOtdqnmjPs2TlWfGeS2bJ3+xCnGUnokmDgkko3gM3yYYA7EEl6Cb
P/Rm09pMahmKq1THzVeF1WPu6UaaUL6HcwgW5/tgUAYlTuga9jvnkBdqO3UcoQtA
fLHKVkDXo67hhsWDolqLD0R1a6douBjrLjFL2hoVT7ddZX85lGnlqFXLMX7CqvuD
MMKKldrAiO0s0EB7iMLC0XPAdBIp2z/7mbQTIkDvw2JhZqL9WoL8fmjS/eMJiDYL
8v0gTRmxQVrBT9elNBphJaYoQ2I3glE/F1Wy8o9YiCdv9SswPjm7D+/6SqNcSlXm
1OQp0VJl+ZUOgZEH0n3WzC/7dQBldJkWRFcAGxnr0YPiKepuPCYDf2YVKqy1XtJK
TyQCRI5eshdenqScEm4oJjplrFPhAf0h40+dFyQ1b6ulXuZxqU3SPPSycS3srWUS
PAQQenGlnQVLFi4D81TWhcTX6srXFhieOIlQUvfSb5e6Q5YtasULUkfIQyx+6Mo+
nld7FIk/1yyPFimP+yrMiF1NTE1rbtRhUxlup/UzHb75ohC+4QF0T3PVkKbi1Rbo
14VwlC2s1B+kvSx6a/7MvFu9QKMXXhKOR4pIgR+9BZ3MgIIvKphfle1ejrIRQp13
qqvo714vNKFocfAft49Nf1LOvDAFhUvm6K4pjl8xOsPChJpccYFHBQLVtiqoNmu1
q2vP/th3GQEtci0dCQBe7YQ4WXFlIsaLP2aeitggFQAWR8bPV1OUJcknIk3foI1k
U5DIHbd1tavoHWcpKpjRapvgOIsBT6JDYGk0HC4XKVyaQulRMyOJ1pqU6w+/Ko7+
jhxHFjItp9yuQ98IsTfNmS1dT+7dgsfBkVYiUf4SNF27AEmv+YqU8sH7hQkR9e6Q
/oKj7txPMHs7E5e2gN6ZLtHqNvoG0YMa/y8IJOtC++hQ1Z6BejzvxRVXFU8EHcnW
5WeVK2MJMUWbYSIGtwKVDc0N86UqhWIg06V6zJjZfCtTj4k9LkglV54A2QdoodHc
gqKO035q1UHGewQX/6DaujfoiP5bCEMOdoaltgmWrDqBcg3UFgJr09SUZLP9Le7U
rON1OUzwi9QMNamXbmpq9VnvnHOWqY1m+NZho9GhCgFzlIpJdPIijFZSIU5UmJtV
Z7CBDv2jgukLNk1RBa6vj92W6PdjH8/EVKxK2HEqymO8OoyjOOvId0zEKOG+6VPV
zcXaKTtrp0ChLBt8bK68c6w9PXmc1Z/hdKFu1kPi8joDgU2bzhS2vwXUZQWK45M1
UeD8bAh2QEYyxCs8LGfcL7S0k+WiYmTq83oYFDTCfb8OEWlqLCNRDt+7fR+zIOZz
UYmGpP2RNClzjjiAWbRbJtoqHbw/QH/wq96UC16/uC5/qafuM1warh4Zfz71D1cP
P+XTZiO2TY76F8q5lN9wsSBvcXS8U7SmcOk2GYh4bGZozfyPEt/DZprpuWv/8nbs
7G/15IPF+mXdmZ/0hSWSsZUjmipc83lBPZrVk+yP5p527XIb6SL1KJK6YQfhE6Rv
p7baVJnxU+TAq46l4tLWVfVL1zEbNTi7jU24CUvLfT/+BqgIeBMU8eGEBbpNsjtl
zpMaXIwpw0Uwwy5qCvN6bq1jRghzPfeTIrIyyCwQ1Wmg4WLLCn5PC6NiUClSY6XU
8ig8OoghOD/ZoCFyB/Tj1yzridhGRhIJGeXeKUW15LVdtE4mkUnPuMfpfGPufMKG
kZVF+FPyi9R/kqcACE7HhpcM5rUoTJm1+jK19iljHIKuGJ5pmCTNlDFhMO7E22Q4
e33r9cRsOmhpaYj+hS0IGItjnxsb7jEsLvp5QGE7RL7pjWBJ3TIyzoNqYkyLOg6g
3oH8nRo1X/Iuqfhxwb58DCwp71U7p/y53DNfRi9KHTrcGX7OW6P/CrSW3IQxuybA
BdQQMLpKqPXMI3/wG2izsca7MMBwDOzD5lBbM78AptWkm8cLpNcHxONAOPeQl5Jt
uWDDVpn3/VgEQiTw7n+9WD+D8eyDF6NEVO3RXwO55cUOi1sip0bFWrzBEBIhs7EN
lAIaHUGI7to1WdSMdZR05FHkcmzuBwOn3okFGkMVmSSaWJ0AaSzrzAo2B4f//aQ8
7HJBVFCMdmRevuFwcoeDgR1BY/Ll3Twzu6GsM3qAe63oywyV8t9xcnwqFl2gevCd
ej1dMdBHDdFup2L+U6z1tVBlVO34LmnaWXwJ6n6FnTgRCNWd+AmEmZFgqjPniHXf
ZsBiljkT89jnYBj2e/MN/sa2s1M++mSL94+H5QbsoPA3Wpt5/Yi3tJf2ibrAa0IS
LBRkXThRKyIqK5xgrHZT4IvN/VRfGHoapSLhzRg2/MUgjvJudKLtK5rl4BewzG9V
0CyRahxl1RPoJwPwoCcQGLrmfUGHsWXxdZOhySdMHR3mCaPmdBSWHsszCYP6mYZH
BvUnvbhUXU7xVUMTj0DmnWLSEVK0qkd/vJF5TRW+wumL4qlT702e0tx9yWo2i/jc
ZVkukE1flwXLjSsvJD73ctIE2py387cbkocFT8ywyg++NSG17dsB2NpTBp4Wh/QO
ThXPkll2LzDER6rtWxEzOR9VQCCsPgtVY70YOywybytyiDL4zu5ay+Lzpyx26QKL
d8cI/28kkh4BxAMCqGCvnSI6zlS36JyA3ztBpxr25nJZk3hujbDRvceWpZvaj6qE
jmxAFvrvMuYuX6Hi0z/r8HmWmLPxTXPkopSg0m6ZLY6o956NLWFrfg9cNsuksr1t
rgxwytTdakPO3JQ94dwwjHb42F5KunrfjQlna+WpuV/HHaE9JX+KDktRAdBQyiQ1
1+e8YOqSN5Cp2JIbCD8E+j2egUa2ULiyL+8xwhQH5/szJ1Skn9SJQ9HLY+sHfFeg
Rsk/hXxIAy5uo8qfqL+QCCiTsbkddt1B7cAYp5TA0l1sPw6YTU4QkSZuRwNmLeCb
zB7GXDx6ZlOpBRU3dORQ4zXMPZDqsphJs1QmK6E4J2DkB9Y1CUaSWK4JC9AH1Nlk
ehmdAKIyjZ6qSXioBQ2deoj/a984dXl8FKP5NyAdyJ/J0W/BWhLsMyVc6rDp6km3
oRUTszVTuSyyiTXwn0GSe6l9s7fxoMtMtDgc+JORpU1t9H9pGWhuXTSN4pPC2k/Q
U+sIrFkPl4H5exw9P0Eert5G2qBkqEGsL87nvdxZ5Ur9VAwpe+wTqysDCVx8ZFvS
oSyxoNR64+r09ZAE6mxvT4pNABiQazjGJcDI8/tobnkFIwY9aYanlMtrOFFkPua8
gelMMq7y5uHMhB+UkGpJRIHwtzCoagKekohGbu82IVzFczbhodOZe3MYgiMED2aR
mPm5grR15yo45uwwHKzvY//o7sEkpOLnpTjFh6SVWu5HgFb7jHnKTIH/cU5dkP1d
PpZ2z2u8cxh00OK0jdHfVghEG13Y7EZQHJGDVCAvhKrNzDwWTSIrzHR6cjUW5BfN
laxvaZ2VNEeJo38Tp2nj2zJZLUeBfUz/Q3v2yqhqYkumLwO6iQXetUI/EHzKKVAu
SWo/vz4gUot+y5klH8k3mPni/rggOGfr5vkJhr4ieaAwRBmMtwGIdfzS2f2Gl7ny
O0nRWvTOewZRV7Lx+jRPNzzzwHScUBsT5Pq+7wsq/teFGuXPbeHwRYI1G9Zf6dPY
1kn5iJUdthNA/cfgkZymAC17QdXH+hdmlyCPRP1lAp65sYTWoPRUdAPIk5Pg16nx
RAmzMtD8Fl0tJhlS/jvnzIOt7EYdwZFuTZNqhVBzDI6WcekXilFVkM60XXbXFvs+
ojVN49OddSZu8sS8dTjq5IquWGwr4U+i3A/Ndeip0buYQiwXTUVtFNBatrRi7L/B
azkIydXmYtemi6HX3TVjBN6m9Lc6kMydYwhhRvJDC76P3Ac4t4xcFE6IEyy/Oa+a
qhydGM5LJCiCpetYKdeJLKO1gXewJNKGZHYfB7t6l8phQ6IAZ8qD5nlWltRuXQGp
Ux98ZlzgDsgMFdHx0tXnS29vRuyumZau2XN8Hg3T5rZTmxzsz8iR/xridY8zkqBa
ufyXXyRaV4GBrf+1Bshj53+3W0godZBaBUMk+5UmFIB6NnYMcyPZLzX0XyBxr2bq
brvvdEt4RHaiydk4abpJQ1eaOC2bnSWuwnBCYep2a+fwYTuq/YnEnZMZ38ehmyC0
nvIw4g+Lsdj1ttFaEgbuxj9eb4iz56PjpFtn/4560B18M4i3SPjLxySpyEkFFN2W
pzeQC3/1ZOP5NeMImWJ4PDD71SMkvcJdRcxUX21/cL3PrJOlvXIu3h0xaVR4jc6J
hz2oCsirkVGNiBxJIjxycZxB8ZWUWu2mRiwS8YUwZtDAmi1tWNUynSUv9cFrL+6U
8mgSGnWmDIDHtqO2Sk4kMfS45p4wxhA8Rb97UzheIFmqA/11z/pyi9z89wlqo8/t
Hqj9wy39dNVfKAtfUZApQp6OWDj+a5d/2ZehLzW7fC372QrxajQLNiZEskPr5pu0
s/6bg9a2gNgsu4VRSETUeJfHoYe5BPQZrjOVFzNhgiNYZmfwTCp1g3zfntyV6GoT
l9rpDqqpHVIS543TCnY61/wk77TK80M0oDMaGZpdlkuaJiC3nTVGV2g/qxFA4VXi
Zl6ilCO0qMeQg6R3ONRnORRBQOga7QXH1G2BEIfKtOGhYD9IBIcedC1twAaQymkG
3WY1bqq1w88HfD1FoNiFFFxlfWOZViU29tnwF//t2EbYW/OSseT+r1gFdG1AWcNX
oZXeeKbCXnJT72GBhRNmCUaFwWZDdcOXUYUSKjCBoltdiMxHVqbZp8deeUc7KcFT
e5b3ltjCN45jHBM86bpbULxAeju2C9uCHlN6jOVuqzfflhVTXukDt8UcjcPbS5PM
1p0nOx6YDznn4BdoHdFYIFN+6IBUhuy5RfOJLNGJDLtyxOqROLwOpOX6Cz+q8DL9
L7z7eT0nQ+phjMvXy5/0W2J77a6E2nn3VBAWacSRLOi+ojlDCGpUomrqGW+gKmdm
gqyvmGeRyPjmgiY1ngIHwY7YCbQSZOfiAit5gFuPR9Lim4HzBJZnJGk3APrzzKhM
D84VpBEVkWW2pkjRn8wzYbPfDjFQRQdrekM89TUW0Z3Nu1dQnftt8iog1p0pV5Ch
9ZlhaWA7NWQYCYKQZNip0gDlTF2QsbUtEtJk0gReHrxqmyzE5emBM3wRLfHbFCbS
ulyJ/pVEUAJGB5ASPobs9JeRL4V7NudV+hEOY/ZMTG+eCEo3Uyzax7pbDVKHlAU3
rPP+9/ap26aQmPNH4DgTs4XW7kjthnE0V92zePNKwHHIFivwyV2u06lqfnIEvDxg
K7ZJ4fUitsQN9C1ND4fUsZKPm1mrTFPymF0DPi+iB4J9IBNJTiZcyGe+oMuEBMUw
qF+IskJ9VLR9EzuAYK+poP5csFo+8T8jm07zUxlZt9Ro2L0Nq0GnnUtyzH3zPZA1
KgBHRzf8pYQfl7krJk/26FBzMb4ear/mpD3acxKYAvYJqsK1WlkfJiqR66GA5ASI
C6DZk/4hdnpmsKQyF8pwNIZODi5uKdM+rMhrzui+58fwewr4TCBl64n+lQjkW/AU
JXGkJbBJeGdP3jjJVcpxp24JZlDQspk9JHgum0Nt+lgmQEERhAoKrWEF7hv2f9g/
gtUyJecZPtAZNeu6Ozb3yBOfPoWVLUW0rQzIMJIa2FsMMTfBt0++ymFlqBq5FA7s
lGa6ZbogoVB7WSspuqakyMRZRe+AuUkRzMXeOBOSn9qWVLiYRu+jA50DnCR0hVJ/
y4YTCn7R1A4EP0RmXELjoRdazH7sXm0I7PlSqySD0RsvakaS18+0rIENMkehqg9E
2/1YUXqarE8cOD4xHDmQ0k0AUQj30YkL5M1pj48/aZWeQvEA3H6/tfS42wPYi/8O
3MP2aUTx5E2jbiIb2joY84J55booNI6/EMzhUnAxuwjf48zWk8R0GAOw6zmuPH5V
usIq+vT+UGyyOI4DEyu75f1fmpHaGzLqaUZF/3j/onUEsjGXR0mRG5z4MYLGmAPn
H/z5W2D3vLIFpm1pJzB1pl/tW2OwAAowjr3ZO0SEniOV4q5qKGnQB95Dy5uJVQy+
yiNbncXs2gt+J1pP7PPwk1D84yJ7yTPy2jiMyihVyPfheEdqQY0C0l92Rw0y8qxQ
0wTiKFeViDtXr/E0DzaqdXcEtt/beY4p1J/La1uIjjG8s5WWVCKOrG4xgBiuxQy8
JcSjKzTzyrZRT7+89E1wxOxDouasbeNJBJbfxJ0okPmOciG06pzTwUAynBF9qAni
CzH4/dvyRfBA6N5TwHajX7iCMq4xLPbteHCTmzqn1cEWlF93x7/qB/iROv5El5oj
fl39Bye22BThJ5DjvGoRDW7IYcYNIiJysoou3xB7biAt4KKmuBJ75NUxbSLajeiB
TXIwe12CbQtMMwA838cMTtsqlB7tf1nadgYwLtu7cQiJV9EnjqF9UH5iHVZucezX
NJB0Hjebcb4I3jPDH9cArkPTEMdRYUeTyfl7XkS2MX0LyzndUBalGrG0I+o3Hhos
T1vPSKdBnqXYtCVeYfwG/fN/xjrtuvA0vE9+2ki+SxJLzAu87nL/5nKXrTzeAsGg
IlgRbzAbl7Y6Q/sTIeol1hmdWXCS7Q+ZByzSmCZrHPoJsJ40n7jUgFH8KqJLnc5D
cbO/K9sp/xXk8OphPq1bMAT4u4VJ4WBuwUGLpcCCpRo9h4uXnD/IgKmRcy9gRUgH
5K5AnwfpqQ3Qk3u9BzTdNqpx120yP0YIKtuJ89Y2ISBgh/1CBJIXx93MshIPaUs/
8Mb7rzQlmPPcLNcqvk25CHjZAMun/3C/QiDAAMNy8bvY8iFcz6y33xdLuXoJycxt
3vDrdROEMGQKs8kq3wYvwt247saoRSyiBdCjaD8RLqpJa5TIthqzquVwRWmb74OK
QQhP2KSSP+KwP80mAI7c11KKjLU28g1uDWFqiZiICArs2v+jU5gLOo/gYqaC5EMu
PgVKJbAydkQu+hlKIigZ/HD4fyf1wI76y+ugL2y6aXjGHuLI7lQqPE6bndSFBrgh
IWqFktvDYiQmB1dVyv1g+WQfXn6d+c4npKTmx3drWfjqp5v6L/JVTE+S8nFOBUpx
rrOzjATKfLkuS+j65XacCsyngAJ9Ugy+7Z8nbv6pBAtMTzHnDlWZhhnmkXQep1LK
bK9/zm6yzONgC92DmxdGhGVNwlVpoROLFyZEoDPSucFNEIFX+vaxM02EW3cYuQNj
wDZjx42bEJR+Yo2f9hLnYvBfFjP2xJ9PgfNno1CoSVDve/AWr0rwBZdqKqp+5YSc
FQlMmwND1tos47BWMCIzkt+6wo11W4GSK62Z6x5i/nDjdalDX9DzUDhSshOGaXw6
mPavX3ctaPunGu7248FaKik6WZUYQiWSWtIJt86edKahwsPieWqoMyLT3TzsoBfC
gJG+GQsyUHECPYUoG9r183Orpt1sJo6BxBFxomWi+Y82jbNn5+IAyuLXSTq4Y4h9
EZwLcrrL089nAy0FRoqrZFkvCGDgrzJpF9UjtZYPiz2kL2RJnOcAvi/tqCYRUVHq
F9l3pPA+RRUGm4SKlL6KFCdRr+SDkQOawhs9V6dfPn4Rvr2ia3J7MjedM2d5Fb7Q
UiIIJr3kGu8z31pbvaYI6QA+b45jfzhXOwpkNebmkVqPg992metWDTYrj4aGqjDB
xt8U8TJqT7aRlIIM6P0lNzyoaGdVA/CI70fP3Ivl9aT4LU81JFK28NaJztMYmGgj
y0/NStZzFveGT9XktuBnWqG6t5yR0kKLm2KLmiCoC4FaOd8JzyiXmjOpAJx3bFoH
yKt57E6UQy88a1Cb9OHma5o3qMZXRZyfyV+f6AA7Jr0puCBskcEBDejjBkCkyOHi
X91xJaHAyO/a2ckwfIfBAQp+ealxVVPBMmKM+LljVp8DhTLzJW9s4vEB7q+ql6HS
mcwGGDxmzScyX8WRlOiQCQfBYpsurIAekeVp5yVOpq5G+F6l7crB+J8p/xUMJ5hU
can1fWy5sCmTEEry8x34OxOgTB0tzsOCM1AYVZa8b3R7dFrXVYc+8JMT+DpkUcQ7
pLJpDQU6LIUuPUy8OxU7F0ckVcfkoiMG02E96Yy72X9zARsSnqJKAYT5wF4hzDBL
Mat5pvZPeKCAWp2KB1jhuSbD6gAhkMhJ/PeSQNjKbrCVLm9WpoUYNDjl2zJYDC1X
gLK9xQyikPkSW4tXjzLrA6F0CvGo3X9og4BMUzCmc6agciu27Qn0h4wyK+0LYKc9
sXIzzoi3aROuj00bBDXh2MlnCP1mGP2J84FBsfo8Ugolw+qbHUoaYWDMreXpHzzt
F04GN8EBh+Pu0trg1o5yEE/6xhtDn7RFmMyJJYVwj8DbcbIIDdjQMbqAs2PsC85R
HzDt9vDzas5ukncg7IW5Llss9ZObpLfWu9MBkyCOFCwPuTjZXzhibVudkL7PLXSI
cY5FigdfNSfGtDB68Kq4Bt2j3kb6u7Iwk76I5ukR0+U24Sm8A/Ylsn3+dVx67ZR4
KcK+ojhaRNdJoB1ikSLVAhCIsoZLlldlIYX3UksxgvB4v+IB7DNm7Pd4nrf0OfGq
nJFXeervelW4juJxB9cjR2AhGl0OslpfmE35nQ3B/dOOGZhFPqG7Rmd2lThODuXa
yj1YiEBRGw3IhADHdcJfprToYiXfVCdfC/77YdyEYlt409Y//rG/GLniktH38El6
teojn2MsJV67MAc3fDWm58pxdC5QPsTlfn2hSbViqY4B4c43+BbpyfTsluTwgLdL
Y8uDaw6uN2Zc/Skp+mxsSEVfcpCTv36RiLgX0AJWXszB8TYQmvU756+f+08lhJUB
7FaN/Jl9En7huz7ihT54aq+0dtGqmytF4BSoqiAofqfF17j1OZfGj0xL7QNDObsY
FDUv+EgCbtK9iAbLJkyDV8OaYeI4TZdN5Bd/QArQBySBR3Z2kJlkqcDHr7ByaC/c
njYxbZKTWCg8oVoJtLIBrYBhQ+BIjWA6hnegWTrARtsL8OZ6+Os1AMi/wVkoMC1i
jIp2Ss8Kghu6Km44j83uSFZjqJWv4CgocepiPYMX4yopGkAxy+iENeVXfQDyIpHN
XV+d7JhV84Ck8svAet9fgjU85preJ9KOPkD1WEhu5LHuDhStcJ58Me2Gtu41EwZL
XJ8AlHxY6d4xGDeewfwJJDTVmEVdBYXr4dvw3cWFA7aSGE5RjL7mOhkupRm2H9MH
yREX/WQVpRvEKIB7uUXoHN/JqT5J3b8m83EZQ5tXjZQXpAmbY7coxfTRtVNAIwnv
wqGYXUnMR1EJksrWPfFIPycAWHxIfG7y66mFoL7VbRPLy3aOthi1xvvaDvnxqraF
fW/zbub6mVMXD41WEQqklyAswbwjHztwsZICm0QAW3/u5+KnbalNivI0ETJ29qRh
XNCZgayYwh8ICnXVuR3dXRHy0RuG8ZaAji8dDqsK6UFPTodx6yjHg/3wTix7QVyp
QmA7RnXqwVFQ6MJfoQueRodg1TnWvAKhbEgILrfHsP4WZ8Dh/zuaJ3wdzsOCOl9w
dxSq3TEaLXKTNc2XXTsmDFu4VpWsmhTItuGy5A8HevUUEMDseCmVLYstBq69kcJo
1EhLtV/mv8oOl3koqQvRidWqL1oieTGo+w4tmjgVNVrAgFg55c4NA9Bqo8ZpUvZn
375P6kzNi8TwJnK7PinngBxlddGFmsmOoI0pSEzQR3lxIiG5pqfNghNN0MjFCYBR
IOVIUgWHebtvZ0PCLKckwZOoV7JdPrsJkWu47MUZOU/ei8xqL+EXkGWX0fmxgNKo
EilLKNVxEeWB5ghKFvfpaUJm5hRSStoaxeySeaCwYqdI93BINd9Ovz+uwLKl/WkF
6uxj3UR2+nHhwZuo5XyZDRl+LnVL7+Z5RqOt4bPV06I/J921GzO6/6KlERvGWzBJ
+MeHnr4cTpiUNAa9hXa0Hb8CbpPaBlqjxmJRYcR1joi4/YsJMCNb+LMYSVlwgKnE
KaZ5RWkoRa2EwPeq1RaEKfvk/pUyjK0ZAMab8rRXdBgg8XTwiJ5DjtDaC6wWloAK
eTZ8dsQhDDrLKkZ1CMQhgkTY+AnJ28tj0BMNariGqcbfNBWE5Ger7XNqax/fFFRZ
HCoMOAnpPngXtkAGHNn30ai2sbvwaGdfk5AwSSqRGwW3LvwSDUnbGaW+JKP7Nhhd
DXqN2eJgijIAfWsGd8real9lw78V0dBCI2xC2zSr/vxV+mGmVbFo1nt2ZBkEWnXO
59u/JGB31wdiV4GRv46atCT3MFxrMWfnrHBA3NrIVLiFL6qLSIVhVUAYe1pB5Hds
M+L6gR9gIuWkM5PFkGNlS9uuYwqNazu1qDXYaLWG4ocXjpdAWqMEdiit9G0oLNy8
JZ5L65tRGD9gW5akWy2o7uc2WTekxhlWV5AhUgy/hXl3ADgSC+7mfbhzMTjfnZnm
RyZWZeBVuwecoGmoi7vFRdLCy8YUGWqPGPhGArmRLQoes9ctaUPlSjBSiuewaQ8m
vLxJxJywmq8+8c3HO+dPHVNlhV8glZOWRKoJQyIy8ghdHU8XJlYL5Kv7Al4jcN7r
6yS/bnAhLMXM+X0RfWMAaC9Sh04XlyDWLLe/E7uDFW2KRIMQAGxLosm5TRFaSLOh
Zd9cukbz6YvX5eIITqCDeBOnv9c0oCkx+fsLnaXwMDizgzMZvVa9GoxQJRWKirzn
ZQbYAgWyDyqAXjKI+KPbrLVOBwV8lphildFDnHDAgm4kukaDRmYS+O8Mc2cc+XdD
wUPNeNHy3LxJ+jL6K6hpVn9s8xoBHP6NmMEf4NJd9OuXDKJRzpEPDPu3ksCyOJK9
x96dCpke18hdSjPcKxd6XRgpxmrfohMwdqbM2PPiZqEHkXGb6gF2sSMD8keaRET3
SbnhzQcmVi+dwCPjKFEjO38hILqfq/LDRhyuDMMJIAl/0avKOXh1qpfGf8xHJzt2
WkcGqx2mFDFGo+ZN5siIoY8WcupqGdWrf5AAcj3LkqGqxNxSMofbfgBvlrWeyiIH
N/OGwAFBWlh+0/qEAb+Y4ANj7VpRxBTG61qV6OkxumP7M42gsrXkMXGn5dsyU3WV
ZakDIHNcURLqYjISLaigpgeNZnxCZObuuo302iuK5OnvOY96hFgonjfqYMcq93C6
1Su3tzxo6M4Lh2XmbPYncnMKits61Y6IgZ3BwGZuYOYzoPocNBTvMHEpCaGpE5D3
GhzFHP8+eeDivhGJ/B8M+0QcWKd1IjCjivz0OcLKSbx4xmkxyxuZWgZD5oMB583u
FpzAR6P0Fvm8zEdoah/9eztqpjdrcIHX5Q/k+tY8SXDeWhzB9WA1GHROU82KTPmh
jgaeRrw/DjpwRvgqzur7JSvjxFH69qANd8RZy42Uhif8MpxHH3Td4xXWiiBbCTb5
pjhTsgoGpALda9oVYm7wGqV1t37yPe+RE8TT5XzuENbuDGQThrMnA+D3Lmok5/JK
gBXtRyQZpaH0L00JOHEzuMDeLh1r80v2ruc8R90iNG487oXjOPbUjFQPZa6O9+Kx
KiOuGSnvW19aCtBf4X809yMCgYmPCgoRwJc9w/dyVMxtb1TSlhwU397qzwpp0aVA
nbn3y1W1besDqZfZzdObjsk2HSM0uAIAoGkTBfmZFOZhfrRUp9rGoMRyzlKJIugj
YzraEvG5MuGboNpW6F+FmXATolusWepWefWnkFv/u51byiRpcMVI/QFwuJViDboT
E5Bjbt2NavE6Z2uT1uf1SENj8+YEnafOnyA3MwrGeJkd8dAyYw0JffgOFpcVsklM
ZN3gpcVA0Lc38nULo4CSQe1ZMv74Xe2OMOXYFTV4kLYF4FdFztde1AzpeWcElh1J
mbF6RaW8Km+mtALRbCMpGIboD8QryjJ2cisIveCKFauN01+XFSfUbnX9mlIOW836
UWKo3/SWny2qbGH66+kUQy+I/rCRM8rxZwIyYz7TE0c83PzqXvryifNMkn1d6dV+
G/4a8GcuOltuj5sIGTnDBG/bWq5YcVn9kPjgYl68q27reOyChuX8Cg9fwovOewjt
E/1V+AP10uTC2PoDwaU0/8Ud37n19NQ0VTBoyZiDEd7rYVnN8qj76nJ6Jn7A8Zsd
YqFdW2+9ZGhEWd/jsrO3D0bgzKl1hH63sJgzRCpZKPzsP5IA4vB29ZJWbtm3vrDm
Wf02DI24NoyEgg8lbJA4s59ixoj3XpRaA2O46DlkmCuObawVZ8Uf/E6cyQzaQX2l
ayJvU0m1MqAyVS0ooZP1eVTlt0pqWGp4sKK9+pG7CFDDVyZWnoIJXScbAelCZa99
bKrhYCZqrC/4VmS0aOVREPsPxAc/wB7Hjo61Mi35V1Sb6qQPib02NhO8t88el5T6
J+jnA9wYk/pLQg6IXU03sai/gPZoFq9delMG3YA4OoyHMfOBXK8+98LW3lI8JcH5
bwiesslPaNCh9ukkzSdE6t/HKyNwgLCNvBTHFaI1nNkbVUs6rbz/WYrSQEWH9Sun
O2UYFzlrpBliR5ic4Q/6sMGMllvIBwqJ9yenhzDf0loYt+bojfHRLItOYHUqWJqg
/RWrdhEHq1vQ65rWsisTzEFPPReNj/Y0Wy7E4WtTtG56IMhKhkJDa4weEF1cVWzp
kaXWIlW4wF6zj2wOF6butsgHV8rfu8uBptMLupDlyu5okD+gbSvFZmSxHuGvLbvg
F36PqI/XBPK3yqmHcVK4JC8K45oqwY672km2cBGwx7Dn0p3PbTKcNOn5sqGjqNHY
5Iu4/OJcuAAd3uxfOm/az0Eg5CC1Tr76cCDUHF/Y5GzX29+d3MvT9+ayLYAwU69A
8Y01CLNR0UPPdUhWOuLJQHFwTYM4zqyOSldbSUr8Db+VefaDxJJ2fn5b+KD5iuVW
OHS7qoe5Dmo46FU10r1lgFmCNaFaPf65b/FPLA1fhPU1yP+PpF6Ao3J0QNkMoaYh
uHI9YsoetmHQiPEMYCigQsbXcSPdSSjE8QoWxgHDR4H2MJPeWAJrCbeSZvCAOcmV
5/LCch7jPhRpMkgaoeh7JOg+ySu5s15qRapVnZvj9hHJtnQKTVhFReClJychywOm
WTxUd/a0xwgI3RubvgQkD3XgCvz3lDElEfiQEVtPlI/i6ipJOs9jwVdUzUylDZ6U
42FeAGBDDywMlUGbS1KgGBcF51HMQs47dV7SNlOiUp/r/IuAXy+Pv6dYCJKMoM2u
Xq0SpixbRBJUIStZxXCOyqQ9ZjqyJfcLNeMv6IVGnP24C00t4BpuiG68pWc0v7jV
h7NpcJwgOK6HTManAteXQdakLcN7jZM6f/SK6yNDO2annAhv1IhhyXfa8xomniAX
VOHx4MTtvwLPp8z7rZ3iRaLL8gtBUmtAfaxxSmEuO1WgN7FD1u4uVbf8GWtkfvGW
vFUNbzewhpQE+gMhGMqzumB6FxRYpPvc8lFG/uKQ1OlhLQ11TELv5MRc4id0s5Ey
ERNORI37HM7Sc2J3dDK8HPPEd03IBOOFYgGDMRrcvVmT3fRLg6l4bsCHhK7wL0oN
PlGimyik7+N+k0zQ6VAp3h1wRiYv41Nclz821p0yOt1iLYd9nMBIk/sLO2styZie
hJe/bprULWIbKmzvxis4LzV7QJW3Gtwp6JJVkDWDjyHv/xprYI4K29kw5iu0qco6
GQBGU/frJ75jHhJJxBDa7RmXiJHPVlrpbj+mkKBvJBumpcpZafSqS5SdPouZZVKc
ldsFCCzO7KPymlwKkWEaq0MGKAm9hKoGUdLIjIBMn63lLtfuY0GDeFcigtklkZq4
Zb0JcFq7yn7niVFxqJUlljYc+EouxuYlbeI6BG0Xld/tsocbf2x8NB/p/rRq5NzJ
uQeuNCDLLnT63AOvfQ5j9DFxCvBz8ZdY0pXKQPqginhi+eLI0pqWgRwdbuH9yyWu
wvr5G+wm/QFNvfg6Vf3Iv8/W4mNCjrN/JvIT7R054yU9/aEq+koMLssdxwtzGnvd
hjnyp3p+04htT3fhADOWd6xR0wY6DHolQGdep454FZ9mk1bg92Murff6VdW1qml1
5WtYFgQwfYbp8GSkbFQ91Z/a9VV408PtlmNMldH/BFo+3dxAHPkaJ2crjg/NsrDJ
O3vVkZMfnQe9PpzoeqXsuNGpYYPGpH9aibuBH34IxMOv5NcCp+tyK2Is8g5CY3kS
LgrNsy5Fm2U4LCvhgY0c8eqtwFAhzpvFjsqweI5PS0GtqP0cBNXht3K7Ry5EM6Nu
LKPcoPCqE9WCMaBKAGjEk/OfHrCI8o4LweVrSzbAz4xWMXIjdY9nkWD2ROLqbMdS
P/TX3iVxdA3TOZNyJuTm5Cta3qRw1yumui1jNeDDXzeDUhl39aDhGUVKVh22nEhQ
iQgz89XkLHTPZPU4GwSkHtylSRVZNKenq38Qus65cKN+5IXcvTSsNznKrO+J8y8c
r0n4H8cSKoC7GQSg0vaRonrJSMXOBkvFB3tlJhWXXTHIwXCLAd5s07S8xc3mjd+M
1mDeQhGZpPdj6Sr0JQ8LHMzzHYm27rvtdPS0d9i4vHY9tfkDEyoc+IBcOk8KBkYW
s+x0JLSFwuWqhSmhIqAsTTjoJnlKtJfecvXiYcQHdsRB4q3JkBAFsvH1tIBtdfGh
wgDYxloA32JojdiIYYyL9B0Bgyaa677kwjjW0gFWUxh4kbnoJZVbgQbblBJteKW0
klBxHws4c4neDHQHIxdM0/C/1KgTDo90sZz26WXYfn60lucds5DPK93cQg3JDtXP
yL6w7G4HJoyxSKrv7mj2NxES5FjawRtA2WoyocELqGWvs+FSDO4cu3fUdhonxqUE
MOdxpReuW7wJqUKgcpdxlfcJhECjX8Xixa6T+TVDjTlekhw/G61Bwpi7nj3Q9CRF
MUYAsKwJIBo+sHR2r1EIiNRf+n0xMIfqGQwi3e4mF2OfPjZ7i+wpUlzf2Oagjwb8
TPTs1Ikn+59jg4pHXbH/BQHnHSXFpz7APN19mByg1BEHKRNDi1agqdf0kEpeHh7c
Kf7UvFHreKAl/Mw2EihuU/dzAcPMwVaodJj2gTl9ENpqIDpvfovkiwlOSFNb0VJT
Q9HWAPHKKbTKLCzbIyunL4CqJjHU9yWGwdHceZkPvnd6uIrf3rKniTU3haiZJ1bB
smyVUaCt/bZLAolgbgW6oAL9ghoonWNf8mhSyJZlm/HzNTXl0bzm1RoOHv4xwXim
K6msw9Mvr5ofGmduzpNly+0H6dZIKo2uUR9bpJjtJ1WHhfr3fMyO73weA+YQaTeP
1g3Kpc0Gmhav9k8LLRzi2TIF9fEjj50U3/L71eLsZiql4egzusO+iIhWHDXO4zrX
/z0Fy0dAVOzEjR1VNtcdvCp6Az03JW0Gzng7FzK29dUJ3pob7O0JRBCxEIt84tw+
BFlFlWhj1nCWSLW4ZQJyHGsdLh1fQrp+SJT1JyM0d2kJr3jVbDD3QZIUzBlp4tUz
jOL2qbWhst3v1lDkjNBQcB6Ynm6Zq6KiziyL5Rq8SddMw5xnsp1Fh1DLnuPUPuv7
hLCS4ih5dLQSGfO9GqeANju1bCfsQXQFDSjtlzolPAce/Hf53jv3GNB/6P5qAo0n
5+hfh3+r2fxvA/CRfRyGYovpitgDBmUhhYrwsi1jhGXXn75yA6i3ahCTdA5k4THr
LcwJxBO8aOC48eouKYKbJz+87oHiRhNPO6LGHuTjSs0Pckwm+kKHoOWSUrW51jDR
ynnFkWHPRP+DzCIRi+aQwjSrVPyVFq8abwv1uDJ9O5YibHZ8uFwYzgna+tIrGvix
hL0k+LIo5Fsh4MGApDjiodUlcZ03M6Rt502hpB2PswVMCML4k3aE4LzKq+WD0kZU
vfmpN18pa4mq6H7QJU38YXU0W5ebMMlsO7YznTtawnqeEJU3fbxC/6sC5HrIZ7I8
0rKo6npxcwqHptUH/EhzLoJtygz38EV9tnxu4s7RGzcVfI2fpHTURaMqC5NjvxzQ
TfqaJRJMN77VEJY9RHnppYWP4rLW5VlAg3Sk6g4Falb5U8/mFhVAOGhmOM9/jbIU
0lx+WIO9h2x8j8Fwj7j8ghQ9kZn4dUzC+g9Ud7vKhkT+lZMHN+z5mBft1/UeuVN8
H7eZ5EHONpW5HZXOO51hRJavS6E0zDR/wgCWQGjHWhea1MXkOiPIKrnwMB0wkk75
op01hPyDdTr9rpdzoewFlhApsWxykJxrPoQsG0svn4XhfnMhoyIIE7ERm92JVwJP
84sh1giB2bDIyD8HDYu1aBgLCUMULXj+f1KI655WgFJFM9KkcS11HdTRZdZn3f58
F9rS0RIvARrBYWD1g1NkmMSR/5GcN748LroUDKKBNB9lEW39xv8iR+BtvbOf/KbM
ae0Q4qFGd2fMlHjO2zR0gNhdG2eUjZjAHw7GNEz5Aubn8yAbIs1ktgYDGIaQXT91
pirTZA5sDRfnzCZXV0NmMb4JZJU6de9RYwzf0+yPWcdc5ybsrT9La2QG1Fs+oKoL
71Chg9TXqpiF6kSYs57x4cvxdRM5oJkpOiXemlNdVgbg7WeUXKx1dZHwvKanDkm/
nPK0xmwBFs22AWkJ8x177utgAP/kAvSPjP76JUJ9ydidwwRs21HwKfl4eIoFeLMa
L/CAsEDY4mB2xrEV+zZ7798uEbmGflfA6iVhStNT3BmVvqDz9CDzp+Uc4IsUrHyV
a7D8ujsH9rs3rVvnyg+GKexYJasmGH+cQBmdvmfK2OjXe3dsvnD932V0TGszzzEz
U98sz8WEwa8YkYW52hTSoe2JrL0Hbjqmko5ai2pFJ7FJf9evL3af0kJsZABQQL0G
VwBsJCbrjkanWrdeINJkmKgYDMgFHs4PSN4mQFkvyFO1zjDw/MDGXeoNJKnbTlVe
oaJmtdf7Qe2YdY/D0XqhI0jnR9FLfhTgmuGS1Q1OEI/95kBXq1goQwcjeRkYWhkQ
c7EPigwFeiOdrDUkmgDTWCuMzW0Oqkwwr20tzea4cXNtRRr6GHXTtfwmA2ZMgaiX
0LtcrUONJLys5I/mHAW4KFwQaqUaaXjjEyh23WsVq3V7SfB32DwWC9IPAvgTjvGS
5RfM4UzCFBPjzTK0mjqrKcF8Khjq8Ko/U0pgTwLM99d4waO5GKyVnXrV2YvMi5ew
j5ONXiUZD+O4AYXNa1TVbImcnUMKid/PZB/4v3fpvF5Vs0fqmk0QX2pO263Vz7Gb
1kRMy+yQcK3iSaZuuIrF3xMpEDuawuoPdO5uQkqfyVD2oau9ei8URv6mYIzN7/sp
g2T+MrEtYD9R8U7HmlbLjzVfPYFpgwfvH6KMYFFjIYv9YQdoMs3hzkCbDH/amqsH
IgyFIsNYV1Pg1E1Y9riCbfE8gVLwIjGPyQn4MD8Z5sSt4D70wsmpn+cJL1eSGth4
32BSGaXdq9uUSaecVcKjR1RXGl1COXBcW8Dfb7nKvPM/3HroE3DItKoAmfUuxVjB
gBnz+BP+x/l+WyI4ILwfYFJZBL9AdGBIOpxcsIQCksez8S3dogZ6Vh4sawrKN8Ba
k4zFjVJlo54oQee1RHt99VRBSlLHF3Lfj9Q+NlXWDI7kBNJR2T5fgC0xv/dD+Nvv
aLexfA35DXawsHsS4vp4InvBrvVx87jlC/srwH9chLz3x4jIFWz+7eTulm+IZ9nG
rcw9wrRkxB73RxSC1C+LeDBlwrbSIONIDDSPAt0DuSeD2U6a/cI8H8Zd3uA70nhJ
2HbOXFni/ZWjJJZbHMiKdq3/dlE9BtpYwENWCBaEmuKn2vFHXY2weAu/bAc3BAXG
A+tv4PmbmXgusX20QQZFYvJ2IWcdKWH1NVy4e5HTGkpxyTMIdb8g3h5ff7zZESVB
95O3FV+h9zl11TSAbZUh5tYi1ViQRG2675FHvhd0h9EjYu6Ws2rVpMi47xXfxe/2
UR0PHcgY2OEm/yB7Zp1zPkIakbresCX7fD6kV+32tB6z6936Dr52YJx3tdp+r5CF
dvqFvoiVGW41cvE1CrIDr6QD5v6rwOEnK+ANbH+IGHcHFLHIEeYZJqbQGS0i58jI
59L6lQTwCe2u/l347HA5sbQot+7VBdctES1Z5nw9LqxG5MaNgNgMTBmwv+9wra2P
qHPuTrLbntF5xFXeVnQouNAhE+GgVuRBNs5ES6ZUMt75UGjITndUH/69S0FNcMOf
BZ1ucvtcg6485iaQTi/CwTwzk7h8cAccpxJPYfmhSlTr+q9tO87K5jqdoj3Rjt1G
LJ7sEYE5h0IOT5HObbAt4FICsn+JDvFVapyo1sY5mFtQU/rkGFvaQUiY2BCVqZs3
eNWw7ctpCcAfDKxa88xg/9zk6HJ6FrCRg8HDpfAyZOFUvQ1ypEN7VfkPuL3cpoIg
IQfn2FM5i2Pgg9VWdkij05jteT2/fYNSVTSVMhuvWF067FQoHtLzaeLIvowpIU8H
T/WDGaS/TOYy9iT4nzzHsQqSEXBc2MCqCd3B3EkpKbF3vqJciksvp1L6LmwbLwop
N4pVr+RywawRD22/2En8DK2u6UMaIkvJc9a+ndhZlS2mAxrl25vLXn8q5X8mxbH9
C1uLEauPlETO7qsZCe6uuP9nTstHkCjqf/OqH5dgSivw53SLwGB+YSbzhBV7Z5s0
owEXnNkyf49PcacKEqUV2f3JCKXWcncazts5IInFkcUoLFPCmocXTYjXE0G5b92J
4xj1laF8PDaaWJDGhCtim+1czVZFLtTFBW1tgCJmi9GdxiYbhWPaVExQADWwzb3V
MixD02hsPvzFbyj1NOnkDi/a4ZYpeO8YnFsW1jliTB32bRU7E4SUL0jM2QP57aWG
Eys8KzRzhBzXqn/9bCml5KFdgBc+K63a4bu0mkecUrnetUEJUW6IrFB/9XdMjjiz
T8gIoB7g9dnlG0OJU6lQpWVdVBofFwsckhW//rJpeWr++5ampG6s9A8JMB1PQtuV
H4W35y6fK2DlV3OTXMyRn8xv1UqGgVQuFef7pZsyhLME1bJKebl8GQizltLt10c/
oRj5AACrFOyaxrzG2ntHWokf3x7TsVmR8dmoTGrJiEevZ4M6ppr47tUGYa8GHNZz
T0IVXUgIF7IjtlZGu51JTMxJX1hGG2fNvAVBwSkQnJzQAvRfb8bw9aexnUdB/2C+
qN6vENh5sXAMeY4NjmhYwprwexmAAYOzxFm5JrPLX4lZWAeBd9OBX5iISYpJF40W
q7ms86MeMhKUKGY5Wug0IJFmp9/qNwzWc2M4Z0GAJHEwk+ErAcwyLpcpKcKgXOZg
m6mE6GbyxF3DiKWRm48vT0doTDBmhQDff38Aq5DqZZd/G+KgCCOd1JdRFHfh5ByN
QMF6QMY617tyaDfv/VRemzx7fFEcP1bPcN50IRNRKj/LiMoWC36G1EvfyCBoc+XB
1JIJ2pwIc6RWXCiHzM3PV5B2p3TaPA6G7OgrWgi9ri9KeBA36U05ut7UccOABtdL
ko5hucgU4zIzhohj80fs4BmKD/7sWJSshlOGwQEAOZTSl+5GI+Kf2Y3d9MENJwId
yKYjZaYo3clSge3qDu4Y3WXpZwAXeUVDzgxaoOTulGhEcVWW01KHHEg+RTLj52VA
l8osiaWllKBCsPJamsRylurnVEEIqzYuehjlO0nk7P9sGHupgYBFen6Ee4LcQTN+
03lVxHzTvA5CfCfX4gp9ZjfFwA7vAmzCux8xWYMKSqdQx0On2wwUp6TqEmcIod0+
tH28FzH3Mp6QHl16iWGP9x89Gme4wZtP5O0JM6y00zbn5eg8vA1srxdQK53KTf8c
de+Qpge0INg3Ot74RXPngTNdZZDkHwC+wQOVefF28DYcwuVy7LcNMnOHIGPQezJP
Ol9mcmekFCaKbzMBFashrtae2M3gfyy2iuuWRnfS/4T5Wgz38rN14+4cQacONh6V
dE9RCL7qCfyvHEpaK7KruVCed2/OYLkpQcRcqr1D8hc2GZRf2t6HliGFhKP57dYR
yK9OH1PHEJtFTzPhn05v1bIYAlLP/el8uAAzNr2SjfqnYXAOGn2hbFSmsou5jzWz
5d5HVUzh8HT8LQMmVjexUns4r2fFhpejcxuz/X4HsIV96RbQi9PINRQd7Ary570P
C7q9DvVgjYBuxMkrjkqXWNw4HyA53jW8uI85oedXS3A/jdP0/K6MLdQZTuoUuRls
KHzyg+Qh9i12B5RtlK+YzpioXJXqWqqNqOyC3wnaoQqxPbuYCH288Okcb6b3+/U+
6eVeIv29wyUCSSytBcxRWHw0GA7XPGeo6/bMBET8LgrgedtvEvd+28ksXUMSqbcw
nqsW1UcfX45xubqPQxqPUqrlJ/SBbO5moCjzinfrJ7/u1V0hV4vvQlGUXvdBwhhs
h4C0lTcn25aJCctEPqR13SieytSw8xUBgDd9d8ApT6mkpzE82YFBOQLNUDRxWDy9
k891OErUqNniZ5tDyJFo6wNkEK5SWRJ0Sjij2C7z6lysz5r8cFzsrBaPviZ/Bo4S
AXZ7QJ+fSkgCxKzIyq5DWht5HPtQXDrC5wZO4/tiQJcxP2RyyM4VcN+SGvDh8Xw6
FKXKGpYbDlyPHSlSBoRKCvH3nx4UV8ZxRaylJlFHmeGZFFjSL2oYbh0x6dBxceR5
uC1xSVA3237Vov/SPlILppZanB9q5D1gZWh9ghOMI0/NtX3OiiHvrC6wgakrgFPc
TyCSdD3qQz574i0iROIIuBS524rWMED6ZMSLkaaWDoOeEITX0Jrrs0W3cZQEAM9w
js2LQ4KFPhZwAH5UxroHG+useQzay00/kgXWHNCLAow/kTlek+7jbELmX3pgZmWp
kRTS/HsSPVo1eW5wIOadv340mp3Gg4ktjrNSf9tn9GcRpeV9fyAuECTMK6muNlfj
FWkdv2avH5ZDCy3/Zncn5LwmScuFHI1F82+T2Okx4bWxl/DkfrxmvNYYiNp7ezPb
MGJy7f0s2eS9UjLFZZzvgDV81fv2Ui+0xz5W4PZ05w1DbqXcCw4AVI/OGxeH7jp2
NddcNqcEZprHguWPND7ozxWwZgLG3tW1EdANIMP7sUjWKplwdFbl4YKf0MWowPSr
SXq09Rbyv7HjRE9WpIeKpHs0USOPs6SRXw+2JbV48OM/wWRdwYtf1xXU9XfhRUfn
CnAt/Z3kAawijvyVyCbsshsODKMnfJ8cVcNBPEosrXpVmVxdLPwJpwTc5EGafuoP
nk0gfTKnXWOvm8r7kq4fPMpb87IB1m1guuH/D4SFIcoL3c8+U72lM0tRFM+kqdxz
jlSXLj+p3otQVNS5k2YItV6EgWBFlaSvO4dDl5IdfrYQ2siE588w5jSNvcJjH2Og
qdy2bQZ46G3wrQ8vPnCsJ0RZmAnlh/d4i3+QkfGAwp4IvGeQSbFUi+cGAOXXncxR
4ngSfv2MgpjqxERUZJbmLy26cQUQampWSKbTTfTldLd28kP5A7i/GgaOd3/m5RuK
qBphc2r2MN2tQgIQNVkku+ir0EjkGcVK5F77shKzmnEGUAOf9aPzLl2mF8cgPk2F
ex3KzfkZE60r9i8WtuHkmn9boYLBBmph1wKZTgzuBIZvzWDRVXgK6VAPg5nzSlMv
NCREPZzfb6OplKkDPsyjc6eGhsJB9OdsZW4+jjg+xYQ3/tytmamV9hawNgbqshMi
W4sZiJIKixHmI9IC7k9b9bYVWpdEWC5sJPKWuQ0lZEl44tNDaSbObYNTKwNUsfos
Bx5YQLC8uKN1qI5XgHgIGHcl1zunxNUI+lG3Nzxjc7tTaxjpsbSuDdzHFUa1KJer
OmVQE59ZpuwKxhXahR0UnhT+wA4Op8xIphXSqx7ZO1VY3MxSUUdvERosh+ULyqTv
1uxow8c6BTajDXPQEfvHqH2s1MmvhNXmZhU7peqPxbZp6rC6AlhDH2Z3b/QF/Ws1
ndXenDaIztSIfQHExEGbP0OAb50PPLNNaGXbyLVUWVLXFsBkevcEKRFHl8DwUGVI
M9aVEcj8Ecmpf65GnpqMjoqrvLsN7Ft/4iBLKEetKYcxmnP2ldKfx0wNxAf173sB
l/B+l39ir0DULkKaUJ6acFCqtPoLKTdmXD/acCcAvIKNvOv7PMCSr8iaVExgvS+v
6uP7ScvYCcWVuTNyhF7ktTk1xKZ15Rf89grRNPAqZ+qWl6AAdBPsltSjPyx5Swcx
vsxI+1HAQjwKrLfd+v7w61lDFygxEnHZwczjmqT99lrZlNRYbUgmYyd24KKfQkFR
JkYYSr9oNtXns8CxIXxw1qJvm3RqkcOGuli7Yb6+x694AU4IurBXBpIeUVpS92th
ZWi28/jHymE6IJjOP+o4z98qsKlaKpW+cxkI8uFK9V8OiJGuHerwSYmegMsofz3H
+J8Qb19anRiV6qp+SmlR57iVvluNXQSPUgFIcfZmyuRzHB3XJZkML4ILRzlGKOhV
1sf410LzHdgODICaq3Xu9ljP3fynwkCcNYZdEGBiVKVpfvilVwWp3k3NrX4wzwSk
bwJrYavFET25bnAKxl7MNvBum6mKnLYc0kY2x+phMx//dMnd1biFYMhvcnkA+u1/
nrIBEf9XtB+2fOkhDpDEwQxNfP4FidyFMFPZsQRquwzZEixdtF3N5BNDbY93ZYIN
FJ3dzeXSa11TUrxXq3E9Jb6j9UAnY2MJ7/Z1Q1JQ23gGgEV3g69ma4OGAmEteW1s
i2K4YeaovMNjo0kbwXeeZyadNW2spfA22AjPnnghJxN/ggIxSphnlRRod+CHvrwf
eOBslsoo87cIsUItto9cDV8CxSTsT8DyYrt+JFQ4lPUh4aNvCjm9qUQQfx7dvTG4
aQy5QqjZp4cXk1b8QgHzI6dq7geOcx7O1w6gw5Aqu5Vut8tHgh93m7w1g1vU6SP4
iWvTuym7u9YdBW8gvFfEHS8AXew8VFY7r67v2u1sCPdm/CCTslktEFyOn+5Fy7db
Gg7DjHwFaMBE1wL7C2/EbWSVizRGvAA3S6wvd/6bFTdTJAFiHHbBi8+2MmhfNtYQ
mYMd3Xs3cL1qvXq7sFRqeo7pdJIbQ40NBGjzIvGNZrL1L7jzX7kiDLcwhQCfsMn3
2IH+3gDNj2p8SWjlzmjb4ILv4WYNh/eVOT0SxfKcgXpEszQMauJO9FVw9daWvFSM
SSZP+oM9VS63hjigXlzvutv0Rm12ZHwl08qj2IZzl0JsUxvAqiX6CSspNeREi4Oy
B6oVXuzx2gSTrKQ84rCclT5oad74m4a9bg4cCkRBCt7lDoAt0PdsCQ6olX077ozL
Gz8ld9EUFa32rntQMWeJDNknxmFH28ah+eiiUWTOs6uCq2dj2MPG/AXXPA3eG3zB
hCC4+YzZWJwl/hroXqtFDyhWsXVPFnkimN6SzXGmqAwvV7+F1yf8sDDkM/1f8WOF
HJN004MjT0lI1CUtB+y6lbslXkQRSo3N2MGU/mLSaZn4NsuOiuxgN05QLH3DbEej
Y9nFXcQnrPG9tfooj9sdGi7sZLOTu7FnMXaEfBEqLcst+LufPvrF0knuSt8rIVrB
bUXITDhza61+cfgkUzuw7qEGw8v1ZU5im59JmQlk+S/8u5nQs/FCI2k7GfmLYODm
hq59Xt3j89pHp4rZHWRKWw/Y5NwIwZ/W58K5rI85acB1BqepxKxiavxSNEhA/AW8
TyhS4ZxvWRgfMbjI5AFZW9+4w1gLzJ7zWqcNGc03oBIzVQab+v1F2C71taepxTws
1vyUprhaXEI5ZgDH/g+ikgeRmAdUely6ov21H13rjY1e67thUPb3esFzNExt9yhG
gEchCNh220ZjZSz4Hy1j2PwVsc0BhGlX4OEko1NN9rWTsCbdC5kvu4KoLw4xlUIS
mzvsR+0iVj6wMgZbf7mv/LC7ZkMVD1BqlL3RYZjUsnKMZtn3LE8VwyHLX3NYdiOr
bPknUDiRItryZvwrrhS6SI5VlD3Yij5YHe6lL08hGgWJaiv3AlDXMXlS+nH22RLe
CIfWm9ZiGWIOK4zvG+hizRa9XMQShc4oSoN3PUEj7bK4k4c5HJ7FOF8b8bNf3DZd
1WsrWErQw3iyzbZsNiDy2EoEaq45ShUtrqOK1xIroa6Ug2EIJ7jOZpu2gI4UBT+M
4aI81pVxvjNiA3sfMnLk8a5sna3nY+AZ44ce/zbXa5c6jg7ySeA2eclag+q+q81x
UdNmn2GOPa/cGgCXjUNHKTpuAO7Q6IBEeVTRO+YIGhz70YBqgagxYjRRp7QX71j/
bRFIkTRjpKH4hmvRQultHsxklvrpf7IJx1G4ST2vPzxju63k9XIMclRH4jZ6dCqg
u9UL0hN+Xza9bLAbr+mUc+j4j18mF+EaNO5B0TBisVOjAwEt5hiGn44T7+0y1DfZ
ZwLQ8qJAC55VjNR01Y2kVZ4jYx8oEyM8Lcbk1R1IJ8CE6G7RHGp6sRtqmdTL16Ao
jZX5dJ/IYzWpJnW+1fI37nSth9Iefb3A79Xt6e7FMOO8QB1Ip4CemP3zytOY5g5+
Zm+/tufwNQIvL6wuNHWRRUVe6JxLGxnPYF0L77GRsUD5+zqNkTmOnGmcXol9teXH
Q9eGmZREWB13qFNDecvQL1ZYvR8b8HiFral4GWzHBCpidW3CSj9zI++G4ALAqm1v
tjkp4mSwLwZXTgGuHFcHQbZ3FUqk7KnnTTDlfbSCSMsLpWaCy8GDnhzSiDWo0QwE
gZ48Fklz9nR8t544aPt7dPNhyc+YmyOwKDtbjA4I3tzmOOSu+4N0HS4udQbGTuwG
iCOwGb8kASirbbxCmzeccU51HoKcmCvGUyoBhP+eP6pr5bKm7AfOqngh0Dt1k9ta
Q7JVAeLvKcGA4GiQWy99JzIMp7srzz88M3kH4iswbng3CVYDNw/WtO6AOc/Nn5sl
PK7hPF1UzKXg3XWASnl9dLOImqGDPJy64+8W0cZfjSzYMJvsUCSJAmdjmYVJKgFS
7XG/u0/gsqeyOSoOcfkxXcitrEkGEs2g4XLm3un8qh+ibFED4oeHYCRdpFowiyqK
3G32Uf9y7Nh+odGLuRPzXeKn1Oiu1lJkEHD+OtR2WqvnrwoqHal//zCNTxisrsSW
u7LhdvFH8HqwBy+AZsrlr9oOgjvMxF+Zzm78TyksI6SQvHjNami2ZTBhVgHxNsTd
wX8np+/5c0h7FY65tme1MGfVRNrZVeB/6rLZwC3O1zKXMhpfi9p3CNrb3fBxtdl7
H97VsGTlotbZt99eRy2qGQQEHeD3Lr5AoRKFp2CGPwR9nwECX57QX5Z7+InPpHOE
EHB8M+Ibs7Mf51jyD2nzZq1rY3gxhdBXRdGR3UaJZceedOHfIWsEpnCM28LDVheM
yRymUExhtMds2IjaSvcCnIl8JxrFAAf3nScndaPidIbxoOScRMuW/9cX+cW8wgHc
7rrU8SWAgOHiQ4r5PMHhkzSKcUtdjHXHmlWooRtcUADJ6wmljBZV6kWRi9eY6CEQ
u7587mo20IDlJh1TUIvbp2cZJWDSHeRtqlZ4+WZlS2vyBS3BpWA+p4MDR9D8CN/x
XMDuEKi7uNnxXcTfX/e1R9XvLc9HtnR/NKIcrQrZkxnotN/fovrAJq9EZ1gG68M9
YCxz7GabPJrK7MRhlIfCRMID842Rb/I26SR2ErmLnJoWMYATPi61XgWDw5oS971y
1/j/GGUEk1rKMxBf6AVpNu8RkF6Xt+LixJEhyOWyOBNexKCXjBeQgl2BimDbPisy
IwN/QSXb1Xsg4xpVi4plCfbVT/7BpA8RZYXCHM4VvcstSjlo3rjgDDEONNJNY/EF
VcH7pJZSFuWVJR+pnGaJiHnramUa7TpYzaAwQxUXHBXVGV5iBdqCYcSsQIowOg5Z
472yT+95kxL+4Qzljf7SY6xDqiuRm4XejjTc4ihwOaPAF49EkXwAko9kCh/K+lqW
qdgU7/doyrfmNakK++11X0W+SpF/f52gW5eOyQ1TsBAvZPdZi6FedfdAf1Ckd4Ol
9DDDbh51akgF/CV72CF+coY8mBpQB5doVNA78xZOfwamEASrd1RLqIk9Ghj/kD0H
fEBMG0rlH6zB06UyoYaOt2JwGz+xX9zp19UAwMfgqXKYuLZM4KAKO3yMHelbzscu
L7Iog4qaRd2WCf1YIxHIyqzpOJlWyoKaBDhhpY1QvSJ2/4nD/K2Cu9L6ZKDltWnc
8W9OVDFvQe8Sjv0mxz5fLddDC+wA01vbS9zMgMMiWZNonHO0bl1qG+Guo9jbc2js
+umpYBlXl1EXg8FW2h0Seq3vard9nvF3ojResnPWyaCtOKGCqrbNKdoceuBvssir
gFn+ZWMpzbERS6C+1PEcM/KeCuMtamNnL4e+S2UIC0862uRgX1w+Vb3aluSWwyy6
zh/6N60EqRoluBRiAVoWJe53DzXydDUV3+gIyo7fI7/E1wfLOSWLR9IH4O4djP0d
DtoIb06Gm+fTN8Au351m5VjRECuc1krAdFUFcKzVLTpON+VTdqFspqg+71bR8AIH
V4xBUHc9O5KJVJxebOmmwF1pPsMPB5OX3fSUg2Fp3KTb05MH7Z2TYsYQewglCacc
wXrh+9eIJjz1vMEk1zM+hgveglJ8ykV0JWC5Di2ukKPeFy84DmvJniUtnLKvxSMj
+1YCgzYBybIoMCd0RyyMiqRQo5auZw52EMA5KJOguT5r9jFh5wmtPX3gP7J5dW7U
YRVzrUD8So6X9l/7RA1fpq5HzSlkY6LFCrfxmCMQb/9MDkGBo9H37ouQVn1gQPzN
471/jxbWOOfmiyCRfPBJIryTU8vbV/MHJKpY0EiNe5c6En/VxXc8YprDiHoDObPF
/X4uqFiuBsoHVtVcxxaO4dtd0bnIgf6m8W9WPj/qWBA6CRXNyPSwJY3GrKQ4W45z
vwVAcMpqGAmnQKwwd921c5sQ7R2AWFAxqrc76+HSYs30FMyxb0IeiRK/nIqyClqi
eiVP6Hg/3LPsrJO1R7/w2IhnWAyOyQKhCHQQPBoCxIgO+8j1TPXxWrqd5W3F6xyJ
S/VwRI9hcakT1m8HkvKzFdbE2iLXUEWpi9zfdAkS5yuLwQ0Jj3V2PvtxL6WN8eR9
G9/xRTja1AwgGPJUyAaxwwWn8GI4oFKD7dFsL1JdTkqsHWXM79WZyi+xw24bW1/j
xAnzRyIpdJyLGmvDtPwAzuDSKvWprz6MjfBnSEXbaPE2x1fdQJj/Z58IKZDZdvrJ
6H1UQDhejVJOZ/9eAj+M0tqLh7MFhAaCMre1oXeOSIFolB72oQelyUzNdQH10thj
2SYmKPaZxCUqv69JXyEf1trk5ck0UWZB+xPyVRzLRm0T3KAO6s0A3Us5TzckcHba
x8VUGD/lFqoC1PMrJywUBT22Txa/QI4OGo3g5s0pIgJAgySDzWJkY2BN4h/EklwU
SHqhV8jnNmGyxBltd7e/gOEwx9NTc0WKxmlfW6VmBCqv8Kaw+kX2x1d6/NTd0L0v
BRyjvLbEn7n4dRSF301TgjKG49vxo4OJxUSmOOQyIyMHz1BbAK1U0xI+72XsmS4h
6qL+7+SBvPKJx523axy1eFElj8i/YwRQaqGdnXWYHEnaeYurEAfAgeuc4RlZfScJ
q5TS0g+vcKmKwDw4VQ5uVFO1OJjQzQ/aGSrInPPS+VrHQuZhXM4y/fgWSYYAVatI
4Eq+tl4C8Hl8ILcCHp4kSb43H+SHZbQoiQBZ2U9LFXpMVEG9HJNhPr3sTXMF4q4I
ukEIOe1Kqf8duO9s+kcuaPKPMf0JFiZg08Dz0+TDD8fSVkL2lFaibYPhqk27cPFA
RyL0+PzVQU7oqVRyrQ0H3cLjW1ES6XDSNhQrkXC2lJdxItPSYFGxWuKm7xmNRReL
Rbd8nzytROZp8xSNNgwqCjs7SUlfny3vuRIunKOoSMV5W4vveutCpDTb3kzT33az
yIuwU6JKnRWabO+Kh/eLfUKakMcyj3FBGLILkwagIsRQAQyk0z6kHv9+GCrldyyO
4WZQnOfjPIriu5efTMjiKzXQm/d/RPYv5gFuctECpF92cPV3xWee0SvOH4Sy97l9
TkJ/o4PIrgxRVxmiicH6tgR3gcMD18i6i8CW78l0fv2xRVqtQGaz0lpjrDCALFF1
PEuHdVW2XcRQvb8nCdO/Elf6Ij5C9aeqe4RBX1rEBSDmc8kK5tbCTG94NfoC/V/s
EsPVbERIpDdAB3uiGlBopWTI0/9chOR2u8xwqq595XRtNeq9x6pSQgH4JtY8zh7o
r5Yvy4hSIgV7yNiMRh/hhbS81j5h64LEOg7OxsIu3IdPtEC8AEfq23vw+MAhKpJc
VGWa7NlKgV5SFqstmTd8bWTJjOmoIVJDIqUDhgthvmiCMlNGfRKdFcVShDGXQZh2
3VIpx21+pyr4C57UgT6YfA2DQMySMYWbYOX13kEHq2eIolD2mx/y4j9bRKrTI1jr
e+6ivTSrDXUjxs1VVoutbbXb2Zw5JuuzDahCrMTLcclv9QaHiUAKtxfyIgfHoQaf
D3pLBXnAEytcgr52HZfBkP+brPt0FM108bAaSf6I83iAxPuoG/hf8jDwtvd1AC3J
j3iBE0vH+QKJ9Jc577vkFIt9hyP0AfvN+OyI+Lx1O19XazSAHdLG8bg6+v2rUOCG
y5SPadvlY73SM3idsGhvagoAem3AGoYWepbyA8rE/YB8oAKzMLlSRGACp0MWbecB
r4E+flhLCOdDVml26jPnaanf3tz84GC9iQjkGSXj5EyuvZyErFzNtA1nSu1McY2G
z4irQ0K99n6oO1T1ieWex+Nx9X/J2s91rmeSh0qjNzYcv/DLFxzTVfU9hiszmLsE
mLQrb3GSHk0AB50MYMeHxAo2kV6ocKrWBskZv3ZUDanxbzQVcmUzdGz5kK3P8/TG
ZYdHkKi404DeEW7BRDp2qAQ2wfy4oTNvEYy0uv7d17yCvPlj12ZxKrO4lewlY2zp
IG5V77ErNZ3y5NfYMBakqxuQed1lM0nxl8ixli9KJIPRWmQLl0+QpEcUbRpdMI4o
VdhaptJCkgqJ3L5sbUiRIciK7drWJcB+W2JsGogwXIb5+lBuvgjvZbDsNcD4xKGc
iMCKwpG/CmNGLgoKyAcdvEKLyVoEDOyFM7yqWd/DoFhAQdBxV6FbdPM60asHXuN+
N/R605Dy4UOvuAlCtxm7oTp9Vr8CxD8So7YEZ0xh03terbPVGUr6tBWNXPihkNkI
DoCLmlV+s8LxKxlyU+X11R8LOCVSh8fEkLgjtyqc0p51kUSY7YoAoBiZZqEs8g+8
qrUHsNyHn4GX9UN1zh66KzHcTjjNMozqeWPIlNikjFp07MWau/uAJGpTQVenbhjC
S11ocbyBiz1a27LCcn7ynUGvFURdrFPKIBDoUS0UH4GJ/S8lIqdI5QZuRhcgMlL5
rfnz7bzHKlQuAOD7fgcAJBkRwkCAIbUIsxBNBJQ+oChnmifnrqnt0Ctm6WKFBYdT
enSDJm5p5ueO0BmGKacNIdVrXS8mmBKJPyK1INPDxQICVr+6mMUBjI76NMc+e+V0
QDoiYofxis7RnwOFzU+EalWiF1GY1226CNJPfMH6GQ4Sgy9z866+q9n5Day079ZX
hspDM2R/DNVeh+HvRLUzb2nyYJ37Pq6+iitGCsPUvvd+d5mrRZzQ0OCIG+4TKU2j
Bmnu1BhbIOOdrIOJdH/5kOdFF97TPMa2pXVoUhHwJeoC/fyXAleTznVDRIkDpclB
eOlgqXweAl2zYQnx2wtbM3rTM9/qTwpTMp/OLV/f5VLP1kTClbmig81rvAGXhKy5
sZXMouiylfvuWfjy7POqXaCS2gIN7lv72StGenatQd69/shzMKrW7RCCwYQQl2DF
73sJQuZ2RwVmEUpZG1vm40bQRjDrP00z7s5uGPMFCQ7mSEwvWUArjbvDAV0v7iRG
fP11zACccwIDG/tjqx+u0NazPCJjxAhRe+VzT0E+I1b8rfYB31RX3B0Vq6565lmr
sjGkui1Axr5R3ajLUtat9+zP/Nj59VEuK7m5m2telHnZL/iZCgIvDcLxAB4/TuaF
vknYLIZCNUTBykAhwQjgcZ7i4SiDKMEVIbZ/OoJDKCPzbRicplkcK5JBiGLZXYVj
a4bhZDrzbaAPgD5xWapYx5M+RWChKFvfSISqPAjpBwwbo7wk6g3Kl65TO6lCakNm
/wklkjxW0gjUQ8t+TveIOp0zlXs+SbAMrUXYxeV4+rrBZO6RkCwsLo1ngfcNc9Da
i8dR2cKj8Nh9rYMDdzL9+QGBeaMlWu66Jaeb/pT91Ovpa9pCPccD9JWFD08wgPtl
82HY4cb4yDi3jZWxC4EAsy+11AdQTM0J+SVgEuKvnpFC7qfHb/KUxUlPvcpnqP9y
6rUJ7okHwFM2rQ/ug/iBk4nxuP8XBABTYQMoDuDaqE80SwGjsJ/im5BIUJGsxWLm
by3ZUM2yHzcSbrD6A/SrSytErq5+n3ySkA8nrZ1VqF2J2Rrm0C3ct0+jumQ0UJRZ
6E1jsVB7W4LuvFaVv8cTZQ60rGAoNar4K7LT9iqQGw8m4XQ7ctYe+aa3X/41ML9I
WqQG0TkIffKMmIqASz5iIkijbZ6+riKTHZkrzMBRc9jE5faehKRvPOmF6B7O3f+Q
SITZg0vmRRvP6/YCnG+9Jr5C9HOgGw3ZSXt6JUjYjmABG2wIySwqgezAKft7fSSu
dw1I0QYACheQUwbMF97krrflmePv/xHzCbDLVEkDO6ZC8K9z7qf45Ga/ejxRalz4
U01TZrf5l76nqkG23fOGANbu/c52LlPMlY/uGFdZhp0uUaWa1s7MjIBLTbe4PxOF
ak1Ry1U6bIW6vUdpbFfDtkbZQRuoaT5MY6WfOCpuo3UBeDJklBq97elAgJKQyjji
WGJMJEsmP8jkVMTyf6I7sM+W82nWYk90r3cyFCcBAbJA5vPI4oRXiAQoNyKWszyT
lWz1Tn1fe5IhNjHKDSsLBf35tiUSNBk5v0fen3Gi/zR7Nqxf9IyqR+jJeSRghiys
uGFVwC9wlbMY8NiDbeU05I0NBawzlc0KpoZ+2JJc0+wq07+YxiAIU7K2qSdT7tXa
/z+86ZuJXQcyoJMPOlNBYsfmPcLZJuf/CP/OJoGPpgU2b9IiUDqrdcvpdFpfUGBz
Gz4lg7zysO3AL7rGy+DT0xWLcW0j8B+jRXpbuJ98iIr9WcAcEJUdhNsQmcuvc+0E
DbnLChWlLtyOLRJ6bMlahdd4FJuroD60ooHa6OnmJp1RB+7q1Op5mngvLEOvOqrx
prqnsTIFwXZ+OfMCbxydSVq7bgIrgzrNOaB03edqg/RCRL8AqUU6r1FreLfeDZnw
uYPC5RVhWZsnd+rDIC6p/RE55jg2DRtjeR1MuK3eQv54lLx2/pnUlWcOCK/97YQM
B6VC95VqORDdJZf8Kifwa0H/dIyYbxXHRiANPBglt1pRklrz7nB6jnha0FRI+JXK
e0gwXAfenGUSyt8ZDXnqZzuhJYoVhy6sDbugiptOg9dQvT/U73X1ZqN86PWy2Scn
6TFI5iKXuQuZL7HpP2RUdcF1BDi2m5n9mVZ/yjpoRSjw8Cose18H16vjd3Eg7KKU
9S4wDSJ1lZQFD6DYjEhjfAu526ZgcMWzqAc/cMHU99yz/LghmhVwFOWlVtcNytd+
8bAuqCf6mAelgsSxIK2WOI2MbFzY4Yzh6VWTYquzuxdfasLc3Vhv4uDCJCYdaeTn
/chMB8m1bjNV5Lc03EuAVsVqiag/zog/gSLq8UOe5B4difgIpvpqUGNGLrRshrZq
TCqDwj817huTDEmgXDfz0IL7VoaCz5fkQVUOmhkFi6lKvtidwri6BFVvVfPOK5ak
jwp49+dAdiAGyneJ77n5st3NcKB+Zy+AdlW1dw2jfC4z69BTHjhyTmB/h+QImDb1
CDAOt1szFp/1JY7g65muYOv1wpoX1U0/wU2EoVS1Ep6kJKT/BL6AgWFwO544/r8q
Z/aBUvZdGqxWpWag2F3ZCGosjcJcAIg43LiWb5GrPViUCob/XguP9pCnPgse9RVV
+b3yxkRmHDwEJGhTgM418hfeNM3eBVv7Elf7VTnkcxKYErPelN2u+Ojh+35iv3gq
XKx2BzqMfRr4XUoVelURmP9RYvsZ0pmV6aRLG4VExC75tSVTj9pfpaaqm3d+A8ze
tfUqaVai8qucQwyLbQutka7Tjvr8nQB2dZC0HI3KYYE6mEOTrzg4Cmis4itLOs5K
iwYtObK7326DjhX8SqanPaiE8UsIfcMbM1uWxy+JlIqEcbJWmVMg+AnHaKsGNN6k
iKtWeBqoKgKd5moDPxsHlW/1e9AjhiQS/qJWrhKSUx94j/cmNxC5rDi6b6QzYUgW
nGRF8hrUq1eRNDTyG14uKiENrZ2qWaPzLML0QthvDs8jDQ+DtFUFto79oWErMdCQ
Ejr8sO7fRPS3DQfcmhrEfNhjI8lDx7lI8CAUHOUwT/FMab9D5Z5Uy7NSZvHWXu4O
SAUMdTtHPEpHP6LJixW5fJka2FjzAmErCzBNpmJdaFbSoHQbqJra/fu5RA8QfqEY
kA5qqBFMtf6PC+zz2wbQ+/KSX+eeSdP4w+/1PWb7l0V4TCd/v6YVZ/5J8h3PmOPZ
VFdbCKRb0wZzBLtPs5SEe1Qt6bHxdS0LWtS+Lpt05oHVm80g8L1NXFEg3cyseamt
gq0ZD4R2dI6hk+IdRp/t0Y/7J3pmLqfJmkjW+0qacnMyWWmcQhUoLdtYqlFsoVjt
h8194z3EqBdefKvm0Zqhra1kAzhxLBdb712gN8CeuZMQ8C8QAaI3SKdmyqkEVzNs
7wYjAoANi357RDC6xV7E6m0J039h9jPQX4TvfUR4iOEIUyCIMaFgY9Z/WHZUQ2gD
756wLs9zPimFDYnx+o1g34SIdyMyMON4dY5OuxUg56vinCH/AQjHbnTqFqZz3tD0
zwNi6bCSsJEPwWAwK1LWZL7H7jdWweEtusda4skqC7wCSFmdzgk930CKOYdEvWv3
DXFqrRlhjO3K+dpT8VdqPWKAmqbeLuTLI4vTbagwjTspur21ML5zh6xT3hf6E18R
J3CV1rYLgM01LoNj0gqDwGXXliaVhZR2UaeNaE+babUvOB2SfX5nFTN/enwvaBZz
lK5/rYEsrl9pe76KW+/0x/54M31YcdmIpWBiJI24QybifHt/iRIIcC+qmBksTBZ8
rjEWUBt7gR4JMkREkexW7BiNohzJCi5z8K3yHTaHydRPomgMM7O7dmwp4B6ABXwy
M0HNuWvcUVcrjzVxEdU98bl0hEiFooZ9Bvj+OZdH6lBc+p1cuIyUxQ9LFACfu9C3
L3YLFIELP441CmSROAZyDOSYCCeDMnGU9dFCN6CrZ8Mxq++1p9ZIuAHq+OWIU14M
lCiVevHqsE32Ou9H4WIfgLjhPNVVekyA5gceAko+neITBZbpVaQLiv15//4sXdh3
RrqmJ2Vgq6q8+yKydrurEZnoLZgKdqZumwnjqPhfZfw8XWKSPcRsfQG6ms7f5YqG
nGTSOy1kM7kHvn4FuKByDXkUaw8ZXQAlNblV06JmoRUNHYZo0YzLGwRgQNaLLpTx
tt/TeirBikJRFIr8ZCsDVq5G2LFM3zfngphBS1RDbSCoHqOy8QOWO1WMd2KG534l
awC2Mb/pWic1JmDi1B2Ag2nK/CA12uwLW/eC4cgIRvVNvRrpM4aAgfw3YX3uQK3J
eSn+d0yfP/uqMlCR2AKPnXGvFjnJHdFUaBY1sXwKUeOglA/MuU9enMASa+6/YS/b
/809d9ANEZu3OehkL6k1nMhyv6Sm9G8SKeXNOkoEEETEwlY/J/SE/XXnchOdk7pK
inM1uY+uCYwFr3Y7JgyDarJCaHYPKOuWcZKblvhEbtzGmhGoKTKRmNGwEejfORvX
7TUC6294l+nWyqXV2x7tU/FS3ogk8uHfEYSgh2z3tOSfc+IP5PrUos5Gce5nsrrB
crEdfHuU/oGMnyVIEJ4cbzBrEJ7IwNocLeXTUmKMosrmdslhWpmWRAs1sxk4RfpQ
h21qHP8CDAB3fLWpEKvxE6SO4Jeg497Zz64O6rxr085pJVxZuXcrJVNb2FEa4jAM
JyuH8NgN35iwoiHtJ2bzYvMxCwZ5bFzFYyFti3PVdKDZ3q2BJpgs/FGL9QawKUB0
YAT87XCWnJS11y94JDdH5Q73FzkIeI4BJJH0WORwb1IHFdFI17wI1NfAUE+XPBIQ
n4VWcWL+ggMvMr2Aeb/Y/uDX1pHNP5NNNSxgZqrp1LcOmJ99jBpPG26Z+5Dqqpmd
KdKj1x4Xf4mYn2sSp/yu5MvehjIOxt+nBk+Vz02x1RJqaNJVcgamydkzNnCT30f8
izYDzo2RpMTw7ICzDpKID6GGvfqPdNP535X3LVCTcHkKa+29IZFSv6hGl11lgDZB
La69redzwAoFwsaUwrfHVEcUidr8seE6IPGU6zf2Cre4necBxvfSEYCv1Vk3XZkc
T1N7/Qk+lvNUXDxSJaoQ2Qe8Hg+N9Ps7nhUNhzHHp6tzvgwsctRLZLOG9QZ7rTHz
9F7DXUkwLGaRli2e1puCGcslOI4x83e5oi3i/IJLP9BMY2mAm4HtidKqpcpVEKqb
pKTWblQ45+GDVgT7jXP7p3U7SFy9EAZPlA45+Mq6zsV9mvb+t0P76aniJ4zpNc9S
1vp4WPF8W5g7wJW1jD8bwqAINTsvbYvS197oSlSPrbHCJncZZYByTjS+FrEcBFjb
yqwwXl7jgQgOhhQrOO8ynCsJkJsdziAUd81A5/uvLoEWc38eiGI8otbYdGJYa3OF
IXYI6btTUtFKHxwHHGjX86MKi9Ah7MmdQzkGq2qSaecDuwZiEObsJ8rR5As8DPuQ
RncaT9WAGoV7bnY49IhpenIc3mwWl/ne6Ho2it2niTGya6RkZF3FNazCcqaaZwph
0wnuV4n5ThgQBJ8Zkw5yR+y3WzlRG1MLKRZC/aQylIZaVnpfGAyBu1vjZCuzzepv
Vz0KqaDt2vSVOhKUV6+TbcO6vJNZ9sfCBY8WyYM6JQU1e/bP0bzhw4oniqqcxA5a
PgSei0sGxXxFoMNQ7OKDyLgK5KxxGMy5JDIs9Q+y7Zlvc/nC+UzNe/b96Sh5dM1b
oU6UnUqTpCBLbIi+hj/oNJWBZSLBERrENfIxGp7FHeyvh3UEk5djJ6psH8wio0Om
ppTudpTeXCuDqzXe7ZjxgZbBpLDU7/ZS3+l77+xQAtC1/lTey2/fM4pnitCl+tTo
8LOeDoRMLXG4C4vFpZtqupiAHkbcYF8/iIBpHKzW4+pjNJsFQYTPeoYuMC9+cl0P
6dbSGL5ZNRnVUP+BFhh+aTLX7sKKAQJ+W7eb21HOfgmRMif1wIq3t8+0X+pTxR4j
BSqDCYE6CcPNDOMRhLinYYXdN7tNJ7eQIbV3YuLWOueM+oIuavHtz0Kd05u53Wha
CTqWJEFKifcq9kBm3jljeUUtPdjHDvX2G7UQsHe+lcbA7zuLyKVVQz39Tqp+Jg6M
JklpKvWlXYgtVmNvc18vuH1QJRrfUu4IHTxb/94uPCHUOLnok5S7H3MUBiJf31cI
e7G7w4aX9QTTBZRnu5YQOWcQ7C5Fb1LDwZSSfuSIo3FK7ixcV5HNUTSh6SAGkMtK
cAt7nuf0R1I600TSRmplQPGG5WL/P/19Tg2RGrM1tz7DXJVvyFWsSwOSm/burwYb
Aq1+BL+5E6LkupTiMKjmW0qMJpHgbNrYN/BXStfamVdRqUF1Go1TEaieb+w4Y0Yu
goQ8q2Go+jK2th84liOYPKfIiGE0z2JvNglA7LDTNMDmLBZt8HC39OmLw906IY60
VJvPezjr645lUglj8UJ02j06b8LtSRy+XgfHC7SKHkYU2jzVtS+I1Qnah6vRoK7X
3xstvlvc5+sl54nWPiSAP4X1mxYpmNyjhvV9ex5ne0fl2IzhcrQEDH8MjGEKzBq3
y7YRVWVr8AeJCFpouA/Ep4WPb7kq2ynDPG+8isKh0robrr5/b33Xd1kvm3gjNtZP
StaTkToKm2oIjThIR2cnxos3hXtJCVe/E8ihQpV9ikHclDVFVzoP4bwHUFuFXuq9
3rBcZo8v4pcxPk+q9Bkgw+AQ11dGVKHd9sE6KhQt9acnFSvrBuuvvRUvDVMXKhh+
akwS8tZRnPfygQ2b8I2kpqbjAUZLc62gIZU6G/cFSmcK854HwjO1lbH/r7fmRsfl
evTr7tWxMz6aG6G/IbzGrIKGd8UHF5TSci9SaTNK8U/1xdXPNvhAkuWafBqQlySO
ETWTVrFZyzqKVSWWYdoX0Ls6fegqN2BYwvbGuPIgxcdU8iKF2n0WIXaVc6qE7SAX
znsTlG6o6pZ5SR6OlVbcbQQs65FJsHWHAYXskPlRdiDMK0h3LwkMSP3kPZS5mzqx
NNgmvBLn2JH5wJtkUnrATXdtqpaESpjZjH+JqYDTmRz/Rgirwm1pdFZwYjq6/nw6
++o+D0Atu799gQRHEMC9Ix3OfNOjuJaOP+A25ZEnF51cmFAWEWAyWv6CoN3Wequm
cShux83bLfgKUWYbpVP29zS4UJ4tO9ubNGvmfTibH8+O6i2/W8t8HGerI7pGUyRv
OrVC6Xf9IcfzcA4trEkjhDa1qaAcCd+zyrwSZUwmRUfA+TQpvbkr0g1tdsgSk79+
S0/L8nKieUgpUKWzToJSsAGD9MTKop3N0Tmvi3oI9Bll1vGAwa/3lRz8WXIjfFgC
y0f5PLrSHQeIhXsfBdwW9eXnA5lVe0xsBA5UThayPz8tMyrgpDIWCLdJXtnlHEBY
H4xH4zSlBmXaGDJfhjQ0BGb7tz4xWV9WKwsTQTBLjjrftfzeh2qy+18oWCubc+05
NR8dl7UFgniGb3w/9rFGlp3oBvlK0OYW1EW2p8nwgpVtTlnDQmDASqqJKPR5IwKW
8we4zi5U9wL3Ncfbm28b49+tNDfyLEE0QVf8WAon36b0Zo4/EA0sHvmA/5yfqX/q
/iVenna3JXWSL9vQB1n8aUpdhKX03vXVnsoDgIN1yH9KyI4iZMiMIS+KvpANL0Ev
Svj3sP5g4ypuFkFTRYxfyRllwxPBnXk7KawNM+S/xgYugYTOtlZsnbkMybHaRZpb
X5ylsLGtN7DsFcGqruxiNRdk+PHBbtwJ6IzSLcBLN8bQ/7q2V9SbUzbU0YhC53M2
rJgi+Na3BIw4oFZu6EnA7j28MA4jEK8ngTCooG+niobpbzFeV0jOwPvH54ALmo2F
dE0cNayacCXIcP4n39IdrlyjmmBoCtPB91PcvJ/YRm9zQOx8MvUYMa6FBYiheb9j
yC2DnjcrjnVX7Rj4lKb/C0ZlkP/e6kwABEl+EwRdjkAoxZLBr3CVHFyLzGW08yzu
c3N09feV656VZQeCB9gJueezkBZUYiliG0Jh37GtNCA2p4uAyk6AfVb8UAqhihfq
TvmP6M4WpjFa7lPATni8Tll1pqY6SUowl/C4yhJ2Uhaj60GGwC0iZFpbC1w3wInG
+/3tUHmIo6ma5jXBhU3FMNqsC8E8l1IMeuh6rauMniCWcUG2hzfFK9yQOwYdcYeV
lb5Lct/8tSLyKuK2T/t3FLhcnVdpOPGI0AbLMVMJQ9Ym0hYNS/3GzC4tmlmQzob3
QUpoS/2X1HGFsgHzgyKUnMTFbdt+Ihjk/+TpmtZof9Au22EJ5PSUm63/qOsUMb+T
wOQDCvJGcLAfGMXslRAPAhYmgLxQaOv2mDxMDz7zUNs8u1NWuRChUus0WKkiskpJ
glJRkszhJa1LR8nzMi/HT4z3SaP0wlIG5dIZIiOJQpV6djCPcibPuLm452wPq0mM
E7tOdixZForXc1DsxUrrpN75dDfNRUFKepzvVnTsAXAHMzDImBkVc+Km8tgy1Ejm
BYdSpVpWq0EqFv1cBpqYNca/hiL1M1vKLOtja4llKenkReVI2YoEzprveaQgWamG
5lWPPhJvPuotvued6PmChDCgzQbz0WNk2ehFSX7iZUMgv6BwMdNDyWAWddXn8Ct5
FRIUefuzXhPMCwwC6mB+Vk5jZbDpJUBtSxchA9uBZ9OvY9OLSAa68aODaV+Zlr6+
2asytCzXF8gmFMtY93XYlFa0BS0WRTKrm0ONKJDcQ5M+IjzeRa3iKcI5tdbL0Vta
Htx+qveqL7Jh/wmteMGKNKer9PP/iH6DazdfXbD/Cb0KdAQ/EKHdQvJ/FUMhF2tx
sGdPsMvB17CSeUgEieXl6HwMtjZd2Ee+PUehu83MIOQkEgb44a6c0qsZZxuF33Ru
5d5SVTgBa7y47khhx/eUi3zfcBKRqMWKc84cru3xSD19rAbVl6HS2/+H/gTpQW97
/ZosPDko6o3uokFre0qEH6zxJcXt3xulpqKTZljHQVIVFCVLMEStQWWaDATC1LDR
QU1ukhIt+BCYJeLAY6FpFJtM7kVUHCJQjWJzf59qu9HMD70BaMWXfNp4fA0elsuG
kqcN+uvevTRt0bzaFIGzZdY/3llC6JpSPvy0mEn6VHugaw5zN8MUzciJBf0q4Drz
x1CwADq4sdGlTXjZrTjm6W9QExLRLePsdB08o70ncRXxyqUOc/poxl9yBR9TfLAU
KODRh9+CZMlgnSmVLR/mkFqvUv6HIyVkfhDwrC504IEvXkphu7r9yKRKpyBGz0Pa
lJzRk0ckm9nc79OITlfxxHjk3hq2sWontIu5Hf3vlGxzcVAW7r9KHR6bNwMgJmd8
IWAnxt8cBqoCczVPl6MUIDVviu3X7U9eqOVUXEt67GKgD34+tYjhqmFl6ZkRAn+T
53tw016GgkDA+cH+wk+02RrdEgsTGSlNjfaQQ0U9wrozAd4c0zLTCs8AK+FgkH5I
Dm88UosVZiHGn/wSqJov6Ux1CoyzQiQADMAnmertotm9aSIYqJq8rteYzA0R5CuI
8vNJ8PJmg+UQjHNGBAc4r+Hs4E1fWeRQ/oXtWKPoivhCtL7wiq+nWQgZjco4LxGP
wKgOD25oRFuRCT0fioafcJtPZQbwYjaNAkFLovgXuuTwAd5oy6NPJPrVDjTxbfcJ
JCsVwLruHy7YXXGtvfdHmSzOR7aCfbGoXKG/BkNOqthi0nlIZg00tNIdobaoAMRE
svfWE9sPkz+T6HYrYqht2dHxprZKLqDwrSyfbYmjBjLbVcOqlfhO4wc6iG/G/vfC
ppL3y9dDQC2RucbxRwMcHl6J7SsIYhvrf+dwToebaiqFLsU3F18ILnpmQ77NyUsn
PQ+GZsDDtEkeN2JCq0tVlKhh3aFdTNv9qBHHFruN/N0Qjxj4gxeqlXLtsnfnvoWw
aDX2BFBcy2Hty3//SOuSlTlraNdHqlTsm+urSJv6o9FaFcxgbo0a1hnzIXRC5MSn
bTolIGQX+GP5HyyOoKpoU1AELhUN/l+Icagp9Sg0qugoY+Wlvhc3crw4DzeEb/Fc
oe5LJ/Jw7je0PGyIl4A5Z3rUnLpZCqZUCIwgFTS3qxZ0f05a4tYtuYpiQ5RdLR+J
A2PbgEKGu9TKvPaQRCJgFfxvlPikJXSpo8CehyUkOid+PwBIP98EXds9iXpJSuA9
aPtaHDwelJ6AX3nvvlg8dewSB+voldMKNJADJM9F5cgE0wwxoE4TikxUIKlrKWxT
pShBbtuqhV0TOFGmvPgMTI7s/KEo5u9/BBj8arOh/How8DIoVhxlb5ux1Hw2gdwX
mLkkMU7uXUDkr3tUDQM8LdbV1Qgg3ARQdalpb4TdOOazdjuTGDaLeHK2Vs33Or5k
BYvsKnmRwIvlNLYMrWYl9Jzsp6Vjyx7iOr7xxSG7x+Zniclau1oR6tB+FWuVD2U0
qDekDmCqKgIZHoUgX9edx/vN49uN1zXbyCeKUoE9Md+DEGeKENRgvC5sQzoOx+ni
4kVTpt9OlWAwdBJpEljt+y6LW0iRJmi3Mj6o6crmkgZu3UW40EmKfLhxggjdge9w
P5UmoGhh5cy8sXGLmX6ADLbo3TrydAnRx8hmPJuJ9/Wda+uyVHVyYgcG+pSyqmjY
qjhtFfvkF4CWjbhQK54ku48BQAl5d/arsDvHFnJ6/QdUCfwpMEHFYVmBFTsIQNch
rOit0Xs3VmNEy3Nt4KKIsTs+/g610f96ZB/20p7W8lQw3zZFr12k2AxXJLFm73PE
lrqs0S9hwV/lFD1//87tg4GCJSYZ3YxkgW/10+I2S6NBsIpI9pmJBqpD1mzpmhDL
7DBXawauzMA7ihVMUZ9RgATMifDRK96ZfD99DlbEGVJ4j2v30CQ2aJTQLOQz8kQV
Ze24xWX1FHjzJ65kQRRyFJsItajuaZKxfXXAyFRh8nl6zViBxF5ZGWAMbrQomz45
Ce1ai7i1pNu0c0d5of27dS8as5TLyfZiKP8nFmUgfXno61beX0ppuSTju1GKfWK+
L52g5Evn8Ob3qtfwu27INgogRQ/5ikCBdPFFY6zQhzE4Hznu7VIES1S5VTwgXwxd
SOwNsGU8/AmP/mPCs0d9gqonEEiPI8sI/7yIpRAgBoA0+Y0LnF5xYBTkUm4Ij/iv
vO3bILtwB00l2NMX1RKrDfKWx8mPCOAg1HBK6v0t7ggtLQGQtBRKdsDEeZSOZugU
yHF1ThJwaVadf6J65p8PGSeSbISwvleouNYKStLfAleKg58TQxBSSmI9ZogUwKDX
nFrtt3Qa0ZAl044L4n0xSEFLOzD0qnDg0DxjpCc6Mdi1H/woBJSLwl9HXaBvihYJ
WYklmWUTJDzlu/t2KUaGmlMhYpk1IROj30nQk3MT75KcX1K5Ijq6DuXItyCyHMi+
fmA/mDiBptYoS0jzFPzGi2KtDU84ASNGH0oXQtZjPhOtQRY8tWwwwuskQZMYJolc
2OVMOaAMFPs3d47HfIhXokIlZlGVyxCyCE6D1V2ixeoS6aur9hqPKudQP/o332aP
kOq0eV+OoxHFpR/PLE5geLeQXuyAXMxerI5m+k2a/QMomHNXnr0+rwe0dy5gxdWg
+WwB2Tn+ku9T1zw3B9d9+c0ltuIvzXCKlQ5hP0fh/M6YmrS2giT1WwIF+tLkeiFj
8fRNlS3gnQ51m+ECZfSpFDMzf9W8bMefOn0HfskBhakmlPFCXzimjt6cB8A84blR
hUr8vwvFVvJDxuuk4SCvx+T0TJKFZl7hrQPJy/6piX6X70dRT4MHyiFc2kTtbriY
/MQM2L5z7BLQuod1IskwJmgjgXg/X+YdmI1OysNqr2+wUuekrefFUWRQLvYofsOw
L4PhJoqUdcXZKvtcjg3luQTn1NtLLsXF9AWm1t1Zbg4bi3bh+TUkHmTMqVBTnBt5
1ion8fFdE22iIIuri0W+tx5sBy9qJM4wxbi2elnNae/Aob3wSt8AhDtjC5o8uYvT
GZhcjIkUl7ouaOTlC03MLCJPCeEoDkLjq6m1ixhO8fLW7NjWLBIDzn5OylYXS3rY
2YkmnM/ZuP2+5lNhkOaKAage1n1590zpIJcbZIxeU/j525hyLqa2Uv+shvcKlBCu
BsJttCupWML4hcO5tnRXjD1VYt2z2TZBVqjyKtlxPb55SLOffS1CKkvYTbtzP3ah
qlEt7PRZB+Q8VavtrvM5Tyz6PZ4WGdlMOjFm70gRiV6oRhTm/8JOZ6vTjFf1N7kJ
wRJPGHdsz7DX5ODBwkpBz+twNZ+hUnRKVJ9YP1oOPkXhL9+o7b9B/LMbn1WoX0Sg
1Sh2seNdCdJF0VPIZFCNXqBmQbzEgEcpq5YBF72KX+rvNNh/IYx5nJIi/0twlV0O
fAAXeDFK/ORtz/sQTnjnvEAZvya80u8fHfJ6xsDZXeQ/l+6YK5ToEAnsDhgPTf+6
PYq04YEzeKKj/X7wvGrp1asUplP65CWbAIIBzTbLf9ms+X7MAa2Nm2dVAe1qmfrO
fIjvWIvw4spZRhRWDFn1blO4FCZaMLg4VSLdSISO27uMUbNKYq70Cu1xdvkwEPLZ
qSyeU+ha9g3hm8fEYKmuNZH74sZOA9nHHrMeiuSLftow1Z9sQjs4CCNmdirE7+d4
i3cPBNyJuYNKRmzkl8iIDRQ4YI4S6EnHMg1sRqbPffq2DEfCLK1bABDywhqO8fD3
OTeuxcQ3Si3DqU0svMaQKXmPs7cyQxhDuf/kAVX/4XmYc8FCHza/Xjz/breVAjKa
98XVPB7h6M/ICKIFdwIRE7mlt5pbkZ83MTrPqF3JvgzkGiCGBF8YtO8KH+/ovg4W
hfLtxa8/GhK8Upv6tFyTPqdhA+p0CutL6t4FYP2lblMmFh3nNP6vMLgosYA4ZoJs
yPYkWgc7vTVWA67fZBXWpB3DSCHCYe2FOub+FVpWOgdxDejuN3I/VYfhwJAyDSA8
BQ4+s4DOuuY2HIa5ZM6ThdIbzrrwKHABdRUjLh7wQNJuvxeqio8QYxArwwaEkVDY
YwUc3K9hX6ZiJ0Y8L4677XNxZpQz+mChQIupHD/NVYeCyHzuwgLn6D5HrcV01IIs
tKoORIGq/eqkna1YUZR3PO/LGxEMmoGr65hLidwyLAGBBR95JBdF0+FZNsHzO+Fr
RkLvJn558Rx3pZitpuuCdaY77eoyPv+6/ktdNVUbHd5zTrUMrLmemzqtT9P50LEh
bBTZQ38RTwe/kCZeLJvGsSqocpxjcX0zilH9/ybvhquE7F5uOsUg4RviM1JP736f
gGqTwLRjM0BJlGfCqf/1FEJkIRejIOO400dUEm6BLSx7T7+iOdw8J8pGx4mDe0LT
eshVN/6dCtPg/FNMngFAMQe3Z3RVCW8avhwIYts22kJf0NYJ0HlPp4vLLmxNy7/i
4WtCQXtX0nu2LBiNO1mtqUmmK3A2JW0zj5evnhzJEa1ACeH2gkzV1C6pduSpb1rC
ok07V0mLpvQgfkubXoHJOWrkFKAhUwgp6SSO4s5Mewh3ynk/JRusFdxlb622YTs1
wKZXW5zkyzV3WkNxZvNWIMrR/VOClGae3mzpFw7T5z/qKE1Xcz+7spBW0jugBUTP
3ALqL9B4+iD7jwuaIAFgw3bB8XW3OHEAihYkHIrJMvvSbhDZnCQBV/XFw+RNF5ZE
seOkXQxTrr6/bx9PgP2hDwGof86+U19TY9l6j3IevOoq0v5UeY3rwa1EnuZPfWod
oCOce5PYjf7wrJJdWgYSIajBIOfDmKLbO0hXt3Mwt5uhr2+Zk+pVc9xh2SihkJOC
Y5lfg+Knm20Xk6liw2BjMw/fRcF3vB8j9+7iyP/4wq1bHL8aF4kBYbiXV0i8ymh6
K6Px7rsOYpnSMjVlt+rdgrtvVpdNY+FfVeKgKh/gIWTjR/SBA1BsHkjy0VUvI3na
jQjuaLJUsSmCdmUis1G40rbbSSPPi4iW7V88ToauYUeVwOxcupPUpAaCLNtFM42T
HLXxQOr8qjzsTaTaATBgBheqPF0dyQyCoxuoVdVUD64EKTuqKUF7yWqT86IKIC76
3NGwKW6O674j8EnpVu34NXKNczWIhginYzK6C0TskQFRSwQStdvZOmN/Cd9mIkM1
IObNs44BtX9b0JY2Supl2MSzKabT8dvp9FTyGaYU7sCuBtBPafRsdGPiLswJi7zt
DyTmVkKiHDlGlgitgBW3VkXpBM3kK6PCIAYCnVmbu0An1f0OGOBoMxa7N2RCyBJ5
xMtXpkjsewuzcw90IgqyetzniMsMb0D+Xn0Mna/tZIIYJI61ih4lReZWAER7H1yA
xBDyDKS2cHCAi4G0DxDMFCTqWEKIYga8bjdNSki7UeE5W1RLqa9p5l6NZ5ZEKOdi
/XfbpCFAAhHLg+3TFstf01vFqbYBo9ejv/C0gOXvoyNTXi14BAUq91uODtpIlkvd
K7nYsIrJZo1+f+VGc/EyKqynAr/osubrUNBcGUzZbondZs7KHcutkVRmsC56aunU
S/1SDTCPK+j3wuYenYh0r/Xjp4rQXOwiEL4u6GOchpFa+gzfsDTlJPHaAo5OlpYH
PHN3mbJ8KozyzAySegJSBwDaceActtSPuwE52EmXKEj2lOSE/PR6XIbO2C51SpOo
2Y3S6zkJj6dBe9Rwo9xc0aYZI2JySPacbKwXOK+g1YnzUrLu7svDbl+uFUYArENm
e2Pm6r0F16Q5p1wTSs920zQ9O6On7it1uKGmQqCAXVUEJG5vhrEZ4pU6jqLQVqaZ
y/qhFLun9XKacOx7k4AA35g47FLd/dl5bk0bKTl0lqvOEmGo6yGfH/gM1fPFd7nG
8lPkziAFUXG3bNzDAaXy82fbXyUDSX3/6YwyIDKf2+gWZMxDO6p06tDnYtY3nvIv
kTg/A6rebNQh/UVEXYPFzaT8UoucZm6lsoN/DdGZu/j2oc+LRRZACIzBslqYU90M
cRZrYhYq3nNHBJbwNTcChk0pNSwMTIHPSETD8m7DsURtwedzmJT0nNIIWa4WwGPd
cxx28Q1hBQCinm5S4dZp8TG9pJpnlwORNejKiHPLOpY4FedkFoiV4+XjHJDqHF0l
g508sjNHyILPurZCk6x+ZpNcCiwVqKGZc1Hbeho2NbdmIQp6S0bvhA8DQHAuq6E2
lMBFp6S6SBiQ0D7kPksVizjZ56BcbPnbR4B+PzRkjswPqFw0vKqxxV40KbP2CndO
zLkKQytMegzsPSIjNi5YQSafmw2BFZeGBQnmDcMqJveDBNWPmX8u3bwtYW2w9026
1GqPQSmDPVw+vvJSl3Iy+qcA3SpIAoZ6KXoPWmpcGRLcA/79G7gLr7sO8XfvtpQ3
smajPpaeEM7j6frzv80WLln7aWMI4W+w9qsy9Lvs9cwqCM+/26urOg86DioVb/Ft
RUtqrk21d0xeBtK30CiYwpaSS2WHCo2wATH0YCE9fPAbFk2s3vFrQI6uzSNhgLiq
yNBlW3MwFe5aOm5sh7OuOoUyCRstKR+Qujx1wksxL1uzMjHRlttcT+7rHzvXO5wp
ezObv/Ir8jOMtwBkOhq/La3CXiqjik8nIdpH8NPYgqCtqPEtR+pd88MHMTpdP+t7
CMVo7F+JQqb5EGlm3jkggh0lD1TXJ7frjHQ0k432PRyOAvKIOBB1b/GpqYadILRg
GOgjBxpP8kOlvlQzmtog40L0UL8+1zNgyWb30GnYgTbpGf3PoWra5OfiQEAnoxUB
Lo0oP2z+QpcESHj/6Lpdp2r2BPuPCKZSQIeajMdb623tOe/iUziCY5EcT9J/AmqT
YKHlF8oXVf27Q+rVCIvp/smGipoekWxDjV3Bim/zOvzhZVQnZBURvdVoGfLNKZqC
Ndao/9f3tYS0gM9HPFgs5vJXCMPLA20SNdeW4ShjiTJ79ONzjqfXucR9bWyG21Nx
IXifaqwVxk5LrW+2QkK3or2B6A0gxZdqC8UF2wJ27zidfbF3TbKuG/hd9TjnITIC
XEZdQwe3DK3x15+D5HE4AfaRf7aN8f//AId3P6rvMHSgxdQI1wE4r8r3d3AQ89IC
6dtTyyVTMgIS86uOQgX/YHYKDOkLLw1Cx6jaWvZ0km8b9BS9gEH2ruLtMV2xalep
Jtx+pwFh+3nykFdoaxVs2fSAmRGL8ACAa8GwtkOh7jxQe6R3QeiQSuFi981wq3ES
VLl6TQ/Lp9xAxBeVnlCSOwTT5KO8+IuToUDvGF3/z4ioPUVLPk+TE3CR1vlxcMmD
vTbVAczpVMQl+eNx1smCNtbM1xHUY+AiTnnNYIZ/OTRGTirrdZBgWxAcfcfLNYfa
siy7UzQrfcKEOLDkoyMgTezUm4GSalms6fXlhfP0fgzURyrh/1TlKhU6TPVkbKdX
l5X4f/1Kg1C4mKTtiiDgo9YKQjtKikTpTwzKeMoMN5Y+ANHKKuX3JaGZmZ3txa+e
y7B9ip06VC5/NPNp9hddgK3dZy7oLCtx1ZMiACwwwWka3fooUFjQel5DfbMKvNKT
zlpnQxcNTqvebUO3A787eY/7obrDCU1ALq3Vy4cEBUAOgFW8So1wtcWTU6G02zPV
C9V2bgYPNW8cYcJMrNIUIA7PhXHqWPCE2jXh+C8f+pPQtGGfasREbb/oXQdfUwI+
JYD/FkbkfFePKHEtZEwqlkavDazCDdOQsHK9s14NOhFFBxDdrxK9AIlMA+X+oSTb
XVnwGRkYiTdtoon3WDMEGMU86dyqrddRleGA3YsZqsbdRB1MIBsVr12gv0fCMA53
7L437kWy5KKho+ZNgYLrxjmukpu/nPyF7Rptb0BxGUvNhKsKlTo8eRLYNpUWw70F
zIwxkEWae1HtG+u2YSO98WlfJTanwL0LCy4nqs31c9FPcq2J7Nq5ndZ3vJkmzk9m
29+q3urYUcCj1Tx8qajVp4soYd3mtVIqveGebx06fsK6vldSw7mYgDDQcGI/aNr5
xOhIlS5CueXckoSHbt63wHKTRmVyQ4js+8bLjxxmX1akaSsgcxho8Bsk2Mtuae3G
Bcvw4z7wgonzEDXvLzPIlW9dIyUsbezYktBxr/SZCYW1J95sYAANULJl4RWwCNCy
WhEGkDji3r1IrE3YNUqkZe/34Lsnm3SfB1SrZB6Yh1zLJ26luRu2SkEstozMYDPv
t4LZwjoGaKMPFLhuXHjBI8ULfpSjpfS2L30BcOMHbvioEUybjsw7oOhhqtVpdU6u
zmhbsPUB+WCCJ56jZUUoTgTssTI7PcVLe3SMLFfMh5OqHH50SpSi/C2lxPeVa1TP
FE0J0/cI2u6VTC0TdohUFfP5N0vZfuqv8Yu+QB7UYGK/KamqeN2aVQvttMO+IraG
ZRD4MNdFhRo/Gw4VC1tA1ZyzH7FTrR3vz/rW1omyXV4YfGcW93wyQMmYMJhaNy2d
Z2OxC5FQ1gYZ1IBvzk+BcMjTLrE9YXp9UJ239DO+KfrgBSiEYe55KnqZ49eWdnvR
/16vBwb9h9nenpm3wnDiLC9zJIRw8t1watl/1QmhxB/IKV4VHTYEADfvfCaol1th
9zV/zyzTV01IqgebUY5UlDPN6aC7fDkx7ExQ0BY6Dh4K1+md20j7I1V0/DmxjJR5
p/tGcOxZ3zrCvuJnek6ID+fFgKxmGieswLXVhEmvIC6XsLFSc3KSrLe8j0KRj9oY
+BO5J+PlnyMxoM2P11HI0yKfgH2h8x8L3HUrlqyrlU876z60W5onXooG6q1ufL+5
Qe8h4KW/suYIG6Pa8JGY95Ssze/GO8xlk5nTaNwLONtNInvIvXy3vJi6PI66ttst
xZKb0UTARphEXi2jObQLnbP0q+S4DxnwhAvx8zR2JHpN+tZM2mKZ72hQR5HblpTF
FV//30qxGN9ZbRTFXGzJg8fFjB3/jdGTMk7dJObKhFP65n981HqCgKaW5YZU4ukI
xdF3a8+ngtrB5E60mHcklOhMa5R2R35z2jIvia5LVCmnWndLSSL81Hzo4xT5Gj/z
fqJS+nMREI1AVj8TamNAcRu+Zt1ZSP3e737DAFjYnrcX65FDVDeCatKP58em4KT/
4uabijJghvxqyngULm1iYobOlq1rz+ZquxvMB+W7LJq6EhaGOT4Q3dKor2RMYFfP
enQz0Spo23ejSSA/IZZVyIdoqYxqHAWeLc5elw305u2TdsE8GjXifMQBdZzWi3TV
oKJJEd8iDAqPQNelQOwiB0tUP+VDHZVtRDucV7ooBeCKAFQbepnPF926Z4mUKi3F
MgqfWuIoKYzmeg3NpkHh9O2iPuoEO8RmisqjzsHraQCdVbceh2assQfnZ5hzSFrH
JPDIu1lTjTjDA+fmOd/I3G7RQIrVP9JX6TpUHwhvOPzLrM7IHLpp5QZ65yd69CqY
i/59zvi3d7noIW4Oc1+5C6VceVDUpJLFmPDofx95cTb6k7Qsy8glf+GCbA5Igl5a
5HziQEeogltGEmbYitY7PJw7qZ4BUIQSBCmxkIWCzVBcLzbXSI16Ctd4Xz7kbPgL
WiaAB9xX1I0eX0tygwul7eFXIL8aSWZBnRRSoTwm+c9uEabpbwx1BsYMYDFNC40a
UYYLClH5+DTXbXhRxQnqAfcVnLcvaG6PntYUQBBAMmNo8c1PyaVWbX77skRTGryW
94CDLJYieqTBAsPWfF7sfZ+ILHI6qFnZVe59KaWj4YYtjAYMGQrR8kYfSgdD6mXM
iVDSkdGsoBQePVaXOKgF5B1ezyZv7ul1hM234V0GlNCMTreYwjAKDF1WXVHcnBpw
E8oI9P0EAK7O8oRJrrFsms+mLjiZrrUDfKuGgfI29nrb71EfRndycFwp2SksaQ56
NLs8AGs0mzkygWmJ2VspdtyiKzH0Sk1QjTvJJ1il8E8KsqvZXgLBNDRym30PbFwM
LW49zS+ZlwlmEB/L9KYiUu7A6oSCI++shIt2QeVvXFCd2Jd53ZzJ+VNoSWaAXSmI
J8r8T7uCCfEJrSfz/icpuFdFoKyvLtwJk/7vD9/ZOvmCFg4aNbd+PkbmsyUachh7
MqQ5MbJLS0gi/nB+oX2k1Xx9CBssyhXYIEHIvA0WL/0WS6bMVKEExgwzw1pf0/yu
gbJlnEwlUEytVfGVsa5Pahx+upESpfd+OQ1cpWv3qlwpVEagSoOn0IaZHYc0aJ7e
/JgiiQTnzlCchBghtdWQvflqf8vARDjEgdHCu5SIHjE5vnZhBE/4fpYx/5Qqepm6
ZyM4WuHyrbV7/55dGRIaqdZOOkB+TVclzO0ibAErYVxsDZJsy8d+L1WtKsB8GEry
75lMtCza/myckdBwcmU9qRsGxMM3Q9plwPxE9MAxIawkp6/8ITcoYOYsaxjsAVW/
EkcBIsolS2tWnOt0/wz8RaykI2PSs2jrFJLEmVaY6ltv7UCHMJaRooR2KiPrX8Wy
dIYK/stvpPD0PlBRwQDA/Pgq6iGsi0YjBk8spP4UjaBTKuHZtYNdwv4T6qDI0eC3
`protect END_PROTECTED
