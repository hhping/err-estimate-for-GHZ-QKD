`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elYwTQftGK9UtgCB5LO/lAZAomk9Hj2DfJXVA3T9Gef8YWv1T73Akvjzf2CTJODw
duP5G/drVVpT++MNlyxTFngU1CCirKfQKzqwRh/R8Ew0y/kGjFOwuT4LOWMJJgk8
ZkGzyyKhp93nMrWJjGQctqht2OJU4Atxre//6hb1feoZ/GDuCB+cKoAq6zqR1oOu
eZpmd1XuWbRaSCOpn6BKE2JbJNgu2EA7oNyuav1YaY8HtkT1manMLfgugShrDIr/
/Y9wcnINybEqMsbp6Wu1ndW4iQXY+FlQ3/y+Xx0zaJcEs3oV9mbHS5J9b+oliIW7
4g5xIWaw1bGhWFspY9BS+HSQnR8t5ZEM+CTTQQpxCdVM89+QuIvi7mfWDjR+I+ZW
gIvtCBAIvnlIcireAV2HUqIe4TScn6V11oV3h/JB27S9XBZUStJ9zTAFUUYOBDnx
Bhke+UNYTjs4cQ2WloJNrYQS7zjGDhDej6gGIozOPSu0VIrwXyzFpxGtGeUrb9di
4OGnhlc+vOoTERwODTJPLdSrKLAM0HLk3/BgsTaauj2fKg7j9K6/4J1zoyJEw3nA
oTmOcfqz+a2qvmmaN9AJ36D2CSyLlz6z9IifGMqEMIHpi1w+CkhfaZ8AwLsEYSZY
`protect END_PROTECTED
