`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8uICNaByf+M+Iy838nzXZhS9aCi/MbQ3nlPZroTUYxX1xVynLZiT2oBhSHmQHRT
ifTv/L1NH+4v1VuetdVkrUSOAjz7X6vZoq/GBQZJ0DItiWAkaMxvuJklui1B5mXH
8KcEqVXodMKcEmapLUCN8ya0OjczOqcEWWgFkytg/HYFvVilje0BpkQe0T22EbUU
S0T3O+n0DfyaQe2mSusJZnbDNzYsM1XmQ51TO9BVDFLLCKeC0rRP8VTOaabPNzer
hOsMRGXdF5upQuvsO6xvXcwBPGx/vi4QYI0HjN6pgB3EEem+Xj6JHOAnPo03e6+D
dq286hjPpDE9UdSBryfO+/UR0YCekxdXsndHLfNmwRNtz4Qmu+EW8Ui/TRbZt8pc
Ylcp2WqT/PR9UJh9bJP/GXd7lIgaj0R0RmIhmKgPvQyB5qz1x3lwmAQSdskHWFKn
1guOmvRaMM/ydOUiK2DSAgv2ljldrd5mtBniuOcXXgi/dJ1cYpFG5VtNQeKN3WEx
Xqhc8+/fvg+tzG77qdMfYgqEt8ansyeiJlVpM8137Ib8C1hQBuY32HYUSnPqggmz
ymXbiY5IO3Es2fXxVRR8nXpfjI2rcV4tmc4HF2qY4bugWTCgtpGyw6hvKzHmUDFu
5r0WsaEVM6mHU1QHPoEnxajG57LTG6n4xUYEqzPLg7Uk8zWbo8hHekRrpAdQ6ALx
rH6OLRlFdmCHsjw23YauWu/Z4X6gnZ297sJSio7t8zY5vriML2Md9AoUeIO1vJda
dbpORwlil48LXajfeKPtcPms1kwtpO7Ef/aveJieezu/NephX6lcCZqVNohfhBT5
ccRsQA7D8DzT/Cciq0MV2EX/h5Wv7cVtfFec38q4oEsesk7KyZO575CRc/qxIqW5
glRfpMp4oF+y1ws0xJbVAUNgyCMlQwk/9PjKkjIG29mpckIA9EDaOjbFk+I2tumv
3oxM2yK25d4aLosuxwYycjmj7DRUwwHn01tm7AGhje2GZ573hMZrjXKDKJyErQF6
5r7+tKSdaEu22HuwPOufDCGo6pOb9moy+yGnjf/nwMCWUC0m8iSBcxN8xcoO5I+m
arls3LnBzo0q8wb1HMThevAd2JZH5DIZUAivQTQRE3wgxM4Ev9x87hqRt4USFAeR
zDILwfmngQxKKlb1bkZfySdDrow9ryhy5PcFD+BREjv00+geulsRZEEmamXgB+fR
MRWouWN0OxiThuiIwpT05DRDdH87BEAn1yGc0Vn7n7A+4Y/cOKNlpODPoPgBncG9
GmBre4xoXDQ9km2A0Fl29TIyEBy9Lhuba0/ZG3qnZXdIhGTQZekSRJ7KIA/Nmt2u
3p3VZI0aGwohrd84jbPseUL0wlcHIBcb0363PVZe8h1aGYgP4PeSDbzljKWpfZ2v
XZJHgQqXeOnKZVKJiRPCSvuyFf8R6GDxqI1e4uo0fDzdea6nDu+eIZcJTHibPn4d
mZnxk184plseU+YfOKxyJbvSW4tia1xAkVaYDlwve3Tju1kVJSR//MMUx6dxfvWg
vXI6EfXhVCC3D1mYpNYRIBjdRajyaNmEu0igRxw09fSG6Lj3d3UbLLlejQPKCLvp
2oH4Ea+Zoq2/V62FHeq1aZUcMNH/pAbTiy3+fJT0/Cegb5Nsi3qUW+gwiPvg9mme
kFU+q1Rnm1lk1ho0bsF+p3Pc+5Dc6AjnMrKaueIlmmO9MpmTYNo7xdzi3O5LcLn8
P1jVPodJ/gmolddLXIfbBA73x54C41z996gkcrcuM94VUtqee6sHToKmWhN71gRX
owtP9N0k+/7yOkvIO4Yny3J8VUNizwLGn6rq2rLVjm9i+echHuqRp1On2K0fxpDu
l5DJuxaSS2oSpUTu3XmpjA==
`protect END_PROTECTED
