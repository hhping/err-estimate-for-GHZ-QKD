`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4iRgIG9rOXx1Fonj42RCgpwJi87CaxW/CmEWc8a0fOgDS0wVYmOxNchtq/2PNsZ
KunXrfn0YgGE2j/qs6bkPvjv+X+rxQVSyPtqsnHz4d5x+HuKrq8pEe4mhXRwD91e
S2/uutBn0ZIUhW33zHXZti5rQqHfIJt2hTJlYLRRsA1zE38OzpuEY6FOJ78g6uPm
/sShV2XCkiCd7LsQZjiqjgRux3orp8eH7GOnBuodafjsk45WFGsWXWfDFItTvERc
/SlW491atp+d6xZMM1fRy6HbZEBvSWtpaZWVD9IBYwqgDEld3PYtYkmFBWVw9087
wDdoAF+H9ICuOD2BnHaNm2TfbN6PhcknRebqLvhhAgNqlfdMediMEt/mo+pe0N2N
8QN07E+PUAuqV56FLBPyflTnBH1Dp4R61cK0GvUpBa5t1qfkIL5/lmhAMjL/Zcnr
vrQEf7NOO8CM14WQDyiVU3kfzOx9M2aFFENkll5pp3L3WCjaRSYD78Zq/PzPm8I1
eWSvmKS7C1dfZ3MQKoyo3vEx/M49OtwXGQfSFwIB66XpMwmwSivpvPHBtUyjamfC
nmm31sO9HYE6oEBoGTCjspAcW4zfGc/3vmMVTBi7EDw7QJiQBJ7hsFGr1qyL1OaB
U4j3LN8IrFFywuS0bX1cwoJbCNo2gw0BDkniWD4BeKYLXpVQIHYjFZbg44hERSk/
poQILnPpW/1CMiiy7JAymdp2nxy5KBvc5bsXCGFjqzdRsVU81iEoFvXKCHnLpGFe
pfm8kHC0UgwKQlYFvu/NssAwP5paz1io2pWn7YCGboR/16qgagrJzfNU70eco/A4
QYsqAECZ9+233Fu3YPpXmPEpVynaTuRwuoO0viA6ZlVNFJmntDh0Su7Nv0EHGUHe
f2vccdGR49oQv8MyMm6YeCkSn3x6sZUTWUATr/RQUJtGzNhaT09cNXmlMyjkbmBH
rJoDYwCnZEFL3qd5JOE4hw==
`protect END_PROTECTED
