`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1KHw4aiJh7FTWyBuNkNXj0enXryrL4APFC0VhCtFJOfzCXHXGX/BpH+kk2A0EwR
rpLHK331CzMwQfxDU0pAj5WoJmzpKnh99n8SbDnVaZx+prfKQJ0xv7rf1uyFZdU+
47ybpiHZsfnEfizobjhD0zikC4xRRklo0gu9wchZ1C61cEBVG3vvFJoEDa3fJS96
fY7K/u11NOiluSJutl4YtX08CnzaGaHEjQmcL0hKVQ+UxWIKGDXMRLkTyet9HiiA
tFbZGHShl1hgEJ3r/pk6kl5kqV3hPNmqIh+jmqjA1gL9in5sHJ7CGRmRqBijLcvX
uhmC6hSJIxwDcwiUUw8qZH4jL/Wa3K/kOzbpzc7CZApVZgKqboZFT+L0DxdwTGsp
shLtKx5S7plGOJV3RtMqkgAvVAf/odvK4p8QvtFyVvWHaRT/GKEfPskKC0bQpCqm
qPgGBe897C0YdGSaHT9YcWoSrV3rSGyqeBhGQHkJ3P1PU4WNwoHCUCL9yFWWdgD7
WpaZmmQI7jC+ZJDu4LZ26BchxbU+yzZgJPYkhzqRT42lPCUW86JqVd/Dnsu4dV1L
NelPIDzHueL4rK3DaFxuXKtxP+yyAzsr2kbuSsaqJ9H0LySk6iNcydEdntVcH7xe
dbXMsm2fSKNDoE2OBTPn1A==
`protect END_PROTECTED
