`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uvAl/10iU5Q0cVlW7EJxLWSjk5kQv+flWRzIBas1fYGRTOfWUaM0t8CXBMswFQpJ
2YqDVHvRFRkVDVRq0Kz3uivrPTtUSrTiazxGtmOxj5JguCltrDf0VacB2PU1o1S0
0pCAmEdgt6dDjh1UFxWepMXeuNaS9GUPQK0XGPrQ0tfCFeIlcnxUu+16dn9wzJ8a
UsB2cq+h1gHRbPXnusoVvYYSq+XSYpSGGHYROzqXA0tlew3JFPua5p4+4TIkrYnJ
dMbD9NpVTlccVAXE4BLS7KWEorSvYnS/3TW0BQpGpJQuxgLIBqQ8OpNeHxPK+DcF
6SxGkF36tdltpZ0lc7zWQpl+2qFYKjjVeOT6ytxWXAYOMAb5FyqdDxx2p8ZTiNLW
vrtgWaL8HSb6+FdewLcWYrXAcFiOSWqC/dTZ5LIJ3fQh3HzPklriZKNra/fRoIYS
8CiWHIZZg6J0Ge1axOPLdWBP04PLTbxlAvMhCo/ry0fJio49kZfPgSvOQjraa50N
YKzm3kRNBn5GFg2Ul2KHucIIzZNi68C+iW4mqAIgF9EYURLnWdpDd3b0eYbMLD0B
`protect END_PROTECTED
