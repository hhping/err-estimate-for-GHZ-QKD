`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdfZAdJE5p+kKkrxwEIwvYvaSk5wafVUt/QRXgxKsEYGt7r1uteLmKb4Sz4FKVBu
7HN4rw3eMJQE3ph5h+mNtgz99Kw9HLqWC8oiWZI+b8hx4S3xBGabqCZpsvBF0Ojr
5kOG3Q49Vydjv7TmTUu9kRejlq+YfAoJ2RCrYFJ+webHxhGcGojDBdErAvdexKb6
+zm1g18YmH+3flAJAQBCkzT74C0ZUcCCkIfLuX86rOnwWZFpmVuWJgC8bodRLbE1
GTDWexikR5S59YyyjH9QNGJtxi/JUvOYLpCFF5kx2OYT4d0wzKt+dHf/A8MITGPm
SseRca4z+gSXM1PPTpFPMVmpsPF9QBotloBvARwmRXyVHtsaE4YkCWHfMj0LDyX4
B1+v03JNmzY+ka+ACPVn1BzJCYNcsyStkNLsJyxDXpbyl/FQoHSMNAxzIKKuSCtM
umaQ2EJnTgXePrraz8dvtT65rlidT7eTgExwWf/QKoppN13bMHM4mbebmcp2SUSQ
GYaN8ywfGBHX0GM1Zv6ekE7HljQJyPIEH4qhED0w8x0Z9bB8A+lTY5cYxgcPfKbx
w2SbCZXXN6mLfaTu6jvOWldZpGjdNxFd0QgOQbIHEk6pfimP3yCtMrxSKBznxh2m
jlcLK2L6wMDZbbKCCKtOZg89tj73dfXsv2s7twOQMgrXcijfAcjOi1zL2Nge7g0h
/j61e1kYBhYxQE+gAffkS+6+gXnxwMFwuPhEDrHAaCdSJXxOEs8v3+yTi0EuaBqC
CI/apNiZO3K9ygL4dh/FJEZT4AXEKIlwFip5ZOnGXyXlkXRgUFS9XSag8roM783x
BHKZaxdondM8eHwtgjmq670+/cLmOsRosbshmu2iWcxmlXvnH/UycfNDXptly73V
9yPOrApKtaILP+4ioaePXALOX9CTaJM9pQwU5Ll3yzJhGMRhA+Ab4TyvjSCvG05j
63k6MzVd6ImpNAdZHrOAT3He9doClNgF6IFXfTx2K5vDP31Z7MSBWiML6KGzWecA
gA6hkkHtStgjtO9Jv1pMmJ37AW58nciRRHYha8EIuD1i4Mku8HSm2KSdhvKG6WqM
AmGDTyqRMifQS+1kNPtHaoxusBzGJis6K5/LCRdPuYqbi6V38WpoOuhfiNKgsiUw
8y9lg4wezpCHKZPaOocyoWmrPT1PNwDQM/uJJWlYFCLJ1LzSm2WQWZmgSkPtOIcO
xUPFK9o0amWMwP9pzMXb+ZsLpEfzyic/E5nPjp72rcLbOlTe+vkWUBaBsLGaO9rH
Q3x6W32OMDrb/Ea1YXOX390qQveElSCvt2rgyXUfMhBBojoNc18iOmAxHZd7MIPx
EgHpKZbokLkGibNA39wKsB3BcZwtDyhJ77FSXQoC5LjcURLSyO7Dp01/Arl/Hike
oHFi83IhBDW1xdHG5foGsXnqFjejpwRamMTCttQB3SvyW1tX4F8LGGwCAXYTmNvT
/uDcyk0Pnlrsq6/kO7n9mfh3BhSb24IeXo7BjlHykZpAEzTyMvvFbCsxbBbqE4IM
HRfM7Bz1aRdCDN0FirfA3fWTI3v9leVTGVmV7K60WtRtvAmYMKwAd6R6roAWBL1K
UXP/P9zjUBANfYyINmxVF0rrvORhJ17H93Kijwb2dvQDIeArXsao68mwVEbD2t4S
V9LzMEqnFTUQKxmugI+Fv1nHnSB01ZiwrWK3Le3BnKGuiejJEQM01y9ceyd7boNg
qh+FAnDZkShwZw2armLnEmEJytIZ/LmvFgSdbn9FpI7nJh+MUa+liFmXMaH/7KV/
Dw8fsA/88RAF4SiRIrl22sjV+UYgl/+xhatnxXrmiv5G4PnniT4TR+bZ4XPP/6nP
66EWaNNWl2XTX6XV7+A0NTzgZof0QoAITc9PLzkOEehYsHrP0RP4eKFY3jqaLetl
Ot+bDCFVieb39NHkpdcy+I8U0s/ZydquVcJTmriMK8VAHQSURTWQxnFPwaMR9tyf
bwkgvkG9V4aoVCpK3HacVuvWfnem066CU4fgI5fagg6sGC0bUU+eNlg9v1BCyP91
hsPR0WbHzXjn/k3cz0iN9iXbznSBB+5nGDAmr47fvu1TK62G/BRQfM+K2qOPkfGD
Gjuq7gUrANqGYdEB6zEpfyGCHNKoiGlMdO9GkKZSDyQvhUd+FvmbybIKxL9oO6yl
37V4bNAVYrittjkk1d62OCWThUyQMwpmWAhhc0VZONzVtKPCXyWnx89gALlynmm+
tG6IxkiFzfWKOlH9AisuRejbqBLg+DGlBhFIUOZzi0OZHYHKVCZcrAmXZCA9kRJK
X2NQW4xdEszTMnZ5IovOjY+gu08M8Dh8fudxh2CnmH+j8ZDY0iYRARe11NfOkc0R
Okenl/ZoXeSjZWMQubfg+t4EJjkE5ioq9X9EC5kSXjs8XoAxF1/RS7OLA7lqWLZy
85ZCEwCqNu9Orq9SOJK9Uo+jWaIMTMXDGjgEFoSkF3k75SKXyh7fGTgqh+Q7vrDw
XTusJEpnodfniXBFsHwNCgtvWagkI11oYkrtgBX8oS9D6Cn8+DG2hEDyqTIkJEJ+
hsgWRY9yzvzbmhCEDykCr9xtYmG5IH/S1nyL6FC1vSZgAwSK88pIRIPBkEWFIdzv
HrTqrz3AUGslF4m1Xcztu3nbdEIUZzZnSGn9jHiasOXaG2N72guMeWDxrXsLKGSL
96JFcvF72jnDJR8Fynpn61g8NLwjaHbnAPlB3gOq0sxtleF9mXtk8p0jbUNYWmlz
k+tUT7mNgqmv3alFkKv66rR5PZXpsy6HtG3wDtbM+YwGswHO0V3nFbh2KTCpmY+g
OjFatAdu/FXjUGkqS0khFPVtcNVi/+aTvtRCbsLAFtCd6CD0ce3VhrpRFK+FzTuz
/7HzoV1kjX7JvTbj7BRy+e+vyCUqd7xz/rrLIyMUUcrz8XWul1boPKoa/HYna9Mv
jD0HUChnWyPqO4zKdIWqPU//jlsx4+wF2D/MCFZJkIh0bkOWnI4Qk5G43BePXn5Q
J/5mYQQoEuBqrh6WBySIC1s0jjf//5Ol8/n+JpFQywJ4EQqc3LAc8JmoFQy3MgkN
X8oHth/era5lCTFQuFy3hYuJ5ondPP9TNisKjeH4MAI8BNPItDm4Bpd1pFYfsyUg
wRPp/k6zCSSBaiJ+jHq8cIS5rQEyNAtWcKX8ZIzTdWPvk//EJP/68pBOv/25qLEF
j2YSqBDJVgDGOiRNkzW6cIeTIFUGLDRce1vMmwAX+8NXLeb2O4MTCzEQtQhuDljs
Ilp2c7i0F8dk181HBBHCdREuIeCWOK1eLBt/M4zYLd3zDNXNPXGkp/AenKnBwEWm
tQzHeMKT41gcziNY1RrAd3UGn3wyhhxga/WdatQWkpL5d3oiIHUSHU4Fb8d+GgBG
Iy4js8mhjkp/4AfEtBaUw0jeAjKRJa0nT44iSAfa1wxPcQzSCwi/3qn5Uu98Gckc
y1r/Do1bEMx6wesYi41Eyphygl2SMypnyarC6YEDNvnSNCERrjVjXFiOYpXAAbFX
gT9myVrUl0dRhFS4S8pIitV+IufR862bnrJOO5TOZHblSe4eJgejFEnn5YhUkMRo
NcU9bvoMnjc3oqWtKrGynjE9vUVeZxr/Hxp5uagLJI6iOCZyQQNOFE8qh0oNyLET
bMDArpPB5xVIQ18jWYhN2KpbcD03w5dflJhR6GYwengntbbMJ/by19qlHZ5nMDcv
fM+WhZjFczAB3c0qGticsQLK61/ziqEOXD4nev9W+3B3CVI7C5UwyEtaCJcDVvIr
7hrBKS1q7RCSwYYy38e9yPU00Ys0c80faNMXRL4gLyJ5rsELQ+WpgdYQCUC0wZ5a
VNqSDWSioumiREr0dVXfpWyoZPgQa/NondGE+P1Q8aj+2O1fEnaWa2LfJ10vc7vk
AzrxbdYkfnTwKiM28DO08iMAI8S31NxFRUJt4z0Klq4ZBecUpvRPt6hn1UENW9j0
H3VrCUNzKl/R4AMFvYpECIEoCwXOHHX4i/QE2q9Y5uWNX/3n+8KfAOfhkay36oci
7bWYGMwyXfRtbz6FfOYrwZd4JiREiZZYZNMNEBE2V4snwFME0pHwEwpKxJmqTsdd
xO0NTnclfDbqqJucgCq4r4ColR3Wf7A7Z9yZ95gii7TKs1RScPkBHwj4Yp4Ee+/V
fzFnm+htQ44uDdAWy5WlEmjwYavi8j6XUZCLDbl5f7qrzDpY/RrTbd8lUD8Dc2PA
Y98iDFJSf5YBBx4poMRxGsydmtboYmaKNN/zelbALfagWOk5rJvVvQ5nwMgoPihR
BY5aWYNQiN0z63JsVVpYIS2WacQ6DPXIHtvPJ9QfT0z8IyWWBPveK1REsgdjlYPx
3vmLp28qdirElMUPLiJ911Q6oIqij3J/PIyRGwZx7yg38uSoaI+niGlEzRtKG2o3
wizWqwQkJbZsyA+KZjI9YO1LlYHIl1jr2+8DZdzSfUeMGK7Pwpn9FGYQ8/0hl6a9
wZVBymPFrBBNl+hD37NhAiyCYAIOxrRX7i5/98eDWPh8DphTberh89gxCQT8d84V
C3uM6Q7qieEyTwV7Q8agP839TujwnPzoxWZA8NJ3HvbmR2FOl77fK6lJv+SUYvxK
1yfzS45xq8hVvjv3qQj86Uw/+tDXrLd86PIDKxm5cZFUhVvjSu4hgyPQAYL865E/
nNOuON7VEmZsARz+lWces4zAlB4ntIi/VE8f6dEVwL8ygF6V0FzcGIKgs+lq70nT
p+ICFASynoqWn508HArGLx/f6JR1PpLyNwyQglh2sPNX40c+Z7DJV1ybJBTTnLbS
+htxCcsZQgKv5iTftO4Ys2N4G42n7l5+SAg06CeYCwtoO5Da6MxW3PDw4Y5YO7wB
+AOm/68/nzsj0PxmH8Yyr867x3fkRnhPUc01hyuTOUkxSE3IGMRLyzRRaU0sMRl9
1qAtpfuyz5yUS3XjMmd9Uxzr7Csb9zwhMaphXnR77Dhmq1CU/fRqwXXQDUVcfzIA
rdOQgn0PebyIGiMFtg/ol7k86tT9pbY4fb1sLFMtslrOiklErdACdAYpPmzeS28E
nOn/VwVb4XUyph31M+Vp+hd/Kcc2nLzyCaXx1Bjxw7bk8zee9nDmZsv9X+pUopjN
lFEE68NvWkZPR7YlZrSyVdvK+5Hz1mCT027RoCRbQqaJbzBCGvWjdI3hhl34Q9ez
Icis305WIEL5JksLx67yviYSEowzInOMPjGGmlzE6u6u4PV5R8cUDmVLfa+hInHY
vhKTvbQ8uLzXjmsHDCweQx3N5/AGaR0/JQuSv02KGP8UHsL6SPhvtRzKuyUiK5qz
2j2Zbuu+maLgSuo2XKf5Toeo6Y6hNuwidp17F5jdJ8yMcjigdHqxg4rbGfBW3WqL
EsFDgjcn83RC/n6JvF4eIXKpMBKUtzNm0kKz9Yu+XBqSNCnHwewJkZipM2DLMQGc
FDmxKKNIrg21Zs+IO4YiA5K7uX+G6uIq4bqo3UcTjs7YtTDFpG929rHryqYhS79+
+eHxj/M9XV67T/70Acbq0yE310JaDlBKLXg3wG5jndI16/RQdFJgP8H8EUQ3XvWb
py58iYXZkzLeRyWM2AqpM1g8mCD87arx2bgPLR3wjUv5AzwRUJv20hIkVNtoEDV4
jtEFUS52RELiKCbAMTS+DBRCvp93u+FsSk0PbMbtBNMH9Rs7WJAqzeS4bpgjhjjb
7zkkzDgO6TkZtHqWpJt0YS2tGIfQKNfaS7XwAS1JNFSIal9G6NyuUrvqHSJSyJER
Chqd4oRHhHgnKS4S/fkaTvoaXP75+2k0D7cVpo1lBEz1H8mQ5jSlhIbXCexpFIIe
Qcu02LKEh0K4Y4KPR/gwi896Py9IoJq5tzOcCFnL288eY2dwhM9NhKp8z2ojiWLy
4VmugH88FCnVxqQztoA4ir/j9EVNNSmQBZJ6stKnU0fXs3lqBmn2fH3PIp93Y20E
ZuOyaIjXUQLqUQqQ/Bco2oT2Fn/6kITYI6uIlOxWIPEO7AzRDqzwdjgZAQ//jIBD
RiwMvlpD+X44Dx5p74sHb9y6cEiKmS2QoJajoD/EsIljkX3ZR1+Va97R9WAfV93z
fXdrkeT8Hs/W3Kg4VIusuvzV6UsbiDDxa63mpRGNgetwoZLz20baBqCLNPGIvu2B
c+0omVSkAlMGXZMaisCgI7R9sqnPPw+0Up8IeMUW/lijvZ5+z3Cx3ZCwkvEGNVNz
LAbz45qjpP/6rJDOudp3eYBta0N2hR9iU0FLNOdknFNqx8ZZoaUvvVUVhgWPnqth
1+x25+4YGFm5Qix6F8aIIKe9bOSRZdHNTCKv06rsY2XYL5jrDq026Mo6cilLiif4
9n9TjsZjR3u36vaCKYPB2t9wSxUTnjeuqYcj5FSXbVtJIGiZxG6k1pYGgPZZ8EHl
AWCWjuQt5eeYz02+aQGffPhl4+8DmLefdAq+qRxJGvaMAylvzD42JSVHJHIYtvIu
AVpBKVzcxN/b6VEfW3VJlvnAzGZNmHE5RQHXfHIWspG+uIvyuU9LFPPMPl6irZkz
hBdZnoBovRjDUmac5GydIgFKAYOPUi/e/UvNoYT4aw69WviOzBhWp5y2QbQ8TdTr
grPDXN+7ZQjP8Zv6RAqR/DPWzFNWpDYbfuChRTE5Jvi7iaiXPZe7SBujn7eh2L1H
o5PRrIHh9S5m4CAXTwoR0L31jkYcGTul1BA2GAp/BE/esfJQOCmnqfmP/HEet2pn
btEfuGerxbs/PnK76TYWc+/q5VBT3dhB7tXep8c4kE8H4p6XKAuvFVfwxYXJD06X
xOl5eTe9ctYYdTyleaa2AvyBJK5ekxJYXIUpzekQlc1IJy71w2MyGJEpCTwLrtjP
r+RzBA1go/CVUfOTiOrW9rXXFtbyAuMBBHsilrgH2q5v8ChGLgHTkBX9EevByxYq
4XCmNYd6dIvFSHoHQmoTtQVCVEjFnp7hweUXZ3B8+YZLgbIGG2/iVDCXRnE4xtl7
EGV+0Lf/ZJ0yAqXsG9TR/fwDAeqUIcA8w9w8O8ewz39D0b+MG3cTutGwd5+yncL6
wt/RMaDGXxUMTZskKo2DJmnLVybU1tM5y4790QDMZ5A+/lRLh9VCpYsxbZED9iNd
PIB3avZfyytijzQOcz+vSbRPJCHa2ODjJx6+CCm/G55o2vU1qXcIyI5ZBRLVC9LE
sGbNB8pSp+bNt+0uP7/udojHgB59Z3ar2th9CpaIZeg=
`protect END_PROTECTED
