`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0chfIoinJo7ptE9Vw10Ejf47E7GmHN+k35l1INM2SIqUyJQoG8qjZm94uCrEt6x
w9V9PFlqrR5tgGE95eCD7KY10sDa/Q6UNIAmsCgrR+KRVz1N9PVhiIc/w3+zOC3+
BV+dcGaAYTJvNRzcs3wIQFoZA614mbzMQUUfNVnnCO6LDwBJS9t8LjuA/onWMDKN
FEx6/DAkbBQbNEOSVziiFYdr2b0AGW6IiykHan8zm6BO5+xRWGPzvpzDBqsAWUjm
uSpC9TwdQiw7NftnvJIMk6XlFw7Jz5hj5HsOPY8xexfDX6dLVIvVvsThacXi3WT2
5QqmQy0KatwZ3I7PhbrhGFTHe3h777F5YsRu0BjUTct0vtVrAMbV+YiMIT0ODPo0
vKb21NO+yGOgUgFj2AI9WEJ9cGuiXawu/vTAF+eB/TDbtVUxdAuniAjBvQzgmb4k
cn5WN2sveCJMGuz57tkhZiaLzUJgYk7tkCt3lnxae3Ia6amrAx1b3z+lSPznw6Mr
8Kq8lZ+fR1sOdefejAQO+5JkQ0xw4kjn8a7N5d1e88hKzeLgJ1bSlyT1o7SRh6vI
VgDz14kZrIjFRsJYB7EFt6Fz5+7l3tyfHKA7noNXoYa3nN/4cQMqdbvrKh1+dtox
F+t8i1V0zDzdQTWrEpfG9L0cEgbh5MO//q+8/BJec8cYgzjufxqJ9HocRW2alJSq
Z8oYfT1fmAr5Q/F8rLjc6WQdvi9lMjszEp1KnPg3+UPW8PHHbHipoH2ArpmRmWbI
rQQJQL6BJn9FXG//Gyl8tGP+FP2dImi7ALqfPOfQ4b6EY5okoRrK14KkdpL8Sj7b
Do5r4sC4CKdB3jeDSGu8p7G0KMoyt4m2iMEqSdq0N8zpU8/uNKq1flgfYpBlfAUo
jVrAv87TPWwrvNhMRnSrk9G+YQR/6DCYhclt2k3d6TC+P93SVJzut6sG1AF5pYR8
OVY9o8bEkSBmffW24mBbCg6vwpmGYMfjjgW0UMkqdOQX7cqUNXJ+HLqgPc53EuPx
k39pwuCAUMYFvsaI5LWLuApYStBXcaX5QKBQ3HIyzUIRDO8pyQGKb/rktBmRPgc9
MxgslI9nKPx5QQE67aQIcBbwYDJfqpgZ8lAtXCaaxjCS1FCDXT/+Ul2LvkhVgzcg
h2KeZMYGvrcoyuQ+l7179ZhRR17sIAq1mFE4FXq2lRfrV1XN/zmWOqtS3MXdC4qp
NIu9Lrpv4kgSwP22Z9EAuN8Gn0j9YG99XtXsixtzg7a6Rf37qpRgHwaR5JbdAGSl
ISu2WPPk0Wj34mpcXQvmPY0nb3RqopmSZbxCRqUVamXzdfIdijRwpKe0WOYbLIKg
o6ZF/4HnNzJ5SK8CUkPxJEWD4Ixmyli2bQu/5TbAUK/IN13ovxeJxGareqK2iGLe
X0DTqzofGp0/iE5gr8VqmTK8jeNmFfNY9rc2u0UP9bS5x5cChCLOHYcUMUv4YNy3
2z+bOSGCi+mCZWYn6Um8vzsUCEMBF8Z3O0todXU1ioMOMzvBdr2ipzCif6eakQmd
bBHkkPE/tI4JhFMAvGL2TuffIz6wGDjlgpuwNAQG+schDvA3cJicWLn8fLnWUn1K
uL8Zz1h11qdm3Cj/RhpNxQT8FSuEzQX3oqsTE4t6TYLnuk2yOHSjjI3HcB2DeoCs
2e1XUoUxrigmo5/uEQ51doqH2dgDl/JIH3DbbrPzCbJWzVerEI5st6j7bBT/ILVg
36npixPXQNrXq25HxpEnAGRGvu2uXz20Tx0GZfghOcnNjww4TInSYziOnOcx/erd
cVnrchEgEXL8gyxNnoFdUyLw51SekzCgoK45hxQUu15RAEujhWbv50YmuXwBGENL
nGfl5CZRmFG+VqDW6cwTy8YGWeDnSxBNjCtv2HqaQy4Ym3uJHF3a/wJMNSVR2Ny8
jVBbvWoDl+Byi7+np3AvwjHR6Vdj9V338albLPWOUJ41FOslvpWZSVx7pK5xWPa3
yx/uplHDeOfai0Sr0bJ/wIxuBlPsq+nuIEU0cfwoyQHSbYZ/huU6IW/dUWgHD0/t
sCwn0dnZ0vn0Kd16iWvJWOET/y5mcnpZjvwhsjAYcmvVI9LFTAvSxxZDhhOW5CM1
ikZ77SbJuRNlVbNqg8fICB1ZcKGjVk4IyWPoNZCd+bWHUCs6jFhY38Isv+8PTbxB
7RrzBlL26iisFOf9JuoSd5UF9MG0pC+4sBLk6AcWBJKWGtbREpkwm1lfaZdOidfm
SrEB4nO0WFySgX8ZvyMegPUOc97Fz0Nuoa2hkaXOgB4VrowEoCZSeIo6D3n8UIcJ
O7LotqNKSGsu7d0AXI3tpWzP8/zZLV/Lka0ucI/EbNCPnntcqq7Mr3cuuT0oIaHb
8R/1RrJMEDM3hSiJJXmFISBfG1RCbiXz9REV+ZiNICks2xSciOLkZN4aZS4if04m
rYQRk4x/Cc4pKdsaVy89PJ5zANTc1CGnuxLxTolqMSI89fnib4egq765mjJTdQTi
KKwJ75MH9qjXG7iQe7w2RGbTWBVaKiOVXNdSDagDX5oDjSCY/62CzJMkWiHw0YtX
gzoBdPilwbVvvMlNU4xtezJ9K+BgzCsulMwc81pVKci47BI0ycsO1iy/kaZmwUGW
FiZ4WxfRM6We6A/oUbwuIFp6594g0xLnZPXw4c7+g1jDCqP6w/ANEViSyAPdejwo
s8uEpTD77PoRzQneim923+IKANgdsg3dKqD8DRfQC7nbMbv4UJw53IRqNnr+rswz
bDlwiDL2gf1fjGWoXeyC7OXNt4D6Loo/DwEe4zLUMAkPoedI5R0HHCvwlsr4A0LD
nTkiW3w2u2HGvc7gEz68Z7lYH7/P/eZy9671ED06mrQUQ2TtXPZs9UIzcqoHM1e6
jmCiE77hcWQL2xwQFmd8Uv60q6ovfgwsd6kX4+d4f1/QB2537rZgu5D0ijULz9UJ
+HVjzGXM3Vf9nO6uuh4y3ij2+pTkQehrk8SisVF7fHCy8+8otXZczOJAOCEk1u4T
gg9SwTUNzbNHeRS/aJTvvKkd5iLI4UzUQseytzvDqlFbHK7R2CRqgz1Sft8lJ+tO
DkHJo01oSnJSP9Yg05dRGw==
`protect END_PROTECTED
