`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ooKSq9s5DbWI0+LxMSQtI8uTuzzbYUNVRfYiZas4zLf2LcSb+3AW4ACczFjypMu
Yf/Em/dWYRzonBKiM+5oYqPtoY8UnutzIOgxZFFgRbbhfLWQnIolQyNwWNWiU7ke
8vItoIfEkP4+NgUxQZ1W/4a/vAtbFgwHRYoKnc71f/9YmnhIfc62WIyBlI8p+K0V
doeTyLOGdMoTRQyW0TCFQAm7ZMF7om4Q+w6T9dBaJ2Ngo7TGS84TbLhFl9Vythoz
xxu5oUeAzpY/FXDEJg97gSGWOJtHBFtYC8+uTDYFkNzvgLSuGlhYuhiisCUtNnPE
3oO2kslkC7FM3j9X0uDsVUb/bSHvPmlrx+KwWYwqiny2aRsWoOLq8PyXZ2cJnMI6
KKfniH3hqdgUSjCrYYbkvzKMKbt6j+mPHVunuD/6jPZEUKxaDIRbnlU/wimVmSPQ
ycYNBHadc1EWqAdszb51uw==
`protect END_PROTECTED
