`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m5rBC1vDa4bYkpZZvw3Nc4ksJtdiqGX6DaFovb1tTspiMoUiKu3SsKzjH8F0elEE
hJC4eTY4ofKJm62fzLl0XObErUDNR92epfgydj3UruJb6PyeWrGEt0g/67Wlbp4N
KSPCun7cgSEJz+IKuUJ3K9a2cFT+9SGDloO0NeWasBOOMwXDsqCVTe64hDFx2WDA
m7XMDi+vWrtf4SoSdRc+vaVKKzRKctzoEB3PifVX6p4lxTmwwGAIf2dm5FuZdL6r
Io5voOrvOKQmbVfaOftuLROnZPh7KEjiJHzPmDPk24MjpweXkZufirrtsrbcw8Un
edvaqK6dN/2tjxLAa/UmEk0N3eAWUpsKfBUZTxAQLJtQT2PvfNAap9/mAqGn8MaX
mfjgROiazfv0wPVCJjecrGPN4+ZJ6g4EeD3o1D1+4qm5wkTdfdBPilvJQ05fNtRN
jDkXbbn9gYLmtAg116gmxG1/X6FWWMKR+5/z7rh1pi98Hjfd5yKPwylx6+PItJXl
oY+NMzJ7lbiQbXrYw5KVh9gT/h+CsbKPvcWX1k2bh6oE6wWpLAJ7PO/y77uIhqCE
jx2UxgaFjF3QgDN9FDWDDfqcr9oRJ1sr3UWC6cC/jKMNK5JzJlKLQ7EFa14EnDbf
NHnyv3OkH0itFmxEKnGsdIPN8bFMD1m9OqsUatOdQzKEUV6jBMLBH1VCCyLyMlXX
VwLEXl3JbtJHcw70f3kA4jbGfppQ8an3KHUfiksCzKnrLtrRFXUA78zsSXAZ+soY
BKMoWsCn5x85Jt2Maf6Zdi8txdhTBtFnYxTgMDeTe4yJqd/8KP+oFrH7QlweApxP
KdS+rWB4NNU77hoc5ycdR1QMS6bNEzcAYhALGaYK3fIhqAxb+ZYhEtjnQ7zmXmoP
O9citZJlIzM3XUFwzycl/cHW0vYWPaHyXCcpuDN1XkLLQR+tZSsl60mtSItNAXsA
gJYn/0fwuH5Wd+rRqrKzaMfaQoZ1oMrs7gUf0izZExxaQvQxT1oMR5VIcug8RKl1
0lB3vk/SAJ9K/pHP+iKXIth4hfnKC0wFnmL5CWocY6u5veG1SGtdLQoRl6WUjB2y
VygbOboWMM3tWs4s3fPnHVpwtSUJwYP4a5Ej1qDOfNeOrxQDZRGoif1Q3v+7DDYS
`protect END_PROTECTED
