`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dea/8PkG99QqJXJAjI3qPgZ3b+bC4txeM/jMZjpVC4MhYEwmNuRamcVyaXTEIh0J
GC5Ea3Js+wM0IcGuk28jmJQ89J0ulx2egBYfYAl/GNshrjsrgbhoQDEplOKXR3yI
9dE7nEsho9KgZzqSdMouu2XaCPgXhAJKCygXHZNX2D84AHlTSPM3IbHjnF/uYuYM
Sfc94I9LDnk2UCwKdHMZJqff6rT9mtLkgWOvbd1FnB5p7YwX6/GzOrBSBWHpAy/N
eDZOTJs8E+Eni2XmpU1tl1+U94pweGQsP38KmwZ2CGvlYXlR5+EzJvwnQY38DcvT
F9j8Kf/U3JLzHlLjHa49++ghTtsLBEehaw0RTvhx/H5NVoKOnakZJczbRF8G9I2e
`protect END_PROTECTED
