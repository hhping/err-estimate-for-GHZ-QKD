`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4vTOhxnZvYsI9iZgHBtXb90E8WhBaYFCnpKg1OBLzr3fearhHWVHszBy3Pqq11F
27AYu6WRqF3DYppBgVA7sqUZzF4SViP/DE1XeNWafaGXiZ1LZSd9rpjRDEOif3+C
cHMnP+IcZw26Fq39g55LTiBd/J2VufUSNKQTLRWAlLEZNniPKFmmBAPkA+xNTd8o
UpCb/vHnKpVicNdCUtV5R0GQc3IRvtwjZlJJ1PR3MNz27kzL/HEX/M0DIRu4Q1Oi
TgppPLPl4Awbq18nOWkC0CEIxMU8ViZmQTPRndQB1VFXzKuRPV2H+9oxTE5dDWsC
T38ObQ/dyVMIGfAUW43t1wrfXDwneNxRWoTH29+e/P5aWGMVcOKARAHHk7qwZgJb
QqiVd6gb9lygrT5oNe7sIrq3+BL7BfZf4gQw7srAgcCoU9oxlmqApOFzYlciPrQJ
a9MlaSGCxtpL/19kieUuck+Zf87fpD6DiGjpesiCA6sNpTif5Ryf5prvaKAAsRN/
J1H3+TpCVPyVvczElvu9s1vE7t+IgmmJKTWlGsztBx3n8+ixqaAp6ENmx95RQNuR
R/CXc7xCUgeMtDzMsXhAS8sXAQIJCeMnv7kfEygv4L1hj0WENJ1nklhCS3fA62lu
`protect END_PROTECTED
