`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSW+t0uQgaXlI1woTbVtV5FJe2NzUlTQZ3JEZO8Iw4lUqGUUPnI6joyTEqaZbBze
oO7fQPkhU3e+mO64EkHeUk8z6pAfA7nkyg4P6VwWH6tj7cheXQe7yW7brJXEfcqH
jfdnL8xFkMRtpmUvKNhkD3vM4ZfGvelZLqmanjxX1h29SJIi4m4lqdtyKP4cAJqQ
53jjvB/aMZAQ5OykoQMjrthh55gXQ7Lqd/v01ke0qTxHxv//n/QmX5vwXmb7jbhV
6cCB1ZWpMnbhf5C4TweUl/5c+bzTOp9kFjJfzZXbSkf8nXdipD8uLGRKkhZ6uC08
/LCSyUiQFotMi0ZsXLricTFk7VJLbnO2CvT8ggA/OQtkgRHIJLtr0WzP0fBzBt20
7/jwvX6bdOSasQXW+s06SdsPnSOBX4y5TbRl1vJMKHxdvFWp3Plz9w2PCgZi1Edk
Zi+gdtXnGA9FTjfcVoZxDzNB8+tJSI3jinnQksr3BdNZUfO0qrJzThv8k1tdob2z
JjtrV4W3HHhuqlaVcbKj7ZY53TAuhivAA5IM6rILWEngKkcpZl6+QftjqwffBkYi
0UmLEqGQYIwcO2/SUIIWwaSw+Lzk62b/K/yah46t6QqfFPhHHAmhmOm8/YSHLcsm
I62wcw2P18aDucFGAOgiLJ1ktANblC147UYoyVYx90Dx0n0Pimr/+C74Ii4XMzji
p7fbqzjYhAdRXS7PVrjMZS0vHzUwxupMwK1Jc4ZnMziw2OIvOHyDJvv3eVBnov6F
B+Ftvmv7osKpcqY4FEE1DiTE4HAgXwiLIn0WsmS7ThY4uiZTSJzBjjtwkx5sWt3V
ShN9sbjxHMVg8mll+WKu9BCAvclCbLzmGQrcc9ZJGci7/CSInYccpvzae2XEY4HJ
pMwStqqC1aqhx0pQFShiyYwoHAhMfQZ5AMw2muUw6EFjiVdQWGpATm2PIRARCTL0
+woZGLD1cCVKv36+kAgfDt4nf6gJHOlhH8PyDFhIhT8es2ieT6oVHbCGNw9QJ2Ii
pd6LNPeXfbqZX+b5XSHERtrHl5Yfgw6S4gn1eS5kbtyqNq7p5vCmGVn812GsiE3a
/yQTHAbauAlYhDH6HChy8hthVUaeA5hm6GhiMtZYuWJihu05ny2znLAMTUqE8bp/
nMzY4RKHvnCkK9vlshFGRDfNpiRXF0SPq/00vjHTQb1kHvsqOkgfWdJHUN2IzYAI
n/mUg66fsmrqsppuWN/gA9nFDr4fOyu0yP7cogsnCRwReG/oXjqnYeTHs3CDtcbp
oZT3oPeNVx67leC1au+BVBi3zYDT3buIgnRHHNsfVlYjYeBuC2KXSeKrXyoTETYP
G+J2FanszKN4M2+/CRLxbrILcRFXIE5JTcIrzrrngzDHQwbZw0dDone8O1fX7kp9
XKpn5Xg6Mdd7UEBg9cyROD/qTtLLG2DPIN6dwjfq63Y=
`protect END_PROTECTED
