`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hOZ1rwJ24RW2H32mxc46ieIEjd+/lqUo/pasWgYM/NRXXs4P6ZwIO7c45fjyQ4C
FXgyljpnu7OLZy3bVi+f7mCVy2VXoypqYLqjDynUVdBwfxB0I6r6fiUOIRg0uKUE
bK+ywObspDgxfh50FB+jedqmuV6/BdwYSlf2xCihiTUzjUargKufdtMMBaW19Pmx
k7Y7iMTizNc732tZGGuauH3+kolmZWg5FgjwXDwAHk1ebydoCeBxhsrma+h93yQg
QzxnFxfRinwMcgyvfoT3vUiV+CTRgpv6Bvn3RD4S+eznk25koIjdab7dWif2U8er
qaEod+EuxeXWqotQUxqDMNxZSEu8qzLHt3NgkIFWQEzJAstqDpewUGUi/lADNyox
FBkgAwhhkreHsR7+wC5KEE2jHsEXMzyT2pJMhHa+tQennG2t9syIOmojaDzt3zfY
KsZmeQvyhYulFZtSC+8gdWnTci9gwCT48Z2XqhIxEw+8V4j9GivT5EjRyAVQTQ4E
oi9zV32O64VhdiVdrOebFNY9hXEp024y+dLpiM25vzLdn6KrSTY+iBiVE/Rzqse5
aPaYTdTEeBoOFxHv19YyaZpYwPadnJfFA5hPKiXrtEa198wtfDyfhiomrd+Y+d2A
hq8KZBLHK/BBhRlQXquUFk5TomFw3YSfv58N+EkUsRmK/KSYizWOUBuZUYSYbBH+
ib4AyNyPL0KpVXpMMpLbdstdB5XCGhkDUWwEFWqXDkla1er+aLmAZGvCfngmZEo8
j5QBAyWgOXpCCbMxL6N3E4spWV3tBUry/zuwpaG9OqIzK1PPpAyxWoai74WSYbGB
687V149fH2H3nab4QNgX4kBFSBIxP7RcPJDOFfD0bhqfsX8IhOEGXzg0Il17Jlhw
2aAKb0B01EjCUBnagA10je22dB6xdSQwFEOXyUGdQ1a4iEjgrgS2Q9exZGmqF6S1
zm7hMmruf1/1f+VCTV+BMb/WwDLJRzK1hMM2+ZSgpn1h1tTBag2nFdqsxsz8VZDi
ovD5Z8mzB3JQYJ6QIP3zTxcvhaIw+POr2NDXpcvc4zju2xkGdPHhpMy7Cfv8NKfJ
m15v0tPU/0oXELhF06XBs+vJrkE1qcpinKwc4ynuY/ZjCdShT7J6KgJImzcjLZ/y
TI1P4iSt2+zbkFvMQZ6XqtVl15JLFmjoz2WYD+aLi7UPArYmZK+V6yT3aVkiT00n
fTT0qYJo5PxHw2ozbyx7cZWhtv3CW4g5KwQw0kNj4g0+mM+yexELAA8V3IF6bMWX
52zn6vzWaaC4lifs4egNlfypKtDfaSeR3tfRl159kjiAOsPjd5s2tyodaOt/0pyN
QDrm2Xr7R8YBvrojMm8yQ+O7F5NoBFpMnCexMCUMn8bACq1Krs8EtsFb7tC+eGJr
syx9h7tIRXzL9EVPxNAnGsyBbVglMmXTgtKuGKb0ifpsSA/eHuBvTAHvTNst3YOr
qlhNYOw2N5QY7udAVOFrhubKASE4rntk9bH6g/jAMbIkHbDYexyXweJBTndX4HX5
h1nZnhjO+nPZn2twL/bMYWDQrskLZjEpZMEdT0FAr7kXORACPmrjiNVLp+jd9Z0K
J48Z+nH+IQiY2HWTw3q3DV8l/TYZDqU5eRtdnpRoOJUBNKFAkw/Fo2PmuwCOGtkG
ydmnYx8ck3hTeKzKGklFAdarmj4nUZGaTFITctQd8l03eVaR30ZztqoqY1OGMJSw
nXFN7Qjs9o3+QvQPkrj5wozurOXlNeS+MRkHqrqzyeXcV6mpRk/ZXWiheCVvk1Ct
/aH6k4Yf2q8peIFiLTqFjLQeLHzUK1E8XkWZBtpJcgymIwiHZ+tpT6E3vBINcI3X
NRuUlqmIl1G94GWveN1mgAX2Q2GYjv2gFXhlY1MzezeupEHznpMwFAZRje8x41QZ
jHXcjJKy25NK9Vi7zSqRKGu66w1KqtMyXxnRZ1zBnrq/Sd7UwuZfVs99wSYkRDda
/Gquuehgb9qmTCRlJK/3y91fvl4bdRRNFx9Coch5R20haP/vUHac5/8fOxz0Exq1
cc6iUza3j+5sqDsK6sCEsZNTu4irAB3qQe3zLxJGD4+bXdyD1zyENJJqZTudPBG5
HwlXR+6ip0Gq3Qv+OAfiMpC3uDAr/RfEZOT+55zbOB7jWglJgC3kKR7gA0cKvcZ/
DBXpNFk/+nQVhrn+n7Edt1i+LhgVGeq6+C9vP7OuEXq5okYPRQeZNrd8q2Puphm9
+VKzGjPWTtM5oWclnbQSGfxKnPI3v4wvoiu0LqDCX+Og0K8nJrmDFMhdB8WYZoeO
gyjEsVbAE22a9soUf/uBYdmZevfqbtMmHR2yRkBJZk3BHzTdd5QezC5DzwxSZSW3
bnJBeAPDBBZGL8k/AyIh7+nyhD9lshsNdOsbsgUOtOPxUSptIUFrBJoykJq3bRM6
X4oXEHlrdhmHUi4AhJOxvPp7dLnhSccqFQXbaNUt1qnm4/AmmRpPLhKmA6JXOjfy
sSZLOMvV1+AqeX6nmzdctHD4dux05Y9JKWFqvh98hdj8Dp5+VWkfjayjuBcmvofK
tFIObeUhH6PPmHG32bkGy2YnCTBrP17kcjiZl1EQTaYuZCu1qAvtMkg6wW/ZRZoy
MEFrbCYEFnDGHpZ+IOBTD2BcsXYpu/3xiUsIkf5PLr6utVpOUwty0FglvOFfxXNV
Swe2aLCsN4ptGwYVvsSLd0oK/H5PI1QE02r/pyiTvT53xvOfzfuVakoZl44fiQS7
cau2Z5g5eqpGsT1XwyTg5lYmlsq0c5tiIBlv0Vqbl3AOWW/Z8RCEMTVWCUNhPlEh
w2SlmNWCZ66HyxJg/VOBqkOcuZXpudmxKrVSZZ77jfyebMO2uK+ctjEqSC5YwKP/
isyLwDq9iKRFshhPhqRyflYKwrJnF4gmJ7iaiVF+hwjc+BKIac2/a089u9Dky/Ez
EFpp142Eio1742LrxIVl2PYCCz0IL0cqE+x1rjvN8vmf1hUSJQljDur7QjfqdLO1
+qTEjLVich7kfkmW6yEqe8S3KXB4i+VoW0sd7k4HsopSzws4Odq/2vyrfdCfvyr0
MpEiVpPKrzfGREVr/62lBS6s9zGv3VEiagWO0ZavdABEf3UPov/p1VmmD0BCIYiY
jTvLvmetImSztfYx05RSFvBoEgxCpcj+CI8uP+4UGwuXhjtAVE6mnVnFXLtE4+Sx
k/LLUnkIx0GVpjma8igmtIV+sRrVz6LniOgZo5jakfXgy1CzJ98WXTPjvsT6PDSI
7qA8g5ZZhTARilSFZ70naNMv0PsjtxJ72uGnEwI9Qso29KvzsYDjQrzZx1z1OpQL
LfwSjg+MAZ9Akadv2vyaURmI2CYbCUNlusGbpvfHmNZ4n5bXHDxKnCMgXNgds/vE
Uin1WSNAYvlYrKgRyJFj7RHPPekQH/Jwwekel89zXfa2SmmKMhIAXFXveltvFsGI
OTVHEdiMT+7rPEHPzOF/8iS7OphArqgq96ngNaVqgmymEFl+IqpWG8kuEqjPOX+x
GOzo4wVc3Sf6QbRDav1QkRldY88PxLlfYOX14KtqYeyO8XVHgjyTsFzQVCCX0QkG
XxfYhDEq4SCBNqGDYf6IzvftUwPiogBI3ahAVFv+HlLz7lsJ08U9EKkrkLQ5/qML
EXm2WvPCJeXND0V7DHOCX3OR2A465fcqol2082bNWQxJOUa+tLyn8o6A2FL5j9/W
QmLuTQmAMgIPl/OXuqe/df8PckNdYz+spjX0sUS+FQbD7cuUiNYbqW4xJ1/xjJyW
xt3AwUD/yVlioWah4GeexE5iOX9rVLTd1htghoswdRzV3c/AW4LDYcxH1+8M68ph
3KpjTl21/7J85jU3Lyy2WJyCwpzwegYeZd34BAV3rqdpFKCYc7mvs1eBI4QnTqkA
TJzpn0u0MbInNtGN+3jOYKiGRew1xBJZJfMrvVsKqJPDAKS4rtaF3FzPcjeD2cq5
WaMjPldGO1oxGbcehgKz5fjr3YSkejbAxUO6pYnRsmy5rqLJmFg8S652vnzpmRSH
C2rm3otlS2vXl+p8lgTghoAZHWB4KLrm6CzHZJWOrLn5OY7FmUnp8YmAyYbj3GPd
eifNMYPxwB1skWsoZVxT2C8O1fHjaFFfbE8Aj071iHlqN+IvHga4ihKkIfUwpX6h
O6LZHMStG5miwEIV68Tq8g3Hcg8XKWIpu6A9atuG3n8Qjo8bZGVoVJtfxAaRXs/E
liyQ8PUb5QFdoHr1XWIqlnkq4CgkCX315iTKe5gT1XJqrJCpxX+RdGrtOuu0kXID
+IUsp8htyhjwk2ri98lDHnpB6xwHBAtFMfSPFEyiZS7J7i6zQm4gWqhp2FKSEdmH
ZG1SSv/CFmTyazWPgFk4zTk/rjfcLl+4ZxSl7CJ+yyJDt0Fcs0BMAvzaPA6QvLNR
UVNKuLFTv7gzd184ZZ2RBUZGnPRYHlS0xB8grrm1EZZaotGTH4eS9e0X8xgu4vga
AAZ5OKRInkQd9bv7PwSFshCRnHadC8L4oThGy8USsYA6n4x3YQJlBmaC5ZSPeoSW
9/s8Pi5+xm8IIqyubeupAvI4GicJqhNTKX2/GDGRA+4XB/xDEXhfZODHcRDVe011
gn8dAekxnb+x+z44CIGiEQ09og9fEPJSSRlWlQzAyadcUgwSiE3u+nafXN/otwuK
KEtgdlLXLDgLqsl2hijKMQF5u/cyjvNBUPM7WpnmF0VRSf4qn3SDHa0rYTDxboFT
iiS+lHg8PiWhArF9NZtsf7j+K9iWxacOcgDuL3Y95USa+YmXptPrHY41rmBjdmSZ
qUgMH9ZkEYQ8mYK7i8xVMsTDC/ODgb30peFxGgTU3XDLZtMzCaM5QMnUw5GHNCqB
LG60R5WVZ7lmTbNLB32I3n/DcUlFf3NwyQqTGY/KxIjSnYTGFu6QmVgY54txexiz
GWENNqeFRXHmlSaSPFz8ZSP6Fu5OF5CQm745VpVntmDb9Gd/yJt0gRW7gUjGr6hh
nBLZkSvHVtSsgGx9h7tWOn5Vbsd/ZHl5QIV0KwWLN4FCMJdul+4vSG7ws4tCCHEx
RFH6i/RFeIyLEfLMrtARdRFMS3y3dQBGY6k8VOVwxeZsSnpupvRcvPaoqpIE1U0Y
5nAdV2Y04UDOH1BZWo9LtnO8WYKOkJJlHGmgKpmXRl4uh3yMUErBupCuANC8kgS2
HyDBow5/iX4qKXee9xWD7rfyhAq5QVMEophzDqnIOdR3/cvY6bdUMa+yG26GFXYe
9ycsHjAU7cCcrLlVhC7m5kbatijC8I9GnAGsWRoWCrRpLTzBFrtSyqcmp9DhilbO
PyIGnsrEStKJEtuei7vevTr6/jt2OUUj0NdD6dz0kJlfMVRB1STcP11rkB2DFD01
d+rZszQzF/xhDpKMTBU21ZP5FM2m63Y3i7ZCxG1851JDWGwKa4cycfozEoEApvX/
iqgX/El/ihm2V7Uo0P4cXVoH07C+9qI4Zn7apEomGjmo6hvAfcEJaF60bmhKVfTJ
jdTJmCfXo/BGSWsL4Qo93UulTLQsDVA6AZLHFV6P/HMp5DypeN7ztFvrp492/hk0
OXCl1I8J6LI64i9BXg9EDRbWLr6yrO0XYWsBOQSiu4US81wljAHg72+IbMe5Y9er
NbFgHF4WneCfqqjnr/fz7Na6iuHRoYtAow3E1sYSRtE+Vgvz6b94X7GoVX9c+/P3
3+8YkVIYyQBLZMZq+A1T9Q==
`protect END_PROTECTED
