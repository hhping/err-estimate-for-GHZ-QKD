`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4XARB/m/1A/kolZDFAILcZcI0KLJQdK/vQWA19U73qwHFnP83Q3+06K4bUDpwlZ
lZWlfaJABu9Rqn7l7Mzjoe6jgnssbtFK7ppsEVTnArz76NR+ci75aD11E0c5iuwb
7TUSs38AT36GJonIR+LHs0KvXTvMNNWkTe8fRzYld5Wr3vEJgoDT5W2NJho/h+Ve
TvdhteCFpIgz+Vd//7zNccSe2pEczQ3jzRgWJiMpVf4PJIwp3E3o4wdY3b8PIWh9
2isXLCK3Fn7Owf9flVTWEtbpxb/kD+L1WPOi2dPo//jnQOGnoOHz8d9sd7/ivgcx
K85fHnNLHWiii2IJ8LwQoZlx2x5gZFjgebMID5MFdVXliX8o23FBDDKWybdW98jO
kbsQQefu8weMbKPq/MlWGb6fSEdJ8rKRU2qcUh3HcOyH/31w5Krvn0eC2IZocgZU
u1I+Mvqg1+Xz/uSRFVuhKYbNqaN1ToZBZc3jccU8y4Fl+w89szdF+0UzQwBk75Ai
f9ks11unfmcyVGijljRKccGJWDE8EC0KiVY+gvkspSpVCpkYLg34O/4dVB+NGzpU
FdlrRuRIGJ5ejM2OUfq3wWOpquoXudge62s3WleITi5RdOXeSP/sJRYje2+jf0ae
PLqPn2TkyH9MtZ7ypJijvzFuQsKG+rcxVYILO4JyNY4xQA+NRr06BRbfu7Rywvtd
1hqyKwVhXYmP/ETtX/JajRBZaCE8BtIhv49DHkMrodlcX2DNiLo28eCJITzA+6uU
RjL/2rHMipUQOuwb3KuNO14zhoSPRQak1pyQqmTmMtUT3XaKmk/zCHwqg2W/eI1y
l8rh0+qWhZeWpyus9f1A9MV5onHToA8qpvIeqUONeY3Tb0IajXutldxV+LU1wJcX
GpG+VkLIMZpKvBxT/1conyPv10IxunRdlij7idwBNP80af8n6oPF++BfML1XFLRZ
+ckzII0uTxti/1rv4YdNvek9LeM1+mmNc6pQj0FSJCTg9JbyAhMgGV0OymDSDHvx
pRWlNht+d/hFtiPtQZ8diWfkdGCj4eh3ZVrlR5iHTzePpDdkXzHgnpKIRjTd03Tb
c+jz4JHXSS8w32pQruvrUq1p8/GhAZv51cjnHugYd4qFaYPMIJIRjHnVr8oU+4Be
KWWWAtV1tMDyNoJZikW3IarORtTZgjnWlEbJKOtV+YvWO9S6yDiM7otts8j1mjpv
P4wnIwvjkhgv1mfF5luR9dMz81u5SjbaucBqLzFhx2hsBqY0YWXEh7qTKD3QdWEe
`protect END_PROTECTED
