`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQHOblOMWrMdFO6dbYksCMBP7yACCMPnYBHqn+MitkHRz+gHJe83YApf/PKmwIW3
Ys6lsrLI2sCsirfnH33ERejFHmk3M1RuSrBV/xn3ClDY9vcZVGR9+9dUmzODGOjX
zyTR0lQGpUYT9bJqnbHIImbzJ23NZMm8erXgbnMflHeHc8F46ekOCgi9Sk/yxGEB
Hxd7JgnZ5sGrmPbZ0Qp/lpdg8uzJ8egcMlNiQ6eKF7vWQAzboKFqtWDJpf3w6LWc
5JkPADGztVOlhaCT0jAFN6l8bvH2iaKZn3qTiS37uCVeeidmPTF5h4W1AjcCQrIL
sjwNrabR21N6y6gXubU/HV9n9wM5UPILOC49RA7zwEEsbJeoTSFyR/akt8oZhW0t
utVy5vQv6nkS9HiLBfUaSNliJpOOMEypyJE1xwXyWcIBQ9do9rCWltrLUiT0OHrQ
VOoGU+aB89omweBjlgzMd1g00WZyZBqRHpsD0E1R5BVxqmrbE518DbbEgKDAvCbs
ADAXvUDUR7yJdb4UxNc03wB73YigWV+t3llCU9wHkWqrbQhBpptmliAAWLY3iZ2U
LjKmhtUQdSgFm2ufnGTifIHeYqqRE9WvwIpLSN6hyhCj7PBaSgVUorYm68FAOcPK
dbRZseti8hmHFT1XxzE6L0uTfWOMs4pBAaoUxUib00bCYPrcXxQ53C8JexjN/sHD
uWsqLx1ZQ9K7iNqMgpF1xdsXftHxTvkIBpT0z+kLwZ8=
`protect END_PROTECTED
