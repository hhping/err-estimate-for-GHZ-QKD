`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLIq6S0bzIUgBqq2UCafoymKAhX+afl1dZPOKe2DiEngGlH5Q9h2vTtAa8ea1zLV
GdMchGm901tEPzr7irDBayjKmtfFyyQffypC4oG2RWpWXOLnq6aa8C1nsd+32M0g
oaogjBwd1Qk0mipT5wrjikz7Dfo51CBuGsb1p+wmdXlCiCAFD6RpxA6w2qk58N42
1z7CtVydhv3HEXHOCGbSvsH4WyXru4rtzvg0UYuT68byUaxoD89hlPqhI8+t9Spm
b1T6fIxIq89RalEhw565SSWXPsCfwfJMNQFzH9rI5w8ML2eW/WuazawxVDbtJOKa
IU1MVHZEt8/VSkibv6StkV8FJongvOishXNWk2q38nlhH2O3bgAMJlA4p5jFTwxQ
ZCkmUD7Iqbv7nrsDOVoi+xhQ3Ii20PiNtsy8UyOFe7qb51AniApv8cvRHcjLR1/G
criDkqRzLSrJX4M/uGf17I39HjTlKvRHO2LUgbiIRZnfXUhnFT8xs1Ns0QVkZMNI
T/9G0sjjrNUSOLqPfqS4E0uxOijFXuyS8K0KMG1m/bDV0SVY1bU7+X8frkLqN+N3
JaghecOzwx9HPoeKIc5biUOIqLbch2GBpKuZlDyVJlsAVRMWszvzaCIDylxM2umu
IzkM8yIrBVL+T3ychk3D8+aa2hFEp5ji3zh0K/HOo4u43bD+x12XaRNuKZiHz+uD
cstg4w1O7cLZXHsO2KHr6vWiFqw4CjT9CnMiryqrbYXibzPpa5d2mJn7gIrgRl/C
oYicMUYUkPtlVskgbb3hMg6K2oYtslkiqJ8HJ5X4qXPzyGgQllOFqP/xubnnjVsK
NEw2Pf8J1PPLoN5D+Y+t1ol6sXnv37TexgkmfS9q3AsLF9RHQWMJEMofGRGXMYNZ
zsDY8Q/aC9KJMVvLZfj7iYGvFtTjWhdfxZAQnN2cH82XkNpVMsYuOjHhHioy8+wi
JLwrY1eTS2rNuSYUAFe7nkXC8uaA7EC8AxDpfV7a0eKolGBeag22TpLnJbSJfswV
yBsjz1xEjEssmUpMmfpoaDTwkRQIYpUV6pdp3N0o7w2ATNu3edZW2L0rp9efRSnq
ai7ilx9XH65UTANSheiZpDaMJNEfGjqPIpJdhczuPxRXkA9pWOkLL9XAhQYQeUyA
pxBfzQ1kRE0Rc+Q+D5Lt/KHoFNTgCLJ3wT8xe+IYPD9XLRrXM0iYqsjbcovCcFgS
GnPstFxmlx7GODaCTN1MKh5Jw3dExrLnt4BH1HSCHzzn0qhLV91nRtEqA7SdWj+T
8kacbFDZSgGAF9HAx4svVI/jCzkRi/G8/UFGvIxkwP0zZo+UNNcSlz1B/wKxMwMg
LlRh1mAPUjJx8WDjqncajZ10whLbSmEnezceOa+M5rFKHUS9jjd+edjHi9WvaAYT
w3MAGL1TCEuXLhGR46Gz+aCgAHPtmhRTD6+mhwCx1C2R6obdTItjUp4T7AAo0f47
MV5FqFqM9bqjm+Iv1y0+4Pu34YYwbRd5sTqrBZkWPQT2etwodgN4ztlmoTAXGZGp
oesDEXGh7a/3FQn8+3RxbhRjlGfRyauKwIQMFmmtHYuhCgbN1YslGqTwt+MLNZJP
pOFiHWD6qog6PsW70Jdj4lnGTaLbND/LYEvbZD+LxYzSP8f6e2Z4TdqHcWzae6dy
z8FYTboHRJk1AwKUvR2e426Z6XWf/z3cKYbb4/k9PoUYB9U923n4RH4ArBo+VPLy
iWOvl71ojkJiX3FJWPc/4BmGy7N1BzK7gYKgHhCWHaFeixDtDVaM2KZPd+TdL4hy
KPWHbR8XryOYk2OjS+NbC0yckS0p6JDX2NcEmGix6a4eBsKXWR5bsVJDTjobptWE
SnZbc4Ln9ssgGCKzEJ16CVCtmNDlDtN6dwa78zawqdO1ZtrRPUWuEO8/Jok6w6xJ
9QbaO7zPmwsRqUtWo+eM05M70I7vHMAsEURCuPOtZ3CjLS+NdpE4jqt9EyCTvTsh
pGo491N1CX+dv9+o0YMaKvL8hfTeMuzzuo9i+f3zJUkq4iQOVgjqO7oGKZ/4Azb4
PcYyjNogSLPskWU4lHFDsVeM0EZdJgAi55n5uLOkHIw=
`protect END_PROTECTED
