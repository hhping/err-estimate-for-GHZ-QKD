`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJQnS/mzuRP8D9fni1JfKK1dIax6PksYFJZRz41SSjPFcEEA7lRy4ih8f54Sa1Fa
3KcFi6Pg9Q+65aLpAlfMOYeZFtcdsdl7bG9k0G5qTJgjB23UpNj/Zrw3YA6sChTq
HO93Hnlleg19zMtqfkRCmlqu/Em5QnAhO72W2SRGZI3uzvpyAFNdadHwHuO39v4g
gQw+9fpMTQxcoL3bsCVSuQpSYo2FRf1q/kaEYnmr/hojpzescV4rhkjuKu7j0LpG
yGmxAhDK+myk/H+tgnb/T4CFca918MgyTsKPn0tnaiOzr5j74OaSP6kpeTROP7Ka
UCuUZtfxOw7uUfN+c3NvE8dbrz2P+gxbutxGoVSE4bWxNJpy8V5LlIXsA380CPRj
nn5hUUMEGRHcnDCpHnV98pIEmCWRcT7VDlKPhIPQ0TI2ZhP6aEGLhwV1XW8I+7/9
TYqr+k8o/FfnrXVvOFDhGzZt3fgEA4LLPuWVsQ4d0Bb4mHC8++6lOrVw/zRDPzu/
aKXTkeiw7cKUnLH56btKrbIh6tQCXJQpqpBPZUQQ8JKitbRsnxfW6XBAKKl5JZY9
TV03JdggiusqcKzWtifMCukojv0HuQvzjqchqgOJC90A+8ii8Uu/c82NzbNHzBml
ZbmnJ7+ctrs+BK/Eqn5qhjji3d7d4B/iCPlc86aREMLATCaQq8XybEcceZwECcg4
4UZwvQDaeujIElqZfzL+3IsdhotIUt0XYOWo8ZceNlDLxPIRM7kltWnMvVvfWRwE
jj6bN6aNN+0uVPANSFra1LxB2EevfY2VQtNkv7DreXKH2nd+Ne99bc8y9OcGqsn7
ufG/qLgL359maXzHJ/wnA/J2KflE6wQuwUD6cFn05ZSJY46o6dZAEwuklNZoIyC8
kwJ4JDc4fxbnX4kVnUVqbyLvJBlEuwzc1wHYssLMBXWDOLD9sr00t1oOROQXKJ3F
M7UgCuMCAmvGuS0Eat+/IFl2+R50ssThuv0oeyiXq+G2fNpvMiuYYVcSrNia8qX6
XEsZea2W6+wkiB4H4F/p3lsLeu9QrkOALAMfNytgXaa0+/eSlDIhqTMSwyBWzTMk
Vto+QMjqmGQ/6DJWMvZZlv4eiwUj+5a9VLnAUneu+1Yz2oC/OIu41AAv2sEeA8Rz
NmCtfydhlCzUQ/rfTvy8HEj9yRMjkyGYVZX57n9A8LCMfTWW9fry8hE1hcxdTub9
70ROQKvnH8DJ1hhXF5tNQVmvhH+iasuZRnt6IpgHTElFiIV/5f88wEx0AAFE/VOH
29hps0fbcc09xYJ34LDKinL1vmXZWwoxEkddLxtpHWlhswyQOlfLBpZX97U4hY0F
3TjkxrbPjL7IhJliVqzJJ4q81Hq/2S9H7Ji6epG+hUwemnFgNVzgZals9tsY1iIw
LlE/DaYwvyrlXf/jo3Z61gBftPGzIEz3Bf+6lp653cJYWqluqE+EgYzNb188QlTS
kPh1L2YfqOkwFFcwBbQF/w9BlFB6ZXGYowadiOkv07Hc/hTt68UTGZwXyJtDxi89
M8vYUIxqf1ngmBCh7pI0kKbWaKDctk9POGPsrvNlh78kT8UBtkYR4fBbxZZPB54H
OtKZmJOSwPkvGddYH2Gl2+x/cwJG+u3GwOWoA8esfzGNteuqccG02fQ6MRXIqL4q
MJGmwBqEOKpATsk4cr9W1usRydCis5Aqww/8MzXFuq4A4NQm1uUp6kG74Jm+SubG
PjF46lXLzWert107mXkfwHzWUQ4WWB0TDEbOREYkHJ0b+eoqwvhGWTq5uHdIKd/j
VDATcZjJT6osGoYWdgDrWnjxN7q/ye5M1IzsEH9+Pej10OPO8fAsj+Ri5LABNUQw
FVmUHoZJpJ/UORRzVt+Vda58UCILyC/BqPs0dVl+RPwrZCPJ55ew2EdipCu0nyVG
t97dkPdrLhwUKOHbDIHqP2/zWImBVmNIIuWyjPbVTeSPgyGBity1Jh3aCWeu2c/F
wTKHC56OgHOJkIi6AuQ2KPn00UcvmUMSUqxEsMyS9XPDJx6dIkt8nR6vx8TGd4A6
6wTLaXU7idu1/yfioCA+6VM3ti5we8NrEvqq5YF2Lxtlycm8uAuKfAprfdS1gN4v
9SF/dFB+4CUg8ROOVxx1kgQ7FCDFY/MD9kX0oV/c5MpxrjyrcBusOeP7S/cpYtec
fNSdQaTs52oB4tRBZvMFY4JW+BszmP2CARcynda9+I6UIeIJ1Gi8fT+XpbNGpXSQ
n6nIQBjL3Khprm4YrYHZZvXn/E9pzISYDsd1yWjJQ2o7nDe+T6Zxa9dx/06yfnh8
mSNT0WEDjWhV4VT8HNrbMZojwCvX+TrKXCY2rxNuYoJCczZtseZXDHJmRaxW0Th1
b90ZNUZQN407wQEvgdvXeY3P8JTgHnulWKUp6AADquzuXzZHup1401H30gA4cSXz
QB6lOaopFfTm28duQUuiwOfjwTp30hYYNmqlT8hJptx6VLR5Jd8VdXOdzhlGI9sj
imL0pkioqRXuWS7S5Z0gSRiSjOaaFhKjH7Zk8dxPP/92QOFitmsPYMXJWz8kIhUF
Lrd7VDUpUBXJ28G3w5u59YcaPcZyoi5QHE1Fe9F6dg3vqCvSbpgo5gWpRGzRm+Dz
Bwr4smaZSUUL9O97vSrQ26/Ebx9M8vykILbhbRZZ81dk6h7YG0iEvOSmJaDEHXb7
3f9CiLzK909ePBowCMaK4OxqDGfwAkJ/+0zqb9QGHPRGp6iGHCzb7shiY2/4rqwq
ok48yvcKGXOb9YAsDMtO22I/C1m1LmiWJOvo9IhN2NOBTyUSEgVklSYUCjAy9qSm
3ESDWy2hQ5sEhE/NUfkXQfcq4sdjW8NRP8gqU6pNVT+vZ4XsF4h5t6tfflwaYh3U
+6ouiRPboca7hIeHAP8yQL2jpQ0Lmu6SI5110Jia7JA=
`protect END_PROTECTED
