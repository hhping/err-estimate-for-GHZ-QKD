`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQ2jiseOFc5wwo6P0NpVmlvhCHpPg7OuheNxxLGVTv+TMl0Y1si6pl3X1LYH8nCl
BOeiG1ypWdUXD8PVM9VTjXB6Y5rTH0bis4J8N1usXrhGy+qFkyaADDY9ib9VBjJT
rCtprSAVCT3ezdP+vIWtqeE+S9RZK5wy2lEB+YMjZaYV8oheBE+TiG3eIn6ETgmk
WbhK5sx1lsv1Kqf+64pWfja5xbyXXQASWS5hdi5zBRUlg22ftaAVSHuoZdFh39aD
Cr3cAICXhFJOoP8+0ZvCaX1yJNBl9AsSx5nuF1KkADDZZFJb1KMvtr3ufnf8tEEs
C2eo9gY7nhoLSGBk0p8EOOtfOplp0KAdkcvbyT6v/9Xz5OTrdaukpByfagp5a7yl
eK7aecoXRtnDuxqGF/NfwdHqZ0Pf5IO8M2eO5t0d/+lCtpCL3L7s7SYhW15PIN/y
+ywsROIhYUyaBMbyMDMLkSlNUeNuFov+HcWrW+oDq7ZdhM3DOCZHN+7Pebjx4V3o
mMhH1JjC0DCAhbpNzZ/Pqmt96ubg87WqR/hta6fPI8s=
`protect END_PROTECTED
