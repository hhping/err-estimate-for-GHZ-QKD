`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
543eDfVonhgel07fQkwzD9kxMc0Xn/sdY5rv/62UywNwYnPGTytJ4YG2mLf3u7iS
hkqwnF+ws9UasfMsio8UelFmg48RrmATrVN/liKJZ/WWus0b2WyicJgb+bh4XIlX
aJ1rNZRcFMTTygvByCb8A+vVjMoP+opjrbUqAoL+9FAf6jyHpxyMH7c/83SBRU2a
NNzUu89Q6i8ejfQ80KAJwQBln/bauxWb2o8DQxIJ/Xe0+kCf6XhGbWdY8KVgQ7h2
gRg433IoGkKQSIBSJNj90gmVWku+nVNOH38515vGPmsz6+X6JuDV+UEid81JMHan
5ZXoRQckztjnXZmNA9Dpgd7W9AsFd18ni0KNJkrXEhBG75tN0zpjlX97f5Cen/zY
AE/Wqj2YKKVybhBDmkpNa0WokrPpVeA1yL5qNegwy3wwGaLQdFuPqqRr22UZpAHy
mydgcMCrggqJ1oqTIwWO89sc2Xn3pupKT9g6HdPiFHr7s2DsBaOPj6i10qvcP6cB
fP6PbBnFExFObhtUIA5e9kYUbXQkE1I00cZxHzKrD7pFBLUjykrv8caSR0eEQenN
gYZZqyHzmO+Cu8meerkt3WtF1c4nVxe5b5Ro6X7aZiYus9m5EkORhU16pfD6lW5D
tdGkYZz1HZkZRAVx1JIy0A==
`protect END_PROTECTED
