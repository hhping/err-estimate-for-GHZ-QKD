`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A90YmOORpzIqacr5yonwhW3/5sWqdKQihPNolV7WNAoSn0jQfUhvYKkM4/+p6Ks0
GF2TMrNrOaVIPErNoFbSYey3n0jX0O64KXeGlqfIOEO7vAGAW9FugIZ2oPK21nki
X5US1oC2UBEF0G98XpdrM6O/Enr74WWNx7LHye9lWSAM69d6N5nlJNv7h3ZQ/u+z
BZqTQbM8lpHDdEHIDTSX56wA+/95zf9BCOLnNa01TfyXjom1teQF+gKa7r+t8kGn
XFbxeA9CPPdSmX1qI/wP9N5qT7CkljCp7EwMx5NArxSW/yswJDag5HLoYjAAXSkd
8+JUW73ZroloN+5FCVPj3vA09ygQyKJ9bTd/lszXNM05ErMr8B1Hj0dA+EkkCvlh
6Dnmq5xoRy8PdenAcrfa6hsm+HP90Uit7LPYifbAL1uoz/N/yOVMKvOvsWQD0U9G
3g9APuCm3Eio+8aDvX+juDJA6tyCGNk4lLnygJSYFCCc2buJgS0iLKzI4rQDgDWC
W0WTRF4Zc+vobGmoN44mCxNGUW58gs9VKbblwaH+HjTH5aVbuRQMhddALXrvwVRz
o0HAbYG7DGZc3kC9hmlxJnuGS1OSOTlCyVQCd6RrsE8EE0nJ7Iwvypury9mFNuIr
bjf/Mvum0UFwUQ7h3I5ef9R+/6ZtqNVMJoU2Bm7s8Z0MK2OJRXMNJ1qq93i/Mh2o
h1LoZcWh75QN5poD5rW2RcSarNTxQSZzh2SJcjjfY1HQVzWFyTX1VklFzw012cFd
46St75Vyn6XwfLd31G7DMIUy7L+BRfRS9DRHvCvvNvndyl/QSlI4Fuf+hXMs1z7a
MnCeaE0QBeQrXqEUlKGhU71CDtaKVFbXcsKgQiHLrCK21mCixRU8WK57hQkyeN+g
paO4TRQeZ4sFZtM2lupZmWfwiJZlteQM2dLGVfK8XknokDmWQghFzgXpSDgGFsSy
O6jB/ee9kX0HKei5XuFBi22QhXgZUfrv5J9JL4WT3HkdDrKQlKNGSE4lYHOTiUdR
hrEEYBfZczgPrxl4QXCvcGiPUeR+p9MoryrdD49mtpkSvSCv1mvoIMIkZFfW7Nt8
F21yM/XNSp6/85uVd/0DXZOg5LhIJ9mAw0b4/sV6xKvm6UXcug5Kd8FvsBTM3IP/
IUq3/HLwcO69C94dHfNxxmiRJgQqRU51QJJUdzW60q7x7sDOCEVn3wClGcA4zA5Z
VhYTv59SKQKH4tbvC5Renw==
`protect END_PROTECTED
