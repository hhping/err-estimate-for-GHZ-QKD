`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4oHHKeL1aAxor0MPsIAfpEdH00VTrRIpRfceI3uRjIVUjbZM6bAX0Cns+Gh18CbR
uR6t/prihf2BRLQ9tEewUZfQ+OhHkHBzxHJ8WZ8q3aEVY6ueHP1fIZ3C+8crQUWP
wJVaegE8rzwxGaACeKpUkQEVAAa3VDWnaFYhn0W7Q87+7Ak3uyabSfSTg0CaHrE3
S3NOvGnP9UxWb3rJ6WyTrgi2T5DgXi4bBcMsSM53v+GOb4SEcoMEC0hh/Ruglx70
n0qhsNn7H1DUDruJz7iBDKWN+qnXY1J55dFV3oNCNZytlAwtlVb4BWcrBeVQlGJQ
ScH96UtW0r1bs4ULtSZZMws34GKnLQ0Us2Hp7rWpE8iYOIVqoxQKhzZNvO9Nzj1r
KdrxgNjFeXIa41nMV/6niQwIlWrwHEME5T8hEntYD9WLhscKhD4agXpHBUijWvxe
ZZK/ijeGJ3LkiD3KLM1Ipob6m8HU4AohonmiDX+F1NekwwevGDNdlCG2+hMTKizZ
uR+5zBx3zaTd4hAfrByML6DwKShAYYKRbo/Jze8EmYCzp9jS0hnPodd11MtOVfpP
Mge+SBZtMsUXOis6IiaDcDWpoje7xybVRnXOQsC2UwFUME02lbUCDHYzRcohYeud
nk/AjiTvLgKDU7qboLXKBPrIBkHs9Baf0+g8TXib+lUJJMozPNmZgvYNdtvdAx4g
ZaJnkgmw5wnldUsTzaT4dJsm/ayOcGrao7pggPqEBORcEzBeXOzgfSlVppLPqh1i
w4PjBRsmcnnd8BctKs28SdAJcUxc3XkWP0r3/Ve4Stt8+/X5yCIgBfA+b8KQfngT
ufJHj13OYVGQA+04KkRFVhLg66eLxWHM7uFemXG3bn/XMiBSqDLFS3P1v1dazEGi
qt/WTHil9zZ//MmcyJ6MbKGBdgl5u3vLFGPUyWhFbeHhl6b6WHzdTUBzv1CgKcvl
XUySWmbKSjB8LNY8B09Elx/FzPTYU8eq5orvU0ueYog8xWNKo6xBJCqxtuVtUCtO
USjCuRgZbPjG3GjPNQ0iMWZQzA1fGbbz7FPyRUC3bOLp7mL2sr3ZVzrNgojCyIiE
yzw4a8lRl6cKfkwWEZy/CNL4sjAqAnkL0n46aAqVh0A4FNtC80JbeKHISp9HXX1N
5bFgS+BNKY6/p+Tp3Zqjt7j2LTrMpdBHaCVIU+O4gRLgDexMAo/6e1GgyldaRf7C
8DoMAYj8e2BpIzJxSJ/IJtt3dDJKLlMemePhLSDknnV2W/EdtCzPBUJzhd6CpFSA
simaGU2JSmr/YJ/lGk7SwAuzNGCG8B8e2RjqikrD4REhbTovjB+glATH60NKLs7j
0FXaU8Pk3YBCStLE3bsz0fYjnYdvO0vWQN3SAZaA4Ylj+zHLxpWJ165H1dBkr0R8
3DV6UFTd/oaizsoFdYwwPj5mxpI/zx0bj4EB9qD+UqYv6DVx2aXdlv1qkldkzUHE
/0V1ItogowZsWy/ppvu+R7YMzFgfEaRG3p4qpMSD+MjczyPb8J44ZnkuNvAY9iOk
wyaawVL2Ayeq7eGreiAozo470uauddVaBwwO6BtSBbLk7nVKGFAOAhIkGen0R9oB
7Uu9Bah09gXNlczXf9eljPK2kWSR70ZIS3VPBOxvGMFZEbjz6o61VvMJm0C3Gdv3
3b9+tmxzG5fZbR6IwgaoaI8qJ3ZdoimOzcmaoisLo28zzaXvzaHtiA7zN1VmvU4M
Y+IJsQplUPqsdz20lfr94RyVKdvhWUhnyyzFcuGp4ScmKcWGeB3Jz+zmWnMouVmG
IPavM0Xpg91OdiCBJVosjU5/4+j1mnpXCUIrWqT9AhvhHM01XDrDoP5/qOC6VnL9
us1RfUvH/8zcaLG7doiUifU/XzyFFcYwHHw+J/ow81wvqtc5juX59bZnzzm4iUvu
lmMl7qRSr0q9PDjylDTvFtMKQn0woo30OmJwk94B55DUDdjQ0pdd8U7OQWl4rqxI
/GChAHKv6I/hZ28gHkjAIz6P2y7n4nncnEHtziAf1vHiRAxYNMIikloODhbCcgZ3
KCE/bcrDPLZxyBmVRBVsFUdqVRFxLEsoeZt7FRR//wNCsRDe+lniXuXcn+wxkj2/
9N0CoR5YQqdkMeG8EHe5lJxWOMgpB5mlUV0VPDMk8A5M/y5td2+5RUp9LHZZO130
hOejbF+sWWyT56p4Gj+1XQS3zu5GjpQ3Ozzgio70A5Dac8oUYx9CER+eE95jjo1D
9ZIBNFsdEf5C/q2XgI8K3FsfMqRlHc0eF2byKkLEPNBogRbjAtIjaXzNAWBq/2OO
qmQ9Hs2MzQXQX4/Szi97sGvewx/xptfq9ewYZxANXxtugqASoaaLl9xCM6X2GjtS
XJhXuV/RFmo9mQnoMLtZsAuc/XskoYlIFXfLIAzK/+C5qhxPqrW26cEiZZyrE9yc
W0bkwmDtj5biPYxGz6uk0nFg0SQtBTkMiGnvxbonKJeSesiI7iCzyUXYxI5Zqq8n
QxwHmvkcej3z/hNzoDJDtzNi7P9AcyxNAGejJXMwyejI0nNVvg5ScMIDexKJNHC9
Ax0mi/qJbR5o//M3H4YMWveG1b1//uKW9UOnSWWAqk54eKS0jYkCSSv80xBxTAXz
zeS+wdF3NW/QiQ/2lyyxbpaAXQD+gGZYuMMPGiEoYbFcXSZ1jgZs6wMVAlbcCQ2q
XHaFlycesrIXUxDH8mx9hhAHVp+xgHgrRGFJEJrPzBDj/Dw28+g7eacukIkmDw2F
2ShPRi1WDegn2D/aXrmbUqAcQDBLAEh5NfoYOOq+nsBQl0p2RUyvpxl0uWEZiXoN
UbEKOP7i20U48ijy2A9lP2nBLoXN2Sj/AyzqKLOAOKOhbuWM6EGVJbKDwPXbqRY4
W/6VUl6q7HxWROh2LMR08blGGFwLBlrzp7zsDiKwkRUgTRawB2rJ83L04R5dAcSY
GzYr+tmnI2o2wN0pvcZN1EU9MW/wBFsHnpSPJCi1Hqqkzv/aj+ST94jwrmcqS9GU
ba335UsjGbdwbqK14HxkQjrtPxfxQUY8hC37whSFPbo2Ji49e18en0Binz3Xo4fq
E+rMCaTVVJSzLSZXRj5u4W8Z97Hdy4YQQ8VUX/QR3HT6mAg8jgvr4lbTg1Yl3FbH
OmOs/Rrotl1zSNj8J+KmPMkB2lnODtPrRxXN+VjU3/U0ag/GWZPZibrpjozyt3X0
NS1CFQ051NtAadvEslGOnk/aLxpFDXtILgw7VKkOG25odAHIHJwIne9UBI3jOl4M
t0zRNmPkjB/gvAbE80lQ4egGH4Kbllz1Dcr3xHL7F0DZpOe9DRbFP17EBQnPnTWd
Kmf2BFOfXNlF/OBqHaqI+c+slH1zE5i4ld+19+Y1nrpbNo3SPgr9LJtkNt3ysfYN
5OZK9nqgrYI46SyPQejEioEnOgvJhYx5ikPrbloTYN1X5Omv81fjLiFl1Ef63Ibd
AwPtLtHCOlnYQINf/Qjx2GFx2Kc1HtFSwWcwgveHwh0GSlX8ajUNl1JKTGyU1s+r
DzakCaLYbH+iJvrUOEqFYENI/Uy2V1C/obxufMfChXZlh0QWWZtL31TMsI7uqnRt
8SAa2HJ+or/Z0wfImghhJxjgVO6CJE/fKj+a1xYfDwuIPYVFpsYL06Z9DkEF4vOP
O/DDQBJkavnRvpCaIAfm9aUZn6NA5MCbIhHbbVwKkru2Tah9iRoHwxbXhiiC+/Nm
m/wej6bQPOcEos4LO9xnLPvxZfFHMpDfix9v5DELCZDjWvo3ysdgfGkB1LdjSlXr
ZVSog9Akvq0EQyNs6JMapquxZJduC9YWCdh2SaJ5ynyGaIFFtjV/hDd0PQXHGjwV
rXXp13VWTDCov7cbmVC4abbhVpHSiqqvLpHI2OgU3EU4gC1GkhjvULfIR2LMAdyN
QpaJWfFqQqGlFSQYXFm9BAiR8woeotWxS7ISJL7CE+F7XJtBsaALgSI6Qcro7/mU
Isd+aS47bVg9jDDMVqe5iXRYcFdzg7G40OacKybbqoI6FdVF1n+h4QZ79hnadGpE
ZbA003dvK4d1lclYjS8aw8MsRrb2Baa830jI9pQlOGbxBiTxqIZa4rJJDFRQKMXR
LybT14AImvLmROjTvu2guGtQEr0/70/VEF8l5gfKuxDyEVhCwZvONwRcwKmEnhkB
v+sObFrLfZdZQboCPB8Knm6Hz0dsCh6QXHyRrOgvcl98UDP86GCav69Wii8zPlMs
1SvlcHaFMIQY0uH1zG+CukArLW2iHZ4XWiGER7IbPJKhKbtMIOv/M7FaT8e0g1nm
eD57+6+dgujKQxjX/Lse8xhpOgOxMfstUUDedXREF6N9nQMXTiBr8M6dr6yYS4r0
h2DrNclxYKoNyea+9ybdq20MBr5VJSJu2UrshzvfBvQ2Nue4oQdrws3ADV+TdpRB
kfwRk5U2KRNOoQJde41uzCg6cmirpSP+HeJr+X8Xco1fj0lbVCOCWenh/u2vkfqh
Anu6yWtzHG++ro0TEBq2JhkjJGzO7dK4U4DzI9ELWUaUDdVWnfDOjPo67bjQTX+f
vT49pFh/A46/rgJPdUljssbuUmCGsInwxby8+y1kMnPU2UaWSrKKnkWwf3sPmeCT
U8iA0HXBT2GvbyQIP0KxvQFmIlTg9Cm5FeAiW/LLt26SBytfCUQRHhDHsevEfkBr
31q0soAujxybMEQwOXcQe/CPhts2JfHexHkaAcDveXkysGkm0ZeDa2jtsNK6CGM6
v5xL9v52GuA0hO6x4b/SEW8uTN1MrvwJQ0m28aa6sl7MkSI3kQaXSDSyRmfKClZu
0A3Mg0eqDEm5nshF6hLZkx46CmXSxDOepia8i9O1JYgzwKWspIhV4yG8typYsIVp
D1+AHegZkG3iRyYLLjZ7UnyuNbXHHE2XFlYSwsyYusJu7dWxvH7m55fkdz+zc92O
uL59qYYGIqARkzVPqqzKfJpII+kmiUBMz8+gocMT2HaBRZiXA4ivCN0oeTYkAG0O
7vwi+H1yMjRm6IGMTHUeVNuiMjFD1EH1z/fK4acIaZoPj9SF1bd5C/Y+a+/myBZ/
OPsXg43wtKSHgXtTL9N7EDcLA8ClOPnctWg07lVwLaPJNsrPBRFhzQd1txLp18Im
EJJsKLWel5k80PqQjtudnNsb1SaMzQeD/lu9fQOTepB2CfQPtSxrND2jYcpwFYm0
XXYYFVNGMkvgPwsrakSrTCEvVQ682fL2QokelypWTpBR10BMP1J2MgbEyGKLu7Qo
bamT2qPN7S6LvIAM/DGrbCJkyKyt5GvtnE0cq1JR1LnF7JSr93QUkmQ3yNp69bn9
FbQC7UQtWOU9kTm2kVh5rvT7istweB7eVtxNL67Ny0Dfmn0CgpbnmKPJUvaD2omB
I5yfqoU9TpB/TBR8JFOkrhMrb8FR6elu9fVOVtdY21pngx1O1qRL4wRlEhWGFPJS
utgcQJMnzwRPkDiTovY8v2AfXIBUP9nOGxigcxTxA/qgCpujObMXVVeHRVXAdEuY
9i+9rpYd0XyT1f35kzj0K1c8tS2on/9wQuVRibaH19C5wJ8kNw3QNzi2UaN25+zR
AGPmwLIyJJXqgQKOeDiWGZbdt5Ll1/dsveo0Ps1hCv1zz/5r8fbuXEiOBU9IUcBe
/VAy5H+Wf4JqbciBiHFGFcHXhVoHJptFAOCMiLa7QSu33/TdMeUzYppTMZUU03qf
U5oMNsRs5dnSbVRKtlU2O7Dwly+b/347hKu5KZfOrtspbW3mWAaQ6eFL4ntCu4Ty
QYcX7J747I9FsrlWw33JRGaim3bBCq0dYgeoogVdWViyT2CuhusyErr+HvilXv+6
PkRIoIO+aT3khRewMoxgiLpFRDyOY7njdSr6Ri1PwSQfoGM5FBSGXq+aqvWaWch6
doUMspzBUGemQeY7CF3+HAX46ve+V4GPS3rYW9AaN99CFpYG2mFlTlQHEhrjm9TL
gl0Oc+Q0Ij4SHHdS/6VXLQba9LhEQU5BS3gnq47U09RF1IRBeCg4u6NPB/V8Tq3f
CvB81j+XHiubE7eDcpaZFrrwyA6HqHyAQ4sQ7ufA6S0CdyZEKBXx0uazzi/plma3
DhB/PAmMCliTbx1V1k4wAkov91qg9WMAQbCqVaNJoB4nvbZbrXUV7BzEGn5v2wza
OEiWJzPlJTe2gSYl+EGK7fy0KgzaEFIauR9PZXTPIKSRHiRBIzi60YFo67SkFRwo
5TijLQjpaOPHYzNT5MmbP8UnIwEJx1EdCQc+uPYELnUL/cUSXOsLGebbfhOWcAF1
eds2C2RC17pY8ndt/z5lkkdKZjxROEoRl+aflt1lYXBBVIM4IZDaaR9FPexuI1jQ
7WH0QZ1IjXsXseBsCc9Pgi30r+GpPiflZJZOqpozUXOGgUWWdOTNE6uahSBp9Kl5
OeME39c8Fe3PHUZwnM6kHsDld1sevUq+WuLiewDs+R4ECmOR2KU64t176K7gMk5y
gkAWXHl+BUxtuYIUeL8rajWuRLE5rAHmN/1mJg1HbDA7h2x1jw1Pla01U8ksIvoc
P7M4ZyVFdGN7C1VEa14XWXIou4Lu+QFGEkAlw9TmnOVi4H3Ga8LqU22FqnRwIRwj
l8o+/uUXgsbSU349ansDZYCzuFlHKUfjXjSb6KbW8T3f6Vm7dyoIlQzbczw5A7Aw
WWraMIizwpEoeeI2dA1xoxOsj9a5Iasw6OLQt6KpUVoUjOFGmZBPjvKNgBdVXZFo
rakNkC4hHF1NNjgJehKmlHENnsG8SP8p2v4z+4TuydgSpz+sAYjsHc1EVR4Oixlt
V8VsWqEUn4fK/1Fmk77ZIzrf92xtTzU06ikr3BkIdRAnEYe5Pp9rQWIoYwQyumKR
70+pTGL1RwylU8JDgPgd4ooIE1OFF0ivwmrEm4SyY7XHvNB458wx50BdozvjBxB1
q2vYxeZegfpGZ/+TNUY0dl+GUWyQqmdjxBKHy6M7C1kQakPb5wJaxK3ALcmjWg3F
2JGgACOdLJolnOWRsfy2susPdByL3sgrdgnWPbhOCNXxMGI6aKsgcNI0bFE1Ppl3
MI697O+wQ1zNYoiCeDP+y0OsoSUBua+ZSIyuyShpjSN0ovhMiqXNWsDfcCg6crwF
H3c4hhqPsfAMLzEg1rxNNTMWeX2dW5fTxk5tJ8LYJwtiJKHZ61L9AT0WaLyFu5Np
HYmPxMsy9Q0kdCRirrsu5I+bRefEITXfvCwnanPYpb+5w/9JKMBbp7unc8QaI9/+
OJCaU2sLb/RFlqCCmQQgOs61/EOHSKqUrtJ+D8N0zGQAucIHhUSSKBrUJvH3dGSH
o1w/ruGNhN3uHZ6NUXKGm8O8Gxs35RXEMdsisgorKuXHXl/sDK4aFP4hKMDLy9oE
gOrKifkQkmLrWo6VpSiB6e/EsqQYxW64l2c249Xm/YODx/eJdQX78UlilzIugJPE
n7zqKpmLVcv2R68Mm270C/GXCHjj6/MZnwYf9YX7TAbcD9wng9NnvsYP7VQvwsy3
bffVuhFvJBynh5btpYR4Eg6oqi9YFcTpm+nYnFIraaciWvkJ6nVyAEFBVXd8jSAh
IC9wUZJsEemh3mxkdOvXRL0u5JSqD7JVDWWwkzO4BmHNv9o70pQfcbjF4+kdJF79
gxluRAQFP8NqmEpGhq5r2IixE9G7UpmOcqrbD4P3p1lu0rYD1pBGmrrpK69Y7Dxy
nLVL0wcf/4UNush2FHTGtIFjRrqxLN3pW4isYD5c3DHeF17yQYpBAUvZZtYN8ARy
JJCEioOXbjHON8m69UGOnCdyrt3M9Gg5cjcuC9f8aL463WQFmS5GTc/0R++QS+45
X690tSTYo15qp9/nSrJtbIrtJ7k5/fLNItAKf+/2uH2wc81i5OeagnD6QwQxiofS
Nw4+pWS8VzC/SKJ8m1oqcx+E8h7OZxXNuId6UzXWEtwP3T6NL4NpU2oOBzla9gYr
M7BRZbpkcchy0tNVBv02u+MwpPOJqgCKkEqPH/PcX5avcKj2s4SY99EybG5gqfCq
saXdVabwSe3lwVilF+OC4/PW6HQPfJKh76efzUhC4+FHFdO6jFq+R2VInSZ9VIQ9
qV88fRXVctXKQQEAwti6AFLPO4anpRIUiWD8ShKPu1liWAQBVVFfRyIot6/iFg95
WjKwZzaSEWzZdL9VHFdQUOsXnSSatJCsjpi+Q5FpG/wr+eFwNHbNbqhGWNnHwv+t
ZYR/wXxrZm5to9QcT5nuv5WbKJ25Mq8337FC9HoL8WDBZThiz1+XHT998nouYr5Y
GxGMw15OhzrrhJlPg7MgAc050RvqRTT7FKURQbdDblHqS39kXNZfDwAnhLATaycN
hVfD0NG6ACjpZBX7qoPUvhLWhIe6t8h16rIqVTA/Krr9X9vNdY437CN8D9qkhqJ8
6b/kL6cMBr9wGS6SF5fXiREKHmFPt+f+U39ci6SfUzsZUks/nuUcHYArg8hJaB3b
0TckFXIQcxFseDdP0JPv1awHnxqnaIXSWzUCJb+MESRV4lR2s9aZIhPOexHoG/X/
O0vF7yV8ydW3eTWcjl7+rWnO3jCj0RwDPq+swcyuQ0D44NBdwHMCgA+B0rgTqNe0
/dhuiUpWht4vvr7TlBunh3oUkIS4he1/lhXjq3axOvLu6szid80QIXjB2mPHirua
OtP3JWY+PieU5pMq7tS06+hZbaOw1zb2uQ5kNgJAcHTuNMopfvGNHfITDUdy3aHz
kkz3xEzPUhFdfg7VuCQl7xQ3rX7Cb87kadVHKy0Tk99ynnsTqlvLXXLl5To1b4+/
FFRgqiKVmzNb0dbNYaM0gZxi2WqIPUxDfLyXv0cGqTG4uq6DHjk1j0FNBbEV4K0b
YT6siT9qmDF8anLsQPWH0oqXIoT63oZUfeDyT5GDBteIhayZj4YykRqvtGWLDdy0
li6Lx79XSEFQC77cak1DqIjS7Uux2rCjk4vZlA6uoIyg7t1fNXgPru/7LujBTgSe
mSlXssvkpBLny//iK1Ae+3zLcRbKSmGB2rMXELkroM6n20X/qegEI+ursdJUY6NU
B7mRjzqYnlXbkd4s8yJmI/KAN+e17q2WoGlr3yRc8WXiw0NKVvXGvtnGukhgcu0S
k51ldo7x1sCH4QMmUaclUSA3BxN2nrZgWfY6cTtcLg3LM2iVzAjO1K1JATYWFSrR
jbuPxhDxNfJhUpWTIqyQROSLYjW4xgMRQwZ02bkEYlgXb5VNIfewt3W09drrdUzM
0VoNcNG3mRuZOeBiu9aY1hEoO2tdWWv3l0OT1HUC7Smd4RCqNfyXL/6qXTicoKUJ
p5vLvRcSoOYRw8QMN4xzmkVisJnfqW1hyg7kgh2/aJYMmcrvRwk9RJga0GXkYNva
ca/C3oFZ3yVDeAMG31sApYA3fHWD/GxNY/14PgHSdCY4bLFSG0JK+e2RLAsdPhSC
a+nNpaRngP7174UAf22BHxDoo96HVBXRep1NKIwAF/nOFeVyxArcngcKwETgzzIc
7XIkVPl4Wq0f0zNc/IUXI0TNHs6pUYd/2CzKnPRbxyBvqzmNijNasTgi8KDjQ1sO
N94DLOgZUj4kRdBNWCXsu4RlNXs8AYlx9VlYLJXkhnbSFHPaT5LnN6hw/X/jWBWT
XTeb2l0LIPgW4uC00eKodzEIwx2wnRZNO8qQiuw2UH2DTNJztrpysH3JbP1VMi+7
9MQNlJb6LPdNwZI15ISK+eXPpIlpcfXYVxcVhJAGJ2MqA7rDx+kEHY7DP7pDk5uV
aQX0f80YqeXn/m2K5oh7NO4gLrl65S032ps/isOPKePqsEgP5lPo1TDu9gD1Z2YH
18fawdhsTGeQXXK+QKRUXKcYj9WvCZj/PU+DHD/pXYdF/HxAKMH30OPB7KKlvJjl
OALeG1SVF8Awi13KALsXcA5FMGxosp/vJ8rNcslbkTB7W6SZ9PkoutQwgSieaA1J
bFrBhCP9+UiglrXfpnN0R08NeyweIwnWGW97YBPlomF9BGtMUKndROQ7UCWuCKbn
Bc0Q5OvHJ1ODYQXvj56UJyvqp+gvBINu4h1c+rGpYw0oiPgu2qGwtSH5u5DnLm/9
DvFJIsyw6TSXQDrZYefXOO0pgd16GE1vsU5+hBU8l933wYpiIOppSRhTsGGsjIuu
6D1sb70EA17Yce032nWAyDAfP8n5AkaKg46s24DLbHA7Qd7zNOXmwDkPXhtwohlZ
TM1pFAje0rtw7jHPuRTPWJk3DEmFhQv+yaTG6xhdptANl0zQTkbQT4Taw6s8oiYU
BU6Ke11weqcNbqOcXe0Cz9HOHbB9UUnuNGqh2IEF99zJO4Nbxrg6VUxWKhX0y1Wp
6TUhCawas0deoJMbbMKfGEp5lQkqKSV4gUnBmcD9Uadz9120LRtbkLZ386CTYnwp
3/yqDBC4V3vA8FDeBbbBNDtVcZB/FcEzLiqsq34kyKeYqs2hxKMVA29HSbEhPiGp
T7sgozprhyIoi80YTcu5D5FmYYvoNnmn1iOkgzO08/yyVlD4F5+M+NuYQae7tHe1
6JA6z5cDgMK5tStmYwEJehguj9Hn6qcpegF9lAjxFR0F7xLwe3eXuWBfl5ud34RQ
IjD5NykaUbP3l6tdWPIDsw==
`protect END_PROTECTED
