`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XXteXZvgA5Xee7t1QdeT6Tqy3s6AM9OTlBN9mLPgjv3lxWKDcEX/Noiso12bqo/l
pYjSxKfCjiw7afLr1H8tYZec+BNvTzw+d5ySqowTAShjcBtO3tIXv8RfswvJGQS6
4LAR5vm0TMBhaCvgF0hedu9zw4HKhd5UTrW5aWTEIjo6uLuI1r5/n2CGyCgHma19
tqRnaw5K0PprvenO6r5QW4ydn7atenE87T/8ZCMFeLMTDadVkDYeWqWZV4RvwfLQ
vZhlKVIZtx2psOs2EvUlNq4n1o74pv+43H48RGc1+dOYoSw9IDiHVPmmfzpFEwku
Y4iweNfaf8Nz1MkMKHsM/As1whDgdWOXP2GDGXPztZQ+80pegbiYzTHam+n8V/Ow
fXxOW8drflTRfvCKvikbvNbnpLXtg4H64jAp/TmUPnbmhzhMDZpdb6NZVevPF5a8
fTAKCO2hkmncX2rI+5KiIJyNW8wWkYJEus6JEQHsD/4VYqi6axh05qWj6fq0t9p2
ZzFLHig1lr75chqhD5+UQYYzoslDRCsCwtj5HOlXK8gemC+m5HditnpcyIJ4zpnT
7eT3+2ssumOSLwABV0ij3eZ6v69xTJguRFayBQfek/XgacgjfBj4Tyh372y7EElF
yxxlqLugjGY5zfWrwjBJTcSqtkhW5+RTZLYp0uk/Zokw/Tn9Olja/vStAAxm9CaD
lGe5aHK8batAoeG+HPM1Tdd+91nyseiK0yk7VFU278B2DASdjwGGvsWaygXroyLc
LHkI+dCxWh7fEJKGLyw3Y912JhRNvmcgBuibqQVWDdoddXGWuMcuYmxfu4TEykOo
nraH+j3rqf/W/lb0p8xIeSwXcWNYdzwpeEeS7wVviKlrunq4ujy8NNxaWJ7d4eEw
lRKlAAbqTg4GiouhuWViORGTGZEGSNGM/0npokdbDTncmdNnXPTubVKgAl1grcpT
JGvXyw91I5Ruh2xp4HEiWnisnBmmH3FaW5To0Lfwh07bJlfCXgLA2YAkSiOoANFB
BYovBmA2LCrNnUaOfsl/LjEul6EbmExMDnUifSuPQ34g+TU6/kmK+h8m1IkAO9+3
NHggqWKmy9xMjZSfkBcmpr7hG84fPA8Ytd7GLm5RkMYLcqdTEyZO00YJRqImwqOb
VjFCDrEvJdI5SzzIzMEvL+kYAJvwwrjdIMzGUrF5nOUDh4S5rwJbR8NwYMt+dJrn
CQdm9HzqEu5oK1BOx7l3JgLtOm+hH8RqzohONkMvCym+GORxIkdkBZjzGqaBPoBY
37alRVrbbf725sqa+QMO6ZRtsmYooVMFESte1q43+wdu7Ix5aaFLVyUwgJdbFkDm
AQkmO+1N0fZ1LbY3Lh8U9QlkevSf7Rd6LhLrp1Oi9RHELSSL7T+k8U8wRrzN/H+i
4ecrTV/rQwT4oRl2cFc5wqUWdRdDxblvCsgNo43crgxAo9vEMYSMI8cWFTQF4pzv
YnoC5ON6qsNp1reyFZgRnGe1tWgOerSfUGrLepYQpS8zeASUH84U4JeJYB+V32rH
q5ZwabF/0S2ixWQO4qrGR3a3rfygnuFQaTCdTfRI1jST237Wkj15E8XZ1I4OTo8c
7XABx8m5hT27KkLC04NSFwnUP6ySATj9ERNh+GLWTBMl/3vnzppVCPPLFhcvMIzw
nlK96HtDgG29G1eHIM8b/YRFTyAfG2u+++ObcbEPVzSSzo3v/gFzRpKXpWn3EjM4
0Zq2DkwHpcGe66sorQvLoKRYGiay5+eEN+sk4EZMN+ptXSkqXeZUKaaaFGtzpvwp
9B5Bc/73y1JpN1AQSDHlr3eNfpQYg9Jl77VVoT8+2+beMi5ghvy5GnE3I7yxkfAc
+O2Zc46sCxD2GAqRLw0FU6QPJOM/8tyWJ7G8+J61wdxAtJwK4pUlLVdZUqGhzoU4
vjoVy0aA+83Q3iBf2POCUZTpknziwVfmC+pHDeqFhwMkQX90yQ9I1/QbHx48h6Sl
QWl8cN31SmGenbpJehzfFYVBX/PsL6ETXO+DSQqnLnxISYO6xw3OJkNsDi0z7v9S
1G3faqVcO3iMaASo2C5Agmsc8C22Yowp1I/K0tCK49m8Piidg7/NSfKNmHSy3gQU
uLDM8DJIwKkoo0LL1pXi0rEt6vJKDvv92GkoMViwQ6ojJd7/fp9HUhdS6R3hopU0
3LhE8mePNxqOZ2sHxSa/oVv4HEjL3usD/pYYwN0hUgvnoEnK2FguF/UIq0BeGhFL
Ngv4z7f9kTsbnIs/0YrIHYGMQjnUFlbeA0lJpNWZy2QA93vmrZYV4+XwXRY+pxzG
CYY1OAazVq+gJGHLBY4YjszUP6mRsojph+t3QqKNxTx0YyZlGB4MWKCIBuXyMNxM
aSYRmOihyG0QIrBLmGGtFHO7aZJThEMNfHwoB6IKRmzxp8qIqx9W2BXA75UE795z
IIBmOuV4846vbM9H+nYOz4tW3WIkaZT0vkKWnPMhrhTq/iP/8RjCCuweZafdTLcE
Oob2NZcU0QTViFxicoDtrZ/G5V6dLE51ecaWnRDmV5oPgymj+taSx66QBagFejan
tcnepNNt0tqyBD9xGcJGpyj50ojFO5cLo7bqDbzV7RSZ7Maxx3K9PHRJECIKhgvZ
6vThvt4Vc6S8M5pDCjCmxwe+HcugMSegqjVoXwOdEbCtJQldHQ1OV6bP4UOGBPFL
NdeD2hQkbvleXwn3FzoevlpZDO2TEYe0aeCGJHKNG1Z4e1DY7iFXNBVAAWoOMVQ6
oQYailM36HkCZXcn2W4tH86ZQVa4yfsmU2kn4bsGCcQflcjh7cH9SZmvfDjiizAU
fFfTkyXoG/qBWuKOtE9A5y2R3lG8VxLVcleydJraFNyba5fGlCvbbRJCJH9vbZnp
pN6S5R9GQJH4TDh35MP03NFKtq4eoI8GywVnrYMpP+vqwENaPcUfaXmXmOnHiiQy
Lz4+FQGKoS6S0Txoai73L2yblVUI8REMnmmVFiZUV/bepsIyv7qMLy98EdRg/QqN
RR0Px57eyr01uzer2NP3I2RZZirQx44RMX7WKLENja88Y0T8xMVp50rIUnV7YPnP
tgZ1k67i1dmcC+8FUgZX6wplmrJfQemc/fEwcIjcz8y8JM0W8iwI+r5wUq1y7y5P
dG05ZhwbrSiWJFxbhrFraedDISkWM7eiCyVzmhO4z164UK7AZ3+wLp8pjR3jGRgM
BxpZnGLeXWxROkAv7+mB16WnllPjObGgL4zIWB7jASv0axzN1BppwKx+lw8Mkli9
FkcLOJrW//yJcJFg8LBtEfV7lIB+5bez5JG982kyMzhG10mlwu8GQbu82H9dbxT0
1Wme/MiHyv+9Hbh2jqp8PSH3xHsqGQpFRY7HxSTRlM+Boj/LCTzWFDREtI6VRMst
0igR7aAk9ZNSfiGQYAGeSSGmBa5rAeKQSAZSIZFK2MYXJS5P6QCvMGlMJAXG96gz
5rzNwUxOapjPDkWeEJKCiiiwKnAaiBYUeNWQG+QY/MCZCbeD1V8EWZvmeprv1H+O
9EqxUak/C8uO/mS+Gv1Xw8pfATos3YjIbXr6YDMzvdU0Sd5GbAqhkN4eDmG4bLVY
SKmi00kUovLGTrSMVTywlV5WCYuy3zZ1eJSNC93pgeJarFapAlDTBzjb69a+d0GH
VkuTWW/oU9rZr17XA7A3nfLaVXvscDQBHb4/RRBUIcdacV8tCmNoQfIgD8ix1LzF
r2UpH/F4rcCR+px5uNpGVY5qza2hS+WwoOBUQ5kxUxlh/FvthtKdDhr0tNVocRM+
/SxtBv+bhCqZuUNGOh/tBIIDlZNTfGFnC1Ydl6z4x2L5+1+XlGEdVPTDI30zVcLM
nP+bfkLw8HHvkj/NSStJ5pfCJRaxpGmAaU4WQcC81ezRxn4VVfKyTy8npNLoS5uG
JjC0YO2IiImkLLykeo3MbcM1cMDXlqyz9ptw1swKQUkNtyLI3150ZYnu7eb79CN0
l57/hHT+GxTDVP0PYED+qQOTcb8hFFUNrW3c5DaAY7dygJG38CSNljKwJNvPu66O
BsqX0fI0yJivduIUKJKhOSnMOaL9t+cklVaq81+9XknaDCCpTsRQ63a0noTqAHn4
WpjI3OgAHyTn0PL/jG1KVwUtb/xtBWrMGVzuaV4ISPzxgtrntihmBVbOqyyMay6Z
uJVPCx2MsqTysqoRgoakZFWhDcB6qgSl9hI9EBublT98F5Wk5ms2JPq6YcRAE6ed
IZVtNVVKlgdl7cZU1zlBtrj8fV9Wj/wtaGAlt8EwmvwmGS8EGXVW86j8TNUNy3/1
7cZ4aLWxbEg1YBRatYiCxDtbPR7Mcm1o4b8fe7RP+fiNzCMMvkiRZM+Z1L5GWkos
el7ywQLCrU0MDr3nxokbhUEJnhgT8ixA3KtYUkX+pJxWJ1AxtuljJRnjjg84k8Rt
mLiB8GP8TWmTr5rcVH/TWG+71DojV7idFf/bOFoio6mb1TtHWmzJxoySRiGhdLDy
6QLVf9w/UaaKJXvUQZqO+BZR6VGvH20I67wd6hfD3fhfnF/FmITR5RQC3rPcqOmz
6mM16dJ2ZDhelFLhLGP72XMcWB3h7iwp9OwhK8/qxCoUPi+S03Rkk9BLI5u0G71o
HH420/BP5wPxlxuhhJ3qtKSxQnYa57tRvZHOKjEmVhEyx3/6t4xoT3wyS0DADR2L
pb939cniZ2QQI+bjIoLyxK3dgQM0NIhbh8Zp5vZPKiUbocAVQJQH6MCn2qWfJ/oM
rYHYltqggjGmPiWqHKLBPkkWitNL5VD0vuBwZ2Yhc4tl27W5jrWF1Vz+G78rnmMj
SQoZB+A3H04Zn1RXFkOx/oc2SdRYqoNUz/VgjOuoWyJtkGjr3ZcB4qsFh2gEoXsN
Nck3SBG1V8FwGMcunTztA1E0+or7/NwQhru73ggd1cZ1hx7zDeMZMiZEEgjfLElK
vOm6KmVlTc00zO/o6SFmegG8gEC4sQPsHDYRAEbblRH6A6YjwV4W4dTGGB7Sa6++
/siMho49/DjTndpIO3lS2CXcG0fSW2t2n1N2s1godHCYSfLu9qBLoCW0V/PwsVPI
x6i6yEYUSmn1JDSklA4LQFZRRKn5BXvlelQXdGwE1MkJZLJ4/gZzZpTj0Ghp/hf3
hYe0p1tczC3WRs/WwwrOjWLEci7EbZFVzsHhc68tOG0qiElB8AmiRNY7sDs4Xodb
FQeUSGvdEnbjWI8dUAxMEVd+t47fGxL9vo7jYEGCr6NWB/ks/Puwx/T+kWInOx3k
+m3+LJxyvAaX0YycS7AAxAbWLtucTG4MrpZidJloTJPf75EJ7s/JEtOFHwTd8kvN
GsFI6Iw0Vh0Xg9w4h8+nxT3L4+MEl2SO9IGXsHlyHAtr6pdZNj2EPnStCt94+lHq
4e01oduUkX6u3eQRfQHD9Ni5frISL8QF84PPoa0o//Ux3Bq1xrA4C5lDih0vmvc/
WCLsgyGeTiQvF9J0oLwi1YpZ+FEUTPq2C+9NfOYfxni76wNYCasvHDDJnSGxLqKd
+bjyZakUSXesmBE0Jq2FWWet8o44FJyUTxBZRvbtJeajnu6/0ezxAJ1JwxoY6VWK
pGbid3YPJhWEWraxfSpPEhDZJBxH/6Ln12DVHFMN1Cu/PzoImtCmysnx2QWrJUhB
AufE9hK2qwfEM3aTlZx0Fg==
`protect END_PROTECTED
