`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdqUP+UBPeKQnWEb2IQYb5+sBpqv9lU/ZIKImJEuNjMhu9SbAMSZ3U2gxecKo8C7
3LHQNc7Y7rawcQRMUDAUrltCp6qqNzXd/tZF3LsfNtSUDFDCnO0Cgqy5SlN3i2FN
YlccLwRUds0qlwK7TzmsiqmGjLHHvk2CR+zI8aRUO4TVnejyMXTEADHvcku541E0
wVz/RltLmpn8zMiSP38zagZQhgrdX7nGFphYB3e6fhmaC2RORufRHvUXpxgDGIzK
whbaXx1WX3CLj8iuW/QaJjmp3gzMWH/JUTzqjx+BIxPzDuwmiVIV7iFpCnFew0uB
LA3ISQa2uWtELHxCknqq6o3+wFPRjEfyOZAo9E2BpGG0yh9twrK0P03EHyZTtH+Z
h8Pkb7QeGUHmy0RlLK0sej9BJZdbMm/G3kcEFR4ttEE+uZdleVlvstQgnB0Iyeti
OKy3DqrBmzn0dOhyY4DJC2mwyVXopABsX2z4ArwUamGD6PRRf7BtLx1lTXMdQjgQ
/S5H4VSDrwdRgs+eqcqt9Evk262/IiysSmrXTYewOBFSfzgRcH2ZVGiVRmWbkRmf
MEfuWE/HP/a6TDwwjc++XITbyhepD4nr6p3NDD+9UxdqtTcgwO/n2mSfUKf8ITDD
KtXzc/ojE0Lx6xkxbEb1UZwc2RAys+HK2io1iREN8rPY4LxeBO+Qf072JP8EedK+
7C7YQn4+Hm8AxYA+DcwRRDxppN+96MZuxFmr8MbWrwLVS3+Cyiad4VpWX+iNqgI2
`protect END_PROTECTED
