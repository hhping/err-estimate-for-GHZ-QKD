`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qX1FVv4ssI+TMf54G1jc2WRfGBVDNAmx33nhgZXADCLOykr2+RDmv8j3WzWpEHWK
Z/6Xu6aiAzoOeg2mlHJXuaML3ouf05KVhY8BA3kc+YsUzTkh3v1D9lQI433OSUx4
ZrIdh8TPn0sY+fdGcElr3eIt3dCfKVjFsmb7V3GZKsbOJaGLKRYTC+wyg1JTUL6N
XaS93yIYYTZEl0ZPa5ciO2lCKKZD2GnbxKoEE1LvuDNHM1K6UDrFsWBy6/uLwZBp
6V3/ONOmVPW9NJjwtGpHlWK4hV2iNJKr3G0W2qSXwOquZrjrSgeCql90ugKIk0CS
xEwFZUIJpE4qIkFvTElC1onF9+IouCHJ0bSpGXfJXbZQd1xt+ba40Mn3GZ5lwWtt
CY/yt453g9y3EN97q6j5C6mScCdl51/zKOsdonGEZc/FulWQDMSA2ug10raX+RT6
o3MPJDpL1fpeowXIDH4i8IQeazpyGUde1a4viuxEgrzmU3FwWKcv89t96+bhwBjk
iIYPcFNbbZ9X8AyTg6SU1RUvIDTD9w2rZhNZLNLfXmH797JI99s2V8RvvepZmAeP
6jIpPxvSgbd7PF2dGXFK+6hHSfGXbLp85tJeNDtPjie6yWkrUCQ18nPv70ZLoW41
4x6gBFWkv2CpEQfjo8lxD2bvpzLtzkDZWo/t2joNm4CW5+Wrf3CeoE3clC+DdVOB
nQlXpFOvTx1NaaHKpQgxoOZ7aP4Ks3bkGj45gQM6FZLFUEk73KZZAZfWM+XQ2oeA
Ys7dWpTRl1px53IQkzbizg==
`protect END_PROTECTED
