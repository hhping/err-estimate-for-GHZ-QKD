`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTSmcp+KlkHggluY7Yje6EecyH1gk5D8kRqz0tFSIQUXzR0EXuQbyEbBD9IZmWW8
1dbU+zZ/90JD2dCkPkziyLIk5uTJIUF8vy3uKV7CLRuTUFLQouOjO9twiyLs0Zp2
VS7HhbKxIlJa2gEW1oTGmN0BoXDq5K5Je2JlyaBaCrkEkQPMa3cN9Z7QoFMt7cYW
d3+jw41MDYfww0AIf2psJa3+zvbE6nC7UtlA5vXuSHEVXa2D+xjAaqHfRmu/90hC
TZFVa34lty6/JDeODiMd2pODjFL8DEbvFSFZuXShN20Lx8vbzCrlf2RCCL2LKcYZ
h3l3Byw+vuzXZcHqIm10DcYa/xplbJgOj8ERgCWFp6kSja9/qTZZ8qupA4ZxGJqS
Ed+k8isllT/+39FNMhHtNElbLYiZLikRuAT/16F7BX+0bMHrP1AoW6+vDyupmfqH
i06KIX9zr0STPKA+imejlPgdrSuR5ssbC0Ej7lDjXqYJKr/aREvXJG2EQGVcHi3W
G0tTqeGa5ZPvwCSw0UBkqJf1RrvOIlFq2lU53F74xoegCU3KmSbDIF+CuXT6xPr8
JftKHx4x0nzLDCaL7mGWK+Q7+lwZE/OxNSPYCkwH7ISw9IXeknJRVfSojCoecFfo
ojqVGIlqGpdcCdM40Am2UhfgEaShcZlbomsZb68gDiPWM8PtxTv3wdarPxytSzGs
BA76mGfTvLBSHICRxHXcWM2ycbtt5ex8JbrP/it4vO7cbi4H3TsKrF3i+d2LOc8G
D0yaLOuI8Ko6Fpx9YlkQpEi8C+7wLfjyy9f7ItVPbPr5aEp/ssgw48PSt3dVoBDV
ayJGaIZgG+Q+GsF04j8TD7SkTWJFXLGEjzmwiZyKBLIIip1iCCT/mbXXDl9tmcE9
rLmO1cQ/2EK/WLtT9OWQz1lDYYMz91Wd/ZqIyjIqcLgzwJhXijPoM7k+1lYsD3jv
KhAuvm8O9B3YrT3FhYSM1m5kiFwJT115JA5qiduVwAcikQCCsjRfPuZ8QgTRRrRJ
dUikw3IC9lmHZaNm7b6fxqPnBAE1HXHDSbNyJIE4RMlJblGPdZdpWhl3/ETVqFHl
5whtmfDL46FeePiH5YLQXZZazQKNija6Lhj0OxeQhuOYizU3H+LiqtbZy45SN3hG
k0a5wJndUKgCD8QRcBi4kA5ZQ6QGser4VtHB1oUdPqhgEs+P64Y/8YnbjqF45OCh
IXSyQSeDvExQlGB3rPB4kZqUr3jcJdjEXaYc7ngYs1VIdiGQUhsPI3DrOqKqa7nr
bvJlDbIkZjioeiz0EVTVu/Mw8cJQe+bWzi3N2zR7/3Ah2c9GjUKUSZ8jvsplUmeb
zysbBHHZushqRtBC0wQ+cs2SLrbJb3kc+ddEHTfax4eJeuUhk0+cMdyFH9GHLv3U
24IaHZBpG/CdpA/8rDIuuBrNcZ6tc+a9vNtcLket+1iScRH+azd0G9jXltLNkQX1
SufMGyQ8n/wTjy3O4GTytShgKs118dBtB/5T3QWy3+CddMwHFUIdOuAAeN4fAJK4
ep6U8SEkW9bRyVspkEe1kL2ZMQQHsKAd5AEuKX+EtBn3a9QPJWrJIP2hK/WWdIHG
ez/bnYodPlmcndC0gsoVJJv1+v4u/I20HdY8UkQLInq6G9DVBK/MipBaDmDDIcHE
uaKxyeHAikxTHG8/ter2R3pWbSmSJIWiMieJAVTKowtmr73k5AZ97B4jrdXB+K8g
gyFo/hSeUZOdVTnyUAh30y52i8F8UlK9/T5HrHaN2OhetzMxuMiJ3ev5GvVe1+cE
/y0f+jAKeOor8MtCR6WuV8k/pPRXgbx/gllNKyWXpnTbw+beK7x/3jnb5Getb1gb
lAKetOvn2pqA03fp9gIax7Z6J0gUhEoS1TG/Dg+o2AClqzlJdIMePe4O3cwU/rkU
Fn2BVXFyod20ZGyaRbkGdlJ20ljc04xDFIoKPHV2xmGVM/g/z135DqGisT1jbNx4
Wdg5Pa+X5vQc2JZUv3e0l4O3ZOMpsltu7AB8eiemAVQo3oz1Bt+9HVW3DS3QJk9K
bhY2oqLidgR4MZ1mTKiG4uPvnuzi4WYcOhlxiUxTvqnZ2jUorz8GQQGyiGoG9id2
VTQOw71WpoHq0VqcDOvOmuM4+T1A/DIvl8Ri1PNuaO+bSKXGqE78rZYPZ+HLKivt
ZulJsxZ10hr1fpSGsJG2W+BCKpEqunVU75J8Sa+On5h3koEKeiyGQOVCF24jtIBK
0Y950Ny9N+hasVirUYgk9wCrj1dHkYcIMSc+MAdL6s/Pf7igj2SNfjAd7wtffSFl
brh1tWepKzBjHJ06ejv6WX/pDpBhjsK7MIsfYAuCUN1C9p4ctb8Qs/pEOHx0sS5Y
IVCF9C4WulL2l3KVRRRApj1gqpflEXRZ7IfZ7L+JTmU40tC+a2htUGDgxDWdMoa5
02N9sC8qEJ3rikUzmIQhXQSiBRV5KiDveAXjZ/6r7mGsDF/8DQ3JSQHRMSb6Sgq6
pwFCc9vDTHOcWvExq8Duo/oFSjgUeNTfFiQAnmvtxfigh4qhn4OfA27KYX7hUarS
D/lJOVYQd/fAxEm5nInJQSPhFT3dwrgdarQs5n6wPFC0Rt3EeduPhvIhyq8CyW3l
0zZlwBiFuGdUiXOLEWg7clb91aL5xSHTQ6knwIy3wVi8WLLuBS4UPh8jQfN6O/h6
DB8bfhjNKsF5gvwbnsOhNOcs1pNTRgY5j6boCwlRQTNADoylAavqtwPKlCouQ55R
68fdlSP75vWd0Juuda+IuD9e0nqVqHkb/fEsMwCMFNhATyQ4ao57F1UPpfL8rno0
3J+L7qlyT07bY5tvRKh+Z9Aufgb1WgzgEFDuV6QKL/6HvdnBItqRnAWNCVJK+FAR
e/+Emv/ZTEalF9uMbxKWgaoPCZXlgLc4hCFR12GcJVBqmQ3YkF4lkMQMtlDn2uxv
jnZ8iUBhQ5RPkattb+EzBaRCec6obyryHFOmaPP4bvDHb0GPSP+YH0jkDbAtMsaa
30pZnf0qaLwr2OS0XWH+iQIwzLCUNUGqj03clIGZN37akqChhvvxuutoy/MJTFQB
WFz9J+gjrO3SHTSGFjeAHHWQh6yGAfeAJj+d0KjEUm7VKVAyznLSzZ1KFX//K++V
Dg2/yBbLDg0TzfnHN3NeFjmfETGxzRReLq2C13dD28PzjITtemu0dyx2rywlWcDc
9ylc+yujYcyay0jKAUG1SrHzZ63wNXsJqr02fkwUTesJVjsq0hRF2y8Wcm29WFGP
NixBnnx5g+49+WT7mXoGgidY97VXkTi1CGg+0axxGj3HdhbQ5gHXwpFZt3ztI5H8
U3iQpr77Ac5WBmSLpopuWsKVUz5v8anUWWAi/gOKxKGP5xta4AhrXKft3bUhTyWQ
sIKchH3kXbf4/D0urAaXXCpy4IIQmzMN9LkcgNeIcyzjL1rMAMM4fcXuQVLryWH2
ljZY4EHT/2tEg5WRmgEDhD9u2wlxE+Dx8vZ3OvkUEWgHzwuYanonkLR/YsG48RmC
rPERECr3oU2w2C43z6rRCrZAHWT65jfX5yTbPmRNSm2XCcbByWeAzFph67/olfDh
1iyVPcYvqEm/RFRectolApLEXFYu+hhCHZqCYxcvgxsFxIE6CJ6igPq1Iyq4FXQe
zgZ4i+uXq6AU0ahvQ4I9mZxY76CluLUGceWo44jlf8S6gh0fqudjBoc7QQs9+3y+
9VMpVdCZd4nLdmXtkiI84wkDRUVsXg3r8ns2xpeWyOHwq4IHhx2/BGhmOshrUe5q
aVM0/9buS25ArurfcsVW2gFJwMeuWp03XOgYjEhR/NfsZhUo0/z+OQq6TBO+g0If
EZ+81uPGHboL6BX58SpeGeaaIBuOIHP98ATTEDQwMbv3Ec7aoJV3sAnLyMbTzIqv
LVh92lRcyCLlpizArzufIb0qGlxtk3EkkkT4GTVuoUV+8C9HGH2He59KZ9AOStyu
ymfLyNWZ+soAXuwTryRLCVXi/kYNhV3xFmpNXtarsykRPI4B5802/S8ZQ66dosfo
p4BTeyO4xuzXfh1TJi7v2sXpTUL8Exa1s9XQI0AQ2jS2caYgipzqKg3tfFrtMlO6
qEMGwbMri2M+UmL8YaanQGOHf9W8y23RhkaUf/hA3RvBBdbV2dBKBbtoiRQrO3h/
83/P8oxq+MKhX6lzRv4XGGOc7MMnPJVezjMvS06VNTpQK65gHKvyS49a5F9qwkgh
0gY6ochfyWDyQmCR74+aAfzPpcVSG8K436ixdE89ZkInvGHQIuT+jEDPNm5QdNhW
R20eXwBHB4/BDOMiD5UfgiyZmCLsTlcJ3htYTn8PnuEw17nROAZdE5eJqozUpWT1
iyhpyzRyQ/Rbhn/NXPisz1GKQkfzEduI2hWFp4igH1iultBNKu2AB2gl6yeG5+cb
3Ca8Gr4IwvVrxv0XgqgxSJdZK4YcUhzDUtMyMVTUMG2hIcPQ9IHIXkWPGeCkziAQ
YmnnKSXpNilHyPOcugKq8qgg6mD/IYPsKUwKfva1qI7BeLv5euOCPEakpfR8DF7z
zKnEfrFXLKsjpZfQKmzHR03s5soORgXpgatgpH4X9RhKERr+Tica4brJ4ibVsqPG
tbtSo2VRGAam1w62kdyRuQP6gD+AY7TbgkMAlpGmwk1dFyrDhcMjAA7NXAXEkEms
qZKxEIoSSffgnbiFPXfbI3M7f/6NaWcbQL4Ixr93ag3eHZNKRCXl3rWyg2/6eNCt
Y1Nd/5ig2lyfLEKHn/51vlMkbpo/DLvFjhGmaGbpXJrjkQfXP1D4uimrDHnLDcVY
cPN42glrQujBDGuHX8iu+2SsREVLJelGvGl1Sf+n1Ug3pv6cROaOzIVfrZRcd9FX
zE1LvxfW7wqc5ljSM6fLCBdBeh/h+2HG2RMKO3qFArtXTQFIVH4/Rt7KnWxwdtmP
8W5/sn/arcfPEYKf0q5cv24yZOoWYVx492WcAQrTMq++AYWEZBPUtGxpy+khqg5g
0GP8fnLFq1BQbewG1dLXTU6LtJEUrOa3ME81mL9+z26/VzeZ8hQ8QjVeuKpcHCMK
qkdJQzKFhLOAWZEkvGH4BWJL+jaUCFQchhUE/mSkpH11KDGHfceGNOza90iQxd/S
Gr+jnK0A1HJHI96pHxV+FpYZEPZMuUOphxi77fyRm5CCiJokIfhswyAtTj8hlz1c
9TTAK1w3wWkGSJ5eMvlPoeEyu1Plw9yfE4eKOsc3CGYaC28XTSSvYrw0FCdqso4N
ZS0GbvHriBySBPZqjRJo9fdMzmg9LgwYpje/XRrDysM9T4Iw2F8bzmb/7ygBA8ws
o+DgTFs9jYHlGiNOHVPXpqsvwKn5Ouy8AZ4K8B9wOL3imnhmnfTfRsAuY/WuDGXj
HNhvKD43TD7d39+0zUf1ILnSk8tXENkB631mqU8hDMk8ISdnjxexIpQ0e0VBB+x7
6iRWlpp0OVcFX2lb2H0IIDujxtNsHm0W7EF1frcbfJ0cQfc3bKxB619R+Tq5aMIE
az4U9kO0nmLM/8cTZ+wtJY3Gg1dy6955rVvgjrULYIi10vohhJS2bSi359U3BmDH
6KK+h9UWAsL0vHZ9864yG3bDehhtRtXTtg0oAdsAKM34i3Vk/3yyFdjOj1Zi02nk
+ZTE8LpdI23+ns4CWS2dqXr2JY4NJDyaumGVI7nISJDFfIc9aTTaueibUWMiSDb8
RjNeDnaRWoAWEG9Mvkb87jbWRPbLyNV013VUK7dBLlohX40MXjt5DT3sEAAwvU4q
ox5UkEVD4sUqjhU4XESJqfjcQY2ykQL7ML6LZ1dwQ0g86qDkEW0GhtBpPdLTdYDu
Mc57BlZtzO/UUrOLA6pUy1aSHV5y0dNM2NUuGazzRRBSyIa5Cd+WEHj+l736x7kP
Fyr7YyWfTrM79w0HBuft53jElAxm3CxfuFOXPVVqenAJr8OWtvvmkHLFQWXYxwvM
bU2dkQqdMvMOQk0NRthhmdmIOi710l4yVY+gmfw+EWEq32VAg8vZNH/YWQe81a/p
ClhCV78SOgAu6/VssctkgsKsiSFDcS3YQ3fYLGB22decWgJSuaHkxKkHw6XMjK1O
nVMxxxvDgyxoUG62/SQSxji1miuseFzRW5b61KIx89XjZOs3JOPEK7ycg0kaX/rw
x1juT58qQjYDuBGAWIxJNgPwy9cgbAoKRns00R1mNzrdafKZ7tEK5AgSc0mkguER
mUJoRLwUQQslr7ZW/cd2YVDHE0ZMUuXx44JH3yHWqmzW280LYoEhIhaO+u/lfGRN
jIu6w2qgJS5KjWZ0YdtvhA88QYZIpXyjd+nF7OlXjurm8NAzRgU2dAgzPp9SbRrR
IaF0dPio9NH2el17Fd8jGrUNxjVZYceai3+wDds1x3Jc/iF5Vsa/+H9Z+UcjJM0H
UHggxE8ncNzJVBpSCpO/rihixV1ARSf5Uidm2/k+tUDte85wFN8MI8+Y8W7SZ/EJ
Qk5MPneqEAWSHO8bgh0dDd7hQJvMc/aSNpNcwPG4pvEtWdfkMtSGeXqMVFpFOCW9
UUB1nJG9fCporDIjIlZ/pmOILwb8x/54Y6cfEg2DsXZZGnxkglul7/pkDX6ekjSG
py7g+zFCm0o7yNfa9+IPfqtd5s3C+211DuzXAq/0AG2HayjOcekpHd4NKi64w+HZ
m+hpfbXISddYRO4jYOv+7GnNV6U/jac7Q4NyGq4wSiQWJ+1TOnNRyXHxy+vgozMY
R4C4vX/9ic6OpPtPH7EPYUsijvSvbLtUnJOy16uPRMhJR4rJmi/FJg+dUd7piPdA
JWi0OhagxbXA28mwappqhqn26zBceOHYe14pKhHyS4HZYVZQE0V7ox2vqaSIbIw0
S0viRgHwEFLo7c/Lbu/d+9i9ykUfuo21i6I1myb+fy7zpPV8KU9RaBe7QzKSoGTz
5Pr7p26a50AIjujzTlHKSyKS0xNnGd7gVOccixfw69i3WiFP49JrO1uSkLZjwTL6
Ru12mVUWmPp/fMGwrHpukkmwL0VZZ+gdjkVeQ8duXp7pfsoch2eFeVBxDPkcgbfg
3U0kS/dVZppCCH2ojWunPDTq7zamko/oa85y4ZTUYFlH2LU18T1jMEuqC7fb5iih
U2wTUJ47/e0Se0s/4VkMqQuvlhVC/OluGhY57vjz1NGpyrLwffZqMo+OeVfMB3gR
Thy9Ft0FhNIHIPfehAvrhdeS0YyhSbf5lYfNn0CjizzTqUabP1pwG+9SckA1oIPr
1ZvvQ3AnNU3GaxaXETTqfXC4TrmptftcP5m5HCNB2MCowZB8a/y998Lgr9qFzBmh
/xV4j6VaIqzlIpAwIEqhV5gO1sdTB9rD/0crTaTBH5yp2a9sj0h6faoV1giSwjbG
s5bNplQISFx4cemaiirfN/664TydmbCQ+ppkKsM2TgUsPoKml9aaqTfzact0Tl+6
qbzJUKee1oT3JXU+TRIwFC3V+LnItJIIeF2GUwbFEI3P3c5Ud6Y8Tb0QTOrm5zS0
8YxuPl91flrRWxrcWjjjg5roCybx8U4JDGRDC1ldESRwrxvot+nEB5S/Ffsp/v+g
ibMgfknd3Wf9nCj7ghhIZ2xIG6n4tTmMVyrfiqia75rAOg7U7Qh7AcHRnRC8d2t9
bEmVEz7PS53rMcDiEC9xhVVO9HgTJKQlbiD7nhb9tzhq8XlGukzka9Wk3rdei05o
Y/RxYqIX5hNtVyM29vkodmpK5J8ckMsj6lJBUrQjyyMIUgo1U14YaH0BTNcDb8IV
G6wN+aO/mHSrlPfFSB67xmGI1ATKQdWC7dUuI0sn9rhmS1QspUnnJTxn8MCtejik
63NddXHQLJWuHe3pJh05q0jg0LQX7yB0caL1bdMX3zdVwLpqDKAf+sIVJOzfrLNb
n2mLRoGx2QOSIbsvfL5/UXZNKECBthnuaH1sZ0TMuoP71UEPrkCGJfniirU1jkvP
G7OQ8a6NKk8fWAnnp0N5dtrF8Dt+N1j5uWqYmu3yvvE0fxx41OCh0g8OszahqFBk
hUMQ5kuTa27LWtKuGn4itg36TyWblMy6vYqG9ezAInby1M5F6Ds9zCK1OB9VJLHl
25yHrUc5lc87NchPfNSxRean0RnmDwwO36i2ba9R8Apu1JHYcwC1PJwkytAEDk9H
IZJjRJD4Gur/E8FVrOeBeotlehLmhmdRAEe4etAjQpnVO1kjEO13l1TNpn/hdgyb
M3nlymSj9aFdmE1OVM2xJA9tPtLBRl1ngZzKlib69aWrY7vPE9kz7stBH5cUpGtW
ditJPw0dXErfYcOeY0fx6f9Rtkia2tIm8pZVw+k0ap0EnCZHtvBJ732GlFwLiCMV
aGjY9OgJ3UpKSF69VtB9quuf+j+TACHhiA6ZmO9akw2JQVM+IkASrCApsRVEQyyw
uWODpqqE3QSePNsHoSir3e4b9F3akEhhtuMPtWq+SkdzF7s6nkam68VeaUgHvL7m
wPnVdwgKHhzX/C0QoknFYxL1tXovZ0N3tDZ/cOEoIAHjYEEzOEM3q1RbThwCV6Sq
tI79hqD7vLt/Q4auYj0rDKzIDur6iTOsc1lxyYiFoSPaWDFon2rvCIe18E72vmwt
qnt81lcCiLG9LSxZCJo+eNvVhwoYXyZBb7HMUnyWgh/iTM9UrAQuZ7DyVPb1Fala
rF/xrrPPhIDGuKtWdxnmhKEkZKFa/saHtxyHKxbLvr20nYVnNCZ+/ltwLvKa309u
qB+U9xXsIvUiuwNyEl4zryFunf0jMjq6Fod0WQOJ3GDkmil7BKTg1q9N9IuP9/Zt
xvOgmsLhaeHxIAtgmCFaHRRAzcs3mlmNoE0xkDm1p+uCzXuUGgrSbm+YfND6kZRv
9XavM+efs6ymju82t5/C2p/eQ+bZvP9f4nNyk05jNGlKKanXcVL4UM9mTaa6HGhl
6mlVDL7BJocUd2skZueTfbBXATK+PSNB00tbA1Zj3jS/+0/wmcDCGEmSNlYvXA1q
5P0UKAcqZg3LZtDm/5a/WPqIf01C2fk4309FfjmBbHqv+QRI26dw0fkoot07ZOrw
lgmczls/Bx4xccBZ49Hxd8/cYB2eIFwu/cWnex8tbui3yMLqHVMbL0X6L+0JcrGx
A05sCjt2au7Wx77TM0t9U4Ht0jMJbxm/jL+4AK9CDQjjYtXsMwiWv5S24VANbqEp
1rcNO/LzOm/bdfX8AADw/VtHALLAQuTsL9kecV3P2OU2Eot4QRbkAxgVeoJ2Egaw
m25CuiHXuPn45nD8aQcyrdrIhOJj42BsIiDqZ1QvWEf3xzhKivjbQgxbfL41HCoB
9MoKHFpP66xP8sCWcoEZ0ZsWdtDqxpJZjVlysMV8ugvqQtrv3TYL0ZgJPiQVBqFj
XWYcGemAgNswZH1h+OOwg18dBvJGZGNJq/98GfiTFZ+AvqzK2xKvW/G4/Fx0g/DF
mwjr2BI74riYvSrAZwlStynygLZj4v190DNO/whSI2S/nJUz40oZsmXMaagZSofJ
7PiMd4QvT2ocEbLoavMP0CHCrxgiU4irSjVrX/QhpX+ibvpawgKcIqjqIii0rCi+
Ou5zqnXCYZwwjNl60kfXjqFlwrGWVuZ/o8mYb4h5d+GsKe1ZETgQV5YeQW8Tfv9Y
zo6FdJ5y1xp86k8iOKZiL89mhfqGU9mj6MSKOq0PIhQHeSV7wflsgPRGHx2+rR6F
ELL3qSyxOWoqS/XMeoyZiIREyYhFWlX56SdQ+cxUs5l0kZSQCpxdPhEF9AjKIQ1C
qQ+26fgT2Xn8LoqIzGvpexw++zuNTuHgJ0fs+ghNVD4pwcyXRB+J+JwCLnQBuw0u
JjPB952X+qTemzEjoE3w/C1tjTJHS8H+zjjBDpo4DFQjI++vsrCbk/TiR/793y24
d3qHMGVYMwiZhwukp8N7e3jjSPHxpr6VrawzXI30wH5TMTeCW13E+WF2gWHW/sc2
pD6RL2lEhJAJm6MoUKleGU9ibkmTgacjrLwMn1GR1bahsoxk7FuQUw3hJDuIqYum
BDfCduIRqPGIQSUF4eGJWuNETcXfdvtOKMDlmH7hUjEUbZvYxBGnZT4QnoDvgJK6
uKvmorsFP3AsgVjFDs657hpZRIjdCgwZF/7+uBC68cEqP64DphZ6zHrDlfaMi558
XOSYNO2A5TE/8UB3Tmu4D8lULNCalL2GXL9giPURupc9XgdPtPfvCtimoNW0Y5uN
o6VetOjGGHkuSrePte9Ql6bMzknDcKkJraxJvax0CN9BQWCE2cSj0TL5O4wNRq5O
ifRsI8VkDRLAnmGQbARrca52+ap8Y4P780rDlbgYDIwpxupks7FbO4dEN/rxtzEs
zEndNH1m55zoW0RSBKowa/Hwo32qySRrYSCtgy1QF3vvxse9RNsW3NIuQRdQM8O+
IJ4kLWhsgLAKstDi9E/OdaFN5lOzFWDrRtTcoOjZyBWj2nVL5jz1fEmFuNhGfeHQ
vNejOkwgR/Z9TTGXt9BTe8DWiQWGosekVjEg4vLDQne+EEUThQWzyqEm86Loda7E
H/mHLk/Vvr7uCpNYmZgDd5Cj6tAjNd1os4QtFFT0t22BQ+OGVzxDUgVPLb+05XDs
dMsjbYpejqDT0fRVQPd8nk3MPUBBqlBtpwYakSM/ucWU2vlECS6irp+wjY/mQrCO
jnYF1ZeCLVp8Otw2UZU4ySw4Go141c/qi47mBOLUgPA9qteFLJiXHPXjY1mdaVzx
/UrvRypvpHIjdE9pNKoY8GUIWztmxkib0pvTN5EH8Lid84gk/kAATpdJyQM0jBzj
ja15xtk8zVE2pehJ1UePBWajJbSkl8MPiuFgdV0++G9sRWrscLBkRUWCEzU0wAcK
f2XAsVX2ejUaB/+78X2WbI0NAic2cEj0BHEhOz9IBqrVdxAnaMOkqq8RzbEROaGL
mFG/XS6zvB8kbB7abh/EZ4K7yJWVqjl14G5Vm7tMKaG8CxBqkTFwN4ZUIOSzXou8
lP2dzJfTuBTnPvtatNjZ/TOXOeNARBxWm8sC1p4nXIHXHRLYM+d2IsdO14PuTk30
9frg5YsZfZJmz6tRZUBoSs+JgCvcuxAh56rPRR+1zQ6eFkdaLbGhespIeXW2o9sE
l+jjDOAyFgiUrtsJoU7DGEMddy7Fu7r9nYs9Uv0GkIicCzOv6o1d3gY7pw59UkQc
Eh0GeSwsthSlZ8l8A3jihDt4/cpBPvqqUrDcYkygNlQvjnxvn8yLojBcnBKDvXS5
ECmhyXjMBdy2oybVgfdZVnKYR0MAnteiqO59fpra0fFjmAxLrh6oxwEpdR4/a1oW
We9gAmg97z8qc9/axCzUjFrq4eiYD+vp1JBTFE69KRA5QSZMANZsego6DDoIVlBR
aVkrRAvWiDeJK5DL87kCJznc80MMzSMQFBVD23GMylFcLZ6ZXEWbYUybloxaMa2n
7Qug8mPOrv8xbvhyMPJPkErHDqlcLnxH5wnCK7JBD/qSkO2dzugTDDtOrt3G86Ko
abRrEiOpFwMGgragbSRBDpz6ty4tOh5UpdCKOuKoHU/7Hxhh7u5pxKDzub2swXSD
WMDKm/b3jQd4XmPAW/NP73cMrydo4Y3Wj18zU666NT2j/CCFliVYj/k/ZHDRE+m/
kjO0t2nJFkJfxBfCV1SYA+A1GGeNAREowrfZzFFdLlBdIjg3TKXoOSNPfPPJSC+p
pU68dpTSNbdCIoc6Ys4awCxhVs+wHMI9DAvXwTO/rPPoXZ96pu0+HfQbt4ClNlF5
6d0JERSH5FDhhOsKpChTunvpzUyIGG0iL+LxSigB8BhdR9jtQ1QB7IeHr+2MOyrX
2OfSFb/eVH5fJa2eE3JL1FZ1B84gSTetIqVCbjO5jrfJiHjwhLzf67JXJG2EyEjB
ChgaBr81MeyB6rjOznr0zcms/f4rbZAO7ko3PeVgjUTLOCbm1Ne04MUy6JGMtAmC
/wYCIMdHOqaDeszdrpmq4h6ltpQB7wH8XF9wJAHuP09+syBXvKddgLUlF7o2MAg9
SulUElqbb6U/KXG6h/jUz9DmeJXUYtQH3Q8djdhX+Xca0O0EpOWy+nhdmp3JcQBz
lSnVwau8xH0G0HMBzYp6cMc+dgSa2NyiPXR7Fayf5kguDPsEsK5Zu452cS/X8SI1
QomcKkTTb7n0Q8vkmxBVl5Ks1B3yqDNrhe3BK/9SZnQvm26t2pPUrOiwclCqqkpv
2nQk2Avolzoqz7p0jm/SNNc6ZWpuKBOg8XLMHL85ukAca+BXhAxafDWfy/apJxSv
XqyZ8QuJAkrjdVG54GUtZpOuXNdhl6V6+22P1HAR7Zwo2fi4wrUBOe4ZPoYugpqO
p7dwnkC8ruGk2VpSNb9Vfu/BvEkwpkiowxAOyPuUV1zCC509JeqCfYpnOiZuR2Il
U2ImRaza24nkY+ER2E4aIzU74ypSVsTSnsAKZVXUHzawbPOZX0uX/VJQh7JMvV5o
39vM+iK1ZyMYovuJ5WxvQoSPw7kzUbHfibUKjUjKShSTABgFMJOd/ksbeGhWZemH
RAWcPuHKUt9xiUaAkRX4ogT1Gia8gIW41U6ndyu65ZG/6DdiIULMF5s2dCHFHq47
KscWQRx9+rKTZtRGzh+AZaAXNEBxGTSnSQi21ulzdjds3+/H5n66gfg4414X5ToO
hms6PNBlDovkY58gExWVer0AD+Hufx01OkZwcHly1bX4CxS/B9+d2f2PfKGmxYe1
09dtm4ZwQXUfKKw/ndc4qRv4Td82a/s3uYN99jjdOAD2mBIHtVc+waY6QTyHlxlU
IMPc1ZmimTMlXQ38cJbmawC5mP2rkLtr8bhHNhZ4OLAqK7SFEo6LaC1DhkDnOrqF
jZHfl0eHRQtw9Fbeyd9VlzxRVYKfdfnq5b4YIkLYrzzGkJY7EujpFBseRWhSvbkP
s4NRzpo4KAP0f/xpnu6Z2dP7HQDvrf3uHQJEUdB18WxpFCmHyQX2rKsKVrc5XrKh
f24DRxgqGm4t30HJZEFGPaiJN8imuCjOiOhRjVTRm1bQMdzs/Rg4/n7bZpBuTBh0
W9B5B7F+sOuOk1IyN92FIuMQEIS7Ys5JBOHlU/VCoa2iIJxd1A9ZwA2BiRNtCfCA
+yLYNth0zz+w7tzW70vq1r9GOnH9LylLvcrCPQx+Xj1Yp6a6KyrX10EH408gLGnq
WCssSpO71PtJZqUwiPvMWuViQ7NoNhHWaaW5BVXQA2fs4Jx2DhcU+k0Qet1Ujlnc
mCpTvOPtIvrDa2JqYB3aVO/xGcr3ruYLCe9MRksnd1esALXdrZ586n2rszZgsa3R
iY7f8gQgRan+aUWQgCvtnpsEFAbtSFRg7IyH2qU5D6pL9mtOxGgvT1XOGdJYYiGw
t763fY7oAypN09CCcw7hEH3ObHF1V5+8SX7qdTN0a7UswctOpdcc1jUoFkAQan5W
uOvdk3ai0I/un7SNglJr3mhYhhXGUcmIdetmqJjA7RQ37pd/2JpORAUWvBxj3NTd
gtoU2wCLCwOtY9YoGo0GLi038nsraj27hbo50sj/wRdfm07heEKUxBp163l7c/HW
z0cb7tPpmF2vh5wTM1Q/zC10xv0sYcWZGLYxnaBRN5g/bC0z1kUgQ4M+EfN0TmWk
hKCmP6ThnXzYKIL22GdwudKwVznZN99uKoYf6WVlOrRyTBy1EXCe7RA1cY7FzUzF
1ZdTV0Nkhs2zfcyFQdgaVZk7DSIQOQF7Kq7l467J9gmTAuKgb9a9Z56bB0u+ZVO8
7/e02WAv1J+12JAGdNUOj9BgUD6MDFR9/Ub1QPlky2MWTQ6Z3NUabTdWSZEFdVg7
HyM2QnHdlxmQjGqB038R+HWQt47LoNDnmvjSbzlsT/oW+y+EgDap0hiCDrhHM0+6
cIZrVJRQDfAz4ylZ4TYO64nrd7MCMTg+xQcFCWR0JWikWxGYvnejQjZ8493I21WG
yW5UqkVqz7fPCR4SJeWtQj5HNM1RSwfIuPUWA1+6Co8r/EwVYr/Ce/dXwz2LHMW/
E2EoNdChr6dFoVL9WBWjZDn+EFS7VWXm2DfZCpoHu5A4oK76O5ff5Lj3S5tqR6iV
fWJ+Pf+Pdn7MlgpYsivzza0cxj9eDm75vqtd+Nfk8VZptR6WMlkkWF0Nei11Yo9x
nYrI9MTkg6HWhw5Sv1cPDOzxIG9Zk8oO+9SueKDJQonqXb+VKL2pUBBBhr7A/3Ml
FDAAGrBPEW08ia3q43T449tg+g+S6vwaCJNfK5L74oP98rq3Ik87oxWIH7m8Fk8a
rJ+kk1h5OqdlBPWHEmpWVjPoVBwW/XLjaYQAPkQzd6s4Zj+fVvAHTJ3h3J0ltW7q
9B3wUY/P1H58y8jfNurUQROECv4d+GGNWEhBQiqXEbrUyMPXvql91aWP9dD2TWH8
Q/G2509e/Y34MQ20T9GxUFBeXwUVRRh5wHTSB8Uq29NqAIxjJ/xlxtIcHMflrwWI
Uzq/ikEiEmLN7myqmNxWdIuRyjFZYl6g1s2ZsAuc+orJAxKsxsHZGHX84JsHkUtc
kBtOetRfciEOCDmwfKyPxhe2wsmGIslqgClTnEWNWoFI0bNnbDZlenHxhVbYSVf/
3POt602nRkaSJkYaK+Nh6NtJN0AIhcdB7PTDzBFjUSes6CKC5Lg2Hf1qYwlEpEN0
hgmR66KSwG8yyh746d7hbPRYDo2vZ5+bnJ7jbUhCZ+9AlXNKLmU13kJoF+6GpWVP
H2jcNrFl2801YpUt6y4udIWRihM3iM3jZB3Zqx7f/szu/0YfSMhWGyX6xqoIoxWz
XpRkLKZghXaWUNCxslgtCxNnQwJ4pMuWJU4ZQHY64853gy2aDzxrgSXkJFvn0hd1
+mxc/XLp0SaXta4bdXlsa4bBn0FHhnDUxx3+u6YQINyCA1wxh/HL2UjG/1hMonpT
k5+t9BOjN8S9NE6BqeD6auxy3WjMjdfSkGtHyTtcs2EHx5g7qQCPmJjzud1i8yYs
UuH34Hn6gEKeOU+yrcs0Mu7+kcjcm6tzoH/Sq9xCkBtlbqvoctHL8mvcND5Vw9np
KtGqnj5s7ALQp0KZQLQC0Wt2FAiWwCwP05CVaBBQIf4TXcQVA48+det3jJpUZWVd
BHTMnGvpE6AVPIi0dp2K2S7ZKcoRQZXTnpYVPPJz4Xw1JcPiQctTpISRhj644um7
/8Vu0p+EGVx0YOWU5+7IT74v25uGouF+3cwnYOL3L4PslxQBchsbx6/eEd/LzWww
IPA6cV/f5HntkrUU9Gh9F5vFciLq03vACVMdSC0yC4RkgID3jLotUsWUEtcpMSKm
pT9J6vW1iv1RuP85sf1dWKmloIcH8CMsZkgHjNxBmkmqqDhyevPLGc8oM7PXPwWB
iR0D/WvJsO0cxQ6UUv0ZyhvNZZ1N6Ts+i8QvcSclHza+F+32ZJNVt+lgf76IRty5
wnepWj5Kum/PI6PkqEnfnjyX+aGcbQEvxGcX5UCHeiS9n/AhmupBl3PjWneOipkT
RD2zJLMYuYwNBZBe32t7I8sG0/ezf3JGqxFjB+YT2HGR+IgsG0yOkW/KL2NUag4t
v0DcJoR8ceUkDyqwxyq/9DU9mbVcfV1epcJKNUXGacLh36g64gpUmjvE+XaGVqT6
ejgwAhUpjj0L+Pp2ndWdAvIboH6hSX/KbulVSYnVbVsTOnTmJDuQxCpn+e5OIFf8
rg0Yzan5Qlak3YB/NYOAQ2aioTZDBpt1LLVczGrjhE0epKuWhaySMHhmtBw++eg0
U4SWdo6A1qEIN1o/HAdDWXq8Hlb4cd8GseRaYQBRy4PH147fVCa+Qm9T/nWG/Iws
ovGqdzN8g8bF8VqWbTHRBcLhAkHzbmhF6tgws6sGFHc+9fdnRPhpTie1rGWr4L7L
chZnT5YAc0kgZBg1llhXJJKPqRw1GI7PuOD5W9dOMZdgp5DUqemufSankqeMOKDl
2ymThjYmfZQlObKlHuNEuu4Q3jwjnorR/4u5wiSBD8t5GmlE2qr0CSF+LXaNFjnh
t7dsqgwVeNBzDtAS9ch4uHVvNgRYwPKqiu2Z1QDrv5kbzqKWEigD66EnBcMEeRcR
SaSa513WdtzOdKBBwHeXAa8U0On0Tv9CXXFApeFWdK4pqN+p7WwAejjN2rj3IV3g
0ihMtOjEU4rvMfiyvjxRkjR1Z/x9kFfCdt3DvQq400/giqmDYTN0OuveBu93ja4K
OiQ9qzG29LYSUE3A31rAvMTxZxdfwgPSwr7yTzDSNd4GlWKPhxQje7j3HHfrl9DS
vZmfBRCEhJXqEZlpCjI7gdge05+6jF+jQSs12DKUaQcKM/glkHXicUHrGYofXHq/
VedamL0M5+0nR5q+6Y4GoytgvnY8//K3vX2dZJk0gRuVHz0QMf54jXVOmTSShLqU
mhSnXZqZ1ufOQ1FO7z3CNpFursEubvhomHNH/9osUZ9mEerWyL80CE6OWCLhQncu
6tw/VqlgQ9ZodKCrO1CRnZoPyu+IZLGJ6Z65Ny6hGjR9vDm06c01f+kykrSE8igb
PPRnbKTa7wRuo5aNjCv4k9AzMbx/eNWLxixm/AEBE7HbzU4cW+095rTKWud3HEe7
O2O5ABOjtF5GN4S0tnvqi5UZ7F+dnUQlse5+Ogdug8yrNqPgElgW5DVJzncKFPjo
AXRsjcmcSOxNy3Su5P6wWYISbazudZ86Wa0IbEvvm1AlQAx7f3wruvxvFgV4yvaR
3uaX5FdZoy3l4x5SIrJnRSjhN0L9xRnZ4DHyjPVl2CT7DWg6TygTSrvCsfZgfALS
VM4SQA0ZrrZBAQBvuSkiTEQIJv1JxolVERa+w/A/goo4MPu4x6Ssxl28ZPAJNZv3
SsDe8i9T8vniyI7k0/zAH6gPhEgmYQeU8Ihjo37E/Xp97z1OmgorRCCSUA8E4ejN
VPu9wap2HN1JalPI4dPZldjB9zTjBE7eTohG4dxQKU3gEDMYckapRAe1sEktGGMB
NGgOf+x4nyAyXI9zP6nAbeSGna8RrWsUL/wvQt0x5bD788jZv6GqqupxbxWaXTKU
sQde99gR64lhvwN1fcs2AMEUBWLJzL4MslVAzHu5Oj8pW1zJPmmIqZJDcRxM/beh
QmrgYS+4RojNnltQQyI+G9ZsP0A/JMnmCdcrUFYVdmZ+w2iEVhxxceRiVtq5beot
TfuPpTt6I8P2Mk5MR09qVr247lYraBzjZZ3/nVTNppcLMSUF7QqqcwkI1+cTUlMj
5supc1PnMlHpfN+Rm/59Jy5qh0Cur7JpXlP/9v+mCv4E7D24HHvK6TXmbiTfwK3r
Hq6pHhSLL8I5TKQ/dYhmb9I1sF0zPDHL2e5NngpxvF0TN2HqQ9vpPo5MWTYKIGDG
Sws7ZpnAiIDkZ7pJ0HDDbWZb68jlURFzyV+jU+JoXwmFKyRiol9ADtaIFEkA21jj
4INr0HdxZcczeiVkcinzDRpND+KfwzGh8OJQ8uZq5Ut+4P/NtcUkqZEcYfD5t61e
LN+MWwOt76MRZrorBrLP26S0jimOiC3AXIIJgPmAgMs/eHbaglKZgsWO1r1KgSBp
mLKixQuodNIkg7caseYRPb77kJ+96AsiAR6eRj43pbCEDyBLr16JGt2rLREqjK5E
7n9a9wIiCS6jzVvag2WWNUaOgXaXO+gTlTL9eNagSyBbsD0rhk7QVZbNmf+sgcOk
hVczk4EQ3Yo98agT3z6dln7Xh4UsR/bK7fYYcflC0kqJEpNxLtmuhWuiZZszaztE
RZ8TDb6hMOHQJe3qgXw5R4fYmT2OKAM50xrTaiTPeahbdKQHb3P0+qHNiQPL3LdF
2p2K8MdYvphiOy+0VN93Ku0Mw60hGfbgbPaP7q/XUNp4Ex8dkVt73IpdfBCX+rIE
TuJlsbUt8q/S9Afu4Kxo29jWGfeZ42PonGuy6PuHvo3QMJtQsMFuhO5EuAIRcqPe
fhVqZ3fLFnonLpUj1b7dBjYlfyJslpjCDrtpF42Brfo/erOnCpNyiUnJ3kH1ce9f
vvnUmGOrA49XGgkj+SNRgpmuuvmfbYCHnqBs84jZzQQVNw3MDDTRGKZbjQUYa3VX
fyykiBzR8ZcW2ZCRc/3wMpFZoZjQSuHGF/uvNgsGoFYjgIOQFuKTxH4BJEA6Jv0C
D6unILoeuy2O5mvFrJiNwFR4ohcHgIB7vHOp9eT9Y2cm2HT19tXtHwRIcDCz51zN
79j7p2Otl3P7Q/bwtI92u+VCAPFw9wqpHSv2LMjt6cX6GNMB0WkxgWWorNs3rkxY
N61JTm59viNBC9HEv0/3Kob1Xn8q25etP7+RW8ZzLBeYc5OBzctMMrLi6KljE+AV
qib4GjE8kZPYHW21MGarnb9MBDaNuwafGT91vsdCO6cXkZp0t3DQcwDIm7nTX6K0
vJac3qlF4GKTlXK5dsa8pczW2EutfaqmDf+Z6r2omxoUHs4zDYTFS4XLqkyM8C50
L8hJef1rM66H1k2PivBqfzlqp/LiHwJMI7oUGeIBavT6Cpol3ZoDFPorpTkeMeyI
Wr8+pv8fduOT3pgZgpOoF4q2JmaTrexrri+J3YAUUR3D6VdvlGMvD2LM3EqE3vQD
SwG2HyuOkzEc5G0QqtGfalCqSkHIwWniJla0WAPFYurq6d7ImBK9IFd0kIdNqsOf
7mJsLBGqrvDiLigJoAdAKYSd2SeTNOxNispujytO+zBeIDzJ8uNsUYk+qIt47RyF
Iz8dEN4VDQGdHeCPDJVklEFmNy8GFL5PoDKbzZOOdH7z8v+v+2koE6sHHxAppg8Q
GVuX9PEkYcfrdggq2cixAuS8CKNzPxQxZOmlpnUwaZenXPlIg3CYTHMvzWleHTM6
IJr2x8BdMDXLVPmVnJMKCCxz6YuxymCW//QjedNMOYhCdd8pwiBx9wU217IqC57M
H8kA7gXO47Trls56Y9K3qkb7aPP807blQuJRGVld9ScQjJUYmop/2JbADzHpP4ru
4jWMO5+AjoQCUSPaJkXvpfjNwm3u0mskpDdOnXyi4Zth86rp1UVIGehwE6TmteZm
vm8T/8y0n8C0z19+E9i0xCqZoUXGM34X0b5/zgOm97jdWTcgOfaztSZ14T9tH55G
r7tkm3kegk724veenDrigl25PUBxzdDXiaz5nGAmbnHwp9FetBBpNO+KFAMKbDj1
tQBcO0hHvh8jalEz9VL9TnROMxMblZGBqCtrr5UcHsy9TWyUG9kFp+Jkzt8cpbBf
uIlD0AJG0wbIKFPTTcCA73Y3ckIpQJpLVFPDueb1TQf2TWO93HOCM/GTn3JQgTmn
FsAh4afdwVtsVUnsvDQh+2PYYwEW44EezEPCw8aFAPNN4B/IXLlDOuUyF/sGXOTr
DXYpdDMuKBhDv1+eeo5S4hCVjmDcAL+5V5p0yvTEQpZkCC6cF3S1gpHpAsLDj4pD
YGuRjGBmJfO67uj9WKZTMQg2M+PqUOcK88pAvPClOgsZz4XxaGnlaYbiBBPrDaVR
QidQi7hfKAIcD9AG1hgZnCgyKaFNFVtHiB3fghTMG2Spwohb7UtvP6asMlv7qO+d
5rGfQS7ECKuiO+WqVvJs5f7UJ8uL+Sqa7ZDbL7CibLz5MVOIg+egURpy99J220HV
lNSsXiVd0C8tFkZPFc66/9g++ksDrRdAdejF2B64I5tiFTMHzlEep7KArrsxlo/s
RRhFmMF8gqXSHVT7fBLu0Bs672QIp7K+6/wQfrFw2lUamuMLU8YxRUgogyht8GZH
7N8rKfh00l0cajeza9e8CFD2neikojr0iZJ8vssaccwt7QXarZeXxxFk+/Byn79m
htJ5ATm010da3vLOoBG+YcYBFZpNhoDRLG7Cm6zCG/livENGuC3VJcvXxHFnPUo2
iu+3JtTyCG7OGGUzq/jWZkh7PtDvGBSCVSY/cX9KVr4vMviA5yqhlNlPp9GxezLI
kUUZ33ATxQy6An0CkKnuoPX4Zy12rZ1jbon9dO3AKYzHzyjL4SszEeF9clNL1f0M
sN5be3bW7ldCAwbnHMvoAfK9efChjp8CdVO7Sc/vEkBRY4TAGoL9PG7yzcBPQg8G
TSr4VUvWYaLT97l8KwuRANqZNB14KrV9yudUEXOYDt7XoIP8eHFyZ94yfcuOcLSG
f75I0O+RrEUjS+OJX3AcFwxryUdzNCY4Hae2zDo3bT9kl0102P2m5Lj1vnBXnFpN
Fi2MXiVyvh0aZiMxH2/iDqDINrGhek+8Sy3iqIfWK9x1Qbm7ZeZMy+znwpHd8+AG
1C0AZaNSiTUzAlF2SNncaBILfmURvGCgPQSDghr6BzARZrk5v+ivwkTQU0QPL0cf
cEZ4sRF0fDR9JuRGzvDl18Cz91xTMEn7K5llFxEts2FQX4RKx6vBQX7GLcNoth7R
V+QorPy5IvccYOVLtVJaYlBZwnMNkxlmbS4swUDbMDcwNQxbq/xqRiWTuUVVbhii
K78TdcxhL79BP5W4TOfzbTQp0T5FfGffpbimhERg/L6O5R+1LAHO6Xjx61yh5iyQ
XvO6xCjlnQzaqMSZXCHtQLh0XpFp2Bifee6P5IkXfvsHBmGgN5JQ7kX+N+zSIpd1
tt+gscTDdWJG5MzhD4uKp4RdbDnc1LwHMXZXk56NcWzRgD7ZJi0Vx8emdZ6f4HUv
`protect END_PROTECTED
