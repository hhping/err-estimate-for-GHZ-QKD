`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWK6jRFB5GXyDTz84gUOMJzqBu1Qqr05I86MVjdDZ0ivqXzGSqCHiH5iyIJJZkro
TfZSqJqPgGfigBxxwmxS93haxWlWPLVifgvkShN2TXz8jEFHWiBUJNwgSunMlZVf
XioE7z5oKu9EqVkUaL9Ogo2ak8F91c1uP8C2UVtn1gAmM4wp8fTkGhbbe/ZjY8b0
jE2XeHNVoDBXA5fh6bWiO5pZp5vpXLM4M/GW3HKb3BLcNi7enmZSGO5pLm6m49Kq
55Rznj4FOlTthaQ4JwQ/lSeWBT9up61i9mzjJ7y1kzZSlrF9i4Gfv1W9VJq3IGMq
Txn+h+ASyoBb/e52tfkFf1x6rGbymx98mtikX9HqBhKlz4KzfQV0d8CPl24tGRmd
fUBU1bYZN0A9EGQ4omEZwMY+xG0VLCmolsDDLF13LcoqYjxCB3lorpxfR++QbALy
GfZ2MoTXfBbuB4SnIkPHMrDavwVpvkyRDLgChy1RC7Q5IklvxLz7b3Oc6lg8TtEU
qcW+To+TIhbrCuyl9iHPik0SwWgd1zDS2NDaysnTh6dKYOb70Iqm3bdKdCHJE8Aa
lAA+/HLm602OVVl4ckl8qw4c2Ap8mf9Z5PPf/+4Wt+g7WaDupTqQA6QSoHBW43Qv
tuoYxKW9iSdjJZ+lZnX+g9J/txE4Ohbb27iFMbbT9jVO2Hoj0B7Nl8tnnMfQ5lHr
dYPJmYwWFBXQmDGthVnwzyzBUM10QXsd8miShJeqPwj3pCe54jXs/6bIFvoSvFIv
1InFbz2ZxHRVq7z9B0wcviMRWWee1SX4CPNXAvVNyDIw14bi5ZtyHxmpzrTtLOcU
6Ggf85IaNMnWZz22RneF8wE5SmRvsrEXT1U/tKyH/ccdidNfaR2lcsLRsPlswIjz
AAJCKy308EMzcLz49KZPvV5vF0MkSmXn46m/R1Ei+k4ysSGB5JhrRMG4/GtB5sVZ
moonEOQG3g8SePZB3HvZaQigrZD3rxpzSgd3/Zt0FmAcFsGTg/Pju+q38huxvf0H
AKvfSKWDIYbjjm6zJYw0VTb4EK4DE+T3kS3feZj44vP6OJzy7RmntfSOw6K2aO2S
W78q3q9du2npfeubSXt8sL190EVscJedwA/o37NGPv/IxXSz3hRTiloP4UThEX9d
cBPYJ5eWd2C5EpJ+tfJXTvtxoCwcpHPFd+f+SZ5YCblHf1dty9xLO4/mTovw448y
XPIEHvmTO/Gz+xrUUg1J8bgyGrEac7sKLykpMwUm+41YF3Y3c8KUZsIf/9a3knCS
5Tk6K4mp7Q9qCNmw7i38COuCgGySE29SHqhRcBhSRq0nij+HW6dJ07sfBiL/Iw6e
naIPSkHJlFGng39BvRLfUe+F4pokjf8vj9t5mv6rDUW7LwHx2DxE4IktoCvpZfYh
o1xGkqheIK1sIC0sJOk/RhE4sU2LWvjvm2Q/wQDiMgg+AiYPdO3lnc/O5MLU5QH0
1zuS1XbYA8HHMeKDTJLzYw0+nT170gJvGerpOg8PawMV1ZbteioUMDuq0jxYOAjD
j2DAFI8Cs3C1kVpJxy/VDrJSAtltzIdR1WEfnI2TOXpZDdy8iwdsn6FXKSkdmXUQ
WmZkeP6mt9yJQ4ApFUcyACvmY3+VHmQEyM3OBklHFH8UoYNBdU4RSk83hHwF8qHP
VNH8+0k/rN1Dl5CCqR+UDbd76u4Gp0bR0ZMOW7NVngz7wZWsxyyRSMgk6bUB3bn4
ZtW9AIMV4AtpBnRaF8pOKpnoVzjOyiKqc+uc2wYB5SgEGLdtq3cmihXNIv8MCX4Q
v19cmGzd4RQQOLRYt7eSqBaKfhVI5ee7mC4E+sb5QNCLTkqRzt6jSJrh9484XzI+
Qu+adYJl4eM2dCmzEsSGYHbZ0UXej1L0YoZn6UZHd3GIgMyHQC2ERqdM8hRp7aWT
RgB8JEcaOGh59piVTJ2F6nwz7rO/IRXwxtPcB5hQTX/oSrprBRwpksk1H7ONOkFF
DGLtajHXe7ZKU4OIDPdXxNCKBDw6dBzaruk9PHNc0664TvZx1QkP4/w3UAk4C6Bw
jg3Z6penNCZFAFwAf+Xh3RqlK7B5qktSJYAPUvhaZnOycc4DZ3DDbRUFEacekzo3
b0w2iTRPVsHqr1eTkycvSTFSSJPy6xaGueW1uTzrCR8W6S8HThCt0qaGou0oBapi
5R96C/lGWdh2iTUspxnjP9z52qNJni2zzuE/Mzp9XHVHKSuhzVCJNkAPT4chPPXC
D2RnRmHXOPKrr33kQ2hT4BYiAzi0igBP1wPincIhq40RiWxijwwoDSKr0yajtzy0
f5WY/DFWvlx+SWd3rmPwqiK7kb2NSrKuhj4E1Gzuvsm2R8zuQzYBkp/7M4XRl3xU
HoAI+cgsXHRhREScyviDrpZzAAKpj1KPHsWAh4JYmyUWL93XpLB1D/R91aHTyy78
XoxOxH+xd+GrGphMXq0/WENnn7BKjVMEZBY9d7grAuYDbBYMu11UA/91j2AOAF7z
cRhU4FocyJxuuBJT54gq3GuIWlJeqUYmKbriP/2ZGyk=
`protect END_PROTECTED
