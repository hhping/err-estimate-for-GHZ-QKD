`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+WWuEK4kbeVQTgbu8D/PIeP5qKXiJ8QK6k2AZa7VCE3d6Kjy7pZgU+xslMDtwKkX
DKx5X6EMiX4Qff7Oq4wKuAi6K1oMA/zBzn7vOmJH3/cHONWF/Gzq4ShMrm+O8SUQ
Oqi/jKpePw8FLVq6UVZC4FGQSqwGTHH2nxHWeDmxGx+oifYJ3rgpk36xv1TgM34Y
d9DOOponAGS/BUbQ6xZohR3KRl4FJqq8bWICiklNlgU=
`protect END_PROTECTED
