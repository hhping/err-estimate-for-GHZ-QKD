`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfYPdiJ5IcnCMI7fxr4MoUFGICCH3jO0voTH4rqKo3EMNwH8GUD2uC9J08IK0I3J
C1VLD66E4WLw4caBQge7DtmJGWMMmlichqVqlak0P8WHeqF3KBWH6UkCIgdIyxpK
2/5uljkfPw65mufS24fCoCHDOnjfozAgBwsw8qADghcwSTs0pwM++Ik6Y6QAG724
CPV9duv+/Dw1VoA7g01Ih0ggSyXQSNvSGoSYGKGkT17GpCtQJ03esKt696Z2QJh/
/TdcSAsnSRFQlmljfqg4h6/7LX7BnKfMG2E0sZSdj/WC2WgqL4ywOHJMxU6/+12g
k9yVWDMBI2UtyLmK+KT80aEtTM2JvmzOp5ZKdM2fc8mP5I6psRIfWJUZ/mDwGiXG
zBl2onA9EOuJTMkN+kiLbSAt8eQjDdwVvZ9y3odepYsd82OibiwrQYNUhJcuhH9I
AnfsCv8Mn/17v38qX0J/DssC3aoRkvl8pod+J6HPgnRSxG82LB4tiyC+2cRdM7YW
DeKL8xorAngcfvMz1tiYV2PoUBomWeK8+b+6Yb7m9HbLFf4oP5ZNCpH6Nccnf5Yz
zIKwY6JGmzHGsIvy6dRLAxdS1BsZOE/rZWfQtG1VoLoHy43BRDokfxBJiOSVLm5n
47zjHpd5eqjlnOjl3r8hzzUaHBCylpDVyUTlmozIFsop2dLQxNtiFT/egz8w35OX
+8UHwaaO99mj1X/pbHq94LnwhLn6Zf3T6YxnYhtpXhfqOPIzK6V3ImL+KhpMJN98
BVwfb/fvOOv7T3gk+hgj0AYzDPNfLQVJr3VgyT/FpQ7pzCWAPxc/3+wZNFViNYlh
7yZQwz+m+dSY1NAzeJx/EQ==
`protect END_PROTECTED
