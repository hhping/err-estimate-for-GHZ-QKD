`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDPtD+98JbONhNYLutkWBzRfkPzM+RQVjS7k4j0mUS4DPbf355M2GRWJMZ8qfGK3
5skx6Ooz6nXjSi/cRJNTfHGw94fhZz0zw+gukc9jK0pgoTECG+YdDtIdl1giqm/o
bZW+ePu1MV5ceDG7qV/PrkHQ8Gi8Kol5GAXjZ4zdTLBdJQ7ahK86YmVpxNJfNQRa
tKf2tIV0bVVqyZHtzxdOXbC1tBkGkslQjkUry7sQnvjK3mwzeDqTfQpKYZr8OqBL
qq4xeIQvwBwQed48JWyOfrW2WM9A4vSs64CvQrFVMjlr4NnBClaP5CvL3SJXSpXq
3ZLv+ALgzoLBurl8urWBYQdhNck2fIez/owNUULY6hwtxKFIHGqsP43vPT9/dR9X
/kGLziez4og9AzaRx6TuhStJTrY25KlizhpRmeUUTgZfmX6lYNk/NNUwnjSmdIHh
DGSI+VZopUTd37+oqq+02eBxXKf3n7X5Vl+dP+pFKW+GqFcnqCV/SHdcvG4zwltv
T1SMdr0CRnmKkCGRu6gUeIk2VoWQh8qvmwf+5gTDE30uzj/SLjXdlsY53C/90yVh
6Lp4Z3D5rbHUFJnf+khObgbolBkiYAbIpuHLq4LYGLGxSsmViC0FbCW5svhSmHIw
JCiSN11UvVsK3p7pwv7FWMLt/BMr8JOIOZICZIOtTooqHBNHQRloHP4LRyJIROVL
59SJ+kl6r5O7cB0hEqvuqHaNdeh4HEG7c/0aJQMFR92kWBtaI+9yvqa+N4Z5X9tY
CHyo2a5QPZGFiBEsrzSaFN15gWKqVB+APf5a2cOLdNS45W4gJFFsvQztnaPd4tQI
sr7LKvpDsngrgZ7eQj2GIdxYVrQFG2ZDxBzXCXylyF+D5ieABdsy3IEyr1XghDJD
NnZkW6h50UktO8QAd6uwYfduo6fdALbUvt7ZY0xavklA/vCxWQkHiMtuUcfydt39
SKSSh1nUon2PLi2IXWIE76I0V3Q2B3nWVSlm0sW8MjhhrhrftidrrFPhBTSapoiU
8BZh3igtP7ssPLW5Pm32pLYrdsei9onuSCC8Hao0dAyrch30NY6xH5bswoNJOLCk
w91kwUoNiqYYIhjGEoN1lHt8zHhsKHWFFFy0jEbif3rFny/AAQoQ3BXCRFS5dXn9
zS3e3mJonue0K/JES3fb9MQoCMG5/kJcpJobZUNAAFWo1Bio/3EpKVYQzF33Zb19
xSGipezTApzSzRK5X6IbiDu5HVgtUQDnPyj0AGmHaEEA+voitJaDmKqmGpog70TQ
SFtSxloFwGokS08TxAXr1fU4RvpHNKybe0RSGrNsKNqHOiBFpNkYUz11GjY/RpWv
atOGIksKP1AWzH65JfId8FHnBt1dNccx5NLcwN5A+iaVFsM0KbaG5ulctn+fMNVv
JAWWpBJGr+1BS987p4d0tEiChn1Na3mecpBrXXk3RgypdUJ5qsD5CpkuiigMCkti
5eFO2zq8DItRVsnbJP0BdZP6i7uOvhTQKPDMlCulpTA7jZxxWcBZD/iu+6aZpXe3
hAsVv+UUY1vpI+fOeYolDFKVVwj/oFMWAlXVI2XDWQrBVcdejakIlj4XCivkb4As
MEEOGCHo9Kb6X1pNIMsh1/mbCD4utxHNOhDHiGk7aOg1PBQ6lBUjYpDvF2Omo9+R
KKl5Q6RU5+grQseJ2YH/b596/V6pP4f5t3ilLTp/xjO1yhxiFs/BEtvNPKFFEB83
Ni2u/a5nu0b5k5BwXeyF0oQW1PSS6Ju1H4R5seidbhP3OZqibrfXlZaM5jeW7z/J
FiSKj4VVYgZavXCTUGLE/013ZuSOQoVCGmjm65R2g21ciLvuqmQGwk4ywclwEble
/mcHV30kbHKdjl9oh5PblCj/Cny1Kwnm/d2IGCm8K0HDw1z14bQqQW9Nv0KUydfg
Mj5saCczkY9AAiUry4U+B9aS12KJ63ZQLZ51sMML9b+6bPRAM9yXGSO9mXL0VL7/
yNV+6+LHOXVuZJJwTkM8ISrktJULU/Y8p1m4er1gZuC8m08vknLYfpkQ9mRhFbNH
FqomILjx7W5EeE9jXsuT8X6SEo+2QGQTWh/kItYdU9Fw66z4gA2WAWfeNIJ7iM2H
FgGv7hyoM9j2bWYhSsIKxYaP+FGhSxKdz85lme2qC3aib5/VLkPoHZtUJznFYX0v
ITV5fOso3dx/8Em0hm28GDPJwN7mojfmsVVH6H6lHeKYrPt4ZLJbRuebJnGr+MTw
L1S7GFTYGOBkqUfjvplja29Uw98NSS5kn97Ct4wGB4jqX2ZT0OQQPFDqUZHn6UnK
xedkMwjoeCDwBDClZ7dQYHxBSLP5xRxwKTjo3ockaNw4Z70kfOgRpzNTvdZtQ8ve
49ZKWskkWoN4ci9FGgfxx3vBX9riNyuwlAiZtv3poWhjwVq6v/Kimp6kuaPRqpcm
LVZ5TSfS1H2EyduOA8BpJDxh44fvUY3OnJ0XIBq2ZllvKDFTit/xcXCxyQ+lPWon
i6RCsHQLFBtL2+PB9m+JBVEOe68HWYo2krj205vqcbSPonQUUMu10kNTsjj1I2wu
`protect END_PROTECTED
