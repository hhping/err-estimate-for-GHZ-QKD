`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpQzGzu7eVQcL2yVjOoc9vyKTGOJADa8/uq58JbDRRFfcTIWYlsbaHmQgIsEGKWk
AkfkKNmfJbsyM15zwrCr91rsrxp6sWRxBFQtev0kBRw2BXaXNRNzb5+klTifg44E
0d3Xeil0bqmlg65sBIS+TsLuTxD8I5S6RPFB9E8mA7QTzqHU1zPSUnfqEmuljzUP
42WnrmjLrJpuV1YbY2gXcwZsYS54kVSVBxWgJCrbOcJKmhts8BDCIvPw4tWreQfc
t396IUj1yNkUVOdjKZRT57IFD15wQU9B2Zt1p0NZbxtKYqvZsiIPsPIHjWXySRoO
dUT0Iya7eXv/rvr6f+yVep0w1L7SSy6CRxWkZnh0Ta9JUAm9Iu3rwITJwcp6wFwF
`protect END_PROTECTED
