`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHNy+C4mKh88B/XGkZhMFeEafKDjlcKpS+TEJVNqgwNQxpJAQwTI7h6Jt+C2X+Aq
B+GckDRH5rwcAs4a8LRi4aTLBcho2FAHmK3OwxVPVqAu12TLobafXvXaO3HlEWG/
KNkt0WaS5UbzhVhwpFodEkbO6a7anNsuntPNEfDIwWS7WEyehwYeYf9sYD3wEhsA
iqrUqraNIEL9Es2Wrwt7mpFijMaoseEgd3DQvGpBtbC+PW09C3OwZO3TME6AYZ9D
qdEdh6dQYAJyM4Mvwn4/+kAB+8VRk8T2z4tADOOYp+dy91d7ObpcrVxW8wI458xz
ao2SzmKJ+sKykVi6Wu0w3zIOElU80CVt+267/WfHlIfoNtIKA28QwBtNE8Y69X2a
4W25Ad10o0OvezE47bQucWcer8XtKhW1DEzTHPjzhxha7oBkaTqVd/AstoeJgY2i
ppFBTFEPSrlU4c9F5ErGmrKqxz8esusxc3iS4jwBpMWVdpmBVYYbQlWip2ki8gp6
Ep7g1x/bAYt6MA/OR+9sdg8DhaLhGF62vkT2Dz1TXjgDJAVKCnppckRT7E6YIMtE
LUFLXyXO2/EDeIQYu8w/w8uUAYTmDHrIsw9d/EiQGzEChnZAH5NebMPM8OIldBFB
FOOUh3Ngp5gII18Pqiq1zLPHa/VUmPdysGD8EhOevRLnPh2ZPBbIVuGLRinMWMht
cgK+nGtnP65gXApZymYNFqlRwjXm38dKvrTPjRx/RaEoZAMWPWtvSDR52efdLT8E
Q3BpCH09krpXKMVTXhISRq2affZVvdz0VHLy2gFo+SA+8f4ORNOi/O6rq7/+b03G
I1h5tCEWtUP794+Q9o9gokd0KUL3x6bacc52AlCSZ8K83jS86YMG2AtPitCIpbBe
Mbz1lIkNP5blVG4boLNTJIfMkv243uk671+zXrJj2Yz+pK5N0TVBvs0DA8v6LHuR
Y5FW94bRlUR89/qshymRPiOvP/vnsQKrneHlwg6Nitk=
`protect END_PROTECTED
