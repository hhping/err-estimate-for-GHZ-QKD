`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HsARV93b7NZVY6XT9BeSFFbC1r/TQKHEschGlFCmYVmt4whl5If8IBIjThR96JrZ
9XPy+7v8heVJ/FcD7tCl++okoVdpx1FACyClTxejDscjq+36yW9e0Hk8lBwWu9R4
Czs6JGx7KCHO08QNs7slWO/SUGujwoB65/kEbYMdSFK/0OYHEJyyTQZhHBG9i+rw
59mwpwkj4hZ6+bJ2b0wOf5OhdvozhGCkc5flH+LN7iYYaUxIidsSUXD+byblo5w4
4CReXFZGjQNExa9X6UWgucJqQBYTl9iTHO1Zl4RySalwvgKkOUBRV4AEXxiQXs1I
oGgcQdn1Pv1Okw2yndBnqdmB40/Zm2RA/76VyRNW6tWTzfmnnLE3iWXfz6ekMWG0
SLdYBnyL760bcXFBwZJYCMjrG9xpBGaZQe8egXwcVr4A/IKFyrctVWVgqt6Dmi2y
K+G286zy9RKYqWvPnDIM4GcmYxCbwYIxDsqxyq4YywDoqJU2t86i6Qus3SYNsF/j
zE9es4bn4I5lhZB//oYUc0U/yM+NxvNBkkc7nnH60R0tHDq3jOgeKiNqIg4lA8ju
bsz/oZETPxu+kqo29TGWiMArfT/EZ0SeG7kOlu5sGezlk2A+kA6F/BDhlha1nwbT
X9DEjfgSeqCtrAV/dFIEpnP0GezOJy2bX/LiKpCMhkTabCUBS+WRQx4KZfAdfxt1
jiI6OzD7XS2TkkJW1VKodlQxLX1Oul7AYFW1u4VaJT4=
`protect END_PROTECTED
