`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWvaCK929mHtwhMJjsGXkHQK1FObD6ELJc2iSNhPyftLvl99FLyFMoNWGVObijsr
ioyxnBQN0zhjz2AHE2Ow6EW0yIVd1oNtQn7RuUwDNwp7KTStDfpKKgQahagK6cfx
niRxhZBaRkRglHBi1Q0+zYmuSlEJ0VBY/AE6qjb7t+HIGz8ypBYolFWlKroQwouB
fsMoa+NPmOZ8Bh9kNTogFqOgebXrwmfeqm7aaF0Qdda44n/KeARcFIb+5diFx6HZ
fheFkEETUEZxxi9aoOGX8x7CfqaTo5TVKru2+A/239YzZohvnZxqfiu3fUstJerj
b4LZcNvTqj9vJSs9pWV7txflmDyweVJF3uXo8hXrKuWWGm8NKKJu3O4w5NgDRpwy
+P2v9EjK+2K+/CecvrCABw3Jdr8/tZuIkb7RIvtCM+3EHHiNtu3Kxt3WV+F/cf38
IznKu6sVc6kmiHkKNSZZt15pnvMceCUpa/8HoSy6CX1f9DAx2QUt4qj08vyQdJxI
EhUOoizt3DkpJZQKDr5UHfwOY1l7bphCPBedTsgpNibicvCfMNNp4EYiAalZ8DGY
fT2nIdMcMjfnwWrlDoPjtT6n96uIkO0HOWY9/zJyAdPHb6ha36/wFsAxi7Rb3QIx
l41MT88NECGyUdFvpcnQ3ysw1RUx+0caWbC2iQx12UCJV10m4+w5jH1+sNQHHrqK
d39WFtb+0FBv4Cb0jpDQZ0zWROiLvcMWkzrM3IsU2SyQYXvpfuF5Esz+KDB2KZP+
NRweEEEmJqGuwUvWtK8oTMdzre/g8gjD+xsJXFVyTDtvk/AWb98MEb37zYF6HRcS
/LaiyJ0qIZ0ZkL0uVzFIpHjQx2UrunIO/UwNmut1DE7UKYgNPC9D5HRpUaznRQWv
fbRakuWzHUxkRwNKxlrhOJrZgA97aGe6ZX29UNp6F/ZP4AMFZP+mE4KioqkZ9kCM
vo64UUq6FJwlvRLlnRzhRdw0tjWb9ZXo7AqVpB4e4Zk+x2dOPDdAs1gsHQqcEyTp
Z0Ik+nNOpGIH/UDSR4nSaLItXlCb5ofDQMu4Ps4/6HsdmDpTqhRWEaViSGmt6pES
O+Xh8TxVVz/VJUO7R+egl9Z8hbKwfaTOTPz4tOcjOjGNVXbZvl/1ylqT5esPlEot
2mqlnTiNfJTl/5HytKfV6baERRi2pgTj1D9Ei9qkneFxarbHHhhFlTyJDvR/zLRI
d5l/yIXZ2U+2mfvqkvd+YbSxtZEuO6K0dnrVJEB5eQxCrhgtY68s4ZvKmk2owO4p
4b4oGNQzFGxsr+/IA4s3U/3jOMYara11K8VbkLtUg/ztCdQo6JDI992XEispQJS0
vw3MlTrngaa24wDHuTR0/nqwEQxvG5K49Obnep9rsx0yl1P9owp4XrzLwpp9Jrd0
1PLVm6KtYBaqO65CGTosFG8AdemEJJTVFp2PiAsc4tBwnLULQ2SdtOnJSSWX3nxq
oySbeIhMnxuJnyjGm5it5YRDRTbYHDL2qz/qwQN6hlt5PAbW9T0lWP/3Qt81isDx
JUTcX40ESXDaDvY0GlcmRcYqkWtcC6kdXdXVzggTAuHEtxJeR7zlVlJrQeFd7Xek
zGK/9OAkBdTmQ7vkQHEgzAelVt12NBGJncvG9c/5wATNxBM3MUouWdWqifGBGDVa
hYBisKrLkh1k3/ak59CfmXdb+cTLS7woTrnMY5zALZ0iE/LCw7jz6NHNXwCsGGIq
DD3lPafXTEKIbtFSzL8KaKt++Y1ud3EBuKrhp+KCApDj9IRch3xYOCEntDXZzdn7
Wn2AHMNXOBIiANswukHWWmjzh3K5/PZDNtsjQca2HGq4Cv8eU1HxpLuwS3iUG12Y
Dh1bfE1BkuW9PysUBEwQQr0dg8b+im6FauzwS/L8vmtavylm4Ct1b0RltaXHXkjp
RY7VZ9B8AVYG80+DxrRub4aYzlrzpMGFQp91F4PxITIWncRiejZHeLoRIDhFKjOo
xqAradtL6hjsemA8ZoqejsUi/7u+DMqcvaksk0Rot52FoIkuu3N7SbZubSi2tmH6
nZvVF00NFCMa0xBJtUkxfWhersNF9MycPOOaHkBwyLS3hGs8SodLFKJlaxmw5bpu
Hh14gL/hlvnshRfrFjpJLDzYGTHx006BsJMZhtq7ri7s4/RaJODSCE2a3HPhKTXv
MXkVCTDmpqDXAFV6qgnLFd/HaIPJf8tEtGxF/rQBGc7bC9x3IbXGPl/NiNeAoYSi
/cns/kFq1Wg0jZEqlFpjdMwABVV8WaXCUCp+qsTiyKclmOYUcg6EfggQ14wMymlr
uwKM6xbEDYzbS64/DSbRiwU5qRA40USa3jOXWzBIqCMxe/K40iCJ8gLOq3YsviWp
pNPbZhIqWfvF9fL38BRVBJzwM2sEOarqhZVLOO8HNgC1678YSz8iYdn/RJCoEfTq
3kVWwEQpn9DsFDE3urynwNJ0vTc5/XtoaOIluornvH4=
`protect END_PROTECTED
