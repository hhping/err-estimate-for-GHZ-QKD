`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDUsR759mz9HeRftal+YY1NV5cCxZ7DxfcIh5bOSkbwoX0zb+s/Lte3sfxb5HaAy
7/EI51UXeI/tH3mnnZwHvHppiSiky+PulzHPdLPafhyLYd2vXQCronc4Ns4UdnO8
r793G0NUsGJNgm0+/GFI+V5F8fWvUrLUtFUNIWg+JwfKU46c2MZTOS4ozpHCXWw5
E/gpuSSYtg32bryRAwgZ24A67RJ+kaHG5ADW8R+CP02CiZDFmLYOioUlP0WGPRy6
ixuZDy1aIDDMJ8chOegiw9txQOx0PNFiBJhdyTdFl3Ri1sV7Dbp0fIRiIO3+wVhW
CyIr/tEjTpSrzkY3CU7EJ8b/cyRfmZJiNSgvvrwoE/UTR+el5lSQk2OGFa8QjioS
GWnjWrnKSfO7oIy57rzyyk9y5LZ4vr129oCbWbjTOQSIzXS0ieIkGA0TL1tR4XI5
Zixp0vbgXhUYYHKRAqx+cfQ2J4zyuRA4uHbjc1NIJChHuC5pzMy6BNBUCqqwOwV8
6DyZoutuf19hBUVTRaHu19hxK+gqLKxJWnBVVOV0cU5A0dW4QFgUonE5J206ZSwx
jiPDTftSaqjvPQhvd34BXH5/R6dVrnN5fJHdz6xk0TGALIwISjKAczt5XwyRNVjt
ti1aSlhV7xItxHla2OQbyrSS022n6N8VBiuXZsjaL+GsWg3Zv5f5/6XppgDa6H47
DlR4QdABCRRvS1gLYptpfg==
`protect END_PROTECTED
