`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMOmtRWaEGPUuSS4bP83JmPg6370DwEokdtwQ9FLJfhP8uqWBkN38KVvSoiTFcdM
MRSNeeqpGyiKl9ayVSwgu7pjjvzCtfCfMweRmt/fG5p07t5wch36Ia2TWhpq69Pk
p0mgoXvliCBFEF3SFEOBCOFPnu6+YZaYjzt2pa3db7ClwS9j6DWkaTXraBoUH5O1
jhwxE/rl2QOHFSTbpE9yUP0tiGGOw7JzPfrc6SWeF7sQjpzO+LNtCrZaMgosq8sB
4Zhl+n4uJoi1A4eyg3X4JztzpEUXJgxt423Cy9hI7ZRM2D+GVxwjyUQ63nW0uv9v
8n0gXxDshYwtlOSdSvEKWUJJsmuCVE9xuf8YWrSqgqLaHQLVx6BKBhIAG5MLPJGj
ZtgHdAhY/4y5M2O5NRFwn375XScObXxLrT4GueP/+KWiVolDM6Lf3rawhQzkMGu3
J8bFmdOSKs5+bCZrToIrafKaVZ4t38peZqsTHyJMNBFEwOIQjZpr//MJTaJL+oR2
PagSYUrDUkgKpknBm2KP4SZESesSy49smZBzCXovqoQ=
`protect END_PROTECTED
