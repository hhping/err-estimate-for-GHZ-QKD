`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdKZNrP/pKbyf7juxASzMvw/aLZTgexfS1inWZNg49rEJbfMBmztCpWE1vNP/JFJ
uD/qyGctf44/OlkyMioZdFzbiCEEvZU5xK5xKtwfppwl+K+Z15QYw8UlMifwdccE
+zy9LcCPowdlcTrLXu5dzcwmOq6DuVJzWQGx5dzY5tEvAqwFtFkvYi/Sxsv7jj0A
qfAGQEKtx706cpaK7aWiIaO3jE423swzdxeFfQ2IsoMLgrvd3NgiVeKsL/dsg02m
oXMUZBsrncJJdwmjtRIYTvH8/HPAz6kf882MVXdJV6QpoaZLrxgVKNo4qT1hkAm9
wF0Ep0fxM3Rbpam33ZsGdfMViaepbGsrenIgSWh2gKl0dlZKozTl3sAE8PcRywrT
Bis3K4EGeuD0HCDuLz2lhrAa7Rbueq3zejM7BHN5LcuiXfFZH56JKrROENV5LndH
qGSltfExY2Ax5LqE81uaq4B/NEAoDws8V8+f78SUSNQt5bah+1RhvEiii03XyNf9
OBWwjGNc6wdbK4VMuMK7GGen1Rl7B5D6hRCST8TcB3BjFgHsDkGZ5bmVjP1yLEim
jiPB5WHGR5D8O7n5+xRiZ8VhpPZm8ys2Ene18fusF2U=
`protect END_PROTECTED
