`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZdPQ+4ClpqwSA9OWMxbnWCF83EdwZMHe6KVQx9mzUj1tsN1FTBJx1Wbsj+Z32wq
ac4wwBLiXtTGQkrnejVlEbB9N5EmDSKAQUouVFLDre+QG5fRZ7QpvVX7fuqCHQ7q
o4PGU3bzfZIanl8bl9BqwQuI4nOeohNzzeS47n3SkiChHMlMuMaZB1n9GpHwnW0f
R9cpnu2R/6sMzv9Kxiojh7K2xJHG1ivRZRfrRw+OcExnYCNNIJGGVH7HDE7JeHjT
CKf/1C+OPQ16W7TO4c2F8if7lAJRpOMpF7DV//ipzKRZo6a6AlyH9WJgpMeNgxRH
1ATSP7XFtEvbYxENRSzZ3fwN23JO9Uc8Abdt454wxtffnMyaRFQAEo/6mrFc+Lra
xG826RWtzhfB/kmhiIGGaIRqKRtd726qMgHNmIwd2C9/C+cRmcHo31++aqE3MflM
gK3ZTv4Yge9r/7m32S8My/I4mbbHCqwVzRRF6v9fzo7UTyDumvNODshx2ursQdVe
FOP3zBOY6pO+3pPiDpJA7YvZP381Hh0WJjZJ13NH6eG6i0oJ3DCX0MLIPT3t1fjM
`protect END_PROTECTED
