`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6STjQukdWecE13Y4cGs3JhoBkfoMiKEfK3IiHpmw9ZmzGmLzMYooQRoMf0CzFomm
z1lzKJ4pjytM5ascdhHV+PChYDF5UY0xVYGAg6M1cNCNu+9JSLIiAjn99GGljIgr
guGcxjWEmbB3FD3giQJtIj1WeV3lKfYkTFTkw+UaUNltJVqwJ3yD/GpWdsUKTXn0
MqLddcmxMvbA74lOO3NREs4wu76sWdlQNS/ZegxIJsihxGOKbFJxYCPw+8BcSvxr
JrVPLqgN4k4epd5aZ1vRuwHiYD1zfFy6yi83n1tTpihq6yu4fmqhMCAQFTkoNAIm
9ouoESH19RkfWpJddHvp38bdeRQguQdIY1S/Co/wdlUf9q+QmeDvU74YSma+iBRV
vaTa5UXED47fStuuzudvXJ+AF+mD4RcwI97Mum3xAkfa3BYU4M7MgDdePRiwGwYh
3Qst7Drz7oBxgwnSxEHQNhmtpnkp48ATBaMkPIMlS7kcci/5UxBb3IDPv82ZdrHu
3DSTZa4gzbNoxxkRhMyee7ysbec8/2rA75l4Vn6+pquFD7RQdWv+vC0LAyb0HY8U
fM678WnP95sQ9SGRx/z6EEyeSRPiyXKLq2XvUbLZsXbRJwW9uq77a8yBIa8vzGzC
A0ovSbHWwPfopqvD3NuWC5zSdtUwyZF68XSeIDbkshawzFdc8o2AQZV4psm3w8VD
t/PhZOlXQVYK8Q74A1ahrN/VDtQbiH/QltHbaJA0MHh4Tl8nsNYE3nkwta+/qxy8
e6LTpBINQ+YizuJoTTn+JOdBX3ot3pzE/qsfNp7vM//7uwT660ahTSBEzPp+/tdK
bE5ZaCXJSSk0lcRoGiHcG9sT93s8kiBPwjdCBKr6oW+mvlqMRWS/acHcj8enS9c5
`protect END_PROTECTED
