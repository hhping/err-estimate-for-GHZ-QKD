`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIciMC4ZWE6T3EV6Qe9ix+1V5ZS8j451NF8EygLNJtqZoUTDj8q0uw6WBsiyhELe
L7q1rwIObpIGS4ast/Ily5X843b9FdGZbiAxHl8eHq6G+XVca77w+OryOAc2dzpM
9X4XjghhrXavct1eGG3TtFOqAGu3c2bIyZ3PkFCDj/R5CyGwjaAyTyRiMDbVtt/U
TXIocTIwUk990ohne42HKZidR4uIBpTfjvROgvC19KmiJC66MaF6hZ3ztVVI2eDU
4cNwZYwrd7dGyI1G+JVD2VjARatqJ6fI+zC7ecnjtd2lrv1zCqy7IX18qphbKH2i
HiAlhZv0zA1BFfwG3y3Vw8h2K7AkfzIf5KdqIPSBqCq06ekPSWKi0UdivCGkMl2N
FtisI+aJyN9vuFpE9iLZNyGX3x0+DVChHPcWW7TqnTudTpC2jt5F/s8QhtvMDEjY
931K9Xeu2hEWVWY+0CD0JCmmUZHK7nCh9G8qZ8L4h7K3fmgP+bRZ/coCmqjwtYPi
D3dEE2Wgc1oFZDDFWzCPYsd/3kGT5eF4e7ApCO6BqyeTGfATpSYYbo885EW8skif
TCqs1BsQKXRz7bsnfQmAwBpoVOD/R2t9hSaWBU68DNRxXiUjzgyc1QLTz5nKq1Q/
u0Dr+NYHxQjDxXmdIxMRd/l+edBAWxoIBtjSv4OAzEe1hqN458w3hpPmbVvpamKH
7fldY2pr1n4rXQl8O3S7bTY8PCWFT3kcd4bMGPYeVoNTvp/NeRXVsaW3EQFdMywt
nPfkYZn4vHUS4aU9zTJLC2Db5SfXQz885lPPLiS5QK5gT9xXiHE6ho/tEN9GPuxa
IQGGObiX8SrhiSPH4suq26mGBpa5RKqKUnWnoIGynovVAKOPyc0Af25JabDhEsE4
Qc/kJpAd99Loi7okEyO7c4d1+1nStvUPhaHRX1IXhlMcIx0+LWSa8MAwnkR2Yjc+
BK0JE6u3I4eEEVK4doJlBA8LbY0yZCo5sziVe/gF0HtowvckgplV45QQ31O665Jk
ufjrd1RlRLYikqI1w9d1VigbcpWODHdP/ytin3CK01j2Z6R4tTV/dB91HSh5NBJg
0dYJHSURcJ6mDmJOeGptz18SHZZ86ids08DM+wtTCuQJ70nXP1T7xEaDx3sFGY4Q
5lScC4+WWKyPl9HmFVgF60LnMbkZmdESMC2HNZqnNb013X4ebQFfIJGRH/ZBST1v
KYaZYOYQcxu3F2gWzzpL9h8UtSY5VSlz18JNKSGWt/j5SjcTSkJQBs1smi+Sl9rU
2KuJiIaVeJKRC/1sFviQNRunyduvBZclxzLw9dab8dwBRvAmfIj5Lhq/PvCaxgYZ
8BDZFdT1manbtmvZ1qqQNm/XMllJe33X2+5XnLqhZ2l3Qy0VMzaiJ3W9p71Eie4u
QKCIBEMNXINGe+8L+w/9mMKDa0Crwo9LEgjscgihcYVXdzIxVCV6f4nAyjY9Yfku
Xeg85UvfVYTgbaw/90zQMWniJgA5Lt1KfGcUd3VXZnLDjawE2WUTW/L4PG1iDGzi
MJmr5ts8YO1m3UDBf3Y8s1HptS71doWAVqPe2I6SdT/Mhz0nEG/hTjhfGui3k6gg
akG4Mt6wv+NDISVMoKeMT2XHFFCig2UxX/Rj3Ev1tKp6oIv4Vbx71a0OfGO86q4Z
kyqW4+8AKfFdAkkEx1K5HcJ6ZCFIQOKf0CG25DZPvhJHC5Btdl6jDvoW9xGcHudX
utwavm7h9swu97iQm+LcAbKHnRQWwtvBjgs3rLrKKcd/xxwO1nUAlYXdryu+caYu
My3LYgPBbPbQJLMAzcIEX5bTTYKCbCH0RKW93RPLNXNMYCarajavr4bPvoUnPnkn
eWhuEMiDEAva6JZY1io8Yr8yoGg1DS2UbJoZAQVPWIorKKlH3dhTxPLZnXnNeQfy
jxfZzrpZH7H5x5MvPWWG/q9XfLtALzxG9djlANeCVtNXskP7tXQ5FKxA0xpH0iDK
gcq0Oc1HGpktDJ126IgbJ3hXhYComO5h94sv1zp8D7l/Ufr4kgn93npzSRyYbMSq
75n1H77PrgmneZpCJ8x9Fwxfm+peZBt+w5F5830EmnZz+AvmBnWs8BCpk2iE+1Bz
SQIIrow2iAdlkrSpJPz/m3Ae5hPp4/RSOHqnZ/0N5XZ64daprlri5sExWajieKf2
tpRRmtMp41ZZ3FLU1P9PryEb3mWKAYv3+nLegfx1N2Q9L55Q3Zd0jdtra6P01Mw1
H7z9WeUJWZVk9+GmpTmekhYnP9454J8IWtQPutheEUx7uobD1u9I50ps2kC21L6i
03B4iZSHR9EdQffb4tHirkehgtww7hRRU3xfwd92OlUEoh1NaoWOWGy7/2VIwWYc
cUbC+S4uZH3IGUL0diUtwZFtxnZHU4Pt+Hl+Ljh0kATmcKtrSxPKZXcD11gLqmjv
kmOgIxH+oNCP7OQ68t4SQ3CUUQ5DPjib1LqtCKBNuFMlNF8Sy0nDxIdG1IUj2FEY
kTi2ZqnL+VASnP4sqiLtBxW6/QHGzP5ZLbPRY3pTrMTx/BAQYCQAh9+ipAuPSqAS
b7t/Rv2XdwnJgoeKlwqlaZr0LMBNcf5ihpWuwyIQv3KOt2xU1i/17okFe2jdgCEg
7tBL7yZVL62bNOq6rYrU+Q2uPF8LC/Tizy3l1BSCDrGAVECVPfOGZIilsZVTBSDm
C4nIbyV44fbOp56hSWXb7J0EelAq4qV1pTKc8jmKRKmrUnFstsTX3Z1OD74L70s5
Vd+WEhp9e+0oU4MLqLYYUUcHezp4IEtnqBkjXb3lLBADNxoQhtaa9VXyRSZAwDJr
40pYje/o8K/YvHzrbte1fBUKXMQo06AG8kHCrmCVKP0cLrYuQSiiLgCiWFralFZc
iToJf71YAb/NOX+t+DgrojAAJjZgnMefsUaKXv46icvluCJZTbOkbkKj7t7C5Qc9
bLn7pZqnD+sIriUzJx1Rffs/UrQndSevwMDVrD/LzoeNUecHqmEJQ0kOQm8HzRz3
NwujXwHbuO8CZ/tMnhKbQFVj7v/eSz7Sb4qfZt4s4h2CUwMKP6Wfu3BYEygWneNk
HVueEmeMODq/cL9WgeElsws49ptA5KpHsfLw5f0PcT0D9b/dfWs1Se+AL8/2b7Da
QHIAIkj9gs+miBaFNfR88fkQN28Km2/sMY8D9ijKECF2xS3RXPwRhuChVZY2xnp/
5ZpK9eVWBuQv890nK1YTNS/iEp/BbWm4H+Ljow81tb2EGn/ZO3CXFXkySqJtxcTn
pdKRwsYLSZJT62vozYxFT7/45sZmJR3i9H5s6Hu7MjzEIfTskEfVdZAxTJ31BovB
YqWVNiLNZ8Ty6jLGxTJCyhVYG/Y7cm5LtERJ8PTQZ73o/UvYftlK0znF3Pa/ltPV
aAynDewXji+SXlE9KW1Mcw==
`protect END_PROTECTED
