`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/dK7oL/dVjeXhMH4y/NeXXQPZi5D7CF5vuCFxPa3OLH3sSaHu8wuKzI9vhUVEEsa
h9DwYSA7dkgW7ORUW4qGF6lq84m3WU1uw0oDRP8soAuDGSZIcp1R+4UGF1Z7ABcK
7hTtx0aXfAlVPfnyTfVaEK6sl4PHGqOt4wTvLg7EQUI3Hayh8/TeP8w8mO3MgZPC
fsfcYh9cdLKLNjAM8PgXpiStCBx0ZGRHHRNdArCOGYwQ4+Sb/KWxYqcdM4Ju6GvT
kSsBBDQMD2jVgvBkBYQo0NG7p6TeK0vFu/QiNBekDD8QlwGTLUkvpHAN7sQbckB5
soO4RsQHD2FSEnCwRmLAFf+WYEURzHVYASNShGGd26lSQ7/uLM/KTO504f49VMd6
FvLXY4TuDmoeJ4VQ8gZopn6YAwxabm3rFrvoZM4bTbDh6IMcugb5H0D70TsKfXcG
lbr94hu4Ni2H1H3KTF0bKYQbizFF3g68WN3BrOgci27+GElWCwXO6KwxxV16aEBq
PaSkiGKpgz+4Azp5x3+NxvksGAvquHq7iaq+euiKe2W1c7kBxFn+N427LV0qCLce
Thc8NPnZ+sk5nEo+24jOkVMXsYoixU9N6TejRt6wJLP3PpMObNdnyDPBQbgglgeV
`protect END_PROTECTED
