`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kP8utU3FckMyG1RDum+KXoDROIJz8gSxn7t5Jizkx3HDct42JK06eTNF9C17j3wz
FMu19YcTuL7EjAaWstTthzBh1kGFLPhAnKLHI2FjYjrkDtoT8gt57FeW1H+/9LNx
+egjQV9Uo8tyKvHyCzsAtDpR+ck73MRpg5zYWChlnUqpWl2Rq/jnQFiVRP+PnDqt
3IKX1Bn0qD6gUEtN90KzgWAk1TSJNZPZFX8yuJT5gmFNxlRgSz6BWzKpsyEWqMV9
Mf1XG+Lh5lwwWPbB+qO6pHoNon4FxaetGgrBTN8WSxcSlNAFYzhXwFrqIxGptKLA
Ga1LfPsb7XE3D0iAxbo3Vr5X0huwCd6EsjOlXb8F+xZr3JpWPpIkhXrf8F03fK68
qdg0YdkUkCTERoLQSOsMXn1Pzlvac2cE3ANxbBSFtImr4B0QG2B9kvc8L8ooKAzR
ibzwK0C/mAvGrPx5P/caUJIDaBMlUw4rT5siJzAhsJc/2CrKhJzHPdLBJ6UPUxBA
myb1ZnfNDaND9Z7+xftsS2pWdDdt7HDvMpKnSYhDPYNa1GFD8i1RC3D+HpLrzUQ4
bKedt0ekuGv8SQIgVyxNLkQkDlIMPxX5VS3LXuuByNuNOb4gIuY7zxpSPnbaEWET
cmFu0p/9w21DU7yFdVCWKnDSEfpjO6c7Ix/EqOXp2jOOHOj3kKO+aE+bUHc5jQRN
s6gi/DPltt1NVkdPGCQZjJyur7Upz+2sXJewWv5e7Qgwajp5vM6++xwUxV6znyhQ
8JGj9d82qEXioAKMj6xUDKBZJwVGom+ubxGCX9XHKfjzV2jIjJn9rN8c3LsXckYc
Z2PlSfEEOz4LwNcPb7Rp/x11bNWSh/O7AXL2fUiAC0Nf6jizDERg4Q4lGZxWhvng
BNGHo8p5k/g2zVuvyO8YofmgR8iQwUfuKE6AjUevAusxcrSX7jO6IgmzaGwzgxeQ
92L2eq4lni+yEtY9HGmdwVbnVwzO5TMmXbto6TQ2MGVDVl2KlodVUWItlxZEB+ok
vf6LQlj5S+4JWy2jLS7ConeVViehnuBVwkCm+wiXwYKhU9frvId7nVciPCCDqHy6
7YUvu6TRzzoP2fjyQ6svM7d9vp7UFAHuJJqFjlVV+TJ7wDdtch0198vs4VmD6OM2
qsdb8Fc3cS4LYahGnJ6rHmlYXvjay8658RC8CBgMFe53Sbu6qfE036PuGI5+yAjZ
ga+yE0L0Th3gnKYy+5emi9MTYwRjddDnzyRVmFlCyQYJAx895Tvkdv/q5IK3ZrEK
ah48rnLlWL1/5MT8Zt+sE3IE6m4rwsPLEPKs5o2lhe8KEUFZsS/Ab2upXE+KNJhS
j0b8VqByAcob55XBHol673Tk013OHAsnRokR+JwFR+dAhbXhCLDi6c2LEJnN3X0X
Z7/mnCO+DQ5BKR9/6UfJhxUlAXVzwjmyJnhkkkaLiCnNJNYbmeY5r/itTcoTU7v1
wmgxxwtQUv69VWdCdDkE0iIkYjPFr5O7Dr4N9Wo8HmBTOknfCn418I+rH28XhmMo
5zO90nEkgoDWWxuWXd3KNTOc2nFo+O4LTS6fILZIIacshyp3cTOdNOsBLrIjhVC0
VDm50eX3Qvyyl+tso71cKAxOK9Zzzux0SMXkr7H6vb2LNmJ/Zkd9poPV+rrUhiw8
WtYtutdBU2METj2dkqYF9N4rOt+n8XuUYKTIU+QCPElwB3NycxMyPFt2oAy4LQYk
cWGHZ//Dcpw/JpvO4rwvK/5tDD0lKACgE4nxnX+kZDUD+Uss82xflamD6D/9rKXV
3PH6dhqdVoCuM5DjjCh/KQA9tOofbysyBqzA4a8teYZYyXR5diFPNKFk3HsWOx7H
NcJh9gshZWFUH0kmbAZdpw32mPrrJ41QhfOCa0dh6tZNYhrywLJo/ASGAZz4Skzu
5yVfT7xgXYetScffRGl4RTuQ0SI6DQLMrmrdJC3B330=
`protect END_PROTECTED
