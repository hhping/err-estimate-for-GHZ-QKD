`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZCvVgszvsgXdwkzsJti/OsPFrf4FYU+kcsTbChIa+rPIcr1NZafIN488AIji59W
jUygG/QfqezYMeSxYYhjpd7WhiZ2md7BZKM3OUktys9qnKcIZ9ePw0KdlYWgRwYN
ShNXzhezQ0HBN34TZp0RCp9YPHDz7PlDxGGbqnSEVRhVeH5xatKohPxU1fTvVkM1
VYHp7bEry6/Hbo/AJ0+34aWqxQEb0FrD3s2ywWamOVWV2/6IBuLaom5VBZleQXT3
kWCit+frKYnOoKdE7UNXupO41ZfUyRbgoyTiHP4nT2qiirkZEPJIjVyTfSQ7gP5X
3XWHXI3lBGjEftslkQ0k+ItujoRGn3pbfB5uo5W8HKQf7kdnRYoRTTZNNE9UP6CR
2apyaMMYwtAkZGLb/kU8iJq9ZZH/qVYEVw6y4RsqSv2vCMQ9hJKXjk5A82KAm3JZ
dD83q2eJbohfc72ppWlE6pJilTSzFWwmQ9trm9KlSGlzHTvoto1IyW8aOCGQTSnP
EOVAhFu/ZLESL57P7I5fhVh3NF39Eu1aeyYnZiY332JOnOWrFMgfnKEGGlv1kyth
VkbK7ODczj+wrCqVXufMeCxCSKq6dfM+71rP9OSrk6w1fn/fl56pgSD4uOtFfLmR
NyDHlyGiv1430wPJg60a7g30wOhDsLcjhv+MT8nUhAoxuRQAMR9RB/TI81TimT/Y
TlKKAK1r++V29nZY2eKm4weV3xOxg210U79BH5w1P4SbNNcTAzVGunqSoOjmjJ8A
67scW3N1KWnbcQUy6OScFMRtZJOiOZkw4uGkJ904wsYUfLglBpgeU4NuPJbOfQSn
QQZQrZPVrzufkpgOkqbazz+Pf6AqXAL6l+s/LmxgDU7+nZFyNVGYbGfmc88mxfB6
PY2Cb23nzLPnoGE9jzZS25mk4c4CWWLLCz4Z/IJmsR4=
`protect END_PROTECTED
