`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99/Rw1pKv14gxTZQfRwfI1ME/7Cc8c2CwkKvxbVBqLKfrSGF1qhlaKJ/lrAc/Yv3
A2Mkwoqr8GjFboWQx9T9hj4stXigqisWHsXSHnJLDtczn+nFp6tUaG917vUpSQlu
o/D/9bh3nHIfni2P0Xj2ZqR3e8pHUVN1zzk0VYscMrlQwNDwIU7X9hvmL8vrvKDF
XOpRziMGTX7rRmvvkc1PB6jw/YBTP/6GFLIz0Gd5O4DklmAtVhDo+YsYbkrfW5Lh
lqDINvEj0QVlvpnkXQh/FwRVEGRh1mX5xwIEY9jCnbrdXQXyvpDxJ2ycTP2JfCNc
xHQR1GG1TFFxni5GoJD64+T4UVYO6Roc560E2KjCSzkH11yRNQYpwpBJJv5DwdmG
PjZ9N+FB80rQ0GpXB6jUix8yQ8lvblvF3KJtZ+/JEI12yiw2C1grQSZKK6JO33+/
EcMbdzpT+tDT3HYOjX1AOVoXOlSsjVjGm06/6XP8/nHqn937mkxEXNh1vMs9nVBm
Q/OYqIQIJBNKvHlNzEdsUAcbViEQ7t7R4vXyyug2JL5qURGkc6ml3KhOa9Wgp/bP
Ee0FYKentZzWXEKUU1SBQhZFSqMCkteepwY1iy4jq9tl8v3g9L+Q1OKK+rBsBHIA
zksvm5Bdzcb9ggQNi/iYTEktUcr1U4q2lO90eWkMIXwwNuLK3twrvJix+rd0Wd5m
lsvUBjw7tquEuwk/REh9smcmaKdvLAMkrKc1UVWOLD6pcZ6zmUe1xXeveKwK8w0n
`protect END_PROTECTED
