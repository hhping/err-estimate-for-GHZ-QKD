`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsSuSzi8mN4qiGk2mX4IuRxk6dMA3k2SaPZ95wNZqchWPeG6UqR54tKEteuZRCi3
kIDnB35DyJIQYcHOB0utKjpG3Eo+zeBvpHZiqCkcpKxV2iKHOag7mGVV5mttHb82
tSk58Iyzh3JCw8A/4I5fzZVhg9d2b3txJLP5XcZizFZg9l7S6I/tXOcsMMfEURXK
6rgi8jbgZ+4AQiE04GriofE+0SMhCPq8C+sVoDx6p3E2cPOUVldVFgRr/jMH/fR5
+R+QEWoo1WfyeZ8aqJmBpCSgyHX94zSeDtEIZZ787oTZ8NpFtlksQkAhqm7IJQpy
gbjF8KqivHmP4WcRxQ8GKsHc9WyEPJ4rbTu7AonTAK+DtLpNnh+ZPrC2F330uy87
uJKf10pX9TOuuYQ3LrHHiN9GYlQYOzv4IeCyu1WMRKZ1O5VJ8dDzl2vrSUCVp5O/
7C0BzdrXK0zl0iqw7Rd06uyo29bKN50NnlqwM1i3UafYha4JLu0Wo4qGk4mWPJob
rLSnhdkhgiEFLQP/fYQDefX/eVt+997RQ/ti3HtDJsm+7ZmTLI6CJPNEe3/QU89m
Z8ICXKLDmMBWQ5iqjujisI7z1nwTiDihCyTsIZTe5hu29U5V9L1hRjKs6ueLfBT9
HjHIm1nQEaTj42SIlNm/swLpngBzRBFZT/+WyTbOk4xLhBji2rbM19Q57C1mIu3h
zp//R/A0jqgU24Eadw2Q99NOeri9bRE2xMmSyADDLji+aVe9jPrTIpBxBX9ZPJUP
v1kE6BFMqarJLwsx+wgK8d0slK4lLp1EWRf3BimGbKVL2wS7rZbuHkex8mj2dFtd
PuK8dpwk3+baJCMxDNRd+6AKFbEuuwqx0VTFkrMHIX3ewSMSEBA6OsrewbY/HLd5
tqO8Atuuq0QIp8COmWt3JtXNq4kK0OKAYCjmnWHsTwnqb5grq3ij1S+jyFKj807S
FUFWMRoK8CwdJ9FODOO1l0iUCTugyyXzi1ggCXOcsWHaCQ92f5cg/WWjyDsHUVnF
I4DjsiKkC3h5NsQvI1lrjBk0jWzNCS69B2SjAw+JuZDKhF0z9OwKcIlH6rMu2VOl
EFA1wmec2ypLwDRIG1pbZiKExiERQfWQZCTv34V8ZyQ8RkXiEfD3/mj7pkO0BuME
+/1Wlg++Fo7mUUmgwWF8v5y4UX/D6b+UHL1BxFl74wbnmf9v0Vt62JaDXo7HuKXC
45flKSVP7i5KNCdmQMYv7sk338PkYuiTRI/VUu/8UijZf4sPLlk6GTY7hSQ1VsoT
eKbeSBCMpnzMypjVUyTQGpVh5KJoeBKegh6sDzdX3C95+0JwtZt9YXmy7LLjyEl8
U3hB9oTW10PVC4wp6Zt6XpcUsKddhugbtj+o2A/jY32BxrWP9wxhhDw9LCBuWgq7
+A0xibHeVkTH81hv8NcHfcTLtzcVmH3YTdaa9huGUjR4bl8+agyr8vdyzQ8+A3V0
Vb4Db+AwKzOcwAPdggatrklcZ0r2TFDKwHYgiCIHTpmAQJi2V2v5fw8wxL2p6FUw
8vcnAT+1ftx6dmawPcxWQMQhDB/G0CEHfFZvvPOicA/aaHVkFMAq4EAm7Q5SRK2p
jXlcz8/ry6hrNLRDwPtYUbBWvaoVZT2eEGpQHOc0Y5g5uFsHe+r0o9mSuRrJavAp
xM+yEWN2RnrCNn+YB2qlheGXasNddC1L2MOLmRhqzi0Bc2ZntYy2W+6vCx+mNJo7
AKd8FO7yShuJqejYVikXKA==
`protect END_PROTECTED
