`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9mnONrQOTIIj+q8WVxTZKk85CZtA+cllM34uBld9aaq9GQIWaW20FDmGC5AdlpLt
8DG81o5JcTCvstKeZyj4vZLH3mIVKGH0ODyANb6REsvBSW4uBl4GYmECwkkzaEkT
eBy02lRE7p+gPAayrQOAJDseQxwVjJMg0k+9EpwlJkmPXeo7qpKA6xIrYkYKWxjK
45khV2RiKOKmUApMIfP9l/cesCAL9w0E1ktdveAdkOArlFKnCS27joip38mBHXtO
9TP37JZmfBF/1GuHbdjGfo/JAlb3V/iNt3nYLylKL8V1b3JUNzDjDt1Ms40mOKyQ
mCHd/ijt0RxUdanqEKUGK3Nr8cBPHYDBbneupZjhW3AufsMHKG8blU8vdFWoTwi6
5kzX4WqETxRnm547lP/qYKjsvEM9MTz+w4priHrTktsjJZGTGrfsN8+KynpVvP69
f/AZ+E3FiIau9auR7Dotj+yaF5+MCUS6CecdAMI3sL9Xpc6pWe0SWG27fu6klX30
TsK8dvtxLYBaOEhkTLQoqEOnDrDrwfFtBgExpsWJguMf73UbVFSPkSS4/EVbhENU
QEgvmxnR+YihsiMAu4x38lyaYGZga2N+kSCmiTuuoxegpXNv5FpeGZZZLyAQmn8i
TOQcsvawf0DzdNQkFv1BPqIC8FYchkC4PK4EwAvH1tirQnIORjCpggXBbz0de4zB
BG3/2zxgPnuIVsCCHCTnI/+dLFDZhqbZ8QzhiMxAIHEQsYOAz3f9lJtF82yyO0EO
FLNxuocoE8Qks9buCk3gfxOyK+rsISPyDpFUECoIpjcnrhXpM/firx/ntfRJQJF9
Yg4/ZVRYLkXnO8EPrVgj5A==
`protect END_PROTECTED
