`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEK0Ewmu6W742WPRMVuDCluFOHWiyXPqdOC3xZPxx+kw89EywsD5jG3yTndgHlAu
ZOr+WMSi/fX1MH8Wh7JP2r+eKdQaRm1dB60stZGf0BRnHh7lxxsoFnZx/JrZiGtD
SVG0IclhwXpdI4OVQHCx0f8SbQrZ8Cv747ssV8j5zmAnAG4SRzD0R9/ZpohIykp1
OtlFEd3P158OO+oayhqWWcgyoqe9RW84XcRbwjA4lNpvWR8ACde1EoJzLusHaVKk
ifksd6mw9iIJk8y+fPU6dDnHq6F9MOi/OGbtHGj6wFrjDdBZmNrnySOejVUXjHHx
syysKFpWZJY4Qc89YqicFJk5Yh5JEFj/uVOOZqyd+6Ffw+9t5RfuPLMeAQgjlA1j
EVz8floZO0aQ90xqaCn25q+UXSh93zcrlymiyQ7TpIcCEFepfQB4f+b+zJcUgt9L
cmztaOjA/nbEgPfXNE16VdhGZ5Rbs8lPQMpSfbRJEeehIWf25VS8dCSlatlR/JR+
dTToy32gpAr+4Ltt1IHR/UYbQqvq7a3l5RkFS8QXGjodopWzxPj4gemykn9DQW6P
L0J6lbNqM7C7IbUCeVHDbjOT3/PgWUNnQAP4xMyTpqRTl+ObytOJfksaawaonBaj
dMyit7ItROuZvm1cgp34MRzhgUsac4xNkeWyP2UQbeHf2F6Fi8FueZrmojw2wjEb
cN7GzK/G1dj15GNhWRIgasLlkHSUQ7q5di7hL9ElFPpnKH6PJxjV5+NYkdmdwrpY
AYAhDVKjZpH+dK0iifj0MM4r+54Ox4Cmx3D/7ucC96G8rnroHdsXTaTjNG3SYTgL
ap40rDNDGL6Q0TX8gjaG+mwwCnpLX/sxst7mBdnIVESij48Ko04+Jf+9CQG82rxR
si/LJI40a/b+hs53Zum1/sgpKCmny9yJXpMM9soWd31jwY6URv/sZhMLjlEuQPRE
CDTHY8PddxsWB6KktEtcj0nASfBCeTaz2qfa0Wl/a0J/ylqXVr+/K2R3BaHGEuqH
c/Sa8m8bWw4NBU/zY7cfV9S1K+r14eKBLk4dayZUvKS6KdrhCRvyd4cM6Wh/cmZ+
dL0A6roEmPxdJgRwQJXT2UT4IJPdOw5WEwD8WWQlXTelk9if8QB4ydYSazN/FwD+
rlR1lMT2TQSEF3kgHONlWoxd6pN9p2FtJiRQ/YlwCzfP/QnYOJVIhAGgZc1+Lnx7
zuw2uPk4vwzUOQOdum8DzdkpqWuvrcHN1TxRsERpxOkDAx8+DZo6hX9uXH01E8J2
yK7Sl2/UnWMamkXE5nVD/9cojMaMbLjUvfwHMxAuNwlEK2G4S2a/MxuyvAOUrafW
H8rMzqtfKpbwZtNRwI1ZHhG/SFkZDVrcaG4mwhI9DLgzMdOnW8U7XBIvli5WPuNT
qap84Az0ZUdT9DBxCuQgLMFbUm8Y9pW3DixgCJb/wzuGCFK/he1Y4oNJO2p8n95n
`protect END_PROTECTED
