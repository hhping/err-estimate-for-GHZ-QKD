`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bpHijiKKMCfFr+dYJVG5SKfr2meaELVbp4B95jDqGlPAfDqclwXrGsvFvHQa5K7a
8MoMJA8ABgzEjprYFcocwlAgztfBpaYbQezr3otxkme7pbdu7MZ8ORV8gn7YexLo
irnU0clB1Nsd8OjImFffWYEsDAGkaWkzwmjlJ59CtttCOLHStekWkBhUTO8nuxbQ
8D7i71MOlnBjUNhCdb3LmkKfdpqGVgeOChNBZ2Oo/xjNTrntPX4ZUe0q9dDKYr2e
et08kGRfdDahfR466+hKtHkejuFisGpbGIzgr7f6nr4CHcb+UP8rXqyzKKXjXIj0
DoLP5wsk2hgEuaVvsphyvPbLHLj03mBMoVl95CbKrwLSndaSR00UT7HZvoBy9nDd
esYWh14OzQFLqungZMj0gWnG0dcwvl0yGbTW9qIeQd8WzTdFTN6XYwlXjigLNhHS
8P9Py13+yFy+4YygPbtsD35aQkMMMbfqb4lP19N4NtWMDNaF4ozeGeyf+grvIfjB
KquO7YZCM5UsktoCjLCc2+dPknG9+6SSjyYoOlbQvM7SSQR4BJ6FXDpp7p+k4nBd
cbiEuFJFy6NAxeG5YcwZq3V0g9xpCXAgaTj+9wHTsR7K8xpC61qRrNwggVBKXEJd
03SwfwIXHLZeZ24RP7Fa9Bc2eg9AOqt8iz/zuGtsjGP56yrDIkJ2XZeq5lerlc76
3z9q4bWei3P+oeiQJOBqczBd9xEcQWiN2eTVSu628ncCeZXDcCIogmyh8VOsLgOF
yHFjQDQ/kUOzuClRxeQciQxfZTmgk3xnflC0T0CBuTRjlhqIhTC3cK/pOm6aFvPw
9YHukyqZHoOu41CyWyCWfY/G8k1mIPBR2xbZU9JfnxGYg1jna+27vzv9sfog4TkR
OoPqiR3nLYMvQZrL2NtwVWOsWlg6oF2vWHIan/usJmDkxoUFZEDadJn0+fs05hcH
UXrWFfWVQsXB2fEkVVvYvuH8xFef9t4Dx8IdbiEbokI6Rk0JeVCnZU6TkDoNMP76
EtLg/fHsL5f+URB0OJkPoKQ7k3ccFShPPucQEyHKBGGHp+tvr7g7tYLI3/UFB44G
ke5g8U2rP/gc/W1wHhJMnJBaSW4A5M/47xf3m8gEAnLQELXgv20cXGG85RkW+WWX
+M+huBgTecxEp1OVFs4Mxv2cNqc1uMV44bxBmpoFd8tBDoBR+iDZnioFsMh/+OsX
hjDG5wcEu9dOfGFW59YTbLizwW8ugmTwpkLBtwgaN6wm7YnGoFNYawgei28BOSKC
7eJUuP4POinXx4i/t6EQfem3WQAI39zb1+DTTDwnQOL7kSm2n38e1KzPKCIXKeRz
VAcYBAopf+t7eVCFuy0ArSq1ikaW03fNymLVIm2kj8SWepkfGKWs0gTJPzFvepDC
LAI0QYHx/Lz5bklN7R9SsOevhkg0htG4+ijzHwp2AXp4bYqUZN4SqJpYMFWa1Eu3
61PJKGKIEyN3m+6f+aL2/YWY5f2G4iGfOqqs/vbpHvKpWTPbJa65zWxSAUMdYtCe
3LlGlcRI3ZEKHTbFhTeJn6ruWmru0pPZbqHHruhGhGK5h14Le+yF6RrC6K7yM6Ru
DiqM5Zn32y+7nQvNantTBXHPLXenAnlAo0VcG4/gU6Gas59v9ght9cyzjnW9IOi6
MgLqy4sAFPSFpLL/UUg8w+unY7OFzOXb9WA/FY3D2OT+M7VJCK3bqwB8I2Kzrg4R
pp7enTWSTpdkNIJ2A1VhyGugZryc85yQfXmyP4ISm4+Z5grlyylbs3zSsjUPDQhN
W2zh4HX+Ea5ZI8HoOpEEp/KRPxPm9mi9j0Q1HKprpSlpoes6JiJYNk+AznJeXMr8
VKA94KiQMNgc3v5Z6jiMgP/a+tmgSULhFM/JcqHFkc8qyWGpoN9IDgSq52u9A8Mz
kUvdPLiK3Aq6nhPLPI05IuJPjLO0fGLmjcB7JrJjb1Q9/6YgoA/iGg3vM31BcnR6
pEAlIcb7tDycK52NgEjPIpzBJpHc2whvi4fSv5bUkgh9xNj3kpOfSL3MTK03MpFy
SgxgmuOEY5KOSfXn7Gh0FUDEh2/aZWN0kt+BqlyxEQJ1Kfp0XzaQV0gqKv9N/yeU
nELMDH7M/cmfEcpOpshuUL2u94mYSUCuaVBqjY4aEl3c9AxKMezzqqJ1hzE7Gdiv
Z8CQTQyEkL8iaWkvD0jXmZ9iwkkhTFvcvFLgsosVn0AnWovf+UpPy8etYFgJOls2
1CAHO58QKmTtj/LKh0+i3J+QaIBPFV+sX3UgxYcdeqKfHfRNTQID+tWmliMKarUY
CThVQWLZI+lrNE3ryyB/M125+gk3Qk+bC+yYHQ/W/K9ASPwBqUYSh4RRxKnoIL40
QgAk8rRX3XtOZflZO8HfRVAi1PUR88BL5JcUEycYtDv1XBRHPOpSrouwvVsOzEpH
oJFxoNRzRXIUEdqU2orIKK0S95CWI7ThWvrAYmRwKZ7ETAXIdgE0xAHkW8hYSlfJ
T2lKStqKI+5CIf1qHasjuy6OVyLGsCRNyalGJGbRJ4I+zVuczCZ+ZKHLF0BjrOJf
`protect END_PROTECTED
