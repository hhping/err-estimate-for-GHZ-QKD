`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8Sv/8CsPNxk98JHEVhFVFFT3o9x/Pi4KKB6GnzfTu/F1+/NWKeh7DTtFF+LEcRl
bZFx92+o8g+Jp7WFBynEekIq04mFbCwJRnww5PjyqwUm5dUDFfFpaX5MGjWj6VHS
/dxvmmpQpCEyljWXEGtRgvbt96WzV33tWZ0H+OoT+uSC9Kj9Env7OaaE5nuh1vep
/Ya/xPUOw7/9R5Dk15P2Dfp+HVwemlv+ZjLnlKapisUEcV3UgkHZGx9X2TkeeEUC
hpe6hBxdQGihZEMddd6Mp5801n75WshkUcKrRtOap98OOXztL+sX9kMrNwKyMgkV
viK+mqJmNTbwb/kGm+Zh0ybmmQfMKGSwL87FmorLnzbnHDcx2Ypo/SicgLrqhq/W
7VGJhyRkyROcIHKjKwrEA/bA5XPEYWs9VXDW9Jt78cM4OTxHUwtwFDG+/H/RJ1Ft
65Gb50525SogP6qVIdpoVGa0nEML3AkuOabIAYubDB+cC4E3PgFzGR1JDlN0AX6E
m5PrrRelg4bTZUg79pD57GwFcwn8cjZnGMs8N7vo2aRUdYQrw2Y5SFQITvTGnHl5
BVfx81ToFpKhhUJSjo7oWa3bbdyJF0LUsWKrRXWTL1HkctJPOL6TqI8OdOKG5M64
WX1bToP2pxOlsr1yQUrHg0G7StDAtO6Mo9X1Jo/9NRKwoh+3vZwJ8g5IERA+edgR
eRqDltfy7rqn9akpdJuBia8kha23LV6vHSRECNx/DS2uc5NoEGJrxU+oUvSrBxho
SjhPLHHyY68nCsSxu0sjpw7Bt/hrj6PVDoJaTxayWh4ZtdnFhgOQXPRzp1znpx+l
6B+ta6b++bjjOicvjuoXe/c6jBHCy2It2tolUqNYaQqonrrE85r4ywgH8ytA+G2F
UuveruXJARKYGBZb17zq6wKK+n5S04eVaAIe7pXXygSnEGDutebKV/tSNSy0Z46K
gWfGQw/3rB+Hlu1P/9n8YvrVE3fZRQn59cyXlfd7SrTFbweRQN1/OT2rafsa+JWt
FEq7yqMaC4+nirx9LpEn7ie377rw3/iDaq+bVw8cBRsAvxBA1ah47RVA/YsGSQPn
KWT9fXYUw/3mi0mGNpH+fqtpL7x+9FbcM/nbaiudPjUJFidOmhv+xrfXp/Js3hI7
ArN3OW8+JVCOMb7cZcexrxmACcq2K4hT+stJxS9bvtOLlPc6U0gXtkIexWfX4EQb
CpTJFp0naDEAL9gXV+1w1MGAlQ2/ePW9Fgq9dYN7ngGsdimiPIIsy5hDhhI7sJ3e
4n/UkXgUPVrwxis1tJCcsVsE2XJVS+chGaVR/LgajZLcrGJ054j8MqBUm+a/bG8e
oPiHDdZGVNJbDkzXTjkUcXmyWU1k3taJMm8m8xN9b5Daf913iG2xBaWlDTPTGKVX
p+4OThZBJ/WDHfMS/JmdEyUU5pTh2zI5E8ikXLfsDrIc0OBPFOyot7/YBa/WT8br
PKOzfPHsThdxyvt2oayt6RcSo0q/HvbJk+4rT5szFD42CcVgi84ZFugUNV8d1gnK
GgGcQ917Sh5vFd7Re0nm7+zs9jsVS+LtXcjnOrGtrJk2WQH7CUPQzkvL6uJ57u7Y
knz4hwSEsrhbU79bNikrdEY7+nzo4cP/hLFBlq7ADpbmZ3tlY854Y8Nio2oQGx9a
J7PjlBTyPkGdnUFd+EGC1LQVXsWzNQLfbVQhsebHZGy1km9vjmVPF0WqK9UiFFEJ
CKgC83v314hkdFpmP8e/TjmuE9L0nPu40rdzofRPR7LJeKLXP724hrvvHHb7KM+1
DE84gd17hbMVLjy6myJ9TZ/9CntW1dfhgOLYzPDfErHcMmVx6xIyYMamQ4nb90bk
XjaXSu1JdthBUnRggb35hcMixYfvDfT/IY6Sf8iJ56JTTAoeWd/KcfRuMVjmmu0F
8USvsJ87kkAxwge7p/z+2SF8Bcvb9hEtaywB2GDU44vRCpeA/KOYE6S0W4pjCjb2
qIuitrKitdUkATojRTFQFzrJsTgJI1vgM52NEPt5Kp+Vea02AmFGsIg5fvGUpsAz
5R/DXcmvpR2E2TFUI5m+T4AaAD9wLYJBHv6kjie8RQw=
`protect END_PROTECTED
