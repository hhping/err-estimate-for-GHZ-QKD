`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqseCRgaR+/93n2vFexDtFegjvQZx1eEBVqr5+DaLdrB+4qZW1y22orN7vSwoyYI
Zq94YPcLM+5Vbvh6s1gXmMMEjkX73zuB+Qe3BS3VWTqqWCQwO8IAKahtc7iwHJC9
5GNIGaV8cB8GmfH0xCxzbdwd+J7jGbKfYAwhYOhDaMg9eaK7tI4jU/lNqmSdz96p
2CYwc9jtXUalYP+bnmGuU29+xRIBzWJ4OzTtTVQjvtGFn+WAWcKEYSi88yCRva+u
Z8kAg9M8hEZVb2Y50QVxv/TJB8qlWMj66ZoNH309x3fyrcXG9G9cp0DOi+NHgNpo
3+hYzXCX47d3gQsWelkPdYUVOvnTkYGTusnLds3jvwi3jf1xqz9CDUxCI0Behksa
TNGU2Aoa6oyTqqxU6OouATwdhxdPvONSy7UbND2Fn8KNyt3HH3UJMTmcVsP2Kpw+
lOGEH7EcQu+MQcqXGY12Zll8DfbgkTUqI2vexh/f8mUlGa1BC2lwDrUyJNZ0UkIX
GoxYc4OaWHDKV+6ZimA7S5M8EQMiKjHSb10RGyA8Hzx32j0KmJsryOUgd/HycEET
/WX2r3RvwHgoDGyaEjsPAGshgdrPbbY/fYe2493hgTnCJqN6oCxVUzvVZhSXGq8U
KBN2BmeCmNvFsZau9ls6vNJNjP6iBS23JTJR1Ed5tBkOZyqVXE39tn9Wux3x6G2L
Yjs0dq2JKjQHh9W7Su5nFzcYzEy6P7iy6oB1Zj3X9iyQ1w8Qc9y9SPYsc8JD1cY4
QNqio8vJdCKQxQHjgpyxgKxSsTLpBsP0xzjzPdswBsnmemxmI0kKBky4uAiJwy5a
23cjqPudqSs7M0U2eEwBDs4IY995k8C2BJiGRLvBz2nBG4tVtmdYBih35tZXCCwL
su4f/SOIG9JCv2/GFbuXeVxWc1dFxxHrAZ1U74HFF+G3bk6hm4Ok4MfnfZzaa0cz
zolbHDJE9U3Z0rh6j7zdlHxCYfU6Vaa1jeg1OopjD8js9XP41jJNeK0ffU9ENtAJ
6LxW7Cx73cIyEvr4jspJduR34N5xGlf7KLZlz0FFWLsDkbh7zVcb0vnG/eS4GKD8
ImGNSSNtfhWigH6HOwllkDe/fMrvLafursRIPS9NzQocf4C+qq/BaeV4Mq05AmAg
csjfLrIb6YNx7Y3n7m9AJiWxPEKAFEnW7HAexeCAI/ejfrxNP7i9t2H+lIrA+kJV
m+RbRvx/K2mYltgBc6AyhH0CHBej0i9Q5Tlg0H0LUIhDC4d9IUKfVQNtNDhEMpaE
M2s/qfTqibTBDPV8kdoN9WHTmPDoCudZbhlB32vIP+bxO5C6Mc3YdN+8z/9PeN3V
l56j+Ae4dtvaO+nxeHixZdRoLBUBUZ9unQxrj6BYAMif5GohCDe+DtE8AjPppdwh
5LMcjMnmLMtMH0BmKNmV23kn7fyE6rDey4kY3bh3I1KSnCk1mWhN0TFi29WLeeZn
oAnkpJJQcPGScH2HQymNQrrcM7z3RVYms0nUL7ombPUtOezQhWAGjbUAoGk+n1I6
AC5+4pd8jdn4kEY5j04WAvecC0rJNswlinfDBz36DDuMxWMC5YwVPBSpBFXT+VE3
L3MDAsZyHInzYgpi4y5LLv1LOp1Q30ysqBZ08z2RU7qTq6fxTciuKB5Vi182Vi0y
LgbmhgcQls9kHAf9eRNDAxNumx+hthou8c2JDJE/sd3ryCOIk4lCEDSblGaU+yXq
QYZ3N251FlxIvR1sj1msOcAA6fXmtGe0cLonHXGii/yyI6grr8zXIR5TCgILqT/L
KZldlfBkD0UCERJGXsN6IZiYOfNBM++/Wa3BYw0fjeEei/ibWUDqE+fRPvgH100V
SR+hHdQbk9MpsZdvpxuEhwkBjh2jOshbX7xx7PqA51AZkM+sE8ZtL2ShZNh+ubPA
zxpxnv9OfjSxycElNYBy8S8DoSAfZK28MLEp/5IzPUhkzlM8ymDSIeThC8bLBp8w
9cF58+Gua3TRF4ldJ33xIN4k3Txr/WyV2b9tqO1UVmumYTbncHwnTKSaTNFiOWAv
Ep/GiJ2ZMIjuP2DKRzE6L/tIXcDm9U5vB29kd6NPwqZ4b0nF7n0AJOaoEYFt9s3q
AO/avH8jym6x4PssPwtyBzc88DP12HO+TZ5iwjv/pBxzDONNjIkOv5sQ7JP2hloP
BP3EF4nCEdOpIopTubhENl8M8gPaNa1EZON1UNcwfSCMSYRLmGrjOIHKioMeMQUY
gbze4/YhkeLoykwO2mL2669yJCz1bbB7q6GVWKQMwlf5qZoFyGQapXgIFD8+8OUh
xRLpPGtX/toAFjY4S4gA/r2bdngFcG/N5gnaVrjueTWRaeVk0uLljTw+CqdUxl6T
/lhoWS/0y1dsQbncAi1w+1E9YvU/mKM02IahRZ7CZzmq4cMXYQo9dJSCQgYtNeav
JkK6a33I/frDcCsQNsCj9mbiEusfT6ABtXqs4nRn59B5FyH4/nB0W++1kHOtWmVf
EpkkDOkP5PSAVjKKyzkG49pmUz2TH3LfN0/ZDCei238siXRchhEiZ4udCP4yp9SI
XUaEor1NxBtuNQKJpf5xtjDaoIZTFMBeeNlj9T+UPq8OACAHhsbsFrHycOe96CHf
WX4w297FAfe+mGx4sOzb0yKxWq906ix7n7WIsqYiFchgwR+c6u0x/1CYKAw8zXR5
yX73oBwt+1fH+ILhjBRMcE0KszTKoJfZmFxKVTTb0/hV5XSVRBxdvDQg3Zl6AoaJ
KIG3+koVVrSzEjOUOP/0WGphz/l8NjzBPS7EF3BhLvmuhk/9Db0ZhzimyE578fFe
kJUZyqPwvdtpFrScI9rLEcbRjwVhPj5OHwYimYIwC33Fuym6b44AiBDZBzGaJ1e3
lLoiPvWcF9kR9kpDJ9knvJJtwsXQvo+zI9hw0mCu16rK8hb8v/Z1TXFWcQZYQUY5
fLPW9B4JS8Rj2O1rQJ/Q4YreGh7OUcV+Y+Gqha3pqeABkUCJD4zwHjjVMuCQIbsY
QnFP+dl2Zxod3hT77k5Notpe2xDhHVDV5WAoIzyGgkRAozxD1VEqkWX6HODEfRTQ
rw6DWjJl1AZuIZU/UacfxKZupohMmGhQWafUxTT5W09BV1YmYJ50ipSq+3p7TdoA
Qolk2ku2xNVVt4FXqMm8RQM7cDSodRYnaGokH3s5RvnTWglJ7oK3jYZWf9Gl4vK/
LO+V7RGMpjwhEbu5ImINoY4JaZOnFcXifwbewvZTQx20gyzOGLTlR2LhKJ32YHMF
EEjM+ujhdzmj9y+CnVg76/NuYYtoBCytxr+4nAR0C/zpQvgrc9kFy/NJXmAOW0pE
S+kOyflDS8+3LZUI987UF8CNNSESLnIINPqW5MhOfpL9ggsqjZM7+K6e/D0bFiQB
7gggxDQO7wpSmi7iNZgQVj9SLzeZWd09k1YL/sejvkKkagc7gwx4kBSaq80IJHm7
IL9zWJNQ2n290PzCcE2jBJL79TRXy3J2SMGdLmz6kROb4CbMt8PcYQnNW3a6VqS3
cCUd5lwzcnCCpHZKLglJqr1eOwO4VmEPygeu8CDZh9vTeBzEr/frJ7faoW0CL0vV
ZwcqMtWf5F6SpU3a555/7OlkoedOGw/tPa3i4ElflaeA2DfhI03nM1XddnTyAlYw
QxhTga6xLDLHZemdvp/8pOSIWX4FQo3HC7u4up+mwDatik9Pjenvk7F2XEyN9LRX
HnMYOykNkdIy38iiUWOrGz8YYgMXcPCqwsh1eDtfC40=
`protect END_PROTECTED
