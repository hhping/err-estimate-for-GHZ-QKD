`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jB+qox6PXQxXp/p525lXH/xEmZgjUCLYHOfJHZ+eAoPkcSqK5PKQfKu7JC+eE1GO
HEe5o4C1eyM2QPKHWjAdfAh33+0SB6z1ZDpudP7OcNH0tOwrPNWESVCE6lcb7UQ2
41pAetdd7p3hm+2vE3+6uPxVKxc0cbu+o5kafPBgjJrG/SVGdsiQxKy1bkQQEgkq
/Ahrc/KiwIuTPp3+TTvfOFmljtB2lGMys7jtahQLQ67u7R0J1wB0hj87SjSOko27
MDXtgYRGS8CLCsSiApDa5Ig7uNa2ty8jq6PlFRSysGVyHhkMQpnRAAZ6d2FHtDki
XaQC406DjWO9yZ1KkXA5iNFWzz9SHl1rQUxgy+poNkRElToZO15bISgyfnK9TXJ2
d/2d4MFUGBrbgJ0EiVNc9pSII4TbC/cvkaVAZ2PZ78aGKP5jIyfNN+2t0BIQfScq
gI9v5//cFbzUIJYr4OnYomqKxUXQydvYnFA+Nex3KH0Y3QkR8GZ07P43lIGJSy4s
04fg4XYMW5X3DbseY459kDZ+axz3Q1xIJa0r/vtPBslUvEz9YXcB3VD720jZVM45
oW3si//LUKFGzzleyMjROy2xWjdWDTSkqzlvYZo0oCgqjFmjsfohBNj6y3XHwb0Q
Sf5HvZJluDu3rM9t1DT+cvBaDpfsMa6VTg6u8GepHIjD5MfcOrPf2QX7GkS1hT2E
lqEEXBQyMYj3knlR94SG7BKgOWlqMJ5Cc3S7tIKzxy+fBfdjPUxbGPoMPrBPzITa
v2VHyrELLMQzpPPuauT+G/nklB9lq1aYL8JAjqdrjW3ryze5Q+UR7+TIHQotgymc
SvNaOZVLEULP/8G26azm97gdoWtzbR8z6HOHSbj4PzRlAGjvpXGWpM/UQAn22V4g
unj9mAaXa17dm96EDdA7kX15GIxh/HU6UOkqNaniCXA4gNvEIdhzn8ncsFVe4XGK
7s3eGgRoPzwvPfPV1Jur0Z95HHi/MvNeQC6Gme5ZNUMxFssTiU4GSibackj7pQlq
yNSQCJR7Y3BfOG5vO1OW8VbgE7yDW+OT8c8fFeq4ioRVcBt9XrL328hpdn+vd1I/
+MyDxrCPJ/VPfS/kDzZKrRcj+4Z//1R4iXzGFmI0lHENYgI7XRlsMh8wguLPYRnL
Atgh3wE7pW+STa2lfLvPc9jnbhUjrksLUkz22wUfHbhEsY8+3vUmXaUknqddjV8K
eaO1EkigG0sa6C1imfwbjYecOnl1STLG6CYJ42kkvmCMo9R26mn8s9dWJVq2jQyi
tBzVgrw/IExL690HrRsxOfBmZNmxbqyalvWsAXrpSwRPaKHsyqqk1vgikD1qUhZM
aDNmkGI/TZlDUFOHwudrSrCxtqG5oxMWbU5DbdgKv2usKPynmGlyE00XCD/quyyS
xWaAver/eZ7PI6Vk7dXf8Xgr6z+IH1K24tCiivDUgoadTCp420ka9mrGmZVbt6E1
UJV2EXOWRWErSag9uCxlydylb1Q3bx+YQ2MpEh0EbJR1twgk9t3Ckl97LyZQe259
Gha1Y4DIOZOFz3Ho/mqgrz0IXhn1aoDv+Zpge1fj5DeRqm9jigSvqAbgvXvH3BXb
lpK1eed4dFCKQtzwi7ct+cL2YgZ5J0EK/CyLnxbg8U+euy2YFkozjHlITMoYrlod
ONE8nOQ+F5pV+FCKOTnQe9H88aabGUmlOjRjeacFH58fTkvjrTjz19nQTLwcoQQh
RTpO1sd5f/2KAV+ZLHikUQ3uMo2pke/Ci0+b2hRmwqhNXugOJZvD0E6g7fDOyoJu
bJOM7o2BUzrGb3U7Ejax+1F6eVzFZbwQlU1hKvvTVvtqrkQY47obRfSXckswXqua
IonO+trFFg3EUb7hCPEvycgJ6oc1aFDA3+t5H55eiXcqCiMLanwNR+t5/GopMsAP
d1iLvZzr/yuh3Vbq9vCVH1kmohHN/oWVSsbZsllppRU=
`protect END_PROTECTED
