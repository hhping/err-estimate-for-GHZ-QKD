`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8Z6npHUHhTMSOr5fN6I9UC5ro0BEI0ZsajLpWFCZJEgO2YAtUur14q2uW+A0Nsz
HgEoj+bx21JAa6Fd1BhZexHvqAXnA6ZSq1mODHsRLrGGdoBoGkLt8wKUU8i3MPax
q1XEBpSP6bzrS29T7EaYelzS4LD80fsy6WwlbiYN14ewMEibYkwAH5RpJw8AVcY0
kHgoYIs9f0c/aQvXBhWDu9lrPC4YFUMBnJ/LcTDPSNtGDk82LCzRP/AnDBI1o831
mI58HV5Y3R5w6rB/abstpYc8Pj3bLfPI0ouiY16fo86GzOuLssguVTqyIjj4r1s2
iURreKOp9MBusLKzP378P8fa68yWmmkCEodU1WSC2qjEg+4IRn8gQ3UoUTbkemTS
FQA5+WagiIzIkDeeXiOrL0iAFuIdrnhoGczkFsr4I/w52TLh1T4PTEmRtTTVQwFT
i7Q0uUJjCuKTlzUmjNv7+w==
`protect END_PROTECTED
