`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Dk/QPs5Wnn5/oGQe4Aybi5ieyktsq4lly9KRlDNqWCvc+C9sT46yBiY2tx6LpEj
0g4JOECQGMZDPE4hniZWAFtKVpg6cwvwxjFaw9D4Bf82KvynZQdk2uRkdg+blhi3
Xp9vQk0l0MJf/ZT89QFW00PheNiMECE0EQnmPLD3gMglWP25N/ahCPWl7vZZr3EB
8SsTRc1/qs7yYLQC8HqJvRaPiAxIUKbeRuLXCg++ZtPL6OTa36AsSpMmuZ+4mPdz
4LY5OdGm+dAfoXs27XPa9S0MFC/fxiD9MPg/KUzyv/1oXNajNaLZ3zPxgl4WJg97
rjTLc+5JkSK9YT6ecdX7L7cbFrYZ02y/G7yZKuxziMtj1CBhoFp+UE3iVt85OQqr
BjoRowN5FNhIGGi+RxzdfkRIYlqRrP6v3+H7ed5TrXUJAr9W/uWk7XvPZWtDSc5n
x86s537jbu2ffojWqSMt42gQTR21TDAm1FiAedPXCGk036AKDoIF65VMwWXH3ivO
XdPSvNS9e+S4Nw+dPRISzM3SZWssYXCSIzpsm2qw2PfAd2V8VrpGG2FeUGNwJ6UM
Pv1BpdF3O+RzsA4LlozFku0v93tiC6thPrbO11ZDZdUJZWcnJnDIakr2uxEiciJx
8xTaNAw7TwjVqzU8XVHkYb6npEZ7kkW+VU7AYJlSD2UgMC4onK1xHtbQ+8hjrJJk
0X102kcGFgbk5A5YNfXiZCg5c0PmI88ui5vxi7NezEyICQlsBWylg+wBF9fBOOi5
PA+fD0OubNbxek4WcxDLBs0/lXn3E/t/pwDyFSuCRpSuhk4IX5o/7NuaIFj6jLx3
zhIgtPBj2CNt/s2ghG6kHzXLnhqOWYMstUGAOfMt+BdR+uOtkuH4KnKQGdINGsxJ
fQrN/OWRlD08LqE1/f4Mp5SyI4Hs46NHJpDr71l7xvvg8UTPyURbSrWhIftVyujV
kaHnkcxZ0zJiTemhf+nIz+8sgsX72KdwcuFQlGYK7YWIPqYyIcIKqR0WGgTl7ulQ
iSiFtrKjVOdym/g0FtZqNdPc74uTy37Op2HPfUf8iYL130rOzSmX9hryH5x/JQ+e
SC2ugqURXZan4DFVd55srWftSJPPUFekHwOOnskxHCe1PM8EJxjxqhpmj7XYoGWt
`protect END_PROTECTED
