`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJEZG/kLGOHqvQzOOYVMdOsd1uWpc52ZEGzoRbZq1GPkOYbaNFijUeLD88BdNy5b
A+bNvqyIHZWEB0kBDudzkl7paOm/po1/tk++TAHn//Y60WqwZnf5TWI+8hOU/Xhf
4wUz/WZCbX67hitrMhaBwLf1N2/LnDkm9wl88duIy9p3+Ned8JjudxCaE3bP9ni0
+aAoGraR2XeVwdkw8gSLXCnx5UJYGmKuhr9j4nVW3jWcECk/+E0Wzm1+V815ibyW
le7ubkfEobOq969YUh/i8ztR06OT4juOnfmkmgOKLuys1jMgcNh76JOGCyYgRiea
arxzq4Ksef4aOvpf3vSEgA+InDBUIB3svBJ2FE4NhDeRwDcYTTqxpzuJAx48lFJP
/FU+0QZEoaavIqKpFFMYJ77yQzcP3B9t4Cj+JCG9mLc=
`protect END_PROTECTED
