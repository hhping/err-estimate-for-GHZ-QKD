`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uaLcbcG7M/IjmwdnhlE68ucHGiasiE0cqqx4ZOB7ey68ssXN3JfuxLJKfHLnngES
6unCTt/TIKMN7M0S+E5AqWOFub5fD5CZoIW2bPS2/DW5/yzuFkPBzRa/Ykm0cleu
rUKf0U4zdpxVR2h7271Io7y0yyb8vbYIIPYutWSTNaJDbWBPAW5lZ5hl4Hrv1UR3
xYcW23y6wDTyizbb30oUpknvPKGPtszHcFxDqpw+INY1uF+4jZsoe6yIS7okHawJ
osElw6G/NxcVGNukP6mj1DJauKnKXggTk+3yRdtZEMhqoZ3btdDI8G+NgLxyR/RJ
TI3N3dEILjlGR8r7kb3hwlUK8Jv+rO6ik+8giG+bofsS1dy8oVW+gEKsve3R3f2D
Rd9zMJFUCVeDS8OBg1Fx4rYhsaB2YjY4NI4vZasCxd0VGu3NtaKWE94DSn66i1rW
EUWeZWb2/JU7fD+P71RYZmtsaDLC2HYwk96xDqi9AzZ9rNDMACVZ/QY+yJYytlFm
Zky9cVeKfDkOIbu04g2GorRX1q3NwVyS5VUVzpdA2Ew=
`protect END_PROTECTED
