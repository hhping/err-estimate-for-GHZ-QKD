`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HETYzw106CK6uc3LyUFQ1podEMU5kURKpAdjhOOcj1O4C+24vX9ho0L9J8E4QvCc
3EKxyuLDy9j3umlQLdMfTX3a1Tq+XwmHOk2nNOWmTpO+fCKHRWqmdeXsqcC8PJ4h
s48o1ZUpUHFhu1m9xYGvaBmUOvKvqeVM/roF9+JZzOvi8WMz6BomVo8BUkS78YJe
ySas/4K8oyLtBwIp05fN6MibTnpQ/+uTu78jp/w8Y55nfZ7UuWxJrylt4NFcD+et
HuuUamT0nY0av+4Ft2ESOoiQbN5/EufWgrhFQjYHYl6mbxWtKMV7C68ucFq2hv+r
iw0FaT7u3/zShD1Qgfc6amXxjNSJOKUB/Ycfb/xSxWuLfe8rnDcJ9VlwmYDYGtxE
or6UeLgFIfoedH3MOjyzZTXJrByn2mPDE+rVbKdu9V1qlCDKTORHIDJ+k1jFNkXp
3WjtVgCxnWRGrDBqIJ1jz5td6x+XW8nPADQ7LtjRgo+TFG0oxCUe/OdvzcKhtVtu
tqZxiZevphzSGGl/K89CGzUku9E1WpV1XL8HZVnUbnvR/zE23Z1b0k2fZGQrwuQJ
J00NVFtmEgPVd3NZejfd7o5urb1PRbx/p3tU5b6mCsb02Ztv3akH4j9FpaA/qCZV
Vt3MZ24DHSth4uUKdTu4fRXzIYZ9WvoO9vCc6pX9Ig/pqrOQkSMnFyjnTrHYY8qz
3WOxxtZ4kH2W7ZQqAnm/r0oGRMscAvovWOtDWTR+Hva0YTqTkeKnMrsygBRfC4i6
c54EFAGA1Zv5l4AXLkx4Wpjwkn7MK3oZdYDDGptQCjzYW1kLvuyGbj74EkDA2ahw
vYapCRWlfw0PT9oYgkY+jFMluKs0suu3UItZLnU4JSzOUoRs4kTcaeMv6DAyjM0L
2oMS5b6EbIsJQUrr0PXKI1X4bwitXL6fn0rVUCA5mrat5yTRWFfY7Zq3seHSv9gw
FcqAkP16Dc1Zjg6gyo9A/uoqvHGPJjStBIOFonFUpAQOROymNjfIsKPsIGrNdQ3y
g2fRxI/fn3a76oSQl/BhOixeg8nvRFC1yPrYKgJBovDyT3aNvsuTKbEkM/rtrLsU
17ltMKl75LJWYTk1J0hYEJ59n4QHe+bRjOAWR2rvtb6SfBtO3mp8bfCLDjFRVN9H
ar/H83oJgTeYfUiUROkHNMg0Po+zLEVKkiL0QgbquFiYytDrac8qW9cxgUnttP9S
oDF1OaPmrHaGYvPii/2WUZwcQ5RrzO6g4t9IxUW7rMQIEOO8YcKahrZwQGewkxTX
VUiNpEuMfzJU5g22iAn7HAndfOyHvJxgEAyE5zL4F1c+Ml/jDnV4e3LSQP17nV0j
ESTfCLN18nc6JafLrUwqfxdDTxQKagCOKaiFQ+5y8Ct5sDUr0RRmThJsRhHFhBir
1cwQvD5kW5OBFZLCUuSjKLagayRde9jIb2j2RqGVd6YI6JYmJjEKR0R5cloZkKYn
qKivGb3Y0n80GEVVqaXYI0wMtmKPiTQawv9xZYQi/UskuHmeZkwnNY+1uz3zsDBL
ysfzW6ZJVPXE3IloTgIDD1c3uxqTpgHtY8IazEO82LarP5L9KdMWNBfV8qWD3jvX
ve1hxKEueZqJNeU+aB7HX8RPdxChJRWfpQqRrmY3HZ3dTWwpEt9/Y5bp1sSA+XRO
TPJvMGhoOrLQHfqGn/Hbx8fPRZUnCZ1McT7+1v2OvUQDPdSHIGWkncDFz83cE2aa
mJ+Efhdkro0d/GldL6FFwgJM/QjnAT0dybnoagGO5MDTXhgu2Hi6OucnEtiJVvyc
6p57oJ5hiJjUn+w9u+gOiuDVr4l3rOCZhjRcQacKHUF0+1DGbglY+LPOWE0d2rgc
BH+9gRUdB1moTtE5Es6QYzoHIsxpqkVltiaMOg/I4V5aAomsXGJiFsRojTodm1GI
YVwaXBW84KvWNJj9wcQAM5ti9k3DN4Bba5TtxP6ejHFhO9zoFjlVvb+sVbgWzdSB
XPTMT1P3dbFMuvosEoveKP267YiSRNO+J6mtJ1pX/HLOPmlNUNJUctAjWGl+WSK/
4xqTgUacExlRqU84olzs58gmePgObLKHkp16Qat9r3v2+5mnKOOkb031Do5H0jnq
0CRsrz27GMFfoCaMpMIfFQVwwCBrBgxVxz9bDmX7J7HqRgthKkgoBoiIzIn0PmLi
3Vbm0dQmgeAprwFAjIDk/1hckD5ywdRpOhThwybxinaZsCNV1oBDpmmsBWE+Rh0a
0avIxP3qg8Cx+hv4WvcKhi3dUO57fuhuAZejHl4VTY2yA+ReaBrmjwlfFP94Q4T0
h/cnO1vb6lyVq5PeGLhbDcYxUb+j268Tz8uG0JuceVZlZxuNDTi++zipxkdVC++b
DZ1HzFkRnwVesf8fchctYp0ZQnZhYlg+z6UyZFK/TrnCQkojq3BCSfBX9Gnjzdb0
3gb9jyzTJgPjMR0gG5qgTNN8CP9yR8STniyOHTjLlytv8qI04rKejjRQ4dMh9kBW
H4R6Y99o3P5GGxpwiSxvAni/eQ/y20wEs1i68uRklhSp6dDaoZ7tiP/yVT+wCbDG
Ufb5JKfrwuyrGRImQzv1Vre7ZtvyyI38dIGqRjbo8AiN2+Iej0jWtPUBX6syi/ge
2dF6cggEMK83szXmM1bLDBCTERfDJH2dAUU16HdHXo97/B720Z98mquT3ADi5j1c
CMculM6HOfzslDFSaPdUqVf1/qTwxJj/eUbvAloaIrCnU1OjP5WLP4EDtjrnAtbA
5NSlMzF2aUH9bHQnKkIyXioXi9v7kJuC9SSs6FOV7Nu+9BYo2OcBPtUzOIgM4Hk3
57NuxvmpSDaSIlaF98vDLYH1QCS3AJYzHije1IpZrmv+hfjGFVCXzGG9E/47IIwL
qV8teNDGT742Eg06rQGzft+VFlyQsAkUR6pvv1yeWB7IuG+5cKl4chRcc+KRA7W5
MPtzF8BqMaRiqNba/EqL7jd9vfZC0fisymLwXg0WYg5PERk5JsfszpcVbbYykrJg
sVZEi1suBiWrW+Da6D51tjMfgZJl0FlEYn442F9xIvAKxwzOam2EjI9N+GQvOSNL
etn8vZZwJLIxf9ZLwlA/GpQPHwRDDUibjpDPJYMChP2U5oPBTS7IjI8PtzOr5iw8
zEGJepSVSCSjJjgO5UammhzrsSCNoECU3/XNzvCzOF/GEgQ0WdKKQ+i/YA1ZzZEE
Emq3aQ0VmaR0itmAhJex2xXGxaEXprAjX5L4cG60OHJI+ekScaYd5Q9dNwrXsj5c
dGz8WZRv4VpKXho+8iLuvantQSZBCibFmaZ/oAyWTjSJdYUdpLlSRAuiJ2i1FN2q
np/TbQkhMh4iHwh+1Xxe2Dh2bXPw8jo0tnO8ea5FC6NVehLTqkv/xGYuQBhHMZWv
/Ayw/VhNu5qpYDMbyt6EFtbNYlD3pbDHIKeU0uYT/Ih6dOQKwb8fO0yYRqX2u3w+
PHBQksXmnXwpZG5fLHJGqquDX54ssW+uGk1LwC2CSOznJsAp3bmsAU0oFi63k0oo
iwLHrQVVS0in5wBAI15zHEGz/NF119onX1z67zXw0kZ0452VxM1nTUxEBxOU/OZO
Fd+OxdA6yoWzO3CxttPBbA/v3SUWKBVm0soFLmYDozZZcDW0x53xi28fIN6WElM/
NtdDHWZDW8oyBIyIhvnMLdZ5Zr5HiPRj3/srJ/GK6EMgNQjismIQQaqoGNIXmNMx
U5NTnUqoUPYl9coDy9bx80vqtaGe4mykKIxDT/9Q/yNMU3a8vzQtUKFfWvgczfAG
dd5sJRsVg1coT3xWLntWv0NQl0Prj4wjwEjK7pxIpeMVZSgfO4/mufbwAjRu3g3B
f0dmIjdFOGkKCMHN4iaVa4zp/GEBsEro1SbNqI2LBgxX/W7pyNzvIcR22iBLT/AY
9XwHHkYNP9L1cUQ9m4o1kmwkYr8drp6j3ku1OxwTVAtH9cMWlXlgjkMOg5QeMe4R
qaOjzkaDLc9K4iRIIED9D39B8oUeojaS7f98JQNx1T0PEliwW/Sy4UnJGOJnO2KN
GVkiv4lPQUAVSz7K8SQl6BL27uFN3me33gc9SN3uMmPuSVuWVDC5lhWm6jBmCFST
QE21+m7EFuMTYYW2Buwg9HC5AiI9OEs4+QSa4+X8lf8jl7kOOD8xgJQcJ5kLAA44
vBWjRveRI4sx6tJ5EDtXZn51QEeJjjrNs9gvCG5n997HJzvDhzJlDyw2F8yWZbcG
hOsmH7zugq0y4b/DNZ8cPuaPgc8IDLZkd4QpMpCqksPPK/ePFanql/h5mW7QCXZd
0dWW/TfSLYFofnaE8PgZnB1LDt0kYzkXEs5K+eB8xHlduvV6LOoz9vJdcTMKTsLA
fAm+eAFPI8csad+eT0e8pwUAebhUQjFP6XGEbJt/L90W7ToD0zyKvgw948rTDexB
w0rtkerqu/3Oj7PjtT1Sxzq1TWitTNcG6Y50heGAfkpRc8H28Y9GS3o+ZjS2xENQ
5Kb8ztDzdAWsR/fOnpUXsI3TOJEOR48jMD3z9hAr16Ho0WFN7MwB5oqcjKNfmyNU
OlIfKwmlL+vx1V5xdJmXFkgfPp1decAGOXd24IUVnNibwLmGOjpvjpKoHPcpr2qo
dEztp+UkwzFnfUK+l8qvGccSoqjG/5Fxv5JMLW9DalbvAzpS+y14o0rchLBHV/Go
Uagyn/t9ecaPCIu8w+DQ6l5zYiCMRsxxNOri+5FeV9AA+cgjT3I0yYhE+sDfDsbA
YujAbeFP/Ij5DVpQaz6xx0F8dQFUgXo8e+g0hk5g96I6/cD0qwUNle4V/eO6mb4r
TSwrlwdEbap3e4z9h9D0PBeHxmGwrfirEOHfrH7cgnKuAfFw2baQGamqMtEFN599
15sGDEaMsn6giCAwQOVSRg5hRM9Gcslb7Z9Y2T6IwwqPO4lfHHITL6+hbmHNhtyK
TX2lbho6LTGy4mejUs9TzUI2RN4mgnms3FinKzrB0V+6+RDsQyL90vfDpO9Fky4H
+cf+vNM/RfDf7k1lGTZSRjRqW6Q4PWxCNLFNnpNKtZoGK3c/ZkcasFF/m+uSe9HO
c2Mvzo2+H1pk1t6jGwjbbbQLY6iefDF8TZAg/ecJqNRFPiV2EItbIHZLNtekPlzH
QGpcTe8zjdIQgoK4WqoCTU0y7sJhqamOjNAuPpfd7NSs9VwLKEXcDZuBfSYGqPZA
6OFPJz4wbObZuc/C0fTXNxQpk6GoYYEvHHen2244Y9yA9JiKlEZXQvNnGnfOpQ/6
v/WDSCxLNreX/ypa4jl+9ktg+ncddyV0S1jGByQj+lUSI0iA+MJbP4NuA4RAt5ya
zHpOBTbbMr1VgeQDpWOuNo3AvSx/jnx0Wy4QY2LPKTTpBnLeecOsU4jAfMfKJqv7
KUJeqAr9eb2Z/zxhWI7zo6RpVEpY0VDi2w85BoT9BNwmWPzM0+b2sMNUeEgi56GL
E6aZGaF4b4y9VL6znBGhXOIo02jGPt3SNEqEuNkSp5AvGqYKFZhKVQX68rmXGb/8
e+xL0MJwxlrMOjOMRTRPp3wSNNXBDA7qwGR9x4OVZ0TE6HBr3FPO2e9pRJguVPhh
4bKPk+JfELqWnqGiNsQYxLs1DpDJwU+FqldjkABLIflgipIcLeRkF8JTd4C3hoqW
nDpbry5Ljo2Nb6JOvzTXl3pxQ/ucWuzqhYdJlaApRso2wVm4J3qqhpBLuv7sATL7
4JFT0Zk/YxAUiu7tlIoap8/pMdw7F8d/pCw6ErdeUMKQNRH4Pqaq8Xims4f5sEwj
VN/LRn6Dc5AFiI45S1FqCemQjs/SuP7BCV3QYaq8dcF44uGpaC8q0tNhNBvEhG2T
mJNTmMn8UEMfThEy1gifGHw5waBwCOEJRd3HHuSI7XUpZro9G3PZdLMhUgJhI6lb
dY1L5bfihdyalUKDABncKbvupF1nlGAZz+wN3ihLWh5Mpgjq5BerSeWiHGo4G8h5
85fxLg1MvfwtveQv7k13bYQkqVhoGEfCcvsfpHVTqj1iS6eSiciJaByT+CEeMuSK
JxCGWmBXWdqfVUK0+dvdusZYVm4gvapskR+2QZWP3FQDYfj7RZyf4rjqK0CDjD3U
/2iLCi+u0U4q9hnfitJlSTEHkw7iazPFCLleqOW+BurN0ottJALGw1vuwrFx38yb
eiW3IXJd3SA2OpvF6chF1lX4wQ0y4fz9XGyjULFfCIkDsrXdXqsQcjIxW8hdYiji
PFP7kSlCU039rrL4oggW6GY5sf7d5N3KtR1I2PTBJA+1aL7HddDm32X3Q9kWiF4I
lBXlEiP68wPc7KK+NheYmI2ij8YLFH/JVI5HH1bo+lQ95NbUmoClhN83uRSQck4W
9Al5oIx+dc5+YetinxGZnzr7jHffnvBi46mLUIIpsi8VZCebktyj2hlnntRev1Pt
HqXEcqJ8nj3NS/ubQW/lokLx3mtS7Goe9T6NjRrzwnGhWXvsJjqN4pwX/J1Qwxxz
7o7Ri8x7b6PMAoS2GUgeu3yhUtQEs8l46xVH1IuUeOJsNbsSHQS6i4eBAhXq2MKd
kjTGiGbxbba2lS6oaIPCokh9lS+adQ/K671jAJ5oKq/DmpH8rM4bT0koXc65brL9
jxVNGPTP1la2Nu327NFAE4G/TqpoIVBxJOloCJDAT0noGFlUEyEgCl2Bu7fv+eLS
Kx5wvQOXIqUVQuQjSbSN5UQIZ1TXN8dUKPOPjfAV+Cb9feHTnZv48lCBTtTN9zCE
QjY2M3f9bzJ8VuX8h/T5fsSKPg+7V2XFETAkfeNejtTTearXjyngQW8JqNu15zsr
7WE2fgoFpwgJ7E+IiPhQM9Rdx5m4dy1oOWydipTDSMR4+EFOCMf7HvPnMpTGSJSa
EMt0i6ABKsPTXKEnR8tQG2HykKhLpCkIuQdv7CMkEuPVILdqoB7bO+xHPSjN6Ib2
ZH4IMFXOCsA5LfvjpUkHhHezZsPZMYHNo95ZTspMuNOxHGkPBZ0A9uWpiLeb3TrA
W0juRW9x9/NANfszldOrpMO5guk+d7aZILwEzNrvluXtfVCKy/AcOkoSeKkvM0yR
xRrC3eSzJ7KGcwOk4H71xkRYpTaASWbC1cFy/nE6L7TK8L5B9jl5hRibHFJavWnm
d6kjGey6cB8wQchHsM/TBw5x4bjnzxobSEdba6Wazj6FkQX1D04+0Ub76gsAiDKL
YUPO472bUcVVlpTnJS3HABMFVDbHRSFNvxiM6J3s6epCtjB1n7t8+xN6iaSQGSEe
IG10ZOg7Yy0EMdqDEmtBztnRIR5tMYqEQWqaZP5ls4U3Ho89jeRkVFmNS8pgyqjE
2x40JK07AUFG5T6320V38gvSdcPzQ7VWTWJJOSDtQW8cjg+nRq9ZAIT3Q1zT/2xs
rRneWcxpuHqhcdRwyhmvSIoXMYVhX/5zw6nRxnef678g94Aw9Rx/fNp5xSM8M6gV
2meITeFHgIlI+JrLoWXaiCxonPrMJG9gGdBPuqvAiAeJLuXh5qxpZq4ct9QQB1cW
wmzLd9yiiLhXwlP6dwU4deARokQ/BA+CcO/bn6rYbYCfqDoniZ0E8AV1I8RELqVu
SwT39SBkTKx34MmTA5IXXLbzgf/6EWFFrhOW3zXircUnvd+5+Dfhl/GYfPftEoUZ
b8oGHPKDZ6r/ORtOoGxTq0/J5+l4TWwFGMDuSoqryFRi9IO8hxxDl2GyAaWTzeiE
C6R02y3XgVl8HFNoW5TzKqNxpNzFY1UjwQmV6+xf3DZ1V7erMLSENKBqpLwtDLV2
SR40WFZxgZGCbCXH3caYbR8DAlpJJKAhDI6sm7hjfF3cWf7WYo0HcZ35gCRGw1/E
JmHNDDxcHwglfTLSb7ELHK9TxzSK2AB//PP9DSFzK1GhqwvuRTtTMBDzWoXLMuM7
7KaI9Cj6FjFpqKYoY+TRZmwk8ezv0wmtURgLubdQAw12PGOBw7Hj6IhTZZ9CwWz7
Y5WMxO9Cv5hUV8Y4VlSzlL1R7usTCB2LcqgS6/i7lApPuyhwDK/AIlXJJMOfE6Kl
a7frrUz0dzNiYnh6pw3EemxN4LWr3kA08GT+JkuLyS3rCtXeeUKyZfy5M5wl9cOM
Mt7QSzrmHbG6pfUWthJqDBu/9bMLSLHSM0mIp6DfZCLPg+VKV3wQs0c7FXJK6QmQ
KL/JyoolRGaShdPASTiPJvrEm31zfgcIE10d6cAgvr8i6N59rQfBA/JmOX6r84Nb
UDBF2mZ4EPpXNAFAFRaRt7eRBjbt6Lg0ajp6iui119cJRzb9Bgpyh9uqVMr9lRxW
cIYAvwu2iA5GTd4zYubj5/RkzvhBhMtM2WxvIjKimKHNow8sOS6niurxZYqsETAo
eet6gazUDk863ErvQmKNP2kzzKyyPtkzjYOVbgBeZK4jpu+NuTaQW+edely2qYkJ
K4Q0gEmxRGoo3jQzLYOV/WWox4gevlPBtdoS8OdLNpzOwShnxO+01b/5t/ycrqKV
jb29NDiyyRcu/GE/yR3JvJOiuE0gbXQyy9nrWfZW2G5vq1VSSsNIbWBfzwJ7dzO/
FKmFsZoveZl/wJqqzEas518INyJ1dr5lT7QTVuEuePWiAzQRpcbJ/wv17zCVEuN9
y6hXLOC6HPv1a/0JOSQTeubA5l/QsHbadBVLU/w7C5yDnjDimJVdYlgHtcziIoce
C1yL1Q4IY5eMsE8r71R4Dshx1pdCS908/0y8BPRUZ4yDFtWyotRug2ktjB1EKbXi
O4NyYLt35AbRbHhs054Iezhj9APjrZDqKnCxkHu38M6em+naX6GzviCy7aDBkIhD
4YKSCrUkqYaySIdUXuYfAFm+p+AJtaUIQGw0OexcA4s798lEUfiEyRo/gFZOgkAD
t1UrPIg8/eFQJb4VCOnQLLyoqkxx3ea/X2lQHODIoL2oGt5n3MaE2yAZqaTB2r2y
3Zl5h+kARkAGVLCM/nqme0lMilbTmPiwqSfh0tjpwtJG67Mfrv9I0g8b+9JbyTwQ
U52G4yBYTNzuBT06Wb1qPkZLz+aybfoPV4W2JsVWX2dF7Inldo3WuMaqy9MZoQGs
9e+xaJ9AcKtnS+RA8UbVtOcEVTSlrjflWmaXolfTOO5juqFhqCROB/M+vqsFsqb5
JDULcrU6uhgwxL58kAXbNCESMtV0Jf4mGxN+2++Bbl75r9IlTMhLaohUCv28c1Qx
dM/uM+yhHi8rQW8wcaGrk8xao2OF411XrJ0SfPalEPmN75+TEvz0HgtqGvYZPK9R
pL2g7x/MlNUd6tyc6/NCMN8PDZT+gzp51sHViSLVqciuxGZIN/0K96oAbD8vPVtX
2qgOpgaTiLwbNidUcD4m46AtbnFYrhEaQAOXVfAujQfMyazYZLgU7MwVfWx3kU46
tmtL6xAd31aRNs9o6udG03Kk4Az04BOxD5E9rUkv3uL3muYDQyUXCpj9JEO+9tFa
p3VSJHpBiKFMoTTYLPzvKgD6KAh/PbjLrGB8bplYqxlVGSa89wlgqtL8hVA5HhHw
GGt8MA1h1VPvwRN/a8SYEZQt6BbEvCxySKbOXUiIZm8eVzM3oYEY0B2M9ovNN5pN
NW74vVK6IOHnAQp9SpqhIra8ZcdISc2Qrafl8o+73XoyURnaK2ERyI/gpOstRQ+N
H0nQnTxxtAes6Hssn6ZvQZBmuKvbI8PmUJ+ju/7dv+g7V5sIv51F9yETXfjm4EG5
pcSBEtqLWxRANoB8pqltsDBnff3hPOWwhcL5MSvvi1xVDDtQWH9kR3bvBaqv7zfJ
ffdqK8+zozHBPRplCj8DTGzmEJBggncvudkQXXcfSzsdFrhz0PlmzNY+5AvRTE/3
G3ZyGSjRuKYcArlw/3SgMlPNMQ9NdnTp6YViMiv28afjQ8PlcJIlyInZwISM4X8r
aEgkOf9l9iOIM4kEGZ6A5qmxYKbEUbDEUrQDA/pOuh/s2X+UxTZb+TTYJrXZdg0Q
2e7GPe9t9zPULuzfK8e4konL7dbA2Y9tyxaTX2VIrdrtMES07u+K+Vr9AgcZhCWb
Pd9Ec+4zWuyCyjX/mtmRAbjZE61Z5KwNkeT5ijtpHCxzxt5X1NcXMzwTR8TJyjeI
BNm4TlOhBKhtNryy26ecwHhO3GWNdg/S2gvpUD7CyI23oCoUfDMN3I+dP8Csvq7L
Mp2qgI+64QilwJtI2dbF9Bdm7ITQcSarsh88wQqrlSZPduC62b057BnLrrieUz36
ZXQl9NyROx8c40gOIiF3B2jTj/egunTZ7A4sLls8T8iTu1lndSG1H3xOIrCQr43U
mGexgkmBXjYStSWnD5MaxGbsbTHsIpxUbr3t+BeVD/5wcZUb362QD39WDcidGLlX
CjyyeJ3Wva20IIJ5zR2ViHp/+hA0IZGBO25HlB2A03wE4bsFVLpFVgDqxxgm7+M9
8Zhmle/Jk46CKdU6kHIBVPLa5yB9sv9XMzOLFHvmeIoAE24+em59f4EwXNUOhM8N
CiD9aYIwavYt45x7I82qyNBsiZGdybOkkWDS7Zmk5xiXzn2EkMHvipYRotp5FoEh
vxXcp2+gggQHbPUVOsZvo+riaWAlNPqBxyb5LjGTGCISfaFwEUzQXocuwkGyQsqC
jY3Qig4SDiK36ZsBsyMOhwDqBfB0RfC7oxmiPfEriuxKk1e7zarOENmPsfw30MwT
y69BNHqVGeezftXNEAvMcGA0HVhRM2IEXPahdbP5z/62F67Q+hng3oPbosawVdF7
SQrvJsTD39sN+q8ss8dcrQupQT+IJggc9rZ/2f0xwHRZ8d8Y5SkN55cJa+9rjR4c
Ow814mT7jYBhNAexHL6G8Ci4wEjB1A4D4D/E1XjHgFfzqBKd7K0FuftEJjjGafKe
4q319RpABTa5fQ5gvNhjL+vekyFE3MabbYnLaSrTMBgLnCdoaCBj+L9sef+PLm0g
W9whdnfHLd8mb6bVSAqYduL+bQO/9fuDtDj1c+tXMuVAmsAtRjT9G6eWSy6oBjbF
fxrwXSmI4vtUsCy/Z5MSKBSpKGwXrj//t3cjaM9dTTC/zsTuA8AcdCd88XTQB2vQ
tN388571IZEPG6kQviqqY0db25zCgRF/sbSwetHpVEAxg9qCLJSDHJGDpFMSuT1p
8so93NwmEGTwrwdPQIDlO2NDmn9hB23ZfGTcF6R9siaB3Cgj1f87p01uWIkv7HKV
9qaVokT1xKbaCGnneZjFkT4//HZTOSTvmDKWzkioyLOG5g0VNH4sEnoiVb01evME
Rr0RiQmPXLgM+gOYP+VP3pj6ys5GOCVEDGCvMkwnhq6Ws9Qm4Wy1pnkmirnMKOOD
49Z+dzxm5gce6hrJsD81Q1kSQQrMwp01gxZohqqLMax+bybX5lb2R2LoxocZ1bI6
umvtsSCpUYgoGnu46bV4aKdVYEeV3mjsJrMz+HNAs7lY6PBkMOgjIOpaks9H7OAq
FKlgCbJ0gyKL31/Zm6rlkjkYtaMl7Dbhk9ZDXyCkXO7AOQB9B8Arj8lxrBtxGvXD
PRn6DmShE815820sZni9y2XRheUno8phlkX7kOGsfyeP1rZ4Is7Kc/rYmsacn0Rf
758kpmnTPEhDJlh5Cyclnoq63EeRwWL8vFwM7C5zR1caLcM9K7bhzeg9XMfdg6c0
7DqzdUe14oGQM+vOO1MfH9ehxA35NvjPDbVJrRw9h1Kot3Vu/CHZyY2KWKGwLDkl
MOm3bV3iqHGBSaVn6wOgIpg1gceEpH2743/8/2vBY6ZI5kXktmvT50YYGjoIoEij
jtgxJoC7a/iMPXvvuaz1+ICFkgRmxnxCK+6qwl4RbdMROq8HQgZXKs5ASSzkzhyk
54ChjALbtrq3920PMwWmK30KPX3st7xH6NQyjYrpFcW3lhEfzdUNn3qAyziEg6Yu
/uBTqE3KwSXZqm/1KY+ck6dI9ZaCuvL6P+KFS53VtPMq2emuKU8bKhzJC5Pa/ds7
/JqHEQ7z6QykV9KdQPoqdepJtI6tFNgoW5XO9JVgrDrXBa4d+CJYHAJdaCy9swBr
9IE/P1ziPn1pG33mUp4/77x8Q9nxHOXMiX+TXGUZc6K1CTXYV3nO/+i2jJX2YhBZ
2sRYlutqEWuiFDmve+IPGoGCSlTYzfSML1p2XveV7XavZvyX+htyXjf7XCO9hmS+
L3XY2z8vHed1vbaRYCdhtw327QZNMIEpVVsFm0y70dy6d1Hx3oq4aHSpKXbUu5fK
HwhHjBx7iGgiMJwdg/kYV1Mk+RxvjfhNQOx7HBimL48b30AFlnIhlR/oVleLZNCk
4PSr+KBRX2P4jiYqFdldqA0r2lXCFGt0zEu8Q1Cb6SSy/JXzOvKV1P4ceIHWUZxu
5l5vjtmdUSktjTZZXTeUR21uECynZpW9Y9F0Nr/KM8P8DAtg2Kd+xMrHAs4mKby+
/Vwpl4Uw7sF/gdgd04HUWLmkqU3kX6kBxwzEaEsVKbsFw04YURQ1rVQJzhSUndTk
CUdEkVHy3gYshdEJcalVRGaM7/8YJ1sFMHM81xb9aU51vsDkE6++DZk6d3XnPlOj
vmMepKLUNBr1hrlaWOXDIxJ8XTXPEHR3HViqLBZE27N22cARf6cuZj47wOhuWKLE
Atl5auFqkcMee7upntUxxfRrIwaBRvnoLFtI1u4i5rkAcsucs1bvOXG5AxvgyYSL
ZiGmcqgh9W0rszfxaNDUMeCEGFK6kwTczPSt4lqnO3LNsWoLCzNSl5vfsO+2ENa0
wCwOLKDTf26v3PG+/m7E89raZ/R+U0Tc9ihowkkJLzNLR5IPXEUou9cfGLzuhdRM
jdnpxo13fBW/3U8u2r9c0EltE+Ogq2ldE94RoYT7oT+2PKowJAnjDt5fYPNeRS4L
Tc9iyerru6YuJmV96YUAf9pzlEjE/lnGG/dwMcHqeINphUTtQPMq5Z/BCMeAdJ+l
MN//uGjK1JAV6vqh3Vz2CaEuY43MwPkic2yXRwKh2w64YiCZvOBluVT7drA0X5dX
ErNJAOltNv6mla3IjZ9sIxtmXcZxH8AP3j/avEyQHBBJmZum0QG6zf83y0mqc6st
MgliqnaxSJta8upRKpbMtlh9EFHY9Fh/E8GD11yBCkgabw031YRDvIDnnADKtcKy
UXUVTyDmjVNCrx0NzV1KjVHXyajJjvIUQoe7LY5vQT3kiPb1og2FEx/P28RZNyc9
NltMhlF2o0hCoiANP6v2K9dJmErs7RA+H2JGll5v1HXpzLvDMfyW9jYpf5HOLWe0
sGoC9SzCj4uELU+y4YtvtC0RsJy8Ee4wBAUwoTtedtT1dHcd0eLcvzrfl4jM81xH
Zs3TfgMZ3dl9RIknm5c3E8qyKd0qlwPW9XxRoPMIbic7plZaCS7gHfmCF1cawkgi
RaCiGufu1VratDYJffTdzJR6+BFoOKumty4rA9lrOa+RLeWibAG8CfggMzBBvKzV
Me07YVJH3yh99HZwYQfdsNRcPymw3E6g2+SCoLfkOU/L3gizi4ud+sy0pzxkN77b
uqg8m7zOFw7ATRP3ApHesEQcd23AnpPR1bCxBkC9JmVxPUWrDKVO9IrSqxaESuKR
qUoMx/JWb1jTI8lsWfgSlarBtDIC9njl/t3hsdj3VlqG41+NnAGhXEzr6hc+xf8j
Bd9yfu2VeB5mXTPcXXfxLL/VoMq/zus9BIANUAS+3OfHw6ODj71CRmK7ATU1P9H4
/k6h7oFPHg3VBn8U4OO3HvvA7T3jmhruxKOWzUHNx3vReImYNaloLN3ohg/z51L0
tCJx+q2Ub8tvTyHx+S3/iQj3H/TXVOhYkBWRrqgW4ncDiVAZCTQofMB4vSLz7YtX
qzhSMvfzmn1RHhdk6Hq/vh/msa2HfY/fnyArantmyOAWdixC9JITnQXWn6qHNgmE
FCd7fYrONh4C+0JaLA2Inxr/PfwDrMxnRnjFUGvP+53JGNRz1OQYmpD+BLy5Y+Ns
CAhlU0WJ4XN3uNyB6gs6HLBm5kUahRaqccZv/7N1gAKGZqhjBdZuPvc7BkjBMGSy
2HVlpMdpHT8asC52pncvCBmTbg23yWZEBaduf7mDZ1lAHJwTBtde8DcjURP5u4PH
awyAewtVWL7YLv1xw9SH9EeseNK2Tu5jyqZGJTyd1fQpZy9P6TxL3UFibsyr1haQ
1NhaoP0oHbRzbRpyFSjwLrT1fLLcsLeFOsYl1LadkibKODUZ6wHUjMcnt6uRji9K
Fp8TtO919+CEaNhhrtkFonpFogXuc0+CmlgGG3P++AoY3Kuf96w95/MK5193F8Wo
bxr2GvpN3k9hypQ6Ld/0BNFIcMpbt0+wMSbbKqz9rQziWjpOVLNtcIKw+bQgsRcE
3GjVRzRLoMtXrNNpnmVntSWkzl/s5tGcTvx9gEvR4i7GoXpy3+KQCpunfKfK0fN/
0UAlU+tiXvEHIswFSMnULdNrqLwwekPsSRscd8AAGN+k40cuN7zWii3BSKZx8Pr1
e9ie0RA5+tdZ8mOt7barYpYDaBKJv0/fHd2lNCnhT5kFH25dVQSQKPoFaISzl7XE
O7CgYhGSUUohMoqBBZuT+f7HfWCH7SIiV8vwjWW0b9DC4dWiVTRvhGi4m6M1ORJE
Pk6c5X42XPSO3nCBaW+TYjtcw8WcGLjdGfkfwvphb3WUk0WBGTkNDoSYMpweMGK6
b0BX2M9Ewc13hvFb5qK8Lv7rYJU4eGBnmlqem1I7JIa3bSqgEHpSsxaZ9mYVe1Fv
aRUZlf0Jka0mdJHM4CelgFfJi+enc6gq/JuaKYVIIRiZXhxrOF7wVlEdHzaYgNqW
hHGVnWCoP83hhuRZLEnLQB5w8TDIi+2di0wIhP3yqLvg2ZiTH0CO//89ElmJaGVq
14C6qWahjESefktnh60I2eGqHhyfsm/uiBy7aaa5WcQLMjk0s5+lHJXIvWtHyc6f
HHpAKnpWPNXzvxmotjvmhok1F0Z9jR61VE88mdRriVnZ05UnkGg9NYTceTr8DI16
IwOsVmVsx0gGD8WfGvB2Om1PGAjstFvdLzbed55cChynEzs3XTMA7yfhu0EJbuQX
QhFBT7HrFwTn5b9cgH0PCxtjRsmRsafylYPAmclnC5bqk7CUEwTyYOXJ2NRgLIE/
DhrHVLzWAghJegQ4OGtXZWil9UdAjH1ZWhqanbjBh8d6S8CN9Kg6ARvInCmve45S
hhbTOSckyW6k6Pln4IVJ6Vb5ITm+YFG/k5rHgH12lsGTqYWu7aVzFCPgI7AXBZpI
Nw620rzgLHbm/pcIpHM/ofa2fyIV8SQRkF8MlNtvSWlcOC4ApAuyNgviiQQVVfcZ
eUslLd2m8aOBYE1VR+8YfsUmCtjcJU+ifEjkvfAb3qWnrc79YzvsYwo3YqRP8ly6
VdVAl934EOJhZnOd/xFrli/KNic69bLVl3aFEAtRn03rovw4zkPw/+jRr4R9LhC4
FdrcJTIJAW876ES3fDiEDC31zccK7bhA3/dNu5/wMAb7bMAx8JwjL/HveQbE7BYa
QrkDWchXHSOOo/ylJ8pPudkuu3B8YLOpKXi6bhUN7K2Uyy21grB/ZYnYfDyzW4tK
tKdW9YLUFR4Zw0HrrUlCVPyVPCcSlfTd0AKu1UN8gK/WlvTh2MOSIuT8PRbL4pYp
Axu0t/NMlIhXYDVoWj4ff36BxMSeAVYb+gVAmNwtSk0pyBLahMqYr9URtcfhK4lP
YArSd+ZemE8ExE+96DwOLIaQdm6sQlivImLTKha7SefySJnfqcrC0Lh5fbFtqr+2
aceDFL7QJM33JtcRID4Lmyfl9/eCBA9oXJLj8l7Rgfkep3kd5W65vV0yBtaV2vyZ
3a8caramakGjXWfEKjFTnLxEO+ZMQ+06OQ+haBLOlo0SkUfgzLroCKcH5f2YxzKE
dshDslnz752k6coyJq76zq7wwTHlbp713+szRLGjoItHpboQvjfwzAJkkKF2PNEG
y/lt3htN9uGA84EOnpuEfMLWZuWbF8qanvLjTAbxBlevMtsK3AvP/2jgLX0jzxVG
OXf9Vb6eQZbOfUM+RTFMIhaE2QWk6wMJsifOvTh6Tz3sSXGQYCC6Esy+ZzGouzsn
mFGxGFOrap2HhXdsqAgCmq+iyMsZ+qr7tleI4WUJ1o6Xv03x6tyoMxe5/8tjA9Wu
/K8dR4cVoa6grAKEW3tiNADyfGCUrBwCLVu58QlkEgeVsLpORI7aLKAPYUug62hE
sbiBpxckRPufMUz7dIoWGjuiE6pX8FjIoZ9u6ZTxpc6SlmthCOn903qKCL7TLJzk
WzT3C8deM1L/m96RdrHEMjCB/V5cgwwJrhksf/Ga3YyTqN/R323CiZHLowKjeqVk
NRaeDf8ke1Fm0BFPU1sg4P4f75aoSJWY33wo7kJu+2fLssH8KMhNOtY7YSa3Y4Dn
ZOKt47ZkAa/xaHWiZm2hZ8YweXxnFiuJylWbj1rS9LlFUfSfxESQTWwXDiqg9bEp
9SPCcioU8gFlKSysol4ES2xEZHNYRqcQCAYKSQVTtlI+Veo2MT8GEyyprvzjj9H3
/LYvbamVT4IcUpMdhPTJA456PjNwa8qbsgZgiFHrA/yUHdZPZxQg9DbqtJWRiWWR
qmqgo45o+IU1hPhbCEHdHHUfp0FdTnxCxxaGonUx2NnPzy7nrhzsulZgvgxa07V8
FKvnsjfMYCnyJHRISVhuvxr09QyGiUt0JQHZwRaxo33MwioQDfn5ZMMlK9dw6dx0
6KByczFhvCdQXt+FTwLhQT9aLJmVb58vpGhjh5QjKjm9Ty56jnIgoYXLnCNNv8av
GZr1gGapHvulKDQpj9QpuZjJxnT4N0wOMkaf7vTY9uMgCUANbbdwSX1MuRPTnqE3
3pXrnDwfkpFYXCIK6ofUhdXs5A7TchdLYV9ZNeuffrS47FjbBVyfGXeASPBPuHYu
H0dO5Cv+91yl+WadAYN5YT6zDxsJgP21NzRbRynXOb9oGeP6U/f1b0ZxWgM2YLFB
Ctok1Q3nr9N00BoiKqTI6FDbZWaVWH2zsQHUvLdQXpn7smtvQxkqt7qO0SMUSXy6
Ix29/heo/3wT/srJtxRvJCHrXEfsYaPF8lyuMwWeYlD0EoNlRO0XSadEEh8m9rqZ
ybmGl+9SXjSIqfkYuRjFJnBq+5xIP/BrD/ErhTW3c8/PDHARv/LGjzoa6We62SxP
hw9iP+UlLubkPISpRS8uY0HqAqexdKXLCYQt+aVosXq1X+1RT7h7/+Ttg79wvaIS
7y1K1W4/Qkn9JzU0xpgutBcl5jIvS+N+qXLJUb9iw3j4kVF9Sl6+rIOEv4AnxJRd
jX69lkB7YUlkgAqk0U5ljZIrfUjAgcvGozbNYVy2MZCkZ7sNN7o1gMZc1btfHMHf
sv7TeSmP2p9CCODYD058bteEJmtct+ehl0maelvFnRbHmBTicAmaTATFMpG/Ybcp
/m84X+K+kkV3HFUfpu+ygHsal8coMVMDQP8V58LH5W0Eakm13Ri81+fxHv4mPrjN
erU+j8Td9d6ZNpUiZjqS8CRbezbzbyGO16jh2wpDtukibn00t2Gg4KYuvvem41qW
B6RrJ3Vye6JTw9+JhzKxnB/wzPdMdIGfgu/uNYe3Dr47FaeCh56SW/BrVBIjiZSp
i9wU/ZaTKw0LgUTvna4Ib5j9UgtppSUy5/25K++0bnLdpO+M80A7BpP2rtLMU0Ma
2CRP/CPec/ZpELNppcL9JIy1oSMb+P1rKzMtCoMW2aj1nOEPomwBOKZiuxRWMPet
93/phUKXxwtJPBWdd1IdyCPbNL4Xab2k7KaI8DiAZtITt2MzvM6faLQ/CRH8uCPC
kO8+W08BGF04ObGrq/+91HutDuxMCvbO7VoeGt2MMW8VuQEtcD8gojHYkMlx7jAj
VrkobIQi359C4wkuXO/Sz/C49D65L/G2IRQykWL6/pOG7QL+lDfMnNrgAvW08oM4
XJguYfc0yHWK/msNnTH6bItYj1fpbJKQdHFu2Xmz/d2ab/8XkBm+Zn6+PGUpot9H
1hP/8MM9C7cKL0tGJpGLx9NOYgxYQ8HCsaeuRAsq0FvHkB9OIRHyag9zP8eav1p7
ygIsx6eM1Yo6LsOyl09lZQuh4c0PpZykntvYLKhLWxe7QEInOrEzRLbB7W746pt4
5T2rFYqyzN3f46Loqd+eTBt+1sNSMEQpEdYQ/nfbFHhDMCI7X9gxIN0IPDFnFlqJ
ynr6argp/U8mzeJUuh91qx1CDtZHyZf3GjeUqCIzvy/pN6U8S3CdQ9QBHGZSEvMU
ix8RgZxARybwrteHweqEBANHUaKUtCRccFXFQv/NJkiq8PJj6GN+sX6KJ2Cuo0tS
iI+WhE8lukTveIuMUvLIVZEqUKFzns0ch8UDJZL/AJA0XAmWIfgvKYk5asA4bCBw
mpLcvIdP2TuY2YxoFJ8PAUW9f0NCh00ZjpAPtj0mcFX0NRO0A1qM0UXpKUU0twFB
Z2v9ZpAJi6Obe6kwIsjBs0COjiIVfVguPlatcNb4RXBLVmKBNTCaKPDz4Z5McvUZ
41Ji2kaAz2nFaIGSFvOJoLf4KC6QoAmKdLP8n7iYpr9C8JwY+ZkK3YcxwQd9/DaI
WIr/H6vB9eUGvwNozwWeB+dUuHSZZvIYiY/4R4k9cdjaXr1u6SduLUkjIsFRgvPq
YJt27bHljQHGHCOggVu7S5qoEq9cKpaGiFyVoBv7khIPGtCBe81nGxkVNEDrJnnr
lc5WG8QkDm19WeyqyJgUXISskQeowzD+3igEs7p9CQFmSn0qvSvaFiMSg/P4qN6b
eN60HXjjr6EtRaDhNhTa0nXtON0Z6lwkoqBM8coqH+NPKn2TMyjumjbZoHxQ/rOd
add3qb7AfWz8VH3UhQ/seUHj+NI5EX//jl1i73kBDKjm3zU9vNEAlJTnN/DEpKpf
5yhoh9PkfCFvNzjnZE+VDqrhnfhgqaSz3/qQvR43jnDKr1j5jKvdeIs78S8XSbi5
vfptRiplFnQ7iT2RGajEkuLyjStRynuKnBvMfweepbG3XYz603A91cPUz2tbHg0x
2wmoo1FCPlLJ1BaG0BesNGX8yibl8JMrKUwQ6sw0hA3jeUlp9//BFaFFN0uE+qJ0
AfpKiW+cQwPwMyCFHAo50kVnndFENIDVmHWR5hCOp3/Lqs28RAuQMj0bOy6Qikuw
Vj9TY0AcOBgAuMbXFCz79jvQBz47lC72PsBbv5aoYh3sKrZX0PtVBptFVQ1j0Jj/
GgotBiR85LCNjzNNSrYdQs6zHGiWJS/953BhEHNkdFwQTEG3OqPa07E3X+xgp/6K
56gg+GDzOguVEllnXCLJfgbUPjWHmYw7PvYzksIcW7p78OSBWZH0AJ+95DWbSuV+
mMyMuOKBHi5pR0rLJKOtKW4ZnU68fMzV6cWEWXs7tciOvpVuJH/6tnz/Y7JtKe4C
4DlFhM35ydYfjNmaYk7oW9XQiXymgcXEnv7sFtNqlg2yFvD/W/2We530+lGp+AL6
LWXLqKU1XIrsyjM3UKICbTu9g42v7cVdbgD4uWFcfbID6r2ZcdUOGBRPq4JkVIwu
kLE7+cbAYuU2NjOrW7dv7AKpkr/2gzlYGGdnnw31dvCgb461VVCOOirKvxziQxN0
wJplEkxU21hQV44Qg+lwye0/tj4GUCDiDlpbxhXMaP/eO1qVHg2j904+0jGOU7Ps
YK5FWoDXO57CqMjgkx9PE34+g55lxrv3K57slmWTX5xojvyDlqe90xJCUdCHp6F2
K/4TWpurth9tl4tQ++XXBKoXXbTHcF8t4NPhb+807XpJXge53ayJm3zSN0cfb/6j
I5Kr36+Asn0GmZ3exe3HLmzVhPwvl2Ehyt7JyDwdIONpJpeClfYi+WgbcyHqiIpX
L+W/Q7G/pJDBKfYLJ4wqfUE3DFgFCUdRUEX5Ek365l6ScAx5ForBdJi3/vfrxFyO
LYx1T7Od+wESaBVPLSk594tRjrcAKBLalZf+BSH6x3F3E4rogCZlPzV2rMNFvIwJ
reCRjtIBf05eVIden/lHrRrNkTEbHGasS1deyN9Ae4tU2s7VBnntE33ex0EppwB6
t5mZHP0Q51sNMc1ryfaexA9Wn5xjgU8CJ6GN/Tn1vgYzCPdyo/N1gPvBxMQ+xT6Z
0FJEBz05nPKF9lEey4NrCRHgD4hAfz4e8InujQpTlVJnFXZ0cFHubS6ztdDpiYXO
vFPdT9zFzySimpskwpm+/HcXMkoptp3kcNiwDl25JbiCBEdDoJ824Er3mD5edyCB
ilQrwcC7wStosdxZX+mhmLHE00T0lLqc6xknGfuMA7ef70es1cihRLfNUXS73fY9
TcwzGfQDsPX+OrKkaII4qZX1lMr7RCNexLlmISken0DIfx1S/G5ZRRd/hfwUmWSv
mbZrspU0FLgfm4lgpF+a6NdkvyiW0vNlEYWVFrmVQPHzXlM9aAvOOTxsZqRTRlyB
ImVFRGw9v9ksLGl5fDfZIvvZ6hKq/7ZxdhCxPCSbpfavQDoqd2seBuZcqJqHVT19
68DGSXgR/S6ChL+Tn2nPQcTlKFqlABsEvySDFY4zxkZ3YDmaPRM9w/EohczELkiD
1FOeA5tG7Y391MhQvuVVI5vgfD3OD5hLEcY0swo4mU42m2uB1UL9BaoJWf9lSTle
j31l0UkrQD6te8XZMlWe84ctHIjniuyI+YCIFsFzPFQQHn8xDcAW1fY1M+rZgc+z
APgHhUaB5s+mtBIHJT2MRS7bVei35becjuNzPJiSWDJu3rzfyzR+4qIv8vdfnvNP
MnS+cHGaw1unRwIirhFwdEaBtxQnw/tD2zqSSKqUFJA/M3YuWJLTTJq7sbG7FuIC
XnIpp6RyMYJksMnXkx62U/QcrZ0IUjk0Q0TgNDkyoEBSm4Orn5pJx2/TjIg21J7s
kZyXYhRfZVHircuHGALfqe1A7lRgqMrF+B/bjp+OE3NypdnTZbPZGGKErUg7tW0f
qhgnue0OYNCZ50pigIUBfq6lpEDxVN80zs0IYaU1gua/QqI7AM06g6VMQUoGD9s4
ibY677iUXcY6mXo2BUNzdUycITzX7cwo5VxZWkmMUNIaGCitCwrm34Y8JqoRXgiu
dYVG735TA/0wB8MxVV1meuIjcPD/xXiYPP46qjg/On4MZhMTrF4BZcr1ZcdGAKDF
xol8FmsB+qEC6FaCndzSPRJ0aBPxUIqAARJs3v6qLtN45WDOetFeD3T+xo+w675T
MG1zzEz9Lf8lbzk3hqjnfxPEXn38hAJxeBP4FTvNpxKk3x/Z+g3seqmuxxUCRedu
LlDrjLtozwdhXyej63Nc6tFnLFmV6nHjp03VV96rrVHZ1ByW8QemJqZY2nnoFqfO
bQkLcrV9fHQQggGXBHqPIewuly3hZk+0fRmw1Tf7tEaepB8rGB4/izm0BRymzs7D
3UnhJXrO+ReIPTxFn7lvct1/FCAi2j+Pad+rtcbb2PfwkCb/ZFALc1CQA/9gol6j
DRO0MWwI2irjRgWxYPmJfiFDjYALJUtBokqgiIYmG6f46iBrvH7GiZl05LfjiRC5
shHnj/4KrRo1462Cpmce2buuYAcOP8ev15sayGuLxDGvyu1HTPyV+A4lowz2b6gf
adFuYrild7ENAA9HI7EwuzphlEXSQZJ4QY6PNIn2iTpnB+M4eIGFkypvBD6JFPz0
x+j5e56sczuQnY+fsnAqrh92bR+/Xi21VXarSwm4AaJobmP6b+1HO5OCJ23NKwt9
llB5oU17zVHcKrGRXzeU98EqeadHiGcgqoenutUxKBKe1LQvZmWbiZF04r9ogmLt
6vj8aw2jN6ChoZ49WMmOtjB2QDh90NOAiO7JgQ3i6IJ8HPpfZmQ0th7vsaSjbkKu
jjf3/Z8djlMRQFkrRySyX4Cf8EigiTgdvJbmg+dlnogL3XcFHYu9YbYokg0DCOjk
WBosxnhpAoMEeqCZZY79bcCxFSb9obw8ladpAiYICiw/953WznQHLHkgZshJmKZX
bB6LX2SvlB+WfRQNS3VHhtZbcrloTeqk7ZWGKXAUO4kuGFaR7e8TndGDHhtdip6Y
L0EqTGhrhzMZydTfdbPAL/iO2SknvhcZKI79e00v5XY2ZBmNtK0sFtF2hyUkWTUh
UT8qrt7pJOYCxN17ovZTYABl+WCR4QCJViPBk4VMARr+YNsNtoh7vgrAIvP5yUN0
mF9V58fM8X6V8WmhfwRdrR4u6iE7SUQtqpF3082TO2ZmjmGiujOWMLT0m+YNLchn
lTdVz29HWybVD7P7yEmGoxLCpwdRGljxFdRXwS7oek5JClt4YgXVjLjPmyAb5SRJ
4IztP50bcFf89IoFNlwQ5kLbB4eDam3twrWd0pgRHxMZr705qo9NS7CzkI0nrNYx
sdfqj55NGWqu1a+YigfKVd4lpQoiV9JYIXMWvGmXRBO5HuWL5+MCHE3gJtjGbYJI
RG4NixHEQwPd3wFSHbinbHRzP+kdWCEbprMyx0AWMfn9ehE+SrjFsvIymlMEF8Ci
dmD7oyjznwVP4ECopLFkN0yDIgu94/IyE0ulz9bG8XG+nJ0WF97cgsPg5VXbg5Yd
fOm8v94fO7Vb/FSgNyh7d37sUqi6+fssWBtEYZbDuzp7Fz3/QbN8uXMApd0baGrT
yp8j6DuyARx/tUnNm+tRJ45+iduFole0pOoOzC531lC4YRmgPj/JG56kwdYv66L4
AIxlAbXN6bJylcxSE9jJ6q469h0QF8jtbPSgfMd/9+eW5+BrPH3XozCai5NPdzEI
c52yP1PHsn8Dj3YRMhmaDAWn+mHv2+S6eWV8Cy1yIbGxUYCzil5yNeuv01zZRRvb
cir7DSpsjX72vx2YMqjOjjKnXPSD3OvHv5pCxqhdfyfFeTaeXItPWXJ0qTntRdsb
iMJE2uexM7nv5unFzlWgNEl/EGBDgXnB7ns8JlS9eGjdEWryADsuDXfeM2yd1J1V
MCcU6+PhlNpd00YaZ5NuwI2qwkIb0I/z7Neuu3FduHouaMaLKSYJiZ4VSUSJyryK
NS4usm7b9z78dj7vk29PoeIP6QToX83T2Fvg+4Nlhyj1ZAhyqvPsQw7wjclINzYX
2Z5IJlJL/rq5jAzokHI05fhT+aaMQqC6f0ZqMTd6muomRIFIk9lx+6wymgjo8Lq3
WWmAAh1vXP1yvRDnwKK2rqLngxA+lt6ghxnS8XsHqzR8NeOm6OfRxsi/VF0z2HG8
gB9MVDhcktwr1CsXCwiiVS1ljWt0aiy39Mfijx+uzrEtI9Iw/lZ2d3WOxOM9/rGy
ehdsRifO85IetyuW7ukzYuYsdf6EkzsT0+TViSYYynjC5tIuLUr+KNrqKebFn68d
7BiXqZ65y2S62IMkfbLyE4ezF1uaBEMcAT7qrxQUbl6dmqSlsEbEKx3owrVfzbE3
vloLGfMmwvhumpb+fJyMtwzaasViQgn5h5cqCd8p372fWX2nBZwRelNQ5QLMA6Vn
EX4hcaI62MwH9EVOATWJ9v6BTXb5QryHsCBc982J/KnBwiMSSLFO8/FjEM1dnFRN
GR4pPQadXPCVBm8Jn7Q2Qr7Q9E+6plHyCSx2MBI8AFBMQ0H5lJO8J0klCqYVSBzm
GDdMxvvddJUE0cX6YJEorH7OFxhk6zfBrPvrR5x/O4yesSHyZ7Aqu3X6fCFEyoqw
wzOPy6OW5SNcxR30cfl6qcmWMQ6d5vW/oPFE83b2EU8mY7HTjx+xxAz/03PJgbIa
vTkLPWt9Z4hSI4R9iV6KT1plEqVHQH1LBXtzilxGjHwzoRRyLuyzrNZnvBoDJbwa
TkbCExR1HaNJo/Kck1frfY2qFdxjVlLsIipFD9N0vbWDHy+xqbP4y8OYaG+caxNN
oT2gQtfw40Fuud+ROm3g0ZytJkCmzsNbJrVCiiOMA6qbqSTyvqu+fzRaNcuQFcdj
FAxz+4dW8PaJbxcSfpyMNsTEhFAl8aLTu/hkoMi8e7hC8JOTT03WILVMBk8dhiHP
owsqY7sa7eSyIJwELePkjxq8G6/FfFTl7UmRKj17ughTQr2qsJnycadHyZwbd43v
EDGPkAyQaJGezQSBi6M9i2y4EdH1PIM5qX3O19B/aSuUFqczC/IXIni/XeVDn2Ty
NI9ry8ehRF1Lxq+jDJIzX+kjMf94I0Wfb1V8b7UbdpK0Uy0lIuGonolsSCXt2c1g
CNhdCFzZMA7iSZZN7JjvaWetW6DW5wiPOH9r+nvg5zhF1v6MCEJ10Jm3AIIjLbi4
x10oVHzyMLvfd9T+1LANGBqccJRYuPmsFIDaMkDrSjqER1QuXONZPsRudyd4FKcI
0zvTvMk20Yo3qMQ/84Z8HertBY7GlOCQ199eGt8ael1pcqhQh82x1Qy2PoBy+3Wn
/UgM+AXvs9iKF0tIGBaDMseDTQcpv2lkapkZYdOtGub5CmncSlBoSoLR/LigwvI2
h6EOm3hdVM9xX381Mg6ayPajuujfQt4xFxHmnE4hmLqUVRnWygpf2zH2GwOxBGIy
N0G3fICEyhej/DR7n7IYOZItsr2CuTBEiWlQGzfNmnxz6u0EOlMmuTzzTKL5YZET
eBfKfIkoFEVtiAi7I3spZQlOM3qrfbzVrX2ji2cnQLOujbbs+VrqfkxlZA9UWRlQ
61dTCXtBaKSZduLLpT8QPHXBtbdVuSOtkKAaOutEsVNCdBmODS38zNhWWJAyEkAI
BCkYG/WrfxAq00ltYpdJvsqmbLXENg6pkEp+j1lBVhUk6rgyrHg+n35VcXZ0gp2Q
xoJ3U/OfFbCWlacDkKdDvwsjoj1D2IbxvLhACmIFMuL7o3kpEmijdjKSIrR5LBrA
sKqf/pvAn4DhSHh2ZwP760cSwjAHo/lADsQQ21Bw4VG0V2ccULqj3gx1of6O31Oc
nY8+SKgnlXLGqTV5X2oVss6Qgvplmjm20lWC6CH1NNa0g8qWBo2E9jH3c+svJUBX
IXTsS75SLP+miHL3ajeq+CpIok7P3zdbhBcaQFRthWRkS/rGcofjCmoYTo/Mg58N
IOxphabVzkComCrXAQddxQgVgQiUUnHBlzyb5yLbkrqzJhfdyt9QU0Oi9xTD6Tta
+BPzGqFDBrp4ejCLnPONcM8NyKwfE7cJDK9yq8rDe/Sy1xeLmtGScSCOIWGnRXz2
KUnc6G5czrCm91oojhCqG53HM0beWYV8x/xGGepy93vsEaMb95UQdrdLdTO+bfgL
Yu9GZ+vEbyqfxkK1MoRP+McAHoAvt2XhU/Eg+MMb5Jf0LrtlutC27mhtDYieufMt
DnZuyWCKGgO+qS1QJsWcbSXP5ynFerJxkDR/oWxnpMM6EWOIsHm1wctm+dB3J3WY
iJ3kZAWjYtf5MtzHM9kTVj/ocG5BCiQwuPgvzW/Jt7tbqz6ZYit5eY5HLi/d6/oh
ALKZo6tTSfD4e6MKKTiRN3zSJaVJnoFqfX0HCgoElXpvk1CUBzaVl4o5DMRRULxu
GQNYdXzORQwpxrBIvp4+PcUl1+liu5gfvqJyGxaKOLzmQFtPQe4JI6gfOWOecMgt
siBSEbyIKxGA/1u7asUvBzGAsSvrn8TimC1bfeuWxBjiP8VNFXzkWgYLrkE0FJai
Qzyn8TFgNG7JPgtr5XkRhTqBqtD9vE/cPTi+oRXqy3eNmG8cXc9pKMych3VirUmm
CkuZi7NToLd3Y/0FZyeXMDlifJYDGx8MPA+KBf7Er5n01C3XgYnnsM+mNegVB2QF
CIeAp5ORAv+neLSDEbnH5FL3Zh0z1I4uKZkfbPxIU2HLgRAPhZ5szfNlAltvxOvv
ZHDNmkaRgD2QbYsfNxwI++JDwK5DPlWlsCMYEKv5hibVYtNQzet3nk+WWeR/kZB2
QOOJ15WTnedkqNQ9K8GlZ11IilxziDdzPlj3sKwl3VU679n5006ArCnFy31NnTW7
xTuckWyUo/hpw7fC8KMU324L3ssQ86gPT1xr0DfcOh2YUjFpVJDBdumXd7cqw7Zq
4xyoBul9/t1FulTpNdrZzUcxJT39bkiDnnJJjMThDxnPiqqSZU697Sb0jCTDqGdN
RQ7v9cMiJ+0yyX+O3qOSqMwxjcMw3AvC5rq1HPlxE+vMUTXDje9ea6Jjhmko/Gpn
havDR4wujhq423gKYsVT94yJGeM6cpB/oJ7QpOl9v1zKgKGBrleGrDL8rOZyfxK3
pAHsKTVMak5MfRdLrUScK5bdkdeTT/9IfWpMNSAW7hz01LShUJ4dk0ZnzTe4Hcy/
t8i+Np8s0Sl0EzySBycm+DpZBSOAFSvzY7d7woon9qOZYK4H2HwLkuaBpu1ee+JG
9gYbX0qTz/JXapEOOeWf2dvS27kbC3706gWyLbsVPtwmbVWp/YXt8glpvhhIqNFV
B1Yc6j6rw6FfG0EJafH+NXpUA4fGNm7YBXjUfZzTqpkXTYz9th7fR+hccso85rQ/
huHWNE1jwiFewqiOBUEnXNu/enrB9TzXlcL3v0RRPYizJE1ZucsuVBJFo9CvVHMb
IIAZ8gQK6pRM6cv0gwFuVxpkF138ZV39ruom7GSnfa/msMxEUZtcZrl2Urjs6XD1
0Q50uu1FuspmehqJrY9jWnDciUCII2UkYhnbdhgqMU1qBabjy89Bsza/fxEoArxB
7inA2orfx78bliK9dfLjvpk74V50/0B6bzDV/9bf2QIj2mlpW6Gm0N78UYzmUkYu
e5JgV9sL8zDzjiHnOMr7oV3I+eF4Ec7JjKjJPfnZjIeJK8qBTxCebEb7cYRxlLMk
MPlydR9K0NlYwn5Jqf6KkFBmVa1hDfkpwE8Dn7va1Ck+XP84Kc1K8ZrTdggijf/G
u6OzIbnB5HlLAY51M7Qg/iesSUlomLHD3s8tAu51tj0jcxYnW0qLztQyTRtBiXXJ
8pAMUcMtXJ9u1YAfotue2H32rkaAc0gv/pkjz0daWry4Jku9hfJu06ICrTeE6FKF
dpFasks04/dCgv+2IWw+Khpbj3CpIa/Qi1FRuOxesnG6iMCxod4fxMFJkDSWi3dF
AuYa8Zh99wAsy+YnkuqQ1mCEXtdkAs08/Tmf6+7PE3ct6usD0FezLQU7uj8s0l07
XOS+tYEHmBHwdh4idLM+tOJfQE1cvN7SM15NBavdtTSf6JhM6/9ogv+aVNOjH7r8
gxUOCqYwo49PHTXvOmtX5uavgPLDRWDjnrvh0R6mjbOp5LgXu8mkT0kGdZ+5wZut
aHF1xoL9Dcwn4iqm4X1nCMwFwJkFCuvDIH7vVSbdZ/FmJpWnyeC5wHHMXaK1pM7d
I3xWj/rNB9xubwbKnJs8dnydmOI2jk39UyoemtIj45QXg+4KBk/dauTk6pwp3DCI
0UF5gS6PE+EWEy9ViBE3VPxHvtKUdpJy5Uzpf0UgM45N8RVblcBOwcJN1ug4H6i/
i2I8qqbCAw+7WtvenCz5kyvbn0NuMq3dw3QgMgUEG9rTr93Ic/O2Agj3cLHG6u09
Ilcgb9gVXmcNxVnu0HcjO3bdMCTAgQK3wRwr2vs/8dGSm36zfpkqAlAxZvREkWg2
EwbK1+X1gpcn1nGOaxym9wZ3AinRuUg/QsGN4zCdHBqzozvfKLgzJaBDIToZNyVl
/IH22ojkrP6lWiOb3tKCzdl7zEPB4udw529uy/vXC/ngum1X6HsqHIIp8hs2P/Lr
mcVhnR9DT69SnvVN2vbCu4m43XJ/apF2GKJRNlO3ubx9dU3Qw3ZBJSNJnus7umXB
IHuZamzMQWJkmRnI/E9JDAiTWh1jXrwts8qmYwmWXj//BhFVbKim5Y6rCiliYrWo
zad34nS6o54J1jS/G8UrJfel963t0Vqtdq+IovCdx5N0Jtosfii3W0uhIKuPIuEg
tXsm/8sc+zA1SMxiCvwYLgl3J4fm1DP05pWrSxrfhmO7b3KgWRZGo/EImDXDs0Vq
EQiYf2cPenoCtqt5ow0pvgk15NFaxRlTMNJw6iY1xg3LrCKKL5um8pucDBs0rlaS
Q1/YphnZyIUoef9sAh/5+MlBdCcuY1uZdJhczXddVa5VijeqNMeWX5Yj1h+p6W8j
RWzOWV198rleFxPbTUgj7DCI/TguRqxmxezTPh0M/cNNFc0ZssA7neyOk2ZgBehv
RTG21JbuMQBAdnMnHwpG2iPxS9ZzA93Ln1kPAc9VQuqwUUqEjDDI8iN+0cWTGIqc
IZ3w9gC5CWDugPLOVDiIdXj13H6dKhHEfPgITZlFqYQmyQ98Mgs0F/w8TR4Xi6Tf
L7APz/WlTzvj8e2B6j0/NtmXduo92DGRNhiUfd4DIwxDk5TaLm7FD9lf1AJPwph9
LILMMIPaE3Q4pVQKR4jqwBsUZUtwBivKb6LBhor+UveEkZdoqpHoc/Gx15f1bgc1
2rE5uWZ2krZvaBn8FhUG3QIi11zhQzGAyKfhvIb+TjqwM0yvts72TBbTiWxJx3U2
Y8cb8QFo24Pt4xE+0lSgfM8a2uLr9pjvOYLLzZ4Fwk+tY02grjKPiXho9Evz8uPs
kfdD8bOqUcZtTuyFCvXglrgoTCZPq1MfswXIjafx7v9m59owsrowxFKv7iv2pD0Y
8gkZk6oQoCcqa5CfnUNkq6T4ciAMB/joaFTXMfAqPfUqneYm9NPzX5yjQ9RPcyaW
IxSaOkgvBQMiDcHOE8y/ADR+LkyznabUrOoJAzQ43bRB62WKfviPt0ISVRySyesj
2Pu2amW5J6IRDpz8pYOpuCjnaMnuwu2NA92laqj7hYsILmSxMBKXVImdMgoIg+n/
SgLOMjBtOfUEPjfiblm94nYeexv2GfsF/Z9BYXUl4B6djU3LTPBGDmE4X9sTY9yM
vFMxzkwskm0wa/1SUPAbYfMCEIWt4QVgnFUzwlkdcNijdsgFdxC+XcUgJdQphKSr
YErR3RCT/sfSpSsitwT5ZahBIuGOfktaPih1usIoMFRheEph0moeYFlk/TIxNYme
6iAmmVqvDFlkNBtwcz1YQb0QQLYH8Xfcb321kBbYCDkzzv4WMEt7A5pmdT5vVdhV
4hAOnIbuo94uZ1kA8cWvEV1fcCjkoxebtgDE2xr3uzd/Io/BwpCjlle+aerl4ivj
uqpnDVIiXuYBLVD1SSvsX8ONN/YVm8X7vlV8xDYCS5QCTDAIJsmH3P4Sx6yWYh1A
paRcAL7taKmPhxO1CnQYW6BUo5ts6ntJcKhCv+/eSf96HptldTPScNMe2GOVK7Hv
rLKGnkRz25yIt57+fjtiBriQ5YTw/YRoDK1cHsP0nYPG5QC/cVNbVLZoi+HKQGAn
ZJihGABy1SN7OtX7CXoIudIff5tYm1x3cXtb1VIfdbSSDRtb/FilEdMbrTsf08Br
DGqjDVaw3l/m/4PvF/SGFvFNUrOYDWJYTi6Bgu3yAAfbv5cD3GgjM8yUVTdl8lW5
Ml1Qn48hnQxnZYPuvEK1f/W3Mw+xJlTUBFsztmwO5feqCPDqYzsIWHOJnUgOgNdg
dWW9NWbW5yn9e3Pz1WlgfT/usrugHCCWzz07yTTkrt25m3F69cxobWqrX7B0l4+h
86H+sqUS+6Rn/F+4PznsoBqbC2CqaiA0iJX59UcXFQISP3L/v8tpS0z7hmGC25zS
1wL9HWvCfVirVGvgxm/HW+88x6tkI2mPVB+ARuvDit+YyUbmiO7OZomHotOgea2T
UrUX+s9B6hTjbCfW7a5LvZE75BOZHlG2ORAdRDJA2IwvgeVyjBTw9KueRDLjcXXy
SN7YAj31qJAyAJLz+Mq6wDzgw2CrScLz1nRqgucTnK7JJlBJXDjWo6A3P2zdfKqp
v8UKfwCzrhmRp3UcXDItnRtLMYR2WLgHJqpnFn7JxxBgYFXTfKTmJFfc55r+GRlQ
OzVvA8AedrpYMDLf3KsLgv127sQ0ew2XJ9kjfi6EsrK6FWl5PAjJw2n0YrGOthdX
iASINd0eC7qfGibYUl7s1v37FfCRBJ5QwFuvPc8gJZ2GiWPvJcXUgxnMx24D0JrV
9+i4VKqqtqcTKn8hGGTX0zY0LEW+u77cyfY0LmBVf6gycnIjxit/nN5oT+TRQz/X
mEL5oq/dCg6+QOMMFvGovs6G1nO19CL0p/FFVWXIKzgoGJP90Zgm8L3eObFz3PJE
UFCNR7Aczj8PzA/NtkuBDJ2SJB6qqzjlTeC1onsuZ6ygKZHBlJubbl5LEX2dm2r/
KYmP6tqxQTOJp2TERlKP5sUdRCu9LBmbdLgwa8lDBzw2qZkHtfczUYDep1YOwyuv
elUo5KnIULi1AgApJpd2eJ36xg5aW15P58tzDNPthos8YYpGVIGJVc1ZncRI3ZD9
CG/tRi8AcrdMDmyxukmnwyAkz7vf33JmaECVGS/nXAiKLxza/sUlZnF/LkStQKBc
mAE7ZoQ+4u1ZOFsW6g5w5dVcf52B/j1UvWOX8Fy+pyD3BD7iuXt/aBlPg/ZyL807
YoJMVtsdWMwrQz6tPBXbMmjSOazf6lw/XBsmjeIzFclc8YIJJlJKeAWk7v7daYdW
oFjZ8QvQxcHht00YAmx7WIQYOrT/FwU9UVuKHaeetUFhC4SIB4soLgQRmX1DFixF
akKw8pZV8RfsLrDgMpoiPKBmk4THvDP4jve3UrmGn1K+gykywavBfv+14wMgWSU9
2se9WXLerlDMCdvbAQdDuTTSXdhTXTiXgR5xtdKT23ctznGqVxH7lo5lyM4DHnuL
tVtrmDkXUn70xEK4zFZzwmF9b1z/55PLQroBSJv34vJ42bk+N0rAzjoDUDBGdoxw
Vq9vpNxhdB//9L2KDwcLQnaiUkPozC/Tc74VJnSbaGjyGVHHb4+OFUQlA+ZM19ww
0d/u0yAwXhHt+52+30cnHzyCh0M7PDY9j3VV//T0GEh9oW3vI+WFKznUro66nTj1
EsV7fggCdy1lSFvRn81gBGvx9goZG8A/TjjowhTDAfp6dkZSKJSmgGRhyCfCTHhH
H6X6fuWdq7o7Jlr9tQlkx2IzDhiXSfv3xbTAG5p+05ZAbasOabPGFgdJWrbR4hCO
LrusK/1zQKuGecX9b1/MaNfXSgy9ILjnyNAZt3X18f1sQCPCNr3OGHdMb5JkaBso
F4zPO9RoZZmEsxaC26CsjosS/vDRZtwY/GsoxYr5ugJzw8wpLmpr3pEFTz5R7nnC
L43yuXru7BKdl6BAXOFVuT+M/71omVIeEUvqFMvdhxHYg4DFM17wtolJzFryUOYo
9X4x2H3whBwyOlecg8MoXRxNFUlhhdCXiBVC+LfVQieeU5VN0IEe/eDiprtVvGdy
6A0u/iwGxuY5xC7GFwn1O67qTJYojDs7iel+2NfPpo8kXwG4guZNoCZTZFjUHTmf
JDV+JI61v+oruPeCOnV/PVfvAi1e8CH92XjLHHVi3Up3y28tJVwSi4t9HLZHeZNp
Mg9WHP9x2gobjR7ERuwwePiC6ifcQf1D9ejDo8QzS36UoSoWbhF78DxkwKHC7UYq
fn8pFKXX0WAnuNu0+f36Hso+xsqRGILxvL7LojjB8QGPMotbNEIHSNSvxRzyxQg0
mjbABDEq4TLUDM54twHEeF8v1cj4pKzlSpUFimt2XBnWWy/OgCGJurStpKznsYV4
itfiHbYGZgttYLXGLKsomoApRJPFGjglzGZP2aLqZDH668UTDbd/T9uiteKBEXC+
WatN8ggvWsOk4/2GH0UCGzk9cR2kn9YsmD1JfuJVl9sHsjplu5q2GKhgpgyXkSJr
sInxRtqDcwpvbXI9QSijycv9xt+pyQdPkZwx665L0bSzlkVCJz3lROG2eGCZnOp+
U8eEaSGCvT/qjCXXkIps+LNFQQ3ZO28gQ680vZ/eLPF0EPPT4tq9ypCtzw7Vet53
mvTIhkUqpFB1j7vH7KZ22D1IZ8Pl+0tCAP6x7KVXaxWo5jADSLEphF8CbvVF/V/7
00J3Des2ohc+GSRoFQKuWbbzuGtLXpKZVM9uCYxVEwVsjdrpkc+eSbSoMSspPoya
s9Spicy2nwMIrg0Lfq6qp9TdoSbKdoR99Cqbeytj6C2J8Cb/XR+ybn/wVOOggueJ
uj9qtCzEelyOktAp49A96dpgGOnwIr9IXhYAsTJmxDkUhkAr2GGA8Vh/jTwUH8hZ
kMMkOVzhTbUk6uBSZ2HzPYHYWZ+80ZVrdUVRtKa43dKMrZIdx2ZudAA6nPYCNq3N
FuBGPVx7WcsPL/OwB0lgbh+2Mhx0yD2O7FggwmexZq17zckg8QxnltvrpdhwYa/e
ZKbP0YlLT5nE0e4JG8dMJix1GLgowhPMNRFk6lobTgsYwSp5vmgvGxu6v/aKVv07
7F7nsuqHy9Tx4mDpd+Sxau1JzlJT21iEYv8u8Qi/52Cgb+bROuTXvgu180Scpmfl
kfAt5mOZvUql2WZiYMaViOAOBYjNLwi/Vr8dM3lqrlqeGHOH7E/vpwUOE3f4AEVd
0jdbUrVxNu+C7EzgI9GBVIEbyTfQqtQsW99JmFeAnONNGFJkg3rznlx7tsj/dJbX
U6lCy3fJFXO5IBHfrzmA/zpmrEZ7ilL0FiWHCcUuV5qTDfHwFBN2AlXr/xAJZKqj
/a33T68RJc4E2Ya9Dcuxa3mTFctRN8onrS7SVh56hzen/PMqYeqViO9QWE5RPqBB
68SWbpepDMNixSMt4qvqz3HgoWI3VcxlEd4TRkix6zer4TqWyPyxl6pOk0sU9O88
P3+RIxtQbEL87L109Vr/KUVrfbIlgEa9oe/ZhpzlWqOQN9icxJUn5JMTo8+d7xko
1WuicjeSIKgayna2ZOhuHBqdGqjPCf/e+N2EXTP5g19GaZbOfQnXoO3i/aB4b7qV
+JFAfvRSV6Mvy1QZd9/SFPNFK+ysED7N+M+6Hyk4TtkpxkJRr3MBo9Kx6mhVy21a
f6yhJXfxBJ2/kM8Fcv5tsVXhZUQE9c5b8BTbeSPl+otesxpUcK1D1H9xFqXOyAEf
rvQh07KZeiVANnLwSaNtqGKDxHPgUj03XaRS2BzMOqFyXgnmxyd81NYo8/k2OYdl
eQLPWylqAM1K+IZC6+UwNUyQ7UlgcInXWWwIyXc0QfYWMV8pByh9yvYWp/SnToNy
PE3ff2jHssV7WJdR1/Xtstb9sdJl532VecRf/U0wzbbpaVLnqzylt0+pRgYA5nXG
rfdsl1ZWl8r931al6fXzlKRoMJLrjUjQb95/eDjv99l1DbRw8zKDvFunyUr4btvy
Ejodm4rWXzHdJZIHOXaZMdyi8hS/Q/FxJDd9f1Qgq9aK/PEA2uSFfYHMaKzxenFh
SH6gXunh+Ej/iVwxj7nsPLYNervfztP/PLfDuu/wyZt+bNqhBsZHD91bLL3bW7R8
NFvXuYyp8xGvMaVPyJ00Y3Bo/vq8p82LH2Elfj/hOc9R7G5Fh2VbE/AEKI9MtCSu
txeFhvSJCBVdKsZHohFTrcqyiBkeDLzFSXeuzU9IxMUGCr9Y6NK/qB6TmtoktJa7
zXx0g7xGtRFVQIzbMuq251hB0lylZqacsjVHeq8uu/NFEAF6/d8m5Ps8+i5R3DOo
odq2k2WmiqFCDddLYTD1ZsT4vYm9xQTd2YCUqk3aQReNx+Oyqj3xZvpJ6nF5QL/9
qhj/Jic7tbJcAxRlgUXfwqnlLkglJXAWQ5s0x0BCltgHAfAgNmgRP4JcNUFgnR5d
FixQHmBotVEGtrpMv9IkXFpZgqxUnF8TMp70eJidSwjvaY8ZxEQzKpIMzQ7Ev/33
4qs/7gYho0XZcLDrr2Xpa8QOjoOt79rN5Pvy60rxJ3A+MG91lfm83c2V7zPHHpLi
v3CTadYlHrGO2z0+zzmqj3531nTwdZeFoRXDH2jOeIblHNYnPG0uPPELb7b1jQem
jZtEk35u7U4IIX9RkGgrvFR/saiY/75dsDM8PsrR8QOZ+a+VUtfAbQhdk3nm6Yym
HaP3gcCag/SinuptkGn1xTjQOoNIlRNbI/bs9FPWf9VDYmktQCIEx/u1DMnNoX5R
rGN31fqcGc9/UP9zT6CoELo7gcY8zLcb2SyBvVyYhFnBxW0TfkyDmt5Xn+CGjM1L
vHeM397WBy6WFDS+ztHWHkVc4f4lXZgKg8j+bx8oIphvrz3glX4KePCXQyXXkEWK
7zhpxCLvCdBRd+7371mffTk5SbTD9Jfbfe/FFi9Gdaq8dmDcKF0Vz8E7fMsuEGdK
efbszi7YKUcK+ja+bd6OZMGE3AwxNB5dQaLCKZX2K0Zaa/jrs/TSIc2tMVoIyWrv
PeD12pw8+eksP5Y6qiYvRgZ/chEPzpu7Q3kSQCFvj8kfQQtYsWHwI3mLMSbGAvW1
gGlhoNNwXRb5yOBh8rQtG8qxY2EZiOJ5wfyCQTnqwnRyRJZXYA4VOAjo7LQ2OAq4
+DTmISzAeZJP7BkJoiyl71FK2DrN83KQRc2mwLgAN4z6kWmOcntsKzO6PlfZ7EDq
+pG43sneg5SaDau4l6/2TZzhqex6GBTZKtVr/YeVLb1XqovbN1Xg8QKFNpLiO4Vk
4jqbfSMdbM+yYbofaDVlKdftuU6+SvBqXWLSzOyXEmeoBmql6rKGY2VkXqOTl4tQ
1N5HHqFLmuwG0aCmIHUtDQPF9qj0Y6Wz0uhg5X191EUbgarf49221WpIh6nnSiLM
maEx73m1G3v9LTSWg9YXMlLsa8Mm9QexitjHQO5HrmK7LIug4LwrPUfxRSPa2VCM
Tu3gqm+X4Y7kjYyyCeYHNQ1Yw78zeFjx5t3Hz7YvrBIZ0Bd6ePzRDqqMFIWksfKj
bj6Lj7l6alcP2KzeNRwrk25qjd/xcCeNBqVugcRa6q7O6hk5DIy39boLvDdKKwf2
paITFR4ZaY8HgZFb4Ga9+MzpgIIyw+KLj6tqcojBdEXhmeSO0YO3rJR+lHkWGzyg
NB/fiTME+upB8H70P/FLfiy4dVsCSm6FVi7fCxpTfqu0S0EjEhXUfOW8vs4aJscP
njWIuxrz4NhXDSSbPtWLqWVFO+uE2/QMuxh0SGMuj5RW4gi2vurrJV0aRTFu7iAc
ifyzi98E2FQM0hJsc826HCPT8J+zpADtOgVAaKR4RjaoBi3yHraIaH0XwWwlioDV
OGp/R6CYetKd++iY7elsuHNO5Nk18vakXTw4B8+Q4vcEmhmPWZGx6998L6cDDWjf
kmhURbzz7lDuPgTL6aPxXZyBrkp6HtrBxTAlUG1Si303OwnhJ8Xf0EQcUJYuIbX9
68cTOb2wiO/BHGiCrfzfYj+2dhep1r1jKm3Xne+0ZBauKH0BuhTsB/VTiIpRLaUQ
LRk72ZustxwVwa2ilNmfnm/fdeIIATSPHiSb7f2blNF7T0+1aiXojCBqpVGfQQhL
kYah02U4yoGckw4toQ0FNOBrKWDQy4w+HvKiTlpA1O+su4L0v1imFYFws4m+CjT/
hZ14GtFF8TnluknHFKd5g/xIqh9o1Vb12QyQd6sLGaQocs302gjp7YjMmFNb4lti
JNmzbf0RKHUcCNw6JS2hqjeC8q5Y4sjLODdu97lqIIPsh59O4kBNF+aVv2v7fAu8
H1mkUeee1yds+B9JNxvAtT5gkRGJqNJdlI2N39NFiUj4JtiOXJxqrkmpWGu5eI7i
gw7JmkrgQz2Jvc4yxVtp69qCK1kBjKUSSRLPB18DHU50k/fA0fZsofJtUAEAsmIi
ucefiOMLeLWaysgadsUogPeTjpF0fb7CzOPx0gql4YUOekJ/P9fFf5naNRE6vhel
j0/KTIkYkEuYZ7JVn3FcTNFypXMwNBHtm4EUq71GkyTMZFiDEXZ2IirFGfDE0f78
aF2ocCFEfpjWnj+ztpEhbbfJwkZuTGFQCN7oNWvDZuhFuMluYiPH7/CULDANn18x
UVzka3U28u3JQgnUlJqtmZHWKkxPg+gJTRi2Zc7tlHtXy7VLiaiw8fYaRoRMUBXr
6srWtnOIkJjPHEDkwX3AGmnAwY/4en6yZijNLSZPCysgmW7ZCSiJZM4R5T77iZdG
UWc0OrsFcLCNxcKkzvbYrCPD1BJc1ZWECnVZBdYEPZjIX+Etl7xs8FZM2avZzlez
UgZKBEMpPZ7/dOVsQ21cG1G30qmwQtvDBTY5PLQd8OhyFG6yzUo5vqPemU+EvCmP
bsMg8mhtXhxU+Zd13ufTlnoTSBMBOk6/zY23tcKyyGN4dBK3Lo5xt3voKrVIpWSl
D4OMUT6+zt1AxWi87AK7FskiZJYIquLjNd1f4PiWL+91y7r15tVSM2kq70Ff3ksv
0CH3tKTi9pNzw6KncOhgvYI4b8MXJbNTAXSQj8mtHnX8SsxqVG0iJM7S9ea1i2mk
N+vJt4v3qZeoNhzohFJcW7Ze5y/CSLFzEj0xa+VPDBwVzZbttbfMx+0hHX/ww9ey
gQFuWs2Unvd9SyJFWM5CJcQUyqJ/qMDQYtm1d550Zq/uBo4UZNBHB54X2RfPzAVc
T/a1C6E5b4U1ptiAqa97H8bPUf/AKXrLYXbUE94gQ+kir+YGmoSWMeiZU6GqfPuf
z5b743f15uJGocgSNuA6wWiWBPdzIu4TavwDcpy0u3rAWBdYiaQ2fUz/Ln/ntYiZ
QLk1NMqsbUZpkeq5XoxPSmnP1PDABz6nm/9ucJ/fPdLNxFsy8plVJfd0r0HoBEwe
GbBA8chsC3fRxF5cCNjEZdVmOkY0nCOcKqpAc2+2I6DmN8P1RLGzwf5hdecW136R
S652l8OeDmP0qKBL/q0vdNIqIDd7EEPaGj+roBNxol6e64KYYA4yJzA9VkYqm27Z
Tpqb5EZ9L/iDBlbDtGhr74GqlwfzwWysOm1FWtip6tyueawAvwJ+w+bu1ix2URVc
rCdYBdYWX4IosGqBfIFrQ4cFzI4sbUULqUhxtGWkRt+uSVM83Wh0F01apC6xUfNz
OVhmTZzXJrYiiaBfLxvovA6o4JLxirmvuFi5rON6dv5iLr9YRzG2dXKDcyscNBgV
Lir7a9CeDQ4xYacDZobIiZ46+1YE2tLXpT0j6ZsWJKi7u6pA59Nosucxvw6unfIW
3WtOMZOk/zRWKsaG2Cne6AuuL0W1p6C39faVzRJKx+jhPl7+wVGzsco3j3H6iOZ2
o0X5dXVZVlE2yBdUTi7G6F6y20Ifec0oXr6LFFMfZqjFPdRx0Iqo1LYwMI2+1Yvq
mRiGxn/zAbeaeASUb8+1imWkMdE0Ol6Mdytta0sCjVvOhTZlQRrcGwftlFzzFWnW
Dxf/k4vkW/XJRm5WYtzr+0jMHT7uAiiY+Xir8dffcI/3+t4o9zzlwD9ow8lYFcqe
Z1xEyKKavjYpy8N8TVAjmWGBfS8rTK/hbsWAN6g6lt8/M4GL/k+IxSp/CGhoRpkC
Si0d8uA8kNyDN9hd2RP6KQ7oQqsyxzOrsT6O1S91d0sKRhejS2+n90i2Rl3cdvBP
2XsxoFBnRecqGSq04v3PkcPSoyF3HpoY5R+C2nX1H4CpXEkR4YSWkiQXSDOSjTrT
mcf6++FVtynp93GZxUkAQO/ZpYTudtYL0/C5ykLVske0CRu2WK1A9q6MA6RoVdlm
ZHZJ4m/kEl2a0sqXR0w0KnW0N/ksoSHgo1Z75LL+L6C2b2xQfBLjH2fBVUh7PIfz
g+1NmNKXrO4+eCfLTd5xwMo8HBltZC+3z7P511J5qjuBRv8hntJqKLIwRpjIYwir
Te3rIhNM0NXdodPrX6wpURvVgcFvivvW2roebjpoeoEnewibgaRrz5V3PlH4LMNj
GQC5eo2mcJskOME5JFpoVSfFm7aszh0sTOyWCaTH1sss7dfT5ZE+JRR99whUte/D
rYQhEfjkrOgrtBW87v7AYFnXi2bPBs/USx6uZBeldSGFqeLKmoM2s8WOq+QAlWaX
rH6hYvQIgQu9cZzGui6pLHDQAuXeE9bParJS31KRzRgoba8Cu3a/flp7LgQmvs6z
3BZo2iUWSo9pcSX6a4nzHdzR1g4V4hEewEwPCgzTkWXzEaj0X6DkhhhhxIamZ/OX
JdnVeU5bEzgV8Kfo2k0xKuOAUewzrp/VWy0P/Sfx5F0VplohSPM2Pn5V4HlEDF7s
8Gls9aV+n6B1mIT56ilNyTi+m5q1B7s0be9FVOEGX+4dlIWGoYXGYc6BW9Db9arD
i/9jmo/G+8FPa1aSCmlbubSEr+QDds4cFE7ylKqdm9bsYCyLjPINbt5mzcE2APda
v81BlEQjGfunT4YbJZqTg3uM9mnq8JELPzlJR73/ONp65jc4GVbgcbTY3M3j7Vma
JWMPzC63I0IgOihz3DwmQPtNMgg4Buiq/8b21O5ZyOPXVQ4801dIjIBzUDEUhbCE
a312AeIXdOocWYCcL7eXwAiOGuBmLakf5g728mi7Us4XzpRiFh1UR9oeaMEtA3Ej
rdFe06nD5pHvOxyUD47+7em6iWr4/mfwk49+NgUSpRL6atBJZX2B6GPuW8fPX/V3
+FTjgKaUImSEIaLHPk7ishjEcWDlPysuC3na2sTJ24raHbI4ce4O5PX+VfFew7Z8
1Cm6kD/r+o0WJMK5wBK6qCAxkTvGhD6bBGjVoHf0L2aDyPC6dqOjIKKgepShcONB
G/sqaDj6NGhsjt9T4TtPYk+6X/D38jNgWfDR+rmQLUk+oNDinhmR9f60Ya2Kvx30
nwrH6FE0fvNC/NdSoe4LMhUoUitLX9sQeqXTpwD23WwjCDhtHpdPdpXsMoVXC7uM
R3/0JQzxFBMrMR/en/0TDZPwIF78IhdkUxtYnsynBkKludtzHcsvPQb2lSe82x92
dbbPKQgPWqFvf8bMU8o701868HmQExp+1X1ChVIdLr8akeOk7aju4tUqs/vF39NI
fYRxTLxqkjVmfHgafG4+BdJEg/F5caw6hSxvcl8CowOsoSg4nVaG7BGvYJAt/WyL
Shtft0DpxNFjdOZxr2xXsLGtgf0YL/ssW+ldlJqfqSEP52NDoo5/+VOs7mGYghDn
TVrw70nASmA1fBxCVaQf7S0o9rGNtOnikgopUj1Bl6vwGEaoldE/jFAWnn+Kw/DY
rO5IvQnMiT9zB6LWbeagu4bdri7vVMtu25EEJPFRU/K3iLL6QmYxOuh0FPekqkQY
28mzVAyuSXNIL8QFCgP9PJ6DhKhE1BgZrcWotPnIlezOn9j6FBeUGrGBHTZH7hnc
hTwS/nRtvyODt75dfCyKB8WXqMit6HWUM+QmcAbcftLno+CsnlaOqpQjjlpMX2Wq
AIlb1+itjcEnojyx93CecJ7GzF90iBkv5MPUVP+WuINol4o/cr9LwBT8VFkturEo
82HuNqo3SipVorje1VpGEQTU2Tyg+CUwzL1JVoWeqb2DBbcfYmoG+S4iOsOFpjW/
mmoB+Nzjn7G4FTRjwdIgY6N2dKrPhlAz8zSv8oDyZPgQFBq0mV1ZfqBLfI7qlzsX
KuWnJCRsCCJv37Mea7TW3WoCkWL3I3yPrtK+dFPRJG79p0cXl03lkqBVv9hQ42kh
bJxAD2d0/wcyJQbowvbW+nfuCgSvF00TmbeqQVgyWVGdm9Ms1//CK517qFbCQ0c/
6ulrM+x3t8QeWLVcOWIeKQPljYTJNjo2sbE0d7Wrz/cIvUJMR+Vcu9iT9Yan6ryp
puGPvsxMJAnsxbaRLBlJDFVEFFyHeynOuq57NGawpeqe1PIJw+2D4A1znaBHjABC
pK8kZupWlLPAERc9i3K0RZrMeyUIxI1Ty/jy89I/kQG6PBmYghzQaYUwhvwkCi6+
Jr46MQs4i6IUaXIz4jB3x/OTbQw7VXumEktSLILRs7f75hlsc+BaM1VNO4Po5P5v
W5h276cqTN75emjKtGsdbTcKn//mk8FYQQgTPUdPjCQf3g5KYq61iZoXErZTUqZ9
qlZ1TdkeTFRtK9XBzZ6TgHhg1JGU7fmfufkd3qBfL72jVVLITLbP1mzswDOhNJT2
L2ZKb/iLx+MBuZvNsxHtQwdf7c6U61AGm0SvGJrbEBd7G+utbg3VSyaBag0JZxAk
AhPLI1D1mX2wHC7HfnmveIAJPz4uVwUXwD4eNn8LIolR9kpBE87ycjJLx3uGaOOD
QfrXB0aGiR0ZC35kkGPkb3qH2JajXEVajzlBrA/8hiz7voq7kE9ExPj1rLX9qS8G
JXDkwvdHY1rnnc1P47av6mVAAHD/qKfbqXG5YTwKejF34xLrzHyoPkR5ITqrqsrK
D8HHO4WThh4Afw+lIVdwlXZ0u0Wz5hIsLthZoL+7ljAflElwIoIghIWJhMRMkJ+/
mL0VVA3/BcfJ+mB4D/26FhGe0XEHGc2Zh046z0mED85YhNtKNW6VSaf8DLgh5ASw
yfwVEQMhaob66xkRp8/zyDfc4pEmomCYlnXmVqVa0Y4nuKkV1QUsSr6+74yxulxk
XOKZxNElQMhhobOODXNfD5gK0Wa/Uir6zwWlfeKusEuSnC+z5+R5/GVHad/mPRyT
6xi0jvYOrCVYMfXh70YwqpmHhPJLlsLumdkXa0t9i/KavtOxXZhYGbvxly1ESEo7
OZLY9e20zmnS28jYKmDeGZ8RI0oCe2NgPbFqp9mRKF7IL9gVn/hs7AZA33DXtcgw
cczrAXN4E1LGkyIsZGY9Bf7MTkT9DITMVwYgMr4NNI3iOc1XOPx4yt0DoVnroBwN
SK/caeKmshVz15pM0yd9b3UVBnkpSzBFT4k1dYoUyt1pfMwGr8108WwxKG+x8JMY
PpIG7Cll96xkRD7aUrjZafjIILc0h0wnEvVpLweazMkTkJ8An2iUetU0ISQpe3Ac
kq9BQh61IXS+T3fWfw26iKKVKad9EPy5R2NLbE9bYO7kQaxltrhjf43dN+ytpv4e
eu00xmXiUw3P0L3AeXVwiIal699w94sYTYfj9z2imbLk7cEMV1osAnV41Ma8foMn
KlBBmDQTG2GfYGYXtMeq0IqCm6DIYZXYFQvN3w5V/4RfNLsFLhFRETJz0Afev/OG
B9Bbqe747Ym1WWlyu5deuZssvQ/qhQt7a77dF1Jx8o7JlPcyG3Kr6xCL8CHQnv5P
4G+lmCzCrlBD9LCSE4uWGYc9cuign5FefFHn8Z3iEm2boDINLuzzPfjSaAUZ27OQ
PK4/RCpvLsmUWEl7edWeLmQ33I2D4rIrxzU++KbCWF9ovQ4+ZLuHXdaAUt1l2iAM
2MwhM+eJezsIyo41NBJWJ7wd2m3nkS42si1psVOrtDN0nsOYbSjaR2OFnlmlzfHu
noIY0GDGwr0fSQ/HCo5LqvvIkzVRCex9QQvaWotv46+ksEiE78ckxyBAaZz3JZ4r
/Jx7r0/3t/3FF4Ax/3jat4Vng4cnTuHYrUbCcM66I91coQeJU3BMxanKt6M5joWw
VsmTGmbdF5WWvwlQ1Wap11gnNPqYOUcjVuDzDSKZFiptIb2Z/9FaHsbco0rCfkbp
XqZ/JXUXdEl64DgMJ8u6GEJG9c6D2WYBNIvAMD6ZnU/oaXVpYFtrWopW3Gj1aZ/3
Gq+3C+jqMeePSJ6TboJ63dTz7GorA8/awW/wAQrdcBNpar3haV/sKhvFkCT+MPcA
DQsUHSacvBaoWyI/ti93ESNxvRYu/piHS4AasyZP58CYdxrliAeN0mKKZHQgpMsc
3zuzog7kIQFuEE3lcOY1OT4JwslI4jrWJWX6r35ye72g3ltgD2hQtK8Qy67TRIml
JySBDEnxMihMXt8hNKI+/dbC/USV6/6w7ZXJflBJ87Zpa9B0nqpBaPPNzthWUtRc
lrbaPyR3crxfVFConhZ+XFzyl+goR6dPqq8df3UIWdM1KNgK1SWQB4LZj6ueP10R
Nyp4fGQHQMDBfs8BCJcMgyXdFfAzjN/Jnyw5hGwFgTwu8SU5VMlROR6NlDYw78oh
qLo0ZwSkS5jNhCpMn23jLIJDq40HXnU8h80BAI0XLl62qNRitOYfo0VazbPeguNf
0N0IfGB9qfM5n5xo5BkeTpAmMACQro5BDTkkbKgeJnhEY9jQmJiL+686trFKCMxC
NA2zSq963kehD9Sx0AYQkR7PJI5UAm/2b1UJmb8qzSEkXZIDoNNsPFapZ7SC+WP0
iMudyJgVnRmo/VVB/DhhiP92pySy9un8bpOCcXKpeZe0cdcDSLvbPs752/6GZxuU
x8T+vZFioRW0oM1k3/bThpSiKnnuuqVueU854VUmSvDHEW9EToEeuXMZkJ1XxBBg
x1zEfyLGb06MYGId5WTq73j37g+MX4VQCnpYVTRUvb7DpxRd8ZeudnGcUafsJ/jr
6PXMgqUEPXZtn4+FR9hLqHYAOhlXPkc/USEkq2hfpnjLmed14POex1DoUYxEvXfN
wY4ae/oR3yLWbtqAecHzw2TuQfwAmVsaduMDjbyZe96hpjNNPCfYQTZWVoQKQTZv
3DNt5g1tzU40fgvE6MXZlVXMgvZ0VxTa23s/bcRLODjapVOrocTlxHtskJQMAyyD
nlEzjAlmJK9Zia0deoW/PuMQOB0jW1+2t3ZjBO94xohIdwtXxtvTDGB/OBsbYQQt
6Sh1756qgTnH9+YP6HN/zQM8RVsK1a645OxjSMmB1a/GQwKqnDITJPmOUiKzQK1D
EMYIVolGXquBHCB9qpQjU7/aouA5avtyeqbcJiMHB+hhZ3yCauKkscpwjDzGlckm
cHe1nIpf/Wcgx0htaw2HRtsiA7YfEMam+5Ed75A0BPif8UrPW/zKCaxrbqysFe6j
IoxcGW8kUAaPdniqY/BpeIrsxXRKL7TKw/zW8tU6vCpDGSDRlTbjWiISeYHmtEKF
fbNCEgD0ySwtG8dO4XF9+7N0UvdqoQPW04Cf9fGdSPtldPFakhcsnNeg0ySLByR5
sqU0u6epeMZGm/6qgtxyTHWpJ/JMysfMo0MH85yVvv041pN0JDay1yyEL9tVhgam
Mhl92CDGutxvOX04FbmKg0YjCLTyYtvXiwRY4lRXJ2YS5mvRmjLqghNRXpG8RSYm
i0VilzWz4UujWF2yDEuftUaVolaoxt4hFpHNMQxQRRMat0HhkLmB2kRs+zMRpIf4
R7XaOcmy02eODm8MBigomvqmtdB21bWVrIrTGFRUqOmGmnsSd6+wymhhNjAABQiE
co5/7O9/EghDHt0t1ki0LFdDdsFLE3TCgdi95P82bzKgPTKeOXPJd8VKl4GjAfxx
5IwtPL5sZlZ/semrK9pSb7FX9bP3bGnS9ge77fc7gvuG1vYoqnoPOl3dJlzdWZme
15XIjQLSJr4jb+iNZ1zbUCBZFqq4690yoQgA2ffX59SP6EGD2ZJhQrWjB70epxs0
BLXYTOGsQcAvVqdvSOH3u/0ISXUj++ATTx2kq1Xj9IY6XSvHRKT6wIWIz0kLlJZz
d1P7hEqjBjJGhuNSyYUUCDOsYAtEmBVmh2UFytaxVUWI/IX2QiN5me7C7rc7NvdF
ntTyVNIb2HkBJuYDRU/Bd0HpE+rZwGYt7ZfveJFoxNskzGeLqwYY7IvAv2sGvsRc
S5GUztL9fJ1NvEiursPLavUsaI4IPFk/ZoGwNw1qvyllvvKpw1Q5xgZGtTH9h6GJ
hJJhKz0YufB/3BdfUTlo82/j2Jjt5efQR85izNYrkrkfZzKsBKw8dDebyUoCPEhH
ohQL6G1qG1yzw+M/EPDiSp7edy2m6lEtWjRw1TU1SZ+T0es8lOhVnAgsaftj7SEk
GGfxO+G8UJUzuDZAZ3xHVujNpYg+KtLCbTfiwHko8xoxLaCec/XH/BTvkz5dlWPJ
TRsfTSqPRROIyRSQnnHWkgOOp74A/PLAkgFmtcfYNBDyN3t7qipQfbzDXONeqGxI
JfKn90bWzll4NTAxg5vEfTegm8G7BnnAZVQCXN3KHhTUQV9z0U+kVq8mXwfPPcvc
NSztL+jN0e/VFT3vorb6C0b7YBs2iWNRdowwHlLlSVulmWE6UY81+m6Wk6b7/cQl
GeNIYIfRDpW9FGPg0HuVq08l6uR4SQD/oNhjJrSWDIOrKlY9KqAB8wg+feklaSOb
pBd0mGGZLknsUcF+6ChHkBtqlIN20rSFYJfzlpYYkuu7DS2V7h1MCIC2fkWsAacX
ACrLRf7d1lvZeg8rGT0QXgeqFNlgtyE5dNRv0fuyk8c+5I/uxjeza5rf0xGt1NHp
E6LZ70kSZMEGUyECwMeraB0Qcg4aSy71dIzwi3+II+5Gcxehk6hD8I0rdfB2YFmm
Wt+sKCIYAsDqGRdcggYYHSwh/mHQkNVygsgeUn8W4Aq0pu1NTTfFv5vlXrS+5xHO
CLR8DSjvegSfKS3coK9oGw9F9oZcvjNBYN3r0qVkoJaL8QPVznAdMF/Bw46eRccO
n0TjsCLe9ReG/+e6JCpz8q8kC7pCvEPCDl50dSdqzInQCb/ri6tl6PkzgGZZsNR6
90AQZkmMVp9NEu2QmURApSA5lo9Lq1RBF0pXKlj4yNVZ1AUzun1Mj1U/RI6A7Yzl
WHqJRpVCSCW4igdP6DBvrQ==
`protect END_PROTECTED
