`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udK8hNsG9+aK0VHCCSmM3o5PbzN0IZBSz+lOWdMYS8CVCuBuOfAn7soDxc4BmFYe
PLQrzqUYhYF5OIjOSrwcHpvPkmKY3w8VieJGQxCWpytW7RXJGBz/fTCPX7ClcxSJ
xXEOKk9EIb94ig76ld9KwEjjLi7WD9JWWf5/9JB+RMHgrFCxzgvo8MvmXX6AAiul
yq5XO9ufNvKVS/0gMVXxMsbYDydXyAmc04e2shCwcZtKzPqlov1RXqnllKdYTpRs
+PU5dvwZCCPeSOCNmPdHB0TpCW2ZPCUDlt2OoBUGfIDmD5H1aH+X8aDzJDrNV1ZN
Iubp55yEaaQM260uc30ithFE1fbTk5zpQqYpJFVcQIW6m4x1vPgc/Pvsxu0seHrR
uu8y47j6RXCvT1QU4BxgQznFDMx7gMpZJcpG0w5lnPSbEsbPBCFFV58OvKTjCQpS
Uutt3k1RkpJUO40PoStqO6RkgC4lCKWmkITuO6u46JqoKCeNAfcogvIETPtI9p2S
IjqHwFNA2aJIjN2wTKPy1G6nW6C4gE1dwKzFMz5Llqc09RjNIQ0decbtYQ/kXIoF
dxUmnHgmE5TmgK8OdWgtsNY60f+IYuOEGWQE59DqVnRsKrBx4rETC1LBkcpk8Way
eeL7InR6nHkH65qIeQg770seD9xuGyXjsKQbIXqE/mX56lJGfn7gyizsM3D4H0Bm
MsA9jaA5qjXVqKyFbjYhth9cHxhqcCiY9KKK7fRX/zpLJ3oFJUdQeHtpHyvoBDwj
1vFbcX9k4qiV4CxrHuoSKo/zOBlAZRnCxeyJddkbJD0UHwEDQNjNJJ2yTSsYumvy
n7KVpdflZw9nkEdGxfUivtcSXh4lf3ix1VTBqNQp2SJLbg/2kzvinkMYcWS5dD+/
L4LUof38cbngiPlD5lvjl3xziRZNqbttlDpM3EyTEnfAlwe+CN/3gj4qVqurFhIM
LHsSuWi3SF1BbvRZCoOAnsEuHt0Ht0zhWF/X+kNqRBNGKFj+52gc16VdKY3jLphd
S3MJ0xvep/RlHlXxJAxd9xQYVz+l7VrJofWIRBnP9xXmYnbgYNSo6UGNrWx0DR1R
h1Ela+F+HH7b71J2PqiKGt6k6XcE9hrqqtn6p1z46zH+ExyjX6Za5rivHPw6u3lU
NuQetS3X3mLB/Z7g1glz183dFBIYi5ksGV9ZF4kSKnoiVp9yothyo5QwA4Ba2+jw
Ypt/qrCUCdyoUdWO0Vo7ZFN+3wly25VRSqsqVDnuGkSWEKG5jp7LJDjNKqGcReam
tXC7Z+/jO1twJ6fYoOFnqx7dniOBwt6y2ho54VTS3hyxUXoLDLubuUKKL4OyJ480
Hm+wApdtSsWTdNJi+J6fcy+Mxb3i3edgZWzsiiqfJsyCcwBqjlLCmW/6OTlaG0OO
Gq+JEa4pJ8mkjlFIHibl56xffj4rYUUNvhxo41LkQKyqFGo1lyLSwdjFND+ved9H
T7bVAHW1689d2hdyMY+UYmijlJyzRKe3s5p4Cz54u8E5cJsi+KBFHp7UVUiyBn6n
6CWpAYpAxgGXqLQ/fhW8VZ9q5KwXydvCYNicJoyGJiR7nCoWDyOWGm04HQZ8D6xK
UgIrgrhxUSxKKSulEAlJZ4C7cEPBZpgkmIhFZKSxLh/mrP1bU8r5nZ80UhuOnY5Z
eQSnt21yUFJOR7jRmdwkgm4u3EXzDVBrHk+MS67ZbSsEonimWaGWv23HJHvyUcIW
3Pdc7ur+6P22HgUpocv7QJEjVHhVbyCFtJJQ/9AZgV5QlnSHsDBIKlLyN+iDhurd
2jV9356GXKCb9yy+Oxq2BCWkziwOxUXn2alZpzn2hq+iS/L8sIZKNh6Eus5RvGL1
twGsZ+VzreAKMeOFLPE9k/epZ9u4rm4Td8guzTd9Rn+upsMVi1s+eahqHa1nF2HP
PKbRvx7tnVdn7mYoZLNAs7bSGiLR3mhTscT7G3ydcj79rJVfzB4dusDkeaTYiPBx
iiyGDXz/J33twL2ij8I+uqYqoEEGkzNvzbzSw7+ZMmLD81vr8N6UeM6h4Roey+Yv
eeip00Bbo/A9zQCO5QHGAilEU9hoJTyK9oTUsD/rn25DKH1wNBsIoOPRU+ggmT79
hgFm+ce++K6bKTXzX9uDhh11Fe9RHOtzR2+Ttp6eDSm4q1EZUPcOsqnzgzt7UDor
Rtuk7LFUqBcbbB+tcIZZYY9ZFLE5p7N/8A0E/5rD5xpQsvGzTSfqu6RXyZmV+ghA
ef1AB+K/hTsCjiwyCPZYGwe3nT5CY6wvfMFm5/nqO5sIwPCImJ3Azg9Z/44GT5tM
U09InyTATKWuH6XviMc30ANy4pWmSzC5Q6YTxRXru5twpfXdNP5tXAPCrW79Vahh
RvluuqeD79azwI6ZUSgWiUE5T7I7lMCTa85aR+SgO18R4uZ4Fei+XKY/dUNEJzoC
jldiXtceTQDMbzeoEd/THVNixOm8gSwUSiiWeLHR7LfFRy9dB9Ydc0I6L300WHiK
pb5cXHt0aacw00JrulPkXS3genGZ5Mi/MCaDuNJC+vJARerSwJIvUdlYk+GXLean
ITK55CO92ABPJ3/6kddWYwkR9L3RuVCGyuh74T4BnmSbPH0omQkTT2Iwg2ph1/HR
lnnkeIIZO6XQz5lhWD/IhlOkfTwYxRMPx8OBPvwzQttHBZeCKpDROWRgwXzgfNkn
A5muy/QuLuW4F8gBU12/2L5kQbqQe3DENLjrO4ZeAfVBpXHGqViLttgeioCC1lhf
aQ++ozZb/ApPll192LdDZA3h6LV32rgv1a0+tnVkHRZRS1/Q1OKaeVQa0vbqT8+q
OakJcS2rniRg0XDdy+jHAb5AmqLCGiNrwSDSyFaa145HN5ci60ABn1YLo6aoCx5p
MvIGNOpSwxb8jPpWPCWDIog/yWlc/KpHqL6LD1ep/G9CEyMrAveESzfaHyK9uEXh
HFlcIwgNvqtYKh33kxzghty0qKTRoX0HMBlyAgzOPkT/PK4oxDWj/Ix60pnASWqZ
mw2/v3ReYIm19a9tYf24R3N58WFDEFgKDGu2NQzM2M0O2iZ0q0TpRUXhLJI5FrhS
CKZKVfD79T2Q6dJiY1Bfig==
`protect END_PROTECTED
