`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zns+6q7rEVY8VhNJpiN9ZWPzdfnSTx33aNmoCPsvLUJNb9hXMnNAgyvpJlgSjtu4
cyhvaX+Kznv97EuhcNCKq7R3dXzPi8mfo94guj+thZCX9dllo9+WTcDX22viFoUe
ay8090Mk5vaE1Tgq3F1BTofpLNoKs+no/17sy91enfLgOx4RQRKG6U1W+X50ikYn
rKuY76Wsyai/RpJDDADXVqUglkgz8scU1TkmCpseMxSHqaK+xNRh+sTH/p9rualF
6QOXRuncWYIB+kocbSrF/oRsSQHEftYx7/GaP4Vu2wILKCH0W/nU2pnrovfHJdL5
T2XsSS2HmHUMueMWDRl11o7pcXA+3POqP0yIls8UASOyaAyvXSGiiVxT+FuH0P64
Y6pOrgCb2aQJKes3pUl9fLpu73QExFBeGs6M8Hb72aCCgolsw/2nk7UfS8HdWG5n
IUrKw38S2j4WCBhs8vGD0E8vCYU+iqEs9bP21CYmFTOql3XAJ6Fo03pvHU1Imy93
7j41s1NqoGuJeOjyupCuntM0u0vR7YSPuN1udeRopqjIuh8e/fF+pC8A9bCdLGjt
0B04coCSeoVPdg16VAHtkeCySlLe8MQyBfHNdHcNOSOeGeuLY9Wn2I4gHrCgo0Xi
mT0vfA2PD3yjcLq6Wp+FTuZ0bxSAuw+0Abbogzkv9Gon64u4DEQr4lGq/cihOx4s
eBGlPXlu5G32BuMTnWVHYqtqnkmuejyNZz6xdBSjq/qdFP6k8aRqer4IM673pGec
ZIlMj1MlOsUejXJexyL6HjQawIVaDOIR0KEPZ+12hI7KoOA4Njlmp3TRN27+RoT6
bHfn2HCNMupScn1ovNfaYOvY+Kiul3vVpdoljRTk/httJb5fsDnym7oeQn1J+q1r
NWEiHOiCadOHmTrwTNb5eSZYm4JrEy0FUte5J2k/tJuik+chvkZnv3A9bEwO+7Lw
z8NneO+8SiqdzM/jPE6wPlcWN9Sh3S8yZ1gSuuf+8aOgLoTb2FKQ0MIkDY+BMPFc
WPIOOcZ3ric63um4JLHOtc8nBMEDc1rCBa/axrJa9x5X3nnd3YjxhY30WoyACpZQ
Smkxy1YeTS/rTG1BJ8vS1QTintrhKKC+2xD3FGAwf7k=
`protect END_PROTECTED
