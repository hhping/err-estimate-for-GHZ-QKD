`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hE4pLnO6m/G44y0ZHv+MJqLofwWjhFd5VKGPtb0NGysYzvW8GAfyjflsQ+B/cDsi
hDekHpx3fcrqGdDRlOBLm3fEVdpAS6vPKiG84sNw531zgl54TDHI8W3z1xk+5uek
cE+xaCEA3m+Y1YZfvH0AvXzJwNVL7sQ38lGmYvnv5HWgoKgacxZAviM0s/fyJHhk
QpsGDMaPucP0RoEtRD4LW2R8ExLXb6rY5VYUeGV6zq7jZYYmXS7ivwJUby2w43g3
LJ6OCI+eaE2flb8Iu/E8FrCw7zZcDYQh+Lq5Jw1ZcN4KamzoSSJ5EclZA1MrVUrE
/25Wq29llUzpXxbFfFvlsuYKpkvkgny7LKHwr6z4fxYQRWW0SBk92w7GtuglbQVM
mH8M2Aor3SSFhVYszbhgpQ==
`protect END_PROTECTED
