`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuMwMiQgsBiqdOrp6H0SEtPPng/uETjOaBEbXJcBRxLv9YRLQ8oi7rdQDthXfETZ
3paGhO3TF31322JGNC+25MX06uSXWRv9D42BNe86Te1+N6oL7Y6WpditGJ7vD8yf
fCHDQCPXBL5OcqqPMaaGHgTMykxQVbzoXv/9FtCxV3Weru4q8N0cILeGGoJ+mHdO
gTrMIx5nS645CIDENp9fGPGGcCPZIuq2oH7le5T8X9goe0tJru6OGmX/dwy/baYu
5iigI4WRqRlNQZOUdKrxr7XdDYYCCOSrKWzpzW7OSMX18nmXV3Db16CAfsqE46wa
jeKyQm0llsqbIx1qi1wl9tSxpAn45slTAUPo44FJGGRP/MLSnA69JRvfpfQa4/kU
eXLwDcPSsg4umaNJ3V06JTCeUIfsEY8m31gKFeA2Hk4ddMfTCaBZxOoX4dTdYv5H
EHWC/8P2cZdJkwYcIEkl3kUtf/xBURlQzh/UbVvdCwbC8t7++s9uXY3XoFW+RTCm
vf4HosQ5quVWDie/bgi3I99V+KPfVQntyXKx/CC5Q3LN+6VOTrxOi/yMJPs/svRx
iJQ3BCkMBsYGj3bSdHUiwA1O+jB0uMc2bTtlddmuqYY2JqX0imNfxEAqJy34iuZ6
5N1MurTkLGOp/NVEp/YVQmcgHCdsFkDp/rrbQeLVH/mPUc/8s++r0KaX3NHgF3Tl
fVPx6Jk0cUYebAH3B8QJhWslYCo10kD2wlEYqDj++2PljEA2pOlV3zJGigLSdyvW
`protect END_PROTECTED
