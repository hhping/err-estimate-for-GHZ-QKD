`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AGh0uv05KFd2MWbEVrSrrQn8xYQGXqDf/VLNEsJ9vEUHZ+n4Rkep76JshE+JGuKX
W1L7t5g1JtwQJdhnr6ltBbdMqoI/8Czlx8XQ9dGz6o6VfdEBGnTH2UYh2QNgLXLB
pL1O6xvK5jqeot0526cnhtdeSxikT6ov2Hx8QFqwHlcxfIa91w5p8ctWL3mWwKb1
g7cCJymIZ4oP3xln/VzvEUYQlyYuiRNCzCP9Yfq8duT+zhk5R3/PMPoZ38UOmvD0
0wo9AFkUupvb4Rg20hom2mbLJYjTDUPIMVeu6PMwfVjJWMF/+EKZvjCQLdQ5g+w/
NAlWhUtHF+IwXEr3BtwbJMyqiWzxj1nWXjPzR+IHcqrh00QA5yXb3GMKeywlvdkv
ImysAm/XMbIb5QeIEC7hcAWj53Nv7arx8MSU4b52lK0nBMpP4dtOBmc7OQT4RsDs
xbaBEml3Ok/wIWSwU8XZncsZKm/y5UhyInr5BX54eMvv5askYpB5tFMB1ejmo2QD
T2xmg5SerUc8sl7CnFIseXTrmhO7z0bgOFamnYLrZzqkXKHXjy0tXZKCpjf+njCR
NAAn1m3ISvhf/dV2/cZFAA==
`protect END_PROTECTED
