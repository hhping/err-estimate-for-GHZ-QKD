`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbX95Kg7Nh+VKreM7Q3PTVoQ0CRpo29OKgkptMdeCJWwbg0MTzD2DD/OsDtFaV5Y
jqzdMBqeJKUibeauz1bNLxk4kwpBNNRF4FxXDbYH394rmYt0Bt4fqA0wtgafyX8Y
eHhbRW04FPocLQdsKpw5bHx7Hu+GuIorqE1f8X3tiLqMNqBGeR9B8xKzZO1k/JRs
pf/ES3FJsUvH9IbNGhTB+hPm46bQ4MzIQSA7O77vkNTSe6ROeCVZXzX1VkC3tQum
NeXnfRLskJe6i7Ut2ACDpFTQ9Xk8D92d/CzHqwve+2JtdjGryRPpgcKFNKFH1YDs
YwAlZ9mWsm+hJLRiHGESq6NO8Ft+/qvD9AVFAq1Qe2ECEiCI9ABREzXYjaOx23iV
+KuyRXw6guXVKTC/kU6bw066QIsCNbcBBHCZS4XTUj8wEhmvMBwAUtlZMxXK4Gvr
0aeS1VRZTkKL25MUvOF8zunsZ6UYYj5wnNRbhGNeZhWo97KP+JAxzCANd6shjk9E
5qHC7xu3lu0+XHi6cfejVRo+H8vpmm1Enk7brh48BBNvUMMCM1OA9SZarUAi0QGS
QTXcZkx1bbPfeFsX8Pqb8HtZk7qvqfJLhoAyaYbc6HmThJItbFNKpuIXu1HGrRo7
rOp+AgxVZAG5nSmyYdcygknOOUxTb6SrCqYsE0tp478tgCQjStYtZaY/VEdBkNok
ifjTQydmech7thQu4CpjBN0cwb6Jzf9WSX8jCQUPiyUBQGpzQdysJIERch8V2cvD
rtNB2c6EZ5WlU0cfKhG17rM9/zzY+G5Z67MEzf0nCJD24Mc3+/n0MijnSScIzzrz
j1dLn2kErGe3xIJuhjhdF+49cP8dRX9spouiRAiPBF5rD/aunCzoTH/HwEfF/mB4
DY/1NfscwnK9iSSguGF34Dj9uNBLaBgyIP47SFQLBzJsdq0wUK1yGn5+VY2CxRDk
9tEClGpUx92Vp/xuWZimoIf4PFUFRFCPUHwIe9FpwU4v4J3aAiajVrEn9+JLeLGk
RqOuAya6iVyPpVXw1cCNsPudt8L5Sc26AzxNBeoBG9SA2fvh0QCgrA8F25Uu3Edf
FzJmt5TVqNLt1j1ljlDPW4iK8BsFe+qp8lHQzRuMcj4oCR0mf+a7iVLaxS7JymX/
qypPDuTbyIqlrgDn0FR9XE6w4xzeULUEDIQW6KpvFLhhrf4VcaCQhSfQ0O5xDT9+
u/fviceM2+awac9UJYVldrtLuFv0mXUfoqhRp6jmjXJpW6cBqKMRbXCVoS5JQGbO
p8u8zFC/nRy+S4IZEM8l39lNbIP7M+MViAqoU8xCcghYBPwc6Dm4xbBNcFx70L10
D+tKocBMcvL0t6w41TPDMNiBWhz9bxttcMUtocVt7IMkQWx+7o0Njs38aPTnHXO2
B79eQT0rs5diFytOG6QWdU0Y4ouT8W8nMAZN1sH960Y/AfbTUuNfF1wsOeLe0V9j
N8alPc+RHrDOMpDuXPmavLVJwG+EznC3H9I3pjXoBHNKHoplXr5YPf6osSVufS9Y
Ji8H1t8i+8GOoL1yGRjWpwliRRjzNkGu/tybQ/lyrRx5ftmxv9YoGnR0U3ixNWqN
uZw1N+4mK73nkP7WcNcmr1NRLawVivLRGc5cxC312iK8949pXF30OCwXCPsRZ6UO
qQe3e8GUefCgLg7gKyYUJd/zRJfHVUtFmEhdCcGkaFLSfSkr233CEgrbC/DY/lsw
/Z/2MVxk1nnlOrztYdVdCYvi0gM659cHcUOf5TOas7g2hoFy6zt7+hqy4/1k8HEj
y9DHf68Aopu4ttWs47Ecpa6UoUprfgZqmRW0vJLsbC8KEgQd3lqPIimRX1nso6DR
OCDj6AXair9RHm+n1H41ek5cUZNKLpOgnMGKmnE91HLQkntVUB+63HU9oCHRw1R0
XLl0bIWX5kaU3PdhDS1BF2R0nwmS0Ph5EeGSYuWTZrMvcko74bLKMdjROtS0xJ0y
Dh1kWv6O8dxcnQsVQ5xamPWX7DK+xfXza2Bl25cLJlo510uwsbj7TU65R8njJCkI
vQAody1A9LOrKY6sHEpCpTNojaUp0CSl3BxgE4wTFr+UNVpF/tj8VHy8Uw/79ZfG
EFKDvcneoVW/5j3luViBYrvRYK6kZaSQ/ufGNidE5fjhcXb6lVHqH0CAnXMQyP+a
O3Wq/lfsE0nXbuLfYrCZul4GTqijGTYwHUyBN2cSTzPxsRwto2Fov5hUCCsk05Ov
OidNJsGUTavk0QNorl27moF6HF7qf33J2ryWoFxGf9CTvTzMxmq7WS/kKb+/T9pI
hRhCFcrJ5v1TussadI5K4J3Mbn14J96VszVAL/vP2YyL8/Ne7dogrWCDs1jwYyrW
mCOniqPUnNDI8koy50sYvB0kaGzPynJeVSSJ0yCkc34ULLQPjgohwwtOTHICGYCM
jHG6wozXiTu+IDeK6XtMhmRU6R0jb12roPFDG/SmoBtJZdVN4Z24mAfOu/8QflBS
5DoTBXEFV83wH4UoObt4j88hJjM5gzFYccd2pn8SoKqyxNbVC69rT0p77ReD4/GF
IVBdBMrJYQFnCmBNfgq+vIG9RFAHchCp8LRXl0MnnUJgcrfHqJSt5Nl6l19M8S6n
t6b2Z16912Cn+8nQEJX1wLaoh1yHLzqwYc5CumgAOvYlLRX0TV0w5q/rXSqKeO9I
00UayZGTe4x+LE6JDrJYWkbP8j/CyqswSsk2YQ6ysigpZYFBKfj4eiOdpRGZQH0q
MHJXmmLB2RBlTPjPYQhe4/gb9QbFTVgEr8Lmk58x2L9tOqdK4y/GRie9depFrKdk
9ftaO5abzGCfzA9MunaKHWsZ+nE0z/BN0BnP/SBmKYHkNQi+XPpax1ULo2wiTwRw
0um3iesSbiKun52J31/AiYy9CmPdm5wY+i7sK9qQJluLeUiGJFURKgC+B5O4H9zZ
INU48PKpQtVCvgAUIu2yLcX+sJEvCWN+eWqJFBPwbwZb6by9QWorNJD00dhPyacF
cGBglHIiBQ9XTot9I/sAtw16orjKoFNyMHHOgyQRneSiYHbDvedBI6gReiwtIVeG
6ezeHFFCyh6wx+kM6FdGq8x+bpwMxdydmA+TxKLjgqI=
`protect END_PROTECTED
