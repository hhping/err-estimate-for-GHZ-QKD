`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zo0yhvehE2nsbR/gBljM6EQolAxxxgkR1tQCKd2jcvGUpEgeD7p5Lfm6ioxQca2
13PyRB/ycILAfT7+a2OZ/Z2RcN5Q7O52QlY32nDvxvb6j946FmjKnt+++16gQJfv
q6O+mTU0GDnKc8mO6bWr9Qp/mX4APscb4CH4kMPwndzOL+gsJcf2WI+lh3rqJnSS
xsYNC5HIP3i43uRqFg2wBgn6DQy7q0r3F0GZ93UFy2SfDt8nNcUs61KiKoeMFi7H
FU02tkmoFgQbAnqcx3UoyflliVOEtErw9RxTJpcj6aakR2YpWpiR21iI+HC6ZenI
DxN0tn8uQFxUgulvKUj/+EtnqKwRfbQ3hhghp1qlmRRyKcuK/Krz8C1c/tnN/kU4
P12j7eJZwbNYFYtUqg/ep76id79a06hEFFmKK4BvKswWKDJqKd+K8DJKDFMDAbdA
BTUR/lh2X5wnwzZ0l+sKzby+DD+xYdXx50yOR2jO3JCrJ6zpJ2F+YicV3zD/82S9
PVee9s6kV9FK5aNUuQQ43oWlfsQUspQgeCm7c8+6QivIqvHxaDp6ZebnAJZ2oZ4I
vgrwZurQRa2v3vUt8uBKAf0cLRXXmkI9s1jQfghGxrxM2bC1hFdtEiUPqN01EH8e
QyqQ8mDz8qsduJIKs3LM6ZSx0JwHFJia8SuZEx2ZaaLNGE7lsDuz32gZTKcg7ayj
myoNdrPI+6e2QWhwZW7kO3gSfBxc4bKFq4Ujkpeg41y1biZhmoubtb/eDvAIoi25
BD3eke4WRMz+1f3q3siz3jC6E+Keo5rbx5raGmllFn+1ak2t5ynT8a5OM9ghPqh5
iMCO0ObEEWu3q2t8jTTvA4glphmOhADAUJp4GteCTJ+X5GOlV75/FD7RxOHCjWww
E3VPk8+qi/4mK43uNsHA+8IjOtX4pnL9nGl8pcp8ehIKgwl4YPOczJjjSObvrJua
6wXRQfJ/niQwoiJIH8R5YqJO0Nk6hVhwZy+CGugR/qTOy34PSMUaQsG+FqlPGKrP
jwaqfaeSnlp0A5yGoylpSqxRLBqnDAO9ZHQAMpw8WsrUi4ySfZISPKfYCjCPrwYs
OSf0mCOlWWoNsay2uA9u8PdI22KDzODMDl4EB+gR9b5i9/XitXlX2+0GhL3AO+Hs
3YTNN7GuQ6q7NWK3no41V/qLN0ANlPnc5ODHkrE+9OQACQ/LpF61cMB9RGIdJS+l
R8WBam6bugXbxiGbv/ZMwbXdYibbH9kemfMXYpSYb5LrWm7545sVdVIdtG1DKe9h
0+Zp1b1Wo16qSYPRLpbIeiWZ/CQVlZR80XELBCOyxTtzXqVYJ7ucpMwuoghL70Tl
VGV5DpOZkV6S6WeBlqPDbli1nLx88XtGXqp+lcKc1un+JYiPSI4r4kdyqVeuQE8I
Go4dmwd9otvyRIhQjPh0osq/J0NxYkoLJELEPuLP17OjELt/m2PTc/O5cLgF43tN
Td76bvdRBGH7HKg3TN8QviaJDHDGA6LF6z4xa5VHgQbG2Z+cM+NQ8x0kIzTE3hXh
peBZSsJSPocfbFZoI9ocw1ZxgcjhsLdW89zSBFzEc6RGrMiKolwi/HVaWp9UAA07
idqjuQT2r8MJFYy7TjJwkjZU4QB9kaoz6IHRBerNC/Oim6uhiUyTqrUYvnVJpY0C
xi7r7d1BNXfvXtvqcRNp1fo/8wPUBeb/MMY/+oGdpVRoqXgtbcB2toctxQjN+srb
EmAB3iHLWZLdoxy/0eMOYH796miBOpw3lrhqd+/TcpFfPDUh3k8IcmYQsQArVv/H
2A8iAIrJGHrFE1zMf7mOMyNVNJRaLQc9pSf6C2opS5Xs3gOIfjog7tQnJ7JBjqKK
HrdOfHsrava7/jUm6aPb35ZmAd+xaG63VT3Z9hs3bmj0KpJ1ZHR1ztp5sTwN/D3T
ebbWU0Hnxm7WAq4u8KFoc2PXaGtbNEZEO9ag+4xprfQgc2nIU/mIr3BmrSpXjgfa
I52E4Xx+QnZbd2kX0mlATuRIlRpgwQfFta0VBWFanmZYg+fzzR0YEwLfSEkvLp3r
HiPGYKx4ocyv0qt3k8gF7LPG4ie73SnXTuNOX+/ra/izeSqYcJIBjr9XYfUc9oVS
UaGkUwyDusSyyZXR6xN0Mj2fV/M8zGB6VPGeyZMbXNSlL/KJAb4ijEcWnl49P16l
oWMSky12G/vhN5VAv7d5pg1Z5zlgAw8fC4/4eVIuDvL7b5ajtpl5U8XsX0r1csNR
kK5JEda1DpF9IVOWn63Ug/pRCRwVJqVk+xxkLsCbi2fWlhGlOsOSdgJKDNtnEY7I
W5NphMRWAxFSYCRNw2obUdrQKT63ZkQ+aaU5ZKsy72e0Vef/W77XyppYRg69ZZTi
wK9GTYOZ7fv1oMbUmux2I3YCKk707acOOtpKigvKFbAcz0QN9BEonl+CsjU1QK/s
8JEtalWnbTOe41WpNaNDyrT08PBxU/G7EG8Po1M2zDTrBQK9dNij3BEADSvXgMw0
VYxkPTs53eTOAy7Abuizwvj1mWwzefDAWJYZoPTpHmgKovkWtQT0m+8TH3993cRy
fVv9/g643p3DAwRgwDk9XUTa13f6SIxxotMboH76HVjjuVH6A5bOrTlCIJnjBWFF
8qfqaRYQfDdnscyj7ex9aQqjg0n+WVd9OzBHSKGiag/763IUnDrg4sjXGjE8Y+j6
zssUYPwHs1zkwHKlf6dpew==
`protect END_PROTECTED
