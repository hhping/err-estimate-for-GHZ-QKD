`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cb35Pw3cDEHsCS7TPuBsqaSMzC+R9Ku6zV91VJFakUwIGN9G5wQqmhbhqzcmtz6i
OBcI0fxEd2DZDR5B+Aik8HVGMNm1OtiwCRVgxuV7afQRdvSDH6S472dNvvcQXUXe
g59qyE220+ZfDelyRNcQ6hoIbLG1HeDOSr6nvjVHPSDQM78IceImOyRsLDcZe8WF
w12U9HC923/si4+nPzKgyMfDxiiRgR+oWrCaPiub66k94y4853VyTg7n1AIU3iXw
vBJOXNHuTGfRYyPVfTNOaR6wfYz6sVA6GcKWmm8Qse2hMFjZNGwLgVe94I2lKgVv
/aFd7R4wqZjmeF/moBJcDI9uYxzb8q+eKO8BfPdWMGfV0t/O9q1Odq3XO8zpS29S
tc0WaFjIkAsxr8rs2yiYtmzWZZOCcM3fIqx1mEJm8WZnYyK/TqKa4/MM+HKdSFJP
r0hT1842MaTcCS9yCcdRKL4IDU8uiryQVAjHcay98X8IPVrcQQaVl6OJZQcAe8NV
2UG0eUBGGuykZyncktWGTAXjNJ7Nd3GP67mKl/cecYqPj3NRZSV4edvYZ15Z5u04
bsgf+zdPP5hraUKVR4DyhRE7R0RanvdYRCVfsbNtT7FbOWyRX9fn8IvA1e6orJGp
up2gvhsHaKlle9//OCs4I72h21rzMFSBb2fx6eOVTao0qJdFhia+gI5ylvsjVdRe
smzyCK41UAX2oRQiWKsELduoYExJEfbpoTp8rMUVxAjg05EEQqtD/DJ/QtdmmV6R
do6zFd2rDtEeoXqHSdwa5K0utGAceVvi11gJXsi0LnfNsMdGi9aWTEEQfm62Jrmn
45mo3rNZzk3UU0duYWjFr/GKl63CkKFIXjThWUnjIyTwcwM6jPORWS8xqQu/3feL
CJJUeAKrWNU9xKXUPzbjeOHt8i0cB54miI3Mmzplng/gCgS0B76Ea537krfokUoG
HZn1UeAIawuYWe+FhzBR38Ezz2fImSZ7jdKxakR5jNexwFRHziBFmrmFx9VeC7oD
CgR23hCgitQQMerEvFlf7Ok8ngD3w9r6Qy2KIEICTdu+rMfehMpApMIetlSils+B
Nv5rbkG2w6Lr/k6npP5vTD3u6e2tnkWDnpEKnUi1o5+X8lhgCnOjHKdvogrxV84g
fuVs62RPaTtY9WYzonhd29YfILqXGAw71B827WB3+3D/oDbFup64elROXcWieuRR
iC/EOWBCYoxR/eCdJwJ51TgUTCna3idfls8/kTsA5gZwnEMDysmg5esWBMDYsg2K
6MI6nRqOWHSIaeR+aJNtRokMo91c4wkaVrMiOKnOfos=
`protect END_PROTECTED
