`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fSljs/p4blEyEqjztdYWadJI4vet8pQzxkDnythiOUYQYled1IcyXqe4ioF1YEg
qrq0RfHFD6tpRYkbdHLe3BIFjvWIunxlmKf2ImbMimLDhH0+qK8pj6W6aHxjxwSp
bejrPlWWsSV+cRPYdAb1oYf4CBMC3f8VQLXPi0jAQGbUsMW1iNOPdyIs8JOZYWRY
mqlfqqC5VT9crDJ071ApTSN+yvzQEl0uFQOxmCcbjenZQpPEOMIg8ttfW0tmMWQ0
lHfjt76G2aJlwRVIOOwQrp9+dXrKED/3SrtYAmOQr9WLH0G3zyXRxepEYbwtHAwT
SITBwT1L7dMMPs2Dui45sxSgf4CcEEhptruu71w2Yb4YnckQkzt+Fi576sB592rc
zQ2UMj23XD99RtbQ2V0J/Nuj2rd2fnKQ+tGsvGXLKNHJReINnAIsGB2vKbv48bVU
QtsdISaPfA9IaZMHXmN7dBYc+obP0lB9gsznnfhC5t9rpaJZt/3Z1dL+vkTXEPvg
RESkgjjQa5T1kP1hBIRpk2ebBnnnswPcUOAR8+g2InPeYN3fN75/QsMVPjW1c2j7
LMaohl5fOtNX9M3AxSamHYELeAm+vdFZ3jPiVyYpgufaKWMyUQ8fXWpkE/xDOAa5
UgF7c66UIcuOkTssX5tewMqqxn9CkQs3XHQJ0nxFxZrRMbsDmPaWeBjLxkdg+s6O
jlhoMUuAjgpsQPeB0oJdYvUwv2KAiOtYXXtolrI8+AI20mzoCyVU7wfeXW955MYn
WhB+zx0gvEGZs37Mh0OoSTpk30NuXhVoHakAsBUcMYsVr/yqJnlno5HYMqNNvWHC
DDoZ7vEku38AxniFAP3tl8npmBoGRfNQ3ZGSCGHjLZvlqJkfByV7JiycbGUJyiUS
LJy7YUz/mJVdfi1FS658XmKQIH7VEFsXgpR6UOk+EObRoE8jnHgCMiR5U50fhAHF
cYejEmnjmwDlEZgUS/lat4S4BAjhNnxaTo+MLDJLt4qIomAeL/lL9z+XpDpRHGnY
1trRKTxmlV2XuWZ2FVWuwVtmeo6M8QpnmrnNTCOHuXgaESkrmVualvp96gg/CFpq
nE5iMQLg+TNSviMRsRtbzuR/HFIFS2myNgpTeC3oClr39GRZ1h9vJXCEWEVF899N
63DcOupq9mFYgEWdFDpE7eDlDWtVHkXx89nYrR/A3Uhn2Au90EmGC+Qgyza9rYtP
o6g/qNYgmmYiPTtNpH8365szGDzlOMzS+1B1rB9ldQeYI+jHxURv7DmC0U2iIkRZ
ItZHRR/9X5QTfQkVGxEPDAwBpxQGU6BF2OeyEiqdB0HOWJtlFNoVbPh61a1juxe9
kIGlUURRmStf6Y2uwX3KeF71vgBIOyPDawiDpH6RGLPeI0e6ulyYB/nEh6iacJ+K
Gdmm0+uEF8czzTM+OtCmYRAJN4aCfwOCMtFJUKUxzDRY9vZPoEOUPinBKmvLRC80
YnLKjlfO1/skXGbgwNxvwTtF83hA8iKm+QB/isWw610=
`protect END_PROTECTED
