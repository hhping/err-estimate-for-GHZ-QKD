`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mtkc1yAjtfDhGTsna7m8JvwEaG1h/kCJlrT1WvQ+KXLoJ0BnIkTBhdaLHSANI6//
PkyFoGiC7lo1gQaXqNMZfvv3HAvC6WI7GNy7MyqAexbHRO/CCKWNFAjrVDYHhmNA
0beZLolTgZ4dbd6cKnaZ5twrrBnBmxU29i6VYH2Mm4Gwwht2ungFhRQPAKSCX9mu
eGoxOtJFYh/08f1Ap2pM7xxcJFxlTKKdnxtWLzlrFJkjDFZRsccZAU7xYvhaQxyE
jgE6d/PDzRo+Bo+cNMDG7EsvdMAkTZp7tpd0iVMyMEJKz7+A/4qJkiQENC3ScSpp
roypor3z1/cCzLeJJuprwNVtYwSOcAGyPQkgPwnNjYIt/fnXWfXXMeT4FqHKJT7i
Gc66lSE//OJETyy2jCUA4fSyhIp5i1z1R9eGJ4vv+/92b8chIzued1h71GphiuTT
A0Rkj+L6vYj3HnB32G9p6W5/8M3T77qEwmuw4L30Lo+16vZ27FIt5rVPBEI0Pt3s
ltQJCyN3EZs0UZ5BPCUNy7xjOGkMfunARV5SAwqYRgcCcG/2KgKiyMabUCgSYp4u
TvvwtbO1Er+YVHmNngFMDdsWG3uJb7EdBJQO6yOv/qat0dokARtc35ZgFSOM9GQ/
E9KEH/oyas8B/dusy7OXlwcv0CGWeImklfgcFauTEnA=
`protect END_PROTECTED
