`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3itwBDAlZqtlCgwXX6HeDJnOWZBSJIJT61oOLlOKOk4y6/6YAuUOgVrfHx7wiKOK
x2ImXLHmgVExeWiYnrlZuptps4Ly9e97ewsfGhu2gLnP0XmDIS17KCM/IqjVp9PZ
Xk+MD0RPqbhZACyhYz2MI76xiqB5/qOXru2UOKLjLr6XT0qM/biR+7XmuqcDHtoZ
VZGg6KSME5B19xIQ7leuMa+cOSJIYi4VKZnp3z54I5URJAyE76B3eNOKPhFYs9VK
K7Be3SCvmI7HvLzoBKrPrJ56QNr/hcoCEAG0FsfAQQf1NAzIwGMk/yYdSQHxj5Fx
0zpZlvfIUYOGPXkOcfkp5qvw7v77RTOeYSk2Z162hs4gzn+BKzF2X1tks0ymFqr4
gcbwKZorjF8b3bJXfZET3KaKfobowOZ/FeO/XlegL1j0vE5KxdclNE0q4j3/qXFw
vMK2L6UFdhc/XamuX/OtXQ==
`protect END_PROTECTED
