`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/rq0iRaukRk499V9X7LUfKfKB+Iu0+HP8XPzE2JepIFjDzjBOLzAFjplvdb6Ehx
shWte1xU6O5/IhgXLiF+18oWn9VDCf/R+RimxLkr6Kdtf/0BPFl4GXko1mcLf6tw
ZaL/yi1/+vkm9twvmhtp0Sv1Dkdbu6bV9XyBD09vFVwDdgMyMuS0Lidjy/diiuDv
Hbxnu5geQkJVvRQ1LSsFG//wvO7RGJx+clwAAmGI/RYiOArVraWaZAmff6DtHs2W
KWcx5ZqCT+6HdJ5HQbAdbPg86OsqH7o6AokkOEOzNNdx40LiSqTAPjEzoO0Yo2jm
Ijp+5600So0DTZTx1De7BURxu9ag8LHHHJ1Rg2LWkEXDQA02rvjQ/BaNZWSTWjAF
66Wg01TlG5Wv19qKtmlPfs/BKaPwtiYzFJy+bJlLp5LfuEKhxNxOm0ReonWbggTJ
GNBvanlKaSAvm13mKwRj1EonbTnkrCeSldSAKQ8hMYVyk9vK1W/eyNZ6m1rnUvli
fw1UuIL7aE+p7U5i4tLNDfmQIUL98pOFiKrjynQ+OU+B1JQ6bucgj7k0OYcqLRqZ
7S3/eiRGkkc4G5tHzN6yeHOVXgVveWoeGr04zfyOJ21/c/KEznPy8ylT7eqV5cf2
mApSywqoI7LZLpD4SVYkLw==
`protect END_PROTECTED
