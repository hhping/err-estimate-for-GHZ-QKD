`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+Y+N4mBnO+L1icmzZMRpk64RQCcV8NUEGLX9oBVjtvo9oztMzdEUr9WpIODVkIt
tebr17rTdY+Z82EvGHSgdnYitQZ9Pqsc10X1IAl5lxc92h/2flEf8akleqQIX+y5
Jut+8R4CWaJED2jcw+DsMBPZIvimIAQ6MzR2zoRguTUDFxdcIYZln0d24cKAqjFy
YfzWHooZVl+K/f+Ld6zUw2A+ptafDRzYogFU261Ek1V/wBx10j7oGHLRD70Uac8e
Dj+N/85uS1ekeZnS8VeBTQaOwxYKMFGM0L7hl+MifHkYsXO//zqUjtIdchxmSLWN
rxZc4DTH8ZzFjqmDEJRYsksMLZT+sFUIWlA2qcqxxuQOAaT3/gb0whSORRpxkULN
bq84ofSXXIzvHzMH0S453rmUkzjp9R+z/eFqyB5ip8M=
`protect END_PROTECTED
