`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1a8Fy2ZIIJOQh1/4NvSabpIBN2mm9OFh2zPQ0Zz21T4U3uyTe8gS73YD+eTlcIIq
3s4IqdrdrWK8YIc2e3Icd7jC5ZmoAZKieA9DTzBUv4BK9sNM8xamh/iO7Zd6xDY6
FRyr4X+qy8AKSrV6KAim7Nghoq2VoSyzCvG7GpMZqY+3+74mmF95+USyzQtENLd1
DSDEGKXo8Ip6YdUB8axIZlAlzABTxGPN6EjkIbhtun/wXLgiWKCBXmb6S7RhB2Ha
yI6DpUMf6hMbx+HrduZaxZLrboVCk3GY4sOOg2XEVKfJS693VmMA6bwouITXK8EX
7PoUEhD+hA8QJZoYCLBHgQfIFYn7bBFZMxVu59lbpNy4Qfm2uMUrdiVtQwVAkrz6
gvO1YS8rTo/gwoFRZJvlWoAB6VWhD9g8EEMp/F2P83CStUEs4AjMzRHtg//BWfDj
eV1WhP3Dv+Obtj6fGHymte1hEq+P9tXHDga2sHDMZ/n9FHVT8RKJcza6zUTQSL7r
Tnuz9PbV81ddu0RuFw+AhVhamm5c617qH4cpi0U7PefmaarNawiwUGlHsZAU/VE9
ZcUtn+c70zA+nnQchOQoi4hmpwX0npD9ZhRe+odkRWUcxAsGLD6vQ71maodKG7aQ
LIXDIEBLdggI/B4YFlBFjyBt8WucbExrguGq4e+OIIYex9A6ZX5sAGaAh9e+HCIh
tVb/UUCU2cnm+zU7rslhTutloqSFLXNyTZgSFSReeQ8ByAMsCiSJ+wqZ7nbVbtqg
muSsMWsWm2jb6HstQrQno42nkV9QJKIL3IhjMHtgeqfMl36mpVS7IANXrQoyvzi4
6W+eQnb7IX8R/Au6Ex9C1ZXqgX5nmknq1mgEdYk1w+A/aii8xzOZlZv8ywZqd+k7
MrGm8x3quksHXi9Q8Ocb88oQh+DXmSiGu1UnZTVNjvR9LzW7yaOuFSjIm9BOqB1C
DL3kzrh3TrjA6AvJOeXjrgjceHLxtAWM00wSga7GvVIMb/tN2C49KX7o1dLtSZJS
LcFyRos/3lfAC2RNpBniT3ymgrZqYw2lJOmHSjjcns8/NzxrHeNReuUOZCXiNisI
F1NpSCMmFwHDkQ17H9wPcnqVBCkfgRtx6IFeXx633kSDZ8zStDq1qa0zuneBrF8b
`protect END_PROTECTED
