`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n7/9CKk89hOef2dkBKTM5FRZ8cTtZ5nf3KCOq95VqHDibBizzh+VizZfgJ3uZnPv
nT04iN7gWbQfwFBP/GOQpbAZJP/6iz7x4vMS+Qh8u0eynj+5T4JD06JrUPanVPmD
uxH3tImxPruxXl7/Ic6jYQHTPd0iPadjl9n4e3ceIk7BNfYUlT7j1ZkrudmVySHy
qn1K3WYMBLMTdLhJhNSzGeJ38AqAQxoB/mGFhDV2FjVU1PifxMwIIV3n9jOXDrp8
icd/ASMemB/TjFncPhXoebD4nvnzHikqnZAt+T7KsSWZLJCiFbjbNGToqPs0g61R
fER7IP0e4WzLaRm/aJciK7oPmyeK9H00yYbAxQhFaUWeSb2u7TUQ98Nia5s/HZWN
4WEbGVDpdXA6GAMh2jiIfBnMta3aJCR2k6dxXNj9GkKlymI0iQa/xG+NkegiVHko
F/QQ0jLiI5EAAJ7EMqzgpDWy83Ie4rNfTS52s+CiieKGtt97UywXEZDdYLYb4uAM
wAFsMnd/2L4Xrn/JW4+CiRbHWw0qe5TnK+NiFFkdu5Yld86Gho2J6ye18vHofWW5
cXQTiscLjwnEd9srBlErx7QrjnqGp+Urh2Ai3lwBefBhYXOtwHKCsB2KJgboVU8g
0843PtAXK93i/SQQ4oI8DKpvpUzunGcu7N1MQlUNv59GRsIegqtL7PiQVDKEPY2a
uaBse1GdHwYDU7CHYwcTdL67yUYpTwV6yjnGjj9M8uFy4Itadi15WJltmGQHUMqm
t1zAbadVlCB/ajXMiB59MvPD51uACRfCCZMzLbJRfMIF985crodGKEGAMY0ISMeY
ngA08x0k1/oNMlXN3qwoiEm39CeTaQEsywbpGKaQ7EN1e89ftMH68pDxL6ANicNr
IfEmmI3Lbny5VdOFWCE/H3hlqm9w2ips/goSXThHRFAcnv3vZwyQiNuAgQACCKye
uDc3OzTOS+xrhbF/iPiFAOsMQnN+nfeJSLPvoTw1il0E1RGlLAZeguudT/1xSR7o
NeUt8Q+JFou1r6RkVbhZoeOc05OYn3Yx/cuZqVsF8Kle4GF1e4BA6iSipKhPeMQ7
dhbh0MKQVhGSln33oyI3lhGEFnlhDRbkM+W0iMZGssE7QyLDCP/QpskhE0XHgSbU
rvFI8O0/oPJjiU0Bm/0OQ0iwd37RbPGB1NCVuibbmPY0Jsb1vM98Q3MGyuDnliYa
NImeRmenFLdHDh7OLdyajVjpPEhHdKg8QQ/Dnm+ZoJ6zAL6VYgcEWfRSd4SYoAa7
+Wq/tt19LKMUrAMKTZM9UoJspAnJrgqKwNu7FaPLnJVK3YhpvJBYz1RrFJcVAM3E
dD5SniSvGOmpOV8kHTyn5N7Z/jLkD6vrmCn2tNNR0AB0ZYAuONph+ysEdDWaw3Kq
ZXXKQ5FG5yvtHNfLvwTI+wm6klz2TSuvm+T+aQx553ZBYDrWERv/+g5f2dGyS4m3
LJilmWuINTqEIoqxX1stXrs2JDmqtuwj5INfZOP3xvD3mWDuNaC6GbpZ+Ai4vviv
sGVPsBG8x7e7GoojZUw/P0F3O/3zFBuSKZQtbV1+yJ+SJKmlx+UqpnsUIxoCECky
SDBHoTJgaD6+DriUrzg0SnBPRFV+9ia5FoQJ+KPgAo6t7zA9biM9grNkQKAEtDI2
OBDqXIuLEqYigRoTuTQEyEju+MT5f4XQ78KQHWy7tkiLYhmcXr1ZbPjt1cAjVr7Y
XuptgY6mKoZauezwMe7N/+AZM1X3+HY85y4zDhH+zA5kIz4954fJJCQHxrVtu4bM
WATBfhpPNM+eLAAQc3Y3jyqO3jMAju+Nsk+La2+ZO3OraKrWAuvA3GEpf1KRLNRU
t/Q99t2A6HEXoobuqJtwAPE3fxSWd0Soib0NQyIPx0a5lD9sh2IxRo69iqcfnHDm
M4yk5t5qI6mBExawf29ZCzJrky9F78H+rGMWsKBLQXKMIesHUk3OAaeGBEbF0pY/
Hcglt9OU+krEe7Ws2ZQLCowexByZpIQQDkStt2B+yak5PIMtY8m9KYjgtW6yaqHH
hWRRK7aU+9QfJ4aGSKNXIRQjh1gRZYBcEAGDjaMar7ySFxo0pzLz6ulR+FMNYihE
CodV2vutbvj/9omF5tv4ixaIQY8ZA7GWIDR/tlchCwtar2IdmgMq/EeFDak1Rkwn
W6V84dgvec8gj2LvVHVN2z1JZnZ7hf6UL8DMm3Dv/Nyt3VfX76f0lHbDDU8gN1FB
tMNieI5PuUsskFOVseZZ9iO/aGlXS1IUWv1/TnNguvePqSyonEDdYkJOWHBKd6o3
Ysy7I/3gXpWGWubqup6XRZnkwE+a6KaT1Nrhr8adPy8AfrsNS/xdZdg3qSVljsVK
8P1xp/MXYlxRUoX/B1zqZPsQ1aV1pH6W3k9+9bjrSr6GzRTVpWNmgV+drDkDmI+X
EOZ+m8KGMlqoVTkp4osmBIM+JWIe+C9v4PReF2pW5yT+IOdZ1y2Gz/l9fQx2Cpws
EOgztVZeFyVNLdJ374sWc285mlIr3s/DpFn86dwJGgmFFbVKNDrb107Of4Aqvtce
wPmLHzG3YQHbHtYw5DklKvjJIy91NCVnJma7Vcy9wEY6LfrTxWwRuTEOUVxK7Urq
kQYDgVVj1FZaiv+U4YBgBv03XXfdBzdoxww8dtWzmUOhbVeJvtWUMqRmORSu0en5
F7PkLoZvzZV8vOyO+MaYwi/csNfaqTmafKuLOSgdW5X0iSJRPot4W3XX/frwaYT8
18lcGpGN4vkVIsikMsVruEQPuplAIKFwEpzjVrGHnAEPklmsP2ixirp1tF4TZlUm
vMegQnmDEob5wW2Ekxuc8HKqqHRTVOoR0doBVyhyztn6GmgVxCvIqAtzqRuEq0Hl
TtDSr3XSidQaYSr6sfiC4p4brN0BF/UPoVhVefjgUBDfzHCF9fO0gABjglDyfzJH
MbpGPNLn5KQcE21YApKFPi17L/dW/aqmjW6qFIxMTDGT+sDzr0YeyIR/OnW0cFEU
GvbSCeL3iWJM+ERrdcYgBYdIrKMsmP2J324J+bLzbZ2UouxsTu7lmMR6nNdewVMQ
q7fK62yPPGaWpUUZu9sqA3jYLTJGxmsWdf2tavoxcApENWOjZy0IXotT8Asgzq6K
AOYsu1smQewHFSpexUjBWDhHJuB5taYpe6V7lAm9HHntJ2mzyo4yaDqSmc054gso
sLZSdyVAv45O36KkjvIubsfu8OCeXj7qFqgMtRfPI+lQWfhKHUvXHevDXdPLlhAU
fTs3cR2eDQgFFWDYvQeC81xBgvuYSAIMnTC3AlKVx9eJhT38zSanCcrTDyHK/Spd
OEvQHlw1fEOwnmM1X/1iAykIEy0ohXcTGTkseS8WfVIpXEjElBzNdGx4UfL9BWyL
9hg35Ex6i/jrDUu86RmBgYPy4/MMWpPDb/xd/KSZyjyr9GYCA7MjhYgjZdGIEs5D
LHE7587KaEJaNFWAybbzKxC2BcQQtWpqdFMDGqr55dejzEYXZibZQJbe7pQHeO1X
GzCoTkMfFIh5n6GD/q1d53NYvsP9hNX/+pCObD25Zge0fvzZLWKo7uAEIBJEeeLm
CvABABZ6Zuv5dCFUim4yKEaBSPL295WBlH63gnP++qTZGhwkG0p+63mHnZP/tK28
DjtIt1UN3jYYwwIvnxKW7q3qh7ouBCKyNo3bf+kozn7EtTXqMhFcL0xXwjW6kRf8
rqy2oJ7R+NVluTJ7n6LlxtGFNPGXf0UDRQUKyvOOty+6W3haxx2tU2a86Afw6x2h
SGXJXbrpWYVXkgPCwCgg77yo927g2VirQmQ0/TVRhr8oP+7ep959Vib1py+Cceet
HsAqyCi5rrB7tZt8nq9oi+ISJvWnlYjRp2bn+pTn/8tc2QOid2Wokdw+j218mZvq
qvMvIwgUAMqHdwpbHGIP6kfkOa6o73fajvjXIjTu/O0+fdzUCq2t9KoYtf4oKRfF
gLWm6AQjthXK4TOwlBIopZFSN/33XKhtPjAFZZhkL8kOE+B4s1jqhga9SEH0Clnv
cpbkPCuWIPE7z35WJtGNRVOkiarstVMwNsNQWdBJ4ey7cUdTvoOKSUlpqhiMM9br
UDGmi1zLPr5304uqO9ZUdEOLqT2S2hHIYDI41iuAEO7hf4C5tVEv3liG4+D89x4H
2/yADgxidqJUnwZbnhPAxzSH1Sq8LCgbl2rD/F+f60FbWt8wcizJYJcAulRcV1W1
1JCfvW5LL67udPNaEi+dm5CYpB0yEfZRaU/UD/yLroQtmroM2kTyR/9qrKaPWiya
jbffWivUL30Pntd0ho51aPegsqMLK2hCxRi8f3zNLuvRNtz0Bff9ufCRTA6zIzPs
5ZeRALdfMUe6Yv4Z6K0qWdCyCgjhjYaWAD+ataSYtAucF2li9Qs0AqP3oGwSF8FE
+kywKE2pD5/gE/hwXR0qyeGJz70vPM7v1q0QwGNOjuU8OZfEmPDqeLcFsWs2RJHF
rIK1OnaWcdr00aEjMQqAlmIoY6R1n8n/KPnSOv1qfL7YMPe+Y2mQFsZKOLqbcmcm
X/IzBOyelTzHC6/8xoqm3CrkFFbssibd80j/WcyutdMAUhixLblYpOHLrOpfnFBj
JCDfx8Zdn0Bc6p0aBpL6sI+SzVE6hO1X57MtEmh1NIjgOoR5KGTkpYtizrKQncpf
RjkcE0mpz5halOpf3khNQ+mto/Wm048594FqRigpehK19ftj+uGJY8ZWEZND+rkc
HjMEGt35sUkh3wIYt7NAxVwhv7G6e8rDnpbvToBjOpF/4/ByRbHnhJ5YZXlZbbSQ
ZWhezYVlPxUno2Mls7GkKBPGYOSSgMYUKootp3isBP081/zWDMjefG9EStHYlKTO
qwmUib0YvfMHbDhP2buiL/C3jKgfuqy9tIs12cpMt70JYwqDz/mXK9QAxNUDSR7P
C0PuxWNG7+0s5cMOuGpTojKOO0KD9tNTaRz0tVfLqutmUKLuaeovRxCOsUz4biRP
Y7hTmaPx8zM7Q//z6MWaJ2xH92PTYNyG21Asq19a0yJIcPkD8W4YvVMBTyjMy9x6
n0Zn36RCbKmKQ9W9MipGB8AdqjPKbRGAWVdAbHZr+b3U6eJmtUjH9OjnhcqofRj8
eMENztSbOUnL9mlrdVUUCwyMwPiYRyB/zBttZx4qO+sWGwVgOA2WSr4AA93NLbTP
zp50mc1K8rZZ39kkdLtiu5TMLa/0wVUpDmq/Nupov0YaAsnwrsEhscKSW/QEy/0s
FJ1vCbAEu5wmqvxQgfyrr8N+iJTbCWq8W5XN+DcoDHu2C8tEnR2FKd1OBOnDZTA0
UONscgP4NoiVnIJCIT0x4tdGu5ZA4Uf/zpGhRmoF+LwV8bZq541sSQ+RmOjsmHus
0J/VDVLVLDe42A8cpJ7PEQNb0FwR9shYjHVrQEk2xxZdFsWg3in4orA3RkBj+Duy
GNU26y7/ZIUmKj9LbAWZ6crHbUdl9LuJ9z0VDW1XKS/v8Zd841p8+QHdeiPWQDJU
xSGs4q71o7iDgO3WZ+Gc4S7oYAY30mp+dlqv4ARqAvHA/lRZaZHDeLPt6aE5ZwJ7
VWYY1pATUFI9WAo5hEpCTiNvg7/1QCl0KWAvEkiLXcog5ajFevLz5kErEBixg8a3
YCIsNoumsv79d1+Qy30KV0K83QLpnA9KkwtKP14Jiz3/6ePL67yQqnF6YQGAQbGd
B1s43Vm6CZfyo89KrH/mf1WudL1SII9t87T23Vqqg1ke/G49jwdtuo9MN13qxw/x
ogHWGmOY0t66U1RXZbjtdKY62m4uNbjtSNBPph+z2sAxuAgTDczNCMlyryVt1PRM
oXSgIGtb5RK+gvYzywkptRd4lfhFLUBbO7e+6NR7ZlUuOZ3ZTg/cwEQlJ7qhN2x7
gtxrn+PRjfEgA/S2TaKWFU7ML3CYAD+cadqUkpT1dWHWooCgAa9IYKJoG1oDscWv
aD2UCHKmdd0riEBcNaiH48vCIfqUWqriTdFpgKquPScRXRyM5D/jehkEnW1+9QkX
aOVii8eDiXOY1xw0xGQ/7OPl7UDWpO0WdX6/DCrrNvPhlD9JlMu1ts0BoexICMZV
pXV9DXx4YvNtB5lnEYF5SClQ4HyOrM0gQjYulWjuGPrslaE3LPOFlGWnbLj79Kg5
v5ELYJih51GkgJV12oopYzCg9Bdsb9DO5j5MlRwSP4OkZXCuc76EIkifoETlF2Q+
FG7dmHwEDw3F4wLvdFKRMWq0UWNwJA6lvJBwEpnS9TcuVy6NcdPkEON7cD8OrjEZ
fp2+tVdpHVaSd8gcjHgWTyNkTo3/AQLw8P8hjSAYW+q/nwjEluiBg3pF+k5ty3Sv
vsz67kMyG02iB1NLNMz4PYmT/ORxNe0ZTIcRTdSir2GlIAhV1FMDnI0tcceadZvT
jn+8KS0OVvwv6WtM2zcWL+R8QWVISONBhV5M5ksQ/bj36oNKdGs7M7MxqyhUpo8k
WAAa8iJXIRvCmDD4B1d1IEuG4biTFJ4wxLioprvUOyiMaZV9LbnelFpQKh2VM0bT
mzQhF8Dgp0dtq72CSeEj4XT2Xz/B18zI2RwrdTgqQu8FORFrNGvH1yEsGIyaVqeS
aMHvJ5JGMYtYXt5uE+1bzNmTAEQjC9r5Xizk6itOzaYXB2iDbY9wzQy9ElAcusUg
VR2tJP9Z5a8l//PsQkNZZNmxL1b55nWmE3PcOGVZeJ8sBUAR4HVEHyaOYliqns6W
Q7CnTitRrOOVsaFuDFuJcFum5TxM7+u5gsus23A1U5dmzOqklXzv7KTjP+0HwyFk
vBPhAMoi+0+dCzH2tElBo6lXa2v46CPtbqmvwOOTnDSZ5O0kA54ECp3jDmjTAayy
D/xGCImZ0mNLfcyQZGvh+6eVPuCPeWhpzqwX5xF8wh9z8uMuB5Qd7ZqAN877CxfK
MWu2cfq8qwnUnqutIj4Sw0guY/Jkx0t7TkEbTN0FVrt0I+/Er8ZCELbTHtiocGcc
nOFtYhhbpUpfSb2BMFu1nUdGCI5dAzx2JMC+bt04jmyqlH3gb2By2bMXMTG8hB/y
azj9PQIvurVS3qp4uF5dGIlxoRFRC+e151HAjF42PP+Jtq5uGwqW+uZLOVb2wj1O
qOWNZiQwy3vsDJEmMp3dx80XORjk2It2Cs/gUHmDzFAUFjFug0D1t9o60MPfD2Ah
793qSXKYJOoUbWEWg1IRh7rNpDJHM/cQGo6P3iZFkI8p705ZxyAur/O1UbiUYacF
1WyUxjT5LBiBm6O21QhKeGALxOFUllQ8k/n6fsEeKpAwbTpkYGl4WM0cyVSd3nQQ
9WYhurmWWI+OKBn7Mms6ABNgUG+/iXecPvpeDiMapZs+qT6UFN6jsyyuNmSn8KWH
HGoxDeA3dGcDLiYXgl2yykEypq1I7urwbDFfbmNNt0sjpvqS7/lEELKAWuaweNTx
W2GhMv4sV3YeBzKtzbuEMv4llCqZPojm9Sy1dijdRx+wsdmQ0O4AWOlfO1+XlBrQ
GCHyRUQE2n9ul9kwmwKc5JX5lceggAlm68mbAdPn3YFHvukNU9/nrHm0YtBylkfr
JbTnKJ2UEkXkgl1RLCJUpNEQEyN9KsH7fLXECUfkbQ0JeSAQut8mW+KmN+1a5UXA
RGxgf0Ub7oMV30UDdk7CoJEGXpE6hGlkR3XWjHnrGzyugQd0hIHhOtc10DtDZqgm
DUAZrraB6mLOKKw8ziH8jukSGg6UqnuI4ilP2j8lm09KJXHzY04xRTrLtiP8fBlt
bb+lPaUjdxITRAHgCetPWX405yiVzZEuMXhZBlMiazDSxliAtKmKNFeZoIr6EJM8
WZUda6XbGpzsdRiqCGw1SVttji7E3fPN9fRl1nLo1yaKrpIUSHACPUBEbvpa/3HV
4sn0hCbe9vQWghY5aYpPFMP2RqoT4n5y65K4TYyokjggTLN7ifiafLklw9xh2Ru2
hc0fF1dMGQRXj26OOVD68IJ+XuoM/X6c+Mmp/hXiXylqQAju8SHuY5nYJMNNKJtp
FzR+9qdS9Ll4c+7W+x/lNGAlq4MkWLHorgY/7vCjJXttxa1T2OLOfX5X6fE9q+lc
78zEUpSD8teEKxfCcWsC9lgrpxHMtzYE6GFYB2DJxac8qjXeR4IyoWtRk3BveXGQ
TaAg6fxqxIOJyBoLvM5NS6cTdOXYr+ri2NOMdYBUQFMWzAS0yHpuzggfj7JcouFx
m5yy2o+1v8k2K5w/itiS8W2SpvmCO1Py/JYSgf+Z0FJaXENTH5hnbCn79ak9rrDt
jXUjsKOfWJwhzjy1uQ8D1Ay7MHqgNrrdTItz5XCKVvYGhdfrvvs9OxB5vNDorHh2
MA0p0k/hC16i1OsY2OIQn/Z1UzV5SZ/tgMP1JjlIZ5xcNQ0mf1gDWDNkqT25nhQ3
cSSoxYbOWvjjeF7leI4AYtDFBfTzzVP4Hpa1e6gohkud+wz3pCmLGAyi5p7KmQYb
ACDsRqTokwgPzB/Pr7BV+DNG8WTEYGiuTwfBukct8/UbBh/g0b69pYAQ359zqMtv
qEBvydsOL5BNjLtv5Pw51Pl7AXrlqVdj5vZpXL8WilaYFDEXwHb/Taaxpk4ulTXK
JUS1xRCB1g8sLkpVzHe7/t2gDnQJ16g2uSxmh3YbZfJO/vvisGfYXTB+IVIph3vv
+nU0OmcKWqszmsn3YSUscE9AZ5dBvmFyzsDqUKiE4CMs0ueM3edGIGlYrrx5MSHk
wyXw97DYa1USgIhcJfIaYoC5DWOtruFqgOfM040rYCkUBuW3yt2kcYJlg7CKhXn4
6P/SoPTzW7YAvWi7B691987ZsC2IGpNsn/Sm94fyI6h1MU4gSNI9Ci7BiaC0QpvA
LRTrlzTGmttggYARO3Gqrfqdsz356azNtBw3Zq5KB+moKS7W1k0HB1KLGEEfjIgt
HK94RougqBD6MF/eG7j87WDUQHyK/WkJw964sovuZXcpcFynPaAj0mbBmjAYLXgA
lPidGwUg+nxkDv+avJ0+GzTaZIk91iHXLRD6XHj7IzHGuiXAPD1Bt4GYQwF/vs7N
YKCWV97G+5eAPfTm9FiHwfo8/ggxbya1wnKb7W/IMgCXOY1dId+Bzt8aZlfqXQtw
nY8Bem82Dy1MDhyjv3HXSbbAmA9lXAAXsk6/HY0Ld/6/BZ5v0075V0AsPalsihCj
Nq0M+xuDyOvfd+X9/ljE7z28uXFGCpWN62NcRLsxygvj2SptR1AzZjnRONG0xl/X
5bDrB8ZGyYA4dWVgozWx07hsRFtdjEpc3zClbUnuQQcMSvmaT8pyTwK+kqxxMesi
iXfzCpZtM2pwyId7aQ8CghOu7tE0CNRg/3WQfE1khBLhW7lRdTDqQ76Iz1N2iViN
hw0HzUWKgzZvD0kAdwQ9u3t2dq8LW3kczCgTawGdT0Bz5Sgtg2fHs6G5dL797JFK
NLWYL4SJjA1MnXdKlFVNfpu4irR041mtamG0zXID0masizsomnm4GBhNkkIr6vfk
z8XdCZNEp5oD6aRypSmi3pzI7cMMp6ATbGDk+HcakaxyprxurVAhmX5Sy3TOAHI5
WFulTkoa7+e617deD6YuUXwUfJcoFJulcvFdkWU7JNR5bZx0+lf5L/d/eo4RAzUD
dJRnZ9epaQ2fmnUU4dOe2qaR5robOxECBGd2hBOoEoPXFYZYNiY3l+XPCyEzz32H
FIipDDyUTCkzy41jUPf9MqdQRcFuByB0XgWPfJL6ciLwMkNQNKAc3WYv9AkgtUQb
qJwaqumA/3pAKr20lwJkNboulfhYxfhqVwXLwQNxL4WPwaTGg0nX/BsjiMpbeMrQ
KgpbucN/qpMW44QbglWov3UJPLRDtavzSMKdNzGWmRKrunpL/YlbOP2mK5zdP3WP
DxQAiwhIq51BsxT1nKmY7leLMSd70+F6A4EVEYjWEloZMOF87bxLzDShOf4FX9lc
v5Ig5HXtHaVVb3uEPN0YxdFrD7eaOGMzcWjwIRXH05qiWYy/cy0tpZmjqXbwDoK9
KzBqNV7EDZRbnFBxKvVILXjVZCswkM2UTYvHgD3zkW6WkAcGcQOi+iQ1nf6UGVOU
mnlibVLZs/WhcaZKNckMlKJzyavlYoMR4ErLRV9U7BseaEUi/IPYNBkkAofCZnyI
bi5SRtVr0VWTHxsvrhul2E+JWtyMfD/KUex+rQ+H56FwBjQM4Y6v8H1aB1iLSRZ1
Jt5ht55yTCK4aIanUwWoWM8QUCcTD8SuykXJF1I63yXtiN/SFseVQLThLJ7+b4m+
vIfi10BzkV8mDpvAwF1Wwb6L1lefw6Nb6OSnn3FO73OHFMG+V4K58m26UrfZ/K3n
YuuU9FO8nhhZXQt+m3fEqrIgOYMVY2lgmET+LOpefyafzd14t5s0nCZmKDcz2CIm
QWvBXv5nKN7rhkL3ik5FZ8BkDLfO86JBedR4Cqht1eyf//KCgvmif2b4+g3F9pjF
l5/pHdK1TufP0nTJst9D9oB2C9SEU0OGAewqi+cpuHA=
`protect END_PROTECTED
