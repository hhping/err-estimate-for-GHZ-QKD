`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRb77Xj/W2kHBqYJPOIzfw30uzoTEUPfWBqvfFJBppnFgJZjexDQORtiuEMm/RsH
gLXp2dHV+4uNggGhL1IQY6B7SgMI3vETy3X17uQgwrUEzHndXTErTutVO6YbWvCI
0/lJp7E8t/3Cw7yRkGT3cU0bb4pupP1ELPiX3CJM4RAzd0gWYn/wblkuH5rktMMq
ryXyxxrXgRyOIr48zTjgyZydBuuzoSHP5csp+7I8sl7Skc88KyDQeF4eE4lDcqyv
qwuT3V6Jtehim8m0EJ0oxR4xCKSlouh55XkRZ1YXUkdnab7h/u8CbpIUoERWXe7H
aI12PLosuw/VIX5wMAkYJJ0wcqGrjLizjgrgso+1CQYfWv6KEF+7ma72/AKxmjZt
Tq4IKYM+x2sssjwhS+SgCWQl98jyl9bv3kfGwe2SROfd0i2EF7FMtsQN5tAiU7tw
hH7kukSdsXR93TkZ7/ElsXFqM0G91DBf3tdS0Hmg1NOUsRTHcwizw8v8/i+5dJBX
N1qDdWACTjKcSOoGLhC83Ay96B88+2vCyZSuA1aIxIJpTvmUqdhTPXe3CnSsvyLh
9qGOjeKAsLytwUvRq5kJ7ZLVZ1w4rRfV6yP/4aV3Vw+udPcG+vTg9rpXdgliLVKD
kcBDXKEXMDGBSQTjtFgCEDoSkxUrHRGgjuwNoiPOzdYKEk14oHTQYbmoR3tmmeE2
3gCIXBz3bi+ndaX1ZiCaWv40NZ6cm90WM8mgk+7djMx6ct3ubpiZ4OKrNJadlRJX
ZYyKJ1XTJOUmtN3PxiCQwy2OW1sHy8p5Xb4+Ne6brecfY9ZZ5lgRVENqHVK+TSs/
WeC+XvmebmtfpoX6ICk74ECnC8Isql4WxlF4jIlXWL/11gQ/rjnuKcOfAxZS/u5y
vlzMVz68rdNbOU4orUT9+ULjVun9xABeiwioT+OPU1hm7CO431saWTsNWUjOCqZA
Vt9a7X0ScDCRa30eFkpjPH1r/qooQzoa9obTYPtUV2wKmOxBCGznKyCUD8/zzRnl
7DwgKGeT6625df+KMacM8qgc0M1FErKvl0D3kmSbW1EeSzrSXsuJr0vf7dA1keMR
6aC7sVCzPQqbV1sIW0S2J/E0NDpQq82+WZCJETTbU3MMnDQpmAAWf5Fv3a3lz19i
QJh9EfO2UmwizEHDQ2BHdpSbLFjdFvjJ8u8wVmjwfW8ldHSnMmMwcGVdhAujhyR7
hlRFcGi8WQfj0S1FezDOzKcySHwHyd+PALEJ51TPbo6ZeARms26knn+V3j297Zny
/KHQe1L1k8hnYK9JK0tT1pKQiTNxI73er1dpb/RkuR61ZZw3kGjGPrOCBZkoqJSn
rhDmIgWpIMs4naCeVwpazJoHtEyepLnR5SBjzPKs/cQNJFS623uGTZXdliaQIoY/
V43gbMDR/SBnr7yzT0tswGC0q1fUoWJzkwmcVMg/FL4cSDXnlnYoVGCTXPe++P7n
mkpcVMR0g+xJAay4cY96qsB07iPT3I3kuKk1QUdiaUlb1y4ZKeqBXOfnMYVHy5fg
Xkex7j1QxyytYYV0zIXPpJyQkipZhb2yu42QJnqa1hD4BDydZlYj7pDAdkYKzriq
hwz3qMy3zCAc1fBRfUiGnqu9fihXiJvZwknc9PUpESSsDdajiYfVjc3NbazfC0xQ
JmgjJQvrLQMEIHOiXeEDobuM0RGuj3dwoioNKbuR4HCSmmsSB/SShlqYcd7ICX8Q
04wl95xKjkjLFGsB4afQG2ECEdUt94hY7KESjc7coTcnC9lIDz1Q9Ea9w7ceAX37
O2QY9af5hNzan691NwK9UPvugS5Wbz6NdEGdGwIycjQ0H3qTQGD2XDxZQWdrWyY7
F9POlx6xKHJnQVQwg3+lPQaGhZvZFEMekm7fUY0FCN1iy0kKOs32z2Dpt0eAIRz3
Ay83VuoxAtfOizK/44bxj8LC4mIfYo2sB3UCR9qCs9CgtYkZ/rT0Tfp6unOQLC9z
oH059PSftas16r5x35exdw==
`protect END_PROTECTED
