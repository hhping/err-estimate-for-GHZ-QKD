`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fz4zxNNqKntDGXo2pUjTpP5OMSkMMZ2XSgA7THS3DSMmB2d9bqStpDe5v02SSmCl
6nXLlUDNfyFpd7Nps8nqo+t7P891XzDCcDUpPvLGfmY7ZcZP2tsL4af74ugENB/n
bYcfJqOlOFrcTwq9wsC7SFfLZo6acbGwBbIAeiTscNE266rtMD1VaVQ1jnQFUtEk
q7zd7gI12oqeV7WNk3Z7HXwayfmhyiFxbZxewq7k8z8X41VDfX1pk9quHiUep9gW
nEPT/fsI1R9QvnxwBGIDHm6rhaj1kCVmvOp/AO8Uo5tt9iNKKu5VK/KXRwvdYaoP
MENd8VSiiRLw76m8z2oY2iar/SCc6xSvqZY5zluvGUB5Mp8AFWEQJkbaGEix8xtl
vdFsyHRz1K3cFX41jilCkjoMDu99yl2THGE8CRQWNGDJOaEApQvWZFgaZeKPRryy
G0n8lXixSnyvtDilSs/Nd1QEp7txcAjC9OmQNJFf+ZP9zUE8to5NY3deXnw0y5as
JEty31QktDMNHT/tUpXGlZPLOYk/WxBChXI7A8WT+Ag=
`protect END_PROTECTED
