`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifcb5dLzCwY1vT98EC2EVx1deC9Writ10yxuwoHU/MWPg5j+2YnhruSboBT4xprq
VHPh5zhA5/ky6NvUtuoII4zbOWgGs0r9nEjS0Nfvu4+HRgLjiNCD5gfauzcNbIrY
GKRkGmlaMkVmOcFe8fJaz40AqOoaNzmnt51J9cl+U4QujMBNlFm6r13x8sVoXf2y
4fWoMSKPVkIj3Oj6y2mObWGSASUk1vmuQFm0kocNIh9ECV4N5P1+70qm4egfOGQB
xMPaQ+RN2jyVurJHpE+BRvhbULjxhE7f3aXg2NxmA0a/iLCHQYNocxBgcxwOAYH0
SMMeIqI6iDhKI4OlOXMR1cIPI5m8EtH9Dv6PFNcwTRnpBB8saaP3ic5F37VQyd2/
6evQhlFziKzaSYxgq8gFIVFp6o2NSk4HnRsm8qTIHRVcMl6rKz0yBVJjOK6sLyVu
JVGh7knhdxtrb4KP4eHEnaCHwEIiIhOs+pkeJOYhK+9o+04bKIlYZOTByqiqLEaG
9Q57OsdFB1WPGuZNh8DlutPGXGx4qLys+1Jr7PyEE8nKLLH5AW9RdB7NtxZdLJTU
pDT5zZKSZlrrjKgk1vuU8b41kNyvdZQLU9fj2n7yQc/80KZQKRs8hgibpfiOiTBw
ZK7gsW0xTkQHqwvjG/EOe9j7Q+Gb1NXcIs+1co0/i/WNa7NHzWWMUmoJQ3lU1Bgi
HVWn3eEHwjUu4JMtAX3Av8RLdQkwlIO+/wCUfSBfrzMaDWsFpWfUu2cwGtyLouSI
s7IQro07HsUOeY/SBxVTQ8r3iiabkbcjBFiqGbz9Mk6+lfZcZAELGnMstYFc5MKE
oOTJFmwQfcA2Xv7GVJsJA/aP0EHjdqsrruUqi/GekVnbxJ1zL8r0iExYunPoduSr
i7oy7B4gAJDfl4WettqeT3V8aCiTBmpo/jGUBTbKehW3+qyYheDvubc021rWthG4
rSAMFYr0QDYv3Xp8DHt8rS39+5QBH4qditWSjA7DtRuW+onDIiCk9XQ+H3gpeHxA
I9jnDAJwlvcb75cMR6yz0OXT/eSyBlrMzyGzAJaW9RxczUZwfTIYuaqcxUYmFJDI
FezJJ6OCO8+TQKCfzXQRTzrHYmF6debO1eBjaTlGAYyd7I5kkXHuUNgVlbyQF5IP
0FnTfudLM/88hzMGuGX2adPH6VlhHMdTxqNIXrtBF654AG1mYlYqlFwjSmCoGgTI
ixq6WCJUlLk393ru9Vo77hfTyl3AQ1+gSV6CL1Uh2fC3RBUmjsRgzFeO4p8I5piu
7lo2c/CxrsQdHd5+La8iXH0xde9/iHVcr1TvcB9bMoyBcAZAt62o5lVlE3M63tDX
DB7u07e/x7VVKg6bNOlxZ0Qd/NJe5SPBQQCRfEecNHFD88z/mnj4bCLbd86F0uV/
4APqBUOkZjx6oKhfNNT7teFmWkWzj/+eDjv9muXLWCA0fLsZgg3ltB8W1UdGEGhK
UBjccP/UaWGvmO9Gjw1sGvBe+0k584femHFw2kuwYsTbo2jtneUvJ/SMk3jeKqa9
laZ7iI1KpCP5BwANIDKrHr2V5B+HxhyNflqsPpScK3yIL9nep3Qxkmak93PJ8Etp
iK0xnz5jE4ap0lGGQvSJgWNFPVZe98QEfiyFyau36QqZ1TRuKEgCD4EtDWphgekT
c0bbFk0vqXt2wuifvYFQc0IazWrFAy6qKbRDXlhbkhTLyfKlE9vei6eUytkxFg4d
Ph1QBUjjzwETm3eWiXkvRxBvJuko2UEmZjeq/gtGmqa8k3Jo6KqJyj2sTGrL0CZA
QzyJlrOl5wiwrM3WyRSFzPGdArCT1kU7RDWzYvPLJVWJHF0fi5IVTdAfrnM1b/7k
OdwDx3OFxJMKvL2aYqW9CGUUUEboG91Nd+p921D6a4YNQ4ipmKgTNbcgR0TCw9yr
O8nfF/l7p5m32v4ykLzbLutnqE+akZlsLTgk2LixYzJvxgY54LX44qrGycCmEZaL
dbDR5mTLduC+Stkk6i4nXMzaia/rNVpkyH2mAspdolKSUDLX1b4fcqJWVMCylos5
3WmloVc5Mnda1fkYzapUHtoafy0jAQP+BiTTwLOM6knzqRzmbKlrAG2FCXXZvJjd
HUTj7MtxiC8IP7/Ul94xg5HtMfBtMfQEBbaOa4LohomcoO9XImcGAJ1nSP0xUDYY
CeT54nqs9fFP4qdvcEiCJttiYRYv9VxyCaK/cCGB8nfKc6tNTjrSPRuI9Fv80IRG
YsCq371wzeg9mC1zVDlFh9fVfkVvvEQ4oZwEkMXKYhpfRjSZ4kZlUEhC60FPUDkV
IuuSDrvTa0RalvNSgBrkSbpvN50FtQCZXLb3vgtkq32aqZ1bXFr8v4HI2gngZKw0
AvWs3PHs7+IpAVjsAtTJzPFggNcO42Q8aDSvRAPOhU3GUkUj3UO8Cia337o6VIMg
MqC9TD2NS3D2ZXhKtl/bOXWZxlWG2WRPBzX+QTZbeEsJvE9CVNirW2uVdr6yI2og
0u9Jf+wJYydPGtvfw1kVeb2tATL7Ku6V0/dRbaaVJJ8=
`protect END_PROTECTED
