`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25lIPPjXuHjmiuuoQylAB6ZpwxWYszWvTN2d2dTqnzLmUk2L3VZigUyz1x4Q37fZ
noD0lUSr6MU/9WJAtus/08tkMxeecnWZ/8ikzaS+uf7t1YJvOPhexFaItOU2Z/mx
b/kLqu+otokfxDaovayBonJnshJ264WYvUdY+efij3eOBEwG0S5wMf2cxnm51e5b
MLMgDXpiAnqiPEGTnv/7wphQjQItLRC7y1sNUWlEb+TXqsLI5SM2qsCpwltUH3rc
mO1LWsYeV4VUJgOzhF6Wr/rA2mjOVrx9B+zoaaZSkLnuFLaIexsPOVWNeW7cA0pa
JgUgCknUPuz75s9F/zcDDi4HAuS1BV6FNBPuwwGmo7gxLvVtV7x7BMxV8n/O7MnM
8ATjHZFSqV1MXRXPfbiRldvqEPmMEQ9LpeDp51usGQUdeptSdJCWbb9cFEcsxrna
4/yedApc8t+Vltit2JSRcQBekFB3434tnRnm5qrNscr7xMgUVV22GxYBI+F2kwqa
Bn0ZSZ9Lx0o7zAm85Ps+W8TjXnIbKmIs6IJH+bxZnafDJzxVhewkLNtfaEPC0+fP
32fnq1QAO5e8t2b7JQc5aRohIKGA6JZ5ThS9b7pkEj+sFgD25HS4Ge9sx1VXTZyo
UrD7D6Xwpp9Deloe3ra6WHyzljuKgrzIeGBBSZyd9K29QXk5hh8Uu3xOi9vXEH9h
10ZUrfmX7doUQYmTpJeHdl6+r4N04chP/PVxSe+Z925nGlL4tBelCeNCWtX2U9NW
U2tMf86/b84ITtd1zcs/KH+5E1hxIE+0571wC4wqkKui+4ArVEmGGuGIhI0g+koQ
ZwYpnDVB5JFylyBPfe8VlTcud/tfFt4n66Nj+M7/ptxZrK4+YTjdPA4SbrFTc1r/
WnSsLHUi3g6Q/f4X16G0nYYIloWRKiw8Gai4CM6JCdMHuSRzHopzsAyAzJdaqjPJ
ZDqcAFjrIisRzsSsUgBNJnSHddH5flKQe/wIb2CYWjBlYsfGuOkTmQhEcKk3o9dE
rsjV+1dO8rrqCrAJoR369dwUGYC9MGM/UyfuBZAMQjGbAYsGR+LHpHWXfZOZ1gfq
J3QK2oochD/iywLi6llpcfaaTL6HbBV96P0R0C5afefC1x+SCNAhzgtkejA3joAy
CHw4VZiYz9xmgsx7HM2EMRwxVJ78zpzLvu4eU5me7839VFJa8YZcmIXlG8gTyNEW
+JLkuNF1nirqEStegqlMbZ/CZyH5H6+WNNNB+fZmPLhVy6WiPAb3KZRaQKLAkDnh
`protect END_PROTECTED
