`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBO3cY3vnv73xdoRnopOFv1B/4DX2N2tYus/3dnSl8l5j1tz63wN9maLvASi3gts
tCUwZ5oEMZC5qNrPAWRCnQEO0jxAgnVm99l5FlW1BtuneKzTnPCcGEOKVR6JQvL+
pSk65fIJFGhqubpoK1Ns7L0ClPmydOjdJcpSOENAGA+hIHxKFtoPbmywemmvDngy
aqbsI3jg0rFtsL6Q8M3v5q+1gDrtCRO/dHSkFjAce1XUUu/LFCJDzWOLBNnUWo8x
MouBDfg9pO4xP3w0V7Gk78rRNCHNIYIC5gIFcZw5TxwjyspQSuJ5nsbgwDt18clF
zqkhfCD7SsNqHVvyUpFBtHf6Kl0G1Fdu8dfNkK8vdPdVv4m2QTVZbkcSyKhDtjsy
Zf/lmEtAri/CGJhQMiI8Yt9gHKDclEKTE8/3AhVVrFCSpUKtdxCWf2paobkL/9aM
+McRKmvlV4TMqsuDtnKHxNL4EqCz4lPzXiyEOaTopJ1+EXRDvvlSFv8yzwH4ncXI
iLPBn50nQNbm10S3IljYNmFP2shocUBslY+L5pTOdOKNWMRuKx3Q/bVCF/T0i6wV
cstrPFF3HgDwQ4Yg2+nNc638u9JT5h8P7brQRlBEGt8X3R0TRZQrqYJHsvgLts8g
fzOjqdZkOamfGDH8pb7+d0mfLr28+zRNsG1nQSf1rQWElKWtSyUW7p+KY+eYwy0q
ZC+azq5+i7iM7J2JTenvpMN5HMXugdqqNpHBexHF7lT7Yaw/rMuk20UrKjNshRCT
c41domTfqNIm9IUyZg5+rQy0bq96r2gCPsgQpDK+1ObPvjKCIFqgvy1Q2VtCX89j
dJpRxkXBIiilnNh0zC3wV4lr9lzbDEx09NHi0QgPZ0cQMnXdpfEp/JZZdQJdDW5m
54nlpsDIm/H0xw88BxFsfF3HvQbNL6s2Nmq23B+tw4CI3ss7jcwD994+BLAATD15
QwalkX71myxdyxO/SDDzjrdl6lQl0/+umtMWqyCC0aIz4WfKm9MZATb95nCTGlD/
eUrtxNFCOAbyk0Xii3JZkRgI3T4fIPQy+so1foBMVfLIa2SwXXGYqG0rnjddpPzZ
xZDLyj9buO6oa2bGmnyXXiypvdqGXWyXyNCv62OSDBjZLwgGmNnfTke7fqRgcvjH
vpo28dmtrD/83Ow+ezNPKG/EJLn33VGg7jiMXBMMWbeWGk89c2dptTC5cIHz0Zel
WFdfGGMMlpNlCcHTCfDUAdGvC07AfWQWLzOeKGs1dUIeK8moHvX3JwhUs9nc3XDg
yOMo0vPSk5pjyyRKSWg+KFbTsF2AoR4H/Iav5TEgQfkhbEWysyFJJlwPzyCgJY3G
ptoecZwKo5aSeV8Chbu067KKIK2okZoJG+fX8Fe3qNF3ntVt86kYnQyqccW25JcV
YyWj6TTozqka9PlHRM2lEZnHulzt/Sl6ieVvij4Jg7T2GlhnucCNVnNxv+hv3aMv
y8rTPz26VJTNNh+gxPwW7vrwO1hSxpSlbhRPSgfWIPLJs5eIX4jIsoPsvBJ5nXJw
tCrLA9N6C0963n9IU4pvpA==
`protect END_PROTECTED
