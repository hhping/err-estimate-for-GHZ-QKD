`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfyMgZGBZFGIo6jFM9+PbwkED2XuOl0/NYcr2JvzImIFg5QBlqzeaEPIsOE66rn1
Tbc9Tn6/gLZb03LEip0Ea2EXZHYRg4yM/HWyK++IdfQDCbz6Y0I4WLk6cpHDMZ8E
0wcEms9IDzzIQI5qrTsO+Y6vjiFGoC+Qbdtc44lrw44Bhr7ISggAZytAT+34L04T
tz1gWJxeTRg0cGLoGaiSagnR/chK+HUZFMrBTSJUKXZHCdDchCs3Agyrg8s1TM6l
yZuAZMWOnIqG3igw5MXTSCuRHk7q8hoJqM3rS7GaeMk4yxp2hGOPqAWRWin6SlmN
4ZeJx0CIls6s6Idz+mogBX/Xbv5BE7pdKi2mpQniq3k=
`protect END_PROTECTED
