library verilog;
use verilog.vl_types.all;
entity twentynm_refclk_input is
    generic(
        pllin_msel      : string  := "refclk0_ftop";
        refclk0in_msel  : string  := "refclk1_0";
        refclk1in_msel  : string  := "refclk2_1";
        refclk2in_msel  : string  := "high_2";
        refclk3in_msel  : string  := "high_3";
        refclk1_muxin_en: string  := "disable_muxin_1";
        refclk2_muxin_en: string  := "disable_muxin_2";
        refclk3_muxin_en: string  := "disable_muxin_3";
        refclk1_tp_upen : string  := "disable_tp_up_1";
        refclk1_tp_dwnen: string  := "disable_tp_dn_1";
        refclk1_btm_upen: string  := "disable_bt_up_1";
        refclk1_btm_dwnen: string  := "disable_bt_dn_1";
        refclk2_tp_upen : string  := "disable_tp_up_2";
        refclk2_tp_dwnen: string  := "disable_tp_dn_2";
        refclk2_btm_upen: string  := "disable_bt_up_2";
        refclk2_btm_dwnen: string  := "disable_bt_dn_2";
        refclk3_tp_upen : string  := "disable_tp_up_3";
        refclk3_tp_dwnen: string  := "disable_tp_dn_3";
        refclk3_btm_upen: string  := "disable_bt_up_3";
        refclk3_btm_dwnen: string  := "disable_bt_dn_3";
        ref2to3_en      : string  := "disable_2to3";
        ref3to2_en      : string  := "disable_3to2";
        clkpin_select   : string  := "select_clkpin_0";
        refclk_2_up_n   : string  := "no_weak_pullup_2";
        refclk_3_up_n   : string  := "no_weak_pullup_3";
        tnum            : string  := "tnum_1";
        location        : string  := "location_1";
        refclk1_dwn     : string  := "tri1";
        refclk2_dwn     : string  := "tri2";
        refclk3_dwn     : string  := "tri3";
        silicon_rev     : string  := "20nm5es"
    );
    port(
        ref_clk_in      : in     vl_logic;
        pll_cascade_in  : in     vl_logic;
        up_in           : in     vl_logic_vector(3 downto 0);
        down_in         : in     vl_logic_vector(3 downto 0);
        up_out          : out    vl_logic_vector(3 downto 0);
        down_out        : out    vl_logic_vector(3 downto 0);
        clk_out         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of pllin_msel : constant is 1;
    attribute mti_svvh_generic_type of refclk0in_msel : constant is 1;
    attribute mti_svvh_generic_type of refclk1in_msel : constant is 1;
    attribute mti_svvh_generic_type of refclk2in_msel : constant is 1;
    attribute mti_svvh_generic_type of refclk3in_msel : constant is 1;
    attribute mti_svvh_generic_type of refclk1_muxin_en : constant is 1;
    attribute mti_svvh_generic_type of refclk2_muxin_en : constant is 1;
    attribute mti_svvh_generic_type of refclk3_muxin_en : constant is 1;
    attribute mti_svvh_generic_type of refclk1_tp_upen : constant is 1;
    attribute mti_svvh_generic_type of refclk1_tp_dwnen : constant is 1;
    attribute mti_svvh_generic_type of refclk1_btm_upen : constant is 1;
    attribute mti_svvh_generic_type of refclk1_btm_dwnen : constant is 1;
    attribute mti_svvh_generic_type of refclk2_tp_upen : constant is 1;
    attribute mti_svvh_generic_type of refclk2_tp_dwnen : constant is 1;
    attribute mti_svvh_generic_type of refclk2_btm_upen : constant is 1;
    attribute mti_svvh_generic_type of refclk2_btm_dwnen : constant is 1;
    attribute mti_svvh_generic_type of refclk3_tp_upen : constant is 1;
    attribute mti_svvh_generic_type of refclk3_tp_dwnen : constant is 1;
    attribute mti_svvh_generic_type of refclk3_btm_upen : constant is 1;
    attribute mti_svvh_generic_type of refclk3_btm_dwnen : constant is 1;
    attribute mti_svvh_generic_type of ref2to3_en : constant is 1;
    attribute mti_svvh_generic_type of ref3to2_en : constant is 1;
    attribute mti_svvh_generic_type of clkpin_select : constant is 1;
    attribute mti_svvh_generic_type of refclk_2_up_n : constant is 1;
    attribute mti_svvh_generic_type of refclk_3_up_n : constant is 1;
    attribute mti_svvh_generic_type of tnum : constant is 1;
    attribute mti_svvh_generic_type of location : constant is 1;
    attribute mti_svvh_generic_type of refclk1_dwn : constant is 1;
    attribute mti_svvh_generic_type of refclk2_dwn : constant is 1;
    attribute mti_svvh_generic_type of refclk3_dwn : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
end twentynm_refclk_input;
