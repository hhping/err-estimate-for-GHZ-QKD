`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7LQAfBNwn+7jtfP1sTAGctHFPh4RsSbflv+1jz7wTS6R9YSIQ/TvFgWzEe3b+NY
sf/yccPhhKTGl0kDcUqy9F7oFarWVryu397uFNeFuKAadgsDPZ7CJtiqv4fERwhG
CAuq7qVgrrPkNLXnOjgdqVk4YjUbLjyjRFwHqE9dj0qD1GGLDHZN2po6seHbYz6L
jEoJ5g3n8eW8IzVKvF21sHsCI/ronENO/C0eG7v5UXdsNy+4QvXq7Kv+1bZ/KBSr
g2JbQk3w6sguxytaUZA5H7RP5kDn3KvODSaYPXaSPSE0r+xQmHGL4g0Soh3V8iGk
xzKsiwL+eBrgPEuMncu9ml4ta7HTZFCHKPW1TZ3PIEsgc+CGJuPKWUbVfi1sxqdD
oc7Z79346rrRDjdRQW0prVhthMze/JTPogy0qoMoYvZBwdxzIbTQh5IKZEQKD5Pj
V6PL7y+PcuufyMcINkwMtZDz86vsSEdfjUV0bIF9r2H36VOaV2oqhYebALPz10cq
8qHG3sLHPTYQj+Oe1Msa0UOA5q4ZFEeCZjUQgHp3bZbJyrcfigLIeDV57ojeSuIA
`protect END_PROTECTED
