`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyGctDKPZh4Pw5guv48p6Ahj0zyi0iMvhOJuuMPCLvqtjmAQZnhzK2iUVA455uAM
LR/NPd6IOhxMYx/XSFivMa218eeM/MVZSU+2vc5Z2OQ57Je9oxuy5LWDIrOdB3Zh
lR5NyzaYlLBBjBQ5knH2PE84qmtnyWExLF8vjK96xVKyQIuL+45z6MgaRiPpYewg
jerQxkPfHAjtAeam+xRf8q3X9Q0quDd97MOfiOVgUhIyw0B3I7sh1O+mXLIuEBkr
iDg0TA66VBzQXvvDbrPI92sOeLUb0nMJDZzb1/3RT9s=
`protect END_PROTECTED
