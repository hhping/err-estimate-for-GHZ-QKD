`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdbEfizxBfo5MDf9yQEen8P+f2NUfqNFoVcM7GeSh57ORWLhQWwO/j7y1q0/5XGw
BX1dlXv3y9l8Jz+ezBVQpe5WVRqUtnqpjEaHDJQyGA8/xBvsNs9jcO7/6xF2VDVb
VmqHZP2wi27uKMs+Exnhwl7Qnt9zOMowz7SJjuukQ/D6lqufISo7y92N0DE3bCwb
qEmfivHTs1VXPwCe5c4GAdJXR9v2Y2QGFmLRJYhcUF2NzaolGJfh0Li0A8KP9nL4
4CPNOMlGAKlwflWYS0Hu9n3LOcp0qZMq2gzL/WTt26xsLkn9VuzNUHsjt63eU7hc
xnpoqRuOYMA67Qjq4G8PqoLrcSNiA04kner99vfZkJznd26LkimQ+65LmwyAAeRn
y1ym2UGIDLf4YY2xJ+ZcGWilDIqUGqDgidFqPwKrZHSjzcngPqYmEdzpqJkMyxtP
m8gVZZ7MT3C0XsTYxPYl4WdnT61i+ySvDVaLhTR9XIwKyVhYUWh00+qGDouxQha3
/jUFZqnZIYzIT4Fe+j7u8WE5NUg79gB0t5vvqNU4i6Ljj5bTyijRtIYmJBtA0p8i
D3spxyKTQx5xNLAdYb3NnXsUOOBhe9TfuqxlZsmaHtlLpDBf5dt32+RqVi8QbK0o
bE3xpL1YfVdicqCYBLkBtYybQMxX/i0a1KBftkybQBboLR0OEZH/9lCwPD/cJebu
fq3lCL19DTDMJ7NrMXiAZsZ7w3V42Rzug+OA6ktibqEknd2uPi6EKvz3enmLgXmQ
/Bgl2xMWbrEhZHGXaQvcOsKG7mkZUZYelD/iMT3itaQ=
`protect END_PROTECTED
