`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JWyeo7ynkEFX564DiWoxT+GRU0M5+GCsQ9fB8AYxon8zVU7N20XJQIPnybIRH/jP
PMGu3vgFOlzsStyc10zHcGs4OIhvCsUVPpDmqT7TLlagu24xaXgQpgry5EFSKnMT
E0ecG8iBaMjaNPWApALauXsOvrPaQvkS53WyLjUhqHkOEr6qbaoHWyLJgBi3zN6W
JC3ArOpMxYZVtH84ZsUV1Ar/Yr+ghhRrywXAEMPu+OidSsBAhgu93CqncJPhaR4+
tL9za5NAzuFAyIIUw0LpsXshpzx15TnPRTT55jMfJmTmcfQkYVBffVuQbE3KKc8G
35WXQDpeRpHcPJbXCHg4FrkUTJ6msE7bSTK4in2O3fy3jOpazL8QKEF3u+5P8hfM
lwsMLJ0Ls2AVbA42mOT0OkTyPzNFBEEhB9h0a0vzz1COVlWwjVeas/LhAoBCoRs8
prjkiBfX2htvkoFFSOrXLlf2pgKjC8COzc+iAddILeGYnKiCSB+i2uRDXKtRNub8
02Q/s7GTt94Wpb1eQld57APqM2hFswDLq3IiLfsNXnLckpjmX3Bes0NSxevW7nMe
JRz//mzHMX5BXnDgaQ4d5Z7yby5G8mhht4o+CNibLl4x2399VvEGl64kruck2JQU
fa5EjL0NSoYNyeG5pln54REqrEOzJaJO4OIhV05jXX4BPS+LYhLWao3Xm600Z541
sI6/HOjpo8Qspqp8mQMFVX01zM+PWhIb6zA+XXDBioVWtux0QlPw2AI4zzrtQpDC
FEjNoFMfztvBbIEE2kVoAdAygiWSmXGtX9aGguBcXpba8qVJW4f2n8pSm7EluE1r
vuZjJ4oQIvzRCrQ0yMY/GSonI8fEg9k+C4nGdKpnxApNtYbUxE3ZCzyCWShq+bfi
NWk9KvuHo+IdShN3Pxbwhd2LdNBmgKQQ8hnTahaB9sl//O7G8otZewHCZqkfG9r0
A7xCvh1rue2PnPpsTzli+KNzpWW7djbR9C8xpqHXxnxu4+pgAUokjDnbR+OSCOgF
dYDckNC8HYzKBKnnNyHD1k9+FXfMp0vixBJyylFOFN6xbN5O1PaQnI6sCiv8MTRc
ztah4QCS+q5QxupSNLgv2VkqCpTLdIutPFs7rMPYufZXcKNoHjM+epy/HhwN9r3p
zFTmxb06HorpKje9H45CYQAL6HpVeClsekjk5RGnWz9E/XOmiiBc9jcGi9M+tdws
oqQwtIBinYDzbrzhzE/hsiFuZUOf2AdDF9mz3P8FDBprsGorH/jDnYO54Q0pq89M
Kt1felxCM6adoKw0TtXZPXjH9oSTIudIDLd8XPo9GS2nb+r0f8OEkbs3RYMbjUQs
b0EWIBVQEf0sYug5NhWVHCy3oXFG4x/ZVNPdCNbGtti+8KqvoFJ/+c382GDl0J3H
IBOB7TdWYAHCvusvoZ46Q8RCp9vOIo5nRG2+3NM50T4FmoWlP0W8lhetDcr3TuB0
agHOIvlSPmgA2SRaWVezk9JCXsdn8JQOtTZpgknFwYgNUXgtFK4rP/58uwGjN9IF
fINVchu12xa7v063JBcZQAILb0fbnYztkRhStIUzMeOzhp909SNpkaXPZLm6Vret
Rpl+9ZqGj++nSyf6vb+RIkH1YGEQ/2HsBp+7alUj04v5b0bqP7gapMCGEW/LAoYF
N8Z/bYj6tWFOAETCuW4pN1qRJFuID1HM7dQCv5vPI5EgLwzUhCVSdxFSzYqLAIPg
d7zZ+GVN0wnlSWyB6UdnLGEAISaGSkvNRrekknEVjezB+34V5EehIzhVqAvMWmvG
F/DKK011hv1pKojoevTz/p6IAMnwlOP1vPtbkkBnlXwqkVxycvMGv1jhkCuZDaPk
6s6UMCpsErHpnpN7iMZwHkUzWxfrIpQi8JUmrtfKTznLrmw7ZUSF5iC/+cTc/hxq
MnJa6f6mDY+E1UuMhY4YlAOt05tlFCJWqmBnhBP8tfqsS3oPEevpnttRGATkjNJG
+gOpCIjvV/oazkJOwwLDUNGI0Dzrz5GXJFj5fnog+SO+ZDLuQNq7wEmg5ve9lMK+
5/zViKlUpNdPpdgZtfpVCF9cDVuZCdll6y8hAeFgVDiwTazAZB8ESl+BTlQgohjZ
5QpgyIeXSmhV/dtZrK+0CaPtT1OuPgaItxm0r2gAIZ3BpZifrGt9aMAbqdgSW7FW
GR4xG8nPBAV8hCXges31uwA/r0mggzTHXdRCUKg88+QlS5gZcd9QQBpaO61TebMI
Gyy9z+I6pzSjNTAXenMJN8PWYwCim+z+pXYXm/1nCxE2eHclO8mnRIGf7pOocN1t
H/RGvVTe1UxblNz1hvzTveJZmXCLEPNtfqL2ORJ7PuwPSSXyb1PUXOmG9E7U3mjM
+rdJf1RR4Go1NWfVwlB3fxb6R7hDfDhUFasjSlvWGygXRvy1hZECJBWNU3k5YyQP
k0idML9euWrSDDro5gdXFh/xGO1zEMOziqnJsWSBVB8gUx2zBxY15R7AptyV0J8W
M/93EDuGWSVPhY38sSDUYf5266edmQ1fbvBD+SigTkcnMo+cyeTKs4bYcLVtXHsy
+8AVhDP0ydyW/5xx17U0FYaUfV0PgG69HXcQIxgSwIlu1toRkIgD/6Am34GPtTij
vOyl0+5rnS9JEAlc30Vh29WvXMPehLV0achgpBapdfaGiaWwBe15exQFR2OWMivH
qLDyFTHRB+Tq9r1a1TRXflLF58t7F5dgEtY/dpOmqGU3JRyWVBKWySydfIU7/eLg
MHKBsMN4njw9ZnswjJnbw7465nnjhkH4D9Ep+6QBKG9kKw5PViDwnjJCajTCuxg3
E71ZfiU2Zf5RUunGBmjoFD3ZiU4ejkdjyMLOkT6AjoI0HwtFUVUDcpk4X2h8UHdj
1t8ypCALBqpR9mNI3eLN062yUryny7Yky/jIn1RAHghM6eAewj0QMLRc9Ystg3UT
ZsI6e97c2J8v21iPmfeEXPlci809l35w6AMGFKCPGJknUTerwhKdWcwDffj5NHCB
hRkBdXy7adPLSNPGjogmnSbzBgSwg6r6uSYF40eYLPuBGJgxotB3sTyd2yEIEhmD
oSVbZCHk7POEWB1ZscSmLKlb8Hpq+VJ0vWuCetMl0RdPB+r8cO4yq3F7elFKyuuz
xsGompUzmIb9bom7Nd+4vK+XOfisFfMXp8psedIal+LRNmlWjbGiii/vItq3W3M4
rk8W5avyNjizZxeLtKIiCKXVMNtHk5AjcmYFg/AHRjNSWi3YrtxkIfkwH0OuwIiz
3/dmVGlbTwOdsxp0GOHNuymyF8E6jQLt+J5EpljLUkhnuCoQBSlbjFowa8QbfFiH
RcYxpo6xIGO1fetMon7iiW235veUgDpI8fYEB3WeL2XrfOy6VBYcJJ6mLcC0/U/K
uvHM0AC1ILqY8STEKHH1eCEe9NjCSevG7UrWJRz8LKq5pnaD+CvR4Asdq/+10qq8
eLFztOYm3p1KMyMllIlyHLjujotA7AfvsJ6SFJOuj3LbooUnxYzRcWr9yL3UqMYx
+MirXP25rDgeWW6IzQ66OKrY9lqYtNUbu8mcBEmw0N7aW2Lhe7vmei3LMiGni0vS
VbUl/5fGQYl3H4y5HjeUoeCJqCB/L0rvotJYachyRvPsqp72P3Q3zlgwxk2ivaoI
+r+tWHGmdCWeINJmXXAe17L+A3HM6dj6hxF+IUy35IbFmaCfrbXApnXKd9VOcC9/
arAtd3xIFdglpYce4by4flBnyTtKR+MYwIEkNIkRvJZIeemwWZ4GhuiYJwj/i0w8
TGdI+SVQQw7xr0SP71dWZzKo7nucQJYQuFB/lW4G9iK6Ietm3FrAo5vZaP93KAxS
RIx/PqeAc/hTlaZb6AcUjpb4oc9TUsKXIKI8jSSl8zD+XOqOMfiyGkXKYfcKCtv9
Qy19lGN9kpwuWYkj4fZtleLGT8GT+jB7WrLSshPSI2sLwTHJHpdlz60cGS0k/LB2
E1hRmxNVA3hfxlvAbnBNaYqbhRFgrQQD/9F/yORNi19Rr14bsvyK64c/lR4fIo8a
Ypwf7kkqktlF0p5NJP18mFLbgPiT52uSMidZFw3t+SEXe1X44ermZgvNQ82xDJii
pfH+fdTVnlLfw3PcCNIAu4UIsbwBZFNswUqxgBl55NtgpqrPV1ZgKWPITDNSZXWd
JyyxhSbFdAzTUNff1pA4xAd2sSLP+doVAhLtsntAJkrNEzdCOrdTyrKBhfKMhZTV
v/sJImC4PwImRRmzUqYKUtt9lsv/4OqO54r2XrFGFYJUWyoS3xctRCS+lGBMdYP7
jxP73S8Dx4bnW4wObFyugN2BIF92tNbnWFZ0dJxl122HKiSIabayQViW+fFDwubm
rlluJNLKI21gOYVGT5039M1OGj9V5RQdWCXhbqNlHLvOro668u6bYMsHO681NqxM
tEScRmvMK5E6N268EjGEj8wz01lK5vFhocKC/x7xPwuOCAmUiKWXUu4q5F0EKOMP
cPC43IEsS0ShsMbEwxOzzn2JZ6aBWq++1wHlPi02xh3onCvUZG/F+fI+EPQ6lI/S
z5TobLL1txUevTYsPUGbsDZ1I+UXN5mXb+aMUuxrH5PAX5iG7/0WCzcZ74OC+2Yt
FjYq4+dWXPYl/E3O5kKFV+9+0X6G1cEfXE1c86lHZEM4Z1ImLW+7on8u14LtHHHe
ddhVSSirGWL0BSscG6GTyzCiSAPP3LNHnIKntRoJgLOE4CDvku9/wd7I5HXv8KlT
6f1Dm0p2xXpuBeRnIjD8cX4z5NgSFPmRp2K+aO/oyGksMh9Vz2PPG52QpDbrt6sn
ZlkDiABO/HgwGB+MaTo0ZrPf3KiDmRU+cJ668Npog7uAgepFT8zfYLlcxA9Lz49y
nKrGIRptoWql+16S6BbctYNYtM+6bjaDMM9m3IF80KVufXC8yAL6u5FFEL6mBhxX
Daw8RbdKbqFBiDRqtlVhWtxdkl1qmowhF3ETlCK4lqj3GmSbIHbU0S8GlPjcJr60
ff+bQhAwCg4rpBSL9ENF0zHGOfY/ZO63RU1elbTTqzt3XvzYx+XXCmPFrBoraMaV
ge7QE8A/kxRk8Sh5MHt9/9RNASL9BeBHYypHhqrohyxOyrxqJ8QdqUegnB83kFVs
mZGdJtUWe4mlB+/Dbbdqf5yte3z2XPzqmWl2raONB6xcSsKhkXbukGzX/JN5MSFS
94w12N0HnnrYAHaxulupXDWYH3N90Fa9cm3VDBWW8eHn+lSSPn4UFE2zkcCDOY0q
7bYdBkyyJ0WCR6UmZO6NLFvnvjICBKocgb+vkqTTzQ44DizaYP4yExd58k6pSYWL
tetbeQizqw1Ovd3Q0CKdrqGMf665mrRZ/QDskJH2Ruh6QiJlnkcgGKcf/IzvJxcV
pru3xRpwDhb/qQcMM8MVNW0mBwbW+XFn+IUpnEfHd5ugaZorvmlh4IwoGNSawAJW
zQDyTTNWadWaZb8WzXl4JJk36NfBAUE7HbaM1d158GkCUHrnt+OtXiKwHyhkmnHl
nBrG2dqvvOLqDMcnGCGJE1elUcOwVBeecSAPn3xdKH/muChWGzmYydbBPxV2Jz56
s2qnJZe8LApUgeB30ZDTQV4iRCTs4RoSgUl5gedHcbxzmHXr1lxA3fm3U+0jNPYn
QwqasNiQaVoxhYDIiX6u3t91Tug+KxXjTDQ0SvZuLVzVWGyZvfrXnYlXAYKJwvsd
v+pHgWvh+ufdbzNnlKyxbnTJaVeQXLPZArKA13m7vffmxdknFYAwQjwTVwlA/T7d
lum3Grf7R7qsz2kaQhNUT4/9HRK9l9MMjxRSlRuoCNEwk1nGnNhVdRP76fB/+cfE
iIunR2PhzrU5M6ItoHhxAprU9tG1kn5FTvi0NcoZS41b5bHHY6ksz0B0xxtF8Dcy
sr2Z0HMeyNjWQSo+uORmSycjjD+QUQ9QDsQqpysS2Q/2YuvqltXfINCV/KZEVTQC
XhGSgmeDefJ54ECVJR6hZ/+QBV9mLzAtk85VJOwkyUkXglSzQyvHZiExHmZTDBPm
Ngu9ur0ZG/DPhTwajHzv4qStZbZoYSyT6UwjREp3EhrMAVHJEyQOG2TH2h/J4rDK
0CybsCk5kx9OCiajdJ8vUcEsOecrO97Ia5ZI1wxvQjFOdR8GdCxT1dBimT7hCw+i
B/Ek5/0VUDpZUmjZLiYm87NDX3wm7WmlpUnhdxTPi1M0N2+5tSk6TZWwtVao314f
kASRnFQ9crS3VzNnZyE0u4hyjyI5GsLMoF/MKwjA9hbEwrSDKrqTTT8nlg99W0ZG
2DoKba05jMuK9YWvTlwMcv5vh7tbGN3IxSkGxrvQRFk//grUrr1bA48nNK0/2LXC
f//WPgJTT5JGcHHtDUB66zsyNsYdnORBFaDMkE/jFhfobzqy0xtTiH8aBQxiqZBz
4A0PyP257k5ZoHtSMfxuwezRSnHJKeZuYmhJUTbZFQXIJwaq5WZzN9sHpETawnjB
2dZpD//EqkJ/m9wvoE8R/vAQfXKiKb8QNgqqW432TW8PmfDYpglDZWpk3OilgyH3
TP/RaXl3RTeCjrlzd5CXlzQNIF5tQQNRscvHiCWt1CJVRtSUOZzD2gUNtWZagmpJ
iSibFN7Cx/2w2jcMjh84rvgInb5//RaVDsafQgTcvw5YXBXVu4kK0NzZtM1GIuCP
TvsTrFRm3NHV1r0B3bA/IyD8vtSmzUiUQva2dZQ4UJn89FUBO5kOu/J7jcdGhaNR
ZcU3yraf3omHx+tFDfO6Jc0Flg7/3WrCfGJPmgc8cNalb6PaDH4eNeZeLTgZ/w7o
Emnhr2ULMz4YdGaKlsHLQZ1UjhBnLj/VaRxRs0OPGLVLTQYH+2FGTJEl2Q3EFQGA
HRyXjCecSFAHmxE7QwgWf6n2wHaHmBfUDaBSgKepIyOLnQbIrY/Y8LDbPp5cHh1D
caZLfhnEBzRhwUDcQiQEXED7zktzidHHQI+GlTTim0Y/Biqy7NF5W0xCK5Dk8uyq
+qRpSdHsR/ZQozOzCPZngLIiChFByvH6RXTevmysk3KBGtijzstJTunOEx6uzvbA
BBu+Ni61xz04xTAuTFNOP38uKqVsWyFmCzuWX0w7+JH+aB76rIUvU+3x4o5XFnd7
yB1zk9ifdKYM4+gi186yDYoDYlq7VIXE5+4DroPUBB5uU3AOaK9GCSNr03Jao+Yj
6xA0k+8DuEmErWnnRmNj3xVhA7hH9vKOYAzDKLgTRD4v+kW7GZ9utxxy1H5sCU+Z
BiS8OBF/01z9P9coXO1fB3QkgkFPLetMDQvwnYQq7QAmSPwfazQYgPC1hR0oKlR5
fVmwgBpMiIDgeSidDF1o6EKIbUrIPp4vgw3xwvpb5nryBxKfJN7MhPqdzOmwkgex
EuDlmmGtgbsFM7jzRM6cCCtx/zCIPeFM2vbzoqgkXL1sJXDZrb+J5mfSu31df2WX
Gl7vIkfF3sB6C2Hw52MJE1NfpnaqKd5Ynxr8X9cPotn/GRJIxQ9S68NT/6EyLe+q
csrA2hRj1VJa5enHPsTOU+iLrI4NiPz+tiA+3DKC+JJ19b928VUNxpBeTTvU6zL9
zzCMz5V2tOnlO5sEuSI2l3LLqui13/Pl2++gmnHddYJwQPBHRtfpy4mp9w3d5Jcg
+oe84c3UML1Q98dXMhpsuw495FZMOgIqCZVwz1CADMGIIOQRVOLUheCUY0dSQian
nXsDhiYq2qEmTsZdQfTAOqqwoTg9mlgehjzqY+inlmphgPeliExUQHFzPTq3V4Ji
h3EofQUIcFKlxy0kzijhNeGQ2sHhAVjuCaz+GagSWLFkfNqT6Mmtjsxz+8kWLTQm
quf0LWaRiHCyM7PhITP6LxYiYvUMrVVjLlyqVemXII6DPJT+FigHUh8u3OXYwM+g
tcwyAGnm6PgHFc/6d8helhnp9/2s4WeBD9U3KLLhieidObgHg+0AsYA6WXtzfRzG
KlCZSqV4/fewIYSl/j9+UVpZrcORNVveleetxujU3CkW7uByhjtFIfkJIj+Z62iv
475/+b9976qY7e0ndbcU17NxY6J/bwG73CB6hFHvf3OouzabIgPJtUQs/YTlBJEo
uIltLzZiEudwjil/xAKACxr/o3YFHN7D+yZaY5FwD46DDAMA1txZGZ7Q7oh4I2m2
MOpmubcZBDNtJV8SM0AVQUL3CgIE+3dKO0fjOjTwRcswdheWi4gbGAEj/FdL7ZRc
tu4FS93Bjn8medNg3+6TAx1S/NQqw7D7LkHnBg+XDLaflxZV6vPqpWUQptNyPvP7
p4NORPyZO9wIUWdWYlhiAgxdkG5dLJ7Cs4/dJZ27bu7px789RBdeb3rSM6ujRp36
BzOvHb+0T8pe5Chnje1LRhQOlFg1qSC1zca5Cmar/ZzeO24T9T1xC0aJDqZA1ic2
lmTqXbrrRkkZZXXRbECevzWNKuh+glZ9/JmeFzoe1oDpF0GorKCg0vhFTsj6BGKS
n4rLhPBWVzaKEGEF8KUDl8g6Z8UsZgFY4ML8FSafrOIYvLC5UsOdpw8NGZVTMqIQ
yweo0t61ql9gIXdz6JhupvUx9Zg4kkZiW89T3jSOVW5l2055aGiuTDpvdtsLyZI5
a+yxv3lpUpycCJdZM59H0Cn21Pd6pNme0IjiRYOZ+ATIbl4fWf8/FpYZpWQVyRsu
19GtE4l9n2XMSNCSGsVmyjJMu1eeMDNxu7c/4eoZNWLzcW3mSAokyBuMJjgATlNC
qpdbDoH9HCRSNb+GQb++dvIAqeBRxdeeuKyw2nJOSzPQPiubacPWkMLkt0SkULP0
N4mMEKONZHjLjRKeEXHrz8WP1YCk5xwSme5j/U5gWxuA+IsSIhNJDc5qM+7QVnQr
h9BGUpYLVyliQqL1cGqv5qGTRbrDX/X6ntuxGBwBtkgAFU3mdz9tVdzoxC2eOn7o
8iRCGFVPzQxglowzOdydXxB16Rq5Ohli3rtPnhqwm08/EGICLFRHJ9CZ/JjiaHRc
C+D+Ck2f3icECxpfnnWyZGLP6oO5rMRYoZAxsS5htX5QfP1kOMIfroOLCZd59lf1
BUDO7OUbu33jcHAqsbcYMJFUAMIdkP1anMlrZXpXYdhyji5I8cOJZvWvJvxxoMEX
vTOuTfr7NjcKf5QROHivE159m5ALSc0GudetL19I1qwXE7r31OGms8kK8fWka1Ux
+05Tg9qVXSJuPY4nrj5AZ3jY7r3POIEbN1HtKX2JA/4XZ+YZ8hUnnhJ1jRtTHa3K
AuF1h+uiZU48A/3ABQU2R/pbMQrM28zmK4taZi0jVGy620INjsfymLx3F0X1pgC2
SS8skYN90lAd3/WOJPhfUiHMSf3vl1E+gxd0b1xlJWuQUHsyTXd5Lz/CqFXWj2yp
YKBM9eVGEoY5Ki8L9YmYi0OLCpWxWuV8yT98HW+GcKR6mJGKPhtTG49pgF2amAhU
vEG2OVPidc61va8LPcbUpMMWJuGBCJ4KRADbGT1fj6heyBijaDxKoZ9shrWNkEDJ
Cx8kXR5q4UTVFhouosZacjT7FxMq7/ovQidnoue//Soy3R6AGHqvMUhAfDoGWRdE
RB/qMEPHNJ64EcmcJnDuG8dtVpoNvRZ/SpMGEd1aiOb5tA/CIOg0TI4FC/ntk0ji
ZNGjA8GtRXVBZPqKvcmt+1BZJecUvmTGcLu4rVxqlzY1J4f2XQ4bxlYbNSJi+661
79CzaKKJGHkSy/g4ARy+o9q3O5nimzeX5f0euJ/3YFoek1oIRapreK4R1JTQ+Sfc
pmkHlBBwGRbf93k8MrsQI88Hf151JjiTn6n+aX5Os7atNjpQaOTAGZ4pfDJYpQR8
iiFSktXweew/HnncqTt8A6Lz7saYBi9eRXC6Pey+Z7inQPBoB1qdAPfJ+Na3qzME
BDdeLgMvQNpJSH0CDsanItoC75qXC6XbODw8IhaG7CAVWilzgiHTpwVShhMwXUxQ
ZUWo7ddgqlFU37GV2a16z9UWuyLzUwh9pLSaQ4dLa1bS0qrW3BWX9MoijjP6gKNP
jT9Ed2M1Dayxe2DRn9i8y6IKeBlyGFqxs6qDVlKJ1nRt010Fo0KbU4oSi+e2TQM2
SUJy9Ws07xz5tgwr9TfTZljuh8CqRKZWBpS3ftJCePaRvuw8wBDyG+LUtXouO5So
SyggrWtEl6RJukNaGAQmUvxwoSefvHFcxmWQtZFDdV5qzwxgKyYvgwp0PVbdA6fM
/AQ4qjwQUs+7MYNSMFrQVsvubB6rECEsHv0BVhALdbOSajtf56UZDuGvgrkQB0Ym
qgO7Bnj5n/y3G2va5ffMXXMaeuSBkZgl14p65njuJ22mYksObtIRMFJRVmF3MUG1
Y/1aEMnp6Tfy2dsnW1EjrGebSw+2bcbn1baeG5hjq/Jyj/Ator7gf3cXkD336ItF
jL3Xl76L+s61nHtaDxyeYhUB/ces0B2pdHsYqXetHCu0RQ620ddtl7Xj/cwjODW2
n+0SoV1z8Ph8/GKuaxbORDvKKnS9RcVF2Nf2amauY4Xlg2BIAM7cO7QRpV46We6D
82CBwK/5SVwMSP5jYNylIetSfgBOxptii6MxZxS4gK4JoDzLM7hHFg5RdyJXtt+4
jtssKM8Y7MJfD4pdVWwDXOyaTXyP3V7veFZ3mTX2mbcEW1HtGosPWbem3xb6B9Lz
DMwM9hhVFMnoGYXQXVtgBgHSV7w37FdimNYV2z0hmEJ/ehntf2sohB7vtXAiatUz
y4ZdS2dyAHCRNLdrxgCjS2xXZ/KgL3IoVrfinqbV/Db0l8K+I0r9oqO6PvIE7W18
DZvIvur2pd9GN4TLmRDnh1xzmdviFTvOmPm3DckoeqEHB226RZFcArxbMmdoXesk
rfGCb2YQBfF5RC043cNJ3VujjXjk4Gm8h3ruJY9oYq4/36cuI72AGDKl44qd+8zh
P1XmWUWHFMfeoziwKgJuO+suH52eDJfMmNtiOKXIgSmFGi/A9PFVJZH7fMBk3/4a
wLo6e1oYJ6H8d90zNDYg/Zyv7RmbT5KdAhD2R/dfBiMTGrpFaGES+YhatGL4PCgJ
dGL8StIs2sk/Jp3Hz+BhmaTrcILP0QbkgMQi4455hIBVS3yu3UuCqy5IJhpmw4ao
KTz/K/hHxVqBUMIa6r4fzMFhDef2P9HXq4V+7nT27KKktbWgyUI51k+ySrKL8ez4
pwgQI6MrC209BSn217A16EcF9KmijoTWO8W8rCBoSGFO5K13qagnOIxWgTWupaI4
OsG+EhL2h8iMK+YiuC3zGOSbg6eR/rWfu4/UfIUySrbt0Pv6SdT4P3M3VS0iBKar
aJLD6LCXiVRypdwb9lQk8LvpwShZcKh1fR1g4JLtRv1dr+aAICC1QLXWfv1i8lrL
nAFplqJFMHUoWeU/rvxHN512dmhtUwrS0SpUnT2x598oevCzQND3fXSkUYoIePoJ
xjkKcF0My6smay7h/p9hHVLiigqS4m5P1JIfCJfoqMfoR7/wLYBoyYV69Yr0EfeR
qVwDJqYIfb5t2Q3h3Fw8HfNYASJNqIHZ8GD6wxLolHyCHwqSiiQHSJo3C/hixWLN
X7FodziLJFaPWn5VFhmkCSx7/QhmOxn7MpCOkBIT9mHetffbUS6OUoIoZ4v30ak0
L0WUBGC5X0+1QdRdXl0y6Y9iLjKB6TyOG4RoSvqT0usAaenBXSc8rHjgL09djkux
RKzqESgT4QI1RNT0ClD0amrUSGwc1tvda3TQsy66qHfJ8Sc5PHcY1qxt6S8+OvlR
Pv4zpgsAkGflu7qjcy8nZHFZM8b10N93dtfcIs/F3TyxpFGXMrN3duO6a2S5hjql
P7S5RNgoQL04x+rLFvdv0oTFWZhLWDpPtLzIsp1dXUKyKA2E/GClbu+QPs22G/nK
e/JaE2SQgXOePObN/q7IAzBRK7heXVOkATAN+Owqr3PfkVCvUjrw3BVQcHfrhiit
mEliWmFg+snw+1e8XVYDonLib2njQYOPLRjFAvTf5u0546zZkhN74M1WAq+Dhekc
aG+5IAmMw4gKVVYSHidXSTDrLM9fpeOyStcMYoI19dRQgeOsFqgKEs/qGCu1GPKZ
UH0FNBwMeC2rh75R5gZQghfSvX7rllGgUEBnE8qomH4SC4qWdI1ppn3HIBwZtmZA
X1BxD/nu1c+tLOeP8Na1Ia0EiIuN/FUVAtTkq1TsH+0LfhdDPlgNhXBgTuks2r9F
kYnsZkGoece30LPur+RqJ6LbG2+EN8aJ6t1LC288Wz9TDIsSkkNyZK74+GsoLvWX
G5ItruqmU4O/cqIgQHLXHXEZ/nBqDh6MldVmXKkD7oMbGGtRzDc+wERAZ89TEvkz
aD6CBbRSkOepzxTMG6fOdyMppCtCEUWsuiUZ0F2Cec5b/VwkwseU0xA7xTdz+6qu
OKre1FcabxSxKLLPbejG0BlnL9t/3g6Z+DmD4JuoMi1FNMUsOwg/EvmA1XyRxiqi
//dAE4tq3i5DOyU+wJ7YB6+dE0EcClf6MnNGmbJTpbaCICKN6ytGXildtZEohu2T
8XH3ky6DRCONfK3grkivO41pXXef1dpj+D3aOnRPWuH5eNHKUaKd/ufUpRZIKiZQ
iedXukgp4IKe/xLF7pe3mrcDWWRiY2hv0IAuEquk6GqAv7nlAao+cHhfC4g5VBcY
VPhOaoWb99pP6FJo/wPBICDyvOXVdONsF7xmH88skJHOH6pzt0CRgxv7vBOJnRyO
v6K9t/YzoTQPqeBFM67IegC9VG5heQi0qxp8kfdbOQyMLOS6XQRd8Z5OHThlIoXo
rv524c1twzK2hUHxc1gaN5BQw/zDeq/uPfJoEEBV/plaKTYValo4VE3WsI5+/HIt
SdMmmUrEVUBDwGmhSI3Jo0jogdcJjDw4QdLUrOWOFBdT7iNbdks8XBIdvQvpYqym
+efaF9+JSFjqh8m3FIRw242q2tPfsYmxHoOSP3i82yade+kEVRD5hPlB7A+68VbW
YWjUhEUW3ZO+6RHF0KbTgiyXyoYtb7nTnW4+81ZU4ijagFfGvPbD1fxowrORKroy
2N5QA8fAmaLm5Z4l/K+qH9oArz1DOMfW77QUY4y0eO6Uu1mX9P9X4EjG2QicmBVG
rQ9XLR4XZAg/6p3FeNEyXiGVSj1ODWjk8krkY6RujjM7kQ2vQ6wPAMfMoYpSCHq8
s05oB51gmErj0nG85xrGR3dFK5BhXMQtLBLnthgClvtKDL0Y9NgQBLDr4VTf0v18
5b8NeCIcJcVktqpT59gRGdm1OTFOLH+i7AOAiev67CYioLnH4UxKdY9DH+zkEB4D
hGxa++2K6YIKXIryz0w3Hg9PFpa0lTcC6B3qbiogpWiQ8khB59ZKSuOXQO2aPsAe
0kyP1RKOuWFuCTOACcHpfC51+IyGnCXd9Frcm9RvlQkXVJ07qxNJjPdwoiBE/XeF
0oAdclh4uMnZBy5H+k7AB/vPWOaR+/LIL+qkUXnd0c3yJuhmgViwFKUnv5qeGz+o
daItD2VfULCwvTe2nTDF6WRNaoVu7b8JwQ6S60E3wRDG6nyf3DrGdB/eSybkPWUy
KSf8wjGjHPnBkLwgXohgeow4aCA36Vj5t0Plcdhmd+vsFNI7OxYOsvsJFl4C58m8
J1bdqZdnSP2st3s4RQYn+DTtO7Xjmo3s+uBH25VJJoWRM3lziFd+ZiY6COke5dMR
wJQcsfY3Xot/tJaXbAYo/ym/O7NjUIWd3ry7OQUtRLQK03C3+n0JWNGTtV0WhSbv
yEzNcer/BGv9HFMlzCWK0KWCRyEfthXRHyxdtRnracJ77MfMKClNYvQKxiRAulZ5
AnBQcvHAmBloamCpeVr53KRzrf/uTJAGGb0xOtji4kYjI9xJqQL9T6Mib9bihnwR
9JNPjjjk4rVUrSBFu/fzlsCWl8nLagneBJRJN3/+9NA43s7PHtXe5zUnJm5nUVhf
SYDk+0euBN10D6FUL60CNSZZwJXmd9ZkvdDNn/Ubk/MK8pauOZqDDvgMSsNoZxj8
wjnjqKAEpTcEp1oV6uZzwo6LavVagggLQUuvHIZduzz6SlhyAPRXyQQb1610BeC9
WpDK0PAD+fM5GexofqjacG596XuYQO1yYNjMuTrf4GfeojnUWsJfQAV8+Ys3fs7K
rMNuQCfMVloSJ/PD1R9E56wek3iFiTwVsB7VSwzMhcan2t4GHzIePd01ap84mJ4+
VuOK6E7UBy0OPgbpxnUWhy0yaqsfK9WYbbgFyOOhCbX4rL9B9HyJjwoqR55JzyL9
CbUP7DtiX6S6SM79a0e8sWTB2hAXYR424yj/eYICh1gUGVyjWYHqNH6iLZUQrMIM
6JAb37lokXRq2a2TCEzanGPPxfma2Fc7fY5EoZFV/YEkAfvvLNPcOdlFxhVcKX8c
idhv35FB2ZyK8Bm9/sWLB1Y3RRLypI875WckqbeurPgi3Ha3B5BWvREdr08Ut6xB
moqb/N3cjcCRufnytRU0cjK/V6ghtgSUBfulSHLo5rxR+GqiMI3NAX+RLjlvtcq0
j80bqbRQgGlLVrAZkOtpMBld4fNATiiYsVPBqI3SUTWBAAV0N0/P9NFanzV5dmHn
xzO6Cseu8qDQTyzGaILLojP6gRrIiUB4cl5x/adniPJm8nTpCMiSzjVBKk3RSuPs
8n2STHwayLXU0gwUkt49VhCfLmF7UR0eTb4A+E8lBmifHKm4p/q94wv5UKC2TDsi
7MuwHfNpjHpVqeohms8rD/dLWGBu1VEWee7dU427e9vW0pTAZBYWckQtpeKxKDZY
dZqI5ypEEa7rvaa4hmVeHdScYl8bB+6X8ACyUGrQ38BsteWndY2y5fvzTnbeD71E
xr+QZTsYyi+FOKbk20KkVgv9uHiRhtoU6iCjS5i8KcGnAWD5uoZwnhJJP/zJQ13N
M08FS90VYlIHz1+VyOQkxIlWJGC1v/K2cM4aTURD3HMF6afAzRuhz5nNpGZ8nWs3
O3vriG4LwRDZNUgNlkINtXf0sCo/r47im8Ji4bS8Ag7Ay/xpGT0Acc4X5+Q7YXg+
rUEhzYKVIfe0I02fIXcDHEBGFSsH2oXQ2jjSm5A+KEY0M5aH5bkz/11LRURtRJo1
WQf1dV+PI4QcI3d4qLkiIRLXYHSedOuoYACL0LnCchYzQA3BMYra/87AzSZ8rWnC
BdFTZArmSSyZ5727WOK/EmKxwmuhEpDyXtRifxm3Rt5mdH5K0JS1eDkMj+6IgEZA
a4xokstWiSaZhITXD4/kggHgrNCZW+ysprt7hDNMwlemfpQeGq2x55gS2/CiNyRt
8AGE6l8ERknTW4KPjjlwbkM2jgsl/MC+Ir1B13mENooybRaNxmLo10FDumywsJpi
bwvqpcdc3ZTWoL4OJXkdASXw6VJEiQrkwPfqAcVyojRBftCw/3dO4NXsuLTnoyDa
22rd3ZJUe9EPc8/HP8mfX5OdSlX05cJoKqAYjJa0bkfsshj2A7yaFNcU2TQqqZcX
TJJtBPUj0f+MBlKif5LBpiQQ2h77Awb3vll7HZX6m7DmqH7HSfbJmbCnc60rhHWb
PHyWLka/y8jvD2TjpjCg8udkEvTHmdI5wytn4Mb0+8pUTP9IzsSS6wDvUAPxw7QH
zpFiJcDFq8aFVC8iHOO5eFqk0Xap9SpTfEnemnBWTaFXwE906OR/svtCxHAsPlWL
qSK0lf9SHJFHbyH6uhFDajEBBrakx9oxN0hXUCdm2Olfqb55Aiu4bIL0s1298+kL
xW0GakGXl4e0YMScpBjiKupExUpiCP4KOxLJ8bhgrGOCfxQL+4UwyYKN3iYAvZj3
HmNGg9lUA3MyUGTk9p+RBLVjjVGYAJvqs3x7hKzHQjKFo4cmChFu8SYuzkpsC5/h
W9FCZfTxro5KjU/i8xcQgub61+HQibosmG3hu1wHU2ByO0iHK0lSrwyYl1Zpp6HW
nzGWQZ+pB7096sWqLcm1Ki1DLlQl6DM/rSEiTGUlsrCnGKOqYhcwNMCz3fVBeYLZ
n0R2i98i6LYzHR/WlykjHfJsQcbn3xfIgjFjZvXsQlpDT+v5k7SRSnPORankNn/6
r8ugec/4G7V6gUxaBmvv5Y4hDPjKYonDajjia5QoKjjQ2VNajO8Jb1aNFCzL0HoF
ku0e46JJhUL0rSABJTGzGN5kfLnILQL0FKYpU/d9XOAYSWy8ga0WduuqgZjdd4uE
7iXmVXdeTDnI3jZwK+p8f18X+ayuL1m+lUTZogL0TPYSHYlXq1ZMe4UejJf4k9Wb
p6zHlyZemlJfKe0G31I5z3b898TZVK8OhLBgMF27IAYMQmjrhRexKzFQ5c3QGp75
mDcZgsTedydYg07wKfW0xN29mysK2toLO7K3Ey2em+wCppAU56LM0eiN8KrvFev3
gpYGgIbnkolYi6T0iwxSrSSCCsfQ7pMxC1kKJD1rzG0CzrDZ32kaUP8nvvh0XBSz
flTAq9ajlLUDxJkQZvsgyqJJwU+/InI/s1YjoYflVHbBJ1sA6uax4i/hLPff7GTj
BRFBQszncJfk+BK8UIMqias91ekWwWRmsOnyX4uJrirfj7wFZRM0KAqOBKIiJr4F
Egm5ACVamlZUB8HZKenbiTv5SBpo0U74ge6GAk7kq21gfXcPF7ttfiNY30Eg4Hnb
SehZTpOEvtdU6yE3Q8dOMLpRmCT5wJfYerXcjT4a6n6utZA9J5uwdEZEG7VqDQKj
D4cdxOjg5ERK+kYn8X0GeNJW+f7yBK8JuXsratJEPHHt6clemmuqAqHBddCDv/C4
oAmGjLIf2xmtsK0fLJif8i+i7WFc31RIZB5BlGwNyPb4mxMvcK/5hNEV+XMmdO9l
afVgvtj9Pb5RYgo9IDGw8CUoIu1bab9taX1gCOu27d0K1gjc5ccrZKrh7feRCCiR
qJhYwEhXdFEv6oW8We/OR8o2PywMtK+IPPy6TWE/4M/Qa0M6hEiFzSmjxkr2EAIS
qj4FKLbFFZ/megiw4zAzXj21uJ7USrxMPGOqWOMQolOtQNjwpMxyNR/6E8v7Pcn7
sBSUc1bo4bu/3bax6tSnOCi87F5ipVtKzDoO1H1g3hXmYX3dQ27TJYZ9QEzk+MNi
fGHz0LscgoKXL9I9jes8dyYpPQx8BTJ/RhUL0h1SiJ0CBcPTMNtoMS3MI9Cm/COS
2sNG7BEV8dwFjb0piDMvy6bkAEO4X4RE/Q8A6+wdPQZVjwFxBHkXSy/z8mq9wN7/
gU5j85+x8cuBTQ3edbyCXq20vjIRww8z9OBsRt42Ijk9fyWcrSWBN/Nft5Cnowg0
29OVheAI+bgMI2pKsadtYoZStceeXboAaGYrMuS53eK2DjymrnpyMThpxk1z4vdu
aUq0JJeU70Xlt3KTobR1qNV8ZK/qmxiIE89yhyVSOtW4TAJHiXM2Zb8W/+5ONWUj
Eaj4qXvuyq6r6nVelTFgSRB+qeaE6iA5yFcT/+immEXFHJHZvaAW2M4j11mt/8Ab
gZ+Y3MdvzHbpA0K+QzD942qufdYiDd4QvG/Xde4lEN/ANwIoU2SHtAllqlSTCpEf
NogR135cs+jard1rBRG/Znz++bynexRMWC3DOJNwlkJ0I4cny/VCdN8N08NeLeKQ
GcsIIZ6JDOAMeuMnjbf+bhNELL2O3das6jTOZ/3eK1cZNOTS45Pl9kSGHIN3HEB0
vwlWpmcOnGB2TdvcS8idH/ODDVqR02xzmP6DHSIeGoBBl5IoWBDyoirAB+jPuXax
lvJe8dLFsTc15x8qCExe3ISyd80bxR0Yl1TdLGtEx1LjCydPOM5Ty1KLGhf0yyAX
mj+NRrU1pUPQd/0yhmjGugZUqmqrj/KWI3dcd0rlteJ78bPNvYnTB3v2DVo1pO8O
k5Mn5kiTCzWChcFeRwdGIRUJUCa0Ovk3O9Ghbf9PBtyqEAvpjf1Qp6N9hG+1ok61
SB9Abjfk3+iYDTNUPACYkhcYpZnDVu8uCTql1uM76Vpz5ObTL3ijmlsde+jXcLc9
IIQiD+ymmpKZxK/jt72J6R48oculI3fK0nY/LU9Q0A5KSIhu2tTo7yU//BN0soBl
oXuJTEAMDp2kMeBhfG7zlbTqIDZ3DzhJx3n1sORmwnF79JY9NA5uUQEeKfmIEagz
VooCQ9X2HM6Nz72RqRr9KvCosLRgR8wy+IJIMYGq8vLWRgZyNlDpN6HtCO9MBcZV
cuCehiWoRo968q9cW0iyTh0Iq4hgJ1fppMfO/fqHFri1BLX0VgpM3r8xCFpjCAJr
o4DgxuZFWhdc+AqRBOxlJm2CFRG30JLVIhXKV5//Eykctac26waGaaLwuGOrwCW2
2jZIqgkuSdCfBEChHY4PuemHTnfdFQODfYYVOGwJkfutYvdVkLUOGtLAkXHOENOJ
sSVdeOehfvd4i/y4aXmRNFyHncC7Ln8hZ5cDXWjHDxvfETBPYGBZePda03DZhs+7
rph9Z7roYabbKvrnqR3fTDZM6wRpii+fVXhSm0riJAz76L+YxZ6zutBfPiagC0yK
vvZdZ/j9kUShxK+S8n/eB29csEY0b1YhWcfwPA4oIz7/EB3L1Ni1tPDCzIIO5g60
JktTcUyNEtZsKRFaqyHxZcXLrNGuO4Kpi8jLZvrotcIBlPgUIk1ya1xDZFe46uNU
2VDSNouq6jA8I1ui5C8Olat/iCPpl/resKw/T3RO7P1sZTFPDukftD5z6YnD8enh
MwCnwZ2dYkWTs23Trg7VqhlchRHflMF6qAArkCWGAO3cAU8OI29iVyiADS52qGRO
EOMByGt0bbdm/fMSqvsvoRV4Uc94fh8xWPol1HuTjtHv+n5tW7c+UZAHErXxR3kx
w0i4GlXDH6iAXQrcagbh8v/Uqc/Iby9Vq3arsevUvhAgefxY+0RhmvJhXVweTqNQ
H1ncSiOr85sW8lvK0TRljCiQexDeYMIQzUMsG5dzbdE8CEHHxFNkzD2ReH5Arj2e
OtSXQWXZlUsCM1oZ0ZAs2lgAeUIefPe94mysq0qbGirQWBOKb71uh40Vv4iaFYS3
wSyf9pOgfizL9mzkaLrS4pUp8J5vhu23+/HMeLyooWOcneOOcsB7sM4dVLLoBVqk
pa4a0ROMT7Dy2+OJeSeIv4SiFOm95SV9LYTagz4sRJF+r+EUIrszd2U610c16PgI
3YCNw0PVRy5PL0zS8KxxKXqlS4FXjF3ZU9AqvP+VDOmYvlfw3+GOEwc2igLVY2uI
HAYjUxDKjWVmINTry+ge5VZsXlLt3mDbpkRw2yRzNNQdkCxkqvxuERQ5EXOaMrEc
mtTFPAWjwRrUUf48poprG9qtEiJZ4e1de51HdLqvDuRFhhPCGlQkslRTs5JBzXII
hjmCVAynzjC50b/I+ZrfcBNMUD2F9BIgXLl+xnt2NDoYwz6ZE9+lMw3YnGZ7ZZse
zbILTAouVuZdC3hCNL8CD7n/dNEyYwarX9HNmzlWHOMR82jEAS2uAzbssHXa6IwX
NSQGyIEw2+GVOtY9vPFQ0vREDwHmYHrSSJZH02I3OAvu610mctfkzkYmw6op/IE3
YqkTP0dm2xcR6p6SV+82Hfkdrpwj/YB8aO4rpAWZz6Vq1Xk8bhah1zviJa3vSEqW
kkZlaI9VLTl5Syj/9cfBZgHaw47JULAW/epTxKNXU6HK4vZIT/SCzRZiPFTc5LRC
FnQmlfonpbBb+PGn0u+31q3TrR+IyD1zuFUiVzpclnU4XjS+ZLzb+0Tjehb2Jhva
NEXEcWrJlOw0yTihwrEQ7EpgFgkL0If36bzKfRXw3yVT6/mUk1KnQbx1d+44oXP6
fMm66iss7LqNa+te8ktDaggeyLdA8ngSbOsuPciHR/6CMWLa6rzWJXOrs/3+vzjn
4dRtivdQl2yHyYP18qKECqBmRzBpa8UId9CU/sSOuuIxA7crJpmGE3IvW+ZQkQ21
1/nCYjDErIThlvft+cPc0NkjHOc2v3e6qkwNBh49x3DKgPqvF4WVfRjsNT/3UIpn
El16yMI01FJDPYXePSb86HZrhosw/Ic3NgpcIIETokOPa2kMDscyQl7TqqsmZ9Cr
Xz8QUKaxJKhy+oAl/rTWDQ3YVd8ZET4I9edHLfDpcvVBbkrR+YMuF2ZWFwRMvHsO
xIN89FPbiY37R1lG6GqMwM08I/J3sT6H4U3S5WNfE6Wh0HzkSkIgZWU62GCxybjM
dsXQBYReCjkgzjHREhMuA0pgaZWVSZ+6RN7nqhJQEoitmsNPUomr8M14oZb4b1LZ
3nR5pIDW5fd5UesROsglc3lBCnn1ArCmrP235Xk2pPfxKNe5kkpyJ8d/ZdNIRTpV
VZwnapOvSJsgNK+VHGkDWvIp6o7/qKfE6tzzkm+DYLkJZ0cXkfz1FWWHVxNOTCQ8
z8lDWdAMpObuxGcC67HUet9OvZ6SxW2OEpljtscJCKQUCycUlvAsCouC7D3z55aQ
AWXCcEgro7CIR+plj6KcfplkOIeOlaW/FvQymH+uUgR0IXMi2nkigt//9aowz7Zs
MfGBtC6sPWMrmidmunn/e70r+bEJkQpzbHYf6gKNU1LB8OLradwlWZ0x2TBZx8d9
jafzBDNhppcfuDJvTt2J/vdf5H3etfSav4gsNegAwu1yc5IquQ/9RVU+5ebcyIMq
7SlSl6FOfRz7Sxs7y0IMn9yvebG76p5I5CFphgep4mQJrfZBkKlDDV8B1D+ZafVk
jzxCF2HX5hHyMxX4cxxiUP9uzKUtHIf3zWYraNGPuycIl9SvuQVXUNcv9Mbhxfif
i+y+y/tMDCnZEXa7eezYyiJRJjtbZBYSpPMQUuN2KhjTQD9J+qPAz4oG83uwEXmU
5vcaYcNF24gW6Yx7xTHrQhkZ1Z3SC0G0GzHwMxcluPEsePJWXzonkmr+PYJbOV3m
AnOO0JzCxPFn+w/XDS9REB17xbJZBDn1Ncx4gYUhPcy4fSMxHE0BBawbG/fgYm5v
DHxiOB7W6QRI7F81cImZlvsuFxocmS3eoInmA6zWFlYZXcsVvfwWnVLTnzTZdNGk
g1yEFi8XPZwag6SoQ1WgokDD67+uFCDD4Xm6toASy3MR77b9b+V43AsSUJ9Woa1m
8BCmL6qJOwHz2bTOcSbsvlX9VnaJHh8DLqmLkIFckSGy1Ws59m+YW9xwBlCcjdvh
1aGgo22MpGG86fhyPE9jWLIlbDrtCDY3A02qjNVzbqy9qATVCQweCAO08KxXGolV
xxBgzq6dvt0aHWHun+TcbnV983+a9mOZwSeyhZjqIJykWRyBF5idkJGNKrV4OgjX
RI1U+KDV8fT1FxcEKaY/RTp2Yo0CedGVj3NiEgxU5scT3Afu7+o1WC2Ful4aAbHC
y0tFsQ1E31CnY05NSSoLzZHiufuaeMA0kWSQ4OWLF17RAfC5xRl3uaIFhTULtBLf
FB5cSqH0CyO3VVvm+dU3ab31lavvwtM3TjZsttPBdoJelCC6NDe9KUCvmXFJUNGF
jfLuRvq5Nw+gI2CQNbEvI/bWaPXRKGMGFZlkkGKgBlKBV7HkpC3xTKUTSYS0WnLU
Ww+AKntPRB+x7Vs4f1tozdeUECVKX9gOiXLDhkhaXYYxKaOynPFsRe1SCyAk2WHV
kxqvbq0wBwOsyJUXxygm/eiEpgEN6b5eK3RiQbwffkw3vRxz2POqiO5ULgRs5+fd
6217P5tyC9A4MlHyWBg7pVXbJLaOq+ed9kPuY7cjJDJ2HxiiMr7mkdyXZsCdOdOe
k75ZKVb6mrJpMZb32njxMoDvjU/zLCFWu0kQLLQu2h9sA8X+ItMn8twWyPbXHppW
49x3QtifG2v/BZjd3bABDSCMoxcIXt78g7MZFNSRJ4hprBs0DLagW3cGttlBRPnJ
USpkOkTa/XOSf9YfFRqCSBit6hgqphQo9lYZGTTzc/XoxwOB3iQVXSLyygxJblRL
O7sI4xwEjj1EsKHFXTofmhTRsooaAYNclyKDl2hBzK48oojpEyOZyZALonpJvKXi
pFlqldfGjD3DAR3RIhf8lmYlsnuffDOuAdZotSWQlzPpLL1MLR58z0BXrR9FtEx6
cppk/L6H1rY1c4rCm4IMNnfw7KeghmNSrBqTZEq9/aBtmnBN7JMQsitDBpygdatt
eSbMx0TjAP14FaZf2IqFA/i5Yi0wpZ8DbmOlOYNuS2wBjQkTy9Tbhd0eGTXSrJzG
bqvOQJMdXIgvV6oet/P3I6X944kdFjadyCTOe9Ub6+Iv2lj8B71xXbyz6mdN4rRV
aLa5OO7SdEjgB7kFGulCNBVzfARpbkui4Zubh1fEnzt9tVPn54c0trS18cABwyTw
Inc1RhI/lMxR6uVUJaCQyHfXjteSlladLiGsRqHm3WFUmPPVBm/noexY7pDcXhHw
dDqRfXG/WBvITyBdpIcd5kJ+EHYJEaDLTQDgJJ7m0LlRBjPiUpocrImnfEZxspka
wNwFBYOjus/+cGQO5vX1hoJ+JVBYiojgTz0BaadM0yQRRPUM82n58kjp/671Pen5
Ahg1iMsUVCORcerQXQPOeA+Pmxdg5rQV7UTfjdpR7cCzqwSGDxwZ4D04isThUqNK
6S3mYB12tM4HYwbd2uKodiBPHGH5PyGHw/3BBTiFOdBNLRQ6MqPJigU9Fg4RnX1w
nl8TyH3A+4ToKhLcWOmhzCs0parRKUcFsvPU7/+Qo1ixmwAwfbiE2FXQScQZfizd
QW8PGjz76HAqlTyHXo6ufoHBpgRql0hGXKrXksuEcPOv4IJb18vVjBT9bZxf+rIl
sXstAgUu8GWstaAiIFiKeqlWcxbXHAdo3EAHIFxlZlCtmHaJ+z1IMnPvsLscMUTl
1232HNBnNTiXYoaD9EUXfSJf67EVE0PD5a0IeeySTE4M86NozPeqRnE6svI03k0V
LZ4q4rVz/7KtT9FgKF5XlAVGeYrxVtk/vpSf0DL2zakZWoHPnhOahXOgFG0shISV
5pOMdykRHVqor8kEUfJbA752veao7KlJ4FJOIFjoZNiFLaF9iN5etdW5Ktqw1klO
Q0Gys5OpNab3z5DkAcRkv6gtmXLJGLW2x4a/3d9h/lYwVHrnYzdScYCo217s+1EL
qr4z8L0c5qif0IxsX9AI4CWIFgndvTT0NTbobZdPv4obvMwax2UrHRrCrckCDlm/
rCxzJirUrfjVTnTeQ4AM+48Ek8LtrfN0tNfknsL72tfaT4rpcHYwu57hiZUyOkf+
CAi3XnbWA6GN/jzNl4MwP2jRRFBGZHWFkNVGc9tzNq2jonHRbdN2tueZoj8AvsRK
pj+zlRMTqVs1dyPS0plsYLRafjWMfWTRxUa9EoiuSSeK35fT5mNM3nDF2JGwW2uM
b/5Xl7A27YrbylokAEjyc3KAbbrx/2gvlTSpRupUnz6B3LqY/WUYuOQ0a4FUaZii
Qbaj0iqxvovUSa6i7s76PlXzFFhq4pWjSaI47r+w5TvmrD6zsIIIrpkx199/TGCS
Xl5QfjCtU1XDBQ5xWcPpK4GxXc0abuGTT9KTk7I4TFCGAAUmCcQsISoodaEtdRna
nXZIYyP7wbVqrTA9egsqW4fdGSPDHZ+wYKOLbIUzwc5Bx1TFAoCA0k5xhPMx8daH
RVRf2Br7K3TPsawlGIVyoVNzGIvuktKrTQOEkY47sS53sZtF8jsoYdPB9hJkOnnB
19lRdezSfTeowAe16s9SYsm5XwFeE5RtpjUjWh9DoqkcdtujTweNw66+b8wu+OJU
XkIwVowvW/CF+RQaGzzhI0uwZ5KbU5jWumJWTGmXU9ySqMSKzZmvoJ9GUm3TwwAs
ZzrCXW1rbXnmV0CxlGqWDfELQ5HWgf78Ay2qCMg2RlOh6t4g9VSN7p3WDHSpyJoy
kAG6JGf41JpoVh7eF6beUaqIFd54z14VO1g+LPl0BqnAxFFik9y8mfAvvNzzGzdS
pXce9RVRzG7rvkV8IRXZ6tTAiGV2v3mwPbbEMJjGBR8SPx3FQ0My4kvFbBVwVayJ
fwzTAZ7XW+8Ap0v94CwY5tzYSkvh/rLMNitSx31odSyi/L4n+vCXf2z/HuaXmK4p
kTipgRPnpenDrtyhqKc0YZqmrTVD/nUJjdaM+lxpeGVVF5wD6QNvIqTHU9Byh67m
PwNQiGzHZZ2+wdGa00Skmsdi18YAD/Qpb3rvUpHgP5XFvUsD3McgZD+7hT39fth0
gorJSFRQaNCUPz5/gfTdSZMoRRU+BUlyuAkKRhrWmacGXfl8vjzVa3mtp/JkMEks
bCN2Ex1eAyWab/Z8ln/rSNLsDqNFWBNGIabx9Q4vsSpQd7YW5xMxlrkhf0BXZktT
7I7ewiFuuw+qxSsQ8zV0IEdY7ABXv5QRWxhclGM7aZS87Wu/wCSnNQltVLDxJT0c
wf3j2qxloN7m9zHNODJ+jFMDucb1cs23hCqwcSaNYEnrP+AdEKeT+n01XIsY11ry
EHnNWCEVvchDaEZnEfK89yPm6wws3EHnlpXZonf0P9oTy7x5BkT5FPZlLvWdOglJ
jdGzUbAtE8Zb8ub0pOkFEmwKNWH4cz4BmhWP6TeHHHoEa+wxQMAbrBBa5nN78Q+v
/l/ge6Hu/Jrt6l5A0UF0/YCjZBLZOxHmd/ZsRjgA9Y/TNuEUDhj6PWi84cAQUEda
iN53dYFOL208x0/j8+jGf3H1SSA82VoSVkS3BbpEy31ybACPe9c2VDanRLXbLH3H
ePbi9I7zeBKt30BchCx5RSaZ+8Hb+m7HbNNJ0xVu9b6dJlri2uEJ+w2o/fJEfSCY
WqFvjSeQk27IKocCQZrI2oAisXV7MshtIUolgvuAUYEfpZ2QorZrFOQfKHPVMyGL
/bGDDgKf2Eu3Sf+Pm8jGRhIwCzsF/LZTUEpeINg2IScyo8n3AUkOeIpuJePXlXdT
7JWSG+DnTvEXNBLW9BFMuuZ39N6m1MNhPsrrNkRETskch7LFI0AJ3OAa5ZNf14jW
87D1ZdAD7KoiDsNlfg73AgL1pZH58ZY5SdxTDZoHtKN5PLQABNG/lPsbgLiYUosM
OGAL5EnGf4SvsrPczMR9p4BLFtsqDf5FkOCEwWemLd0/y+05JEebZZDV2pTL22Zg
EBdg8KJFR3TJMlX3EBOiPVXxo2A+CucgkVq1OW1xla2+APulsUDDe0dqt++mHiVd
KtfPwuA3Vl1lHtxZa0IPEX9/sSdwSh6Voi5r64Xb+DuvPwCAtvKYaXH4frXdBulq
s+hYRpWvCk6KAJhJbdgKgeyh9c+Gy9bRNPQ1AY0NcSueUc4Ub9nM+6sI4sXlvidS
PDdJG4Pqy0xy4MwbB0Wj9bmhTQNs2lWt/xRPOrSIIEiqV7dTmI7IfFdWWvRmz5GP
UbqpWSVHAbyu6o994mAQhwuTNoR7oRaDaVuwaIID/wwQdW1Eg37r8K0QWbjWado6
FesTBlX1aQ+PjEdUtQl6v8L6+iabCG7kyWsRp6ust3vlsCQM0mCF5lNUEOn0cd3D
aM8o6f6iP1k1VEclsd4/F5wgd9kMbBEPwpfwG75ht2fNZgRBfeQpy2ONM0PR+1ak
Yt5S8/zVLkwwlZ0fvomBOOjZEblJt9WBod7x5GX3ByDelqC6HWS10g0CJ7Bqh1Os
nYNd07JMHH2F9pnkrSCj8S0xdrykzJyBRX9JZKpljxLtEHxdOdcHKtsaWhOw99At
5qwCSDDbiy8fA2pEsG/+KsFzn3ksLGcWqvY2AyaMwORkG3Fh3fHmwgKdcQoqx/ic
Fy9zzlGNyobYDEbhSG1ZHzEgxTiSL0TpI8sXJhQ7Kp5MM9uh7FF6oNrZQEeXAJ2Z
tOYMeqUOorxrhBGS7QyQxOeZ0H77FfByPHR4HcOLFKQ1izUkuIRk/mpNtJhwRJKU
m3rA68Dumi5Ik9DQSfA4a/tx3/hewm1qxA2/tdMqHCKglnzW4gF8hkwDPYTVBxbM
Uaips+JFfAUjdlQ6yYCjDjjqbjdnUojTiEBfRhyXz1zxGFkONHM3IATQQeTxtz8Y
lMc/KN1q4BpgT2RFZRnMfmWV+2ElQ0tigu4ibuULlJUJiw4vkHBxWlA3essmnYGT
7SlNuEuVtvHIGUjbCLR4kIzT6ldLEhc63soMWZ9caaRntPiozTriLmoR8vjh6uXP
gyaVyc6YfHT0VdKsJI9ujKrFjDqmnW6Si2Icu0jZz/op7f+O1Iqp48thWjUPX1/1
tZmsb2ezQ/z8B0JSJ535N1voNuoYABNcfxdnAb07eWuQS7ay8u+7TSQi9gkiqk5U
RejlkPWnCzXe2q8g5vAtSoN8BfxSQHzn4fZSiShy7p8AJOSq/Mc2Dq4B+2nL+lj6
g9o+cMJb5wySpuQTUv4qUD5GywNs3VyVi//wxUt2cmL2rg1DF1kvWZxLW805YWDk
ufnUveP7qOugId/I5DTruz7cipShUKNwIZrEEhMoer+hCjvR1tGQazvykVHrjybK
YUWIDGCBradivhUh/jubX7XlSacjNRdMLv1I7r5r5uL8935GIze4cc4Tw1RaM3Yq
49K323GqRDzUhG1cay2lD8hlnFSLEkwXxLeK/aUlC+hRqPMg+e1u2EV/SkdwFTx3
RvO23i9bp9jWu+RdepBdMYUgJGIkXAHB3yIKX3p6Ap8/llSFNVU3ErPWqrDEA3Rv
1K+u03vdjsM0Es/NlI58BJkFzK5w5oqayAbEO1g1FVYmQsyfOxbePT8OEslHBWlq
QSr+73tmHNfSPTgtNB+iozOKotGGMGnA2lVuNqi1GuMRy+w9eGeuvaXBoVwZKSAG
dFEy61dCB75HmTUpkTbijLHsWfbA+Lc31ujy4IsZKfgWXaIdnAOS0FzcsSQdP0i1
bAt0lib+2feea2a07kej4ybvYmB8fq4u+aUflI0GnqO+FKdQfWy8MOPxZC54zM2r
MRnAx3ACPs480Yna3T8lWrQN5Wut2jnwV0XtthGsccPI+BchA+2iP72gb8JahqTT
8kp0QsjN89C9cR5UOnq/DlAQGUlDvwX082Fc+DV7P7veywr3orFBcYdCteGWpByQ
waWYXbAGdLoYj+bgN7S/XTiGeJVtb2u7A2e7BKiRjJRAxK+4+PMYd9FfGRceo7YL
Oucz9hsFA0MoRGHH9EbvOzuWuOK6K/eLcUuM4BoEWCx1M2mZLWM8i3DQY8PfbjCL
ZJH/o8svGPUwwqJ53YHVerlU0bZYhejBbZj4RLpd5+PdQd5qz3ryF0e2TLIo3mqb
GPgMHeyIkrT2gj14jNT5ywzCbSKg6XNA67sREFN5T2yDwyLuGHVcs2alZBMCZI4b
5+RASLM6WyRXULzU4A4DubsQTC6tSFFuXTdzmqbK37flQsN9MGefRsWPRxLI8R7L
YnUFs86OSGbaweqY49rfDD9Gj9OvSx9N1qrxjG5rJkHPpf38gfcBz046O95PLKNq
JTujRIm8fUhtXAv7+e7FQP1NqOmHSrBcd6ta4lJx8oMT5o/e28gZwFlo7nHzveQg
nmsssYqVVuLTny7UHIJYxB4jxqAnhAxkFNiXcwq2+c6fRJ3YvtPe0WXzHES9gJgy
WFQdWRJYXcpjBHdFwrRPgw2hUODvdESAwpsTv7pTvuRfC9XqMim74maRx3KHT+mt
AXZ09dcqFAHhl3/NeGj8XyaWoGKU/sVqXxXMVQvEKQjKMyZpA1nfC2eUFF39cNES
wLGTTpzESHtFVx37EGt9HattUR34KrfkI1ubO055zp6ObYVh62TUIXVtUa6boOVk
xgrrBkOlSWh+bYGzPTzJmUuXhkZRcdqlwMet+t8GbynrCfoZIe+MGBTpqYAhtRy1
AJIpkeHetqkZMXF48aZOMUa8ZZCqThjygJV1AgqZrZGYgU1U+J7AlDB9bl0XaUDC
adiU+gLSZBaXxUg+9M1nAg8s7nHfoR1gJFbPq2BMAPjO7YWKfwGfA0Iz8zrbBPkt
u8q/IkvAEaDeeoFDIJxlQ4DnWX1hgI+uAIAd3CMWs/LlXSUzkSQJ/l+g/SSodSVL
L/6yk+TTsrFUzvbZIUGgPnANxdzpv0iGNByROuO3IRgTTB5ohkz86TWEWVShkgKZ
6JyEKXDY5O9FxYKiYM2c8ygt6l0YT9/33M+OjaDeCbzoY4C15FW8cZzGQMpF7zen
VcxJ8h8ZU47/w4P2NJkJ+AU/9th6YYBsqLWb06sxpjbszNyap0Gfy5b6jg9dnIIK
jSW3edzaMQKqERHgmnr+tvP8JQwJoB+Gd0ztVsFfRAW0Ns8beZUrIFwnKNLc2baD
y35A/QuX0LUfcZxvVEQPgkd0sM9Lp70B5COe9Lr5RUGStw2hPnvo6Xc6mipQM4e5
WMoXLG7eZ9Vw+5PU1dpOqrYlP3JK26jlC/d8KPo+M4OML5sgKSQktwY0qtwJYXwL
VQhBp+iedPdnyV3qHan3seqAeGUK0nywLnxJNEMQ+KVqCKgjqtyzPFuuBEzTLYjd
Msn8wfRqBGKdDBfeE3GhTx+P+zBhbsUMQlvmfr45CNfsAt1+pK7z1TtFV+si7iay
UiEznrHqgG3kdRsNwligjm0RRjOBWdSAZxpw+L3fVCPXlfoWcXIq4hDtj+onlmz8
vL01fys7WNRhuA3yHLS15ku2SEP2t8OQPB51dKqfOdSNfxLcWXeFQzgK5BQSN+Jr
rEnAfv7f1URUPQb5OP8L9/3G1ES+2pzRIs237OKEduhjviW33hILF/ww9q+zHJNy
ZUOgKKMzehp0cVKHAevNujpMBxw7z8a6dicAFXLdNn5ZBCfQ92bqsPaa4Z+EIKQc
BnVvd4B644G279sCSI/ZzCsNxxh0PVpsVBuYdaKCeE8peAviG2FfgMUjYBk3ooZH
IewKmRs1fCoIwqB3kgdQDwcAWCN+7PGqzphKuINTowV1ZrhG8H4Xb4IABT4KnbIw
S8Dnb9NKLf1tLX+9eBlhPBo/AGBkH20vrDkBXAp4U90eiRshPGHPPR8mHY2jHXaY
tfWMFYb1P0ielWkkQAMByyuwglfw2bKtfzRsRXpz75m+Dc3wJfDKI3I3dcqa6foK
+VHIYnNYsQ4Gb9SebFBkK0A+HOiN/g+yZukkkarGJpBMxBHAGPMiDlDeWaA8pO5o
NyOZ+gYvOaNiZ8ogSP0B7vybBhr5tktuNk9Lx/5ZyiCeVoHgP9AYbufrru6z+Tr4
npgX7DkNUzlm28QMT8wKukjX3l3RNkRUddkbQVuWl33tBvbQtC/I78HGuZ3z6/O6
tq8dwmplTCgbd+RzEhCJ4b1n8rQYmtCd/91f6yt+fG/KERp80q01zbQQEF1U3lEj
QIeyTjEHfhj5gN10CMFnHz5UXQmPfBqrDPcu5B4xdYAh356CAEWTdtV78apMORiE
sFRiQ8ioDAl9cv7Gri3Julam81tPAIa66waNBcZj1nByR9HvMxdrC7AzRPhj1DeU
7expS+IDZaIAs90Agq/Z8e+2N0xERRKwLLdp18aW8PiCUy0T0SLRngVN60FD3emF
nq9g+30L+dfwfX0DTW1ajysB06CQIAgfFzbIPkjcY0E9VEFYxugdyRWDh2JyqL5h
D1/QYLiHhKWrqG+dlXvtrFmM23XpmRqGv2pazO3WsIRZMXr0aP7ElukhKMP5mdwL
CBZHfHyndK+dH8TJqzj8dYDULRsD5RQrANGmV5zZdJ0DcGaIBuCTYrEKknTzW6lh
dy/CFt9x0bdlSJajXxHwpv2jrLWyzQdsXl1OKP+xeynGA/jHX75dzDtqVbKa9XXw
ArvA2XC858wLqDF7/OjaEkw/AwjAPK4QJA9YeTOVNanpyX0bZfMQnKnszqkJTKd7
/GQVwLaSc3BiZbpDjxoICyOnepaPHVithV/BfidYMJQ=
`protect END_PROTECTED
