`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSW935ALRFkZ7ovyWUtqysTYDAYXhG0bUq5sCVuRc5rVeoBS6ciNX5OeJg5kYQWh
jr8jNiAtLzVCU2LXSofEQJd/soSwTu/o0mLnLPjXv8bsdxkpPiqqdqJRX7C/g8/+
ZaH/1uak2C9zNi1Pd/IeegL/OC1H3fhyJIr9+PcuElVGz+H0f4Lvojb80t7ceHAq
eK4uQHR/+hK1Q9kkhOOVVbo6swT8X3XiCPmI361na2YJ1mg1PYpZnq0poadcaokt
c1S/ss22FblNjOjopCYaufWLnhE/f4pO/pBShKUdbRKVOeuYg59MDFGyaui/XLtN
+PYMTLi7vJ8+9x2gHP+HnQg8J8rvJRSN8lJbnz/iQO5cHTvo9Z+P6jGBEF1seN96
/3yOTb1SEB3yeRbK9fv6HnM+2D5FH/8YE1MYPrKaPPp6kxd+c7nclDXFWL4NSwsJ
Y0jZJyuB8lgNj/ZJqBZDcwu5VaRC23lpbSN5DukWITnR59sar/bMrp00fovw/wGs
2cMDJzv0Nv74XDyVFn6+eCSF7tPFmWhTsbJvR/FV13z9X25FyMrdX7N4BrDPwqHr
k18m9qtOVO9OIzdHomxvp4BW2QOCr8f0cXxozzkWmJ75UtPafIoNT1aMraiQLK5H
+ofBkpuXgJOpMjJird65IyaQJWfYMH7YrkSbU7n2XYv5nbvKkItTQd4ZMPT1tO1H
Efk0nsMk3I48eoDKvJCOJZOT7OhMITLmp6aIWVdYe2rR0Btr0M4P7knAIO5QQ9uh
HOtQ5qY6dCRDqyQ8yBl5pqJ2qL92MuFvh9kJpnFoxE75dsrn1Or9jegH5hC7CYlO
xUeJ99uGWP0KbRcweMRPhD1HnYGPbeTzcYQda8KJiJmTMedQRdWEvg8OfQC85WYM
I2vbglqwiVFP/X1XzOFG6hJga1ZYv6KzEIE1gT/RAQF290/YqsNzIjoBAON3q3mL
KFIQcUIeTjqz5rQjPYIoekJM77AQktmGXVG+OI9qdd5mvrUe8zkw+vLG/d6E9Odb
SOSbiZLWBq06O2fofyqQs2860TtAgr6eBQhdw1IRqcfMurFUAo3DXYbJXnwdpCnU
F6cifx8rRsvOnjIlrZ12TCaP0kEptNFvAggYWjffEQaoifEaeGR9ndp9A2V5Xt4v
6TB+hhR2LpN+owBD9LcLyJiG6wxKWrdWubHuFOv+p5I86/TKh1yrll6z5abBxsbu
FKFXNufDziYnXu3dwpNPdYVC/U1YbFjoc/WwBGuQJ0eHgcTC+rOrOX2i6k+a1kwm
obDWGmPIu9GRo79i/Ix0BFLBFVl2iPh3sriR8YNQJLiLBDk8n+OyhtDAChF85i5s
HBLjG0TcWgMG/fDtnsj+aT2W9RhKi7zi2c5PaDi7mW+uRLorM+vRVNT7dIAieUMi
Mhm4lfk5fpJj7o+WVBWhbG4FR1S9jNFb7PBesdR3Ol92hAZwEl935q4lPFz/M7O2
quwjgh8zv7iHvL+kGvTJVFjYJosDbO/catM57Tg6cLm7RXs2+KPEubAueMRgfe22
GeQdPw3TJnsrRRvFhy3BB8FbiqbqoKYlnC2AmWKc5bydHI844QqhWNJyMrJmuZZs
p26BUHd5HDV96lm1H1kSNoXuDTGKp9ev89DNTvgP4p7wCAJgywd8eLdoqNwtdOYO
UktKFgx7tVQBRH4wN282Bc7ZIQzCcdLzM2ceLem+HvL9n/REIK2g1ty4BUwDoJRo
JKLvGvkh62jNDBeI9cOCvDeMUjnR/ezVbbEjcOkJE8xRC2cmPy5NWSAb2mBBKJLB
aCuy/b2/nawr6DLh1jJVXwETL2wjyueKXrzt05Cum3rl9TLV3pQ6NyedAQ3kDxOC
GEoMUg0e6Rm6eE4nuE8JI2aSeyk5gd9DK4TB7O9HPD/kQWPrGcg6nilB7LgCSwAL
dLoKKFxzvzoe6/FZlJZEnLGtJSq3zjZ814MijuKBc1CqAwuc7VUJ+4A1KmPxN5OY
Cu6aTdR6i0hWG0FSkloxQUFWI3NdtYE4FGEPTBmFNhbkxHvM3oKDD/iAQg9ZP6Xh
26fADTjezQo1NfMVGetw2/5obuuR7NumkZqxHZEkMXs69KKeo+ezwaBEgKAIsqDD
VRANroMMv+eBiXma46Ng79BNDqIGxJQA/wMM5zemBsbAGAcfPh1zXqjSk3w3tk24
scSh7vmm4+29iNpFzO8jhbDDVIALr5ezSBCBBwNFNjYHMzVSS+JJCO32BzX0TZf5
0ImaA/Ioy4ApXQbEj4fwWhoZhtENoIuzxVcbDC1Ll4GXouBTZPXNsA+bKrrjHp71
CIj6HkeWfwwAus+sO0UlmmRzwzxnVaiUhcTtFCDpYCmhlLnshCL1+n4p9U8vSxv4
YyP5mu4AAHRtgH3VybT+WKcGj0vwws8EPHpi82nQxkbNNdjyNJb7U++i6uSCNRmD
l5w6wfcE1wvRxstzWvXZDV7+34ydqez+U0nhjhn24RQOj3H6QE7Vv9l5C78ioqlv
lwdw/LaoYmHD8NV781almzB+jKYgXmJ8i3WAuaXpZk0hUzVZwFAnnbZEa/2ycYQ9
aB7Z6AktUQ8lvCg66SALPNEouKONWg8qf+2esZnO5JmuV0jjNmsYfFVt++sDpDs8
bQ6T4wQGNe923PaI1C3uOhuFwMZj/91DEpt4BbYF4mkbmtxJxzvQTddY517u4/D2
D/VPrq0k341ebcWZToSCZviWsY/uNX0qOYLfXdmxPUSn7z+y4yGEaa5/OtAaU5Ac
SAgueidjFlb5bU3379kyNBxpsZV8VdB8dAC/qHWertTfBxev6iHLHUgOB37ecwh7
Bxi2dOQ7bc9yJKbNDuQlqGV6v0jtxgWDdTlMnkqy0SgsKf0OzKv6BFlq8WrKmTwp
SpFBI/pDvLL5K1/+4pO8VcBTqg6pnhaEsXK3gLBPU+1IwIuuiPQZAKRXE6qYsuCE
7H9Fy8CtYJUZTAumy1bDojzJlfh6vXRQzx/VqJT2aGBgun9yxdhnMUqBW6nDdVMA
P8Dxa5Po7o0sK+s7IxxgaA74LJel1SgB184IkLt7RgU37rXD3iFtLPg195jSV75+
iqZd888Y/LgrTLvXGATvi10L1YSh/4QiqlUHLHvMRQwuPzkH3B/wj17DUtqEdIth
t005bU/TBhc8SG33WRkrmFUs+BgD5ydAj9H/PmYiugRmrycMATwPFNB1uakp507x
SXqxBeRVO6VrGXANAaHr0aj/SrQJxzjPZ7lvjKbwmlypKfUEJZUItu0yD8ktEU/2
Xn44RwJbtkShYoGDIn8x08/M1nvAuUkmXaeg+dmBo2j1dGtP4Q/1rOlrTWBWwHAa
XFkpClJyz3iDZ7RQSE0yE9USCokce7HmK/YBIfXwfF5eI96lINyZcu70uPKhZNFp
VRbid4f57vFhirlilgGumtVTDSKFmk9SxnEQ0FGaJ+k=
`protect END_PROTECTED
