`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eV2J8oJJvla2gIz11FZ6eSdBVlxjos6tyYgH4HraHjn+bkQVCoVbSb+HAApv8UI+
plZYLBKQQpWpVr4KD8nGIVqrGWYj8J0ppHHTb6m5e0fGd9Bb6X+f52CSgxeC/4EE
gD4Gey9Ieh6rk+8BjPZpSj04EyDU0oqoSOBz+BGT2B7RE6qEPiX6gXlP8+o1Fzpk
Ws5P3t3D/amCsizypmm38VNzcWYkzOouY5n1ARzwpb6rmlkWtytuDMXTN9Ckx7Kg
//A0O8Crz+D3hwune3PMZNjYWsl8FPsY930HHjLbIMbpa2YmYzM5UHgySoiOyCkO
ASiIN9mrtD4K3TNQtOPDZ4D5yVqNIwE1ipJLTI0fWoeXsxVKhh4gDdwHxFHQR2Aw
uSEXcZQOQzMp6MxYwNLJMWpa0UxNFV0JmKcwduWM8T5/bwhtNa59aExW+3Y8VG/W
xcvSESQMBtDV74frk79TqACJvx5oIxCRw+2TMVwE4ImPiWQoCL61t99WIXXMW/ZD
GFAkLfYROQK5VKmr+SeIjH7XKSQLOIOcVt6s43SDfsOYs/XBEQj/m9K6RuV3Kovh
DH2zmddeB4lN2Aul0xU2AN1At6vyAsYHzIJY/MMj1R51NnXn5zWXtltbIFAcbgUj
cC6ipRXxcGZcCVUynSs/qW8IZvy43RZQ8rsNzR4DU+Udji2ZtpDQxo2qbfcQvHRO
Je9PxhvDrEoocawKrb9x5FMq9xyey6pJUo6NukF5ASAd4XSGdg9mY9iM1mnqHV0r
oFMS2GarxRRPIKvoK1aiSq+0H/wDsPy1ovFT8laSDNEFjVAJSR/mUlg5IEqTjHCg
Kc4o+jFo0HsVwXsJveSaqPXgyFsHVmhZSpMhJjkApQZ880KFmRMwLQ2228fhGkjU
CKN4daTPFPvhO6Uz2N0gb/3RZOVvqCa75gxjwGzBBNwnSjA+HyCxEoF8dx3kJqpe
t/hVaPQBB4lfsSHd5IGcjzzKtBFXPAnklGpLqJLC5DkFfAKM7t7w3G41WRhd4UUA
bWucvWDTpwOUxqMAfLEB14urjEzDhG/iHXRO+bC/YYG+zxSqyaBBKF/bf+i5GVcm
T5TEMlVi/I9dZynxhpNkX6prRCgxbvbcXX8V2Cy/4vpVpgNGGRMMZ/vmbzBgGTZk
G4B9Hi23Nq0SjC3nTRugxpZ3p2Mb+AX3u8fzFu7fQ2zYeToqgVHEzo90968xNCW9
YGC24JMipvzg1BqbiQaEW3eS8/6NA7LULp7wxxkSplkfXlKmaZOTs5FDg9vWpvdZ
nfqCdebAz8NyiyRHPc/owF7bn4+FdpLUjVEbh84/YcGP5GiHQ81PhkJovExgOmdz
jBS27ciHuw8GJB9rsqQBj9/0doOLaO0++jxh4WQu4GFyLJ16gOKeoQupNLOCPz18
bO9Hn5rKxtSVvKsuZpPH+17dzxTPK767BxvkeiO0nV1ldqQEpITaQUCZP5TUz9gw
oFcRV1UR9i/9wDKp2RALbxmOoVi2Q113VEhUy6qOSvG7KRbAm/rrJAQIpacJFslm
CBSONLU9q4ldWsYYfe5AGINYu4eO4plzmZ6c2qWd7KiTPQIyiCzSRuOFznMzvcMo
PVE//awoUqeoJp/VJNnAmGW3lhC5IaKjPXfLHUSfkiHdaGqyaxwPU1JtJBlIc9t5
yk1Skej/KaC0SYGGVop8f7BdJOK0J3FUlKvZNoESo4ZhXg/qv2yL8hwGTq4MuRDG
JnGSNHVz9lPrqvkwURmhXN3U9B6r+Dy/ls7IL7yl2UVGd4UUNyypWh+W4USp5ccD
AOQouMp69UX9HAZ/vNzZ5K5ncVgS6nxA8pXJWsC05kEodNRGMNX7DbAGavjA6qj5
cP8tarbkGHqrXVujSyAuNDrgb+6jbjPQRT7NGuGGayLX8gLgi2welmbmlD7NFiuU
xltNehwYTxFwyBbR1wUV3E7GQUtWC57HaCyeJCPtW8bWpQH0gsBg45Sh/os47jTl
eR5afPTSLCg6ewkP2F7NA9SEO8/D17rCFxuFyD9jGe2Of+iFGJnfC8/WR3FY/R64
RwcDyJjSlDeDMost3fQOeCYmKuODxbcSvB2NUziISSYLONWzSsaJoU9Amkl+T9BG
rUSAETviFry1EDTos8ngs1hQ9yzTEN5swAHLAZXrWWtTwlZpnKOaKvNcx+q7Ynna
ItyldQ5q2g4t1QuZQpLe/oOIsQLLUjwIY5igz3fbqE6QAUGkPHmgHsCQbzi3Gj2t
FLSCNGgS3BmkfK2Lipdfu2hE5KV/ZhNOuXQ33mq+KB4gs5QfLHg4G6YwJ4v4UW/3
hhSpbt5AN5VTnpdidEhkFDMq7CIkjmMIDBo2QMlp7dGD3x+6mlOAE8ar63XnAj07
TSCcthYYBrrdA/wf64S7AdKI3O2MURu86UID5z0EkkYLq1j0gUXQk0igjB0aqZnf
CQTbn2PS+kxmn5Fv3lbHPaTgkJJa17IFzsz7ru12ox2WvKbSVk9TYWc7BKBDW9k8
mAXzFhZK4Tdt/sGpjPHemz9OhEt4SKXh6ji+2Ucpk/GMoiKJoI8YPej5x8xIsnVG
AXMxQ/Uz8QvWGNgUWEcJKkkXjAmwDN/ad0Seevtz66qQy1fi0IvJpHvuDQapHwJR
EBQsn289/5JhQDA+HuWi8xpZ1xX+IF/9qAzYnpZQeP/Low1GVWPAv2vkIY5ACfac
wu7xRf3L5zWLNOjXkzRYCGqF12a8HhhRkMJSUOJrZnjkZdv2Ge9wUeha9WK68EKX
VkdYVACn3iWHPqIW3sDRcJNFgwRlSZcFyrp8dvTCJSqwFKoNG+JStXGmeX12Jgci
OKXOffoTDqJKMtyxtAM/H8FyQ3/iFvcEvwvCpOGJ1jjWDttFsgk47/27HfxnfOcF
TchbrqtJnBA+XEgRTP+PQahtkHQHBsD4kMspD72uqh6s+H+ZkQKhEmQM2ecATXWs
xADCd9dlMlfaqhA5uTv7akusIE5p5Lj3+lQb+dACEOz99dKEIk3jHNsUmaIFcz3h
zN/kSnJlt5uX8v8jSWVXYTK7mNghcI+psF80YrD2PTL218bjj14qLZiKywYrGZih
btyxPwz7l1focLeppxH68hD94FeH+wLgohOp9m2dxON9cBy4bUqqCkoxivdZbUhG
06swAD1TbTuR9WLV4jpjoHP+6zj51fmKRn0X5bFCZsdoFVMA0VHL0foQURloTquj
ZSIEElt76f2ERl1Ia09qeKLxI3oCmDpMatiyQkmYIpbOKvNkg1BP5FogqYQSvLGy
uSUURBNIW/mmdEK9bQOH2+8myDR2VUqCtm9lkQF4pp6OE9fM1gxmJFdJiViPcACi
E6STdki5heLtjfoqGd0gccdZ97DKwgf1+53neNpqWVc=
`protect END_PROTECTED
