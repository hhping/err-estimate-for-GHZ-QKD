`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BmvbhXXQi40W5vBdEuQNPYFvfA1Kt51nXXENffiTbGDB1TKLYW5IaPeYctU93qrv
lx81MYgH7r2Cci0GJ35Ao1fqrwKJVfbjbK2QNhQgeqUhoJ24+h5IKD3ReSYTzExc
1fbIviiLuYo564fY9XB92LmqclrYretrqYcJBm9nqtztnP5JdndW1v9vFKqws34y
E3oKyxjP210Y9UV3HN09iANM50CSlSct/09uYoarl3W6zU61GimcADvBH881aL23
DCTLZu2kRf8z5BKqc7labrDv2CTPQSbHXcNCJL/yHGwkBQyWQwgv9Ji7AlIuqXbj
+Qh/P5AzY1AFgNYNSTbZy3pmkZRERNY6x6em3BLGQKgWmHvEUBp4paD3nb9779hr
ZfgGmX39FyGI5t4KsH0sNAWwCZOWjnA9E80SHEZLikrOpTRQnehSnOlECePbWMl4
oY8BqR6V84irH4+AiJgIrgbDgsPonc+qdeh0V/Ag26hwyHGRc6YeBfEuunoxFfD8
JQUb5MusRx1FXsWyz0aKkeaWLvj/76ktxxnRSr1LviH6NkzufFyVXS+Dw8s6Q9hJ
Xl4lxW5tx4EOTLhnhi1lmTnXP92kI/nEkvY4DwrP3/OhMRPa8M62mubaQybBRU4l
1RLThWgeYSAigYdD1ZeiccaRkZ7pL6mcks0RqyT3WCwzc6RfGnroxjj23UadBC9m
It2F0nMnlmlcZU3o67DaW9D5XcZLy+VCz6P7I8lZjt5CQZV5vOouXMTdaUq1MWMt
r+swQKHGfNaCaq3KVJc9ucbhDmhMkV0EMKduFJB7XYlGj8QvAxTV3VCE2I/+a9VW
BYnxDBO1RsDP1pcSsjsygvMWyay+OWcbhnuQYWHpEHbbtyfAlemzhnNGl9H3x3nX
u/CqNYbdbue1V/mieFp3J5wGcEAm95ra9c1iFj/KlhnTYkdGkIjBCOv9M89go7n5
iqKQ0ZI+4Xj+ZlSs3xwvL3VkHcj5VVAphyXaJ4sgzQgx2ijf31ktI5Cem35jgZxe
ixuNqxTZ3cWmxmuw3ov8X6uky0tjWOyVb21n4Hh214ESgSBoF2zbFm3ucYeNQRHQ
ozV3r4Lo6sm5OcLGOcWpR2Q0f3BqlWG1eE/eonkEAb752X6cjVyeCjOICh+iVzrk
MDXL8k/bfvx0Cronz4NuIPjRA/h1TYHzL3vZh1DhRfUGOHXDV+sgBHIUboR8mF2+
qgOQdOAdm0R1JaQkDBlNQTt7h22NNSO6XIb4p8HAKmKLYzPU60RV6MTSRtrnOJMc
0YW6IgiS9FiT5ktL+wbwCEo/2fUgkVxTqWIEs6K4asm6chCmW53gWkFm0dDa00QI
U43MLKPRJyzE2uAIjEpr2zxGUJ1TVUjottrwB2FFf9PM44nO2Lj7M9F1uKehXIXj
xBnlhl7ZJnfjMEqbiafOlH/zXSzESFZ/8PM8F3xkjN1sK1xgevhffZAt8gE76ayt
fEnrJ4ktB4cRnJeZYJWe4Q==
`protect END_PROTECTED
