`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0k/nVzHDS51kuQkU82TgTJuHpNfLJ0aIuphmeKxrD3cnh168BLiv6rdM8KHKoGv
22EQ5y/5DUbhItviD3yTjKQzDkPJeVXyrQ4bfc5SIc5RQNwtRLn5sa3zOeVdVFQl
MzLfkdwz272XaM9KUkU45elsPR3wnpyngTu9JiTsqDXeM07TDcLY9R7F/0Ywp5zq
YQ3t1lM066KCWFI+xvgHrpGH/Q3B/oxGrDJh+8xCJWUwYiXl7tR69kG+hZ/Lh9Qy
qP/2HAnqdvq4UDdIwZjj+iQE3/jos2+pGAKl5N7RcRAsajOUCLoUuZjpjUrrYyH3
UlKF9JrzqRA+4KzPGnofPrHhnaH3iuVVqmUSGBmmU8QCMl9M5dimVtXcOsHZ70wA
qH6UNLKZ4lh63Q2MhmpsNVFbneaykkegxwV/zK/JEZUCwXVwkdE0gUg7tjZBYYzn
sKfDyoQoabv9qGzyRw4JpGUpjNHSLttj+dPQj+UNJYbCFL3YgEyMN7Opm12aIPiB
5j4oYd6ZXuc7Gd67+y3+IltFHFHLoRMuYN9NwEY0Z65uuG1hD6Tix6PfdIbzIcvP
VcHrJhFSzlxET2Du/iFthKCna2lXc/1PVQEMc6ht03vNEIe5bV8tbBS5cMkAeZIg
0HfMmnXMxDW2+xK/A6a5VNwjGONZAvhLtJux/iQSTmCuRNyNJ6bacplk1yF04pB7
tbdIZQCv8y3LA42ld6fPzYW6dBiuOmCVEALFvjijPv7sprr64ijG6cywYDqlBs5Q
D1zzpUvgMsrnMzhAKmePjE6aV5wB7F7KeSivRqR5U1NLRQjQ+Y5glBXzMw3hlzDI
+ren7EJTVuaiWbZYG5SJGvszpSPdGxnf5LK17LfPTg4y1DoOc/ASu5BOelNgQB5C
o/DBJB+Zf9zLS5MQK8B/JDVuiVIOMh3xKcr1bldXRi4qIPeb8y2KNtDhuyMFO6Lj
mVfYSORxSxt+P2GxoV1u+3Fg4KpSFp8GpGCXWM0DhaiNjIxA2Ag7R+xmw5TLDTM2
HCDwuKMkbBCzi7wDkCLvudo3yXEVED0366SOYfFUI1Ij9ML+FEflH4gtBF3Mrue5
8u+rskTxP3FMJMFu/ilyigHz1NccWOxG1wBFINDJU8Iy8V+sKTY1FVNRpFxhfFwS
irLXs+vbFnRe6TJRSarslsYqctFlIAsu5nom0Te+SoraXqXzg0SZqxyEoHoILUaT
/BmFfy03nWpXy31nzkXFk1w93J64fY2EGLuipr7rxNHi2/PZfgf6t0G9vws26IlG
Ra5Cjif/hRDDzCEodFf4Aw01J3KnfbgtFKJYLXc4dlRIOmpreXxDCJkcLsS/jaAE
5P8bTNCyftShZkn3/1HVm2ZBkXMsh90T1k1G54WkdnUe4TyyNU3nSvGxjAIEMTE4
CzBp/FkNSrp9kVx7P7LIJYG3bM4m1gTAkhRGjmII1FwmNxQKjxswtmDRpXgvzD/2
F1HkEYbbyFGg1ayS7Q++W8mMFMiD2Qktjie5jiHcdwan7x3hSwSZSYLlQ3IwuYPU
qBoWtSrpjiZRH2LZuIjsx9h9Ib+tq/gpgVP61JYekobmoMPXQGt6thrLnCzOGDYI
lr8AbeMNubG/MLQ8+2/0uP5IrSbrTcMcbNWnCgfGd7KtNchBLhKJZjOpCP4Kgi97
trRx2/uTpwDQzeVBTlnnv/KMGURmvVnsiTIEtAxSCx0bMcV8aGdAYXL4//+v/j6o
LKSJKgABu2byFnKQRqQt7uSTD4C1+uOhguSQPfJMJDPprxCfOZ4G/6pDDmUHSjph
jsPbrf3GCLAGB+voyAXhJPdOz4hWxFVHC5KM1eKr31SYtjnOG4+3JZBh7k0ccon5
cFHQZQZHem52ZpHxtNGmVrlzjveAQ/+PIHTUZIBaDrIGAwwaKbZ2PQxZo/e1dLxp
2vAXUMnxa+DBmVmlL8nOhYfQGbV2IBorDzkHWq26s2zQsw5g3xDWZTrBiSFFPGoG
6e9IBj4CxkGo0As0tFk8w5m7BvVbBEW5iaZRd8VBW1+yFxrjvGENJIgaiqYKgruz
laRm0dUdfYlp6AZcdsxOzvdNtx9mMMVD4h6nlk4Z9/+DtfXpO3LSxd8O2IWgnqRZ
6GWLht28hcZVNO5qteTJyKqP35HHRNEjjthvFpAqkBml9iCZ9EksCYLFZy71MmSX
xaYiMmJ8n4eHLPWVihE+OjBcuw/HgoP4Gid4l5Osf7njLJENl0FI/Z5xJBaHdgI9
HI/ABL1HaDot3T4HTE38ixUIRJ3WA4wf06Pptq9lt4mex9JeURe5AJi4i2oezNpW
rMOP6OxAgZekm+QnVCakjMInHgVOzwLCB+DvrdQDMdRCBgXC+wUax5zRZ4WmtgYa
enoG1Ik+GpTNEpgVNdyQoLuqwdpMkvLB8N0pQch9tIPFhn7LjwNPxAq04BLjzsDl
eBokftOFEDFPL7OAwrm4dA+0WHN2sHw8R132jfI5I6ByvQxTjIPGzcY0pPKmXA9j
bLf+rVw9pbj0FfeFiYnNwGJ/D+fSXW3X7xQUKFXmRHK37kjl9g62EaXYc2hNmQUo
mbIqLyENH+Bb1mxO/pu4hP0n1vPikZymQ61b33uxVggMPYaAMZLtSxx6dBP+si3R
tmm/bGm7vSlNgP3n+UFx9h7rcsjyQdLBDOFHd0OmI4RQZ9EUZGOQSBwXBlADLGsU
lWDdj2hsf2bGft5nbIQ+kfrmAjOL6A8xAw8vZfwg2LzWqtKO4geAVqkTNxDSgNkj
Nbwl7IaLzKlVgZRK85dK6RQIob6vbdOklKikghBfXBh1wyjd9XB/9v7huIrTAnCx
Re8JpIcCdaZuqWqxOWg1PSSnfrfh3HNKPFUpcWZUgcT4jT16GhISeXAcrrRcksgV
Occ3vEW7LQEGuxBODhUqxKl0yb/KILe3/fEwA1qnRk5p/lhtw9fSziOC5Nv+YrZ5
CLqTI+kLFZm8V3ygWaS4/K8jlCNslBJ18kx36ezBg48C3bCO24sXDOP453BZqPx5
++hcjXt074zKAs7ElOGbod4oKqzleN0T5okleya+4hYM4pQjXD4zuuq6okyQKxc5
h1i6EVLiMo+yI0ajNtCp1bTw7iN1ZyynTL3oj1zQbD3LAWOJDZ/k4seRxMUUKAYv
sJxcZ+3JNIJNbeFtBmLU7rcsNgKpqtwKkr4sB6ENoF2kqUr6Vf3Svg8yvhpy52IQ
ddYh0ymBSR1m6lLeO3L2EQ==
`protect END_PROTECTED
