`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2meXKvR05Lm5RwTsAZvr8Y+WuA3GX11577zHZK7W+SG9rPjrtzP2O9kep72h2Kn
9WEKDqGq6YXblljJebNcEfScxikgb55COiNiuTNRkyt1vu2B7YkDSFc0JbJad5gj
vqrMGK/c3F60hIAB1QGqOhLZDrvo/3K6UEzgjUyNLxpz2f5Erjdu9eO7/4XmhZls
m7hG3a39tgCx0iY93tLLVjnGfT4Ndv8/JYj/WZwCQTEj0wZ1CgD9jcG5f/LPs2pw
KrDdgf0nmKbMJfWKHE6KKrH5mslkhjbR6WJJw4zb/j0Db07dSBkf4AeXDSKno31L
oCX63xlEzt4BmYvkYejIT/yXWCIExNZpCAQYKRUeTCH3bdg27bdo+IReff2KkcgX
HZYZf7pZvUUSh0i4nbWNmIRQoRwT1pRzis/JhoJZ5PCIYO0lB8ZFQHVZiJIKjvu4
jiW6Bgm29cXAYHcqidI167AZvLwxlPTh7/2LdXpXNrM1E2n4s90grgpXxWQHefUK
zEAuu/mJ3ujwLF/J0aG/tX9C1tJoX3hMHFrc6kz++3Pz82XGaBGwsvX71NdrZsdU
GzijmjwXs2v60aI1vlYtzPLsNQ3ECYbp6otT8ukF8zqSZFW7qQB/XB+IkFcSCdPZ
Ngega3BewB7jn+VW3sQHFStE3XKsesCSH8VfnQqePN7PiNrz6CGxTv41JgbCYkFD
HTN3VQ98g09xQoeB1oGkWtFJNsYrl4FwTKVaK60rY2yDactcFEEcqosHsIEIu9EF
05zR/VAVKtDa5L4RcCH7l/Kgb62v93DoZtfUSVAhLLUtzCAnvptEg4uXysSbiitg
qdmLYo9PChPVq48kqMPo/sFsrbQz/qha+isuRxHljuoaLPK4HCUdVCS4URNrWLLN
JuUli4z1R2PSkhY3yPUAjXl9XkxN1fSMZXX02Awj/0dccMJMcv+3U5V2vhW5gC6A
qQ41daD3QhghgGMV55J87V/T+ViGl2qZ+2cLHi8OLXh3IIK82IXHAlNwomQh601q
IuaIdLBiLBP5TBUCf6C5wc5dMgEWA8Ei77GUu2bZwBs8azfG/KCLEygZy70GFP2/
CftrU/7unihylEy5CpmL1jpB2mqN67N5NSKd+ErF7KBwSJbcfx6B8FcW4DT20Y5S
dgZE8XEqaQYNxwwq0HLG8KZhkX5hViQORwxgPSU/KL1/eWITphVA+bimz14CsJ6C
/+dEF+381L3pYe3Ix34y52IgjxVg5GitZpWTGNOO0ltOpLrqiirjlSjxueE4cTvo
5G3QOHa1hWGkFJp5m+MeLEPSSzayClyqMoYyJENoXtU3RTwXnFNO1mzqrN+zkbSM
DIBWbiCivum1IVg+rAH/6ruxt9BZmk4b0Rb8xH7To4a6HvK/6L2hO/t36VOli84I
Vk0nRhYB8Aijyn92ghby6tbQpH7qKj8gRD6E9GRwOvz9RTU1v7b0bjXKHb7ZFa5o
F+Mnh1sYP6K72zwJS0IzJ2XeOG4Y8yNzzoGz7yOBW18L3j+qiYsFPWHQuxsaP1wZ
wxRMAQrIi+LV5USTUuUYvraPEiXHFuujfjQCzLKhINTS7eZHHPvaRxts0e3rAgR8
zXzqElLfZBovnNky1xMFVo/tAcR6BP7MZmaJgu1+Ps5g3NR/xN9EPdN7A1AbSxCS
SFkd11nndXLw2AMOLoMWfuaQzzfIiIjkm1OCJwnOPKFtl9Y5Vau0TJv8AobiQALd
ahkawyue/8zFx/4yHlGjQ+BTVQjDMmpGCa5FmewH1Idx8twkby+dQHgswBY1Ypns
oDM5C+thVgabzU9gX6SwGEUbccL1erxnCsdsqrsnZVe/7vkT8FzJopLAGbkRiRVD
quzhGBKRI2jBsMoiAKUxrvVioMVp2caFyI2svbn/VQycQwPvRDa4yFIRoEUtRUui
3vEvbp6r1QjPh5wlVz2ggQ7gRDi3ZLYQA8sfqAwI9sG5n+CCfDL7p/U+kWV/5gM3
YqkpsvXBezglb/eaEN6cUYgbfqfjiqPvJGAhpVK/k+snLnu6+W44qd93OjfSxCQl
8AiS5iCafJrJElVx4t4Y1NmsRJv5+W/y8jHGvQiytlq9JnUDaR35fGKJ/jEnjXFW
RsU01YUBNpxlnLqL9kapa7ukK8+vbuZBBdMvQqXbx5A9RH59Rr3KM4LzEFqx/3ZQ
mDhQsOVFQOD9n7rlFMyjaPlFrjIRWchc9ZGiD9R1Q4R7N6XlqRSZg0nlrd3Eog7g
NIGybaXcj+6UhZ8+SIW8yCbPWG9dwBNm3qXP837TsMD1uOEHpaqVXrZUOOHG0Zmy
7ps4PJl4ZQaaUeDqJvENHjLT+vv3ZkT7S2/Gr8rXRYEa+dJ52EcJ10brEm2Foc7m
cnDM8CR/+x/nHwko3+FXj65rhhLC11noWO5S+5G8rVScpOlPM90v5ner0foiHmLS
UCFQyosJpuZYPfypNgRbnv+m5QzErpzUv6tqAzjvY5UcWCVFw1j2n0YtDWQegSEH
6veevFGTOMIc/ytt+ZsN8iLLxYBzYIwODYFH7yrVy60Siol7IOc7G7LhY4/quxT0
AqY+n850AEIPyGggmInl9aYQkUnoe/B5ED+5rODjFbVccwXu4OJHOhKzlX5fVqpq
CtxZRr6QMOwGATDUmN3iQ/UNaLy1UdewGgMd9w+lvS3wyYwcl+mpLGm5qqMWr/Zx
JrNyH1UEQ0Ru6PS36Opg/JGe5nY7SiyPWeuP+538kRNNooVok/DqzixXpbdnWaUj
wFsKkZVKISxoHkkWvtLj78Q/887mCrbYcAR/E6DLWW/f4yEfSw9VJ6TU5x6JDLiL
L8enB4NQ8TUlWMcNWYjvNX/7WJS6vPl0v4VieZFm//QaBcc5X7F+FicDg59Ag0wF
I+FpxWeMKseTOaa4KbKIopM9eOUd6LqEEzB8qD24MaTW5YRcr/XW9Yg5YqA9wlUf
blOehzUQgEmdX+S7/d92WmAKKQ8S2yUOyngPy+9F5FIOO5G1bjdXLWqxhcPn8jmp
535DqcnGMA7Jspz3MxPZps73A/19uObK5M/stf9/vi3p63gBWlM0fOiTni865Nub
x02nLPNbKUtiafaiPJPQASeMA5MsY5+OQ5yg3j2YirceECrDI16J1oci3ClBDQ9g
F44XdZXtBra9LmiX9CJv4PkxTRCKcjG90aPrzY+HwiQPFz0O7iFDGxFkL5sau8sV
`protect END_PROTECTED
