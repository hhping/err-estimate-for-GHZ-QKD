`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4qUnOK4Z+tU3vvNMLEU0K1U6NdVKD8o+nhvnqv/7KW4OQLq+sp4R/R5vGSC8Uyu
jpfMTTjtXjpdN1SGjiFrobrBurhEWZ2jJoIz1dn4X5HdbDlRwiwSRsdlbehQnyS3
NcTHQHrD2PK/Dd0M2O42sFdsL9TATTQKA+O49I4NLVuTAUmj58JYKJ4qT0Qlpx4r
2uSwnJVv5qxEcPttGLL2tcYqlQhjiVmct1J9LZgYWcFTvvNU2t7pWEAnJdaBuhSz
IeHhLnoO72W64lxD+3QRYxxH/HqZNkS0DkcrXpgN7GRWHJLXPj5CpvqB3+59zWbV
mUyooVzlxMWPGElyT3cSAncT1Rc2CSNb1/3QCiEjQcPw5bmnMNKX3JNSBpFYWPsY
721jb7jLQ8UogqcoeM6cMKjjhsfqX/6iBtlOIVs4mO45Bj/myMae+oYZU9Q2GHqe
G1C7fHGjs4xO30I1mifn8nZDTyAtvcBxLu0VeRcuNuRb9RNO00/bCLf1ZXxg7Cag
AdPXCi48VelOzWhvnIe/gBAyTUPTZbypVfvoLydYP3dDjHH1ADLgZK6VFKbh5vi5
aZXVzdmUkfkIVPJhINgMnBBLz/Nd83PL1pqjL/PWdpZ6HtMnHLRy/1keHgQhjT1/
8MAFvdsFWxKDjgPV/wemAQim3f2nGwLBhpYydyqlBAYAcGaknGUZtjxOqhTEffUP
cF3dQS3AKL8gjPO2RwpdQPfIs1Xx9ME96iWidSXA47yY5m4JDYdWiAceKlUKkWe+
`protect END_PROTECTED
