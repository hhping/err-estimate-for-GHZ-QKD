`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vAvhDlZD3NqCnRFhQu16dR1RFEOxzuz71wTnvVrB1pM0tJYvyjsiz/PyJcAYo48f
pQGEkhxucntseWUfneWp5JbQBJeAFVqAtTKJypDdqiu0MKxTz4wHTwo7LyMpU0yy
XzBYiQyiSk3siGfMtvoOnnjiPdISs6pQkQXHMHCxrz6+lW272XM1d+HCvjVMNKKV
GE7ZCYKzXGCNprNzgpE99gbv5Y9YCOz1pOLV5JcGTpKNuVmvagfhl8TnKp/4qMxx
P8PAwEMmTNA1cAX7PLmIdYvNGR/nunMnK3TA+PbEGoAiIf49bfDQEdy2GOH6XqNX
FtHfNKsn99PVq+7i440HIPWh0QMRA7xbKTF8kUNag9nhz0X6rLOR9pXH3/fyIS7N
LXPLSCosoVo1eZVkJhykbrm69ivrjYs4JBT6hcUcIBoPuqja/lt1ArQeHOZbr1uI
kqEQZu+4lOGsefkn2vSkhUJu8iIoHmOZVjlnaAVfbq4=
`protect END_PROTECTED
