`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIRw3uqi9yYyTpr5EtqZaHIyZ3cOIMT8ISDvsIuwMwDehVVwoLMfNjwM9HpFJ/0c
hcWrirpQHv9XLsx2hcLtl9dyn93mYqw/zT4eZBWRO9jyMutDbkp3bagHTzJiV5It
5EVJO3TGb7vz8THp/TaVZIbL9j+pYv7XsY6BrLloFLfzKVXZoTVdvtwgdiVu145L
WXUd1A8x9FFcdrrfB6wM1UP+c3EBtYL5fjcyVt2WuMQFCFG9FVOIcI9b7wR9zYu+
TwXiPaNqT2xYr0cEPIrQ4Xq+IPn3Cd5oWtoNxxEdlDazumWQJVYUs4QOGkdDJq2Q
f/rBZ59nE54h1TKC3HMp80qdRo3cYte7WlwwYL4OGVehYhef7MLcXsXSl2rfX0IY
oofoJiiCwi3/HaFId4Us/tbmH8ArtGbzIoRyC4zNuQbK30etzZsgqyuZ02MH5imn
KpCRTLzTiOsoDU3P2JQPHnrg4KVGwK+yfxB2zKEVaNLDaacFeMq5hzNRg07V6Uqv
BenvDJ5u0uXOpe5fuRtu+soE8Kvy4SvmdLOYEWPSdTooP0G/FGaOkjvI2LcIOlg/
N6R9VdkBvxe62w68YHm1CLXNi54Xo7+l0jUKKUlOe6g2Dx0OvBpMOt+UYRinIw22
TxZw+HNN6Ipydx5jB3wvEE/PePhVY5sooVPEVlk7SMar3AvYVMyu35lbK9vYpvcW
OC/XbJJQaB21mNsyMamH8Q==
`protect END_PROTECTED
