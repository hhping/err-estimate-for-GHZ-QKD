library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_10g_rx_pcs is
    generic(
        enable_debug_info: string  := "true";
        advanced_user_mode: string  := "disable";
        align_del       : string  := "align_del_en";
        ber_bit_err_total_cnt: string  := "bit_err_total_cnt_10g";
        ber_clken       : string  := "ber_clk_dis";
        ber_xus_timer_window: vl_logic_vector(0 to 20) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        bitslip_mode    : string  := "bitslip_dis";
        blksync_bitslip_type: string  := "bitslip_comb";
        blksync_bitslip_wait_cnt: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        blksync_bitslip_wait_type: string  := "bitslip_match";
        blksync_bypass  : string  := "blksync_bypass_dis";
        blksync_clken   : string  := "blksync_clk_dis";
        blksync_enum_invalid_sh_cnt: string  := "enum_invalid_sh_cnt_10g";
        blksync_knum_sh_cnt_postlock: string  := "knum_sh_cnt_postlock_10g";
        blksync_knum_sh_cnt_prelock: string  := "knum_sh_cnt_prelock_10g";
        blksync_pipeln  : string  := "blksync_pipeln_dis";
        clr_errblk_cnt_en: string  := "disable";
        control_del     : string  := "control_del_all";
        crcchk_bypass   : string  := "crcchk_bypass_dis";
        crcchk_clken    : string  := "crcchk_clk_dis";
        crcchk_inv      : string  := "crcchk_inv_dis";
        crcchk_pipeln   : string  := "crcchk_pipeln_dis";
        crcflag_pipeln  : string  := "crcflag_pipeln_dis";
        ctrl_bit_reverse: string  := "ctrl_bit_reverse_dis";
        data_bit_reverse: string  := "data_bit_reverse_dis";
        dec64b66b_clken : string  := "dec64b66b_clk_dis";
        dec_64b66b_rxsm_bypass: string  := "dec_64b66b_rxsm_bypass_dis";
        descrm_bypass   : string  := "descrm_bypass_en";
        descrm_clken    : string  := "descrm_clk_dis";
        descrm_mode     : string  := "async";
        descrm_pipeln   : string  := "enable";
        dft_clk_out_sel : string  := "rx_master_clk";
        dis_signal_ok   : string  := "dis_signal_ok_dis";
        dispchk_bypass  : string  := "dispchk_bypass_dis";
        empty_flag_type : string  := "empty_rd_side";
        fast_path       : string  := "fast_path_dis";
        fec_clken       : string  := "fec_clk_dis";
        fec_enable      : string  := "fec_dis";
        fifo_double_read: string  := "fifo_double_read_dis";
        fifo_stop_rd    : string  := "n_rd_empty";
        fifo_stop_wr    : string  := "n_wr_full";
        force_align     : string  := "force_align_dis";
        frmsync_bypass  : string  := "frmsync_bypass_dis";
        frmsync_clken   : string  := "frmsync_clk_dis";
        frmsync_enum_scrm: string  := "enum_scrm_default";
        frmsync_enum_sync: string  := "enum_sync_default";
        frmsync_flag_type: string  := "all_framing_words";
        frmsync_knum_sync: string  := "knum_sync_default";
        frmsync_mfrm_length: vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        frmsync_pipeln  : string  := "frmsync_pipeln_dis";
        full_flag_type  : string  := "full_wr_side";
        gb_rx_idwidth   : string  := "width_32";
        gb_rx_odwidth   : string  := "width_66";
        gbexp_clken     : string  := "gbexp_clk_dis";
        low_latency_en  : string  := "enable";
        lpbk_mode       : string  := "lpbk_dis";
        master_clk_sel  : string  := "master_rx_pma_clk";
        pempty_flag_type: string  := "pempty_rd_side";
        pfull_flag_type : string  := "pfull_wr_side";
        phcomp_rd_del   : string  := "phcomp_rd_del2";
        pld_if_type     : string  := "fifo";
        prot_mode       : string  := "disable_mode";
        rand_clken      : string  := "rand_clk_dis";
        rd_clk_sel      : string  := "rd_rx_pma_clk";
        rdfifo_clken    : string  := "rdfifo_clk_dis";
        reconfig_settings: string  := "{}";
        rx_fifo_write_ctrl: string  := "blklock_stops";
        rx_scrm_width   : string  := "bit64";
        rx_sh_location  : string  := "lsb";
        rx_signal_ok_sel: string  := "synchronized_ver";
        rx_sm_bypass    : string  := "rx_sm_bypass_dis";
        rx_sm_hiber     : string  := "rx_sm_hiber_en";
        rx_sm_pipeln    : string  := "rx_sm_pipeln_dis";
        rx_testbus_sel  : string  := "crc32_chk_testbus1";
        rx_true_b2b     : string  := "b2b";
        rxfifo_empty    : string  := "empty_default";
        rxfifo_full     : string  := "full_default";
        rxfifo_mode     : string  := "phase_comp";
        rxfifo_pempty   : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        rxfifo_pfull    : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        silicon_rev     : string  := "20nm5es";
        stretch_num_stages: string  := "zero_stage";
        sup_mode        : string  := "user_mode";
        test_mode       : string  := "test_off";
        wrfifo_clken    : string  := "wrfifo_clk_dis"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        krfec_refclk_dig: in     vl_logic;
        r_rx_diag_word  : in     vl_logic_vector(63 downto 0);
        r_rx_scrm_word  : in     vl_logic_vector(63 downto 0);
        r_rx_skip_word  : in     vl_logic_vector(63 downto 0);
        r_rx_sync_word  : in     vl_logic_vector(63 downto 0);
        refclk_dig      : in     vl_logic;
        rx_align_clr    : in     vl_logic;
        rx_bitslip      : in     vl_logic;
        rx_clr_ber_count: in     vl_logic;
        rx_clr_errblk_cnt: in     vl_logic;
        rx_control_fb   : in     vl_logic_vector(19 downto 0);
        rx_control_in_krfec: in     vl_logic_vector(9 downto 0);
        rx_data_fb      : in     vl_logic_vector(127 downto 0);
        rx_data_in_krfec: in     vl_logic_vector(63 downto 0);
        rx_data_valid_fb: in     vl_logic;
        rx_data_valid_in_krfec: in     vl_logic;
        rx_fifo_rd_data : in     vl_logic_vector(73 downto 0);
        rx_fifo_rd_data_dw: in     vl_logic_vector(73 downto 0);
        rx_pld_clk      : in     vl_logic;
        rx_pld_rst_n    : in     vl_logic;
        rx_pma_clk      : in     vl_logic;
        rx_pma_data     : in     vl_logic_vector(63 downto 0);
        rx_prbs_err_clr : in     vl_logic;
        rx_rd_en        : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        signal_ok       : in     vl_logic;
        signal_ok_krfec : in     vl_logic;
        tx_pma_clk      : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        pld_10g_krfec_rx_blk_lock_10g_reg: out    vl_logic;
        pld_10g_krfec_rx_blk_lock_10g_txclk_reg: out    vl_logic;
        pld_10g_krfec_rx_clr_errblk_cnt_reg: out    vl_logic;
        pld_10g_krfec_rx_clr_errblk_cnt_txclk_reg: out    vl_logic;
        pld_10g_krfec_rx_diag_data_status_10g_reg: out    vl_logic;
        pld_10g_krfec_rx_diag_data_status_10g_txclk_reg: out    vl_logic;
        pld_10g_krfec_rx_frame_10g_reg: out    vl_logic;
        pld_10g_krfec_rx_frame_10g_txclk_reg: out    vl_logic;
        pld_10g_krfec_rx_pld_rst_n_fifo: out    vl_logic;
        pld_10g_krfec_rx_pld_rst_n_reg: out    vl_logic;
        pld_10g_krfec_rx_pld_rst_n_txclk_reg: out    vl_logic;
        pld_10g_rx_align_clr_fifo: out    vl_logic;
        pld_10g_rx_align_clr_reg: out    vl_logic;
        pld_10g_rx_align_clr_txclk_reg: out    vl_logic;
        pld_10g_rx_align_val_fifo: out    vl_logic;
        pld_10g_rx_align_val_reg: out    vl_logic;
        pld_10g_rx_align_val_txclk_reg: out    vl_logic;
        pld_10g_rx_clr_ber_count_reg: out    vl_logic;
        pld_10g_rx_clr_ber_count_txclk_reg: out    vl_logic;
        pld_10g_rx_crc32_err_reg: out    vl_logic;
        pld_10g_rx_crc32_err_txclk_reg: out    vl_logic;
        pld_10g_rx_data_valid_10g_reg: out    vl_logic;
        pld_10g_rx_data_valid_fifo: out    vl_logic;
        pld_10g_rx_data_valid_pcsdirect_reg: out    vl_logic;
        pld_10g_rx_data_valid_txclk_reg: out    vl_logic;
        pld_10g_rx_empty_fifo: out    vl_logic;
        pld_10g_rx_fifo_del_reg: out    vl_logic;
        pld_10g_rx_fifo_del_txclk_reg: out    vl_logic;
        pld_10g_rx_fifo_insert_fifo: out    vl_logic;
        pld_10g_rx_fifo_num_reg: out    vl_logic;
        pld_10g_rx_fifo_num_txclk_reg: out    vl_logic;
        pld_10g_rx_frame_lock_reg: out    vl_logic;
        pld_10g_rx_frame_lock_txclk_reg: out    vl_logic;
        pld_10g_rx_hi_ber_reg: out    vl_logic;
        pld_10g_rx_hi_ber_txclk_reg: out    vl_logic;
        pld_10g_rx_oflw_err_reg: out    vl_logic;
        pld_10g_rx_oflw_err_txclk_reg: out    vl_logic;
        pld_10g_rx_pempty_fifo: out    vl_logic;
        pld_10g_rx_pfull_reg: out    vl_logic;
        pld_10g_rx_pfull_txclk_reg: out    vl_logic;
        pld_10g_rx_rd_en_fifo: out    vl_logic;
        pld_pcs_rx_clk_out_10g_txclk_wire: out    vl_logic;
        pld_pcs_rx_clk_out_10g_wire: out    vl_logic;
        pld_rx_control_10g_reg: out    vl_logic;
        pld_rx_control_10g_txclk_reg: out    vl_logic;
        pld_rx_data_10g_reg: out    vl_logic;
        pld_rx_data_10g_txclk_reg: out    vl_logic;
        pld_rx_prbs_err_10g_txclk_reg: out    vl_logic;
        pld_rx_prbs_err_clr_10g_txclk_reg: out    vl_logic;
        rx_align_val    : out    vl_logic;
        rx_blk_lock     : out    vl_logic;
        rx_clk_out      : out    vl_logic;
        rx_clk_out_pld_if: out    vl_logic;
        rx_control      : out    vl_logic_vector(19 downto 0);
        rx_crc32_err    : out    vl_logic;
        rx_data         : out    vl_logic_vector(127 downto 0);
        rx_data_valid   : out    vl_logic;
        rx_dft_clk_out  : out    vl_logic;
        rx_diag_status  : out    vl_logic_vector(1 downto 0);
        rx_empty        : out    vl_logic;
        rx_fec_clk      : out    vl_logic;
        rx_fifo_del     : out    vl_logic;
        rx_fifo_insert  : out    vl_logic;
        rx_fifo_num     : out    vl_logic_vector(4 downto 0);
        rx_fifo_rd_ptr  : out    vl_logic_vector(31 downto 0);
        rx_fifo_rd_ptr2 : out    vl_logic_vector(31 downto 0);
        rx_fifo_wr_clk  : out    vl_logic;
        rx_fifo_wr_data : out    vl_logic_vector(73 downto 0);
        rx_fifo_wr_en   : out    vl_logic;
        rx_fifo_wr_ptr  : out    vl_logic_vector(31 downto 0);
        rx_fifo_wr_rst_n: out    vl_logic;
        rx_frame_lock   : out    vl_logic;
        rx_hi_ber       : out    vl_logic;
        rx_master_clk   : out    vl_logic;
        rx_master_clk_rst_n: out    vl_logic;
        rx_oflw_err     : out    vl_logic;
        rx_pempty       : out    vl_logic;
        rx_pfull        : out    vl_logic;
        rx_random_err   : out    vl_logic;
        rx_rx_frame     : out    vl_logic;
        rx_test_data    : out    vl_logic_vector(19 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of advanced_user_mode : constant is 1;
    attribute mti_svvh_generic_type of align_del : constant is 1;
    attribute mti_svvh_generic_type of ber_bit_err_total_cnt : constant is 1;
    attribute mti_svvh_generic_type of ber_clken : constant is 1;
    attribute mti_svvh_generic_type of ber_xus_timer_window : constant is 1;
    attribute mti_svvh_generic_type of bitslip_mode : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_type : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_wait_cnt : constant is 1;
    attribute mti_svvh_generic_type of blksync_bitslip_wait_type : constant is 1;
    attribute mti_svvh_generic_type of blksync_bypass : constant is 1;
    attribute mti_svvh_generic_type of blksync_clken : constant is 1;
    attribute mti_svvh_generic_type of blksync_enum_invalid_sh_cnt : constant is 1;
    attribute mti_svvh_generic_type of blksync_knum_sh_cnt_postlock : constant is 1;
    attribute mti_svvh_generic_type of blksync_knum_sh_cnt_prelock : constant is 1;
    attribute mti_svvh_generic_type of blksync_pipeln : constant is 1;
    attribute mti_svvh_generic_type of clr_errblk_cnt_en : constant is 1;
    attribute mti_svvh_generic_type of control_del : constant is 1;
    attribute mti_svvh_generic_type of crcchk_bypass : constant is 1;
    attribute mti_svvh_generic_type of crcchk_clken : constant is 1;
    attribute mti_svvh_generic_type of crcchk_inv : constant is 1;
    attribute mti_svvh_generic_type of crcchk_pipeln : constant is 1;
    attribute mti_svvh_generic_type of crcflag_pipeln : constant is 1;
    attribute mti_svvh_generic_type of ctrl_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of data_bit_reverse : constant is 1;
    attribute mti_svvh_generic_type of dec64b66b_clken : constant is 1;
    attribute mti_svvh_generic_type of dec_64b66b_rxsm_bypass : constant is 1;
    attribute mti_svvh_generic_type of descrm_bypass : constant is 1;
    attribute mti_svvh_generic_type of descrm_clken : constant is 1;
    attribute mti_svvh_generic_type of descrm_mode : constant is 1;
    attribute mti_svvh_generic_type of descrm_pipeln : constant is 1;
    attribute mti_svvh_generic_type of dft_clk_out_sel : constant is 1;
    attribute mti_svvh_generic_type of dis_signal_ok : constant is 1;
    attribute mti_svvh_generic_type of dispchk_bypass : constant is 1;
    attribute mti_svvh_generic_type of empty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of fast_path : constant is 1;
    attribute mti_svvh_generic_type of fec_clken : constant is 1;
    attribute mti_svvh_generic_type of fec_enable : constant is 1;
    attribute mti_svvh_generic_type of fifo_double_read : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_rd : constant is 1;
    attribute mti_svvh_generic_type of fifo_stop_wr : constant is 1;
    attribute mti_svvh_generic_type of force_align : constant is 1;
    attribute mti_svvh_generic_type of frmsync_bypass : constant is 1;
    attribute mti_svvh_generic_type of frmsync_clken : constant is 1;
    attribute mti_svvh_generic_type of frmsync_enum_scrm : constant is 1;
    attribute mti_svvh_generic_type of frmsync_enum_sync : constant is 1;
    attribute mti_svvh_generic_type of frmsync_flag_type : constant is 1;
    attribute mti_svvh_generic_type of frmsync_knum_sync : constant is 1;
    attribute mti_svvh_generic_type of frmsync_mfrm_length : constant is 1;
    attribute mti_svvh_generic_type of frmsync_pipeln : constant is 1;
    attribute mti_svvh_generic_type of full_flag_type : constant is 1;
    attribute mti_svvh_generic_type of gb_rx_idwidth : constant is 1;
    attribute mti_svvh_generic_type of gb_rx_odwidth : constant is 1;
    attribute mti_svvh_generic_type of gbexp_clken : constant is 1;
    attribute mti_svvh_generic_type of low_latency_en : constant is 1;
    attribute mti_svvh_generic_type of lpbk_mode : constant is 1;
    attribute mti_svvh_generic_type of master_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of pempty_flag_type : constant is 1;
    attribute mti_svvh_generic_type of pfull_flag_type : constant is 1;
    attribute mti_svvh_generic_type of phcomp_rd_del : constant is 1;
    attribute mti_svvh_generic_type of pld_if_type : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of rand_clken : constant is 1;
    attribute mti_svvh_generic_type of rd_clk_sel : constant is 1;
    attribute mti_svvh_generic_type of rdfifo_clken : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of rx_fifo_write_ctrl : constant is 1;
    attribute mti_svvh_generic_type of rx_scrm_width : constant is 1;
    attribute mti_svvh_generic_type of rx_sh_location : constant is 1;
    attribute mti_svvh_generic_type of rx_signal_ok_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_sm_bypass : constant is 1;
    attribute mti_svvh_generic_type of rx_sm_hiber : constant is 1;
    attribute mti_svvh_generic_type of rx_sm_pipeln : constant is 1;
    attribute mti_svvh_generic_type of rx_testbus_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_true_b2b : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_empty : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_full : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_mode : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_pempty : constant is 1;
    attribute mti_svvh_generic_type of rxfifo_pfull : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of stretch_num_stages : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of test_mode : constant is 1;
    attribute mti_svvh_generic_type of wrfifo_clken : constant is 1;
end twentynm_hssi_10g_rx_pcs;
