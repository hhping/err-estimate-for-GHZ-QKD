`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJOKTNzdb6dwscRptEDqbcn88egMjFbnUZbz1icg42Z2rBwWslwXK4W5juLbB/OH
8cL92YwHyswOYn45w9wmQ8qjytGuBIVfFFv/b6XAkOVdbvVn8gc7nh1tGNHsloux
celnj/fJT8/OMR9DLU2d2zvWUpiPRJmAxXDDLDOTFobSgPvQILomLg3/xbk2L4Q3
r9khw704JkznBAyX2ODJ6nKL1J7J6tUikylOc5Wu0dfvMddrLKJrEUy09cIakB86
tKj7V1xgSEyqOiYJ31ypcKdsAmEZWw+JgXQLDxfGXmMJwsjrmeNpw+1y0ytiZeic
JkGHyPYLf+50nvKFOnS7sT38+yMvpZtU671cVrMe7+oL1Iks8KX5l4vX1ZfaxZIC
dGFxYz0F6T27G/5iTKSIVig3q1T3MpmsXlAYKxXrNHEuVIfHEPSLwDso8i8ceU2F
7r4TXCHYBer0Qb77G7Qh46/iiTRtvCOXiHkcS+A8wCOcVMnD2SAFFEZxI2wpSP6P
p6tePy8Wzou0A0aEYy1sg1BLV+xyuebh1gicneOs+FC4q7YxjHYBDV3ocC9HnIxz
882cIel9Bduj/HFhpg/gX3vW1frzTU3fdDGQy/xzFQtisTNZRlzpBLEY59hUKhkU
EanUVwEsMGTBgC8gTpy7u82vccck23TNk1vQLEv7N2MAUZbHl2QO296Z2HebAGl3
LaPCU5bx1ZgGw4JuAtxQPM5tTTdJLJ5S1U8GoYhHzFGAl7waijYCBABU74cSwT8x
KsZI1MyjlYYGxL1FNsRh7BgxnSX8KQ4otWv6qziBiPG1TDkjbHxqrmOiBVFJszW6
cODUu8Y/xeYWp9RBHdsU6AOKG8NLSgtZoQnt7thvfmMFDSaElNO+6FQ9OHho1H3c
IgJAuqG0vU67sFd8QEK1zLjsY8M9/CrDQsH0Rd8OFgS8oTM6OvU73FjtckIX51xg
JbelmVTvsvg+FzVD2ZR5JcDYD/0pim24dfyMr7usNFk=
`protect END_PROTECTED
