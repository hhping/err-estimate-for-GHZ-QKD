`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v3d0gb3xhv0p+nQA5dnH55cV+4UjTgNgIh5gGFK9IQZgw7O6Qr/NoTMBgmpj/0KX
u6UwWbKK4w9sxjw6T6+heUYUNHtGwMGxEaMAMpCAj3aSg1OcdE7b52dDCLePZLBp
GcAIHcigH3Inl4TGZvBvvfU5GSJBS+6YPkE4PUgiHesKqack0npxuFmqVXr5kjQV
hFuicL5ukf4j8Av6cBIKZPJdxv8oAAQ/EcLHzTfBrlb3Go3rX7JBhlYjnH7ZhHEE
M4YUKGHq/k6j0Sdrpqjl3ObVkl1SQMb7Kk2W1yCaPOWBJIFMlCXvAKXnuVbYsxaw
zr7ylp2FWfIToAPgYe2VBJ9LVsfqCWYp0wy6IJgxYwOPW4cZOsAaOIsj/Ps6eP20
U1tfwi8dCo+PyRowWDakrJbLoiC9751jlZgJzIm9dJrnFeAGkWLn3wqdQr7Hz7Dx
eWFAozMjz1D4221bhqxFj9yZcuKhU4a9X3a6rgfeKGuREPumxceZXRo5wsyvp97z
qcMchu7Wss5UCZr4TcqjNK0oUDlMe1VBBPIJrXDVrJI6m7ch6ud0hdd5cMrQmz5O
`protect END_PROTECTED
