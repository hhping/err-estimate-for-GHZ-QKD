`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BwAipYQBdu8Nrr8VaL1Rlq4XIW+FTlMrKZUw1yo69FCNI3lw6a6A3hyv7pxu1C5
q8ACLwgHB+9ubOtfLJGuTod1FRPwsog3eT4KeFScTTGneruGqZP3mxVFZmovxO+M
QgaWy4f1XDFkn9+FYXkIEc/9yv77EIjanr4wibuDwZIacbrpUPt4nsKp/Sx15qyY
pxjH8ZYyHj7yhAUwM5IBVSlHcT1RTXdws8OfmazprMzm9rY+7Xh2b7ljQJmZ+2d3
LqBkQFat89napwFgEyN3QjWL0i/cePXrHwQekEPE6S1FFeQuv7LmNE5ltsI5YISL
MOL/qxA/52TvY7AqMr9X5PmzfRP613Ml0eRD9YaIV+LM8OTozCqnELL+3PvT2OW9
rpQ++wgdP7AtUvvOPzXTbhxy49v+OMn86cix7MMH78detEbpbX0Vj2G/txQ8ljHm
UxiqqvZ8vs/M0sbNIklDsbKawrVlfIT5L45xwQbTh7VTWb6ppk5cXECdy8Ntv0Zn
dIWzOqCetItDdjO1TplaDDLoDKmW8PaMAF6CoCrRygEUm7VerXl30xX7zdCavXnj
EN/8fEM3NdFRIXSSI3SAjknHLBv+CEHBlyCgpr8PCys315xf2n6VOyR6I/Rzgtpf
A5ZlEHJvgWbudAjcZJTtvVXE8A2WG5c9v+MZJ9D/wn+ed6p99gPtPBJnpqCYX57U
PVSpH0k9ka4YcAmDRb5DKlh9JqhltHyJpVGo5V3vaG282RFEWtK4gb29Jj6lfudJ
TNNfKAZBhE8TtjLuLtazXtnm2WmcsgYh4fOXuVTDgq1OEZB4JtMi8Ur7807fUuaK
`protect END_PROTECTED
