`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBjiLzCUHX2AQOe+IRvJPJUMZRAx22ak6JargFJh4klH5hNumJK0LnrN7ZAOr+m9
3bNrODZQeXpT+h+q0jP+8tD6KPuknmJ+b4hrgr0hGaY2e3wpg9HPqC5DzqKVQLwa
x7+yh0B76vRSpfXrqBvFHprKc0YMxb23pHU/qtinv360Rym/Rv7rqV6RBBy0q28F
UP+qg8de+Pstif/R53XBwBzpZh4rcx3+mcbBtpquSLaBMQAce/AOhU556BTwSn8g
5IOoUt1Qzv46PXbAyrwfnzGXpIa9T+a5pPVyc8OnhHCcxpLlHX+M0fwQSQlkgiMb
s7BB+y/vkFNxKNTdcoZQIlUo0ih8MRHCKyO07GI50jcx/OMh9IVQemVI02wnpjth
Rvz+3+KVctBtGOpO9BkFWbhFvJtXoO6E9cUCDBLZP4CjBeADUBtyEXrAkq6wX+OH
BYiQTafMylvXY2ZrCZrCb47+IcJrIA7FeQ3JE/DaOq52EKdQlDEwxMezpg3PTc31
MvpjAW/qExbn/r9fD5F5/l/SkFiF6mVcxx3dwC3GEJ3Px0WsiWwPNvBli3bIt//h
UTxgGWjCQwdzE1Hfq5OGMRgSlGKnK7D8i7cRGFGV89hY7taOMmDS0VP0r6jhcEUb
8pOfYXwuA+sVMcbvwymP/AErwKTpKqgZjFdn/6PlFH75tgS4wK7G8TDtWaYISfQH
shrb/ezRUYsgoh7xfb0/sLGJMMxyzR+UtJpDHfNvkjd83xouCOu6orYAMHSfj5A0
cA3iRZti2AG4LGcFWvF9cv8ACJlom1qDGoq76+eJ+fX9I2duSef2TTa+zPwGxKq8
AQ84JWnbJxmpTxTnSi/UTuuaoRBMkZRgbaJKyPGbScsp22JCkgiEwaf+a+bEBQZo
i7w0O48BgmrgFHsiCytQfIexFBzI25LzK0b0nmkWRAeB0KG7l1Og0KigAvlKQjST
/wzc5V8WRQUPeHyHXmB+gAmOUh8XkbR76excpxK/zFATcGxaTfKBsLOBrxf4+E3y
5mectvjtcvG6lKAhFEMBeAiMnlVpW3Nia9U1GIdqtQqNamoMk6ct1avK66ri129N
BknQxQY0hYdFZVKOfSe3IjLxqlP1dIVGlpWMnyNOrlAiH5byDYauGM7igjb70iTc
XD6Tte4lKnH/b/P3lCky8XS87kMtKThQmGf1ESOoqYb3G5XWBE4fjK7qWjqrxg/M
SDqtwxhf/t+gMNT6hIIcdnJtqtkn7e7H6/7gSAJP2tWMBaCWy3i1kY/Q2FmkR2x2
VSk8mNDRhhB9OreBf92XzUpfd48edFp1t+fc5aJFuGWWT/xb+ze9AmKIZKpfpkcI
bUuDoXQy2FmARPNxOazkCv9GxZHtbigm62CfXcKB63nS7pDTIz4aZnw0+hHfg258
TKLzyvoEk6IWosgjqiXbuUyEfuJBW2JDBmcKFwFaOrKRcK7VQ5xzNHRzcVL/lyZk
w3wCW7h6wg+HGSWgnN0tGecvWxGsiZTVtNb+xPoCCjU/zKaWc5mNibhIje7e2zgL
J5xggCu2H02bYC6idgc9HxzjVqDYfReWmgopJG0S6ZvFETBItlGAd/tmVYwbex7L
yAowoTkcaBrzic3DHI6D6vYtPa7IRlM4bahHVOGDm5YNncbY8yMgtD6JCBE1ZIRl
yYhQRd1lpvjwbTf6LiJvn5sjkzTgzJT+PHCZeEwU5lVZ3xRVXHSL90CSFa3Zi8Dy
HgcxFSDz0zWAAXOQS44RWtdHp48o+Dwa5Obp0nEOTTHZDnIx+azzDhFFzXdBLnqk
mYdVaOELciWSe+Q+zm5PlQGtEKPVlPxrVQu+73kVNAjaJ5mAnI9sBTz2n4fl/DMq
qaLEJybrJIZ6twqtnE3uPTakl+G3YtgOBhs22sNok4iRCsOx240//Qb7wQO2QOtT
AaXC60f/bAdZDJY7SaCHppeok4e+6xX/Qh4ORjODXURpIK5buG1A0FRJdNByB2iE
SaBdtUQTrzDsa6MWzmVb5idHkCbW+d77oXzwbNuswnSaSnmZ9v5vdu4NM77rX7uo
0t+ir1q3U6FlJt064DnUzKMDsufPz76Lk0OnCQrQ/RK7x/s2/Ba0bphb8gYeMFxt
1ZCHCvWL+u03U/A/HSOkAMkr0UJkbnrvmy7R4NBGPAc7+YElrILiCBMj0ghXwL1u
ONdKcMqFtSVOLnsteAlNTspjpl7McW2l78JaP4FICe+liw9XKnRzwR2pQ2SY1ZP+
2Bhng5sENyT2lNN7Fhuzq7o9x7wKXfbh5ehxTA4v7ECAkaci73SMCmC/vlQkfmbf
B9TkQeVzbgKGWYsGNrWzI5ghTHx/0VMyeXIZZBYYEKEaBvZTvu5XT073/b8CBzw/
4sMEwMiETo1sZLh7TunOQN8aPCDPvsD1dRrKPDqD5R8gxWkm8DbxsDrK9aCr5CgN
ojmGv58W6x27m+h3CaA76cqTpgmueeW7gn3LlnLNgnjRRCMPjCTCQ585slMQ+MCo
Zh2zTlRvDuPGullS+GupOHXJluGFVo/3behp3YdXqOUbCwGxzoknaNlO0h9OrL0V
MX4ptc8qn6lbWjpMo3JsoI4GTwgbBxavQ6Qtjg7MLlUJ3trQ/6KmwA1UMUPkgBwW
xg2ymWRhz0RLd4v0j0mqU+1dzpVw+a+VUqaaGR4IR7MyEIlR9/ZslTG+GqWNwMo8
jeliM1B1F2MW+/hzj4mZjB9h3AL0Mp7hTu2N46P/cLXf+VLpXNWXkALZ9j4i1VrZ
KsgH/HiAlkqzLmI3F51ry4c2kQa94UwqB8GDBvnXkvHfVKlu7jcXAdMcVZNgfEmL
TTv+1Wkxo9/bZKi9qvl1qjX7ROjGemQADahvygxzfsYXNc5ByQ1/8OSAV7UiGdzz
yOzd/71Bdj8yRLRxQBdfI6Eyxbk6KFr3mqKY6shNTpeIFULFzTw8WfRtNNAiQt80
4Qq/oAi4LJ5PyIeNZAnZzpzSCIrSFGS70guJg90WzAZ2BQUASjkEyT1AQ55CMxfy
/Rtjc+7SowowkKRIZRoOxuErsIzG4YEKZXOWORJ0TpYQQPTyuXIPEDSr8TKT3QW2
lEK7o10YNA2DuqEjHBBHCIBUT9WfJEoyprNYlaMpH9IrW4yyN+1Skg/jq1bnTjoO
S9y/gYn1ORnJl8lPetWiTDAgB4HEQy/+1LmCLGhP8l/nu2phtUVee2ga7+sq2Ke9
b6dc1mPXjJHkKohZzCEowdvNDgzNG98tbZ1CB+MFhGwG7lQu4q6kS0oNoGcf2Llp
X2R8pKeP/gt6F6Q81TJWmAWf1m17AM1iXqQaSAWogKpbl/y0CVc1dsLhJbZTH4Kj
sPpYZNEjo9d9JhH7KHDJL/DWy4OVckzEameaJ0ffFhmxrAznvzZkvounMLq/k/2n
RwOuLh/CpRqtAXlZrPtDPEzxSk69Sws/5retgJBz4p9ux4uvxtKYhrmbxvmlS+Y7
wvK2KkQoQkhJatc9dQVgU+I8V8MH10BVNhHg9dO0byDzGLXNf9PYt6m8F64Hwdf3
pXThU7jqbQQ/MAmwnsiOWZB/mjv476xO0HcUvEtH70JFmouFGoLxE+kfSlR29Grs
Ykhj0ThOBWs4Rsc6lkxB1eCUOfvGcDw1934OW4tFxmUBTkrQRGyC4Mq1l5fyZWC7
SLz1rwUoU/jZIG2FLSfWJQFdYwJCuUQfeVKgfbwntK0xXcAMeLXDw6vaFQyZwq4u
Q1Ul92I9aqUd6hmDeIM5GUReL5+S2cj1Zsb4bzYhIy2S7Lu0ZeqfE7Ixuq8whGje
iv5cT8B8bsKxsbFl+f8mVZoGrVBRB1GZrc+ikPRzWLzAU/ypL1Vo89AGc4ZyGjUE
GlW5rU+oJJetn4pltoNjRCuBJPIo1mFOmvw2XqTgo/tBwOToWi5dRQN+PxfyaiFO
Ie933C2tPKsjNO6SOZXQO+yjyIIzf+bLn0SqR8hBM+/B0xkW5f56Syg4/PY0KncN
i2dTYxKOc9HSAYJjW610s6+uwLkEkxikZaZOaripbLGtTbHHVzpolr/dOc0XVq5o
C6JkZP71t+JtIo9Z5JZ4QI5hzCxdPs+z57cYJVQR4z6cE4/gUTKkxQioInTESLpV
XRv7I+vvo9fDIr6WHxvy/oapjzDl+ck1Mu5L5SkkaZCuS5dvIA4pFq/FYn4oiL8E
EvzZjCFV00lYvBiw4s1TSy5mE8F2aYnVfMrCARX0Kd/e2lYayK0Ug6+Gzo3gdwNN
YhPgf+ain3vrSXTMKDgbL7aUEEbORNL6S6cQ/1DltNjMqovVcrHKV9OOlOD1kT8/
XAfzphiav4uPlvJeFrxH49tRqVERb2jVZKHlNRuYg63IE5GJe8fXTkjHex8EnsUR
y39iGGsyWeTREdHWKst2CI9ok3j8Yy03Ap7VZ2Kf2q0=
`protect END_PROTECTED
