// fp_mult_fun.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module fp_mult_fun (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire [31:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [31:0] q       //      q.q
	);

	fp_mult_fun_altera_fp_functions_161_kajft6a fp_functions_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.a      (a),      //      a.a
		.b      (b),      //      b.b
		.q      (q)       //      q.q
	);

endmodule
