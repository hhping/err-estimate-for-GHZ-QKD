`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6cBK6RWbjnpqRrZVOjHCKG5Hov8RFnCNz0oydXg0yK+57vQ4L1MZRKQWP0CpynA
wmhI9CMsAF3aeizA9wXNmI9pBPvQne54Q1nJph5Uj7FW5A0oNzyjJBXP+luspNGf
HAwNV3qdhRKmaL5Ig2vjnZKYa9z2e5saWvZbQ/NPFW61TvcOUOMjLS0P8Vyi/6sq
+t4+maVp7Gw+ZxCUqdvpGOc1R+0PaVV04VemU+fFsp959modMzXqdh0PHN9uUClN
DPqGpdwGkdVQxzp1Epr8XBPS6byYqlw/9Czks8P8TTM5LrBtyy8oGEIN4yMFpg8m
hibBiQTZQVyTZdqr//31VJyDJbkBn+rbV6JbWCnjBOJ5GLKkW3gpdhoZ1kJV2b68
6nDH1tUJd7s6YGZsEAzbme0l+0TIC9YmkeQuokqivSeZGPY/DWeijexGrHW8e7YW
NYp5Jlgw44Oir0MilJp3BbfINw3S97V1aIVcf7WrbI5gz/ELbt59b96+gyw1nZAb
ALolOdtADrKiGwwNwYRwrWl/zOjRzwrPELqBw/jwF5yfhWHJQw09NhqtsHcGvrSG
ZchNHoerGxE5mWv8CqsIPFt7iMk3FEzzxE20nrKkVAwnjKJTfvAd+ulXAY6vMDgu
aDbxK+OmQUnDPirfB1QY1FdfAmhEwbYbdNzSFGcWCWkKxHsA/74kw1TMWsIwpScX
szOuaBNuWAu2xYOIb2WoKnh5b1tPuTIFy5q9Fz6oRV0Qy3zq5A4KX54Cvy4rqAIN
Uj1YGyT+z+VvTCzLQOBOs7rAMTJ7ofG9n9ycOXevlMJESn3ADokzdeyozstkozf4
whqeJwNg6Ok0lNHuL1zYzndeIOW7qNdx07wn76X5LgSppa5JUrwK4y90k4lJwNFd
r5EvuZrMczqnleo/oZfWKE5sRXt2DetEFVs26wF+xZzGpGZrwW+XFai/h7ORJ3F3
7Nr9V+e1QO5zzZKKLw2ztfMB2chAIk8Eqc8cIskM//GDJGThWMK2AuIsICF55Avk
KlBuX5Z/z8eXPsqkJHDS0aUBhdnl5tlJEUEPfy6g+VuXuKjA5foq0/sOJw/zuHkt
WKZHPfVDZVDv1N6t0uVBZueOzM40fzRokGex2DToaPzWIj1i4Lhrtcye7pyupnOz
DxVuaGgl9zifuO51Ax0ZlCVTHr3g8EBNn4XclHgNwgbd9fkh88Byo5ZvS3t+tO5V
2Yu+dsapgH/V/c7sJnhdSM1nHNp66pkN9G9oBBD4WRQWLBjlMvgl2uT8jKsV0rji
BpPTD8iajvayrkULgLnu//BKTAPV2zsj0EnYm4r6hyCLBFlyX1xQN7D/Mi6UglUB
cR3GmEtqV7JixyTjrinfxzYAMpc5thHFZOBOLXEcSI/N+UqpTFMIZyd5it5MviKe
gS2s1p6a5aaMTWGz29tEbN9ynlfL7DkVMz++StQY+3F7i9dc0OlrpPy2MJytj9Ic
0LYer22dkfBzgTiht8GAMy7KfgbKzJ6vU4c9TF8csRvwZF4leGKi8taaMkOHr/2B
P+NUueh3I068+DqOpRRXDMy+o8txu1A9RkWRMEP9yascnLoR0+zwbothc2mxLKMn
NhVMQDMm48i3W54Ty9IGTE0/hq1UKqxCH4VAm3QY0rg58T8EusoLPSMKcWvBDhIp
4vs9EefRuz5H3azQ/KaI7XGeSjL1jdwR7mpA258IZC2de26L416XFFHBuzxCv2AR
bRtE7d6ARXn3piDBAXLcFU3Q0aW23P6Ali6fNl/QJTqrH1X+khU6kcJXsOO9ksot
xJuGsDJfsb+NclUYX8bzoSGg5NLpoWOOg440qwjh5esBDT+XNK+6AZkUgqtcqhiL
52DlxHwGqolsnOssxSVZu6t0Ly2rkm1qnQaYSOoknVF1Vxg9cQIWHwfztoQKlNg9
14lMGOTDchRK5FEeMWTV8j9hV20D+UMkwwrdUL329rtNlVfoC6AUprp97EhVuSNM
LEyLmWmIo23+DFRHKvzp2+OV0gitKO7Wffvc5LF68vgtQZ0/+MCAdGFssFTVH4Wl
sD9JXRodv5MabTtehcfZvMKEuFXowBYrcZ9zENAig1YWPgPifF3bAauKBxgzYVGl
2wUDRDX93iYgS/PKWWsi9g7dhS2xyUvEd4huVkDdFQNLSghXsz2swPZlzqe0vJsT
9Ttc665cXGAM15RLcsNL43WqD00nzz5jxRKuNwTmvSTOu85lRnyHCJsBvFk4kFsg
GHFWSwq2/oaEXODly/z2UhByoZ0D/h96afjnlBZyZr32mLnIrkC9pIt/jMcVWQAv
MHdOBGVpJoiq68T0s6qUL2WTjgZqgkzIp3qAObgZIj+7WNKhEGNlEEZ/sBngA0fh
fZBbd8fBSeE6koKjJ7poZxYrmNgBDSmcbJTCGoDDKPGecVxsRQH2kuxhs/WB4TYn
GZajN4Q8MrkzJGNJYWMfrRiFVioKGS1xRmKQvEPKRWUYgpYMm7pydx2HhfgKpJ8C
J5McngacaXpjrf1Dz0O6Xc16sCO3drQIjWy/+X/tyT62Rol4wy66o7czod3+uVV3
Q9ENlWZoh6/zVp4YpPWQvmF0cCmies11WQyQ58f/Uw5WRG9zuW8H3ZA2G9cof5Wz
YinqZYx60QQdwAM5BrXjZME8m8+WU3i1u/CkTGjJ/u1+MEkqHp121hk9jGBAIeia
SG+bYKvc/AgQc+qe2by80uUO8l91/MTrTlaOHlb3xSPMb+JfDzNw+ESxjnrzTKzH
Y2CRC8Lzk+KBg7OyElHLBkSk2DYnxgsnO6aRhifxsYJjcFCpqmaqxJiVy9o/mekT
6DmO4NDOnjoXZE5xGXcVppAg9H6JG6yL697q8TQ0s7p36mXn4nWRmfYOM36L779j
xeE4FgAkg7CEwjZdBOkqVTXAzwrOVmX5VfQFrRAn7l6g7KEjL1aN7/b+Ji8iP2E6
D3Ag/lckA4IHp7bJzKf4ci75k09uwy9DVpo/7SGKotAxynn3AJOfvZReDaQhjWdU
5qkBcxS0Xd+Kj/lub7SdQ31egB4QLZ3S/fzmH+CvmrMnlFxa15Bcr66wbH/ryhQO
xo0FQOGosO8mFpMJMPyKQrnOc01RSsHW5DMnyZT1y1QCARt37dSjsWP3QXgSC1Ni
mCSuS1xNYCIbM4sfQri5k+IsY3mqq8EfnAXKayGJ9sjNdY7M3JtubUbDM7of7OVw
FxfYJJUvSh8aRg/Z8p9U92xSPEdokeJLtR0LlErK3diLi/UFUO5ogf333yNWtZET
i59C3kta19Eh+lQx0lcv5397pUwUoFGswMIMpOjkT+hqAnA157MDcFXwHddWS2WO
`protect END_PROTECTED
