`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5GXrF7I1HEqM4H15H+IizL2j3DuN+jPMaRcUlvXI4gN7bm7KL4gctR4qPkoaYCm
nf/CFq/+On9hNkbSwwlRWOlJ09Bena5Fk3Hy1a0bIwCxqam9IPEgpdRAUXrcAPT6
jiUSP4gdMPNF7yAlwRnVUjYwZAvUJ21Bz0a2kpW5FAEGS9D+1zt66RXWBnsblB2u
1aOGu+aV3QXfBNDNnrFWwZfvDOmVLpPIs9gjdhtdUlR0YyqYn15YZQrzK0L5Vx7G
0NwoVLubZups1tPf5sAUficfWwF/zTrIuu/VyqNE6oGWo1+jnXd4cOMOByTDpd5G
YVHZUIpwKzvaDWHbtKtoAEXubEev3EHt3x9VUWowwnD5nzZb5fBBlw5NZ9xj6PJV
dUb7lcNstrPDa0aocxOH8ia/3KWCSvxuV/nwa7nafDLPdVrlPZlDDpJifRV2a6jn
npqbcyk5vhKcqq3MU43/9XjcS4X9IcRDBqjb4DtMA07z2Kwymaoq5+PuMR7ttIap
6ojCA2Txf9FfifsSvwqVVFQ4KA8yqow+rlN2xe+To8/HstLE1MmnRHYQ+wK8Svr/
wRXvelygt/Dd+E1p1pBQOMge8I0EMqaEY2GpYy+GyyGygX422Fxqswbb/L6ObmC+
amU9GqS5C8ZeIHj0Q46xNk14KHeT/velBMopb76OcqUABYK94SSI/EA3Pic98UOs
eO+M2IogX2ybmdoBExGE01PekJWnKbMGAgr5+S3e8MJxa81Mv+x4DY8S9ZWBLd5d
8eZgYK/+ZOlB4+HWrHUxCiG9o41RB23YKibmAgusaMpVf5SFR7VLZtmcFjOz/ukl
9bvMNruSLjoCwtuwtworj9XmohImzJZzSceNrXgqver1qt6Egv3hd4rPSCyGG/0a
Lb/pmYWXF+kgiNUN8Ap7+aE3yyhWz0/y4iEpSZVImzW2ZTibimOA7Bf6ds0dUVEs
B3noHkBXoFZu9YwHuhN94ypGbd5M4HezAFhQ06IzmbgBzO8XKa3eApYCmMjSAbRn
19j4Ls7zcPv/ZCWK1EBmKzw3Qx0BJeXyEORdo1dgdqssZfRlSB7xZyWiDdXaoktq
UoHhG272BXnVCoKVPQNsjtMA0ZVXh0qzLjFyeaa1RcGCjsHaM8SSKuRjLenN7Krb
VaJSqFFyEspcYYtiw5wABxrVDv5J2H9D08FNl9rQ38/cJ1RcHnB8C9Jolfk7wLrc
7KKion6Q0nyyGI4KDhxCZ3nf8WA6fd0Zodo1FN8pS/y6ybM/wIph44cEqf8jV8gT
hRNOhFtjrElGrjaEGS3n2KlgiclvqjihZqxIa/AnYWxoanpVtD4UEh8dD48XtQe+
Z4zG8FFfOrPVbTeZlpUTd90W2hxlidXwz3TTJ0EUI5rB3CXQJXxn2ZqRN7Nj89+u
SREXSBj1GWPHuXMzD9oB6XcTFWtA5hcDEcoNf0cujG7k9WPjYYXD/R/8EeQLb9v/
a8jTps8x+Z7ONPomlhMruSEc+S/Gh+hCrGYiTuwHklix3Osquvg4W3C4r2OCJirs
VKLo08s9k8LArg0lcia1+i0c+/qh/5GnAf+Pg9kU/ATEaZRKgXINWD/kTdvYbLSn
NjueU+KPttqX0qxGRTtZnlxdWRaOaGtVL0fyfqLO84OcMduMiT7YB1H/8zDvcebM
vKraXXEMgh6IZQ+O0NKTzKUzRmxw07/9xkAXQ7LeTkd7YbD/CFuBJZSTjnllA14q
ySXr3zZRq3Hq5By5ypUUGInUZIAw9KVUAOezHtw4+TUH4K4mEeFmAkhGVH2MLPMd
6r9djeBmNLd7CvGxSogrPHn7hDbDkYY0pFd5p2FJQ6+3VV29O8luLi10XtqHkPQW
r9lGAusKhIUmTzsfJUln4dTvjNyJBH4vPtr8HAnMs3Yj/pCBriZqNpiiIKNPIReJ
6Q0ZjpV6WE11M73374L9Lb062Kp9cP/+6Sn/Ox7wSJueD4TyhG/1Bc1/XaylRk07
uliDQ75KHXpTFZDX++/A9RCmB7dWDZ5YnhRdsfyRqUt5JRUahSvs+dGKhT/5SFwH
5jMRx9A+AE/GW5hG6m6NF8tjbnqdRCUVfuVt9nJCgJXGr0l3GWaBt1WAfmpcCkP0
cAJrPQfuKiSr/zD1hxRvGoJM/Kx3EeVIt+udPNvvVUs6B9Ts+7kx7rhSGjHGzJSp
qzUWG+p9DHloLNEPqyKnAZ9sRgFHZwyMd8PztahwJvd3VbbXGkvnOgs9KrKzq3RB
BF+J1PsaMKtHe6OmC+84Y1kgf3z+JUcSnXEnTWZtyO+cdDwJpwUpIJNmYJbffrXR
QhSNkvv+gjzBZLtXCEr67gzxlbam3QaKv1L7Mq4rvx2EIba6asKPX9G/GoxwtJ1o
WSilbEICFCbxBNSskvyte7ay33xi72TVefSphJVf5pOuYy18atiwD5RFOZ2IIOSM
PIc62A9oAfMwPtbY34SpM96rXyXam5VBX4b0y36fa6SQlwY23U1DqjqOhcrDjpNk
f02aP9uM6BxzzpY/eDpn4g==
`protect END_PROTECTED
