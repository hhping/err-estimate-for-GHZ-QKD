`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uoA8fjqtcLioajLn0ikGh1/9mcZv4Kl+7Zz7yT7FrTUhUSPuB3iVG4ii7yHKGkPh
JwPykrIl7imokFPW0WZWBSk/L7Z6FcNZgnZCB/8mquMzzEAs3kMlPDXr5gLdvOpT
Qc5qbZJT27ZTcFPz/9n3+C4Q+dLc4gHyVdiA0Cqf4MbQ0K09K+nSIntAPcHHvfsD
EA+ii1M4KiIZPvp3f+6Cx7uqA0iRmbpntIN3u1tWlM//n8owr1VuSlcM8snMH9IV
qpMUTwCh47An3qaDRlFc7RMywbX5nVsT9BHlgFMcjdNY4uI52CHXnXPr9b0mAggP
80s62DbxzNHANpY6MaF5nylVl+uItoDAMpE/y5CBVLnfAmZuXWSWXmxEvzpy1nRJ
9lk6Z4uCR5+Bin/s9vBPaEdk/7vH/TS2EvQJFzaTC0JFsW5xoXV1bOymePCVXTM0
8a0i+OhTjBWhdkJ2bh2a9m7gEQeO6EoVKpI3xjsfunSjDXj8TYuYr20AJXFIrPMF
F77O5mvr3mjr8teHl+A7kU6L8krTdpCUFJswrc9qcB/7xMyuTT040sBbef4y7s5U
rYUcHmvBxj5+3B6JKv6DIPfePnJQ13BA1+1b6hXi+HU/mEtkt2YcSqiOCuGCPy/N
GjwXzL4XgQLl37ZG9zn2pnQf0BMMdiQXmwWqBtV1C3RVNrDNyDunETHKF4W7kDW0
28lI2DjTpE1cNoqt29LMzBkh8EFXB9H0M+MgcgRPK2i4b92OAH9r04o3nrlqBMDC
+m4elKdkurJQGEtdZe/XxgJ0ymr88E2jNERQSwxk+zY8XkFXFi07qZ9+0CXMAAcc
D4uEEMnsq1jAsaAWK8G2DG4+2Z+Z3XQKJeQp013QnRJuuHSXSuVKe1I9yvqrzLKw
vAFEUKftRyx6J3Iidqbv1/L7gXRsy8KscauezwExNlOJEeEV2DhTUf0RnwZESL/h
GriUrWh+3NFBiW/Ebw/nzIXZzxRXq2gJT2yh5yXZ3ZTuKtYp1Aa9PDb6YqHuU7dS
vpLXahksG651G6i2GBzLX6IaLR1mQi0L32qo03Lf4zYlkg3EC0L6Dj+qswklmpdq
CvGRnqRgW0EVSR2XAq6gy7mdHDIQs29tUplcoPIqwCS+Q9+JP20FFsYWRytuuh90
EvdhY78PdOhhhvbUkPFVlQw0tcfQp6XWwWL5jhJrq0OclKnAmLNlgqEPcac7mlAv
9cYtsstW+TpSxKVaZs9pIh3YjV7kZCvMbC+SKnh7iRaVdWlSa9rhp/Ysl59no2Df
BNsVMRk1WaE+GpoBJ2Nyh9W8OE45O+kR50GRhv6Ln4yxeKBTH1vzAjaMMB4UM/9s
383eH9J6gtbc3cZbZThju+vWzAvw1FbXXSrIRE8NbSZ9qLHabIUFQ8JnxDeZj5ci
QU8zl6m06/hHOlflIuehSBNF0USU8YhRaEUqNWqrDrifmL9O2c0eJLnzFy++sdHO
385Z5SXjLM4WlBkxV71QfqMLbJz5EbWfr9pes9AsIN5ZtdFIKypO8P1OZoqUfGpk
7CDHaS2obiCQ1WBWtldBUJ4qH+zbaiKVK85ZIWy1vZ3Vp/1JuQTfLB4BQ2N6fWv0
jalcy1XWomgQpH3OUxakNoyj4XoFCHbnAyJf3WHFhsozQx8hHupfHLT+TsZmrA/s
jpWIU/piGP3TUAwPut3BXmyRUo6xKShTNOm7TuMmhF+G7aWeHxqdaRD30hvA6vl3
5XXxZwyoxvXHNWsflyAQFDJykiA0kVTH0meH1VHHFcIZdkgJMEZIMB0Ul//p9xbK
fA1sH2W+lKZWq+GPqgihXjUEdWgGOVjl23ibEaPf0i7ZAHDn7ZNtXRV8HZr5YICB
bU6DQLErhhO366XlKIK4jPQdj8o4/DISsPg+JJBP3O2RvhX2zO+YC4OzbY9FFx7D
UwAzAB4NZcVxprg9QdZ3VCP7Gy6IHV8boHGIAZ5G0i5k2MNtUdkRAejYli2AwcYV
DaKfAaduC1Ju5Krpr+lB9tztJf53nbLci7ZsJ+YbpXCjnvEM4pv0P1PFhtBvfAhu
oNPbSJTkUJ5Wfe15CvsNwfBFtNWSr3guVKfJauuOkV68bXfR60Ca9ie9mwSJmSb0
Y4bouIwwpubL98FGZOwOv3NxxKteg1g1MS2gOJkM+dypRdEzJeIxczRJDAjJ3tBJ
n2HhOZ0Evi3eIqFDv1J8JxNO7lfh8iUVzXyggwqnRCBH9kqCDOuUA9/cxS57m2pf
9jco8UC9xKszFV1r/AmqQYj835HY5hGjVNIGJkYLRXmq/qvNSr1Rmtzw2PbOS8Zq
SnmaRUhD80EWuynidvtBX8UqwNTyTFVhrIvlARANptvnjjlfGSpwFPr3O5I+Plry
Hzl2LzZq4u86MYre1+P4iOObXIL6IzVRbmRg4APo4xQBDaao8knHNyOVmpAK06gn
uLHTkws+6PZuk5unDVZaFJ7YK7x4+0/w/JTpXBzXGtrwfHV9JD5v907f1TVouJcZ
GYpZi61K9Iw3nrMQnstG0anyODfBv7obQAl/Jn0+uIK/Ua8FoizjviQe/X9j7LKG
m/1yfopEgJkElUPtplr4U/TLh7dh/dPr6C2gST9ODbqG+gNuIQaJMuCH1Xr7RL2W
14kQyhvROYFHStK0kbUDyBhfuVazX/vmWry9t/2KcxTphHdaOdqvf6VPGqHr9tyN
k9dhUSfF2jTtE17Rvj6NKL92vOyCWZdQ0z1fkPtRhe5Cnf+miJawITsgwqnc/NZW
0Q3e8W7vqXA+NHQi1+K2YXo2Tw2nOipLdDJxl194mNafWdIFFqzLVfrxs4nNWKs/
rzU1WNytH+G9M4CwsclaIgmScN1Uche0+S8jBZe+ffSuPSweDgbgCgxZc7g72keQ
fBQxpYrIPU3dRSFNNouqQ7MH3L9JnoVFGzFYFHcFSqU52rfnU69B/pv0WsupsEI9
EoqGUmzX9ksXt4AAX5/lux+Y09jlinDL5cCZatgty2nqWhIlQubIMEzolttDY/ck
xAj242xJKfX3lW8sUgkTGWCxVUBvpR2jYBlU+/zek8qeRA/l3mfWsZf/AIWq1HNS
UOr/WHzWIbwfU68KLsCtowN+hmJXaA7w7OEEbSx0zl9sTTAVBizjZrObp5SVGSrv
DUbTkFrhpSIVb0s4kVr01RJC9y3KF/k1+ep7kgL7U+IumycdBPOJgANfVt0rNbnz
CWxp/lPYeP4LgmCVaB+7lA==
`protect END_PROTECTED
