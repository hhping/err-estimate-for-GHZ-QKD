`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4dYkZJSKWvrvJbyMoZwfyWrT9LVU1sYtCO8m63aPtVty10OYfRXN01TZCAzcn/b
YIqZMyGymSB1i16UxEbHaNkG7yadsdlmvhz60xcCkSm83AfHnZle/UAoSOuf4PR0
KaBFJa2smnQUsQluiWHSH8aWb1o6ezy4uMdTYZlOHvxIyr857GJ92pmw/wLnPxd+
+FOaWCiEILHP9aue4KsZcAdwtV0iHg/uUtU9L8WiEPnIdyZkCJ4uNgjOf05u7DO2
D3wCXd1zcNcwvceo0y64FCjNl/wBGO0/FqDyA3fe52ghlgcpXWrSig2XIo9wxaly
Ta8+CQO+ZmiCeKEV14S3hcoNmXSEXmaUkIunRn5qudaxfNzUO55toqRBmrXqKwai
G04SxEUsW7yUQ3ByDrBHBK9U7SM49f5WiCGsJspP4uehE2CMS4Wh8IHcptmFlus5
rmw0XnPmsvO24rO/MtPjgWEtLBNgCPv21A+vLScIdMc+aP9krAnSpe0Rdp/VR+ZA
MLgfTgysyjhdeeQwsZZkZlFaG73UfA+ULZizprtyuSnDTlp/k9wvXBZ8SLWBlk8s
ecjb0RTwHhBXQBr06H2s4VCStxqCzJaNdTT1RldJZujWwDR82+x0UoAdWjovYZgS
g5zlGuQsTv9J79k5ptMnmgbfgMqQ0ZFicDbc+C/jyPhwAhfzRAQe3iBxuGcLWkET
YCzJHmYai3l4Ifvn4uL8NqBhwD/vjM8VCAGqNPCMUlDa80shg4CqY+/jpS909tqg
3I56VY4Wbw4dKCWIXIu6OqUc55l7Bn6EnLxUHc3lgx/tQB6QWGFaplCIWxzC+Zqs
/1RJd+a7GcTzjBgwsfvV/wymFt3zUz7jAu2/oVwOaiH9jIYgQ0IOZgGBynnb0XEG
flscN1GoXmZvUO6MW20PFrBO7ZmKTpIsygEp+clISposR5AkHv9jQH1v6JAsB/EN
IwUaobfP0sQ01xH5QlypdbwTB+on4rGVAxa0foj/5N06A//7p/Y4fleLtXEZi5gO
s7TFJdmLr4c7ul30d3wQRj9cLapU8Wai1oac1ZqC7KIN2klm1CX5CZ9a/pMcVhio
MBTEBzx3BeMqqhK33aA/s8geuWCR9I0zWEVUkYk5QWSNVjh2L3osLEFgdCtMhehL
3Ho+mcenzjPTxkfANeGfSJxmQv+c5TcneNL+4sYs4N/Fqi8+Ouqtlx1p3FMJjrmP
g8ILqIyn/mr7lfSY3k4qXgwxDHZq6LDhKgMRKGGNmZuyp9r5hVFJlOXbih4/xyc9
RCV5sGV6ua9OBQbl5cZBWT53jfRx+yQ5IfWZkh22yzHUMqhLesm+JogYvfo+oL57
uAFfdoVVv7zMhiz1esf19IFGM7RdJWWC9ftW8scgBzoMPJBopA7/iNv0tf+zzqmd
r4BgOHca9YyxfC005rDNW/3lsJa6B8epnJE6+y0BiIEnGsmM33JvG+42kzbiBl63
0Lu/G+qYZOFVAzE4Qs8UlhAewcqb9nco4O8y7o4CC3R9ZAk5EFvG9l4OOVrC1wGB
R+F6nNIl1+lLBUMNhOPMyafUqpnfNxixjYXCLAZIjQ7MYRlHJEo6xpjk5mY/Rirs
AhMKYN3OQqtJXFRH9WDyAgbpSsKDey8bB0l3vXET77sbxoE2i6vFUEQUFxJjp/aQ
RJmwP1IYpSzWKQjTzHusHMe1BEOaIFCTxXRH6x+D3G+eibHM7p7F5+6tSBEW4RdF
rHAraIDMPYJZnhkzyz0q6IwaqZU2+WAcL09iNiKA4WKA6Fz6f2Z89C59eURTZerk
SO7UVMH+p10rJVtJfibUsylr1lLC31c3pQHFguF3zHZCYoG02dY9nrtUMH4gVvpe
tyQkFl0pSNzp0r/XaZP21ezHOqT9o6CRu++sMm9dQlMEFRduOtsruLwL6DgwNA1v
XQvXPpQz8e8xNI0SQB61T+jcEd9H+d8Ny0M8wsaZwhA=
`protect END_PROTECTED
