`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0e1VOFCTI10U4w1WLP87xEqStND8/bz8jYo6kzS/VphHOqiRhgd97klyvX9tukeu
URjmHExuh3N8s+rYzsBpdhU/4k+B8WMFSVRONJvAI20Wch4aG79B+BwaJCxBDbZy
FrvKbPpRrkFTJxYHb1hBZjMa0eBZDlwqoh2sJw8WtXAplltL8hC3jWZ4mvUjPX7e
5frrw9XgMdLCQQx4taZjjbj+hihgHBs/AW0VFe5CBoX2rzR6hW7xfQS7sr7802sW
RpYsKQxnk8xES00SPjCxILgow5g3CubdpIhS5wE9plkzexgxVF26H8oi/MhOKPxA
zfEvbZiI0aGBjs61m7u/coHCUpng2mwhuuvnqrR0AZIOMGvb1ObJUlrktLEzlzkN
ia7qLkK3trtquIinlxW2uNzWS7il+pynQGNZAEzt/6cSyBPgBq76h9awgmJM1muD
V4/b1fb0babMATTr471R0T/24CdrVkA1N4XdD9sR+Cj0IhQeID3JZPEaaZLpVW5a
vyth1V3bKxEuhsjvBcm7UJoZ0LTMH8R5TYMufgNRyXbEHnuErOeHWzHuQAq39KU8
JlS+B7Ozln9I9dEwcEr9zE28WZz64NbuF3/LuHp2UuRGgeUNUEwkrtw4p5EuyRbJ
ZJ3kiN7gyrw0mIuhVHwYo2EzVGaFzF/+ojDGhyscz3bsVdFuMPnxFjOfVTc58LtD
TGgo6+TktoZEqM2jZ8FffOE19j8/p2HhusLlNKqKQ8Y1dyONsTgVg/fuz7uj21+f
2JZ8t2/Zxl7cX4Zju3z9rmnbdYD7ssv1mt+P4XHweAd6CuwgV5WYFpSysKbmblBS
bqMAXZX3a/df/8M0G07JDT54WBNyRzEhI1j6IF8DNKKX9idMYpaTPjlc5U9Yv5Dx
NTNz7pQ+8uGAKYs18fl/ZD/vZ6HUm/+nvyUOLb1KIOL4Lu57wVud2vZ8uxUPS9Zw
/bU8XjtAf3TMTtmc/34vdQ==
`protect END_PROTECTED
