`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WkSCCvNozfQ5GfyThNCJtbKR3zgNwIO6SwnYncVbe1iZE6V1+ZadXinvDWSR/PQ+
T3QKs6XIwqOCVuyGVWjxpB6Ivya4UgjOygqpthJ8WjeJJy5/M8XO5XkCBNeaMFmN
p5gN//f2753wYFkri2apASF5Fn5SrWIxzhvImlEKwvBT+YwtgDuNpZt/qerHyJRP
h5XYUTongZxLWiyxs7RvoYx5T/Ug+TYb30ZQ48sl+gD2a/mr2C3USL5ZVTvs7tBZ
oB1xn94QyAQ7B94q/epuK21Wb+cvDrAdMCJuRr2+0zQJ9U7zADTLeBSByv0Bv0Ss
7ON3P0AQpxbhUScGv+qniW0pYjexkMwwfC3M9XmODR4ofym3Xc/wloI3KILw4Qnf
g7a830QCwERV2R6Yd9CwmLAyFpYXMshRHrKysQAhS+fbwoEynAXyTZpDRJyHhdV0
RZRcAk4lhJhlf2heo79uN+eyQkwqtyGus6FKaSvbLH6W2iyvqFYrOcxWPYQ5UOQo
bumASa3WVz71d83wbkC+F0iLeEnAAJ7DiXwb2Qa0/xmpnUIbxbutnAiuSsXmcEGZ
J74qXQ0Y2zlID3n2fWPC0QHpTXyxxQzUHdtv0oJgesHQM7GzSYn4a5/izHhczDkD
iSfUkNR7hdKbKJSCSrhi/674xSeHZIG0j+CKVZIpyb/wGZDLbasSBeYVwqZ618T3
pMuXLIGgVNz03iprwWOijGrXC+KYJxyqHsJXRLfP+6RDKoCekpFzlIBagyIzA7+3
SB79jDdAm4eJQshfnKwlcd1e4ArmO3ktICbmk9Jozz7D3oGxnPUpB4Gqju20hWr/
De8T0vWr9TN7uhXX+hfOtSMSENnZzgF/m2n45JbC5H8tkVVjCkcuUYbCvlGWeXNe
K9Yz0RUUi9UqxSYWam0U+UFY4tLT0KqnUVJ87CwIEnb7uslcI5bvS3QWdbKJZf4o
8i5D6RTlNVppXdRFcs2RCvRNeKae8YC86ptGy7qEjYUceoR/EQBXcO0Q2HXM4gE0
6wnKcXhxoJIkMAmPBCpmQle4ntcOy1PJ2y0bv6AehvLpg/On3lnbGLKPzQMkAWcS
5zSxohGQIKDbk0+AR87NntP3vBvdt/TQI7cFspeiD5O4u3MwqSKTttLrlwJqsEpE
My/t9d7+5m4Rpc3uTjLDI9QBOoc7Y+bLuKmeLTyEYz6OodMGgmF73tBehONLcFnC
dbNssKXwQchnastjOE25e5PM6i4bLIntKcP5jrcZaxoZUMTmVRbr4P+Ab8nlKH94
CACsW8NNfkLzeNilE+qqricaCG+9JNsQ8/nZAP0XxnQwNnzlmifJ58Sk4A/luAFy
VRO2qn0uYMJqm5ZvCM0vg+ynkSRnnU/KucRNfKXBgr5P0aV1f54FnButXoHko06m
5Yik/JxXqBVDD0WA3taGDW+v6kJkkLXZSdq6qP0hljGcFkhZosDc+d7RRRv6/cSc
6JzXEiikwq05LGIJkJBU80wvwtMxYsDNOM/ririq3EhIXqdwc3voqei0ggPlanHe
INbxAe/7yOFMPIKt4POPVymJPUbnBGDKvft5pQTqT2toxWUhV2e2/GDQGYYTy9eo
5O0VVZwRhhYL3+FEE9ByE6zdfkTl5+SVodTWK/2wf6N0Fa38poqAuNzXatpdAOc0
4xinSLfrZ3UOU5Mg6M7Yiy45ep5fIP9jNaThDVQW2D035m5nBGGNBsJpWC746loE
u0RLxKmPOgC3rSv0U20+amEHM+PHnD59gvz89QIvvkXZilsnO7EaOogLbLkdtleP
CsSKts7+2HR9tAP7esT0JcUBGOzJgXBiqE6EZnkIk+gCYbhMTaxmAl//KUMIczKz
JKDimGv0OM4ROxyeVg4zJ5xwsykKSw6Jb4aqJtwCtZSKZUrIx6107qU1nIDPnhAy
elPvleF9wFU6H+so0A80tK9rSkGurVNO5606VLJcALoFi+1jp88cMqZVnemRpm4G
OCv9wl8Ckw+3IQQduwI/8qWa7ZwyChj1h+gZ/ICWHHY=
`protect END_PROTECTED
