`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJ0YClvlg6ma3vFKFjJGqY+6Gle2sdhLced/6GHtL48bb8noj6gbxo9zl8BegnAP
StbEoQVGqCeKjUKZ455AbhNM5hA4+fJwRrjUkLQCFUjyDotx0swuZ+qWqlUT5EJh
cx+CBwZMICtpehmjfZzI/pnaUAbRF7IMUILfMN4+Cg2o1lSnaZTlfs60F04JsAO4
zb6L/oK2xA3dsoBqORVikEyy5GlUKSUdZ9Zpp6K1eFDfKgfDT/7dcTNlCmmJZxSV
1lorHCIZ3mc+ANMZcWwDrDHMOqwHyLXSSa9cz6akJg8ZSD+N0AnN6/sb4Ry5TRt8
j/91vQByK7leUSwkJQEvDo59LSDIcvo5vGSP19RKxmVwEnyLVng4sEA54G0FsJqW
31nJTT84lCtFjKu2w0yuoS3YVXLccjFooycxyQYpcXpOZXez8hadjVAl+YxCjDxR
L4V0/Jj5U4y+vdb5CbUjPNqfcLe4dRmusl2f8D1lFpRp+W8JkKlHBUMnG1F65fdi
j5tYmfz4lxnfbt+jhA7ToRCkSxtnsOQEt3KBlDhb6ig5/3zHLoNOYmQzAWCbX2HV
8zU8Z/5HRhf4WEjq6m+7GUbBB5bz5V9GxE+M9R4tlcCZEuTNuZLtAp6AvpMdkNWh
oRAZ1XhbTj+VcHwp68Ppq72MyY/IqpdMpLSvraZaRdo87XoTasBw6hpLE1jaeuGF
GVuSTaxlztX59nFcsatyvG29/eOd5+OZS3x/dd9BqdLtX5VKj/05VoyuQfHhHUCw
krxUtAJdI0fVYCqIccAA2ff6YE/zNyhGQTE/MWCjPRcwko/QPrENIX/9Ags0j74w
+PdBFgj9VYMoELEIZK04leo6zmluQh1wA0lg3bjLK7zHLvw1KZoJKdQmZk9BEmz+
jwNZIs9HBXcQaHU0N7vd7S5KnfftrBj7RX3Er6muNe8FzLzAykJBueFQTolESKzD
OIkUJaasS9wmimdxgxPnG15q/hMu9GQFw318gUupVPTSlaJY9Vyzh0xMfIEpHwTJ
4iMQ1XzbRtNJRsVz9qFL280lmBeowOeKYelPI8hukWBEUhIkPzBfnMha3HR+WjqX
q/2KcdAFqR2A52PwqszFJcFQlvRzO0bjNj8mqYEjEB76dGiE2/Q4vgrV6LOVpFDm
TEkGcNeHrysAxaoz3Om1gFpAjlgIOoaEIUjm1CfIyDhmxji95e7+zU6D0JUwYj0D
pFIrwkDMGj9xpY49hcr0OQyi1gxqF8VRik2WIhjI6yR7QDIcYRkRi75ZI8P/Zv+Y
Ih0tu2GzxvbIEYOMHajKScG13cNsyYBM1uZ9w5pJ2eDxcGpKk63COY4/YA4EM7Co
vHZU7UZoDKNndJIxOE9k0o6D2+IwDPLfRnT/yyKrpfPYuSsBg54x/vk/kn03srwn
eOBiWG2e7Y647nZAvaOTmwg37VVNQLJUfLT2kNGHC0j2oWu0nh7J2+xXwhAlotxi
zdwLddYaa6SvFx2vqrz+9YFnevJqolbMPbkxLNYsAZB42uYYU1Cxti4zxaCveN7H
irl4uWV00EB63RXTF/JHKOOob6bvgEKqjuiGhSwJD749fEuKJmciYkuGCQ+go2/N
Y5VNFV1z9a/KN1sYgLu1zUR7eZJJzn0x2c8ukRZNg/lCgSqYf+UZJEEn8cvmDHTB
so27N4DP9kHrzYoZ7V2yWThgOGdZp+HsAew6ot1NNtePPnqrxB46JCnVaZe3Bn/K
oRFBLTKY8BN0iYGfKyS8FQMCR7nwanMLUw06ru0nSJ4SCFgcT3LuqJXZafi+viai
AzYoAaiLJfZhzOlCN2JWpV9V3NfTnqEV006pZ4foUH1pf5ENb8lco8amLpcew5dO
m0VOtKMEo7/74XbIzaBiH4sF0G4RgeBdYr2nmpxiJhi2XS3oFerKMOo8q1p/8Zku
8lAZwMKKV0ikuJeCM41hKXMfnsqi2SOQ1NEO/hrBF9FDNPX8Lo2xCCtYTgpf9+wS
9D5IFJN+l/sgeYid3+OW6fzEyRQfWTG7R2Ju33MoWNP6+QiCduDaJSdGhP/O+3CC
3CXet9X0gKImb8X6Nace7+RyjQlhOVq2aQVR2G6anJCB7iX4IygeJ0FScFNQjNJT
TbQCqrDvwRBEB+m3li/e2dSdkKSzjukw6rCM5GrhMMDMmGqNNU0PZXfUJ1FwWRnx
NW28672p7CsZNkZ7fFqGUHW1r8XWKi4iyskZXAPWzJ3s38GXe/Pnv2CCBpBNjUkv
BxBXaSd9r9ed7fMEXePd+88BlYbqswGf8IsTDLWmO67zpQmuZxRAb8XRAkQaC8wt
WZCaWfeGV2K95EvIEYzq6r6OK7rQ/LGLd3PtNf8rUXjMWUTbcgrSSSpY7iDuHTwt
RzAnnSOpa3zwGBm7uRxGm/KoJNuTrJSeD1h6IZYao+S2Rs0KFvH4i7CPekICe9+9
TsWfFZOC8OkTnbdur2s7OMVDoGKGlNQCuaR9O7R5UtZsCK3I6KO39817olXQ8As9
vu2z2Chbmzi/P2JiOHZzEQzBfxO8+PHFFJN8UgyG88oiOgpE3IX3IBNbEniKO7AK
uwmyl34nicD7nvxUl1/zMqBbNtB6tojVPqW+BxBA3LuBrL3H+53Bh94OgHXw/b8I
AYHHoKqZfITTykwsdNZLHVt2YktHFtC9IkGWgFPszZf1DEpNliFOlGU0D/UGTihZ
ODZpCLG47CJTFGhXIBr6T2HXOZrAglc3A3BUonGZAgdjrrLdXBR0fq2Lw6MbfurT
gQDyDspC3dr2hppDKyJfPllYUHZw5Z2x/zfeH32b0+mF+9dh7MufDx6NHv15ICGH
EYYz/pTH5snSi/4pPEJarqDPH6vxwKMLXzcJoPESnYim3SeAXS1GbrkkKuqV/meZ
K+B7pNspjajD9n1oPm4hDaUdGuaYsqrHRCkdOckZQ/N/kPPISebqBHEQgYXSkucM
NMKWjS3j6zdO98cUnZyyuduH8YmDdLHq879JposL/c2VWqdsQuG+vt177OUrcoyl
pvss5FkARgEsXiuULhanh2epNmG8bUJMrN82aMA8Q73tBStBH6Wn3eZmSPCF/qVB
eKbtlDonA0anghT24Kc0ZeMrw8QL4wPRJBor9OQXuzcwDL8NyupFFm0QZEf/f9lK
ufDtsKwjDtumzvq9H9f69KFrKmtjKUD1fRsnW/4efuQHLU/N5dWKVaiSnsOUiUMr
4gcYnY4KOWbvhGee+H/6R5TmqfIhZi96xLIWyDeAuTJAMzerUk9TLfA9RmwKX2aa
2jPUKoCRmRo1PIU6WZ0haYpNaBeC+M1AnB7AAj5xGLw7Qr8NSM13oLDtKrq+X8MC
xiSUMTsn0Bnjd74pch1IV6KH5EOhQBCbEak+69C1I/bPBR5VrfHI1pfuhfVpD8F+
tOqRw34REjGCVpPdVgxVe3r92SlhY8dWaWHMLbggHNQ+5Mp7jVlOGwOX5KdOZWxJ
+X8NgezOzNlUVswJoiu5nyt6hDa3k7LVcz3lHfFNvSui5lQhZAyD3HZxkdb+e6lL
v1D2rpPDi/OQgLoBvL+QkTb8/cpzhsjNwQUY7yd2d/+6qqPG3Ajl47HSuGUc67e9
Qlu8/XjXTiyf7ksMjidmdHiUeCPl/xYPj+pSTJqC8OrBoby8Hd3Y0zgAhj3O7agl
7Rn2n6w/rGDisDhrQMR4uktQki/AEF8vwJnoz1GSY8VYNbzH1hD04grP/9mc9nM6
8w4evjS296XF6iqtHfsmLNILzHEGnysq8OXUnYAh8EywmRsfIVAMv3GrBGwtYNJz
VlApAaaa/2oVA40Ny768hPkzADxcHjHw9FfWdRlgy9ZLIFSE0wcRwrLmGV3cCQuu
eyHT4aCIW4yYb8ddRtpMoz7JRatjau7BuhBaWw+CXLmleYpNU3c1Uo6R+YYaAjMi
1GFccZaY4ntTWSOK2D+sfLvN1sN8c6PkJlEWUjLkt73epqvhlkVLSRC2v+YaqesA
US1nRruKS/uiQy5FhfqJCQ==
`protect END_PROTECTED
