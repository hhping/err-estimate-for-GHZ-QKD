`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHSF9+F/stM+h7fTV1up8MSSqKr6zpRoaa5Llf3vr8zbXS4DeqeAIDdUxtf9WjNz
omu8duo7Wb+Z6ZC31dYK3lTOmUvwsHY75Ac1eJFEB3PlyB/qh+USSHguDL+TKXTi
RZrntUJdLN8uX/15kstboPMGSQOkcD34SqnJvE+DZboOl04PP6JPuo42pudmdHOj
7x72UOn0MWeaKQK2S9FuXVVHZsc9Ve0ZDj3T+ONvKC+aiNbYIVKkAhimvdlf/lMx
ZHYBH7LSuxmJkpKds+NmNXTO2NHMgg9ARx5b5U9k4bVUw3tMn0FwMQMUasN+WF7V
ZSowDVQn6WHKJeZpdiGZ1LBxRnp/044T6EYDwj0dwsKveFNtcav4M5ANx9vsw9dW
ioZDf5WoKtClCCQFRVgff317NXySGZDPQem/EwzN6Ybi1N+VS8tcNxT4J1TkOewx
cDzH4yUOFnlEdCvazhjbLuKcV3MgJE/l3dTiCxOoh+zqH/9NpdVv3ArLzt4Qj2B4
jBjJRQYlLbwibRaoOOx1YPQULjJZK1XjzJ18v2Dz+TQ9PgytDPKKISr4uR10J40D
ASLzkTr4KoaKOkbb7gMopZVGDON7EVfBHapeixBhUW2TG0JpK4savWyl1hqlqDQ3
KKSEM7tZu2uZh3X8ZI9kv6DjmJFEL+rHOf0RWUNKr3tM2EpfrA4567d0Iw2xzOm8
OfG3E/Itx0/0Tl52dv3mUC9rzNLlAz8M9qIpoaD+UPPeYId4WlPrrG4Fac3wPXRB
`protect END_PROTECTED
