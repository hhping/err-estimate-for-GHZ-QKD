`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfJLZZqRjRUmfN58pE33EHmMvklwZz3ZaqVIjTV+c+zobCcFVqukh5hqHXrEuHk1
9zT4CnrnnTchxbQ42vVznnwGmH+DvJFSF78r9YXaVOsEA+vpUEMSbS3JP9oE1rGP
bRoT9buuWEpfjGmxn0nPZDtsGsVB/ULQ4TsHu6E/AsxSNezVPxY8xglIa/f4vrkG
J+4zIG1sAxWnm8NqWrPhjJkbFhGj79uFVOz8sZIa79K0ohQ2br6ONh/mYQya+DAE
KlBzLGD8khARaxy3+kgIHe7T8HqAmCVXq/ytDaRJWOxvKyyYf2sISLqXxI3bZEUz
Ti19Vy4ydOoXaVYWA+9U/TKDSWqrP30xG26NHbDYi+w3n8/xBuYT3ycyIvL7JJaE
mslj8+ou7KohB90dcdf8VR4ykLE8fJ8Gpih4vMAPlWT9otpMHldPfmKh3+R9voKP
XMQ27OhgMgAPR0TNUo14U0duSiSRrP5jkhICCCQB7Q1vLdmm2mKSNC0TuJIrys0X
wqCP7XAMWPS1OQyok+YhQs6olOM+e4o47TpqTjwe5j2MSxwPRdCH7YPLk8gwHwjf
Xikfrw/XFXyElXUYyUTFuEnPSdtjPMFg+gNwq8NNN2JX3jAaMd7njM9zdLmQdGZn
6mqqXV7xRWj49Zt9cVkvZmdzd7pJzxxGKb+BMWmjS51k8K3P6Lzvmj7Qn2RoocnE
SnK/2AEX1CnUSbdHaOHFNa3CNaGD8N+DU53hTF4UmQcvoWWTHWmznPj28gr0Udv9
WGfrPnlaHZ9UXowrcCr08YD1859rROgr09FCVTH2rUjfHOkrTyUbiAXWGoJU1p8f
MjNF1B9DBcNUgPVMyVHMeA7kmHsOLxr/OTUT2sKfOdTVpPu6VkER8GQg2k3FFpNu
vdISBpaiiqbuirNgShZSSgx0LGOUSLt6AUKB/Cr6Om3Rc+yCn4doNnqqmeP7eUhT
TR2uVDhgEnwwylE/FNSnaYYlcUQEZRT8fssKVc4zzyeObGaOhrhEMSCA0zpslZ1R
xpmRIY77DQ4PIImUrojXAG5rWBD+RisTpp75XKRm8ygb9Hi7k4aSPnOr/DWd8alo
cma/fVDLiAXNle1uhc0qBD9ukj4e1Zk7vE59mb/AM+bwLuQIumadIt6DQgE1Hwtd
Vr7jUcIjQ+n36Iqd72m0vwDFQKEsDEa9tdQ37cNanmSw1bvFZpeDRSW2CtGdRL4k
nFyNH5ZCHROOYw89QxRZYt+UjWmtV7dTISjDMAJoPsFNMYqzv1g1RqfZqE0JNJhL
hDTwm5l7YysXtKTLxgQOZLuDbTnHunx7J93cCPIjlM4g+MjgqP7wi1TFQtFwn9OS
M+sMgwvZv6bKzHah9C/Uh8abiwjwQjyCCIVzpo6Ctm/NmwDnIWmknWKmA62rW+NQ
sdHRjm01LuUcYy3/l4xWLwRz2DoSKGYo41Jbb2ByGFFO0fRKQA66aiOpd5u/gC3W
JLUNB7MqbdVyzf3evX8+sho+9GLMoiAz2u7xRHqPiKAzwu4r5+i8SYX132HP94o1
q0CO2TgylULi1Van9wzGq61/1orQSpPOF1TbGvKly0ycy/+X42PRed6IWIHUbpq2
HOgQRhAFM+PRuyFvlUcMg3i7o06nxzwDrDyFyPetfUYTeDVie81FiCVHjVewbEN3
h+FVfFTyFp/t4EX3f5pE9FM1tmU0A9tpwcn5yxdv9/MfMRnWyRHBzD6Y+OQFr+tt
pWDvkh76lo8edXNul9ACLRp8Z0THChWodk9meTQ4px3b5TmtvTiA6512eiFi8Qyg
vLUvya9O0tT5WvRT+wTDFkrrqx30Km77eDEg9H+UXM1UcJhXgXUZ6SMo4qibQdok
sy8t/fzgifilqKmTz1EshgJ3ADIpzLGBUAcLLwSnxmgPW7RM4w61Z1T543vG8nIH
JdRc4AGpguVMBG+e8jdtA51olRYRdy9ckeIpn9LPbc2pbpkPv8NULa3u7KUP/ulM
Q/VzFjUDE5AyTpa0KQBBeAo5NMoKjHSY60xheA8mxROlZv/512uLnUAMdwTqnKF1
SgBGT6nT2XaApw4pO9KSq+NBNLxhxJ4bVTUtTwwftQOEfv41jdM1OefsEYQzORT7
nHQSFJZn1aJvY7v1oUyanAz+ZVOCgnkLJNsFKEAznZTRFGAoIFszoaufHpXTHkZx
abYjU6QIhPqKBJG9JFlpB3qHlLMW32gf9mSqeX8rZLm0pnv0ewQ9CD5bXQxT1ge8
48qNCOR5b/ey/kck93XONhHlxacFIRdpUQ4EHQ25RZ0dVK4A4jmCEMfYLTRDE+9N
oMMbq4rrkYGtgE+uAEmAqE8NZMYrlJg0ml7Ey91eWZz256OKZW0qQ0nfhTOyM4R/
O3YR21sWIr2p5E7PZk9fX7ye1S2DyU/UrZD4ZkJwZ1f73VZvStyQU5HpwC2MyDtf
cZ2nCANqpN3B6ALq1EPb4st+iXFMcvArk+qhLpPTj2o00P95kUFk9fUeCEWylXV6
HfVte2/vvgMWKhyI7nP9PPraX1Ok8tTNLzi9lcYwKD9zze3HZDjiBW09ioIXLQSR
RvaIEt0TTMspWsaMy4H9kVDLXwPxinWmwlGtAPe39rva7jDPqJbPE8wKU9KTr+hY
FmKIVLf7qRngi9ABDmNjiW+YPjVwQpVll2y45flfU7fWUnCnflYR5QSGEfuhMUce
qA0H4USyTX5+WZVh2PMJlDuZ+rVVUCZrphvg82vf7SAh2NRxTF33uP2gnjHvTnJp
dAlDlxytwZ4TW9r55LzkxquGXIyFMth67g87bOBQqtj102lQPIvuOesF76gunvwI
U/Oi9/hlPNMD9V0i5qC8iEA+zLIhIyh1AC9pt+gEunINixfTFGRYqByNU/Ke0gHk
vmaLwX6uixHcZmrF5OdkXDhWpt7CnWq0JTwR7FX7zTcJLIh1di+Yas/DdOxdPxAZ
sEZAX4ForxpGY7eV5za/sy89gj7z6PAnrAinBuzkGuLKMhhA0SsuYABf3mfYRNym
bMNoEMXiHzIh4EGYyTRXz2WAndbYYDsw3dWPWh83J8wE37pG+ej9mR/AySaagolC
cZ6HjPFegQ18zs+Zz5KF/76GWHxfW7WaEgLC7/ggl865ccHUpUHbusaXW+X/xMxJ
IvhF4WqPyJvUtHXvigauLCBZH+48q1TccjmWJNklYCK+eyNeYQwXmmszAxjyC+gK
y26NEIroYR3X6u+RDowjzyko6s7DCakylKxDL34B599PbZKDiF/lJfCQ+lZP6FOh
LVbL5PnKGZfNb2GKVq65EIbAXVUXPdL6TWK0lDk0xzCFEfUzE24wzj37WKf9bSB4
94ivM3132poGTrBGT+GAGqz55vSZHFmA1rLjHOg+YD2mdOolRYWh+MUypxecnqoQ
m2HtQJ9FTvNKZ0EdG08LFZPaXw5EUCqhXO5+WuKMhYh2bKOeO2elkPbnd8L6qbr0
XlLn7AEJx/bvRAzMwFxaTk5m/OrnoAWuHFp16Xg+FRSPKYMNyst1ar8f3S7G7yJx
mkLrJxVl9EKr4NLfMBHS+6XTXBGJynI9uag5WIfl1DaI+fzYsQZPryh0eBGDWnI/
fCIoRtaWX9ZNAfSMXUg6yIKa9DKXvckwGhvJMXwce2/GtYhoFcEtsjhQ9EGsEU/6
1EO8z22w4ls8CBTlQH7o1PPKAgw5SaUvyccAR29nrLMF1hNTfvSP3+FuoXP9AVDm
JFsBJFXdvCG4p0UGwJhlZ1C8hx7aaU8lqXCxBz16Ub899PpTG/eqJWaYMmwUaEf2
HTyfNbO59ie9zj5KjwpQ031wPZoVDOXKVhVJy4M1vU2cSKJ2VchnkIbdaS2/XgQn
GYmO+Y5s9OoFf9qQGuOVyBQiblrZ7qkHC5WM1M6og7s0G1Mx2Qf+lc5Dcr48BzBt
EozQExsmz0QNH8ZDwar97ItIKStLLGP+cKpkVfo72cTE4aeTUGIblPGbeJaYpH4d
LM8KaET9Bzx8MAKDre/N54el2FswUFAPuuTRI6jesz2Jesf+PLr6X9dSGuxlVvQ3
eanZfS80m6P5yUohF6Erv4C1DP8Uv5M0ba7lwP4y0vqWWKFKyfrIuTqXjR6hOOBC
N/GgWj3vTRHwcTl2K3jV73tDa8bWV0Sw215H7vac1m5oBnfT1RTDVzrSvhtHTn/R
eqACSFvhNiFyYh7c/Kts7PQM5XQ4U02enMD0C2e+zUrN8QGK6hSgamkm0lmVWPIh
/8aOndhei2Z+9beIIiUgUDNxhZ0C0vhAnZ1xNhRAaAbiQCdWn+aH4F9tJzXDN2BZ
IYAHeDj4eMwvKVFda4rUs7ytefs+qoE8dxNpMI2IGqb4HFEb8H2ucM2jhXr4DqIf
2e89l+MhZbGRQXu/EBk8GpGu6RHjSlgCsGA9jqmsRBv86DEcGLJqSsQqgTeBLzdK
IlUdE0ctVyOV2eeWRhP/SvH6260Qbo4OPnvT4ANYoTvpBl5xFY62SuJV5IaMm6Cd
2r6xsQANNfay7duziwzzrm1KOVoOT9AOKw3uz8uyMF8vwz98FBqmJRW11pv7DNmT
pjmymJ+AdJhZ59eTXT3+XxV21BZg+DueZTwgnyGRlmnU94Th9UYCnZmo3Q0Lk3qc
RN1WDneLMmL/BrWDuHoAyfmU2Xu47KO0icUsXwSOOQi7uNmgi+40VivcMbpjARsK
sXA173s8dwJqwbQwwLn08ss21AyBmCBlOW4n1LfUgwy5CnElbZJ1ouepYRudHr15
wX5Szie0izAB1f6+B/vqmMHAhmGLDah9SiD2wUVFtIpz54gj/keYZILEmbKnU7wc
k3XXI2PCbYwgp+QW6q2xO/2UQtPEZG+QDPLV/k9jmsMcWrO70A+hhR8nzJwJZeRJ
oIMrKxxaZ77wf+2W02PXxQlXm/B7UsiTgZDBZEpijVd99qPYrlOXwe0NDCCNbfjn
1NzSZtZf5cxuW8gMlYBaWGz2XI8TgQPa3JLhQ9PoQBS1ZoxvKW9gzXnYgpTqDl3q
bVZv6k2uw3o3YU6zfMpl66e3MtjzZycUhaeBJMZGGNSAFdWZQJu0k5EFnmMtjsEn
+cTyhYY6ffoffY1BshPNX4DcBPJPN4G2b3bx2hsshEef7qM4HQs29PYvjSorTTa3
JJWIRfQSDYFz3Xx9F9hHGc6XEOIRD4xQ9CGg6lG3sEC1Q3OIsFW+CJi0SrY8KqUj
wuFXoWJ9xMNAH739yijHrh/T+IgTrP7WhBkKDCNQJkveLzTQ6ifgbF3dmS4VtRsk
VTAd49LANGAe97Cq46otUAin7lFqaH5PGOuI8gCN8z/zEw94q4rnjp+3S9Fthqh9
JwH1lgMsR+3BN/Pkfuxu5JtVFEz2JfIOm9LqfHp859PIrCjdNbGGBXKSzJVLOJN6
ByCKD6FZ3Esd9umA/q2cQL08OvJq3S1m7BmPYNYm4Js3/z01ztbW86O34t5CRfww
Qb82EV81CTG3nlh9twRwEn9BMADspASmCmewjcuL5FH7nwsDb0yC5yNDka0Aau3b
G3VEldvkoZ4w8vmhaXrf1ZxXGEnLgkNzQdx+o6VRJ1mVUbLNYVCtObt5Svjhxh0p
Tpx3W/c6Ayj/jvwhmI/JbGH9C1uoIGwlZjPxNtv/0w0eMJl6n2lZXLT4swJ3DUD2
wQaA3i39278Xbiqdby1FRSJ2GUCbAjM5CiBZkxNfUk+nMlqWhqHzRk6Gi8AerUTA
w/5FeVw9YjMBblvJU6VWNwlC0OlWoDvyGNUijL4MA5WrFA67KiX3K6nJVo254Eh1
dFNUq6wOHU76lijeJ1+pX+qUuStfpX2WR05c6M/PZLcO+vkD/GF1cEB/U/eqodZA
0J0qaou/XPv/yGdKEJtpl4mJ2bby5VEjmqOoYGHpokikejlsO8t8xMelP2+KTADS
NmQ5Cg2IXXtwJgqQPLg8HoAt7/U0MHFvLfz6dtGtuOubbwyQk4rBzA53uj2ymJls
uv5OC6K2s4QgbSZRim+fyL+kqHmYxtUZaP/PZslBzHYcLFlylMtz97Xj62cVvVyt
ySuNG1mQ/JYs0W/km01h1qyPNQu0ANcdxDnrcryJqepyM5i4MLnyuj6VdtpAqUzO
KzO67kd6Q88rxdS6Kb+9T49rxaj4F+F1IAiBgIdjZNQrxTOQaEyKjYP9GJ6w0pFF
vEv1nhmgeeEfwxhMMUjpbAiZFRp7I+Ny/br8ud4rsNeTG9meHJRfJZqJ3zhb4LfE
GwPgbb8PJlxGN+qkHbcPsbyRhHW/8ZsnVIcOG7zxAeG+AzJ2qLh339nwDCZ1dKkw
cE9rWn4NCOpeyLbO/cTih7+ig3m11znDoFlPlqAxig5fUh3L8UPRvPKeYUKbVeYz
st8zadOWiP0SBMruu6QNKGXK5w/3I+pp0JvfZ+DVJNWRrh6BA69n7Q0aOF2dW71c
YplBPbnmzv/fiAAVa22U7cY5pnB1kC0H335LBqlevbTKL6eJbKs+z/X85xK2PESx
wIBqQUvqjHjmdT2bi3Sk1hnXH6ouJDZZaarAc4frCDqMHUXh/d6wmv2viy+WFntk
dBK47P8wlmYmuoVnDpfHftFJ+efsc1VSOH90DDC53NFHlXi0u2dNPopfzT+1iR56
ZwXuKbDItfSz159nw6COlT3VZHGHp92yhW4LIm15/ZE/0mX/ckkXRBOLiTWkOm8d
cUUmfuLhTrsFolPET7vM6+cYaSBSTsiPsgGw9Y3oA+cAdfMTMwfFF8IOp5SxPU6P
pr89kZjSWa+DH0Qa0rG7ZyF/HgAz5B1YbBVIEGO2ErWd8uBkBxC+mytex9cnNA4p
Zxis+A5cYi6shEoG3FppmJxodAdayg5q5ws8QiXP8AIiUVQvs303t1VHMjtjNReZ
TZGFEr9VLPRWsRTrwgOJ+17bUA5kJguMO9Gfc8DMGx+uOA6wSlQXIme1A6UeuoOq
mwJQ4NmE1jD6XogbyN2WukjdWOqawsbToSOamNyk4Qp1EWJrzHvxr7KxWA1PT9ae
jLe7BALg0AVKTiFztPbu0rgsumHTyg4JP9ew+ulny2XFqLizoNHbfpXwKR/Srp+j
cG66Ex6iGRMRqXQcS5FmSugQaxoAmOF/oNsYPNsPeshKmGpTJjBen5zZ1YW3EHPF
wQUIjPIw1UGz7gFlMB2N+Z4TzGQ7G9WK2Kk1lsbpfNN08Jov0LZTI+PShOmuXFk2
lfgTMByzRvlhloyt1q6KKYkBQOhXwlK9B3kGwfyqMF79BcfUsljm6BgDkadgWoH2
Csumn1E0zM+HkF2zQZgRp0BgCDhzxA9x6rMuKsAdgQ5eXV7QhnNMowdBpdBTR/gP
91hZtjHziNGYxEjFRQ3wo92gaigCOFYaQWb6mIedL4QY3JuUSfpoXhdDHhNv/pfb
xYAHwMYXNPkWQD2rLrdhiEn2+W9JS4W/KRzFoMY6hc7gMzT7kHohpUq7DtwOUgmh
R9GBaOyF2CbwAYXBz8rYyg3nuKFVzjMS1Dv3LPPyfBpWXABesm2K4apv2DzYoYVV
SIi8h3sbP1OlP+sEn8czj/fr9KjzpeuKRea6HqLZkF2DGwuCgFp+Xqhl0wYMIIQ3
2sBgEHKYVtEOGUIyHcXxzqvqmsUbp1dBXrWs7MJ7yuk6LQyfxmZMS6ci3It7enLT
XOj9BB4E557EpkVrwcWHMZSyLynklwVSQTaN9nwAgjo8uIO9AySiN7xJcHALf2eo
hyE0WwKMlELjyN3Rg8/qoUNonsLqsaTwL5WMpCxwdGw7luS7tWkaG33bB6e59egI
rZNOfJ7ubWyQ4qoWF4XIUNBv1Jq5AcU0KRcbu0ikqAKE5bWCsgHbipsCC6udYNpV
KIkoDJAtjXgYvRTcaIloO2D1KPOwmvOk7VineQ3zWTc1LjQwGlJKW8U3gaF0hDAW
JMJyhoUIZmyhxZ+2VNLJug0JnQJyKefU0MfYnSyZ7kgxZPJQ5lvv73XVOBpG3xLs
Scjst6Q/+PFt5H2yiEqVozryN/wYY+e89yjsnKSKONTsNV0RkYeQIHtoE/qSluZp
TWfJOayo1h8w1GsamF0eXMseNKGA7tA1dN70OSah2PnC7tur3wcH3uA6G4W2rV56
tc6MbfiEk3IWzDDlGl6R6mOcG3LrBpTQZiFrVzZjbd+bMOtLtlbHvd5XLjNp2fND
lqYC6ePNhXI05EW6mn0IM2jHcJNngFvekj+YrILiKEAQyswocmU2I5fIlawswHiN
tk4tyq4KABNj129wfgBtvgXeu1dV/wCzQdA48d8WK4xbzFWgCv7+7CDbFs/3Huyu
ADNbyk7vkTK4fDFAxpMlSI9YEKbSEPrDNmXrMFHD9Xn1MDndm65QB2VvvUv2CNW1
Hh7Ee78U4Bni/zWFae4bW79ZSBmuD9Ha1MnBbztvxR/36hhVE49p0dRZsvyPIf7k
47BCNkBTY2Kust8QQmyImPNBpueSLsgsDF1TjF4k6GBJH/2KS9/UMVrac/8u35td
mCXqvuE0B3E78ck09KsOBeF9pey/XGRVWtVyKzlmgNbDNdTntHrYDX9+Y5JuU9s1
B8SiYiACw03WuwvtCXxvIzbS93QLiLRDRqIe3i3cs7qU7ILxwszcbHzu+3S/h6Jm
ENpIkXQFcipuCo91uNGs0t+ngDFrWUwU3b3RN6icOU4FXiHr76aR9Gmail4x0jhC
+kd/4loj2aPJgIJq+zwECraup1GhMo/7J7fPwOhHvt88cCG4nIA5L8DUWU/nkifr
Olig/pQZ41oHfywchS3Ed3g7PWqJYN1l8zgr1Zs1yJOJM9H4NQOSa0eBytK4Xy8D
L+aaaSlvHUMHi8jyHrr04ETgT5Kp5wijMW/VvzXn7sq8SK30yOLtfN8q2HKEcktz
P0i5OFqB2MV9vE8lzKivSNW2jfuN0G4jv9NYY+qeza/OPyYvg4xUOXFCmclD3f0Y
Afy6wP0XfmK32q7jNqpIsF6arYhcd7p7iMldogbVuGzdaVnBmEvTewLHvsZhRn2g
qVYZNTf9jmzxaQ+4wlAaqIPuMIbs86lm7+QtuHtrWRaM9VjD0Hgmh7zuLwNlmgCp
SqulIT0zSBNQOfdlpimkfCgv5zIKIEdhdFtSErt/E+eDpuLbRwaKu6wLLYJd87ll
EU0oGZnjqd8G+bKQdTGxBD8yOqfcf5oDTzkSbMBlI1T/2h62MyDaTxzPiiwQYTA9
l2CP0lY4QSnmXZa8UNyBODVYk/jBgM9l2JR8Ek1BzghOEL3GfqMJsowCBkBQig81
lxLvZ42Db2p1xsXZkuTj2YP1kkk099dljObR2FgHyTgLPLX2SsvVob9RpGGl4+rN
4tXSom3OaC0ZtVZzmc/3T5JUUK3wTGo9WknWb26jDNNPE3JpkoqZxg2U6LbnB+Ar
Vf/jNzbJwgRNCoociW1KYebJknXSjCuigcT5YKrjxjomFIKiyar6uFyV6EJhWY1I
37GCOVZST+VmJ1+GDsVmVTjcc5Z9p38TmMGOqrJfkRTztQEViTFIwETUgtzAyvm5
BiWY1ltbn8v5LP1AK+smYJ8u+RVYkFhPzI4FQZO8uU3oubC5f6BXPRYxto6BKq/I
OCsTARljkLXXU4swJCsSof2bXuw4rV2gMYIGo7Ao9S5dkEmU4V/z3kAJ0Z2Lshby
oDFCPFBK//Uhzi0KKjNC8+IEd6OvrukFVr08apcaNezUUUve++bVKbvtU+tBeefX
tcONUmLEoziLQ5NstbVHtWYMYQaeFbxLZ2VJBXd3/DuPg6HWPUmlCA7n5FIFZCxM
HpulScFygkmayLnrF9SWu29rZvRcLij8lmBb0XPOcGcD0m/oaExeMScK8WnuAnVu
pWsUhmys50QChYEtM2aKOQKgtzrrTcOE4y8l2rYn7eUe6v5OE0vsSg/ShM9TLtNa
WTPwZWObeZYHku2Kx0rXeLrKrJ0S9omBh2n5i/RM13dKlHbunr5vzVZf+TveAVAh
M5jqBj3icl3iymDtyza8aLp3cmv2e7xRCb4NzdEuY6Yd7L63LQfhsRdCUUH818NZ
kzYalDlRQtaMHsSntgcZP0DYYDqxX2bQqIpz2fQFaRGG6I+jPJMT4icKTBN+JcDr
5JEl2syl1PMUNuMLygh2yEsfqJaVjtetGef5Ap25tKgMTMBdORwgAoItoABy/6mo
FYZDJGlYmeMEzVL5qsiLOu7SGWGd9LKb/PK+Y11DTC9Xpv6Jm3u+9kQoXyQbCy3m
hJM7ucvV+kRCBF8Sblz7gc0m/eu//Lq88AU7uKB0O7cFWQ+IR9lIgD35Ql4veGqH
3OePcn35hXDDLX9B9QmOS0GWXQpBm3Y81L+XTzhQF8TT8w4gkYpta6fGmhocn5We
0pDFupLhBt6roUkXCBEtIU35Mv8aDj3Ree97XEg45cqIk/f0jbYQDcoCrbedpJ4C
VYm/3Pngzb9HxGSmDTTASLroAMVWSrIUB+H6zlqmvYEtQ97GBOyQlX4jD6NCecdL
2l6u6YBpINadnIiJWmLVvZBdGPUjgkrwSBMSgAs7e5POGtNreuANmMAMIW0ky1Ks
ht6kxS/lKh0FK/DUEEdoZ+o1y8wrqQoLoeLkXmpFa1Twunaxh/M6YUcx1H1A0/fW
P0CmECdP8a8SnHd7mtBPyc7hw2RFmPxzs+QyFN+kTqhFlyF/X9HhOhO4Pe9Cs+O7
s6y6fO+w3qD6zJWpFjJd8NP94dybca1ThoC4193C2lYIDpc0yo3HLoJC9l5i4BsY
PIDOyV9lU6Om57iNeG90XQf41x8dQ0sYReNvdQ4nupaIy9N5sF5zLW0hgs1wM8dh
nyaiTAy6tbdaKTnJEXBLb+79j/Dy55d7OILJQrcy9fBDQe59idynsqQvKUS8A0az
hKOtNioJ6cYeQ4Qc2Nymp6+fF0RZJsvOQ1jXdFpvdrqcfKzBZWOq7XnLlR2sotrM
LYzvyLh3VT0H962wAUuyHiuaKuNNcJMO/C2x4athQgmUWYEWCeXQoV1Esk8EpMFm
w7cTqz/OycnYliue5GXdWbB8mTuQQ1Gi0jUkeTxcjR4rM/K0HwEMvLBnLGv3ZhuL
IAgT7y8iR5mJPJ2xqP228lBq+4199h6hhI6Geo+d96dCADJl0s19A7DKhGVP28Zz
+ENAG0n9kaUiF5Tp/kUDcfT3F03NUXNO+7/2Ind5dadB3Crv4Uq+JDAX94dAmh35
HQDQtloG7/qClEyw1JwqrA==
`protect END_PROTECTED
