`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6Mvmq5gVuPGE26u9YKzgiB+IBrO672gQaKtiKciEokS8DUx6RoX7FFaeflr5eYp
GFXS07XNtKrnSL4yofGyoNLM0sFgvCyN/fL/+CHElg2yLo7OnRdMNYmGRdzSLjUB
YMhRV07H2P6usD+TUCPiY296JJFqJmXV4gUSnytTBjMQox6dNhkVM9kx3QvF/ko1
jyk3FYAxZWoBLGY4BD+4fPYBTKt6lFWBtrC/6mfZcM7aACuZLxkodkHK+TtH+Ljj
CC2e2ZDXaq/ILT8TFsKbkwBpzDomr93POY3+ahNPU9BmvQpp4EBJe1BzgHaWTtvH
qSIc+lVS4A/k6XnpGVoaoyTQaR5f1RrVJ/DNKyQ6Na3hgRh9cYy3DuixlZq9wOGE
knF8H09ZG91ZHSH8AcYBsUY0+Ss8SJl5MppuyY+v2TQ4IQLZiwuDUiLW8BoLwbxP
Pvm52yetVyf60KurvDLFwrmUZ6rZ1w5waVC6W23MT08I/ETggyxrIqDG7bLdo4Cv
I2dPviA9U5Mp4RY+ynP4WakV16Tdkn/RIxZbQ3JLzOvYWd5r8eXItTSDfRQV6cXj
9KJE+M+bVOHjPJNQ5rqdQUrPpOr/5rLfyq6BCP1DQOigTjkyg1NRuBg/bBReY5bR
t4KthsY8bHjin5rikJ+1uvB0qvI+FyKTR8guLh8q13y1bydZinNDhAmNDf5WRq2P
xwaTbF6WoirdxuXQctb4H2juFETWqSPK3Z0jdSJSlMveEKltrpaQ6dFuKn5KpZiB
qkUkqYjEdBTriLO9WxwRAfKFCHy3Gcw89k9NkLEgtI91CIss/TQNbI/vBpu+DDn2
AgZmQF4CwF7Y1T5CojBNiwjiuz2jmHk9ZRr/HIJ13b8+/rREj2nPwoUvcGX2e1Ig
JOce+wcQQbthvXP4C/a+o8vkO+9aibVgFVcv/pTD6I7VnKP1h6EQUYkCw8AYg+1J
GE/rLJCbMvfGMp38Z5lIEMTR9mzAU9bfCD2pvj/s8OnINFjoSIBB4ZwGFQJdVgrB
UAYqTglJ4AbgaXe0/VR65P2OU9bzUyTHicgwL8jo8Zv8kSTv9i/jGQRixwi7MgBo
iPDl7GVji7GTpY64eFh66EgkDIU8CSJvr6aYjC1NyWjipIuq6+0YpNfnGX0EDjgY
ozxAavDLv3osmnjuVK09MoN33LQWbQJYv8IJTFz8YL0mUE4BAT73RcjOue9voKGp
8jVBbIhHggYhj/Chb3s8m5ho5vmbpyhQZRYV7eMCHjMq0cvESvqRTN4eYDfKFrZY
FqgBRs7Tq8zNLnSFYCTmJWN0EYvyQ9Gd7qFjSipd6wukVn8xFRwD8uCDVLT2FFgc
j+CvjgMNI1PcZhL3C53t+ydHjZnE4/z5hnuYusnG7NoovnsBTa4btfuh6hbXZ+aN
mCiZW+loOqEeCLlOVnAw+rjaVzJhBxk+bYl71YUiCGSG60XASIwA/pEQwHskJ02J
Nu41QwwgGppAO4hBM4NTnW1ah5paOiKa1BKkUieIhRZOxB4XjPY2lN0nC/hVuGwl
SJu+96m09s8p5BFcAMf7eGoqF7nqQOIn7pgY3DLp8krodThaPNVSAKm7k1YemeD+
`protect END_PROTECTED
