`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkAB9Nw2zso2Ja3NB+WOa1YOArIBNne8quRfxgXEBQbDI9F1gCv1L5boQktLo6x7
FoEFQj65Qm2s5/zn9imPzanryQs8FOc2JFg6KQn37UGt72pBAbIQ3XrhXSSIhlu0
YzFvhrWNwhOr9NGIat2bzdXcm8y7YOyPa4A9AJgE57NNV8MRhf9rqeg5EbekyBpx
iCXiOMbg/H98VKX4SA27S+Lt0Y1fC6vK5tby//uPlxhKs5ZFIwhImfQXPleTXzDT
uldUweX7SGEC7gCszHM+obk5Ehvl5rA3XK80ZZPbcyKgnJP7hxT7VkqMx3Nz2EQ1
3HSbPqcdUWry8rAd5byGOM8lcV+0974j3b1ERakMEZvHzRJcNlNULSJp7OoAd1GF
Cxsgh1QAeBcTg/pSPxb7yqOOIeTlwbzxSqi+qmx5q3aV75CvGfRH4GEolD2nTkqR
5y63PVSR7GBuD94cyaSlpAWQLVSZ+lWTCUUvlQtULv0qV5oIVmoimOHGlcLbc0ZR
M2MAUUeoib8veGcN5sEXymSoqp4nuJT0kVcqS/g7+s1Be6EdSEOXQLXnLV5GHiJ1
pQ6hUidOSTXwrYJZLNdqQA==
`protect END_PROTECTED
