`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11URdZ8Rzi5nMI1EfeRKXycV4XgjfdtUWVNnucqRdp93oJ2pqThAWazu6+kYruE3
gNA6Q3VtGvbsv/zCZdH4wmNh1+IvTzc0lm8+lorlF7PGGdnfsj75uQK30NgD/Fcp
hjfUJ/6QmAd4kn9WDHpPX+lAZwt1MzWopNvotlnb29qx0NlGhHbHWHdYhi6FBdLG
r8I6q3WCntkFnYzFPpvS0ptj9vr5zEMrsm408erVIukwS3U4x15ebUtwUI3lCxu/
HTIqwXmwyxXqP9oHreCY/lMlpbsZL3kvYtroF/Wte/ePjbKa7FmOYUA/vK718ubS
ADeRK1z9Qmt2MDoAzJrYwB862DdWAM8jMbzKMpY8qN6yM5+RpSxBn4stgSWQ5Dov
uw+bCKSHDGrLc/QVbyp/NtpSZryQawVQWQrzYgP9x9UrYhWUpFTbzjBt5TsryJIs
mh96qkWv0EIdOkDUC4xKfQBTeypJ/AzpOMcixMq4Eo73KyGkpf4A9iTzCLjaKWRJ
NvJT5/gEbiyjNyWNJMULu4rFa3pUwChZkhLgxs73/2xZVuvOWa9DW4ffzVhV+Eyb
WC6gykquHVzgCDpn8oZ7+s5R1zfWQZS3/ms4UsHlqBK7PCYjuXbZ36EALC7CW6m4
MSvzMxN/2QNOclfAYZ/u8TJke06eJdQO3qUIc5Nhj/ziM7EVV6QuC1GOoPjlyjEs
gEQB0I4Z+8L5xy6qdAmZjx7efW0eGxtIdVvVu5qkS6sVFpG4warlVQXPXcaPTlXI
PhqpIwVn7PwBClYLFfwgmxHJ31sj1SK98Pvhl74o2M4OhLU9CB/gRGn27NJ/KdmA
2KbR+lsLizVMG989I6mFgJJuMNoIJqAQcJMv8WXoepAFONBWAVsbufyrjdqEJDZN
rqN49jHtYnzAGIljARCANaDxpKI5FVgRoi5JqZZbO1tEHwaS9IpDb1wJAkunPU3M
YQhjFeej1nvp+NpXnTwjKGU9b2wSDRTH77cjFUCwHqB627dIewP8fRoXDhKHdLC6
noL601/Gg7CPQc0GAboaat23F6e9uoaRhEXLswqCsnM=
`protect END_PROTECTED
