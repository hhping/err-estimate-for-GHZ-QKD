`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1BU0uNoJ8/ehFRLiQFwviLVXN54gNIqKKhVwBDTaifCaI5lIRMaOJiNgUgrEdBN
Vk9MGWjXCI4uY2hJVMy5MInmUsrxxYic9LAOkUivDfDN1zLlPF0RBx7K9V0VHIaw
eduVKYVnDqiIw84lFEOdGw2IArUN0fGewnK+qONLfy8UebyVPqHRRLkG3gIlkIH3
uwjbG3VDIKroMV9rc/ep9Cxwn+b6F8sTsZ2r/qB3+3KZKvN4gIoqr5cxT6wXOI08
MMi3wJbO5MvlSwzgvAd9nj8ZoKEytQE/SvRD/4RepcXaX3LejggSVQUoMx62uItL
ycb1IkoC7XDcO4uxOYjB0pUtZRHgKYQpJuxZFp3wlK1IaEsLM94i0DUo85YNaszZ
Ll3/HtF64lnypdhIHd+bfZX7VQFZV18pzjkoAn63CNGSMoIQYqXfEUHgbDAm/zSF
klhrh+UgNw4lIlnohn35HReFifeQX7+cn/PMbzsuTm5gE87Nip5endXYGWOCM99N
tO8sj2mCidZ66aNiEvLkyUUl5KkmswvjPIKDU9pfuksni1X4Ds+zA72OzVU1Fb83
jDDijw3zK9nlFp7/Ia3loyPCd3ZpQ1yTk5Iosgs5csSBRzD0JWt2MjuqOPGsOg2d
ejhXIrPdImxm8ms8GdY8J3F1Rmszw52UsgYSBZxBmLEARJw28XXmVpa/tFE86P35
6OfUY0aNPbpFQUnZ8Y9deNDmQK/QVrySdD+eoMBG7y3JhRni6eTHiA22SclZNZa5
pgPgKExUt0h6XO9IY4jp+uijVI2xnWA/GAcZ//ihbWfYiG5JT2Qxq0nFEadVAPnN
M1zxeRBfMFfsi36oR/ZaXYSF85xCLKn1l4Rcv13rj5vYnvOPIa5kMz/DjKrRtKr5
5rxJYqzLR9TYtajXM7N+7gLzEc4U8I3UkMR1g4t8iLZR0mDyOvZRqVfytQbswIm0
5zpnjsokv5kQLfkPB5luoPZBUslbE/j0ENkC8Kojyj7QayTf7FuCehIHHqKV4dzP
0M5Qt5GeIglvKvTc1n2Z9ZaVVdaVafAVkTUxc+acq1IeMvbzRdhR67lUL2tz41IH
+i7bJTGN2sE9yZjahDnCZrwgdYqKNtN7CiExMYjfPFkgNK7XR2bCjybyg8+VlQzS
4xN0+Ztw4uqxuoq9Xg3O6ys5UTDqGYLKi8yiRXmj40e/MoYM9srLGZRHiyFeUWSe
G8Wg/SG//Di/EVX9QhLjm5F3tC3o5OMUFZWfVc/bk1O+DA9U/sD1nYhZBsqeXzDd
Ybqg/dTMiGydRfQBsUOLWqlj0hnAyB+P4cXDrFpHRQLF/1kou6kT2vph+ce9g0QL
kWT74ja3YtHb/mA8uTBrzZnqVNIzNIfqIxr5rspO9Uru9ey1cVqiZ2ipkX6sdOvS
4Sj4QWB/L5pSPGrWx4xBh7ToI5/5g5NYL7iYwgeGms0yFLI2TthNT0tT/refEawE
nC5USql6PhY2kLq4QmS+ueErjnKY6TLjs/DvJl6S8PdGf+o0/ocbQvMU1Hl9RGUq
1ZsLJwKoJP8hXdGs6b5Fs8x9RtmHk55zm/qc3ggvcYZUX6Wt71m3bbZ14oBjIxj8
6hDgbhwtvAJGdrwVoT4Q6AOzG6yUjk1vg6MN9eC1XEeH/eAHqtwtKa4yz5TB2Toe
ZbWUzGujM5/xCKaJxJvlN6mEaF9gDvForgmTx1E80X7/I0PYwdASbZm9T/mG/Mxj
zTfoMY98vT0ohI3hrayA4rgzMfsn3HjBlUeqizV4586vLbI9hRlV8BvdRO6K5YgZ
YNxtMoVab0p2EpjxLOou5VuJHucmkMHwgx0voO2QZZ7MDV5GP0h/y42UmMcw3TLY
XuKNAoqxy9zCx0DhpgXH+WCxGbUJzJcerx36CZvHphZNdC4to9hPJ6Ede1Qw84t+
h/J3SLjIHXL5S8FzRHTQwEOT43IB+KRI0gYjaYwH4CTgAQ6eKie7WDGWGrRBqbXb
lvAtST9d7h/Fo3DMk+m5CbS0t2tS0tLujh2qM06lFfJpB+02vY0eTHeWG2+HDmOg
H7nnuDzDT5rNS1dolyhhUkxhFjU2NoPexIxrd6pqvUcj4H9pQGtBcnN2DQxeuw6a
iYpbs2dQ5ZI9NCr/jXaYXhWt5RixBCtJ05jHiIurimQUCk2CRAhHdVtHYH8Fv+GV
Llbf16Xbcia6WZNS9qqRd/Xgl5u9el2k4CmfrPa4Ujxj4IPanjOAff5vf/kUcVVF
LZVCcrWjKMG3YvqCWl1TgtEMeYX/Pv62iVP17OQoricq9his2ls7yVm7+e1ZStC/
WNjCQdvN9/LeCRL1RP+c6QVDtigEvzgVMrrBMx3MAzMfhn5AYMv3ktyzzthwkF8W
TjIov7/3TCzXiT0++TPNKvRa7Yx9eURAL3AiyKcSCqy2NyQPHIclhu+6AKXhT1TV
WZZt4RzAwZePer6tnx2ING/jiBgHsHyiKZdqCTJCDeCl1SGukm59wpnEXA+EdpoG
F4Q+3DFeNWFNG+d/7+pZltGUjiu8SwNxVF4IAwiOaqXewaVqL1KcsplnKPIgc9sX
BG3RkWr1gOtBte7PnmbfCaJaq52fgGsNr/1wszZb3Rigj182imTVbbZyVgvDHZAN
NUP6SrpEZQ6FuYTrTeaARtkfgv5DST/JT25hm64xhgIhsbLnM01Bskruo+CCAr/+
gJvUttMu8SRfWR18iH7VuqkrAhrkMX0E/Jc1+dDsZG9SndBxPM9HMyRVY7Oglz71
skgNcRVdCJN6/NS75m5Nylcx02Y0EqP6hz6e9RK3MVAm0iE6N8aJ4Uzl6Ip9aVti
3IlT/Pc5kV10xoWryUwuqi8emvmK4kqW9Nh+QI5pY2GxnaQO/QxUDLhA8uGuCuDn
B8B6Hta5zaiBFr3JSDZLBKhWoVJ2s7jqb9RLIJDw+NjVOa3Rm6t+PO2zTTXH6pz6
ppopygFJCH0jWe3KpEY14YuLuuGb7LdhJNiIBOaZEy5pRrqvbV4YbNMHaVlE0ct1
zd+KM04n3ECS5FCkxbeIzPCF2FUnFfCbYx0WWo1bBE1hYxyXloAj+e+84twHARTC
DeeCyQl9kNSQSUEH8jq9j70NgqSGVUq9fq7hphZqN/udaVfKE02QtQ/9dPg5kutW
gkqUh1S2Fgee98BTjw+/yHsyrkPoxG0HCkL9QVf65o6H/j98nWO3K20cpyK3ltpW
nbd14hRNDdGOz5YBRVB2DgLBuhfQ3PYBRj3gdXlPbfF14RneVyAC79kvpZj9rHJL
rR4zeL9B0Y4RfOYs7ViC2E7yaTatYKSANjalxtVCdDxTHf6nEM+NeG6asG36T550
TdAwY+d/Eb0b+r+j5jsJMPKEhBxXMmxAfQ2KFq5U+++YKZF/nA8FNozMk0lebhcj
LGHr5hcEwGwxYY2sLNu3CuHK4dUdVm+yxFtT+jJj4OMGaYnkQ/PW4k3tXjnJkvpB
CGpyDHd99IS/DOt7uumZt8GNQQBVjUI7v+NYW0qTR1eMudZh80qWFZWfsHBdAtGC
F3Y0PaSnVRHkh03BLnGynaWeFyXICzTl2363gU1FIpADz0nU/Zkw9qPIgkLgM4Aw
VkudmlxVt/ZXhjKFx8YBgtelgyVjdNJ15YtknIRP729aIfNbjM1LGXwa3++aIJks
Gf1GSeCF/btT9VB1O33qgOvkSRzGgJkGorpPgxdyCpK/fFJ1HdCc3eZW4cfJbI8g
QsJLqkxF4SdtpEfd3bWFUAGRBEOQPMcyV+yresO99qtK+qdxALTCtn6HgRU5Undx
UfFZu72H3gE12r7UXF9u0WitPPRyAnCEWwEMvN4pKlTxJ4vlByy5STW/2+aGQUJ8
zp15I6f8m3cCarlmpvUvmfdtPGSvZwVZPGoGTGLNbOiqSWninxoWMrG+jt8WWhea
/ny1wTmLHKfLpTB9zGBJX2xdUO0OgK2h8STztuhNmu73HJcXICOxIQ06twTyWAwv
r99EewAWDTPsIGwbAPKDqiqatB+OATmN2X/YMSTtLiR/3TuNwEHWc/86j762Jgu1
2AK2YJA7L8DW8SPQLU0oMcFOjpYm6t11eWWb/6U87QZE9piBHZiTJhzkSMciaKaW
VvTMvAzXdibWrFKQ2VexH7wPMuAHnBIVupbRyxxxH4TsT4yoEPTNxwv3WLatnN0x
LMfbFxvI8fx+e+ufuJ+wbkI89yC41TLQHjA0cYX5BHnULECLpZWYFTMpnGZiHxSP
oRQ2DfRtc5B7DEU+hpgl+A1G1++DXNtCuy+8/khUXU3KN5ouhYfzs/EHXkrdiz8D
cor6pNNkSiYDWDjmf6z//c3M2XJtcQiLpbOB1+oUS02zPGHRUtf6fzcdcAl3grHm
+oaPqfTNljNtZYCMnYhOmV5a6JRUF+5tHq7qICuC7xfhkANhOtM7VQ9SuqSZpLXZ
9YBuhdlSmv61bCUDPGAMAz3PEHO23g7tOuwJ6pz0AdFnOU/OfGYRPTHpgNV2yOqA
VA+OgGHPNmy9Q1wXQYiSpNTgMAWbxiWvrgtnV7mU5Tz2wzEggh1AxVX1eWJzkJ0l
BX735ZE0ANPAfzY4ayMjr5hrI2mK7U4ndOrMlt5ipEfUe6Nq2Hbdai4eOy1E4Kwc
GlgoeCCNZHMo972MALMmBzG4IJj/ZwKAzGRjOIJU5/06cgZvs8FcEB3OIvc1l+mm
j9r92cHVCmYSn47/D3sq4xbAvN6gdgJU5TUoRb9c/Pgudgi0t0xdPFGJNAPLVH25
VkHE1hrxgnzVwKBtuw9ubeCs2s1UqYygBbwH9hO5UJYSU/ou/Bn960AmhN40+w+l
wWUzCRxiknVOYvv6m7U1u0ySoo0/dL+i2KkZaEeW8edqySczmqcYmCOZQudtAn+D
bkbQjQJqL9SX+l62Boh5Ru+Pq4zyWbm5/1I4kHJWL4CR8DfHAPtUI+lcTNHiFAEN
hz9ODKVLSoxdWYbupU5dpQOac30g7uSFgds7BCjlkxSLF3/NQlFhMTZdZiNt7a8I
iznTaM7fFes9mDT3ZvV4AlSffNwzK3vG/6F8lZ+AJMeHRj5jV0Q9DsY0iXoDcMM8
XITKJzDWhs7EOAmddEzT5ldDxvGia/t2W/IsNNQWaH+hkkh4lwjXxGK0g0CpY62W
bTBxI/PLvIkxl3bDK7KX8ktJU5fyIFUU0evjLnorDxHvqrqd+TkWifXasW07bRNL
rTgiu1dLfpPpg5HLlHD3BrBIijEk2UGRBQmCZMd+GKdJ2qst2QUlcvDhyG1fx1Yh
/+XaGbDKmfOFWy5UN1upDEYWMGazZCMZ7g2IgJcZKi9xuSurFcx5TBl5xMX92xSj
zlfXMGLELWm2u2+NeEFYg6J9Nl/tAOoCOPGO2tAVUolDsCGTUjb9Gm76BmVKDLTC
NIQsOeZByKLa6A6iCxvWgyTLqY5VYzoUtti2de9vRmMRLatu3A+IzOLsTRCC2Yfe
L4asWbwsp8Xt5vFsvyWoNKSBlm7mVTmDObB45TV/HViy1rV8LHh/sJh6G2HkmKTJ
3nivXLL9fIjEi58dpWZydhPIkyH/Q32UKcBRDvxPfI9SXUttLSbR4II1ZvMTDzNV
/erCP1KMfBbNPjWiHaglLp+1JoGqjGWJtNKbd3QSiz8lktJ7tCffrIKQt6xaP/nF
qKyPUDZnh4JCLzOdHRavOS038sLagmFx8bAfNHNVNYPeCm89SkvPt2FGmcincPnb
Vy3WV1cB09r0HtSIk0InxzRiQGvDXoOmUlGlofyxSI9mc/ucm5gfq0R9UoFL706h
PN/fptGCVum86xNRddPr1ismBBUR8E+KZmWQpywiS+dSD7dGOCI6xb4A5r5kAFEy
Ka4l7Zvp3knzCvjGo2I+UPnLJRUUzNnlqpgkrubI/EQgmBUJEHZ2On+338kFCUIz
ixAUwnVrpqJ9XiX4IKUN6yLEFKNm7VY60IEXbGEVWk1eWGcDHUAiPG+rcAQDszXW
7QJRbMper5DQ2XPAeuJy7v1YYrzXA79Gc6bVafxKevOVnW4ge7+F1EsTUswwDZxz
DzeQYzB8X84wEGCxG+qJwFPKdWdCAKU+CkoDG/Db/YaScdGLSdopcQTSQ6Ho83NU
uOpPnEMi1gkFD3Rlkz1udOkPFJVgqPOmg/O6ahCKBrdVPOSxccwMrXbFPs0m1UGT
BsYWaegbXTSkn/O9P0GMo/fgNl/d1ZfVOz1STEnOWpdzjJsfu5hGcnFcJpCHdSo1
U+DdHzXFgjlBOcEKEm5QqHQGGQzjmPkso/1/GM9KytWsBxtINs+/VKFgF5VaSIjq
GDK2VlKJnNtcrA/BevGJNjS5CU/fYERRviqjmGvdd3uZHY6knH97eDczZNQhxpmN
x6tRXlotuHPzSrdXQUyKeHfww7GUv7VGV1NH6GZOGZmXOX8oQ7xrkYXkRcjXd8cn
bJzvYAPO1L2/UdtrdTNQq03AuLfm7e+QFYcM2KRuXszHK26zkjazorT00JvrFI8M
zKMZKPi+FtgwYHnI1+G8anLl65X/k+kerAFkhy9Z5k8OJ/xer0202CGJdrpBkVNW
pWbSn+PF55Gg8iAqb05c1m9j3SdeA5+WRYN3+LuhMG9A5bKU60o39FjgrMFcBj2f
UX9JIIUgEQjNlOrY/RYqxodSltHrkQoonbJfRKxRtI98cO9z7JA7DYWoEPN0hyj2
29M9MXlWrfJWfzsOEYBXW4R+C/bvfr3nc2ag5xDzE/rZauakdxwtq11P6Oed0OTU
3CNTc6qpAUPKWWM9DjVHPYGaOgZJNrEMLPmygjJEKmOajUC2mAhFlIUZr5cS34IF
HLCqx65uf2MYovkPNOarNLL1Co41eFWQ+vg7KTjJcrltR9WJ/d3OmsuA3TI3k0bY
wvs5M1vOGaPHOmLrjlrIUMT/CnzTQl7qAts+78XVFI4UjAhuXKEF1EEkn6SFqNIn
8I/YGp+spzNRi3d7cVfOet7YZiZPLPkCJWktFhn5KNKeueXTzGKgBtq+EgpSJ+HA
3Yee5LuAPfO2DbXIKksNatlRMGQuO9i3y6IJriCAkuRKBaUwjtPWkkMdavL5U6HG
DRnPZ72bZzMFqQIqEh7bdcQkg03m/NjeSCTp1HNZD/3yLzZlbdVl6loq2KQWgvA3
uvhX4jMON/jUJUm085XfQLPzbDHguXWpUVV171O/kD95HyvdLdOdvToobKtKd2gQ
bLXc7ZbKAz+E/CKPFwljFI/1mtnEwOGFY2q8GyY4VGLwg1JW0wVKlLHJW8SnlxSC
GxdAvQI3LHf/ub+Q6RTuBJus6F5hyngay32zNFv/6lDlQuyea5oMaFT1agR9ZJPI
4bpHA9DpxF1Jbt1JoQfrJyRyHDl1OSZSuoR9IOX/hrHODqZttUmhReYcfZDNPURX
ZmtMwOOH/1oe+4cgwsTv1jcGsh3j8d6NIQOz86NcoCfseOmplausvr31DKJfUIrj
vJoShYHstLzm3/Fk+4SIqppRLgYqym0DqzRSM6croZiU+el1sjVRILNwh71+1ZMN
qCVr8fPSaecBIjzLTWa1EWEL+r2g8boWxEdzbe6+NExRGGw2Tycq5+KE+Gf4eBbn
YV9OlscDx7yiUHT3TFZLOCIaeCLW2SRrjUxmSQxbjxgXg+YeDrd86o8Mj3ysdeUT
/cnbX022KKlTFLxEAd8rJ5wqXvyHo6i4Qlj4mASpttPyMzeoDvjIGEQreNMVsbh2
mEAzR4XwCw0RwuqKn8r1lzyG/XBhA3mKuI0qWULG+hIPjoN3NAZPEmQvOUP+HzVV
f/YCatUCjKCApLBBi6FSehLI9J51zhHDWtfu6KdlwARLHT2q9zbZ43tgRSkl9q97
25MSUDSzRRE4PxdUTL1vQvmRxcSsFkkNC2C6Tw2HxF3YtCnxHDqAUd+GI/8gFqnh
r6dRNCiEEqlMigRynGV2vKEiH+G/c+fv1b77W0lpVvcJFjQD88YolQDUZE0jmrDv
jTqOV8XcdwuR9ecCJfE2rZcDGBs4F62k9QdqlErR6hOnHDz0zHUhWnVYTCR35kRr
/OwIcDuV9dHyKJRBLMT4ggzBWeyj3+OMvCQ5Qm+BPUxHnJZQJmV3mWQH3In6hUIY
4ItcC1lQD13343K4UAsuSs+W8JLJnvELyANIrldd5V5dgRy9N5AqdZKfBP0rR64D
CBnJIZGg00//fsfaW2slONaeEO4SA+9CaDGzzuYtjItjdk/hHEbzg4egyWI6eeup
bgAXfveBMUKpjY/oNzFuFv4nzccpGmPLMYOUm1Oa+pI=
`protect END_PROTECTED
