`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2bcX9NhfHbB+narpxdlOdDl/2cNTqnIOzpx45uHUUbvi8klUwiAV2l1Bg3/Fq3p
IqcWfz/LbkRjCznbYeczIJjgNHV+5QCeoYt0lGGdCndsAWMop1c6IQ0mY2YDVQqE
4swmAVQxJFqcN3gbgU4iVDOkIQ4PafWd+gduncIp5r+AzIvJ1DY3j0uelpeycdv6
3E27c08wkQCaaDwVYJe+/V0jUL3zYUsfQmJ4DIOTpmxLP5cj1REAf/ozB7ZURA90
fxe4LBpw9N42lI66X3k4/9slqup6CiY2cp+ijAS17ukyzPtZKpeCcAXIrdNoO6Qq
DwgMgG0jppkz6Jeqa8OU1zLrmj3CzNkpkqGemf2JRFJRNeh5EIQQ2kvYGq8I1+jo
B3Q3DHxq++WE+hVb2B+kvEYktoTI6taZ3NBmss/vf4k/5V+NAj8XCnDhnZb5b6F/
BF/4qpc/3k6uq7FK2qmM/QibxwjnfDAhyw33ahd2OJUw3Z5g6MND4XxFHM4IvB0n
3DxYyhBkdvQcGLVrtNWmxtYZ+U3RpSdu9/ZZS8P9V5INxI+qcINwmEjD7ZCHLgyb
AZn8SsebYtAvYpPrfa80fam945pc8kx+Erw7NEr6qvjaZZQOglBnHT8OFRNGyqJf
DvwGqX/cXkiVgb85CS435lyAgOcDrYT1tZWCYDQ3Xpn/UPzf9jAcMH2ELIWwWZZY
AeFg2Zy9iDBrEePGfg0SJRwjumaMVJ+gcNCj2PdPU0HOFz2/P7PLSd4TycDDo+BB
fLzjNIYusYF4OAVSLHuVXmiPjt+75+WJ3KFhPg4y8SP83NCx4S/TwU+xatI78O2R
unwvAgTXFR5UnNdrmm1h9JR/1ZfcRO1VmVXZ5kwWHUQna310zoG7/zJ2jgPcuemG
edtGlSghXyoNbrJsZHMo5MnwEtkt9g8vC3CSU4MzplgF8RgozndBRYByD7w6lBsL
MRswWFRodNyiAiOSCg/YIIDHMryU4nEVjkQMo+xTRG5sGmbSMIEHfZtg+k4/Kuqh
Ro6SePN+22I7YKeQcycE/HPp1zy6xARL5kbfZYJoeJLG5ejQnKnmZUgkQNwIQThB
bVeDMONNkdUGGVZyPbh5hpAB7nVeSmikxiWe02UZAWQtMf1gY0Rhm6giOl0E5Q9A
ctAAO6tyB7NGuB1LhLivnXAwilZ2sVfcBykvzBP3HpU7TGkDIzBr9vZVpRryivKd
TruXVPDMXZmOJ7ts9qPR+n9zYnTSO10gpS88eSDVm6BOPwk7aP/r1jQ3nUpR1kKc
BHlHicGXA1lowYgiLdpR7kpskazm3RxOgJvTtNTI7zpWvi+pT16GS0Jx6t6mycCf
xksQSFA4CfaQ5VCaYLn/TPhKg+Bx5Lxs4prwnWbC4Y5tSFGtQj54SY9xA6fRWYIr
YJaHsdTiqHP6wNIO5UUrs+pJ4bn0Ywtx+k4elSTpghcu+ZXRcy7L3ucnY7IuEUVB
ubCqEsMZXplQcgzfoOVxj+6+/2xyahFhaka5ocrET/faKE/4ThCJw7HvZixRPnEY
mW2Vn0FrQ0wSxKJmp7d7z4Bfi+6FNwJLOUvnne/HmHuEdBFxBRK1unHw1/tcNutc
AlhViTjEaXrKJZvCt0QTPS/MY5P+jzDQohRHEcBZekwqT7xvzYLATj1VfooQes6x
LSvhDHqwg3Kyd8efOk4V8udjSvRctwnk9XhrnP7fEAOV9tCDKOeuHX3JycQxYBbe
b6TxDjMFs4BRfXG6YYbOxhOKcBkgkADP2sOXmZrGHpb45VMbEo0y0aiwd1oXmWXF
ieXzXCpeAeGpSDq1dZRNQQ+E5CIvG07kKFJoNQ0EzJAEf37mI4KhC3imzQeihjhj
QDZGn/83UTqIoyMDg55SHtAKKaP/yDSsCoub9P/PIwuz/Ew13IroLGW7xEP9517/
WQE3vmLgA7Q9VSOXQ/E45P/ReoPmeTySatFOblHQr5nlFOayxRVdHqwBo0lpT+Ur
kluikwKKFOWdCjwMg1JpqQ51mJfL5v2NqLLHA1DG4XC666rvelOcQLUo60fSruiV
xKOSq1Odt0kvtAX8BylHHiV5oWBR1eio9W2zLHtsiw45gqFC47HAYZfxLh+YdVfR
pFfGlPy7U95982TMJjJT8SZ4OkNN4yLcUJDnnlDYzRpZ4zPpSlBKq5n68S6ZvoqQ
O3tfrnGTL79/64p83OyOpIyAsokQf7pVOYTsRv+/EKqosyljEPB5LDFFVWBl/jyf
pIfVTkYUoJjE6Hq7+cR8uCeFc7kgjXP1VdnmhQZ39Mh7lapf8bkS9dRdJSA29inv
EPQhPLYqVlfqESsRv+tk4xN9CX+MRf8VILvfRtcZCFlNXDv9Rg7OJuUPQFmxR4Eb
uquBIBNKssCF3w79fwnTvooyUbz6dTnKNDYhYx6hyF7E8ldwQNBRqau6LXd6UQph
odlrQT4gaukmR+fs4MaEXR4EVfkDbr87q7f7u1I6pRzNgmpjkcni39ckPPFAgxiu
6I/s7bwOSOd5okRs9JfFC5pCZOfvQ5QmoGyRac0c9l61rj5OpbLVxQdXmM94EvHU
zm1Cm/dUGly6U56fdYGATeb6jTwfxjp87hwoBRD3lZsva+TYGXgkPKztRVYFdEnm
qN57G/wgQ5jrD8oYP0UusTLYoz5K3CQB1tiF9QhqjFB0EMg92vwHXrh4AeyiNCRQ
vKGLUBcXYc/f1CAZ+X/296+RcysSoZHuSybVNEl3U62vv60ZeSrVdvalBlqEu1sQ
5njwhR+T1IaU/JA2Okc2ZNa6ITwf40DKblaHfrJ0oeBKZcbi7l9nusZUhRuBZh1V
a0NElp/MBmwI7IellM6ZdZZAJ8Een6jfe+g9DpLbeFVYpbuH22MesE5yYjM0kH25
McHKNOKwg0wMhBDSIB5o3WR+chTNOLTHypEfsn79npo1lA+67Ubsfxl3VHPvtGBx
ewkFh8eay3eDB3+O87PZjHFKMpeo2nZwv02/dKBjaSVkeFWUiTk84t5YzQYBIUnL
MHC+Q/7JiT+YM3JE779cObFVShyTVnHXfALYMqKJu5r64am1lVT3ywouSdC5haNA
EEZsZBkqI1WnA6cfBrowwqjOJlMioslcePAWWWPjhQnRze9e2+UDPrk9IJlIMAk2
La0N7AX9YxthkN7hkzabfEnkM8HugbEgyqISXRIfelOPtcHPhj3jrnylJmdsa+L4
JnVkaI+Y4UdcbN1MUjPGiIPC3JHemCNzEfWytZa/DuqZIonW/xskLrk0GQlcoV3v
eoqS2q2qJ0jVATZDOVzJk6xLFcNM8Zj+c7oMTOl+MMh8VeIy99fKMbh4kQridPwC
e5lmmQlOWCXF1T8/FHFk3i4SgAvpLFT/ZUQ2XqsVLpikl8T7lNtqJ9WQ/muS678L
pMd77KyrQZ8+ttNTZ5B0iNbubfrJ+HGmGRHLYR73wjBhG+ZH1cp/L5hwWMNtnDG6
B8j4QTwbP9UojUptWuSDJJY8cVW4LdURGMXhmVQuF8g9lIXanqLjpzWfNAm07CA5
n/SKJ+9eDBhiQSVqFx1qU+JCzC9j9jFzqtjrkLSKdrhjurs6jRX3zanoOkiwe1zH
3nmxT0qe3zf1tZvQrnIxVJJDL3MYkZ1GhfcVexWXxJcl5XD8C1meHNNlDkmYBqzu
G6kFMLAetEInD9ERNWlffOdn0DszeCWxC9+NSYCAOZDdZcFlNa5IixImM+6fZzqg
/nXhRwkGCw4njwjqxZUuVCY6xnR/0qvYt3h7WdMSPisdQbiOsJc8WckikOyxekdZ
hNj063JIxnRgixCnpfDw4lh0UJslclS701KRBumpLsd3GwhUbKgZgUoO3dYeCLYJ
53SnnQI4ppQKclKQ/kHAG0W/VLtMQ0zjXDW4REKwt1EhNBHLhYqFsfY0FOsIkMsk
/x502s9JCnNbymBZc0wJHQpEJoy8yfE4uw5KSBVCQATwLP1gHz+PXM7HUSvG6XoD
eSGPJjk10ErY2tlWBz49XsgJQCnhk/NpHeUTjY4TfzsM8z0Dpqn6h0m8d+TE2xOJ
SNFERarAeRbVux4JAukpaA6qE+tgfLN6b9d7r3ptPpS9x9febmlsd7h0x6ptZJx6
nrh3d62JWrn3/Q2bVg+O7c1dqWdjEChuqBGx494UIPFx/GFc6mSoRFaT2x5T2z3y
O57yjuuYuqnLZkdnxk7qD+oxpkJ9VJc3rtkAHOZFNhnwYgJJbYYy/A0zIkeADAY8
obIoMkaOVbGeQbpEzVQiiUF6//0g6nWzkhe6KkL92kCTx0FeJpdMYFaAhV6rli7T
28Bwu+RSZ4ZuI9d9AI4WTamWTLhpHE9YPBx2T0nr/OiegB1onJtG4ikJbI0YS8AQ
jKPELfd6Mgj58+xkARKYd3h/GAEpOjGF27iNAuMFYQk8ucwd+XuvRpc4NlwV0Zqo
yMU6UF4vPgKW/Ga6qnMCvyLPlKaT9vBegIlvWIp7lEEciFN/NBd0ilMs/exPXXa7
JieUbTMfZH7iv+xbE++uELOKtKMrohUo7Gc78XJ49h6sFVKSWL4AcIFszT3qRxIL
Mf8NhDFxJ0jZzU3xYuzDAv+TfzKaoOLiX59OMcE59ZHhFPxlJPdGVkOY+/1h1UQ5
tw0Rk1lGvQPxRwnDBpBxc3e4yJ906cENgxYS5yjcXpqAt4pBtALtlaxTKCrVjieZ
BuqIDLq6wUCbpErquNmzH7DYarUxDxn9bKzIgz8zyeooZ0FOPBzu1fqsRLl22oLC
Rt3zu39ZX0O1y8fRgk05qaCaKfjfRuMhkvFULqwdf7+Z8kYfGiktxfsuB2Zv2trh
qjMpUzzN8nkJerA1u1LkoDuZ/KV9hQN2M7LYPqx2OdWmK6aTKto1U0cP7AFZQlaR
TUauI4MInwt1VyODr2W24rK4nt1vbPebyoWTJHr+SUfG3vLAVh58nzMB8TlsTiIH
ZqB8rrlDz0lF9NXL0LwZnGoDXQFPMsp1Uns4vdakgg1eAwqptKQ9xL9X2a/oMYuX
tVWUDjUM8OjjOUf+ctQAjHYdDndtvwtygWjdrbdvjChbVMDVVCL6pUWTrBNxdRLL
StkwGPA/2vUEb7GE9Xz7Zjam3Ia/O7TXm2t1cbMnrh83XT/Nxkvq4mDTAuTEIndc
uUzYbmt+wtiOwbWOcNcSmQr8ubQdzl1tbSaN33no7ICUu68IlsRGmup0AOcpCQvo
PYGsvAu1jZt4957Gi6f0OJVNnY1m87RbUW5YnD9dKNKQB1bar0IcOjOnLdnff/sW
PJIDYXfCBh7wE2gELB2eY+VqYtTIHKiTzNuyt6I0aP3BTLjNB8o3a8pmVStsxWwS
ut0N8h/Py+2UtKentnw1OGKebhz5mqYfIEwvLXSM8QjAaT+qER165q4W9MX8LcQK
5m1EITij4HJQNZFUqGkFIJaq49c3YF+M77kco4xYn3KowpYhSOEGPrgDeEXWLwX9
FvSzk/emf/pMoHE6estFQ6cMzlf/CsKjB2R3IkHFJ7dA2vHSjCGfOjxl2KpjAgom
q2L9lmtAwturgJ9y3aYQ5tHHF3aBmpPTchdhLeg6GteaAwtCzkeQ9ab6zBwzcV1H
uDmsV/SsULetJONM9Hxup4VSVJqSWBn5wubvrTSKb/3y2B0Z1kV0vxut2LRxpj4L
netgx/KXls7vz5s5kIe1U1OtDvg/7Zy5nXcrmfLtCp12A3lyrqFYJQflWI8J9Bqf
meRz0aqX3q8111MrRBuhtGHYbJUFiEek+etGBnYFpd1QMuPrY0QqdKVqsAEL8jrd
HSgzbb3XihZ8Z8LXdSgXMhPF9Y5nBvqxh5rPZfeoHeZP7MghFjww/tXdO3QeL5zt
y+M2Z7Dej3nRtgw1c3E65xN1ZeWn8EW0hm7REGLOslRLqhbAbSCxzft/A9oGKg37
IvTd+QdFNm+xNpTY0WFOINRrTwcwkh2t/4W0a89/2xOa9VjjdgN9nqkwoK9Sj2TL
4p87vd+u/CYt6kH6fKs1yUf8zdZEnhfvLr7DYbj54geJ7Ams1l+YhTaaFP8+B8L7
XuB77sVX3vEjdMVCxQOW6N2bnbYdmFNjftb1w+Q1PGV4Uf0aF7cvruQD9n+KyRQC
yo8kkorGsjRBv6oUcw0iRsibAInV2nZQLk02WowkE/gi6ktaAtkYdvDSiq+Etk0Y
nFQZQW5Db8C4JWYl/xPmyzpNL9AeKgbz6COStv1NHHd5kpG/QCeGzKhgEgi/+S8Q
BJW9Uyos/hUURF9EkFG9ZsHoL/OslQZpiIdpsUrnKzQnQmI70M9r4TcUKlZUzuL9
Ywzb6hVpYLQ3b3Q1TmyqPPGzUWhF8b8YaAg38K9mQ6R+snn6iarMtY5WAAWF44hE
OtDrI5sDf+jznHo2oC1GusZWWV0lQS86Yubbgo/UmZQR8Ux0fsWGT+4b37MbPmFU
UpcPRnXBqV54SUVgWwCd+DMjiGoWowNSdIRnic9WmgpAz0Tr2EVmXvDa1oyRU5jt
U1tvRMGeL0jglmicUKc1yB5EMnNCuRGAKKv4v72Nf6tekXakloJKXZXzLIFx49x7
i77gZ+1HsCnN6S+l/she/AQOHWh3Z21/bz8vjabSZ65NCTvUMYpc/WGs5Etp/Xil
4Ki0MZ0rOB84jMnTvj80EFfNjtiHOA+053Azbph1C8E8dHP6Wqzwba0kB2Hm6TbB
ViwZCDZg8iCbDxiC+xBjbfIimwtN56R+ARPMERJo3EvvQsYGVxsV+rYS9voanLwe
2F9t7PSz4r8JjqFMoHzqoZ6QNVX8d3eePR4aUcIj6MCLz8OBzl1SOC6tI1szR6No
ArcOLsaBDFk8gAg9YoXevcgF8DLgQ2f9G25bYWnrKsjnzekuSRfuCvpL2DK9Qr0P
OSK4pa9BA9aC7Kq9LW05sGpRlyib1uyr7xTaC53XBb0MSLDUt+gewyFqT2gwjUgG
tYABqr6eePdqeHc9b1g1jeBozRkhLGFEJU9Xv6C9izECf90rpgpa/xwqwYs894UD
tRXpwQRRdFwCPPWUjdgsAhplrsNYu15mIwehJbrYPot5uOVYucGXIMWQ9iCy1i8W
f/WMkfleO5oU2o7xCTvwZa61iXRdTODtHnw7TX0rAPDlEhGtuBYy3LoX5W/lUU07
M6taWZdiMzPmC9nZolB6D507lczdB/7ux/mRxIBnxbATgsTR+cpuLdsECCM2yMwQ
xG6YtXdSvcCy1kpjP+B6sjl+kYpCT9rQPaCoa8otBlma/rAFHUsNX033FXzRvy/W
0xktqeJT3jSAO3KgA+jQKTCCFgn3heDcBCmiHLnCsGvaT86y/J8WhFR8nznD5Jum
xQ+4pkYWO5MnHHMhXtCWP1pcLT1n28mO9ysKgAo0mwU8g9W4ELCkyt1hROASq95w
TEWaoAUweaOUjXQqIbQV7ux55RDEpSQchCjh4f3MFva9DXo22aPjrDK+yee1A5+1
8GLO2+4ArVUJajX4UZi2Vt31B+eHqTgkgivdVNzLY1TD5OLVVaT/79ZyrSf3MMC5
BNGMARMF9+2TWzMouLgTEzrl6uRCirv2zTY6vwmapOs7Oy/PoyyD8ObbD1Lu+xLC
f2ZZ5Nc0B/dtCd+TrSnZIvbjBD5XiyyhtVtYFWDMxDcACyNarBXZ8ebpTjNyQyUq
c6p2dV30rCGGBtQVYmn9dIlonfOlZ1Rf/JPxswtcBVLju+jj/o1gDHteqFW6JeIm
DJ/p8kLK+/mPh6Hgo4jVNEAd5wwEPhBrUgyRvaddjwQLM7oUjk6ITF5eQkNIf9hK
Qx4XDhfd01qGMZdEebpWli6MCj8ZjJI7yWyRKULlhG+J84oIy9T9y2OMaeTjE5qf
kI4nZFRHgxPOv4E/UtCLcl1PpAUQOpVHuW1ASP69PnvNFc3zqBlVWiBf3koEojuy
+h09M1X6HctLBuA0YsQq0jX5bDe9EIUlG7TQrOe1cd/ZBDvBf2SzlPib14eLLPOU
LRNOO80qc/aqKokKiFNn3ibGqd8Jov8iMupYAEW3FhUpPJlFAE8I75BhMGKeXmnF
uYLUUW1S3+KzasUMVy2lga1x5T5vEEEKrScC+BNXJknouEMzLEe5uOOGlUuZVpzj
2L4tS013yADbdP9izCdBDpBvattGhHJ2Yg/u03NV/kfpLI6HMOF0gb6wRdl2qDoE
NWYNahci3BTWzwH8Qcy9v+8d3b7fszKOQ+O3WM33cZLObE3kIhHdNpxy5JdGzr3x
PZkmGmocGYF+sHKRCoCq5g==
`protect END_PROTECTED
