`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34NWNg9aiXEXBtxaLVehFVuX5sdAxejezs8zOSw5lRAsalJeIFy2Pj+hLXtXoKv1
K72kZvWZWGyIMQiX5UOsJNqWF9hMxLaHLSHNX39PxpEWVekc7WQ4qZ8h2abTH6NB
xcCvzbPmy51+B80bfaCHPYkGgnA7IQE4SJx4ZB/WsYCYMWv8NzsDFy2Tpo/xmh4L
JQoODHR/k8marxSzBZdDKbugzKusBgAsX+Rn6wvOBr+x/91f12EfY//0PYcMVNfm
cxCpiMzxgfAvU0OzcQFv/K8wiUQI+RS2SYC5GVqsSdpRAyg6jiUheAJT4tMEKhXq
rXqUJ3oOJtTzFR+R+AJQGk3XqTF5U+aGRPcGzgAcOQAwkUWDoAIbM8xQtsjOcXYO
Z6dg/g+Db32ljy1YlBEvsqMh6KUTgGBf9egBENZ8rRr6vCQaxylXN9N28w75s2Y/
qCcXEXStIhglUpYnP7e+aFA+457WHdofrv3KScDGGYed21zeId3sIw5eCCeJ7FPT
JhVT2ZnqDPzmFKjnlkR5GAkp3laww53UXNOmL04cSsKvC3teom03NwGa37s/BFRk
yZ8gSnHHLLBbP1mXZ91mtvxv7toDQoBjYB9BTpymTFTDYI0k+OUXyOsO89ctckzI
eMt0lqd0aYmS82PTp3VOnSSbnBg1wbiFTcfP1YckSeBFFc0mSN1hhn5K1lFYsjFZ
TdeGdZ0TxVJKyN90uYz9+KM6ilhWSnvPZXTRLTVgDH3fJwvEZRVICRKh5FwhT14w
fuJyPmbWXunOPuKhSYKAfTahUBt3+0DF2hWONKlN6pjR8815K1lYy/wCK8Aecgbh
sVm9LW0F/2JurnICum3p7X2xItpiiHqH8LCUKBOpwGd04VY9STYcN4+T9XqxXJde
0QEalTlolXotIVAzayk8JJrBpD6qiup0ynGO2EHlN4TZS9AYFWXdj6XViMLa4EVk
0OICV0lFhaciUi/iCSxoPDM+FNMA/CK91JA2Oe70LuYF1BUE8w3a03umLWRo58TW
6ivsGvBTsFIxXTuNGq1A9w==
`protect END_PROTECTED
