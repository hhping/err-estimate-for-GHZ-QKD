`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfvOeg6VnRuui3qOu8afxgVG6Llg5JJ3Z5tehYdFUfaexdoQdJOBXMMCozcvvsif
jwshD6z9nORzfDZPc1dv39QgiRG29JvGLfs+Wgkaa8NmKYrKwdsTcdEknP4a64D9
0Gna/UFLRx7ExPuzh0hTIGiscAHO/8TNm+OWfu+8kdxMGxRBbYN5GZXqCaXgjNLH
nbXJP31AZC020jhvIBAMVHfrKBvJMUdFi4CQailBvqpxsZI5bZiVwUuleaGTUIOq
ItvC+rsf9Vo3lGw3s1jMM3gMxbY54hDKr3lqQ6qg8g9Q8JAlNUG6BtemTx9ioAmw
8kCKcToW9dzrh4Sg39O2AmV/AGMNcaPr4dcDinj2UCrySRBKoExg+eZB/SQzFSgX
t1S+y/eTz8R/E3djN6YqBb5q8QnaSLD3uk5oIzf3Lt4oGVq4Ep7Duv24H30Sw+Vw
NtcU49KO2dLdhZeiyrzGiXvhmrg13DmSi2jtfwZ1KK5iqYh5fYxlf2Jr+zkKRFsp
zYc6JIcJlLA7C51pDAVE/3riVVy5smJ6IEMqo0HU3VfUhFgT9RoDJsJOZ6vuf7lB
S2KjS9pjuY9jsByO0tOuc6vG18vbh2afgHG+ia6Ywmg0pc6ff7NIlFlkIXv1h0Cg
haVQOSUwCfnlvQJsDmt9icsJB3zwH78610KivbgKJgUj//ngYv1kL9t80zE5NogD
f79VANnhDVjaIhjvBD/xjGESPeAgUJbeVw+SrnZxfRXVSJQI0etjVha1/BKhQnge
f1xaZv6EvmU3i97QcgpADr7MOUD1S/n2WQy+p8dsHafRXPlFdm0PjjWLWwVINbS7
iRmF2i2Zh2FeXe6DG5Kv1UaPIpwRoObFpAebcRQYx+2NhJrzpCOE1Ys9SuKzdAqc
fZ/StvnqZUN9LuQUsmh330DFoPBiyydk69HN9k7Php3DFCSSiVZZPttPKGUs+A9F
PJyNNXGfj6qGWj3PE4Yd6w9hHQZkoAiVuL+GlKrX7wKFe7/WDLoSq8Vt7+q8AdXZ
M1t65Qbq+3Jru0Pn1XOAz8hWkYpgRIuix9La0w32c03DsXwRpOxptoqADrdBmdN3
uDIXy2MrJXxmiYhKttqQsS64jz7kJ84T8W5aQ/IngA66YOYm1i02cTKTyeBmmwhX
I3UTAg0FIpnjjVgD+QBkX6IlAVzgXE02uR5iZ11fsXbnVX93dNrKbgqFHYRUrqPs
C8/CH/NQN/n9V+Equt2TEC3rfRVZ7cD8PfqZ1iSQ3zpM7U3tJ2lhu/2iXTJmMqhr
vv0M+9TGg2H18HtUPINsgjuYyjTUn9ZGPsnGOIhZO8RCW2JfpqYUXZNPSWDTJJpg
tFeokWhjZJ5DQCtLjIEMz8kdQvrZxXXYyEFoRb9R/6bAwZfw5jqRzGtZcHvdcWD2
3biV5iJeJ0dJG0v+DTczBT5P9K91BZ3lW4D+bu4l7P5hZuZpTjYAB3+cX6h/LGA7
dqWwc27bqMovt7IDsBYqiGZevdBLYBfgJDuCR34felmO3qSxdUl+cSp4QN+PO9QU
tP/xQCoEvvhC0AdF/drlXu1Tl4ICon4yD7Vjge61gKZmme4uLktZfWY7savils2g
qqWBrLsz0s825ZOzHwLxMjwJ0A1YA4kQgH1UiRV38S5ldygHFFY8lnXbjtDkSpXU
Vy0bANc8p3oxC/9BGPQErlB7SPrrmsf7FUkJefGYjfN63E7cKk6iiR5zwbWa5BhD
aEUNkMZY2QRWk7Kjooe12TrKLEyTPnyNFMhT4te4GLJ5y/uJFKIkbewliteQYu7q
4n/J1kwhGhThK3WE5sn+0eCod9sT8YlUihsUmeb8g1xlopxAMwTzwKcvfI4Y33F3
NvO544Jm3aeJhIfDFiwx9Or1NRAoAtx4Y81pCGhaB4e6UPqfAI8sD8bktq+lgLhi
FjmT1bd711hyWfOwJ+j/PXijlOnfKn6bztsGjZRc95ZenlIuEQ6ZWJsjMvSHLuVQ
EMSIG22VWCspBjrs72fzSBDjQ27YtWpS2t/afS38lt0ebczfcVE5wYulpKteUZPc
UjhuIMW8QwN+tmrX6+s2BpDxfe/awWbYwZQhKviQI/l72Df4+8oPf9KqJGKbNoyQ
THzh+IOrEuZuwam0JLjA/byPRLJYPsn1YcbxUwf4tGd4dmCa9PseTdxVa52vlO82
+FZ8QNd4E+a9ZEwE8hITOEf7l5F2RbecVyCmRLnzJ6FtHV0u8X+BXytYn7r4lIfJ
TYPZvniOzldfYXs1VG+I40/bm8W/LGp3iNWZtzW4Dj2MR151XiAND269MrAJH6R6
O0AaHIbmSrcB/s/k2e+cLAtbXBZztG7FuO/trTXGtY0vwA0vMzzKJpRz6yeFmT5A
4fG7TBRIVV64LWlq9qYJAXi7tl5oxoh9E2dMB4k62pNl16BhRFSfrS4XLVQKo59s
h0l3PQ4NAZPXRc6saZyzI/3i84sFEsLSLJkwIaVKK4ge9B5iP4PG752hNx3LSMJl
t2A68xfD+O4DthvHZug+Pf1v8PZT6RmFzRMB+xIh+p1nqo+fFQiZRr2ufug+bIEp
vReVRklJNlbEQY7W9Xpv7/UooHEKsrgc4EUWYF58z2VaPFOqBCwWZtzmWb0LfFbU
GJSsyR6DivSG3ra52i/SmAJTsXH51FEu4cAbxCmlY5s59nZK++BFJbJzXJiUQLWV
4+u7mkbh9Ge/o60K1vqrPmed1bcngESb1ZuPeCrT7Pcc5fyP5a1Da27H4Q4tOERZ
Ty3+c0MinXe6bP3I6ZouEaW/d43zOzDE4oLwmnH7QOXuFSnT3QDJLFKn3znyj8oL
mc2FsAouxFBaHst/EQxy9hIRbvzJRiwumsdrGI2X9vz/OK99Nfi5MoRyO5RONz9/
Ftpi7tCkdTJr71b07WTfLd9qOl+YuCEkYINNCoHVjyaZFXKNjV+IA508wbm3d7Ri
Ng8jRO/31qrWrgVMe38si9VnuSpHhaDDK+LGrTdX+BExqoSfRkRmshw191eauzhU
m6xJl9RV5F62RRNDojMUFnmDkeFAqSx5hVjXEDU4It77OiWXfLe0YwuRJFeJT0TI
FLin0ZRqVUYJe0esNCaQnK8A4Lb0VxjL13AaSgANF6aJZ0I+OhiJtrl61KCGyZfO
BUs2Bk3/gxgJP788nSqqf8I5u77k36iDWCufUwlUPvPzw97yZGqfV9lAe4lZ3X6a
cb21imp2ua8NJ0onKEHxe9AfGySCTNMAhrzTAX9fZ1JJu6FrL86uQlxudkTjhC/O
VVQRTupMJftJv83Z17VJibDyCV3P3JKswwDh44+nKdBXkEmCTCysZUj8w2rF/BI9
RTOV+q5B4H9t78zkKQrrW4sW4WQIvu/GzN3+Alwv5jCRe5Y71ztbYcaM9RetHDtY
VPXYVYfHpPCSOBLy9eLPx2XnstaAFTNS2v25t9XmlLBF3Cx5CXPc6TDK21sXKqt0
MBXMLdeUGsJmiZx2opQ99Er27aLD/d0ywBrYZNDBHy4121TQG/j1iJFr5eTq7NS0
9POJ22969yFcOKJ0KW9NtBlqGf5w1NJ/Ah8Exsu96mqasLCRSuVJVpVIj5s9YyCd
aEWfQju4bj6aEViR0g9TkmFkTwKCKg+RNU+664XEzikyQNifusvUG1F2cOVZaKFl
es0HGUHJjUEfuUsqq9f3v72fHw+jzZU6E5FgQ9gnFXxI9BVLNOG5eed7O8qI1ZAg
t7XNNA9oFjN2ZgEcDNfue5dWw2bxpomRTsg4XmUhvBqXCNA6dziCgy5CLKeauCdd
agxXBAxOqK/FgujXTwcfXvAdoLgESibzRm3Cy/q+C0oJHTIQfGdTMnPcX5J0Io8t
zR/SmpMnpgyhPatnAYt6MeG89Ex1Y+1VgC6FSttBHprXtACv7YLLxerFGHWcugzr
0aWvdyR/zUCJ+6yHv4WF0shh7tkLC6oPRS0dNaI0Vby3sj7XKar5IRdhQ81pKJG5
53YyCmNhE6XTz4K4SKqxVQiSQ9ROkDpRs2KTIJsOLYuy67j7WSbY6gjbF9fBN2Fc
Uhmd+vCj5nYqRa37OIpQAleyQaPYKpv1sJ+q7Mg02yUtoz6iHLPqPh0qcCt1+cvY
ZxxXHiRnmtLkJw6RUXKtGO2hujSzhgWypGjjOSlIJJGTVDoFKgOAOC+UZzB5uKHR
+LNhnno4jgHS6Zdw6pjydwBk2iBWXPYyrky1trm6dgcrKgMXdWEVdzW7wohK2dhW
T7CXPFKHd4aXwZfphRD71lWnAYyJYPIYAKBLWWATd8wXtQDqV0IUDonPhrSTpk/N
CzOpnyZfbjWtmIUyLBy78iLjcULfMVBAAESS0uOraikmNt5zq9ROYNXhkmeN+i/i
IhbMuzP6mLJO2WUnGNuPgHPxft+5WTjswyQQd41x+ubGL9MWVH2Cw9ZD60rtu9mv
BRQftepRSBV5Sfu5rzKJXpwPssZ0QV5K01l9AZbhyTZ3yNKIQKLgMFqF2DCB3rQj
SKnfM+BlAjchUE5Ai6KSQNaWhvc/r9otE1HEpb2yTKNALQw/0f0nGUSjUcbq6ZlM
9q+Eozjdxci6c8yGNnkihtdDsDB0n7bVqbd9nC1+WWBXADTgRCeVnqwDxzMlglUW
vHbBEUP9nYFnnrfC8ASwhbZY/n8kvItkThcACMMB9ozKJZWB5dPqb6I6ymoh1Snr
TivNNk2aOl1LKmxi8rE9Cq1odJIEU8FPVHbGFonEvbuVCnfpCrLkYrD4vntxOivS
OasMlo9j/gy/YEUaT8wtON6epdqPeV2IoR8Dx/jkkJXOOtJECGdGcWWLxSzYSzIJ
vuR+5ZegvnzmM9NEpUTB68YDaaHn9B5ezsGStfZ8Ix8dyda5Stb2MG3koFFDt653
kIP9mXIKIghHbwDVZptqBCFQzcvJ32TRdv8Wmk3NgWMavUlKR7mhDhSX1v+VjnVO
OZJTrX6vrYKS1xcY86SRJ9rJ2rZgh4i1WZ6j4KPueOswud2PBUsvU2ae2MW7ksRx
jBJIQl8Fb1do+8nMhV4zRlyWwItEbk3crlIms8CM59InwPJM/DEPvXSvhIt36OpW
smdcvGrl4VjPq1RBINzwBfQpDz6oMyFx9TZ+A5Ey+/UKYc/IWSXMIwpHK9H2Dua5
L0ni1fOfnfTVKB9y6Bo2CBa+52rXI7JGfazfqAvMZAekoxuPCEY2/l3NXAMy24VS
8HjBxLxlGUi3rogrCF53H1eM2t7DD4fzQu2BrUu0NGbwt1UW2uQe+NN2+ne6Jzcz
j727JIz15NN8FCvMe6e0Zw6EQJQ2FlYyTYkEvXIkgEd0pkK/4lsCLYRza3UHoHeF
A1jttBvGceyqg9TBjo62VZ7yhx4bzWm2sZPl9CGcok+jGbAln6ia11OZxUUvn1pV
mIX52KMQ42hqFJncjtcLlFt0WUr4wExIisN19Vvc2+6j2mF+aCKUxxwmmopr6wOZ
kQK17MGp9PUIb+QINRvmh3liK6s3yH/SSCwvrjqonJPOlJLPhGZgjqzy7bLkglJP
ECiVTxTVFUqFgu/rFbjLTIqqqv0XcSyoFbR9H31WTlRMydZoh40+XNubQ1VNxDJF
h8lO73lzXHmWDCpHTmIEb8IMzNeklfBILk9UIn7kVe9tzniL2f+csOil8UO6vqth
Z/Qn2bekv7J7nW2eWrx9dL9iE8WL71gNHgHytVAqTQ0iu/qBTn/MXsvInQQRbSGH
B6UZhz2sU5WeP2p6nLUAWuwilGNNdJqe05MX0k6gC1rVecIhPiHN16E3lDNjaiLY
zvgLs/Ob/mKW5PA9PH5FYK4EAaOLcXRaEdnAC5JHiHt9LIllQ27fBVFu7erf7GpB
2SBAn5tOZi+wMxJupA38Jm+O+9C79iY/tMbPWsQHDAv8f9VU8GB6IMQGbel2qINJ
yd9gzOPyzL7ustMwwJFESdihNFaucE2wmvzV6IvNtiiXCn2VmUzKkT9zQl6Uff2b
XC9juy9u+yS/D9F6kZ4ZAmr9oG62HQTvFu9jlgLP2/BRz01ZD09rRqvFLjacs8Jf
35ry+EgC5YfpY5mxDtd8bAXkluWBgGoNtU8YyNsn+SViyW/jYMN/rBAFXsmYQSI9
6EfA/5Tbg6QZ83IEzgOkwv6Yxf80QygE79YQ3cg1H4gkoc3hD7vFr2ueEPP3Lpt5
5k0rhQOYScX+J8buFlBeGbBsrxViZg7vQxnXGNquavdhuvTHhHaSJzFT8YbmL6rS
Hf1IOo7oBOSDmIQjffW4vGCKMAj3e/GgsPEEasI0YyvgdQDiq+0U/w38e7rypjHd
4VSv90Twws6DC8VbnWtbfCHzUwcfIj5eJEPaiEct4OSzrleesCdKQQSL1bBC0H68
3VcVgH2maIllKfRWBDsi+LBmkNUTb5oZD22Gjk0Z2c5g9Ke7y+TAjcerX2ZhWzLN
JXCJsekCrVUb2a8ZFdYctlEmM59AK+Dj17+nd42H224yOtS6gg/RFkjSd2TSyDfo
tSlzIQC4E4IsZ3Xq5ku++3puHdDPe6Z0+/m/8sq6yRg47TLMsV92G5EiJxCiw2Mx
GVEX52CZI9zAmw1LKtC9w3zkQH4XMRVr6T1Vq2S+Mvl7GyfmMyAnrwGryYEHONwD
smo+Wz9OuxVNvkTL7uIspw75POMYQiKUwl7sGZAokZvIBIfcjNlg+NsPBPJTU9n0
K7LVcO8tjgoQiLQ31XAsXnULHqk7GvRjuLyLdyYvF3sWlVJic8g7gxu5ul7SsFPn
bSAfM0/d5iZq21+ErmZ6foDrBcYr7dAct+Q8ZR4ybxj1122cM+8WZslWJ2oczCi7
ca/ST9hPZb5NZstH+X/SYwkZHZfZjaOaExkEnkUoHmt6zID8/3/yqWMJhVfH+RCQ
jZhBAMfoE+Rtzv8A3VCmCVDl99nqDmNeWBtXHbR5u5SsMKotgaxfsp8qqqFT+42T
cq1fI89BxDWkb2TeSF1C7558jDWR444HBgrSZHoXP9Ik3WsyH+eOqNnaRRZUNKAI
8VeLEYg+bjtRNpa+MkZcHV9dXxqXFSlj/eDbljNPEiL1cotoO8p5NTZ3kYRwDD7X
JJCrvL9Zbhq4lpQjrx2M5S3qFHzJ2K5M5iBhf2jH7WWmJJqG5DzYpKh0E/SuAlYA
wtCMp6owhO7pQjU4cXWAS0t2h6fFpSn7va5Hphqp+7ZetUDxGldTrnKWJ8QWunHY
7O2xKsHOS+PuoiCsQieDg/iBDHGR3I1Xe9oiS9Pjbg4e01OFEjGhw0f09IerZHm+
sWZPo3UznWDjzMxTqE5xLIIx6WqF7hKJVpzoeLS6M0szXVoXNALQunE7l5WCKDzW
MT1ExN+ObDLdrXH8gmTrmvB4FpcZcb+XFD7UA8U7sI2SBmPwkU8CjfZ+5J+XlYCj
Jjq3Q1i8DfFZJEHTB6yhoAzZ6wzfJ1IZC13pN8gYp8JlfyjqiSfWoRQwCtgv1LUG
mt+lSjOhGNdhSliME9CkywrwKWnM2JMm+SVzrYqL3cegybIAlAzbz/fxqxNs3Z+w
vDiJtE0mT+Sw6fCmEGYFnZxUU725BsO99aHP9WDwku78fN3CBraewmxR2WxXkOCj
olMBXY7tukcX7/+jw3RgQGdot0t0jwrZZvZ3TQfRyNoxaXgUFeKgzISoSALPKs1H
81CZiFOCMM+7ncZgaXtDWxZj0lOgQzJ9u28wWJazds3MJLff9b+xiS7wtyp9cBWr
jAjEyup2BGtAa0qVFKoXwLnA/WD/F97CHNgnVT6/Ch1P1Ajv3jtyDrdOgfMalyQc
Qd4dON4R1Azze6Lt5I9FqdAgE5TPjS2pw40ba8FQnOaO05toPm7I8G9w809k/Xyt
IVNxff4nZitKSsd4mz402K9FK9kNeVI1Pxx6KEGIHvgo6XvKyPJl8BwtAHaNWp2V
FCi5+0+p6561+hAvZTWtnSx+RT+1CYg/02cqKQl5erhmk49di6CeNOl5eZC6jsWW
jPgsgPBevk4A4uIidUijXtT+rf0ACPzxS2Wa1dBDlfuu3x+ooQJK6e5aWqdMUava
xn62lpasmlPY2xhjkNW51R3YImxK7F2wpgG3X2nwf7Mw4/4A/t7muOXmFxW5m13G
Uqzddw+cjIXzaHVM0fqicNGDWRirtqKTnE+LIU1RGRsQTTQENlms+RYGoLy4nYo7
0AT/XIbrUQ9WKgJfqhOQIH3BoMpdW+Y2EtuB14qrNvr90XOGzMrXnBeFECypENs1
FHG1vVThLhO4Q6Uv6FcmhKIjZdyzJbkF2qvPdrRGW/E4kQ8m7skYR275RKOjOELW
NbLuZko/CLMRICQYZfKVAUbshcA+3GwMtiTc9G88+hsA7v1vhHCfnp40VoachfeA
hEuwjuY1anE94t9ygieeqaobWjtQsg2G3CUEzlKPI5T/JRsl8C30bGUSymPwlZaW
E8gebXYbaLzv5WBt8AGl8WtwGQj5uipdwpqDRXmZfozM5edANSgDdkOwwK7zP2a6
3s42H11vUzISwTSERvRymKR913zPFrN2SQ0evEN3GQLULQ64YRV+eaPMVDbRKJG5
z/ZLUb/XAUDcgZywKNMbA7gu3dl5sX7Sn3EEqHgRPd0j3/SQTuFBHleojDIEgncj
u3FaN7soTRLCWqVsHi6w2oaLWV7pIrwtzovYlpOXlrWGk3eMnnxN7SzUHa5Eqcm/
HN/KzltRTubQhW4t2gPE6wa3sfsw7Osvk/zbPHbwA6O2gp1oyney7Ncisx9uK5LC
U7BcausPMcCgw/ILe0aKnOoIgFRKGluPU3jIJR6hZfZ7/E+N+znccZQefWGR3Fkf
VoQ+oDRmcwI+y9aEMDOJ6gJGSYpQM4JX1O5ULvQ84XlD7gfFXwcBV8mcxxDKdhsZ
iUUj3Pers2xb2b1dRYMONX6t30mDoVpZJwmCKakcZZhuo07Al0C776oiv5KBsde0
YwLcRoM8sIrjNtpCu73dEUNfuxItOmpmf7B4hKhnphIruypf+tXyz/3iYKumkqgs
5oPYzPqCfBjcqEI5jPOoJxs1NbPOrygJCriTFSEB7hRaYUyeyCIlsFc4HfW24FZK
l6TcePgdh3d5WYEWxFPJNKTDcN88v8oUHJ+f3pfm5OQ=
`protect END_PROTECTED
