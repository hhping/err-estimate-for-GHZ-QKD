`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7U6zP04vWSfEGyD+eLNiMS6LSLMPs4ifPmZz+4KtQeIS2N/mFwXt+N13HZFrkKm
g9KcLXt5fy8UurmrcO9SJRbc/YF5TTfRWGDbT2kTTuPl6820Kdxce3LQ8fxq+42M
1QujY0VJKK258d97Cum4tgUqGyUEj/ak5SUu7LbCdRjIBCuN9C6tSti+wfpUljR/
+S66I4UaZx8mBFKdCKKJUK/biLtz1IbPfCa6bvug/xiFIhAohiOeNlmsXaSuUJZ6
SGXDxGxIRRcKrstVdnEqcM2pTHANJ+oy4oWoNGtcba+Ms0PyjkYigsg4x7ny2/Xd
ykKZIlX/5gki/OOcgRGhVv/nhh4sJR33EwLX1TYdaZyVA/WqTxgqHcArx5pARRXj
j/RcVYp9mu6eD2Rraf0S8ukIxFmv9THK0DA/40xfgmXZ6G9Oh/FtxEzVamjOROjq
09bNlT6i+NU8NEtiON7k9hPTXV1yLmjcgRp3Iaix5lmqvSPcIA2UHEFeXXlPZsrL
i9MtZUZRYGE7GaFeekiOwqDEbXQKvP1ra5SifeaQGU+ZdeUvJGhUp0e3o7ny8Baa
18HABQMloOZ/N5bWvGpm3H6oyjLTODjsFT00Q3GR8vOCdlzGMSi8eFzVtwB54xbb
MeHlrGpS4HOO4VygCHZeAUpQEHYxDtI7wosTEJwZoGcViehyVHpNC5dkeqCdIDlf
U7bqgSBZcraJzG7qa7pMeGlqounZ9QDKzFDGn6qgnGvZbfSoVsDnmCgVktFp92lg
UMZ0wytfGwWf0dKOQfKbxG5sdbmBTbs1CXyDw4vGi+r67dKTav5Kj0I3jI40m21+
`protect END_PROTECTED
