`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j10685wL8zKQ3Ej4JTR7aT2Sr28S5IVzS7p4JRzWA/z3rgplirk/1q9v9985NJS/
G7Gl4ZEJy5XNTDbbKXGu31/obI1W6kVZPSnQzxOg7sxl5xWFlGhMiXIhzWg9X3bf
Y7zhXOiUgjQALoTmUzqgImTET5e86+MQIYQppEDx4jmRv2tQkKg4GssGsU4gwEyM
evLEEa9Q1mlubhNwqXMMuCHGBaqrbKDadLQxHqBII1JEPwhkTGXWtsAs79N70Gcu
ikqOG2Nhu7FXgETX2Q9/AirWSqsyvkIexOKEOYq/gHjjf/juO/5R1x/wKfQkckwr
lcTa6rOUSnJ2NGXn7i2ZMjUuntsjUrOkYEYR8PVR/ZbyWD6LYm0p/WNdfulRhXul
Ge/txApLxJ4CSIpTKuj7thzbZJVvFBb8oxWRTgCdJ8EZR9H/qcBxHBFRE6Mw3s8C
4xPESqnoGBlHZPjOfbltTYuRThGfptTEsKYDXIrZEvXVD0FHsmCSq32Oe3B5lzpi
peNzZbcT4Mcp9LnHhWxb6B4cISnvzbP3Raaw1z4tXLQHjo5vMtvU41NKHV6Qw6qS
+1WIJ1/YuBdhYx5OBxL55dqfMh49jRiVbvCL+A6xPgE1bgCWihtu4uKDosi8FltT
AAtUBoDlBx828ELuSJ/lG3KeLPuhKqJYtqELwGAXgyDHvSC+7RPb6CJCWiPnzaC5
kVVkHqWtu18F5JUhga6GCHa8Qls2NGTZ0geLViRRPMKaBvxjZ1ISnhfjpcjdO6GV
/HuPCMWnrhBOCBHhfdhd9eaJaconKjZjnAU2ghGIMblr8wzHBQRKK3ilwoyPjC1o
pxuq/aFdWjHkrCZfWdL2QCmldAemBNOugGHOfvWrlgaZbGAtG4VRKwx7f+29X7KZ
I5n/+dacACCVtF5Jn68rgyq1V2DMXsmHYuzvZS/Q35p1piw7HAkmbGbP7kPxW3Qa
5x3IDmiFIJqIIZebqR5kChVwxwQGA2QkFW/y+NUWo7N9e8oqy0Ky9lf2i48Gy2Vd
hWEcr5PgQDaxetgOLkmKN18DdEDdSQxdC+QeUyEV+MM62cKZRqwGIMFgc+rEwQ03
me+SLaxQl0NMjhHKwKQs4Rvsg7SJ/ipMINBDxJVt50PY1ceghiADi2vbGMUlsoIB
`protect END_PROTECTED
