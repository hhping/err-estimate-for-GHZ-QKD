`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohxj1/u2Xg5TFmPksjQFlJKarhUA5PGhyO/kunuSAXuvPBqKtqIAkAU1W2zCcWfQ
Xa17W8nmFg12Rz9W6IGleDNIgttUrVRZejk9Ef7BOCDr3erxnprc715VlwG3U1/5
dCJxLfXpP4ThHsgBgHjCelnTiUuHD3HbQhTHsq53OZV8KEjZgLMf5svF1sC1S9DS
bUbQkhSXZ5Kkbq+KKV3O0uKf6gNXEvBHNv3kyBzoS50N7m54zomj+C69N58i4ThG
WYx35aQe14BshIyKsChXUOsZC7QMOYmixgaNrc14HzbpqjHkm7RpR0UHz/bUSVks
bQCuKVp5YG5NcBuyG4rjKJFNqWjGxMo3H1VjBhcoJfpjwrLbkXBjW6ZMvizBXG2f
t0o8Zu3OxAyrD67ID6deZd9zb77hJaLECwTm5+TaG9JuO+LbT/WxwX69g5XD4PvR
qaA8st0UMgaEvbzVynjpfZVfS3BZCy4uT4kRynY9y1K2wnSmGhGvEuNIgR9R+1b5
bFnCabWajG5l0TLQNt6ySIo4lzWpRAZOjwERb4vm+0td66oY2EhC92EqXEPgV83G
Rvs4jxEgwiQlZAeXbQSpbGJXgnVEv1ArmScxqXYrXU0ebbYheElhbOJDySVsG0Kt
rgFDdBSm7EVSPUDMYAN2Q7CbRqHuGadRZYUKngonfsSzcaSecfYMxbDGJX6wH0wY
xVirNyMolmDG42YnbgjfJ9ElQHzbzhnYx/HYNitfQ9ZcaZTLMY7py2iZKiTd8hIn
0TIIuf9r/f/x9DO5wngaWNVfoAAThBQRjASyCF0tPSe5pBgxY4kkAzZHNZ/m9d1D
M9nVj1Z8UFpwoTRkQDrzjmEoj7J/D01VJgKkn+THYQU5Sy2i22NG0yoZOhtsloS0
+38sUvuOfme0uAg9pJ7JsSBSkZDMtTyOZdnmCdLtkn0xVv3Smfy67IH9j47k43EC
XGndyJR54rPlvGNJiqNCBvzcEO6RmXJs64WeZnL4EI1RN67o6OD5K14aEjViH+LY
/Maa1vB7WtiWp04mBL9+NXwT3HjPOUOxSTeA0kAYqHQ96GdksrqHm3TAx/UpNzj6
HSOjTjv8A1GZ83vni4CRZDuF2PKSzaKTxmFJjwF8O36wM30Xl7CRKh6f6Oh9NPAz
acL5DpnsUFnFxWIQUf1ZarzsWklTDp8IPrM9jSAC+mjlJe1XjMDXN/HOxi8Zq+Vq
NpWLbrVKaDaVycnzGUUWvVwNmoN5sJOg0SAKINKOtVZU49Bti6Aj0RNv4UXmeLsW
v9HUabZ/R2FOjbNgEg/CWXkBkD/0T9bYc9h1eemrdzkQJwtSg7HAwyygLtuY46Jw
PvrXnPOZ2p8jxa48zitHZ+3z/ngHuTPdfEz3tKj7ft0BuAe8xEHZt2Ip2q7JHMW3
axiR0Emhpa65mGyXcvc14dS8DC4o9zCLHogPwCJiDC/MsYIXjH1ewOtOalZcIeKr
nwXjwSSJCmOFuaSg4OO+Nyj49EradxUW1r10GNT+q4PWhrbaYKY5sv1VK7it+tKX
Oc1vXli+deQNmKN/81tCoeDtE0f7eWj/lecpC9SspqnNmW/sdvrh4p1qSPAn/AMx
RyB5ZeBDPmL26K3v4xxqc7gLbrKicR/MDIL9gZHmHqitplbl2K9BiD7+XpKh/+58
+r2WZTl9nrhRHo9tzNPCgZDQGz87VOKAk/vmWmWKc7qvUtbapV2NqWZt53HiBFEm
FSb5cp5Dvg3X1zMdYjxiyClkvzjHrxOa1GxRpHv88YD+EfaxB+jiDcDCzs2TGdhr
V8u4KwNYm5p/vY44FfMFCzbvsBYujrW4POXMViHl8Vb1gCP8+WL0RTP5FOUt8JY2
yvLQZcT7V1lAaatntIJvDTitYzPyokjHS+rD8BbDHB3l7H4eRW3dwh2erT2cCADK
HHvdZa9DB/w5YBCrH3/lSHET1Km0P3uu3dDpUJ6ztOC2yRmf5d9D5TeCIv6GV79C
zLdEY3hQ/cHSVcl0EyiKDKBakkFlOTMfWIWbqTJxfclhyXRlgQuvLg4Afx5Zfx30
Uky0oXJ7SpYDUkbtWcFcq5kG1zxbet4BSRsFPKjd+Dv9xABfMHaJJE7xnHh6na9g
XBNaVx2nGu9m5tb5Wu1mMjHE8uNKrjSS9qH6jcYjzjYFpEs+ip9TxVlOTfmdEmRN
DTXMrnXbDDofJFrpYjo57CtoXY11cT2s40uuvKVm3ypxViCf5S830xNRvwZNKVBS
Y6ZLUmNT4N60hujJYdAn9QgOKcqbq9VF3b6GqwhTkS6i+erWSGi+0fC0N/6lx/Qy
UsW2s7pZesIc+6ZBQECR2U7A4dM5XutiUndYtT7diyi8dldNh6xijhWWifRAdCVE
uXu/MBNdcCN21Ab0s4HA0wzOUPAhsTRxB92si3Tmik09SOj39xKHY97aViatI84K
MW3WM2eeILAFVasdFfqDVtxrEuyDrkvokFR3WM0WYpkFqBJqM7+7riz8xUHqUBRV
NijjqJ7X4suC5GpYrR3GpFemz42o5ZsdKKe2drGnDJBUCttfV4dIhl9yhuuWjBOW
kZ5BN9GAKn4JvDzF279S0pEZ3CmDMur8O9t93+tegB9dxAY5JgbtKKgCdgL1ZoTX
ZRK1xTRa1/XCaOLW4n/Orw==
`protect END_PROTECTED
