`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBXwXIg5Rc+I8EoLBBgVqbJnqLje+gMu17IzSTU9ZfFUHNrkOsK8PyCISXuXluO9
NqrIWEnfWVW82336aCsrbmE4xrWCrhhJGS45AJnx7i/g69Jx0YhAIb6fDQCMldqb
1aWHoHCaZXT++TKlr2yq+RvfiPgyg4hvqCoSOCGaZzU23FjVa8O/Ioe+Jj3wUs+r
cBu3t0o6pPEhvIT8Tz2u/mWjCT+gzXLLp2Zpj1HS9T3QPsI0gG83Q31itVReJoap
57oGYzQvRSGhn9l6Vd466Lm+9f3ywisIaMgeEWnSKg/MnhPUh9j2HP2CRztmR4ON
UdhDjhwwYYFW+86yL00Nala09mi/5tnZ536Hlw6X3Xg4sSbC8sDtUtai3oQhVR7i
XYuILq7X2zlbsQy/T96H6H8do57LXR2DNcb8Puk+czAeV2ywZfsdDW476zsq9dU7
v5ia5W74LDRYKufsiRq55NRtSZ7RpTDz4/KvAoWmpTl4E+ZAt3Hk7O9WsJumhLbD
9hGhF5ZSVzOVtilB+/I01zb4guX0CzflQ8sIL7XCIzL01GdSRGvAgCfMyFROZatZ
TcZUiQ2bLVDabRPBL1YJjNp0ZNYgamX5o/1hxEsjd15UYN3g4/eVn9crRljRm1Em
FmdYjCe2ZLgQg5pp83gO9w==
`protect END_PROTECTED
