`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T7bND2emQAKKcoh+HN+88gJYS+V9BE8hyW8NXp32qr7o0CPvGiJahbC7S92udl83
FXKSS8WCAiedVVPb0vRDkLSXWlLodEibnDZ+TLEa2dORWt3TK52zFkt9P2krTgnw
rIZS9P55UEiBmIe01hsclYSyFZYGC7GDRFbF3BaCr1/vfKnGBisJnZVW1JUO7HAP
8BwkcDd3+50hAETaml06X3iv+cBu+BTgTFtXJWdWzDPVvi23l362mF/ds1gpvA02
vDNfXhnpsT4K3/+jGib3TtwglPexF4nL/NmSZTbuOqB8Mo1k/CzKXJFPU5BnopD6
2zlIcfcM70/AAQzmldFxNG5zOMSWPeRkaS89L2pjJU0U8eeIN3SOCiFO9CNSGFA2
6ydwGCvjchH5dMgLtCcLw92dJ0VQEOdAN0DAruIsjo0y4y/Bx25de+R2Cj/FCvaV
xI0Bg+UFfdVqkFpIgyZ8WAYQ9HoXNejOnuKK4EHWDvGCzEXxh4nAt8rdw5xfID0N
z1h9OyQm1ZxmlHEyrJFso1+iSUYXjo/c+JvMK05h6gsdRIHHYF/riqTYMTY4vLte
oyL4NlGT0HLzvSAXXysvEApc12D51ztoUi/9/A3AyPC4O+D6NmijJYWr9z+HIGe4
X4VhEeDUFtGefR/i0lebRBR0/XhOndjmGUltoQ7bOjGg1Cbh098ovd9S8RyMP8fx
1jyz1t8WEe8AuzajyymEGSttEGmen+H59IlMfg+jJizfWcDDh6Fh9NNq/xo0xG2E
BzTsNbHKmUic/BIChHmPiB8S8AyoH6k21vM+0J+VdZ84G1R19aBdVwh55o17ZZVD
`protect END_PROTECTED
