`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PW8XZk43SchnaPLMInBTmiQjPQrWgOF+IvwkZtdNGEGyo9TApS6kvzek9aYI/G7
sAA2bgRq/dK5aj/XkpHuxXIwHuZa1G6lawAQ+3VpxH7EQ2jy08eFyRtyB/mx1WLI
OCZkExtrANL/GauPqD5TvrxiOM0NwuPch+AzUG5HaDz5/XJ+XTcsxxCXIgU3tF23
izvjU8h5jbEl9qYV5VBX+Y/L3qS3mxThD7sbaTbw4G9xOkThTgLZmCHFQMfzRR/m
Piui6gdlk0LLX8CVXH2T6sIKVHsRzRg5Db81du8mEJmg8924wkh/NyMVZ6PypeUI
OWb8pFG6InXLlOixBeB4uAfcYA3rxXISFR9gcBOJiUAHr/TiHiJ4gTafJW37LB4+
8dOh/4LvKhpvTGiso4B0A26ojXgm03wXQVC5muG8qj+yTrYoVXKogk+va64aYbfs
iTCY0zar+WiL01kVMNa/x9ma5UltEfsc7k8ECXBka71KbZ2vo8vsdnrebxfjbvZa
kOcw6thyNvtI8BtveRgcuafvg4cdTQuJwMrOaaSz6LgZi8iFDTYrnzE/ITX5V2LA
hqtLAesDEOMfMAvNDdhe7UYKgeVeIDt/uO+RD/ErZjCdwfA7ORWogMcKZDLbeXzV
2RYLtVg/iGp5hG04ORBJKsy3GCh227Vfs3e4p3CBz66gldd0owMSmQMZN1y33y4t
I3k185KdZde29AXlWogQ+W1P9O0aQUOdVFYgiOLuqhci3DjQ1IF45L81Pi/1xrXf
4RjEoArYYjw1IUWB+DpneA3pG4FZ3UbOF6wr28pOmvnY5EZMlHMRCy2iTDt72Jpt
08i1peACkC8ind6aRnbkfCeaiXBceAy0lPooR/z6uyh/2o3rJxjeff7tR2PAoyhd
dCSn+AXxzm7Ih/kJgKtbS6HHcY5mxhmvMLKOBub586QWVIGBl5pRIWNGWziZRVWO
WqrV8qJy00/YoTBuwtp8YnbtkTjpGOycFCwiKJ7ZAHMW8Bp2Zpixw29Z/k3nZI53
kW2vwR9cteuhvwcVmJG1wjIJL7msePv6fgP/j3aNGkkMh3b+A9rwLBizJU/Yc/a8
XdFGdSHFHV2ggwRpg/iMYg==
`protect END_PROTECTED
