`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84rgAeUhx9zcLrOai0styXJHAKDrhUtS5sEevG9txAZq29b35/8k4pKWCsj8q7sO
fmXOA0U6rVbWHMLIYkUzjQFdp+0PA31aAbPhRPcETU4MzjSHmwo+XizYmL3FPgzp
fN3XewyLpuTaCJTopr/m003F0mC3xtzcln+rAaewGkmFUiPSSUaaBGr6cqh6IQAT
Bkvr/tFHnZKhxFGTIz8zKbEZVeDDBG44okMNd6AZQo0c+qB2aUPi4NhplcP/CCNL
hTx6g4eKRoRlt6QxX9b+v7lX5bMyHvraZpG1BAF4G+7K00/MFuBU2rYDrQfOtZ+N
N5rwWLLNT79l5lH+81hJh2QxjY1EJwEcdV8DePP6oumXEZtCJRnDJeVC+StMoZ1x
i1hISAq/9Fn7yP0ORrluMkETwB76GbLVznV1ibDCmB3cplCa1JIuXWE9sCdqMx2D
DHbWbjYgQD4JP4kUigfjR9UsXJ0Nr5bEqWiClXGMDrouF2sNNQix4p/Mo2GY2bhm
NCBjii5iX4J24HovXk3wCnzhD8FDyI4u2RdIlUD7tgWgNs5P7YQGb7xQA/34wKpx
dbNON80RId6P8RTnNJaUkNFpX6DZC/9TBvHKU9pkGN79FOiMOxHH0avEld6ooFug
r3lLyF/VXfRSRAVkl7R0RblSRrm58LmkVWsSa52K4ftOGs5QdimhY1NO8Z1n3i2t
5DP89SqFsswTnvvCDAWIg4n8gYXggioJAT49nRo7X1OLlzZ+nE/IZpLICYIoe5tI
f1FtXbHSY7a05yErIorvMNRREhqtcUskqjr5O4vxNMfAHAtTmpMZ18Hudj5Ztbct
+XtBuEZYmkWcAY2mExGUngXzxNRvLP0QqIJA/SnZ4TbLsIrkYg7VpN8qzN6LNu1F
FFLkCXGAol92s6fTyfK1jXgSjhka1iDsG7DliDOXWEmg/+yGJPZjnArcBQRSMSEW
ArNPvK6yxcifGDkXbMFTLitDXT1E8+pthbEuW1TeiMbNNTDatOslUacSMgFW79gv
QDQktimtd74E9JxPkYxFythIVcTiTWMDDbpCeNKHgOYz4SQa52Nn5GneIeyIqDTe
Tx3JuLcWBTmO+h2/WweL5NQb9dOs4JK3ywWMoyxFoYWoflkQ7hTzcBDL5jHdCFc0
cc/p7643Ghcm48B7ELS75c7W0OEuKs4w/TmNJ6njcylDvrZTgcbw3hN5Jzs6YSYt
pLxHrBJJiGuBWd/Xa5mBZ3U+nVru4Cn0tlo69uKi82lBloh0y3fJyG7rIXdj2dIg
rIyDTYzVZD6CV8XWAVMc8M2/NzVmB9XgQcnVvpML9sLuz7YbRx74OA19L0E2cmYF
HrF45c+a9bUnhGrbd4b1gviPSoW7Q6e9u3XiINAYJ6nI5/714mfe7M/5PiWsb2e2
OH9kL3pX1xR+Dryj486fQ2n3hsJH4CSg4HKMHigUKC0WZ/9dyQDPH5dImzN02Rxc
Zhe3k/2qCr3wx+zw3rmWVT920hMCQr+HnKRSKm3gHpcnywlMp9MwgGCJ+7lhZVH5
YwaZo4SldIWI7l20xZNiBIQIlnSKP1dnnOEy1tGBNauCMMVopCNhJB5mKXXNsjKr
lF2Sdl1LQs4L/kgD5URoyrh1XN5zLG7VCaxIwR/6wPdZlorCu1tL6OSqd4Ab9eso
JGqBz/T+T3OCjlF9Zf/6By297GCB2bEXoyA0VBi2CSCJdCCSrquf4cuGC1144/RN
k8uwaLoG71ZWW11WNWuQqvAMJeSWMjsoxQLt+sLDg5LIpQ+Taerv44kzcSHEfwKB
x8RcAzAStTErYlOysaj+0A7Fb4sar4P5N8fkfP1lFigHcPMSpeGlSAEchNnzlu1+
Qb7W/6lG4H1S3JzRf2EEEtC8STwDjsEQYOp0+uqG+e3HfuB9p5cntaJFdbQklxqW
PcrPqyDtuL0UkfoDc844+suZw8jgXGw35B0MEQUccKHAJsKRKKuUXdxVIlfMn5eh
ijx5/AvfmJr2EyvEr3CZVpEvDkIiav8e16fFotw4+WFiIa29LM/+XjYps1rBKe5X
oo0ahB0SXfKD7xpRFIoo1y8P5qBmBgJQl8t5pJ0y7GlICYoWaAeBCPlxtgDR/FpI
QK2TIrWDjGrWQ0yuqHh7ny8SRMPxM8n9aj3rjUWPx3SFixVk9HBPSw+JUZj+he5S
1XPWv/LLJdsGKv2ihnlDXGP0IMWxusvyONd+vxs4KLSQg9T3vHXR3Y/mrpOnTawn
R8VSPKXIobbuvWxmpXcMdxjBNygsGd3tcUvG5MBRAjT3mOBqzbItlkIBUGl24XVY
Iinx4ZaiXBmLSmrAkLrFPA0eTWOfCf0QsEQi/mKlLxOsjsp5f3t2WJshVvhe40p1
n+W2vk8HQiLBDXwm5ocJnu9WU6yQRoEbG/QKAouIiSWgXRefP/GSIHpeLXqLBY81
jYT3JA98H9EHVbghQhHcIS8fpTC4VdiNUyvn3Tqx8WfZ/10b9YqFFNKyAKMXpnxC
qTiHOig4mOi4puziYlEEsZoF1vaazJ7G5lbxjqatElhd39QfcxHuId6YaUoh5O7G
ghf72bo/wyrKhNNm68H1nKD0fp6bzEE4dxb0Ln6PxzP+yzleE8uwyUd0Q67p1l6W
Rz6kQLl7lsYXlKbyJeNr4vBTzCuyW0BMwdHIokl4tgpYdfHVmmyUAfCXgybycpr2
TW/0HAmacmsaxQnOPs49MqyV+dY8e2iL7fQn/0zP7yFRzZKNqVplfTfoFHF28SJk
1aEbkCZtR2hkJee1We7n5t+2KZccZiZgHim1MrZlH3hDkfA0MMAl6mjB1zRO2+AB
Q2zWDdCt63MFFe260Mg/8dZNwQ37KeuqfOwtf3Wd1PvhHF+2i+EK84trUE6Au+Y3
u4c9P06ZLGw9lpbKNuUJlcu1OzD67b0O/W00CoTtkzXbHnAPIb5BkziVfkts9hI0
8Wg2T+F81nnUvERY/ObAUgNRhbCWfT3jHdpVikKt4+Uko2KaoduKdzwvcOvWAuSQ
3Y9hcCEe6a/LSoWahQakw5PT0JC4Q+ND0xUuYR0BZ62XMAYT2BU24YD/ZcWP+lT7
/jvOJlruSYh3Q4F6bpc09eGABqyaDO0qLHNb0n44v3nYpXxjawgPH8Sa28SAbuPM
kedkM/Qx5LLi7v0BU/oNORQYB3Tfe5qyfVP1PB8TrHKNo70rJYD1RolUT5Nz3aF1
qbljPo6I72A4ckvBaU1f4aOk/eqNCrQF7FOEQUHTnz4Xzbxbd2iznWIWPUFcX/Xc
NnsLa97wFP7y30y2Y6mycDaF50u2GQntSeonNC65IE1nw7C+n0qv9NqodRGYF4Nu
IjcDVeqBdwbVxRWAM+3ehAMME05iF9eXl6n9+sW0u2Ujbcmbjnh4HN9cwgN7Veaf
ka4qpd/fyFc+FqgRbAUjp0sL+C61YaqtJ8Tyv2rn+MhNGkhW1Mj6vSHRBcpzqjRJ
Kv9BNYvPmfw2pAeDz4IiOJfWP5oKeqF1kFMyAuirZeXgnKdjMne3OrU/On/nXYe8
CKZFH5BpKdoMHEEWWnPHvS5nB/99qaFLObKa2BSZ30a+pomv4CGFybvVT3IgO3DX
WwxmTBCxommnbTW3Pj+kG3r6WRK2p6gJdwoY9PADrX2iV6Xa8ZxwPxTbcMoee5rw
Qftl7XNFAO41ywlSTeArFoLxpR16DgQzySFIHLyEJo7WzPCO3j4vvwoGiHDiB2ha
B/Sr3kvxOeJhLeHmq1gPv+p8l47DGXfhCRp8kg1fQZZ20jOJ14RYfHo/B/FVVB8w
tsckPp6OLclKl73tYutH7Ae2nEbss+dvaDqEDIXZjzVVWfG6pe2OIU5WWbMI58cI
xSPRioeqbNJQpGBnQQi5BrWCaOyyJA2tgPuHR7BpSVLYHjJGoNPFDPhVpqg8JD2i
QZSm7s6kryTkRdq9oeo08AeGZW0boLmFMoPBmQDi8qjqUdHB9dCMEUEFIAmeajcj
C9XmdAiUN4JvNKe9O4Jy9OSt/uwrHTHHlrC8GyGoVBjRW81dRC9pGaxld2a/21ht
fJFGrl5th6MJWVWKrFlLK9aHTevrLvDUCP3damRmaTE3gOyC7z0B8bYkeq6xuGwR
`protect END_PROTECTED
