`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PI3tZTZIQwVoOCDv3My9iqnKKCuiHXm1aoY3Z/12kuRziSIZ3kY9AmIgJeN+Q+O5
+zpwPqBrqlaBsOQ6R3jAKSfhl6ctpMXA26BMGqYs9BZi7sz5rbz1cyevLj+ShCLL
JXnfH+mqlJB6ZnDE/g+c/kvhHI1BJCKtF1U3mD58nFaT9Fa5vwR/7LipN9SQuRRo
BPLvJyBLqRQMlqCfqpSvtw8gLYpXuj2vXA69MYuXOo1RlBRVYlykFTAqI3S7tEj3
mrpJm/h+RNdynvNL97mCupWsUvlGGPWCaW/RRBbPg7fGZBvvuRRQU0CKxxHavWIv
MMG7IhI5dnxxDz2LSYXgFxaPyCGmMWxGH9/qyGASBlC6IaefoiPa1Wv71e56Zo+M
BNdPzgSAGEivMp6AbzRyI9OfpKohuIjOnCgxNc6MOV0HjO0PbzonOdhq2nYEgYr5
QZVIDzv6binr0/kmS3n5heHDkerzLmjPsnnVFqcygPUxPWPFWAJ8aAjJuLB5DgL8
mY+ykQoi4zN71aIQJEP0jbRCd9Nsyh4o57jqBH+Pd/JrGjeN2DdaaLgdWq45VUOi
znsTl9b6kmUWQgwxOJ3a4A==
`protect END_PROTECTED
