`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JO/py4Kq6IKLsjWD1DYma5F0vHpLNN67uVU1Sa0O6SguLvKYrxu4MgQ0COKmG51v
SG4UDXsnF1n/ADGnUfUZgwtC/YxXgctl+KblLm1yzWxCrsbZZBdax/78wCSMca+r
zJMyQrnTC79ZksPy/6qQmOtx0MjYSLKpi7/7d+8qRZuyQWbCb+eHBevxBtW6KKw/
Jl0Ns9BzMzIRze6//CFnWTfgSn07h1EBEtzKE0CBw2y83YAhsWBjN59BrKJhNtby
oa4SqVDdhEBmmtrXq/3GdLb1yzCuhQhIEi/bXw2AG/s/8zq7tvQEQWApvC1U/EHU
OFa+UWTuP8vaPj7exLIs3VyI027pEls3oBIYr0XZ074uvHUCT6wFV4tfQk8zQZj5
SGNxvxQGc594VDwet4cPxvxCatPxYhq42WGBkMj7ur59ICEsSXlrjwQOxPTco6Om
1HIXyXd090InAyecOarCEwHt6RQ8cyO5ynFKOa4/adHoeohL/oY7T7LjfBms34hL
VpiUrIV+RKITg6Bn73SOy3OT36GU58hqVDXp8eUd0v2uHc98lABFPdFoekHjHBUh
aGbrXOD/jsBF1IM/LEv5lXNRbNwO7HTHgcENRdgTNa0NspJf83itvwgD76rzAmqy
alftDFfEMYRpubyc4uZ4s0p6AzE1GY8uml9SFfTs1+Znl2GvUXiA4ipHN5nl2Jv0
eRIwnUwG2rYxx7srxyOxYzrdiKQGEGlnbdM+ash9hIOO7YyGfgmtDHVcNPaOcYuF
sAdXGTkyZWrSE8G721kAQfOcE+CdGe7s61tXsfYR+MnxVXRO4uuuUPyJQDZAI3xp
/D1DonelM8WHhcx2Ys6BDJ+CynkNcbZuWDJ6CwJ04gZNN2AXIkns5W+CFoMbZ4IL
yMNiL+h4F09kYwS/j/q/hfmOdMJGryI2n0fcSCjti9C6NhFekmwUJWsOLnt1fymu
mg8HlUPQtzz8vVNHfzrrEkpQ+bTryIE9iNuNzCRdHIEe4n0wpFikHMM7g/am2LmE
OR6Hd4+COxWfVdAjcjtAEV7suQVl4e6GonLB5DPRFxTMu86/RkSdvTif2VKohv8r
1stA25bCbpEQlTimrbAhqVasT4Xyy7vLoU45jmXFEATZ1oy9xsv/wdZNFq4a7HMG
/J1NUkJmvxo/6NofA4SLc98ukH1Wm6RALYoRFxgp1wbZccnQDXYTBp+moF2kTAYr
7b/hbol7oP4oHOz+rTx/RO7h71/TKMUPu/GcR5QrNf18exYISnXoivKnztV+1kea
BuqvF091abHn8lThKwo4HaF1qeKrII2uUuaVR5mcf2pF4lgKhpNF4eHiQHEwVdpX
suuA8M6XFl1GlSMHPV9C9rgNqE+BFYR2LkJyE9pLh+PTIKhmiVpYo2rw42rECcAs
UmruS9As6JxeVojxNszCNZxOnZtUBJIFjhvMiPjza6O4X5I383pk8VA/IaGBjP14
sioxjkGGopdTpAkWKDKN+Ls5NH985lx9xJSW7/b9htlFubIJpimzpHIgCSrbb4Ww
/rBiPPWHXZKgHCW85Wv7xridE5WAPqoEZuonVTb14MYiN9Hmr8EN1khuPa1R1om2
BGjRKVEPxiJsHwA5u3+oQD1abb1hv2Ne6+onBBRhF+9Htau2idOzcFpbQw5f2hpL
qIQ0Z3uHifCdbSAnf7E5NP2+v6tDol1SvMC4HRTNWQmkYQvcWuUGID+hXoJFNIzV
YzEaE8whI/B4F33f+UQOp0jc4zKY4Sci8qpuW11PhQ0uJyZ44pJbf7yTmgwY7wEY
DS9UdQ9JfJmK5nzFmWT3wEWhlqTVHv6/CkZ+zJfhGklBI8Wssx8lfvEVIAfry9MZ
k7GFsYJJKzqPJxBZthmZEF1AN7QxIEUXYKqefELCfWOaTqrjtg9yPlHQgM2DVMrj
e0wNoNVgN5S3Ufr3eFad81nZo6N1WkjGPjTQ+XYAc/YDvysWDgvBjVjKdkQnmlPV
L3zXS4SihVcrb3qwJwTr+37MGGYQEF4XQRyE2QgcfG7fmsVtJkVIiHWNyVqSxI27
E43mZKKbW2nHduVzmwSuDK0Oyou4ttERab8dgmvO/WLncHlfrjPdkO+pK62S+UfH
cW6LSdgdqSbMoOlyUXTrBTurexGOuc0kMTFEc4hAvaKIMK7gPx0/5egN8N4sPXH7
XqWNeMHsroNFnyNT9fx3h5GhvRxyzV25fVRydpjb/xoRleEP8BVv0oEiIX+uj6be
V7yp2O7kaD0TrtCV0KByDHJyv+JYfzEAKMR8HrN0QLzI0ORANph6yyWsNEzP/kdE
UpE1YZe+4ogm5S8h10YQrc0e083vguC1dq/yOwmVSOiahZUAnUknetXf52J4ldXc
InCyeFFMQmarUkNweM6goTCYUsLFE3yCwdWr4GqQpBdyJEgX4dMlLgFwwjTkt80F
FM3qYmmBHsSUJEi9gqwt1bkA8pnak2V3tgmT5LpZoqClARrxzwrXWQVmiliKEpTI
hCcghs5xQ6CGTkre1yVcAuk7YmnpoS1PXRip/SVYU036c/hnBpf2diQfxZ4TVb67
+RhvuDSPjceRDWKdmWjIHLFiVkPP90beNh7jvNClffCAxelx8Rz/0JdySPgo73a5
44SWNAW1uFtYWd61CeScDBiEG6Z3jfLVpquI+e0IPFn9QfvLon0eWaWbHY6aLXR6
4S5wrQ9OBRE9oF0jNW+wE/MgSUjPUTMclrGs86sAGyF0BjtEy5Arf11HOsbNCGqr
nGijdzoHk1zBAMkTxA4ZnBWzFafnZBM8H3Ar9Brmb0+GqFZfL6EP/a8s+Yojb1AV
vSTqYVPb/E3ptBeyS13xQEf3eUJYevZfoW6fap3ptshY9KCNi3wB3wcnkHymgwn0
Of1GVegiCVhfjRg8ezyo1Rif5caVOUWfiOESpAaxMHZ0dRddQ3rjo1tWSfUEHULM
z8p1Jnj/MV2I8jo9nH/DBsXH6G5Vwm0amapTZTSMyTQdTOwFhivRctEQYbIcyz0K
rieYSjDmN2Dq4s+cZF17WcMO4CGDMhWZD6/4VtfKu+PxLNeP9MSKnC72YGMDcFMC
GdzLq1kcGDNhV/aEv7fxo9arPOhORzWhNzPPJI096H8NrVJGXQcLuHqMNE1fy7oI
f1Zx+alP+DBiydlesDiIKTvof6QfOAJMhpSUY3vsqNidnx4Sg6XJmVhb3aanL2Ck
3/QA6KWtW+bZsB2kYEYWdNM2plfvX3nvum3cwchmxGrZ/9G5QF6xy9I2/+Kb+rjz
/7bibMJn1TinzohwhT9V7jG3fkVMWxgdmxsIKpB3cB2BfhuKpnXrVkG6z/zy0DWa
tIHj4S5nzZSI86Ox+84ZGCKZAR+9ur+kWGKEL9aGbtRMZSNvRVcwvSNjsZeyQ+Yj
xd3LRQnOmaiOqsHsDSpXNJig+bQ5gqdEIs4qp614FnSaDEHigOmHbC8e2h0+ZHeK
bsYQGRJ19coIGQLO0zEKnBm2XDafOyxiY/GopnWes5iNxYcpzFnEPRC5o+zL09Zt
ZWiiXPxTaU7N/tqVEYp4vxLqXTvLdi5RL46KdIiQex2ilbr2zrw+NZ01rJUwMSyv
nhdd5k+p3OpBhpcBKJOWm4z3mW2CDCdBEbRTZIX5D3LGLpSSddf2g4/GBWOxt+2G
uDMWKZo5cVpTgfUdNh5i01lh1CLCLMXgfO1wu4R6/n6+dYMOPD4I6ObmR10z9bXd
9qgM1Tu012+XBoF2jrhPoDYv13U2E9hge46brLf0jkTh3i8x+b4Y4teAQ8FWBJa6
x+HhQC9B9NdsaYFT0HbeJTz3ez0g2IDiALnc6nmSxCoqRsD0Deys2IgFMPidelTX
EPbaRdbuqAwCMRXTcLP1ZlFta7dswtLckDAlC5VdFNszrIRTVizbxDulYhfU/pS5
bs9Q4yZHEl/iizT1VnIhAk8V2scMi3s63dHrNIyy1oY35MHcoR2nfnURmVGb1dzM
WUqxhzGEqBD13nlh2f4AF7f2N6uW+QFCeZnl9QrpBlStzboEcJMvod4goth2IODr
TrGoO6j3fWa9wTVOfuJnoKQO0DjjEORDXTXGu3RF3zrBQyC+uTdpEhESUJ5qKHBV
rbgOEU5J1XFVIoXsTe0tgw+lkfzAUuMS2deebmaPqkK1SjCmUtZ6GDH2cpoT7xq2
BZXcmwFuFI7PoT1AvsMRtIb+k6SQTA1FUllA0loHs+WE5B5UXwphYggc7PZWE1pb
FT2E35F5tIhYhdvMvLqQAm2995N9lJI2nHMAl5Asv6Xh4J1gR6CP2FqLdPzZDOq3
pdfVtMfhqYeecsB2baLf6S/s8cCSewSNa1vi22hh08qVQtoN8kNhQc2NmLzKYqu3
6Hbi/vsxaIQTRFt/IZspZMHviHXuGVWXtEIU2B//+0en0tWG0Yyf21OdFaYojbHA
vLhWaKPCVWqYt/F1Js9HjAqlN7VRu2/ySjtv8BhHdCFQ6vRezvsVllMK7JSyfFU3
BeY49oGwRyoGNdKtewk9Ye7Su7KhC2N42Wgwcen5V9PLZWdLw7rZMAYBgL50GVuR
fpJIFWXjrDvO4884sksXaRDWgSSOyQIu/3VAqUhjHeSmvVHiCnDLubga1YmjMIEb
0tl4lmxLBwZVshr3jwxP61SlfkdcqZCp0o2sICSgizNV6UDpNQ4vTC562qKlP11x
YWVFwM2GtDiehcOV7QVLiGNMfBS898TeruuITggUcfC1xbZ7DzyME19L+kuCFcDQ
qGutKRMrvSV5PYr90eQ0xPhz28LX6yU/iGm803i+AE06xq593E23T51IjNl60Zns
PPBw/CsOH9Spxx193FIGXYpU+axycjlwG+UY/SYvYWotx2YhuBPnnyIsAoBcdStM
rCI8lqjmbYsZtTPSN4pAnun6naTPz6IOQ22/fRvoolsz+V5PC/DHmWXwB4Z4j+ut
yxFOJLF3HwlgIErA9bCQdTQ3hCGPEWaf5VpVLm3y3xjt2nHDP+mDeeYPzDxUmv9N
TBZxe1gsTyfVZYaffNvbvoPLIXM0Lb287+AceL1/4JrbmiME/vZyw0TNhl5hUf6B
MNrp7UdLWbTCJM96vKvKk2LoYti9H5WehN0+MFbG5fOAVFfOXGfukpaJg2RSrlY2
K6c/C0CUv0UICYBKuzvKKCvum56+6juwQKRuqrccG4Y3Zppdv8Cl7h+bw6rN/MOq
MhQ1l6fBb6Ik3DS6NEJyteeP0q/WaKY71RnIjysU9my5eoepgAPd85LySlhOGG1F
pysQT/jevP34RzD/a+SD0E43Yt/g49/VsToy0nebvaNPP6nHNKQGZWOkBvejgV3Z
TWdV65kKf6srYnqkTTqWo3bVEyKyLuqqV7BqlaUNu7qwp5e97KuhARilpXV+S/2D
/iqB+wp6mtP5VbMJWRil4zQn3SsCn0y6iu3ezXvh2URpzesRYubBanyILj7R3V7P
uRnWE4SFCyciyKJfXIWrQuhxLiaSAMIDIrPF1J6UxRwV92bl1YCLY2qW8wiAL7vz
PzDGRZj/FRDj6OTyTcpLF4uhCrzXH4lRV+7dQZ2u7OqCnVriniYB3sR1SiHIaFRF
M/OCBhSZhjjJbWmdVSM5OG/j2DTaTzVj0qtal5xUiMp0tkNtbP39nc9cyW5+dg+B
UltVDaqH8DUorxm+DY2EB1iwWajHGNiu8RxKQdY1FqAKY/yVENz8R3CHz+nNJrMS
hFhP88Jp8jNZ3ZJOaCVX8GZPr+zWZW03HDdqXQ3Jb6tVNcW4Xd5aKsNRdqP0aE6D
thn54w8fTUvWCg7fP86qFLkxclLgGP0/BUvORFle1B93UgjoqX3K4nJqQWFAM1i0
r9+3f5BQWJqkRcg3Iy/9I3ESE0Go3PdgrbOMgzE0j/8E5wpf3eL0w7xgD+yGEzNm
ZCiINSzKFUxYATyGLwnIFcz0/YaknVT4v+GUdCRC7owZA+zzeKlj9PXYv008Cmn5
3WGO7HE2at+gBWHBhi7vDTr3mFcAT23n6V00VUe5ldQVarRz54UfNBI92mHLvBqP
1W1QNcijYWzNs8CyoaJXPC6S+gmhUr69qMO7X1DnCdtyqS9dtIObbHnHq19WB5qa
1/XyVOiyj5zj9bl8UMq0HJ8MdlNVfM+n4hDSxjJyZF/sHp9c/popLXyIehQIekhL
q7te7frTs7jUH/2dP0a+bdI135aBmz6ic8m1x4lqjY9Xcgkd0VF+rawlR/UFxwz/
gDOXmimnoY3evjBvwxYimffy51iSfuwtXKoPuIL1YhIAm+z3Y3e7oVYtiZz01B+p
E9Vd5sTqC7pRSrwb8eQIXLMqita5eB5atuz9PqHBzJACAATFc37l8xuhN0fpRVq4
FnEyLo95r63oy5Bn6TQpyc0nYxSo/0MK9diwB/J6iH0zULLmG4/jKoq87ltZrwe6
fcleZiwhbZ4bgAVLjEcoShFC2zYD46sb58G1mbNwtK+86G/Cb0rt7GHnXc5syuzA
BljGD5odkpnxIOhOL2tHUwmSVyKsJG1mCpn2upUb3sRCPEkUHYHibakCAD+ssvlh
c4sxcYKfGE9thijbK1ZXisQQsH0Y6fVtRHku0cPwWaS1t+/ux3CzZqZ13VBoE8GM
PyWepIOiWZkLDapJdIV70Iq72Pg/d2eVxTtjfLHsV77Uhl76lUUyeEr//aFkQPdK
0ng7y87ODIVYygu39Nd5cVDySSFCDoeGtrfZdPuTzjv0X124zp50/1s1MSU6DEpU
EW9P07j2FmwkRn3fMmXHx6E26Y9LZ6de0wtV/L93H7uA1EZrclB+TfSPhQHpmHgz
IlKiuyPZX4bWcBQLroqnti0CwGDvFfLUevbBRNd0QotDcwKYx4+WZG8Timwg0Zi8
KjRXpIXBoRhWQAx4T0DxtoimQUgNoPCTDFsl1H9RKy8/0v7EC3Hpb3122hkdATsG
y6SwojbYVu1dhDtM54/x85hj3y7f9hda0Tum2tqkU47j06DmhfMzfLXUiYEbtTvD
sKVUPv2gTjgD0FmDPXdIWTD1fLmy/ELjGBdSmCUmoFtpErqaos8pDubqkew7Zlhr
rCFibnxAXDOeTlCEQ/XownkV6VGyVeMLCDmIiXGTIdvwYs3QZfV1roMRYM+mV+zM
`protect END_PROTECTED
