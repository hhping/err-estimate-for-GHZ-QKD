`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKMoFjLmTnh/izQXERkwBoAwciPOLDrZibEnH6rwk0WBF2rl1MLBQO48+WBYKMua
joc6UIQWwkXkeVMvHmBTVYIGnGNzMatLG8BhRK5xFXSLeWUOgcolxazKMJHdfwoS
WqkRh754YS6X2Q5s6gzdVzM2yUBGsuRzxnMeq8p9uS65Y/kkcco1CyI/E/iaONXl
hbMGSYe4RMApnjuCngXolW8Qx5XPX8ke/h1e+RxJOhQ0erk3+yqZA0kfdg3xOPMs
rfV3KjSfhC2VCAxDV7tj685CXpBYkfsuUpKpaAthvOcyd5F+BBNmwV79AdlWfI/c
beRREEOGCtthgEREC5U2VsDDvn1DuO0l+dIv7MtoOg2Fq92uM0oDdQVrY9iGWmJZ
vltCyy5IlhiykJvl75ukkA5odtkBnSiPK9ZyJdhmxpNbEO0D2/XMfQ6nsJqRv5dx
vANnP3a1x+MKDD4IQw657p/i12aVvCcAM9A7Rkx3gbSeot5uUa3NwSkK6eztjBP6
41NBohkhKdlu/vrL07cdiUl3QmWCt6I5YkNBXL7/XfyscX911t52sv05cpMK3i9S
2qbc02pjUktw9IfO+3O5eSkv/fkfVif5WuhaBjJgUQFEmg3lzhp4q/RBF+yHizP1
BZH57Z+P0sWBt2n1gznkFkgI7PMUZCfmPU+x0Hm6nlhiDzwl0gH8lmwxOn7ghAz1
v8Z1+Yoe1JE3LGEykxAOeVnLJNKBsueRm+yMl8c0gJrtmXJI350IWjej2rJywyY/
V1yYD9klK4eqXyaneCBtJNWDdem+CfmSs/TXpdROaYM8uk+p00oV1qkvB4HRamcI
JzpDhipbpgAFtN050XjUGHWONopLHzCiNwVVGIs3lq9dAsuU79AN44Ses4YzrGjc
wmh368z6ydjWGlFpKt7g/XsGPC5xiDeEE2/JFiJo5XF3kjAFP3Be5ABAVO7osZNN
8bBAjkxneWxJPEmngEmyNBPw6PVRl1b22kyUb/ist0Cg8cI3dhEEZ5wzkkRXPRTJ
1HPKVsI50Sr8eU2xEtDjpKRx49ftfYVI8TVQuaP2gg36A3HjPE4Tvm9UUcggqb9X
0zv8IVU+IL7LPJu9PdbTWcYccu9gWK5QRLbF2r28hHAV1AcES4r5pGBBdmsa6Wrl
U3ReBVJCxEnyCLtQEAlqkntxWsLXEoOxQzSdD3+YNHWEYzZnguoEI1uW30Pjl/IK
r0AVCYE3pZdatdumalo6h1VL1CWVr9CQkG9qHltC4ewz0YJRxiMGJh+Xv15Fi7TN
ynxaJpTQtpkHNk10TJpnKRlA1yv4kVJmfOQs+6RQdv4FI6v7baHZPMJuUMeJjN7n
InUOIiToXSoAqf8XxDNEpSvV2Q+Yz2A9tcWOS1OSqoDJJbtB48rdrBNjNLwFyNtf
gFLz6Aw9ibh/Itm7t7/BRXMk++Q6KmViQkFvGF1IPANZM6ctwht/HaS3mR42uIdj
+5hQ6S55lPDAq9K1HOKTo/eVenjhOJxeffwSCqgqiNrmOFB+E1gQk6q3ogv9ZRXG
vC2RWJalgHAq2S+rN4JsudvtVzwQ34NViOt1DbfizUuWKuUauj8fEXs9xhZIKApo
byBVVgRqye2u3Bw6LcXlr1Vzb51hk94yaHhMJ5FdxwOQ04vQaPRKPiX8YmmH9vj1
aEP0lAN0OVrWjN96vkujkjAGLwccYrqDTQ+DJdwT07L4fjc/60FkrMwZtBwxRT7q
nbqCSW2GmYH86JU93SGSNZVRD+2QVOc6aIp2wPfZIQsqvXhtLy+3eqCDQDl6PWUc
hP59ln6ZLy3n7pY5oAmFPvhC5mKxnD8oz3xPhjw4Vc5mwbMh/VJK3kFC+OludvTx
FjPYXpVpwZhGDKkzHV9O/r9v4BYEIaP2SOOMMEWkQOiNBybvHLFQDlgXF4xBD7pu
Iu88Qp7bHc4h+0OisI1KT9rXzE7htfgqKJ+zbCJNML/gfAsISNFhgKAK78FjjqEW
SefiajUUySD+u/F3BGzPLdPVarcD5FRTlE/cQ0p+kqaSzfqwzO7gi/FRWOSxJjFv
0gsphuy5nbPfCzp4r+cq6xjdJg2UXSyfQ+ka9vXB4QaMaBUj885ALZNJV3R6Bvxo
Ev1P36/PMGx3cq7r/+BhLMsXJFAvyer+B01uQ3O/OKlYAD1Ty7/hYAgDLPWMqxJG
eKBdz67IV/EgYlHMOkV2Rx4JA+FC+1fldoxUFpcfwuaTTdRURwBTu1mMYiXZA2QO
V0CYGxZ3eWughgFaGPrmopUOVzLI+YqTct+SE0jU3EY2BIMh69rxhnE+FT9xyhcQ
5vPWwwjkI2Irqvi7jlo2IkFFy9ZIr+5e+WM/g7C8A52kYmrvBH5nn3YiLw9zfRzc
N2PKl5gbPy6wPgPpaooR6K22KIDYJdhJBZVKX5aRv9h50pJbuLB7SUmWfA06mNya
uE9xnv1N75YzPx71u6+rm8VKCBN8P72WZNHhtK6NSLTvx/ii0oenmjwpcNjuxQux
5KjfpFihZx+ahdbdfh2P2SURLWAoGfKsWtwNj9+J7Jovnof+VGwwc6aHZO7O1eoo
5tjktV/oL7nmaQX52bsU50QBqURDCw9P5uQy9yuC8SnF+4vUzqLxO5CXKVojrmkC
9TR6gOey2n5J0PussX3WIw==
`protect END_PROTECTED
