`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G41413ZZSeaEUP73GQAWnjJ8iTeOY7fHGumoKM4NjyXgl7sF6PoaBxzTSaXQSXDX
6HMJZ3lRhhQOHQYRnnODlEe+LdQBdOiH/ROLrX7B5a8wwkaTXfpPeC9/xejP/w/d
Hj/33pF9sCNJCIopREE9bpK1YOHyhEqt3+3Jtrh0FUjnsrDbJa70OA5aINdkHo/X
RodsuqxhPpXfVex8vvJxOu5xr2CTLgEflh8co+r6GtfrCWHyfG/FK+Y30cG9H3Zn
q1aafdDNomx82JHTG7NE4I6M54fV3J+OXwJsUrDrKgaK+fnyqJuVgZZPx8hZ45FL
aElfGdqNIQ11eVhT73hwP1hRI6w9PRxSbWMdzNCtsgYfC6PcCNjvITp+tZSZKkcJ
flmGHYytzZT1WhztQeQ0T2MQg/gQbtUriXDpe7X78mpuwjTC2cAAUtuMIFHjq+1Q
OOVTU0Hkvwm9iG84lmpOs7sDncrDFnlRdYMJaI+z8UH+a28jaM83SX0ZM0KF5nGa
IG7SeyMctmDJ6VZEzcXhKHmIJH7a7DZ8J3+SOhWc9WtACYs19xmf7Kru0JUXKVOA
oYLNHf27990KNOxP328RTKQQ0xudn9Ix/exQak6KKxfVppraMnI4Iz7CljQujtRP
RfHUqPv65HZdsk6AmrXCszGPMDQI0Iolf0zolAv5JJ+KU8tVa2qg7WI5t8FU5Kje
Uwpm7HcvG2n+ivxKSdtsBU5m6HQNoMuXfgARwUwCwaNRS3EXpo4+OiQlcyFqXWtk
LN+dbpgoJ/FThmbpjMzOkoCu0HlTn0hOPo8wOH4leEl0zZ8tlT6ZQAnlabgOZ4d/
UmqUY9hUrkIy6xlYbKXnZHq2tH9DgKei+Mu0ALoWlWFWHYts6Bzh7JtxR7yGZvvZ
wtLDHZEuQ6LQbTYY+ZXEMw==
`protect END_PROTECTED
