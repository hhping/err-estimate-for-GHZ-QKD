`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Bq4m+DXapg3xMKxRNqMqhSxARmw9/DrFo7qJL9h4IACm2rJtRl9kqex0ShHvma6
x7Bp7v/RdYcI+Om7fMD53Cv3wyFq6twrYb9xXOrP5VDkhc5NIaxxJ9NeICJnYksv
sLxHgp1ke+DZNhCxciQS/oKGuDqdE72etNFYoe7dKrNgzF7J1cAK/sRUImVSkIIt
ZADw2VHoPz1M+NtyP+JPGWDFZrN3+4Q0fOHPf0z7XUL3UJwemWkQqB4AZeM3Htwt
5gtvkGvFclgqYgRUsaXoYP6w2YkCU4q9WZAWKgCXW+jt+sq+wHi9kImOa0vt8vNf
olN8CCMYBqhwdvRczcHzdSvsBFtIipmDT3ctTw7+N6zTrNc6opreRDfM3q7piuU1
hnIs99cb2kby42htnkJjeeMPjwsESDbM4uFkJpfTy//bhlZMhmzSUacJliyfpsNe
p0VHD8/+h1LDHAQf6OX82pSAEUa1RZNlkrYsq5Ln4Pfu2U1P1t87odM1mHl2BaGs
pxEuwVxsn8nlDHjSa6RgpBC8hvvfCopQc10QsPDYejxyXBl4H8PAFvHBKACjRNWc
2oJrXvEp6bkM+ihZQw4yMTIEfgwXeCVgW1a909xGT3VjUN3qRuaX+O0BAWbjhN8z
xa0sUF/PAuowhSD1HbfAyULsMUBCfaAhugsHjdgbnPavKXPdYyZR0FXo9QbKISuV
XA1dR3SrPIv/4RfId5tJMqI+/p97Lds94B7GBxvWEPiCnMKPThd1b+th5/AtFVjD
fBZZcwmlyBtq3zPmJJd1+XpQklnugIcRssAjoalbfwRJR19Oyl10e9hy0PWNQ8KA
nvfEz8ZC9oJfrXwoa/DnXKIVcwVC7+vOO0mHUkdrxrjWQv2gzDbxmnMvTr9v3uLD
9fqeJ+cTNVV2+WjgCHx9/FIzRK9/3cXGWWwa+iiW8gWm585TvYj2/OPEbTEj5ZfW
ilx6+SCaneLygOHafWBNhuk58/qmIlJsP2TnSMxlZpyw5veqc/om2yzM9JwoA0gV
tdRw4uopKTRpogtpAr7l2Foplqz/wuG86GPD/zXtK/cihcS11e0gncTGttyQ5idO
nL4H8BrafUuyC2vEg+9IysoDW3c4JivFNsBSOJnWBnUFq7JDy7mkYpwzH85utvFY
FCwPUZyDG9g2rCiKgMAxfyvUWuC+Ej6jUTd9tcfUh8AicpKwNpIcgvciXGpJXbkK
+9H7iF5BjfYUpKxO5BM4PHnj/6KC1TekyAfoedgpncOMh+kSnEywbTEI7n/oLLRP
x/iHeJW1AR2nwnJV+o1yOBRr6JMfksu1tA8/Vj3yPiWQOgdvEZB2Bj6k82nJCOw7
Kr87umNsmlvEwTsP+ruLDbz4PAgO/4Y/uQvrRRRu+1SN5q3fYCzBQWxVcURr8dFO
tpAYII20kryjlXdB+Yg9eqGZAy2dpjzD+4XkMU13vZBFp6KwoqjaKeNq4AYv09sg
qZQD2eoX3FJ6aDPdZ1wBVK+IonhF/DlfQn/2HbYV2OW7XTKKtHOfmYItmEC0D39s
H1Pw+VBhg6aSCvKmG+zwCFeUll0IQV2aSkFhB8BoylVRVx1FuHHNMevyQv5Mu4Cl
`protect END_PROTECTED
