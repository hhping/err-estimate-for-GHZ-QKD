`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKfR0suALail6bRXu9sJGNRsmKr7d4gPLmebDZ52sZdIXTZVKIS12gaGDym4YhJ+
2J+tdJUxdr+tkjLm1i6K5yofqjFnIi96L5/j+prS5gM/5F+PhJ1F9nBnz9WiLuVD
y9azThNWHBFJNcCsNDRHfwm/uxc6MzJuc45kt1kOv1i7ePxVN6yLC0IWsHviS05E
xMHwqm06P0vMoslgBo/7bTtnMpNdM0yOeexj8QX9rQp6x62yjkBdgyawveOz+2Kh
Q2G9+RDq3TW4ma8bAe6mLNvHWGeb4qXxBgXuAe+1m9hyMghhY5RrokAqFo21qC6g
MLSIKTVivn0Py8U9w214WZyo0z4w1MaxuwX33f522jJ2/Oxmrqhw0g279+cIwI/E
gNEfU8sgfr2AR1p22ZILWA6BRDspqKZpRhMqJnkHXkonp09S16FVvlKnriOOt2mK
jSm1R5WQzuws107uOGMhpg==
`protect END_PROTECTED
