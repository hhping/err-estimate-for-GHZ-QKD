`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uTY1qpum6pn2tfp4LfyYaXTUgErIEJnkNU6D7125hIrD+TmLvbM5YfwN0s5LPurS
rc/S+Yv9e5GdWOfD1hl3uxQu16XgZgSZwMMvulbMiy8ZIk0QWfooRSYf+cqIrXEb
YrSrUfa2E1hq6lMZT0e6Pqj7vkRF8dSSsKegYV3MvIn9B7vourFcmbrc+LOLvjw7
LywAl+6C0B5fWaRttb8kPMEXjGVSw/9q9LIGHmM3f8mnEO1OZsuAvzObZO4Apnid
kXcyCFOkAMpMgv8sgh74rkbzwpHPjNkC4rZhBqNgpJPaO+JTGBvXxXHzdZokzxwt
pCIdGNa/lMvZRJVTfuhdriJML8sfWNmWusolCI91wM30/6GBx17I43xmskSnA8N3
H5oF1Zj+XPgSfnHehPrPUzQUToTZ11RRQ5Cndp55EJW6osDZeZDf3KCelKCAA1ax
Ldm7M0qPykOyVl3pTuZhVobIHVMAO4gll131/m4FQXTc3GZgITTyAHtnQwmE4NrZ
qjhru7zGnSLK443YOGQdtpq/czzrk/d2ea5hx1WGOksV0a1OTAyzegpYzHfFhba6
Yx7vt2efoFfoONm7+7U7BwLbK5FuiJzZl5hF1na8ApUDFKpFLwHOJ6oEd1EpEh4A
IED+eO1ZKMGmPNhlQSWRWsEf4gC0LUtSUpuU+ZosU1F2BkYNFfVKbf4hiDKFEATX
`protect END_PROTECTED
