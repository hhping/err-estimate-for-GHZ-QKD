`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24fbTYnjpKG6Js4OiIYjcYbvw3VG/+5rqYZDfOBrX/L6GgQ7VAvPoG/wYNMdhjnT
RKwFDy026m3jddxqSD1eFMYTnkyzn3Q3xMHSyDwHhcC45Bp4EBIcJEnoStMJibS6
WGfEJdC/9Y6ThtYgLtjpMO0a2+ky5parcsW70eHaYqFMYU/Ydi7Jfnr1VzB58ODZ
XFwz26GkDqvV2nprHgoj+kXwlWzQe9oJ3Hxhu9h5mcPnB0WVd8ZRiVq/QVdAXOIH
FRd6tPDSadFHFeeLaMutIbWBzlNISh/nZPSsckm0LUpXSKigC7cHvPJ0ETPfAeMB
4e0qIeOgCZTK3g3NSz9Xwvz83FPDP3xiKMctGbh9PDPiO7ekY1iLPkdyJYKF5Til
LIT4z8RDusGlImQ9aroG+DTozMTE5Aid/d4oPfMoa0sK8rkO+qIjmYSLZFacFAFW
74Q58MAnvCQKDBDl8nkqqge19A7tINktvwfAn2fgMv2g0fPqMWbGBIIIiJ+6t5DV
IujZMIOKxP92G0wWdQU1xy4nrgQ/xQZZ3w37jmd/obN/SFYH4AAGvuwzQML1hkQn
sYbGMSgc9CQyXGxQcS3E6uKOi2PTVcGyvA2qr75axCmcZefpIbh1ZxKW0TJA/d/u
v1MrvzX5EOUjzBpTWXjw9Pv1FfG2zlg9wVXWe9OroOJBC/pHB7UQ6YmRQBGIKeCY
ZgclRwGTCWZS54Dl68hKiezAGZrsu+q+jVqsq1td+Xzgn0imbgCzuXVfFy8ssCSm
h71iThOZC8N7a53mSMh55Ji2GigzseDZp3h0GIv9sLi4QXJ4Wxav8OlhEntH0XbQ
+k5sPmhVg8K9WHwAEfDu23llzHHBYKNKp/y3SJ9rXbRy+ZoEP/rTlB+cZF2akaHW
iUxb/f0m8pww7Xd3juy25wCQRZuw/SR42Jgn3ZIyvJP/7mHuG5DKxKPXDXrhZQmK
DvvLjHs1wjVdv6a4Q8djTIyER3huINL4CAKkG5MCWUXwvkQ6L2AuSFPWKtLHRirP
WUbUt3hrCDewiFrXjHaJKiEKAgoCULKymQ7cASr8Hp+B8U51OVA2EKLvc1TYaC1+
gbTJ/BsdR3wkQy/gv4eMjJ53fznMdVpvF5FgT6MPa/2OvzGQiLXaC0VYOde25vzo
f/4XNYrn2etjFpxB00n7IlSrPXyKrk03BnrPbqXkG22sUPi2bLCIUoc9/5pysKi/
WpqxaB6noOwN7JvjvS5EkwdWcOZwbfY0FkN0W+pnn2O9+06ekKHsrXaHzpJ21EpK
socFHpD0bvZJ4ZnQW2QNIM1XKZzT2a2HyBNliIvRYc/qlxGcYCEVavko33GJFrKc
xvYwkNnkHpFoyNV+Jfeo63pZXW2CzhqqZPQ+sVVeDrHMUtaqHB9OnVUXwT1cOcBt
CoJ4Y4a+20V5xTGmjxCjHBn3QsLzadLq+tXdQeP3ARrmgYwOQ9Gv1vTHGORsAu7I
fYVkgF/Qcm9zzqVlcwiOZinXXafhz/yAL9cwX2UjMI4AQyHx8UPIvYD03x6aXR4p
lFHe9gSwTN91KEzUSBbO91WluyTCCajknsmpP1LSJzmQuN0oEoNlwHSgVjiOVunp
hMBD7XwVTv0Zo+LW6LE20MFcMq7CWrCb3LeddloUGapa4xYYnXoArDKq5JPg7TYE
kd0IlnvrhvZv2jBBSH6kF1vwx/JO3IoWi2kF7RessEEWUPhJGAsdIBT2G/MAbZff
LBP0OxUMMX5JFwqpDg2vYNltrahcb41v8Lb9t1/D7A+MJ3R4QmJvbX7lJ/HwafQP
HA5hC6MAnMW7zf1/Lt1YoAdpZaOvnMAy8GGEnO7WvlBpi46b8O/XtlIrrV3eKbKj
i6AFKrNRS9ajfG4oqvOmWHHwOFHTvH1uOtL2z22d+4GDtLDOyitltTZVe5HEIvVa
LsDiSrc37+mje6QVlyKmzh+5yB9YCX9+6LzgwplALgJJBI4dXcufRR5utOUaOZ60
ugP3b77SVcJ+04V9z2rrvgdgoXar+bF26dlrZNBU0LzGQlWUyGzqDveP7/Lnemn7
sVPBInA+tJRWS6a6dN4HLEbK1dpZPzFXMTsvJ/dvhLrlIE0PpclBrGFb2MHOsJr4
PvUyNa19OdS11/mKEkmVM87AARbCAAlslvhstswfcoAz7+tGwgRhAaz2A40Wu3Ag
7VzovJ9ycNtN7hQudtT86zmDfrjah12bQ9JxDdgkJhJ0loMYvXMnB3LllnweLjf9
Atw+WUj0JCEIxz1o8xniY12kxdFs2HcnFkYCIx60nNpPKJasv/R9XYgiVLIGDWQ+
tZA4A09VzYunHLw2m8maGICuNslQBZKy4djfQfnDrnvtU1A8YDuDd4TofThwqpAS
el/+aFI/A0fllhA3lpSAxxZCm31Qn8eqzm0urP946POz7q/3AiBhetX+ci47udZ2
U3ErlP2jjfl/ubkIn2/QZ/0vt1AswLLQbaAT8vTsO1ySj5zR4iSdWW890OU7yIAv
yT+ph7W8BQJLzUzVSiwbEvsJw+GsQZLC7sOlWT/BIyNN+tl3g+8AzgNgKbu/DcFX
G4ZxWGnB+LxPzNy6C11ThUZHX17Jh5hNel4ppERpVqgd4Jg5n+S4n6VQq711S7P9
l/xB9Cfa6LsXYQTkHKyTLqLQvsphfjwzLrhYBZC4bTW9urFKULePxzYAmGQBVyfW
gbCv07TZdLIE8GQsfMJYjbLTu9+7qTrz5uMSIOMA3zKtCQsASBTs1FOHxdRj+XFw
C5hGfmFRK0uQjTBCTf7pgeFV0U0RsWMS8q4TW1Did+Xjra56n9CioZiP8cuTQFUu
7efp2TYf+oKKGbgTlxRDQhZtwGXvOy8EW5yMJ9ZnYTrLpsogTcr2tjoTd0AJKwbN
eyKC6J2HzmDOdN1YdyPRETgkNwBEn3yH0oSbctNQWR7DeZDNdgVBnUMtxMLHpHRW
yqGE3IaVQL3s5d8pcPHRZTAwYe+WdFjWp5Wpr0w+PLjw9kyknlg+tpD+q+bxJXJu
Gt7fAe7zSxCWAFxYOXR4eEl3PE8gOQcmih/wLXf44XwyaMbph1hIQZO24G/txUw3
W3fFnfomhW+0+YMRsLIocXJXN4qQ4ZCKdbwLoH4oHJmFV7kX+nL+G0PaAm8ip4dy
rhFG/tqQaefyOeUWpaCQ5AxBfns5MZLzvXTdrKZiq/lfzSo5CelVPVd0DyJ2w6+X
6Xs/tti71sSv0vlBCWAIbTNt8jNjgRs180Zw5IgX6oO1Y6X2sV1SNEH8wFRltWvj
eFpDJsCm++93qTocQn0V55oh/UWbzl4AOZtzU6mFptBIUGI336nqbF7kLdfTsyFp
bJg17Qc4EP3PbxO9YfTcCeN+5sjgDYEOlPUJEemXCsCI4F964n1vzjyv0MPiFK2e
HFPz5AbB+lcZR/cPzHYQb/YxtJyjdwXUYHpAVucN324maYdieas5t2xHAhnuJiLa
AG5NlmopvXaDi6wfezm8t2RNxdetVjPjTIkSOckHvddmFK32+487uNJQFQfKCxij
FOR9TAX8dwxBmShIXW/plQoSls3yQP4v31ciC9+amoLR0lBJwHGeij42N4fsDTG8
NYqA06C0NHoDX7KsVNnaqDt+nIEhcQiOVa0KsTa1YTw1frdgvEbh0rAJAvuENL91
fs3P0UxEK220bMYfmBzqWpbf8GrAY0TCQETQu9X1mUuwtpaFomc60MZWa+vFLhJ4
+Pse70UkIGKDSk4TSkCIdJ3l0W2c5a88ODaNKvTlV0Flb1IoKTt09dVxKXx01ql6
bfxGz9Ha7ItcJhZecGK9d+lfxtcc06iKu+V3ryk6V4V70tZsbLBBosQYAnjJRTvI
qplmw1MZmGUCkhMSQ+mO02FZd1Tlgz61pb1KQp6CpcMqQV7+ExpYe4VsMMweGppN
+En+88XRiD1+CsR35Wcq7V4/2cdxEXBqLSACvJcPSID517ccxswCCowtmGx5hLtK
NQxHo5EWOYIbJG8cZm8dQEugzPlPn++Rl5Q/L+jiV1ro9JYhj/x8hO+Jan08japR
hr6IfPRhRnTUgMIDeSDCyPzexzYMLSC4Kj6Ay+8RQX6343L/B9IQJwtN62gQdDNJ
PH6AL5FMgIhNvg1hvcGt02oIfh9FQEyUWB8o+3ydamljYzuOyQ/2lZoBzXUcXyi+
04U7RTZeujfgOk0eg7D6toQXVNT4PdTX2prCx34hkizBCAPgiaiqk6yXgDHpxvvh
KfYGDr+Vr1JZH63palo5CIdMAYYjF1BZGHf1hBWYHiLg7EFsKRoCvNc/JX2mZPKq
hV3XvM2Hk3ThcRnrg59+FQ23MrXB+meOpgaMpwUijlFqQTd/4dUet1nmbTscullF
EMSaH1R9gFmXs/jw9C6l8MQYBL0+NsjoMpt/dRuh2lka457Np/Ce67CKFlgAhh1f
E8BMCElwtgjHKzDBSoDsYFPM1KOHcYaHUDI6AczPtYkSrwBbNN06Nr3AgKlZWg8X
FZjwRkBgt11v81rU+M6h9stypqvdunMylgfOJnRriTR/GpuWEW/zkJmNVdSZbiZx
WJrdFFgIt2YjDQXlyCKRLqo9rISsLy9NNo3eccx/M01dwZzPbQ9R0Ykz6vtYHVXI
qWyAPRP2/Oa/evWq5PoptHGl6bk4Tjgq1lYyM4OlaQEh20tu/bXOT02CxTSP6gb3
zfp2VA32kKcVeLpP5B4LhNlCLSA6oTnUCaYPCY0pUu9ksv/UYggAlNHcG/IdCLQf
9ItZXTPnHbb1Gct1CBusNyOyIkZor635L1/PNcht6EFTEUEoYj1IKsxTWOFS+j2b
j3HkfT7AZj14SO0aL9qwJ5vorqW6CEuPBzPS6VVGLHV42ObzO0+LW9MqC8Wc9k5A
t2JfhNZ02WVcxAYgC8KFMClEsNsII0Lr46RcOYIcVQqRP94zz0XvuaCm+o67Yc6F
j9Inl4IY2HVST92lbUw0fHnScq/iugs8bo2627c+STccK2q060GlZjQaQYqNAQ6i
qPmQOBBnGKIBF5Dmdp2NlQm9vsL1NFYqPluQzb7Yg29HupOJ7c5IFUI8ym0BYutb
ATj4JHIQuezNOJc/jAaJN81b4dPDrpo/XaW1B3B0iIJm7fz13AVn0UK0Uiw9zDc1
6+aAc+zNqmBJQEFryAHaB6uKYU8jrPyMUSq5Rlnho1dYpLXCxPaVnYsB1brD/+vl
1rzPd9Y8E3dpFUcYKSySm1Efok8QNEhENxtdrGXa1xwp4S+Zd2ulPj5uvSmWuEJ5
8mXw/My7qtTbuz5hkYRPDEbsty8GWwOFaGwTHkKSPiL1sgHJ6EHPvUglEBwZA/wk
xE64DtNVVcjbQ/QKHPMykGIxp3keezez/kAq8Dot/KPqBhjzgemerGXGmYI8AO6s
fWIrca0YQhuMUpxKCVv8PeQe97FyU21DPFX5VdG05DAluMs9OiTJziut5u1Fl80B
+uv3juyZzkdz+8iQaJWfhY/BPh5oPI3n1nwaO+t7VO6aEGVbjnYmY07wHPj5fGaj
7h/tz2iGjvIL/0XlJ3Jedl0Om480tKDnf7+ic6D1Ms0mfwPlJbFr7FJNgiEtIp4L
zcLLKiv5NE869nFx6erPTsYAfXUj0O4SQIhRAhrbRTNl60p8uMLfnO+DGMp9qtMh
vrI9yIaBIedYBwgT+aENzzPPEMnKtCy2gBbKgkbFP9HkCjq3OCqeCvEHCOVzs6ET
k1AMK5wpgajod9w40Y0OLEQ/EajC8NlqA/DPY5aUDnBJZ3xtcT1vsJ0cBePxKBmy
c/4ydbZD2Haaxxq4XUT8E7AzBiX/aqgrlWH5bGGoD3DIrrrjseZ0CytOnZgU4Md6
kUj0ihsySkhphVvcnYU+eDJLetNZacz8HtEtWcShnHe/zRkKr3fT3kmNKjs++stM
cJ2RsLK3dsYePD4TMRfabIRbaBXps1Z9x9FngpPYnKv3+3WMg+ZyX5icCvcVC3hD
yaB6T2XT4YJ7NQnT/bKDhp3fVe47foSiCSz0x7qy4nHkYAD9E27VX09Dmprr76nT
FqQCk/jrKJ1yfpHqfMPy+Jqxe55jDeZaH1f0tfsRdQpWdgyg7JiJiKxqGcfcnVoo
F8Z/BsiS6hYDUz7BzQi1yjb8hvA61iwSJG2efzA7IYX1MVmdN7BNHoinBHV95VQk
vi/TP4wR/2vpZ7ZGatV/nx6NJG/Fwsrkd/F5Ho9dQ640teb4mK/R2Br4ucgOaB0U
uCHuhej0mBWGoI3PEkaIBRdRqwLcaxIkDmPzGBz4tB042wdUS018ywRTO9hWZUP9
36Xpd7c4/ZeHVl1Q9+1veqiA/F40/WkZm+uWZiiI1nBhfOSTS4RnsLwucA/uJJb2
22IPqyuGhD59APj5ypfOwC2cmVN506DRjtIMpJHz9JePEc6PfwzzSS5o2c1KRqxS
6flIdpyHRYNk0Jru1lVjg3n82bcjy1/02/DGinJxhfMkzj4X/jtp7DY7hhUo93AE
OecsPDUQaoacoZ4lLiorkE77YAPYrjMQ2EqCrdUbBeeX31FDFt/1rAZ7shaiY8bw
7CL1nul1Fr48GhuXqmpkwyQlJ8NHIRHJhOZJjQYjBPEqJYnIyWFu6Hu4QB82qGfg
TeSY2C+3k2gITJs/95o9BVMFS7+hqFVyDnt1lo5TjoYlZBc89L27coZBCiYRqBbI
UtyBm7tD5kMHukA3TnawFnMWEQoHxIxozHdF93sKsAGIib90rW7SpLoPIaRO0trj
QM0woM3NdStdUYCv6WAYfGuc9cmtppIyMucWxBVwpMMqD8V15cgrxp+zauWQ23n0
SEw9sL2n35tQI5XeccwkEcwIlp6thURJ2YSf6kmfdFaoEHvMRfy4hmVOWGRnBOsu
sufYe9E6T+aug0NrYjgn0BD7wCPacfNjzy4PhCM5Kp9y9NL8Uu7P0FjDrIa+/5WD
TKIaeVX+sk3NTsNfzipYMdrzasOfpNucN/uZ6S1/j1d5G6d2/ho0EKS/q/Tsw6gG
AuJVxgSqkf+AXWvNnSlEbXOuOCIJ3J1OrO8+X6aMjnp5ClkMNU/LYLWp8vjKYE6R
LwmSdhA3H6j1/+tn99uEj0L0b0HAk5Rn13B95rGdBX8zQOJ09zAqU56+00cO6jTb
5OV2Ud3PC4pEkTFaZNdn1XsVEBtaIffMnFwuxV1VxsEZIDYraM4OE+De5YrpIe6t
V8NeLpvT98o7TMYgo+KGGcPPOECzqJBPQrBk53z/0agx5+d02vmarSxab519LJWF
oJgbrS6iamNqwP0PMjkxiPIj/j695GhpjwWf1nS5hx9B9rMb2uOBPmcrLcOg3V/J
kwi8dGLw8j5cz/u2eLV7CC4ktFuEsbQ1PLj4gbBEnZDDmsc1z+s3citoCZd3bsWd
9LWKD29Nf2Z9L9ovmpDlfk8Qu+4uenXuDQTE5GBbIeOzEi5qZSqIJ8MiYfrCW3o0
OtlntP5PJXBSpIvn6UEribzam0SdVDyD2kQa2i/AwFBGxnW+JURj4eC5aW9JHTs8
jPL0EvbwW/Y+jYByQZMc139mT1W1URjz7x53ViLIz7omMoGiQ8YpPqjnzQ5cQrWS
I8zfzKwuylnOgxAfwzmj77dfskwfmTqxMrYJXfM4eweOPDSBDRUOra1ckNi2azLv
qFKa2pf9K8p1jObRfObZM+3P6PfLEdhccQWq3tdraUbwjZ8n/FG9Ew7QFpCs2td0
fTmbq+0Uyp9BRxnOXJ4LEH924OCJsZtoC/ObkpRkQsleyqzZmx6zIq5WjGpUEyiX
tVUgL5c9kpv4v+aTecMITB31Klql5c9gp7eBAX03fdXpOgcAW1pXsWqSe3qip6DR
6h2MBWv/rB0AFsdNmNCjiA0Cda2cf5DtHiVSzammz80LA9t3teEocyY8LXznU/5n
egfqGFttjo8kjH7wA8ceNxv+WWLujmuSLmfRN/+ODckPQF9p3+nD0gZ6oIxSlyjy
78HsuILiUVCMNjAyXFmc0S1K6IVNohOQUUaKzLPAu0+xmfcNF5dusYjYgDUxrfW4
bmZefcb2sfsZo20Ej5WxTjipUSdGrwY3pOBbK78BTB6x8bWztCASkaJYHmWF9Paz
xws1qI3d/45Y+o3cAU93+EQet2jlVEkMNcNEWebTX2QtYQZwMCudnUCoAmuE5r5S
rCSVjs+LDc8ngSu8kdM29nQEAdtFQKNqZsOlYc64fc7biULlXrLm6Cf/yswIh+E9
oo6w0zhO33vsGDZrHNEwZMwBIcDfSyROa8C7luKFlOEX0DC8kZh/yTM3RA1Xcch7
HUx0+AgkE6h3fdbdBUaUcTvFTwgncBziZXTQz6+npVE9ZWwCLwGTrW5XNrTAu3hD
obWXyWc1FQJP6zq8NSdcBerD2dtT2mELEIYhjp4WUVOSRAT9G7bQLngQ0dNk3Fzt
bEdOw2XVFoz54ZzY6TkR9gCxJYcZ5Zelz4UU13puSePJrARCY88c5Hv6MOwsYH3k
G+3YAwmUufuHOvoR+7J5LS3FFfKExGizrOe54szkqpdys7qjg20nu3W7McSwmmI4
gj2l6Id2YAxdeG5rWofE86L5VCnSwa3t5mnQuThFUYtv90Rja0D3ZsuAzIQ022AC
b8MhcvDq8MVwbAmL0Kl5tF5h7xZ+E211fUMknwbaYLIcR2FIKOEyxNZrizuw4kM0
u8IYse1mUJbgNZCpLcDJCKiSsA/N1FRbUUzuuTHbNaJMs6VqrC9o8T8P/LgDIk84
W/6ktxXxjWe2bQ4wzmk9xrIf4nsOQh0Z7J1XkimofZXSX+xATDyddX6S/XbxWlPO
lYNLfjG+cNfzVyoQZXJQIudZ/vyng9FuSKMZ7G9Kd0/CGe3Q5Tp0glZRSMWG6UTl
vKzIK7TwUs8HWEgMs00HM+Zs6e3b4SLtAB0Og8ve7yRHnplqoHuXr+ACTyhz33PD
pJqrIbLnL6316tg+fodEw7EHevRJYlZUWTvJdWitspO0ufmynNAiaL83yGSWyMLr
1VvQY5Hv55eXCd7mHmCzDqo/ITe9Ru3PrMeFp1FvthNUdFBiWKFF3ATQZgc3p3E2
LMeuQ0hAEFV7xDYhiHmi1pUV9nMxNxDo84/WwtjCLwucKib2FENZICPDTV+xp5Zr
/OJIhhM1bJroParQs2UeLKXEta6ufoD6HGasQ1Nd0koUaGjO46VlXmEICIkleMn7
HsjVqNm5/OG+OgAxsAv3Xq445LU26zwiHEDgn0F84FoRSc+S2uXoL6D5qwer99x8
Ibr5l04tJlKfIMAVhn8ac/MSXC11ZYQz+YmIWy2ABLJ+CwWROv8j/2NJGRMFCIIW
cJpp+UKaMxFJU2wY1bHGw2l2fuLcF1d3P8Qv6w+ZHStGdTQBGlOY/SY/EZg82C/1
CAAiFQzftV7WfhjcWW9OGZcHJFwaDv143xHKs4IOgXdCewxZu3fLVccMh5sxpFAl
1WENx8KYyP27o6A+QmS94mSAtoCC0hwD+lof6RvJBGEf0jRx6b4OKyMBD9yUnQGL
2uNGxpPuOAyYiGVjZEcOp1xzsq26Q5kKlAUpsfVE68ikNXgjwWpCTNzVyxyyiNWh
bnrfZKD4XySonEWbTlP6F0Sh0B7UFeOXJduArnFRoepKK2zxqIQDUKMQj4k79pGW
jLuGKNYuvNbUNQVDQgZhhw5e0k1qdgMaUHyDI9gPoQd0Qs+QvWuvipkVEM5hU4VA
giAoZshNaSnY9/X4PaiZ9pFX3K8tw8YLSOcM5LRBOkJ4lM75yeslLfr9ZIp5cVXU
M8oP09cVzRXkWwRofQv48zHUYVRYMaSiRkgjr/JlZehO+bhOu8Xf+0FRMsI4Jbmn
4tNxJwv2mmmbMn6qoxZWQDQGCYcdfj9bAbtTa33SLnP+8e7LKtgbnNhWfRa31wBy
1VgY2KzBBN1w2XkNyR4psIQzJSmG4TfS2ahvBaOsPf77SSqkYUhweVv9JW3EEwbo
D1pjHNNM9iqT+iiP4ho6tYf1V8DvH6i/ld+0vBSC8LM6sDcbfIgHyxLFsvhqDHL5
dyx/a9QU+yOx0lSfMurVtrijJinzvT/goNIGW5okiKZxf2zBQs/gTjNC7u+cap1O
yq8478vVeeJNEYw85IHw3pdnwRH3d1rCorvfQlL5kkbIJAsgSSejqJ+Ig9x//C6F
IHXcEJoHtHTDkfBVZeUsUjvpCBVpxYyItzcs9iz3Kt0Gs/4tPAvZ7Uxej/GtGMLY
w3V8JtLhzDsGYSHTTtIFuy2rAaD2FdeTyjo+G1FDKeZ7b4S539xlfo7hJ4xcUUhQ
RUODn5+Q43vs0LujK75rE3n8BOGI2LHKYoMmeZuDCLn1wyhSrKgNiesb5pLcgfy3
xoZh7mOEAbI04/IxuqWXapjuEFJu1YpCtuDAZePonzXJzZfAoumgWnhMHGQJVZKt
6vCr3fh3CwQ9+vIARmO4g/6ijcbziyIP2XoLdlbuOzLbDDvGWbE313jVVh98cIU2
wUygAalWd+/AGCUaGWmriK5fkPlsy9DZQI20iaPRyTLCoNuzwHK12NMiyl053zTs
M20sXyBXR2OB/bwNylZZRDx6GoHEAw5yNsJmp4KQlrlJGdZTNmL6jyk5YJwB48IW
1PW2KNT1jZjNvIlNg5YiKDk6TW+/LaufXoVN9fJkDVe7+I+kJ2jPUIhc6VhZEkOq
SQ1mRJpDrFBtzQ7GBu1DqbjYU7PlGXlQwKG6ngX4HFQ4EC9x11J2gNLpV1vRwzQV
b3Q0413oX4ReAaUldmcJRaQ+tFLvIi3NRRuPk+Cvley3J5jC5P/aLIOhymTPuB4x
eNMPvUQ71IrQ1y6hJ2dRQ54XTJZk/c6Ua5hAK62q4lDmtZyc7ky7AzDOZZFAUl8R
PV9JX5fQjQ4hk1m3CaUrzQGqY5gu/iBkZTmj2NtS5itGf4Mqmws8U+nj21o234vY
IpW98zrf27hqaO0i3ktH5YGkyFENLoSZTwyL5OQ65mMbdf8FOtwfwcvek3i9eB4W
fCbGG+RtvNUP6PUfbx5Hf+9d5P8GC1UG5bPZPbqAM8kuJM2a2/hwjzlZdVs/3Gkd
jXC3LcfK4aSZCn7cioeABo51Pk+KzNsPBaZ2U8ANGsMKNCwX9zlYqR/3phD9mIxB
LDjEt/688zGBIZRYDX7OyFQH5iIScQLozlCi0nj26G6g7SPolU5iyM3UmTVkmkEv
PuU7R45/u97u07n7gp+ruH+1zhKiHK5PLKMe78lJ6wpWkIXCITjNbOcBS3OJV4Qa
8egpONbfVD/pHqlnXkVy/EmJfHWE23WjKypVbc3rtz+82eNmCd9u0x50H18ov9uo
+Db5hamZ6h2y2vDDf7ir64gQ/2Eyx9TSlFX1vGeX/EO+7dur+Lfgm3VklzNBCKal
6/ofuWEArCTJX14P0D/cPcI5TsoNslyP7XRqaaFjzwsTITy8LWLYT9/ybC4Ge1xI
r32hlaZ/Evsc4jFw9P8ZRomKUiLYeAJFwjoLH3sKXA930pfpvCDQJYs1BfDtUYmx
ji9ixtDHKqOzkjUYzxV/jJQjc0UcJfleE0/8rZuh2m/iy73xjc/Bks4PMa7luTgi
HBl5mRNO/qsp6jX5fc7e/Mz26qplTu7WU3SQh65ncKNtsLVh5QRzF3wB6JYilwOW
LUE+FfYwNoKhBvr0aGwKf+agKB2/HI+2clCnipJgQZUabiPH/y1YTgvL5OacEz56
i3q/r698osiOUHBMWF08Wt3rt2IL0R2F1/wbPWR1HwisZyTNF6bgQb3rXxar4gxo
7f4x73bIc+Hmkp4Qybeugj3/InZsrDyldLPh6IlreRRK3ULaU63BlpzVRqFqhU2F
YmPB8Ls91Cwya7xIZjL15D2CI/EMInyCy/ALjPTh4JlPlFPYBK3zY90VXbhpJ6m3
oFgxSZVWvQ01G7QfI6sREbfWfZgWKN0u/KCH6PSQGI1xDgBM4xjNcPRWdDTvL/nj
BTtUU7dfGO8vVrvHEDbsQbhhVbccdsyNsZSdlh84uI04ZI1/3yovzc5CnNtbrRbU
pzyQK5kEHCNkXr+OypHpe3NmiU/MhKrDMPOsOn4TVsyAAPkMbh4g5dFtEbro0Q+Y
L7ge//ePMTzmUo59U4/kzSgXZ3m0xZJhGTgA5+f9lmvalw4bbPdmrMOFfFshmdtH
JW0oY+2vd6uULgtgNH/z3Do8J362na0WXZpiajtX4HWY1FysQEpUFACcSD575QO3
fuPIU1WiKvcSlGjiHVpEuOrJdIjNKuCPWxQYVILTXjx0g4jhQwLm0agho7PjFCUj
vsYwv7AOYvKPQcfmSoMN9W3xQcmzFOVaUMxfk/IaEvqVbFySSsQjzXHrtPqznzM2
2XsSlKfTq3Xdp5Zz361p2vVUYcOmwUgNVYiVVRWK9chLs4+gDySydv0GJoG9lR5k
zx7xbwV+M3bA+hyIzrZhuU82rnZ7cgJO1C+xjHHzPO2/dPkynmH1hM/ZFIhN0k0m
6Kq+iKFZ82gJfyImxpwUMyR07NwcAHevJ9qpAnk+U5OZtgRCZRdVo1m4fcxL4Vh8
Em6xC2yKhCGTSYtjBQInBlqQH5ZFkCwp0Hti+fjHjljHSLFR8uitn9in7aU48q19
8ycop56bPVPmQ3/VC5rhCeIiTw2H5ZVnP38WNmUXZ7ZJ49j8qqn3jMwwzv42aWzn
aZQQWHfJcnGxVazo+nC1PkEFBMkIfvRjgERMDWFJWexEFnH6aIZO4iMN9BnuD/VR
vJSwCG/j0HxRG9z/Ct+FRLuQ9CV0GqNi6xyjkklJOQ4MVgG4bRPw9VwWh9L90Y4v
0Gn4orjigFHznVAD3LzkOcffg+JuGtsiLXN/yQ1JwcsXFWbRjY/S76ZZgZtFq8oL
oPhTP76MVuX4wTtbpDWNufgV32URx5CnTe0yGETf0Ov9rg/sMjHPYEPFZAqkoxRr
4OpPyTsiEFL6/KkOQEf4vljdQmTep44+0saxtyKG702S2Dw0p9tWdEqSThKWZw2x
ELRTlPkBVRV1tFDeQZEg7B76WyRjVhsvzEU+i27eiHUWE19Kx6NtvLoXmKS4swIS
hf5LANJi5OH5lF/JAlpFrFmaoS4qFBJYUdADnrOLeXmO1Yi0b9I5vFp2aTs1hjd9
MLWe7nopUjsmyENjRfbARjrR4oVQ6ggLTh8YyJSWQGak8xvK4f30gerNOUna4huq
kzma6XxXtGCvhOSb4FPrhTiu1Kdzna3nwUZffA4FLrp29Sb9RCpXnSQAfbtpQ8Ey
pD/CEDTom3bkE4MekqhN2wSkb7Sv0UhQ7wgHliURHldDqb5tFBhQJennQNoYHRS+
bNmV+LFFHLLs0wqpVqqjT4DiNVwBmpND3SCmFfdMZf96VQEmAo3vnTI2LV4Ouw6s
lw1ShVsFpcTpJz5umhXuyBsA/hsJP62XO7rUcYwbtvb1YERr40IKAnkvlFm+V8jd
P7iyvJElAKs0yLSKCHE2PJaqDQ1/D9UdNxg7m53DzBfFWtwJwrG2JBN/JWVWRZK0
B7WXkIY/WaqS8mIVUgTEmTirnH/uyJNbHwhAqOLC2xEW6GZm1R2E+eKeO4du89YU
puk45Owd+sf75ce39mkReBBgx7YG6B7NLtbXg3v+/+T1OuUI/hD0gsRY78WTLOYR
aQ4fuYxlwidl17OB7L/ER1bdBYgQc08mXYx9nmV1R1nDEexcXvHG2Fw1j8VFva/P
zPcMtrRSoJ/xUqt7I1FMWvwnlIkngMpeN3Qkg750iMSgzLvvpmbRCzLyUdxE3PZE
vgcRuxW+QX/qWtSko+KtoVQtCeIJ/BlMozfQd1hFucyPlx2emxLHyEDby3pp4VAE
wfH7lgOkRSvtnGpDmAMZLOzfukSHbFPbus2/HpaUTVT+Wj2Ai4UoGfadxVRPw3nK
Ok1jP21lQD48QzC889hznyZ7kYomhB3G+Lo/JmxE4+ycK+mlmyClWK1Of/isPd6X
fR2EqjyvzDxgbA/UEWUaXTjU77yAv6nE2iEwCctzHwAdT7tET359oek2GAHQdYXy
2BjjG3kKLL4fJ4uHX/O1N80rICLCtDYu9tujpsDiucS2ZDmUfPCjN9vnsgDmjQCA
mkn7NCumMZzihdNiig9KW3xKhdmy5/5it95vj66oIrtBqCLYY79KbidAL2P72OIl
+St0FoMHwwAPekPqWaNnhk9E9O4yBgsYSo0umDOGaaplZOhOONikcZ9B8adbHcqQ
7IYquzUUdul7/7l8QHMvEndsp0sqHsxgqiIhigZzKBhkH9NfLdjtk0PFhg9csnUP
JAG9Xn45ofiHz0GzhS7eGQ3DqGKDhQoXXX1JspXRz9vplo7PDeOSECkQWTDQb/L9
prgNIGhO9dVxiBu6lhD+++Zh6sYCOxbt6bH78UZNhHw9Eylcmxnj+/VMJnw6/cmU
r7nbasNzz3CrYT4rsGyx4RqyMXAV4Bu4ehE0+pwuLCCymVmfHO+mxyvW6kwac11R
lWNn5y1oj6xVdmUdOVjnOZROZEJOuRJRZXvP9TG6bMFZMDOHgrbwXOeyALcxD2TB
su+MwWYqlAP3/yV6iOXzRaWpA5rDYshTouUyG8kJ45snRoCYz5IRc5A4SiPiOKCl
0vEWDOnHJohhvOD7W2fT0YwAUlFdC4Z8TX/8qFSYom+HAhq3rbz0+xqD4fR7CpBN
4hBXNpOCf1YbkNRO+V2sGXeLCQKItJtcgY++pOlztSQRkEKoQYgdYhUp1J6eQ1lJ
RvghUWCaI48txxFhQzf7wNOlfm9gEOJOiccFXXUdvdItxWHqJUS/WdYXgXXMe0oT
+Yqg0XC/d7aHfg1QALh+2T5aFe/6OKDCsSmL0m76XnJUrLpWaTom8v/IeX860mnf
AiPm3TfX39vImakMtfULZuO1RqAJ+xniV6HwuGNUTkFWpx8FS6c59iahh0uj0gxF
50SZWtidAp83bYxSwnO7QOk6G+ZeLJWYF+PWP9ZwMvYTLjldHMSQnYHaebRuTyLL
K1FQeox1bd08NKoZ2PoRkNiUV3OlrjCjr1WXdwz1bTlGrjUydkf81AiOhpikVUMH
TxEXO/08CSztKzfkgdtblQuYuZZ/rBIKecdutSJiZz4sncX3yOMVXnNMMc9pgXCP
vBwS+2J1fImW1GfPBu8ArA+Z3mSYjcbt2uyn1FESq/NbotkfRT1muMhaoMcVxOGO
F2fRNq+yG0kxwvaNQz4WYeab7u2p67RBJCZjYoK2c/fk5wvoKtr+wyU9xN7+2/v/
xdf3/gdcF/xaZmpUq75cRA+Hw/Nx0Frg9/bACz1SWnyzT+cLPIBkf4k7CGf++Avf
hUFvC+5WXXr7KsHsn8Xc4pY5aVKnTBaewP+QLfHGfnq8hGeEx8hf5Hb6ChvMfzK6
YoYUNhy3iHVM34ac24AK+tjRHoQA/cnSrieXi5wfNAJ6ZC0dVg9E9rSe+rqyG5N6
gv2CtaBDmaidCf5+I8evVBw9dx85On2JBbMXMko1MnkxycpQQg71kFfz3oaRCrmk
/LLcv4eoQhBGF/BBl7ekLXm9JMtLnUhNFlt7V2buTCI4HjtEIY5cSe31s+3J7GDy
lDKOzNUAWtsc8JV73bWtr30uuwggU4bHwwWhMPlNDTjbw+wjWYtqHDtT8WnG8/ky
vKM7Ht6sXqADxan5zkFhFT8uiVlaJdViXwBzaTTPF6WFKBAnT54Q5g0bqiSbgm73
7UWQ8MFmvgipIp9BZ2m908s7bViy8i2xJJ4I7TE53szZWzryStX0XojOU1yTuwO7
Ti6fPpv9ZSdHu+amoLMHsIi/svtDsupbZlLSc3QBT7Ra3rICnJ2KCdSltoCMsv9E
Z4Q8D3B2LPL3fR+pamyhnSI/QHfRM/IfWWBBUCZja5jHIkfU0RpL9tl3EPz/CII7
PkSj4W8QnF5Njz7HC4dgwZlx0abhstLMYH8cIICHYuOO+9mkqqFK27l9x/YgeV0M
lslFLfMWXYdva8hw6tzSAvs9CCZ+otQOMI0DrQxJHgQhFJV5i1DjeWTuul0Ij1Fp
QBuQNOGEtU7MwmcA90TVKNz80ENnG0jn2q7k68ycrKKL+YH+e7/kJLZ6/UPNtDna
uUzBeTsFMEvo0BKvgIZVWSFoS9e3bBMDl+vfKWust+LvbCK08CcHW0Q1i3NZBqfo
QtUGgTt0+VCSlD42bUL/+HEbgrCMqcEt0+fDFrbgzzAvKf/EOHOdXFfya5fgaIHa
LC7a4ckBk10lVXPmr+mMLwGrSdPbli6p3OCqwB8mGHEGcC7Yvqz+qcwSSKBKGrdJ
AUYLI1xoTYQw6wwl2M/y8CbHbC5W4Qf8fnDsyTh+/W0efrFqrO5tWXxF08Z+053L
TkEeBxJ7ceNOMClrPKZi7mKWO94GToYWCC67+WeOb8G6UEZkdokMW28w8KwX5dw+
hKwaEkTIyuerlrbrArgjk5HcjLaiGgfD4bQXYiiCxi0c79MJ063x85LBlI0+Q0Pu
9GVtYHShjABneWJZYQBV+5mnSxXyJ9/1ZDQ1D90XArcGYExtOI9j7j2obH+SiG6l
H5Bb1Ctt4oIFb35mznClFF5BLsjlY3T/QxDrWl/jvawznKMBYnmHnQOusnTT8/dh
2rtsAcpQgTUpXVCm7tEvSUxzSocPbwS9B/emY7/yuhePz/hZYkVXj1y8db01UD04
eWGAF08cRL8yY2ALHFh2VNNEbAMNCC9JnahPsh8/3SrpOoLWgjHa8OwkPrRPjfYT
OgzG6cD0WWq8h1enAd74+UVIk8C+/7LlwxseYsg9UGjQL6j77XcrvfCFaLddQJNP
aqeIYlc9KQyF+4ZKqVqQUleIPQW2zIPYzphRxVd4uw7P76zQOo/kHgj9Py4zz9ze
jxbG1MmjxiqLSZKzE7Y+xH0pmYxx4CD4XrEqwwviqu21xLwCrM13PvMRyhgoYdec
Rr6HueYgXdZDt6zT18zHZ1IoQxJQqaFQiQJsIT/8W4EnWgFBZRIorTKHXn5AGPm9
O04U+rnk5DFBoB/DRusQ3vNyMVCYoJEHD0PRiaW/hiq2ocgY4DGGQGCFxyOr0QMs
+cwI8c4ct7UR+UoTdl+VLYNtxMKs3rZTap/OH92/iK+F44YQo1iL/MawkNL5Pj4N
n6BQuiugXgY7ioLzqLZFfW0Fn8xPtACQsnOg9k/47IA0zNNlVqYQCMF05Rnu0nut
g4DgBnyCm3DL7VcyCnoqJpaoVQHWP+k49HPxUCmUJUczRpQ2r2PZDWxtG8CfidxP
Xkq+kozrP2CVHntsgXPfWOaqi2yNl/4S+Jh7NbN7EUUN27L3s9Snw0/JRJZyiz0n
HqXSTTAu6uGAcdEUEqfq7hTUh+Q8gG896OArpr2wiWMqyPkB/r/G6nhdMk4lgiL+
57opu/GmxMWOUarXaBvMeXVUn6NIjb0pIe4zyMBfQR7WDFnxGT1on1/mKFaF5bq5
yeRzUGcsY1MN9CW04EWIxe0dLJCB8VpShR40TMv2CxbjKby1AmB/7L7NFrrOTHRg
WA6nw9w8Z+VMq7H66sWjd6ql1Qs2X1myl8hUct4UE4mBb5e227qYdYveiI70uLN/
EDD67QFG8Ws+5hMCzlb/I+gnXoLoGJ/CF2kYqeAM5RDyPsd10ndFgAUWIjRR7uVm
PUBARYLrwiv6XgJRN1LYq6N+0kIdFrXuqJ5f6ds9AgGdKDD8LDW3JOgguJ16r4nm
QfUj1MeI3WKyAyJBWnyS9nesw4p/THGmul3Y2yjQ1G1uvEzWzx3cIlIteEpWDNym
EpQSYGXVY6vYeXMPI3H50JkxYrX1eDtK98QBD4vKNVyw/IF65zNcTS+5/+ROUaiv
+lXDMB7v170GojSSyyjaic8lX+fhEl2Uyj6HS3FSpxtDLNEXcNi1YDuBZCfGtyB4
Yf4mE3CEYi/lNgIN/PFSOtL9Vvv1BLu1WFTNg9+Eo/Fk/FY+XyqGxQGMkXpr/slg
3lbnYaTLAMEWwlrSMxBmibg4UwtrWK6/g5VYBiGBUgzB7DHQ9QeoDou9b7UKyzpc
Z6yt9PrVUqfoyi+pISwAUBYqtO+1qpEqUWacbR5Xx8WFMfbsySh/NhxldqH/y6N7
RRQ1FzUfk4ek5L/cL4Hf5N6VUuo6TJHdSUpv97aUYCeZG/Eb9qkpRA0/e6z+Tfsh
mQzBKAP6+eFKyFkq9R5xkk23Fs28aeJfNZsDAH2nmtFFpSzTUuQqatT2fzokp9++
OjfW9Ieu+yRH3IMhy5scHaLhn89M8Wj12FxGaJTjnrm+1XB8wVcyoiPVgUz0sBR4
ErODueY/93j3jnL3xkuVvnJOTjo+RBjXxp8rc6XcR0uLKNmLqT30kxub8Kqu8Mmh
uAjPvDUjsEYvmt2HFI7SouFEIU6N0HScxfs+docxVUnKhCjK6F/RWys4eCmBb4PN
HMH8j3o1SVdr0N6gM3Br93vDX5Tm68Bl/T3eMk6aCo0YDXZ1PtLlQ+cVE8tz36wY
PvMxIgOlQlD8/0/Ov/Ld3oz29W3FG7jhQ69Vb0bdSdVhihK9AaHFyKQ1mKzMw5OG
Mk8Q5pUGfi81HrEo2Mjmb8bfAxSOKGpm6lnZ3Uc5U14PUKGXkUFYNTylZbDESM0g
g4YoKhO+rX+MMOx4D3rYs4JonAu/Q2vEHjPJEeTb/H60wKVG7q+RGxo3pkjObuZh
Go1N9/F9E/0gVlCX3emejS3SeefdVeZ0R1LoVauS0cgBBbkUiWrGFHV0+DC2oHGa
6WP9JuYUowwqIKit/KxVPaY/EbWEOFTVFCKDS4ngtaqDdfThTPYSLaCvspkPtEML
fjzsA77NlHgqR+5bgGapgQ0z53cQ+fh0LPMWAdGtS9J3IlwjffhiNa5UXGKm/Mne
uAzwXJD0vahgtNkBwOzdMMBtO+186O+lK4liWULwuch8i/xvy6yk9uAATeTqjfcb
5DBAKBFSN23vhmuCkB5jLmeW/9k6zZjNUp4b9QQzzpPdm8jAVVM1WPxRw71ycXGn
egFjuQE0XKrG6QDuuiSRTsrJq1DhDRECCm5muY2tvqKLpi2ZaxB6DGup9JQP1jPw
D+j+c7Q2K8GCv31NAgQdELQ/XXgcReX/OPr/VRvnHWoIgTfgJSHqqZ00uGbi6MlJ
PrpGnMWtqbRCpyy2iTtJJZjl3Gh88AddIdy4AQKmYf8xvL182AbzofOk3JmN0UN9
95fotY28L8TnvRzU9KKAiL7l55qcJ+rNjJo2ovlsbJJ5D+WCEd7PmC822lowtum1
WAtee7e6+z+uVH5ts+ynmB4xkBK1JrB7B5a+e2sA2dIi5b21Q3+g58ZY2v/VSv+q
43pKCJN1/CMt90B9445qC6lydm8rZLtN2bL+q+nloMGvFc9p5PHYljY9PmSu9DNx
gmaTEpu8LLjSlgGV2GHksi7oyrj/XTQ4F6Yqd9YpefStcGOePL4IH/DQL0UYI9Ra
+1mcld5Y45yxPtVEbrOhrR86o5Q65D9D8JqTrlqWe6iO+8DIU8ZSZMolzpH2LKzj
1Ga6/I8ZPVmpNi+Enu/IgzasSLNMxMKVZkXIb+vUPaiEFTJG4q/4qWNFXX+UCpWj
T3zI47pTiEJoukM0z+r7Bc6c7jiB6f/34w6WqCq0YODApQGzBgncm0RYuPJasWQI
4vUtjkTpx5MnpxK7bHlJvbq2/L0i6aTaaSLLuoIsCQ3q02kff1+2f8EwzUUXGNu0
jd5/2nIhauw08fl2Ctz32kCaZwmePSz3lVbl7D6gz/Oku3BdXtfsV6AVF+ALfcLn
Y+VwRyps6oHdFOytB/kYs3Bds1w8vyxfdj8JBqklsnPoy4NsMSjxPAid2fYq8Vvh
eZ6ZNexfLl3EB/lcBMjRLJxlg6eiGzfyJrbWYRbYaSOfoCwneDSFGPHdTSfuzchS
nqhILXw3GccFZHpYSZe05PtEieHpNZVcB7jG5KSwOEmpAIQfGO27+7bLCCtFEH1r
WXE/IYKFVYBc6iGjBhLfDwZ86T9MVg+aGak+uN9IxUb4ExBvLNO8+vJMiu5Ty7K0
j8SPC33AavgAW5mWtBhmNh5qz3w824xdZlxme6yK6TeczwOQ6zHqtXo9OJNZ9Q9U
HE5ipiQ03pa3S0YPCf8a3/K2FKfeOM0e3XwPhR4n4UAXj8IkjA0rct4DONArhm2Q
Q6QtkvdBKP+iWKtRgjPWIG7XKHrT5vUIf+sxR4Ufnnt3szVnzbbIWqHkxCO0hfb8
pUS4fzqVqp3HHrPjHGz04o6uZ5rLr1yj0pRq7cFKsctOGChJ2XfqyXjsoYFrH1WR
MC39NfcVXpl4n7r3i45rQfGgyBa1NR01C7+Zs09brGAurlbKk6HrxQrvmNfBlki2
IdgZ8LS0ULYwT+NTX6X5A68lHgteSJr27INzVPc/zzNn/uQA/wQ3WZrAr10vl6VU
1Hid5v7Gc5Sw/3XI2SqAkQWDeQgWs6t7tXH8AmbcBQQmOhfq8eKlYKhVxIqXOBIF
7q13kkBFMmoi17huTLpMPruSV5mVWk1+MoXI5OhxC04UZXo9ANIw3Di376legSdu
p+oKc9jnGHlHZYud3GM7Cv6xlml9E9bc0GiqGjjfILRHo2zs8ks5bNzoZ8DbQ7Cg
4zLdbdkblvst8vfQMa4j1LsWMYq6E+JhZJ4LQggCcxTUZNcDGNzxnNiSkOo00q89
+FE5ZRwRy9kJfRru0ciz63vKs1OTOwq850OognAp/utYC4LxzrAQnHJtkUYwwg9z
7UC3AbT6dniE7puIJBBtgJON0BnJx7pGa+SrTqhp0jayhMbVAD7Ln5duzkiBKIYb
nQ36PF0nxDXYcwO9rKLXTF+Rt3QdKB2fbEe9/Sw5Bwu66W/oD/1OvEAMcdyy8ImQ
ZtudX2I1fVPBeY8FMyAmkN0NaHwxmMBH+mtF6sAG2r4/ju+mcpKP/bUBCZdePmKH
CP+a/5NxvhDRvEsh/zvz3nQTnONzCP14IjIabUjvpKOcPuhvpZwySiZtt+jJUWlr
IHgGEDBvhlBbfXOUi93GBTqfDmv2y6fQ5+GYS7UdOC+bbf+9b6qMRHs/dFeMVG+8
0sPP9Bea4P5Ss9cl1BI2RiGqvwdwV+Nh4LluQdXFv3YS8XwXefjkD2PskhGuUByJ
wSQ0DvOU7aRY0fmFpZcWWZq3LxXNaKLkDl3c8PnaS2/CkI05fvZ0a8OQlUKuVTRB
F5VxQ+LCSjVyV5VJIeqZorTcDi1/X0UrtXYKitLHTXtFVP3qYxaYEiqHp49MD4Vw
RMV/sbgQnkWAgEPnqnD8wmPPRYlopwg6tR1RcfepjUaQBokJea8sWUTMbUp/z8vh
RDAO3GJPmUTlg0GXz7H81mOfqrDI5WM5/mpcQilXtK591Dk1r37/QnYmCcEPvpOo
/lzLBL1RF+R9MOVIkvKDdXHQpdrdL10uXQ5fboK3eHxqrwvgKs2Sq3VZJibPPvdP
KmJxgKeiuWqNRUpQhtP1hKU2fxYuXn0N9UNIakS+dCdTBNh+9mIxSoW+P9Bt2BaL
6MO9eEnPj5VeKYHgwLShFaewBebPLtPXa/QZ1E61SNV204qQol9l53RCAfAA9hX+
od6c0kZdEre85K82u7UDusVal9ON/2lJgEtfuNvE6a0EBWvjmnJbHkpt7NrmvEBQ
NPMns++bay+i2aWf1DuS4DGF9D7sFBjbFfSZnBeJel5Lr/gSDmgPLrXwZY06Owc5
aCBIDSjB72vjL3LTqCxkYpyzo4oY9X+w1kihoDxWQGxKwIgW4U+6dROTRa45KQqm
5IKLcYxWyIPxkASBNBrffnSX4FOvTvVSXf32hkcAvPtTLLfItd0qgbSwckO02FCh
W4qKu8FoxK73HRpQN6ooq/wWOTEg9jWRM4/0gwlKuCpLsmZ/llkTqm2NKDt4YUy7
7R/DTD9iAskXuaujm6jZNsZ8vgiK6s1fKvCT7EDEQqv/VteaLMWX0gfWAbE9ahSL
QzCZsQmiWNAi7Wy2LqVPkMbU08tyi16K1p3scBW/sK8CU/A37TdNe4jjpXGSjiOw
kv7cyMuwuhzqdkglLGbN8lv3bDwtxvpAOtMdFmGD6aU5de/KqjWYd+UT6/wyx2+6
x9kGC+ub5XGQlURIqq8OIoeZo5N0sA1oxB42r9utyF4UsbBMpLTjSrD0tkOdc0IM
JQlDrVkT2iD+yroY3vltylEwxUJGcKDwBVb4cco4oUscb39+5R833R/3E3tIXEOt
GS6ZvehXwi0I02onJ9fayN5z3LsV+VeWXEECS4lCh+Gs19fINqYjn+32kSXKZ80h
HPMVEAoWDNk27zQxlJZxBnzonyi8oclsqnnRL7A63nw7XrZftN1HLD3PEhXOGyTy
LSXeCtLxYLPtqedsTCn1B3z6UHEb6HNv8v+UYleXYnK1fJjOh6lAqC5LUP5o0J3n
F+a76h27VYY+dJD2Tp9vg+tTobUUexfzFlR48u6hGEWRQYaI23smsx45ysvX5vds
q9SSYVSVFIuegftAeXhcySVbx3wAZUvebtdwcI1HbD8JObc+7f3oCveRXLqvBH7E
MSCjqNOHuSKfvPIw764590HXHEcroIUiJ9fxFToXZEr034hiZNB5xuJWB6+0RJU7
fc+P7NyskuvIE72HGgC9HCsqTtw5Byr+tCQTNZIIeTSG/TSWa38ywxMbs0JMAZjC
PMbvQN882oUCRb/x6gD6dIHMLmrV5cQBUeziPZnePwJftnnIbs8C3x9QBxt3Lv6V
f2YQk8VwO7r4WwU6ndjXZTeSCB5VAWlGlfClLuvGJfwLRA8w02FKQGOFp6ngKVEY
bmhA4lDYabXjkWPdc0R09Nei8MfbEoBYL4IXwkuAy7V2igAqH5XdHtRJqRtOU99K
1G1kU7vFOAoeO+JbCqaSgZHYCQzg6+bjEuFhvoLPwdW3Xzy8IAab0rjWEEZdqPcO
SsWrWXmXS9+ichjPQqhGYjgnuA8UCX3yeLeOPTGDsjXkSCmYz3c5TqINC2a4I5J6
dbzTtahosku3JVyVZEXr/Lw7XrUwgzkPitSKy7/dySL0RZKyvKoAjnnUmZiYHUNP
QtCKb5Z/+7Gwf2na7lbLfGHo0daVYZtVKiPOVijqbKtLs7uXasIHGHHLZfDUVzhF
Me1U59AnniIqvpruMyBWccba+L3gl/smGlkqkgCTAgq8qs9uI9MKmmg8hRug0GlY
uYQjxvePGz6ktpA7bkvUwgLm+GCjt0/mpVlXsGY9g5vSm/9gYzHl7o75EkHmS+n+
kwr0IXMPbrkW2qXnGpkK9tzBidr18zXEg7ycxQnKAdggj3DbBY5hXZnXn5BlL/dA
y6JJXjcMjh7AUAoB/LzohfC4n8ja260nCI/0h/P+KI/WCGV75sL7GkQJXyWxWYie
Se6HDgOf71G92Eo3yMSNuBy3S+qVu1due4QcwkL6bVfVVJHuSh+zKwtjPUfKSB2M
gjRWGKqXkrM1vAD5c1UWel3bfVI6hJ/KbcUwGL4KetspbiAn/xklKONl7sz6is9w
da1wvm8gdel2mzIYyJNmUCT4iiA7wUpvn9KifuK8MBWJdZ6tpxWhPWt9CprTNAbZ
rwm8UgJlo9HGJDTchCaYxPpOamdzzYoHmvicJ5oXguIdtFVIhOA9C2/y290sRttu
ZReadh026YRwFuhZ8iYE6WK5yZ/7GSSYHY104q0vRbn9sztNSWQmxzYiNohgyjyE
TbWxNi/o9qst0++gHVt798gCGA/IPqRJaOpWmSIEwTBihJZUyVOUpo8Syx5w75QC
Krhq4eIW+Ry6BbUdw1z8b4jax/F+z+yWQcDZa+k9brmw6Mwgs/acxlAP/oA2jTpS
6K6oXFshJIY/FqfhZuCVeCjFyhOVCw/9CEAPXCspAzuRz6lKa3sM50GiNkz/V2O1
BkXJjVm862hEIVish89EEVmZOv23zh0DbQxZxNEaXpnT4Gh13G48+wAQ0VgIS27F
ar3KoTD2QtIiM6MtqTl+eZV+bIit1AyuIDEDNzyxOT6vOxia+0bRL47AITZTkjtc
6re9FaGDA4TYlajAkugdbAmh25mu2h+tNBztcl579eg1AXPTPisHTHTHWEX0OkeW
XAa+UgkkccVYa3Mz5M4Khsoau7oMESWjFLMaxxITDkfx2ByWNOhCtCHIvqUX1DK/
+gPZxTkAUSGjrMjVtUw01KWMPu0sqaysfBpC2pId3jyjAqIiJiAzfRyHePOQZFu7
lfvdU3xAAQ/sMpzf4ANMVABCxBBfbV+0UPjXT0obyQ4f2HvQtSCdQA0dJyuyz3jA
rUuh3ijvIEgh7tRy96F2mV58/Or1hy6A2E+FdSpr54DMpyV1SFv6dS8AlbJ0xnPU
bkxD2Vl9cWvL6H2XtNFXpBulYAhAoj+pSQKh+FLaT+2U0rCSoFIYCTg2Sp8GX8Rp
wFNAXR/2I3foW2GGd6Nej2C1+Zdffg4NskxdOj86ZjWKAoTSSCCYEUeYRQSrTgxY
ROPJcLIGa+lk5TJkpsurTYgsrgOUQbdyaEqN9OligJ8O8i6JfBVrf9PkNNRQk/KV
mStOlM2Db7jURDRu4neaJpWY7hSwmhidrNYdJsw89atPpAxK/7Ssf5whe2oFDTJt
KM43z/uo8Is6KTpexoYEJ0L7NB3Wdmkpl591SwYIqTIThGXca2AW60rR10tFbPRf
dRq0IOefOVMqf+tZRWBBppLpwndrJZ+7+vP/qJcaC1NbAZJ/XMWw9MYkKYgDEvd8
SHPNTzNNZ9fqurbtPxAlTqi0jPvXWnCocipad3jDid0KPzQF+ov8lHEcy5hp7N9V
y73f8pcPt1aFD8gd2TO9z1iXI29oRDxug3X5CjKABvwxr2G5AToLg07RYeNqioXe
NRK+CUWI6iXaNSKWtMlZqpVLTAig2miFogzw4f+K5C3S5u86XPqFzOFF/ybgTcVY
xk2YM1ENQWOrKj5UW0dgd4ePdoV1HjKW60BeulrFSdfuVJcJUL4z1ScjQHwFPIY+
5SpU3MXlQxfe78RFt/MRM8xTl0vYw0+MAgB6qM2/B81cx0Mq8JpoX2uPjdFGn0K3
ubgR/NVXcNFNByS3KmwjrT8pnxdzojqSy5N5qZxmSvDibbEBOKZsbpL/Ex9MtYC8
HYdHDUSj8Ifp+QUPvQnLHpAvdtwRHeEJnr16Sy670SVCzg/QxNJtdMdLqGUqWRK5
spCVbt37wfPBIEBmeJRHqYklGAyWSgFAbSgLHevtR5IzfCmMynNp1q8m0Dej3TdY
CYgLFvOoR017uhBOUZri4fuNjs+ul284adwNdX0+9/ngjU3fmIDlcZJDbFmZzaMl
3NGxoNhuEYZPll0tkI+ZBQgx46hTYrE001K2zowpBxXpQ1RHf1co4gz5cPsB9XVG
DITLq3GiuMvEYU/zpv3yg7fWq0HzElsD49T4koinmf2inBPZHPuzjzsvpyX3BOlT
vBjBoPr3HPuLXjhfuGaOt8Njn8TWO0gar1WXfb+MbDR+mm33qNCgJ22cauE+i4T1
quGnMBcml53TGih6wsGoG5Y06is6AHokbI/oV6ZSJNHlekr7Eat4+kGOfv+zD4tH
DTzcpTWggyPvI/91NC1eFz1XXnuwg1VhiF4z8litpJdRb8kSlJlXks3z109Cnmki
f6WMtu817con3VGwOjRYA56tT38Pn12QywiLsIxHmq7e0k7G+DALzWSOmtnKdNbZ
Xq9NRiFLV6yqaHXeftPBsnD9xSwghW2u/NCBs4usNML670KQZrHT2rMhmQciiJj5
w0XmGkpL8s/hCZIYhm0Pf/0cjSGbZIQIUNjwWRuMAKAIcADINKluNa71meJU96zW
BVoNEQBNLYTBOQyO5hh+UmqJQIBFQXNjBA/4e5UjD9u5iahsmwb8M3tTF2SsoQ8q
gY8/zeuWb3gmYpM+P8UDdzWYRwJKrnBuxO07HN5RocER9uUPVx1Km9Hn69Qfq2OU
ufdRcbHP/m3FwxiAU4n1jlx/DcgSp1c9VOpcs7VtD4vwYSV16EWu2QmGC851+I/m
PVnoxBZO1WBGQMHkNDR93F10SWwuNt8UQRc/ut4pALXGGmeee6RFFwF2zd7IpRoP
APu+0O7xTlnmkSreSMZ2oaCxf4itcxWjN8OyoF9EwENte7OCyR3aqCSJP4PRkJCU
oypPo/e7X1w6LhXb+pdKY35YY8vhsuL98HMFOOr1Mqo6zDPtjiTzWiP3MzChklLJ
r06Duxqr742I+yyJTHmMuWnRrkFBCvdX5A2kxySZkkX6fpY8bsz6DJsHy6swho4G
sJT68NMcBYmBm+0wtXBYDPu9Hs7R24Rl5BsAdfn7YoaMKiCkZU2G7YJDCmgzX5Hn
PAJzJsbigHIrhe7ii/1Ir1L0dbeShDjXoZqJUR7WTr8ILtX9NI+y7HNEhpM5hIl8
HNhuriOdDrIBcrVru9NfkoLEXKWEcGvMj35Rb9IqsAMppyJRKYDS0sigq8iGUEoS
1acKg1HaGs6VrKJfwcY04wfXeK3LEndEfDe4T6KOVIjmNo8/KyhiAyPBVXOxsNzT
uufllOOCdd+5toWQBpzu3wb4Si5k2K4QDp/nOtobN7ZgtwdOUxTjO8z1VdOEgx4y
0HO2FAzqQMlDniv6NLCi5B9W4aycAytVwdGgEVBRfiD1gpZdvoQC0fv19JEgNpiB
DnFdE9OSje6C5/Ld2THFhxh/rDegAJZtdMxJtrLNvo8/6Az6GzZE8/uzdTnZpByJ
Wfd6NM0+Zrs2iihTmNIGjmAOyYOxb60+aX/psSLy6KMD1G+geK1mMaAkuAaG6gMD
vZ0v8r1kY2tfpqo5n46XMnSeK9IHKeZIEoD1C5rhvY9mNP0h9DgNLKGGk0ENJjAB
rFVDlx3oT4kgSU5IdApuOIbGT6AzC7QYC2EWkfLZd0hBDPZ1o5bXkD22taYsp5A9
Q2DXYc4wGmTZayKE7zbRYxaTPnS3yfjCvAic39iF53NyWyQzMbx+rLbZrvTwnCXh
H88OhFzsegdwjulY23xxD+RnADKGuDQ4wKXXVcfbkfg9bP0nPA3TnCdp8AE/l0bO
09dJL+Rlz/eLvTZJh6A2MEBtI/HGucIC2wj51Q9CcGkng5PsGAs3DvxhylS3uh0Y
VgWlFreNDuPERgYuZkM2PppqOMrRDXiGPNUhKYApGODDCim/RiJfcKSKUkh+niHl
QMPa5SkwlDGaCh4hr87uecr/3UmjzynLu3sITKzxG64er1Uipz2yE540cZxZPiwg
zNKsWomGMvhFA4lMU5Xwhy+29LKVfMRNH/ua+chIDw2NXjKIasw+IBqYsyR70+jh
6DMKYsnAvSq4i6iYCep1aevFMEpWXeZp9jQlJ7xrrStTQixAel91+U5XwXLf7ES4
ERohspXz1+BQQa9ebMhaNaevHdxiuIbW1kfAHFcb+Yq/VPquv5LYMMkAIYMbFmir
lee3ySKM4BJXdGU6KZroKZ7n7E25EbWDejzZ4393/3FqnIKlRVM+saqdY80nkGFM
F65AcqtxmUqPe3sDgLBtVa/2Vk/gFNnl7XOip6sp5UPfHwcK2tYMg5J6+IGyR2dm
cg4lwJpbqpNHdnVh6Pysv5qKbju3upOEoEI11nt2xU8iHPLXAfC90lUyxOY4dm9e
go0uoZ27K5JvlCDz9GdRa64ud8AS1vClDFZvKZzCFXbU4qyq6RzzYOfGf6c596L4
uWwjjgU9MbQvO6ryGKVPLbT6ldD9wtSD2C3lx1sr9c1B44p/aCLqJMdTuICCQ3Te
OXUND7l6qxkas0/znZxF0nKu5txFkspPus7kxIXD3Tcw0ajJc6+gQKM6BPL7M0Vx
DBHzH3ckxIvWfwPLIzvPuBD0xKyBs2DTbTYj/AEhKUgJPrlXIXvEveId8OZbRYUz
pFHETZ/OmZr2UR1WfDQS/Y6P+blazO9r0bzYiihnf1NVB04Zbk6XjD3Ext+O25j6
3E//gTkhyJjxRMtwALvcxlDZzhIgPg5dAt20y9USR8weE7cltwt1LiD/u+0PFKaH
bWf02ljfPjUepdCWL803I3PDrVVgL4a8mZeu4WMhxLPJh2U6nPm/IFb6TuT+KgEi
0Sw6bt7Syyh6RiWIbu2LUjpX5dqbmwy7ng0tkhDTt4PFnNCRsm9vJgipkqIYTyCE
f9iPbdxqbKM6/qQRpS4Gq/+J5HFWsGYZfZXavMfCuET6iH65WH8gnHrHDzs84SFq
cNAC+gFwRM1ToTCk/Oafifcx7vRTxzyptV+mSZDeIXai0X2OK6YJjSiAL60CYKBi
Sws5BM+R+Qgvb5/LTMt3SszAYUNpBOofg3DdXtGmKX+MngrmhitLf5Ej+UvWeKIm
qxnrchnDinwLtmEWEIG9K1AmytD5JZFxjoKHlOr0Te/LIp03ZcByqhCAz7wCLGOw
AzoXv5WKIy4fIp/+8+SYYnIkf5QE82kMapH8b5LDGlUF4aB5elg5uH5sDbYjVsFi
+q4w1SojGsj+dgxtUEzPYDAUoff7xNwr4l7A9l7FBdPbihh4VM2lgCHwva15bL6p
ZZZggnc2+p/UGV3TzIEAQbpy4Vi5ThiCkTjSYTUNmpsyYclOg3x9vMq+Qo2MGQaa
zJQvYQ69zVYDL0kzmZX2Oe+oFE1QVOY6OyggjsRIYcMwdSYrwTZtpGcn4eVDYmbL
kzqpdvbAZKusgsvAN5bvSmgbzAYVusztnD0VNYgwNiQQedbrBDU38pljHXHg1+q6
Pn1j+49Lb6LK538HmvEkvqrdJEeImZrbupoPyqkNOav5SoLd8OkOa7w5VApZrQlC
EX8p6b83GhWiMT5nUmJva0KfZCmUtsPgPhLaInlJXRWZx6Wn7/ElC5MwgMdbNByL
XqxmmTuw0tLXrQCMSNONkgP9juJbL/pVuhhjy4K3Or9jGoaAA2MYwF+n7nxt994f
+jdUPitQFEUZkQJQAbK/HGlle5LMd0JxIyHWoodblhSdWDAVOpwef9zXpvLFE6ph
6DjTAhPrbGSBUp5DxTrI0t5OWvUtPEkW6LF8XzuhqUPEC6ACHbt4sNGTKghw9tdN
AlDkMvkMrjoSl2igE3f8ZtmivYEn2H6OCDACUHHzwL6FyWf8++dCEVntsOuGMlE/
grN5vvFo3SSMf3LFaKeshWTz8hGYHWda1TM7pS8urNCp9VlgVhcuw7EX6r9D2p7O
epdREqrpjAPRwg5yW0A0lZX0sQtNEvyCoHW9/vGgTi6RQquwG9TDjJw/v1GtViVi
/r8rVH8yYUjMGERaIkRAP90XwlzAeRq6XLt1ujvIIJx1gEuu97Jnv6lAO86/3qOx
67KTd6ZeFiNR8CMIgYWafdnBlAvCR46kuii8fcyLAwXNKr4c8+cPSpwxO1yi3ln6
IkH88mWroz7/w4QW7G3prXOsFXaC5FpeoHSztiP2za3wKwHUf9vE/q3ysIUHOj6j
/pZixjq9NeDm5cJW5LEqsGCQJnpyUNrChdPzWUhjee+B5xMuus6g2ZVytSeAQPf2
P2fuwpo41tFWCq8vInz7S1jA8XEsGttZk9RLExgvxzJuEpO3NyENrpbsQuM8eoy3
47MzxPqswtAUouX1ry52kC78MlsJ6TLYBVwf65aLOMNSVGguCXy2uFh8JIT17oYb
OFyLjE1VhA5JI3ZljrlttvIlqJ2GPYrxUvaLO4V63/nm/oyCmnyM9wXByB1i5lQW
kPNw5zLDSLPArYRAZgyb8d+YW1Nr1K8YVwGAlYydU0sWhamh8GhwyPpLG/cK9F0/
SSfeQaN+qrBXsNXJYMb7mqQiAka0Qqc/VhdnfR4sWV76jAXtg6IKWvS5uw4uJg/Z
OSrsXlURPfxDdihyrS9iTr/t4OfMly2S+M9Mv1Xmg329aODiNduJyKgvmm8ucBwa
xl3svkfBjvB3YzlRJSBDZZbIjvBxX9k8gFmX3uFocBaBYgVYyM3LN0kPdfOQMFo4
83qhxv51OwyA2OukqbSenR3k6OI+z9LT/52ypfxHAzMU8smd5kr+AINSNHyTpNLu
s1MTQkQl0b3LKheDCooj2AyxeCl9g0JHE04YmevUqkBJB6PlpcA3I3eKH8vctI0l
iwpwkFuPOkjnO8OlZ5akwPqUKFB4mhHlBSvtLh274gQg38c9YZHQZXFUB887bC3Z
dDsGGMLcbH6Cp0JJ3TbZOg7ONDBcMnXHgzNbElvuSxrZvt0p7+c7T8Ne0V4S2/IR
Nkt+fzymAhb7u+4vRRhaz1ZghLcp9XCO0LRhs44ydWzxylz5oM9JxgCHaIJFjh7l
x3iPEHSpgi4LvEN6AC7T1bMGd7YuNfmIOR+CT6W6wHZp0j1fn3q6fZI4n+QiEZlp
J1zy7roaoszhY3HDF54B0ll99h1pKndRrVoti1/VqOWwsi26DnOH9lch+2aVPuNy
tDLqG2iqBY6P5+lrp3D6FipVaXlavYKdlQCBIzlNBa+49B+3TlS+Z1Y7tlKj5cqk
78PmTA9Cn82KIN6puKxiq1teYYDuhmMwjXcv+qTcl+tosMEVFpbaTLfZO4hMqRch
qrWa0MHs/gq/9xtjPyALZ8Xky6/K7oNFp2lQLVqB0ktUtcrBnl9hCPlfAl3HGMeH
CtLny5BfzKa2r2hFxvbVG8io6+GEuGM+JGVDtTMd0r2437cjJb2jY6uMEfN6WHoW
V0blRp5kw66y6BMlMhowE/XcX0w3t2nDFNbT67prhxGlqc1TPcwLurETy8sgyzyp
1UMrmDpVgrS6MNjzcvYCWm++3MQ34YfkGpj2hICmMZssUDKnpgXwR04rIlH2xHM7
Ky7E2vPYHnFuLEIO/mr3fDfdF44RwDxUNh9QpcMcCRrgjV3heSFS7QCH3xOr1e91
jA1yHoIsf8o61HMdu0gVnWkY/TLEC+S5xYIRpSYo/O/GgZayViG7Aw5VOzypo73n
/qAjpvqhZFEbJstogh0etfmOLsJKzrUklmMqJz8o5VCnl7G2wjJUcOzqICOvOA1C
t2NXokRd5hd6KAipYSzlpjcLK38zUEulafbi+HuqQAlNBHTH3xKMnTC4YnlNiJA0
29DnKc9/kDTYVnFzUNtCO9m0bjXKpT9FaYaYS8se9C6QGcwaaC874Q0aEoUmpcS6
sL961dukk7S8HYuWNYnQh0OCkqGhsYMOdCctR/rMSYA/8o0LZAQqfz+XnqwLDdVM
wL9j/T0ePnP9VEeGlhfVWZ18rwvPMUn6zd1R2aGCmo864rK0f+r0a2Eb/kC38EWS
VAx4IKmVnCeJh/kITMd9UP7nf5sN/3oxrNDH/L8EJm+NYEu+v6FIXkZasrsfAdKj
y2Dm8qTeGs/xkrIpdc5vmuBxVdvzhfMGCi08fJP+p+fJ70jcXuJW/+CbsSQgm/Ve
k50dawaLXKr+4ZoqqZJ/hNotUHxev6jO0mz5LYkyY3Ji993dpO/lh9MM3PZfRfcw
IUgyJSONEMT1V1c7gU/2TGw1vC/rNMWUywndEkAx2QiDkNFCZrgnrh0IjeZUhJ9A
CLEu8m17bQGJP1gbuZfPtH5sEhqKx6J+9FNx8wGjbhrbrlxxBhwxikNXV9FntHMv
HJYilsEjekNGDSiCVyevk5tbYcI3Fr9WbukNOxKNMzJIZxj5VEm+/fh781DYoo9G
IQdopKTEd6k5wuGjhxLX4EE0gr9bwAYqSlVlEe2/OmIcEvRht4BiCXA1aHUfs4Il
Ql1maceccEeOFSM7WdS0HM3RkNhfFCSokgvF+zISnzevtCrkM4WUTPxh6D2/a4d7
V/W0X8NuOmGwEs6ilgdrnkb6+dtr6bAdS+NHe/bxBIjJ/8vwPuqj6tbCyCpB/LJj
xYoVccY0Dqa+xGG4rHwahXRyMTBnFbvYrfRWAeoGNbVgHoiCQVLWHP3IEXV5EMlm
RoHTUp9xRQpZrG1zcEeDW78lzABfVx7TnX19eB4hNsx9Lkjpfv6BXO0UV8tib177
OoKAak+TVNM3GqPruBjEdWuuSPPuAs1lDojhNE/3rTFQsHmOJaUvmbAXsnz0OfJU
+WZGy/bGDTUboX9IpVBgC+CzK8Z6l+S+XGscScV54oUcD5kcHve7lUfqCbUUmhDw
rS/xO/s7DFbxBO7gpZlXIKoHvxJotW4fUO2ybkjMx4MA7A9d8/OPbhmlRy0svvQI
bokk8zIsiQSYuWqLUOO6T9XCVRHPg1vmqYnnUG1T3o2lq/H5b97IPqkLnYKNbR0n
OAuI5feNU2WilsIcNCnWJRQOGXges/n/x8T07mwMLZGnx4x7uMlAFIDOWFsPyGI1
bZjcVyZv6Wq2z/nF8yIRGhUR+DqxXy0Djn5nl2Y5WLQv2eLGysUjZg8usvdMSSAA
FWI+/kbSow4StyBKOn7AxG3Rx1x2WTGJGjrlPf/0C5MCj+CbTv6FP0j2uCd/tl/6
PncVwzjpLre9CWAjsiuPcjX91Gy8x0LYkrYEo3sPD3a6OpXIeBgSQcjs1shpWg4Q
pHrHffT4L1t/G4WyZAXs4jkQqa3eWAG97XA8Gu1a1jufZPviStkXV3ZT1mebdPpe
v7UIZz+nIblwL/T87FhwUjrE20kISCPSCNyl4xMfRumN3hHzwv0RpE/BEYZo6LMo
AouVruDBmwz3cs3rRN//SVQZLBYemIR+o6t8fhq+2Nh6EbeOva+KE82cKD9uIFm0
siFk2FTti+THYFLBx+KK4Ti2q6y5WAdkqMLL0JKv7iMKDTJn3DtpJl4TvUx1LYY4
GA7ffD9CIaP6XcDjSIX/hQe37bhBddX+UVlVwqJq3Xrdb/iGUZNxC8kjQ/cVd4sJ
B2Cm3OWqPwmsDTVyVWH3eV0IMj283F2R+BTQ9hbE3WyeclG/peAHzCj9cpRB226l
xvRrWFRL83qGiyd6sk2nhANqf5mWZQZKDvtPOJwURKXv8nzzZ53ZkxL4GcrhsJax
9fbjKxEEo+g0/Qne8iDK4d7eFE0OeWECqy0BjhEAv3V2nnK8deSYSC14J0f4j3Y+
dxxQWXmtGAogKHODQWXx7WomMkr1U9tdcbn4ZOLQMtzaSmMotJTRy4N1Se7yfi5L
kE0HAS70r5fjzJVGP7LivHQnTh+tM2/PbYDhAY195yv5QhrzhepPoiHwSS7Sjzf+
d9UaPsDFeMX/XOqXg4NadgBRvr6OcHmJ+AokjrROl9S8kGIQjYsGnEH2UGsgKrhi
bC55UTQ4aGAqPBZyqvxrUejFJPCjmq8B+rgQHteQwX4Tnu/zVAz7p7v3f5c5LuyT
3K278Tvk5+u5wERW9u8iyrgA5T8acAQuHHmTSsblo5iBQcRSrahQ3abiUfk4BI9f
D/YrBtGFzsYl3ENoQGBXrGYWE/lOdunGONXoXI5Ow23mMwYW/02GUHoA166S+vt5
g4eoT/ZONQ7t2s/hKLnM3k/T0+JAkWT4Dr4pnFw7urri3AKLSQRrWa+FL46OIcoC
7aPJbXFxn5pjBbrgTnzUlY5/1rJwdqHkac+kcnTABrx59KSVxopG3NLE4ivG+iST
ggzUO5/jB1Ksgp80t0btLhyOBc0l0MOcgzGDTWp4Cam/itNBahJzboXrrQ01D+ZT
0x47DDaRyCZaI6sVtDsD46OK/uoB/n+3HPiasQoAfl2IWwICM0fXrDT4MwzCpin1
wi3LslfF5hrq0nBv3MBV/mFrUuUvmkeOPnIBUFmXAE8BsTYvf1dj0T+KI1TogdMy
y6j0DsSckey11iVB7YzDTDBXz2hnzhkLzQAFIRzdrqaq4cuaA1odFUCbpHCpGpHW
r8lDidxByILRHNdFUURMYoLP3J+eSyAKIiROap186P9vo7yas2Yu21CNtzuw6yA7
llHn+d+nLu64O1n9I3gDbKQNwENSOlHqwuMAGBFmACW/DK5EHyZ9q/Rdo1OjpDyz
JZQa/n1FVJWas/Q5RBBAEii7IyzMGcD3lL4D2Sj/9drRJmvZb4GLaaexIV/4bdcW
KWiyx3ym5XkJWUaxeAb1AbTjTmrjEY90Uw7nqMGJiptaIet5ZeYc4Ye0zN7YYfkW
ZBRRjen2ZW/NOF78HSYTtuIaCBrqKRkeGTYgModSqEFjWhxWdnt1w2NLxetTW2n9
C5zeumyOIevybWb4xFOuWEGvVFs52sfPb4ZYH35SbkIvKqIEiE8RsaDhLLNpQTc3
9VNiWhrcPFa2aa+MjmHUrF0SUFB33ThCPNxWKWEfqk7kE3rfCGcWYevBpgeUdu5Q
kS2lo0kpRhf4KyUd8lAZUIWELiR3fYRRYvDknDLrvd55F68QKDEWXE306uo8v7Jq
5jIu/0AcqoU5VSsy4CT1H4b8rA1Ptzupb8wBdaMaru3p+DnXv68LBb7rwaPjws30
pRz7eqlCtlJNEhYJjq5/Ak8c55kpzbZV3UTrCQma34CNYaZXjTapj5MjEIYuNpNI
vYk3XYbV2HTJWmPM2pW89+bUkj8TH+2G0tkx3xvIAr2GYBDsYfxPVbFHuLAQ7hAt
r0/fQ5JuU1owDU6TrrnJpHPYra7q4SMJY3pnrMBcHAENV6JTJTAHhIvNH3JRJM/0
XbVe9+sJPO6ejq6JmmQ2iVfnO5am0y/JHU2k0gawEtr7HzoX6ALiLBBjvJQ7GybW
64BDuEc+f4eZiNpI486LVkbkTHn9q+pjpePIrsdJm754XHb1dy6mYAjdAiUpaCJ9
T3ByGqOYVQ9mDi07vI1BKbto4/eIJKAdPUrB0TYNrLTW5HIcr2C7KjY0Ehq7O3Gg
lF/XD71oU3KJtggTuebrh3C4JocbAAbTBUPXEZrrSRTnfE3tvCCiu4cCxFvDjIMQ
8AvokYmAG7tO7sAUBJJTG4Zh9bXnNsEcUkEx+TEHIWRc8aGZ6hUAbCmEcuePVZDc
g9tHD+C3YWh0RqBh4JSkE51N96F7dgvHpyiQRFfqsuC2sRHPl/Me3JQSvkOwAZra
la0kPyDzBg4zIY86iZ+C6yzwWBxisS2ZisM/YU1JwmgB1et5Xwpr0FZp57/9+xY1
HW9qx8giw+YMrOYnYam97VYDQkwcnKM8tTex+/PjYU/AaW0XP4veZtRZHbIM/Xsi
u1q/wVyuFwU/9ctJFjPwnN708pbLTKLQkUewUZOLWMt+yeRHBY8prTq4UKYAKWDg
AzaXH9hbgjJnimil3PtJQlQbNBiIg1GKHeaOvAEbn/NylxWY3xOTSM35sGl+kyZa
swu02iRpKqyTt/9jOyKvRCaGbto3E3pOwojilV2kL3Uq3seK8Nxr3MryBEExYT9x
tsWKcek/PZ8cXYCVAnCiCjdfAbUp3PopdpBULSjHpsKl/yQP/d5egDDlFkvYTFyy
byvOFkOoWDRkdOscJjcBo6Envkw+7NY8Vd23iQY3viS0m/lVTS8GwRyXSDMHXpkL
x0f8WnzACst8Pcu8ijp2s70oFGV8uo9hfA+4UX0rMbhcnRLr05Nb5k77/Qu/Upjo
H8We0B7uCMVBwwC44kTRiFi2KVRNlLXgmKYZUf7WA5XjdoR0OJYvmxBG/mfv1yNS
YJroazz52wC73kkNbk9TGxg8oVlc5C13TvaMj5WOOWLb6TlPNFbpw4k3L/JyBJN7
VLezf5MW9q3DrnmNOXOBPfkRLi+id4drBYK9oSE0jfSmKvWVl5q0J2PKf0WnY7kC
/gJBrvbvPPaRMn1ruTHNVBpo52/TWije4eq6+HqyeGCkci7kuMVudLpJBokdQA0d
7abuqrvdTSGLT1SEfyP2poFEfCdwl2VV6+b9boK4P/cGajiANsGhGY1lijEDFfvB
lWY9FHJxjz7dUV4EjHy6l0TymdG2mcTQ1XIeSE0k8nEqe1TaHID6HPCk0/nZ99Xd
fY4cVYjeBIvTbBAw8RaIj6cguZhf5J/WkrWk8N/LtoYXHz/9x2BjBVjkqn8S/sVj
xhunUAzdxleuvjk9NRAam6pHQNnd/uk58ObMWPFU+z821aP0T8K/1Eb2nFgjProL
QzjPCPMFajGOZ/NkbrgM6vCmxmR5R6o3zXOVIpGCfQoQ6MyU+s2GaJMAxKaGmck8
BOFMi0S4pTGSBaf8iiDb7jp2qaxW2RW6aUjTXNMLUxUeBVsh3MMCySWGuICBJH4E
tGB8eqJr/ja7QSOqTOQf7n93X97XLFC6P84qyEYik/336JRrcpaYdHtcCArF3ldR
UM5rogplYcrSb3NUIIApgz22SFddtcrhQSHYQR2f9vErSia3l17DcAR8gMxot5V5
4tZTfjVNvacIHUPtMDR7P1FO+rCvUAqnleZWILJ5LpMbMDe8staAYA6ThoZejc+u
OG+C/WcOUVusJ87pnfJW8xW7dBPZ3gQ9o3eMpDfJqvJv2ZDcleutTN4Qkp/bdfWe
nzA+J7zbHjDs3vy1hFfJ7v9uw6PTj5LsmkFJvxVwNeCn32WzQEN/LtAwUCJjmKre
+RMrYSq9lsBpKpZlLIwmumX8c65x7vMpGsPxLoGj/HQdfAO9PGC88rrJQjZwW2tA
eAQhjKATwRfl4MeBL8j8vk0EuDPKGJ3Hj0vSt8PfHKNtyxMAs5S93Yd3SEHt9U/6
XgzNXRrhht/sRrL2/tmxt59AKxuGP5p1f6n+0rV9dGVE0UO8lHEgdId9viRfkVA7
NSK8sPvpZ+DV9z7hL2sZ3owl2Fy6Tfgxs27Uljddyi8Q2+MbDAdtt5zvYmJH2Hp4
HIB/71HIioxKWj5kfAqzjN25ZtQe5ef/RYoujO4Dc2Nx5zWkk8riaFTVHyaymEBW
qy8YuRQL+lGXt+elkL9d215GQSM/TrCqgIOoYuOGmOdijEb1T2RxX7iIqbYp2Elk
bcqOmb48ceSGAr5tPqcqTn1d5OuhJjB7HQpnO6JnsCJMIKbslMzKLIcGiIW+Jypq
gVuiF+wbXd/MCYhh2AOFp8N8IQaM8X5C2jTGtZ5cG/iquw9lSj+LYGJtyBsCDnoq
kdZdhFOIkQt6EkJQ5FXng5M7/soO+8lkbyKLUgD2CEMldO3feeVDYMvEtaxSc/Im
/+MlX1CRQ2fhdkC3zHFNFHrjehro5NLYPNEuASGAJsh9gaIf95xefdIKVSA3k2O1
kzkx5B47U6a1mzRitFX3PHmmrzURSIYc7eqD8g3z+gIbIhpjGf96LPly8ZtlLadG
1RJ21k9Uz9favyz8nRdT7GXXgj2esRhO7SE9iyIHacIIrLgJJNlWL6VpBVxyLUQ2
HcugPUVITQpI0SKB8JMG6D9gH3TwUcCbAMmKrBO2vUJuA7t6nMUKI1cGS77zym9h
f/NaaddaR22squD9MUb5Ycy4OjolF76b65fdRmVCp+thOTZEY9onrUdqGEJ0Kkmi
47imuJze2ns8JFGkswMVUDBahObqrIDNW578SjksATf8bI1kzV4/hti2+cWremF4
/CTtmdDcoiQIwziP05S+X7RB7x7p2MYxC277kEgyhqZZ9DfYkJntjPoTa2CNTlNT
wf6znttGY0Yuw3mZ4dNsXsVwzeQxT7PTCSL+M8YW5E+tFA8y6klp4pIxZi6YA4w0
lTnpLICGpXwU1xGH2CeUw6V0P9aZxxHfJUNf2eJdSj9G6gvgn0tABrGPZvcyu+hG
yInBNaXn0O/D62E50vPmrlFbYV/D2VaOZQDH1eadX9dNGRWGmKeLPJ/EFHKwj+NI
THUnxiRI8D60h18WXLJkAbCmvB/b6w8H/vP0ad8rAwJy6Nd0lBfuggl5QKbmrsrW
843EEQouiebYbt3REKWE6YbNmkhF/OcbXK7PU4kJgW4G54UkMAenFwPV8VDqpuOK
pBF/E75BW3KDTHF9s8KdKD0VyqQwnD6mu9U62ujpbVa+8ySXnDKipiAJQ4odUF7g
XVSazSXfN06a9/raJrMYbKAoVgcFLZmqowIoi+BlqxJ//V7gyVK0WsMy8tlro+d4
7npgvMNDb4WwmHVSzm5IZZr4vQ5IoawuGUbV3cZu1zMHe9CpxoR7j5mZpfZUHh1w
tYiD9yGRL9gilXaqoCiM8UsVGN0a66BAYsibyZdxLhJjdWil5ZK6aaAu92krQCVd
TT0FSgrpYt49urvTXLmK9fIY9XShPEW/6zJs5mKV/XIKjcaQIzJu6lLqYe6UTjYs
CnQPAh2QXBBGOdaFN7DDFjR2+f1S5R+oawlWhTHZwUZeH/JBsNU5EbKucxlx3LGn
G2eh4hXD9AG7+E56v5c7CJJ2cC3pF2cLkf0akhRRhHStVqqz5k9lBdlY16SAlsb6
oXpnxVlrQeMmaY3fSXDbwuW7uFmX9izPfu/hSsNrwepNx5+QUQoQQmCQ2Hg9Fv5U
gKF16qVvYLg4c3PGsUMdvfmCarJCXUnFcq4G2m4nXwTvuRNN9oKKaUv+5gs1r7WR
x4pqPeazJTYJCIX6wa/1Uk/hbvc45vj9/yS2UjPcm+Cd/LngFVMQPKdFjso9TMoF
ZHcUXI+bXtx4Fci7Pi21G1laQqC8RPCTOoetc3JCkw0QyeMYVrYso6xvrv3GyC/z
soHfvSZIasjD7moG/fm14SfkJmtcPOW4vwevSWhVy+T/N2Eq8vvjU9eGsMZN9XJA
4dHxo6CY1u4isRtNdCpnN48e7JzE72HlmK3173ckoQ/oL/HXBywx34R9GVpoVlUJ
lQsnaUoN31DNGudeIzjK5yXeblmUvziO5FYYC8hSR6hTv9L9hSGErepaWh3hJRTp
2riP1qulp8fs6JbCkK+5HCxFkPwUJzv/jKQAGeBgAQBq8RQDCdvOvobONDFLyxu1
RFQPbQhpqS7OzPdIF6cNVyj+R7782PJf+qe6xVdeJCo5awOygJuKy2Bk1yZ40BK4
a0qjipiXSEdwbXlKAg2kdNNDJFZKpFwtoaRTak6D9gcW7XHujpCcCVKV4UfxRuIe
SDRQRXcq2luoG6SmdqyvJsuW7uGsJsJPMLi6bXhN5SrqQcsZ2JWTRuxj09wOJ1tt
ft0MJgR9tThzNxrDQvmVF5trHwYDScGDM/DOLn2xuvzwvq5f/R9PVYJDPCvku8Yn
/b5AtOpQCOMF9yluNXrmVyaE2nWtMrWTJctyl6xOQUZE0qiE22Co4skMMN0F3tA1
xf91cPaX0rxSzlooSwkbjLLxeIiZLIuvxevnW8QVrBw1CIt4UNy3wA0w8bX+tuth
ZrJD9BnphnYjR/hxIPFIHTvF/A04JySVXBag7M9Efwv/eEIzMHo5SCCqQ6Lh8DEV
xFBglsHgWOkXvVtuIGIUY4qR/AudJaiYQ7M73jDUkLyDl2Tve+l8kIpXHvElx11q
qfGPxg/y1oREnw/UuckmEVcN8usZoIUGd41y7ylQvbkm/NvtvGQw2GNnyz+NOhhY
Ce/9bTmBnbHTz8I3qUfByBXj4a7u4R9z89gY83fWTJySn86dM0N66QXI51kMs7Yw
gJi9VSqdp6dL8w08QX/I8up4bTUOo9k36ztxpdDrjhrrpfFLXkUhaGbQtbnLnBDc
AvZF8eglnoHMtxhtTxKQ8360OVEXywz0d/drujcv9EvAuLS6fFMm/JR8JCzb+Ttt
du3HhR/wsw5hyKKt064qFXgQAS26M+wYsgT1XkfzikXXBFSAD1LypMsx6fbY6PTe
jjS5mpPgElMwd/Qo6W7MMV8M0DHblHyzpu5vl+JAi43HT/ivMBGzH9TDRH+/DSao
WV5YaRno/5N1p194ZpCwDHuKEkdtus7KmJA20lfvb65/XBWsRVG9D7NaOoZgrqpF
c+PbDHTgSjRix9wkMG9EscB7Zy4eVEGWfb0DjT4X/E2aDuCb/shxRHA9UakIPAB6
GSk89vQfKgrr08220RehLS0fJA2GtiucitT8p13Ue81ZG0ki9ae9j1kZgkc3PCiq
nh0P8VKf5T8IwJg0964KRC23gLapg4t94nJWzo574gIYBb8ZkdjOrRy2eIvgbSnS
3Egu6zZdGCUnDKW64lnge5XbpiCv93XstchUxPB5KaxuaSMgarmzH8B4z5xy5kZU
SklusYP/jyjECKTctM4f9p8R+fb0MhYR6QP6nOWUpjSV4dQoVUEPBk6cDQFwtQiZ
DKc0/L2HFNbemfV1dRLHpEdMWmIgXmsvhhiUkqaLhMtv+AY12cPYFTfNL9xi/Dnr
TPJ2LIxy8DgTERaCA/6ZNSveFvnoSpzB8Ah6wrtq7X2NJwAiEjl7ptb43vOn/XDN
NzLiVXD1o3PrrQGUufC9YvKo8Lz4UWRaI0m3kwsYi2KlqmKDDhB5yFqrZPiNLzly
KfluBa8jn+cMWhvJDQfD36eOm/iXZTqcLvMaHBbVtSXz0hWc0fzMck7/kzJE9Aor
d9S2oyNrF73axDzeWsOUEVn7QmyuTjPFfRMRAVGdEW0VzLTF3g1uMI6XibKCBVmh
PxmJABn2O9QsJBEtZzcZGJCZ8LzN0yxElO0ic8/YPPmQ5WHEiFbh52iMNsGiOx0U
SnwawzQboNoVt/7GHlnyxETyD9t2mQnyRop9i+qCG55QHdViIqjcUlENLcX0cJSi
GgRTM0AiY+q+qnwsiepiFxfjXwbpicQGzQAUll+4hEsOe2MKyDkVCUr8ezX7qlty
Xra781JZHX3FwcttyirvW6EY68zcmTRV0fT2F08zIwebpF3KCCeS8NHcvhoEQEI6
Qov3ALugCENR/1nOcRzn5XXXI4OZjBbIGb7Onu8QpzS8iRSRnWhXUtk3Zk+IhRYN
qSuD8uhQ3x2B2DpqTUqb6LCPnWnqRS0soH3YSDCZYCetI//6nOuRtBNvt/rJnw43
elkwpa44sbHDVRK8/A24AyGsd8izw5FYfWwxdm316LGcP8az3bWTCcGT3uGSQj97
djtw2Wit/l/aHatTJC3tR+67ZuE/mun5ZQo1wIleQXDbypT7UvLFA3Dx4BiPeElf
B4bmKJwf7NYkjLymnsmhDOY7BydnWT3r2XK3PjQDThgczs5ei1mIRL0Z3sLESpEA
wZ588smjslU6Ti6HaZ1VjDqg5w7ANkUrpaHZ5J8Gz4S3ct955qbqQ8hKKL9tLHR4
SSeQldI1Ul0nYKrBREX6tcb9kRSbmlwjgTw9+cI7Pzbjp543tdmo5R0psOLpu0WP
t1CtUwkY5mokdLzMBiqlsNsoyzOfg7O+KCgq3J8NlAlt5gk1KipnkIThQ9pPaUzj
wn6VZKJwn5RGK3UWCVreJERPOdaG+8DiD9Z8sTNDkfA10mNRL0rnhAfGs30eAnpJ
p+k97KIdmtqXlZqv/DKpmJK+nOVhoCGFYg6bgs75I0BCTfUSD3mX66mLDmwU/kp/
Loesgzn4HT7bzy3x3SLZFwMUSJG3yhzvVA85/Zw2rxsD5WjI+iY5SvwiLE6QdY5d
240R9qN5ov613/4eU5GYO2nT3807d0j1wweOjhhoUBUBH5lCyHChAvyZbCKxcsNA
rgAi944/RZpVwG0yohU6vEGuikdQoCaXGxdM2aXHKV385MNknzh1U7RluItBZMql
M/8i87W3yS/2kl5AItEzTHptsD1iNnI5awdeIDIMBC53FBuunQUsmYZOPNuCXjRz
Tang9p5YU34ZB7nAkuPgcIhtPx6xICyVeqzXBPht6B9I1nxzAc5wPVOp0cEFwvku
UGHMBxgP48v058IDoWfYpiG/yZBKIIOaS2qOBNolJcsfAnCvsxYW1IsHtaChz3K7
j3fm/krIPN7v2nVr+p2EvrZok8pI+JChZxFBbCBDymsPDh4ZiFUYNsoGHVe7+ooH
T3XbQbrrXf0uD7IMI+YTc48O4VceBFjwu3oBbhYyiH4TmZhIXlAhjYyvWRUu/nmP
bi7cQLIAYfeGsWqjz4wLJyEeLsH1Sft6XuPuJqtE/Mhp5ssnor36AmonwgjOoJof
ItbDz2en8uv4hTtQetcawnYlfZ9XBjgYUVO2zuBVF/sZnY+Tn8oQEARGstMg9kjT
/gEZ6HPt2icLx4FEbAaIpB/DjANoaTt5Z3KzzjixGW0KWvfITOaK/MdOu98qWAPS
MlUI3WROEllyBJ+LWHpkB+asMijDRr7qHKTe02+b/yEapMdVhUnifgqll/A/Xp6l
hNyf71/fgPfD1pdKekasTKB1zqpdUX4wsHnPlIgxUY6j+/EZumtVcnC/mS2Sdj2D
ZfTEMyBFQT0811zpypxNBVRMCxaN9KxNDvEnayvph31/7Hw0Tl4DggG+gTUqeGQb
4nEtMd2is8U5dGKSDzrAGfIjLvLmViMkXeCTJwrH5KtDbTvtih5nqepahGEGpF4L
Aem0ELb0TntC69nFh62WIWAwM5z1K/zFmvWtv0jVCWPgNtPd+RD1pjXp2vAiGQDJ
cW7eZ5GDb4rVQ1h1tBkk7aHOZhp72WkW5sMRqS8ek/ynZMLsE7C71eGHJRzIC5OA
U6tOiXo0+WGvrt+LWxzKIjYJzbxXbeEUJoMZyznTTo+jhlmimwq2s1QYZ4Cht1b3
vmS2qsYTArr6MG1BgAWz0OyU9wJh/UaSeUS/FKkGhYXjmdJbDvdhaOuzESQRD2fM
CCfnuSsx6r05M+S9a9ZZf5yGVCLYZiPYQDw7R++D3bEsRs6AB8RNmy+rUsi2o/MH
Ik6w++/o9j3ROQ/kbonpYyrLWcNovEsgU89wivlgo2mQNKeVv9JvpKUjTzIO2TtT
c8kyBJ1lRu+sKU+9kIFzSFhXcZVZNX42nbAyA8eZ8oiWQ8Lh6UlihjBhkNOfj8BX
z71/AACuFdIfbx78Af80B1K2X9YVqE++dgSZfyxjV+70BugmNKxlN+5eA4ouqqu4
YgbghJnyWKiYbHjIaBeZmG5Il+e3nmRnLukyWdndSX4kwYE/kzUGIuAAgPMwBma0
rInOcD/u4Mew1xwZ+Ocyz2VbzWbixcbtlgTPdsM2p0L7Rb7F8u4NCEn7L7Tbnzs3
xP6N5bBBQo5bsKNuKvp8+0pe0fUhtoUiIGCv07Vcbq6FgBhjsLjCIi/tLn2T1iCf
Cdxdm0rwNCQly7SFAvsg2Zyu2EnCjkSo/CuscO2BagTf8fgiYoDO1Jo/iEe23pna
vtRShMZCydq2KtQ4LuonlR7mqLkssqpNYYBYQWvbZC81wUFZTsQHqZaJj5BBJXKR
yhGaYt89DeNECRljOpmZCaNR4DVIdWbCphXXs/7lg7jspAvdHopUIFkp+bWcuAJR
VIRplG0u4oLG9WzGl4WTY1362VNwLbxKc/M3sDvRbj8YBUcjd2LTnMrqawYIfT9t
4JCfAIvqnxUKnBTQBf2dF3SDm4JNO5iE4E4SsAbvBC5CxDi0mmg5mrh/z3UEIpWT
5jSvUtWGYYnvK3HKQbZ621O83brtNZ+EjWr8neZ6F7dqyiG7Q3+NHLDYm07irPQK
RKIrEwfGhYOOu3IBd8bry061bgweHejBcfau+eff3qx8TzS8pqrEdC0hHg9yXkQa
I093uCIHPHeOFmMuv7fh6iMvExiN+sUeZ4jpu6RZ1Nk0TkGeq7CUvu9nNYfbBhks
dYXM/mXvmxKrbrThS8Jd9985Hs9HgoMBqCrnWa21QxgN/iEd2vZP+GSme4RgJk5h
u6R+D3smzbP0dzNQM4bXlJaApGnTK9MblBw4D4Tr8JsbWdCAGXmbY1Yz1qs6Vpwn
EIQnw0D+ZCpuMLDbC9n8oKtHnjWzNDNu/dYO4Uwvy5uRzJ+tHTnqG5ZlnkJiaqZQ
28P4NCmkZX9z+XQ+eaDnlpZK0cc1Hrzr1Mwf5XoFOqwoOQrTBDF2nGIErW0j5qFl
v0WEqtyoTmKMkIM1HUThO1m7U6v5ZXhL2UPdiQJj4cAJLC/3Za+Cs2f+jgbSHqhM
1q9HSjJD5gOhQRm9z7gz9T/xHnHigHGaN7Y76lpodk/Fz1PdH7yLvELYrAyx9eym
i9pNHqbT5/g/aZ+MbPlAF+u/hKgV9FxUfgockmDh+GgkUlIxgYpy6V4EbhYIaUSl
21Aox1Fvlpl38U82/rYwIbpssuq/kvXQ9YDoLHeYEq+pGaFbAvcuizsC8dgNXXJ6
wfR69UnGQuRkjcLKHedM94WMeCfqgCR2jPvoJ5HSPGS6BDL0pFYDt2LVsBcYoTQM
vJjRSGw4qXrhwm3wMuhqaPTuagw3gkguJRHSKyMwUeNovM+oeH1zQYym53UZl6rq
2+yq/45I73uR6sxZPB4OXtWnuMONCXaoonZ7G3BR8M6HcUSAfKCUq2pEerHIBq/o
1lrUwd+IMYbZKAZKL3U5LUry/+XXTjw5tqapXcVMqVS/+f7V7pLaWB5IDQOzRAdm
M+9DTM/12LmKi1nVzjc/Z7eIkqzf3/XqaLI47Ypi3pfJ/y87AHQuLNO5quhDNT/O
EnLaBBhPkVJhRVPnaPgBvVP9O8P+DpV7BfQd184ur8SCAJHlLVRztt602tivKBOQ
upSJQij72/ipb45MJpKYggtpDxM4HQA/MPHwRd5p+0FV4Mf0q3ZG2z9gelF17ag/
PNkkp0J+L2U9cXsWZtrNt9y4pEJRGHLGVPniDHIEUAWuqKSKue/SZhYKNdeLihmL
nvrzC/vxKpMMgA9NnfwZED3DGulxeUSeHhSZGDC0XMuVylWUPUAo1dE7e0GYobny
4QAZ/EVSKOb7POJzUoCPMZ7gRzpDFsJRL8FkyvaO6gkyi2b50HQJI/v0ZPjzIGjI
gy7dFME2Rt4TiPN74BbrmFUDqZFKT9aDzMLtlb5DTV/0pIW+HTZHYKpJ0UetUXqm
aw3xAxde5Q+VVrxt1iauDtf7BvaQqFBovLRIlVlhhNZRqJWkNdCer8drScOpe6yg
VMf+n4td36TqkAcidVl74cz+UhcXy0xI1G5Sz3hNqBXYVKROBU/HniiDYcWbHS98
xD8kSuHwXHQk93q7IQvufQU84oaYqspDvc8GTw+pdSWFRaVyrazVLNqK9HOzY6S+
WSmEhLaPc//RrtL58RrJ7G7yRaSNiGe4kjXSM+olo3IF5pTig/+eF57gXuqpb4Rl
fao2FYXgYkZbvIwmKigW8jofm0to7rzAScmeESMuUpT9XJMMGsy1hf8QxEpJt0ag
IqLoowtw/pSpQ6JWA3lNA6AtepmaOwpg598olETS0C8w1KiL1o+AA+unqTMloc+W
0be/q1aVDatOIIV94Gj1F1ZmE67n+zBcqfYWwxmOOqyP+qg246psasAt2fm44Wi9
+Ozi/Zfbp9V5jxGrq15R0mi11jMXBfPz69jX33IM4ojGba0EYjv2ak6Z2UXZjxbu
u1tAsIlc8fiy31ICD09UW1mBrSt1lCIVZ8D+YnVhirzyoFeP5IYWkgh+aEcVU1qN
qfX+VnxXUM1B+zpbEQG7pWNi+UpGg1XvpZSkUIEQg9dNe3eC2Mrb+KorsH/zleSE
VGX+DJBieEd7g6Mp2digWC5X24fn3zI+zbv1FpHxMfSLQBHOJv3VCvWZSOq/f/r/
Xh9YV1RZhtEOwnGcpe3PREND1xjdNEEEfycN1iMu8B1ifo3Htx0swXA8JTwx3PRc
+lKt56x0hpNG3W8E7gwK2xwz10nZ7dSCMMIUDbxXhph/mwv1kfx6Wb/YvavXAFBf
UCtnwyrP67tIAmu6nQVYGNpCnK4QkI8LaV9CQj8jq19CvjfaxDqwCd7sKM2heGuC
hR4u4/OmunyCQ3/kO0sMEoYoCf1kko638erppmcLojy0BLacbLdD7yJz/ZFWP8OB
L5petQBu6nsbaAkp9bYed2tfiWxroL4zJEhm5+hjGse/QJoOs3Pt8GEFW/zTfp+S
gNkT4urbPmELjQ/OZSR7kg5xfc6WubidG28Vt0QjWn007J8f5jb1c+HveXWNZ3Lq
6Ic25FL7ZVkU/S+3JzY0la1kuMfnjh3nnmbdAi4DPwpbUT0TBJU/b9kNhdVwJBEa
jMhMmvWg2MZvkF23tsGI0Gce4zRg03lha78mAYVEi0/OAQWP6mvDKng73pD6wXXK
RKvq0JQnnU6kVGdaZoYk0M5f4WkCDxEZcmeX2oCYmq6+hOD1SAtHFUdi3uYZg3lY
LNi+6phVjlo6qogDQFS5Sc5CfPRrz/ZskrMsPoyko1TTnnOTfXr0sryVo5aJtXV8
SkMsLJhnVpDqROoL9pSeXR3BRAKG4LgPpqvnbhSFC3UrcXLgyCDX0psX6OtjZXec
bh4rgKuJigwELRPrQIglxf4oPaF1q8wshM3ybqE8Lxx2D8P17cK5e+fEI8nBIVB9
O2ZoCZZ3pwg9NjVEBnSST37s/gX7j2crRqZIrKUADIlTz5LEAkyOTsU3+dlVvFfe
EpNc176Nwqo1ITxKj+5wcYxtvny2MJKBu090tCHl8PlCOvaYaROC7CbWK9YrzUL8
qjrR5AMIM8uv3u+UYDgRWl+kmwVReRgegTSA3vJU5CFOmz5PtdgFyu8LqhvtunuI
ZRnUJsv96EDT3Q5JtwhDD367Nfu1q/KK1MEo7A9YEPFWNAGDdg5hrfpxfnHo01nZ
kGLEgy5HxX1YkzlWQ4QZeS/4mhyIDgdYD2ft4gHMyFN9+9nUyd09PY2e5rhggYbT
hWrASMxkicXuFzD48M85/B9RCQ/sacCCqA3Fu1PKrC3pNIq9lu/szL+bMUG4Fjx4
hyd39pZ2bOgh7GMyK+Xn0ICdIymFRnyMvOVrvCZPfiNDto3AmIap35FJ9asjrxSg
vMmttkVWyIl9S+pQT8RKIvvfsuwIfSqtTT1Ay69x03alX88f69lLVSsSECp0ovHd
BRCB9KmrSa6Gv4qXovjH/PIna/jTUOGEEA+2uiVNeKC/WnIOLgo943FOzWwf0ELC
7WDGsRaCH+4MBUg/RNDJPNOObu8is46he+2HBXvF4wVuui7iftw/8VEYlgUDQJgY
7pxDoOwkO0KMKVdYs3IZMHccz1m9362Qyft7VOaSdzNkSvs4/ekF+D5Lnpl6xd+0
ED3qxP8eGZLGASto2DFYB2ypCql6CSnd06bc7vNips5DMEMWa1yBEtPbSRk7tCMN
OfIRtLewDA49/wnVcDBGqgdagP6YcJnTFijz7YlC4LnxNY8ssrCC8ChTdinFlhhz
ywSRcx9PVx/EMANd/aqgqlGcUa0ehMkjE+9G5iO7es4MC/QxqsUsNPDK8VT6uKar
6dHewTTh1NP7K6i3HQAxiNGqfJeJOzlIXq1eH9KvC7FkkrJdkDLMRbesN54D6A7O
MEiceTRsU9dsyxYTkGF64e/PpbE05EQwCZtPmmsVbVeGcfhjHefh4RjAOVuW3G+b
dEX9/qlsRPg7zogGfIONVKS3ozd4oMfU+ZTvSIjocJZxYG6YSYOZFigSFExfYDGo
InGULfyGOP2C4WAU0XT+acW2JdYZTEH69gcmazNgtAm/VbMVqZ/eKuYi58wAd+kb
A0pHswbn36ngBkWGu8Dmm8CYXYu0BGI7+0Nonu1xdQpuhcdKMjEuH2ixYMIIFhIJ
CmxjReQg/NsFXPCAJMmBwuuUKLydUazWM9h2nBBaWveaxPWmVeaQjIr84lBrl+63
KWjCVN/fcVcoW1HR86ujnQw5Eaw6L3UHnEC3sKcj3fpg/zYAspotDqtTP363VqUt
L28Mqgu0FtBv3xk6Mu1UqsstshgWEt7/Ymh3C8ZXKElkQ6gbWLPwTmiaHzmiey3I
OoEqAqam2gxU3cKK/ocL2y2ctaX/5A+/wk/PdEyVmBs9h/gscNo2KJcEzznzrFyr
b4kDN3IvrwnCewQVom00Iz1zwY0EWfO8AIsrvAJETIy9Tzrt174cbXtcNpirsnwU
i0TyM4xCv2zUxFkxsPO1LlEWJmhJGGXS5ReeRhF+6ZW0P0CDaGGwdUup6fI5sjF+
k5CQaDszdbUsg9uhVK4dVpAyrdg19PnqApHf0E7tHwmCQLoB4q/89OhrO29bFVb9
Byc/gI4HLcUAGOM5yS2iB98B+p4+R11nyPrO+nl2JKD4xtOLftN+7LeIOIlRIMV/
68u0fXtA0/BAZ3vN4qRDd7l0W8DBii5IWcFQloFbf1KwEV5iHmKxQUhYxaIoRrO6
BtZ42sNdaJG8EHhL2xLyy9vCtSU52sDlafFWnHU12zcEri647nmGReKayAAe6M1E
TXK4dSF67jFQfY0XR9F+xTEWMM2s4V6cfBsx91MutENki9XgXFZBTSXsR6EuGkKY
KWwHoP2ZHbDaE/3xNznreWnS95XgoR8fekt8N84BAxdechvgrNR57g9v6FwBcubf
jCZqBPkE1D/2P32pZp61YKZXCbQhcWFWSsSZeTsqmUIyq9aJsAYSpKEKKnRlKZGB
TLYII6g40l4Ey+tS6mXzJMW81OZTwlGn7nRjwHrhHOu31hgIr8wX/YMu7dMzcuf7
BQZUY30HYfyydajxczEFtUr9j2S+AqnCPt+WN69Hz71eI7hXhhrn3bThVtLEdEPm
F3GKynnEsXB39G8ujjGpghW/2AX6BZNIvkXyQmfFfSkLq72UL7IMhABCKKE81s0q
qrjyMjEzYqDIA0MCqLKU3fwHMY5o7Zqe7+WXYivQ5HQlHExd+KjPYf9VTHK0drgn
xK2sjXohxl7wNomqDmx7fM6nCWdF525xOSosgdaKx6VQ5zfn5rtc2XEA1NlghQsw
vPXrasGmzHTw1dNn0BykwXhj4SH3Omxe4jzRUBXsDxXJq8vXhIlawE/3/VXw6Qyv
E+X2pw4bGIzxpdDc0C1ukCHSFR5M72gOR0ahYQaJW7TvCUMv2xO+fOicJ5mc/mpO
/C3xt0W8xV/hK3dLqdC9lWUoHu1hzgjgN1i4bdlLj89YROGRXs2TRklT4HltJPxn
f7dmNFZQOss+J0WKMf+a7Cn/PzsnLO1eLor+4RNFXNW1qCrJQSXxCk6hpkIfmUkU
dNwm1T5dEzfsO5Q6cjKWUa3OnzFEy/0NX816FjYDZCIiimdyPMo4Dy+fynqAJIWn
4wn8gKd0rZ3uak8mKaADjc/a/LCLFtucsr9mxQQF0I3njaEcz+Nlo1bP5XKAVf2G
8sMXmVxwWCynEfHL9kObem3JWybhNHrHk2hUdtd4rI0XldfmJ5DKrzvRTAdnOUHA
a9K5GzYfX5IPhGw2JSWcioEMJMs76yq9al0gf7AU64duuhiDJN4gV/fmyfi3VDOf
42mIF4kgX2Xs3MHQ0FxzNm4c407wwZobDFEH2wevq2l0uxAj545L9i+yFdoGw7ux
Q7OZ1xpMPYYRH2AtklrU31D1Aud26MUWRioIXeM4T65+Y/Y/4voKI1I5rBkPCZZW
pifWtYS//yMZf1LGBkLVkkC0SgPNsWkFy5ypYyr2cxQDCOwIO1BhjHPn395ENc9r
fzFiDkIw8hffq/Hqat5WQlYTHJMAaahR8X6FnkS7uXV4ZLSe54zyZ31DWa7arL0Q
oOSEpQX7ciNzio4gbwRnQYGs3JvN6oF3ufVRbApkxxaI1CPj8O1nILIpy0imtPJ5
IleIoSC2zDD2srFLVNulwLzrs4gcyxxIXbmPjmjFYzDRg2g2eQQvC2iDzOp9RlSc
eVscVdCV+Cq9AO328c7MnK7zKoxYYOB8a7oNBur+FNSSmAi+Nfp5tXXpyQfUSg/a
lF4RF0UDl93+q1sLoOEG8bjy7iXR8WHLEO6ADD1ckLewGu94Dp0shUSbAbo/U01V
5e30vlJS+/Nm9gkkcHil/IpSHwiv4RUcTtdmAaEAM3JLGgYcMHLvsG5JmfK278dA
x1RDOGY9tf2zssSCSIXZ8FAwR9bxsOW1LoJkFkWIm/GPu4qn46NA/1wXnQOml0Nl
RBr0uL1l/gBVYBa17KqnmmW7XCh2ja7rcjPMCcy4FxwEVWFXBQzoRYRbdSRKeegd
ku5pDbZ3sQ/FItbr+yhM50mwECimrEuvEJsytXIwWffFbDF99XLbHaNvCF1udmic
i4EiuFLKxt0nIdm7jAUukXGqbvt/GopJifGGiu/vsdB4Dy4HuypV4N8LmJHJMN00
Z5ONWrYDqV1JxJuUcmulOQWoVGlNq5o80P/lwsTsqrUBijGbgGplCv4Yf99y7fN5
suDF8/NeJ/PL/Vn7YEWLbgReolrpf5E7xvmzJ0TeQ+/7H6Z7+jBgxQceO9eEoM1o
pdmTS8tiU92w9VlxaXfRuYbOMeNEvktNWDxjZhF8IIpdtGgLNkjvRF+vcK0O8RKp
Kgp4dTUaPrg3JNv1ekrE/I1Q3fdCYNIW+ayygIIy0Iyu5qfkke0ppoWH8iaZEdyr
lobks6MUNEbpuvh3M5+xoXg1ci6Pb8q8azzxVMaH88jZygJcrmtajiVgHc+fkH79
AALWyWP+xInUy/916TYfmrRCnH3u/MQyegF8k6+sd80sz+jxfIbBp5ydINJf0mUZ
lg6SqZknMhxtdLYVNMQ3WIQNITYWnmRfbs4pNIBvm1uwNuhTxBsudoYYI/tHcnr7
jAMW2y2J44mL0L/8763PSVNty3FWli8qGVsApUtlP4CfisS4S3mUmoKvULZuXpKI
KTK3Fion81AXo+UmCed+ZerbC3jT6KtsTOW6EUfi2Eg0lszvc/g1FyBpasdDDNY/
diShI9SHEj8XJqRexRpWVf1fT5pemuQGsdJ2/W9uyUYUSEfx142N8DxgpYINmQIp
QOGW/XxbfaASSRLpjsoJD/9OLDFfPN4CsZN1Nzd0nBoFh1a9vuCnQTyQo/z3ViTx
P3t37sH1bjCiruZW3S4uv823FRbpBAmNFSYMWHQs7rSTBJQGmeP7kBGRRjaDIs+i
oGrWVtJT0p7wsSt4vmb9wtjBiT2VwhpvSjPHnDi4asoWqcvSKahGy4oK9UUMDeoS
5uThS3JUT2H7mwFP5iJjAUb/ZH+4zf2NdiVLpxQNMPDF8e+ODTk5TcXTu6BRCRjy
JVVFFcPyivzS7xx8YIa3hoppK2iGBvxUWGJotmgKtIpyIc7DJoPTt/qcNHuXA7hz
nzmPbHljp7SN29ljidMqMGzJ4VlVCLr7usBsdYB4XhZxg64AFE3BizZ4OLnD4c7v
TYQ6Z15BzMGKhoX7wezhj/LuoSK601pVsd24b0s0MsWG5Q4yzTg3evDrssYRyfSa
L2dD2Qc1lhSBdnc9XD1+6Fc5TRCNraphyA23glldsjKMByj/MCmTHylbkk6YtEoK
/wNCtWt/NSv57+0f0kQqmS1x3NpeotqSubrCs007SGXDjZmFTob48GswabMdZLGR
IXsRi7U5HVL3DGkvUXrAX1kZJZaqG9LUPHqRXHhHQl2z5xPpFtNBtqDfScvjvXzs
kJSdvBI+maZxYB8/i5N8cDEU2GdQWGnEvisWAuqsNB2YgX7GyzFhdnzreR/wfrTe
iVunjRn1EBwQ67XpwG86ECVXJPn72l8sNzAyvCBW0vSSePkA1dxXR0CNKmFDq+SR
dBM1DRIxVDv+CqMTzM5MPWH7zBr5HZEmElJhYPEfzGAoFUbsrEgLRilvwkLFdIzj
KcfhF2fCsAQnyJyg2uV6YKlq7YWAecIttjW8S6Lc+eO+KWZfJHuZVM5QGkqOZaNq
qS5XY/EzJBqu+GlxFD4kt+HhNE1EgO+m3l8dERnM8HO8hXIV23yaSYbt4+CxiA1t
McadEO0rBwwl2PUjh2aox+m2BP91AGsAwMh5NxJ3oORYxdqrhR74bzMudWt0qg9i
Krx1Ls9f6BkVJgE+n1LUIoWtCi9ixmJo23hSWSI1DI+ZbJAW0n28NgW8kJyttVNV
Ayr6N5TpUsYJ8nHfWswfqejA0fkDriQHGU+M25GsW/gHLR0XSWqMcpph3KUCxsv1
Ba58VdIebJ9hbOq7O+6+pFCPuOOKLvU0nxfXrJJ2RIttR2Oq1wstO0kmFKTW1eYn
T6Q5ANsYHWb77VAoRtRBf2rlQCttVhACYDBC9kQqgKrPKk940gULjAKusVrdiA9C
As/dh6cPgcQ7dcwv8iv0zD5Xm0pw743KFfgVnrWVRB1A5qivooKxCXmJdGZUTcWa
2n7xjKf7BPKSaYxeTxQ2bNhV0qIW+fXkqUoOcm/mkSbp9LF7OM2gQYvGLGm5Aj9Z
kcBQl29H4Vd7QIEohMsU8/7ozbypejF28rMNzpgb1n75oyVbiH+eqifoVzjo+jJO
Z+1Bl5Kx3YcgULdIV+TEDtFRw0rUG5bZ8LPA3rPLf924NUSKeGXhijR4xnaDHqWS
yX+yyuJtepfo3rNqGDG6Y+QKRGo6ySvLJ/tbDqwlUlxeXaAcdbgWqwBAl/HFdWS5
VkE/QtUB76aLNmNp5viMN6/NqmxL8fE6Ya9HnrmXHDQdev5JaSSLwiSKEx/5fnV2
LGtakVQ1nNHG9DmvvUvnwr3Z926uBklZ0G0USyJ0tX2BUXu+S1TP8+VfOWwdHy5v
yIQc4rrRJBXd9YGjLTsPlTl1WSa4MkmfnbUNZY/sC6b+CQvtax05pK5+O/l8ehLR
fLnyeTFfTWYX4mDmWIbXgA+2K9YIEQ8hRcI7U92/pRyKxkhCNdSzSal1aEeE9G1L
s70BGkLmvdO5Mce9cY5TP+SlPvx1zF6vEx0XfHe3eOm1u1Sh+DSXsXN/YQL+RmYM
iYff/xCiw0QQ+ZJn61VsptzuKA82f1a6XqufveriRMgF2MNsRPjQ0lC2mRQdRhw3
uC090ypyaP9BzRpdJNHUPS1dt0f3sSfbDWqYs/w5LLlzR3d0ExUDzR41xPDM2JVT
B26cIklBXL4UO3yhTZ4T1/xAo6UHSlamibmS5ATWEny2FVZ/DLInfIxg2DeJ/KzD
zr1jAUl3W7HI5vpQFA4h/kKAeAcS1sqXnGPvCfxm61VlZWPVcDERwphv/pu8UClo
yFkpdDtCi1H9TLIuin/cm/Zb78EXZAXb2TbIsp3uzz12vrERb6Zrei3KWVSF6zBk
5GBfOD33/J4d2xIt8adHBf2slib8X6B3sApWxGoh9Ru9V2Y6HEaBDbULzH+f3wUd
X1FID4rpciG0EBxIaeF8mShb1CrhlUPq8+1g96ue7X6U/nrMW/n2Oz4dQtsrPFv4
S8+KzRJMypbl2qVc4OXPNdqrNTouafu3PC5khkHJ+8xD2p15tQBji2R54VZfYmSC
gTY6vAK4Znkn/zpvYffsTvR8BLLfvear5ApskuLaR5MozznOC544xdq4xEqrGRIJ
8xuXOwm9yLKV4UBxezp5B8mCY/9Oa1V4kmIsapNbKuo3TnfMZleCtAw5e21dhyGi
3hVn9R6HsUMatPS5w6z4sgBWiFO0fGEetX84lb0Zy3vPfVt/MLeSU3uieneMEaia
JLxxyXk0v10BODu9JnUYz5eg8Eivhw7NqV8lCndyHcPr4UFA0ioFLIoSWl46nRTn
bxpMDJJ8KETpgGxBMMNbfCw+MGgFV3w3T/XKSc63tL7VTU+UD/cEXLZ2TQSxMnv5
CJwQJZg4WAuiK305SrwhBLV12zM0KfflIP32RHH//gNxoyqbL2JtKijTp6+sW5n+
DH2OhKcPZ1syZxTq3DMH2qLhY4vifIUNMbIIa+sTQ27kFB2YLEKAS0wsyWlhdLHo
KZ2bz1Dyo5giiYTxoAr1OFRyLCdgajvjcE92E/wwUWfrUbY1O42Ic+eUTI43+jXZ
+yHKzr2t6nqyuAMy09ul+zA8q+b4Oh2VWN2D2qI6fAUNPJ8NTzufOLnQhX8GyRJ2
+TpRy5KO9f7Vos1I12HwtUBAlJ2c05bEtR4DoIASGrjJpnEBdJ0ei9p5waoLXM2F
w6PmPjCE551xdAEbXeIBY43o/OhfeIUxA+18q5+oOTo9cn/f6uU7GPaSGcI1Y6vn
SIGveV+FMsCUs7T21ZoJAXSejNwdwbKpU5aasjv3kIpxOdbh5+o2sl/5AtdSH/6+
ewhRFylAKoVYmCm8keTU8+oZ98CM7GJ09Tz+HUC7JNpjFc7D02pYQnE6vu8SNs4Q
3N8FulHd0fcY8vmsPvULuMLdnpa9n3bsi60e0u9gfJjMM4P9NJQBTrub9MwvsSvo
gYqHmmIFrM/ilIldUkow2FDj8nlrE06faAG8txlgEVnvE6zFUKUHVQwU6teoe3U9
hgCLJLA7MERNXAapOnBpHReJUv085IZcj93V30vrx7/kNmG7FPzBtyTFB4wC6W8Y
7CFykFDvT8n3E7iBmf3hRxMas9srcOC0gyKMuPA3ndS30ZO3Yeoj5aBkeOnaeuLG
yDvOw575I4KzdOUVlVdEgt8AfArJKbKLbVpJwI75KFI49yFcdHuO5LBXfE78o36c
qTElwBsmKOAXY0SHMO2+TjcLxmGu5/6Ye0kcBpTG88HZQkCKkhG+afugY2B4/CAy
PwIsJiwqq70qTFnU14D7Ug/TKiTxJ2J8yPe1vXqZdU+my8f6TpKexPTwx2svqvSN
EpoT7Ob3uflI3mRu4ldqkFfgHWB4krlq+rsMkhUOmpxGWX8m7vObHUfbor+VUcSX
qgiK/dz31PMJbd9Ha+YbmUEOuTeLFiavKiTKccdrhGCojc4DiJlbfPNElM4K3tm2
sWRx1GqgZviq28k+3VGUSxHQMUg4HnjAXYm8o2x3vPHYrVzsGH02la9fXN5A1pK1
mN1wELj8PMuc6v7UF36g+TfBpCTQg0h0uqBdkasHYz2hjnwI1FoNAu2R1wxQ5dAk
1omkSxO6sCFsxWADhFTDtqyIlL9HPwtFZwHAulKnaEACLaGqwNNSCjRUPO9LwaCt
q89ToEhiMvbLnKTJcQIXymwe2qabuZv3MJhXAMieDt0iLgIidB29nrGAZLC0AZO1
Pf9rW3/IyRC19Z7wU74bcNIprdaqWRZycsU+nEsRORWa99Dtn+2iw+n7by9qgVg+
rce8EeyrZAojYoOR2u9XvhhK/lX/LptHKTt6XCV+MKspy5UMlshJdYH/ycre2fLX
HAx5xkkxuBYozTHqOEoGarq5sRGGj9ILKq1843IlphKpKwuylSaHGCeCbtPG6nzT
L+W1+0Cj/GsQvg/5ttfckm8Qn5qvViWfrat3/VaZCNxi8hxzw0bRGN+NwLzMwwIC
qRs6k5UCNSYlfkYwCyLAxqro61f1eg8YinXazM3GJYXqR1dV6937EpOC68Pw1mDF
SQPh1slsiePWYWY2Flk/MESn82OAGanVXTqJvZxeaoZEifGZ7rFeaeqkZP7m1wtF
sdkQrdI8WEEm3WFrd04KSxlHsXKehqhO/f5RP3tAar5k+JNZ87nbzqiPTz3x7jI5
GptWrwQcJPJXRQDB4x0IVDX0XtcmJvMpKz8Oc1B7wRF/0sm5yNHjNrOgnba6CcBh
0mZYrWihXxeyfHCJ97eg25GNl7s4DmYwDUv8EZnxOiGi1wo9OMqdlgZuZP/+K5l7
emlM2qhLDnNP3V4w/00y/d3wlY4LYKEIqE5CHxPn1vLXAF/HFpDQ3BMHTJTyvM4j
jQ+aU24BMp/z57yab2t0KhrTvrJJr4Mh5gZuMfdDE8H4/neTJ/H7br542pMLSKRz
zKK1IPrDjTvcLNcnxhpSYmSVOgXUPN0nI+H1rNugtg82+Z4+YdT+8iE59phj2hZ0
9HcgOSRULioDiSjh+DeLmTLLRgsnvCryovDTnUHn54Q70ejnY2v5v0Ce8sURL5lX
CGZ0Ip28Y3TU3+5BxqHjKmjq/nuFcTqibOxfMmCV9T6jSlZlej/Mq4sbQgCb5efr
ppS8O1OF0bcH6RZXU3e/YnkxycEEMH+s80hp40gA5xLD9IjIH6D131oHXww9g8Wd
gR3o8TH/C53UT279XTlV3MxjHwhYWpjVwWZfAcWqowYzjHR99RX+A1GjUU0V4pWs
UL251NhAQvsEeht2MzYxCnV9E3uz9vEPYOXheyHzcL3AyJNELRHsPV3bw8Pmbkd7
vCejRXDwER264+o25po8NaE2LWbqOltSFk+R4d9rCEItxfuSU9aQlCutUNYfJYTi
lJarUsB6PzKA9UmF45MpVVnQoOVr3cA4bEPkOPgIYo4jZX267vAFsRPP6Q6QxzuT
XTHRAqg1CIYJX8L0YCANwujhUMV21y7qszlpuD93TWc4nRIFHqS/h9xcfg9KfFyz
NI34J9hKjSBUA9vSyjTy06m5baUdMBtRApUEQw/lYUEYSqMnLZiMHY2wINp1kaFx
8H2/4Mr2SaKoGgOAOw/oyEX9JFowycAb+tVscNgoYlGGb4LOdqoSsT9Uf2dafmLn
HddDnVOqW0VisZwzApwOxjNK/5I2bxEhmz7CbkrSzlRF0HfXcxoMLatefRrteEht
3Dcgsln4q3RDBnlyguiznprEr1zITIoqhTwGm7RaM8guYD38s9YIQsLlrrgo6x6t
V7DqLShGl3X1PpK2VziFLOL8U8aFEqImn/1rf2k8bD7zTY9ujnaBWGxKmthJrOWC
rZF9aUnr9GPUypBoxDsrsA2mjK8OlktUwUKkpUvsUr3gMhxF22SkZMSn8e+oQGzU
uU7Kx002szpSspdojZ5GMUHksq/w4PQ2IH39rZrXefJh1tAs8KEmEkXHoHz9JhCm
V4KQfV/ppqMkoHeKzx8ik89Myu3cXpm4Bd2T4XBpvDfaVyWS7c27IdxSEzm8LFhs
b/PKxGMbVsAkf8FsgimweasZn+mEfFkm1ucZYL4HLjslsV9Q5BsGrCBgQorBEfSV
T6aoHL9n6Ivn3PWBgqaAXLwDfaJKN1frVbhkniL03PKcwwIFDZIVwWfS1q3BBvWe
tthtYpFX7eJlPR5GC+ZGcu4ffE5/kzYcQPbCVknxXckQSq7hLb0soGh3um6askIc
Ac2qDlgqI7pKZ4TQNsyMV9IZWYK7cpco4OqJJOJjz6WYEEq1M+89Ue26GtyHf324
z5r8pBRXJXlm8YfkGbr0Stl2PrBJIERE2DyeL0Fw5ujTNTgcLfSWGD++gofnzXo1
OhgbjVzYUWl1tSUrZbU1uq3tOibbrqr/YW3olsEnXX/xCDnK5mAh6qnau+0UOkjl
YJmsgY9OD2r1WXpiM3btknAuL2Ck5Iu//MmtCOxCKliksS5nhm9QXGS70EcCZhiB
MiBX5kzCaDYx6qiKs0xppDqbAGo8jq2i53WVmq6k9jUTEwF/rNNGoKXYfH9uyM7l
gnr+NBSBfH8tcgizyE0zCDUXb2H4edKzRDq8CWVf97ewfraS5z/x/Gte2smo764d
WCK6BisJVCdlPcEEnOnvdOE/Dt1Mj3Ek2bmA4A34y3mzewWzXt6FJ4NqqOTtG62E
JKypmJNWUe0uO6vHvWZ9MazFwGW77GQCn2NwTrIX+Empj7yp3iO6swXXMEfHkMpm
2TfTyabedyQcSAKlIKATZMe3mfsXsdgsUiUurtaGzmsO4cXgb5detCqJFySVLWRv
78YPzJhW70BEEYXMaGomqF24UParTdi+fl30ZweeZAjrsWNvDJ17pdMa68O5yiDt
WrmSKrQBiqNUFDbdTDQrVZDUTDxrDL7hen1eb4Rbv2iEg2YAkXwsIS7g5npNajvb
IN4qfvfCClc5R8QUQZvpBtgae9lxGCmPCTxAiQp6dDDmtOdMiaBp8QxhdaD5PJ2Q
kNrECbeVmH5/k8UfT7WJpfeKpPhm1yrJhrIIwFKdGvaB5BdZ/2XsPf9Iw1dd1Bfb
mg8ESShSZqkZdzF2o1i7jkI+9sxizEkcNWvVl51T1xEyO9GJE4zqIUrVNj2ZLohH
GajfuRtHPa08KO+Rp87mqSE33Zh2eTxIaBlE+b0qHqWP0YBpT9djrev0P9ZdHGdS
bkz20BuF8i1+paY+0rKOv7bNP0ftTfcfwtYMtu0s7952gXgYVzayCmAHd8AVimyz
dRP/ePA5b5aqds9U4TQ83CcE2W3G/y78NQtCOSk58MGX+XThd5vCotGjTyWKVWW4
bqHKxIXB9aVsOp54HjodfTdAuNMfHd+muLLFksLg4ubQL3gKqSdC1mmgdYGjAkjM
Ulbz8KZ1HY2kHARAnCZCLW9mATMvFtLlP8893wO5aGf3pAbrCMo34QageoKISMwa
M+ehVMfC0NSVVvvuLVUqp8m+MSmgFhZDv6mEJycHxJ6fsCpbLh/NpheCGoF3BJkA
HRMRb0e9z45l6B4ZgA0SRB7Qnu4FnSPzePdG2epygB3/wjo9EkTXI4RT58ykyBNg
P4YxnzOMcvUBcae4E8yjBVOxzaTJaT62vuxy7wVWkrcBlUV3C+VDl0znba+Y1Inr
NekJSotFTIiqPgS/rofBiO/Si/5d/1NWeO23Fw3dp9IprAOisSx3xgIoCJUzLkWl
7ld//o5hz9eQU3E6cVwXoftoe/tcCNx6fukIMrHj7LipzqVhrsKLsZ2cuwc0pKgD
AHeeXAkRDtQTw119Ye1ZR84fIGYb7DxZkEnJmio03AyYLzc+P7+r876K54lUJj8l
DTNU6ppSdyogH6tLPIk06/MYQvySeSCwO8WtkOjep450psbJd0/6EsLybjiOGVZ8
jtKwCH1KZObpsX7PZ6lcnkF3IWVLV2G1HnM/xHtYIDRZtTPcdyffUleqR7QO/XH6
yPKKLFrIYAY6K9ucWe9OxewV6dWcXOFRPZ4IsjDItaB/KEwaa7VHzh/8Pcb40BK1
JRxjmroNMjuFowH7m/Fz2HCZI1fyNKwzogQX+HzrjOd4EOqucZeuwQOTFNRmK6Fw
sDVR+kBxaHNKxsZozqrmhYA2h8CHxKjsJmA8GlSNVYcWbGwfXk+uXRpLxwmgaRz5
ad0sOhbAKCVLVnorTUi8VC+oltgR0pTTkVDzOhTjPzHLtEmCrcwm5kFb1Zwd5g3R
HQuZaP1TR1JXtk51uINAhpszJTyi4dOixybAW0QKCWtc2V4UbM43e+dlUix3TyrP
kkKMng5e5I3QTT+UdZoVD0UKUT3LQ/khAErsj/LwCzse3jBwDMmn1ALrDTa24kjM
HIZQ+KRM0sQdcTjarDppX7yDIOeDMh9yq2W6ee1+LkCGbgmlcOcxwr6Pjnf2hoGQ
q4GDx89DRhgTSXmrk5xzxZRSCtJiwn/wyHbkiD07/hTtgl2XUxWlBh3TGlPbRbDi
hNyv+qrXhDipTvwKhqfuSEpKkgIzTaCfpsrlE2Xd9wtKjnmKkTGVOiN+EolUtvfB
0ibRRxga1jMzyQr0ubZqs6/IQ9livGz+rH39tHSZtcXNrNxEXptr26Pj/p5guwTt
xgszHm0Nf5ombvnV3CPK0ucnauBntVMuxC3PfADTJyWAh+49EPpdpxpVGTB49PLA
76f7Ko9oLgvRziLx48zhiRVtxh7qCG/ufgNEyfM2rikaxIcrd+kpbSrrel4aX/hL
2P89L/YpmUY4llz2axJ78w2M8PFpAMZ/oTF1Cw1D0YiIL1ZSIf8QsQ29OXjubzaw
CFO2IeAzBmlDccW3IUkJGxW0wFkEYeBBNw9M7rPStQUjicv1tX0jKZKLD0RfswUW
WBVsV69QItNW+++LtwfcS+MlUki8Z8WrHRlFTR7ysP1MRD5wmcGZPcZaJTvdDd5C
d2hbWhRvhuphVTVpANEvQU3nfmeR7bMXxRNNI/cpGq4pPBY9k4JtHXF3W+DKoLMV
5F7EGA+GDaaP/paDAVMj+6cCvfFTh14gXXihZJG9ZNB08DxiLGjPEitIz1VgY1jy
jMUMdCGAZEFC7CEXMIjqBUQCMySFhFc1+2e5NmsuQj57cho95W8DnogdWJqQZwiI
eZ4ByhcHSNSahcBUhMcNLZZKZfo/WmEYvUOCSzuv1xxN9rtekaQ5J0otUlInoyrW
ZQSbl541J7mdK24VWnZJiMt5ESB7t0Ay4ZLO3Bu8Rx83fb86c8owUZCJvGRewz5y
7Lt/OG1OJKjG2EwzhLNhfEFuz8fNV6zOm0/Dbyd+6zeGDmt9UfxvbC6xtNF6+yU4
539CGWka0gnhHGO43Prc23HjLyCKf/Nm4G4V8baj6/0SzlhRSTeL/NS63/8aYc+7
mQFg2o/TObeS+/5GoXqyeQrb/je554af5wlxjIUJOdXoRsA/nyeDPsZobL40GP2d
1c50eE6gyH8psmlw1s12IfV0pPVKp4UwOu5t7swTevvcI1K8W5QUFCmjujvKYPx6
yuEs3Z4GxgJ1haaYaETy2IzlbLRe/ekPbFlV/pm/115DE2KjLNBV37UA+WnZfCEI
tTgtwNqx8jy/P0/LWcfWblXKFENNkaaexfNoID9Jm140i+U0P6jVL5rXeC/xP9fw
YILhNmL+gmOYJ5EtUKRp7hftfbtPWbAXpVF2F9kEPe8rdxQbZDNM3H/VuuHPeUdb
A9eIdXr/5UWrwkClMqpMItFABoeG2ka7fsIxOphdary31SceEKWGja481qYp7c1M
M1+ciwjrHKKznZMYTL7ai98xRPRa2mk5CGL+pzIPz08akJL1ScxaVXjn/ixi7RtS
n8FG8ycfGrRUOpAgRbVjnqEwJfN6KANlfATsB70bhgh2+tMuXCxMNBpmGvO7Olbx
hx5smdh96npCwf8lseNtBIgOM4glz80US1WaOlSLykaXZvtK9dpRj3BcBUV8ElSG
0TuzNZl896pOgXHRvgzAIwU4D+LsVontSVNS7vrcoA8QT15TcNayFhR0t4Xg5L4P
EsEZv2zhHFQZcezMP8/mqlySt4bZ2l9RiariY4Bqr6ohQDyuSNSTwtgH7I7iHJNK
ywIXj4+BeI1TzWKSYOdGq9epKmKhV0zcvqJpgfTtH6+KPOMAJ7dvHTeSCvNEedMO
oT0SzIFkj6z3SjEYJyTgkv18OV+wqUWhfQjEeAmGmLkUdVH+lsvfk4WoFqC/tgF+
ECiQw2ERRe+ycA6UKTRR0QLJamXxAYLXW97HO8qtchrEjeDzf5qncFFo9ZRrq3dk
rU6zBukTojSC/nhTcFtg6YbOLv+FhFNmIPYxMx5erl2TGnR5zevT5poX038bk4Dr
OIUpUJMq8D6+iIKpRWEAF88aDxLZARtdCI9ndeXL2wr6O6TJKQu4/o1MHr/SnStu
gu8Ex8h+W7uUCjBN7r2mi/YcrgFkY0dsf/h7tZZ6u+85zKYr1KfvPbDg/4WfvGdX
VhtelHCSwIvPy8wxbb7mlBDGkBUXUxzsgM1eo2oZ/V105werP1VqrbTySRfIAAVZ
sYwKsK2KRO9T6SXB9SbMsCgPgPbZUaUopONvZz/0kSqJMnZ6Uctw0x1/sl8Smg13
keBSW9Svn9tuBf+KNQvPiit/ekaS+ESUq+VW76lIe5aASxjVcHAFtg5eWVOKIefn
BZ/njATdjTf+bG89nxfNu3J2SybJeTW1z10BP9Mha1LdeObcYqBo/QOQ6zLNgv6N
R/8wkP0Z1sFzyuLHepvpIggAt014CRz09HgeGGUqK10JW5hsEw7b1Kn9TTg1opbK
XRtfXjMFpfwOlvBvVtX06NpO/0TGXvRNTzYnOAE7KQE//dJZgHx0Ui7d0wJJ8g5u
QnucWyYJSQnrPuZh22FEmtkPs1h0DnzaDLlba1wSQxViutbYrjYFic5nD8EQK5Lp
dBUIrcvAc14eUa5yWndxS9FNpajEphqQX+QkonrA0u2pdPW5QVRwAZjqFaSN6aLH
OqorChGposmGHgyUzV58AqJFzelRATfJ3Is5cQpZRmJr7xgi22ayYIfTFLUno8Jr
7Doe4sBlXZjPGeL5L2vwEckX2qvXGGwlEyBKF+cs59SJhdV5WIcGrSJcZ3N7K0xt
MPFSYMcNiXCGuis8kRzDoMEzM666tQE4BaVGDWTeM0A+/9644OTAQbCiDt83bIxD
j2GEMF8/eyq8zCP2sLCvCzNQox7gfKgLWp/RjQnlhqsXphoBpO7iK+snJYUYVDs5
Ra2lH/b8FIoExY2Wqtda/a9tU5urTcbOT1NJjuy8CrGT6QXbBD6HUWNKKAYLBWju
qYxs+i3YNz49VzkP/jlfQ2rGOWqFUfkS1HUYdYvhUjN0mtaTK1sUgEwjdi+Jpuk+
qG6Zv4FsJflIspVhToo98NVYlv1bHVxn23QBxuP3VASEn2l7ZeoHF4avBfpm5u+6
eoKMaauvLIUCgCVv2khrYED64mWMDqAa0wPQbzM4OVFNTGY1afi444ansTwMHYPY
Vhy5aEseRn9EtdGyq0EoPTu+NBAvXtrJHUUOoDdrFDq8PvbgtD5t6u2LmLrUzbk+
189mwYd3GauuHurcXWJKZHnLCxEEGhCPmlkMCIsZE1j2tZ7CbAMWtxkCo7bZIttG
U6JXPK5sJGn0NgQPV87DWcbsvhZ4svczxy2erzGK5qhJZ1M8ThV/Hc8ncgvopLS2
69qZRZ/zBo/Gl1IzjatHjoBYHpaezA62NuohqI4/0pQQI4zTbQOqyeSEmbSlEA8+
/4eFRmFlJxe3kS+XYIu6EvnOM+vSmE8Tbx5VpODg+osDTVMiB1cVmKVniuWy6uIW
ZTx5EOMSgRfWBIsYvQwew68aWc+mM8/i03+tvpK/J9EL0CHMqk5v3KLmM6QAgeIb
FEqVMgDlfSYFU9+IWIJnFeuBDyXFIXKep1TspHG/MLRofx9QAck2ln6JjQKBKkva
0ZKCvb953AUFtIyqV6ByKH2odVZ7KBJ4psnkAy0/AdRNPBaXsRMx7lj1Qmo9Nj/F
/dcFYTaENZW8AlZyXz8QCjg/8CvBFhVgfTibFLc+q04EfUnKhOxSTuEARZdaYahI
AdyUNTFBC86Db5yyZUmz49/l7n4esBAhzWXjx/AGcmkKlek3p+80wMae/wxOHR6M
bGtc/dBtAAF776Xo4+jHnQmMsgOMCtUNzqadeql/USzazuAP5zheTQNyClicEJG2
5Y5gbsVckc8dJSJ+536E0epD9Z9Pcm74J/W/SAAtNb+Pvbq9xuXF3qFpounCVHNL
M8BZ5sI15N+tcoNmiwsMkEdUDvOeX2NBreavknLgXLlzYKbsEHb8zjy59ajD/kPK
maz69ch3ilHbVefeGbcs+ML0E40bAWf3hdzwksy4HMt30UD6A19OVYFrkJnEtWR2
Dn5fysys92TH5RwhWTlGZcJFGs+WyL/qeR8OMrpnJlVql8cMCYPg+PH9S/np0eQ5
23IAIelsj9TkdOUPxLEsPPNpAm1isAI+JNkaAkcC1wcFSsfb/jePBGiCYns5fnCv
7DvAarnTw7xiewm4vyJTOjwPEQEeWfOaiXtROud8oom/5lGLLVbvDYHu7r9rK+6D
VhOJ+fzRA46aanDD3Bce7IpdNUZrFkKBpb7uwNTIKhPNbijFQNbJGZz39onT+p4k
2Nl4iQ9ztEiMUlRVzuedgIeRty1BMpvjnOow1+OPx0HcsbhJT6aGW6Qf5ymxE+hN
Qq0jTqpWIUiW0m4uYwN42PM0vmd1nfcjxg77gO5SAmhB0EoWsQuAl156C31307AN
OBh50OgQFtyf4yFFeKjwTREheyvlg/VE90dqoa7ENSPZ5/btla17Ojzpkg2rqK3W
bSsFy9EVJmwDvdtzeAObA5/a+fwwkffdG3roR3PdkkFDGXM2EuE4atlmIn4XmEYd
72IHdplm6v6MCA4eec/fu4DhO4lf8XrwmNHEVZyhYZMaj9dDEhrHqM/K6T+jGTYR
HLN8H9e/U0E7ivQUbAFGYueTeOizgAiNB3Ti/GwsIrlWUZpjUUnc2UHLferAjf+8
krJHLozd3nD7TxI3Ks2UKsRBszrXmkaUBni/Duelcc8yYKjScA64T/HTf/Tj5s/W
cm5zzGzKNd8hSpHwVy+0zOgKgUUPRdBcV4Jk4jI4O5YEHdJsns8piui+f3qTxYri
3toow9cN/JVw+p9mKxWakjJSly32m0Gj70QJG/TtwuFRoBMS1acvbKRd74jMdw5X
5CL02FxKHkxN5V6PNx8oojB7kRTB0mU1WDu/uuNB+Lg=
`protect END_PROTECTED
