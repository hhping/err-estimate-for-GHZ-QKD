`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DwJOmZ1gQZXr4gqX8tPVewg9u1s+c29htNtQuilxLOhD2lBaU8HBo1ZnnD2UKcsb
MJC5ZyktmeIQ6mpSzvS7FwMQ1KFzVUms4MzHOFenYhtcBTfRMo3daGxbDhYKwB4d
q3yIFm0xYRMwdupDZDerH8ihMsQk3T43fo7AnnscddbwuxRJoT/m2dn6yantqKze
E/nf3VCJeGfs9ZztUll3bISMe72OJsqLqpuudToyKTH2c2c44SrdGSHiBbCaJLac
GIXCKH/9wzmgyn62nRsEk4aG6wQ/IipBBKYfTQ6pnDK/eNDdHLdd6bQWlwG/Rd1n
1FhOIkkeux0MLit+MAWcRYSWwy+zFuvnPxc1AlA5GPb9Y7wfwDxgm7sYVSd3Ak5T
0XleSJ478p3/+unbZDViNWuzq7Dc9TSF8ASTC2+iv2+ry4MMa50RhQdOPgMm22u/
f2ZmL9c5caARZl9h3U1e8DNQIQN7X7i8xWupvRu7xlToZcuBMHsffRwIJeiP+Uft
E+sNvdL4PtfrQzQyywnM7MKErsBDOD8LB+6Qstdhy79lJ57ActBF5T3lBsHoxate
XypNa6HRMPU4ClTDYJ7KBbFfCDvpLUSjXtjIfJeCtEMLq6KOghNOspI7Qe17QwQ5
R7V6090NV35GPZkhfMRKcZ7+yzlxQfWN4OUFxa18GJbiTcYVk86Djfs/D/3ycMl/
7e3Vn2+HTt6O9oOU2pLwVbEql3Webl0QUl55vdF5AsDLwyiwcQ5cukswLKEfqmQd
fvol5Fy0E8JiLKzHl0Gasnd2GaP1bnM1JQA6lVlIU+ZlPs0jzRtNel+IhLHE+CLV
8eqd/c1FkXoDR4SafPF3eGrFyxm5La/izeLcLg+qmU8lMMKLRYIZMGbmYBMDZ4Tm
GtZLziua8PDIEx3BOe89dpGND9jcAfsPMd4U5G8SNY6mEESITXYOVxXbELaTuXyL
tc2O4U6r1vVW7/BffErkSuKYBnz31fcxH5V8Cu9KIIt89bOGXDtFS+PD49yeMgPF
6jG6i6qeEzAqdW5lIur5RTmB09zSAVDzGDEJG8BXSD/90vxDCh34CuRZ9ufFvxOV
PV+onwsA36GjrGPWFAtLfR6+HSX+P6IrKxSIVItHdfWA0zelxKjEEFTLg1zP7gLO
xEY5ikL9UhXwi8lZqmwD4TtpaoqA7iQEPMiPOp7zInyvEUnk+2cO2tvh+CIwnvAS
FXM0br0DdyQVK7JN5CtpZhR6GdpeLBn1Kki1Tmkwuno8eTuqHQMer5i6aKPcqd1W
6E4OTN+Q+xtkgs1P3y+6ozjqlzHB06LF9/2SIGUPUkoqPbangCIcHbLQBhbQI8a7
YVWk2QiHgDCPgOnvbxP56uiAalvM+htvQJJvBbKwK4+I+pXzQoiGMft8jCZ5LsJo
UsjzBIMBcJqCc7dc/cW9qVtBfKoM2y3hmsxqHWyeZeDcSSQyu8rzr+TrK5mkHKdb
yIjbbf/NlvhwDxALQRaiBkgljbVqZn3IxU6m/FjjbdEDnucESYJkxgN5WRQt6kzS
HpWnopVIr5BsFpMaHHkQAg==
`protect END_PROTECTED
