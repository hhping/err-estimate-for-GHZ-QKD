`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YiDuVmoYWRymLyFqZhZgtjhcZ2taFvybyRBs6ot8N8nzXrorln64hI9mGhUIkzwh
g+8jcaj/KCceYUkL7mrZnoM8TLlAmGFUAUNhHb94Y8BBerOEDJAhTBCZlwfXmx8r
k33K0fE8ssl5O8gqYmSebJZur6+zBn07qRpRuzTls9Ms9BH0ZNY8LU7Rn2CkEQHv
SqrUW6AzwyhrkL3OGE6KImxnu1ZXPD0Ky1QZrNLqj4EMtYcB3Xxgse+XniVZHy/d
Ip3kzNKHMsEJJjlKEUFcseZN/wnSyvZ1bslfbwBzn6hxolMFa2oXN7qheQW0BpUq
iDy9IGOCwtpN7Bp4tbXNEmVOKUZFSz8mqCNpZevIG56sD2Jac3WxQudSxG9cl+Kk
IJJ8GyJWExHr9w3s/YlxWyegpsaJ0/RLbvC4+oW9q3Nj4dV/oqJqz4gfWm1HM9Df
00qS3Kh+ilPsUMynWRHlKyDzgPo1e8LT0UPlXtZsE4WzeDJ+pOgZLZU5wwjpaRxc
IeudAZnq3q7/fpVymkQ56RUH2a2uWf8FKRtmfJ4mC2mBlC3w19wv03Ni1UkKyyyl
QMapGuXAPbumZZUijyXTxTgE0fwuIHcxWHC6H9faRGsqqVNN8z4Tg3Bq34s8qcsO
P5LBDaMKUVSxNUF7nAoJAAb+dZYwFG22sPQoseLg2DxiYNE/Y9NzvaGuGuNLdYj1
XbHTzJKSTnh0y7PQVTFpHcS6YQ9YMykNTC2Z2C9HZK5H+Z9gW9vPyw1SxJjq7r/N
iVmTWeXn1FQCYfTAt+CKIGwEKosFW46wSU0qSL8xevMR+4ALZUXtSUJO7ViY7iGV
GkqgoEIqy3s6OAa0xaEjMg==
`protect END_PROTECTED
