`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6KTNvtH2hu6Ahz5Z8eBDht/xEEK2lcuKgOLUjFwDKCQ9AzI3TdjgUFPfsL31u9H
WPoKfc/2NYFIzXHzfnU0n+W7ZnUvs/IoiRZMUzcLUK7A9Yn5jziHjKRHLamY0f5v
KEDBW0QE9S4aYb33pH/L47gY1s0mJX2ggXUsG/xSIlIKhKXBPKNQd9FbI3/XLrJD
CdP+8wWUhpW5Pa1MybREgdJmKwsoa71jKRYwUZbVHs6oaSjibkayfzzjxqRRAH1E
lGd+8gbXomQrqv2s/xHHJa3gXygjeGidKK/GKOEW7EfucG7MeuJXaZBbQPEi2o1z
87ixsFC37RhJ6M/HAatwmLykCg5sA7wfsNV10JdyBj5GOESLDVRW2R/+LAyODnTi
cOiYMKaCf0+YfSdNl4aOYtqCvNWxLTjO4fXiwnw0ZHfuzS8dkTSS8q5jU7wpFKwh
`protect END_PROTECTED
