`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ez/KqFdky/6TEkiU0ZmKWlpmEe7Tbtft0YAVRwgurSy6eEBD0xkIQznnHVAdYJJN
1kE74XzhYuMP/XJJ8EpsfZ7UUydhTsATihF2fezQcc7EGQVyLTorZm0WSL29MwmH
y2uTi3Bv8E40IfKBtmXEElzgIMxkqDB/eNPVBMtFSA2Jp4aOHSaNIRkpNkZ+5d73
GvHuVZeuemY1szLnTlS3NAIZQ9nqS2BphQ6TvWnpXr7W6nmkqxrUVPpwuODDFYrl
xS3eXuknuhWTTheVMFkIV+Y29gp3qTlXizP74kna9f/fWp16RQJvVdw580SjfvhE
dRKsQbx5kX93jRW98d2r+iXThU0nYHoCscszgFaV4VzFGi0qQIPK4AWl6WRy4am9
P7M5uJ7f7mI6NPU7R1oLQ8DlRoQnyXdi6Hi/KGpTlHq/VAgMTLPRdVx0RWXkP0j9
YZwwf/tTc5fH5gYexI6zvn/4gLU3EQGeuiROcVqRJvF/xYOYX+tWGBevYpkjwX3l
i2Cwk4Wll+TO7AoSRNCmIzbE5yBLxburh7LypLY66t6cP/b+A8bfBNzkV7dtoSAL
8/u9Bv0BbrO2N3qpO8Ca+hC7H4khOgOsh5ql3feBnZWGdmr9w1LVwWunUd+PLrbC
gvHf8fgOue0onKE6uOvwfXaGWtQzcm2k5dQ3i4SnSliYggcq5xVxHqdbc8JxoNS+
HUopW+rIumJkDavc1XSBoOaBU63XHU8RfDUI/TWjQ7P3Qp9JQjaki+JDiToh04ad
B9ELDZsmjS7zjq5WxxNwCCqlbuVjhxogO841JF695FaO0xqCgD7Td+7tGbG7d+lm
FpHsYEubd02zNCyZx35dyLZ9K7UA0CXRS48g3PjR5p6U/+qVdd4Ou56DVVAEp79+
RaWWY8OPljw9HOOSW6LDrwH9oiOLPR90jECswbSK8UPGjWAx5p6KyKDp64z2Rs/l
c4bIPEsLvSZ93Glqn0R/7cyyRpUmveW6h8pARyOdy9gXD1Xkq9fYViI1JbmdFuDq
`protect END_PROTECTED
