`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OolDRaccUrfQEvWjlde1K6V00DAc81m6zONYias4XTuFEzVaW2y5SuMXWcj6NytK
cN7iC88a8ZFw0BNll/hbSXB0rC+Dk8k8RrYp8pycNZDnjjxM6JiSzeg01+mZPfg2
o2m/z7dhhx2TyXYr6uZdKhIDk/kB1zcJw/3rDQCULol/c/GRtAqFOWQhFXXQy5xZ
2qXbmpGCvbRzE8OfmqOpu59R95VIwZdfrFrodM7laT1M3ejaNf0bZTxf4uBZ8tv/
wjm7j7izy1idVvuPrsN9zUsRSgqgsmeFCd9/3U1aBxKyiAp/e6vrwuHNNKsKrp+y
h2FDkNgdpcF2+D3IbmF2mYOGk+euM6mGVWptspVnuIU6HxRQmTt8NJIYyoNp/Tl3
xBh02k4AP2PY5lkTV4W13FBWIVHgOfPRCOrXpktVX8Tjrd6U9qgTnR1ci1Aoeted
L/rSDrTaWidHJw7k/oZqvAAe9lDkg/MlpoXm9x2qvtpPymHjVpaCwmmRppp8PYzi
jC8OwfC3rM6n3UkXYOOTUTHSffFm4SXZZiwzMplD1AcvlXEc1FrFt7WmAQcjcn8a
MNU+hmgt93wxF7l8j4ayWd0uvJc/yTYPgawujp1k6j/4DKHSmP4W4K/ZwAJ2/N5t
CWIzIctM6lcP7lLWA2GljrcTGY7rcVKOk7OHVc7pWZXE9240o+zMtWg3l+lUaa2q
CF9aHThpuqfRBRbVUCtpuxfvPg2Ca5lm72Hkc5fEl8sGgJitnSOAyauDYMcOcWrH
SlqcCm/bC+h1+lK8EZVp0VJPhygNXLkxu+9xyqEgbwZkeyoS5OaPQC2xLHrft9+k
dAZlbSou4//1sqhZ+TDRvLagtLYff8zVsW7nxXMF5l0nmKBdzw2K+8OujIMOvF4T
co3zQ1WLIaqzQdGiv9Ng01MlSqraS1ZPu0LVHG5OdRnMIj0t38HzIrH0eZS6wgdT
EZzAqXwx/0/VoUbuuR4YOPxJMQGjwHxA3ZVoDatbHs9XT9ISbRG5gex1T6in5oAe
5QOPC1ndoB8mh0R36EF1zR3BFPJvc8WjYqf/RP82MDjGf5Lv8DkJGzJgn0ctfu7R
xShF+rOBumSvBK6dB5VTvsokntiUCflE+Q/soUh74ZQ1CsBOo8isJTeick6vFfIT
R7SpLX7BosRFCVn3GBegHEhhAkCdT0bozk71huY2FFN9+PLdBbXO2MRCZ3+cdSCI
rkSPYUY8Ytlg+elG8qTFfTlISKmCH92xQQwjQxETCPrsdwAwvSJdrJdjc8U1NNy0
FkJ2kTKepksiTZivpeuIC0+CRjCWUTOTiPmKlY9dfpZ+Lyc0YC4NBAUfEi5GfCXQ
`protect END_PROTECTED
