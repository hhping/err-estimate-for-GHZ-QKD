`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzmQoVCkU7aT9/aRPgnnCM6KVJe+cl3KZYTnPHb99Fzs6rB/xxaxFYEtDmSPCL5U
F9iUAtf8ZkhHyu8+RZy6J0FC+Z0xeAhanSSoD81SpOqZ4h5cd3Z5paKjjOjeM42+
tuyvNuyIuBoOSnnZaQnTedsi0HkCc4hrBOZ3/5WyfoKX/pv4uwMZBQO+ubuCWCdM
K8Dj0ICsdHmvNzWdpHb03SObUwR61USDe2H2DDdCQbQZFAyYl+Zoowpp5M4r9qtz
iej9mg2MP+OorwhWbH05QhedrEueuTqLyzClJozQz4oaGzrUJC3bcRNmwwCTa7+b
LHRDVom9f080GkdVa21ITUNKwLziOOlhC/+yEwBtUaWqC5CK7Cqahp2j6+yF9THX
VjcnoAjV2TgBrCmdtOLCkC7nK6vNmYQTLK8a4Ww00sGuK0Iqn8k63AXN2BkTDix8
Ja/skS7gQYKQL3rtZfO2sH2+oWbVK9lqoAI7eHjOm+yuS7GL+68ociOBSP8GScSe
RHDbFG6zmGdnw2l+TA3KUu2fUrIXUYu1oga3qh3nUwbdfBUj3fxAV2L9GzoM9CBL
q1mY3fURnpQajpf+ZfFesO8TRqZCzZ/HOmBeWbFB8zLglscSkKZxtOijTjwb2pBQ
HCwe9k8spkuNi4amvJagWBxEu42wPA9M5z1Ncv9Wtzq0zDRvj4Ec/adAI/8u53PG
JJelLMmvpLp0dsX0PU9+J+MaUODkzeFJXsc/u8lVgYDP2TT909FZ3UuTjEfQI7LA
Vwljm0PCL6Z3lg0tGs9YKbfTvtvoj6TnK0JI7AngPUPNiBZxU+dirojmXKAe3Pfw
VCULM918IlkXVcVY2MGi86ukVlB9Bli7ucfHwHszVNUcm3tsfGRE8SwuYSUqVaIu
oX8lsCiPOhIoyluO3buMnugT63QbPH23S1ulaI78pVIYN46sqdgAT4BrwyqXvy+V
3HK6V6yP4ys2a5bm+Qdw0Ro36r+PE5zrAcB+3sapuulfmYnHHvJz2/z3+U6bg8pW
nOMAO9E+rMuAuEWxoQawxlZtrr6Nu/fnLqCfHYryteZBVYkvWDeTvBUU5UCERNNM
RWyp9BK94bLR+03Jq0iTGgaEQ2BjBbYnS8g8N+KQBS92qJM7Ez9v+F26SxpaczzM
UK6ICwT3cf0cDHhOzMg1Ktf7JZSULtAx6enSK1M68Ol6dzmu6bqm+ljldOc7EwuE
d/515i/g0sOFV3rg2auP36fDItnzGLHQxEeljDOb0SUpNDHWeDsAVmWv3kdRug7H
ROZeG/aVh2fAwxrupcobI2eVoXc4FU0bNNC6+nIeyDEiMz5w1OYN0QZAHzIWablU
sMQlW4ZluqdtoKCXB2QIZ1TxiLteZ1g1qM8hlqWJhB2zu2WJlI5C3axAY4wJQDoR
GV8zhlQ89fgvRwnJzgCz0mVUS6G/5h0sADW7Xel+wMZJ8C1UnVTV1Gcvylzq2Zy0
ga7TLn9DEwRjH0LSbzPcvSm44rFoQA2cm29AiHyYLn5g0pezqTBWkHDkt/AewTW4
/rbP5aFi3RZjCGtXiC6zeykRAgwJCO6ton43Qmb/7n7W6i+mC44vMwdSMEV04tkk
0pm6fyCEAk0SFArPeaTCbmR+BH4Z6ElRQKd/0a9ZRTaUoA+SZRtIQ902HRMd63aH
TECcEauLZKEKKEu1P6LHLnAyAL0jqEszaKB2bmXB/H6IhvXXW0cjW3iAKUYFJj1h
`protect END_PROTECTED
