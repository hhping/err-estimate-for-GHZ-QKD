`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zr9+ToriKrH+pLOQ4kBNFV6AZvRwhn31BuDNfJderSJQqMeMy1MOucI7+M3TNto
EWwR32nUbVbq+dvGb1qW/Li2MgMwv9WsW9MtTBGL0zUOeNbXbhsBQOARF58YwZiR
G0fMH7yW3g03sIEcXKO3BJaJi44Yka9TssZcDlFIJy2uag6v+lG/jmA/alUMYnKf
YBQEbH4ydUl+ADt7o7BvUl1PKkoRt7bOkczTNKYF1fvm9Mu2EPCTnX68VMiVtYWl
S/Gt+afd3QZSQqeSSI/QU2CCRWXkcz+Rxe1pfbcWsCfFDxBq9hSh7t917Q2iGKYc
H2EaMbrKzEI7UGkO2VILplV5yItT3RyMsDe/B7FTeRHejbXLkarjfga3TqLDk/ua
tSLSvIh7t+eT37eUIF8tc5W3jHFFXCqUF4gR78SmcrI12Ih0gpxcjcKyrlnijH3J
HNPURaJU6pD8jw5Xc6LxNUz9QxIxSjnjdmHrlR/JO8B2dOXWEFeYWrQMAizBrNlq
4m1ZyXNzdqg/ieOnFn/DCZUPQJojDWR1IPs5B9+Zlwc1BskQx+Q2xOC3fmDG1/zq
9zcKEqneBE2j1iqnUALve3GUyslt+tz+Q5udRa9WZBso0OazIOaSRzEfrXB/UhVs
xAI8z1b07zvgh9TBVefyOVm1EjOfkEX5aU3b7DXoCIgJkLdymg66NkPhczxnCSjx
qF62cjcfrdKOImUDZGlAcOCHygUszeQw5e1nSehMro9OFSx4ZabTIWt6+iEbHtcR
46f9cRrCCtkdHxX05zUcXNRDtCW8j1ayB1S2Q5/uspGxzagu7Pw4d40XiKeTowyf
Awrr+/RqcnV87VxTJfbsIyMQcB4pCxffZTJIMSXD0bCctz/viTCBFJJVVMp9l2rg
oZFeCINixjWbVTeaw6fUnifheENbqNVmUj7zkyrfio+UVY1bfFpFhCBMr9lT5BQg
vVxGElakACDgGVeFNVhtAMyh3C2Y1IeqdcoAHhNpIW/CSLzi9cDAAL6d0UcpZVqk
8nNeVwTT20udvAo89+zDIuBnf278hs3Q0xVBEwDohcihOjaBQV9K2oSFGXEebxIY
JZw1rAOtaZsbb6i8PnLIp57d7va2zzFQO1QrulThZm3aWqFATr0EkSUGaG4ZfPev
Gm7vqsvp4MFblp4YB8NvkhXsOBrtHa0BXDq6+Xaadpz+82hfFHGubo3URG6c7LGD
vyZEHKktres73jCcHDD6XizAWwEVDP7uT5hmShEz+8bFclQ+UJpIpKKiFjUbEPbF
ZNFWvFxn0aS3xIjXjLUsaQ==
`protect END_PROTECTED
