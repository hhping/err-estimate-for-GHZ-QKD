`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Bd8VLXAmVLHwIaQUBU7DO9mTy5PQpMDNWopPQMk3gYBd2paomRPXOaPOhHdqRw5
vHFVbdTY7CL/ycBrGdXOfIyZlyCl+tCPmU4kigdPE32LGgiD8k92+VD425J0m7ph
/vbRUCOINX78J0ibTfjvX6jKZJ1W6HDoBZSCUHHvo0lAvbzyY0oocT9GPhIu2ImP
dgdBFGzATuH7cidpfp+aSmIALC7ylxWlU+8AKxuUB/nfCepP+6I9yhHJS7mGbkRp
AivbaXYPvR9lz2Rey/KzrkoM/JdOo8A6YU4GuAvhzTynr38MTCWiR4KKnOoujxgB
dvoB4k28WPGsjhEedTJGTBhhumL1VVbHUGqiRfmExkRg7eOh2p45KaTnuDIxTaV5
izfeXSNyevRMoYQhYA7xS2aITSEkMAntipDdgvk8AX91RhLuVbw6IcWrmF53gyGW
8N1wvmkadnafY9GS+vQzJhbcXCVUxzdNz7smYFohumJ9Y4r5WC4zU4rO9h6G1iAq
5YQrrcpKH7pQrebVDlBz0NQKZhXbbtaclIZfWuSQ51pUJuqm7mf/SEXVg3vvcxCI
s6iEm/8/C1RU/WwfJoqv8zwMA/r3Unw9YtK8sqsx2RXxLopru9ftS2nRiDekWpoM
nP2nfH8pRFgjm37pu+hscrhV8CmL1MNL9zVEj7kyUfOKdsRocFB3JtXMRKO4uozw
rkKlSXgo5K7lRNyqwSXRITFIPorS+iwwqWwQEsEbOVsLSappvfoprKT6Oh1SeeXe
X9CbEm4+UncxHR9syMYagZjYlwsekpN0t2bOZVeRdkcktccvuH2PC2jMDqk9n8EF
VBIE4/vjPWGEyHp0UmYIMLFLAoQLNSSh9DsFHAhOmOxY6BCBN5902nOk4nFlsRER
LDTwoVD4/pBKST9+owI5llmap4C/rGiGkJqwWyPv4jtT0/2AkZGlZ+x9cTQ+kvGF
zi/8sTue2XMeP5r0UqnDNI7a9h2TV0fBznv2icRUwT1oqcwQyfxoort/H8oN+LqE
`protect END_PROTECTED
