`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CfIkUekslQrkd02cm9J1R7BltHsjXMLvAj83DzIbab5CmciVLOOVFFoSQ1jYnQaO
SyL78DYS4hT6Q139Y1U1k3rkg4vD5TC3wjw7+0XasJQt7ueyWCFOyWX9ILx+bbbn
If60ZhoAtq1HvohwvL9RhGQDR2N9ShLchMmrUYVxbZe5o0Yw+5ycbHIQxi9V0D2f
V/Qfe7mAXgPU79YmUT4N7cSGnYLPD1++SlRrQ1H6eGsV2bGm92NBpgCYoB73eFah
yRChL3/xiQDsJhKVc1dTuc8SBkIh1W/p3dfV8kMsX5E/RBO8e3KldO2JRnlm4N7Z
0jSYJdSlHbn7LYoI5v1TwPUZ5tTE36jNS/gc5hG8SWEw+n8UUdu2lYnVqWSwtDDF
DFUBdf3Hv/lblz3ySQtjTPz/Yt0x+lpxMeX11wQfVgvia5YgaUclbC5sMe6G5gSi
0PjVuFLTP4wxgO6RVZzOk7jfYUwk6nj9nlgfLc3HTE8hGAThOI4fPG3+WMorH8YW
0TJvSpaTm99Kqcki3CL9JuZTZR+7al9gmSaFhiqmVDct4TojWfuwD+D4+Cy53iBS
6+qhv/PMDgpyFL8SBvCtsJsLYTMpTTAprRvnByqxdYwnqmxwEOp4IY7XJo6HlIlG
oxxYatwSFV3BLT3uBmGs7AXx+R3fO/w7taDWAVa/8kAMd77i9HCe0YtNSHHWBbxE
U+l/2SteAwiEEzcoTK0xfml5Rvz846sVvUZpbYIlX+axCyp0yi4zuTru5bSUDzpN
kQh1pVf0k4msA/4+r4JBzpsHksno2QbN0wEuA6ny/vCuAwEJQTClJ7FIjhyJRqzx
mx8utDd6YyY9rNZXqVYHvyjWk3Alhuu5vE5CGe/XArB6ltg5oMPTEWN2iR2/pCEL
FHn8JqNWQ82aA15UKod4YZJYo7HdS3LXrqKeyffAyYiM+YD6EXI8FqH5Sn3kUTKU
GCz31APRspEFeD7nVWsg8sfYsso9TWCmsM8Q3aahdLlADM+sQLKxoNbjnL8cSxTp
WBAm+H9Wqs7IbM4zRCpjx73uc267QJwzljzn9Ix56+lWblby5UEczIGmuxtwAR4R
B2zBVbCbVOBIbmnxcKG8OTg51LfR+xsFFe3nFoGHsIfydddxpoSFuJQqn2ZIuda4
ftTVOBE3eWEx33ry+T5XSHeRb6b+r/RrrMuP87gjK97E25dK7hPH2HDpT+odXCMP
HnWk9tveixHcMjGcT9h6pcKJKYkurJUbn3Aklsn4E9Wo5eBsBoaEyLVOrHDiGPN9
4cTqh4pkn1H6SF+1/GZ+rr8NuB6AJeRPgxf7NBOrKhTlY3OjST5kLia0imHyJnzQ
7hlVXI5WXky55nbZ+6AxJnOr/g88GocCWKuWe5kT/ZK90UO7UVlyFRp/j55qn25A
YDj3oYFk1q3rUadIysHAPtEQY/HvMDJFF20CtbSbsQxP15QA5fJZ/4+68K8odICl
BZ9tJkA/oJmzaOCZqY6uvNRWyWBWOuX5F1b4eG8O9KNgto5YQmY0hHCsfUKzkj4c
MfZmOyH6/3t6fkfQUweERg==
`protect END_PROTECTED
