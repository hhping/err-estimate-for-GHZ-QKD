`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+j538WrzweB0Zp9nLrq/VssrwIQjSDvL1jzByZVd8LIzuUXXqOoYmFrAWoT8IHYz
OxDrhoG1hoM+T6zymiJoGEUGD9qh5t6uECb2Bo4wQKOACYQXfaoUYtgJf+DMxfBz
m0zJUH1moNSeH9TEZAzRsBQgCSZPDlnq05YtVXhQz2fdyhBwWm7l/2O+RiURIVAH
WJPdcMPDc3v/L5ZuMu6VBlpAIKtBjOEN59DvjbJ4DOCf9V3ZN0R0APm2utAxyqSV
T/jwORz/YQNIXyeBHJGJbCz2RQ4tBV/YvY1VPJ88lQJbkn8Yc6BvehIDfkZTpdjU
rFY8Cmvv+0RnQ1D2Omy7mH94TqnQjEi2ojiSk/Hx7xe2+EnpIik8h27krmIsCbHL
H6Jo1ID4fZW74QEaQhSpnkPEssSKpw0G8FQBF6bIyUIKIWcVy0zLKnBbrWzcmsk5
5NdX1nxjNMFEkZuR7381YbhWt+BAFEXli3gGWbsYh4NVokO3K+xZfctuI/TLl0wF
1ChOQxahyj+RCbubnVnuOoRCBfqDaYceLn0YNXs7yiBjzrtfh+K6ZuwOCt3x17OJ
v1Gp4O+fNWOs6nZw8fBpS14QAkW5+YLMY2TBb8DXZzyBqqcfav5GRG9Snx2i8tLz
sITowK2zHURghRPmRFC2BwBZ9dVTloAkJp6F2uadUpg40UZZ1FKOAP44u+RFDicX
eeWfWaHTSy25QijjgQzDB+6ZuS+rQsnKs0+sYTVjVA//DmiENwZYGY4KmCnL1i9g
UTFP97RzifmEASppv9sOiVcuVzjKZ741O7s9ZRBjxnLCyNaCgrqv1GIFJxDRriF6
KEWmULZdRutZh1sCyND44vgSAN/orNGwwZuzLUo+3N1O9sznzqMSrzhuWeMKsSru
UljDJvFaX60pBWNdrr0j5w==
`protect END_PROTECTED
