`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuLVdfwZVGQjFYtiIIpw38n9boCn8/6cdGThQrTS3EuUBAMwbHfR7omBORBvZVnB
nsS143FH+cf1eh3AWi5uAmoyLx59huS0IlSzTGBqM5tXWH1FUAk7krFSYruF4lpc
DYwAdYtTn4DwCmPxw3amLXtxU30khN3C+ye8Yc91H7F3tWzm001HFF3KVDkAOZwR
HK5k+CaZtrwh9MMtDtIh/jCUPhcoudDFUxyL9sslCAGyselAFCv9/pc1i/ZbzBrY
3jdx/7t5rmjbAmLQexbIK4B+G7dOVyO7Cyx5h/UN+7dXI/sycujasVMLyJnYnM8A
426pwCW/eMCO15p4fZSZCemcywW3WRrmVbaK6rfla5LnLippQomFq1/OZgSScm16
dHqS90kGv0EWTjL3xo/FLw==
`protect END_PROTECTED
