`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBaSOvRHSDGEiBJsNA5yorCDXDoSjEzCbIhM1fKw0aXB0xhJZGn1gBAdMu1JSzvp
ejsn3pWWWHT4TmS35kdOb+23VdWfknBY7X0Ku3cHFewrlx/QjlC1Tk9+PfG+fytu
PGjrStYHkHjbOcQ7i7AuGW0MELEfpo8gDXcgUizkMwo8ND/XFQWlB9rziZ4G78ur
6+LRVFy8SPPux0K/hQwNogCqKSJSul6NyTAzQHhTKDt7IXBrIC0F2EZmLjzYJJRE
QLJEWsocIDKYxLHGk86tDGEOYm/DZ+1MXNn+4jLBX4RBtCT6He1ZKulSBp8URpyR
mY2ZRvKNAxYpDNh4uUcVeYCfEI3PlwEYm59htFgB/NXORcx2Gpiw5Qh4Vxz69sGn
mu8zCwBeINEK7I+DkvJ9DzP4idbcS4onNfi7eFySP/E=
`protect END_PROTECTED
