`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjvZ8I2lDyZdYfHl/KzjAx1oX/qmHnSDfagHUQ5lktxwAYWzRj7xNgMj0aZ+COwc
jnyNTUWPopa6Dn2lqw5Mkc4q8iTNKGFWnUaE+ghOm47wIfnbSkTYtmnz7EU4KGhs
KjmfJKZHQo7E/JaPbOsmeAXuhDawDgQYjlQBNElIGKm5fNeMy0eEyme1l6kbtkOI
sfyK8fwIf0U9hx1v2VoDUpLA+Uvii2Df6mcDlrzs3Qr9OAnmb8PZR/gBwFUVEL7J
Ci+v6N6TFw4jqnGjRgSgEkuVHhECWfUpaGZv4MO0YNxxUuQh2QlqOkjbxwgW+kWw
fY+liNyh1RBGUpRE8OBLYybvYdQ77iOejZd+OdtP16ryvvECGHRzlzBI2CWLnoGM
UFhJED5oR9vWCTPZYJ1K/qbB8OdbBRwrwHirMTuYrwiV9cfoVpxz3DZ9UeN6wtM/
Glf/YA0JKM9kQCqK02v6zxhtuzEjrtMkf21DoFZtUI49RDeWyp2TakZyIOMN+f9P
XRM6OZbfCUfvhiXGG1RLbx3/4z8jbk3QS+gx8tV1sW7+ttIVrkHwBs0DhY4+F1Jr
UM/3hoSFbgtFyik5gsYt8lK/Uv+YWGh/b0B5e00CYG3Cw/Wi5H+E+3qLoc2tJS4R
lueGw8DNBLxXleSQDu6hzTOkMO+mHXB1O8sn3cgX57eMgTs6amIWauptl08Hw60+
PUlLnRmLeDcUkutT9hIgzp5bRXWf/Vdqo3yFi6lRzId8b/rFs/hWEp0Y87GiHX0z
Gz0LyTkB9i16d9fZKGl5o9XpMkVEiKi7f4pZ7YZ6Y4RA4gbdu/JKbTa7ZhT+8U+W
FOsBOxlr2OHUwGe90cMwthPO9dS0oVZhPk2qZ8qJgq+Lzivtb7Qe/hxUrwGGDKJb
gtshSWv7SPP6rxQH0AsUReg3D0pvcS30S1+S5AIxwrMWzE5XqiBYdiKxTK2NRbwR
E1oPLxXpet/mV1DhuLbF9vCVgUEKee7H348207L2GcvKoACTCYWo4LqcA6lHiH4f
7S6zowaLCPvv7tHLclLS8YofAXb+dkNBBPegFpB+CwownCyWtBYJ06oIxttZ6sp+
gG+FhIEkZcnAbtUDvaBq1WMwE2/IBVwIzd5SafUCxT4wu3QD2vzTLyxdSyuIJrnB
A1lOTh89yrRxkEytRaqBHXZyqo2cxYMU9YUQY7A2aKBbt0vBKurrbNPdk08isFC/
VvanL9AkNB0jxi8J+zuX+udU7XSqNgYvIHX7NYjOHRGZZmXrEniOjX+2izn2n9LP
baPDsGuBAT9/KsyejsGpoGRL5muTiZJgrTjXxCxvxsipDJDYubD6g8TjXYkKa6ir
BmnXbIQWvJD059mOubFUaJltM5T3pHcaCuvZb4LJKXpUfh/Mlrd/JaPcZLmuQP+x
2s2BAccn0pj7mYQpnqLertTGTdkiiitBf7BS3WD1WGkILn5Rq3GMSWi+ziVwDkkQ
wpg4VNZpqMdzn9tU89IhVVT39oMMjWpzzpTyOyPNLrbEiTGut5SUKd4vZWOZeg3W
UrkvxCxhjoG8rYIva20d46mj5I65ilIpEcAXX+7ytOoxGh5xyldcBEWByx8TmL7+
mgc40THyrgJYKweCVKhVnjtbFepm97yXfUU9GmUvKbTF8qGfrjhFVZBJB4EBZznj
Oscffg25PgQlxLLvXs0YFyHneGjGtattbA1YYrL7lrHpl/82GGKRXr2z6QhTZ2Gs
y4HAoXmhMdmEhAW0ZPlFoU+DKWSwheUi0H9883pvRZGVxJ+GkqyGWELtuaEKpNDv
CkQxZpYvzassh40IvvIPHAPGET5qxQJ/hoWPEEjEmYrc9N6tiTlnv7uBPSwQz0sx
js/sLper8Zp+FGlQ5jmjlG5g97yDG5cyb4mhdX4x/AkXaliVmF0QUWyJqqezBJhl
LqmgXiHPxh34i45rrlMZS4oR/FF3DFtWzIzmIn7s0EYGTB030RH/WW34iplDvUwB
gO9vgkrqH76pQL8eo03LKzmT8Zr5UACg47i9YroEjaVgnRRK2j4cqScj7lss+7St
3y9UZaMhyHqxHikHre6So8b2Ks/wPTEkiQpLCXiQszaHwoy4CJC/70TwMU/MZSFX
HbEmx0jg3Uga4qFuJLgVdiqR3AeTfUEdu9NwX1AJoNDoeueMaso3d6bIHfi/nzmJ
MjHi13MK7dE40q9bFObPNFgjPFkZfHQFxQCnpRYPdwTf+myMa75eTIOnbsSybJGJ
H0RpOxlk9F8D3AODIcx7/xzpqZSJjYY+ERb0db4M0Oa1NpG6dQEt54E0GDzwMZXg
cpjdvx9BW48gtYFMsavrEXUdznprlvqwBpgDBhCLVQxKeWbng7O414CEjE3TsOyO
stCAqTCAxrMCoz6JQmNLGDv3Te0191xsDQwJ31+bT/+6QWPYta1j+812C9VrGSZx
zUh4pu50NgWPJ4GjnGPbyUwF8FBYPrv7XkCeyZpHKuHf3ldA9mKfMTRhGHLhtivl
vYhSXgy9AVNwR4LeRt7cCV+NrwUHoObML4L5/UxK1mfN4tGO8SzvYRk/RLTa4Aov
WxhCkm921a0XC6Wy8rhGCoAhOEKICgvcEeqXT6m5mEzWjCyVwCstgai54CjBWgFs
KSkEJI9qEOHocDkWVm0BIYnkfeQU7/nOpKOMcPtNuolbTqjd0AZqghQHmV/j09QE
tP5ouZlxrpgjZkz5P4YMXyzN+F+aY7FAC1bYfhoOTNCGcilgr+4Edx20KMfoNQaJ
2GU3jCtR8WsOXnNYKLtMEcOzJbnmvW4oUgpRe3ehElnClFER9r64FhwUBbwAOtOY
gLIY9NfbJkMWM5oE/MTTy+AgTgL49HwZbxmyrp4JPDLyudmxPTVlfRVeY3u+UE1c
TIpIqe2cK+HQz/ikiZtt7pxUffogUwo5LGjrJoX4W8e4z+23k3iduQH3FQ1kP05T
WEL4JKS96NUqps61+8AIkvXmYbQiICyaHOzcXOpCl3o0mB1ZtttF7Gsk0LlMosGU
`protect END_PROTECTED
