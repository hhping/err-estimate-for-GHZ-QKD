`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pB6ELDrxOl+UJxi4x8huThF8OEn6uGlRsV/cEMhJN5FKIbNsaGhXSIZDWkhtZKKp
ojrPXagi5D2nLesJstg4KuPSL9F5w6J9ogsERpQ514JIp+obawG/TGFYev5cRVfH
tHuuqT/2j6BvMWSvvzXH4wWceJI7PBUSf47X3/sPfgGrMhI7ppMPtf7Gx7TgNmtG
mxcFlbLyLew8xLJ1at2Qy81dZhZQjg0BuiadM8flPDxh3JpZD/0KNB6ebUMccuj+
ww2u5ENXptPOwjzsoVlWHIDvpbajTf5NWQc2iGlDdcZaiFeLmEyKvwx3HCM9LdrE
A8b66rtTl2jQT+JLbfUaK4NExMC5Ob3jU16vRJavlZ9IztAWbkbb4SHPKkAU3yoY
DLneFg5AfocX5u69Qd31aZzQ/35C40gzqMKali6orGwj/4+n5yU8dLU4wjtTYqX4
T6s4NYltYMyJfdJfQzSgdKWu2P4Y5SEsZadAnuX+RNIUvr2yXnXT3yZ+ehwHLRWg
A2QRcawip2g0QW7E12Gde3rRYd9uDkMrldhD/nVkDFUdtRzM1Af66Fj8y9e7T/aQ
UIQYbFXiNxG7lgvG+h5f42od3Y8EbrzGTcYLf3d4+8JeX7tciFoGdXb8ADKfR8Pa
ewvp86O3RhzmYs0UWP049tUTuUqETK1sHFu59G+XNUYEOSOkg0T1pBhQEpMOYmLs
XW6UQ2iJYZg86FJKU2AxxGrE6kJbR2sQFsRh5ycQeMRwmV7KtyualgHX/UexWQqm
qpwxR57FHRwwP8YspbTiKztqsyzRS/L02XcofF/LRiJMkWmoKRw+xLwgooOPbYuc
nyD66qvRfnXxXTIbJunqpAs6JvytrYdwKn9D7R9uwSC0wQ4JltU5p1cwbnOvtwRH
Zg5AQI2OQFdZ0YgkGIHb/Kh+i2wduwIx2UdnSCHkyF3Dg/5jit4psbc1YEfOIG3x
XEX8695kGYi9CmRNTf8k4vurNMlR/OdJQxP+qVIBGzd3duZ4Bhg2VlxMJ20TD8l2
r3yL+UPUAdEEDQUtlwgFJX9yI1mbHue30Q8WCNz0kAVxGt9xgVghw6jY4bVfWWnf
s1AsVwaffSgfcct92jROKMbFZnADCcJB9PsUzVAViEfPpp+eKDMib+p0j3UebmpU
ZHhKWekf0TBQDbtAu5Xx7nffFaA6C8u7ZUJqZmd5ke+3iyZ6RNZSEOVxX2fnE6DS
MZbjypc6sjsgqRVYMkW3ji/8X/9FP25RBAA8P8BVThPJ+YQ1//PGPAmM9NLGFR1y
vPjmWWppqxv1wAgbveUh4rtk3T7HtxzoVMZ6znA8t6LtmWiuYTczIXrjT+ra9ZjI
zskmbY/VSoF/zDVrHYFFcxSTfp2DbsXZ4yYewfGBvEu6xfOcl3DBDqVRcn3yV7Sn
FL65FUIZKLjvwGiIPH1LXF/LNZ/V4OiUS7QLL6nPlVWNXZqvkUWsspzGDCZwMMqb
AcdtF1x40VRyrfuLRxdooY414gYXzYsPb1d7PuebQjgbdtaZWQcjDm95yOnbg5oY
al9mxyqI6ors0eB1hdpOCLSX9iiGCZ5MqFruKX1xOVxwRjMazeEhcqpdx9xkErvc
tJ1tlWmcXhUuq1B6Q4FIZPFsgKeD93xa9woDV/QIzCjKdEz2vg892vE2t6DnVUlO
0oqyE8R36k8byui2/axFkJ1wML5vLwulKuZgjb5OaM37nEH9/PrZJYFlUcH6cjpM
2U+nQ4SeyzLldep4CUmNEW//XpCJfiAcq0H4ceHYeJc3/+IBLgCdAg1Udfbfhulj
rEQ0e3e/u3L+u/4bsT1yMurJKHNIXFJuWdkwfgsTKXbBZnBGEL5QQZx+2e6LhRAm
Bmno5l4AYSsi3PqHlWPgoyA4DrX8QqpXHkp2BLblYr5D0IESPWA8vqmWQrkpLDQn
P6HCQZznepk386hPQ2hKib28zttMmM3/9dgytsjMPNVUte+Bg0yAcbZxQTnwAfWy
vYuvUFNQYbbcUAgvXkbiUAXV3dvTbO2ZAZSkeEzrrw9l0A7HZrAmBg1RThMRc4sf
gvCdqbTbqqU6Q/akEEp68QrDpPhnOOCktFIHv2pEuCYFdeU/HU44HW96hgMdkO84
SPTa/HIrI7h20AVEBBfY5qnA5ZE7ZxGkXxsKJutrysvaypbRNL6YLTV3YUe22gZJ
QSRbcnulJIZOTXjogmV5hF5dRy0O1kvjSZ+jm2ZVX4t2g7I6lH9wzQdWb0cuK3vS
R80mBLDowbmcE2q4qVNjn52r2g+KvJb5RzNLNgG8Xq9o0EpuI1UHiYNLDsnT94pV
LFA1Ru1DU+mXGf9hv3aICMoyIvP7FW4H8HuPUtxIn7URximDHvfDmPgYq5YJBcwH
fwQe2Aj00bKU0SDComrFFxyix/2QQ6Obr3ZeBqJLcvHOZclu1ZauLuG4O3Vt/XAk
OM/pcx7otMqAs4zG1kjO7Oh4Xd3lyKhN1jItCTjvSbev8lga7MIyjzEbaJfPBDOR
HQ0EeZIs9Y15iZQ4zmH17WDMmqdGUK2AX4Ii4hu66n39KsGLWrQELSeWH5TT+WbV
lswYgZh+EZmXTw8AdZrzI4cV3a1vbszN/7/zHERblTKv4R93QUNmLUzkd+iV2kfJ
jJCbCCwdyjrdQM6pgtcH/3ZQzOoZ/+f1wHklRsfqIyDO7245JAekUoWkY4hdAz/h
4iblhbI+eFIABiWt0jqIzUFCvmmJCOI2/jyxgFpt6gUBtEYaipoRo//aEfH3HX4K
Mi8cAnaaJhGVXfQMGFvO/ygN5b+OyueWoddYS/IZcJqHpBrYVjtUh/V2oHgJMC1r
v8ttHjiAxVZ2ito8o1/mckOJ1TyTBpbNPsLCv5ELgTmfVoj73oERQD4MtlBr9H1O
hl69Pzax7zDd+5+DPh0HaWtPajjMjjKirsrvcGvQnrImCjsmWxoE9iiqUdKL9iim
0RwwLBTjY9ZmHs1YQEMcyb1dTtKvgYgrX8NcpM0RauzvLn1ejmJuuWrrZqWkAqDS
ywQ/nkfHKTdWDwpgHAE2JWNUxHuN+8LPt00RSaGvjfWziSR4Is2+mhS7i0E46jzP
LXxiSL4BId9LlVdAqLZvoIGVn1jHRqqFZuM01E9vFxSDSXAAz6Mi6gOqHO6gL0iP
BWG7vIE2ZlRX2hxzNXuYyA1Ms0BYRcK6qKzJyoSoTbUSbqF+QwLv+voEViuHZEK0
`protect END_PROTECTED
