`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqTFt/06hNjbhLH2ucR7RosENgHuRRyUPFt+Y+gg7LW8K0/267euiY2BDcI1MzQ/
WHbodmAQ0K6i57uzT/1OnWf5aekfX+dNbIYM/BP7M3w7yeM4R3J4nSmhBPLqvbDD
q/rKBSnKL1i8Mv/blh1tQT2d+5ZQDF/IyFG9bm/7fqesxM/rezhYvv2i+dO/CqFx
UsGC5B77RYgf8kmtjeV4+moXg2rNbJUXRnfPv/58Ek+1w0blli4FptlAoufNTjXg
xr1rdeBzagdm5oGOPnAA56zfXUCeCfGjSE4jufizmOnqVFmSspFR2KVlA0Q3Jb4/
BZuMF4PP2h/gEI+Dc50VAYmgP0n+zRyPGx8Buhjxg7y/zt6aBLSStQbwFH1ab071
WxfX1ns6GUzmln5lbSTFclCxTgYAEak/3Y04qCH7rcMUOoHwEhjAAmMo1KHU2Vb5
qMA3GdFWEzq/qbpDVrrhrnrZCzbbI574LOc2dzjpoI8cR7ZFHXtPsnNblBKBVPPz
bTUds1UKz95C3fFN8QqUg3apy5OModjf9/GLwiQHekMl0CAm7B+MdNr9LZU4wafn
wWfT02JxAdmS5dY3NgskPuEfnqcrAEBDjS5CYDzIIrhq3Whjpq+MFQh5I77sJBc/
PiGbD9Y/jUFJX4CT4LprpaBmA5MQXa2e6oPNn0h47cbripQPZZvWzTy+HF65pEYX
deBdtL4BOzgFevgrbUJeoOdfSwKGHPmVbHLDdeerS/jVppMahqRja9bkkpGVLCMx
9Q0L8DHSNl/VsqrYLqQl+6GdFNaNChrzk+mL9T7YZv9P+vln5BC25Ht/5lxXb3QA
j7VwnNjbmnEw1Ny1ixEPHDA9RnUKeDyODDl64bsoDNn0YqULjF69kn4yZbT/1b3k
JSFjVKS9certmiPUBAMau9xRBceZilfr1YPzwxOYoXJ4niW9ZC+PDtOrypK+avlf
knW6HKZstRKnok426wMxPx3ec7xlTl5M+7RaPszypu/e4KFFMgaNVITFdJXepC1f
r1c18PpmB0nT/QXoULZSzx8TDRUtDYHs8gG8C+F+H7JExTqS+UiN5NVA19Nr6Swk
U4BbsP0vKNkvDuujjI11aaVIZQ8tfx9jzzo30VzOfvbPM887JAB99l5og2HFsSnV
MWt34B/Jdg4Wrrbetw3UXwX5LwwY+8ntyYQMohdwa9eTvKytI7LQ3hyOCmt26d6z
E9c7TDRtFeYssiycjr4IClM8k2oERqxYKuMVL+UQWoVNFpRik8eOFWc+eDZAmGT+
FLCZn31wOETdeleT6z/sMYXlA8/CUlV6NnJEdCYNSCb9eK5DyvQyz1uT9GJJXqp3
3cOEuglUaPcFOUIRTuQeeIwFc4LS3wItym43PNIrEKV3J0K4nzbbbDYRmaT2Rnyf
3eTKX9hh5MzlhPnX/Y7k2L7DB962y/pLSDDEctQgrVdTqgNplkEzWHuk91E7E8zF
EmfcyhXYrotvXflp6CC8EOkZfodGTQHGQJCqjISygZ1goaxqQqtF6DvHQC0y2V9d
59LYrCUwKIj0plEvlXlHt4blwCfKHCaL9fxi9+RDCL8XKwRFmXhm80zfMikwywA9
9gWqq9NWt8TJci53Cli4jn/RcBXdnrWDewmlojC1Oxp0MSUlYMugyfQonqJmVcwD
6rFAQ60E21w+eAp10Hq1W8sh2XsKb467lUPpJchjnwu95nszRzqML4a2zLZcsRL8
rQtJlWnfhjiL4j3EgWbfFTo5YrPt04wk1fCQcRWUPxrviV+1X8epmQCcZP5GxeUv
js3Ab5sGIxdRz88pvZFyTWwfV1zyjBicN8unPm3TX3P64E3vjbXSDDGTaahzzQdV
i5+CfJXOWomTQ5GtamHQv2bQ1nU9Ema0et+a+9VnzknEy0plg5jH5AQ9pIyUL2N4
RVKgob1XIGDkBFENN7k0H4AfLVzm1iTuiAxR6Z/3YttBAEozjejaFOTpBew13Ao2
ywDp0wXuHlbyTvYzS5J+c1o3YYIQ5vyljXjaUmBmgTNigb0vV9oseLK8QSucYe15
4Y1G8D11Ytq/YiH86ppw6+mFCsWGjileBjV98Bv0liLcTA4TdkIoNFczuwRRHj2w
TQsehvEX8nyZw/+21EVvqi4RTWQy3AiMxGBMpS/pAD/RwXUtoHnSEBTQDn9bN4bj
ads3Of/aRIU04pJeOiQVjVTWEgeNLATJYoqwwjTsRmB0InqbqW4XzeO0rCw/MEGt
qNaKS+XIRSMnZ8VRdhdsEbCn2U/hdAFNadY+uqMUCMHUGzspyGPmW5ZuikhIoOzT
qiOQDgmbVb96TfsOMzPeANtAibA+lpkMTK6nIHitMDIgsDhAzkER6XPoFEdaVwl2
Aos8RBR5f5S8jEXbYtZUksdd9PKaZP6dMC2WFMe0qbz0XkYoq1PrbgFdttezJKkb
GItEXlTrzq/2Fgk9J0Iq6dNPtH1IZgr/xLcLgc0Y3tnVyczB41Y0JZSRoNieVy04
ZLD7PapBv0LB1ynT1vO173vKNd6VfJs/sVOCP1tA7yFnSEt+5U+/gRrfH8b9Ks0r
rjDVU4EqAGJOpFnQdPtBup4rrU/EZHncJ5MWSOYgabch22EPKRhbwuW2Y/xvFo3m
IyvCji9Sh2WyD75VogDKyDA647g6yluRADHsxDMRo0muUY3Xbt7JWaMthld/nB3P
XFUIBSmIJDAuf5WXvsGJ/mS1Ycj7Xs25O0J4xcQrincB04T8a0UFUqmaLRHEbCHP
ZIrT3mxmRMXHpMkaa7aenLTLV53OVSqeLCxDB+wXV4YVOXF3eadNnB7tTQjqInBv
WMzXlWq+wxNvhHuk8mLnN929S3iY0lIabZj48o33R8qggxqr0Pd2QlNjXyZnoZz5
L8aX9W/DdlkGiyhhoU60keT+VDTYaTRW+0HQbdBvj+KGy/ZDdxm3lvqxb9ZEAiCy
5GwVFt2KFm6uRQKsTOMOlczYyqL+9x7pa8L1euCf6/HskNyVkbtWKRBZMAnSsonr
FAAqdWxxFPMKDrSrtHzNQIuFonsnSfxVofbpO5vZLT62k8pEZGJKfarFF6WptywP
BjIUGx66Wfycm2a09fAarqKxiMo9wxPwwmRlZKzKpD1UpBmW5Zd3fBiSAE/iXpvO
PX02j1XpGb57RqLkT51ljFgKmRpQRVJryX8z+uMBd31ULHvNoNVvwRWg7htg56/a
/0QpBmnrPkGeULnhMPPXCdzCtX1q2zvWV/9mm8eF38dO/Yde2UtwNikj7Br4VD/q
6cPDr4Blyi3rplgkchTTuv73KCM4bAawTheI4amOQLXwFcO+wNos4px0dfgEiEys
Cjld1ldWVyXRl+k2kPWrG66mVXvf9PjS+RbgL6u2Wg/rohoPA0HKA52V3HdFZDgy
0qUGobrZl2ajWLQ672UPiI/JxuAjwY9Ggb1u+7vc7lLMUBQUHSO8SYiepNKMEQAL
7Cl7m+kFkE7QxZPoi+WpWflVgatmEVZWCwhVshKlcptTZgRbAqvGCeW65FoozoxJ
Ur4gf56d7t4pSDykgZRSItZCLZ7vl+rKp918eoiBnOJ0oJi6M0Pyk07A3dLGHtfF
bvgYTsUS6cDc5V6p4qEoddVdYRtbJuC13T+aQFWKYdJ7JvLOxfm+Y8O0w0ZyTfoq
xwGG9VHCcHkIWqil7mTPPfI0cgX/voeER3X1Fwi8LPPdU3CzGdRYCphnfkJ8RLDX
OI2x/xjXvapp9ysQgs1y46cG5GFXi4YGcSqdVKdD8446aYzvLRSIM1NZI8fyVgxK
isG9obIJSO8cl+PcqAyUBGaMMjYFs7JpacuObH96EK1l9rkOn6kwLzG8y2eijqez
4q2FsUh8FULEFJUJYvsNZfsjcjEu3LwbAI3BkdHJtF9rzoRMimhsHjbfRIar6VDp
sqvA/l5DC2liRVulLEKJzaK46vPoquvukjsipzaVBkKJ0V0RUpjuhoSFzU9wnK56
3rzPj7Ghl+Y5Nc05yz09oRkQ8duY3j/efwjxQJLKi8HvPkjISR50fK3qZuSTpK1A
cNEXXPcFKFL9gUW5DCg7rnuRoy0Y7dOlD/Lcia8sEHPOMVpLkZVrLiwBIF+jQ9qP
SISytVRpNDKYubnOAVzwL8sNRIgxs/uLR7zmICB7eQG2c7JPDfVC3rHRAiccpkN5
xCg1OOV3Tq1eHHJJZ95tpljbHsqhgUs6xRFz4QrTgBbkh1Ta8g7BbSIWUTZBXlw6
0fAarU2MArNPYsidC5Up0f3qDg7Uj16uKo9ZHrhyRgzwkgBSq9n4/qpyPB8Nm1o7
eByYMJ5k8kXfUD0Eia36j5+zHbIofd8SjpO0AnplepUHv59YGUIhhxSOdjasq3J4
+mw8FcQ78X0ThAChWqHVyjwPAN/7xEaIXpwIb7Di36r39G9+UZZ+48sLJpx0PRSx
zrxTPZGdaFuFh0cp1aWwMIpAEyl9xlIOOSJmi/j4ClhrY8Aq8PZCAbklKK7RTNQE
qywGtuVfs2615zVyF8yLC5qN8kbOzpPa1MhzwWW7QwK0liYrw2cwirHY4svW2TV5
hIkeW1ixnSU6D9PjwWCm5VezjXC6OvNMHO5P9ZCsVTotTcoOMCfE/DsMZbNTbNkK
GHz6+T5hwYJRazHKOLCQBvQ5HaK/YRCnkGlNkMy2BQ9auu05knajLAxzvivVAiuH
IhtPXiV6iROaiOp1idh+iX8rhA49kfTNoXcN9G1A+qtqFiO110zjix9FpOnrwOcF
9g2gUCjT/3+fEx0HExrKD8+BLL0zpo0CO4gf/wuCAZiRMvUSqMWJP6xtVbpXk6Kw
QUwhLPnCGiFnpFa3+iAw4nmo1Gf0XYAI6nliDNEW28DBf+sR119H34/jDlygaVFY
nosmu/Kx5vwEHJN60XJDiryzo/uQFXMnT70dJXUxakGo8fMe2gQhWkPu3fb0T7Kd
F8RUBuXGsisJNqcZ/5y9fJu0y+HQB1l7OWYM/0QUPnhx5IabhKqh2khavbgqj5fr
zVn1QSpKPrpZMyXRasyeAb4+3hdNbi/WTTWuTzyKiOlFx07EbXRk/wXRUjIw6Wk4
4UJHG6hlj9dl45ZZJz94Ml3SSHoKopjbdNpfgHrf53O8YL/IkuJYRZRwskfcnx7i
hHqQxxE8JNFTabaGPmLTwDGpCHGgqfvdPHAa0zMrRY/9q/fzYFO8o8AKxqj/rYkB
9Srx4AzWpxAvkxwEuqh8+ORfcmGKX+wGVDC3B1/+JV9UUh9u8hATve82YHdyslsF
C/C29bg3PzM5NTnlrghrhDeMRCrxhu451OZdX0ydV+eB5LmYMTmrmVrODAZIpNbg
thGOtFCuRhNI1+k6r22Dg4FkysY22v5kWCvlVOCIXfvCg2F66HUdeefI9FphhdjJ
M/sbMUg8jtP2AD7VzwvLCflSL7STZbBkXXSJfZKPwF6JMdv2pDEvMRYK4fFwYoIT
G+/Z3WN0Kvuet62bSbnkWKIflnEFpCsDhtg8xdfyubxuPTV2FY9IjKA+JxUeh30R
xWfY7I14rgJhS/iUjmbDA1MTZcs4kXUJI1BF2rJ+qqwXmkZlwxh0KYzhsESZJezP
zchPia2oTcpdhlQZJSRmZ5U4KN8iwQBfwuj1ZbqxvYDUT1f8WT2G38EPt7P0bwVX
igt7pkDLvsVZrCUqdOMeqLKePcFkN48tX6Yv0KzXyyF4MWvTCc5qDRIjxCSExxAl
utCNvA4jmUhcowprmQ43JC3x96tp7YYo6tOk3OmqA5sVKH38BSCjKlWrc1OABi0N
Nac1pDuT6vktnrC3O9peH5UggOancHYKRUgGKIB5am5W+NaLsmI258BP+XXWnVDM
209W3cHrDZYjxQKsGzsC6v58WY2M0biMWEOoK9QPjbVoXEr/WY0Vj2Ntxnof4H14
4nVc8R1gAYfSpJ0oA/d84OJvSloj2vIaiD7UII0uLKRfMDIWNrq4RHEWVJwHYDOI
l++2xEhYaOK9h3L6y+u5sZJfQHX5q1iqoQTafeGS+etx8cUMweSt9engkU/372rJ
VBWQLCG9ngLnIWwvw18KErlc6p8uH/7PJsu1i3rRrKF3P0fikVZZo/Ad2Dl+Q/63
U5iuac7GDezWDWfLfZ6fjH51YAPu58BsmSJnq5J6ya1Ak7w3K1/ywc9C7GrnyisX
ldaipt6eUj78H+9+Hw+B3vbWQ3TE+1mTfMfw4nEp/0xl4I+np21e+SX48nWmAsf8
PglA52mDtw8FP5i/PJZimVX8eP5o4Rc4lNcAfUrFxaabl/nBe7PVH1CaF5iHSJuW
zNW4j1adCsG3YWkHnSj4old/O4pKYNUWJEK5gdutQr+Lw/zlvT1Hd7iI+96zuddn
9HuSEpksVrZzdKaEYCwscRNIvOQwFs4bIKag2fndNZELlt1sMlAqinPW5lTlOCBr
8lrUf0FU7xhwXJzeMTCGQw27CdpJTj06uNbDtsGdODRAZddjN5FecdbgHGmQN/EL
zVzCaSxbHIJxPGBk8LPD3IQg/k8qKNoJ1QekWsC7a3iqtNjz7RvyhMtJMmi7QPwh
l2xLG+22HvKqed4gD0DOGh7kuQ9qq3faf0TD6wuLlX0RoRN0B5MUpP6anlgXQ2v9
avNrfPgJWNZcfQ+qc8V+xeTmgEsjPNHwM59+yqISGHD5TloRNJR7+LPe8YhP5Y1f
oCNQUzZaIt5yc8kaDreOO5l464t15uZ9HeN2lMVFECBO8bS7N/shQ3jKsg9kStkP
bpUK5oqyh0H/+hcxIBWlP9LtDkWhtDlICPvwtVdv3miSs7PoobVkPcNEdpQjU+8H
HoIFnKeOpzKiV61qEqJnOrE9ZPGFdF1pTQ8cqIxdB3QUjfpc3AqtrUmlY8QBp8sp
x/Fip4d4lvXSFkYfdchNyWZp8B37qmUrT5fIzdxdMs/SKdHElaK7U2DP5OrObQ9t
80TnZ/1fYSZTEhwMteBtR5qRFdhnSpNG0uxHeoH77lu0yp3tcNtlewCKhPNq+BkK
GzzE0gdsaZDDa7xnhiMB5B9sQei8uEyLxKO0WlHG1I+v1JM3CiF0SmJ5CAKzV84w
WUb5XwScifR+o0Kdq7M+Nig9cZw8L/ir9AUvOGCbv4HBSvoBINrR0R1gTtYkyuFy
IBBGN8Tx5B6XRUZg9s2jsRYE9KyKCJh8nOrXSxQPIpeAHqM9u+/ppUKIqXQsC++Y
2Ah+T6Jy9QbH2hGRD2MgT23wofltxu4Bb3wbqbhsnAUvimPQfI3aHQO8yxKkH+om
kVql3gRcjrsHrpJwa9KwPg==
`protect END_PROTECTED
