`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WOek5ubs4sDfCN0tmb7FG68whHE2uD8HXUXxw61/0PVSjkP0InLETo5hbd4gss47
DGi3N/SudfDVCddWvlaX/mulimyqPbcN4ioi25U97uTDWsNLC2/L6GDwEISw5bIR
fznwe8u86Tfd6Npclu18MNUfbSoekfrIXxuPX7XcyecpSXciGfrKfI141KYgZOX8
a1EOC2t4l3A9ULk7UY+k+R7cWB0GzgkwmHDQfWsh9mPUwg4KSih2kYwCcTK3PA5W
wOhBreJBZEaDXD+yb0uGTzf5eWLNmw9IxmEuBIZ1SCc8+DfRuuZpFpB+oX3FGT/4
p5yj3Cme5GhOy1ooXlHc+Hz8sQePAcO4wxuCZ0oP5Xk=
`protect END_PROTECTED
