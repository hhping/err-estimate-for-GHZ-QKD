`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2aJWFom1EvD6sVRNYCCNr6XkMeKcOd/iTtBTqZRtIl4eLM4MfhG5ffibN0qcrbc
CHTR7+5XBHajhH37oBxOxd9A/1kGryHSI4jmttXX6FIbqkfGU9XnMJKRwYdmlhxX
rCLM2QR//8LFEf4iXVCi/JU5VYavpullMIoEyeqdNTpPBHVfyzqy+9k0wDM8ekWb
WWINaQnjlmkacazBGKEmZp59R7fY96gbNrDf+y6JL7Dg/7xsnTrIVirj1wU8qlCg
CwLxEnxqLJIvgjPCZexB12zepYJJLMJiU1fVtwvSmHK6eHtT3IpUbfRh1UrE4BkE
o7yBHsyz7/yvCAHmy31ovV2RFznDeQQPcsx8MrY3m/ISrq/ko/mEkFEHLF3E1Xbz
T3Fo5iuPthefafFwS1wEnq2pPRioW2aJNs3Gwhra/CvWKklXrWNyA1cEPw/JNeZP
fuGRR3HKRgENl41rc2p98Al1CfMMcmaj0Y5q/dAzO4lAWpPOFwNYq6rpWq8pOlZr
63B7+tFPDt12sMu12eA8gvcArT+R9nIl7Gcj+QOIWf2nL5D9KEPiujYWOIHHZoEU
xX1W04nUhMi1i7PatP30LOYU2SOvr9iU7bWTGMHy6Gw2oDk6VrHvx5+/FP8WURk7
XyV3fGfp2AdwOa8y5JZ7sapZaMwv51f3WonN9eVkRL2z41vtQZC3la4jyPh0tej6
1YSWv4Ne7/1yUh+8DPrWn7x3Uddf0ujnhk+9m4UDdznZJ2UNz7LIUJxF/cjZzYNa
SyRiK03PK0cH1CDjNJz3BGH8hf9bgeQFWRmYV0aScIFzHn/NwxF/zjwWb0gVFMnf
/fcSGED3vQeTzONxy39K/13NOn6FHGvj+7B4QTjcdwXyRdgUpk9mzeeraBEuq+4M
5ZB/yzOb4D3KkL0+1Em48Iw4QjON6h8eiYoCDPbW9I/1aZPI9CiLZenCybbzKmER
SlPkwn12kxl9gfFKzlV5bDxpPI1yxo6ZGXCzb45Qwuva+RXFfTjrwL1s1kilpoj3
E0GwfxFKPMWzm8H64Sb2BrAmvhcEcmGVc7gcJAyyKEYch+cCEG+Uz+JO8TOvXYAo
hm31sslhbnpPManH3KjtIyCvJr4PkJy1DtcgQ9R3pGYFzqvBfU1+nFzABsL0pre+
/MlzYOJu8YvyqySnBKsdcOSf+myrBYg1TR6qrzllb2dSxON2IDeQhkhFRPI+TQUN
XylJqEynhwmyD7/ksdOV+5jtFkJr4XyzEZBDFDgz489JNfPUDNciETExKcqqAi+d
xYqKQNkfrspPw6V/ehwb6GeTMdf7jkMgwJMYDMweMuYhVjgjxJmsa2sdLwOCFRFA
/YkqOzDg0j0O4majazU6F2zOQjhPkbSdQ+fuQg3LOY582Sb8DnkcIXyscokZmnkL
WOUjAjZW81ZxaRaLgxmQQyYtlUlAuUXwM47bLOnHX7+lvfpf5iW9h11HYf3h/FoG
+l9xMWs9QgNJ2heZ/FIvuWj1ecZkWRe19VtqRNEK7/28zI9d1ct8kSsnylK2JimN
5r2Bj+rxfiNnSN64lEDfYvuvanWBL13/XTll2gge5b3eMhDM8DucDBw93jFxsI2e
55dCL3h4AJCy09TnzhbMnni5g/dBamgO4fxIrhxESYEEHRnmTRQ/Jt+JA67XQ1QO
vPjzYO3WHYNAMDjqhHC+Utjzu0Ef5KRorNXrGbTVvQa048EgYgqg5tjfOsRuro1H
bEJN0v0IECHoxKwfsie9K9FpuS1F4epe1LNaG6tkFl5vgcm/6HTxb0vj34XYxUE5
REKlB/FqbpCGBexTF0OrbYfvxo+HE04RcVGDaSGpP3flROMHRBk3Fw9740uutpDZ
V3bcws4hecczwB2P8VAYG4JTGczJ7kEaaMJeA7m3R5QS3zlY0qEQobkcBPCuHBKJ
kmSxgh45Yn6oFX3oZ4vbtzs3lTky9FSbM+OmFdUo79UE+az018zskKkqOgrPkdPZ
9lT/8p8Js59cW7htICyRKIAfvtlVQ8XZD1dZM+uUfCPVRB3yp9NX57KmEspbzk/S
m9qEg/3rwLKSU37TAUUPRJPNmZ9zzs/ysssjdjYtawhXWpo7AC7NJGVgKLPoIQdM
YP15rV25MHz3feVwrSzP4xFpP3u1p1Gdu3FSqj0OXJhK7BPekwjGNSNjWxul2E01
+tgHcl5Jf2suAz87i66La0QkWVDpzsEDm1+cwxfy/fAkpu2UYOfekoY2h87NLizv
46eo257SMD6F7PyFDhQWK75BR1/qWP2zFl3JTYod2xy4mh7oUqMY0avdQ6KmmPkS
W5K685J8nwrtDkJnzziNZQlL3m7KY2HyNYWY/HTB6hOY9zHR0tM5ynwcuwDvswmq
LoQjCOxBQqPnHfnOD8vxeeNDNZmI8yYAd1a3COW/3gWoHp9Zfp5tdyozE4I2pcEp
nireztQm2abOEDqkrQIBjNoFYmUBfyOQhXsoPa0eTH/WHuo04vCLQs037eMMuLHZ
g6e5+pJViNJZfQ9xQAyN8aWsKJCbPS8bNCQ5vSmKsk8kLOgHtALhiRlRo9Y/SIUa
Ani+o4UAlt+5UjVW08yVzfyuHRY1Vu9OemHW+tUFAjKRcPnzy1R7QB6D5EY9V4ts
RF0XyGs3W3FQOSTJPNKvOoDbFX1jLypd8iLidu4WrJGZ5Of3Gk/Vp4YBRnED7S5b
1RHNBr3xSmFpwThbB6UNY8/2RzT2lRly+547BiVpnMLL0+f476dGW1CW93H9WkeX
BsJTeG7RC/EPCKz6GBbF2GovzoAwCkpAbaJtoqsx8NpUd2ZHSreJeHybnEE5jfuU
3CMM46zGEJrSYFgoAqYVv0qWuWwFF5/MNDV2KXR/NGAnW+bMYMI0xD2osHGLSv+V
h90DIozojD9qmVaWO4MSFNvQV5YIm2yHMTQDPAAIsW6dlqqR2BqqrvNV/+F9Zhtm
xsC7SzlwWW5kCqMPJ48lUubPz+sO+gLmiRuHzbczPs51v9UuwIRQla9YB80tJU9q
a8UhfWYpi1Ze5LEViY29dIk/u6owYgDdV66e/owIQJIvLDDlqaxaYbYhQQxIt8i2
9MEI9s5++BefKU3VK3us+fH9xQeKM6RJeAf0W5sXR8LjNh37YciqNuEI9cja3FQe
YCA8rvWcgZ4zOZkYljE8F5uLE6q4DVoIDD1kJFSzfeuIQyIBpZT8/TPD02G6/T84
kaupaxf+ljETztpktmY5WUArIfettiJDQeAcYDtO67wpxzod+4Dr4/lQfvtsDtPF
ifcYBQvpuM/5R/xsBJBVKUn5EUKPKZR5yR/zz5rj2+zNpK3uTNyumWVGM/DPRz80
hEvr6dQX9Ksea9+iVbNTtNxBAIIvXOnqEs4vYaPxB94CRPo6lTZbu114MAmUPRiP
A5TIOMxn4Q5u8ViOSmdizp8FZgKuJWnxJiarur8RNedmBLJSBqHz8lVNeFnOwe03
tNpObP3fnntzDip9waRhVApoW1jPi6KXoe6BH1mOt7ORUJhrzPm54E7hme1Y4TM/
4biVvXG43/JeLaQyAT0Sut57mUSicElMyW2sSuGow/BAVzBj2MHcxHSl2hEsEkXo
tRngADUUSemwUJ57jTq8hGbw7KmfyEk0for3slqx4vUKXYIAFQKeBrn1+aeKBHmg
wtXPEx0UA6vI4h6aznE3raiQVbyukKzJ/K6FRNGrRih7sDQC4XQdSXQjbPyiEvE2
mQ1XKjXTm+qUMnz6w0/ZygvGy0JBJ1QCdUmMtJ0CSzueNz55WC8A3pjve/XJkdjJ
/4ilHDPxMNds9FdKaL26Fpz1hbYEacd+8Q3Cote8xq9gkGq9A2YDILIfnPUlRXds
ng2P3HYCiBVC0Tprg1G1so9bHo2d+L8p8d/n3EJxkePFShrqcdmnJIe+5s1ngH9o
wzemGKa2BBhGrVyaNWchht8yxUvyk1nQdfhD1/UeP3qds4WP1YKaVfClyib7Cd7f
n+sW2kkJpcSRPXMS1eLLGcHyQB08dAutA2wnFE/jZxAqQM7RYh/TfguFZqS6lzsN
jYkla52t/oQuK5YdNBy7PIF1Qp+/bqeISIb0WM66oLxMYOXI+W32a8LUptcfZL25
z7UXP6Jju6jGi5YZLz/Z6zZVfv71ZIwYB6PQrPwWRiPdrzf9zwLdIc9pSrHzl7ta
5H0YetBTMhQP29MIurzhDsz8kbHbRYA+HgNICpCvTqWWWo+dzjVi9C0AZwPeGt4p
ZUqdTLOh5Vhatr6oPdTBp+f7L3bRjYPMmbfG39gWIUSPkYBBS/PApB+Wg242WSoX
sQDBKgyE42sfxqiN0MpEkGG33oAADM8aUvuYo/E7Nt14Tf1ACGwH36g9y4GID7vI
pvBQh3TI/68cWin8jyKcpF8qvJDoO475zSDgfEViGInQBPSWSThr3KcY/01vutu4
CRkjMBIIMW3+AE8em3xqeC7NzBGFCZYXKXnocZxi2AxC8uqNQp5YKm6wNm7UdsU3
F0YQ4+xCyav4texfRADLwGL0iIb2RwKxx8ZaSpPvxdYgqx8hLP3jfbNWH2xDs8yb
lzJlfiy5riKSKaKOV1N7NIFAxQpPBA/qDaK8DsxNRIiPrAdtxPoWQVdhgc3Azolm
FhRvJr5Vc9ZLecqm7kSvy82amlMAVTnggYT0Rekpw1rp+Ef6xMRMPt4l1pRkLiXO
88s0HjKC0zBZnRRDCIr8Y9J9WB+FJ5CmpK6VEKuUwfB8dZNWY8rqcZav0u1gK0hK
RUH1UWoink9vkX71MRbqJVciMpnsbyjGBAz78AmZitDrT154rOoXCVtngBUhfvvJ
gfoc79bov8o2VpqR3gEg2SxDGmNyW9IMTKGPOdBt0+mJ9f8MsX8HdlobtEARqPmI
hd1meBZz+/DHb4d3+BL4YvBYo/Ky/8DbnNW5YuoBDD+3X2+khfOBzDAvXDjtHZXW
dYa9GbuIHC5KBsuD85u3EjhOMtsCo8KSJzsgQ66C4l8syVjCsxfZd7vcW+8mo+pT
AxJHb3ly7sXmd5AYNgo+TaSMlY3Ce8VbkwdhaqlBOFJdZVcYrR9X4j/KFZRgoEAY
+vs6qCqmLtAX8QQWsTkx74ODQHdumTxhF9MHjoniWXhDLhCpGrp/C/ZOWzcFBmzr
DrfM+Z0HHwoLM4MAkKCVsWm9Jo8HyRUwjwba61Si7JKCCWdSqAwisy98dYHtJUsS
6mL7He1SEKckWGvSEDxnuvwvu62/R6WncU/3fzR3lvGmFpLuKjlHAaLK4FewBD9r
SPiBPLJzNIbx2uunJfTPdGGGs1CcOn3/IjiNtcMTjyQADgMI60CERBJsnpUCuExa
GMJSfYi0lpaYRf3kB+yVYTNye7zXKhLFyu2gPATBiOcbv9L/16DvKI3rUDR3cdKY
s2pOsQ2jM/z7e4aJflqK06Z9ugswjytPpq4Xw99C8UCtlhOHKQcmAGdC7hEn8uw4
F0T8m0xu3ihx33YWWAy9Ga86g7RJIiR91Lg7vQY9bkRRrIx4zXpcYD5CoyPXm0R7
DvMPNPlbbym7j24zOkmRx8JKISGbCLgjp42kY0pk+c6rPHp6emxVX2sWFA43+FUx
9YR1RMB7Seo2DI/T54bQ2EhRcerrW09DYgj28ihDI8Whi+fe8p+mO9AYpsMIZ2nn
p0z/JA1/LC6f2p3ZjB8VCvmlKxOUutnCDAs3KOJfHqHhjMf4c/KhvLbxydLGp63o
bhfP+eZslncf2aldo4iBx9ortqdBAuXWEMC0+75sB4d32Gn7p99Lk0tb3oIGN1Zt
0yrlIGOCJb5WpiID4QqqEUKHK/RQTJg72udeDTD45fbodK9p9a/LXe9gtVxqetfA
sYaX4rYnYIwspDz9/NlgeLnOYy55rcR1zWnKdhhF5KTmXh4SPxgWPTDxlgDptb/s
YI1+/dMsoXUTxTqgQAshzhmCw4JHIgNzGZv200aRZeJpKCAUjgYllVhrk/Mq7xir
SNGNmQkG9+yxCLgzYBsUpGhkg32KSSNEkHzTyqlpYzjw+izZceWyQuMZOjVwTX4+
HOo5qvtdx2Uv2LymxmD+5iwe5VETQLo9kNeglKjTE0GRiEm5+lgTsXcTtIZmFQ/z
bI8+t+gGzQqBZ0rPF9CFNrCjI+BBxpJ2qMLYqAe5FUX5oxxLFLTnhTRfi84HDp6l
Owl2SIwoJ3GKYZ6a6xpn1zSBpWUNZblBw5DZ+yZnKOD5oTf6T1KkTRMoq3MGb65u
O93TJJGOV7nascKpF7yGTEsKK/cHBW9/RnW/YDQwF2l7fQbsf36v7fBadjvQhgiN
6cF66VR2xvamO7a3ic28baV0f2e8Gs31NjXdwDdY1oqV0Tm3p3EDv7JC3OrjU4Zi
U7uSdLOJGYNne6w+yIsWLtL5vmQFOzLrGZzTmXvVFD8OcSQxVJNj0hoL2xlKAo6O
da26fB0mLmF22MglXtYRKvEE3M/cv1FBQaI7Bsabroe8MaeKPk08FyEeLVYIeSiv
GNazMCXs+hGd8/RIvBNHFr1bCXnGpErr8RuwIgWvHxu9ZJHjbehhd3VUaH+bT3fi
f5TvF8AaEAYnplImRTEpNeR3ImffiftRTJ4xxjzLetRtZvbEteDeqAxK49ihTrxv
CxQoW+3W1xkRxoQXpRnJj41oZ5kDrxG40XZD1cOME+yt0cS4MLNIFzpRfX8xU2YG
rpjEAwmv40uyNUEkifQxNA+kA0W1cpODdbRhvOe2iB+awlxx/HbBnHOdyH3lj4Bi
bljFE7LUr6gU661Qt4zoSzbY2cuCtIFkX+ucLu9Wuu2jo9gtrhEeWLEroDwkSq49
o8j1yGxi2/YPOOr46yIdBWI3/YfzqTzNhxwnU/VTb+fFSlfNIP4W4g+akiGEYxDq
6pLrDKD98kmFJIG66ahV+1naG5vVDeNBcWRMzVD7BYgI3GgqG1GGIriLpPxcWoBT
GA5UOoDcTLmOz33doln/facairWoSnL5JxMC1PtI5Yw0w12IGccbKmHoTAWdtGVR
vbD9MdwobTnJ0l5tNJcfkb3FJu8N3t5Zg6/22kiGV4rU+BlUQ6h9e9QRO+gEGFT2
l9GgtLRVlBBDXi4yA9JdQ8CFZC9y2Uqz+rRHpIpH8bZgXAoDd7nVzZd1f4ygo2Nh
g6eTowKbQylmLPFM2bykwd6U6RGgB3j+16F9D2+RAgqEotg0EqQn8K2c5eqySfFZ
PvG0uVWPoFzqh/3qkyxiYPSlAmdkI4puj7plCuNXprfrpTejwRwjbpgAE0Q81h+0
/u45VRoNoCHYGbDcgBg7fbWXQw1q/kEsekC1+tcTTovsynyP4MQDoP+XUyvN0xhj
KlffVy8plxPCvNSuGkLOL72lbdUQXQKjc+Tl/3pmmC2K+WNaXBwfbr6TQGDzKAkc
kbdvoKHOXYC8FsR7hjK8dtMcm2i/L1+ucL301iQCkUzQYS90J8+Y5lqmZfkccAPF
iV5x6BY9ZkST982PoPEpsnHFh+rcZHTP/b5woMDxFyrb59sU5UXXDbj42git/hJi
CJEH75WpsjuE8Bgg1cEeGYV6YnXuS9ehvnDt7tETbKE/xt5jb26r/tDewmufmHfR
xDIMVgIvKdvq8e7p6MNMMKAwlX2Q7B8z5iBR1/6HnkSVsj6IAarcGAdyJSIvaa2S
UL7CkLVGT57rpiEcsdInFDgDpRIfSK7A8rWmf24ozi6yN4Xhb3tDXqHO3g6EKwC3
YavkgSK80KG205TQxDLM070ZLCeNyrWuPBwu0as3iFqowx+AxNod/Y3BKv0UDyWR
PmVsX4RiYWRolqo0U9Gu4uU9ASFe/kocdoqMZAT/o2VlK5ZdPCP7ghRwpMvWpTR/
VZ18M8pXvmQN7JyficzD0By/lRHyE1HsD+z1lz0SwTY/EIsUeFK3gF5FsELipN18
jXV01SGV5CZUaLZGQl5lGkEUl0DWPbbJqe//5IE5cV5oyLRjeSljPrUwBOKaqKE5
HjJwhF0GljiMBP3qyiXlG4cA/nBK0Fj78BNvOmvTOUoP96aH4UjUWM1CRSPTlLL0
Vwf+uZx79m1kmtaJDxBOGggji9FoUdDuOKHQVuM+rC/mZktTESd+D/tuMZTipdI7
sCvmfU3ITNe8SX8QkQeBcZtbNhemkEq3ii72Q6v7+Q2eDeJnL1DxjFpKNREA1u7A
SBA7+OX/bqEUMFvi07j69ElzAzykEZAntvp66JTNw9cwNwT3zLJ5raOqrBI1T7Xl
oqBVEGu/e8lLXeAXxb7N8HI8PUWCJwxttKHFNiX1jqN4KLEjpLS3RgDe8JuTJ7r5
FsDn/lJTcHFt19PqruA3+mO4UX7L1tSF4WaYUP42mR/quyZDBJBg+IxCo0Xs03dt
By0QCjMNDUEQme3k5FJSoLZbRwOV95Oxye/9x2AMjj/TOCcmFPBqL2hZE0Wo8now
2SuIUl5R25U+TWsR475VYSfiLAeaDpTTqUiIIin0oIjo042HNriYdxdvyxpN+VUS
r+JVL7mwWZlVSnSl2BMnvksTW1XDjzjFov0LIFL+jpxyPbMQqD+To0xoR9l+9r8u
r3NO8/08rTjUfOUJBgIBUOIZp6xTcT23nX/2WkBW3X+uqe61WzFbN+1EQuEvu1H5
yp4YaQI42Zod4zoLxc+LB2i11FkN3nK7/aNVCUu+TY7YIxWkSPB3Nwj97fLL1/vD
Stqi1Ym7kwvMCbrGAadKTvSJu4mYGhrqiv7215uLI7GC2q2xgWGUnjsu2Y2QgzDH
UMxtJLUCp1bzuBrlo+SuUkn7cLURX+ksNnzYK0uC7hzHY+lknZGK7G9QecD5n8D1
lCVtO3BTCgnLPl1jW3ESEEKV0K6rTrwGBpfJvW1DIu6adWW1acbFG7YGkSxCHTgz
ZpjUukUzS4/nEpEqFRPvHP+MLqjIZRqtz0J4erbEkrzmvkd1CG5W1KbgqtDu/Clf
gpzLRv72uV24GO5IIdJTEodQLDkwz3JG6HSUw3ajIXy2YmTTVn0eWpiKWnGAYal2
+zaWhsptRt0JVJZt51Aw8SR7Wd8nlAQGlFmooOdZ1g5tHIJ/ZlfyNExYIxKdLdCC
N27L7KqFQNy1HVOldko1Ww==
`protect END_PROTECTED
