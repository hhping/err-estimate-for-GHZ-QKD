`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGvDdNNZSWfFzeS/v4Zi/81LY/Xqnc/Vxmndp7Tk5F4R5IRJHZ48jAsH5oT2NJzR
77GaOlMFLNM+zICmd27PT2R6xgt31H38rAenmZhk54fltkxaqL652bwme8Dtd8WI
KfoCtK8bsbvVXMmt9BtwACrXZ/lGB3OiAAurAuAmr974+y8LAADtBWaDLdLz4JYM
RLvByS/JaOQZmlOvBaXHfc8vQQVobuthXbYHse+chW87oXJTGFbP16B9KOB1tThN
64EIRDyTro1UpaBbfI+pOBbGM7LOpovT56D7/qM98bszhLIrwfi1JKTBtUYfCXJf
fF7DI4AZ4aLCX2fmeIoD6/BTiD9X6bNdD/Z8X/PS4q4r1g47l4EwJvxOBB4nmADG
4khf4/45jXXJp1v1Q59s6ieSd4BbVr9Ne5wfWPn5PuetAdyiWIzVfEwmL76cDPYd
ZQCiD1TFPajUsmUq5l4ctDnzD29TTSEEpWuQ9Q3wkpoBMxMI9gAUxW1nyWZC/fUr
yZ0Q9yRn3YJfToW9/pz72e0MykymHlCY/X6DU89t2hNNt+CX/wczTZ6u+QISXaV5
SAMBjd+ynIzsNpHz9nBDPMi50IfiTRtbpOhFe+lTflXMo7SMYmV6GK3yXrxFStQN
o1+q5W+QPMfK9dck7es+z0xT83ifbw2aPPMlLzPw3AciSN0Zdo42hcIT/ycKfKix
+hxiA5ttsFzpJ1XxaGcD8XDey9Kq20hQ7GnSINQgwoIxh58BrrpZtSTGc/FiCf8h
C8k/GhzB72UP4SQX5TDO6QvlofaSwQHi6S95KpNxvL76PQBoUEMZZqNL35PkEAyt
FfOKq56AbAGXiMHieqLKVejUhktNKMlobRT6/AdnX+UvTnh3BfY2kx5zlXkRghM3
Cs74L+gAAKGUBjhrbZ8KDL/fwfsW9huL0UZ9GGWqTkd1X5Qv5rYT8Y34lU9w5l8l
GMmh5hFI2y1P9iWjSR2MJOqm6RUtKzpJtYBwXDiBM8uU/9MaGk5E3JuD+HrK5yZY
2UJKGWF+Euz7U2wqC88wEwZa7rItSa2n+t8du/goyAU=
`protect END_PROTECTED
