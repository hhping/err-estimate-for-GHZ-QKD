`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4HZDNGDnrRWRKUPrBw1YLUbqIK0QTGO5kZDJgyOfw14OnBjJdoy0UtzsIFi/Nos
edn4Yy1FKnkRXKkLt3NR7PsuSASXvJd9FJT3uhK3IPNK8gQhqlNps4cBltWZLgNN
tITOR29fltqMbOsokOyeOB8Aon5bg85jOo/gjXTeJm3wmAb0dINxMAkl4nhDNUys
BBfHXQwA8jtjSCQkq1SqfePIMLSNhe1fC+PUb2RhP+nAux68L4CbtMxCVB0uGsLU
TgqloeVYxigce3aysTcbQ1eIlsSW9IShv1rZAXimiBnP8avT8dT9HsjcNKkSW2Pj
AAFihvIJ0pEDMJu640xxIIhRnAg9QiixOnSGH2xCdploVArPOphlKO3Ql59LLnqi
q6wwKMQuoVf90wYS0BxRBUdBaQJzRfXjnmMJesH3XjbMvG2BUZQkFgA26jajHM16
RI7uOMupA8oDVouwZdh8aZSQlQG3kjcrt6kX6oBB6JwT92MWDyRY07B59wWHDm77
2hP+3MuYutPCyuT+IAbTnkwEeuXIZ0gJCzd+R6xmri5ga6tHTqoh66oz/hNPkf+Z
+ZYDV1SEWTNnLKkx0IaJ1MqpicAoTEnmKac7qeYVxULQIaPDt3k+P+ggZSEaUQPU
cuMST7n240J41+gZYEkTJ6hESne6sWBo8IYhEBS2MGxcl7mGdoInoaHN2TAn/5r8
NE9s4N0lxx48e69NB9A6LnnBKErurE2fc3lEc97221g=
`protect END_PROTECTED
