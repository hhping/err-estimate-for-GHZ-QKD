`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JtlreFuDZhRihdXPqHW4VsH0e7Okp8RrJjBFjGCrx2iPN8K6SMeIUHtTV4JhCSZI
Cvd8lIJ3YQD97dKhoVomoEHR1Pp7+e/FyngI/NJRzcfJLR1vd/ix+cPtxwll0PAY
AYBjEmdSYr/scbTXn7aaYIft3F9Az9lsH3dci1k4Rgy648kQMRonzYAmaOqEn+CQ
Lq1JvHya4X1YI8fnLDJw/MDgmfT0kVgvmlw7d0vp2BDGUSdIVOMO+nfpk6t+oRmc
Z692RCuagjYCl6gpeulMZ3U6ccHRf04GeqRmELAc2+5JcfeK2/0t9+KkLj4fP6Jr
1fBzXhoFZORhzDaNIv5zrYBtNOjqkDP9IMFkdFEWM//XY4AhchTGirPlEw2Kmctv
I36bnWS9LVQvQqzVkhGE8ejOF/HdLQq+B1GQxLj1l1TSnIYltMLamlQy7FiVcHkP
42VCI4qcFM2+0Os7jtx0GQ6Hr+v9klIcJRWNpATTqZJfa7cSjKyfbL/dsTrLwtRD
Yvmo5ONDufDSNfhLmdW8p/Cn7wwMJaWkHw6uT1ULZuLgyqsJmqQGOoEjYR+VExDF
hHRTn3xHRjF8LuxBsPiho+XAlsnIJkpSAWjifqKxDi/8u7xPh5x9yPRAeCem36Ym
NUXXv23DmAjE8dgMnGT4y6IK/oQFFOos7yzxxG7Ku5VMsacSXc6/nlkz7/jIGpsr
qqNoX5SSsc3c6VdahTE50zMDSyGJ+uzF4j08UalL6jNEqeLrxGxe3OYXOT0VsHMP
lSunddiMIi5Sfg2g0M0sCUcWCi+WZRZgjuXpcqvWQ5dfysBetn/G0M3cS74ZsWIr
EMbkik/oNkna7mgguEOYk1B5i/nc5E4nWiy6D6dxVjuPw4fkl1N+rkalltTaRd2M
X4gnNmy3Sf3fbpF+JFyD7L0LZAndeG1iPSuOa+avLxWUweXDkJWCWsIcdLLL6XCp
Ep/Flf7l7P4ubwRpP5CgP3SdXcSwiru10RTNGtAa6LsLVhecdZaP0Q1Rz/kJL17E
aRs50pCwM7k0d9mkVrxJcctwPagyaXlsyAoOGey+n2pkoY65FwGlFTsa7cOVbrUR
M/ak1ZSERWHCxy8VeHprfnrEL+s3BRGJ9ULq6pQFhqMB/5Y3uhnfdvMLRvozFsBe
pvbCbkoCaPXJnBaXPhAiqbxjl1kyRGY1B6X4D9hWWrszKSwEDWtiaDNWoh8Htqjh
IF3nX5hVCHvDWDIzEntdB9p51hYEKzaUBPckEsG4657FfRH8uzH77mfW8Iymuo5H
AV8W7RmgP02uPx0qQzgoL0G9p2EazzUtO5639ormfbbkirzLR4kTgt5vdGUu7Vpk
HNAqrCY/Z3CXCp85fqELsQ0motjw/QMT8GkHs3iPEgE88kgRiKvyU4l/VgajSTeX
gZMsZEQM5xn7kJIYz6ab9lmt9N5vZa3KcjYCRf9OOb+Yj9MAoS9a/ItjrIGG7fRB
KXTyThknHxixx2yozpn9awG3HKBOhsDoONWaWULMSuju6EYIHCFwQltJ+S7ZfNp5
m7kN4clZlt0HU4OR5G0731vfHGQ2unODsD0BBNtfJqo/FmWdaBiv2XREMGEP4cuq
m6LyW7fVQBNftDgLxBdYDNy5ij0ZoYThgPhsH4UYkR8sx0Y16JntBwVJqoZVy/4o
5VC4/DO2X32RdCpisfw77GIAII6aQ2b5j/cPBW8Wf2dCIFw+Z1qWiilRo7Hq+XJC
Os9rG2yXlVAKG+xB0rRqJMVLVA911Gbek+SJDZJ1990DPz91CuZWslFEjk2CLOjZ
8UCg+fqtXIlNckX2VCOg9sAqZjH7FkZ8g/KfJ3S03qD3KnL04XijkovBps0J9RQa
+MSQl5gnrmwakIOAba0kTQ/7UMH7nAnEPxvEfKQprs6FlONhqTJr8GhuqIX73CvW
oDDT3Fz6nyYDvrAqaAVeXN/aCUzsn3AmqCZU3ZnAyD/LExDxPxtEJbSERC+b6Jye
6b+BoFs2iUVt10s4SFQcukoEA5sMBm99NbuBPQdGvJmryHW3yqBDeXwuXX/qig27
/TR9tT7PisGKF9Q7xH+dsfJ5IRlFdJNDxQFaMZ8qJG5NgJPKTAy3euZXxer93DFX
i7PguglFsZh2jz5sp8Sr10o6C9U4Ry7IjmE2TfqsUwfFtLiesS68VrmWVWdJh58u
UeQoA6fJ8RfQrzhIrxBL7SnUvyq9q++p6gLTxQdJXS+MnPOIJ9m5dycDwwbnCWlp
rF09oX3qDmb7QetM7qeaa7PUEVoYSHTacDzzTrVUqGqtx0WRGoWlL+kyzHdar3hK
mD126WU85Q2DFyFfZwnt7Wmf8UghlozD3ivYqoqVbdRLCTS1dLDgNivWMew6NIaC
d63LQbNcIXdsKRfzChz01gQusLYjjZ51arbj5XdSjhFxnlAJt6oBj8bkSWzoYXeS
TaDndHl+44EiTeHvL6aGkaVVx59Rm/viZ9LON5n4jd8n2oY0J6toZ7danqgAJyRi
Tmkq1orcgzxq8tsBK4742u58DATHAmHPa9FBgb6u4oanMJG9ZKU19ildzPLvcUAn
cTLeEvdtiiWQNYGgn/SxSckbLfMfHS7QnsYwDWHx+9fdKfd9bchuL4L09CNCWpwT
BmlykfCOhnWCSmgpi72fPGoG1OWY28TF+3DM5CT0MS9LEUfLcQCHjJWqKFmfGzx7
rdjkRRhCuKBE2JUxg+IyvrFkv5M1W6cpP/dSzkKpkjY7AnJIOCHvq1q75sAo5MWa
GRbc1JWqT+NQKE1TuggGn9vnuED1xlthnIMmHFbApIQOzRq/eMlINKYdbJ5T9ETN
ZN1J08sfCC8Kw53Lc+eK/W701kn8YBQxVqNy3zzE1bWW+/bcC5kfnVC3oP+mgPxc
6sXNXXAkljlNBQXZls2P1/ANim3Cv/u/rtk1wYbP1ckYz5v8M58Tt0epyPtwxfoa
ALRXgFAu4QdQCqMAEpjwhjcQlbnuBsDslep3Ca/WQHpg8DEbhg2HY1hkULtQwmLn
zHT7K6yZBeHfLlIcDG10GAEeAogD/YedS4sOO/1w10E08eyZEhQWSGrul4q+uAyg
fXwLPPg4xMKRsBdT0Sdsfafxb/ZPDDh4ZMrn02y/ulLeiHsZm2y/hsvqb8h0N50B
HgOm7l7ZcTvvYvSQJtOcyFgMlBDwDsBiiWuLhsnmk+/JqtfkRPjx6i97tf2LV+42
VZR6/8yLhtP2/IeTxexd3rfLUjUwdH3nFnNzdkwogVycrcTs6k7Wrc5KTd6vFdAF
uDGHop6swp3MT+Ar6QAh3utJQd2xfTVbUbnlMadZJ4feNtPMStP7MRHyRo8YAh2h
bkfQbUy/+bzhIDJNw+qKfgkvcTDuRDNnMpOGc8URRMUQalQ7gMs2C2EquZkdMayQ
L/aCNhMawgCfa9FuY+zMoZ2p0KV6jYYD5g9fRqpUizda6lNYSkbXT/gzzUt6MnaD
MrGtGLz5UtYVpi7SR4mBX74SbCOdW3nXC8b0gaUiu1ZlUnqAeuCFnNavR1n1JJfw
5oHdU2Sze679W6YeUP2ZnLZBn5EsxTWxERGuPW8bKcCHXBIE02LxT/sZTBlChmhf
cNwOaNd3Y3eFvTwVBFUP9zb4iqVapZ3LrDy8HoP5to3YdlxbjlQWXV9qNKQbNMM2
Q+Z1G1auOL54aXZctZyjAB4arnGt90SI+kJk4VYZ/Qv1DTCY1qeVxQkKZ10qhkWA
IuTyul/dduerZ99xUSh5u+fc16KA5L/GzihuR6TFGKLlg8PqA1T79T/bRhhrPWKu
NcHRB4ycnHNkYGb9rC28OONrbkqV5MzDZVemJSnlUvr5kIucMgRAKtm0RZW2Prk6
T/mcc9K1hJVNc9suTBUqLADyXQDzrEtz1/QmbDcle3mOOLNbC6hfE2EZK/7a8CVE
K9e05Dt34hJmpc6pRPEhQAv8yip3vEL4iweZOK6mzZ5hoKifyj3jZXQiArN+3eao
+qfPQPmgQP4Hg4ZoXSYoB7hLmtHO6s3OPLyXfBgDcMldbu5rhrYrPDJs0vap43xw
JeiCjeW7PU2QnJuUrM1498eTVudlrINP6W9z8OxXJnsvGJyGIJfYHS/IJ2D/rKtf
QVLQTtXzKQNTPxrDcNxt2rl3HHfoO7SS5V9x8dbpiTzElaH9c4bSCt85GpWna9lK
Mwhrk/Tu4KfKaebg77UQpZUNry2HIwL/b34ztLJBnUvvsxEoYAq4ei3ohk+EK2aF
3op4tWYDBTlXOCwlOm99FsAHMwEaqZV+mEiII1fT4r2Hgk04wwusWM31kC/pNCJ+
Ti10IBgFPVyKgcxHPxHTRPYyI+ddT6vW1OiMN/46qyeKq1miBrK6TDNdmSFWj1fT
o/F3NTpy3SD3Z8rLfZGg32pa1ODEnbMHUM+Qs4NCOiXdiUcxBskm4COyV/4Gs/I6
Sl/px7K47uTYTdzie1qThtdTwO4PvHTPC0h4/5jo4fkqBBJmpehAYtk1fhBwxT4V
JntAPUe0wgoQrcBlWjFOHA6i7m543SLV+HYeEN8477XqWA3vxeHUV5thQ5y2Qisg
4h6klkid0O4hERAK0gME/2r9p+DWQeAZNXFR8RaskwEk4J+Ulp77fhozJ3nLGT4M
bt1XMeGEXiq1G4RhCS5SUSlA1hTwloT5+80Ezc9fqJ8bQGCEsF6sj5sF1jAM27p9
LF5ybjnomRkL8adRPpP02oEBiXz97lOB/LZrE+nlxtj0hscGpCyhzmekA1pXD7Lx
2+kI6LTQIHVH64wgvCf1Rweh8K3vPnMpDoqy0DsPqyXiloXu1OPNpylTruWRw7Uk
S4RQVj7KCEOK/gE5H0oxKDvaHtsQzWBpkCrItsH5gJY6wqlSmlHRGrDcP4MAAdIU
MyASnc2iC5g8oAh0tbbj3aK/1uzQni75joPPQei5+x+fBNbiZEmmr3SU+aR1T8il
/vLsQfziGtYQ1S3Dj6A6f8M/iwTKQ7iNx/PYq8L2p06VMx54yjvcgI98PzAn85k2
yk3+IrtXVMK++kIoG1JY3mrF5ba2Do/bn3AzoHa1KZoVMF00hMYMrZYmeAt/jxSs
IyyunrLgWJ3QHqWfgMCZtxlk8fkiyH6SzEEzSGKQ0lIepqOJVhQjRiT77M58xbjC
VTMKb4emhGeCf91Br0+gGwue2o6RCyX+SOvIAa32Y9Dxj//hRwyYjo6r9sFtOb2m
HFbbefJDBtSG0SGtfWtajSDFZPd6IMjf0dC2R0WJGTFUikGYt7FjMRxufnEn0Cl0
kuNll/Ntd1YliWU4fqsOiYl2fwCY+K0i7V6ppnKHV0oV9B40Gs6vqNIq8sy1RmYN
X6U5kRDixWGlYR/beLnoWPTLLh5oYv0OdYnIHm7cS41ipp510l2+ZBfrDD6x8XJB
DxLgtfmO4UmJwhVXeMlTCKLC7oNQAOBpSa6Kwl+km2dqZJRbYwxXDemQzk8Bieid
5oCtx+WF1m2qkfEKbmLsZs6JQjw2+YSbVjoq/orLIXGa5fVyBWlBnbphKWhxTSYS
gMLqleVA5OKfLNpxA7/81Mi16MY8vcBrOPDZf3GrjvmUEU9X1YM2t0ZBelz/CdCu
u+SEMKsS6NCHs7c/GVQ71YfV/oZ4UgvMcJj9TrTuXLnEhajeakcAwIkpGM5I7Hjp
XG5Pl41z2nF/a2Ai1dQtp8bzg3LVKZYqsjHxuFWO5+PE7lfcfYEP9M13VzUzgPEv
zs9JTM0jbtfXOSOBqjReQduNAgCxUT7iGEraJySgb+Cs64ThuuL+4xDAghVLfir9
VpYd2UdO7TEoJfIu3nKwhvQ3a56FuYC5jsmEpeiNndN02pJwtmoL//+lhjuqF7/k
uP+wbhtXGCDd65XGsF8BQ2MRx31aNLhCsmcIDe7D/vr2UMJapuw4D3Ifv+Ofuw2D
abKlxr3L8dn97TGspkw1LLQZ/FOPsNnBxyBGUB5wrI0mdHe06dJnDKuXZM7awh65
SC9IKDH3wxkJdSc4+CRatJ5WCW49b12wCigS5W9+KNgjJAI8225hBTmc8WR8Y/hB
CLaTQTnhSoUFUhdiFkOhujHUb3wDZph+Lv1zfXvtPaxfi+uKbRpddwAZsqtbzu90
SJOaqB2UImBVWe3q6F1LcYHJefTL/sYbI2HFFjzBsreZkUfPNkCpgge0uq8oP6c/
wWDFWOSx0AIBeL1dwbSAnOnBJTqEyJRXGi1ENOCeoSBZhCOwQw6Pr9lBUTA0bHs8
KcfYtEULO0DaFole5DFGVuU+YdLg7gl7aiv/gwr5sMM2QTXuuyAqPcQFSgOBHtqV
lVirVuuaiA0xUuvr91cYQnVXczpAmOibWkioYiPlZvTr5gfnYLpw0ErC8RoruClF
KoEIwf4E39ET0DHG9CQz+2TYDQ4bSwLeev2hS0cq9IPpKk7YV69CZb24Ugj1Ohr+
tTfEBgUW3+qNN6g0JItLCEzKotj+lr40rPQwJeKMylK6JwZPZFLwDy0P02E/GYKm
O4EZZUTLz/L8Qhf+4o4lFW4C997CnuiL1IhmBnndtiaxvY3bUVTUoS7rL7cYXjUQ
lNWu89DHX9tjRgLKiRb/TRLaW3npwUUTdIaA8LCC3jLb5JaHlEcTFsycHrSXzcgy
kYNOX6jenZsvbUSbICyLi2w8Q/l0mmmwHrPTenLomNvvI3UvXMyiwSMcOimyXmOi
kjOp5Cn8zJXciSdTg2V8PxUPCINy8kKAHmPdOUFUMpeqcXLfP6XRH4VnhKKN/13+
/62ZK029JT09k0CDMDMM/N0PNQuWD3ojehUYL+ifVLtPhXd6ItrfrGnF3HpYtiR0
EY3pHffzm1Y4gPmli0ADLKIh/kYhHbFpbR6h6aX010xApkc6jzV/+5ylj3UzkDVS
1dmH+k44o48vmFpOIfnpDk83Bh/yty/oaDAPL1KCstaZhB7LC+MNfAE1LAvKNMXL
pNSiug7ur50DdP130sQMziENzCMPpdMnC8tX7Jiqg0Xz54Mj5JD4jxz0Fns1wQZI
tDEBY6pan0+ehZBLxg4QiZbQtLA8K9iEiAXobe0vYqH66t6PV2B2bKfp9/09zhwP
+Mz+UTf9qF33L/PZT+octtxkpi1OQC6FkQQGXauLroRrCtN4RNNooDADBt6PaH26
fS+zw48NcvhO+2WryCjQtfF+oB+2bozJYJ2f75ZYQy8rSc+/B940wVwr/BGyYUbX
FyYa/C5/GpWeM7rrLQHg2TMqA7Kt1krEqHZCIsV67+E2i2SdALRvdURKDtATm+5n
x+t4RIyZ92IH4BCSRLoMzMTgotgNcqsyp7pOpfj3MA7P4osrray5FSw5jt7ltika
0Jq+qJYPSd7phBgGYD8Ts6mUBBADynFNjRX8bqSwGg6+knxqFfd4JSEeIwoC6GNn
rvh7rOKXX9zKzq30YMA2IJQffqMFvT8F+69N9mkNM4zryXW3y+JV8UqD7MvDyZ0R
JPRD5wbtSauGUD8a2qb06FRx0Pm1CC4FUoUSSyV0NcBMcRY87jLXqlY/dtc5B2T2
3UDXwQ5GKNl5L+ZN5y2DvQ5uXLU/VVsVcjpirjQlQL3ITtAeFxOD0vvirHyFdKNj
dDTndtvWLNAz5zldVPgvalr30UX4eswnW3cDod9EK6dDScIYvMnHi9I+gEtozzTc
8NzKF+9+MGl+l15qXkjsg7yCM1HNIr4uA5W7MUHw1bXj7DRituJLc6ye2urnEM/y
UUsAIcR7u5yRfuBTO1nqOgt1IFC0fPszXacxpMmvx0sMw61dRqsQ2WQIssD1AEvu
Bh1j8Tg3X3dLjxtosmjYSRtDQRKcJzPBbu4RnNSY5nJ0PQ09rUWt6Bm5bu9vPeb2
4XEFW8DOEP+plyq03XAhMR+5rLSZjewnjVhmSLp9oysK6gNf7gGmZjR331gcwaa2
3NwOP6iSsLYRccAd1CPoHRuX8cwMeGlnLfNEMGmA5ZXyyTw4LiakPy2VlKOdOIgm
paakMzF7OMwcmIprCHeEBi42lfIr785/ZPnAbFWpDwRu5htNrQtGXw9iuiPCsoKD
SiYzR0wKVHbImAZrS6Av/9fR8gEd+rUFoJ1HSNPlZpZGiBll/Py9S2ezEkS5IK+k
BugVqCu4zOMppl6aspEVWt9Ef5x/s3G+3adYhzKl9n4tfjKCMcg7nPRvNP2FD9yp
N5YrWKDARUHctN48gzRRuh7wnKKfnJRpsNKM3zVKsUnogAmwjUV4M2JaGskz39cp
Bz7W3uoHDreztHr31kyqZeSCDiTiCzSwbioFkPJLIJb2VYEqDCgtwPpHVOo7A+Vy
XGpNR9v7rwJQyGeXrNX96kvSK7BwkbbLxOTUki0pVtu4C3iFbQ1plDnkbaVtqVmx
DmJp8a6dvq+d7pCYf9+j2QEdPF+DyU8zz37t63ffAdo1pGeNTkE5rzoW6sA5CddA
wg9Qfc69lSATJlv5/0sNjbJmWiQBdS73O8Smu+Ayoekv7IxGEDn3dlVLZp09sX2I
ExeyPr0wkKPA9sgUI7kUkbhNlHgfjqfA67CUkmN3aseYh6gVOYHtc80fRoUXQH0Q
hRYByLDzpgn2pXA8k4h4DVpQM7M6CYOjC5XXfXNETMkaa16wPC6RkzY6Qwo+Qz6L
BQng7KuhdC+9cPI3R2e3enQvkNMFlEfLNIvMoOYBZrZEf+ka+Z7WF+sRJsw5vpWT
R08r+FVjer9Vh0FPbCCYyXwTK6XPs2Wqv17iG3d505SmwH1R7ighsFMUIvZrKAEx
Zanjt87j2G15Ew9jJUDikp332mMP8fChhFscTP5U1OTYo89RY7qi1Qk3tzqh8qC1
rVAZxMU25ZFg9BKwsrEUrtXM4ebP7/6fJb/int43lfYGwBv3EbOOriaIhH40OEkB
MZCW85ZWkGLw6cR7qx+JqybxFpx33kju9GEHdkurIg3eqUAQNbAfNPUQL+94LlR1
K8sCT/dps9oy9/qPglyShEFxebcAnOKOF79UUarrtJBEagtIF5XhVg/WqBCph6L+
wb8VcVbblvCq+GjiNTf5IPzmeuPvOgSrUkdl71gbIVE+BoBZ5TmskwTIboQWSHo4
BM+iHoh28NNVTzbDozXyMoqpne9qdNO00nygwACvaXkFWArNHJntn5nRmjuWG+/R
3/Ox/If1xzDOS3EcMLUXpwB156RfIfD9zruRN6lBh6ngGGAGpf1J5GuOXtqYN4N0
Vf831Yoj5/wZ2OyUWh1syobitISUazxE/tMNq8OnlkSb9jfrb6dZpI2Sm0CMFT+E
IYAk8IB7wp4YABCFOE45IgzhlTU4MhnVbcqqtm8Zxq459xQ2s7rAyZV3h4SWz8ed
QJPsqtXuW3yKb9KK2VoxoPF2wIbjzNbjDvnznsplvg8l7R8k5ITQfZrFyj9CAovT
399kf6sHQw1hd+vxBG7ZUNlqhPm2yt/6x2vDfydIMh+5WmQE3FYq9WkUmrDWzN+j
4QYP5MM/dUpKMm84v4TWV3KVzQzoVuRPoqCtYFX4qCFaYyEuSdccoN3XZel6Q5PR
c7EhGtvp6SZOWnuJGTpwNYghqGeuz5SkwWwEcizxNJvf338n8hXclej3+ImYP4SI
aW9X+wz49q05tCpcxyVu6j9lrp9QCL7w63ndoPtSEP3uBVTGuvPv64kYxBfSh8gl
Qe5QKipl0sqSgHxLXFIo8LMbXglWIJWVqKPDaZKMfYQ0xUzcSdOUYScHlV6VexDI
aAWi2suPVO+MI90sC3oVuHGAH51+MzdIHp3KBgx/CT29i3bvLcAY7kdF8GyeZK8m
xJR/69Ko6M8KBRJa9mHrsSlebHMT3LUYvqTDbsB/LDquWc0ZqdWNuHGl2+8XRagR
TheK1evDdNcyYcOkCVwgwVXb6P8N9P22SspnDfmNpoWRkiYOz2uNz9+beW+nxDX2
RG+pbbAqxm4MLPmM1JxwD2CNfPtIYDmvb83XUYURFCV5/TkyPQc7JaIwEfVl+VJR
x1HP14Dv7KPgnI7ZC3ah1j/sJzhlEu3pkRq42Kve4gTofd/481k2GStzJrT7P/5l
62KiQHTAV/vNOKvn8P8tWiwXl5w12m2rt45RIT7uQaBAp3w85Gfk02fX7jYNOwHN
pKtDIiWWi1W9voTk20JBZdfK85pBA4LhcMTvrB7HMlA3jMWKhy6l/uNGg52550Hp
sEj3BlMHmB+sNYRu3YrNcKwf+b3GQTGgzPnPB5LUPyNQVtIBNKEAfXxCzukCR8VQ
mgoQL0T2K8S3FrQMVxgW8DofoDyPeQqgvluV8k5NMSyJHW8lrkW7J4D6JOqCENDS
/+pkFDoOAjSpB2I/WifWTSEUrjTFzWVqO6+3SnzdoPEoOEauSpWhHF8ePMNBNY/W
F9D5jlcjH9Nwojgh3mM52/ySfNWWCagTPKutiZddFSm4b4kK/rJZB8zxszjVYk6G
wcLdi1aR8gSW8/vQFEfO774mMKbnqGx5pMgCvj2qJte14+urA0vgA27haflui5GG
atxl+VgMHaodPbNTT7OMNoB2Ps9w/HavwFfDjHAoEDO74hBdAXlbCtGA29YRMayQ
UAKQgPDV5RLKGpn/FFAQe5rUteOx0n1fKZ9SGICrjJATXbU+UjH8k3+vQvNSmiXD
fVqUDK70wI8mzeY5tfjZ8FGRiSm8Aug/whLqmoWMilUGiTy8MF52CqEseBNiVNJP
Q/sVlpsNFDBk983FzewWSsxZBEe6+6VQR5anAnkGYoLiHxDyAh99hvIEmXgcMdjF
SKJ042Wfgh3Q2eFVpuV+bHFK88KYHWv1noozB9sblMjyCwE0aK766Xip/yM7IUba
KZ+pb+pAfl6pxb5zlT4lmUaMV82uL2KGR9AIwqMHi7E3cerPDbtts9utiw6lrI9d
HHUSkFDZfT09B7Lu1EAfQPbdOjyBoEQYX1eQKfpXgzufhcB6vLA50o811dMn3RHN
w+wo+KQsSDgkAtwyTYXvQdCndcsAmtGyDmtGAE9dMd6oCCQi8k/f1ZJNm2loRue+
rbvR3WMz7SyJiAr6tkEuz23kRPhKhwh2QYjQRSti/wbKzgnhd0rlP4nHw6xfdOqf
d3hcooFwD5oJbWx5UuCZabvLjoTVH5CdqmNgv5C+tKfvpkSrZ5alze2d/EyvndBe
df3LpJG0iz+Ck7stKrAfSAWY1IGF1fJ1FqYCrM5yKHX0sflLJFQyy/tjcovk+YSs
dFPvIVNgAiTHRZbdic2lSmgKK8s9VManzUSi6VZ/HQk0i4KDoE7E1YE7yUWYNQnz
7FtdZ0VsfsWuvNRj9UiMtWFqBLo1tl/eJKLl40xFAOP1YMZCno55aMhWPv1XBIfe
A+E0EL/t3Scp/qsYXuU3lnUExd2BqlZKOck3V7wJGeQoS2mKJBJZKPL0WsiA+4eU
qqunXuoq96OUER0+djliJWUz9TXzbTabOdetvEBzS4zLA21nrYNxX5VOIdMg6tiI
38PcKGd9a+BUAAaSgHRwP+it0INMLKMds5dzSc+spmXgMFhmJaI5FwU2X2quMDdT
kl+HTT1o4WNbK2wVbnjkpKOcumbyfhjmyVMsvun2IXcTlyqOpiPHjb+DsYZxnjyT
nDojYfwpDYZio+OKI9vYH9tLJkTj1K92upjR6Hm8uNn7HEk0fG9KjNh4TFalKcg7
D+MuvdNJ9gI8HA9/xm6Z42UZwtGQMZYNm6SpSTEl/GOkPaccj+wI3t90/urLMuRb
uO03+FmRTuITYH5TqcE0HJ1zdieB+hk8W4U8xZz+T5dMksIJ3ARtxVnIC8+zTRTj
eCo9A7C1lP14u5rwDubxu5Stwn8yZyozv5o4mAtZJfKJlIQ6UuElBPNaaaG9biL+
QwWzqNR1JP789tqOQPbLKvwb79C0mLq7wCIAcoeLiWV2ry2ApJrcQ+IxJLy7wLmx
H8b8xuVM7RM8sLvh75zUlRXkb4Len3S9Ke0sH1y9d65rZ5ko0SDtAzIfl6Gl/ZcB
19xg9ylqlxrhsu/7WH2A8S+beB+9UG3i7Vii0/33C33zqwV1oIGwMwkWj3GtaL5X
tRCBpQUTNlr0NWoK3gYpUf3xjpinrUmlZxCOH30LjDLenvfycdNkFOe0jntfJmid
NYoojbcf1/4hPpwucfNaXmurxvE89LrddGWjB+ky8Zt60a3qF827zvRZYCWwh+rx
/aAaVzUfkgGA7jUihnzXvHcz4JG0VuTAh7MLCAinYv7BZzPQoX38rqWYDXNdglwP
UDzanHYym8YUQ0SJs0nBrjUP0Izjz42tbMfWiHLtGt/kuyZwXLg+YBV8iP360BcY
v5/PjjMB6n2epuB3w1/+sWjml81JnqMRRVZtcqEzrod5gjJQOcqAImuOdtgNEqfr
0OPZTGQr3HiiHgQb/l2iPeqPZtk/P/RGqBZQ2zmNyD27J/NncyUaEd5p8BzgECea
G2KSoDaFXrM1N7fLgxVU1noV2PU/SO5PIjq2oFjKeSG3t5NB2/vL7mEy499kdp12
otO3/2N+hGtDY9/N9+MkVw==
`protect END_PROTECTED
