`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QPHU3LAIu8CkEVvibaRLPdf4RE4Wf+burYhykcjFoUtcMtKBvfgJzMA/sMSwW7U
I30Rf3m9e1XFAbWN0/K6SaXIYxCdc9f9LRLng2JU92SHtXEATrgrvO5RNoOFQFhI
ZIRiu+YmA29Y5OEvUV2hHzvgofGrYPk+uyCkQCskDNBFL1W6njVk/cIgzIn4xi1k
wBiEgNn3NvOJuHgg16W05YZfx9lUV09JsS7sdaC9CmRnGrylca1PRWFY8j5VGdTK
C8zfJ9hdI9EbgDxsoiPODH9IzvNIhPdGdmHvPI5ALn0acwr1oJr9e/Xx2usU/fkr
DGK3sZYIdY//J3BfEKomQm5RpCCz6XNKhZQMPRPpn5QU8A10JJmfQCWPeOt0V/nI
8r22fQqRyBfN4Gd1l9cb2oJQkAnPHB21BYEkIyNF3ruJCQsXsr3jBHrLV8i9qmxV
HoOFlcD+K84UZ10d0hbgr2SUGzhQoPZkuN2lYZqraYfRVcXn3k73tLt8PkMtP8qm
uLriRLKP7wYBKtMSDi4AO74gQppMbUdBP3ZdKzvsELKBKeGVViRgRrG/rw0fH4X3
oG2tb2ivWb2UqHflkO3rkU6o7SXWSux2v/sVgkn/xpf/mFnx78DkHeqQ0nhaNftD
Kj5oyr0af+vi/E0I+ukgfbz2vefKzFOx/41+olOYMIkH7p3pIY0xAlHXLpZJLs4m
BM39P/2HyYw/w0XWSd61pbOqwMbUHVIGV+FzHFUOOP2b+40xEHSY2+UotnUV8YbT
1MY2oA24dAD0Fnq/mu1DDB4dX+agtmnlGY2ze8xR/0QwwmWy63GJtom8HGcbaH96
qKazuQMXNGDbSYZ5AhF7kHN0AxcMWGnC0DW1UWIP5WyHIC5znlfzmJl0rCYl/Mf9
3WVradHBh+eK9Fyj+IjCJl2VOn8qykyzHQHo/ZsyG0YS41Sh13uc4VGvxkx9D/6l
n/MfZXNscaCRVoTo8xrB1E93LIFsFmEf7HP2JV5bQHlEs31oMLRhzdKAi0ZW+B7v
x0RcgxUmvZJzIyJmDx5DlV609y5ydsfW6YsJ41NAGY7KlG7J3Cbz/zOq/p2hLum/
fffWQiIQxQLarGai+BdYPAI3UYbKiLkT0SWZVLrOcHUTClbfd3/jiF6VsSgNir8A
J/qNOnzKR3fyhxMRHp+3Hmay9IPvKQsfDVISNrqh4SxfTvqlaEc/4x57E3EZXvru
KjH4jSSwYxCAAeeDsxaaPht1ESxRKZ52QVeAcOpjB5HP0Bnv3bsCBmPjEanqqSut
QBd7iKqn+F1Vr8B7NKLPMsDQW1L5ENItLc+LSzabSAKFgNiULTI7Hr75rbk0zwKj
hIJCCfL8rmM1jnvPyrIWdP76jxGkfW6OJanfATEadZK1/37MygHeb4bQGsbRjhiS
txha2ryn2UcZDLY/n8RppEWH4uf298N65AlOK6Ilqb4qmUkSpUNuCEVO5Q82DN35
4JoqgAf+WZQcVwh4otjmDciFzvqRlH4WJ9i2ElwmmJa970wimYrgJf16fB9idYtI
iNWUyMTuocwQnKfL81AsdCEJTPE5Wr+vDLn6t/rTn/nD33n7jflPKWVL/ltDF0Rv
oDy6pNqSMSTOZmwsipWEiJRGdQOoDV37746JeJdjhWPGy+J/ot8dmrWLqzSX42qt
IQ13rTMCXrN/GMk70CFlqwcSzGoCit2rr8N3TU5pJCpD9+CILR8g3odFOQIGElsr
nskjI56Uafs2M39ELeZ13f4zKsuVh4lmOPovGaEbaW5fA05NswfWSPwARnq+jgNn
DPmxCb3L0M3Sa9jF/8+kRZt+ssHHMb8TCilnBnc+2iqPgiv1r5A3mZLY+4zspiqM
Kbhueuqn88Z9oMHMhwoSJAuP9xZ+0ZGjRnbNwSNIJ8QDr/WfzH+VuBBMiDFp8i4w
lwyTGX5a7ggIJspRRXA7RcUtutO+7WZD5CH2N8FVUKIX0VbuKvTzdXCZClJUa/bW
0WD2/PDoYKAhooggncfo6RayYzTPmsyIv1SjxbHPlE06E8jQ5VMqpbF9Qfp2uXvM
JuwQ1TmYSnRKqIO0zfc1onARAWBjTK2c5LlFFjQABIvDJZTNlmkSDyjidRXUOZk7
X+dtScrvW/wHNANKsY05Pf/xZCiYQ2fcBPdFcTDcVG1MQp39rHAIGRu7ScL0aHG2
X2Q/o0GX0A4EuAAkiPMCx9dgUdZ0r7yNMaKXpm8j9ipJMQFp7M7cKcPZ1f0azSi5
pQJDJLYM7SeWUvx9ZU7ziOTR8x7XeZNt6uUuV6GUZjr5MrI+LoyNqm9/JkNqDIGD
WFKX4CKc8HHSMB78zw5BMkf6aCRrFe5wUwJOqFRm0tRGubztw3rETj0FMVeglsSr
D9kA2GQRIJBaiwbe+vPnKkkX4CgL5dqfbrKWTR39h9h6MoGe47F9ABDqXajDQWJC
tQHEEfvFz3bhRMHKS11g6bVcnvFNrRGmNaubinphP12/Ikiop+Xsu9JTR/uSvnNE
HR8sYIFExFA75J5hJq6yVKOz1R152NEyW+a9PpPnbh3OyE2Lms6NdZQyaZa+OZFV
xt0uY3ncuNmBllLsb++dh7y+FOMwdR7Tmc7hPbwd8PXOe1c3kK1FLDaitrYuisj1
mvqnr8dbHY5CN0eeRHiCw1TEkDbQcPUUwqP2ilDHnYO0OM1ytCPEK7kgzW2riLfH
qkdN1OuR1sTQJXr2Ti4LmTNWld5Gzbl7syvPMDEKLl9tKaPsL4NLTdQ2pPApHRuF
qTA4tI5ncGXFLqu1CXoidXT8sfKxA30FZa4HQDtCedDpSfZQCQOl+7mN3f0aC7El
i7eyy/9ETUaTZIO68r/hHvaMOvYG1+pk2yac4CCTz2XN4dRN7Oug8AUSOkQWQ1q1
U5GQERngv8aw8ID/203LRPa/QgYclwhK/kPFo/643nz4IAznWcvdXPUeE9KxM6Gy
f5YdNFZwhPbQITHpUKOInXsB9cvCerP59bzpnvCbGJe/EhrNrXoFJirzob8xR13w
rovUaUgOpVlxRIrp1jPdRc30x3Cx41GV3lbASU/lv0WpORVYaDO+4wTzGLzLpDNY
QCfc8nfsUvbaXXKsreZKYwzNyyHKB1TSbGb76sgz6biIgu8Xz6HvuMb2TdcLU/es
cFa6oNDFGU1qGIGBjFMyVJslRInfp6tmBBYqPg43f2aphrxP1Y8W5Sa5B67sxmxE
FcKn9josEXsxpruyuWP9dWerc9vVEEIXGJLL+PH30BGd/xIvB9SwEoSjXcQQvjYM
isAe5wVxNfSC03DfDLaWluSZNWfWoNsQvIYwBnwupmWbmRVftPPlLgT1CQFPkjrN
/iunqMZ4Y+cXtdjseC3biVgCjFdEFj+ha1ZgbjH5v/Jr2v5bTL77KXpxCdGlfv3K
Ribc5H+u28vExl6VAmv+pCLMAuLK7PENnoC2n3wOX+BcPmPo2rExld/4kzM3s8CW
zhKppp1he1dPmmvXcxpevWGJ0OReU1+Zg2ZiVD3vvCMxle9gk7u1wNzhTyiz28u0
J8kZiCq5Su7+bzBsfaEpTb0cW/9wlk93lWjDlP+qdHBIS9hd7RgdY3e3b9S3UlD2
aOOs+Ao1LP++oosRf2sQ7EXIj6Fjtj34j9woo/31qX/AV0Wo6p8N09xSgy1Fb6AD
bbwXQAM5WDEm9+/dOwuXxk7vIZFqzv04On4u9AvCBxZBhIm1DmjyyIkie7e3uydy
gQRoTNLXdjfANH5nvIX59DFBmrxBFWhHuKrkVNPgGnHJtc3irPVXziWAXaBrhRgU
T88wETkQEyP/ZnNP6YRoTgXC0WeojDPvqxQ+BGIj9sOQqyWvpnPao3Ouqp5m8vML
f8Ob8YbRr7e5Eth8zWhKfMzGI1XidKFxx0ctPCdW0ZJG6uYZTEJbRmMES6mWHruj
7QcTYDZu773IHbsjPLbdCIVOIpvtxh211z0hNtKfMlM3fvPVn5D8vfZOnsqyoCZ6
Tso8O6SC70m61EpYXO7C2wYf+mL8hL/ZtjtVz1BJiTptgbOJu2rFxkviBnXxcC0E
EkUjZwCu3amHFRDw6iSbsAZH7stUnHxVvqWjifjtwySCbD63vwYOUB46lt64iGCC
uaOSgk+3F3PIv8Ai0ZlnsucXcpAL/ie91V/n5eCULTiWKh9/C6AcVOcM0syJeZeQ
0iKonec08xa99lwNe4VrYfsX3FTUXISbnBnUHy54Pa5J4pqMd2MrAGIjitgQSimP
df8LAgHzVczWMqfVFxhfDTltphaBVByBFtJdAwjZQvTIOBp++fO3Mir/4qT+Igtd
H1XXNh1exQB+tOnzBGzAISOQ5jSCeCgPDTzCbkzeu3F9b+lTvU8bHnQGGVE7qGfX
LGKhIb5Lhors0gO5bOG3tE0LC+ozY2qwOcByp7GIvLCs6K8BQf8M+Jx3+38zUG7f
4MxDKl/snJh77k46HRu0rNXryZx0DJTt4yGu9PdZ8B3zHPy70O3QqUsvpVyiZDBW
iH3p43H+v+goG5QXnigosX/wbHv7IOv/xZF82tHnd3AP386VsbI4tnlAEHRQQgjH
KRwXRsZ/bWcEJgnG0EbHHTccY167u4AiQUW/qVqUSRYB7KyhgNGjWiGRvLIzQw8u
YXpG03y7qh8Q+Ntac0hLUVBHa9wz89+ud67Y//UlDYeYjUMQBoCWBoGxUHHo7EBg
I75Z30RHoDIW3r6Uw9xSIw9rn+gc0FmTwlbgJMWRyU596sRRKvuOgqT4umBkioEL
DJY5EKRljtFUGmb/LjerKhJDgnoqAz0P4NJrO3QF0ThZJxE2S0U/FkRlB5xF4g7r
j+QkC+QR08HNDt9uOv7wcW27nZUDNW1uTKpVodeQEa0TEhIVnRYagMqO92gw6pdo
LspqRDhp2GrVwLrAkutde3J/l/ZUh1caVzaeuUiqPmriv7pMO6HO640UdufNCLkg
AQ1uSWyMcPx4KewI74KIQnfyhWnGCHLsNley1HJO4KJ7kvDq0hTHpGwSI267KGyk
yFKFqGT6p13TUf6io9CvC3wn5uZsJ7YqyfG7i8pGk/i+saDXXuK4RvrSCOT4Vhtd
Q3/fvSDTJUzkG5Tq1/P3D/KJ7sFs45NdPC9HHOwzHVeE7hZNn3pzGS0XS/AIigSD
mSC0H5rwPUqjywTAJx5eLkpBR5z2XLFG+niDy3EDm71auxf+2PRT/nJaya4L+Ipb
szTVR4ITv0uDrluwpa0sbvA5daofZCr14UwooxuDPEMqYot2fMZasApdr/sLeN96
pcZgb5Jrpdpu24fVAlZrufIs9FLjjq+5YxCQrv529LYUeQdWPoBMbwp+jtQCX2g2
uNEZNgt76McombWCDjGqATa6Uz7Gj2bN6BkwiMOEiUNn5gMxl6jDLI++ef58J9LS
3r9MRWfHKt+/Lr7W0/7bpPLFh6AGIbUSSPgLnbB9o+KjPdOvkbu1pZW66KJIksjN
uE8mHsIhOHmoDsqp9kWTIMinQuDYxGXjuyRhCH60hz2hjGFRNqgkb5hdmULj9hYB
smnVDPo+UC7c2TB1fApnvJa61us0AMYUwPadYzY5MXJ6aartolQCtgyCTl2ofcF4
24doyMS/W0ip7hx4jNU3vOUJA1Xi4w+hFy9oI8fypAH8+/zUhgLzTz05LOQ5aAkn
T5yVISkLmjQOZlgi6ghGDj2qrzcv4RKJkKNoEVqh1R2hYxfNCtVKdjHwhOF2h71c
+GcIZdNEWKxKAniUgvSfUoQhvyMZuhL19j1pmLz8yJQf2pbF4WTph8oVaw4Sbj8O
V5WnaeajqrEK2UaMzt9tp14Cl/PmIHEWTkMnxo6vHG6MeKS4yz1blWKFMBdXYlnA
IEwPU4JezVeo2tyOi020AogjnaXO5Y9CDTkEFp+ekM52cG76/XU53T03voGhmlYb
fyxSOG2zDzv8bMqbMVAxZvH5ZPJKs4VnrI2n2JVhZDVEP1ORcKiLF1U1XMU4pb8b
H1DUyVlMMMI3TeLz7P04/ToQPyQV+tHmVty3zvappMVzUw31s8jhX5U2ga5W+qn3
qDWCsxI6TaODBnuq3E5nnMMlNAf2YhQCy6+Q0TjOBg7BgsiS6wIMGzZXYOMDX9NM
n+Gr1yUi9stVuMa0Ep90Pc7eEwsnDotNmcJsDsrSPUXA2Df/0fEaCvPG6B9IaN4T
mhXFnxo0kN9Yb4B6AMdmgyN62glLS8XN8FCPfqZSVrsdVXXGdVuikiHIWiPhcxUq
MYhaoQVRXnaUTeO5dhS2tExpB4Je86ujqqum4aADH38hGDxu81YDg3aiSWNyihoK
/E7hffe/sqe6qCpHxu0o85Cchnly3JzL8ayRr2ocF5gafjB+qwrFtxDRWQ8i4dbQ
UWjtX6NSbFPZWks9r/MLsdLj3Pd/1ZINIrFkVt22cFn7H3Nba/Bx6m3VZJMQYqXn
WlvbIkmF8J7fiKpPVlCgckU9D/+HIFZoqaiQGcuea6TwHVYi4U55Jr5T+MbxjwBe
eqpHJo+sYUufjimdSFqoFpsDMknFxIWPz8SxuXJJjw0nCEFxXA5Zq7Jj/Pn41bI0
3qwcFDkuefnrKSZ/qm4CSkwwrPeeJ2HxFX+SIJniJpDF3X2B1DeaHLOzEjgIDH9s
so4igLg7kYsaQK7Vl+oWC5fjjxEV2sTfPL+8W0I60kSQWNthChc7tE/BPFIZUlWP
laqa+fAhr35ANoqilJsJ6o7JQ8k+nZIx8mzQ74R7nj5EBCKubHidrls9TlVVnB2m
TWVeL96P65/zsCUEyL/Y9TumSONgg9CISALGO33kWlEE2P8w206Bjt7rvuEl6MkS
ylUocdUsHL0J7y6mPr6IqKhLeSdW9H3WJvg443Ru1lCA2hMQFDx3mA2asuE+EMV8
J1xDiR3Ay1y3W6zXZ9QciPE/niwRlQlLUaN2+ScVyAGzN2oll4FQ9UvP9W2937ci
B8URVs90+1XhA9eILirhCznKnxYtlnIG+OGRi/XGeBM4ZldTJleSzcLtg64/JIUR
xY74AkmunwE9P0262m1+bmARXndUBeuXl1DYzVHQQBHVQ1XcITDnpHr2tSbPTQIF
M7IYa5fC7xSgXZJ7zGBJDL+JcKGtiuucnyWeRy84GEnAKoKG9v7bfAmDGqzfQpun
lZW4JC8nDHaRjQQGZzgqKkjjWYBXTDvlPKOXq3dACsHxESogOY5E5bo3mcW0k4dA
wNbpOHIW/9dprIBcvNSxs5CtAnAKyI1YFqEtGJMeHLEBhrG0PG2GCdjIWYNYKEyE
Zh7fHhn+rMUGR5LmVGlpj9xo0ThwNMTi9K5QDtqC3wv+b2XZHiXiPsPmDY6mkwyC
JrCVxuj8U/wrDZaCQ3DDumLfRV2Jh9deIk5oAmr4TYw8/ahAn5lZSG3Uq1zARwBP
SQU3y11V0axOepSX2hTxskw11kp8eFXsS7ssnpS+pCZM4fYFtuLuFGOI3myq/9ex
jm0quTuG304Uqdg670NXj9kC6hgyf9VIXE7b50bhy6Co5L3laAqcKDC4wASvq0iA
EDPgDfutHsxY/5aYfvDjdeNlSIkz7ufh6lC43+wPHysV3YMYDNetiv/aBMUFjvRn
p0ljUvic0FOnt3kqSKpQ+9bwoiZL6KoH/mcT81Kaj7p00TGZKAK6MMSJX2yGZ83/
qNr2OMVteMrr7/qCm4IDqQUU+eRmpEhyS04HBLmx1wdlVzK6pQKqwpwpOXfgbMGp
ZbUJsu0Ne4NsRYdx3w6jj2SDmbyjm+uZAMo+JXRL1Mg7eQ3fv1+tJlYL7j5kNpNy
QuIcxO/zkLATkLqvwUUe1MohGc+rJmHL/RHxcksQBOPsikJjX5RBcqKJYvReT9wj
fGVwM/XA8hz+hFCIV6WVqezVw9gRnkvIw9bxkjvBUdOglAFNM23K1OoU7mQWO0tn
Fj+uQhPy+HLe3X+sVdg2GNMwWqDA5Rt1eRXhM+tE8cmpzwzfOgO8vZjJYl4FKBF9
dqlst4w6IsaSwiG/7Gg48S28itTTK8Y68rvfMzMaV+iK00puxT3QUiBU1ikaLWdi
KhypHUveS0z+aHw4Cgu6ilDKLHNfe6z4RGiIPlkV+0vd9gbmtSD43z55J8DmPFkY
DXitJXS5anJe7oxune4df/IYRToyrz3KmrqdlrbV4L9YhCyNDJkfH9qSNQkzTFat
FucaAG17nFlK0oN2U5wD4elXgQ5Ut7YWHbpuGahcqx6K8/Rc0VV3/t8TJJO31/MX
RIVS+RmdFL5shWXfpA36stELikseK/3WyLLUiV7WzGI3vHuFTl/koba7CPP/whud
6tjEHcjMf1GExe6EXSt5vvaJZbUGHu94mKm/4H/UDhS4JTmZFDjD5Mii9MyDNOKY
SYx8EWm/6LmTgkWccZ5RFbS0mp+zTFcviJMNQAUPRcCdmMNFYvEpAoPWza0CfdvQ
wrbieeMjZFhjhDxROuxxltm+4BHrBvB3IlK/hcwUVuLSzLrsyg9coYroukiUe2WC
Hr6KUmZC+zDp742klRNCDGzHw9vecqmCgUeNvP722C6gUUqz8w/c2gOc8oKVmaIc
YCc26po1zdO+45rSUewDtTrWJ5S7OBHI24xzK+/7UMC/Vjv996XiXpwV3KhSUP4G
cTVLRzWF7ZIpL1Ox0QAlpzQHnyli6su13HAXf4eNDMQpzOMZ0QaYagpTLutBz9mo
Ojwn5wkVKAkIUcDgQ8KzteRGffgtQn88xlZrTL6fSlorkzp5meeGlF1+FPLcCTjm
G1jeRlDzO00OiYJucjXKmVQugH1jdE7scd5OodIJw0PwnCSWJ39NAjNtPeMqgW22
HMQzsju51GlJ0OcAjtZ7Jvh0v9ZiVorXOz/iw3LeUUtpy+RXJIxEY4LHaNCShs3z
Z1r7JYAidSyaLLSSx5/+a35rNyxXVji+f6IsTf97TB3eg+SZS7o0mXrBSACpk4Bl
XxyR9+aooB0JfpzYDyM7sjxWxvOzFLSkUcT9dgArOcWSwPRsy7x9AzDH9BgMkzc2
e+O7/YjrNHZPhd0pAvEIB2FoWdGNIua1d0whkOL+vemCYTuBkKO7Bfwl7l3++iOr
PHQkR0xcm0mNFzkoaA11//rXu+CZOVr/KVtqYxz9CeeHtpKSABH0NoxnLfAb1TVy
yTJqwFoqSKQCGacNFagbVFAE10AvaAm3sUDTnzTAo8YLE8jC2MQl1hrIb7FaSLi3
SHZS4zNl6DTpj00lWPGxA2yLCLp+436BxMNoEv7tzBU/0DMNgN2SJEUs99oLFkb5
UTz2YyFn4yo/pZihOoHAS7qM3ErnRRmBkxhTEhkWUbAq0px2Yq86WwtcxlX0X0l5
KBLJSTthV1qaI/din2URPF5+zvXfUat9dPc6ovPwA5PAY2PGu2oQIIJSIe5jmRSr
VFgOsSv/9iI9WLXntheVAFkzcXMA52xRKtvZbAUnO1ySpM36SrR0A8zQy96cmSXB
xPnzwv363kyKVIWgUekaxESOtuylfqyDvhM+Dqp2gO3Em6CzOZJeRn6bYytVFfQ0
StauEMFB4m6lIdvVZXhss1sMx8uqEytdLuVlvUV0Szd68aPaOu9FL3gxh+vU92hA
OQ3oFqoPQZ+kKMDnH0aoZdIf7pUBKYhRQ9BSOc8NE6TXHDIxfz3k2qTiAuA/Hw6E
ZYdOBWozTdEsWiQXPzcqxaES5hd8THsvNcCGGWmPlJ5REYqimBgiDlyLfZLdpnU6
vuemEtkjskTdWcuJqGQamaBVyz383IX50Gjuc2Xq5UGG8lTP1Ur77DU7KO2+QfWA
aJtaiYmeCUX30Xk5fmtDvrBEIjV4xN1+B8w9MdBk1fihQW01UoZgbNP36mABjK7H
2vROlFo9DeUpNiRPKJ9xwrwa/9as6sK8EPc3MaiB47iGT6SyIN9hy+4W0zc6iYWd
rUtJLFPtcaKL8lQ5eH9zc0y3621Brwa61lAg7AhlykxrG7m9gUMoBNmRlM1jROwf
6ZCxKpgU+21FzmF4vUiD1wiatdmmU4i0zsrvrAxtTeoUXdUJm/Ll5GhfH8HXypkC
/llSWpoQ7r0qv3vpOxVLTNOl2pm+yc6sBC0GEwLkeals1i7ai4MeYSe/CqQYA2BH
1nswY4xH1RGzokDRd0VNrsYmACJygtTNHviP2yGRH5Fm/StL4bSUJ4d/DguDSdkO
7ucVt0JDeMLlnU9cB1hRnP6vpPkoCUPbCCencqNhmOFMdzUDywGSPbK0PPLUSe9Z
h6k3jVoHWbvd1yIurFAv6AFQol6REI/NY/T9QPbUWM0AsJea6DtF3+QYGbUPlD/S
LBPjaprA8aKvPKN6T3+fWbhFG+Vo5oXiEFjBrMfLrqfSpGRhIi/YivsZFQu3mYFc
akBTabM8JcY48zzOBKqFyfcvyHgL6mWZrJLVrB/Bhat0L+6GIacuBRwfAPzuHSwm
sypWUZoyvyMJtG38ATgDSchDUhIwUpeo0QYMN8QyHtgcRikQWwm8YHAB5bHJ1tgP
/uawbE7KC5s3ebCCq+b9ULgpK49LNhi3CpsnfS3KBs+YcXccIOvYuj9LA6KZeLoB
Kdyv+BHc8cCEd2WfHDUuGO8ShK3p9wETQe9wWdjHCb0skNQvnydahmaYa5KdYuO8
9s7oo60FcBYW22R6SrEOyK1iwhrmTuhmCgDTfoprTYiKdRtxNu2RUHSH/JG4LTeu
bqCYbAQrnoj+PD9oHbuVEtPvc9EmU/7j7KfHyXTlrUq2FV0yS+o1mK9zyviQZCP0
PJreM6G/AjEf3sob1k0/TYxbxndzMRq6S/dDXEns+VZchE7/Y5q2XujWsgtse9cg
WmGhWDqc9xbSsphg4F0D8QtApSyUOpV4YjsVAoW6AIP69zJviKjeo/aEIc5TX2Ug
uvTWpkCHyztk14uH6XvqwIZ3ZuA0T78phLGYCNGTeDBEofHxS5+pZGjPLS3VvX7y
5jZEAg/oQmTZezfMLYZNvWvH+niQgpczpFIXJMdIiVrqOZCXshhklO67wV4exnFU
Vo/9GtXBffM8VPts5Iw+cYcZ8B1WUpHv+Tr2eMdFRuIBUZdM44GN3DXc2FWn7pfo
7s26VUXE5s3PUs5L0CcSp/fPKr3t25dHcR8dzwuHqD8jV2fuJdKLPFjHX5Z2WbhJ
SI/CfWNv1/DhqO4IKEz7NMQCNI8ay/KPG+Avu8VtFMWpZfXSCm0DZZj2NXX08mRO
NQ9TDYZu7Ljm27CZecrpREobqabFIewnFuEEQVyHrTmO4X7WpFEk4kY9cRCgQLaM
iDIoDHKMHZpzwKUo7fxnKMfyvmaVEPx2fqQC2CRGaD+lHeNGp5TbO8hTndC5zvAo
+rG4YAzVZkB2thfB1gD3CNlsyPQyrdwmKTi1ITNPoGIoTOdr1xwqsQDd9Wh3cpFj
JVAxE80vbGWPzRAerEMALgnfNFcTt5KiZsL/LyrhC60l7KN1y6JtQb2yfCtQGt25
PyjcrtW4PoV+NziSbjxqQphwV+71Fld/V3GvnWajdfRc5glxBzmLnNjvVMLNQCzb
rOixezBZ4v+FBKd206ZxIISIesuOnltKJwRS7cBFIjhf0HuRXlXuDxHsOH6PWeCv
/3Pw3vCjrVdsGK7VUplI4W4tXVzowywS+f9Oiw5WR4aUj53V+aWRAZGLGoOJkQ9H
4FfoQ4g07Tn7nyGJAM5QX7hx/mHiv4mL/NeY7HXPvL9KOo0vPhjyW57qEGSrYgX1
wQUezY1/svqk6OhG32qabwv/vflQoyWsvDV2Ikx5+thALLP0H2fucxyJfrBUjG24
8ibxf+8FCbvQUrNivLTBCq04dvvom/3+YmfcV1ScwwwJlLM83Fb1he2VxN3EhWEP
2rYGJObbzzq2+/+eQg88jfLgCGTse7pXkL6bPGGDDdabJAxq8FrrcuqUJsqU1ts1
ojTWGa5UgEkV0gVSBOwmpaEftuXf1WHZjFJF47tUzT76jA93JoWL6+IBkbKV8pgm
qkiEE2yi9zj8PYbTMyVql+m5d1Tc2vDnJK5Ftgk/INnnydd2LYE8KDxVhnSa5elF
Xc05mU8/75WpRX0qyVmdq8aNZCQkvbBOu8jov8T6Ss7iJVEJCZkA5boQzVpAfrmm
oW0TovGM0kZfTXqbbzzDLP/v9O+Eo5q3gcmUuBVBf1hAXXOc+fApYrryGuhQR7kk
AtBUT9l/Ept3TkXZQqMbg1h/ZGfPgu6lJo0/7VREAdd3IwguYJBqhiimHXl/KMPb
yLuEGdRiOG3CtXnAYGiwMjdozODI5Itg2kF3DO379ckQ2xVe9jjdj2pHm+2Zc3n5
xJRztmsaPQW/vfCpoUO5fxdzxlG0SroAEInBER4Pbj5VKxynZ7i/UgAXHNSgxVa/
zi0BNfYozkPF3p37MTDPNNAGmK5irJf8+8V7AervxWzWurqPvfZFBIuSEi1tuDkq
rKN2QafruME+QAlRlbxWzGxvqIYdiLLund8JVzdSj5Gvp87orlCXU3wEEUiC9gI7
TT++hZjktpDSojb+SSHWGHXhwT24mqFQDbBNazDa/xY7xl1V03j/JRT7+VQCuhgP
HjxrN5QA/Vh/eAnCFg6XqkNqOjeF69mU5gexaRcnZZp8VDC+5TVWitVMNAzyCZvi
cM3AIy0URAEb4O0zf8n8J1PEc92k8qN8D4y7hwpy27ZBABKkWlUWubjLI9NFgkdV
9l2785scevcFKyig/0OW2Ed1w0udg0obstK05CWMXiPybZ5QanQw7kefElZe7Jzb
tSyp1mUdW07MiwTQcTiKNmWXD0eRtCs+ITmGwE9ArCLRFlXbFoDXp2Aek+lE7CtQ
0VmijTgj/qEOXJO+el+gGfpZcI5vN8K9CuXRQmn7LylnwkzfukRQ9c33jfDnA81S
b5eLY+ZJhTe3sRoerNR0xJ7o9eSIXNalnm949DC0R9ED2+jHm7LMHL6YZTSQ9W4P
pXPxp4+kJhtjR3Gn0iIF2cihpIZjb3AsVA6tZgM+zL1UoEIO4UlnGAf79ie0tnGA
hJQXWSjScItNOKNVZreMakt7xDngsYCB/Z41nsyay8aGMvxM91D8BSgMYSYkbvIO
Pcn0tnE8/5jOeDE+0CNeG9+sdWT93x3K+WFCs1TIOOELS3tFJTXZF+02fFBSNQU1
CccDvRexhG9ZfBZFnOjI1imCLSVMeQiWklyQXzNc7fInilnCc/1sghFQSGdJe/pG
HDdkE2EVuhTeubQXavXvGQbvmeG+MoZDZjXpMlbSyKc17PvbwfZ0jDtxhX4Uvg/H
fcElLOu4eJXx4Mle4tVJcD3K8LD4fp2//CnS12vtgvEh2P3Z/EWxzCM2iGtdotQ/
7D9Z6pm9Sk9Z+QLUKRSzO1J8BxyK5Dlr7A+AMuvYLczAcl5cJG44OZNfoGeIVq6x
ZUx661ZEttFKU1nQsqTonc50Fg+6EUJtnoGmDWi1ctwblGDP3nINDz7gHb+GH3+7
dX6E7KS3wgNA3gc+diVIHLuGiE4pppAIF109CCy3vlE8Y6t88Ol4DrFMg5WKOExG
7lgzRIG9RbteRjX9I7sQQ/uaftOTDN1NIs4Od4yynBEuRKDqV22gYU1PEpQO8+vt
0I9LaL9rNkGbsKODlBsnZTvmU7vVJ1wgsNg6b25dckqBYt31HI3vqOWlpW2s8BB6
y/Kd6qxbqCGIjBY75/MMFHa11SA0mfwpzQVf4CLmuGiW0RQrBQHNocIFDSrahzBs
3cyzRn1Pp41aZek0PAU7FWZb2wuLcJcCF7U4UQTKDmwG/ZnYy/8N+K226jq7iRKJ
odRVms2rSzIb5w/rpzIm2Jf8ZwZcrWnhVhXcFXE+29oOodiu4z/HAAQxHVrXGiAr
FBfZnlxKRMx+y5hTE6pMTETI2w49dQ75xv3PsiG2agrV0/q2MnomDoAqT3ZKSw20
UcCLnDTg0I7IEgMDjT98eqq3WfOtPFi9I2vPXRgpnexuhs4d1aIJkMLq+uIC6HM7
Ubuunp68BQtoQaQmJarXV7v7jaUavHkqPNbmHTtAMZtM4A+DhoATAlCriFxxUMy5
owMY4nSLSKQKr6V7fXpT2uTGAFIcGRpMWyItfqZ5DcIgOWHJAbX41o9o6fVWfdan
HUPzadqYystBuHpgjg6zCI5LDCphtVAlhUH5z8FJxA5BUd6oifweBp0Dgr7w7oZT
/RKpTM77GLekDm0EJ1/xqGwZUYRAj87KzQKsONHVf7/167XwkN0SNo9Clfv0ms0e
o0TZ9yHRT0lNsNlXcAW0dstTNB6596JgEA25wJX1RYkeubsEEZB54RvROAakJerJ
jHnP/8oR9rA38bcwsJBVCYBqwgNfQM757FSkP9ao2nE++NR8u7uvgYqDfstYaHZ8
cvV0WBqJ+MGGPSx1T50O/dBbLK+gENntECW07ADgugf1pQzRf8/5y0ZRaxeslEtl
0cmTLPIpajEKkFkGZJs+ibZlCJOHqD2nPcVqvVcHq/JA3tuKgDh0f2aPA3oLrBqy
Mb4UC5Z/6DtFPYypmJktZL5ZOgCgfwWyr6TyEgLHhDuavax6jyesASZHq/5kOCfb
1KxnNrN3eP2JilOUXcJrxMJBg4wpEpf1B9IViCuMdzm4BgxyBrES/mkUHuQQbvtp
dGgm8bfnBgVHbLYEj+XJjJhhiwU5kDIa4ufWPG3rGjDZG+AXP0kkZvoA+QirLWyk
RcIdSAD3ZeSjzljkv8bRYRFOI5jXCXIkQkpdMd5jGJZtaANz4Wubt8POx9gsKgxD
MSsEq7OmivbgnuBig5BTkG4hTbHRVnFX+rkICIYossA4OLOUBcmuZ2SIvAEjdGd8
o/MDRNn/YSRxLwFnV2zN5aRtHLkDr7YxThRkKSVQZwbhrfM/VCnl4Nk9ZJWUjJ63
G9xoDl3wjrjnAHuUwr5BA2OI/knvZjMunSSwUJN26dKFl/7OPxCFTQoBxMy4TZAp
4WIxfmfA77BH/rxOyc7IcMSpowKSP4X0ukwG8RL+3IBSWYFw/xqrLDI7CbVLm42b
8rn3B6Js6x6XIhfjNt5+UGDBDkIrO4n+1AM3zWGEUBaNHStcxQ7lzxF2uORZ5T8Q
fAsXHrK+luJqHHQNKCvQQVcTwVXzoj0qlTORVt/+A4aLTnjx1f1Y1yFpP2dyvGew
MMAK4JrRBTdWTR9VObcKmBJ4JG/df/l4Nw8tFozKodJ6RnF7JJdU+oZom4HTIDPs
bqzVqIwNQcdQN1+BqL1ioigFro9GWj8q5mOjbtK+2DqWOU/QkxCSw0bXmRGVpzGo
ZGdEWylwov85J+iTEHhFfH+gYfJTtBl//1pWkoAVBqf3Hqg1KIvKvOwyE3WUz/uG
oSbBUr3WN+LGoo5B5MSBjbR5XOL7JEwTtVp92NYBgN0hxISXUwreZlhFDs23+B3D
DR7U/jHR8d4PWLEb91OMFmVOBJF6588K+qn3E9gK1sChTF6GUA7KZmwUHSKFdMiG
2OLptTv9NC/QMX4JcwRNU8jOYr94rOTluPEuIIDJEqw0u10qiDAomubVqgIFm0Fx
I72Sx/2dy43j0hPsryIOoppx6ii6Eutq15b+0PcLSZWyjZaK9rRaweQQL7gZzt+v
CEC5NtvOFlznBhrfHZ/jEIWpu2OVwJszBWTJUTLx+4F8CB0AzhnWU4aHlhhG2vUh
hLxXlBW+3RdyYkT8YlObXzpgWaSMpuXyrbouAvV+Eb6BV8D1pxsBYiDkOgYrIt3L
F0DJ4aC4EkmUsDOaXAa7l4GvzEa/iiL+gLy60XTqgWBkCNMcRR3ejoSHvOhAgMtl
OYouP96QaaM63Gzimhr8daaX444NBl3YYi7sP1VVVJfc0Qc3pQBUYwO8Vb26S+3E
BcNGFz39hYe7iPRrxUxA58AQRBEarAajWuV5iSFJOv5D6XyZGdg0NUgbzplflv7d
BETpV2fx+ea721W8ZOmf4yTgRWxNY1lSCBvsP60ZIHfRCYX6G43jiJgQ3eclV2wf
8v+FZRQhxeJsy0XOaI56jNQDHNAR5mjnsclZDpbfLBYEgnDfj9UHk91Mp1Lc88BQ
aGeqySankgHlojDCuGOrrQCjT80ik8yBj7QW8MIvpYiwAj0McEPLd3ITKLdP4fvK
qxK88Rf7u9051LDx94QeNGWSx4vfp9fYJsra6ohUdkyTArISExl+MYUz11jJpFNR
rGjmWxt8RwGqQkKEaic6dQOSQThgll15Zu/unco+liKRyggm5W9J1J8XXZSykuP6
H4u8WZ1HFcNy3TsFxcTcs4eVpuryoBgbUIY9BxnxmLF1hAu50HI8umPmSJGk+sSV
+3RZVji6nSCaxn2zeUZBlUARSM2xO77QtynQugTva9xpS0RreFZ6uNH8SSkS1y5P
Gi/eeb5FY3TXe+mnJkThe+azQs/ybJYHc+hLqMd+6yhNtVKB+v7YEL+Ve2Ts8ljH
9ElYJm8Y52thm0Al3TFn8TuhBXBQnx75L2KPjpIJP9vz3koz75oj9xaUgBZKRFOk
kweHoYy2JXdCG2onR4CrnJ4z5ypS07Cl/xQaWvvymsirzqaId9aLXwuwWJ9oRwUg
gopAEm0/FkYmci7iio80ovu1XHOtlcHzYSR12Rv6ZS8G5EcfK3NQJRrs//yuzoZC
DE3esxEAlwSwemstt9dTtEWZnPqN02s6Umt+sxkTLF70iFqxeeimEAt4J5zNjenf
J1LX7tJiQTBJ7WtV/qatc5c96BDbo7NIpQBKEhnmqlI3rXagseQViec7YZYwEW6z
PRsNQ3oiMDJP9qqXwiZWsnO7F4DnBl5Y/MY0un71GfhE0Zyugtv5Wzt1LVscZjQM
V5CWoMuqgDDy2qbFxhdvBmrZ+vJhZ/fPyELHFmMZ1ximbUT42PPgSCMiZe0oMTNp
FJjfZM8QmoASkMbWkZhwBj1p59THO6qjf2y/orbfDKMXsXDuF3hx6oHi0kxeNEPN
6wGJL/OkaCHaN5u6DvgZwkPktIK/KVt7pJUHkQBixw6Bz5atvXSuzHz0D9U1II4g
I8RBFwfksOZlCitqz4l26quWdj1UEDAohdfWzBa1ejQN05+OcydmDSifJ5BYfO7j
7pNnye3OotOOnMVz5jrMP8hdaqClNK45r8FQeHpM0Yd3xQ2aIrhTOlQYGm2Em4Zd
ZfFrSY/OUk948Z3iFNvGcYj/lY0+u/H2rCYBTXl5t5V9sTqUnjhAgMS4+tyf/LEk
12u3pVy7pwoLDlgluG3bkY6NfODyNuz4ID8Hq4Pb/1nYTjmdOmcaGhXEZvNLdgsW
/c1aIpRU9gGhkBOR0S227m6E4wyC41Q1gLowHn9Uwqo0HvLDPPAIMBQCnOVmvmBC
fQxD6fVnxDXxz/8O7yw53rFlRv0MUMNeHsfDf8DWd7Cxzlb3vSj748iPJWiqBP4d
74+ZRudg5OkTFvdPmFdhoI62P6H2n3oebVEBaDYaSR9MOEwZk/bwTrnQ8a7Dz9Fw
T8jatdqRJTaTN2/YuvlpXcGdmydduwsEigCJdNRLTbOZSYCxjdTWBxr3rL0X0eWb
6tvMCpx6Qy3kzXYPbud2ollqz9l01LdExD1/s4KfGz5renHunftmejqptKQaWPMy
9hbUVhM7J52sxQps9NLKKtcXTP30q8Jh1qJc+xhAmZKuPcZULjSmZUwloQbfxTFW
8pl7pmIWE1417MYARq+PCdZbmP4b0NQgX1IAXjOOaXrNDSt0v7gfiYSbDkJ7ds5v
jSSCbsH5HwnecmkWzeFnp0NTRB2pDqa+6Bp/2HQNrDoYBzQ8a8iaLNHvZCvLBlTg
HYCFv5NnMX7gahq/RwruHb4s73h81XqMMJofyGQJrDW1RXXoh4ErRG7eoxqW83fI
ryo2s+e17tSDfSg2ij/UlLDhv/M0eej+r+saMdJl4e+Ok2t7Os7RANX6aB+KfSpM
/Mdhf6HONZN35JhtN5XohWPMtD9GkdQQH+oBlwdEGGBAJIlStQdPevU8KaRoR3gF
UpfZCehqJ37QH0xEpqik+u13hc/q56jozyaT7x6P1AlFiFLZCSo8EaK79ghRXHje
BhcdTp2DsvbdCkkmavGLYNE66N39yux60C4Q+zHCE+2xZ7UZtNZdDrp/ZC3rV4pL
OxyruD4ueY21HHR6kF9c9KKp/bqtFZKYjsXPYBIBhve7wnKb9pcByd2MTJ29pnLl
x6nPHdRmTPxgCpsiglyg7hR9yrrkiuTlr2Eui8/cKg2iwthSlQ2yQKohBIl6MgcV
GiC24IadEx8qVjdwWblUXKBb2Q7F5TWjsa3yfn5aToSNJeZMq11NmhshGilpHFLR
xyWGTkAqFmkW/b4PwoRd7AUJQr5Y/GOLP3cw+0okKg0cEriPJRgzyOx7p//6PC2n
o7oAdrn0lCjeQdq7S57U8EY0FojRlBwZPGAnISqKdcwgMaRVGVC6vhRc3ktdysCx
rHrbSsxSR0LRLi6DSZRRpHKDGjqAg3mfdU0F+GSw9IseEbbCOQLgJGOVz/nReMCI
nDsgg+ENzdmfYHQ+kv6rTX0BTH088AQfwYbbCz80YWDAxMgIsSIr1y6kDyW/oeo6
3ARkd4OeklzkXuDw/683eGim4uJLxDEMNF3S2oxsbhe+ISGYiM+Kba7pZkxpizyx
NJ1lVJoQyrmn3SPBmP9YrB7DmL5fhb9gfjK9RRqSET2TQaIgAGU/vW5JEUL56GB0
vkvOkQZ42r2XWsSgsJpO13mNW1nol6WabECAs4WKg6bwaNebSgdz24IF0Ds6TGQk
J+VTNSN6cI1T8lpduP9yzM2FnhVdi028NTVTGHPZCQkj8jKKe9HqTLW2YqBw3ZGt
XGiSOUKqgn7ozTkZ46Hae6VaC8PYsg+XSX+1GWKnxN35R+kA0N/ccu0ibqGzNzKR
xFY3y+bkafELx0NFQFgmcF3eTOo2MVECzS1iAqEn2HK4DF4Hj7YgTVd0IKxPc4uc
0kSR+chcN6Z+eeBSZWEHUyepybBWGrQ1afrdJg1qZF6MTk7v7cSjeqmpUZtV4g4h
IKg/Ba0/R1sZmjpSUo+fKWFczrKSL5q4bKbIXSshflx/rXJMPG4Ky5++bFP1ufTa
cnB+RZDot2V0FPQ79s4N68dW2NYroqd74zRRuNiUrPqRd7lTOfQfnwDc38alOZAO
xubhzrm4FLKplawsysOu1WYr0u5MF1wIWCr0aBDGYSVB3ULePu/53U+iSjS2GqeA
DX/3vqnlcDgDgMJiYZdjKa2vIwZlf3gtj+KcN5NOrqiX4tKnXeSuXal6i3gURnhD
9VrrijP/WhfMkpz6Xol0RN30vKoIAwyDncUQsvA92yRiY9mdMMyGr0SB5L9Go/1L
f7kBY4HJPqiwx4MhQYCEffqMFYec4tW8fvFmudLOblZPHPcVe4z+R9dCFDjCzMYP
nThrnr1XiRstP7VXch9iCy0xsiF7RSCTXxVcGw1Kg8v7DRJW0L8CtUD7WLVCnWSh
Gk+4MkNLI0QXbNvzb2ncfXK7PL75S7NSKgv7BRz/G5rcJ8nQSHy1m4EIrrU+HgE/
kVLAsQtRYkcEmk6wA7gzZ2SdWjO1AkhGYKjVKlXeBtAOepa1yAfFp4AfKDDbAfKd
7+D3DnABHsj96ApCuxUqKg2vailgShv/OsTDhgUhUqWV+z18YdHVFktcJ5pJLJQ2
vj+fPJu6XY06o0D4yTDGmZedPkPVt9IC0MiCPT2SOljxvktCeLOiblGTqio1eat9
mAVugqIs5BzMq9NPv1KXrQUCNZdb/jDfsF8FnLouq7oxntygH20GaUkHYrQ179HY
Z2EqrXLk+JwpjeQo48K1lw/6w+0I12DKa2dAgWiaHieJl3PeYU/p7dm7aIR4+bgj
N8PDyAybFDQ0VfZSZykztzzU5DfjSSK0AlBc9n0k4c5r1P1LeEneaGwFnr7kUepg
41BG1MpiV1AKRrJzTktWB4qPaaEQ1T4KreJWZljzF+FtfupZZW+diR6gi8jRompQ
C4CXc08/uTP9K7462biMsh64Nwqo0pDnIwsoiSqgS65qAgUMS4kPCUjcub+jMhvt
Dpag6zjerBQJEaTCsT3kS1X7Re87MC7trRQplPVXZaISJa8Mxz/A+11FBnEuXN3D
907j7mYCa+lQjnwbNxOcpp6tz1iiPlF1toDKJj8xfbYrLtcu2sOz1gy1mM+i7b82
SYLZiTpyCsMan2NYwZvxeROv4IEpwa/UV0LW+uQDBhOtfnPXP5h4A3EFrNxtahcs
gWLfC9S9MFU/dSSjP2CIRXhCG7QXBMHucEjod9CjL9gCHoD3ytu7TzwLq/X1hSzw
YvZwkB95JJjUpnopCmCWpzEhAAH8h0c5c7eCAmsccdQ5SwH3Uir3hbE8tzpJqBWP
/cSvpxcnB68MleM60a91rrGAPGmBYhLHee5EhKTX6rQHRCLzPv8zAEFnYuIteN01
3et5p1at/s75Ijb6zbmX0AeHKzHUDzKifh7a094cH5AbYRHD6jQT96BhyRw0Lov0
EkTdJLvrovyJ+1ox2O9u/V7Vqv9Ew42gY9g3ucSuUDF309wmDEG0UcZ3TYfFJhtw
gedelGDn/E3lu+b6oYCaM2WQXIW8gzmapwp+eMyOSs03zHI2Ih3CUOmYJpYckrGW
6zC4Gm8auW3fqL18U3WhxxAofXJeUuaKM0PpEoi/Hxy0w8ItfqZ3jxwFXllaxJ1w
zFpPxAtwa9bHvrqVI8Wyrm89qyUyxUKeFAD775BpOwaA6Uq874fQ2kxLX+1Y2nhG
vVQnHYaPnVPyMwJ9AV38UNq6wmas2EO+q2k/LsVA5sEQCvDwUusOpc3Ylb+ydGBm
rh0IDQSAX/pyt84Vufik8UhOSHtoJ8isz1H0lFU9Dzuc9vx40rImCs3jYoUxYFaP
OrJSvj8g0/3H0C8h6QqD75MPNLrXpAUeJBRyWHmUTGKJeS9PJhJTnkzn8WlW04N9
gMWmdPh7XRisenmJrOE1zjEDyfmhsYJAFvA+xawg+WL96ObVMAUo0ERaW/Av3Io1
9XQtnytJcDvVI8wZ6DxaJUkX2TyHayNztcFUF+V6UYOIGu/HiRMJJwHCpI1w+yr8
Y4Vyfw3D6NMPXJp1jKZ+2/xJQYMl9t/Pf82IyBXwsVy8Muh5klwjHeOzJ+lpeo6w
2t4iwRMUar/Js26dslRoQNdfa8YPo5eufvc/DqmtSG63hhO+/5muebR5Wc+DZRO2
wOPeHbtL/JxqUIQvnwJNKOBONwRI6Zp9ur4bVdEDI7ooajKJS0b6L3fUySjVw3S+
w/thgQ5XCn7hmQvCti0pApshxp/iLqkWyqDrg0LCnN5OldeZcSG43PQMEQIql1/9
nmzZSfmqt+dvqVHeJvAr5ANI8IBjt6izCCYR9xg2QgabnqDhViYwSOuQYxJaPfeT
UbmM+GKcxj3nnoCeHljsdbjyjH8RLQ6OvSf5HoSzpTvTLbZdE2sxaKoUwwhK22Qe
mhogJXOZNvTcF4braOHPprefB6y67B8A5R2vYshEOZpQsa+mF0ca0EaLEGHWfUIY
gl0Ok1KlmTa+vqZatwsL7PLiTzFMIwk6wdO+uRi1Nxu1pVFoOVcKxU6VOGip8e2T
gSRfsW1pboHuMKkwP8BVEc3V8y6Kgs6DaVjAFEgzPknWQTEdGIKfpO8H4BRM72z6
R5zhvhPAVzhudIWGkxzQj6f/8yEtJdClFMmAKBNk53ZTtYKWyROHgUBSpimlTZgg
Z01JA7tjcweGHguCI6JErtD5HioUoe2JpsQ8BX7W+cgegXs7FgLQFEHZPJ94K92i
8q3EWG9J9k83NUgO97E/wfBrVRvltakEGX1SZ63gm24QUjCkJ/2cPGtb3GEgL0+p
BWbOFYpeyL5FAqzYGpQ0Bif4p3abmLrZKSVlPMFjL6HyqmKt7bYGNEgHf+3W+/9S
UUV7MzV8cI4Rmscmv8Yy3xVuBJlMPsvTbBSYToobwMBi+yQR5Y4Ow1QUy+WvZBBN
4O2dpoASPQIEVo+Ks9kpIHZQbL0fjCUekGF5deP6SaYxZv/mGDU6gPL7AaR3//bK
un0+dZeovXk4JnxCe32znm3ml8eNKa5w3MJ37Krs0iK7PmBPUrPUHjWVNNU21poo
T9M3muzvRpUlNcQMb98B9+DgPUkjVIiEE4n7JwJMib1NofCl5vdS7rUjpZSfE4qm
B2m+Hkk/idxq80R4yX9O+0buDf8Jk5EyUadYd6KtDrjjyWGtjFKVnVmj5eKmFppH
2AdXe2rdSUPwPl++fLRQ3N+iEv06lTH4BFQl+nRZuwuPu8g0dP+KNFl24tEb/UZ3
WlrzeQ4rPL/ckBYuyUGfRtB2yEaZhk1kAQdHz9vEuKmb7/yz+TzefK+E45Zx43dk
IKft9gBvnFubqtOvQF76KWPtfDa7S7/hDfBq/6Hef2LqKnPMFmtIYIYwvgJr99uV
D0yg/u/Fbqqnuq8jPNuDhuNwYHRQMRSZIywIImDh7+25ts2qkEq2/GhxpaYmahNr
uhrjMsI/QSqpXXsjxm9h1g9Ue0kWzzvWZX+olmBYQOX4ayBAlUINJhYf8aihT12X
aNOaxRNmLG/o0RGT7bfG2NHGXg1kMPmtCaq9YNMdSeBrlD8wCI8kQlHsntfPnW+m
1CXiwcA9HweBRBKaFJyDcOD9iz1j0PXMscwcBeZKKMWUJ0lP4pVdbTq5WSV4rEn3
kgua14+Yli5Msy+GdSIIBfCL14pPhMkVMkX0yFYIbvF5mZ9LqgPnS5t/YyXtaAiQ
fHqTLSi5cRX3uSeZfYEKy6ZZ1FzWQg+Bf0cloquPrMuyIOMhEOENjNHtz3RX7bY9
weGi4zzjLu24QE7UHEaU+lliRy4mNbRT+GVFkB542hp/qergvQLIsLiPsgKgMac8
RpeRTSHWLbngSoaFUjGXgbHTJEXW2ndR1vLt02aH/RMmWV+kwfj6ZHCa3tr/EQjb
sENrLGaji/K5A89/RclJu4xhrL326Y5sK/am1YZg4gXvWN3vuWwcAC2YPPgcRhEr
5+VKiywdUSz/u0dzExw3c1geqULlV4QEbL0/W4qaRviya6WxNCPZ8s5SjzNsG79T
Wizfqk9Gz8Z2dhF9dQw8Z65iSYRRhMS3a4Gg3ppmX0FWpGP3XPweX1IZWiMmf62i
jAF7kZ3GNki22ReCkcE7eM0uUTet0WWOMA2pjhPkLelb/FRNk+JnV2k1HFSLR8/w
YvUzLtlV0YTeRPiuQAP6xF5tOB26h4+SdbYyFKSSlMHbVMlUiB6IZOHm7L+oWAsO
aoZRyaCIX5kua5xhDQDVq31VLn1nL+Lz5P7M/kAIv87ZfZMsLjwuPCbg2vdkFMa+
fNTBVRBEjzMdeO5tVpgFhPRM3J+VqsdFYjXg8nvcmp/4EaPTg3rnyAjrGGYudeT8
4VCW32/gPX/TjS79B5nQ3rnJSxKWGe63qXOybSQKZwgnbktAOrGWrEN1j10mZNFq
B8F8IV6NKqMTiUHdSm+XRFjjYqSx8ed5E5/4e6wRyxzXCLnGWxSMVCwySgmclzSd
5VbiIUjjiGQKmBGyB8Gzt0mMBx8kFsgEiycb+EqPpJ+9Yi7HZOMjYqESxbBEhtLc
CRMSVtxeupdMHVZNxvD2Ihbagxevq3J+NOxjGAJezMX+bQb3YiQAs/3OmRq8FVTX
+wjiTGO73t/GHQO6+CHwlnJFXvgdIDG2V9KhowHJtNCqA32qHm4ifVenwBMnJG/K
ttdUhcNQaugVZJibkBWkbPpPlQDmJlG+2+s14aC+4Pmz1JxqRvOnW4UrJVZ9Pwb+
tGRtXTQVQQb0i+Yg0M3LhzbAG6NOnIYkWebzzg630CP0TapdiBJWSMpxfQAaAB9S
/2pjyLj86ld/jBQYnx6GZVV0QIzi1ViN63CAHMXrSCK3YnbDyqxUzflWCLG3HER6
9+iG7D3uxZz6lphZug163jtoqqHAGEmrNlthXsQan+daS1ixB7e/ic5iBPnelgRC
PjvHOpouEvw9kgLlBIN/hN+htXPZUTisq/nanzu272uaLY0wHnxuC1G8AdkHPvNR
RvT8YS0Q5X/E0wdP1EautjXK+7SKIGQj+PxX+r0QOQb3Sv1HRlIZSQ4tRaDOoLMi
poJEAZa0Y7TerAjMVw5AW4fGPWLSyMmV6SqvW7LP5wO16j2EKreMCLarq7gAVyN+
h2290F2JWjDg215aTD4Zk068/w+d1XmAAnZhNFhWPzvPrDMTNFqA2P7LBHnE/vfZ
P13/YUf9fGJjAp6OKtRMsncb+ZzCaNa3a2AJUgQE/710YnjjeoA45f2/jBgvjBgz
oG9dS06LkPCDLIdTst8mr4L9LW6Y3dTQa3mnVptmFvs0Jof4cn+55yjjeb+BCd+3
w808IA2DxjEtEzEv30MLb60N5l3vKadmd6lJL1/C2rCSHqNsaadqaRWKYIlEmkWq
qrREPfJMKkO37VTHWKPWYBDEVcTw8vxyR40nvRj+FW5CYlFTxITZt3myJ4/33cK1
rEIBrOeVW43tCxr6VDqy27t7GQV9/j+7sdFbOxPyCYL81iVR2eoclt89ylAeiFIH
7ZXVZsiy3GV34Mea/QcswtuxZE+We+zNAeeyviMeN8jhXOecgnu6mOiYrkokX5dt
U3MtMsvmyCWRBu7jyeI+tLlP9Il1XAKkW9gVk4qfIG9NM44lL9GcAMJkN3o3NBuS
sM2RnBlVOlwPpVPlBhy7DfllBfOzU9tWMhF9lJFWVcAECGZfkix+/fYkVZcOrKhd
Yp5Tkvy1WuUp4hSmgR3vSbOtVHoUdkZq4Pf2xVcIr0xTFomW3zb9VR++ZcWddr7d
AuFGpdvKHo8Fr4awxvosAHrOTFSb7WzXCRYdAr/NRuKDaZ2+mXqWFFyT64xa4aJu
3bEPPxpVTHehoLroH1JdlxjkMvDb6H9+u9ImqjsnZdPdwOznat1Q9RRfUvSeTTu2
W0uzxPQvrN6iAoxFhmr7bhHW//rszm+so/tX18WGPtquQgeNwBv7vzHG5GFn/qxn
BMgD73HvtQAxJcHsDHkK9Ki3MjIrHL7vIhSyJBD1dc+kawepmcrciT71KTnktLN+
hQttpjr28jyoXmS88hBKhfsmA7as9UBl21s0GkKKTVPj7IOrcJyRlC21/JltQH3r
pgHVZaFBp3HeKUQ/Y8bJX4KDkInHO1+sl4wMZ0W9xeLS3g0zevkB9HEr9/tsEbtZ
3jvwFFuDQOHt2PozQNvb7WN15T+yjCc56N9mwCaMC04gZR3WKCBB5wGfrzmHBnXJ
Gq4k3jiJKI5EsFplgurkbJBMF/bPywl2UWlbD4qJ/8cx1OM8re0K0z3sh4az+19C
YtBigmDmSXPt1neSQVqKSMJikMy23QHf4KCerM2CGEIkUVPBkIpq7Vt/DP2gzpLJ
YMI0ArWWPHpVzahovdr/4u4O0XwmGJjAdrsZrazY1GkmbXlmZZ+9U2LtGK4/6MCc
DWUCUtmNyMgaCVq4UdKajDqBdE8AuKIHO2BhI5qymHTaZ4Q284eB+MTW5+oRXXeW
zLOb6D5LzLMPu/zsRCiEg0tW03WEWJ/W/V0NaPFv5J1ghkDBwROVHFze1uZZNy5L
t50foWPuLqUzxD+OgC3csoWKvY23KoW2xUUKQhS4e/1tw5cTWpzspj33NZlVYbEF
PFkqWdQHzKOzUquB6q2YMDI2LyWQY29vLxWcNJOj1tTLtGaDtpvCGzt9O8UW4h1J
A2a6wo3NSuzoBTGaNnhRSrfDUtOYxmts9wUXVOyjFVf4mLkev5aVHiRVlJchY9Na
6eb3RbTQKaM3W4805k4Hj5+8f1I0DJxD5jsufhoeDr6QqPOvy5zq51pzyaiJDKev
BPSCzW0pNiuO6mibMvGueXKbFNJhLUcamXq59XXzF2AZwRa6pU7MRrGu6wdFalX1
uz4xAASV8lh6yuHiyQET9IT1wW2DcZYJk1zIgnVhSUgLrLo4Dhm4MhMnvfAjfrB0
YQlCVmtYhAqk1h6FsH1rx+PeFWQsfIY+hSMh6EoRFfB0b0AQy7qpnBMbj9mk7qck
tr3ptZsMAFy3YOvaPfdnIGlLP22EuCsrgGDnJGNwJPhmNWdu3X7RsMA4nbkIrMc5
7HeML8SF1+S8XR7ION8Uxec5Fh5r/kAdqhYsJdAGRVZNyjyQCMQC31SP3XzYRIRF
AVBorttR9S10E6q7tLiuhU/0Ijtrs9C2fMKPn4SXAooHbMizzm60eppvgrswTjXS
xKuHocOO2PtGb8xTqgSWgVqvIlLIShIeyVf20aSUUSsyjmL2pLw2u00QqdxsYWdd
cN49Q9SrC4cLZxPLZy8dMdSQybQUiA2ptd0NyJlZxgmeY5L4GH3W9pE6rKcYOtmQ
UA4GTHxoqzD8jjBPD+ehq5A2XT7Rw5tDzrP8AaJRGggCoWT9zcJqkuhJ1VfeJnPe
HYY8vqJlN8xP1ho9Tva2eeJ82vE5o31yv23caM35RcEVBewA8/ymBfPHLMR0QSdD
niijSTtEsvNXN0ooL85/lCHras9WqnSMxR9WZ1S6rFyRGUlT7Mbp/fOVt9A3f2TS
U6RLmZzN5hPMMXs8Hb1T5q2CS183qmZG1GOD8CPI4VqXDbnNS+yV98moVg2G/SZa
niGzReJrJ6sxi42or0hX88FFZwmYx9y+73PdXHoPP3r2WlW7JenZOmj0DY61kNxf
kTOVjiSmtlUR/V9aiebe4FkD4yn3FEOZ3PwnLNLlBxA2hioxqivLzQHboY6docDV
v5ofYoJ0qYLdTP786reMj94D5IPxYJWRWnStfcpijOD+KYWqL3fv9txJJ/GnGiXB
xFB+EsRfjWuwJ24eg6HsvmgQm06WXA4anzVl1jxlywuncdnZGC+MIT6Dv77wm+p6
5eUSm53A7HleSaI1T2BgeLAqE+Hwir9cB49GPyH6NIQdqYOGml3bOVsqm8A+GGra
Htduqmv5OQpUvAWruVM0ef3h6b8QPBdiIbgkniNTSY235uGIB4Qurw/VrEXBhb+u
f1RMiTDtLG+4uVKdaHOy/rHqHuOPb1uC3B8CNbeCfKYSaRjTdOA/S3dpvQBXqz23
icBPbDa8Rp6Pbjs5dgW0CIdA8aIxiKog0V5qv4Ze0PQFPhiZ00uK89gPvxhZBn0y
i99NhzNE19Ir9/TPAZ+kH8RMPxliwQPQTLFT4q7KN1wflK8pt2PBfUM+3g1ZkwHO
ugl/RupG/OQie8VH80b5rLUY2lgAeJfQMHDwGu/V2IX6UwcENTyxqduWai+T/L/z
tu7HcggADr+17rDYwMobRS1/z8A8gx2ceM63Lla0x5hoCvAodh+xGMHRlQZbGBRY
+xs6z9q1yZN7z0gQiNuyR/Op9DQKOphaUPuYlCAWXo2OmntAaNaKR5RrdJ0SQNWn
DnZYHk918OINU8zwEL0n0BrAMoaGdaoPMOGQ57/byYsyKpar1MwFAAwy+3nHTDa5
alv9c0L2lvlLIJNz3a04Ok8EBfHOoL5o+xiYfzPyyQ19hbsJwi0UzceKvZnPmkvM
3mN+f0rr5fPeQSpgfz4LW1oxQebeqgqnRbtWmt0iKxYxCQiaWM/nOvDE/2TMRnQO
yr+Jll/Kkrv6Yd+05cqnWLw9vgm2sHRn2PBd3KClm5eRRlFhPkZmzEp6vpRxD6Rf
zOLvVhuP2vCG1DW3z0XSrFXjaD/hQSRLMIT26/8B5mlpny+JGjFjn9wftaN2H+Jz
Sd6guon6IIBJOqeL1N3hbBQP5bsxl6WyXEMUvtYtkmOpCJg27gBd4NYz6eJvkh1N
+tkQGxI1TTJLVtornydhnhzNwbNTEYxYNMZ9xRBUj1ZixWPumSbT8xQ67iviosHI
0fb2rARtxXLhAaj2ngDRt7nHQM6L4xBqQWQwM2oPcRpaNQ0Ft8o2vRAe4zEfUBtx
rTuIvq/VHBWDZ5miMr42qx4UP31vV9KRhBdg9Kqb/J7/Nf4QetRI4zbZkSWfrVPj
zpEwnnyCdYMxBbXFvMd9ezsVGXK0YJFCESuFKedmqbF3D1etUMujZFdLHsGsTXdD
GF51uvLLG/GBohds8ofEbH2EImSzkEJaA3MQMqkys2GKvYg4xb0wbCk4cGUccup0
No+NHMJUtU2Avl4BQpa9I5kd2k16fbgwpgSgkvHoKNVjc9ROVibaBRGmUgd9jiTj
6WV39OJl5vcfkSRFGG5TsT50tI/Z+svfMV82YVnEYeMCk/EIgBam0sbPe184OtLW
47h+W7bINTp2eUfOb6NoVFW74TGv8yCAemMDnc5T+r1nUNns2L6xUujO7blirrK1
xQBHVxTiXwMq3E+ZjDBg113l62C5oqLfOLX4muX/G38tv5hXYqZNycld+vj6KCJu
SkYeHc8Xv84cbHBs1qXQwKWxt3FQJkfsJ537RjnOlMwCh/tbJDzAq94gbiE2rXHr
uBmxiDPgh1KPo08Ub1OnLM5iNDJY4mcjvNVRtI3Y74LGZGT1Sb2LJXatY4q+CwfI
rtqlJXKHLSTZp9z//KZUOf2ZCCAs7F4ydxLSVB9qyA8k5efzCKIlRO++1XMtseze
5/1W0Le+IgTjk9Q+i19VRAjDIB0t6yVLIPzy8Jj62ZNzm+8DABZ1WmRzB3HRsEk3
6CApg4Lx4cb9HI4F/IAdtaqvDvTOTlYySQeUc4W7Y7KtorYUld8b0QbuFj9aaY/g
x8mhM86ek78B7NdKq4kYkA2fB8NbZx9LDeQwaKzwWrgtDdN8RCMRftKbt3BROKQV
pZUQajyxXE2WEw4u3A52JGGiGIx1uOGbdLPZahrPWx0stEmcedk5caViGy7WlOEc
EbcAtC9opJm2rHtHq/P+8ysIhffr8UK9f5B80bcEwb+oL3JjeyO/VJ0IEUDFwONh
xetG0TCrnxowRo2asL0l2nlQiuP5sjJCb/JfiTifyGKxu+XuxkLwCGLyuTn0opoZ
vx0VjbN9layuCqoO13vCXYP5IEFCOF/6/fCEPEU6c3LhcEEKNCt+eb5esAAaUlfP
eCk1axcPORwGpv12CpCLbsJHgCGWaKO7w4xkIjIhLk+JAny/hbaxHI0tMBiy1/Ss
HIQRF7mPI9doqIPmkDaN0MYDNsJTuSS/cKUsIZrcPKGip+dgI6+EJy2xuhNp78HE
vjQ/lDXY0vT83c888Nd1WsOTepr5G9x1TTwrZJcnlK0um6Qw+1w9/D1+4kHmG4pJ
yzUZqwjY9d1eqADm5mltSBv5IA7zmvLXYOEsnnlERa7J3nz1qmzPnXzA849eSv/u
FtTEiRLquBOkEvR/BseEsPRFjCioZeyTQc7qSDVLAmh+wwYX0drfzE6qCCmgGo5V
i9raThhuHADtmaWLXqrO4tyq+vDkM/rD5OxMGdPQbbqxnJRLUQy5JUOtBEMrD5nU
OHE9U4QCTwW61n4dFM5UROb2cgH67zeTS9zsTHEt9jundIjB8WXcae79T5R0dHbd
83xl4yf+BvXrOKj3kV4wSGc/XFHv0UdFsMnlIVsV+xIFiUekZLLj04y08FwI0V1M
+LTWUliY05j0Ndkzf1vwf0QZY827UPgcdedvinbZ0n9bCNUi9kqZr8o12itM0C+b
SM1Gtt5T+wev33/iqb0NjByxn+S0qLsiJ2J3J1iRaN0XUS+IpPgUwzgAbEs90W1K
OKI+xVLRh+s8mp+tUJdYUzkfCB2oryw8XCpDwKKjS1omYeU7jdNrvo7rsfwn1wZf
O9DA5hbIPTcMPeOS4UnbCsnVaFWZx6lPWjn5yVG2sjhOeucBKI4ssvt8Rn1ypZed
MIH+MDe1xdFb9qL76KRfrl7nNDYMYEd3NY+1+5TDedR54bGR3EVY+r6hyBPvmGwc
q3lW49AMye5Mod7VjD6fog8Hy57kI4shFyncu5uad5BWRkTp/GHY1xKc3gbNtmgZ
VLYvKmYgcMs6cMtW6rleumDQimQOcZPm+yO+aj9Umfw0AoumxPGAa9YqjDLKnSq9
OQ2GOzMUG2f7MxZcm+rgIdDOMlz6i9tOstK1WvFd/8wg8iiV9MhPRK/HY/KhDv1V
LXS7M1o8jU+Vnv3goLP8wKym7aKOzrgJU9VlJid5f5NtImu12L6un/y8o2wSV6YE
gRp0Gj0zwlySuJ4Xy00YTUx/CkMme2YZRYgWgZojTLqnP0R+bDoESTRC9mhzwUdP
ki/WJAqKb7U1fsC8OqFoHNjFbA6zbKAzZK9SUZMR61wUzIpz6+/mHZ8K3g1jOhBt
iONl1scn3BB11lNHIBK9+14dMvpn8P+CVrq3TgxvuTajGIOcaUBEqIQtk551K5pG
7Vi5MbqZIiOmSGeAB354CIAOgFj4hBW5c6Nc7Fo11wrX3Y0Al1oqooBaVC2jjr60
qP86VtsncT2kw9fojPhcQWUvg5da8veSfMoZRkg34em/5D2DGhpBtZNUkcgpjwQL
KVTaarJxh2ZQwZ156hK+Zvw0N7Z9nKmok3lLSkrUqBDa7zFsZzbx/XsaI5RcdeTY
ombyQOQw+u43u0UB3bs8nBKe2DomVR4kHQN9dEC8njrSLcMAgM2FcdOqvpIlX/S3
J+orFM6AX8dmJeacJboG0nRRFaImYodI1u5AltzzFvRa5dFKQttNpeLO3nhTcoYT
h3OmLT1pawDrZVaxqVRhmIfCkYYn/S710GcLVjTgOC/AKW7FbBzt93ezK3qp/tEk
/eh4kLEAdnlqWjpGsQslrcIornoh5F003jqRSiGBqESytPMpeX+RV9XruzhoZdDP
4NYfrDHlA0gfd6mIBH8tLSIqQ3cd0leZhReH6p6ttE2XzcZjCF0XmH4UyU/f9q66
iXbmUsN9PaOoTpuytBcn9dS2V4DAM818iytRqgRaC6Rh422msWH8IQWAlcK8N2SX
FcbvgCHwjezo4VujXEuyJ2Q+BHT/Ifhp9U/9HC6bGbcexKVLWtcSNsn7OWJvjs80
wXg7dDuP2HsbIiR7ru6eQMuNcvBFusUx8tRfch5xjlrVfeIpGdZu5g6P4zd4kDeF
1JLFnJotkpKE5+mZ69u5s0+tLWABzPpc55Kjevr+liVKL6V2BK1iq634Tt19Vymr
P7vvbSeyjpXnPtMYOYronhqmH+ifHr4fPjhf7INR84mxLm+WYkOHdOo3bwogvdaK
KZyH5+aUYIhc3SwFApyxKfjxQttJYf6kIoaA2UJB9r7LA6uNRdNpNf/KGlFKpnyK
EwLyZYy0wtA+ol6hjmraQWvBpgz1AukH2Ttm3u2IZFcIh0vGJd4E43b07gNUFMf5
U3ZXxVTYoDABh6lDFFdaWC6vmn/Ts8AsA0+tnlNqvY7tOOeQvExSBh63XXX6soqL
HRpR3Uy4F1SMgHuA/KXskW8sLtU+BSAuN/IghQ6lCoFwvD6VCtPwX+9dsCyzRmQb
qqUtKooKkOTOASLheCV47JM3uhEype1UzoNcCmN6wocoIKgEGGC5oY9DZZpI7nEb
ORisJ98nvJobOQyfih5w53mLtVsdl4GkL+EbxwJiDCJ1HYCbDjRRiIS2q/XtgS5B
4sf6tzhyZmDJ9SNi+Si0CA3o7nkbGPh9lEbW1ALHDuNfmC15/RgS+rXf3OdsgPOH
gMrnc8cujbwpd1OCcHwiL/TpUNUVZjo/dyEKK+vujyC4WwSRWXi05Mj6vUKKlXX4
zSPLkgsTV1l3QiDQ3TxUj/QyCKuBoA9LoKEKEPZxMof2LRK8sZbW4luQWVZdbboM
JqJyqDt4Nqphmzcuw6HYAJI5a5OHjgP9+J2Lex9wVfWe4Tq40SIkM24MC2NI0MeB
oO1sUOZFP4R4VEzkTlnV2TdYuTHWC9VzzzRDl7SJdY0KXQ0IKBGpEckh146TLDih
8EhzFXVYKpajZYeWBEtLsunb2KCV0gzdigcUGKzOdymjzeVUWajaM2e0d8a0SQvB
O2uhqFpELMPNoCRNgEqnOfS2oRAcxMuRZypCHiTUx0xzJwbh/XKAGCm1W2Hr6fQy
4uBJCmUXPHo58XR+E7T1iPGww1YtWp7f02aLsOegA2OI/fOxmzyVwYm81uhLWvCI
WIRlDpRtJ+IbJOTW2HBNWtfbdU1U7IuRlSRf6P0G4qjminfaQV4cfrrN1fjC50SA
3Aw+vQOUv54zVGhaSSCNA1WJZ9Iht2439z6QJTHAYeAvWLTNFfvY4MXHQF0AxGXH
FlZ9Brl8875Qj83fHGMSrStP3Ug1rnMvVTqy+VQRYExwddwBTP3zEGMnMbsoNuOT
kIHqI57d/RSnCYQ4swk6HnFPGi/uyCjbhNR3ZPJ/WM4/YX7k6r6Doh7s5fKQYeZH
noE+3qIOECrzhx9dqbehQ6lvqQFgK3/Pv/McRDSHW65S1RbLRt9FQjHZwAy/4eZk
brq9L73b3PmcFzz/Q8j5GSm7tNN0fa8gS7nEWWt1Luy8BqATsKzIMUP/2OLo05uL
QcvBR0ZLVp8W/5fhARLnhIiTdUAWoLdbM5zYe55AML2E1ChhGVmEvM/jD2lgC2je
+uV+Sz7WmoMQv/hIHcnRkeeUaelIGlRrPB87Tr6ZHWuLwU22GhXQzi1hoxnpTajR
EVlyNBl0ITmtmv1DlhMCYTAtLJvFYTur5UW9weaaEVgQDLynVQA9VVaik9ALxQK/
3lOyBAaTt3m38B+qLovbhiuJ5+IWm7WnOsJmnHFT8B+Lw3XBPZcc3aoFgXmkeXsx
K+c2ZV3+oiWZIv77bWHWu5rojAqkaawwjBd2nwqbK/5RQCIB+GoNllE9z9n3TTbQ
cw2cFWpkyxKou1ymHkvYCfir6D3PG/rPm0Dz+45VeEvSNzbYPLMrnzVlzCRbe9tu
FoVbo2+r/94YsFMzkBuRbsPJ2hVvMbA6Icx+GzEOxIDtMOw9WPUzFGUjluv/s2lF
PXxKF724flupuP+KVMl2kXqjEPDlg7Hqv/7ptUMoyY7hDl2ZA3L0WaXG4BmFXrYg
q35nxnzQX/eGOC0rryr/OgdEQASQvx0pLkFxUAFqiv329JoGPuZ9wBaCRsuyIkpA
YB3pOoTFKw2dc1DnspE63UmQ8qG7DWAXXJRAvoO531xd0xzGtF4OY8SG/dI9Q6Hi
SCLmVOMffJSsP0dT8COFD7OitVw8nCissG5VVadhUijyJhVpCa8mauwPDt6eib6P
BLG2onHPNkmrTZ/jvusCvC3+rYxyx0trCH2g1hbNx4fZ/YvrurphtcIts1MqU+1o
IqjiPoPLcVQ7b4ABnn12PZr3WgMF2X+eQH8zlHkVUiGm/hgXmAVVTZyCERJF5r+3
SDoWjsiGiGukZsMfbh6giRCRFLu5sxzBDuTjxIzA/tm/S1WTsMMUVG/K6DbVovaz
246HTlfrnqMDlzD+rmc0BFfS4AvCw24rHn8iKHuNZ9kbomjdPbGCN9Qg11nDCP++
nVH2CzgzSmSp/To5X7V8hI1QFmmIIyl+hZ8qeegD17hUl470KWLQUJhg3HqVzhen
sEaOKTuTeWiiA8cARPElUuUGg4asHohTHP0iUbwEaPW9bxCiFa3uY5a5nXr/Bd/G
hyzBr59sa8XCXJ/+C5g571/U5vcojk0otDBEIg/OrjvtyzURgyAeahALn7YaeIDf
okMpz2Ub7AjaHS3l4On7WQg8HNXRyRgAvdLV5YmizrLQpwk0sXYShZcnQUBeqFEa
Ox5GqYKnyd2UtMgPbLfrC1dFmOU4zwRjPIopYy10ozL8azWR2njR9BtKIgAwxX0D
5Q+Ox86PNqOuEhPRf4A6eb3eg8zgd0W7usjTsFe6Rd1Dov9RUGt9DEtTA/Ob0TPw
UaiILe6lprPOxT4RYtQFvQTqOcrGBCI5pxZKPfnGVJdnhoTk0uNeikE6Gh6pdz5h
V6xhM+xxCA7FrPUnhtfXV1mjVAu6YNV9FqU8+3HB7gPfrNU6Ganc4Fw4D6F+XI4T
4cAbDTVz0+0fC4lzsqVLOyhlqlkvqzMFvXfUcp/39sn5g7jl5gDwW/S1QYkj2Htl
Nd+KNQ09mUYqUXJKwqO4i+K6Hy6Kv2ZQPLNQPn2KwOEqVEO3eHicbfOlm+zKiITT
vScF+Bkv4bThUyZ8qs/2LfRdBF1PnO76QRWTEdvYnaDidziwiA0OKqBjU4lISrgq
+/JHpPFADcIZYOp+m2N9kFwDP8M15iLuEZCfkQ09WCeeQ9ooDFYZs6D+SP8bebG2
qjnf9kTx0mCnQVOOXALDLH2SbG49Nut4Wrvilbb+edkqlnqe5xJFPLN68ayf8ZbX
ykUeG05qxL6HD78L92+9YhZkDzRtaCX/1YMjG8S54LnbccyoPwrLzgaEBnQsYz6j
/phFEfb1/BDHKq5tpfpTF2za+h/1NvTIhzLKIrnczQoG5hWQ+UnYcrL6hkpW85LV
C1PQRhKhHCq9rsJiAdWbSd0pR4To3oj5IjMXpBdyn//qn3PVdWPB0TcEZ0GZ+qxx
H2ZCnnYqj7Q5IyoEeFT7RUKm5ElxF2aZfokbwmCqADiZJVsScFhE/Be/v87Af9cq
ik5XUO7vTjwjXY2pC4VjIgy/8b2MbNWvTgD4cZ1h/Iaj+u26v3bIvPoyl5UU/zgt
wDGw/dEYOG5SO4w4f6uMFdAc2qI601o7UM8uoOJgas8IIeYXXiE1bWBs3lJLFJeB
VzDqpiVKfGRRkoCekx8VTvB2Y9lhIgUtaFdZ/Zq9N/d9QqGE1G+EQsuBojC4s/+M
rxxWi4aeryyRvEcd5Ntxbwq2FPuFqPhGftT0KKL+xSlYqRIycWO4jq1RIdrQhDA8
0c/ot9mUrzQyqTqPvC53IJRRj1uRsZpBQ/7BhuE+Tdp9fxOHnAdFKsNe5a37qSGR
gWgwAodK7odexGDsHiLMhzv7I33MyHvDqbYIVBqVPbgNq/oF7mpDB4NcxVgWUjb3
cke1BFqBtUt4C0RczuW/i+GFh48l6e2cHcw0HnuDsqDlkRRtGNQmS8JoYT/nlklb
u0yq13y2yotXLwvQ0YVTWIy1Ogqeplt7V+DYlgup2IMjUzfoFuZtZuI/mm0vklWF
ttJ/p/mtqpLzT2QkmqROtbEqU6sIk7+z7M7TYY0XEV73xduxhu2dTZt8DegYHtTk
fTKV3uCj1KjVfOPI5r/xKp+jVVoOCJz0bnMaKTOjxNw//JcIo/uRBEQhZa8QvGkE
B0BSVMtpMLTnUH5iudtNH/cwjSQwjuubGAH2jkIkPwJL0g5FKBSXSkNwoXcmhibB
NXQMKWziinATLT0y0mQERKhS0lRrM7Ba/7Tza/9bB+0DoPtde2yPOclBj6oXH3Ac
cyyIg+sF0sVdD8DHLIT/rm+gSsW+gVtqjMzYftYgBs2TUX5eVpESl5pQuQlifpYn
43wgUMCggHsMWVCf2vWQCvzGeyOLTsbO6jJqzhtgzRu/U3IIZj8qTlyOk3LCW435
QBeF8zJfSfgPSwvEFFHYKgO2QtT3FC0vlEzFudUIzpQaxgA9UwEBoNDSNr/jyqcL
t2IUWGVNeSmcbUkRnyEcI/etTDQRKuyvS1fwZttDnzvjHBM3AZstS8mIekcghqCO
xoQGQZI/Hb5OA2km52dHwjJeF+o0JHpLRJxU9cdfRriAcDYQ+gtn68PD2kyvMydj
KdBExDfsIqMxH32yi9CTEpflQVbOZbCsRrYDL/ueQkEXZxRfBaRrVUPDiELzwr1g
MgbsB2tG4BNWQlNzQ5WC+hS82tpRU9Oavlszkt8sNW6TJ9rAvTuB/e9QU2e+TRaF
c9a1yPyolYdLKD5dTjo1BUTkhtzDEjz+Pvbid1eGZ5OA/c99WRs0SMH6vyKA49D6
+UcT3eoddslKLaZqy1ZfmuNdesFASyz7LBS9b2Fx54XA9sXc89iuk/kUQ2eVtS1R
syxwWIpDlRD3bQoIy9bmyXoAyNOOtZZ1FdRLMybbeImvoOwgnHhLopBatQIqD7oc
xp9x6aJl2J+VsVlReDTgn1LaFit7SH7H05jOFkBfHUciYrKoSeZ+pwjLWhMBzjh/
GkeAoqNNUZobI/6D8PsMAHZ16YKuCMXdP7vGf6Tg8jlJlvhfJ1xw8jDgpSA/p2Ay
I/LFHHfwEEqqQ6h+ZRyec6HuBTguFfy6EFwMI9vBP3pPg4RB9vkQy2LGTY/gBgkB
5Jo0B/xWxqPi/bZRcxV5GICP28Z+lnWCXoXg+woPyaOmNRVN1kiOKiQFZ+G6TfGq
FwkouGzZ6wpUOfXgCbYO6oHXSyYkguNyjop867VyZ+1hYmvvoYipJGPglI4pIA5F
f7svppIKgPXK0WGjcAJOHsuM9rrkxpetw3mAbZKuao403MD2MoeOlfqBWkEhA+WE
01mBhW+Qxzu0f++9E0OdtKgzt9YzLabGZpO07nWXjOvF6mnqXN6gBRVscHSI3KUW
NTTE6iDXSL9AMpsoSSVfB4f/Ou7Ot43FnMg4LlpHgsWZG7DuZX+uJ+pO6r1dxbwY
2Rj7L3K59ekB+Yzuc9Ubl8O/VFH4W58EtyacHJ7za7HlrP3dOommIWnJ8CIhVnt8
7LXg7qSA+fNBxjTzYweaik1/E1dIfQ731PZShnVG2W9lSqTU3AQC9PpMd3Vv1AW9
s06gpuamcfH9aQQZzoD5SFZOIPPJtcAqs07HZlM2oYc/4zcP5tKgZeRk88prvz7s
1lDeWUKlfdaR4FxbBQBS7D6AQbdftEfN5g09TkIjuu4a67tpx/W5N98SRqSPvgHD
dCVT9a5KUvS4OVeXZ+4LsYdzsCQI4ytYbtbl8KGfFr18zevcdPwoikf2LCjhiQbN
d16ELqDl18M9I9UuqdhUYDgxwYcGRZ+ptcehtBF4w5UXjsxhH93dAczccoAXjh6P
CGnlJj8iE9ZU8/64Si5fP2kS3Oa5ldS2o9kplWeqGV4zzb9uKuBNDw+r2uIYk9wH
LCpB0kAYXBQQFqe7dBV0tfTcxAlc5Ypker8xH6jUT7A3jvowepy6HlbiotZEbJWC
1wAstw/b6IMrPI/1PA8FGnmpXe38IrqnXlE3EDUty6uoZ0QxJokhWpaPKzfHhnyl
q153q17V9QEl0KpaxjQLNYFV4TGIwHCIEviTwLDwQvdi49IbLYdG4jWRb4KREY0B
OwC/0V8yKj07aSqvKgDDsNuaOZkZbUPC/olDrlZXHm66CyZG0aFdDAhzLihmrBTi
SEWCLlvpu6vB926bV3tXeJOfYV/tCPjy1HZzG3XqWC+dKJXvhPXixkSS+LsLp0Op
eBZVuCa8y3RD2Qpw1kQneHu4GWc7KnXVmZLTnL6xKPr3J+rw3jlZRNKNJ1rM6hEd
vsrJdxEUCM9XM/AJqk8uLo4dY93uSbo7QBfes+fp7wOlOrXpWzV9SnZP2b//XgUT
pbM6Ixu0ai1+Wu4FenboXTUxRbtMXZjssTwtPTI7QBvAcs9fZM/wfMYVy6gcDryT
4LTT5srQ/MZe2e91IWo6hprJJBisUJplIUAvljJn5fiP6XAKCi7RVLc1QENvlAnz
IK4aKHb0cm14q7HvKBEWSVTZlGO4rYrW28ZT5lEP+X8GS6tL9f1BHihhpn3Lwo01
PaKG3vq/PZlohzY/GHsFLim7VypHJanecbvZzNlYXDapkzc/moDNSW6x+NV15FBE
F+53pQKtXo8V9pNWXSS/iiaxbqu9IppP4dUUbUsCr5Y9bp55FvU3XPqudWQNFwGR
57bDpXd7Ke01AFN6/+bFuZVBk2PYe+gOWgdmXbyRpNg2PleshRgdIOsr2074B7pi
0HF0I7j25i6l2UNAa42uBJjAgNJYLdGPdSsDwU4EW4j7H3UA3zyalu7/kQTARwZB
9e2qU/545titFs3w7TpBVT1RRLsvUUDVEjQz//51JDiFiSJiTm60NMtw1w1AUxDP
+1J2Q9h4hLCOWPRiHqIWI8x/1SnTfUoC/5MJZleCv4rU+2LtKhJPISRDRaaazNy+
Kd70R/HV5VEU4n9KaExAB0+COk81rNxgvOQKGPI3l0N/YYss5GU9gcjegJBUBtZU
BS+qXOUDtjB3LDRm9Iqqloy4A44QVpn0tPPzXF7voPF/CUJizYsb9zdVJhdczAJI
QCYgDhRkEzDzD9ESegvCUYyqmf04eRkxcoFwqVbb//ka7xGO1yjC8EGrPvkL6+IJ
9BDRJG7bjykjC8zIyAxMSX80J1rNWfdVXopbhRckHZYaXJjVWNPVsjigzkBx1G6k
1zlYYxfNcWLuYQL774j+NFBiB7jN7YFb8mr/nhBv5R4BuIHEegUE0Thbtt2G5Ohl
pM8DltwCAsZdUQNSUF23yMlFY1pLDNfA7Aad54Por50mpmPPIXry+9jSCQ7B2kPd
ROmWYL4urvfejiTSI2NVZohO7vyecD8hN+erWgZ0gY49iIscGyoNidrng6eE03JT
Q2ZS7FnOd0h7gDrXo/hpLIqYV4tr0fcnKUOj3kXJ/hLlvi+Mc1/etwjVDJuWzxJp
fDNmKtmjrVhdYe7GqtW92ymfGQZVaIfPUb7W4tW9XQNrNfXKo4vXJ/Jp7l3h884X
RBMiRq2gkudUT12Fcn55W0gi02V5XDUQQ/BlMJlSZ1+nVNLlPYXK+LlTopukxmsJ
HvUqBOLuxUFwkrzu8BHALBpZcjCJSP/aocAapRP4jdq6Q3gevgL+Ygs/hSKFNcDO
qxCJM1RgpvMqzv4L9hKD/EyeaH9DqfsDN7re3rVWq4co0TsqCzJUSyuITsYlSQX4
V+cPnAPWZ84QZ1BXsmW+/fsxJP5FFTAeVmEjfERhOdSCk6fovh6ICsCo6al0KG4u
bpn5RSJyK8noIdOeykwhSn9s9OZgJiIOQHaP4u6oVodhyDsDTjV6GSBq8rvfY2Lk
2SmWYeFtmaSK6v+HPZ5Sod3YDrHqYCJkSWuoMLAqjOzmcoHIokJQA1BdB0jIuJdS
L5flFih5nxs9cSByjMlioA8y12gC56wT0TPQUpgGFPdScny/HJg3FE0xQA7XOxA5
+kkvDeXL/eHK497Bw+WYbypeVz4nkmWPTRCNwhPI/YpBVitVX+BIodPWrbh3MrAc
DgUQ3lJL2jXChCxVm6TCp+JocfPQJzZKU51HDghdCa4SDzqg9qk6ItfL4maGar49
Z9jA9AzMr0Udb6qtVU3LGXqHklXi64bTbxpBQ2ykRFSWFpydw1Ki/WBeK6ZHhQY6
QAU1JGnPYJ0q1xEAnPLqWlGG0kCL2ZGDsMk2Spes5VMdt+D1AySYPlubX64aSsvi
7sNNIXbdJ7Jr+hldGLMLVrtwGwW7BbX9kwtES8Meg8Qgs32L3vOWkODXFIbzhgXt
WxBU7r4Z8W2KWJLbA8c7i7x9eAPYHYnEVRtGSfIW4aGUuM6otzNSJFWJy92p3jfO
Wyg5MjoqJLyBG6PcoNS14rUDsapqsv0oBKRx9KZuBEnNGkqRXL/uQn0/hJ3o6lPr
QoHY0/8b7G8kxoQSP9WaBYFmb+BiKjSQWb4Z/N5hfkwNfEVsJr5kXqJ/SNvlsLOV
BpL3fdhaRZ2LshDKRSN1MeThK/rY9UegH3MPDAFZklPLo/6fsL5drFNmnrXmwMiI
liFe/++E6BzqMvt2FiQQOmT5Hm5UV/0MUJo8Z4JJXDSz0U61D/zGFODzNY1MZuWD
k96sfyvELSxu844LlhDVEXu5DMJMh5yvoFhYuIO9ynKAsQr96paFXJQwvzehf66F
mR8zwwATFCeE6MXbKbmhsB1aSsTkphr+gdk/jyacQPHFbMpzKno8G1TKff2xLPfg
OSkCYGlRChNZChOuPk8Dc/vUO/A1cQfDCd7M9gt/ACOvfTCLNVForaHIMsQonmmC
M//4jbhBtDfZWG14zhb76p50VRLrQvP3n9fNMPbGFza/kPVl2UVE/4joXSzFxojA
LPJIkOIGRxG/RlyTjiJtamEIsausX9RuZAP17Ibj1L86oLeZc4R3Ztkwr9yEdJhp
LGpJABGDMQqf0d+WTdjBWBYeFlehnbPO+OaBSU/G4PhBedpVDi0a+w7JM6b3Y9DZ
3zGg77QmCnvWpB5/1v2dKLWCBDIGRCsyDnYPK2sAtPPk3j2k5ksjv0yI6xVJieLd
1NErFWgsbCM0gO4jWgDQNnx039BG7k2ejIq4mb/tEpXulKoIZX/eI+J3woKcA2Nl
EWy4N6OBc6ONYnpQku9qY+hsUMucDjvL5193Cj9iBKZOxVhPntFrZsRcIkQTeaog
H7nQC6Yt7OhkHFcQ8eB2Mm7E6cFFfGJ1hXzPxft9CpjNFSsFUcRR/e01DwRTysGG
QwusTwn1lQXEckDPgDLQnJqsGuXh9nbb9USn8bz11XIAinXHsTCeih2sjJmO7c4k
qhbX/UUULsCzOGPXiXkaYaZoQ2wrQudsYDI03F8CeMbuYC/t93CPFMqeIqWpxB+w
30e7nrHdAoGK+ZO8tDPXMQXaKExeUo6RECSnig1rXD/wo1axrIpq9giGOeDWxSqe
UxKV5N/vMXNipQg0EcZ+wkOhZUKv/r7r6gLhBGD2ssYXHiOKmndJMJfkoDJOxG0C
kv259beF6K7dgvRqXO2LAVEY1yXEZ1nQ6reFbgdtTlsddZ4UUo288d4JOvBxZs2h
SEiyj+lWOIbTfYfEoujRfWSVcHTQVrYexAPEaYfIQu04fQZ1D1Uil9QfExxPajh/
+C/ZCBqWS9+E4g8ISG/neo49lYI6kZnpBxGiZnhBNP/UnbfcvdY2edui0/SY4S7V
vuyjJvqf2TC7GSGCASlrgluXoRiTH3f71GnZIM9s4UenNTNscDmCl3ghkiVY9iv1
p3uPBgmfusexR6GsVuPZGOJVMLjk37MqERLhqnEZNeXO2e9OX3DPDP+gLF6EyUMU
VRCMZVCy+AjFGZiEFXD4yOTWZFuJsWZ6zpILQ447JEYjcSWwo6I71ddaWNV1TZDK
nV6RA12qPZnD1xOkvGdeZu/Z7ZQxr30BWxkN7WP/WcveEvCoiMFQfDl96U6+7Uwf
9ERur1wg3uGANP5C7e4Qy3NV4vgBUJiapK3zQrHHE3pBN+RDRFuJ9DQJ7MYW9UMd
nFOaBtTP0ffF+FpTyhR58yZ/17/ptsm2AObgudUsWSnsr/pslyP5PJhP0NG1ssdA
f4W9uZhDKJUxvB+Y9YZmHPRRCLKOvdCdsQnHXvEufxcs+WrhrYqSkOwNA2mh25bF
Y4MrVqlBj7S3AdYHj18VPOIimjL6Iz/aTGZoMuvLMVYHfNBvYxfQ5xxzuuuoDi4m
/IJBpMx4MAN26Eng1TLpx8vDeHzg1CVNF3K6dLafvSmzcEVJX6d0ieVdF7csGSnE
EonuFoXOeuIKEVpxs6h4sgeSDa5JRoYd6Rn85XMBeh1b+KdTReTaIl6CwYZ/B4Dc
PWMXkpfEDjqEDfOM2AjZ8iUxGyVs0/QOAk4rRpfsTP3Yd2ng+M+dYi2aG49UXx21
eR/cmPHPXue67glTVYxeFtmoGSiHWe7ZSkQV9dlh+cwRjUAXl4UNMC46QDroQEzA
/LHzw+AV2OHZ2GKLldP8cqrvw6EEek75bRzMAKgTjTwQNqwdKDoKhGu4XuYVZmut
yyPKOIEVNJhZkx/AT/aAc38KwBgcwWXYzFdTIO1n9d/7yr6WucN8EW8EZAb9abtN
xMKsDYN1ejRf4QVPe+n+d0TWdYUwIoFXsbdHZVj+JffGfs5Wl7Imzqe2EbVp6H+p
z2pjzBtHubpLK5+T+02KWy6P8fD4xi0koHJ72HEVDingNhSAXXitgtb9b7tXGJO7
hdrO4A+XXJ7g8jgwahcBz9AxpCgkjfl1MTgqmm8KL6mL6FsLWXK2H0S5QEYrwCEL
uVz6dZSTM6hpzaY0tUYVkICUVBYV1eReuCr9wZLQFbZSN0qMHJvYaOghg77g/6da
ohnm0/t4wbpqmOE5YeK+PmLmnX8VaTwv8P3ibNtSZaB/MicWo1c5Op6XduPSpM1+
yBQAcL1Ba5g1UEjGuGcn/hvPVcBAErF4HoA+KRdOCsIRriduhorDEcTGewpLREUy
InGgXuqZW2aOzenCqngYwMK5BJoYc8u/PZuA5OLl42eaok/gJjf7h+1T7ZgyjosB
CzmQJwGJmtkFZiXfRouzHBigLIAf1UX6XyUMLJ/Up8aD+vycumrGhV9wXv8Zjuas
d/Menx0pSJ8Szg4dkXZkvS3tiDewbfK/S6jqqnefMRF4D2q38OLPISFwoM3DOQC+
4GDMZFsVDypPNvcAAUZjIgYRPAKk01fm4eGDEGI5ZN0Kd7n0CtusgdcYxSWefBm+
pTsci1DlcMTWpnP5qySzqRWXnaQ+7WJuX1HZL5ewfuG/qwbcl/2nG0c81DllQC9z
MbLmMKkX5hXo6WU/bRzv96xaep6jdYS2XFe9SceVrqc4ucHWvZxiKDnu3BveNFmY
WgUy2VdQYiJGLdP4FNecsjeuD4k+nWmQxJggXNVpUmpFhxQCAGAx0tPFm4/hteD6
20+qBbkvlZA2JAlsi2prUaVlySrO2K0rXn/nPB2GOj+bjuV7mXL76XFywmvnfubG
9b+h7CE18BUxtjTCuAlHf9QtgseSNkHNk4voTxjHxUDe1L6pxzED4Qp305EO9T9U
4Y4IqBFB9/xOujPrTidY/QKX7bdIP1ZxMxKMjy4VE+/mMY2M7VCXtvyeAHLpTz6C
YraobJV+u5+81k1WgfVeBmPcT065JsLp6YSA+lnGb+oaDoQwAjFCkPj1e2BxrgaD
OeN1K30xSs4Ku+LblMpDyBKFGX3+vZS0Luc24xXNaIC0yhMKHkhM8EHThZq8aTzE
VoUcR+ZFBIpUsckxajVlPosPc7bYOfn2NeENYcLv1QgxK7Wbi3OE/V/YON5BbaCu
z308YnMjpWFNr7v+Y1PALt8iDrhyu8DjLFBl0jAf2mdh+kQBE+yq+vU9NSp/r9EI
W24uvaRpAeKEE+GctlPWS9Mq7Hl74wnxVUHOp+VZbkmOyhmbp3MWofoUtdZPD1v3
Ip90RCDRibmDGNaH12silGG3ruzgyrRbDOFZkooQxVWUTyUqEDyKJvZU8z6yey5m
WC6qAt3EV4szoA1/RBW8o6a8oquUPyCRTdcjmvwKwo6HSDY44KusGaR6Um3PIDjq
HtP0ZX/okBQ0qcWEstu+QaArumc7HPzIKm+mdypluRPv2u7CAOvzZOWH6WK2XjpM
C3gAkQmkMOIAp2eioXQ1NqsgmNVucrtuUvNyU1czn4oCFFpadbkXILCZHLSUPDKd
zzndo4hpxBe2BMkFWf5uvjKPPf04ngrx5SfWRe2QSbWU8rVYEJRz3m6/toYahmMB
anQqNrgR8dvRyuVw451xM0FRMsTwR6ZGDke6RZ/xZRD3W1CDBeUlOLjOLMKrUyGu
juZ9YuYQRsdBYlB3pHtVevJU+c/p3za/NrWSTFkDk/FUvq3Xdjd2rMISBiN6aY52
7siam+u5+se3izBCTnVVzrzOriYTgznwQ0PFTNOiCg6pmhJP194NqPXJUnYd76wU
M/TtBrwWafNf3yRpvPXxz0fnYvShBdCtZqGAQhSnWaZZi4kuA6vNvIzzI88LdUww
sAEJnIgZrzc2jXCqtQ6Gc01hLX/5x2yOvvmezF/GFLV7UBr62vpDWz2fAkEw2y2K
QRyIzmWmqJqs4Em80yM0bYkAYduz3Xx5uszdHOCktFCuEsrB0r/spl26z9Hz8xSR
/3gNTaQIqubGltu8QhP+9mEbrr2kC8Ja5bN9rpkMrCP1rOwNEYBUhX3gScOYMoZg
VO0IgzpuRSjSutQprLGyqr77z3ryoBYXto5wYZw0eAPG44XBcw19tXsQkdUYcXBo
6qDnWPy3osq/K+iANyf7v0iHk35ddFLsB7+hNWBjtJcds/5AoYgDFhTOAUnyP4+V
p6PP72H43H7nrbA8B820D019gmckgly3Snjg9ubkUtZY22PP73cJ+hRRhmgOF8vt
xT8cSxPnG99zZIGtczisRicmXogoQy78bfFGfqMSXSdaHZIu9MVSji1jTmC3Iigr
5cn8NNQ81IbWiaxIIBaVK+YbfPIkvnUzhUdk0KxuszjrmlbzMJLHe2Whvl8wbyx7
kUltfQQwt8vrDPlXcF5lHj3/BU55dycD/Tu8Q9mQcrtcWha+23gBIkeGeXgEJiWa
MuN9HGtxeUvwGGVlbJtahCH80bsfGTa4eG3RKOdf+2w1MKScKQM+dX8daIvyobzZ
cQQGbJfQ+4pFCzbzIwowIo7tx80Q/IPz6GhsNaodYwI6Ru8S8aKmBUqJkRQgJYFp
NPvdGkEgIaMFAvsfgizJk+iIEWBu2pm/hObiF53HIA2StpxyMZt8Iu8GtNfY77Q5
7H14ihf1hCXQldbv7D72SBArjfWdIlz47s6j8xNjLG2jR7QcsTvSYUWNNjY+AdDn
5L3kxdWfRrUV8LIsmPk44oc3XZEJepmJsvRn6mxE/kCl3VenGztCFoy8GsNgEkIW
cN5Mp6gHi1RxOohHfV4cTyD/sEL/UfkWRvAOhRlyp3sIM8Llm99rDSy92N1gExph
cjCyFOo1kCGnHgFSSE9Y1HPzo4kJeiviGz/1C5Rtplf3nKtNvGLrtwBD4FBGDDWD
lWI+rJwKMysWZIWCXe9l2StaMCMFxJHxBdK2gG1ED083QojS3RiLPMdOhK2hP29r
irGxUs7nnJbK06/3g/XV06b31lHBqkcQ90nO1uNhEnNz0CczLr9UXv6a8V5PANS2
oNahu5FaZeQqux4MAGJ4vQdaTi8ycmt1bJQbu8wHr8aEF/UmrMC9UxFk0MuOMVB1
0kbu9isgA8xZVU+rdZleTbU+W/VIk8blkC562vq5QsfodzTVS69LyIqjtCcYZH3z
eAPtYr2iheqOli0LwSzPXXzT2yLq8sTflU3UJZLNXaEButLCWAyHO3CiD8SbP3Qx
M8p2eeGnuC0DXby/NUSEKBzYGULCDoaVnVJrk6eA42BsoySwnki/Rk+l3IlXAp/V
c46PKh+ENmkDHCDIb098JxFLJXACTPvMg5wKjbEBnNIl4UJ0WHsSoqlZDCp3x4Xo
84lIk8J99ufsD6QHQ8T8BO18fU7FDIMUQ/EONDluH74ZKUKCfHQtqoWRw1WQqTxj
9GSINnP3EZSDlo1xPw1/UVartg2S6UQBjeCZzXjipjkLxMLu8Be+royZuafXnt5H
pE9op0YlSmo4TgajVbjau1hHjgi3iUHsmjDbFrtweDS5qS1T/6B1XvaZSxudC3wX
o9kWZgcza87lRVfuDz7UM3MfF8SMk48HnEa6H8Z+hb6TSU8YmogAG4zOdzaHKq+k
jIXK+H9NbbO7jsZ2cX0X2lnd2xTp1LhxXxbWfsZfd2mygoNVB18cnPzs4yrb8PHa
XcjKECJ8QP8UCtL4Plko2ZX3JTT0WRXLRmSsME1G7KWfpR6M9IqepkUFz+9IudUk
knePYZJ7ZWGrPZ1N9lZQ0Elwz10l5+95IbFRKcijXnmuZ4VbYRgyCWo0DHLRNuEA
1YHLefZtXbs/lN7RTUb1ya+lboy/hPi0HEtdyqLfXqC7DP5AD9iXzy3xua5swoIT
19J3SGtok8ffc5jVqQxh+LJPEz++gFTfTXe1M89WQJcPqOmigG6LWVbsO207OrCd
bt7x3dLi2oQnGaM6kwXeWYGIx3sPdr7Sj3wgjsRzkiKZhV7+0NNAtM+WTq4i9ryY
YTjbQXRpb+SFhJnOzcFJ6gidzlQS9dSg5k/PT1zOF1X/F4UM23YTzlGkV2OLKOeJ
7KYR8M9BfDspMbcxJ5BnqV9YAdjnEujH0uNyQT9L0oWwt4JbhIi46DDlvv3osUHq
EdnLHdLV/UCNoWZmOg7v+FyeGs3hjUHRgKuRmb9l1m5CF08mdtURPPtEQS0y9iCZ
UbserFy9y8BvTSWwOBq1sPBB5G/yOhNONmVvaj+VoT0mvxPmcIXW35Bi/6qACTA0
SUCpEIGNLS6ZykxPr4bnwQ8TNi8yn0zzj1F6NUb6pbPFahQE/WQVMwOyEONyeckG
pK6oXf1DE39tUo0xwnHWwH+EcH+rFuxFsfMevDoriM1AZrOzUcvfo9j5IpjLdm7x
6fFQyx3W4ADleKZcXgBBV7Q+zV8okTXbp5MjflfFqN6Vou6hRxLEmwXFJQ7GbhCE
c1qaX98gZNeeiYYb1U8FB1RgfpC5dGB9jJJBWPXhI08DapSoeWM/T2zJQ5//8zPn
Yjp6zdyYQwfpf6g/DIbGbyA8l/d8qtZ88DCzxtXoS1uTQvs4Ag9SShPtP4NzSHfa
CuR1uexxBSYePlWBOWeGQ505+VSvnDRCcLU/eoDLvZMgr3cODITcniKsiWcVB91P
CLrLW05q7BnStVduHUU7cRWayc2QkND9ZSThKmP2+sbSaF/aZKC9l0sVoXEVeDth
CYsjtsiVELL83TBCH3u5725frlXweE0HwaoQYKT1Lwd98PKOM0sqJMIWCX5ylJEX
0Xbmht7NXvw8d8vsiBTKLTW2TU18nf1SKdafRJloRh3E+soFT/6KvkgglMzwC8c5
y1ZnPF+4XqMjYbHJYaXmk92ea7KfH//e0/V6/NZcPo+30+jnBtdjwLYqAzZVxicZ
MLZxvMw7fylVkUqqcJsugU8Qvd6abtOzH4Kh1QJimc9rwhjUCgJDnIywVHDJrUJ7
DdFCDyvMAjCRzVo1DGjsODeTA05b/CSNyc6oLe0c+Mu+XsqdeLBbwJh5XuglIc+S
y5G+hwY1a3BykHnX1M416h/7y+Dm6yfjYF/4VFHYQofcA5vVSiQIqszW9MPd2FKF
VKky9RT5NvVAmzIxcTIpqxSLy1CqWl7+2jHyDkFOwRMqc0FZHQCdQhhOS8AJtHRf
TfUkX0zsrPMVBx+9Yof4ex+xVxODpYuRjcs+pzvgjDI3c9W/3BAWBarH9WY11QSN
2/8oAnD/J8zul3Jj/6EEGulw58cRUCzzeFRlK5WRRlDI/GTy02W70+JnWRBmZxzl
PjB2wtTYVJfBEM4Lwocshvjh8tTY7piZFQJfdf5VN8my57U5kCm+Ptl44lmrYpx2
k34do6WlxD3epCsjCqCHIy8LRLJO72HY1htgxGL5VY0ifw0J+gCd7mnjxkdnK6ff
XaHDKGPDOeI1CUHpsc3TLqAw0R8HtW5Dlcwy/Ca80+U8L7gAXWTZSWvkGONGqkQy
+/3HZ7jIkimQWk/SW8qqtfdhzmx0bGvmHBKxWznZFs+kq+VnC+IFtxUI8GIwVUHP
OGbcaC6kwLIfx5srDguyEScQPDY2ANJ26+2pLJpFkdPM9+u18EFferpJYSuaA9/u
yw1//EFIDWZDnxymd/DJqwT+DAN/rHOhnvPX7UChnhfOG0GspOrIXkOTj5n2jKbu
jXOYReLabxkvsp68mVQtUdrEsXNpNIouCmFE8Nga+JYQWTWjrNo7D/XIsT+gySc7
8NV1aorhPU87NGBQXacDpJ+A4PVcNXzmYcVKh+6p3iGFnAGpPFjdu2OaGDzLA4aB
LlAnUO97kpmFKNlvlIWgBAoqoDo3L79RXZU6Ve5FaONeWTEphxJ4cXGoWsI2fc6C
2lofMro+427ux4y20PWDeA1pRrGO08pq9dmGKPItduYZU9Gd4flBa5KK/wGgOE06
CSD3SUCdD3gl5zvYVPDWTHnSfjulL6RnouS8mF5wVUXoBOJpj1iQ8WIACTrbDMBx
8az/vS0pZkMFnhKibr9Bk78lCjwJ6co8nc1Ci1hdTfrXe8SwrbpCr+UuYjPTxat5
D7AgfajYvQY5RhFtHcDbBSxjVjETAobl8BMvEVw/H56mQUCSKJwlws1K/qFh986T
QoXwNmkWpiNvAh/1k/9BU+FfW2bFO9xXA5sE4xJUd0EqZNTq7iK/usnyWsByfVZb
s5TZ2dqclrw0M6SIiGpG1DsOXYHbd5yRyWAEc6pdmLopBDqKiRmD3oYZsvNK09iX
YZuY0RFJVgaGt9yTUXL6uzPbxqgKrdejmzbQ3ly/dpEWpUOCIU8mfX8mlUn5n4VC
Nkf2Xcdiu+YNO7RFupIHNBHa5inKqGLkxnFcouDxo0Q8ABvldkfKO224iRaaV0jz
y5zQxiFU8heSA9c1qu5DwPbRuTWeLQeNJ/a+Bikjf9z6m58y4ZFEqJASbMY7wLEF
TcaJNONz7FzJTfsRLT/EZLn7E+jGoEXEJ8MYlq+7PhCkfQB8x4Hizm5QOiK9cat5
h7+iCpHiXBGVuUo1hTkoz7mCw/r3wNncWb3FhL1jn4XmOvHvsTTERUbk0qlXVfGb
6ahu3M5UVHf8S/O2Epcc2eesPb6cc7SuNzYDfuiyKtMyHhloKutH24lHbMll48OJ
LIgMWLxEoYw1DvLOlVyUrAwWgibQHgVQb/I60pUIftgqKdhb7clcErbKoecX4xjt
8MaVf5PXdPQ/IbJ7o2h/18b/aUkM4Ppx5diwO8hK/2EJbqxFoJWtajIReHb1mRmr
D7uLzadq7PQ10ODj41AE83WGvlzKzfvDF2B6GNEAgUSgYvfQtBSkogeKXaG+4aiq
7nddnWRpoDFgxGE4V3Bd/qAhYAMrp16NZG9xazm+giRFYUJFh5uD1mfOp3NnnYtS
1XKyfcGlaoMwffhJNGdr95MLrJTPse0j3xvsOXHIBZAPJ72qMU5BQWM76eDQL3pv
k2l4EpVc3UAQwtNn9n6iLAvOG16osEul/HL48JNrpUUrrBDJvAB/cZTwp0AJ7hZv
hQu8RKWdny4HBBajIKSMCeSk0Otemq8HytaAxmzllMkX6JnjE00TnZKVWHNjMJfm
Gay8aN+TN5o2aSdpKgUu/aUWElgaL2souRTqZuby/tCBiF7Fw1iv6zKTRe8X+23N
K3oFAWp7S6LSLz1hBKDgGz/IyrZnJggDWDlCtxlnZU7YOqeP60V54ZagKP22Qz7U
afMyciq4cz1I3A3UCGTQIyl6uEF4XGNKuFJ+TH445haTSf900c/uVuji1ZGDy9Cc
85rENGEDdiBZldCDnYtMNEkxjcTLJqybKtbQl7aE+Pl2QfsWLW3x05B5ND9Duos9
hpYN+ZJT/l6YvQ1hVTyeogBNsrOzVj8sz7wzXDQLq+JPzekmdU7IWlIAgR5c/CfD
jJeN2CTDYeF0kveEpmXRE33lBKwXiqBxfFbNtdZadn6NDG3zw+9HwYY9WN/dmeVr
M1bCIIbSwc+pYOdHtS6JBPIc2ASq+DrQjNCdzrnzIWOwuJ44hEYdviftCaTxl+NC
zgl7f3P0a+JAcf8ZbuhKpq1xu46ea6yvetQIl1mBJRq03WHxJk2F5aCAWeH/1TGu
aQzcDMfc8tVXHqciBCxucqT64+tvUj1wbOustMpnNXsqJv0m9MsF7t2l/e6Ejbva
vbhzshU124pQRHWxDEXjh2RP7X0d/y1ffKg4me9d/DvTQm3ggUOesfvCi1yhLSc1
Qu1WPBVyBcwX07EFT65/6VU/bwyLGoDxhdzNJSCj5Hld6qKB6FkfrRjb1P4pChw1
ffdcaBQ37oij9eRRarAt+yWPu4Rds6MuIyjUUAFKwhS4P4+2gsh2LRxKVEkUwKvi
4XU6Zg/Dt3YtCZF5G1CvoCnsVhdbBDnxHTC8jf0jDoA0x2SHnePqW80UZlpDvNyo
TESV3vlF9AjuC6tsPljeXMgM2/7Khx86e3SndGrhErcO42ZB78+b/5i51Ih+UbL2
eiWTxoaYrqRzKoD8lD84emRjTyXjkYfpA2g0glLK6J32wdUyqp2ek0aWxOBsFMU4
wNa5E64xt0ZyqLTcCDV7FO2R2gOWjDeDKT7CstCWg0NJac0n8gqMz5uqLgCfiQvu
63qPtzv0OZ0BhV0hA/Mmge6dbg+WmssmPrQmqo7drHWBEFrN/EHiD/u8+oeYtL0Y
8PL3/Ltoi48JRFHkK/VcjiJXe/Zbsy+4pohOR6uTilNT2SfE34Xcx5bNot7UYRMN
DVmiu+j05AXslYI9/bTu2nripvevdxcFNhmEyJsVs82Zwkd4Xo27l3lt/UtfxcZT
cI/5esnACAmgoJjKVwaFhOREae1z3k4BnNh48eHyylEHIynSt8WuMAJJZcw51e0h
T5cq7zqBaRs/qvycNPTT4J/uDbSb0CqRIYxc8aSCS3zCx6gej8P8Fs1POsFtBBOB
JlJxtla9TiqL69iK66FBa9QvUy1JLEgwlYomQPIrxpzc834Ag1sgPaIQICgDz0Rx
pv7igaIp3Je52OyANCDjHOvdJoNHSUGAkGErz1uTtBQg0+F21HNmolnFfz/QSQ6O
XvbPgwyryaJGYrVZMwSaBdiuTJ7LkSOAf1lAXU4BoZXLGHbVsXvv+qKzq1NSDVye
Onjp9ftpEcg84Y0u7S8tiKwRz5usfYzVWayw5IzaewnTAKD1r6hbOe8C2EQ5x1oa
DR6cEI3hFDuQRImYb1ZgO6EQe0zAIKVWbrNKWG66k24wJTTtiBWk4Cults2qGBPd
Bm/qVJ4m89h9byT9RZ0Qxgbs6OplmZ5mOZ818T3jC0ImF2LWfMYaKk0BKkHdDIBW
Sco+zbF7DI5p73Ex3CH0xtFdbbL667GNk+jQ9Om8vaJMSNRdxyiQbFogZoG8nP5g
vJlaoanL5gp3TAgRZVT1yP5/SIma3b34N9aukglRlgUFZ4NasSudPGtriVFbvPyd
8Nmu5xvxj4iv2lmF2oMQeGRlTnYFcHFc3zlkWRYcIYtgL76yefKno1jjlSYu4HN+
UAwK3GNK8Qwha83T/Rrzvgv5g/wgEm3Vx4fcnAcOmyLtzGmtFkhWRXRqz95sh2rR
syCLEVtDboNixWJmK+9u3Zd0Eb6Lyut+cDb4aNJRfOtmIh6t1Cq4/pfJ9fmLk2To
m+jHyGsKGHtAL3DEH+EXJm3PHmtn7+3DKMnFePLFz+uabD4pkBH4qfKkbQo4tUf5
KnJUWkV3T6xOIyS5DdyWMIlNbLLwGKFpdoqLBn6E5VJ4jeSqU7uCJ8tlU+sUdj4q
5eG2PJUaweAuhj9bFH0oKquDCDypsCvgq+kuuEpNJmxqDG9Dhiq552YVq3RWG6Ao
ef3TesOYMHg0G9PuVQ3IsQyxmiTtfUsw71iPJbPBYh8b4NYLep+pfFQRZm6/ZXfV
obcwhyZ2KdjLgeJrfdTdzSKDCwaGFM8cUzDA2LaQPvrK5kmZq0aGw+0O6pd3rZho
2LRDJKuiPS0BD6LJBUf54CCxGO5Qo8Hpk3ENSURdTt5b2hZ1fPZ9HXBxoXZiO6/N
5k/9ZzVegaV6yQ2B6WZSpwbYgNClOJ7wMlsb1AgQtY1oj8Sk+ejjVvzHVem4RrDc
GS1DQ4QkeTNQqn163DftEkPEhvQVdqFXj6qcz0qCISIt6m95EWn1JPs5rzWWAcpl
4PyAWLJPYG2orXrkiBPD2rs0S5j27CRiAuj3kcsbtI9s3OPzayWef/gb5AWgqj8o
iPRRBemD9HPi7pb3XG2bhh/ib7uFIlCfLw/7Py7noHK8NKTGd/BU49JjV+DfsD97
QNdhiAv4o31hrDLXI1UEkvnP5MvgVZzuQco4oDtnwViEaqePbo1vWT++qzQ5oMdP
Ypaa4m1ODA+5FmfuF0/ZqG8UG3uS7oAlektkWXhYiQHOoQDf4IV6bsQFKy5VWdbw
bxuU3DOV7t5Qx6SoSUyTK6A7rLmJd1/FzygKpMdYtJvsYrOCTKvNi8NMk+o5m58o
eKeyh8AvP9nfehcev7nNVGc3Pjp2LnMvbgPWxxUm8PdP7md+9aswTesy3Sc63uCq
OM9LRu3OZMSNqL6ksLUT1N1/Xs/HVE439eJ8NRNYOsPkWvszXLB4+k8yzwyX4jTi
vdjOpeOb7iij9zUCjuXZLcIo47pEZjZZNXdrBdH11h9wNaffpZj0vvuQTdX1nrOY
F8ibbdvsO+qqmnracxpVoNcQHWLcRF4yk5FVOHQRD55CD1wJVQvoialEPL1lZOVr
wK8IEc5+nrzswxrSnU/sku5NSyQ+xdh2jiOHUA2fhAxIDki7qhE2Uv+yrjWWxK8a
QL3z1Wxw9/3cn4lxnk0NPMhZhYogcXto5ld95rs66iNs6X1ofn4CXgWJK18FW+LL
21Rt9gGEsrBcQ1zdFqo9X+kNRSq+AT1Re9IxLFLQpnaZGpCUdwpAQptp/45+umhy
dYMIliQHkAC1K5yrwOusCqpPgkc8V4AZA88YxPAzBGjae4is3yO0O9wAsrrZZhzd
jCYRXYBKp/gBgS2fSuA6/Vy/YN3MPT2mW0KAukUnFBCXoE3hYNreEog6UZXgQHag
sZCCdWgJstHD9x4QIP/pBRycLCjx+giEYCBCk61aLqMuI58JakpulO7h2BRXHRFm
m3m0CeB5K3EP1th8bOeDjvaIOtrkKTJbxE7XqPRjNiwPRkv/XW+tjxYRUuv51eaW
jackoQOBbnHpm1as2TNQCQ404PKZtLNL43mcvlXvhwNQtbgrPyCTDG9cYaWOeLnR
DVc+Ldmci9aeLlYL8HjbMdiQfq6oW8fFsIrmdGG6mcy2m+nzQRzW2Dm1CGTSCMqP
a1xknnZHkBjyUbVhO+vgjVYd9CIf0RyI6WHC/SOm8B+VCYmGw7Huu5qEenuX7h1t
O7aT7Dj3usM7qJcCx5u6J/kx/7N6PJV1CAN0Q+bLrS7XoI/eYoTw4YPc+q91F/1L
uN6g/34G23Km3Bob9frRTH1SU7EFfPuL6e5+hG0k8/BUiBDT/GKL7rnodQ7kYtPd
gX9JW/vSKjJ5SpjgrzBFMsV6E0XUf/7KvgoPrtzmACAnB6vR6gJSiKN6Sd3pT+8I
HP70o4ii0JiH3xlz954st6JYyBowq3wEmjkP2qF8spmDqV3ifosPdBnGA2UUIjH7
CJZBRtEAMnUOmxifmwa0uVg1YeRrf+1jPCi0SbxMWsdVwh09MX0muT/gnN4gcgRL
MeL2PqU5s20Ugio2WI4xpg3vMNMWNCCdpGILYO143iT639yezPioZiVQqFFO8T+B
mIQAy1wnDhsrYG2v6QB+1QdG5JgWGMzUN+yMjBm1BFZ4bXHeh6qW9Bz8Je2mP5bT
Rtz7Socg+qxFq8KT8LPB8atw8q+9u3tnSOgDZhUSRTc2WMPlDOQgH8uD4R60vW8b
UsWS+Wv+LOwfw2bCTmJPMYjd6C+oWINUR1LrLfMNJupnsMjeCJ4+HDZp7LTqMMfQ
tvvfTHQSd0CcoO+KtSgkAKvX7Fi7hn5mdpv0muqpv/eGlvEhPTba4t+6UZWxHjlA
ahrXypNcUb4eDcvkZMcoMu2ey/u8V9oUeUTyDlS+4HHQyqsf+Eis5r286wqay9vU
QBy4pbWx8J2t0inyAT69iF4wM8Xzu8smvrs/7nqqEle8UEpEhF4ZIyGhNwnv6tDk
soXQjHCWK2080LkpQ+yR7tJWsR18AKg9ykzI3nYhbKMZIynRs7H8zUondW7STa/N
rglEjMnt5YBmpuFWMy4+60I2/bY6XbSNQG7Ys7xKFVZ+dBU+gABMStBwrpxNfaLJ
F3q2E9tIkcCn8GgUKuExyxEbUkD8v1Q112O+qlrAPujP6yjTN1J4oUnDQxWN9126
py3DKV+b4kb6c8HUS5fn/tf+IcikYa4vDhhltTlpqLTkBAgmsYzpGprQfkh6y+XG
7FCuViKQ01hTHdiZErxt7hSGjiQomDlFBQUmkFtw9F7xOGfc7BpMY7GTcCgEaKpn
4qHUMGz6nLr5emZzl+K4g7MlGb9/65WX8D8RgaQ5J/xd/76kKEkCmqaExkCjDd5N
85ZddaKhEaC/6oQJiE9AdlMdBJFB3Eu4I4U3k+cQZX5FYKF62bQKOdWcDavw5wtK
4L1SK2IB1wzOQB9xRBs7vvlZ036gdNEgpD8YF1WTjf2Enf9+dSlMLgh78oLCVQPx
Sn2FLjBGXEE0vI9YRCLsDHO+5qCG6vEU/ZsMz6l2/sPwWBGjWWJpFE5ObxpAGFm/
ANiwbwO5Z8FA6mVV+rgTXQ3rEQjQ5HJTfAPsmW6W+tADfQ9zT3qXkt8C3vfotBIX
ySXk2HZWhmPC/YDCXIlrcOUpfGyF7yaqSRPQGEcopv1rc/6alZIh379NB3YHWY2B
aA0VLsqCJhKWzCZkGWKQLduHj5qn75ZbcTdI5K4MNj72nHg7AFm0VXqaSToSYGdX
1TosKMY6P5sB+ST3dEQzMZSpM/dWZRbcoRHdrt8MMnhZtm4jPl9xGFTswdTuYANP
XgLYIKwo4apn+k7WL5i1A1Ok5uD5Is4rnW+Q9lXB9Q45Vr2iKnTYnyya7xQhZNXV
JQLlgyYWT17nahnZcnMGKI5PMcCPO1knm/dTpM5T2k9uVylsgVQpCuspQCyr5Rwt
U9xNxHL8pQU6qLPolAjD6gvBc8UQSSG9p5YoyimESyW5hEtDOWvj5SYkAi+M4gf0
vsl/FNSFwX327NLzD9FyayU5W2wbYRVVXzBmpQk5ogBupDU1j8sfAzFGk9Iff32E
6EJYRc7h79xHWC33hI/f4/pwelIJSS/RFu1z9zPwHNKq2t6LmrtjhfEL+2WboTT1
m0f++fhsnznvvrZNwHAEjYr1gUbyh6BMmJn/WVPX0AUOcFaxLWW94cmNhvtsP7jl
CQgClOeY1Gd63mGA/7YSshav3wyi9vjfXKxzEBfA2zMzkJxfMqZenH8u0REjDc3r
MglnL0vMqEAT6qLF4naqkOpD7RWxBjLLIY21/ucn9RWAQpNYlbdux9xAzUuINLzt
Px9ZV6uxFm9h7GM9sRX96wvPSuzBdqzNXOHkWbyLUToS/RY8fSw/h88ljERk0Td+
0NT7BoE2ixMAEWDFdPj0H7b+wyR8Utwm6jUiYCVJBb3GNdhdIhX+q2TK3ms0IcHS
k1oUKeKrvoOB96RPjHP9QW7+47G5J4h4GWKBXvxkTWNUyH5khSCPxKZ6IZRL+xpm
QQJweDnb5/vGQGd0wvzR5GdYdC6O/FmK6Q8gDlnlbUrQAqYhYKFSV0czLko2xKWD
mZaYceA2GdtZDwX5ZYkLobDANoDHpExE/nG6OmHCGPvKOwqJeRot8Sucfdi9f9gG
/EtEYEz3DfVFNmZnO7CmON/eJuFIIYho5xrmgf+v4G1hDqYGwsHrgp9V6CB90AVA
ez+Uq3oxNZIHeFPZ+R4inrSmTUs+qGY/DsCmydsvSVXD7TyszYH9dCKoUm5ndKZ7
Hy5WpII6ne0e0nL6WbXisGcHt3mEZGPaHcIKuPsixoEMccXUrkYMNBBZ+cM5a6yy
cavBOQIyjBMuyQi8ZK8mrtvMbkeoTJab6yHgiHD+C+Gdp6kTb9bXsSMgEKqEiZr+
PHLw2dkSmwI5NcvvK4m0SvFX4yv6CdO9FDE0c0zVczl5C45uvPghoKpnFp/zBWGX
BEDXhuvTZi6hgsCRA7fERiWImXm5H7hM3ytLFd0SGCz0E7Gali9eIKZDTDZxtI+q
ucRNHhkcahX3LJnQcMQhdrJKb/hm4mnMp0u9gBB+X+R4/tbt2CDHDpuayjP4jGHo
FeWQxsJY1r8hcTMJmsVdQx0jPAfv9xKbKnHZVXMJL/I7m+FR50hw13IbEwEmFscs
SFD8c6VAlTq6GiJXS0YYmOw0r8W0p/3PeNFG5c0QlDv/Qiuih3FIT6Eqq9AIaZDz
Akd+2sz3vL/eeW6QRm35R9+dUMMUDyXXFp3VXVcBuD0M87ijwh5ek5QZYq3vAAKD
YTIYOrP/TvYAnxWUJZeLu00Sm/Fu4AihebLdRNMlIls230oLiGvVwoG9D1yEUk+c
oILa8BjlhFE5MH07XfgkYm6ZEV4OFeGJuyA93Rh5wWzbE8A6WpfwHxCijMekOcu+
AG/ViwpHiqrm2uVUV2UvwFAeK0ZCJQ3WpqxGjLOmo8DY3C40GOnWAIgqFk+uIBBj
yieY2S3vU7mSU0+YjuG3PFdXdc0ZHed74yMiLqUMYZv3KBVBOKnYdJ5Zhz3n7qwP
Hez18meDHdW6Hiz8r9Eq54KVnv0iBCPU1ZEWgob5GEm/rzcHHJ/I1uIx/bBJeI2r
KrNYbZaHAIH6OPVnt2ZqGSEzasFy2NlSsP8p6pcOEJAwi81HNHjRPVJ3rkASwNn8
z6tnKYiBZsmqS1REJWdEpfjf4vapebNMt/OdWvLWkga4D1WJv+rmnZtuAVF0670b
5lHwatO7FzdpkGKyS4Omeg5p1J9ocEWV2oyI2ec6zIwkj9fZTtbFjrjvwz46YATM
0wOeACoY21ld5gyZIVC644pVbrOQOvhsXI9UgjLsxUeTTauD2oOIrvrCZGgH4yhy
1hCmXKpXhpAXVoBdEcX71KFyNwnMoDbHfiGikKjgJpzvLBv8+ZmEDdmkLAfBtp53
GshL/7G3m6MIMkvo4uQHNum3koW5VqJqzrewGBeVdR01E5Mj80vaWNR8+FQ4z6EO
1gQ3lVxY4nTvPRrz0//y0JBHGGkUyVNWYJO2wh4CJ1CB5gdzm1KmTH4THKbpyRS9
bcrtR24X1zSBDPXypYBK1eNS81n0HzNPQg+28JDhfY6nzuKivxxxQ6vlXIBQLPK1
/+U7S8xAk708wqrvbVvmhiOMp+kKkzhr5sBzKT6cAsNCVepV/KcD9wOlB3BNJ/qN
YDtDsQ8lX9jl2jNTIPgoNvnA2rOQEcgVl7dqYMW8Gy2elDq0ECooD31SDGsPr7Y6
Mbm38HHCMz4xejJ/stRkEnRp+X9OsF0ti2ZxU0/TUhNQjccK4q0jBCAwiX9Ar8Ok
dlvclKi5h6VMxmRVoVWihqlolbinBY/iQ/328n/OT0qEHoGyrdLKVxTgjrY9yJo4
uUkU6qFNvUj0L9V9dX1u2lm5i+Vxy/BjwgDCCKUqcsV/eiH48iSuP1BGwVL2e1z4
eao5cIpn4axFhcbdPGAEdoZTy8CFkKHtrcibMj4S35vI4/8CwFtxFyQSQjg9gqiq
l1tg3dzH1Z8BmnKq9iE+LRdilqRF+0/3t/ovIJ1EASnC0Zr1nTL6KRxFvRmXQtjM
oRcwI7QA+2hQrVjMm1n4tzGpG/Kf9nsaUDwlaVsadx3/p7TzA6lZUK9nPI/I0ot0
WgYKGA6xpWfDIHgjjKWfvjxyHeKNggJyjP7lQu1xvd6nnsgBlwTb51chaJnrYMoH
dpcIlpQI5/meM2wBlb2vzZ0ckIno0LEXsz0ucdUFRSmecUk5/bFT036A62RaDz0/
7hbGhanacWdUkCv2iY61CcCZod0Gy/HAJB44LV0xuKyFqGWifn1A+3tbV9S2lgp5
kM7kakWwcC+jZyLknZInvlCl1J/Vx+kODmwcZM8boaL+cvc8EY1t6QSswckyPt45
8MDa/w3RPZleuCgDHudLno9c6a1skq6pYgAjiwnyE4l1u4ZIjZ3hriBcj0EnJRt6
870x480Vs4Ok1f7tvsd/wmVhajiszsc8dbWgDQd98wHeMZZQHA+90M2oHMm7AD2S
uM6O0S4VWHtpyNN0xPrgtdyCbo5jKOUylInit4aiSOTR128wM9Ia/GYwPgM3VX8a
m8kEjYrP/FlImnoxcGXIp9MlpuNSVjfXJWLCbHqDX7+4r4NQw/Vds5GTbsuof/oU
YG8Z1YK2ZnV3WlPqsR5HcE7Y+H9fUtY3+dHoQT8YxoNeYibI5GxqM/SSAEOSXm3a
DQkOidicvWJFF6Y8okdy7Ree85lVwfKhiC9ge6O1CrYPSZ90L0l1ZaeBaLC02rI6
SRmEBHnYSK8JqticqWuikFZOqdyaKrtwxgI0ER/gtEOWs5e1G0Fad8vPU/esqAzU
n09OqXUqv22h9AgogNf/s70os78cDFkdljuVWi+QkTw+SJ1jyP0RDU8MCs9Pruo9
YtqFOFgF+PxO7OB7Qhyv5xhNsO58whVioZgZSprOSQxrWo11gUs3bQY+ouAOBVRU
3RkwRoioOnDHV4jzP7aW/sCcrH8fTxy9bThfXPFnsKf2WTZD+ztZQhB4dgskNair
Kpm1BU5CHmkIuSRZwxiXjDWExOhV8R6gDIqc96hdjWsNEhJhux+mLxJ0uCT4h6EJ
619GG3j3tsnxk9ssXMK1+6Y0UPbeW8Tg3DVCrynDfHSu59UNCjjXaJXPzJJo0KDP
Vr/RiTHBRBzEoz01hnJA4avU+3XyZF866vkM7kDKqgwyI8qxmgqqS1/05sZ2Dct1
ebEuV9at9MFigc1GhsKdu3NTMEORGS6s+EdZomNEhie7FaAvbCB1sAn0f/Li2dkL
5DB37FFVXxpH3AAo+RjqjoCPBmF59utbUBxd9OwmizHCEgMbd1eQpph2M98yIqEo
i9dv4zpggkqXoVbTuCMjoIuK8C6NAcVa/d8NSA1FSFyuuizxtvi0qZoRAaIdDNZm
MD1Da5iCUomBzMZ1QOO4/M+mOvKauQS5HbxXf0LhS+t9l+BSKRn/wr81hVZAwKQ0
utjTDDHeTumfG/wfF04zQu2ibPOZ8ymBmHJzmbr5h5ho+n3GqBhTe55FVghKu1yc
RBZtK9upm9gZXlt60BuieiH5sP9bJ87r9AbKvFLMr/fli1qShEwagUhm0pAJvO9w
+3Wu63+4rPKECTdXbSeSgDTx3zHiQEdUptj9WhyVgZIC0LUwro0j7Fw9aiyOKR2D
t+gK9A2yfaHQPurHD7ziRQ8zHB30ORYsdafpLwrsNQ4eqY2rnOGXmU7ggQ1unLr8
EGpXYy2DwcKMGu4Qcb78zZmtwQ8wBMFfGwZUxcsit573EAPsHN7HusgtNwHIchXE
kwFSCNlth0HCcBPxQ4VJFO3wARh7CLi8AOb0TN3uLUY+eWGxi0zCXFm/aJdRwvgv
tFGPTPcn4/wHFcbV3piw80mwbd9OUiRN84cXNHkjInSvP+DBtaydznC4gDYYMRoB
PdObjcy6xQR4ssQHkjcp/zSxdHb51rz+LGcz3+a3+dz09C/e7tLcjDUa1P4W0FA5
xBUo+551c74lYXswLdUw7JpbcOyRrrtQg92bi21+jwmbIlkTiJGRw0TYVpegdjRa
ESMhFGTjs+onThSnzLPoZqu+zFB+IgvLmMX103ov8rQQuQcWvlY2RKL5BhYUQoGV
ck9Yf23GBa4Vo+7rskB1Q5xkqIPM6MP4vroojYbCaZzKsL0MOjLMi+pmkBJHAxjO
WJsvR851ExP2Z0tzl2rS3L1ne88EBAxltceoiZGADhjKPbKtaQQ/abvbU/jRLIi6
30RJhIkVYtN/YNJpplNVQynOkf4cs8LBzMyH3O7pMAbn93J8ZnurIa79zWZRgtaq
8jP4cYH8WUFtdHZyLVWQ6IBm3oM2SbE9wAsink4E3wna9D6AAm6AR0y6oBScItKV
SW2pL+o4454aLBr0zTvONakjcSLeRIpsTRCxVZJYqlWBdepGKLB1+RnzpRIoa93C
wjtP/1f2Tqm8ZOb9Eeww7wpQmVVuX3LNApPQy5wVfcHWeXk89DfxrSiiwFNGlZ9p
IslCIPOHu5fQuhblflzm51YEtOA5xei1jrzGm919GZH/lQillUfH0aiYiBZPfpwX
lM2oFPcG2KghqIgWvw+vkoI7YCXrhRufJ03fgbVYeWVnuhCjhX5fW62WWtKRNeTb
9UEPbdp0YyHhtdO3bJYtsB10vY91iPo0jJLqFSHNcBZNd/rLutmGUu6AbhkAGako
ml+cN6k7Dt/7GGccf4QC4lDJ3gmQK0MgxpUixJrE/R5qjxPhYmxd+U6jvUkcXizC
/yKlYz+pX6VRyy6jLFWnihP0ouXlp4b2JDi4Say2oh6SHPe6wGoToKxfV64AlueZ
zzCIpgQEwV/9OfOJgv7FygGB2SZBg/JMfFH4PO/pYvhFtpS4WQTeMDBCCY1CA9zt
LQKbt2Fxeub0QVzHnX2321XYp5Bbgt3HIqskIH8t89mEq9o0xykWV4rv70fXbNnV
o8SfoNUkhiZJbcLCgLRwJAfvjSWmKtWW9u6n6KXhe9Fc60s7BCuRjnhcI97QfHLI
Hmq9MLl6ozo9QfuTb41fasEcTin3xIdnWvtV49THxMUwjCNQ7cq5EvjwwcAHt1ZY
l+5afUmw8RnOfFCsKb76mfsSHHD7eE2WqBPq1K+EYoVg6JM/u3grQ9Y8EszeGAlB
HEbm4mHK2MMZjCic4iaCe4lKia4nVlv/B3LQfQU7MJgmVBxSR0Urg7OunSiqjVda
Xcqogsq+hFow+7ZgPXtHIl0JpQS6JVP8stL0wGgOW9mFnNjb7fVpNvCjcWlfIhTH
jYt05XEv0s6FfkPBeeSmFvPPFpvm9+SD56NyeQIvO9ZiP43MQDTaJGu1y6hIyCIG
vyhzoXQAwh4t6T8Szce2gsf+8UuOt21CS87HjX0vXJNQbonQxPDIOnAMugutqLU0
bJb0jiHm4I7THAbeWbTSDr572IZInTdoJuOH/vDoAv7PqCWqCCPtpD6RciO1VjrG
GqdH7OVNJKyx2QwtNvOo3GpaWWEqxyPs/VT1dJOSlPREFVJaf6xkfV8t/XKITOeo
alrEhZBk1jRH6tRnBKjHimLht6fhGa0riQmUJk4lzEG+uy+bOG2Z+rW6sTxvg6yZ
VaE3DGx7UATQOB8BpdBsCS+lnwbBj7iykV/rYHdbl6vfNUbpwNeb9NoFYhl97H81
/vp7NrRrTp/YChQrnF3sK4TjFQZH0ah8k/tB9u4LBDdu5ZcDGpOKMWIjphJe3Aks
hknqur5Sz02l/A/dxJZtL0qhaVt3h/DABO+2YljMhnP6pxb9cIhbAWvLwEiBKn3R
3OFuVzmU32FB82m4NtoNEMRpwlb7vHuzlrhMNea9EgIaakn7B1ZFfZCL01cXRTA4
xzubQigPyZ0yuDt5r6njPOfal6AqmPfre16cfZEGsgV38307FjG2egARmT64mizN
f394lu7XtJSxzodTixIW0eL0uMdPOsGORh2GFN5kKhV0JHDFflaLoMjPP7pnL142
23agac244xyVuw8ZKQ+h/TaqPlC1qQJQjUjx+8hiW5sCsgiuhoXgP8CssqRdYPQ2
sWJ+6gimz2ReI59PI5zKtJ//0U8T6dO01ti8smNsZjPS0zcbP6dAto/qb5T7EVYM
/awsmyWx//L11zZaUmwD3l82Zi9BN8tSZWYGz/xyhiHlQeI4vZTmT/ZQhKusKVYa
3NcbRDfywzHsbb4IgXMeiLdl2zAeHQBsr6ZkaJ5yMK6r4diIXl0rzM9MU1KoIavo
NpJfZ4O4xWyeCx189fEr5fBRGxgZ1nXp66mc6R6OhqUyFKWs3RVxSgPudfvEYQYi
GtTiYTLokwMy53g2NCE4s0JPCHSOXLSvi//mC5cmVXm7iUxORyVO8M/BSrktceD7
fWz2BGPBvcEf1adeOo71PBR1BUaMV4zP1lLOQPhMZlax5sQ3EOWZf/CA3r5G0EWp
O/Fgvp8RYUgqI2Nkmd5jnzPnAnZvSwiXzlWcUR2Q4YA2Q1673eeobRp0B6OyPLDg
QSlwbSxOEgK4xLtL/H9+1T43MPBXCw5ikvnwVDsejntkFLl7dNIUdtP/7oV5DpqG
jlqbQeG58fmBcOsj8LuJqRbR8LAzsrLOwQ01mHLStmTT3XbGe9bQXWLZH8Ounbqp
4lhoXVzUrr47fmSkRiRK0OugPWP5VD90mVvHP3+1erg2KojcJRjDQHBCsqQFH+xM
VbNn+7c36qc9jgZo2YWi3kVDuSOgM8Mi8rPoVYNYWdBt55Zm87In8gAX1kRhyYN4
+8JEne4IiIzOJN4Ij7E/JplMtmExf52Q5Es+NjtZTzHfE8W8kSLF6GAJpWtzJ/tI
+J+Eg4BFjmAHmSbfRtfWJwBBuKoqw+1PrgSN5yuhAaWZhLTAxkBHpSOzgTfCKAE8
Lxc2HMtMYEuEoyvIfEWO74OsXe2S3lwUe7jzjMePAabirdZ5g6qP2HI/KOpOjClc
vpGJuj7+q+ZOYnd6LVF31AIjibymscNAwSRITO4RdW8Zp13/KpFmkZcKfOsg66Pv
FBjplPPFOH/JRnED3c4GpHMymm848zVrdCYL7Q3yew1sJSaiImIO0RiGn9pupxcU
rFSoueVH463VSzWA/jg4RuaN64qjGuiuqvp3XJofnfIqTs88RDLRtGmPsK7pzmXX
kaa9FXjkkviQ4mivWy7RFv5LLEedyFvwxB53M0ECOZUJcvQgU+Hc/aBDMJHAdu+m
76Avygqtcowg0xh7WEBQ+eeCYlxMovspWpkH/N4gdyqhzSUugDFvitKTw+t8TRAc
X0ColVhiBv7xYooECfojweLv8GgS4fnjW0QwkJeGmyFak/MEjD8SCum/HnxnbdWV
LMKhwJVEwxojdEyhrCjlT34/PlGLTsdeudrdjzw9TRWCWiKK+eF822TtZpqFTh4+
C2BUh6VscTSNrnf5+cC6TghzbERs4dTp8jplSIkZYno5lgm+lReK0lLcvYusOLHC
L2VG3SdWCI9WVvLAp/0I+y1DTcywqS+qXRuryPD3kyXiQT6DcbpHIOl7eMfynwO3
eklqbUfI1azZIwVdrqwpHrPYRQ9ytA5X3D9BlKoDQdp3MarPt5sNJS0i59OHPCXg
eUotoBF7od7JAut47dDNMVPlKw6N9hkBJ5GafpUWEXPU13NJKtDvLul+q8BqGpay
C4lGBA4s0xVr0XLOSr5oe77+NkaZ6QEwNCYUNSlhONUVdGa+rOucnuGlO0QDXoTb
uaeSXomhRFB4TV7aS0Sd7Dtr6vj85DOlsYjJjyCYbzCYb8hmg/m13J1GWB25/xGj
J9aGDxv/DNZO1MZFnTDDAo+1JhxpmnQ+SaixXlLunY6a7iW1MLINGHttfk8UGasH
sSkEX3bmku1XJTNRf5diQRhe2pV4w+Y2vZGpiI7qLKSaQTKdinIgbJflAXSlm2/3
5SW+GRKZuvnCKJTTbUhIo+x3xPQRcRrOkh6+bajG97HOqA7agbCBMcDeiX80hajG
AwFiCHb8j19I/S25fgmKQLzv8sPlAS3vAEReaoe/zvKzxFf8+/FVKm9FDsGHfJnk
NhqC0/tGkXq9LO4HSdNNL2GSWfBt36iJaqTnPacibLllIqfB//dNzeCDXg8AJg5H
ZMTZ4JztUjj62HA0S2d2aQ7cCoLQl4jIsYUrnq9MOBplS+8kh8+fhgueIwCyu9Z3
8HD3KUps9oaKQ0KRpYTAUVQOjqAUvIwg/m+bFXP5U4NdhLwL9JonfQfzK5aE+K4E
uHDKVGLZfLg+u+LfPRo6CcYwtvltmtMOsKOeWNH8EXibdGy1TvnEn1pe3KzCm3sN
SJ7AA/noWSVoGxtO06fpO2EThbOdH/kwtMTjC57M3gA=
`protect END_PROTECTED
