`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7iOZw1pgb7mcTVfxajDp//71eO6xKSXS1DcJjqFuxrX5SN8Fw4g286B+J3y8CvOb
73t8eKWJnmJYYTLrsome2/NrGAkv5KqAdoPcMAYLOBYbwFd4+l939UWaHXKJKgLI
iyt80axs418ixCAM8zioP1kK19jNbQ3v4QPpaUx3swb6w7SpSkmFDJiDuBqBVlL4
kmcZNr40O3q/mgwQfrhWzLvG69ijTUXRdyS52croU3TBUJTEgJlnBChNwhKSb+kL
UGme6JLY/rYBQQkgk7xPm8WIPD8iCuPXfqAHiaM0DCHMSV6GX2TAtRDtbQB0X+53
0ooJIMpAz4kzFcUuelUHR+bnvfYEBQRRDCcIClPSVeCONDYA2JPNswKM3gyHxHkH
FbdBuUcOJkiAdwt0mWh4LYlrl9dBxB8ttbkKEQ2BLzgk0Un8tAZ+zgndkFMJL+aT
F4qi853oGAIU44vRZt6jz2nejntSURBbLG7Vxu1YRXyLCcWN/fHrCIC9jAg9DVCr
gHLPUzcCBjIItxRcZf1yvuoVVZHS9jNw+zoU/UaHnzA+4S62F8jXpcwbIBy54yKF
e4M2rb5LSiL+H8eeK+/indCTyWWMOCXBRDtU8yGlhcY0MSs9nIF62wmY49qXvZYi
fPT4kRZussSdVMPncCyuPrZO24Z/tnBVh5U0xLVFK3jgItrxQTKlbLNeM+pwA6OK
WN8ssgwng3LgsbC8sguyvpXE9kIoxXt0JRQQujRhHT+p8BwoBa6gxXD93FyoZ3/n
OkEnxexGBB9WeshzH+h6uw==
`protect END_PROTECTED
