`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38lY1O/u4KuB1BZ9lT4QO75MRtdheZ+8Rrieloqr0feUMCGAuvSY8NwKBEee1S9k
Torr8cZBi1SlGgbtxigP3NUfLie05epfGJCYaBgcodveV7YBrweO/uustJ1wludj
kmGKXq6fLRlohk8uWYS64w5TzPkN9XgJjRVcs6xTSRUtlftYe+LPNFr/VKPu7eMm
0ehmr7o5pem+AH8IHNwptsinvXlBq0D6V527jYtrLJdjLLGslkEKq80cAfz88w5e
6SpkV6iTK2aLJRMtvrDpLbDftnAupK5n7wB4mzi4Sr53ZZ4QN1ticwYR2Ot1rrhM
EMOpWL+p9ARcAIqrNLZ4kvM909FHjjqiN95xEozA3jHFXACTDsGE0uEG4pjj4Uef
qUYWM3ax0gRfrGSqhuMYmI0DUhqMfP48XBa/QaOKcJNRis0oQBjVG/1MuMeRMewj
cyOBO5EsPg0iR7qPpoTx0axuXMKfUNvqkDhT+9wo0CaAu1hMC165LiKVnGL6Bt73
J/JKr6+Kv/sp9xKBfP9xvsd9wNA0KPKhwoD6Ikh25eg=
`protect END_PROTECTED
