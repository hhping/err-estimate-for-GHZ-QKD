`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abkXrlNIp1yzOpgNqoGTKPq227e6ChZUDCIlf342kkJQj8PFy0fltHnA3VAjB1Vx
10rlpgDLQ9UOnOlEge8H1DLafRJp1EppwSblW4RGLFXb6Z/wtHgT+qPxrSE7NV72
xcnc+P2Sw8P52STYMcukxjGKilgZq5GDoVxODrIswJ04LWjXa4JM6xrGkXgcba9Y
ULz9xP6w9NuuqEvfQ/wP5aA6682yzMdmCwbWH/cDS/WbAr++nWMDxTpseHNH6Mb0
IzEF/EipoWTtaBFgXbtj7wka1y2f8zoKGTFqeJgkP8jU67/AJYiGDHVEQfLMwx79
ZEj7iYaoTgzW63PYsJoNFbIICRGZo+oM8WzlHhvpaJtvhTLO88S6ZNXgFG7eFl7M
fhtFEjh42AdKbSdxaJP+LnRSo+apDzcDSrnnQ0Kq0jPnxVYtoC3HsWt0kBFt28kc
STLfS4qFik6hr3UZip0FiVMzRlL24fbr6gA1BbHYZ8CP9adMxyob5GtGe+fiO3yv
kr5PAqlxXO50EhRznRSbNYDMNUjHRkpRnPR/hxsDyP3pQlRAgKXEOiCIHHnZCjOp
Ji3O5l11WusTLprRWraSwQJ5IHPZ8dB9LD8qXveDOjFEsndPKJa5Rsdsr41wzhGm
JTwHv9t2nFloFbcSz4gL3GrcjoZWf4n4cagMP9DEJZJ3lmxaQDWhnJ0zUFTJz4UJ
iPTWJJkqNxF30MQRVcSk2KiI43AxgQygAqW6Gm9Jtr97QwDhEs4JJETIEpOoM1Ur
pnT+yHLHjSS4R46hbuRO0UtrR5PLzyLYwvPZLuiU33bbY03oIoQEpI/a9EEiqTEI
RLdkQPkTezGgz+uo4Z4oBPiJujIEKQgCgcybnStE6EWPaz4XBN4ekJU6S0LLXSJe
iNnak75JXrRCv7XdTpHHojwnaM3VCFqETt/cKAkwEVjOFSkuqv74JvbvpuXS/nHk
2AuBdYS19Kq4ferBFQneC04eNgZZbwim8MaHBILNpFnEuhy/4SsV0OiPG5ryJ/sR
XUutEi+wRKyXK6BD7PK8k/FNpKhnG3edU/m1lyARewF8Zzme3F2PRGpxk4Kw4+PM
h3DzjmtdMD1CJTXm5ul3NJDpV4yrAciqr81gDWy6iTpIpLft1bPH9LqFcUVpZ+1I
Yj+KkfaQL3gaTYGU5BRq+xUadDDGHF3wg6hQiBKD+2I7YdhLzd9hZtsdNUFccIR1
66nxFYDtSw20ARhWwtfYfilgUWKkzeLZQpso/X6GuCC1seci1Zbixxk0TDZZql5k
xPp0AXk5D1sA0b4TzQwAPoIvFcsN7IbwaKBFQWHnvAxUILH/yrRqdoX9WDnGY7qW
q0I3CISZQEphhV+l8k6Yc+o9+ow6oAQ7etP+I6DxHiXM+Kh+Dif94oa7vNNK+Sdh
6XyxZDSDMHhV5XUmWhAuD2NKNsmSfC5Y0Jl2m2y2Ee3xh8uJ/NybUa5UqpA69I9u
7m7lGrhAINCpLGNiwp/Bn7HgedXtkBcTkbR/MH/jm+CYnDyzWfJzb/IhfTAgSIXx
Qn4wv0QCJGbr3YIltypqrJaPHqK0kR/PXNS8DzHZkem+OA5eN/rOUHfDKewvdV7P
9Lxvhv3AwREy0TjBExyDdGy/HctVBeOCpF34inFYpfFxlIQ0S/hPNIwJ7PU0re6I
HtT4Iv0TfRao5ot1BrvUbT5ncCBPAJExJIcSur+zjxpuZQEK3DV/tZ9wh1q3J0TG
1d5LdBsxdxmx2E1Az7Eo/HT7C1Gvd/8rWz/1Yvgk1YN9L8lhmRqZQWZP1atiWQ2F
CmuahwPZpaGXfz4XmPuo+FERGxOz5SQI59FLKjyLtjt3w6vMF9FZu32Td2P2QySB
3AppcE5IfrYiSpnJKtzqdk6eXyg1E9cXvfpEO3LklRibSJw4f49SO3R8IvFKTzwL
kOWCxgLAwuhaPsZp6ORa16PwWGMU7Ms9swPiWkWaTWraV52rj3QDD4ejygtIlXtF
P4zckUmh4Zp+gbD61Su+YfyfKq/Xl6zTDPiuSy8nXCRTSxiWiue5T3vuo8Fxd2tY
mtx2W5GRu5uiyG5Qxblf8mgCyFKLdXiVQ6huVHAtF1yVFZaxErvXr0Ut1DMn+hcy
jiGdTywvjRUbaZqnzJHPB+IEcCP790tZOyhamHcYXVcLISl5AzJtQEVusUPKlxRr
gSAH75OsoduSjTRBw7ZOrA==
`protect END_PROTECTED
