`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dx67wwZppvdHsYHefwjZ+aKxhWMq+RTUtv5KwSp0G03UXmyACs3Cx/50NrIAqArz
iQUF/z+j+fp+JAUQUmr8cdCFzxaaZ9yRBj5PFeGejCESdypxTir4HIi+UyhVR2cw
zbZsxpyPYlrlDjeF1B2l9VumTAevgn0MvSwjsjJuXystYcqdry+zX5Gy9eDsMoL3
6xMyWrq/owbovb987uRmgzryv0APyh0kY9W+LbAOolSjFbxBKugdlOrKqvPkrDi2
a9gPGuecFXdDfJhfNS67iaL4R3meV4MGmRbEn3l8Z4QO0/ms+7lMCcxPVzyM1NPl
t2vKgVUkN3Rgaw0xWVZCTDK89DEDVLrl4Pa+B2IYydRMgvmbV7K8O29iRh/h6CjS
`protect END_PROTECTED
