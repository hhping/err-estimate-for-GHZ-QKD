`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFVf7uSdvztx4W5f9HmCyVRrW/DARvkHWgY0/V5W4HBN7xBsBeARIFL0k+3aoAXc
9oy8foQv8mgX54FCDqqvR5Ad/sO7Q1lS2hTGln5MlM4cAy0OuqKJCT7MmUlFW+u0
NKp87mmQcG3/yXfbZADkAo+9F3jtXAgIxIq44RlJG5zmDt7Xd3l6ZoMajZPsMyd+
Nuw8my6C6zLE4mEm0rOsACpIPEsdyKnr1vURYoOdB6E1fxAJCISz86/p8xAT2n81
m4yb3jzoUCv6T5BcEDA3kT89URf1duAD3jN26OojXS4ttRWSlKOvo6NnGWDoIFAR
C86wIxgHB2/aSwFUT5NUCxLgssFslLkAgrlckCFjG03/FwnGOn2ZSdQif89Waklp
bD9CkfiK0+IItCZQeBji80tdEpUtfn77sbVCU+xRrqxkKH0S+OoiGqOCQy5ilKEj
X8QzT3ocPp2IIMRzz+ImAjncVzjFyhrqycagdORGQp2eQmjykl6qaPC3DUfTIGk8
PBfbuE1bNGClT4CM4S2nTfmzHaKsZ3qzEgNmdMgJrz41tsI9NjYUt7MRJPkUXvDo
5n36TGinbC0tHgqUNa5LrPQEA9VYsj8KQ/gc9JmkI8SDnHcs33Kyync4/ptod4xs
/fw8ljVS9W2R7XC38bEgbGwKsEQWydVlMYOyGulfrFxKTetGxJvd8A9HABapxtGX
`protect END_PROTECTED
