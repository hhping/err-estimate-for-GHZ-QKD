`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01iZlsX08EU1xhjWi8wTBoX8TJT79fa/3hfSyLstXZeKpt4VmGHAys2DoniVlzOC
tXRK1Ajm4ffH+irEnCPuATGhLeKAvZrDWxQIFi5P7+qswTmPVWY9TlTufnPWS3t4
/vSsIxe035Kc6dQjEhprNWWiYK4fegx+NaD6QKghYCfcS98XRDCIhGqpY/uED0H+
pZsN/oGWupQ706EFCwdtoGddcZy+SqcQdQG+0uXJqyjWguCIGcfwep7YOkP4UcXe
7ZK+KJyIEu5v9+42HFziIwB5Qoic5OiBgPrkCURccBRQd84JNZNiQZ5UkvqyPYzS
s6ZcpSHjE0pmoKuopi7zs9I1GeY/RXJZOgUdenoeiMOaWD7hS0U9T0LWNWNwAKnr
z8r+A9MQjU4TNC+u1vTcBi0zaWHP+BUj1vvuIIYY3MWA87tRCnf1oOan6VuhcECk
IMcSzZgXa08WS721zU/5uJGm9y4VlMp9Cs3ztCrx/XpgZQA63TzOytrmQXpuNS/Z
JRGmwWXv4mayjCEJ9s5NkuJrU8RZJ/ihuCSVIw9P1y5LSvRJESdydG6W5A+g9esj
SrY4rNwWJEpnmSUMYHiX40CB0b8KO0AxqHUFDDS3810kRxKXufmUvxvs+e+echgF
atyboZfE8pYXyOGJgjUJMAZrPqfWiq2SrvvAakUdNhW+BKUIxnUN6T2kK/K6ASkQ
WjFgfxFhU+tlKLEZBoP779dEfeIfdzUv6WWy1nqq1HXbp16cV5T+YXv+xv5BFIKY
4SVtyeVmyHmfLf4voEoBJXx48+lrpHxUEfZXYvlw3moQ6EVlC+ealOV/scJFclXn
cb8ngGMzuq/bjEbRxQrC/3Jz1rG8mTMD4F/CvnFbI4suVMFUen1IYQbyZmiiq8Xu
PTIIFYmUWkWNIwngHlq1wPaFljXZY9RlJvNojo9IWXA89Yn2Mwpb/S4EFPs5pJAn
CuDahhbbSXazEi0UWk219vFAsP9cK/xXQqgT61vZy+wsayzBxMEQYvJS8/nORk6g
M0cuiaUKobrUifTw7mWcvWPayYhEAXAKesgi9M39AcqM06UOQQF3VApCGeIDEX0C
W09ukrpkoc7hPtt8mGInmeX3Tyta5TjVRQcLhy+J7Cl0BAQsYiTE71jVGCpIMNqs
kaE3cWWwmuBZkW5ElWcBC+TCD8ejg8z9mdQW6qCJm82m+QLY5VND0Tl7Bt0bDjnQ
IENVFJveHMEDL1oZ3O8suj7ua8r3XQn4CJqoTXbwkuVRgYUy95T8XjpWf8KScqMT
tNbiTugTrdA7WoBgPz3qYxPH3EEekl+ZR/KXvKjCSp08hFZ1dqDTfIoaeKgRrxcd
YawlSCSG8sVLuNMulk7rdD5UdQNLQ8DBu/9d4sjuVjDf5I4cY7rOWW3+K8y3BM5m
xsljwHLo/U6tVEV0QAtxRNL9G4DshVav8Kq5CDJjJd/CrzJbtGqnhPKzjuFoeyQY
yraZOA5Yhoff4rz7ASAGF2xJsBHTlId62LBouiM3HlRSh5uxan40ZXyN/A5fS4wl
HKv4RcUkhag/uHoG1rQge8xieUs1HzlAqf2pr34RHeGIixvZ/3qRjfPAD27aO4+n
9WZVIG9Cn303LL8pRikyFRHwPmr9wnR9jk0xyJWFYGVtq+gaotn75t+6ZQ3YSj5y
/js2XmpJtdbfM8ZtJX9T+YP+CJJS06Hh+VRpQhiH2w9s/bFzVecRlsuSIXN6GEou
szb2UHbeX9/h0XjprXpVLGCfVQNbxy7TNxVYqmTbRhCbb7JeJGS7gNLmp9S/K42w
AX5g8jqiT7YelYnHPxZFk+RfLcl1F4qwtcd6Vtg/boHAVeh3UDnXxC6kMQyZuSo2
4VcNwacni9A9VjMXFOU2HBLIdBJItLgbV3skXQqOor6hvZ3147qRqp0oRRTfywzA
FdUYy0y/y3k/Z9IipMzpTk949i3rmAmNokkGIlniilL5Q8nx/4JHaq09M1fJMBFL
07WPKdxV+oDMQcOmGz5DTfUofGgHlww3vFFp/ibJL9AjjRZTxhzSQLOCGTsN5jfF
vbZTZ/NYyXE2YjVoJOAj0yjXjEL7ItP10M+2d4HPy5Xf7iNMi3TD5HMiCUdRXrzV
SF68OKrCeNcSwc3IyzqsYMmsJGXd1GQoDFjyd39tBgFLpNsDAHWKPcVbZTwmupCw
RG1eIrJ+XsrGAIrz2tj2JpAekDBnm9Sgn6LwuDRdu7Z9cR8RhJrNsUVh0TY3vh9N
RKP0NgnjwhSnnkIOs7neVPV6BEVT+uG1L799ilsu6KFJp3YpLwYXUPpEMDxPJuV9
uV5ZZZdHj1KEnq6fyRRDHSWo2SRYwzV7axesE4IHgBM47RImERuIrN38/kfgb7JD
0C4VYLaA/q9j6lAczQGVqJ1bDqWUZ2eeqdacJae9syQUkw6ouFUuM7hWtxbUjrou
vcnhyuKWF9G9EkMzGAyelAGIK6PlhKll0pe1DcCzGC2pDx91lAPZXwTE43+DLVal
Bijp40eTbIgmImMyA9v6dxMeRr2C2NZvgTykuP/1Rt9beq/xYHcRc500D+GDbz4a
Y7f9ZGGujdk0jclXLZ0ThQf2myAkkLu/+MWQpuFXPlm4OwfpSXaXPowXFG4i/sTn
y00tTiSHeZOU6wjj741Y7KeIfdb/iKFJ3D3UpajpPgma8so/n2YDaCoDntreYWYz
bt3D34xTv0F5baqT2/MoJLNkSH3LM/wClrvJ4CpJ6zLn9JCqhepDYrW42ukyRfrS
3gFcOG90gngnxKRXG9wv4hkrbeHn60YpVmcPtPg1wnoiM6HV5cgh5ZLCwZXPIquP
QCqPoXuEWZCIgXsFHuhBRZCiMwWWW5epR+5nfopRIMjn3QDBugPyv76jzwGiHXBh
UTTK4SgEQO3yoUXmgiO1GFJPswq4Z9nhYdc4Y/4iuaUefvWs0uQc7gnaRK79zm4r
G0wGmWflbW79X+iCo5OX85ZZf/q/w0nA76guWgRWly7BGrpuLB3FlXGB01+Z31d+
vOu3XSZNYTkPI+w/ckzC6gGSLr/GfOEws3qjK3t/bij9cR/MnMTZu9MbRCyrbuyo
WT79zVRoX3vR5PcP7RsBmyR+DghI/0a9NgOEQwcczh07b/9H4zffpHjYEf3707I4
7He3QYNq4INGeSk5N6q1I6ypj1HPUqgSOHhEXNmZq3jQU8kOAPNY4vw7KMjYDHhc
jQc3kCJiJ0EfZU6gOEG0RQmy3tJzpl2tPW4m8th5xUtM+lNLPle9wbndY1J14dRt
QLvaw/+Zz2O2ZtozxbMaR1B4Ani+g2OsuYjS2NdoGh7XWL+arSmhChhJMQ8i6qFx
4mA97q+OxkyJTKHuM6ay/SNcRIfYczl7BnudVIRA5R+wJ2ikIaMr3AMyO1HLRNjb
wxsFTCI41BjtbDve+F816lK/RSBUa9x5dSgdUlQOQ5xCoZYppUwFn/w++OgzF3JS
hq48QVXfD7/3YLhm/Tv03sbkNQ46F5UlKSu8sNRNoMR50PXPaoAyrHsCjgMHaNli
clWdjhdMLoYnD4FsIOPdUkj20c5NfbRweoa21vxO5jb7jxfH9I1O+ZHpdCh3vh4r
btknEuKuklzYqsCMshDHXKD9OdSTFptx0+erC4yneqhfpXC+CF2ZC78qUmg+0hJC
JVhQorR+sJzrV6H2E+SVj4XKZMlTzmBSqJo1fmW/gKNB7skRwf2htwm7yEmghVgt
P+8S5iI2PjBoTcBZwvVhee7aioZ2+k5u6dUQr4m5tOjOqdDXB7XFsKw87hBa+rEI
RO1XH3ScBaySf5GuCpU3WM8Cc0DsGemmvsNNpK0gYAEKaTmj1eC+tjjs3BxIzvUY
StiCv4Xu3KkTBTQ4M1F1CIkowt90YjqW5ySV2K2hcgMfRki3OusCmDm+dtYn/vc1
aQbJdEJtsCtIhRIKdaSohp0mteDwZ1U2kUf4nJ2vk4Q35VMM+DFMl12NSC4FlDnK
XuyuXycFW6QIevMLNWd0NS89Kd4j6Jk0LY1nNE7ubPRHf6XfL5kExZjPXYPe1xlc
cDWdzN6WVgB+402yhTxm7Wk3sNOzDkO/71vtykyhGuH+W14CeCgoUIPyPh4LWRYI
02yMYzAsG+ojt+qTxkCq13sRgUMYDZICo5MwDcv4m++5zlRiVXi+Z1t6arXH0bwh
MGZxAzyveW1pOs6vmWwATNd+7K6XXx/lMA5whbzy1QX45N+QtJCVP0o2nP/eG/uh
+sJ0Tz6QecoGhEXVpcupRNKPlSBSmov7C82ET6MEptQ14GPpP3gZmGxxRc2YVoDC
F72PYghoU4kbZ0MD1xhlVgwPuu49AYhpB3ua25vI5zhIJg3lxW98Kj6Gs/H4NgS/
U9EcJ0pC/kKYKsYcx/yrhzzusQYXGOomzr1yjlKv9lHlCeja9BmWZRfXknh+BTwb
2+F9cd4Hvq3i/ea0f6P72oCQ+iZGOP3rgmWF1nxixzdg2g8WCDgjwVQNU02JCzp1
tjzjuX0EvhPCG4hoXNi4BCRBA2g+Al5s6fBteFpjwC4=
`protect END_PROTECTED
