`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Xxov5xCTWlK7aO56S1xeMAqcbXbpY0gU+8E0QAFGUTnSYxuN4OFIlD4LiOtp8QU
CsV3rbAO6vgohvDM5tc46+d076lAH2k9C4IiegTpnZxeCGoUkwQn+R5olukYRYl9
HcZAkKgCtJvvrqaZM2YRLM+ssOpT3QBSNOpV96WmStldIJM9DJgs/ebeWto9GQsu
1GcSZxgtk4yd6iuj3YUj1UPvVFRRefo6jlWxikeB8fHTQRL3BL7jtzp6RylV6OSp
yGhwq4goR/JFHOvVvrlFgbFDH8oBtbkwZ2MKerdsYBtivkPPDm/wBgUNk9oR18Pu
hw1hUb1ds5Gr8K/dl4yB57RBdBg5HtRCWHOBXUM9DsxZmliR0FnicsTzseQRqAHR
Sv2u3rB++gLMgTSqKODhb7mv5B2QD1FawzGcgAsdyk/Of7Miyxc2VP1R7zmlOd74
qywmU+dP8qN6l6mQeJS2XwqrSeFaEBXV/cb3h75XTLw5tQr68VcYeXHRTEw7lI5T
3fiF6xivwFr0kQvVTULHQ+gn/kUlkxNUoLsjZKVPO90TLAZrEVU9DJrEhKi2fsyf
Pmm8KQXBXSqS4ijAiQE1hsDll0xRNik+KFp51Q7HrtgkHg8LpMPDZngSO+Mtbc5z
4nfdw5Gp2IXE/ftgh4vmPxBtxXskiECXWH2OPe6voKYWxOJ6baJIh2YY0N30RnB3
INje7eX4X/VFGh9ITgKQw5tYgbGF3vlLdzs9qOBNQJOOspXgz3XlLAjxV6aD5zTX
zD4NsU51bQpFyynYxK7ZINpkTZz1448BswYG9SwGVGln4Rmsm6l/yASjWsjxfUAA
5HoJMwIhUzfrzStOXbJ9YTUqznwU4JHLM80ZSVnYCQwj878D5qikrMbIzCI6hWTl
/EpJKIpSom8tNIo/Cf8rtvXgyQZB0A7ILxflh1mxY8E4ZTS2vAAAuq6RjLHsa5vH
bK4IIVuuS9f5HXK4y05ogFEvFUtAQd4BIcbkV9QgHIsmeoQJHFj62fZOWX56gJGd
07GyKRB2nT0akibezwsAz+cQqGaJYCW/mAwWkZBZUXRVFzKGFvHgEZzQ/ZCxlgOb
GvUrCeqO0fHygXXyj0IN2m3+vnhh/9nX3Jf79gTCg1WXHy06CiXNh/N93GcScwgK
ELRKJLsJpy41zOXWw1c7i9m30168F+K341kTB3paNTijESqzdbWIgZZlxp0bWP2c
bfye0gbW11ZTgSbaRN9WLLQJ5RpfJvQCG1DbA2FtMYXWh2OnVGLQ2uZjNtDBnEiB
CtIDrIWcSbnZiW1d/wxxAc91WpxJOBAqcsAyN76uWGDhtYTmnnYh+lJxmIrIxUQY
0GeA+H1RVVi/wW/Z2vML/Sm23GRpvLdB8g3O13D5BjSZ2YiBPlL0b3UQ+woUVVEB
HhSBB59PxbeEA1D9vpy18cTQ5ftqLZnTWKqmjnZqVIE=
`protect END_PROTECTED
