`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaWIO0a/OAYldcQr7zaWMWZH+7iNLwST03x+1bqo7aSam81s7LfPQYLpGMBKMumb
oxJcyBx+LsMDkeA7ZG31wAAt+OFr3o7A5+J1B2fmPG5aqf90WuTsGHJ8mhY9ijeS
UNAOHtUf171i9jN63X8O1/f87I3Q3fAidsPaAyR0IX5NnjSDprHbKvtW/7LwG4fx
fxR3O0Xwg49b5MRKxT7w6AgcsqbY5odAJ8xUNaQCzNjJeuWxjYhMkZvh21+SulmU
mEo/nBnwQtWgXjEN6sFX1hd4CyY3mJgnYuiz9dGVl3SRxUBZLLc6o5az9LqPulQp
+1E4prJbHub7MYwP4MAzHAi7TO+WLOXmllLrx9U5GLihiKEdsLnzWJkGuUNVP1EH
WLy2Qu9Xlap5KpXNnsYgqMShU0s8JHe9gpjvWClF1FLPwWZmr32hestzlZxBFlKi
IOaElYlzgKTIBemhjOW5Rc8qkQRPjOWnlf26Ejv9yWUfxeW6xnNJVvaXzaCdstF7
dERPF9BjCSEYuhgoRG7nLGGcgBP2w/o61D0cWLvvtJN0A5QdY11fbVeW+kSS3QDz
E5ENmiKmw1R+cS4KxPBXS/UROwe20AI2yqgmeY9Gp04sk70IT/KQ/LbAKusIybg+
/1cuPiTay/6NGy1usHgFFD/lTJLCbA7pA5hN3t5kANL6ulv+ofnsUyK0CpBfija1
aYrTr4oilAPiijVFAimrpEQNfreKejM9RCYTQcviB/acCufmQaf1Xs67yAU3gPzH
RA9PDHXMA+w1S6YSTRxvp+lnMuwT+bTflIfS6POQxDejZuWnc8gC8UXC2Aryn6vm
qvy6PwEsrD2dcTA6Ot5XLgHDvtvahJh+yqtoyhHwrIhBXXJ3oV30fzMkS6+z/+wQ
bxQg/rH4gy1zjaGNRdg9PHIBH9GOMpimosrhmi5O0H/lyPStjmULeVhvhya5mxw4
IhHiZGaS0qZtNoi2X0GHeOt0U4dtSvB5mcVNlz1w6v8/9PUvoCKimSSOeZwYnUJs
C4nN1FpSBLoU9sWFelp+nFJsNjmFb3gIQdWtItAdBMNG/upspdxPygA42xvqryps
ZPor7zJRkj2N6XRJDzoX1vK6JVewMxj14oqVGBMu79IBEUIMGlgB5HJPmtPNAOHA
2hcIrW/+BAYFklBfO4rcXV9CcKY7dFIEuJFaxmSMQ5PLmkbx1xP7ZnImZG+SQY+0
Yt1a2HQn0LWZDa2+jf8jbhQAhViAvcxft5lQGj6qYA9Qjl1tr0Rtgja+yZ/ioBhm
MuezxuwlIR/RsyK/pr8gk5gm+aZIiZTCXLZYH6zuR5m/EOogfjzg0VEkJAlcav6K
DS784UrtzTu4GNI99qlBN10jegGTqCyuB53j4GKdkoAe7gKP9qrpLBoGtYwHokKs
IZ1b62HJw/dE9bip+4KitP0ynZPBkYz1KRPuWL+uwmafZRyS4ocd8VWbwkkLlQkX
9XAofVOc0pYxXq1a+3hQN4CYBQjKt2goAJ2DIfTe2GlN1dVfAkKbYEUYIbBJE9O5
0gtc0/LtBXJLLeHJblxXk/cAbBMjiWcQC3EAYoCkxo/4tivgTvmAA5n53hj+HHcX
c6EpcuFn5sWvn5+xn74ZlBNzzjhO1+IsbWtjSlQfS5pAxTOjHcm2RaWc4qwDW1Tk
qyH98FbgIC4pwlME5zbZ2to2EKrtUJa9S5ErUSw4621rj9/wejpwuXjIBlXaJqNT
pYEj/binVHzYarFtn8Fog7j6NbUJqHgRFXjM2UIPbjQiZSbQLTQQE39yj8JYVWVB
JL/qlMqErgC67pXBqWHpNwh1o2B3wPBrLZJDwhPfsmElsnsP452+UHT+nnooQa5c
I8xTYYW8KQ6cZtba5C6Yh1OMxkxdOXVUrlS5KiPWpovqOKSNo4Eog1uM5qhU3oH1
7IZg5nT1+JUDSvQDTrW5QXFyCn8dqpT+4vfNU61O4SlxYROToNgxMcpC/STAb3Ur
JJTd0q75kwftuXQrK8/nSmMhIupEXu8tJJ8f4uNPUk0uGhYQ3wGh6/QdI1LxwVYa
g2sW1vnDOtyAeKQe9wDDrCVSTTgMBeAFj2dEa8fnck1y2jXZoOB8HK6WLWINC+ng
zKqQVeJ12n5Ny3B7nBJGjEH/UNOxWxTE3Vl0IpeEypq9HFzOxKxLF2+3HweH78w+
I3xEppJzg5yJpZNNd3dvCBAK/g8zk2uOx6gSdJaLUUO+qqtrF0DyvKR57xlD3AhN
ToAL9kSe+FCTWFrPELLhF1DL/H74PVMKCD2WTZ5ePhD4QInPgNo1gnX0K4lAK4Oc
MdG9KTyQam/XA+g63jEim2Z0hFw7nCYE3zNOVdk1CNjmI7YMlXpyj+GQvVtDg0MK
tJrKK/VH0xLuVaz/0x0jgExfK9Z28y3nq0upijTCvDD5HMS5gzeVp24ksfiRQ6Bv
nrcMR1ctfMPC5V6uV+9koSqpEI9SPc6f0rufwANOOIxN3rlyRf1QFvsXchNCZghf
aNPMt9tfr9kZ63sh2TYOQb1CGxI629Stz3CyMCE9O+QhWba/T9RI4TGy8/eyQkIj
ndPlh+mt8aHXa5RH0Qi7tZ5M4chwd8IDP/mgoFcrD59/CrYnqO7sZS7DMeE8pSY6
HSWk7iMYEBWacq5PGfF8golocV0dcwiUZWiuvunP/6PskYHTfriUJ314YaRPZBHT
sFB+xoYEHHSTCj4YCgtrJB2vhAUrJ1l3oFZvhI9WfFThea25aFFOfGaIuBk/2qez
Co7sagQClb5dgY/FMLxyM3xSpDbKFj6TEcZQrrbp09Rw0b/zYf1J8Gf0E9xhRolc
YN0prFKYw5Eru2Q4VdqzyLq+O7xcmB6iVh5S25IwraTo3OALt7Q01UpzUGqsYtt4
u8lTzz5l8PVCL3gqzUklTH3OhfJOMbVbzou3FPDSReWI8OoenFblIGC0+Jku4bd/
4KtW6hbuA9eOwdkWDP9pmFVEJ0BiEZZkW5owTUTFtapSNh+/EBz22JnnQSl/HPj8
Te4frcoFZ9PRepOqIqJ2UU7DOU3+OvEDUHEtHZo/440XgDQwwHBaRpt1d6kDI3c5
Uu+crQ55yBIcYk8rdWCCNbioNA/+cp4m/WeiJhJiKg2F+nURtacnOCQkStZN6MM+
N2lovoWx6+4venRh3t3fhYfWUGUyya28tI52xEhokpwl4ohSO5cPHEWuRmcwDImv
88VMkrp28zOAQrbilHhqSyiNI4Bdpum9wX6w5Cy9rWymHQvUZSEOKFhQNWUf2w1Q
LrKHqjWVe0w1/+rRSGU5NJAB9rDJj3TE9zBcOn+8ThkP3WsBdhFHDoqwWDaZJxQ+
xXKN+xarkVaVPogkaLIZGf9CcMZXPrW8whThBz7ki/b92zU7uCS2szMIfkS6scwr
UXX2rPDSMiU4JM4C8SZqd5bxCiUhcJRbe/To3x2KjL4tSrcs/jX60DgMQO82uUqN
wLLgwpmTDl3rtbLAatRe3A+hswoMlhsCvpN/elpTommBf6TkmTVW5SNRTJjBC6WV
DmMPdeae7e1xwsbeMQWJoO8XsbqJ4KJY2R4MIuGfP5e3/1SvD2YqR1nngh38uBet
TkkEB3EkxHT+xaj7QQd8lmNNg2MOWwV5nmsxyxWbFaJ+MHtHVQHoEewbxy6rz0OV
zR4Thi73l43dhsUE1WpWYYRL1rFn6olqilN8Y6kfa+YjMjk6IgqYva/hx0ROfLdE
GgxRjMEgVWiRPDxaZCsLo/opF4F3yO9qDeDziVwBkkkkz+CAtB7SBp8KlMH1kwD0
SVL2ufljP7cj+o+n164NgcZXXKNBC7Y9tfrQeqNXJX6w0ZcwbK9uTtT+o4NfAPKc
kyfQsz7j7jQkoN23EfFlaNhnwJqjCuge8Al1gF3DMCh1Uy2Lde7xvtZBPQCNKDoE
vOygvmK0c6QJU/srTWmlhQYWfyumdGtgOl82EeYOQq0zMGwD+N+GOpImOZMxwRYW
JeExvAplILB8XUP7VTujhFOs87sDbPfk7s3REWE8HY3cG2Pdx9VHr4s+f1u2SJaf
x845glN96ANKG1QeVO2kagrQcQSQ6eORtmMrFtYMfzaI2XVAqHZRbQLy9Xl26GT/
h1sOnC7WCzrZCan3By5rPnonZNYzEQGs6vLLmZfShxAMSSQO7JhVc4o9Z404+ckD
RfhhBAvuwqYbVTHWDaX4BEHPBCFRgytkLoXSmASZOsfgPiNmbRXRko2DqOQdVxP8
v2Z0A15G2A4xg9tVyHGrxo8fGaw9rRX8qpXLJGmCPToHBNzcDwKzy2SCKukCfi41
Z+DhEXlaKxWx1yCdOxNokditltWUWEk/QZ+zyIj30SuNaIaghglxtOANpv/Zvv7y
p78rTeQGCVLZPW0qBEvUfJpsslY+eEvXblBGenVjfk0KNbZ3fwCBJFOzCKUtQOIX
pir2cJXFPvNh3G93Lg4BjDcXyWS8yyulH5kbgt6CN8VeSPNQNu1lkeh1aJyfG3AB
FKHtE7L+GsYCnGy955slsJDsuTdu5qTLJj4Utc8JuKnGBxfgwS+38fPcyBtPAbZJ
rTfrVZ/aaTi8EmHw+OjDb+n5aPkDAW6zvIodNePDEjYNEPhU3NNhsPvx9aOeqaUB
FZInr91n00LMS96tj2se67peNagAcuUrN3TOolN8YgunWMBFsy1uEiiwdaVRTV1A
0KISK0hlZr37jofiSTaKyRcrLGVd/XXuD6p6UCXo06AY7nPRjr+GsCw+0dmzBFg7
EJVl0DaCMrEBNWXSjhE8u2bo0vXaZpXG9DXxjkyO/MeeV0tiycs8z/q33wL7adVN
8QjO0rq9e51bVd6pP8b12vuKkthT8QY578ZahSLnGrmoTNlKW4YQE9tpw0wpTRC+
JdtWBkCvE/6pBApddFSsnx+YrQ3gRKg0ARNOL4NAXD9ERnwNBGSEB10M80JIdkv+
awSwZs5xjhSDF5VdoutZpUOxIOSSnMHCFzy7AYdCadAVPpBkSw0SweMgfd0mReVD
pYgSiBa8GDYb2acvnGkgelnCE6MC3gbLIgUEDS+Ivb/KEOV12L5rfAxtYJY281ZT
jlLBL7Zyw3AasSDmSh6LJ2F86fEDGnBqojBJ4tXL2MkWeVJwl1ANNirVxy/FzFIf
PnP1/Eib2ZL9lr26skfBwoeBD6FCKp5RAyBmMbi2rVMbBkjxEp30TOmmdC2Cluxu
Ry3B2SLCyVcs14+hVo61arXXXwaYdrp85tGehv8CDXVj8xykTcVGrPq5qF3P7vSN
HWLCoa/Hp2q30exSSPYccPGqi22BRfHdADCxKpMIdqY1Bg8CO6nhyghwLe/u18G9
dY0Ldn7eBC2GDpTQl689FtDQ2ogo4grKxhnvLmp01CsqC8oot1sA1UapdKqIA5a8
Jl4VdLV/OA7xtF15gm+dI9bJijM2vbSb73Uzric3CQuwvFW/oS1rd8fBKMO4C/JP
rngZC6xNJmzKunldllMxh1upYI+O91hmsMntbvJg8uqSlOWgHKvqmxwEqi5pmq0Y
/qw4ii4NyThzHIJxLmAE2q0bIBb7u7roXp9Pn2PXP8LqDgePbSf9tk7AD0xD1lxz
9iIGpgQ54sqwzONxb/7tCx3zGJmvqVXQ0bpEG8o5vpEjawIG72QuCA+967P2/aGx
j+aPfPGFpxc6sNWvJ6tjJCd7HI6rtaOIF4wkXkwRZ3gS22cMicYoVeeoZLU7yRJ9
24E44baIAX3MXu666VfMc74OgJ6XdNi0YRdGQvUUFNevFdZ0xoPJtepCPoOeoqrr
x1ht0vGQiEoMJRRwd6Pr676TUMpN2PwLsnHLydm1wsuevTl0cC2LtV47FgrPbT4M
QkQlC/i1Fp8i4iyK5VxVK7y8dJzgFcQiF52QPXwO/Onbs8zKgOXCJ9Xo5rCWZD2U
J7GNtAd/khU8ZLLyNh1MUSm+l5JXOWsxWW/FnhNED7gcXe0qx40/gRAR8/j0/zsH
SkFHF64TxiRR0bBOK3z0CWeEctkTIbRXB7V+l0cOjvY1CvYfG6catQlK9y72Gpju
ezlS1bM5SQXxCwinyT/TMJmWGpMphK+V31Cfaspw4bfOeZldJQCHqMyJmwT8UZfC
/sV6UjXh7HS/Gg5edBKZRs6QuW0RicBJNa+S5b4CzENgqFdK22rieUygNR/TGd4A
BWQpZANpBmJ2h7L8TGYdxUdGmIRK3/NCDp6npFZatnZHXBO/bJMAMRAJvOeJDKF9
agld94+fRGA+hnPJxNzBouvksDrCR++DHCkyuFhEc728TVsQR9j7Sr7hu4/JlpkM
8UxEs7YEbAtLKIbEz1EmsFRdJ9K4ichjrDWdQaknIVA/kzncqX6wsvzhOGbUooHZ
7pqsYpcimnGZNcXkC9TBe/xruWnCStTQQC8+YAJyC/HEwKtwLLiv3vNOjUZKHFXd
X/lp8udSDKRZ80hENSxsZbDimSiRsUWqQjFnE6jiZesYP4BTYBtM4OLn6VHrJqG9
OXHbR4YezqY9n5Ry28q5qSox1ansmEAQ6Q9NgFsWp1TosYyfuUr1ckTTKJkPp40L
HEwxH/gdhWQ8ZP08RCMuuYTdbnrueAheGvc++hPQlQDIysiwx1LnqrlORHRyc3kA
q4GOmGbU+lMoVDcpWoWg0IeqfUPoGfts0Z6q7rg2ZdkOwL2PsQ1Vu2y2yGXvjnX7
W3MIPAWia3r2zDKvJSuIVkuPcauP87p28LT1aD54NP3tg/4uXH4unEuYRrX0IDGL
RFnYy3IQwLX1Dvi3psvgMH1Lq/eq2+6mlmFgwh7ddKF4eNYWBEk5iQ2MsMfut4nw
NJxlwH//POjHPCDr5U24OU+zSXHcQ8kJJu07p2kjk5z0fvrh7aRR6x7ILiD2WzEl
C/FJGSceqJYMWgL/ivMF+u2JJNzqF3HXsyql1K1AVRcvTytNhdWNMhdFOTWr9y62
Oaod5SS11DbYEi4oafN3wIF2xTrs6U+O7kyoYZFfu5mHVovRcPXFsxjtgIfSEdkb
brl+9lbWzNGSHgMRP6RFc+65NGru020ulBC2Gv6H8lwo4JLI09zxvaG8NtdDPYdr
5O2HDMd7lfaUzCK0Cmj9t13eApK1+KrWiB3O3ZIHRPLgGQRGk4U5TMoOjhjylerx
D18A86jriwuZF9IhVph3PwTHaUYBHrs7rb8dtqs9zF6DZvg5jyHDnXPzjSeFurYs
X0APU4GAC/2DR5XaVLrLKzuApM9WigvH+nC5SsFOfZafvetA6vnSQFM/dIhFALrR
7Y2DAsk5rzuiu5xOyi1E9AWlhrZ9XrdzTkAKyjBXbcZ1yid/lc9oewElKfGCpP98
ORBeSTNgCI5hEfzzo7XR4O/l2CUHe44YLBnUHUTNX6GwrIBWqs7BYoGJKMUQbxBk
zVUVzZXnWAxg+U3lBVx1kBNfyTZ79IPosPPAnoUbDx+NZUZ0ApvxCrTs3skLEVab
cBFP2F9es5wG5KcIfJ1sI6piKe7HCgIkfdvNIS+ATNzi9GQ3yBEty/MIC1aq0aod
Z+AgqDd/VDmwX/bjlMWmvrRtwFotI4DaAFGm1EYWlCkF6DH8FABQj9iWTBBwb3wm
AVN4mKULfzdhxdPlQOf5EVzHYZwMDKpJ+bctXyK0/wUYx56QThzEtaz4HWYnRGa6
typFljmEXzX4l5Q/9ZIfAGbZGYWg41OEr4sczc5bngUJE38OnWD8pmqPDVQcLAEc
XowO4w8JdACXNxzXkExsWaUsbnTqNi9KFLbGpKSyI0LY7cDmlbHKvzTqYCxlhhjx
PNe7VFQof+Q8AvA7KYvPuHG06qeitdW6lK8nKf0VjV1R61y/hlbgOSb7KKe4rxmu
ubHkykY1Lz1eceIMopdqyt63wgBNvMTh40DXMofO2yDkHTUJ/XtLegMkXHgxJw12
grEgMu6zrkX/46ZaV68TyP/CTBgG4zvUZPrp6HtZda5MiFloAYKByBasftLGO6Z3
S9+CTAaqD5wuiSgQo67HirX+qxaSpRZ+Foco1ELRIy0p7MQLbToJFtkhWsJ0Ls2+
AUKLoH+0swjxyhZnm0sxaEMtavSNO3KlbH2Vbv4cuM26DcRWoJ643v8sdeTxjYfi
SIcCv/mvHqTr2XOCb7qOw7HGh9Q3xfsLDerYwkEPlOHkUonbF+REAiPSIG/M68Qr
d7UPlaiNzm70BgBVbiYksIugD7t4dxu3fzqlema9UbPvuD4DUPmj23Hb+YZqo+S3
zCe1ezDfYQK0wdmgDK5aXXR9ONdY2leADVk8fBh37TyHQ9d+coKJ6bazKJ5MOF6H
b+G4STuFtg6eSKBMr6PtJxdDbGLMYkj3rGvcXJZJVAVbxQG3uS/o069V11BBKYH2
2w14vElwzebjfUjXcNmKAot1Dbgp3RFbXAWwrKjuC3Az6g1j8Zif4I8t9jp3oKyy
ogeIogriZlDqgSc4snFyUbl0vJqo/NES4qxk405pKM9brTqzlk4XTV268Zo3Cp4F
XxLbNb/AVgYoVhs9j6E5EtiAAANJBn4Xoj6e06/4ZV4D0/poF5JQYcL0WhcQ081V
dJlCCtGpd6boz0FRnmV8/hyAgJ8+2o+HJluTPQB5Vs6j6rdXkpJaFYlO/x3OyagI
Um9zWfhhosOVjp9CwIW8X0ZGZfjHs5mobyHECuYhWXdE3jrbWAdGt/k5h7BlF77K
QNF8Xh4MpZUzHy1U727w3+S+6FBs4ObC2ZqOLbhzjR/FrsETLJu1J1fyhjjcl9Qh
lyvruvfVVVGlPWKWWj2ngs+X6o4czTBndVYE2EwnwhtMG6roBFmZkDXIpjYU2t+W
R9qlIZ5K3wZ1Vswly6vhYKMZAX2BKAQxyQ0aJbqOypX8avUfTieb77dtj1gmNGYf
2VO3sPvdSJ9lEZyCR3oBosqwUzBNIUNyPIAheSoLGysgENQEOSQVG0e/RWkRWs2S
PZz89m4eLKi/515ukcfEwnIREVTQoJv/NHTRxwPdWgDLbp3GRvJ5+dnoCtIopta8
jY4t6LDeRX9gSgEVbuTvW92fXTr2bIhAkgrxs3QjTr3yOX9NZO9Cg+r3f4mo2VE/
N+xBBiP1MyXbHk/4fTDZpWAYKJBe4+UF1IJqjZeGkRxRkv2fiudxj8actWZzHi/K
vuRGRupkJJFtelFLz39ewFrCFhLLX0eREl/hKWxfjxsFmBhbxPb+Phd+05XZHTxD
VzraokYjKNvaj9bv/KA9+CENu8AhdN5m/xsjtqV/iszKmLjTdX4d9Mdi7kbLiHh9
bVoNmJt2nmuq2BzjNUfCDSgWjLOQ5rKh/oaWQwKOIoBr2EOZU2INIUhDTRueU5HR
K9FInIB7pl4lWOBDFoZaCfXr3XUYmJR/YxAdTZfscYSOg2e2fMDsRX9f/YE2pUgG
BqfCthIPnrCwm5WwzQgKQw1+tV5N4aD5iZtI8Kdw8cg3POeclGRdlrHs8hHsAF26
iXcoFVlONqteLJn543zBhk5xWNwr8TSA3dIhTKKmJ2rwEEC47DyuqpaYF3hWo6Dx
b6P6NmXuUyMgzWIr93PA6kuhFXMP2ERBkzqygejNgkkfVe0bjmjtRt2lZ53sFbHj
qQRdG8rtdMQ9X/fdO/JdCak5CroAzwhEScfeBYZe5oit92TOhhfuFpkX60f4BIAF
sqlQKJIbDcKJSL9X0azhKIdU2+yeUAXU7seINXSaApHkLwZwFKvP8vSX5P097Zci
uKBImPPNnBLIdQM483liLdy5FPIHWM7DbHBsZwEIYGFDWmmxo3ND1avTSNkowiof
ETC60lW0PPO4SkdVNKW3X4Gqx5jw08Z18MrsZzzMgIa/qBg+wjgxPohyaGJGv3lb
HWkmiBClTFQ/FbNcIu343uI/6ZznHF3v52QdShFUwbHoWq2dJShRM38UGNcPWbPK
46qWxg0uo8EfdVNOPQqHmo9Jb15rUNCRAz+oyCM27KlJuuuMcQx3LpG4YvpAtaUg
bTtSEOn9O4/Myko2diOZp19H9HdTCe9WsgZdOEjeplPFuGzKumaYTj7YGXTeS0tE
DEmtB09xeTmFie061+/JRsGv2btI8SKv2wbryjkIjKYo1y9fqTP1tFI5ydrmngDo
rsFRwfUUCgd/mBc9rFyxqXSt6jLqoSG0HSscdZlSo21CzRD58Pa7ilDJl5uMI7VK
QPozOvsx2hVnMmIoK0pC7eb6XYwPQA1igP6SbcT7hKWwNRkhUhJbwVzMSWAHSqod
ve8hhF2idu5cwLJPa8vszOuhpmraGhmZ2nVdqZJVfPqvXMO7IPapIRqp0Dat3FJT
Moiym+9yiUp+kSmNT7PPHG1gpu4Up8QvIIpPkLnLU9BNYgBG39hIsLdkzr/PtZi5
Aqki3HgDqTzKuIE1jgFOrBitJaMnm8g6/MYgXW5Xt0QNmbbSzzpdATnLb/VTpnRY
vD6GzU4GiSy0Vsqcpkw202S9wMoDRQEKGjyK854wSJ/OnqzNgIbsYNkl/yrVRv4b
k150wJ0qDdvjNlDs2R5dvE94R31Yienkxrs9BAO9ld97y8NFjCzoNiEUY70HYOZc
ZWoXPZM3aDC9Oj4YFT+cPuPxMiu4vmw5V/A7Uye/S0eS9taIptTPFKkWhlJtBF7a
ddgsyTyl+x0gcFXEYPB/CfJ/1YgAYEGLL5eTqQpmIDoQn4FnV5ke9UExnWK40PTh
DL+p07yD8nBtAzD9fFWe+8U6UtixP1t/4XFZA/JSKA9QhTxtVQo+2lAgJ1lnK2GL
T93gcBICye1k+fQvsTzGVHmG60O0WBKK36tPKYtcGR0K30tYd5ScAeycUEYzc+BH
E9QDV0qkME3DTq/zUlLQYGTOCL8Hro9yC/M9f4ijub16OfCyeZuC29OvQ5lUhJms
FAzPT0bjhoTQ1gpvs91zX60XCwSuwHd/g0RIUo8cAqEj4CyLkA9i5BQf/puvZ4uw
VWamCNW1e9ygAAc9fWC9/ept70v4mmxvrBCWM3u83BA17/4buLHx1LX5VuXLBVPH
uUq/L5B8Xp8zinvg7xhwjcQt9rjFx3kn6R6C34quy205mb1Osn0yGmnqh5F8u350
sWULixTYNDtYXqkNiHomZ+EZBI7vsq0P7yhxLXkgn9TX7y+QcoJTorpiqbbPsX1J
MyJKaSioOJwcm2f8dyIPe93U2nIR+AUY3O8WtP+0FIRox3ZfvJXMlI2wwzOklEvC
MKXUP7NfH6kKIl8E6e//Szm/XVJBW/g8+gdfvmlCzz5iKxMAlzuddaBSX/zHLaR3
BdZIPgUVJPpHYr01t/E+/GCoE+krnQ/TVYeBoYWKG4ZEsVgzVplNRIVXPsKMj6tR
7osH4OazIFQmpEHAaHwTjlojlu5pSWtEyZkV6VO5GP+eJ8FFqvCEu0L5p/LAujo6
x3oreOGjAYqRl/sXOwlif2oE829F3IVrLL6wfZ3CkHHTO2dlqH3u5dpUZx643V/F
tzvZ0lBQkkv4TEbaRBhzC6YaECGYB3PU6oJfRyaRpZOiIKpQ8nD+RNeOdQsk8B98
zA/2UBGzEAkY7jtneQ7XVGC6YDxpet/CARn7pOsV2/Nqq30vwN5yfblx2kc4CZVA
90T0rJz5o7jPrWcDtH/AES6iI1OJi17e8rRWf6cBzSpONUFbb7Vr3kyrLthTqJKV
1wKuHFXTS7aZAaWj+BSnaOQCkFauw1XzwNm92hD0P2bA6N3QWMCnbhW/nSVTENg+
S3z0IuSOaw6GRhC7zZTcs+Uwf7FhG2RRnUtjeasT83e2YpWiKF0Q5333iEWADEhV
HPLSvabOw2y0U/myQQ9z8RrZ8i6g9Xwx2iELb4SDQL/MW3hcdk6Bwq8EBJ8e6D6w
JYmAWnHgCv+wq6dOXx06DzpWyTRAENYCwP6SdGVM4jXmQqwo7FjI98H0NLU2Dzi3
vhWmWqqQ73qwguXQVW99BhuxE3mtjJGbIqSN5KDLD+dMbC8QH0jev2u3kITO6dJu
dGDGuCQjxyOhxcK0lNAb6QEWj+ZgPXHkxnupD3IRO1WssePkO2QuqfV0JRh03uIJ
AEoKd6dlLr4Amtqn0Bzbvx9g1CgN990Muv15PuT3Z6bRWXGxHGmW5mXhgsH6pvax
wgDDaUrZfcaQfnLd34AiY20vEinCRyDaOfBqGc9e3ysnpdfimIiH9R3A0nciSDOw
cMS+XPmaleSDGND8guhgxfSmNhmojpMsdfHjez5FB0YcE9OtBefuXXHt3Amasnmg
rqXlXbtIznIov3+5B/68bXC5bm6Sv4I72pRnDfzk8F7E2A9jM6/b5wE/1WpfsE7C
Yz7OKE+lVFABAPC9XpvWLvPpqQiMMBy7GJyogHMo1oPw+FHC8+wRdwf5uRaBShCU
FUT5AC34FTYmf5Uqj+xTZ8jbv2/xYY2VdZ/C1tuNTa57IjlFd9+IxEkN3Dqm1wd1
f7dieKl71LGucW2uelIU1GvfTto1I2Dy3Sifw/gQtvf49oUQbFrmtolf6sNtVfBH
NZsV8t7taSMAOrk1in5bWuv7Nu1+7xky9kJc6NcrziVUcIs2wF1NZ5P9AfndSyyh
3vU/zve0qk7mS9SfCmriUnACVYWyHfXNYPS2QMDAKyGQVXIPUoBWip+0bGEzo+jp
J21mKRPkHOuf5U0jyMyfPxSetFGUgAhCYnSNvd/sjtUi2G6EcTu6xeX5vJtvtyAU
n9J9rKYF+35o+bvVwL4bD53agCLh1+EkJ8UJplSlW31rc2jVx7RRIP/9yRBcTXWA
LLrDV3os75b+Dw6S+exH1ku6kmg7dhfmeEHAO6dc9KP55do7jgGGCeNlZ9JAVojr
TUraEIq+xoPbXUskXA9pMEmwoIhdy+O2QBl2lbQ7Cc872mZz+1XfqV0qYotPYsUj
d9Ru+ylmh8JZ4icfmEchXh1aqqo5VReuU+lR1AK7uWCxTYI39ejv+Hi9ENUMO8IV
c7UncnooRpcvOf8nOpao/AsvcqCM255iX0S/XobK4SlcVm7/B7WU1HalmfDiF7DL
MwaD6RYvDXX4Ygp8DVFRrpe3zDOut8vbsPKTIS7kj7e3wgdbQpk2fB1O5hqmblAu
4lH3mv2uZIW/wovm8dj/wMz7iz58DE5Cz1bnDMuZIL4i0nMGGkiPrOvgI7Hkvpgx
zlgSqtUajCbgMUDcJZb9lnZSZM7eQu1/0su+Zr+mFLcTvEjzKRC1mZV6PIDRvL2Y
/SrBNE5WpSzsC2+xQUzAWFuszKCnpFVqN7zXCazMgrO4Dbe7+WnaRSr6qUfD7R3H
PjuVDTO8FKRliIqw5hYH36vlaI3sxLbI/zn65GFwdrz0ltj2Yd6OZdJ3YRLbcTmO
xHkRB14SThBD+8RxQAqiOqcrI+aDjQbdw4+qPXDcVY34boonk0P+g8Ja+7tDqxqz
A7ievNX7NdD0XkPMhiZHeEsCvEzTG7ilNUOKwZrgK5svPHnzFfdrBY/sCEQqPlNz
ZwSz09RRFyyNTUQWQVKcT0NmAxOTYlZ3a996GpWK0bwscQFyjRtbYGt95jHspRc1
gpOGhM+DovKHXWPE/5BWZDCashOuty/PxqLvLbuRfNCZ+bP3nAWN0oqvrh7uexBk
hTgvXWNdvVd4CrrAgL0PpMIGcM5ALAIQ6sEoHba1h4DkwPxSfVN9mjHOeFf+mzuu
b5WgiiusZ2fx+7JilDom8sNHrkRgeYhxN0eG8mbnkwWO2OsW1TMe6r5Oe1s88H1O
kUjJQ9N6j8XbJ4Gc3mJXTi2WeT2dips5W5m13W6531X3Y5un0YlqBaDQVQtTBMKs
vfelX9nxgkQTMt0MZd6ARBUXZsdn2gw7ufKm5AgdhKrG8vsO6r5bWawnKViveH/M
88nAUmTSj9oWSpgLy+up1yGy15u/TqiHqdJZA1Z/d/AiTqHBcc+81BEmMyORaVge
X/Jh4KiaTZXgr9KQDDwjXTN702MHSxgRkmpYHT0RjySBiPOH4XKgINB1jgAa5tZn
VTkExoXDRmZkIh40UWTkix8e/d8NezxmJ8jQMdxzCwL5wixHu8CeaDsVRHmcCFUb
mdrphmgS7N2XrGr5JQzaGqRLuRMdatbEoD7go+WBfIr6CxL94/znCUAXuoZExT4o
TsAIusZ8fqUoct4ghhNW4YEiiC4+UH3tJEu1g7stqdsDvVNDXFO2/B1t6zWfbAid
xAspaMTRS8RrBCZNcLDKFncW76PtUpjGdIBicQQZ9xyGbBOq/3eymokgt8oJApSg
zOTxxTnOllB7u+B+ZN0FcWPDimr+H6XC4X4wrRmv5jfMEKlIXUZoeDLjmsnCS3Iw
xYj3I8PN0fOR/s8tTtdmMaSIC8bpP/s86Nx2meM5yHSQhtrAqO1ZF5GwOMd60Cth
P72H0w8jpA5nA9I5a+HdCmw30ow6p0LCfEkcHP8AvF5UqN/gmQ/Z4vnmMoo/Tb9b
uMubT3TrK++g+gKAS3wXA+9GvUSPXOta/aHyHUAertjFNTdenMdAIaLwwEPnwZmb
ga/aKaBhVooXHjmLF7b/i1hpESiURiGslEGBBmDfO/vZ81F+EvW2TIYsgRHQ4m+D
/5/pDR2rMp0e6+GiZsBOh2/aAqGrgwb1IA++8Wy43YezE0lfCE7QDAIkDh0CQ/0V
0ean6LfN55R8dRpSkA+7RkTkfL8sDalzAyb8hhcXZMtKttyriFVySsI7TkAxhRQK
UYSE+kRg2aE/SCFADh4Rv5AbrdLu2IyrQq+V9BDGWP12ApiVivWyMClC1YD56RKg
73m84AO3jfMn8c2XEP2zDz6xq7LktwrnTSuexblZrTluCBdAVE3vbLu6mTCA/myj
7o8Y2N4CpNKmO8FcvjX79HzB1n/PzHw5jSIY9Q91vIRCVDj9w77ulF6C5g9Uw82M
J2eM5//BgZQNd45LvepkBbz+SMKAonmrScSdaVDC6jl4rOhrzNyHl7FgSCA8S1Lu
7EetWA+vEhajUEvCi5VEW4HNj1Pj67EaUY2bLHeJwe+KlcUEdesuLK1HfEkOPLnG
3DRDDjYu9eIuadsc2DwnFHZpUeOMS0o6vTLe28GsPuqjNf9ZitxegoZkl0Wx3Msj
PTfGYpbnJmBbjIBdNb/VHbgJkWE5Pj2nvGy00ecUAxIeaqs1NKI/GcBp0PW04bys
DZF2vugpnN4KjWjKtPv95hfP2ck47/LjS2H0hgaPA2HoMM3/QokSOSAE4H+1ozVx
or/YxDkKU73aSlL/pftJLD1xaHucrX1T9RuBNDlltBElkSxFbgHhqrSu9USJBWD0
n0d5/LL2avMo0AGzsU0eHmFAm9vKCaxTLYJs0sld5uZFhYiiCmYwpQ6PdiljA+1B
kVmjn/vmTjO+hF1ZManZcWPL99nvw22d27jhpL1fm/cMfc0Cf0TYBasZ8Rk8kDkC
O9Ei2D5kezKgkOQle14r4m8fSPgbFbZXiFrlL3BV1V7fm9SR/3d/Rl1eQCno4RZp
iHA0jqVbxG0zFotEQAXmQ9nIjepTrbc4UWgkbXlUkcIWEWaxQODWJGt71nWqruTE
oPpnPdnCisAYO9im3fpSY6RT35IkKW75V/AbetoFom8Q/oq0YQQBTqM0HAD3scfy
3lfMdxNSkQU3305zD8oQFfDl0rIrosks+xtiibFuYdbJ+8uXiRLn+bTJlEptoXjG
8NEaPBEm1w/1zLijLecJq3e2Vv0bAkEGs8bNYskmpyfWSeDvvISc8Baa+gjlrhkN
OGn+ezzfw8XKrWDafdnkrB72Bn/hJrFUuAb/wLyyCZnFMjM+9GOej7Nu1Nkgrbdg
88Ou8yphe0Wq/A+vo8QFhEzphZJZF8oqMR7J2ab9bA/wQFd3CU+n2pdkXeM4iM6o
/Y0tNNNFvhN6Ndile4fIMqfzKnb32BSPkwibVVG0qlXxTG2u5Q917urPuBguMK12
nohk1bxkeoIuoxJ47b00x5VvK+GukJt0mt9C8H0V1/ztEe9Js0AvUDNFWIUKbRJB
E1nz/ILMzfywS541u819509/PvU9xw6H/BbJTUZWFu6XnEEL2mMy375B40IfASxG
voua/hlYr56yniqTXPyBANIkbTyOrHgA56b1U26BJpEa80p9We174j2LxnTPkLQ2
fwfWinhZ6vmHjNDTbnChpy7O1GrS/G1u5V6f9s7wf5cPf97QT2anHiKEtDfO3nEO
+QCcn6vf9Q/+zGi6GyjO/3QjByfbGNbFQKLwT4aSP0NfygSAjvizZ6fJrNDpjV9x
v6NA1kYx0AhbnQLPj5xjarWobufnJsN38ZWuW3z4NEjUC/JuTzpZmXtdwhJ9hwcm
iQriClW8UwcAsJgZ3vAu8i0wXHQk+DURsqmUjBbNbXXjzUsFHDYze1Xx1EeA1pkx
JxdmN1/WjzNG2X7YNi6aHzIOgNFVHqpLTh7oGo+2JZeBPNSk4mcNJyH7YdT7pC6E
DkSrheVYO5kPEpp8bomeCjMJK3oeT9c5RtpEjAeS+6ICSOtlBW00DLJvI3k1l1Pd
+JhBzjHG51QO+ZF16rQp3Pea2O72KDVzpZ4qlXTQ5sfVQRuYfnmqh638n8ZM45cN
2BfXiOPHM5eHvLeHd6i9geXKfPuZ0YFxnwySrTncmQYOcA0E2QvunU95nTU+Xja5
qgWA7tBeXIphd3YQt7gYfRbwdRcsvk2tbcwh4aJQ5P6q0N1ooK1xDR49wdgd5TE7
u1admkkJXLxzqWwgrmyU4xvxk7q7jTFDENlLZZKoqjA/aMeY8of9F8LnSGJ2G1MU
xRoYgEBBqVYjdnVo+WsaKBsW5z0jbKdNsBHcrxYgI6M/4it3VZTMNpukUWiMemVt
HG6IHtgGX0nG7+UaxBBG0HbOyI/mgwhdVf2VWBuiiIXmHQlY6oKLpe3aoGb0Lwfj
yOFEhhMapLMLuBE6LsfD+ts5RW59VuoWhYBiRAq1C1dd6VDsXp1KRLgF6ASS+V4D
TQQ5MA4fcwpWUFryJrku7CkFpS7xaR3mWcqj2G9VnRnzpZT/dKIkfr2PA6T2W6Vy
HSrj1i5OOi+Wbd9Jc3gIysuWB/XBk5flH05idjPeQF9/5OzVWPApWjYeFaaJthVQ
ZMF9CqsbGteB5z5EIHXTN338fmBgkJrPrMvp1bOKdTRU6gEdNXLrwZ4dypD9wOUw
KllwoGpAWFRsRPic9MsjzS1XZRqdTb+1Rkjo4YmtBe7NXPo4qnLFQ76OcpGeF+pB
iYNWWo5iHJ6yw1sZo5ixvRuG4NctFr2jLLmFBS0rJVonC+xpV2whkM+XoPCdhKlR
VM8cRAsUDtkGR2/FiHzd7b5GsFb8Z19M7odn3E/dCtLx41cZKGrMd6UU0POsM8p4
6erokhrvyXuDS7nn/oOjwUV+LcccHkQuICuil72Z4v7XOCBqpM8/e0g2vwwD45Km
nd9rxItFHFZJMGxBL94DAZQaS7+sA8fk4UOUNCsP83bbuoanzjjNrFks3uSh0KF9
rQTiamr3wZSzheLWT6IEGp1ZbG5OMTwXyb3mYVIRdBwDcVXnIhfdcJysj1+3bOth
EolcgSByISP9s6vihB1lBlhXkzmMVZSUKjzEHXyzdUSuXzTLcxKuPS4A8Bp407kX
FTY+JZ/XR/4okA1Svb3OPkakcstJnLI01VfUIBNC4+RTJN3ha0O/Honfw173bT7I
VR4DTNh8ozGTfZHkyWU5o/YzdMig9J1mIhXYYLt1LvX4DguBxZXPCJi5RxjPJBtq
RKyuRFOtOgMr/tzckcBrHRwJWsWq1fBeeCkerrvJswZvBzw8nxR63ER6j4F1aezc
AhOdwrmMxFuSsDO+kgt/xvLqEpUd38OMr92x1FsJm9dBU/IbHDQ+xeKofHV5EbTw
FT4/zzj1PsTaZnTV0E4fqkF52DNmp0TpHKpEx6niQiQldCfIpMagExuvyywcFZQq
ZhxN+ZKpB8jkUGQ05FVnBJyBmZFUeD423+INSYfzyzNxywwY4nB9Rh1vmhbi2tf4
yrDjt0sGwj+VIP0+afq7kDS4gTgJjtC9B6cngLSL3+ZQE/IqXAErlDlfS8ciAhV4
B7XMkXpO+LyA77FIWPniHqQwnfoae5dBiTpoBeBEyUjjK/ShcaDVyIKSjUjXng4V
0VuitCpW02hRyFwjyHYx634ax20i+EERGY0qD+jfEwsk1crjHA2i2gz1FSZ4b3/d
6bnNo4OV2vYCN3fVrPUyo3OMKFfumPMCtm2epwhT/RTD1itV5Wwi0QHxwOOYBSx9
aSHny76K2h8iidW94zyoVJk+eqQI3nb998gEkbAwIyOU2eh2691/SN8hfVd1CEO/
zIxWhhVXhEeEFklP9fApByEA+op4nyGg3Pe8Bgjgt8ybRL7gM3Tv1bwOCEQELT6u
X8VnxO6g7EoX0985YzEDLO+C6PVICPcpLh0050ItjcvczOmlHstueXMBWu1Yjxd/
hb8vU4QJJUTSYWLb8XV6ofB6ZxCC3i1qGqEqyFiAtGIEzgrSwnWGyfQ8vYftwlIX
dR/iTumYV81pQQ2q/z7C/fEbrf1ZABBs2D1Dr3vk6N4uLW62FhbHUXPDNvcv/OTI
yfjHBF1BJNUEGZ9SHqrmha8SF7NMYCWsLjQYmNvo/+VR9+oka8kHDWNFw6op+YrB
3XpVlhJ4HLDeMgSDmZ7paVVNfVpM33GMC3AkFK5ofNvVy6BP02pOvK/ucd54YbjK
MMeUAJKqeRQ82TqvHFb+dRfLYr/topzsr4vwRYBB+ogFRW6gBnckRBKYd8BdkmIn
vrLKCuIjuV1fgg91BFbrJXIjLvtdTPvpkxLsf9sCuRWwaJlSFeCW+2WMPWk9IAl6
CijX1N2VKoZfJ1FhJqlNyLrpCyI/ulnmpfvEpchOoFqeeumFDMJ/gtL6AB802TyO
+MxXBYNl+xZS2c+9Z6gDvg7NofmwKYVs6opSOFb38Mtrbwu8JR0ieNAQo17JxmKq
Lexu/yP4v3eWnViXdkCplKQlR48nw6DVPSVvd75AhsObI7Uw77tiH3it9aGK4ZM9
F70iph0wQU7xJB+OtfAmK5r/NB76zsITpLk5exU2jsdAxCIwcAh3lj5qAPjz7E1N
LUa23FNH5JcTDJOHVBmeVwuqdrIIe5D5GqO5/qBy7fjv9TmXJ5tzQVC1sMhO+kMM
MGFEAdEH/gTRAm/o/0x/PXYnip9IVpg+2wxhqRiBg78XhNPEx5RXhiZHLeLHprA8
Je1V5lAYM1ubcgPQ/BF7wVj+McF8c0+qiTNIxOt81d645R3GRVpX6KfVGsDVn121
3gweMDl3MOc3+aR9zny737rAGltg7MRPXZbiDkUROf9qwo3hF4B1LYBrx+wkQgFK
fCSvb5nx0u9Y91U7h+QVUb4MsJpf0CmPyk75TU0cC39rt+6Yp9ClWbXw5vlYmSzk
Mw7YJH4uckDm2p82yzo2ZUOySaGM8BRddQHN2PAqEz8DT1i7hAuSXB2PTTXJPxmG
p2ym2PVYAWAvnrlZhJuD9y8GijOkoUSIv82ZAQ7B/Cv22G00DtfgE1t7718sRS9/
rO2peEVrgBOjGsaqIKUq6mczaXLoXgXh6OKOhUF+edfMVIf2tXIljddB74DNzLiM
2MX2TZf+WPD9cfZHQ2rLL0KYUwZAnAOWKttALbS/C/fP8zNjEcEdhnHWsJSMUxY4
PHuTTbGXw9vSt8D7cFxAA04tVECSG7GxafBZoDNY5reCODXvwM89j2E/NWBJ7HWp
ufVDIbWVItZHsBrW9kRwsVKHCtQZJwo3BhERTep6MTKOKC9QiK5tV1lWeDD3eI9J
v9T6dlIH+GUU8zSjC3yqEsg6Z+sqNzupBTUmhPwJUHei2PpkGZw5MoHIKEnTTRaI
GgNHKrkuIXZaweZDrXxQvtgPOWEfYJmfywR94VoJ03qIVpZIO/aSbm5t+lZ//ML4
pMb/0cjZA1vqN4Tq8Q7NzV7emBh7sAlHNsWajzuYWfIa+8VcsP+qmuIkYKb5FZOR
HXgDFdKiydTelcZEFHLQXH5s15lVJx1jG59P0wxRVhI7JLTL7n5hL/5bZuOOjKmt
q0YgAwPiI6Jf2JK6z6uErg+kWRHu+Nvb9+wVV9mKyBrWDiegtlO5yLPugzZrsD1g
2g8/MyjRC3A/VDSRETV0Tm7zSKqUFouE+oBmrL55kPefOkaM4XbktYzpCEKaSN7c
5//g7kayT96Lofs6f6tt9v4bYOjzgknl+D/CqWPa7oalGBj5We2Z0dizqj49ORAc
1xex2Y7VPptEdZTNmOW4nNnU30z3XFeh0nGG7Z7M7qdl+/Vixo1st+mA0djTWxkP
H6TwS3z85vUEzl9GRXBips0Q+8N0aG6d0udgbEenCD73m5btUiuRr2W0xL9mtxJ9
5IYMdZI1CjKb3/BDDszMDAVXDuBTK2t5rTinnA1dodbqa/YkN59loVwVOM0lF/qM
kAFsaIy2o5AffxUppo0fgN7hYq17LQirGLplkYk6/PDXz16nqkFBUmqZeZl039FR
KbA8u5ib21oACa0NhNlewJAfDq1UFjpIeuTrIYYGVGJfNyMoag+mNmiYUY/mSlft
LJiEAqe496RpYNhe82qOpTUndXSDTvk+OtxsSVeKHZYinJRE7SSmm0BGGoFR1ghL
RHA0ipRDlUBZE7JYJYB8hbJunEk1ytbZZinNgh5GymBqkyNnTB7M+2HO93JUi9wm
b5ZBOQ/pB4RHs8gFPWrHp5deJoBKH8Gvl/QDpl9btg6ch1U822crNLdvb+oGfaPF
8tWd8ZGafBL7oAbH9hDJFcj+Usz4tlyQIREE7uvgKe5oiLHSN/jyQwcMDoM+odBG
MLl0NxTTz7SGVT6xwZk14/W+Cyy3Bo2FY/+3sXVc1G8EDsQkTQT0XkH7zwOtXqgT
brLhrOOumi5dVJhPA8Kfq+TvGJopXLwuCdli5qyWlpqdnjcx1HK6oohdUaDaZTsh
SjCDWLURDMVTQLHzsIl/aeY7ZxSh7i34ijCK4PxyEvjtaqBogaoe2XVffdCIETep
gVZYKiy6hY/YWjtBnUB1+G8Iao2IWWqJhRiYYvfUqrLzCCnm+kC3rHW5CVrh5DbO
DjNYXpsXrAYM4/JC4inJbTe/tUJPD9EdcW3/5uKCNMDmMyGkqIs/tQJaCJXMrtHB
3/VRM8EdFyfcKsct22sD2pWiryS6dwTMy9nJA1xLaIKXecLoP/uJ0MV//D5jjwdC
2s1aRR6DfMKIwTwj8p+UCCb2dwr4LAIPOy9NUecxRih+89rGLRvjwtSJ91VAPlMZ
XauH9/Z8fD5PfYP7EUECAt4Uq0ZcFJxt1g1ssSCyOhQ66IvFbcyRhi+gKdCrUrf/
uyepkSm/mCgJCQ2oCm4tCGLdsT4BzS8TUq0wX7fnjajsnt4rI+Zrt+msrdrAVInu
xw/Y42G05mAD3w5BD2S4QRo8z7YiggPtJnK8FUk97xXPSbpJNxisGBtPzR4XqsfP
SuPnI234h16GKZzkv3V+woZtc3vMudZ6Pid+atB0hkX2GlD0g/eSB0HoXtPq+LRE
giAC+sdF8Ro9bF/dl1T6iJJ7wX/o21DsiSkp3eBBU2pKI/MMPj1uTupGuW0Euv5A
TXGfwOLVNXPft9n8SRwr3+A5y6nDSOuEdtWk/eIJq5PFWbZl45f5uTy7O9QWk57a
DKsZWbGI25BFUjXRtlwvMb/yNeVmGdFMubdSwP6A9lrpksPBdyprGPHpXed3E+qn
QfKNPnhbFL3xk3htKQsSVDuD7g27oTVYaXmAZH5WepTV9bB6cPHAnU1dS0UOwWbR
xlJxJAmMQEgReCgCZWGhCiYQP9dGrGPidDFXAcp7523PUVAO9WQLBOxOY9RrBSwl
pn2AH8v5DjdqM4A6w+aUPHlZUNv8QBPReOwTtsyBAo3sqkMTD3AykCBE8Kynyjzc
qp5D1GXPTioh0lnrfM8adUH7XEdgU9KDsW1wtRea6J5Ad1ALUaMqrDbMvhxGwS45
ZsqA2VYMRgxisrSrTSIVVGTVIHRYOHx/cHka/MgeahdOLU1vIfLLSV7aTmmp1+cM
U82fucDr63Y6ME7i3EB1m62wYzMY27/X+GnKoW2o3uJ/eKX1aa2XGwoT0Vim7Xjm
t41fa1woYurt8USWS6I+7WMxaIkMGCgvBYQr7L3Mfbxnflm7v4bgqH7izoUJLYg0
qXp3xSmC/JiXfrASQQXmg1h4/o+czzPLDdj6XrbsjnsXBQGP3+AfYbD+StyEbv1z
AKzgupjUqdtUx4h0+EdvTSSdAXpueVKi8V5+Wg0G7e1/lsR2W1khtVaRScS+LUj+
UVGvVvy3/x9N5dDaN02wNNA4G3bZvpQVRhyVTkSszNsOQBPeF7B9da/QobvB0kNa
sP6thiWWYstt4KZaK8CUaVikmE06XgMVFsOrs48kEbNvUrR35lTStP4Jow3trl3b
oVO9NmF39nNCLEYPz6xf/0K9y01ku8tlcjDnlsRiXzsKcAjRxOpdlXe7VzVVfEgd
EdOzA6kCe28rEAPJ/8PmPofAlqI/SuMBnvQBniC1phLbHaodgaegqNASUmmBrkcV
dxOt4Gj/sX7wZzORf/EMaWQNILFGadtnz3hHmpmsE+kk3sOKSOi6sEjDPeCAhd9z
nH4sapIDqqceS3cYBsHB4oORJNRrZcqVTF7iDL4fJZ2JjeDMfF8Wx98N6LKVKBT4
LsQHf7QXQLTY8kJuwULzRmg1AEQbPrQAheoX8lXMQp5NkdZXDNxKomN7PsXWui3D
90fTE8Qd/+xBbQzPaljqKsFfG0lAQ6q3RS7e+47RI0vMpwfpznpHUO8htACmo9gt
KwxtgoqH58DzywiAfwJZFp7jkfxEG3FJdWni1wdJiiUufgJxotHuwg5lh1pKvqKq
R7LgIe1hpQx7ZyZ33Qosrl+sWAZdjWoK2ZOoj6w8dBTnGQEz3dgluFmu2ixrccKV
M4FgbRyd4sL5hWWtX1vxLI/CUQNrQmxAasA1HS8eewo1kWVMLtxZOmB/QRdtlyKo
wvgtA0IqmHg98XZOHikvZ0c9kJXnS0hEDpWWXa5ECkmckx0UEljmjCOjez3NPZOQ
CU0hvLVtewbZTWRlxn7d14Du9l+CniYCuMPd+ZOqJ09YWcc3mB+ESqs3+YF1NdSz
ovvrxls8ygF1p3fCVghIVa8JCpGqYToBVqMlB6wJDaefe9QGrs1xYgwDfDVBwgl0
sUDTjdc7BkimAVloM1UKTmY865gcKumuFe1hJmWU5tEqaOzkORDfZ9bItF9tHYiw
Wot1ZrmOAAeAV77sgU7xbR452XRTUtKgnrCHPS8k0FLMookm3y4IagFb5rthj1gI
K7zPYk3T0gwylCguhfzcioyP93jBQaxl2NRHtB2EEtiA7Bcvn2T7Hpg8JwX1QKb9
rWFT6M+q1Ia9ujdyAfZAlF0FwLWzEfXcJqTL++SpIWbHuDLWEAzqdH3OmmYjAJLF
6MBubeFyISaS8vaGcS/rHn+Ezcxy794u0ZoFf1W0fRUlTdAjnF1yPUQ3GmN0Esi+
6i5OpbCV4NygN+Ry3/Ezl1odB4oPxtosX7RKqfnCwgQJHqW8iTCYcaRfkZcodKjj
x+Fc1zl48mgcbz8NvSYMGi2qz6hcs4UAe1S+QyMXmTMBBWonz6KFiC2ma8W3QH9W
vukiyz6Js01fqG5Fcjsh4Q7JqUDEyqOnCIK4uLPYusLPwi+Loq2+/SNH+oJodlGZ
3joMgA3mIPqsrurDGrU3kIvtmCN2VFa5aQpItPgOPcCW95R3D3gdO9Z/9XzuiBzq
g2Q7cjmo7FwzMPGe0A+aB5lHZO1IsDawZNJM6Du3d7Dg+nNoYNP7hgBShe7E0rCv
Z7waEBCzKZvxF6BrxvEMY7EO1P/XXL/iHtdeE5oM6w3u8yeGQCcvloFUwv8zaYMr
ULkYTs5zM8q6JLS35IpV24+ZsJ8XTgWTPJ1zdRLmOkIZ2WIog2PJo0QkgaIj0jkw
cyJ6C2LnvVWourCVWihcUSBDa7eL07ut8FoRgB8kAmTcmW5eVz27gn7OUs7C4sVu
70NNyQQjVOAgB5msXJHmiuHAsoPRStD/Kcca93YMiypbqSpjN8fTf4LRDBMFBHx9
+n0+QZwf9TR8ftGC2SkpF3LogFM5BtpYS911T9RS8Ah6gCL9ydEzp6GuRpYGN4+N
+hRgUD2xOneQd7LDeVo7DvTmTWxnrTpBgpAuIKU4PJQlAzf6BscTyTBMxS/xuDrU
rd/uif5cP4SJ1VJyzXpwfHpiQ/BsiaUVpw//rIp5eMiRMJwejpDDfFsyC5BUDBqU
Y0kbxLQoRp6XRK6v5StLQn8yxoE1oZL88cLOPBCTT0vSIMlnbvOjihdPj5IWJwS4
iLSyUesA0xZJ2shILIGCOYpS6yJEjy9zLCG6MEBNWN4D8/5J5m7n3Kk85/cs3Od0
gAVnvX47fxPBXnp6uuknXak1TXafKacQp3DLaAfwTjHuzrZKNJghginxqcrGfq2v
3eZ/FOWiokBFV2Bk78Ul9T7L8H26WfkLVdft3lG9Fassmrc+I/QpbvCf8kIP1v9y
Bid62Ug5TIpOxvakomAkPGi4Tl80rtfHfB4h+CMMNYQ3TWbWcGIKva2EPIJDSZ6i
LeyucjviPfbnSYDGQF6Rk+BPyzwZBSxd4kxDNmjxHJFi3VSgCxbOUamf4m3XCflw
Buia7oYMQ4cKdC+tPg+aVdg+CWY0aYk2wNrYHmBryDilM7O1Y1hY8bTc9AkXGvcc
x9aNM1db0y81JpcPsyhisqLoTGiRAIIDjSqJbZKT0bK1H29AQ/pJM8UPdiWlnAXP
RN8cyY5shkVc0wly0thVzpW4T/o2zLgonmsncTabQnZeCTBk1szAoGTLOE0wHpS6
jLwVuVFSMVCjvkLVpCa4QJXZolNZNP9pTU0Bbt6Q3e9wYOrdEgsxRCZCp6Ax0muC
IWbXsboerbTX1xPhZo2kyCfWLex9MJAxkJQmEHk1+ggt3An9IkjHDrxwWNe48L1/
wTdQpSzmZsQSvOnn+Vb1rkX3ZiFGPbUtBo41bdPXk95oY5bGHWzwzlea5Yh0qR5V
pzGQabjlbN2/uwzb/DnphYMteBmk4s3i2FOV4qKiK04Zun9NOPWsyVe5EY+UvAyz
DQ4jgXmuh97TXvFxUqnSNuZJoNpu56MPaetOPtFAHR7puBwqSK6bzONoUq1sk//l
oUTgcJDfYf7mvdKW5ENmInJT2OyZ5GJo63dXARUpRxkdyfeMhYDNSExmroYhWCYm
uG4MKfGjdLDRLBdcS5OkvDcgFUQfcVhBpvxhId6Ygak/+N3xBGqJwy7rF/QBIuMP
gPMp79Ck7x9MU5Fa87bnv5k6Iv4VFZjcr+EPA5s3pHmEo5TjIOqauoteEP5yhpFh
D6Ed7rYQFOjDkLU7/bViEjgMDEUtCCVDFa+HMclx2ofG7ZG2E63Uiz6k1Q1p+Buh
0hGX176CATa2jFrNvPWhY4grjKIzJ+48Qfgx5H7CopML+z9BgnmvUVQ5fct8p4xE
gWLZnXioIR0RF+pxDuE5Un93tbfIntniuzZ+tVKfKesKLT6GFVPeckxSBAOSRnTA
eKAGU43rsj1BvdD3TDhOE2Hs3UMNtbHwRQm3TRuWfdsB0e3oM6SqTZ5Af0DdQJqc
F/aF3isfsXOvINNUpaiq4koD0A525S4/EeY+EV09DaHmICF2A7ihvoUGJNeu2OFR
IQBi3A2uodIkKE9s1k9rjfTCeLzYEAZUktNRJSI4yA7Ohh0F6tYRJM0b7KFoeNLA
oGdx+V7H5osR45AwdQ4Ha64vWKu+hdYbwDwW2pZz6/Jn1JHMavUwgg5QjzyWEd4F
WwYKQyVtdZrIiPnzHimdy1+QMJ8yAKPzKs/Gb7JiT0gpwQrn+QDIWa8jRlAuB44u
wjalsNrRLv+C4OidkawFzToCSGLwCTtYqgOz1gyt7qM7B21m6wFRasdSPDuw9e69
t8cPgBu2s1CfXCAGTkdzW1235pcQXI6DQCeUw7fjlJkKvA3sQgMevSg1NLMf/4YK
FBAvbyEZKgcx/vSlpisAS11m8wWFEiKEl4VPSbh6gh0IQN4wsP1gm+WnuaJGhLUI
TShkCJ2/XHhsZ5V7UOy3RmSE0PZFX5x0zCShdfu0qblQWtnWZDye1Omm84JoDztI
Q55Q9evlnPOAuHPW04AMQnK4D973FuSZQEVr9Mf/HnZ3dWCyqyDwdnRhUf05fAxn
uOQ7r/6Te3TLHtN2XucusSMTkgM9FDDNViOhoDT9LpBW2uVZDsfREUTUI4Tltz7K
VVEiv60nubeC5G/ogGHtz9fyqpvAYwpUgzHC6mlfvrEyaRdsrCAIwxYT+nqObzJP
D5tp68M2GD6aBlPUMl3CgQYm6AcgEWwvlaXUV0WRNdqJyDbjifvTW6IVADYdo56Y
qmREdGGsf2ebaW7/MsEBS09tEPhi31P6tY7lIXPcqEgWH+0aFBO+0AxetSKsBoRd
i8WZ/7bsAGYYlBFRBNPxcRz3l3Gz7Qrgt9M7EXVam136/EesL4DZOdOjoZ7DcYnY
YxRD5Kgb6PaKAkLdQV90EJHgE6Pw6rJsAsyIl0u3pwrJWONbazEkMEUYwYvIVnQy
Of7ojCqWPirJN3P3Q95z0WBvWomJXrCG1T5wFBLzhrbGvRPPwgUdR5N3kEAae09W
0d+GsWUppi1jFAiF834sHTFzekL5HPbwFuQZoQJyY+o0vD41Jc3fPh8NMBUJEYgc
dPiXkZCYJ6DPFr/Swdw2LxpfVUIqSBA/TlmSdJctCLVMHCqScWxAR5J7NnRbe8MH
j+4YJ8F/2na3IBqxBgdNJfIdjhRyYkRYiGMpb/v871/O2BF6AUitxHQr8GQYbO+a
O+QuSl1LbAaPH+9LOp5K0LqX4cTRwGc1AQHNT7hYNijoFeAhxe5Le6NmwIyKPgXC
QiUiRvDTl0k0G7MDrAHW3WOYmNFlveuS4tBZZ+6T6MaKbJJh9vlKhsu1lx9jkR6M
jFXyRvYHXBUzrDeZciTcckjjEcXY/TgduZp3yJ8VZoXd+JoF8wz98mJ7CvGAVmov
MXmvuUHYRiAIg7mJbLKaV6f/VF45f0hz0JsBHngh90CEq2+OzrH3QQ11fEkVn0EJ
rmWkYhqw9Ntve2rSOME/WeIcR4TTY1ER8bXDaC9uRJc/mkM7JvA5AY3dXlS4kusp
xdjuVZis3fwWskQy0CqXOY2pXe51HEOk823se0UiL/HaB40Zgktn/3Ycm14NpUKh
N8kX3bL2VhCaWZ9LQTFui/GzZg2C1wbxxb5geE06e+ny4XF8ecqD3WCu6lkCGFZl
NV1UeYMxRrHI2tfWmnO5o12pKhGLxuHD6WiRuwyG+io2ZSjizc4oU18nHLUdLWan
uS1Ex2+sFYpYxz0hhxh6SDgGY8ussnnO3DHSxJ/dURpiiIjmhG7j6sx58IIqq1bN
1cT7S9M7PSgShDWlqwUUyXjS1QMP9BTsnxVsKrwUoIDyrTsVyS2E83fH5tLlFBSL
sZVgfuU2stbCdRN2C/gZu2d69j/skU1vI1/W58yXHZZ7kiqygGU1CIMyHEBxfyM6
rMcaJSIJix3URpzKVaoNiF2rTsH5pAhXSvDDGZQgs0IV7mFtewIWVjLmoTF2vj/p
IFF0OuD/Hc4fUT0FQCDUP56XkBFNPFMfJvi58Y+RxEvkh5YVC0XZJFqhK5NVratB
YZIkYYSJzwLKjK9S63kNLRF4RYMNM+6LCRHMNYru5bR4I5+R6khjYWNMe1GzMzom
jh5UljRlMG6s79vZQSv4657Otrw2gL3LcjBrbimJ+RTFgPycfvgubGKl+ytmsaa2
2ZHJYMk/5dISgnogqwhXlwp5M5nsch7uHxb9rqKn2+0VuTLhbFbmsvKcwCPaEDDZ
EPz5GTQOARvCScYKG6WLUta63yrjm8q6tgSvm4iEcPyXGVtkvhJOqGssHPlvu/jC
2Rqd/EDTNwVZBYvEP5xPN/GOFUAhFJXbzaB3jH+yzsqIQ3H2a5LS7rl4PJICDgOJ
rbZY9/qEpb/TDJQ4v+YazX+mHm/uiAK9DWgBjdFRG8XhDzi1VEnzd543iT51ehDi
aEFnfxHfy+bdnSzKzTSx9LKrHlwsqoLiqPbosEx0J+fsl/k95BtAMDBSVppmF3n3
17SbUchGBSSEnm368AAwU7pJ02r7JVpJP8hpn6IHenost72rwFa/FIcKO6+T/o0i
8Q8FCMyLVZrcpKjEt+A437TesiXhIu50ss8cpbE9sJqHoQyuFrMUDz9YrwldSXCE
oXG/yEvd+D/VJyEPAoMwS/kPTSmBPfKRd1sl+MA2m5HHxaR4HPAZX5rrqdJJ/1ce
FnivbyXr9/Xw/1Q5czYR3E8+30d5amiwkk2DjdfQrHrI13R1IoXBuxA29v4kzjTP
c4HmKSojZzmUffso8+yaUf1MAHxEf/O264dzmSuQ37tPOw2PvOGBDaHYokCqJV4H
P1V+7b3Iczffb5TXhxifpdh7IcgVEiW3gTrvr/q0v8Vl6ug1nze+m03XXv8OJm1O
rgokqcDPRewnNjjLtriwcvdZ3BZcGCP1e0R6g8XLUZ4wQspn4qgkT+vwhe3Vnbcr
5foX7v9aAwsjloBaX51TysCgRgaGutTR5XICEj/w5RNlZb9xS24Gn2kiJdUfVS8j
O3Bzgm06gFai3A/DjTpRdIRcFpQgCcPdZ8B1segDNoDwDEYVtPCUofYByVwVwC06
2sCjbzt9uMiTjDZsbL5MbyF8rLYFdn1QdzgcpQQpNJl6zV07j8gqeA4XO0s5Ad4f
h8JEhXb2RvHt12dL2V6TdUuHD0gA0t0reIB5kPHaCq05gwH0aM9R7eM5Pv1RqDZb
KQh9ALa+in3vlYldYukvwyyY6tmafCb/8QxF7wYE7WMKJM5GtpYWRn6scM5sg5Kg
W8DmGb/pkDejSRkzkBSD+OlyMb3NtnbyMLtVzxEGLjeWFYBHnQsReWkqMPwvtmdt
E/RoNsqnpmS+E5UIeUTRwbFsUNx/nO+kzJ0IWUWnDbfBI39UVhhcZh7I1WnX+J2j
uWPhYNVTCJ0hEv/xIkihs3SXZLf4JOsiYqX6fqfaK6olhP9LGem7LLIy6OpRtIBY
NSi/Sg6kOdrOPXwHdisuyYFmR57AjFeBmbPo9I/4Mlst9s4eoC40XhRFcmW9jePX
5VZeIcypoLZSviutCe1tq7CqPmQ5E/5fqTuPLtQA/iFPHoYROBPLepgNQ0C4VrdM
VhHT9vlpcoX5NQ15xMANROOcZEhtBy7i4W9VX5iFJMDio4YedRftFsawUrmjDFrG
cvpKWU0b3Ri3EfP/8LWlM0/7c0EY299BrHJF3QR4wr0PpagoOh85ztE5irvb6kHG
M+aSlRsgdfluypBLilOVW/vRC3/pbCXt/I2BscuT28L1+WZc1WiVidMGQ1+z5knc
CDVmpBgLQ6zOJiTZU0V05CvB+JLh6+4sxj6JQHnKPzcTHmsIEzabcAj05UdzMNZj
ebbkBJZKkQheAwMz3VY22YvPfsULBODI9RL7KTlRee3/+C4L2cpbUE5MkXrVom5k
jFQ/jRUzL/mceLhU1Of8YX8Q2smKE6UQZHCJCDFTTkdhorhEUl7geusHNtx5jzMn
cYnd+5N8+gl/SXtk1ftwuPgGq7BbyPp7ZuY6e+IYkAMBUTfvHYAICOpgusluvT/m
rHD3BvmQrgcfV1Mjwh4bqluv++FIKTNFPsaOFrPBOw2RhCx43n+jfmzOo8gKsBtF
zHS8c3MG+2WM4r9tq5pndj07kPH5uI0RmO2mr0Ha+0yhtf4kx0a0cBAl3SBOqhVE
F7WrAGDO39oiDMggi3zpZlgQjMnaGa7+KxpHtkRq/QmbmCZtz5lm2NrZ3NPMxyRa
MmFHMTmWF1Wp2z5Z5K8zWUZ0otwB1zfAG03giPEN20hLfo9chBhHxqe74lalcmot
rDD5umILTMSE2S3EkIZfMUUDjtjJoz9mC7JDWJF3beLiGZjUEK5Lb/YktN4GrMgd
46jCJkkiUmwZPb+DgJJb/MLKg0FJ7Vp33iKGD1cx3I8ntXabnSlYNzVQtC71iQWv
K1gvCNGpijMPcsAwmEhwQEPSUMNlkL7o6zXO/wt4quoIoK4Gr+CX+Uq9XVN6U72t
JNBS9T/xUCix6SR7Pjy0w20B8h5WfcZgplKV2vNujhnEWmtCvv+48JnPTFNNo3V8
z3u+VwKglKh1/9WSNOnPG727lCJr2YTmHPGKACb/m39Ya9w5QLdajSXEClKlGRMA
ZCYKftB9e2Wua5X9jqdb3S3a8WfSmke5VbjYm++IjPjwns4/PvDUfeanWbbgOzDy
eW+qFJlb/xZImqvm82/M8qQqZL5OZd7KcGv13xtm+ZabCxRhc26+AaLkTLWD1SaM
cPR42fQDhI5XQD/CEKUk6vP6slnOokVEKWwX39ilTKTXI01XRL5mvepQyoyFN/gI
TcPAI9QVK4MnxeyIswVNQWcSz45rHSR5t22CkpbY91BsSC9dCs5ejNyeDaXJ4CFM
0tYZqbnHKGLSnfbme4MXpFNyehwGssf5aq6kzX/UwiixdSaSqeKeG/7g/sytiYlv
kFiQXQF+99Fg7gu1/O+0xmq4fPeskMSYJZFR46x7Irg9SHzhjMKChoxB3iwM6O2g
pHmddBmKZFoeVuAd8mXUSi9R1NDoL+k/+ZddGlIsNn/0esK++sxsr9gFo58To6So
DBj91BI7TZ+GLw5qCnhymTkCL4eVAUxqJyrOGbdhLT9i/Ng/+Noowum0KQlFGLoU
pZ6qanGUs72YM0Kc9sj3qFjYR125hwL26nKcCOeMZ8AdICz5h27B4zW/+FwSBuPW
RTNFDRgb2P40U23mIYgNVq4JMiUfXLMQZU91FaZgT7sDjF06lSAmXG1PG6fzzevz
iqeFR8tMteEA5i6Q7TnmRKeuev+POUcCgZLMnvtIb94q3MwOUMraVkA5J+fkC0oy
874qxz8oqgE3ks3tSFea3Jw+/C8MlKHRS/y0DQ4T5kYg3Fwk4cjXAFljbHU6Wpbv
cwQJmhjrSnX5JQnjeXDYXDbIvOlwU1TYO1NB/FhE0kEXKoe1H0PjX5/nA1Bf/3cF
9ozOcW0gUstz9ZjBFzGZBxnhyx8mhexpZWqRMM/Wm2ereyOv5TNB/bQ3+Kf+lWyI
RIAPrKN17hB7pez5OJByv7yTpqnIWecXWEWxoVCXEXFrpZaA/aqIWPoY0cg9+k23
zWTn16OkuijiYEbh1P81RdiwDTnV8NVcTfx63qFWzTAGWFQqvEpeF2MJ1oHuyR4+
oHD76u4RzLPc5FcLudqXbpms6CHw9Z6azAgMnugfd4xxyioYbr0YoUxxBqqmLiG8
K1NGJHbXugWrodKArsSRemGbRe6sBNZNd3vYnOolk1w0Q/QgVv5KKF7NSLyS+P0j
SGynv+6N14o+P9r76h6you07hD91EJaja2Wg87d0Zdw+4gYYn4T4OWRQMuqB3HDM
AySoJGmZt4N3Kh/BAXTczeZ/na5kostlKAfQTmNkPvBMyiuoXSCX1bT0hTYmXSib
WEjMlOu/X+e1kp4x9tUzRkTE5LLWkL75wr4nv9NZyRrrqr8JNKyu2Hry3C7ZoYh9
3M/BCsGRlBeL6AsRVtat8mchpocBD6d/QcxWKIiZVb/g29Q5TX7ZQQvMyABNkOAP
Fk9Kz5WJAAoMeRSCGXxAdcHYb5oPyUZuHXta9F9iH74zAYsdgEYT+NQs7VBXTt7w
XkjwUm8tu0uWHfJ/w0JMu8j0DfS+RQSz2/EJIsl596v4LaWiORrPMwiB+JfgqAnI
Q5Gv9hfrRsTXFyi/DK56W/GpmAkhNBHttE2hJ74eXDxdDE78YfzK6gmiAFCDGXoy
z8IkLDAjkN2mAwJwF9Tlx3WHSsqoXwXnRvPGYHGon8PhI0H/BgzvvaMA6N6iDvon
+py4RtVeAK+818jfZfiBlq7FVE3ZfxTnkyAZ9vPRhKmJlanpjh2fZjdwPracxvuA
rr7Y2yFhmKY1ftQjLn4IqxswB4F+fW7piz/OGDtz2XEu+rHekb7l+w6MG+DHMPiP
iJfmkrI1dZ8e4Wk0XBjciHrlpYM2899364jSgIeGxqECcY2nrdvv91qIi2jLI9l7
RZhiVwOkgqABIIpyRPjvU47/528//3GBLoq4kc+Uzdq4G4+mLg6+yeCP4XG7/AGo
37dI8KyezKY5gnsk6A7dT1TzJohLEAIe9hvfvDjMM5s5e21r3UeUkLZxL4xnQf6h
AUsdXubmaT1xbrifXkkoC3VvWDoM+fqgTyZrJ5V+URyqp/sDbxrDcQKZgMvEj16H
M9vF2vi6XM8DH8jnQkg0LmFUCK8BPRZ0A1n5EgDmGg/nrm0lZ3j+m5A0F8Fg8Dwf
eIXuFa47RXxauastrLDMqW9qeMp36SeRB/a8XGLzbixQi4DSNdrJOYYA21Qf8e+H
nQnQkqXyLOPJhcAywnCZCdYbIwTO2I0zN6kI+nHzugWCyK17tpRG2BNHfWhFv01c
MG3k9xYc7TCUh5isVNazJJfqgoRTd1VvDEbdQ94b3xgm4RKPvB98hInzHRaro1fc
WuEbS0hO0ePWksBeEmJSx4+/j6op6nrVg25C+Fv9YMok8QMNHmSzC/MaaCOPb5JU
d40jMY+xaG3jEM7LWL9kFaTkm/UCiKO0TX0pUGJWLdcbgOjNtDkGqxFL6G4zmtOK
3peYzeHga+og507i6DqzLvKglZi1EBhhLCMoQq+QGeAeGm7KSC6gtbQu62qrNQI6
7N6QSy68a6oPfqBLopxZRt1Y2PUh1amjKQ9b6Pdaobi3eI8X4q1f09T+9rCOqX+1
FtxDr67N4QU/cWtVdeIrcxnOOG7RkKPvU3BTwR1HAcSgN0s+ZK1xQcO+GehsIg4N
XEkOByhtwhZO9A3UsxjAL4xSOrVa4lwQKqM72x1q/2WFKoGmZpJd4dN9dH3i+9ij
2z6L48lY2ytE+ArkD2eVgu+2Dilglk+zZ2HuvIYqc7gJCJcZEysTs4bmUN8b/iBS
+xojXOiuUu/IuEmg5uqsRnFOW+/kr+eQToyL04rGeUwMUXal8F7qZH0kke/0FSA2
5WvqVfDribg572aH7r+BEbkL2YGs9Al/5r9RexOWOFYQaoX75LEVqfTDIfFKnprv
hm6ArH9lQXE6Xeda4XadiLBlYobKe1ymgiat6J1T2doOUrDjfYU4eWtNh0wPyDrl
ZzvvYjmGw/vysbsCp67FGkYF5I5s8Pvs923zokCIkDKgAvsmRYdeGJ2NGiWAVBSb
uhk94hR4/rIQuqNxsV3y9+w9TsgKrfjm/SLLTKHiIT+7x0UuVuZLJXNQLBGWQYYT
SCnkBLUX73d3C4GO5C5DKVyIOstpvtA6KAqKfAyOK/RDLH9/T9vjBsVhyKQzSt7+
KHNS0miYXMDD9BjlWWDSKrLfwH8a/5N65r1MdgnyL0el138vrb7BRJ0qTafOrxOb
D02nNwYxDrkZw9fBiqJ6CSOOodnjjXgm5pLppH1dxHEaeA9Qj5C4Z/wuPcydLZkS
UtzRMe6eFlFIhMJFhA5Nbemr89VF1T/kDmC1z7/Qbs7oHiHNt8iv73QPcvWGYqUu
PXB0dnjm/IzFh9uIqxoSrbKn0nnDxOP+BSN6sZcNwgb2bbjEtj/xnlNMOeysOKvl
2EFyoDGwJwbEXTAc4A9afmrFAohDpoDPDxnvculgSSGm3mdOvzaEMuYUb1nyTorS
JEYzCHolw8oP4uD6nBYdH+XG7F7YwCDvaqksytqtWHHR5Gu5qiT0F73Ug+SyDoor
XKTDpa2tK5MLiI2a8MSJrQ3lVz2nbGR4Q1hrWujF3o66S4sH4+adNPZ+g9d2akoG
6YxY7dMNQmyZDRHrA9QrsHTHWp0byWaMXI56fICQgVEcsRRKxK0rp9ISKjprXKfz
8VcD9YzqiVoWOJa9txY/A7RaZgSV/5PbZlGkmXuwCQ3A3s5KY9FEPoLndE+lEWG3
u4ABXRBe//F6G2lgbkRXndWmRakrkoMlMAY6OO0pI0upTcnv3eLJbaEUP+7nMVCx
wHYKoWZgHTaXzYytKGrIBXR3Q0h6e0Tz4T/dl2mlfzzwyLfiMerTBU2uSEIbdtNF
DxT+uO6BJRY2nrysad2n8dmL4takrAjZz2o3S6/fe88jGz6yZ4l9boqWcSJUU6rh
pVag9KmMYRDwHpovmM7cusNH5n5Dle6d0nYbXm1oxFgmJ/t5aC5mWLZES5mL0eVg
pTt5DubiCaYMd8RIimxneBPCSGdDuIME2kk0CJkSWC5jejTqgzPuYPxep7rG3cTG
iSwAL25TkeBfWCeuRZPn53dnVEyqoD/5RB5kccmI/VnR29g0fTmrUu0tin4DpJAh
4mM54XL2zET/T0mVW18lXO2xnX6PtqXSx31R5NP2quSVv3wLwWfpzvghQPPvCXdH
MCZp/DiTAEyN1r9pGl39aFgON/BjJ1ZMfRwx+QqDOkEH1ZQMRq4LiWn2cIUznRUJ
oOB0pBSnYkjPoO9dSfn/PR08JF5JB6b9GyBFZzwB1ipUGHYzK9x3+Y5S6giKtknj
9of5cdjHLWjPCOHUrjNehK6v0t6reec665GoU+HAdQC3Aob/jkjWqxgxmh8WACot
Oz9xhABXl6amuF6uwSmhcuqmdpnjeRBo2vTnV49sjUTxQCyF16GJEIAO+mgETe/r
3WyjYmiGpF81duJta35aBQvfSmW66rUT0IsXazkYQiJPxfU+nVailejeipNiFFXp
LP379VQSnM+gu8308lkSCdQqww5w22W+C+PzNjR80SN6HtRX4hBJPXs252wePBQC
h0SRDAOWyZEctgACeY7HevG6dCYorGaEUxXukgjBSko2BtQAa9bbgV7Ee7CsSbsI
phRY7Z/vHTjwSzPPpfkPC6uWCAZReoZIc2HWH1RSsYxLSgNfF0GeMkfv7G0ZvnA2
vKd3Fe/cQjDUz6CZ7S/QBNJkqlDAbXKmYwWGjj0UXu/QxIwI5ACtbCcAy1I4XfTA
nu2NnzLSzyWTSxRT3+VL8bpA+SNSsHDiDodBp1KKU1m1KV5JcXQX6bJIqsOhHp10
cNpFHvV6lXL0YbqqtGN4es3K/q90g5bi1pqtESDd2keg9h5tzbwucIfClOLCJ6Cm
5WdoimPDEM1hl9HD3StzStOWayaHo5VhANCFRpsoL225euBibayeXhORwXN3qeMm
KlvSHZ54yovfIUlv6Cstp4xEsHPzTUqUZEhrdBWvBv4zEhb6O4mvTk1cBRXNjsnW
qS9EYpWL2RFxQJEVqoROHVWJQWmY/EkIYeV/YyHWtgq9mgW91kcMre3bVyyMWXWq
dedtW+gCF4hkk3INyxj/p8mXGv7miDdhcxAe+rvtPtjSwKufRK/fCz5Savef72F2
//syTT2t3dmZWWV3pMaTLim/ouOQEp84wqF1Ctan7oUv6DKEUsyXqYiojM6Z9qTq
A71X3eGRWy4OMK6zwdTE1cMkgVLeC45DQyB8NsYnViQv1+4ObbZGTHTDgVSyAW2P
JGNt8deu+yuss3bkAziySLqpeoNSVielorgq1o6ALr9+tq0oSwYs/yZRU7j8zHNr
n/IHwGjbgdUrnfcot7U16rG3GyLnTrKq07M9CnhxiBNhgholJnpceRhhg/9/Krk8
tAxEV2ASedDpTDbrIlh4gyqB/jqMvlBnK1rGiz9B/yCehe8eNUymfh04gw8teHCS
7oG3zdDP9owQWNxrHStd/OUez5d3LmFomqBtTFOY7vSebWGSK5tWpu12IXMCIkW3
nGNdpz4HQMQsSDgnhp24O2knz8D+mIqdSAQUBubNggnB093cLQQ4Zzlmt/suaGmY
7QATBDm+Ec5K/ZFNagD03YTJkZKPFdYHqw6sP8a9X1EoLmFuJILhPX5l04ZmjNXm
5+Pc1aioxsP6LikGkX6I1Q/GtMpJj8jc0rtWPv6hfgAezS0q+iOmUYZEE8HYn98X
TCj37y12b7X+e+7SeZHBK70zfp2yY7o8qJcO9GjyLdOuni5lS1jd4PbI8rGCN/7F
5+g/4B/WSAlE3qsb/w0zAdAImJ4hAH1oYhIBbaXL4bVnC0A4addhPmnAi7fvkz5Y
jVzJ5Wvi67jacHgdwO9lNDr8ZMN/uJoUfcKSUsNLsIHNYs/bHkdW7WyBfm8AzuEx
yJKyeHMIxbgZyiH3/2ObguEeshigQWmJ9/Qu+UK3H+kXm1St/LPRCqImS4pF8+TW
J0aYGsswKBr1OR3VdGD2Ig5SLhP+F8+apXmsJRG/9KtGP7WR4utwgnJYuV+rZ5gf
QTN+jnpWVf2l10raFWoObh/8dUCvQJDepI0NPlfUAv1QpmQYR4uhfyHPE8d3iFOq
PK+5hvh1cp4Urv1vTeQbpLkUbnEBCC3JSwe4RWYEdOGXnZWTW7yOKdgWuLurwnPL
oaZHX4Y7xbu8nq9qfU19yACtldDxnL/rtCYIAuD1JKzyH2Neurzak1g90Of3PhLy
3Ct1wpfIGyWf9oLky1FSZX/CRRwipq07U+2Bl8mRmjlm2QuTBRiNVfeAsluIE+VA
GNtblQPpYhGi5pHBFweHBpgG93B75tEFcZpdft8z1WJN3HFOaCzBDdsKO7yEJm6y
hmmqNR369lHkwrMy7p+WIFUPw06jUmO/9r+j6LsRLBeY7sIEfTZROGIsWxJ+3nmR
H7wOR03jQoMfHQ+SmAMLmVDnJBfQEWfvh/+RfgUPt4bBARiMuV+RZauopSADgYA8
jqNkO+jxV3L2eFihbJJl/ESBlI53fkWwyCxwWyCII9HN5MtS1enVORLY8ty2wqwt
becVITY7YJXw4ptYQeZQyvrQWrw88ztPtlcE3THeSuTZyTBa/j8JJcvbf7Ypbw3s
5Rw5YVzPc+bWf7/b3tchPXBqqENRFvxiKKApK/h6A9HMilKZ7qmEcl/cAmvkbC+s
8sd0hkiy6EDXq3+HX8fiYbmvcf9mj4g9IYSTmHr9oEA5OGXcgbQgZiXunypEOuwQ
l3duCFHC/7rgfDqD7Ff/thxL9KVWxKiH0G6rvjo9hUl3WvAflqxFf6bODVuR8mKM
xH8tVPwAZXspWE77VJfdt3tXhZpK442IxDyzeSFi8+L87WisiOeWZH81Rw7hftg0
haoVVg7VcPle36MMUvvPSERnTEZyNKWq9KVhLsSMhwaZIVroKS0iKdTbGYYJuLom
1QJj2kZYjG26MxOeQvASbHijRtmcQIs6MMyG00cwGaf5GSOtQKf23iq2gXRJ50Uz
N4TFSWcgXZtlpa+/tDK0E5ue42i08fJyB99skFneQcKx2eo2q2pGv/yt2o6cnDZD
qwfMlG2SizMqNRoffQ8Dwa79/29jdmlYuW5ERqB9WQDOSrOcyLgBdv8X4GblWskT
hnZ4n/bf6Ypfzb8AO17Dy6vRnb+iNw1M5i7A3z+KS5aLsHvZNNlzPhw8M0AyA/tN
LmjcSkfnI60w9OOz1Mim9t3LXcSnCe9qU4np83vZx4cQ+b2RraXfdzlNePoD2u/U
OYnc+BOrRThv1IW52oRTpYdeTc3KipFPBghfx7J25+JbvGdjUAaWlVcvp9fjoRxA
knIjSXwyWOKaMwJpQwVI9s/eZCkFR/tgkUDWBOdLZe/nnRgA6BJexuGu1SNI8aTM
31xt3l0g/UM5xLHcIJB2jzEXuaML7tXiUUFcpUZvAXF9PuFtuBEzHcteJHTp7tQg
ij2bQiVRymqE0cFGe4EW0WdQtD1K1uCuVRsOQbdU/w1ZK6NWyNa6Hbad11iTltYa
gP/oWAFjvKCJjltkYVzVXuV5NQvae9Ndi6i1Jd6Va3VgAJVJFpm/+ZNN6m6XSXPf
ue5F9I3qEsS1D/1ayK7DJ98gzZBxCtS+fcMl1XEejphKpGkySz16FEGFPXepX5JR
1yLbu40xKw+f/Mva0/sHl68NJTaQKKsvxkEhgWt/sIwvMAACd0HC+P+QR/NcfyiV
qfStUP93hogkpgVJh64Bdxd0DCxEz7Ncc+Nq9RBylMBX4u2J/0p4AVtUHDO+oL4V
ySFsfCnw63GQN914DGznewWESgL0d1GPtzDcx7Qp2aopfaouOwcc7YgvfgUAjPU4
9PYtRSrvyix5CTnLUBQXP5S7lKSvx6ropfvcUAbtrZDATl+jVaTZiydA2nEryR8w
l/KmHScHecLPvBiC1ToxLCa26sm+JOSyEm0GTh6qDbveg63pERZYQSweER240Ort
ocB+U0OoA3D9dYrpMqbmNSjx45IxtyGRwnap+wvDQ5JBAueRgvjev0L9jFxSGUol
cpsQiEI25lvvd+jlawQ7YeZf87gHIlue57xk2NZp12F06DJMKu85OkYhjiPdO7AU
vQgKvVqCWsR4rDw6kqZSrIZ06Jb5y8+MTfvV617XzdWz27nC4FNJVKkAKwymXBVz
o2H7hHnUkNwVNsgD2SLs9wpz91mUoRgveoKIuurCA7SiESfpJkjRQIKrP+fpUNii
Qa8y2Kf5lcVOvNJRd0qbV+WNIQRCmAuWJZ6ehfLto0TxpR20G6zdIg6NJl7h6fgv
n/8kg6sVF8NwrXZ/jJpF+BFJ0ViPacwVp4k1tIzEcjqPCkugzua8ztxbJN59qYSe
vThKT4g1jWQi6MIpN3M1iAfRI/zk4NEos5aAd9woVOfE3VLeU8QBCwzbhE5EMoQa
LsDvr387kFdsHed4FP9Kdms6fh4JR3tgn55qj4DTQoDe9yjONq9RApQzl7n20v+3
zr0T3aaFMwljb+HVdjcvmEMku+5H2aJF1Pn7Gr1LdwSBxNrtoTo1b/Lg3JNbQPdg
WxmsIyNA8QegRiwofhlBytvZh1ooaF6hbRolmz6ltkIWRwHdvJzpRK6YWmze9QZs
clV6FMSBEh1YbjZxqETBSUe7of36cNUs+osoJxuFCFKae2Vrw7nC29EojMEzefqd
Zq5Uj3ep7p2Tku5xrIqb1OU1rAfDFG+dW9hbG8UUAYBm5OJunZtIVt7pqRR69GIN
PjKQ4+D3fE1n9MCUVXnM56w1fS0F26J3BLMQrKrcDGTyzlKb1bFLhGNVtgyyPJ+7
14CTtGRPcYH1wR9dlmDYg24iO7ckXE0T4AnG6sA3nKogfPcj0QwFyjMhPZfiUcs/
dnL2757wUdHfVidIDFpeTSPONL6BFSc369jzGEsOnxRz6nKdW3BOGyHJ04FHBq0C
VeKSB8CmpPOTjWqKFi3JnoZMmOne1ptoUu7F/s5rMjmC6uMcUSBs45blw2cmhQS6
MKiSgvDQEQCIB7R237777xbjNjebzM6M4tPAAKNTg9BzzTNlRzW9ExwkGMm+wtCh
NVPpirekCijPZPcDODlROY7M60XiLqOr73f/L/Nkk+if8gU7jc5wskjKk8GJkyEg
Ti6AhV8ObXh4l7DbJZ6gXtLX67BwyxSd7Gcqi4lYkkjNCEYJheOggfnOfA2iBkD3
VAB3PPTPE6WFP2k0N1oNmN/ro/HDwbe/Hz4HVnF79iy1GoG9MeVP0XKUCGJPUBJk
y4QpCqw0QklYVMk/9cBz4/XOnwks1HMOIt0CbqAEBlFI3Cs0UNk+bTlLJydkUr+o
mt9bHXcXrwfDRuMFX+/Oas2E0EKfJcwpcAYV2RZnIay7jV3a+eZ64tQPR5xKAVqc
qZpi6Sz5jhF54gJhZdpbyn2Dfl+IJ7hvzSCqJk5tWwCNoH4HHgBNNfWp9F+OgpXK
SKPr8cFztEgS9xmPRbhcW2ffPhiUuxUxqnnOJxiUYjrxcxn/EmtqMm7AlkoiLhQs
aVZQJF3dZ8ydzrYVyh1BeL+rWqZznUPkP24dLOMCUNbT6seQr/f8UVc3OLry9XzW
EqNfzM0CnyIkQ7zkLzIT1yR/jQjkQhIew1mZSnqgc66n4lfDjU29s1lc9CfXNHE8
uvAD/qqVAy8Zb3OSQ3bwQb6c/2V+QlboceMh7rYODsp2svLaFx9jgtw7H11ZQHRf
/0WaSWf4D+db6C7CpUl05KK0FaDH5YCsBaVaN3se/GMYNOMsoW6at1WH+gkFHsln
/ZywcKyA41GwHLWJJZvPCI1t4D5lnjWX5kj/vAubEamBdUlGRtGnYGD8IKFJQACS
ghyNzaFwTRvkO2E4EfeK4XHmpg4tj0wWWhm2y9K66PSdeQayG+5bDX2D9nGivnlY
n9q/cpEkdVTObUOeLktC0vD4FQRX7YyTdZC6nxDe9S+PsaPyqBV2VebBiyiihyjp
e28ukLVMxLGhpjkPnSyc+hk86NX6KpRcguJMa+8VotbN4cuiDk8w7O1vFsOt4LOY
4Pu3g+2avFudUmUnKDItG5bFk5rhCFTqrua2wyiVX2/D3ZI6lZUEegdrR21WQI+9
udX++Ah9lYhgRxqWwPMkaUfjme7+V/TFaOmogakVoC00GpUsjYrsX/6Znu8u/Ilk
vDxy7PNv49J7ihgGiHjhprUSn5PZRcV3Xxte3PYoPelsGJX+2Ls2LJrvluwEZosD
3LAmj7ThMyZ6o6My4CPaZOzGV9g/jP14MVNPAlsmh/hH93MTZzmL57aYTMGNoZuN
0paQdsxmLzksUs7FL0qtdlVCVcH9zu8QOGxX9RVVOFifzTBc3ovKsqR+TJfFHdUT
WOvzMEUaPj3P2LtuvrS+/REKhx8UhMpphUY454lwxmavKayW+Vc9N2ZSo21GyHRh
7tEHMi6CyFFBk1FGruIzx61p3bcvIQcrU++aE07zcAhaKnB7+1gcJBXDxVSEDW6R
cFHcy6d1g2W0Gv25NUbWRrnsM/K2XHv166I5XMe6OUn0FixHWRHi8gQpYSFKdGBX
uYd+jPnRR+FO1El1B9Q4upNlqPrPqL5HMxFqaMHqI9BEDOLrSB0D9qCd0hnp4mVh
Qwyyp02OF+sXiB9dBb8zumL/TzNT3XLMV0YNVoAjTxHZ/7vxEpxiar3njD3P36Ww
xVzK3pa6zN1K07rx+IOFVdMIjialTtiixGyijGgKE7ManSK3WEhl6MOYGOwbC7uN
jtSwrM3ZtheB/UeWlwip3ZS9A1IQ1EFcwCdySxvtxK3OSltelVaB/9ZYu64Qw/xu
VzZslX1PEqh8iysXJHURiBkgVX6E3LA9CZJkepZHt+MYm30mn/KzTGMMrwWAxQYF
gZKjAK5UbvhV7lcqFrz2sMhfM90TS1xLosDL/CoOaHkzKj4dk8OP9pgpd+V6SQxt
5zGOqzIFLIKdz84hziWBfngoB6JrCkqR+K65FU2M6S00Wtu2vjcR2nM5NZnTley/
LqfQk2BTEqPGO9UENI7mGYzQgT7/Rkbt0zLr+V8iRiGBNmKqD9Mog7k61LMBJuJI
joa/sFG3RozxGTTOJfWwibg32h/ulMQONGa30aPkuyZYjb8VJ6mNb/lI6QE3jcJa
FvynjQBpN9GlI9IIOI2nicNHzSKIysTO689KI7D9AOw63IE2T21jcSFMQbxOYMXX
WLW13j6IcQMjdTV2BKJulmI9a9E41MzfDno0veM/vzpQq7Vd27KT8997xVoTsDza
YFqeZ9JN5+paB8oxHRp5qv/Fu7FM8PfcyWh46F8a9Qt9J+p6mQWRQfQJrprNYEZH
wtUiYNNUIciVhSkTLMwRj/BauX0OG4KvEbe5zv0aAcTanXHEUBUo5j3mS4neKxTP
wy6az/39PElnT4tfpD8KXhC3jP4+TT/e4RFKPJNPqFvPmfKcTgWb8JpxAixkJKFV
xUYRSaO7wXIFsIcb1aGCWku6KauFAeIFb6w1ki9pJqf4xVvTvA4vmyLZNjSsvEX4
9zZ/3IrB+Wbw2vQgLHfN4vMKdjqHItM2hyaujr2uAQ+CNM6Vn7sDPJ1TBuvbYE3s
BwEfR6v2aMqHfPxayFng/0O4dVCPZMFMfDRJo+93PIUSiLM9HeTrbdrqnwvC1WIG
z1Iifa/hTbpPwciMNEqY24D0Em0NVVsaSsledd657JbER0gCxpUqbChaNpcr1Qp9
fDc80gsilAAIioxgWwB49wu+aY0u6cl1j+ILClHyzVxurwGSNBYfW2ZH56g9ilh5
LUNHmB3E30AoizEAWJLIJ3daSoV6e2KDRSju6PdhT+4sF+FSrPYr+qz0Smx754hx
Es2re5F8je0234tfVbckncAKFNZVdY++26N1aJ15jfudLl/rVIldwisIFPKixsKk
KRZzTKDirQSeKzmAm+3g8/A/3Mv/FH+WcTqwNc3ADwKFWwsfnkUaNAAEIv7qlKG7
AuQF2C34LjPzCxN2K2OxIa1xKammjBraJd8RHgmjIjGxNKJeTKQng1OwbHHV88sC
HNo0NipARmF5uafLBQ0inEk7n6VAhTtIyOs9qg3Iyqf8CgXtu5BOwngViA2Wy9X2
f6MnhzAFbpgCh0eT6oxbeh2d9JUhqzEa5ThSfAa1EZNiXkOIYQAY5KhH5xxEip1m
LPN58r9dAFwniU+GCdPkZXZ1h8Zyu9FsRnVGxEJXcQznl9GxDBvP2Oij7YMq0WsF
VUDXG7ZPz/eSFYxZ3EodPGDXAuMnWE/7f+VyDTnLaybkb4FFR9WZmiKb5aq2ifbt
NpEFkIpc2I2G0BftXPF+xCkiUv/EH9mJgU3mzvDZ24jH6mUn6DhbwZFXpeRFVg5x
k0RL1hx7ArPZ7vdgBjlWdnKUT43bMlpwkhxVKkPHhKbOKLC/7m48vTtyeFKwttDq
6GSXS7U5mkh82I0ZcPF8AOMGY15BQ7zOqjvP6DpLGFmx+idaTf0ywMVRqTc6+EFH
wK1/SotIKX0QqxlZmk50tXzfLv4irzce5p1UAe3B0REUTSRKSd/ne+T13VadUH1/
p4kZNUBVZpRw8FBiRSg6oI5jU7MHdaVUMepm5FuB1i/LyeMLv4LFSPUrLtNX8kZd
0DCQyp2MxSr6S8FvS1EVIHGxLEGSvDDuC/qZXkiQr8GMUdAmRtMIJsanGLfQftH8
GP4DORcEhzX31peROMFbqBX0Zur3Q02WpFmj/GKHyD3qNdjX3ORNXspstZfYFQW0
zbs6iRf+FU45YoH/OgPUC46/Sw3FOkpt2UpRofuOtsb7EuH5T4tSFHEo0u3kS5ct
pRVW5OfgncSDcAYgWpn510eDUxcSrwCpaFgcj67TS8kAE7KApD0J3Lux3Ho+04hY
w54/DiOa0Mf1h3s3/DPtB9wtl/d8rwbxvEgUO1iuXTVwON0kpndpwVJ3EBeNW1Ig
1doT0xcksuvYVBhfTg2RB0alTKPzX5OSbm5yn9OeKXGNQOQDY15CQr/05jv8vRxE
gRYLhO1Qgs0Tf/3X54lXUgNWVqjAjW1y6yFsZ/uOmrYGeVQ+qCpRZjWTiRYCRm8T
tBrTntMWdsm5wQyXb7f6xq3uvDSt7lRTeSBjhYERaz8ARXyMFHmJMOdRe21mybYD
Wyk6QoRRNGtt5zSRhXotacKVVFa+T6Kt/0fTv4bGc9nd9UgaBlky6pae2bGw2Dal
ANQmb0jBiDDd6CTEUvAfJzhwUXiMTgfrVaORUGVR/1dqARhZf3uPx9eoXbwXzHvF
m8CzCd5kq+/2ojCuqJ64SJuuncZ09i7yzlw4TL98wIOntaa2VUQE6u8QhdV6NOWl
CoOfYuLqTLoC4HSA/ueDqAmzwvKtwO5IsXkkFRJduQNzLFpzvy7oKAb+qL4BovP6
odadqB1rt5CBjt0vufpeX+OksJrm3MQeJ9xfZMcg+cyFhOpYBLUNzWauwEFPNMYm
MdGYRmYhfiiBuAjeqQDYIxulihrSdme0pWOJI8oh9229P4dZvBxEJoj1xz3JT/v/
R0/0c5w9OFzREgCBjgHYsgAiXFvNMDKTQe9YtDBVOc42fu728+OgjSVkC59kDbMB
teuVjj3OnMJByGsE4wNZYWubJh4nojuxc4nAtlp+8lnI+e+550bZODvZ/1VHibKR
ENYEb6XNlZHF9hFK9RSTJq38sPVzWU8nufJthsL1ETP5s0eNrW1Zver/Zl1+/fhh
VlEOlKnUAOx3N6u6jXs0sTIuroExcev0NptJ3Ool/FeQv2D30ufrcdusjURdP1EH
bNF/mVbKip7WT+1Gu3qBhWm908TkaM7xYRyV06lMiimNBGTm4YdA2nwyaT5RYqP1
MCRZ2WVJxm32LxlVWhE/k7HAzFIseZlv8nM0uAn/0glqOXz1FXtBIgM5SfdC3Xl8
i1PSbm0rjbT1TFnDEHy1/5IjotMtIOF88L8YTq1Qpc+Lpluneo5RUtjTCJPs5sV0
dbt6Du4a2j6RG4UtrkivHecMXoce8I2QhpH8dvaI6zKC0YXaYbF67qL9IuRqaoov
oaaSsGQeur8LIThVRxsxj8jB+atAPsmdMa0KxMe5hfrdLoLYthKt5rOI3/CiXFwh
HKw5O2agEV8Dh5DOKct/oLWcbRA/rz14CWnDq+DeqaCZUk5oCso9vBgu/1MaQjLW
33VwPZnodiJ+J6QEqfMC+fKdFwdOFqn96KwhhopkSpjpn972THx5pZi5VOu0lf0c
yE6ww09xgujUmlhX32hL5jRi54WYDIFc09uM3IIbWOXEdBUGuW5KqmIO5zXRIgrD
d4LBVpvrVqc+ppZo9hHNWt2Bu/R3t5K1cMxNEftXN2H8ie3XM+Rh98bI+XGgkmz2
Z2ZRx5cWsJaTZxeAn8ksqLA502v+cLOmjpELkcKvCzsFPfiD4YmHF0O/5cWFpzIz
q5ya7QnmmsITIMiTKZa13zcGcnoH+TSHoFWMQqhJMMrkmQvrKJ5IqEkdSMcy9NmW
Eh/4cZQwpbzLMdt5tu9wq/6NkwHRjGf8YEXHETlz7cNsaPHMrsb8n4LEDhSiMxXR
/M68KAnyN0YH9KYaMXtetQlJ83lRNWpeUTKPj4VeW8P/D5nt3porsuzWZ7rxtBsj
3Dwac6WEUwMbz4UCYAwKNeSnsAbLb0l5/82W596quyr6VOn2D/fF8MHgji8FllV7
GOKwDJnNfDIx5aw+WGX/AfLspqcHZjFxddmg1Y4YeGtgusvzbYwAc3fQjb5y+cTK
GwIHiWJZSdbqf0klMjCPb45/JtuU8v9hzfkp1A/On1Jw8pHNXc6XY6YbIA9WACPw
5al5hXqXnDip02/8Fjvqjw1M0/fhWBgFgA48rXKQSo1DuNMKuw23uTOuqqQ7dKj3
yRRbQE09E0YxvXm5xuOLPiFDnxQymcLt+GYm7wu2pOCYms0qLrULRGzEjAoYdmxH
KrVV7SbOV7fdQcUYQMd4rZmbA7gnJJF7Lt1SFvhEOzPr9Q+btsHovQ/WNXUUBTse
2eh5eWVH1k6uacavCxMGvq7dxx+PDB3fKPUf9n3CSVJa90qGQqq4aJH3eJQRRb/g
F4uo4ACCfdowHLP77aScQUP3ZpxPslEEk04sfGXKvDTsCNyiJJMxOZhCKDLSfwGx
tIWRPOPBj6yAjcgW/s8VHl36tDBQt/tTXenW0rTjAL7XHjHncT4A8Sk7MNbcRlSV
POKvBN8OLHWJ6/GgTlKQ5jwdJxj3izoGFsjCKUZoVxWDP4s647OhKEhn3p1T3Hjd
8iPZqLAefpmwLIFCtgeGyAkitIS/lcmxElyURwB81aTnkKK27VWEStFwnuna+tPt
BkusIrCFJ5d4fyDD2/+qZgrjpODBCO/ss1rre43r9nCv0zajT3pkd7NwhnDc6cyd
xXVK95F+PTVpGNExvYNeU3pTUm0TsgtmitIbUM1+Sd6VhxjjrxEafbAvYuOEzp3X
mLvWv8dbF5Zb6WZF4VZyjLoi3X0WsJQlnD/kiWypwV34IslpFlpCQDO7H30vk+cp
4LlvR1eC/u7w/D7WULuo23lYkqEe8v/H9DYYQslAk9sXIjLFSMSHGVYrQ4HIzX6Q
F0F3BobZyQFcAnFOimFAshshNDih7AMfCAPRKZ3EgTGa9qGxIah8Nb3WcGrHc42h
6xHNLTtvGWKm/jZDginoiFDrbR69t3uNWJKvh4O3ds6rA4lJqomtRSZqAS5cibbV
JBdakeS1OnP0sW+ou4z/asm8LoX5fwn/v7TZ5pfxo0+7q7QhJlNHqdpxFmjz9Yzc
NYlMUsFMXshKAXq7YP6j1PlRtN0ae2jo/XZppj0GF2k4gi5Pz5FEG617/dkwjkeR
Oc4Z5O3oAMUOpG47MjoHgkzku0PajbvJrXFjvkPLV87GK/kUU+dCXl0b9jSGOxvG
d1bo83x8+5XZ0KglQX6Hb562Xbi9Uv9BDybligegdq6SH/vLEYFPZchbMM+fQDSH
tq28/tzSPGvykQ7u8ynTHFERE/QgveO4fvfUVXjRASlHiBLXXOQM6t703+DpuHs7
ltv0Bm+JYh9eemleJqFLHDYtZu3RJSyDtMNBje158UKemLG89XHyWjLQwax6dNPr
sItpHwzMvDINlphOdXadhuFaVTouF82dJm6e7mahSRkTjerenH2dOB4v5zcm4Dvs
STGw19U1hj5hptSIxXwmRFULfB5CqsG0rnmepI3nvzdMre0QT0M5MiDgbM2bkcut
H+D3OfTpjnllhfXBCykTWDlZLZA033QGkvHpD6sr0rk3KRwn/zfiKI4sfxUjqloi
5iZ5tS7vIfjGRiSTU7FtGcb0ZB/KL9djbZya7f5ra3oFVvCEgb4PW5bBZ0j2+W+z
/x0/hLkQ8Pq5iH2mOolyl8Mf3OUKl1/kEdD1JPP26qi6BLuLs7mEXoQgVqC7lAYY
npde16Bdd3vksAEEgerYwkHoRVwZ+lLfIgTQnkCDxDZOqKVCtST/HW0kR6hkzpLn
uOpLfMOSXIvOUahPsurRuD3zMhYbUm07MhAIIpQPjQDBoC/3Fg2q3rsytRP/oozk
NDHi8XD3N+56ihGe7NLPrhN6pwzDPKOQzWvZ/NDcMvSJAz6d+oPt/P9MGuUVvck4
RXNJyA5dN2oul6jjWWQDF87rzzU0CtVKMDi9O2QS0AeYEGS4WR+JhW6RUbQIOiRq
ZPakNp6ly7gS2jlJ/dYzi7HYkf2vtpxGT4eDEiA/k0ChbEyyhS/Szsvxf3yI1m9R
cC6y7wvPsUNVXLHV+RbZ/P0HqnrehiRElVXB4id1KcoYaTK/lCzSdknMBymw0x6+
Y0Ct2HCs8WFf35wo6iyUCSKwtoIwoLvak35Q8S906Y31/h7jFzqohwKNI0ydmBJa
5qCneT604UMidy3yxrfK2ggME0FnnIbPZNC3oQ7metQVHqtvPboCXI77vneR2xqf
YLeYH9DVd4hHOlYrNhCo9Guki+8fGuJWLoPb1K//f3So6Bq/r0c0b3VfH0kg7azu
ZV4Bk6SMV16KhEfw6cmuqzWCEcwJTxJu12Jcco23khSZNpBnRrwnD1SNTbgShBGQ
78+f51l7v+hLv72muPZRBKkUVUngWK0773j1aK2LF9cmZKGzHLaU2fSfo/5ospMZ
tMwAHn5YN1N2MQNl5rP+QArtDgwhMTEhjfU0OSHTqPK3PZSXnb+oqQiKpYr67+c6
TXA/URBJjqmjFvzuPZPORu0S8FvHShD0+86vqeFkd3Pv4kw5/GRULuTLGZrq6fKU
7Z+/aTUbZnyKCm8B3Etaab4+dSHiAFDo6kmAZLkIlASQnlJOhIIh9xyFtrW5Bcqi
tzwrTjayTmztAdY8fhwTknw+Xk9qu33iGH8RFH8bVhmlP8dcuV71BEU7wMKA78U+
S5BSu5qNCB1v2SsR0/XlpRHTr23UsivKRIIog8GjDu9vWUP8FuRUL6gCx4IHbpLB
e56Si0j0elmd80i9fx2d/D2QMrrtb6ljvSpU7b13jxIj66FbNlsUEUmhYTBO441/
RNoONqL7V9607cXtQYbkt1VWfyLdo/gLdvjE5nS8f4q5V4XzCCu7OFjSmYrVAYiF
g31jnEqgLGPYYyva/lUmhQlwv2IqK+LCITGS/IqneRurYEtM8mecAq7VxZvTRZT9
EYo07fmu1/kcEjTII8aG+Scf0TS0b4V+a7m5zPNIvD7TUiWoeZyl60mhfqzwXvZb
ZnbaTmjc4awo0c1xHfd4Vv4d0oSKHgqSZEIsNhqvOq+IhboJqc4a0XjDQmzm7ZpN
UAtSHQyUKPD5NVGso+c9KWkOfJoakEHQpUrEpoyi4kz+1AKhZLhmAFlWclLcad49
lttMSXKjm9DShOQcWfdCSxSDNkA0S8Mya2AxZVX+vTnfUFpL0366r+OEPSlYA6AX
Z8EJ4par3TBDI0rrVz89pW89GeVPPdFGV0OJfERiHQAPGGbr/EeH2WCVWeRxoEMK
T77CvH3dPrThDSbYF9ULeXip8gop9G7wqiR2bjs8hsa78x3Wf2BVHjA9L7yAEUbP
dXC/QyqhbauecOvY0eYhbQ+vsm6i9Koim6voaPGqECQi6qmyVPOYhvs5II9vGfTU
E4Nb3rtGamSn/potEHe/F14oBDncMxDOssIwSxfWjhk1qhEvNjnXHsBT7WkZXDt9
wUOdx3zU8Z2frjw2kqq3EG0ginuCoNu5270wzYapjNWyP6KQbSqBe+4HF49xMI2s
xR6xrifQzpUJMKh9el3drkrkfJnYwr7sYZJG2IAcP6C769T6O/i+8AkPvdkWruGg
ktxBFh00jhpgR8qrjYgn3F5rsAZ/5M7CE1gPIvZ90knVpV7CKgCE/MuxFlFrFxno
R7jHvmEgxYrXsvmrFeKxizW8ZdQ7lYVh+HGfDAS3/MTWRYL33eq4s9zx2xUfw3ln
S9RD1PcXZgGXNVprUg9/84qgqk/ocQ/o8CTuC3Ybf+BQcZqKXI8c14h5Cs0ZVaeI
n+SDzO0mjLgHmhEYff0NUd0WrMdwttj6QgOsq1OHSQSJPW+L+S2ja+9Rg5w6PcHK
iVzlu8xhcXeOaJmmWeTQBiO6VXYtmZqZdYhr8vQFPXmdjZmSbqZg/bSPc7ucw61S
kkneY8MT8+D5v8K75bnwWw/n1E++ecA+j0nMMQ1lAaDyTXCdkcfE53ZIlozmL6Au
Zu/quf8mFsZ7m7xtjsouaoPEu/WIc0I8ZyOOYlTO1+gWZlCOeVgJ/NFSn93iVyuf
1vgWB4cKyMAKNijpRnsSCIG5CHy+hpQjQRyhAYlhvzKwAAtjjdSgkqyZFITIbF+F
S5U45NgGcbpuEB0MMWU2zpkLdu6/BUL6IYaraNZkKplkMq4WuMEGUwpexpAR2/NP
HPAgFahDXmLWePhjZ/O/3ZD0ajJXngkqHTN/RIfIKnq6o3dGQUZu9EUe0AgVSXYt
WjDrvuaY2gVzGpaiXj2a1l6BTZ16yGR31YBWyxA9fpqrvY+RDWXfJOPMfwL2m4Pj
GdoxGsMArqNXiaN3qL3ladDPCR9lh3momQ7UtOHeUhmVsIZs1LhV0snjLxpmgWvH
67B6FYir9mom4R8RAQ67yXOkHiXW1uICu45jXq+SMNWj/RJyi6eaGlqNlkijBVrK
htgfsdTHpchnqH+SO4P/gzJ4DSTUN0QQLP/WDe3aqwYxMJH22hpRwKxz0MoKitk5
cJQdTbhKnnQ3JupJQCKbwS6AjvzPsSzXKSrSJiu10Ra7kJzwTxeTgP3IoyJ54kcV
hwxk/Yu2LH/4clEp6E7E2dkwjW2iPG0+LFdEvoK7m+38xoxypyuo0KQMq1ZoMoG7
ZSxJusS45Magv55Hu0n9KbBLZLEfKwytcuPx1LEs1vwAc6Dw64NiOYDU6damxJ7U
dRaqNzMFINX5sPRWKdGu/G1PT2y8Ffatw8W9/Sf+SqV8Nu0rtyUjS+bKajFl93UD
UZ2BcbUZidOpz6AM6EOE/fN9tc/SR5mfh2Ntr37JhMPVVTg5UfDxS+XHBw8sqgVj
81kH6ix+6Htwlc8oqKhvfdkuibuO78Pcgo1i/ksxrCOjBIcPGOi7bZUOK6cTuBF4
/QtueKjOd+0FGY4kCMndAAROsvoHQLF1D8V2ltePuS1vKV4evx63iVMO02pAPfx2
ijW+6Xtvq+eTD2j31whPEOxH2wX+9FVt8k6m0EHmv4upJtQMy7yOTj8wxen3KcVe
sXVAU943SYuP5JMF8cuOg4JoR3vkqsJwV363dRxZpby0uY5P6fSGV1gbWok8HUAr
8ca1JlSWN+BdopQh96jDh1/7oAiJF6oD02ilG2NTMkrJtfKZ3Be4A4U1URdxNr1s
fZoC584ncHPujNayEzX1JaubesrcAnfzwViM2pONCmy2DDcQBogN8mN+GzXgGw/K
Qbolpq+0XLrqKgus9MLUKVyv6LmA132Liy6Hxo6AYMhZG4MOZWwxWDcuJ+qSNeoU
H2KaXJHwjVjrsf42mUhoe1irVfYLkSJGj85hN7Ff6TxM7bw17XG3R+cn5Ed73R9f
egebT/N1Zea8sfNFBbUnY9hk5wv3sOFnMcFjePT45+cF9vuLM7P2TmgICm02QR6B
mxR0woTyjGibd1fEE65EA1JBQqtQzeZ4tmZ1ly3WNGGcby4AXwYJIlbGUgj3/Pc+
i7aB/0hCvdwOUIAtQTKDWJN61T2VmJCeI4LYcoZn9GX6evrjPFwhe6S8dBO/RZG0
6GuKJmYZ86+8ewECrOvC9Gztnllg/WaSS70gQnwLr+jEeZpuWJMf+ugyuw+COpik
TUqzRJ+Qe535/78DZSeNcUsUv0/j37ndLZqNL4fL4ebvZxnNW8Sg6uzwqwTMBWMd
rXHl0ZRG+6I4FcMFr0A7M5YJF7+eSIIaADXabScRDXTPg/Xqt3cG03cPPpV2cUMH
l6QjWIgaxD96pSAmmNUmAdc5ntVSyI1cUSn/p6WCwi7RWuXZi05PzmZ2mF2cP00i
kwxw0rLE+oRJHFF713ut2ocss+RxAquIlxRGip1WPC9ujYHXkob7PUbzW1FJzUYG
gmDO2xq4xJWeuCYrO7QG3kmOD6mRC8LNaavvLasqYLMFK0i3ov1HyB3fgD+hG6KQ
PXEh/qTaH1kmkZFWCZa08dVtwBFF9dcceX78N1uOsaSzE8s5PkHyprHkSOsdqGlW
dTqg6wqszXmeuwiKiDeUzDXAELK4Q1mvhZ+RiXIIL8KH4hAsWe6K+/YrlYSpSdap
Oyqk0W3u/u6JfaFgv3YADLy+wpY7IozPoHvqs2d55zKZngMBoO7Pd0L8mu2he1rA
3xDakgiLY04Z0LXRzmi3ov6FGPHpUoeAfyjEh0vOWCZkhik2ZJ3EdMXsqDZVnUnG
pRFeH2UJG2rk6b2gueqljZ8YvadavsVTLZV7FYZHQ98fKYUWAgWtXX3eH1BlwwuV
vIhXlE96s5rUa2FF0le1nMYTL1MRmardPEMNoyOZLJwQ+JcAfciJoUs1f8IEmXWD
Fhq4+xYrPQxVcIt+gu7RORTTcOyL4V3Q/6cpvUl1rZ7k94dxYyIqegVgdb33N22r
ytynYCxygd8dIZXL5/kzGI3XSfH5GxzR2tTrj7JHE6gjZqP+lYqmLi+ZwjbBHvaG
o12hbKFFzZ332X/foh4zJmH/h7oeHtW/Ao/XT+w5pse5NDd5y8XlfJFKXmG8Xfim
nM64mNSsMPrXvaszWL27GfJkDajltUa84a41vDXgrdyZjybdnHCg/thWM3yA1A6z
grohXrP3GK8nBCZR/DwvMrLWvqLRl0WLznL3eTiTyGdHoWkcF6Qc7I/mc3aL/wrs
KTJM5FV2F7RTOTWzfTLqHenAfcSAnNcIGnCyoEupJpM9PAxseECbWIAN9ti8vlpm
83yL1EIfC0vAWI+0xJ8t8989Ofl5pvMZ8dAJMqo3r15pBuybdIaTgKlXcCaw6WPE
8jqWUacBs4ESpHMRTAgS/XxSgHQJ4Ud7xFUcY+KW9N5d0gIGGT3i7Xi4PxWl1ur3
iXj7QwFauybzgSACiW2vWj9+SqyTi3uCUaQUqO2POqDVsH02x0bsBEi4tg0yxkvx
KOptRouuwUV8mWFXuLIad7JUfPXCaAkXe/9Z1aPwi8fd9nZt3ZY+xjEmkJyecde8
oft6eP6zfL+9stO0Kf/shFOT5ai71hvGyZEaNqdLVDWun5zYyOqcGDSjUzGJZAOV
7Q8iIqjtce0+dVsYeQF46RoSNER4f4eOO/93vHjLAHPBsNcosI9GKNzCSSpTtmfN
wIe2FOmqCEdbkUDq6I5IQhlAXoCQdCLhNRBtGLLrjLzqqobzRV0ld8VlHlX3nVwf
dtAHrQYTdDP8fkO6YPXb5tHkex5d/J5Ng1FgqfxK+IBiVbbAaA5r4qkFXdhrTvnH
TkHNORga68ybDVXJNRg4NJ+9zZ8JbfWiiLMeAjfofXZzyP+CBmkFCYpyJ61lhszv
Rus/XmkN2JVs2scycF3ACd9Xu0OIJplRzDag/+jj4uKuedDwgahk/vv8UJH/0o6e
fDMy8TyZa98xfzsVhXxhOfCuA51WmsxEGzvZZ4WVDJJ+KDQxWe3DjAdlollsp81Y
aNeBRYKN1wXUTuVDzE2I4Gv0g9q14FbqaodG/+2adVGMs0sli289c/SmUNmFzB3n
++uy7drSZmC4QO01vPembVVdiNUVJ62cV86I53deFyaIqKD5tXxM/Oev03b97qOM
B96DVs7Xl/V4AIld4NUntynvHkc0fHtFuZzYiuqHkF9uGNhOKjFULc4Xyod5BInQ
RP7ncntbvxYb2HgbNpxQuQsc+OuapSMQQF/Kn5eip0gVKYtEmK1nvaRJAW4ZkD0V
55tF4f6VGrr+bjcWelDUyWodLqFLyYVrx6rga70q3UpRE0OkFBRY879ceDrYpcpC
BcqZ+EmireDed4sOXVmSSZT80DRxegUkZkUsQ0Pbz0y0vXt+XHBGe9D8HJ1hyKKW
L8oX9Zh5gNzKTAhvvz/+P9SONchkqPYwxLVwJ2f4i3PbNyKQm7bJOT4d1A6lNog5
kYpQnCqK3d1xVniZYInbOJuvgxFoMlPT0JViAa7PpLeo3igVMdXi86U1eilc74F4
kvTeUU0L2OWUSb11BomSV/5jqumBQ1afrB29qvqxUtimYekHBtU4fO6bKwUZh2cQ
O8T3T/HDXvkSXNwipZERz4vqUexQey/iWEbkgyq9QwdN2QZKNZlTUbmn5D1PlYk4
rK/60r711zUnOl3+6XWZHYJv2EGrQcgbCEgWZYwjXck0aAAmJKCLQosB9SeDJxgo
cIEnJyrX13JxCTNU6CS/ZElTR109PBKWSVz/8YFo2qv/jPWakV3mClOFssf1K9gH
6p2GEt6Saa1wa+u/d/VEE84WYea9zBHbFtRzDjGg383mDfAfO0Ybh2pJ/aibr8qs
DUbvj+T0wDVeuBZQcmAyW/7TS2gnK/cFXBrt5THd7xkE1wKMNpxIWv0+eng4Cn2u
dnWVst9bK21uZiX1j19LJXJTHsDaUC9+TmwiQHvWU9/10AA1Tv0M7poi/Oy8MqGQ
K/1jb4RTkr1WQvDBAyvv6G68kFVTHckGXpV5SyPyAyS/zi3Bwny6o2Sc/WWIADgE
IovGzeQJQtVhxxLHa2bv6lxjfoy3iMfOGKKX/xSqJfOJBGE84c9dM0PPcCozXbl/
jK/qzWq06zsCusr5lodm0koWKi3ctGAHoJxoQeVJXNXSvqHs4em2L36a5I6o9YiP
B5L9YhUMgvWUPxGm0r4aMwd9JGLUypbTUawrHyBQsFP4VtBh3LZvYltGfKG8PzCj
TDtjCdLG9GJCM+O5LrBegWiSPcqrVKfStUOVlRKINJA7cYkJWnEPhW+K515c7NTr
XMhk63yuCdFEC7a0K8YnmWwxp2+PjfIRqrhX/exUi3eUvl0+Ra7Iux9dzVGJOYia
ccljl1PWLiek2/4kr08iHBhhSSwHHfQV0b4JYYOH/oSUh/5H+tHcIegOm0cU+Qfv
nObKCoibq3Txlge4+SFzryAM+TmdBSpkr1AvdPCr6fTOdj0ATp1zjy6ki+QV3USq
frKWUPzYy0KLYKPZ9LlJVd+6L1zZ9I0BZZfoThyCk7dH22CdFIO0g3jGZt18GMUv
TW6umJDULoZ9uWA0zvA8D4mL73XBlboO+OZv9uujnXSgaywxAA1ay71O4Gi/3Ynl
jIe2L9HonlN3xCQeac+cFD4em3ggS1vR4ypkOHRz64qbD54tWAzXOQp4U0H7crDs
79aUD0uRiXvAa7tQOJSdb7A9U4reYZlZ1QuvrtEpXMSIkDHJcDIHY38v8sh04qIA
AXiTs7It7L1Z81xLHobgcTv3UMK0zm6BaTjFJ4oC92mctXz3PrH5j8fQsGwR1MYh
UXbxUYLTYXWvwZh5BPOw2uFfJ4y1C6NJRIKYnYm8G+Y4rwW6jBvuoiGAbHKqrvSV
MKioqUcTHBovC9HcwJqIqdhFn31x16O+XQHcxV8CddX/ASolfOOowwVCIx9XGcVY
V2GQBsmoDlprhz9Jet5n1hDkE8CA9pHDqgJFPlNPFtnQyOkLWRN2kkXHlxjVfnaj
gKdbwBgj6FA6KtqKirbTZC9ryC4jU5UO0trgabbM650AdMqdCaxJmCOQGs9doOEC
debyqWnKFwjd02LzDUrQWGIbv+7NyAmTJvg3HKJJkBDTD5GnA/x+6yXUDJ5W0Dh/
yqDoyVPtWE1qLlq/XM/cFFSGufVBE7owGcHwJn1p6Q0Oovpfi1MqjDdyQfTs1q1a
C4FoTF6DP4Puxcl3oE4t1aJ7DUFF16qNIUXguTZ57GM/hf6C0T//nd3njJuMyOdn
f4lPunpV5UwFNhRoMjOi4epuZUBNCvarWbQ8GTO0lcifh1IX79gQ3jLLlbIASqeu
1Rw3sG0e+dEcH2UohdvLuTa7hVIY40vO1+bL+Zu+bw2IrIfNhrENdmM3P/njIIT/
sKphXSPyECAVh44B0jyDLoUKO4Cti9L6/GpD4wVydwPUuF5dobs3rGq1i/mzMaOH
heFl9VEL2yAeqIZGPMwXW6JR1LVFnbwzWQDO7FTWKYfgEJaXoA9jycoGuikdi9C+
gLqlg5LSQJkJPd6O0dJq3UEPlCFxYbt+W+Hvdx/sOPHFORcpVy9xOEDnnLHpJYcI
QV1HPCoz2LF/b2tObb9R0BPJ+KbD6Llow6nRHW8aqz9WUZ7WrFK7dcxlgzG/Nb4q
UU04nDNhBrNX5YIYixgmro7ixfCoRZ2iLL6Uogqnd5mIiEwOHERu4NCQOkgf/cYq
nUa5r37PW6W9CGsPDYJFn/hT26eYwjJAZCtj0OuZOOvSxAan1Bivia9sPMYYd4iu
lMXS+z/8VA+XmmhP5DAdkSZ9h5ZwEwzBsyhjDonbLVD+UwLSc7KaILHtltrGV5dZ
oTrreIa32mdloEyX36uQXebb7nI3/UGtQRg21O6vc/+OX6H+gJDC1ySmxAvlNfi0
vmYvNzkLZJzVXbwWe3qy+/7Ljsi1OMr/c2BqCqPuyrYLjgcZUzgSG9Ctgnfp2GST
XbrsvBAxQ+wM66hcTztkuUa4JF61caNwitHGeU161/uDSAiZ+pb/T7f+0G2h3lOE
lo8KVSOrBhJ1ehDZDWBS/q7JEx6R5qVGFLWGtyI7CULiWYq8PtyfnFgmkRiqB8v9
Ni5IYUZuK5p8jBUqMSdLN7laUorJSNWhChUf8SLMlmGuWj5OLAZB6jGiD2Dyl1yf
ls2pOcRqiEvOx5vRqpynuO+2ppLi8pBkBgf8j4DDDiEPJHkpihDz/SUuCMxVmdDr
hJ7qqxohkzwQC5rnHMNh7KlOX9oWVwDFe3s0pz3sn2HuRLxGs2nQrCIpduNrR4YW
GpzLkK//AiRqd63pzMeDtGOhq9MhgEJI7LpgZm2cx60YOUC6HpZOGH1h91VSBl71
J2gfgghPIXVYNX4GwrLCifTGSEQJkqmDuwkrXuWw7hT/taCQW55SthRa7sYJwhLY
HOCBvdFJlg6jvhjG38WnnTjQmPumEPWV2k+5PWMyKkXshb0XMbGrBydywP7cNSiA
zOnlpBCcze/l0cKCB2JM+zsdkACqzkHy5o4Gld28DE7aLes59bXjJ9VpnKCklGuW
k1NN9zBBj2FlqjGhGnAzKnWR57NEKmb7o5npI9pxgRnUvPjdc09eMmFud+/0gSME
rZVH18YDSmps8zA4m1CrpGDcGeDcUOc3GZOXaDnJvFY+gin8IvwlXaM/b2fW4g/m
ZtAJWda9q9sKz1bld+RemKBc3r1jBcChWfnncTSbdEGpDTSyWvFMi5NnClANbzIN
Pu7gdsDjOvWWtkR/6YGfb9RPFZPTWtltk+fboIY9lmumkLJIw60+wooj9yLi2KXH
2LbeP5pwFmV9+NGAtxWRID6vF0YcsrMSfCCsodeywGMJnGnZCciDbXfCOLyoaMqD
eTDgeSF0mkth+fHHTAxCNUkv37bu7HLt9WIuPJ/xJ7pruf4f4luz0UyWAN5WBf2G
2mKRwVakIJJliwXyR752599PrT3Kv0PAX6g00kPS76CeTKoCHcJXxLS2I+kEn10G
kKK4Cv1zXhNgpiJUQODrIIqrIPTet4sAXLdXU5WRu12NzMDqs3T9dg22zBmGZ3FC
bD5mLg1ivHeFYDm4o3WoyU3C18FoKaCjRrur3B7JimowfXVuU2s1P43VtpRlrCwc
GHKXpQQHAs2So2zK7Ct6r6kXkqQCRt08zujrF9A4/60oFje5JYdolYDNJSnAfkQ8
O616LnmJWUSBI1eEjq6kEz3sXg5MX65RcD5PGXWi7ovFmuRJ39XrSApwwqIDj3DH
M/f6xap3W5LCJdhFB6qTCwXYRuHGi38sCZPbSBLs5vCI3uD9idlGAlYoUIslkzDW
vudk4PKEDEpEvxrQvoRJLhWoYGhgcflLSWZYfpZTNZOQk/RmAohtrqTLn+rzqLAc
h2tlMCz6s+CD0RTLEvkwcuJWBgPdad+gDUtfll8MsxaVLUJiA/0/W7TnjTxNXqei
js9aO7LgQRsj5sx93SXgq+EaUGOiX8i/Za+1uyhESgjjJmK9zPhL1QKiapN+pQyH
zveipMAXyrhZ3xrrIKxhtyFTvAFOIpE0sDIVwffLpHUiWpqGLTSg2jxil2RcsjHk
rWgXuw//o2ia2OgW7Mv8ij4qL1ihChBikA5u6hVbm7uD98xGpqLHanXY0cgREoCc
chJavi60JKV2JFMFawCu/txmAlTWLqLee5Dhri0YWCk/lOj2Bzho5D2FFez1n3iC
L4X23SkI2svWLgRnJ7lWLP4Mzf4q6qaMwqrTqS3m2eMcw0MfyTslhi5XYst+Cg6v
tbo8BD29EIQPN7oQgsjPvWVlE45TjAKFB5pIS25223qVBGhS2IVfjgsC1Yel2cXo
897+6wh/55+hhDQK/4DUxWyNdDNMPM646A+tR2L3dNIyV5FFym2neAru+PchNtn2
V2aFbu9eCVC5mivysd/U8hY6O6mIp9lv6kmDe5SsVXe4Gk74jgnXnrqeOFblYN8b
1DyXrmRJqPFdVXZVs45Qw562r58Al3/Sj+aZta23X50r50ZUd8JhETAD62SgxmAq
+NhM80Bzx0pijDQK7KXvMq+sX0VsCP89nhl+aFWBTvYkUtY4/HlCuWzFc3DkenYy
reDQflPQmZEC6XODLv779VG0uiP6/P5JVuA+CdFhrgYBfa+cP4VECW+URNTY7Ltf
EDlP3hzR0RJxVaRLo6QAA+0fUPhNrXhLh2EO9y1F+WnViAUJnTBgBowBo+K3LUJ3
ypODdeUtvzBaI5lywEBtW3vSMcwe9QRMyZydhVJ6IynU7m7lR4a5MJc5M62JZJPW
VwdVurPHHJLx+FkuN5SXbLlvgQET0ZfqDW0LChLvnK4m9qhnGCMJnogx8X8VH/Hz
FUa94Ti7a/ypgBKQAO3uyQqty1DxC3F/T6V/rmVN8TFyzRVFupb/lus+1+yTdei8
N8YvkgzwRx3kjzZYrGvBl+E6w4lbhKjjrH4L8zWx/Z7nmQq4orHw4x/Na34L8fUc
OFpEAmhiPY0YFAS9lE3bKrKYcUo7YuKJK7LR5b3iheecX9AgDpnGbG0Bk+kSk0mN
63SdRqjpG+SpwwgEg8Tk9Wsgg/eh8Wsbtnw26vTF36Pq3h7k1SJVjhd/FpwczeUm
xO2ZvUccohy+D09h9TKT/RSfNE2orPf7v//Mgj6ZbN+NX305ac3EzGSwlkIOEHn/
GzVlV0T/BDtGMlIpMMd1N4CzdoriH395vVVseY6lpsrjIMAaZoJJ4Ecj7za8cl3M
H876oRb/fIwSSfXmL/Of8xBDK043yb2yT0eLLyIC1JB0+H6fql63brJWEYL8WgD7
vrqYFgPHnwtAX8J3eMOhzhSDL7OQUBWQClN3kREHnDC4cIhZnYhO1+mKfx4TLrzH
/VfQ/Zn2+oT7UgRV9/ILIEWr6ih3AZOg2zYuBOsiVOv1Y1cCumqCReMKDoogdOGd
sfgDXACVaA8Hv/X476PvWzgS1IwX8O10VB/duuiI4qLKeicKr4TYIBKjoOO2qC0a
HtuENXLPpxcyM2QO/Wr6OBTmIqKbqxOnLt30uvWJa7PhtgGBKDhsNIyaRwYQ6yDc
t2MDUePnzwYzdPJencVTy8bhQJMwxaoj/e3doTTAAU7vunWqTaEe/xz20qBW2ON1
o7MfSoTQRUjoRTY1cjrrkHdRUIu/j8OlBADGcSnKeCmtp7oQ90jqr3xyi2fcuN6l
Aq13sKpIrhZzOHqMoP6bdVw8hIJ0u71mE2M6x/BZ0wYjCHT68qc08BBOSmXNdRCe
mx8w03gT2RWoCFcvBC6UfwMpAZr2W+BylEh5ZdnDV9uA6Z5XPu2KeKGVohR8El3h
29eWD7MwYyQ+k2teCvVDUX8guLYi4tSC05y9tZ5PzaGhvTEUksBk984qWlKmI4o7
y1c8HpINCHDPlj83xHzMPqedtrkCWZv9JwdHoN7p6CFMkNMhPORnXBMFk/Lnx4UX
Vs0duttmdbSRMNWIZObC02R2uODEOfPnvGpioeehnQwiYpcZPvLrqSfVA952PJcx
0T1/Nv2hq75tO7BnpI/p5G9Q1o3g83x9DJtidHaXSMrG/1SwCg/U4rFXW5VG2xRx
4guwoMW2GzKDsCcdm+IRfEqgMjTf3de6MSwRua56LdRl5OAZz9PyHcaYjQRH78ky
LB4Ukig1hLpsPEa9rpVo5h/gcOocr1FH9vQApzFM9zXNpCa+NmPRXwDObG17jk/8
iSh1nBSC4ijZYNXerreh9NU8ETYd2DC7qf3HW+soArPmPpE+8JMhdg6sOhzTbSf2
Wt4l1OnuGSEEV7wYB+R/Ja2ZRD70+sNY8mBhFfL6YCALqmPzp0JncVOm3OUZRyrF
dXN9UWguecV/nFWSZ56Ii57/VrXGcg7+zRfzX2w+uiSmGglFw6wcMkOQz94dYZKk
21cVUpGMAi2Lf3q5jSK2uCsrkOrQp3VCI50Vjx1XHbUNmyTJJaqSgZCH9LLoP7Lh
MrtC92md+oCNQ4AYDz/V1/Bu6QHHCYnU0PGZa333+u/UIhf/yVbUe9PalEPHwdZB
cbPuf4mkuawKFX/8xGmCXvjkik3egxpZSPubKh3lfRx40tRi/t9uEoz2KFX+mV1q
F8Wury1gKEjnjo4tgWugsjg8mEwakvZW+92umVnWIaHnCCShbRHW88wUifNdmjWt
ynPfOW+CyNzm25omeQpM1u4cs4PK7oAnhpoYViEZ1cdjmCR+pvo1IQqAAO8AE8k5
7GYoWabP6JolLgJtDgEuz19FnCqxco3a+IggArkgUaYKAQ4fs0/U00qEm7vOHFDp
updpj6d3BB2bfO4svgE9vgeJ7p6qkWO0frhmtgY9QUqeF2hOlV1p+NbR/Uoegwlk
cNQAB+pKazj5vzwkYLUC8jKCi8Ee7J9oyz9VNPNIL8jeCKQkXTiNRvYhRE9sf6NA
lgblCDKohvqQ4gufmO8qlJNMvPGt0d8SkVVS04J2Hef7UBKUTC5BUTqvxvinTH0m
ENXr0gTe4wKimQhUYyFLh61NKANj8zrd6SYjcRfNbzxEjVdfwEHT8EYBmcaBJIRN
oXapGE74flF8xOXaWQtQJQ==
`protect END_PROTECTED
