`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/zBSsBSUx3MPSnE90SAQibSTuIndIny1jNuYvAZeisKEm0PqO8HUnJu0ag7Ciql
LabFbbCx9Q7dKsphpRDJ+MOd7gOEec/xuvZXegpGzE7LWm59uDwIHrAMZNAjtqdr
sMKYpE3qeXho6MpFACzL1+jn9hXzjeedMIcmOjMF6U8Y819JaakH3yXonTDzWYFl
RJgYSAcxKEEa8pMMCTbl23zSHKgeB3rilaXT06ni5/7yE6TnH/a+TE8dlOsZP8B3
24L7H4+Hop/H/Quf6CI2HAlvsK+T9o8jMS6VBI2OMBGxz8sxTLosobL8qsJj5WXg
B7nxx7GEUrILwLOWqvaQfSEJvrQQ0dq3jTjhSM/eoG8sOdDeUdp+wK0QY/dBMIa9
0KiM2aVo7aLrC171rVcU/o2BWKpfGEzf5SG3UQg8ZEs=
`protect END_PROTECTED
