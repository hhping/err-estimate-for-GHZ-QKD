`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGcCXX4cZMXHwGthfetr6ezCwnDHwXjWfiaLySJ8/KAgQSZK0C78Ztnn7JIaAAXM
fsC4VLSHKIfwWJdaDQUIqd2L3YW3jnEnnKajH68LaJpruW6bujBoLv5wmI7cnCRi
dz+DrCdgS4HaHP14glHFvJ+8F1vF4EffUn8Cnp3v1PkSyTkssVkHtChGEWfxsr3z
Gtm1U07vqLRoKM0a1yxwXgNkH+12EYU+WEvFMTjVU5quvSovL2QYu3yLp9acg3ZQ
VPXv1F6x+Y5rRxjVSneHGF2rnP8+0qG5T82BQYGKU5LlM4kBIT4ISWVG0b3DYXpI
fkiLVdse2ob2ySCacoICLzJDitHvY3c9n2sUboN5X/qilC7O2dkhbHixbUjXGFKw
2ZvsifDVtYF3pTYkJqpTCObnvIMT8acOaACSAhb9s1wY0KEeWmJMX9627Z7Zqpah
IoAVn5hwDrkRd/qwv+/gKFqxZ0dlSKaklocof9qP47jf5HccxAwpawARTbmLBCu5
1bosd2dTtBCEfr2uUT/Xs5oxRQWcm21mVhsrZRcx7Mtu0eVhX+Orr8UJazOC2bUw
WZBZ2RfKyE1XpmxGJvqXjGE2YOdPhzLgM/UOnDJZhb5FIWS1mfR9H6vab9kJ71H9
D6euzZS/wx+Bb7j/Zhm7xrPZh/VvlTKbWRxJN6DZ3AONWi+1XuLx0SQf67EIcNOH
7ne8tuBC+RdjX8yRZChkhe51dX0s3+t2+Qw0mzrCh9xyea8v0kW4cSdiYPM6zg0V
vmzUlnwC5wWlv9j9t7DPAKJofJ1Ezsxu25iTlOnBVIPOJh6iBzDgJBa7nkwQQXTS
q3TaQnbEPd5XM19wPYzsTGxNwlSCu7nDuq2JToIBh0CMkIYZvfj7jI16yAAl47pB
/lO+0bw5Lms92uJI+Z/Ky8h8iK76LsNdOGE3G51pKm2/ggauJSuLn3QpXquunWvS
ZVH1W7BU3k7/XiHccR3amWCR2izFxFfCCVQ4j+1zLqN1x7utKopY54/aDWPvF+5F
47JhSQqK4OYIaSnvw/oRrk+vUYw58P5a3dyicYQiYDbFwKjLO6aIK1LDtflpyXO+
SdZailXT1nD4+knfc939I3Af/8g05uoqlCd9WNkDGxP3BssFs3iP7e32BVzJTU8C
dFpQw8RTF5pQkT4zey0B/uLxI6P0Ln2AJkjATugSNp7pS24DKuJQ7Bl8iU4Ic1LZ
VhxpFY262kkw+Ji//5uupd1lIv6F69u7yz1X//UTpsgAefhqpWwIvcs2gDp0L4/C
tWoRCLidTs6UfWGkpzn5jOhSEjBajg4N1Sc7qBg9ZvTScstCmTSX0X6BJNLA7Sqp
skiaWN3B0Th/9WM8OIXongx+0ZkjmLvMjiI6HhwoOLBw7rsh82/QScvjzQ92dEzF
uJ3TC17JuKxT6YE0aM4W7nWS+cZoXdd79zmLyJL3ZyKFGXgO1rzszGNXebXeZNGb
+PNohUVISuhrHzs3jBND2Br6QlBX3bsm9Snd7PzcA1b2i5tN3ttLy0USLrUfyoSq
gnHn298yc9LoCtKehif76xNnVzB1f12uEYJ3uOEVZA9jehIfwdxLMRMFtznxv4dP
D078K87x/aqr60HoyPvMW0L7wPkSxX+uDCtclX6dUmbRNPb2nOA+4at4eRGq3AAp
y+U3rekj5tAd2JGhUKBzjTrzLySsCGfA4xelFxaaUuQHXP0W9+dVDPo33C/Nhez3
7V/qbt8rQJ+hh3GYAUlvkxs+BUVQZAMvUI8D3yXvK/ajQ8Wcp43m6etI5PGvkhLj
OpI4+xbTDomIlWuNxwPs5v06+JwpG5bfeThupZj+r6HKnhI7Z941ehWh7StC/Gb3
33csGeDFpFyNehwX4gthGVdDxJrTpuJgzPiVRoqUKFKnQ75gsmi0eatNrn0LBoDJ
b1moAZ60WNd45YRTNe7QhzNln/x4nq7I/E9f2AooBx9wb9m+qvDgbsVhBSR3Cvso
KRxpJAUglplJqxzy/TUlXq9jO8H0bDD9gMQNs02wBjQBfXbjpTc48KZSP7ZCha+r
phMliNImpNue4UrUNqkIzsKhuvj6Z+gqxXrMT1TmmQM1kGxqabpdLpQA3Ni35oYq
vPuy3x99n1Mk7w0+onzQOa9aTsbwgTdNIQZuf1XZvJeGW4ModPApFz49vYQKlN9/
xw5anNqtt36Qw/Gs1gb5FPva+ZgTJnhh6vuQj231jnU2UkDg0fBTtD8Xts6UzeGC
aPD4azska/eUi7Tqi2UP6sqqcGjgVA7m2OV4tUjgBnyOq9PqFm6RwYBGduseERVU
WzlxflorUdcTEPV/rxIc143xQtxxa4fhX2pPnio9ZnqFO0lIII3qQUzGjIZONocv
o0GnCH9dbpJwGj+PxcMtqqNgj9iadlZ2x+uxkaCdo0NpgUYmXIqkjTCZkRko3aEu
Ad/X922DiWjVxWKDezYwnT5B6cxBdWPZBNccBnZ07RUOKJUMl5iQwB+26jKBFFA6
`protect END_PROTECTED
