library verilog;
use verilog.vl_types.all;
entity twentynm_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end twentynm_routing_wire;
