`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y9XjJP3ldFMM0f6zIXnzTS6suX++Gqtb+Jpn1IspWJPejDOWWx0RkIb/iahloS04
oYivOO3FTDD+6W5yDZgkpWIYUYfr02uMcQLLlZmq4QG7kVV0ItjZF2T1mN3ho369
bdwA1kEkOlWXXbU/CzjBXmHHBgUAvcaUbQjJ0ETXmQ0C+OH1NtD9lHU/LKyryRJ9
W6AnueZkYFkcG6+LM/YPd6ajGniYuX/lo2QYNj1y/mIjhFBE+Kh7MpRGQQ4J0wTn
Mn3D2ORXfjOppA/xqMGGlqNs5pTBQwWtOr4/iYP3IcUvGCxJnLGT4XNjp2aS4Dch
gq4fhcClfINHFJ6zUffzb9M7+Ao3GF1FjpV3+maU96fxUoHQstBboee5MAHs4fMu
H17pdSK28Edl6H9TYuX7JYQqYvu8k7XBi2fyzqLQCQE6Pc6nIKLsgHxAVKDzNw88
ZYvSO+bwd3mciT/zzp3axu30GDQBegVG48jePS2kPOObDOea2EPagq3bIL3QTncS
e+Ejub90bbCcJs1J4zIcHdcFDUtD1mkrfGEkQlDZlCDZMEl974NUB8q7dH55ggO1
N+4PB2xjXv7LwE20OR4IPquivE1mMOAjuPgBRgbSTGmiPw5/8mJ01uYUZDNxdHoa
lfklCI0A7KkAZqaXb42zICsGmHPOmrWQYEHVDPf6MqkUjtGJ5CrMQfQgZCPuuILu
riw+2UJXzY3fe7fmV4lMbKuiGRXyx6iy+PCXg5utWjgRf12caaJxL7q7lKomV6Gb
uPiAdphES1GX8wq5J+m3YagqPpTe0GlZHYDQNQfH0Q0yCRgK8bOtZNLJESuK2X18
IGXMF2nt8wYEtgW6sIu2MlL3AuzlfrbGDZ5FbOXdqhdRuAACIdZGZWY29A2eEVA9
VZkZ5YFuoSQhljA7PMzcR0qo1HOrJWyMaEuygrkRVKBULFLTnmhqfLgshPO782DB
1YNYKXOfPl0yBrDrT6OyCj4yiBj+INGcMcGA0nKnSgn/xmY8vALct/6l/fr+//KX
Fg92r1dSuS8iA3VhkCe1Ox4bNZjZeg10/uKDLvg27bXMLAizqg6HunwHQQwQfpm6
Kr2nNc4uhi3aDifNrUJo6OYECZKGe4GqR3yQaT+9jtJAjWluq5bTw88WtIJ2aDfQ
umVT+FIl1gmyvhTkgbskm6JZItpHlQlJWaQM9AdTfd5xGSwAQ1FDYFKp67gGwaVP
NxQLi8DBTI3Hgyo/kvhbRPQbp5Nc8NRWuBiKOm3xKlptoOBPfx93bz/M5LbBbw0n
sQFKHaqFgyK7BqSbYHM/q65/itLkzQfZGWeBC+yLo36MS33zJyJUoaMGRUXirL8/
lfGF0nueertAefSW1+Gpbx55YK/b+Q4X68j6L+s4IuRxOwb0xbAAJHoFq05wPSry
YoOU9ojguwc6040iqesMQCZTMTFhOS3+KMG8qVv/Hhvsaea5FxpLWqel3WU0hp7M
YTptnS6NWf58Q2VctjxihSq8/4k0KGe66s6Ap5QvZ+vLS7EQzLm3ZCYu4FX6+K9B
2LRLCcMDXf5iJy24fNvKywmRvMkCwBxZnhc5aYNIkjrKQi0dAYV1ktKXWOWgsrgv
dXeEHqkxSJL5Vslmcf17VF/9qqJTEfOWRqliC/r2BnUECT+ABmSSnNhWiKKiVuOL
KcVAo+Le7dJ0JsydzT4IbLcT11cDUiotc23zkALzgMal0JnRw2/03tr7OveT4ibe
eN6rZYpFki0pSi4jS9H6Ss5yyoAQK3iZSZA7QyZ0ypq9Th7/ySUPlr3o5VvLDYEo
LFP/FAa3V25grCUqIx2Bn9MzC0CFAObSkRVyZeMHnANbVAPtA/Vnd1ouftwJxqsv
UgFvMDmDwTWOc2wa9mTh5uw8YdJcY24iLwl/XfDrrPkxFHS7VvmSsachoFNCyx6c
NxSUXpQQpZgw45mWkwGMIyRRK3s8y2yPrfNRFS5ze0vnaKmrQivsjIqqiSBmkDLj
91eQuhEdClamfcemqL082jpsZqgjW3ogR3dkId00U5cbIujy4ff4Fjvqgd4R+byG
Q/lpfjmUTZcHYBB8Nc+ifCfo1udB9yr5aC79lDKV8U7qCmqCukjX4/pOzt7MBH83
fXKabWq3ydQCO15+ZB8xR+jt4Un0MagkxafuQXx88k6Ht2EFeelj3yAUdAYwg4am
7x8BLVuHq8g/tQzZ1+uX8h88uNkRgkpPiAJCGssaBnV5aSxjVlsy+9TxZk6qnYUh
a6PsZIbiPu3GwOxEDujhnn3ZL9BsgfZxu73+Gbh8u94HAVT57Tv4zwpadC+ffzeH
WeqVkSNO8uSIY5A1+cbsXgP8ccq0eaOKU4oRvq0sjAATQYfHWRrWUcfsjqmgW1qj
plYVHN+pwQneD3/yPPsbsI4fD62VXLij4LeAndFp/MczZnmEbZ0V3aEgcB3oNIjB
eZ86MmACET2pJfoBK5vb+DwzP8U2hVTwZVSSRRgiYWe/e36wd2rqHRxiX+qbwM7i
hZn5wP0s7Q0cVESLTGmB9J4OPis+fsV4loiY/gOUr+ADXjEZRgRqSOgEyiGXjCD1
zBG5gg8O+naFIWW76Yc4izAT2jKJbFONCZbDzlCl4Egjm/usF0RRm1tBSJCaHPNO
O2YR+Jq6+IjleDtsxgXoGiPC6sNIZySBHTObIbkTPaYqf4zJidMHt2J8S/YFAwI0
ZcFBfeETUihdhAVNJ0jOV/Ww7XZauTUNEBtdIW/RoCoSaqTqxf5zfRvK7iVfTq61
+GClq2/W1imRQQrziF+mmdB5lmVs5e5l2S0wEbZMOsKaD9BjqN7jTsNU8XSUDFYf
cCMzZ0Rz4IHtNw6warSWVw4Kl94+DYUo4Rgnr3V1ZzBikfkKnp8WzJNaTGzxmFYi
oiStp6615AH8VUE6q1K68NUbuzhOskBnB5HBJwoIH9eJJAqfcy35MiiZaIeDE033
1imDVw6rb29THyaFWrqqab+CuGmuHT1k3Jps5eEZ9Zj/7T4261Pp7pnb0ScvZ//4
1ZnKxkti49H2zNvhBQ2v1A0QjFijDefkBzOW7vVVvbGMQRDIk7g1tnd1VHm3yDhz
ueC+TJvDQ7VaGu80OjG0nJ1enVPy5A7NDtnndkBcCttzmLHZQBycJe3rsk9xFKC1
ac+sEIoYtgr8F9rGdbq3RGhPYS2gh4qFNi7sHncgUFHmEzKLUhuRb3cP6gyFMnX3
7tcA4PNQ7WWD7/ewXQoR8wYqro6hTgCDEasys1U3eKWd92kQS52a4X450b/azZyG
nLE9F+U5qjn6lQYmwigYQKRoNU+Vob0mRI89O5UEiX/xY1SrjIv+HS8Yj3HdhClw
mHQVdGwVMYvjXbrht5YW8LGU2Wk7KuJMNe0vyY7zWE/0PfhJdsjKG/GlFx26Td+x
n83K2w7aOMC7eiSbz5DsRkD/gExfFfWa0Xu25PFYVcR7/mEU2q9nfb+2RCh+ouhW
dIkmWCkiHjw0UcevhnKpHbST2+aJHK4sduNtOf6Q4EsAzfZZpxQljiZ1tbOMgpFN
WR6rhdALUgB6aENMXmX346ffVtXfm8IWDIFCfw6qXTlaOS77d50CTiPHh2MNo+R9
6jgmvK4fkFQLwPUhWY+gHvgSSFKwh5XzkUV59GGlT0e3g7mk8doHqxpuB/Vk91Km
MxOwbzsSYPG8hAdnl07XAyzsy/xiYxjAMd9FJamOukPL0XJnHbdLrlq8IC78cxxT
azT4lohL+6nnRsiy6eexXyghMa7swpJ7TA2HCZbyKU5HwTO0LFmAsB6X4SXnAO5M
NqRYkH7GmjUmnM1QxFDz2z1mMT6GphRUC6YS2s+hukV6VU2JJ9ViieWNwN1pILs+
gjuw727wBfTbtxnCqL86/q/DT6EOr3T6kmp6GaKxFpBd7K2mQWx3ChThVm/2vP0x
afmytJmARea3zeuUYYgXWTGo2hIMoY7151iQlsVpQRKPci1aT4t5cSboe+dFsufL
8yzCizwyF7A1PkB9sznJdXFSHz/Tgl0fJvNbUXM3m+zjJx7XA+yZncF0CnufH42x
BzIJnQuZHK8cdEtsa0kmO1ihFZG+uqAUeZDeXfncodgpCe04RQ+es7kUjI+D5Pxs
QrDjKhlKAQgH2ggaibVWah4ur6xlCwko3tEEARKxehWpqhWdU/fQrXfH8XumuM+3
zhk0TkWt2CdH4eT3lETJ8z7NoA39mWxq9TCvKJFAZEpzeg/WH0VgZ/rFizQ/F8NL
GEAcpLnbIQNamYZGFMtk13bukMuBu605DKNRssOR9zmliMdyQZKBJwVs6dWjb9G/
jLROMiZphMtg9ipr4GV4J+scUJ/JGXrsbI+CMO7B5rzVxAc1VASuVwwjwYx0Qt/e
jDNtAexuG9/bFUMovscc2uCOVEoHkySy5UW7w6HQPPtQuT00O/aQPPUHWM0UZpWw
+ZNohqw9Mwi3dn9qRXGJK8nZ51iwPNxtUwGxcfbFG3FWmtzjEH+HYnbCsRQF8j7k
CiGRxHLYMv0WnB20CAnTr27bd2o+XfRSIET5KCrFXFjOweE1mdDXAzllM1/q3ukd
ugn+NHMn6P2Os6WjEO0dSoq/iaE65OsQBHO0v4CEPAa4adGwQlR3xcoVB93dv/rK
wwufSl3FDVXaqruFlcaj/MqDiI/3itW/9GS3KLrnGj9ALC/gLgv6bagkB2ftWjcF
UznIjit487cF0TvrEJisal1zRA+EW2xl/PYZSNpQTmUp8ZnrAM23aD2qqHukC1tF
dC/uXcN+kbftZ3ttr3xaSSZ65IImz4PRQLxVBthX35/Gd7X9pCWCCdrJGqJeZDCA
ThblpjAQh7JOxj1GTxeW9DqhSymi0h55dK828R/uTUr+8uewX2CVK1taFjo3L5Tw
docTPgg8ZAIFS24peSQGXLVabt1bVNP6EnnaQVAFAlJ5bjt6iA2WSdbtBt82coCa
57rIut+jks1VDijZh/LrzlFEOdbbdC3J56iwgc6Rw7YvNBYtmZBq2JbrwDhLZ6qz
iZdifnR7PRiCSBYUv/vbuL4nB4EcT0CPMMoynvhIiNbUKu+tmjiStwigcsjtAatS
/FdosLdWXcNo2pIAM/t1hh1bE0m2XgdJcHdCFV4bsWB8eN7BkkauEmZIjRmamyM0
WmPpFOTAegsgl30YF5myeMAW6Ue8AobeqmoNUeVb8aoR5yv2B6dszGbNwiEtyzov
Ox/hSuzED0jczwsb0eVYurYb8G8Ss4D9sILvgUanwNDvAogme5xPehlJ7HmDL7IE
TtDzfOW4vuJ+TmdZNGTxo5ycxh1JtNxcbAgkFRtEJnRnuVh95fbeCHwOwOl55rgk
C2yo36OoIRzCIgWKPyvxpaHpkIAXA66sPMTV0ktvpf02g76FjsktQfIOQQ8bNpaQ
dFtcohgyWlEJWJna0bkv4zgKH/9hUoEPP5W6oibHtSLHJ49K6t7w2DblN8kAYm+R
gcuALl0Dkq6Rwx3rm3fN03B3LY+r6HQbcUkoKYKaUhKuU0H2TV7CL/X4pLLt1YpA
Km5ejXgVEgx0TvzqiZsRWbc7qhsBwh0+5gZACvC5jCkyFMMsg9jA0aqf4nk6rIh8
B9TXROsF4SAL5mzk2KRSflD4QxFryHOXVrraxd4r1IcnrW4VVbxAkVPoyDKe3jjV
KxY6SIdBNlkvM8+VdBarY6yX+kr3WVJMzJtOmKp9IxP2/82hKYRwc/eSx6OND9YY
4IKCcVSw0qmvcd2OVOXdwsKyUVrl4LoZyxX3+nPOgieLbVbzA0eTZMZiUKUWoN+w
I/RQ98KZACKz3rCoiO7g861VBYGe47sh2cMPKQvcustK6rAViaBNVjS1JIBodwx1
MIX6z1el4/JakD+9vhQkRuSzl+nVyKW9+SkrzQ/RbyvvrAsm0lwpNItdV+gaiRwv
ipdg0+7RvAXlkTPxosmbxBUGx23KMJiibWrzpkSmwTSHIH/Ct+Fbl2A7MrIQpIPw
PjOh5DcXRbAIktMM9A+izWHhzk8zpOOAGpBloRsCJawlsR+XxglrmgmqrjhChnve
+FMQG4OF1eF+4o0AMsFlpELkDLc96nVLi1bV1Uip5kwNYbupVO/ME3IGToAExhwU
ajMEc7kKaZmS+PBG49ufnFjo19apsui5Sa/akd2rACo3YGdrpjZAwJvQaknMXKPf
TMncBv7T1la8WMM4u7SKLyMxDG+gg33wy6ybvfs1V/dFYzA1lbsBwzzVWOHWcy0A
dUE4P2YU0aQaHE+1JqJ4HEKOsR0cARtNCS+PQ9OnPNmJcCNY8fKfZjRK7QV4GXXD
TwEj17gRmlgC5DAXSdSUzbvUnpp25X2rXJv3McMAI+EbHacykvM23BByYHTAK49M
+YirWu/Bf2nGRp6Q4jYNRgXonrQDRoVg581s0FG1YMtnJX6P3GnKjxGZZnYZ9KF3
GQxOeRMAZQl/xMTgO3CdQW18WjM8bcgll+oP8QcmQjohLVl6vcEbduczGZTgO7ao
KCBC2GsckyTYy6dsaUj5q9jPUApMPIpicQw+ncrz4wHBp5ZaDozteIHfy2YN7jgf
WZRDh2hnHK4jJUxjTwlaS1VyR8abcxktXb94y/QAljVyaVMVzt5vDKrZl2IO5Yx6
Wz8HsILl8Yv30LQOwlTRA1F8pyLMQ4csq/IepLpOVya/jzHaIWHpvg5UZtQMI4ij
u4PuVfTjY7RNAAATYtUWwPAQsY+lpMWN8ctmfKLL/Wzrf1nt2vutytYV6CY5e/Vv
Es+396Zh3ebeSzp/TO2ZSBkRnRY6QQlSPrUqfNFSLsa4aedFOMiYuvrv4SPXkz3I
oJWuTCZ5gc5Mu5pR/PrUR83nb3Y3mFtszX4FrD7czofCyojLWXm4TFJmqVrfEdlI
p2/kdSVF4i/710VKAk469U8IQsDuaxDIPsOJlvx6HYHNn7p4eZLbq4MACTRAP4z9
2yQiq52iQ358ZsPrW5ee+AKr1SbquM+FqPnblg7RK9R5Uz32N14qHdM/C+nf9/5e
d7xrjASWc3yB0N2lng5rmjMvpb+9UGH4uqLtW1lxUNVXcwNXqMa7MZop8OK1b7Pc
fPHLDXNLjmI2nfWSLm2CrlyS4rFd/1yW4/T5SI5+yqJiWLTEMYEnrgjIbY7kkldT
twoXpcGKloQqSEDIfsJ13YMbt5FkoMP41LU2aceWs1v5j+2Iao7vIjZunrKQsEH8
eZyoFZsEoGO1H8Sl4Pbla+48mx59mzuwydndXLMwKXGywtrXG/Ug638cy7WHrAQb
VhgWbT0m7+8Qfc/5GeKn2KdMjcJLlidvQqB6QaNq/liLxdJNKCv3cW7T9HNfyGuf
qy/GH+BG+DKK5YStoz0k95nh3RHxNTYm0TQXcyqqK7YpGzSUXLt2/OjWbMx5SVRt
Nfiw3z90+4xKCkTiCd47fzxEUTLx+glBQ1fvZydpYXZa0T9v4RJ8Aishwo3A6+0S
TA16D6oOE9yh6DlZVvtvMaAdT+hnNcrbTFSc9byKoD+/Z4JtnoN3/ZlG+OY8jlBu
llOBgabsxx/lHlj/4rYN7MufvSheG0XdlT1s8tDVzWLMtHfzku54mEg+vccGm2Vw
n3i0S1FCmjQVmy0gtQiKgKWdAUBeps2Akc3appGt/xKQjz9krMmry1yC1SK1nIJk
NVpVeeRHCyY6EDpmDVyldYsvO2ADE6sKWUj1RU2IQoN7b5W5mVEJQLA719nmVdeJ
0HDff2Ycfe6hXCE1wlcm0Qs3l3HEToLQqDy8l4nJKQiY6D8lc8bmWnEf9gdn+FCk
4/AskL3MYlz6xPoUkUjrbq2CqsX1xTjVoKJZwiDt5uBOmOeZeT9NM+tIkEHs1NAK
mhlCky/X7jQLJisv2QZQMtzVhAPPKtCh4qK2kmykGYZ+ZnXSqZvGTRf9NnvTa7Z/
Ye0kPhMvcpIvuRA9BPrl8kjnyh6NVDQCUZzliS7LN4vUfYj1ZTFxhLoaVxcBKisY
iRgWElBYNbxeCZjHV93yCqmHqazlKfJ1qLciZCFPolF9AmA44gfaopMj3IzxiPqH
R5QQ/XbLt7texspmFpWztID2AYNFoMv2XPeH0h43ypW8mgfEPUObd3D/D31Pm63l
tybMS5BfOYL4HJn2OiOL3TaSrp/7mLmPnb4h2Gd1V0xUf+welGwFXa80iOqhkTZl
dkD992hq5PTRm9DbkD816Jbv8AqtH+cU9UDh+uW1xE+d7IofsELAbPpO+uzXIqpI
4ybzPkRxx33LcQ+5odvg+jD/JB7XJnQY9pkBBeLhgvEstTXA3Jeco6G4HJnwhYUZ
Ir7ei7RdayYfo2gn1+ILRCKUk4pfrLdkYX5/ku4ZP6q5qGO0X1eaPp5qXiVcAC7m
DmyrgIwJIPxt+cm7aXHzw7BNvpecFJqgGtUSClG6OYlXVpUfoeWegy1SUq+PFGfi
X7nsqSTM5s6M4y16hVKMwG7PJRzznM9W/0nuAzyOrEbRMgOINCBksu10JAHhCqzr
4v70mc/nHss06uVlQXiXOWVsKJtAuNBKgrWGqP8zRTUECY6JMYskIZAebYQ7AMbn
kT1MhmI5hUcaSnMsam6FmdawexxX3uoXJI+hO/qDEmVDOHoExtcFYa9ARbu41xsi
YWlelstrVyaCYRYtFFCDV2sdF5fBMQuamJx+hGy3Jci0gKF+IcH8tzSSE4Tdzvbj
990kvyULwrdVOLPLZ/TiEnybamCe0r043AB0DSGmyMAS4WKC7432C66W1WLLIE/n
8GbtIfJwTkNcpDKhQXfiuZAVgoh66VNDFJNd13/hM8hZE+DIrWRZMvQXjGrUz/oa
Nx6Yg91vrdr4xTvvNxpxWbp6Mox2VcHvjwve7KY8FSGfpjw7RK/VgczFEeGbN4W+
2s6aPekvy2H+08jeygv1VV57gl88tNw1QHWm0AODnsmkMMPvjIs/C9brs9++DTpl
UpzjR5Gkqoxm+Q5RCFX7GgpbFu4nZ7CEV+6dP3mOqpjftZYVDgrfQgHAoQnsOnhp
T7B+/IHpjn9mQrpVhjVjiV7urLfMJhcccK2rBAdxtIXN4ad4dfz9CIFuOTAotvXE
VFMjvQjUd4OgOpLyRIChpdlpnCnVDd1resQEg9c342i0cTgdI7WuHl5cmPTbIhJ3
Lyv8rvEyOeiRK1npzORZ84c/cSD9fBYrHPcYt5cNOybbwti/hkqHIXgFw87Iz0YB
HdsnQh/akVbf85ZQsjv+jyDR1tfYABOKJutFU99HQPBDhKEQhZhfShH0twMokwda
LOdXatI8/sjlK19lzelewHGoQB2gXYDwof8dErFVpD3baaOVTBGvetk1I3FuPIeb
CAoCB9aQ6mQj7dTyeMikfP+0Y9A1AJUHtKGw7dhibMgL6OulBxoPNdvGJl+YTkHg
FG3hdfpa5vsp8BVbPzH9u9kC/+vIoAOwalKq2aBghescg3SpKgkf4uGKgy2dxsha
Pp7BNvbr4KuClUWgqysUmr5ZajQIVljJfnj2ATtEIeb8XFtBXk/CML/0EfR1Y4fE
Q0PL2OTe3jnAWsF+0jtrI9Nzh/u7bA53+kpNX2BOYi2kgVWT0gs1X4fedjLsoTff
dQNtK+gVleV39e4tEWhVBnvCfHoUa24XqxA9MJznhV/9pwW5xEejUUfG8cYbN1BR
yxPo1EQX1QNHyEJG49GopxfOlYs5K0S6skfcfskuSndjgiWR9ISYfc5IzYImQ7ff
Va1tq9Rgi5zb1thS+EHi9QVd9w93PtYNMwza9v+Un+6wy1pQCL3PAZT+uF0TjNUW
N7OajKnw4hiP/LtRs8SxfVrmPw4j0O6UN/lD65qd+BCC9fT0/InTSz3JBnho+2NX
nN15XFyaoDm2XAFGh3Jrsug+O7lemqo2qfaihlfq/zA8MGLyKNf/jRvI3RxArYA7
7l+RH3ljIcZh2Zi0XrgxTkRAmuF6P4JOfq2kuzxQt8noyLkPCis/boyN/hQNYYGU
npz1Llzhk3tRPm/FmjkAhTkr1mlqC/8fLO+W81o82CK+m2oENpz08WdwMJGZeCKW
6LnFqruDaKjZJ2Qjgt7MbQRNkD9Yip4JTjCjFS9OFKWmYaiM2dVrpSGCNq1QMzoG
T/Ja5Na3EqrSSuk0k9W2YCovTiQSiFL9xXy02R2I3RA5O7hLczNNOxLy3AOgfEuM
G5Vaven2ZsjgdN97tgW8gChc0N5rz/EwCVQkzDiDzvG+r+YdOvUWssOf8bNATVvK
iVTJrxQnlzL3RZao3EKABWuBfAQwHwiOPhypy6ZUwH96shSluVNpFIEolx12gkjB
9wl3vXgWIgEAw/ZovPHKLNSuuSi5pQTNkpv3bTwY8gB0uPNtUJS76Dg6SGZoVLJ0
eWFKMXmUDVyC7FY1eDezywFy3KJFamYK0dSPkPBv044Ce5fjUObGjaPQqt1A39j6
RCTKZOIlWRItgKj02JnLKSe9jN5yMdka+/Tn6wKgrGN6hZKkO+snwlkVwdPhuQB3
HbfbYSgT0oVVgWWUvjAQVhF8h8lGgzDHO/IXzZtRtvPnGjBnQT8e2gmP1xsXBluC
I7JQHiYzbQhG0RfuGUWWt4g4DaEzjafTIRlsXe/OeL4e/FWOcTxqG2uOcugwO3th
9gAu5xT8A6IIopkxbFtr8A9AcnyRw4MMPLrWSr1z6TpQHinmQptl4WbUgyGbAi0J
SULEP4i2XIvx4E50o33vHr76Rjb1SpVNR4tloct8GSNMX1y0LRmnpodyIY8m09yt
wcPsSPpYsIEDO5zQ89rGFXXuo/oJceQSITzQzvi1M+bwkn894Fn14R78GZI+45z9
LAiilWNd6WtRvjYCRudbsLlDZxeQw7fSev9769NFKYfHnFi36uWfxAdjA08CSEAW
QSSzbK/8D3aW31imZ2Ib66da7SW5XgtAQhmGTtd5Er/ci1KuJrj2mbgZdzka3v1s
LN6oNX89afpI9pi9+4Y7D2bEpR9ArgC70Yn2fT5qFKRasp9uifaXytvJ3aKiQKXS
kpQFzEB8iyW0NrRGCUM/PE8UQsDQg8m93v+tXar5rkMpAjbS1q0AT0Qe3XU8lCw5
JZjuPXAa1BDKYUCvdG04jb6ORiUhXPtcUUe5Q4JVh1amotKvUK63eYErB5rviSZV
7d+7007UqIngCIC6BrSWcE6ycK92KYvlHXc5hRK4mnuuDEghUBxfb21VuwIR9zly
ANtRcYIbPmZeQbfhvAv+sxWhS6R/WzMOd9q76QxuIQzU7Z40kWuaQjpBQAmLQ7ha
vCdMLppW8p0/8icYp5RhqnzxhAX6HiIphgYxwSkOIzblxGj0PD3+WoRMibWVAifF
7g7As4v6g7LRz9WhPjqr8ZqtFpXEpwK72Xciabpf8Vgek4VHEtm1NiYz/OJbw01y
LsCCAu8nFm377PJj/3/LDxX1GhhA1/O+W5SdskqNP2Y91oWt5IxRAr14o+P/Ug+b
fTIju9NbGijVAyYYZq/fBsOJ953k0hYRapkbdujAVc4kCoJ67b+H+fEAIbD/BtpX
cpdWNjSZbcpBRd2nID37001XK59nCGb1CCCFXW528vOcIJ9l5x0GqTnQ89TxG5eu
Mznz5wX36mQ43alEmCWiLvBml5LUE9FPBu33Nv1d1ql/03r9abKHjX3Y3J2oz/4f
awCepLOEJ2wRN73X9k69hEd82rrkIs3uHhw8zGxsWu/B5Rmm77zyfH44YtyT/Nap
hLr1C5M2DHaOKs1J48/yyI3Mn1EPiAOUnFH8QRG8IB05ZU82C2xI6oUVT0zVuwZW
FliysJ+WOPX0bTXWqR4FPJQ6x0nErmpSXBJcgyD+5SWEVcPx5pWFxMN7cNAzsKmR
978MVFXK/WLHZ6uXEbirbz5RWK6a26WoZp4TzaTq9GgzGInx0mMMHOsmC5Z28A1n
tGdiQtDkNpnKUOnuIVCAFUeQk+2LkBwsA4n1+0pClT0F321+3xPw5yvFMKP/+fG/
4C0Yb/WME0YsRda57+ovbTrB6qGsyZfs2/xStGOT9K/FNILAJ5fNXafCws7sQ83/
SlQecHzGHJTWj9axqtvnEpgCTJmqYnqxIj7n9ZdpMdoAvXyhWFosfuAcMnNe9b8x
EiNeDyYePFapuSmLT5uO15bIvty0ozxVI4pb/wPa50NBfvdByP7qJ3eovAEJWoNA
gOkvrKTtU0ONaggJgA4z4mUVPcyeu+/tQagC793kcCnqX1EZqToS++v1HvS5W4se
F+u0dBMq/7QlUfkU7YjVWh2LGl0ZkmTGMjOxAIFnteH0zxaQtpOPwnc/7NpcKly2
0lBAa8YXN6iM24Xk/a4yqlL+/Pp6SgoEPcOCZp415lijdhcvCtk21i0A7Locp32r
E1cRb1+wW4mbKXGusCwD2mcxyYO/Ls5oMDls7g+bRvgvftvbQNWhuhxP6NakNY6P
eqLNr3OuS/4diMayOacul++O9APY5xBw/lDoSPSGx7XdF7UfjWXrMMqV5ZvTpHR8
gzeSdhGcz2vduFEPP1Dl2VOJxRui6ufOi2jNbwfoqAqSDjwTxxMhe60reyBgrcNh
BcIfzCf/1dfjASb7j41eWSP8TC6b/8HwtOyow9BGFI8nJPfrJaOBDxnXjzCGHvk9
fyeAVxiQ4nTlMXwrlmqZmhf0B0N/zjiF1FYEX0h/qg5vpGRRlyLDDMaFoCErw8o/
qL/NVoqN7Dl/oIW4y2NO01NF4ztu4GNBFnLjecSsevkoS1aWnXUif06g1QPmzqIL
IntEH5pptMpD80mGZ3CQVpG/hLy+xXmYt6Tk5Q0BabK8/b6YLtLEqCE+G7UbXgE1
g8/o95SFu/W0AtLjW0qj1L786lk36rGkBrgZK4EssWVbFUUxro/asgbgpwVN5d80
OQmrx3NdBT/cQv0m426cz7AKIWSOMXbz+LB/8cMpSwH1j0rdsqJjXIPgbOGPtt7V
qcZTgkHIDGMHNcRrek1RRfTcUhCzVTowjt9fhMd0+I9pFKL/6LNI9zdnnKHkONvB
yEO1gnJGrrWIXOu+kpQH12AVvg0G+8K5Bd9PDWhUTNcdegp/lnUDDlSpr6kj04gZ
ujcue9DmuLpqmsmb9qkKu7HQlaLAYu+E79N2gfKyjbUf+JGuRet5n+Qk2kMfjCNZ
1xugvHb0VT4DEz0esxZpcknNJ3kAsfRVu+/vwxscjmIf+Qth1cJw9qTOrhfijO8n
r3mKeQTACnyL2qgfWA1beceXD/ONKgnTHA4XoK/fV1DfxBudEHmCrQAFVQTKUb49
Vymq2EIxh9TyINgqU1Mpe/C3JZllM+m9IzH/spZMaBqii2KxDmlugOTJoSHI7URl
8KgxjzZhWeXXc/b61k/LkUqywd2KoxJkYU95LndHk4n3R3Zqx1wDMNMbtrIwa0GU
DLBJq7Xj2kjz5plTrHw81WBkt+D79ts62cqsBbJBjfEJgEbJf+OzNo0g5sCePwuj
WZ/XNwLfBgZw2Q5Wg/AGE2+8mAHVINjO32B/6t4O7fnx4JPdxqfRu1ptcTo3Ljtv
gG6xWir9h5DQZDidJ8JOv0ycgx7tyWxjRFRQo6luiqYKhIc3loCp9j3/kBFLFbN+
Jg2dn7HunWU09ti3f0Imenksj7ZX4ZmyeaAhmsKeKOiU9h6J7yidd0ytiHu7Y7cx
ysdYxB9OvqyXXY9hEorGQNr+DtsiQAgSiEeJm5hWbc3aJrrv9hWjj3viRzS1bB6i
4NJgEaCpcsW/t90cabD8w6TDyQnameq4AdXO29+StCoAesglxLWgSk5PPDhHo8IH
vEwL3d/pdwxjNVPqqt3py90uqQTiEHShU8zB0SV7e8ZzWrExx05L/XAfN9HQo/uJ
ysTyV+0n7r8ZPNVF7laVdQGSkU2xeptHQP6YloSVBIZ4JMqCEIAgCaAgUpUx+Piq
r0y2fsVL2E48FLOGa/f0i6brF6S6zyic/1N/jS1Mv/rsEt67l5JlBJfKYbOgO1fM
3tfSNfnahuDkUuE3ooZqqR4b4m9Yl2UhQUQWNYfesHLkWTYbHIOONr+ivcEzZwQ2
USZtzYswtsYMWxoF1OJQFRbGULjDwIUMGib8iOT/Sn4nfo4bXE8LvqBwkcD7Wbq9
6Rk6XFzyKRCY35jeUpoJWuuSiqsJklJE1aMLu6fbraTKDsHblVSJp8lJnOZ5D7CG
GNKAVnaD2qxuxZOO8Rf9tHEUX6Z52wUNSwFyTSyAPRRdEsOIFI7WUlvX926rSuSi
CeImOQ3rA4LBjSrYZe19XROIWN/uF4f4gpks6pj67wp0wzQu0up08MS3IXwDYb/d
u0uupKMAWEJbqth1GH92ztunsNhDd57EZZSs0K0am74vRGfLhYSQHpLmhk0xEZK3
fVrgD8pQjOanjWz0NjFTWWh4pUT+6aQLWd94pT4Q4EEG8thOTiri9JqNQNNtiO0d
9YChOY2XGRrO3S2+r+aK2ctejSOcMqj3cSIo7yXsxSMq/MnOuajPidiTS3dLGhH2
/Dr2NeVwSCH0JfrZEt7wE+9Iwhlsb6MS2mMmBRXL2s4Ur2Z9aIkYtMxGXveexskX
CM0gubbOgj19cRgkLfW4RHaSZaKFOt4M/CVARDYlVK9TBvNFxKuiebs6i9MWSPRQ
dqf39Z9fRONuPXplnQyjCxUeSZKm8nHf6RU5rQ6En6LgMk/tIHACYvLNQWkTKHMr
8IQ/69Kkc9MAjGh2dkOh7J2DcZ+EGrbqUUIbeRX6M1FgZbyye1sOfOGA+MbygRHR
EEZOcmKfH9NU7VPsx8o2MOyhTFL4ZoDc+VbuNgd8/d8RdS2/uAc4gCSCLshidwLx
XVmAxQwiRG7qtn8NNs36gs0pKcsfTfopxeQYTj3b4Lkr4TrBauIAxr1Vb81b1B/R
ev6u2RRsmCcaPNw70b2kLkv4M5Dd43CyIBgRQMTHT26lLqIDsJP4ohfq8wGqeB7L
ddvr8AMGAyavvJo6uBS0Br2xGjrydi7nXfdQ/Tp7plX0W+b3XdKdFi3lB1NLHzmC
uf9xC/QoW3OnlRFVd9qpiuVJrbcW9amYpXqW0KkBTTNvaq3iohyYnd8VyEPpoTaI
6quK4T/g3Xi1TPOy0arfUnX2Y1bXe1LVm3xAlIMtuu1bPMBRYsdkhB3aRPLi9b4U
AFyNjfcF03bGcEa6nTaXpeXItHA282SJZ6Rwf+YjF14BhULw7X98Atr88N2NWnN5
Aancjfh6DlCEhsJckX28rREmpY68K7ir0q/Yu/Ei/VQrgXisrUUZdf4Iy08VK4Rr
mkjp5mNzSN01nX5yJNQFj5k/9BRIOEd3CQKV6vUIAujYTddKVAZGOlxfYjLn3rbn
Q8HYBHwi3PdMeLUAfSvdSgw26+pgrBWcIDtc+PfnmWDJ707+rTxr+P4zCDpeqtaB
VrIy8ut8k43xxhx7PchOEXrloJ9KrpgHaNk6kk7MeSVqRXpxYTwvLyOBtVRgEfSB
UkfyDSQs5+Lw+F6shKpnJeKg2nvK4cR7i5wFBAwxU6dImarTSl1K8hEP1x7WP+U3
nYQuigrJmB+whTsRH24QUCCXvJ+nTPeKAHbG09xfqlakAqePEnlbZs3sorWOJViP
MwMihS+FGN+PupSH7gwn1F4DXwDfjxRl4KVAfVKRf2RwJr8DZKm8FoXE0nsks33E
G4qMEmU+PfP/icihordWp+exhqCZPs/9fwuUrlI/10Z3BoQkrCBgLNab/4bHlkqp
0SQLOhrm66Cn8FtuTlHqgyDCI7n2WF5qvVjAVAtD1xQ7/tgWaY8H+HxtH8YXmKuW
vUmY6TCLz45hnmpsgDbx+UcwkzX8HfnTYPRVenUltX3MzDNajAEhaCVfEEL1X9nx
WecbDrWfIIM7TifpOlMFqklXATSYVTa4m4fqeGJ1iS1GqUa77aGhbsAJuZFu3zHG
iWWWNoR5wGJe+Nzkgb+ifg34NNLllML64L4GpvghZ0X+g3FWtjqyBYx9uPpv8+yJ
3u7m4qySipkR2g0U/03sVdlrJCjFhvatNDVdGdiGwyEeKqDysaidTk2On6PZ/aBx
EuG+R4NeGor8kYiKCWmE9+W8oiPxTtnoWx/Ky0UjRzQsiZHUeOD+6i+Mfj4+llbL
lfKs3H2Lu2P4e8qx/k2rsuVWrOWFgAPiFozRLrX+aMid9sjFDg1ulSWv1UdKDS1e
QrOYD12xwcdHGZd8NwnlJFb2ut876WEso8hpGfYNTLijrSZ/rIxxuC37Jrofwkkz
vUQ514ei7RuyeqI7anr5u4uM0iM47C/+yMTveTN0484hwYmSzV8CwKUIfUCDWIO/
I6RHgcOk/+Yv4/JmHGOiAGcisZRtGFc9f8exi5RdKn1GM+dnwA3o98lrCj013MiX
tMZm56AhLMYlzdBxWoj8JUMUUMp2pV6eT05CnRwTLQO7oEeLGOltIkPLC9hE23wu
iLQKmr5X4qTlcbxSSEfm8EU760+494118Owc6uzgleD8NXlY+990W2tl0Ve93Qsz
U1cyUXursIrNQpJdS/biOBW9VcvEaswb1maRYNQqIgfcJXxY14kbYMglK9IFqqZ9
lzNvsNYaD2MbgyFODxpgDA+zLfiqxPVJNC1M4wU07f+btrLmXuPSRgMVQ+gIJHNe
VJ4TH9iIaf5mVdkgNKdZwvnHIUTOoVl0EY4RFi3nLJ0Lfk7v4df7KDaq7frLQ0jq
QXZXIhY4dQ4HfYJdLSNb7CZeD4/MQ4+d1nOkJrLs/n8cFrlc7z55aVjpYxy4HQ0K
Kn/VKlnyafiUQVBXf6lOfoEJH/1yKcbNnSWmvxi0Ggj1RCVcL4d3gyNLdJaIPpJc
cmxq3OzFiFwNdLGQEFlOnqADTtXRhPG6B3I03AZfmqvHfVOyrEgifdyLUxBVTZ0y
rRz+sCYoKMmc3vWCrc34/E2mfnevzQu209Jl1E7xzBTC/+PcpNmLe0g26Fp9kP4A
SRgYt/FjXo56J9fNEty+5aI7TmzdxVD1x9zgRacewuhcwI0JerQbV/eiO5U7J7Ty
/GegB2mfWXQ33SCjC73HoIzWu6dobvWNUrI2b8aTBXeD1N48Iq1xv7KwE9mQbNpJ
foKpTpMdBtKWEXkRroQXIAA5/zcIcSKll0o6vAYAYEg15WbloJAn8X4Luk8zJpmc
IqYb6sXIiFaugJJV1i7mgJ8LQGhSuVjS6ZGeUCrfdJgHrqgFHqaKnKiK7uEOnOP5
zVoK1MOzR+b7ZkTvqhHqVpLSv31uNZTNlrWzJQLK1CXCwvonGPvaa6wW99M0RltD
OABdmIe3szl8vsGMDk85rsb0Vydt+t5ExvjToZpE/ATZwF9NOvrhPiTyvT2EWmwK
3jpbh6IZi36zC7g/KJ3uGILVZ4ri4pisE/VVhNQ/Gd/K/rCL40H5rYx1Q7Zc8oVK
wk6N2aizpdkfa7rbYoQ7bpdPXP/WKnKi/HOLYTlBJJfilVHoga2ud/ifltzdbiph
sZB4OT/fZwG3vv206aZMZlIZZHqsxPAe72cw3qTG6qRSJXufzdK4KB9+R1+4pNDf
yBrr8rVfJaCgD81QuZIMkdR674u6miFbui01tONW2JRP7hc/A6H7MnNZOl5aJF5v
p3iStcWcGxcQbXl3XWN/j7Qq/89QoXMZ8c08zcR2w15ZHYv2vsNGNCDGaGILSkr3
dXAfWZrDppl/J0bzhIwrFNah6U+t76nHy93sdyonI96YWh5BkbPFcBqz38g0bI+r
BwOSKEh7W5tewDH7C4oDoHzCrBaBNf6KaSSVUgMRaQD4TGse9+HBc22yCjHXkaXi
YmXC+D62Ewe8+E3bNwaNKj7u9fJJDdQBnBNLJQROJ5UFyMDXachOCKwJmdkHPMUk
fXuVA2LeOSRKRa3n+GjLqdJlDHf9V8XtbD5yBd8mh4mZJ9oiSm3yn2ycDMBfgOEp
rpog7AbZdmrzWoGooEbTvkPKpjQzApCv3CaVwW74npJPdqr6shvb/fsEPuZ3ZJpK
uxAmPbhwkvUsq7vDqkoc1sIQphexQxeA4a1HQsRXrtHQEBAPPnMU57BhvCVgGCqj
b14xrB8+Px3T1K+NOypsBGEM45sbepI+irJjyiy4hZJ8dNESYMBhO+LlcQNt2+jW
PLKh8otswCMMcwrb5NTRHAZXwJrwxx+LUNIrRZ9yaa95poYLfqD89/NF3PFZDayx
9VikZZ/BLk4o0NEvx8auN/3lTLdU+yy0zYRjikyiFmVdf9G/3/WJMCBLgRh+GlBD
VANshv2OUNsQezFdsHCY+UiU9G4fnaxCuGP8Xn4nRBQtLPmmGvPqfoxtlg69RJJ9
jXIzTvfYweb4p4mXXjwr4shHTUN8R/pA+n5EeWRnC7lXljcmX6Zqtfossz8JfZOo
/2fxay6zHZ1xJZ4OljnEKw3jiCSbY2vmwcFpYvg1YwmJXEu2q6HEo5cT0k9yTSt5
R1DIT58ZzI4O+jpXqzrWvEE4qMF+a1WYOSxYfvrsuiS/6WD52LjBGZZH0fOmhBLt
WPXL2YVTFCrUYGmG+NDN0ShifHro4VRBUHgvKqkXIUwTCGI/VTDiSBTKYm90ytEz
JnTxuoB+WyLt+ibBtaDaflNapKZYg70woT/m+scfgIk7Uyr73rpY18u7s09hmO9L
g/noCAV7adB95SlQ6fUB0T0tuFRHWHtXtNEW9Xe0LBkmLcwY0Cch8zS4ndcrc20E
GUGpKLGw18/2zNxg6Qnnw0hU0KjxK6qpt8vO4vO1nqklpWbwHO7D02BLyPf8vVZX
svx0K5kqSXPgWpHvhAc36At1jKnMEsNzxoPuyAs66Flaw4kEe5tfeFAhrziCQwwS
cZfdoRDadG1JNu0l6RfdOG78zLPO83vpZLP1QRmLtffC3suMO1eWYlocQMWr8o26
3psMMXeC1IL+QCbqcfVVEQTQor7oc3jo7KVcOVnr5FtNHfabToLYGd1M3ErJq7pB
ieU3JGdSLiDnscC11iIW0/cbV4/wEkc3s1YyFAnX1L5tKNNnL7wkX7rnnj3eHKRc
hArstvC+5MNVtIZ5Bj/XLPP9QhH8XQ2zSW+MXajjzgVm09cCrs0rCrkPXYmbnWuz
y3KDrJgjEV72lqrGqLBgRZPtcVWRACXklkg5WR/eRcy0vdFDB+iJmsp4uwj4mPZ7
wtVCHWQc62ETa0pVhqfoZs0wCaUsAN6B7vzW48WrDDpcIFwwYHD8dw6DIyQb4BOv
7lPKMlTIvu6mMNjf9gB2ErwUobQfu2ZnCJfHqMMfC8slCkFhisuvXzMW21HvLLFh
nmrTTjNbKwCX835R21tnnpPuJm+RO38bUdNgjjLzTy/ivk5DEC4XVkpjd5VUjB21
YGXoy1s2oJqYONAf1Uvbwd8ppevkjoOT4ss8aZkatfhB3VrzPqlFbbJzX/d13ZQ3
IXUljt7UJiQLmIykZEnMas6fExGaa6AOpPZ5RO7bovL5nsYhNA8K+gIj7VmCyr/0
w07g21DL+43vTXST+O7yJL9nYgi8P2CTwzz7wd2xBOuXxroXssp/uA44u3ME87ng
q2Z3iI6gd6Jc/ErjVVnYATEii7cG4qavYs9qKtFCr49+aAU/bGy4apfwLnR4Guno
AFNshOyKzr2mpNi60XZONIarzKkRk8htG/JrhrY9oF43/Ixz41p9LU7V8laMfQ7D
DzeDyh3C2YCXDQ0zXIs1fDmY0NhSrmrPAbcjrlRvQDb3DT3E30giGUHT3iuouAJX
372X2jgkUeJSLoN5Z4K4M4H+RtuLLXhtvIPTML/9o+SBaOOinQPyR45+04CAcdWp
G3yfcW0BGHNl8la2ATGiNGpCxCWD/kjMhtWllxMGZ9nxGfCn1UDDH/PW0XOk94PQ
BRFyD+OIBv3IysuFK0fa4YqEvbAPYlR+SlVQpy6xQEuquoUX3RmIpShlOoDvHlGX
pkRRtBHpavP4XvKBm+5nrS8dJC9Abs7dvIxidxEMkJIUqiozek/bqmE2b8VGZ8s6
FGDws1XAfON2NAP4POCKvEVAeXBPozjvwnd4FRAKjhcXIhuAOrW2WdDjRIwj/VPT
8qjyacdqNP1iZGQN98gph9PbeG9O7AqTK/769UBkEP2hJY3OvTenc2wLmwzmPjOM
FXCkRtHb4kWLbEAztbS/9/xJtCZBdcqtWmUtpgLbfC2Q8fNUzM23e6SUa0wdgkRZ
z3OUDdMR8qNW7JmjPJge+MxtqDZWrt/RJ7Re+Kl/FzRJ27DrQweTLoZuNagjs5Tm
JnQNIFpcUNLImhdj+2XuJ07+C/MT0KSXBDvyUDrOgHv/AwFi2bbOcs4uzAhyz5I8
Wvcjb6iSE4HqxoSJVwhVVv9zEFNGmz1LugheoMfQ0y80b6/qTQqKu+tWEizTlSwW
WCEStOGUYj9aOyg8XQWSz4IRVIMbBS5TOJwtIZHLna1tIVP7G4aXE27HphZt6utx
Jcfc7arFIinWS6+dhpr4nj10xh3oz4jsw1+J7m6SASxyolMq+4vkRJ6xBXiESgRK
zkhCjAjn8MthGERTYfAtuxsOTfqG1KnffIcYuNJhRB4RHGUtXFkusJVnF5NjEqsT
DT7wFCBIpKRH4Yn9fMxnPIq/nN7sta5d6owA7yrVtR4ENxMMBWClMOjBhk0xEkhZ
IS7dwxf5p55f1jZgwZfRAzZVfcIHC/e6tqp24egYCmMXuuajkUMp5I9QTZlitzkk
IhuNdh2vX6IZvU66cqUcq4a15LUcYQIdlbVUgyi+DxGf+nYaw+aECxjB1VqvswpI
avnlotAbzJ/oTFlXR2sgGaugdqund0DLutm9whqGrwbYQi1RcXEl8mXhC+XXAY/E
kUFvQQd+plaSBsf9N5g7Mjxb30BPSYeq+nL4mUb5HE2M1TWF/8ELHsmE+TfWGs25
eGV9ZVtRFraIT7WpCn8rGuc/A8p35TYmpfslfJaIxgYPfvzMrYPdsNSd79f4A77S
tAohi+HWT2GL/zebJuvKRHYAeZyZZsqUK8uOC03mCDIfj/+KTFaAMy07YVVifLqi
TCAJTDLCsGKSNNFpAM82Vm14YkCe51kXWmcAt4tz3kmi/v0lU+kRrcPOf/rJEsUL
hTFvapkMsPCmqpC2+yCDrE2Z4UAVEDs4tUnIXOdr4q0M5NINtR9bWw2xQ3WuM+xp
/w9lgtjYIdcyph1IQkvuExb+WPDx4QaDeAb+H22CFh2F4sqJRsfzSiVAcmVbDxpN
mW/Aiahish8Fmqz+gTE9cdVAymOaSBNayuoflAIGNQ3svvnzJLOloCq5lMwKSpMt
woT+PsYjj53q/+KJxHhZSeO9fYIm54Pxha7nCxS3Dpa8HyAYCza9FGOo4f8hYtZ8
a0amVX0N5vO1bVy1+6ErqV9no0gbYKYwAIRbyOezeqVU6cptuM+WU8uTe6+PYCzk
QkWur+ITzwFmeaSftaJzIuOwTVdlevAl5h6rB6r9niUUezoll0tm29EX9ubxz0o4
fctUn+5RbSPKShOEqOeXUJadfGk3Y5bGHm21P0aYG/5kZmES4nyg3sjtvOxtFo5i
hol5Y6kJ6Rt3SUN+K9aYbQaYJakM4tk5e8bur1Lr1zHkFw+cb/RTZsRMCLXy/iH/
X2aKMwSXm2axQ1klSq/1CnwgpUVhj8ZVW4nOc0xkoXCmdXCbs+vKvJVaScU+4v6L
n+GkGXYngjyneOTc8+S/ymH0n85Oq1qYbGeanLmmSsj0+a1kLXm8v4BTt5iOWB7v
92uECbbra66KsIL/ALc4cuxe+I85ALv+ZCS2xaRikGBX72JC80+vmIZjVFASgxaJ
K5N+VftTiWHKdCYYy4+wakZTKO0W0kX62rP3pcUzNFu7dnzQ4gwLamNpndEJbJtm
xTbmJvjycQQZznOUxG75BoQZiNsJkhuAuTdJ7Czh+zckZKcxxZCC7hSCm5a1aQev
MsiKoQ987dL4jaIx6Ag5I5lZ4OiWma6FfBvx0M2yaaILfjwlC0GTNvNUs5XogbcW
CSZrGZlLFRexolThxVKYn/yNGyQX6+HWozciK0F5N5OBaLJSUXduvWguvGfM/EcQ
dNyfPJlENmxVlJuD5jbCUgPoi9Z2UvrZFCZawfH+YnE7ngfkXHoNIBqewUm7pOMx
T7PKTEt+pg7VFdbG1heik0YU3RbO+EYgV+in4zKQPHWbiW4+JIi5rfGmZplUncZ9
XI1XsJSSs/gaJW5EBeTXcafkaK/OMXB0gfu/BmoO+5kO4QBbAWB/0uZHXd2cGpK1
08YOAx2oqjXdqgghqvPYykLyxvjUVoxwArOQDxSoUtDFDp5c9MWRmjHoMs6yiW4a
Z9JWPKvGhepQoaEb0yoFx6/HwZkvsvVejEh/TIObe0ssBkWG7lz4nfthgrFxlk5k
M9WTJ8j5NmLPwul8WRgED94x05Dp8DiNgFoyaEdQnjV+cL4/m7W60FQ95JkxODS9
9cmG8+O5gOqMGnORViobfUKjDXvYzWPxvUH8uVMu3MQy++emymBMbPQwolWbGuUt
1Sn9mDIgDEO6nfP4rklETPco5E2K84Y+DlJbljkEZ/m2NtuCOFJHVjo26qzFMdQD
pm/GF2QATHIl1xSnZPTX5NCuzEtLaLqYiQAKyggggVbf25dslaVoay5X8CoR2Vnx
MCJV//PzBDhiv+inwvjsdTqm74xxQ96vf9D47yhAPelNM/T1JVAbAdy5mp9KI56v
B9ayijHU2fJYB7ZWDczCNYzglFEah2sMDusspu1bPaS+Cfwe7jy5dsMJNpoDhYKj
I3t/5fmUZB9Of4JXqLwqS21rhHb9ZT6brcg6octrdWBqIFNzoXEqfDcio7IYYffg
a5PCHd2Dm+Yoxk5laXjKHyPtJU2XGTBb0CDVOlkvLjglgua6VRlW6bSESHNoZSoF
w5flBjfFRMeXlRFTr5iKCP94RbYUroEywRfhSSt96dS2h0J1JdyPIzIxsZyjfUo1
0gw6qkOIQEhO3W9bUS+lJGqLdnsxR+kO8Zrg+Qa5Uf4tkfH4Qa7b3R9HPEgEtdv0
0bmZDGIxjNBnZDacfKsf91RBdQvLR6YDZOPnT8xonvgMvbNeSvXCPh5UQGTxgc2o
fEKEMzlKRTUxaatg0P6kQdfK5r3hoBbzKVDgNWkOkQOnN7yi9/8GJydW/2UmRno2
Dd3cN3IaSopYLRAS1iIZSM1i47MFWMvc2NaqYdRwnldQwRggiYO9eAxQFR0t+w1Q
Fl55qmH0Z28zlAkzgvCeLpPt5mH023vF2xSCtMVpQ6CDUzx1xQ6+xazm2huiKD21
34AJ1HLcJlhZrD6hylFgeJA0Fs0Q3j7uMQFkNn4uK46vzyVdw+Zj9RKthjwNlNXw
DSIjWIanuGvR+yE4qWjSIcNk1P4kXDfaqgD1qOr5UTcsqJdafsBBo1UbTt4ap2r2
U7/PMKfCSL7hTtfynmOini361OzhjrzRGCZakoq6/xHJsq0bak2mn46s99ZC3pyu
R95Lin85Wfp6jqWCPQAqyfnp5EUYeHwovCDxGkWXp9sUFSOhViyx3GyulchaGG/V
R9M4mxVjlUN646Tk/Nh14imB0nYBDOYGsLrUTBBE8HiEuUU29u512hC9jOMIO+F/
jD3EO2pILuko6rJxEWTEjrGVh0gcitqFPmYyOjFx6xYWQMxiCX+mezjTA5mY1kmU
x50bKCzYoXWTPA9xKHHreuvtJD75BjJuDvrIKrjYdNHU2lQ8/LujguvIDiR7g5o4
5nLz6DEdIaSVwP/qesVb8veKw2hVmzOw7mU2xJyqKcdXOKcdVG15qK+kQNRm1cEo
1umVZcqCX+nAMhFTrhNYl+VdE62YHS+MTP9u3YTu1YxdFcusA6Sgwz748o+0+Y8h
C9h8utenYb6T9a2B02T49YJ9EAP4kNLPBdXn2Pxh5xKgyjQ1X9KybPeij9Femjm1
hRJo58znkImkzGetCwrhY1UdYwyjqm3wUJkW+NW03CIzTtVbiknV/M6QabrwmArh
mR+e/7gOQ646qmXVJYBl9tk/J+sXFPngV+MKpJj3VNWUxDJHoEY0jouYqIMy+H9R
U73Fp8bN0hAn75goYZ1wdk229/tzbpS6i1Qq9JtjXKsoKgaxMLbsiblfSj/NpUU2
Nsly0k2m1OQIde25EE+3e6tIYQhk45WSeOmxVRfpKoE8hzXXXlEyDtR/YOUE1RD9
mA4M9ZppaI2VQ5KxBBR0bF1y2E/cImZOhBdDq7DStqwHCEVW3HaBgRdsV9DsIMb/
ZVMG76+edLy7PDboPkG92R25mTyYKnRwXNVEIWBBh5SwkosqyR/Gs1tlbgMyOO9W
+1vVD+jV+oa+qrVC22bESC28JLgNiq2/OuctIOoB5FK8G/7UUYDu2rjIT9cRzhuT
gnZIOk6gvVUsc8E7R5b8XAyOBZXtW+eV+FI5E3cANysrlz4AlRtvGhfabXdJIEgn
2lVUvBZAu2mys/DyuKkSmwlKZqeBpmPonPnxLw5R8LI3I1GErsmQ8j9G1slDc4sQ
uBI5rfxrjbWYe0//wQHA3X+S0A1F7e/5TOhKtvAswdFzcdSgRTAHLNManGeBFMHW
E2RBTD4I8beyzten65DWIbFEQiGymVkAkSB+D6fCiLO+XTw6sxJXFmpfOAoYe8wv
ffVkUyypr413RkWumfqMJeCuhD3WJWoQJeIyqwqteZX2iOixyUJvu0A8Gn/DsaoU
KE/eFdy9BXfAU+QRKp3PYNCI8XrVmd1gMaQZaG3JOpjKJkvW5ipd2ajPq58rqDGJ
b0EGNKpXUBU4cdGZ6ct3vfuJ9fz1ZausZR4TUedVNtlx59muoAowHkDNYN/LaDRi
Z+skXWICYsiQPCWkl/4oImE5qbLY356foPBYZlbTT0Iz6s+mrLQAGSytd3VbSH3j
VFwirqfVhN9OoPu1z31P3Uem5V/PErIwfzoCrOj4asg0qH3cMcyDUD6gKdVX3og9
zd4ku4C7yJWaAK1k7lhXpcUYRvoLUZQg0p730i8z1Y8kGFkhM+tDdAVRUVU3vq47
YQDk6Zf+Ktd2XhaZtx4LyO4OjN/C14pZP6CSzHa/l5xLGFqRG+GcTI4mhwQCK6UX
ofWB7YQ7SQgZjuq/AsmjoAbdwzT1VqTnRJZhv4jCCX3lCqPV+QZTpChEs8hElNoA
yYCdAnJeTUZFAggyLzft++pKeOGlByYxmCNSIFmt8nDtTeTpoO+Xc9kTsYhi5CYF
U+f3AmdIcO48o1lJcTWfjmSMfCA0BDo2jCLeiutpKnZUrUq04Yyd4Kc+0u7JNxPX
sdWYvhRkVQi/Vymb7tIHJgKtLZymD45KnwYpLFrqk07Mq2vgxyB/8xZFKeJeXwXV
G+xaUJU5XhjpEfkg47HPOaOVbbDboIELzDm+fiIKMIjzHg1Lrd2LrLHlhv++FAvw
20wWiNDoZyptOlYJx6DAOfEjNCUmwJI/2fmg8MZnj3xE8aUqVB2rpcn+qj0xU3A+
auzuVWcQirOxDVpTim/pkXdBYdCTrxPR5fophcW90dcIpd+mUqAD1Kej1iyB1xmj
xGKo+nwm8Alvi5+uYiwtfV0g2+P4DetrS+MjEnujB5VQTifb62NuLL/tNqDX7xFU
aoLiqES6sGPXkRWxvPWbvewS2ynvX/xK+dpvp92AHmU+cuUEf6qAzLYlWodXLuZR
NDEDd7qy5YNm9IRBK8d+PgiGj4xDI/A94eXPdlGvtqiQ3Cl0vVF0Ps/mIgndpdYb
QyZpDXsWzWlOqfA7f3GvDQz02iVUCiOYMu+/BvYWTLB4mTiAXdT8BemPHasWuUMq
6bkNrQHUKRFADi30gpHqFAfSIdF02z4qbAonRvpCCdfw4YtCRzMreZHJkViPAlvj
U//0B0JZhX94PiOwxbnF2iyKzkpzYNOiIiX2QPTvTnz7ytN1iMpCXnE7wL/K6fpm
4M4HYdp7F7mONyHz0uwC8dN2+hEjijkfF7VO8lH1r+c6kGOfwM/fDHNSW+L0E0u3
CkbCCf2FOFomX0uaTi2Sl0K06DhoE7MBTZW4QSo7Y5ZciNiFj18cyG9lwc2VIHIu
DkCQA3kJP5326v+ItIBBM+GuW0KCX0IwHGexKhzKItKsOao6pNgl/AFy3+aPrTZQ
eILwFaARyCUE+0dZqnNDv3TAB2YRDPgB3SnUU69q/dpBTaLxflLF74wlDhLqYrqB
0YmNrIvPhtWsoZ23vIoIwa5BNzNPAqSVYnWZ1nngZikkpWagdcTYiMweEI39d1pM
VXXZ4FHLpQ81necHJArIEcoSl63IvH2kMprbMTTJqie+TCt+RrL+VwZvL5bVqOZj
6voj/yhgt0vEDlbTrty8dw5Xa8QzwyjY63rv7sF8Il1RB+Ru7BByUFoNV+YoN6BC
6C/bu1MewedbaUlw2prh5iHTnW2Ao7l2Fc1taXLMSgDA8d9NUohdDxQcj9GgE0lS
Qr+VS7sVyk7fmxCF8qXnCobXN/a6LKwvGTqRdNB6Kb3XNW+hDCrjQCFo5Nbv76W4
Xet9aIFU/1zbF7xLQ8GKr2tEvV9D+XnJ/ZKLjMDqVAYGh63kMZEPyv2oM3hMUOOy
ee7SK/GNaNFnBjt583dQIRnkbIHpwz9r1c9/ye+WkgzctikMWT/3+ftD3qiFNMcT
rac8hYQslaenazmY6X03b8UPlztrwNV1Y1LpdU/RuOCn2ScjE5Y/etyaq1ZUt9Vv
lI0Fhkc6n1P0GVhZDO4whtvUKkWfxrRhzT/KAG6VqvG+QRrmAY74VPC+e9fMV8rH
B/0B2tt9/86wqNyk4fbmShJcEhFIB53rtiPM6uaEJS4k6xrYn5K4T9yVjESvFnAJ
EEq+Fw04y8JjOYocD6YAcfg7kzVWHjnnezlrysFSgcICXpff00ijNpkGU2tZ0IO0
3MAc9eFRuMgPWZYmX7W0fw0RmPQDJsrhqXWGjkSOA8OXXzsFa7to7sxnqtn8tmhN
sFMYlICYQ6Yt6thWYkqSCM/8kX0WemG6XQGmTdtlc7mGt35ItbYGkGNuyVwtC59K
Ff8LU3t2rLHAI+6GRNVOw82g24e660oIFpCMZrlZHkpW+9wNH2kzoMGEnfAnsg26
xN0a/KWoc9mqqUCSsIJ/PhJJcrohm2HFIzAwT2RsSGpaf1nmp+RntgW5oYeyv3if
Nr5/NCFJaUq13uK+oVdIIy5zFKZHy8BnvkhpSGP+sbVwO1MlhroltdCmpfrjasiy
zUTxcPMwi2gFd7Cg2nG1mJ1S9GAigIykoX4VFEEAAAiA+oeiQXNMyGTM3b5n/Co2
Tajm5UG8oQK7wBzf3sQnNd++MvIAoi6mQabOVqeBU3e8jvmJsHgODBV1gZ3xUoti
SBxXS981njN89d4m4ZE79n/wNyNBtZAp4c2uGuz52sn1wFc9QT4REJpQZODXtuMi
XxenqbTjBvGtzHb5r7308YNBlLFiFwGyXmjVUt5qgM+AIg354xN+iI4Ex7S8KMWw
0kpsnSj8mf42Bi7KAV+b+UBBb626JX0pbIK1xKn9liMeGaIG19W70qJ8DYk9vV7i
AjRTJfQ6NLagWOsJDn13tIOAgTFRFNHoQ+5qZfJVUwVpb2Xoy+E6Ya40x5uiQZnF
TY/BKQySAwe78dwlGve8Cg7PoD79Ju6NAb4hWggWqnStJ01EoDZmac0RaMKUIvHL
2w+jpa/8ztYOdTMoVNmNNFW5ls0zfTVFWwN6U+/FHXIwA090ynedZQSyHOBsQtBv
0pHEKBUH4NAbkE0MlTjb6rB8qF07yIhALztAjCFqwb8wCFKgPSX252QORa1m3Ygs
Frle6Ak8FNsDgK5RtG/nUgoa2oPZVllv3bfWHvHc3IGTVI6B+Mi35WsKlCV2crxL
3dPQaAe5M5yx2RS/f3TKI27ia18BpE2luf4lBaE27xf3W9nB/aWsAXzPrKOS/6Gr
Ri4uhcCb0jN0j8wnOufviD1Q4ExWIvOZpV+BzhGeppYxW+ope3MaRIZ+QIhAtmp5
WO7NkLWFLk0Q1wI2LWJjrBrQP9mnc+AYcF5tsabV5Kw91nKf5isGevPpOkSfxqGV
mfVPKwuNkn5CGBOLUfi3kEfZ8xCOFJtV4dCeKJU+/QQZrsRHa0v03YTWchi2pUbM
EqUc+hIbiyuctjeEpQC6lvUW2RUUrnGAuudM0/axAO2+94Q8Ay5te7yQvHWU8PJj
DfIbSMF7Ynql1RMaxvTs5S0Bxm6ki5MwgHVXxgw0qJWOicAeMs2cW17OHgscMgM3
t7dgx36nNAhjOdtHCGr6pQ81nKG6XatHOwmLnQo74Evp2050CwVKfNxXVXjsAWrJ
okcqZRbCFFlrGR//1qFWHi6/gljOSVDF4hUfy7NnJxz0JoUVpwNcMdKFlNCSBFS+
RdgMNQm48Y8INLpDm+W9ftczSHzocALCiCshFoFMVRqQXMZRRe5tFGfbD7IznnBJ
qbvPffnhyTMRJNWOggCiEzXA345/tYxzd9eDhVrAz1CEDRr1ViArzUKWsCO69wem
LxrAYtSmAYWwGn3+teWoBlvLAJjszP0jO1Lf/CxrCzG75xKPQLX/cog1YlR5T2T3
ls7SvRhwUPhcuzSIlmCXDN4YGVXgHlIat1qCgTRjM6ypyKRpoViAmNiSuGJftAL3
E5lg38pToKCDjDR9rwCcLqRVQSQ5qeOTjcrdzIV/KCq7nQfQgbz7O41iGFIQrtUN
5Kua4mivjpoIyOmr+TxFPukc0nAJwv7UYuJ3zTALIEi32Cyh9iUf4UWMcirKcfac
1CsIN5bxS4ouuSTk8K+BOKGpN392AnxJMVDIE+0Bu7BkFS7xXSgugOucv2H5Xj0d
6JmP+XhkYhfyyiyphDVLsSiobpiLcxATB8Wth1ym/sTr0H9XIqfwTAvJ4RX67f+b
jteuJXjnl9ffIAwzz4DJB2AMb6VoLgvNwJXcGtKPpr0nKB28fUgKYWGpFomIPAAL
gUJrR2aaDtPS6hBehgYMqyNgSGs3kuLYKxCfiVL5g6uizs7NdGwt/pviOQ28oeVS
A3oElzO7yiY33P8JlpOYlWIHuUkJauJ1XS1qbQsoV369fVROoDos7Pj2uFmEUtEl
9MeE4DtOu92By9MAw98Da5rlUw0/Jp4o/XAPzPlc418iQEH4P2VOkGGj3k1vPwQT
AAZjNUUOClkaOjjXKLOk+3Gz7jWnJpsJCkiTW8LnpKp0R1CPQG7SkmDkGNyYP9x1
3P/85UFww9UOQeFcSXwsJVnq26xCUmfWhDMHhcrCxQQKjd1QBIIGF1p4KXLXguan
XXwLWDwyUeKRwGGopBlbverl9hOkpjupNX9q1uRbLViqpdCcvz+aLS5eE/x2Gjfx
Iz+eCHZZtvJTDDpKGThcEeuqSY3sjcUYKRfW7RR0bDvzkIxXI7uvOPhESdHVQrPq
sJreC6EvJTumoG933hS6vJxf+M4GkgSWzBP0guM3jC6ZTWapBA2pxGrr4R6yazLF
3RFMgSQK107Iz+PNtQ25MH6vBHcx4IOeWMfzAnAkns2lfm/vAXRlUueFzZKnuXOv
8jfNONHj1h/P9inh0fU+7kx3bGTqrBr/AhsKm9e/4L1vBPwuBfJWUBzLZKusCLd4
ezsYiTUCC5XwVndcH5R9peUEAwH233st0NwvaZyF3qMX3aa349Sh/dSvoZaiV2WD
+fiJUVAqGgzdXt2cQZiSdePCYQ8z+HAZQ/NF4+4Ofc19QyBfrNLZ3iMLCh+dHZMb
WkLARfQmGxXDGDd1+7JC6nmR62GIU53RaPZdzXQuBrqPubfF1Y3K8gm1we2emj6i
HSgEBYw9GPOfFNQfMgdGV3aTEZnLePuO099nXeRjRSqTkZJh8kfgJtuoweoZfuyb
dzneFBmEvnoQEnx3rcJHqkTcMJP6M0DuygAeQ4be99lhIUJGFjbSBRHiTSamce7M
8XiadprhTtX9tv1NhIlnOHXb97zEed5372DkOPaGNNhgTcnjv+JLNhj/MbycP0NP
uTsf/WVYuA9Wf6rh9HOtzdiwV08jSL4CPfMSyI2TWlNN2/DzH30jYza/b/EGXKEB
fe6XNcNYfN3qsaiH0xic21IEiwHpfqr9qmCp8hblu80ddzHIScjrVrhldUwu5kuh
mKIofVaF2A3KbP8ZbdrpgB5GoZ1JVBS0Cj41kLnPXIdEf0OwPJEbDVaMmLLPQImH
AeqvEWTPzDl2owxi4eBPD9+nT/c6v1adDj58cG+9utFiXB6lAQC3OsX8BPFb7bPA
uvR6JrMt9B5BKTSkhEk8sEnz2tRsfMbG7petBgtUVCjjz8GDOfyXl2ptc4OFYXwr
54ZvO7sAvgc25H72G1eklgcdEmEEqECt1+hUmkHo8z9s5ASlu4JaF8P0Rj0xLW7e
PJU9AldXSiW4bZWZLBypaW1jb9hEws7Gf/YLNlkrgbU6cnbjoPO89y5QWg76VjVv
PpVq+G+ANUcYuTHVfv4Vl2L6ffhuPYfQcH/6BLsmfaI80w1TNZj7sENcKG0L3FZO
6STe/REMBlJSpcECK/cMtG22xXpmGG3NdvQxHnEchRm0qIa4g9m/Q5bf9ZhsWDh+
bsFOKfgdxhqJok0pi4RioZD08MWFYyQP6caxx4PoS+anDfBGPlI8d8Alsmm5ijkY
H53EKmjw3X6UB3adXMK9OSjxZtGl4qMzBcsJ2gTKFm/v46eG0BLoWE+ZPr2hP6fO
+ftiu7480CsAuhVOYK6nEscRIbqMc2wl8/z71IqRk6gG46enGW7WRADoyWnG7yDZ
fda31oRi4nXLpv3pcwOr8kX8NS5uAVsYh+CDIKU01tNiMHjRCiR5OWzFeEJoURZO
aplUtKJ+/2XlBr+Vh+BQag5QK0tqhS7l3tawl/t3V+HsVidhn+0Dn8gw9houRWa+
k/WrEnTsn1WEWJqnOEfoRKOVfeCONmOFmHnx3HMg3/aDVo8T5JBqRA1zn36yCi8r
PoqEENxMiVpZRrz9RjJmWyU2cZJshqM94Zq6wzm8uhU1OpKBwfup+DchL+5pr8W5
QTxdaocJz2aR+2cYTHHiTCNM/d7iUGyqVe7Ba8jEJTSxu6ef54ywOhdIeEpDtfwB
ImvNJKqbZw4jfR2aOywS5byb2xzTlKSDOQghP+PKFCYzIGx7evXbeQ+pS3g8X+Lq
bBR6UqmqBNl65mei/jpT/bopeiFYSOLSiiM1xrF7pCR8GzDcZAZqtwUykV3ZJ6+s
zBBIznh8jbf2teYAtc+zdfgC7GTOKhzqxoX7UOguLkQNXcRoUTKPfBWdp7WxM+ck
bf6CGU5X3zARDikJezjYTkT8Gn0338EJEISFUsTzMf0PaFX17ilQ7R3V+G5Ebzbp
bOp83D/Ew7wb/c0IQT29MWBC/GDQuHXG22U1sg5Umy2oXqS6XQDuOjsSHQNtVxX7
hUFmXMroApJR6z0SdJMnlqgFZ3I/ZOsdjpkpYus64as8sdG/Gk9C987NUxV+bwjQ
Q9ICMCt/YpsFE1cXVOunDpPg2J+PEWfEdnuIqy8x/khWABRhxsww3tzHqQS+j4rN
Cca0I+X65bEbuAI69QEvSjM71qE8XtzeD+t91yzfTwLmHP0EANXCzpvRu0079nqm
cTL9xmmLzCKLy0HsCfwabr1KomHDf0eWN+S0IOHpXMT7F+2ZmzWPATYtDNVfOPYF
MaKfde0p8wKmpVYtpkv1UQadAhK5TH8982Gm8dvtaCkIFDB9AXUm7lEcGbgQRT1N
uW7EyibV5hKeJQGriCryAI6CYvx3PgJxTuxtecNKtjpdVIGD3guq6V/fjlB09Gh3
vVSrYRFOwnZN6W38AfTSUhfl8+WgoJNz38YZwXsPwhC6rFYutYYj0ytc9+QTZ54n
xKL1+21pScGQqqyVZTs6CxBcduf8q8vQwcgGrW+PJyEvFm0vS+9w9k4FLfgjVZhJ
1tZSSoI+w0AKRF4A/Sq9fX9AiJlG/FPmq3vNK3NpLWoSkRBsJ9hiJe+i/qi+mMk7
o1eOmuM24C+PCX219IEBhJ+kRUv+zfQnHZLNsL9jWU1h9J1RAJ4U13OEdJET+uxh
8I9cDfQCpVqFzStJQdelISOlicAAPcbbrPtR9sjPqvFUJer6uqecFK1RcGO2Mtz7
p1IvEybJFlEEqjYhZ+Beu9HiT5d7knZoC1wKTzCL965EJ0eXAMVHvEQMiCWxEpw+
tiM/1pWAtLzQI/migLnMs+iKzWX9JCjT9hG6yyXbxv12KEwVbcElCX3lChw6umZA
Z3AQEzB8/yyoLnOdGLwaNISfDRTdkwiztYI+M0yiSsaYMtEqtIdZ8yKPvDP3kyDI
twoz0RUaYZ+wnfwreyGhdck8AkYTULB4nVWYAp7R6X7furFJbLHW3IUCEihY40n/
12gvDpE5JiSmJh7t3Sr6i6y5OuMERv74hvemYBrOhz5YQSDRx1WFwLvdw2dm9vXX
GM8PY4zyfolmlodvKGx+1gNs1FF4V2piBEB89h3+AuQ6zSOk/VMwmc7/Ls6Joyj4
pUEG6bNGbhisunvVhGdIBxJOVzrB9SxIlSJORAu55n4hsoq83h9fcwVvkqOrppq5
/YrYGJZQbFBw0wp96iD/2muA8wshKfARUGjrJIfL8uRpiSeQC0FcqqKtgf7INIV6
ziSjhidD7BJyopWDk4lxnUNw2ChkIABNIg0oVVG09yeyaMeA7G6bICfwhg1a33ph
qLSsbt5FwM1eaoRB8CeXScjFO2+N1ktrsAlWNF3b3FTb3ny025GMdaDRNgJuuYvS
9AFmoyTwCCu/aQoT6rpZUdpfsBTgApo7KFET13OWyELtcMU4sALeyCTwhU3mVvOc
oSD5qcrKRZAPFHdsmxDt2qWVSXSbIfOOiVBullK4ea9M+QeSvWb90sNcwN5E5jV1
j9vMGq3k9FkDlmO6okGzO+P1zKPOWgt7kGaPLMa1IXa5ZrVwk+H8VBN2+8zADJih
v2u2wtCbXZzRYW2LoAL4HUSe+MgFJR2uJZy0SaUKB9qkvW/Z7EaD2Mhw3RGD95Ut
5NpppB/UdeU4xYNvzYil+RXOr0/DlELgyCLOdnYWVDaJ/4lxw6ffwWj9qeeOu9Aa
1TYmEjjJv3DCZEujdlSiP9lZCott+9PlLeFBGjfSCLgUjhcgVm7Y9nRZTW99YOtL
bmbLeKM/NohRz4EumLogMpUNH1e0ibXv80aiBTcZltHChz+WhF57D7F8BrNiU6yx
ZuY2Swio30PSci+2mnYlyd7MQ2XAtpxJydQf64htl4wX6d3XDugZej4C1Ksa/S+0
Iwn6Wd0V7DxwyTgv1zPLcDxDdZUa/ch4My9P8Iu2F/ZN5WJ/mtC3Isz7WgzuqNfO
/SXbshtywFvjmWtSk1oZUmHcy46Ei2G1DQf1JM9RRS/VMUpj+xek/bvez8tIvqoN
AQqbvi9WaIOvLr+Ioe9tP3QZjMAx3kULJgHTTaTarwvX0FHntz36GcEWqwGTJJoz
2t3tbT7IwM6/sxAl0CN37tp4/XepvMXaTF1zJOkol4BK42V8Py8vzQArK1dnGTTk
y+IrG8aB0ZTU1VXJTME8PY7lBh/mswWXBCaa9pCMGNZHLDqF2smP+srSYSW3jmLt
qZ+Hp9wBBlDpT7sGBJVsM3cClCfgg6clKYkNdd3mq+YIZSIXhL+wGbZ7O0tue4QF
5d7BYjfakOXnFxj1JuzLc7cSasG7KVveK+f8V3OWzZmFQg8DXA3lXrjH2pIWbqy+
3X8/SWGPMuUo9jt1gMfw3AT0t9bXG0otxuA2y8rz6srA6CxWQgBudll4dEhczqAN
zgRO09UqRg4eHjTOf/DeXf8HNzMPVRTW44McITcJHjvzfiUeYriKVBcEUUp6lBFP
bfEBpmrOvGFWy7JQ1MqY1DRHtszMpfFcvcyCqVdf6iuPIcK6rWbBXi9E3d2B9v2Y
TxQ76KwTjTkzga3kys0e2mUONskPMSaBGMAjMk5MfMgNdXEy1J9BFzC+Jq3IwZDX
UW03i01MlV7o1KZguZE9iMSETJUuTULuYnjgRWWeeA6ndCPhPaJhW6cgabgepf5N
SyrOAiuIfuCMCtANMSq4BjTZeiyYIHShjPec42V8CL6QFGNQp3SrAKv331h10rYe
12mI7YJWvEmAdOywaT+Fvv64FJ3yPZ/zplLodLKmILA6TKLlUmgZEM2FIX1DXiHb
816q7L0tN0pxdsrdNI/72E/JkVioR9CuwRKvT5RAtN4uvAp10dm7RXhyUndImD2D
wBjTUhCNDBEOsKw8Bb1RMiHGlFRCQGvnwdCsic9JxVejRjCAINUGP42ViSrmCSXl
Y4BgkVHEmffZc5p9T2OTbua53/vVb25LqmkktKqaW27yly9+vFnnfTml4nXiVv4x
TAHepx8kcgolq+Ooys1Lz+Vc3qq2tvTEVAoCyS7EKi5AUL7GfxW/wGRzMdpcOb4m
JVU2BbJNxgGdvVZ1U0RNX7eCZm0MHmjreHvGTPn82jAbkV5ygs+q1ZCPenJlMmkK
5ro1trSaiUAIvpjFCsvvrrtjNUdrjZsvmYIao0hUrGmQmVDG++2yHiT2RsAvPK4C
3bAH9/lY91N8iiE5SWwUMcy3hhEuQQv3oMc1ZDisA9iSavGTGATcNYJcu3eUMZZ+
qqOvIQxvtbY66LUZcEnqd9/qLwSVk9Rq7Eexl2D95YGTDVVta7G1vulh8v/avHjJ
W8uWKZ1jqL/859d9Xv7PoKrkZ8LSYOWpCUVs7uU3dVMd+T6oJCwZPKhQx+hLTFK6
KPV7+LjNqQQcvNTDn/qc5zyyYBLp5zJG2R5Kkp4JVGjvbDkI6OsN3D4gmqVfFUji
r/uH94yTTplBUE8UudrR15Wdn+PBa/EuuY45MvRpy3tZs5NK7IpDb9xLrRZXAWlf
vzg2nV2mk7u4+YNHL/IT8gM7fCbK/9kZoOt1U+t/Y3iLXnp8WSW9uaDV4yHlKwCz
+E0czx/1wu3E9A0ubxPLUPP1G6mKo+NhCy07L+IJjGSEHZsjMjw5p1iRblD3uBTL
wSkYspaPAyCYPMOpX55oILesjrw4VGtB63YRs8fIuIbfFp7+qIWiU84Wag0RHeV3
F9oUzf19SZlDXOs+HjkUIlN/BLLlX1QADbsUxkJ3KHlzUt65NigxFM2JCRrUis3Y
pZZirAQ3ByHKdmPdF8zRUawDnJY1T6Ad7JozlVLjKw6n9gdfk2N9A559ZspJjs+V
LweosJQIFPwXYI+GlIYofnSp75ihkkcXgbphHG8yj8zyG90ifz2uoBabeldPpIwv
YyRgureYFVgxFZd4onKMLaMkaFLl3v1gphPL1K4CMvKtUqnWuMS1Xss/Vt6VvRcc
UBuVNsEmgRY4Xw6WdaB1DLuAc+FzRvrPz6c2vSTzNnPMOb3I4ges7whMaEvsxlzg
qIWVkQaDZxa4kbnH5V0b9ErHmAJrg08xAo/EyFlwo6BlY4sxsU8kdifXub7GcQwN
pIG2J3HRx/zXRFdaIuYzVg41mm+xX16yGBw0+XgZT7yY/nOAV/3R1skGxsIsTiml
C+KFOVSlX5+t4jrcmILpWRJvPeAl/3+zGMTLAuK9P2JMbLU0Qt2iHTAd1kLfSTC0
qpqOaZ44MiY7JwXodV6tjrYjMpnCGlbJE496HXpjJz5g6DM4NP61MpRhdZafnwOg
LwsAMygfS8nAl8/IROlNTwyL+Y7bRlmxVsFRAjOB07Jr2vydeE+Ddk5RdDF1LKEg
kbgiiyN8kTMNo4BlxSwK8eC46whaAxOyEyZR2hzA/yaGJ7ar2tGfgFpjck3Xr+Gd
dpZvB6tGJ+Zm3/sQNVOVIzOkrUsLquDbvtkyDJY2/ysAMSTbJYN8s0vtsLc2lF+n
QK8ern4yl5GUO8fxK9oSht9Ry8wQYkOjsthJZuF8mbzxYmmE9e/vvQiHP7A9ygFX
QoBVQ8Voz9WdysCrCUNokuqtpI1P6NsNwSJy5pwZNnN03l6Xd+JHAjUcp0vnp4Hg
HJVy03f1kmMxHR4Q4l46cMYTs5Fc/xzHmNm51qCgKn3DODv2GqACRTnfvg3xmFx5
WUsqzQ6DKijzr32H0mfxf7BnLKqTn8mLDM89jb9mv6AAEQIVwW42OnR5QIAXGZqf
fHiAPNG6kqL2JqGvHTpCOIbJ7HRS5XO7T04leIDH/iFkM0vF/IvD3OBF4XWKv0Mn
qxiEvnBjBae+mlwVvqUesi3FUQQugGsVnumJMkA4uV3aMY6ZjKg4q9fuqs7ZTOVa
cT4b3MzI86euh2JLw3eGrM3GlzHMIhaNb7LQ5rJp1kldZwp/ToPwAO1pGJawgHE7
vms4HvfdhO3N6qasVNXKTz/rCU9sMnWX+ro6P6ZeKZetQopiyd0Y+geZ7oZjzUjT
cubgH6PnDqwZlDv3S6tDv1DBNP35bH3uM8oyqw7WoT9jGrV7OxuhOMPj6gNYz5op
NiW1leeSsJ972hLFZadrNCaqUwI3z9afcilxSglb4B/fEns6JAjvm7SHzDoq2S3g
GraD3JBTSuw5Ipv/RVPNh2rkfCp0ZyGGZNTlCmJ3vD1ONHkV3z8M7gRnJEZQ5VDQ
RjNl3URfs251ZzRdecA71W1AYGimQnD1xh6IaCmccM+SkinKZpIXCo/viHjIQjG9
YinrlpGNZBxGwmyHRGn1N40lxB4G4QPvzLrIfqvL/BA+61oNsjo4YdU8AmKfR53S
te6YF6BcPzzDFI2z0jGCgaLIlnGyKvBwAc4JunmGTq3UnvvfKzXfLd8F2Eu3hisM
Thy0PwRM98j5sYoxaHBpLBuKDlIBbbbAJScCbA9AmzlySA6ulJXrFVhU0ykVVykK
Cpz+74rHJe9EnwOBa2VsZmK4iRFvLIo96qj3ofy80kvoJnLMl6Qpa5FtlrzuyyNC
1ucCja4F3R9fmNIuecVlom7ELarioojsaQuMi9CPT8MFeqt6KNlkWxYcWzx0jvgN
I3H0BZQLNqzKPFIYOV1uo4TCEHxK965YS2R10cvJxqrozfgxYMkz2LXLAKNDhYC2
E0WDQAC0YX6yYoYq0GJWxGCCUUpBx/zRAX14X4ApJ1b6NOUL7BZT4mGo2LodPwfq
4Ta9itwhYoDPIu1ChvsYpp2KSDoepWQ9HMO7aflUE7mPJv8TlzaL/W6X/XiAt2+D
UQ6avvvThOovQf0f2TK1SnfKhyMJ9zJmANhZyguyu4EeEshu3gvv+tUeJP47U+My
LiGZuFCjg1eJVrFYn13huCkv0mb9Be7TsNL8smx2vHlrGHDgZLOA9Jgsdu24hh6F
AUXoV/M0R/g1Akiqi96hJ7P8HSh87FkwmEgQ4mEUXIogAOnIdD/QqSjWu2PQTtIH
/WSAhBCGhC772u7rTU74VeoAmxYHTdSmgaWGLMQfSuNkrH3Pez/WlyR+oZ69NGbs
s5TFtanAk6JAbw8i5nk0CJmfz/kOpnuyR1fb0pY0eVB/O/OIeRDitgsJKE+yGPAb
K0Mojg/Q5+yNf7TeazGrUTw16UF+HFkpGCNu22YJeXPU1LzO4rOHU6b+IVarN6j2
L4vovGCDKKLy3ITaWTRfysKBIqhzk6LvVBK2u5gS8pDxllkdXX5//k20lffpUMRv
hSGXgoEvpQr5M+Z4tC2K3MzfrdHoKDxCdmgPhmaBihCSDC8RP6C2BJAxMRqPJugW
OJ1PvHUI7vFgSe5lUeHLV659kHSRnSUhmP2utjzetRgLKiONdwO+vdmBznwn/rFU
OpdrYoD/6VnggyFFt3wW4sESM1eyW+ekIoaykAJ101YO0YwWXIwEFOscqlqwLLFu
RNkpGxhea+ixgyu+kgfqxi6u8fkeMuYNWke5QSVP4DEOs88HbNIHIgL36tB+tiRX
/runwrRwCXnziT4a6/A5GvWXG1J5mDAOssEksk/qB23TEhY0RXZ/hH7oAwy0IPon
yuJek/LS2IwM4JoVPWQiLkOwi/hZvwQEXpEAlw5REvFs9luiwZlg77ZX8UaAkFz+
lVrQcZyo5FsntQ0d/EjHnxvL+Tw2KX7HVCwHaR6k54bOGI2qiiVS415GoLPpNGAW
qsvKjteGox6JBEXi2RIk+ZgcOqGxK+jn8xBGWXoFIi/mSzE4huB2PDeWEk6PlSNn
uo6RLSz7nZdUCsWqwmn35KrD4xlaIKhJvoSCTkp7PTm+4Ct3w3Si+wJ4abNqYRk+
3DzSkQpfoLoKLRTeudQtyHnjqyNGjSC7euq7hBJRIeSsPZRNuOTJ+zmBNSIQZ8UL
/N0m4o7RADEnXF5/J2OM2VRWIE2C7fqVXGOAZOe4/BL8/NOFoGnKyjzK3opuRXqb
UnmmCU0JtqS57iNQjZ3ox8Mu1IiJ9A3zVRptMPvutPiQB4LUUdJjehbwjiqmFlL+
a/W8a6BlEYs0kVTYBREcxttpjSkEJLEkZIpCBk6tWqeCFq1Pl40VNMoW+9hHFeLy
xMSTov9yQqW1GUDM/NzHtWW3Jp9taQD8pHn3GzZ9V313YjWZ9aCCODNt4mUwlrF0
FDEQNbrX1j3Tb7T+17u9f1fjxuGaPJjUigpv5QTUr3NwdQZh7jP9GTzkpbj0g5DT
auLh1ebvcrweQkpFRKg8ipPylMigOdEoKe3aDlWG3EgDKOZxeep7IZ8QF5fSVyEB
/AGM3GmOpe5KYgh/zmN2T6vEfk6uJcRKmAb9JGYfNr+QZQhDdM1/YAFSfriGNIMq
nSX57I0swqlvudNer2Pkmm6lvXHJA/aKThobBAhiWHdILxRuEj2LggQf156FyynK
bfwRnaAbzEF8DNxtR/nGFEN/RIveuZq3YolnfySc2CFmggun/yb0dG8ROV6VEdhW
lj15YjVVvG19v9mWOhlh2di0j9pEWb/VhEBzqJvS3/VXz5SEFdagVoTLb0mRx/Cd
ROkf64y5AMogthYP8iF6xn6A3yqXP3/lbGxWB/Quj7f0wkfXDT8Ui3AeZwSRqfhH
20P935Yw6D9ffRwy3eRW72D+fJTSrFoaJwKnW/N4AVgMyRYUdARB0Q/Qiofn9LI1
T1zOuhVlwUNGUCKqfZRG1hLanumz38Y5Za/K/d8ksI7CO/WXsww+jl9bsrwKL0Qp
1BQiJM4vq9m+A5hxCjZeca4wZmWMOc6RUgxAAWESMGM04bAstZRmvZxB6jgOc0pj
9pxnWv5M+CiJQdxapNfRMhTFEMYopYlDew3dRGswU0gWj/MN4xuPV58SiEKXbPGM
tcq+k/oUgcWq0XpBdaCLv6ChhfkcxE9HE2MdwLafDUXKHDDSWxr840J6RskcBHc+
vQgCDjbX8hhQba3ZzNQE84SuTipqyT/wphV/C6nNquR0NLEMXdl/za+praqTsyKs
37DjSqGwyJ14vC2O45sr8EeEtm4XNtjHoTwb++hL2fTb+PsqsLc8/qhEIhYx5vhC
zMuTut59YXG4A9Q+qdd6E7OnpfWmu5k0NXHqDtYk7M16IBbYukJgmD9fCN8CkIMk
KkkuoFt5SxXYtPSJXE3MK15b6b3l4xIL1bwX8HK6ME+4fkJuqc5owAOMqZ8F7Zpf
XucdmgUUoUJSJCVx/zeK8Gsn0xwdX2NY5Qd7aDH+LzYiSOfsHTjkjZraG3woImuK
fatmUbWG25mbY6DIpPPQJyENKqVktea+G2xZg7Ed89+GKB/PhGfdHDlB4q2QjDqS
DhuoAY5Dx/ZjdgpbKqwIIe7gEWemGylIu4CieZpGZFywfuojt4Kv1rtRSwLSNgym
OOAv7+xUbJ7PcDnuLLsLDm6W9Yy7FUbVpIZyZMBLJc2UsqG1EDjA6k+jGo/vBqLp
6XdkpLC2WRe+HZXZ//B+01uik+lYrVGnvqO7DdvErk88Hts4KnZ8MlAnZp3uCW/Z
E04HXqvUEh+s7LSWmIP3HWfVtaQLug8rFru90UYssF3PW8JyFoVnUv7z5btSASLJ
8fwR/jtJuCG489sGh706B7ifr08w8CC5d7h6FHyWigC6xHk3m7ec3d1p/6FObYAz
tfuWNeOBV4PIiGQjBqdUSG5sSRbVB2d2QRFV4nZrOGgFzolfQTrXmwe4d611lstr
qXu4CHF7OX3moHPhuSjQsbVTKicEFYOhcuRm5soSZDdgvDN8L1bFxUcexMtT4oDG
/1am1F7Q+1rX8q6oBQS8EEgSTNMMTMbW8PY4HEm9iG8Hsj0YuGd7WWWx1LW4kaVP
FDxYmp62gTwTrzrvd7mzLVcCB5MniQySdgLXioW15jbOTIgv4FGnrcRyrGLkdftv
oGGuLLf5/N1bnQ1ljHueYnxfJaP4sKoWnGzJCi2vH3L3ntfZSj/apx/Tm7LH0nyR
pzjxXt3Xz2DVSGR+sIaUhFTysmyyHMYksDhQAZPPcqWpO9R2OrtBHa+7RVGobgVY
WEzk7EiGa7J2cm7xbonZ9HdMcTZys2ZeLfI0XN9zgXSb6JZRDnMpdDSH0tk6aeF3
6rlpVROPgQmCVhbnQzPHNKNbqVQIgGmQqMX5Nw0vN1TZ+BSeTL4ehSVhhc2SCDys
xAXA9RkWp2BUt91tiF2ItGYE1iWO605e2+sz0iHRLrs1z3QdpiOcXd7TOgmz9czR
1IiZ8w3u9z2d83g2ny6S/pGJENKw9NdpQFWrYrNGEIgbe+R0qIIXTjWoReV+EhV+
SMlaNjOeINNjVrqPZH6Kf5v1ZC7RpZkmbDZ5bhVmU4I06LXVQKw67YIPq2wrNPvK
JFNxKkHfTHkJcNyT10BLJR3xAsCX5kxb5cYRoCmYzKwZ/kFB2jB+hyriQPjFp1cA
va3AdX2Uc4a2jUtQu9SLvAPmR8NRFIqk59f+NKDaVsMwy6xAjPO+PZSvVuzxG24B
XxtWQ8zgfHQR77kEpEGstl2UH2fMHpvus0dgLAw9xeuFF3UQZkvMn2pDfdqkYTc1
DXVsYJzMMy9UctlNDv2h8SdtpoNRw4t9n/dP3jWOwzm03PFb8qMgCCdcI/pSN1GG
ao19ASPMS/9i+X9D21gZGZwIZgTld8Xddtg/TIcyTyLZs5QqBm97L1V9qqmxLBg2
t7NS7IIcbfoD4M8fgIIJWjLY/+XfQSu1Fhq1OofEUHDGTHvgeAXVRWqAM+HThJD0
djOYfrFx8UgxBZMYdIMn30v2OGFxbgFbTpYhoj6hsyPh6MLkmHk18wauXdbdNAFu
pcRHm0f1UAaJ55A7AXO8DlVE0aF0GIQhGMVy54aX+nQyACLRFe4/X2NpxjQC+b8k
n8ggnlCqns+OwP6VlEJZth2RCp2wsh12FCDdUHYcOljhs9qQLOeQSq4UGsAY9sgo
b1etCh3o2rN4+YfOgnngSWsX+viFtSClFJZarSXryVs+uYmDYPq0hgDreuLazY+A
XwZ0bpBT/aD0Su5v+7R7CgT7uz1VQ8zM4UF2wrtZauwbOMFNPRcMF7qcCJoZ4aR9
P+jfhnFk8INENiBKzdSmC2Dm8g0p1U/l2lVilhD1VyjgNd7m565rjf9+sCPRlaMa
4zYbOSrliT9xn2aKv2ZP0i+c92tA1hGT9rCbWR1uIkHiFVaFdezQpNkuu+zz4jBH
4aShnvKEuHhQhR4YXaPX9M2mREzvK61IqSLYPDmJeZRs3ZiKEZuqjpdbBeT6bYL9
jgRJ/kqQTHy+qqeAKjcdlrrJBB1yLA8YkCPG60xjk0fQH1N4sKgQET8KpXsNFCoT
7PwDx6O2MURrAF/Kt/p8x450DHrEBGfpEiigDef51pDdfRDMuSfoj1JCmT3fhoAZ
xSBnhi1g/UT76ww0b05SNlljoQDM/1anz/96pVQs9nnQafzwg1E/IpRI1ydmtNmd
dxoWrvW1BjG5E2rsr/g2TD5eYC/DuMybMNa57R/B8eB3tm2cXbIUcKHOY5lm7MTg
Hle07c3t9b+dCumDnJRkjDIZTh2CbmFmmCnPvBUpEnbbAOngitZqiW6tTwgNcvQm
tLaho7KxEmLJT9NTBFWAj3qcFI1OZAWJ/LVN6/IuaxJ+NI3jr5Lk6EvO1Dhsfpl7
6p3d+rtjEsBcr2BH1DSZH8nhEPg7vDd+68cFIL2URrkomtRQ9pSWpEfocj2QRQvg
JqJOuoMOAeURIOraPZZ4OSfQkf72S5mvLffTEbw8UM3bqXfaXjUjf7vLFUbeOPIW
RmP66R4aJMOxtgSq8+rM8aO+ep4x90ILLeOXOXvvNbE7cahl7WcHs50xyqIaRQpM
i2HQ3o0rpIzSkxrEwDLgJGLHEqOEPdw67P3h/QkHH1WhQOO0BlSwIu9yKy9PPi3p
yIhgWNQ43FlyVHN9J1kenFg2QLf/R0WIpsoykVf5IlRTl/8nwDYx2IbdZqgjGNSo
f5ygBashBr8kOC6FQSl3S2sZO+I7dDq6qgIKK8GCymRguGUsfFhDcNooEkeQPi73
PrOmcC8p8erkevWxpmlKV+vzdn7cNSlfkj01v92IRgAxEZYtiMycPDf1DpGu+VLv
xtSEDEMKDr72cIdhhpz47urWEE/TIAbXR/E7wPi6YsrFWXnGgomKpBlE7wvKbqmI
GU4y3REg4hHPShXNtq6MUB6ylUjRPChDmAVo5Cr2uiW7o5+7gsGReU1ZAhzvV2Dn
EBDRF1xgssTseoJ7Wez8s2DT7uxPWNlsfszdUp7SK8SvDfrxtzfuoF95S04uKD6t
S9JZDQLC2BNLLopYoK2NVrO5ovDPb5TJzlIaQpx7o+fjpU5mPJDDvhzyKKMhpKMl
q6kAKMuO2ZkcGm+W8y/j8TK/HzxaaO+QuWUtV54+GFd2s/5Turaeruk4uptGZEKq
qzotWXwfsST5ij7l42owTju5pl9ZtHOoX0Ah1MIGegk7ve6hoj85WP5J4FQv6zOs
u2WcwAXA/fBSHsErefa9Kd+QJbK2TeHUiv9iCkhjMOIBZGvwyMEdnVDPeofdtqBq
vaGcR6V1u+gnPqC0xx/aegK8D7L0xprUZY1bCcfaaGQdoAhEhmZdxm1JFYZFDE6R
VGzdpnqrBXTi4ZWmDXyQwf5wrqfL+QQUoz9gkyVpapMmxHuvBvPmdxeYtbeoXh2W
u2Y/ArL2ek0yTI4bP0cWvmL6wyOCqharjnLcUiF29sE1jrASGkn6hJvnIUIscGrI
mf6dv1i4iGrJjbIPZK/BHvdoyc5U5YhYFHUHyQej1Lts5ozuGvFI8GiB1IO7RBOl
FLfO5/ioF1LL1Vj8PHmzAlzRsURsH9n6rAHMz8Ci7tT1gj+SjdrjlaI2zYCYyJu8
J80aGBReFcOYFd0J5UBfbpyCXv5vAJGW0TrZVxDL8KvN07GxY+226wUOYDZfMpG4
DZx2By+KnTh3Q+KFIH+1VeLNhuFfU17CjEZn5ARD+BOC80R2jXW3VxmHwHZ2hN1l
IXZSjHwxtot/ZwiRvH9ptOlMmc8j66rmZW/P3VFz8TiT9NThj8rq7NfxDxu59RVP
DXTX/1Kl2Lvdkhfvl0nYdhNLPXfGo5bUCVsl5eSODkXBOAseKer7J9Bp0+jp4ZWj
m+y8HcsUMm/256z4pDXUxA7+N30rrkqIbrxZMFQkCf7+Qe9iuH5+hxddGs//CphF
eZJ3Zj72LiZyA7kx5Gx4wtYL5uLAzx9W0TYT05ZP6qjV8s14Sfj2TlwblHF4PeqO
5tZIt11SpBS53b1Bha6v6YzPP4fTwAseoKFAQHoVxiCzTqKnZadKLVRrnDFWYErV
1glG1Ur9yJUXfJAZBdib8rM29kjrt5xzdK2AoH+YyPOH8GAe4ZdFYnb0ftFNhamL
Beg7QbxJkEr64Z9zzyfwZMsYJr2GS3hMDIf15fYn2aKglq3IlzhLAlCEyibI+WGk
86qZY+ilJeN/lFx+wcY5EDEeRy35asX5K+i+1VdXrT2gZGumxYfcS7eAp3EE2Djq
Er9OvQgsER+utXciE0c8sV99oVkZBdr4+F7+2fSq12r1vv6Quim+nGuJzokdmJXF
EcyJqgA3RzNJ7iyOXBimSU1MGlqFzNYaww/maxtev4EnYEtY+Y1a4x0QXJ4NCPJd
i01z+u9pAX+3OnVUm7DF7t0Xp5lZ3Iedh/jvsi9RvJfQW0ttHZTi4HRO/cO8vGj3
p5LLIpWuy6LM73qkrf2A+ezUOPkM3qa8C5ZTQOz+fx0eN8yw1CsfIIXFnZPLncH4
dAbpdIumjaMSEU1EzaY7MU2I1OD21T39bIZFo8eVpVSqrFIyCDtmbDa5oYnlQ2kV
bgaZGevRsGKO3vuELDcgSfiIe/re1Qp6gPEly0pjZkcvAXexiNs9+7kuEwn5nA/4
+f9bujg/O61GRCUqbrtBtLB/RgHayHoVSimNi3me9or5h9OMN+oMuHynuHQOBJQf
eoXuVVnpnSfw3ixOhS6XyXhDZDh2EEz5LH2nYNwZeFwmJykDSggP+ZGELxFKAU5k
kVcrR84dagVJOdprXHRRNLNXiHeDF/8IHl6EjyqyyswVTjYCvEU1+DxQLO8OXqru
YRmZrIrhifWE02SUp/jMPSo0jwohCJvlKsGUr9zNOWWm7RnYC1V9ElaPFwZcuEpq
ux/T3FqfiAlbsgeMVhumH+H/Kv8xaPpQ2X9ohJBOzasL0DaCuN/Ike16xLWyCzAY
CPgWRED3iDPQM1aB2ckKg4nhStGiPydzykrxckPtsgqnbMOiWduWl6OgL+Uc5l1N
Za5FQTRc/a7CXK04boqJeivrBV14KP+SCBYwXpolr+zflRwhYwa0P3hOzqSiXKZx
GdMMv2ALqhWto+VScGstwXOaPmEhQ93pwiYUdYP3KLmHQwYsaEjQlHUSpT32pHbf
FGU+RaMIJ0pkIREwZm+fTR+bMIC9XEpOYXfcFbryBmtmttawXvcHLs51csWUXx0R
jf9PRBOTZTl5zgbDV5xjxIg/ahidWiWzELGwXpn6+UgvxWTA4MPgIQzh2X4cJADK
s+RnGyYXONgXdDsDoBM/MvOiZ7M5BMuwo3Namfkcv+myAHWla2hmUjjRGykOxIzE
fQzwMcsPlMkKsQ32xI4CMX1n24ldqSexKP9VhBAgsQWIVyZAhHfG+XCgsIGUyi5g
hhSV+22r6i9GgXld6ALAQ0jMcKxT++8KGK6KpFS0WgaFr8GLgR+GsmSHrjAdvaSk
UkHXzUFpZZubrAQtBSMbguxTMgoXzlgq+dmvqX9Q6wkWw3nRURhdyXD+RzL3O0dz
gMxqgpIS74TSv4WpDdbc3mJNXPDIuVDUOt3RlD50/eORBltciMo1tq+6b7Rm+MCU
Tl/QadqVoB6ldXLKuLnHXlOFXa5vo5FPPo2vfF+lHvUydRTGt85SpJTMBJfBhGbi
rE8q4oYPonp8r0Bq6nOn0ZsYS2B/BJeKC3vH/k6tbevKVokB9MOUfgtz13Gd7V7C
1PaCPsPdPuwKUwttw2SLdrhPapZ5HIJchFazuRhiZBHvuziX2MD8raqqZbvGesOT
ex4gKUPIi/6Giu5ddoC8XcJac7YFwD3PnkRY6cEAxlKWZj/S3Jq69z1Th6kcYXzW
OC+HrrXYAUvoNNq0Deugoq5qmpHSgzAYZMkLOaIrRSA5AgBK4qPeAUc4H8D5Sufz
p2T8PZEpM5GZOVNi2B/utz4A5jRAZc9TliMnfp9+uuaE9srYBV1rl2JR+kOyGnhz
KiYNvA2xG3/QUXOEaJzClTqZS2ezo2Utjl9UxVGSHsGxr6+Drz6pgpGEyRA4FRme
nz2OWJbrd0NHbcy4UinzcZOTbthoHjtwq7SYjP3+wg+Y606DibDOGIewi5NmHB+U
erRkyPZH5FQQHAKLV/dZJQaC0c+luUeiZdOLPp8q/bukpyp8qzcXwV6Qw73rCay5
B3Q6tyzlrECTZDxJKzaLR7rxHfBZsiEuUuoaMSK1YHMSME+jPT38A9iMYWedXcTA
TIH0rXTeKEw4ihmwEe5HXkcQaV5rFwTzxrx7U760C55dE/ga9BKG+FAHop5+mTKB
RueBcPXqmigLyZmuZXI7NOS5Ud1wc1xqGvxqyn2uJFnafVb1iVDzw91UPeEdDe+G
/U9lLRYhd1qfR2eNKDYAyqV8hLBK3cqRT1Wok85G6+umOKX5OAHO2IHNpHd5lPoc
fzPebT/tTpnMRrElO9mMK+UItUBgZu7Ti4Vzl9he+rB9e9SERLFQHMqNu4QznLrq
gWdgjky27h5a0Y7zqAmELPK2aohwSXvUxDhz/cnbf442yFOIoDhoRdS89bpK5uxG
3sSWLHId5qJE6FOahC2mJjohXRJUkQWzmIOqR+yI11LFAXpJ+bu0PsMqYsx689wg
6fDKzt+YI6Ctkgj4Q/M/y3UIrGY1lPznSwTUuP1O/i1GO/GY7sHotPmJ3+oUipZQ
XrllfzftAcrW2norUSJ7ok7nEU4NTjB8r0x7TzvzcsddjXgcevHfl1yDMfcqfuZi
iVaiyUMH1Y14a+yIkpOuCvoj1FZxcWZRMJ/wqGHj3W61c1x+gGprHXSgL0nDCCb1
2IzmM3JbrVGBMsGZMxweDzjYmFKfOZ6tmlwkQtqu1F5Sm1wVKe+J6eDzxYOoF26f
ny77ALzTZCntEMF2jPH/vqoHdqislYf4JB5btyswaixKGdGoloG2vlQ3b2AopiJq
8/r7L4B8Nu0JwSm9FOq/IXbnTg+Ssrw9iYfsbQAisSDb5+Qm1JyuPqdNLPoPelfO
UVCw0ZO9wLmzWm0BMhatL3BskgKZ11iZRO+S7fxNOKbAVMoPKMu/oRfWDiyp6Ob1
pm9+O0qVkgK/6GYe3c/xq8mpjNDuKLxvCr6DD2pQ72zQiu6bf4U35HdjLdv8dEIq
iOEX7l9T7itom+oUkE5fHZEBkvwAZZpXTLrTN3/gcI5saRaRQfaWS6fRYMI5G45p
WJnDa8kp+S4EYQJ+Cfa8Tholg6QXkg84cEVyoQ0mohIQcm0ZZd50Q4V8IswMl+46
DLQf2jtEj80JySU5KtI6qysRlXh52CwwMkKlhy6eZ4UZb4wFE/Hc9TlvdpuUHFaE
rRS3grt/bMT4eAN0JKEmucPrY2jx0yICZom3RzE0ZJd+nMwyNv4w2mCc+ZX8+ZxU
tb/y4Z5vjUTgnWTO5S43rjF1Hnq+sxkYw+hJLwjJSEt9I1fJFgX3fwEFZu0vdDB/
fbdKPxQ644oZkbW9o7FuwHzW/m3Y9JlcZe8V+z05P3vXBmVs2oZxDqa3g+XAq+I9
KawwTXZaBMG9b9qggQ6L5l4MqrXtezczIJimZuaBrV13/+m3bREWUThQ5143MTkF
nDFctL+RcMbrFmjSOoxmQXdrjkBZcDxOuficzSrveVqeaQnP+5odH/HLQ9R3Sx8o
X3Kgrf9LJTpFmoH6pkZEbuETNR101QhVEeIzHTpDuIC1RZT9vBJxOOJe6AaOX+Dk
vya7pAlpUPRcU3DLp2shVuQ/KpwvAJw22yI9mUAoKVEZ90jKggNFI+ND1eaut8IO
nU+AXR7A8tGi3e4Ch4oIX317mt7jNToJz/fcZWeTFFfG2gJElvmpmZzrE+ZfwOZU
TZWoJIlICWhsPvsmuMt4hRZmj5x68iqB0+RjfzGd018iEZSf9eBuf0Lq/25uYQBU
qzsqpfTbQRVNlQm8LEzse8V3oFPkvV5oM5Z9xICvoI6I2ZFkkECfOXOAEyos1sap
IWpIioqD026Q/vM4aL1+crerSQwxNlopJPV+3XvByLa1ZcMRxoOEg5kLfYtT+bul
eH62lLCoKY4OWf5pmI0cwynfDCuPUSPGK19Oq0DkUgcb7ADQQUwyRYS3ML6AcIIe
G89+Z5VFyPYrFHnzp45HGsNo0EEh375P3diuv5DFjib4P3FI47gx6UKFtQ0iZQHA
7Uks9JXcUgHE16eelR99G2991g7JakdVJ2sQIiFNquiQ3T11tD+ioVwLqxBD1qPO
2ft5AQWLJOynCMJQqRTpouWV37QEIGyd8cRgVER/LjAH6eVMwNWhAICOiz5WxkGM
fTdiPXNB+uvArtuWv1sz3/Myr3RCDeB/yDtE0/+yk/h92lMJ8RKy/Guis+YV6f7R
qUsQTLCvapj+AsjuP81K0G8wPRfj/e8M3y91ZO//n6BVmG+t4gi1FSDotGzzTZE5
arIAocu7zk7Xi8DO5K+t0L7FL+lbRm+KoA3d5OyUKGHzauCauP8I7FRqnK5ZAK9o
z9Bnkm6qqjJezR0WqfFDpnogyqqwZyS1FUGlttlYLBnCZli7tz97MfxDlajHivDA
FhmWo9nRZJYAkUpAxOIo0f+FW2klY/KhTckPKNxfkUP3rCDIHhclLGrmMTF2mXb3
9HjcGm4X3HtGQ1ALfK/t3fpAZfHBjjwtoReur2ZDvnIsW5X88MLian8E7hxA2iyY
FFbPhYLd8FIYAM+ESGKLhv9YY4/HaourWjsdyRuCO1Hoyfaq1TJEO/z6Umsyjo8c
cgB5z5olivFrvN5N3YmkPDMnheN19YF9ooT5yJArZJZPNQbzFtSpIqhIfKvtLt1n
K1Gt3PASuOnBxLzGJ3ATxPICNKCw1fuHX9OK/u94LiwwrI3ZOMh78IRHBmVNWA3x
XIFHL6t+1nPp8L0dHG2m2DWW1ZcnsAFwUzT7RCL2RQjkl1377xVufJo3U25BWu6a
1RP/F+xYMWRP4cG3hVT/8s5w72N77YnaEth/j/HKbCPIkW3AxHMgy6kd6fC6vWuZ
1xbfi6QW0FvW0qvZNhw+X/WvEVcTucSmLe180PDxt3oYvZ/6rrx+Ua60/xg94ZE1
uxafGnGtFIDWy1KaG+bSMcdXrJn4x/eoedDTkDFpdr+jfnl7SxZDX9ZpR5+z7CV5
dz/4t2or3t9Qby/0UnZIN9DuxBd/JKdQC90xh0NnjbT5giBTYYtsTK0DZbBFfuD8
eL3znbpLR5Gu0nXQCMJaduOD8Mt/j9jBRfFb9YDv9bmCntlakJcIGnBZuofJDpxh
R/KK74Yx8N0BPcaaaYFtIrSq9RRoI79eo6hOiEn4As3OnD+9GDMT2FVuXxcVrhWQ
tR3+/CuihYHOihWCfK/qnTvhkZrzbtAJlr/zm8iarZ+CldHuHzUROnNQPCTlPPAp
FxAmDJAh3TJsMSuyFNuWkJl+Ok2XSKW8SZyEP/EMd+fx2yiDf99NvTjHofaUVqUy
p4z3E4DcswFeo+WmBCWBgMwqWoygxs+VBMmdDLoVFBGN3qHTv9Ox/G//WqkdYlv9
UT9JR1krulgNH1nKfiQbPdnY1TkwENzleyUPK1a0cHvr9wvuaP8niWPZzX1tIh4H
ApHQEAQ3edMFJjJcfXDVFoinWcoBtFbsR8VmdaxI7MtaXUY/823O8suFm7osqtHK
d2ehHvPzGZLPgkRnxh/v64VnivjleDrbXF8lsksN1hWw4YC3hf1tXOXIFQxXgRhW
CsiKAfnHR7ub0PIw2B/Oo6PIWrMzkFKojeFD9/s+z7dX3MqUhCyKiAAhDC+Y7X8t
Tb+5rcOmrSykKolAZGYWvHrcKlMLrl+nUo+lxg8HCAsOzvytQYENXCuqcbB7M12N
WZCti7x0uhKJ1z9vcRWEF8CLzr9hVYp241Cm05PirZ4aWop9XLC7FgnLVebHPpLr
iZKZHWppku+Z2Jp0o6nRVgcsEv2c/jjfUAaZvNzY4NKOgu9Vy5dT6FgAS0TRknVt
xFluB5O5CMDzCaKYrjfscJlr0vJwd0KrCbndyr0Xf+6+2EZkt6AQBghWvQmnn28g
6FsbYbxVw/mC+D5PoIIEvi0j54BC5SQA1nSYSBlngZBpBQDB/tPeh1QoCcOaHlNb
6am/sPxIvAwna+OE0D/QKdv97Ysbb+fSg0bBE1rp+GqmbOFSDPpHUO5Vc/xeb8+C
2h7ISfaCtvOWULqWBk0u9wDuZAD1Ita8xmLElh8tEZlh48mBa1gnYzEivLJOvCIm
z5AYMAVgWvgJnt5wRvctcoZrUr5rX0bvOoOYltCG4IRZKQC14gLwOjPOL+pFAC2D
vcWvXMcSdfr3pj17JR1toUTLI82SC/QRGWSGPy6MEHHnYHtB4mbv4bG+mAYqt0QH
xC6Sj+Ta9Yfo5ErrYieOiJ5mztcaPrrML9gm/n9JeedLZVIsMpid1sQTGCoPceZT
aoZp3+qKLbpN9VGxwY9UY/XMaF6/55A4qqZfb8X7kfRT696/Myjrg0/VNGN0alUG
2k3CQgU8qtceNkZVuwnmw01p3EUxrKdh0SiLjQcwh+nCtrBxDCGcAXix3I0K7XB5
czIlAFDXusHyDiTm6u1Ob96kMtEvrZ8ukIhsuipu4cAcZzRDESezFKS8F0PcjjVk
oaXccfMBmuTeoP7ibWk5DtRx5UK69qePOIc2RK1Jbv2y6OmNXv6DJ3qzc0gIw/ZG
tTP9rVjIAs4/uSGZ8cV0rS5zqBzb5xUtmou/V3Vpp0Qyn9CADP7zFOiDnD6jKN/H
POijaBlfqhrzSPAtfDk+ZO1+V24doZ8D/eeBUXOvIiSZ7Vv0ZOwDjuBj4dpRyZK7
zTAW9hwpSkAAWsyO/dsfMqASXGTv5XY2tE4yhLgE/R8GnBIw7+BOxVSXi8tWIv7v
6vD/jFEWu8+JPTJiprgVyWfX4JztY2lDwWpxGRFAti7b65iXpJosRF1Dw8RULTbF
tis4wqY0bK/pNcTSGNZRuov2cdYHZ8u+rRr5NM4kwJ/W8RBxEudTn1p8fYiAb8f/
O+bqGr65ZmpCD8NHx3YM1JQi5sJhxw/T6EyafIuaoh4x2GjeoTYD1SJCdngAZljM
QMEHqGZLB/QWpT9x5glcvzzwVjLyeV8/SVz4nsh8ujLdClcqGu/SU+REcx5CMRnX
QpItv1ZJALH2fYD8Sst+HH5lt55tq/TGZKoKGvQaXAuIg6feO/9phL3kUoRcrf6f
n1JU7hGPOhPoUb7MQ9kZwB+azSOXB0vyFiovUHu3JDbQy+H+Z0Dk1fUkFmgn4Xwr
nqOYaOsp27ppi/nFbinJfvNpImQnOZuHJcugN6GLAL3WJF4E1C8NzBus+KAsB6Kz
g1nXTr6g70lJEto7HHv40S7v23GM+L1BFMNrDkknmm3DCsd8l5kyhVpWoH1rMb62
0StoktyB8Nmpn2G1qW93yGRqZ2D/zY/Io9040IR56DYw9JYw4t5q/kvJRS9zRyNr
ZknuGBvTddbNyfQ3XJbDFoMCAMuuE2tk13V9Jb+G94xMDWMWizJ+B0zF4azLZ/Vd
rbOoxrX+EwjI2YOaQH3jyBGGVXyuWo+AzcYT4dJGVA6l79NTI0ict4NSEA4H/oP0
JJYHyHiuXPfFsGiuEe30agTry5nHeWGC8tiRcKEIXxSMrcoyNI3L8aC/0o/Pmf/r
VFdMZNW6etSQ+J4ZfJ2UttVAwuC/SDT5wtBciuNze58EJq7wmuhN9DOwuLzjTb71
wAhRdPw33xgx0U4bDqspdEIXYvfxlsNElw0U9kspjn4MsTlGliFAEVA4ASNpkuoU
QVZu4s1T1fc4Dk/l2tbXvcDhJbiyDPq4bYxiOXQRtljc370hBUxXAoyStC9hgAQM
giWOlNj9pBCO+ulUiJH9bKq/pH1GFYXDOyeHQJDyJqGahAn32uCuLd2IgljJvASe
dzny5PRImKK8zynMIQfjq0/sSNBjfwgkp6LyFzEAwsTnsvb4eeYDWhuOhsttaVoR
GqRj3G3/ssNxdxoSLArQmB5NyDuwy5TBbIP+Z9kY3h335Ei4MZWfcBt/SjgZgofS
0+0FHny37oxP/d82rmmCwjvRLb5YZi2DSMdJGFDugi+7t3bcNJuyJ8r8MlXPjRLw
vns9kVuP/yz5UqJJ3V8ZYgmiU2jPnhVf/Kv2nzva/4CMoqQ8RCpaqTdjIPQ3ia/J
cBfQV5Ysfl814XBXzpzF4wH8uRhISVI5H/lOAppkeH8wVxypuM4tFIVDbZhfvxIi
N5g0/4ULVTnzzskFIzO4rT9faaxVRNNu/p5bmi5/tVEspdAbYwDx1ocSRB9TiyFR
nz/DI4n66kvF4LeZtwnMhKu3rR+Qjos14JAbjM96xYwftX5mRtO9F/JbHpum2fYR
ozfgWoGU2hnkZdq/GLZYjB2V08VQv7iQVmVbLt1BynzSIwGHrLJQkVqLpAkAEUZJ
AjyUgtAUqxwstSHd1Nn3+2u/j+SaU7blanyC7OhBpXCuUTeB7z7HTkrn9UWfezz2
gy7LoEv/ygQxkG/ZElGfvVCyW7+kWlxFz2S8fXVeEFf438flRwUgGfFfFVSPWx5d
gS7rdj9Ew0KONb+oJZqOH83DsaUwzi2zjltSUhvEi9ChlYy6Wi7XRxFQs8YJHEIl
5IYY2cY6s/YAY4OxDhM/Wwn3MMg0UEJ1fBaAQ3QB98rqbwWzdnivBzYWjHCFkDuW
KG26tfjzm31A8V8RzU3sGWrDWg3yWfca854I+1mGTM4M40BivlR20JNUemx7MxFs
6vEdL/znnX+cg6dRyWlr6XV/JIgzze1DazRUb2Y1Y1b8l4OHGWNNsBZ8UlAiFZeq
mANSGMeoDDFyTyJQ+xrJQFnEFnYNhCV8dRYDL6RtoSLzCR9HCc1Ap5EsGFzFYj4n
vp2LprxKvx9tC5xa1s3Baqax+5UhVmGmdM3/XL2VKNW7GXWSoovANvBCCJJ06qvD
VjfkbI6sMWwQ3GTO9us+xRJSsywivd+JHshVLIrVMDx/MOiE51bBj5Sf0KQQQtNn
hXtdiJjkMN2+lMEo4Y41JsgLWRI5tmKxPDlHfaxhCDuCVjIL1rd/rrBBx6Dufz9P
nvAj2blTDdsfCu5zntbi8EmnkBOTjNNS7H11oEaG+uV3YStfE8FfV2OR9ZG//VGa
i9GsIXqLkVxQxAtgTxl6raUSRqwioM9HOEgRXVmS6yT8dWv2xh6LqfKrq15yFUvU
5a6odwR1D1VfPSnPr3SBn1k/qfexFRSVlXstA3ITTlTF2Xxvlh+Ph4hzEh06UUqp
xsFyUKDFtfzAsMM29/5A5ZfVy+Bt35AAo8kreJ+FUSdxi+O7BkgKx8/+OGPqqcmP
7mNJPJIMcbRtNP225JeFUP1qregljOYNCLtYQqEQXRP42oFIMbAQkoE3cA7ZroMg
S6taOKF2adtD+ajxhrm7JahnQKOnzaYurEI+iklFMmctqvLzEFU3D8ydHXlM6ADx
dRjCBeAoFkubuOnuxYyF5tK+/AXdslCbEF7dAhTs1oxgL2rXVze/4sb4Izf+jXbT
xh1g7iyV212A3fUnmGr8wCHpDHZFNmfWndxyfsPusLBl20R5bmTrtGZXneO3TV4i
KVXM+qj8d+trcCATw4wmFJOJ7Ve9Csw2YalLu+v8vAutq48Zrz8I5nUW0R3YBZaX
KCljplenuT2kocDJ+IAo2s3HKj6BSGHxdW1PNKoJznCrxFJMMaU3sS9yZnw7xoby
Hz/aKPG6k131ndIAJvX50TNe0cFuwo5apPHsl4HWcL3Ni1VbXklj5NyZ4AO6w0Ov
wZm+zlFwOwJe2xa5i9vANnjbTXvKt8NBM6NVDYcYzU57VNyXJu1vVPo7W9J80fdJ
43iy0pRlI5ib1GwCKHvUSCMEVIFRGLHwuZajxT4+AM8TtxChT200vAa3xqGjBQyD
beJlhDUDlcp40c8Dc7ZJn8twK6SYGK36jAvgukUrHXvOTdM+ekYTykOGTlpJCiwW
yYKdsXp7f7upsqG+YPmjd5YgZTpEY8G6AYtUll2T8BRb/FKNTp+8ngJrA2Zdglr3
+CC3OACT66LvyD6ENcLC5ICz7QLJYq9rsdIy/3ueRIfeszSD8KLEl0JYZrXAk74e
8Mu0/dNH0tkWu2IhyEwE6CforiC5dd1ro0nXhJSvkERPviNzJvZsmBAbeENhg31Z
7eQoIDIRfAl6UmUsS0f1AYtyeIZq8+vKoKOpUpEYDkdNFGHm5TFZz8QSwHu6U8+4
ZPSrm/WjEmAUQ/jEIynurfhPvuHhSW/QI7x4LLy2iSvZdpWiDOP78PycPVko2L17
I2k/hdlhdaLkVNbNm2zc51QuhHZeoZWzb1apeKbr97FEvL7XUyW87eBnwSWYmkve
kbV5/nR8alb2nWslsQIrvmp6u4gjo+x1+jl9rlqbz+bO9cnqNbQZPjAl5EDT0SPj
UHmGipkadWy/YaLkIRp8b/KqYPDQHoU4hk/jOsn8ycB6DPd/gcgoNtozJFbcuOaE
AkTtbtfnhPIqGE39fRsh0IUWk4xBHu1Iv//lqFXCl6kdkdqmmZFyLbbXdbOSrAoE
VaysSrD6GwSv0p1gS0373ehRhWPexPs0xqsc2AH/hxFDuo0PToR4VdR7XeiwPbSq
LTj7MinLblb4/wOv5FcZSTSIQOXQMwqNZagwHLKySug3TbzdfNkzEMhaoP6U6fMg
4WbyPK04PX6/NB+4wnyNN6PHKhfPwSdkircE7dGqDj/cDGfKlRHuf6j/Z1dHJp+6
DytevdKarspZdiJmIF1QojtscMJVloKgf/tUnplIBlDZSnGWD85mfuL63UhDpZ4J
yHQNE6wbvTGrtiAvre7C9Jzyly9JmRfn73WZ4GnA5NPRngFdkOgSPQa8H+2h30qB
7tPa+0V2OVniqGCnjuMj1QljCCidahV7HXbayiTbAzU0rpMYsqh36Z1Zw254sSBD
2Rf6ejOq6hYNkky6QCF9jOErOft0VIgHV5sMV+35rUsb86CTRCBlwLr2igV/Ok9M
5tfTLHVty1D/KqEU/VJwAzM1DFmV5qFpiqEK3T/Ge1iL3Vc77kzN88SJYr0Nzm8e
1dRR/I3Slgbu2XDHI5GWd65CV49LUfxvKa98sWmkDVwolLbswz1sgFpFqLTnQA2D
fdt3yJzoHUdIQ75j+AWPLs2DPWCJw1XqEgzaDa+KIu/1IS30zoGUXUN0hcmf0SU2
zoyIoaiwCVNLb83gbvvQmChwS87NauoseNncP91mjTG59DM5qmZk8JqZbbGNiWVP
TlSSr+gMzCmZydppzJoqtpg5mW3NZ0xm/4XUnA6KBl3zOMZ6+6U84I3pfm6fBY2S
SQgDFdMmCWzCH/nBMyVULFMisiTMYgn2uqy0JR0sFaUczMfvhUKuPNmZId6FAFgv
tJ5ET4+ZbDbzWKZiSgZFpyzumQ3BWJDRceeU9ymWZYhrlcUmOE724pfJnP29uj5E
LyCFq1Isykc5i3Kd3LNuzouXQrsigVbcNtzD1DzrcauIcS/eXDo8eiQwaH9/SK92
Y/KnHM5M+y9QnILqjZbO34KGWWZ+NXccmcOxZXkG6gn6Y96dCNeKkhTjXzxcPUGi
z4oIifaISBYq32o8MZ3ofu+ZqnfOcVO8Fs4OUtMqvqSvAmyIWzZnHSIpFLdmnmzn
5cVpTIaVUh2+Y4YKzlnogxilbNJnwsYDu4JFUlO/wX3NcoaqO3kmhI9uq0l0SuJz
1n4uDQ85TZlRgzR+clkod7Gxr4syoAdg5YzI6qMMBvPaKChEM96Sl4YwgaeTj+3h
PtqtaUiuMnolKW4aWDrFar+XDnDyv1KRCF1Pb4rwPFZN4bmG2DHS832DTfsLa1zL
iDPp/MP1o7QzJSPb1Wq32qMj6B7kNieXR8HdHQ12zEFtrNCpr7WBKLWDo/aIA0Bd
gXEmsXrI+xFBawQdmJYeIuaGO7gnKgF3i4AvjNMDbOVNUpzLUiElIZfLlYdMUTrK
PelYpTbihna4VSuHi8v2bX7JHMGkwT/foqzykAkydEEkW2i4j2hYMYxdnwwukWxA
TM+jyECsliS+4dZF19zNJRwuky8p3+4Ads9aOe+RghXkeUBN3j2Jle3DHrYekK3R
gHRsMYQeyT9/Q2HiI0J5vL4fSdsiMvCu49e7Oy5qa3DGY7FwuIcGB+lkNZhNgC1B
xZ/ftIqe3HMrJFcsaXVOJEZF3jGmycx/yJmAt0bYxpmc8F4ErrMDwpBP6iYaswEh
wgX5fyw98NqXIBHpslq7exs/o8xTjqdmaW5zUPQql8tZVzOkwHOiUjdSSU0ett4U
MkB8HDA9Iu99RU0jR7bYti34NmOC77iOdojxttIPCdaBEtYpMZ2049y3NN9PohsQ
k7GnYf7FTFrn5pbikCbWRu1bSU/p9Bg3Q+S9L1bUgVyKEcEA9SNBN6hoYSrIErHl
qBXAhMCsRu4gFm/HEU1I3SEdjSmTEjTgHqyM3zc51UZBa4Cz1ARdSB13JBLphLCH
uN7+zJhz5Dvs38PrPAvFW/6lmgkQrMTAk7WwwVI03PmCJ6f8XR8FMK6BQi9ny7/D
02zLuv5Y1PQ8OxKPo1xyn5v+myEJCLEzuezmsxWQ7mw538FzbYCuCpAOJ6mMVuas
vWBVSVzmpwCEmsyE4yVAArQT6FKOpvNyH3YUYlNz8G/OyM4a6kcZDwt+9gDHDl8Q
RJlnXUodDkmQKxLqIa489kG3LuiGxA8Jnl7udergsUdRjWwtJTYJT7fr/NfLB2C4
bomZb+IfD80tSQ7ikgUXmM9Jr4UbRM6b8cyjK1xcK1PVrpzWGRZ69hKLVHVQZYXV
IKVkGD3LsBenVC8fxZlC3F/c4PaeTEWATHJxvqD4vodqNkRLNOq8ochD4RZM3oIv
xRtAohJiNaO4VjZEp7UEpe4OHFDLk1ICKxFQyALe1suCaRpQd8JPoh+PpUFRL7/3
WtNjc3YGeAjsu5rrbtKzRQmFlGR4O9c9+Vjc7YFeCGNRZEywlXMJ24DJdw4JUH9s
PoQ2GEzUOFlmxn97+/FGm0/qni2lj5bMErVnw/QYMr+PAgqTvZa5AZr+CMLGf4IT
L3yDJ17A7brH+EiaCrNzEU98XKBYAhBpwOX3/YX8bg2QyECZ4FNlZ4k2Skazcrro
19xeNtAeMOeb8pVUnhN18DXwbGqKv+Ad94fIP0uTp9caghHnr1Ipan95sPelMkzW
BqFospbBiiPEvUJRJax1zPw7VxXKcfSbFVDHt2S+l9+OTHuZtuWJLYiFshk0OkgN
DOxJB7VBCC9hPWhZBO0h25rcffB6DAAC3HsOGk34H0uuU+EtYhA3nSdl3o522p48
2R/6mytEy+j4gGhxFd3h+8XLvpfnWA+WSoe5Rzrbdnfc/C2iGMEc9D349E7ekeIu
vKSb15HoMBh7woavvZEh0M1E3Bb8Jnm9n3dK+7Oa3oNyo/chS/TVncUsAAiWMfFu
gNeB7/CXeiiKcgY3qG8P8L9YiBw3HaDSTodDiR/DngPk/JqBpFfKus2ZEJP9aRvk
Dus17EDfVaN1ropl+W6dkxIcOvNg4iWieI5kLp9gDuwIkEfBA7VALVZtluXB3Lu8
iIpAhwn9XkKi/CLrkZSFTB9I5ch08Ebq8a/GgWe6NOUHEOeNhGa8M+WA1hDlM+vZ
ga2H90fUkeei1AkYnVcMNVbldgIHd+mO2r/TA+jZ+2WHtx+ChHkWARTjicO8K4fB
nbXqUH+SmEM+M3nQPuE+6BY5samuJQHfirwOvIrj/aTTyTVmKd/925OHsMROdfa/
OM0bLBZuTaHLWANIs4m6u+Cxs5dxgvn2W3yVi0WoYGPkbA8oRicZ0lIKQKHmaBgG
TxyiiKoLXmbaSIQcbLOcg7RT7Dg6SjAa23Z4dpaYoLodilIeQ/wLKqADVKBxVHbv
gS11WE21LlIResOKtCMueylJOP8DMVoSKDSZk+r+ldoPrlJdr07NgyihQCKiB11p
inTc5+QYb4itCe3a/F1FfewkoRdZ+oXm9WcuOQ6l2TFKSyHl6hTG91P5Sx9YP55y
QSeIoZEToZtF/Ravl2DbbL/KXIEFUFvQ40/Do6N1BGDiEANKB8OmD8R9FoDzO40M
60IGV1iTdjYtzG8XI3OsOwobnhbvyHGrFOiPqWDivHtOccq6jIJIJ4tXOlDZv6jx
EsBqKogJxR97I1dJyeuNxFQ3NWugSrfoFPBlZusL6/1OAJMF5IIETku0aqqnegWP
DeCWfHT/V2eQT18Q76qjckPXLZ27rIMnYlMiHEGcUJk+hc9mBZsJtkUulQ2W0ONb
JjhgZez749aY21thLq3LFaLJmjEK5R+qo1G/02GyrwQeXSuRFQuRVN95lzYGEx3f
WEAMdVgO0yOrB0F51DuKbB8IdC9V1sFT5bLplaSNO3SS9+t1FCEC0jVI4Cy4eSaM
EeWyhQNzOimEL19/1KM3Kz97F4B7iallPWQWbTc18+0t5fOCmoD+JuDzfiNT+3mE
rtcVUMaFIJnG3/580t+eSwSe3rvGxS5LMWox4SBJbL+bXaqK36uSjgjgGRI+CR8v
WHlv7w1+OtpZAYionYxN+ByqkzJUVHCJgfOBHgXp8ZxL/LTDtQOxWcayQv8V3GAf
anX1knodGYCQHfIK6jAZO/lLu0QFgR/GvE+ZsTKFVkgd7q1xS0ujXURZKHftOJ0a
xQo20IpxsRCf8EV20sCkthGjIVYI2IdzLUnFfuvLtVwkRCE66fvJj5xCxrIbxCGq
4deiP9849JUxGFIvb/ea6n9wIGxe+5hqzORs8h2a+FTgc4gZsi6JMzbtpJcUPb86
pysd9HvnekesahgPZQy5nrkcTVdtx7hFxxJnzjVfUdoiqCMJbh9h/yPqstq0XI3Q
LRprcXqxisKTbcV/d1lmuS+XirifVTD+LnwBnnYmzHSnfyNkfQxKWy8IbVKlEwL4
QApK8W8OV81TjlkEnJY8huLEChY1VUGhx5BWfJC6caAkxGflvroF5gBHLC0YQm8s
GhiYmxRG+35MchCrqJtVsEImfGnNnOL8Yyaj4JSoirFLmkXJ1sOqMFu78WteV/wl
iyDgVuK+jOnYan10ZS3x97qkZ7Wrb8BTjTH38+MSrWLrkWkslMbBgX8WXXvfPJpD
EQSDbLgpGbqRLM/6L5roPvVd4PLY/jrbUJwbt/bLr1AYcK9TaVDCSDz6B4Nva1b6
UTx8pQViJml/xIUGH4eTJCjuY14cSs6noHXA88n9Zv55tkRI61YlRMvqXbvC30cK
ecpY7H3f20yaS/1N+eRfVjnH+OcT///4mNKw5mPbn+//4nLxp/vJsoEmTzda9z6G
P3O/skmQEJnDob1Lsgi/z2Lst22K0yyLVIugaaingjeIP0xxbYYahO9gGp9vThK5
mfZnqwv4JICowZT78hXbtNobNAWf/1NZr16wAiI/SEoIy89yDhM3GduHdVpV1L7s
bQz42073p1O1xgbzBBEZUqDqplzyEOPEix+qWp89Wgxwic2gtELYzuSbBM8HQCds
2MuDT8KWRGJpxvsOKuJBWds0eXHW9xSA5PRwhfR4PJJZTZfNA1AplWKrWN3IMQ7N
qgwPs6D7JFvoMGL5dO9m5MBO3jVojpiaGx8EJjwTJV4hJx8DI5Te5MgOC0R2eol0
ri0k7SN+WZbKy838LToO9iXWFp6aMCg+38TW8c42j/Yo+3BLSzoXrmPnSlV6SV1b
ZzP43Lt2H/l36QpC8ndpURfTEajcegur9njPIJY+RtSXd6/mL8pCJMg/4zZR+8ud
LN6chSZwMq+2UhM+TbcgaIyKAZ3HlnetIHBoCd568ownT6DqfjGfHB77WGfD5Nv/
4EBaYcnhlo8+/o1wlbUSdgz7T52gnX1rJeGjXd0KX7w=
`protect END_PROTECTED
