`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKhJv+mWxIzGPqTDWa9/E+n4TmUgRqviMunq8QyqOhL+L5cSNbd+5IR8IcHwPeKk
1SaS2ihZn+8q0KF/D8Sw7HntfcMcb8eUHLlXMnfIGM1L81GEya6jeC9wGVpYnxx5
g5R0aVRnTaMv88C2rUsmN/fPpEg8hor6mNUDAYVM5jIhh3G5smmKEpWXrBuxY7wB
jG+ZlSL7JyTO7nOwE4lkEdObIVzxZMmUpu0BZBQ4ghF0PZtoeVvIVFTlNYwvqiiK
2+uMKYaDlyIqT9t2bIa9Om5NP5ShqxlpWNhp36BcksLMK6x/4oldU+vzXvzk4yzL
yKUNXbq2gFQ93HYgXhNjUsi22tYp4Cq0SV8k0T3eKJwQ0ph8CMV/6IN5v/6sLDW5
yGq/Mk6mFr22Zoj6abof62an8iQCebXn2XPcni1Lkdp2FChvm+2ML1Gx+FXWjyad
CaZAfPG1J/nd4morDZtzZAeqXDkBSVMAKwbxBuOzvn6uPHteyZaXKQnpL9A3MISB
QuQ1Hqqsvd3CR4SN+xhof0CD7nFXiSl5iaTDoT/Sk7ZRQMLXDl/bYHEWxj7L7Rzn
KgBFMQKvEBEwCQYC1k+3I2j4MbmFD4djK8lSMaeCs1zPTzHGkSXZvRRcjoVjMwGq
Uu/e+8hj1DHXNVC2jyy2m9gT6ivflvWGCrz43FVVlreq+7pA+Hx1ycTGWsl2QN+k
0+NAKqKtIVg1XmwhuBIZUnVnOXd+eBbxaVTdJPon9nHAri0/Ebsrp7X8QtrEb6pd
wCSbR/wv/UcM6gC4+xiG48MaTdjAZIMvbT+C98jTdF9cddhunxWaS+XtmjGgnUe9
s0X6XYI8Nqkfub/gRo0wJmKL57D3qGTS5q8K/tbeiTV34qynrEVEbhJXpakxANbE
Kcq4eQvezZ1rrLassC/yXj2R7Dip1e/uu/d+V5mNUBup9fzWhL8yYf3zGfrYn/CM
65riifvwMAZeIsrqUll6gwW+8WL2rcQJK3BOj1dHrCCOfFW/SbBA9i13zf6wnNRR
gk7+t/FwT/66hIO/QXznaWiLxpV7D3gsDtKjmC+cokmeXyuyoI05j82BnclS2Qgw
dP89Xf6fcYEPylWSAMBCzDST8eDMq5YofFxvGt099mgNAOJ+ws2OTmDXqb/I/42b
81kiMQbAGPfdo6NEsk5s5ynhpzuM5B/DX4wb9HMRfGaquS03BT8YsH2Kk/Nep3Yj
t/cCFL1vCvRuxFi2dB2kqwy14YytkE30f4txty7B4irdT/7keCz7XaTzArNKIeV/
IcVIHtBsKn/5TUArJ0I9SeEKvkGIsvB11VhiG1nbl8zmDJdT9OeIwgpx86C8z3N8
SMvmjG0tlNsyroWeG+oxhlb5uuAvK0F7eHp9B1O9pusnLGR94IRCC4zL/EBpHDFO
a03b36jh3E5IXBKJKemlXzStmU0ZJsAwMpSRKCPYKRqtmoDV9CJd3SpjozdiFrO6
Zy13L0WiKDN8i325e/7n4rWQkzwVeYWzi2JadG6wWOFmpmueEiN+15e+wHezZPGn
ex2TxcLdCvP0OE1r9WFdSRKxiBl/B0ovbEf5VRA8ZdCTvrdqUk8ppH7Tt8PVVLV6
yHRORlQMXMoeZI42Ynwyxe/0x35svx318mJnmdjADjgL4cHbiuFfFAz/nsaAdSiP
1/uJwHFRdxO4MrQnOYzbGAhs/epK2oFWOoqL5ssu4e2Kvo195n/ItNWsLLlUK+F/
931JuTYESKvA7Z0jN/gE3RqhTIih3+dujh7wn64HtUQfHd649lxIyXDXDv5Hj5vz
AwRDvVeEE28PB6yYm9ImVy4pyok7+AbRPyud5czqckoTYXnYSGzWU33BpX8rJXXF
u2j/sORi51nYVKn8Exuy9ZTgUGHaw4/ancUAaj7KEUMyEz/McNwRf91xwvopeW+U
aZdIdEuWuOk/H2QpnFmYI6s+g9LIolRqIqTBmBQOSIEdpVtNiERUb1OkxtY/CcW8
GonT9UhzrIcbjsL+RXf54RBCuFh0yAngl3Zlucn3H7xzyl3cXdMyS1Si39oicQ7F
SDToBvX8ETNfHPSyl85x9BjmiTGRJnBx0NxMLsiPmIlN4OprW1hXYCBiUTKWD3gB
5lNeY6YQ/uJeu9qQSgo6KhwAy+yvZIG5v6rj/axCQnXnz5aLky95b0gN3svhN8Br
WKsw+R6mfA7LzQLYlNCa7AksVaBqOiZp1syVjkAxlkCB1FVTybKnRBTHqJAA5w7c
s6TTyH53TQK9mDto4678VjdS39MZL4F1cjL+hQ5A0KYzzQmNK1s2qNUoJ1aUNRSf
xkJoRv/b5roJyhDN73exZkztBxMPHcEFlp0DSjLb37Q2ev0BXbBbya18bobYnD+R
3vuKODnqexLOp8CslGnHgnOZ7Wh8XKztztSjYMgmqtCdOJLx5jdJMmbUxcfxqYAZ
aL94WxFoGZWJNNHhnlWZJ0CfXth0NHKKYVE16VVOkacQjidwdVuBpq9cuQCx7T3x
sVaFkgNcENZCw+KiLZ+JQvFEZr0fiqwc2M12SbV/sMUL9cth1zyvfWZnC/Z/qZn+
dc+RYYbpr5GVyhLh+50CSlleMmRpo2lUCUufTkBhQ0hFxC1EHpPYZtkRqTcXqkw1
FUAAdCzhIu1J3THCtyB5PReKk60xHY2Ijn77CDZX88df93ZVjWPzwOx/IP82Y3Zw
9OX61TNwNufKkSMoWKLipoLwTizGIuhhKTlhyma1ZdXdQ4aLuU2/J/6Udds3giP6
rY9uaJF+hcPZL4FAsIvwem8Z2BBsbVd+xrJRYn+ulSfvhhMkxcfy8zj9Sg1GIszQ
pfmP+NorLkQEUdav7iDSm0Qeh7s387d/XXoIZtdhuew9Lkuf9n159cNnU2d57Ere
oAO/y2pfV2WyAGLDjMK6aF7C7q733M2MEhgr2HiAk4uc+jykq+PBZecW4QkrJilZ
a/kk2woWKj7WmrJZUMzqChE5c16m9JQj0uXEfbzgSFGCZJMGeDsKwNOmnAs67FVh
eLMMiZEQJLC2+1+qlHdHENFXEe4RjNK8lvwP/HI16iLDaGLrm99pCArmrRQ+6SKV
3/SpieS+oGDMqZl97crYWg==
`protect END_PROTECTED
