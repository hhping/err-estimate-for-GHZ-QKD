`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eo1a6zHCEYjYTXM+QhZquqJvVfa9MOjNjybkDc2EvnJeoNglYlSDnllWoCqbSv5p
MlTwsIS3QnQJ9d2HooTlKxcS8/P8NDED8UPaSYgqHD/WAHN99oZ2c4FUxUdESGyd
nTY/O0ZyTLG5FBsVBF5spFnzwEJoNVcesaiMfqXPzeIglMeD3zJ5ceM7hBJodvFy
QDsLixT1TqcMk3sbYcss6dKFe2bjsGxOPydxthSHfW/wMPsZMWR7RJgyvU4IrXZC
sY6Hv5m54AUJzzFQhKYDba7carmGZ9SjBejcPi4eiQLk3lVKqeVKTlW7gE/ba/Ts
1YuBBj3TA3Ge8Evp5QgI+sbRWYhDR+xja0DYxiPi2TqKjVawG3c8jyqdNSa9zMrz
xYVvnJKGwtEdLygUXL37VjoRB/GolxrRI8bLqvzAfU1St+sL7clyFuZb4xWkoGd/
J13w1nK7U+IEzZ7XJX1tbg2+qICyf2IL8uYBVEv4YwPp4ob+m4i1qvGXihLtFZaH
nDUBOmnlo6hqEBrEgA9DYRR9I5tP2Q1k6MV9yMXiYOYYr7P2DqArYMmmHEBc2u8R
LoEQpyVI9SRaTHnOROB/LQsqqjTDXWjKKDn1OVRMEyX1j7EX7LDzzwtkCTxHze56
rAYUM111Ks3YIfr7VbkOk6n6txkSl8jVxJD/XQaYPjREyYkWFaehZAAwSNdWhgJE
7z3NtRwr7aYMZ5fQeppUQwF/2T9FANBlP37d8fjXGyP9sGY7ehYa+rStUNVQNqAf
zgq2xx7GHx2HckhvLMOdaur0R7BNtdVB2rplPUHP1leUYaR3k+BRzvzkn/ZYvcjS
gahKlFBz0cvqJQbQ7E/kdGn7y0O4EppQ3sb33tAskaeuNWQXNPnmAzXhunkb10uv
cNk+0im9zZVllpYrhnUiaAwP9BXuq4swq4yTyIWkEnrgDn6B7KfMyS14w1RN6mJP
wUY3Eixj7YU04rS1ZHF3jeOoRH5F6yJfEpjR0HUV0p2wO4oo98FxrZp/YLIrAEbo
IqqDHrDg1iQUN9DpZIJaCH07xorc2XrmWQi3CmQGjicalaK81+8JKYpq8geO7DqW
vQjmzxN6WcwGPGWhWl0rGtQrFkOaMIqDilr9LtlsPJtq/n1n129wG3PVQA7liVuq
zzw1/u5eXa0jDuUYYtZGZZrZvOiJARtXa/Hw3jSdMHxI+H7lhpNYXISmHQm9jhv6
Cyppn3zD+WV8rsebo0ksjbgU2x2BmwY4V+1g1QJLaYzodk5km5CFSmDj0l79/SyU
6rPKL/gEyMyfD5MUIbSYKzM+JSUC3XZ+o/T2rNSIr72x4bn6dUDU40d1/N7Ne/o2
aNfwcjy4I+QHDciRJXrhaFksO19/jCwpqWWnyU4CeGv+neiY1aYfNn3/7qXFEZek
HqmPE11rLssG9Kx7q2b9xTsuBy1awfvpeW4lkpnfrTy+IcgeimAZQZY1yv1dlcf+
R/2QKrynLD0J7kovf9ii/M58uANadw1G6vOp2Af8ovsmvGEtuhrgH85Tq0UV4UYP
ESQKsIXXpEZD6Z0yd86OkMp1vD+YHTjesWS4agkQi5pUQrxaf31gGvj7taS3Pa3D
SqaYj/b5UjctXJo5wmKGbCqLhVuDDErsBIxK0pRtYEyixi0w/+upfSO3xqgdf2Ux
+NiLTE4dENHn2TphZs0hqGj85U2fRZxSIxGhggsUeW34EEFOtd79vEJt1ajnr9/2
430ZxTY6U37vaO7CEUAt7wuMBVMYhJWzP4d9759LiSfTjScimIsOoGkZL2JciJlp
t5xGMVPfV0OVDjX4gY3WOr+Ds+ULh97iEvGBdxwTjv/aokKBiNsS8DI0pPyz9ZTe
tnzrz36lfRmz3JImBOinBNoPUOk2NVd+DM29P7afX6KRaNkRMV8MaBOElZyJ/AmU
P4ZoMQltbl0/hblDb1d+uWiQ8blOIbY2mManBAic8VQ=
`protect END_PROTECTED
