`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDUeyy1bL4tV/bk0deGXmyBJr1RejNj01sDmG0UWxceHrZIrDSmWmQbEQ9XJ+MFB
gBkuSk2bKFINrPNofyyz0sMltmNRn7YVjxKlz6d4OsyBGyrXab4yHbuGIrm/MD9K
zuF2sV4urS2vON5zLhwjYi+dyl8B+qe5E/sbJPKPQyKSsimCGhHqWx73kzpq/08U
YAuh/EM3/DFgjQ2yNLOmyU2CpOY5g4TsvDY0Ub90KHlfcyJV4UyMGLEAppBprZyj
TQiJ8i4O1yWKAy+hU48QbYyqUTSQfMHhCXEYOaYLC47YUKgv989kGcAvWoh7muxo
UT9E1lgw+VHojifHa9ccfkyLwoMa5Js8p6XaWELsNb39DIeci91gZqwdvMtVXFg4
09f1r8FsFr4pJmKopRob/o4Ng4fwNVMzsvjnUr+uXwBny+ftF8MIt+DChSUEvSZ0
RZJZWbsb/YkoiYD9uEhFDxgnd+qsqFK2PS/Z+sru0ozR3NltG16HixPrmpDUTgEz
5By4vHX6espqC4jVUERaVT+sfzh5tyyXCt/rYCYWEsiYi56rNC2lBve+DHPqBJG/
oVExmENypcWIRMS90xb7O/n0PRbhrfJJfSbCwRP8Os7TqVa9J3368+cVBPReOpJk
uomxRSiUUCT/aL3OpY1LgS2tt3vka93jEIlVNZbsA9bL7Hb91aN5kz8r5D32KE/j
SpMEGZrRi/CXyQxnEYdIR89qH5R0+wsYVNpIh0FPWe42ETU/6ZYQaWmqSdOZ2w4H
PZzJarTnHvu+F8x48zLox1kuWNhH2kZLfGMNGI9HY7CaRTOp15u03TA8CCn39YbN
D4yw97qYVA1+LNaEDNmcsDaQhxHL0Zs0svRdslvE1tDVux7cFgt4nqcgM2xuIb/c
C8P+D81ph/PxlzjqBXoMzrQOIpuRU0qGUB8oTVWJ8Z96TmMB4EmCSLdlViiEA8V8
5aJSDnoj2Kh4UJtk3YYuEMXBJS2YPTIuM0UQEL6bgEsul4nTdDjPskAOxUv/w+Dw
IKD0F2tKJRmhsLOnM3mDpIiCF1sHvo83M4QSQrn8t4aEYHwyWWxYN+u1hmdasJxj
PH7URAomRf1lcfFowH1Sag==
`protect END_PROTECTED
