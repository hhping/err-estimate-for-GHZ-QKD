`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mm4z0i8jH5xkzUMSu8BM33PVPGK0HHFc76dTFtf6CaLVjfFARFemL2Lh392fs3tC
UZvczyc8YjBkxykqsytP/UHgEbQz/RpUVkRGyuBQApCzKFtB2JrLcf57Axx8ImET
qvUbEDmlEvXz6vSXdUplDLFDYWAxUsgwe/wWqx1JmpQXwUSa4ppt+ADgoq+EEY0u
kxCZ+b1Sdc/izn8o2e9gTBOusqt3c2gcasJ4igB5PoJqEAjDg0PJPhunclqAsJsV
Qx267F0QzQ6AOLMAhJEcjEC3nb65NcZ6rUi29MMAAKA=
`protect END_PROTECTED
