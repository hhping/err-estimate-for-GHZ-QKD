`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3oMEhjqwsasQGov9m23SPwNeMCrFJ/qP3vDjBxgMWkaZZhkeCqlIqcDcbBG0+/4h
2rb48mqM9THGix9j5zrAX6K39IJg7P8HA5suwu12R7Km4YoN5c1rz2CEf4jZz8gI
4fNC+r1n8OdJKVvvaMZUhREFEI6gKSqE56/bkiRL9DkEoVXOBdYIf5Lrwppq8u3o
hTDZigIGOs5O0QwFGXRVhGNEu2WhGhbXROr//YPcUzvfPqIqb8/US2AwAiS9dvkT
v2dyTFbyR+ifObbFNeYzc14+Uq8h9gq/6on6GPFcIkHworU8wcw849fRHQG7VcW2
NMnTYqgLx1oN2BmEJIoDnUluSLSLm3qa3nloAowrQ+vSLrJvOUCILmWMZ2pnMza4
A0o/EnFs+SKtiEUqUEvr75DXfRIXvEfrplbB9P/vaNbGcBDmDALWD22jNrF6M8z9
atEEfYW01apnLCe+S2dqYE//m/ONU6HnHeFIbaLphxl03CEf92OFaSe0pgtJpZzB
1Ced9MEBDKYzmigfCrWw0raVcYMnnraCf84T1TOPgcwd5rKXkplhRmmVybym/4I0
8qvYrANS59RrXniIjV7H9Qpf0JxPcYJEK+GJWPUGyc0+DAur8+2/WljRq160A84G
f8jgFg7SJUXyPWxdAJXF4hPPlgGBQQmcXuhsBTgXZL3ZSkEGDMN1z2HvjXeDjw5O
2eydqDF4rexyElJeISml6Rs50Z8XOkFEjxg7ESFxUf309bcLkIcCpXPhj7DBPcAc
JKDRO4mft9NHnZTICav7w7UcgpbcdcqMUIx0VtMFXh2vDoinVBs2g8QnJ7q1C83U
g+IESAdWLYyz3EaoNdAKNsPSr66kBUEYEmQ0A1aKuZwpnKK6pOa1R1lEWyAsufVQ
9XaMwK/CR3B610NBTJM9Z5uNdWWW4HkozMG3pA7T569Bxzxp+BhyXXM1FoOMZG6H
EV0oJcEmJvb97TOBW9wLe/PmBPx7pf20jMai1vJv7YnE6UCS6A2qbbw0l6lgJVFV
0HzGbix+X+l2pQmKLagB7IfcG/SpWRTY78sW67eaZ39FyXoVccUJJ8DnvDvANe8S
RLN01qUtCQAbaVge6Oeuq/8QM+ZpflHybVoy4wbjPd3f4u9V7JthdJM8O7T64UAj
dJc79Xpz7CPw/FOzEwfuXvc4w53doXdf3UC0MMxiax9vBHVYAzQDrRaPMw0mUlfT
MFNhVCDGALgA+SwwkeF2RhDXX+kpTmpYfog+vgVEUvMt/I9cwZjo+4PYU00tONQW
2LIZoWRJc/ZEciZBnc8z6BM6XAlnZcU/qpSwoHXeNi8KT4xmxqiNEB7cN58mX+hO
kXQtx1vKC/43hJK9D4fJ5Y16JdyF2mozx1t6edo0xjWsr0WwpqiWpZ1u4uTtWTkT
W9N2hXjuoIws1i238zCNpWRFVezaipm/3R29GEckGg3ltnU2OBFD1rWizLWlELCG
yryGnMYSK3yEWlwOsdxcTI0sBEytYmqu569fr6y/d7cPNtS9E3CBbJy1We4w3haG
3hrrgpibMTK6Oa4HDZx81qW7zqV/BL2kK6rKxWQ8mnx5oqiNl7649jqtMUgGxXjk
T3tbeVhMzCaED9kZd5WsbcK8UleiJz7CtPzc/geOok96PC8S8FoQzfjSTFHgYZoQ
PWjmQnlci8j5wrgM1kUScmykF0eVs+EbsHpPxLny6Peotlj5IGJiyH8IdZhdpb3P
4cPr3oTboTepA59DVeLS+B4k98JI43+0z7pVK2tUAOdKKDbGKMEvFZofEj/8oFeh
3SPTAliUfQfk8u4XlGP16uLjVyxw/uVcDgJeGJZN52B3d6k32tmlS2KiegItJvFh
sY8BgcXpRiZtVYpjh6uu0ANrd1RR4vbQiTEm2HctUD+deEULY5cxPEWetgdJ/hTv
FCKfMv3zkoJdTexjav6zqXVLanC+GknSVECJiYRPPQDzFHOqyrOBdQV0Oc0vep/G
KFdJT6xV498OWYDfWvIeP6dHzWGxgcccxpZbeaiBKEeF2v6JNu6dGv/Zs2VrREqw
rCh+XML1yZU8qssGU/a5ZMwzgMqPCy1wES/RAhIh4ZC2jmQJMKlJNFBfp4u14qEb
QXHn5TH28QyP5+9iGDZ3Wu8sixqegrXDgmJwNqInIz0BuAaucQeUZwK5guoyOz1R
OqpNqIh8+I/7rac+N4ythYepFFvrr+U6D7hPqxrm6dXsEWmVf2cXDzEDmK6E8frw
kR3hEj2R5g4Gm86ulp9iQKaVtr0vw54SdFOqnHDCoH93pOq88+BnF/uQ7PVF95qt
OUH2eh0GPnOhW51YhkUvWriPPunXNgqhsd+yUNBFduUzYpcIl1pkRAJxwmoS9AY2
eawyRVTaMZSppN3la/NRf6Q2ChDiOMSSFqMTPugiTxhWUQF+Xsp4zAY/G0X9/qjf
jQb9HX/ZdJpqQy2uN8KRsz1JG7Q5bAqZvPdtgAykmDQN97fmfA9KmUX78oH9cmVH
SKe59NyPK6HcViQjX9yxOzTEnEZhLQEumdY7nNlqk9VXxhtMP+MPWXo/sluGl7BP
vYLXxoxtUrEHohn7+DytFzSxs3v3Wc8geqDua987rcYzo17bVr7FtPI5cFlZz2b7
qMYWIH/iipqFllBzg/LYnG3qyuFVtSbB7C0DwzQ1zxFxc2TOCu3Q51Rh5WSRYDJt
Mz8XXalHIhJWBjr89M2IGMW+TSB1lJmH4EuaWsiV5PFvmX8Lt5RswJzMcAkE3WVT
InDmyw5L37/tKkbp1mow3evdzBoGpC/oAROGCGgJX8is/7MKBlwLbE3JDFpF1hMS
Ed+xF8Dl6fWpMv9E0VQrCwTsB+cPqUQjmle5ufBhgeBEW4ppkZbdYO5ah4CNnyG0
2pyEzOBg8JccESwycvc9rq7xbMvq+9Tdyjj7f9bYdja+azY3/szkUihxbNrt6ZaR
3+Lf7FnocSWCNr7caR9gbaFwwQpB6uUcwDsrgUq85yae/t78AOhG+knbJqUdb71M
SXs2CBYVK2lhL6w35dkrqSifhPywmoUoH33iCvHmdEfLE6oKVYDvIkXnKCJu32aN
vcX3UhNWX6GR0STqQBOYDw9J/PDgTr8ycZRWDzMatDBXYAYlgKQ2eajqScjqmia0
Jq/Q1J4DLXFsyoGIo5EsMs8t+t2IEhJoduZgzcfZFTcXQMpviecQX0Ss4KSeBi9D
zzEmdrVKq9Mdnpgb/MiBiQxyO/eXZE4GqwV4Ga/6JUYvDWyEVzDP2cJrSkuDe+ST
nH3kwXAx4nXg8CPnae2/GFAGeO2FXS8hZRq67HnyjplZyeKcopMVRxQiDAj3Crf7
ut0muFtg80Ed96ywVV+89L9b+d6mWNz3FNBr2oMUTV5AO4jFNstT3eIGzzv8O0k1
+43YrG+70uYPyZ22oD+Kyhty9s6sFb1TpfDB8dpi957F9n1tCBiY7gKc3uxbfbDU
yaPGdRmn72W1eE4fH3YWMvN70bqkFn2DH5nr7/RabGuifE0xSHK6tcUyVTsjxmgj
auT9JlXNQpvxsb8o6HIafNMNmw6I+lJSJQW/IZXEYZLxtznXFrq4/heFt1SJwEeM
GPTwZbv2h2AWe/p30HtNFNgxYwz0soKxGHj8txu+KixOMB6JfGOaFXF3qz3QQm+L
5ng4m3WGPZep6bHoLqAczwQhqZrh0CzjQL9J/sjKXhpgUR0DJ/nZhwgkpfiE3yD5
gILNfAPV8ycp2/KpfRYVKIK0epNrZpvr7+9+E550Q3X8ELC2zPtuRYoURUF6eS38
WZL6yTVWPy2dOQDEVsSkWo//c+oJfF5Y3hmOPl3slPI2DjRDSRfuhyvXIDET7z1e
P/C4HMDz0q26s1jQnNEpN9/BlJi4JyEGSjsh90B89IlJy6hOpaXCSIfLhE3YmFvc
se9bhmo76Z9PqIru7Cs0ARmXr3ArIAXe8B/PBoDRHxY=
`protect END_PROTECTED
