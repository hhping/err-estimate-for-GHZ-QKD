`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uemyjvNoeotJX4bX5oYljQTgdOnFMCR6V4W8YMCHJoUXuvdZ6hfHwYeN0Y8A0ye6
FhWh2qR9P5XUupMFqCbG9Mz1+G1V/hlT5qgGO25gyMYZq9+1LThyxnJq3EjD+RYH
wLq8dfmPdwemIocS+QuobK8RBGDhQgJ4Yy/vzcI+g8vTgObrc32Dhj9FhF/xJLTx
rOqo1NguARv5AQw6PKMJ8sxTrcl3L8T/eaK/2Loe+xwvi5O11GWjGXXxVOSil/qs
7e03/PswG852NK/EJHM5mIKE8qnapoWU+pc4r4I8JTsTclaVbIw1QJNCv2X/63Os
TxLVTJlfcCw1DNlSishdjBA3ZZXSfV/Ver3oJTQgdbPDhNKj/Ejsp8W/kPRk/ewL
BBxhh3+hwpLpVf00ZdEylxA2VyBBBuK7BJG+PIKt+HWetASJLO8YyC12+KaV3O9U
Teb+IEq6H+wPMnjT0X2nVcoR/23/uhTBQgr7Pv4wU+K+HZURPxqm7xNM5e9nLbzK
+WhpOVZtfN41Bg1Ddnh5zpBg5Tq4alr30KPqmcavnwEADiTO3J9XOdNbo5cDjbA7
70i20UjIxTTPh55ftmGme1LQfe7BriT6KCSvNGHBFCu+n1ipZu2yRThyvGLqQO7u
aSsI1nO8NQlzDjvN4zBRF3osW9l9BlibzFIsZa0DMeC5IMGjrJ0QxRKx5fCNQrw9
`protect END_PROTECTED
