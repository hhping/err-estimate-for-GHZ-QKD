`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXLb6zf1JW2VCBBnUCUwISAXlGKv4LGiMynGynlE9bVs9ucbZG/IzbJCrTCvOQ61
ALzQuxtvmDfVmCwk+pnllmSJDuE4tB2nAQFt9vmIT2aZMXrEgBuRHsUaV2xqROyY
SwQC+JEcr73cafAO5Qc1nhBBmVw+BH9m16DGoireXhlgxtLk5pmNC377QHOpmE1K
3XrD1CMkJp9fcqBlZ8f9/gDrlg4h+PamKSk5Q+8nVbcqSGLjI2HJRS0Yd71mfh45
NhBLRaoCuTdvulep/s4r2S7egY9dpwrR4g3UZ0bDhX/27Iw6xs0pQ4+zb9QIgEf+
8sZo6GkKiXyMJDq/XQ/LMJAjn/d9rnft4sxfOesoAdZ5VKlfiOlJYOYeIs1mo6MA
u0UG6UG5bAJ+8GSFV/bBDqUa7r2Kno+4jL1eY1ve0Rcqg39eudf53q++GGjlNoAA
uahB94DvHZzcT3bwTGBEMLQXjnWp6w8MUV95I5aB/NqsINd6unWkrmjqt1frH986
HiG57hzfxzWXUipN12/MWaRfOIxImWSGQdehqsKPjFhOlGCMuZ9qgH+OVCxF/Tl7
0yw2gm32SIchFTfwKGnXZEByTgG61Lyuj80uLLEjYjIUVU8mQlRpWKwowsYfhjsG
G5t7wlnrmXBtBlTY3nHphIZb1lSMNtrdtX+TU0tsTrmtalXqYMsXzbF9FM3xmuIV
xAF87xHB6U+N0jDupQJcksrYEjBLKhYXzwNd8XBaXaNMt2sKrJcGv+wnJfMdOLRa
cNF7G1GBfWZ7K5RDk5NtDwRq8ZrCU+ipl0oQ+veFGoOJ0DMdxRR7mtQ/n8jAhhrB
ajRCtfTJJk6t1QmHDy53l5FpDyAZMyBop58bruF0Ft7KivpD+YxN8J0AfMFZMmyO
8FIDTTye3J/jImyls8uBtMEHsfjOQsiJwtdeNacBTZ0Mvz6fpcQDYWgZw9tNg46C
dCiI1RLbzV6YlHpyCu13cdHG2x64T79BzDY4cd9OVMU1cYjh8IOL2Jkl8iFkIJ/P
V94hTYQcCHxcW9dJg+4dMXgjjz8AFV4KMwFs5yjxpxObHVLoqTe28ry4Gk6Kc+61
5hexEuBbFZeQ0ltXIfK9p1LaweJ2brY/H/rP2u5YqrrfDZsYBz/s6n5glbNoFHUc
PO0udxreJJMVef3eOcU+fcXaZo072iNSsy0Sxy/bPN+LwUjw5BDpnBF6ImjQtEk9
eYs2suGKj+mHsxEg21WKbCQxN3Cwex38dIYYg897uv7CGXGOIYKbY9Snf1tK3Xr8
BG5wGzhnnd3TZhlNTgAByip/bYgGnzVhsJjNT3HGOLaIAEtyvS9xAI4y5+Fi7dYq
iIhlCJsgVtBw0ux4FeuFZfkN/1MvQvw0nUFkVON2dDPuk2NLfp5cUPZgqpD0GFyf
bgVkCISzZWLfCCTLstP2/t6mXmmJrP89aS/NOSOHMWgJVUis7oz5LddRohl6hypr
o6sLhx2ZKEvfjrjnFOd0P6F7nnmtStwLFOUPZ+UHUIXjowMQwGQHsw8gvJaWG0xO
svzE34EdLMVIxURVoaizslKXUzEWzv7rByEXTysvXyZSjCoJRHhgGrSjnTsXWEX0
GAJcVh29yisx+Q0iu31FthrQbs/df5aT9s/gj6UlkXmEV+UeOebbRhsavrV3kRxW
Dv/dHOnb+DvLH8nG3kv7QUiyFNLyvrrUUREVrUUgRBDeRxMgIwSOCiVKAFPaht9+
CJep0cFlRuUwNsJnoOKOhHSIuicad/Dw+jGnMeB3tFoDAAEpUl52CpyjS1lKL9KN
YgPqxDbjKJQznZ2R8Opog016U8kqQ+bcbXAssSEfDVT5iNpYCwR28voGbqgHbm+3
5y9wXQjr3Vpq6ieMktwd/AU+3sGb1CFxtdRTgnT8tIIXFvPn/B0LfLxVL2+1b1AV
6Vpz1VEW5mg43fz4PyppSHGu3PbVmgqR+vyTeb5H8cKvFMxiCIStcJBjxWnUjEd2
Hc8SymhCjG+SfP3CkotFQVFIWb5j7Ig1Mq6ke9KykJXIytibW+4yXfziSJGUTmFU
DslaqXScBd0gjZOBcRd2mXDnen7kCMUySfz1W560HPZclD+9ZTeRW4iObZZhhnSm
Gj6uXdF1Oy2MEbZw/6glDTiNJx6QqA9Zrw/en1gxiuQGOvpqfgTtJe5dKBeCzos6
5ZkE1HZzQ+QhtyFiQD9ahL99lVq4NvATAI/d9/5S3jfBDQ5/gHvS7YHvuvNrXI/9
FrIFWfIgUdXFPg8g2i1krZI7jtoLNF/1MJ8+VaxWpWlALEUmETbaZ7+gM6oRWA4c
J6c29TRh+E1ZVH17FDaxv0uN+0DadkV9xZdY10QbvfqimUwM1SAWQm2ylatjwaZd
/U+daPE8Tz1O53nYJF8kUGgyt6SGZDt/yrkKBYTHr02za4MvQJsWQtDziHMNrq4G
ROvGApj/3wORzKhEraw0kBlgsOznXkZCPwmVB4OCqRYk/ALEUOWL8LEP360Og75p
Zdyq8gf/5Es95DaMiZ4VY1mN1VE1KwXLLziBfalGQ59rlL27PtGGVeIcwl4JdRHJ
xfb/sZlAxTURJ7pm51gS1E2L2XOgiAMnSh1RCFAUBg6mIu/2s4AtqkLM41fGZihP
35/BSdqNUoldMVrc82HZ1T0xAVx+8EePugX8Sip/OrunraQtVrmSTm5nYIMmbPs5
OIROI1q6d5bic+Z4vqTde8KLEVAsyOfEo3SbacC2+G96iYCALipGf/mF5pGf9SPS
LwMXhO3OgHLmYmQV9qBUF2rb8LxbmQHHg7RFsHIWXOluduQtOk+PcPjntP6TvwcG
s7ukZdAPBLw+TKR+uxpK1F+TBj19644k3f6EHW0rtzkxeYao853Yf8B2NT+IJIlL
MMfWaCmAgqUEvb38b0/eMu9Kcy4q3Dj78Y8SVz0wJRKynqMF68T49L32emap3uLU
jjKKOD3OvLbeAJW2LXDOtipWIpBaYii6knSagRFUMZ/JTEMPIyFNE0bYOuRX7Y+c
da0v18/CXA7idv7Q/0QrPf/Vhc2/IBxs2yWQWADsQf4cxv88BQ6mroYvBsEo1KLZ
Eq0AJr6Yy863Q+YV6P1R1Khb0U77f1OGb3MEcDPsDWh4AZN12UCaWOL5FebgyfRj
xRbm3gckwXelJh7hj/gIELBmLm8/cTJ0pLw6sWxNHol9wCrRsI196eM2mrHrGrg2
R5uxW4iFYks2Zxb58FLlmke2zUaWwouKvQi3fBlMX21nLlU8tVl8NpKlL+GL+Iw7
tAkF8sj4cdWBVndoTs660wnQF21dJwE7dOrNHaUqeqrArR1FVZNmCnMtWyWtGl3X
CWicNGRapWBOome5RTjKt3PXffiR0Unuq2LxW3xIEndcetDWR1KZ6sbQ0aocdh1O
iEXt2PPsqqBnJGOEJZRnPmxuo3jCivzk3sKxL44B1RoKmYpqtmUSjcqNGh1VJ6bN
94+sPgGyS8CEkna3QjTkK8PL+lPQAvOXUSLvS9qFSnt0PQy0ZTv1UqJJDcM0LF84
dTZU6XuGNIh0B5ucKWYnsiAfB5bni8T2wyG2+/v+J7WLFHYp1v2jwjlSEACVnmsb
jOjn1dWu4vieHp3MxGkmXztdpzj2Dcg2vVv+yl9rCypMqJw4dkpmCKAnt/7tIddj
34Pff5nhzw4bkiopzCHgykNudRjaP2T51z8fOeQGKx8ZOI6Z2yrcgvnmCJ9iBkP9
0zVVtEIfDsZBWXiw5vxeXXgzL6A12NIF+mrpDYFxuUodwe61wqEbNZMVBtztvMQT
StlNt1NE5WRrii5uzWv8Fpzd35VbcRbsQL1OmRASCLkfcN1Hchg2TzADDFTt6Ix+
MGAw1HZKEwrIVHs7wFc0TwDvBvCBCWe04RKYf9azRyoKTWsaCBOVBqir4oJIMSmP
JULUlbSNLLxDHjoGlvUWEiCB15misBvz9JEMfZRjQU0irfqKbko9+WirueDopbUU
4PvhwasLZDeFTaQVSWVhMsz+VGWKgyQjOe0g4+PM7x4vwsSYvLw5kx2YWTRR0+nS
lF7Bo9YFrJqMtCmaCHJYb544aKgkh0/TqidmK+NAgd4vA4GkZ3PRAo2xm21H50mY
/dnKdo2UCYPZ2uoKlzChgV6BiubNYXthBZAGs4ErvD/Dcykkxbmrs8SLo08uv10T
BQXINB0/dMwJRrllPuaiHrog9QC9/Nb85p2IBON54iX3ZyCSHJw2vlMOMkyFxJD0
3+2Sp9ojtSISnY5ma0U7EY1O7Xeosxc5pe6TNc48J8AiA+q+vQXx5Lmk+O7C69yq
wwMAD7W0QfrWHb1hJVm61mkAZ1IpMB0TX4x7g2tWiIYSsmQWt5SYQiLTyAtNrZzJ
c/6+7QiHxXZtWW36rj2DYjDJ7Kn0hP/yqiJYE/FyESA=
`protect END_PROTECTED
