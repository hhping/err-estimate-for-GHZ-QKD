`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMw0+ceA9qglGA2cTzJDOs1jnLqj1RVhl8ZHdgVa2GmtL3sw6/v8E2sXO/AVirbT
4gHqUYJJlDCPq/aYLgU0YSS8s5VDmxLmTT9TWjQIgf8HaH2UhhQacmgbP6cOYS5o
eGjV/C8sdugrxqlQDLdoLnMKgFwFwJdTOBs4dnxDO5zrtUDkhboaG4XSCFpNEM1m
tuVWYWyUeKQ75mDDUBrvhQX8N1hdadkVRqc+fV27B4Lnz97fQ2Ao1xpiqDAoYpH0
yy+fgx3M4w3pzUEGJI7i59mmSKGXcb0vXNjeJXAbi7WQQBEfECt062dohpgN8uCk
/7nFmh4WshTUX6WQF3zE4S8/WqDd0Lhn77/zSsc2WLSimsjfTcz8tpYuKytUzXh6
ziEbCgULEoNW7Nk4yVviwxN7U8nvQwlhQPV68hYX5KMamdAH51rRox+j/imEckGv
YiBGO0tNjwT9prXzpeAta5PxZAKmALluyzNxHWEH0IepU++oDsXVn15Z0O2lOg7i
1QQ4WrYM+TUQsXz4OnmcXYrh4zfhmoqtEIwJBf+2iNjGvK3AvKpGRCUO2IYBNwEX
CoAlmraom2xOxMPw1MMNcaE2AwQq49STIy2n1MRbG6ST1Zapmyj96V2lbb1qV0Ld
`protect END_PROTECTED
