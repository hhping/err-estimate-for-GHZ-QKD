`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFaAffvHp+sgPBSSLLRHk+SHlUiQ4m447HoLswqjnAGYt/lJO7KFdmm/LUuoQk0H
jsj/dRdNEKhMT06/NpRlmjikXGSajK9ARzJNNhARK4xrIByFuXJIESJyw2OAHOoF
5lW0G2HCdp68zfwHZ9acZErocPg/w9kUl/Bs/4ZdlTP/A2u0Yn29QJSjsL9mw2kh
OgOadBbAPJNZX9uh68ivCGLayib6R761jzxTzNCmAOaCeovzhPyJisRIF0nigrLi
vr7ZuxOg55uNE0TysLc1WgD3ni55tn5hjOgIjEyWiQLcqbhUNA1Mw6ogpNTPAna0
PT6eUZ69JdpRKXUNEpK1cxn8QEikUr4g7f18ycxYPMp1vPb+1iipM0NBg5hQ9ZTn
HitHg3M+6eWYsBK7b8db8s+6KcdcLXSoU7O3WtTh6isRStDAWKZhnmbhURFHg3D7
dPryuSdzTRfOBt4mqbWSeC55OB6ihjcwI7Ls8vVOneAhnA9BdHn3B11AtpDxOEH4
firQC5FLrMFgCsZKxW/EIE4sJs7iByKjOsxPombnC9gZ0YLhnxZq2Ll3lc3PeQ2t
Snup3eALt9lyjMJ7kYRwUPSQuCXZli/G8uPKYXta5LwW8W7fASx62Om6cqktyg2R
Dy3JsKwbcxn9dZ/jMqLrsmisSB1YOumDP74cqPfdsbO05UkvPs3YxyqQM8uM+g4n
sGifT6zafMd56PYTDvNBevES1TNLmCDqVQLlVpzDDblRUs5jpgePjksZZw3ysDsw
E9Y5I7lLwxuJlh7Qyvh9gyZhoUhugOrkIdVquQmPrqEaPl4eLhs76kRPSZj0kCil
oXyqZFEalQGIC/9CCIJSx55A5S3tplJkuWQoFnxvqkJuNQaHjt+VW/JN7kGOu38V
9a+RT9RjhAIAqbbkaafPUw37O6TxV4IOy4cEfy0WZi9TxVOp7XH01FVtvU4+RoDO
WvpyXdFuWyhRvX7W3ayBd2hJfgIW4kuzAGJpZdme7KFWsjFfEn4rHwJ+KnW6R8Ki
HKWYU4wRKYmvHCLdnc1PXzVQFlZbia6P6MGV1v4qbqgMGO2K0i05W5trOAHVWKpt
BEOEG8984dbNdaEkTGfcHee1ZefN9PLOHXcKhpvsMUB51095WBFP6BLgVajYdv5W
qjK2v8Vl5Qzx4lZsiANj71SHjLVdNHITvrYjjjAwnivIXVAtYqbGac7B7whtRp3d
7KX4s0W4V94v3tnYvf5E71nQQOfFOY1VZi7qjioHHJTxiksrrcVVr9I/FEPTR3I4
1nJkwJRUJ/tjVZOqZmQF6d//BkRFCk9EdYY8YABZ4jVrSS/cSy0npiQFmk+d7Zy3
TdPBvUMK1xZrW6g/uZYo7trSjFTB9d7yAfGF7Lql9TtSY4AESJ4n+F+MESkCtqhJ
4bH2Q+dvOhGkxffzMp0YY/XxUmw8tfxMXwrRhKnz60bqhHkfVH0P7UWwYD2vm1rC
Xs9FOBsKigYSyVmqudZU+FeH2HjELA5feWSvQtw8kHqE71jDIlxh868DR2v55zjr
6/luLh2M28hQ/2Kull6XHRpsphlp/wih5q0/2E85tQyaHnJLRDFHyjB6cU7GbsbI
uNhpLB/12Vdm9qoKw1tYyDvAHyEgJTrB/98WATr0Geg/I+IN5jlKW+bdwF/MS/pH
WNvNCEsIPoxqRP6yd2++vLRtMnz6v8AsDIlE45kYNkB0rW8O9dVPlYsZM4zGn6Gr
G/+tBICl6Z0goKTMVsbR3rXM3YUMOW7FdqOFUYEzaPx8DOXYOc4fmosjEUxnhqLf
HS+5OUrm7qER/6Vg106Qa5t2hvEiAbAYbwmYhYeUWmvUH3Z+TggRJray9aDrO44f
XqUqpPRwsknXeazd+RQpzSD2PcO9rSeRrTfrKpKZPE9C100GULRh4Z50fQUOoVcL
2gnboaWLdZyvINGcq0ZHBdO22gCdJAVctJlOzMjbtSzYtOEPUrPvNcaNFKF/OY7g
9ey7mPQFi20SJ4gu4cB/X903PkODIdmLOm9K2W4rUE4eaN+DeULcpfcaQ3iLDA0H
UxY3tOt05ofHvM0T5+1oxrwv0XAXBfpBJVAAe4LMZq0LQU2D8QM/pac2QXfdPRff
yY3exlxAtRcW7aSlYzZZWHLeMHYYyPFJO8TCdl0Vu+Y=
`protect END_PROTECTED
