`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byCVg5Odz4CSPjsL9/AAPUAVqvMQzgfBwYxRW0eLUHrVoCQaVzzw1TUoMZ/een64
rN16HYCKyusci2Vt7s43E0NxkB6m03VViiqgoNYBio02q3QBUhnqfhyVIjzXVqHm
/rpLRRwx6LgRdDNQrlkDiPyc1wuzG9snhrrsZljCHQr83xiopvaw77dC9tSPLYBN
SYnRnZ3AFM0pGOt3KELzsSGaYA+RQU1GLmnmeV5X3H7T5lvLbFFAv7CZjm5EJwTj
Uus9TZdGMCaOZsCuyNa0mmZrs5ml9LlgMvXDionP1Fe3UQ6yJ+sucXHOKLqsr1+g
rJdFdV9xtTBt/FmUNFypMA30VlSR2n/bk4DUlDVZ/l4hF3YBIwRXDwzMctX6/+rV
IpZtOoaZ1FTTfRmXqtDXZEA9lfUN+25KXW/DS9wr2SBry0U9+E+XASwu7xU7a0oR
vrqgLw/Vlc4lxWBm1T2WWlXZHdIBv4lz7Sa2jiKUMUFAaeK+srGBBfu7ZZksnraV
RVHToO0TRspjeT6zBgCVCU/tsp/oRNX0gCHjdc8PHSFyDX/TPVIFZ4vzBbJsXpf4
8fdxAU+Lb89VpWE84Vsg2ZbQpuUaoRdrqAOUvONeSTj4Mtk3I8nXHBpMd/5UyuEO
qTKI+z2HghZrh5AbO5jbt8h68oGAqjSo0J2H77ycHWM=
`protect END_PROTECTED
