`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzLxmtWUYFGU94AJWecT6X7I2DYHLn+ARyYr6viecqQDJ3p0lrZODbcS52JpEw2S
KyJ0W525a8twXi0D8hKzyBS/jJ8424zsHLMIO84MZp77quDcNaVYIFfTr8YCRn6m
iwCRtfgiV14DVOc8W7AaERUUJCYt+6z2PwzUOpVRe1kKAPpnmct48MQcbR/OQDvT
iQHA+XdFx2piorU+eI91E+7BR2NxwFjbGtnYAUb4Yhqh5B9crLw1Ktgk0xnnaXwC
yS+ovT0WMb9Chc18zrUq5zOzuvKr0w8rEcV3S+ykzgJouc8MPFuIbQsy09SHuu7M
NwpSMIBVPe1tBGN6UPsHy2442pAqQcda3Vk/f83SH0ponHs82cc1Kq85AyMnf1S/
Ob/rD6VG+juap8YdJZyFf+pKPsCddpyxe13xuO7Xg5y6eS20cf3D/65ui77eLS1Z
O0tuTcT33+iTBjpr4eHNf7lYczJksIJdlxfHz24FjZxMCib4XCjmGH50Uqi2dLc4
GzaH7++2B9BHBTeeBJMyQF0R5YChk8ptv2s7egQxSlznkw6QtzkJo0ISu3uSrMvI
X8AtwXazRBF6o2yq84UC3d1YKgWr1NNeXi7hOzZeVKY+aLA94eVrxW8SjSW7A8p9
FmFXQuaAbbUzM8NezOwFkSjmF4BEdFqaMtk6gw3fd/+jXLwLu6TagM38lPl1Rqi8
8TNYrtQ/DylkLvNBXx75utUkoCPOoOfeL6zTTLDDWqVupRZUgFH/LrivYYO5kv36
pxW57yN9pniqty2JLYDXY2bZhUxT8xXCVAKBYIwCrw2zl+lZY68rHjAnIEQLXkdv
njEnCV/J5wpiyIY6hcnThbVTo+f4VpR/69+yJ3U7cxQmuBPeLvestH9Q+UOr/RZK
`protect END_PROTECTED
