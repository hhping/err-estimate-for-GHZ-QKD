`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
la6FGZkUTIB+L59TWN21o+9MnMcs7btgAhjgaRYHkIi7Q9drMJ5bpyo1SVrXJWCa
EsvwrrMSUgo/i/m5FwOY0BfOLAmFY+0KNz6Vs+hoQnPvF3FbYLKIsqkbK+OIGlyd
9vdYFVtG+sAYCoRNuM3sF2haPt4NcAXbsdNPjr0tcFv7eUIXDtihzSEuUeADf36G
5RyRFuRRi3SWLMNjGVV8+9uwFLo0y6NCLCPfxqxIgKHvmeTe2MggLokYGvI+8JVs
xNT2grIrCTNGBCTK4gc4M6X7mXREM8AzuYNhX6gcjX6Gi/rwQuqtsj1JR2gQT7O5
aybGYV/f5mndwhaazOVU3NiqA5vIrivJyCHIaPmSDfxtyYoVIkFWC6QXJFwHoEtZ
+eXEkj/9B2tCyLQ/lMY8k0WCi6c8G3/Hnzq26oqE8Ta7NDCeKaoBdBpK5Q/dJZgV
rAvsBVObUmqvFGJWYwuvhY7ltFjxoWwekaYHMrn/v5OrBHwiv9qrfIqLp/R33EH2
Q60dlN74UjD8Y4R49khv3nAvfQ+k1lifPIj7kVo4NGIlomfdMOn1KBd5xTBRK8vE
0CXNyoH3E9lkjKthT0r/3CkOzqEoytHe2UhoBr4RLoKiYvpkzB6VLTN83sg3OU72
FqQ4fPT4O6JPMV6jcyzEq8m6OLKAYTpplQyjo0kXmOvNznkQd08J2OJYGCmmWKJc
UulYAEPhDko5WDG0pz1BE6jGZAynmKUZxWwz3cPZ0+fUgzBO/YYa0a2LCsRkfAZ3
9aCPTzHGtv0cRbS/v//i1YaMUmmpqbErlEXRs0wMjTeKd+P2qLzeZorXro87eVbY
mZHARE6DWYWTxuM0HfTzmrpkdJznvy7VMrUXMaNUbS5kyzxISYa+p4CALXPChwo8
Xq1OwDZ+HDhLu3J/Bs4t9u1T2lWTj4Tn2IyP0KjVe1pQ4LnPVYhnNVqhApMx5mlG
chDZopaeQcNyaXIxqVAr61SXBZFU8dY6Wiu3a1SK0a2vdckDZJWFsxLRjVlg5Esq
pjuFrTXeddIZZBPXutFWP7xN7cSg9VW6QnQTi/0ntver/OXQ8wI+XfwWvJsjOcn9
BrGuSuvPkoxgzWvOST5O3tf/rcMu6XIrUXYdVFHhU4aUoyDz26sjGKebGX+997Yj
C5syyhwDGbMEnVvr4kRz/TSzq6UcF9iEKX05HS1MkI36VsXz6Bw+BLEtmYYJ0C48
BYmQyUVJ6bpT05rnkdYYELBdtzYXNrHBS7JC0uHXG/d/nrCKh4b4YZ5nH0dYlvKc
1hFKDERitvTjd7FoO/Lp1S+d2eamkkRa9pMR/bsLGYfUA2tUyq4CKTZH2NuCwVUD
kH6DjaDP4rsbhmlVTwiRdKYo4BNkvB1VBiYp+fp7PsytPM9TyQeloHmDtLWwpxTN
9G/RcLdsrmvVqi7PJVbiMEUNY5WeOigz7Z6e+5YmsbwLOzgZ337/uHWVDlzgr6V6
C9+R32q59sKFCKMqiZNt1S6x1C74uS1N4cAFxtjnYk+PlFYceDCDErHoyCjArvWR
ofkEPUciNR+sWIJ02Lpw82vVYGkgFIjl9vCiPBBsiF0k4exg7VcXh94Tvcw5QDJc
v2UPeMPgw0l2pmAIp196Do2F+N2goTcIMuiSu9GQsn1RLlTI/pzjsJr80/9dDm+W
TmuJx8a38DDy65NZw1hsQ472rvErpC2TjmA/zCUKHhP2MTvqdH/a5oPVtZh6o9Gm
YH+FjpwbJp49TtgnGnhZ6uCdJj4jqeatn0GgrGEUR/Imxdi9D58oUymxlLSnoNq7
akY6m7oUju0zNVem0WqhYuNWv5Id+c8lNw+jjOWU47ByI1jSPky0Wiggr8I/ULf9
LJtd3xSyCH47nXEuipgHtRdgPppDdeoMyvBaqBDEzF9uqjH3zpskNn0PYyTbGLDr
KQLVgs+JOqDuzGorwJvqGzRfqEBZxbapDuvQp9TAf7dgOymFRT9Jlc39VxlJEhYZ
vqQjg6keKbULNYuRVAG3xD4hxJD8916OjhAcLCDyT0j+CliHG28GioeRwNhozZSQ
F1DTUXyt/dTC0Wv3ad8dI6K1+fLe4b7RDivKY77jz3C8DMLSVGW8lGt0dXK59laE
gZ41llGDqa2T6KD8U5ghyhN4YllkUa+LILoYRmhh8GsTtT/Jt4MG04qciQ9SYRPQ
HTTHBG6ZJHspjIRksHpr4eQ/067U50apVRyYAJGukYQvmuTBP6C52NmNj04REJsB
5QJbSF8PW7UCjwVN1566g2GNoAEmXHYQ/Zsdaoqgl6cdl1v/D90e03Lq8NTIp6G6
TsPZ2k4j4YTzfhK6NRX9gTwzr9DPYeqYthNhnChffoJpRiBENq1zzRperAA3Cp3V
+vOradyz+iJB/xdeYs5O/pTVIh6YOlq07vFzkkjawdhUzxQRBXHbme1ohfVJqBMY
6wVWcERF0xBkELB6LqNJow4nsf8EIppHpIh07IO3cCIozMtalbWvSemQPKEmlX7D
d40L3BcCj/zZNktRr8pgWMNwkJyIh+IGBryNpOvpN7cMtLfMelI2LxRU++URPliz
sIb9Xp7Jmmcli3gGWWIAa3navgtMeYFrye3ODQUgk3sIAQeskaI0aF2p7RPI13OP
3XXjnVxIVLmQqGCAZbWSb0mse51Zo1GxYI6fCpmXd1+V9jsdraYlAFtauZHcFpFP
WgY2GVczUqdN855d2H98RngXSIdlnHlHevw4YcsB+QWntKqprCDsKDM4hgU7eXiQ
OwV3Im75rHJkCRqIIft1URvEJGC1xc/Q16gtNGkyRKjHsS9VOE6bNch8GCfZ0eXF
nsoRqKSEdCl7yzln2vkZ9noNoTVbV4QINQihPNKYrf8WC5ZSAL8EBZEc/J8EhtNt
VcWkae5AFD44Mei9tUNPe2wNcj9AOIQ1jLkyGpDb8+118wIvL/3ti7iVoEkCDUab
0cFy4HrcJcUE3y1D3veBkas03TTGO9iC/SsG29Df7xuIA/PdhYrKOLe94Z/Cp8ix
xbb+AEr+qNKZqvejKkRbL6l8PymJKmbCUJ1jPl0ThT+eD8tW//kmUiBo//9UhmVk
4QboivzxKUJKP2lDLzvh6KU799YfCjAKzU5daKUhG8jnmy2Um2AESepjpe09UVNc
JJXxNFm0pQOyJ9Bgi9/Q1dsRdXVkZj9KZISsfoW74s0r604CvsCe4CbbsJxdV0Yj
rM2OXVtf+5/Ox5EWCA+DrcVVX0fAQxBTp+JXDC8H6Cb+ycqbRSsG/xM/+1OFsfuO
UJnU/GlWogTt+YXtWffo4Uu22b84KD2grn4v/fBj3pPm70LPunCuYY8lGifrkMk1
dhCfwcb40syusjCufDIXYpN5QXPbeOAlmXipQhFzeTwUpNP9UJa7SCLtGrlyDmsr
zIAmF10v4+YcFstbvtSrZnKbm7LVysyPr0ybHxHr2Lud5g2S4mgTCgMhQyTHj1DL
Tp2pgYOKizHQo5zX1lM0/kSaILgeB9eClUm6elH2FNmhWkY/YN5QCNJj6PPw4Xl/
InsABxTsZu2dCPkV9t+IHCLQCccJUNz4YU+Pu12X22TIPBNogafoVLjF70LPsLvu
3DcONPR9ekr1LDss7Q0TKNWVZAS0S4YVQFX5e0ei97o79MOkknfEMKEuKabYXoPX
BPdSzfHEiQuh/jb1HhESX9Vb9oSi7p/gNaJd02fgiES8Zo0ztNQ7o51IZfMw4UdO
nRCNpLb7qYYVgoSeFCY7zwAJx6JY2bKzSsLg+7Zb0sE+sFDJczLWJ/rHZr7FcAuB
vX9o2r7dtqa/MXoY+f5iP+F6RBlRAYo0Cp0hlWxLK9yPM4TR9uXK1IF3G4edCWkZ
wqe96qEQANrWx1EENGqBVo8hMLu5JwmRPcXo2DtdIoSjihDEvvF3SMDc8D9O8MmP
SauzXHVIFrLYl0jOaQKW0pHZ2OzIhTwVZQgwbcimIEI1lm5QL2D3easSM/w/xWJQ
689o4bZlZWzrIZ14qPsz7YU//hLc9uT9N4tWIBcBu1X/McG+1Bdr++jHacex4UNL
v9pNyiBXv2DNq7BOSXAOVA1TlhZ2jJK3zl9VdSwDcWFJd2atJDdA4/O6jbYrJYSD
jM6JZRqhWEIXSnJFgUvnm/uP1AC9V3xAZiNt1jQtONQr4DlynVje/068rmEDrFWY
D/XwFYeCVoQDwoS7YyQ2wfB/q6jogYDIp9oWOwzbkrRRLp24gWTDZFdh0RqVwYZA
qMGHJz9slwt7pgVuKoPThu1Gvj1IF4N3n8qEkbS0RnsmwKpxR94JftkB5MixcpKX
522pH8hoK0XrzCoOefPmpvwAGpPJLtF1WfQG4t88aDPdBs1vyM1JeytnJ93/RMY3
HEcbuhiG+j2Ms4DwrkTEbru5lSthgW/ziSzUgHIMH4EE18suLTQl/ggx7VOqzcDe
UEFZ4IX4J5qYZVx4DYTRRxG1OXLRH5xCRx3mPOlVrYZt/ELGMhHx2XAm6JM+q2k0
PuqlZJhUusxHJYMSSqPBT+MsLn9RRLiO8HPTf6obXOIfe0LuFlaRzbJT0xybtoZH
mMAqQ6oeVMWHX7IwtBHVJTeeyN21j5+YrI1JmPlTwYqCAiP4rfpw0Y4xqgEnUFBi
vQelz6DiLWaXpthtgoQvUWCeqqQ+31a/fo1s5FlMTlbn654Upyo0UU1W3ETyiUqK
/Iq58AG1FMZnQa8Sz65nLo0eRZPZzFZwNRht3sl2CxMG9K5k6ONbPyVnnyYlIyYS
mqZDnzakO8RLsaNYOSJvEDcGviR4k/8T62fPP/WJH+1ots07exOGV/FHn8jXirfg
zFQfxibUlDvN5BaMazGxUDZaUy5kieP3VjGOcffAIfJZ/IOsc4dbIWHs7B9bRO5T
fbR8JhWxvUeKHlmeikZ54VNmJVsh2H1POCJFfFJK6gjqqJATD5pY5ZWRRFcFI0QN
6O1fIajDv16CvKmVwbQL0gIHlEsiMSqH7/qbZB8PX3ChN9r+WOY6Ddpe5k2p1YGr
v9j8RK3zzQGKaGpGriQYAMSBoxP8J+MB67kbN+GGT6HNHHaVK1hd1KqyPKIoB0z7
wDvyxMKQsCaCJtoxFQHxb18cfj2ntV4l/Pc9d0BDgIl1QiI92+QKHsEHqecD6gyc
5A3r4WzVc9PR0mUlJsUQkTIa3Hag9ZK5f06tO6r+Y2vbUhRT+J+Th+pgNPhPKARk
u6Z9iRIM8SiZEvMTAt7RLC9Uag/2FJXwGnOeraKtDxoRBCDHSUcITmhwp7F8DuGe
kXi2k7cYo71fhqo47XJYoYROCpa7/29C2Yb9jRzUDqfgKgF11UL6CUJTCYVyQAWx
ETGoFq/AjCL22116jiNyofrZvLvdbuiixnubCYyowSacGQge9MtzQWe5yvSP0tfh
iX25+r7jQoYcElEZ2pamfUXkxO0f78H8RhcNv/xPwceAY3mw/+67WCYvDO6tiqDi
EmsmSdMc4fT8+zHLqSTtpM2HhFaXaidFRk5fp4grx84NsjQQOLMzHrclohPHsV96
JA3k/v8/mmOmE1EVTZUiL3KLIQOFOSlV0YnCumo3S3WzyVQb00N9kSEIeY/F6DfS
SWMf5zVH041voIxKKg+yM+C5J2OzdVObj+jVZAMk+7bs/u6v0mQ88Ru9dKuKI0xY
Js3DGkzeyhPG/WTMbwdv0A==
`protect END_PROTECTED
