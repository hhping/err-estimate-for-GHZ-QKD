`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTnn5kKzz5sq73zFhfp5mruZegy65HW7uznBcde3UeGvb2kLglWoOQt6wMQ57my6
g5gb1CDJNcsyEoT4BvC93zVtjG5NhcS8CHwZbIlPCWX3WpZzvH0kDNjkYqc2rR5m
BNmqZwrD4zm3GgJId/BZFGYqVN0oA71fj/UsS2a3LhbIE4j1UM+OmKeuhC3d1KMX
NV5e+qrCrzUj5uRd/OLGpT5hfEp6AeLbhH4uF+32VpyXZyqlOfu0TaNmFbPe2A8u
y6szgSi33FJOABCjZ1pgRQWPBT+8ejvkw6rQpBq1Vm7sdZvwxpf/GXRzxF4sn19B
s/S0Vgsf+NkrkSi0icm0LCYe0xz9DQ3wAHeechvAEkoIva/RXkcivaM6Om07nlqe
wFNLIOseVyKIVl80AabDomnNBgXCemE7+IoxJPCK++iRgvslfFOPN58aT/UnEATM
BnfjKafzOwxF4lPptIVgV+eyQEGvP5ymM3vdUTltsoNn8KBPPn79HUgEHkXRbpHN
uD3NuYYsmAefKhQEi6F4hj+kJi3kiiVCVsXwA3QmiZjI41XlL39KjUb0O06X/ngV
9ywDN1y5Pr0ZIoOyp9dGQfFqyh0LTEcw4lJjT2IHtsBsScgz2jrB5aJM4m0qKwqg
+vXdgNxEaCVsApmqurYx757e1WvzIuR/+weP41AWox+SUSE+CRor6pkAl9tvHBGy
HOo9ZCFTLLgm81VcQVTJMiAlLZJxctWT4lTpdnnhGLrKUJQjKG2DBIIXCZ0cL+zz
sDMsNPLewAMRx1yaq52goSKGR3fh9iESRr4d6sxCMyxDwTmzFbk/025gLtgOieuv
+sCH+zk9t+9y88veKNKztNMf2fdZOCKts6F39+B3+tLoFuHe399EsH+j4Xg3NUOi
drEZyLUHaX+ggxVQjk1O70JHrV4UJ/7M2T2pLLjtVn90S+9g8t1Fi3ZoOVpBVmJs
MYVROO2LF55Fi+P93pV8rb+Mh7BTHlDkmr9Gd/qxa5fbxO+R7ylM/+RBQh/TDeCK
RROyLlVesyruS7n9bUTeFELiQkV+4QCbFirqs0NQmS1mdW4P2WUO5MpGWMFBuzoV
JNOZq9rfti3CLo79dUSqDFVjlPUxXQwyrDUgKoNz71v+VsLyDvt7BEI8fq6HWOGD
ZrSgALLduomXxWbaB+fhJLWFGGxx+E+Uz3E+Gr5XUrwG6Nruv+B4lHP6EYjzGexh
MXEH+4BLQU0TtdONikjzTw2RNUAUGyeiPFaJx9Vw7GwgKfCSco30YUC1AEuKGcfq
FQGlDJTQB8onL7HPy6cntvbjKZbq+CdCwlI1j27egnUKptH939vmDEMa8f2YBFTZ
XT1dmfrSNiaremmxj2W5v9uiRYpxyod71E3lWsY0R0v+6fAe+FkzBQ7REyAnseh8
HC7Nr0HwtXCHnfMrBxWCqMd7hr4v1ArG096l9MIDoI5kgNV3fyPel7fDutLsR/C1
1BJ4olqqeR/EnUNZnPVvDis9IUNx8oj2RCCIWgfNWUNsjs1HBcfbiHXvOLeWVmgo
hkBaAA6hLSUdgkM+gs89VQJZ6Ge2449ZCLLUEvTCq7rQblnMkEdrCp1H8af5BhMN
DvyJS6ib8W9Uvnshmc1+xkmoCf8cGMFufIVWRxeYlMReF9i2TBfzEn0tCUxSLsYP
L9hpj9CTvN4qRaAhecjyB2DLxMMN1mQ0zqvXTTYtwOf3uUhlhrZjqzyLe3t1YIqD
6eyPiSngXQLBeVJNlPNTmc02Knq8ZK03kCvWUWXsyGCVJSpx8pBi/YstixZeEj+4
1UKo+jpGb8SVdNq/06+HxL08Pk6ycQXM5ocTHxKkx8zP6O8muZ6rV+dCAL9AGm7u
UJ9PxPt3fzj4uV7HY7ysVdWu8LNYD+EjqbuXYCFxEIzzh0SYI3gPnU9UGXkZu4Bg
6cOhNcpeMvnNsc1Pb2aXSP012qBmiNGtMLK3SFolKpMEfznotRiU5riSpiSS4Q48
gT/xwFfkhiNzQsOCrGGamH9TihyRa8I+liB+nqQPLve5wHZZBF5fhFNx+6eYzrnl
mCTQSWkLG//Ww2nLfAoVmp8LYZYyxGROfmmBINk8qQtMYAtjZdUV9OHMMP0Q5mR/
kqISp2s5m2WrqzROAjjURtbT8vM0PVYgvI1in7ZqMWXaVxvjVMxAjbzqWzVB5V8v
zGdbv5K/fn67ju/dsYgqFLgzPrF8nH0g2OniW6BRmY4qRqcCtE5SBYglkBJ653nM
FzL85sSPgDaHO1h7oj70Q6msJFKY5EekH0A8LgBppFHbi0VEDz5IcO3qZigSCX2N
dnJCXIuHJJ2K1QrBnG/yXJEFLICweHqTk1O/WXhH/dHb1mSRDtZOzuGvVdC8fQ76
3asCwgWI8JFCZdtqU7KFmp2/7qh0bBrululHTCtaYIXVlbznvAfWDr1XX4j+u9af
k3IE7zBYfVfG533FKckby45e8owlRiRlK13vZz0oE6YjW/GEq0XkPPKu5HIV4lfz
57e1IkBDvFvZt5utgzP3DpWLidL0UXP42mpvBuU6IqYHoxgpqiIlI21rslLc/y+O
nno5BspJAuLFj4FDlnP1giA5l2X5N/+msRBvzWnvUJGr3hqHyn3ocBD2/PkuKDpe
eHc6EGEOPAjoeSISsmrUt0nxAkoOKf7HWwiOGrTazh49Gc0LB6JSUgPtAFAK0Ex7
/lb9fvgJbHWsXc6OJzmuZrWlyeT4tVUmoRJ6U399fkSqhGZ38Y+XpU0WO4orlegk
p6B6HWO/IaD4CWk+KMNAz6YLk5mQqTAF47BUC2Jmz8RpbhG+wx8ERkGEv4jWYOFy
yrTcdaRCOfB8fFAK7uTfAYbyvXaSVcDFyPqXeoI4FMSv6pzpyn1hsuNT7R1x3knz
44KsNwFjgRQQgfkpGjT+DWvIcPbon2jJvwg0fay5ymojDEN5HwFFwu6vrVomrYkl
sHveWsktnxogkvX+qJjtST9bmMsHiD/aEXY51zgv8+17LHZV9Towq1A+7d/fuuWL
w17CbqH4yQWz8wwPqfFYu4esSDE+cuAEmTHSkpQZ4mcZDN3uj5louioLTUFvS3dP
T+8GBV7hV1btDuUgLdG+9wF6VeRuwUyXgCEmfiao9QMKUKvCacA8zTDgRrmySFPj
tHeq7vhjPRy1ZQ+xIbAFrxXQLG8+JunB2ldQHTWzixwCeNqjcyQqYvnYcGeeC2Vv
kHjxMou2V2pVs8OqaE2NkzhBW0pZFuBkg6M7NEmvVj7RMMZUqXwD6CJm59yrmZYE
FvOc8F3VY3dxfKnv7xBopaQ27IOJ3UEo1zNq5S5KjX9q4xdtCF4hHzo22ywUdgnS
nE/cgE7XksUYwp+W99UkuUKv0+YdzhIwk3rRPkx65B+l1T7AfCgOR57wzhKaOmmv
a/lSpi9RjCm394QzqNhxAoRJ9i2x6Eokv/orbSyRYZJWNv5Fp+ctSL4u23sYTk7h
qcIWB+U4YN5vOvnPj1eiznekfafcY7dPVSjpWZY+7L4/mZTcEUC+WDaEOcRwAhIa
LCYo/hWDHVIOOzDnV9rHeBb4SurGgOSD9Qxkk7WI+tLDDPySA9FcLDZWXFNfGGwn
NniQRCqXvoFmUAnbx5LycX9ZZVwmyynmtmbYqDlErt8pskeDE/U7htmPsgD9+Aim
0bmto2tr0TXL6yDqoKHm537UuHNPt28U8qhzAjiY2XoupIi62VKETxnv+Sc58BfE
9u+X8VDvXJW/WO/QJh0uwENqGfsxtys7ivu96uU2h5Zgn9oKZKe46QaSIfxvcavU
SeO0cQppsf1W/pUsgzXPrKywysE8pIe2P6M9XR0UhOt24luEyphORRSzVgxCTQN9
ImX74Nf1RW5g5OnhFdqn4JrQ2Yr5ixjNkVeCyKyPVW4BjWTBs1MaE5NVxVqFkg09
QN5ERlmkUEyvNLBBZe0OPw+5cc6XnMTEgZ3QD6K1ZnYvCebwbC2V74qhqzudqew6
3R3amx60Fcmb0SzLcJFT3SaumtxmnuWVJh5SVxfvrFqXSsI+6qzzdHnsdrnfLp76
x8s5N0dL5p3lTPpouNkNYItlJflYv1V/pq7XJxoMoljqsVkLP2oUwDNR9WaZQjhz
so0IYTrso2I6WY5FxZzH0XLyWDFxyJBH5fqNtvqnh7gG1rlOojMD/V4uZv38ZEOO
O4E6QHLuZ0eeN4+ESAtrE59W+QfXC6K4cT/3Df4ifKucGoI9i2iOA1OJp19EkNJD
NCGYzg0pVSsIqJkovQAKSsmsCQJNQZvMwbsrJZ2c/6k09DqarP7s+3Mm016vDnWg
+UD6W0tdh1D/v0/MOxjOjPpaqqdMGnShUDNxaZ0/W0VJI11S8zFn4EmQnxT45x3j
2sa1DNI9kGZYRAygyS/JmOeXGXEz3eLMMXSs4dcDSzYjm/OyabXVzJwHZSRfAPGZ
f1Oa1vNIWjbeAdsJvoU09234gP5LJGgKRNmdRbb3UbrlhfF6z6KmNwTh7aheV4IS
o9oiXClAQ85HEES03TBwGgWgvbanG+c8Q3vMSYW1bRDBW0MCvPh7eCITJ7x4moIr
+5TI7jGQ9Uvc7PWE7ahROkEOa3n0UjEHetVHW2Lp5yRr0NOV8rSEu5+TV7y/qiOM
USc0IfWDZr8F8XNaMyfGP5BnKe/Bng5k0a+z8SDGu76AMcpSU2EVYJWUCJfEhkZ/
2W86hX4rtamhpsU0ZdEyuzlOr6aiYMDTrteLZdjGTWrDD+muNdfBTq1x8iYMQTdb
NIq2T5sbqCBtMpIhxUcgApUNn89/OKddrn2g1YSRJabsNYbo2PAy0LZ02p7QxhNs
oJ9/L22mjLYfVDOpm0ESufuarS5nXzCKngNDmewrdvEvErdE4HMkXl5kwSBc1e8p
fBqO8uzTIyH2Mhh7R+Rx1o//QMLD0y9SZsfRUTzLgq8x2Ebjbc4+MAaYpwczlzON
noyEcVpuumx3ilbJGaGaEuQnK/oymby2YoVAaFD6I0k9vbCP8zWfSpbJXwdAbI18
Fb1eDFTXieptLCNhVVXAUrKTYdedKYiJDumWzWJWsZ1rNsgXWn1rH1uuILp+qqOI
Qrx/kxGrKLgFYz7Lk9+aK53dyXKw5GXsShfMajgTY4a1dgEXDtftINhpmHFKcnLF
QffECqGCGfo+Rw9IF4sjHDsoj4d8HRkFbAa/qkd824kAMT7jjZ6cIj7UOdrDGndW
7cklpCX4bbYdlOfektHcmxqpXC3vf67op7KIoIMTTu6K1nrd8cNL5NPbacOt68UR
hmH0nX9VACqfnMrEhbZsPoUNwzvETGkKbjHSjLc66B4VtkzS5puMpGfjeFHaouDF
fEWXcOAoT3DHadzeSPBrYp/MZISdFKsXETzYrvv/vUchE/JjMUAKK39WEjYc/QZz
VgcRkt2+nXS/1fPaseqqlM+G/6zYGlWUzjbzgffv5ADHjJv9fuhwzd0J0HZQCdYf
0zneFJuyNUwR9YTaanYLnK6PEdAqDm4uSCcYSqQYI2DhMTe6RK6Ab12nCAY61hhB
CHqLy7UPByNcJVRiYCIZc2zI08LL1PI1UayubORQpehE/nuuXKy8eBSaBoBTlAuq
OZeV3nyvTNYrXnqiQT5HPuwmPJqa/44W6vjBUDKcPGitYepko1haFOsFU+/Za9D4
QOk4JmTmOJ9dJWwzliiRPCFIcAxB9v6Llrx/NuF7/72TFIUj0t9S6OA7q/W1HdXc
iZJ1wL8IbqNxqhV2dURBVxrdR3FVxsNYkp0Zo3lvJp1snSg9ZyPho4xhDCoRuE3L
FlBoHZZ3h+r8YItxc7eJp4TdT5dy+lVfgYD/jlFYd7pqIF03jkVByrfwb0VavxvH
FKGm3u8zuCToXXwIXIW9RFk2w8vXHKdIXxoSSksJ/jOu2j77+gs4TE4kyN/3jjT9
SHTCcL036xsNI0dchndyYqzQxYjJP8VR7WeOoyQCo17AE8eWliwWpMhJFz3r5dun
78xWCQQooptye8dMCZm3Drve25HEoIpSq1RRHmxsxnjhlbDopE1R210QKCJRmdI1
1FH8q4PbpNhWyVfBAm7DBe9HTxkVhg4v7HThAPPs7+rgjgdQ8FsWQiierZTzKlin
n2kJDWCFU/xCWoFPIudtKJnPaYwlCKfQvPSHc1xKQOXOx2pk+y27Y6VsTG3TVCTB
Skld8XjgCYE/qima9RdGawuokUZwcb1y1ozMQaMTXW26c9UCZcTlw22dxxOnl/OG
5fVNjCFxS+S76LOAuV6fUfWx53Vhv0EBz4XNX8OcUalSMhOP/bIO3hxdlbO3IsHY
CyIRH6sEt6J4TmSMNQePA92YWxgNEME41UKaYqVxHNjvTgQRRwt7u9YaqkixUZ3S
Wm5P5Rqt0bFhw5D5qcVMp1fTXjykVpC2shv9YUNUPr3+FTFsT70ESHyJAxo1ph2P
AOUpffj+PT3NCG1q7KmswGeiSq/p8vaenPfKD4i6yNc1FByuT1pDKPaSj/dF0gg7
dUVo16n8lgFvkcQrEY3mJhj7eWUCwZN0IZxR5QAJrqQIgxKXIADb89AXtWdfsrC6
cyKvWKzOL1dICheJxeqbVznF5pMo1KHKhEc4ugo31RieEgUefzalaKASjb6Q9x9a
pcE0ulmTfTNFBh4QbZuyA2M1XHhcw66d06KKdLU0LcK+ECQgCBQkfCl2CC8Jbe+2
CBjLTms+LnvX5VapQUSoCIp0pVSQCI/WqVG3ld+6g5vzRX8aNGNix6VfFm+TIjg6
NY5AVMK+vxZY7DUTdgN2NxAtjmzv3PlPdHXZXYTBFdqsPPqd1uCLcSjpEIO1LFYs
m223kL/ksanqUqxmdNicMNo9CpED8+FJg5O006T5aFOVzbVhw6CXdySDCdidPQqU
/cM1xKF4jKPKp6Cp6vLMg6TFWc4pQh0/iWPavq21ODqQiJwDyTam4qjdYS5Sj3qP
svThqxtfgO4Ym2nORqg+KIAMSeDrdjkJLrgw583SfxhzrMgVVEEo7yupgQVlbepi
07VOAIqCtYX+4inLBPBEjsfBaQQ58MnSjg/6DM1wxBWuhAcllqCosfb24zinT46G
dkMGenabKzM6twrEFqWBFo5ijXLZk6FaK32Wsvi28D9jyApyZ9ja9+AsuvL6jgcR
4d+SV8naPMaJBn8qs/qnPCQlqZJyE2P0kulBT94H43jCB1ckc4qTrMuXm/ybL/T4
BCx1fjuHAg1Rprpl/YcI//DDco51jX4c74ktSvXExIYNsMi4sAOqWzz4AYgdKM3E
n6Ynj1nhMdJ8qtTDwxbBYKZvCFiFNrsx+7KPB4P/UVNxp9PWdHBo5YjmlJRpmRUn
uewI+R/NT3XVk7InYPZHiazTz2K82p7XKCtlJtjyrb0chzr12s73QhmpD1HTYf3w
sr5JMb2hERBHo7pEqn0EvDFuaZuPsKDv4Urvv9kzF1KZFiA1zJShEblKnQMJ0v3s
+ZR2IHHHI/JKWbwTmt/GHe6AuVHWU5m5PRnVv983SgcyucDgjJn5/XPtsceJMZnk
5Lbho0UyCcZW6sQTyM4vq7vzh53Uw6IOazQqo3e33vESxDUDbIy2pmQ6UPbPFkDR
SyGfXkFZkUwOhYNdbjR/5tPlqr/Pa3EiEWA6OzPmLymBFZlN4cWse5OrNrUbGZhx
zJEDFpkdl0wsd5z2M6CdH8Ec/Zz+q4KcGs93Xv1E2QlgeDeabLRvGbFvu4AZjibo
RS4Eh6PmX9E64K/dVr+SvlwnbRpiQeTF4O/4yDO/LFOb9oIsBQjEQYcjWSTySlTg
jYi7KI7t+vKXlYp2ZyRrpaQCoMTag28L5xsf9b+iy0mlnQNC7crabhpDV+Rs/sNt
m7FntbEFRLLnS9Zyoil7DuhABBi3bxJeCQnriVXDvzDkKMf6QGxMzMltuy+gxAcH
4juCg0AMubMqhHnO5DnFna9mx2S9cDSsesNBdxWnItHH6RcOLbenkqZqXneawvc7
dE9MAD3I6bA1rJOxCKPAmOTCMgSw2urJsTKCI09krUANdmEYL2J5X1EiNcChfGOm
cprO6Jqbh3V/FwkPWefs4vj6QqPT4QeqQqIYHaB78A6bTHth2PgPr/+hrQbofsRh
AS+MiDRLKTVF4gRNi80BgO6tmTPLHSW2kUYdKKYliBOLckOICRbvVEts7t5tivvq
SlGcs2ZLvaSoHdJSIWYe4GiITMe6yHxb0j9MOTCBHunFMoQfRxBQSiZHupx4R6Ne
XS8QZ96otyILxNCL5EvSq5Q3epmKD+ofj3CpnbdJqCmlCVA6XtOcf3K773EWdXG9
cWvVh57c6JWXhuqwqckXDBjX2sO59hvHYEINGQqoZhzw6CmKr8cgiGCns2/7ti0d
cYxNm+qJM3L5rBQglljWHWsrWaflmSiNEH/hgnaexWdu7tUubUfovcVQHLXuoy72
+3mC3J4rvV4TjYGu7eZttfYwOTGHxc98Xnqqwb4Ii318iSzAZeBQ/MEP+7ZBQwLp
bmLB305WCb3qNP2GiO7R4K+XPCOYsqIxwPosIELQnIzwAOdTjM35+nN1J4OYGwar
fstqdqcsPOCGN6rD/zRH71DxzVLfsNu+g5qp7jKp0FczCkGZdR72/sdOBRMjOZGe
LUh1BHnbEe9TSWHD9xdWdbecNqs9Vi4SLLg326fKMtlLM8NfMK504PDNnmPYOFRt
fZCRKtgESo4/Q50mmbp8Jr6if58vfK6p9zmYf7zrZh/nAa/03hXwgvAhnQXwH0Fo
hKlRzax/5QRMDAEZ3nkK4Kg0DsZ+pG7tBqJfPoKOmQYs2hERHXjpjWPx7tat8wA8
gzfkQO09LWd8cQn/hoiqrSpCK1WZV97pTajoGbSpDiJWO9bhI71aY/vJHKHhxjua
TNgsoA+ylYP4DN3Rm/RjiM21FSElErQUfckuYcCQNfQ2kNPtYu86bWeAEe36gDkn
KKdaSCdEa2qZ/cf2RXorMF6ib50OzLedbMGcyL6FoetzqxR7+SPPqssJqHqaAFrY
wWRRSFq0SFa226hcy3A5fBqMd5YhWTz77fdo04OUG4efqffbE9tav+6qM7QOaZE1
Bl3D+HneYvnAEEsPX2Xj/C9soRpJo71l6DovGG8K962ZgA8DobwifTctp/AFw2Rf
y+ap+aOt5dlSjzRsz8slqByUyLkxEVStByVLenRQ/SopFDMexot9Qsp3m0SRb+SY
0ysvV5/qufIRcwvW6bcMvM1aFoJYScNg2McIkbsTZ0aWbj0zdqDvIhZI0VJw84yT
UWMrnmNKBjMJnXsF5lw6XIYUw7VTCT2zrFJwKac1/zhLprS18cHZxuvhcbfrn+Cr
+0PodWVhQOJU5mYkQWNK1yOGVn8h1QhUkNm4u1b1+wulXGI9ASy+VQOmZ/aCKdTD
t1sVlKn3Q1B1DymX2tvi3ZnL9gKbWUJXxquZ3QoXnu8G5lrkIBhsVCGD0ZTyeflq
i8LAdbNKY4i5Z2NRu7gpLVsDHZfqZapGtb9Een7bIKByRS0f8beeva1S9HzyTFs/
XhpiNWJr6VI/OpcrpJXxvpssLN+ZrlPZwhz/8skPk8+rwGrza2Go44Szg3i3DOiv
7YD0smw5U8zggu9KjvhpZDJ/QsA7zQFtgYDPTVUfJDzLfZN2P8JD1fbagVVZuL69
KqHOiSM6cgM4lq+R4RFCMATODeSjpnlT6qO8YVl0K/6rdqFJvy5RQqcHoL17BfY7
lT/gtFZXO8FxABz0NrJuHG0v4achHG9IbfHwEI8zmuvGw11mjsLDL9uik88N0vVa
0VsUyhoPRBdRDcdJEPFW2+4G1LHB+HNSBGlXqeCBzBxLjKPywEihX4YQOs0jifax
NcmiOEl2WPaWltXg+Zz7kMfbk+yupgqGW8jW9aPcNUWXVZYXwa+AwH2tvU2rlYtE
6WwdfBHg27B2890nMA77Ay91skK19hhxT0rVgWhtS/MGdk2HMbYunh3H97v5RwrQ
cAiTAg8kLNOCfRihappozTS4GfQ47qytDMzsLDIJsGOoHLRVDl+KCa5KoQJKdyc2
Kwkh4UpEs1yF0fGgiIa7S/N1NvvD+aS3DmxQ/lLnXHjPcogbrly2jHrE/WzL2Ls5
28JFuSVrEELW9uClietoMPcwahTSs80H3r6G+ZVhzX4qHVIgikY/h/rKf3JvKZ76
dTBjhiXCZtGOqPIVsphUF77EscTWCIIWzSYUfQg5ulEzFpWKhS8/d/6q0Izgl4Ek
XfaJPK5dj/w2f7SwgxNDLegKuLkwOriAp+rfU/iy31KYKoJrd1Ju03AYrDFQT/dj
Uu3XSN2Vp2q4zVrjwp3SxmErnJmzV6Ko3TrrezmuoHCSBT9bGUnMyV6LhqOYrrPu
1Agpw6sMSEMuUesZKme0h9ttpmilJVGm5zDx5auRUIQogi0ys0hW5Qw7R03Jpt1h
HVAZ9Qa3v/DONAQbqHfDJDxHS06YWe4MRRJvoggqWueLeepvS2Gh6UdyXjE+N5b4
25iRyDPn8p+MMyBQ2bn87EQkHwDgWgInOtoivvfgcvuYDt6rr2cf0Q6vXB+rFF0O
9jK3tX5WfC2NpTUM1s0y9QKurFlQ6GjWho4aQAuscbZn7YcQmipTUszqqVHf7N1i
BgzvLjzU6I+QQpea5VcUjTj8Q4WknDF+5i7uQ4GoZ1FTW/WpD+YnAldcxyx3gRdM
mL+KJyP38iEw8wLp0hTJx82ZP7RNGVmrf4laCHZWmIF5Pcppu2Je9jxeGz8gD5sh
r93F+RP/W0rLQUGcqjT1+u2nwm6PjOO+Y/2HGfpzWowJV8vlhlGZqIwRk9p0xJ14
J337vxdpb0bI7XRVViEZpEYhi9kBWXbYC4ql3VN4u2LN8DYkCyMwVlTWB5N+y8cF
8Ybs7slcJh8viLo/f5uqkL0z+HkvtE5oBT7MdbaSwd9N13/HplgbqYgDZTqptfVS
gMDJibnF30YWN7xRPtaNVTVpcOuL7Kbf/bZFt9iAXt+MjIr3EhK2RpMOzMmADWDN
THDF9VKU2dwFTFGRH7CuxRrJKQCGlHDhMMXPNrRkcQi0z2ieteOuv3OSQvSE4BlV
DpEuNpvXdExLnR2tjFq13E3Z8L4cPihU2JY0HiVwke9q+D7P+NiTh76arOLWHGWs
z2TmraiO4ThOGaai0xzgFdswMEnbFWGnJMTnVuDy4KWJBeB+e2Iwcy38BpENYG6Z
dqhbVzv2g/XL+xWIuZ79BFST9QZ+XG6dArA3AJHvpGwSw8L6KVXrFm8T0JWb0WwO
tnqcvPpmISiHU7TOV6uALFeFle3Y2O4+gwFwmzoAiB2e+UTSY8K4VfbovcIaCByD
diESFn8SSU+UA0C7haLTDLIarqk0PxRUdqpFNJiOXg0Ql3uGDWhfXdkVetL1s4Ae
XJRNlDW9nAiV/JZWk7PBWT59JQRcTU2yr9/7PPd5zjcgC/aNwlfjDfH1KIVb+srR
YSWWKa5oZYAk6mfTmnPIyY09/dbW8k4CcrfWNJCasuN5UPNWHbGTwNpNLZ/LMT3Y
/KJugoumysEYIt7UVCvLNE7hqvc4zVyVc23p35Gb9lv8K6tio4qmQPxltoI65gAR
jF7pO9PgrTKGMG+qvnYJB3UHKEjW8SF7petFiO9MKEiyB/G9C66acJbEYkVj/tmx
l+ggyy+Iv+seKfITG4jb4hORel2Db+YZBFN0+6tAyYqbaBK+n+ruOg+4lXO7d72T
JkgYmGBkmrXN5pz7xWl/CSTSQaC1jF9k2i9fovz3Ald0fnzwm+u18Pdg9qaVSKQQ
Esr8XttKmMvyHYbkjBKUgOyZ1ob0ay5w0/c5B2FCajjI8ZjUxbNqN58ntEMHwA44
BBn2gJxM5+E9brykhzIdR4yOwxm7ojl7zU8GgXUx9CsRN96XgoboiZwmfK4L8lqf
gBF37ByLcxaUYH+8THAzqN7KtmnSINS6VV1sLJ7OaezhXkHKZwKHwwmaxvK3k2NW
E8LeD7rXiPBA7+ssiXj1xTaSfBtQdu0sghhca6/7qpWv04gIWH4iP4AZTv2kN9Jz
gOjumLhaIHKTZfZ/kH/XBuZ26AeeAppezrtoX/L5DK+xK7GHEP8dsoQbODMz18Wf
xYPKoD/c2TnaVzWUecwXW7qwhRjaWhm17vgt2N7xZO5KKTVfzLGe94BQ6hqNO3BP
9RK2WPjdVQTxc+Sen/xx9zJRCR+cYACksksWpnFiTyNbmwwgjMMcXD6crrPe5zBC
4YRA7gfY8SOqxqBo7iHI8UAFn8XLaz6IRkOvOzr7cGeh3go/WsQzy7BuyBaNol0A
8kiJz/j8isNqoBGj3hGBKkyrLpDhz1fsP0OofHYKL1krDY3ZbSBaI8aNZ48MhhNl
Vw7YthyOuUymuqNIq6WiLWTSi707d5FRla8jBgZWXuomjmXaLLED4AkoJ3ljQ2zx
Wk95Q3IU1AVO5p3yWaEggwVWLTJQz+XAGpH//3/Y4JGCmlMGO/Q5kRrSpdeOkGQa
I9VDjJDgpqquMDou9ZAyR4MrL27+Anmor2o6zlUpMtnjgkTY2jYSGCSCdOASAOeS
1Q4uFDrQmqyQ1V/47xnWU4q+bbso/5kDXmQav6iP5ICCsu4mVPze3YvlAGrlb3Lr
LpyJiAyIMNYlOK/u+ptN69YATpUcqqk4QMoEcu8Ve1MzjidMqTLfcUaCaOMAH5FQ
oVU+nPV70awjfrEZ1Edr9ANXdnx5HFaZ1svRUjnDqTgYJZVsUHUp29wO0xQZJmaQ
ZUrVQqW1HESSLv0djnC9gwk4J3ywp91lXxpOGh0YL0ouupFElfPZYzu4jlMBSgsN
KKTmV7L5WliFZUuks9rYrS9ggtVzxtVEvGJpTM0BH/B+M61tNAEpak6MlA8DwPRK
0y+Xw6Qqaq+Y3jnBNT8h+CBn75XF731uhkHIxFZFs1X9Cxn29jp5pjHKQoW01Dvf
HHfuJKVYuNr0xV49JxDLFFfg6iJZQbM1vZm3ryn5Ok50ULgbDjxEsenJioWlFYD/
3J0I63hnz9mtnqMs9PQyJWzAo3lQN8jmJ9EGro+/WNUElrYekjMAW1NMihgUttZd
dRRZScDfWPphQus/aucNgQ5TiKizEFKT25T/iKMMukrlcO0adS17MGz3ez7NUKmF
cO2z4/EnwzF11ufUqWDgAK1NIG2Rj2LKoOvvw6QYWNJ3orCYORQwNFyCx04iJQ0z
A6BbNw3X7XVy/o5DwRKOedLrN+yj1IMekATeHu6r+GXZ9fpX7rueu8qGytl6SEXO
VXV0eTwfsnkc0FL8D1gHM51fUHaapvKoRFBRT3d2YNplzCQHS6cuFYM4E1dlhTbi
KoGk3tm89zaDzN9MGdsWvnPrJhJE0golMya/y8A4aQc6k7HSY3cFYMx/KB0nQ7kK
/wADoqtDUyTuNbVvyH+9CLPkBzaJNYvZeKFcG0l0AHd2DxutkvLz7zF5e+vPUlUZ
cCdJkiQUYVsXjNemN9f7AbXlsgnUY9fDXRIf3bNZzehjjKB9dTMke8p91F6xNx3b
Z5oDBqBwzw8WpeVmx0MRJFibnvBu4+O9QQ7kx98sugXzWQCyjU4y9FdDmWmfICLX
+sE1g60YAEqWv34cyGAdyGgWZyvq7k1nj9hVYjOWFbQF9ZVFUCS9GahtgGSepAhm
sGevwldUb1ECxP2O/XwOVjwHiWQ3e0Rn4lhfFU/rmWNf4AbjZDiqE3qYaDs4Z2NC
Yr8DYf6xPYqZdQXX8wUVAUqvBo+VjtDzsj6PXti3VeWIX/ciaGHj/7+6VwxV9SNp
CSHJLumbPS51WE49ElOBU/Z87HIIEls3Z4EeD4j9NwY/vV9CdF4wqNDfoDwXP33+
eB8sI1t54RKpnH4B0GdtsyGp7sVjl7Rf0TTwO+5t2WhefJf1U7IWE84mRaWJKg32
rytHYnsndjBYi8yJXbo8af9bTv9x0s5plE782GdRgcYyDYzmu64PA+xSLdiN4mih
+kl4LdJbyjgoBTEOtl3EkjmqEwb61BKdr81W7LJcYldSLayXtjTMmdFBbrZvuof3
TKKUfSRu6xtTy9X+PEKzVt2kqM4xH6rJ9na/v3w+VKGm9AQdojHQ57jDc1cOwxDy
WXO798t5HU5IV4FzNBN/khLBYvhNHLVNuq3213T3cngKahn6JTbztyWiUe+bHOlp
Ux83HFZpz3HnR6nSiwoensPSdGgscT95LJekndG8yumW1vpbwwuGz58yg84LM86d
5UclCW2f/ABL25ap2xA5CKWIfE38Q/UKnQdfhWi3/ILGALYtAL6uzyc2gIPseyN1
0oY3TdlML5IhmK1ZM5qMn5xr/WkTitSDO3mjdrGvKB4cPYwmHPMHxkDUaoeAiL0W
J0uMGeoKyBJSMLcBYUN7gjwIbqBymUAqym5IJ9wMTr5zqINbvHmVSYEhUifS1A8j
1Zq6kBSgvG42dez3gAYBk/fX00JgL2VorORHLWsWh9vCBVo9zKsF72cMAzPlTJxr
nH6Ts4WRQNbVxJ5YPPou+r7lxC2rhHc3Xd464ttJNbDgPO7Lw+HV78dmVmbqtSRC
eMk9l5XzvGnwA742BIi5W1TegO1Rs7am6s6PhWZPt9d0+GpCrl30UsCPgo9Jeqqw
yiTWb3mReBnv/GgdFpk6eapH1ZlXvWHVDSoNgxgd/bX9N98hV9Y9o5M72SWZrZJ2
LaZXM+QoEKsnNFIQIrbbDvM6wgowZMTLPvYpoWbAFQUbIOKMV/aggyUBKHUaB3er
bPfFtfM8zVL9tYzmb/a7Cgk/yet+KN4dsC2196mHDa+GbdgDQWQuvUCqll7bY1sQ
EcVXTU+Rd+ilq1du5mff17mWGTbmZeMXZEvEHqk05LewM5vCJASpKokbRjdiJRaP
6ItKi2gm4sAc+7YiTNDetd32RvlcKoG1t108iKIT40ggC4wCcmRxu/5mpWZGUi1i
eFWJrdZBZelrjvKeN3lBqnHK93cjXGv2L4Eri9saVNpMAYhJayvMQs4gC/mp8/Cw
wkYYAUn2S3p5luq0NJ6HeTTWpeyeT0cd2igjV/ER2mnJKLyaBpbmv+LgGHsQH/Fa
HkPsn07Ak/8//UYenUYbU+q9PxfCdiLiH0fEtx52srhDTudCjqBVeUg9nyPvLkCL
L1dOUhpsFux3NbjmvbF/Ikbcc1IF5FjbLmT0rvBY7RpHGNr7i3eODbcFQEW4/0P2
7dcm/m5WmqtmIl0rpPiU2xfqFTokTYngEcR2Pax2jtMCQ9xUVhWO+Is0y5L0t7Wx
Pc87cyPx72jxQDngY5f8wcElMpbPnIsbTWg0plKXjZzIl8RFLHv07mj5xJlrYslB
1WbtKbCLfAsnD2kKwMCdTPzaZ0gMrrIQVkdwyiYL8kCnfArVepWGLhA3pOk4Lr9O
X+XQs7xWIUOIlHQZzHAxGN9qwiTefABAQRqevPbuDI+xl875JY99cnl6646kgNyc
zHgtk8Ps8pZIq3hpf/8+mpi6UH4YkPij9oR68VieAdialbEZ2C6ZWt2e0tKQFfBP
Apx/aG7bXAlBgvrK/dqfN4klh3GGuQs9kwSKEEMFgDmH+fxCKqfHhlcRfJEGlwd0
gJGacXyYLGoIJbzhzw4SdtDJyJ7LRaJdwGHQv7S6Owc3OMi4fMN5KYCMnvAlrkkY
dblzRzzt4bPUErHHf/92ZoVnko0YiXYajE8YGipe7RkUjHf6qjQ18ecO8kgjZHEC
ILiGG9tNoVVcO/LrY1/9u8+2rfEFztf2d2Hnk4HSXhMGz2ibPTtX5sOtEt7EO+yg
Yx9CNyFQtl6yANsqRV9DbXv8ab5bqsCLXV425kX6SBAirrYYf2WBchFOOCi44TAY
qcepa0mfbyWCaF6Qxr/jJQKavmG4wRFTqiEsP4CEv7ChXSaJIX2fhlq6AhgUazo8
DfUYoTfLLSHVzWu/tbpvUW+LzKfviqlnVHviFJ8GgIoKg2a9nj4H/SIXyp4k1FHG
SJRC4L58jerwdu+M4LZ9exVCVShf9VePWjJjA80m678WX6u4bVkvLszvUehsJOZm
wmklshS1aa7CHJcPypzQfKmu74ohu344yS5pvmwiJJUSOjuDaBOU5ugm1PZVkRlX
c6RourYcHyY0D8jSZmqZywlIl45sMwO6Z410y04e9iVFvbFIWt5s9HIHnzQVXBC4
3RUauQe2866E+gsfdR00DggRUhxG/rBPOynw1Lbc516WpqimGhL39Zwmc5NYLCZ+
J3D2582kUUil5zFRcRDfzNrVcFvo7kILTyesyP8GK3DRyPfAOEPO853Rt1em0qFa
ito7ZUJ46prHw8bJpqlvHg0p3/Ht/ufEoXXuOkqlMNR1R5ZRP/salKzOnz4L8yeF
jbJ+W7f9oYOTihggyIGClWNz6CQykkfHhB+XbUKB7s2siun8/2sKORQK0B8JuZvY
h/7NvRGPSRdAgGsjJ5mS+9mM2wB9f82ysMGV/chHNFE6kDzCJf0x7GF7+/n7orb1
Ar7AXZjXA18eJTq8tifL9RW0DNi1+U2nPvoXycTg161HfFFEZjbehv6rVysVsCMs
q+iSeXsLx+fnpNmWiW+VDHmMi1GCDr+wmWUd8Uak02n0vvur4ZrAFfreg2ByDTTn
KMnS3dE9IYhONfebBHpPmuxdxjUUmEtD2ABLT+FVbzFjcMbCDCOJt0VvHsIpSRW9
jUN89FnmCUwsQxsJ4uPr0A+WP5jUcoxiQmGOIHBvxyNvgEMgw7rqdrf7bATN3cki
r2n1vJb7Ad70HQIq0HZ6z5ZlKoIxD69zrBlLu0Aukf5ikzP3UWRCJRdV/yEIqF5+
nTVOAjpHl6R/n4I4o4i+z8Sg23x9+fWiufQiSp7Tq+y7ZdgGjyFqkD02i/ApEkl9
EZRkAKInzhNEfKUnCSJILTh694/AojKK0TWWPXy7dZqXDeEphpI9J/sZKCyofral
WHaalgjiSJhCm+3XTKTyhHvxOvhFBeMvoVsbpg8zNlPkb0ye/GSK4tkP5KHwEqj2
49ov9pmX49sfjVzjX0BIjuWjxgPX2ozoEtYaVO+al2nNQsijHyRyuGoRA7dP5Pid
+m2JfsAD3Vf9i2E2Tz1X1QHqM7d/d++mw8pPlJjJOGGUMObRTW79iPpqXoABg8/u
5oCJM77Q+RYytNehyqHoGAZmJT6x3vUmi2Fpfv1UF++ZrHrAcIEliF25z7NkjIFP
V90RTEk6zmRdh3KmuTs77TNUbS9o+tnKhZ1Rk1XH1EwINtzLuXn7JxTje/3qj38N
B4bB7Vi00CWbZFUjy2ys4mVQUmeUk77EChr7vCZS7IZUIbuEACS/CGHzaB0KQ/2S
ufLNKkuSvfiRMZuKWw7hPasnGpUZLxGS+Hqb/HEtmNvbSKHLvn83n0bQTzXFBDYQ
95F21tTdcLi6bdP6KHtjanZegRQyZn41snmBxQzDzCr/4ULtEdyTY62A4aO78wSG
6c1wCBqkjbyjlFV4xvB4P77hYU+n6yegDy0NT71l0TzVprdMhjHHlFe1wBVs4GNL
EBCaX9oWbYmQorJ7Mvl9jdcFZYyWIis+/bJwvm0LLUu63c4xfOkLTX5g+wHjEoSQ
LaEoSaTbaRSeSFZYVpuqpnejTvXs47TPE7GSLeZc36GsynUq5M+O2ikyJwvbQ4jn
quIGIOejL7QuJcvg+YgnHLw83NDcvIZj/KfE76L9bzqkSRo73UMGldK+uYiGSbw4
ZSX28ZB8IcxREUegInK5ofzrGqTsSf9lh5kJrgFOCNgmBCiS5tKGPNL+Qh34H/yi
uNqm1EtgUrlyhoRDUBNrdrYMv4JYWmGZmcOUWsmG5AFcSU6W4JnN4ACRlG8PNkvf
AgJiENibtEy7xoGCkEvBkr+W0BGBISzQEAeJYKecojHfrFM9ncdtZZ0yuIzZ4H6C
K6uWbrBPp6afqAVLp5cbAFx66VP0XlBHHZgyT4yLqR/qHr4AAuRg4P/Y7O7vMQ4S
JVbo0r5d3MkqNig2Lgbz1kqi32MzKLftCC1G6lQMRVyUOvK5xDyOfFJV7pLwT64/
2SkKhuI6ojaQmZ14HyrsF5BC3k2128QkZgcItEJar+qYYrAoB7eaqq2kkvKfhFWo
rKZZyxELaPfuYsczb6ABm05X+X1O/uFBHvBIu8Zpzpn6Aa7gN3uKX1BZs9FatdLJ
kcxpTZqH5zCn9Dc7waGh4bu7r7pi21x5njdtX3GjeDm7dZQyzgub6EeK+BPrRpf3
h6IsBQL5nZEaMsXAmJ2WALHPSkr8PEmT5v6GsC7SATZvCki4xSq+UtSQFXxW7O4y
LNziM5myLtR/cpfZbqobMLXRaBJy/X2azzI/QqVOPZ7e6FeLrfZckQhO+Wda52rw
QbYsO3BpUqDfD9yThGtdIAbcFGvcJk93j138sM5Klb/kqtLyjQQk3k4Q3uwwszAw
tITc/KHbLdxghoBw15USsMAcserPGfPdoIEGzmv4nUoA4FlJbuYAkjj7uFioTuoH
PHOK/LVT1J0w5z9f03PTosSGycxaUaw+KZzwMoqL3ejFUsprMb75XzOBhf5JlTqm
9CmqXVhZcWA7vLel+Mk3loUVoLc62SP+cv/fuzTICJHTE4LPTkrGYdclFqiHWHzr
vPN0+QPU4kbwJpIwPWsQGl+yNgLHkozYWA6Z4ZHWgkIERRdDpungXEiB9pdYMhYP
d1+o+BnRQs3+84k4GobBSW2SSozkEqsFrhrSk4UZE+Dea1JJwvYgQR9JaY7duTqn
jA4l+3/EZt/MQuoH2l5/VtBd414DQ3GJCG1hX5Z7dkuImweM3ftz2U6EynbEl/7/
9/K1ymOA8uQn1Z56DOofh9q6IY+fthh/mEbli40Ya8Uc7hqRTWTflNCBPAMjN0U0
5UEXCmwBeX+cimtYJHurRQu0qdOR/Xdsxz3Ms2mXDlNq9fG5fopxnrFpVbXMYRan
HM1VR/pqtywjgOwZEK5UfIbxVhd13fVyEkKzFEDkg3OA7JxKjaU0PvD99z+xkFgP
TIVoL0zlzWuIumw13jDL4H21ycC40yDoWSLW62YAtFRL0LWZNNnOpYrtJB8pI+1+
mgXhF9+DEKFXZG6ygn8zIHM3njkGPe2Bacl4TgDBdvOD6rucK2+ckMovA/+kYVPy
TNLFp7t4ITXBtdaqn9YBHfG6vVw6eYauowJMIX0318C8Zo5nHkKa/TW/EfhVztLz
11hQJ1Bc3t1GgMfXhc0Wq2c19NVNeYgzWctg6jEGElL9ddlPBXkFcdqpjOirZmNX
6N69QSG42SaaHApD7LQk3TUiE//t8sWfDTDmWckDYVDldlEnGyXb9LQYuNec8leF
x9LF96Za+PJCzc1Znwew4kquqtwsYOVt0568X6Gc3SsKrHFHxp17lMBn790tvX0B
itpfEbW1At4eyXyVns0CsFRpJb1XEpEGcTCl9BnVAekqNYfJSMfa+wO6y2v+QLlt
OrqK6bbkn+wJbiDD9FESMbR9oHyVG+gWKwSGkmkHtOfnAk08XVTcyy5NpN3Syc8A
JUWADcnOyBYseHOOsTghBKFZwNbeCIstRVqv+3IaaNPG4YaOvs7WbangpeT2CvSG
89Ecnnd/nV3uM6rnYJcLe9xHigHIxohfQ8Z4/nfe8PMlz6d8eEFMsyKKkRmeMsmv
N4IOVlu+yrPM4MQu/++JIGkawIAsjUkHpGsbDqFo54WIhExb2gvzD/YNjwCCEDc3
0FBi1vfWuNXpjLupe9njfyRAy+BX/+skiy8kcMttOPMTgmNpehLgQbQz7zwjLf0Q
uSKIBajaLn4A69+5RpJ2OW+RinA7iwudVDmwcZOK6Celo/FSvtQl2tymh6N3MR4o
LJIDchZ+EP3WFPUcIchHMewI2/xLqgiwSDnynWuo19nB5XeBL2DIykq9JDrCUEdf
FHrSOv+hcACv4Xy8/Rj2Wzdv5gCBeRcrhMvmotVQtIhgBchhefVwFzZ9QCqH7CUf
cZPlsV1fppcc8qEQu+w4z9PwXz6L0vOGh024mqAgbpxLY3NG852Vsf73LfOVMCIX
wK9BHyVG1u4GGSkaxTpD2aKyDjVSxvsJmuTHkeRxzK3PglW8ZLs19tR+85CSXupr
3Sj8xJcJM9WxLNcYQbqVkr5ulkZof3bd5JvClfn3auV8salTZAMwxvGbRXLva57y
avcJMxAOoHvqmRFi9//utVeG57EBKaZB/Mpay6ffXF0EwTxAB3MfQoLSwsMy9xTQ
dqUG3e8DxqBVLjhl21IBQQ0Z3jKxY9kPdyDB5F7OBX6El2TY8h0qbjjgT7skP7ua
kpLYjSYVCEGhmOkCc0PjeQtq1b0+GQ7BemuKsqjd60TSiGhcs50zxCHUpiwL6/2y
/41HGcm7CXZncgBdwQPunLM5ewT5j59XPv9IVjUBS7XZGFbTFm9vtM2HHx6ORJCF
cO02QxzKHBmvp+0UybMsExVeN6lHM0/Si4bs/WyBaayEtPQiIpmLvL4w8WAwY9CK
XehfWGMXsYN/QH2CkJ61fX4mJPIjG3lSoYR81HeArNzQdz7TM/JS/ib6SKUJGoGz
k0M4XYmC9SmpfetRCDhZGtPzt3BWqTGrDWfg8A7DBL5zRZi6dcUTjcv+UqNOy3N7
mQZUTbfmwtGmPviZS0STQpu7L04Ues8eqBi+4E2EiOJkrduTWh/OsycOsL8SAutF
MpcjLUqcOkSIm3olx0BPNg2OARDi9WeV4dKUMYiWdhTfCI4iVlSKanmjYSArz/Ge
PVrtFp+Eyy9jbFMF7OxvG1X5w7xyIlc/9GxqTpcmDZ/80zMfk2V/h4ZRDSJyGwyt
7N0czu/paZkIkUo4SYPi+kRw0EJpLGTj0x2VIMQ+EeBIG/CRgGUUX8tA1jzJ0aiv
h7qP8nmFwVMIDnI4EVMvGybyaTld1bsDtgNbysBqIuX6+NpmJD8prPF6nkkm8iIp
O4JD5oB7iLsGlzb0Uzld+X3zcIYYe5qCQ/tozEp3oZ6OgVH8/8TywJzTzJRHgk0d
V+Z43AZL+GAx6qqBEEozlBh/2M2P74hxEh5AYwb/HtP8odkwQEi3xBFXQYozUa0n
vBidqQ5dgr1IrBjDK/e5yLvQwkWTLuKMxav8qDorEpAy8FjwsjC9+ZQUOa+9rrUl
YZCRAVrQ/y9T5EmpoIdb/SyRDkJQXvmTnKT7KgWhrhvlzpk9o/pqC71M/g/Fud38
/eTIF/OKPlh8bLtbfkY9sm9DDNgMK0clRi5eJ6JpsLvpN6f+3y2L7nxL6POa2tYb
a8+3oiK+8ZRVLV2CDXC1OA1Tz79fvU3+L/0NDUTEyUSKIeup4R8HOuvk9pWNr2XY
0oq3m+wCT4tdXCppHMKvL+w7WXCOvi/zl6bMcW5OedqIDzgab29sVtIZIGv0W7ht
QnwdoMeV4AYpXe+QrmiG1+jNQFhGynDtUzdGrYRaFAHD5SrKCcRgnChIBbABc2XD
eN8z5pSeOFiMQWJznfkDfyh3TJ0NdOJF/G/0E47MuOjkwXqO9RVokp7QXb6V9+X2
lzsApwH4Qqhx9QXVS+dEUillL4/ljuiRKj0B89z6z283O7kBUmt9f7RdlrBNOLtu
GuQ7m2oIA6P5MG4jJjtSCA89WofVkIlLImwVClJvOcS6lqn1aCxgjGEjDOC6D3wT
Zih/3gZKHaCjIib+Kow1kJSmMe/M7MF10tPX3lfKJOfhNbMO2nMGH3NwnJkdmR5P
p2FPjKhwTx+7LOq47/veJwwQGakU3VAw9oekIihafyApj1AOqVt9DNJUx96DnpZI
rnxH+XDSRsxZI87m1q3GEJn1rkul0m9s/HHG2OIlsCUhxR7XM7uaNbSw6VTMoxmD
ykK/tflgWojRyniGKt/NFKVKcTC7SRWtc3x5uF+x2R1T3QGC06jTd609Q1BnxIaG
BQV33Mm/xa5MsgrSGefzUomu1iw05tTG6PvmG2nF0mhnja31Rk0akE+Q4goWVHHa
hQ8J3noaP3okGesO5pecJ0eemnwmDeuaVGkJWKcu++oQiu+ti4zotyJ0qI/Lb8ib
yvwM6fvNdcJc+uqiXCx23UcVqxmAtP/vIjjL3aGOgLQ3j/isghxGhCxpB1IgXoWo
jcSRMINWiDnYu8omKQ1f8VZ0pziWoF+RGxyKTyd3VTFLyd+KDXWn2FinFeUWO0I6
Ymkf2XmS8Ck2H5AdTXy5kYpJHr/fLrxRGo/MxPozb6Rn//wra7begJMg2kTsyIkB
WylDZnPJ3eCmJYQ+vds8jRzl7MLN/gmNkO3Bye3ctWzEq4ln7E7gd2eQf9qyefM/
EEw8f3beb8RPSu5XrdkkhUEbk8HrSETHZKxraJMa2Z3OwVhl93T2qgrMZe8mNRHV
1YThssAbIriwkW7eojKEQKs5XfwdLoQRqHvlkqD/TPr2PESberZ54N5THDb7PqJH
WyKMSz7G8IWjh6u/JuZsy0hDD8UDoe3P5YBTEfaIkJkEnN3P1LCmlwflMqobl5d5
y9eEQizUvVJ/MmOVSTUBHx3hC5yu9WQkbc6/I1RPaCquAJ+e6j9KR5odmB/jjQ/b
cKx4ww2+mKZSDL0opflIVu6+cWs1U9qVvb/VCfa1y72nQEaVcrBx/eDmHouRLhso
q57xzCVmz71dkgtLRSRS6WWdOOBSFoIaWVD4lxwSpnXAyn5h/cpp4ZfUTUw8MkC1
xADAjceojKeFDXgTh4nPQCipFH9fhRTVMTyYJzhAEiP/j9sXxFpsIDInGoV4cg5R
encn4he3fOiHDSGaMQXmNGFhTVm7EiRfLUJxaK5Exyr382fKtl+ErS2+PW37+7Nv
EEzjsoSNSxrL5pBbnUafKdBm9x9FxByazQtJDMDkPhyc9JxLArf+INxX3vrgcL06
EXTcHvx7tbU8SdK6/LJNYIIE6haY81LgmagbsvweYJLqe+JLIZeRux8z4fXNdZZd
Nnv3emrQKC3TEEa/gQylRCmCY3k9ZaLialo75S9BzrFjqFUzcZYxMj9XK8OWLx+P
wP5CKMNw/PBFIISGZEYfLZ0Mpkf+6lN0r+P8ssSWYYDmhVEgE2ADLYLPPo4CmxWq
hfHNMQKLGpHhNtD0OgmXpjxqEcYHtheM3bNvrHAdDPH6l4wIH6Eb9je83+hqHZul
BM7M0nPmTyfR2FPCFHLFHUHGD4RY7flX/oGjws9f8FUphkRPxFTloQ/s9uo9HLPG
7yCkQHoKTraJBRKU7BWl2jgwDK9Vv18nfiQ6N2LDTEr7eTKrk4lxhV/RUN6lTFWv
ZezJ3f5hVIQ0YUlsApdMBLMc74zibycbAbS6wm5bqNGVjoIhRjkTbvL5QVZnrTvj
da/R+bMfCnfSp9Ojz0hS+zqBKaT3wKvB9x1bbq79Vl45jVO5AEaVtf6YHLu2pPjV
4aI9TFeYuZtpMyIHC8u0/mT0TuXu0itI8LxtRumnnLRo+SUe/DG2SmlqbZTaaDss
FjTzxkV4b1cId8o+W6apCzVctw6a9muJgeDQwRRXioUMGfmU+cKS1ahLfEyxppg2
9HVxO1JNGbxGDP+aeHgrGN+sWm7xJcY5zcojZ0agjlv8pFIouYcE0tRmEduuKzHt
0lT/a3ZEoeUxsc8yorYMYW6PzOMaiTTF/YIS+p877iR+ZpYmcFQCe+1pB41Sdq4x
fkrMzBA5BYNIOi7gQFVIunD1ZntzHs2WWdGGDZ01kkWo+miG+C87ZJjsa9VQjK7A
e8AHdzGjIYBv0cHM+2sFdiop+X2igZGFVubaFnxeGJLo4/Fj5Fp2YNhOfnhNThBz
T4bqwPylZ2SNzG4YNy+QWuui7c5ZRGCEh879uiDZt/oSnImzTFm64X6mJMe4pzQN
kCqXXRKrnaU+6O+0Ql5G3RB1NwVa/NeReyPlLwL2EmI3RfLbfSz1VkPmf8l0yBAF
Ya5NeGOMZi7N7qZkPDhAXrT6aR8NdlJ+WAzpE/Ff8vIFdMwLykjV2CxrLn4OIp8Q
n6TZ6UDK1uSmHb1Yfl2q2OoFknLeS5RbjAHZ+Z89mJTm4cebeiglAAJAGhQaFtL6
S88bSe9HD8ZBkf/jpCQzz3z5zEImDRXsdmh4sk3JB39+NtoyfpYzO6PgyP17+0hN
+p8DmP9p7bsch3brNs7hOCPdHbNo3aIWY+S19m+fhsdc26JIM7cfpbFhS7EHEJ6O
lMGD002MYGr7aBQNxg29t5Y10gkub2QkxlwdvIqQ3z2V6FVPryG+qYVnM3n7DUy/
EozqCBKWy/yDS7T23Mta/iRIj+hjrDYI0ZYIw/srd7ufiG/Wc/dr8q7s/qRB/aT+
2KF5pj+OgnqB2FQ0/QteBudgzucfm4rYnsePX0vHtb1mgtTTrj9rMM09npzXAOwH
GGLMi4Cu9PGXQpTTMVw2Fh/Bv7qhJ8G5W657bN/z2NaCQ2rmdTC2oQEPoJdZa2jK
1zBGIcBYqEXxzs8BVkOKf27aePhVUpPb0gyDWJpoVtBEDZNOjvYFQ9Rn3mEp6AVQ
7eJkd1oY359V3PMPRtnO9vDBeLYi2XJztlC5++wmpv84ISBR1OSRVWViSXFwSMB1
iKWOclgGbM89MCVeaAhpBTjvz1PIYkcZ/6E52Fl91l11XI8ErIiNT9OaG10B6DQM
CQHBCuPL83ETntvBS0Pp/yRwhkbnKdRamty2gOWHdtnCjmVDmIa+bJu95typsxke
TbrfcLLDsV4tYkTxWIugm/53MV7i2FqktFRZZQjQPAsIPDVE8LzV/Eqliv7jvZaG
SrOEaglKBv7svUo+TPKpqX/EBxyj31Sq4hbEggeGu9kkiCZTchl96TpyEYSOaXLA
Vl8AVwaGkVnl/O4kU9Gxq3316rcQcgr0NgS+KbbRaHrbSCT9yTAnA5/xqWSdHwkL
5g/MJnN/UYnttk62DaT4mhMaMvISgg3FE4ark04zKD4oLz0YjTR2RXWa8OdDLWNB
a2Lpe8cPLH/DWckAjiQe3nt+MAFBahc79nzasdjb3bLJKKZr6vOULpKjxpi9hntx
UE6wY7ZPtpHbMttw99Cnf4b8CsvOnMtO2ObQM5SK/cVKhx90IwKf1x+HN8fngW9u
xj4HD3TZQMt6iNW2clMDsaoIjxn6e9amYwHHY9T/XeUc1lHB0FBJAb4vYNayG15Q
LQBeBOk+iPc+oVRukUrYtTGvUrD6MAm44aMA2stQqYpPc5uaB51v74LJ5N+edl2N
czGMq0HvcNQDPEZTl82lNqWTPvn3uwE5vQp1PvX6KSLvY98slRsCRAsxuECInd9c
/vo7JMdezoNmWoYpvHFBverJkwE4iN7k8i1BkpCZG8X2wWoIEJcAmahZdaF1gcaE
qvj6Rbma7gvWDgf7CDW5SItOEy2y81qiQKt5moGLzRz9iN2h4g2jDI9B3QfSJ6WT
l7yE40WBhht6leZWwdqyzFNu0uaLSniIk+i7AU12MKUO6Cv1P2E+s2xP2cqygA0x
k/by9z0mGFw0QHmNYZcBDpkbXsjC71uIYEuqbmpSBGF1nyuO6G2eQ52Fv7OUW2+/
5vrh8y/KLQKf2WpicAIoahir7GabOWFkPC5FtbrTLqpcMf241Hi/+zSGfegXNkvF
Msziudmw3O8TzNnaWoJAeVzbJwWkqA40QPm26G5U3lfrc8UBjtPBZrZLnYvNLW/y
gjlH9CFCGTMNX+syV0xkEk3ygWGrptu6xYLsDuFCNXneF9evaVp8Vx3shoeX3jMi
r8+UC7qrRcG8Gq5K6d7WPvqnPxad01yp/mobiZUJiWMvW3kERK3hfTkYDd75FSky
FhD22rKlGVUgY1EDoprJE3580ay3eO9TrYF2jo4yDgaixtgUT1CyMVfDiQZwptDq
T8BXsC1pQOM8/WSXSPB8vCmDRHmdga30pUlMY9A1jak8E96cZDsGK6if4mrXHvkh
Pi4alDywnJmBF2nHEFWz2gJxgJXScsSUGs3WdnhuWHaUui4YSKxq0yFW28vwJ/qT
oTQ6AyeHKVxoAobUcSS8ETEfwqe9TNjQ2w/3wCDR1JcNVW96Ax+Sfm/sKbH+Fyzc
enfyxIgOltTqLbIK+vU3wxQg/ug+bRFc5CCQVjRy9wfhqpEsKePxyVdo2lhvWmfs
uuFWfyCr/CpKB0N4WdvyUlOQOWRKMUkDXVE5XRLidpLIW9LrdKeYVVhCDrIC8sPi
ty2lv6rhpWf5//Da5s8PfmQz+VFdWMhqe+HHP7qu0y/WQgWb8NEQ2ZZBJjeFSMXe
I96kwN2QYk/VSB8WUDxxECdoY+1gj4uGqAWDQ5dUZ3/4MOmG9VenSwev1sKHa2SW
mMFMmApF3pJ8DThC3DAp8dzVRpKqSh5wmwce5JkgmDuKCbA9vGCinhNylmHlT1HT
XzvRHPhJt/hC+qyl5jsDb9S2yoEgBIathv7co/8LtPL/O8lI4g9bJDMlRZAHhSyR
j5CPwEeC8WgVhVyIgniIudUzPkjjKW9HdNaVPYyyUC3Xd9OfC6TOIFiQ+J/krthJ
SEUbXFc8Pj44D3Bju7/AdWWRxLYvgAZhD3nO+I5NpGfgrR3bqvLMiwJN19/dscfY
b8hCRzRo9t2VM8w5UVOqsYcLjnMr7EUgaAxMWM5O5VnY2i5wzkIgSwfmNGsZFZ4q
o8kif5ScgJg2i1MzLP4Fjt3/GnkMNBII1PcHduf0DDWVLE6WIsUWPGEn2xr8tW+O
ZfghFOzzkCFVhDlZB87oJH0S89GGjsyj7RvbczlbSuev2GERmytAuFh1XsVWcAN8
hy10IgRceBfYD7fx641bCsL5gjDWrp1SgTIDFIxaAALjB/NAGdaPx7EQfWHLlnCi
u8W1NqP1NLpwoEcvIsnc32WpGQQmX+rK7CwPxLVEcIxCbFUrPR1boDAspW8Fd4Wy
s/B1KaLhyHvDawisa38ut4Atu/vVU69PhnBppRzgnYyaxkl/7vfVCV1QpgkIM3Aw
DnoxF5phul1WRDwgMyGi4nGi35uKDG24QdEA9UDD7kOSpWkPT+V1U8PfqZ9trLZZ
xTNYqZID5csQCOmTjIU0SNQuOb1EVtdrAp3sr+iHa58VTol27rUsSfftDwstNu7R
lyy+/Mw1B+4xBJPzqAIDmyKol3SccZX4Hs/BdpLmGC+sWArVldFVMFUjbCLNaJm3
0NS2NQ+fgRKPM1XcDN2iOiY+MFghHqmA9VT8pG/LYyYoFtDuua/tA8F/P7kcf5rn
xrqq6fGjq483fHV5eCRI6xYOVSwa6hp6oduhMr2BtXKdUgNM3r3Jx3c1Um8sFN7t
f0GX7b0cjMEn1nGDPmWmNsbCcKxyQoOyE/5ssuNipUawlMahe81Z7feg5m8bt8BC
nosuMDaU0rx2x4XiBxEPHfZ4h7YXWihBUYeGnGHaSoEW7End5gK0rXMGcjw0UIrI
UtrJBE0enwTIbq4Gu0i4zhHra2TkguO03fPXO5DR1sN6doXv9f/RXFqmQ+1raUoX
t13RivqgTs56m8ca2z6nxczwd1zcjJXeYw85L4bMMh6W46svokFlGBkx/WLszxJo
uozl+u7f+zqd3wvKtq261R4zWAof3YnJrPes2ul+lT652sYXRtuTRX1USwodL5tR
BXI6MmI8wjTiqd72SJ5gwPedog5/7qh9tsCr2y8f8EcUIKrXOrTKzoj24tTwaPfz
Z7tVQDSYAvOocw0DPgg4UipBUW0htD4bahUcy7XwtEsYeBzose1YbMEjGvdc9AaQ
UC5+2mvzv18Sc6JEjoDu/4g6Dk3EOFHw5LCtzTy6wUS0gegnLRmjXbDdTb+ErNVf
bomUitDCMPpvkMNdWBf6I5yjkmM3w8ANUn8fM2tdHY8g4sYAUHDJc/2tX9jeDf+u
Luz1JHv+M0AuVrkO7t3gBQX13xNlCTqIVapGdwI6pS1sY4MurGxu4wADyA0faPTX
m2qjdMJ8hTqTWbvaR9VR+zB3rH7Qy8CCwz9CG1vblVUOC+Er1C8ZztF4X9nIYDOU
nB1UbfVVb2+BD4ViDIui6E2E/9XEt1XXfby3kZlG0eWG/pHxHOpOH3cY3prB0j3G
bMaSvwgMYY+yb5hC6LutU5Mt00oV3/wQoiLdXOIPRTLH9Jjvk57sg0iuT7rbiuLC
ASgrLci1dRItB8QpxvrHlPxK+IYrHswuDPz3D6yVq2RH+lHR0R/d88+xxDJ4EXKP
wOJufxn2f/tf7vO39ffOCQbKTQ3EIKoFMk24r/9S722zKVlj6oSqziI4dupJJY57
Qu8USCJ+5HmcscVt8oBIybQaL9DMCAR7tikAy2nuBTG48JP6Ur6JyRml17qGgm/i
NUgkryqnNA43evYqCU1P+3tSqXhImkk+flXDEDkGtNUoNlbz8T5N9m4JRDl99hOO
k9TQ/dHy2eP+bszsEq23gS5SbWANdPHC+00nRNKO+E2Xuwfump73FAxBSAIoZTrW
IyqQfik64AivsVXDXFOEIrUtF0sBXSkG1J8xEnZKuJ3p+Z2oJrWmEACrbEw8T+zO
olkIIjUkcpKJQi4eNCg33Yw+4L0QqwRElKOJEDn4b1nFD5820ge4NMhy5JiXltmu
Hf84w3zfGvNhzBaI4zXAdsjPPoI1HfDFrYNHnlNKTBkA2T9CUn25gVR3OlECYIc9
9J//o+JhSnCWWJQEQ0hrlWe70XZAy/tphGyVZw2u0BLjmmdwAu8cAvOA2TukpsLs
mrCmjjJgSCQaKIwVNBE8IXv+dzDEF05BWy2Yj93oBud78ScUxbrAIDYsKIJotWf3
EooWr4YGyj+ahMFQsaXbXS+m+YaYZKFBxjNCRhy5f7Jf3skQ5BnR6jdrGhtKAofT
4r3EPXrNi4mw40L3z8g5bULnCUZ1tDWXmulDsNMusCFMDAlpXvR/6wEShqrkLrfB
iTid7Z5V8d9jMewaG2wPpynVGu+CBRGN2Fs3FCDsvdOuiFu4SXv199jJXZP0aIMr
NMy/pIktA0i1o0oiIBFwH7193uXdfh1tzZcecWOxsLiGr/GdYhfY8dz0SoMUQKUg
Ilg+g77m1dHLIET2GPboPCrVwMmEnHGS/Jf0Klk6aouWgJ0lCpRXb2vGv+ZePeI7
B/UR4CejQga3xE/dsmpdsI2qkmEn8vTGS2EnN1EUQBTY42ZOXzQIBrYVf4vltnDe
/osqf2qC2nwglC0q+j04BCGwwuItBJ7nEbsnKGSsqeZ2v5Z6p9mzvMHg2Fi8FgPH
XFzjx0G+io/kMZCSOlEb52RTC8upS7eWa2CMC5rcKKlcvBLJpSnfhiFDbMj9Tt2h
9JwaJmfgn/PagCdYEjLkHwzS3f+zlzsQHbDs8BqcMqvAYqsggVEk812KIjCkAGsQ
VuK7pM3kpoQcKl3n/8XKxcJDpWzIZELJJ0AnRySJ6dtqL8aOdOSpPnExd9MlPz5R
niGeCFF+YveJvJ2VPn+YVYZviYf2UJIOcEAqj7zZOc3CDAUtYtxM2EfSflk0i61e
5gAeyavfjntnL/ZztbUpAOKVs+JBuMp7QViTeiIgDYXbs7slfwP9R09faVfjjgSQ
LLDUl9KZJgAK5b2sKPbKcqF3sqvkXAw7yLbIFMTIGuym6qhsZYCwTBQNi0rp2+Oo
aLOQzRboV3dRSpqwN6uaXGMB7c3ILaoNOdzwZErO3S07oqjOjSDSgYYqO3zOlq/C
rnHiS6gPtYt0wkQSN4QMXP9cxsmVRxnJTT74aC+l/PqmTcRKXJ3Cs8B1wg+674sW
c5maEaXF6V0y5ztrbKsRUmmq2r0pISikHeIFNwfzMT1KfY/DjdrPH+ZBMQvHf772
ihu7/jYK9o7tGaEnYxJdO4z+blJjYnO/X1bGjoXSc9yDXweLf286V8sedKXPQ8hb
iwOpstoxQHlqfyzJs99S55OpbtXNxkWvh4rPEgNSRbDe9uRvDQbMBrPVekPR19sv
GO/u70jI/VJCSIUhPEFdtNqDVY+/y0Z6FqBdyQnowniR2VqUfBWX0FB+Pfv8dEXk
1Ps+aP9PhvXNWQqpbRxgamm69CQziKJLgGVGpIX4+ktcl6EVnMCLZ8xUIaSsxeK2
cI3FahflD9G95G4OtTCEyaQQ3RMdLgYyPxYBcJuL8dFV8a+K17Q0cip0fO2l8SKH
hiNXedQqlnxPRVlYcqW0sVu2YXCI1Msk5Idc3S89oSzJx89QXMDFeaV7s6sRybNx
+g2rx/KexU5O3FPKWquT4x1geayPSvK67CDA2ROz44fOwB1xmS98dd7aG/VgYbRi
cNTvXrS1xf9a2NptLqSeY1a4zptwjA+dfTXwvMkvejn8SpgfndgqBOK6qG1P3NZl
2bwhHtVpIu7f3UrSVvBMFpztTbXCbJdHQvB7+q4tJkCGsEO578ue6snxuntyv6bl
KGp5KOSaucrioGWlJbwosuGa+sZ/sJqg5NJ7B83ImQ2wdzovqJEwYADlsxir1Brs
gWUHwfBYw6rslyABkmYeTWPy2sOouvFPn07rcudSBTSM7NO3GyelXzr6cHSnOP1y
KxkUEmIt1uEddZrMbwKUIxB/6hF/ximn1Irs2ULC7Ykm4BbxGRrviCxe87f1sCBE
ORQtKIrBjnC5pEjz/RxN8jL+aAbRDyu+aE2rm+35nadrIXAhfyOZFIZRxWPpg/Dd
otu3ZD00xxcEMfXPiWT2s8cofquU1kT2XYnXIoVoJ3bm/6GMS+4KMfEnGIF61bvo
FDO7mzOGpDPfYxEArxVEjj+ArOMPYzTG1aD0uDlyLnJoiuI5xZKYQMTZGmxOxBut
+g5D8FriVwdYXwGphc/mkch1p6breHS/wHVyCkrh8NUhAqxoNooRB9zqQ+gpCH/X
C49Ng5rzG6BKnUXiQLh4O5ETJLV94UnowI8OmQVn1w75GS+jIISgq7r3ScIdCPAj
g02xr+EK3vEaGseecyKOCQaEGXxNoskRhRRlR9tqK9Bt3QKVp7lHU416gREvJMQH
LRuGh7KGIFn9qZNNkdLrKDL9j5dPQHq+s8+uig7SLqTNTl4rfC5SAxyXTqn/x9zj
jVQletunlEYMToWAAp2hw8ZRiJu6jnKHrC+3Qda7frMCJeQRgxxkjPS8z52InFlj
/VFXmAMAqkUbG37I8fb11Vq+oYH4TU4NEMZJ+SeXZmgbZr7B6w2FvX0wpmNfZE2x
sUnBjHEa8OgYnSGGSnJHuGGt22GxBnZZOKBno4F0XOhp5fsEEmJAz8uWKYAaWQnp
5rzqTsaruiqkMzuRxXTQsBLd83Vq5oQM8wzX/S/2+8VcdPaz3AtwZlhHHo1gAGfX
bdiDduqoaqX2eopJHwzIg+5+VkarOG7/R5WgNN0joegZ79qeFOBMyqA96+Gbpk20
fS9MsL4EgoTyyNwc4JKQ9W+9x7lTdY8lRxqG9uYr3ij0lvLYKHAMnOL7LiKBrAva
7xUikOsUq8ZBTRIvHufiqt9TbKD4390PtaLr9LdGLzIkYZ6D4n1AVnprLPtxJCVe
d0qnYn2DNI5ohB9R6GXzFaWt5Gdt+7xLdiOQCMIP8Yrfq0qD7BnHBjEgCzGTXlcd
i3O6yVCLQsMqJPUs4rED1DYhq27s4WTreiZc3XjB0j4jyjdOXkdnPS1Dt6b/xDiO
AbJYuZC3dPyUgzJaIB7C5LV7hm1t0RljzH9GCLpb4SQGEZs4kceSVnigrxbfSrm1
a0EVTTYyvHtLs/4i9hMlwgQpGQjd0N4hCN/xHWS202gTgxbQlCtjbwU3tgdRYd+6
XJaaDFvASBAPX18YmfpK0KuzpybQedrNhZ3jIhRUB/Rquz2OVefy3RCrQ1qy+rNz
EQoo9pSLJEiETbFL+MUsjtvc7Er7B3L7Dbji/MQVa59IEcLtmO1g8TS2/5ZOUDjL
/qOyl97F+90xye7TaOJtGZgb2xK99xUe1a/lyBvlW8qHKqnSy2MsyvWIBeMIkoBe
I3MUUNwG9UB0IwzoVR5mQeU6XRW5mywA5rRR2S/L44bkfcsg2zvdFrUx5nDZnYlf
EILjrX208Hg0Pm3+yUkeM4lPZCUaisEaqWoJ2PdwXFqYf2s7iAG1GwpIdzmEY/bc
eixchkNbqPFtFpX0JBM5RMp3V4VaOy5lqpDXdU7bJaC06fxJaIxtl4cTuXcPlhkL
WhvCyG1pLn907zL/jJp+4yXfYDiwGdRs7ZIvH67j2TYoF5O5Qt5i5QY29Rki88R9
BNA+w+v33kd8oq06RGJ9hXDeHB6H4f+/CMkcjW7g1OusjEmspg657tU38NbWCj2h
YteYpFiNttUXZDGszlKMCaZWOiaqi/LK5+QDQq+6aoDFbwxH6AVS/P+NjXbd2NH3
dOBEaQLUJY3Nb0+iqdvsMIIIHSJ+MoDxUPefA8YdHTB6vRXl06mnpJxOr8O5BphW
q7687yxcSG3TEvQ1N5dka70hufeNLLCgclAptyeh1uhzF3Q8kvQATHWrx6maVmYQ
oZ3j567FssIhTHQC+cO4jWWyG0p6ygE+91hwx0d22d7Uf29P2mgip8IFov7WsS9l
+DvLva/x6aXEq1na+FYmbuiTNAHYOZCa7NmrjKjdvPTRhgIOEfFcML28+qmK7rrm
9R7Ze0q7SYInkj859VeVt+BFgdeex3oZVfkq5pOK7XBC06zFHJyfjNBceyNgpDTZ
0Sz4FTB/WgLWLGv7B7i8YKyLGW7tOkOndjvKeOvuCaaXw6beu8MFqEHVtrNjltMR
ohNv25nEHALSLgda1UyeRIyIH1WpewKpMnVWYc393cLh/sZ1Mne/eiPeO+JLFTU5
4c+R8jC9jBUIlY6ebWBGsO20uGooHvu3OwiVaGIKYljpVx+ASCx2ggWSlqmPDmtC
tPZiqAiT9gwIULgh6w8Dz3d33ZTcXfn4nuax+Em+0mqRANopV6LQbAtHax2dbhVJ
9tEtb6Cbd+SBcR5HYKqqgKWWozJzdMxj2f5ue4WgSfLxSiX2BE9+Py2/yxauMUyC
7bepMoc8rzTUg2y0l0m6Zga2hHNiosaLgFeTDi479ukAEvhefuPu+1BFezlVZGSN
PX57SuLtedWWPVHUsZGt2dZlSu5/Yk+7aDbY7D3kaZztc7464DwjVVz/8BAWuuKG
VxekV56ykBlMkzWvqQPTx3Nh7j+nN8WV7COkuQ04h1k69yinEHq+NzPl+/bN0flj
9xbz8szgg/iG6tRzKphUOrxAWt/9jNr7jW2wlQSuvO4+ONpgRMJF7Y+EolkYWcwm
nWyAJWXfBA8WmAfsGXDo+ZeDS9XWkrGqufIcWeKcnrvxlE0PO3Z3tiewNqlubgwB
QXNSiZfIvKDXMczDmSM5q+pRE66xUG6FAqWeBGD+v13sGywpyX+004ADclm3Jvur
fjXcu2WjHSg+PTu7+dUiTb+nQhug91/qNoNAbJppizcIXO9u1b0YFBp7sy2SX2i9
LtagG7lA1GPvgPNsArvHIJA1zRCRCUNBNwEfHjRAlMtbOhbGAIob5MY7ViJvJe6N
GNkoupthYh3Kj+4R26m0X16MxFtXTyzWsyXyPPdbMeIVwJAr14lK6lY3Fhqu6prh
52PrmFv8LkdHIFudFD3sRfjiO92k/ROKDUVc2iSthweNiqqQwG7w+/Epj/6Vcq9v
JJT2YD/lkS4cCJC/jkEuMRZoP0Vlb3OfwFPc5f+Enz4G0PJ8cy/rL+4mLbCi51w6
14h/upY+MRCU+coXB4eLUby3YLcIQTdSJ3HuYBVGOmWBTnP10ReryCK1nv5J9nQD
7gfsepC/aO4zj0FxSoyu442CfqiP31G6hK1rOfCuOPAghp8QwvUAtA+TdKqbRqom
PcCAelfTmmJou076foOkU+OYCo0p8s+sLiOmPqUkVvmDLGrneuHjEps8R4ppoYgZ
Nz3W14UNSRhc3x6nrWe8nJ5N0Iv6ZJmnSuLUsTI4OQax0Xgl6IDcUTQklX3gKN0a
j+X2BySMRoVbgckf6Je+81BpBzo+4pDufla/ZAYMXAy4ojmzLBl/emHRFJJyqkI8
1ASTKkYmD4a598GM6UEvXJJ3jzj1CcqzvvKHhvcWf4URmIUwQ3XMDzLYOJ/vIMNm
IhBhtJqRX9chb/qS2vLZEjfD6Lig9mzGGHQjBlqxZO5G6qnOmzcScTRGqNxsP1FX
VrPgbDj14c5C3jw4nqxm3Gx1OwlpFgfkyUWK3uQBgv+7kSdc/u/Bhy/Hn0BfIHmF
ZAmNGN0A4nNwBGKBMv6mTifxCtZkVZwOpuewpDaCgLBbUWDHLfvAseX4vvER9g5u
74HlgzpYIxwj9mZIrZdhZ3p/dRm7xSmImCGXNz5+Xf1TGkFvBi2jwRz+zgNry8DQ
IqeGA8Plj5tdp/7Rj5EKpq5feeOL9OqRmbQb8svz1WsRa/rR91EbbGwRad7GZLQD
nAEdI+YqP9Ks3mnokiCuG1s1PMZd0EcGuIOi2sAyp0yevkYH6hH+Q2BcfKEQYD9J
J3AwVykxE8855LJuAn4PndvnR+NCSg7/O7LrBIE5Vs0kpHI845qnZIEv+PIjtOCa
FnBc2LUvSuXqdRk5whO5WysU8nCuEmcGL2D8kHl2kucTTWPVixSFpJkc6SJm0Ysg
uN65YCImjjXOD+Wu5LQBH/95iyyBm6bpOjZqcHIZIdJgdOt/JCdRIRFnXpyB2Ohg
Av2U/G1s4jkncfAGgHdB9DvN9eenIOk+AME0ZLIW7wRZse2UIPmBpB97H+d+XP7E
ECQL50wDIi3KBm+luz0hwrYPhOO7gkSiyCHZIWN5xOLhBIRpEmuhHdyGu1F7ZwmL
TpPNQO32DfrqbQE92eE1tvpk0hX+kkp1ocLEjv4SUyvpv46Qclkg2YXEWVOmGLO0
hQktiAXVP/Nzn7hl316XsEpq12KSf5bMKwSBBWY7usOsUxoa6Hshmd1gVbKMVgqS
ZaBpquOGzBpr0EXnwwNJtXnNlIem0em+CCo3iOPF9OHFfu3g/2PpS+ubOG3X7J6K
PB25Wg5Oqg6ZDxnf8jB+sV/KAMtsPf1v4x0t7RhmYyZsRbtUxRuzkUXPyj2NxTn9
cBlIuaggQgMSD8YYyRBYjxqTBbTWGmGkQ3bpLluKP2Bfhbk2mbx524Ixg52qa4oL
ZvbO/i0Q6M1q8Zs/OQpn0LittYX1A2eS/TLzdEqxm+WSpb2cpgQDCH1keUO2Qnfc
U5CJBiXu/EMI3aqLELBRrOYyWhrI7bbivSGI1+bBaWv1MZpE2JE3ohPBdB3OoxJy
hUmzPXRqAl+dSZwkGBZgNZfi3EMBd3uhyaLtpRPWeCfnMdRNQZLhXB8R5Vl9sB3i
UMkoVC2t95TorMHS+Rmebxo6+N4Le5Sbiy9xws8UXuofxmiCWqaWZEbrP9F/49Mo
HPqLVebtQqod0HaFDSCPKIjLFLeIjp+h6GCd8MVXn45GnKhqcwfKP6DLtKoP1XVi
/h46b2Q5EoapQJ41XC5IMxjxitJHr8vbtFdUADxCV73Uyl9IFNnT8bbmqDC0zrzw
PgEvWnom6alv9obWXUxuLL7AViIdHP2PLD5IVVEjN3SbgUuVzKGi6kxFtjnC58jC
wgE25ZLRF4LUVY+lTxMcThxMDfqm6cuTCbus7s8EmoFJrrv/mdqIkKRrWmemK+P/
vCtDmka/W7iEPJ60CPHCI3c68+c5fbPIWtwrGxgGNBgY4Q/HnkGgMLWvTsflDTZh
trH+tVmVNfFdgSEdFA/G3VsgOBh9YopIeERicfaYIRlcxGJQk0R/TmfXYgsi+U4W
PMG4+k94xU4hFziX5NYLCwOQGI3vpPTew8lmXmGWWJlxn+eKM1uDuuqKOkS4Jqkv
XV76zQF6XVFHPKMIJWoI0Mh3GuVT5zhSVz1k2DC6+la7kc9UwrBbCAKRXj40w6N4
6kloSM6y4hpHLY31fwyGSaJaqnJhS/hHPaO4BO2nTMmohZbitoUmSYcJT1ihejaO
oi9PrOTxJEO8kuCLZ88ZXa1LVJRMYGaopvdkYGeCXILFYSQhL7igAOkhuf30AuVR
l/CiV+e5WlSR0HvjqIMOnWWyRgxQU2lGkgFKubwqs9qJ5YoOUEkRaY2wxBy0ThOs
RHn93rwqD+asWuAb8DoNXcqbs/cymbOnh2LGeP67BSAOrinrc39YaEt/OMeUGyWd
8GKuGChlgwrHpKP2omb4jbTSN+BG6YLWM3KtnN1ItePssGJLiQORacfdmJ6oMcwv
Fi/j3YTACajtmBeFq/kHMKATQmcYJdUEXHJz0OXb9Mi8Q64LVn6i7IkW7r3RbxnE
0/jqNMAkr2qJk5kwq+FkxCMTTgDcwqsKhdYN5ZZb2oeMDYoMv2oDL2f3PnZ+zH4n
cpN5GgDtMnDlz1jJYkuHcntgX8Nsd+ys5Y8lWowd/pRnwjEVD88+G9ysb837x9/s
LWIRMO0M+8g4cgNWwe7Sz6QOcksCZmZtLrEjYS27NB2LW0DG0UDc9KDpFkHbUA03
5ihJPScwHor1J5LljAH+VYyGgPvzzVt0ielFXR2jIXAuatd3or+uZ7mKcGsMn8/6
PKHIieLqii84aSjLZrhrPw/JeSF1fp6iiZpKNWsVZHqcJRTzKEUYPNgExoqhtqrY
F7XYSHp4MXprMzuRwlCZxB05Mer0ByD+WMTFZXVE0vdpOqrTjFoeGBGqA1s9DU+v
I4K5O0YnxdVI1Q+EIgJXJ/ilzruXflFoFu7k4QEwF4V+9b8QmkFJXdCy0zKv73/1
9669NweW/pkjQw4DcQ5K/w1sRXf4Pl0ImD3RGaBjEyy+LVvHt6lp2cppSE2RXwd9
yvkjQMPpa2h+p+Px1rqJkzwH/attjJVfckkgnbhn8soCSxfBtFywTiLuhvxmCz5J
8XJ6W54r4efuaMZDGy62unDabj0IZRc05402XBaesAS0dbkhhxuywdFc10LmOPPu
sssKChv6d+mZNo/IUco61W9Ad1N4s8T25iE0y2J8xnEoxaWhJ366cq3CCDGmGvBR
bofAoplpFVdGCC3RXUfVPqkssEpebxT/1nGXwIbH6Wyo8y+rPbU6BM7NHULzfFOG
nzxlRqGRAQmmoMMK3P9hhOztOT8rG2vs/ldS6E2fqiPgjM7v77UUmku+6mmFyvSP
9W57+6eYcZYJ4/F7/7ptA+AxjUZ393yuVff1ebu86qBH+w+7mVtds1IU7NWXUx8m
0dCXx4zShzzTdtW0jn5Kv7Vm5uhhEfo1i3WGMQViHUb2mQ65oTdf19AljJ75uZtQ
ioA0U2002K92JAMPNEtEIV589goFKhz9eoXgLKNrtkP9KicMwlEmXuUdtI6Gh8TI
7+cYDPEXZILSmYfNa0SQavG7LOE3j0Ul3ENrB7jQVQOJoRYiVwwP5u1QPLrYgTw8
lRJqbQ467xDUnNTNt73ksJn/RvIL9LUBFIWyEIfI/KxREOoMscol4LFgG529o4hO
5K+A6dM4cke5R8N3kyKpyqnuBXci89gKcnXRpwWlmYRhmvNHhgSFHEUnbf9g3la6
p6g+S0VDRlvofnc1Xw3s3S2NT0AmoooZZXCjguD9bneqy9frn93JfyWpppFhfcvh
B880kz+/+0Gd3rkGnvrOkalqE3qPpG3MCLjUyKgkcf7HooWnzIZt76ySgRpeGjt9
55zpBUO2ufLCyc+VamrhoWoUO/8kcWciXVF6MOP+Qzu/NiOeF0qhRflGVMnJBx8H
deWSQf5Uas17MCqyw19q2ZH8v5PMJkM+b9cQavXzkbFAHuTrgqwMcqap4oReIsa3
dcwqpeTO2mv9QA6QTrT2WZx5dDjn3NJQG1iTlytUmHJH4/hdA01oczX+zz925cU0
XMyXiKwR2LEyIfChaZ8+9JJqKgn5EBiwknbbqUxrqC0OaTgjLoFWs9thzOjS5lhh
5WcGuwjzeds+Taai4wzKCSZYaqDD2bVzYlOmd3IUwY5Wsm6eiuTwYS7c9z40Q1Yz
Cju7gkkpz0qof32cIEA9CmD1ZiUH7Ln3qFhfztCiEbCKp1VFIyVSRJXitsu0T9wc
PCCIizd2ka1T3Ot3GannkG/TaFTbtv871lvj4tzwq1QlGiP23K/Ols9Cmlu8UhXJ
G7MMY4aEB/e0ywWJGK3SeGhcI/u7qJLC3h8EsNK4QcWf7UcogV85PiGvzjJHi2pf
wjFq07BXYR2aCjsnfjVERYriJYlbq5Wwy9mqseYIfmtP5SfK+fqQkC9eYr9JZuk2
ZBET/AeFChC5Tns+qG+DOMKEWHWttSD06w5mXlk37kYu+boJQJ0bVhnpPURkmWjA
XvRuxh9VjqG529p8M1t8mo20WYHXt9hThSyBmNGnA/2pafQtyIQZ2WN/8ys9haI3
C0vkYK+ii00bI7AiZwEmQP16qhr/Es9cjvZSHafg17LIQj1Gl+27PxafWZQ9b2S4
dT9Ca7aiIGhrCp0Kmg7ZTRVFWHS8r1/gzcRMzPdK61XEtIix3dTDox1rqjPHhRcp
5e0RdTlooeuRTod5+G+2aSYLJv25X0vGMV1gBVy3QYayJW0sgHJbAMJ0Bafe28Qg
DZ1aZYHZ6rBENERf+I0Zgxlw8H3WhvGM7s3gt3u3KmvvwpuZ9+HLtbrIxbGjNVFS
tQrZSO2DCoU5iDlrUFb+QwUMO4MYTDaCGuoCaQOaDEjTdtRRs1lZGwgt/bpYp9mS
YIWfBEZdc6mkw+yxi/Mp2k8+ssxlzyXovG2IPbUIkqXXRSx9CrhsT2CiCI1QdDU0
dkc/DuCkJidQY7r8I4gCoCNjHbOuTHsvXeKmSmohJcX2sZGItrJEoTR8WTT0Vn9C
sGaDHIf25oCzUhPeSxYpmAXN/LWewowiuJ7s59VKQsK5ohbUOTmmj7opgmX6p+XO
6nbHonjTCqhA0UeHCzirhtvJT9GAzo90nhYvHhZYAaB6GlLA+gBBm3fV+075uiye
gbRJYJejgtKwDs24vE+rrFzxmZP7cOjr9IHdjBKHcJBdnC3YcwFzxsMdXLN5sH8Z
+54OY9FYRM3lCcipd91DebjDXWTbASK2cLpSIFHc02CcxUsX2TmNhOe/QT9LbcJb
q7RgTorieT6Y3vs7pdbuAclhlCuG2hLMyM5rFMSP9cfgxXzhimZLR+pLFDphidLc
Eq+mEFtlDA4dX3aedC3ML+dP9PYsBbUVKbxWdKgRWhZSJ4H++RA2XTNIRgpC+rph
FzCZUco0YkeSnvixcAvQgog2Ty5HyPm7h8EdDMh3PG6hg2JvxYP5kw3wBz3sG8t7
F6eF+gP9qy+N4j0335mQuf48byP5yV74HOjygZBnekLi4gLcI8MXgI7qan4qd8Rk
g1+DIKpO6yemOLYP2rpLmXDFXX5ldw6fipg3YoQe9O03gCAmqfYJ1pjTtWg0yHFN
jlJPHiREs5OpmCs/67EFO4z1rQ07JbCUdveG65RoXGYCGEGJJmk/VrLTWxwPfTsm
YAuqwwLehJu2L/iTbtmyRDRpMItyT6boAGU3qCHIeQmQbkjVrgnG22N/X/BAsKeu
JLG525dP62WsTSHNcXdqRSYuEdprRLS3bv2dxNTLS4lCPjZDBisDYN5vieJsw1Km
JpIG9cIT9t92gkPDFQ0IkgFgKg7eo7o27pM8NsXYZYUUoVEyQT389Xrt4BiLkkRo
ay7qhMLDMx9xopbbmxpXFFhE+crnNIwO782EHwxtvX8IaRXNTu9DKCfkA3Qu1Y0z
J395SRVJDhT8+Z3iB1VaFTDc/+jlqZc3FWTVnUbYyzRtNsAZCJwLRQnObIwrepUI
zcLXlWe6yjVcg7H+eUFQALbxfjh47Feez8WiKvcDl0ZTRG3YEC5IXoELud9tp1AK
AWEUD+tUh9CDVNsw+MZKI5lBg7/ZzNuQF+G2EVgy7sfi2hw/B/1vc0/ItQRYwV0k
wdHlCzXyMtr8125ATdLyW+ibXOQfE3MDKk0K40P7it3yVMDmkmqf7622LTgoI+vR
axKvEGDIkE9Gd0Q1ltHYkL79RWM8X5U6sE4vtrThFa2ee86BGOcxHH7Oik1IIjUq
2bRKiysjx+aVNVMUrAEL3HyLkHCS5PPdISZAC/dfQfB32PzeXlJWw+UdJWw0V31W
46LwpNhJiZvd0K34kHm0qlNGPuAs3BrrWzOeC71D7X7ZWClsZvIf0xEQvaTbrRFJ
PPZrrieD0Nc6tOHPHTi4dOqat/xYbqgyF4g8azVZEExjlm8HOSkd0e+GzwIbaYp2
lmtkkT9WlBIMxp+2lw/ELNbNA7Ev11sZbCurzBG6e0hIGWYGLzesXN8Bj0qseYRA
LHYx2NhiGTobD4JVIlhQRrKdbFmnoxB4nUGJ/HuUwv78HUQUG9qnE/33JGJl68zz
g0Xdx4POOSirfcXkDW/WTIdHby8XgromxQC8vyKiZ7ImgQJxmSvwv7h+71btvXFo
Twjf7aPHnDYKgmNo9Szkxwc8TQORbVfuJVch6yLUvEbHkrSpzSgLKxxIZbjkCdyL
XXTVx0nn2fwP9shRDi1T+FC/QP7QYZo+m61qRAH1IiNTXyjrxBO6kBx/uzr1mXJH
mQuwphwJ+9wVlDnQRmc5QKOBPgml+r+MlXQEjBmiA42XyiSOVRQPaGi6tmo8mxas
ynyxUuUgXoS7CnXzyuz/4Y6zZvcmp4GmtOYRZXWGm3KP6VjDfFHB8PNNtj+QkQwS
iW+1W+Ix20QPnIkqk9ZRZGqh1HJL1T4/iDP6XJ/OX7CCe/GJxXPEf6zKchix75tg
bTeN9MC9zo6OqTorkFYrZ8Ye4BRqO6LdBryWsi6kUl0kmPNWd25jEt/qCHHRAlrp
3aJnjH3iznF2S/mqWHL6MrB75vrK7eAUZMCp8xUTO9HsCXPyIgYdcAZW8tJhl4E/
jEss73SjSQLH26siWk7ZWPyTQwoNlT2zbG5rlOC7XN3PeUg40QFFY608zXl7/KI5
k1fu5CVGqbViueMuDFctKietruK9VuBK+1ou3qU/v8awyphBDGMfcqtV9qJoAS97
P3WhhxSlM7JqhufYbsRY/hX6IdXPFbmyUbLiRuX2FCm2ntwAru4qFVQPCh0b2+Dq
zyGrPDvI/8RhNX52yAUaSXaLVa52zdkwWhgvmYOrEHAhfTRm5UKtfKO+VwWSv3T7
fGbjA6yilik5PuBGN66/jQCF0tMQed+t0ThT7TSceeT/DQL7ns8OVzQ9/kJm+0K3
CdmXeQjO83WUV16eGZJgvUuQ+z1NIByPB707IVjVV8IPyQEjgsK47oWfs4eZpkg0
0Gm5+yVzpepBTLkbcs42Q0ltdfgFZ5Nqx56Gnugl7vHASgHOncqhpHQK1yru1QPr
gQQG61rpyypoY4bO/vHEAT3gyq50yKtxB80GI4pNIA3qysV5fa6NjRxbhXCXBXpR
ZYAG7h7jHQ0RY4sUda3tcW5ByY2hZCrZa1bttWDGZQvKEAMWy3CGG9ObFkpNEQ9o
geBBmIzBnsv4QvebmltnI2SGLLvAkHqAIsAsiK9FWFlk5uPb9HNTp6OK9e0eFNao
FPnOYIlnl71AMLWoT1dTvBNgNorBti+mmbYT8EXKP/cBb2m4cwZ+gObqeAfT5YtN
xfKUi/rK/HAj8XXdWR+jUdL6WI4dbfNnoygJiCmrElAHX0Su09mzP3dqjqTB+UBU
HUXxr0n5DgpbmsZBycwlpbNMxX4Bd9rGcxqhz/syRSnsyVnh5ndXLizLY9x6Jmty
53seMxo/wtgnILcyu4I3iuziNEmOqiTtGvagCMgxMl0pQ0qggWRw5dGdKq32NNvv
4lIOYHUj5VTHHIBNTPz1mKfqAQ00s15Tio/CdaIGpojZOEXVSzqs/rKrz/4XLcn8
68KC7cO///ksc2oxibKUJiPD0jsClNssJIu6kwQNI65J2xJ5fyyLnMWCoZjZ5U6E
sj6fpBy4FJfmUsc5my9A2pKOC6dvjfQZnP9wgkUh311nWDyRZ36/yfXV/i766hm7
CQ1pNdh+yNP1cksPwRbRN2CJedurtfZpOcjZRp3QL6OHJcDlF3iuQIvsKnBsGA0a
J45ccyjE82xUcD1o04u1gHDNupRZeJNDPayMp3/n1t9mU+UCm0j4GCT7qprKBW1D
k9No85Dfg8dvgb3kDn9e3A7DBzt6b/NXAWQlIGXEEgHlv3PIHfg//kB8jbvrIUEt
A4urnMl1Y0YUVLI7pg+cGJMwXDH7XNorywGEgt7yCTtfVoXNqrgpCEJc6r1SIynX
BnDWe3HG9U4BOfsrjDOGE7mTj7RxRWJjcqAlyK2E+i6Yrg4gzeZzerF/a4lzjshw
ncMwDyfWsTLPD/v/47bC2yyBTFhtjDIsK7i7la6I57JK4f5XrJhpQ8te+tAEPvQt
Ax1xAV6pCwd/jXHhNAxGntJQxVQvtyFJzFTtzVFWCqw1b1quutEnYBPQim8nAbVJ
29oKPtsdyb/CXRUz+EE/tEyK2o7FWmDCbatp0XxSkEVPq/ZeALqfUmrDZ3kWO0yv
+Bs19++NekOR1hEfygmlC0F/MbHPSHZoB1AOpP+yEfkSDNq1XBjmqaE4CCEO+AbW
JV4ZdFgx8k3Hhu85ARKgwpcczcBqDkRZNN+nbclBI83gDN67PvPKQ8pfOSd0TgSq
IVIWGDAWftXai6eku4QeONFAJwbmJHacgEGhZHIZ2OSgyBhoeajVPROwuYSnLQs5
LCTMK8DmASBJBGLovOfJmtdiOjSGEnHv28yrKU7zKFhNRBgHJo/Zy7RuAGPa9cVj
Qy2T6gsKfG3X8rooJEoMl3xUQMOdv64yxfQUUPB3pSj2vtJFmYRVx44uVpvU8qUy
V4O3ILvNp+y8sqzRj2fLvMJWwadMw6OnTJG3Tqnh8EVaCsMZzoTEZsGTMe2Kt/U2
Gjcx9crI+iOGo9TDQAubnPwCi55aTo8b5NUDqHCYmxOs0vChzALsNn/4a6j/2zv6
9s7l0keUyx0eqQeedSlS8BWiMun2CcJ+JjJO5Unk7cNourLe+LFRIAlJeySbvKsD
weG4RoHbrqAtepIcL4RN3/jGg2abyuZmtbyaZC+KtEVoRIaBhGaBsylXUzKmiIkG
A5fp67fTqGGTAtZB64zS5A0HxeYB7CTPj3xNaOWBON/M6N3+Zef9/kiGqt1bdqa2
98vmMmQYr1DYpq++flZlnUSkJKAMgweqLEINLAr/Fh49oqjTQI0R71/eZGDqjJtQ
bG4hhr4hiZyuVM1t33dB7idaJTznHUeE6EIu2ifvEQDgqQsB3ifHIYNlQ6EeXY56
FYNeWGj1ugDabyXcVRz2dtzEeBDpeqso7G3wf7lyvd0TnGPU+QbIWRuBD8IKiZ43
KywI5vdUOzgcLgkkAeCnXvwvTvi+/naZ3Rxa13SrogAXFX8VKkuudXEgnJChCtVI
mee/9PjXC0P+B3fB/htK3VGPuB+nYOgP6VyYN+eTIt7tf8x1IQ7spWHzFbA3vFOC
sxl1xofqAsq3OW3GhlMT3NRhxmtZbRH3qWhMBc4J03v1P+GpsN1WoyxWQpo0M8zp
wUH9/XEFx1MkpDY6lEt6esKIB9l/fPbE2sOnMzwCK33gDI+CLX7QxAr4m34lQDxI
7q+06osV21uLus3WVXW2qJEZp7XQoYv65CASobaVhZ5GKGUcOrYRv+ti7Zjhy6Tu
D93rXUD3GqQwxz7+e9Dz1JU7oNseBz6Li1/fRGTiEZh6aN5I8Bty7AWWw6oIiINO
GgwLa0w3kPloE2oo3Sd4rOApkk2PPPlleE8jWNlEF2pX4733Rsbk9U3Y/22sgLZs
/9uiflVC4AC4zFa+dy6TMsw03UX1/X5Eb4qkTNaLm9BnXejIHXVVMZvEBl2B/lmM
dRUn9Ma861zGmNULOEFs6UANFfmvL5GeGPqNp1JAoBWHGUvQRAggHEmSrjJq/S+e
BdDk2qjRITufDDYp5XvI//icFrpGIdQUcF5ss+erQnIQ+Pqj4qBQIAvE/mopcGuB
qOJBgGjUMhzwqN4/oeWitrxGE1DYLEAhntuClv5jW/ANcywKRFKvPslSyY+pBhlz
2cWYvTx6+SXGcY/4gEvdGwMJISPE21tm0HhlCHq9Py47tw76K7HqiYGP56+0/2ps
dwKAZCl6HqCu19sseTk9hb+YrWneGg/t4+WvaENG+/rfb/uCDDJ8Pr6rhXx5Qylz
vlWgvLINnwAwF1umxXulNz/pAAmyrGxoFSAzBa94STgpzbp5+38g9u/LtayyhGpe
HdxBs5oNp9o883f8ySgmAj+w9L4KQ+JQy2GsxyzLAMZTnsrT85kuO9uikfywWmkw
5LZl3OeReErHa/6nU57cU6zzvcljmrhDOWzWj/K+zgoGiFVu3LWthjWe3fWKr79B
q7QxQyMV34wDurOCx4Cnl5fSjDfdjB7nV9OCdJz4CCVepaWZyZ2J2D4OWfSPnFBh
wdQWQgIb1fGNMV3CqLe/HASnXZJEBvzUZIsYRZ9ONBeQJBYyj5ZlOG7ZQ4psG/I8
BLBXAiGjoXoAMNLT4OsE89BTc3m/ltgrjDsQFQmx+AWfurYaxQpr8YJ3RA9fZxvH
Uaqh3AIyQ3CAqsdPoqXlVsvMx/enn7fdOW3j+da7H2EuJgg/NAhp1FU3t9+x218K
CStW4wwtVycyveG449M3NhXmoQrLDVGiRj+UF4GWThxCgq7LS1zFAXwZAMYW9Aom
YAcMKr41XNYnwcD2w/1kCP7xI9E1M7HjL7KqMmMkxRtAmwXykmB9LGuXjFVWVy0V
mYwQlt1ytcyBkQ1n4mNcvKL8Mf41lIxonA5z+cpwQsgz2Gz2yj/l7SF7LzUKmfyw
rCEw+npsw/xDprSPa0eAnT8aZ3k+z2lpb+r4/AlX2WKcPmTqXZFJQgJHorAft/z6
W32s+82ifT2ilboecjR/Py1NMj3bYftAhUFsJ24058E2EiN5Q0LzB1o1YJlKp2T8
NcIuVM0bBXMKsO0Oinsjb8qx61DQLPiNza5trhlpBBjq5IVscvUuvn9XmLN0ml2Z
gH5DcAggPXO21RcNAOjHuhLdMA6BDTZZOTpaqsKH+Cu4OrnWBh0u9TMsOZMc5xsH
YbfQu9RBoU2NOlV03GwFNqyxemMsyw1hBoXxtzRaaYhSUhDQ9R/5mMDvw/5Qqcmp
BFwOyodxaz4rkwBXN2KnjWyaka+apt/snpf5eN0qbLxS/cn2+aAHnHktF0YbucDt
0Cb1NwAYqvQwlTP1nebBYW0n6/tfdwociS8SPsZniZjJ7zZzLyd162O42oXxi0Ym
oZHLkEQ3ywEVcKcn0jay3/lbIdXqaMN661lYzVvcE9gfHsnkswGMOMYLYCMaMfrc
JhWPa2dWK5JVgUVrNUPIyvhn26CNEtr49lyTHTIJCXk7EhM5ceuFeTyStwfCv/nC
mP8u9VsvJCOqgmDmuSlkWHvfHGnJX4pSi6ln7NC4zYW74xuuVjwFUEIhTjcPENQF
xnnOOJ2DetBsyXpbjg1R/2ASCgNs6Akc8zYJtw2PylVw9kzNdHXeZWnv60G4wsqZ
2FW9gtUCyyf1KN+X6EmZ1SW6JWiwAGU2vAhLuAUJwAIYpYiJySjV7iOk6P30YEw0
OyhO1+PrWGjl13K51u/EdU7ONQPIb/LdfsTntkSiYXYihQcdLP1nmrtynVc3cjaD
+dqnspG1VjKpaD9JFigWoFwnv5am0JvXIOHd9fSkCVLaHgC0IDDVpv7DHM7owM9N
AZU+dY4lMR66TW4e2uZaunPkCbc9cocD8wDA2evB2xZwfvgV9QhKEshzYX34wZFN
SUXF3eJWOCmOtaiivvf1t/xhuF1XfyEGELaet4ln5ChMM78Ihqc1+LpRiQ3m7hQS
cJephQJib7Fo3gY9HI80UG7+J9uS7DsjzkJYHKhxW3DhEcs+2hvXwWYbXgbFSwPn
09HJ9YCFeLvi7lE2olUQe+kbjSjjJtKKhBUaL0krIUHM/jDHDdLI8eb9aHqOC15z
O1ERrrD4CyZvnw+QNM4nkmYrk9rCSGya/XGxVhMZ2zfqG4k6RwRhGloYhNMDM6AS
TSM5+3b7lMobih2YQlKsUe7FDc2d7h/r2u2xkm0K5/U9Bb6bB7elHVHAB1beY/ED
Vlsvd4v1oTy/FcaPQvqIDRu7HDj/hqfcZ059dgXzKvNTFD9dCBscu8yCq9tvAEWV
39cZvkAiL+ZjrP5gH6gkuOpbUdswtYU4LCWvCxsAFmwx8oMpFZFCienzbSYrqv9Y
ojR34bGsMtJ3iujl33RHn+R7bhwtApuuBS922xCkRzH01wYQkWlI9SCejLzyaJgM
khXHXOo+XQ3I6y+uX/kWT27EQKcGvnPEu/E9vZvaHMhMAA4vhNKIaCOw9zZQPQTa
9mYsZ8Sc6HZh3+dxTIhRBchqxp+Aejhpnt+VTU+t/gBgy01PdPvCcASYSN/R8nuJ
KNUEIzvZ9GJM8TgSsY+qvmhBpwkLQ4eFx4LUOGhlMnROVm9AjsFUF4boQ38unBwZ
ULoKgQYd/E/jh2hYwbcUljxF7YCdyxhUQWG1CfxbifK95Oa7ldCbkfodGeglVAPS
7I8Feh8APIi9Wd37Bkg1tFtYgNGG5QREFHm0/K5T3FYTmdE64LJpAXUEhiCE/qry
q8oGAk2a6ibAQrgye/Qj2VY4p8VGvqogYQQ7QW501waCvbkmhORf/xeWfednCKR+
IcWgmOeeL79hJyrpiEAiydNTxMmszvNBmPGJ/HfIhRjNAIOy2Fiy1b6Qx4WzAFcq
ccAVa9laYYpKLHnOhskxJoQCdvSDXgJBhw/DybMPr7QtGz1QpRlLwSU1nIFCXPa2
8izvKqPPBcr9mjVMyn+dNmoF3Ot7Ffkh7l+rq576I4t07Y3Lnxbwu8uWgy6ddvA/
xayHaacfgNaZPDM8EpTsEg5ugc1o/NmC8hJt4e5dGIhc4NXnlDwRuNz3SF+whQlA
445LVnTKZGc5Z1SasgH+/s4DWNkqtQLnKVAIU+TuFwcrHDoewLbLVjLdHMHQyNrM
AUeaRfC4r/ArCDg0Tar70nb3xPFU7YpLBbKsThZOvAhyanJbxPQmhjMNx5wLCSKa
SAo2ZjPh117/i9sbZG80O4HbMHuASFZgO4OGT7UmwjCRcw3OxMN41see1/QOFzRN
EgHhx3uRSswQg93ZDt+YTLLyjWbqMqrB4RAJRMeTM4b5cQdNpK/aClu95HfiLtYH
tccmS2U3bnNT8tWgh1WgmPkvtNIdQTfLNtpQ+JLrfAWJ14hWXEJEoU7Zqa1G3m4T
CHnCV57+85RF8ZW67aVedw73xrtxLBLFg9CZ1aSUga+gttSVt2QZdndwXpvQRPDb
fS9QKpxYwslyq3vNeGGGnWD3m6BWfa1tAuAIThS2Hiv7GxtrhkgkxCtu58+vKmSp
zuS7Mc7vtWqNpvA2AD1DfhIODDwiuMQADFWIIA4OFoRz1BUUdhZKda5ConHq9LEB
LdSVIyiFi4LQmK1knHzp2nImD3z8q4TKaHDCGoZH/0gb3dnniruZC9izvmmHIvXB
GbKMUzfoTyNhfoevkXhdQzn9zET3P1deRgPmpyCtmGAklyw3ntXI5o/ZfE0RGv6N
wh6cJyDEXTl0RjGM8IELjm1k5cUEBnclj6ADY6nQiAdkMOM2T7O09WAoGXGX2lnD
5fB0RP5oSKF43s/w3xpF7+1ZoPWanA/J4UctLuufZfmL070iBZQQgq3frv3Y1QMT
Clj8u9vQJ1hSSpZvHAJarVTwccl+nRM/8RxIhr8TzUnZHdFUs87glf110XNsxDw9
czYwbY1Lb09XqJl2CWMaeRTzcg3kfviSOZisBpAZvY3R/tRpduxZnbkkupp0HeLo
8fMzT+TpmxOLzewW6j/aa/02jD91HHptWP4kU2Yfn2PjpF9N1sEKIVbQD699vIMx
1g/ud2a9lgdNG7xic1fkUsYJAdz6Q1+G58lAWB5k/nj+/sit/IB/Tc/g69VCtf5G
wNqRDyCToHTEU3gmTnUB1/hLk6DxORUnTM9jUYxsFcan3VBRPENeA6W8rZXxGS2K
4x9YDeFjKYXOrUYhie5WTb8FgE34D8n9NzzrsCP+kBuXm+mkToe3m32vkBCr0nae
xRaVnJZ6MSCWwK4adEBivPUi+GybpHQIcjZzECe9gsO/f90dJ4FS3oPAibpKWEQC
jHgbAFiw0+SwZV3Sr18fh/veLn/UhXiWkJtTsCnGKl0zE8ZFGL4YDBJkMPXqa/+h
PvmdW+b5S9lua5x5aEPfWMDbUYgQLHVqBLy/FlO7MBjn7rA9ISw0QKOLC/hlil/2
cn94VHLkcmCN82zCnFrVZzV1MbzZWByQSlrrYXW+T5Q0saOACFsYLGk+NfJnfRgX
1OfMXwqMfxeMMbSPqGKzjlwo4GEzbS0WtDUE049EjuDkXPmtS3t/GDnfKSnR5Sdc
2MyGfAgwVolhR8B2CdLU88nhR3J7h+pDsZLPuaFqoXQ51UMKNZThkUG+Quo2PG7S
YvL2kAN2WJbkgZylI/bFdfGrNFtY1Vj4IxRcCBixPTiiIlvSRQ2YvOs8UOJ/WIIM
DjeTHS61kJioTtvoAkKbOee3sFxdh/6Q9eAyiO/Z6MIYa5c5mQ9S1JphCvUgLbIa
IIvPBVoK+F++YcZD2CLgP03Nju6Hb59PfvuvSgHnI37v/x4gsseRivPLfD+xmNFO
49RCpDpNpCQ4nnUarliBbFc8vob8NFgyDn6Mpy+Iv/2lnfT+HsYEeA+o1R+fvKyH
Fg2QukZKFgbR9bUnP16q5hGuJm/Jw2FCG0vO8Y9xYiPdlxKfJ85A8wQj4Lzr1tbm
pzb+4UcUlG1126UgzYcy1vd1YvUnqz3NOEmcoswVprNh6QZG5H2MoobPlCqlsEwy
p0H4SMcoh2Pnsop692D0H5T8Th9kWrWLD8QZLqALc6UTnw9eNdYSrd+0WDEkjT2d
uGoz7vREeOaRPJODFAWkKB3yXe3yT6wFWEA43hktLVaJv6FxfczxaZpXt5yEYZ2f
kcUfUZUm16y05rMUtw1Du9QqMinhwAVh6X02ikEk7TqcXbZa2SQU51lQYzDNpmL6
lDbfSBMA9eW9V+M1B0rIMSWP/4n4vh3cQbIqNp6mKM4/azjrnuHeK29eYatp175G
gc3aNkS75XhHYG+SPg4+YoLi6OyHMsvJp+swEMTBpAUTo6ZtCL1KkAV78UOXMboO
Dugx45UX1JaPged6pAl65sMGFtt4nCGcQX+P2RpOQNkYftqrMBDeMHRTizxVBAIg
rTDuqyE1Q11yoUkuhLrtnkuv78S4yXjNB/oPTy49T+ldwH/34URTvcqGWR0CC84A
PM8um3XG3/QrDvRyE7C4LOm0jHbBaWZHLJ6Wh0kOJPL6R+x5oRd5lf3jIS5pIJ3o
f+DnzoJBEL0LF4qAtH+TlbmoQ4A+M+VHGhg6AtwEpSe2QemVirhxxezIUriTqoHv
9L/egnJnimvyxBdHvrFvRBMBuQr1zlE+3v+3NKz/3I3LT844gKAErIIT0ijghjEr
1QbTaryR8jFqAh7BzCa/p6amqCu8R2SeWabTcwigzR/6LaU2ryEHmpHhku9clK2j
U4Czk/SKCxxuNbIBVNcLftz7W9zp2pGUPT7z6OFxj4KHLXt4LStsIgtwC2jE9I1S
yVbdBoe7wXMsfPLLPkdmg9hYt/xjALBjmMMt8rphVw9IR0cxI6OBwPiknADwSrLh
AMkf7m8C1TCWRJ/FpFX3ODShalAz41R77aCB3WSqCkTQyGvVhbAQ9CRubtRAV32j
M4dQfIQyq5821ifl1eeTMQKFHK4MKpKvnRncDRM9yK1MMCBN0WndfRea5BsX//I6
kV73RUSAhRbGmZjxoXqUZtH5uCCErxrCxIHNkY/KVvz1rwphFLfbrlfnFlr2Vtsf
fSAx/xKCTDmPSn8r1glqmQxyfKzkGjvrAHuXUXPIjht+hzwlugdM2YneS4uiNHbC
9KoB3va5HVImaKCFKK6sYqBR9+juFVT43e++ikMOQjZJsO/me2Noh/y/94ysxslY
CS3TSVqWK5gU7eUNCbPNRtdKoknoxPdgr36dlGNVIWGTg3FlWtAIOlI85hNfGq0q
pi7xWDH2AkY+kdV6oIPLtilRrVUtZkS3WAKLG6vwWrBJKik2ItMsXudE1ogoRFD5
Vo2RjKMRk3MhKQMUWjrEeSQ3ekWw4kcPITaf8YeAWVxLqoQSm+ItSealwUveAcXb
47bvtYNvW3reeiMhObFJVqEFMYYoIMvUnLz5q4dlS/+xbXvZOOU6zKwnakJzx78G
Z7hQ9mdESxX/1JiZnz2bZz3rEPfFIn0c11yLhQ21sV5XW6CzT9mDY1sQAoyzTgCs
TslWO79/knKHPWFd38WJI3hgM0Kd6yJzXIDmxcbhVkEjQk49THU78uMdSdBmh/8A
lpPQUTnghuVkMOT2sPE1IuwcKKnDXXGvsvwIvcNVrrlU+rw135+Gh8LWETv3s/Zt
gmy2z74HI6UTa69ahiytvc3svDWzMdVrOr1UvIZ2RszXLS9xHkUdZd0IKh0YCEHM
vaRVkkymz7lPIsxr78hYE4q9zrOLYZC5wnAKsNOvf/wZbHwX6vau9N7RTmLAlUBU
0c88jeOL8HcqAl/Hw96fhJmDQtuL8mAvn1s2brb4CT4QvoeYc0AIwC/zPWn4SOk4
yZhlEF3Kl69UgCdhUZtlEfVUt/UrBzvQTF1YWbs4ZskDutAbnEEzIfB06jA/cVAa
AFcHbgryGKvIecYaXtspcqtagui/9dbaKDiLakrnXsKo4k7d6xYONwyd7PraYOQW
JYm1eKvyWtxfx4OZF1WTnMYVOVbmWkt8l0doaHLCI0/xBgJFQ8Hl/cnXxRG3dy/W
4ZG1BkcmX4PTEczmxBSFv+L4wTZ0N9HBBqC1I1Y2Kl+14+3WvWZ8+83bBCvepHyW
wrVYikHM0vsQ2lGcq7ySPKxdJwf8angd0DVa5WghR/w7aH5az2W4utj9YP/IMSmv
2eISCS2rpxigNuKVyraegdKCjg+d1hJCXsRGX/0yfrTZPWV6Ad+xRbVSSS9CKoiZ
7cJHe7g+GVk42VaABAl6awYocE6DyhedZRLw41mEcDFRyoBGCWIfA5ZCmCZ+zrDr
mpur9TrQXvIQ9ZVnBMHb80rK31oGwycfZinfrpPpsFvTVUQftEizVV8FxO7ySlGq
p+qBxAq5MA31FuYM0VI/2pAO6HztDejbpKd5kONQCAszvZQ2aO9RX1kOQHn135xR
1tHHK24WftC6xce4GmlNxNQ4zt+TzMRyALR7+4aY0uzSP868sKKoCmLFnJ+YMm52
1LSUagxA+UUYOUgK8Vga0cJSXDY1loHJqdx71jNXtYZ3WjBEIkeOd7PY4lKrtMH+
bOycF+Lc37Sd8W4lOcjZEssNKL3Zxja0Q0PxjGNPuwlLK/S+8JY+u4Airm57yBQn
LT3eEbZSZXiFn/5ApjBa7DAFFFkCi6lmixKIV06c66pwx2wpN/OBVoYkXaDakz0h
1JH+dz8z3vYSWb285/vwvVezWA07Myub0jIvGQM2pdLF0gSQeomGkKnEhy+qal7C
2xuS9QulGQRvgFd/fvUz5wtx2wOJOWrsO+SsJFImskL70oj1qX3kZ/YEAeszYDZk
sgP2fsQlulwpUKeHK02jsQCe2CdtVljGOj7ykHqwRe4BQ9tN4gr8GrLF6ay/1pja
a29gHsvule42vKnpCKgmG3bgXRLpwY8uEENB5fBva03cICohV5ey4QavZyvzt+B3
ws/WoaqugoHhlRE9B36O7KAz7wHAVm/iks0s1HzzkAbE2RlzCR3F9yQopFIPmCSi
7LQjxlOxCReElijRdS4VCT90cF9Jtufd3391H42Oo35oX4Y2xoUWbp++iTc86B+B
CBXXJchM4eePtJ8snT1XIrRoHO2hyVTLNACfXtIfRxX3O7AnuLE/W33Djn8+iA8a
F8Pj6EqrhrGjfcLJ2kmmPOUZcDiQrAez3IONdc7OqW9aJY/sVKYq84Pio5fPe/nL
p4ckwp3zbJn5y++roonWGSrY/Ny41aXXocHlQspXSidLrDs/3/FWKDFLysMAlJOV
KmyDoenLLvlV+6KMCyd5wZkbm5F8OoJd0egc63kpwIWsiK758KvYYDaCvSATQzln
1Mxc/lVv6UQmLEmkA3e32+lRkg0WecMi8rCTAxPsgMs90Zz0MVkrdKKQBkuoXECa
ywy5CALoPnkWL4YdfLK8IRLW/AT/njXQwBJ4yx6HrXHyQdwxL8VYzENGxuyJKdSA
LjePIBNx/NPqnV27MR2Y7kb0dGVqU3hAzmXz7+moBvAdEZIPgYa4pdey1zf1SUHk
QXNrWPwDmBN2KFssS/9uABnmURd6bB87NGCALnfzZgzSP09aY5iM81MRdAon/mu8
S9t0HXmtF3DwPE31QlNt0Zbcgl4QiL943gErjbvM8btNBCwylwKafqHFFK6SQA8l
WGrgnIWs7qFDlhP197gwP5rBnUW2639rxfgQsm8+/gxjXCLBnEXRbUUuUIwZSmFr
4T2KDZFf4NWTiilfw6MGMIFMXmLxG26MMrAGWsnvHJw3m8t7DgVXze88lW25PMpp
JwI7tfvD0te+j5Sto0wr+pEWlPcnRjV6pozQuhx/1wKaiHxlcM9cH4PnBdgfKHul
t/gyUgbgn/mRChaGgqjq+ff69XPzsKPcbIyKxJSUAJAYwHDrS2z2iyQNTv/gJG72
Iyvd6QXR7vWJZQqepxlUb/rrEXhXdexgsPwoVmtnnzIaqyytgMOQK5m713qL4GXH
Nn4msTfRA8Qo0GYnpYDBY5GCytAkuj46gNq7PpSN0F+prG3U4u/I+1dwxC6tIVIC
gBL6eJY1F0IqhjkSFFfSaYvlpIW/AJgfyAjWYjAftU6o8BlVIqk4W7nzt28vNO5I
h0hxM4zaXEJ3IylWA7TU09gG+4lBOMdLrG3727MuYf9mm9eTVciRImAL4RDS1Pdf
FM6qgz9WjQsajIZm1JH0pNdY4qMYmg372Hj8L3814hgztZGpWU65v09rQehDsiKc
bJtO5NfG+v5/YFe6gk8xX4XzXpHirqOJEpl6hu3155BcDt3b5gnwIp2g1CxYKsTE
2q0ZlSClS3EwLXBhTim+h4q88wg41PdXeXXsNLmnGkjoYuPtuhHF1CpYUdVunIps
A/NA6gjGRitzCZfo8FRn681fnRqgvkc554Ra8bHe24SFD/64ftts4sgm7pLPWBiU
+7s5tzRelFj90wo4IMt0NyuMJNWwd1MpWkdmn9S6YkUTPXPEIRhputdE1zSxyugy
2QL2FWmeVQouK81p7mm7VhgHYZ0s+ZeyJnfwlLTJlOAxvpyiHJ6Jh68JWqPivGiH
524k1wzAgQ00VKIRztrl7BbhBt/MmYwOWbHaIaS+EZTN930d2FkwFEz9ar1o33Hv
lhzr5D8a13VTQ08xObPuZTgb6qoC0SnzINZpxvdiW8vKpcpqu4eKQwF8qG5SP8A7
6OKN3EIGTHlHu8pJev/Q5hBgxyQWJ1FCSs4WiI/tI+V+YcAKwBf8TGx9HEOZf9T1
GhV0SMMblZl/bqc22B62vpxQ7OsKnPa7RKSGWRfaKLgQZh+TrfKB5mKsCAvY2krO
pm3n8PueAHCOn+5De1QcyrnXGHuVCPXJm7JsJWoJLSW7zPvOiNBxJwY3i0bBlUSW
OlT+HLVKNhhknqxgh1m13utgjUBGJEl4vgi7WCppUVlPjZHnYjkNBQap9tPgw9mI
+AzWTa6cD9j/VJvFKeToCzYHkBlwFyPhek15lvpu7UOO4aYYNZJwsX25N7PBGIFv
lnS+auJb2p1TfrVyrALa6oZ3dwtbctfRzI9873hO87ZDTX/CZAjCmIIvGI5YwF/b
/zC0UpJNcuFBOhuMtIsKIdef7RvhnOzD5DNeblzYFbL3j/Ftw/0IKP1d5VXHXBnG
gqRB5chY61cb8miQFslNOXoEkAMMJCPGVS4iC+GSFOJyW1ssis8oIRoUNCd3Gjm/
x5aiROPfczJfD+7TQX7tCq9CFs3/QLKEIMnyjSLNy0sXKw3HbK0o7G25BbcYarWo
wsXlRupO8KY3sfx//CILyQ90gbUoYQMuYddYfBziviZezI3rwx1LBf/u0D7Uf8Fj
UqEKeB0KV8l0eNRwQe9R4Ipw5srlvEOLe6j0GZxeQuljgujriFxFqZI2dreG6/A3
FoFZNTxQJQrI5WgrW+XQLWZ8gOzMn1jmTNMOVMSnwFznm83gnq/A1U9WfwiZkteD
mS2N4FlOpisUtI/jp8ew6rjyiAgNEAPxvl5Pq8wPNu6acdJCa53JjinKKHHS8/9P
EoDAR6cHUUiIN16AVtOKhsAoGycAR/WdySwTf8Ml9Aa4b1loxK28Rpb1xpwJOpxJ
Fv5iUbaNnpSog+9rr+5LA+z2RpWXQThjsWcTesptRKf0UOrhIJvD6t4EhR+bBjqz
TYN+7BWoRobO7Z+zmWaZLraMzgQRy6hE9Lwbrc8IXgGzNvWQJSVqX0bIydEtepvX
nupGWquH7pPlriAMxNoRlSWvE0cLtMns8i8Tnbf6VzrPSwiRlzlnSLz5oPFfLIQh
xRNO23Ha0IJAZMvQ4K8YIfom2t9U6YtcfnPgMT5esphY56L97gdYt3v4o8tz9Nnk
NswQP/MJ7/u9/Gp1PNAl4AF0yPbsVb30mgiCwixUkTppeQPXqJlS4uJRJ5BwGoff
kQGwJ2BHeCFjp5Mwymho7sc3Y0sN2wxwSLl2/11RbtVcnoSyozBOrJzQawj3BPsh
q7sBWFIanYRst7BFGM5pMFvw1xurgSdSR/ut2FVn4EBj8iBm+GKkF2tR3Ifqv+pQ
F7tIrwbNw75zqS5sjhGbu8E759Q9QAIamHfASs1zCvuPxR18aHiMCP+yq5e3Fh/h
zYyue/QqgC8ptuHnutbh84CEzIDBdK+Me6SgOIdNL0jzeMlonN8tkc5yHEA41QkW
lNb5B76piSKELrbMnT7AU3FOrRWTgC8z21anO2redAaSsCw+foVf+6zcvGedisky
UfyddQK2ndsSN0XGAX4yOB/0pb1jFJ8YxlFd9SkGCB2FLR36EvEnqbi9YxuEy6uR
3sNNB4Lw1K5WEcGUgRytNPm23Epg4WoztzTRLiDpX02K8GHc3x3i0d6XQtvQtJzA
gdgOBpRSOk/r9kFRY9ZNEk7Ot5qYh2o/QVFAFd/LzFKCt0/R7iXi76idINz2EoS9
AVwiOMXfrWqadMsLIOBc2Ko9Pu3l4rOMUiDyBJZ4JFimo6v8xivmIlq5tLpri6hP
ftjJoBwPJdny5034UledFGFF9Lj8eNYsHdeLdMq2pn0/Ag5cU7AZejNZi2ATdFBX
EcH+Ow/R5ttoSa7nlZSfP10EKqnrhtPQ/fxJEKhNkPjnLnY9vL4pGO91FXPGdPiS
QkF/YdH2GvcY8OhB0VQqvcpOSOkIptA2WM7jx4l7y2WVEmDV8gqcOeRAFO2wwl5G
3ONE9qfCtBfUtcIgAuAaHAV5gtc30iEIiYoVU6LuirZZxGZ4cUO65n6q4iv6uc5j
9aEkdRJJ+x/+9ECeZC/YCnd59PI531jTbWWFHD43hX/4c4r3oVYNAqIuw1NP5ykM
F/btw5cKEwprWKShUfDdxLsAmikz7dxMigcSbS5zoDszZ1Dva/U4VTpoV4S9Z7wJ
SoQg2jdlCMo34D25H8uKFaif8v/jOuW+IjSSEVJAXNrs0YrYGVzdTvE9kCifVFeQ
taEgX+QiFgiI51/Fa2GxMipkrreqAvpHP3x9/eAw3JGfhQfDe0wWT5DKF/r3t91T
EfHPSkp95LowC2AW/7wD44CjneV1gf+K4uLo7rGrZi8EFCKCrOER5HrKynDaNgJT
1FtLoCbnr7RjA/gxegmeoztxEdESxxxzIH29NVzA2JAswa/ex3Hlem0B3Tzb6xFt
HSHH/gSBqvIoiQd9ZY6dmZIc55DFdS51A/jr/Qodc1/n9gfwoOfyNlOmhR+dd8Sc
3pIWlYKb4W3JEq7EpHH2PGw3T5uSFKUDi29b95CEsr1fjyzhG3BgmTVB6eCsvJeX
yYBSJNa7ybdiDrTBvgNUJuKsWtm/RgE8NroLazbKsrLA6rWisCVSrmUh3xuyU1mJ
BCsM8nv35Xbe3JSi4CwE7k39alpLQ24LBy1Gu3dCaqy/5mP6P585sU3r7Jb6yJnB
yjTzxBHP4z/My06C8/37GJmx/yT+bSm3ScI2yOeiZO7V4hw9kikUMU50glYTRGak
0g/LmdEBc3YPBYbmOonAleTw4p4fkjGR1Xc3R/a6ZZyBX5fva7wAASjZMHHFMbhx
j2oHeMbSqnyvbN7p/TCqWOGdkkzod6NofKoxeJMD0kG8wc2996vUf+DBaRs+C7s5
is0pZJp7HtoVy+pq3gczlRQpBYE5KIbWpkbBt+thg3uUm9FjlU/Y4SHzkwq03SC+
JMezR8szGaYGrwSULjP6OpzxE9jsBtRnpR/sufrsRyM1FtsvIO+oBUcu39yQvA9i
5d45OrEPZToSSBnQwx3By1Ca5ZTIxGeHDEVqOQHBYw57w+vdIUjN71H6jq6+qOeo
TZMW4sU4AuhNIVsnBLLxctwDalCSv/qFcec1oKh4sBxBt9pcQHReFRj6UKkeNQtK
tOXWUXDHmnEW3F4v99HojdpAl5KDhKu2dXyne6HgJIGi8jhjGZkKm3/re8QYQI+J
PfVnLykZGdKSVpkVrOkcqUXcOzaaGRaL0fMv+XprMRxDWA5nOwdlbQuYPNmVxN9P
B3nxqOhZlfNF+TLWrwIdzvRZK0+w7on7VaPXM3u/jy+JRrv7kd8u0FFZTLfwBlIy
8QcrVzrdRgKoJJGDtKjAnjzNf1ubhQSLTtDTns0rDUyYGFfRKpL3IcYzqPUpHD/o
7nsCW/WTjuyD0Kjuq9IHM5AWwrGpCGqQqEu4G8QF/p2Y5zSlDWeOTMz/9dVKgFrK
ubJmLMXrpfRbX5TwhhQQBZMevPOiVRaHCvztLf/4Wa9yrC/tt5A+0Gu2LZM4mg6n
CiN7X3nDg+qQKCtHoK8EouwNQJJOhcKvDXXW/ygBaQP+YOQtGCs85654loqU7ilW
b2lxp9IFm7XvaORdvS/Og2xXFKCbCQjxuq/v6Z11AvKZMlqx5uJzwrgM+oOn9Ukm
IiwZ9MBpehxnnlURDydfAvT3UBLKpQnQVVdcqSIW4HO51qyJ/gmux53+K+Zw6m8I
OiZ7mqCbLH1/myH5eW++K8nXg9oqa2fF4YWFHHzXq25voHI+wYD01vQ1tG5aXRn5
G0haAhDHk3ezr2UCuJnNMNKPGlLrONQVEc9AaoStsiaW7FQnmhE7SlpU6NHbY2YP
6T+iDwUCxa+q9MBI760R8fhfTs7JNKLwOLqdVrgaQITAPMnx35t92AQ+GsIAGF2W
ZfSoNY3o5pBjak5GX7gPRbS1Z3Pwa81aMuQRftKOcs3iS1xtWXE26Pge0nsG2/1E
aoir8hyt+WFqiI2xMVNF5LKI1q2NQNptHA5V4KXrawzlo5mBn29HAHDjTPmqSaX7
iLFjecvTRSplabR92E+4u68Zf7m1uvNWx+oMsEPS4IyAM/Nlaw2T8BDJZrR571g0
qMfvju/eTEpJQ2AwCcCfiRxwwAHstWuITbi46yWuSKEoEkcrhEwj6KZW7Urp+86f
rzpEvLBLKwwfxcvG/xqMixrZbsbYYFKbFOnspVHVaXUOo0ksBQmbxVz7Kh8ACf19
n5IqOPWVZGmr57g/LHYi/g==
`protect END_PROTECTED
