`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RhkeAScNoP70GED76ftHbuqTwaeVfQfltKW8WuoNuI6Rnl5yVnZRPQGgZwh+YAMr
DuJ/pPbZwVnOBj09tYnjByh6EZ8XZ5jBd/F2C/0+sTrt5sc+zDZk3AtvmFO2/hz2
WNvHiCP+52eVywkkEgVACw9DpcIRxFyyN7kIjyFTDoR6+HR2ZeQ/eoQEaRpfciul
/egE7OSMYBw7Wy1Ad8jvkgcQEs9UOW0mY9szh/Epyvi8g1ExoXhY4f64ey38/wei
kpn9Mbr34sb9ixVSRfNW+rVQAZpVBpAbyxI0D0fuabiSBXXjaey9d0IJxLZehVJL
55Q1qVGzF+Z4bl2+pUCeFBKLIdqeIBZ3wl/0UZVDsUd6nIA/954523xIfF+9Jtxe
FAtwQdOjccU4ek8DHkNRufDwYvHLT6/xwEP2tAXNGR7U1mc+jc8CmpPWZz8O5XTN
C9Kp6PxifNpBsN84gceFtvYZv4kJODbz8mTPGMvqjMg2FtLRiT7eYZpYZJMV2Ter
aNI20B3XYgjwF/jMnElJ7ZyveYg4QaQsHr+yS30BiLNKcyqQA/TCO7r9gHOHYnv3
eWqQcrodIAUUAhxwLBJIWvcuk7f4x1Dw7CjlJEkcYDgzNyfVIfXQ8M5TVO+VV2J/
XudggAy+12QhybbOMBCiF7PaRj9U3Jg2OTxbCzfpjhlteDMWhaZOJUTnsSFcraVF
MU2yk43l2NDk+h3G6YMxWFlFGHaUaAVMKjiEP1H3AmNTjQpQtkWjvUxyZairT1dz
yg7SjcJMiVc8sdLB7mGAyQ==
`protect END_PROTECTED
