`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3qt8ymJDei+SCd/YdeZckOfLd5gVjh/rfZkk0jbb2ofFZMBUa/Ah1s8WqCH+rCh
ORymd3oe/EtNdlabzX5nVZLnb0ZJacL8P+ioPN72QWHf64i7zArP2NIykD37WLE1
P258d060kcy6nQqdQEHsC+NvBCLxpiuBI1kQCTLpF1hz95BbNt1JzM81nIg3wMSk
qAVty/nTdA7b8niRlUUPbVLwi6UEO68+SPyH432h61E/V9sIEJhF4c1wpmFASByz
kES8aZpWFtk0BsA81D39ZLT+cS9U1HqMHUbYMFykpvDDYj4ISuvvRYowOhoTD4LW
3knUaTiDmsgP9VP+V3XiVgZRRzy7AaeKPER4AIHnaXwUH33YhHErTyPSOWRiPaio
xouFnSP3yLLQBJGf+slnbAZ15Uc/VRZXFkzKaDD+aw45Wn0yydS0+nAjNE2Kc5Tu
q9yw2MMVCsUHs7glhUEDJjrTgjAN5DC4/NXDIAnqpmByZ9K1Nyjfa/NhGbH/gb26
6xC48y7Nf+5yBOyWa3C0ZYPjP1NpEbhMsoETAWTrerf4BVJESYTBsJGCgUVPG1WM
gaa3JgsvbIIRfj4Z/dpU0XeFEgGUxfvrWFGNKJeeGiWVDgF5x3W2J7DAeuBQNkYG
qB2jrBhQoClhiNbe/hmdHvYUibjzWmULZBXbsLIYyQgzwlONQgZeAmmONK4f+GhJ
FYTvZgecFw46ZvLY6ANn1JMwQU0V3FqDZp7XH5Ce8KlDxdTLWpN366cytIMk5ZPy
nWQ37gjRoJidSEenIxVgJU6zsZAbYcNhCCsJ2JzkOvYsgTA/8ky8pGC+PyXTReaM
FZjBIW/Jv7yPbcFYsI4jgcZ+m9xeL4ecPHtFxfo9pGUBGZTDX9yj8XjQFCV3H9AH
fd1PBGpRMC90S5/vF6dZqhm9AvMt/Rri81hEV5VTWU/QI/TKVlKGookEwi9aX9BU
EUmgC48RExoToiDKnFL7XCIkrLpC3R+tr0pFa7Ppe49V450ThSGTWVxkRmRnv6ru
6jH5gaMwoGE0RVAD4skV+4YnNYu18906mzENBDBFUoPamIl2Yq+q2iYo1beRqOjQ
aR5J+Np9v94h2K+HdJDwOvcrGF8hOi2WilwLf8pEKIfOx6W7PXjGXR1VAkmsXFyO
u7kBbSTrZgGcZNxelJECCIeYZQupaLEG0b/4YDtmlTRzZzP84e2HarM5ogcBuC8D
YCbi7C6DlBm6L6PDbtGiytvUYlGZLLrcUoBMtmNFxqGOEEvdhLtF6wdAfZvUd50q
+OGyup5rYslGbc6L/Km9eAAwz02RmzGOZqA/0LuCOCUrgL9WprupKAS5G1yA89UE
aI6RYj22BOfizr62bPHdjl/FbNs38rfxd4Ud8nCgNLjkOpDja8zsex+iRDBn7g8N
mkV0eciV2RSLm/nT6hoc8rTqN13avD3LcVQHPG2eTyuc0xfHutgokM04T/0/eEAv
rc6JU+mR1QFm515jsLjInCyCX6wIKZN2FhX3WPu1KH+0+RWQeskSRifbf1nDezcv
fA6ORwEt5AvD3dTgsu0aaA==
`protect END_PROTECTED
