`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XIMznGP85lGlsxNn7E1y96Wgeau6KWgyUmp5A9xpA6k5fS3Wza6KlyS4KWYGh+YE
y8jS/jLDf6r3/yMa4pFrUgzfrfUsDuFhB3PA5EUehzNkt1O5FRCabU2sc4SPOGr0
puEgHsBwIFr4YkLW+WVyqSKT0+S0UkYU002gzTp2LGXSFAD59Ud8jJ4Dh5cdS7JB
kHfIFakC7XLhD2l8tjrGHAEDbp9+kqbyAAKNZdepmEoLicDF6TR3F2yLsSXdhN0v
aH6yqs3mGT5HWKurB1RVHP8uGFc1op0Fdrhms2+bsdYwGOaQfGZeVi+JuvG5kMtP
wX+VroXifWRvI5Mt4aFI74OHE+QEeoSEQdOad+UMSd9o/Vji2BLqGUKssIqSDxjN
hkTBUn1i6PVw5OgSsRbHPyCuLuWdVwaqDuVYo5zu3F2OSQ1bmFIeYKe8tgry56SW
v/oNIh7RbwRjVOnC1eGNZr6/uXD5Z6A2ciWzpdeuVIS3i9XWrErpEjl9nZjgjL5K
ENd7hlB5IDBKh32yXU4vW0QGIKnIy9edTMpZQiJY25E8KbfXx6jGaIgPGotQ/Qn2
uvn54Lfa34PZQHWV8s+ogd+Vr6oFgq4ZDjZpgPw2C3Q8OYgALlq3hKzchxDr7X8g
mLw3JS+IgG2AsZYDZQthir9iPyDeeY8WDLhd6lMvFucM9WBg35mToPdVnOcdWjfL
EJFFUMn0G6ohiqXImQD3sPeHxhxWCvZuKa8Ts2hVU8VxhISkGh8Q17DRsporjHAY
sYqKjKRrIe4jM+HhBpeplhbmF4u7+0NKK1xdFSddul1afUMUzWXRdakV6DY0lOEw
4GclivvPtJnG01d6om7/ICpB3goaapa26dBcCii2guiRj3/I2zL9qTVNkiaOELBZ
PpxOUAcqw1DZ0r1Z6jnbf9osdA2GkvAQhcupiCd/yl4EddxX6gyhf+o3KlxFOh8z
Bc1FS1GBrSp1A5P+2Q8lPSQEJI2K7GOx7Dfcg92Grx58C7TXHhdGsSYalqMUn4gP
4kiyzKguvywyxI/OUilxF8Kcqtps1jnkc6EMgVcO9ZkheiduTEMWV9RWxF48N3p+
z9ouUufnyN1/is1lRhbKBnl7bKlbc/rKMVwtrV78m+rpNDAMhNKghny9iEDPT+fs
F1md+R4SRNICTUyUysKjpQVtBU3603eSgov/TOY/axTE6SrRKjmIGMs75Tz4lf3A
K8xPJgNt2OrVPB2QWC0Mz6sggxywo018oYpIeTnf4m7VLn69ny1QsWtNjk0kYBjr
6x0EF6MiNCg6YqfLuD5z6J3RTp8bXdNasTuFSYEEqBr96R+Z2QdkF8amAlGGsZQE
y1e9c9eXElmgL6uu/WLZh1rOvXVwy/FjK1BfutrlvBypdUTEhqSrjWL17+E/iYNo
M2wcM6xzuwNAKNpQNORI/BXS9uMvonuzqLBCbTRY4w1V5aCPkqd5YHYJCCe7mPPC
iG3iQhm/+ETQyhoKTtNp3FMHAXBE9XODIow65JXZ9/x4gkqQuZbhJmOKYltHG5K6
lK0Pym8+ZOz37TC9VXvL7UT+zdbo5/qoET2rXeeYuglPEmgt3+gzFD10rMnj36AQ
28X++hAXeURxXY7MfV1HCsrtTCvgKAiLrLeyCjQ+br5/1rSo4ry26amKnN/Bnaz8
K3dSlWQrnzi7hxfk2G/l5Z84x8gSnm7m+srOeDLEkYJ1DTtfR7jw233iROG3kYvb
/Y8NVjoL/Y0mCTiYGGdu2ci9U6jfiOYohAaWDsefFFY=
`protect END_PROTECTED
