`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1KpXXPZO/WUxHI72DJg91aOd0daD/J01uzYHZsG/XfJrOKOF0AmqREVepTJGjysp
5t3/a53ARVW0e2w6tByvDtFTtlefgpf3qhNZ1JBE5D2HldmYlhhbrWp4Ss4rfJ/o
HrFlGoNpEAZ2EFl0XCYuGOVE8J3INC6Z1M/pcBfcLeTP0N0eIZO/JsjXiWv2xMOf
+koExQaOfCHQETXVlx54CJrwqDmTot3IPXRFVzgRHHOMgvyTPFm6fzevx+jy3Ytl
x/6hemiKPuRVZjDFg+gpR42y/J+SXRayH2NHvgrB4v27NKTr2A3Z6qo1tcjDJq7y
LIU+MGSFcEk36Cg2Bs611VqvKXcteF0+qWsfYacXFoS9Z4U6aSN2FwXTOl+f4pFE
GenUbNhSAoXSehWvVDXp8x5OPQ97B8MCZr3TneQCXD0Euc77WFePaIwpasF9+63P
r2wCuJc+hPZjKgUz0DT5VZm4Qt7Ylig8j4Sb7R3M1Ly/Cdb7kg45ytf+jdkrJrGA
uyyTkLtlyF3IJwgrVx28PATcyf0kiOeMsjV7JLD7fQ36z9D3XN9JbLNpuW3sCLTo
bSGqblrZgE5wwtCp0LsDViXlOr+hkltcGoHN4h5GsfXK5Cbj6MG9JGFkin4m3Qmd
LJoxDzVNi6+MJO0afg+nvmi7DFMxA5fmKoYZQ2AQenMhreMsvyLPY7HTFdZO1+lM
4xRKeaJuQYVXyggGS+gfPQKhjptd0Y/6YkuaxXhP9vXumRxewyzMbxi+1lZDY65q
2aZl/P6j8UQidcAQZjgpxcgAvrrmfeknSmdrml9y9pE=
`protect END_PROTECTED
