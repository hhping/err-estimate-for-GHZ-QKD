`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fjroOl+Zly3b2+CGEWilt0SYM5wWnWuU3BtSlj76UqKuPSfZnAIB/hHULZiKYZ+
i422rKjDfI6aPrVqlDKf15CJu7d4xApiCikhcmcZgoCNh8rL03rG+ZEzzO0+PGN1
InNY/LV3338B82nkHYOrWWhwlkQT2hByWCwxXgF+GMRtaqDuNIusapOl0owt3xcr
Jgwq4bKROtMC2hqIrZQKOehi4uQaPh99Db+E/ox/HBNFQg0HYrQjW00UNADFk3jR
IRS3K7onK8JWqVWz0dJKnOdQIsJwLw8j63w83f74xry1iHH8+tgDR07GXyxnvVth
RySKgoQicXtpdO4+0loUlavNRN2sJZfiXWRIHFaVTkTM63olDaHGPPHuUlqwWZEo
i5NFgCXlIJw5rctynMOXAWbAsSrKblHOR1pC5o9UgQlbzqRaxL3pmNB6fDOaBBKA
FrNxRs/5HsPQAsYau8/PyPjSAH68046i+7RuG8QUyDr/lnPJyiXVqRT0kkk6DG3I
wnTwgfvvXefwNMUInQI3TtoNOYsAHne1EEnNVPRPO++4bRORZ6LbeurFk4RVt9Wx
AIrcCtxuTF/ITF89IrBaOyIhXjuanwP+WXqh0tdy9QylMpwMPEMrd+nLzDE6n5eg
JmNofbkxQtzaLgSSK2EGGMxOvVa7M85t9BIbOf3MAnLidCSv8pfrSlEE0S+GVSrD
1C/OZbDhgmiJ+JUK2O2nzp3QuX1aFdC9SXEW72gZk1lnicI53gY/RuIPCP3X/5cv
fQAAD9Q1+esApFwonNtwA8Eudcm1stlfqqI7/ffQ/H/+R+SFc7yuAFZKMcF6VGJF
Vei48ZCVmChv5Qe8h5ITb1LSNYrckg4V/k9HuuFMC2A5M0KSSnL/xrEqgJs2MmwI
Sz1di+Ns8EHxbCOY2hU/PqnkOCh5dlPvNOE81B1n0u/7vIDS4WSGWrDTRUV6GSxB
mxqNVgVaAsxxPRf/j3e4lpqnz2eVNOAHw9kH+dZuj+ZgZrtt06vSpqBOvTC51sP/
U8OsgtIbWH27ERMcv+HMU9k+woHYReHx10JHmJenj20EfYxjyGtA4/tbjI3+MJkO
h5jJeKJW0/vUEPzzZ+vCZn62GxpdiH+5oE69SEAN8zh/0aUYaPSdSQjy3LL02psN
fouz28drgbM8VB8dffri2iMkymfz1riBRIRbpkWxIBGQBr0VeIuur+TMf91bLcg/
wq+GvWQMgoNunrLWFYUVOf3lWYihGK2/Zgrf791M+7DCKWsqatnlQNH5QGvol5UD
x6DXLDI2EI6e3sq5lLPiBhMo9qrxwsZljjjnldBrnXPQLSxk1O5lz5WN382Xqjs7
`protect END_PROTECTED
