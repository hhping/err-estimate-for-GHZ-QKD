`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ec4gdoB/JC8w4wcS5MrmVc3GdYw7nJHxFmQrmZAVeMyLwUkYFapa1t+DknLjPWOW
p2qlY3NeOoj8yUkq8lzbDNttNMZm72YNXfCfxZlqB4GlYGehMPsFWBczJnCRyYCr
Z31WCGxv5oVC8s7OU6ITxgtYejbzTqbX7Uynoz2wmCl8ZNVfySJWpCmy8FoQBkX8
HYulu049obS7UFXw5UuXem37VfjoV3A4cp9Q+j657whQamz8qd5wSUoD0jJmfDhf
0vfxSHdAGax6ysIQwvkE9moRDa4LjhvRLNYptnGx/XloLYLdVYJumA0gsxi8VWpH
/xw0wbDLZgNnumok35dDo1Mw9YrWq6cAPJk7aU7gdcUaEM1uutVs8ByJR45djlXr
q1xnQmTwEIKhBKtRs0Eg6Xr62RtinAGkhdNxUtO5jzK/ioMh3Fg3qoAQ0zZaqMYC
P4srA15KStr3SdWwLNlPhGEj8TFF6BrrbsasaO2EvhaQJizZc01aAx8PoOlFsOnc
JOM2cErNxvSG4D/mA++O0afkLjK7xGx1ilXJ+en1xkPRnvIm+2vOTH5lzbtg/NPp
mCn/Gg2NWA46mUtV5YJBgPvAlnThRYlPaMZyDL4feJonvumxUhNOo0hz5ryT9gP7
kb5i3l+6aI2I4vhlt/y4XxdZghbhPbafRNZT6YDSfmoCUOB66CX+ON5UuKw6g2ec
RTm/OlwAKs0b0zXdXBD8NQ==
`protect END_PROTECTED
