`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrvl90Sf3ryG1sNlMCgahU5TARbY6HA0NHgQfubTRJsZ0ubP2eHasV0+VmmfAbmg
MFzuFLQKeMLL+wCYdb7Y2mCGEsgymsg2nCVPyU7HqLSuEwwZpXTxlcifIqRvjd1F
2k5eoHKUXcDTJuVZg1fxWx5fV4TXBzm8WLTZi4Umug10KME2TzSVNEkLF+xwrsDV
2XgrsMzdAM7bKFypStXABc2hGUJMbfFgOyp5A4vJ6KsBniCM2PHC/3qY5GJxIExx
rR4FumC+FJPKakJ7ZFkeZGjenJ7fEUuHrauCLnpT2fwzNLlHqRg4SeCs8myNOc4O
l74yjTs1+/cRELhCTqwru/1hC1Tgx7CUibX5mEPvwwkCXUO48IRCiwIVcZ8oRLwb
FfyEe6jtFQuk5KM0/Rz/xwOrNkHJFySIm8TEr+lPwxU/Md1VXHf/miz0hszT4aXq
IxuX/kEgSE0ZSC8dCtOj1AQDRQjlbOeKs/mVSySZ12fM059LGtitIKutE5JEkTHe
jFI2bURHV84bgfGO9KSNZLC4KQAN3LCkv0S9OnJa8xt8DRHtggm//1uzM/Y+8Bdj
3ppv3y8fMHguE6rjWSpwasY6CiozA+LKGdvsJTcxD6oJ72wRltuBTmhq8+cVNu5L
9ce4RxfS9RWMkCGC4g0n/fzSwhCIwZxvOihY+u+aYIAFcVqe+C+NWme4gm5oDIun
wShHBTr0isnBP9xVCBMaHNOJAf6iCNS4T7Vf5YWRjODz5cAiyMVLntXC6uunZ09R
iNHCMoO7cK3m3twpjyDt2nn3IgjZxiGv3z59CoAzhknIrEwIad3qL7bLQe7bbCsh
ueUixuwadYKtD3oczcjzCX7drdAYpyR29RXGTsag8gf+YTf+YKxyUgNlGQ8QwDdn
L3OIS+Sp0Ln9ZhqsKXNFXnve2C3xNnvwR1O3aW5Sg4Z9OOLDOprbGJKISxQTscs1
zqgchWI19c+li4vWHXrjUtjUyR96UxynthVksjiZm3Hf8KYqUrNdcRCjgVUn+ayk
TAgx5uvplbqZymFHbtgREkXCW62cUM38gdOD5bu5yJQ9sy7pi8y0J3VYy0Mx7Qj/
uILE7ChOQru83B0IGSG0KRxCnA2Vase7xbvlnjV3hnsYm0r6MA3WXszV6enFhJHC
JmDw4hbO6S2UilArJLJQxdFA+Q1esljeLa9eQ5CRGysgYm/Pw1dAuD+QA+hsnIme
WLCG1AveIdo6GWFJNwjdpuplQtPldVjI8yzLZeoUJxglTZXbJa494whghyk6ovKM
VFKAtgxfMswi5Wi3Lcyq5JdeT8c8z7o+vSKuaVKcIdgEPDHAptxv20ol3OXxq56N
BDOUDaZh1/d17wtmXt2YfcD8w81hvINAsgN1/o9zy4aXb1V/rdVNpxUBJfQ1xNAD
nbjusKLagxOUIw/8CkayaEot+c1G7u2cRtTS7pNRYhrdU9luVmhQ9kSUorUTNuvG
Fumrb53rhft/RAvlKrE1Px8j1kr42QK8VMzYb1qRJMqrP6ZnS0xPWbsr10u2BWJ9
mzOJGARs0/tz3/pfF+edaZ36cVb05hAiEdQnK7K/3AnLQw0ZNXm340AnaIlmrynr
0SGQlgsdoe9+Zt3WuxP7B9GX8Yv+ked8DeJvhYxx4cbsTyNfFZMEPK+9BmJHshPf
KZ0m+TPEZmK62rInk93lMppnFXvh8yCkKVbVy6zUKm4lhnGo6pSmaa10xhXL2EYk
llQ9TtjCCG6YwhVRA4gXNQE9n3jrfSoxAoyy3NiamUJerLnhZw1z3jhuIRocNk7P
RJyWGNojqWrli2MEOZ56N+HhnZXhblCU+TJk6Mv5UUFM0eg5zDItZ2mGtmVMHRnt
vFtHEeKdEjXokvgGJ9Ix3fSDbU8MVf3Tw3/vzzgzR9j+OLzMV90+UbquoVn65UM4
FOYKd2QyqVkyqC1Kc17Noo0uBTYJ9F+3HcZnJYaI912DWgS90D06WGf6QlB1guAM
DFdi3YGFaisgJ7KBx5c8pFlU3Wd5RchNATtHLES+fMgizI31jCBu5gxaAwOnRUbD
OPwpixV79Ef3MZ6tuVAu9dIknq+FFTQiNlhHY+m/PW5ea6gDrOJfo34CujZO7n5d
XkLu+ZdNaG8ZoEyANt4y1GxDdZLKktTt1ubNGF4vJA0R3q5biGWjmRlteRuzdyKp
qmTCABwN9rMgjmhE59wjGsCgtbe9swdLyzn6UR2urDZBtFo65ru/Q2fiwtJ582PC
NnXxKdhUzQZR8zJp3dni5W2TWyxMHbySEcBdVmR5yiiOHGdTOUvaLi3aahM9kkwD
y8l/RyByoAliOCiYxdwwy4cMQstMjyPj09BlGD4uetGcL20o1ILSsaRdHBDIFzj6
kFGibRVCf0u9ivGNhCp3ZVCOm951a3YtdTjIiyUVNSsXoyKxio2baMJVnhjhT+eC
IaGKRU/K1AWNHyjWMMY71mr/gup1nEhfBIb95eGkJl7FpPaXNU0NTlydM9U/V2iN
T8RfQZV2GbVR4d6iWqvoXEEmcYSZ8c+/s7tUquFMJaNfpBO1NhwyGm3rJ25d4TX8
r6Q9KJvXXuy2QEmEj+mI8CqvWLbw3gu2QV9c4eNQofh5UXUHws7oNgNo0ep7G8ck
hu0VGky8sigeq697KAfxNMHK0P7FYamFIdocCzftN0Gp4DgqADAinFB9SewHCZs3
ZQAvED3FRvPEiHb4pGDIVA7n1Y507pLkuh4NvUagjVEhxA/8QbbppeuQcMuZjGqU
20xjON27A9ivDkmVCSqVX1T+9byZwK4sMIddbq+TKav3+plU4yi/h8OtM3BR4tvV
SVNVg9wsXx/F7j8NuqFPsKSp9+bdwdY1xaBpafJRwoXahV4Qagc0JRpIUxwpVG5h
lZUbNULyXz+hwrpRp0HPp7zoDOnNTmqJko6xhx/49lbc7nNXM5JXsVj32oBZH8iE
NnOLwlSqanfA7Th0r2oHRa4Sax8984qZer+SwcLMaeQBdFfL/QL4BYJtZnn1K0Vt
H9aG2ddoB34XRVG/MIcHow==
`protect END_PROTECTED
