`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rFsmWs2sbIfNuzoDsDjipFIAS8jpxFWScN23qy8oIGaQTfS013lxB5im+7FNoxw9
GJQKzZcp7v0UVMIKuuFN5rr1ZVkiLiGGGHSyZ1aBZITPpZHSPbnyTYwoNkaXWUKT
FzajYdktKCcqECR0Vw45XAZN9E2ClCtn+U0DbPFaBudTxpANV+mLRzugq+w83FXt
/FgtBlt1G3v4EFprhmZ+2YoMb4p/+aKU5L0dOVzn1ltdI3KkEWEyWKhMcs8/AnsX
dFy+I8YDT0KDgMkx0nkxcogGa5x31cSxsrIk3RcXK0j7bfKGOjCH7aAGQfvBcCIa
3pFFGaG1KrOBpRgzsgAmL3hE73B/Ygl24JhiJCqy27I=
`protect END_PROTECTED
