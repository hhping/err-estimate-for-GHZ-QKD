`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YflS4toSe6hy77Jj34Z6l24Y/PSN00G4FrlnM/QdIy+ERQT6/3KOuqzpkvnZEr26
iv1cCRXFOGTXEWIFNWP4Jdgusrj4S1tpT48v/NkCcJ6Ky/quVg9DNZ/LIvC0qKIo
ctAwdTScWg4jPb7mf1TYBz8pkkrepE18gmUmQTdmGLWpbWc4H5DIEAiohDw+H5Xj
2bpaUVjjyAtrnXGcj2Fze7ILdr5gVNARdS+TzhG9BTZGn+Dkydp0tUZVRGsn5TrX
9AnkRkLypU3WLh70e7waV/g4FpzfhLi+BqxASnbjuMtJcgbTu3uC64mFcSNSwjFr
CpqDPvzYQ2Yfn4/6CF4GM231KmAhfESIqgqVyErZzrLd2DXzCFiM3eIu3yaZt4fP
AxGSh+B+MhjKuWrquciXfNa5toATXjA3j0h6YexyVcYZyv1UchBxiS6uBzlBTg77
b2uaFuTvDZpDu+D3hMxMhE8gxlRxE3lVD2qWuMAIQZ/k5TOapqIrXACCC2lWu201
z+1/T+chfRFn9v4D1lZFYC7pcnH3xb16swZ/9yduy20xNNATGls6DGWieN/oPuhL
3rBcpHnlgEV9oPHguFRd/b8fu9LoHedqAfdNMN9X1vLkXVR22xU4rX+/5wNB/N1e
/847Gh8pL8OceAfsR/WT/OvYYR4bPt5jvrWWtRYAMRR9DRSQwqdzZpJkVe8rWlPd
wgNRu+T/keNSauO4lhbngfvpRnH63LsLZjPdjylPnFuwtadPN9xi03LSxz0Txs4D
vUx8IJeYBZl7hCVs/4UH4XK6voeJuJV1viAKCTv3zkefcoG2uRbqSupRRO1P7rEU
T/LcTnK2diqeNuEE0dTuUR6qaJgbr6BddjFIvnSRdlNhMZtmWW64/vh493C/GXrm
+HDeK19WCYvt8RaXtZ2orT1imaGS+ekQ3oJSq8yMHs1jVEe3y0s833ri8SUZcBOE
uA0VSnwU12/WF+giyopYTBTwzP/fkF79zGTF8lbnKa0u0hxQjNDoFJCAOE5BKllw
ZqEmVTERz46MB/AVhl+sZg==
`protect END_PROTECTED
