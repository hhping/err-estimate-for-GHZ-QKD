`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGUXr004QLgVJjloqd8+SjJ7w0YcVXAc4gi094N+uDbBQPS6JZIQHjd/udC6kxgL
08EEC6R0qZFQ66Ep8XLg7o65ZIVXXoZm7/ciJQDeMC4ZtsAahqgAP8WznXn+Uefe
2sGqn0qk1HtFnqbeDqUW4EOAbJhHqpMygOa7q9fU9VxQT9gxg4pHgGM39AceJgQ/
y7N+DOyDdkCSbJVDShplLGlTEEVysrlq1CamzBL2x2ypqQuOEUI+E6YBgMPvokew
hthsZx3NkMQd88gY697TkXMYlu2jRj593ZSAtxszJ8QWIQfGPYGBfUmrgkeE4t7U
9vWp6fnvNXi4GgHWco9SlCYA0rLe3GMWT5SmOX0KOq72X/YfJxAxIm3gt70nOBT7
f0qv1YVr2rHxY3VK1/OfDQ==
`protect END_PROTECTED
