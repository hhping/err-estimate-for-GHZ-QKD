`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WAdbTn46oX2TQBPwpPo3nNaL4IF51gR/I5lAkBKksPayCcrCduz2u/RwXAqy8gmy
2B110Bkxz4xxroc943rSGm7ZC2ykp4wX7MQDGN4rjhFLBoE7ZYDJX1vHLlRm4ngv
xggnyNA/kVlnqHdV/Nbkg8o/CblUskrSVjafpv61OEn8S6esB67Ed35MxrUMifMG
5fdcID+HPrs56UI0XyJN/oF80zp/Dcx8VNojGNPMkfdaV4oSGo9v4YfmpA1t9yJ1
Rqia4/P4FSdhs9GpRaakx0gKYNnwr0f/92sY8b5NUzvzCYPO7Q3S+XTrRCOzcKv8
qFwY9+IkZumRBTfebYfnPCUIbGz9cVvgJiFtmhM8QLrp34eladDgH3q7v9imtQ1s
0xAKbfq9ARJoHisrBOdmpxY6MXfdJQKS4hpV/XsGq1S7iPsAGtsOPh7D5iwKrv5+
wwdC97QOvfczDkiWnXdbnaTsYsbu+UjUe6MB1R51CoIJDYbPwnAvWNrVWK5txRR8
3ly2ei3mNq50v7Auc8LdFsF1UdcoNdPVYrif/pB3tiB0IiK92VhutFknYH7n337g
H2V9ALTcFHbtmD8t4i4VnxlOZs1K5V/aBxPFA6hIuOdg57NdiRRJG+n+0jJKCmCb
qmhB/emoMeoIV5T0zqzgjzN/0O6TKIG6h4ijClN5AMLFoHhqMh/lAdPMxqXr5euH
wxR+tkLLOu/2vFPrREBUcjAKV1K4X9GOrQzh6HD0jalkwY+FPBIPKvTbDqQ3boPE
n2VHOUCsDeLwxVXzWsur+qCmPnFJ7YQQA9CANaTsgQGYMn+qNnhgGja/IdcFZoPC
uyk/8OIuFJ7rX+HVyiovS4/y5DFQT689odf9c9mcLIafxI9HG6D07MAcV3XyynLN
As9HjkPsUVh4hhd4qQvxrg==
`protect END_PROTECTED
