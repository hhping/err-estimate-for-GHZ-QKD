`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yfEKq08ypvLlMuH4DLzLl+o0U/oXDTOxYSJRKS/IdkOITm8ZdmnAFPaitDhNeEs
7xZAwp8eqMsKPwzeIQ7adx1zeVZfutR3oACBfNZjthh9GjyPY5VnSzpsGJGQ2/tE
g3t77+ORivwJ64YifCehQEMjXGrou3q22Xdu++siejmkdRyLylp1OrrJ+1qg6jSA
PfPZrNFkafajkAOFtL2QCr1TO0BEAWWINnvWIGLQim3gA9X12vYVGGBmPtiJNz+q
ihdzJbCAZ3qyhjE38WT+8Ln+1sjICOjnQ8jVOi7XvkkXdunpQaR1A9Eq6oZbaJXQ
duMA9YCZXbI24xwxAdNNpKdb9jpNICs2s47kUpNrJJn4X8sLvJ0EKaLcMn8yTaIo
8C3gEgTEjJxaqDS5PbCDs7BuWi3L4waPbBeGtLV39i34uBJeZidiEMVkIWZ6p50I
lQ0qH5NQTUaAfm9NdQ+zOj9DnpiJwtO4jMkSr30CdCsjvytaYK2foVtKTodGkQFY
hV9yOBfTjRyJZSUFOqBQxihO2r2I790gfM7kNO3myadu9a7HI1KDhJZRD1FEe3Yg
agV+XkgQlJebgy1IpPt9kdb8zrhSpqWnK2CgxE3imXDVy7iQoAlzlK7z5GKPTBzN
q0BDbgaeWlw46moI3UHzrqL7R1Jl8wpNuRRBNnnDBTvul0GCJVd0flfmzyrO7K8P
xcVislqmZXOuhbMJ2+r7qbqC81pjMESMhYlAaFdjuSFbBakWwCBdufIVKxjKX/ec
ynCxkHjpgIuhF2c4EuQi8JPqhxBLGJrji3mxrU4B2I3b2FImxjutKICdAtxlDdNs
LqzDSZPMQW4t1ismg/UO1lmtfdDlNF5nZuZ6/44RRGqJV0G83Tyj53ppncMBS5Fe
Uob6ugkUeT8Kmk/t3ITE4VzvwMAngMo2gnTS/Q+knw3CRaLrXMCo9PY/6CGwTrM6
lUajPw2KxmloALpaWcySIpsiNyhTKW4Dp4SHKzpxRQG3+zYdoZ2ynTzu12IHjfqR
7qI1gGdiuDsuaqYJlEb8XeiJVIHFGMaO15+9dkZJXChBSrmq4YXUBn1ZofT6cMXi
BpzP92iug/udF3rLccsquAPmcleDIIVgVORV+0ciahqNnnTlfJSJjcW9S3B/qU+8
A/loDoAMumn6ziNxXT4pBEqnLhleZm4+XZtLeBsj26XpynOy9eGB/LLAM+Rbk7YZ
hwkcSsjWswtfVqYrGdcClH9IKWDCix1uxkjN9YOlQ29iY3k9/bMR9hgZOkyEvqGC
dxg49MNgY3oi2pLUry6RItM9kC0Hhu4DyROQlGvAtJq+54UZxvCyqevhTZxMf8V0
ywORuap2dAFBiVTZd2Jfn5bVKrDoywC70KhUXpDw+ZollO+Cq5EdND9nGTTIZs4b
tKbOWKMgx2V2tu9j9Zk4D991J61iHK2nL2Ekbc24nWDfEoJ//UamKzhcy3TzemTd
fYYw6VFYFqIolgjgJVqe49EHItg7mc9/1DV83vsOa+iehz19oYF7QXKue4DpuVhv
2/eHOSyxyDF5RUN/NqJN1HoQenSFBrRHJgDu052LU9PnSj3I29wgw++Iga903dSZ
voeN4OByXJP/PdxXYr9MpMT3dmZieVEl0javK8l8NSklIdM/Stk2muyShQmeJZK2
CVFnsbfqnmVtQkEQMWlt70hP8s0t3ng7Z/NfEzD+jzLaptxTn0mHPxmNop8Uf1j9
2WVY9NohJlNHLALX5OetdG5/83Fgwf6ZksmIMYJsx/sqJFqrYklfTm/sHHAP+gG6
CwP1CJFa+aTjH7VfbzyWpHGBS96amiimkpJGesruE2vL1ttKrfddr1x8xZdmRlru
Fm3J6BDNI6byDSAZNIfChBwbJdIEBwd7B8BQPs2o513MoC698ivo1Cx+9x29MW1U
jczc09/qvzeFhJVDK8RgcE8sCLeTGokbVqOUfSrjM/Jrtxdahk1mWGJSX6EFDAgW
zdhbI6fUUrbfUJ4l/R12LiDC1aD5BOFSz5Ooj18M1P0XbCDdwBGyffTKLflucrQK
6KdgmF2OeL8GNLcXy1PWN0kfUfYAIw7NdrhVdnHbBlRfLQSJMN/Z0rc6BUhrbJSO
e98jnD6JYUms/kcQA/QJ6scl3jqkhjqKjwy/c6mFLKTatkZgPhKWH/KdPRXOGElF
Ltb7sjKm5hlPJ7rbEXIfO+Js0RVfoZR4CeBiYr0droR3XT+bzLMmrouyOBoURqtt
0dqp7Ej4HweRLp/qD9rcN9FAf65vSHSK7mB4ksBCjKR7UTzWh35mDC+pW96KKK/+
xHe1OLYRhysiQF17wEM/Tuw/mOVXqZGhQJAPT/prVf2rcik1OxdFD6xKXSP9VjPn
gZMkEAOfLn21/OAc0g2L+Y579njY4PFg3qZE4QzxkuQakFpf+gHC2JPSYktwa5zz
d8enFNR+sZ+Sce2eZeVwRzFMY7pyW2G+HieZvU2fHY9kp2scrCKQfp3vllfKHknX
4XRp9jmIIG4UVwhBKXjpHWjzrNHTUZVwh7be0d75uUslfXZH7i+FYGOyF9TGM99/
YHSFe/FO5dwns5tWqrIFYpo7/7tbdyrpGoJvRjjdzHSHjBVg2DzGB1n0QJ10xlQV
WQgN9/G/scx6hktJ3PoWBzyR4B3g7VGp2Zh6SIn9HBKhumWkglrhYERNP5z35Rpw
iCVaR123zipV0VEU9POnW2IKCz9son3P89rhivkAdRudDUg3S6wrHGzbtSfnUmhL
NRdEqlXcl1xDllokkx7Et4bPGTIfGRUHgwySGxC2FYNHBnQU0l73tcAf581GIHtW
7zu1ULtH5Fc8MS3Q1HDpGVELYBomdUTkIyxqv7x2RMWd4MbHLVUAlegwiQIRFY+S
AqX9WC4J9b4zERH1EIe90qd+soF8P7JGmzxvqQa2ZlC6ES7gztr+Tijmi35FwUcV
K7S0TefHdn2OP8j/ks4Pv1967PdQXLYJQx+ihcJnq7nKAAJBNuk1kGR4NfyTjBLE
GmXVV1Y7ZZGCGgs52p8lhYp2It60IUqQBElTnR/gBsXh30B7JaTnWtYRqrdl04Xt
G2Cm3Orev8j6THM8kqv3KbMX+iSkrVaisYXYBJw0b3gCLmkFJFc+y4/B+blvXpMO
SIlWcpVnh8IhhqszO7B+F77pP52F1uSSvrNLFdVV8wwa0jNB2kF8Wha+wSQCKBlY
ctd3Xefq7wEP14BOsSxjwtVk+ZG78Mi91x6KmaQXlfVQv+qlsQnF8s4X+UNTaqRL
tXxhxrlw9gvZbgbnvdhhxqVb2RS1oQBV44AZUSmDza0nJMyoqK1/iMa9XpBthclQ
vJO6TPQ6TwaNzii8+DA//h8enw6p2ha4yqCpUUmQEE6CVyW5461TjjgFayHtV/yV
awHqBk+4Szcp5grtu5VKgrEaMW+8UbTvqyWO7DT90XlO3wK51sG5z+25U+A2J038
NHzN9PfA7jnBmtCkKBza88t0rrT/JCqzRfSC0ao1X848bab4ukC6oFgayP5uOR/U
41N0mbur41JKrol8faLC/22rDdG45oSpvnsQpLU+J+FU4eUKM6L+bLg6H+6aNoLC
ez0z9QoL9vYz3/nlvNCwP9Sud3L18SEk8nL8tmAXVSuqj7oxvdUSNABg/8VTkuRC
85XM16w/hF4TKfG7njhnmcNXCTiCuwFFCy1wvMylLjqAKHz7OsecRTJ3thi0ujWT
u3kdPJLFWd5dZh9GLGx9FB3q3dZKLoFfvfULj2jyOqYQFUIegg2iivYHTsHxINdY
w46AzNPk9OOFb4e1x+yXGwNVhPsFBh6DxZEHgx5oKPiIwvCAwE0KV5XNn+bvUz4s
+9mi5lbQPE9LN8Zc26gYxCQxMdlvyEF6Y7WhWuf+jC4aNyibya9NMGqTz+3UepjL
9kJgUUQPUEW3JU165qpXQ/PdgMTWSQRZ/lSGqDQWhHb45Gods5pke8SCFQIoO5mw
gRg5Hvxmg3Nyo+pIY8Bx5fbO9MI+QFsCf2F6OMMcCW++xPgx64WVwQVWJe5dad7E
SfIvxDUTUoXcT9ROIM2cak6lNJd6B0Qi2UfzscpiNCmfRwqr0llRfJYe0JilakT5
p+Gz1oi8CTg61dcQ/yNlwjENBz6MB+h46t/eIPPR+6EGwr4VwW78JZfifmNrHeai
xVznOx2FWQNNxS70qYxJ3wVp0NN9XSlKC8GqNl6k9zTD+SZdqFfzjDT/M5zz/h/Q
Ubw/m4DlWO5aXzy3YPRqi5jk0njMxU5LeTxQaNU/zAuhCESo+wp2zVmS2mXvC+KI
8ilMvOdkSrDz/GOvumZiaI+YHDmstiwXqmh60aWILyPmVwSmf6DyJf65yetMnefI
LGCosHp4SaBtJM6VNDTk5k3L+Lh705dFUTgifI6TO+Hc6mBscoZmccaRypzHga9C
aml/owEptOK5ZQF0FiSK38ZGXy/dWTKUGm3LdwURQ7tKqesvzD83AZd3oEBlxG+R
Enw6keFKiB5+qscvqJmEG0KWRsPeW/HuEC6KPr7t9u/6Z+axBZMlTMSwXx9j41v9
hjaqIpOXzx8pYI96K0+45f1OJiFAsiE3xwis/Ba2E1x3BfpzEbun7FIcCwBANZIe
lK2y506Yb9qZ8vc5bkTXPqREVyreYrLyHaBVntPTsKxu1HMenXbYzk68NoI9tk2v
8tpG5rp47/D6u9A7JR9HX6UEVrOBIWn6q4zfb4VZu6s/SmS0mvdvklQcpx0U6sJA
WgR0aB4UtxX49IuoDmHjYa0lFI/5QxY2reuHFQECD89dSvk2isTenjDX50Hj99AB
DCVeB3sqrtxydA0I8fATQBo46kYSuyaz1uylepvStth2eSt2EdgOJmYbaIUroh/B
IDfEMFM99Hg51y1COatXe2ektVDebqpTjOWS0vMa3cyMNA/yRZ/x6iYPw3pKa+ht
Jn08/U8d6k6cLaozu3GUe2IxSU85l6L7s0lrSYfHomOtACEobQ7xuPCIlam4idos
LrdnVOP11DlySZDuxbrqxILnyyPG+/8ySwG6FBZvtuEQlMJKZEMNcvBy0H47t8/N
D4d7yFwhYTms0Rc5MgbbQjyx/lNlLfHtMrhRPOyWmRgg59Ae5W24fk4udmimcxzM
lg7BXVSffyAozxbyT+UOD8+2I7sOb6IqlkyAXLAOP4cehgpohEqnh4E7qeGaGcVY
FFcXskdhCAxHsnbiG9Fdrn8tWDsZhKnrCkeuOQGauIMR0eGKPx6VNmCxrx6VZ4+S
kzwlzIPI6BOJZeyeNo6PLJviMYg3uk+llTpPBcc8vBj+psgcNjNMWdmjuBqsUjLQ
V40pVleLSx5W5NG8BRxlUc1mtKR1EZHXlcetIjqV8C06y6RDftHYILXGL4fsa3CB
U3CcRCeloiAIt9WUETNxwUYaPOKYk2wPuD1rjeymjQcMzCNFbXZ8WYmzfCj1pjs1
4aWisfICTxry+ZplVvoGVStXk2P+M5tzhEfrISlxZoEi6IWEF/WA5I6kVE1XooCu
bnaI6bS5Pd4tfufN0OvjOlYOl4qtek6njApzZX/iPSOg+5BprJXuKCqkK8VeYT8z
B0FVQG2Ql1cOxBi/AcbDp8pa/cb4otcLfNDNks1IvsfCP8vtX1DoOya3PYLUoKyC
pljykQdTGADZu9UTenNdxXIooxNQWRX/r/VEFY1xUqDyNN33pXlEFfjE3HUia/fD
L2z/CxgEHjxvnuuTu1VufdDayy9QW+ylsPFaIiolBYpg406E8chJD45De7MdWsq4
+/4YrPdQ0hav3Ubh3YX5ubEMJwo/77q3WU+AwannkgDu/riZXReYiR+RqNvl0CBK
YwTJ2ABZewFIs9PKx+0NsVHdA+lSWA0StzlVxXfeY2lOQ4pYjf6jBWcehkvNB+ND
xX5la2gYyQGlodqF6EflSw2BypSVhXs0KYjFpkQM7EgZqIGcsY4vMSxfRmQ55gAo
el/va/LP+o2Eil0sIxsRjtSGPVPh2xB0OXGsRFVCc536mLZDcO55eZZY5jaVr4bN
Skf9HfgaRNa3IRSHjLBzQlo3v720jOy4x89C1AgTA3XPbSFSG6PlAy1y4daO9Nvq
qG8rGbVJ3Vbv4/Nw5HIs6Z7EiUgOuzqtEffHqdaDV42FX7jFwQ+mi+vUEG7Yu2RC
ciytn7YRCMLQDZPlBfJd+KcJndZF+J/+N/wixeU+LIX7KZ3rCs+YEMVTu18WB5tP
Po/NZmpwikeMmqWoeoIb8hG6Lao+9XsoKQEFQKX6xjiO8iwdQZhhD/smPWM3TJDU
O/NmaNL6yqOdMB6ZIx+QL17fWUZJKl6+O0fCzlHB1CNpjgb+/m6QfKBb6TXIBpUC
rR3fTq+7u6oPq1PZPSVeMtuP0kSrtfZ1UT7L9rehOv1qSYG3Q6hC4o3h0SikNwQw
RyYRKgPvMc4bBF/t3EmUYo4rRq4PgSohf2W2MYF2CdjLtIVkiHNHUfPq69huMCMt
x617Mxb6C7RVsuE+IiFXaE+zJTlSvgH9iO7cEVuDbUhf3ndl+oY9mSJJxoesRWLP
ldw0Ntlqk2AfMWos7CXBEnjuGM3FEob1+oQDIiM0v0BI7qIkEM+q7rQBmIEBG1A6
n5PQlSXCb0wOfauZdIuD8dXEb6cdm7cm3vn5tHudtEcnyRi0ng9NWqAvXMC46UaJ
oCXh7lf6O0KGZWn2GrkTRSiqJh8bxnEiMNfplIVTycWWU30bfU/ClEPuTjKpDCxm
hh7ekqh/XaXjehPqliVleLH+HQeSyOqQYVGyDujsIGS5CpBeaDfkx8fRLo77i1eJ
GTwcrW8QYUfCCpB6BdPFXF8/vR4EoItRVxeUq0JWMkIs3cvnQh7kqdN2Wbb1NF/F
MbcqVlRsmLO04sdS8Aw4hmpoOTy137moUHcoNZbBgm6d1wL4H1SD5GrUJlKLWWgJ
eA9gG+zV0vQ+yE2AAB95v/T8a2qxytbyAZMAyf/Q9OrhWjypReHYaFAX1YzgZ5EC
Kg/zfVzUjb+VW/xpSzMt9v0VNO4yz8mm/CK+o8jP5ZbhabmCk2wC7KSaSE78oC2r
cW0GXtvZbAaozrcqcpogT4gYjEHpDjAfikMi6kaQbLgfSDwfzOvsl5gIf2pFWZEj
DlDSVMW66XycrH754aWLQaumIPNvylPjpAAPZDc6b9aU83dQgvlXJGEY9BfmInnL
7StYDKvWVk97g+ofw1ouInz57Gx/7O2JVaRGuqtP3VK9bVsA4v6X41y4P1g+IY1/
ojsHs3vTjJnlKzfM32P77UlmkzTX3rzUzkCeKbsD+FnmTGIv5AvmtB1hVqwEsaZ+
UmpdsjBDlBb7jrMYjVfjkLOPx4TIJ48hR6cv86IVhvOFq0N35wnK62+usQHprN8i
uaKuw+5cGoU+kFRhVmmnvldM5pzVRmY1MSMDKMMOuIRilRj4Am/JC1lFhNYBY6XN
BomXJg29WlODIW3TUfq5NQR6tnP9mxhWWUfHLI7V1pNwe35r09D8WJ3wS2SjBUOH
VGO2dXrW5qv+r7Z2JQswLRyJnNqBZlVoPdF5c+q7GE14VMLqT/quYvnrvpLB1i8u
GrYVSBsph6pOAf6kn3ch78aUqffuRBWzDaDTuxDKSh+L0ituN/3bUuLia0zAvs6N
n6ZuGMFI7meBdfetur3/NAjo1viNfF1CHL/le4pu5ncp2yyk5BiSJ+FopXNGxE+w
arbDbPElldIczKCXCYQWplVOvB8nrSphohSj1ZrrxeeCu0lXTg8lt8lqmzJuTEit
JFMxRHvBvuIuhMRjDWEovCxCsu0AymZCquU98X51KSGSA9J9Qgp8B7vj3dD+fTG7
P8V4DOLpfUhbGNaxYUcX61T7y5/sRrsoy3V4h4uY3UbyhW92m3itacNBq7lqlpNU
4azzJnlBVToUv+FVa2Cy5LiN+V45z6J22LqorC/7lSOpLGvDUPKSURI2SdJB7TKT
GIrfQBAcuttJUP5Ri+YdztI8qRkOQhqWGYbBTGLnCmo/8ONauxyeUaKsoLrWi1r5
P92EAHLga2/AII2P2oDh2iITYzrMxakNrIN8+jvXJTFR+d8sxupQ5x72h0b1rt1r
Y3a67aRh6sHdbvQVnqkzWawF2Aocaxv0S1JmdX69rqThvMtY6Fiqh3bZPW89p7LL
d2F3AKcLbXoRGHAHnX7IQ5WcBz0RUg1zjo+zYYeaUJ7jfal2CHmK/8O7vRUGpj/R
9xzwQKWHdkh7FI2NZ10T2XZUDylH4TMNGCykm3IBCUFHeW6fktE2SqUv8NvNZTZP
zTr6jCdJGXoQMquFWjfJG3gAzbHMc7w31BdT2PFc42GCFJPFRayn2WxO8f2Ppjei
VUgzcPFgTPw2cFC+VsYMTr1GPNzRufbMTBqYn4P+ZNY5ulcNMS5XERjnnWMyH4Sa
m5s0HTvR/ZpAd2Z0tBFatiYJvedKjUo9Vj/+lRna54bTvNSE/E510Ha2lFORRE1O
nMYu3FMF2W+tc2Y1oZvbB3X+GGCTushQlop3wVxm75UJsiwTOIu/p7y9ZNVy1hGn
W4s/EUjLpw2dwL17eU7bJhPj2HO25fVZniltMEfNhdeayaUCza9H6Y6Yi1UOGWxm
fwvF5KDTgktvhOmmxnnQR33xx2YdtcnojqI2GwYkHBMxXmXjU/k8n+70OAgweYQ9
oY2HShdONCMkN2v36skppVw7NGRP0nRJUbk0z1ZNvacp0dSLgz+gCs4pztit5Hls
KVYaVxkundHYi/d/JgbXFjjnHNs9QzZCmShwsHUKrlkTjehjtxsThNEqS3sGtsM2
A6xaPL0dQd+6HbNUjrdmDWF6CzCt9OqZpCdgy/noR4tnH+NH6T9LkHVEq6GhQzNI
j5Gwe0EOo3w8CLWmgWM54CDXjifAgOv73QcLlhayYkW1Cy8/C1kDV2ROPMruyEcD
U+r+UMCMTk7xDROe83ze3jWUtBYnUKHZmS2tWBS6Kf84I4ybZ1hiqropUQplIakq
glEcsBWHdgomsYqapi7wGtucbWHgxZiaYBSp1hfLXzkxvMGrokcFhdXKSuI/qNCJ
sm4BoEH4h2DfLKNgr3tMt0+MZsZgEcOhmzaoMS6heM7IHL/t/hi4S1v2oIRK/Etm
CXPnmckhI04r6fwzhLrGJls3ThFvPZ91rLmn96Ki0XHykm+9r/t1rpbMsQgB41l1
IsPZWfYy7jtNOQsgTRsIY2kHnVpf4beZeaCjIYznKvwTJpaaH1dJE/P8ZVAMLZGn
NSUkdNPG1nYrsllW7pz8SMzVZCXcADY3FUnsb1KjrMTtfzxwQUGhDTr/+T/OgDTj
skPqGZ20LcY6Ym4+iif4ne77ZTXgvAiMolYH3L1jPZhNtuN9yF61h/BRIIBG9EN3
Z9d5ULi1RBYrrCPAvWRWHDVh1oT+MK/JqA88vX149O/K1H6DZRCzKG5WFCxQ+M9H
JFTPcoWu39fMqm/kyGQbVflA6HPsON19dZwypQmSghZOpiAIXTvflscr1sw2k90i
Zgci1psYP97G2O2sGY9nVaXrMUS58OuKtCVj7qC5MCvkPeKXXPfgPNjtrvzcdQ1p
odAQEjTi9yeqQR1uBSiFWgpBEF1fEpirtnsSuWsmDBx5SuT3m83HnLY2uPP4AuNu
ObENhJFjlKkgq+ZIQNkh1CpM3KNDfJL6Cn5dw3D8QPnXInUmsaLygeOyE7EOd6UT
ZXBvAG6BasEzuSmWMW1Nx2tDn7M3LpcORM81xV3NYtSFTIHCaqtHu7NedUDkL3JT
KSPY5B80ymIgL5xi6O+3MGkW8eCT/eK6teBTxA6bj5biQK8iRsFtqrgDn0ol5CA0
7vAl/zSY/0ESXrN9hKqlTo0s97Hk5HI+UgJZ74n6IShqi9Xs3MbgkO5yVQlQVHdf
asw7YD4/zLslNArgND0UFm7axNsmi3o5nfH/Z2JCaHex+Zcst/XmfSAEU5q72uCx
mP4NFDdmUz6IVhpwzFU1uPSYqxxWSKWpxDppCuI6NmhkO5Z4P6WrJzGPhbyvl98p
vTIPw1hu6BzHMJGPJP3WFSAZn53GwBcTPaNtyLErCJWt/5rA3lTLuWiLaASqFdhR
jDWw18QriJPhid70Upd9IrvcxP2PitMmzd8cOONId2JgC5JzfV30+NRt3AUB+n5u
Hcc1tciuI82f3tWIokzswEWA11Me7JTovPJRtk97l1wMUvBxfb5qVoVwh3PE3SdI
gOezfRACTUJ/7g+TkVIbLpcsz2KMlJSrfvijtrDYWlGI9STWeBpTFJBJYdfW44qm
9nSY0GzQOQk44Jf6vKx6iOa7p4pm/nSNqMCvWjgLXZJUBmhSs4PGneQOKItDasjD
Tby4WTaC58/J4+G+9C4BDcnfBeNgo/WMlCxTkRC5qS02XdzaatD62zy4UlMw9XqT
a6WoZFOalu2qIMor3vKPRzfzTj8pkqp3yVO1HawdoNPLdGMCOgRDUk2UKuKok7HO
tJWH4qfnLrG7qq8TnQVccHxNQed4ogmHasYmRKCj4znjWfkxUq/aH6n1Cw1PleqX
`protect END_PROTECTED
