`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jV2cmRKoDLKMnag7K/IyeVaaaaCR+3Rnu5hc4lDPOFHnGkMGWKRAwSn59BHhYGGo
Opt2C2r/fH9wPdZbAOxiXMUaahbyP3QhhIVNMHq7nwQy4xv2DQzxdSgahcvg0Kyw
zP9xnwyTLzlBKA3VPHkrHTsz9YJRpXEwsEz+u/om0wRjr8gAtM0afi4z7Q6Arkzu
lQK4Lcbldv/+zMTrMYCKZlMTl/AgJy8MZNcWOQKPh/1aHPg8p9CdzdAI/4OIp8Lv
OX9Zly4KuGihZFWQ8F9x0YrgJROjh8gLiQUs8yNU2wck2Uboe/OP6xrWW9m9kMjI
wUy91QtWyS3Ove/6FwxDlsAZlvydxX2cYfTrO5lRoB9mSi7Rg6PruI5YmwAFVzv8
484viqfmnpCgpGX89e7cuKkNSKKH2pS8AUN8vZ8WYF1jjXAMwZRCjzPoyrcB/9mv
6RpwYDnvKpP2ktSSGtYkniyKIU8Vq5/ALe2GQKkKEw4JLg2gNs7r3QBvQGscdEY8
/woZ+HLtt+WBib6262VcmQQsEbTwer3+rhAeluaC1qv9AR29tn1rCVIuaZjL/UlT
lWq9pMpBQb4/ndaPKUjXM0ZQ4yzhJJWMdQ16tX1w1vY=
`protect END_PROTECTED
