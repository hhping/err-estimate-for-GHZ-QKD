`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0QY4SwZ0EW9QRY3Izn3AKZug7AZGi/k6RIcg/2JD2RYIVrD25dPTC/tHarsTc8m
X1yjuBN0CWhrkC0iiMzu+Twj3ok59XrnVhcxMk220h3gs8XX60SruTdXuv98W+Qf
orrT8NFRybPkZ6Z2czAUIa1tEyzMi6UzR+yNxg5g7ijD/Na61Ohr3CiC0C6s+wlh
OBxr3kQkaerTDHyVEsc01v36bjvfGGiM9dcS+Gks2rDzXgb9ZCGArPhtv62yu1yP
qY5Tt1HBRl4rC+1V2J1eqhVvZk94M3PE9hshiHxDdgKhaPZM9M3836KseDj/r8wO
BXFC5uVzuutYuivO/5+tuUswyGZAYg1UlRsfh0lzCso6eNcoqOFIx8taqNquQ86z
NcMh1Y73QuDad8jwT+GwQE1+DP7zS45eYzHfJh0Bz2NW9eNjoHzOd10GwszxAG6B
j1iYTBMI8GyZqXh0Ury2Xhvmj95AV+6oJwehcHI8Vx+GcdWDR5LithuDahE11dLT
IBOm8W5jW4etc4W4i9xDwFNBSc8OhUrscy5PEFbvqTs6Sx8FiHwUCXBxpFrzta1y
IIj7tNzyIob+cABL8FrFkocAwHY/4vACH0EGm5EE9TxvGbZ/w3UVv8mAI4e7d+jN
1cPTrlIbBYObkLeALUelbMexTR2fC6NAf6IZ+w5+lGGWOjILaSe2kqGziue3vPMx
ePooHyUMOtESWUCX0Esa2D67h3uXhTTuNFD9kThnFQ11iIkKs2nrFXxFrRJD4eqU
d1epcMz6vC7ijpGvD4QqQ6KZ/7jbNCV+ZBWwhfIBlW/o95H+qzNunDEkIGP5R2LL
DSpNAqv3FgWQTy2uq4FkgoTsc29Abg4ZpNeAT/B/2BYwdbwK/6WuHWvfy5Wy/4Qm
JqTC1dN1qcfMsBEa9SnIiWaySJd4hQ826u98bkkKVxtn8KXzDz9/xOndWcty4qen
ED64KfOq3dC0lb2htnjEAv2JK0fA3on5lwYjm8BsRDAV1WHxgkpUK5/tDMJWpyWz
`protect END_PROTECTED
