`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
toS7aXgpL+pUWFm3rQSaG2FYjHh+6A52jG9LaDN2kszkycIQg0sTyttLqtB08Sj/
CNCzPXjEPK6lboabajQW/1CWdMrTwoVnHOrRX4Y4VN56cBx3YsShjdL6o92GBW+e
vjovvO/qkuYVf0Ufs+y1VmK5KmGbJS3biw2a5I6nkbgwZb9AVUE22PkcDjTh8iak
0icyxGKeFHzdBSR1h1EwpuJsJmwLM6rq+HIqvvMv4RiFiUfnDUR9hnvpf+EBAnRK
YZJMVgNuAPzjiTCP5CfdYsZsMoqs3kc9mPu1xdEMvHSWrpNV3j29M+1+xlJpo4BT
ksDWlhOKxaPU3j3CPrXkNbOpYfnETNx0Bfvkk/GvgYADwUqgMmlPsS6CUrBz1rVc
HiXeyvnzERa6y2N/iL9snx/6tbp1beMNrmp3JIHJ8phC5EVtlX5YiRubw4N3heO/
IWWmQJuJlFst/ItDIp9UbwdLwrcirEHLR2whOgHdYNcRdnC4SNl7ufH6ElKYrtyc
MTKvTQ5/K8KfL+dV0Atmtn6jpqAdzsPBYtbDFihBjEymCpBEaRJEH3KVKU2OUCZa
kQIj8HnW+Dk99FpZPBkTaSqK3iZAOPskUiB+fuFU3q7Lh+HFzA6yWDVI+VNbipV4
CGFwBd6vgCK8+A85RSEGgJhE/B63mvSfsYF3XBJaXygl/LoC5L9HqukbInbIEIEc
8ai082ru+nKVD5ZcGyVqayz3diqHOQwdTqXxFpUr5JzwTzUeyEXOtA6xH26TGrZl
hrPCpv2s4dEKM8p2sKvFsu8+wsVhK+c5bFwmfnB+MmNNxCNdLo8a4WDmzz2NNTBp
ZQYyzVRQc+TeBTMCJbzB4G1p0oiCB7wkngzlM4T48S6PLGfemq90+S1yYl5l0wHy
h+9mBXaHxjStXNgTcSn574j5vQolgxue7KidkZsUqS0/PLIPCzlDyrN4zePysORQ
EzVeLWI59KNsbCk6x0yPcWZ4gw4JQFXUIeZmr5LTtVnq+JYW3EsFfAHJs23wVdYf
VrVTB9bPnoa/fA4y0u9qmaGq/wwI+83viP/Y3M4ns/PfabhJaCZrwL1ntXLxiEYd
oXECe+GRYoGqCgfONf5RITVJJQtr1nlwUwI+9ystnGkt/W105ELnPSouWaDjVgXT
EVO1oaN9zyOst6HNWHeypIz1kU8RfjFpzejXZiyvBHaW/2fFE6ideSKppGMXrU4+
H0uYT1bYrQkyN9UiSib4Zu5zsH6+J8YqnpwbFy3u7+vsfWupiRovwYMWPHv2y74C
zg5mMKUijoBbHy6h+nT5OTIWt1t677dXyRXG3UKqPiAunwtfvN1/2bq2b9J9hg1s
uyOucpfi/YOOtvFwZSnQLsht06eu+ozh6x6uYMpxLbcKAe8RW3mAzrJwkp4T0vjN
EOywpEEe8eQGHA0KMtnI1YS1MwSM/cxrZx8ckUfr2AB40Y+gsYo3YLQjMa4GTScV
Am8aR7qrXJRB8jcjGAEnU85dk3Zhd33+qMGJCE9fBIjoQlBYbEeLmpSWaiyt5EYa
AatT68wyxYZFMumbNXUP2o7jdYPt/35JBeCca/AX66sxaD/UA0kkJ27y23lODGnr
JgrEhpF4OWmy8yoESDBFvAAPwNq7D1ABLnFtzUv2MtFfxVEw+lSUQF5H99fg6IGG
AWyWMk3YnGOj6zJuS7pUR7iPeFwu5+oqgke3BeqP+i4+0/wv+h93X7TkI/5lPSuo
oLaXHtzJmUw96l9hEMO3NQ==
`protect END_PROTECTED
