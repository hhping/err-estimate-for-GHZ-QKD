`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVmpuOyPKtHl/CkaNCZtapIVL7cCJMySP8A/d7LoeR8TK5/VMO5p4k8BZESFhP1W
8F5fYCo/O5auJAVINN8Ox9KSeYWqNtgUpdITZzUhnmfm2lz3dHIOu3ambPL2g4FH
7GAMUY1FALDoByNdEnZvylNe37O0hHbEBmGR7maKJ9rZRBdnY/EdxmrLScViYguv
wgwlpEVQ1U009CyWDpEFXFCtb9ksPF0AW6TyNwP/0NnKvDsl4O3S/y8+Ex2LHSg4
GjWj35ZL7Tiq1UhzMdheAMRO9UZxT4kGFeJ82bnqpi9T6syb8WoT/dheZxVWLdk6
NZpdLkPVm70jkLpM98Ina3PYRGuqDGM2ePEYNKD16ec9PZSiZBTRv8ogVlJg9iwz
DDCLdOI/B7T+kiENlnMbI91Z+59h0T5gwvj2ARl/v+ok/vxA0EPPY00X6SLhkF1V
r5kUa2IKWurlObphuvWXFDV6lFEZ4bq3hvG+PQ35nrXOa6j9L/DIYM4skXXZjZnL
4K72FsJxAR9+YK01O3pZvFNNwBuhRYmehuGDf1y4GqrlPFAn2j127IPndAeASIi5
VD/TXgRhP211rmusACEfK1+vNAj10V6bAHLgQsQB6b7fOtSZMmVNn7/3s4AHFCFJ
8vByHNd5j747kN8fCd2934bjmcIkTr9Bf+PiLECbI0o=
`protect END_PROTECTED
