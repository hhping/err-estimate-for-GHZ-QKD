`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6oHv0T5dN4jdR3KBr2wwZ0qMAqsoXpTclPKYuSFAkU6EbXQJTJJnNqZYSyAWRSV
Va0S2OxFcnQu8NfZQiIhiMUbCjnnSl8FonC0N8LB8RwsYw1D9AD0aE7mVwhK5HCT
EtAAXk+UvHxCS4qq3c9dTStOu9ZG2GkdOiMSD+MiMLwsRMMo3z1oHT5//ME6kysn
SqGN43/b/iFW91AjQkscRCb1kqbQ4DJvymNOsu+ANdn1z3QVhAqSukRLPtbJT5Qn
d+mE354MH2EoGd0dmMogbmko5Bb7ISlQLeX3N/7gJ5UjeI2QmG1ouWM499pIwKgM
YQ78KcOwQhytaooBAnUXSLNj6/zNixpJcLW4dsy67JJwdQV4c3lj4kUTH/6ddR2E
Q5nUyfxGYYt4AmxsVSZ6Qg5/QUPhSyrKaVM1rV2vI9VjNbS1Bbfn373olZ982Dtm
pzLiOAF1Hh0np/HY59iFkGtQLicfP9PlL1LgL4HckkBh5vL0DCr8SJLFkxf9cUXo
ilV82dD3yom9kcr3czIKwDl8xs2gFkoCL9c/EpMVyVSuusUOlWKegUsFNvUI3FDS
lsfCZOD0L3oba6XV6NrkB1zYO/G9wB/eqfACjc2AntlLkjqrQ9C/6fRwejf3yxda
K9mmW+ByT7++tZq8RfOrMIziD6rskINITydQ11fpvHEKwrSAJIrnZphwnDLoWN7l
As58j4rPLhp+5shMNFgusy4UtMnW9gDmurnKAHzS6aPW7F0R7nisY+5SX2zZI2ss
kFlGIh8uYkUfGVDQ2Nlv/2JkSTFdNZ7ZjkfjiHc+NEJ8cbYW5djb8ocEqiovX2Ld
ZVc1DI5tbfIZzAYXZlvtyyrwL+KCZwSQ/oFEKB7xAUCHlCniKqnC9rY1WMyWTsR6
ZVJtZI3Eb7mLe7ui22mWQMLwLqieWy/L9zVzuN1dAj+Rxu2v/J69u4fjoXsjjMMV
sKFwO/PpSo2xfCxNr4U3WWZLxRcHlUntZG+c11yP+DNNw+8i2iE9M9pfD9sdqLS7
tXquxKvopT+qvY2OtSjyypvmOn1laLx2kVSr1/BrVUB0x8DIGdV1O4Jva4CWJXmE
OK/2BtZAi7DzgQqp4hF5qBtFfjd3GpzzNUKLB4q0LiEDJI4Oq80P/SRIasRrHJGK
YsuwxOCsxhXGLXj5rkE8FnhPPZF55+N+F7+aCoN7ZQ3HFXJMDInR1KvE5ClUtKp2
KP1ZvwzgeiBr7FAZr9oFdaLcTUdsKvDBHXdWd/7A+rZ5E97gokQdNmqaZzA01tCL
7f6htwzb5FMdicfWuFAFs3qg8AXxPamnAruO87kukYDrR9+nk1qXmNw0V86/hFTc
uCGjRz9Pz/qw2WAb8E4Vj22efrilu/uz4KEO7+0Q8QgO4HUS3Pz3zfM2xZnJra7R
loMpwObZwQIiQlq4Ouux3h0oXoXIffODpoCx2Fb31rLS4eI+BzIhxH2vV+qq2NJh
QfEqq0PkUanzrMghHDEHNTypr1H1PzzE0B+at+dbyZ5KKN+CMmOg7bESJME0TMGj
nl2djqK+159/5VsbKmYktesNfNNBOyhIxC+QXbvBD6PdXb4w/D6fp5gryISq0bwW
dOev94GyMsvuWpc60GBpYCiA4KZ/o2xHR3sr9VOXNx3cOPwq1FHZhi/0A7bg8LHq
G/w8Wgi5sjsZulN82Zwfjwzzzc9Gf7+Xrx6bKhX8hhGDtC/SRpJeujrgzHHxkMCm
ISH9wfsBVksk4AtceI4SVFBT03kM3JxBzJOxl/X5bjlOX6rsRzWU4Qx4ZQ149m7q
SdNoZm6Lh4WelfQ5qHtxwEcigDxyYYo7urTQ8vGWbBI=
`protect END_PROTECTED
