`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZmwnCCtKPmSjxI5BE3Pb42avHTI3HKt8raE6i4jKxUgQGvlvDR3Te05BD925srQe
POPXJsoaNbPWUPaWXoYPlR34N2GBiUR34RSh49YRSnn9ftoKVxDFwoVo4XYelZ6Z
SCLBvn/TjMLH60DouEZsSEi7uqEbFCD6Z4B3tALAA9GEQdWdI3AxNSTTJ8e1wJD8
j6Wo8MVe4tbxEpjZ62T6NWScxbPm0iv7mgeYK8cVj8q7nPrWWm9uEnP9WmYtCDKg
MMus9JjstAydc0voNyboKKjhiqh3k3ZxpZynBV+vZIBrwUm7g4WCQFBpzMa56wL6
cxI3zomt9z7/xt11AlomXEN+OODUSgjPFlR2JqjyXuiVSi2HltnrYM9kd2nbzvJH
hq3yxt52KcelOV5foNdR264hKomXohZB+lv6yoceGBYEKVcVKw8y2DG9xbM0Ppo1
itwAXT5Vd68wVG/ai8sbLhT3udOoFwOID2U+bpKN/DUNcsRAnPEtrYT0rEEBjbqZ
m5ltueh6JH6IkLuTTSw+Fg2yw5m4mZuSdz6iPjAuQcL6qMaB6UsQIl5yVvmxtcuj
B8IIu9L7ltPZwlZHw0+4lzd74VHjn737KkWkdCDd+ESQ3yWoWFroZ+K0cLmgyg8h
JKhsjKoD49PTs5FWkeoNu3Pbf6nnNOOpkVI/fQ1DDxCJyF4BrPq18+0ztPXI0u7j
TuLAr+9vq0OPSempZSR4MH12doHH4ir0e+vt+JuiY3tBnovNqTFdEzWYXqpCvwoD
VaWoIVjJm29QmcusbXhTT3Vv4NLkNfbHq/NC0nqTfvOrNVd2ANosNhEYW0uqYU9Z
SCCdNXoacI0Dqrw7bBEOha4v987e2mWdk5PqXhc4eNl8l0eGcniIZ/dZ6gDsRTID
Qxgx3JVXjTFAxvTYF0D7wmf+8TDrxdW0MuFYGUUEoKSbjawrFcmwk9Y9Zc1eNfMu
WCspa6quynVy0CZVot+n/gWRYNvsj1Y/QiqmrsBuYocr00V4qZxs/Mmh6EKy8K5e
nY3vFXWOg6P6fFriKK+UWnKTEpV49hGMu9OZYKpuj+M=
`protect END_PROTECTED
