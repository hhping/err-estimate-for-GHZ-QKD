`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7umqJU/HO180BUhEyPy5Kcq1jGT08ees5kp9ayn3iUKKQMx0aj05iDHcLTqWgFKu
zWKkzCH0yanwGG7JnjAYgahs5qCNgboKp/FxyAUm3waIm0F0QISbgR9acV4Zl4N/
CuwWelHd+XKmKlTEALlMaeNhqjEz8pT8CDTwHw9oDMeHO3Y2ARyB0xXaqa67REo0
i8Vnxp6toZ3tUbGT28OQeTIUhUH8R4EEBKvPn9OPzW4r/UPN2Ze/lf2bI9EbFaaT
zySweEPfeEdnS02jUoBasA63375WhH4dapZ4DZ2hVCB2Rdh8+UT+hxjSkBExuRaj
hnDowucllhlTglNO9+KaaaNs6yJqng2MZxg7fs1FNE3rRR/V4thOTZU9CFBo9xuf
+9m5CQs9RuZJYOBUaV2SNlsZxscsZaUvO7P5YQEJqBMuzStKgsx+WtOyl4tR1Gr7
Gf61eEpjRud3f/cNj7IiVPzehURCNmOOeQXnJopcJ40=
`protect END_PROTECTED
