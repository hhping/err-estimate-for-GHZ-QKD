`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/eL5CmEuaJ9USg4RXRlKa04MnglLinP/clivM5zvjFRvp5uPrTstZSHAq30wPyM
BCdR9N3zbze3MXn4SjyQxlRHFL9hSRnHgQNqXk4BB13MwIbz54xTPGs/xv3UprR6
HVy1JN8uqA8c8tROqX1aMCVQjpuwlDMuKIYd7JrtRwArg2KN6EZ0GjfKg0286B5D
heai7SqFn/M0XQALxTc/MBik2S4UTdTYaubnbojhVxwNIrLPy4nPc4JSSHvx1al/
XdtfzNFNysv+pm5xWl/sX8COMfMPPtAMCMDwdn9eqk1gm+GLRBqI/EA7LYUhMmK7
04R9FzRY12pOPAb70NRy5u0xcgOoWOeDiNcoEZy9NpxcMmebQGIJ+Poa3lT8mPEI
IoE2ti8kv/LMC3y321mOwtWI9Tl4Fe/8pylgrZfwYoBXi5YJNy1chuO/MXbDMG+o
S1vMKloKUwxCHNrWpCXB9dxYrowdOgruGOYYrUe1ExHBxzFLLmbhIu15fp0//sj9
o6UJvFEBjzItKpzK/2RcuU4AV3YpGFtBGtbhQefY6/V2W1l45VNOva4S0seG8Zgq
slsczKPN68nA2MuUCnP9kK44VtxjNr8pb4NBB/drseEBz3pJdMZtOQB9Eo+wmnf1
`protect END_PROTECTED
