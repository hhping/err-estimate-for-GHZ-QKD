`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZ/moF6CbA0CS3+BmsDzbZYkhzbf/3sZ9yuBLFNKZScF82GGmslzm0zdexI0CQVR
uGXPJhVXUz06F0p4qHtegTRFpfknmr7QM9G5CO/QB6AeCcG6Wg64ipvzXdOd6OHS
UHxGSJUdHfJ7EroLxkMZJvPNyPdOzDzvxWO/Rlz8C5d03rW6dCdOQmr04r/TAH1s
FFJDZmQ60/kcz4dkUzHD8V7ksmvA6lt2sL2b/xHGOK+vwM83DuN/RJiXRLRZW+VF
B0bOJ5E+0jKaDXZsQzUgZ88fUWiqpYjAjCnPtjx0ySPk6opF+e0k30iboSlg3ASS
8XlG/uKBxEKOJYSlwLju+BSxLVtlhGwAJbU0/3FQb70YR+NNCQxNlJFcSXjlLDti
8gwdIboLwFAn0wJR/bOk52rRAllJZPJhN4DPK3mWZpSuVbGmkvXFUK2EqW36etVb
kAgRvTRkmwvi1D9ilh3wLpWOjNzvYKfbn06UvRcWrx2hQHhTD11HwpL9TW2fdY5z
tp2uc2InKZ6NXrOEhtkbHFAqTE0IUscsKEZEnGXQb7iW0ubluiiHdSF+rzgSZTW7
KoUJEBIgKxkhO7+9PuQTwPOnxJAp4mbWogqnfGJL7eNDW/uuqI019oSGeb+mGFms
kx/Xf/HI0myXka7aSyH3VEl+7kn6hpdqwVPXUHqoePYloDMWWoSmo2xlYmR3Be+C
AqV90nm+UoB/UQ9OShcKRpzyke5a/XVggssZNc7pcEjXOuGBkB+rqKu3/hJbPX9e
cmWNuN9PrjBFzvwwiV/PRCUt3ptiHRrMMJ3X/J77z3w4PZI35hdmyU+pKyfF/MGK
/z/9OCoR1NYvB56762Aus32gZOIOHUvr9zHNX1jvwDMWS/GHo7n0VFFMxxCq3OtJ
NciHsJVYKSxIUfPa4q+JK7Vqu069EdFz03UiCC1O2axjtutnH3fhdWi0LNvktT//
UobbkT4VVgQx0X99DYJVG789xseZb98ZlAtXDBknwInZysrGBHtAXDZWYCFadIXp
G36NppG88eKlt6RsdpILKuBOJmv6v/7r/yAzS7EAowEVgCSqiUOjekJUW2Ape/Je
vkpu8kN5kxvS51qJ4s5iv46H4+HO194uZmQpNel/SZvbRMakkYoXqQG43UGr9Xi2
3k0zElcldI+rMJK+9ANL0yxVcUWxFSFm6cy2UsmGf1znGp3pt2XpFRsOag9OMOHB
linbhMUB/lBFB9RxbpGn2fYM7PUuvvryyrsvNU1zZx4dP0iSkH8ruedSQd7PzxMK
p7HmAFwylZ4B8ULv+sCmA6DQlieTEcI0qM9HoVyXwYAx609TCJBmWXHM6zVxhSeT
vJskCVjmnFWMpmZsGCsw4icBsZa3NE5Q9mxkPrpbFghbHKjoj5nmyRFPdsWtjV3W
pUw3hKVQyyB5Ph+Y5iic9jrIAByfS2/Cd9IZWQi3frCKI4HVBrlnkkI+ss0HMih3
742Tt/5FFavXho9hlxOW0uueGI0sZ1QEba7d+IUz7/lG5etODX8ltTJPvH3DKmFB
nvrz6THuOyrQHP72NI1uY8CuPZ68kRohwtj77jbCuM8=
`protect END_PROTECTED
