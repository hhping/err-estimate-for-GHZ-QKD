`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvFpBRvIfSHhxqDGb4pu+MsNado7N8+ROi9pU+PNLXQEy3j81nfY4V9ws1mQRbsM
uIcbAhB04kc34BTnVlDtWCt8ccGLg8sBs5SSHGxZxuH5gs7HOnNUzM2ga0O0luJh
AGilr+4P6//aZCkSxDO9CWmfsjrTEBhA7GnRncr6SJmD3AEgEKWH/3LzmlY1rakQ
N125U/oXZg1xpAbwvjsQ9qav60rk2d9xSnPXESy1RLEujB7uggfDIRLfPmq031Us
7lA9bqz4V698N4rmeV0SScsyzIrZD6OH1//M3tMQVACSw+uEj/adl6vYBa17wxC+
EUKTdTKuXYxtM3DiJ5SHycanZp+uxV0dtkRz4xmcDrGBe83NvB430yDTvuNaWP9q
XaC3vnW6+91fSjWAfC/TdWgvLaqlLOuofavf8hNHb2dUPDOMOFomUxV0po5TxMFJ
STZ9iLV7GcL7mte7vLrlv4Pbfn8ETdwgJFIbgmPMruA1uwfJ2GohJx1vdAX4bLkc
oqLtW9/U6TiT9LqR+QWb9/GecR6Ofcnottg4aXdxzzyWfrmspQJDFM3JKgMhu40a
3OCBqQRf3gn2ZBWQT6JkcZjHPHpm0ABO3z7GjELx4RGIzQWGeF+kvTgKH3yN8nyY
o1aQNdP9821LPmzNEETd0PZ/fsYSUWPTC/AL0tTaS/zARcGIlH4ERyjsM6PRWp+l
v/HGXJf1rhzOBf7p+OH+dTdkAdHZXF7QMzC2GJAdfXSgqp4Tcj6h4W3Oe0BttddB
wirVA7RFU8K2Dv9fiKyySdgwdur1CoayDzfJW6pbTZkMpAa3kKpF0SbymPAqKA8x
kePUPnmNPIm3j7JnYK4fYLOTRJZqxPVGAoX4U9wWizmwEjHQQQeqOe8JVOTS8+ut
WHxDs+kHZi+3wk7ZHozutT31YdOj5LpPgLknZeJZIdQzzODc/iim4IfLY/A/AMXW
FtNYOOXNG15g70mAlMERqfqDsiiIApITGTV5pMG0P/mAonXniMWSLvgYan6NLTVO
gupFwePBO81yuOkE3TPn9fqGIkh9b9y43/ogHeTl8ETLxSPywpru38xJvot/o61x
8F82KfRnatdMnSMO1hWSOe0ZBioIRw6KT7Y+0G5whsEZt7LSCvvUtWOeRwZ9L+6r
3oXYDJ9o6+CdWux7NkcB6vBnCwfa93vLHT/9+hdQ2bV4/3xGZXWlc9NEEJ5shRBR
8aUaKpiJ1GW0C8wlYx8UwbAMcuFrX+c/DNZnwGmoEivV5gdE99KsEnbLCqJy7G1v
WXsjPFyB9E1KEHW68ndYko3sz3YJZx47l/kGXYVFLLQj1y5UtkKVTQM/p1nftuac
AW5cFg+9rch5tMYwHZFt/3+cvPEf4kWnmP/2mhiNjxaohA00N1LKutwpXtQSv79E
99CRAb/YwiwRKoNzH4suTGZ12Vrjw5052d4zYktm+5FPhkQXpOx1GalvokffkqgD
A2h9Bhfr69eiCDR2/ALViDSjri7i/Xb3K77nzhsUz2nfI5Axy1XAfGeDUGbWWEER
jME2XKwKryJywYTUGAEIIeuUO4hH8anLX7hHwDy6WDH7wSHFF/HTKIyj4OQCw/WN
GUhdlrCs9vKrWAS7jmBhWqNbsatiR16/hjMgRCIeUSPZ1uFh3HV/4KuyRQ04x5yU
25hq8dpA8eJNcbrS3i5SGwQbnyFUBvZQpWz6O5h2s+Z9Vx8wbiiL+PdWJDo1MAI5
EazsN/dPYz7tb/g9xQytf8/WK0WqwSbcdncGUQu2Ld1sLzlua4WSqDLHFxiDC1/K
nbKgjFcP9bq8SX+xXf2jFLAj76uK2l+IE25GWX9+kXRvlTuXotWOO/4kGawweRRF
4Id+o/LAsRykY/ZcHPB7PEfYxeSpGrqOsDOoewPnjPIU9WY3Y4RFvLYKCAA8ZI+t
3Y9pqswFjfaey5Zl4G1bfEoMV9agUyfjaucXqcSIqQAMyJrOkrLQWtmm4LyHbsMY
uwlr8sM0xYodUj2EZnEDyjSWY+bx3xhRqX1Vm+IyN9g5PO1bLlGYHGiLPf7z2abB
6WJli0Vl0YaXXy2zzkk4GJMb7XTBEKXzn+Fu/dF61xh+LVN4zDYZazBCUEX+ONcQ
3qOG+78kVzoSOKAtJ2wa3vUST/E0EiPyvO+GHqmDv+1iGXAXlpjtLRq0rpj18vdS
1HaJYHyQJvEKOhdYLIfQaEzBLOtFSaeCQhplryVQ4WEfcmxpBCRre2M9oherWYRI
GgYYmm64hojUjcp0q14j70bfC5N33dgQnaozgYb6qkRr/rrGUlGPNgvM8mawnrSn
SltIDp1FHfL/ndNb5BWAiOam11VoFD3xkYvu3WSxIV5w1TMD+aP9PtRsGg0cDzy2
s5Ti7PMNVnFpluSar5UnHT3dU9oq5iHqBNZpa//YuRmfctJFWp5jxblNv4RaOdkB
1m+F03M6X0SSI2wb4jJ3FgT8sRuEyuwWNmEPn6fkNIHj88FFY7u4NoJsr3S/4XcC
eLwXbyqQHZYxvrxrlQXCjVjbEuRY1avbG+gWQMntA5VcIkN/PDb8HDALWNCeWIuW
tFp2TyhhdL5CFsKrV9Fg6/5gOfunaG1k3nOLACOv5QeLCA0tk4VQW31b5XgG/TIo
Fnm1yOgOAZXvN5/+2J0v/CGW2ih3DZmPB+mqxE9dROckU7FaQ1UiEYshXv2qecD8
6+O9/7aFp/JfQPBLzBlHdIIgO3F0LvK3zhiayEE5u4HXrgxEBCZ2pagUc233wKLX
x3lIf6BO+dzOTr1OyCdmI5WYgwZywa0xQhD7pwd7FfZII530yT5lLhI7j1j/sZUl
wr2vR4V1xGzqFYBYFTcHXsGpzP9AHlUglChB6zhwXeTR3QSsHehLjxFKBq/zw2y7
jBYpKYDUUSdGoJf6qsNsedmx1GrnTAOVcovnJD4erm20Ks/kFPK+PyFeRCXUJ7j2
Ah0njlHsLeHY/LP06lhlp9Jg65Svc6Kk+9+vClx4xPcpI5JzCJHIPcm8kp2zfBS2
jm5IpmFbQNa5op5hlG/OU9wGxjWpKY3HAs6ra3xqJcCdbrbHdcg5gkaIFTNwsmWM
O7phSvTMMGy6Mm1ndbgx7SVeBxEsribGuHwzSGY+Nc4bImgRxxmYF5Co9m6HXq1S
e8wiAAfHF6exURLa8Zaqv6hbJg4p/naMLXj5xNCAVZcfClDci7MehKOePPSut/1X
WoiLgbqliAhjzSbovbYUYoNERGCD8F0dIxee4Ua1S3BUg4YUZ8J4+VsElUba7XK9
Z3YxhhoGdSZb8e9sIWc16/oaP2M/FrAmbJeXczxnKmf1+mxLT5oqXg3DyQMvxPnS
2npRo6cFWXMUuTKYJw4Hinsn6fsX+LRe6pf6W/IixljM/RFBOGZqE62chc2JTj7Y
mLUcZN52G306s3bEvUbJ63l7n98VhNkZlhOK16UjN72hMdy93aRy4VnDOCJMEqYt
fwVYSfmuJD2T7jwx4iENhO2E2rMuiyhBdvGC2lnCfv54GsjG/8XHrpoPXpd8DjQc
t5dBn8x9MeL5N4Sjnp+5SwhDq2iNc4444SEMS4MdzS6dX5QgqNezP5gMrBbtUmCe
Z/7KJRnP/GKefaDVAcjzklnfoQuf+EsuTLiAqnWOMPJp8RjudctOHu6N4IhzacsA
/r/9cNbwX0oBFHxrD5gP7RDG79jhlmdkhWwYBTIu39l05nGH0X44tNskEMn/xIUq
rFDM9YVl5iAs/iZm2710n8aRilHE97hfW7XhOAwoP9UCCmgbIKAfe1RxW37m0wz3
ZVAR8OGqKeEQlid+3MxkdrQxQTnr3caV7KQp4mMu6rqBE8GVg8oQAHzPcnP9sVi+
LGrgdWVYVY+UdrNlmCWVYp5eyYtFj+y3+n64+YxfQ8KD+kRu7q8frRFYeUcso0fB
JDy673eDy2irDCZ9I5oaGJlTeqfS9PXAqnKV09LtQGoGA6zfNB1BA56QF0EtlIb8
4ItxpNq8S3bzvaoCkMOaJ8IKWGz9XoshIzPRdQTyMEOpAz/V0dtyksz5yDO+mGD8
xNn27iT8My5diHAUgbaYtXLAZQaXPi/hutrQzykzzDU9z0Cz9N2Mn79x9NQhPM7P
q7SMPOGLTW6RYh/2oqkncqutFRiOZ1xNOZZeWGYdj5MeriieJOWE7SfQeRTrBZqB
fZC404ImQkLJ5M7W91f8OFhGQPtOgFxSoJRnYMSORSjaEuwrtK9PvHSXQIj1u+oy
cr7GlH66Xm9VIbnpPKYrlMkU/MrsGYu4YEZLSk1sb9GkRVlJGG43b+Ejxb1LSNob
Mez5xeTF0KZIIBfHZHJ/RNr1guh9fss/oRfdz4m/ZfXlqu1DpLUZdoKl2rV9Hhdk
oY0G9ARAuiSY8pLmB5YQjWUCaj+NwhuT/lyE/BRuU7aNUey0UfySizEyTRAXFfnp
XCd7IP3BEw0TYT27h2AXV6gsgBzHYgV2mpATI2C2cRO+vv6ke0Ckp73MJxnHYQN7
CkxCM1IlzV8ZYHNl9zwn8v0Bkitm1eyFp++IkoDWe/Ft8dGzlrPn0AMGKrRIdqGE
+Lk0l5DYrilzXpb8fOMo59+k/K8zyvfYeYPiFbyjqwYXlun+RZ6IBwHrDsQVtIGy
6Jtt+bmaDxnLcBEk5U+tw/p1GTpJ2lXlifhODwJSOmY88tVNvk9eiyngH8tsDhQ3
GdtP31AmGwFHm9l8E44fq1wkpL+8IGUqwWS9M9KIMbuy6Ny2kcPY3MOrWACjHzt7
fDpvW8s3dro0l89vQHU70vimv/rC6MuCt+A3LXtBpZTNBMKJtObsCz4/ks6wCPPK
6ZPzQ8nRnEzeW0nq0P1d+Xy8SAYcebkAxJdXh3pvO0zTTvlk8i/lGo/T8UT8BGRz
DDxbpUu0D8+uC/IT6EHuq8Zvmhf5cFtIr5S4pH3Hf+8VSKTlNVBSZT+93WwkVjbC
t2YJjB5k1q7LXO3PqJjNZFchEb/waTqyT/L8iDu+Aqh4IE+musqALOn3+KdCPdMo
BHyIl9UqoNd97kKPAxyNizBSfIbkGqoJGRgqy6dLip4phZD9W51FjxFPCASa0ggr
u/nuw//YRxr5kSVV8ry7kol86d+8Hr+HDALwLXNaVbA8IFZlHdhwgwopK4Ya8zBO
JVYps/tf51wsbqR+NIeTz7fmLEswVK0s3mkkGcfVo1HuX5JsP/nrZYz82ulrn3/b
gp2Ivo7jGQQUFDjYsH4qKOt2zU42C7DOtVyqCLbdZ9BXDoCayjZvKcZIQjGoI7mN
/xPKT6GUI/bgOHjlFqJh673DoXTvgYJvWAEUBYG2gNHQwVYohmG/fgeD73Rw2L1p
4yB24CdyjtG6GiWQrH/vSeUctNI3hmkuit7rg2972ElRf3un6o2e1Db6n+Wj1b9x
vBDw1yP6sDvhQTvVFuqrNmkv99a/5Gjd7YXzD3zjl05fzi6AsqFmM/74JAZE/+Ul
FakM95lcbHLrdz+DYHT53zHt4CZe8GrxqqyWmGvp5TgQrYP9XOgcqQfTf92VSh8z
NIYfIBZ3DDY3ncl24gEYAZ6QxbqvGGWuYwDfYB5ykxhw3gQpwSrih3bl7MnGC2qT
1mVV227mhEO7u5o9eHIoMVxQLVELkYOy/ZXR4e0xBoPYRLzlPHb2jGjWqaSpvTdm
ZmdUhBIA7d2Y1gxIvy+IF9baEriGNyTNO3aXtBnxD226gEwEe3jITxa7cu03Q2rZ
F6/QLNYDjA5FR46y46yYtzcd3qaIT8NYKN9CdN3vIITSKGKr9saHWFMx8rjM+X2H
b60ZfbI68KMIQJWbymuHU8ae0iODMSDhdWJxf+EG8rFMxb6jtUyVwqlDM5m/uYT7
YkEgNyFx6CkXIH1SG1lR0Rv00ZBjD6MZSAmxUwuzZOQbq8plok5f0PdS24YZnI8U
NZ5GVvo8RhxGXc7WSLUljotRYpPPMe+Wc2t/wlibpS7JUjVwuDeFovDQfScFdt+9
SZOMFllzvYw6dl77X1+zgB1R0M4kF5QWzUdV0ypTFeKpR/+0JRWsM7Lo9PvJJO7r
Vsq9En85NiKn9T0EGpwdfTDSbeptFaIoWcxozHnttrMPNc+9HFaXi1Q8By9JWp9J
xMz3Rw7o+mL/aS+dMHX5fl4+eX6lIUZwzy2iadYuN9GohIWrtKCC8QgwHd3aCGQv
Ww8kF37xmdyuxWPhj2kIpW36h7KwNg0i4m5BDKhwFUrTHQiP598sQIMessVWVHad
T15Ejhu3Jhe1Aaql/S1BnNyQMiyGTyw3KiC9jODFpQVLID/lIFsnd1HoUxSilnhP
C3GqtVHDollTY/zkUqrvR4BW6kLXhbUBbiSkAgc+Uy+vXP3IyD8T6agIPFR16hYO
yglQkE2H/7VqI7h3N4zKL1iq82dEZTZGppTD87QJ18kR5k7GRsipu5KfbbLH+1FE
r2R1co9aPKLdTz3Y0fAxt6v+uqCnY6CiPvIVofslokj54SoPaRiKkz3HHExabXG4
3tpgnGqFycWISAOBC1ioUa5NV2+GG2YZdQ+a0vKmGbLeBaXbxnNj5P2XgSWZmk7M
cWjp4s2gprn+Ji5tpsUgHwZuKIsbDtJFmSg9SSRIazZsH99CEnr9es3LRqIOk/2G
Bcn2kcSuKIsMWiZTY8gcYkCm2m1sleqoe6BkHa978L+zVnO8EtzNJZv3i23J85kc
J68/Q7ZvPJWnR5rCMSgg/oseiBf67XJX8OmhP0UMf4qwVmbIAjK9qGSrwfZMuG05
gMM7lfbvMRrfPsF4Ya8nGpBP6KQfZK5RSNjbQjzIn0iEndUKJiihzZkXGjAohXC5
C27FJkT+8kayaCbTe7Y1c0SryYAXbHHYg98IihPD8GSCHQRGfRu49QkStbHN1+sl
HzXfNVi1rx5VNX68zEO0R3hgoxHXy2ayKK5cua6ilVGOL2MGKFb8lqGB6Xk1lBob
KL42UxxOhpZPlrBdEWrCQzfPrbakYpKVuIEMGd4H/wrxHReRIBI3fJxMY86DdxTA
P87EY6HGr+AcghBOEV9ejaXJTNkN4VdIcrpSmGSAv1aA7KOuFn3vAh03+yuTPqxG
Y/Une6SFcA1imU96IDZLHNqFGu64EN0/HBJaE6t7WERUDC4a9m9sQLmfUuEHnnVr
xj2momHVqHDG3TvgP+p6SiFHgn1VJlLN0hIXIWIqlwz4xSRE9leAlEcz/9oz7x95
l9UZ2QE9qE3jW1VRL2Aden6yEXlaazySE7orWxrbrKrB7y082kkUKVDZZaeNR9kg
sV0qQn02Xev0sEYFihPZmhU/KWMZ/4yFsinSzBTC3ahtjN3FOCHkwdPAahCoA2jC
lOEaoK3D2JZGUrsrEenjeIZ4Y5rC+JIpLm+g02EU7QRg9jc5JWJqC0xA3yRp7ty/
3ARQa8MGEDhU0Zrw2ClcSNE5xz5LYPM7EJAd7uQdmK/OemzIXt8aKtVV8XENYV6e
ywtxeq70OGTyeaaOn5yQddaItS56Isp+fXLON1q+8MIAY01mQLGfvxidSfW40HNG
wohyvBscjW3LDpNFT9LeTUsAPT5MWwOPUhSoXFz1wkSQnoxWkl3cSWGFU4HeGjIe
hnX7hOgKEogwrnm2BH6fC7Ok3l040JVIfN0b1rLcJXCsVVhDg41sLonF31ZWXoH1
CMHxe8y+JxtpMzWOpJmUTrEUYq9ZkHgIr4I9ErQjTlGQ3mZ5Fg0WwNk9fR8HEroF
jO9PKSCmi1Gld82Th0LI1HW2oy0kiO3LKDInGvwnHpvEYqnxzhIRdIvycdc7GrRZ
41+Q/053FWgRzf/NTU0kIbYPieJYUUf4T3CRIPlPb/PzwWhw0I1QvT1erqADhUuQ
lvr4xHnl73bJdJrBUa1JJR5IyMIljKdhUa6Yfc0xvfW3q/dRScT90qmK8/k4FcTs
H0B+F2hKRTNt6ePW/DtgGCzR63yonr0zncBWxNyx03PghiHBaSxQiwj4nmHZ49pq
tC/xdKWBs8RJL+T99/sDUE/9NLXZDLwu6si9TqNFnh4iqBXr0JXjF95o4OD4yWdt
EUq4g+89aPt7J+Klzay0iAiAjUzUIZP33s0XCnBOnehcxaiNqdutQdhzOlnm/g5W
3ykRg61p/3JWrW1LyZjPphKxG/nX2GKsGABt0SVtfIQoQnKcZ3l/ThhzKkRT/EK9
MAK20bbV0nF9MAzfrrxjkBFcGGnn6zbv5S/bK5HtCWDyWn09KmBMlevqZmTjUY/M
+UYEDIEa6IEj0xN9NnY/JsUGXDVmDHoCZhSUTrn3mMm+TBLr7XYL1KlWxCanD6Q6
Bm0Hn0p3wwi0YHriOL/h98glK18Bs6Oair3qmxHNztBLx3TKP4wDbC1DxB9Ysu68
5GmabN/WmrzScCzyaMGRgU0faMc8c8l9Tz8NXhSGh112SkMJq9qvOf9wAGZeIphW
jpMgQYEWqxU9BDpH1Zaz5AwfqN8EZ5Hv08hj1e3kruSJNvmt/oPg+gQzjcxL4ayk
5apbMQLXcU2o10/m75TQHFXcrkpyNpUN92norpsAVvlpHftKNV15eW7qirz5I15t
n0afbtrgHn6L057VtliaGBIHf/cLtxultN6t67zeLHMMGRvjbUcUhvtGjzibDGLo
UGsWS91aS7hlYu2Ybfy3RnePk9PoJnDZ0CI1TlTlBjMFTPTDV/rm0hZshHleKtsM
LljQ7Jomvr0SeP2/Pwz+BxC4S9x8s0fsQLbTvtfHC+iKeXzGrXDp4FQdBQGSWxcb
bXSsHD3fxx3sV8hNCzN9k31TddDDyhMxrL/FuIo1QSJYEf9ap7bI+ZEnyA4jenJy
pc3rFqdjFC98PDxe8xYIKb4ZlURKxPgOd6uAMN8GWKOduYWgRNx+gB9YRQy/C93d
9PfAq6A5PzBWWLE1T3Bm5ZsLHTTUOXNGVGiUJw4OIj+e23zeHcwGQLMg+rSXhFxS
U4dmuox1/4hpanI+iYwjTNqfO9tbsbOeVvFAeCLyXWwlEwwAitfoKg5tF6zUsn/j
LaK7EKY2HPnr+fGH74PQN0lWEQAkjO2Az45PooPGm7B8VeoXTLDpNfFSX/PvVlWe
GH96N2E5KZMylUJsYSRTKjPPUKHn+sa1wGdfm0YnZZeQass/8qQiCZZeNa+fE90X
3TE1p+peTgEFfNewdLbskwgig3TKgX7PNW+aAoBa7cfZ985FifYkXawpzisQsVJa
zmYQjRhMeDJ953MnQvlLt3KzVEqW5MUQD5xZqz6Zq7Z3zXkmK//NfJ6E3kMH3DpG
9Ahlg78gQMxQI3sDDQ8Dw3ZV7T8o8BGyPix7T2osHFHGdyIdRHzQ9slWLtOkDvIL
a8MRf48zD63pj/630bvk91tZtaOHbciqUGS4ZU7t8lMzxdAI3X/oBJZIeSA/hK2W
wkBxAT1+wxXY5rs+40Px3Xj0VP5nxYQ+g8v8vXU4anhGB52v5eZ4zeYBepSAr2Sb
p9lmujt2xK+Kx49Upwxz14QAIjKQaLsgiklIpfhH/LSVEPpCaUCSQ+qhKPQlnChA
g9zzKB9a8obEgcYWcq4TCTGlK9AnuyhBhuFVNrCASEZwZuvmyZA+/bSBjBcoannK
JK75sblIyS8FEi0S05flNnwUbCj44pWtH/JaIsdYoNzS0uZ4SrEsPetWxfOWkcr5
igCOPP5fUbsAI6VqqaRpGLm9HEYBre5M6nKBKqRxmh/LsqfMq64qKa/YLOtModqO
XK4QpowhbKRYSZhWWVWN9KcP62KSZKzW832Uhv6QRAe2slroqacGBY+HM0zZ6FEb
EGKN5ADbCHnARQ3zu9x1kKZZojCjER091IUhQwYnCO/UdJbXArSXRsE+agGuN6IA
QnzfFCuHpfHaXkYYEWWUmfFyV31O1rAl1ZP8a+WPzp8tZ+aHzonWgtVWPIJpCECF
3PQGy0fbdJ8CtqJckd8run5Z4+QKajadRb6eYvzF6sM5pRRA7L+naIKlmmVfdz0w
tMprFToZwzoBCDUsnj6afVJ0OLRUcp0Q7AIiGfyRpiIVmrKy/bqOBVZHsauFRdPM
AXpPmoB8qr7QMZW6pI7d4wWl9QregCbjpU10vVBGwbv0VQHvoyvO1SJRxWgTfP7N
GM6VWaBBfr+lZcIfrEASHKWmmBKE1iMIpdjeq5id/YnijPxH9v9OsnDpNubY/wkh
hYGEjn1MrMqLOHhpinJYZNUN/Gopz18gLXqeZ2vbx+pqiwl7gsm8C1gxnJkR1nqE
PGKtiL+dpYaARfOuKeFFIToD0NYz8XCaATtTzwgZgLQEiKEZRzbH62QEoGmdj44I
Eh0jYFDKMsPp6XRGVmIS1jiUDSvWVWdS1dh9I3ybkQgXKUvdMgejbk3B7eY+SSTg
MqnpaKLsEXYNBrZogu7D0dQFydIphSUKfMVx5MclX1nMjAYvMKiC2eEcxacoRAk/
ig/Dac/W5hy2cnmpMta3yPM3EmNHFlc8KcYipmwMMemVUAE6hIUMQiKm1K0QBND4
IkFgmlTBOpK35j73Y1M2+UHBn1h7PFGXVWBWrfjv/vUszOwKCmEPG8PWzER7QkhS
8zoRmsQhXjnvKUrdOj7P0HOeEJiw880YhBIOCXbapi1DUPi7M7LM9t0QAg1eeUP7
L/Qy4jWPrPxGdeyy+TaTmIVhilNcobyq16KrQn3Cv2vcak+wNA/wPxap0O3T6HKL
mVcLJ4egH+cwmI8VpWVE1Br/r/H4HhoBc8dzi8MH9E7J+8ENtJkegAaVq1aiZbXt
d3qHb15Zu8qHAGZRetFdHlqqxh/UtBibHbFfR/BygNPP9zGEFFXw8lS+XCUZtQmL
IQuiv4vOfZH6kA5qr+Sk7tmEBImvZ81UHEXsuheBYqMjDxzEfvzauolC95K7cmw6
0OGol1i+WIZNkZlH2/GazXBoFDpQ50f+maAEBZRTx8Y4tFW2hsmSUi/6OXNqpz7J
Dafi1eIu51iRtT/0O/SNnhrK43xkDNBW3fBqbGiDN1cMXSuvQQ+gMEZqMSpWYx/W
MsrRGBCEh2kKAyn7VM64l8iM9+RVJ43ihI3lxOrvesBmElqwYGK9NUvOyPSyuD58
4JcTyf1QDZzotilF0z+0tErO0wTiHUbW/m/LnG6qoXktrXJj/URajvqeUQP0t3cT
OrQHhqOGqYdpwdcfU4KnmItMnPM+HmIksN8KPtUUfwz/L6YRSVhRtgQhYarY0OEe
cDQWSMW3bw7M8bB6Lrk+l+vbDrILO74uuu0HNTsvtd/dUrLn8WjecHG2HVEoEe5j
7WMyaW5n+C50TH9HExvxEF04VXJPiKiIleFmnrRns21ha+8aKnT2ZE0BM1QKxlYP
sPoga4dc8hGzZAnUnD0bF+YGkad4SSDLFsI42pyEy/H/LRGxf6snc23W0rChI2Jv
/BDQa5w2wPMQDCKfcAMyD08EhhWO9xtobFtt6978dOnlWzJsvw7SLau1JTmfWHhV
pX0Inv5qE9FrGv6HlxpQ+tJIw44a5PaOdHgbnNRRAzd+mFdtZKSglCVyI+MJ2r3C
wPzQypWOgm0WqRaAkkQQjUVeEkR202M/VHCQLvRb9rVz3FoXiD7ZM2DU/nbG1orc
lU27PEkB8oVCDBwvf2hP2BlNf1xyWNICrT/C0xGKJZUdWp4la5ncpgpBs9mMXY3o
uwVcuC70YmLoMMJSfvwwWYdF0HrEgSZdmE4cbOnaABnwmu7Qg0jq4It3yBcpXox5
4RoUEyg4Z5jyenm6npNhtk15SIh7WHYpWMge1xIeUa1nuA00yGpuZOCok/bKdOZe
8c0E2B89obYAjxzp8cgNH1cdAuhOJirkEuW4pF6HlSv1F8aM8+MuuDd9svDX8hha
tCIr06wqZYKH8ZZ34T0VICWnxylkzeUn1Zfk4xV2D3R2DmOvB6G2L1teHbfCd8mj
tnnxU4+bHh+4kdt/YTQRrg6Ht4e4SVdPcXPb2l5/W9YCX0azK+KaNi0dMTf6Pc7G
ETlx4eROyDmfAyxLEBKK2L5idsi2ZzxSToRkS/Po6hXcEJ/TI/1VTKGzwGDx0SWf
GmbbiCqp3Rgzz1QYaGzo0fT1wXjKBLvNX5Bthu3Vse83FK7C0PoTOdZ/NLM8WZXf
lUuLBBqC/Aowkw5CNW8geJtOiaDYiJma6sChdaKH0hz3UEJici1LuTL6WbIDpdbr
SnmwimXNcaRRrJ62FBActyfvCRl7dn4EQMfq+iCN8J9MOuoEkhRR2KzBxXOH3Ztj
LOT9eVoEj8nV/cGodfxOHRyfpLM1QUvA1rjOSRikmxAp8+upmu+b8FExR/G9B8xT
5yPwB6oNs33yo3Nzxgv4JKMksc62izSmOoKdDjw9gTzMEtCa68pp8trDYHLZd9LV
SjlMsMiHY2V/4AFIXReY5AsXlXozqyPfG2Bxv5eN8lSxAR3cYUkmGtJk4LnMeWj3
uo7nck+wpbWRSfiDFaPvaeIktudpmHSIS4uDwLtTQTeAC5ZSLjyBHZh3Ftq/7uOU
j/MD911MeKjpBcXCMYjtJu4vwLmzGtnuzgzY2COpj2wH1+N63YfmNfoWLtYhrAgZ
rkdhfw0wmXpY2VLWsyn98AFnQPKhEJ4+joBmn0BMwnQAhYRJ0Yrji5rYiKElzqqO
WzJm7tOtjRqBzGKPEfXjvccnlgsut0F6G0XJDrBZjW7Rd8ibuPFmNAuQ1hDUHseG
cays2XClo+FjhrAU7dWaXcLj+dDQPiM/Ov6UTB/tE3P6WOHGRAW9q3blRZKlbaPx
AnfOSphwnQxNSAWSoit7wv9Es2KU5/ESKrPe9SiRmfWaToP7DLNRW9OFDZ1n02aJ
yX4//eniGqoQHRNT1zhZBtxbT9KqF0AgV8B+fkQmMwxc5n44U0uStPrSDvgMuyX1
nfjjuAXxzN8UmpzsTVY5jdS97UU3Vs4/Mg9DZp4yN12wXvWS9+1uyolwPQkw6dYB
PtwgEipk6gcMEH13TeW0jnfeD16XrQyP82Mm/Gn8sZ9pZM7fSFmCVTegOx52WCmI
Z/LyNm+mu886v3+cP0ltaypgAR9JZiG8eW+cnsyu+RptmBUZvDA97j8JT8h0rd++
atPzd6qj0F6nxfwUH1aO4oJLREJ5yLkFG/bN4TBOxUidNpTVlJWDNllNnnIh+G47
7FDCKC2hV8Gp7r1lbl7X+1mLftQUyjg7iYDUCJeAWueu/cKCMqjTxHLvX8RCXp4w
/1etCnu0lMTzTdLp2rNAxuLHw9kRdNgx1uO/zFscs1D6b2VvanU58Nr1X708tWMT
77ZRELCMAajk9TyIgE7TwM+pmKR6vjLePvZ/wAeCYesHrOXq1Zrx8pD+O1ABrzuv
rpu2SlmABBDl60zsQdjX7M7eHXecG64xHS+yU6lQ1mpSuK6uUfZCOyO8hx1BVSzy
tmC5fsRcxF/kaxUWr8biokAnIGj4VAFfIJOalp4IlqbeLey+sgrWuMRaRJndb5O0
4K/hk1XXtEyL/dObD0Ktc0S53MYZ3y697zAD367gOIN4Clf0QHjfbZRjOgxEbUBT
l1NbKcRVeNEAQPLltQXN8hFgXgj1YHLDy2Db4kQSjPW04KUgzgyEnt+0x4U1d2Y2
v25r66eu4IFFcpf0bVyhGzjff/y9BiNtpglJAP78NGwdKiDzjsmiAQ4dLdIVpquA
JH//vMgr+Zz5OCHPRNUsMx+NAi56aEDVM171GCfTbB84rc+pZB8gpR+ICjhXlRNs
ks4EV5Ww6VO+Asw1RksSmPSsZVRJ4Yupt3l041BZ3xebzX7whu2CIL6aCY2zlkdv
LgZ0pGRpu1naaMAB6tIaEhb7Jl8IAmzpvzBezN3cvmwm/yVnxchf2IFfvRObJN5a
mpaSOk5Nado1Q09fh7LJLZ9W+NNjntmci5vVDAfRTmf1Lp8a6+bdWp3bcFZJyMDA
t4f+XGwPyWZMiA0D3pWuu5X5IMgHBsozO05JZnAZiK2UOKlF1mC4RMdVlAO91KKa
PNzAxTIpNQGy5POjeiqSdEHSD5LszfOyQ2I34WoGDl+hzTNN+FigJipYhdldDHup
QpxK7dp889KukjaakRKIcAnGOXFiqwwe2voFra4wj4Sw04TuFxVomAkxN4EGPxPN
7nFsPYzhFJDKLgI/QY6k7zH94+uWbSdP7MnUfkilpY1Fu24f6qpP/UjPpFytxBNU
XQrU9i9bCCB2FRcxXcVefj4faQK+tr2S7QkY4EaCzE0/RxqOqZ/w9pVAvvsvesIz
Igt2y0KGYfgRgEtqQWr6Tpxasr1TMJpJlx/5R5EkD0XC6lUI/z1RmEBROw9I8LZ0
1xJMllY5Q36Y8SVvy0jHZPibX0mqar1wisx/W/uWRbCA2iPrhcnnd0Ed/xbxmHAY
Jo77TD6nSYptRyaAeIT+K07XtiNLJVFhbGqR9S9zWpY34SVuRQPUurLMRpSePvA4
ntK06cm88iPWtEy5bZIjrjX18QzJdFnylgj2nxWkod2VclTOHaNOEJWSjAsmWYcw
ojsdZ/4Y4pzR9pj3ORUVA1ey2sDGRw3goFZFXwWvd+l+09w6V0VJStxgxTca4aUj
uCc6Vm1COnYdJxgFC9jIb6baYQpFKKAS0+yAyd9CSG+Rcva2ItxIkDvRlUi1zaTB
09h9wON4WgixvGL/2HAQYMwRqhyqIF/aYRsxEjl50Agmpbud21J0bOa6e2tWhIap
1EXApEuMX75qzHBh0tuIBHhbQDXzP3X1y1CvdEYZsHRn/VqfkXkCOAEQeR05bTqy
j9G+UHIUdqsgytdkeumw8VdEVYpVA9RkZxNJpgI0Jb2nG6JqjsCq5rUZyEKGwegY
flbqcH0ZAdoxuCYzkrH5BRMEOXj0wa3fuB95x/L9m+VFpttNRbvHfiTZf6hDUix9
qMoM+kPf1VOpZMZ33ebVQ+8I4ETHLdH5ff6g69B7Q5HL9e3/IOuDOVuVcuf+AsWn
W7GmUOl5zw3L4FMNLdKVuuwrg/P9b9xXR0hvdDyEBXyn6zThAq0y7ix+djhL0B99
5r9LlUE1TO2Tv9NQLRVIiJQK5/1FEx+DDCuryfKfCc4WmtHYnees818H2vSUjz6Z
7WJTNaMJpMTN/SIfVToejiGbtyy90U1/z7ODPACuHux4gPIeOGQoin/2j6+Gxt/Q
wejO+EMQh4igbiNJanlXa7t5MZUZ4Dvb6wFtThkMsXbHCJhIsgqu116tfJ/+7mMD
iN0wS5bwMiMlI0ZI4RpdFReEmTG0rNbU2JtV4uP2du0ZhJUSsPMKTVVn5gqIhdyv
A0gGQJya6ElyHvBnyR5AgatVujwhx3+Qvlk/ATet0dporTZU6VBRsKQoZYYmDhvZ
CvwG3NIZGcQ9M3ub1slWST68GXbAhmvOSYjHPL4Wk07SSKbkXZcnN5jcpFCTT25O
86HL8cslsQNWh5mliuz5s2SGTQ2woJ7rVKSk0/JCUlIzkZ7r0SC5IqwwXpjTCtpL
PAWM+UM987OeXxBlf/WemNsJYg3HbOZtQT3udqZznOYB8VfsWhNcAN0ULbRYYmNp
M/YVjNnfBEjmcBs4D0xLzOjAv4Timroy9qGIFCZiFtq5l1P7BPg+lhVsVtjjmT3Y
hNFODgMoyjrWzjBhKr0lY2MOQKMWAlMBaD7q6pjWMcV+RPDQT5qqtDKO1ckwzh3p
ImKTL+BgfZRSw3nnABuxcMK31/a3yuHaFycU7GqY73qI0oSWP4vlDm7tnRKxVtF+
osxkXumZ06Er/LxnwbWK/9CMBbdX8bIJ5wiVRSsJ9wLiy5IumhpzUzFI7t9KurXM
2McieEkEsL/qO56pdidl8xSsIELesVOpIMJK9ZOVWfLpVGjwKlr/lHotdoL6gdIO
DtCkQqg4BgsdAghgE1dLyM18pU9KfA+Xwix+RY2qRsNJMpFs4YW5MRUQE1gK5kjo
C303dBTsmcMLU9eze7rAoLEJ/bjZNzn/4vi8FS9qZzQ11WfrobBXyiSq2Vl4jfOt
C+FUA4x3aJMM3xNMBNRzDS7tb1bhW0FaozTujw0J6123/c1N+JM2Gxs7bXArCqcl
oVo3IFcKkD6Goi42vCgtAGRJj6SFO7YPzo0ZzmNkyffYXPcVa4mQLp3gEFY7aK2V
k/OAiRr+xUtVV+VMHidRhicbNSWdR3qAxd/Q112xpX2BMPW/oF3DNQguFxlgqrAs
e4/BV/O3vmnrpU85F6dH2lI1LpQPZZkY8sw4DPRbJA08bf4Vlo80AkFGy99ghlX1
cRaaCJIFXMrBvn2WjBvmr4kXnZUnY0GUqR2zxC6SF/WQbOLucfhCUHd45OTi9pMc
k4pSlYjUKfw4cGP+Rj90Q+zqRSVnWeASq3aFYVRdpUapRu8g5qx8qpddhmwjKiGB
VqkRGPdzIjILs0EiKLBNXYrAWwomd2HSZuukqpZTbeJ81zgAtKJovL4OrlVoyzTC
AXg0/a4TKdnxGg4asBTrNw+liI1uXBNvYTy893bAwf/B9R0EBCsWM2VSSboLHllq
Uq+Op0mKZRSDNiXAIstI7UtxbT6FGBXxcwAR+qyStwyc0j5yWtgfScsAx5y1+0Pw
E/6PWEnS6lbqW8bhc6awdMEWC4HlG5N+/5+txdM+1Gn+8DyyTkCVr4t4jw83cTzk
kE538xS5ogPlLyDmfTR5/ZAZGSw0dM2520yIFpHoekc1s8Z4eHurg8VJGXHL97eX
76Cp94OEFY/j8OVhWs4CDgNgIb6LoCWyhBApPYvMaLpV3fSPrDAtG8oWKe/02/dn
t81kD0j6WLC8TkAEPEmpKe4m8qFyx2w/C8yTGE1/lqGfgRew/KSVmo9idLMVvIYv
z0Cq+vhkKPQZfjoldYJKp8uv4t1rqR+3Ta3h8CVC+B7eklwOubzaErNRrV1sni+n
TjCclw7VC6uFGIU1B98Rzqm8IPKHWbH9hdNnNHaQgw29/w3EW10we++NrtmxPyoe
/n9tB6PJqymhlAm19R0CZ17w6F0Pgp2N6VDuyMscVyTQLrmaGh5Yr+FCvrC22fBf
ykTOhIBxbQWaN5wqB2NKdjQ7b76A6Ph/F4aKK7t3O1WNejNi1ZRU5iLlAirJmQkh
uQZ+OnhNE8AOWYGymOTuJ15ZYhdvxZacKpSYz9fgwsjp8on3gBgSPnHeURqTEjZ0
YyHAa/9NIYpVS36NNAkuN5EmBdKQIMPphLwjVJo8d/0WXZOMhsgfLZ1iSgGoftXJ
m+e6FoXcL2V8khPsxkcpWYBAq9BJxA3kZG/HUsgShdtluslIkKCXnG0p9rNBajGa
Ggxdp64r3/O/Fjubsa4EidyOri7f0mb8pUhj7gp2pVEc4KqQS84ADZo8GR8XtIIX
pbV6h0/XC9Fp/qVg2jUbdgjJ+Hh7akpBGhOcbbt98Z070SKsnfL9QMjPtOOmo6Ed
s81xCoai0x+HYcjBB4Xw+pcQglpCNgOgsvoQJ/IMaNqqdOCgOsbgRmB2VzUF2SMH
cWLJPz84x9wBIccVF7W1aDyJWXX5uavanRqMM/Y+CCQAxnoelh3WlZ+9l0R49NYk
HH4wDIvxuirTw/7Zi6sjYZViK+uRWKDf6XkPQUhrKlrxQoTJeiIRx8ZBvuh4Rb31
yTsstMAEMx+57+UfEuP0FKqjPtVJu/RkweBkSVVqCMpedmF5s92FjSIBDYHv7Uby
QfVWbj2I9MBhreMiZzYPV/kaEaobE8pkZ57mubS4h+y13lHEQVel2BP0oWRYcwMj
ePnLxm+C8xvxBULiQoEE30tZtDKnEDwZG8y7AL1Zc8Lra/rjhvzin/c3XqWlOm8f
WGcV5Dom54GsTlgXOYJXf8KpVVxMQSh5WixdbjAbqqYtF1Sdy26jQF1jZchKUM8/
zst3cWd2Bg4d3Pelq9I3vEj7YYAWiMZF7/XtvFZcn0SbLp2zrn5T8BbeKgeljC9J
iUPIjJn+bxPyHaGwFytHFiRVek7ywIHYfdTkzjjKAsnsYS3vQWTiVW36sDnk6kvX
01le5amv+Xn6w93/TN9luJgOKRglXy8dgoWZzSYKkhjXdgSltg1RH7CVYUorckuU
h5YNuDoidP6FCWFisPxtorMIWQNPhqa0OGs8LE4kVtnS2ME8cTCrGUiQJ+KNYZhx
hX4LMKCjSyr1xDGpPCzUBPuEfHvaxSLLo4fTP0CUsvJk1R4ITSd+mZg/y9ORIzhb
j4DzyMjp4ixlEXW0vLQWJce004r5C7PxhNzzqP/De2/7MXLMMadD41ThpxQ61Gt1
pzIz4r8I+6QPN4aYSvxOStFmVVL310yPaNpIy4c/qXVaMhO0oC39UPq6wbLpIDOi
t6FUY09QlwidE989quuRdODDNeksShL98nHjpt+RefX4ibtuWSambWxMxDQlXSqc
qnCXVAUt2LMwHs9T8arUFNcyVuSSO5+a8Ws3xcgCyMWzh1t9s+OVGhyfcvS46E4n
Xm97fv0/KwMCLEA/l+x0elWQISvclpVq+y9KmwSYdNMmSTx1IKpW5vAAnkK9F8VG
oZKNNtKGOUuMdC9LewjffGygj8Q19IWjas91EdLZQtcpBR5j0G5L4OFWC3QgA0uN
TlPsiZiQdrhKgx7shXtVIZWhUNkY6MGhMXIZLqKrZHQLW+eBiew0EpNWu+T4jHqo
ffRg17sQspZpHlbjQPijdz9mevqdPnlvU6QUUe4txhm9AyPohn65npNnxYwGtKYN
6KF4oTDxWC6qBkZJvzt3aVTOsZEezGBUPAxFbausPX+UYndh3/CS8LQFBYI6Fgec
mNOEIY7i+MX/p7ztFLvXPNev4nztFi7OspKfYFxXLRM8FjfNZQLw04WSJBkMmxJ0
3U7jTeqBvSsK0O9r75SOwtvEZz+/5PRyvzXDo0uJ0pc8456L9vm9tU252Ig2EQUB
8QJAEHnCRFMwUKJwADXKVSELz0hMQzp7Xno1dKlpZ5jQsD4wxS3dTDA4g1jjQIQd
ayiZ/rF6Cob1DKHDrbnRLZeHDJPJoh1Xdr5p3VQ2tkZdwTSVLMRPYljcn7kjuriW
UjExjfr6xBb3J7x+dqTESfa7jc5AZiEXyt4gJV9zJn0yzqR4ioCVtJhBgRfWgWtG
W3Csz7xqldB5erQgADWPf6BnHtsWfNUanT2StyGj4LiA/wlFOqtKap0JFLCJ4eCT
GpJowrotV292kfIHQq0cpFQJjuXEVS2zolzDQCehPWv5TwopS/0Bjwgp9UsXFX7y
BFlIQL1FaRgFRnoKGQNjbJurMLRpkKhAwGNAjcybY0S7P+eIZT76D3clPaS5CtWy
VIkcViKj4DMQ/jpp70w+COG+NX86PTawnYWavg3uueBkJFi4+OABxT5xP+S/LeBX
2EhnPbaMGkxvF10riKgM2iFiMMRZXz7JzlP92zGeCaHgQd4LvIJIeGsXu75fG44t
I0tbh4bkQ4W/tIt2awoqA5w+ecn8Z5xR4Ml9S2RotHNAZrrkf03FFl3p6Bw4LSyl
Eiz/d88B9OCkDx3dMWmzCyHqSy4UMhf1TUbPtJeZWG3gyxvUAmR/+gTcq+QR5Xsa
Go70/wtaEkn2LadAYwkPEH/KJDC7ysFJIqQj6QVuVVkMxHMfTA152BdJjNoQ9JpW
J4e/cgGpNTQlML+cdEryXHDpOQ1jQG3TGVmyjK5N9TL2qHN/wsB3ym80BvPqdVdY
n5nUqKA48TgmvqKbCRqw6OjB4wMHQMhHeuVuHNPOGo/C1k3ni9RDkh9LnTLtuyYi
KEqNuj8EuuhwpZjUZeis9NSZ3pjFcf4JhY06ZChawkuBaqn/Fk8tPlfb02VqOO21
MoMGd4ymhvHxIC/h6Yi7D8Pe9GMGoQ4EMN/ytwkyAA6dvG0FGTIbDf/GlZ1+L6x4
mZOml1bsyQPoD81dIcXFCNsPKDkKyy/wC5H3fwDWEn48GhAPv6xOkhEEhczbQ5Kw
0vymuZ2pvMR1GQJMkPR9KVSVR7bYnWk+i0wDZ1okSFoLYZYPORzI3+GR9JRZYKg6
en6n+b/z5YgNmRvV57CY1Ib8aKufxqs6DZLZe31wsz0P+tNGeyw4SPQuxrJRv9aY
ZPQEl4LSD8BASdGKo8Pco0n28wnSJJITFz5VbKBtpN5BpCI7RZYDnmAUkdtfsWT6
obqLq3DO2LnkJFQob34SNJ8TMNW1IK2yjCrSEARHSRRmBEnX4R3zVlm4aNFTW1kK
XPBG7O9SASOcDrTvWKtWEZ2M5+q0+JFJ37zOzUvBn0f3F5x1eR/1JiNE8aMySj7q
c2VnGzladR8DGeaRSLKqWKHPGEcjUEpzEf4Y8xIJEG9odtWqkUK9oGlJ01xX5c9o
xln247odMSyZWf5L4s7oeK+tfvuPhMUDLFqS/YFCmR3MHOMtYgJDvmV8AkSf0PMM
lJzDBx5Zmhlpld8ZK73qhBYPoBx3OXcy5uvlbCpDm4r8dJtkdBBXWC4CoLwhzRgA
0Yv+Fb57Sbztv4h8x4no5S3pfx3d6xt5i7ygjvObK+q0+4u2hWao7/jib1UF9C9b
p+Kf9+W8AMxqwEpuDABEIuuRFsrq7dvxjLMPwKH/9ZRe18xQSlS1wp06xHfmOrHl
gDphkihFaOHfz1TflIQKXcDOGmipg7DkjbNKrDf9//2yWvZwbZGw7brpizzhtt7Y
y56h5ct3E+d3rbc0lkb0MQ0BVCUMmthTGvrWGz3UQ+Mgkkl2Jkxiid3rGLGNGygX
98Z/oQRk2D3qDPKMVs433LgCs1B+Jt0gSiTyOEgXpg2G2xC1h1JQ22dSYyLS6Ok2
aM6VaDfmaiSxY9/Of+krQvhYDy1Ovthnsu0v63JMNJLc7Ke16Xh6zd4fWBW+j8+U
wC1fXiBY4sj/8dqpiegeKETmVpDb/hFtB2JSfgBtn57532f0m0lFS2yybLU1cS0q
ILZR3F+v0/BEGpICfISpO3sjPxNNHrKXNg5Q5cDftX3hu72sNB5wTyHa4Pu3c50T
QmMj004ORG72wcXZTNjS9qzU7FD+La9wfh3iFMPyeeJ3iQ9bXgsUXHkAbSuEGG+o
lhvHJuumJlh7OJxFfkhH0XWPImQRRMUOpBfWkrX1WjRZ40VIU9h1IABR3fQMmPg8
FACoRLlV/beJbExEUmAPqK8MHCodJmlEbMMS+Xsx5hQVUrHJ86JcT0JtXqfvwdqA
eRp6ktkAePPSGnBue84KvM1L9Krl0oENi5sdXDgjFtYYkJVV556I29I5fWdliL74
RgwEMThOqOd07L+WhF/Tb5mR1zulszq/JjDxJjLFTRdlKhK2MGya4cK1I4rsNTwO
yXAcrTskBjXvOo4TdmQ4xuQQHl0cl9wastuLmNIRCFcdmtVLQsYuIhjAOXkuvzt4
jb1nVAMC+IOe+lgEtMBhHQWrYtAT+qLFc03d2T6H7PggKIeU3NpqnF8fLPZr8sh5
NQcX1pUBTftvoXgsZvHH2L03ZFJAWa+25D8/s9k5P5cDYUmb33emVXu+FhQ73dqR
Fmzvr7n4XrLuOVXjMJN8KDMhPT4Trre+vQ9aa7+DQ+L/aXjyWDV3xV/HBH6FsStM
+O5aVbzzX9qjsJyngUgJCbDjGbUlrSkmzejSBriIP3mtkOwJyB0fllcFL75BZ6r7
dZUQ1q0d73VSX2NB6X7PPFG5FxzaDpT22mcGmvyZ5jEgKImAhz+RrqihkISoA+7w
smVz/X6ug1cVLvuwvkT6pXWvXJXa+v2mJPC/uPZBtcDSZYoTcKpvxseswRHrm82l
DLX2GT3oavL3PMlCebA8ufJE8uRQb1CaRXv5axMkg1pN6WAC7RDlRHmiyiagHqNt
u51WudT+4U61O8sn/rIqbyhaJlSJK6Zm6ocgW8HqMMWNbXmKcSggBd8TSoVHstH8
/aUAincN1cRzC/8sXbmtCtB/UhIIjCX/NJB7Yl5DRCk+chtuzQHUjY1gdLnslcDa
ALIxAWynHrRICbURqE/wX10zVuxriBhhghxltbN+WUH/gh1VC2EuQeqmFm/+zvcu
s7eO6CdqkfhdTrB47hUosXgDwLtagtnC4GKHpPXYlJatjH5hd5LNkefMl7yLldVX
ShKPoV6F4P+AG1HLJjwb320rDszagu/Ch+1RvwwkxpiQb7mRr65Z4jJ6787zHhRC
sxeQ5i+SjoDcCMs0G4E26i+UguYz8Z+Fsfw8NLHdxsYZ4XAUcMDCMxPqapEdvt2i
v1cjT5mIPn4zlPlXirbfWh+p21xffquYLLZXTABWOmdcCRLDTe/6KPsWVK4T7BRi
1J+MBRgQ3KvBGxQvnjAbNzGoCXPvPmGcu7TZ2XpWHYDeoScormUwYcmuISa+bI7L
3mlUtOIwDt2QPsrXLuqDWhvGLlsKLizkCVWt/nHaVrqum5Dx+NMVGC6VV1PGO1EK
reNVDGEMyHwEEpGSFIOuRNuJe7k2OHnaf/QQAQ5m/kUN5K+yzyMGvRpa0zTaXB4u
aU/K2hiYrk/IMXGVF0fIPVoE4qffHTWpwHtcmtU/A8cvE/bO8OGsRm/a59cetEjj
XJblP6x7nUTwnbyDlXgunPPZDTsnM1ice/014dY8L9JNbqKOs/JprYN/ANoiRi7H
OKuvpPYtAaDDe0MZ0P9CAdV8lgPuXDR+OHP+akT980ym7oiWI+DBXZiIsw1GForj
QnHiiOkG6RPkjYkfZ7rMTbqphI6v9ggivBTb6nUP1P+CgSYfQySXC58uRmsgkvdu
vomQigVj+EqOt9QsoabyJx0sZJOsjNHdyDRcFwAgC7LcdtND7PP9OgOY6KyWA3WM
l5aCOu/opKKOjno7anO3lCJB1FQFyyBLbaJ3ProHPAuCm1DFLeJ8q7F05VVKhgB3
ITnO9u79dcw+85ayrkY9k5Jz2Vl+WnnC8A06Gh900zhZWY4Rhe6y3aA18dFKQ4h3
iE7waqPoukb+t+NjZ2jNzWHawZxERSe5+1fu24c9VPyvWEuMqn1GOjmZtWuzHDCs
fklXjC1lqXJpnMd2ie7Rkd6zvyrQqnIrncgoHKsIaJIaR028ZwhRQpbzTGXPcg1e
YKuyjcy91LWX8mL6vuZOpdFBWRTtskxUtECaT0BmPbvEXj3Sf4odYLuN6IgNv1J0
EYGF0uZwv/kTuNDkI1FHD8G1ySxfih/6yjntsPfebiRTiQnG24XtkdVL2oy3GcXM
BOejVCnml/SGShAclpVSqg+JNeHd3f+oKjx/S9I91KiLGzeTLvpmLyiSU53jZW/I
+jTOuu7itqvrWVnZzCD/oOru1ycX/wYQ8t/Dh97bGsx2FZeg2x3w9BybOiQwlEde
9mWzveNzq/EV3ovT+zySUzFOncOJjgFnwWGRjRfXyBfy5+JCOQAyaFQswDt2bYSU
cviWESII8LRx9hZqVMeVcWBZ8vfGkE1eoPQzb4pZYshyb2IKsK0Y5O0ahrNGNPWi
IjrqxtHqBUwHaQZXyNG1pJXwebqYOLwcjP3j2UuhFJHl5EpLhvKfLibz2rQ1mQu8
EaeTEStilpMPof5yOPvTY9JTMXJPb75cXg5r8jBVvIKa9y2Gu9g7tYtdtwrOK8PQ
NOEQxwol2rysf1XUlZ06F7gh61G0DIbp2+NMISrdibB/xGPwK346cG59WB3Jlp2h
YTLm6XF0M5IRAvBoj7kWaaG+So3RVBB2jqW2eIuVbSFqvPC+7ksOccC5sDVkykzG
/0Qr4oY4YeTw9H/v+ls7tEulS6cZV4/DLvahmoCsmGogmHheTHZEH+R+8cdPZhS/
uCrOv5UcGqzhojO1Vh7DX/XdndIO5th1GKVNkRlf9ibDwzB8aPpZUqDk2de+tNUC
OUwi89/7J4RbhL6x2q3gDTZIk6zyi8UmFgDqHMSQX7k9/tWXeqIVYELbwXApDaPp
Kawlby8ymlywcNPw1I7lIz08wAsEALDNDpntetoQyUZU4KZvd1BJTQ7qsN6r16dy
nRnvGc9hBEglSoAheFXgMc0i/7wqYCCVVEQqQINQdQ37eBtENWy3FwucFISPRf4u
ZwvgTYW3Gc/S4KQTeTafaIaTvcaMOGoExkMjBMYWBmZmogvi5KQtIgrSjHAiRe75
muMNCzt6I3XLnsLOmHskM9JvW5CqavZetbqpHWkLj/mN/pPq8xmIM3yt4OxTPaXW
JLj4wNRclfT0pJ4CntrAADWk3fcbQ6I19A/4lq3abnsNaRnUAXQdl76yDBbsfv8i
uTq70dtr41XtoO9PL6BMc1G+Yjow3GZ6rYG8A1myaGffOwSHabrtfZ7wYsPazWdI
DS7ZRe+nZZ/wiv8XzAMCj6/E9Ey5Ha240iN/1HC88CY8h7ejO2TfiipO0aHq42Fj
PflIgTN0AmHO+n+Nxjg5/WMgP31u05i7yg3LS/VUdhD37g42xhjIblXMMZJ2ZYFl
k1SXEQ/ORa3b22+HX3n7IJDEjiqEMdqxelU/gpmi8rmfhuv2xni9P337DX+sxrUK
7gA7m9W1zAPgoKiBQO+PNFYZVxOAjuA+b7APHk9hGgcMz6+K24NslaNDCoAjGiKn
AHPp+NSPgfV6Jxe1M6jN/8KXYhkfbIIU/uNRJaNdLvu9Vp2BI1mf0qKT3Ui023WB
xf+nNpexs0hJTziiS1JO6r81KqblpUeNjXe2qACMPXuF9aZD0IB1bu00sqfzM/Dt
3w+MpV0K6xWzQOKSs9ZqF4zALIlINmVKD8etevwso6bQVmuv5dKDER8xuQuu8qlE
TVb+gafAAm1YpDBwysxzaJ/ebANNcu3+jHnaZ5ILqGRqYbykcX+1AIksweI0n8hY
MgVOsTuVRdfXvtGcpaM4TKZNyU5z8tqyFBsR0VAUjAwiaNIVg7vOwAVscsukxziU
HWGIE0kLIKz1BhaPMALlzf5XPNohoUDp/2LvBQxTnlwtwIkX0rBTMMRnpoEJcyZ5
eYXjIFrvu3dzNhIxs90oVwDUSdpLKafNHuR/pOtv9TQAafkmYlaQCnzXaoiCXyMf
jn4WAMr7nbr3jDLnHJHQZofdHri0H90EuqM+n6+0irzCtQlE2cQyzziFor25rsXy
03PEp4W+6rtBncnCfDe5ST+Vr1BmpnS7LfkJQePYQtCx0vLUy8IRUpETHCWVvLXK
yLy9JlJx610JrENheb0f+s6nbu7YKjd+j773bqWPBMbxHYrWub/TY/1iGO5G7sdD
TDbZn0/NRipIZV2BVO7TivJvyQTiFvB6N+UQ/iYglhqbJru8Q3qXtDsGyo4pjzDZ
C87U3SPP+FsHF2oRcwHGViAzzQOgotahM/5gpvmNq367ZNjZGnvSzbwqLJmxXOPF
toI9qAltcvPc7iHb4LQzSgEmSQbtG8jfV31HOQx2kFNFGff5f2MiElGjDrv0pOjc
6cXINIGHXrARvo21vPzUbJJtm8EHBbUvO5XjH+wgwTPduMnFu2gwGFn0aGRgAVoY
ouGyYIdSQwteS1Um+83pufcQsL6DQeFTz3cTj9XI9smOsjib66kYEZXhXQ6PwEq5
kUGHRo4vjrBiXT6lbIb4T6jYaWfcLDqnI97bzsp3Pa5jH2SK+yBjdPXTZiJhCu2J
xxZv6/ZuPW7CX6v8yYN8TWgIho5PWp7i7Cly040w357tHDDpdb+Ab5gwMgnDDK2E
jcClx+EdMHSty/uj0ibnh/Isyl2AgkW4ukQTLZt3xXlfQabby36lGffEIT+0bXnS
SxZ0dO/Ks+FpGHQP0JRreenx4v60ZatS9dUAd198XaC7JIGY19VEJRQ09lNpvTTT
i3WvcUpfAT6AsubW2XSV/GGWo3Mc+sp2pTo9mR1SshxKTQnobUSwhwnS9pbIk+uO
S/jXK8m7FDsJu7SqdsgDws5DX52BlW4+fKe2dY2ME3nmHmoXEFeCy3nBlrwZPQl9
V6gYpEIawCv408AdnsMlQxhOyKeI9XDU+fB5IImlcIfVCNyYLyhacfjUktaisuDE
W86i6FCiv59UsuTD9mTw8FD8pXs6Jyzz8IoNxZDfSfayDxOMS6iHvZGJREh1p8xK
245luID0w8VrBIu8nvpwnBjly4OBT/OTDmuOxEqSR0ibWu5AR9+0Kq9ZzuYYbiwj
UpVDoNKZtxHkzNoMMij5RxdTV/mVQPkxOreq1WdqBfzebUPqUhux5Cd+Luxswjv1
qTAt8aA7LQC07cdS0ZkEXZl8g6KwPPMF55VI2a0Qocl6k4lqj99Z1fEkSSZhhrcZ
Bf7XpTOyQJfaOZBJBMQ/SXC7o0es6B84Kj7fia20u14lwos4yNh1EUcPYtn42RWM
tV3cDlYTazUVBPxVKCZcdvTrWgBgeNLVs/IyX2Nx2uBLBuNQpNmdDRGGyQl0M4K9
tpVvBcF4GmGOp51s0rWYBkTd/WqwYiTp07DMDt8+rmhKPqwYoDJJr2Z1XIPJWbrN
s4K3G4DE4gMxpGepDdqpreu8HDmSbwaG29yGerwasqDU0sNm5r8G16U2UcjY+n8h
LhpibF/Qxx16vZpShAz+OCslz9KbMyetGeEoe+j3IQwhBttZV4CZWXkD6Ru7HWLN
bQdOOox/fp3ZsfBCmZILG/EijCGCySDr3dnJZuD+s7+WLglFDh6OwwBGcu2xPJBT
XUw5jC+vVwMdqnhzZoVvjnsGdPmTBCPH2qht01dwR2bjtD02YyVjv5V7ZZ4hRjdu
Z9hpmJK/7YtSSXbU47zhFPf5Mrbz2eOJb2IR6UKoPHsgQDhFw0zUyvD6WcGhbiKQ
Tcr9osplLyspD6irBA1qeWll3Xc1LIbbZS+79EaF25dx2CEE964g3fNjuA3tPMCk
0po/YT08PQREIxJFOrDX87+3dpCMjV6wwgOX4y3uGgRVu/6IRITe9vpgBtM67D2S
+py0gau/0cLW7n0L3PRiXHGVYq+VCRf0FmgEiOIN5ts5w3bs3m1nq0vlP2+shbQA
eAuZ4L4IrU5dBUua+yaec09xBduJ4PO93HmJF3CBaSxbyLTrWJ2TPNTxGr6BGHYi
edCC+5+mWKRnM2A96boc2QJ7XtN8ffs91Gk7jjUw1tAeWBa/tgQSM3eeucr3/fCS
fvgdGo71ikKdcfTk7XiN9oqcNpLhx5k4tE7YRjSrk4OssQDjfYGcC+Sbn/yh9Cyt
ZFD7G4Sq9WN+3wfd+a3fD/WM7bV8A3pRXFKTYODm4iI0RUXtmCCrvGVohoh/uVj0
esM4ITJZ/UQPZX2QMomseKIoPtsrK7RZixZj3W3dpKfsvHv5FTsoyvmh5rkjIpVj
B51LX6s7pnJb026gL0+xgPGol1zhu4Kr9Pa94tTSqTOuX5MAI49FSonpP5fhdD26
ospoFKyK9NJ9lGxptvFRBh/X0XZxopg2l9c8Q9pw3bKNdEp7gcwPuefStVfKKg8j
wkosqtadJBf5UT97Qr45H9NHAH/oft9Tql9XVWQJaU8908ld4VQHQ+VTNOMU6f/G
xU9LnKFLa+BHoRD7Y22XhENhDKK9BFHlDFuIk0oKl2Xdx2C9KppbS+SSZ6iOGrHP
3tjj1JoQq6srGK8dNEaoMSmpSydZrjAPwWNCHwaaRhSbuwvW3uK31qchFqfDSVko
mBQ6GyVKcI037DTAVk8CCFSscz50nQtmTBOonVJ6yB6qog/MmypGZOALokhyUajp
LG2Wwhsp+s/nSy8gkMIpZJV/1rH7hkixJic4DyrjkEc8E52peJOQrqsn5On3YHh6
jJ9cPdVvd07Xh5u9TtamMezpOyRs0smmmZ9ULdMREkODD9CelOKFPttcdUCQTOwu
A1Nvb2PFErZzbOGa1n0v1tWmyf7Z2yXJBFDxzk/qb6rdIO2A+OC7ph8cOZrZTae8
Kn9wq9M9pdGt9gw6Nq1OXjZa8CBkWmhLAgz8pK47lorR6j/meLbcUdhsRCTthXDb
VF0BN1xiDi1mTiV9nYpYYvz+jtxQo135Xj+NorLOSETd0ktZ/U+cdZSvPU8pbEyM
qV6oYEIUrzhPFRWlOp1RlyNriZxTyRR66nSwtZSkwujJ826khVHXXTlEaGp6rbZl
J2o4YoUz7x2gJc4Nsi1lQ0zDcG5juxCnEZN1qhdU2nC8BAJmsJgJj7LfeYqn0CxP
HgjB6Q3QyCkqgxbYF3WT+tpmWj1FfrrvFodvblM0hHgX4wZoR0oTd2jwiGIQCTcd
URwo6AHwC6yxFgnF7ABSh8cW9myuH6188eAj7NDmk06y/jYfLCRaikUQbZK+XjOz
h7wXvb55Ffsa9Tx79NXSQM1EoapU85yC0FQHiuP1DC13rQf1lGlc0LJ+dkBJFEY0
bkuUdYvIrQqmpV5muxV1/UoNpeTxCqevqdMzbk8UEkwsaqpBWtojGpz32jriyHxh
RDL2eA/kgk22eV6ZRkesggYdtsKdi9HwrzDXUVqcHYFuEMDxzl8Y2SpJSTQWSDCQ
KDRTtR6clGBuU60KRXB4i8+7mfpfcbPGDOxOa0uY1nvOS+IY2h/4VaR/HMybLvUp
u05JbpQegkC3Qj2yBXlDeKGzLcRrhJGXduNU5t4cpRE9/7ChLCWd1ZF6ghW7H3W6
vXRTkjX3VU2N6eOBDRTLd3IsmER7bf9BEcMmRWFsvOQmtHhz49h5wipt8LhrdhQp
+hEyliGu71QWzP70I1FSXdauarscvML2W5BNifT7EYdhwlcSjjOdlerpH4neNgqO
fPwpmZVX1iyaI1ni7O10qZ7lbTGbzyoZUn0qgenz46BGodLKixgnF0nMsEDX30AR
DlUNo/7bF6PaL+8MrDaWXg+QxWtojMJN6O56oWSGrVxUAiSPvOSPYI8EGbjcJbyi
1Z703VIg/E8FPdSG0LC/htgoWkkvUGPQxOdvNnpKjcSJ23T7So97XQNtw/LBvDxb
pteCCMnl3wdxwcliuFK6aFMQTiVdrWRdsqVWJKhVInKZNGzD4+WxI7e6pGUIsv+U
21U7SZNhzPgJtGLN8KjdbcQYwk3R3p7jl//SDUkqCl2ebOwcW1njZxGRcP02PIS/
q8Uu15NdlgsVVgsPhRQzDrRiG220I8YrurCWLZhS7B/DW3yhEke0OaUdW4RNQnI3
9r7gscfRhMGdhqs7ELlw3pTLH9IeuYgRdG0Z9kiPXrIRAjUw3L3H3tmBnnfbplHI
RsDGZSMyw+FJD8AFfHgpmxscIvTUufByRmyk0SbfXMPHRBjhLLqZ6aDG9ceEOhDG
tc/Mv2PrbVGeX0JdAu5/r+Cg67iu5ndv62Bdj3ZsT/ybjuPv6hbOLQPlGAq5Z4mM
CbJopIMuD19M92+YlFXdpnP+yj2XUfgBg+L9ja2VOoS3lyKaTSeTtKg2PFjnOeDO
yW3KxfpybCPvkWy13Q7VR8Gi3oM2n+1tnKkoYQIj/sPJqBvaGB9f5lHZmMVBXidB
ztZvwXJdv9FjgTNwprwono4TlIJCsDWiQYxh5tgkVK6sAmtVpFFKoG6lA6sgSMJf
HA8rvMUQcqJAyAukJ/AmTJc0XcDIRkjk1vDyf4mY6dp5uHUEBJiXm/BITXuf9/Lw
h+l8gYh2tBAkXgunquHvHuTIPVZuvnnvkXpnJTIztsTSG46eelSWZ6zkxgGFg4xE
KyLTID3UO+W4LbS9Roqt/PJL2LImBgjkfRebIYqqvZgQ7f1wo2kMWwwij+p5/Gd6
0epByR5LAsWcxxVkKoiO6/qvCI9qLJqkpdR0bDvo3luiNIkgoWdr92PAfoUOQodH
ijP0qF3FKLnRI5slMP/8oAckrnEqorru8rcsotE/O+OZ/8DOeWPVzL4YYUny4gV/
80zKzd7gHUXPtQL3y57jLwPT05SARVcvZCydaHw8AQTYmJpoO494wGE5Eoa0o/Zb
ii1wY1OZvEO75DzTCXloeone+vT3XQIRz8KZ39JQXJCTaJldYuHXzr9EmkkN6C8k
+OsXknjOGmn4H6PAg00Tksk26dC4IpgCxdaVzb88plv4xqufKRQ2cyl4vrU4K0h0
9AXIgbfxu3HowimZEroaNr4DMG+xlRisOK9Bru4Gx+dCQJSlg260Fbc082MoRn83
gDEMEUZUyvGV3OB/AT8KWjBP2pNv2zTZGKKcYHBx1aGBlvny26iEp43JS5NecHer
rYYMWZMdBJmpxL42LiMDx8yHpuyKxC4rawXJOVlfgLFTBmb5F2B2K82n7O+eMlmv
xD3vz/eu/1F6dHM39TX5ujg+BIa/1vgJSedPFqaAyAoC0RbM2jzNiUVGm5jtB+V6
bWtPqnOoRs7psqr6u4IGcILeCO7VGBlkbwAbQ3QiTVaaSm5zHesPzS3cep7Uxswm
5z+2Sr9yS9IY45mBGxAIhm+aS4UDv/2/UoRlD3c+OZIYodHrOccDOoE0pz1YE7c+
oI/ItV02wx56RdYLC62DVTlJ8EXtTOKBKQS28tIqTgV3FwRhlvKFOJXEbDLlRRog
HaLb01r0dE+16s/aAbTH+6en1xZ69yGmjlhQ6w5GZ6wogkhsZTAEXYvCnU/JRPXZ
NrUzz7iQh9H50fjWYv18RsP41VPshHRrxVEwGuTK+272WhS4yriYSZzUzLt+Cjq6
mXayPM2fTgy+iMe0QWCydHViJWhJSWDeOyi+HDNy+wQ4S7b48ECaa5qDiHGP9SSq
UbmVFrs2Vz6n/uTFOEvJpi6MR1ZB2yje79Q15424v0bOZRYaQFtSsys4b7f2Wbh0
6Qe75Ug/SJQSooqe0XnPjJBXiL7yrr3UZsEIpUqRUR2V6RW3WofTk62VsfmX4aPm
P1YtoFKs5/UZiXCrVksQK2Aol9XlKfx65gGXdTMj+eHr+/XxEj3HeBd2Nqg2v3qa
ItDE25UgbJtKvzskAwSoCDHF+LoP6ppugzuDpAoVlFjb84/mQjHSRUtfFK0OA8+3
nUyUXhJe/2pWoo7vObUYjfTAz0303QadVCFpZ45tBpW3nas78/Jy90JCj2xm/vFW
B7x3mKdpxjkQiBs8uJ61dxviknXz3jvO1nLnX85AdbPu3JZ8o9bru91V9RnuB5GJ
pcV9+/w9PBUzpPt9UBufjJgLfrolHkGbk6F4KqFM9SFhaE9U+x/FCLvP1k1yI7oJ
bPLDNB34KZKHxX80M0RkwbqBCIRVwVR9PGT2YoHLKJ4mRIQdnLxWavH7SIsn91Mj
GWZ8TFZ+XooQ5w+O1Uz5DQk5aIcpdtqfMxFxc4vd4a7ArSHuyp1347qBvHmrKSG/
8STYRH4j/gEZUbi4gcwoorah4Lrv10b5/JBWB0zrO06+X6iya4FU3bvefEHUYFfT
0jyURsmLJDB8VReAypnjIlWJUvTQHIPc7Qm4YOrKp4OMwA1+y+ezK3IGCapl/ykk
F6L22XkfE07dN357KoBRhX6R1sth/edpxAS2UdVSFFE5DbV/ifZOoY1EfaShTCG/
OfrFFjKJTs9HRBi6g8iy48V7IE/EYrEMiJW4lIOwEcRrrJ3uuIB5KLX5WFq6+PJ0
vw8rGB9w59nmGqf1piNiklHSf1a7W1EvwGpttHfT+7+xZI3vGKrcH/tYN/plw/4M
qH5y4C3mc7i40htVC140LT5YpNx+dCmxFiND3Tq/bl7jWwzrhgvv8tQns9oTR3Q8
shdP+KTl6jZI4cAhJswC2nk29sRROQoF5nMC1FNgs24MXVu8mIJcmWRzyi0P2QrI
qEzC169WYp7iFBMjSNfnb4SAjcsT+71JUzJMKhIZk6LwHgozCnxSHw6AwRsfhm6I
ZfPJNPBL4sEQb7dLLCzSTxAfZOT29J4tSEeo7ym5CVmFbo7rNtKtyh8upzeu0f3r
o5d3bnsXDVw1zCBKPF281L+ZXZKGuwBcqHxk9mXeuRuozylF21bxaIzA9wV4SILh
bHWbvt0qifUydfukZJxya/tiy0btqqkAO6MhXZ6DZXVV/9IZsBA8VHFWvxw4JgoG
6gQAICSA7gG8Sc3l9Q7cYGZvfGG0TT26SuKUdAf7DG4JTRfBxynjoN3/rX3UCSwu
AaIxo+6HJMrswOnghqUVh0LpHGG5iufBoMRp1ZOl9CW2lfc5MYksHTrAOXX86oz7
Qm6f/OTNIfJHtt8sIis5tHVt24Q7y5KMSWNs9D/U8bdp479Te2W+aCpXrkIEsikI
oktnVspR4IrSaSatSRO5Ar9gMxnCymn7sReYqFi75DU3WZd8L4uP3l7P47metY8M
Rt/D3erWzVE13nUWoxZgMBw5vRkAnIdsIFAweO57VCAgza8c8lZq3pgMYlx4SXSz
qaNBENntOay3mWKpNG9O8tVJ15JnEHDz4x1SiTtYTwC4ux+4ZFT87+xhQDhK8Ohl
SbLprRCNIUGgxrKoJfg+BrkdE0EqImXeKzCX+96nWTzX+zj9gVNq6A71QGUvy49s
M7EWKdFIlDWQ82eCdY2kblULqu9Ait09Y7Tp0MXeHlq7YMYbt2v27IOhRWvIG4pM
cJuRGQqawB0HV4uHRrCILRLWSA3+G/z42CxBJopByta9WUudgAos9F9VOf2OlWY4
Lh1eA03ztMYsRK2VyY3rVkhjp0EVEHioDZ+1jWRa9yMWAH2/1/8UFiAKtwXt2yWN
U065ewN6yuf194R3KNhP7Wsbc5Cds9hfzIZsTQvH0EJ20DC++V5c0GkX+GxTthPw
5xCcuteGYzwxnpaCaGLAdpeuws0fQMvbZSdtwtIYaJM/p6kkIkXjgDkTTQk/9jtT
53TQW1In9V9dN/81WNq56OKBRguYq9GuLH83HaRRvMi5pSC2T7LZC5bAsuD0/moh
G/KJr54xYD8miGeUZaQmQkj3GewF4wqtoQKFWIwWcbS3dIe/QvavK27cZekUBhAK
pIU0GaOwrVYQRnP+DNhLC5u5pfqnANTXTXcRyQShrXoKXTMcMdikEhFfLvQWP/qr
/rmAusfb9ol6+QARZh5XzoD7TkrwOlWw10j0lhBP8LJxX//Rc72DVTITCB36bfd2
Dgn8631uVXuxjRQCuPiYcKaBlMd5xk8w/an90hrjldaqVNfzoR2YIunB14Dal9eg
MVf9S8iL4Z9PaaDtrCIHe6XyIlDl6pRx1tkffxdzjnUiCnztBf7qgwU/mUsR2FC7
kZeE3DAm0eeVYPWmem6HgLaJLKGH74zlmQmz3V/L1Def46chi6WInk4LOwIMr8Q2
ZvWXYtZIOxAmnpA4S1alr6Iv+BFXSf8AqkDSlZMhztwE9fcuNxmZ4/wT1/UTcvyi
pyUEIVxtVsYOeR9IEyfuIRayL137hwutJ7gFuX4azO6vOkoe0mW3nMcCnPXvIyAU
allUtQxwHx1tpIRsf+iw673zAilt5SDrqAcgBhU2mffmA6FTxcsWAtwSyk/DWS8T
/wHYUCLQsWGVtsXe29oIf2RR8Re03dPy2h8mAfdpWi9a/Wlp0IEUJa+Nhf5ACZrl
w3zVyyYwfjN//rbyaj35xXhpaBIWK6QhaEYRc1Y/vw7jj4hh/KrIurcaytSP2ayj
UE68QdLOfysefhI2mTWKau4bD46yRWzYthSh4rG7EAw+S9O8MNYfrsJo5l6p8cGb
Fr7U29dpXWzzdwT6BWxOqsQCjpgd5fpbxd1tgWes7hsEQqejAeVlEG/raF5NCMAG
GRUDNAeE+rGLjHIzyiaE7y0KLR0f+NAG9kotFz1MESuYgGEcDFZ1H5TjZDJXtlSl
W9t6MJfRlQpvqCWggqmy+oCNHABzRuSsIysbc2r9HZtKqGvZADpCLQ2NFM2dnpmx
flQmnkRt5nHDvcpG5rbyRrbKa65h7hLg4+flUfYCjoUNyfCCAfNGj9RrapzU5U5v
W7Wjeod00iV0zFeLLo7Mxj0AY/9CHQiCLuovcZsKR2LrgdZ/CkCiLgMr1X7ShANm
0Xphtyah4gpdD8VcQ4SsQYcTXf0lu/g+Z418sCdSrw9hWgnhC6Yvpzxnn6KqMQZF
lZGHmyeU7NgXaCu4NkwC45xpi7z8x6Ub64K0aOkjPQLWA0nY+XgrN+q2cWtPY0g4
YG3AxOxZE83G4eK1572CHMYcsTkau+UuPX/Y1XbrFnu/FbQ1Y7XDl9RScIbIzVP5
eVJ3ngaCTtoSSGwfy4NRXnBM77uvwdSVK5S+b7Rs+ywvYy6ki9wT4L+4Nu89e1lK
CCadJ2ANx0LHe+kHTaxd32EHFiZv+OYD2EZb0q8M/kLFz+uwAODRXE+Iti0U8312
xj4rOmbHLpUMEXEZcstuJRqSL4oZt3bUmB+fdQI/ajtx5eIdk+ZHvV6Did0B2Yn+
ndCDSTgX0/YDFq5JJUGc+rqa3pP+677GaqAMzob4nk1jg4H8MFOY9c4yBo91krPt
NkHaP+dj//gZa9X3/YDBXf5LliUY7zC7xKK5fgACtV74ReJ5qvKQV1C8aFyxO6cK
PAUT029P1UcONgV28ZIp+zFKv4Tib+0Z0N9pO/TZiGtN0Y2CwrYYZunfEERUIFrC
yGEkWWkgaty2WQPIZrvQ7lxwwoAkTIvZKvTwi3Q+Paml+P81kcyztr0nXMmfQQVq
b3pyYmCgDWi0ihLwgINizfo2mhleC4NeYsgvaSy5taVVTKxg6doeWtUZqYtbvF3b
3fKMye6bk4F7g7YvPVCJDqJt6JKNXMEnxB4KHPQqrRrI5uzZqKCz2zSQgupKa1bo
VwF/Bg43krnpXFg2In6tQkm50wCJW1XEBtxbHclXUxdWE9Q8dMA9Yce1A6wgZ/VV
zZ/tYaSJX8FoaWtul50elPY+Hf0Z6N7jsDXkR0AxqeAGKTyEGm2+Tt4QI1GqmHSm
tUJa5Cfk6mDIJP1gqWU+uso4qIRDK3pr/8N95dFUG158wkcURo3XRxfyxWeZ8kQU
jB3KVIu4Zm88siF36BoNUQ0+msyCmiIRtGYx6m6j+PXBiR1/JwoHuq46rYcUUDS1
iGVLr5an5RjqTQMPtogWl7rjahzNxLNDaXgqRBWqYXGb3bT1l1LPDyJKWNne31+I
GbQSRkKJYrT2rfFvZTVUCh9ucKalWsSJkMFtbQMqzK/Vl0pJJvFoX0BT6gD1eMPy
ljzO4Snw2QZxVFczrl8VB22xf8KnHcfko4xoJjhS+nZD5ITUL8xh/qqKk5zhj9R5
gJvArWJIwWRW7CYxj0236mGyarSnrFwDH9zlgMQbpMM0hZb3DLHgR0Np01N2aPnT
4WkAu370QPuZHWeVFXJEdpOuaU+ExbhtoKnY5psLv0ySNKmMZziVtUX0DpbkbKxw
rg9LKrNxfvWrsEJBPlH5drcTt8viekz0s/mPn/Vmmuz/iJZoSrW2ydb7WnRvAgNh
GBZ/oN3UtpxrtqOOQI1eJXhv28DbuLupwyCo3rQYgtJpwYE7BZMQMoQYbyDEgzXo
XCDbTBmsvkUnLYM6ynqCLXSd0QwDE+N0xySfAETbnCMk5zpyIbKcOJQTPkCFPg3k
sBH7gykPxdbamlhR4yNgczovFSrnVxaFevOC1qzWVLkUQaV30TXV+ZSnl+nRX9eS
jlSqHhOgMU8kP6KWFLQLP60LeLnva66uoyS3F6oNb2MxKTSuVxVkWAc5TKh8pJzl
3CMR/bYyirF/C7XBQmVzZyGuNo+uR3mFBr5kjKHrtt+fh3lQEkYKDIpZzX/fVgs4
P76gF3Ljk5qWGM5KVxBGjRE426yEKGkZQ8PeKIh9z0xOm4sm5PB9ks6oYsHWkskN
m3l+ZrefWyy5owhSgme9KgUQtIq28chJVTTTzJn2tfaY/YGazsDR4ziHkZfhCSgo
SEKO8KB8shGgPMY4gs9PtF6jhe6FRGgAE55vD64IHeXoEeni69zC+IaeFDFwngDS
usFpsgkO25otnK4/TA4Z7L12trghcu+bH6jXuN3Jzda4D5fxrlcl/xmI2e9oCBKT
U504hsgK4AKa7qtUebvf64Bg8/ZfS2MVliclRe2kEZMqEKbZXJY4RWibEZSpsldy
NGn/FeHHElx97aT1l5wvDewLx7r7Y0A7DLRUaaA2jnKDjJSpciv5iGlJ/0dSoMoi
NBfmL5vbp49t4DX8UTqOh90dcpB1WcFPEJWLxeDnbhYJGaCS81UY9okJX/krtWR6
ohjIKk8qW/4N0Gt0UYSyImY8cZWHHiZzI0SA66QpPBLsst8GUhD356QdnInHJIqo
VayNz8xHCcSa5fhPhpV19b1hEhGwNB46zJHZrhgcCaHPIMptcITlLXYL2oH+BFpx
12+6NsyFKqx+wWRaLitamkDhb4HXX8uKjba2jXjc3RWIRcNIBqNXOM0RaFo9H4XS
LVtDB3U7g+ryTNS6YTzj+f3O2SuCN8+447OZvdiur2nMdy5gXVErczwnlOEtueyI
m7eiGNXxs9LxYlZLCXj6wWBdMQJ6Z5A6hxXttfLb8MpvuQvWlmmXYWwj24OkgmH1
MRpNehNvpiDYtiJwLnkuAaSqbn44wynn/J89r5TwOcCXUziVVG3v0arDjosyD/QI
raF0Ta8E0zem4ysaxsptQbDzEg625y40fO8T7tVa91W2eFi7zcGF3zF6Ry6IEcrl
LuV8Eg2sGgrDqk6IaVzcwVihrKXyl0CYuQYch85xdn3uaGRPOVDw1XeXtPhH8p7M
tf6J9o7BtITWwSgzesWMSfq+dULorf6LtHFDZWaTrSBWJ5i9ynQS+NB1naHnY9qe
XI1kqSymv0Vf0xsbc3UfP+18COTKXiuIZiCup6cCgR145Bhx9tfMWEcL8/AqaBgd
mOmyrEO4nnY3+lD9wF0hUQ3sq9RKKsxFzjfsltwtc7FD77zD7S/3RGyrExD9leu7
BAjd1LlMkeGCeOrd/TrvnqyOfAVNjBYhQxcgo4HKd2yp7rcqaxZ7TVx9EzQ+5e9/
+QvG1rNPdGp7NyxCZuHx3gBx2eYNiBa0aMwL348DhBG+7IrIULk7PiVYIk2Xf773
F462ujJG65jhBHnf43E4fH9jfWeJZP6FlVUaCUGSf0CZ3uclbxbLSYT4rMzaN/dK
0WPZWpCpyqw2v3cm+otRDWeEvq6PT1XusIkhEc0ClRI/kCgitFOqS/eQg7Datsa0
4FklN6M71/Knwf2omkGgBTfP4VQj6lgkWq2eVEiyCyBv6zAPPiXCEdR2bnFsqCBW
bwVavXrA0NPFpfHtK5p++2AvAgrE0KFHeBv2gO5ISQY0FbDuXPuj1PqycuF/DSUM
LFo58rwn3r8Aub/UHuyOOMBZI2fJPkShTPDTdnZxQK+W0XSFTdbAwvGxc29x90wC
oWwMw6JYrzDQExlYLBeySHiWs3285bc5A94yFyfbadsYOZ0Y/FSCFw5JC1+d2Im6
P0qxB6Az+6w1kPx7IZgtywK2alFjLoHi8Bz3N5KVMIqE6/Pst9HPQUJKH/UO3JPk
2C+ljmXNSPdk19YxlTmH9nSSu3JItlOuzdZ9C9f/J3WpB4ijD8YOf11HcrOtUsAq
x0TGAtt/T2+SQWx/ge3EXnobi25QjlxWAyPM+Y4mdNc4BMO5xe296DTwwmLyilA8
L7K8QcNiLjiAZ4TSNHgiNw+vtreNJVqk2AcDrCrEOB5AuiTdmvzoPmrCPiU3vJex
P236LwvqF4o+oEyqqGd2WvV6YyLsFtaTLiy/ibkn1Z9IjgFeVUZUMW5lhU/tEBDC
KR1KJHgqP3r0bL1s30giMl/ThhM5ebJFx8zK1KrUPTxCS0MIolEEGK4K1zDJxZCi
+yC3UoyiDB3qgLwy3rpDDMetGk1tJ0ywIbw1gysB0rbhIApO6JFlaE9Jb5Y6bPa2
LYUOqcSofl5liUSOA/m9g3bqtbKO1xEBnmhrGzqfcGrtMW/qR8a+AiyIRxcoDNZu
qSfdWc2qxKHAmwQYD2z9WMDFPCcirET+Hn9FJPXdsfkgq9FK1MAnq3sE5R7KDVV/
Kk88KsvSo/+e0sGQohFDab+sHgLckW3Y4qkFRp/33mRGLiq8EwGLch8d/8TRV8US
OprvktSMMhQ9sXywnZFwZ6fEygcEv41C0FA6V2lp34GCmrVh8b+T9h7X8t18zy9h
noBqE0f0IbDIKGFCtLhYdrcK0uE4XCXFS0dTFDLgAlJ7tRxrekVlsWsOYqajMdam
YtcTvLhF8KtZ/765yJ6E0v/KYQ6ykwWZD3kFVxwwrqBPTw4n6x1k6NYRC9yCA7Ta
7fFcz5iNla3MSS9/pMzt8gMS63egOT8zZm+vfwU7Os0+kMtuUtUsDMRYBRqZVplJ
4+kCTZaAme699jkqMz4J1RNGEVWg1TXumhyiqXuwS3jc/fX3UF0S5DUJsR4oZI76
SIgyKuiSUZOhEUfMoaVIgVuq1qpFMre21t+8qubUO/cT2kNtOzzlMnNeWdUDGV0c
1yjRrYGkG9o8UsjTJBjKlfaADMR6FghR5ktE8ip8W+2qUqxZdAhYfWNqDyq+VtwN
OX1TNYQYub6nGI/FrV+VPIj8FKowGMl1qMJAbrcItS9u+F6PXGAK80Kt39a2io7X
bVahloQseG/HOfCV1gZSeojGFuuUGRaZh/adX6crC5FzmVZf2kpjjh9biIr9r3Ey
5Drq69FpX/mgxJ3QLX92FjY8wDFWsa16HOOho6LpFYFIWbJ8m45D7UaaNxdl+pWx
xpJKgq+V2Plqq+YDf0rRGJc82Hd2xmaiARQSLLMq5qDp9udfsLqoUMHJTVLyJKx7
M/5UwCVZHO24IvIKL6xQSHGaj9QGlOVOixu/8y6eeCNqi50pIWq6WlxcQ1gyAnS2
XBCNjVTfUZYcq527204cLgvVP4w1/OmFwt1s3eJ3Ivu6xbp9P/IIZjbmK0OVOgag
FlUcHfv1kwK7TV1WjsAMBZ866BFKKJs9lCReAdeaYCz6y9tC2lv1V2RacnzvmyYH
gallBszKKCrD1MdYtrAByeQ/aaKEeJbgFEKMqwKAZSuhREuY26Svc6y9OBF2uf/R
1SfKO/22RooexP+3oQhASzWzlmASGncJyYbYDsJPs7ui1CObJnQ/TnKEdr+4xqOb
vrzRawIweTBfIJWFNPjq6EQ0SkeJgLVx2hVtojZ19SKqpJA2ivnHDPC4TiTZO+Xq
FFLidJ76rtd6v6vq5AYKAdPCJwYWFLl7LRHtoEL+4PfOIx6tbDROy1nJdKUQEBg4
Y/K3TVdyQ1Jn7roZLAuQv+aGTYRh5R3VzBZN+l7Cq4djkfys3LcuYu5Q5B0f3MFe
r86mjt6/zpEaFAudaPehUo56o3Dou3WqEte97C7KE0GSOR0uTzLD8b/1BIAOBDMH
c3R3IgTjNYIplfH3LhExX8pUi+ck5/ZbYhGvjlQdAMjepwoB74dH6E+HqAMvsCJr
Ox7TnPdjP9THDEmqPGS+q7dWLSHGRJJsWq/Z4tiuHexKKwMpSq/GCKCCgFy/mcK0
jsN9FeJKOBgMSSNGgJEExzP4Pe/kJwOSYG8aiAIRu2hYz8Ok2Wvu9ZeiJdQto61K
R+fvTj56HOkn18Iviyd5benqLceuru09B2aGN3Rklx1gliCRfr49L6QU/0cnZb5s
tRQDDCGd69ioSx0rMm6CYJfqb4VVOViyZRPUIgC4C/eKkPqqtjKCMkOFeiGQAL87
DitgCDElB8CR7qEOk33usqcdmiD/RBoq6gUjZiVYVWKV2/wr2g0N6AjexV4qHaB5
ChXrVLAPxhzISDJtYMXGIEizdzHcepuB14f1+eebXi7iJZHkPQ4aa9tyc3wE+hu8
3qnyACUEeCB0EmWkj9cDmnrqGseECpUsKZEfBBUry5odT2BN2L5y+Hiw1UpOybVC
ftzJ7uWogmadXEaHzkUNUH40gI6QAjN4XmDB67qHO+rGp3APhWaENMy6skBATyY/
TwXLsQDqTTowOOZhpPiE+KsXqZACfIFhrY8HaI0E4chb/mWcjXrhfpnvYnyl/xEL
nGZ2blX/uhmM6HLa2m8d4Qcm569a7TWqZxORIK5KLZOi39jqYbJdYfInS74QD9X+
jHrnM2gso6eHjLTbXSYTae/lcITrJOYZgMdFBVSZftSPMomeUZaJHRWxYzeacpBz
IScxWFX2lQFy4JqmpGopxhdr1hEcY5VcPJ962W4Zal5Cez0Zyurmi7s2mozllBNK
S5O84n7ww5UULcvGVISQ6sSZ1LtLrY5GHAc8HclJqUeKMt+mQ2P8wS+obJSdgSma
DIUmFCHuO7oouaOQH9VWVRNhFDH+MI1wKxtJ7wGYLhLmr4iqXGePQefEOctUXmwa
EI5F/4sUXALN/u10GhrbmX8/5mJiBrjtUqH2rqpl9SNhNzXFEmPZxHo6yHB14Wzd
9zGJ/dXcKNQlkKmG7gCuGV+3dIlugZEmPCeoyUth60Qxk0eUwsojPJopAzCUvt04
9UPEWSQUfhMeVftdvIEaHkWi/tUGscDRrExbR2cSiQEsg/ZrqIbWEXJ+quNVD6nz
eK6gLraz9SHxXr1YY3aRXSy2lT11vr2a800tFcPjeqURNMzz3C5di93Uxcyzw+PX
e0GxjgnCZZLLKjQrSR8KV8gXKN3XGyS0m2qeuBXIyC3ajT8e1hlxhxzH5K9utPHT
EKG8JyQbv+HAW2vg6iOFuNiCs90fvNDkgRTU+ioc75YCakoJ4G6x6/yp7b1fPxY9
XiyssUsmRBo6ghYucHf6rC2YJ/pMRCYMYinPstBqwx3ESl68LRbJJB5H7/WpTTfy
YYpeuELDFGeHAwoEbrjp798VyLWG1chnOyBCOebu7v47XGq/cuoj3gtFG4yCrbfO
Xw0Q1oOMOIX0wWmsF/1JYU5zz0agcXHOgR0Zli0aTE4WD7J2dGQCU6ZgVDnYFyMI
WHgp3ahY0pHTBx0Y1bdYtyqEyLH9w42fh/tcy50ubJYYVH4Il1RDknZNUedXYTla
L9zZKDjSXtbxyNDPUaUrtLFMjVa+1Kzb9lnXtE5d7Cxsz5inoj+AfWkepAqDcxkr
VQibVRSKd+lcVwWm7bSQNyC0LGJHv0fYj0fFGZiFMnX0Zi6ijDrZ7xNykZwyftbV
TK9iVRQ+fON0pHkBOAnSxDBQG6Z0amc6KM+xmPzAv3Eiq6wFV+cjBVdAh+a2cjYW
/RVJRDq098jS8tzWTqlWlQBJd+SYO3A7/DrCxdVQTA8BLuftEoJDQH3RfSCmNUDj
XZRFjXsxNcCRKZqMU2Wi33qMnoF+KJ1u2zQHu6TOtuKSFITeu2uAL7jdLb4+Lxqf
t7ajBgQgWT+22vxPabxp1EUsv0cz0GDa9xO8NfVDXC9Z4XZpE+2UNJY4QxxX9nwo
VUIKWDhuIfGr3otc9Lz8nrSNTlYZdWT4KsYbEvZs3XiZq44/yJYMPUOH8Kdxq6kH
bNETeU7SXF3VF/OXv/Ws1/BEMCJ2hrRbuL4ZixTP+5ENNiVK5Ihftfk7tgDhgi9X
J6qM+kFfR3v9Y0LK4mbuDvViandHaazPoKQZpva8Q5kegjStDwl5TTJ2t5FSW59M
g06D+mGwfI77l3zvzb8U31nMfp9z0VfDu49SBfdX7qc9c23+D6eKaIgHEI1kdgBD
LrIsXroAH3UR+/0UrRhMkr0nNQzZm9RGtn7Jbi+nhoUEjktLsNgQj4JvocsLCDLy
3zGidMcsTm+CssY9JHQKB8JHHtbLORqyWrv5d32Kxy7FLODrREjb3A+V4NRgQMUR
ddjsYG1912khMIVYnXwQgysdzZneg8bfriQU9R0hJPOU3CAPFfrz81xmIQQIMwoi
buMSYsiO/yBe+5rj+jHitcso/rqWThDttPbVsAGLIzCI6M9e8A42lnQ3WRwclTbD
Ycb2uadvaxpTJPwM7ogxvARgmUh6Ak2qoJjRvWTZ9rj7YujK07s7dns0Rh0hWMeh
w6USH5KA31oKvhWqgOOG8ymj3CiJtsmPIk3cpSpRABofD7iNjLfLWhOYQeGFt9J5
eL+3ljB+zKUUrsCpFbyoqACEigmqjTi0lTZY0S2Vpm3N/GgUygEgY+3FdM7Ru6LF
tMv1olXwyYvO4f0znDxWdWPvNMYwoJDVe0Wzon/pSnh/HwxHgggLAQip7Yz2TykT
gxOhW1MdUjRlBDhEuHi5zMWO8f8yEMbNLSqjCShEPt0oLlKCU85sdbrQjxlPW1r7
ATG04rYbvgvBhzrCYl2hWR6mvT0c4dWay7jl8M0LNVMystakKz+5/8F8wO0XngOc
6G+/JBj/VVMVYOsPWQbwz0PE9NPKCDA15TLeErxpXYJpJ5nSlYwvXsfGB7FYL4sc
jWaJ5gN2OoK3KjDRQN4IKWXKZEknh1xR6PPJMRtlXBjqceyEHo1WdZteIWLR6djE
QVKnsfQQ6auHRkWZb+EQgOYbTdKI17iH+QGx0O30cXHrtBj+wfRFUXUTOqkeCKWn
SQZ68AS9jN9kPcA6GmF+2bSk/G0vueER8jL5vtoSLsxjCNhKPpPEEJ6ZAzAW5x6V
BZhX887u/TsJretA23FUqXPAbM0/ipJzOa4NH2b02aWXLsQySECq5AdLRLvXGrLh
gX9Ri/ohVa9FeY/tdut/8IGuoUXWJvMFcEG9cBui5VKVBupW1qcw0WLFsyBiH/HW
cONM2aoB0nBI23YP3+mnlDB4CpDsTip+I/nAS1Abx6z+kftWBO+jgg428FILq201
33UKLfu19JLStRPQAsbILuqxHgtJXx5DG/P4VstY31GSlq/hNlBw5ozdtLSONm8O
H2WCRhzcCDtzBuyPDB5zyXsJpHT++rVqQoe6v/QjyaYYJ5o90ICP2c+w4peAMO3c
ThTm+ZN/0RIOms+b3kC0SMbl1es4hEJ2nhZymID3MBAPhBHvzrlAYOZYaUarXcV9
bPTEP0eQPsSvUm2/cQfkYH5PgjOvKT9Su0zCha6xDFDhORjfT+Qnhuo6+fc9gb2/
FWH01qrjbHko46wx4TUPtciZYcmNCHLhOWHYfJ/jgS6lHRE0erAdGs/7hYr8Xlo0
s0aLm5LTeNt13JkNcnjxDAg52sxcCHTNh/eOLFoo/vY2RJ6mQ5CqIjTRkTY2FMsS
fpXrxRCwEdLfByGvXQ9CPxh0dXUnTsN+GFhD3Q5c1bJiUHJE1G4wGiu3X/W+uhgQ
/G2Jvqef9S4RJK2Lpgai0TdRI6QF5VhhIok/V9apUiJccFzistJfImjnnwMBjj6R
iZz6KM1/70BM6xk2hhWdLr+SBCnnWYEDoNMswDtRWf6F+0yCzyOGz9vHC6gGWKmV
pqXJtofxMkIecJC6G7v7E3OuGR/JFjDql5oyrKo0x5MPEezyV+88kDmhjBrg7j+5
qoUmG2FaBuP2sT59wPke/9PvNV++h+LMNlFSyyHucOzuzCS/9c7A6NMjqx7D2SkJ
9g1z+D/+4OC1l/iz1IcTGNq0n2xzCqFpZ6dVKPNVqFH2hvRLP1Xd3aUhdqcCJr8h
4fvaGb76VLLfXsOcqR4hUkbUeI7mfz2/6VSewIwiR4yIg9iKAcWD4RQNl8qZtPHa
JTSPrJ+IqTHxsqlq1V/suv8jQrU5K2RxpDgEcB2Y7bfAfZSq6JlLJGqitGcjmRTO
l6KtY38h+hkn/IsxltLsq3c5vJ3GDu9mXnYupy5/p/1kn4XzaV32QyrL4w/yzMGu
6k7Fq74jkRUPfzX/2z5quiuhJXD1uAFBbxCNCrGXbaVmpTFzVUUDQpGzppKfG+mH
wZsSvJk/VAQ2tpJRhug55ozt4aV6XzZ9+f6zWeDiDe7jG4QQnFEjQOPlVbnU2I4w
dzGgbvRx1x/CGVLhQcIwy4NBi5a0M3ScElAou2LuTm7eNy2ueMOdmXEEmYr1wZO8
mWXsQSmm2ycvf+WEsU/5bj5yijd+tWh/Cidx6+dVweBiRkUTE7UUU2hZI2qL1zDq
7K5Ofhnb9vv2ExUQ6fGxwt0d9HvDbpQuTiuntG+xYz/KvOTmpHfaiWlE68Lf1h3n
wsvza8auanCQK0CqiiL+fSH3kGCB8UbuaJLHnWpe1aPGJ0xGUfMyZEQbEX7DFs/x
PTFBC4NNDbjwljZ9Ix2ivXVLWDgqX3UuQG3Nvl8vy/XZayPP7XR61dsbZUyaDvT+
bV8GXifCzUQijghIl8TrDB90luWub4aiaUiFAeNEmdayo+BeKMN+BfO9qE85jiqr
umO8t6Q/v4dVtoLdcGTg8New8ndxpTLfunvELE5jpXj5AUly7N43l3IsSiV9rVbp
5v4TUJEy/daR1N2lTz9KQQFYQuQa+Z9FqlbkljXp5J0aF21KggBkE72dAYg+gfEp
mwt7bzSaIQ9M3Vrh5HnX+tKVeBx4FHGjeUQaQMYNyW43pM7DQKbd2zuxHHm6EhEf
ZCG6CzjPoEcPSfSUX1pEL8S8FgCBi68ig6vz1zz3Nlfopyv0dmLfoYE3+5OsSIEu
BQt526Wym77Z21Iu4oxF8p6mQz+cLVFfA0TTMEn6XMOxPDVT8OqNcYMozFFWG91D
rASLGxxUKySxzEQ7ln8OGOXITsS47BB/6gwqbR2uZ4CtBPpsmZFr+h/CYpXXZXOB
KP13+Ja4qA3SraBTNt+ukAMqlDJrOteNmEiTrkOEpuhhHQ5Zexul+/ozx+ZO7Cr7
g6oxHOxlDMtwkPQt3uLPuU/Gepd/zNcw+Y5WxEeY05mQbiiS8tpP83Hmc0qZuvaq
V2Ge6/aRyqhF4/JofJI0QSYGFlpW5NtrsIYrWdK+IrjbUBgBEdNcpPKNH+bvZTCV
x1g0B/8V1p/79V+36EAS37050t53QnM2E2VeltEH7gpTXoTq6feCGx0RI9MHkd7P
dbQspFpmmNIwghO8cN/BAJqb/QSVGTPRClRKkC2ifqoYOPYPyrWrobVSVrb4XQLt
FCTEEV6Jf69HledbYhkbj6qz2HipeqKkICcgA9OAoZu4UYDzlPvhHT1dFfBLX1f7
dGxtHBGH1Bkslk2NWQIlRSzLpqS78s2uOyLby9S9/u0oGziQ5hCDt9l/WcIPWMND
NTZ16Ek9DvkeLoyI/FRz2zEgRV4VuHaKDJ6grmXgLZcbbeef8qjOWB2ZutqXOnTQ
bAkKVL5EQhwHVQ5AoIJJS6VS5Hbv0OY1fqRxgFFDOuv2nhn+lahDbS+gMR/6FhMk
0AGIPmMSPOv0LMt0Jox1bXUDnBN0k6gB5f6EVGVmcIsTG4ZVedLAmkQMk1lRlonZ
fkfOwvdkX5TCPzn3bNCnBGS02psZgUtfFKY0Jc2Kp43Xus0y0FY6r+Anh0a2sjzB
IXebc9Z9jt8q9VlmzyxEKNZ3mF5pqlTiwZqDlcsw9UmvVZSqZndB2XhEE6el0PAE
bcH3qtWol/c0ZOKVnepN35cw686ST2Xmn6fssqE6+xAeMgyzX85ntp5O3t+R0NPF
tz0CuDnBrJsDBkNBuOZInIvCUyjKXMDP011Eb8czKGzvOSLEqDeQoKBMWZ0Tm385
Oug2Nzmb7k5XlgX5nNTDWMhZZ2RGky1uuSOQOjxe73+2CtY2w/9Y+nubvKfFgc19
3rd1jCYcBsN69EWsxEPhsiJIaTl5UxfJ4pC9FOfnxFas2OWlLwwZ8hZBXvWuCgE9
6/Ih/cLwN/Mn7bLxn7iFNNmFfBaCXj5UrLIWsWn8H03lTKOi32Yekkgw/EV+H2WV
U6YvtsBLjtGrnUWNhTEQ4YWb9dLTAipR94czkl1w2O2aQJywdfYmu6h/4wbfYaVx
RqRJEVQnfqFqgKyj8UnUX2i+TE0VwtDpF3fxE6VKnEjKF3iX/RZcdHpYxsAsAKxO
ebKUEWclfsJMDz1mOgmPt6G3L2JYxDfLN+KTVr0RGT99IOuRQ1zCE/4zDgdHNc1R
t+2jrku4kukjWoba95k+ov1gO6+ZM3W0BB8xz6KolxbohX0HQwWDKP7KmGNPLUNJ
vrEzNvZM+KPfweA88RYRV4bnYdaLaSAj3H9s58q2sLXDv2eTYWPnJ0Wl2d73cgwZ
jxB3RD0ZmmaOWx6gbsS6St+OMhoSsw3VAtFo2sbymA2n3d4EF8YqcynozSF40Hym
LimbL6vMrpDYvVeiG+4ixJ5gPmla1bfciqfTk2+yGWYRiKZYpMw6Y9S87pCB8Irs
Ifc0+pjhLj9Namn8Q4TMAYk3GaQi9cX0cabmN0AY/JGCmtLGzVYMixxUYmURHax5
fdzz5s0tElsUJlw+DoUWa3CYqKWR1SlzEjd1ZgCgDiRIYEk7UTiYoH997ZfbiD+3
EB8tLJFE13yjn11Pa9oUixzY/6+6pkstQ8WJFi4ZDkkhxg9hkETqBNiInIcCeHdc
pd3Sv4FbPMKIjMyUT7s2+Tf/l+3Ed9ger78W2ExLwhxpNmMa60UiOYOCcT7awybZ
aJUnoC+QRDkGO2qtaoyAVUMjPabuov6o8u7SyvvENh49RkPV+MEdLupIXEp4momF
ZCQRdG4s45NInF9l99neofOLGPAsP1jEq2X1RhM8ovCP4QufFLZ9Egn55FgQNh6u
gzEx3KoT77xOTzC0p1GNa+Z5tznXWXr82mCaex5mdgWrJEOq7o4dV5v+DFannqyY
Es8OHgTg3G2VNIzsP2p6UVrDWUnYcaClGVzC9EnJX1ZUO08d8i5F9sF2IQGHzMv/
XLKlooy2e8LMJv0/uZUdIJ8iOF27sJLCfe0YnZZAXwsYNj5YWr2wCIOageN32KYO
P0pUDNYZnVj63noiraZ3izJuZDuDr6TQA+SSUCWiPt/2p7Ez2IT248nVmM6X3RZj
VkFdkkxpKaz162Swzk/li/5zJJQ3dsJ0bF+O0E850s5prcH66FTpHQTuUMRTK+vu
ZKxXM0DcSGG+tH5o+d5nGiHOIOBsPe3mf+G7yLZ3u6s7nmH9zkoAHieWz2l9SHgC
ZKjScCig0/jCug06xvtonqZzzqFaw70R9/TEHLAfuNIDmMP93bDHiHCMKaxZg6mi
dop26DdXQDJPE5ZBXVmaJmVUjb2Ahp84qz+fahzmAk9hzkcQIzlaeFjMZASWdkxH
YvokgWMK4Aa6k495oaBZaFi6hgbxfbjUCfkMltI9oyK3+wmz0qCzCwd89Y9g158B
V38hg00upyVl+Hif05K3opQh4OuVDrdD9vkmpilQAJoTXJBGTGeret+/zHCEK6fb
sVB54ys7hSibhogpr8cQ9cgdcoHKe8bz2e/o1DIkzN/jVKRHpmGTjbL5N2JeaQ1o
odFakYnPIEKuJgvdtWmn9UdhUtq/Njo1yAcdhfJFo9fN+N0lxB9o1WE8kpDVY8CC
2ssClYu+s7mABM3+nvFz2dVHmcfsjiIX2vQa/CnCYJ+fa6ishkJ/oGOv+yHJxxpx
6RDBhiusy82MpyMsJlo3Eb3vfmoMro5aVtv7oikNQhL+jLiflI+Ygkz/o7zccNp0
Eu0PfWuKlPBC9vk1A1wc2IGZ2WPXbyiyfHkU24X/5knavCbObJZ6nCu4olD4sfKM
8BTzcbnHkGLgyxifRoQItSUMU8ThdZd7K1y8XTB8JTi4NNbuYtp6QFTfPbmSSUar
AlkI5+cgcA8dBchuW6oxg5S77YBclKkjSNVKzz7PtTdBmUeIQbrudNCUIofdXjZt
Ql4TkLoOztDrBvH1G8RyqYAewT8/BE5ZBL1VLze1RYJ5iBj4eto6c3ZEH5u0lyfa
XQi7wGS6p+YsY6B8WCKlaWd4wkHLSLU6sqJKaOCelWcuEEkhPSIsFnmlusIfxAmr
Yn5lMplNA9AUnM+sNhBhU5eidWGO+OY6bE8mOYPayTpIoaNBwAeT3jbZu+3XavWe
JQhuyOxmZ001IjcLhyKZHyA3lJSzvm8zvMp8qVr1WKAX48YQBsUAbt+hrxviOULr
ft7DKzmDI1Yrq6PFdFApdjq+veEu94ZdVnzO1wdBJP2Ao5SuEJAhTVMU/s8jeRSI
AZdmc5jwKWoA9G2dTfP2vJ8IOOiP4FVDmj9+JIM6nT4CSU3LCgRH4oxP3VTnEulD
w/4cndFRlrBZOMP/MHwcUVGDt8Wd/zRJkIoTzO89bbL6k0vaQjToFKoc7yOZ1zw8
xQSsZ7MHyGqEzo42hwRZ896P7ccoqCGhqumc8vSW7IZL9h8ERexPj19lN7cZ1eDX
tjrQo4TitHtc9xMBnu32doRgdnWamHwyfxLKn8fH2smTp9TZ2OoeEIJSiBKBoDVt
xGWIF4GZOXm1Yuup8tGjy5e2tw0S6Zv3bDPrzbMbzS6bA4auw2+YmqXNeS/padVj
NdpJL43F2qzK8Wf9nQSIkqfTEuffdgKLUKdC1RWjoPwyjOEliSW8LtX2EDIjXW4l
NczNZp2PaLI327eiSgpeGs7xR3plkN+JIYxqF2vARE6hhK79fTW3bq2SwAv/kR2n
09Iu3IklF1ZAkP65qLU2NexImBgL18oQcWHtelkl8+XKb5GXElRhqUG61fOEqR8I
PnwmLoNQk55qGA3osivUd0rfUFNHLsgLrT1lnlS7zV3MlIjSyEStSttv2VgYWtew
vviRiT3zA3IyJfbIm7tTSJYoiTdY7BudNDPSes9YcFqWmT3/rwIkLJ6KfGIyqSF2
AgV8xCbISkLtAyxV5WSzwJueqAJevgCoCMSB6hiyAlGC+5QeevNsDF3kjKYWOXKJ
CMRrCMNy+SWiQ3NsWKhId2Kb1RCXrlyUIEk+ruBnzYdtXaNM+WQGPENfkWljKfor
B7PqpYEwaP/iYazm7uaYD3FD3MxhNN5XqX0JmkoHNNLYON0iXPIU78d4clfxJ3Zp
zNRSqW9EbTG0fao4H4YKWcAMihBtEfVbV9Fsu7UR4rIFmw/zNAUYBisHi03mZsHH
uqbnTihsdxuYEg9kvOf8bqhePTBZa/DSab/CzbhVsQlzBSswyL02BdFdc/XiB1td
iF3S3n0kxAEVyaDi61DA1Dw66twmzMaf6L17gAjru7YcXIOqrHvISVWp+nrr+jk3
p2Sqtd/kuWsVLUPTG8ED/OPwHG6SzysAE+4t4QTeoZKaKEJDml3UNtGrduHGZiNx
aPj1FomhSlaAxKO+zsYgzJ+uv7+Nvi5Iqz13bk9Goquu+0czR+S53mUJtUqzdvau
rbRrnMBHU3usGRJoj7THVgt3bLtiGQE2XeU6qffqkvm4R2z2GNbHmWUzOMWgK+uN
eRdHwoBv7WmU2gIc0JqEewZCk6OkQd5ym0BCbxD0tXMvPe86nmYt+RPoYFPnM2f7
ozEIdRFeELmB4FN51n4YJq+t6ewsR7FvAlnh7Ck7Ws5sUXowESQ7jvZx/6V7lLZz
hsoIAcjQvP9dZgObkMcLXKBNk4chH+aUqlfXu8oDLBJoR8VDtATWNK9xGYL42nGh
YOPJZbQvZdPZZyJCZ03ofDnVaEs7k77Heo8Iw0sW6SGfjmCxXycVkfvfMJZIeoH3
ShY56Adlxb1q8j9Ta1/zzxON5x9MQRM5Cp6Ze/fZ0iKdXJ5L8PI8/3ZrOEDP2LTK
84QEjYHLnxw428sMdgcg3+NI9PHqFJe8TJqnq/aNfnsbYt/EGD1h8emfYnUhz028
inL1aeJItQVTsV6YYUTz6JLy77s2E4KxB60WdESaAUjNWNOleltAow+NFdipPaqU
cKGqMNjJs1qfW/9sHc+XyamwPDE9ftKKlnNRO8oXMRrmPnXBgGC81yqcFhAwfZoM
Kd43d7FOKgTwFrLQDUtK+K4t+y1nPflLQ9e+IlwbUUVfC2KrrbspQUTfqSgQSSAJ
cSUviZsk93HxycvfdFI0lFRz6X0FCShwlMR/eTMqf6K76KWdR553hYxP0bARyrl0
H0hQhDAsfq/qTgKWKP/hJ2jN/KcK+wd2vaNOk32lCAPnDeMa2piOnX/5HzpMu/Ct
2pvT7zoXGvSieuHq96ajc0taZYnzKjQa1IFEPwaJ3lTq5BZKRsfHord4Kr0gZGrF
PciL7RfUi1rIVURN3zAK/aLPRdj7stnaJc+QDlFstFJGNOBpReO4kXOi44yLT8tt
xQDr3Wl19oE7nQjZwBn8130dPeUs1ww94mEdfeEE6k3jT/BEKRroCWIOjD1vtAsy
AM6QbNAomHebgHyjMoeeKfKLNSdtbQSjxikhEK3M02+Z4u7gKWP0PxiicUAcMEKi
lryJH3JSO0SJ5xpXzZTHRTG0dKjFpzAupIEW1tj90lCZ2+Nv1ley2LyoSSCxsWT2
Qs/5CuoreBg2evXdsKpkwtLragWrKorI/sSkbU2Mva3ldHVD06z+juAxeFtEthLI
bD5o7589UCoF94T3KjMGKlAaUM2gUdFGum+mA9qZl88QIqccTBCbrgb5kr9KAkYZ
SHrw9+Kr+iQHAGi4XZ66KcGaOK4R9h709/rdmKLDFXmEAzT3ZxjUMZSVMxW5rIxK
d9ee8GfmhKs/J2TYnS8B3PrZsEfg0tKiVzz0cz2s7sJh17WQ6sKt1V7HJRva/WUD
1FZ4A8ETSYwF1p0aV5ow6uDPBA7fyfWgdDrPKUvMUaivtL73D9/EbbRylJnM1ihw
W4mBLrSxk+e+UQidGz92Yz3hxsPLFb/2BprEsUb3WIBo8byFi/aUCAD1MUBYDtQu
9n/de4H9ZQZ/wFH2FT6Y9QhcGudxY9txm8i+UNL8hfovLKP2tzzjVDkQfXrghUyr
nfh33Cx78XDW3lcQNxO1K4NdP1JTNImnb3Es2cnVFoN/I1s4NdVEOHq2d1rynCUs
678ZivJO6Ezget8rF9Ekwdxk+kWQEkfsLgc4FKHFjWsFQrPrUoQ2dWZOEKpQ+YuF
QsbyA1wCzeXLU6+MRWc3UULlMNDrs8CV68oSvSMvUipb6wBKSofG6ee7rXgdI2I7
70tRnUuoTtUs3WiZRYJNTNiK/CTuxJfjcbsgrFs4CfXerLz7Uz6cIZd9Ui4IGfO2
rqprozios2CGmMSbfCpGIPF/GZ5hagSij5U3dq4YH/qvOobLN+u0VFKcOuo71a9W
TzTHISiNbcyds+K4Sqi1YW5usuWRtqtPvLeqy7K3ny5id85Z84h1uzzmPDU2XeaH
/jnAxByHtStbBlTTuJ9P4MW03EfIg/OwVIsSlk8OAL/Itm82Yqa0g55LeV1c9qjt
UKOGOG+DGk7koWDfTVoPHs5daL1un+rukK1HGxHE3PP8bEiVXFWA+8t6FKZBaf9o
IN60oTblj6ek5TiW8FZPLwnbY0rKRUO852EGESWerdDewwalR2np/8dq7z1RM+HR
YuCberkeMdQPllYY/BQ4LRADLZ8GQEr8C/2PwsaerOcrKW9mSCV7sychb1etMS42
caPsNltA0QnuAFil9Pv+o/ILYS0M7cT1HP3K0Ta/x/6RKMRS5dL8qpGX38XDds0j
g9pnW7CeQOxSytxETaicScYC17AUNWnXXa/Z5fWn1pFmJytihrCMVJaqwskbfYp4
bXAt64DhAKn80ZSPSXbKxnlSKLrPdaEOIULsRAWi/FKXmnuxmEELHn7bkpfYsakB
hVPLTKz3ch33Om4alQj8BQ/6aWK2vTV98gk9GjRq2S5Dyn4mCXVygvy6Rswwizn+
C2xLi7muDfHCDGYSfcrbprQbaeEAzynt3vQE7dymoOEsO8VjqyBgEIzgFR/zU7wA
0OltgH+5p+YipODEWtx9kr2BHJFSvIWPK2aREJvRrizkttaebSMQ5F+gQk8hMx0x
7U3MMj1p90mvwEvqecz7hvMnkzAw0PA33Wdh5WR7cPjxcOsYXFbzo0jaGQMxyvRY
crpS9tSs328EiP7lCvuIylpo7nMkpbpokCAkNgvZxDyBAVVjBaNXZztQThLXtjjo
EoAoKXNdMMM13iHWz+P7zn7Mb28OBf2/HEXnwsVnpAyAKknUjT+zw8EaPiaChe6E
UKcXdpkLrzD5Pyozg/oMqI/MLjUUPTQ9hEV/earejxPN2h4r3ROVRTPC6kqN7HuT
qPKC8oHi7envI9yb70PUW6PVe3viL6farwJzwVw35TfQVCtmYfO418LuLJ6eiTrs
zh+fzcD5NXNUA0fRfaDfvzXoPkXwEsgU+wTTkMSb30SihvPQNyi7RRHiE9wRkTbt
oAcafWFz0wQ6+XHw4Q400SaCBUddhygUBhmXhKPT4q6R4Ol0s0/OUNuZM/v+jj4r
7YNGrI0E3wudf5YPAgdN7wW4vIu2OqEgjaYUp/H7W49NGo8Zah3gc5/F53E4IlNt
wxQd3e9uMIs5QSCenZuquQ0PuUMLqqG6DTkRx46xmqjigT5PymEoUiHCmW5Ceigo
NkPGQ2lDpb18T5fIdGAPIMlSF40JgNov347ONWoC7igEvQtFnK35+C933ULPhj9j
ESr7TcPv/45gbn3kLwCEnrkF/Ba+gCSCyihZ7dIPDT/47Eruj1LgCifsRu6CP2xM
nnPH8VsEYafee+pDIp8VzKzFrzFZuJp7uWxYKgsX528xJ4HwYWR4y/5am7L6O192
AyiGzVQYYX+VAmDYMjYCGIv/mr5/zRL0HAUg/JE0bzsBTBQe0YNL/XtdEBPWFzRu
gCx5rh/sJv+4UCoES6MAzSCv02n18ouyyaPLljVCKnfJPN5aEdg9JtnLpTVjicbw
y0iA7wVYtzwmct/dgVDUd0LHZ/gA6WB8KIYcZ/mIODEgHqK8K0bXfoDguxfSeg3e
WEU54bswsQW0q7G6NtWL5DQGqYGx/XRb42/2S1YutPGz7wOA0a3Eb2IA9Jb2L0C5
HKiwPF+Ee0j60+CZiqsbTi3oK2oCKG54ZWdvUb3iwpQOiu+h4QZN3oIhmMsW/gIy
xNjXRT9I9kBL7Yx9YGJnkrNAbng1q6lxlKtBJt1gTczVaG0x3IA67jznasYHWHpE
npS9gx+fiL1qB07OguG2EHjplvGdu5T9oQUXFVt68coXoKXjW6PpZaN9I0YCqv6r
pDe6fNxmxlzuC/n0YF1VoSRIeOfgUHW/BE08Yup1KAVjWyXzQzBIERdkUCYmt/cT
Rww5JPjgTqyuY2hpVH6z1hVBlAmCnoYL732xQ26gtb+iOLrBI4FEfQQV8gV4IoRr
TyKrWIxEFgLSiUU1yQ9w6ZJgKpZXKDJhiGfeMmOE0GMkz/6vmLLsab2V0fR2TeDz
YBtJ61b/zcqR0bl/0Wp6Sv/7wStoJp7oJacVPp5zWFchu+d2GJgAqwluNbddYsnR
/oGieUtmlW5m0+K92hVzmWc2T8A5ykuWI/b/SidialeQ0AJNw82ApnyaKtm4dSDJ
a8G16zriqNerWXx4J872U398vK+8XJ7Hi+A2F2aZs7odAxRGGXBsTJYh9Q825lar
xheP0w1e0cDAWOpXyYBqM4JHt99UJ9JvK9uIKpJbqD2SaOjhCEkNT2IUEDT76nRv
kzHpGWKig2qfEeVC/4m0aO7bOoOC2UOBwL71iHCXA0KbiiTYib3I8+ei6tf4i/ur
Zsu3nnAlDqFywbBmnfat38hzmC6cU6iqNcstA3NMIwOjXRRbyoC0mLw4e+hXqZ1E
/uVvhGQfRGSmXDgC+2CevqKSAU97lNxWUuQNGoC0KyVjRLxc7lw9H1+/fQNy2lYG
8Y6N4inH8Tb+211ojWPlsSPA+yubi0+UcmKxms8o8gMjiMhQs3zteJFZO0fruRyO
iWCg9lyrGqz7C8YDDdNxiWUMq9SOdJBO2zvkIPZNd3JHqQJaoxitZ5ZKDwJ4JYFj
b38YEeoWzOFgCsbuWDNADfhiORYkHtBY6hg7lew5gpYap2S9ce26ziXDEAHJhWI5
CXZpNRvyUGSHBcAr/bpzsBQ0tgE8xCo1IRaC35YEEJ8K/Rxv6exH/0KYc0I/K17S
q/+35mIQy8/X05SpHIgv+yZXYFA0aWtKuTS+TwDVXZHb2bbOqK+6sbYynlR8CmLi
fknJU/e9DMyom6JCpqqa9Q54aQWrhv7mvYGuStnAIAE1qb7GqYUmuUVh5tVxsevK
KtcKD3nEfgRbJPW6xCVDdwwJDcenuiJbaNwJj9bSHk+p91xR53auMOC6fNNcf1Ds
IVge4NWjvhEzYgqJLnZP6IMZBPtiPfLamLEK2Xt5TmNVfmAVLONEZlOTYaNgMDEG
bYIB8aVDFctpo1ZPolfx66WcmAq1ch1S586C30DW/b0AQJPT7a5uEJO6GhHD00tX
fQtuHadpg5rEathkWU/TBo25AMTIgtcjVcRO/S/+c1NnY5Ti8q2360RmoThFji5S
K0AGQWGXnQBwFaSe0q8Uw+5NULgfdYX7tG3i/2ESbhmzrZg1kg72ncI2fGvUFZxW
G5uZ+0ZnFdJGQAoNBie55GmCamz0oPgqg9MSiS877z+q4NxaAG9zyx97RGZeuMfa
3ztZQl2+NBK4vK2q4+VeXKcO6fhER/UEZuoVBYniq7rr3UTeuiZiQCuF4GpNIue2
J8mbj68h41JIShkfwqhiGTDJSmS7zwc+kpdIYHoNLGS0otk5GNMyLlsOTaCCBQeq
q6Q+dEC3zYwOls7qKmR+05r4ohENXXV4uFx5GSNwL582HqUbGNUV3vbuRH4/lTo8
DsUXYDM5NXIG6LBOlh1n91Z2GkKpod0Kxfv1RI6bjwi3B2IReLGIc/Fs1uk6bCPZ
CSXTPNY3kZFxxUSTv0aQ7hBW/ehqylhYFp7Ai5SqdxSvT3f5PmQcxSXa3eRbCvuv
eY5T15UHMOvERlPpYvb4MMw0YW2nLcjztrVcamzL9eWlX6kt/Q0MpTD7xwfwIR87
b12uHMQLw7WEsXouigC+KzijTQaPsipeJ0oxdswNfiZHSKcvvEa9gRvM2AbI49WO
cbQclQAjQLrI8TFa2Zysvod069k232XlMVFlCXDI3W4yXIz9rT5BlCRofgYop8Qr
N3lCNb96dkWt1FoFtFCKPvla2a6JJwmXKMAQ2qO2y2zuIYOhxMsy4iIw0pbBbC/3
aGZZ0FhFX61ZPj2ea/cmaNMiob0Z5kuDPm15IxJgshr7y2YCfPRFacrmupnhrkg5
wFD6sBjzZZ91imyXPpLhOcnI71CpdnmBCKmMPl63x334kDauIlkJey/rpb7GvTfV
av25M1b4Cgl9Q91Cj6UON4N7LrUhPYd/1p/xEgWnnqK53UXRLh/z9wGmZ7BEn/sz
YEd2iQ5NmZejhrGlpWrlggkpcrIuVLjee89COYHrtYTrn5WwHbFw4OG1hqvaBaid
wWnQWgIBM9nv5EiQ35rHfdSfEnNHkHeXIOOfXpayvXEqLybV80qmQtNKr2DkDGnT
MHkdAQGj95FPeI66NV4aGP9F/P3GOTJP9xwfQokfgqwEighffKnp2MAc+PA0HAg/
nHi33KTYKgUS/A3qTZpMv9e2ddxfgrAib51WWyNi6v7vffZRwdgTzYoscPjOkgsy
s/J6odZQghO8i96bRv2mtNGIRommGo3ecmCcOL8JKDzTagY61UoCRDUeUNjNSbUI
8QGLx48+pnjqb62BuiciVU4v38JyqWvHCM59VM8mM06GyRzLNrRfNEgusFq9N1qH
QzZZqGUGHialdG5yMQ3ycGoZbpYbwS1Ab69ECsOOZ+nOVZ8FbZ4nLFFfEDIP6SCz
c0JWEoFhxkQ8xnoxNe8P68LMBwxz9nhrnQaVaDdZXZ96gMftHo23xyt9NzBc28Yq
zsPmvF/qdhtp10lj27lNlVnRCP0Jbd0LhlalzhXsPKASbe34UXhnD9vQEc/dPGGB
IF4cNaHewtAFqaHBZvPR+5gIXgRP4tGzWqxoR4D4bBnZqLooytk8QO3gRzfg2Xw6
frZDh6P5ttA49L/sZjY2pQqagFpKROlC4yUzHAVM2TT1PqU12zrfb3YSoaaUhVYv
VrtrzWIhtj7iVsrFGBIsQmdlawpPQSBTHTj42zBqW/BFTPo2raABahjGze+iZsx+
SK15Pkzhulb/Evn5OTdwpDJLQWWvh4JpAcUqZGA2fmAHSg9eA9LZj+fC+NEo8MQ7
/5uudoeTA8n+M+jVhJa6fpVcKrJ71GTEGj5NFUeTS1LLSivbfMYWlY5mguFnpAF2
6Orl9PTjNod73KM2FipdpiiLJx9oe6JrFDiq3D23AaEkjcFv+zVFw5q5QGmyPi+M
o/nZq8vWAADQPe6ZNQ//BX5mvN7s4wRjHNx8VQC47tdIcnyWZlOJaR1jUkTOn8vk
rTgiiL+Aitiq61jdookbLqRHAgPNJuJCbA2rKCZmYlPDyg6HvjKGqdfpTQUJTIdT
RHx/q4TeohxSRYHjvpRmWNo6xUhdoPczsO//ANV9yLNqpEHsU4LLxa1jGsRRsD9n
iKOimWyZsIL8LhJbuJXcJQy/bBkFY8j/xyQsR7Jma6F43WithhexQ3QdXtj9zNfS
biPwUh+jGA/91v0F1tkd3e/5DweFUr21rTnsGI0sgwj8MrucwXuC5YLawC5HWivA
JNxs7Ta5Y2e/HU4dkMJcQ89zwU+ec4X+kUJPWLtQmZRcZirYK85ZODroyaqigWca
KpOI2CfyH1Sodb7uhoAbOAuyV90XXoR25Lkrx13hfy49fANJQu+mctm+i5KUgocE
RJ1tAQbeLnKME9S0XEO1O9fi227hqKBwjDTEwwY79bCd8vpeumjWH66MKik8ORm0
JrOVpIoShOosUpmLcYcsy0AqH2TbEvXnsbPJ6vTsRrTQXWYnOzH/AokUczWQ9nDt
18ATmpmAB5P7LqL8DibTcYfi52acvewqofFr8R/s8pJQPaWr8pS2mNLbEUqNmhFT
kUCg0k/HBfMkQRD+FYDsg8GSFgSSvXhjp0ggV4ori+t6u+3n/CPPeHHWLLU/zVZX
aRacWnhlR/ZcaH/wtOZ2xK6hi8W2fSisSUAgO8c+kSQbjuIRin1oo+Hg9aI3FyzD
ZE9B12pUms60bKZ1FkPmOJ35p+UW0EpIhR18Fd2QWJx0dAQlfZ5yPnHvrUu9lZ87
/EHR0BtSE5RnsGNEoxnaDVVThbgscVIDpalAshtM5RTVRPGZBSjcngn+RXybHqWi
6zCOan9EBPgzPoQmFLh1I79sw4rO7VIwsNJ8Ks/xaCK0EqGI+UprR84vKhAGs80U
KuTnL80S0oBRZejXQQtb8W6gIaqRjeCKxDCI77uMuzj8APDbF8Be7bL9NOa1JZZa
Cu9lv45055IpHVHP53tEJYfTmK9KnFTan1YsbvVz8DH+TfGiidfehuGd8qePF+t6
4zoAeINOksJkLbeMeqE6K7Qaof4oM3EDCKy4pU8RoVHHWyrlkcOhDQ3GT96n5FJW
ziAVcyhi44m8cX1dEYirZXlJSSe0gh+4a9TwTZXTc93205KBgegbQbepch1lYQct
wrir8Tat6otTXCpOqRAsMA048Av6r2a8J/ReTsc/nJ4GRayT2qTsyzc3YquK6T8e
iJjGtZpw17ukOgjjZyOLo5axqGhOaLhgjeyMlX0NmZ2nvw7VWU/yL7IDy6bcti2V
dqqBeiKVcxh5mD7BRRbRtbDIDV3WTMW4QiW3AVrmg5/5xP9yCtFIb2Qisv/NTuHT
MZ7nHvhy/28FLUq15rFc+M02frAlCXd84EywnTWDy6W5E+AtOfuDUUwGXD2/lzdg
2noPE/kbFnSL/SeluYi5+NxP70HZlqxeur3wnkU5Z2jM/f9IDqYQ7zn46XPSXlgJ
ePXEsRVMNgMvg1UD8lmZpqdqotgmFuH8Fi5DxmZpOj6mbSpr4LQiLSkvWA+KIQW/
GFZ6Ifk9xqDFIoQV0XSjdb7/bF/YlRR/UGIhquQfOBGpD3KmfhwDzcqZo5Z3kKye
28rAmQGQ7S48ziAwRAKpThbhRH+HRm9BE5hueAEsHkZZGnGEGA7PLZlXsM/sD/Vy
4CVFLBel7dtUCDSW/jFodXFdiAZyobZtaJgmF05renQhhg0kmtF4GHMumj4mmnr9
LGKMdghVMRY9ETj+EG223DTbXENc+ChHcOxvNSwyzo0JM7N5fSrwqJEiox+p+3E8
IZWbd8YkS/Ft5wOF7YAJgqwCousxFuztNd4urSpyOvr+5b21TLxWInkKtWfAs98/
/+HZ5Xu/6siwetwDkh/3ld2VBQ2AoCgud2PD+bqYvu5JH0GOaCZBatrs2zuuPlw1
NyCBkp8sq1p/e9HwvvXakAya4aK8Zhuzjf+T+UE6CLSSbjrAMIg9fHIbYZLrPT+E
hQlJV51nhwOuGNQTXOG++4pgM1Q/ShkscAyywj5D0Uag5tSGPf3mRPqusVglQgm1
4J+OwxqgUC1yklJmPOhnH54h2PZDukkLc7JwVt3Hcq+XtFbm52JUhxB7HgTLM4Zp
f9z1zdpPB0GPh1SrN5xaS9/bxYy0u9NEi41EHpaHwXUMJF8Y9c+JNKFsb8yRmwti
B9Tlkk4Jp9wPe+CYw4E5swf1+9kjZEtNVcctrqC/+wDAtOM/SQSAHFHIW8VNFSYN
OMDrqHlshrY9D/jxbH7N+SH7Wpbx15hC5Izh+xxHkImDgvI8NnzXRJMqaH2qnroc
MNCL02CCUvZlRVDYKZew38LhP3y+8zB5y7DxMv5SlIGlnV9M2ibtuyPcj7P+OXXu
N2U4BwNlPaZkpK5kSHICZyOhpTK20XjpjfcZK7ayYc97TiasjQR98IE0ZD1GufHa
XkhjEN4KA3X8oA3nnkBAeiYCRlNW5gBfg2pzc/Peq9x/woM8MHmq6VIOnz5iDeKq
yBQ6Z/wEDfBpQ+KWsRw8fls3kXr0Yj45f4qfDk+Kazla7mKY8xakzfe0o3AoxWQO
XwtOEJUEWF6iVlKSIDyRHlZu74myswjjQLA9D8kIR0UXD/xdn/bC6DSBBBvOxNIn
lLgh3Ru+KRj2qyPJhXjOMAJwar9XJftfiW9igq4iS1FLhUVYQX+BEV73gpxeV6YV
JULNrg5vauQ8nmV/tcw6lCXBSHKaLdgGjWLkpNewNyzylPJYY0Z8gMJZXkuGCv8+
UOQNM/9KcjubvzMymL9dYTXyKmLK7mB5ofp5eEyFFqm/rHsLzCwp+6M4waO6uCzI
wXDRwm13E0Tx9EpExozhpCNef4qRP7BoN5gDLA9DvsL7M3tXCL9PU23NoLtRf3g7
PJFmWe2hjc0vcTTVLydjdKv6byYrdObXWsUpmfaTGhbdmJ07lDsKIwLfh1BcQ+TK
wQIOG75yrDjnnilwfPvpx96gKJ6VlcmtO0Rx39zwmcbshdZqcHO9nUIzbWKFwciR
sOT/sFvy1CmIhnv668XnNbR0A0LgTcPUTiFpPOPUHr+RrJcjvGKZOJcyv6iwtUCC
AsTSG6DWAjnX2LrqhtGB+M856dhD9ZrcloHNodHBNq6ea2HdIi8P/dPWlBkXvfJS
CTiJe7U85jABtCO1lrX1wMatA6U6DspblyqQnmA3Lkc/aP1fffCmQ72PBgOdh7ks
Us3Jy7N7qS+fxOGqrFyJi/LboE/Me6xSQr8TqwoHS9dka3RuSRkPKAGXd3IytP3N
1S6SvVgjXzqM4tK/6XIhDZSY9TgBI3pS78SI2xEwHZOCPkZKS76xkHXFq1rmzfac
yzPoLLBXCJE/Rl7HU5mWbyHhC+zoHC/0VV7084V3KGNe4pAcCfvPSSKhs4t9lXCU
NtzeQTJhz+CHHpYpHAqTpXro37u5gg0tSjmoxZQE9x9rWDYujUOYW2qQ+etbEagw
VgDOrO3MoJZ/kRjIujWhLd7QUtRXqXLjHiHWaPBXMXbhr/eQglAUbN6UEG7Zmiy0
ImNGvdN4uhA2bScn8MuhsF0WYdqBFngEr5f9Hi9frFGKePIW58yJ9+kDuo5TMvEd
lwESH3QGOZiaMDiBA1wCXYOW7Alh4YdHtjUoP83nZVB7YcTcoVqbjIGnrsW+kaiS
BNx5HIgj1IEgLyjxM3XSA0JG0d425HNlLe31cIKi0tx1UAg6FSWBeDHJtlm0T6hU
g69q/Zi+p/ocUw5dBMz613qlZVHJXM36xe37UOgXSz1D4PUhNYq+Q6/+7vjcE9XG
Yya3FccAy++XlHA5Py/RcBiVrOfku04Qgg1ILF1RAj4jnH1HENsCEFZ4Khim8CsR
Ax9UMJBnEF2qpc+a5bgLUrlO90kqqetoP6ZjGVeh8cDA3fIfc+mDMUImhR0y74/N
/wYW1YBJh8p4nYvxEQVXIbBY6hNKgo3m8QrCS5cEXeke9WA0cJgnQRuSKaOnIa1p
xREtARPxpA+r/9jvLhyW7TXiNtyecznZAz7je6/qzgsLNUcBUVhGPC6/9YExuEiH
SwqOR/MIdt7DfATPm6MKBmIE6pQpGz2a7CitLM1geP1s+172lACw/RmGtrvV6g9M
+SKbRGVvRAfa0W+5sc5K0/xtvxZq78WQcjbuPX+Rfl90YCeXczdcKn8ocx3Yrslw
V0uSWt+AJTbN4Zjwa9ujriWSU2ckNCevkRRtqs/yuqa2SphxCnYRsZ1fFVvzPnFR
lk0qsYCbnufiIIg9cO/9hfi5YbtBkwMJYzrOafHI7sVqRn2XQqQX5gT5mYQ6I3Nf
bmnFqutUPwK1+va4B+gPMxhVL5Ns2qkDUJtyZh+YjDRrA3kpHXHdJRj1WQifBGG/
9Y+XJwwZDsggLcVBerK/z4wjmK4Ue3LkcEyGw4iyNp2Ue8ykfqeSxqM+yvkC3nwx
wW7i8Gag1MJ05EWWeFIpE1HxB0RuY17uFi0DFrqh+zEULgJSxSHW+8TeUZhlaEnh
T3w0uMEvgB2LxJ0tyVHnzf1rWvG2MtXRyuz65IXQEPu+S7+OusqxFGuJBA6Nu0FB
h4B6b86RuRNaUvAzYZ7rcL02Tfb1tltbkiL+WyDqFQraXOxfRkAUmv2ibFm7UNnh
uyetxkZHaTD8kf/NXnhM/VY85eLD7eLDn5wI9KyL/o0lHVbQPqFiygM+0qXTfrws
mE1Ye3QGgejg+RHnDAdxfp5ZywnnqxC6d+jXEhiP/xMzshCxOlyD8gG7o/pcELS5
u8ejE6795PHBZulkuaNawEJkxTQEJ0lQRnLlDknYWmonbq9yjqNe7ziOmeJJ8w5Q
K2eMpcWNtgwn/PGwPwRTXiMBbJOD6l0Cnx7LF8Wnw7vvJ0F3BsAAIeuy3AabZGFJ
cIb2LOWSHI5vlIK3rK4AxnwyjWBmWLrAhLggzpPeenLuZ0pbIvtDDSlOvrpIkJzb
jr0XALfHbG50HQPvEq7bEel/8qmhN0g/yyJQpQFar7ZNDBMz3b8bdTOGJ6SIA3p4
tCYYdG7gs7Ka57AR7h7/BWWjOjgdUit0kmSgX15avhCU5YnlglJOJdwu962TON6I
Dhx6ePmCH+fi9J3AbxP4LSpcQjl11SYAEbp6cf2nSIGR3a2//C4tshK/HMbHTws9
P52aarGYoK0baWbvadt9M/GnB9ktyEnRrNujLfUGwX59yXC9vM8nfFtr1jHe5TPM
awCrHHVuXQpn2cZpDbB9SNlz2704PF8/t9RAjV0Y6xJ4jxmnboX+ZOxH/gq96JRx
AcTa7AJwCrpuOCf4mfVrIjGBvEIsiPgM7UqcStiOg+FJ3CmqET/XmbckP9ZjDwyo
ZLDc1Gjx4xKJn7r7P9qa6e3wHgfZXWl/8NPqbDe8dK5Xs+HQa+PMjezjpOnus6Qd
bsD6zc0J8MSLoeG+U/wUGl7hdBJDs6octgvsILHD1ehLL0+0U+gwHrY83XJEzsF0
xEsqzgRraFCgzuAwMixwTvWe6NeTOq7MZenQLqVPK8+o++Ayloaf7Pc+mVXMPbWU
/wfAqFbJl/UlBgVMaYSXSZ/NBZvw7CteaqenJs2hTvwUEd84j9KfYgMYagqIV84Q
WyV8O67GFjgkCrsGKwJSRU6Og4IaStdpQKWzxtEHCDOw+lUOX3/t5rBdRAh+cMk7
98UcaIYk6zo3o31gXw0kfYCT7VN7L1PauQeidbBpPxEYSTWfJxthzl5GSnmSUOPZ
4eEL5J9nq53tjEf58Sm61bJTvXCxhpuMvYPCot2bOVBvOsSZ0RJ7Nr9e3NOqldRn
/sKe5Ta8wfj9GjaVpWDJk464/084HK3za1R1cylH2J185hF3yKKJKCGEwPWbz2L8
scnZdjdPHHYxQHPfgaEFpXttOwpWvviv28P1FO5MJoOGKt/Khg4qNrgCgZ4StF4s
yU5zjJBWarFrEpL4GbtZ74Kz1xB1ptHbGqAGritv6jJQJ1Uhj4JF4otvPTLVXQ78
+6khUEqjnQCpxA0z112eB4/F1qu+r4s8H2puvzj4NazXNkKK3eFEaDn+8x2ydR2e
ctR6XkLtVyO5I63m67/Uv6TuEf6S2qis8JOEd3KycO3oZFWw4zzopyPFygHSCiiL
mui3J6jL5lIHJDbv8sV+VkyphrH3jWMblWIEY8ffb7DAtHIiBtpZvUEKS1GlXkzN
miIZ5281hciJ2R460tdk6KVqH9W7hDuIcEdhW3R/ajqSN0GbyZWeKOktbQ38YaLj
X3iwCTb9RP74MT2RC8Pge1rks4IaidPJ6yjnZYK4IR9TYKsp2z8JkkiURsr9trUR
iQIBl7RwuiL7KNNrIuhU/ClqRn6VWivb6zeoFY0RdBB3TxbUiDvRtNcGqIE8/Nd+
YtyVSBHUNvIxGXgbU2O7HrPhs7pw8/cAH7+PGQA2uqrfWk1ie39HXmvOvyD1bRYA
YsXcPaV7UpW0Y0ANUxjysulWtEVhq4BeG4a+ZXCcFTget8fDBDGpecHKpiJ70NIV
XI6BmFvdlM0rJkPIwAornePlwzxk1XFzyz708/tU8htziC/CmDplqE3tyu7FtsD0
0oA301DLS+nBE71h/qEkOgnZQKNkWd/QoBS4irJw/BHDjdctcCehyy7baIKWQDua
Prqx6At5+fBpYu8qEE3os3KlQkHGdBLkLP5nEN3a2ofRirc6NxxhL1cXSfFGFdMV
O8sjrhjUbUqHA33a5i3EIa7BpzRLLE2M0bfic2Zr4kdLwDFFRjNrYYdz56gkQDvq
yirlCKPRnx6Spm1WHlHiYNe1/FhcxakKruOn+rpQECfiCCZnksMnZcaDHCf/gAWu
sEcT+On8iFf+Apd5yyfZDfLQcQngZq+YIXJvI3x34X3pajxQrlIRPI6MbTAwd1K1
wMJARGaOtuYMoLq+Az43/2loVq7HK+eXNmwLNf8vRBt/NU/k5BxXIjdzX2qe8wdr
iJfGQdoon5FHwJZUC44kk10njewamYuXsPkkvFWN6zCYeJV4CxpmAMtMxvR14QIV
UNe5MdfYJ7ghbQpeCyxcVhTjiPlJsLEmI9o9b5mg1I+zZnT8DZFef6BwBGwjbV6B
q4zPC9GEYShE7GNz2VNuhtWlvvxm+PwmWwaFTAAhAYJPEh3/WRBlVmP4tRiDbf83
goVt1JPq7EQhHGSpf09GAgA5NfwvTvbofxQJ1BHR8aFaKufb1Xsx3HVQQX+WdlpA
Kkw8sKmk6LEF42/hGKhFlbBpkENvkf+e3ABFF6GSQKn5DeuKrH4akbOCt2+ls6pB
VJ6eGHY3fMqKFEyZ2pDL1Mqi8HP0x9ATnFQqLMTVBedBhFFP1gN6U5JVeOtzqtm8
zT83FBWGyZN8RtqCLOMCZ4Rn7xM5EScxx0ApJlMdH3kC7hv6r3u+t2xvdwaDX7Eb
5kGhadPNT9h2ktcZrgNmUNCvLS0PEe3mfVUog+Kk8ZhckVy5ZQHspeq5GAlrYUzH
MDiGNCFejY8e9RDIPOogJgGJKluDknrj2ZFyhQ4wIolw3zFpiNfKy9oqozOqKC7/
dWibabHR7UHGP1V8pJUb8o/yuFdcC4UkcDQtrXBnoEGFFcS2y8dtZDk+ooUVIOzR
isIc6H178JB1abhcJf9P5BJiq7cB4nfLLs2jUPysiJ8cS3vByUaJZfYErLF5maAJ
t2qlqaTUjnQVBSubfStOHvB9j6iYLHhLkZJu+59nDgA349OS2dnVQ/0aZ3Wxli1w
JKNroDdoLselMJfGF09gHXW/5bW58hfz2bYCxIWFAKf4ysn7xyiIYs+QQgp1H9Vi
w0bboTcmUowwXI1xPsvYvjHE7AwRCqVQdgQ/6skKbe7TGJeRzjm3safzlR05My6e
NnKk52GfV3ASB5tFxyeUyzL0X8+U1aMlUAnwPL10UkVzfMf8Y1EFJ62WAajmFbLZ
D68pK56wml3oxVcD2HnicNwqAZtXa1u2BLz9xDMniW6Ju2hhcCWiY1euasZy554i
9zC6qwsviluQStehMQ6XM7D7lv5KY1uibScGjS+QCrzVKntCj5AWqlkWK9jFSIEi
xsX4rC30PG5yGlBoA90kHcWSZdn4rfqg8GK6hwCWHPG/sAqXDBjgpnHIoKmeJcoW
W6uvlXImKr8wT84PRPX9FR8SED7ogSlLJuTFN/URBl5/twcNbdbkMkrm/1h5oWoA
JNKH9UifKtLWGzyVdOKXgO/Xq4Zj5Fz2efdwfjnnQLEMUy06/VgZjm8igbEejP+S
cmtEVFkVUh+9/HbPuVuNxIHTaaijLZT+PkVIuN1wYJxVxIdeAyPhTI3S5c1B0MdV
AdpUNGIv2dxWPII3qAOrE5I73O0pKpuP93X4uUBjq+zBlW7Yv3sFtCIft5n/X1HL
fzrYElZW1+W6XbI1GPZdvihaAJFCRbd1M2eyEPj+yNVjrWsde7AU5ItWoz6/hOsd
bszHWMNqFXRaSp+QCNtobKSJ0NTBo3dP3PRh4WzzX5gRXvX3t6mNx5Pd8b+9ccYa
Qq2TP3hpeG2f1V2HTAVxw8cdwfWzDF3cvh8QuVPbgc2UKtDzXIDRD0CSAVt4HrJj
YZVW2N8PqkPwZmK+8X5xbj8y9H6TADO3QAv3ZB5QdCLJ0lz8KcQx6F8f6Xfc9zh5
ksBCYi9v64Z8FM4x4DufFPmKoLb2RK4a0J2eAov6w4JyJqFrS5kKF9ZQJXwdFnZw
Z8Hq7TgdTOStxrksSQKyBnYIBWKSoDuJF+mXVr00PKh7h+RfMPnfPqTPDrsEgcL3
p6sm2vNDhoAgV3wqYIdIG46y4l1UzehFaN0JhA/KmIisawuOpsUZ6AT+jjcCt5vK
7zJwfr3NPliQKsbrHIBFQYG0FNVHLY/ubkIb3EiI+d1xvAFlR2pTSQwqDM9opKNz
0hlB+4PhVnS0k6g578NO/9ICiAcZlTyd8G/A6slgaIQC84AvLUU6UExUxKfX8c7x
+3W11POZtu/Vh49pjcwAGpqDgum380CTteIlQiRGPw6ExqFPp9ObWcsHfLq5eBl0
0Xf7ImMr1D8jDj7//u07rg6XemLXdqM3J4hU0W4uN9cnVlvFXyb5HJC0MEryKb8o
hWoaHAEbANkpSc0/tpLQgFNB4LZl79Ez/BUpZ5e6rLf+If1bcASwma4TUDEkCxA8
2bbDasjATd/hlCmr3b0K4YgJPS598MXfJXByCiaQH6HVPyPaXnidlGOvF3JRiMc/
KB8D74EGRwlkLzOJIPuSLyWD0h/QM+CUBaMK5Er6TveAZYFf7GQeNuu7Dp/wpDPj
1Rop1BND/HLL8dE+qjx42k95CpyMHQt2Sg06HXOCKuYHyIeNdlxfX1MRIy3mt1mO
kavIJ7ZKUnmvqugkf/Vr9/73QQxMpkR4hsIXwZ+A4Z0ZEiiB1qnDoXiHQjke7Ylf
lg300GrXfQc27w+wq6tO/14UbXVP6Y3m6nAMc4w2qb99kUpwNOhlkBP8pflOIt4q
TPaJjnPDT1etcXtdTDVoruZxN8sxOd8wp+ZpMtXpMZt5regMbawZVh9Df7uvKvdp
+MO/S9OHAwdVCeGTIiMor03/ncLU1aOqm9seJr2we0T8Tj/9CSx9vvsA2ju3dbJq
Se3qqxhftPL4Z4BLl4pumpkz6RFuAcntFtwTT4YXoQnQZsqnVcivn+e5StdHU/bT
Pmvv/tUARxR9Va4ueE4toGrtjvheuA09HHOcuULPY7hNxVIt5PV8VI/Q3/mLGz9K
Z1FFHnlrAUirUE9tZFVxKEz5dbisBqpdqiwbhIFKZSPgI3vu1iQYX7xgAVFySNlY
U2PJ2DiVk+uOh88ZzqlIYUEK1iPD/yu0ifGRNI8ORPnG9Wl2e+9HMkWQ7C3TMrQp
KqhQErY1T8+XJ+jMttEPq7Kv+uYiIIIm1OX9Yhi8f+MaGZ7g4TzhVpnc0g0O3mu6
oOaFEeIgDvZCK6ORjzvnjdhFJEacah/j731cQ8AkNDXS0bTPh4hfW1UwQ/i4JqeT
2MGoYTZ1dG4pZvcYQeY76aEiKAn+cTRUPLn79DY8r/hdVzmckSrJYe6Yh5a4AFw5
zPGyA9t4hnVgMqo044R7TOdvL5SyKzDSXjXKQYphatwPkEaEfAWvfp7CdEXvdg4r
wepuXR1oWofRMv1E+5i1+SMT3wv4PaQ4oXyuy2zdnz2bib143BFtgEfiuFGd3ptU
0MnOeD63rpK+CJDjY44ynLbe0dBk71srqiwkrJHaIFGZt62UF8uBPJ0EmMub/uW8
BpWcRRuLhZYd2iahpmHZCrI4cXX9sV8maA0fcH9eCyDEVx2hiwnzW7cDZD7xDVPZ
Yw2SrUxidTES03jj0bE9s3eoiFic0h03AGYRlyH//OhsaaZsqRG4Jd0nWgLNv5R8
oBnwq+HR7QB4QxWIHFNSFkF/komyuv2SMlPZZ4NwkkA+c+r10sBqrKpQz8JleS3Y
ar2+atlByZeUz85G35XGkL6Yd24W/L7529LIHgi2cfK9V/bR22vbfNjW4nM4IPWe
SMBlyB5rJ1GnIBlCXfZZR0BPi/JAA9K82D8Sm9NgooC8dZmQZhr4dCDoBUv0o7ge
jU8nWraxrBSfyEE10ZaZ4fLe2B7AdSv61ejgGZVx4+vkoHtjRXFz+J9ywyp5PTc+
PidTb5tlGq6Mk8FuqdXf8ZOk3rm09JQEHYsNlKj4NYjSloTRxq8dgvr6J0GeWw7K
Zrykmrzo7PoStMo4xevsJXZRMSi6YKTljEpcUhu2fw7y+yPhoiSsDkbH5vo7Tokw
D+wRpppNMPz4+s3mhf8Mpx/Vn8Wo/XL9zK4z6PnuEigu/iv48MWpSKK/XgLEYjz9
OU0/x8Uo6rcOrVr6nJkrlaHIisRXH3Udt8nW20y/l0BvBpmyfUUEesuoKJQCdWU0
gntxdCDCPceVpZmBbp5JBULvH20GSXxDHQJIIdvkUr0B1DTAjRhbglamf+FIPz9O
9nM5V5uhpOXb/Jak0aTpHUCn37eOlviyGsIyqJY7bmXvRMyvOx/Dumn0c2Y0UK2s
zSGs4unwZtgsf8jwYMohWJgu+0dij1THgL7BGTqXWXD2MPtkK4DjUw/Bcs9iXGc3
IlugxojD3qhnvWA6sDxQVEc/4TZ3DnTv0//lx1clq1TNRoBZwExoubdRkkP5GR7L
Lc67CGztveHTKPBRAZoLM/YK28AW11CnvTrSz5t3BpfejgfOrShf4NgFdRZeajD1
jrModJqncBMeXbY0hrHUd7e88eBoWulZZ6vTt3oKYcycPyoTnGuk9sDvxdvAT8wk
QcJwABPMlx5a3vPJIMagOFEkYMHuI+WKiyMlimkVNJBBhgETYlZF/kZmn64b4LlN
85ajgewjwxPxsmFrDC/f6XEDik5+V5R7v0AnJkr+NvjB+eTgi3x4rJp11bIfAzEp
vfx0UFQkrMgwyOYjuw0ydxBfK4xoeN3GNAO03AKOn3/mDnsXkYpBo64rzPdfWkc7
Ojc51GCN5Oyx9LjiECNQLxxcpVWh0Dat56mmytzQwKDnj2SheWgBJ/A5BJGNI9DE
uqhxXi5Ngcu8aVqhG9YnKlg2ZghvcAbIUuKUi3EGYOq075XQVaFldJhMaTb0LKDB
GjYZbwSgsiUF9tzuUrHXWeT3JZ7iKhhWqygAbUSLUcPIuuMmPHT4Pb9j6RncwPSf
mhXbwMaJ2y9AoLD/CPTfWxP3uOrFVLfNWHEcITQ007+Wuw+oeBhwnvEFsC/jDluw
YiX8qZtLL/8Gc5VrASpMWJLmdPFFQULlxuTWyYVGVjnFJ8rJRyVnVG6hsZ6wtlNW
vL4dWAT/QN7rjRNyZCBwBZXVtyGSJsRzoDiiaa4V3oUK35L6W6yNiFDPbWRwxGxk
OxaRlasVM0QKMZItNJkQodmdcCAwxGvZ4kU/3BptLivWcyZJHB/r0HZSx4HZh+xn
TdtUB8ltNF/cO/oNymXSP4MEVyCHK9quWQTfvWrB2ZoCIAUmn8hZTID1MdKMly4n
jtT84I1GvUBAdAyYB+C8YDmxcx64t75uThpaoTjkknS2G2owygfsB7ZoARoQ9law
/TWI9VffRlVi9gdXaw3PJxT9KShUWXQL8RoRT0+oXjuy0BmwRT5RS6z5GT66nIFO
73T0c1IUUfbIOPb7A8KC94ev7Yzt/mDpctj4tSXi2rnCTuzPrEXLaxr5wllacn9Q
iFlX+QhWcdtghXO08aRG/pC9HDwlGP9kEYk0Y0SHZKxRCeKOCLOHnxhptsIf2dT6
SfF02KWGQT4I2/AIUuvoDRqH6MZGEtQRzZ8ATyDQmTxsR+zlbIzbfcVedo/OMvex
mfUlfKWTra89XUSFQTrfToNuP0yOoumepYuKqAV7PlA4eOYVp1nNyG/oyEJNkkgC
lGjZ1lXnmRP9RsRUc059C7hv7Jne9hSU6dxtS7IRgN6qYJOGKhRks+oCFujMK8zV
mcHGVP9mDcNAC44vQmo5N0/wVMv2hrB4H9lSt9Au0Tzf72DpSPKya1qShQh6UACU
ZQIbvbr1BItZQ6krWWSV0i9nTbcTtgszAl5FfoKmA+Qm2qQmP9jm11w3UeFkMoSR
aacb4LFTWzEa4RT7PXqEA12m7jwzOhzNPK6B5dH7pKUv1Z4iZkHWa6dHqGzro4aA
3aBreOVShHEaN587v0FcY2bi9d0aStMPuVrNDnDhD0JtXhmOCvY674e1E90deYCx
NmTrVkbY3tWBT95zArG9h2IFZI3fX5P/5ofAHY6qeZOecNRNavxBTfa+3JK4in/1
Lg1uaxLwsX+fnpeqR+iK3zcpoLg4flv6QM6oy3s3OlhadykPS45iChyLr1dE+/Vt
BTpQFgWDuD5a7GHKeF9CV6mBU6DgB9BMT6VoYtiqUyeyk4X4PIodVTPaFjILplVk
4mJ98QOCFMMQk6EFA83r/x3nXnoJGVJRBvZGN+G6oVeE/z5aGyzKYHMfP4MRL8wJ
hBxE7wrB+azrBQBS4AprR9jziJspitCocqqVf68MqcAfWSX4ccHl7scLKg5ndyA6
89HiY5ECNJM+FPQ4JJoM9j/qaLejDI9vj/T0PVIsstakg1p9BSoi+rm2WW4esGuC
YAERvmdv2R5+tspWlfeGYqAiix/pT+kU1I84xc6AMWpl7ckrPwkHPbUp5dOjiA1G
e0p91c+x+EvKaw03XCBQ1pPYAyjiQm738WBNDZQQ4xYZ5TNnMzY5y+RbjA9IoMT0
RB1Q2tmrtwZTePp+JXB8GWnGOZL8JJJWQopeyghmLP2KbXqnKUj2+QQ1w2DHwJUS
YFCjFIVD2r5pFZaHyJ2BbCoPK3iCbUz62+gq4oSHcKK7zPORr+A6bO3iq5S7CXsH
8dG9ycs48ZVe6ZxDh+yCG107JqQgIG7nNZVqBhd+SSjC9Pxrj1e2ryUmjXPLetB1
LMSmz3sOX/d29037ceBlX+T/itEgm+XwsPavCFV3xYTlJygJb7R1XvdyxxDATkw9
tHm5eV5DJeDCgYxj4xNydlYopDar+qCOS2TaseUKluwsxE16CKcmbgmKZ7r+p4aG
mMImvRNBw813+1smT3DOdsYKAaJRJXsOAlpo41zjWVD0v/x4PbJ1mfza/oQY9fTc
2VcDLt1/sX1cpLN10tvWLvkiCECZSXTknrFJdQOcPfyCGXvuDVAUM+GPdDAekN8h
+mS+dSNhrfb+/i/TyGRCsUz0xi/+fF60mKm3buw27Hz/+15M/R8jVR3H60MlCEXj
YMJQ71IsB5jXYngST4bpu5JqvlQv995qMUYz05Ilzyo+BvcMXpD1B6GUFC/2qPe1
QDRSJVBmWQG7Y+gW1PVvB/VImPzeF2sPYvtSQdNrybgHSVq4vyxGh/6uXDjX2S/K
g9GN2cu2nVsHBwpdGWS7Qn3GuC1jJodeBkGdmbmYEEyvGCjniCI3OCzC9RnbELEa
G/Gnea58PzM2nGiOyPY7C0ax4uxBrGBr8G3KXJqWyHJ9UtX7f5RsnvbPHtid44Kg
aXca5ha9wH92Udv8WTW8D5wqUbXrXbN+rbKojw10AVYDPkJT6saKZHIMwcSpNNEy
f+8GtLyHotkWI4+BWQq/C8VB/q6/VkEJ7xCygKDON7GqzCT9Hv9CSFqDq4ZyEKqd
sAg1YHvUKsNvFiviXaiXIWC52PBci/mXUeUHBoi9AQ4VBxIRT4aukHixnduYgxjL
ne6kD54ShzfgxPF2hqU6BdoLi7Pf7e/E5Kz0P3AKZGqSECWDuxvPUKuIvGvqRqYL
NoAtABB+bDVCGrpddqsZuN5J4kfDzjBYEzVbfPF0aulPDguGsSqADfQNMYF0owmX
5KyPl0ilkEFvIK4ZLmAeWU2FsKq4HwN6wxmQdoQ4JGTurGQTeME9Cq9ewKv6I3SX
NwROwEJzvk1D1/lNQ/c0Bfu0dmyLNhKe5Zv0ld4Mbx+YIoYiXrfF9z8AZAFn2Lxl
H8i1Op4+qA/jBF/W5wiByzeKIk/Ad7bTJ9J24H3rOCkJPY1flFdkhyB0aYEKyWQJ
adJsWlTfvW9IRwjZiHBB7Mt//PD8RBvjJ8xqMyMdR0mouncRQ7Su0QVTLYTgZTXd
n7WJqQ/40V7aspGcrFsfkmIcx5eHZW7cJo1cPkEjUdEyfytIDS1QXY8GYuOCLfmP
pCrzHYgzuaVUeh/8oKXToThrQv7x3mP3DJzd4oudwxCryDbCcNWBzs1xw7AO/M+U
ghwveBlKIpAGvhX/V2C7IVId9RzUm+0AGrCeuPY2Dfph0y/Nn/9Ock4KPBctvPjh
Hw4Sh54P0+amHZkzjQjMXOawLhF8HZerYaju74mAUmuh9eLoLil1YPEk5NciGryY
IFw7+2rOqiqcgViH3DH6wPhGVgPccEGFTsAqREAyGt7FM8ksRiMuwJKaa61qfYkx
4PQUbB+/VR8DMOpkWht2c4MLJpENOP10DvHzJEEuRX7Vm+MuCTEI6p1gdUp8gG+8
T1czDcKvKVjtM77ulUEMgyUgPVwcuU9gvAMlUMqNOQXNqLJgctDsLF9A031rWo5Z
nXmYtHbsCnRNtromzJOiTI8Wyt6/gDp3w7XDu3uF9fq5VD/zJAWibjbLTLiyEeSj
0AlAXdXCanv7wLs/ClXiHwnFLqq8cCVn+emMaZLgCGFCF3tRigQ46n+ws0TYVnbf
VwHQyXkoTNwF30+RbGlKd7YfOfkcIxfWXxuD3eoRmIBhm7/pQ/fifrJwNjEZoxJk
CkGF3yyIQleDhXBCdGtJEcoGfj1lLmxFJ/N2ep1L/70G1fKnrDWHEzi7wVSxUfiZ
A/xHWuxbJGUEetHilzJO+uSvOj6QLkoPMbp9wqDdu+ouvrWy2r3+3546fu2oDoWY
oRHH8lgNiu6JLVfHH1kZuwAGvYezjSjwwEE2gOBgD1wdW0uWGiFulZZniGtDNkYs
X1lJXQQ/8V+VU3e6/WPx6cu9aX7GcVAGx+oXv1n8iTabTSBnO+LonasidPJaDJT5
oNwS14j/QmCpvmkX+QMs+lCX+cM+XU3qgbuzvepb1EHiO6PL/60mRPrmFVhrc3a2
ahOQqG63XwgXtjT8Sgc8m7bf+fXi1Zx5bH545bUzy7TfgfKWYDeRhV+zWkIsajAL
P+8/rDHJgW5eIdITa77ucM/oWNjYAM91pihNmbDBNDbZ3lmO5AaQO3LYZ2db1PmW
jbuPs7EOO3TMF5QF8uKdyg83pB3MqRv7vL0Ji3xqaRgyNscud5RkIgTfv2TxZWan
jIPd4BlAsUj9nOK8LfXHqx4X0m6PgbRq1FNNGkpvEgrQ+3UpXfPtfkgwqPT+j/+C
czpHmQidgCc4uzIbKbQLwcefwBfQ/HqKORre0Z86K0+6eVKpLm1nStv9dRzDv2nh
Ow8U0+uzuOJnc5+c7r/X5nuPYhuPBONASVktkxGC5/wNr3AdUP8Sog++ONB3o/qi
qXVu2u0xilqIgxgOaKWmbPUZDHg27Pl1wdMZxuyieQHqUSVuBlV5bBOEDXgk6ftJ
CMuN3HWs3MwLVbCi2QrB3uaf1rPMvKGn9Nmi2bQJW7JxUwYP7YH5JBx65PXt2VPR
HBp79JIiKmXOpCWNrVERx3YgWY7zut5/gTLs4CT7RTF5Mo9HwPv05Fcyki0I0/CA
HundhE4rjCr2UUdFWVLDGbOLOthWOwtAq7U9d2qmIbvak+9HO9QOP88/Fbg1BkqS
T0rROrjKm5dsp7vn2PxJhj85BCctUOnH4QuDe3EtSndS70EpCJYTvQVf/cXC0Oxl
mnhCF9zlydVG6RU75s70Rp3EvAtRWz0101eFxcGpfMv6Z1reuJLDNQIkUjc0FFcc
l3R+p6sVBn7/GhF1Y0UIGJIYbLzHWHWINsaCkeymIMc/JDJwr4VOh835gPloNKGq
JlcVq6wpEkL9NjnV781bK2t9J5V609KTvzOB5lnyKZU5Zou5F/wZ8TskhvgOUH4L
MbtqQNE/DwEdsZQcRbDC5krNf8eQQSUWhbrJVdtJe/qlJ32OF6sbfKPsd5hpoF24
lHG1y4Ao2a2/DLaryRMjOtwcgiZPJZqETasZ9mj1ugHqCdYPUv1PQSoF7v+gQg7P
MKoaJeFuH5jUOHe3Y/WjDDrxC40F0j+aH0Xr8SnsrchkusJ5sjiGmFpyf3CPDXFc
HH2aOpaZ7ySaq1wDMwMDNqV4HIWJY4jZbVHpUP4sTkPD7s6f11yAVKLI2WijINyj
Oo97Ff5gmzI+7wnvTq9MPwR3JmIfFYBQjlHQdp8042Q4VbiCWSDRLap/BuCWu95S
BaucIwuzfK3hh3Flatn3YagM5U6YuSrwBTYAS+Olet5RmnfuecZ0eYDBI0MU725L
SxNoYHh+9ns2yhmzkgsVo3welAy54tW2xE/k/LNAVEa0IlGVFhchTZaqZf52xUCv
e+iArQ4A3vcJMZkAabGat6J/66yURlXTdntTs7E206bvc8FVCTXkZMxCjKVpTvra
Ee46CMV3BDHdOjuZSNWkC5rhND8ehFP/c0BhpprSi49/WPk0PeQ5m0ix1gFvIFok
R0ewCrXYjhD6vXEgz5ySd4Sm6wptPzW9q5g7tFPLCthQCXtv6usd2mrWkSbCOhhC
sHBD/K0wG5yeHEvBgvVtmcLmnwB16fcuS7Gul2XPBGBRCegDN0QgAX00uTYXw6iF
hFP/rJRTg/qlI5nsFeWrDml2WdhHo4Uv2OKzgb4DtMXpvwPYi0kqS6FY30bozmoy
/3U3ExIToBlNiZLUfpJXd8m+VbplJWMZRZdLmElt/j1+8/kJnOrsV81ExzC3qBiM
+lUdXKIKVBEsle1MNFVOTD4woA4bKqtod4V/yZuMH0w9pZgZptOY5SOz/pn6owS5
7eVr1c8UJFCvsqdbuhBwXi08Nk0/ZBREJUuIhFF2swBcUnONukI2wr6nH58nOj1c
zfGH3s1pQjWlQhFP35iTK0CIrpCcZ3xkiS2q4IXSRYSdRr4VnkIilmWamEgPabT8
s8JJVX2ftzuEZRr0s5RZJ4Rzo3c8ID3stmsovfENEWQWtkMhgNlqHmm4az2Te0ej
lBVdjTGmXvjcYaPbBPCV8yKiHWyiLQQHoUT0PjzE4hH4ydrM7VCxp40V6FR0f9dW
Q8yUycM8Wah8ZBw9i2IeRCKG0tER28Hl+jdPAIBROafz4GA63B6XJ6qRKhDRBA/i
cjmLOp4fz87KkGU9cTtFWB1lqdKoQQCojXl5ZGY8UvHVqqDT+9/fD1eUq6Oblz3f
n5EgnWBlf3jq7kplmh/XjIOcepJm8zt6qJkk4XxfEsIKCbbxjUXzpDdoycNC2WXC
ktaHeDlAVNt783DSlurmZLeVrkxzB1jiCV9tPtGhnUuC0cN/ugmSRGXOUjwgzCLN
XqzM/AZMgJGFdwnUmtGhNgYJ/SHXkUpwr4ukIG0wA/r9Ft2v4T+5EcsjdOgp9tfq
VhiDohQWwTjZq5fzHA2thXMpZNmf0KqQ7/qt1jlckI2lYpKCp19XIqxD5n0m2sLj
G3+LOzZ73HLG/iQkgEhcximYxJmwCoOOgm4ZSrt6yOahQjjLOfRcp2y2wjn83L/e
cbvo+td54JelPMPGqwSYOLy9m2etJDvJRECaNlmmwdQVgiQPXDmcHAlFUHuBtdEE
Z5cQYgoE1SOcMdPc+VEZ+ij4CxmnhYPU/B3MMOhf+XuMXoOHgvioq0uPF10yddYT
LVxrbPdbT90NyTYOYM09RHEiXOY/qgpmYO0xRxhRpXtPSIuGPS7H6D3AS0INjX7w
sOfn+5NAf0g0SePSC7EYsorq15k4Hvclh7SUHWdkZeHpXHIiM5cp+m7MJuLjFbIA
IZMmW9wl7BiwzpAr4Hb6WmFJ2whvwX4YgFY1zrpitwp9NoxM1rOxpt2KCfTbi3H5
6YGAPe6RCP/2cAxy3fkn0HBmwPWd7DzhRq7hpx6H4tv8GSIRxU/GKoXrSd6vZz5V
tp5rlbbXIQJAHagJpWfwtvfuHh2Aqf3SjBmKMU7cllenr2iWAdw5QKiO3MJud4zr
8BVofQPKz1oWf/kP+8Ydmv8t19l2xQE+jNL6aVOIQi43D7k/d85WecNzV9dEdJS/
Q57YXhxKwzMIhguiTJftGlLcMH2FikdzdTn4141B7fyKgu/T09G875iwgtgTcCtq
3g1hwDJjrY3HxDIG4VnJMgRuPvsrW8Vm/n1bZJurvCb2pmrSFWfh9YzmROhOrixO
LUfA79RYMMzS9wjlLoei5t1zT40pky25RU+QlPDinEWmqkjA8KYjwcJ3Or5pG0FY
VSCppXrK0XJKdtO9upoBk1HfyyR2fHS2qjFGW0dbuV5g7+K4I2lROhsSgDayxYLY
Q1Jx5vu4OZvFQrE9Oz50ATR0blc1adA5YDUkkwM02otpkoA834HEJWyIfTC7xx5q
GkjAYU8QUnDhvei63tplJu//MBr7xn/JkgpxmliFUz827lwl/lokbecBOiraYZil
SJDPiKe5iCOHPry/kKCPpWNkD8wP/myaO3FM7XWrZ0HT/HD621tpzYSjAux4qwLH
ghjZykjmbDmBdaoz+m00nyf/66N5BBnHcoNofxTnmW90XLc31hKQzwlNk5pX1DCc
8c0mVsQ6S1BuSTHI4HjB+QAspp00o/MvXRr8/KzRTH9pdR+ic5JYto78owpqaivd
urTCKBfQb54KhJX2MvBQKQ2d2cE+3VUlY/nUUr7iLTs6ebVP8bA2C3zJtgqrTKs4
q17g+IXgPzsxaAxiSl3V54mlXV3zdI5Ue8d7i1WeU3RzcnChLpYLPa2K5IzpiFrZ
j3cnDY1/nemmhHFzC7apFn9Y2xCUPG29herl+EfUzClbIn3ifUqwXUd6mWs90Z3Y
b0XapC0jYRAWli+U80p+1aOGb129iVtndOczCRWPhLJBMU5FrpLbemL/jZiv0maH
QvZPNTWjBNi0oobkZEtJb/DDLxuA7/DR+7tJMS0+zqpkx14JEppx60EvlUoAhX8Q
coTsG95lHYPKlTRLMN7JWNpoPBiHJQzUE948IC4gCEDMpn66Ic3xkzylPvViw/tH
BY8SwyxlN9Rlk2xg0iJiiBdBjjf52Wq8QB6BPUDhdthvumrkI2TgZlpPvKjfQpwm
0pqccsOXpGPnkNgKvBD8rTFBDaDP9sxGp0qzKrfFJa6F4ZlVryT+8MaC620e4Sk/
nyt9ybsiED3cfq5RGZyxhwzCN2Rb7GXmgePsPvRu/XwxivFVoxdcNP7HxWKEGFfy
dcpLq2BdBEKvcqeJ3cUsPbKDZYYQg6dCAi0Y6I8jCX/wYYfLReO0PlUrAoBLgsZz
TX/ST65jGwFyZ0jCbxQm54biKuOpyG9kAV7MYSylyGzkTbxluo4TGAPhsezw+tCl
bJRQnmwpMS31c+7oXHSLvY1oOkMdRm7L2MwBhaMz5MYRR9PGAizgBNb6KgqQhGnT
03xG6mi20GkvqSHYVOFFEU3mkZjxfFFKQarwyqsK8Y4A9K2NonEiZFn9YMTW7JKA
RRmCxmgDX25hgf3qRSkk19pm4hhJRay/9w5nUVvys6uFnQEngdlHiiPMHlbSOaBo
dKFFsevB6uqeApJAEzXGMlYsF9QKfDBsu/2RRZnD+Sg3nW2a8ZiAvaRRoGbDFbsP
l/sIaCwVlTI7iYpem4b1biOjvM9HdOkXuRExLzBECytWwsiQIWKuppnmHhjBMs0x
VtCi723oNxLD33TWbcn2VRaiR+/P34z88mKD/I2aIVWyug8Y0117HO6J1zpI7FHM
AyLLaJfAMCJqqoAfHw8xrBBJhuDkqqADI3/vPmlOzv3GAAz1VAhIbPKbHDalMom5
iVqy5yy2Gck/Y3ZcaANo29KrqUk4Jc6xF0debDtjwtSDYR6dP54d7vTn0AoD80Oa
Tp+cEjnly6HL0JFpHzygeqPFKIX1igFnJCPJyoI/pZuitYrfrawA8fazgtiMkeOR
RvUYfW/dUKgyyvg1xkszaVPgD7+kaiAobCjbwHG+UpDnxo+P8pbAeGSMuUhNjofZ
RiXAULPe0wwIBBl9KJbF800whKtroOqtLZVOvLD4KJ6Nzgz+kG+fa/tVIJS2bqcb
zo+2CavHAcj2GlJ8ep675bOLIbRcaNut0j+V//8fzZC/C1b1yxnALLjCnnjOGIPs
8oCrTkszafgHB1IhXA60VDrPSrPjUcrhPz8YL3UqYj9TvIwyGf0+KO3geq7vV+v9
TemsuYjXxQV1/FIvF4ArllXUvOSfpMBAfdniYMGAsei4KW/vIsIU03ZqnuxP1VAS
MN3wh66yibV13ch+H0y232g5cz92ZNVqEHMgCewDOWQWyRl9KYU7xtLwFLJKmdpG
nAytjVQZT6H3oNSbyyZXJAvKsPwULSWspnkzm44cq0Sqt2fjczX/J65T3aWSmAIJ
d4CWvDXV5dHphrmvohYdPeRM1QQzcIwJhb/GgM9AL01lPMHtB5R+uaZiT5qni3P2
SRsvt/idnfl0vk4FzRaJDdDT97Owc0S2HAl+13SRpII6Y95clxGTdjhcIdjs9kG+
oyrwkgvsE0C5b6SHAyAvRTBgK5wIhT7pDI3TOH83qs/GCXaPBtiiizXpGt99JiET
KTVfRrbKI5WVQPIaRCCoJEjkDXaO9jIqKtTyrR+qHv9LIs3k+2XNyjdhEMKs/9ta
2VXYRcbQ+ebM9wtO/hK3s/wmOE0qWbzjpGO5REOLI+7Us7p7AAfVZEQFuoLb+8hY
hFuzuFyQ8+5BxUt/GVVTrQVL4DEuQmkElttPHak2eahK0YixaY1b5R3wpm+6plCH
bzbo6phI5iiVIGwWwqTkZzqLjLKI0sjtRwSjLV//1qzK4PS3IIvlbB/izPjMlcFQ
nytEdhoGavf9LxHnqiSoV4KprFmoxqhc58IQyE5QilS8mTWBpcWZ5rmYfvP2Z6/g
EQHkmo6bzh8fPfPf9xG1mEwh3HwX7n8Kuvl8ONN+VFCMYYBrfWQTNA2JwQJSDygh
Ybr+NWuK5VZHPef9XyoHBLmyhhMtjjipLmqHgmkLZSM/ozMVWVyxCIWZe/+TAuqX
UWld5tpAkML1EmL1xD4Zk4wi6SGdVbbF+JwwBbOW8vAIUhLDZ1L8sRs1Ppbuyccy
ZwT4K7mtSRgBNbQICf1CcYcMG8ZJrd72yfWYmXs6TM/mDJODe5MdHz8QArK41SmM
qsAi70BH1+OSzSC+PgJWoR/dUdq648v1bIqIP5/u2FD+t3M2bNEHaxKtSC+TqHq/
2Gb9zsA7R0qSAbpHfAnft4bcgr/5fXKXJX0ySFHnYkyCkj73t3namwOrZ4zg1369
WLjNSSPLmkoq2LiNZAWD9LLxIXdC5dQ3pEzHrT9jfKQ3gbJWmgGapejydBgFhPd7
YgJWlkkXh1apd1vQbIZVy5iGzeHmunbH5bOxZDjNfMr8JT4BmUQZDpD6DC8OPN6U
RrOFnHwTr8RxKpalNbNFLVjsvJGY10144a47AoBAVtyguqPj0DLcPYC4A3vsZ2dJ
dFeToTrAFm/NxWcs2qMBpQfF+URCtEOpMNVUb0Rz1Uo8yE3Le1RSC4xITMdsutwH
9rQuAcRPmstc8UAadipe2tfGDHm2FNo6irVKjVOGq25OUsI1SRLNeMsMr/003HrN
V8iuoBE9axwCa7EMpjMx+9SSXc4SckusM6LPBNMCnXTjZwxatagATf9O+DJnC9ui
nXq0snnk9NqW20GBc0HkXf46QJjd/a8SlMu9+gBqV0fYralgxKwhYMY460NLfHU0
0rHxdL0xUwFgBYkZmZfD+hM7Yzi6psxqd5Is3bZqLZbE+pu+x1IMbxoK9+vm64T7
hhZU7fww/cDFdeAfvycWHpJFodztAvmul3iEZATpu0OQNEkQw/ANuF0oOXT8Hmot
eT1lkDrNuutDCmwH22lhMhQKptpYpxqGAUnSAa/igRfUsshwDkhXBIYDlkmzpnjU
OpLoW5Am2b2MIRU0Dw+xzlUTlYdLhN6oUFR+ViKVj9FcOqXeSaot9VyEjnSka4yC
HlnQC864PD6ECAfIxFHlGmFtlHzkF2hpZXdubb1a7mrQF0LONT6FiGws/UEiggAw
Z2byX0B+tULbtYjqPxzuRhge18/xrhxoAnkqizQAXGY3mby8T97wGawCjsXrrvwQ
xztAgZ7QP/oTLvhbsBluqcu62AEAISStVRKfDoDYhSB7w5zHGNjnsyGhXX7N6gtT
YZSSaA+72Ny1cZ+FlA4yztNTWY0AaaM9LgwS0jrur83vOG4ESQysRbE4AnDR3MoP
McP/6eNh7OnJlu2dKMdzGzCVQoz/WJCFxUTL93pK7Bl2DKKgJFy05hgkfEFLDYXP
r8013vtkBd/mewjCeUONsxz/qjcYO/Bgk7LT1URa2IygnDv7ZYJwBAhJbP3FWJJd
CZuB9gdhCjWPtGjyKp4/h810JVObFMx4pbYFaArgmuEz9VfsWnFcl+Nj/vsgTDUI
VQnBgMzZ3xFh/jN/VCAflqjp/DZpuv5VlHJQp3X/31MdJ1gCt5CullN1P9XdBcSB
Q/yIecoI+gpSjXD/mePvpmFSZj0UXDlrFd7swyQg2uiZ9ZBqe57IvqMJnAyxdIWs
+MpfWaYGv9XHWssB7I5wujUGuCyrnGr9ZM8iSG7BmtLGOfo6MpfHUsANcKA4CGV2
c3KQq4xnzILKY+roa67LNc2dghceFrq6cDRWHjtmo1AQ/DZpMFDw/pOJAF2q7JhH
9fE1fs0NWvyTmpHTmpZQ+PtC8cJ4dvSiIiHyllrVUtSIxnh0hmRTsF59VWgNwEuD
57HBPFWirJk/hio4Ff2NK+2qJUMTqM84OlLheVau3IYrQmAcKqy34f84eDdiJwmJ
m/4/aecvExfdDQ31w/T1ME4u6VDEXc4KLGE3KWU6ohxVLOl2odSqZUzsrUSh1ta8
i+L2xDgxO5w/1UpsXOhAVWIl2pXP2RlkgN3wnPYI4qsH7UMZhaUF5qBXsN5cwkkB
0XKgdZnWtDImDjoK/mZn0l864Zj9gtd/QV9b+JOr0Q9ngKr68A2pGPAxnZHyswR7
mYP+1BF+xjje6LuSH5wDu/3kLEodmrqoM85NiDqGMf472gX6kUd8ZxYvCQPAoXsX
XA2o0X8wShQCJMMh1mewTYuUY00pvkGnC1XDCW231qEyRSDmyc7heNf7VuGg0ZuN
yrbOugCiFppz527Lff3jMXlTVu0411femeGPj5iYHT9eeKrAuxRw84zEz8s03IDd
nyhLfgQAVb/nI0ciDUAUfllv4sIUujrrIizRziFI8gCVTnz5oMRWkGOWIdD3A1Bi
UR5+WzbiU027yQyodBwwTyl2kBqgbpAaISqV1JTOGgbknQ62ji48bRpKyBOwjWfI
WeKesa2amJ0R7hDewF3+FM7kxNKt+AEu0goAuSFqO+dZaPMrdwFMcU0Ggkma6gNQ
2diMl9QdMpUAVIZGawtMfXqWr7QBGQaEObCaAvJGVoKVVGriRxgYioxoUXE9rFqm
6KbVCYYRiHJKNoCpgKR4CbMgwvuU2kxchISfNQKujAWLYQINLdjBWrYCSoChqDPy
D9/pJ98CNzQN23Ih3510CXrm1IVzh5DX/knTE7W9b8BqOMHkDp/fHeJoqr+eJRgC
KXDTnF0y5FH0zxZR5n70MsBN8bjRW1Yp1dRVOdw6EpE+W/w1KGDF2GZT+FJ516IO
W003AYHtyR+by2oMy/Qr9H0WohluOh7feuUps9RJ1KDQBUJgzp8Y2r6gCZVJUoW0
4vcHvONVAtOGTATd8pKBaV7JT9u3fZmaUIwyeHaMsFdMTWU5dHGc0evKaFVhOEb2
k33FmIfRKPjVcrUgzqE8oSgSk9ARosEObCakRlKR0xF3X5ge2LSA6IToUkywIPg6
LzdgSPHBfbjWBLAoNqsqr+Xa1/z4sKf9tu2nYiCzq6KZ7rpxsBcURKr7pxYEMcn0
6UKkrffuNGrBNRlOvgv2tLuRPH/NJiD9uJrDAvcNghFbDDBNAUtVGhgTL+EINCz0
JLclZAvJ8DHA/WlBgiicAgfPzG4/qo+7AnC3/NbOB+Rz7t7Y4rXxSey4kbgh5mMY
o6EAPfD2OwMWaw1zyv2X4lHZ29CgMCvmOaMHmgWOj6P2Lgl6wePJfO7E0dsJks/2
R+7J0IWEHR4gFk4b+FT0eDuS83bji8BOfRI8E0IfHQp+UPv0p4xNZ9vDkVxjo8Bc
XaaYkdWWIrmAVFfsBRBplCcbpj9avKv6eiVyRESEsZx4ojyy4trVG8xBsWBrIxoA
svxMnySpamb4W8zRr0Vz4FURbEiWH1dNblYPqo84oAAw2kMDprib7hPKGlDEOIbT
Mla87lPgJ+HZOjNFgFWMuqPSZ9Cp5G5Fb4AbnWJXTdYoTOPU9X4rz1ilKb6t0kNh
nTM2d0rZjOSBwsdDYP04pbguv1T8FHgZao93YEZkS+4LHk4pO07tCK+HucdtM2+D
GPY2l2aTqGP7TcrBvs+3BuclxxqPr9NjEz19X9/Xfn2vrL6WSswWXr2mTnc7HWQR
K0e08UqHVGgpA8f4omTO2F7SczYClPV6JFWIy6vzHe786T1iJ43D9/vHtAXgmq3m
WOut2Y76afAIe3vWDvfdrwuCG2c3YuWOOP7QaF97oW7XWDn3V3XnHkdRKgw4lnyd
zZuohpWtTgt6z34IGIiW8QAGnlsIdusDmiZ4fDJIJ8YLETUKmY0obGoC2Kids7v8
Iu351MPV0XSOp+gFOEAq9fseiBuvYrjQCyKvZGzsGRdytackjwWYd8MuPfg3DjnX
srcDBEt1U0LW+KJA2PKGCY6wtEcJEW6usVRx3oEx5BCavMCeOWb10gjvyC9k+tOE
f7vZ3DHqgTxTL5SD5jXI7+lfSsg2I5rqO+OaheaQsV/xgSIqfOVW/4ScvCzS4bWF
KeEcUt8J/gn15GJnYAj5bIQiVBWGFUCZ4pzHhVwVxOQEUVFn8vVLbnRLq+RNgOfc
NicJZd+ahSxE3hjFpjvP1Fo2YLw3snyU/EjObpxizrf5KmwFwKbGhx3/WlqEyOSs
5wSBXNzbw2SSsruem6cw/9xzOPmFsKZXXI/AsaLJyS6dK5yVDOW+Cx6mOAjM8InU
vvQX7vQlNwJTQib2AavBR3Bb4Vbqp4M3pna2SFlZUzG4ikQDKcA+7mzXwCvWSp5z
5/b6HKwn1vm/IEl/+3Zpmy5t40Ff0Z+vInuK8ztDbRhrcmQ4ZhN8B6qN6Jz8Vc3N
iMO7GeWdJ3GZG6j1ytQUeSxYXnqrBnu3oZ+17156VZdEI6IYaLZTvFTYa4qB60NR
+3hg5BgsuM5+VuUWaQcqqkhKZkWnIXqnW1cxSWM8hgcTxr7zay7C3dioWs5JfnRC
ccOwjcaCV2hGUQ7KWhYPK0hzhoQ0GrgCfsMKGJw9lgYtI4asUaQgrq5e1o9VHfHG
mQm9VRSXSc1pSElFTJ/rOarSPP/sz2eEMQmqIEgt9UxJTvGxf+c8cpKy1h1FUD3N
PjTpVPso2f/OegmMJVRG7UUSKxdM//e7P6cVt8DqFIauorUawWOjoGe/XR0WataX
r7gPye9RaGOJRLrX44hjikMZaNGZGaLcLsatWpNTwuIpeVfHed9T0TUjZIcRgHpr
rtkKCQr4glrS6Fw4pqmPT08UltMOJLouh69ouS7a+OBRWImcjZ3U1Bc7eqAskmfX
JEV0xgFyEd05I+x2p85iEiF9tij3kekKHNTeDabggvKbRx92w1c75WXgqoZgD5dh
PE3PRA3U19u2S1VhG04sF7CSbhr5HqNzdKEDDFuNp+VYWo9MRisoPt6EOAiQh8k4
IfMxkd1UqhT+bNEfrkLROX96HxM7cPI19z8LnciXlK3/t+Wqbf2TsggQbtOHpDB9
pIv+FWvoDIGxJA0roIiZ2M6Z48c+J1mzR9qmbCP/Z1HsgtcYQhGyo3M3GB717oCy
Wd2QLdCDDHxvjoeXqCCOEi1DjOMUGoGIIqjywzVvSkUh3XOnRJkCx7Lprrbc0s9t
MY4XPZS+G8/kJ/IbUO54Z3BoPKoJP3L7teBRUT5est7h4sI5vXtmCwVMEyZAlXZG
6Li4ztuQDvXAlUxbQTpqZqrLSKz6vJV3uW0qm6JqkFWqtknjg57zh8g8ysqd4lYQ
LsSkbVwwXnKsTMgE7I2lIX0XUxH9IrNHxKLFsq+Q3/KtGiNSmSdAtXnzGIEx4akJ
r2YXAHwjurk2Swo4xKZDpXwA+Np8WsDbwjb4mkMfZxsY3S0lPf05hL0uwplG6sX2
uxpH0O2MUxG4i2r3xqCtVRet9vIKAOkS6+JpYxxVFlCmv8ulrKKrhQi3tu7Nq505
/yyWd8UpQGf+GFtB/D4CuckiXMzkuUosvywdFjvsYVT3cnqUCReq5Rq0Zvyz6xV5
Ng3ZtrayfoLHnWFxnhaUBQBPOvsZr+sCp2KwY/s4+gvXb6hUrLtkzVXVxfRSlH/o
W9OVAxCZFy2U0g4eEFFqP0rSJeZJ6dpPTSc/p+w8jmBwgGGLig2B+mWBycl5l83a
mOg1VuTeOWBTDC0J7aQH37hjb2C6r/hodYK7l0zZvQWGTOEuVs5mXuHUV3MEA9jG
f85y5Ms6fnzTck5yRGm9QvJ6U5iV+klyzXHZTKj1DIIIrpIDvIqbt2Q1+U13x6mm
3GZzbfXzdpoA28KJoJGxT50b1T6F0/FwThKd4BSV10ZKMFuentWfZYOQ9c67mh7b
b2j5+YfU3CVxGryvGf11zapoXtQq10IWxOfxBQPKs2qSUDn8ga/X5/Wl+3lxkDFJ
NPLerZenon+oI+Q3nS3+eeqt8Y+3R0QPu9smPbGwrwF7vNGFG8fiIAY+K4nw6dlH
qrRK86aYBKn5OQWDJBh56Lh3tnYq5fKZHWACrdLbkYlIcYQbN0B86FD1wxijaDt4
+1WDvPbgEjCbKHPKNdrkdQJAFGPEe08VZ/GTCjzUbyQ3gjK6kiRvHwjodRUx1BId
iEo8jmhCK8LSrv2g9nWT+xvvEKA26NbrF/p4ZrL00gFNVETLoz+PKRt8aMQ4DVTR
lp+R/XSl6iLA+ciP2dX2phqq/+1JCvB5MOJJ/E71rx+J3O/LQ3leEKZXHZ/cP0Lu
pbpjuIWalO3NTlP6T5oL4RHKIWcUOzL7UkVmbhtxLgCNlaisaEX4aiUPNx5847f5
hni5qe9GJ/IFWEyFGOLQd1pEOuNs5q1ETx3xxNN2CKTNTFRQdiXLKLGFVOIztB8m
4PXGZ03Ie70KhWX1NmE8HKpXdXZdP/Z3gcg4p2HoTcC9aAGUbHdUMCsP84YCuYYD
5JV/Ndp4cC6mI7MuPbwapngV5wo0wqJuBjlGvsl5WdCW8/lBNNkNW/sLfHf5QNIK
XrpVDchWxbgKN+5oF334/rjRQrp17iF3euqkVueVmMuubblGR2s+Uno1gz93/z1g
YpHBEevEwhngySnCyPjYPsOSXxtqSKFFarOg+BQB0oqnfhDBIzErAHTv4rLnih90
6GulK+1zlAlxDF+G3Qm1s6UcOOTkxD9IIF5s4U+QWJx28LOZLwChYqP0fb70GEIM
kin2dZGVwnaRyJSZo3GQyKdhmwk7auMSEabnYx+wjX6OKHO1qgSlgsL/KDGoREGn
6o4ZuyO4nyT37tBd7NQmIkmvaS9dD5LIkF+4b1r8JebQQOAehDf4wHK+mx9ebe4r
bj4HICrheqWZUj4F5KXUDmV/eys3y6F3RjmFnDzvn2tnFWlFo7DC5XUq4MHwcAO+
8djKiCYHCbfmsy+fv30nhMy1yVvs6Zb23mfHhYhK3Zdbss233MgqSQ9hOTjXtP4B
3O4x+lW31hSXUoXuyeJ9GXp6orJd+RYop2UxuUapjFh51DEyhZeCJHr+rw4buLFg
mjkT5AV4MWRcxEJyGPbNbO3JV7QYX21F39PodstQvtR2qFHMd1l/1w00XFfVNuV2
30zzK//TE1UkgweIt+RabFg/n3kdmaQ3RvH0KN++O8g7xxFa88aPqsVkM+cEcJFs
1OPwhnjJ/riRlLJerHnR/mtTv9o/Z839BDS66Sff06CV5EgQNSP35sd2e8kbugaf
EsR8e/YxaB4jdwCtsFf+eRwIWT2BAffDn16gjCqNJO2HJ40FuAp5yoxTJZaEp3aJ
JSYvdQ0VXi6TQL+lAOt4nlIBFfNzr7BdYjpqhGoLOTlY80hbiUc8g/YWkyYmQUw7
+7RNEKGWIXKDBpN9UI0g311Uvw9gjU1T4B/25w+ajdSU0UImJ8k34Dfk5hcWUQoN
Z6Darg7y+o2AOv6sCVTdMiTdwpEYvB6M77WfSXO+TrQSK2+vGZNEAij4I4Clw8B4
pTa1wAwtInwerrr7gvsk4yKN7Nc2YDDyJw1wruDAC44yXbC2wpwible2zlWh3FFd
O4dnus4HwnRwpHjZ+M1nqwlVYkCrw7r6QVK4uJBeMHZ052APlMIEU7D0hGv5uCbC
AJIPL+lTqv2cpeZ7GFkAn5NdKRrF+BH1bEN/SzkrUlf0WvFsE5O7ha5rWjH46INN
81SVK68keF4RDYspNUXIjFlsVAanvn+xAuAnTmjr951nSMMZ6Eqt+j+GK1fcQ4v5
wTJnbE9xA6yV2Nho/ahOtmmlXYjvJ12loujnhsrDdgC4RKQek2Lhvr67TI5LqXUa
uVZtgjPBJCvitjh+UulNkHkVp5C5r6jqeoYdK7MhYC+tO8+q9Y9rB/8DZ5U3EA+z
4Og3ocfe3w1r3bDyML+RWXqx0bZ12jBsp94RWcHhVRM6STRh/w8BggLlve/Km6x1
MSTYlTRyxs4kNcZMg0Te3DGIBrdd8PyU0IbWM7bgPOMFKSnOo45+jfhG7kQUIzmi
n1vHb4m9lXZiyIoHSMWMvdqDawqMU6a4GNFf3Bq0ZpyoHvnjcqOcfPyHCdMcqJn2
a4nfguEc8iFVFqM7FLbAJWiHcdrUfsnG/rSKS5NWAOReCrZLddy1eKbKXR6l4bj3
90X1apYUzWq6bz9saWoEnbNkFUBCP+yJ9DVtjMEVYzj9MixO/XNUQx6m55pLN2G6
68KGaZjgbOZDXpO3eP9nQl7beay4HXcy55H7n/Hp2hKTbmxh8+cueErQ1yqZBGC5
nQqUWsJm+WZO5wmPLGaScmDqo/7FarXEgU5loxDujAmmLHfDlu1yvAntQNXK9Y+v
Pb+/9LZJHzW9VPhJt2SDpFggjVLLL3/EKzri/cKMg4Ssg8qh1FeeQRJjTQTlpCfd
Ky3A7D7dZGdVGf3/20gcNN1F+EtmmQXe74QTJwMkk3Hv8fEOmHjqc0QZN+JQPSnp
8bmT3TqlY+1WRxtMPV/re2IRPd4/elkphPdPfCG6X9GSDNArPdUX1/5MGd3Wes2j
8zUTOIaHGdyYzDs+WbW3pUTYjuy0u9ui4kTecNPLV0qaNv6M80bG39oFn9J8nX1I
4r/wp+E1aIumAbwap17NpmpJhuDyKCWWg90rh3PSHQEw/6gNLYBsNOXmiLmu+J8Z
v1WT2SIR2N9hsPXVT/3UAqZtRf2/A7c0gEhJiR4E7UnZ63tFfHpSGuM/rKNKwM+v
nkttzlgQjrSJHbt+kY7ygEqj42y1EHBy1tMBedV5MV6XIUMKC8swB8ZGa2ReOHzX
USgr03Bg6WDKz9mUU1C0Wfo0oiFvu2ZJITPVfYEMpfsCAJU6lP9qgBAww3r1jttI
DkUtgnFTSySmHPCrvtg601AAFUjVhHMvL1t9mkkb4sA6Ru1Si942FSDhdSJ7URPQ
IirDV89oTN01QW3KHk70xSqX0FJ6LlAbVoHpZVQnL+K2pxaZMyQH+6fAtKA7uUib
xKji66FfDFrqLctrNveUiOxpHeIg24EfmTqZKoE9JS/gOwf9hhIwP1KkLrjX9bE4
PmfZEJWxaSaCyJfiVzDPLJM/jF0lXoSqcWIZfSB3+9eyoEdXzd5CUdnzJ76YDT5+
YRL8/Tp/K6WlI0jIL/pis5piaAcxuUsc88fPvZZD1hy7HyBeuVfcZirjzIgqPpAB
Cr3YrzOJKtDuePWgAXvCQzc2uHLbbNV+21qOzurRFkkTOp0qfeQHMdmOXX59D70Y
PX/BkU3Po0zV79EDBl9kMY1AxnI/LJ4IY01vu8AbtdA3KieSyuB/u5QoyKNvF75s
zfHlkeUwxZW205WlBKJz7zEzeXXFjgUVbKhZnwliNiYk/VEY/EYCdJ5YT/8iFEon
D1hRF2VRcQ3n6pNd6Bunovr8zSPJD2RD+YJWh1Lpn3KBLsVELcHWMokFls7yGGN3
9WLkhbzwX/aznt9TpGynRSM19U0e2HUUsErsMrCzmmzYLP1lsL4lLPNrYS3vuvrF
8la8M2kpGOcpAPmxtkyM9IkP9Z/cuTm3XpgxkFVa8Zu371nLFdIN4aOrZxgNYzhB
cwGu6bg4C5U2KlJMzau9D3JtiLkLNb8pbEG6qP4YHAu2HgB8VrsEZjJMKyfaTL84
kEtzVNZs9FnsmQ1jt6pb4qlciupgzMfYO3DCWH+Ldyj1wJ+X5MMmVBp3wZ7nUyKe
uZieww+6UMmCQqMu1Tfs1yunKgSotxGM1vTm1arux8EY1ckcejo9c1JGXncwWdtd
UotJQQEopNWQT5Enevb3jpjqLQnsvlH1dCn4ljftTTvasBtgEdmmEmheadh3QngL
hc9Rrl2Hj5wsbrKCxuyAqsHnlyxnYR63mpBB1BKREEuAETr4rLDaDKXa6l3PhOVr
/FIJPBrghfx6aEgRSeWK7+Wnbb/0oCQ1bivCE061pI7dkj0fgTrHueS/fpqmYdaR
U9J+AjmZRVVLbYhy/olNRrXl62v9R0ZTbrN882CTIBeapTelHaLNevtT8fInplOJ
BnNhHexpvaTebJfF3AcRn+dEDMsF2ZCIceInoFy7nvZS78ELElgxDzTatJMYGRvo
b6S47AFWJMoD7kUdAmVjwmgJL8P1yyDqdGP0mdWBcgIjKwjfLQfj6m6dVfEnfEAm
+LJFatuQqVBat4hxnLjPWNNJFVX0YrgFwZCA1yaLv6nzI3yQZwLrRfiR5PxMhvIu
pkT80HygqEbXU7GmVRBRT+jsWtDa4sD2t3MYYddg225iPuBDUTqpL2wFyoe/h8W+
nrUjAqnFKwmByICBuBu83j51STp0BvEtn2PBvo8+zAx4xERZ+lR5x68+gHLxBa2D
VbyifVLKt1Ggj8nxXN88Xl1f5KeMXkkNxqMHJk02X0x55Fad1DqJAGUo6tt7GoMC
Sqav7A2OKczLCxiIHQCLtG/xdfGhsF9BI5lGtLPI4MsFqQOCQoglcXXdOGeRbPm0
AxzlkMGt03RfLJdTdami/I8xOkQ0FPRdULMB5RiGGT4kvJQHOi+BuwglMx1Yvl/J
AS0iGJVjv5e0Y9+o4XtLBjeIEwFyey0t0k/drxraxMyUWxRDkT84mpSIc4dxqQzx
nTkQunslq8aIwzTpz3v5nYl+qc/kf3t26iwmp0kw90Y0H45FUklokSz3GV/fySA4
524FAGE+vY97rWuns/0w2npf5VItd3u9N35tjWn9h9OR06+tizUVY8rLMjz/ykzb
rJlKlQXYZidShjTGdFYn+4eS45SGrl1mCeEpF5yg0ph+M6Fw9EUzPQ3cQiEbNcL0
W7bTj2gzX9ulBvNQPL5/u7vDYj8jVpnkyqAMzF9OOoVM9AxdpWCC55kyTeEcAmjq
HLL2qPVnHrTWTPbevqK4uxojTk7TynmvXWPKsYW3sp0odxe3p3NNGgh9NwiEh+v9
kX2J+c/8FvW+XR0lWzM9TcCkY+YRnQO1YzgWrZLQeXmGSEL3c9Srr8ntfpRl216a
YYnX5G8pdjE0X0Nrn8fkWhpolDDtC0Aas96If1Fs95SmWsW8Aw/Ba1QnxaOGu8OZ
4dHnJc0xtwovp/m2aIaXzHbtvKqL/FBYG6WY+kyD6UaG+SKG/HUubvEdyGy8ri74
rklI3BV+gZeNBKg8YJdWH3gLI1PJSN54WeGllLkUFFicujZilp1hSzny7QWrUY2L
JotiPv/HCb1BDz8zVe9WAav9W5SGiQS1yMxdrFemXud6e1fNeKRUU69Z9Cl5iaVX
0aAtOCu6LyWJfufPOlLI+mfDf5SS9WM1EnaBDle2JnbjbYuSLKolUfoWQtKxzF6K
gcA87gileq4ZLfI5UvlGDyj1B8RUOiXSONXbiBXnbBlWBsNXAO2uQ9d2mbz+LCyE
OAy6E2aG8PF3sgXgBGFLQEjnFaKf7NqLMIBMuVqh/kd0QDxyYriKCzXQ/GT3AOuJ
3Y7/fm1wyv6vCKrwyW0lZYvrrLCIATMt1TYEM/4n6KBLG945QRM4otb9oZUP7oJJ
rp5L5107fyA5YZ3X9AvASvqG8hKL0hyYQ0kMtuVl6Fx5ZXf3+eojJ3eSlGVq7D0P
6RDOIyhi5fdJ/7jM3AUXWkfphKOISDvMgDBGKWWrbo06zh8g0FGl85C0G2NoFcb0
A43cbSB125yBdPL8URn04eyqs2rvPqOHdEBawZW636rIeP/fd4eUmPWCK1zdHSa8
zz7N2PSPbL5TGoqCiVZf6yGi1zx85sxpdr3+yVt14QivVwzkjKqkTB/QUerMNEzz
7W37V7R4huNvVNNR7NghpAjQGKmcqBEQGtF4rRL1zEf2WhVHrOYSNEXPY837Z4lJ
yKW0LczDLpVYVaCD/d2aUV0Z+EA0efwxTEcDneqtjvSnQkvxtq2TFbt7BVQ0e0Xq
/MxVIq474e3vaG2Axy8tZCIGUdNl+Dx3ZFEAfKpJWjY5Dv1R8+9Uja50Hf9K3g7T
EagYmQx6NUMzJKWn8nHGAeRhNCp5bUECJlV0tCfM6Si92c0Km/yR4uxAx0f9f/VT
CWirQp9kYiqE/BZ/6Pm3l2eTRr+wmk3K6CYNNIc7aW4PChSTbFREkln+yHBLXFVR
Jlw8dlgDnfR6EkfoV8lRTJIqgCU9wk71qXderw/4xTRbf1XIPt0jLfyoASNCDtcX
tMOJ/ICYJCf3UD8F7ofA8YrvA3+iZOiCXPaVXQkJsbq0mYnmdx9Kw5ou2/poH/6H
P+G1Nk8+gCWAjvcBzUF5fqOP7cow42uE6Re8UkliSUG+mZfr8U+U14zsqcPhhVjV
jt/dOjh9fTwJMuIAteMAtsU1UKxr6me31fric+0N/9/Dmc3mJnGSd00hl93u85H0
rr4jzVnNVVxnQpqgX0Y0w11YW7NfBl8E0+XgYNGCycn4N9keEFUTvcDLTPGRPKR0
If8UHoWoC77VsIOX3eoGD5rH+KhBL1JLIMhrNyEAlUCWbby20h2/lNSmXe/McQfI
e0Bjbv2hcoPppue9f+etUI7XYOUwG542DZV8oa6Q/CeqTXssj4StqG5tdGTiKy2u
CQkqEnC72bK/5bEeuJrJHM8StgPT07k/atA0LX2XeKToopF2MUFQs06EKqq7OS9Y
wC7nvbuJ/PJPdsoWMxthZMU2RuDHicwH3zf4JQlCKMpG5OsResmB2Xktr9u7/y46
n3tV8HT8YsN5wVgm6NJdFIPFxgopjBtgnfnC0qUh9/67BwoApZFG8ZHfz0L9yDBI
ox/g97Fb5+pgIJp+FpyA+brAezH31ypi0ktmd0NfveD+LoVMYkK5V9Hmkzm29cza
nR4RE8NRduFA/eHl1UY65gxsR6mwzXdPjkYWHTfjVJDDx/XEVH6CrZnEDpoKXs+p
fTEb6L0txbfLzEVUasZsYagpKelmnzX5eTAqcYDfQLSAopkPJsAMoi+qkdR/CUFM
3wmgClBG/XYDRz42nP2qtWQb4tfM1S45tK1RoDZM4ypWym4co6xqhH3swOZpM0Ue
/G5lH8t07o8exV8vuPww6ljMSIkaA+xztf4q38AguLXTkGtvmHPbpslJ3A82uudG
zvI8MFtHHjaW/Kwxa7h/MHePLm63JJSJ9+IrtKy2pHUn5H/S1eidLfMoPpFmgulx
wjHAqpDcSC8h2o7tHW+76kLdjK0nmKQvqdDAt+LpLphEHS8DeORt/uKYxTn45VZv
6zduhBnYM3I/3y7TyOTf789vKDiC0wqimdFR6F/ysKa4Jkjfao/xdSD63SYN/p1u
+YOs+5tIjpWY3Lxs7IB0cQlS6hkRQIRl98/KjUYSq1xi0YjLlVsJsEJgMz91iRq1
kEiQsyK/hYroycSNap+omjEzjcZmJ9vtOWIe4nuoTq/bp3r3lmlR86hGaezMvoM0
uAsAZwWzoJuA1cH06IhjVtPNTPWWJ7cXFfGHA48MO9IljHw71tn766nHf5d9ogmf
lgD3kQxA7swhsLjgbL1cqDAlgzLV1fI20l7GwHXiaCC6PRzWA/d4ubMCD0VOmJiN
jaCwXuS4Jw/GvbxV0kMuMEXNllE1c1EuYHntFd5/qemLVrlEOie+jasOyISn7ini
gXVIKPVTfuEBdRBsxOvPIiq6YwepvpT0eVr/2OdMus6g+gbRvpA0xb3Kix/ItVv6
r7ZiQw/kRX+BBZR6XP5niJ3BUTeOL2V4Y0M9ZcdpC5EDRQYJBTn53xcyIKtdKXL7
EzuaXSR185zLCDmGHbC9foBoS+qehkgKVpp7NhgGnVV/L9KeVLfBrPJq5Zgq1c9m
DKnYpVjnZuqlVZ82ZLwZYdL5UYtkW9TFK6Ci4dvemCbf224FQ1kJZsCNjHjvHTs4
mpwfHnyjnMnKTu7dNiTw6d+AVFZ0t7tlkxXKBOnoFL1b3XSLPHyvw6VpfKK/IBL/
NcuXDDT3tc390lshLciqsmCXA+Rh76n9Nl++Gt8I8AO9DL6XbytPUBqtlcRDyEGT
eidFqPurKHCTeLMhPpc6damdBIvizmKIqaThlUUl0qDGmy39KINhTiE0Os9GEUUI
u6NJb6HAtCnEGH/uwn/T+S+zZJUQW//rFADZGckwJzLOeXjy5HnfuNmb2EgOKBxB
C40WvA8CqeNoPTZF2PK0oQ8oUkKBV1Cf6K1c5DZ2f4uzJkY9fRBVXJHefFQ4ubch
JRA93TaCGX/Ezw7bUkAOKPn6wwD3q49RdoidWlHSVVPLJiJv96KI+tVP8z9DskQm
R2t76yI0ozIXeO/lYEqEDUBMUc71RHwo9HnLb6XbP8Rf+ufyLcZfqffYMCvqyoxr
JIkVcecNeK/5kQH49wxbATYThrBlBKFpH/wvXwMJEMaUZp8nSBUv+GlJyfeVRsK6
LdsJUNtpM4J/S6JPcWymzqPJK0qdXKACopQqoG6ppE6TjY0LkgG2QT7bOaXJy2sk
CIZu6jZ2Y/YJ/gJxhZUB51NNqMWb4rAvKE09pWBrCvr73Rxhj8y0r2gW/IlvKWNt
/6t9bDN62Q+l+8kBKwf/1yi8roadIGppQGhFwQW3dTpWK91auM78eia0NT2kzSyX
e8Qij8WaE98Eit99YEgVSqCUu/wfH8jC1CCqX4xUNySVLEASzSdnPdbe+Q/uIsS8
J2+yG6Z5AyCFFfA8lHP65X12a1xBUU1NKYMGC0+FVCnLyjewAvmLJKG0sOvfILVV
M/B0Crcnza0b+QJxaG+8fPnwyTXTztKjm7hCOFm7o0/tegiaiq9aKvuvXrs0PO5d
n27iK8J0NW0kTedH2bTojAKz6pOBhcEnVhq/ddQJDMXHpLcLkxvwKWZkCT8pGoLe
fprz86Y2DW96wTBCLtyZ8x8iMa3E35i0Ct8CMz+ZATefn5O8souR3jJn1+lfuewP
Cai7UEWCVXpOstMdm1R07ohYbLhDKlp1/j3OkqmMUrWG/od5CfzV8bfurjQMXdpf
amTM3sU2JafTYknJFwpT1B4+5WQgsRyUsxpU4i85gN8NSK7OYK4gv7shooTdfEGs
VGkmRVwslN3D6lusqLA+VpmCt4Nga41KqfBp0OU/ucHxj9+DMAOkdUv8YcH5pXXM
TLH3ZX5HWdwiosWfdKj1sIJJZQ8HRclw+6l8ljyOJolvppb4584ObeY0MqXavsJ6
o6fU6DnCLhHqg5hdKiJdjAGGe70kWnZ17Hfp+HHEGW1y3yWazOBHS+ecTfLgbZo5
644dQz78BSJBnge9yWzgr2R84+lXDrnqdWKYHC2Fr30D7IMcC8AmPuuqLV2Qe8jE
O/xI+rpo1D6XGW630Ql7M2JnxXRD5e01JZJlnZJncV9KeKJyjWWyxkuVd19DijW8
eIv317+if3MhQ7VIae2iL4b5fk6mCeaIB9Tp6h/stJIgTIeTgDe3GbtXwfkIucg3
8/oa72JcxocDevlp/pIhzG9MOQevygUc2KycFVonvdEl3/5euShnmpY9oBXkFbBs
lS0XVRWc5/7KIqQ1d/SCd461e1tBn39qpM7ujlFKDE+5OxX2BWXGOERw7stpMxMa
J8mUcrvZWQS7K+sWTq9fTURrMJr06VGK2JG/AlsOw/EZtqMCQ/S+HW6oP7TrWZOh
hy6uotzjhrB/Gk8/9URpfZ4/ywaPk99Lvy6j3qGnXoQTSHQ1oouZtae1DwS5VHe7
enXja3br3dwbAEasYpwzJjdMGtQSrDEs2D+lIH+y9gzCvzQgglzjJ4x3HlmTjxEu
wfuHUG+iMzA8W05Q5dKO+5G0nEa5WxvYkR1IM8z4S0+9nhDk5kWvfnf22ifzWMsp
o8qJSW+JKqBIEBBR+NNCTVuVdrC09Jp7E9fcXfLqxXHgdS6TUGIYUQDgdCq6wXS5
F2eOGEsS62AFIS21Apu9rrlVsLn0mzB56pj9rfYfKIbW/wdXEaQ4WisuV/CqHBdb
5jIhtNjFA5vlrCtiZRkhuQpRHyREnocUyc0rHJvhNCsxym693HoDBtdn6d0FiAKf
e/gCtdVl3yvRbvNnL4NcYi+PbPjzlNrGOpjiukEAHj1i9wbg6fiibF+j98es+RSM
x0ZPz+DLQ3Fy0UzVMxzwUIPh3D8g1UtqW1jPIWtDGz/5UxbIrcup2UZqLhT2oscc
HYYYD9+BbFOaUIyJCk4fEMK5nqqMG+wz9S0ME4K9SjIOoyROq+kdtcHMjMxwCKhX
UYTv2W6Wqk7pj8HVq64MtuPepeVIvySWdVLgobGOQpyWGRTftu0qAnUJpRiKuAQ6
oQ7JD+iq3NdE/2FN1cLigpgbFO6HJKEPF9Kb3qT9Yj7ClJOKGxjhpAm7jOOGVd53
iEcCLB364xaaQ22iJDxyg3jemGGY/6K3TiHxT2Nk83/u7HQH8Qdsy89IyNuGxSMt
UNaqt7U3CrrFEgWXjEs6uHOL8A1RoIziByyXB7vIZxfvQYRXZfAcsBI8gWS4nGDh
LaZhq5JPhognNID8RZKRhWnrHt76X4xX6ChvlDfBEiNB9lMFrh1pNY8+3KFf0+zN
mrV/013Gmdst2XZnt3DZ1eMhg3Ti+hNonH5mz8yN+rWKfAPKYIGyRmKhAi/DLg8Z
s7/Hz7QPK3Kyw0JNLnub24N0pQ7xTkm5cT55N4IC5R4S9zOkyfQCUEPsgjs0Mvgj
qHRwUeagLkDgN144u+h+WD4vvt/+VM3qmWGdvfvqRX1WH/NFG2n6uamvSmHSB+He
KjUYOyuyrQCmhNHi0AAEvU1OV6u0M95k4PVhC/x0O28OeNSicaTZpcou7JZdRzqB
re31mpW16YLQsHdR+KG3wmoOIhYDQyFT9eh16AcMXNm+gVFrKC3IeFBhtuaUXJAp
R/HYJbizS2PfQ9p7UGasQB30xmZalQcJ9mwbKtDkj2MFd8vdsRhIDN4jcFjwMa/W
brYxQbLS6qHpRbSXNy+2yqGSHoXf7K8Dbry4ELFCC4rhm0T7BLnPGzPUWWrdssXI
7eMU/IVYN1or6q9aZypql1mmGRsqCKnHPfd0DoAg3GotdtAtCjp48zHG6n3vwTf8
sIeVvCYzRPp1di6V6bEtPue4zPm7xG6OR0rIzLkcEuM0oriPQnHZtQQIXBqSdf6s
vhT3w3b9w4baLNIAYGPC9PWHAHBa3AO+BffVdWpdT0O3TqajalOSZJqHi+FHUrK4
7tvJv8o0U/+Ql2ukTk1l8KAfD6BlOIXyjK+bmkM008o4Gw8Zy+SOBFAiNLOvV6A5
klMjrau8zo5GyavdDuNr2Fg5G8XOogj1rNbUumtYlZFBem84RW9ywHhzwKQ4NDx8
`protect END_PROTECTED
