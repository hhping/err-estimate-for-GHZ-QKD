`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
926smF+TopV1aJprMdqY46A7LLG7jNYtQ9OQvNMUe/jPCPTT+s+ulRnSF8FSd7VN
d5UWVwjzEryQbzcUMf+agZWFIYnSTsKfDFWbZ6ig1QhpA+GODEZlErcGxwN34Cfl
6gLhjQDyHco+eOtBVZzcHreCVCEZPHuhb8qJnXC8cw358NTc0degArnDJXVR2Id6
K956le+RfzdzvDUQwXQidr/+zDKkgpvlv2ba6ekwUN1kUmBOiJLkMCaNRYXemU8o
3uuAA41i3eRBMXc4veWfFYB1fYv/5SdCw3aQ4nn+/k9w1oRV/FiUDLYo/aRJkBwv
2/NjhOutCF/cVZZ2AdA0tO3oOy14tJqgNJNL62sRxhgG+/we7V2OHIAj5bAWwnxF
OLU1amtIs6wK/XAWyTJ1NxQHXVIl/OFhOi6tORefsA++tqGMiRfTlyVTYHsd279P
ucYLQXemC34SLqR6dnWjq/CACKICo7l62HC+ETza5QfqtItINJmqXCG1gDGfIGCP
FQqPCJW239cS6mwVgKCq0qjbZV0yguXcw33TQw+ZN6eOZQakxCrhL0WPM4aZh3AQ
kJAM6MnY7GizSrlvTeYW2h1FQsf+llnA3PtnFc5nqcX/QCNXTrUU1K2m8lOKXPtu
PxYtz4zlxOd3InDH2dXq8gXvpa0bzKubf2Kju2UL1qQVVbjd3FNzx79K788KmP0H
f2ereAaK56xJNNX81Pvr+6VbnbdCWSb+Aeigvf9NJ22YMMCD2jwxGBzpB4CkdLg0
pJJjeSQmIpzzAoNPsqr72KizznzA85FBWSja+SOOf34NUtG+Y9220z85Xv9iVNIF
kJgD+q55g+AC/5FJfc3twGKTqnQ7UHeh56IR/ES/XngHcHb76Wo9aWPiSgOSf2in
DOsvA0fcFeLVTgOo5c0RmDkzRmrjzq6g+6ngjUnsyJOBP/2IN2WkqVaGw46H/aO5
ZKsKSF5p1JP8+cKEj9/P7a+98ytoEr7Uge8f5752cgzdvEXs/l3nf9miWIFw7Jtx
pV9wNjvVnpLW15ehgu3nUIKcuQgkN21VFSZv/mLESy/3aCpDUb1qIipUm6ABi1no
6F+h8xrf9+K4bmI4ZUCHfhOm14nctYthy+sCXmuezMoKd2L57jNU2oTKq8nufrPa
cG5TVPbTAiN4O4ejgB30OyepKbK0OlIZb8jN3gVh02okjDnadC0wsWSLGTCZLwdj
Xh5Mnno7ZwQV3rs4jUyyhueci383ZVd5lHq9ev16JKaBltVGdAScvIjhmhs+0yQr
y4XXWxOwEcJ2PkSmAsUuLFdhmKTaWuNOsKBHCSv6uQY8dKgEwjVHSWyUD2n8XGN1
Mo5qH45OAwoBWDm0//ooaPCChdHnWoJuBok/vP+Ea7idz2ZiYoZwqqe8OBQ5QUAH
AKIf2izGTyhFz0KA8AFzzVDUpk+IhEN4U08uxqkrmlpwnqscQVwwdTjWxDGO22L0
dExBKbnzyjMO1GvMTrlIUnHGluKuEXVYU0uf41nve9bHYylukxUmuF/YTjvc/7GR
`protect END_PROTECTED
