`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdNtVrxdXfd6V/GSzuTTMaH3uWi/KMFbfZVZgvqUUV2QJBi+fCXL3JcQhL0vfyUy
Uc9J8GyoKDdjwWU4TMJ4Sh3znKmKXcQSMNgcSxdZ87FltHROv+P6Mx4kY0Hl7Dmy
cNLvMbjbJenFYVEo3mf53YCZm+6XidzZC/yEdQFVj+Cnn+Q2TU9Hrcl59S5Sl4D+
N908zcbGKXbz3Ahr+t2eykNiG3FkPUh4ktPM311C7nGM6f2USKjbZowD3Zahk6KE
jkFvCazmDiw1EexnYXqa1LQ/P4fFlrI15oNsU9v8JUMpdzEOEarlH0TRYCKVczLD
QIOBEQuY/rXYhbNgF1599tmqbTZCkaa2aUjJkn/IIyhNN/Ep4PFA0DwW27H3n0XU
SVAkLyfkBxZG/ZuDxBZO4AfvfMbhNM2WXQF3DOAeb0iMrha9Tgm5k7wTFgxYJrLo
zhUs2yPhj9tNn0FdNF/ZOQC8AXk5pMjDQc7Gm9nRW3MygBy1SEwFbuWMrJSR9meU
cZFuaq800zQ83Iyw9o44GzPfaLoJD0ztt2XBQVb4r8GIQxpDT9HACxyvm8s2BJHD
v2yO7vEZ0m2JAA24gTVjd+z53zxB7d7AM975dTKzqXGYKb2wANqnJNHswkiXn+1v
BfrebqR5fyUEFEnajk6sc6YAZB7UFhQSfrTXV8DV76vm/dwBwdynAzHWZBGZuGlr
zefuB1rqncTUUW7HkwybQlGFBpcgAhnQdUdWM/JcP25zlHMZnK6FAe1Yn5WKifRX
erDjvlk5HDAbV2agc0bhOBZA0gL2n0KVUGOKnZzSh9WOdD+FF4B/EYkDOZxcKggU
bIug7OfuiJZ6QROcMQEoEAORF5UPThqcVgiU51fgbdfuqP4IsXdRpwiJWopSIckO
e7QCfPp7eqMet/D/rEVFIH6amq8/Nx75Jzm34RwE/59s7Ja69/vrQG/Y1mtyG8nq
2gx+tpS1352iukeDeI1+16in6B0X7kRrcZD1ZzzrqECWeKCdVVrg/cJGd0txReeq
3vwiLJ2t2j6LreH2mTnkAdWevY522/AjCEpcVPz4oZ033BSfy7K69XAVRImBdyi/
Sd89QelWqySDbmgx/TUq1Xmos72kz7ppkZGWdVaSaPz0xx1++kK+ykO0WhfbOwo7
74PHpPYUy+9GaC5uY0pifN/FyfVgSOXCRyreS+FlSUr/Z1qV3s1qP7g6Z5vk1Tr2
1lblVM45zBjnIauBAj6+Vcd1qR286Z9i+dpLOllg5LAjRJfn8ctSll5Eo9uRP7tn
1rkyKHvejO4xzBoo1/BaxtCvgqwxLiYUlEShuTv4lx87FEUOBRWPjyGHL2/15SWI
d0g5Um8kXHujyF8v+4s+Le8rqmNlxceDNxplOZCsEEpF3e44atdipYB1zomGQCL+
iBo3EbwBsmLoiNP/0/gsaflXguTijTixMr2uPoa/kqBJXPmu8EEuieX66TBbXruE
XXM17FgdUJbn+Dd6CVRy3supEg2dckHHAECcbABqQliuCQn+BzbsyNWtexbsL3HY
WCVXmI7d+38TgGQrYAP6mh/RcADi+JbmNXmkjp1DI3kCJI6bnfcYCotss6gLo9K9
H3H+dtKixRM4IKg85Q0+tgpLLo0yLPcX2M7dr4FAWqn/a2bpFMozfkhZ9kRF+tH3
`protect END_PROTECTED
