`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wksr+D1Wfwv3Zn/Sj2pb0xI3aceLSE2lIOweTZTM0rJym+2fg2dG2kXZ/njoib7C
NHKrKDsrt/6fwK57g1Fy2I3g2tTfyj/G/D7v/oJWjuikWJ1L43LVUGfPZnyn87iT
TdxPPEg41SuF7O5LC1SzDxW5s4X3HsnVVClujviC38Je55Dsna7g4Oec+XKHV6mx
hkjW5U+i/LH5zKBOkgUx844l+iHwhvAqC5w/RLBVql2gNkQy4/NWCVtgfpQSqviM
rpEjSxeTcBA2qKqDLrCt6N9HsifNG8EfjmtzE5BDJ+ABNlj03NCRQnL3xliOPsd0
ZLhrV7Nad9yScqtIeH4vcFOg+13gzXMAawrkcPt98/+dIJlxuMcZ1UjEm8xZOziI
7qNShyEsLrpx4b38fj8E7abRTVAPkQUiH0U3lpdJ/AnkCh/HCxWevwriqU7rvSWO
vLKETvoZmBokONKoQL2P5HyeV5dh6R6AokmOZXUZ1eYhm8o5wBfFdrz3T7csLxAN
IHHEKZBieg7djvKkqR+8L8Ij9kR/gybyN3gELqZ0Qs9WDKmzsF5tWxYJtBGbxBaL
FhmX27vjkGtAa3UcF7JV1Znm7G9P2pp5Elc/nkTjFdwy6TLCQAUhT4KyRhB2uthK
cPi7DDrgCK5X0hxuqRYzjClVHrTSqCWY1iBARtcqXUWbfDWvYSDV3apOASd0T0EO
pLOd6DYcQ9QNEVd+P7jlQzx6+NHWVX8CMvZfnFMJERvaNuEsAOUb++moUC94Vwn7
EyXRsxPjsQ9jiAjurQfVkmsWtp4UHpTh+ROXJ9Z8JT+p5+zjYvO922InKxJMCuCv
Jb5jT0LMLs31vKqmYqpfBP4Y1i21Iy1KSrR1h9GiJHGow2u4rjpp4NTiXaKjumT5
o9abd7Py+xPkXH1cbVBovQ8n7oZDqgxQoo/XmLGEQ8a6Ei810gl0rRQJgD9Rf/EY
IoCFh/x0p+ZEuA7/5a9Q75ZFtkHvWjxfU4EPBaC/50kuYkQGLEbnoMqlMEyP1KRY
jQBMhRs1c7J7N1rredg7NON4avVjGt3+m7TwvJJ7zriWqq/ER0Tz71hTJFdJT458
SDLR31Okg7JU5z3wtQJGs+/A4HBBOPLoTuydjcVPraHe6k7Ot/6lYMQ33Y59V0EA
1T3W9OA4YYPP71le/2EwfiyC1G/atLyDfW+M+jlFbpKUZYbXOcBKtmaBGUcQBm+P
G2yo3h1FE+tUfTcmHDaen7vr73z1M2wsPPTHTc0X/FW70fZmax0QTbo+JzDhiPbx
YfEAOWkzIZx3upzbdng+VpW95zraSUaeJ2+6YZcoNvnnI9FYPfuzis+mZOoKHnDq
9K8s0UbE+mvdeKuuvcItT6F+9k6c5N92wBX9lMhErHoYrWBqc0n1HfUdoiRwPeVD
aqbQ+L1lqaeHeRJfqYS+btuxhQXm/gY1osv53wSPu2aBaw76tDeXx4ciePUVIqev
31p+3sRYpV1boKJ4wVwJgYjy/3UGgZ3mebFSm+dSJWerY5p1ls0Ev6u7na4GncAQ
WatomNKg6aKoEzivnUuW3jRyt8eh30gcKlCfvLxp4Bg6KbrZTTFx1ZDUTNcyc7zW
OGg1XsN0xO48G0tMRo6E9t1PRi+prPQClnlK/UCePZ+OQxqThZoH1LnYEW3ue2Vn
eLcVkWIX0tBCIOXvoovqY1fCCo8t91IKSaOlUOUwPLpX5AIhS1sMkhDz24L0cagr
SIHIrK2gjJk1TnrCFvFlOZhPbV90AzPaPssuzD7RtF+w02aW9+PsEv160QmntGYb
ZqT8v99mcbemTFKiO5b0ViVz1NIfEDf+BXtxUHW/Gyy6x5iIfUyvg4U22ugITcdT
HOnFqei70+og/OXI3ZKRGYNzB2PA7WjBO5Da42/6xrb7UNpKPqLbz7S1Zf3umKUD
2HgvOaQ0Z/mMKsa3wI0d0KQmt9pViv/5EU1bcoJCrd3zWvSR2qZCz8DpkivfNylO
cT9tQnKP/PKEdlMHd8eeXWM8Ho0zcqRlzUarAYhnLV+s9kZo1En9r0vXyXyzqfkq
YEJapkk76T1WxRAo+PtuBRj8vWM1C7rGAdSxu6+zy+9QwFEex2JWvHtXORtmJDu6
Q7XQEIhdtOaW44buLYIEzEBqGCfMIhOMAwZjiLnnButtd/1Y2zRqIPoQU+NyTooy
WLrjkSjr2iccFixAwfuD71U1e8Reev9aAqO3HnIkiusLclI9Ndn49XxJK55n+/NG
Y+X0NRBPlPUgbDfztzZz4TKcp4v/T9xDN4NzAnqdBSr1aAkE+MDCUQ1WJTq2QP7t
voL+7AnfARqPQuj3+t2Sd2QCW2Sh0dFc3Eksq9R0FPxvjXf7MKS4ycDl0V4HlQTa
l1qY53gWxd7vILMVwpAlKTokqiCZYgS43MlWDgWQ56vy1RvY8ntcGz2EfMZUcHOS
TEk0fgSAAHjlvSCTQlkAPd9C+bM4pRjyJ5esjeglAviv3ScBVrifpieQ2E7WikRa
mnbXatP1WSMljYaZ0zSKfTQ9JpqUiYcNklAZx4npVXXJMLIGRK1lEcYhLP54+806
6TQSKftqflBM04xHsTEba9nunCqG9Y0w4p4Ptiu63FB0qdhHuFw1f693Eb/lIG2S
rlY244wFupRwQ2IYVkmutFXS4xVajo68wzFIGEYPtcYtZJoIgVYtqUVPoKWGNywv
REve9zDcq0PpV9+pAV0xrK9/iAnP75iQgdFjl029Voi8Ah5Xsm79dnrM/mLgS5H5
6uNTus2iN1sX8rQVo8vWK2M99dfVfDG83ODLerkKWX+KQABgQzNj3QDWWJMY6QSN
bnUgMutzYj0PlJNTxGt4NpUytHqYZVeLgPzXqDatM2m2wZQ+tRElRjDZIA4OkLnc
UCZtgCF4rWj+Yyq87Eskq/Ib+fzEjL70UNYAXlxC76p1EgBlDQWzVT2MUzJhxyzs
6yCxjkTlyrX1tjsVefpqFc5pkZog+IyW3ZWQkeleZBHx7u4ZFk4TT01JNFeK9hea
Scl05QJTv8MgLJ2J0nSUDZ+z8S93GMl06iBuIPg/pF0xfnGjMQS74OQOylgopnjg
CyMpBSQtLLs8/7n38xdRsqB3LXLPtrdmFBbxujUAIV7yCdaEHybte3tJ6zqxLzMQ
SLeomWD+x3XcYwGAe6UGPdgC3sfoUCvoyNi22/SWOLJ1T1mbzHpBB2VyGgyZHdTr
4b6v65xM3E8a0AY0r24Pk+vUY6LIMW+lIqrg3JBuGRKOKBKL3V8oYR/8BpXK6zhb
xcbGST06PXh/CMpixkj7bj8D1MwTIBwU7oN675QQm3xj+lqlOhnnpizWhfwEi17Z
FpUQewuxknuS26mzbetrgmpfFM/yOKnhbn8eATLGqi2MvVjy+jlynRNA/iItj6Ux
TmwwY569nIjRp7IqIjTyiQtnBSEGJObvVJQbMATr68kZwt8PPobRUQ2FAbznXdd6
FmQ7GEhx9+4saTzkH3gUSgg5brkd9cF5MPTxlNwEwYrxRB8A8rWLbqhgO/KwSRd9
JJL3Hc5Px9LIGNhL8s4gTmXO1+49nAnePfsqbZgovaMvi8oCzAE9yeAe06uoYmEj
RFJ39wj1iJ2LPKQrSdPvhI5nOGMdW8RRt3ys9LhddW2f7E06e2pVovtGNKxeGeU2
EexDVtHZr9rzRkrb1rjiltkXZUbyTRKdV6+32dKZ2KCxBED1PtMiwmRHWYpThUnq
0/ac3r52lfbLcZrzU5gr8UbkKw4ag4YWgm/ReNig2BKsKulZ+uCv8YF+B8zLg3ho
X/nmpVnG22InUcPjjX3lMMVTedCAS27qwggjtPNWEgSrghLzYnTj/AkR8NcrdKnG
lR551EV6t9sJvdzJsGz2pfAK8LXtHOIj/ub75i7t20mdcOXMzEOL7p66wxI9x5As
OtejRFUB1+8TfoRzUux7BjKHYzFXyt/l/slMRlGZ+QwFgPcMYWRF7zhCVCSQ3xR9
7IUsj2f5dUU71/csHL98IHkxAdVEn5SR2F3Kd6IRugM0NFiXvQYRvN92QO1mgBz0
Q4rqevE74uKOFt61hU8MUq4DgZCfcagq8Nd/pgMQIQG5fuL9GNnqrWx+vwF6rw6B
42Orws5FA+ihwmJxeQ4qvccXdTjX2rfVcRmwX2x56Nv2RepfMWM1fz3EXg24qC3o
ebACtZM+hNZI7TFa2qoXRw/MM3+BMCI/W0NKwaKnLLQFb8qN6cmzzUW2rwGNTvsm
532/EC7SMnkUiluP7yi3ccU95iig7yNGpwCYfrXJQ84HuLS3yFcTKQGGgcprJEMX
LJw0AXfYkTzqT86s2RXdTyrYUBoeDSgNvOk0Vxmh/s6ptVKe4dw3YcwCRLJp5RL8
jhVGSy8mLVSIG3X2xeEKKlobUjkQZijVdvlX2zidTEngyfZkkAlSJbmUbsuKkvZ+
yDtWGJ8SrwouxDvksIvc/oyeYtJl1c6YfLNHwmJDZOs4QP9O1GcfcqI06sAmwgj7
ZOhS12vXOHxCwF8c5BYUrUA6+QYlKH7HWshBJVp22CB+PZq9DLhXfOC19b5klbwf
D25mVwVAzz2r+YgFuWkI2eTfZlqLddZsYZjNhSKHkCV4fGRltDGGcVym5+TCuQpX
TfpvwCQJOMehdeGDwSdYDx99xSzXNlbt333vaXPhnk1XTYrvHa8DeuNqIh2D8NS+
l9p8k8KoJV3+t7Gogy1SAhHtPdfsSkAnZjRLQgAES3sIvSbjJ59sAEbrqXZZkOlh
ueS0OAWs62i9fhV+C18UNf1kCupKDzF3SXU7KbUBXbF0DgTfvsKmgESXp7WMsS6z
a/33PuhZ2JVjSrY3+UIiHHwJnUVyp+ARCkQAY8/yXWPAVU9Dfo4uU01UuUadR4ml
eYsGvB8uLJ06vUwhFWbq5FJa1i+F+bx1dCYFmE7mas+5C9AmrffmzM9PfCT2rh7B
ERL9u32ZmKwGASQy6XOBxKjeiPgUyD9s51rtHkUv2h5Q6O2PKr+W8JLSv5aqVoNz
QNs49Uz3gZx4SCw6u6rYKfR/e/dYbB+F4pq2CN5LJ8a8Gp8wwbGamnnoFZTA+8ra
O9fYUcd1lm4UKqi0PN7XD6eVCDah8T7KchDjZ9GKUCvjkWaaS59A+xlteDxRLxI7
cZKDr/0e6efMII2PMBNFERvZw6Ywh5G8/BwuVKrv6I461whYowmcKH7LF8Y7OKfV
WvNUZlm/D6a2BkzGHXlMh5OpSRQGE/DEaPWG+gQgR64cNBRLpSi+925Wd+arPj7a
JJZfI7DTBRgWS3kD9JItFfiUlD7/hWJalEAmN0b/rtX9ijKZTI8tY+MQNyPshRSN
VRY0sBb71JUe3uxxHquQba2LO19fQRZsS33qgtn7RapVEEw59xRtVLg9AgK0o8ZS
gRG1l31dmxO8tzghR2aaBtTZ/mqqUs2q6ROQRUyOkj/CqnlBD/Ergt3o52vc2wTk
TzeggrewhqLWLHCDGiU3JZqZSJTPbBmqXfGX14/ZEG+aDnZbcqx3BRacvtn42SwI
Mvk/oivj7IBn/hk7Z+TMOfrA54hfd6JrOjzQ/i6Eih/OJwHWeIEKO/647mqp8/wo
SOFTHhzt4FZo0+vVYiRILN/Fe2CqyfgiQyzL1pN9jKbHR2/AIL88Nn7Qxrixa3NF
11GeddqtG7iffKLnY0f7Q1NOyKmCtJP6lRrY1AJx87VmmkostbE3y93yZcrilBME
/UX7bQxzRvCfXnumWbNc/2ZOCpA97JdF+AlP4uOeoAkj+QgO9YnR4LXTi6gu033p
l5qQLNvPi+iEX80PIENN0NZxjVhoGZOcusc2B6twwWiv9/YaM6KZdocmuxsf1yw2
YUBXwuVcr9jax66zZ3XsNlf5JyQwm4caMIPcxxI/LtJRv5b8nZzdswlGZThNdhw1
w/PEpz/m496fIow29PFkgFvrmLP0kPHUwzTOXlwjLv7RYO5qgAjSgsrG+d1rrGAQ
0s8NpXpUGlvdtwTxGRRtK3mvCGuDf0rlacodmOHFzSqcSzZrpYEQxNxMFhSV6ZGP
vO0zbqq2hyiMazhHXxKvl6t/eqfyP88mOthrg0L3AU9nMRdhqhk4hevDKPnNBqJz
0DTlOG45kHCn1c7jCWsdg0wvTxB1HaoY68Am/PpawpPeDs+yY26IrDn7A8KP1jST
5TIFn3qBN34CllQlsFVSXhZn0DYRdr+x38mVREUIYpM4Z7nhUIjf48E7z93X3wkI
YYWY8avJPLjLWjD0zn75pAYeaIP5SQFWzIwHvOOLKOiSf40cbHHbOYF5CqJMcAsB
YO+rEif86tC9WkNrIvb+Lesez1WmBsTuSzberuQx9kxIjcVdXCG2WQ0WzGfxIpdV
8xQU047Q1XIomZfoeX44kIQnYCHLl8JN3QI3dEJnBipYNaHkops3N/pVIYKoNhPr
yUlxH/hS/9Je7iM7yOOl1hXKLfrYGtDVzPuzXo457ITabMAKuQwrcVIzuKmvNwel
ouYL+gY2ene0B7CZ7j7+gSBce6RfTTblYHW+15ABPDh95fgtsiedOhcte+XcaNTZ
LMSC2KschGJORgHqyu9isCgBOKcnehN70+qf3FAtHxnr1eTullhmXWgcBpuVFlA5
HCk+ROR/wnjzWME9kEMQMCN5s2qIqVJ0p/Brl32hJopaJvKYIrkzF4gFG6bsHiSo
D6f0HBVUPeOUlXDV6d262Bp/GUajjjzLXu/G5Zqr9K2SvfwQdWR76oc6pke6Ztlf
UXsNWSd2fayryP9OrylwrW7hG0BTN7dH3yzxp4yWOWcPQLi//15ahz5R3JSwsckE
NHsIJb8nDB8TNyVvhbMa0zKHZ/3egyxbgwRtg8fNXhIUkQYhfCP9r3B0NRVHUy7f
gSzM5mAPqJONNjD+29RJXLRBDWy6FAqqleS+/21OfT0vNVdGV1eKmqz3Cx45hd4w
5ZJWHp+aXgO8NwkqOdsuEhQ9hUUnvzfZwgwc4E44bol477z9/hzlb7RO8VmVVkvg
irWYcUOqsU0+GPGVzu7vXIpzvaZRJW9KTMKqExGa/v8xVlarZWFG9s68f4FCyVU7
K8nBlFSUWsPt21hal+23DOOXcC3G8ra0jFFThbJyVBLMPNLEvRBEKT0IHKa6dugd
WUg4WCzJhcuAJNn7k9j8N9V0UhhBrgc5dA0Ka8y9IPH0DsU/PfhluqpxkOD/Ftoo
UQlhwdT9xIe+u5qiSjpyYfZe08uDrEgxc6C9y7hl8hUyd5Vr+VhdWKWQi3TLZZp/
EzwX1EnjWYPKxPvEcwH+dmatcC05++Patmx8TasZ2aD+oL1leeEACO6QonNt0A7Z
J/JBqYYi4brUhBKzWVQBPs/N6/33AgRccvN5vahQRlALQSTCZsRe0DJjS6fsRZvF
nku4QH0plsemS8WsW5Zxh7tFOMCKpmGGypQxDXpcTeF1kRWaGVjoNPFEQcl+/bEJ
cmD+7siLjmlt3SOtPS6Cz+cCHfyXjXl0iqRXiSacYrxT79w7ZpGpBBWEmwEaSUbV
tsWfWZTBmkryOCEvFrMElR99zftDdTWXFYX1dZrQvqAOmdRvR6LrwhqVN4i7ENxF
lqRdcp+HCvpVWqEHPdGpmGMswyajM34rErbUIlGJvJRCt+GfmilNbMFDHeVMqY8q
sRh9ECn2cFMPT9HjsQxdRcYYjW4R0GuRCzepG3NXmiHEFM+7mYg2j8De+ykAUTXN
p//dUq+Om4jq7QAjpwfa6EVmlGN5FuXgn8uso3O/kt7pi/fAgi14cFoJX49FPIJV
UebjlIX9k3yuqrPqJUNqCsydTEawQAw/vaNUu70osPxknQK1prkUmTULdbZzsZ32
HjpEjot5bTKHpNSbE+AOYtKARqiWbvHpSYAoGXc2r5N/qJVK0SdsqULxmHnI3SXs
uzxIvbdFZJEMyzVayxnKLPLMaeMWdseACei56Kj/++ywjBbGz7B+5UBm2z3cvPp3
tqo04OmX3Nx/k86lGNRGI+iKcYCxbeILTPGtrTVdjQlZUYe/oEY71GGqOrr9d37L
g0EkVfy/jEwQPJxG/IDn71vN9ivPuJ7vSeqXPcjcUeTElyw2pUok+0P+GagWmYZ/
bfWNhQVu5S5xCNRE+AwYWJlfKTeGdjPWbDXHfgRStXqcmcyw2BqLVxJ5XGM79baO
TQ+Bq/Ah1Rh4zW1N+hQQ9fzmxSFFqXAXkaPVmfqgKv2r+MG3qWO9wtx4qXZxJ1GG
eBU7CPqsuj+qZTqYYmbiGg1vmdYVXKozbIjfFanfGrPBascaovpX89iSND1Dv7wS
90mEEvLwVSe4cH9YT1bEiyjdIuz+v98RsxSsttKEq+EKabu/2CdQb0ia/qWbFkoW
H1vyvskWp1rWx9B40wbEHP4ejtKI1A7sugokVTPrOX4ixvthceCboy2aeaJFMtoT
6MorE1R+au2xpOw2H3Vym4Z/HVxIlOoTEnpZF3le8BnAi9b/o09nvbaKe1p3NGO8
JNgFg20xFsatcNnbT4zqCR8lpBmzhtF09Muy3FvhG726L8ojC+6PxlrEwwddB+QR
0oxowOzA5xCBD3ane0To+8WpLXSw46tvy3qFMT/zxEJyxdFRu2oLPMa/fS/9QOQX
Eb63i3DNcjl34jDADRHw+nup3PW3LMco/P2fXmJ6ntJ4eC6KA3zxVUjSJgtU+TeN
UFdtVxXcr2wZpHj8EYPMIjV3L5NSt0azG90UFRE1na+mWdWaAI4/9H3rlp+QUIyn
KdbSujrNKtzO/VeW4zsBTr4DAm4p8AN4GEc2FWVkudQJx+1ZhiO1mDJmxacVrVQ8
dAhYBVVBCox46MqXGKAE7X3KsigTvAP19Qu9uO9DfSA+XqsWH/NTXaop1BpmzdV4
cnaQa3oYt5ummxpC11xGdIqZKaLiQsdMzxRpjSnEwh7WkErufKViZSMVSC+RdnE+
Hh3ITpP53LOOoxxqwrNs0AY6jQiO14dzz4rrGvZWx6gMWeuWpkqb7eekTNGSb/Cn
+JwqP+ELn/AxzvjWIeSXZJmhqb61S+IOXZDOmHb1oaXj9KmkXtLpq488pkWlUtkf
X52SXYMhxQ7kxXXa5ZZzjzxCba8xgD2CJi/bxb4QMaN980mKY3t0i3Wcc9pc+jkf
PuZPqoYN0bDIZaKUF+/gzAxKj9Y2SeEqvth+ugVmMeJn8rNWlKuiY+q0LN3mDAKj
kfq1rF0T96kom3Vhg5yQYKRdKwIJKT1fP/UMvzMQu4KEgy4thlscdDNaY6EtA3l/
7449zLPgPAwTBWvhRFwy2Cq4Vv92i3fSoD7uL3lg9FHK5izHqhYNdO6SU3baL8cW
yo4nd+XITstmOeIGEa4CPwif/glBZcMPt41H/+9uxRelA5ysEXEhWq39OEZIMJJ4
Pw1bIrHAhl4b+OaXpQHDlOiV4utrjw4NhThqx7UEY/sSXSwqr+kgCjTbgV+tMsfO
Jm63JhrNV9HBnQS3o2sqR1CYovNXdJnSdj5aMO07Z+UIFw7wmELMP70N90h7/dNx
ya0ZBxv1DoA0raQsEqh8DP4hmOfPrWK1BBZPtD9IU+c1h8yIlldisTdhceq1yDlg
RnKXhvS3Qk7VnHloNZOBFABQtPrcRELiqLFCFVLQdJ34dLtIQkEkqjlIIyxr6NWu
W+nGQFoBrPqLfZ+hO0eehZt0givYW88c/BXRayaY+5gxjw1Mk3G1uVYTM8ssggn/
N4BdIprNnkPVK1mQxW+hCSsEi4Ypz1podPO1Cll4MOBOS4sLUoOxMHIn5jMRgFnl
FHI/ZcTCOXTqIyQBxyDfrqsraAsnVxHXadtkgMEug3q5bZTts0UE8FTcM663mNGl
91z9gYtD+5khfjWzERjhMb+Et2L0gcG1bsdlEg5M810ZGbh7qvtkKBOAKDbLRTno
SBZ+w2yQ7IrJ8uLF0t3yhr/sLGPDsXyhZsG4xfgDATQnPA3M+EzYYnHDSYAHv10r
yrzPJJBCPKAYK2uQklI7ptKCAxg84S6Q9ynX1NzK6u8YNY7asv5HsibzwPi2ppvP
I4rYWwcwo9Zj/Ghy/wj2vHNpsC1tGoXi6wi7ybP2Wf6VB6roRqeH2QCutdtneuRD
ATP1tTf/e9rwCBOn1Tpb/41wM5RdRUkFm4gDiByUDtZ/IuH+cxMWZn+QeNlx41Cs
IvTUYQfC9mXV2FFmI51di6MljTq9bdR4XD3Aiso6+kCToSRk+exk1D3X2yajQ04P
KX9g1pf3Bwrwfa57uanbsjcnsY0YdDQaHXtw93kFJdZEfTlB+Ie9vbJJDmoISXQI
0WQtsoBqq70Rx3d3viHtqG3QA38TbjoMjX9nILMI8tRgiDPXNeHvzY9UXTgkOjzk
q/QaV9NbH+PL6OuE9vIy1v1KzKhglN08vape908z4YIZWNXTEtsQU5D2gUxg9WRS
1OEsTc3FZqDePzOyxm0nWxNU8VvCpP4TOcTu+b9o6CTPViqaNJrRaUNynl21qpCD
z9IZvQOfAEdXFgrukI9ABe07FcRAKHl7inLtl1ZCgW8uzHO3mESQjIBuWqaeuitB
ss/Q1eIzBk/f+ZvuSdnUe+WNro7xq6UahuYXURxUVK2If2F1vlItQ7oz1naGnlp2
LNemzsR6Y5ATKZ8Z7dv6VK9Xz03L3OeKqFrdEDxXuw4wHsci2aASBbU9mDzZ6Tab
c5Hx0vUolgrJZ/7SrD1HyhhCj//mOiP9cRuBAS7BJVvaBB8cbEDeixrPqLle5TkI
dzPShEh3OdUQOMmPQPmdirdFnqwlI7iaO9B7ii5MDvr9iiNanvYmbNi8f/ywD3Si
HJjKp0RIflB4wggrFDwZ8iPuJ5RSZAb6pe+vuStiOGXweNe39xNmW0BO7krC3L77
A68ymvBUGPm+SZcqVQk37c3dq9Dk/aXLduwg7ucBlGzS+b7tpo7e4VPrcT7eF19r
uWX0HnwqG0eCxwTw3AoKCxhbZw0pOxMyPHZT2qGCPx9m4OqDC+P/HIjk/naMoolz
Nk4JofP9mW1ByF77I2ZF539vBFbZ918ajUYmjs9gMAD+aqRiidzDD824AVKT+Gtr
tY60FTfB8MF7eStpORDxsOWPB9+Tka/jR+0MEHQ8UgNsnf/ONDpxqEp4He+0lrKH
Tw8GmTHvltmMFGS4KwQHHOQeydxkI3Sx2iLRBPu0Q5mZd6Psrv5JqVZtUPA/vlWr
EGKXDkRLV2ikkjbNOu/xY52CsFvFO0m6aqegSRUNjHc10ToWe8kuTYG61nnkwigA
vAXgABv83zeDvPsV8W3DKNSmdRtJ/2wE3Fin4nES2QGABVpc64jlgYOw8srGre9N
lEylPzYA4vn1d+XPt6fvehqV/01gtLhb9YA1V7D5mmXjI/cRMBibXV6uDL9QoLad
7YpZ8RF7lrcuETe5Jad+eRnxr5vNBEc3MDmt0x96zJOlt6VBZdnJFaC21bV6SbCk
2/5KfWbZWz8d0T7acS6OQoOGr25gOdGowDzK/w+eKXOlzb6VNwe94wmQZJJVjw36
iYHDQbtB1A1XLFBI4JOILH+U8ZZvblex2LJUCYDfy+Hmsl4LerpKLWl6kRf3vS2L
yBBjhJS4v+CssF/G6+IUCl1fsEp6vGTI/qUuMf2zyyoohT6YIli+D5l4VEPSoHpB
UJeTJU08lYIJcJYcceBJf3cCYEwhXH/A9ua4zzvmIvk3VESF3hTx/0vtiUPMudkI
kCqkRUKHMmaYAhUPXuNjKyLxY68Gm5GnhNULsh1taSUZ8QBB+gvA90APxTGmZQV7
Y1XbJ9gWfn7c5eCmWLjuKZ9Wr31gV8Ar9nlUvro+Hl2po8NQvaH5tVjaFXDH98ek
8ROA6ITx0Y53Ph6FBEcNxAoL2dXytZhef9gjjI1+jubopORtx8minmEVZsvWCbOB
Ulp67iP0Il8cYCjLx0QrrzGkLerzaIEQxEvYUO7E0Z/3trpOIVuu+yPKpFEZSE/w
YPYi2gOJmvjxAlvSLmCfrb7xFmYUqIS1s+4iRyhe2fN3p78q4PSyYD2O4hILSsrb
96GX+sjBkilTp1DYGnYqObSWL2Sg5d9UrJ2aJztawBdOY7Mt3ppn+tCWpsD7YxxU
CHHg/DMj/xKAM/utidbIk52IqOb7Am3trOQvfXrPb4ehurCAZoLMB7yVt//r6eht
EyVNrUd4cq7KM1DCdZ0m7LnMrs2eESZHw154WhPnPhV3RoMl5jBozLDBNUBqpJKf
ulAjIbqUIrprYabdxvTJlIo83e8CTGhyQfV1ZczLg0nBkJWUuNqZKnBX0w/Gx8L3
mFcLyjmEvCJp8ieGrKdJ9qmZZwO1gejCGIT/NiUs5hs=
`protect END_PROTECTED
