`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RdzGv40RLUN6eCNRjZShRl4pNsCIgQ0HRWXZyHepU3m5Rz+a6QKx8tDbR0/YeRZd
OOvNk6z4rqMarWd3uaIDkMvYlkwn4YI58XRVVN1iZfLujeSck4AGRRav1y+XANB7
VHesC9eCCm3/VtKIGUvfywQm8k5wxA6cVngoVzrsdVcknXqsn44NwpBZ40qzPaJz
adHsUmTqpj0WCKAKuflq/85EyZwwLnLSQkJXW3AoA8P5UCA4U+FVZPiXS/ADlRCO
lrygLmykw9WDoupW3z7K4RgZRECHx65g//BHHv0lgAKg1Rg2CRZg0ghuK0JMqxzh
mG2UpzsK9/S0ZJb8Webva/HjnE+y62sy+t3wk6nn/BT+6koVF4PrnCbrlLsn5Avp
sUpsBQ8OddDhXHKluL5v9Hnz8QZ0iJL+W1fOqsiSWv7hiBzjlYYaLgns5PxPwT73
YybDmfw5mqrBlJlVJbwPhVpytyLFzCDIR1RQqFZzrCksKJAGzscY+c8voYUj6Z0A
bcTm3gutxZ95uDYp1uUNne7Y+dXE+NvdoeAXnyWKZW4cXZH462kIbER0TOh3gOx+
dCeU4rU8q+9NmAdvx6hxRjDmkRVX4Ly3o8583V3v99Y/C4LlHVqagN0UDlmzRB2O
cIlRU72F17IFKT40pXtNefhXAJAAdBbMD1xlwT+HgxXa0bHP68hbJQ/Quy3SvB+G
WUWezlCdXp/Yjx4wjLgjW1eY8HUGSVz/cGFaqJd2bBIF2vgjOMf24GxjaAk6I78l
HTVTPYd2zgejBtuRU53PfwFF0Ybxu66ROjEsJiuilE0+S6vLhkPAcYyP4uxCIj7s
KoCI/RkLS/NQ7YIeMTAhiYpzZ2s2Gehie+A8BP97N6+7Q80hUxiNuivZtocO7bCB
9z8yQVBFOvh0dCcn5ztEo014yQ2KGroSxxjzjQXucuRMKY7PnzKZWIcYqiCq2gZ1
yZcb90BszcTZBS3HbuD8SpL+HGH5dWKur3kR3oqdTbCWbaeqRStrTWE5fOnOAiLk
r4Xdz7WVls1ruXp3zRZexg==
`protect END_PROTECTED
