`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PiHgYSu7Dfp+KOKfVY5F4G1pvgBnN7e8b/fFc68XvPvTKxWjPBlhlz4lV10uL7ue
toNHSjGHnznX0qzGjP6qgCH5c4yQOlEVyH8THzhAVdG+/12bVvgDyeMpRQO2bDYu
5yy7TuOgVS5K7jSNB3PC30VBbOWnTXQAHP0SzxYvzMH50pTMgg9CJdTiAfRNqzj2
odlTcNhd/szItRHzbJGl6xTl1REun/GUHzPs1VB9HINGtPUK13pY/BlnVr2qK8xx
zBseSyWMYVWmhAJNBkP7LwSdQLgSQChapJw8cnbsGnWYAAPMdtOEzgW2NFK75NtS
bAFwxLzA+EZAkpL4K/2R5XYPaLr3dS9Of8ihXO15A22f1ionMvCBiRrlqfQMSCED
dbLWo6vWVuGuB4uyj7pAMG8Lb9R51AcQm+bd6vX9LyaHlKzwy3a0ICOMszwMsaKl
uFzgv+NQEU/JWsHwfhaxcKnCgOzinXIyAxS84XCuNikIXuhswqSqCgiW9uKPpU4f
9DpSMyeHsX4UhC+h0eNNPnPU9mo8IofSWxHBzqnM3L+tNnL6K7A9BetLPa+SFqoF
R44z5CmArl9r1lkMkQwgVESlpQltu0ePnFq9cjOR5YZbzjJFps3qmmOnpkwN0H81
Ob8yVEY5jsx1s3ww/fz7kW7usMZE5hswwZzRLqFIglIZPS184oH4FzyAfLXVq9PX
PSF1lWbx7LKm22eqNwQ2hp2TuQ2yR0dBEjp5/br8QmrlztdeNvq9wbh3H4ku12sT
1L3hIbWZHeaZ/PXJJcBTqGE8HH2D44dR1iTV/71bGW45yVxWmyHF9af7ae/7Mqr7
vrqFzEZ+bDobGUHWwYVj2wlsshE55Yp0jP0xxD/NEKWMZ13g+yJwCRCIEIMWGHvq
Mqqzc0hCjfkm4cdUgt7F8gKDaKqegBFafDo62tSS1J9HGomYlxyMeyL4/8fC70Lg
D8qQ55MgnxhMsEvhgAyoUuD8jKClxzKNvJUmP8WcRZ8pRKCHNi6yVKYyChARKDAy
MGKLKgbTOFORYo84kzUyvSB28I+K2bRVW0Pgiz+GQmVEi9Fq/gLdQ/Vv8F+pGXJ2
JAS9L7v/i/F/kCMI4F51yxT2u3i8YZTSid1hbpMW4D+HOqt3dv3YVSiton7YQTCX
BvvbeII0nB96YHTtJpOsD+zNojhtSVrkhvwkPiNSGE10krzh6ID4sB+8U8EZTEhq
R4Rvinl8vNBHCL2UU4bdT3/F9/VnaZdjFefF7zhEYIIs46uFRHU7tHd4p92p4gGw
uS7S52Sqg1qRQqb/YPsOUf2njYvo02wG8lIo0IFrQCs3KA/ZY29oKCXYTI/wEvXb
lIsOgzSK7tmEiZgutxCQ8A6FSGBrueF/ZOckd8m+bQ7v8P388J7zpLXdjpSnHO8G
VHTrWmdutTK/T68ixzhhzgqv7v2Qt3EeKJnBXdiBOtb+MjoCxlQAWpV+H67DpcC8
/LUhnVt1ITSJQ2qzzmxbewFx4nR+3TLSd71ykokZ0dsbS4aAMqseldcg7AkF5haf
cyh7yCCoW5jDELL8gtAUuuLFGKYD5wg/OQBrDMW5T1iL+WOrzOJyfc7ZyhxZ+jHa
G7/RFxrbruscRLaPrNFWhEzUroBJrRfKclqa/jo8LgUlzuFZPp19ETOyeK0hcOjK
KAV8A3TLxp6sVhr9uzxVZ3L4R2KlNrQBRE7h5/iasNVy4InJKDKTl0day8W+ADea
9TRPrsAobbacE8OAt7N1jA==
`protect END_PROTECTED
