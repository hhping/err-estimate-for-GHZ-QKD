`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFo/E2uU3gF5QaI34Y/tyrtWOz6Wuy8xLQ0Df//Otqwz7yOqYgeEKFpbUtK2dzI/
lj4HR/W8M+RMKfXgZ6HCWJhEApGBrrC1drsZKBBzNpOPfXVHwoRi8JC+5mkT+YWh
rIFC2aHV/y7hDeCtFIV27Rj8NDaUAJtWgenkRclSovmErkkV+e6x2tCXZJ5frbpp
KSKsZHa1SxFFzkb2JHmrd+KONDaVYJ39L8ak10ei+M/Ed51smJYUkqWjGznFcJ65
+mFMoSc30kut2lmXT0HVQWb8B7aWa5FGRZbLNhWbwz0h5g7eJqJfzhl0E5f1mMu6
ao+3Amz1HItFuX704mbag7Ezp5XnV36CNKTGhWQndXT8d5lqR/gZRsiCVxesfz5B
9EDVir7Vh1Vj/nsnjCp9YuQ/vjjF7uIxquqf+RltnvVx3/pdq4e1ROz6uA2v8kdy
dGcFMZJcq2Pt4FzhWHPyuWxc3mmNf52BpsdomO7y89Jx9ylCN1TdeMGHBLBU+bBC
8iuoYTcvkqy4EIHVzkFCw6fg406KsNfEvUvIVdK2V2tyIrvu0u9rAYHeqoJuu6QS
0Rdt52XGLLXhGMzaMX7vY1i0iQymfmlld4NwNXxnL49NHyYNEHRaRTa2ZsT+uPFz
`protect END_PROTECTED
