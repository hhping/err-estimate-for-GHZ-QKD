`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9D+vyME4hLPWtdqpWpqk1tuCBFD7ygnyUwqPtnqB+9Q+wlVOk2ayomBxGqVTxlv/
1Vq0vqjDfWKd6//OQadxpFEJM4i0nM1mHg16lmIHWILxInlwIYcNPt7QgtrzKiuw
hZvNhBFvNQif94ohpzS5FRheSxywtsvKeIU0nEXJC2V2RLIhtB6XA0ZBwaZNvH+y
StCJXcoaN1mJyEHQCifqDWcGApHwGmkri+V0H9WpLUstKGC844qPNxzWBONnZlJV
lpVe6konVSGiLlU0nwrF3ZvzADbLOLhPNYW3YdKTGH2vZSRsucf39HvOgYxRcYPU
BeKrpnlEeO05fLcblI9z+QSqFlubptjD+Vj+mrUMiSORs5q5myrP3yCijNPh/UZB
5jNroKeT9YRJH2emLdLef3tAVYIlI1O/ytoR62qRe99L8LPa5FDTWQg3r5a9k3I8
NlntnavJQ010c4hHdOCUBa8nRXrb5AP1Ji2wpRvNT8jxEPIZJmh3V1wGzDa2uk0u
v2imF3LdTSRTFmjQXcliD+vayrNP+zyZvacQCyZtJCsORWQEDKw6VtbaqPIS4NPE
/yA8fLQK5DnONXQnHdpE4WRTN8tJhtHjbHjn1XyuQIna7mWHyK3jX+rKBldvOrEp
ulODTa/BjMv1NWImHyn5ae3m/vqPe1LtPNs1ZerkRINW2cUXUNAoIEbr5j2Hezcj
jnlWOvgcGMnE6CHpexSC7g==
`protect END_PROTECTED
