`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72g0NZXEQMw0+fqTotb159uGEjG+x7/UU8e9tNLbOGFBK5FosqWUXX967fB/LWzo
e0KZHlZ/v3YwJIEDEWL/0H+2R7H5i4ve5pu3oGb7m6XQ43lPrjL2smvbd31p9B1Z
RzFrZQZp2U8FDB52nBzl6UifVigna/cyWoj636lFLXGtSRMf+5qU3hO+vQgDK0x2
M6DCMfpYBuMxqBazz8iRx2TdLY7g96cF0FIcdeO8/SnTs3mUeBH6pax7CUdFAq1k
UiYcI7sGQKcqqW666DLkOxqHOaX1wOzGqTVB7kLMtjLI5FGhpV02HgQkL4+qRa5h
vN9qmW17gpQ31adf7ufUcjuwW+iPut+Lscihg3xV5aULSZMoqF7OjcxI03iZ0xWY
ThGCnYxGVJeeYQm+W/xXu26gce7UMTh8vrd1eov6sm79aemEV+O4wC+DS96tD+8K
zHpXoV2uE5tpEFWhoAXObIRRx/eZwLHU245x0mWtQC2wipdPeSO5yDfVR8wbe+oo
upz/RSgu28hEAKfuQbQhdX2+Mf5EKHhSp7VIke73P9pnvGMp9ye+tOF7H9tHtHdD
NGdjyRN/m6meODwzPdJUPx/tR96pyMPWqp5gemgPrcRtzP++CbZTzkSCLxIFtL3j
xJBOIJ9yOPqM3riRF96I7yjZsbZIWIZAQYuBKLYLCmTt/vO1dpmVIDZNbCPVpDu2
evfeoZmhqQtBUsxPBzt5oUKZYBlXaVnd98RocpVrqsBcimaULwEcrIIxx6E66+LL
miEnIbBrxXiJywNKtueOGor+lK5bM8SA95EnLAnTFXX4+A3Htal2XK2/Eb4+mmxj
NqS+vmLXKdOu1h8IvOZKzcWA8IqIL7ARRtrGm792OrWYsPEyqq5tksVdZ0QCuyMt
vIKwF6GLzR/e/a9AABdKkA3fdQu8dMhqLkC/P5CaN20p8kpeTL+GDgYRNDX26nU0
UnF+/VhQq0AqvbJ6Xa/9j4203mwcOwDBlwNIBSEV2NKnk5QMkivpcTVYIeDdC7MG
saeGns1DksMSzL2FbprdKpwO/w/E3JBGcnrQHzIfbr+zYSvvadUhnIzXxO5j2g1u
enDnUUNE1QPgI022eH/tDpnxneCUsu5x7JXtx4RGgUj+6PCudWBWq9hvFo/ukFU9
I6620HzsUOlcjNOvlI21CoTcZLySefvSGV8N2ySrOCNfpSgvMGI5HBnHywU5LMfV
3wdIswXjAXiauuZVukEI2SBT2z3/9ebt+wfo9zdctcIBxqh+kwhsHT5Fx7GFUnKb
ok0PRG4G9+wrfmHPt12DFudo0ue4DCmBzHcXNNOHk4gxqi1V6EopK1MFXKq25Mng
Bfw47qc61DvB94nlQJnQdruVc4Z8wK+OkaliD4Uz8/cZXEjZ0p8RihVwj/rmea0o
RCumReMYzLLoNA26w9TbpquVRKc+cQqG/mvLzx8HX5E3swfcZjuAnEpaq8vkb/+C
dPaDyzVgJqkJAcAvcgnh/q1/cF3WDaItEjvbxk428BsZHHGK5CFJ7ZJu7avU5D8S
iljTexJWao6CxmmQLvJ3x0YLMCIyZRKE22ZFMJ0GsALt6ltfEmXzLUVyri8YhfTf
8C4PflTAkfNeDgK2EfnfROR9PR11ibPo1gNxKFaImEGYdXzLoMPtTlzFqDoZl724
j3hsekqsdfmMEEq1pYsRelqRTexQ0Jx03oGi8G6YqKnxklbJ8zyht2c3+5Gio4Gn
JLVhcbyOK4jkcABz2i5RwmPN4Cg74YMLQ2EG8vGaGsx/fNXzCi7gzGGRQtPNu8Eb
A60Nb1GGdMZ6QFIAkU1BIGdFSeSeMJQ6Gnc36rmJ1MLi7rsWuNVvK7C9TEYNWx8S
PYK1DgRy/M8z4wUJmVf03BtcvxCh+yebqj5uPXK7Df8gErRkGd29Uy6+RGltWm3x
UsL5+qqLLAm6JsvnuwVhmsPX4tVcwzYbE6VMJ7njj7yQOgkygaslYptMCdRswvyS
lub2oGX1OH8t/76sQsQz0LHellwJ1AgOuEnH5Zjb+nPTAU7IsZ4xRs9SKqeCgOtp
IBuVWRQ1qaEyww2FR4a+vahd9uyB4cSg01kw64Mew9ESKCV0TTnQoQbQYrT+06yt
EnCvATZlIt0/NQBoacZZtY4bi/6LgQSG6eZ7qJ80++SymQ3smePOfe+Q5qFEPGmV
pIAQ7NKarU7pkoBbozsQTotKyzP4MiB5wOVgyWbfGQ1LcgGuUbEmEcL1zB6Z0LDt
+YPCvCx38lgpIAsXBFJaT+ZmUqhqAh4HX28tLKduckpmRtBZeXCePQ3k/gwaiVuT
9P8SxyV2P29LWgjGE6gx1eKaV1pSlnledV4eQazeWqALdrZUy16WmkCt40sm2Jni
hlQtwywoFI9UaNbFCfjZnihUekdWy7lWqmKM3TMUjKPyI28p6fXP/5BjiuaVhd8A
XCoEUKV/EzmpJqWqi+dn+aI9Q2o7gWNTi/M++CsmzBrxsnmZSjv+vGTHrGCBgoRK
2jNEmi629ar/vOKmx1Xk/FzrxFfTRQy0v2pG6ay+S2UGF7xH0Z1Ri8YfFGOpfE6U
6L5zTt+glTBOMOUIiw7PqJaw0wKYLaZll4P+71NiuZ2+mTeK2OdPGRQ0KkNipEov
TpGw1T98QPYjZCct8/lL0FTW9OoS/grsN74qoz3H/c0L0fpsUgRVoxkrUEVTAf9L
C8bYIfTSFSLDc0cnMPUXZA==
`protect END_PROTECTED
