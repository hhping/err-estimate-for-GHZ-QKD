`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1a4X5/1Kr8H0vZ51vEkHhli7rGb7r7pw452hRAkvZeurnAig+XzDZ+qKz4fps6F6
SG24czfMnNSRWkiCPF4NJA+44j/XWkchjJrryJtRojA2F3tNReXO4Su8oAwRcGrp
PBIalYf8aVoLKW8qJonPEPdyJNZJtGMtkTS7Nep/qvoiIrTQBZhvBVrCJqP6r/97
m6lUhYVDJ/qhNYKIb4UEj6gV8VfyL1t1RgDjBZIZU3WdqtteUlGQLKv68UOGbEgC
pCMKnXkyshtLSEFQtLGhwRLuVBacYC2z7bnwHxfgr17QH1eGjKeE28Zsl5YgUB5A
NlZmioLFSrhDJglJhZs/cXkJfMWUJQPKk6ewdlic84JlCEXl47dHdGeCiihQTjRZ
taiuEgEnLJDLUL2VKQ2/EfR15GA69pEJNAa5T+rjdghXwf/pI2tNZrgkKzHt33+T
/3bF7oCmLhYxl9/aP6+Vp88rSf3gFSEWAGm+36eWGaXgkQmQkRDyxx4HbR9aUEKy
PReNVzef2xOV4CX2z7mwGlth0xMFzbC1Ae4KCWxtwOPsxtzmO1thpdb2s2Wm9sdJ
MJBiu8IUE9f5f7RYzDvyOqJFMQw2FvBvBFcdNvusZJUcpeL4Eq718GKO2/h/DQMg
bfNIYxq0naDg/fXh+e8GTHknr4MMvF03I/OwBbgoV6yYvUGVvNtVhji8WattU2It
7REbh0rlO8zfhR1t/jW9oJiEo/8hbubxnkYF181jKuZpwNQQ3NAM25qIiiKus9nJ
zEsBqkj6uMnrfotVjfy8AD6XNk3bzxrL5qtQq/OwhqQQ1pt8WRfkGhzS6RkWqxIh
vli0m/sbBrctQ7GbIHTwJx1qs+IaAcmke2UHEzTa1Zxn8S63yazlB8dMdxWnAXji
RdJARUZHfnzerU8wSgMmvX3H5XtH04KEvtJN0eLNeorj+uxDE9qw8Kxc+4Hl0bEP
OleMBlLQNE9ApeOfecylcuLDBJ7/HW3yiiJMfeW9GxNS1qY00PL5frEkKMJlALD3
cYnZcympGKK0iNRwFnVqW3k+1nSr5kpze+NsyTM1gEAAWVWrpvNuxcA85ZlGCN/O
dBzF9KqLtLRFE7dYqzTfBBhQC6xWZ7ifFrDZq58GJi3vMbsqgTzXjTxDunLmkPGD
gqAb0/sxCxX9fleJlXdICtC7OLkGqxpDi3atKBR+APSUrNnLAd/BBp2pb5FzzU2h
oyk4apIjQGMBbep4KaI3eLJdedqePMtQ5HhS5jdYHW9HkkHT8b4Os72b+xsvf+tO
6/rR5D1fQm1PavBpAKL/TwmHIGSGF42UEOcuhDPHGfHG550P6OJH4D6hF2X1UnK0
T9hlaqysf7cvMfCCNbwmQ06ixbGNispteZuPs1dTAONhbV/GmW12weJHGpgZraG1
JFQ4XETzUxBybMoKeVbSH0z8DdGWVaj4kl+HxWCEjaP8O2kjTQJlPqByqOpmmQV+
VOdZk1G+pPYufXGU6iRKnAhSU8b6BFhNTsgvYjLzX96d/mVzHj69CzoIwBWcRPsE
P/LlRBEEJ9khodmEtHTIjZ4w4UL/elL+stlse8ij4Op9QKljtM13+NEUgQ5sqYt/
H4Ii1dhA8EvLsyDsl/X6j7hHNTEEUbaaDwOF5SvoNweB1xCTdI0mODQ4hRTdmlJJ
Vob73bxpf42dn/zMKFa+KE7dx02cr56VrqzZJVDe30RnkAaovKiFjfbUKH1x5uZt
HXxLjLClKGCeuFy3t9JMplxDq96LPYEm6/dYyO5T6XwvSMWf5KGUPQMDgCFAq0qO
El/yjcgZGPwJk+fHjm9PB5jYzU/eSWUNwxOo7dYs47dXg6uQwUhBUqrRa0yb7hEP
larpHyR2h3IwHeAZ1adGg9NTwWJXUh3+o0oUSGe7+9VD5VoC3pjcqGOaNkrDcT9d
K3no/A5APZK2AvfOwAHCj/cXbabuLDKbmIabQMYGltn4EYvcQMm+39Tgenq1pS+W
bCOVtDl8kxnWPlohBhB8t1xFY5tA8f9Ubo1pVibLhc2kABBWfRWCRIoyGGZo1i04
iv+yeZzLT36h21W9QMx7WUUaCPjXRVXIi/8/CYEkzkKnf0/4e/78G5iEj9cFLRSn
h2iEKQ57s6pdT5j0LI0MDTnryWuwzp1KbEN74++6VcYx8b/Gcx9Z3FjDEJyPfcTB
ehlmggV06WjQKdkJ3iFdbPW7PB2cT9Pk70Tu7bAd5mnxC0l3dKofhIiMBaRSHwWf
E8Gt+C9K2h5LbyD4o37eqyaf0GauzjElv73AfE03q7HnpMZjqaEExPsqRbvWx5Dr
2nuv7zAa+xr5vz2zT8bTy9ydfnhnD1R+GLUa7LEwC9oWVkLjhAvG+kCp6xrurIiG
085IxZxkOvusrd9o6l+2OUALT3cGj//krumyklqixeiQzbgl+BmsuTJEtea07Zvn
8JDdbDYLVs3SNw2Gl13athWjy2AjEd4Ph56fflNJcToQ/5PHWfWfBs5fmcdZnIIo
3HVuIwx3rYtARbY7HfqR78wEoEWzQgnoKpkILUoVVl7UIuicn3esfyfpXElTglbf
RRizps15J6PDkra6Gp+NOCnTTaFru3dkjhCTrKsegWN5VrxMD6UIyXGFyfr+dOG+
GAyNPznzaotxlf6gMt9ayc1hBo7dXhmTzc6F7vNJOu0dDKddaFi4tl7SW3ga0frh
A+hkI5TlV6b1hpSWP2/W9qi1dOmR6LtTjOI5LyA06gFHfgtYKfp9YFnh2fFPxg3Y
oDANQjjE50VjJ6ndwxv+iTn8jBKGp6Sr3cWHz6xPdTQrAhuwVDPuSiKrKpqDkWBa
dOfOvKoRwVsBjdqY9nkv4VmXBKEI2CWZFSqDSPoSKiqxq5uIGnRm0QNqVl0YVkKX
9mOoUmrb3I9pZ47tQqyxnpSXpGdM5LuNbHe5Izw8DNtHSu7nnapQGBgvbW57O8Hp
FdBeInjWZOqaS3lZnXsAbONYA3MI6K8oq+tSCo+DYGWpRThkncJsfI06pvkAin+v
IbkJvnpjPMvXMwSgB+ae73E7jpMNysYo1zOQG3anZS5pbPYlml91x3MbU1D/rJPJ
Cl7Y0dsChRn85kMvu7qYoNauNebWBwW3/iKGBuiRLvfznV9ta4xzKUiDTuRi+0Yw
3SkXQrAmnRT/kkMdDVDPzslFztLTkKnVOhsUQCe4XXuZTuA7AoDSaq5n9EaDu5LG
41fUudlj7F3aqzVr4ZMXW0/WCooNChI09uz8/GXeyfKoPiKCNKICIi3L53PEyt4g
PxC1YZkZQWemzKp3v2lRcG7i6851o3eloYN32cSDKCP5Xs4pqq36DTzD6XCgxQbE
MYCju+jy0W/5kvsdYvuKt/qZCVggD5qSfAK8WQb2Gx4qdj8DjgLDlrP5fwj8PHvh
vjyuQzAidad3CklqbSQk7MT6Hud/XqztomGETxi/DpejORR6jpHUxY4+xCteBBon
41BOZy20UnGFeIZysahzVNg5m7GDrLSAoDOH/z0aYt5KBvQAMQC7mXSven6lM6fq
xXiipoJUiUMtv83c/UqvomEI+rmM2jVljijyT0V5qR9/P8dqIhecH+DqqyqMM8j5
vH1c+ZvVnvIqo02s2MxThZM4U1HukJHchhl6H5QBVxb+fVTIoFsC/2xwKc1d4osy
q1CorgY1tMkwCWrlDEkjamkUuu100Uo6clX4LltyJk9/kU4+NCdwhD1jWseYt3xg
NHcpt4i8TZSevuMNQoBFv2reJyuuZlu9/op6QD1HDErs17q+qzJUsoqx3PYHcFzj
TY8Qvti9oq2uBTE0lF91UY3BZ9zGy0dRTMSKQhqIhpFuVrC+lDICLt4WQrJNRhuM
s27f9X8WGdQMCBr3pe5CQrgpAMfSxMbPAd25NOJ/ZOp8IxpDoFLGY9JWPC5ZyGyH
m7awUe+GH1vw4CTh5SyAS4x9wUcNZqmG4Ktz+xV72eHq6IxEWhA6iazfu8QvkwOT
Rv+jSaXHsLhHASe6x70dQdnf0QuI7euVvsz+aUDc/Cpx3Gh0gPRJ8GoUOSCvczc1
7c/8y09wFoq3xtZNlTMhqQio0O/VvTvz8KmfOIMAF9KiDQd7d9z2V+ApVk0rWLbi
ok//uTTR3FsDa80gUdPUALeP93LDX8drWCHRjQ2Q1YoK/wqZ+NIaGVhN2NGcR8RQ
Ha3VnRzdwKxx+W7rX+xdthuo71XSn/nN5WpelQ3gRcOi+ZsrspvG9ZQYWy/V2/Mp
Se3oZFHOUk752qPssQEKAcRwSjAZiiI1DNWkO7MdE/W/fVtPsFX/b/eyGUhhWdAP
lbAtlXJ5h9E0LXsSL7TZv1eTa3qdU0nv2BhneSbPMbqo0f3O1zPn5DCI1bGuWwjd
fi1QQXDtcu6wWCVVdoHbNYRZDuBYtWdL3QGWtBsbWhdLZ2juYNIUMYNccci7hqLZ
Hk0jG+axkkxGvMrZ6NQNwGQlxjSBMBPJ7ETDY9LRLsKXLavZNrCnLypgGOKBqByK
6erG/jVbooszv+hOozL1Q4HFR7wHIXej37JW8xmZvKt78Gze8tzrNWjFDHE/WNBo
a6NUlbt2cqAuO8GwnnLk+n24A/Sj2Tu8N4JngzLsN6xJ3wlFCC814d41HXJaeCIq
B6QaLdwUrvg4/mzEwEe5FDU6vhNW4Jo2lJgQxnSak3yrUg8e3Xp3LLv4KFNGslMy
9WgwtCgKl70USfor6J+ZWCrKLqLY7fX4wdfnbCrtX0QsTwMbLw8aS18qjmUF64ep
KgN5jg9Lch1Md8+V3HzGjIuqjej0jfvpOF8vuQmFg+dZDE+ebegnUqn2NpiQuPv/
IGOkWUjAhEbuB/UunwvexqlwTwEoOoYU+0CCwAI96/y7XE1lPl1CIJSrdToOlF2P
yyYVphcDuDKsVCRTW5m2n+6AkGX7WFzdB+AD33lHB26LUkiI40GzC3nJOxHNoact
DF+7TcJWyNIgmPtnmoptz9PlyFsEsHB4DDIPLOBklzaKW6bHSXEcPoaxZ/1X1vsE
eh9ZR+Kh+IJQPrugqZX0chWSbUXV9I6sszvS+UIEnTgatGNPEU6blRL5/LvA6zA3
ZIqxAzaOED9MO6yg4gWjn+uCAroV/q1/y695z2Xd9cDGGTXUC1/mkg3oA8HQQzMn
bv88CFUskEF+gPMrULvetcZUTvO1USzA+DZuomF8xbE5jU0QhPCUIfsHs5fRLAK/
N07Ka5HAK2VKF39R3fNNRNthtSiY5pP6Vwkmh2q/aHdpgQUp193H47qa3Q8tNJoY
Rt+8HI2WBKMekNUsJuHGGKr3zfMNSvcESjf391BsfFg3URlUftS/6VkUrr/9/9g5
nNRZnKRnAZVN608mA63B1/wsw2Hh72FSyUIxutx44nmX7+2Y4m1as+XoOc+owsrj
B/H56U9yGHa86CecuDM/cXQhFtaOcUayKqTJAoZaW4A52gu2R8fu8K1zbLo4YYnd
N4c3ZMEVls+tSQ9NPjrDrBzR6vcTeEzIY5mbN1KWYKtXhTmbVGWrID96dQWNEfX5
sg0f1mrSBrG/zXux/a5GhlFI2nvnvyCRNwKF64mDWA/0xE77ds78D08gemHkhINM
ZfYVhYqDO0InUK16ZyEqblpjwhUoShq7B9Nha9j3nz1yghroEOvJ9m8Ng8zoILl4
QdlurrV/trVM/aYQ7HUqBo5ggQkjOm50991fNkcW7kT7MImvfqLS/dS7SpR6xKFh
ruldaic+dHvMvt0iJ87frv4x9mslWJQ/fhNT06/eF+/CNJKnofBjy+BY/SJqNe/Z
UJhk6cxff1RKHrVC8ZKdc45UB87fUdZy9yTDmbGQQWiK+GqWxtmsRj/p1EoeV4DP
0H3ql/j4oOQufg9wstdemq4nHJb5UizHeRWcsPvL0whK+0wgPRupCqIcnV3iedi9
/0N2KyxxsCF2Nfv8QkgreiK6YtABKloDMyumHctJcmVpSg4XCrHWi6aE/6EA19ta
l1MltEquhMws202PZN0U5Q7O3Yw0LLkDYvl9iQCj1zc=
`protect END_PROTECTED
