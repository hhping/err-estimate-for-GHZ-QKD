`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LKPQ//L15V18gYki6mVnDe1m/qmVfrCiK6tDJkI51FnpnvQ6l4JLgORe3FEeGxu
v05GRratpXEQQAW4k9kUQoSyUhRU260DJHNx4R2+EkBNUPx4wfr8oSn54OXH7KJx
FOWEuyWthsnVYoAMS4UogqbnV9BiD4jdEa6zzULDHWBGJSNJbLvxxJhdARH7r1Io
c/nenSIJMM6TGZlF+M2a77Fe2nayjrXxBFRmZImfSjUMGEiphMs6QiaKKDqkyQqh
wH1rWcgFHI7azXN2ByX/LLPz8WSC1CMmaMCwXDEtWWfBJRkUL8xH+N5CmAplp0dG
lCMy8utTLUgbrMB7R/Us0gl4/zog2l+47v0lJRGQxJGz/g2nObRCsnZuKLXKmKbx
y1xWrumGhN5T2OlNyT5TRJeDwWR/oFPtnIQ9cAWVd67k21lPm0NNAS4zZw1OcS3U
WwSCrCf38/pkiobU4UfsG5VGhcVhgDmKURoy5BtWFE5qG88T/qJnD9I8E8iXxd1m
WYQWFu7GV6gf/UkueoShbeiid5Jf5LQAQ/Do18IHyx50tniR7TXf7wg8Q1b+URiK
64LPXhs1F+V0eujsMV+bjVhwpTkqv89pDQ4r/gVdm5aBRokBUofOz1eHTDI+5Uhh
np70cso1Z9F77FVHUhVCFMcJ2XuzzB4hSUmKoWBBi6RORdDsWLqHXOkkjI/WB6vP
uBGkJsesVyA1PN7nhyRbtHz4iYrItbWZG4EOQm+BgfcXroGKQxu/wbWRFNZGaOCa
r+ramdEXUyed40De2L6/8uTaXQr7LcwlhL8f2dq+bF/fjyGBPNYTvZYzkgCRPipZ
Mtf9Y6vMmthrKPxLHL/gLJ47tv6CWM6DiPG2fcqZBPtwrJpiwpmREwNOwkOH+Lt2
S9H6aiJqGEmSljZOw86rTIWRhZa0nMGjzSage0HvuPZ++NorarfIpwgihOZFiQIh
isNRysSPeCEAP/JQN/aU+g3uCZ6CVbodIgwIGkU6t50jfVWJSVehmM7n/OHPAdY0
RbZlTDNXP4OcIIlreq2K3DYdBLbF1izTPrnu+mf1MTjS88EJcRe+7aZfHjVW1y9P
jJFHaSWusw9a4xO8jf71aDL3JlvHjUH5+kYyeXOqEl3gOgmuc42Xof0m01YGza5C
tky2NTl35OPI4QzZ6XcZO04MDiEGTItIfLq7pUhtT+RmGXonkfZ/YbHaY7NV/txR
r7na2oBOARX/BvDb9O3aRYKFQaw+gQZRmF6oaWHmCG9cTQsfmQ9qtpWug/DRbqNU
/MXk9NAIyNxSWT2T0LZ9NIajNyopmi5bJEy6Kelv37hLz7cxGeWACkyINv5nd0g9
TCJosbMUThyUivRLGFuqGnIKd0OM6I9Jl8Y8ZWnWJGJf+Ec24T4c6UMVGDliyKpW
Bsrrjh2kAo6qZ4W0VuRpzcbcvAtRnvJexZC8tdMJqoOrLUGAlhgREOPWRxV0qRM3
o24czYhoqo+ACFQlUWSpx+AmuH0JbwaSpI+AnW+2s21GBaUgXTyKQm57VTVgJtcp
SBJLSUXR5kICaTR4drIwJI7ppkudfHDC5oz3EFVumNqx46tBczOnJ7pY1793ew8H
qY2sXl1kKttC3rXIeeGwdsTF7we4S0BXew3anOdJ2h2JKrMklIB+Ucg/EfnJUz1a
TbAJT/Oomv/R/I/KO/B+hcpcq1sp+wYX1c/RRLn+GPLndLXFIbnWati3WQwFYrFT
2D81/N/4hQCRZgdj9+fY6P5UprODsKWS8ahswPG6CJydBT8Nb3LcgrkAimsgBTAA
5Un9ve+SshkYQbdpVUAcJoWmWiiWnVpiH+NtrMGmC1+hz0ayX2D1zcTqlnzMtG79
koptlmbtxYVeoFnOWvKrenXuLVKZPlIM1uOAV9JifHNy9EtCstaL1FwR5E4MhXyC
MErqZAvWDBGX468CKOEqFlmk2qye7szde6mYnyUgzYwIWrBn3aKAwY5Bs1+C3gVo
6wq/IuhP4VP9GDDkHTEO/Eud3uoQaPQ5vKL2u3fYLMWPl2bbl3EIZoYu3VYIFiDb
tc8Vrj8UT66zFoYoNJxj1W3KZshJQYNXgxzD+PGgIYgUjlq+bTlyEOVCxsiUUcj2
jx+8vqwEPNDwkZk27qyVPmqgUL37smSKdDHGkGTsAeyxQeAvoJfznNgMipGvIMfX
46J2u47+Rta1P4RFYi1YhNojTIVy6J/mM9SmmUyV0I9F08jNMC4i3Kmm9jUBgIET
UKhTOv3fAsa4u4n1dFYbF4o0HuEjxtMSpk9OpNNycUwrIsYYzESAF64SFFtftXD6
CH99b8cUCGFeAFZLTeidHqRfBglJBXWV5K3dhgdouBg+WkUz2Pq2THiL5jOkhox3
9F2EENN1uKWbvM23OBnPCdCj1A9XAxBThk81qg0n0wT/CWifNv4j/PbgAZAfYdYv
PQKcg+ic+Bk0o7BrnJbSnocYl5jFKUPKq3zZf5ST+UJtlmm4Ch6Mk3ms8bYMu6x6
NnwjiQpwdcqd6x31I2WY83e7DlurE1lEFkeUsHgVuvxBAs04Fn2O+Giz8iXtgLma
0rdwLZAFXJOqhvwkPfKNBsGxyY+9EC0Nf20HRAm5l0zpD+ltOo1a3owrfEaIjKb1
o/DV5G7id48LRBoKaqBDcW3W+zCjaJKD7xBUxe5fFGGfUaLHJi28SvIUquSRhP+b
SEcBxYkWQVZYh0Yrc0Cqkl0AFLF+LA+wgsP1Pab7LyA1tSkqcov5kVoswBlBNZ1r
Fz4OFulYL0qbGDxcaGSrZC1423CGZiHJS3bPmoRhCymuI4MNmv6ylkLIwOOKdJUI
XQQQS25VNjGdJzDeNJBwSuJUUJD+MvzG8GhXcHy9se3o+UqQYBonGORIBlLxlfVM
BSvCcW5Aq7Me3zHc23wcYPJUW0FjI+WJuQ755bJXlMY=
`protect END_PROTECTED
