`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0GIuLDa1QmIplnVBXXtpsyp6/SDmamPnvU7/6uu433JEKWE44EHURy2OSUfiEVA3
QrqeRb5J8SG3H+0beP5HLDCfIbaYrn8J5JX0PZLCvHqBecis+A8A2FUFsI1PjNJ1
hDslXFelCEbjUET2m6PWrJ1e9z0Sn2tKtTyJAVER3q9KV2PtA7tuYbRjDwnfcAP2
Y+AjChdf2UESOKtXbNLHzS0szCQQEUD3084IQ8s8pMv3QB+cmSshZll7/axOAnti
EbMLrKchgzJ0MWhgwbbA5FKk9NAXJqJBQnisRUH8QuoYCf/5ihpZSwWrlyAtb7hq
dQdGvxIhD+aXGSNC0nJK5kiQepjSvYraDVz5kD74HTMZuGu7CpU6mSgrvDPh5aCd
WsQEzkWQhN3zEr1BQ4WF8YjOM0w5AlzujvEo0KE6Cw1za0+qSZ0p1FF37VWVcWHw
Jy4xRYo/DHT9UZoRc8avxlmPNseHgmUcqxTPLMuT15Zf6LCxwUhiWWz7pNYws3YO
8Yr3A7uxKsFsmMvKdFs0HFr8YXA8K1HIxqRnY5Tt9OgNzykSOwxs7TLOatghDKSj
fkANaCUZlMH4Oy5ahlvMR3hiaWliQCJMMCGIsb62yDqbGFqzy5eTAnMrt/PRkq5S
ooRJNvL+5e4hDgQJynsHzHHGtEIuRsRoELsvT1wXK6WBkyMBJdzQduUWM98GI+Eo
UuakbUkSICAEQAfmM31h9JPmc1GShRjxUWaLfrqd9Dv1g6hhtyuPg/5SsHJHsv8M
s6L6C/hQUXklfYZwIyX2c+Y/0wDfBcGN+GXRftw5iSx5xrGHAetKw1KwrcM8kzd3
aIvwDHfH7c0ORIeB/8+ArPzdUdcd3lOl6nyt8lMN/CTzEymNEhREQ4HzsaTO0PNF
H2X9h53hD68hwmZHtIJqhILUsHQ35/mR3O9mUJeIc3/wqv5sW1jxrG+VmpIBZ0xG
E73rDYvBISWuPUcALWXKZK3PH7oNPR7KHOupkpA3FzzRc9JFRVb4fPYBogxKUpIu
bTi5s4iOQUywCUhAADTSu05x3IXvO8o4411B+uN7F/BpUSEhTUeqr9c6HuHgV+ws
MHRF256JNRftxuJKCKzg79hBX+DDMW8iXJeB+aqbPjdt8gu0Y8Gov5sFz5cIsAKp
Mj7qqZmOmSXQHsb/gVK2TyudvkeOeQF/61pggf++O6LNsDTBXCf+nOyUwd2LlIy2
VTERXL/L6UH2SI8HXRZlWd0oEmGKZgAOwYVmQiC8TVgz9eyy6D2l+clML3zxBURP
4840claPhbeCRhpD3ZTZKJmgAIemAqk1L9DyiKgjgoxuK3amPgGEDJ4/LAPSifPr
GwijsNjBCwT3T4ee32RVxLOXEwAhJBsS5FPd25wM/Bq5aOa8blAnQXHWMMBZU7QF
P7qePdH6e9z/G4lnbbrJDCeyyN7mggFbFdz4/AUrsr34/r4LDaRYRt9zhMnBC6Zn
IwH6yEX4krjAhUkynotaR3cRVNrvJ1D1n5j18Y8aMMVn96NoJlerLBi5UAYEVfV0
zpZB/tUG8/ckdOuGaYXXIdyyvlsKbqit3CYy4EmfWyIWrQB6ybKyqP7sorb7b6uQ
I6+R95k1Rc9NcFq+hGYaM1ZfLDiuzeEDM+8tvUEMVHQARYvTZbKPncX7cUY0WEVg
`protect END_PROTECTED
