`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qeO6+Q3un3r98oo9Kt/o/fp87/jiFbbeCXSu0xZCc303l6zfsqMxF8ju0Wr0zSNY
KW1k0IryLAI8TOZMa2luI78uqxDnCK852upOufJibRaE2B0yNGXnH9+wuQ1ehbQ7
gJXtDCvc96OCjSypeyxhZfYNGH+tF9BaVRlX8MvMQ4C8TZzr+pSFOChupSM+VyQC
GYlzonytDzrpDezZsS12FNVZaPLp1w9JRfbz7xjSENBACj5HTBAuws4NXMMQm6of
rAVVIX3kJqsBnvaS4h9NzlD3tgVB3k8gcqunREJhMV6McFsX7ssjt21XA+w9CgBM
swc3vbUVFPtTJO0CuTL0jW7tXX3p14EprFz8MSqtoTXntbme9j97bf7MhDTts6GA
vaoPfLJkj5XUXq2SKS1zEA==
`protect END_PROTECTED
