`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYZJjiawl//DSd2ajNAxLvI5ZP3DGZzUrhcrA8IOHm5uXxgkccBAYMJXiiWEQA53
ejtrVZZuZiWIkU8P0PiugO61dJ4+7AR2QUBF0QywhugW8fQAIx802uYWJ17j1U5h
21+4XAqTKQmo9rrYtPH1WiEG9uOJfxQ/nGj8rCULUazOhgvJzpcnssPEKZblevc6
+FTa2EPKE/4WBRVgfsQOjlrntBjQXdlwgFKcuLKLOiaScpI38vN11ElZu/n6/yUy
7ETxbb6rbRenqTOk/oc0UUwk/c2rsejNT14Vy3onOFrttX1bnD9wN9g3P4PS9CGB
JoUF7wpqWYckz6bJKKnpv7b0HSRMYr6kDnW089pAe10bXJEE8QTxd3SO+xsO3AWF
vfF8AIjKeIj4yEWfC/ktGMdmYrGfabh0yiF8x/vaDvua6yjD50rJ/Chjg+EupwiU
8Bx5WRAoFCJT0dqh0HP87PpvZUJU4VvxTxHd+W+aEXKjTgCMVP2hn3MknSIRWuIJ
NoKD1SMd4LzpaF7IoYlspIxOkCibHtYRgOTnFpu3E8lxR3jg6TGNhaenGiFvq3ZS
YAvnz0bivnSFBINI9IIny6dpBS8OHgC8vdfhNZPtO4P0FRRFeB1OauZdijvKE8D7
j3bdgTudD+mUbQZpiBae9UPxCQqIOou4tYXb++WUxHg11DrH9lucAA6IPaQB6spw
9nJAB3BgggZpMvIU09C83ghOhAgzlE9KWdPVNlafRVT0s3cNqkRsEdVqVfdN8vAP
8MobQcG4M5zfTevqbiKPkWlMEAujVS/0u9p0GqvpTp32lgwLZq41/G+GrQv8lQNH
qyNXPWC9BbWZmduoYRk9ur3KC4xgT7MAdfd/TDWdBgo3GOpGN5Kha4HTyNfuazFy
IzBh3uiwwDtxzZJa0MiTNKSwycHekaSzfWBMX+B43j9xSD+43yaLGjhBoU8pCddI
+AoJg8H5JnB9i4QGoiw9WVeKqp0sIxoqND7rAT7bLci5ybJI9pSXio0BJ1PMrOru
mxUrr0wBhSMEDWsmphGG8y3knBs+TZnEzLrZz8ft4N+SDD43bU4BRe/zuacoByYA
qGX0ZVmXmEiAi1EMOBJa96vaOYdN42rIpo8QBT8O6TW9qbGoFQM1n2uX+d8aVzdo
mZSaup27JwyHLSchr+Hxgl3OtheTiFHC8ZdTedmw+N0AE7+9Ie0xYPSkmgfMz9hJ
evpN4bODaskvC6+KzRcy1Whg0wcgXdZm03XF4wI1tmJHqaLO9dxJWQSsryaiNGXs
75zFbprEhPfOIq+0vp3d/1aaDLhb5WCLBerT4qlPTO3CHiJUlmmXyuiC98Kk8nnW
9vmW5flOpQoQ6kC3kDJH0quFuESFvAKBM/Y3e0zriCdj3rDVQkrvAxFqiNtfziI/
JJh7LsPpbIqblYTuq9P1Nywr2e/nJJWLhZlxJ0NS3K0m8OQh3KVGQIcLmHYnttC4
DLl6vRfFW38xPbM9Il3pNjk9104zVIzJsQzja0YHWNhE79MbbiKtIbBw3rh/Xduz
yN7k9pQMXRhh9T5NnG6rZCYPZM823emaPiTXR42Kvqrw16lZNtz9Ki8t63AmCrSl
2dhlywAu9gKg+IRnndAOMnM7sdygGUZFcpuRbsE1v7xoaplyg05rYs/1d4hGgQfO
W/0XEHIVazVddKNkJM36wWHpiOxVZB7al1DV/jtTTwGk1PWfPM96+fxOoZ86YTWy
mGCUBLh0WpC1pZrYXuoI5r+jpE+xsNugAPuKsEbmjUrk/ZO2mQGO0b6SwrLOnYpG
1sdtKkek0dE1mKkvQsbxsYIMF2rlraEfz1t8OI2+bDrM7uoG2qzltgSD6nWgOuTG
dDxO2dNdZKm051gWzXXdtQCoS+zrMejQZ1xAqBrjyIpdW4UfaKdm8BXoT0PZdinH
PDhx6vCKPsEYb+2lmKr269Nrs+BmulMt4W78C0X3zhBqGI29CWIhZKrrgEl3Ejmm
EDPwx6wFumiCowFxAqyVv/uxLfFcamJBEOGVPnbxB73IVR8+ifL5Z9YHswp9wPC2
xHFWr7u08lkvlJiHSm/aA45M2jjI6ip7kVa24kURtnjUKgHIq1A9FfJeBNIZuCVp
dJnxMzd7BaiaUsbwx6RW4AW5+dHzFXmJg4vmXSbhxlSrYgdLEZfhWWKUz4VyotX+
onXd8GL9uJWXsux1ibNj2CgZ3m1aZ2/5KSXf+SY5KQw2SYZWqOaatbWI4Iw+/V4p
Iux4z3JvqDE3fmmncHR7mzQPKsJomJyusCCQEd3E9JCrUxJLh3KvPaQP1ic1fvcu
lStNlwKLSRieItOk3gVL/rHX94Ol5LglZxA1ZLGhO1rI/+yWWPCdfAHfE4zRE3oe
bWXEZ8a4TNAz5rsibbUYKQBoGdtux+p2LYZ35UApucAE5Pf6TlcSbfpdXtqrys3z
73t1WTdkHp8zwzFI2E4bS729vGEsKvDAkNH9WOSeb5N+ICCz/gLLHPakjchgSf3+
K1o2YZcIeBhdsVD9f0zwtqmmtJ1jfDmqe5M51O7DIR/ffd2x7MbDz4q28tbLwPU1
Zzl9ezjNpJXSzFsyJF+HFqXHVrNz98M0PfYfdBR5/ouTaw9erQTNJP8rzz4Ie2Gx
WsItDmosn5gEQYDOIygLXsC3O4BAPG+oQMGHLEWM4MuwfAr9kEruybN1uHGaydGD
66ky+k+ewKrYShM8ZJLABwgXVm6M3Tk87QQZzQvDfHHzQNYFqNu0UP3QlznF+LtQ
F21vZvLJgKvCFdRyt6g8R9antoD97m+PfujvKsHlt8eP42paNBdv308WP8g00vrR
VcbVKeCqJzBYbVE2sLbeT6gTkI/qGHCVD7yhQ68sLhpiH0DkpHItqfz4iLC2H22G
FNycHEEOWA5b74lptLpIOFT1GNoK01EuN9vjJACimwc4SH9OB4ayFCsifp21bT4i
zfX6cCTpZg/d8uBnrK1xBfAIIMUJnrMR2PAXsGDmrv3/h2U+yuAXe7jz9UxI4n9A
l/qN1P3a38FZXYVFDAA6ZBmZjghqbdNjFhgcFZR+Omsfzg4tfvvWetE4tasp6SFS
13CqoZaw2QfXsDYjpUyWdK+425qXdOREkXpj8eCkan+G0LqlgJp/RBMrLX29eGih
wBcYdQpMpPEtd3DnhBSM8RhQbxDZpalH/tkG4SIltU+9jBkYAYVQnad4L1lSwJv9
BQF8MoIL3lIUTid0GcoeLQ0XXaNt0jvK9c605YpSL3EEXnv0WtZ6Tc5+huN99768
NFElvhwqR/BuNHwLAe6FjmwTGsjZp26mRsS053C06MVrwtfPIkG3Ni/bpXq03k7s
ElHPTC0Pt43vMJy3iXaxq3s/rCVwZv58FbFG02ci3iPL740rmnCxg5PU6K6xWJ6M
8UZ4u93X8IIpQygdDHYrKT43JgJzPqTJrozINKCEXpqH4Ksp9UOkW0bor+l2tJ0e
fGdqdgIPk/UKib7Fn4Q3gn12ggNSk/txzo0/R3VJKyDKIxtcywaVElnmBET/EVvP
cvYOCWFCsfGPf1YyOu+gvSS4uDgMQ+eQC/YwDjwWTVMIr34W3uLIv6fy21Tdm1jA
OTGAcfG9DccaHOfXy/x5CKxlaJ0HCw/Lldet9YXYpQ76m6oe1JqwKQwm3vF+CvhZ
Kxwgn7gumln8EO1ZB5MC4KKVwJ/HLtk2HbtQkNFPgFnGfI5UXR6sH1Ad+UHFb+WN
66hSyACq9I31thG7ViBvthycVMmUNh80VSrNLmkjnZUWdg/EWkBKpI+Im/aCTrk2
lcMhdH7EIEOojL461/4TZtPCnkKf+yNmRLF3oxrokA3bzdGB/BPnV+ZB6yQywTBJ
01Gk93QUFssA1lRUqzf01ksbeGeJ0HfEG3WgTJptswpGGibpXeXhF8K2jTrPuHPN
6tPMg/2VG3Yj24LWIt5RA1tMCUG3uIOXDwj2VujYlMOA2hdvRqglKoEGw2cZUQKu
OzfDkaj+KVzl1pRbG3bWVqIu4H9/u84qJuQUz4p4KNiPB3e2QE3hfNqP3vjqtHAV
N7u004IA/H32zyWg3CTdFiRa1mii+6O48ZdWX33ZQNx/clZb6YRzpNyzPygXPB8G
2NYZZQmWtp+JFA72tDxK3tlJqmduJkptalZrvFz6kUbCCfGCKlIACWL2jbEi7RCr
ZSfdJzd978jIMK7CzEDflCKDlQvbmoY6cSpxuvmyD7uB/dk2SlvlRbFoWGBkpZvp
HOmwMrlb+kfUAA7bmITsrzErNU8I3Cx5t9iw+aGGaNV35hrFAWsOz6N91kgK1cSm
MV6iHR1NnRWvSalrxIxhdg7jQsTA70sRDKTnWG9YX1gZDz2iO1UMgiJzt0443F2r
OjPncqiuVLzm28EFa0onk14RGwhBHmwkYGEIt1rfPZKEI/B5wrwWznBge3inUfRk
GS06QFquN5yoNt/S3lz3GG0XBNcoiSep0Mv1aXR5XFXzPXDkKI2ZVMc4Yoz+CXm1
tCeHlTxhpTRUJzmGDlc1X3jaKr/TX1rp8UbEdv6KQaZ2zZ77gJdNNejxBHMm17We
GKq2XlIjwn9vbAFcAmBx22KmahLciqKpyyZmYugd+uXA0O5RFDo7D8clM0fOC/bf
SWojIK6XPSQKmxS7uOWR6bgliQU1fUJSCzf/C5cPxjeBzYPxGQKrnE6ixxtixAqj
vbW0BwXH00CP6ZnlOODt5P0oBEDQnOGzE1o0m3hnJ23LZt0oJsOihYD1U7N/fQYx
KpGOyCFSs41RRJlLPrQ2WAxSSYed6gmpPN3OSW7/uRCWbG8fHi3dM/fLa6xzjttx
7J2O4417a0VI2mMT8A6se/pXPs41r3H5dQim9pkU7Vw7W50HbcJHrORcn1eHZBdK
UfxYIs9X1CAPUtisx5ru9xe51aY6nLupcOLnsCLtPJs2NyL+jWLGSGSEKdginwD7
R5vlFPBr5sCyJ9DN3WatxnQUgs3nyTcarMjBraRof8K1a4a12oAyorBd6GrUmJ1q
TVbkYBwag0xZJXMoBk+pZ5rAt09ofAK+1f3F46jfL//LPH+LVutEwa4rXM608xzf
ZBCbHG8e/wfzHyVQVXqgLc9Pu9VqJSvMlAjXv+MgSjhwUT5cyME2ty9EWSE72GbF
qVU3pHXXQCV3xA98rnm9AuibnGyKPn3OKnFVSu4vyWC0z5inDhGCm+2wGhthC/+0
hCyMOjsgv+NtVelvEzn2fkE3iOV3aUjQiyevY8jqAr0v6B64QoouI6UJVxGBTANM
kK6up9ZUnBnL+5BM/MjzxEofTKWLCQ639x0oUGiWcQb3KFbGeDAWpCIjRHhjjdID
vEhel9m1uDvDOCKKt2V2lltl1bMf2IOLoEXUX+hdmx5j+XGfd/xH5iuXKQ4R+OmD
8HtUOfqwSSsOm5bx6OXWxFh2oMX3HhdjfJITHT6Hg2BaR2/CerLZ/eIsG1+U96dD
VA9+yWw9VCw/6MzI6q/Yu5vwtdB5FYvK9G1H4m6RW9FNTVyh6DxSeoJLjftI/qbv
UO2CpTy8cSX3NhP2/5z7GtMjGS3hWXI3D5RkbVxlcAih/APnALJQXX9YcMlYIqE6
b18X7zUaqyjYhjKcjKmdmikSh0X+VDwoHXjut0pl3dz6L9Vrx2SWNcQjjUNgBA/l
pwNCzBUjONBU8i21vXDjom+Lj7uLTqEmAY7uj94gud7BXDeofAvkCAjuX2Pp5XYw
ATjosjnfbi971WEaHhaSdV6VMS0fL+Q4F/EY0kEhsrEVm0S8YueUrKRrsw1KFFYl
eYKZ3gCvloyPOZWy/BoErrncl6UhArdozy9I7bv1yxeTCa+U4vPzBeSnhnfzdfu3
yzB0K1asGnfekAKGD9AmmUuQLqWojWgcqfDOiG2okeUpqYNH8g3L2IjITSQ1KPO8
kP68zZkoY1WDQ7zmTTbwOcm9HdVcklYlyY0LlHHkSE0ESu/Z7f3mmn49RS4LZbSr
vzW0OUpTMy4jQNVG1tWD4ZMuIkV8QchwCbaHsd9JHmZgm5bz5LZ68Q74EeudaYST
nnBZXI37k6t2VcSO13MncTDUmfS26qO2+PeLTnkb/Pgn6Rb1iXjMXBrOBM7WdlnK
bYFmAQBw+F5fSSL8sySv6pnHdkpKp37HlImvQeTQPKqYLlXnjzQ2VAC/ZT5Yhrqw
pj6B8nmfIxXKJI9KvYIf6kSZnUPZID9JKsmeTr5j40SZ9/naCcixzADS/X+2fqEN
zAIM/qcaO9uV9TbTWI2oVVsNQnhP3AUS4iqDP6TULXcJR7Xn3YlKMp0/o0xPTpIh
+s38t+rkFyPgQo3+DMazWtRiiDMBauyfp+kPN6L3Lrh9a/oQ/ZG6HVfHSvzKeHPz
uzBa26i4i/MvgRVPUxlJjzjWt6dvf+ebr0sd0x4MRoFj8nGwXKkrkAvFL574lscu
E+888iaO0kGI6L15vBO7/eijW7lDEepZPDKi64UQZXEmRl8rRM+d7GbDfnAvzEJg
+Np+ziIHcDhZh1pxjRm0W0C/Ep4qqX+ARZ8GTOI/kj5zL9430U+0N2EpcopKKDaB
4dXnWbckCVMH+S3B1461OfNu4o43NHZEhaHbfm9BeKKjomtnlR4tOA3ijwrca/E7
YdtY7X2VDGwZzpUCZr/IQz6V/GOKTC6sPq7cEy31UbUt2RPZRLUmp00tiYOTf8I3
wsJG8Ik+nXGxSXTUaEKGK3ThZObB8MLWxMVBcXDnfnhmGhnwfWmZ3KpnEo80fE7J
hAgsggah22Z6Sl9jxeyACgB5hTWx1CSxEkh4/R00kKmlwKvC8h74NbZakQXodQmf
hLR3yl31kIJkKLdkI9eXgrua2hmamPeRrmL2hit6MqkisUF4BTlc12S/9fPLx5QE
CCHYyflBu5KupRY41veM1fysLGR2+fAX+sUTCfnzadJznbnL1+cVHSVLQavCHAxm
/imDvKxcng8OyR/qTjXkdwbPcip/1vLRGv82iFGiaeLXYyEHTBAN1k3PTiY09xq2
daRDfaJOS92PI/ZQff80vZQEo5ymrihUP008IClokoh8f/Z4moaRphr1USK+1t3W
HMao+AEcpefe6/rhLQjh4nV03zrU0LTM+mJA2cF90KQRxMnqY88ZveLe22IDp75d
27wUAiqATdE01J7vuYHktTUmcLw2bQwAildnRHkgfXWacT9WQiVc2OXconPv8Bt/
qbg8oyBtY2pqaG35ClwlFefkyvzggfhyKDlQa5E/1l1uDXdqHbtpgBD2t59VuWM/
NEoFdSvMm/3rAbdFK2zkByNjcTW2XFpoCIcVJkI2eN451HdeXRGmmA356MbGs7f7
F97Vkwbg6lTOD/gqKjT5pFESUcXGbcSpNAZFjNz5JEyiWK3Yog5hzFpR8t34/exo
6wFVcPHG1oCEi1Pnxvqp/HPVYexnCWqHgziF999QI2CAqmKImvx9MxMvLJ0/nUYW
Mnj2kLmzHPZbyKxUCBa7ShQwzVcx2yTwOA+ExaYJ+0OswbrFpn2ZLeD8MkL35w8d
BnW+7MaXAdWrRajYjkzIuzOkfBOPzQ1Gbdk1g1Ttp99xr68xruWAlcbsmoL462ej
WN9FWhqWGEqoRjTBlc7wCckNuYsmkNM0bUFNfTg8mzDNQGVi7pUGv/kOK8fSjoIX
IY5PwkAPhX6rysxVv7iNIY8p6YOr9NiP2sp3nJ2zUpL14IwFJwmO60e8f3C6kGyb
l/bkumYK8jhVSqMO37v3d+Njo9+IGpAYP9WsmbcK4v3w/q8biksjIqsggXmkzonT
LMYftMJx3kZTsQe1O3F6C7EMR8Re9FDcd2IsvQvxBTND2qxNpugKOkco/Eg7o4/y
MkbYcMqczrayLP4xruqsRDu6JU8ymCkLmXu+r0oWQ4bpQ4ErvPQt1bUOwcosH2+V
rSHGjAKJkTchD4StZhozGHa0XxjdrtwDqDKv+9rQOB6d0pF8kwyqLpRzJ3PEySWx
FwxHdhQPxfdHdmNZuDsBzDYn6H560vmVJHd7FCmis5FT0a6Iz8H7I55FftC+XcUW
Ipmuru5lu4IDxfR1Hq692FGHDCGmJVrcrWtvB6P5zfpAG0rkyq7sQi/YkMWEsdyJ
VvoM0fVm+PDpFGdPfbCPcq0sERb+ovT30xHktcSC9Gf4ZV2w5OHy8yr947FPXpep
7zU7y0b1hoTtNmo7GNcLNfr4j1bEsfyFmLlWM9MpNfrpnalQO5FJU1EUR33cgtym
n8eXlSgKAOg7rOpjBnDsz0A6V43NNnIlO30ezR9iaC9kQkSn4YN0OFX2kJ7hhoF4
TAIVdMW8+06ugsrykIL3viyovB9TLXjiMjkvm2czOguziDsdsbWTzjOglsZVnELy
G80RYd4j3LGp3qKbdLwmlEClay0PY3skHEa/enAy4W2xrmlfmt6Si1F5/KYhTTBb
tNnP2Jdx+WEJcJQuQ9oAyEdPqJ/rm9Sh9YyLa4qTNnOGKgKrOeqg/+rXYpu11Hte
c9AmI30g6Am15c5+uI8JID80UKds/TXwLlUpR3wR5eKfabQXn3nE88JKzA8n723a
PDcJLmOtQJYcFlifKigaPwHEa+w1G12WmzW/Kqbnm7yjkevOzVWnYFwfDjKdi/EL
Nrj76o+Ys2BVRw5VvYqw9bzHqLuV0LvjIXCcIwYpoh4VTk/HS2gF4AfTKZYvQF+y
SP04lvyRGLxaxCj6F23Pz+7Z/iJqawHoHUd7IzHMv5tp/SpUXJ0XUNsgisLFmZMC
vwwz0AuNPIRwhs1wiSw1CIKcX6zTUitTqpP2WoTR9zk4OrQSAHpAdLSbp4XMEI4Y
qc/v+N0hBp73jrTFO5Wh0iij2ID5w/ooSpiqwXUS3lW+h/KAqdwU1ZqHp+plmxtr
QU7F1OXfQRvodOwHkO0aU4GhdsZ7yCRO9R+2WQW6pc2yOLC/bdZ/0VL4QQ/VVpSW
qbY1bY+d/fdwSAoIHolLqMj7SAmbAMQpYttXV5dvIldH4MuQ6EhzWgnbL4SrM1Oj
r6KT1FmmrmoJzKt+qzsCHWxLICcBRlPRkbmieIooaK1vzgJmEUz3si3BfbtBoli6
9xqIvj4rGgH54xwPKdGA4eKNZLjiUysWkozQ4UQ07qvBvaQHJGKjSQyoo8Wzmiom
ek62KXYwaJa1+K2iJYP8iEuSrx1nsBgXpeu+pYeOAzkWCfdctcBig6FSDz2oUQRr
mcz60CkT8LnvGSZBGYMkg7CYDEs/aQ/tsLzbKTAyTrcA/9WIKA8a0U0AL1xEJIIj
z/5ooFnoUtwS5IrKmtEvyqh66GV6ElWCow4gfDIt4mTtS2KyndgDV+wHxxQQv26r
tW6LvafrW1uXmIF9h4fylQ8o5wJNcxbn1atffFDZ/7X+Ismrpwx6BzTD31uKscFj
UtdV4PAW6bQfxmpc1Q5N3somKaLW18JDNe8ckFbNA478Bb0My+WRF+nAY6MJXp/p
CW6hdb4hfmJ0LAqezoTTgxf04hMOKIrGqJNLNEPT5Yg9Qhv3kCR80WcAkO66JryB
PQDs8UTVt7omzFkxw+EciLT4oK6B881AnTJRQKWuEuJeZVc7tQX6zSp/NhDuaf5q
hziUxxWSTfkh3AfgFej//ZJ2fOk3Wu8Ip6Z6vsb+rWbS4LaVJja7KulLENR9rm9H
aj6aparCRtPnF1WUl8hczFFIWNRSTxoZU0uia6GyRMsxG3a5+K+vbwLOX4tOqZw7
iUNmS4QfNHi6sg42ePueIoOCKxWfRG5AB9fkInQfbZR8mlOVT6zpIDetqLtlLjIJ
KA2tLu3q3dvvFaWgpCYFH9wJKwxjs5IvPMJf9dMK8JRshlmjia04tiQU5Fgi9fFe
ex11SYJMTYWX9CyCLxYJi659yiBef/fCCWXwT2ODNR2K26L6Kp4HVZ076hCPAWPw
V2E/Anp46RsxbSvO1ty7b+QkTck7y1IRE9zQ2WXmA5jgF0elrll+rZkGYG+0tV59
vsfaOkT/SHPKUYT7toIXgX6BdXUPJf2JNlSqqCsOl14NCufM2UyQdaMpBVo4QF4L
1lL/EJZmM6YT5Rh+ArBP2k61tX1V1nu0o98N6vR8+IXgIfL+4lteXihRkrdNn8v3
35aU+/wJSwnY8liIaS5wnwyUgIfpgDdbbd1o62v8IBNm48jyZc/drYBvgK6UzWdP
1jfH9c+DZvWmYG1J7VRnR/cQS/9sG11TQK/Az1tpGVWmsA+tBZngYx0qKQ0HnhyO
TL/vYCSXNwQwuAsRYCM1RFaLPpxGKDIXZPPBSiNQRnuFFUiEZv5+WasDVurvsAIe
4hW3ku6ShPaFT0XVKCsfe0so1Y3hePJYfSrtdpmYI6OHW/JvVCYMmdc6VXXLBSC9
zMs/3x63XnqfEi3qqF6+hqfmqiwOBwecOWE19oWxPlUjNhh/TCHbPmBJkYfKKenn
HvNv+QJs2/yMHnM40JNH5tmdNeaXLceeV01B6uLQSyHHve0/bWY4jn1HJOICrW6F
ov+4odNIaJEsxLeRfnec9iMprzd/rUo/1JYbaMUlLoRIW1ayjmwNJ0Zxw2rCpreH
Gy9Q4gYmKJIurPpnMWsqgm5KRHPIeYkeChbLQDWuTHyeyMJfxSbKr1w+nMPS+40X
HAKiNrDEvyFr1xkyzYinjtVBhkcYZ8uYteZFBP/UUR4q3P4tbIrxnwLTZ3uYJCj5
mCnal0fVzptuwhVy/5wQtl4K7nQsOHkhOUMsvIJEbQ/HlZU/kjO7D3/ZQbMPQmyc
j6On25b9UdKkPVh0h86CpJq6KAsF2nyGKrIVHGsyoUJGNYb5Vf4g+yFPWMHQohxV
prgZNFcxmLq81HRDDn54Bgar3l3/pshPv+hhmYiX9fm9+/+XZQ1ljhH2jxtuFbFX
jQ9MKATR3PlIhF6eTE/U9a+yO72dhIShBQm+mzYnjNXQlTMeDPpcnw1ADZ/+ydxf
Vee5t9o+KpInZntmnJrYj+zMHcXeZ+eBoqrtfG75rAta3bbvbNpmFOuLVNOjuHLW
REqM6nuoB6rI63izZtrTbmK8UwlaGKOxeTl1H5XGmUtaG1Rp/2Tjjq/qWSI736Gx
mAxxNu76uIfxy8qoTP0wi5Ia10l5iaATb/5C5VRoaLZFdfjnvQzRimXl3WyTDpLY
PjZrBhciWLiyEFLP+ZiZe7Iac2TAOdHbWO7o75hZFphb+Fxe6MA6foLXCEBn4Uhg
iTf2FusOSECmQE+Ccy5hKau7SLnvl8Kl+nQK6+aNoXP/S6BCAI11Ik8/NHYuJuH/
kT5C4M5kOYSqwJ6fFbP/HWgKWbj/FIoUx0Lt+lfhtgD6UjvbPvxRxKVt4zClCWHo
3AfxUdShvil3rjHXk2wEa0Tdcejc6swKPqb+EaWjHGJmfJNQZWf3zgEHpr4u1M9k
0LCx/1/E9kmfiRdn3zLdTe4JNPOzRXvBswsqJ/MM2DsBuPK9TZJdNEflvAkvYROA
D82w/j+thUH+eV3+nNNFn3mMR1Vgo+yOWNXIsrQQd35eOhaPj2HobvAm88Q/T4g/
ArnX6xkf1qHY6AYieMWJrjnWyh9q0C1XmsDpiMLAn6XQ9oZjlzZv3vCVxpMhFsl5
RLbK19Nww3cic8NWnmwIsroGePz0U2uh+RwWo8G4OAKgY6aaHMxw9i+CcvSDIq2o
mvLXaipH96lleEuIlFZL3sjwqtjkNGONv3VgPfFG9ZQ447KjmGiQWUabAf7cFTeu
0F/W5PCbJyWjPyQRtQXXq+WUI+QB9Rr//rSDeiLlDdmw929Ny349IiwG7YTaRYs/
q6usC/6dZ6WRhSUv3lyt2GH+GfHbUev7vU4Oyg3MzdpYvzWYq+GJkUjoSR24PZj9
kg5elNopVh7zVKS8R6BFKNzo/lbU0jGBvWWhxiUusexULf2YpWH7B9BlEYDdXpMN
UbkaNSOpOAcvtqdRQvzWRtFe+6pnJH07lG1tvhCw984dfaLHTtZf22ye/rI2SGXs
Fk3sT9eMLwets8w6aJHzRXHy6VmCqChaP1n0dZe2kphaEU/ux5lAFAoW+J9DmCkC
2ZBGoRPBGh6rdEXoM9j5WKctIumIeaT49CwrRlER/TuguwLq80OJGxcLJlwJA7LK
D8b8HgLuOyn3JJbCxAJBDxKtQEKvRIWKO5uAj1RFK2AuLsmxW2Cs0r4SZvEPYkkZ
X8fILDUQfBL6Wg3i1vwHcvaf5zMXkSh069KGpGhdXE21Q6uRYTllG6XmdQsSubeB
gUdYOIOHfuoVat1rIu7wAsJv445bjEjgV8ZICtw7m0IFrLskvk/zkfBJlzaF4ck/
7YyZS8q9Ktbmj7/L6UvXwyyrxJ7D4z1TQIv48YNP3/FZ7TYclPXp9e9DsH0YW/O6
vIrvd7Fnok6kHYMT8+EFquv6tPIVPhIRol6Rai+4rZpoKqj2jXR+6yN/uvyb+XzW
Jbv0aTL5qHTEqtDSoX9rs5nEWGqFSb+BHC7WkDF2yCiKLT5Aqdg7KSimj42lv0WB
jQHzvyY1K3bUObdSKLeT4CxJ5TDnN8zMIaF7pDew2lUVjTUT8XU5YLZ9UJokv0Ja
NIfAM0gbsfsBVu2KN+7dvfQV4doskt0WVO+/B6esoEXbwbhNey9glazmYqoyaqoI
/dZTb+dlrp4tUQfUOQR/0gbZI2Zdjwdu1aSDPRH5ZYoU87z5oHkq8IZEc7qZqueI
vJJTlh5M15c4FVV5b6jnv0l4auNrONYHh15Oa2FbAu2lhWwsoCm9LXf5438ioecX
TtpARRRAbqzEJo4EEa7n3qtwq3SOUkLNaKYl1hStNCD36HikfE0pWbMC7sgmV6Ge
ckNYROX4XgNQLCzickJ+XaGukv6cMSU3tRaDG6/ydhYdw8NA5n5IW8zD5o+JwaUL
rSaD4/iJzZEBWUwYIg8v73c2eDF/Whu0y8MgWxLP0nJGSZ2KH5Gi/XzqOY3lhgQq
Qcy6KAeAwxmPdHQOGWjR3BPKiO1kZVN3RbauR5MLe0K8twM5JB3juev5xGElRsYu
ZevXf0MwM3UWvxA2Jk9Ifu8Rhu66MpNRIIKNJL+MiwmZWPpnzY9mNV/xB5uS5c+B
duHJmlwzJT8zMJHnh06AXOAaSqMdhiGrGT3XWSiKY2TTb+hvr47ZkFazR2s5fG+i
NisceqJczw+A/4FtN02h5u/ZZPU2TKT83LdqFTePOUFmfKFg2djAotAI6hc/ZFYs
yCrbtDE4ERI+9pTqgKTbwwfWmvLY3mjZVtlmoK+xmNK08kHYTpF+mBwzcDki/hzT
7Vo6xemBsWp7/sjRJePlrbvLQfqUmkeRzRw8HjejpAouOXcKmYS/WWE4zuN0RxRu
LvieqMWgm4MDg2/uV1mYr0zUmIOoLobyoqFsuPMBdTk80bPX1x8TosgLAFILjTIY
x5noxgnRd0Djvnu0oZObv/K7Bk6aXw37W0dtBSjBvcu/LNFFlpD21vhG09H3RdtN
fxAXahjVoM93MypJH6H8bsp8Q+ncrHPVkkp4l4yBcwPlu2HuDHEJ5kKd6mNbPYlG
Gabjhrfk0x9OaV0AmviHSS8CdOK2zRLPXN0vcYH8NNgMXnWcneKRrlsc+SP0cnuy
YGcQ2NUeuKByJr3KGXnhLUTdczXQ6JSc+YcNSBZlI0j6VKsaIvuNTH7Y+dv3a1K4
bgpOxxkQrcu0beG482Wx//MmEdD6fyPMWdewvrwl7wZ6dZLaNwbny1/yeqaFTeh9
LvorXyUXVJw0JBRdlTwEXSzxNl17b38BpA+sqKOzB7werIeYoGX6aZlnlZPAF2Tv
4qhPlkf/VmTb06S1Y/tC73mIkdrGYXiTiIDl/Br65kowgqOxhdDDKGoNrHxP8ihB
43VH18WC8UnlzrsGr2MYOegFgKKU2ytyTB7CipKTuwTmf5f/tqckHZKiyVdpr8xE
y7pC9uA+bfAhyTxWp6Ob65PzbDWo0kcrKZKw8PvSfq9t9EaN5LT7Gr1sNK3FZuey
hZYCaHKhs11NWFQqchAweRByI+7DFJ0/g/jT2caWszht7GI/qL78LJ1StnqPvqmS
fyqOPH4KMPK7FWNXpbLC34U7f7mEFCWERx7YzwRfq7bqFfM9qc94HjgIcw80PmeQ
/gHr188kk8+/ACvXhGNPymkMLAYfNYn7C/qu3kCC5zwYoSMixbPcS/6ii7HGmkJn
7W4tLMZki81gvhLetb5DarsG7zj9uDNv/uGm1p54l1MlSyfHSq1tRowv4hoBY8yj
fmBPNBAzdCxvH7Yplf6qSIIlyvHNAzQwxOQexX46C15g6qJ/JkAYWoyTs8LycjuO
oc2rwrRQ+jsltP9n2zcaznFzKOTxAqS8dU+NtOJVKAyvLhmt109y1+270dpZIG2O
GQff49tHzM95O8juffzXgg4tScFHOFRhid0IyGWkM5hmamUOy6c+cKzsEZr74Hqv
Ka2vJEIYW5tvmMt+unZZ+t4gDeVzlKPWSFbO+XWMHzaRZ2tJYq+tRd6upLF+8quS
IiwROCeP7kLECw25q095EKPoXkMruaP5LJDM/BeVcBfZg4qkresZRFUO00Y+eCOK
AR8qR9sDvJfelJji5CBH/CK7pG7h+ekwdgGNiWFXf4EJGZc6ELf55Z7fqSn3luet
cUyIyW8Auaa2aAAJFMmA351aAW43Fgei6HmtfFlBox/rKjOexCAIb6o00o1T5BFs
I+R7C4+Dd2Ls5B6v4A2pUPIt3oEgoDmSMw75zoaKbNn5QPK0S5tmY8zC8xYAG7UN
jmZ6kKVRw3DaSkTRuModhCfH7m2Swmo+7/+b49QePGrPsP2C0+suzmTRFT+Ntljx
Ze9WbkbErfJb/7W8305xur3p5x2jbPt5rrNWhYrQ3xcpmHxOEG8tf8HN1OwmFxMX
Lp8dk4spezvtEHrXvhkdSLI7PmbRKWuMqANIizYD2Vl34VY1bZMA1qF7x695sVWe
bowiNS6UnoAAoPCI1y4QcQtUsHXt1GaEJ1U2+Dk3hmqiNJv1OJPJsKpbVy4sudD0
xIzTxhXihi21aJ/o2OWQ2mn24FXISr75VvvbxEKzuN+P7WJPLFd1uOZi7xp+JTqH
MfUm3mlI7bUenu22YmlzDictsOnHbKEJdY7fMH4Wi09pS/nJydCG+msyS/WsqpGg
WD4CvBEexAvdwgLTrpSV6kGyrfMHUhH1fbbrkZgYNFJ/MXxazh8C3ZlJUYAOYR4H
Bk347+SyJFdDQHeX4623n9OXT8Drgao9pn0NO9PKMFpZE+v7yRzk1GaWRdVVSjJr
Cy3kjjxosu86nWVafrshCTrtYd4Ap6CRnb03XmjR1fgWvZgxqE69AimrZq9vjODK
j17dXrjAUdHu7YCiAFY9vODzIa8Gro1zszz+OeB3k50lrNzaGhUHOq73fJe6OurS
6rOEqF7/AHOVTQ0f36o1T/eCs2qhF9WlJTD/cr9JdGtAggxMdueXA44rmEH0nYrE
uKa0ibKPnGpNHrlqYljBCt9+ILPgM09D4i1Ndt0rg6kDR/tktvJS+1jE40HWlbCn
bL6Ma5pd4s3AROVTOONbP/orLqnAqHveSST2V3yPwm7iXAdhohtbjlrj4kaT4hcr
78RVncHgJQxsrwHJmWDDn22OUPFfXG/K00ckPFooNDVspooAK3qQTrocU578zmVp
MIyKlGkV4v3k19Js40cIQaeLAxK3cSSmfPpxJvNoyiD8LnknfdJpjPGFFLvAUt2X
qyRP3UIxaP7Wzc0wLiMVYZE8B6VL8pHAh+47NrC3MrLtwJRrCAvQs5PmFxSsbwKF
xk0IoXstUgCcIihJfinUvAhskzzyYY0s7gYbUPzyOw0HWwtg+XvnJBt/VVhdjmPw
WbCmivQZuhwCU5HPosTFJbQd1uDr3VSCZHKUTQXXeK1qIsv20HAQYLjV7YQW4JBb
Dnlz9A92eZ8qeaG5UFFqBWYeYbGWNlVd7FawnutHmIHyESHIagnPdt6rSz4W1+4J
5fY0r3sQNLWUMNag4r4YEYZeWsn1FKYfeSMs05CskpxnwEiircYqzEUK0oTzZQRp
qpe49DfH5VOIonSan6LHBheY7s7W2StMhi2r3jFM722lu/l+7micEGmIxBjLO3e8
rTxNfnXcGkIDPl/1y/lZlhQYRTS/Ga1+3mYcZWP372Vfidgm5Q9MAeK5IZd59kdm
lvxlfzR0TDtzJkHECGNpQLi4J8CcPDh2It1IUFxz36DKiVBcxSQm16Lnfhqo2/Bv
xlONF1fT0jSlbCAyf+2kixN0y+noU0664dVz99cDSa0MEdvoU1hKN/2PmymPBLrS
LZYZuU7cUIlrCTYoqDDxB9/l4F/s1us/J7XIToTqcTSSVNrVuuWjQHODc91NiW0a
A1ODH+nCbwC7QVq+uLYtRdhnQ9PyAXNvB5G48VIv36IDFXk6HSiEbZHZ/INz9POT
WNNoUsAyQfIat4vQn7yfWmpUm+rfSlbYI7pyK5XdGapH6nEfRhKKjGS6Y8pjJ+RT
iExNAo07qh1rT41RKrWI0xyMaZ1NakiRkA2cYVD0lV3U+O2AjBiB6N07/cLB9Ykq
IFGLP3H0yCj0NNcbNoYm8RdgglK2rxNHWc6h/RB0v8KxSRDuincNVvnsmjoC1zkF
As7zYAE0jco7L/ar0Hvf4c9hEdHr/Unjj7BRvtqMXkKpz/dnBahB+QkVOruikmTg
02R25JKy9T+nYR+7v3cuaTAAzfPdamNM+y3z8dM2BI2rvRwnTx7Hb3/p0Qd5XoTG
JxYWBybfAkW9PTzLaJMsPM7W4iF+krKZGKvrwN43XExdAuXhgd1gc34efyUtqg89
bVATJAcXwOBXjqgYhDUorzgKaQ7okVHH2h8sQhMhpQeF+N6yltXkRhwtBgvIRVB+
zI8UdrA4S+G868/mHOGdisSIRHdYCJdfYicgLH/zqzmDwD8sirrBcFlAT/RAcbuj
nI1IjmvC85dfw8nW9sHxOmuLomHQCYNNgHzCXMBaMAeZEnjwM3w0U14Yzp9WUaKz
Kf4Il/FeHAwkljCy6y6o6c8QMOgS0Z3avcojkuPYMmeqHbyJSFHQY6TpvWvl1Ftd
6lEi9LCn/BEIJ7JldPypik9GPJmeBjYB6JeP0dCiaUxDNAhnyBq+FjM1+6pDnUce
jpi3sDg4gtkV5JChl7t6rdCkUoVMtd12+32IQAwsRGoSV/iUMidlRZ++im9mjF+V
xM217gSb04E0k5sKIDVvnzepLmJL/q9gbOP453h0Odd/lh2u3qdaqF82X/whVhqc
zpNgmbUsKwhoB+k/GKfgQnZWvL5oy1N5gqxXVTDbnbJr8brcZ16oMPxDI+B0HaIx
lwn1QxtV91bpFfrZsfrFu/D4nGVsAZsh40f0CNngs1zGW40bjLbW6MYs7kFqk7ND
pi499kYdcIdjG6+IAAKN7wE8zdSbkTUiIQRhZO8Blu3TQcEEdVRMhbMR0Eaqt26B
lVoOg3snBHqtvwd26KGMCKevDv/rYQ/EdLSip+3LILtTAdNizRmUyIjwGut6o7/0
cWM6GF5euQleuNsQ83eANjUQeTxWO+bgQVP9Ijjlhc3EcvWQZbsZkB6721nXOHkJ
8x6Jdqb1MoenpOnX8TtB2aSuTU7OZtzvkda+S8Vp34gY0Vnhwu5H3lQrQ7sZKh2p
ETOfwwpThcocmlc7nAg6FUeIolJJFyCGXv/8fAFwwP6T0rcKPakEnZHeDSPEmHQS
8uKx2JE6P6OIzH+T7dWdJUpO3Tc1GWxLGWw8R+siRRWTUuNcQStDlQXwUe/cdGCi
3mz340PbMJwSUoiHcr6Wfx2tdjM7s2Xmh1UUlxw4jL9RTlXi1Blt4p24rXrwRGFS
L2ivCJqdXyHs23DOH6e+qqHETQhAB4fpN0c9hAyNv2N/Qea0Aol0uPfrF6/C61tG
ta3btw4QOR36G21T7Gf07HGyK9ZcZhdbLUpL7ym4s/qhRTQlEmY8x01EcWaLTqLI
izu9Gc5HCT3XZOQt+D7FF4Lq+maB18H4azWSHspd7L4sua4hWR+ZuRB3fg1KdMNr
nVKDn721pMVu+Ym2+lx7g5oY419fqZvi/zL1onxiz3aWdKWqEXyd+3gNvD2+hMd1
TSOm9fuFUPdaWdGJ6vm/KCV79vp0HENFd5f01sihwIZT1gAPVUUyXyE1zuwQQjzn
cQWKPAJ6vmesOrK6qlmGjMCt6xbfze9WWs0B0yC6nkIPCJRE3UEdW4RG24AXP0Bf
eSOufArTKZrQOJxUtJFFrcRK+ALqaOc8oNGF8Ghi0DsCGiE6G40al+0tcJkXy8T5
sWh4bw/Y2Uv1Z8vzxYxo8xiEm8a37TUQD0aoBg98/COftdnkYZsGB3kxhxz/Hw7K
0MDAg5WdNoHl7a6CMITrtmsRDLZekgIvhCL+EDasBTXd3ahuOk65JxdCGqoG/qgo
J5ddsseP8XeyLbjw/yllTiin2/mv/zQAVtXDC9piI5LLKTUUrRPYeV0aggN4R1vD
TllupBgSGESXFBR2nEsEXa5U5uoYhyHaBq9G7rJY/soHv2FgLvqpTTPg/hnTbLem
3EjJZFldkQLxGcYqHI0vhkexmdM8YdAIBUtDhuBl9Q7ude0OSp24Yne1+Ruethwt
P4+qmTFd8gGjNF2T2b3cAlEwNEuPlkdbcin2llZd5H07acbQrLq8tlQ3RrBZl60K
PbZfQtFFMlk/95wUSFTk/Y4cD+8HPkBmDSBQ+FuQxu1W9AzGfsA9xyLECptbN+EJ
x0BzpSBKACqLw2XfG/laeEyY63gCpAp10CMfUt807Kyd26ewP4h8mIiBJUT0l1jy
LJjxPv88i2E2hMU3l/LpxJigOJjaVZ8mwWA00kJof+1oBQOCNl4h4mCQr+wSJc5p
scVFOBd2yugB2iRwhpGE+B6CvYoYX8vPdQPvcphOACYZymvSrRXe3Zo93djJgoC9
xtJL8kGuDT/q4QveGFJWRteyHOUNdoH4R5uuTlZS+SBfVf64O7GwCvc1LfatEDZr
THMkayAniWIYTuyctzVbgBhG2Dg5cA+H/jpESt2g/p1ANqbQkDodnqs3S9103ta7
pVRTFXDymulZEgvsnMT3WvXppX99S1HK7h0wdR+7vWpWDTmr6om3jTS5peEIEdnH
1fED4anJ/PANvs69MA8jO4dPgtJCyF7giAfchsa5xKKrwx6hKyPiOwWpRg1ZeFf3
tVciWYP+hVYEYaoK7nmnALVnLxMwb2FICmCjzpGc35CrQwcuv+0vmU3I/mWgLad5
j/DvJSSE81AzYfnsjfpw2Q0xAQrXy2Ezb8CjF8uCCrzcPlwmWHk2Q69t1s0S0JLA
OmhKGqzUrLZIHHjgW6rEFHVPZu8E/JHV4ladE+3CshxAbEePmiljnejj8kP7DQb2
EWgiaXmyScaC9K1rwSLjhZ+XhHU5I/9lKOfoB+BVakMAN8Jb6OMSWyVQP7wroxqg
JK9LDbBnFBuKrAbmv8XfksppV2uiSbI6uP+8Vwcp4CkCkw0kQoebXO2vDUeRes+d
wcHudCsdX6BypA40d1K2pyd6cWDjSTBhd5MdkvYeb4qZ48qs8catkb50qy01GxWu
Id8bjwQczCCqhOpt7AlC40RuN5hV451qEK3GHQOsazaup/0VCXgUXMfmSscI7f3I
8jGjOwJgJ1Yf9VbBeEjxFKdfZg7i4kNbaIN4ip8BnK9fWBtVCjCIrOEaQ3fUSDYN
TBwCpgvRVZf8fY2Ll1bSQemajRH8TiwVObx5sgvU79uTdqcAW1+uQcWNKGQQ2I2D
zXxJW72MKpGGwoHdXzMDhbsVKDo6gGS0ekjwwgSjpKAtS5oIQc7kI6gfNvulGYa0
1ZDyAjoaHPFXDwLbrhFLMRiI/XeAJ4u4GPCuop1UxasTRAyQhVBzFCIii0k/WJsH
wE3ao8m5U5MY7b10HOkzmwoAbUMQ91c/WmTpCsGXFxkm6qBxqLkp2Wy8H+DsXeBV
3v7Dq05qLGNk9jweTZtskKjsSkfG4BStoXWSkrowWNVIZ0j/gHOqOEeH0x5JomHa
g7ArAi9FUc8RcTpbFutufw0PBDi6yQB2Ohosq0iZRS7bzIrmm1wR7tUdv5aZbPsH
jXu0qa4Cw9Rx5Rds7FHDKs3PymnP9fBX8mp7haroOIUcmpI+owt5ynsBDPIUBqaF
/VuJnALzHkyHfWZeQIvb7Zye3DOpBqVZEjca9c2Pplmh2Kw8MlqjfAO5QJcS3PPu
NfJWh9b2q2pHET3KNzHXxGsR1TyHRPfgHVOgKaAT8Nw1t/7eyW10gXgvauvnqi+v
H41Yx98jZdx5fsvrCRqBvfwHh5VHmTTKgGfHa9wWlFX/JJ/1btCgig4C5VsPQ7Qc
TzwZ/eArG+MD5mRytte8F2IwTMgigiRKVei5YihbF8+xFSh5Ed2Dt6+R9NJTX5He
j55oKERZhnCE4YN01bsoQ4Xt6dFkMDZpSHoEvxZMzCfnEFjoY8aH6BNa3fO4K/Na
9010SDIFf0i+Xux5aUpTuOuji2PMCloGkgVfs4PydRYajvlZM/qgz65hHBhCjj4g
sWjCkSeKR/DB2VY9dFOfSYSxUEOlmd1B3w/FmxOX30UKVMSX5kpjga/saU0/cIG7
IbpMBRvFxlKplOR5OPqE6RXL2EMmLdcOkfsvNZaWAG7IUOqcKo4LzbYF0wFJE4f4
d2wAqhIVWHno8/HQW629USYf6BvrMfE6AUqivb+mDqicjy6APEv/W879QpYmYigK
Y4IKDNMiCb4tebflXRvPhH6feDw/CMoN1Z4UNH/1jI5sNabxn2kuRTYeCPawMHWI
Aj7TtP/Es/vlNRQtNXbaNXL0MVtfIHFgQK41dMPT+IZ2G8eD9WAmLfd2hXWljVcA
46hM83Nl/Jt63d3ZSuMEC7Di43j0XESVqTGaawRtjT/3rxO7DczC3Y55ktQMvhXN
O6IR4WNFimJAXDkovRaoUUeHSVy10cOvYE4/Ps07q8nbWacS+UgNfFeLdPjso4X+
dDnLg6pRzAboCUDoNExVAkDpZL0TsY6JuksJ4aqfadLVhO51JA5nup14AJjXKDFk
Lx3ua3uH5mO4ic98EPOJ0Rw1ZWw/dS7JGJiGNFDZAowQSfg/8OI19coLb1fDAIy3
KQyY7kPdsKb+L33zl5InKcwfVoUXOJijfWv5aWar9vQfNpgjNHP0CW6MVjZ6vpY6
aUBQWGaxLCHUMjAE1Raql1I8ckf48INwGxmIn4fWrbzh8Cc2cp8vHK8+As+V4aKW
BlWwZxQYrzh26OgYO49GE8A4gakK5nLaKKHwTDz4PA5nWNmRcwEtCpCnyRY44X8m
rrkoknxbvGfc3Mt5GqbH6OAn8464a/fTkBz/YwsOuKiQoGRRtEDFqD3pCvfrMM8+
UpVDpCFab6mO6SK8Q6dAOwfaLNM8TwgfxlN9HQ2oTw0kN/Fq9tNFSKgUyjuFge9r
ysQ9wdZuF8Bpuep6VPwHyRstuFf1RKbb/Ig2bbrwjqKoMsXk3b2uPAtt7PEL2e1Y
Uy6yer619gFoJuG2gRZaYKlpBVZKNVSod+gmbePBhKn1KkiDIh4Ksg0redvM2u/A
NoHIUysNRetF7XJQkp+PHZB6sMBth3D818WxCBDInVZ/Iy1eprvmTkcKrgz2fpNz
eCt8iI2FYZ1tDA5rS3HNxb3FQgIcxeWrCSu1CtEiXJW+pBbLQEVKk5uyaVPmogiQ
VxfIHfSwOqT+0UtP0kUA8XFeJhl4Z3AweWDCEHq6yk61dhOyqLzCWHt/NzVBSKLA
8XIfdU5fzrUCkH+PLPNkemxAyXyu+5HHZYkHJd/cvRHtKKaIUBRwfBpLuIZnhWmh
v4XWqRJ5hijMaZB27Ul06aXpUcloZu72yChOBy8HHyFDXSPgcMFfdD6IB2JW4G7v
aUJN0sH9Nk7GNgDcnyfWaCNSLUyuAHQCOw+/VNtJFqeH/QnZwo6uzO8b45GrHlSY
FNSAc6c0s/ySl0Y9PAni+hb/nk9B9RIPdkoJ+qXiX+S+qBvlfr/twA2NJDmQCti8
sQXYI5TfcHE1LBWssJEtP0OWWDVKic3l3lN97CKP8R4Cd9sg95mQhHT01f8ssDx4
30+gTPTh0Q7GVeS7QwUiYz288IqJzVsbDZKRpNAjUNr3cV8RI/r4YBi6AAXZPHsE
jtbSANzE7hROAIDYDWvkGtRIs8j4yw+CeEsxWKPyPnxtV7d8ZoWjPSqk2LbH6Ig5
DPQ37rzqq6cW0fA6+PHiVMZS2YFo0fPL1W+K7AY1HmUJKGXOdmKg3QW3nl29sQsr
7meeXPAId50aIYpR9FPVf7BGY4+9mbt7SPEgjKAep6pJgPbUZ+jS/2q3TNZ+hvnt
PR3/GMyinlh0mSrUtaw9a5D+VFZEcySnwCHUHkgu4OSxyTcdwaKiV4Rxwpv9aTgH
6W8CBIJlkj7TRnM8/ZHOEtzHeZPaBnScXzp/wxbpP+xGdC/2aYwooNSyYEmiG/XO
v6buWSQtv8uDIkmPUEWGhVL0Ksd7iREivMN/mDYiE/V3cJQ0vyDaANAb03BrtCr2
k2A6134co5wpiDgF1JM7RUUzpTEnQNEgW2ZRSkht6W5zDEj+GjqELxJHiq/MOuLs
0NjRHXVRk9oVi1hizU+qVzgctzkaZPRbNg5Jri4qE/7qgDFGv9xeR6s0Tn467FMp
mKZjF3XsfRrk2sTfLYE9Tswqt5vQgvPhYMbaNz/2BMSsUaUbDL8yVy8raF4cSBSq
08L8V8imRkrJbp86mnwNiLp++OjuHNTi9b1HC+o7vrrTjlg58MjEAIIxdhiQQO04
NI97TGwtxw9LWv2OC3+MXE3D5+ltRjwZ3fOWfMSYEss52WCkpmW4be2kJs0SyO3p
TTvs+SOTLvGvYXrWCrOzegmU99fX0g0SvOAFOMavkgfZJFPJYNid3TbcdvrbfOcA
+lMyIgcAd/mtK201RzCo4+HZXXOwuVNtWSgvEW1xU/nMfnIPRY/nW/AkFbGUjjTl
UHSTKZNkVg69yVDeyhzQsFTc1IeJRsazdUB42eGY6TOmc+8pE4wYtJ15sokKJnKc
eoAbv2JxgklrcvHPCLrWreK6sWuoQQsRT/Aeo5Var7Ge/nMcz6HccK2XRUFpkec8
o42OdKxVeFCicmq5pWZUj675TmR+5Cqh0KwAoU8itvn7a4H//Uv1K69Qa/a4rhzm
bFyZSIvrFA9LA5DkHfAxaaiO1u5G03YSffN5D4smfGyRyHFDo5KfEF8ct1JigmTI
TkZkimtDSemwqSniTQ4I4sTxebP80+BjSpA/CWzUU92MyEXuTvlkYaEzFNtAU2Bo
fIpil/yXU87Hh2YVEAe3fdZbEmGmF+M9xOZEYpg4izFq2vo/VQ9dmt6qQsoQHPeK
/99+Mljtpl+08VlUYCDu23RilnIfX8+IfCfzcvpdqjoOEg92by+3vtpv6gxiRJWk
5b7H51iOS0c2FqDDnbKXnb8S36WOA4J7vB/OMJCqxrjHH3BsBcuAJ+ovOLepZAws
mTMV2QKAv6ys+OHEuGxFLJmd9W0Na+UjIWzLBJGr5KB7QWR84g+HSJ+0HL3aO638
TzhvNW/I+Y+SOR2lc0hpUn4m0ZO44RFCG4SrKtKia7/Z8qeSM5DHIkqzFhgpXYpx
yXi7qZNA98F//eBb5fDZvIYmvSSgvmf40KsiX3odsG7PMT0mo+ZlPqSpUUvYLnQk
22P7YSySga9GcIPb3LTZm4LSC1EGuDt2uAWGxipQ2CnbNzagriZodJdH88RAvIXV
RneAG893Fnxk8XYm0IyiD4exDlx/OdYmwKvLeslmz7QnXeGsdFjCL8LUAQij5Ezs
sdQq6mb5O7N3jgrAZrEug0Xeu8K4Rjxta0+GH2U9XzpsBkvEhpMtD59QKveh8hkv
OsAG3q0X7dPwKdNFO9+Zsd7Dnfmhp9n4RHcL2p0rqWPBNtKkcTBpk91tyTk5ehpp
MCrlZWOLA7n9kiCZRNli8rBAiQcd7UVN6lJikA20MqJWk4BWupOaq97b/EAM+46X
uZj00Kto6ujzOKA5AbndWU0Yre+jC9ZvahqLbkUo5Gq9SHtJGDfI/FgkmUY/rvp3
CZYXbttgzTZ249AZhqX+4UmEALaWWj5Zi74ExRwfNwvIEq26gDocT1Xwab4iZMoK
MY42NUMw5IYwNhnW268yz/Yn3EFmyc2r1da95LVVs+Bb3Vh+Ky2eY2qbkJy4cVm0
qaRNn9kkgN6DjmmNAPJF9DU/uYuCvvX22iJIsaYxDrDcdjnsBBM/u8gwMAuT92VK
zspvAlHPXptcMhGrYJM7olg9PEmLBKaSh+NzpJ8r9AXv26ij3pdH5N7msMx4rNWC
jU+2wbdut77oo8L7Lq4J/5bPaJhoPU33FSFJf0tlgmxlx3XXTlQvBnm/l7rLIj8m
+akV1c2YulaH0+v4EUUSAjuKn9jEFFPnB6ehrX9H0/Aw84ROifYlqFc5YAV6pHc6
IsL6T7mJEKoHY/qnaGlT9k9/6ywVQBvgSJlVITuL39u7hZG/CWSixA1GrwSOeH8l
9Ii2eBmiCgVejtqqRro6fkKahGKi6dYsYB/8JlrEzDPwkNPO8T463EezBL/+gTw8
b/w8HlYQMAU44uyaoRH4B9h/4SBwLoC8NQbK73WzIr3FlOxc6nQNq1UjA/8UK45p
59Bza9+/mOSJVnhz4ANP2ro4H43kIt5VcLXrYACt24p/dQdzzUmtmmTLQ3MZXVnZ
nJp+14jBJWiuPhYvKyoY83440eaFYlv7AAStLafgaWBa5vv2QxlapDO6TfEKWs+n
7KNHqQ7lzfGUpeTGLvY0vBEFK6bnAW+ZOcLvQlToN9ANC1fD+Al0CX5Xb4/uRWZs
y9aBXu195GRxU/MVmmfHtGbNaTSDYifmDF3mQFP/paN16FNy4VQRt285srZrAvRT
Vur2kw2VjARs7AsrkHWAZz/IxpBS63empvgoFIPuaJRyslEfsMoJiO3SGw9TBBmV
0PKDx1PQg75Qz3Ge7tyr7uigVYyAh56uaCHDg4Bwwne/5Hi3ecPnlMCV48jDaLsJ
lugClGuZojOQs0NqFVjB7Hk68lJee1FZCNThstdvVjoZ5FnrXqkqdzFFDIMEZ5dC
UHRYfPekrxrpnwX4mcCK+x8NOUuQhNF2h/n7a9D11vQS9AQEFTouH5px4dbmAk6F
dRADJJFW6jYVDnjOYJCIYDuhjf2WEEkBw2RSwydoUJ3z6ecgTLNzHnKs7NQkHKwY
egiQ98f7iYxezex7mq1vnsVmL+5FYZ8ptIlmUJHjU63B8Rtjr6t4S1M5yuXYD5WW
io4oREH7BQ9LRuMcpTcpY2S5PpIbNuLfVNteqwUFaBYBOW7IxOkkyIu//L9mZH7l
Si/NwS4BwFjoD/Mhlg+VedzXc8F9CFqx3XRrKu0JzZleoj4Iwit04IR7d6D/50AW
BqcmVm8IGoclEFTHLJJy1RYU+knbeB64FnNpNwZtwe7Ao4TwD5mc+w+NpZrADDqj
/VRpahh/Amc8fTc3cy4KpM/0WxLk13QX6pDoEXpjwLDAAmeCceSMiRX5V88eilDL
YF+QfD8Yuh3OKLhzHbHTqHPSFpr1PiS5HDAjiCiBd7sFmTt++syrZKJVCHPVbFEI
F0Y/Tge7i0qYYXbPH1M1+QQNyLEBwaQKLGulPCZ02oYrKYiXQXMNLJVQM+79BVJ8
eC7F2cCpYsq1vu23uK+SswegC0mXsZJkDBMnDui94lXqXxbLyOryHz2pyk6LCWDt
9AgXoXuydbj4ZnF3+3yQVG2nnL67jqYUHBJp5VS5N46/s8UfGyLRrQoWtmlV0/xp
F6nQgOpLCyIMBJJc0wYoxSfdh52MSoQhw7QywS21na7U0TXSEbh2qtaQN61hRrHT
QJyWuKI0xRWVR2HjZfGtmBli77/0iKIy6x+CdyuGaVOMZpHM1lF8lpfmdovoaqYB
Nl4rtRL/Pxu/bmNS9h4iedeIBbL1si6geyZE8F8Bk+dZYe3SQe6CidnrBmrEDEMj
hWnpUQNjODh3HaAQz76lfHuXwCAxU4LkRqFf2/G0xnqHeDUFfoOIU+QPnFAPCf62
p2BaGbR+GJ1loT1uaAzrD9VC4U5Rifc8XCBeeTAhtW3gosROnNuXP15XrHk0+8zi
q5A8V7d+JnGlBZIK8j7QExyjYpOuqwMplolnTtBeh9wMEXTrodGRTbY4awSk6lCn
w4kRWCjWo+B0BxV0MF9XP6Ca4ph/JSNqx085zNItJ521zdSAWhWVpJNxaMU716vJ
Mf8/KhUnQdyYTSyjNXiNv4CKAQ73fiL09fWnMyl/kSZBXQSnBB/WPkNyuISttkyP
9QY4lMfvhiMO3tHp3ApPg3HPAYyDgUrtKhc5jyvfMYqBC+nMrvC3p96H2jjpSiMZ
xfMLyLMXVS8sOh7ryDUl/hOxcGh4nX4/nfMPVOe8SoIJiPV9E+5aAxSfz0k4fef6
x48QZldIs1rRC5XrazMm/m4VDNwslvIsNjgGALcqs8R+uJVfK7kQFTjR1vpHBedd
S53Qwaai/Xz0bAACIvzgx6O/iEq5kxC4sUeFEycJgBMbn0yLk/qoeuR0D05Y/Xql
E5Iaxgp2MPW/F0d8Uh6UnlNjxZ8J8lU2CHkDbfzXbPKyKs69X8EsQQABuH1ysG3N
eQ0IrqHvBRkKSPnd9ZqcZL69KDiJwL4JHBmbzWCewEG0D53LQyDXWF0GzH6rJJ3b
L9E75h2N46cDU2nyM92FDu4zQcG619cFyrUPrgOH0W813ryCK9bTpFpQ7HER448L
Bez9rNSig/0cru2OJkvcDJWBZf1aZgjTxd7VksOFQr6wBCoV6L3MLnxtQiWXhurk
pjy78H7yd2QtG2AV7dp4KkI4zg9llkKsKUq4H4jx4JJZIjHSXndZuKVCZiKT+q/G
xk2rlDus++2PO1YqvGPp/g1vJyfxJsP7sz+L4hyRGK1TFxTG+g7HGjyS/hvm/88O
42Tqs5HQfHZRb2QTBni2zPoFH0Sonr+pOdcibnexXK2dqlx0j14BTHpYP6FvidEs
E2KFy2AGGiig+xMuvovgeUla69izbRGm+5vcQQVUsvo7aGFSwQ1c5O5/UZXbLuu3
b1bKwXb+SwAyL5eawZ6nDwGMObi6z4Nf0YZBIAy25BTJZDQiPgyx3eNbO+ceHO5m
jLmI7mpxiQVOqCpEEW0q+ag+O/LDOC2B64bPz3on9ZWbkfq8wPyVUsFl838Y1M6+
ZKe36RpJPHcdRjyfieKby2lt3cWeI+TmEchmSfXH80c+2+RbYmBAlS8v5qPfS3Ac
33ZzgfM6CB3NK1g6/QvEJQuSa1c8uG+soCZHajnEr9c18SUlmRI66hDN8kblDkUa
HO+GQZ8qLZnytgHAgZivb9DV4W6LY6S95omJuZl6iFQ+plovM44WRnISmHMBuoY0
6SDtdGk0Q9j0/x1LvFSCRxxzppxg7p5tYfjq3UUEykeLN/1QBSJkZtfZb5J1sJwA
66Nz34WgQQLgNMYqM0g73N+fOji8KQJpoRXb4ZuQeJQAiVYWWWeHnlRuI0r4G7Ph
yhwH2LdIUqvJwuJVg64ORD34vxXGz6ySOTPBaYqau0O/qFyugXqoo9q2dV/zjZ6a
linhCxzFzHnOxM5kCHhJaJNKcIK5anYCvsN8FLh9P1yxcrSsf12bVqDO/c6pgEsq
FtFUKpMB7ZeZdoynEFqE+i+m1/0cD7/MmgK0c3DEWF5OZV3mLogDoNVVTtUcUqLk
nCrCn+2LT8cpq3COXij5FjGErnj7JVLbTFF2TFYOdOdBeIiRqz3u8L4FrWCeMGIJ
LxjapltTCqDSP1xzn+MIo3dLp/rxNZs8gTwtQUasruWTtUZZRXVLAIncCPkwWqNM
MgdAr/Y88GNPdzmnehTJVqpFJZ/eSaiCzelcqP3hshbLH94DgwLycZz6kc2o+C1B
n53uSpqDjrGGoFoxypmkrIzqZDXQMZ942WQ+Z/gtkoGxa7IJ7TqT5PE0dnoslMx5
0Dy0UTWuVUJdS0OwbmGhsrDQG7NwNqC1/VtYiDcEuHmcJiy5G5g2NQmgmgHAcyaY
FF1VocuUsM8eICQLD5xfSMFU+z2XG7H3/9Jh2F0DSKloaPjohZLIPigjDQv4vVvi
0S18Ljo5wfxkpje2HTBOPTXFHueaSMiDp0m+YVl5Mih7l9LULEo8sSIu9VgZjNkD
7K1Yv1vlZE/4TUaJifMqmWGepiZ9grT+pJ+Xk/Jd2kpksVi7fDrc8H97ykkvATJk
V7C6/S6q3gM6oD9oB9QAUAwQUShY5bk0y7YOuRYqjlsxxd56HoHIFdyp81xnJ0Bn
El+syZGG9SvabTEZXBZqWWNmyxbOLJGTpFxAPG0o54rS3WTwCzMpbr/JWmgWQgDM
cVrjQCzHQ+dKI8zgmaMuf7BiahOKa2/irKZAFzbGShkBx7BQEtaQDD/pikdKu36E
nlzQXxogvo6+JjA8yDafa05QcI0Vq2F9VNrp7NPlCHmn8L2QufWF/wxQkcavA7uK
0DZrUEE/l4MQAeyp/Yp5GSMKLObZ76wF3yxr4U/mxOPFpT2Py+szW2DoxQ2wws8G
R1J5i5cX9VlLg2bOH5if5NxFs+qsB/I4mGVBa7hC2iwuFkePfcEp4lRW2OznMW7X
vvaUaDl9GnIAd8W7XrMAd6UNis6l5TlPXO2nDNINvpwI/HyNKSx84OYTFi/RALTk
hH9TVD9qmq9EUn3igatXEJvEEcEdmgwCqTEoAZ/suH9SzBAmYmh38UMtIhK6Hh7j
rBBd11vTOPP/o5vjG6vg24dVL1EzVCarPnnLaMBipz3AHCRA+/aBVQh99uvyEDiy
wCNrqnihpEn2uCU7KmBb2PzwBUbXynZhzG1P8n/Ex371FoFALB5PUQFfdM37zf2y
OoGhxKOanR+PkTJbrScneKjefWnJvA5MIxF+dN1Si2p3eQ/2p2LF/aJkfVqsniYq
pHsXKZ2HJC6lOz/nCA7El08yB7ruyDm7LGNuiSngaEzlxb2FLzBlBx2oxiodYxnc
uhRc0RzMoKGtRgmQi5ey02u/l8DpSkL6w5lGH5Uetky55Ti4PTCTOkrZ/PYRG4kL
jXjoxcVRq3XJw9Pn/18fv/Jb05ifvczzEeuPBQv729I/68sYI7XR8tmbV3v42wcJ
tGwJZrBid0WMGLD+/TOUMYUStjyxha15WP6kGj6qa7eSmRNjQMGG286Wv9NBsc+w
DGJddU2zMTRXzxKem/Guo8umNwgsjkvXQkHMbUFAJMtvWEUf/lwECmIg42SIYc7j
zRFQRdrP5Fu/8a7v1gT1S4421V9sCT5XBiW8vBDNfQw1r7CFKb+06/tBNSumhisJ
8gk8qFAvMFdCA+gZzldAEuDe2ZEm/SWJnj/mj1D7/s9SMsUF0sVy1DKgrLm2dBC4
7tfIWiSM29M4Wry1cZvDZX36FSln1iNuJ+AdrU6Z3l9izaz5+QhQ4a1w86KgEeEs
RBxXMmEMFPUV7dhhvJ7DFCBocPJwztjr0ZWmG7yHR7K5VDFCYOpyQ96VJb2nZZfU
Cr7RNNB9ODuP+2AJKOFpxO/vVszYKypjmv9xdqfrkA1AIt/8M39PzUNjDe5HC9vb
zCFrBczCByre4FWfuLifUqfNOb7oYtzofqbf7prNKjzPPVVxH19W0YfG8P6Rt9wS
1fkYAW3YwpjT74L5CR9nLrjp5VADWACKPhGzSvXpxVQia/+oYlfHUpMdip7QVJV5
PVxcnrO6ofcQzcketat6Z5UGfQDPLT9JRRI/n2w7G78A6SR4ifI+iPqAX5NjORbC
W6lSGMW+2cnoqxYgprCTBL1mKsh91a0l4ttdKk3Rtt5bIWCo3k3AuJQiPhouwWZY
rpVDP8wODdGRVANvIdO73VxMecq/UbD4XYqhH6FwkkBvGEICWpC2KkfOnFW1tdoH
XQ+DSgX6148ELz2Rt8DgcE7hUts2vA6T6JKZCTcoMrCS2Mdfz4HIRDoL2PelUrSY
j5aZB9/KcOzyTE1y7k+HX2ZhahuCk14Nkk3ZIgdx0YnbOUthz5sZHlqxyDDzMJsy
fTgbzkLzQt5pGh5V1lc8wFwGcInpUnf1qxJlX8+At0WKlYyVZph9zAcvu1+KSx/b
/4s9d4iDpqyr7ppLe3+cdKj6PRBOSuB4sGH4RHrvO+mVyZoJz8UhFWnN95bpRu59
t4OKG+Bfpjia96wnu+/X9a+e54SaGcYHjhETtYxwisSmqWfqAKpCxu20A7eeydbB
upSDBeiae1pYopi27apD+Z4qHfA+ym6IrqeySbJ2HWSoWTJ86GWliaiY7LKJvXHx
mbI9mlT0dotdlAYgosIrBTTrpiY6T4bX/jBnNb6dN3TOJUaCxkgT2wGiVuYcKIrb
sR+lh9Ae92V66tHdZJgQ/imQcPLb3yoQmm++F1HZAhIHSlxb8I+O+yZ83OhBCqlX
lmZS+8obwpkLuJGRaMjrlvLnhbZ15OHT73fwOjcRzfV0L9IWUnmTYySuw1gSVIjD
3X3t/dR9D2qjkHLXyK+D3ifZvTqpL90lFY4AjDCC3WbSEiqLKDx0P7JsPhSQfKRw
CNSNVXkWbYn5TjIPhnygj3U/HqJtJMu0zlR7O/F/4kJsV4rHphrIBybDm30esXt0
wU7+tWBVWzo87JkgTyzMw/VloTLPRxqpe6rsZuSkmHPJodoLawC0wMP6jD5sZRX+
Xi9i4oN817+UietyiNFDlIdVw9xlV8XiAnKx2CxzAIwsyv7uaIDbMcXDk24EAsrw
Y8GHmL4XOkp+59s45u2YmV6g3PglFs8lS5TPj+8LoAPtDhao2tQ/I7oXdv/02DiH
Oh1/Gunft30Xa7ijR+5tpdWqtj6/Y/u0bEBmp+5CYJcy2pboOVNH+5ViTAaUbdfk
7BCLYEUfS28n0ISjwypXkTjcSqsFbiBg/SS+MhpSj3PCRW0Nc/04dkX9+uorT2yU
HhaQ2p0Hwk90mBCGy/PusBJf9pooODqbSialxSxffUd3rlvdl1wPF5WeMjKRCGox
XP9sRXykcXmLMvYNa4y1tA5lnbkkC6Zde3fZA9KOElJuap9HeHex0tII23aU2U93
LQ63aSnpwvKo83CyrGZL9ZUE3t8PSMvTRXZW4mKww8sq8w4CGojB0iPXvqcERb+i
PR/jVkfsgNSiiMMd2tVFm+HfdDumZbE45H6f+cer0Mewvkligv2Z8217QefGBBYf
1jjWEhT0dl61/J3IurERsaF1fCVKRxeyFhhH7dtzvCa8yTAwftvl4GT8h2MitXTr
E4XbAjHB1BhnNnLwMuzC5BJfiYBsmgbfkBd7qyBdJtrkHQdcuyvqogKHSXRt8Zl0
2hy7f+5cuh0j/9kE/pIDYkp0O7eWorw1nZiKWQQwU+KvftO9LS9BxLAb4upzq9Nw
efbRCLRAQsM7RCpbQQwIJWEO5E2GDkzLyOlOZermXNtnPudW9GA1r6eYCGFxQkjo
kyAn0DacvawP0e7VaHtm4KdawHpskq3KRsLJE0LBfkntLjv0sLk42nVokLAFTN43
cXWQ5yR+FpxfJ/HAseW3eoyf36nz/2fm8QyVBriNipZORiwpImSNAnRAfBJ0Af93
xFD++YmW7uXsq0m6P0IqaaMx/rVwI9fFvVNkpvtB7903XGls7xUPQz/4epeoOGop
KZ4kDapj0eHJBDGGQNx6YgYNgHKdBTpksuTC8Me6L06zYi/E8IrZDuQrB8SaZJ8e
93xi+SmMTJ74qER/74aqE7xtx/LznGF0qn2lCJXfpxYNlqV025u0mLAgV6vqwp5P
fn3fV7DRGMJsaYkAZizhFWVidvWux+SL0vqQRG5IXRne0UJob1MBbVe7tn+PHsjU
fpLdLa3770jXJFi6ry7qgINtmxonkNtsMBKOBj9cvD3fn4w4oh3EQEvsJKLUgkYk
D2Q02OxLIdPr+hGKWPlAeemN2dROvwuOy92CPsI4AL0o9pX5oGU3d/cZJAzYSdzC
DgxMN6cZIlWEzbfY98Om1jdF6i4JWCTrTZrGz2b8xG8csDPSN+HbA8ooXtyJHw6w
ebpAyRH4pIDbTB4A9mctd5vdxq2gsrJ6gHlwfEb8nsJiiKvnhfasQ+up9RN6zBHb
smKXzAcUh4qMkrSDz7uqjlQKH/zfQ+i2+eMtLEYAilEw8ZQdIARKAVla+RjxUSsT
Dy6iLqnAErcBxuYKO5yYpPRvoMFpnKfTAT67nBUUs8BysMNVqZQvEW6lAj2H7IhX
P+gVSkJL9Rzfvi+fYnMEMYzM32Oe5xUIJe2l0HSgFjJRRyd1ngowzpiZxzOZKvoi
ty4nylw0rqOHxRf2B1Y2TSuGe6oCSIecU1cpH+5ealcnd6dT5CrhdRQAYnhYhfWq
ZDe1ONS4t6npAHYoOZpxuG0I2eKVH3qchNkIb8MUFXFKWdEhPiA6BcN1EZtrxv+Q
S/zN+l2zP8mGg5o0/m+ioVlubeNI80DPGQM4v/lEUosXNtL0t5SrS6LCo78dwJT2
8jt+kJ8f1bCWZUjhkP+G2pf6YEcSDaCqsdwcXRZ5KQUj1E+komlgMFswvSYI+d14
l+b6KN7SQDwIQavMJ+w7GAnaxZho4YW7RV1hNcHpuNovgk187LBCB1cNc4z2+hPI
aSGBzwT9sy05ZzQFFjnE+CUz1RY9IglpGpBMUxbP8D3p8L4zpJDT/HJ/eaR4LFxJ
3Cvt9xDwV/RAd9rD7jqVWzMzY6qUQgOKZEltE6YEuvdIELEc+SvxafOEUkAqdqMJ
duZR9TWk2dZg8MT/HG31T7ON3dVF71lRiywqH5WK9WgT/Ke+hGpwFfJo9OUcuhPE
RJufxp9hgTRief4Tf0KkUMYVf4bQtHFpGZRiBG7kqqblBu71Lizvl9wvvlq2mSIZ
t8UjEw2bp8cmAaAFPVzqpOJyf3Iqeg/GBjlOe1hnBpsM9g6E1ZtDfD5LuKmrIB0g
eMiBHpY2D40ZijHU4V49O0WXptG9nNnYBYRBNeS7LRnph8SqrVH5PeDTZUeTnReJ
yQ94V2x3ugPmKu2AbQMJxIlI6aVi9Tik41aDxfdcKoOeHkG/F5CZGC02Pv4X0eNt
JcIT/hesG9W5slbYNXbtlIRnfGMXni13F6xyB12obmuZQg+r+yWrUyWHZ8rPB21z
4jabNc9ZQLyvsVIeqdXYfl+5MzejQBaFDjFvGDSTMjUsoOSxTvndaUXBbs/xEG18
hw7KOt0M6vDdWpqJQsQ8/A4fEAOjNhMYVBFHqvB1TvRvkES1OSQ3512OKEQ9Cm2P
bvT697HZ6kIxEfCZSk+qrUTkQ1ync+T2xov2Dmhp9WfvWHUUOT+bnvyLxaggZ+Ne
AEXFJD9CQIYX3XQgsqwHpm28sFBYlE/rFe8b4xO/8VFrFr0DvcU4ZMz1uuw2JU6C
bMCrbKNy5JtMR2b9sch4oGiZlUmYst5X7I8cucUL6wN5enZ7N3wSPi4KU/vtfJZd
nCfTS+/Of+n3/zZXu066PoDfOssblUYWZOCaBsAw4J7UTRIW+jzoMPvl2uOSaRxd
6sFzsFiCNiyKOYeU38+htKKQacVMR2VIJJyHHy0nwNSacKLxZgzjPUa6SJy0bX8t
H9GmyskKYV2NIWipRyLkRQ8B98443BlwMg+HCpdLDl/HSZ/IzRO3i5mm7MvmS0q5
THLi2vyWG2rRUAiUe5ngf53onxL+xhFm9qxkE/4Z2d12DlL6I1fyevrGFUtFoHVi
VcwqWTS+Gc1MAx454agaVCLpNImAeq3TP5QPj+oH0QHV6JUm1sUHps6oboPZZnlj
6EqoaLLfDg9vi8dmsHc7HSOmsavcTQEysB3b3N1dD7j9VWjQoPfAOLaCi/xRm/Jy
7d9pt0KRZjs3REYNncQ4ukYj9YYi5EgmLfdVUYdh3u3Xv05g6rvzRlFavc+zR3Z6
uNckCya1oQXSQgAEqVOgcdrITgHPAEF06QohIIUcdwrG8/+vlLfhNBpfjvKNHHA6
OU+UtvfheB/WR1IVR3Ma5HfNo4fczHXw5j9/GKicKn+8XPlRjLtIVYfDxCZ5WNVk
YzCYjYchfq8EL0FWIn9GbtaTb33rsZyML2fsz5rSKTQ8/9AxjNkCfnVM3xay5g0C
YGMKi9jLZpQmrIpqxie10m4SZQiATc3+lNyQ1bu6bCi/5cglyRsi9+zDuN848L0w
IE+vyS+1MwRc7kpalWlS/PYv8O2fyaiLUJi92ikV3gTawENQaVmhqWDA5rc94nT/
a8jyxDu4riR/6OlkeR5ssfhmwVKRsqe200Tc35eiAMeC0ztNd0j1TuLNjSbx/YpF
Pp10GxRlNM7OGdBeZ3NhvU0gBoXR0vsaIS8YfN3wBTt8BS57rW3uPhf8AQt1x9q2
Bwivb2f+TZSdULt2zjMiIlQjUtTtX4ucPDCkmNqrZb7Rm9qDMwNnc14EKYtMSzXZ
MBZStxamTTs6GpjWEsaQ7myopSu5wRbLfMz146FcIPlO499WvbOXD/c6RvVrFV2k
dqfdU9HULD6lKjpA7yKaoaQneEjNqIyPR5rjmO9wftulN9HxyO3cKFF8S7Heyq5G
Rio/Z/ax/smqZaxNyz6d2LmpPeVJiPJNJb83ZqvGXlmFmiCZbL6zB4ThN8bIYwUD
Il6r1FAjretCUVR+QD/KRPsQc8r1FYxECaEZLQDg7SoXRM6A64n05xpjoFoQ1Xr+
uRBwVp7RcxzgWwQQKDBkM7BqT2XDD0Fi9xfQ3kUnE3vyMOVPRJYbqgt5IZYjuyRF
akfxAp9L6TCjNN3yOIjvMbhGTRq1PF71HPV0L831H8l64QSz/kGtx0uoGSJ8tTFW
BaM/u9VLBigIzoM0+9+JLe5b+yIc9CvMItAp8bJQFew+OREHtEyGY+MAgXOMAXUt
6Wp/6sVm+k52xwqKn1DLI+R2ZhSL44l92ovd70XIjICMjux6cxy7lYcYUN9NFdFr
2aDDJpIy9RQH1PVlsSwYAQy24CAPhxMCaksw+ap8y61oOOWJEUw35OSzd5OqYkvO
bd54hJoxBwOKNh3xuHF4ULFgn7VTBU2wHWTdDvNl/Tbf6kQ2lTlPQ/zrUev+4hXq
3vhCvzPw4FU0Ti9g35VPu7CoQYYJ7UAA62PdHkmO/Tx+/+tTYZkmnEbovDfYXf7p
zqWbgejv9w3tNQD7jkObadCIerBQ/bkHl7sGdqHXXUGuZONJgFmKU6/FFXlOIV7F
1brH2qa4o8W6hxgK+slfk9TKcke6UB4bzyonOAcRmQGxv3oBL/ed5Jn0oSf7VaWY
GGqgWNzObBwCvdBEjGSh9jF8KHTb8CUdEj/MjH2LXCAJ2qzjIUlNfVySKIyZtSBg
8aV1qg7jX3yR3lIbEbSE1iZeHMW6UWb4rCzE3BQ5l4S71LHiSvm5ySd4MKwLrkj0
6R9WD0rj/zs81br+MKzy6zE4B/l1Kp+SM60gwb61U8EqNr3NN/KLep2+HGn25sW8
8X00pQq6DwtJU6Z1/LCrgymFE8A+YCX3a82VK7jwi8VOxdqmF712JEkEub/Ydye7
AC/cWOLcI4vB2QFJO2m0YPwP01f3VlKQqsfe8hm4NWm7sSull952bCu+6cy5tizk
pKL86lkeocgmZP9iDIXJ0QpgbMsMdsWutVwY4sfzkCcPGC65pzSRVWHM0X/k7LtH
mA4cuLohSwv0q6Du+kr5ACU3xeBPLfx07FKthdpQR8RZjCA2l+JG4xCttZ5ljaor
Zhy4yj/JaWunuczhlYIPI4kb8nmM9LjqucQMuySQde6OhuBnoNvoEpXBlA2xobYm
dnGcgyXoiLcU9HdXyteIhWJ5ljBWW44D9Vjbs/CQ2gB8KMjvbsW5Q7dvJIU1TBuT
V+ovyvVtupeIYv36fuci+HFvfnMLyg+K4b0gtPI4M/HkYcSR1RUmL0u63JCxfEVi
GsQwte1ImL5kLWq9DDlGChJVf05NdOolEsNuvas0zkxSIG11qFH5wd9lQ1uAYutT
wBmSPlSPr2OB3Vn1tAkOzdy5yjdcg/bnHUVETHZ7d9nf1AFR+gZKPB4qhfIAE6AI
q5tI/xjX/xgAtDIOXBgjfGuMjKx+cyKzGRx6rYfwQNyJfZJun9pNzZ3r3bdMn/aM
6+LwXKMWyPKkbvFyJOLjASEAuyR+bnbKgvNpIcH0mHDH5jFs+EAimQUSGbKynll4
jniNgFpgtD3daPtUOaV6GOGSZC9MGuZmyejNCnr1ywArk1hSLQQTOXagDjfWw87n
jC/PaW4Zq+C2az22cke+0jxmd96VxS/CHalBtP4r9xsLMoSByp1yBh5UyhA/CdwY
j4n6GmWLWtK38re0Km/04sSWBQ+DpQJKXhT1XftR5paYO4FoRLT5U64ssiTGuGdl
woSlRLPiML1cF/KgYi49TmWjXvgLUHvLtAezdNjuMKqf5CmuDgrS1ZDErK1pouMi
vkAxTbjeQq0WDMOGp0IGwVSplByWD/FhmSJLGpaIypbKlp6tPm/QSHlKpCiP/Hw2
uirFZiBBtIMpk62Kz63d4YQUog2+ATuuCNI5Bm473YoOqKrGwrQal9HfYCBUpZLI
0/afJU24JHLg2F/Tr16TlHDRh6FkXhT09x6OAew1wqvSfQs5zA4X8j1qMSD1Q9Vf
/i5FhSDICdLMk8y2zbYIBqLlV9EPN7Ss4irU03VTDq2fAU+XFT7NRGJdslmhG7MB
r6TFuP7MCs8faClmcE5THCmAMF5y7yjVIqtGgEudUtKT25O9hrmlR9Z6dByhdsdb
XlM8dEwYbYiyLo1HWuzCU5/zRqPiVvdOHc0JI5n4p4kWMIIHZjsxeVQAICwn6PBd
BjBK6C4B6rcofT9i8h+ERadwcWkh6mxEp5bTlpJ9qeIMypvlI1lV2nTXRYS9Wt9H
wqmoKHKOzMgo2qGFXajvPAYXFX4ZAsbxEYy1OOgkkBDoA9pWU2sWkn+AY0BIX0G7
6rgLJCy+qE02WgelXuzzdh2mpk+9SsqxZeHFMAs6JNXSUMJeMJKMt1TsWePg7t5a
FzryR4ohTxECmpuT3c9Ie0QA5vMRaxWaPRypv1haqgph62AcQHJQMbNYT5M0gg7O
o4+uha6mce3wzpVdlqzJvPm7E6HXaSZknzzp2Q/K6wzzmvowaTWn4XbU1NIwW5i5
sJZSzIULn5IMzBZkdyR8AX1gmO1gnNKAupgS3+kS9UydGQZCqFy3iZx3fi7qt6eo
MX0bQqvbfc3nrlPFKwcyvO6tASrWZus8CU77G+MKsOj8KMfXHruw1+fMy0yuCjXj
DTsA1MFxabqDvJTv/jzlCLmVDj1DAm715DTGL3QFG1pS6kodmiXojjt884/Sw3AD
kYURuFK1/ArY9w1KxPlu0WYQ2WyKXDHWmhH8crEFLPfOAY/4wU1SI9uo3OSjdKdT
ZB/4GfL8D/1MJZ8ZaDOg6xzm2nLJNjThDGpwlj+a8puNzrXtvwRcq22BzF/q/bol
NycgdlG/WNVDLwCLFs8lId49JJlSBwhecsepNp7hPgBFH5+0DbgiGoH4ixq31Njh
04cAZ+Aq7e4+xH+9GepS+tyvpWBKdQNkXZ+gN6oyvrQ1nVURXXhcYWg+xg3JgnqE
ke4MOx3uBVU04jest2hhxXG90Dr6ctmfO8RH0qwRkJpX0f5NJkoBW4JcZgpWdiMa
qLmEQ+MD8y7lSebkgQY3FtP0Ir6+IX23Nf6SsIpWjoZG8ExOmWvlX2HEXZrJ9MxU
zIlyrp0Z3Uot9jCCjMjeCryfJErfrZmSIZd3maShQGoPlCMf2cB5HzPK5nOEBH8J
n3QNciGc+YA3vrkZbYPZ40e08LVoedOlEXnxWquDT637C0VbvCUq1a/4Re5W+kn0
ZxG+Mv8u+RnyXaJsCGyE13rJx4Fptb1cIVDywgx4lJ+FoP+CMUHbJl/W2eO37l7h
8MVhyE29ecQ2NIJv5bq+1a5vuUdXW8OxHQ4i4fcM3ZOVyjEfI44cFVMQeJOJZ3jX
oa6ehXxEPW45cHsau1gH6ZmCCRL9bcDNV8Ij3ikIuzwAqFjp1Irsj5vhhEPjT6ey
xVrelHvPy/l9OtdVBKpej/x/wVP/70uJmk1BBvJyJKFyj4HbeMl0YoGNO11j7rP5
u1F0sLKwqlg+noZ9oAAtCc3Cl/pV5aVcsjZCHaP+rFpPwbDb22WKlxuSOb2ZQpJM
i1FsmCyH6L/a898pOpqwsDS9tEIcTYLLEGAwvFpbsMyB4eZchdN2InZGywFZgM23
Zn8W93IGn5/H4ltAPFuoIQc8uugswJVls9vdEv6n3GodQkhM44EPkjhDc/hKHBN4
UfDAYXwxEYG9N+KOJUCSJW/i7D5otAXgghmpdEXqCl7fEFSXl9w8cPU/5eNSajPb
dKNMvWBcaAMIJpW3OiPqEPNUjSlAPiLzwtuajsqWU9FzTMknqlXDDWlhv3ptLoxv
EBwMFV3344vcApeZjG3BabQgrd8tyx0QxCuNSFIKemLmZpqZMxK68zvf0EIEtBOj
ueVVdfTdRa5/45ypROQUfrPdpYaveNgjP9V+S+bgsOFBy23prsxIVHM2HyBKN5hp
0+M5BJOl3poeB5M4e4G8BEp/rPnXhPcox3wNU3Har0uYBy/AZ/mb8op2J0+qwpUn
3AHFMy1ZUnjpRE9sf3ajku97KVVca9+71+HqUlxJFKxz1H6KSbFd0ynUjNfeSWiN
bzBo1r6/D5XdDGrRhOHKK6d0S4A1tOeOi3J9xiqf1VcdmKQfjH+Ahxt2yyFRiFrM
jUOEguAgvCxbxnhyaDYdDBiGBwuufeI3y+Gqfu0TrQI3bkBT6TC1peGWDzn6/iwl
++skUfNt6YjmcZA0RxHbv40VuOz1Y8jpkB/Qu4xXoUBrxRWlHGbM7VqLV51hG8+h
o55vLAxrVWB+Vuohe+fIA9Vi1vRHQsDQJVh1SLWdntdR0LB71h8vKtekTIWZfM/J
nKyHBS7vmOxejEwHV98SN0CMfX9Be2WMmTkXrwsPsqJwxj/lcJPMMqgNWlvI6818
pDt7GygVAupGVeeyhoQdsJwzKPhYSKis55DVnbXZVsS1pqLlXOfRyrI25bkXbCuc
yoP4lhEzj/gZ9QPIDxtWqf6RzUK6CwOdifkCN7tSRMD1zpKYbIa0bjzEcItH20ep
ReNEwUkQ19yCy6EvA8lnBebF4qIm3jwDkUxKlUNvOkh4ww2KC7x1WZxVlp115/c5
mRZwtnsVdCBYwm+wKMDg7Gt13PFhoehR2n5lwFM3im4j+SW0l53yejzThbin4ikH
IXOeSm5RmXksrtQFicr/egcmOdKBE8gYtE6BHl8VDayFhYYWYVDe+DdwNSUpnpqk
2wDkY9vJlNGhoW05xK9Ko/NeFAMTa93PY1alguf5LbTUJEqukE6BYpdQy6sefhYj
AW0mrj6YfJFeHmaeXL5K052Ol0UK929/4M4M/OKO6NNKiHj19fV1fVRY8lUzCgap
N98U3SXSJyh/52Gue5j3NBH6ty1ukbaMCiOsLFEsmtNVSKQZroBkuJxUHwOSPTbG
IdnZvL1Nkw4UG1USX5MnTZ0JXwc5oOUVTIzfGON3b4rkX8r2F8AzjSFx1rFGlJiy
uiS+/ly75Nj3QAl8nSVVwXAwh6sKGhhNJFRG3oNzsPEto45fWC39A3nDKzFyo4S5
Rp6yICopNngup01gVG0N9B4QvtZG+AmDMD3KBl+wW1x1myVO8FUyHIQd+4UzJpYm
VTAEbLkDqWJVm5gq/cN/3Cpo3OHy2G57sF4igigEK3otYjSWeiTuIH8XNxWfc56X
3vuMxM4e6RgIWjXJWjYUWON9nEec2wm9MqKWqSTMOA1rwrtlyum6yBg7AKAhwfz2
59vzxcGinHvMk+TTqdGjbguyY4+2/59uKIqTl4tFr9oOPNdy0dNohFvpNBRCTwKr
hjg+xrWih+VtgP/xa5JhSAI9zkm3/zi76qizksQ2GBwXbX8D0xeRbBVjP1r3TvzG
gFgwfWMuOwfPr8yqqYODR6lOqYF+jhlJwo7CK+wQqpuw7KApKt9dMrjt50JJHPes
nqREA5mlm5ikx6LDVSoMFLB/5ncEW/fuhAvo/txkU5nprHOXSWzXLdYLZc6axXli
9d2TQ95ogMY6962iqfGgm/H1z5QkGyrUjR4/ihPpzVX502N005Y2+ApPSW8pSCPR
DmiZ/B4op2uEYF1/TfwEA2/k42BaxMlPJaQXiUHWkzJgdcuLsjd3VAu3aLzieSb1
VT9By2fm9XHtVWujXcEAuGSVMdIHOcCJKt6zrWpb8RtAaWw8D1l5MckFtImVIZlx
7vri/qAiD1hCL1TbVTqEM5Xk9UMp8SdUBa8n6t8oBjwXvYLarAPNNRVdB18WiT4H
t+L3mLZnOA37UJ8G3R3Ljqu/+GWDhVY6WH3vLtY/V5Ks20HKG89QmICAVWxAZqB7
p4HHmn1e1L5ro5Fu206pl23/FezUvPhq4OIG04PztdZLdUCHVDdYaU4qsms423/9
tGe4ds9cejZnqLgpCArFdz51+0nwAVHTiVuvEh2nfqhlr7jhKRMpRo5myeAgsQEb
J5Sdich9KDQlDAUiz/nZONRZEohWvULVB7IuSAqhb1HoewqDv4gcPAKXk9ja/k3C
hKYKsZCWCDtBHfrDf0K6OSnsVcTu8OEOC0tVKB/z94lI+jkAS+gZIWeqUtJCL88L
t5k3v/O3RxbuSDL70Ro9zyUckw+ssCtwsd5RibPS8xyvYdT9YRGOg+ZTTQk7dKW5
9dsIgm+9qWCCJsi613EBfq/Y4LDPabCUT10El9O6REzVltgbI6mdISxWJ8GA/HmG
ZkK+jI/DQKlh9EQBhWinx83Re6HI9TW8IJi+E8gH9agegYHZ503WS+oo+JrAqY9K
A7P6JCPAobVfIxhjNLDOjLuYmtu213N2EH3dofckd89Rzi4dPl1cFZ7AwlMg/Wab
27M11D+Vfu9GWDsNr2cTuj7przupxtDc3u1BgTdihEHRRPAeakxi+OYIStNNQopS
eIlbKWAWBmbQ4mFSv46OZlZWjirNagE7PLX8olACINgbBOBtkeAlrQd/ISAmPUnr
oXP1EwVhplfhEYOq3LSpNK4+4DjMQ4uvfhRSq9XqQeqG1780KkZUCRg1xsaSSwse
54N6qjCf6CZDssgISupi8KEY16JEbpmR3CRKDgFjmQymjn1t677FxsUOEsqPFs0N
DVnu0+f9cV56a+65s+aZkuK3ru0rBa2w3ksOiFuKQy3F6opd43EuNw5GJDgI+I21
vtQrP1BlSWCS5kQu9dEWiFS61FcDDbGEviI6zVjeSM3XkA3SDJPA9GlfoEmWhpUs
BAb9UYtvpQB25VzKU9smxu6UG76NyZN76vJ+ltopvUCdO1eYR2uxXc1HsqLNDXQG
5LuIIj/5NBWZE+/kPCWrmWLsFMIkVia4YEPi5kRpYJL7BOjKrfxo7+CUzCbel7f2
gUwEe5pSfgr8ON0Efpi1dhiyj1VCK9rLRzDXpCGrH00T2vtpA3Z4Dy9D5vU2mWqh
18Nn45fEih0bzeoFxhxLLXVMDNeEayg/F63g4HvLFeDPbUidE66gsyyb8+gsULuf
1NH1Il6FfFssoU8PrzCJCmIukgomr7fAZpmjlAqalaTpRWqipDZpqhZ7tdcaKXSK
8K5y/Kk8OFP/+72+JqouSZJds2zBA/yFt60OIp5ba11dR/VbkwzeiYUH0UuaNby7
QAgJClvPdE6Z9IOIiM7w7RtirLh4nxuO6R6YNk18SOdtlDYVz/F2+9+N1hcnCmCx
08yYbQ4bBgrw5VhpXVe/e6LCJlXhSRQOcMa/v3bvL0ua7llP+tFrqXMQRJ9rnVbZ
/dMwWtcpW3LetYuimRmNWExnapFOZmc+6UFT3RaI1Gxgcgtbbq+TaqVmcSE/0eFE
d6j8d3QojCGXxEwrKtAvZ/OBXqoHaA8IYPH3LqqaX+RL5gK2LmMiC8LLMFLS6ynU
8x/tQv60hJKKvrwHcum/z6B+xjkAy0o9GODS6t2c5ibiXm714Ra9J30TGGwxnCEg
4jcObG6yEmwDFJ0rzq/pKJ7KFLqQdi5Dq1HsGQxaszOulvm0oRKak+Bqtw+ErNsw
KAbBzhyih77GHsTMQENq/h1yNP8HCpMVxDtqCqDE84NbmQbeJoH2thnFyL5lqrF+
R6c4elLXjPbxbKk3+vrtBV5a6IXvtyuOvzSYn7q8K1JhiVpFcboBMGZ7OUsXv2mk
0bOuonx2SrII7k6RV5Ad+t7/8GByt+ap6HVxIt7tCGNbolAWLFhGu5ozZxqxr5uO
nHKcvbpmXdP/XL1y8CC9i0x7s1wbuo+/Nl0TafISABxg3LVksapc4aCxAAxVCdjR
IeGL11JqKx4As0gNIQbmsf7Hr4bmU19qTJFvgPulOmdPtSg29nkDQhUYXt36GGcM
Y8dkfIIILTiJW3/H6anx6Izxiiigso0UsFj+UxkpLpWXX+W4EkOqTC6ekGl5WfwI
aJtNG0S91lwOZJliBcDU6/ejbTeEvoQAgevzgtxylu4jrNrPfpZDu9dodw07mu2G
+mlgC9cxUk9N+VJvGiwhBO41ACiTH9Nf9uIR6T4H/hv7LZtgjnW2RgJYCti+Z+c1
rZ+k/9CNXGT1VcVDNyHFRU79rrGMtcyKuodHASYv72lwGYe1S9m3Or9Z9P2A9/2w
sG+aPmLNh1WkowrJI05JSfLkluZPH+MRdP7WgK5JKIwsKBV0SwrREBgNPOaUvM+o
RHQ3Qkn598dEqtPo4udZUmCbINmGVvlPFJ9Im/MMBdO5Lvfnx38Qk3j/ygojoJxi
v5OnjvkQwksgvAD87zkhDq4mSFI4NN18JA5OiCSDNVfbAVJMuV14BPtaNNnV2N/F
c5ZmHQvma32X3Fpvpfu/mR6Gxs2iQjy0kgkzKpa4j+l6nyGYXhALh8KaqCV/rykR
Rd44O4os/7FMTuSeB4i1c9vDWNI635k6UXocdVDoBfQf43MznFIeSWFG3rZO3G9Z
jq3Pr9ExU/jMZXfwJJqdriiifgRLulS4tp2BesgIJN/2LB1yRuSXD/HlEE3UMRqb
bNXtIssKPBimnW/YimE/9ArTrhhZXaruL8wAmiINQRDZtsLe3cEjRX0cNz//uh3t
QsgMGpoojZxgW5PChMJ1ufjC75qunmLeFJmCJ14SOvxoI697FMqlhWLKRLy5fvnO
WU+eL62/w65BcW5w48KjGin7DU78ShsSwy3nu9fsS5qAk8lQbW1txmkzrK/LOog5
rTAKkvKhnwJwsThRkN2SSA7NkhNgBC3v7tBovJqaDyLaMesbPkP0xNlCcTr13xKT
I11SamqlzoUvYJsuzmg6yWvLwOzIEcTdhsnbdRn5TQsZPkAkMJcHSZpwE0lrBN/B
t1EXZ3yCdXB5qkLBSQmG5DTbpugfjtJtQN2mKCrO/T42iDpcIHPQMoI00s4d1t3a
X7dh1SGR7tYiqEvOFhikSLxosRO9uQe0PMxUbUq94tJfZ4vEjnqwuMpdi9eiCNqM
8baUbP/VcYPMSVWokI3Im4cYVOJUKrZoYwLycgv2w9ELOWKqw+RZ+8qPctg59WkF
cKxJniI7Q7xbaBxEiR1VkHLcUXiFUID91NCC7WV9hRW4ZvPkAe7PvsjmnMVDTqgb
B+qh7ObHqtvn7MjbnCnx1FDIAmY5fSFy+JXlyo32jP/ipUBKsWx9UBndGE9t3wXA
YFKaH8HYgh/O8r8LO1i6Wfvrs4AHOt8FHmASyHNwqn3FoO+SBL7XRgckCpvw0Jjm
fdlpnv6cmn0DPw0d+olOoHKDqnoQAA7Mqx4o0Tf8qKO5/P/E0sxTnRkICLuT5sgR
oggQsskaQ1vZRKOrgEpLZnQJdE1zRxyzja5u/K479izJaiW54BJ9E+YcyIF0QdNn
BwfvLjww+6l/DAXsANazBGBlOIPAMSbd9/UgGEpUcz86U1wNInthSGQe7qf4A+7U
qvNxG/jCW7Y27dK7tYwPzQ8joJbcE30nS/bAXL/XVvhhKGsARSLBqrZFVAhB/9/T
ORFc8TAbmp//ApsyPKJtoxb/pO4bQfq3zYN7NZGGmLmC58O05uomqB/TliBCC4cK
Q9GFqfIn06cmE0SAbsmBnDRiJGMEeK3X8AcmAewguqP9ojaQuljQBPS015j5SoHq
aW60K5UqJRfTz5q6CH1GK2Wjh/M0I5Wsrk4kBeryvoBfC1/ebjKXULhTdtu4fm1k
XJ/Q9zqE+P8NrShm0axYfrBHOYTrDvPO0SEEBZn2LP2j+vv/SFcn2quuZqpo+M/7
Jj6OZ0aB2yRp8548TuM4DuYHzI5C7JpGsJA+OaKiApP6QlMAJhB8wohujNisP74K
oo+lRoRLWUfMqo772QagcMLlnAxNDqfGIULI7MInammhgsx0kVtgTh9QkP+1xUE2
E8AUulZ3Zr5SmKYl7hPGUvxtDo7KriLzzmf6637Edh/2FaNgPzj/EgQfKzTsHrqj
tAlRMpFtoVYl5Qd1ZIJoJsjqfKfl4oAWKdRbfExZMMJtxoq2R5NJILB/Cgj6KWHW
IZUPBXajw8G4CjH8V+rZwqu+5ncEuPbWgAHEMITZ3sKOnu8Vn+ci7w6h5/s6KGgQ
NVlC/nikSi9+YQp52Cv392PbLo0imGDAV71PZRyLQPXdnvAONzA92POQGs0AF6Jv
V9G/ySJ15muVSZlaUXEZx7pjyT+8IXYSux93S+wvuvCktXyai1eIQMT0ZBOEpiql
8w/L2coYo5yWACxNl0oxqELHuXq6jrSD3RfIwVK+wW4Gz6H680lYOpJVkPtG/uMz
8mYkhl/WBcK9/5PgsxFPJ12F337V7rvAX5czuWsTgr25aGK5BOoBQYBoQSgmlV7i
6Gv8aAnWHjkcED3Hjbs0Lud9syG9LifNftnRHmXfbvF30nvT1DXyysgi6pKENHUI
+FgOMKdZkWHbHZE2R8h1RNpKrCtKZpEV73TxhIk+iDJHE29MWLm1HTICHPJVunR+
Aja/anOtHyGl0eDMdWOqapI4+MypF4Kr3CneE9vXWuYvtDVR6WsZwsYN5ikNofB0
Tb7DzVX+QYL45uZ116/sj/l38XMqCp/mrHO4UP9oS/2RogH8WVki3Q8PxbYqnMVY
uOrHKfas21ngSvpHfn03LtHfcFy7bxu9GnXBGgsgF5aN0ZGGZJacojg7FeDG+3BZ
EjvHUcEN05qk+3JboI8dBYTIlbmyvK7NIJoNprm0B3JNx2V7dk+WqFKMwV3yVyM+
A8VWDHqUjZY48LYbUHrHsPPxvM2OJljhz5gpRESIUZUSIoBh+8JVzeyKiEBFw26Z
TD2swZ4FcZCGfUqcB1nW/E/O4GopheOYYi7OR+r5J4QXuTRg+qS/73pz78tpat3A
yrigsFXny6XjoHU/5mZZicbGvaIqJgsRd7lvpbA13wuEjbmC7uitzpGkgS15R9s+
NDhkxjYjA820kJ9Fi7qkigR5mrnBfJkkTM6N59QoXFKXk1ZVxn7BtaPDgnTLuhIt
atrcz6BDgOWtL7uNh1NVsR5yjzIBjCYF4LJ6EcPt/EcesoznjRTjY97UkRXfGc4k
rlppTvGC93y3YRVyo9+Z0qc3dfA9d0HmjFoYksda5NaW5iZvB3JbRwqd6Fz+pVCu
B1lmp+4vxDjAD7GnI00Uhl7zMfN6hDNeN2Q8W+qtQueMXJ8HTNU9GU/Xzi16LoxT
naP9jjJ5GXFtCEwNYhzqfYCDeTOEJIb0Xje0Ivfw9N+uXqowxv7gv/Z14zUKeoTP
7q/XMODMwV9flT/sqaXshADTLIKmpmJcws8Yxn3WICQ4Lv5QDELqY02T6umOH4Be
ZfLJ+xiemSJYnblxYjHsUe5/gp/2biwEdpbJxPqjcNN7fNuYPotmAGzWue5MZpKk
muI7qovpEspcbdkDoAUztEPwQZOyWGVIXCCWlTxJ5WWwf0+B6gBlie098Fdnc2FG
6Cx0ygigQDDR9p4kZGJbl1Mau0q30jAIhwqjoziZsgttJnjtLwhtBhnE4GcqeLap
dhuVRuLmV1JSwK6fNDYlBoqD7a11i4ulCMj+2rrAFwRSsZlcqB9YWi8v7mClNW4o
flP6svmiIxw2ZY53bo4iizwhNYWKSjljzmxY9ekvKnekejSyfHnJKtaksq20eb+Y
+jnSWuETem0+Ho9rBOtJW/N9qTqUagj5uudWQC/YPAWF+g+KyGIcFPgqXanRYGNp
qqmtfmY5Gnn9E8DdNHIDnkIYgaOOb57B8UXoNZo8tvDrsh+Fx1+g1iWoRO8cNgXo
0o9OkNYW06ZY+sslnYUCOGamSzPW5TXvK0f0+rPNbyzeCYR2gajGNyoWseKBAyDn
hYMDn5I/+/BZp3CYAjC6OOIbZZpC0Y+VdmTcUXebHI93RHufvwxUWpFNTmq1iT8t
8HrQpg+OnsmX0j3vCAUlTCUDJ0kZVRH4HiMRkSclQ+f2hJhOjOogiGfvrUKIwGAE
p+Gw7AKLmQHhRDHCJTV2vLE7Gfk5FD2Ay3XlGl6nsnx43aGaQ4c0RjPQ72VU9/62
wxQhbj0h4DEWxsrepJ3I7Bq2+tJkNyD7JSs9Y79eFpOxyUp3W00+lcHOlV9e2hMz
f6+6m8sgoWvCvzh9iVO1d7w3hJz9deQk8doXXFIT4Ecc+Q3NqBYcDMx46ocdjou2
gG5zzndV2RCm75NeLekxWM8TotzNJdUYDnKxmHq0oXBrp+1qx3GSoGZ+5JjKpQL5
sHaDe/LNTn3JnKkgeiz0eOnIr6h9tNIW7dC2T9X74QA/VEXLAntFWQkSHBV3n5uU
6Ff2N19v53DaI/4gCSW6d+O/Se/Q+GdM3LLzrLBZwZHiUtQipx50fGxFmeac9bhp
Mk/BaGPH2VACUgLQxVJL8aSgdxXj9LqdNav14Ih/SGlZ5C555851ZICg+Xl4kIMi
XF5Y/I64TobtP9P8fycacS9EC6AyhIqpT6o42atZDgZw9vuZR9XDYvDpbj8I6eNS
tQa9wMs45ihHM6yDYgSRcqOA/KFRBo6fpVCYMIZGqWtIz+QDFN49k8zXyb5dQd84
o/51b0hOxt6pQGAkeQWcqC3pkRiEWJg7TqGLpxeL+uw8hZzeTzb3zBSZcmReqS+7
c3XN/Yu3XvCRkVCRfThY3pCFxOoCjtENtGIn1nNPXxUMNbWcueM+vjTfc16wREpn
6lxczGeKd0TZ/MwR98zcEmsI5BiD/4oDbUl7c1mupe8nA67PAc7tgTyh86kllDUG
LMayWe7B67i8LCuSjon9qryNVql9bd7wF1P5UvdZsu+1PAfd751M/4bto0oLPVey
WmJREMT7+dgiGc8QRVOGB9GQ8rvKXr2Pewnygutqea8jzL74rpLbM7NK78VaWDTS
9o8HNcIVL2PP8MnB0xAbBGfi0XEmee64egsq7VlCTw+27sZGT9WAfmSEnZFzItXw
XgtLNz5aPomBSFxi8iVpE6tumzXIsjp30vSoO3Rz5JSoiHraTi3eovI7B6xN+tpN
8L9o+S/hPLJiXiXtqXqKTrkUf9vbh967TJQHaHuKA932/Wi1J+IySqzBAhRML/bh
kTxPAD00DeIYf0nxAmpt0lhLp2+kwtMv5820rEe7th4nBOZ3vl8rB7I5ZEkA95FG
bID3JRBD1s+AdFpLi3Vdh0aN2oWrrj9ANPHRGC6vQfC6RqSuUFHdgL2mHtwklwN7
dxF1oJ3kVhrGYDdZoHfdqNLEN+KXo+tpVOXnSjv2LOW7mTymNVogv4KwMqBdnGRr
8HmGcaE+ThFjF9O6rBdx9JD5Bd9deFdtcsmO1WhZfCFdcJkFOdP+yVet6T+PMiSv
Djax0y7fKKKAB13bK89/PmS7tY5plu9AaV1nRNGgaXjF/wACgHGbJbiMsX4IkgYA
oWfDPBoGV798u5+qPE2PYSPjlyvCx7OB7Fq68xAr/e48VolCDy0cSqRpyzG3tpRI
41Yckl54G4vzYnscH1U2SD/Or1V5KC0/KCtnak+T/gyr0u6HVhkYEmqgjyjeZlaD
jxb0+Sac3ICYYTufKoufsTeL1+E/jZKg+XnHLxamGyg79yajIpGDR7jFqPyhQChz
puRuE4PskLV5lHoJitQOdoxNxeYSdBpMG+oLNTkgB3onoI8m9kLARMslxZ9CSmMh
hWoMsp3dVLrz4wB1WTrBWv9Z4F+tQLL3eGm9RwE+YFofyxVf9nNx5Cz6HhtAUYI0
1xlxK2qh7JNUZ5smUJ2XeZyggpPqgE2TvBgPK0tZACEopje56PLGEtoxL/vE+ACu
sXhy9G8OIxw9tKHANCgJqNOFHtj60iz0Oi+tKbLkO24+Z8XXEmMpClZK8/53cqsb
hS7lDru8Qs+uEHmAwtCpfPYio+bREhR1C4UO0BnAv7JGIvECZhxDqnCynCYGSJWO
QHPNtYss+2iOQF0uQgJxv6zKJL6946SAFuhmRsu4qrtDNRxvkUFSMLY9E43Exqv5
qjxSBY8bv+Pg0YqBlW3tgEf6Yzr2OY7LqwLhxpyMmT5fyeRqEJOniFA0YqrysaJY
e2R7ZeCMTl3zh4XR0nhg7k2jZ/yvFviKvo22K/Jpf5utcoiC4e8CE+Ee6mnINDyw
W0CrHALZ9j+tB2gOVJ9OnLSQItnXz/PHwNlqEKMijyo9AsAxjglxXaK2usQcuNbA
8AXR7ystU6oZaPMKhuSqi/VQ3wvSAYihUwqKWkvn8s3hsf57XaomWKQnsluEEMtH
67poaN59dCt4rzY9rRolRBJBhpxBwQUrVQmlIIGskSPpCnZ1K6t6TODNM7mV/V5j
IPKnziCz9q5XzQ8gfjJiZl/soJgEzL1wmrvfOS4ayXlXkZu/0EGriH1FCH6WPk4j
0443zt8JgN0dyU55A96DxKlC19UntklUqqtLYHJeTkiQB4VMZc5LMQN//yazeoeI
iFIeoEeTZbb2Feo5HkAzxFehWK1nnAbYERuDWpIqnqpvfsKLwsp/hxO50hIZZoqi
uxdQNHu5SElSUuRO6lo3vHJndVClOnSl3SEfyWY432NXTRZL/z/S6pKrCfsyE/1d
bHN5TVzYrNdaUb9BXow7h7G17U7F5CM5BQtSCEWQKa1X3hkmrEBUWFT1PL8N+/nY
Fj3DWecChwNBVHLhKm0Gn8buW6uh6tZWw4V9nUG993iqlq74kSXk8yk986RDp+wD
Yy2ZShH4a63OZiTrviQySGmou0GCbHScC7GrJ/bZtM2UrZjNnVi7GqAyn1QyDac2
1ZRLurxcSxU8LDjKHjf78ha3h6qc3m6LhNOpVXWuwFmflm9z3oTztBWINP6TCnW4
03MfNmGETJhnWK0uoVLqjA35p7ZU/LYu88Hn5MSzo7HBXleL0fXXVRIBy8Wo5HL+
F1+2V72d/Z2PiFTFrJ1VkLVWKd9s5AT655KRY7nJrsuCDhJDn7Ygw9sTfMoc5haM
pROqq0CH+mOUc0+gRWOiTx5wNjprVfZrOQc+QTbEuukwAfiuaxNS26itJA6oXlk/
8wz5sxgvUyyJDZtaPq+GT8nLKu1g6IAMghpefbTGj2MQXQAD3zYQiWWGKT1Ylh9r
It7AcKNMZ0F3GbwA22rZYEqW2mcE41pOaru7Juzj8haGr34Qt49SoM5kSANGgR9B
yqx9x5gY3ydzXh20yh9LNFrIMDISChF+9moTH39fd2KSlcbtMuny4WLt32Wf1dg5
oaRXI/cDXmdNhh4DWfCw4IBnOnU9JZ6eaJejK0IlKcJOAV2WT/H7n0u46G9ctj3A
ydkCd5nQmnN4BjZmptQyhFOB3CBsSAfzeRO3e0JVdXrfEttFgILBD/ERLb7heHA7
yJM9ys/Qi/0g1oktNGzlJKg9zd6hZ4ikTCJOu5vb3XMwaGV6ZrE9iYADbyuf3MEs
AOlnTQx8aUq0Ah275KJcDLBsGY5QACF9mq43xBsv6DVyNvTExQJauwI8A/9fgd0j
SmiQcRX4WTHBHDval8OgJnqqhr1TnbW6cDC2fJ8jAnSXxJ0zC2239OA0d81LsASS
xSFLY2CLmwpj66ySZsr1oDLFt+DRvQvNJFN7LWkdcOt+LeoNW5VgW8E8w8Udux/a
i9Hiq6EdT2pl0ywg+PgHsLv3uk1fwSwBF5BUuTT+EUUJd40IORTltnILK3plp6U/
ws+e6PUaTH+besC9c6fPJ4UUjrIerbMvFmJvQWVywngzrZFcvmmpMnZFBdWoFn9+
oWNCSq5elh/m5eXE42CL3zgoXsuFZugYpXB4cUknDe/S4Lh6mDjpnXy65sxX3kGs
1aegi2pP0SfnysSFx0ttEBIMrsb3BlEHhjTq8F5HfKLpeMiR3VQZz1hwUyeVo+rS
RGCDl822LcmwMMRabRdZKDnrxFzgoiOrvQmRv9bs4tyjtb7JXVMItGzjzI9w2HUG
Bcft4tYaBj9BRCMDh7AibKG4IyqKdaf6IltoGeu0kGV3tX3diGLZReSmKCYX6i9d
OAvEjs4V5ltQ7MsvYBmWdywPOLOK5cQdM1hPBHnQOVewawAZlh8ouCWCwEEPJdkP
5lW7GPytrUdgW0tSlW427YQS9yN0EIpPnBO+SuVXgf71BVBJkjHGtNDaYACyTBV0
UiBR0csJVYdiA6QR/8BxslLlekfKSBCPt8ejwHwTOTGqjCLxiOUoFpL2EFHAMCQj
Laogz7pR59ZKcb1u2D+njb3pJ9Eecuay00h0QPfiD5BSozCeRxNbuXRhUBMNs8oQ
Yt9r1OIsYaZ8g4oG1N51jfCc85ircQJZUBsgszqKoekcaozU6bo1QO81X/R4xvHK
gVHIS81zyC8ce33pRx/VqeaLIpBh2s2/FcptRBLmLSi1BlMtgU17XYfGO3hFYaLf
+9CymRMgITzH6Nm1ePFXbC7L+HOSp5vYgxIHtPjpOuJVuqGaq4KLQCztsPnzAvQS
VWKhL4U+JlatipzN4tCPHYGgm+eJoNPYXn/xbyBPdIekgJBeSuNGx8fx80noO8u4
mvQlphsMTLCW4xBa9AKzEC/HQ3VREAyupSq7+K9AimAr0gb0sOKp1jd5EV0PmldS
chIFLVHx7ZzZ18wXGffOjjoUIe8pVGaOaBp9yUEZmVn42TL/4TtM3rZWGRRXfNuM
IyBimIt3aEfMbgm2cPDn9155kHN6wYly5WqdOpIg9DIK5F3CLke7h2MsdrcpGuvP
naK38gQj829ZO7f3AAiaUI6gaDt7md9tVaUbsuE9bhQU0chlzT4Xc1rhr4Vz/rWt
irV8liwr6qsiQ3cv5uE50nbUZcAJCTp4YTgMVlGZZWK1+TwGqSK96n08JX1etmkg
4JiYelfZ2lKkBN638Zs7EWlTvM8cdxfbaNaKpNQt9gnz7cBDw726TIgzoxQ+ncPV
7WVD+HKh3iUjctUpOE4mNEhbrdbk8dEREkbbNJzXmFhUAi52qAX+yvbIzDONOAzA
Bd2kN2c5ynHkuAY9XYmpdhpxsougvKItIgzWLIHkNQii+9d3p47ucXhLGHW9LEgt
Jiqb1+mqFV1QdUArZRJjYiKyTmNYejUdWC+GxhJBhtCaAZlbpdD/qUlJS8du4w3C
E56mYLcRFdWiiTrfOH8wiQXSXx196ZxR/0MPTaFwovlj7Rl/tm/Tbwni2CjcKUqc
BaaFxlwKVVwimV7+ViGMpQjBIzBvFhRsysZkAf2VBr4R6s7U8qSVwS6jO8ue6+AZ
/uG0tFn1Ds/DO9n8ucnt9lYsGpTSm9LzQljtRN1p6NB606tjm64rX1Xb24/6Csqr
g33OFc4cLKP5KvBGRLAJyQGB/0w2kzvpCrZr5DF8sScI5ptByY0VEPmpOZoTT9mK
5eC1OGDaFTh3yYQ/tFHVSnndrK9pCa1A8+8Tr9UlrNJb6sx7xh7LeOUlZW96pMr4
t3JqJV5JPAb1CK+H/OZVEFLrbCFi/z9Qf1oe2AeESOG0P2sQokipGPJdeS2L+K7A
Wlw2ncpIl8BEssntobjIlHNiRmnn03ozwpRgMrfl1M7LJK7/YF4+h5ZJLrkBD3vE
ROcuaSq1+bc21P/i4IxpZZzScK8r5myLeU3GwdT36mOP3pytkwv9Uj7y0QzEFhZE
0DuuTlkNQkB5G+6+0ckzuAw5a38iiv6AWgG28ESdJAtUjblvQt8AnjKrmA6i+aLx
tVuPnPaVKrl1L/+VPVeHeOdT1ejRsjyV7L23yEhbbNIJIhE/iXeo2T63D7JLJCzs
6S2yFGYpFQarhIovTqFc+DNI5sBjYBEUdovScwapFda1ZZbwLiQ0nZbi1GfQFeyT
MlQ4VYRCBUsO4Sv7J0jFn7U6zO4TN77uLZPz79P3NRTGbjJkLTmsdmSWGDdIhuDm
JXpot8tX4T6OA1NgxDKilNu20dTR9LYQZAR/PhoUsU+pTeunTzA7MZDVUZfopnan
4iPgPixwOhP+NkkJg1GWrh5IklWXRHmTLp+cIyoYlfSOmLkEPPkhrQDnjIJcFO4j
PMPLlzl/xDKaB+i2TKkRtTqfD+UlWhU2wjPf/AbkjBCrQwIPEOepq1wAp+u5eyv+
q48GoXvufzAeXEnCh9hT2JIVQDm0nhhgnh4fZOEy4xHw4aWg0t5rOv7gcPLj3r/A
Nl32TPMttgBixJ4bRNmJqIGQpPqy9cZteVikb5ZyGPp6bcin4AIAIoADNEcR/e7s
XXrmQpmoCw0tEVYhbsACu07p/8Esy1Z9jxv8TEuxmB59iOFIVVXCSoycdpa0taC4
6avJGaffKK5NqC8QX3Er7rXhWbwnrTDHQ3EsBouBu+waydrC7OxJEsx54RPXfz8v
bHPyFSii8BteGoWz9nF29N5kutCy5arb3tMfngK80enkp0wceKiQRBol4tfa6fUO
Qwr8gdcLoiNZlYo+YxCPnTpxOYuLn3v97SYT5DCg5R8GQqgvFDGivJA77i8WjkuK
8erQgOPRUYrGV9WAvgo2GQTNXOywfGP2lfJyGxXe6Ng=
`protect END_PROTECTED
