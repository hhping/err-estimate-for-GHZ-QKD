`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YzNue7ClrsInFIJB5HItGLpDICjVUJaQK/Hl16Nei2sYTL3YggTvGpY6nbXG3muC
W5A3WgYBz2sfEaanZhz7Vn9Dx8lk6574ggjWJeOH12WdtHbg0fmFwnLqXS6+ulQG
iuby+tqwdJDUIjbwSshjJHIDyr+PgrOvBzLh4+GSAFQZLx7+7prvpboUCPW+Ltmf
Z71YAYpAD1fY9Hb/tNd/5rncrjzRLAnMlApLnFAGnM6uTvHGb/vQ0ReuKblDYNKo
3fMadNlJ/i05hmpriV+DlUvN7aw5VK6rCBIvLKDNytCGOwruxnoQ2CFa3jARUK2j
mCszfmAravPGrIvcd/dg/ZDBJmKYz0qse1/+cD0TFVFB8zxopi1/sM7c2nZD41DR
r+DyemORxqrcfQRK59c7MzDHHJY4outpjVWzJoBY1eNCv5XgMP9aZPCs8p68WyXT
e0u8y764sL8jP9eRA1fbD4OrHdD+V92s28ljv+LwWaV6j2MTh68sVxoEF91dsL6Y
tY4i5CvSNNvKH4oUJ4R0rb0UB++v7Ihn6fKpzR8ggSlqsFaJfHZkbYLOdgxT+uIM
`protect END_PROTECTED
