`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhBAiXNv+i/7BRO+3dyCtq1H4y+yHQdMbzcztbOJAkWNX9oHT8fpDPDVP2TaakEF
+4vRPic93lwPVLCk4Q2kuGvYLPj9fgcy6AfYGjPuDOr+2sEkW0b8DmP4F0PjYc7f
CekINzto8RDIfcIgE/G/9XHk6blgmw/ijD+9fcgZiHdnFFCVmpc+vtSpa/GUz9oV
33GQbc57/AeB6z0tkdwb2Vuqx7t9d46gYmv4xf5ZmELj7qNt18h3DH1WEUqa1vDs
aAo/f/QsDXXCutX4FQe+bpIzc8eg7KmdjYmM6+3EPWHIzTLf3nX0EYoiiW3Dvnng
HXNCjtXVYu5I8aZEcC5/l5IfWBDWlj32r8qFZEAqCvBJ7To74DbOF4U2wPqDsAdo
mt3iPTKO2K9nzEWFkYU6vv2InF9KLFYB/ku1PV2lm/IZ41T1edr4YVqIrJx+d5Ad
NUZcHWUDfmBeTlMbVKKQKCQCHXCjVSp7lEzh5jCXskWVEQ7hY7vIdJ3t5Xzae/u6
TnbOFTcK1i/20eqUh6fsGHU83Dy21aG6F5ImItmtnBdc5DooCJLpm0HrmwWAfHzG
uba3NxcP+vox+iLH4HSw0M6jIiFJXn3GXJFD6LASho3K+YuT/7ntGhvDTGqxJnOI
CQaJmSmHeV+VcZ3R+ZB9Ch86EBtV43OO1Hw0SnE+rDVwVkWwQ08a8YnAWtshy71r
qEt4z2StpCrXO2UvnJV66A==
`protect END_PROTECTED
