`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxQKKgGAUFV9Dl+DIqNbBF3+BVqtFq290UY34TudAUXvwasaetEubNnAJHIt03FY
OlXcuBdJrcArFaWYwaMrgZaYKNb69+b3GVmQil/0xQlTn1++a8CMiNfnnZK1xe6q
RC0AkEsCDznJ7R0ozqWQszbSiQTUduXBfGzq59norHU7QcVrETcJH1frgoU46NdD
ojetg0uemZpVCbm3cNS4FKC2/u+JZ70ShDZBGP4Nq9799LcipCHkquNgjfPCAt8G
DtxgGPyNNEkE92iGjwiBSbDGRF67el1CO4CW1lEP2r5cNxMi1O0BDAhUYwCFl6V/
xaCsVcTO2d/sLADdzl7wnRfgzzJ960AsUNCRq4ZFsxCQFp04wnbnBnkJLpM/1ysc
vNFESUA3LXIpc4YSsFG6OqlZuWe/fVSq+KCrW0ndZ2NlP9x+st6DXxMK5toSTSi5
4/JwA/6CPQP67LGdtgQJU6ppa36+1jRkw0Iq1DX2GtFEwNdR6teEkmCis/+UycJN
gE09QA7RuKleu7q/11KOYIKhAXDNow2fc6AeJEV96DpvwP0WH7FYQ+ZxCRSuLbC8
bPCLJQvpVbPC3xd8efSZ+izVl+FvFKP6TAWqpwLM39Rkh/r5ph1juYzSpF3RY1hD
GKyDKECGYLE44mFgDRL7VhgkZKqzl2FWTGkU62awCce8GCSKq4D29fzzBfloRf2h
Wi+HVUxjLJlYOhc/j8z8iTazD+fqmiMWYro5DgqXkb5sg6+A4MQXkSF86O+K/byB
gIW+Hvplp2OOVUdT/T0jhV9wRVAxZgpuQNo+jf+jvZQbjGP27qnuOEn0cVNdZi3j
ZV2FSZJVNFUV31lg4BlDRtU2+x0V3vCTYvuurUWlai0FJHL4C9Z/vo2hA3UcqSz0
t6YLvl0YbPLEb2aNS1GIwQkk/8sLcpB4xdYakFPWrNOcXzbgf0UIxvBWlkOW2Vq8
O6GhungANA7WGUvLdQyS1YWHMZE0c6ywSh6DF1C6bEkXmZF4jyGFjXTZ58pQsm+F
qcuqqDAS95ofPXrdyMxKhmvKvQ9K0jTnuiShZ3+orfQVPLNQFSDMvWKQK78YZuCf
CHEEYHZ9TbB1XqLTIcYgSPZnYPTeFq/q3g6XS2kyHjnByDW06JTKVTLP9VIrVmQx
A6EUoDPVp4k4ATkDKVIdQtFdh0G2iDYbuKWQ6c8/Gw3HOt/6oRJeIqY6GI4L527k
iXTO3X/ZwuJdNaAouK+DmWwfjPBwSyL5d+7K2MOE5ze9+ym8rrfD6Jd/Nt1EE8E2
XffU3zvpSJYKpHZqBrXT6aa3H8iPbaHPEy++rV7N6mZ5GRojlPo8k6R9qRpo0Wdu
o6hYG9og0B7D1A2ssUxtjI2VkDIJXItA/FPqKhWDkvuUyYFdKwZZwEQCgE8kCPHY
qjiXhucWfuDO0QQqOP/mJCBgUQIUviQq2Un9k8CA2dgam/N+WotAlg77oSB/JBq/
OEDMi3f4GWWALUhiACMx9pdYB2CYDEkN3I1am2gVYhBf/nfzKn0ogEajHphWycTo
LJPQeLKxcLEi5nNrqyu8rRedZvAxwOD5E1UoWeDstQ8ylqqpuaWZKs+OIdqu/19z
PpztsdNv+WzLmj3ZARKL2mfcbMaQcE8daUYz+GxLLeqhKO15T4xx6rVIYgzg5gxF
tjNQu85+icpwRe2gQa6tyhkToMWo46WskqhRIMILuQFTWctTC0m7uKUrIZwo9Cib
iqIY9stKXUSUdcGytz2XO2gt1p97nkdWgZovliHnbH1afBPEnb59F4BQy+3EGS/H
dB+hXsauIaoKUe+Gnt07jfGimpInbdWt8gnaOQc4OR6nBWdrFv4wp1tz42mXiNl7
UE3TqCYBkCqFGqWWx6J1zz8VA8RPBRS2A3u+jmmqyP9KpoApG7T5qyNA1XhQDQaH
p6VkkSDFAXJ6b5cvgfZvwJiIIeRxjlpliQJdgRvC13E4m1hmpJxIcWKz7y8ye21I
JJzWqAYHjqJT/eyij/KfLpCtHCUnOuxEMtrOUp7h1XYKgOQTBza7EPLP8KxHjwtk
qsAYxGixHpwK82QTN5tNOzqtW1Y9UE+/tWrVDxnBQLoG2lpLE2dy0b+Ixz5TaNUY
PkVNX9MpL2d4LlTNj0DYsMVo0LTg3U04fDg7Pf3zgpvcvFw2XdLRsoVItz7gb53g
loyv+BBdFO6jv/yETnkN2uWXHyoxc5bKyE9VuHiLKp37fl1zdVC+4iFZxp+3YfsG
vE/74HCHjR1D12kXCYHPwYaUAiemqEHsv0jBXXcWoM42c1MnqqYOwXfRy1To6pQ/
1hb9TxZvTvE3zxSBgOlTifGT1yU0GV4Pt2Q1Cz37Mzok5CV0ykiEVmzgN1uRE009
1KV8Hy2ZTD27QrUA8G7lVLtCPGLIlCajotqlrsw7PWlYk6RokqVFo5ljuMVhhtr9
AIIWtmD7io/a8EJTsjEqpDX3AKcUgdgUjWe7Tm28Mrjcy+HK+NxzXCA0azBMOtMd
43X29xl/b98YniW5LMXV9YCL9WwCWtc57CTeppqvjVAcyP2eYdvZmJuojJ3GNTd0
cav3SWSbXq8T9A3HoBgYcbTQXO8fbPIxbPJYFaBoaiZovYwoNWaiiPiWTaQDikG3
iIxEOO3edAoH6Ii19McJqjmmn5sUyvaFS3xH609zOXRObFnAkO4oMGgpnaPOGa5l
pAFU5VK4+48FxCOSwcw5yra1Bt1AnaUtAw9qtINuEJ0gnRhBYX1Cblx6bT8i9Osk
fIsEwZdnULrwuH+I/vgJ/JZOy3vsuh+guqGPtuGYFM/3svMFXTjmcDvh6ESK3fpi
G8p3OhBvbVH0jRl4tWm7hJqmKrBQoLuvqzdjgASfercPX/JzPh2hlRmsLZy9PmTg
BEwgQF2hdg2cBh2nLDVjTa22TrKCJ34a8A3us9jb1mzSPD6ACBAbGsLQ+OK6shBT
FFg6OUg65tADtzIHq6Ftj7yu2yEXMQ+NTq0h/KKKchCLR8YvRkl5JLY8fMXFrWIu
/goxcnnkm1tOaWXmW6GCvIFkA+ED8Mkg856QI6e2MVvZEpkA8dRi6ZMloeZWF7ew
32j1zs9/U33jj4kbPne594A3IJboaC9LCABSJMyfl7dZsNWysz3IDihc13TG2yl+
JYhfAsnZQHsZRXknG42YfOZwDnZWxHeS7bldWgdb668logsVLQH8xouZ5oia6Ofs
zp+Yy/K6lPTlAmtZn3zlCYcoDZcxNNLY+wHY1O7Fp4dlFCnyQ2+HQTAkRGM1XyAB
U4PUzBslAJYCEFy7zPFMMcRAM2/0GP4lf9zaWKvhx7j1wU3Ke1s0WfXkXkV/mNyv
4U2H6IrQ0yeYe/3qd+lEJBGmydZ1EmAeAD8W1Ii3xIcIFIGhz+jZK6FRtlSZi8Oo
+jcIsVrG+d3OBs+m8TVRBCZigq0tOHedsF/7VupKYRSA1dDETAOFu3nC4LCju/eF
KfSU4Mfh0OjPmI7LoBQ+pwDIerapUqEsrJoVDaelCYYXgSdRLv4OCQ1JN7N4o6is
dR28jpfHt1f5jaNf3t6KztU/4D58VVZyxVuFYOmZwvE0SCbhodG5vH9Fcl9eJrpe
k/kzvWzFhaFo2pi2PyjBMDRAa6t4ctQzknO7qB6e98M7QRy5vBs2uq9w4yA3x2or
wt7egVlXK4nWMiRtavA36VTPSE91kyOgWt4gCOi/o6NJ6RoACcgiSqpc8JD9BC74
QlEG++JSUB5JfNMNlileoCpPpCsLI/VB7Rsg8pzjZ9c=
`protect END_PROTECTED
