`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLF1trlTQbPzM1WgqfKBNOKlRLp7Q7R/LdXVISWA5ZwntVnZeCpRwY0bUx6M/VeB
RX2nxXSRxhU6jMRtMrfSzbFDqVvPMzEnqm0ye5q0eqYvdylLSDIYBAN+vIesI/r5
gN5VBtQZTF3r1X30QGI54FLBqP3JEs9vTOSAEYwxuNUrlsLh38j2PVMhMjYSPQb5
v03VTBTBSunBvdC8Zeo1Se6K6B/hauzbDU8BD85PHML1y0dtWUsOYBN/ZC9kodh0
Yv10Rxg2tpGWrBSCNwyPhd7q8/OEP0xqhOO0Q2Ugofrl1JfD5ZhVe0lmapabaPHp
JD8Gg1DDjCCb91Rgr1oSJ4O4xC8P4GmjWHC9VzV6T9SVhCB/bTqhadQZlJhGhDNw
Lrh8znO50QEZ3/DyCh0h+QA8SF6awzJlY3CqeRm97mPtQd/kT5izAhIdj5KOInq3
YSigDIEqFHhLbsMuspQWRS5DTlrsC2SZAMMKCZTQa7bg2lcK8tehZ4crd3zGp2Ve
5pzhLzaIPJe6a7O98Kch+jhY9mjQULyIzRKKnv3jDw/YsPaWQ7P4OL8HhhRRFTSH
kLUt/R2bkitqU99Vgx3VC/FEbKPJTW0akbwFSUw/hQzXEuiJLTQnAOaYQhgDaV41
HQrTr4SGPjY48OHr/nUZ4XNSEaRaIFzNjIiTrR5aFewoPOlU52KsK7gSZ5dENd5A
xHMjDyxHp392zLGf//CcKy3LF6qqEbmP7LvBEzeMX8a5zguMWobdv23kdK0PYb8y
zcUJMhadXVURmQqbNa6pLXxA+FMfwHiH1SyaZTiWPiRfRpQ7VsVR1UA7HUU2Elaz
F/UdAPQ92E23vcM3ORL31NJkAdKf0T+JbbrFW0n7ZrTK0xv49vzFgnr5sfY3+tOk
GfG8qKbM32TEtlWJI10ZV8BLYN8aeQy0JJ/NZU6wQCgTJJr2GBBAZfCnM/Wv2Y2O
k273z/WPR8U6AQjRP20QXu4WhJDf7R3j/nFv+a06/24/LYYL8p68SeGZf/Ua4E6t
k2/ZcAV4wVDUk8dyi/6QWwQG8h/WB6Cqiw4wgY6FTkN0uLAtTRPvXEuuoB9jgB8C
/10om3yL7hWAjvEZDbYAlhOaZpvrAJFfzyRyhExDCWuoU+0hHlOWoZquFlekPA4K
M2Ux3k8FOKwA58p5mQx/77wHZaFTY59JMfDHolnm9lMPDMpFdQuU8I7xzfeDh6hv
4600mhor80P+WLDwE6fkCpC4jpglXfpFuOCYjO3VngGxqLxfuN5vdqC3Icu9LSLH
t7cpJtGz6H7F0C1oeyLQJSg+X6I8cldS12ryMiGqpPpuktAXTpy1PXrViFxJg6P8
lLZB1gtWab/AaoO64Z0APrtNZonpo23ZiuWuDJ6ZCNjKjlcpPhBzIVjYMNScUW2K
aGyTCGNVHMkIrl7QXUdptfCvSb1H2sZuT6FqA0Qzbzc/dfl+YlGU6N0J40Raf/qk
oKxgkhqfcDvlUcGY1O6tv2JaesqvTX18H65rcsTl8Nrubk9xH2WU6HHrn2uBeDrU
4fj50lQx6thQVhdOzs/oHHx3Zo2OHSO3GMFvT+PmQHvLGkOk8Fh1isTRluFNwscj
dyJehtncPQytpUEmgArmX3mdxerml4nwK/Zyb5awTgU38NkuyscF9IZhk+O+sSvm
/kxA21AfA4g+gR/MXybdiJJYai8oHE3VjjxRZo0hnh81/ad4Mq2MreaZZuOHCs5W
lBR+fIJZ2/7x7NR3gZZKGOYMaRZUuI89BQQrB37GdteYAlZ7ZTRbqYlthb3Phi/A
HDfHBsZBV4kbOFi+Eyaaxe2YP0Ll3IUYO0rEzPtn8zVIMthwEdRgbxiWaIKQVKDc
8It9PvH0XpjcRmA6Ttw0IVNKy+q+HtlfKRQXMpa07OSsw0ClJQX9TrtSFZYYM9w+
PMnC20jn04rKNZflZ9/JCv8lQ8wMCdUfXM37oKwqqeOr0cVkkVBVEggPr4dZe0rz
pzMxfvhU5eBfoXwYVhnR4BJLF6YqyBnzMJig90B4V6VQ+kY7PGPoV5PV/CpCUAtg
SqL2CUv0jKsaWMROz/quzDMg55+P5aPgFCqUMpPJ7F/l3TKrNkCTeC5vzUnkxbia
Y3EKtBlVSgElMgnLYfRfse39qN523snL6kXRCNnaypagtSI6wtxZedQK2CnXwZmX
/J6BhIdaIrR2vBAfj4/XWqWPh0YJ8n4P5KkSbB62DDH77L5iksew1uEZcdMYHvAx
z9xBmom4uMD3e+Wu5mmUsmO6sOroKEsq8xmAi9zMsYJXIfJxIxfzU2LquBy7lQet
PfTE1m9Z8uv1cvG01KQ4uJynd8+ANOAbMbFux8OV0+9HWtaEYotW0cC5xc3iCy4+
rmT68uehqmj/dII02RY4NMpFnBIY7mAkmLstK6BJK1RXaKMdSirUFBvDyNjqBP8X
OsYgXq9/6FRlxHEyAPFUyB0IjDT4Caqy4xZH5PpLYzyaYwGgZcwzdwZWJprgIADk
PO/SL68a9VLTay75bjkNSAFtjjqwKB6u3bz7XWvZ2xd6FKGh5BtZ4vz8GwWQxbCP
ALOrQ7FBdvsCeTOZ5qJp8qXB2V8x+KISftuX/T8hSh50SDMDxPePo6d6S8NQdwLi
`protect END_PROTECTED
