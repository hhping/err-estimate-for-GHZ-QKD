`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vV7D86hnZKRtqiUT2T1xJ0XHzJd7YSHsufb10UrluVa5Enyi7wjhqHgtyVVp7Wsd
j3xWASEOZqtgm/bEE7j9dEMWevDyD6qk51liqbtiDnQSIY6IaLSk/Auk7YtaeRiX
hdO3rzaDWRpoifr+0FC1lyTXi0jt1cXo+D2Y47KUYsUwZ+MBqpJ2ZMH2ebCgHT1u
aDZQHSdc0WwkF3sEcC2DyRN0N977ouJpc3el2pxy3GtEnFCOSA4AFd210RGWo6Dy
G5vI/EKpSkbg8PX+KEhP9fI1xYj4R/FOY4baR/RYqkAmzCXVgW7NU968Yo73Qtq/
beaxjpVtLwI/zIsSneRzHEUvmJ+y6A02fJbItcj8bp61T8+nqTExtFQtrgUqn6ma
l67fFX9Z6LLuaFT1jc7+GjO+aMU9D0720yLNAOjZFZ6wmEixvo6kEqvHJ5jKE06h
b9kHUQXORgd78oqyOPf6tT4nAyCBSR+xzmiE5wEiS/EtzAkFRjrSLp+KWrJu8sgX
xl27k21plsd/rrQKnD/BWVrr69CQmxjCr7/UmOIBZpFN6ZSSvwMUWuNOXqqwi8f6
PgyBQoefJcWeE50r3QBk0UrffQovGlE6luiUA2YEUGcDTD0VIhpCV5CKgODdX/zV
tdrIZHsiEZOp4itCtpm4lxFkqOilITIpwgL0F855Un3wgI+ilwH9dm+0B91WV6eJ
fiMLeUr9JzIP7WxTmz6XpMQXiXbh1b2Z+0//BnbN0bykC3Bw7LqnV4gHJ0hiv0Qk
lSGn3Dv7Ee5VNBBTyp+GvAKaFwzDzj4tcpkJYo9UEAbBbf2dHd243Peg73y1HgPB
QZEParlYjudUxx2Q7enCeDU4rrWVtrl4EOYhpv6EQ4kG8+GnB7w1Vm9PRVsbNg8t
SDbOaW5TnS04fUYxjrjIMfqKfFNaV3rSd6BFkMelEN2wTN7XAkGtXfD4r3yOuoip
oc4zLqWpmywwW8+6YxPnxNIH7+dI8pew+Cdhr/aQmV0Ps2FN76Y4m+rc1Pij0W9s
9GHhMYdge6Jba5DFEN/aEsEUz7Bjqm2kmrBKlV3lVHEgWwH9UBIig/okyieqjMuD
sPPCNkZY/6fJX314x26/TIFZj0Ld9Ibjr71DUsV734aMcWLrIElMjTabFuB0K48z
Z5GFlj0QyUpQf3rQWZReOWsP5SShHntWr8Lp4/O7rGuo1FfQY5PzJurp89LQ4iH/
RCy19qg8iSsJ9aUKLkRVNctnPmnKSTtNgX0MZFmW/xelps9vQiS5VEfVlGWFGuyx
GumhIJeePMrDOV2qIbX5p0YAE/xppu5EH+6MNtc/vh2KVO4JmdzbwJVcru1W2MtU
4d6PW71peICF1fD3Bc8r/uh+D9IQCvnCrC/tj/aYM0gw4aroj5bBZd6nviHrWgN/
rFAZoCowaFv9Vn5N73YNWJNLmenUvar9gNmfP2o3La5ejz7FlY7D9YkLUDs7vOzt
bDyVKTxSgJqpsm4/nknNBx6NqeF+fdouBNUqUigSbdnF7/A2/aG/gZ/fcrezhx1+
g1SQlcsIJonowUAHxKJUlgjnDjmht1nXQAS8pWko+iVShy68cZZh4A/lc06HnSs4
GuBbwz4kPh5LHzlAUh0X+Yvy7C0RQNy79SeFPhS4ZX+q8Qwik9R6QGiazkOWcS1r
N7EIyR0O1WIor+d8ipIuJd8WcrFw4Hyi5W2lo6Vi75dwklo0nzg2TKUwUSPvW9jD
9guhD6QEs0gmzq8AhWxVadUNYAH00ud0UXzduTrp+nn0PBiiSOZ36Z4US9DYOFQn
j4w+awS0wwae3zsCdyN/wLJcoI3rKktPWDStHpuJxyLtieqkbvMmWVj5owvGeyCb
FXWzuECQYHz25mpnwrlFj7459WSlzY1/URruwYb8rDCBk/PczOhG43hHjaX4dyr1
KluZ1d/3igBZwO0csZjpf4nSGhcp/KgvRSBepWVOIgpiSQWya0jLQ/uebk0u4B5q
54UlbxztoH5ebSgxVg3OxURu1en7Z+IH5GG5DmSEdFFQBOeUhVB+vZG5Vh4qBEou
YKC6doRfOsqoo2bjBZWJpxEGMIhNgpoDSYhxXrC/T7QnbHhRk7HBvleHE2Dqkc3O
5+n2OwZFc4RirWjUvMtuKDI4q9rGZ4ebSk8lMdFDFj+n1CmRAELCSd2NL+OsXX4b
oIloUxP910YX43p+VVilxqqT63VBGoLUiIOpv27yj3Nl+uW78Qodya4Kkw1ZFWrW
1I6i+DeX1acZNdjwluaF7KZ1/ZcGdYKK34Lo7bkTN8vwqN3+2mJ8yrGvdXx8ny5z
TdSssYZ5c7ldvd2WAvCp35HPuNpit3BizJBbSPT2fq68lQWBgfhEOSXyJKTyvR2O
UrF41EusGh/ilvV5IwIOnnOGYaXnjMs90cYTEL/2IcCgPLc6UVXoiIdHVAHBi4t+
KKmlgTSwWAwb7twxxWum/vTjy++s0GWkuchOavZG3NOwt5GjVplD6Y6R0XOGilEN
dxk4ddTwtkac6wlNOReIeCcrJZ/2prG8k1YgBnJo35fxDsdJ4o1sotbKMEo7Dlgd
mOHHlU3q6aTiOsl7/KqHBTmo4EQhXV+rkoSZ7I23tnHyvYsXYtYkUCjiNmfQL7Ik
KQ2pUqLOigNinZd0+OFAeQCD8RApuqlniyGKxzm845rcFSRO4BP17Mctkhu3Q6BU
SjJY6CZOslUkAlIwHXS6LBu347Lsy+Mf9pcAT62YIsdToTZTKSBx6TrgMnnX4tbj
ri3/ageIdl8oIv8MaT1YBy/o79TSHTwFKALWlOfC362rAZLTdlI9GlTDsH9xoTTl
xtf6BHRoH5X8lNfyJD2onOQVK136nMNgqjiMw0/noQxe4UcFH95/lbUEoCvCZtCW
Mo8a7E9hV4ur59XV9BjfVJMr0uzs1/6dD4BoBNiVEXmOsg3W39ti5prpVTidgTxe
UOIctl7l3RtFqSdjolivbY/ZBbAfrbCt7zqf3xvPD0CYdNRBvLlYdjpJBKPgC/kk
tFSxl3KvZBloLqUAd4CK0hBmgdUu1b9AHXtK+/zZ0wHvmCwlztFOwYdxYuJP89XH
NUMtcXj31aeJZtBQ6aojsqpyejXpMLtutL1E1nbTNpMWTFPSYA2dl5tRdXAm72Ya
OXrD5HvC53ba86rYgq8RdU8s6j7T18lgd//MplZkCjG8j9IZ8HYbAAf+5HbMJv7S
yccybrAanjV6LlZRGXnJ/Sz96MGFnbL/PQChAQwCNv2EvNd4E3l2djBBlMF1UeS/
udwWYaSXdOWrToHHxcVQ2b6HbfxEuyG1VUpZIo8NjFFqVc++3WUZDtAT3eQx1Vpv
8vG4o5cpV59WNXf3iYNq4ZIiXhox2Ycq64uRzxzV81lapdgqd7Si+xLL8e7Hs7AU
qhdosYeRFFVw6mogZBU6uL/iTUkOJiu2WqLbpLKMIRLMrWfyDS84KjiLaUV3d6Kw
OvZr2v4G6AxWLrOmk/gDj8QcgcBK9cGqndpBQc7NsMZSfdttWflzwC+J9YlDivzB
6ROdHLzV6iG0mGIKA4L3s0BEx9nWC1Lt/xjiQ5tEUW2cj5PbMCde9niTxF02+iBK
1/LaIuy9TMs2soQcVXcjNiw7Q7GXdAZ6Orh9osTmb88AIbNv6WfCqYKxawJXBHQ+
h7v6GtfZaP3flOKKpl7pXyxLdvOwuj2Y/k6jIjQUvfja4a45cOH1zwRSRzkbbeHs
cgg1X2hRiL2LbpSrWWlPi++QJDOyjIINCiO+llpCvSy9vhZStF1KF2mGPvlsk/Cf
68QeC6TYpZcYpS4hx7elkjztkxhKHnTwBZ88ZDnqDz/7oD6QI5lIS/fWXPlaDoG6
eEcedz+Sd7O7RiW4yAWJjGTVoaOkdKLD6THgrpA/1hixxpag+8cemR0F3h9ujdS2
tZpMS2VpBx4eC61PTGcKNrPlSbcQtEhVDdZBKGwyX0q4LJzy6Rtd+A6SlIk953/t
/KoS94B3UkO5j3QGKiHJ74yion5pFdW6ZT5MKXdUojUgLIh0CETTgSsH0vKqUUqR
oxjqb+69LmOvdT2ritHAmHdLER+wxfDNLLfEv+MBtvHxD3wf56oMLX2Z5aJw7v3e
u7xq0dX6dFAE+ojv2YXOtNSS7tSeyJgEjFD7GViVoCE6bRsse9crT2Zsro/zNTgN
AHEv4BCh99Ea9OtIJaPJhI0/0ABFv92ZQdHMGjt6lf51P368bslQrbqcdy2TBWVg
k+/kPohexm1fk0HOtIDIH+QbcWCwFNXTObVFKhhhjVL/+Mb6oZNDq+PqsOQCSL1g
yFLHLonJcebxd3tUtal/osYhddGwQh8M2+BcXPZJvwn0IPSBTAshPMJ3V3jOgD1O
aq3ScLIOscZaEluMWXnVX/HvfWj304ePAk+0NAPlsVpz33cMIm45rQfU32DJXW2N
SmVXWWVrh3UKdsuksPkldBNs9BYrjyiJKsTrvpRP1Bo=
`protect END_PROTECTED
