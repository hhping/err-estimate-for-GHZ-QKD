`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BmoWPEZO2/XCMibu+rGUnbmZ7eWHYEYy0L0otOw4CwY/+4DGtWeTPb0n413GaDcB
QfAHeraLLZaTilJ2izKtuYgY+lhf0tcdq0wJMg7ki69kTyNnsVaiH1nYH9Qa6Q09
McVHgXm8pdbFRywYUX0TsOBpmETKCx1lqdFjDC5RPtPiIeKxqkP92L95duo69xK/
Kp3jzl3KOTV7ucUKHI5ZGAKRcgqEakGYhxvcpUkMIVI88GUdP8AePAdOHSDvZNHo
psCWpsSegMuBv3yVF/Di3LRONBP7ivze0vpC0D467LjUEe+dDIUhqA+CkLcsf3xz
n2/4Mp+4K46N1cIvtU7CxRSPZKgWCoRVBtTshZQDhuFPGdsZUeJNpqoBVeYFvVte
rxXUy65Prof/9BRD3m60bI05IpPXB3cNHO0E6co4WFVdzPwVz0enHHsFlvmub3Fd
gSBC6cG7qdz0gPp7PzpMF7tDQP3BEBZ3MGuHvVCkL4E5znChvXicoOIenEV4/dr0
e3+ZOxQnoYja9U/oUYNiadHp6nzWhIO1m/4R9sJiyQiDnDGIyDALyk26bhMfTpQb
qG0tnTceuXmbY9+1T7doZ4Z0bLYGqPBNWL0snP9WyEWH2S1Q/6yYCvwJJnFN/dDD
ho3il6kVYplNzj4oh9KrmpECc24J3w3aQ/XXiSh/H6mntdcYXhZA2ixF8Gv4u//b
E42NWC9ewyou9XYyfW9zIWBGTsrKeHMMtPmYnkwAuQW0MePa502YPBN8ZXNBHV5Q
hXb2r8yhWMNz//QrSdto3AHCUsdccM//GXwyzgkylL4EAyE9uW5BipSNvwaXa7uK
73I8EH2tPJH5q27AoRpCnR4hRQZLJ8JGO2JNzvdmJDA5JYTpmLiBn0VTYvM+dtOh
KPEgBKRPJRPl8L8orX+HwR/k89VCaHSC/4jkjMoNjfrNPWf0KXcINMchQEyAlsN3
asvV7NAuUkLs4MxAgz8TVYpju4GjOOG2w3omiO71IHZ1XWt4AAJCvrZ/7/RppaYz
kA+0EE/4Cjh1iYBb1tFkKzytYyCYL7gcJtPmBb8KgJTKwdHIahzOSBpLJn++z7bq
3oWmZjXDs/7eJYqSkNKWLURCZDkoTXcuRaYvJVugMpkvruom1A1331FYbbz95kly
Qf16Kb4Q/x6kPnIT8XrHFt7Orb8qvQv3cz/ke9COyIzk3bPZSqK+CSObbfnKkYFT
nYZ5FgEZjr/hPeZOuPzs3mJJq7n1sH/A7xagnxoaKgZKhmR/37vp2C55SObwetYC
/nNlBqRUsBjPtTmjTFtecuxCaHuobNmqH9LbkkJL3Vm809t1chyH3DpQccU93GCH
sRGyrrFv6/Q+y4NvUGlBogUaYrV0ilyMwuaK2TKKfkcE4ap5plASYCp1njjK5gJ6
DUzxo2ZjssUejMFyiQKLnRKpRLDUKI7f5BIHQVXQVhhiA6b38zbQk7hD+qx6DKoD
nGffDsoZ7LNBLElIzap2RMwH3Ra+FvnqbsYRxmIdP/FlYWIFbTa6UNafVqVt/56F
Hjhnf/zUQd8OQhDvPYwtRXG1PKPE4tEW4IXb/1HBtk+vcXTCjCBnYtKPVa8RvUfN
lSL05murnC0C59sW/3Ukek57Gn/cyx3RxTzOiwgnlIMwmk1F2eWUGRZs2ZIdhH1k
dR3ztO8jy5onInvE261OZHT4lFiL0YQWR88hHJTHe96Gj4M0tWO3kUw2Q1obftUF
SbBtyeF41+Lo9U/csIE6e0iRqSFg9bOAmHM+zRsegiWu9hnwCGHvZpg0dMMbFla/
kNYxCGgnwmF5xPzBwdmqtcmcgS30kmWcf2LExTu3pqs1qZb2j/m29yfwa9dXz5o3
A/30SLfEphyTDb0UGTaAA5/FP8y7AmX1ZHy+eSmDWvfiDT15KuhRR56fYg0b7y4Y
iD99MBJ4Iy5XV656b5IkAt4YaQ2S1jA4XleOJ8owEvf/66LERJsO09jCcRhNCWQu
Aoh7YaTSsAtKxVN0jrZMY2afor1tDiestUGIivYTXhs2P0CmwpUS8jtU+Q9qn2m4
UJas9QJJRIgQDzd/of+6R0qcWy2OaBg3I6eDmuReEdGn1s2A7jBSXsRYV3KZAKIn
TLka8kAwH4+Ktwa2l83rDG5Aa7ZQcycacfxop9n6dV36o2K+VugKEdHYOxvm+nq+
DlCje6P1N6RVFXXC8rWrzdmcnlpQKHry2Ij0V9Dxyz2QVT1j18u2MMLS/Wi813xG
`protect END_PROTECTED
