`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BhDDq2NdIvy7qnEWv6hQeAaeOrCFOL58t9onIqFADc4WIVtQaaIHWXHVsrS30K7x
JVGcrqPB2wgMiuoSnv6Lpo4dRZcCRYaMK1R3GIssAYT201mevYm4TrA9P5Fg0RJH
JXT08ldfwdT2JQjBZtiZ3WLU51tRHjGhj5FHQmxhA6Nos72mUPc6lI08RST0BbtW
NVFu+i6r1WFlGVOYsD7yUFnUXgQqAoW+leHguikYomAwpg72JkQgKeMfbv1GnmBn
v2KggMIaH2sRHn7RsEjnww9Amycta+cxfDIbhwaBkQNcpWHpxXJam8+4O13ziP2+
tIenIthMLVCrGVEQhz+N74syrusAWu25zCSI+SFujhbac0prXW0Vu4d5V0VNTFfF
M73flFdOdLKKd2G0pEFC86nmBjvERod6pUK9toRxXgaq7nKK+v1aDJdWSY+UZkIx
+tzuX15gsfVg7d8pGsjJkzv4Ay2MK+oxdKLkwIzh0te5FA/p57gbhbOfFxaOkllZ
1gGhBCVpZ9MDyHMjvaWWLDet1XfQBL/vXMxEnn8IRHQQ0lZrqvk+TXNRRIr2I2y0
c8WDuD8/hlKNaVPveuZYpvZi3XMk4FLRv4/kN7JwYclhwhsui4XI+klE587A9aE7
5NZuAsrIAECwkJiCw7cXU1IsMiRvLJz9Y66eYZAirB0CZ41ekBVPxxMB94BAi20w
ZkfsDkgftE3Tyl+rsbNBzrgxjQpxndejASZmOFpwZtTJie1CRMYu6kvg9eN4BtWz
gz9oVz5omt9J2CN+u6bcCNqXWkvfFt7RcdlmK2bKkieXJV4Q9r1a+z28x2uWJAZM
Rwz1U54IddmhijcCcuXzYQ==
`protect END_PROTECTED
