`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wlvnUwtVA7jzPGebnPGxg1x+4Er/2Uib8qepAv8qggoRzFuyTgsmuWDGdU0JnU2J
iDy5LOWiLzhiIsLywMnvPJTF9RSf14L0+Rmk0NQYvBvRLK1OUT4rWbbrDGL7H8f2
2lLnGctXxViq3OGxnL9JqGvHVajj+JGGoDOxcdipp9aL+YLlKHFUKNiyI2GwcQBP
EM9liwYeeRQNPWAN5+421brpgjAoarmctEjA7s2H41pLvTc0YB2QBTClq0raHjMY
NN6p/QL49zbs5SlwXbQ7FaDe0sSGJLsVqaljk9FjWcBP24tLRu2cWT3LjqzuQ1g7
5+UuKozJbBbiKYvWZY15YCz+2A9So3AF06HSc3K0gqUvZsSJIr6lf/f3YGn/QprM
mE3t4bGrf5+rE3FHNwMGfRk8+WzrHa4lhR3ALC4fvQQ=
`protect END_PROTECTED
