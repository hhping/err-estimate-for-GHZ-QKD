`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3/n6cyChu6X8avytDKQnUV3JKVcNo99ZmINsgH2o4TvKL1iOP0aK8v70ILFg9+Mg
GB45oG4jwt9zAPWH0qBPrD8NhfOkSfWqb2VZ0JYOooiUdrnENWMI5CCY9M1ml6KR
v+3MC85MA3L1y1hwyYAj7/rvP7wDs1XXIF2Cw/OIv48zsqhDuN6+3hokf3rLb5bL
bLBbm0LU0tOhX/VrR8Jl5FylDPosb+wN3LFpPVpm2jA9d1NXyW2LxCJYAoe9Sl1K
Yb2XsZouS10ENAzWxLphizbXWeWWmMNHdojUe4fAayUtwKvSRm/6Ro2wL/+8I1DY
NyAIyjHksrsKv26j8eEMd8ruvwf8PokQ8wwq0cSfIof3v8jrOc36ntKlkp86TAnB
1qktouA1UGaTH/w+Np+gf4K1o8xVzkIXJJPiORBAM19RFZSrQ/ScHbVwOqTt7SRD
EIoQumJVzOPxurGEojW0QNGXi9DG5p8Wa9rNv7Ln5DDGcYk9mlPyRaxaWw+dsJk1
6540n368YDjOHEKm8JztBDhk/pZpZSFlRykGUXaDVTkpp5OGFlHantjzk035nuT4
778bziNVHGFhUMAKsrzzq0dfuLJ2RvooSB/TtblvNhACWSAodPguajinIZTQhejb
f4NI6vmLrDiy/PmX/lX9r7sgObizu0q+xFicbiKMg3g7fxTell7Z+X5571jOC+U1
6ljpm2j72a7kybpvAYxFbrhgPm3fTFKAQ2jw6WPqm73zdsiuRFUvOoE/StnetZoX
bP43WQkQvCFkUilLuxwCvVGeOMVlA7hSK73OSnHy/U6kcpd/9XJ8bjy5ym2fSktE
woP5FIfhjigdzdX9XrFYDSHxoQBvsGO6Wlu4MDOzQi79+J+fV7HRzEl+vGdQ5Gwf
ujqF7xAq+7yJ4CdFqxR7hB/vMkkZxEjAuIRkby5t0FSBFDApIQLKPacFeqFU9KJI
5srmFF6iCPnZq5Uj98r9DILNqHBqNEwYpkS9TSArAMSLng/DGDiCGzDco+AKlUxq
dQ5v6CKBS/S4CBYuOEkxnb610eblQF2CWpTngrgOGTuBFNK0aB+ICCtW777jTtny
KtAYdzjYSDVgLXWzSVsuMQj38mFRGWifrVvN40Ib/R+qditUWJJ7vJ/WbitF3Lru
SLQ+VsCuCKgIhrYAwovRZ50z/Ned9S7yBgbRVTawlbgAzGhLiCRV7WdoFuDWCz0V
OXJ7/phGh7tqu0X++UHvwJG/C5o0zWUgstCbrr4ewRULZoZeyu9YmY0pKf70Aarv
pzhmOv+1GXhR1+VhzRFsMXE66FOIklpxd8QFAWpd6so4tf3cvaLB7nVk7hiUT9JH
6vkPb5fy6nZDAwonV3XVMwEU/z4lLU/+OeyJX9CRnHfjxFI46AtOxzcHfz5M0cHN
fhHSyG97/yxpQGlyV1tRhfj1/+GXmYmH5lTh6uAYUG2bRLFEy4Pdaqu0LDjjBujR
g9NddXR3kkUpLh0+sIE/YrIQ1SMJ9MDQKb/TbUD7r9ykCPgmpjanf0rhA5Q1+Tb1
X4SbhkMbKz/pP6Ew1k/WaXK1GbPtcpJmWkM7ZozhTxP9q2RRopRoXsMt+D/kdS5a
uzno1WlpHD/vvFcKKwcw8Nr8UXRdp3GfajHtCG9fW4yAacXWoV+iC8s0rIMFPOOO
FC5cjEJ12nX6D7b6ThdfavyOs+2TDe0ZxoyB9IYxz02qtUfPRET2fWz6/JSozBA0
h1bZHzY9RIFlfGMGZ/GCUzeZZLVz6yfLnHiIJvdR5flCQUEtVpB6utPQqjjyfvel
UxIdELZmxOFH86z1ueM2ZwmmhffViEk3dIzTuyRVl8t1dwhoVUMbYrkOtps9WCP7
eRwBKlKftVFZChcDslrLV7B+EI5hlpUALvDLH7pQHNDgApDL48rDfxXcREujAqvz
VA289uvrYYVsBFarjdWI1P5G8i12K4gVtkIECaxWVYPEst3+h/PRVAU8lGfuKKDr
/WpSYK1xMMsnpwPQA3cRjj1Pl/H4zlxz+KOVI6C+YJSmy1h5xbqd+ZuuMEKKp/It
AKz0nVp+8IG2yLkZQLTr/rxuWN2Iz+MePzSpjgH6TXE+QYa0DCd8nqAE6mHYYCz9
Gse2urftWibyIS1MqDCn3RQXXgFRMvM/U6OWGSPPrpqonqNIwe+YaZ/dg4vtQlMT
szG34Hmby0PA0iTrrcycky9oQcuX0kare0B9QgxJ9Wc402ml4+v7VjyeAsoZXoSO
vq4S0tiMabKAFzGLSjUjMebm1Z4MbQrffiGUyipN2LfZCDqVKlpYkr50GTbsx1wI
GeHp+i/qa/7yT/F4v7BUQEN2ouQic+ZQBY4JFIRLg2cibvcDl7Go3gVU+D6N03d1
lASizS78TnkhhktFbLziLgz+WiLxpWdZDEIRECXAppFZ1B19HilksSUH8YHtERre
5Soto6tBD7RWDzY50nmEk3QbHK63+/xhMNC1D+zydKpbrk0Fxq8u5juiDcPD5Xj6
aSb2gH02/ZR+zBN2zcRHjzLNkjgi3aaGkKsNtULRwGHk38Ngs0sk+nRKjZigT381
4KGIOOykGA3TJzQaq0nlk4e0TKf67qqbu0qweH0BPezj0znc1T6i+/1J9mIcj7k0
XEL/c0r6l1y9knrVGQOKJ5A964wntcnkx9xsaSQ/YduPG0tdF673km3MFsbx8F43
k9KqfVaYd0tOE1dHooRJw0J5aKh2r/og9bOmYunDG0QsS9klVlTn2yd83UVUZQF0
2piTsWCRfv1iTsq05duJBRLVdWjLWmoVk3/gIEuSAxdrwYgJCdA7Hu3CvMN+V9HB
Hs6J0FyNmuE45s/1Zyofr9kpf6EQ7t2C5r2QDwtSk5SmYTvRUHpKlnY7Ptk1azoS
WtjmlY9u74PtkDfvoZeBevD1zbOlQnqGS0HHxU2ba3paUxc+9KP6/iTEV22TOZgE
fV8VxAvV49X1qNTX4zdmL4MoKwX6X+y1NKQB+yRYWIxwkPWNmEF0YkHNgznqtaN/
bvWCqP9oK/cd4EW7pEcC3c5AfiM0CUuu7Y7sxg3oipu9h8lzGqTiW2eajlEta9kq
Rmwh/C08V0JTsoKmbDrkNCvlJKoryzxROqsE22UOPVTndqacTCNQ32l57ZV2YHFm
bt8pLKeDF84b/fIbVghQA6pFp12Y0/XRbRXXmmwW9TH459Dc2iPjz/J14kpQsBt3
Ah1e4IFNTDDMMsV/80Gl04pPkycnq4lluLcKU48bjYAWF0kFqDIdS4UKwDnX1Dj5
AQfgzyOvE+sDdZiBVM0yYptkpUTyDOvBt32FUlN/ObGOsqHP+tBvVphS+ngndc33
fNVGAZZDcPK3cJ6xNWBC+NINyIrt4zLFa0l3HwcS86Iyhj5FgQ1+RVK0rz+IbJaO
bR5A6fG/I3uaQfN+OZCXOw==
`protect END_PROTECTED
