`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGr4mKWVFT9T1W4ygSDS/7RYVu/CxX5Iah/LnQRP563eqiS5CGHtHsSnyUJZzmGN
eIOgYRxbfq2olwYxTHupEKzSwgUejL/KJXBXTiyFaYWjH/bv+oTXe6Sjq11SXy3O
vaN7AU6PWlOBJGIibNH/2TGmY51k2HP2g7ESK81zni3gNDGE+TETMG3MfWlksDHP
FFlw9ryMYKLV+8g91PW9V/CWidXYlFe09lLrj17PT6eOz3CfhyXgV4GFyPhRbb9J
xmdghnZ0Kzvt23jBNg12NpDTELC629p95TtGnV36NZLIQLajOGTNWitwq6CgIsAz
D20BkbSr8Vleq60PWBmcO/J8rZB0IDQ1Zl/DfGdnXPLtddn9WhJ0Ng9SZcwg/1+s
nZz5E234x8Tp9uSEsLH9v7gklbsnnV/dM1RGVBLpeexDm5xx3YDnFdus6XtIM6cr
XJ4QD6W90lMAjbShozYz4L8uwIqcjejIxZ0KMfax6kWMI2YnP2ecbELiM78u7kZl
5mZUt63on6L2ASLM0u11KKy0rfaV7wHfeAly18NlkDlblRy9AWpw6nIBRnmdrzk7
tK9NaWzrTXBAkCGdkgfDnRd9v1MdVHc+i3bEHvDBYRPMRxTXlUZZMWqtcIYSMSdC
oMmQMUej5iTO2eiyE8eSjo1QzZnTlZPdLNMSgRsUEqwlkmUzX4wdWfLYdw7QxqZL
SmiGhp2myTtER86ttUzWGdz2Sca3qbyiTRk5OsilJ/bgZPolPHF0xJbhwlF5QESY
j77P1QNcIILZVRF8gD1BsMSnK7e8TH5JYn6zdHU5IYbuap33Z6pBLI34gecbMCwM
uyZtVtJkvRvxN/swZPv+OAWty9a2LKTjon3DxwzOrJCU1wt0rULClG0s6PHclHCO
wYY9IKGquJR2wpZEmq5NwXeyIBFjdabi1leWD9L7fLcU8Z7dOduaV6cOoWpfp0G9
v+i54QqK6lAv/+BdSYiBeECUhjVrIg4jM9o3wOhPn+axWU1z6CMYTuBMNx0t5g0s
yP9Oj6vmAuD2RLRQ4rwcmYKXLn2rdepMpgdPtmxLOEf3PjvzlGM/3WJWOoZHRX/c
sbKZYU7jtt3mUq6kg2VSLYl5lTMMd2YvpCkolvwbpd0B5GmvDXGT179QkJZjc2kQ
bbtOaCBP192pXgq3HAnEK/SuBUnXuuquaKQ8e1MvbjO1rbq48fsPVXIxtf6pX85K
EJ3xPqDS/BSgk3VFQTsk3QkXnkHwX5wbHtNA7DHh9C5sH+yncDEUhsbYIEQzvhqD
W5v/d1SixdE+ZjeX3A6C1kRXARfmGnvD/jzhN3LNIdIsddxRvQsMeTr6mYv+AU40
VwazLnMMXT4yP9hJwCpCWMbf5dNFd0gvAGl2nC6toTRsxrlzNhITOYCGAWGc1uc7
/U4WQWRxtYLgyWEFORgnGvsTqoVF8Jzj4FuZeEoWnAGhFFbQ+lEBGwfOjgUQ2rMa
CsOZVL0ast0hL8x2O+EetArsck8pOP0rB8MW9tCYsLpvYGFCKu2AYuvzV+fkScYY
fpi4eohljuapQBHg0j6SEGtOUfZ7+mWL+Bap18Zh2fdxvDigIbJLzD+X5wR3CPA9
9fQg0ecL6Fwr2wxaXJXGJ1c0wpUwOZ07Je7LhQMRo4xPRa/buY8dpG6OoNJ9/WNU
HCXhkqfYTW+Q4eg3hvPFfkhw7vucaAJFMaDcQUTLyFmZtrdsV+pI8FuS5OGswFj6
iy0vC7Klq3AGiqDZuIdnt2KPJjtAr8/J32Xw9i9rQyx5624dMLblDWgbiN6aZVjt
/z3thY78XWlkITL9ILeVenAO4goJF7L9EEtwFEWi9qKF7NlYxn+7UQp/VeCwY0/N
ffsqjSZOHK3zyq4fp/dUfzERSAc/HTO+6yizFQhXCAho2BYJFQadx7sJLf96dFcD
8/YsYv1OoR6+mSLFN1ZAqZxL87He6fsp1CWZlhypfGtn1X4RYuBJXlmZUrCJXd/e
7Qdyq7vgduN2BZWyUFIJ5xNx1KKpFDGoxTMdEmGsr9Kf7OkBe5n37oDd9mn6ni9O
KLEoUvSZoCdvLNALT0/4UojH3GZRW0FHTv8nKijYLfRs2wd8/NvBpF/AidoIUkMR
BkooMlW6zKkq3GhanY+ICIecCIopGp5Vku7M33tWF4RdsffEEr2Eoj+brz3kvg40
l0hiBrTw9FFHkK/oUUaNvtmcAdBwpWVLgmHaFv/ywxwNhnHoKBZPfPsEp/WVO7r9
89OcRzqoGwH8IJkt3aRtqCZeG5HM6i7ktuVZm2wBVCWQE+aMRikCyr0O5Hh8vPrB
L8BMXJhOEcHyhQOCMh1APWI4ECl0ihxqhEcWhQ/Iszuev0Y2ES5Xenvl3nF9whmK
M17T4mMwgLEMqc4pdGVGtPKB9JMseYLYZwNdd/Emt4uJs4FqLXYPBjm0pCpRwXWU
x7Bo5F+hUL2wdUjhSDwEorLHfZQ3RC+Dq3u2KQseC6y9YQ2NPucS/OBA/w61Rfak
3ck+Q7pss59ROPUBO6TB3Q==
`protect END_PROTECTED
