`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0I0UMd/px4mjn/Uq6qV7wnQMmBrX4oHbBqgNOHYazu6cIYM2psHOBCPXcs3M1jg
2WRhRxbX6LIsoj7VmKyRDBpRSbOSP5BqqL+2b0vjXt37ObIWbuISS8yfUFOXZ3IU
jXCPWC3lb1GC1gak4ImghQUbLWJDTMC2o5zAtYmKd2/EgaBHHSuJtYze53JNygZn
DqlQaORZCFdrGFR6KTtCYK/sSVhWoV56Z251ve53B/r3kiM7ZH0UTSEo+5EKSSvD
PdEQEFMkjqP7I/PgPvwaLOX+QqWGT7dw6Tu9YglO0V+3yr0njdVnlIWj2LnFrzfr
pQLRV8Q+xwOAkOIy5KVZuk9v8jV2CGk5lUqz3kAmncnViVI61B6vqoYu/4zZxoQO
nrLLOwPHk2SyEGJhxb1Hg5qq1ypmEfAqpGVzdez+FmhfTdan7sgnDq9/XQqPND3G
KEk1CCqQH7HetAmmww8vweYwlpLSqqsOVrLnccqdsOipA+Nx45/ROdqutR9iubPg
kgjRkVGL33dpgb99xrWsvOkg+0UFrki2RxXDdrKoTxnGvyiYxMa9HOdLJeBTMLTg
DFohpkBhe/WoeCh/vOltYsc7Tn05iCAgpMqHJH0BERJIAvFQnaA3zrXR12um+aaQ
RMbfKDetFmpbJ6p3a/CgUb/ynFxaaY2CaybtyANWE3xk9c0G7kFG2wj964of7izC
VIcTB0ims6/jKkSKgB8/PD50mwgDU7AsFcxczvdDFVAw2PB6OQm38TbmEpJRq56h
mNfY3qeLfAq2HNb/QWmFXkAPuLlu6xDhpg76BADeH8581R7p089qIJINiT315cYX
aF8vkixMNQgWmuZnhxe/z7aiHO3MN5AHf67MzmuGeNI271m21/7QVkOpDXbwhYdb
soscQIHzkG3nFIqm/i2LCo3i8DasQKqMvH0+WPN2hfPawSHJHdQDzvSr3wsV/XdF
WvB5SgQq5NoypNszIi72+zVQ/SmuSj7+jJXlh5S07EVsEhdu3ZhmyPeN/T+q/mC6
Jsyv9EfcYCvgJfxU8VG/7dyUrSFT1L8OtvUu4hRdRIO6VhAAFIt/BhVFhptcXc9e
VVzusFP2SBc25/8rF2vO/gN+7O6BMut5cjF1675kD/aptQ35eB8nxyxvOgkWAIcR
szFPBaIuGaNsWV8JgOe2SVaDWu3+w7VkYUT0p+UZhNhI+PxE6h87AtZKOTOhpJCj
Fx6WJuOri8LYcBdmPzPZ5e98phwrn5L2rz1OtH+tHOBrUGWNaBgD/LH8iuhkid7U
8jJJkR+S8uQWdShkG3WRHVUy+vStqFLBdr2qRyJZNpiJyfwnsyGPLt9JrmiyLBo8
eMrYC5FlA9buz9TL75H86HpysKgjSeqCZcXdlXKcAbfpVPeXghX4T0vdoL9hl39G
llsbn6kHIgV7zKROuf/cDXS3nTYuKRL+jeYQT4kiXJB3Gf3ngD742GhjQTEErX+5
tL+KlP5Btxri17WHT1iR9Ycg3MwypD+bvPKcAz6xmZDnLzggfVFeBFrhz8kF2F7R
hC0lZNyo20oCu5CMOgidXoJ85d2sQYA6ya0/YG6k+3B6cn974LBjGTJ72RnBlRvn
mJJjlX5zNwu5JPzfytv8+U/VzVV1IKuJnNFERt2I95VQaClw0Z4PetaVeFjoo0Ah
IoV/GVjTfruSgZdVk3z1YRMjosvVRuNfusH1gUPUa/azDN66b0f0IkeJaqBHOCwi
ILXlOCO4TgHYcbSHqoij/OZ9UOfOEvtXg0Zg8HiQD2GcYo8MaZ58OjOS7Thci3yP
KyK2NV7D8R2PvW3QV15mwDNfnwZMe07J9+k6jksYLzp6c/bC3CeUw14h19jN2a6/
/IRlYxbXA2lM+3aCW7/jb4FQPh7g/RWfk96Fw77qm9IiLYRmlUNbjCua8MSYkoUu
Cl/6wMLAwWBth0N2VoRby+/JAdxznNGnKiBNY1k1Lg6sxtlX7UUdVX5KlBOm9nCh
55TMLzSyE3ATK3BNtsj3ovJbMKmXOMWXufnLx8pdXuxJKRF5vSVyT0qEtG5jR4qQ
2GOTnzC/EvydBvte5xFpXMOSVyrf5fplCh/KMVQRLgwJBBzWJj5U1V2xKd8bWJBJ
yxD4SiqFDcALQfaJWQXj6+uEnFrgNtfURU7p82k1zfFIUfbU9HGAZTtRFrCLhB7p
3VZ2wkNFVR/N3oZsVSTSoD2rfNvpTdPRVbDDbcwzT9ughkyju0lbyBWtwJJ4LUtM
HzksuTvpmElHW7wc7g2jH4N6eFwXOfkhsrN3PP9uSSytHm3+U1rZSuXTpml91k2u
4um6e+bYdzEDD9PPDodd3+sbXCI3wfEya8J4VzHSaBpZ8/jcknz84jqu7rQHyPMH
nY4aIEa+EovW1r+olJo94A==
`protect END_PROTECTED
