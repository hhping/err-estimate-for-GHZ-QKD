`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7Ap03WU7/knt9+1IQ+exW77FZgqGuYtJFV/CRxM+g+/atzKaubgPvr1EoLbUpJM
gTRWxX6khYg5O4Ka/HwocnCKuKhJdi7oZiuZAiibPzu/Vj2K3M95BwWj0Oc7tiuU
hecmkPoFSkjF3T7VfUO36lIAEHPsnlfP3Dwc0XiinrWG4S0MTQ0oviPJ4Tzj05FZ
n2f3BwlP6PBZLFkyCZZMKRrZi7m3YDQGJWdjtndL0+cweHWLpbCVK+wQIdel3WzX
MiXY5vZZUfU3RQI00L85rpZfG5S8NJUzw3U7BXRDCaqPglF6WkOBUA5Ke3+8OlG/
itZeFFMtxqt2XRt/NMEwyhT4s+eLTnXyWz+0uHmnULtl3acSvA0I+ylhZjJwtKN3
Q9FpJTrQCCwPCDiHgfv4iu4BsXyvxl3MLLhmF00Z1IkprxxDy5zqBlS1nyJqH1B3
KKzLAuTWNOJuqMS5/Yv9JZguYa0JomSbZTLhtTcCpjXCOmsjIIn1fWER5dPR/6jR
`protect END_PROTECTED
