`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DPNYdv2DV/4Bt5K05xs8WMkP7PfhnYSLnv1o6r5g1ypuOQDyLuYYM3gIeA0H03Fo
meJg9Ez2nbaH89d+TgCIw1edfww1XkHPqNBpMTEBDFNlixsFLsYlb8WtLkgfnHys
WE8sZyUoWb/vBsQr/eFu7ZmaIl+UIgzFDHrs90jpNDdcFWZysQWa2Pq4FAllyFNn
wknbhd2CilbSV0UVwtR9LqOCPmAkHMTCjQd0CIsyLQ5bBGMjRe5LPywjeaBZ3iOJ
Bm9pvpuoITDtAfq9bwRPQD/F16TpotUb5oK+eTCQT6CfWQQnuppg/7sLvjWMypfq
HBxuDA2qkaRWlVGVEZGDOdBFuuhaQi85CSENxuiCD1cCjSXblQsAouFjFq22tqfr
FV+GRnuidwqOXudBOOc3Plbi+WFUnBRf6mCzp+hLm+wnwNaT3a0Gd5zJFBR8hZyR
FzFIbzYkWAqjGH3oq7M1r76jCaYfjlc8c9RR5Eo4BsumTZ+53nXsd5j76rVtnOyk
0BR2pOyjrubXb1U1ArJ4vOlkA20h9v0hKG2Kzv7mgbaar7VgKtV00qva7A+DdlBy
4EqA9fwlXJQtIHsHZsgWtDkouu7J/Uq0LGvYZorVcTkegLoyKgAiYNUyjvfNxr1h
4LAZiH0wPALcBuDmHuyzfA==
`protect END_PROTECTED
