`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHtbt6GcsWVkKqBE0QybJ1N7Ta2BQIuSfVNKtcWNgxz7/waeTnWTU9BCVCx6NA8f
b0qLx6HgLv0vvC2doAEPaGSTKXvNe2IC6fNFAFFomTRr66k73Hl/mlKFHMTXWbj/
j7IofN6LYwKQohcQs2752fQ7bcTfvFqfLQ44KXQ3MxjF3Miwjg5XDWE+VMB+YT6o
vhJceEQza485PkrQCbgcZDqdA3Nz6PBldjNaVasMqSlnnzKbJlQtOV4tJsnGi52t
s/MCvMJ5vpIce13f3zoFGPhRGxDuGvjnH+35OIn3xJWTCmN2jxm4UDzUrlmtBoe2
A03hev+wKMHFyOgYiTpIxI+qbiNuAdZ11SJ2z9AzReo5PWgJ2Is7wJEZDmoqbhU/
/YU4ZQxBcuBzIffWX0PPasMF1/xJ2w3IEbqLrZVhEKO47o3ug7CGxlUJg6PMupob
aDCQWtwAjk//yt2I+9JjlICdgk7OuTR0T1M0zd2Yy2eWdHBHf3TVXJ5oGAYjMSVq
ECfpxUO/LqKHLCx2qPbMwXmQ9LQ3MkKo8jwcgSQ86XgBhBRl3aQ+tsnpjI0LVwoZ
j5B0HehSBg11CD/EQ1AKiitX+lCElTH/2tpbLlYefN3rN+vHP7he5yMFFrz1Hwk3
O94ugkxXa7l0qSr56GlkVtqzLfuzsNz03mjk9ayNJhi1eINQM9KbqV39sni6ojmA
k1DpwK2CvXHSt6opuiugm3zKgeW0a3rselF3h4ERV9+lL+QzfiGv40SV0pVlF9Kk
q+IDnyHBC+R9fwc0ZupcGjmqRm5frAN72xpD1ENzVx3M/L5/q/sDPOwMNYpmic7n
m7jeBRrgqFvlIyk8x0jnhStDY9bqKxRZkTuJM80dEN9/pWexhuhmks6jnjjZcDME
06GMJAWQ6id5hYy1Y1eEObFow1LtinoK6zj+o2EcEyMZIxXsLrE73u7aIW8q4AN5
xi7fvFS893RvnxMLgvEPcNQd4W0fM+Afrcn+wZIO3Po3gUrCSzhjjaQHglXqaD/Q
CtFeIMZIbH+/9PXNNgP33PIknK48GZKHNaAE2uhyBsmV7ot5DWP/b8jBESwq0g3S
AXtov1MU0Ni/zva11gdrzpl6+4INh3jjhdvrAr3jFuFaEAVENzZP5rlndLBCVBZR
kCAaB9kJo+89v6KzcZsOE/a4+xztbeVxg3RP8KOOWAhaBZHBmN6K2JMfzG817pMA
Yr/RNPcI7Ax4I5ZtPgp5fT6lfWTmdcL8Bu5e0WTeAiOvSuDj5bGZeGQOttmsJCbc
4XVrFReTRjwKpVhP2Acd2pUjjs2mEz/MmnSHSNd25rbTvuhT62LH9ha2g6/GHZfG
MebYKu/4RMjSpE7XV/eDit3PXeAgXaRSYOhnd3OH2eO/xcOMVCzhTyYsrNp7ue4a
SWg5RaKQb6k97W8FHjnXLBgxhnFJAE48EHojeHaeYNwVU6/v/iNZ8Uqci/wJW+tC
frVnALoa9nK/9F7rEjSSQxDg3XamKKsGvramX8bCrfM5ovTjekTRIxDvkZCtglA+
jxoMN0SPxoMwWhOUH5iF9NEy+Lm8G55DegKK/OHDUQv/Js6rxjOxTLXVT97ykdah
81E/IfLQXZyP9TgNfyFJQNZ+pcXkEhlT4VP2/BcQxd43uiB1VGSeMdhG44JUEhE5
cIKo2Xm3ntHvTzVomQEVgTBpvByv3Js7BmpOwW1PHgHkcS+44HmoBlAGJySA/cE9
IhVVdJL/4hSKIDvPAwu5X+KfhAkR1ePjT0ZW6K0rReVk1EEaxKPn+refISQWD6qi
JDPUKoi+oirbcyzMaqlc8LZsazxrwy9i5Qhzm2yrH7+l53LNhqJMs/KhDJEPc998
LeXV26UAqpJ1rFwsS1GOEg==
`protect END_PROTECTED
