`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxJOONMWL7xBBUr18O/kMOj5RGa/EIv92xgEL/ujGO3tskbl6QZFEGpeBSI6P3p4
BoxeyCxSwdubITssOGlmyl3FW+9uK9PpBuWXgHhjBghlS2/b3bDhMkml7mOT5NiD
FoZL3ueLHQogr/B9DgaWArElQ0pDfarDlbzx++qApPMkEGYJUNBzCOCjQwTKROMO
gaSMPMAZUlHI7RlBeJZKXlBWVsu4MT48sbNL2/NMzcQ59Y/0cOxhOiU6vREFfQDT
5RhiqBWEJyRm69ywvTb7s4LXjUnK4nmQTfgahpQA0v2HOfxQmmMotdmK+15HoE/m
Ktv4BVqdgWlcliKkkNgcUy5s1ItKfN3WCI6/NKfKyJ5CcUSoMA9r5gEzXS+6TwfA
REhT+7TEDygxnoMB3BS+o+HzHOMQ03mhjQU23bADaDaGTZkwwZWouRzf7O5klrES
zBV9jP6xA/sKkbQNDahAc5OUJd3c6IPNljiYk0tUBOXiY0+Fvwi+g3uV6/Fvy0A0
lHyt5e0iw5ceZVxSgN4MW3dUOEM64mCfGGe5QhjqaTj0ODiwIXOjCVyb+90KfU4c
/fp9XLei0O1x2tsZfAIaYB8MaH4O7H7j7R/cDjPPB5+e0L4szz4vUc3L5eD+P+IU
lQXOxNof8hHAEfm85xQxtiV8vLQG8sgyfNjMb24KW3LtXrsVE7F3vX0XH33Rnluo
ivQt+4TG45S8v06KvZezAJ/DK5fd78VUxYo0Tsrd+rjiNJEeP4HjvOiusDcFqxSv
lUlpQ5J4MANrzsDYasmB9PNoKtS3fL5iUIlAW6yO5Ir/gyllpjmYOf00qsv/p72L
pjsNA9CxnwldaTscAEavfUFS5uRoMoYgACxRYy8Oskw1LIRnfLa1HTP3OThdY23J
aDG2bz3tzmvTl4eTSp+gFCYLP/Tu505/mwuvvx60et2zHfpq+CaWdwm+opQasBsi
14PMRaMc5Y+eC8C4+pjRYYF72CZOnn+89vINgZLq9AyxvzP5SPBwZYn/eFDA35O0
5ou5axkraPymoQlw9ZAZC9MGtRiRgYbmUPuDTU64td4Nhp65GBR2qwdfW5HEuuSL
QMlMJv/fgn38xA+jxdOBTHrgFCOfQjiEcavbt10h6elmoB7Hnsr3QjHQYOaPcjSu
dgjFJwER8xUPjr57ebIj3+YNcSoC4f5FHd6UJ4xSx85cTuHA6euMSNddZJJOpy8t
prabRZjHHOPNe8MfKI+n8kLtujdV/jpFYL+yBWfZzcD5dJPeKXxQWiemF+76W4CS
3Z+fQtLxVQRzSPlFxrm9iz+XQvf4d66tNcXbiD6dTsaO7GhkwXoGnDe4x2+GdGGi
LpOMbJ0eI+HjP1gGFORJ182ms6xC4wmFTvAT0CD7KMMTk04niGEZsUjuTmdk2Sm4
AJMAsiNm6/jqYMOfMXDCZ5ylLHoWYz19NScWeX04m5ruvUZcb6NIlzBYeogMLL/o
Tj8m4kudCJr1cqPo/bYQBStsL+GiyTiG/gCh4F32IXa5Xbe6vRaHx4vBSShUcELR
5R/w9pKXiLCnejyGVfh758U5bDls8xFijqFLZDvjWnE6bAC6iG8gYgVEkICoprwC
xI/h4JLNE/ht03PLZbO2ZRdF6c1j49rDeOOjDaKzCY9G1ybp6vFJQxBoTMGCDwkg
1IBh7IWoOvK0/9hv5br4KBldC9NZDOGEKYt8jCoyGCILhJEUXvfs/lpO9vKDRaH4
9BknYdHNz3VVuvelyLZHApvHGoz06iqCZdzbqq0uAOUmHPJasqvJTp0SMq0s0ajN
KzpZ+dsnmfWUo5mL0qao8Gax7+vbWjI8nNDsLnDVeFXRAa64UuteY8f/ilcufr1v
U6A+2A8laAxQXA2TwUfERy8XfPTTROnTUZnKLC285btf6f5jvKxN4lEGsMIqV9TY
b6RmIfqk/RDT0SgNco9rxAWOiMn1HeP6d9ogh62cDGmS5/hnJf5bxMqLW2uN2j/S
nI0AYJRko4XCeyGRjkAEyjngxSeTDQqAPoXceyYd+ONI4Q0ns7VdFiQ38DPWUX4u
vjxCyZSAVdUOxayzukE2JEPhZfe7eDMbOvphVlDRQBlgeceyfvXjkbQzZWKDxWTw
RsS5bE7yFphIdr/+pK/XuuLwxS5aF7AeW9O6kXcYSC06OwTlvA+eXT8DFij6fIed
4T1Mb9EODJN+b4E3JBGmc/6cRMr/AamGWeNoXUy20DjuHEcZJuhNRbyfGNwhDIgg
cfDxSaeEx+A9uvcKjYhya4NHza0Qf7CqHmJFu4j5AKI3H54UjlVfww1ftQBTC07J
xs++gABKXEoFjGdBkAIFIV0ymVzA9rq0Iy3tuPCu1PkbjAKeAydBENDeXxX2X64n
kurmXaBmoNzHkHQEVJArbbz0dTzZd+lFoYQH6flar8IvF5VuR6yYFQf/S6OmMeLO
LWgm7qmbWrqOwkb1AwfZxyDEaYJ2Lg1dHhAVhEmUmnPSH+Be6WqIcNT6keKhiSb1
WMUfRk+A3N5MN+cJIEqB1/0Opo41/A4QdQ1yPKttmFzE0/ol80AQGuqBxstq4nlL
2X1cFABf+mjKsdGheui4rQZ+r8Rx2yqCiRUSqoibIXynwf9AvQy1mZcFbIu4TCR1
GFz/ijhXOYjJNhfRery8oaLycpNHq0fC4aVzlOBbK7dGgBhrXwdHRRbjWlXPi11v
BB6nx/0hlT/CA5MjCZXe/3WVR6ZLrM1DrVMp02IYwmMuARgNL8OasgMLykO+5kqD
IMsD7RecgoOMTgwlmGaSHwASa8jvg8raq/w/fZTDK6b4WxKmeQ8MPgel4abVP8y3
dVwniah4AtreKl6dX4xaB/SGfZv4abeZva3PEw8Tp8rCd6shdih/4kA6YmCYtaDQ
KpDTqZRL4SDpEW+PbyWLohz/fb5HL8aQkIud++nFdbc=
`protect END_PROTECTED
