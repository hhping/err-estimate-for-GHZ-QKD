`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7rstmeatpnKFcmDDDwoQkgmZCs8fq062/mMQbBUhUdet3DjKSCLcMmyfWm9xVgj
Oq+AXbqBfhTK9jgeuOtDyuV4Vq8tDDkkJvbnc6tSpFz9oJ1jkmzWOorD9aPfcygV
846kC9P2WM2v5QESOTpmaaeAP58IVf59ReG4gNPenM+o8ZdFFkqMluF6EZJdr00m
pAuqwbOBOWnCddpzMicLFZqtXmFM94M7933EHlnKYtaqPLW2oZBsAP1djsTe+Dge
7ujK+XsURVDv/bon5TN6AH0bp5UOoBMImhngIuqYqmHE7RLeyH0BcZgWOCh2lfKl
R40zHYSDf+7SGObvmcx8ARkomt9pf/yVnicj2Kmwh2vpzUMqV5KLMO2VhZqfOYK+
iI+yet+QPRLiKrB8/d40NzACEKewOVH5TaZTHTJS35TEwV5MvdBulhNblmhgFmiM
5NEZRZI8QKazTxP3EZxr6V4TOa2EjSI3TrLlrEHlaTjZQRIWS0igUld/1Mio0+Ix
AKxyYk/Wy/4uKmcLA07TyYlwxejpiBcgGINdfo269tAgwRA4Kw8rai+Sax/KGbpc
F8MbzS2ZNvIvA7UdbXKO7mdUpgmwBZA/voS/PtIsPipmeWyO49X7TjK0L71Zx9W3
dmitDJ+vfavBYdA3tM25bFIPvrnjM5OuuOc3eVMBdDUI8U0gM9xkf6Spz036U8e6
ixPjJhn8+35poyxVwuKVwtRP+xMwqqmwZk+DIXij+YU0ggYiG5QPdVEyogmSjCuc
UTh1IXTJp99T7/R83zqPVBFnR/v2CTwNE7uBPsNlAPXsIfRRqL6vlfXHdfRdW1CI
Udzms30IWHRzfyQ5tjPdVrnt0rLC6fDGWkzhQUNSZqg1YY6OaqGGNnd0G1SRhzxk
E1qn4FKAPpYEMUXZ+lmUBvgX5bVabKfz/KsH4AjgNsiLJFAqA1NK+2+SNjYGGnZ5
TrZQR3NJRUW1lTxKaD5mpd3lv6fmRBcY9dpO6QiNoFCTSIlKCucxK9IAmbtPyexZ
3Qiq+fCe8/IcMhD8MKbFSCjVLaBorEpeEKr1Yg30LzUq4E4Xww85xAXVfzChMRK5
to/HR9Ots5KX7+3dR8A5wHimC5CbQ38bLa8o3MM8p/4wNnVMHTvFHjttyWOWAYjL
MdU9cfAk9PZAYjH8RD9Lr2PYJeello+jpZfO35BDzInfO+GlOpc25CUwwHGJAmQa
RIyX4K6ci8ANrnsNbSIYS+6jmlllQzf1LwyIN5oMbdL5jaCfRrxAK+09J5hkIwr4
oxIsGQhcHE1hY/gQNe7yl+8181GdmhfZhWe+k+CpeMD+2JuBCieRc8zIi5TzHPsE
5PEm1O2A+jK8EJmHTLN4+UU60yR7lgNSSnmocCGf4hqFrPqAbg/qm2QhquYYvwO9
vqK6RhP42PqPHFOscFX9W6eWaoX4yTXRBU9anf283498bHuUh6piK06WWCZuW67V
8KZ0ykHCoPm0K/15itjkSQ==
`protect END_PROTECTED
