`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dbDLd+8KOCtQWY1Xwdc6BHMLDC+/Phc7VfwtCg2QT26KAkpQGuVZqbEYFSG4WPlK
qDvCDs7YCtauHwJwJ4Ft4h8Noe/Zh3qVjX+MGcpbip2ZeW+pGxcJzW7i6YF3E9WS
rR480IPq6DlNu1nsNqmfRFF4jEpFSCmgVVt81A5TTxM9UbN5zklpO4rbvWiuf5MY
9fPkukkwtw368+Rz7WoNWU9d+o9kfYaqn6ao4feJJ02sks9kB7MBv9PF3bEdDxS1
+5oHx3ALz43q4e+ENeQ8MYoj+wskqWGcS8qSbDkqnYAGnSOdpLiBooNBppS1U8xu
4zx3YmKL/ddA5of9G1mGC0+vi+dbeP2wePUS3XSiooUUAv+kK/AE7eYoAYNzt2MV
7eotZuLjC21Y0zCQ13omj0d7wHcZm1XXQaiwqnnGetQAzo0ZCXbwSXdKuV+Kbesf
ds+Coyyggd1Z5ceEIK8AL0bwzTD0RbcZofG5eRyE5dzuWIvTqoUBNip7/lhbC4TY
0scx+kmglnkqbmMZg7XoNUyIMjTqdzKFslqWtO3+PyXFjueNgkCBOb34LycfU3QP
qbv3dTRywXuJbpr6YVCKLX38JfkRqxnSqkY6rUsGt7c5CvqQo/0FoW2JA3lsSLYw
oIFC3hNXnytpqIGAipichS/zR02fqWoAMi1bTXDarWfT5TiyQuiO8x0ptn41R1pc
5qfijbYkWgXiMR0JcsdalmQ8DsFFXf6Tao+nguTu2giQiFER1ULPmGHH9s5EuwYs
hWNTEie6M28cR7bfpJKbMPRzLAInA9i/jm89qh/gliJL6Tgg3XRoCo5ApDbBDsen
JbdHwIMAW2rFv1W4ArVbh87lkKnO0RkW4QeOpBf510r6YkAN1PkFXnNcl6SgmKuS
sqbg3H/L9xDFpCdWMGB7pestJT/FdKYNZTbf3I3oOSOGkY8nyYl0o0YhlsV4TD3O
gJUovz/1xhluo3GJxvznT02bbJZgLcEhBmOTd0YMrEdLhn9+CiDaCkv/yA4m2U+n
QdofiHcq1JLDdnacTHy1BO90ZzHH3ZvQH/NrkwJb8NNv0OGF+sd4Wws5/g2oF3QR
8ft4UPXTLw8bqZ8YZKthveXyMayXbXnDutnIYHf+THbN1WPySlDt2EodjL+1uz1y
Y+T5kBSJTHKr4BdEZ29lW6PHpfZHJ7zzrrAAyE9IfVkDkEsylFTWUNn1B3J4NDRj
0j/YSk4aoTOUT32LNLpjLZtCNqtkrh9t2ikFRMtciS1FoKCeqKWCg4+NaH3SLYu9
hHP3naZrxtm+0rgG/5+O6Ztd+790361zqngz+6r1HpkUNWDZwwTzuIxNYVAsC23Z
4EiRDnLCAc2w2l0CBu4oA6mu8xErWxYql4FLwBeqiwTSQRbFgb+olAH7C5pCrKtE
juf5pk4OTkZtlmhQLjfjVQAH/pFHNAK80AKRnbUoAst2NxQ0JBo6ddfJApHvXHCe
AMbdlZ8YudI8p5NOooHmvzSU0HI9oUbOdI6WHFSKAe4FRVbHd2FyG9SbQb55px2G
hGFTY2TFjN3AIYfLSqcNhrfmzLeSekYOfNsZi0B+oKFO8HsGVbmFoRF+BMA7moCW
3QpW75vB/bQOV1LCT0fyCsTJhlV+9vhe/dwu1nTGdk4zHL1qB78bL3YluxmKCFwj
o9DFVA6Az3rUWPxfXAjtbJr/lZIxv1Rg1yCBO00io3R7ykvpD2hFDRAsaD1ZZsXV
QnWClAGcA+9oCEHpMjpQ/UrG9/fUArOMQ3cT0PsVxp6ifoBdupgfEckrFYme9G2J
8XIcvTwSo87FUdueRql2grfFJwBmQIYrAzkGpa7oaSHbXzKbrB1uiXsaYKtekCIC
s+v0JEAq+Vs9MXqvE998Yof4bRsvm6XStqogUJrbqvuopIJmK6yx671gIUj9FXzW
8s8fq3pGDYmWM+RuvJ4jtKpE7M4pdEbtwFYPSh0+RdKUxstq23eFZaWUGr7lr+Pt
4nHDeC1oEqYWLf4gy4KzrDZLxh/MLX9Zj5cOyyOd56WOtdImzzC76A+fjov3mEFW
5eg4TWyPmrh5bNv0iP+aMpehf21a2e+F4NzTTctz/9eTwQRb73VMvTBhiRw0NJnS
q+G/KhQQMqwqCtiUB4qqXYawuiSkY0C3oz37fGckaxCMlymVolsJ3D7fm+To+N1W
J25ho4ctU+h7TdJHZlkSkQ0X4RuMT/2gnOVe86Fa+8hGXFc1PJ3HM16lajSu5OFc
13rbIS5Y/Lpu/yFOWMaksy1o3WSwaQ8d4wa9k1DhtyfYBxd90x0C9BnI3/HXHQtN
ilOgtSF5N/VkSr0tCAValoM/MF54Vafcmr2R8voxBPu8QXFaoZUpWlL9YC9QJfba
okmrvYm7hx4UwCgPSnWSwb73lJTPj5ep5yujmRhy7v8PBbhR0cC6zmarGnl95396
GseJacNWnI4hIYdYuZxywUnDjVIrCxZ3K7yCvNJd26r/Qx2dmZV15LO2cO2yCtLJ
pvsu/Cjjlk6ftZHT3WQu9M1ngvn/VhpVe4/M+4M9SUy9wR99GvyA/Kj9h1CsOmo9
rcgCf13T/Ggsh9TCCdrmRXWxYh/2ntOgj3cYj56tn8sYmGBSDt1sg3L589/hrkVJ
ZLdwn0JCBpXc4QJ/EHXVDeGOPzRpP+w2wAKsEkXhq+YcgbgFSzdXZ2dvYmh4sKRs
pnJicvhz5ZOtrNF0Xq+i0vrrBbrYyc5Oc1LF4Jd5m2klo07HTnGstq4PjPLt78Ts
APxspyq55knlLnjSL4Do4bxZABhWJ/ESFGHcyMsPnhQBTzvIDnPhh4CDn4le8Gjf
mFWj1WY9q4Nfq6nS85Qhh3oGs6S9i6VTQZ3N/P2CT5j0Ut0wEArbfm89a2Q11MoU
sS3Oloy2CqRe4TnIcCiO97yq9t9vPRRjesr//LvZ0eSy8nsQ1jSNh+35BMxtPxGo
BWTAGGArQe2PWGEFL+4XyfVQF1Hy+W0A6bJjkGRabea6oebMkFRYcX41Ww6Wo+nz
37q1Sa+JKkiWq5MIz+K8kwZ5tw8+3EMnYZdq0v0788yHrk6V7ZUve4Yt2kYGodN+
IVWwYkJQ+P23BnJZy9sw+2z5TmOvqJ3+O4LqNCH5XjWsCP9+ky7lPyxwTCGYHHIp
i4E4vs5NflFxN+uggjkAB31Wq1aelIUU1uMJHBFc2D2wBJa8FjcqRaGK4RFhQd+x
KMaqggNYZvFcq+WUq7SrRXzXLb+cF4qzyGf1e5CG8fLWB91jT3eFnw+hT9rDK7Ck
7bKK6N67JhH6cYVVBL76q9IjCZtISwGa76PYYaW0xnM8kh/hXlZU1lwasM2Va/2d
my88oFU9StODx5C9QhfLvuWy8A+htWA5U51jx8xdbFHGOsf22ZsL+cdo5cmCmSuk
2KSwuXhozi4OtgX+vydRtiamMMzaRjP/TorDhbVcebX3UrqMr79RInM6FyBqhBD6
zw2I1MkzpHVWQwsNPyrEZxkQVxsTJ1fawaft9LjyztsO5hfMxfzPKIzxnEYmO72D
DK+EnpW6IEtTe4h6gi5ebvsjcBv70s9SPZdPv05lh2IRMPTP0SSuPg5ekCbTTIAX
pfBezoZ1ca/RxXXndop2tO119NicCgFAxmRv2Q/PH33udUYRS8UmSmF1oYN2srS3
6zg5IRx3sndjk1gUCKWhR+Bqfyy45xe9+cfbRzZEJpsBSfEozx2F6P2isAILdHgo
O04VaHCSAyaefTsd3OgxdFATyP5HNrsuA2WwVSHY5N/FbCAWK92uzRdT+LW9VsAs
oDJcXwHMuAGrdbEQje34nvLLaEsW/r9SkTFC572OAMSkHIetnTvOmBj2Lj8fgOPu
SMZTmyAyPV+N1aFCoJnsp3/j376HJ/dKoH5x4z4CV6Wez12OFgaLbV8OBRG2ETGa
uAnkdW3wBX3rYsqBKccZaTYYoUffA+cbS/iF6gF11Q+kBXjcuYylpXZapf5UigfJ
DsHyZxJSb1MfjGn2xRcIGFTaxBeBvI2RQz4yPEMmgiTMKwdraSx0kUNJgy7A/hUy
MJTM38nnQMUHYtJmn1Y1r4+aoizzKN0b+mQgOCEUd6QLaMZYuGjr4z84pDRIIc6K
ovYvWULjYHHOWYwE0SCyPrzWf5y5fQddilnJsHhM0fa8O8JT+cr0gLsAXpmdJyam
n9AbxnEq4nhIIr0LwzCRjl68Axi4mI8cgdr2hrNo+nLBh69SqoWN9LshAxiZAL8F
/QO+T1pYWk3rQ+M/JOy+a56VwCqFYVL+JAzTSjmEnAwErXIYYi8bscvZwCadDsBs
9gmX7FnJk1VK2GNxKUe4BmJS7fzowYiBY9SdwutO2YQ144pv1VefmeMv1QLhy5Ig
1x6duPOaJTfoscmH0nhdXS8UnFe7jUlnhRytTnMBt8QeHG+6DXARqpdHkoZkIa5s
KpkdR5Pp8Y5xc/qe0bNuvScsQHSsonBUNNmvttIeA2DReniIkIF4eLC2HpsMXslt
QmCjIAEbMdr3EbdHnSiyJgZ3XGPZFWGXrrluCkycZDBYP6xMXJqwgqSWHrtdD0/w
1CCs26G6lQBc96vkjvllMfr3DfojEASoFXlBuXoscqNQKwuCb+cIrLcjmx1DeVsK
eT710gKhRiIrr3uqXXxQJQ84CSkF3lAxtjQ50hY2CugSgT5h/ob2mGm5hrb3rJvA
ZmPrP2q9w1jNCpumdCececjikQTWnJe/OUCgzVSgelbnfGNDPZoEEZdXfSCuXxS6
iIrxJoE+2UYrJ89ERt0MGo/GZYaUAk4GGjbkDHjIC54+O/BdbBbQS5TDhSuUajzR
6BOYu/R9bWhrllTekvk5quapPS6cmRGIJXuAREtnGJ4kvEOn1eTofmL4ndvdXpv6
5T34MJelw1gOEhlAE1I6agVj2erA/EHooDIv+MCOmvkzvsv/rauAZBGQxJ1d89lc
b9lEq/RjUE8DBQWn849so6koTrVjpg6soZOrd+JhM7ysJXetUNo/rY28ACp/ycNN
wNaog6Kf7rfO+E8PdrrO1oBKVBRRHP+AXgxvQDlYQyVGDmt5dcmauYFcuptphlQ1
/3hfQPf0ZYvdrT8wl1x+bftuDSYBjG83YZzZSekDRM8nek/mZDyQjxPkwB0QAJIm
dz2luywI9RcbBY0eKqVupgnn83c4DzUuSE2+URnvvKWnAPMOVD4Oge0EJb0W1b4c
KB0+fYx/zLdcOlla3yryoXIpxZvvE+hrDF/qgk8puofaX9afwy36irGe3pzr0VG5
vtnmJvGwOZyImQIUdZaolLiYkm8Fu14RGDc4UEDObfCf6G4yy9jfpwJMfx9qbR9g
ftV9mC0+LiA5I3D0akE1/GWsww38ohtvPIkeqYb2NWaF4FBQO920kTT+v/K7AZng
tWCPL+Xv2l9lKV77hVVZSfEI1fz+JsclnriBTwX9U3Rx7+JwIlgq10VMK+iBLGY7
chCGe/sO0QvYveNSu8nldbOyo7/kr1w+8WVZQ8+htHmd865RikZyJnuAoyqH3egU
IiMDM7j0tFFqKchFiX94z2ozVwA14Uos65qvP+gUpwBZpODWOzI7qFmJinnl57DJ
21XOdqTwWvm5Src+3lOuXZx5dbtjVljfTxmPINWOXoT3OEoIBEkBU8bZr+F3/14v
6BkL8QGPzmoXHJK/NcNj6vJd3LTXi9GHRPWEr59neurncHTGXF641sA/uSG0PmoZ
yKU4C39OWe36ZgNue5ZcL3ol3/Cu9UCNDdcnVYNuIx7/VxetG2Vho0OfZSL4CdNd
apWgqRxp5n24StQ1XllF5B3KM42iq6bCu7PtQYCLqzrHpW2NctiSNGaqYXiSAZcm
cNlZgiA4Dxn9tddVxBIA9VLSo958tuHDPSxUKmgwru+39VoULzsJq34u6urQbRqk
sxj3dwevv2+J58TfUK+SPLcXGuCuP0e2L9tu1Hmo5S8YHiF42Ddi+pXYfTLacSIE
SfPWkS9QRLuHkHlXxjnbNn1OP1e//t0y1XC1XlI4iffvJFe0nmNOixvo6NNPqsij
lg+b9rWB/PyPJ4Xx1Aj15GE+YIfFI9KBGooZQPdW0b0TJSYLfwxkZNEJvzYjsHAv
mGBNsSxPQRS33SafURBwQtFGt+Khipj5HXPzvRO3cMksliw25zE5+PmU9ZMam2YS
5yDQahaYrPcSiwiQOJa5InKNALZWgMMlBzrjiqHb8wxpKAEQe6ONzivwj7UVBuHF
klqpAH39tlsYpxJd4WrPfhpWVQq/U5oHke8ONp4HY3h2Ifuty2sOSB4NPdwroeBy
GqsVmNohTyxrOCQ1nrcPVW8o22pG5WJHWTeFrDg3iNm5RNj4UpPWqvafVOwTwIfG
39UR0A+a+ETm5wwkictODOUX84fcem3D+q5m+HMKfnOOc/G+pqP4npd2WDG6JhSC
gG4Z2NkRuYPuq0Kr3ttyXkgONoJEDwaAKLeMyfXn/PX4r4iYph5QXkARHJMCz4ia
ID0EX52ybWf3ib1dE3xveQDrP8t7BIIR2jYwXRgRNzHJeSqg2GeTn8FuyKYS99FI
ldboTkvb38jKsTVjftLWgHIrxyfxC4JcfN9uulSA8ewB92DSphHEcxYHMHuIv6nl
I8ywWjU7lSkoixNHdSpEJxmY1dz7cw+NaE5Kcn9rPhw6APGpKftFXnt3ndxha+hF
ub9h+zxOq8AVngCFXoP9DiEP1ums8FPw7J2MntZ//BWpuzRh1pxkh7EB5WOyUA34
po4CS7MU9w0H6mOfMmuD+4tOT3rLsKI2a/pX7wo8OlMEcyDI+yCcuUaHKti82VHX
7Hdj2f4+8clrrlTkJMjGpXh3tWwYswgRmvCZdCY/bqSrrR6EpmkQoMMtlp+kjFJz
PMJFZuVYcsxGEEdVLFWCSaAbePJKEOen3A7OT2NzQf8cmu89L+gW4FCk0eL6CkLq
eewq91IZXD80mMPAWg0i/ysawVKqWi9uQVuPlygzgccbJUiVOwv5Yl8BD3hWLgyY
9WGxCbRXdGvTnYqaFgk662UoGS6EynZGNuKqZ+vGZ61NirZV3OMPLfcdoR7QfyaW
jnrj/ZPGmXbSTalNqqJ0+iKKj+M2TPYmpyl8b7HxOOckANS88YDU0Z/a87KjGV6M
93mT6nuMbMwm0ojYeDnyz6xCUT2vEHtNfpC5fTlFe8fs+z9rBAFpBVI4Td0yOCU3
9U7vhXURJh2riS1Np0cGwvRIaiuX/KvX1N3XhdayxSZUlSR9KbSj6o0QwnP2ghIa
P2wmEAyUL9tmoisWUjRTfi1dksrqJ0joj4nPR+fIKLHeSNoBTEGI1XLxrssKTlLT
xMHlDF/ubDL46/J5dde9wpY/au0738IAuOceIp8pQ2DJVBb6ZFEoocywnf8PzurI
onVbB646JTM7Pd0PsHUU9ScU/VuvaYsDA35uhi3H8rZNVb8mturiq4GI2bdFbyo4
0YGCyf1wIY0B+xlmHakgjpgoq/d6+R66FFY3sggTi3aeXOy/Hlg+0rbO3RMFyd6P
+aletvhSZsOeBKaKAPp1P00QezH/w5WfDt5ZSLj13T9QfT4X2LzMpBMHa87jxHeM
cp6tfWpy73Poyc7gj5Jo2f1HoLsZpkaLET2YzpmcNLE0LxJMWHXvb+nIm5LXT4ga
dKUmsKDMkH9MmL91Y4YZkNEMBbSsZJxgq4qM8XgBnnhB1AsXXGWBblARtg6EDVli
oStiPHtIzn+2OzIf7WpK19WmLCtNqTOej446JizZES/tTZg9wvNZ4Rc6c+CBtNvE
0Vy+gdL4gly9MLbT8+LigafCqUfFhBwBWYglmAdhq5qP11httyx6suaC/Lzz0465
A1Ln+MDQYLOd49dmylZ5JkuYMGY3A6SDcXaOw0bOyOgl2yPe5DF4iJGMuate/Hks
YcE6x2+yGQ1DsTwjg67GIM5DxryqEqEdENep3ZXOvn4KP2Wxu7lK2bp76AdvpInE
5ZdOSKjY8T57HYOPG0fwPXx9whEtoS4yb3GGKj9phMFmKfClCoTotWMTfws6QmiG
WzGQmLzvJVJA+ShbbyAo2/QwhD50V/qzqGRbb+h4QUsDPuPgHW4hkrIJBTxysP6Z
mBRMVFJFsAJSgJnQkkZc+b2BqJNCU2WvZO0UdP/szOCgcOCNNK/iHDVVrFwdwgyM
G7SuUyxSbLsmFj7gYVLKc/wnZqwEVHb+uPvt4SKcNoFUyxhTH7Zf7xGfpL8s5PwV
Bsqwm7lYLL3ZOelaEUmgtkCmbtIG9dBi+vyiJBcRfdN9liwULEsCV9Z6OUaYo6jB
4Hd4Kko5kY5MxGToCSnteJMDWu4gawAqv8d9nQCjGrCyq05OyXbEfs6xQ6aSzNOs
OTX15Kj7QGqaRroHcZbFU5qAPPcb60S1sfHIpvNXxMIYdWCLsf+g0qX41248shkl
8n+MrFp/oTxqWoV6vSLO8NbEtIjplMWM1WUhn+Nj3r8zU5/k6zBOYdM99GXds7Yp
dHZc4IjUuCSroE6zOaJ9mvwlh+bSS9SLiYlZ4JjCZp8WqcRCGe4QJYaY89VR4MwY
+GdSQDx3B+vpJxcy7r+L8ohAdAv7Ettd+eWsxIeEGsdaTb9atuXbvxFvbhx1jODF
OQEZzJxgqzVV9CeepWLOL6leqt28Od7igfwtJjStol4ajJ2sIi0l7ykzLLKQwWuP
cXk7tfLXmpRj7LZNOfCdDBajAXTvuBOg/bdxJ9luCcX/PPjhikZTMQ1uTnz4rdtv
I/nM8tWijSnIPdvhobr+HEcpzV7Fxr03R/H5IUl+V2t5uuSbmCu+YokRcuYPTVPi
lxTQRXNymZ1J53VEAz6H71Hrf6bhXhs5U2VYGFlKe6LIbJSQupASRLTEiOeaznaH
yyxv/c1T+v3sAyKHO+FC8MvMOnVRPdQK2Jtve2r0/eWrP3OsWKfrOhzbGy4dOo5Z
nbnJy6Z0XOlPA7kP0GLeqH+5MZdjmTkSDL+JSxgua6c2TwGFE3rYgB6/NGST5BlM
FuMB3aDugdSXa8Yvlnk+Xb6keyUHrdJIw8Dp/erTGYnQIyaVfizGrduiyNuTzLzo
jFZy7pCsWmcm9aSbVGtho8u7ocPeYzKrTf5E5UKBo0GFNJLYozrnzM1da7hOsvSF
MpMwcxKpeQPHeNFMW/38lhI4qzRzev1wAghg5A7Z3SA9mwgrhU0aOPzQt0ZxGUhw
p8AP5nyIkTnvRysA9LZP6gdbL2XQjeCBUXWyf6afL13JpTBJomnqk+nsZm8FPPfw
AaQrZYa7/kTW2qPpCYG4ccdI+ze2kxEcjGPI0QakEaZdoBPYENQ5x3IAK1Ywby+b
3l/UAf34ptcxU0X6H5O1ad+tftSfm5VLlHK4EMUzp/xGIhvrd/aAsdrKJi70QHZk
A9vLNniYwKKocr/XwVcjG9jTEY6BtmPb0QBp8o5TgFhlmF1pSyUns/2MK8TXNlJ4
40I8qSrYuEBAF6IiyZrhQFedNr6naJD2zyAN7SrccghwKwV5ybS8rwoL/g1YxPCW
U4uFIDHikKdkV3BD/zcPpdWq9kTJu9FRLfXBvIJCScccNttp5mPUOhISuHTgVkpJ
cAkfeDFo5ZvoMFzljj/UTMf82QTgXF4vkqjTbbRt2FrvPH5Cg14WjuB8CxKIuek7
zVC1FPM/KwBU2YMiKjJoKFz4AoB06WXmB7PepVIL1gmpONuUzpMnxEuX4xzfuTEw
GRgiLiWXYYnUjQ7zD7UCNpu4ksZvnLOLIk2wRMnI1JqueRXEo2jJYcdroC3pcMfg
hrmHpzsUQh9o7TU+LyUspimJa27vZkvhfeeflbciky11Iq5mnGJQ4iGbX0FjUQ3J
GxkT53npwjXa0ifM7dRfq39uFiAuDQvO2rR+tmucgmapuPuatZV3AMGFULfyKVTj
GEba4vbNXXqB0zvaY2KSdUsaOPIPEOrrDXzyFv1HvcjA4SDZ+V/if80wIfgu+Fde
zVQ2cFE8CwTP8M2hch6Y5PfdE2/PKlhXixmcmCDKwATwYXr0DWXSpvD2EMUou1qa
LVkMpX26pUVGtk6zx4oQ9dKPFRPT3SGzSOVNotmOlPhUkoUqdv5MQ8E5+lZLa0Lb
mETSe5BOlBYlSVAZCk7cPJyDfhm/eewKY2N05KVajH1uxPDXbbNkHgMz+nJ2WgtR
K7cLEBeBt34C8WPHUDlzHfMy+CBYfiPywVrGs6TM43BRL073f/yjYQb4DpiydVAf
SXYGUzyCC8pa/MuJx+VNc/g5j1bAUc8b5xhHAKvDrJpcv09VVEn4hsCd1vAaL9RS
+N/U45dg1EHCxyMdzlFaIP528CtoYYtsT9psbWx6Y8iyYQebCyjXRl1uM8DtMv2J
+aCLSLHgrDgozt82tTELcOq8pFo8918ruw91bK+p94Zw3P6vxjJ96KMXM01592mF
Lt8EZifuw1fA+hSw8eJF1DcCgE+QdpgBQG3yxKYTRmMq5jwbTUmgJ9lOHdsbDlek
NcIm4VVj9X0myrcUkx0opkPoy91S0GWUs1LP932Bg67VthchLhCDJuv4FKDz2I+X
pkaXQedU+BqAGFvi8/JuSeFeTGPGaufMa1n5Q0OswABibbnRzkH7JPn46WrhYODj
09RF/tbwtYOnnOhLdY+X6qqcuJwwxg4wF4g3xbYoiMVXrJw/l6h3pw3n9LsxGLca
NlMQUoB6xv+eTub3RbIffzm/X+jz+nZX6B3yLuaj0wTV1T88iApd0GcZ3FGIT9Rc
ERv7weoxGwl4kA9tBAj6TlzZQZAE3ooG+R0+YomzUiwG0USrPu1iZZD8Mxpw0V0H
ZNOdLsOmt9fpKa6/Ovh39013PxDb4ojKnTVjP2PjJxjknxF/oIDndmt9ep5wlWz+
ZRFSldyWDP88OaNGaxhkp44RBO+gl2BHtddM/YfRCFuH2HYwb5HyNyFL9IRty3RE
6IgQ/ToGH7bKz8QyilwUjaaJ7qCgW/0tgsJt0zk1rEHhXRxJ4j9CGqzbo73zC2dP
9R51QluxsxKN2eoT+TYo3CqWJIGFVvUESce3EeThJ09D41j0b4tKZFIXEpQm7gcn
1uX7vtPqSKWSNiKbrHGQkP8x2usuD8yuYO6eQVLwhEK+7oMJtBsE+0vQCyaW2KyJ
UtMVI8PlHSNvIcDDi0tc7tAHVJxcRZXaldDck9op0apPca+rJs4WsQ1+m1hrQxQR
wMhtI3MBhCpWXvoTylJmlUll2Tl+OKSb3KImx/MXqDZYTh2xd808I0QWbjx20r5P
KmQho+vUYtDNs1og5N+e1hHUozoKCZMPkwihcxDu/IKQIeW4qiY52a8PnqgjPgeb
uKATBO+dbX6tPcidj/unmMo6YfvVflHm6zYlWmKBAHIhLmB6djtJoNzdoTKCtkzL
gpiNqQXeo3mVoZFOcKhMmfRt31C03tBaDxs8psZBM9nozB9eCZbNyqpzNMRM6+s6
/JNdg4gqCfgQxTPQ92MjBSmwTB/964Dhrxt0CJWbmSOzBNe4Dbxy914E0iw5e4gE
gsir4iezInd9GsV90z2bUhn/0XF2L9UBAdn7eku6RoKAiZLpIclkxvNdOmegwExL
jf7hi1PqwaMb2KFRAFFSWVs74puQHmuqqGTb2ENj4lE1aTfxyoWS7VMkwtd+E75j
qRA/Rp5/8SnNdd0DH6pZOPdMWAAJARQt0Xv3c0uuTLN/89PRi4em6eCFFo8rYAhs
IslxZpatuFW2k9GFjKXVCV2PVXn2u9u4RyFP4bQozmJzuWDbnLjcG/xfW305UMs1
zkBGte9c69zhwPUsdlAMlzDMCThTJ/5zniy4CkRBqUUbF8KoI3PsCZ8y5do0fNnP
A+CF1G3ov4tWZHLhsKFynT0vvGOtSZ39/9uVQIgF683hk4KQXfmcdrA78EfNcZMD
xuSNKWFNVwv9f6Q1rSNGqVSwoLeGxJqEhIK2doSCqTRVAEk2SJmqEK9IL9Y4CJTy
mzLQEhAQ0MkEG4NeClwIgKvRCq7q4D5B0qZLrnjET5Ak+Rrh0YMKm6bOOhhb/Vfa
wcl97/0KOWGVCbhSM9bepvXpxy16D7qZKNr9cMMM7ffjfljBQRhAAybSLSapjiPg
BlyTRsWZRWRhCLEPoxS3fMXhG9hstYbUnEaEv81uyoDmidPs+TXAfRhW5O8UbsTZ
ZN6TbYp5N2vP5JcniJf+T8r65TRBi1iQWTw7F7cS9lKswm/9FYCIb2dV2HC2mIMm
z3JnjhZrODn1niiVrcLMsV9Us/Eykty/kOBO5lX1z5Zhpd5+0m7n5GeP6HfJqq5v
oLZ0FqRn4P6WQE+SqJuChSYn5UBPf4z9YX42IzdUZC+nkOXpF/HblKisVxHLiyvB
Vh8bN57j/RP8aD+ihlomjOAcbzrCHtir5kzMzn8M7KP4u80tc/1/lV7Tr0k307WA
oHQ0YXke4KFeQBMcDqNdoPHfDAt3rDyFk+Pu0YZ3nbc+/8fydRokbkWvWP8X28GO
HDzMcXoB3EdqG+8gHe81Pw2Orw/thokkPUrR9/sOgRKDCQ179HvOim3XIOErACwQ
fT/dSqd309oHf+4Lg6zxCwrOhXoUx92CINjKZvWljX0FaPpDW6BPZqbkpafOcUMs
dTGXPx2h5HWsi8pz75BxzVBoO1iE4JBp/O1ogxQ3l27k1B2pn+2uAzi9Q3jhWw7+
OdawYEF+xzvy0hPpQWY+GNca+Fyeo18ejdb0KwzxLWkAKC2E8R877PFm7Q3WSH0H
DFoR8SIbllYI9W/8lSzYTEIcudhmfsxtw7g+rmludVhb961BNGCu/yaQou2IbRum
RLiBhfKKmrKqAhmQY1/7jHN22y9bddArHwivxX8yG2G09yuPs8twaug6bV0FjOGb
hzMDXgB+UUTg7k/kDtr78tZs2HIcBQ1tr7KvCz8qu9OrE2reL8ff4vz71mpTPlcx
mAm+UMv5cX3Y66CPYu2p0tGeAsxOrmu2gzDCU5RdXgViXG+TxDYxTLKFaDCQJupY
IPmnBN+rgHCgj7q8eG/fWz8rBUf2q0nm0k89WqW0NSqcap6HTVOY0ryUOUw4QHp1
UyCHYmcApF4XFSewW/z86eoacsXv8Edev7vMn+cE0t35hP8Mk5p4IOdUhHBzUMyg
P+Nlu7ho0j6g9eXPJT3YLPinGBOHlOTqrBLm2CgBPNHseX40Ml1Qvb/gLLG6iQNe
v5U+JJxgoZCu3HYVN3KkAe6OGeZSDLjZUaOyCmg5docXHfxHChOHMQfGGPWnWz9o
ITzpNxh9M+w7T82BEbY27vGGxD8JxQcLye2hiiTzbEY+F+qTvGKk1CWjKAQnKPo6
rg6QvR4PZTqswwMb2FkwN2ZJz0CKB66Ial6t9NPor8K6uHnRt+EvHDbvM0TLt+Kd
XVvDa5TAo1noHqRKN6vT7Lzt/9uLaz0tWJN3O1mQGNuaUsXSV6udyMjVbqAvi3+N
/LKpQnN88QZFd0Ge7mObQMk9pRfA/8ur9sk9Q1CEVfaxCD4IlypyMqr6qIQ29x5o
nP+Djp51Mb4vc9orF7Ti6lkkNpO8Q5NmS/si0uIj/2cdcgPCCVRDlRnq5VRJM06c
KTV/o/lyjja22pRzRIOPFwnZeuiDTIYmR/a98qCi1XXO8e1HC4F1tixRbR/Fn9ra
k1/1hK8myFIHA66mkopFlQV4tsRqqZZuUFAQ9Si/4U8yHs+8dKQXcIEFB1h4QgVJ
WwpMeErnWFFVrt7qfpMRE5MbLWaZscwX2jycxMMTinAkVdV2zfnigYs/1FQtbiHR
E7tUSzO0djErT8eCvq+/28TsD+h9L3gDBD5LA+vaFS/5/L8tNs9VZ1+LwHNEoT4b
BYE11u/B0ul7dSE1egsXGXvkakoHK7KeHNTP4oKXyMN4Dds1Q+ecLDoMXswwWoDm
1FNsmEqXOJ5QAkxZPi6OL1nO7m10VtgCsxXQy2c+ddoCKMbyrSfuF8qh6yctmKoc
SeHuxfORvshcanSbiQj26wr3g+LWfInUjye3jfDtK/LndvVBzPq0BkhJNWLCj01J
SCPE5ksZovIdcIwPXOQrPPEqy10xzyAytdgegCHRaLIZveTQK51LiyVMuqLzoAxA
Uq8DYQdP4ovLgwY3xP85ZVd40fr3yAuwVvzoywO4bO0t8abUlCe7F/8CiwRC+byO
8ZbOvhyKmTdUcGkMhXx8p+1IO/+T398k5mdfao8DWh0RXTAuEsg4DYiiXtHnTmqZ
ohG2mOm9BNq08+rG/GwawONJxofXfMzrAh/l012a22xu3zSMnlxXbGbuledCl/sA
PfsShrQ2j1G3/5jmggiAtToi0UfXlSKy3mKs4rUips9FI9Zy6eLBqYycclCPwo8w
K4au5Gj/ozOKQPHGREGzMm3IbQCDJ5z8K3KLVQc9Ei0WWLzEjYK1sQZ/lN4Y3pgB
ekJn5ZK+fC9Ua3EgKVVhDLchdqG0LeyS1iaCo+MA60GZGOt/W4T9HIfa86u/UdH1
ARlDp84Pq8ix0w87am1r89zDiBQb2NNE0i7mdZyaA9YrnHZuqQSakN0sQdckRR1h
2/j7lbKjYVHlMwcxV7SGY9HL4/5juEsPt0mzEIzX+szC7O5qwK2P8O1rmzAI44Uh
kDHEuk7oTrznODGrnnAwkA83u1c50X7YET6wa9fZYzGTdJJRquEdvBMIU4g18aEa
4I69WMWYm79MSyS8hBixWT0cXzpa9Vd4XD+3bf3MMFJhVPO/64ClN4pP17g08DpF
xassRnqBlGm9fgoKvtkgQOWQBKtZqb3qhPDGX9709JZevR9K/y2LSPMTfdWR7lxU
kvAaZ7SL9Mz8FqlqJt4QB2Uz7nwbEzWD4pRd2Hw4F/YPChvUJ8JW23J21ad1A/Me
fJXOW3DcLfc8QjaEfdxk/Wuz/tcN5Qfv7HuCbHoneWpPeuzl9QJOH6kaII/gTEgL
vqX3Fo7vkrPNJXXFMUEU7EoQCYqKsqBHbwYa1c0SN0NVbo1p2rvjHcKaHw3y/AZB
2mNh+OuZOpA9pG11xPBM3f1rCU2MsR3Idxz8L0uEnmgCSJfAKMkMAnVakEc7oT7i
fWvX5ntcnpPwyn37/SCcDShZDq4oYLb5zhcnS369eTC7oVmdLfp73iTCUJGU+thj
uAVYP9ibp30/6k0gNb9PKjf+m2gkd+0w/kyMhUN0loIMXRxxuYsNtxjUqfeK4W2J
IhMlvircpPY6drXPsxytCnbr3ZLR54gvafM+PyBnmUcVSeQl2bAww6ac3zRDLFHJ
3lDCfXoEDgM35VL+ZsPgmD6C9um9kpBAYOtq0lNjFXSCM/Y92jIeI5iWs0WfNpeT
2fLTurAenMCUHrnJALXIt0+GSJqsF52Y6XIqEp8PNOoV0lemPfm8xAfEb02WKVCj
WQ10DRoULgi4WA8snj/Ks8t/2+E6sMi+omz4vYhpYJcQSiteUWAmMSG/uMfmJiC8
jJ+GpzRuXvPn/lxNVEioBJCBdpJTva54O1vQQsMHrWh0ebEQcCnHphyElZRBC1tW
MKyGwCVwzBAkRmDCKbDXV7yvWply8mk6Ji4Mh3yg9LFEMYRhNaYG5f4RraDzvQsy
EZ61gV5fmhHT9X5QicJms8NZxX5B9VY28ZX6K0BmWK53vD42gmlr/mMo+nnxk5hE
Cn403XemMbfgNEWACi3mO2shYISH978j9d/kxJ1J8s6Swg+UPFgtA0V7Jk0woz4v
2XXNTep/hLLAL8O68EOAtnEr7uGuGPfhrWAI/W32uiuqQz4/mjeSe70XCCI/Jf8Q
TkSBOus+Du0H8zJT1lILNocTh7kwxUrBHToxsT/iyizs+FXGBm3NDenwNREqEF1A
W6dTLdulclr1M9g/9thY6HnL8BNN1U5Vhs+KfkyXdwQk1S5kpLy0g1fleyf1KSgj
5J9gsVvtKg2tq2u2RwSbgAo9X3Lusr3pUB9MW79j4z+Ju3fv5P6ObCCCQGt1vCg0
XqvVrPMUiQGbkRWUdlgVmGXoCtWIi7mF3Wn3lPeqJcL+4z++BI272mVDKRmsMnsY
pr6q0KltqWC5vxNTrEnhyHTxYdxsAnr8J1ADUO7pdVytT5IQvZHaBdj1KJYE6Okx
MTKg17+XJ952PCPQTJPtlhkKHEDBYW06KvVmXBOn3Mug+G2PgKfKY4TZ0X60Dp3I
YOrYfd5g7EqZbMWM8SXI1ozAL2vEdk15jXEX/PmI0grXmfYneAeiCQjyDm4mZEkj
PmYWM9CIHsbHHapoYXs2yGWp2/u3QOpgbHzBXu0yS9uFiTpMrTfpLEFvdtYR5ii/
AoH09eZlskWfqFnxOpU860cPB9mGtp85x4cUqhRi/6HGR86hiMggzgIBLfC9mugf
/TXWT4+SWlHyArM6DUc9AOnnPWTMldH6EOMuqrjqhoYM6qN7mKaR7u77hMQvOEtg
YOa3KSfyYoHywJ2avyA3FlfAybSbQT9ajN+lO7hJathW/BYC22s3k+jRGbPgjsjm
tNckIYF1u7uD1NPM6tcCAKlY7LzcC4ET2Bq91l4a/uAklU9dPXSWv2M12Q7dcOum
Hi1+gOr9grxqlTetXF4hEJFCTRQouRFQup35RTyGS4p+BUn4BuxEoydjd4171jDL
tg2FPIS3oK5VYBS6gPYnVwfAQcqzPq6BkQDbyz8PJpdXlAcYpGCbK5vzP8454BhN
uNun4wX0N+GmIuh/B3zssuysdpvaQcnDCYWBxN/MAFMe0mGZvQCgBIBcDrOrjiEU
tDh5a/vB0vg2+7/m2nTpbbbtsYKWxSBonMZTc7e+t/HblngKovYHpar4NAJFnMjh
1fga9PR2H/IrwZUfBQi5w0kJudBy7mAzn/DytgzIcOPws4f8sv06ohwIsabdSCs8
N9/67Fy2XLUKb399+R/pjsaJ0+s62+km5keIlFiQPO5UPupjMWPeYh6FSO4wkEhf
zO6RcK4UZNFJDwll6+uHyvZSx7Su2E8LbE+EFDTFwB4KoMaYWkcYRxaL3VbMi7wN
v25zCId4DmKjtL5Le1o/DeJmsIHgs/5FoOVcQzv3WC2wBo3PM7shDUboODg6lWHZ
zfjGZvyVEuaT8+esPntXciUlGudTnk1Ri/Tj4hvViGphw1oW40cPn79sJM3LVt6h
SCQpTJhdPMpZpcF2KdoaSNQLmn6tgm0ZkyZBCM5XXWgz1zft0xTWhTOBLdNktvIQ
GEbA7jglvbhf7pO5pOKSpdMAQDSkKNhn7GXg5Qh5HhGIMDh8NBA4zknOVz2fR2oO
bt77yR9yqyG/XlFVt/D5zyIFtmGUhTPBt6/t6IrM776Qfn2c/gmrB0+GU+CaRAy7
1bkainA2XhdAilcDx0Svbe8SKjeqKMUbUgP2xM/89mWELVTDUpm/trDFyn5jb0VN
fMoPaov6qQLFymcH7Cc/6pq8OZUpHojAffe7QrY9hMGtjKft7jDrMCb0YvGBl8BC
EO67Pxo1/lj03GlNyjrHgxtmZs7lZyz9p83QZfEBqPoOKOmjkN4j+IQLoTBiQ74R
rhkQWiASE29jMxi3922DZqdv0sM3FFuSyGJSuWZXByB8Djzer0qyJMgfVVXGMgFc
wSPTtfNFmOxfEZ7H5bjQKb+KigQEjmtVy+5jiC/+K/um8P4Z12P1K+qgzbHpeSw8
iHJo5XAmDrLhz66Hkgdd2J+jisUQuncZ4PTChVNxpBpnlubE6oAUH420FtpiNOBJ
rGfDtc9IRgL3sFa1Xv/mc5u0FkBzHKuYUirqtbwu1krp6fFOpdJ+sSD75HPkKYAl
72AA+vLrsO1zKPcCG4j2AOguBa7kM5EyMz+hzlmxy9f8RT4fboNvLfu2/oB2hJFK
ZvEv53NHFCom8lv9nEIct8BwTz+jsVS+JdU9dI4+GrUlgKjfZe9k0R+8iMcUG3CM
80dnI0WiZbya4UCVZbhdmBr29Lt+uKSIoFuqpNSUNMG+S8xWWno/burYbZLfD+Xt
eAFHPLPR0BcUSTM3l0WcSIXgR9pDc6T8nIlRHx5W6MBvPeEVRk+O8vexkCB5yEI5
sPbUD958BPJ4piKvYI/k8KmMLH5jomZI5+T1SHQH2k0sX0ktaoJVrZlbDhdrNPwk
yNIr7lZ9q9sH93OZc3ASWFHS/qFHeLueHrlhplhcscHaRCZUP3FmVvsZ9gmyJZND
dXMRpe57N+u2MIfhWhJcEItSjdP0sDGejK2bswM14yMFE9nArAqp85oiWWRXD19H
Zi5sAkCxlSqqzrwh8sRec+LuLxiZ9CeNLZR76XKMubJvWeGp0+0yx3DWFluNJxPL
KEM8Vq5kmdD1v+T2C1jpWIDOfAtIlLtXSA2ZZNgRign23Xjl0Onpx+KR1+baqSVZ
fdiV/I0/TzOBKF9G2WthnBZxCv1cSukg2DLImmukQwJ+HG8XrmELqca9Q1Sx/lsr
g27nW9ZY7+IQ0/PaLqW5iPFmifhXb67V4XvRk662T+X+PBtpoDcqM1KoJHNBJJ3a
Gz1eMQwYgXldlarCaK+JT6l4eNRDZQMEGc0wsMcssqejLmfDydoOD5kOs7hgJOPk
Wdgyu5k4au6hcT2wZ1dNIke3rdeAJ9WkQWtKlkwkfjhHIq+d0qzYmOofOMktP7sF
9wzMCPvQCN+ryexg94E8q5eZUWLsG0eV4Y1buZQCT/UwLDBqqgpikq3q0r916OVN
ubaCT1rAcl+soIvD7+bpzy0Mif/RQocRAokmFHDCjj1XdJpAf4Lq2h8S8neRpQJX
QixCAJD4RMY/cZU5fCb968K0rNhJ9sMqKD5D6yFkqZYH0cXf+L+ByfFf5GD8iiUf
5IC0QKkWJmLp1S3UuhjD10ITVVej8lb1g7OGc7TzspZl53xqdHPfC/PxCJ8abPzg
fJpWKJ+ywOHLqmsnH/1zD85mlQ2w5oziSssjhzBSa49xlrN206hFNOPhlwh80+/f
oybUAqoGdPkQYhQ9LsSiuIvr/qyAuCrIvOgOG5RzSDNLEnv8/VYc5U0BbwDM4P+Z
FTZPo/BmCfdzb9Pn0PaDgZUo5bx0fPxO/NZ0n+NQqQs7OciP2J5y8CHBKI5YWqdq
kmAwzyg/A43e0RCO4hlZfkq/2vaFCDWNMR3jVk2RdBThbd7gtcUSu+oHhf1BSO/z
na18XYHenG0RfZ01uJo1aE03t6OLxVWiQjqI9gqJVZRZbdDJKcXSykqzntMI0wZe
k+18CQsdnGhT7YFJ+mQBd/Iok5DvHFQijvxM3YQfj44lBFLY/5MC4g9Ybh+3Zlds
r7Bxg/Oap8Vq0Cdot7MiuX0e7RY1vdozgGR3iyazMvRjGx87qNbkJNVq/7DKlIql
J3CI9mV1RlAtBdHIusUZgpxdWWGlp4q9Fd1M6ZLuZap9Tv9LDwJzu3D0hss8IxjZ
UrH5E4i4Mzrlqh9LVZpQoK0WW4fegmX4a7YVZMDsL+BUvGoYMN5QZmq513zMZlIA
cvn/ySlhXDlWxy3dVxYTyIJwNWR2VehjUvoyf7BNxoeL6Yf4BljrjQxRnQ3A6Fn8
Mf9YSxyudLUCVmj03hfyKd/RJjdj3ZLDbe4OBKggLAe5bgdofJ3bN+Zb4D0lAGDC
mksl7nYr0fXGCBDgVMGQSONuGURBE3JQtRxAQGTDOgxc+4lEba5eq8pCaDre+f8g
uFwwtM+yfPOorfltRu1VNkg75aWbwYNhkXFE+NESBZiqSdpKEem0Xjua4f1G9TKn
Jq8F824Cmm46m8vJpRGLGT0SK7dd8fI9ZBq3WKy4fD7GcJYnwvBet8F5f7Ti2VIn
x08j9Yby2/UIJH+MqG9/XulZbqZBcWUcR4NBB80fj64FPKtfyJfq0nrAASax7EQ1
r1n2v2JQC5VG2TfgMoSNrcq74hC8DgReDdeXFsZcOFi5l7DBq5em37o8DYWkARHT
QGls8u3tRpY4LLhPE201ImVcVnIhpAjCkq69X5RBTufosk3vgk48dNhVZMSS/pRp
a1uqagNeE/rF1d4FsCa1fhRqwiw13IxiDJLBnCFGlpPpjdKwERqR3ng/PwRkT8VS
bO+WlfuFEDM0bSyn/atdLB/W0sF9PId5+yby0hdl+KxNxegKswVe/RTZpdclnK44
OI5Z91OQeTPiLOUjSN4goPEvRZn15JrZEjTy24zelUDTa9HTpxf2x2JjZzVepS7O
oW4qCRvL/PE6K9bZicNci1Z/FsaspT4FQrlUIpac2g+D4ybxEDSUeDl6Xj1seB/Q
mndJ1UyO4ri6hKsEGBVYz5L4A4p1FFaQUkQ3O337iNRcQmJ3S1TCFJuOVmY5DLRk
Krbl2Fq/6WmyxfNK8jbHbq1tomoMbNWyfO58UAsfC60opajZh9H5QmAvYPXzLhJ7
M/R0VRdMiK7gpYutpU0sjhhRCdFIAoPPJpz9zCO7UluzBveTbvl0WQAfwfyJu8h2
6IipjGU01PkdZ0zRMhcJNMv979NFNHXjbEebz/2dHB8Zjj0/eZETe13YrwCSlDxf
mOQpph9XgxxOaGAZsEP53fuj77AQ9q2husxFBUd30dho4xK+me64ZbaBEXg+6sTO
+TgIFcmENH784h3QTS2Oh9x+uc2KkpnwnTOg0WeFOEZZ/ieonN/3jtFf/aEybxCk
meZaHW7ll74BYdi5+XU389M5FDUqeNvXswxzBnr89CJcTCm/T0TZieOMKyTdWRLI
Wzh//qrjhhySDnIVi6SBRo3YJw2KLuNztraSH8FQIHq30cMPRtXzZLFCVyNGedF5
dXCXJxIP4wN/6PJjl6elosqT4PtQKW1+iLUOM2vzvZQNNQnNbh2vw5bpJdSmTOuT
qPUmKKpnd/8aLIGOY1FFiQRRz4PdaRoZekWQV3NL3uLLGHH8gj7FvRNyEoW58csR
3lwAKZMvXG5UO2X5nX5FARiaqJtrvj+Pw5NHJtnkKFvl3YhhQlHMSwPF+9pUnZ61
m63hxPo9J/tNTUvS2n9s1IcneptbvueEFj5i7X2VLLKkDkRKcRuTbQFfSMqTL8s6
ar5Zbbds5bYrxIrCciZIVD+vsv3+21FsKkML0Ct+T+XkH5ZVyebq33oE48jS8OZ8
kHRvSG7wT0QC5k+KuCzHJJaikHyHCnRmOwmYmvY6y2ikvEYYVpNDsNAt63b1k7QA
0DNiEFxOXA97MvaTDbEK+mVD1igqf6dCHJrsFu73ngBeTRTe6sP8YywDxJ8XXMoc
hFDXvz2qDQ/HYbLml057rZ01OmdcUqfYO0fTga2DO0Cwgl4s5KVtRdAW6dTkTRRr
Iwcb6fLE0DW7sgqui0t+8oj+kmJFzyL3Cf6s/Sh6hTXNie8tQvg9GRogK59GU5sd
qvNPORTTgrkr3oSGCgdMDer2BbZn1Ip6Egz2SOUQHpf7ugjpC+qYjgT70rDc5GsG
TJFKZFPbTZcsT4uim+qb1uZuLc/6Xwjz32DhyHEiOx/GQHf9jcnO1iGEwYbQS1af
APOSU6gb2csNbGP3yFrm9JnksHOXKv9URuK6PBqFSZ66rfsLjjvCvLsvs6hh205q
sSei4fpvcuu5futkK8+GBpIntzhkmYgcxl0CL20OQF/mJJUBx6BTAJFgBeRNB98c
Fr1VYFK3eGeQf+M39+uQOLzHYjgsB/4fy9YbGkfuSBlVRFo+C2MSt+zZixMqBhtz
tkZR8IyaIzpqEkX1p8G/txWQMnjZR7zb3BWBbK3tPzYgrs6p8f2EW3Fmd4tRzUxO
GAmMy31pN2KiL5zzo5q36ececlVzB2o6FYVO4NMBc8kr5JD2lEayDOVWJZ1ltJOK
cePpECYRNesMsuIRfsiV/GTYtm69sbIeYVh80J06lsKE7V38tgKVf+h+R3lVNHZ3
GZRbPh6R+zlI8QMydnNYdyg4iuuksrVJCiLfsEi9Td7TPNLOik6MMsb6AeQTV0b0
QiMm1b1qxsG35MxQuxLS+KSBJahTzD/qjYPaG3tN929bsxZ0XcIdZaKIVAoTqILK
Jze8/0vLdQ6PY7a7rKaYbQXRSaBrPO9m4M0zOo4VoFTNbvmPq4CcrbIRUSPKu/mi
7xUG80i8XU0heaubhLcM90nmvTuf/U6X3+6gBhhbLVLZj90v/hPePqTX7sDDNPyK
PPXroMVKnRDNPJq2+AbYoBIkisBzwh55XERdilQSGB+6CmbI6BH9U+vCW22q/Tpp
JxAUbGdP6Ix/PRXTNKMs2bVcY5kS1tu5j89oIo4OXdHAOwBaKbzS34dNY3E//uUP
sZIsrLxZWDTh1z4g+4c+wBHZUMUy3FpY732xwyVKHJRtOEidPUnMAS/31ngOdyIz
PNOQBpUcYxGXrShK8l2cKlPdEmOc2r//Cg7SBHFh/ymlBIg/Wh79YMuz+xu7Y4ma
0Zo2AI77C5dccrmsUZpilyQCZI7CZvqMtXZjnsoNd5pqtT9XgDtZVAXCe7qBiMGo
6EJ7tqe44ZEzsTwDQlCtDJEcZ/mBVaZkO6acSoZxVQ/4ICRCKhbYUTrTfhzSVJI0
uAMU8tKLsr2o5HQuM1OMrDZ6b/cu5f4Wy3G1M/oWq5Uc12t9LyUXRxduQKEd/m7K
gJJsukulC88HvQL3XKGUC3rh8quA6q+R3a1hFdznfr7egbVmFPnuDcz2J5ydqfrH
hjteYKtgEj5oJKJr6mAGc/fGDu2NFeEKMkIKQ7fuY3KrAYwU2elSFHFmZ0iw7vwv
YwKq9TuyFZANs31wkR5tokDnaZJfQKQiOiL/ybSLLz+MSbHQ8R2sQh8dRoCE/JKB
+vRpfXg1gsC4ft/gi0hRJ1/YJvStpY7J6vGFrjpVNTrIwO7fpq4XRk0Q5w/4pbQo
EBLPMnvc1xiY1KmDZPZe9ohb3TGcjIfoHk8L319dXOzT+jgMiVL5xZwhaapaqDMs
cn+LvzCiGMFcbEZqYr0ExfJz5zHNQUwkWKFTQqnPXkZP2OO9UQhurkI5eM0f9+SW
pH+/RnFGiuNCjIhaRV2MMvTX7ypSuSwA3UynkUKyY73LRxa5VsOO7V1ljDmPwi9l
TGJwOUUe0xHWtSC7PgvTbgildSLZStNTOPRJJAAIw0T2S2AZehOLJv4uHWueWWMx
LOfQ2nW0aClmxjuE2awFZnYWSlGRRDjCkj3m2tRZGiCdVD96IQY7it3mGTsPk3Hp
JeTk7lzZuhsthp/9Fw+AB4ZEO99y0hQEtZZ6GvtLE4ZLUJEi2daCBDl7Ihb/ZBFx
6AXeb/o5CuC5Q2oiYZekGDCUTevs895zeHhZ9s2Z1mejE2vdRraYLBlrV04j3kNH
8ik9rGmdzlSWuZllzAP/F1I7tqFwdQg5/Nq8nndmVaFKc2dTNMxzw1ipnz679RpB
MvV+9th3uRLtGI9wtTG3eITU071JkGvAlYFvVDY/7VwoeM0qKRLqzEwrquLpqkqM
P2u94VZT3ihs19zd1XkoA7h2xhJlVGJZUUarMYsfMZqsdRYSvb+HnSYkHSSeE8Bz
m+pC/yfeblcgC3vdUb6XVmMi/rCFir3YWqN0EhpCLagPdysmeVQGvOXlU/F5xYqv
W89GBSQ0WHqRvEVwnzfvf/NQXoXIsUo9gUq6Y3CxwO1M/YAEls7yxN2R3AfcpAH1
s5AkBswvqZqvPueArkiFscoKhuUTkgqTTXAIwI3x5g2gV8QBQpozMv+DT/M6wimc
lTo6fbRazjCOzFG3n1ud/qUTzYmfYyaxQ5ZcSDrClgbEqdXJjkLJ9cTQ5Ij4CK0x
9XGtVjyzpjDXwOJ4QJ0EYiLoELWMw9e1+OYf+KFNYa9IzNF/L6phjyjdtkf+F1Zy
GkcUViiWopKaYR0Im1Dxp9KtLTg5VE/FlMzuQ273KfmDqXdUBWOXRiWFuab1bTYU
K8HltaZIzlLY2w3z7zCA/fup2hXJHAphmPNFuE/jsO4/nMYRWWrTMDtFuvvgigmO
u56C/N3WNUH0vkJG+607JNe/XYEYORBraTl0erypqUvbvg8GoDgcUjZIf6NPyKny
FFDqiRpdNAQS2gvtEfM82peZ/8o25coFdlDnBCZWMDRaSmXTGny8BCT8y8XF30Fx
mZey33la3sezs+eIVcsN8ipPojF9OhsuGejULevYA0FxLavkjd4CASuH0tqaDhH1
1JDU7QrQvRIK1X6p4k2goU0kF7sARexSZrOJuxWKuSVyfmU+4OMT8jTJmBDkzbcU
sEm8KDV9FvxZlMA2ZPC/8eXd1WTilRnqEDyY//olBtlCM2fAkU/D74XZfKJPD/Af
L148YEQk5ZaqJgykTE/+rdvNrnGZGyR7wgI3JudLymz5JWneTSuGqPd1FpNy3XsR
bJ1w8O/MWCcclmjYv+Mfi/kRFfvqfwHRPsaQaN7kyUsPGPYt2h7L6gsYoh9p6Ptd
sIISjq3mgUTGAb0g0EXaHgbFZ/dl1WU3wx62U+wDahY/w6IaLWlv0vwEPYBl4pgX
UDj94zA/P0kmIzMAl5ARCDMjJkdVztaK50qvbLZerxy0iUBLVKTCpFKKNsi2QY7+
FcAJUQs08JLCBKylsTxRGM2UBlFVfI+CN3WCXUCdrteqA54Bs8kZurxtAO0lmVt7
mDrlxhoZowYTsNwgcxZGtCM5JO9pp523kMN2NJ4TJZ9HssmBGXGHa30mK601ocdf
XW08xVDBvQVJLmDq3YJcrdZR0cDdga2pTaimVddzDNQRRqQzu40LXRmaTUBztc20
+w5Uhr1+c91bpHGyCFUKKpKaVpU093bN5Xx7ZPqxCzOfLQTVIWFMY7iffQ3KEzw8
5Ewlasd7S26MzIdUs4mfW4/lLk4Auknq1PRJxal651prnPUtBfP1Qu5QWkGUfq5D
wAejZZOh5Ed5hUgaHcBWJIbmGOefzVbxUP6Kq5FJFItoNpEDRFzFE8366lpCkfrO
oxXFsm/jlsYF5DkUAvN0imc0Oeww99h4VMnYtF17d6Qk5gmzhY/sOYCppUUIwwOI
wBgjTrF9iQWBU3xgd7MaepFneErs1zW7rnGTVd4GMjVxRArQR/Us00p3OIsf7Y+i
sUrz7SPwxeUBaLVdT1Ih9f57+aada8XfCN9SHcbba1zsTJbEZVj5i5mP6J0IPkON
qI0k6+zwGEUdEiyLcaMAx1ZD9/WKf1QAcDsl1vulbjj1IAbrPRoAOY3eLacnovI5
FZfZKblnt1DSvCRE5GyAUibd39lyKI34x4M5bsq5MysdtXsZaJSPz7VGD5fqlEdG
a5SlH2aK8wQaKt6isEyQr1XAcA5eU66quKXqEpAfy5KRmnUOWJsGEi372mV9nsds
DcRDC4tPDXAyOFoHoOmimEfVqTDozxvPDTxHD6jFZe7DAQ59RXciXVHGPtuO3K9m
GLv6e7d+XtgMMLSr+T0AXQ7X8KvnS+dXgTLkRA65ZSdFSE7lOfIFxiwx2ckuxk42
pXHQUXp7vb58n92vp3sgZT4wQzL+GCNeFhDl6zJVvhtC/91/ONGrVPZOPSwYD4g8
n78fZNsXgOFq9yqPPXYSJ0JOb3a93cW5nqkv3xEh3vD0ohxQvsYRAJXCqhRkWm6m
ZVRG78d6hShUS1ne+blbXs3DZ4BD2vstvAFzkXemjbJ+u8CURuTX28NcF363ZWDK
mTUsod46qlBfStkOGxAr94pjy/QCAMMubJblcU+UMbQgm1H2/UxEN8gJ06sM8FwG
J4LYp8f28xVX/TeAC0DNGiYZe5ABJcLmusxZEvXXRBxfF3h6KeJvkWtlsCJD41Eu
u7tHthCpJZWsCxOLMCxATObpw3iJHrxBAtWjizK5jZAHhC9aIsABrQoDJbwd+JQ1
Lo4uMzlyZi2DE6hYxzjHcNXPvC4rAu+vPjuZcbdyAYkgpXZ9zOUtK4dkJd5jS8mw
5KqdaKtBQ47chCzTVzsHB3Y74Quwcwug1/nVpRGw6CWHjiLqJp/W0e2pHlaBshTV
eUDSRenkggbVknpa0DY4GEYjS8nS59iKc6xxVltdqnJFFEpurda9dVuQ6xUsbicj
lc1qI9acViXRllLqbww6tjGpifz8vng/pbmx+GnSSQu/Hp54VkolLstglU3W1/6U
J8hEz9Uq79VeQ6qkvjAbacGr+Y5TBoc0oyd5TH8M/3ZYBmgYh9vJlc7wWTEgZi4O
zhqaRCqXoXKjISqEDtsAPJycceFfA8UIIIMa82Hv8loTglfCvuVWvt5nZ7otLqF7
7vqvV69xneLwoXICJ54DNfhjk9WC7qZnqeWKyAER68EU9qRJBZMLMJgFaTaKboCP
VDLfvTQjAk+9CZ9BVeY2mU43tapsUVAy+o5wXn/jZ/zzWupEPXIC4yCSuC1jtTt8
lWsaWeljqeyyjU+8+GJzUe2K1J8nd/T7ZJ64BCkph7cny6W4z73/BtSyAzLJnTHH
DTrBbFMGPdjHVJNTZylkrFb6NSh52F1+xXnn37LSEqTP0/IgmP8nTYiYcVr4o6yc
wGOqzXXZFzEkLeSkvhEi+8WSOl/TPiGSSTpsJHkbf77+wh+Rv52DCMRND9+G26b4
O/WyaIsfNhq/Yb3qpyEDdyi7vToOeC9yUtQYvYa4AqyD0XrIR+SjvUKefH3ruTO8
SSHWaKx9yEJuoGyuRngkBohor8GJETL9GQJpLVE7V3qL9HbOgZs3FV2FOlin92IU
RzwMWxZTTUC8WxOQLS369lVn4NRxa9hHkGCJlPuC6bfit/+NaXGYEigL6Ha8A/9x
nZehTNZ9dmUykoPZQBgQN6HRpQvmjHtKJqC5DvwpaheQVpXy4BVZ1LzVNPsBqiMv
epzhrwW+j+onZgez8kWktAbtLFiR/RsuXt0fUvVLU8nzqnReE1Zcq/DzfWBxGnHZ
1z4l/Tn1G/z8/tVydeqc7Zd719FPZpRX0wUMNNC3KOXwbe1BD529GNqooac/hUpZ
MzXSOg/EC65WF+ZLDmdNgiO6i9ZLOHq0KAgHbdtioAdh9pXiKfkgA6+/E7JMbLep
ipCKf5VC6fwlsPbDr498t4nQaVgbLLym2qFgoEWjJQdAMNWrwZ/+A8DZEP7m66Ha
vYw9M8X4XyAnMF0gjttAkhq3MYa2WePbt+8J1Sy3x/3Ez4dKIgkGuU1SWH5tHp28
rmKd44k283WgvyKjMM7t2avSLVxnSEbXZZi5CmHWZ8AAdMTEVLb2+HYF773ymh6m
ZTjtEI0i2XT9DvcwJhtMAekxiBwOe+k3I7Nv+eofEoKzpuZXRZM6fK3x5zRNOdhC
ZmpvbyvzTDe3cGO+ZdGoxte5/iiEMKv3t6rvbYKCW0nUoujrUlqEavFWIj8VLXEr
j7QlvlYPz0lZh9D8bOWVoRequqn4ufOPL7hlGKKz7MTIGVPSymw9H7QtBkfaYD52
Bk2GB8U7OHdQry/5kEK5ItOkCEGxeY9+JvvgbjADUZDIhBj4KvGA5Me3S7E+646h
+ksVRMqYpHvcrMpGuC89my7hBzdi8h29Aeo+xWBbstZ90e+U/c2A8kMC+llQUzj3
PYNyhUVmih5y4/HXCtovpZIEA5/pAzck0pe7j59tFAcEKQ2dyVqzm0bZEozYIXIW
kTdxv8JJgRCbl2XvhuexzYZPzurKbVH3ToclXDJHJrXcPByF1Y5+hi+y65eVbIeL
8Sf724jYEoaPcy9d7Or4Ywbnh3iaJsfCm6Fs4LFMYzKW30EwlCBU6hmOE9BTBlkr
08CLBn90TR+U0QdMfvJIbmrxqQH0X/za0W1g5YU+EBORcZXCrUm2nfxUFYyPKpv2
m80P+GfO5Ib1Ec7ecSEee/FM4sFsSTUvVGX2dFXoOhvklafnBrcNScKPI92XfivK
6yUZ8zELNO8eiO4vFY0yMFRqCTwQi8xxcbKxRSrf0UvgOZidH3pHQjrbYqa0NSe6
OGat5Gd7KotRTCRVJN/m/mTNOySpE/2FeqF+izG4kevHuD6hMHBEa+LjSYafwD8D
aaXvJk2v3FZs4c6bPwPlI+y8GtB2jfWeuCaCeb1dDHzcWZ2piId8p6ZG2ywD6jhi
puWoQkyPyH8rnQmoJib9uvDVMFD+NTYa9PyZmKi5T7ppuDAZKaP98cxEcn5fCx6I
EWeUeb1H3v7KM5DFoj/tnzhdh/Ps/FkWHs1Is8bMGA+J15zezMSCsk+cjyAVBnQY
NW8BgEAgkFuDxdMYNQ2NF3eLUFZBi565biwVt0GJ5FBKTbxCfE8bSbHBCqega9ZK
XKtdp9wpNzXaPpNhE6ynyUYYeZGVhd4zEPF2ukGnUtPzcP5asmf+Re8HYz1/BlmP
8imUBuaUDfNSezpMxTbZkS+Bcjy5KYAKX5NtdRQTi7uboFDdLhx4mfjm5hUNrlfx
tj0ZSj9bSOu39aP74JUtV3ODkuC0ugWWoFW5lT9nmEqQgYd6TAkaU9zw9ru/VpZf
VhjzGxsmxfyKIegCTWlUDr5vlsCRwduS0FxKfY2S8IwL7/PzeZYHDLQukFoYjMux
1st8U+NPZLB77a8fvJcD8werxAArt19JlnQHld+dwJwg62SevnP+ib5VIwKe1UkK
2b4BwvPBRgOY4Ixo0AUfG6b2XoXs66mSYPw5XSi5vd7+Tvg8CpCUoycdAIw/REKj
2+I+Fm3ZTdgw1sllsJrNGpOeLPbG0oDCcTxOdBbUslf9qNciK239dRwD5uvJs048
XDENP4QjthhKitARPc+P965oo/jhij444uuFQqdkARG0K1YH3Kj4cAQ9IV4yZMPp
3IFjI3ZsaboRwJMQWdMKkv/LJTe3makHN+NCl52fnSbpUPGIXG1VhzIcQPwiXogI
uWpvIz9Ox++Ig6F2nOzHdkIHNnRJdmf33eViT8AsTwX5ZxBzEyj31Xd94UMjr1lx
AsFDZoeAZII/cwC+YzUyWPdIeITguoE3S95W9Yk9PhylLYA+nLvz2yb3cNwABY+X
Dkbuea8eAFarqxyFPFD/UIz7MSRN94mfrwHCKdXXRojFNuZR0EESo/CB6FrO6MsT
pmuIHVqh7Y7qqVKffrZNWv9npMfS8iy79wBKqDMFaV4g8xelAiQ+yZzvZXa1OK6z
NIMxFKqSV9JDCdTfTpcrOVsc1QLfYhkkkirFUMIvl2UjXcoN9DdQ74FGvQfkyeEx
8yL9BnmmbZySDEQSxHedh38ToDvTb25HT9G6zsz08PEGnfW743iEtnsrHZEmwfb8
ABRpXk3YX262vNHb21Ir7qq+ungDdwTs2t+2NZ7GwkM6IEeteie4oYpQq7D9MpWJ
V0ZBpccMy9578vywzEBoKc7YWTPXW9Id0OCoPZIFu7XP5tUvD+yX4Tb2MjMQy+fL
gnx+KXQfJjSxng+zPRM5inA1JgSftV9Q6KigDmMnufvH9bB7NrVulRqFZtHBRZIX
2sDbaaKz2DqqGKeGcVUAQ1tw5TGB1k4g2I1mFBzZQZItZMQcXFV160gHNCTwVDYL
75C0Pt2PD/0AmuPoaITEZQfV9mo20suqZbxZpLz9KQ7PEY79b4uqLRGRQ7DanvLr
mcxQnDvJ9wEEc3rx8mic948FKkdDg4XklJosLeGMfQCbKugFxI5DKdtZYwcqY3Bn
rU9VooAwNzK8HVOlYaevOxs7thRFdJu827X7TsUZqWunGOLs8wYXA3XYUEJVRJIq
T6kPFlScsXTFVYO9AsAe/VAfY9I/hoGQg+GMj2qBdt/2TKEODze+cW9EMOdCitpe
R7DzGq5DKVPyGaB1hRDmnFv/Iw3oFM5qtLWtpq8/yPPfCc473ap/fNPX51YiiWsO
gagRoI95woMWmnSr46o4q6nGKpgYuHYGPOSkYGsBmR+M+wGdmD1OyH6pbk7/bJv2
Zjeeo4tNFFsYPymB9ZVI+zweIWC5765OAxwU/kMDTPCzRn+GSiI5sioMxbHxMhqq
FEmM+FAXc83QrNYM23yP8DKOj8wXhRA+LinwYWnKJ2EQnTajTqxE54tRHpooORJV
L9PLNIDStUWNEE0QIeaWNDALfyjPr/iSVkFssp3498QNeQTldbrSKsFcgLHTJrfh
1cHEP5GbWJsN+LsAQFJJW8ttcus00P2HPrhJp/EdX4jpkFBLVxEI5solvZ/u0sE4
0wm0QWBO+X4hxDluFUJ7mOk1qtxQyeFw/kLMuvunWrnNroEaa6qI0yEGjCN4t7TZ
Clpy2e73AXBcsuow0u4DdagtNeHRvbALZw9MGB4BfSJzz6fsd2HYzBVLb/kYYbrY
dK+tawnPThqzYQ3oXR7FnFzUGHmZPX8n6ttgrd0M4uiznuPDTEvFSwdB8E/JgSwn
8Toq8hQrQynJ2p8hCuVhIZTGzDGUPKNhHeKCHl+nQF2TOxAIy9ZKQOX6tvtuKsH7
tGCynpRMOnMP486QhruB0CEYsh90VO+ggwZR3R/bsDyejMa1uyfQvSvNja5rFNWx
lAxCpeY479hJLQZ/ghlblQO4dgLFSHJvQ4YEvtdWxeWSInniLIieyVuB9VZB+Hxd
Ksjq0P+juLxQHJ2Ay+wOXJnVan7Dn7uPTQOWdx55zQJwun5VVLEFXQwRL7gJEET+
jQscvUGBhXyDpWZLJ7Fhjmp+DA355whzrxTtBjWn13Ofl4yqdS07n2mYOhojeXWu
OLqrZW8R2PHNCReXP7GnVlqlUyg56fdn8tPYprEiAHqBGmQGNU1ZDN5Yjq2cvkBc
N/pKm2vvdnDmZjF1hhOSnoRY5matfThnaapjmjmqp4ktLZpSEFCwwmFD/xB0SJa3
SmSdBmk/WWdhcoo3mwsbXoRvnuOz9DzDhaQETNBD4f1d3E/k+7Z3wwfluyhjS6AH
z/qmJbxHLJ90D309Bs+WHCDafiW/wzpxPq6AnBN4ZsjJtbd6ulK/jQJsQMJ+So/o
cDsRnSAnnt3UXbrUf7rvS8YYDpRgjb2udmNVk3nMykomUuurnDGk9eVlKoPf4469
H0dMT8LUoNybJJPE11fC+nY+pPfwIymckhtH2+EJf3sbcgwqMwo+gS2CNPei+AVh
hTcHs0ipDKj7m4cNWNqxe2Bw47d5ODV5jJ+ggGgohmMBj4tzBnPB0xOMcw20Yk+t
TuvE0ydGUy2bhBKgZmcjd+VrCdXJJBbM7eKv7SgemaRo2rj2T0/CPJGM63mnPY5k
H2AEfGlSEIhyvHmy6TtUZN2IcwyeRige9qAeSiGbIPCU2/eoFrflIHXPsLszJ0zf
+7JW6aCDEusoEtIYpPI8K5bdpsMG1YOBm3dZsQaUIO1Hzvdfbl2X4K/WcLPzx9zR
aA0LsjG+eTRD5wKWvGpsayXeAYRY4xjCLSC6Kpt70TiLJGMFCAbvgxTOeR3oXnSU
SbyEemtfUFMHZKxzhynZbze42hKuOYOghIFMS1jvkBHADR2nQabiyKQf/ahpkhAV
yZVs8jl8cVZ/y9zKhGASWAtr64ZqZfznjM3FrCyfFB/+ZmOvWX/XvIyxmk//OflP
ckrqTMOdus6eXmUcJU09jLs/HA8GojQv1KCsayOZskwzCsWLG2k8sNWRolLHAu0o
2IwVbr7EYI3GxZvvc7VosvtDDLUG6rC+m+kR3ms2Yzml6DY70b7mVvYwcb5Q8WVY
r7t7nWWULlVUatxfrEzp1FVjSnE2OwWzYMYs4x3+sXPYx2PflBSwHXi+oRzABpUG
/6lr8n+JYQ98ZknNq0WMCmil9EymMwcyCoS9AifKo4Ev1FSpAGMawxbbIQcFQ0eN
Xb0csjdcedxDCSjv9SUb05PZDcyluVO4G9+bE5z9kxzEbmN15Tnw30IC/kzHmAMq
mA81ltpbdMxfzhXoeA3JBlh7Xe4R7W/bxY1k2N6pFXoHJ/v1/gOfyatjnvXyu9yn
0vMIXhmSXZ5tYvUwPUkKezY+eqqnTLYGHTubFAbEKZySrg1g5UTj65jkImzwc+w9
0riH3nRuIBjhc6Vfmg0uAu9Hmw1enbfApQSr0+3iLPeasppbs0P6wAMJbvnVOAMD
J/O5vWw7urfs1pvMqdbXhI4NnWr7WtZmZMEdFmOVgABr3JH2O5cOqg1a1W01zfL+
Dp4iiBPcRFXTY6JjYdwyHSuERSirVfSnhicCumNP88TG1ozaexrhQJ0q3HLD5cec
uc95nkkr2C1PBR+Z3XNUOqizGgPUtWLhVFIAfPmRc7sNyLE2sPvqazdK0OjVLroL
s4ftSZzC2hMWie+GMBY20j30K8iYlUji8PeS494zIDVneZhAKxCZr/eGkCMsto7C
UHzp+gNMztirAtfespiZhKSBILrzvsO9a8FLHvsshocbQdl5l/LsxUizUaiam7Nz
dD6aoxKZ6J4JIBC83N28XYj1S9XNMfRvTPYEKSNnTEP1OjHZN7z0oskKcEwfZ8Z0
P043Z44WNStzjFpcl4QghPDqkGBrvkxAVCvSjAAm1BRlPhHGDILwfyDOr/Q0CJHU
yVGQ5fJJ0YXAg/nRrEGY5Y3YSJ20fug1AeGp4S36WQsUP54IfWwWdUzvjYndj22D
RGY5cTUdejWdhUmvHdipMdQuY+AU4HQmfzULo3YH/KlZVYGT9M79UH4EM1nCZSwV
yB7WwghNZEpYxmreQCsYT5w/r86lVxFCBwUgfz3ZdvWyu/bem7TvG4Gt5R9MvIOO
S8nR1q/sRhB0PWv5ioZiwcfaMn/KfQ0+okKgDGXDRbhfO/6knujkbW7sQ9IL1Mdv
/uKQmzjJERTk7EAommog3hznRF0C3cujMcFLAOOFWmZYzRwpLEZcJkOXWBHclzDL
sIuKkSz8C07MEdfScVwphfXznokDveiwsRmvR1MrzDHQb4NT2MoD0zAZW73aja7J
q36pOv5JzauWtQY0T2CRy0Qbl+r4Ms4+U3r6rpGy+ZrnwzqbUT98yTOvY2BHS4wS
+7HrACp1ljuyXgAHY3/eqSN5tdDJKkOMIxBERQT8LSs9S9yUN63IqAei2kbnp4Jj
I8vzeZIMtfeXGVdJ/+HcktvuOmhU50TkTVuKnWuYrBDjb7q6T9SdBJpnLmGReBDw
8C2Mp1F6nguptJzITDWfKpmIIFeGXYFOLKzu6qL2eWPyxzsgPgcxJs+rHJvSiExn
tFBvcz0vpdkks7Cf0z1o9y1L6u2sRmJzXeWB3r3wOEOiz1wbTF13nvyOlymm/YK8
FfCXPTjY52f/7pVhUjPr6OArkXqVu+/4ngqzRklHvcFUCE8xvWBrvn1vNauY3K/o
Sq7429IFPdR0ki2QeFgAyB14yOw46D3GkFoBxzzX1onwL+eVMPmQ66/DdvRTfl7y
YX+csuAJn7qhLvqM2+o1NkipKzY0Nocw23NdLeiMa+qgWn13/Z+b0oqjK27nLnkZ
H2Jh2USs0MyW7LzYrGJNrtAMcde8DhpVlHUF0FSiOh8gNmpHfUY3Q5vP4CgJ+tlB
Y5zYH+PAXaTk96p53MHvxse520BoaOWoqbjk/woAGh6qi7dHNEDJ/DhJPQcHzArM
GA6Lk0HFgDEb4MkANqf39T68isEg8Owy3N31cq0qRFbiLM1sDjIVKasRQW36rGT+
jaVKl+F4q+mBqcyMr5GaqvvOPKh8VPM51iuLQVWEf2jiAhm1fFmi0CEgUxVLaOAQ
/PrKYfkKHLQtgEEEt+xFG7XQkZTxGOTR/nd87E5N8CQMlhkbJRm7zxAVTfkjIgS7
CWOuHPU0Pw9CuAihKnAIASls1Xkjp+U4dm/PvBgTKJ01qHIIhfG3EOOWcNAqkQ2r
+h2ASDXUhbTuoIE4zlDB1LL5aRfjR2YuDt7+KoQdBTQU8DaPmXJHFh0G6qRXX8q7
K1vDVgHMrPMw2o22tHN4tK8sZl8QEfAE1DxfdLMFnaxlEQGFMvW7+mKLHWlnsWs6
F6Iz7xUk55J9u0JaCmnwUFFHJbbmsOH/8DQDsheAO+m9gChsnnt5VAbkfzCF1OZN
tbyA1xdahcUZGrnEMKbKeFkWKCU1XEAQDV+sAfLAs0TImdbNHd/TF1AA15GmSZuw
SxQS3Y1vTRutRn2eVdyrdGC+DGbujrR5WlxvnHtVe+1VpQxWAytckQiYr7V4S9E1
IwunNvlwdQHVeFRtsBqUoieDgkPWzSFW1x0Nm49lVZOboU6+3WZppInfKt+Clglo
WLbm3PawKwI4kIzc7Kmbe4vcDY0JiH2A5sX65hU8bQ9Z7PfqjbshmiAJ19usRmMD
m3VJL9JhHTKQZCDQaLKeRgNMPWDWA3o539gn3iBQJNo/CtzuE3VCr8QXkNIeur9o
/njGHLaZYx6y/cVPNUvRMpChxJDCtO0udP05bEDWKD0tBAKJ+i07cP3a6goWbdJD
iD+W2zjPoQBw8ZTk59kBklhMJBufMAvLOGDbn/GuO9R70Yb9Ey3ak9HoJkdC/+Os
8LFTYGau3BJrVBjSuvFGpo4PtuovvjcD7XgcMzyYN6wrFPoCHSdKVvtI/MgeFSNp
88wZ5Kk9CF9cAKC0G6UOeJ70sUs2Ot+jvzQ2mM7I5/KbO+5Q0I7drTLxGgUnhCOC
hZt3wz36CxrXpX92VqbaoPkmQHTnCeo0nAEzI5iiBrXfK85/N5bJx3Jv9EHbV7Cw
F/RsjedG6UXKNnTBrqsdxBHNddV4I10A7ZTCGublJdFkIKR3JWOyEKecHy7exi4y
5TOz/Rjl7//S5ShWTSG5SoEfYSTpbnL4bc6f7KZLLHOZUF1iCt1cMF5X6syVvjxr
rLaovr65+z5k3DycUDmlMoZiWKFIRFAApUhjr6wCeFZpV5rtAL6miZf2DokTokk/
1DLAai7F/m/F6Ijqk748yJu4J2anhI1jlbd5EZb43u8GhSo+Q6K5Gk1uFyaGNow5
+/GGoRgkcxuhS4cP/rXehoneRU0oYPPguKQj3yhYH1xYJVpMy4op/FV6RQgH3i2I
a3HhUUMbvCj7Zi/7iL2BLPcpGY7W5cq5TE19sgYYlA3OXxXu+aTeqEH7nE2hU2ih
D/6JVb2h2cjie3/WHSTLdgoKkLYMaCMDTBHoFoqtEl93hJH6G0eoVWvzMJmVM445
Q3xahIqlYU4k4KtIqSJdGToxwsPXXuMSbMd0OfLxddhTZx64j1Xoj00SIDCI6Lmf
EcYAdv/KQWC/9VFFRCMgv9LhYCYtkKvNCXtN1Y0lpC0ZLny+/LKXGBc0htyYDwVJ
Wm7DuqabS8V36vT/nOoi2Z47eIj9FmU0Gnr0pPiL+GLozQXFCtKvRm1UImojcZVS
cmhuS4L+LJhLvkJL679nTNFtAR7bUEWdrlbG81NTPlhOT8KkKBmT92DgVZz/FWso
biF4vrXPsvYHUo5lBTRB1nKawm3Zzc1gFZq6FlcBoAhT+T7XiYKFWhMpyPXnfi84
1zNL4fiUPR1m+dP3v0rTTa/HW7PBF3Wr/tcDA8ZUpjcmVDr84s2AUzPLPx0BBCiW
j/8inSko6/1tL8LUX5icl9RGcm7V6RybnXfcO31Pu5zfFZX5OqhyorsIcaTWZJKc
yzUkRglkO0XEwV2OofSUdO4GDa3IVldsUxQl0PIJyBXtD4co7qwtroHRoJyrpFXy
uGrmwTC60xUcwFycw+6rG1lU57cNULrnk8uz9LTAmgmLW4XioPm+F7P5ejx9lQtB
Zs8DRyfh9dMG42CvmjI6fOu697+BjO3trTCy96uQPmrNewgTR0Cq4B4frTxNGKDZ
AWPlPIASDCfitkI0B+qaSur1aPD7RotNFXfFQPx04loIvIAV6prh7VPTxatd9u7I
JEcZ6VZqPxzmQBe5F9ssHFJ4Zf60UuLTcP0MkvVeIf/Q5v6T9YqIBcCuTHXIfuVL
ttvTB0VeluEGdH2pcbW3wxLVpUnrbOx1VQ099x4JN0EFEJP+yTdZePZbmhYHaO5k
+h+ssKOXV3wUOjSgOkCqImgiyBdZjvX/3MI7ITer8yiBi47KKz6n+4fcgNj/yH9z
mc00kqW5kULqpwg2ILi40TJUVMYohRfDUUIvVqPSbCUfXgHYOu6/mUvWgLXCt36k
ErJE6/Ld5qfd8Xdu9bN++VDnReSoDXamzEzePQHoBl5uxNFG+qbuJGJYousgx7eA
QTPDm0X68/wPGkLxEtRNDQ8XIW24haxJoCL3eUuHJ3QVr9CAyCiYKldEhqk+4SbC
m0q8rxNleNJqd89s30nl2QyiXpo9E6qKyplBvAzwedlrgDqQTAtuWZ55D9Ehyt2Y
J+peTXsJnnArj64o+/ARG7pBo0dVCXyR1+3H0rhf1rJqv8VUYRvlbxIydVcWRzPy
GQoMZmt8NWj8dmHQjWYpCEdYRZWYb/kQDkZ+nu/HrzgSwW4aredAmaNCRmV7czSv
oP0JG/DyUB5Kq2V+xnTwx4mUAPZU2S2G4XhIvsGMSFS2tYVtlbfb/yftHXCuHM94
ymfWg8ra5oq+7Z1cYnA3ZlDvGL+vqgeBgIdQ7XzSQgQ8PIiER+X0N2iyNMUZBJ99
RwaG89717gftxRhlAaJ3G02dYVy45h4MA5P09dKtml5NNccDrsy19uIZnEhtIP3+
6lKidhmOELlZZ5+vXA4Ax4uFuijkEybambS0iVZposkOVPS0dcbvQ0X5j2moJ9YH
yzsPJILb3KW5muL3xsw2ukX+HsU5AKAH2ziIGXX+lz/uglVV6w3b7PjVCHfKqfe1
t2DTd7xjywsEanWxbRGScat3zysPZXw/p3dT9uPh5kUgQS1yR7nA9mwcvcqTlBoy
AckcbG2IyvcGahykpmIkKrd7JTloB4i47Syr/281sx3zjivJmimLRSm9bjT7iS26
qdxakI3uLvIATw3Mw5r0+t9R6yLBNb4VRJk6eHvXXRqycA+0cnL1+VZVmx+wTlPt
3ojnyQDsf6HqnuniGGwfdthyiqqkAD/VVFz4XSeh6paM4eYoEIFCYz3J5kbuXu34
qsY87Pv66LdYRGo7NrKHJimrvAbOVKVDHgfh120ZIXrlL3hGOxZoUPHiFs7Va8Mb
UDrYtM86gBBT+ICCbon0C/LR8QFTyNiViQmIhFSkbWz6newZuDm/NSivehw6JuO1
eddvtW4cV6rJWF37mXUOvrg6B+sNx3GVYvsGRQTuU76Wvk1O9FBkvVcrak1erNgG
YqOl4/mU28l55OBrtx6Lghqk7c9liavvsx7hA5EVvUno+3ZuADiTJFjbnOS1UuQn
MfWR2Xp/3fhG4EV3zS7KXy3jo6dzn5EwKOot9bscP48ppgZJ/SHfg5fa5abWjSx5
ZRwjhwc/fcIOwq2gfqxfPSmcDzzROgwTZReVckki8FSENL4rs+QjhhTBZgmIsRY2
uB7570Tt1lRJz0N2TpsI4WsLYIEKg8RwpzRc3w8jIx7kXNXNI6Mts6Vf2JMy/MmR
MO5ycRWUql49L3hej1cFBVcFb74xGH0B1rQ8go6s9wraRFUu04OGoIUkW/mXTUqm
QsqoBN3XlQFWmDm5Pd53MEko8vb4jP2XK/ORnLoy8+T0kq+MHwTcRzK0wy4heEHZ
jlGzPQfyCEzFUh6HdCPwBZABodvLZeordVjmK/RCfiOKJhNnaIfItyg76JAYWkLF
IuTdgU2fLLj/YFPl4WDwLyErLzz6thF8Bqi4Rt9R+JKgBRZMMqAs97yDcKdcOeIw
agdszk3edO29eH6yt9wx1Kfqu3dDrnIEl4+8uWTSy9/nEmJ7OWx8SFR3hd8kxcxW
n2FblbPQQn2cxboScoUG6WW8Xcoxi2cS6QC7Yecca1JLOK3gmrxKeotJgwVHbGGi
XNZjQxcowMtsLTEUWIN6TG8Y7pTplySC59OiaXqM801KyM1AieuwRVWTjJ1Vvi8J
KeT76N+RGV+aC+WomJa2a4afQ/7oMqnYuXQn+xpe0u5sA4l3nlGRrpd5RMgJXnKc
WCyCwOiHmcVO/1rznXo7/vCOD58VEUH+HZTKA2N4+4DTAEKlDc+HVOPtDc80ldk6
zyww6bCEhCkBiY4v4byK54DtHg4ETGUoDb2Wv4VZoGU6HCh0auhMLBjSXN0vQKC1
fd26WMkXXBissPMICCYNrAHdSj26ucO6F/z1VWUFMi9nsIXZp2tVkkvGkA1yIOXs
4azpdqlLcTIlKAzctl7//DD45J1KeINF5IZ35HLNvZN2jFo7DJ0n/xjVj3T8JyWb
PiIQ4WJeu6FdCgEcnFGWxiUtkcfnqbVj/jEFHmLmWfCQGYkmKiIFKBKmoIXSkskj
dLYQ+zSW3f4QlpEyQMi5vBkph81BEhJWQ++01TMFGCHAIzfsmcWPY5fHUy5QRhwX
L4ktv++JX441dlDmH6w0a1DMdkieVCqkPlJMXjju+p0JI9GI7n2fusipa9aC+ivN
g6HfelFNy71MBgYBSS5VA1I+XlG0JAm9WCI0+pBqjr3cr9/Ymi5p+td7EvDqTOt6
/FNH9xZN3cTnnV00gmD47QW7naXUOpA/LNs++y5QgxZ/Lp0hSnXtjTZ+T2l08AbG
BTA/OWaQI/ZFHr0MRy36KOEUz9NDYu2J+PoVgHX7QqKuf5iGiDf6/EfmOou9k1Tp
8hwGDC1BhTNRHVdJB01uug+Dba7Y3ibluFd6y6ahtOJPePtwK0CgRBcrJOjpwwqw
s2/KVfKh8xH/GH9q3vFvZ+BkedFNeTo9rNZ2j2Mx//4c9AzoxLYY9BtwOCaocQ51
MctVYpjyck0HrHN4wPNsE0iDEz6hhB34kZdYsPa3TMKjoa9GkJ3H0D+eV6EKKgJ6
I1a5Px8Lnwp7DzRVlFAzEfF3Mn6mjU0PPdNfNgace3VAZfH2ewRftq1aFDkHm+u1
zuv7RkRElEPFN4UrHbxmTG0QgrwdhR4LVHIsbfxQieeMEkNg6CHZhW/t8pNQtibk
K7SmckYdYCl5gPFyH38d+lawUY19bKh7OAY+m5CUA4xorUEX1bJRzu69Y5TUYRtG
kt0WQzaHt9nGL22awmiiAKIxxr00V1s0HVGrtyNGabPlqN1Hl0roKguc+IyaNlL2
s0wcq4A8AokO+0SD9mpC4JoMtp8YcIXkfj03g7p/m7tOSMToNZq/uGIKkoto2qLM
FlCo95ft5P0C4Bmh0Z3teLKb+x1if3JrG3C6jGe6sIwlt4jLfePc6c89m81Qs+Cl
O5zAUQhdBm9xZzqWkc4m8casMLmz18rg2tBhLfZY3x/Z0ls3k/JaDfIA2U1+JcJd
0MZDo0zBB+CcKxhvd/cv0VwcSoz3gI9P0Jy4jDK8eH7xqlZ85UcmPuWI+Yn1Ubl5
4LWD4qCF5WjlCgd5jOhw8QSU160IR3UXCukJMdproTmfoZQGzodzA7PRof82ivUe
yvJ6MLmqfTeshWahv04HW9prDqRMaj2tHC0TwVk+aQK4XW22KpU/ipcfzXP+fpTY
S/u9fUFS23AnBCQkTbgyPxxJ7n81wqHYRkgRosOcuczIk1/ieVS6VN9uTnEmUJMM
193e0Wfa8FIMEZH4RBQ3J+KU+PI9aatqsdrgaLzavl6vj1m4sIbKpSPdft1zjkYR
DGLVWnMkoMGU5ORQCPFnehnN1YdPwEGDFJxGXBthU8d+8+FNtyJNUkqwvDiihqeR
FNzTBXFRiLdIqADQMK/QQC21UYZ8RV5BmQOxa549SVsspC0pMGoROCwvxamXFveU
xI/SPfvEGAsVRU4rhCrHuJ2YVBQoCVefQqvtvV1iRjH1dHhWZB8wzY7Y4eXur0Id
1CjxjMaT/KU8sFkM/P/k6AHM+xNCYpG6k/Gp+SChsog9zo8EEuWGiP8TcUHcgFdB
5t09//cX5H96m/Slah2sI/dBY22H/SSOvtfA3wcFT7iGmOvUvaCeL8GobErQECsn
x2262BOatfcFCLhNT3UkEFYme5ZizLQBRruysPhq1l0RUSs/nJLOezbzEC1SElBJ
qyKgfbYx7lHFzvmRIEf24irPRrekHWNjRZnXIQvy1cXrzI8bIWzn1JzUkD5qZ5YV
lNLjKLknpNUCQiehL4F2UxCQG+hf19LCuphbWLEF/O1HVUyqGkq4/JQn5FyE4ZdJ
gx+qyO50UVjkpGJMe0LUoW0veyJejCUm1562MLWj2+sxsAzQebnmsnhiya5V+a0U
jc0DwPHIEqxkmUtpCIAiLddmwnYTeyyO7/V7wVVKmKl0bSqVUbFVvX6jgGdDnSYl
PiNCLRwNNli0cgUtlB+j3O/3gc3HwoYX9Gj+AisJbeXRSV4zhTKyikNdWyrQYFHV
4ecWu7Qx5g9bITvIjfMKQrJ3zQu8c65Rf72iGjs4/Hnwt+P//QdUs6WfO12Z636i
A4plsMPuqFSkMdX5UpmWjI2aTo7PWFLVRaKGuYaKBYmqB0NrLjrmbsvAxsF2KOwm
5xZ4cGySmgedUDeOjhZz/KCGsStIpp9/jF/Kt4YiiHJG+MPovMVIsGk8poswVg9t
Ycsdbio/K7vmSuTS5l2mo1bq3KXyFYdldttkkoLPjDbrik1JiIf98nzmyRMI/XIx
9YbOkz8Qu/ZwXwDenVGYv4ydeAqrQcgeCAmwMXH2/8DhWEjDxYP6g/0CycR6aARy
d0pFKyPlfjpjwqCN2Q3A7L7Kb2piPndG0y9FaNMojhHRW/mYAkxZrPtsjiqv8ll7
Jd99KxELUDWxCn31isb0Ogf6FABbqQW79DtBqh+x1uQp5kKBHZnK2Q8K4XBG5iCx
BbXPVqY3n0L68Elq6FDWGIvrRONlD5ucw3/6E4we88+x/FkQS9T17uKsq+O4bCSe
UmoHoSM/7Ypcy6QZYkoEh8EhJc4NyB+M8auPVTQ3SE+MkrolRUtEtdTSg59RwADH
HKjULjJFi3TUsTEPWQWObMSUSlAPnYKlbcTk6gJW76MDpYJO22j2i6GBPF21on2g
rY1scGCvq2S0HjQXv2mYkDSK2MF8KvNsEoj0qI823bC2fnDdc61krqIYa/0basQf
bSA6Aya6D45fP1kBwi592mliAh6eNU2aRXv5RNl9pPrKmcYlpxhxMlJEvgtYtiMW
BQJncMTmnL1UD1wrlKw/AoFKdk2s3C1yrrrl0voMNxxefri0g9tA7BtCBmOqP4aS
Fh6IbJEOF4IyiAmD/fBEkRztV/tUve1tWumSBIa2tnJsDI1o7fKQSotSLa3cznap
jmvppNKEpOJ4L9T1k/Xl2npHqgOuiRZt7SHerZDZalt5K/f9JUaAnjKBAJXJgFt2
3TKX8wm6x+D/RCehOfDIMem2ZABBcD8JzM2V49SNV8JlBCjiakFzn9Hpv3AvDzLX
ZswOzqAO63EZNHSylnexAfP1Hk/lwFdRKVJotWWsa2iKP7CKMDVLWZpMlBUuqt0O
aIw/HiJcpPzxEedCRqrymuDHP5Q2BG49XULLMjZCOaExvfeDU6dC9RsfrX35Budb
z/qPFyB+GzcbJ0XdazL1TBo9ZmzpcNH1sRRURZephv7O0PpHlUIwSMsYxuMKOQ27
j0eF/Q3U+CywNOyYVASo/l7oce+BZyCc6vv5omtFXer22y81N9KssdWUTTWIMvlr
Vcph7wKYy8kZ6DWnfL5/CGtpCuHLOub6TvYwmDZAy8+NV9yu0pJ6iErWNLnSSbzZ
QiAYDw8x7gOsMe0DE/3+FetTWsgk94sfMgjEqj3qBKXRidRl3/gfqMDYsM3Ng2Ym
m2Ne6drkPROQpFR4MegtpzsoUXaFNCR9qPs0w801mkGCmpv/pYjMuw7y3SYrrX04
q8jb+yflePGjotLaAnqyCs+a/+s83p/fYpaxDKLaZuOb9oYP/BVkjmTEBGM/0XOX
0F/i3I/rdHEXtogexhm1uQMzrMRLywxr+wbNObnjpZCBAMo2hpyfQ6tS+kjohvrc
kkME7C4YiD0BnbOYyzvo+EIAwsbgOZGKb2Zl/G/mXkyCLk8JaE2Blo/olZGJ62Gh
5ROC3SYgN+YCjj/J9QFJG5fi+A6igtJh+jNxILueFUIONgFkNj62IPB69Xxq2gXP
bIsaX2B19zpZtBcTE7cDjQHpbCmTpQLsRq5A+ZWckYaiY1Jvvok174lWlZj8Fw+a
QO97Xln26RM8j2Es9jMDVNsyIFosucrX4POaOBuPUlOF1F3e4E3epRbn9+2HwVAD
kiTkoeNoW0vWvM3A1Rf95BRRb+gxVIv59KjKWlheHNxX13CEN8Hsy0W+dPi9FmqJ
9Cs4sPoVN7TXq6hOF7ecRdZLHwoXLU/uLPMK3b95Fh86/PO7gzKPTNFlab0Z5Hvh
SPR6HfQOyhYRNbnBYwSBmFGTlEPwdTNWUp9AQME8rZ25k82qDSnSl4BjkmcSAwUy
S8yVNYoNHWoYdKisTgqPtpgzwWo61FxGtIJvpI01/aHwEautuL8zBve87jOcitlB
3/py3Z9z3q+Hj7H8J389IY7dlh6d1bwnY0fu100/axoya/QdAq2lat9IQZTiRhYO
tTEEsVjNJkIICUM3hWhYI+nWzbbZ2WtlQ2q/AHA6Boc5dZrpCO8NwYRyknCXQBWA
MkEgeGX7AQYDv6HOqGR98wBLt41zw1gMPRmzvxOPRahU+lxqPdsEBovPsZMEhhcE
1bfyzeIzqgFdHiwVQYh/eUv3gL3as1dm4pq/tujjZxi/xnSvvrhdF+dpzYnBH7JC
pCVTE0LJm2z5e/TcOhWtoXNzbls2IVDYEGhCyBwjS/RfLFj0uj699fafoG47GOtQ
JkknUo9V41sOJMnpkmZlszbVo4q1VrBSiel4uS73L6kd3NB+o+L6kxw6eiMNUP6Z
NfVh2JtD+qcqWM3yHqxWdmbC3rxMvQY2qTBUUcqRizfTiwLRP13h13e7oIfPScWL
9q5SpAQDwLD6jbPkS8VyvUURtg7CGElhqBZERjKEeWMJZA/hDwnNLLZFQcJTmMBs
GSZQebaa7kpWvZaNQkHXkqIfoFxq+X5PJefSfVkRrpiexEn3sMds9Fj3o3LLFIaE
uVahb49iQacL5Ibnn7W145YZIGaP4cxqcbCEs88IrT9z+ysbeeTGHeJvT3Rjv1rU
gt1SCL/QuY/h3NV/Kc8RDNU5RekpCiCO7J8K9sU6r3IetGfMd0gW2Q6X1bF8536L
GsYqzXMItdlyZ6F6NytbSYfal/s4onEE8jNgo2h4AS8dOD91dGY+TqR6TZ+l2SYR
lq3W+V80kGTDKHo/lI5pF4bKFOYUL/2sZ3JXWbcCSD4MXs3640nePfl1JPuMdpF+
O73zrWEgs6OC9p9Xt6ZMOuMbVewaIvH53PoYj8VEnu5Mkj2fcuzbkaKZjq3OXBeC
HWAGPybgPFrqWIcRvWWGbjL1VCDCikGHqJHoZ5LfEWI7jipWkaMyuj8OWALMx+QV
9X7MNqn25e1JVpniixHfmwr7UJccDHpfoyViya00LY85nGXjz7c01b9OttGWnHpV
EZUxZwXpLY9DhZYtpWQPDzXFkN/K6JtGwUCNlokDns941oqANQh/8OIbR+YjGsg/
vHvADPIzxjJKFZ1Yhr3dbf3T3WG7S05C1QxQHiqDM++tkLTbxqqlykUzQdRT5TRv
dpq4T/z/fEAFLHKVKeiZz9YQxdtKJiyw/3+3gEucaWDIKNxdiA25UPzFXeYb6zfi
hk6uePvqNxcpKEV4v6hugYtrc4qUT1hE6DkH98N/6NZKs4Dxj5o0xYKfwhETFtYt
QtzQ5JhwFSPu98r9qaR62JSaee5sCwq2Owj8vZktCO4W9DOmnlbty6aUY86Cc2Su
eetzsNr5J5ra93XNaYMyxRFFQTkssbMJW8Jwmn7QKdf8+31/DLNEBD9H19h9wodI
1R4SX+CE+NNWGEdmfAq0vTz1dbVeWhYK/f4GY3VVA/17bAwMl0twC8ST6x6PUo7T
VazmKbrZmVFjNbXf05hZGnAyENXN3zlRT1r3D6X3m7qDUfwqGxAy7/OrfXK7tvXc
AFZbSN+sDUx6l3ZHbFD/w4eD6KYDvocmIQdOiK4Huq8SqCqWxqxWQ5nYMWTsoVgA
RDYaieb9rArNy7eismSP5zE7RekjmPYMbwPQqtZhEGy4uBzNnFL8ELkVEluyi/Mj
9lMpWuJs6krp8EOSLLRlZ8wKR/wvtPOQWYqO4jXNL9fbO2jOQdB7QBHEMZ4vDDaD
wdS4pcUUG/HBVM9XAVNTClIMEHgcsS4GCq6CIp2+22kfQ4ey8OJIYqCNfXbVH8LD
cXbjHD9bvmO8CfV7sT9bcwhfHMSqvh3/uj8XvLIsJklVyHOUzlVkp5QH4Xv+SVxZ
2AbkbYU/+8Arg8iWuHXiZIoqOBaapB9BV376BmUL3IPcZmpBh5H6orot6RrpBP2Y
2r7kgVyVJyMyHXdCyC6OlnFVPq6P3VBQtNv1FV4iFn4Hbns6+hs5dNHTRfbad813
c2Ca9lwuOjqS0T88DsES/BV7JEyJ5hIDozS53ngK3UTzf/IzB5uX5BULqQPzn4eC
r/pSYYHcxjH1csiV4tTAjvJFIEyp1MFr4cKmhd54drSGRn2p3G4FnBHXZHQJScki
AzypXVc1ZpGQSWhal0UiHTZgoIuIxib8PXJDO4cSgJwmuYfnVib0VAg3NJ8uXEUT
//t/D5LcvhosAfNmkSpAiTq2zWMRs+8hR6NECxoivF8r/veDJgE1RY1wWMIXy92h
IesY4/5qXa+dGW740vpcMnN/wE7NmED76aTbAkafO18u+rFKmkji/dM+33wSS6rd
ITdN7tpOmig0h1XBwC3WaSBaG3YpauMjun18Bj8erJUHZGGyGQevqNVg1oYT0sgl
74hO9HcyrCYvajDaDbxFxvweHX6jx5J4tQeFKrVtPKaeunSwRPMfPxgrY5JGSpIu
FEeVo+gHvYDvlaUDMnrXus1P4sZCGOkIkj8xNY+byVPMWZMkElMK91LodNHIOwyh
O2nqIZ+TleUMK1hH9pUF3Qvmz3zS8n7rbctgzz+S5i+2XjQdy/qlkNSVAAVRflCM
aclZtB7/myXGwvxma9/mFDa4ShqE+uT9nKtUJ+lMWd9ppOauMqju/VM1kZWeOyNN
BAbtb7j8SdnKyBcnqcNMJ5l1nOnKZxXmQp6HS1qjdDiC6g9B2aYbc/tDxdChKV2V
pzwBROBwmM+w8HYmA6Ut+iF/a1GW9EuLA86Ax5dzgCAedG5bSvm8AnRuB7BUUbRB
WJjLLhb0bk4UHRMKS3riDa3aXhn99v1xNHOsmDAEnh8wRMNzKVff5q4s7/99F+/z
9saZd6Ue0MbtZh4l9VXAFgSllksEydC8DeROXR6KZ5csKRdJkps6QxQ51DFvuCiw
4iRa55x3NcqLCQLySZ3uHv+rwAMryCBUoBK80hBeXaFNirwYOwq3zfDOUHZYWMZr
cSwmpIRuJ5nDBe/DnzRRam7dposnxlDciu4OlPevZu5OJGZGolQm2zwNfAmhIKvC
eNK1rdNxbcVbsUQjkkzWlxikw8Xm7iEdxlp2m68FFCkIfecS1ad3MUFM3Iitu7eQ
Mitz4aJsbSBjELUS5v6eBYNkVaepDirGYHlFn2GKORefDjt9BN2u11v8DM/tnSAt
lSGxJil2J6OOdF3Tg2SmI8hApduxWcRsy/uPGkUKjiLyLG1ahDw11gq6mB54sekD
r0E/KJXrTnKcQZOnReCAoY7RLsivJ9nNsHP+dcBQDNQyHUXp1chf0zdiUsWleJ6w
nUkvBtS/yhsIxwN/6Gpp4cOUFimNAfrBjiUcebD/CrYmsddHpyrSVCy2/sHdMAER
SoZFRmN1P292HVigb7mR+k3VwFrUnuhPRTvJuhQXXtdEYfkyi8LfnJOTrf9vASRi
uIIZMn8ekRWNH7vq5XIdwxCdGHS9i6g32/yBOjLWcIINVxA8K9xbqHn9hxmL+iyi
GwkdIDy6xZitk5rRoIwehukxsmf7mxS8avf/XDSH7t3vNcpswCme6sLznU+1rItY
huHIbVdtHui01p0vqahnm+mHLQv84fcXAkp/NduC39XxK693J6x7yiek/Cc7J2FE
ihMhhFT7xLFgv9mKNPL/E7lvzRDlTP4KuRnhH4/9mr18c1O5fwoRO4L+XCnGpAMa
tXLgdVvWcSSeF8MgHIvP1NxCNwrsDebaWt6sJiQeeHCNYvbYSac2fsNI/pOf9q3T
mYg17aCv+H3q8QiyttTUjI0AfoWS2BUkhctCoUvjSnC2JfMMjnxyAkYHLnEgvCQw
AQRtlmMUqf+6DnXtBwc9FfN7wM8SM9SbXaqLfRIcD00/SsAZvoiKBgne6kIclQw4
sM9LNeh1PqSeEKQ1rSkdV9b7SGWmVPcFaGVYBV2T/5cdKuGFmYTu4GOUO1qdL2dn
8qHBk8K6Q7QU6nzfCZt6PIR8uwAt2IHSZ6J3O+5UrQnEn1EGNJ7nboOb4mt6yGmS
70t60jXsNoRCIwXnIka88DIPyh/seaselQGyKfwP9IDB8rdfaoD5Ll8eXYQEK8Ym
BvZF7uSbWlC/D2tC3wsJoOHF0/0QeOGkhpMUy5f7AgHWP++eo0GvZ+B91toyyOaF
D/gjZDJt+bYgqL5QYkNtOEUpZ6Njz+kO/aalxlfuKTadrR25XTKje+FSVJ2MzdGX
kvI6lyiqihHVOkZIKEKB0nNrX6qEb4XGjzLszR4BFo+qvZLZXC89YKjL3HR/8mpQ
oF6qrnmc/Sf3fi2rQNv5Zm2J6PPFPxUWnCBSaWhHdBAH0kObq2LZUphz4SbEKEqo
bMOtN5TUl0xcaGsDuSS03qjw7JezZ6uETKSCjymDz+go8YhOjLqHNP7YZ0XtEUmY
ToF379wWdsCmRC2yiq4IvYuw6vlzRzvmrTjAHLqBLxQHImOvAocLOpFC2gDTCl/v
+dV9jn0z+MDh2esRfePkaPAtHSoQ4xhH72c9gFvRHvMfEf+vq10L/ytb32yXC/qN
w7aEbxXtIEjw3L0jVyK68g0uaJ8SHpvIxJL81qMzwtNnpvQEbefHHQNt6Wbq/c8H
9NunlCFKwfxu9Q/8J6lCvzTZbRPMLPuhpH61NH3/+nB1TSe6ft86y7BamaCevhPR
qYS96NZWKI4/RZw1DYYNYlrWX4XrQag4qUheBNRkFwUBK9Z8r9NPPT29vM8SyXCO
7iS4ZEMV8gm5X4Ks1f4uz+svgeKpO9NghcuC9B2UA+my0oVwBEoDIZ3r64RYx5jh
VsrAJ6Aq0Jj1lMVpMk8wVux5ud60D/JcPswaYJvvGrBBUPQ18JPFos6kVOatJD5T
0knW8byYz8G4xyAb8J9IGrKCTmeUZuBj1saBErXms6C93tNDAE9rE0cwHe7hgE4C
J6kLpx9nM2DS+ZINSiuULvC9aps/pvgCUXhfev1e/qVMbM48aKHAdxtz7LsQoOAC
k8wuDTx/00dLz2zxJjR2M045Ow+2iGn80ADFoLFMPeWwAs1Tf5O9O0BD0is/KsLW
ajJUQ4qZBcmAcQlygXCtXn0+sdYfdwWEwf7CQG+XQgzuVPeKFQtuo9Kgmp0dfBlY
isbi8Rdo/QqUYAjRJkru4qfuTnKgDbuHTQp+S+s6oPnYZbbxEaqJCe4epALap0ry
k/I2fK8IDARytM5/uycp4FxhzAblIMv/PQYIo0ZBvDAzjW0msvDjABJ1mdNBNnTg
U4houMOemqOvfWezKyLeJ8yRepXz02rdJSc03scLjIUhNjO5dqSKXAnBW7wEiYiv
zrGyQSylGp9fCUVKUGr3DLF9p2YY9cqDvR9cq+ZUYknLLKdH9YQ7ZVTGaBQr4cdH
INfPPLXBG1TbClSoxNswD5vFozNFQ7Ssr1kzEZ6stz0rmKluOmoh2j9Dhp/kYYaT
10rB0/k4VS2YDHqtO+qh6qyTHuEv+9NiYYV02Bc5G+qutjAhcFmGh8XiM7VYtRbx
zJG5crO9/bn4abDfrKYOraT15KzzEy4I+q0m5x2RmXkT2Vlpylw9fwRkuvTqd1N3
STyT9Ocwm8uW9exAbAqaR9ATNTMfRwLYc6RgPtZFUQ0fwu+84k2CujgMseL9ZBzy
wrD/s320dF24Pbo0JmC3n5mY4xVei7pXZ5hnYYqd8ayK0N62pgzb/Gbo2QpzAzW5
l0MlcQjfDq9CrdSunpWa3CvmSi4T7iA6hm/kYWz9S1d99wwRrvs+05zdQ8tV49mh
CamudL/qVtfh4QhSamiwxXV4HJVPTk5iIToRdvtSFCuRPVUH0Varl21zsKTnwUpk
l+hz2NhPEworT3CScvFuFu45/OF4O3DcGsLpTrAhnoOHaBwK1JW8gvw6KNdlw88f
qVTvFGEaKmTbYnLeScZFk7qQbxrmMmjGuyjwNmBPpwzwsAnYEONWyQ3YFPV5+BK0
4anMBjBAzjd8P5EubkIQdU1dm5PUMT/1HtvoDYjZaD7fHvoD1kVNZSTiq1hc/3b5
c9masAW+OqmDTGQRk1XHpBm7A/kf8QapomCnurF56dLcA9Z4EkTbcrWoNbjFpKup
SmczdEhJhuanWLAfFSgOvy8CYqE73HWlNSfDWbBIQfLfT+wDd8hyfS1Z3MyCXBbf
W7TlQhCzYJt8brf/1vl/L69DfsWz0fHtzxGujylWOLy7CQAblclxvOjivEHzwAOS
BdWKKZVzbI8//hIye2NFPjp7AY09xd3NUtl8QvMHFpVEEwmMwzSESGsSJyCZEoQw
rNAheC/D3cj6APVRY9OdyB8MS2sjzoQ3KVIx3z2glYHjNbk3Xo2yWBCVIuBd/XzC
+q+mvFZWuE+v8Fq7z7dLIzKEKoIfdXgKnpfgC/wiWRQw4NirDJXlJxlgTL6H8hZ1
rd98kRVl4NMaDSGJXjlKfg5yCW3OcH1N778niHVoZdtFzS4XomPco1Cvm9VWY4Gg
vQo9lmbEinIbtNjf3VAk3JVkZkA1IWz2sXW4+w+/dPe3DQCDtZsQgPRU7ClgMpi3
ljADM6zxVBGh8a8GHkclWIdIvsl/OJuitRrU2jqcVu9G7nRPE1EoyJcMI/pkcUXw
2vu55e5nPBbpKayMDntHcLntYjLVL2qy7k2Zt1As78S6yy7Mv9Lp8+PFOEu/pC+L
cyXHxN/NCNojvEW+dvyz0yO1mBIaHK5Y8ksSLckHXq5ehU3HIyFxZ/M/YywcfwKe
G1vBi+nfLG5eU281dVy8bv0nnOTzvOzFXODfp2vtU6mJ3zl7/BbWUePxj7EyO812
XRc4zq6cv/lH/uZ8qKzdwezpYT6pWUtWn8roW3TWedetdf/5SNUvW975e14qfhnC
phI02idCUG8X6luYlVO63DJNnMKHOkXBynrFlj/N85HcTuefm+an1q9QI/wGcLMY
fcUyPhIKPbkccwZmcUD1jAgfRgUR1BWs7iG93YG6iBA6oZ8KnQdsp/WlLCMLwR8j
YdlqB60ZErsWPYyuRoAJ1r7wY9rHY+8G8Zl2D7Kp65JQtmM/+ZcIIittUGx2D3IK
rs8mGmLhWcValO8qsi8OcGkpTZO/bPWjpzPc+a2d7vkIVEv5cR10cbKSLGYc9ET/
E9LuSqVffJCn0AWC72nphlHNX9SmFOH0uCXoIsAOtL9+ESscesbl0EqUx0uZBJ3a
NK+ZW8eAiL/J4LAM8cQvx82qiPc6IaZ2CdGBvFEW0Z7CqUAwLMxn+tAcbfiQ1k3+
PDjY/2X4fJDZ9Yfe4kAuPcox65rHvISBAz4HmLeHGEbHC+W86C9UowEoBapugE8Y
kIy3sfETn6/jExE4qRI9BagJhJXw8cV+rouYyfuKr/Bh1gB2vrosFy/NKPGy5akn
QV/sIEJFmS9TG9iukwP1m3FIlr7M2JMq8A4ad7UgjeKRp64b24ViBaFYQt0JxBZX
OUd+0gxJptPi9bCgtk7WfNBNPnx9gZ57bh2J+CTVDdlqQ8rUiCgOJy/tpyxrXfnk
dk6HhPVWA0/kme5c0Oqjwg9X4oTimlQl9ih/eVVM604VetQcrUkrxDP7PIiGOfX+
6nk3kfqsdoVuCScYTlopl4/ikhX4M4zYQ5kNMYbKMZmHyzIYRXPh/0fmNypyRbo6
BELYE21q++6GVsv+IHuV8NDGWc6/bSg3rpVeRfL6skLikfCTrqLCMF1j0AOg1P+m
rEDLw5YjP8W3K/HHWcNYWOCkHFnkgZzgghdmLquug5TBtTWHsGniYez7rabF1ftF
S0c8ni21IMlSMXa8WNdxMB7XM2ERrG1rw8vFcCT+RP6M5HYKr09dFanSM39nZo7b
x4L9PKKFXWh3oknCY3TNpLgm1JRVBAvF3pme2j4YHQr5DuVqRZgyLZcJ/uCLEwDb
MDY96msX06vbHKN8zJ/JddddBk8WsWRsQW8Ib7HfIWSCzKJ/ZqJUppEkx7ABnlR9
A/NdhxTGiezp13Hem+qhGCtqHT2C4P11iAQPFHCh/kJCZd2E41R6u6x5+s2+IqL6
18Cc5az5tJd6EtKWzj91fwXZfGSdWcH4tzXgYcHgAWU8+EaI7JlL5zEDaLmWM1Dw
Nr86WOZ2IEFWpMtiKDp2rxnWuLjk82yg0f2tvrEIAas5Lk/nAA8zeqrYf/t7aKvu
IZw4nBsyJYiSNE4PHbaDCj6QhDGXaEZUMTFpBqBdgycGVMnOEJj4eN9+RlZt4bbl
JqdJ0eEIS/CAQyVvoJ9oN7VA08rMyHEi1H+71sUx9qqhlTaaym0hKQ4itEe9i9Rb
hI+QfI4uOcfsNFCgEyw87ohOcEJTBihupRB5wx6PHhHWVHuKyZS5r6/GS5yWu3EJ
0TX+A+NMQFQjevgusmz1N7tDqSWiEa4DMbRzGhFegAlFWskBFHb7V2C57vDF/dZD
QkwT0aJaJqCRBt5yyZz4se4cjDYhjx1mf0menzFVpMdCx2U1+ciDOUkF62KSLls3
Zk06E5wn2iHM0HpypjZhkzjUC2kexPN2/wCtWIs9UXLwanG3RrTMnGh0C8sqwRWO
1nZFvMejTby5N5qc7Bd8grjT6OkqUXB3hPJTsYDixXRDswfDlEFRmM3aYDSvr/dr
10vlJVLB74cmXOTdNPdTS8/BxiBw6arzls4k9lIzbcnhGazs0nkFZE4xONavEUFE
ftyXnkeKYe5ExxiyTDKMLYaSOXGRcgxVUzX7yD1BO7dI0XmS+DSv0j+aDmcjwcC1
gUU75CQz8t7pKkyBsV0Xlqn16w/brtUHvXzQTg59sI4mIhji0qE+ZsFDAYO0UrNL
JWZUqAMDD6vJrMWsyC8BVznaFugiymgJoAIZdNAQzS5zyW8WHEzDleyxH6nsDy1Q
lYgM78EKS5Ro71lk6RYOnG8+J8z/DB/8gIuwN7n5iC/5n5dDg0M3SxXod1d5z7BW
VULw1Cnev8u8YQZXqkfFZdyx2+iCbeOQZ/9W2afC6EHXB8D3plCAglQvFLwCTal0
CFw6kJX1OwKA5VzZQqPBm5R3uiAbss7TQ5Fpj7EozmV/tWs1OeRyzgYjtRmbbAF6
tXktBQme4jIxQ+QjMuwjPT/lJ8O8CK+icEJT44xGiZ/vhBaK/DMS5Ji7u0FZtYhn
tFv3eTffqM/N8fh30iOVeqmfOBbRE95i2CZjH3O941667eYeoTt9WPNhF1pDIUDV
8h+yByrztraZStGn5gwIb5667+8ba5mt8iXRSx1dyHZjiWoLQ1T6uyPv3QVzNaAS
1UE3wo+lg8UUnZD0D/lzSHwiWCvDXVhT+vYTEkP+MPogoZHW/fd6BMUMY8gx3LbA
JlawGxvDHWpcIRWU6hTFHYWmMzbB9wRybFf2O9Ipss9PRbdC5Q373cPuHO7c0b0w
bgKjwRx6uyIxLKjT3oTcshb9VbVy4hvQt+WWHrDliPsnNKe7H04TBsBYqVs3GM8B
0sgr+VOlcDfvwTvRqeDj6n31WRPzMrp1jefin/yOc0wmASAtA7WDBteq+hn8o0hO
qO4urjQKWy9ygHB2btX83Ji4Gw00dreCOrX9jvrEQC1Zk4sfvrCTXL2skbx32bHn
+SfcJQwLfG2IcFA+HD97xVdP0RF2RrHBtr3AZpx3WL8KSjxvaFY/CqaXV7nKduAA
BTv+rMRe1YvpiDx4hEfL1kIz+bCfCyqV6QBSimVp3Z6cv7pS7svuEwo8WLZxFKE7
5rhTbvsURtNOljt2S33tH+D4rZU3noXzVWTe3Lg1CLCNHBcIDw74Bm/1Ae7peL2f
yhFsPSSiysXUJxsze7UTL+IL+neR9P6Dh12pY74gjI3F+oLqhCtfl/TJtgJVcO1n
0d8g8es3oAlccnEc7hR0Y7lcSYHsgbHAqTiZvb047Cxd5uqWKOXYKu2aSgVwoWzH
Y8A7GX2BM1BtlVHaiU74CXoOSkGJ+TtGP4hYI2MBxKINfMWw9pjqjgvyIfYijH2i
bjLgOTCziMPKcGo05GDqXZdgsRxbkYYdG64LuCshSW2Dt+2KrbtkasJokAPDrkxO
omiVCtgxie4u5bVdkqeLkXFkV01UkxrlOKtj8Inbu1sX7OvMODlt3lVQd7XZPbEc
WrTallaRT3c7wkdCCKAno1jOY8zcChooAMsqfM5hxOUrDwf3lhXrOk74Sei7D5Ed
WQsdYaS2ec5wcMsHRGJgZDMOJbpry2q+lB8841hCvVcW4fAlhfi8j/5iURRCnskv
YftZEz7N8g6ME3WNABmEQ50WRf1Z8laOE3cGnBfYqV0pHuCEMqwUXdLGb2uL8jS4
SWy3yWSFmYwbTemzIIxI7rQpfq8Vn5Af32QKYw9oIcMfuXdcKEdHGFTEdCR+5FfJ
xkB0rw39MYmqTqTC6uNpSyqC8PaJNi3Ksu/7GoL886PrB7PnQve1O6a3h1NMP1N5
olsqIMZWyQkx+9qipWCLlg1VMwKsu58yF92EOvgaD5z2gqCAvDHshay5zSNSBcst
RJV/si8n963x5qJNbGq7yI+uSlt5/FsjID6FOjeWN8QsRgnsLOZ3PN1TNn7lwQkW
pV9vokybZCGdZ6ndzYYIjZ3Q397P0osxVQ6orHhvqHc1M/urUBlaj52Gd8U9drBo
mNJdKYbOka8NPR4zWPTDMEHFJQcH4odA3+U+Iv9ieuBlUVSLLhqALZraAR3KLrBe
kiV/KZxOW2t7+FZjEVTUdLhVp3J6Vxf2oZbegWkZzJpHW2pnxfbwxibJKPiaZtcB
x+lInQ7xjiyjOO+CWA5AUzVcD4fINteM1zvuiAPLzKgFj/0ovhbR8YXhB6+ynSwd
Zw74wwGNmgYghpJSwds41TyjcPPmy8/D5XDwHbCv7K6UAyAtEMTVmFwjRna1j75D
BQd7RpPZkBtUERY5AbzzNOWKzvHKQikNpityzpjMUe+zxmGbDS4bTDP8Z4YnQ63K
BpvarYjRQpXZHhE7L5hKxwyoDoBCmBHto6Ayv/Yjv9KAVtGAyWFGSfNMXvYAQFdw
XbkCKF6cNOg9Bt3OrNbFpe4et/Vqd4MqK3+S2T4X29vfNARStihIILv31XBh74Fj
M6TFuhnFt5oaWV1gko+mE+pDVbUYOHQywKuPwkCxpFbBYfkJ7pzfq2+9yjIB1hxq
XlXHgRK0wCAz0DJGpMEBFrYL/gC5RXAPIawxfgvUWCCDa0adb/rOXOc1z8xumRQO
4zKkEvReUwriJL3rEk9u0v5uQFWEWCYeoJj9+PfjUvYMaAg0sKqze11YtlFdfqyr
Pb32+h0nMPWsoZO3Uuf/bANuHRbhO7qrg1S9mrtIRaUXEsJnED3BoQZtkPp0Dm1O
dRQMkql//cWXQxxPtoFOWZT34hqcx0PDFF4bAOW0wqLAeFtSGW6uYr6o6VeJhQfy
9lq97ZAkVncMye4ez76ySRoodG8L0HZBzRfPkqy/DiQnN6wNUazUepkm21hjsSvK
nMPvSfAmQ0nHlbz2HQwIoYO0q9RgRfhfCltX5OiUnU++Atf9cpCXirUnIXtX/dkq
dur8vIxjQDD+CaF8X3BL3GQnyAVxUrG6kep/aiklJWm/zYSS5DUNVEHWwt2ZYx35
j7z8y63EIm4dBjwBeGw0ptfalTDnhpQrSLeSGU393DIpThOQKsDfnKSpHspNUhnH
WAj5/HM+SXoMCtXH3WpbuGxq8j9m7mJr8nyZ3zB0xVWp1a6md8mKXQZ12bp7OGAi
O9+JDeYIx4kvGBPzulbZp/8ddS+FfYLN+9+vIG/NHZtP37fOEu6rTU0zPc76+drZ
SdDsqmESKcVx6KBTbzFKtP9H9TB0EvlNTspt/UF2/j5Bd1uu4+DqFL8zpabC+/sw
IKw+nAOlJZrjSSK6UiJe4VDiX5OwJ22CyC1MITfvkbkWGdaRMxt8QkOtqsXzrE7o
cFGMFMLrDzKwrxpCkMcxMWbmsHSFyhXbTO5kcuDmOhivFMKxOPuJE+ZKVCcnHUg8
S5/DJR+Dsxu8y0T3lYmdzxnkM6nlCuiWpNYRDt9Gr65XALfE+CleaCTnooSP63Mm
10R1+ERhk3m+ZeTqRxy+jlsKZLhqbmbfIsF/HFp4Hz/hwWxfXL3MLuQKR08hXyf4
/HRdzpQZaPN++q1X2Kp5FLPK5jm/4NfZQx+6dvGvONVl/yoL5etMxQhdjeUE1sq0
XxJONbsZwb7Gd/Pqo5eqAndDMZmqHRJMe1LrqRHAEbbE/yLIvcd/Bfce0AunZO+Y
76c2nWpIwGbMGFmndQ28Y7JDYNZ+JOAiphOr8FD65kMDBAFj6R1fcbjDh6RhZk5h
RcciYObe/7XJOmgwTL7K06jiHCGhcA04yvzuj7UVUIIgQQdgfNkdWgc/rn/RW1lR
XBTR8adU0v1pMIc67dwBYBsorKJR+RAj9ouSSzPCYLKSoPcURhX3z2TVKB2NNVny
lDFQvf9FjAI6fJ9mXbW4ouM7oI0XxQXIf8aVcoHBVQvuq1YO6rGvKJEewIe6EQ2b
PnH8VNuHVRuzSnOyhmtR8yUoTi9uAGY2S+GqP4tGwTwV4p4m+XECHS6uPibu9+O7
2tfID6gcoPSAuUsUTiPT4LhhteiMZbL+5a4ihKqLBDJTorpA7KlGI9hIourArLPq
U2AD9GoMDY6r5w7jbc0SATRivd3eAdVfabU+cttvvaFQqHYLVTxbDoIZgQ5MUr4G
FFMOwPdmyyX08MwOZsnB6QhnjGrn4e+fx2sxHhOxEc6mkO7c1nXECuSZHCOtl16q
UbHpBL1qnSnJ0MtFbyu93iOhotgYTDGdRCULkqElMxPgDWDIBJ47GalTQI2/urFK
jEEHXmfuBay8JJ9HkOcW2oyb/8BQ65PViFkk8FridtgCZv9by+a6i0IT8UbwfiJX
tUb3masw/xVTtuvBPySG5Q+Wc030PjfgGbicZEDWneq+y2qscmeedGF7UBlbk/jI
76WMsiw61dzDNKDVEgaWtWEqOsUEMQRNeCcF31jvuExA1XRlan6X+Q3tGUgIV2It
IzjaVzS5QuD8+FT8xkYcSqFT+Irc12PutNa/at9n//w6MxHgs6HOeBw2JCbVzD1b
hXuqUUXykEC7RkLQ2YXJDa/CauA/fGoCQXInVs5kA7t1RhXkHwVxE0z/VRDRB9CO
HBr/r4UkD230bI1XtWmdhrP2qZCU4pDQKvEY5qeIhl14ODPk1+dgGI3euUvUM27+
wjxDcL89OVIcMjUIbFE0EG8aTNS9YfmCsWOI9JVN/O3TXEwjJHw72WQNlhIjz9Oz
5PoKUqaL6HXiXgaPHV75WMhMw+SG5XDYPNQaWZUIlio9P8nz/DB/a9G0pNVc9Qm7
rDbPozStckVI+VROGVsIt76OtBr4TPyIE5Y4NJTUMCPL8zgppQs5XafId3KFMunA
LDexoZK9LufxbF2uQ7lDwcnXJNAWuzfSLPDrZn/JgYGWi92rTFMZlo5l4o1GWpx7
JL7zqJd6HqlMUyBt9qyrvHRZjWUd5iH/M0aBKQhytLcs/CddVAEG0y0egOzRSriG
VVFR5traaKZVZKo8HAMlzUgqaEfsLAZ7IauPZIUhHkQdnS6GxIzLCvatg/HGd/2d
c9/bRcw/kZbAt8XGoz+Ush0f2Vf+zSIv6HoUs3BtcqbwrhZ50jypQrHplmnbdln6
G0lNLaZRvsWy24r5RDJZYzBXSnpyTGnwf4SmWA3u41nZ8c6UsokC4ZrVj0h+ThLR
rD74d0gY1OgFU1CHb+gx28Z+E6kLVcvCIDjuZB3FwgX29WbfAjCfdVxum7DxJVul
qcVAQ+UME3Wd82GzDR+cVFGOnMur2u3ZFOnJeh65cEbSqGitA4SYkE7axbJkwdq4
Uz7kd81UsvtLatek9Q0f2k56kxRxR3u1zmXjNPGc3j7NgWhotRteWSYQqAdWj2bO
1339+j1hFUUWL/iJGvLTgxJVz4at/ryb2by6sStaP6x0GijNM7oghKyRAH3xo1kV
uwXD4et571KvNmpeAnwJGKVwWiQSXsVWb9XGoRBPKnEBzt45+QZLVApSy5Gh6zJR
hKOQWipCDHz6OXFe3kia5NwckKK7b3sBZwATuTsITNV5VeIOfxUuYZ5eQedtVkba
zSLyVpnou4jMhTdaXbr/I2Z4o9sVJSYYWu3kZmXJl5uJhE87QOG1rf+42N906e8f
079agWvfBGWIVYHf+TKk5u2SutW8GJt1chAjNlU9pge/Wt4Jf4JcPcjVF94Yy43M
xaSpIBJUGKcqLNKnCGk8vPXGgzF6EruoSeVOr8ctM7BJw1Kcpu7mycBkm+5TD0CV
ANJesYqujfl4g2bYkO09VJpJWRCdaRhZRwbsyoHPsHN3OMFCYUchOPr2u/YEkGcA
AO5JsWyFIqn15kU2kAnMnjQ3jlgqK/4mgsAZUY7CFWx7rvK+T8SU8xkSp2oQzAjn
oIJE/BAqLmnRL0Jq5FPcV1J6sKlWsYzImvRxE+oKNBjvPqIrE6Q3STXSJ5ClW5e5
3KNBgXFludGgv1RCCbEKdCo7YRtXpjjLiRd9Y8B5YNvFX5hP/YnfZqh9eRoliMB4
ko6zBafiZI8MLExGP4Cewg80xk3btiTy08e1Qt6AqpIQmpKuOoBLe3TSxFa0w3tk
a8MkQu0W9bTRMP2LxPtX7z02hEpLZwUjCOxUXOLj2R8daVo+mzpvyRK1WY1D+2Pr
zS40l9BS+AgV523QwADhnVb5Ore5Hj8Z5oGZy/PGA6PqH60cucJjnl0VcSfBI7vw
PK3LLl/oIkcZl41X/9C/NEvIcd1pZSHLxglJXcBLE1rqHVnYPpd73V6dfY/sWEog
C/FYR7J27A4NTFKsslokM8/zuoled1ko8/pYynOkSEb46U/Ao3RTE403CxHGE9n/
upt4mQhpC3TdgQw69B+aEyslQf4KgEuOf7msJ2JTDflQ0xBrbc2eLVTqlHuWnrhL
8wE2uP8a7aQXPTYO0tWrPBa+4vgLtCHhGWktm25H0RrRhJ5oWhN2gPbg6qFK+gjZ
fGBElxcC2qlaJztnAdCwuGN3Cg4RuZNie6jd6ZvZ8ejngbygPeVPdxb/agLGaJHI
lAtLK45O56f+PvnTueqzK/cl0FZAZY2SXsG9utZ6VyV4ZTLg8rObD4b2absaM0lG
sRRi8RvHIjhGs4YetA8sd83vBjvnHbNn6UUJedpz0+G1x48GaVn6o5zv8SUNeeot
sHZmsZesK8vfNNOkBpBWwer5e/NQSxR7OUCbawMJUX3m+AjS9hiuR9dW4ZDFFP+K
kZ4IaMSs7DmHUAJWHzG1nJBBN4PNRIF/wI1j5jKNFQ/Rf3j90ltBjhaQZm2Hwrs5
ez3P8fcPwN3HKPArAfecbnHSzaJ2MpBYaeo+5tg2PFLtBwKRBZsGFiQ+USpvGDea
vCDSwOKrofx7Zb8VBC714fE5ZYFfpEaA2wPxIqerzGJtnG2z+w5MbX9Qed7V9b2L
4dp7KrrKOr1YIUrRap2N9it5sFtw4BS+98PO6AosWGPZDHewUao99O0YfZKC9sus
t9AMz+8Vb/YVSctDIJWCwd5D7WcbxxOhOQxOqi8nVAy1/sRkdFW/zX3ejuAM0Xgw
RZbQ988SY8nQy5jxgHwiosJ5z0icDLDqi92rM/8fivmlDKKRH0BPXtd3XrOKvoun
0uATzKKAFGG9WoefwhF1EX6fOXGwAyTZROa2VqUEDZ4eo0DZbAf6nD3Ta0b5b19e
8bMoqy2ihUnVsjaj+Z+gmm+MARjf8VqVxtTR9rztPhlZVGKEmPUne8O133zoi3GA
3SurUGLFptm04D+mS4ErRoPj4MDkfqgpP9DGtxfg835OScZ9rWHchiq8iqU8xBD5
q/c4PfqnGftFnkNURQHIs2+XevELNqtU++Iulzn/T5EGr0biu38RlT3pYXy/XSOO
41aFyvVNafj2x2R0VAjDg0dL5HMndeiPNuuoDm6mBosnRr1MwE3ZtKkFG8LUOh2W
hXVlbP1u8BQPHTXISkQyQbWxop4jrhVEGhpSfYVr8qd9WWKs6dX0wKYtCRoyndwB
cz/13Nk2vFTZt2ASh5U3tMDOdE7+N0tLC6ezfBJceKwGJt99Dd8U+fmjQI3b3AZN
Hz7pAPAqZci+xRhTnuxPTUy71VmQTiluEletyCM0DKFRPSaL5+1dG9FoOvbT81gI
LlWD8k67Noz6OKrClcDG5OPX49Z04PhMgyQkz0ufM+iLymYZxSvYjuZ9GmDKrch0
u2ET34T7f+Ea62Fof1aKifG7Vvf/syFaz7nINqo/GdynfKA/k0XoVrxf/sKJRh+d
T/d5rHX2tlQ1+qxsGxpNos0gLQC1ZNt3PRVJ7aJIAcPxCrsVEBristz8otPwfmBd
Gb238Y1//ugWWV1dWzaR099+n18EkX8/haNUkP0tq94TYcyWlu2vRnVySez9VqJn
LINuPiy+V7//dZiVzrcVn+PHRnfhpu568zbCt58m5U6LGA5W7Ac4fNTIr790H4Sj
n067ksZQG6zIMhjqVp9wvYZCAewMcxyYBQ0Rax+Y5CEyj+8zgjQ83l8sNOyOIH9b
97M+N/hFe5rAgFs3+UJ6iKMcIsvCGrapYpFTczCJUNM7J3EHOSnitmd5X5Hn5+wC
7l1fb8gwPxqVHZdWwc9nC3VvYot6pG2advqXMYphh6SZs6BRWdogsBS3MD/CaBJ/
qnYokyAvkkcDJkXKslLHX1TS/dcqA/ex6ymlMzfA3VSyAiJb4tTbE26QjSRFKDEi
G1magPMI48O7sNE+vLyKPKuo57LnrC75kLWnPwSjBuEJtkOHkm6w4s/wh/39tlDL
O8yb3vZEmTFtYpyzTRcA/MHeP2GI6nb7d68iDoH4Y4mDHRz5mrBQUyyEPoU7Ggx7
HON3brBgK6AJzPxji7JQJ3I57iNC1IVrjaqqUZL7Fh4cvbDfH5oH93tyQxSyu6Fv
RgktSUGBpnzt/ZVtYZw4IgR8AXManZrErOjeCS1oQD6IbjvBg9tNCgC3b6pK/cbK
1txo9+b2yW6sBY+D3nanlAGZ1BIxTx3UklIiH9QR2g/v3D6hGW4ZkGSp4AudDiqb
DzS8yx0YT7imefPvy6PVU4mXUo5pFwpWXUEUMEz4VfTRHoNv8yPsslrmXrRrum95
XIvMX8p+bE978Cd3Hu4+RJw1fzjFE2zSVaohcaMDAawzYLnvjxV8vpK3TYhIlWjE
QPB9uoqG7VmTjOUuTXQK+m+IAnZ+MygouWGX2q8+nsGHaneA9dHr6KAgLXgfYXnS
ikjFkXLkcZ5So51P/D0gAJ1h6f+XqyXaTJKDVd9BRtCfkMK0ZTdWCwTvTQ/K8OWu
9XVDaDhyup96qltK2+HTr5sT8MbY7TxwP1aEkB2uBNVcB75LDhp1V0jPVkM17bMV
6s2wc6GjPp5zeraJ07/PqJsuXg0/P2EdTx1pedMVUfbswdYEo6iZvrx2zGfcLSrj
Tec2kY9JA5bwVJOlbT5SMBJhGUkPGFIRqqxV7ecWvSv85WGwX2+jgNQj3Vbh445d
5Vo3knYcU2YqxXsmrEreHu98yBP2c1+m47LLYa8YpB6nJpzM5xbvIkk+wA9pohQT
Nj/pvWiDxZbJbRJ4Z3J+ZY0/8RjVvLBi8x7VjkOLKHiB8qH33b+x8Prcs7fU1uLT
YOHcExvyeMhDNfmHQzCHoR0plst4YKt3Gjk0koWKfQzVh2rU6wt6WIJMnKD5cFJc
/E9D9pqJLpEbBuuB3SC7qYdoj0MsTE0K8Zi3pOkDGqqpww+sBQiddGnmq2H29fDf
s4+Lniuq6XIZLlPZfw1gfVnBVsMJ1Mm7hsfusiLNieedZfg/MKamELIcgi6DoaU6
7nbt8I2wy0wrwjQHzA0aEnG0K8I4CHPWGdNDI0F4/qJVEz17xs696K+xZYzC+SsY
9optW51OjZTmauDjkqfm2zd+lCfRABIpisDIGaTFTvdm0jbut7IPBudejDyUzkz4
8jdFia8D/zDlQxpSfeV3PUXCdCL+59AQcr4bASMDCri8nLHoCGFylseIbs45o/jS
IbeGaHJ8L1XQau6VCaJjTB9DtQxKXx9mczJG0nzIUqBBSMHiZgaiFm7aK4pV782+
Vbi/72m70W6VbmK8dq46+n8kfuR34HXkyFcBVHZ9axXMv75E2Kzb1fd2Rs/xhZPj
2+Klck1rlZ3ulr5ehxnIvYOg8WE6vxxa3SqxkaRAEmeYh0zKvrABujjgEo6hMtIs
cwE+JJMVqftgyuCuHBdnZ8cnfXgSZNeUw6Zw1xjO5BD8jTCr9Qi8+4M+ABpvySpz
Qa6J1O8TXTb4geAz7fmrmqxOC27li0ogr2eR8+OabaCMvW/i9CN8OyR0NWwFNddK
TcgL/OCO/2rwy6ZZugnHuOmJOZgIq8F9yePfiNiqEGGdLo7Vg3AQRDDt3kwbNYqE
VsKaVyZRqxt80mtDNMYJFhZ+TrFjfcmwkvcgl9ABcq9aIWB1gk/UE7P6Nqi5765L
XZGy68L1ERlLQJycbfCjoeQq6unGRR1CeoLgSIXaNoY/WdnqfNr1ve4ShZi3rsjv
bw3otig24eD+wJzSoi4NWOmEh1LNviScUzo+UUGIumRFl65tPUKuGoyc2gFW6l0T
1eEmrQmjo8bSm8VpxHphkE/KFMcNgG9Y7WX9V/yosH8qZht4Dt4pFnWZYmDdq2IA
BW5N8JDDaSfHLiM0EVQILNEKSnVBki05GfMTHp1bP56dfrU1NHgLPGKEZ1Gc0NRq
sAjkQzf7ACxHiWgcaoRAmaevLLSExlJ7cQrt5ISiOoZIQi4DWKRmtmYRJy3Pko16
sbBcRfMTGH2Xjvs76ZWPPypBI1xShX88wvZvlzkyAykvX2qb2vtkKIWeUY4F7SP3
mBjn02KdgU5j4WaTnDuiP0d854yaXf5iu52D+ZKddMAgLIXGLZ4Lo11XUtIQObXs
F0HEjVcarFzwFVi6iHEWx+TqgOiCJ/gT24i0JRni92b/xWbkEPgvcTWA4NTqpHfo
5CNReSplGqOnnR5J154bu/0Ql+fM4DczzqGJkZ3LrJRqVsmUC8nS/UN52E2zJsU2
xN/12inW2wRwrzG7wE8e8qzaTgwXcNnpG1SxaIpgnIYqKdoBl9pmduSdbO9DDBtk
y6I2Rr3Z+2BuE8jKTneajvSrjpt37aFq6hFihOfOXQ3T3Ttf5G5ISG3a0MuQ7YhV
cIl75jIN1qoni6RSHCFepe7UEuL8UYw0W7n/o58A+60ugsOk5vZGdaeft6EOr+h0
EeMJbq7iUYKe0UetJw2eMoDGbdHN5kIxa1cS+dGvjypI3Sa0jtF3o/QSrX36dFVq
D8pLLWDtZYs8ihvPdB7PtCSqODLW9kqFhGJ52XqSh8ehrxLjBQzGWaFXc0S7nT1L
uu1jLh5e0ahMgygbWslIQ/8H19xLOpUVx2qhiZJz/04NefVEeuiY3bBdhx2qT5zz
BQA3fIWJuzf+75IjvF39NUvgMZ5KpkSKGh7xKoE5a/pTnxnGKgXg80Lx2MInev14
Qt/0sSi9U8TZQVnyPwKXTaz+zHi5kqOuMe6vKb1u2KavSAhMDSobFBnlPF+QyY5h
8i2rIDnZiMlkV2Py3+bHsDDoXAw4XwH6iHVZEMBcUQmEc/WfqnuwYrF4VJlnMKne
xMlMF8o/A2hOZ0WE2dHQ66NvmQJDC8HSpxVOSbynzAqpzKucvyWzAj73rrWDn1/A
HU5ibWhGRDpzGH0+r/SelfKhCNNrbdRQ6r/QTppIVsBGYpuXo9vvzlS//rH+Y2X7
ZvwoKQ+g+o0QxDi4cPuvoBzTsjKNRo5SqpHdWIk4QTHbIAkkQaCzQ7HhKG6lNlX+
KJDYdYusUE1mVtZCbcCGQToBHxE4OsxY22+zcRdsB8qgRIobviNkmJRw3BmxfCbS
fA0q6Jh3MmxnvwPXH9ZO8twZmb5WXJAsRcBjvGOHjkpkCCp1cY1lU59Fs/hkMALv
HxZPmJA9aBcSYAQq51NpLQyqKV+u7prVPvqOs/AWNX4Qf3bW1wgaAQtgFmAoYfi+
cLAI41DaE19GZdEqe8AHVbkpaSIAzE13JVpwEYzGvVVhieYrcy5T42LTzVlun7Ph
4zuPvBDo8+fy0SP77oQOTAPJWTwXZrHqjqrjhVGNnUb2gtoAqDGUT72UHBvmggWV
NOCi24TyMO62hjQ5m6oLyuHedA8/1alv7uabgq11B1R0XkqYj/PjdVCTAlYEisDP
`protect END_PROTECTED
