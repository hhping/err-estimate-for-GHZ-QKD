`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnjCVkTr0BeECVSJIEBPTydW1JLADcUZup8Y8K29DaPjuJKjxRrW3c/qMzQXHk1K
u0Gw1INZ/7QFRyNaBy7O6hvTgH9zWRnzjTj84Ee4gvgnJCEmqy8ABek1txGUP6Gh
Mk7Gs9TVt2LOYMSLc10sd0YqmcanyNB7sUOhNNs8gIXHHbXayMM0G6Tc/q/Mft2Z
5OlLsCnUr8OUUj3LpU8+8mv46prnQMQ3N6hSY4YYlByZWnYFQ+dfY1xe+8WW9CPB
EUrNBbg66roj16FanB5gr7qXJu/ZEGuFZH4whFRZQxmLGUO6RiTQvmsuCyIoP+9l
6l9G5SLjYuMwZ7Sn0LoNNqchb8bJTU1b1Uzkx/4idfjpKwZvpX9FAlZufu4F0L3Y
8Wf3AzsJiJgH2mnAV+qVJEeB9cuOtS8G0Gg47kQYzruQDpTpanAT1Pf/PgIyJgY3
zHYVylqRtZECLEYT7JPQTQ5peg/1+W22e44WP0N9HKdAgkFz8VB+tD5j9k/Co+Qm
NUJ6/9EIU8ZBw9h6K+Fmb1qRJ02EzByOJNtMUPhxpZX/ij2nro3hA81ALdivE0LF
5y2KtT2TDyRWvfgAViQfbtcpsMuaJ7VX1qKdLJXnF64KC9vCpY3Vdh+uMbQbI6Xt
jdj8EOn476y2o5J/TQC27g==
`protect END_PROTECTED
