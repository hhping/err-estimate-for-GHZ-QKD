`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qx5FX036W6J7e7VSfyMU6LJfT+AqaYPFl0r/XN22fj8kvnP6bkNQxwww38WqExJn
VEdHR5AKLn7qKrnnWikKhNkYmQXaAVkOIxIyLQcBtsZZ2UsmoddBjHK0Ol9X2Kbw
3TIKtGmbUcIWrjn9/bobxLGLBxFTdP26l2ljSSZHnaL+Ddjt5FIPnT+BMli4Er+L
R4r81xGkessQ3IStyB5/+ce2pBymYdNCxng4w8wVwKomIn3g4w2SOp3IL08fUOss
vIzYAIlYOsGoyX5AtGAkzWTqAlNlBujB4/OgfyjrNKzkLpMg8fELVtG/wUdPK4o4
2WMmmJ6zXEf/hFaDooDj7Ei8brHKkfbLqNlwvWETLof/1SUk7/U3li60oPUVi1Fu
HagluE/Miy9m/Am1H4WzW7EZF8pl55R3hVpJ4qz3CVP4ufa0BYxE12sIdZoxBRy4
w398UNx7SGFH/WJQQchyo+iOVRMzJ2oqba9B/NLIfDYlao9ssKmhavkRfZ+HDt4T
Vk9SQ2QsUlNgXiRGrmW3cFe+FAxdaAAH5s0Pd7WOyHvccRzw2RZlWxA4KiiHuWt6
FZVzKzApPrQMguYKQvt7uqhjFze/K7m8Hr5xBSIKyNm3R4vqF0kUwtswP3UPBibg
pOKdHMo+YqjCscMQh3ll7O0wXoJWrPtXJtwckWa8vTg5ccXizXfLYrz3Rz4TxPUs
oaMZuF0T85hCdM4SWPvAWw==
`protect END_PROTECTED
