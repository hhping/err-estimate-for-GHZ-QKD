`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWoDhx7dNrZ5JtBW6bz+ZlIbybawqYpisPGNilENVrs7i95OBgrsRtgGBdP+UON5
VZ1FkSZxzV2+2iVZZs60yw7L+DnMDFyA/MqvozXwMhyqICt/3Ssw3AFsNHiKBgim
34ewnA/QHAqEmCL/u7yjnSmWGep0mQxztVenJvLOYKm1mpEWyzzrQDbLVdl8BreY
uKmvz0pGyUdslMMAqHSyngaoPD36T3N2kZ13Ui+ruk/k7xL53vBGhTYXkZkVp04P
+i3Yv8WHOvQFiCOw0I4RdDwgivgycsX5A20/LMDPmYJ2x47GzwxKUpbajYCwGxkI
wzcNuwJk0fFSuTMe/OpPAGot35qaiDQ6W/U2/+5I1bqfW/s6+ghbOc6mbR31g53v
ElOAEGAWcrGJm1qkKJc/g48uJTgzdjeamS3Uaoo6aF0IXJZoJavqAM2awu5r/EV1
/QzDkV+yCKyF/jW6QyJVw5IkA4hE5odmUVPxT2dRpAkud2+u8DXHrd+Kow89X7Ab
ZhjzhLlJrVSb4jGgOJSFQqCW+aPCiTShOfvl3ZaWOWpvrRBCnoIf24fLoZbj1HHl
Pb8RCvtPQD9hIJ2EbSkTC+DJLlILS0r2rweUTs3y+s7Exvh5I1LkkD3rztU0AS/7
FvKJcY81z/J/6ysTtao6AJaD96I3Fx5QDFEBBGYgT0Ur3blaxhNg5dbyGwO2eBtV
JakSMv/mVUuXiOtmhHBxDl0ZSYoQbxaMGID8/tkGn0S6v+IyPQWIWYQJGn8WgAmo
MVUfg4uu7wQnMWAoxmYrjuxf5widmbRviM/Krwvjbfx62pKGw3tPfbRF9rwiffFm
VsUNisbQ+ek38qgrx8NsPFH3IxIaJYBvpHhTv1R7IuTTUVn8Cs3NBZw9GcVGfBwZ
btBASnnLo5vUPxtpZO3LhOaubqCKcYZTtD9QKU0cTQzj9VcvtzmMJJwjsZrsv25g
fTKUnSl11P0xQGgnHnZMBBaNqficP7TEGdNha0Qp5YHffh+npwCqTWtahtTGdRUw
EqFlqIoZv9dixTjegQp+ZswRUj6fyuu5jwhxhQ9/iiBa/OQRmDsjrt/sDPKpt+oZ
rbtY+eNhvOdx74YWKKzlt5JxzvAhuvU/ov+5teDYJD/tlar8iB7ELWdt1pLAvcW3
1G39IwHP8S7ZOSyklZcJwlejwdCMrvo+GYfYiudJhxfvIf+nKmvtrw6hyUh0aqoQ
XdPOyVb2eIFhglynMfSAfLK8M8No3yS6x7baTJg31exGJKLj8jUVVTT6gWafiXd0
7iQ/kaNg5BRF3btOdPh+uck0ET45E244+zX88iju85YyJVYCgv4cohR3+rUnRLLt
T1H2gZHR+1fWdEtPjHRQm6k5kcDj7fRWSR76K4PK/kY0l2rlAd20anb2sI9NLnPN
od8Dh7O5doW8GWMV/IBP/fLchM4dMsEBKZ+Vvjy5Lzt3PslsK5IzwfLhWNgz8Nwl
gB5wjm/AV752aCCydlZewaYfwcH38cv3jx65TiznHjjl/Y+g0eqM5m29LJAo9oFe
ruSmzODotC5pKW5kuTNOY2suEJpZrlhs1/YI+83nB6JQdkewFjLJMN2SCmBr54JE
wOFqj+47r2WoVqCwKuJBM1NC1xVzXA2nAlobNOWRD0StFSTtUC4yd6cVctwqsejC
1h6/8WBkFAeFhppnSaJ0goRSFI6INm7q2UQ+ABSCkX2h6NJrmd/7GetbMQM1jVxq
j6On1xR5hl/oJR2L3VGSaNHGzP1vXF/5UZeXkU+w1WPmJ2R1n6Al+hlvLLCfkKWm
vK/1X2QOOg9oUrNQgKG1015+W3nH9nxqJUeZYgY6MhNUsqbOtZtS/L0DfC/KoBqS
FZ4LZvPORsC7WEA7zhGSfg==
`protect END_PROTECTED
