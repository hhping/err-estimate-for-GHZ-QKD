`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L71k9khUVFlqJWA4iEvlDgKypA0ketRyodOZp+KvNVuLJ8smr7IOzoRo4lfg8HxE
ibaBfB7L3Cmr9ZyBYPJHbv5DQF+b9c3oifGPSZWvNpl4RepSBsGoz7azW0GlEkpT
W0TmaMhKAzhhzUqkS919Lvx5jRZuejIVnPhNHOZUuLARvjS7cgdfGrsD2JqtjymY
S40lqvcaDL7PLfZgDeOBp9+Zt0AOVfWZEyAFmuyzFjU7Kk3ELSUIEmEpYRXOfSDo
HCAHNSpo/S73kztTuFV7v++5XVrSWXyQd4vZKQs6HsQyL+RlCNTjEx0vM9epDUd0
KZyprCp0mQgOpZoAUl0ECxw1iwYZQV/FKOKPPmrlvMXo6cRWQpRNcQPmcj9GjTIk
oJtQvr0jqIqZLiLyDz+jbFvICB4nWv5sRaSnG5iPK0ygsW0TG1nAbQXaUYd0LHxv
XIPQHk3rAbA+cj098eE9AsYhcuJSQ9XKl8TflQUeK0kDZadt7n8NDfFco/4CAtMR
EXaX+kmayz14ju07Fy0sjVGVIUwETAdVU8o2KadXVqt6WE2VFB00HGinUKZHpAud
89gwYH2st4a7TsY4oSE/zhgKPDzlvLYlHYwL1FXfHIZNhb0OEZhfucSseZY21l7C
yVc3pNW9LurEGPKKRQuZSrYn05OwhX5hgpLWwRusbpIOectmA8Rme5AhRVNwLetn
ldzL7LkE/b1TfRQCQvpismpvmTdx6HqZHOp38oZTBse7g0N1wjXZuOGe+BEEPJXp
pdDJOQXdZCh510SD/gCnmHQbjfxAZ9FDVKrfH7brpOoNT1asaySTgxZBAW8nrArq
HWBVszyEsfkzbq1HUwkPJ9DDRHiUcl5kYuM6KLcYdIMj3bik/e0c8xdvJPIkFv43
NJYFUxjb5DmgG0WBCEgTOVUoZEtOZHhLIrs4QfjfL423N9NspmtXUmo/9iHQNRYY
QdmmYud5x5mbsWTZg/xqCEoPe064Hxhx4m/HpLXcOUXK61btnlbE9opmqNRM1nXS
TTzIsatFs5hvo4C0czu7JP1QwFpp2lXqEkbxcFUnXBqoorE2x3bIaS4LFQT2lvCE
0GHkeXttfM2Wms9ySzdINSHYdDCCkyqXUlyQMG7KjzAQxrWuY2w/Ldlgc3IwjVTL
FGhSKgR/cRL+q+cPiLiYzsjgZawRr8b/QP7jzNiyse2uf8DzrNJIXWJ70S1dcx4a
Tu4ZLfX8NGYvzWXbStTECyXgpCFEqWddjEAtuxT/bfoPzgLMfruEj9t3MbXRXD55
Dkqn131ZDkLln9vDeeN6iUAdwAnaNECwdVFigLDb0C0VkqLa/OO4o4QJaNNqmsb/
7D+9Ic3vai/QCOXCvXC+vTve6IHuGaWVDgtn8Ah5JVbtgSwRXDwKh9tkGQELhKcc
uA+yBQrquTmyPzrRzxoISffi9AYGBdGW1tiemlGDKExTemAIJ8F0Q8sdUCi8OaDF
MbEwY1NKXJaAjuo3qf510TY3LGCuA49edra4K9vAu4TJqeMlYyaL36laspaSl+1t
IT3VB5oXhovdkZMnq5UoA1KgJgJOajhgnsTq7GoJ+Gk6oKOwBuZ3j6bMEZtrImms
9KB+aAr8AN3wyLpN02cuUdW0t8axsU8zwG115BYMkX4F2++q7QMXJ52kIj036t13
IOGTeSoTHXpJVUEY0UqbUtbepYBCu0UWTL/6iBgzPLjhoSX4BEboMkXfo1x7noF7
PR6/Rx4475ceFIKlkRqqXSIg4ypJkewDVX3P83fhDw2lNXlTRaGPEChQDnneB6ZC
UVYW1Lmt2PoNA/rO/DdbQ70xJEjMJJ1a6X2tbk8/O1UFeuFTs6X2OCXig+l4E5N6
S+Lt9LqvS8fSOFRd6nLLeW2ahN+CKih/YYF59qBKa+m4rg2cBxkGWFMwfBCvsO9U
8EbSXRw73EzkU56+yq5Y3iem5T7+MRdYCtj07H4F4Sy2OHXPS3vZySP3bI4ZIe1C
meDLYu8S7Cy0dTRev3Egm+VAVqwnIhEtsNRQVKsm5EYjwbPq3gcd8AWJr8/nOZQl
x1ICFqPiltcK+Ya90sLBnr3fleFKwQaP4bk7u3/HLfpu+dfhcVm/1Fjy0M2zJ27Z
eu3oozOTVeotwE+5Lpwh4WHF2wSCpC7Qq7tMm9Zb/3momQADUR06O4iAjs70qipi
zZYg3klsQDPEnciB8zNS5g==
`protect END_PROTECTED
