`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yh9Dq4x6yz+m2B2H8Szfrup8I/Rp8nj+Ci75Y7DbcbYy69a1+ZiHaGq9PJMIQq0v
zq9rKB/U39IXql9DKJKeYgnz/ujR/rypXMikQhzxuoCd35B9knxSiERbcBbC9A7F
LvGSJLzjA0olA+P2NM/AzUX5IsPDgwDcQanoM3HUm1lS1r7QALxiLSjKUX2vLh5C
pnsTj1DM2p0x+u0CK0COYdZpo/FNMGhbatKKYxz54CqUpfHNwERQzMlTzMPHzcK3
pstz0Dzeka32pmWKCcf3vwrGEoybXGlQLi1NZDM5/Q+FMYNVJNTAx9jTNc0GD+/s
liiCZ6nkIA6tfcvTY03ETG6c5s1woTAnwafY0PSCpRqNYeLxjc8UZzs2Ukddajni
IsmKrK5t5JpOtmQ8QKhbXbkXeqC48glqeSbF7Fj2zrub1D63b3u4SwKSBMePpfCn
72DjRcEJzana4CrqR0FdfJSkZ/rDWf30HQnk6rGSfmlJOz2GYMwyhHoNWD3nRyqE
QdSwfyfkXbjqsw36aB3i62/fDX8r11sJWUIuBrEv1fSYvvNDXVAfAy0qzNgUIDtJ
Ru3OMqDoiBZUBFU/Nd4patQwV4IDpSi3y0GpO0Vd0I81eV1FFeK+2gyV2H3+q3uS
f5GjUjIYkPuM7vESAJl2mDopKaXkoCItqtIktrPeshwTLpI7r2pWoN1uGbIZXCmW
aS0RfiQwIYfJTmgZYY6r71Sw+M9aaLSz3Ecl+zO1fN3ztRVYSCJlLb/QGXkDN4uv
bscZnbOMOShWDLpu2Eg/h8AJr/THXnEpkIGqH4rhnm8Y9xp9+uZbH4J22qz8G/b5
6i49VGbudvjzsBoV6ZwhWz6g1i2+D8hGMVwTlgM2k5BrSTK3Ezv/xzaU4phJ0fEM
/a1/pC6zfUkxQ/kFFQSeA0p0x7hN5J7NcwVnGcONl8Y=
`protect END_PROTECTED
