`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhYfI7Yi6gKJv0B4rUw/sHNJ63Z2HezYikvK8MuPgFoPAwpz2RflnCUqSAAudZ54
3gJa9ZaONreHmtwbHT6IQLbeSKO5/K8KfkaqY23QcBm9i2qt/BxObZNQReQcMtib
dqqjN0Tjr7ZMlLP0bi0Ij2m39PC2sV47zUedaNVqcGXuGudp1RniBp/5lCiE57E6
6/27SHzMiL3RhVGdS2Cunf8////HqyoYynXWNpQk1OeEvzCsbtXlaEEyYSaixdZd
cjDdX8zHfvrntRBy9uBcnch4sUTL9Et1aL9NnQP8b0oVH0V+ysYgZM4cKDlZtmdR
HLkRXnNwymgVmxa/WS+taviksIWaLdsJFKj+igANqAZmq17gE6eSvWX3Tms3kLrF
V2K+udiz8W49HGeyoSbTaI1Y/D/6ppA7aaykidS+CsPRINW6w+QiyTwPNJWPVAbJ
FYknG6JVcYez8S1n2L6TZ0G9acmPSpYixVxtxLn4FdTfGXo87nz9shrAZjJDbPlP
t4oNIsPxWkWgue8aL2hESAyYTlSpMdYMDQaVMazB5TQYFI8hnNuLABypzAbRc+Qx
9AyGqsSfajEPwPTusMD9RT1ImvmpFZLmE0fnVoheAjQvJkPSivfg35Qb0FMlNwpk
XsmLjraHxfJZrM6HTbdo7dkK/JeYlTItPx2XCihm/tZ3J6+V15AGsLTnZZ3B2opt
G+ZLy5olj+3ymaEMNGJB6ERrE9a5M+hT3ncnQEvT8ph1dAsuZ9OOUMgTWeHwpaHy
2NqE1ZIhSq62kKft1bbibzQIj1PrHmzcqoy6IoR5g9d72thifyMe4LNw2lP6Ggtv
w1bt4n4Kgn40U0x8HJj0a1V3U9jW8YczP+ZkyU57Tj4H7BLj5hQYEbeYRQE0lDOS
wnDv6dGrzewZ621e8T+Nd4r6uMzsGvtdDlo1BnHBjhADuYXe1th3GCRiSGLXOpjK
tP7Wrs/Ln8Ef5MaR7LbMTEoJ0NqIPU9y2QC+mM6f74j/HEQRMXOMs8Oi6eqKYb7S
nnUJfu4WJext5DtmgT0TZJklFA8q/hY0INjISLTASguW3OJ1UzVaKgfS4CkGcqK3
uoCYX6SAaUvRbspNV6wtj0VqW76SQh1MHSr7TIOqUHLKGe8SLzvHlt38hMricfNB
6XlRZmpqGPJ/oKMZOjo/Xo9VfVuA0lEKRir805z0eJJATk0wH0YUSbi0gSu0ZYNk
iIi2WyoFNLDF62DLR2rtFaaUcWoZNIRCQip490zJj/cOjrnGiw5ItfcpU+v6dPje
l+k13ckQpBn1uR8wyxt6NhgwXs2WSfWbQFr6EF+mu9jSZVBvTY3AUsNOAELeY0nk
6NEHfw3EHqBIzg9iBzglGk6/Grc4TPQmaA8vqPRsrcnpORPgpCh6sjqim1jKNvH3
HRZZIh9NghcdGS+cvf1CcLoleUeeLZ2DFYjjAH0GFnHl8PIJKkM8NYmW1jVsSJW3
dgNf233hShhdyBoCr+D2ZV0m3lCZpjj1IqyEld824IIEOetTkRTPXsh1HSf9OgRD
UiGIMTO7zSEI2R3bQvVDNNYsg8z/dubcrtVjtHe3qxSfdMaOjp9LxYpSbc7gZBHj
13zmd0Df8ZtzcOhCqIBYOFbFxPbc39vN1zZ14cC2jqPKlV8uo4jDtiSEGHpeL9yy
ysv6a1kN4x7Ljm9CXOxGR2yMwdKljbNwUVodFm5YTnGUZ1nLX1bWsIzOcCkJj/hN
Bb0A3OWfgO2oHRvEvTmvsIisixGrgVFI/vmEG5QBuT+KUOylLV+uIEnF1VVDhZqg
0Emj1iv5wUfItOhi5KyaeId6WjCEkSqdDxIGgOJi734i13cV4GOmCSmk3h0lVYow
qYb7itX5J6n4CBRgITub39kq5miSuq5fiKzjEUUveclHOe5aORvRvoHvKeIyKowd
PszgUwptWhwBzL9bF3Wap0xqBq2j4GhtU8ukdmhJL4jRW9vCHgR9PvCFrQ93ADW3
VFYKKrgxTWrRp0K4+YMvW0upn1hmC7g5GC4ZOl7DQqL+TgsVgEXK6gQWJcSdTdSe
Ch+WSa0TWmDG097le8aSWCvzweFSMO7b/LnVwcwt+9q7LZpmufSHNQLfiOinr88j
BkE1GAk+JaOVdqJ/DEgxoqphHycl+6T3wFD/r5IzDYSUulMNiP8dVxaVKcqQzSJ+
3Og53xqrsfQ/0MwWWVpjJVLRlsDnTmnPwIszr0kqLHeLjdgaoK0OsUiMYxqWheTU
XpOpwcpg8sowASNH8jQz3AWxc8D3hIlxEdRrNSk93oIjNqw2vpQAca4eCDDRDdzx
4NyPFVJrIrkaQ85YltFq75UnMd0Dj1MvseY/0Rfl1T/KAKy1wVK9yaUTmoc04+YY
nnUzYXZRNki+c3aZsopux6xj2bUpsPfJNANItWBR43jSeFggvcT7oyKt/2y6p8OS
cEPDCBNAjaaMBzhawB7LlYCUuajo9/U6Y2T2UKLaeaHI8F1SW6v85R3lEYssKRfb
hDFrrZQ3tdKgCylH2YMU1/Uqj2WkmDZvDCFg4km3noepkB40OLOf3vEDTPxr4Fwv
bVBkat2BO/WF34d6ny2eGBuLdDgec6kbBLyI+8y9i0L0zzPEBbtLp7bMi/jiFy1r
U0RYcWEum9T1Z3gr7kHoiH3o7yPbY+9SvieCVEkG5Toqm8/JuZ2Bxit/fXd6dIvj
S1Ub8K6+Hgi9W7hzBVQzcIGPEyGEA+/oVhxwmyj1PRm2RSsPqXGmiAjGshoIpUBz
rV3RVU9pRpESzaS4Mzs9bM5GwHA20yH+QTxEq9lUN7OAL+ySCzboSCcQe7guB+uF
WTC6wgdZThxkgDhSa2qjg8cpMmJpvDZCReuHtm+2ZxUpmDfjQqY5aTZ4ZiNZmIrT
X02hJI4RwpO2wlnlWmRzEpbcewuolq3iPGCFgWeuUuv476TZsv/bQ3scUupQRVtb
KmOKv9+9N9qygzn4MZwwZowVIwWM2k8At91QWU/SHL8McFn3uHY/RJ8EekcZsfRQ
WxQqZp+QQ4szV+hfX71sMUcC9cZXYwKMItXdhoZlNwQIBIUrs8YLcIM1BHOngrAT
ia7YNaNaSbSe/2EneRMoEo721vKc1G85NvYUtIWyp/NU8EswSj/zvM3nDkU6rCDf
NUsCU7r3Lbjj4O4R7NOr8Plqf/Kg6+BZirw7/dCWoMHECfpKbiv/CZKuzz1DH5Eq
WJk/cDIOzUsk9fHpAXbFhH75d4wvsY0zTWJqbcDh34xA66Pz1N9CfEmj6zrYpc65
aACLNNpRrclic16XGSWWB0dEJY/gvkP8i7lqBa/j1hucUhS8FhcExpYhiWaaoUVV
TilNFHTiR9nXihp+U1pJqHF4QUSvzbQMLPclJRVUjBhMG37OTtUyebp0xn0IEqT/
1tpOWbG+vcerJkYXUrHrKUCbRME+mw1zculJbjOlszjrY+ycA2eQWKGVMpGQYmbN
BtTZI3ePeo4UIs2jYK31HFaMURNmjCzhaeOyW52UyDzpKnV0QfAgPwRAQ1RS+2+h
b03YuCit9Yt4Wsi4gMJcRQ34LKPv5qj5n9gim2+iJ/EH2mkecctdl1Dlu2sET8In
ev9EgkXO5UfMi91l4Nvr1/x41exTokOqpEQcjP+vfSCUi2WT0czMYWP0/Isx9Scx
y04+BO6xQitllEj7OMeiFfboRSlbU+W1J/4eZa3xrd2N2T8ZCzM6Njz0U9HOHTx/
qrE52QeThQRvdveCHZki9fuYHTI51AtoSkmnS01ETKRFRJUQSYpmIUIFDrFdhwmm
u/p9Wrslkf+z3Wtq4LEDLSBzdVdDWhJircnFe9qqqNRCb1PULhZ9MDXIvstjK+vp
hUoNct7sI92cqz2BxX1cXQlUmGpTFozpvxHK/fZCiEOZPWStq+fuoThxKDTUSRsM
X2mSStJe2lc4//P5gGIpdiGOIoYoDnhcKRWjzoOAW3P3DJHOxzmTMpCaLNCUUSc/
McxT4kRTB1MFKNswjB0vNxSwDnVVOYmlYuSmIn86PCyBib9vX2tfVaQKLudjbDdX
gSIBndxVprfRt88Vki7NBvRUcrneCNW7bmH17a0Uh10=
`protect END_PROTECTED
