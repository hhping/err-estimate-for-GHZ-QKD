`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIiFw9f8IgA0UeVugn2JOsecDtT7Y76ititdx7wWu6AETeiNuLTo4e3wrTHAWeDt
bGpwGyHqg1Xfh7okX3orWTJbC1TqkBHExit3XRTwCu+q3eWWEQVDRPMbc49iOHBB
UhUPaW6KWaBrFsYGKiLTCx+Qv7Jwjtum/7dChwNuwmk2M7ShanVlCjm0FDaUTK0/
Ie+OYXocuA6S+G0J3hxGzT6oZ8PvEr7kVqRKZvpeiHIxavBd4v0YiFgITgi0+19W
xlpOAtsUltchZr12c16XtNHfhEPy6em/r3Ns3aIP+SqS5PGdnAhBxpur3O2jII1u
7K+UXWHW9Qyb3ntLV8b2FVoEGVeQW9DtkrtRUThi7OmUX5YzxG7/gjtn7JILDt0H
+ohyHifoP6aSbb/+Gq2bI4zzDOiFU9gKSP/AWK21jaxHDYRcADzfnaXoZ9U+Rhnu
`protect END_PROTECTED
