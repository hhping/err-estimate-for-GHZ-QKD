`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybKfyHHtjiBVZ8yODJkwoed0NFhYShX6tv/wjmLUOzg+L8AUxW7nnMCLXaL+KMkB
EySfKtnaYrlj86hTMra9yfLsrpqsvny+7OuXArlAe88TK37qR3JBhjjsWoH2qyK4
9CYQjK+HwEepNrQ9X+igoLN9Nv+UivkbEvdjsMGYszaaaZotcR+DYCxwYpymIDri
2aJDIcbovCg12JsTmhobC5tHsD7l2eK0YFe1f0q0pl5rk6YTpVBbL4OY9D+1ZMt/
1gAYb4EwNwNOQbEaezzDzzCEo7Rtu1MIN6Tj9cqo9bxR0mO8lhhjeX+UbA8p7YU8
/K4McMXQzpw1HwxaucKaHjXsaFI0gwyLXiEeaM8pjTPxy/1heFMInGVbA90AfDU/
pSOFJjbXG2CYofTYvLIpdi5EJbYz4cx7KX79TLOm8n58AmNm+nbnXdHHiz0PY8Ss
yWd+eFgZ13URWweXIeqyHmgyYjgl5hT73KG94MhfU/JFJducZivP3+/YSdncBZ1i
qwo696UQQE0Eyiwvo2mjgRrp3am7sOkJq0krd7gRiET73YjpieYmBHpcrwglOfM5
geAO4D3EpFfxFqw5y0sc+cWNf2vmM3QCj2D1SJ97QGtP66uj8tjNYfwj0tSPmEfG
ZxMR/DYENTCgZWtdQKfel08MCDA8s1fdOe/AVwQCDU0j+q6Pb/XUqm8hWOfuw1/h
zWh+X1XPBaiSpZP03JFVpWp+F/AF/BXXcj9EEqY6w7RXx61fQbp9PUheQJz1nK3X
aN7KvveD+/cBdEc2fZdz7M1EDjARA4rVSpjRqacJXhVc/QSszulmSIrGXHIs/0Ih
1QiCURUkicEPH2dEd/50kxviUyDswMfLqRlguQMLzNUytp8T/Ziwu8s1J333Au5+
48buHOUwKFNf0uIDkngG3S096FuLkic7LIPJ7yg7qYuQBAMAfrGsU55rQhNDVBFw
DPh8MpJ2e8B9AdQkaNBXtCvYAvdK9TwqVYW6KQwdg1yLkPmKklbY6WN/B2BC+uoF
y1BOqMcsrJCFARMd8HR7os1zhScnbYpMXC5HgGSrQvzn40g+QC2T3b/y9cGKPRcQ
WG7f4NER1DZOWCiaDCxFsnuWLoJ+98wVPIPwPoQmqnQvmyvPs7gAQrC6H/eg2JJ2
ifQtwsdAqCbBIBp9O0m84+eGM+caByr2DbK9r1+EroCPi/0QtRHLdqo782kpmEzS
EsioPly3qQ7vp2FKgy0vot/Tc46f/1hF6Z1olHSpgIZnyX1J+Bs01XOW8PlX0OVW
p+sdpBl6etUTMuMVtvIoN+I0FjW3qPlT5Xg2qpt6xQ4hkO04hI8qUmCDhpaxQlJG
EzM1mNW7k/4Xq5SRjYBGewhTmqG1TSo9lAAGn+4pu72B+/kJz2R+SJGQMM9+jwbh
4AYf7FL6GZ3Mn4SOF3S01mA7rcn0QA4+F505kxOCLZRsdF4eDIZEGtuwRIQiC/40
hlLsNL3N/n+KmduK9EW0M+TuWgnFHvTnO1t9qMvKYhppDafcf0SLxH2yt+9+kLNI
GeGFej4CTtp1UbQr0WcVcfegzpssGSohDj/P6jmxo4BxY9pbjeXbPV7bZM3XJduO
vMp5T+W83xXydG8BMD7iUfxElM3Yf95RHYfDO1hX8zn9ASYKhVncdiqkwFUgI5zf
OrYPXdIiL8+rMAznihfRTYC9p0vxafTWoZbQbzpnN/fgPfVBlKpDTubmbnPHXEXB
h5ks1VW4X4KjjAKhLNs74SCasDMFP9C7J/3sTkRE0Xebdma5ucLLnVd7+1Cr7mh/
Q0GnpNeSGUeD8ALmCaXosCKZ5V2n9OIbqd6iDAJqM7kHTfGYKw7yLM3VqRbl9uqE
NL4kFQDFOMKGBQDqheJrB5FYpQJq2mlarN2ZubdqPtkvsk4sTxOfx0IfOfFq6bHB
LMM0WYWgF1XBzr8z9U1IqpWvs2K5jpDRFKOPuzegL4s3GffUoY+vPUS4ablLZ9R4
DPAUg0KDgOyTTVeC1KvJYgtGczdUuUC7tL77+tR3iBxrv0JzFLAOk/0VKuzYwi9K
MbLJOfIy7NTdoWJ3j30pbi7tekQKBL9sH5yCw1hc9v5hQ637bCFbAeCOnDCyqvuW
ICtD66l5lNaQshkjoHX2jsu0DiIcZ0JtYiM7HusjHOq8cSXe/sgnV/VwFiqYSwnS
bHZ6+GHAqj73ne9B2+10ik1XCW8dKmBXXLcOua1cs3l8xmYIcjsW4SKAkCCTPGml
4cZ644wDH6WV0jQbOj7uj9YHpA/pevtC+ENBATIT+P9G7cIhSaIsoq/6vtGHlGLb
lFh4LzTe0hXEfXiC2EmRZVBo1jhPQFpbxwZVRJUGlTbJJzrDJ0r0+ZzqxXfka16G
Z2S35ZIxbOYAO1TaDrJc9UfhBwnz4rypTUbSLMLsFrVJrAckg4Nkaxnlt85pwmmt
MVuHrCH175j9B5M8CShL//J7V0jYfO4O5vrddL9I2M7zXaz/o/7IS8xu2OgREHTG
BKdPrlyvDfDOIOhJNdwnAJppzasyKEpJp3bs6yU8vmXOFs3cf7hINnE8D0oGFQLS
kYu2xemgrAid8EEDFvDB+tsqnDvp6066m+UKPpoDhnUPoe41EqTNepOwxq96rYxo
UYqrnzBrRE0XrvwpL3NeeH6KvSYMLx+Qmg1FBRWMiAaGhf9nk/wdHhVZU31gEpKK
Y1IQCLUFe7gE/uqJI6xaoEpTInLbF4TFwz2ndMX7kP4rHb2tCIiIvdyTYJZsLMif
oukMyZ5pr8iRFvmqXvnx5uE7nBf49wTelJ+BdPD2uOpmkS/aaN3Dg9jpeYUAu8ws
Lsr6LPhz0UrreVJppcN/lCzz56ho2omJYti2OiunOEN/o04w/XgOESH2v/si+0U+
sL9HBEJ7LvgZJBi6xKL1FwCB28yIup6Q/ZUboJbEu+Sbu7zIL1ws6pmylNjiV3Lk
6C9uSHfrN+AfKLbmcx7NO9u9pWsU5OUNeEr9axwN9wuIRoWoV0goIcIIe5OdVx5F
T7il6EXoF8XDzSCxSDydJzheh79ErCyp7xzh2bItNgJbFEKyPLK2ZCUFCAsSE+1O
7MoDt9u/D7S/fyVo23h7KZmrlsSkr1azunMAxoyo0+d3JfeipgHC/Vvvl5tU/M+f
lE/5jg6ixXa1lYLRYHj9BmXuOwVPQjxW6+FS0HeessZ3pzEalZ4w0YWSDopMb9rO
H/Ky4kzBnswwCcZD1cazXzmADOPvh22zYVMELYLC+QIk4xItyGGYXdEvxkESAqFA
kSJhIRZ87iHrnNpx/GuGK2YtU/LV/8XkupfG3V0PCGgmWPjotbKkYvEfMTeZ2z9K
JcEvGMbluU8rjfYmcu6/Lnzqo0FxDbVdLTTuOjahNxXJBJb37Ilp3gBmhVlN+wv8
AkwHgvoMYe0edBu/JizIBqDvezGUW3gGNAUX4lFytr7ftaMe68PLLJ3uV4L/5hRG
5zv+LBfLdHSNBeAC1XVkeuCmbxpn1WxVVhFL7IneVitdhjDxVCn5gTvLxm2bNKaK
eNvsT3huyNi/DHDm2hpL7m6QWJMUrmDwuvtHD1lO/Qxh7j1KvxfIhrWsEwSkg424
P0P/RYQ5oQTFbngyZpwIhXnKw/De7v7xln5E1on1Zco1Css3r8Q4Ho/FH/zzc48v
uwu1yETcL0diC0Hg4HJ9hLgwhNObpx5SXCGwR7OAuMV8h7I1sAGm2EXWsKwgPJ/p
RZIxPhv9baMzhY2K1ruXP+4ys5vPWZcQT75YHFgNCoC+NP25SUeKUBRIk1RMPKJt
F1bUKh3YMPIjX2ir/4zk+RSdLOgj75hBwKW6bJpMRbILnRaN0ONsoQCYNdrfgNWq
K4sf1LsXwW1Z88ybuRlUNDpE3n/Cfd7GPKpyaK6P1i3uPoRuyL9vhdRS754NGjC+
ZSFMkKTTT6Ye93nsFO71RvYJVeVQGqot494UQzBVskViM+8XZNUUy7v+hp9Kcknd
n8qvMkE9Hc2e1pWGQssNs+tZhj9fLPybm5iaNZ/hKKYZph5sIOorb5T/hJvc5ipF
hNujGy4JQsosThAcVQe2QyXreE6IVmJHTZ4XqqOTW5mQ3NJ1HJPGLLAHVHV1eMaG
SEJBguS0+cwOkvOO4crHrbZYYeEuoU78w0SFHXq/+2k+xtfB8+NQ5KqN00mHEujq
Vjw5Pv7efj8ZE/q13NRy5Qb3Zy4yYJL119g78vp8L0w2YUKHshZIsMidbbJizlFU
MkNV1980ameZ6aVudo4WO/a4441Z1+r6jxnNnv04zNcbYDnoj6UNTbW+fnA+rwCc
sWkEW57NuPOZgGWSeuPvoNXtTrzeWQvw0pAL+2dKsy7VIl6cemAYiwllUVNMFBlD
PjUUeaXqL8YmYwiIwQpDFV7iQf2paxZgi7lGKvrmu5VPRH4ZxsLUaENpuovjQ2nn
MCcFOY/38GpGR3HAj95gSGkeM8pYRBwKuuRcx9ZhotXbaXJGHXpOFyKEMpLdVv6F
f9cWyMA6cy2SHubWBz6PwA==
`protect END_PROTECTED
