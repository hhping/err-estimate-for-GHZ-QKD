`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9wdcKt1QQlvK0uu1m9dpOa1F2iKXgKu1DTNfS+fdph1mt30CeP5YoQallid7m8M
L+rmowv6vhFlUsURHswknJWDmv7e9lig5fLUPF/TRKNYTd5HFdqKydUPzn24ChK4
KY3GJaITQALMgMcRnuJlA5TbC4u6fac/u1wZWg+fCQm4baPHDx6Eo6e9woG+X5Wo
f67GoIqNhaEHDDnwHueLFZU2y9Sqq2VHZ+LLsvFgsAKlHNc43d5HdvazhaJOO8hq
dUgDgri62K5RE1k+fq0nM/nfBtWJolOB4xpdn14J14XATB6PV/A6N5/2Ek0AZMom
C/Jt2DTPBXSLDXz1jLlc9nsXjpoeKmmgRO6+8BYpI+wdmJ2Uy+yjYljPcNAu14hf
z0GD+xQaXf26HTu5pXDfaUuwVAyhn3dKJKQhNm4mlhnY1+WoNTHNJv61wLdiMGMM
ONgH3yZeNK0jHgOgf6vO6bMIg9GyvBhdlXs04D4IFvU+7FqGU20DefzDSoijH8fl
f05FsArCjFT3lyJIiE+jdoB67gsVSV9/KSLfxaLUjpnfnC0A0wnN+79ruBY0cIb+
sUZ9c4GX0LXLskDgzZ3mSNISR85YMtqdceAgnMqc/x8BY26xnaAPE2tpVeexRjJg
bwRM+QUh4fJVeoiVNEEbGhcN9vaAOV0YFwJ0w3PIiT8sK45sd0BnZiaVzzV4+Ixt
Vo9fQI6EMvhL6iYfGA6mUigE0QsUVld2qG5uU0wLKlHL7XfImF4lb++q0ukEDysL
Mm9SB5MQc2ohb7UJ01REsJZ8RgCVImLYqB4BbCajDoOAB/LrYEVpBzZxWxhdldM/
E7RVIbCEAnE3NHLna0+JiHwCZr55asl7evmQ8VfisSY4vTTwte0XnOYq5P1/xTKg
kxwPLxfUS0NYgQ4QoeaXMHjXM3ZSmjDezXDyQAuCUg3deVsa6+x0tTokkiirVLkO
bcd2N5mHKXCbpLb1q5Yuz20XWi1cFY4MkD+b9FTuBHCjSJ951jpwqvq1Jqo/xBNp
R63xOYpmMD7iop5NOp8eSTHbIYLDkZtas6V2BEnCnJQtIp8lAc8swxYoJdFHY5M1
+/nPSPorX1HzOdGoMQaekcOS3dNi2rwmZYyGg5e66VAIEOXtSwDxpqysW1IBClVA
Z7bVqwUHeAwKVlUA4JZQr+R2wSP1o07peCrJywMgbW1nSvol1wJIElRYwMoDxcez
Ots1PL6nyNJymYKpQ7pvCV2cvwknhxBV2Hop7g/emeqDDH8aoqwdvcszXXa0N8m3
Hd3G87woSzpBc5pb4Nock1tnNwSkixRwQfTUvqvI5I1+mLU4WT/DxzBTpF/gZ108
E1Z2BD8rvMGh8y8q2vO0QcWK8Sbdatz9KJ7ppzJQuRCYv3oXYkjWpR7KJM3hqCQF
pTzlX7ivNEjNLH5mFtb/Z4YASYlm9MoJ0j5OXuX7EMugrC5aKpxXNGJZCS+o/9Vh
/uaBe68qB6SDQAlHJEQeNPofTreJh7k/LUHxdU+NDCvpc2A7nndEY3bZ11cm9CJE
PpxizZfS4qlWFtLeEWXYKskj2oDZ9hmjW6ri3N6MMDC70zcUocwEIKHef+YFH7mu
GDMyM8tFya9OZhWkrFIKb+n8JNSXidKyR9oXsMrgPHe5NM+IMjmiTck4Bx1xe4bQ
90BflKUK6wksSCwINVD9rCt8geLVhPGcnfLeEVSGEOEfQ1tFs5xVmB5Rd5lqT7Gi
lNrTq69JmMFlydQvscY1VXFgA7XiQzLs7HUgXwsnY4qd/6MkLVwpFNRmz5rJ8st+
jgDdK76fM2EJrwsX1H0v6OzkkSUcWLlP6LxzNJM8l2isplY94qDQew8wC++TEiDT
HP51lqj2iwuXI2CMUhqRgOr2U8e36BoQd5z4wzfUV2SDoYU5lUTP4zZdMFCSS8oc
1k5ScOhA/fIElN+D/ysBzoMRWDxMxbMUrL7PyZNn7fYNC463/fWbXigfA55lj1zb
2a3DI2LL7VvdXuybBjfVqrigpfj+jYjPeiGGHOk9UJPC68/Fo93MxT0vEwiWt0Yp
6d7u2EQVsFxCVwLWsNv+kT7ZgqBAOtLMB82xsf1KJim55jzD4x7YC69GlGZ6Esud
tX0rPe2ogsiekr8lA/upW8K59ubsausxUP6Beku63hADZ82Mpo6RWz25XpcaXW9A
fVEPu+l3zDNw3ojSU6KxNi4gghFlFV/w6gaWlCdXMmZbzzHdCP/XuiJPVDsQtTdA
r37pCnGu4LYNR5rrJ3qoZWVvgfQep43uYmIx8GDn56F0iyWVLSkJW4JYjIgdp+GF
/lySATvuNc0KDYRVrY0c6JEanu0RxLHkzP0upBYgmk845Yjt3SpMMLj7JZBJqJ7r
68hos/PSEvPMzrLHm8p8RxIfzBcxLWyCaI7qeT/M+A6R6vFNWrd2Tz+g1fdESUWw
MbJ0RIu4jHcaCKIZOPJWn5KIOsDM6N09+sh6+h2Uz2QSipn1QBat9jpG2l5VmnaA
BoCzDrDWtXS/yiB75el/Aaf2fO2OwTADzi6W2cgP0Mn0DFZHvbkeQxRDeminTC5r
9pwEiKMIubW9iya8cX1pyC2ImKZJyTwaI3XjUAPIEqhc50MdIUZF3dAd2y6HXma3
fV17YyXkwL0qSbP/kTy4mSykkbu43TzbG3vJusW5DvZjR9iMRbyGgoRzUzeeq1VV
2Yyx6HBHT3DQ6epApm+hLdCbl+mtJixrhNQX/uOeOkzUuIyxrWWnD5LRb32WHiz7
mXN08ahlShzMydC1hv0DPoiVX/HyEWl2uk7AYmaorCV8VeYLZd6u1JZWIUtdSRM0
E0yLQuOy9WoqpktGFYbtSOLmCU27DjCImfPS5LNmGMNhkeoeg/WNjELhRU1sSGU3
B6Ku/9gk5UyJNBC1ppsXA0OdI++SK2RJDAQ/q1J4n3RV/3gRdKowSesui5krgbwC
h8zjwf/oxp3uniSsEBply/mDV3WTYQFuOzt48g+wJy9m53jkZSl7oN9S+UwuuIvV
4oK2upVZl9I4g/DAURYGC5K21ZU8t484ngPQy6f3LSSlmda4gQZBt9C7mIcRhTWa
l2EfTYYxiV5b1K/tGYu/zUO+nJmK7fTXoyo+SsqlMkQEKrX2p1978zAc9jRKL6QV
cHHWqeViYbemZepip7FOowoM0BI8aCWbxUrAloYVNsrIuOUvU/dU1YEOKX4khKFY
M8fQgDsBpbXMYBKYzaT2YecKzTooG0MUp6XFFSrYZPsWLH8ctGXMr3Wo5eGbjfPy
HFq8CxPbS8RRn8AZfSifVR6Ao+vhfVn09zVU04PSTc0A3/cTUechkRwTeq0l7gAD
KYG64RqXnQhAIPYnOJ44Yo/oy7Bs8hZxsO6cDQKchGiLhyuOIofCzaey1WFgYL2v
tlA4izV2DZjUxTzcKvbJEvgUUkyRtYCRGwZ2jPbXobT+Z6aOfZ2RrGI7Zufc7P5A
D+P9xrM5r34v0jpuVlyd7JREJZkPWQOlAvmTGtDkjCFQPiLt9riTnwDzRVitWe+U
rqLeqmvugaP+7GKVzBlfj/FqRZBdir2ryxxSSJU/YniFgetjAslDT1+h7b8aW4DO
XCCmd+8eX7aiWNurHnw+zqNYeq7Cx2PLNLhRGZZ45Hps00hHO8apvT23XY7xWtbs
Rf+Z97N1WzTmyyR8c60Q8Ivj5JFhV1r0SSYX/+pwtz4Nirnpxk7LUqMup1dyRuUy
nymcJDv24yh150XhbPrb1BLX6C9ccPRKGsYcnYHJvL9buaaGcleU2w8+FWi27IxH
rLN4RK7iqI4J+N/041VAfSGkJ9PdtP0am2HHwAYgj/HzgksK1UfYTPAMtHgixdl3
CkHxpg9Mz1S6XeS+JVrJMnl/KnUEkK6K9pe6Mhvq0bU6MJi6iaTfBLERpgjb60m/
S+vNnvJVOZb1iVSe6pBkqUqZAwBY3tYqEhcjpTONuNlXqukcR6s74f2vO4KvdzVP
3yRbIzZIj/+x8VTpfZupVM4nxt9X4T+o41dTdM4Xzz1LrrUAcp7TLEoB7ujMsdvc
FA1RmXopMcF8PtgdHphvMFSlHfsULvrtcRjW4vg5D5b0a5VP6z0QaBkg33VhIUdD
yGivathXOG5+zpQfDbX4Xb3N0qXL9K0/6qrzhHpJ1p4xelccjbdIJo5AAQ1odUKU
awb7LK6hC14xp5yD4jxRVjze40LepR53j/KYuiPNn2qbEyqAnXVvScSEZDDYRZfs
KWYZzUyiwlA1kIItzpCmFJt3ARivZTVAWAy76/Qs+YM0uWkT66x8asw+It5C3Xa0
mSu75xNyZE45CfkpGlGwqZBjXDRdR0XjV30ene3kLmCzfmkxOj/sk9RkcNrJMXtj
iU35OxBjKN3Evl1eeHi8ZuJK06EvaafN4aYAhXkZVNOp8Ltlc1qDUwjwsTHpbm7v
GT2bcMTggczQt8UJp3cbgPIDp6A+HpqF1+KAI/xdIsjioRyMGXi3aIH9112hsezq
6cijWKzS4rf2hqt6hOby4lE7ql8346/JqXw/cVk26d7PzmlBibGa7Mha/+YBTbI5
3IObNJVN1khYFN6IoCHei0GmMzqghuQWMAIkcDBp+BDKK7ytegCOwbJAUoPY16Dw
Mzou4VplK2a5y+oFOvcpc5N2KYRESz4fiTbfdRc3P+lqycuIQLXCgiJESTQp/r4I
CBtM684AsH4a/K/F/t424CySBLiSEWNqqKVcthTU1NDZZ6kYO5RgzuAJRsGiLnO0
83hIAtl96fTinG0mRXTgHKpwzZARwV1awqyFK+rc8h4zXbUFPj5qX/FTG+mz2+LD
FeaxBxmfIjeFcazo5yVmsyWeHN3uzN/PZcMfhI9pk2g5wC7epdiuNszdelQhazki
xkiqnubyj/KIyP4z2AxN9I5vSC3zvucdmo5dmTFq5HhA7VRK+5Eyjs++RWjXbpdP
iuXXn4eMAnFiMaku85ef61XGks+iaVEb9f9sxKmKr04lavea2JAKMp6b4B/LahzB
6ac3Jd1Z6HSB9vBuKdIlkiZ/9F/QQg+w6+q8TjfSc5G7W/tm6LEutYCwZqYisryx
DCv/xKdPduR2DSuzPfuWoXQL5JUOCkwC7NSpGbrSdmcELm6Rs20IlqmAyWUZ56bG
noj+/ODtpKGolAmjzHbWFJU15yd+hSaeESw1vB+HJi4eaXlu6KNUx5i+Tb81VCFv
9H/3XrX6kcdqMg/4mRX7QNsIBGLMFApKkuGKQ5clvbDaBbJzbyI/HgbCiw1dkZxf
0EB1e6iIIEfw+Br8i6uiJluImCGs01IKhqbT4ULivQRYfNCVm+2gDrRGAADJRKxc
XbU/P0Jv326tt4ehxVI7QEDbieN/Ukf/k/gGEqz5f6CnljQ01noQeUARjeKnXqqD
v/I+qGIBiwauTjTjAucg6T8X+UbZCzx2Gc/cyoIAtJ82n0W+PfjICo1jbsNfSfN/
I4fWjxyV+7S16/ULfRm+Pn+i+Yapep/e6C+HsGvZJpKw4h35Ej8BbtikgZjQe8AH
2eiPPPOhNj+Ux8ey/jjsEvcpWeNTEIUOxyxHuY7Y9W6sFVrx/grvToimI8ddf/6L
UD14HdgeGd/kjSZMDplqPp+Iga5d+YFWP9UiKMUAntL/lvjTSEInpB5uopw1Un7Q
b1t9aADOKV6lBJPwjzZl6EenW8XjfQ0OMzwKjT6Qupg55fhlovrFIUgMUUET7Row
tCguwUa9EZoUvIh/n3aX4snssXMeo6hpl1b1K528Elq8yCdFRtJIOnt97smy34Lw
kM6kGNbVwzr1iX7M+ltx+He/DqosZTZlLtxpOI0cw+2PrkIBrm4H58t2bXVMLV0I
TrAv0C+9UWfKTWueIja4pzcSMZ1pctIDe2sma6YrxI3nYxQLgIUDwr9tjJ21UUqt
/N5BD5bdWpKSCGfe7vuwS6HbT/lboz9LlLqoJ7SBoybZ0ugsHegz7bOqmAyTc506
o3aeaxrCzi7/lCz3I10nc1fDpwobY71h9eUCicaKn7fkTPjIyJc/tdJ/hWdqj/He
N//kyK4KAD4V6gST6oaWU9j3axxX8PVIjdT9kipxjxT1ai8u3bUheCwtkd7XFhfX
ThhkcZwnxOiQU8tUp544PVF2oOT3WZkEZmJgicm2ZMoQx8zsIEmNdkEGc3Wyumjv
tW5dUoh3lN34TMromkBE2AboZ4oPx9BwoSsuGKbA6dNReyb2g6QSLOnl2iiS5z+l
57CV9Yuvm/lxxJtL2poiyIE8H+s+fCGmLkS9aXpCuYjzjzaR+vz01a924O6JvLb/
YkoT0qestmlwRjVZGyuRwEsW7ZFg/8vvbBH5xGM8ZhMA6scwptBVn7DS5ORPmco8
pIhXL2qJhfbI+OWyjuZUYZhF84QOcOQ8YL+OJEsy0u52WBKkOEE8+VggeW7/iR6m
ktk26KtUnUKciQ4JHMtVHXLJk1gVnyzKxOAs9IM85yNCJQ0vIGOeEOabrutVAtUl
MmVXUr7OdkEp8r6a1GRLm1ml/lRp0KgwnB/2QsxNOk7kGKMgBD7lWKizDTnMd98M
XtEqanW6Ncm3CQrnueizmeikxZo6FKoHdyf9+t24/TOK6jAzJFSamTQHYQzN41zc
6rNTPvcEznlBxwx9bW01CHE/9MPY2Fz0zUVo8tjEd6NC0BZYIN8s6aTvN4w8EWeI
avunaeI8fndC5ii24pkucVxuv65YvcUcb1FWi7W/PN+6SolLf0klex/lAvgE/i2f
kXKmxGmGkAYRby0NgANoo6Lt7qE/sPUhqp+DkbdsLo5hj1Won3yVTPBUob8VXHKT
koWsEF+6W1Q5NHF8gue64FHyN7VuzRDGgsCwbmyeXHCxRt2xuuGXxWL2TvIneMMa
FSi1Eh4XAEp0x9z751/mfV55LMpk2YTlsqemq5e+LEtJr1NxbtSn8gTI6rOpGXW6
OtZjaALsW9Bq+W6Xsy9rBMhpj3XFcvCdc/znfzW0kdjnl6aWekkB05ZkE5l6eoV/
fErM0jpPiOkRrble74OyIfNPpb1UTRUTcu2Uq5F4Nly46ythah9wUoB1eG33Rh0t
oBc8UpBx2ePOxwdzUItYn7pL/5irqYkGJhN+SyxapkaYEwf+6nLihUrhmsFFCH6F
j5Z/+ZQD2iKtDms/dcL/lmeC1EiNpIOWjIWjqIkrWy02WHBNu/tYIzbH9y2W8awT
R0n+TwPxWnI3AbBiOHqW7YA5a0mr2k29vTOjLA6PGV3fUOlsde/W45OsfaV7Xpgd
l5zmDu7SXlxK3+ZqpaWlL5QFFLfuKXh5X+WZL2faNX1ewTYmnUtsu44ASTc7s+FN
ccIt7yD9HDQV9e/O/52zy1SThjWog1iHK1mK4LIRq94sDKmlkr9euqQ0OvgCO8OB
TEMUrFMJRzp6CL7EdoXzmU7RbNjfjS3PXcStFIFQQPGB16Nh603yHcbc60RCkmLy
8TWan9lsXy9kiWlXtO+NB8po7UwnRBiQKmDD+SIE6O8brDnDtZowu8WD1HNY9ga8
gvpnTcyQoRQtCnXKR9yFOYNDikVmbIkx1qzj9NBWUZ88ulqo0bI6jdgsGzDYvFbY
IjvjwSTSTl9NErg3PBQxj0DhdVYDx+k+xdcz9/w1jootbm1CaO+MVlFulTJlyOjw
Uydl6KttZl8ExLzXVlcbOpJayO/KIn3GkYZXj66oqkm7e2e/9zXInmMMv0iTjVcA
uNIGU7Ev4yalz6jkCntgIDydiDD0PHdmv75yEcsc9nXhgRmxXEiES9qVlWaHNSEB
7Jx7ksbHM+K8MBx0hZSNvQHuzlJ++o+aEBT0qaOoSN5PEjw1osFW3ZQYcrTC3WvB
z2p1BoKxRMFSzS2V1naCu4WpEYWsTzPxeSiYI3qiE7nA2CpyerZ4OyP44zu+ZeIJ
V1Z5/fHWTfvkw/TUGeixgbdcS4OUz0+rabi0RJMOzsqYm3PkWvB9G0yG3Rv8m0dw
kfFZHi523q1mJqdHNABkiMpkWsQ7CyLqmwEW4elhntTedlGgBs8sHy6EtcTnpJ0J
mb5TBgA4nIxBpKSLtGHZBhrH9fWIBhtTvzSloFqcJ3PwIQeCoCp2KeifvTEDjBv6
Srt9NHvl2pc/MPWkZdNvYsYTilBUtiEiptW/t0mvb1BaidKx6v4wrICwARZVuBEb
RaDDKriScrtJ1/UhT0J/NMoZ/vYOd/u34KDsMFIrNaHKISOQ2JwLGnHM3YvIwVyb
cj2I/8GlhwLPQ62zi39Qk21LQ7AsWmJEqq9l1q6YxMclBMONKBPRrY9nlgf31y8U
Yc3+Mi/CkK/4Uh9Y/LZbpscoRUPorqp7blH5w2hjRd6OPiJ1dvEjkZ9BhQbum2gH
AI3o9swfXLJeKDwBrfribV/8/tvKdyP4uV9qtQzTxK8DHrjJXHM+hQFU/7OduWIn
sGNHLXOl7upCYJc3fpVJWKNuZIm5Bl8sWAVYjJH35Zio5PGGPwqbxSXNNFe3SWjw
+I1ktsbdEQtXQQ/DgWK+xMutRwchv1fjU4TAAuwwzTH9P5GH82B5hpfWplbWQZK+
YejvAR3sdcxG3WzV0aF9dH5ccjGiQyt6TWXDPSgOLmetcj2J80C04z2+O8Zv5lUQ
KgCkyFcgK1B97CtONXSgaKAjVnsu+lHLFs7pFJ7nS+yPNPdTei1u/6rr2YZ2hsts
dnpjrexopIFTWII2mFuBPXxs0zLbtT8MveXiwqiqIZkqz8WDp1B1p5trnifPe8xa
AFvFRBgKruw38q/Ymx4GpCAy6BR1LtmZkPtLqAaZF071jt8dleGvYl/ZHchXNJv1
5AFyYxws6VhHJyQFHtqY1IUWaIKKKLRo/En5jUqWCIj8nQwS1Io09TLYLIFIh90T
/zroYLkrUGgvbfjyUcv4NRbo36ksHOayOMBzAUQSTw4BNaSTJ9T0KU6bGfWzsMGf
yO6n38zcCzVNr2RNN40PRegxgaCiQUzUhS9YKaIBy2W+xQB+gOtlE6s8CfC8tfz8
lfKRaMApRbzwis9TQsxnIx/dpm01WmrRUg3iFxkT9/CziZ69fMOBDUBwJu5E2DvX
PVHflPryj/vm7fSI61a/Qb3z0jrPxpnL523SM3M4TM6crFJ+VCJBNryYOkRX+kuW
5Fe7uP06WNcWg884I0N9P3GHaSaiDI7UX8YDDpXkhN1fwzBKW5qBfX5ZS7MdsgkL
xzs62ou52YJcZxs3uXzlpJeqqQ/q6czzxwumMXD6Tqle9mcvkl5sbKLwOg5b9cNa
PtyiNwDhMnyHwwTiXiZutf2zc0EQ2Z8FeoyEFc7MZ6os5wsSwuZTdUK5l1hAm6vD
ZHifsQ2TMzGjAvAnRKWYWFKbB8EIMxvGPzTS+mx79zWUfTPBbKifvepq/JC9C6ne
s36OqbIf6hTs2NJ3RUPTs0vViQFEuXVicvg9h67Ussn3IsZoo2WdfWxZ1TcKvw+y
JlC/uqgfu/VHIrmMxDNaX9a6m6/9Nx60YyRhIQkgdQBc23p9FF+PpyKiZc8ImRLF
XRgOzIRHWBNMPnYWOs1reeZvpfRLjc6nQH9Xd2q3Nq9y0qRQcEpjq3Jv6vWV7Eks
HTfgGHHTJNEut80RwVcWxlc82pgnnc+5V+XGNmjNv8A4dRTe2Lt7J/JpRDlXFcgC
E2XOf5qtIbVbovQoE+5rNlwIp5Ml8qpv07tkYZsZpKyQ+vG3m6pD/wzvqwicMptp
8P0ETaH5NR9OFnTDEu+7brYf43gr2Ud+lZ+34r2TRQ7pH/L/SAhoJOTkchAmPZnq
3irGI1/AV7hXc1gbkYq8ADTXBwxd3MFaHIeFGqAzS3Rq0tXirjnigb/pR7o0UlTW
vMpntECh0CIXydOmRDRFQD7wYKmgVOZ5HLN6/dmIh9kfkBx05XoXItutcQJ3nLkr
t+Q1d1npFPmoNBzFonvIGZO2sO6DfnkxyUcmOjiFEQhuMLq5sofvuauIp85Km78Y
6kgONmB3SuxE1/pn6As+eoXGx5R4KNRl3A2OhA92bMK+NVE6Izf+PNgzJvjjcUZJ
lYGlW5LNsjEwSBb316B96EmhKiiVy6NYnK4j8LHk2i/nCqaJsrYpoknDVAO5s0mX
1mo1evw0mCpTgu72mAiprmm50sI+LnCHSXpJNsjGPm2wBjRHDvkqP1+tosj0aIvy
mwpK8ZW78DuWx+WhQJEgOH9wp1/NZZrlFolw5nN6Jlg5RslZs1nwLbTnsy3biQyb
8rcF4qSmtdkxKp1FzQem7/8ow2ODxn1b34TgNlKe4Y0jgWD6X/yCI15uxsyECDln
ocuGYTfq9RUg6yv6I66j0gl1RficRSrFQQgskgmjy7Aj7WDxZkXbezvSg81dlUGs
WIFCOmMYWwml359rrwVkT79Vq1b7CC+nN1dXK3kFWJ//KrOy1RfSS0/qj2PXehuj
VRBwl16sEPyvHazWD4AuFjg8mFIw1jw0gUk6naW5XEpvPtLXB59kP91iszSYXiOi
HvcjIf8hm/86ipNAhIGjkVT2AVZO/5MoNd82R5ZAYUVi51Vpw42ukey/2mv9WOtr
oD1bSa4f1wUqHCGGODaAsSSimVtXaCr8CsJOj8Mo/lUE8YY/gZYqUOJ0yMjSVQad
TFFJX0F4SPRDSkDsMBnzDpREowKci6EZSVqmTRsdpjuv9kj0yA1MNoIUByZ8sFAB
pA33rLNvjRHKkb7qqmSdDbCgwWeFMflswuHhXY90Xf/GcRlS97qWBTk5bSlQDJEr
gNbwdG8uRp5Dg0Iz05AHPhtUukBcHpFUhAD33Mp76z1N62qB/w4duAQ/S3/PoCoO
CO0LkeYlAqmwofuyOj5IC8olu3OhTAB3hQzYRXox/51sMSEy36H68ME522/L17OG
1opndQyopUxuB/9enkQ9mtYwZ0U80r+nzKt52LiGpakcw+xOryqs5ho32oxVJojK
PjcqgnYhIJzvfaAuC0UqB9dLpHrtZZCfgIzyvx4WmmNxgVF/xstyIhct7UYOpwTS
cByTR/yHhspqUBnwzl1TOcqRydNZCsL05J73vgmFGDQI86+Lb6+PUaGfIA53llS9
kdjfYdeAMv7mjdaEkDsA+8jkKQZP6utFBIFhwvJBEr215rJIMSw3LVbdI2q2UsOA
MwDcWNdrV4Mymsyj8Z628dK/9xU1ytOqUqW1/V72IL1Ck3Dm/AAn/eddqJ3DQLSj
SDT+0tbP+CfHUIl/hjMV3/ueJziHbV6hZd16UyiyqNqFAX3QLWTyZaCp7AAuI4o5
jYJdUJ7TOR3zvUvFUlhRWlDb7yMj6kLUEhNq6JdKH4jetpWYRSem/NGn/4LTJQ4M
YB8qHSkJp1VdgGygWKbDaHf2YZKieILRZI6UYa62IAITJZVwY8UJtSN0wvzCh8BA
DWi6KLU9LyKsmE33qzy5Lo8lxXcSujfQKyATDI8M/76OCDjRtHmow5B4ABOLxeO5
sO5BTeIfi5sQKpqrLTPR58oxKSBAbzaXmDpmBQsPDotpVAvamC0akI3pDmSRIrKh
5Tpephr9bPXo0rWmnXj6shveIL/3NjS9Xck0F2qauG6hni24hA5H9hg7kLYMfgDu
DPfdkBoXUlMR+eqXIMsGFOk3saZrqS/G5gd+MfnUhFO4JC+4eXVvw5jWnpAkMrFh
b8crnWnUky5CmNYr9v5Lschx+Apr7AzT+yqT2LIRJPm21wG8SPz8SUYZxubJ6UjY
s/M+f6zW/0Ws1IJAdtUOKl9aOtB197gI5k9RJy5hYv9RbPKSuB2TMYMNmQu39XsQ
9KAKcNiceCabCGbFXH9LhvZEpd8fGwJ0yB8eqhooqniq/S4vwWfhwhvg64ghVGSC
hcAZhxbdibnA2a6Fu7Y7ASQujXFzTd0fkbhbkgyxbKnfe+GZvSHpOnuYRUW2RvPV
1WTLKE0GAdGlqHjnySWEkQy+4nNqD0l4ga35FRH5IwTPU+KEspH8RfMqhtGcVTCN
tEZwLInzWjNrsp4ZVQg28AShDNiRvGNhj4CsCFwiJgdaSXhTLs+M0nzLSEVT8nPF
ApHD+Up2nUPlI9pSkGYzYj1BwV6tdfn5ndWXe9GINVnZMGQeBuEHs2pSqqwi0/Cz
l7aZoyuHNdg6C6P4OQzoKrHnWQaO6bxpP50R+SchCQbsbLqLdL0RwElHnmClBot5
v1uCyhSmxCjFI/S9Keim+8xAJCqd0xlPXI+N5GczjRZcveIDX8dEeLejDCqQwGtP
UrFaRktpXvlXWxnneTql+xdlr9nrh6Y9lOe6ldQIKPt4Dy3qE8BWIzHX0Ty45ZYT
pMsdAF4W0kKW0QDm3seIoFe8ssNd78vGcg4KkC6apz8S4zO3iDvTYXNekzJDKW1Q
x6X6KI/0XCEoIrA3U5Crsm0+oPsMyiLEkwkdHBJVEB5x5dP9cAq5RpRG9/P9x9B9
J3c2B1sz53pmJqcFKd/JKX0tzKwG6eZYZamA+oIwia2rLgRgywcHCchx5mItk/Df
upfZv2yBmM3f+BgB7b7lUl1lY6Dufcq4DtvatovnphTvGqkQ3Sa+cMc/tzJE7sQh
bKzvyCSMlVT5ua4P2ldKHcjg2awDgu18wPNH9I4hMYprslXI+s1+bnEVB3Uo67PJ
jfdWTtoiARWuFGpqRrPvR7FDSrqv7ZvYrmqmuStT6vW2vw41QqrsKI9586V/SVzR
JK84jQFRd0bny1kAS/DvWv5XBkPRvEuAt6VgslLjGAsCbTsL4b+r4d+BPU7RQDMW
0JR1OSbNYw/bogVwYXd5V6hE9zQnIqLLCOZEPX8+tEpPm0G5XnsQucp8G2QZHwbt
YdXtWlDYFeR6bCohGEBXUQv3w1wJgSL7VKAm0DFupx11DeWxdgKNAMUXHOpoYP6m
DOyxWwNRsV37loLRx+LVJstOTDA4HyRjkeHjFNwGLb5tOdhMxYI89J0v3+5RA2gD
ITCt7XIMX/Uwk+yDIlqkCWosRQv3Kzq/fxSD1BzweURm4QD1BNAgxBMo/7cDIjrw
4wK3U3KsDdn+VUlt6EXCnufiJYjjBNA18Gm6EKrDy3LmjOr1DbI7mPjo3kG8jTwJ
gCcv+ysRbyrYhAC5fqd8u0cOz9ROTxFI+Ih6kxNfwcWZMcx6gaR47olKlNlHC6Am
Jd26fEObT23UiqSwd3SHkOY/DrnOQHdollOTj19FaKKRFwY4U/jj4xbuTMKfCM/j
Ks1jMoLqyUZJlxqJOXr3LF7GC9cZH4Jr0e6d0W2NAiegESA9XLOY1m61U/O0ZhWI
flRt/VilCQUcTojjrDHHjwfk9bd7gDSrSJOiMrUeucUPjdnnDPiv1hPvHlWIl6bS
SvrzkPa9EC1pn3MfPhZODUng+RxuMdTfxVmEDFs1SyKrbqilSDFdhzDGcRZxJFpl
ktO1dPVfM4/DOXIWHgCKSHvzmP9/PitIECMD4W18NG12jhZpLEUbBkUtLExlYNke
dED1VGmkoADq0MG5IjwM0cMNWkjt8e0pvdYWwPdHHM6hVw1NaJTfl0xc1HdAXjLp
tw93F5XY6/EACLqCBUrAIIsAJfKKCEtIgApxe/Jcq3739iARJqBPZiES+S8SHTvS
u9WECVheECSDx1/VfzV0NctowYNIhjSQTJK6hn5ftt0OV3fi3xFeL7IAGLmMcjf9
AtkO9ylULYdjvc9rWiR7qJ9sstKg7lTVUggfeBODnUrTatu2bg06cIcLFhpL+NwB
CoFhzyMYnEJQElTdEPWp1gH7TNnFK3VeSwB32ZLkMWZClk59fZGDFaJJvWeqM2m+
b8aNPiPIlfN6farpGwYI6CyF8Kf6PYVE/TgcknjB/mcLgGA6b0IS5F416/HrSLAr
xCw0+cZU/No8iQbGuKvaq0RWGwXFlFYMqK19mHWU0YqoAGMbuDedc/HJE2CaKIe1
ifI23E4db2rUATF/ChFlVI2bQuFDhv3JgHjYCWsO+gmEw6ylXhG1JIicmtZNdegi
1RDsw9Phj/LrMSNHhZc/s1XMUbjtcdadOR+Lub819HsG9U3ThTpViYqkw8QWiJvK
NQgETG2VEPvob/5it4tYxrjfgq5dxL+e7wM/7Dz+1pmYqhyeEXdJl+jGA4AIpXOn
CyEpngNeNmNC0FxHWidgRadZPYV52w0t9ewfy8B1nixX12KsCldHdvZup2FkfnSz
J+etA3NekRqNIBtdIGG5qhhnFZTXIr7AQjxNEPMdzzrvNW+n6mrV9VlwxjCRoiUC
e5bEtOoXHHgGJ045nxtVD/Qymn5cwOoCz/1tfRXojhf+qWWsoItuMRmoNDvX2zQF
rQvsA04KG4Hf0bPV+DJM4Q5TKrqjHyXs9Lbd93jHsnjqU5kpIYOQSapKSBVmso5b
3xkMCkD9gK85RfZOM+T55N0rZg9kJCWaSb38uccbGv1/rCrugiPuC/86D3s9a751
pN67QDyBd2orOGG/5SGLzDk4DhKTQ9QWquPX1GR6G6j2dW/rAoxEv2VR+WDQCiWU
x1TZ259PsXwxdSOJOfPlrIkV6VtPh4KIhDJPqRTYAHmCu741Eb7lAIHBr8dVOCgv
0F7fx3/LAN7n74GQAEYDbjz/2qVWkrVPECqs0XFc4O0BBkGlAmb0Z8d3G5uh6VS3
/rFtNHLLGr3KYEMWtg9xY4zvI6akjqpUrAcadYyOKZwoZzzoZy79O5am5OQDOKoM
t8gCKzC1NlMU1TLL4eO3EbX9sKOa/FzfPqMHpZdqaUggOjrOCbaMP/qzEoy+aeNg
vCYksPp+lSvp1F+pHYhwHgUhCGtxC0TaW2B7N6dembHHQlmZOoEW47B09hTRyYij
QbzN7Z39/QGF3vnmWWc6T6+Tj7BnKGiHLAK3tji7P/np6gHlFO34LEte3nAbLayM
6/dHjci48G5AMrLJdcxXRe6jhWJug5UZ9S01in20hVfVjOdSkLHGUC9Y0z307x4E
oOLOyrj/pnzG+UJPngypAYHQKOystzD98rXA+PghIOt934zNS1ZIVfo5MHOyYTrn
WaFwdToq062tXVW4gUlnufX1Yw+tvPbzha5PJUhYKF12OguTj9ShgsVNNj3Kvil4
tbBeAekkU+HCZNStCuERt7o87t3dWtXQkNzP1/MSf1uSkVabkh5Ay9kYxzc0xGKX
5rAL2bhcByly9caT1r5z/eAJNfNSFv8+BbnFG47dspQQ5hWbS9Q0XAn6sK97zLkY
nsYwCw5j7I+ZZzpogGRN8P5neQ1HZK6SfiqFpsWcyLUkrsSl3lV4nB9OwgzyS1kp
kvt01AXkPdTWp8N0BYh1hshw3M9E17JOneyPwqKbRb/bjSLd6f2qGWOWkHYboYX6
ZEPM4O6ojAkUSkDelm52coqUCkYRS4WuzIQktblI7DGwgH566OdC4t7gMw8sFp9M
cFFIRDmzKMNO23xbzcQVedcNkX+FUdCvGVWBqq9Eysq7/ds6iWBSpcqfZ9K3L55Z
EqjXdkSF7utRPFYvwVTRM5Mjwto7zLZXIaQo/59kUHKVSzLVe1K9uCVd0zWqPQFG
pRb0xjplJtUdLIOK2BfQERl998lBpQfizIIBdsXDIIIwm+TT7yYgtW5V0cyWYIyK
5pStJKiH4g3cW96QhyR5Pu+hSgJOqXJg3UKFS+w8XY7X2bE/ds8jh5Rm/Wh8dFyP
ZbOKNuwWWNwjxEAzbQJrbfEg8BAIAAffdyUlix4Hwt9GOERcRRuCyr7U/QUtdjSM
JSEzz1iGgNCLamIEW+tvNoEPl9GGh+Ne7sW3zWGQyn9eZixrCwdggNPIKVEQmVPT
FjewNyNl8Nm34RLFRefyyaIX2wVv1fVXmTOwTn0Q8ImOFN1ESUiVq+grNwfk+j1T
aQtzPN3b8BPaWh/fq9LU4EKEVfN01RIRXzSg1+35Tz0PgxlwVEOMCYG17GKDGW1l
DJtaR9ViAg3t2XwgpQnnuWsrAWN/bf5gtSKhQeeFcOi9mCV5MUTO+hjKJ6SI1oG2
BhYxSTrDANHtnxxV5uPRMj3SXWWVv3lcXJp9GCqYPfDWFwhPOLCbDEMJ8W9W275v
LUmGUq0ra6eGxxODnBHbP7O+rM85o4S9eDLF1x5BBbT+8anjVw7RNy6xuoNL38Ep
+rhlZ2zLjE7zn6PmWYWQ0epAhUQnOqUHRlmNf/chPqEPUEnBMhn7tYcdrmRbFbun
/iJ+/19819VmePnov19glP7CfPs4cZB/mZVx0JShFocEaPGp/Pv4OFuj+6urC2KM
DHHhgN81kQKSsIlXNWXt8fOo8DpwNWoZ3K6Nl0wktBJNbM6iW0Q1X6+qRdOLm+zg
oBK4011FFPGax5BTpyIZ0xqETiS447JHXc6UkW2YpH0TuXXrRPPMnLzs+uboW3ai
dVtahrtmeGbgqVuTOjJ3jqNla3QVLRQMh1EvgWCHjv+Pf+WcU+0J+MOHLBCfMdN6
EXpNf+g3VGhhBeYriWxceAPa4hubz81Eiifjxq5G+tTZIcFh1HQGWIN4nQH/oGOY
kV9csgnvJqFqSwfDslHa0c7id9c1sym5f+IX3aLqJic0ES1uJeY9cxvK3mT85Wgz
3n2gPAfo14KPxmx4htzdlxPjdTQQ+3nF5tRd4IuTOgB7vC+gL2HR1jbjq37uwOs6
iLSVpJhM0M/UUq5FDHAMmj9KxPoGxZPpRcIacxtZnP9VxgrBYQnp7jUVxzf7Xp5a
RZ+SJcB91SjhCyXGjKJIr7guufUkKrU+uqjP7fhlYAbqd19rKq1P+u3CjvEGcfz3
XspQi+XZjNXx+ni6zj9PsiziH+UfYJzx/aHia/dnCPtYulNojwIMU94hTl7lXJRb
Hw13sTSyPy7V7deqmhT575cfHAO9xgWtiJWi0yUTNJM/rlZi3M3jXbRFfBJRE0Qx
wl4qNKD5H8FwGitoFv2aC9af11/+X0aTbyW9OMG1qds8WXPwDD6VPPv3/u9d5WpL
8UL61AlW8hu0nmtFTkDTDxSGac0RPe39Pc5kJ7//l/8c5VEyOQNMBx2SDTtRWbPE
aG4eGFCXDNZYXebj/nH2bgks6QnqyTxpcNaxLM9Mb7NiXeKJgL2aOeEhT0B3Al3D
qLtgR5FuNGRYsD9zC/xJvCpQ3s50TT+zu+EPy299MBQ/mZ3MJCP9gzI/qsqRbsID
6gFlU8IjgY7aY1dilNExpxthS1F8lEIVh+yObdETgU+825tVN6pGQp5oiKtL1Oup
Loe/jQ+I5Mko4GpFxB+FsBkeoiTyDxDJX6LwXhfRwbi28FgxmT5Qpr+tnE2/NgZW
czP1qn/efP05AOwqk2rVbvfMC7sKcNG3WinOACj2UflZWmw/G+US1FbxVNaAzXn0
IQ2JqY3mOStQi70rEJEFdAoxyQRVRpiUbaVbsLjYv+ibDRu2zr4iurfPwmCHJfs2
Nh63fuAifAWiftRNAyFhFCWOrWm5hnXXxZbcizHhMdi5vx4v+2IZLzdoq2EDl4JA
2lI7u7caPr+Z8lE+K/vcbqOS2nntciuKwN9SUYSRua5JXxHvatcZKhgjs3KBmU/H
TTR1hIGNIA+hkbvIwZAJ2arfcDa+f+NLtIG6MBisxsedt+WjQ/po69JH8DAK/ohC
YXUMIpXT1Ve0gIjVsifx5gpwW7eYcIhDLD69dialQuV32zWkWbDQa+eId6erWS24
ksM7SykT01NH/GJyLE1bnVszwmZiXCHoe4ne72BYCr2jBtCDyqjZtSRTjlUQ8Kuy
8Fnx7WQBvoJnWK3dAJO/O6FcU2umJvxkLj8HQjFcgXDom03u0HdTXllzy4k3BHHs
8qYcED0lQH4uZdTrvYcv1G8fL0F2dtAisrz6ZBSrqDLPB55BatpEdOfXuJty8fqA
plVSB9kdHdAyVOJO6UCl1sboKKf5xoVKse2AZ2PkpbdNL6wBwXYHjzv4E+93Opoh
JGm32UdY+Ly7OaHy/jrIrP/jFkEnwKRX8VmQ8Vf3NEM42XdmXq5+R/tQAyA5qtJw
uPae1BOsUj6YLXcJgJN2Db7b+/jeKuAidBDqHnS4WciLxea9+XjBmT+OD+LUXMid
dIkKyzJpZcNgEh7wH4ZrirwZvYnJFnmn2LKtFvyeX4yFZWwBVpN5UN76DI5noqlf
taRfFkFZNj+irDLqV91KXDolWCj54jdQVKGbeMJy6YMPc+GfgrXSR8UIyQruGfbJ
Snwz+4MgH3mWwXPBMcATC7MSzvSQtKK8eyRHZggGkYw0RB/etuyR5v8fuoBha5dJ
dLGjsP+zuAc4SbSESKU3soRHOYFOY/vuIcSv9t6xatR/XzXsSF8QZR+heC4Cg9Lq
dLQUelcAmE/PKDgtK+4dC0VuMDhhGmpun+t0eg29OdkZLLZK/G4LOqd+NO9Nx01c
kGvKPJwEyCoHa7H0/dvvwxF9UCgD/S+W5uCDk+i0dNyIWD9Mb4Uq9BWMXfEB/qTw
L4t+0f/og9tMvnq0gO5VDT1igYtgCTzz7SlIX0fP09/qLi/UPtv81wd27NV/vksd
0klkyQA/9f9NEBZEubdBDgd3HZJ9kqv5hIfKZ/QppgtFYJGh4NbYrw1P4kipDcLJ
NIqAzcyA/OauMuQrIjSeARmtJaCPX9CTPXc9YITSzoyou3GYzDowh1VmywkVwbxT
4zhGR70cSJsYgOiobsbhf9jYOJ4BSC5wKVs0YyF+xNuszSc1HEkjPJ1mh4kR+yJB
L9A+Skl2V3+WL6dNRnPYtygh8Shm0F3hc4inPAeEz1MtOKz2UInHcDLWfHDziqYl
m41dm6pIGQv4CLH4EnYbGiiSbjj3hfN/UpFCxNJLJxZd5WfkCCzwCoRW+y/lkAXb
SdoUlPwCvxpFhGj9Lly7EQVVFbLVR0yVQWvU0zhMLUddR/VK8LVlXCrJGXiClgqH
beMXxvU51qu53TBufpYBUN8R8mgYnggq/Nq+Qva4iJb6ClYgmP+3OJ0CQDTwr9tP
5X/b4GSZQNf2G/nnpDbAM+qjpMzubZPJSm2SG1YpIDPmmdR+Yp9lYsuwqhHu2zfS
+fRv3USFzV9zU3E0rbmtW90RmYf9NO8QUtQ5oLnVD4Eenz5Hah8M30fqrkaPBHmY
bAc289kYoqZSEOvfuzJEVBWT3BdYMraL/6LUHYo1utBCEHY/O8O7EDyN0yLrZKbF
zsb/Wd1Sz9IHE3BZTwyppi9TOPKA4e5gIuSXizjZ/K54qWZ1t3iaYpMB6XYxcSq9
CO4gjV2Vvi/Pm2bzXTn5+6I0uwAVW+1P+XHKrVb6EfhH73HSJrlSePGp+0uxd6+C
zn+2Cw6SxfBCp6t4tFvVGalcqUf2i5CN+DEkIK+80s2/k69vAgF3BfBoDWWD3SOh
bfQvhCeml/pLU0RQ/YhKxFNFpdlnYFPKku3k5iuEipqwQjm8nhCGAz6dCL6S48xA
6pRXhzMFq5EsjeJL80CdHXi8PfY2SXL/urAd7LUVzR4A+M6+J+up8AF6XPRNsino
tmMsCot0UJOvTKAxixUQpwyoZAi6fPFAcdRMDQN9aj/9RXgUr9W5SbSgGBDgK4wN
5Fu8nkc/eASMjD46qML1ZcWlt5BmEmZqofup+M/EGP+vSAki3L2hbA78iXOTcgZ+
GO1BjHlgDH2wPLQu1R1r3EuJlrU1TXQThN3UdPycjeVHmlCxFBJc1e7hmqAxsUFW
ijQR6Rf8w2I68Ov2mGEloj0ve0ojkNfRLjReGUvnp67nborMnkcUE/kD/JC0ZtUx
dQbAKukMI6EYVgkYhnbolyenJVBWhbIfP8Svp7WwWFpq7RCTBZ7xtbTNYPd4UCo0
yBE1F0N1d16cDAah/1wMkUraQVgpsQgBLyj7c7Sc3aFvMWo8pPPEL8Z/j7H/Noaj
6RfuguuDkMzSODKjd8gZIZkZyXyA0nVE3L/RWn3lGwKPpamzTWy2NBbYJ94g6PEN
3T+TBNah7fVIQ4iyjLVADKRgZZlDBfEURAUHXKkS6g72gTgs6zohPmNF/XWzx3pR
hRTHo6k4ivYhjlwx/x402DHhUMD4emqZfEhPHjZ74moj0HewAJMwEfwQdTLD0Dmr
HasnpLloI/QphlvHia0eSMSC1gSvG1yG2zDrngESYT5w3Ej4+hk1lnoVmmuT+X3k
3F0kRcD0YYgeu9VEn39GjzvD72316CmDgazk65JP3GR6GDauGeQifFmsbq4CImyU
wtdg8EZRML4vgcJ0y06lg+cAA0D2ZA0IwXx+MD8OkdHsh0z564WNi6vVHmOEk1Zs
6uukU5S9TZqPxoXkmn3UiFjvT3HPzhuPlbDsLCAGxLLPqcIYYmIrBHuAPftHmnKg
105deF9dLe54SjNWe+vk10shf2TlY/5M62E8JUwVca7yZAEtLqhJbkriYvtHR+Op
UjXBq/n3nChHtspMZfRiT765E6JZgKMooIe16sBwCog/af7pqdIm5pzT5l/kGmPK
4zaHNGDJZTDKn3b2JVKz29mDHbC/+/RV5i9M9CsVsWVuUNWaYQQhIp/DpChJBPI3
B2MW39oiP9/5Q/64y45+m13hO6vYmG4XYc3nSJZsJnzDsmLKHa9dCunLU2Ugzaoy
i1aOrfvwOFfaJcjBXYoSfzcO9mmZvpRS3njl8mel5qzB6LevMv1T7Fxv2oaHlMqO
YyMj7NKKjRHEIi2PdV1VybaFWvPLHXI6T9OQ1djzoXoYn1ofPpyqn5l+KmL05nby
lJ/60CfgAfDFUpxfTNjNYzLcMuR77y00t6VRLgOWvNCpBsbEIQ0g02++vmGAEp2W
iyTkbVt0btGTK8t3mRr2VIbaWBZFt3LTFIQV933buwMGk8JM5dC++pcG3kkIwQ66
lcAC6ghj/6V20okwM7cIB8JQQeTEfvfK0XtHN+YfrkAUnmJASHkODfLRZG7E0C3A
12iVQDweP/pqRbp43RKfTa/8KI+IG3JfklhiPKJmrokg+83obEBMlw7Ps82198am
Fj3GppZAnx70D30zVwYjdLiRQiTUQfPlw35k74E+QSeKE5fxjyjMwB42pjnl/gwQ
2J1MomwBszXHPuEPxmbATGeFwNf2jmMmKC4zsmCvv6oNgiF1McC7VFo57T3PcAyP
fjOJ0kMEpoqQArGOd2ftqvQNbGvx2sQRU3bHtXRAQX9ebmQJxn6o/Io3ap2LcCZn
PKx/zQfJazK2ct45R2myEF6v5NRRWv7Ty1hLeY+I1ZjN30qO/sRWROnPgt0ooO3M
gO5v5YtMB0ukUx/wip8n/THeqiw+sIJb4zqQUmUJVMuiItTkvGQ+6QsTQtCuGKB5
xGNAq8dV9u23dvJ9jzZdkdmUy5kIUmKpHZ+xbdZaqY4bpm9qDuxzW6TebU16kOL4
eHA4Jl+vU3gF8eD1R3Se6sPYYXN08r8yXsohG0NKCVugLW6IkpsW1oReClSADwA6
w2hY2tvZ81wc+PHHG3fVLJZKVSg52IJaGlwn6mrfiVOjlEICWteEZlq4DckVg3Wa
PPUJvyMtDlGjqmZeAlKKceEnzZcHiif4smoAs+uO2VzLVjRqyDE5b3YP3gr3Y597
D+zOxy2fGXE+Ty4iS+bddeqv5y0nu8AkehBQCnWJyBfEVDjCRgYNGGR1DMz5GaJN
1V7UFvJz6PrnWGAT19yHVNC8m6UY/PqruO1wRuCSouk7nA+mpg4cs2xR9MnNapwI
ifw9BdTOpvGqmQ9TASQq5EkEubC8efx5edIxqOjIPHvX85S3zLORPNgEropQRoRv
ppPfhAt7H12kio13HTYWckqxBmJJdp9pr4CXhGrWuN4S1fU55OjZ8P/2jkcSNdiE
9d3nLkuR52aC4w9LpQQ1Y08qaM7y1dMl6pAFj5X3QXtfCW65p7v0Tc0utZeRznF8
n0wA2go3JlSxDtbVEYRgId0gbKo09/KvnWiVbS0uUk+dQc+xFkpGRfkjR1UHZNeW
6b0F4e7tegykAVr31cNX8y+1GWFW32O7oZqiNH09JLzra0R9w/7pZiIF34t9XVUa
BudCajwCyYF5q3Vz6gza0YS4QqQLHj2lEHoUSsW2OGrUJDkjr1NDxvA+tcxfMWFH
cOnmJQkAt1ue/67qFJxZJLI0aYJOp9SbWOFqLcotqEkPCXoKTYEloz/C1BeoeokM
QTjZxQeeP8Xlln2wdVHZJADPO8FqGfFTQsJftr9gVaHaDHPTiW9c0UrFng6wTY7Z
TMiZqhWJbzSo7T/SPPEegIC/tNyfHx4P6JoOpDUvbkLWLAhQp9Q3r1/rQvZjqWHb
fFMcWoDsMjk5uXZDUxWzeqN9G7ktLSA2Vdjr6aOS5DWhEPVwPFzo0jujysdXK7PK
/4dUFuChaNUDRoCOO68AOTDFG1WWYCTD2R0cAOUDHMmo9+vl4/F9Z8ojKUXVG5wX
L7VYbw929CTjxUytnHwjMyji/qQL9yp3H75wcH73wSUXHV0XLz5aO31L2ZMB9gjo
03aJ5rCC58PED10+vqYEoMh/omjNbus06aaLVI20u8TMavBL/BDEfGDAmZhq2C7U
tG10of+Gft5QC2wpAv70O6yT3vPGzCkzRugc3f0P+ZDUogR4mR+W5voD7AuI7ltX
U7sIfoTYvzlwLeDp/MEXgVR7FHA+ycUhotfNdyVS+6FOgedJfjhhC9N/eaIcdaSl
4LEZPJ/Q2Kr1qw+Uwx55NhJ2+hvybCUhr1W1nZibxBW+LyjdyLKpxbw2mpXALN30
nqU4E+y6JLWycww16AaB26rt7Ookwg7tghsgiVJm/GUDrUCdVeMfCduTcJ8fD2Il
VQbVatKtcaLpM0wHcE0AW6LI6hPyZxJw3U0SpqfkYYho5DKRgFio5BHHQFMFgY6B
izKyEzs8qYDweTdBdAt/ZzihTFCZD2HJvzqkzJCJ5yZrM+GXRJtDG/Y11WTuR3K3
m6JLP4wnppUGYCuSKLlbIHbIrx+FN8oBWylhln0/ZM1SOD1I6f404odS6V3L4W/1
84SF71bkxPUWad0MstCiJiG2M2KRsGIfNlKAMKZdOjolTFCHNmSIP5MZOJQHNK2g
WyaaUVwSObnSTaHfpOlkFZF2bOyBx2f7voWXyWo7XLrBz0pbRtLs+D33ABFIqmZT
ypP8av1qvJy6LpiLIDs4MFhuRmYOwajPTCn7aGkc7ZSeWOwHqeZiAfT+2Xxuvtpd
aIf6bx2c9UVYLzqpAGN6wGj/qPJeljhlPhI+b10bGCB7WpxN+0+DstiLxPTz4I5K
10RHJbDErOfrUUd+hL//fk7IK6lEx1zC0KEdRFwDmrqFKA0fSNEvibATs2Wm69Od
1ljWuSrr3TMpmJemquSKQjMJQE1BrWr0hENzulKOPS4HZhBGagY9F8kEb1S1178v
QxV4bL3ltmr6SCqBP/QGdAz+mJ0b/t70WToehdlaoYmgsaJEzUZjocboK5rjarys
OUY1RqmPXtBj4ONhVP3evyUBRYipCrNEdDd+8HNn77rRcbJyyRjYFi2bkHKXLviF
2s01MM56BIinIZUC2B6HAlk4xIq7Muf31xk0zeYQQ7Vkl8jTUWdiOB2qOb5sHYAb
oZivdu0ROM8TmjDzmNkw+Twk5S1KYnJ6Vr93gIXAoqRJJ79idfWc3XY0y/TsTqNS
LndrQ5SUazJiNbFaSAcZWxmdghlPnpJP5ZkY3A3tisNXuUUeDB3zra7T7oU/gSqs
KOsh53GtQ27uzVoT+cSyZv7jHO0mddMyh7hJOwt5nhVm1sBT080QYhyafqpfgY+W
2afMiRr9y+yTscbtGnSxxkRl7dHyNYD1gsR3dupISu87vyUy3SAUaeH1+GrgmLTa
SZRskoKkhP17VS1rIALlOUE+wgGtSDzsQd1BZiSVuTNA/JihZpl+9hmE1GlhCMcm
G1fts0aGGssTPmA4ZF5v1nGb3LVC+pO2ZR0MGVtlR990+pGP9maDg23ifHOHUPYx
HkrAjSrLLNfQpOVunEnJ0u0YVcrCFHu8vpu4SJpLgtyThU6sY9k4PWwcJGWxNHwS
P+JvEL3CEbmPG8QczpA/FykiU+sFwlHymPTS0enqEy2CHmB2GsLi0x6XO2K7B6GJ
Hw+DGpvCZpLisqeI4l1K6FjHQ76wUpq8rhQJ5JyvzOz8CoKS2XaWirwac7QxdHXM
VLf5Qx21tFfL1tD1uQZNBylG11+zvudNRgzYMkQgjCvm09tcbKqgiafDVhmaLE4G
tnrzc77Bgf2ybF/TKQ+9Br5z8PGR5U8r8IxZwj5KGvrVjAwMR0x9JH8+9RrnWoUy
9y+qiMIUiNPwa/NKL2mJLesaAb+RoImUreDB3hGXujouCW1Mrxa6Vr57DYe4pHkK
fvIYeDEIKjuLawBz+I53Mqg6j6Uew+cag1tDZuArnzEooBfRp2qUC6g2oHWM6tHw
l8UAUtyRYmRG/yl28iwfwWXwGlNxEM4Q3y6bC87nk4tAKPnLWwnIiqtW+91qJtAN
f7N8dF9nwiOHGQekdGijEKB/NiPKirXZ7CLzpadK5jjoq2hr37we/9djK8EOOsUo
wWWAUIuBiF4bF9ce5uMv/hznzL/PUZk7lqsXcKGhewjEAMLDsH6N1kDSjtALV5Ng
AEPKCvrym52czjhBAc4ZuWA6VqpIZ2UqEfHGk8RvrA1H85OcNsJrIbf49oecxQvW
jwtRl2elEKn87yTnVztNN6T7Mu0nxTuwUwUxVEaUrJBeFIbeZtCKzV7ls0d39+E7
ct1CEQAYbhx3FwwKJbD1bCABZwIWG096FO7y84aXWRyAypq5chFyxogi4AjzcQrc
YrNKzYF92k2CQPp6e+2ht8k/67Da9BeNg+ZNXUMgzeP4QiQrkAsMhnnyL4MXx/ix
ikWebUqc9dxrBy8co3gwuQUfVH0S9ry4tDjPBTri48+vG/CXDODZohlXeTxU3x36
tiQNkLcjmekTIWnFZ8OVjT7kecMi0cDJVlCAvxhVIMayaggA6+impDA41nv9RRUi
BGG7IePuPSamp0YxUPY6k9U6wTaCpj5DoU04vD61r42Mj2HDB3opXOEiUMmJCzYG
kRGd7nO5ASpLZ8P8Ri//clZ07hwCMygTYsF8wiupIHQAIwvolPg/m2t4i0yC+Y9a
fZy9d82AaKq6Qihbp/OyKtI49Rr293uCbxK8kebyF6G64fr5p7jzyQoxdsBlsEGc
nNTPNi/fTi/160/BpqWrRPxl60b7xp7e9YrE/oL+vF2xJRpRCJnqCIzWHxzWkp5X
Uag9cExYuJe5PlJbluB/PoVWpWdSc+fpko7jlpX3/THE5wHADi38xja3keabH61j
4m+kG6jISCLBP/cyhnZ2LxKz4NJhHOgIdMU8OhdVD+K1zWs0AW2TT1ahVaayaJKD
aoZ05j8RY6kmQDekSX/ENnvcPtDXMpKLkjlllLCUTP10382LIS5QC3Q1C1Bg04oH
J74kZEx/TNsGOzXbQsQEj90Z7s4ykQX+I2bwk5qPHBSGPKSdPBFbbvI2kXw0wt9i
P1k5jdnUjliW/LnHaQgJxwsj0UbJMxc2jkw/g1LqeGx6qTGsKP0w3jPx5ZvnaJIL
CDjUR9rmc9T2M+lSnty1464ODbmhFAvVFq366VhveCcLi/o7w0AfmJDVO2LvpeOt
BGnQgNwGgZb3OKueNkEI3DpPSJgQ2oIkvrU49P8iDkbYo1p/E8VLWmdnibLBECDQ
WvcPsOuZiLZGmBprnd40OoKy6IXfmL2Z1TQCG5+SM8GCyO2oFdt8gS8ssV+0QBXA
UTdg9buYR/QKgJWmJ0LtqtdtxvyDJzntKt0T/L2aH6omakJP59dPi+J8Ie6hLcEL
MJOmRBaF+Tx+16+SPqPkISgfhBOByGYrCOkyF2xUcZQ7JInGdFlou/0mOr0az8QM
SMgG3Iy30M8AF0Hq3vWZUA==
`protect END_PROTECTED
