`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qGpipEwLDfEH3Q3Q4yz1sUbOqvjyh86V60A1Uakh4tpfc8RNferZ+OJ6MS8M0DH
X3eEWAs5bH5jO0oLaA5FNWLbA4LdlpGk/8nrO1BEkRJXyMKkGFKBqiWGqw+55i0B
73hmX9E6pxPEYIcW5/1uzf6jM2a/g9IEh1xTDQZIC8cVriuviHBsukKSF5/CYv3d
BGI7SfqqMcXkQoM5/VfCqnSCcPbXoENdH60UAmyFa2fjKRS78/J3yW9mm2RDk2xj
70AaGRxTMQzCjWZE4vEwP4+5Jx+T63SseP2QpfZDzUW6Hazms+aYvfKO/46/97wg
Z8nT91g93pGndzGfuSEM4Fkkou10IhFboEv7rNNP3qrFoTSrEiaHwKvHYDxTRmxE
s/Se/e73uiHPe5+VNyqwxFUyRvtt/TLmOU6WzRV93jTW0u/5vmmwq+bm38Af4/d2
I9w83VnlFU7z+qUnw1IteQVRESEvkH3T2lCDsoh0zvN8X0X/A0sAr2QerEloB7wW
coLjO1ZYU9vINJVNI+n2tw54fO/2gZ09fqFKJe6jck/YvbTTbmo6D/7HVHYTc75Q
rzv8Tk9Lyev3pZcTxnWU9mGo1KTbp+9YR7KqBoHKngDhjMkMNYxJ3MBfr/Y/d8b4
BmItG3nvlqCoL9kKZRM9XEX97Ixj8JA89BzrWywnJ9UsAY1xRlNZ37fi23/HeRFx
ABPxQBffjMNpV5uQRpuiyN2QVXENJtkynHV5jFwMKQ3Ok/3RIp9NpLCk9l5bDFE7
cD8ICjMh11+4BekTYSNTFQ==
`protect END_PROTECTED
