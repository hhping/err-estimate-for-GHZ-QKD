`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YygRXanBJQM6/j8FFFzVKgr+u2EsT+DyLKUcOPAbd8IVo5zm69iApGuyrBRzMap0
5U1M2E7gjLpsbm03fIHqfEqUO1GRTvSCLU4HthOgo+ZiuFQE7L5KT++PRohbaHeo
kQBiSgSsfmaLD6ilQ24j4ODVxkyXw0G16dIRFXNxXkZz/nnpb/PZQZDpf7tAE5HB
`protect END_PROTECTED
