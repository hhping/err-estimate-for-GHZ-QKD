`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmARAv2FXHxoBn2XZGEP90LEExEzXHDmOD1EyWfXFtF2m6iqi/h4unUaAuSM8Wi/
WxBkA2eznAymnR5q92oGpyxDd7tcS/lfwxD1gt1lNFb54NIQYPrrHU+ZS3JqY1HO
QaGfZi9XD/kVSy6d+i8NIsrn7++QHt4kygDmew/rqIrIUFKZADAHv3ovOkAlKUhn
bJyrp9q8oZDC/En7HVW4QoTL7AQsZrDEVQzAW8Hr7rs7FjeIrFgxjPYcU6GlujGQ
BtAj8Y/F9c4y9G9ElU0mPAE/NMg5U+X2waCbw6yL6NKNWyGBZsNeuRwWlcbJkp/j
Tb+SRUUguwlaEzBfrQv49iaxRCfpAEpN7D5WeTvzkzxjz3VDh4xl1iqfEErnx+Gn
M4f1n83zfSF+XaJHgBOne6rXz/3TpIta1HX2caz+JxnNUtQmALXY4+o5AhF3NBo9
5ByaXgvjd0TPgINM/VRKwfPtQAobUkz22pMdEtQksx6Js86Ka8NTSQ0+htafhXCg
3CPJKWktPjoaQJB+Lf9WDnMjKNLaPq8scsTiBPtqjgDhji309a3cLJZuk2N+l+Fr
RkZxqw3fDq04vwghFbDx/+dsmjSmRkO/mt4/Wr0wJDoef8QXO7lQpw+R9Xz95ppB
`protect END_PROTECTED
