`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sc8icd8v+NwHrMvBvLkMZmswNVQKHDnOMai3pryfwxnmgdKbo4Lf7gD5Q341mz74
Xp8IezsMdsC73KaykrkTFc0Qu1fc5UtRDvJWaMpRnaiVoOR2KKn9GUO7kp7G9GCY
2L+HCBTkBemfNQ8uRKXzbMSN2nMp9wSnf0W3kKHxEfYyGTOejGYJ5tF8y7+wtt3k
Hn/L/DqrgoRw07vzEY49sNyVl8wjQDayatU/ca5dm7tBIGnhhOBBMWIxfzMoA/Sa
vXy8OKB0tiBCDtOC8GQbeEu9gHG73G3cMorg6ANPPCRJhC5ohVEMOyT+SMk+/Ij/
xByrnCyis4nOaWTvrhF9OA0rAJ1sFE7RdhDtlX558Iw4oOFTlvKRQoe+Ji3DtC0+
R9wCMzde695lTBH01xaN2rTHZY+k4Gz2F6dGUd1yHQpWMLmDfyvKdnG4CJTKpAKT
ybxEkyedWUaIUqymOUyhCLzNJpnbMh/6Naly8+0QZEnqVWovhzzr/j/cfdRVbNfl
4IY8j8DMiqigy72LWxXyprsEdAFRnK+P98KG78VTE/pRAJc2RAfotCGvzWqacRv7
c7D6QPoFELMFCha8Yd2DUd+otw4zX7lhvPDFPFMb8uUQ8uZ5r74AN8M3mtF4T9Ky
R6kxI8n+Blg5K2ICPGQZIzrN/vYC/yEqHHnr/To+i5Beb30TwaBJGyUwhmj9XEN5
623sOpMTRVVOsf2bOjDydt+XpSgbr0rtkuU/mDAx7MfRlCMrkX+NGPEsJmEuQIYS
EnlkMakZ3mMKWPGHe1TYttw8p1qvLpTGNgzaSsrr/3d51xv3CyQpIWUZfb2mTUm1
0Hdxaehb4DbFAZkv466xrshppjuIz1DpKG0jyWjppqM36J9xLOAE3Hqv5+6M/XuB
`protect END_PROTECTED
