`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ifZwqnPEUGHGpWqUPjxaSIv4H9mfgB5cOqg6VIunRvxoLd3311uPOpjfrAFF1xX
pgPYq7Swca0JeaZQKIhti64ax6+05/YUw8s9Vi4EnkXW0e8jI5BJYmHaXTnVkYxD
lz4vhg/t0TX5k11GIf3mA+kYMIB2F8RTx1bSnqhyU+Jq1JgQySjfsCC2fB7arPiJ
ePUGy/uF8yBVRxXlwDAbyyPPXJJXXTGgvnEQw6PKTJW4Er3mokUD90PuuVBaEKrX
Ybo8HBZex+IUmdSzWY/IUOCNtdlQsev46hPv6xMBemaWBTay7HNx4W40JKeGjyIB
szrWE+a1cZ22iYN7A4q677RFl2gmMtu+nXhMh9Q/ddOQjLPZGEdhto7x+4kuwwq1
yFpcmvr2aSqJ3+HBcmWm1bgHAeXSBSBrfHuiUhXhaskpTPt0P0wwqTKjCMPty4FJ
u5/4gH2Ys4f5sEQR1Xy8pvkA24Hg7KqcCrgu9rduiihE6SUBkiQYUCZN7M7k/wUv
fgyWijUKQTiYEzlaeyeHjA==
`protect END_PROTECTED
