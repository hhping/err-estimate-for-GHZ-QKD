`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgcyKvbusop8seyCP4x7iUrnm4L018P0kcdZtLiKODmlqiD41ndpqQVnStfOcF0V
W7hFCR684NvuCdxHpZJb+Zcnq4ZgBio3uMZDE65JCQ7Y6Le5V4AqKDpUkmQL2L0i
6OFjqjyGfB/RYcr1avWathJzA652AacvYcXMfwLpWLTaTV8UiqM0mgbzNSaJ1K34
ryL4L2u8DRkKbcrVdk/AizDkwnHiS7hDsMyXJv9NE9CrmRCEMkiNQVPKd0c2/pdM
Mz7OCmX9mTCIJsaafeM13rT/8bjsZkrkFq4HWkD5QpFtKcPxOlzpJ36WeA6fqjff
dQBn1oYJcehC1c/8o5IzJv1Bx100pQFVyI9HTqfnNyRqOtV9foZlAudPn6cNfTUI
l+0XFxoX8XU9NuV1hggEHu4igdW1f/bPtBkT3UJyPy0sz9rXQ+BQJYMG0NJV7+hP
pZ+IpmONRSfHrgh69w5KELcnjg9xjMGhkQK1mu/IbKZsWtzWLTd6LaxBiyVlyT7P
Z4YTrxn7bB53FCDM43CDYDdZeOqAjEE3fN5HA6QmtBuwX/lMcyxbrQCGV9QJX626
NFm4Ux0I1cnVvwEp4I8iujGXb5n4ob+QA1fGDgsBsfQtz7NfVgz93I+p4FnJ6YjX
rT8YXMtS7OQ1UYoWVqpPYOFthG/Vphgupl8BFeQ2REYhS1oNTyXF9hVhL35iDjcX
3lXrI3diIxFqFKFuhpfuGiapEF7via/n9cXmCz0k94fu3+NjpOsrJUajb5h7x7NZ
TCm/UyWpb/4C8DJB+kCYOdrbYofPAUnVSBDOJoAl/arEwn8tGq4nkSsmDgLIOWGD
5Z/ypeuERbWVzNAMHkwXeG4mwhAdrZxIzI0cm7JIJ1ycyt/WqUXPkXSLdKgOIKKo
VeEHygEpGv5Zk6iLXLL3oaB+FSBd9jsmo+PeYl/gX1uHb79pChS0BaBri3pjXO4M
zE4LCkCzACn726FpS/Bn9Gx8kcFfPTqu4thMuVRKBfJx7GYiggw2cRSePiEXNWwy
EmgymgmQ1WIwrHv2f2Xb8RbvpmsB2w3X9KzwiVqyPwTcEUeFj2EApbwwMa/04Yvs
mGvc8IyPH8TfbVEXzZYFg8uFgTGn3oTu4ChPQZPt/axcTpmD+oDgArXqmd+3OXVV
yxkEmr9vI0hw7HT/0a2EXY/jdZ9vjmmkOIXllvhZxE/lSUEWeLSMitKivpUfppMg
zYho468jycwOAbxf5B4WIhG2cjvlhZU9GTymkzZkCVD2+QUvivWmyzxl6M+alN9f
pUA4Ll4gLZ6DFvweeqKWomWe29+dMyCqycz31FOXFV/+QpYHtzQa5TjLRPq77JEF
`protect END_PROTECTED
