`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
48lPFbXbtM0Bksa+aaELu3wfS1gOf3jMp1k3EBHHLbzqQjv6xUp4ocFa4L09ysGx
u6zZP61VMR351SENzvnYEXB6ZwvJBLBCbvELMv8inaLHW8uM2byB3en9Efolns40
C0bKxImwMXt5rDEmBsJPks+LojYCAWfav0H1VNw6fZyjf7PAb3fU1HmaU8Uv0Rdf
Jxl1ytY4fwXweyorq7F3FalVw9TZAn0TsRmkYtu81ZOYPVq760m6kOytRA+028G/
i+FANSWDN4uzRlYMe7vAb/W81bjza4ZtKW58e94h7utB9paCWYTIPB2c0nZ0pk8I
+Ll5ocv2t9MpaVYAVftE2sVI/I5pXeZsjCSRDsnw7Ovk4gC800sKOaklKUWQ82gT
M6KetreRGS6t97kQv/u4bzjhhRN0x16ZgJCaybop4ZDmVJ7MGqSBVTR+7Il4D8AA
Iw1gUvjGcB1a7RVRvpIxSiu3E47rIg+pGImuHj4gA10aaDd2PcocN1QVLoZKC23W
c15sq9KCR1jnMu7wdTsV1PtC4HtZ4wfNYdaxnV28mv1F6fES4jhBph9B6nZPZ2QC
7M9eZvccmS+0g56WR5+7pWWhDEhrgopK26WMqoCFafA6H4vuk43GQf5/gjvA+4Yo
0uTUJspGfz8jSxXKp2HituUzbZAWZZh45DcLQn8+FJPFz3Re+Wr5Mxyu+CGgmhCt
XV2HmsKEKjc6SPNCkkpGsq93yodVCoA+kOp9h6iMkV+Duk0iyef7vg0YpdLT+jqN
Prz3POtmzaSIP77++W8015gOMsBgE0DpC+fK3iWYXdagtyeFxiIv/nliFU91yQxA
rY1ung1R92deJYnPu75yGLXjCmCwjepEB0nnqpY6rlsMrV8+kIUZjPlW7h2KzKAv
S8TS3fEHz9553UPWgAJunTwsNkLv7JMco2JIgzh+KiMYBerQi77iRNrJeQGkEUpz
TUHWNVvMgYruWyYd9Vyulpa+oCpaKf76NsOKqt5IKkhdL4LKIYm30L/ZyFDCZqS8
FZ6F+cRTf4nmuZ8hheu432f3xf894zO34tfA3LSGJZ0W0/YoBYY4UbJUFJa+ykq1
r32zlY0pOTtOxnUk/+rO+sMPE0UTE9yWQvbxHSoelg2cR9FVQSyTyxxoDfDrD7Zk
m4hDVhYYlzWs9zmd/rVZx4RRECd1P38N2gKCkay4BCPVl9k8cpkEH6TS6eb67As+
OE8QnoCoGZDutpjpJdDk70iVsfs2iaqS+DVzr9kmaiicxLw9b1nhoRNUy1xxIJ5e
Z+DJIpMVRchlxv9o/KHZ4BeClR98W0Z17shBvjs3n5CWKAjzlJqSy2bQmOGmqax7
JggreHZe37sZDaI4mEc2L8DcRwpyQMjC/Y53Y46y99066y4xCd6MD7lS4N9Pm8nX
sds++IJdTVVSe+Jqz4SrFMEWpt6FN4lx4BcDGXo+Te8Q8lEm+F2oX7QD9uJ/VKKC
gs254bgAVD/Y+bKSPSJ73srZTDSquuTSgOPwknHtTPcw0wSCzuMUqdERZB8mpFi9
0fjJcnAj9wSetX8rWFzk20FWe3hMNMNv/xRNIhwTTzhj0e3JFGVEP0n9gJfnVBJH
i9Za0fqcCoFfrXuSClhFWVJ8N32Gy84NQTXrZQQHhGDuW1XLZS9s17fiT58lTUAB
wEMsM61K8uj4P31xVMWnJasprliurwRhAGAvZba3G0rLLWQCyWpjU+saJEfxioCo
0ya+2/72PEheO6MW7nmNHpFB61j5w96U3m+pnyNLNaZkXxKISsq0PrKkbkzLGpL6
1WJ7aW5eK9xvfzaQzBZ10rTHo5ScR5Cpekt8TLIfbLMMn+maYKOuvhwxUpO8Luwt
YrmNjYhVMgetpXk3hLgwR6QbkMNY4wHgoaXVf1+OEGinWz7h3Q8x2Xq4JM4FWm2G
UaTWgdR8VxJLpMvVj7G9PhphnKFZsmYehCVWmHMj+3q3mpO/fyl1ZaBQMCs72Dhy
oPXB9aRCNOvyQEAAvNBTyM4NddTRLD63TTNufUVjmz8hpmEbZ9di7PK8KFpSZV18
d4a2zGTf3iMYIXumcGWlMp5Vwun4vLis8RSbuxUso4jbaPbLXUosloCCARIgIFEQ
Be/CLaQm3BRB/nb6jJPzkAw5niBiWkInYw9+YxC/ATwi4/jLZUddgz41T6qG6cwN
y+tLMFWy5tkLzmDjjVSlO3kLi/stXsYb8o+zZc9TagBB+lm9FOGDSPjpWmoyseUH
XFfYPdS+dQ1uYYSVoERN7gOBoO0rZYAi1H75a4jkUaPEjz+mN/9Hzcg727LEa9xy
Z4fl+bKqPiRpl3I04WBYdj5/gbo4AMxHziMbipk97S62JL8mF0ZavSRXIVOQXAcJ
RlOv+a8gPtlE4FG4Iwws3mBOXoVq1+ENms/c4ARAKa5+XFzkhFgHbtnzf8qOGN/h
ISHWLLkfvqLVnleVUgKbTh+IbPsknPKM6naSdPVSXqrCPm0hIvkoOVJrtrlCCnto
50+VUKeKLkoQlXbLGG79LCb/Y1r7JjPyofB1lmrgzmcv6n9gGpa1JD9zz7zLfsGv
6l9UxZj2RNqdhOMEApuOYxs2iQPjrM+KdJX2r21QAwwSjmxaeR1eB69HDuuj43ZB
Bvjrtxz4T82zA+5OGyWawPXHYHZSQA5b2B+jsytA0BTAiz1ZZ0+vZBC8LFI2hH7L
/D0M2Kzd2imqgQFMTYzZQLD2vOxalduJNpb32jE/5sCelRvSTK/UOZ3td2T50dbT
bJqr10vHBPVRvk1H3gI3dPzKIaQg0sKFebZ2wcmz5Y57SQkXLKBo8QZXQePn5lVa
LJ2acQ3PMI23dv4QcfyT7Bthh70rId2SJkBjmqf+J6U=
`protect END_PROTECTED
