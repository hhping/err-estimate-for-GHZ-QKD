`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/94xx+Ns/6dvVKJT4k3tiebQOwG/spSBL589A1FkqlYhJ9SqoOPx0eIZW+5IIaos
9vNIISE+fjiRrDg/IeZRIHUs0h4ihOwZmFfZE+qqQydRTXuOHGgPEFLGGAwGLs+O
PI+mEGf8qx0ZUTMjc6UB2bA80mJ+cmUR0ZdQvfHU4Q1b6+xFOYrTC/YbLiZqAYC7
hU5AZ9Fw3wfSWlAW3SUoG0T3wj8EE2rZOMvKQ5ECN+zq8S2GCW/zTBTgOt18qnJT
nK0nXbgrV9d5dSlEsOuP0wk+NVK2239D5BNA9dhWNM+J75KRclAfzRyjsAlOJfnE
4JxvyLtSSrp9glOif0B1cFNe51DXC5g2Bfi/aUj4Wkqi8KXsZk7zA7wp7NeHOrNJ
ETWc2ffhRKCvGQr121jwRVbKBt20gJ9Ut5L/Fvs/T5CFJI0C7FgNdFyDZO0uuogb
20t4/aMRxqK7//8Voxs0DxQIPTqQ+T3jeD494wxfUCza3Lavfy3i6xr8R0g54ghn
1xEUO+xOkNMc2wHKr9ZLwGVYNPt0KCkau+ptsY2KXPf9qeAJ+vTAqP6ogDYjYpwD
JI+FV+EAOVWxSRDDWV19QXiuo4vmpEsW7O3UYd5VQaL9JsceUSatms5cCW+CjDYL
MaqHK//d6FH+vHwfQMQnl4MW13vcoJQE2rPqyOaBgEBa/lEP4T/cJrSwZnBhnx6w
JpN+qWuw7DXo/EjBUD1vLnXpGWmGSIwOPApNZjKtmxh7XcIrzy9LO1yeCeC1zt35
9GAllxeOyhfl1PsLiTM/JtHN/Uw+z99d9aHza+s75anq+3I/BpGc0agGXQePvIKK
TjkUPLyBy6ru3GdJ/t/EOxCOMMTj9XGT2Dx6UnNbt9hxQ0UcZEjgQACKLao9QjOX
8OdrQRoz6E1SqIAMLN0PQjoCRxJP5RPLNo7GhXU2zlb1qhCFTwKDfQds+Rzrdvsn
mly/DC2ReCmL89jtfAaCW/CH6uT6wLUisC7FKGjbxhN686Y416+IRmgvFkNbt+an
EevTLw7YRTlwQyalvE0Fsqww8g+/CmSgMBf4s2W0Qm+i+DekSihrcdBEQc4DBUww
Ogn9fLRAC6YrH0SsODanRk59IV5ANSehXMNKPfRce/7Wr6HALfaztp83alnbZmjJ
co5+vzPHopzLmibVi25ZOAoDREqU9hM5t+bmi0Uk7IOkUDGp9SYFa9E9hCN/a/pT
Ot8Du5m7neL5HUhR65EVWqD+sq9L5C01G56epLdDLsL2A+gxiIcHAqE3XDriXZfe
SSyYOtQ6HaD4ZvwKBiyRA+aYRyv99UoTBK5qLgZ42kPTb4Yit4gDqQD3aIh7wD0x
ubtJwCo0b2rUaA85Lj/lHTkepC/vn0BI6bJGsx8RNZEmj3c9JnAUubftaGyJWFFG
Hyspp3aVen+Cb0WCYZp+jbqhhDrSrxXlxJtjxQ4fHgWZbDUm2nuYb/8z7gXa+2Jc
pQ36QiZFSCEvVQ2yG+pZ9GGopKaKUvsRvBOIKPUVJuhC2+aCG9QG0rVFAz+iO0Sr
9+wL5C7C+qFdRbgXSnb8hVxRu0Y9GWbsLRqiIfpnkruPcW+ea+x3BemoNmTD22aG
zKmMEVO0/wZuY2snkt1tkSH2rqg3i46RFv/9K2golT5o1ewxVypXKJi1sr2Vsi8M
DQ6AlrzlQza1Ul1aGY+pNwq5tAwp/CHKFCvQVCCpFTlqkt4x9z5kU5zmIx0Jj9b8
wofrYernIu8zwm4uoaDUN9q1UQdx8J2CqGHolh9y3/eFJgQGDYVlUtBo3+x/CENf
2gaHFblg+g6OwKY/GTletEe7Q/BuD2b821F7krnH6YpocqIdsYKTTOJleRCj0AFR
vzaf4nqmNQt1SxL1c0C4i8CU7INzuhfILgTf7M4tuZX2asB8SF9+wq2Sqoc9VOsZ
nrhU/VqHnCNWZmq1duBcM6hf9oBGxshuFqPTTc9V/H0usLfWYkX6PShTXkcm6sac
2mZCtqbkWm/16kVHxRufLDKVRMsWzX/lfUdof29fE8+dU3vf38CXEdhCAzUJPXNt
vkr+4l2I/3yw1kL7JYkaY+wGv/mH5NRjb8zGnVgZgzPruyQtc2i0zUt+6aTGrvQd
9NwT6iAtmBz7aYy9hCDJjhiHTD65LbZWnveJvGl5my99yshqD5QbedgKiV3SJvRH
pR2O+6ZSCj5g0mN/0RUjVJ55NBqY2iZ0aVROCIBmvCBhvZR3L+MWCHnbTHk2IUxT
Tv3G3x2Ge4Gr1O53DmAd+9ZSaxYZiG/pn52drFJmA2Ud/ENQIKGREkH+x2HnBdCN
eN8z5YV5UBmTfw1QxlvR7sZkcOmQ63prKoZimtLwyYcJ6zPUCJdxo4QujggaHtqV
fXJgM8hCrJBm2K3oKA6XH+rt7clNjniY5H/ZpG2V2Oa+GOHk06N102/aHw7y2fQ3
l6tSSC3c8HvUf1vlqVlVN1ezzUrmzV27aGj1slr+Cpr4EVT7eDijUgi2pul/44vl
Wbda0nvzVKOW6PpQ2Otn2rT9E7ZtpGB9Sil3tfURb73FDuxRmuaxmt3zFrefriYX
QBpRl3DnOldPmhoH7XowCLJikdCou2/hye5ZJueh7p8QFw3O2FrGuWzBQAX6NgrT
196JlzjLpK2Mb7PmJe2A59fWiWs5ZaI8Qv3Vik2L897ENeNe599jWiddyeb0Ab17
+W3pYMde5XCG1WWkLULlGR3m3H25ChOHegWIxKJStF4=
`protect END_PROTECTED
