`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWPo2kHR+AaIf659V2xOKLBAB6Q2xHR7CcKUwr3Ge1bZxbSFdXjG90DTCIm4lc9X
+Dw3H7ILJ3jnEyV4QTdLoOLGZULQvehrR8XcjGB12D3IuZASVvFk1PXi0bDYL7Ik
sly7lBiIUFLMTpqq92H9OLVx3XIo1xbDnDwljsgkY9rFcW77zs4HfmjIRoUSC3tu
o8LTfo40Y/1SohiVKyyK8Lnu5HbKBuB+mR+phq/+I6UFfr3r2FXv670P0btPFa5X
/ivSBuXWSoXPfFjLjch1PBpdN7AMZMd4t2jaD9r98RCT1TEvAEepez6Ogb5SostY
g+Fwb0jUdn2BDB9P6xNIHc4YwIfgQucMHAnWnfcOBA9ISiTkOGLEwh5vhukZWcP0
UrIbvU77BSwYZa+Al4+jEIZq+uX3OMdBEcdE3r4o7P+o5M953b04k093RIB6b4Eo
35AjuwZ7Bbc21+RWSaGt1BmL1IJFM420EvBKovz5Pi4fQPSYqwHUmIwjVJWOhdwo
09+4m0lvDUB6kGiNNvbRdYLpHCMx8yYYueKdNhfMf4ayqSnLaEq0xojbP1gyymlb
zfpcoEDRpR5yZqWBVjSsNKrxqbQwG3KR3XzgYN+9VVoE/u2DEUUkFBU/1tje7vSM
olm2YYZFKbh/eFKEidYwk7MMEOsmKSFn9wJ4IYKHzyVp+TLEwvPQbbKosSo4TMp8
eE7iV4yICqRN+3peOcQauQ==
`protect END_PROTECTED
