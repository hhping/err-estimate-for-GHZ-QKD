`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AraxTAyz7YlnRnQnRYGOEcFtfLG7O4dOyvTykaAUEuDopCxtZI4gEGq8WCCZ0NqB
STDe7m2GfgWPkgcdg8OhCmljvYgYsgG22PWQe3dcGBRL3Ih/W4cnaOPMlgx3o4Dy
QMPQclphI7n0FO7Hz9Q80bx7k1CQIwVu/8wbLV9djNY3r4DGuY3K9mYYid5huE2P
kbvRB+UurHrFtNK8nUmlBDAvssdvLyKSXyOa6dgyILYN8gI6pPjRP66sBMRI8nEV
Tkqbd+lrCAjlvMKe32/HdhN2T0iZmMNbzTv6hr18Ur9+bmsDh91oqfV4NNxhfIl+
+p1HBHUP98Zz1X3qsgTa3DUS5qegXFzdSfZBarMN6LIx9mnOoQxWG42bTg3A0tm+
gO8q1SEPRmwPW/dG7y5Mcn6qE2VoiZ2QJr+2EkDOOzaXyTVCHo3spaEeF8cpfuI5
6cuXPv8tMN980o34RJ/PKLrAoP7EDFnqXAY1XCUAa95Jk4FMDNQX51iHQJdbcpNk
TZpdBzD5E7qg76ef2mvc9cM9luABn48GQmVXgv7KJhQ86KiGDU8BXlS/920IKzyS
EvpMU1mzJ+pg7UmZbjJIO1X0sqkoBUTbRPaDk2cVb3wD5wenPIkyfpnpHul5sjXF
FtJaE6zUcCyWwAyLREXgt1GkLmSEi0E7wJGWG6uWBwHrRImjIs/GPae96MftU2HO
i4QyRqoQfDCyAp0xr9q0Tw==
`protect END_PROTECTED
