`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H35/JpVB7RxwVwiwjwd7Qnktf0KrECGPXhBBcpb2/A6IiItmbC7VQXstH3b784hX
yj3W5yg/yQ9CjHu1KjRqhyVqsrepalX+cxN7urwm2GVGHtfdPj0H8ZbZGqqlKU7Z
sr6lu76CvCeEeBkbR7VajK/h9ysyHoaks4+Fz41Zphzk9h/xMqnDY980W/lNfTDn
gQ/ri/YXgiQ5GZzAMxax3cLKrPXUEH0fn1yx+p+/1KkxHM2Y1MhNI3dN0sFs0NUO
7hfiNAvpA2g25JhZ2HoSEmIE8mmoivbtrX6fVYXs5hwiYJQE+nC5jh3vtFX9PcYO
clkh/C05xXCI1NdsZrXGrPGCt3KgfPlShN7m+N4rAPLxH7FwBeEL4xSdLeMx3oR2
suDwhLjF10L0WhFx2Pk8FHg0XDDwo/MbEUOOMScA7zXu8b7eHSyU3lSliPzuyrIS
qgERlPTldbvDID+hgFkLj39jresn1n49QsowM6+GOSwRjgN5L027z+ZGBi0sLe6n
rkt7FFeYw2woFzBBnvnr6C/ucvUyCL1vlCzouKYmGna6sVS4y+FOK9Fjm0yjOaoP
ce2sw2xKJrAdiv5DK/teLIhw2Elkd3VVw3gDKcWsBgLk79G1eLRduZ4V/la5NCYp
wXhUX5RQjVYy/jXpVnFh1vFXlBnJ+N/qmu9kCObDFXEniruCFkOKlH6rm0ZX9i+/
`protect END_PROTECTED
