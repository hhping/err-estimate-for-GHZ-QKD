`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJItJKBgmkWcyVsP2s9GXd1c7d75r2CuQrScIF1EQHVpfEYUVoWphUQSFzTEww7b
ylKnf3Rl4TJKxoAE4/HUasvRmAfgKGA7KwMNEoaFcYCTyKSExL2zgNVaMqzNziDJ
vbV+S3Sdk07TO7Y4VkWllx0FJH197vnThMfgUfcE5SGAR0+M9OlNtATUaUJCBK9N
e41A3mzG98Hxbdbt+Z2Qoj8o+Mu3dEbArUFvBGbkozUgLMdpukldIfGfvvklQ/AZ
/u6HLUlwAYNiTlhoBtUMVHS5F/DYKqFzAiXyPaAOLc7Mgxm8bES/OE/p7moEKvFx
8luR5LpZyjMnSbd3wNy76B6YDvJ2lFj3Wx+UgmqLxrL//BNizKiucR2nKSvKlx3y
sUUQLt+ZNEnzaNiK7Z+G1gNlLzPYn7JtaN3DWekGDzNCnj3uYCTOmMl9JhDgtmBc
TjDxQcW4LHlBRWkpgkQygSKnLufEtzZR7LpJ9roYb0yfkvwKAG1qWlp/dYTb46oX
+Ul82rt4KfkL3vweXsWSzoGcTrTyT5SmDLj5PkD6TA0ibTO8Y7g9gsmFFYJ1MaFE
Mdgoj1uQ7pcezjq7Q5GpL2VpTbKTfv7eBZg4hMaI6V4CB2wTY7KLBiPS9VQqGrvL
N40jjn3gLF1F4FDdBpOH9wf7QT5iUCTooL1dWgvbeKZtoGOTIU5KGW9znXQzjO/V
FpGzWu3MveDAosX/bFIpwS14DpzJA2KQb3fit4JdMoFZTEY47tVQKwgrkBTqG45+
PDMQOgRYc0ocJ+rAEmWtX0qAl8boRsXHCO9otODWxmQjI7A6fldeTnqES0oXAXIg
51XnoRpc3yvMKgIGyZmCXJyYwkFAwN9Bfba8tGdLQcLX923um+YIhxEb36T8SRvG
sKhl30yNplWLCydnT5jq/4rS/CGhpYcY3AC37YZavY7nBeZ9qNQqyb24sDaYZOHv
7inHyWSjig43yka3YwFoHSffjR8ZPgnFy8+/2zOMnDhmMgIHFwiNU05RGRJ/HUAT
gWRUQasslHt8SNG7yoTB/KoozurSeGMcK3Z58cwnrZqC/sC4pjmZgl7zm/FKD+2O
kZSlxmcFgatVbWlm2zlMrqiAW1UAiZWwy0ax77HIcM2jihkf/wVw2Y96jUH0u+Bd
Azg9yBE6f5HkJzn68ci+lCcqPYlm732jZRYrFnaCeOyS1bI+uGKoWhGUBYsGpR8M
xTHTGxKSevTQWsFi8ekgoBtO1JC9XXXl689s09xum5E9xf6Ziw8hekiH9Y+PgGcp
cCbuFU5ZoSvpVhQlSDQy8k1GQJoV+zR2W47sz4jzmI0=
`protect END_PROTECTED
