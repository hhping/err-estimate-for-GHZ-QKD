`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imLpfZVpcnSxSFplW8QJWRapcsvjHnmueEORMEF+6UyCMFb/18P1SmqRByj0ZPwK
EqGjxwfap6sfAfKs7NXoURTzBB8uIQZMq+L8Jb6/sNNHJRWhl6RlKnpW0hoCK6VV
4NRSRUvPf2dZWzQBWCboRwh6voMyD4weidNMJE5ql3iFRC+DV7uZ8u2LvB1d/xGt
dLvK2T7/y2FllDNujvvtsKFrPKwYU4FjR3daaZQUrYF8CRn6MK3DEDY/ZaYRFqlY
lggDWkexzS40jTEWGk5TSk+P5r8QhJnBEgj1iqgxEs2Xq4T/0WAjc+ot/0ht+cKu
9GXR4onWsnmERKubK0xPScs3LfvtbFNlVurmUjUF7Q/LzZGD4jjSXKVZHuByZZsH
WHv7L9p1I2zL/4mg//q5ucMgPI3oiIrXUujQ76xsz9+dSa+JlAvWN3LC18LfCd/r
2O8RWkDOszkuiGEfNDUjliGI/MDGij/aPmt7r2fd2as+Y6UwjnKUIb/s1YalhInW
mB6/LOhm16WDUlqPGm8t/BbBzwgyVwHj8lZFJVAMEc/BE6nU6r3hIto8mp+VGywh
AGrMA9aDwJC7m/25P1VgoSz+a2tqxQYko30SIlmWxVZt7kqL8Fq1Ak1XqU8Tscvu
JJ+APfDDoyEZYJ3GLKHtvHehkm2puRuOXW0IHw3xStuRQytc2FxVwlGmmAVaxtxI
4hKrUXJIaIp41mpZQrQ1KHUrBW6rK7I1dK0/nAp59DSZ7WCq/T2rkK+d4ttHFGRP
TAIHpBkzDHyJp/BgAwryMXEW3QnlOf1ieGuaHl1dyDPq1Z37OAp2PSHleXE38W6f
mK7QGnPfy/ywXD0E+CY2knUnqFTaiFobsPGUuX421DAt4qMcfEQ2gJHeaMsgzvht
/xn1zRvHYz29PqZYUuO/EchJd5XgiQsPGGXF3GQQlDzCovfJZ8RLxd8WmRWm4FdC
P7UyKcK7vy1jqO7my9YVgQ==
`protect END_PROTECTED
