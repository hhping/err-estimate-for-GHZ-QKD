`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IzjOQSWy//JLi1icmkFDqQQP6bjlLlB6wYv3NL2rFB+mVvy0M7GBvoUDYbOt4gNF
woqN1XbDhXo2yEX4ZJkXJnc9hPTc0ryMcKWa2tPrAR7dUYcGCpNicb0XxQKLEig4
0+INAw873YiG2OtRQkmtRNFIlFMMbynmsMOkokSZqjxCd0Ws+Si8mB2NuZ+no5mf
joQq3hlX2FFNaerGPPD1CQ4mhyhWqWuuNY/upovni6976BnNqWQMrrAN4PV/ukdK
gt3DYfpzWo5WexvPPggvjoZZrOBvT8mtpwF2YOwif0uy5M8DlFDbLmzl6NwkxKuI
J1G3IxX4XsfXOa0D4Yrv9Q==
`protect END_PROTECTED
