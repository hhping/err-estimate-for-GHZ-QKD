`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYk1BSqYC/wSHXA7XzRPTYGWF8VsDGuyuHqPlDmPpE1xDwY6jTYVHVBbDCq3mPy+
uGr9QmNacDZaChNWTs9Q4XTTRatVWFGQCJ7GpuVclQRcRByAJPaPmbadngdqGuHE
hp159yYJoTCrjrbASpuN/jLuhQWd1oZ1/+ofQfH9RoZihtdH1Bmto4OoYgGPbm0e
mXu/C4AM/u1DDuc04a1ocwr+UF++3TqEF5fBfTeg8+g9IS41/+7dByEWTGj/uqoN
lzTH4eQeXpM+wsEmkLEy9FIBdI1KVSANOMHRp1EQfDYVqFew+wksSboo8ek9bmn9
M7d8zGulJK//MnFFAWzM+at7gyjkgarDmHFfIUjTIwEkXueOnku3StUlqJ2sXFw7
mO3j2/4l+uaJ9Y9r+NL4VmCLEsZjbtdVnhStafMMMg5LxpySL5pusHNymnqBhJHD
jksQjr+DNIi2BrT2Hk6KLlfLV2rFkrDpwQUktebBEo/8n105v/IX50o47w7yXQSj
3xG4yuxRWw75aa3UZPwnQzN8GUR7KjyeDOo8YVxWIhAPEaoh3ILLEoI3Mf/rzcuq
TTey994j56ARd1Frq6BfTTESwztNI7mzXhmHLRHDYdsFnccWl/gL5AbvFTdTl46a
JPSNEfTDTvlCwAXqeIfT8TcPMurXuqxqm2ItxKdyaA23HhwV82dBXbacNUzIDWkH
bj0t/oQsftA3JGwVXDJZNQr/kze3eVAIfs06GYd+tAg=
`protect END_PROTECTED
