`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRfdYikoPETSUsSc0S3EywXn+OvkAHxFrYasccLEkoc22h3PG75G2Iz5L+g1rUgB
2wSNlkkH3r8lF+L4AOhk8dLX+nILq+IIOiwYieEmEq/uj/AFlsnQVUrI6rm0NSHd
1w6AqGMbFPzbCb+cWDUTOjWYk/iXw3sYo9mk1+PVsIJ/UAbwPKJxDIngj3miYZX/
wwoCwpyU/GhB2AYDm5ywQ2sLtEEyxoFDpt7asGiZ9KbU0TDQfmlQCaX6ucM9YDlv
fjX2i82kFRrLOa+Y9+GO5pNEY4x838pjVfK+GLpVqPhNLkDkt6ncegKa+LAeQEJV
0hlvesd9vpnNGp6bpoc/p2FwTK54M5mqLGFPX0e8nWWkpZ56P1uT8Rc5t9LEMA/3
Rda+6aci6qDAk+vEWt0JkFjF0qbZXA4KAJFJiTSluPgK2E4SQyqd4eDWc21JUroy
mtqqINSW6UsXqdPXc+0VcrVj6SeElqmMZDGn/vF5MaF/1Oc4Dsa+RQw3sUZhZ5gD
xh3+QnjqkeZyMUjWBpiUDP4Ekt+nFQ/ieerXAi0YnGlcTdPK0ib0Qq/Ahx2yCMKX
OYnf4L4DHEWIoR3StouQAOv1gmq0fveW2qqB9kmnZIu6PAUY5h6AE7PvvOuFY77y
eJql+2nCifUlAMeQwndMkdsJC/4lp03AkeAITrVUCrvR3gHr42TobLyCxjVuhOZt
s2jBh03oArz/eE7LFPP1XiKY1TxXSBsDehMdJFToFh6JOfSFnPygKCFK6pINXR7v
Zo1Qb62CC0foXxJsQ8EOebdDAek1KmS9JdPQ+lfHp/YG1+itOOdHM6Vv4GXsPRTn
RblqWAPzjwOBfb1LUePcZ+ftSSKj005BfsUCACUI5kre/pnVjCBMM2hT0TK4+EOq
npmnBp6OUBZ8ZAvERf3m/wH067aMYHl9DfeeaH1uqIxDfbStcBzNwv45WCDsJVls
ES8lSzyj71IJYiLFdY1NBWrgBUETSN9B2fdscvkfGFNljVYg1TEpjAqRn7laU4OP
uYUI8zo8aiinFyNNVCXzXRX2FU//MJBG8f2QiMeVBNIOG5uB8wVZRcSteZEn8Xp9
XVw8X9IQScB0C3DBDrVK6fdMd/DudA6UJE6iFRctxYgg9HEe0QeUszifFcaB4cfq
HEwn5OPZLLhhekYNm7WT6A0pm9qxzb8mvamYzkPhSzm/fBuGZ5RaVu1kjMWEry8c
bvyIGgRA7bdXM3V/OFhrntls4p4sKiTdAOtqTO4uFE2CgVIeDj8+apnWivfwLTDm
A0BIKvz6yjVPYL5hJbFYAJtsWPCD31szR4L9InpiAaCUQj2vgLBAXDUGJX0WOx2B
XB7q1GfVDSxbpQe7G68G/qXu60+xqniHnoL8Xauf1onY3FIT8mz+shlG3BO8x+GP
05mgh3arLPyOadE392JqjQ3UrowA7APGvwjSnFY7PX7LbzOtlcfu75W9pSyFOlv6
34X1zPptiPG+edyVg5z85LswPE7DuXDZS1ocS+0vJjNcXcz4zOlMbKRdHtHWmFlM
V0mKd5+iuu4iehUIq+o7EhEutAN7GT0XgAiRRib0BD9gVfrJH6Ucr4nwFRTqpnYA
gda6AYRDanXvt6udDO9tpCPZ3kTCNgTwq4pskXgm+YJVbvDDxz920QYMAEakK5P9
BcmHv5HvF40D0wKRlg70c8Fy98WNktP4gnsWeMBENNTzamukcdX/3CNxJwzyRqNG
3NJYErR9ocWSkz5NBxA4RILDnUy/j0Zq2ujEp+24P5yo4TEjYNc90LtlO472aRLo
iT9ezUOtr6EWmixVvqSmNAh7YN6+9I8SIR0D/GU9+Lzr8i3Z6Nin7liBdjb5QTKH
kvFOymhXNsUDeyA62lrtVZBCNoLl/uBqH/4NWkS1ANVZa8dk8Vp72ygLQtBbdEIQ
FFEXjvfhgvtkbc/goiWXoBMCFXQ6YQ1Sy2OkWBBXKxIRknGJCLutlxQ3cRk3cskM
zKOTJdHfD0XAxM/kcHyA5iixdmpn/pDdbKk8bn3+/UzjRz8rgbnUq+Ft42pzXVed
Y01ii/FJZ3YTmeiBI/dw8D/ttTID/ff0t+aQecyydNdKsmuZlcE8RDwEo1kwnxNL
o0jczuu0jNGPzuBthVmI05s86SVz/j0yECbbhclYubS7b1aVux1Ttb8Th4kAZBFi
eiHNX1WmuLppGode67EUobeHnaLeZQuMxCRtSKG0uY33TXf5MWluxRag+wAwP01s
OR27PvufjMtGcVgMCEhcPrqDI3b8f2Gt6RN5aiYTkGni3QuMoox4UTyrnIduMQk1
4uIF1Yl9fPrQkwzpAY/zKmf0e2NQBaPpYJw8wlbI7E4AWfZ4tIMcfBGAi5Popawd
hqtv6MoqgHHMRjc29nz79T3iY/Y8FsF6L/T21x5g612pTZL/xbYX8UIbx1Pg2EiD
odjTRTemyFKOOSPZmXcpFgUa1nu8sDQ5t+I8CYdAPNqEimd9emfGh8i9uYP7Eb6M
2lLcZOHmiIpk2pmlG8pJaBDWHB3VWWRyibex0liP+mjnU8DSSe7JOlNCR8Dm0uKO
2xD3+pNquy5Xup0/7/v8vuBP7t8d+0798jKAjMZzYksTVmbgnAQKqCiE3DeoQzCJ
mMnDcBMJTjPEhsgxDHPpXM1NspQjg0jTM/91NCBOnha3ZXRMtz2YwTEU42PnMhuZ
k1H44P3mFzN0z4hjuVlO1m6jRvzaZxf1kSmI45dbXsSHJ1IF6aIzyIcWIAXEv8v3
uvQ+q/yHsAPB3nsVPAxbU2PC2yMJi96Lrlk1528SM3imoBqznQERXewbxRua/fXk
xYBPNMEL+MUSNtF3kvllUPQoJ2fhwjDhPq4ni129EWMHXTyvTcXgj8EHHD6dKiqg
yf3WFOBuzY6bfUR7OZBFMyEFYzfCyY1VG30PHvYs/6ytKDZjlh/bE8W1mPZMq/j3
kmc8hwXtjjVlsaHlEv20c4ZKIMIIzcTInvXPNegljn+2bMtY4cUUJMhNMsMJ+K/O
n+MUsPMn6Pi/pvDfYTi+0RA11Ng8n/qjTg/XvyHz3mxZKZxrws2gFGuQBUvkwP+C
tProysJ0mA2qa8fc/klxpDibBA6Dig1UN+HV39z2ThOkLvWVVX6jjMon8HKJg7Fe
USaONYSrKwm2gXKi9gjQYqYvYzL5t5I3mWUBZ8ZS//gsIGsnkHugcA5qMCRW0wRR
xFhhXuC7PPYnMlvVdMakORhrevBv7H5mQJKMvNHtaq47j0TwIg3ZknNQeQjLQPQS
zfWSCyn30A0+nGuDEcqU52NTwpqI69MiXf+aPj4OEgYFr5iAuk5kEU0pexw6wK3H
eZ3pTqdZcQCua/0aBTkSJQ5xoX5MOjOwnwkAcqRk4rHx94VqU27kXk+8rDY0nCtd
ggI4f4UvtpBCxUk2KGj+WC3srb6oK2sd9QJYWT3ReYVGcKJqqKLo6MMnpzO9BGv+
UwlaLHs5ylHJ8YOjZkKV+xgpR1S//eoN5ip3DxPzsqx2euriYKdijgLV8KKYmGZ9
fTZR/Fs/h1WbyyE7oEDNGvw1Kzxf/5s9/67XoADiTfaOdt/IuWSMdCcLi6fgDtkl
Kuv2KUD9HOPyKfaSAWZZ7pCj+zGScm3yuARDCgD04MaKbXHaBev9x9eTNLnerUYT
pD4YAfhmHythaREmwU0ARrgaam8+kmlj5quRLo4648M1jGdQ1KcmG4H6CFDiSRpl
yYxWAdWMw0d7CSFT3O6iWhyvxfl6eXDDfdsUCbFiHGvQ92ZO7iklJF6q1Hkz1LBk
bbqsR2Lc65B8Nw/m5DBQIaqdKTQhE7btAaw96iDHkfEAb1fbxSZ7ZIlK/dcL0IfH
kcXfdnWWPclrKILlQMZtwBB+hlvsKI0mXg74cO7bQc0mbQPIMWdLSC/N55Fn9GKU
Yv6LeRa9UfCXEp/7JWSh9vhsUFtzAhmM2iBMgSr7xMvMfkyxZa8yzBrFHl3SBA+O
R39FCbzf7Yp7OLm3BzFsWIpK7KBoo8I+N9YFV/ksEcLLEkyxdPOb9eM8V8NHEhli
ZtwZdpasQkEBW9AnIaXx3RaejVJ11PY1Uvexb9YZkElq5MXpDT+rmFXNXRfgfYl0
4mkEDYmSYEcDv5F+oBsP7A0Utcjpos+FH+zdq6ocJCuJTrX9xbQzQ7KXRnF+WuzM
TrZjxv5uoT+/ReoXajDOeNl6mP5SgWom156bp+zhv55DMO0+8YHsD3EfXLqFtM4S
xJaptpeYSJDb/2ssQcqr/o9o44WmImtBfPly1QtJLeYkSUimOlyZQUVq7l1+LYQt
rFL9URiMtaQ3vFoeLsuxjM5UtzSkSI4ee/ftp3WS3FuOz+MR/Xo8WOLJDuQdftIX
75BDHCjVcVDHlzBpktBgWPXG08dofYU3WZjlnX5owWvz5OEvAEBkPCbLjt/J4hE2
Fa/CRdVRueIIZ64CmzCJDcTbSwDRi2oiuBMdcpsilptnWP0z7AF99lMHFS+y3pQN
/Gn8B4lc+QkIBxO8lTA1ebGCDUP7duyFMM9tvLN/LftoTao1IHkvb7w6D9ds+Q+0
CGOLahAj91P61tYasETKPYHvwu+Idy3AEQZYUUWETjTWGhyoEC3iOMccrzbm+S1E
CjgqRtz2te5IkVdRsaZUUMit7Gx/GkW3D9MgFSmqRUwNgy8BUdZTi0JAFIvN+0qX
3G1y8S72RWUK+Vgn4LaG0HbgXqh3Nb8rEDf+WgNUkI60Ifh1nAOO8WCwy+cHmWUk
1WIzi89f6enTIIy0INkgtXZfZZcxpVp8b8/jnwVqmDbg5HTzipF49ZXSUS4e06to
RP+jUh8HotAzUL6n3ojby6krKS2ct8XwaRIPjVJqWGKHdiiMCl0qISMbpgJINSEF
UG19ILezkVHlHYsqWJU7tjjCx45Yic9bVxaML/QNTqGiYU0oQyH0DSScuFzecdu+
OYmPp1KN0y7V7NmbdMnkhAg7rGmIAekHQhudiyJILnSmZUpVkKiQAYvqfvS0iffm
cN7rr3qVOIPl5BdJuqwRxVjXjWtG47lYqPzXEe1deO4UCv6Ujl99MUh14PpMB255
aYvIALF2h33Pxzi+l1ZOSqHMEvJECH/RIWIDRM25EhBhBi0oGNzJt3oUjiILdStI
Z059G1PhV5DBXjUDOdnPHl//dd762CxJb9URrDsxkfYlrcubiSjn317G2YbOlpwT
RzKOfQ3KC5qOfFubUxAXqtDJKnrpFPibtJzURN24rS8cRhs+ASNy+oSKhXxBD6Wq
T9rsviGF+MrzIawmfkbxHebuJljZBG59R/a/kXHUwfMeIkSlRU4xaD0mGr3l/Zur
GaN1o/R1gbH1MVWeByMxSUnYYf8gVfGeeAiyTuFo/rn6whWpwoODf5bNNp3Zn9aI
Tt/MvPfDKDhU6oO5VQwpIrVtnz0Qcjhj2fF0dEGxGi+WpinStBPjqB0LLlC/eeS7
eA4oJgaeFipmEUBYE7DbY//TiHMgyoKMUla7zudrlEH6Jgr2jyHRw059+4kD+dtD
pcwBfK6HW5j7osCt+1S7GgRW9SbuSlIZahGEdICWaOA3DsTtCovvrp95vjjwWxj1
AlNubKWaKEHYWP6g52qlZBesuYAAoXzh3Jrv7CkDrzw+H0s7VWMGvp/y1jtQPFjf
w1fULvWpSC61GBXeDZMdBA0tU8H8U2e1zs5KgmOHb5X/RIuDTCZXldSCIUP/B+Va
97RCgW0IiKZ19HzFVRbSAq8d1Q5paqikvsiw6tygbdL8ngdzdawmB24QjfRjTDPI
CzM6vejRWxKl8c4GoKMdw+VMczaY1DFawjUxuzElzi4Wbuh8p+9HSd2noiRjAByD
oCCIcZ3nYj/WFEydaQbuWrQyDaCotz3bjk92dg6oDLCVzMQ//9lVfURW72x85cZp
EdOQ27AguXzcQ2gTn9eIYP1PeMSP7wk5lkHcL7RE/orTdoh6WVMgqW9UYA/dznb1
JDwXOV5HYwy7h1zpFYhlBIn8/dfWkaZxeYeEHLAev08sfENZnG2NjFW3rdZAoJY0
q7E2jbhwl+ahsZqxGjuwkq4JZjklAMqcwReU8JqvAjANoTVEu+cvgnflfDGN93DC
wqPjSJsbKGb4b9+NIt/oIadpkgZyLz3OSnWcWHAY+MBYReZADEozf7WYrjgWa0i2
nTucqD5XkOrjKngGIzqo2EOYIZIlmI4RMrLd0PZZzn0k7lajo5kBB/qhojPgQ0km
IN/zwx5Z96VZiWzqViDeKoVbp7k7TNj1osz2hXzSiZFEL1kMiA1L4HFJO2OCeu12
1a2DznbtplokndOCD3yZUb+1xjz06ontgV0P2JWySpinEPgbsY5C3YpWe9fYdCfm
buEUjxATQ9d7jsIwh7u7XKKDQVHfipNmwZ/BG6yqnlS3huBtXI+scIgyxqRJzqwi
bSZE0rblMm+2oadvpsmIcNBkfZsqBncuWhc2lEF0vEh8vGqXKJIltg6nJ5zBCgMv
CX4XhZCam8KpuZF8m+6KrRZT5h8oClxGWombwzIaHzrkX8NQlXTX+OkEhzZZ5pGj
/8ElMpX5DJH6u3iI9atcUiQYhScUGmsPs42DZsEf/wyC+3Arhg6lTSTrxaJ9jW9E
ou+QZtu6qZ2TlZvcuq7xv4tN08/SfK4n3gzIov9CekcyXK6eh0z/v2N59nSxG2SY
nOu7Lh0XOP3C8bmalUhFdMDjUvleB5Rn/5a3vkOglS06ghoq/Kmc1ugm/qApxz4v
/cm5p9FNUyRS484ocHuoZ8a55WYp7s1TXTmrvSOQuQ7fEOsM8MFu/fARKFlT9c6w
OenZGY1JMDfNeiiVPuMOnU/cCoEK29Bacb3IcJhIG9SHek6sdmnCvTo+/S/ouYJi
Md8oxqJvLc5zWS+wGUviY9mbptV420OVa5l+XtpxbTWlQvlUJpalr51yWefNryNw
0xx6Q1urCbsG1AR+3GCdqz1g5Kpx9SBq6EE6iQDEk2rLqIGdwHfsl93D98Z5rdUE
vleN1LgD9DiNvbUxLptwxdBC1iaMMg5y2ArpELi8QnC2HvmlSC3nEpRuJaJV+H1A
B2p5xZ6AQtEGZPJlzWlwvVGMG/hbw9awmTMDDR3ZW+xChstHKRE9BnHtAM54ZjyH
mCp8X9C9VgY/F6flbAYFYFXBCSndF9AIkyuQrGs4PVOxYl+dSn3Ickl97Mo29aPP
f/9g2l0dEBtzvghCEAlVO9SOj5GKzb/R3nvjS2rMlWqRODbm+LFh4Kw9/SeY0wGx
R1cjTEmmYYl5iWsFbhdJpbDq4jPDfNxtlnZwBN2YitsQGDP4ybZrKlZeIPnOLsPE
lZzXmhHqjZLtzYkRHZqnJz4GDxM1lAD/52I2oJTmn7pDg3DKtcZ1BME9Ruk6QR7o
2uDa8UAYUftgQTdGlJJMlSBgj5/EuSVaOMWcCFhtX4FHS8mr/BiuKVBwIY8hdulR
GFT56jpNXG6Go+v/Lhz9m/LDWbsCuNzw5Qv5U9jpUzUMiU4lL6u/s83bMn0/uwVH
ybeMOVEpMdcynh15bF+39xX6Dgy4v4AEd32Su8xko6XRuhVi1NEL5CmxnvoWrvy6
8Fhswt/Mqh7SllRe6Mr7mqCY7SXN7hHtdkINrq651t5MTh6odELoKC76iI3kRN44
QHRoJVrDygzFkbVgx1TTujqVqGvZ5JbS8Zrctg26SqAEGcGEJdFUU+WmuJsdi0FB
jztd5yDiMKdhvsQDYtD5kulMW/D/QJlTbk1mb7QtFhuWFaeoCyRKnJ1dq77+E3/1
iJZ/K6q+WL5+GUGOXmxQ+rVFRB6cvOWSF456h6tTZQFA3RX0EHQ7oLjZFPloY9zt
qxE2l8MQs4T6Rq+fyTenJVA5tSkECUy6bqPiYUVKK2GZwH12Op1/ynVkfLWSfUpR
HBF7kBfUNtsq29431oBHZSxXyGD9UNvPmrs8fabYxs5C2DO7yG+WeELw1yksO1Um
JuuIotxnWHWgNX/OY7z8RP+zntzpNjSCbKhdxndiQ25nMinsDjUYDimJutNpc2zs
Br8GaitwrjlfqCwNTMXuu8PfGRr420baDOcIEaOnfKBCqMNJ7sf97QKOQoipsXZH
4wwNggx/EovEByxhoNOWiWyA8mEaoTp7WkHzhG+lnoWVdFhIV9S6WQrQSK30hEJr
VGci7/EYV6ih84dDNCCO5/eFCMo9FMaq4mySrQbC6czCxoCFQ9lyoaucCIIR3LCl
EiVsWhjQr0gyQ4G+g1zRgjNTNb0ydvhpJJPmAw91NDbvP+b3MyiyP/Yirj3OHDna
1oSZUgTLBnmYZ9P0yzhAo4F3FTG3l6QkXWTs776VxrotEXjUXR2EBg7TRo/ZpcyO
ujyBlBZEYzIKiHJTQS1dfJxZ0Rcrxi8s7KBL3jUbKsTtUam/uvVkWpctwqYd+9kD
MP0eTDm1BA/PkU6Uvr4acJiIQGRfN503S0/73DiuJtrmJ+VUXMQrPiynS7ALYedU
864xPVSVX49ykvuoKH0gU27bWdi6lQbTMBgDZBMxYMaFAb6bFshslF16KrjNgtkr
7ZTOEasB3r9BobcC0yCdK/TXqfb7Mq4lu9J9WLtBVeILZcdzKt5BVYwiZLxiTY2R
T43HLIJRngH93Pv4ywBfK0YwKF4YT9CyCV5VMcMG9H9S8D9IW+WJipRd9eI764v9
+Tpg+DvDxBzZfZZm3EmTOGGB03YBShOKSpoM9jCIwgw=
`protect END_PROTECTED
