`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jp+I9pZvsWGXUL1hBfpDyz/3rqx95wo6s7spqLnyIXWGwg2xR6e2vjY3EHmD+sxS
hDqeWsMqSrPsfoMWB4GUYMA8KcBBpqOj9nOAQObf1E+uw9npnIyVUsJ6DU9dM7Jf
pSx2mhosghiYyozEExTfmggsDWzgEkJ+phf7ya3nHMwQhn8Iym8bw3kS/PgTLMfb
HGKa9YH4eyRJximDoGnEGESxOI/K/xFTvKMGHa+Q7ExSj8ezua1m3zmluXyaSfxq
5q8P113nRr85nfTb2DdwKMkaelSln6pA2us21C/PSBoKwFkh+sru2Jg+FgBg7Fuy
7CVJeCquLnDGouwFzgSEsSdHzIjnulFnQ9URBuCpFOtavgTbfEKZx14GW+ywaTD2
xyCZucHJlBFMnFGB2bJo0jzxGufe0C+C0de7yVMTkSxccsz2Ic1sE4Jz40mkYgPW
wYxz8gTaYYFmLUNL0u07M6aCM9CGz99nJdmNkDHiR15ZPXZeDQYxyro0zsBl4IYZ
47hr5CDJosKGSfj6JY9ajo4MhkBPQuy3gQBLW0rOknt7xEIQGuJ8cmeGusLXP68P
VZJbl0rQECKuQgShKAV5j+g/vbp7Dohe4O7KoxRNwqY+ZPm1aUNdrYukCzpiyAnQ
jgh4jAgOCXi0rS+nGCqB9M6bOQMXuoXtLs/ku084KsQ/FTtvdvnOtACBfvWNX36a
b9MojssHiInk25Lo2xbyIZyD+BleOebFzhCY2ktPYEjx8bgxahzyE7vEuG64FHn9
YkeRfLQHC6v1EG0Lo8hw+3Sz4xmzkT9YmFMdbSmXWQyaMBmp1ZNvHEk2Og8++J7Y
8hMReDIa4kzKf15tP4itUp2tQsQg621tqd+tH7Q0FuVIjgCqwXz90TAvk10sn1Zj
r4Ct2Z6hhTaskL7LYBtLMEPmBOQahP39SOA1WOqjhQkxE7M95NYD8YggV6rJ11uC
PgLV12+VH7RMZVNV3fYIC1aGmb+8K9WOoK3WfGucJTTCCogCgzcoxtccpI0wUUT1
T46A+e5QdPXPZHevFSwq/CLTOb9Aj56sTKvdGO6/ifVihkZ5Yk5hDnF8uydKc40p
`protect END_PROTECTED
