`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEK0IqH/ZDN93QWhCOLXgkAkl0mLTwJm2+Ztic7+a0x2W7pa3GAK/Oq8ylubO+v4
DB6knzBMR/F6EHI0W6tzvLhuY/pAdlHcx9D1sGcZoH61ooEpboauw5QJgViOYbFn
Wc3PQ9NUnCI4Hii2qky0ABCpNPy68e/ZgXbTECId7al7p/3t4Wm3S2h0mUzYFnfO
5YtSW910UNNjExQvztNee3vj2Z/FBuUSVwWhNOdzNZXLVkwEVLB+hLXDmt4OvPq8
g7rp7EdGMayW2VTwnfA3qwUJpx+qnB2uk4Z0ZVDqL/lER/KmYmeLSQkVDuxmF3KC
4PnAXkDz+qAG1gDim7qvtZB0nJ8CncSWhzMSI755OL1vH/CBwbUJOR/kuasmv0JF
7i3YjguS0/uwJRoYdkyX9xRABZqFDL8NDPgcA3BToFMPtznIbR1IVEgNvkQsJJ1r
Cmr52Hc88iQx9Xtt9W3wtsyw524p3DQ88O4qKhUmRKAjeN4PuX5DKFC0dRTYBd3o
rZOsWzi8FXmobgoqUdvjEuGEjKEthiZu6UU8NXUNPCecVhcXrIZ8EHIojejA6fgM
G2NIPB8MKDVvrS/+BfME2ZhdM8gsaa74sse/NshH5mOo6CRGr1OXpxcEiZmEP5YA
uO6mAyKjlh4ASTxNgddXISUvoqFVJRwmhQ7f/ZJZ7o3/00iEwp+LzVlQsE5ytsLc
ZiMJO/x5z5OC9ERuqjzG7KWSdoAcG0M0enqrapm9AdZ3Z+t5VrwMmpVXET6U/uI1
wCvpG1jQcjM1UqdDgmBDFnJHIL012Alp7kn70ogvWCm+DsiWBzXrLffn37bxQxOy
lYJ2h7uYMjx2iYH62bw2IGqPdLUu06ztqIT4p+VlnxOjj79hDfSRH8T8yJN9a9yy
18XgkCtFDqJKJg1WlvpMKuSVqiEjibbyWLakgUhysA/JjTpkP6Ul3EpU3g0f532O
wFvwpdgjlMirSttx9EHUjB6PTxGU8zZmSsti8qa3F7pHtxbDY64BNGt6e+a+WHpW
UAAteXuP+dYIfeldF0iVBFJxh8wXAlCLDT5P0kMu1TxqIhevTcRXxCky8d9yESQX
fXTCbMeh7gKt/G+uHQutTpHX+qvDWihIGJV0xkPtNc10Pxrz4IwHTEKhcP3UoX3v
ngN/S4TweWwh/AOshysFillo2feYQ1SAzw3zTobo4weDUfEIoCYcm9iYTgFJhEJa
df/p0nn2hL37iSC6y7lse6aOOC22gMk6GeuMo+3mUp3jLc6x4aRJnl6uCmyXnQDv
qipLf4Kp8OFuRT6p1hdrHW2am+l/tl4awg+86ubTRzhoa94gwC1qGepN444rApau
jeWFdnf3LL1ycumgn5jKECDqhy1F/3BnNwB5epC6g1DV9Ch9bhsb7Q2Dkz7hFikA
NEi3AtDE3sestvYZUqTmK1PHc1ZgEPiG0MA2H3qf/DCOZ+CxwJR9YMA6QMD3/8sC
cg0jWafCtNcWbZ5QyNZnq4utGZvDpoczbkazfLcTJrsOr5yvNxocG4cxxdE3xcXn
Ti0bUXxLPLO38rcsbP8VTn9EVHeMxajrCmNvlSC1whczWrletpH87ON+K/RBqUHf
qwy0lRO1059P3e/iuiqzB0dA8AZ1AUSWo7ON6RaFKEMqWA09myfyQP/2FHpM49rE
vqIz6YHkGIHpgtbZppKPsXXRPW946I/k0z0EbXOTtB5129DgJuW8dfMYVukyEukx
5kHWZ2QhX0IAHj+w+YtZdrO8TffaAg0SVAPzYYKfc0PvoKwth+RwFAg0x23NZtsG
qRAOYPQAiKPusc1dZOe9WVUJh7XokSLnAzmrVQ3T68PT+J0jUHfZKYsbInUV1Xdh
hecKFqWtApo+1aELRtjsWzbaX7aHaZT760HhX6hswZuPMyDKpq0ZEN7FBkrvPn0U
+nLA88QaYlc3QQqqtkKPrdCT7RFozr1xcJ46EUEjqGrZGxKq0OTHGXvXrLbDweKf
axGiM5UdbV/Gk6+wrqOvHvmGwLNhTsk7Z5YQpyxlCysHDvztyM2iyWlceflsjvir
5fl2cEzPc/FRE/9vPEGVh/NU5+/88DSh84qZ6dE97yU5T5a/zTG0UQyBfTS9UCoe
mRLOQ9X5sgztkYKYGpCigTx1Yt0V43JjijGdNiapLi3TCuiM3836eHyh9YWfC8Jm
qA5IHQ7kWR3MvxLyBzF6+p3DCLcR3V9Ts2+xW8vymgZzimng66mq5UcY2+tQUXK9
Pm12EnIH4wdXDx0jx8PVbpK2dIw0qXqcCmEzsmM64IjkdQmlFXYniW6x6G8ahsmI
lJn5gVBUXiOq3GNfAwzOOt9yveyfsFi4SOG9RRvOVF1xgw42YXICI+QtN3qrvOxv
9ypRJVYfZsWqflgIQSi4DORGU31QwqxyNsJmI78UeguNZTT299ybv9hwO5L1Snd7
lkRqtD9YWHakpACiGnBcY1nVdsq5Jdl1cONBYIb4CyLU1mD1J9JMigErF6aQziuP
DgbIS9BhILHm2gy53GUuz4Z5smpr96kKm+gLDTCF2YWZM8ZJJnT1+6qTq2wGIi0v
oln8f5eXcQY4CvSYizXVV7bwYcZQXdknQf6wiOiLm2xqOOzFzp6LA9Dl2/br8Nqj
SODxKjT/yzEdmNmk/QJil8ZnbblAn8T/bWeR9+nCbrA3wfRcoA6XGsW5HUFJVVmQ
od4nHBx7vzOKH4vch2lBYgDnhYr5Tm8XfW0ZFp+edJSUiJTxX4dpAZN1Td/sgKXV
e1ndYMg9MsP9AQCLktMUgrUii3GNltmUCacqs7urGTTr+WFw/w/DX6yClMJdkYp0
kgqB5yKWx4B7R1tTCQXEUNSW0L6zCtIR8QpqvdUHAToCsef5wZDa398PrIdzEoy6
BanNUgYYvvNffxxiAS4yEabNywXjntnwSdkJrgeMZ92Qxtz8A7IY6NQn+JJ0V3fE
NlH9/YG2Pq7U7WJb0wAuksswXqXtDf5Z/tho0/GkREXYwSklnrX1hTxtTiKpgX8c
+FVRqLeww2jHf+dKBlCpntIKXTg7ZbHSOco8M9nKGWv8Q4njoYmmXf4+vfNi9F1L
/n+GT0qWZUY/xHmqnIJpUQPKQCAh/7EtAaYWVxGCnq4Cb6XUt/LvdzEJEU5Drq9J
iz+Jka3R+3t2MGiyFF0HZJ968U+GeZYYL184+tYoRRc3lF7nk8ViZdm33bFp6KqG
n5M69GPINEID0gW0sXw8+EWIg0va+G/wat5fnWwVESwyNCaM4zUiNQYPnawDy9Th
8ymUpTauwgRymhmAgaQ5vNWjC6+nDVPriaWE8F9mis+4QB3OLPKT4+lTiRFWQIgL
H8YwhOrgSks2FQxB4Y1OsxoZUhV5CBSof5SScdMecjFE9yDwRNSiI0wzyT+5nV+N
rasxFBApmFpOcxmo/jEpBMbPjbCe8g6f30YgITE1vsqIQVLU8mJZfBJ5ylZ85N1K
Lm36xqTe4yH8X1jwkJO52Z1z2uUxH/vjGXI8AOf0AopIzSbU97A0pHXNOVBzBP66
I4w5SuBhGhHWbdClwIGifm/y6u+ReeszYE7FOuFkZUYyFJ2R8cFoM8jlGyj2ENiP
9JdCsgBaApi7t91BfyH/Eb+fH9y2TAArnheTMJ6l9iW3Hjy6cTHTeWWUxTUFEDpt
GH6EHbOD1sLK8lrAQEiS8NiXJoG2TTh41MADJEuQ/HBJQqeknr/oWLexf/t2HZpF
9F7E/VFsgE6h4oZGxRG6cvi/nGjR+F7YVUk0Uzqbqv81aaL3R/+ITAx/91m1x7Qm
9uB1ZOxIrYpPbHBUzpZajs2nfOPH90UcepEPPz5nLoC62NIg3o8GrZ/HFD/OC+Uh
eKLLN69fjPJ1R7116vMpdYEzAfGtEomAOxqpBFLP3iFm+6KwxFN91zyJnwTBG8WA
cJFcYKUQ9iNDnoqSYY55wBXe8QsQ3C6kGgYfO5wlbp63wZ8UNJKTOG0S7Ju7QAE/
WHZoMxWs08379tycbOupcav3SlAvjstpdWzbpDlqR+9Uv6R0xwTUCN7R86Tv7ox7
YQU80YFNapA5JNHYM0E/v/XgutdYLjbOrVBc2FVkiZMA1IKu4xB7fbtIOhnvJfnx
e4hDQcMTyTbU8F1zIlRPo+3XxKsXyAOEKC8opee8d38axoLhAfY9dL+BLCElyTwf
usuKDjRLZ2aPa4yz/GKQtFD/Yxzk9YtZEiBvKFu2M0fth+og/1I9X3MDDXKj+UbW
DF+EUwfYgVHHdeO7Hk8wPdU1crtpoiu905VHFnYWEjtcySt2BMyKAss49t1OqDYs
+rIFgKOKVEj/Zskg5UC6/U7DGXJ4hjeG48fS01Aw2zTNKlX97Kr2WywBoTXJ4dom
jrdG15xwDxGIOxcPXjm2e11c7dey9MnF3lT4eY0njTWCo3YvW5KfSKz8A1C862IQ
+OAP/Q+RElJrlYrR38whPbYPu9A25S7Dtaxprla/mWTSBRwgXY/PjVtdokHLcG8V
+H+m/Li7gppGhR0tHh/XVOTyE7MNicLdzX+cgG/QYp/Vc4uySWVzCpBr9ApEuXzm
+DjzXDBMCq5CUquF7FmWmYwFkcbqlJYD13OYKW5J2+CoJRMNNvrb/61olAXuGFdA
4kRQVcoG/MMSjfXw8DSfmy5a2JgsFQJ3wHquO6lcz5XUmW0hVkuSa+kJGzPCbubK
EfOdIVNRefiXwOQSOgAaTfW6a5U6Zc3adN8rYEucAAaIPI6A8/UZGFGi5oV9CBt5
6zYDEouIrGNIDC7ayKAfuCq+xaH3BP3nDTn19Q5dg3BCbkihzmY1D63EFSyV/LZJ
PfImLoPy6d+Gyd28xQvh9kNOVJSaFYgr7A8yQlBkRcOb/iFii3kZ3GBEx+wgVGLO
tgkvVfGRj70xEkL5jJVKnzMTXLuzyYVAqRYFs6xBMMEa4Z24RVjofPKPXWD8V7k2
YEDb7RBYF70c5GBNVrjhbjTqJYNhbjSwXu+yIjVzVhdptkRaprGxKYaujuRd4rCW
A5+q6B9FF9hvjJ0++N2hNfv7DCl4/xK6c93rFD5VrotI2Ry5ea4vAuWbL/cgWXOS
fTt0lkdQjoH+7iuynHOojxzwGeos9Kk2Sfvdv+RlnhA+MzzIEf3h3tY5fjqiYyxy
gxrONLbekDgmdcyvUzQZp/CMOSHkSJtQpSoz5YtEQeCjawhXlhPxA+TWq6zeRsJ6
VrREm2x64p6kNbNdf21s3bqPljHuP5ssjTTiIvksGLJDxtqKisNS2FUH4sqTHC0T
5FpAxT1H72M+gFA6fV/CHddNKDE7EXdiOaYXCEPA9+mm4RovKi42xSom5eBBIlcq
A1o9OfnXbGfI8yVYli0utCPJ3kB2hpbIVxWZ9XsuEWfHWeXaQ59bQ9TFuqWaJwSS
P5OavoIMzRSFXedgQKf6DC0K1OO8TJMDBo7IAlRdMW/rrOgB3iSDUgu2cBGJX+nD
gkVtemSIEeKbjFTQIQFygMdJ2BBOr5MEogd4W9j9kGBAPp5YMtnhIw0tXxUMwSNN
YZLF4jt+Qox6D9ylTX9BnvENQhpH/SvETOk8/IlngU/pRiHljeRNs+vxsPSQu0d3
SA7DolVa2olUF6EJBihejfMDgUt5NTAOaEO5B0cuYcbWYeTalJm1FGF5qjUth3BP
+Hm+4oJxGglbo4FWH5unmrLsyGxkAhrUHFrzq3fjJIYiQLlCy7piSq4Gx1cEKMjG
b88LtcjQZRY2w42OYbkxiB8B+TCvkmeR5kB0upfPMjU3SzpI/Q+LdPov/4zU33OO
rLJlx2Hq/WXI3oVU3UFxAm1TfXMcF/7FKixZ8WOdoSGZghVZrEUeDD1YmLNP32Yv
p3o3aTMNAGsouDRVRqQkm9UAhdWqQLRgRXaZud/tqLv+8f85pDWRjJP7iPRa/O63
EEygL9MLo/Kp1eiS/AH4Xk4BFiqmlXtqhOur/WSOhfON2/EYQj+2AExRhzjJ291d
i+BI8casg7PsSVFslmJdfRuzWsPX2uPs4AKJ2tANgnFU8qXAOgl3hXpsE1R0P4Fy
kCELVsSRopVVxEUKePhE6fI35flRu5gJYwxVd1ifrDD1jT4QdMQkkPxpFIcm43xP
2TizjZTnUyuySFs3CZ4/V1oV3Gbnu2fTtFSNHUDOz/WMGUvI6EerX34zVT2RTyQQ
mVnz36GYiftUHA6/zSQtp1NnvnFn+kSiEMAu6SgMrm21e49PbllS8TUgetlTXlWg
mmLBPYytVYml/bF7bCglD8Qri9Y1yA7Mwk/kqiwu2XKcTb8YA3xIniXmthKkjrJs
MPp3mZ3EdOs5/Jpkai6pRruKyQzIAoAPiLkgf7qptOILdlD8Ov20DRpLoROd2h9C
4iXj+v0w4Rwu6yvMCOTlVC0yX/tCJNk9kRVezJsMElnu2K5x8DmUnfh5w59ZRxbI
v/RzyRU4GWSqMYPYQ5zds5NohR7phZ1a+dIyBU5DYXLCRV+ChEd0pMRrJJieiMI+
TdoNgkQD9V7vOxTQC7kUYcOJw85NFv0tzp5eQq1/y40QGmtFXdgyLO+m01Fl5uB5
0ZIR8/WSo5oJtKeVY/O6MjD32GFvUdO+71WSFOg4HZQVy7QGRKpMmJgAdBxACbY6
RgYz4wKxyA1QC9VBG2wzYjQrf3otl+/ovc6f1jh5AMCV5KVk2NExk9f3POJ0qv9z
gfss1TscdKTgsWIIXGYsW7zxgMlivR/q45PvFuZr1VVNtzIBn4HBM/R0CfLRSyvB
A825QiucFWguy8EV/GvoAw==
`protect END_PROTECTED
