`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q40/81gqN2Bc9kiToLdrYFYJAUY/Ct4ZsTQeDV/aIkstsfr2Yb2/8VZLLc2br+va
5p7zfUstA2F2QXUwj7dqTziLUmWD9ce7pWGmWziW/N1NKcRFYho5PyaHDO9fH/mv
ZTZZM9cCKRKeqsCrzXHeTzXF9O2wW95YcDPAkkCGY6n1WktdmDxyeuUjSPoK0g4c
JQDBkcv20uk0S75CsOf/cddu5OEhNGMcE+ors7/xf44Ey/ZYnJ0g3F1WBEvi1XZj
hWk5LHs4JRsh2Z6LWrgUvrghD0zKCJzDeTwY0HatAGvcAw5dNEq4juyImy//D17i
ZH/F4RFajE4sJiWEwpvFsk3pf8EWZ8NCtnhQxqanYuoz6jeS38RK2q4r3lhMFPNX
Kqk5rbNopjYtyzWuXd22KKrMVwfHIgDoUlhIPtRs11UgkcFAT6jaYcK6Qrm7q7JY
x+REDxw6YTCmTzPjv8srqDD6z2/zMSdvZbvWtV48nAW7MmOrirlF//3F97UsV72f
/gxIZehZ8rTlRbYhSPjngqxAUSL8VdFMuVnBHALi+xKcw53lRiRVUXN7eYDzUU2U
mdKv78PHMcZ8tS6vnflLv1S4Ygt1z9lXb7F34cHjFm4CzyactJ/qjREG8pr8dQZS
9PCBtNQE5K/ma+Dlu7OZk/2WQBOMXtGAynJzETabHdjKDykJrMb9ywfhg+/+8SnU
khjWqLpleYMoMVLnGORqRYwddgRPoq6JKuFyeZWvvoC5dw1KVMdF/XEdNwnpvP4N
N9Sp/OlwNp0WR0w0tsmzAZ+l63WK0U+6y6S6bsj1JCFrH6/KiyP5KrN/u1h4aYV2
XmMAYeneoWyH+IAz4h57QjXmUPndR37vY/XVsi7w+yEpGh94gCBWeoHOBwrst0t1
uCqBEQTi1Bk1AD2yiv8hB1sIZx+SC0/C9284AJh0wNfkPJgBK07uY/9nVDbay1y/
U4/OJL/4WiWHXGvD3qZuQ8IYd8kfwDQsVGoXXRy69usNHjE5FTS5K/bmOm3KyxX5
Lrn+fvUd8+nVjai06E0Ph87AOH24d1gc6MVHlLI2fEFe7wNu4zeehEkdwAHr+rW7
q/Wk+vXFDIaknWQJNXpzoK1I0ObvTF+qH5DsoSAZzn0C9F+UzOIRrZ+2UuBlEsqk
tRzTTbA87akrChlFd0maT5xwEruEk8aDa59lOF0ttmqOf6vgaQjJc2zpBvOeMh20
Na21dQq9c8sc18DemQpEJG5RPKyhw+iv/RlBGOoMxWdtbP8+zIGmXOxFvRUlK6Bm
iO6dsawImH//joevYiKWJaLHoSMSYn/j5lzAmRFE1wN9o6lL/HlRTBRp6L1oL1eU
MEgw2K3jIe95Aa5626RUGSBJQ8CCHGRP1PAs1fS2kosB29iCSULUh2shVJ9EGzwU
DGQgBFjACXcumSetZZBB7xsLUtNuJJ971ipHYa/N68uV3WbxSSODmeQmTmmKtiLT
zBM4fRdE1P8fKsGHxN+Mim4hL7G2LAtGb97bxlqLK4O3Sk1t7n6SIWNNgRlV5NHB
fcTzChQKu+Kcgv3kdy25KtnBnG7RrbYeThMGPFGR3cpdVV4ziSvBq1LZ7qY/WfOf
vEebC64YRgDA2EvGV7/slUr+qLiQW0CGnQo5ddlclTqFbOj1MuTLSvJiklgE9Ghj
MIgfAk+evxhvg2tqN06FwqyqQx+6QDV6BzQRPb8UnSj1Wj8sCSyLBHlT3Tz2VEOw
I+xWFNOjaWz0Bhq0iZ36gNTXboiXMgAM159jv3RQmt+Dgs7vJbwEtpEB1znJ2Zr/
PCNNLYHvAN51/yd5YABU0r6XNrh85tnQwnWOddSYGDH8N2b3izBN25uCKrghwcNW
C4Ilp356eOUxMkD02zdbPinxuzgyJGxwjJR8bdBVtWw9gOyLu0uh4N7qUqRuhCOP
A3AO/E8U6PNDN9fXfveRRnS9aaq0MZYWEhRsBeAs6qnehqxypAzZXxhoGI89Tjc7
QAov9yqY50gISCpycv5n6NtZ1rA5OTdxgjiFFs+3FyPD/7CrYLAEgQ0UIP2xwbrl
JCcl9ld7yS7oZS1Zez3CpzB16szkkIkaJVOuetSBarwTIjSgtgtcyNicGiIyzGJs
wynup83m4Oky8lfN1rxnL4XkpnRwrTQbS5JccSErSjSPcWIfkI6AxD2OpjA2FKzq
ep8u8OMBn/AL1ngnTWyKzjg8Nq3ALPGABIQ7JP1um06Mu+Juhxhy5t8BLdkHmobM
oyg2mnUCMRJGyOqkLgeumQIOra3cKPnekKrxV9G+3TXRbcyahYPf4fPLzCkOfNdw
LGgWNcOsITUk5+SMf6zxbE9TXe+v55uoUK5im3XvmxmutYENvYmDkCFn9WB/CtaG
Lis1HrvFFPIKZii7Yv7kw41yGVyc2ABWQRom85qb+SzUyz9PypJ1S67SyP1M16Fl
UUkGarjVN7odeLYoP+K3gGwEfpBDHATQDRlKYkVRaCwr7o3vSYQYNqR2+u3oDQPJ
hz7k/IBj+Z3Tch/wRupDweVzc2YWhKHcKBQj34fH9TEXpROpxDtnWAV+a+XLUkGu
qY4oJ+iq4Ec/ux2DWTpL1GN4KN4J4ACQCaHC14w2Y6f4dgELtM3b4aQ3lQTCP0iv
QAKmccHvEookhvWwjX89NHUrPiFEsp0v76DCP7khizy40XvQb4SgHrsbOn7qtNe2
eFxQTBrcV00DlF16j0oinsnrUHnSvC/AC3Af7K+cUs3M7/JPoxyqc1QR5DGfab7K
H1fPLU/FpHffNkBwQdyI0muF4vBp9WPWLv0IAsYBYfdV05PI6eZO+ln7uQdCSy7f
SGRUdLBChVNpws2sreMa4IeY49bonxoUI2uKQuuqSWiFmY5rrnmXn89W/F/Ccjmv
CjAQBJzwkKaLM3LRgjQ3/jAIGt9qJAPAbc79B8yc7eM=
`protect END_PROTECTED
