`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQEUp17buQrbO14wgpVxzdrSaZJhwnoP+2edUGoLeObt+mymepCL5Zx5PZgB38Ns
1faeib7txtZDkXRankuGKgTFlNuYIBTaixzhfpuZ+0y45lLjKSOg/4tDEWCfqbSb
Ut/dhNzcuybEWpiQ82eSI7bkK0IqwtRNk9pRJGmXOh8JTY3JbrqEozzcrYHIhQNb
g/B4LclkUStBtHgeek0OLBNrXbwdsjIRxjWv3pjKuDTGcZzXrllAE9c0sdiRzNLu
tExzfbNieL88NftNCO3IBKK1SWane3sulVre550XMbovYVUiCoEj0tOD/4RqmIIV
SLpXcTJlluoOHi6VwSNEFYP4Fr1VZJvlGSzpt6bRzDI8QRWV2bN+gii18YB1HQL+
FyLnl4ABAYHyiB5ooou3k1d0XpgHt6pDRcaYvdy+D93gtW8ixV++ZxE/jbzkpDjf
QT0dxutbC9Fm3hr6W7352YYlqn6QSQvzbFVXCQLdG508ueZ0YdXZXqBx+5imIA9B
Kgn7oibj9odv4QqyM+EbUTKbVgf0A82vd1eHMFDzBQD1McfgsJazLN8K+aPHzIYT
+CY61B3Hvj+XzHbJ9raf9JzSg3GM9PGayEJ4BFj+3RvJodllQUrndZeAphgzmuKI
PDOQXUeCJuzi07qrBkrctu/u0Qeuerp9BGEg64ZMa9iCnWO+5n+p7c3tZrjURBtX
NaDw5sV5MThoLxEUwPHdO03xwyBbdCadGOrU/Ljot8+IbMp16ywASNFl/4w+rvF4
21vzqR1us9olBra8KAe1UcnL8FLb0Pyh+u8rgjLvg/694s6r6fa7RPqX13sV9Rhw
42R4kBjHIJyAW9OFWqglH4OeYgG9N9gJF5vPRtwIWi3qFlulI+ePE3p5BhD38HiP
p2nCIdUTsJtjE6ruqWbQnOTVR+QpjoTP/HbHoyQbkyCSczBAoR2V21V+8S+2/xXM
qdMN4Mc/2iDXl9P7Xmlg4Nk9kdEUli/OUf2Dd7oBAuC6CDBUpZnsDHcb79ac4P/L
7pd7XAf1zPgoBje9axFg7EPeIZsiInW6cecSA0kijOK63pnJHxbxHqZxqqYeW1Vh
1x9FgLHNi0fK3HLXSAiWzoEVqxjx84A3A8ThodL7OhubhDHiBI2QKWS5/Z8Muqch
LgbJIBJTDgXQYedS+rjSmZURk9F2HnEQR7zsLA8jpiDenv5bHYZ2tzM9NPONwvbV
rMj4hD2rTUHv6kFhPGPqWoanVqsrRtJ6n/0USaTdvzLTIZDl44BcImgK0MhamnG6
bvKDDVVl07jZE4E1VZDKqWI9TgIOYEQTGzmD99QEetMfWMTgrHrUhxvlV9Q/tTOx
o2rY9KrHgGQ+yKJ9sDNvSA6sKX/0FivEC0TxzENGBdu8PnyywW6XdiQi75t+9NIJ
HIIC/xd7nPXgzyRhqSPzJFFFKertwttvAh+Q7HGgnjpVD29ZT4xeeCvlIFO+Cw3i
NfqL8dAIV5TPsOqSVMZPX4FRAUtmQke2r+jfxVThKON0HTt/29yEXktFIOqYhvzD
oXfhYB2dQKeNE0q0CMw5VlqnoHr49iH7t0+OKWMuEq6vrE4Kg7CBMC3AXH0z/j4Z
9RjGHZ8QBPO3PxKr0rgfNFfUWHQjhRO2vCyNAgkEfZ5cygzzl4pT4BNFJCfhnAPo
6QgCaLMJ6roDy7jxJNvLCeAY5vmCR/aprLJdmlpqFpcD0lLtKoBqSC4q2Q0Tazwx
VDCOppYt758pjZXnqwV5FjYGUdXYGYTKsKqoQH2OoMqXpKF+cbaoA+u0gTn8uC9p
07u8hzkWKD+U6pq0Kjo6B9+mnb5Tn27ahtXBx6lbfyqFfKLFIwyT9QB2Tq6S+NLt
SiPdIgvNjypTroCzFXty63K0Izlx9fd18jjpvfff9mD0pFs3yLKkqBh1YWxuN7lX
C+Pi7whGviZNwVzcOUZMwaPJx+1ia3Bvev3fXSgJkKalzDVGpN236Cp8LLQQEnae
+X1bSXVwS3r4s5nCxo4cDQEDTAAB04/9SlQLA/xpgWRlHymbQSdoDTy0DEr6E4/F
pcclodUsQEshbWHKmdid3qfKQ53S/CAadhphElgBvUGpap3RwXnu28eYlfm/DUBc
0Wok8k7Uy5YAJZR0xaPkIoC0+aV3UI8Yw1VhBhgTe4JVsnwwmeujxAY5hkRGqF9s
aNlYIad2/YUUQIJY5FXvH7F1Tei+I5xid119nNSDZRwf2ITiswOw5lJ24qyJLzjN
gCgOK8qhSvkPJra6celZVGmEU7m/K4Gcasv+2/WwJlQhWCFFT1LLn+bI54E5OJq4
Y7LpveRDRwQFvzcFFv4YmpCqOv9P5I/Hf8mcgoDHRykjt1lh3wKsDM0sDh6xTkbE
y86AvPYQmRzrXWBr/x2a1JoYZo1Tts16HMUnBzzRrTdRIoeBp75m2908uCI1OTbm
7lDfkrwTT4jW06PbcAOTwNfZQChU8gP8nUjLGK5KbrhgH5ZyTLIV/RTs3rlwgWB0
C+9AtmvRsdLAfTwkxYQvlgxyelCNxDca2BNUB1kPG6Ur/gagWUtkyCwJG/2/4I+0
MA66qt+j+oqzou4d3tKMr0sMHLnNWdqkbyHBOZkUr4z/YEj871NEAzZhbZp1yTMT
7oDHYz8Qzn61zt2DXFThbED6qzpGyUFadKjUeEEXvWFYWGAIERyam5C9UqCTUL9+
KOsB6KJTb4lj9yyfDVwhBio4yaRc+hXh5h7M0bIzhIhQbGJA/VZaIS1ChTiASmOp
VoMmK5CjSNXIrPzyRmyLGkerkoTbE+cbxVTFQ+fueRAgvlli/x1MsjaS3BYap2q2
w3JliSTheuh5/n3wS1tVp6QBfO57UqIiA0byRD4nAYHRI6sfGZlUxUtal3ItSrVJ
BAMhAyUrOoWG9WMF7GHorBiYutKjSIB7B5BHbGUIf2XTN4fDaiKjMYwyJiFOz+e+
xVP7jd3Rcw/7tvi1hmnNywBplVANjQvIx3kvag1OWgigt3tb5p0tgajzNSuUuGb7
yypPyMQ6jEhU0nN2aB9J2O34Rrj59YECBFxp0kk0NrvU1oz1Xel8MTQISgNTEvjw
rtbexHD5ZVZvEIvj/T1LSU75M1wJR7nR48XvwWcjg6x1eAmr6RB59tOB1kmu8ZLB
+zOotgkiekzJRrfCi+6ay98hK5Xy2dAjx8VUAkEpzlK45vijBgkBZ0oTME6qXqNt
d6ZC/0Z48BkeV/6qDaPcugOh28OcinH/ZHow/uyz7C3SQ0cPAuNcyGXtLQBOHvE1
45v4p2bYpoP4OUnYjXLZsbTfAXmrri324NPNUioEuSsIbMF+QNcTL9Bm+DHTH+AE
BkjDgrHlj3/L3Xzz8RpNgS55jbAQmPX3wwNmBEFy6MgFvPZ+hXiY2GQaPSF3cBLk
na3CebSVmhN1HKS2jTt4X+D8vFzG/fkyJ/E28thVfKxqPSFaLC3xNVm28+70EAnM
nJhe7vHq9b86BqYisy490GXl4yHzCCCTmvvLFOUX1VhTevvGRSY7mSM4xzYhlrN8
AQVQjUkezqMTDwng8VXO9VpSdCAeJ2NNkjzebFKqugTWZ3eLEjU9PwlFIkKfL1Yw
swa3DLTNpGjbtbwkKJZtBYsA4TtDz2RIJTYL9S+ja0O09wT/rRKGfffWe9bTTerM
tpxklL5bhxPpQlP1uDyChX7U2F0ZjK64w86ApbmRv3TpX5Ftq5SLMWieRh6AcZRN
en3QMKAhRigCVEiB0vvvCrevXSF8Kza5hNDG05vNllL6xhn6uoGHhdouaiUOSDA2
FEazcOKfbVBgJR3BhST0Ox5OmADv90FjzvTxM7Mgzbqmwqf2fpMXD5ACWRMRlEvv
MOZ+z+r2tAIRTBhOIDWCwcCRtftayAvbkbPz3m5SyT/MtNh+eOYzvMYyRg4yGspK
Pzm5wVjBiflqaMw599AmCEbubXMW3Qk8qBaCPAxPXaDtwJCn19NrTeO79V3Rztyw
4bWVLRwgcjPHCId6WSGLt5txkKuuYWDoIHDtPtxOpHM+QgIBumYm7nC66W2+Dy4/
TLqQFLIdLq804apL3KXhHIPDytZu9MnXCiooNEEIiuj1w9rm1DtTrVwfek+C48Lm
ZqJwgTFPPCeLwAYwsGTXHQygdcUv8GLFi5FE1TX6uaytlSqNSWKNokCuZHNOvMlx
vvQPEQvugpt/3Tyc1jKOJx544duPaseJ7qkFTnAnia6dt1B9yMsqcfLRS2Jr1szb
eN8gTkgJsyB0beQDiGxbgUgHin2IA6m2Sbn2QuFf9LzfBjJCSVHZDRd1y2bo95ZL
k7nWYe0zAuIVynrsAZsdviWGLO8tIGUCbFesS6CR6AkkniPWHFEqwGS89htq2YlE
HGB3toAU1fAWX30Ak00IaA3KdpvE0tp1al5OTJ5AVZCNxAb1hPi4NRZYGdv/yHn6
91KZq84GGXABt6vlzskMyjDACNUiZTLHUs6ZtPmb0NsV+3FhRG7Gqfon/IVsjdA2
4d6vRFnRGTnYuKBKcbfyWSLEws1X+U9+CmUe8I9dbyu0TJVaZ5GHOd2JUHIjsPyu
ZZAdAHfhSRB0bthrJNsoZbchZE78g2jnOiso89tsTk5+3YEQyySrtzTZu0ga1u+C
wBJX/2IVkratrzXyB6bva1wRS0aJf8TjR2QU6Da/b7L7rCt1IZXq07uWOQgaenoL
vFzE0gnnpu6YsIk+aCv/nMOjhD+72rrl2mFqmMpmCI9B//qnSb6FtObARXVynHyH
udv+zVbWD1UZtHoWQ5KSMfMxLPgWQhe6hWtNFyqBgDKZsRo+8v8w+Uh733cg7f0x
scxZH2z6JVqwY94F0npequdIphLX10SG/b90V9DjWXJL9cvi08erzZPmue7khmyA
6O5ocC9tzdXhvg6WzHTNHJC/h7hIR6oz/wSLMkveKj0YJumIqAY3Hznt6VNW11Ie
/67D1WtSG2zufmyBFcJg0Tj+sVqqKdpQfWq9+m6a+lxbeNKrUQEhl5umk+XdgKsc
CIwmFsVnxyMHWNgVpztS0QEUiE/peG3BOHCHRzAwuVl7El9Nq1PN2HlT8MkgC/nr
GXd6w0yc5cEG5F/ObGAjjLyYLe8GEWsWDHH4IGd3tavQfu4AuiKk3qbgzNSMO3Xk
maiWzAaltyHlIoluUldoIEumEnfglOepKlrAUzCzGDbt7Dnk2zZo8Cr1ih7lwPa4
o10lsV4Up1PuQpX3ATpSdwDxqBozInQ4eanIpHbPgl83EVaCaQ3DZwcNI/DWrv1I
05JlPbSDjC3K7St26ZHZf8XpMaGv6S2jjnq3jxIZDAJkAxMq2/JhUYY+LJssdxPD
kXB6NICLbTEyUMwobB7XUKUcRsbGe9traIQT9Czekbx4DZ65i+SCA0R3LMTXB+CF
CTqxPpOxqfw8FoEiJrsAjvcJ1uhnS+q3yxXL2jdGGJ4UoBhLdl1v/U/jjtOOc08Z
qJkVC/yY/fYQrAKGLXVvWuHDlAWlYXNIJR4vxycRuafSuhnB1ZbkxlwdXqntlyzP
4dE0FKyyCiD6V+uTsRSyrpTSAboeD/1Dh5WgC7D4XH51E2WJ41JQeECaQgTcLbvY
pJaOt+28+QeI6aIa6asOy7jdA/sh9eG+KNoDh6cOr0+/sNCorl+TILvyVqM/tthX
fGfuDzYmwotEkL6bUHCpx9uvCQRWrXp3gzDgW/An/jzTwV3l6pOjT0h28N265ukc
F56R2LcgwQXx1fvd+HCOTAJvHDouhKKmla93LAcskhz8Czq7opJvg/Zik2sAdT7A
0/5Z4uMfAZ4MA+pL+zfody4qWpuXmW4NOyamG64kpkC9NNXchqlZpL6tddpsZO+H
zLploFY9veSYerXwO+aJawzJYAguPbg5HSa514Jp4uNX8zbrZTIMm9GIZgKfw7dH
lElRNMlA9xVbcTqCdxteqb0GVkxRoPHaRFl+oZZt2PSbx5SqUthfx9dStWmS5pYO
7FQq7tUcrg49hdB+A3POe0Xtxt9HunXlJKR3VdsVOTeSRq7h3AYZ7FDXoIZ+ow//
gnP+TaDiHwyen4k9+B9jqo5O3csBXmrfkM7lcaZ0dISURnx41zooIIhFiogFp/Ao
cJpmYvaypTgz+hiD+GDF69MqBeFjuw1KBrbh2X1DS/tgOSyz08Z2jHdPyI9H/cHe
RgdReuqLz2B/WWuVpwOAymcUIuVINaJ+CHV9ea6wWDhJwSYciYfKHpfX2nez+QgQ
e5NsTW6DZQDAktalm6FM46eM92oSxxugbojtJnyR80ujxhJTUbZ8+HSEcfc4tjZ7
3nQl6vruZMOLED0so3Sdg2iw7fHxUXfFZFpSSxEUc7nWscpDl4nvd5hqIAS6Zk4a
vk8HosyHWO3NyFxh633nBtmrPYrlwpU/gevY8YF8nv1YeTh6QhYb9hMFSpx1k7Yu
uB2TLMPOj8Yk2fK7axW7XDR/w9zR2LGQq5t0VXIlT+YPwlILO3pv2gnZ+Zw6ieMg
USYeZT3aDZkQhaOK1ocGVq28IHUFqW/ILB2wra0TCp+aM7mhmg/hq1JeDHcz9Tmi
1DI7qKWDv2jMPeTscNdq1IyaFGerGotUtbKuUoINA83WUP5E619wG/VaIrlxQiau
OaIrQibyUONSfcNKfbuaR9ITn1JEqq3Wj+wseG5aE4uVg7LxvGzoCx6DnMmfrDda
1INMWpN0h4JNxjb81EQL0wTzHKtqiZ6v+a9LS856fX0NXIKgVs3sc8NCmO9JETKv
OKOhXQiaPAz6MfgcHred4Nio9Fad2dH9sKPkslk93XKvrgLIpullIiR7GUZgbKGN
tPnhBiJ/PccVPf/Pmd4gQUQ4S+YWcmrwI36M9GP3EZ3NQDrbLERKUkJTd6zd2WhH
53F2H4wQec7BinCbsvLefUuWFIOZPYZyG2tu7lQ5DKKdmahz1HvFn1RmVNyFvhSK
OQz5/o/b1fNRbM1T/HbiVsIl2sJYslUEkKvSLnuxV3dJFkMr8i1I75bpapZpaJIJ
8s/M7JMeWz/2mWxTwINPmurjN4J2oBt0zJggqkb/VosSSCf2ZXBZ18ExsgMGSKF9
vbf2f8JQDM0HhVakr0gsodTlHdViexqQrqA9WsYfT+Bf9XRdeWSOSPkMFEXJk6Ul
oV3avocTeD992Mnq0xY1oEbV0ybL/UhM7MjWAYdWl6BEFKdUGei/t3GkQl1yXya3
K4KfFzVm63fhk9gthTGUVCJW4rHmXulnL22opOfyEDDPKyMJVSTyQYtEEHDcRwVq
8i280NHUOxi/cOZWJoPqE3bNHl5ofyBWlAng6c/e2NwcxvxzLqBae3vmFt5eUn6j
IbgZnc68lRpe6oiKijxbLnnISTBMZFh2Pja7Zyz7tSl3HcBaG9zREYAkxTauJUPW
wyeezNB5aOv5Ppqh5wRSAVTkuFn6vSOE1uyjkmH1gdPp9wcSrncRLFO6s8i9Ca/4
MZx+SnhBaDb0KjlBBWQTBBe6FZtJDMVaujGcbboOBaoqiYAmiqKJfVOUN4GI4mJ6
wFnUvYfaNC3S73eLGZEnJl9j6Qx/WRRcUzuwOY+4VsQXEwDvS425Ch4xg9M3bjId
R/AEFtJCdqyVEpKY0zcAP/o833uE8BTPy0OqUtvSlltPcv51qyNzE8lpPnm1ZPRf
UXPfpM5gZoXZ7v42TlE6/ByZVqPmBx1uLfezYRDnKPy5/wjKzWKB09VQz9tgUQFX
15CYUHZQwIEzV5mv9MfqCb21fF1b4Ngg32LGJxeT7kyj05WeLZTux4P3rXEmh68Z
bNrJd8BLEWOckldtXMH7M1wRNGAoZVdKA1BA5YBktL3Dz2ZAcrKVO2TFeHJSJ3Ho
xrkQ2tBg2aKji0VxNKE2M3T3pTk3bYRkK+JWxJejns5itXu1l/650p9uyNgJ5owG
Eivo28J7VX2Hx9gvpHaZULK2SfkDez+csQfph+fszKRfcApBDwFRc1jqdH++SslL
TAudJoS+ZcKSLcxH1PkzepqSJlj4Sq9NNjOdDNsUsNt6zuEly0VMiUdYFPVLXP19
/Eha+i8ScY6TOIzgBVcvcbpUIwTN5qjJjBb+GS2pwEsXTNrcIl07OFd3yUMdlvT4
9m8vvP4G8QQqk7nQu2v/uySUvDZvhiiMMhyMRgG+B9fAdCc6YkOlktukar78+iIW
vLd+xHQvlkBcZBSx0zTFS4mZOHua8B6a8Qlt28yEU/rG65QSIgxJ8qUoMaXg2hnd
KiOJ3/GEF1DUd5UQIG3P2Dl9Nk9u80bFRJ9eGmesEWVJAqQ4ZhtyK+BCsaTVzhLC
vx8tU9qLtfAHW3D2ebQjxOQU4ww/e/hzgVqIewqSV8pILLxBbVXAF3r20MQUSP7a
z9LKQRgiN7TfExMaWk3DBaj8mL7GSr1D+ixD+sR51qARPIQdWsziNc0JCZXa/x1/
sdYII9Kxao85QK8awADfZ5+z799Sr3T5iFY8lubCqcMOlhS/7p4fy9UALqpM0UoW
P4xGebJceqqeiVKPzT4mmPkwkPOIxKkUJjJxUcYvTaMZYuub8bek2GmWx5+96165
VYkzZM3LUQWK5YoNVl2/4QRPPYSbt3ocKYeBHoPVRdLvw91CK7GacAPgtiR4BcyT
GcLxvK/KXRYcpMw5qJVHaFvTajuPFx78Ok/bcDLOgFKeLzdyCbZ6IoCwQf6br/Jd
n8Sb0pheFgur/+WLB73BasxPRDgP4sehaJUwfPWcbeS3ub/9GoY2Q4fGmFsNhYuc
BFri67+MmqZUBa/+V0o7GtZhNYzQq0GQUwccki2cXEROKAJqtxFRJY0BmUbRiOqr
YHPfh1tIS9uzhLWzaFHNleOVvYZkenBO0qilOD2KO/5Vh7wNNXjB8Jd3evfruTR3
t9DYX3xSrGhozOCK2rDNP43XCaLxj53dJrWOYkfY1qsOtDMJXVe7B4ghwwo+dXjq
M96PJWD6e7Ft6BNQjEs8PV3iXhNOGlbzT47WccX19u4D6PJspAtuy1+9fDFsUvHK
jPl64PQwwIsbObztY/zknvrreI6DtbQLlB5ciLd5XyXpS9sYnw1nw0L50Pm5PPRt
lz0vFNW3RYmIZg7N6IbL28GqgNMKHy+nHtzTxkn0sxb8339IDCNP+MWXgwOWDajK
7tMvnuKfiIkl/IqWp+mnxgh2wFH8v/nMkQBdMyobav7PB6122u2871vm60d5dDz/
iozXUGx9CgEubfTyPOF1QRNXg5tTvA9z9nhQIsqV4r+HftDyKb0JhaKAws0j3WtH
w6E2udwR+mpY9Exqb3eMj07btjkrvHyr1ZtiwnhNwTjAUuzT790ImC+mG9qYPp89
RxO0i/RdYlWiD09HAiGzn3QoSyH3JJ8CeA9belnx/5upNREchvVm/mTtnB7yu0UP
sFavQqq2gAB+N06qhfuOYTbtYeUALnbmG3qIUU3AecjM2ejauFkDU5bjkbhbEIa6
CkaMOBmuWszla24OT51KuuYQ7+6Yi2nwB2Taccdt9wQg/8Osrxn6JLI+fOZdrIlD
67oA2h3Pffc7JX18ZmkdorkAmkB3Czc+e6KeEnAMDNOVEscuxcWivmyk6hI7AXL8
VB4UmQxLmTU5bc2h0FpYCCA7hIPsrqudfJYMubDBVvhaujFvbWcVEtSiZ4E3E2l7
rh75RJ9KHWAJ5lLBwXmtQXsjKMw8+1MKKlSVSLlF4Y7vFDw0YYnKIIpTmYduU9qC
H4WU2N4U2neA1xYbdIHkK8R/sv+x+K1NA6uf94I8nQMTu0z1ozK9vwnjaMyLWQsC
3ghPlpZfCURf2HlBMkJADD0lKQ0u/ATfnxOciCvz3nWZCdqVPr+z+W8LCa+yYAgH
Sj0OsCttL5VeJvwBPYBLs32Povh+GeHjSFqEZJZE9PBeYpOHkmvb07C4MY6+CmSk
Yr1JM8a+wbI+ARhefLVNM/YJ5lrCZJp9h9b/D4Mu3ixl5IbJo1vHsmNPcaa61Ebj
nJFY6b5oZizItoqrfoB0XbFtHltr4j8Dc447dSn732JIfTMj5arrwieeIlmNTcqU
bmHmtCmy4I5BraqnCi5qHnFBGloHE24qpkj1jcHLr9bnzVTf5QFCLowFtHJC1l4d
OAfqQdm2bvvk+HeUTndlOndAzTZyJGyjwGsU6OgGSUo=
`protect END_PROTECTED
