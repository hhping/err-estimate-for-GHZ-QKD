`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlR0v4l6ZdT4NvLBlQrNyrkLXZq0FlzTvUDpCpvwQjyTy58PUj7Dy3/wdPFuCBan
6jlD10BPIM4xqDcblZXbs2mjkq+39pRbboz/Y1NLUIj2kCzidePmvg/8ergonzx/
U8GQkBx4LTEhR8op8mCs3qp0ItplsXOt+9pqRUutBxWitkqi8WKUVM5+hmL3BzJ9
5BNWUVyd2dtQWHfBd7LMLfksAKzJHm1XjJR+x7Znzbdgd6boorLvY+ut+5l3AcG1
6elkUqstham9hl1y/SE1faj4/N18fSW0gyzkx4Tu1RJFNtUnHT07tL6yOup+aDp4
o5/2ZblXwfOYRLMEoG+vWofD2UwTVyIK3cZ7mJX5TsIWIH+rOs5grGrEJg6ns7Lt
mNdxtVc7V1mW8y5IesZ2PPLHd8/d0//YW/9LAAUJsmdarFYuXK6FzUmkbFQnwqHl
8n1NngJDZP81esBzuhjjUSx6zPe8Ekwh+MGVYGlVwoGavvDOCz1qUqF/iIYYeWEb
GpeGz8HNA41jv19wd7oDCONT8/xRQi5PVcVF656ydKxQW26E8evNUFv9PCR92IVX
IgzxsXsqLQXoSiTO4xSBc6QTujpyz8xmTeqeAUnXMZcr0pEoEUe2nUlHi+zbek9R
d0u2WvB2jl4ST3IyUxneCw0k/3DfcSV7mCKQ99u1VMC6jwDMegJeIFdt6rPuYDFT
Wm6XWSgg6HNAhEhblQX3e8oj3L+I8mW5zFReB3VO7VkRSAUu7BEh9+y6Ctm0I25u
3maPZHxdWLVXKp4Q5cNV1yPmeuIfZp9fmPbr0p+AASwGlyPDhLP0ZkDqPg6Gokch
c0aw0hCx4YSf3VONL6nDYPIgwVrUG0tV4k/I9YZ0N/UODJ9gjf/bh6iJ55avviV2
TyGZutwcZcMahoKvNikfpcGLBW0cbT5q55PVxBoTQrV8/4bMQCK7HDLlFznSU8vq
loPziv0dovVFL39XASeNGTJMYmB7RTQWRclKzpX0ewUVjD89wU+tOWwXcJdYC0p3
OOsk7eI9LYKysllzMxlChl4CJqZWjAcuETFeU09usU6KXXoEGdej1KB2JfZE1EbG
dE5GCQ6+osaFv0TPvVq4hGYwj/xAzujQAWf3W1n9DFDg/lxEx6NCKnYlO4vTqKIM
lYLaCbyk6KzfTb8p8T9T6gWbNtsRLSsBR4CZCiExiNMrw1Nv+4CcEYLbrPy+8aBq
MF7NL6lkzt+iKdvjYLZzFC1mwwqHhAwteTkSKmI6rW0HpqgGPGrT7zRV7ExPQZ33
KSQT5glcNJ1vX85VNd52AbRzKeU0H2OoYGtohPYKhWPVAhQCel7Suo3aFrKzedrm
51txIQy+EM8YuhwOu4kSvC/3iHX380QIOrF+ZTMmh/aps+/jpyxD6wqGavnEol5O
j8nEe/ctNlUO8mYWyAK31JYfjztmhZfR0DQC7bnmZn8hZc7nJpi2sPsPRO6KWH2a
aIWjvsxNrPO9DXDkag7tmSq7if66YPOezwfCqIkI9jEdO1adWGOlPn25AAkmFmcj
uU+gGx3XE2A/m9B2jpUo+POdegMqIq5Ov/RUcVLKY2+Px2Xt4XOzxAWXVqKdll/2
u+tOAJDe8wHeewpWV3U5I4wBbBJTRKX4g5r+71EP4Nd/0rzeGpNy+cSAqPDclZxd
0SDtoC3IDf8nNwUNFl5hbzJ/PtxaLEk76Yq03hmAwdWI79/fLYKvpR8bKTnBKBxT
VJPAw3Q6QjJpgzyLbutMBB1zlOMzqZ/avhh5RvBOF3PFM/KcqKGqYXOjA964ZhR/
ec/pMUszg9O38PgIKFAjXgC9Y0q14jDijAnky3P1R8LFGxfWB0WMFVaWmtOgB2q+
IofawkL/yGuz+rZdgvZX6mRqOnKDceRlWqE5YBzOKHYbEsnQrPRfotBwuS3uad4q
i4DJI98Rs/R4DA9mWNr26wVWwQTwjrVcGOTb8+SFoT2Wn9+owQgz2RcDGke/qu1m
Bof/yPnPPgvnKzIUY6r9oWBjlA80U3n7qWAnEj0BdFv0FUnetx5NTwgDaXfOkvBx
kn+YeRKtYU9YrTe9RiK1xGYw7JNYT6xzNES3hBqwTUv7PDK3G5f/Lu6uhaj/qoU/
7Hd+upmbgybehijOAOlliasSsbq7kAmcWmEmUwfW8hc=
`protect END_PROTECTED
