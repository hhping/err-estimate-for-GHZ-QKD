`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcvbIhLXaTIwGaEZuVgBqUSr+ZnT1wiIBShpYwlUmNnNRmqMnhYlZ7wItDu9thpp
VNtmwbXspis59w9gYkV4lCqF09Rb87Z3aNkCKx5dH92mrR12wB68rxLNml1hE3Sx
dnn9KjGz0sF7ye6eA61MjcO9dvkjhJK4mGwz/rOMT1nmjZRzb95a3x3FYIsGHo2f
sVtCXgJjFbfy7n5wr3M/IJAR9/e/eV9AKUsfDRktO3R/bVFhyXa3TxuS7UpLjku4
RWIWoVJdy+C46QpuO6taAKaI73PhgrlHUdGcIL5mSe6h5/JhYqsq9mt733SPKyDJ
UxNd8iy3VQtyDbsdCcaDlCPmVnT0EyfP2KxNMsZFiypSspHsWFvaf6P24VClCLPx
p3qrl8Zinynl9nlFo4ALNzjgUK7jVT2aPgzVpapuF53PzTz5ituijO3p9mQPBtN4
c4JZxRM+CiMiOyRcZDz3mMuAfz2O0JKKdUpzDfibQ8eziW724IA8VchjNVqU+nKp
b3O71O+WuFyvH5J8xanQUlDuQZpm6awcSf4cUgUOb+flDYmD5WwNVKONF5tRjdkL
tnN6lsBTbZDyx4Ocj6A6qkA7u/a3FYAmvFofQdltNbfGfS/A/tm1BuU5zn7YHpvA
X/fcnj5K29uAIiUkaPrRqXrcK1cB9FjQXMj652yz8Lvt6mOWP4+51Y0l+XKq9Ejo
wnOVG7JWgiAQ8YaLMKDKkxO1Usqb+OfzPKyjionLZ5Aixi0bMa8MW1ri78GjyQ5G
ITXezqXrUtcg055GKNEvPD/9SBCGoOZPDQsBqCoOyCvYCC36NybXGKx3Dj6fSduk
mJ+MGTmDlVGEfyYo+umy3vod+XSJbePLBwMtBASHVO/XCWZknsFwhlGmi6XYV2bT
OzmJorirel9CqbCVrBpwr9zGqqpGGpZsOIpXJHsdYIWGWyPjevuACiljRIWCJuo+
Z7U2RskG4WN04+s0Xcp/JWVX/N7Dx4/oKz0au8JdynQY6p379mW+ofpeyEROZJ5z
63anjQb0XO41991YtNEz9FrzlbjoqSS5N48eHwlKbCgcHivIRcD8PetQev5JlCRe
ZTgqZeNjOlCaj8+TtdI8dPqAQz2MIY9XGm90XwMP/zhqY8P+5k7QtagrSnCq9Pj7
27QlIgmnYKFlmveiwxXByz2feElCVX0Jcyv6C4XvH35bFZ6n8vQR90J7lS3roSrB
jhyvI65y6YeHhcaN47xDg2w+b4Ucey15o8tIq6jKVv9+4Dg6B8NbXE0K2hornU/G
Cah+rJaDZPb/sRv57kH1rTSGvidkJpRHIqvCXKrS2K2gYF0xtqhjqL0/mVhUo17D
EYfvpUDOih41HPTBo7jJrkXKRcc6CdQ1ihHfFrdty+H/MR5litsWmNUxAxbX8GIw
Cq0RQg3RZEVtJ8hOjBTyAcaVKP6MGmRaGVgUtCEqK+cTyPnWweU58pfxIxFfeglz
UK6jKlxNYgLWx+l6IexAWAz7pkmy9W02lxxBrAHl3jNl0Cx9s6jo9MC53MCzMeHu
yTw7TiZNYE0tadkRDM2T85AubXzF8+mZXXfryXqsty61v6Y7meQsDW5ClbQdZm1M
mgKPnRj4QtyctBSuv+D0gDTHmSqXqZLzIc2RHDamKzljQkaMB3Uk5Czi45XjBaBY
cMIPtbwl4iXwqCSoizh9aOY5mPvvX72zy7AnctylLZWj1iBDqljw5tobdkuhBoZu
vnw7S+a3hxk+b5g0gzjcB6b+QwA6h2O2yWMMVpeTJjKCSYEspQsy+j+BVp1Dh1iz
YIRTtWuUlpB75cU7NDOuQ77sp1JAWLNV6WBvHsSY1B8J23ecCTtVZitmjzwGiTNH
82c5a60fU0cI5S3mCH8dVNC44L0QMDPUo5+lZgP5DVC/5lxype8frTm8Iy6F+XB1
XGSulfvjvl6ZCVLe1dQpht1rX3HZ9jMQM60tABnee5zcnGnF1enqR/lROkXtN680
0NfqRE9g5rgiHaNN0yg9UJ1thYcnGofC8MFX3Bh94Toso4jdtHDBQbgf5g9EhCYc
qPpTD9Pr/ARgUhca/+Pu3gtGukWMm0kpxelm4FCm+I0E+aVOlh1vBFiGCvvXlUS2
4sbl+8oOeU7FKfHXaZg7SHrQYzpU2rltVXcFG83y+R4GU9K2ETJHpP4pzR5ET7No
LEMQA2AWd00XSR285s38gYym44INQyFq1BcFh9Oiohh9fJk4SNfjgOsrWZlYu9TX
Ky6dXD4K279J9Icqv6Dhs4kjChQBkBEqwmniWSJtMyhHPjUaiYB9r7HyY5leyHcX
Mps025yQvOLRbg2IjNwTynK+Z2Vi6XGPVERP5NNxmtGEr6by3cZvmwek3dYc9tBL
eriphoaXiyj74d6VBuX0ccNHdvXJxOwfs/A0mh0IV2hLG3TTUJkP15zF0RxK/oCb
vRBhJv4H413a86R7OfuiGvxadIsDEWJakMfhMQ1JGMn1eQaqirLZSeHtVvRsKbv0
x5Gcw464kodkFVNpzQdcZBp/aVjQExX8HCbCMor+jLDq+OHH8DknmEs3E44qcmbN
4dFo9610/YJ3RdU7EnnOohBdfIFWpkIMtySI1i7flhF3VBPJNsAyYJiuzSD6+5n8
AatEUzeIPuS9fm76XQHfYzgyjbdEeaj6iJe3PCpEstFozW723avhxe2a1yNJ8s/s
dbXw9VE+QzyFm1l51C/st0Ak22f/s7E8GNbJvRIDem8QDwjd8tfT9Cdcoaziuwt5
xbpbyjgOWL3V52xVdG4xzzd8RMoKsCiq9zBXRVLYTEhEKNcQM/H0M8sS0t6qxQY3
nFOjy04/LgZwWiVGZ0CCe6pd7V++mnwd66MeFTMO4CAeqoSz0XkxTqpV1iXylcds
5iMLtRuRRYUz+w5sHTMWhb3imSru4rbGCg0zfhLJL2JzNcpLPuvRso/4Z1Ca4agu
oYxqtwoQNFAz2g8iWrRJx134FD7pHSiieQOR9QCpmcxSY7IDZVgctN3Ie6sKI1+y
A4dmpCKYqofovzaeSM/Dh7KJSIG7V4v3vE2uZFKphMYyP0Ns2TT5VrR0aCKHa185
C40tMj6yEu6SyB+HljavT9uo145RoZt4/TRmIKGTktWwTq/Z5wrzZ8lxItOTtKcO
9ILVx56DQc834PndqmLKvpSuZZow5tYcgUi/pip5e00PQK1juiwEKPlJJQGQsY2s
12x98YDeO698GJ11wOMeBKlusT8NBqkZ0Ah+Zt1Y/C4EYjSqhXmOChKE6p4BsrY8
eOWiKSgpEIW75Tad65AYOXAh7uPj4Ey36cmdWasahF1sK2UOmyycKzjMGXeT9c26
kr3NHlQLdUkn8OwBwBJlD5zv6ri2tRBIT2h+nVMThScXJRMVdGYHSuerleeyo5Co
X7Qu2muceAqn7zff3rAKgWeVdCGwdLGPOM8NAsIo/O6AjSzjyz1AEOEtqdV8UwGC
TOmcPDQn5V9AVSDMjX3NitqebEoMc/amOXs/KkIMEzWo/Dt/pJTy4XmSgavetHgi
TyJO7tf16tslYDpsLggNmeO/s54ywQItBU9NJH82iES2mPDR89vz8qsBjXQnbGMU
QG68KuLnf3D0TqrWhS6H1zMeUm2nzl33/64i7Sy1f3A9SRdzhoDUBaF939Aw1w4c
C/Hf/LvLc5JrPXjccxJgzHIKZ0IQKFPzv2PmzW41rhaoELaC8Qp67Osr3Np6/1R6
Ve/nm0eIotDH5EVgn5kYU4rZlE3DpeOL9oY8rJLaJDQvtw6ZTkrZCihAF+CT5iui
eKEGjgNK9ARpDRTnitXC+BAF9fceC1i5rkYHiHNb7D7Qlugs6JoZDHiRUZbGyMOi
RH7n6FNe4cxOA1Z2MqrmvUR2MmD8LE6XjRP3Szhs3sB1CcRnShNJpkqiquEqVK+x
F0hQCs0aDiVqICFx/9Gb5PIuuJdZs+QRZW93sRHXB1TPQviDFfqyEsx16OPoCdAi
bOo70l8cagQt1T0UQcMmG00sYu5qrU2QXJBtL7VNaLmVx7WpKuhHX03Yqtt6/vff
TSm7BvYxQ4H+AWn72lOEMUDVnR+BKrR7oKEMvqGoQWn6hs0kz0I4nXcBlKpaYR8X
eMTI5TT193zj5SEZzBxiJNb6dgoplDta9kgjOTbaf043b9GQNglxuDL03twkD1C7
gCrL0+8ZVs2iTkMmn3os4iAZExMlRgMY/EabJBgdZseENPgwvSPhpTIdJmu9IgrA
eiVzZx4ec61QoRhnHprcEvWFOqXxRONCK494OhSA90DFijNq1gZj4EhOuuIsAfbI
YIlyzbnnxBwlOZzhmhn43qBgDaQEHbvatMgpHjHOYTgBCDseomNcCA8shAXdJOk7
jO/8sox4GBUJacppiaxT0AICWW5360uPy4+qMnNAtGWKxjLxWOqTW/HV/YnLiqaO
b2YymUz/6E856CNsuchrMB/VxwxGNdbJnUgiP9Xg7/bgEdlnQgmANbb7xBk0ThWi
Xp7Cl+YMslcANMiI1oQxkn6xId6/lSJAdgJWyNmdLU6n0RSpO8IMFpb1WkhLBgD3
dYR3hgQb2aerOwCc4HYLdEXc26dKtuCs8hVS3Txu6jUdgKG5a4pagtQV8qlrmufO
SwGYkoGTYj/fffGEa9OPcveKKyM4Q0o8FqNY/ZGTrc6x7f1MAWX6mY1Mqpbjn2sk
dQvLEXT967qbpSIlxqU0pMjIHphUl/f0xZoNx4pfjOcYw9D69hGp0Hs/8A24rzL4
ycQpZdurjyQf8NKa37l1tMLSw+PjHiKE7HlZDS25ZG5ysBU08aM1vj6IAM//MOPL
eKSA2+pbMORhsHFqmEtF3RZGctmqqLs7vz5yuU69NO1nujqBhs5MMq4IV9P0IDcx
7MW/JsVnhdgCRUtpU7l1+NZuNh48JsMPgZrnX73Lz4CDot0LjbldM9duaHLdLG2K
DLOQJuauyT/qj/Z2Nc6OFgeFOK5XwzPlpg/q85F69bVfjfpcY6D7PGK2N9fAGyPN
SAXeETb/JGPQHGW7XSYOlB2kJ4hkRH3LVK64vZd2qOvOcx+rGz2PmojM6dN3o3bK
KveDnuHWklRjBfPLQm6QEkdsg2OReSJb+P+bLfsNI6/ZGlfLj9FQYN6YbF9dLSxL
q6JvHD8G8VjZ2WhoiqsZ29ErBlH0Cj5sSho1ULIyKdzawIdUc6y+EqnMRS+dJRG0
dDtl9PTDvOIL5SBusKX58oIMabcIPW4zqbZ8iBrNJumd0VSF9Mo5OOfw9N0+XcK7
GJjYb4uMJxY/eGGF+K6/REMjDPtYUJfGgstw/XJIsCSwyrc8t406zqI2LbDwUOu6
NjkAEFcuH7rBYPhOx/4TU7cyNL8pevnPIr/elbnRB741YJn9Yth0yJRW/g8Yh7ZT
j2tucajwPgB1Abf1CfQK8aZ7jmKXMntaOnPP+UwFm7Iky6ICxN4NGp3KZG0g7i6P
HqBf6cqXg41GwMfXqYX0R8VLQVdGVaBiDAL8oLc21UKM8a6vNMWtYfEWDnd0KUjm
8V0+B9RsH6y1H/heN0mzjqtNEozmzeUijrEYWz+lo5AeiDkQhdfg4lhIPKF9nD9k
QglHMhiCWY/wu0SXtnRZR5fyvVDvm7XBIopKVvydLpwnayDDUYwNQ1yzoMDgw3T4
PaPug2kihKmmyamEsOVrdIxY/+NyDlDedmwgzONMcmwOPkNf9F1rwN8Y1g7of1Mb
4DHsKdQ1IeiSrQKcftKY3AZ5GkB8jftA9xIxh5MuijlvJYr0UFO8+cj3Qfax0tHo
U2R24j9j8/XVi21uCrH2+gdqM1/q/XXH3NglfZT+PmoLI0lmVphjxJeM1fZPOQN4
ZfgqSVtnuWisXZHiZYK1nOPAEtzd+AOryj4otsQpmk3aDVXkXgl+YlnoKPv+qs/K
dG8ZwyL+atS0HUc6w7D1b5Fdh/CBXeAKuMdfCMwD9o7jwB7SCr92TIf9GuMAOa3r
F0vpQ+umyc4WeN6eKiW7jFLTZ1PYMivykgLMwZVEbBqQuRNadBhaQiWsnlfW3LTB
u3de8ZoJFvSadDYN7hUItjnbJP6NFG8alGmHL89IPl6+RlJxpVqxnXV3XkrXCWtl
OcjJJsu1lf2O/lRW3gyJNE9gqu7RA0nsac/Ejno7vcmiivD6qr51BTe55uVfMIyE
PhrZ3stl8a+ZD1nBVaLIPhrJ1kNCkb2gKWYyoiIBN1yZItmBG9zJJI5ihJVDc8FO
BQJ7J3UcZdono660TV6TVlehnDJemP27KcupwYpt0m/7wZwELcEw3IBSM2Klh83R
o1sjoq0ZFv5bmAy17esXiScJAzcEd17LbOgCH32JGkogmtNddM31xTkAi/1FU+hF
OwNMmdEj4RZY3cn4laT7U1KmZCQ58Lbb+BS//DlDfl5dBxjiVoOw5OIfUnIohJ/u
2a2cpwU2BpKnt5UHwIWl721W9AYyq6DCv24O/lZq5uhg19pUE2bBKRHTOs8I8HKL
jYqPYmq1wvGFfhjxqluLcuBgr2269dbUQ+mNXOBOX/xQRLybkY5MSbe4Stkc+cgp
WRmZCRLJ/y0gDQPmKWDEAEbQT4ElK2DXSKc60Jgd5frmQMhn/eDz3C/kzs3ql1o7
Say3DPd9xwFhc73rb/VCBdS7PtdjJI5r0uIKWx6ojuHQHZRnHffwVPnJIUE7BKL7
f86mvU0jYFk+x+Nxkg9umioLQdnsFi/9523/girJ9wxWs1dSrsxN+Jn6cxPcrTWx
z45/VR99VdGfKogYTTjJgRz6AZWFuwwLipwScQ2M6xUurtRK4W/AFuQXGDKNn4FH
to9DfRunKPjG5yyJmRYahJVbvzDq4xTDYpwNC582QYSo43dVE0tJdC8enqP6Tniu
FT5t5vKMu58FrOOaZ+2qUyw7KAz/cG0RBk3LDhGG1sx28oOe6hJir/W86kO4DBlM
jBCRlaWKBC3Bg+GN+EepBXGJYynTbwD6db/PMwts2LhrSADVYmE+gqNssTvCqf9w
QG5LNGPk66TJjxUlYb0+m31khhACY2aZ04IE27GyFEm3BxfFraENsa5RgYjsqohS
X0Qa5Eu3tmGP3sTNl6l2T23bOZkX/fTqZT43mcDFtYjvbHraWY9oUZJ9cABOZ2zP
OcYSOCoxZ5omw3q4DR4IXUOVd4yaQcUVN6NWkdvZ876V+DjUXyPvRwP/bC3iwBmT
f9tKskq5JVcbISKUCcoLjs5y2HWLkq48vqeyAqm5p9N/3bdWACc0iu9uFAAtubgM
zmNC+K1XMf7qjI7fYwQ98ugehU9PgM3iwo/KhM8mX+2DA+otuQQ5nA2R0ds20abe
+MCaQ5avqh3JFKwyyZUBlQrLBb9tm8nJibGiVV5exuj+xV4a9aKdoLLFvUrXGKUK
g8NzFwY315944WE+1aUP/SD1X3WhUso7g3eMrF9Cz0QWjMcjCPtJHaNUTF7h984i
9Du9eV+GLcK5XY2kpjOPQwymuZd7XUYpvkwfy90gXRLnx7k8hOBRlpLD1/o/juow
55TREG/xAb92+b4E88twhwCNXLkBcb2c8zct7WRgoIVmCUTg11ctFbQFeWFl5Nrv
QHQafqGAeHHWRzwaMGpEd8OZ4HNki/JMUlpV5YLFl8mg0DtC+evhI2Rd2rnSK1bd
DrUJA1yrXYLLTRJZYmiU5XGe5Ky2KgRTiSQ14NcDTWUcvl86mhkFOnOraWweWA9i
MuOqyNiGQzCDzw8g0PfF8Oa7WTP5ejaBvS9YVS9H+hCMqJtb0CRqpKpEr9DQT0Tb
qHpKjdqYS9Ljqd7aQMiWlu4ubW5brAE9+BCuKoXKlvcjKcEjxhFy9ltMRVgYT7kY
ZRnvuhUzYzSfVyNiKqk5iU6oPQB6sJtGLFqjeSX61ZrnkuzUV/6K0kAc0vx/N4RA
wXnTP37qegBWxWAfIfNfPte3VKwN4bRxPSMpFXYf0tN5T5Rm/UAk5wYCM9YHKUhf
Z4EH9CBTPPmAtZUsbaH0SaqDvQ6RYVSMHCmyxjAUZFa+5UbbAsQ862HRy2yFA1/p
f4Z5mlhJgcAoRMYpkdmOlnYNUk6w24wpo53RB2doJ830EWc38TCFD+np+lOxssOJ
LgURXIo4qqQo2PTcgqJfk2fBQSbsaoD3pqPxmsZYrrICvGAQJneqQhkg5x7VpAq2
BSdY2gehkHgI7WEYuI+/OhoWEAcvu9sMKwsCz/OSNWAkppMjlvjbQOfU/8nzByRs
TZ829/fcBZAjdeb4OgywRaAAW6JhNXag5stTT4iuXUhcq0fo+tRD6PJ/8p4/rqP1
dqANHMVRXnnf++iPpgmpVFlvsrhgeI67BPrkQgP9J2IRw2ln28PIYwqZONNiKm+V
b0osP8mVJbVHkYqzvoJVO+gMB5TBfJS8fSiZm4+1Hon1aiNbHKQe4rWcsXmPA4RW
HD9QX47A51REaTzS9OlfOJqmJhDWc/DEPPvSsQJ9hGPOuQyvMB6YhUKUbriTBZ0v
Z+wfe14uPwGvD3kNn9KBOLLtHdefxNpEIcs/eQ8s0O+79wudP9qzbiDEgc9x9qLJ
qVQnnVHg0hom51saukLowtlv8M+lk34s6KmvJtSCZZ868l5tFlCM0LckVM4eW2+U
oP6P2UzGFHkdlgFi4C7xyWP69ce0gOw0tUxFUde+tqRNgdi1+Iq7wFMWYtr9E2Pq
tqHeHLogvYk8Ra1v6snI0n/1vMkUNSuggfiLq7uAlj3BhpqQArcjR/UhHwxFRaKZ
I1OyvcHft+vfrLmL9+tbHzBSRkDF10i/utNdcxdG40mv1LFkOme8qvkBw5IQtnXu
JiDiPdQWX6bE+WCbpbEvei0q7b7BtHKDooUYi3djEDAeEF2QpQTBE7JtNUSQR6Ia
HZa7pTnEFO88/qrvi3zXZFNc8EHpmlTD4IXSykLyvqD4IxLP4mVRoZNHWmPoSBve
OkVTFgfPd+8KsnY+M2gwuqbFmaxpGv1JU/V2CJ2bq/VSTpWGj5NtKmiZtPXfJOFu
kW6TeGMFRGCGm/4uTK34lb3wNItLDS1jbiKujPQdfWY5a8EfQ1vvStS5bnRb33td
Cf7u+VqVdJfM1A7vKEHwjNQfKz70PSLKWG7p1YIBy+BL3ePE0TPzcs9FhwtN9Lte
8GeW/RCMqSF+q6ojrOmYNUDdjRnOcvkg3sMYTIgWjOdNZVn62Wtygl4SQjnk1oJ1
x2p8mOcSJWGWPZPhhY/9YQLciN7zzcy6ZpzdFdTf11u7/OQ7xSeFBi9S47kah/cL
n5wD4spChduTG+IwVNeSJN+jmHP9niRS8rI9yiSk+S33W88UfqGQ8PVuo7df7GCg
bQHYHshcSNYOGoDuujC6uF73uFH9uvWKiKfDvMCEpVh6YW5VUsSigCnq6Gefv0Sy
YWGXjJ/9tqq3PmqbZn84N/hhEp0ri+AOG2/+usZR/TEt3qXtP/B6lcdH3uUCyFmx
BKNwXppNaUmR5z0vxoHjl7Bi+5UdLyWaDwP/LORHWVCzS7yu1lxtJIUZKB7KJIwe
5mpFvTgYRvHlB61SbumFDzUQ3eZb43EBrfG1v4R60R2nEoDfGe/E5NORZHTFrC9S
CgP54tC4anOMkfKmn5SBFYouoA5eUzTOQhs8hsAzMPpDoZTm54H4yFvKrfivW7uH
1kBeerkaU92c8ksYnQV2h7IRmiu2f70VQjNv6izJ3LuMnXDJA3DHezOpqxTG0e79
3L06WllfihuwOVLk5TaWM5Zg5her4oZGyM7JWlD7OWw0F6fN4cCH25Gn7ADNOJsx
iVeuXkSKqmIflmEWzaNUpJvh0MkEpy1HML+wgfrLGdAfw8uhgL2/BiifbbXm1/gk
h3/u3UrWZsgcbHK5G1ZhyBxRHupdD8JjQE+eXc21QIp5oE/qAGfp2qF1RHUznNFL
IOzCokKjJKJ5IveaYhbzqzUuTnKa7xPK/jgsiViJBL4V2h7tXDDHFxFwKTeSX2YP
uLJPNyVLqpDgTm5ehNIPqs3/uYXVaD0Ue5P18rCmAwt9Rdn6zwTaofuzoSaAExzi
Rrh0/wrRtRSxQC2SbP+7FN0d1JG1US7Wn33n6UW5ahT3hzM84cBjq4be6+dIkX6w
flXppkIhcYmYIUrntw3HrSnxWbqbz5kcxvvu/DnV9OiswEv29AGLnS+qIdCBeqGw
24ps41aOPtq6zRkYRKas5TU+fjvo/my5h9y8Z7NOclyaQtG44dEXCT1xs/zrfcBm
FCdP/w8kpJqsWd8abHxqZrPhKhZuhGD/WKJHGvNayGsxAs7TFfB62b418n+YHABu
x/jwByOYKLKOHaiQFIb0YD/wZhOJFNHl7prGJHT7lp5NtCDy70l2lgi5wp+vP+/E
RsWwZ9A86Fq7NqUI8ALpClhUqmrFiYAmOU66PyCwRLb0Qc3XA6jR45VNawI2ksxD
+ZFLXIndZydFwZCbL78mwfZPnKDeuXEIUO7gRMKDzYwBP99gyF3m6CNp+Ey7fiQS
Ms8h9r08lw1IpznYJkR+sEzWdSXSp+MJpu1k9l997Ia4EQWJaYtoYrFmrlGJdqy8
TrIjiO//JJmPuRL97fWtEFaW2tRlQou9P5neph/OpF+vlcxNzVr8gUEuGP/u408G
xS6QMpIY8FVE+AM4sjDqMdEUcNmQnfkBy9Ccr9DTwG8QRw0sQaZRxz+ZGzpxujqs
xhApQBt1zTgbuFnLVaaCd16x/u0fBlxaVzoE23Jh4oQ7UTbBOqPhuZzhOp7WtGmf
lCmOMytM6fRnIi4scbjP/ayi55EqRFjUodHLlCoPgMM8VktDIhRa/Mx7dPVeZwKO
37Nqi/lXjO4GXBB6qj7wfrBO77l8yPqRXgDHZFEwkGmLNf+W3fqrKqRNv6U3SSBR
fGaRpkprjoERsIioKF8OSMy2Hagc031EAIQBI/HLxfNBwXY7Ga1g4uYBPsbObCoZ
3ohXPCYjak5J68hStYDRK+19uZYfTiMtskNLDnq/h1S49Iv+KcKGGLQP76LWCo/Z
3iF93urqR/A6Zb9Nvo2kwck6pwoDb540wKcXuTflRP9kiLs7R+CHAW5EUUHItsoI
fP6pAwW1pIC9vTc9b/s5eZuW519M/qhIVzjCO9uAkjwKqO7/WKJ1SrvvcHAw/UeW
WZSGnPn/mDznu3Dprw4495ss7aZJ2GiUD6+JntKAb99yA5z25uUKA9pnrZ+pyO3/
i/FMd5+SPajl4+bko9eQVqaowrbSJ97lLSqRDYV07+Ips9kvRMihnPdO6p49jJCf
HAgu5JzxcekI67h1jwNAJCplGKi9E81/prjvIPjFUF1NyFw+Ke0xREtozDkQnkbY
TIyNv+c3usqg7HXkIOGhnzksl2/hgX69wDBumdEjWoy+ZWYwXHDWTJY4vM+yGcVF
d1LDoFj03/QlnacavZItSWpK09udOJvjw4o/VLqAeVhgU3bOZbKormFYJVKvvujP
ZyUhrvYhBGKDn3ed5NWANexrEjAIMD/2ZCuBDcINKtoekAW5Ar4CMG5nDkjQUYC4
LbqesvN5wU1eXThZaoFpM6FH7qnWs65sC3HSiY8q7sHnHRrZ9VLl93s5LNox/7yE
jCVcMpZj+b5cxcmUveMncxEZdXV4DK6rxRMV5RmVm06qlLyOhCg9vtW+SeDx2bmY
Il5vjmzR8NGj5L52F1/OFfw7KG35AVtE7SbaOBf6skYZh3y63VVp5hC6NHXKjWqz
5Jzjxp/w//ALmXp6G/4xe/VZfQq7gt66aEPPlX8fXPdpGVjHYSbrzNhx67GGYnvb
oYZuFsjFgEpDvQz4+GgWK7Ns3okb5OlKIPxFbPlKyhMLqQwtcuLzS6Va1BqxadXk
GzW6sJZln6actx0jYcr5V7yFTG29yjlvuZaEaK+7xAU/PA+mWwH+KWiwm1OIVf9l
LL7CCtsH/g2uI0lgWxTOTDfL4Y5tPqBR0Y5g1jyLXXMGGx4aTvXAZfJPpIIWsAgU
WLmUpK1cjKaVT0R6bQLuMNi4lTN8W+fQYdJKRAsWG9iwG4vr5hZRtcX25wBIJwaI
U0z55kVVhotEH9ErWKXKxRiT026upYRqN3hju9kFCNxNNe3+jkeQ2yo/4il08Apl
krK1eGhYJmRofTZh6dSwdCo0v9pLevT6xfuNAJCnpb1xTNDGvt5LqwvGWJwbAtbQ
8RR36lh2a8PFq/xp2+9f8iMF3TKy8KgRH5ebRob4jnfpYd1KyKM+6zbvxx1ZhMUB
3a/qKGGphb8YUMT9gYpKqSvx7TMHqUNOUrXiyq12zx0zCL9WXEf3cFNCJDoGolWA
BU381Jj65vKJxaISWGeEaQ99w8gxPkc0mMnHd82KK52+f2aozGdsiBUKO/2lsfmb
j23l+jz9jjBIq9Pzeos5VhH1ym8bV6TSZNmDfEnNXAw+zAjOp0sEmpKjfqsHKEIa
jKZivzBVy7CMD1n0pQ/sDigo1g7RMvChikQ2l7/myptBX2Yzmch4/JZ9K2q56tXf
2FG5gqYo3ev3njLuPS+7sFH09rnMub3foZinQpxbywF/1O2ko4bc9PsxrzwJb8L1
DpwK3c3Bxp9JtS833weixgzZKfQtWGLydYVdx0ji0ELKMeaAVi8+zk3KDrJeVWj7
c5xxExVEsXr8g64jdyzbQXMCG+qv4Tan6Ofo4N8vVXKoIZ7vl7FUa/aF2Kk6dU82
2lEKMD5r9QFo6wtIH63jOdrUhO3Rx4tIMubyfYqZAYFujtHjzH5NpmBlkKy2uUi1
zUrg8bvn5jFSAf50UZ+7JpcBZjBrqKzbou9nYRgKAcHIvVeN0Bx3eJKZ4J1dfBX8
QYqtFGN5Yh9tjHOPDNTNmSN8MPCuMFesKPGlQ3IHY9jNX3yc9aHSgOLkLv2kZXEn
Jzd/i14yGubB3kTGVEX0c40OP8KHCuqujeuXXYKCGU7co3rIUIK2Z98dMpgEbTKj
NlDwphkWzerdcpS4IEzC5Nl889ywPJWK9fKvfel7ryto0NZ4veKYGaRAsswSDcHT
GQyGUTXUOfoZtKTmLKcJniQUjVf87V5Q0ZGmucwlkZtfyeVdCAwiG/kdQ5+s0rrz
gJr4kQ9jqfRZDL0s//kmXJ8Yl5gjAuH8fdOX9xBjxOrqCaSiogFnn3BArx2KE6sb
XQMb0bBoXsIIzTyyxPztBrZaLaQbyVR8hSAYghlJkeT5LRD+p7wF6fypUUsj/NND
kYsgEATffE1RwmWlipzmG4hGxsb0uHwuwVtZUN9CnuqylmO2Tt97a43j83Q0gTt0
xoOvvWMzukGDSwmJFr0gB/TD4hx7H3n3ipn/KmxRETRjdfq1Wu3S5Wd0VyMUPH6j
B4Yy/RFckKq3cuHkgAUXgRS2bYnnsvnzOUB+eCo8K113q6I0rqNnL03CWF8+WBCK
yc84emkzna9luqgXML2g3SXE2qhniMroqDTKz8C5nmnSinLQ5Z0d0OOZYnu3LRvh
VpWyugvnhf+gRRgDyQvVCSgDDVd/cRfg0hqNR//G9x8QA3jgTT7bfSJWEa5xwFSo
u3Qb2j4TAEY82aWBNuyvBU/MWt76a1vblA38rZXv5wyU13xMCPSlGV5rIhZyrPE8
l6/J2YHP7DRoZB/aCRlM9P1g4oE2K1lctLaJ0xsk8BCM1qkMA106aXj+izw3LGFZ
e7H1oeE9agNMY1iGzOsQZfHI2FohcCAiypOBxBsx4tZmsUjKPsHHXl42zTQzmDb9
uonXuJakJwXPKmqHdspe1kHh++TixLN9LmBAsMZJdciLu/tCnA/saEngxIcumbNs
5CSGWSgZWHm3jcSDbBOmiB2KCe+M91jfcNR4YnpcoJzqMnhfe5+1nEk4MJDplvh+
c9k1sS44HnhKztMgUoJIbdk5V/WvlWi/fXeqwRhW0AstiT1Io0HDHWDAFW8544Uw
8Ns8CnHPpyZf+I262Gmp642v6x4YSxOKSss8iF16cl2aEIIHcF7qdnc6B8+6nMAj
V7c1i/4OgUrrBSyVe1bZLIRSGBv0zROtmWn5mCVAbTc5xrV7E3axUC8na9sAHsGS
DIJCUoS9XxVHGWS/VlhdIa8KhqlRhYU5wBzoA+oz67UrykZgqIMmo9NVfG6onmIy
PDB93sSCnGrwZUWe4JBdYB4EAvCV/hN9lsIN9HsaSQvtV9bPBbif8CLcdveLqwip
tYHlf6SNj/SsAJvtd8bRNdOSOUn6lCs2PYd/bDgQhJOc6R1fRV9WZspy0B+gk5jC
rHgCQgKXJ+l6QfguV/wF007pwK3IGbvs61GZy5p/40Q6D+t/eOd/uWCgWtItVaBq
eNUnvrCkLrj1JbA65MYt6v+btAHcr5rqV9iYrm2ZKhY0wietY7B9Knb5TL4Z9WY1
Ay9KgaYDVtuFKj59gTgfmMkdevj1s0JQqJSaB4xDPrzRPsJ6Zi9WMG7V09RDPCXI
uI1/zi6kJ2rx5o4TWq2pOe5vF1aHF7BuMdTx35gnPXShfH9Famp58ryzbf1tF5UK
UMMmUMgmb3psuDPUGbrMQ7QMoMD6O/MTPCr3tmSBKlA4TWGYFiP/npBxDkOg+ZIF
prrQAPSLO1H1yOsc1mlaYVhF5I7yPiqigTXxYmFK7+hJ0Cge/DAxebeCUI/Wt31m
dUkvqfZK/HxuP/jyjgXDoKikKmq0n+q6hvTu0ULDX71YzEI9VEcs33DlK9Z5K8NC
91LkX5dsjOwleV3B7h5EdymXiyCuttRQ3x7zvxUsM9CqSDf22VnNYlYgXjxUiSFt
BXNeF2msjIwgqs8sDbI230aORsoVbX6E7gANtyaeWxYkKGiOALMZV1lz4xVjdTXH
h6qtqpnVTT6AJWA9z756znrBTDcFBlUX8Kc2Z8IwaItnveOuTnixTMLJSQpUc08Q
uYPOpx375Kzy9JPcy1I18yd/dnzVdxin4WLd0Y3uu+bKnrvo9YPdnsjefrXyn+4+
1vEQL3BjkB/1aiDiFYyGiN26fcq7n2lA2EZwaAc9Ud4OZ/l8t09Zl5dAqs0U/7bP
Eb/INL84FEiqgDG+yQKqnfj1S5bGevAFWprsfUpg3CJErb8Q/ouoUaclbsB/zWzz
+AjiHSEX1sh+SCckWZfQ/vJIkLS5jsmMBxtDz4t4jmy2mvZF9I9FFTPlh1bb74gM
TkwqSHTs776NNNcvNMavEdwmUzZW1J6acmrFsgtUcXRxRCZLzTT11tByWu5xF/fu
5X6P5c4BEV05bc2TWESNzFOpMc+wEx7runSWMFnUfbm3LeZN4r9ldFC4gzS0EJKf
GV5WjwijLQMGH5UC/IQi/m0/j9AfmTCPWpzq5ZWoFgYxKo9MCIEjvk645aMG71K5
IAJWFhPlGUlbBstKTNlOgpdgqUBeTLIaTz5gLCtIF16IXo/afP7lmceCvhwZ5Ts+
9UrIpyVD6EjI7KRGmtt5E+KU71/KIi3sVCjgV0OjC5xdh5yyx29I0wTvDmTzAAO6
H19b0DhUU0C4ltkvNatvkUSDTr+PFb2/X/v8uA8ryRJckHO4t2CgPdwjMdnZuk1j
y9pwM3lvloU8L8Pj5g+xVmNj/CQSaIUvT3UMz5nxIMq8XsNc5JFwzO3QKaHFndpk
wF9a56681m6KzRlqbIl1M9vhPa6wG/EzxClAX47pk50QU/cfAEHyl0DrJ2Smd9VZ
hJnCnCyaTA5G1LQ2pLI3bRP+MnZdvmUv2QT/fX6B8YHkdyxFXLA/pGQYzJhCOFLw
i/px8GSbDx/asMMnrkWkS1F/YC67gvExmZOmwggKHJJ6hrB6ZFBQ9sWdHscWASuO
3rcjH844MzzGjAuiAcu2z+ii7v2tFweUhSH0wuu1dfhOxAilnDYJ4thbdmADFi0P
OJCq65uF150iVYlnUELgAAGHlAkTcqGsIG7BtytKcYFr43PGY1RC9TttoN4Z4RGX
+xO4+jDr/fFr9kPRud2ansbkkiBjOkT5+fSLDMYXWfM8y5KEKMvIsWScKI/2SzdF
0+5ARGI94fu9bVi9/3NNGN9k9ilT/ABkgwKVI/+FBKYhHdNHnZ7Mj9IZ4ZmXV/pQ
VjxX5yEexLMK+jh6ho8KISmLZFiZj37Ew8zp6nXT2f/7osMqTQb5RNQzEaWHg2S7
9IhZnHmKD0qJWfkeFsfN3Q7lfiMC/dnZYLb/l1PXiS7gFasMVcCWevO4FsEuDLUY
cFoYtxDzueeaxFpTgxTx1CZ6FAU2XLs0fl6EnqjJ5Fojo8QNca/Db5l1jRpX/zqG
M633O5R99oPTHrLYtmomxKpPIpKJo3KRUiNxLLpnuuf5AuTdEWLyh+cihyCIopBX
1ErgzCfEzlZamaKG3fL3yw4KTL8nk1TLYOWtaXWjUrwlfLJ4cbPE7elJWhOHGFaT
BeFJCH8FTriJIVTGyGH0N8dQ9tnUynrthxprwy9zYp/WzaPAIAL55pGp8rKhiT8u
jeojSWvMjPQIOQIojSU8jcbvB4dwaKOCDDYG0fC82zBSTBoy2rHUYB8cZVdwcaHg
kgBiF8S6Z0WxK8WVtTslrrtu6/OJOcK+gBLRgjL6Z/OU5ywRSpuVR28d583Cb2d9
kvAXwV2/KFi2IKXP0dq0e2WNcyl5uF3sp0xgKZDbsshEjoGeh2eHN06FMty5wcpq
oCopwB0x9F7yGPcPXdijopKwcZPeTdq1NpL+rEeFgJZKJHNlYErTjAGTJVkGQGeq
UT0j/YbN9L4F8Pb9/SvA9cbLRvxvl96fjnpDfIJvm4E5ml4Anhjlx2uL+fdo/9zp
Uju8EtvASQnJloCiUeiucWbrlX5yFvwiyNal+pnoWLnAeHR11TKnXy3S6EUW1Uep
PSpxQQUG1ACUr0iYJmio9Um2cXf88acDJGOEkbGjds/5RRtKHvMXA5PidaV4hx4U
J16TAUswKa6q0Pu1JAi+UaW1/YDIEaaAaguWqCa6NA49Nn0t4nk4MRpXy6B24u1M
NtOcW4b6IqdxYDyJDbgcM0E9aSPJSi7b5pH3bqlDDhq4/dVHmXbhXtJx6D5aqrdp
Hg8mrfe648kN+YFNx80qjUNWkx5FgzEDm+stfklYQ/2hUyc+2yiaSg7gtM5GWjvO
4fwHU/wnoqKWh+5Iqen9D4LpF1Xxr22gXQd0lY4A4Wq0/z3UcM5KYIrGQ909F9L4
/b9iFVKcJp/Av5dqoHOI1XhgwA+xG7rLspZ2JzcV1uw2yZjuMSof9rqUH7stwAkC
VSORZk7eHvjRGQn9bpl/f8OzySfe9HfkD3CBMvr9I0EL7lUabY6dAJq/I88phf09
ZPKm24DA/hOGCvHVCu7QKkzHpl9R2gXahj+83biw3d0pBTVom55nUCiiGHpqpIfp
SLXKIbO46JPpI2plVBK+LkaUEzMcgeMgFKio0V7YL+vw0Em5+Pv+VS/yQaGYNwB0
b7Yz5rp4D8aWwNRedS3a/70fjItVQjyuSrWNudibKNvF8B+WzPZ/jlkjenEYieuT
UcxGOUz+tbGLQe490ZAuOdPF1BEytPp+yWEviM0UHDVuOrAbNFclHEprIPOBhsl/
j016Fb97xSssQyIFvXyWBNSZRzWeObJdy2f2ERy7xPjJGRZu8psfaHIb8u9N5yjy
ryp+PyLhV8hMe1L1iALl2s/XcA39heeIQ9qc8HXYq7knEJdS6sJl1JCL5egLP9+I
Uwo66ndxqdTAonab/Eh5pTiqpP7bZLaAoiCHCFX8omakhMomd7BSLPf7FCr7VU/B
PGDYug07E7NPFw41dNdQnj5PO8zBEEOd3blAlKC90koVN/rI9mlMhWrifHr6iR3I
6m5qwpqdlIzMBHt/xMoeEAP3uXWvih6zQbGsLk2y2ddjfjVZNFEsdll+iCePaa+O
BYr73slRcn7RIiT6+0Scv/TrQFdjdBKfdocDQ3HV+HIQTwKpqY1IuseNUBvkAfoo
P6ijievB6kleCvIYCEczSvAhar5LaYax6H2Ghh0oGtLqqWVqEY0tAXqWG/Dn55hm
OYsCKuaa/moTt+t8ECKdGq7399RRpj9NKA5Prx2BtzrMxpdQKhCV6QaUbIerGkjC
gkGO1ZB79G10GVeZlth7KDvqaGniKe4SsEmzc/boIOzrzMpkF+PoTSO+GHUbEXtb
FjYUQjabyhj40nzLMGVI8zVIeoOoUjDOZpWxdo9vldVbZn/ROECubmaXXn+LarMe
7FH7QyunwYdW4/magl8GoL4ZCcaQuTVsQiRhMnCExSAnkddKe/AH4hfOBROsQ3Xt
UV0WFba/s4Q+s5WeYnaG4L4QeFQgeSSHWHCzo6biiN/N1RQJN6VNkTetrpImrIy+
qRmpljK8DlZ0FDhGcgpTYSLpHmrpodLZfoBM4Fn0tgpvz6aGqP2DAkVWaIwgay7f
OIVq+wItWfNHXQLVSjSLIMjdT7dIYvMwG46LazAGiYNznK8E2A9AU1a+tp3Ec7MY
mV1x3DokyaF1Ghy0YNCx1FIcSXEFjQwqZiDIqob/sIGNcenrpa8SSXTMOUxcxD9F
tQQF3cFNVWFkSxfPGOGa7hM0n/dwkj2J9JVe2gWDH4/PhLheVxh86djjRGlt86q4
SsYecI2Ge86+U9qDX90DFFZ2/PpGlvRdrxcv1z1foyh9SnmxZbC3PZXeCtIoYq0l
LqQSkH131xQ4MT0CBtjPQ5FJckJhITYg776m/ccjnDYaQ/uSmi4Qo/+Rrzbjqq3A
3sTOIkxkecAitEjq1A6Tmo1Mqdi/g83dY5RFzCtF/H0dCOUe0Q0AtDNdHfNGil23
wQkayDSnRgIEeXnIM91Hq8ZwJN2GEDYi9DqVuP1jcySlOEtHLk2bIOSXTISPWZGM
YhHox5ucLSMF3uwdp/mPX3t1k6wX+c6tDoj2lw0sqokzfddZLN3OauX9EHS1TOCO
RxdLLtzdTygUVcr3J1lgDywa336LUiDdnYpBly0tcOIPNRiRRDi/u5hSKJEtqon1
iK/BHOBi0m3pk6SlSQSFT+uiiy9tWags0TaQFbaeDI+XrYrRADkRJVQTpGzKDf2s
diCAVD62lumoRoujR2Dmb11SoTNpViBf4MJ9oq8gTzEUU7JNNtUNSD2TNtllwBE4
uu/xKCoCwWpSSJhO1rPVM3W844wCk9RwrbjA9902TeTHUdSkAtTFcqFw0vGnSpYu
ShdVruWQAhZ+mK8zPzeXofUqOJs1mMfGmb7WZheNUybKpAvp+J8e9ojPiOhOSPfM
GiWp2trxr+tIlfaLX3x/x4D+QA/tzYoET8/ez8A9wzypyxFxkdy0yyClDxndfTIG
lOx0qBAaWR4RLYwakYqHwHjWXfQtJ8yGNxy5DblM7mGapgryzQ4PryApLUXHlZH4
D9xzRdDNaIvYT50cU0eEfoTmcrCT4IQzl8Ev/Ue0V8KSODq6rnCQGQhg+f6du7vp
4zZajh2jTLEDjGS3Wv1CTO26ZJ4RRSyPvpZohDkx7KEZadZ/zvjnNSmh11DGlOsD
ZWitmbs5UxibRnFv4Sh4TzXOBMpOgkZQYQuKL5qq1autN5xkY+D49PhtDXu/0oRv
XafR+jKNv/QV407Ue/UwxU4J+C7jW0/ZBqq7hB/0osi2qv7AnkOCulDa5kRQsSBB
veWsSS/B3A6mE0x1+yqtSoIegDhP5eiasaQpIwMqSmqarzsZElYWnJJ1ilf2+7r3
KUT7X394xUOdxjWviawTuu+axxg02z9xCLH1lz+cayK6RMlYTxEGGTiD3az5FkLh
dwRuefPmRAAkGF1YOdpG5bcWIMrsKGapYjJTL+PM4NGunezPInnshNnOaV3s3UAh
vISoQO6zrseg9d4HbeQjPvARWA7R8xpEqMDoVkYjHGLfZg3UGG7zP3uQ6IKZKAxs
pFMVcxtS9mfzEzJF8sUqFvhjFwzOiHgHAX0xRS3UBuoykpe3Rin3eDcoogjuk2EY
CU68uOwxEbLUFySK5snycHzdCXsxwhXOdeI5+vigEpWB4SFXTPF7Yh7Be8mOFALQ
JiWEnvEA07bm8z7IFl2vOPhP6S94TLtAdfA3LlCtL5p1hA4PiC9C+icTnPdZZJsM
8DmAziuZFkq42XnDdlb0XzB/bCCuhSb7AAXLWzOU3XT60ONg6r3Ch43SAjaR3G6U
oYyao8MjhJLYl284ztpbzTYPKwX6H50kc6Rz+fM0rU468kDC6zTdSyLDXKOMVdRC
HwLOpbUDGeux3/6AHBwDPKdQrtzStf8R/cxmPUjjvzJtgRzXQ95ZPbo0bxeY+4Xw
R7e4kcwbI+DWeZwJrNfai3ljdYXvynywdcYvYWS2df9WaUM+yykHYOQnHW1HQZvX
/3skz2GaV+rbl1M6xdNLPD/yNZsiALIRBSV4Etzi4ZY2dF+uj8aR8njte07h4Cf5
Wqzkz2mfQw34X8aakcMHa1q10uxQ0UQhxr+8givE85PNVF6OEnR4MnEj8LU10XTd
72/27hNcdEAYCMesiFvWYbYu/KWlMasyZu54t7vT9M5PJpkeQu+6emWFk0kEG7L8
lmmyRwM7PFO8XQwWp9OsC1hJxCgvyAkO+WEpg53veOY8we4p7vUZ9P3ZxPJe0M5Q
b+vtEczk4IwXkBaPkvReKQoNHeoD/IXaHV6+42cSDM/zZzrgMD8ocUTeAzmtrnba
FS8CBrobpJmfVJIXAJ0EeNPzeXw/QoEPXGX0hoaet9qFXmpPmGwsnr3KNdsCCe2W
+F0DktMLlEbSJpswOCPZnkwipNUweYOGOFNBy79/rtZNbqo7fvJM1f/qOSxNEbE9
W2AL+IjtJ9ffGJa1yw/GywVef2qliRgcS/VnS7vHf6bIY+WNpSp4NTB3eob9k91w
BVCiLZxOIJFIoXc22lTMQbcfgfjh7XLR4Mv3iEjgAN6FsI/m/wBWqgFLtHkwX4v3
y4cMvw5CmZh/2AkIVuaSfAgFJDyb1+qlI287ua9rIcxi+FE44jv+JH510Yc4zP4/
rFL3j5+Zb1OchxwqHNCjs90dTVMYEjdC4CbqlArijTnWt4QQX3ePBp8yO8rzA55v
G9uMZywSf0P5QAHcYX47Kxd6nxc3aXvewuvzx5eUQNcRFRK7Yk0xdftEVuSzxM3N
lA1pyX96wH1MQhDed0yCyHwUsBSwwOdP5KKTk7uSU4x7INsaUAfSl02ctk/oqNMY
MU6IjoDm86p9T/hod0ULVk9Jb9kA65bEk+ABd+swlwBLnKS3b0R4xBbr/R0Saqzp
oK7ZdoP6U9F4PKyPB0wSeL1W6FqPHguhEJA2zMO33b72IP4t17zhL6puMniZeCuh
ae9XY+buXhnPuRh6p1Sd+81B4Gfq9XpBYnGDzemENspSiIJ0XMf/IN2Y08b4ofXJ
8RWRbcQqTEXJ88/Hzoz6UkKXaBRd5XeHBkWug/JWFWwpM0GypNq+PTnDD0V0XgtA
1VHXlg9zYPKyG0vsPWlFV4YANtFX/nMabKYdH4+Gl+qkgYiHoIV3/rSQ3evpUpSy
Sph0mkGEWPok/ksmXi+uZ8NGxSYt+eIe1Jxvkk7SMAK+JXo//hgURbZ2RAMQOi70
8puK1Jf1QnsmNmCNxE8Z6ADQXFq7eT6xt5R4xeUzcqjpQtrJVFfly3igT7o97Zpn
3WpwL+B9EXL3ySvLj6gVUBwbPmxeLmm7+cvPa/ALhHtAHjQ2pmf1CZNbaRHEEJsb
qrXWgOHD/XOKRdb/90zOtsDLOzS0XlEuYDUZlCwxtrX4WAksfpI1dV3rndMt1jee
Q6UpQ3Ft4k5Bg5dY8UJxeuJwTVsosHGfPcTd3D/VagDEg6FG7Tau6nUg5j11v7Tn
9fdaofU0S0RIbCgdIYRvZxmdFUdD/O6TYeMqdkGb5iGJdeKKITluWOWGaUKV/1X1
EqImRPPNeq8ypPTSPQCtl74RZ5BoelpX/0JHsGCE3GZ46/8TIzdQjnJxAZ/JqOHm
TXIshg+pH0jkXIXh1i+PRu8huVPdzA3Xy50IJp6f0GnKQo1K8n6C1ViI0N10h1xt
hwGaCOIFYnm6eTnZzYkW5vMwCODT6VLVtRK2H2wxHAJR62UZ7gJr4h47KYwaQAZD
fqxcOQ9USXnQXNlt50YqcBSjXeRjesC0i9ok29qFc7eQCKc2wMCGtS/mEUaJXm1y
vGaxouznkewkSgbUMXULU9xaNWRJ+SMhIHfNBYfBMhMo9lfX5FgaBrVFPrzsKpeX
JTOgQ0lYSNFepG56Pf+rWGMZYI0QXByrbjAKP2VdEPbquxt5dslB5cm02AeeRVmf
9gTiY+CTMeg2FbrnSIiM8i+eGVLzEhO63jBFSRwETG6zi3wPXY7xuUhjYouxflYy
SjUJecZyreSf2wu5KycxRLhCmaSuYCvPLHtQqiGf3/3zb84aISRpnWTuuwx8WGkD
l1VcNVZhQEKMzpn8X6YbRVpPQcAS0o3tWQpm/0leRBCrc15Z0thedGw/VknjXpxv
Rs6GXhJzpkCEBfjrqXpzzSVSdf2xseaUG2VNU8Qy94TeGRn6sshG2hlXZH1yIvI/
AKab3M1NT8WksOeMbXq0H/EEJFtGg5mynK9VDEaAyJyqJiV7zV75FH++9e9NwTn+
Q8MspW7lMuFcKK4GRTLVbqH5mF/I/X5WimIaUowNbNuXo5v/9St3yuvowEDGU7oL
zX6n1R5I2QUSID2zeKpwxO0YzQvgwB7pNvaqmUK+aI7B8gUVnNXPTVysWDj1ITM7
Q4ms/OuS8G2ai0T+0zWVrPYR1945ZYycV0H6k/Q0oWWsu5K6cSvMS33c5NbOlX04
SkvB9hdtNZ/5ZFHFewRMM9L1OK30oi4oyLFA8zlQEH21A118GIzUs+mHg9G+jqQH
x03R8N0dzxOIlw9UfXYjtLEMjm5o0sH7/xnzeTMweEcOYF0YsqtIPdCDIrrzohoQ
baF935f/GWMfKOLzsxuJ4rFGJo+P504r8SWdtbH8M0TCZcMW12o0zdlEvn9OZ39d
gOFdCr8C7IabeHBbRwPvVX3rzZxWEMETAiR2HSDGxjoX8zpJNaPwMpIK/fF/Xd3a
9ztQ0FLOloJUqV4ALj9k5gLomByVcNDWHJMbnEtiZI1+11nkphz3lJ8IBEKVHm9f
hCYREQiWqDa24co5MeRkjZSgiIQspGfgVCKWksVE2nnz4neQWIgw/QxVeVVjlR4b
fAZjzwEuV9JVK3RQ5rQMrWq3efinNK5xak+YaaVztZR7xXlsyBFuaAQ1amSpk52f
rZnGlHaHGu6py2MSUFeC0gUzHWbzRK5G34JZHHRjTqhbSGXTwc6biBmuvnjdgar4
+ea+to3wy2zbCU6eoNsCnPMg3UbxCFCTtYPPycFN7XahOpOECrHdxrnjeWvCmbmz
IwjFvZx9Mls5m/DkQPbjRMOv4qH1+LKG8g33M8mDO/Z11e1D6llrH+iaAYxKjgg5
xFvfGM/dznB8WlEbYQSp+dHnfVtY55/cgVe3QFERvQezNwiAv9kfw+TR/JDneP9U
ebFlzhSX5Lr+7lp3ofBnCjB8k7Qb0az1+BR+S+N2N8b7tleWH2fnAGUrOnR0pkz+
N4aZHvFQXuwU1GTK4qBHmF4wkxCGKwZRV4GRXz1fH8GTbCo06tGEFsNjLtEOBxAA
Wz/zCR0oW4bOrMBGa4Q4bjpmLTGWpQ3xI0mutcKsxz+a3uZEd5WOsR8fVLSJmwM2
Kp9AcyPxnUtJNwtuUr5altTm9ezU1/neet/Lg0eomlQGcMUTfRjePpUUCx75be32
xJx8FQfJIYa9KmlGWxm2Ppz19kOPyZwvRvzd3AU3rXxaGI905EOOslwZGSfpcR9Y
hgd7jvrleLX55AFFeAJddbDu0q8INOL1aZ/Sj4gaBBCMiuoFpgxKUsi1OaIDM6//
G5VUtiDtZ3eKkwa+km9liThXHRNNllDPMJBbRg8kY1D/fZxAmCNQgyy/hujq0048
gcKIulfU7rktqeeyemQXm2OLwe2xdkXU67Q1H0tGdnslIWgboIT07bKm5ghSeMUV
3Z6TXFWlSLIzBF+f5q36FLlb+mnPEaevjxlud0iIn6VcHqx720RhlRJq90CocYvM
S1KFiSaTLWBpEAmGPqpIrpnDYOUgPrh+CgUjkEs9GJ/pizp8Tx943mO9rEKeM9XE
x5pMZjIvh//NWiW/h20IrhmSaVTBTiC2xsoQU5RWxCuw6XUFqkPcCVajrTR5kBo5
OMF58X95pOrEHRRnxXQfV6FWh/VycNI7lQe06xLoyXX+gZbX7La/EYn1Y9LqxPgI
bvGOZZei7DmzfbM8vdczsSAH6n5IyF7b4RtVdHKJsBV+VBAESzvao3QqjBmbpCre
dbjU12ikWfEm7b7+GAcCVWzXXtb8F2sKQKqY2+e6IZ9LdYtXBIdCqnngXCNBrWPB
FctWubG3LRQOt77/Duvjs/EdBqjGglDcOOLxKm07w5Ykdt5M2ODF/5Dv9+ihPuV9
4b7qJ9QVjoMhmyVe3bZFAoe0lQZFx4xQISp9x5nYbvTgSQlN0shSa4+noOP6xHss
a0d4laqZrlx3xjPmofj/A9ymW2jCFNJ2fnmqVFTMuwppWp+AgCCCCxctsf7UuCvr
sdJ6A4GN7EiryKO1cr8T2DdG+eyawbN41RKSOd+J3mj6xyMCKhZQNBLmKUDmOgG5
kGjlj2QgvU2DCXGriSrmSzKJCXwtaHP7I6IsGPNyAlqabfR85H0CRAErSmlmzq/B
8XDv/gC5May8UZtuora8hnRSUtylt2ocIkS3npEAOJrYphXBkEJGsT35OjB265MX
gzQSicYz00UWONSgADmFnjrBkpjUSfGC0Ln6tElgcVPh7qj5JSS0/oJG2cVhOE0n
2LSAqseRGWyJSOO3eLNCLWZ1R/nWpodLr4eX9CgW0u6In7hHwYUtZ8mQ82LGNzyZ
dwOwKHOteBEVRa3bZB3+7+3LotR0hGx3IytN7pnk/CdYsbLUeLpdZuGr6VHmmTh/
oRtgm4/cm9vvDg151b/gBHFJoBQ48wo+PFuoUnTkEhD7JKj2W/ziz0QkVg1c+4WZ
xybdjK3XvzpmKSo97Gh+i1PPoIN6scGxc3lAPkVRNxdaQNPzwysS3hzPXnX9CjAN
7W12sxwkP42xIDyHuFqog6TBcVkH1ssTtKqaX9kfA8tsX36qai3VU13OgvsLHUqi
BE08zbTUmpZU9asftzwO8UNjH4bWik968wIrSK3el+++14dMaHnCF9aSTYcXLQt/
9Hj4knU9ISp+KIsMNArqMxi3+LF+R53gLKdc31txaKsosXuJEvgcLkB8jBFrM3wS
8uwx/Ct22b2idiEPGek8NMcU1KzBPZX73A6R1BcvGghJkufK9+ZcUhIp9ItT8FGy
XRgVwIBIhEFcTTqG0pzGJMRQtlF7vvGKmXMshl58VIeJLvXW9dSc7Z0A381f7R8P
CAjRJyI/B1MS7LjaaP+QAKxpa3FfD6lVLgHRrIUaFhiogrYlVMs2dcxQudS6lzRd
bWby3A1m97IKXDpLBUKVDj9ZfxhWrFaL4tUPmREQvdTRkojotndbRAPpzu11rAud
mCOaD7eCQhoeZaUTAowyFr86Ci8q3HSNS3BHAc5ScZkg+Tg9Oy/hH4JxRtCqxgL/
vEtqPPOpPvcyukJHOfRLl4V8ee94umKcHW1ink0DTuovix6+T8uFOg9gEcoMiX0m
5lwk9keh+PEiwhBVvLQHqwhW1inpyBop44Cf3YIHQspavXuOqcQrVouk6WA6KFO0
v19TSDYJ1y6T+FMDaDjxr8cxR0MUthR5oMfQwnXpaqHugnpfvPb+fDo1NxR4+T/D
wbgAlF53pvLVoAE5Nwj0cF4Dg/+trSBYjd6jv2Sm47vXE/yokVvUsIiqhN86jP+x
FbSvZnHNW5RRkDegLLhLFv8g++NbLZe0nYEpVYqqqlZiPxbocGuBMeM5Th+ZABA7
hY2KVogXwXKzv+KLWdwyfspqDHbMDgI7oxITzXwP3ektfX0+QG4zaXoqPaitqdAp
kIMeVYtQpXndbhx89bzqoYTUguoewkyGfnATOKRtVlxwYlGgL/BjE8wgSiLgWBjS
3RJRQgEOiI8SixRq3b9YlullcemAaq7oFMTJUjJ9G6+xq1ouZNNcBrrp/Y94y7iY
FjXQ4Jm54YFCysg94/jBAESL2N71hOYdtFxf6zZrSXZeMhi+/SUhBEcXVdMryCHa
AnQFfs3C5iMo1cw1LL2lvezdE7SZuIsRwAt/cTZF7HHCgeM0hEqwj4EAgnbAYBi9
j6aTifNqdXDXAaMpEg3/XDHqm1mw1F+sQbcHLSiuMFF4BlgbXF00QvkYbrpadcPH
aJvkCKHae1s65UJtT/aNLYA+Y57g/2ehiCiYLmi3OFZG7NFW8eNZLf3f3sM9bjlI
eFAQsjwJfvcv0J2w4TJeEVd0P9NA8TVFvH3cLih7260+aZi5GSMxI/7kgHsLWR44
jgEjkRkPdaSuegX+Go7xn/x4ORH27nw057rIvzTau/Ca99o6S4stNfOa1dUBxTaH
peIcizjfVnama/+ICK95fvrp3G5yJQ8+6HvL8MaUI0UohELQ2OhnWLsnDSJR0JjX
xt0EPXGRrhL2EUAa8/cCRbsst2RiJ1nSKyaS+IFNlehSHW3He3zgN3p16XQj/O8o
IwzeS/2Q32hiPOzoMOINwjZVAVQLP+Jg8jCjCE/nSvX8bfprpe54c5qIoAWSRC2G
0m33QHpMoyQhcT6iDWp+6xuZ8apHSwoCpOXYyDZaVAmM2iqXOHmjup7pn0bYWAqA
1Riw7beN63dpDNvOwK+JdzDMCRcgz8zWa6U+lQ8004nAZGAZFkbM34QD3JSTgRK6
wagr/5j3LXC4ZaR5ERUw2x58haCvGH9IeigSatMgbuuEBuaI8TLrnUr2auCFGi1/
hGc6tJF8uFJMj1n4Siy/cf7Lo3k9KQm1rIjuCYhneXIJESmi1YnG+R9BXWIU0WaF
0zxAKRjx914dAjpslaCeVl5ikpt34KbUK5Lu9o4L8Qqly+a6Ovube+7i3HkWvMmW
DENSARa/HfO83n4LAg4Dz+qAtpsi1UZSEwVSem4rTzVMad7crJawkPIv13OsY2zB
tD3aUmq079CKK1wO33Dn91WxOrTCF0PQsuoU4R2vT0QSWkQ7VXcRNs6TqgR76TSc
CtCZfdo3cKLkJQS83t6DuJ6CY7cnFFhTLkhhRQXZYNKM0MVGM4iLhMoV+ebvKz8F
PkFU/m04qLXOndMfxWd1YURsE/EM+VEAKfVW60B/rGHNO4BXvD8JnvZ7NMC8cY+d
Y7bzH0DWeNDvBlAypAqBryxfwFv1EKbuQHAMH7kXWDMyKyn34+LCTOnQZNIuq1HI
oQwscFTNBfiOTx3eo8s9CtgnWng3X5cxYP15/qqoXKQHPWVYYrGuc5hNycR/1z4B
xWQ9uhYGTDFkMMqKcZmh2tMis3/gTcdo9EdKjGbDcg2TnTay30G3gSAYk6MVqUZA
RDUZmLRIpBl7nGzXkYblaxIYVh2Y/qxT05NixWarT0Q2+U1S/0ElrcBzGYqVKzMR
aclEjUkYPlTRanIflRhPnHTwwqWRbTTeaVdR14I3sU3LLaIR3y7QHQA7Aw7NmCrE
WuxEQhK1VrQcnVg+ucZ4xmhOLUS8wBOnARLvJ+NK28MIOUKOpZD8yMAkYqvncDxQ
SfvaSINfp+O5UGJ0LRIfULvfsoRWdtjp/rtsi7ql7IVeZeflHMkxpGCR6rNeZrW5
iI96bIfQPPO8TivN8ox/r1EKjz8A5oLNGnkSKh0aPn/2EDrXaxDg5LxEIKiUVU84
nbLgEkW1y2utkY5K1xEydAB0cqKSLQfnqim3ul7+zGRCKpvAzx9GwBdHuCmkebAI
shmlqGUKbK427lGY9BHhrsG/c3att6pTk3W3jDE7pqjajACpgcBqicASibts6x+1
NiKj9LrWODng420SVsTB7+fu+9ERLS4V5hnIVk9RQVdb0W/4GmxSvfGbQkznhfb3
ZoWw0zlRCJm2r0FyAi+qn8eIX/MwDy8wv073vX2ay9slxEYUnmpwtz7B9mN5cqyB
A5oPUfnhH8QWgdqPgDDoJwZViG9m6OIJ97oqezE6c8PZItF5JaCvhRXZRI8L+eJo
Hu83luNFeKBpdr6IC9ZlLAhPFUpk6OU0G5BpvJePWt/IIuigl74kS4dE4c9XuG1R
X8gZ/qxeNo/Wuhvq7Ef4lnaFFb6PH4efJjpVQpJevAb6QoOiOAmh+YS9Ch1Ns25X
nfeQzIqnEc3I59h4Qaz2LYFLEkier2Oknylet7BhpbV1G7Be2/kNrwG9dyfp1Cc3
DHRTUKE4hmZIy/eKEftYV7vIwU4h2RYrPMpi9vizppRQx4WdyaVLapCLHxwHlR2T
ArZS7Ey20Lt7i5jMoeo/loeQRkMoO8CedbOLP/G+ncNxRm63J1EfJApUUBcSpHEK
uXVGTGlttGHyKewLVIsCQhnUCXxAol8MVPXCqNoh2At4+CHK4aBMeaMcZvsUUYbB
r2vj5bSouyh6dZdJKVOhZ0AeR8ViY9acCVTRbB1dVoDWw0qmOxQOSuhJhimadgGA
ZIQWELdw1lTwfsRdH3oCN+00fumwxCsm0bLUjM/A0zJ3w9Qtns3WZ2yJLcjuJzl4
1oh86dFM/oGYfeoVHz3N2pFBsoSMVNkvZMlaxhTR5y7EP54ftGU7eOhx+N0iedXu
eRQxzMPWbbH1ZQmuScbm2YtCkua6gvjckt4ukEUil1KVUgAjjhbbPQewZZbPfW5V
6zzoQMUlNHF+3FN1GEJ5Rcez37d/nnLY8ACcpo+QZ4bLGIiaYVfA3zHEYd4mz0Iz
QecVQHbBsPaUZamVkrG0mWoB77Zk/EgMUw0pocVZFwWnjuz/X0iTTtgWgJPUHmyv
qgIxkRq1bgPidQ2hmOjVoRXEiImhEfMqqwmjMygLUbszurvy4PHvF0mSNeXXjItP
10VBsYZ1ugDuhGMpnOohDVWkC8R01unZyfE1jUOVh1D4EdbAMXgpQWD8EMiEp6yd
DEVzWLSYP+wOj21PMZcHPz3Vo2XqQeRM3nJlpPBOvuqOMtlBGPZ9gi7jq5O2AeMm
zUeKHzQSK2GWfnt2LEs3vABt1dUmU6z2D9a0NRN5+wAIP8qfBF0qIzPMRYdryt+g
IJb2eG8vnPpVtwJB59F6aSK0S4/YWtVktnhlltNA6d+cm29k4DC9oE3+1Oxt2Mr0
BTJsYHSrUfok8rxmwDDc2ehPuRUp9oiDFEtPFiyuIz9q3+Yw94yJ9wEPKSq5gdRM
0QUsBERtGoid8qhpsdQiZ28GeVZHTMa2MK0Gk76iPfAzGObVa2H+EaASHFht0xYM
k/j53THWea5rJADbYbdDXOmL1BWXrv4hXq09CKYXV1ZNPnLkLCeJL7RTPKPRj1ru
fEjqf1NlrRiSAOEZucH3FsVzlJZYXjoOk0ozgHPYmXcymFfIssTCom0Ge/5uFsgY
yR+nCWzEPwjc3LIxpjktBHCtQlvhZUUxKrMokT+MeW3lGJgyaVNhwp9SXW1vKfZi
MzNzeBcOGnynyGoUoDdHhf3BoVKpo44jNLTDMzotifk5XdAWqtLo/RdaR8kFAf2j
aITY1ZAzloiSU76eMXRCtDbUO6sC5DAoNe529ihEY5hYqA5ueSID6qzeQkN2MWY8
f9SOshZ8b3Bpb2UcujCHws+jiUuA5Fg/0CLcHI+GTKlzwVKBzmGtlcMcTqiSDaoo
KoSSHUgllkZLz1mn+jx5wSiNtrJBQ0jYVhrpS6es+gr66VWNCEvukRVmUFOAijCO
HgsC++AgRd3rGUIiGp2snPo97xhBZBc4yiIK2DDvUhM4GOat1vonL2Q4R0imSB7d
jZyynqZBJxJFxMxMrsbGpXkUefsJw2nuvoJ16/ybaewlEF7PeOdYF59xRR6FXI/w
akjSifpkHco82mAvP2PMFEwRUK9vC5qBuROrkE5cD01LmBRsiTZqEYsL04iC0IWu
rDdnQPF2d+bYLgFLuOo8Iq2OWEKEHRXht87Amkra8S01rykhCVfbFgsIjBdr7GNF
xn5owijei3D5TOBViM2XWRrsoXuSM+PFdPVKyrzCe/zMr5yiycwYtzBD4M5BtJVz
9agWop3QNbfQLv8A86PgXPQHDG25f1CMmIu66zhj34xFVreQ6WgekrNjx1uUJbc1
5oSLv3Sv9rvQoC2IFBoNgJy8oy299B+qc+Yx+RbdELvTjBEuA2cbNP2in4vyDQiR
y7LTfT8J8G9a/ODBcBk5A6CMNzJqBxYdNRw+Iv5awqHbYNOseapoZae2nssquosO
R4X+BnXZ8BYcxyy2pX9PHevvnjvqOvRlLOuXCP7gc9WYSowaL3m+boApQRT1mr6F
ziyzy1pG2jH/6rLhjJ42vBlJreOZNOmNM4zluTcBeZgi3TqHy1ANH8sZ8z6FHlDD
GY5lXLcF/ieb4mCxUWgY4FeU/Mod7IthzoHudajmgesPLr4ZCpfSl0FOINCOkE4Q
Qg1YmJbY3vixXawyQJB7W0iTgjWl4AgobYytiOMJ+v2Yw2hxExE2yUshsFT3dAEh
l81dmzyJGMbI25KkEEiqSLYtEAZZuhDGac5Q7iwzA+xEEisEPg9RJqUgs2s22ZEJ
oflbs9Te89cEOe1BJdeuRAUzLxxtHGprOb4Gz0pRDtQg7g1nqH9naw+XNgabaWsS
56hd112JbCDZB/u7l/y/QzRxOGAox/e8sWWAlBadBeTUgr8q3aZsShhvsIG1jT6x
sYDS/LKVMCrKgN2im95Q23UAnjerEX+/BC6ooQNE5QxsFHaS5NmgszyPwYAwmgCX
pM9dRcVfqGDOM9ZAhB93/5OAbvDyWHClhZ5LmQ91RmxB/LUD0corpss3ipiK0q6a
eduewn9fAP75IgdHEA4kJe0kNYZFrRlgsXdFZVlQ4IbBWV6HnCVxQlYUCyDALhz/
M3gMYj7OJbt7U4Y+w2Lm60OroWyhlz8DyQQ/Ud+cnlgnenW1oLIREBygxjDcyIae
pq/Ab2p62LJbJMh8+KM0syJdF+MCv9OvvR7r/KqcNCSgPRfw3MdsudIH/dy0UwUP
jPMdvn3NZuC6GGIT5WM0KXHbjCei9/EWBftDU/0U9vJR/pKZ7A/jQt6fRnPl1Zur
NdogHeTPSV59eERxMkN5nx1/FjT0ZSRbpnzjnlXhcuP7uHXYIjWTbvGuBTb4Rgx9
o0K1Ijz+Cq6yRG5io4P4alnzazhQa6QKb+muo33+SEA1SFhHfQ+4d3yy1CJ0URTY
cx5HbFR/D1THkvxUP0XduHPiTfl3xQ0MWivcm6sX5mdpHNYB9TDazzfwlNzUa/+u
jT4aYjb2aW1uf5MA73PXYdjTnsAP0sRl1Lg0RFkNelkPLtOzgD4BaHdtyzMRndAZ
nVDZmCOD7ls4t6BHzXOSPa1IGqz994WrJgu1M0LztM2gHmGP9UnRvfcH0ZRFitNo
l3Zvs0J9en3xhKpHJXFJOBQrJuvGNxfXFzI8X2cARLkr2HVMd7PE6HgRwkmqzJ7c
XLaomXsEk/joL/BaaXMioefX4t/eK7BdEnzfNFXJV78YZAg7K6krmO54lIEED8iZ
sDAzVw/C4xxJ0lecPprRTq9MvholvSw9Adq5WOQaPgm938inpQHzZZ0FhdzCvomv
vLsa3YwW3a1nTmuM2AdODE4ftY7rv1tcVdv5PLsXR5+qiFI3WHAynkeG9FwV9SBt
lNr7Ga+gYoL/9b5rZ4B+RY/ACPGBcd5hk8dqd0JvDmNax8q8gAdP9PXym0A1JHTC
UJDb58zlxdRy2nRYF6Z9kCfwES+ACs6l3f8i0YG/F843SfDtp4kkjIq7Dcw0Wk9F
LS95iS8/NYK5wWEI/OdN0zq63sJ7AjWsgyQ5OVyCZqn+fNkwhOKTPbn0rV/UQFgi
05imkUO20RRx69WsT+6JIYYHOz8sV5TkTwANfiZNzqIYALOZr5Tu63F5B4bAZZqx
ud4e5KZoSVONadSNqsaLg4gI+EImS7fx8GM7N+lZMzjTPBCTZ9qkZV630AQYVqU9
3/uE23AQ8AkHmqQb91AgRPOVdNuz+oD1jupAoJvnaEScmiafKT7GrC6VKs7/6ld6
6ue0XpLJMZacGjlgbJTkOTcDC0A1058iRTjp46cNwll+9whyaikpgEASMdTVcDZ7
nDaMGvhWVsPwB4BJq7wBCKrQclczFk6+Q4LPz/ZuT1xDWcVcJC4AuKRV7vykT71o
jwa8DW2yF22vnyTakTdN8YXB6cxxtLGOdJs5YarvWOHCKTeGng8mDjd1+ig/lOun
PGM+6gExgwpLPARM3ySXmi/kzZ76Ljrk8XPfKepZVbKzttTtsWuwY7OfK3TthC5f
0tSWwNF1qX7xfLO9lSNDBZ2Kg+ddANUYazcJccs+eEfn8S/wDEJ8HboTvD8I8dct
CG5hBigfXdWwD9ldhjaXy7OCirsihgnY5kU/oYJdgr7yCXMYE/I4uQfYFWjmjvkF
Oge9cMCYTQxTnjEp8SAK2ZdDN7m4dligHk1W1l9Ku9Wo5PPx9CrQYwLQGefnmquc
Gxwt0zED0lXj5alIaI299ie1pXG4BcZi/k+5qPtY2ZknSnMM4G9QsAPuJSJtp7ki
IRF0y1NRCgrJ6t1ymAsFD5Wh6cl4KrKOEo54q34XnXsH2Zi0Xiw61pZb/wNYezw3
AVHu7fXFfsB+mDoffL2EorIPesz+xFqVdfeCdF3bRCoqaBPI1+xIKxK411ZD4zTY
tzdB8iAJaoWCQnLluVNkey/kMBAr/u0v/ePLA0ZX0IsdqZoM7f3HJotW8CLLlWRB
efiV9Ys6aknTulIyjq3uqnr2HibMYX55dCUCAVR8thGSqU0XvkbjE+fH8RRfkQpJ
HMlkf1hPq2Wymi3XB8hxI1Clz1i6Tko4N+wOTo0zhML2utzQZUa9KkSGGOgU2fzi
hB+rA3o6qP+NPrrvRWDN8Iq7WMqGxJlx/o/CZKHs2Tueg9Ioak8RZ1UWDG001p9H
Tokfuh6fBNss4N+7g7mUHyqawwxrH6nlYRd8x3aUI/1abqdzapV3vAjj+yYlq4Aj
rODal75SQS72X4fu1V6FAAbLCWD6WOIWByvKE2Cd45L34blntEfkDf4NqfQjQdNY
mdqGm96zeRoa27guFXHVZQtf8VGmVtSP6J6H5NEUBUvZQX5Yag0s+rPgZfbgd3x2
2F1IAkDMUstssTpQhmvjmo+DyV0QC8NdUdCmm6bt7EKwW9wWskazZRlZeSOFVQBe
Xfpk08XscUIeiriTBYdbgKh0j/PzzV9HWqPhalBDMz0xq8dMjxLTsnX2YSw5aKLw
7n4jZIiC/tJto08odEaW+YtnZsO77KX0VV6TSk3VcwxJo8RvqOsa/bNXTUBHvJFd
3RBgmcX5CubNfc+9x7fdT8t6AQPvI2I71/+gcNVRYCDR3lXP3oGz2ReFuL7j0FNl
Ulzt7ljiGRFdPfR3CpJf9moO9utHSWaZbVSeNZ0rmu4+tc0IMo5Rf5WrjJ7HdRd6
eXqop2CvpGhKen1buQQ5KPYqW+zuBgNCPuY6pVHDKRcQVG2Fhp6OdN85FnsTTzuS
nsoWJffok8XzMNhKQ3WESVS1iRQ/kNzUdLc4gutUS6bWLLOV5CmHkoPsbPki0CRq
5mfSHO83wyZ5NvNUojRholbFpQhlLx1p9hl9jyq10qyWkm8pZkhWI6MQXwx3Kjmb
jEObJcJ9ByRO+vW8HbAnmRjUONRAzIgTdapXlG/tXRSF922BK/1Rk1+LBwjPgXfC
qzwr70iCkw92LC99aBs+XWD3FJgxlm2tI9nBunV1x4VriNTKyR0hLq53BbynRTFB
wwq5gxcLg650XsYNj2y6XqKqEboQxOxaxUK1+5AbpHt/zAfvk0dPvxjhGH35laZB
fybgLSgqVH73/lw4nyd22a2q7BxIXA8ED4Rf6Hr7Ich1phgS9KmC/xiiK6D6eMVh
z+RlkCKVECwmS/oddiIjOCrTmeKtP1v2OG6yzjI00uh/Y6sn6T+IIKuEtAALh2Nl
plw8aKsSRNBAynTKh+Kog9vmUqDKgQf5i2/vZJ5IoeVOEz04u/KyvGgS1SVgPWjH
VBC2D/4maxwf6HdwI2fGGWqQgGTnCKiC4EoZ1HmAES1yv70wacs4tQxa6qcfNUUd
f4zgTvyQgtsF1uMLq9psDLAdFh1GyNFHQPVHdkl7+FVyutJOHFFXngBTrS8glqb6
Wq1+dyrPzcNQl+Ou5m+JOtpzeV2MfJlOB15cy9kK7qJ123msYZSuKLFqk2t5zq8L
7fpvzbtju4zXVzKpKy8zx60V+Dg+pryfEEm8vD1BB1xl5+MTow6reY4sLDiAtO7f
8ZmolQXMT8BvbhKqpo7W2Lua9jJWK50c3YvaPq5XNGgTtQXRBb5e78wfaKUZsPfM
5HMdjVmwVRUmxPZ/ZyFxhitU7iX1ivfwOSuFV0DcYY8X5fw5JT5BbhGkJoY7AAAs
1sVVs2cHCGUDgkJG4a2ppKSP6cQcHNXEtsTaUO45DywU/w4f40HXxAQvqoLPfCQB
AsIhAm6ZXVMMSBcVlC+R76dniTHqNqMpQNoNLpLQGkYf/j+A1IBt4z6FvBO1IEmy
jeKkxxghgiak8rYrJYBujdR9amGjV2UggvIEcR5q30cxGYZy1Zg5KrWGiooHRHRj
6xnk3aorHL5YAQ5g6JyMRupsnfaiLVj0ZephU4F6XA29LIrs/bXAZEsf7Oph3dsc
GKYeopZSqFHuyGWVZiHbwCZAxI/u6V/o6QS9ybYmydaZsg3s9VSENG9C30C0pf2s
NOTYHn0CAInoZQcPBWflYQLhYZ8TE2EYqPOOeOg4IZ1usfeSOrzCgdDhPl8Czs68
symYiZcSIMTKaDgKFUGmOyhdeSCeXjL3B7lamz1zIRF9UPBHlvUywKWKKkf5zzDs
ZDoktw+3N1PnC61ny3SC1P6oZ/DrsbBlBPX1VjGLIG4cFUQLoS0w1yBsPD2nwCB+
/294TtklZM9nmGjX5q4RQRgZjuBUUnAQ5i1Fl0rom5U/PbjgMQeM5biSaBSsjy1r
plKll/BoYESDwmvHRpEe3P6QQNnrDumqakW1BvP3IGn+Rmc1xcLURMjAa4G+1anx
fFsGihekWJ4YUlJV6fdwlBmPm4znMWLDM2dwuwmdLQSAZhE2mQQvSHhMu367zYC2
5Q/L4bZqcD0kplOEVDac1Wb3Gbt4aVuqCMr0ZQEy4cfFvPGlTUdV9ZTB3eiorrEp
MA5feBNpzV/38Eo4E7j7s+HqX44zLG1ojRDtRJKQLcY4oiSk6vZcoVFS4MkU6q76
f+tM1bMdJB1mpHN/TfjJYMOmiltFaLHLofwCSZrC9/uy0mTNjleHWorgrtnjPnWQ
Ld2sYqdQq7NhXFj8eAZ5Ma+9ySwvoWIUL/hfVgtBRAyY/Tvf4s1mx3m2BWRopXzY
uXo4AJcpyJwWte0SqpWVjJVpeplqS8MUFKzaDVKsqAyL2nFwROnR2DUZJI9/e2xH
tGdvzsFFxf4fO4+HlAsjfva51BJxmSLnGej/T/vEjmtMhkHXCyB/QlqWWGRPcEgN
VJSWPd16o9fGULwm8yu9EKXfGraP99++vBXqZ3YXnZJO0ZavINYzbjDovBDdZY2c
5keHka51DfaFKdw9tih31t60KtNAkLj2HlO/xYHAg+h1gbeEkRB9YVw60zUDrL6k
oSG5iD/Tqk6eipE/yazAsvaM1HxvyenZYyk7+v+EHCJt7xd4bq61tm5Kgu0NeTr+
gE7kRW4eVzVJ5CY5X9dXuCpzlwF+stbANGBQ1zMBD1MClY9sSCzhxqkV7gOA+C0L
zu2shiPJVQcPDvLWKbSIOJQczyOVf5REOIe6cs0ase0n1g6LkJedgW5vmd6nvN1n
v2oXew/Vy/Yzt4D5LFIZ8DFkTETJdkwXvf1iqkxPsBhmsMU3vk9wvHv9w6TPBHFb
8C1ccYMwbDlXM+puB+yYmI+yzOaMUDLe7wn/IGtwW5HRwOy8XcCuXjLMf1JRJOBn
BDsswEGjNpBdHI2N/m63b9ehuiw8YKyQzNIEWMY5KSjzd0g56xNTZ5Ejrn9Fmpxe
NYWgCta8emT7CUj2dtsalG1eQOM3MOxj7X4Fj26gV8kKZplWda+ovfMhmjGT3sPK
3szmXx5A7SAds6nubxtBPFprq24Fjkpk9kRF4qmbcvQR2AIdKcIRHzN9oPqlBnkj
WC9h04D/zFK6BJwh+51lDaQqfgPXyS06drx6jK/fM3hJuJEqLevx0vyka6Gvzz8b
aTzs8ZBMQLgP9I/2nXHoeZ80+E5eYRnrYiq1gBqpZHsVZK8OvILkEKjwdIvj54YN
12gleufqJ3Y4MFhD1qXG5I20lIdKBrujnkEcFPaASlkrdJGN7quIgMl2qiw5NfKk
k1U9VtYzk51F6gHdTXLMZBWlzRhXeaofwTGWlxGn6jac84ngG347/qFClTZ1wo9N
ynJQYBdE3OnvQ1ZgxtSADG2X9mfEplCewT6XmyyH+nfPiXIZ6nnbykVOpSvajPPi
gxIgnnSOPWEayT9mTgj5StxGNT/njtX6bntykaj6ZAj9sGXiyQJEkvH7udy22uwr
YNMiUYlls2MATqRoIYrwYGV3UBNPFEv3sh/Id9S8Mn/qfyH9PzTrz9BZRcwhYlk0
ufy2WVG6z/IM1tZpJK6jS8bnssEbNHGAX+D6znGXbdgZk8ajd1z95o3MGlo60mb/
L51BEcyeWSwxib3Apzh1Fl0iTkHjLSBob0pg+Ns62KK3U580yW802n6HPW90IGq3
EBobQq4p7JgtLzXiu1x2ZLlkuWIHOgbVsJPiQsUxyusSgUrwUJR/NrKPam55gdov
IlFWzQVf5heruogU966ET3mYYD4FldZBK8QqxE2wBAN8t+1i1frNHz64pSL4PG8e
rtQKZisavuLrLwDODfqkipDSqOj8IXLFfexcgQ66sw2AveSFOAPw6fiIIQjvWUwV
R3aUKyrC4EuQRkT2VuMa54xzzPl0DKLvAnkFnmGKd8ke6eggfxatdlZvOgBSC3er
O+uGpucmE8SDqJ/8eQlxAPPqSO5uHzPjCgfpZe+GuwF1iaZk2g6OL6GmheiNZnKv
RX439KNvEZbm5vnsGvljMQH62BAZoaWX0m7pKluptQ48oy8TiDprwkxspMn5Iy+I
hko2R1BuLgXOuj84Oq5RmLIep87VYc92ZsIOeaHd0+vLxzEvaxmlnTjXUisROImY
fua3qkrUSTLR1zbwXL1eEcp2dtT5Fu5LaLisXGTKurrnMorA5c+DYuj/GrBOBIQp
BepHT2ufb6pusV2XNvSsW25GCReiy3eX1s1UhDtupJYr699jHZknexG4pgwbPE+b
YVNJ2YqwUy+TkeoigLEL5xBIvClIttjiT7KAO+2QvbGFpHRchDNdGunMzNh7XNPr
sYx7OvUAaI3vkzjTtxf7E2XrLohNcUalR/156gE/CWzVapG7zAuwZXkep36Zt937
XYWOLuNLMDDOH6Li6I+TU6LPS2AmRCLI/srsYcSCA3hkyyxZQN7GyktwvYtjbyNi
rWWOGpZmaoHdmJrGJXXaoRTFgkAOrHaN2NTlpKlrnsx+0krt0elshj1n6Jx+0CL6
850NdZSbyZoCF8OpmTleYC2haDPwdRrRubrILYAlfS4NEKQ5wP+Dsm+nQbeP7sy5
+w5NC4TVTDs0Ln0++s014cHqsURyawFqr61gpZWV9JiDXQ4Q1E8ZzfA5KEOQXRCl
THD50/MWey9L7EcZoW7akWsQ35hWyTL9+dNFd8psAn8Xoy7C3PJEJakZfJ+w6SLD
+LnkAfK47JVtMKupgeQ3c+16+qBiPzYPR0K2DlMdnDKdOMDJ1B4bOHUGmtb/yV4f
zmxghC2DwKMFICs3r3QY9oF6yIYX/L059ybch4hBwucshoD1T7Cu2BXZntxc/pIN
nnNMOgfIs9iWHXlBFh1/eLgCVkcskQcm55QbH8aczKD1spycLlKxYwUeK8XsmUMk
JUj1idLmEHVzvBqA25ZnVGRg1XnAi0ZwIb71EVAGd/VtLaeFj9iwGgnasH3RuzU+
sZdcNnyNy8NZPOFx25WUJxgA/vhbg1AkVSUM5tXAowXDiYt2TQq4uTG4CfRGYVKw
t7DObPHbSRUMCayvgUS6f+/+QY+0JLfWahJfOeby+wPK/+H6G3k9Mfhyj5il8vhR
NMalCGEKIprIIUHn/BXhzGaK+rOwNrtmjknRxwkXVBWM6S/WjhmH6wOfMT3XuIW4
iRuS8Tdvl9o7iQ3Jgn201jpwFW/FqfEPpt7kTm8AWSLDWsjVE4KhpFhkB4XL4qaB
jCWcKuJsakC+UzgHlfl6WQUMMcT2STW/L6XI/byBGfXAQ6mQUEHlaeBIsma+s2Tl
odJmTkgHyhnbinRyueb5cGhQ/OFxzOejZYnZFid8hnVGOeNvCGz9dllX/70MMirO
19mpXRqEohUB8njoe90zn8440wS5hKzHwILn1mJ7LunhpFS5dgu9U0HspVz0wCFD
MTQXzU8sKzqRnwE6SrUtpdK6GC2vDJZMdIESbrGIOpwEMhRnzzXLC0stxSHCoyr0
wfNgiW4nG71h8R7ocSaTvyocHwW6qGmZt69RLGAjclTJ2RFCA+yR8H8hh5SaZzX1
2y5OczszkwvdnznXeePEALosqaq2tnrl1dWAx/KV9WS2g9zBbmXKakGt4VZK3bSG
aGVk5D140E6qai4eXFdIVvL2bL+ht7Lyj5nxd5QOn/v0SB9NjKfXJVXh+JDglVzp
ITMOWf7wVTWBP9zfcfZfYtb0jBQfnUD17ZcTLmhxnqR3+OaEhY3uuY106hZfD8We
5ByCkM/5yVJZOYq72JFM4eUTKclQMSY/p7iPhoEVT85i1enOJTRhjjAC05luLxWw
jXG56kbhH+D8c6K2o0V2i6K/zR7Lz49fuAtRq/+1URwdAej2DU1P9VBTIa3ZyBUs
84Oe0dsflO9Dz6Id9f3yh5vNYUfZid8KBBNirW38PaKRVPpaIerI43ZKHrEffSjI
amviiYfeMLM1BJaKBBWoSFA7QxgRBkCggBaMNaYU6rYvy0o0smr1T3PiygwBAc9K
OEIjH5FY8PIk14R3Imfu3ImPGM//dDBGZmH9dNkE/9pWMOeqUz0iyF5SvFnJmB/V
qlosmV8xNGJurbB6aVlEBinow4jUofAJ3SPenoOzVSTgFfXgEMN8vfB+Mg+J+18N
UdHZSl9tarC2eqB016zk/WkdDsdjDYrNr+9NDyUxPwmcyHwvM0YWA3pGqMwAtrcq
tO49PrKay7dIBgC7+FvrIYOw9J+JaMuTTsf7zaxpPxrq8iCfnLWDXmpzC4B4e76u
VqLMVlQXxHcvU/vEXQFvaasyaZsRqCHXjwtoUW7M+wXOh6G/3SjYvas2CJuRrIPu
UnbwBnGFyA8j6jbQ6OdDSpe0yO+eFTZ3DAgZE7FWckL/xpWztEVT8hThSBKrfh57
xo08Ld7tz/S6szGs4hAw99yHDBG2GRIOsHRWSNR+IbiyEH6r2E/E5K+0Ql0LfnnD
wj9A61l+KIaGAdgNJQjafomRdSkbEisyABQqEKyyOXr/gW2oel0i7Vd2R448h7qz
09Kp+Q3klXqvzISazqNbN0Ex9FOSlM1aBduuAJsIRbP7oqHQcfsVehKmfMfmwlmn
1euInqWkUyHiwY/lmgci4R3/i4+giSVKuADljjPEsHtq0vg5qSM2PSFc/RhybQzz
yMAOcaS23Y2xbPAOuwQ1rHVu2FClc6jwxMFFWbawFUGy72fSy0IV13o5b64a2Lx4
BpRlQ1Niq5gzbjQgUoH/mjE59mKeB7s+anilmBmzMoT8HXWuAABiEnyyHObqe5l3
+rxzxlJYmpo3hUXyV0fMUHXz+l2f3RqlBU7T/yKHDP9OXB85SXIOk90WMiaAmr8e
3RuWJvpS+LFRJbluoUhBCIuW25z0BF0E+ByKwE0Xw4iT/gAaqNCLQ7rWFWHmdo/u
4nSdZEUiK2zNcajA4v5plU0wJ4n9JgO4EjzhMhIm7AwcQZqvCANDv0aGfAl0/dF3
Y60F4nBDRMMr+FdWa95AGqsGu0R+bKtVkC8rLnynVGriFa+feZmZuQuHrKyTia0p
ISifw4jOsTBX61stqz29GvDNENyCFfWRxWwxR3WpieSn8B1M49S0aUTk/ljIQizg
+fF8auV1De2Phs1dPRrcdZ2gxHBkUSeCuQO5reTlYF6bXoetnp0aD+TVlhVWaKeH
dwi/AKUMDgIH4U2J2FTUTJN/DSqzk2jVl7rC0thFf+5mNlSnNj4GUFbyeLSxdzzc
RdZb0WsE7lHF2LNMUuVq2eLK1QuFhgNxUZYentL3QD2m5zP1kyzr10MEGEoeq6z8
m3lfjUG0KlJEdByKeIiH4AAbscLSgAyacV2ofo1A+rB9W0R/hAkqIZRgY0J5mRRR
KA7EVcB0R/FtyMNiO3Tg/OguUkKtKeQOtkaIyjQadrNiH2nayKewfJTR32mXT4QB
5WYymMRLptFSBgPCIUAoUtboyfGLshsgba0/GVWeNliqqDKUAW6vsgUF7sI7LF2Z
FoTQdmVH2mewIM27nYfQih4zsBQRVqc+xinqXOnpn3LsbyHICAO2nmcGdax2btOK
1V00CoG8+HUWeZgeviKfr0BO+3r1qCNms7qMSiPAaCiSMn2zQMqSLz6AOWXFIKqy
EgaWBHe76PzJtaH7eXzT9TAlhaNFhzNaQyL7SfdZMUzlmaQ0S6ziSxXD+ViNzZlL
GprxJN1iQe+VwDdrkQOMnE91FrTH8DG6hWCJPE4SlxqPi0rNceSRssisZ4iJJFs7
K+oMBLjR3Ne4EMPWpr9bQQqH2O7vYJlY7+RwulN5A/kBFfPNX6ss2UF/XeH7unCy
0uq8B7Pl+2SPXfveSdGOt4N2BgKZDL+yvkIEpwS8Y15LD08i8dA00gtkoBxkJSWO
NJMybjgFVVduN8/vsOlBvcLKjS5arSeoOZTBeqcG46hT8z1ae7em2UkaLuc65MuK
mj1nDI6A+ZYDvIY9yJM8abUZ+ODSbB1dnsK41fPzSOcxcDsGCfleUywTjh5hkTe+
vz1x74RkypbF8zpW+o8WysS4PR8S9BPsmK0C1smRAFLVLBLvcowqVgplT8nVogbQ
0gje6GptaZEGRSdDvOBuVWma6L58bkN8IlZN/l7VVtw+0KKhwfjFB+MUwcKuQfFb
Ez54+OiH7MGyAQJSGIlbAXjdhE/XXMjSQglBo/4wuqF40BVG+l7yUakxfcribnAb
IXSJ4FqzHlMqcSfOo6nCTCJv72+1NmBWB3tJ0QAiwuvYjFZs4Gtqp7fgKsm7m66X
swBNriuZOvcilgXtsWdwJZhOmtCu/mxleM4x+cHUiLYpGUR+Vk9Ux8VPfAt/5im9
zhBGDPgeTEBkn1emPdxHmdIHgszykEyJLpDPxMTYHz7c53QcFJzoMNzD6EqQ3yuJ
IsrZfp+GuhIfQfMF5mRtnUKbeuwqryfF8oOBpLKXCZC1ic/NNfrMfqYtj328NkGm
1eYKg2XTl6jCSx/Zr/Oqad9pp7blLmZfYAGMieXtOh/oJ7dJnyk0+8E0GLgmxwww
8kebz9Jv5QR5qIqkE1PIRv7xi5kTJfCmvP8BHr7JbJbGUJJd8L5Gp6yH5H1p1tH6
ZP7OeQ/yuZuxuXEZUAlF7XQeXOhCH3UhVik3vvEUj70st2vPIP6f/v9m1H7zErwL
ItqpguatxeHNij5YnqbLnMPXa95Qmo8IMbPK4fTkw7RvVSrzSlDPyv8+6j9GoD5C
+LuOHIPXqQPmcwpijMszz95R2ENgOME2m/b61efLz+reiFQ6ej2Ed9qVWhzpGoAx
gYU6l/+tbKrkCp9lE3wWBYQRDQN6ubpXd26E5J73G7zcbmdRmtEvP8C4ZDHbYoxO
vvNnWaPP3duwRxiCbKUDIx6V/fCVjxRoKmWcyg4QC7JHNF88b3iOS2zAvmoj3a91
KdelvYqJeqjGhsLJYx82Wx7L7oeOIMyZbIMyz2AG/y/QmA/PJyhvM39HlkP9J6op
TygiS3OyyGNiCbfudW9q+t++au1mvpS290AbCTU4VHY3V1xSUwnH4K8DAk1oerof
gOexBQZn3fieqRafoAvKz5zofzPhUyTzKoqZANV9QPyqKA8sebJAtIs4KjTb8wfh
QTxjHP7hmMWfUi/RQSTrKmuHRy9T7w2cUqtUdBgbZPc9/FxnvmwWOBBCISSsn2mX
A8/04IJkDofUoW1nhX6dRwd4YdsoG22VAS6e5jknH1LOe+TCN1htHpXdqMK/aFgh
vpYAyePaDJ1IdPsRBdfWiTCxYrvMU2V0IFsvycUVzfniJJk6VXyllPJPymOWs7f4
SEzCx2h9Qyw4u7qC+xyzFxaly7kjTbQ1jzfmB2p69gRDKnKcS7RPrhPXXAfgg0zf
IWeRUgLkKUyU5ZDL17bSmyLiYL4B2DzKjbu2LYEXaiK14v/jq6zqoGbVJNBP/Oze
F7qKIRj/1vFWG4nHPs58ySRmys6HhrvxjDc0scoh+WyDms1xq7jkTRhSMwhg3pW9
oRz3avCHQX5HbDziQOio/qdccvprAYU4VN6wItKsXloJ34j/BYfOxeRjK/kK2mPI
MXXHnFc3OaD253mW0eKFXpbx1/yIQ5IBi/LL4fSyVuGXCVx+Ujt4D4OR24Dgjjsu
srFpogaU2sxmoFEdhwpWrzm3fbcSujUfiTniDzIHQEnql+kaAbbi9G1TyN788Mkg
5mHB3DVGny04OgTGTTi5ofvrpONhFzoHD4BcFCtNS28tmzJIonvOhZWgXlfCp68R
uwx9qN09hEkhWefiuKQ6AFN2oWdZwOaiLEOT5OuM3ERmaum3Pvx9L8SOr7usE06f
EHg3gTsOsq/vH525GI1zyaaTYp1z8Gpda2y22D7Wr45XRb9TJiS/fg7zEE0eMSLZ
59afRIwk3lvK5okD92Z/CoEH12h4mDYD6bBArwq/SkvNmjvwUD4Crbgrvh0PCyeQ
LCOYdKDwcSLgMcuzdTrBR6vEMo2FruFakU/dpfHNwxbPmn6g1OJ5FVNC3U4gVjrG
ACykRybE6kYWJBbqDm/Q99iHTdSg+gut3ESYJ1Bre2TtJzTmHuhmxgph43aUfJQB
nctQ0o7zsNU+D6FDjg+JyxrM5UbXAO9DSdI4eGfUz/WFUH0aXSGtkVcaUfWXJZNa
EGGWKvuLnvlI8t2Jc3rp54x2cXJ5vKPPGEiWfQz9l5EgfFWKCblf1MrkAA6uVv7M
GvuM4+VUtBL2pjDPoUeQZOqCppEa/uHMf3YRQYnaUPwP46X9W6x+/nqwEI9wdR0O
Jy6T7Vyhr+HI41MeSK6ZYb40voMPY/ntFtJEkhk+XvNBc2fxb7NByzqp9r7WK2k0
HSRY3Tx3lAgzXz3TKffvWb1kVQ+CEeZ2+GHaBS8zYJ49gn1rhN+WORlb/Ds+GOJx
q8ZFJZiQUhntd9+p84SlYhwu7+bP96FGuSRMjp1FUkKGLP0lRfGzik7C2S0CifGV
9fOrv/V9uNGJbbs8GnnsiWsjbRNo2AivdhqjfuZomiTkNDGshipYlh58cl3Vuz7u
XoruzPZiw3nQuJ32C6xqfF/cT8I9rDtd+ege1mTGu+PBXH3dpVkUN63JUxj+LIye
3meZsjj5kNaovamXktthlYumSv5s/CLY7B+5gWfnPL/+RNj9aBvDlDF6W/KdTQd/
9pLBT+wkcBsTMpeVxjb9a8V24FGI+UyEp+kfRzoJ6itZDky+/wHGoJkxvXENCcEc
Ozb4/cfkfIgSURErKCqZKt7ThnC9pvOkQJdAcl06jsTZsO5w04u3sEoU6HcbrUsg
WCR1aaNziG7ajOlVMsX+vhCe+IlFUAy427UXIu6t+3pxiUvi+fAPevo7lgFlsWce
PeSKg93ojLPaqj3TkJrsHqU7NtZJtoIBvESnAXq13zIttletJ8XupIR8rFoR+Yt4
8mAp5S9ZgRs7mLghaTAY8FC1+oA09Iv/jYGOtUXv7uPg6rMWnrnCnUocOdrRwONL
ywCnAImxx80DELn4AOqx95t+weqAzn18OQqLt/Pa3Pq10XKZfcgVATKx9bURegy3
V47uIGCXXuLvbeI2I9+sRlrKqEYGwaaRpeJNXhTK1uHPsSXZ3C9kwbkuc2sUy+Tv
xvTIvjAHDgrZuXemMtfwob12kXI/nKY9rzuyrc/rOnisiZqFEWDnwE9EpfIA9ksb
KFrX9m/lkIgzVha81M1uhIsxUldLYydMfeyj+tfTzNBBHMjUds8gOdHSwOsBP/6J
IVxkgJ/pq4SlDtFbdz1UNYhAGnFCNRgFR0HVQI04TP8BDd4rVH6wE5eCriXwcPuv
xSOn3Owb3tBZhw00l50ZMbh248kt4E8vocbxrwB3YaQxDgpUE5YiOXGd1TUDuB9j
NyWE2ZDFFSdif69DnUDZdFkbpgTjG2ldVz6MVBQycAoL7BgyCXmSNdbxQFWVkGg2
9liCsJdxMGqFwNI+RcH3+QxB8fzHyqnocKaxyPNY7CSoVdpiBYJClO9IV5yNnG4J
KwujMztH5zUhEhol0wdam7lgIiJsS/cdnRl7Gr3buyz9pNLfsr49Phroq7iwd/mL
KkXECEozOBpW106KLatVB7metnxbEvzi8YV4qLu+2/5yPf23ku0cv3v8UDv3X+gf
kfNK56DflfhnUUoDjNiG5NiTc97BJ+5bot2pGB6I8a29VyiKifYTU6X/88VHIuEK
jsTYapfQNbuWfPTGaP9bzlIFNi4nTS7nWUvAHGErDEkI8mK7qBiZwU51BTziTDkt
on+hUXzV+PR7wvXg0b6WgmOggHHLVfSLvlTjXLRGvLsnrlwa4cYzs+1cR3Kes7Xl
QLYq+PB0iruj9M7uqIEEziYWli4rwFVRpDcVFhREZIEZbJQVlCVhEcZZ8ilcUx6v
s36rUNxZ/s2Yc2epb4Dv0hXg9K6x24M924Uc5lCA6C3N7QSgMbJo56+Qw451XO9i
TNGXXghU8elusugit2eN7wOw8fhEBX+Vjs7K1hAVbN+WMhGHFnBsgX807SCFmNKn
g1UU7CY9yzBbQrApj/j1bJhgOFPgl2j6arv0cP3VxkCq4Uc4sSuAHsTj7ju4gHF7
MBTtf2GFNBmMAV/pnMkXD7I9zYloG35t1xCmkwoxtzHN1ErYMXLR09PPwYX9qipc
ne/nLb48Uc5x0558YppazUnpa/Oaddebv6o8pdI9+TWR31/BFK41KinepWnREDmA
bdI3UQ5h4BM4yz2woHkE6G/PFJsBxNFy6Qv8Hfu7TSeneTRzFIZvIX3NZPKxFGPN
dC5uBTQDN8IItxj3NnfzBYrmi+gngZeKqIIXMy2iqZP1oZ+Y07ZHNggdQsMdVCIV
D8roHCZuYO0M3nK2ChJWUGMlB2wl7Gq6c9L9qBZSia1iEO0zzLrk4JdxXsqyGgKy
/m8C1F0Ftw0qVnsWwsAJnQRethRWbfs6FxntWKAvjZJMfDcPYfRam7DNY/MjJ/aH
EJx3nBggqoU8kUTs/Rn++IcD5fG1glknebECarzTUJvxL1Kmx07VVPgLVO0Vl9Wo
odqfForXnnEbK6i6z4yotCsdpjGDP1J4KF/WpluHsV9AFHF5wusKTNKzvgWpYODz
vy7NKXWNz6Dn+DzEIxacqavkN9/mScfJhAYneWlSn9relHp+lBn98/UEpNDdgfHw
JcJnwStXOW88Eqr6VDlEosCR7dKo9YcqxRTY7ff51+YM6LCaArZsXPvWbjrSh+Dg
7mzDg9SrihbMOdzwiqa257MOKuow/RGU3UsvSpkDawkD6WID6CcgxffCy+GBc9oh
XTkbFYpW04OKogikeNZE5BEAYZS7u6HN38KrURW6F0JIbawnXPMKdu1b+JCxA8uK
DWCYAJaYJxgpahtYvi91bqaINsMm0Wepe7o733gAhgNIt5Gyy9WoMYVqzNTqmXfW
NdO4rxPSAjoclBrkHD+No0/8DenN9Fr9FAYxU/Q3jWpOjOWuG0e3pC6u+50E32U2
CQAti5pm9lllIH4f/HXPuZ5bxz2z0pbagpsjIuYLKN3ihldXGHI731JBXmavAhUK
IHPcA6iwIlqabs53GwX3qK/9ae1PkgCyhqvXAFlnVPPLwitRdR0K0o11BjntBiam
Eick2LF+X9P9Xf6r/Fs9WCEZq8DdRgd3g10XE+Igo5DRMyp3oV96u++ByAGhoKHl
3E9sM6aoZnbDVgpV3QwIFy+mZOSaPNEe08EwXBswDL3PUsv8QHoKLMmQzxqklsMv
4oRD96OTmg9okVIKhJ2Rh9nxezSTGeIBExnwsACwCEFuHjEKCT11JRIV9Bib8ea2
Ex6iK9hPcqD2i+05aVWjzM+3l+f12TpHChIpqmLtWAovYURNi3MWp29vLGgooO60
iHYEJilTWXHGAyJhda4d9UvdGU383J3T0O8eEmz7rD4ltSN7mb8+WxvRbKHguXg4
ChKYZ9vIGbwEa4uxHT6UzEHfVdatsMFzl3pcHIEI9wkLI85mN851DRWAx3uWprSE
GlgrUdxquIoheZWEw0dzqOP3Talq4ehL0h6+kC41U3VazPz2VYQ361rg8V2DDsPY
KiC8eXAXmB+3dMMZ5ANOtFk8intLogvqMn2f0zlhorrEogoXCFQJyBWElOcG8yaW
90y7kfGF4gGn7SwzwlW+jgsfBAhtHguVr0wzqtpRFCDPa/6ZY9X8UX8xZ8YYvb9J
nXFbBXt4tlibb5br3TpH/UIT2FDK3Xvakt6CWUOC7ptylLzfwkdSebDGuwvilhZt
TvL08Cmhl4f8LX+3vb9DXJy9rKulR/oMQsLMdhkBDAgRhYzdFPgYljQNP4IMyNtu
bxnQcB7wmDYhc83zYGdyyecf7C3pMRLm3BlkeDs0/NUtq/0GJp270F4rKzG+54vL
GL2904uxMlM/9pDF104JpSbs/jxYEqBx4aejECXkXeBPtZANlWqnztsuIIwpks+g
NHXGBnqzOOJn/39jgDw+QhNYSljUXMUFMcFd1XVQSrJZ8uVgMijVITYp624gcwrn
Ki49UA7jRCVt1N9F/8S5KztTUmUySYJ+6wppT1eYeu82TpQLudmV06LgjKLKLkdQ
+5RP4wL+wEHRCi7kzqsowVM5GHmoe5sH7/70S8XyGtkCTs2JwePZ2cxzV18Ho8bn
GNDyFOioJC0pkxvG1FrnV3vYVtBvTB2ANrMZJXG3q5K5ybQOfTzXjiNF7OwLFsbZ
oJX+oj//anZLCBkozRYvosoTSLzou9Gqaf5dN7Cs3YFaP7aJGOHmKXttoU6Akg48
Wb1Kuz7Q+lWsxcrgJkvd1LnjjMt4EmKgFSxQt55JsymT1Cri+WAYzRMvUx6s7JFr
0Hg4pxn4Q0OCJDIpaq42boFyMktivF/WjvfdcU5XEFUZ386Jnqw68bBbmr4VeBs1
LFuvKa7C7H34oKKR78dRq+YNawUnVwUu1nr3Sj2oKZXksQRWSEx3A/Wu+Pv22YHl
6arXwJxCpwBUEdnZHZoGMsHEmwMqsMM4uMBwF8+HJtR7eF4TJhE9YIa1FmXtXzxi
1/E0nwW3B5zmF0UkgAJ4oBpUZwiEIJgOnu0tFEaC/pydym3xNYIRSVpxDgc1t3Ri
EQvRbJhCzmCCH15WXN8jUicjdawVMmdBYywf02Hnplov+Qp7pXyoAZBu4ArJEzYr
ytAG1SN824ju7W+9JtRk7bm2iKsJ7RajIeCU4YPrGx0eGSYp8yDRkv38fmlb2Fa2
y3ZN4J8jKKCArasu2rYI5DCs6oYVFtRXnmEjPQlK7Xo81FQgNBDAP2zHnQOJ76EV
26vxD9xu5jdIXh0AWtGoGwJN5//sN6NomilmW0AQ3Z7DhpLQqUU5lVVuULK4K5BL
9Kn60rvSFc2UdbCqNhAcQxKtMndFaU7KdMlmv3TCWRULlm0z7x4xPA6vgewLnNPh
QG8jFKOgtCvUjx7qwujEYGxinxrdgxF5Z2/ysJbaB2R+xNJV9AGNHgGVJebVL9yR
TzfqDu3x14cVGIvYZdkT+7a6XK2mhcQ8h4+kGPYB97VDGho7tXvK7FOCtfw5AjjR
Lld2s73BqHwQt3ZPTA+UkRMARS5JL2NRoIzrj1MO2Ts84lWah8ih+e0JcqXgmB1f
xdkK8CWnjYb7ZxqxYY4WS/Ncmfyc3bdX2PBoQCuGNNRRHDlifQX71ei8LW3vPbQW
XQ+8SWFZzTdLOywyObZl8+/Q3SeuVD5jiC0YjEzMU7Q/ClYkaZhl4m2R8aMuRdZc
RAFBEw+TTJjIBGGaGwepiLUmaJ4ifWknneTyendr2KYjRvtBKZe4cfOVr5RvtKRS
T5XSBqbJl/5ZZ/aIiEdKMYBnVYjCjIISUQ+oUd2yxg/sy4Vowqws9EFHwkSQSwA/
vUQNqOvje2QSLdx+ju/zffwFYG/tyuDy/te3UcLM6fCKGbJ4pXgIRi36UdCBqW5g
b75aVahaJbtkiWWaCSXE6fNrcgEvdz1gypO0gTf4imG0P7og3VpCr+Z9S4Tzb6/c
YdCMRKeYtJ2MplgclDjcPoE6qe1OTqQSqsDXItf/J7j3b+ahPVLyGENPHK+c3xDV
O2d+wnDynflt/a7wRCu7qjgi3cMejnTcWjDUN0UuGSZUgDAouBGx3x2Po6T8uE3U
Cq0QDsjlu4yR7oakPjPT5ChDnmpxenoPpw2Vy8LqgbkQ3pusFndiUZ+JYx2FA9yr
4sCaETWVFnI7MXIWOJjUhNQiPRdgvmSC23zoUXGHPlcMydCJcnu0SlvJAFryxQ5r
Jku7LS9Z7vpAzR+z0N0MCH6MvZXMizuglKHU1ghVZIY9TXa2KJL+ysA7XHTZt9yg
JaluGs7IbozWKq19VbvBi1Qt7kAn4SBm+n2uymBQ81uX0y3F/C/ClceLVv9otvLr
FJCCsLu0rAsbpCgS6YWvMklJBjhubL5knrz7TQabd5U4wCKMiCwK/bUV+LnFVMnj
68mf0LNuX6ckRuNGheen5A3y6FJZo9f9iYdcn70+qAtwVttSG0HQLeffTQ2nPSJ2
IUkR5bS4KBWpf65QklwZgKqaPCDbaGcDANGV4y4SBDx1ugnDQYPw/FvS8fOvf7g5
rfZDAOQGMu4GtQ4lOyJO1se7IGarvjkP02L9grublHtUIj+wsDkey7cIyhlC98Kr
nwEMYQzvBjuZgjvMZyp24ZogWk9OjD21HNygyNiRz/mFEL3x1DYlhvnJCJS75xC/
AEnduxF+M3G1Doht8QNX6M1sFwX3Q84upO+j6uQ9nXOnkwXzwDAy8CSHG6j3n8M4
CFnndQF9Lh1kzgqpMC5QR9XxeKjzeGx5h/u9yDF4KmpisCACd85TmhjH4kFCsgVh
s+paewPye4A8cnyQQ5nKFzAZdFXAMNHRrS3U27NTmEOEMXscedc9GJt12Wt+Kwut
oIN0TGSBog948DCVmo0TOrtYZ+bBRMYXvk/J53kjJwk+pLrgDZ8OYH3iHHsdf4Ky
L+LLhBtXrcfdPkC1Iube5t/UUZIoN113esIT0Ryy5xWqUYC4O9vi0vouu7FbZxSH
aicf9JebnoZz8TB/8PDSy+kEPiwYq/+Lz3u+bDhATTyxauArZZY76uOw37a0ILRp
KUtg3rSps6JsIyzXWZVkXl49uWx0+kKx/qeSsJW+2IIOQYzun/chrSN5OZlUzo5i
R/gqnbyr0kAYEgFnWnbT07j98j9eSLBufG/PloH/JNIzKb2ArH3Gh7eOQyIHi9xM
RS8bxDRFArx6sT2LN/UWzKxDOV3hxUEPJgNNwV80wEyQuTPVR6GMzmeWXEXDDAIy
Ko59E91nHZV8aVefOTPBORBB7VTGqE+Yx3V+qqbkwtQI11euEp1OWo0RhbgsiVdY
eulPW+i4QyJc1PKmL1W+7IjNGzbMOW9xo+BTFYq/jybEg7t0Fy2VHMPgs92EZEQ7
u73leafpj/HE5S/oO6co/MvzZ+qaGCiwDTO5K5QQwPoarwGPm/1wBay7e6vKpOkF
z32Ndig4Ay8nqJjnAZLIv1TEDZxsSejG9pwWJhBW/CKyf7G+k3B6IEAtZoJRmd22
5tBgS7VEMAlVgvzJfRSPE35bSuJ9CXJKeBkbKc+x4QJLyI7CzRmFroHseondXVQm
CH20q7z7JeKKFOiqQ+L38cUk8KNCH61++GZFX6NKqN/FmQLSDdY+UjQWNefQ6z5O
s4cYwSZM1xaHrQmCZtj0tmgmdAyXj/IYr49+vkVeQOn8iNCx2IlXeohHHzYRpP9g
eiO6rDutwbKHhZmcAez/FAF78hA2qVjBvBmC3kNOb1jEfVrf4yMf4vOId2l7ULgm
a/5wH7RCTb9hq2+7oLPTSxjp8Vf/HLhJr/iW0xqhm0NCbWrJFRZio9W427k6fclP
PydAcnrs8tXVB4RjDFX7YRzjh5erwQHbBQLl/q132qBPzjxoyThQOahvlGwCTenG
IHhDhvQ84f7qsbpITiq7x7RyWuaE/xrUVtcVorLVPe5Sjt789/PxUMakNvtkY3V7
V6KJQaOl171m6myZjjkiicI8bPsGqmnGCVGvLroDOZbhgElfBhztoMPi6alzdrZu
qJqIRlRhnsfORm78X/Ygf8vNBg37ddCyDZEW1c5fv2P6q+8B2AfEWKe9/uAcafOh
1Ot4nP0AMyBTMXDBkY0ln5ouqGmf2zTCAUaxNdBlvOBTL1BT0pu1+8Gz8RavCPWg
RWq9Wrk1rv0WyShK+2oKUUY4AE9kArZ0DtdAqBo3eSJ8sFRRdaswGVkdtYkd2Zwy
JIUHc03YY5csRw9EqDOCkxJwmMV1XBvNd6OZ7tJJXCeAw5bjlSMYURgPHwRvNtvC
YcK+haJeyiuU8yWDTH1opt8KvybClK+p8mfNkh/qOS9uEqfoqw0TA3drgPLr5xFj
lxqyCOtD6Mn6kZ/vZuZLNg8faP5A5fxbnRGv+vekdEgvoUJGBgrTj86QQoZtUmgI
Vck6M4K4zpETXfsDj53cwBdSfd3KfHAaFb/04NDEj5ioDJ9MoPxy90dT+8VI1rMB
uFVx1N/6HUWUl1cmRiSAqkboTg+y1HCR7Ivz/ddXmBqXYqLL5LQyIAbYJqdXUdJA
WROKObsRVylIxEsnTJNXl0L8NYk/Fre3ytxokeS8+B0tK9uwKzXcROJxBFvkKdzb
DKygFBciZHDpnJEu5UMh0VejJj8dYUe9HtvNkLYiRLiswfLrgeGRHgN0fOqEaA4d
jMFBkPBoel+ehRtNmY+jf3XPWoI0PSKF7Hig3eU+LcsfSKjBMVvYlERlpop+zVHl
1VVD7s9rucBb4iEbpLdllbmxZTpJEs/APfICeMWhUXAgrnB9gWwKJKDeeZhmdxMC
gRYgw0MSkR01DxRCXsqdnkcYkHTK0C6O0AbxhYhjkJBfrjWPJ6iQ/QkhenbO0gx8
TJOJVHDXsmQp4Tc2nw6mj0J0gioMWLu7chGzb1yBgUMk59glzJix808EhM+Gp58X
YY0gQHiAF4ZEg/mNVwTpvPe5b5YZtgyCHAcg9auaBxi7mZbGJ8GVHGzQGW8nhdDq
eOIrEIYooIQBm5TamiR6vLmERvye1SmPvfzjbMExX9dk2i/p74B7T06MEKHKfneJ
3ruaQFI7rrrljSw4H8eRzLUhHsVT3+x+ZiohYdAroOex7Vb3JtmmHcw+vBxcfVHE
YgiFTEkjxY0Vf2ZSNG1vNGst2y03vAxgUUWijgdIrcAcU6HGMwwOSlJlRBeItbXW
8VeeU+AqGAjdYRxljD1L9Pv41o7N06jE2WWCEI3B/6/XSWKo+Vaub8miwWYb+iEc
Ne/igXQEJhKM1ofXM6Rc4Vh1d3HDK7MijEUSv8MsvgtGwfO+Frflfr2JyKPZ2T34
HVCFb0YIIfpKJZkRVxDbJ2HB2aHfTO2wtKys3rUfufmimcQucbklL+aIUX5u8njG
x0U8osAfAe71jO2uq+Q1s7qAI/G8PSdhJNu2g+Y4doINA3w2ivABHjJ4hz5aiUoE
VLcwcUly3g9Rv+3JOhVr35Ff1IotcQbBhYqRzsDq1BdBTv6aXU3ur+DrGvH6rgNj
9HncJDmLllBN5FO6RDZLtYXvJhYGQ5jm8j85STGw2b2NWrpODPbujt27Hx3g4IMd
CPJSL7skkCVsC3AqAAdGRdhnLc3IPg9hNX8YlW6o4wkBpbLnwnxQnsxkzwWljDoG
zLzLd4DkKvEAUCr/Hu4QzcbPNsDrKgk7HDoR+7HMR8d5CyBZFmFZvDFRAN9GOMn5
LJvOoP4leLyRrphkXhgMPihNEPr1DMkGw7v3TCikf8zlKT8ytJ1V2swFLZ5mw8+r
2V2E1HouuxnKjgH9vKFkzsyGQWGsA2KuPTrgjaB25DbnSE7ZHM0/U0Asgosw2T+1
5Odt0R1Yg2hYScKSZazTbv1nbydyFz0zSBz6cGqz1H6WLr3frYK9A4f4BJPvBwcx
3Cw1CYkrq2gEpWTiIqTg/K9q8iyS/lag575FzUfJizEfS/6VLb715DJIETU4YBpP
8RbB9YDgkc8NLb/7eEwm/fT3PUvpw8eGSwRnW1s8ANrRK83+9N1uJILeJupzWqXv
JTWyi3gJNlpr0cK5YSG2Ar3rVo+8preDzntAIk+pRrV64Qza6+5Vgx3gBcL1G4yw
F1Y14LRQuYi8XlM4LIb7lyD2qocIjUo5MH90aYvBTyuR1OuWkX0cdIJQQmm1X6fn
pd1sDkpEVP1tENvwxclFxNENytBv1h8jGYEMw4drpLn0Evhg5yhWEh7QzazHsTkQ
//tWFE/HTQDep6UEziJfBPVp4pLyXGbiLHH8oisiPjTK2+NzgJglcY2dgThojBIt
OQIZQ4GQTgxANlhyFaBAQtAH+9fFgGG4HST0a6jNwzUyZsH0tOCIxSkB3WCjtKkh
wurzObV36cPG8ac+DTsMAYBo7wOOYewVCL7NeI0RJARwN3TaYXzPmfEc7Dx+i/HY
POTpg72ZyZb6p+UNOKRx5KeVvyG6wv6z1k4afBezuRemxUDsQhpwP6iINl8xRI2d
65du2x+nr0z71WvAVDmyDw0STun0ucNNVR6oBB6jjgNhFkE8OncIzVQTSNP8BDLM
mCjIDMfZ5eLIcjZDVKp/X8Cwb8GIxdUdIMPSj+bKVz/d2PBt9JUo9+7oFGMw7ko5
qHJ1DId//qTOocwAVuQfjhLIocWesMB9jSH1p3TlBk5RHkNHwu0nu2eHs2lisiXh
o/xFzjByKXVan/f+oSERyJ+yF9wycGKhUiViDMXUC7Z2n2IS/oj1BriroXm3xBwU
NP6OFAycppARtWrhyac7D7COhd17jipU0CndBvjrZaWqrrBJ1MqbGGb+JsL7ABFZ
5p0oMyurm2J0i/4xcyeX7Jw6OoEZ8Jn5eTchIUCvmj3iWHyrV6otnQz7yttxE+eo
FtYamaYuPMPkTSkk9FPiw0LP4trp20VD53fmysuKg+zt9HZ8l9z7FSyauXP6ZnP4
dLPMkbw8jSo9ej4u2Ix9P/DiCOLVZHqeGY+R93mjTwqIfqf1aJf4OUMnxrP+jD2s
uhmZ4H6/GGcaiciug4cecyr6q/kaY9OKrk/5v+2VeyWpDc7N5bfSQpfp2iinBQaz
7hOqKHFRxDOaUW/i9kkwjO4F1s0N/xeUyNj3hw2iCPYfE2nWZFX7Dc96Mnd/quEA
jg7Aoy39OK6c2uku0TRLU16W1AJomhWX6P438iaotNqJ0Tzkd2RZzOjYI9Y70hgG
HpgEC+AX0rRGoun0eGeV+4AovIaNTPoYDfAQrdWpd9qJj5kcnpCMcOyaDo+x12M/
B5O2G/rZ4osA45w7FDjBieZRL1ZOxuFQvDJgu1mLzhVsgmt8C0BeTy3QZwWco5E3
TcoNqz9wTZmdp/ptios9/ZL+kpWAdsiXJFOHcGELxY0dim3URZ59c/eowkAf1Lcp
KhTvXtoI0Hsks3vBZpkxWBDLau2l+wTLMCByBhxnIKbkYI6vGPkv8rArgSguOp9s
kAZHtaNFreBu2640MVdOu/V69MykYs33+Lo7J8EtbywlJfouPKBuGlzjy2Pggmuo
TZWzzwR4xrwhBLF03hLBoJKAfDgVfIVvEbH8erI+Uk+PKaLSo93W3Py5rpijykOv
NtlXCefwgxEV4sJjoXKdDoBfJtR/2Uzag80ShPLEpZWVH8gwkll2gDrDdqOi7ChS
92gU10etdKx6Us400A3mUR1lQOz0+Fex1HvSOf5qHqDqzdzWmyk3jjVhRHgcxXTz
kLTGJE2TqFXU/GVaNfLGi6Z6FQpoUoSNYiWHCD5t68GSdXtAWkWQIzP44620hRxs
WVj9Jq2x94IkmH0ipb2uoC4+2U2KPJWOTY2+pc0nQZaZjQVflAKKJqAUqtZ2BCLT
gU6lf05jhJcnx8zPe+00DgEVAC/2/IU02buqu5UYPt7Bhd+zSyHBXfSEe0kgqDkn
greGA/ZU8ESJEbh+AqrEJlMglntSnATSDoDfzwCpMd971Lc12U/tMzYA80F4UnYc
Slc1Rlv3XHu3LbfEVHFh7ALfixMqUcoLgOPZ2mnXoN3eYRwT+zXARgmJQs3dqLX4
i9IGs6Du1qSMotQG1aN0Hpiyjozx3AZtqJl/g96/JX6ZCU4xVfXdCvyQpV/LkCnM
a1dYNUofAoB5VRMX3cHirgwtyVXX9571EsnuQNnnAeBMgSoekK7iFCqNpqHT9CeE
KOLkcvEcrXR/djH0zTsQxV+yTI5yU8rWiqCp06Xm2rfGGdNDZTPXUC4G+1lQpAks
W3rMN+dQCWxadtOSx1nOIYYc5jq/t066LMf5p/ieTVcphYMq5+JB5bmBoCa98ZvK
hJbBqAEPlhJ6MfHhD/Uoh10I4bt07k8BkakI6M2WDE9Jv3hCe7NWq2MDwfL7v1Im
Yugj9MU+lM3NFuOoESb0B0PeWmMBB2UjxRMxhctIjcp6AARNay0+KuT+qqZ1i6fl
Gka1GfQo6k5sXpbPtffZZPQEDz0pg17+K3lstreR/Q5kJPWADHXBfeRplXAxkjdx
baHrXboIltW9ONeqtj3m1bYH9JbRV0RwwueEZIEqMsta4K4KbSam1vVcWPbwK2kk
i8v+sJ9LtrzvqyYpapTaJekdFenuEelXEbJXIWkXVe+Z7ZdFUkF45n38useZWfqB
2P7djFJ+acvw4CUwvh50jn43VhcYZMJ0/VYuSnhNfcjDJ0ZbUTbX7JcP/Wn80wMg
PzYcd3OUqeSq7+FLRRjV0ycxPGmRvcRVbD7bIygP27CsxMQCCC/jszCihH4e1Dfi
mHgSRIjGbmScek42uOWYk4ZcQ83gdaSNdxC8xZZA7+MmlpQDj3yz0Vw8HjFT823B
tkX8ASluv5qq760KKRHLtBijSSMj2T8rqLKWM3uS9j/0FiNiIPXP4waKN8oUahvm
pTBEkOMFGlOCNBUQ7czfGZv++ryo8a8oElXLIU+79QtVqbY9tuWbm6xSusb8a6z6
6PoQJ+qh5Hcf7hSnthLwRgDvk5/1SpfOs3xz1BC2WYZX8wu/5iIHspUQJRnFTA2J
OtTVDgEAhrqHpxBppcugPT0qUs0o0FSWolY4Jozgehy1fY0zwbQQlD0vmmI8rnhG
RguQxN48sOBeDoZyQFrx4dc1JEesEPERiHkyKnzfdKug08RGWE2HPS4sF9/ZestW
fg569MkufGEErCzjk+cAfojvgQqb3iIgLBnHIfsjbYD1G88Yk7nTlncUxTPrOD0H
vaYjgTbEAhSFlidM2b9/e2aAvkWmA9PkV8s6q4+itqz1bI4YAnUh5uRjodz6SQHy
fjkvC5+iTaQOuGskChOP2k5f7VJgU8ju9pZ38kX/STIxfoDhzgV+88A86LiTsbe8
HlAe0Fm6j2BXLerfDAiblZCBVSsoOu5S8qc8ki1mw2sDw2sBumXLw1aCXL4f0M+c
LbarHgbWcva8BJZPf2OaLPu35hJZHbnyAlpBlTyDfPR5qMl67guMr3yp1y+ePh4u
8ZFpYx+8oj8inr8l9kKTaggOEm6VWp353arToQMSwR4/2iLsVHc9CgiKN52GVgee
dvVqc2dcbSBo508991ol9whPPfBWUNBcd7FxOGSD7t1S356DObiNv7gXMxOlmgv+
kvQvb3z529ho0THmQcLqEsPI1jFq3APbzZQHGSGGmEOqRKgOHL+AWUwTFI/rwolY
NRKn38QbtmZiuUGnczxzTL7/up22PxbciykQHHyVR0qNfaVkleKtpnp1iKnE8L63
SNb2uDdHGwLDvKZxLlHkSCFdxI38VeUpb+v8kuJ3Cda5KNWECTarTRJzH4WrTh/B
Fq3EjaaOjlMXMqEWXnsdmUXh5r0XQYehmzl8Wyp704YET7xyDN3SmZhOgLWMwTCn
jesOnJw7llVZmEOZVns/TdDfbAGV3JFU7xX3tn7FlqdWey+E3y/DNfOuKlw2LMVq
nhA6YCtCmxtf9iDIItZ+X4vaTcRA4FIjmF1LJ9/RwCEKB0UQcZB9soHLw/bYx0tz
+JAsI9hHaVVG63r/lHnSBM86YsuxYLBOSqXD9dXlM32q3OqbSvssN460C8TDuHrG
dNnRsXIxSBfyuCGBRaTDwm1MJ/oinpYc566R8TGSOd04I0/aQY5bmdrfRg8MursS
BbrhZncP7A/Eovh+eQ+q1l8kkcVKW6sStZe2nmoV5dWX8O3TOaxnsmfc1QAwbQPK
egPYsTzFqKvN0w56fCn2ectn4Lcfejp7APHaF6BClLnkd8rewq3t0HXyQDLVrAtS
ZSfi+W3+dgmvEHIZMQ+TXozDfXUslIBFMxHRaZy+yGXsD4c189Tv9k2NwXrvpoSJ
9c/TKfEtuF0BeRxweQEPn/NwwOlIWU0HV4R2jYZXQUnsUpGog7rryBTVeEA+m0PR
uiQQx7AySBB1wba1sh4TGcGSOjHRNvBqT3ZosG40EcO+LkiQsxZSpMwpykR5ORhW
Og7x9EdrHdyhiar/cneSLFo4pmId6BfV/RUj8D69jpHvwQihNNi8sQiNsDxPfZb0
NY+MQOrH/sqjaLksNzzdFxwr07FjoMyPCG6NXMHxTAiEzimgrnUydwHbrB/dOpqH
JIEh0gWS9FOnJudPEa/XP0yoTmpE/k0U4wmTEqFZQa9bEK22LCjh/kqL62TthJ8Q
69qXfDJQW+XtbST9oGnLyifFaIqv8a2SUzbf4FbOCFEawhk9XPZJFmj5cUYO4aww
8IQg1Q8E1/XpdAqm7qyk7idu9XUqnNTWThBq6LItuHReyplhrfKDctXMeVVMp7sQ
hpevM3EcYXy1Yutwn//MbLMjSVw/I5bQvxOqMqMN3yX0kO9BOSWRBu6gg2AAuhzB
J6VzsEsDO1PBP3+qvDmZDHv2OIiBosSOXxvaz8swz5ujqfcF/NMQI3tNQuSdvLUj
bK8h05agM24yii61920YSbjF1VJA7RpeJyX7f0crzw8mYSflZ6E/47AGgkCgLMrh
zqfq0JlBQ+ghaQcVo2ZUeC7idJ/jEkSPLOzx8bzx/b+cfi+yp17/CBSV4Vk4IdF+
m3DiKvH8yB+/pGiz8nBDioM3xe+GL8+n3qWxIBXkyEdxnnaZeqGSezTVvBFU1q1P
IbnIx+WPGHE4uRAR48RBa3kEUH5CvCRzpbbNCYZQFgRy8kN6GcKL3shwigrLjobW
ldPuPy1D3k7DGCd7amNecmMVydbmU5oK6x3JafcLBOHIZCS6q7e7RS3g86HKLABO
ccN1ugUALqwoJN+THgZuQAW0WAjPq8rAqRqGQhBHvmQfkOZVdF6VG4b1c48ndAl9
zt1pt8PruQNRwWEnBK72rxewopQBYbrJXXigaXIL+tLEisazOemawJl0lDuJXRUG
mUwadlfdWpkc4xmuxjnOoYWb1UzuoRDT8/5lrWaKvUTQGrMmvp6tvJ26MejNs6dB
8TzOFSjXFiMxrktmdqZnt0ND6QeEXNg6WV1IXrIyyOMCmUd5ZtJTL4oDqTDZ6q+t
rTI3b/5mCj2MwfL4SeD/X55p3Axe+KYTubszOExlNoNit/zocwb1oF39vrnPizlr
YtCKZYFQJPVwOQjl/j9pNHasRcMKn8sPl7iGI3OCoyIEI23YWCz1Row2lwH9k2LK
fK2IylZkEDyL7a33hVEfU4rhglo7vsLVmSTTe1t635ksLzL1nudPwsOG5nrlSqxF
xxo2k8UDvMiyWKODf0x0wQWTDQ9Y1ehe1KDFebtI+WlwK52wEH44WkV7y6CG7G41
30ryuk6SWZgXs69BD7R8Ouo409wqjLihWeEOLgy921Kd5ReH93tDLTmWpzjG8zLf
0fMEPUKrQVmKgdFwrY144i40QMqwJDvysM6QWL4Apc3HCbBewmv4FqvbeB+S0Cll
ZIynVKY8OeJh5waF1hnh6wOlbL3YO/7qerDleNkdKGXresarUct8q9OVrk9qfkTf
l9jZthggGT7zixzC5VTNCYAn6Vibf27x5dF/W59DFNYESgSlPgFjwnswTwiLf3Vh
XIDOAgpdbv1qvpnPW0WQ+E7YhhryDky1SUCrpk1iG164R1NgTe7OVsRNOkbeK0YW
AaLi4+KqJaHcx/UyM6/DB7RT7KkHGdOGdSkMSPkq/F5jYREs0kUlL2OEAKhzMWCs
CkioVhMy8V5xHSq8VFGEWirPu7ws3Bq1UZSaIvZVoUG0rpCVsOESOhXBbH9poT5L
Q3lOv+DydcFZxJUssVY/ZP3KylrpNagIN9inSpOtcZm2LB/b2VSFb8jpjakIpWWF
ExYQeM71WyPfKR1bngWhD4IvVBuG16ROKPtJW8qZlwk6njSONVMKp/tA83UT2ITG
uAFV1C1KNDCNxLJhzt1LSnAHUk7goxaP3hEkaf+jKYuwWeKjjCe0o6Tz50glcalx
aP80aoyAX0NtjB34e7vRwJDkT/kPl8D3mfK0TvqXM4wZN4tnbV/A5Kt9tGMIi4sc
mOzV9BrGv29RAKTOOAhiqB6qEPYDWP1txR1MiO9YrUZO4WJROIhyDhYEDTfhjzQe
PWVav8niuHxS7m6kvrWwAUJBMrQjvph5tWO5sufYvbeN2wE0eRBQlgEtEew/rXKS
JdNQQK8ye1Y89AxPlnyQyEKgVtwz7ky91cXg7EG3xMp7kHvE/UrjelBxAtal+QR0
JlJzUMgXbVm/gTWUrkcSjLa0WBvdJPtOKgBDRcJpCAi1pXWJfOOAE0X8jW8nYWzZ
Iz8S2dbB967uwKb1ffycOreDyr6B7GAvuuPPJ2pVyDIllrroHncvTkpp2oH8SvbU
8QAkH0KY/W/mWXvdZhz39PFWLLLdq2TPhbORtj7/9nNHMd/6oNGfHrug8Z70zYp1
RxKgIFmuCuiuImjqrerY4Qy7uMrPLXMe4ELpgl3tJ0YUhMk8ijhL9RSsTsBiR6FX
uen7W9tk4Qh4/t6G2pP1AkSp2ZUJmTVghYi7yd1MMIp/8B2QOmHtHIqtEJdKB7lX
oMgNtZDslwG2tXcxktDnCtDPhEGbHG1h/hr1LsQ5a3IC/xmsporgJ3sNmxX+X/zW
0h83/QCyOHQHOoap1r7etftGFJKSnF0SG/EVtUhVJulbduZ/KkJf2ayJzhdFAkSp
e4j+tNmCyV+OKuiFMm2uv9CBsGIzMhstv+9ml2lSEgJka7ZKwPMUNEDA7iSCg1uq
FnTX7tT44MdQUv7jxdoYEEHa5z7U+6dRUW7POc82Sl5LPurmwHIqE42CPkH5BOfk
AEJbgbWchG+RiXA2Xb5VULiGVLoMlMYHOy53o4jg04dm6+EIDPfzQkx6xmt21nyP
zcrvXSeUwA/2roUamweCb41CS0MSZAuGHQc4G4BaVPRN1eKWK2s3ZseB3iF2G9UV
RC1qjLOhlmKUGy1ZLXcV+Mja6LqG+yXUuV3SH5OnU2Y8I9+9BYAt7lM7579DBBhW
Jinf9TvGMEZtC1urA3uxkGK5wQIk0wcMV6q7Tj6iddEPwLeyUm+YE3N7zmoSF/8v
TDsQsVxQjo73TneSXsEgxKkuZ2+xYIIXKur73JCcw08qQ6VQqStjlZ4TVoCE4HWK
l0dAbe7IcLfZgTYw94Bq05FugzNWyQpTPlQicNoqN5k5zqn2juqmBfdcgpG/Jy8E
SgamZeTjyzhR+4rMJd5vkSS7i7cXbwsg2wmIqcWS6E08oSSZQ/AksljIRYqLLnyc
1qBYKiygkcvKO2Q9r+iTC6JqhV5aBfTgt9x+9RBRBergOgGe67Ot2NY9mjVPQRkq
Gagq3VhEntq1u4O4iMAehsDlgsXh+DvNyg9L6R4vkFqlv/geH0rX7AXGfdwb3ac3
uxiyNX43qc+6AxgvJtATgU7SMCfeCgvYw3sEmE707v0IFuUkYMvQ/kbR9GgZw3vJ
NAL+xP8l2RpmzKT4f+rDL2tAPNtKdSJQjc/g/tkXXB80IjYPI5s1SFdOHx2GNwLh
oGUxN6EdXrMR+au5SowP6jUZbAom2tw7nu2lBsxOhFISOK4owFy73XC/2LTrjLz/
UkEnxoCZmghyrJ7/0ZJzN0ghjSm6LgTp64sH5rz1oyqPOXq2NvfeUUavKdNGoZnn
bH+ibK0RgeCuo7sUV+fwlmEZQM9/08EBSGSBj1amxMx7KWKJgLASFwh9+isvO14d
NEDA6Qk/wEuN32dolFSLNa7lXqsKwWMeeNQjkvwxMYMTdoqRn9x6kO0AZ7hSx12c
r+2P6MIXhO9b2PnsslGD/tcNx3FecW/3D07OqfS1X+A+aVUEZ2rwBZoohHLe2eI4
/F0pKf71WWtmtcI8/8q8OlY+pSKeW1TeMKCWTDtpeKm3OJPO6K+QwvfxeRvSAaah
+LU0H6NR7XumZ3M9d8z/8e6SOz7ZXaMpKoFC66qQUhHyMZ91AMbZYN1ROJ/PAaUW
GtBCTOf7G3AetK0Uzue4H6Iyx+yf13kKQLchmZ5LIgEJ3mHhUay8U3T36fldPBCs
ZEe8BzA+RN1PhrvC8kFWv//al5qdH3+QxH2PFYeE8i4/ptmYgtNGtoGsyq5lITxk
qbmxmCrQdg8hoID4rk3omo77mZUf3Q4P1nJJtE11bybcjIw1Lhugt11d06PNIIMX
fbg2hwUwI5F0uZoZLzUtay/atWPZ+5i/mRrQrk6p8+GeocDtlMpjj0bBMrachoM6
+ktVB3cnRicBeubIT86FdXMfMfI8qZzMpCnqmnOVgCmXwStgk0z5EahyS51ywDXD
lwMJQlAkkUJIZRq8UaPM12BOo7h1o2f9yVfo61HpemcjYCfXjdBf8GnOlQZJ1par
cyEaFiQWOWqssCMDXOA0RM+Y+jamzNT1z6KwGUA3VpUx8wMJM9eEKU6ezvfE40mS
6FkS1617uO7NhnqEUmrLPhcM+Wg4ObKKMyhvRBLjAsEmcERtybH6O6LcHnH3krzn
tcdYFuOEGGL4mcecP8vCckWzT0PHD/975kQe4Hc4EigNnPRlHifGn9ke3cTE5vw2
t8dyITJzkvR26H6QE71pcHW7pmosn1EeUozU0GS4GVTcQHsHA82903V/ft7tjN32
klxcqw26I1LQcuTeV2YPb9NcfL90M3caO9lD1nHNlzNnfeBbvIZDyt/IRnzm6p+p
a3uOvvqwUGI5jm8P2NVhwFUetiCzCdeTsluYoeXXnElQ3h6x+5pbPEmlokOnlkNl
lQ/yr95elTEpAmWE0GsPTrbJ+3vbOdVkpyDUCG/+7Ftq1l/HzeQRSKsQMEXnCKdz
tu+k74adhMUZiObpavJ+ujV8r7A9USr3sxKO7jKk14zArsLeWNcEXAdAJ5k37t7I
vsXjxKWMOh2RcmHH3N3XUhYilmvKNwxB8+rj7eMX18GyBHrErioh54Fu9ADO00bY
Ljw8G9bry9k7vCcRnSEXGNp7VmbkVaaW6rVRxUS8WWSTkwNLFsHRj2QlkyOakWDY
Lu/t3IFKQcxNjMWUAx/C7i7IGatASDbCYIueqFPrL9rDKxSWmRX9GiKkag2DtFe0
yh9oBVf+DqKE+UlcpG/TyTxl/DYWsL4Sc6NqisZ4qF4dQ911WZePDWRsCdsW7NZ4
uuP6pdyORk14FnqSiJ5kXUlVfjNR17WZRl4BMaTnvryficHw5YIQ9xypKM4d51ir
eaJbcFafqAow1etKeFn0SUk5sazBLMOTwBzOHxoIhPBHwB1OHvBHHgENmz6B2HPr
e/gVnVXPG1nMBxH4X2AclekUJ7m6ohaCPQzMiCROchJOUf1XHv+1ity/F8wg4Vr3
ylC+1bUyVBZma2m2ofAQhQnihV5Aonqyi4uL5ki08uMOQKMs+s/E05EIOw8aLfGJ
iGYSa+UTgL39v6yStEfYZrnu+n02YXDODzWvHaZ0nrdlNynj7yRV0EmKdVxyHTry
5yeLFLVYHqe/CVBIVVZKPei3tyfTD3ycjuc8qCPceZTwZ+iQTi+cdPyQW31h2r3Y
Fi4fRW8RPHa8JUP+EvzZS4De4g+D268B+nIKqAPT5E3wq3BHrgBnVyIS533Id6dw
dmNQk7JjvTgs15wp2GSicS1Mlqsmyqif7m/sSf+scLpeYgN6WdS8ZnPcl+M9n2sh
1neEitclvcmkDHbNpC/Ga//jV5yTtjx6sGXjxLrmaKPrVpEi0miikT6ESl97xTFu
aWVVstUUFbdxbMZQdwSks0guFV2K9s6fq4aKJ6eiY1e7iJfTKeAwcchSoWjv3RzU
OMo2oDB6EZjdgLpr/wHUEfVeP/FR0odyig//LGXYRnl6XgYokt8I1MFf3GNC2ouv
EjWxqOuMFz/jqFnWkAYzcKyQofoEajuMBk/QDXBL9Qo5yw+d8wiaENtSXwNodySk
dVL4ejMfXhl6ntm6XEPah62SJ7/ngmYvVKGjbTKYJBaS2JZubAkKPt9EhxPRfx3q
PiJlA6niXc5EGL7+F4Z1lGTJAa2PZIbP5PHyyS4wbrPH0ZlbY8QiGxLe7Z4JX3Zr
7fApAVUt0RKEl2P27LFPeuO28ST349hNM0yfqTV7cqSkN+OSIP0ZHyUYnxIgrBBo
0hOEUd/TwU86p75jo085t9TQcigCLsT5T+8EYt8pxA/EBb7l+ixVBgUVosZbOPh2
BXMyvh5oyNFsVVmdQ+rl8nn3ot8awVkAuZ46wNm//MFrEtIBd/oJ685dvWdfnPS5
3ebLrWF8eyqhiluf+833T/isgJa6BAFZcjGeAvGbZLdA5b286w3nWaQnFMBCuto4
ZYEEyH6mTmEZJLjKZpMPe+HfeNbeepryXOACUbDKhLEufZ3A0D9UjFNBHMpISXja
+nPtxfpsiPvGJM+5rcAGVScz+YLKlf5hwct7ZTU0xQbBYOssjm3Ha1MOJUhbWqp+
VtZWBDXrBUDY8DM8z4ieIqvRsmb/sMX+nSNjEFO/alpzkT7CKQLv8HiwGH7uOLh2
0mHrjTb0GFrxB1yKnlC+tLK3aNWsmJ5KgDcqiAVOLLuevMe2Cbm7c/1L3mXHuZuG
kHyiu7m1Xj0dI/HmIWNTWBF2VSe/MBNXR5frvLWo9etC5SEllW72Ew8O4/dQRrmW
jwClmgX+pkEkMwQxPE062fcR3jjH1Cd21kEL8q+fjElsx8AClDFDYUdTvfi17kYl
gtVMnGSvZT1YcBc1i28Lp7P/J3OJLUd5kBKqvuJT6pl7TS2EzoRI4C7ebbktyUfh
InbMNMfU9UBMG0tmooO1TEQVEkoQKiZvNn1qiT6XbfdgNoRbH1h3+OelenK8yeUv
67jgPjNoDqyzKDo0fuZzBsH3rACEa77syDcfa5vctZUSvbpy5Zv1WEyNjW7yGsCh
RI9fJAjBj0LNDo4oISze0QD9m+WlPoeWf/Cxs/oZFGWgYSVJ3HRg4auF0nTMo7W1
MziFLlDr7omvGuwNmnyRLwbj36BTul5Yc6cjqyL+6JTuJQ5ZtMpT1Ys9H0yLEMij
v39+GdyKDdRMYRSAl8FO5kBEgTGf+CSJunn0u2pHWklCSbSiqUQHRzxfPsGPx2wC
yrKKsifXZpT8tl6mhwK84/gHruv5AKsOKn2Mw4wRYZ5XS80+BFEQOznop1+BURUd
E5CcTSA/xvEFNNPNdGKFSDJniNDYP3djl8iRy1eebHzCdrwJ2KJbCV9Bamv/3eP8
MwZDUxwtg1sjU1JujMwVQ3/jRhAOGtGt90gblsapbQ/8QYzjtGURcqFydhJombs8
0nxCErxs8z2+aAEDBHz18ZAu5lCQ9+OQ1uu5SgXD1G2Tes52Zg15oMJfsQ5q+CDt
CsnCgR71AUlV3pKkUg3++rlnClktEE7RHyUWuNYsIYOuQoeO5FLoDU2Vdomolcg7
62s6t05v9BUK9Mwg7l+WOLGz7efGGw1QjiiDUWcxR9giVhQJwsDggVcB8Jz7O1hl
3rf8wi4RsIqugJvwugfqAkiPmnYQcjCs7mNykpRKRlsCpPBJofwU1Covqc6iVcOD
OQP/5Jfmm2V650uwe79w8vvZbOkY3ieO5fkBtOCiJbQ5yixC923qbpx8FwWrzI/S
6rt824W5eLLT8MaNR8cxvy+apcHf+lsNqY3m8x2b+OpMXQnM016f3yZPbqIwszbD
6sPkSgOYRvNu4Km+b1E9UC/d/v4Be5mYeDTOk2fBUKGl7Wl42J8Ke4qvLfZYxjWP
EoDiVCiR96ypkLYw7WVI+J9zc0Xfi6Se1sl4jRL1GGCGhHoXu6MNh7lB3j53KGKU
K84kkkkqHYqHO9yfUADee3/u0kkWDs86Wa5gZth4oGOl4E5s/TjJ5TVHpk68+888
8w3XLK7u5sgvW9P+U+TuXtcX2L5ZHqt6raSaFGvdNwVt12ElAnNEfLMsZUoO+lv5
NCLzgSPlIUAE8ajnTrUmHZwGe5G5Yh6I5k4yf27PfpBdHrDttCEhmesqwzf1wsCa
ZBlDsVZwLLhG2xXaw0qYfk24k8Gpo01QxrMwdADkmOSGNDX9VrVdZ3QhhP77xyTJ
k3jTS2eTDtOhZfIQUJD3w8JhSstWt5e+D8eNrn5L+1h1RPTZL9lhtLuCQUsJKwbT
ZqgSRdJSuKv5BdzmtUADo84ZIAciIdgMOuoUV3lqI7kOSP2GwVxbJ3TQdWtU9/Ig
yV8b3mKkhjXRnxRX0g0F7SjOIKiQsT4i8bsgdgWBgjmYD8WFG9iV9t7OzmoqRGE6
8w/JXcRMIX+h/4Ru8csIKxobuYxOZl5cVMDClRxRmCUP7w+3XnJIyd8w7LMhuzWa
IyvCIdsN80aA/3cx92a0c4RQ8E9fwhkyEafu0sm51GDk+z9Qy7rBMBNK5TiBUsdX
7BTJpgfF92rPnDZYppJ4RjfTWLF573D/iXPUUcxWFVeFmuTPnS5Fp1BPW4nGIhWG
bJBexfS4NE89k+JcAJI8f8exnITkPD57AaltehmtbmR3HPW88/PbFE9ajJCFHRnD
kbeeflFnHIyGVPvpSm/uigzIAOoys9dOaRIRnsR/9/GOeiiFVlZdNNIwHPwjzj6u
z70ONDSdzDXuL8hcigtQPCzcjOxBh8dXEPz2swEvVR80bbf7XP0o4oSBHAgswn2b
t0vKxAsDWRDHV14b6eg4NpHzZ4pYt/gV8ymE9h6thvAq2ZoW/TNJMswZn5BV26R5
H0lpJedFT1DX583CCL1h4/iw6Ric+ZOr+BBOcoMOViI8sJXW0I2itdYvHQszKk0B
HFlTTkmXyabLDF7ZyNd7Vy/iuoTPLuvrjoJyO47hA/dAnuqCeao0QMJEedo50dGp
K2f5Lu+OjbB+DRsG+feJ+2IRncVWLuULwuaa/IldVrIYQGkDbU6c7247oUA1uUaw
XuUq5KT9QoMQA2rAqBH0q/iJLYi+0F/yJh3AUeMsuj2hUub04TuHq0qkG5Jwp1B2
7SVlXd+nszLCmZl6wOxpXtmfVNimuo3NLxPA8AMcl64eAFapz19/drlVjGJ4Gsnt
qD31O4H49I8C+0M3+N81zbvCKBOIh3TmekEaWiNTf9pougSSpgpimF6ry7e8C5kR
EdDB5KSshfCdWFwtcIdbV4Z/NdoLOcCskmkXyZnGO5RR7wDyqtcCtDuqwhbgXsk9
suK4jr8+RgckFcrml87yOX8v9ALiXzuwFsY4dMvlbmbZP5Hd1sAD8NNmEtwtKeEL
XCf1pm3CzuI9VqeOK/M9hQPiIKpYsZi8tEaAWsCBFCpCYsCzeFlVcMoNmVF5Raz0
JJ8f4JMGQMROYQyaIv52W3u5p+FcTVhypcWDuVM0gRQaeBAx0GCbqeHzLyIW9CCk
tGp74Kvk2fAZUkOw16t9Ncx0Vz3UayPZGqLD43Z8vIhPJ3VJq25TaXwXWMhiqET7
/ha+/DmcPW8TYBxN5tvMX6T0cOB5/htsGP4WhPG/WglrvnClmvUyyz0KVaFl2PaA
4i/+spmLKbSs4XQllV5Dfg7mmk+Rf+V7u3UYAS1WDTMmw/tloHvSBvQJl9KRK1KK
7DdPlDoCzYloI/bAXhoFhSPCoxSFWsovIfRxMGZ1PmKB7TZnYGVbaOLqg+/4mssI
hVrtHZm66c1D3r+nCbILqlJ1HMhLzGH5dbWJjftmvF3+MjsU871E/kMtsbFaTDOY
1ct7LeBhadiIv8fSSSCjQDgpPzpACZhVGoM8gROvu+qwS7+RJWWRZ4lDkOwS7573
vDXLRZOGIpFld/JM6FzwoPbsl7yHhMLc/SSsLm5VU/wUmK8FiYVEmfbpsWygJQYL
sD7hdcfMQE3WpadeB9Ulojwr8PTbYGtEUo3X272bcaBP3oEx5xRiHmCyDjKqBmlL
C47vqL2q02FJTLcG0gDaODWnFX5fFjMRCTotTjMH3zuf8aBRX+Y9yK3XdsXscoiU
n8BtW4ESkCZ6rFpR6OtsrKI6zYDiaIxTySLZSq8qvzLIyLF1+keSartNxvh0gjaR
wJENVnYMaX/99BKjtyMsf3BAE+ZXfYPE2ISEHQoW1GuookhBbfb0nV9FSjhRv4W+
O/PDHy2lzSLKYUTepPBf/tZ/gFkkdyFaUu2Q20NpD2IRarC6NdKSwWpMJu6pqwzb
S39bPNfUV3Sf4CdNS0TEQDPtJ6bqcOVXUtWGny7OF2JcUfYTBjcljvlWDnEHRicf
Ckb+2tKrwkHEy/LayTwZG2NCvhQUOyDFqmb5638jHTwaPAMcIbcuNw3mwPwKh/Qs
LSCdkUtZNaN4p/mNiTMohN2JL9bovQrKuEiMcE4HYkcmDOpxjgwXVRuE7DagKtYt
5tXvpH+dc5sEgIEOh4Ba+XYs9X+MMahmMuwzfLieCwDb0AWfxF/1jVaIYnh1u4mz
mTHfQKMkoY6GpV5hIdhgOi8HueqeszgB1gEOXABr9bnD88Rh0q/sL/LaKaipPhji
1QaAc06nHcAz0pcd9YTfw5Ec2IWVqIWJq8V6iQIkRjoy9tC/9OcpEs8jRdpjL/ou
acrk09tVckebwXr3vNvlg0E7B2+WwHPdSu1FBGx0k2rN8WsVvjPBy6C17v7xx4Al
Ch7Ah54SHbnSTkXXxcrvfXy6VziOdMz59h01AN97jxtZRsZvoFLVjo/YrtZzW+BL
BTZ/PMWsgx3kJ2/GfxF3ZjsP88/wPwUdQ9nFwTUj/d7S4wHV83lvlsNiXOTq+wrs
8amzQ5w8hdEvgGTZYkZO7O2561/fYpjxH+HIGUikYnsdlBZ/2og2XHfV2/pefo/z
odOMzJlNxhc/CJf3Ac+0ubWn4ePPNmYwudb/F0Ia05v1JSORydVLrk5S22D+Wzg5
YBlRGzZIriuj0S44P1sZ/isv3Y2Tvi4xnr/9919axXFJOIpctDEqsh99MhGNPu/P
2kv5XECfRT8Q36+KQCeAQqZEm85aEOOdJH3Eu/kKB/3UmykJxS2mO14olk8AVj8Q
hdZHXSeytZYRCvBA++Ay1so+mgCTOnmQsY4KaFTXEsq/25XVHO8ztVLEEKKOOPCo
TaRTPDlI9XLXnWeS1EZpsitwn1GQguC+TXDU8RXBW8y5xpcdKex/7fbk7dQpwblL
epQFVWcPE5RwNFCeqfM9iMfXUU1FkcP1YTizmpvhvQGXQ9LBqnu2XmojYbjJh4eA
OTDj7JDeepqkyZDJgUC3cL3Xt7WRX0KQ1D6uLwDDxLUS4evlPoxL35TcNQ2cYk53
Sr9v/5L186xib7E4xszrBL4JIlSUyTXrU8t6FElfgZyY4+1Y7/tvARoyWB9MqxLw
y5+Ox5sBijhEuRGfYTvhQiWkUsrqWT0NQs+InvvSHh901TKHoEB7NuflRhARMv5e
8gFEj+wqMOmhX5pf7zTFCNphPoU8DT3SvWklHn3TVucPL41nK8j9ryaL5AelqQNw
cOR9UFU+V4T0dhJu99hGmh1grUep+h93xQH90NSAlQ8D2pRmrcFbxebhvhn6Ynnk
WavAE1y9ny461NXOHsOWcAuvALj+pduiMegAifU3loILBZVGSyG8KhYveJYK4GXQ
mpKabBZeHjsio4rr+i21CPhiM0fHCv4dmBUAyyCKOdK2yd65y0aqgFunqKUCHYlt
x3osU5/q0wut1WTExVOqOPPnQRNkaNYHt10tEWVbSTSugm8pz5TNscU473qu/lCt
+Ca5rjNgYZjciVF9nsrhMPGLI1bDSzYLo6+SNaTwgYG8/IQF7aZ7GV4MxwQaV8M5
uKJeQ0CK55w4y8JYoNYTsAtl7zYBUyIf4yOedQBRzBCVh50UGLT5Z+7MUIQtwuR6
HUVKc68p7WPtKohvnGj16u40MbD4ALSuA3HdCv7CM5YmYvyeP2sJlsHKB3cy/HKB
Y52NyvWpuGS1xPZnF1+mhIOBDHqTxwekoGjYRcjbzFedznh1mta8equFiG2SqiDA
oEJt6f28pBS7SlG26UBUwfXXOcpyg851UqMp47rrxYbnjQNf3zr7ZfScBp0lHwae
nFWzrOGSov4lgxXGcn4u4cz1eGs29HrBC6EMod4kE03HfW5RaMgP+ykusDHm22Vf
egX0/BeCKoSV3/MbYfS/EIHZZm0S8MEtOpu9f8HS3s4Y+T64xUaKh4GQA8q5RbDf
BU+T9cnLoo9FMhVkti/2xV8QF5+NMgUOZmJfyX7QxDy4SgiHvcwPYm7ndkBBe6Mt
Ut2B09rFoTflYpjqWyykshFDa3pA6mFHxETR8eG5XH8jZ6mBOGUd0GwVObOa1Snf
SehXOPU2spisV+4vKFZzrB9c4juzBhIRfkp0U7GznyL9XNcmctQEE4WKL3DC+aW8
H2ZLalYvTb2BhqK8hQd2B8ErfakB+HJCzXu5SB6/zguAKQDKRwuejjZYP0xl4dJb
aG0zeJ4ftOAqBOqP2TS0X7Nuk1uuRFhkL5toDwOm//h1b8VnanFxgIsRVthY7ZPg
v9nybCIfxFTIVonyoxSxsYRly8Ct5f8hAhxdiP+pMCKnTSGe2QIlmwQIFmHRc/Rw
HxMExRfmWWboxcTPrCHBqbfyDYSwiqRBqxxyOlo1+MdJr9ElUgIxzy11mbJTOu6M
31VbkP+Z6Y9xmZyrrZX4CrWHBzPGULjGroYk2ZVQsJFx5asU/ISdzuJ16HdOtgI7
+4fejqHewIiVr/F9LXMP/AArJhd1x0tnR+a13Vjf6YYcWLSxsd94/kKhXTZFV9g/
VWLzDIOtZLSRrYLoEdrcydiqbwi8xyvrNvzGs05aGpcqcl/6FEyQJo4TEM+Zcl0i
83Y/5zzJf9aEN/oNmTJleud172w+zeX6xe+UwC2iSx93WPpA9GnpaBYP0RbCI1pQ
XvUpgObjuNew/cbx1EHs2NcyJTiaJQ3Gw+WM/cbdetG9niwRsqq1aJ7wL8E0POlX
4EkU36BIN+4BEYPPueVmqM4X6uZl9W6/nUAKrnnKdN1mUSRRI8dgFbLucaj6LC4j
QYz33Po6yltEp8wRE8gqxHOabwCBj2lDJqvZMJrA3dI5jWIvNN4SMrCfNowK/mOY
952fsYKQmaleNMUeejJfgy2g5HJqRUufQb6de0lkvEIyuI5zeVU3HGKxunxvLSpV
HY3/UU3a+89KcyN22+UegTFoK2Il6m7q+YmsC3jL59A3jSH1JCW3GZkQAyGKZSA1
UxDTYfPkUb56lLZ0k01aCyUDSWASQrf0Ji8lN33irlhPjf5e6+JZoKoSKQycqAhw
fChWsqH/jArU9DRfROoWsjXqj9uwTJgQlRFlTZe1zc/MT5VkrnITjmnAxHME4y7p
NmNVGpXJr+NDbiy9xlHdgaMHZUuy4KKFM5g7p3t85LPO0AUHnPb/3fLQHnBskpH7
9aaSOqwxdiZ9eqQzFWz4u2UVBWngqSPDRJ3TSSKvKvGVPvzH3yCVYvWW8j8SDkPQ
BFMFISe2Rezg2t/IoYk7z9W1Juzbybr9pt/Au4fwIaBlnmSyxD9lCS3WjEJDSG2m
gCQnDrI5oqH0gY0GUAT0dxO+rfKg9HHR3qCsAUTAlFM+bYSnflSb7DxB2aU4nzOz
SyIag1q9+sBn3/V+3bIPwZ0XdeTZMjYQ1w4pZ+q+Zmus6rw221nz1TGdN3CQ1WkR
SiDGZM8MU0/SEs4tLqPQNutFrxC7GAeHBiNmZU0i/dXURc9MbQxiFPOfndCN9Al6
HRw+/qiVDt269VRl+fbNo0U9fPyB4rJudAjvidSfQaDJKDHY9DO8dAjh/uqu67Xi
/NrIggd/Hmqumn8WLNnuEjkTFOHVeCENGYNrL7K1vOSGZ582Om1Zrrza3cppeV6w
VWZOwVwXOWBv4IpOa2SpbWHuq+kvCKII3A0d99pKqWZUGPPJmTngK6c0YgDIHjGp
oUJTVJqRQZM6HUsubn3UmnwVsSSSEsTqP1y6mPehvUpXJZd18pmGIWtXbiwcXNhK
5TvTrrgs1qVDdcfpAVIYXkcPyxeUJbpu7ikSDsn+0CYcb+qijIKE6BA0WrATHz1D
6Js2IE28PrOzcocwlvT8XTPjBWreycYToPac8OX8SSTSaw55qP50koYzYdEgT8Ml
z6lPR3C9Wtv9Us1ptvgXKt47J7O9hPBHzj7Uo8e4ZRPkdfLg0mva26MFjuLI2pCZ
y+I8I227l4n5LOB6atSbl0z2yuK+HpjEVRCZuMfKHywGbrRmI2+UTF3wbSfzEYGc
+9wU7v3Z9u1nZbNxL9ciwXenKoLU04FCKt6c1SFTV2hb93t9aHOlLf39RWAOprFx
q+HYQIR9flyx6bEEu0ZpYYft1Uzwmj0aZjMGCHqP5ehZrbirfLuPkGRAuZc7DuNI
qh4+AQEcRuFz5IOh7WyFm4dAj8A4Xx5nm+Yz9x68H9hi/nfln3xl3YPqwYP9/6SH
klkheCTUpzRoVopvdH7bEBhWOuyGAoEX/krM7uPp2tPEILSrzxDEtap6MO9sSb5a
qoOfE0A3LJm9G3ENUqehLLeHIgGoqjhXeFGxSIu/8Bo5lyJR6z1VHSY99xF59e5r
Xzd2JTUeOg/gSIfjr3e3FnR1q8mOe/4Wjsorta/2Z5g/WKjYWu5SNrrIGips6aGf
NMcQ4Gv13LJCeL/+E003QqaiLIL74ReTf7WYWTq55fgE1a/iZsCOzIilKrCSGlsi
SLZBcKdzIeDbGOzK7Uvnx8AWfangGhtozjWfcnm2GwBSYlI/bK2JvSNEfVoimp5R
kClk+IIqt73Xu4G/ni2GFCgrUt2yYWcCslRu2VaZB3U4AmaXJ6eX43Yl1AlRIv6S
Q/JXOXt2dHSR6PXevJ2K8chASKyZWOKonvzNW/z1O12TyC3BwW84bB3KBAmoKX50
XqRk56E8pKgq7LTpsCKVRgxa6pUgfiIwUfGfQbhCUajwp8a/L7YUMNeKEpZpuP9w
/3bw6KYSQkXbBwMk5u2rfGGP0u67SyZI7B2i2M3MLQHZyow+Q4907MXTfkuwvyZT
I3YKhMCD4Asjk0fnDBDNTR6Aj9MGOVKuC7woyvP+MBHneKeRZjqwgBzI8aXej4WN
uOYFimunuITK/2BvkO0OHtSSKG1LGpY4aKobaSQC5fs2jQ0Va9A/KN2po4GV0tL9
56TwwRrgTkBjQtoLpLguMguxOLlvAYg4rripPwxqpOWnV7N90fh70E+SrC0BQPfb
/l2CofKT/6/J/Kie+0UPlZA129s9+x/wvEg9AfbZ8YQ+2m6+gY+sphV1ibK38QYy
5NJjmb3FbTubo1HC7u30UUIo7RNhJSrrHdYdrbQ61sHAW5DtodXiZF9MBT4ATfVb
ugzz+hXbxxfguPF0ggEsRDkqYKvPIzZ1CpirJLtntxWiqTXH9BAfgByHoUGLzFbW
sveGA4H15AMgatSdoUFlK9w5UumLUaB/UHVbcYYt/XLLFUV2t8OwA01X1QIWgo9H
TVX62m+B9n5wTJX3AFhwuLwOGmd4C5J5cYnMV4dQA5jieMcA1A3bAlqi5v2nj/DI
i+fnYJQNMDUVGBYPAEGx2HiWO3BkT7HBrb5TM+9Ju45/KGuYY+9o+6LT4slyuMYo
FYRsl1Sx3XQ3p8mT59xLFsrlqSwUhxT5jXa0TwL0OE/BvXHomB57GVbVTXUzwtm9
nR+80bljEOd1l6C1xm9Pwo5OmmZB+QUwf4lx2VSF1M70KlEWXqWjZHdkHGRQR9nr
D4eAyRvR3ONkVvNSCrohG3G33VfoI5HAJhZjQzeErN33biti4jA8dlH7JESRXwKg
qfLfQt97qhQqC0AHN6eMlK76a+LN9DXmVGLoiG6pwKggP3sqbj4AaEfDIJgi89L3
JD5LTdXij2/ThdsaRE3wbX1RCWLPLsDpd+wyyFmKXkp+tsVqldwJu/9vjdejt5tn
EStv9epPLOVnPHy6uOZBrpzxdTuaRC7swOhCqv3W9TOiVl2ArLTPtcV8W75tlJgD
fZZ7VQgJ8+GiW6tXGE+mBkqh0JeZY6CEh0ZDg6cdqjkFvTGTjVBYTxgNsNRHBoEt
KdCPwTeqLu8asLF7MG7v0HZFpQgEIL6KfB06epKFNZpTfHPtn9GkiQ2C450MEn2A
Nziix9mQmW/WDrSQc/xRNyt+rz1N2iJT7eWLfaJRuVDzrDkzQTcEjM43fT9DO19E
RbAZ7u7PeUIBKbUUG+vAUCR16p6Av5QXR+vjZrKiP4aUbezPPc7SJxT8apxVc6fW
KDo5Oqg3jMKlHrJj1H0sAWTfewvUvzuR+RaqfzGcUMrK48Hcy9Jcnl5kbRliXE55
wRzcdgCfNa5fTx235oYUxff7D3hqtOS3yTqMbYP9ZNBb8SZQtX53HNzsDxxCDXTa
pc5RINoL/HUhnk9mCPXlmWFhrYnQET/IjhS1DM8VsJGrz3ksuW0kMSdEAr9DPKCZ
F30M/1qU11uHj+OP56BYWxoEg8sWwfsNzQxCPz0YAkSa1XOYiqy1bzX/kgwIyB6N
l1DeddXTJxXGWmkdmGSIkrvwSyGf+iOk473wBbF+8QY497lkaiFkxv3agw1mmQ2v
Kn6S8heUoFO0vtvsj/RpMfMqiWgO21ZPPELr2BInYqYPiXAQSS9yFgMgE/VGmFXY
Zhu/vy50FoMjR0x0e7o5xQULdSAczATIuhYeJFMYZeGBoDsvf+YNyvw57cGcTXS1
UB4qaj5dUmVUhc1IaAD38yy75MpewtdSZNQBkP+wgLqhIcOaylfI9QAXf6VqrVY1
C/Y4ycg0y30a8ttUCQOkjq/0GHvyjMWVcW8CbvhVAz3/EletOxRS70SmRRJZ1k6V
AHvJUYbsVCYktYnniLoDUK8lqbwbZHv0NnrceJoJGb8ikuyJhPa6f3mko+E7PIIp
8k7TwCoeOjnpMR70282O2/H2p3hUJJp5+wFs4ajIFrQkggEibeGH3SABFWfq6KTx
Yn6l8OyVJgGUsVgmsuO2hLWHA99DDALH7k9BqdMklM+1905liO9ThFjZdJBKtGht
HyacGR1Eedph/hfZ4Jt9j8RWs6O1ZuXehtwlKtt2Fqw8o9aJ0D2pHMDE4/0R2qkn
HyHOzTjRJXva+xl1BbKfo6ZleQYy73c4XPayHIfQlNcVSsZF6yalygatvXtxKqna
8whNpU2TYMl/xVp4tZBboAy0+PM9kgUI7FEdtytNVi6YvZwBF1CMstdvmTL2SWQv
Woa6oA+e54qg7DpRnYYYVSdntIfuHcRTsTgEuXAG7bNeRK1Qgic/pqMkouaUmdmc
MV7s2Rpg3NnOP8bO3v9QZj6h7dVF31W3opl5pyWB52K+ci6vsQW+lrWw2e3vDHK/
SoWCBn212u9KEH4/8cBnK91ehSLd/UlWKP9Kh6B6frEns5s6W+7+VXd9QFWIPs3T
P1PBuOzkKoQ+ji5NBh4+2SNop/+Wo2gXszdiIjq75tPGkkSByYiNwgoP8NNQvN77
1Ou8Olcq5yyO/5aHsaszuYO+rr0LchbzA/n0oYRM+5Cvc7GLnlKAIM/SuK0xC5XE
uJzW5ppUiWVFDkJ2OW7zcf59N+HYzUNeEEsfig/2jKW83KSCGntzo0NRlhxhEeXq
gPhQBGp5mMgSammsEmsk+otIely0M1d6ThUqZgtowSbE2j1slDmgFhAqzwl8cWmL
emJFpkGqJ0kDHVhCl6uVLcls9WgGJS81aCsckIDjynsdATrYzkx+3it1A7Yt4Mh8
j21jb9xxZaE6s6DZwyRMOPiVv/DT4GBK4jkWNC39ZrcrCCboAxsmhmE/LilTYN8p
SFUgvSyQfyZm94aJ+bFN8GiRBVksq+keImlGA84gXhxHvMXy7YJIj9J4FNudGq+d
DciIqp+bsb9Y/sES1jyEulNDOoPUsMQ1SYYrJbmWTwCBvUShdMlLxZZFVgNEBf41
k5NnvydQqboaH7AiW9tm6UySlF+eB57txAFb/Ey6Z+ew0MHustlJsUO/wIbtWGV2
pivj+tBc27nK8h42bmHup7pJkBDd8dxi/Pg8TVcxFNwTD9oKcSfU0kWKUvY4SDzM
QmMsZtVglsE1p7ubZM0N1tZAYNvqCfVKRgKRGlZA3bRvNCu8q+UdVdIrbVurdg2W
OZ2X1XRIJ8VEqCGWwNoJeaoL++Uw0j21PN4EkvP25kjds6vZiGAHxrEYYRQ+ODk6
6wz3wWcP/2pmtqTUaxnOy12uY7roT3O6l1d3CsbLMkixH9xoAkx1v32JKjxXwxq6
EyhikcdwrqsuuhrHxcr8hTQkcVdOIu+x+BXaVGniAP5RVTDpMU7mkn6Mb+FioeqL
arKQbk4DJZFeFaMl8Rn7703H1SslbaPLtb+CfEqtP5jwPyYOjEm3+v8YCuM/c3UA
s1w90ql7xperSdm4WQjgm4tZ2zA9J0jaGjjXQX29O0IvMsoOPJtxUBI57UCd0NWL
YkGX9CmJ9r07VxDt+TK6QSRBtuZivW3MeuLPFuOD0U31HrwqF+fkT3ZDiKDOrsRE
3yS7DW2jJ/QGY7hCmzBB+ZftbWYDFEPkb/tvFkNPJwQXIJqxBhE6aTLPdwAiWLW5
HZmGqz2ZEA6hSRHW8FSGhuqBel+yx7T9YGXIiQb1iZpWaWyn9rWj+yajzUnqKn4p
FaDvWDJAazaLxcXcG7G/GbqPmbE/cGoyR6AYDexykQfWHLVClWAWe/naVHVak+zo
FKSzLaOvWo9Rr14WNH1EACBJt+URDfbttBUBKswIOvHFZmkKIZabuueDBj0mIA6f
Cdi5XUlZ4jpm7L7VFR5zZnK/I0dTtGAaOLZH+QStQWTyuFJzmcqW9IQXYoPaUxOY
Ku/uDt4P4joAMv87tRn1Yce+6+wRjSd0dOX41oMqDQHX4aZKJuF9R4mVt1vtoBjU
1YFfD8DKxV2s6C3ybGy8v+cmRjoV6G7auhgwfl77sMCFX2o5mlMe9A6weOcfl20f
lOhXl0bAxmj6d6NCi72KHMUiPI0sxxwtMRsz/4Ssr9Ib1sHnRzRaSyMu59cYtSoL
bp9Kq7CXxGqZZ2FkscTsYG3iQqjW73Mj/6THDdPwK4Iuc2kQ33p4Y01yXEsPHe1B
4EdgeGnGIARETzbKgxZ/L7xi20TFxyqPhOLSJPAJJdi7swkqwqCbLMefjllVQ+W7
DNq37GYOXTYPkItD/p8FbRrw2Bi9WxPh3kx34Z5/o6fy7cOOtKTyKdnGDMSu5W1x
qCD1gwOF7b7sCepsRaEl6isKrCI6Aopm71BqcxpncAqYPCzzWGG04wz3vYVHtDaU
TgZx/3/B51vyl30bPLA2ssHXjbgDKGZzNB60u/vFr3WywrK7erphioTEgRoJTmvt
h13aeovQZ5u7kfGRD2pyRcOyVVA3Btwa+3MTKfngn+G0bI0OKHMV6C96Fr0OXk5l
JlYRnTHaHfVXjMI4mFUy3WgZKyQ1D7V4rOBfo6XOx2dBXUDgJqxeez5hlpDkGvcK
Hee0w0ng/FWs2sfFtM3fjJrlZWYLt0egEYPMAWuR3tPDEb1QbmbH1iX6hF5iFEnN
HD8L1kNgroQ/jNJZ329gW8DIuCsYpWcSXq2bpbbCMII3r6KlxJcXmeDxKbdIj14B
367cw5uEnqO2O/E6QeL6aoJ9pjYA5ei9A9b0bYuDo82g4wkF5D32g1Pn/HRQ1gzK
V3DBe97Yh3+hR2mAn4Uam6/hLVVGgXVbJu4ZFuZOEdlKkO0M1y1xHfZ9Q2PvG2Jo
bnWivI5tClgTpKREw/GendtwnGYN1GU9WDMV1VQpZjadjpS3Q3dYj7oEu04BzHLR
NJ1yBokP7A0WYnuZO/RRmVYCEk8geMqTPsJyqEF/lLOF3rWtQJjvhsUTRvnV/H28
TCsCImMgxhNdH1qmUmwKwA10xUWQbiVESW48h1mR7iZWmvFzwnkmIldjDJ5/Aa9f
vus/99zX3HpGjf9SHck8Zjcq4aGV08EoP+YVbebkjCw2k0cyaRs1ile4pcs+fHVu
GDNzzcfVaccAk2QWsmXtEZM7zT33V5mq+tcyeBDzvsMpkKFWRBPKEhyXP8f9/2J0
+Fm23laHohtPEEty/wm7r+u1DB/odgPCHkwIHR4B8A/iz+bDrB/Gsn0T3wrapfdM
Jx6nA5wRFCoR2DcvF639jR7rGggW/3X8e5trcTT0FHDQW/nVQ48Et5dr51Q9zlB9
xPcfuOMCU6Yvk9UHftT0CfyeURAeJYfW46Hiz04VWvg5UO874Ql6RxsUal+IpVNJ
2NJhSGkbmQAoD8Z7ltyCZqDo6xTYTY7aucVmqV87i61vo1l3NK+hZielCiRKi+YR
RCdPec8pkXW24sWuqYsOZyVWOAJEjCRyk/6wV7i2tsewBDp/Qapvt+ULPb9F70k7
3MhQ4O0lqgVmbAooZIlXBwerIuMYfjy738lTdfPNTtTTlDDc839zm4A6NmOInM1S
xMctE+DVKopTjZ73TFNqJHW+Hvz/6gd/wA0omFyB9PaW58TbhmEolp0ZMIKom7eV
7hOPd417VY1LeNPTMkaibppXbsHKJENNHudu1JETfvwy0u8MBBZz1efYC1rrWFST
aRU1BfF7IJlN9x7URT5ABvBnfUYFjcaND35yup1sjTeD49ose0CZ+Q8bmK1GizIL
4spMg10hgBi3Gdm3hvEidf0NmUzPSygpRGRhmPc8FoLCilJTm5a2Pa0vxU0SBKTA
BQYjt+F5SvocLokLclgw+K14fFzdZ3Fk3t+82DgEv/td0esjdl6DmYdOOYCPSE+b
8HiQf5weJIILzrEh10QNWtLKHbcwBY0j1M9ZoiH3Kkrv58/GHudwfueJvrOlOlKy
N2423K+0mGI7+FXfNJXbO5sG9iW0C1FwzyIxhoc7i4ParGNzPtI0aO/61QQ1h/CU
YmvhP/oFBM3NHqt1VroIfPOLj2T11Uzc5YnpIA/E1jAKleavz4O4cVZLCfXQUjlZ
h631S2o4YLw2rdLUvNQOTN7VSmPV2H9+qW4CIieZqyTXbAP8FpVZthNQTEtK/4NX
cmNqdKmxphxiQzqbdbpmSqL8fAsR5XC1iUjcxbq6qk/Qs1fZ64rQDcaz9g9R1zaS
9Atm30AkiRGF+2mD0kt495RFYufO64nCRM8ZLnsxns+5xkm4RtJu7sSwD/05eD4+
XtjafY0G6lPnIpJn6sdSvFL0kMhhsjDy4/8NAiFZYY8XLBhjroB0B2qPq0Btr9gs
6+wCgbf61EXCbercr8JAfJTug4Tghtv4kfEtUWNK5/iWJGjAYaGVeWNSYKcKUdLv
gclK7mDfLnIKzMxYbp57KZzJzVKm+wNqW3LAbptZsYX18EpBkmAXsIosu0e7S29j
xgczs5gVmPxnYyEo+nKDl8D9pzT3qnrj50CbH0Ry/mCdQj80X0gTl1sHSJdTF72M
eNhg8jpM/c9cORLeEEgSs/ah6ZloYTAt04Dz0xguK4sFyKe4NpUWD8RpUB2VRpZL
rV1rMppscjr2M6JF9jEDG88eznuR3UthgkwsLxEDVyFMxhGOlvjHZ+B8HZzt7SUj
4LFo0A+YiAg8mwjehqY7MGS8xvWPdYTd21TI55WuvMs5aYjJstrg8h2nEBusb15X
cqm/pyTU/sORV7i4LPfWuU30KWNM+qcMRRoZ0lcvwecTCdkWHUTa+XtCA9S6Lmrr
pdv7d2vUupdn4Uqwn7Gbh7/+ThiHa4YY2QK34/R0sA4NY4nM1k7CDkCIpfetoXBG
dVcUAJimLdY01+1F5scPZOTDUqXRuwKyvAKK7yoDQ8/aapfP7rqni03F4Suv2ZpH
4qByTCzAioHjXDh+cVIGih8pLrpFgeKlltd1D559CQP5T+CRZXZtT9VajO8jrm4o
TKismOwTCI/VLzc4ihVbP9ZqdhDPLWY9qUZAAkb2xbJFnMqV0mNjXj0sqLUjjjv9
pyi1rjSXyHWTAD6Y4NNcrGuG7mp5P7bJfhuU4t+ztCcTyC3HAPfd1Y5wdKz5fF6+
QXKaaUFwga6SCR8aNdfTiH/ih3kFxF2zqXb6sWodI18qTue/kcTlSqPtGdxYaWbX
JND0/PGnhDURZRwtpsyYL+JL5C6xQ/C7W9hT1ooh3irjsAYN9+qCunb2FhYCMXmn
oXDnhZqJYaOFigDG+qh5bMJbAmkR9Es/lDxBLOj5eyLZKW/lB/ttcUSNRYRgYEDd
Ro7WcDvHGSAVs3u9870bSIaLwwyTGMUiamp3ecujfuu1B0gGAeuozwdr2r/G1fdI
x/7/14cGOZB2k4G9MRVzopXgcrFS1xx2nS3XthGieolYFaoTFZWxc10J3x5cRE9S
DBye8T+crZjaNi6MaRTf2MZQnSqF8UIZKYjQ5cxGxp3rEAFHole0IL9KRC2exi4K
VcMOb9++ew2VlLT6ULUmgCW/YKfCRmHEDev9s44C5JVJ2HqYfDU5kofjmCCNnfOa
tgCOvzhHrQTzUaMtFpUS/s6MrEUb0Ulc294E1u1leJNCGEaIm1LUWLNrk+0qOKTq
1AlGwMuQagayON6P5nOpTYbTcsaG/tJWTsXuFCBEfiDj1MNWDoLKlomnQ7GkkPxj
YSAjSe016WyPZ6k0+fUCtz+UgQPCxd5NJTm/M5sobW9Sp3tBJc/mUNP5pK8OBT3q
FMOdw9nWVDy6iS76t5xz3Lh42Wjkov7mhtvJw8ayaWRjazdCwWQO/AFrTttewFaL
lokMglohbSHYI45muOd5WB7uO1/GdPRBoVGQuDhTpJdg4dEzCha/Avndd82mKvrQ
i5Rk5+OEvKdHepB8KPOkMy08Q0zHRwNjVtuMmokKzaonNEA8+aFpEoVpfCqeVniT
OWTp2Rq3NgX9wIa7yy3845bPAKAQhgiViCanjvkHgY5kdeJlYe3PSCVklGIrIPuL
tLeMbegmxuS+jYr3tqFHO/6buAXXcZ2bgyLmm6HOHLnbDPotlVtbDxBydbsr+Mu/
IQCvlzwDK6Qlwrf5tVSqVpqHFtyvpJLJr5qe8t+NUZi4WVR8mSJ6MNN+xVaqNTdF
cu61q2bht91raA3QrWSzAhYgm7lM3/Pa37qkTw/OKRMSKwc4nHVmxxKCqRvuXE3G
OWiU/SOVtL6RkTxZyls7Ly8Xre4Nqm2l3sC+REXUZRFQFtuDHMu2jUM61U9UV2C9
AQQqMLX2LLqb/8kWsx0gQ3jGIoeC2uuoiHv8qoZeUsCawEiAl+7fMOdTdW9+dtjl
mNmqrX4KRP2LR/qJoNKOOHTuZ1K08QY/4DNU7zgEiAklRI1Jcdf7OIfvoLa7vl+N
ob/W7SIcpWcK0i/Wd+IEE6I7sLKY8FKp54d5dBnbASU4xCjMgPA9SA4bJT2v95BH
GHvgk0iAL6leGoJ5HWb4JrGUqbwVumXNIdHAJlafPFAjw6sF29ok89Jnxk9QHw/F
SwjO/Xa5+a/GcPy2TMM+vgXkOdr2VsjTn7hnVkGmSLowzGKax7RztV/ycwUJS05O
avv2KKup9O/vJTbbpNT2MdSMZFToHtPPqNFf2B4sx+yPS3DgmE7UuLFR4K7ICVGW
M3yi6+7YW/zJUbs8HOl2THUPA+9R+9gLHtY15Ul8zsFn5QUnmQC0leaGb9FadJA8
zNMZ+8SU04C3Q25H3wSFuDFsQG8voMPZ0EphSnMYvUNGQQNh2Kbe402eioNuPU1S
l7eDgpFEMTdoyQmwXdbkq82bpn9C/HGyNrIRiRT3niz1Gp1p0SvTYk4drwTUwd0X
zD3MUUfJJXHKOnCKnu0crRfe0dqxMliJ6by/BTLyprwaqnF2M7SIViLRrAkxtRWM
sIAGvr84YNHTZB/MGyLtxt2Mk4LIJfkcA1RLWkMUpDgjxDEDyQVY+hma9ruMTO5w
2vlYYEhm3HboUruInVfUvJFEfi0zTVoUifHX0sPeuuiufw8QqvFE2SqNptxFTtCD
IjOIPzDedldODPeAn4p8z7t2aqG519mBKZE7z012DK5qrUjcYcVf3rj5ReOzBd9i
TZXaGMVbzMmfq5tRM8rlDAvrMkS4JneQXkJQhAj8hxCbzkkdK+w9XanW5Sqj1ZWB
BN9ud4VG6fEvm6sE9vSrvr2AcV9WbfzuyuhDHksRW40lK1SiR25TMNz7PZchyeyR
OmxemCSUceB0Y7wt8YoQErU2b598rzXeDtiXKwtbiYhedmo7ha44Cf4imVmfBCxA
WJXhsWO6uQqhXMDJyBZOqsNOdYXb5TEOcPFBzWaOXBx+fJsvJK4OdMEVO0M5NNXN
e0xwqHaxSwXZnCwccx1ZlVwoM7xQCgOMvwG+QNz50GkfOSbMoh6u1OYCXpKpV9u8
MAXXoPgOOfbOp4q6ZQfn13LmsxvlpvANwNGbboUtT9GcpFnx3Q2ko7gYty+/kDSc
I82yn0Uw/gzhgRYox6oP34+pQdeDSXBIitQ+bktJSxNqyXpOfDxK1SS6mcWm9XlX
tontzznpxw76ddYToIPyRoKDuaKvMVFvqkrLU50YeEInO7IsHL7uW6Mt3R7NAn1o
vZifqv8krBIcYuCKKUSJeO1sPlBYMXE4CnlQXhYLojm8KgHzy/t94vtW+fxFuJVC
gvWJFoCJxOMjBUjR38gtdj/Un3Jv82LDjpjnieHcYZlTu8VgAh/mAZR9ZexyJ81o
cl96xLDPI1X44K6TImiaMGYQsWkVaXhiqEnzB0jJ2VxLR8kYy4FefjllCI0mwicK
rxgvy9luulWZSTyqEnISSfL0i8uKra5hVpqfhcfxcaI9QmC93XLcGNi+4ILmZwnA
jwVE80GPHoXVB7h9BzZQDpZZOfe6+TKy1RBavnbs6ei/fhWF+I1MEuTixo8GRPMd
ysd/Eb8zmE7/rr3xr9QgGOwIGr1AkCH6TIRens6fMo+ZT2wHzSJ4Wco6TjpRj79Y
ELSAxXMMahlqud5/TBGYmVzDrdHpbPhONpVA2k08DRDbmnvL8GAkvIuQWPm93UCD
4TW1eSRwP+sQrhjpl7Hvsz1AnDzb1TEWCZCgctgP6J/OvLg7w5EdovMdC4utmrqv
b/9epFXbvtkY0x4UZ/VwrKSHHlAAVSyruC1gn4Gd2/QfX4tUPQR4XpACVsZ4wnUn
ZrkxL3bmMIwcBS3iYwIhchkrUtTbvPSlEWrvLZOR/wMePWfevL4TBbsTLtDsrkC2
5hdX7MIhmfk2sWDTusnjV07aqTBnZZR6DvzNfDfcLWDohhfEIGlTjlpqwAbySQZx
fGi8MPagZ9Eqo9EXqqFFAx/vToM1nFpbi7RQx7sIrFLuIqDIyVcnfE1sv04+ts2G
t3EXh/aEJJNNqB40T8EIMGoT/DSjXjDOZ0ou8FL0lbLZp6P8BPu7tLDojNCb/fAJ
cJA/Z26oNmxlMRKBALWNd+EmlykL2IQ4iiPCr7Ll6syjMGTcXjCTOYhZ98msHYZM
dpxdps5xSxR7bszElSfasfjgSJCeQshUPWEO7+X0G/CSPueZO9+k7XKuV0a0E+c1
ANxiswYyH1TJUwLhajUf5sR/ft12m3niGAk//sW6ULove6ow2bDuzF/7e3ZWZA9Z
biB/1QSW0geZH4eWwneDj2eI9KVXIXv4Vttsrs0PniCi7qzF248ABbpRxD3ZbzK7
5NlZdboLru/mqJobPNuAwQCtYcy5rvfl/IGekiz2dnTK/+p8GsgutTwenG57qGO/
GobVxblZ88R8fjcZzyxbZVRChjmOG1kmgkYtnqyY9m6KuSRm4+r5H6tKkZRgtSLo
r8UyRURDVWetj2UANiy/CFDOxoBsa0ZOtyfQQR0+IY48plbE/odzHHTiDr6/7UY0
BSUWmQz2oXM89kJVrPBjxELp2cq4qO2kF7O4JmvImQjnFJsokWXPiK7Xpcxxx5kq
6ltuumUWp1DniYTe8caRajd91i0EiDngLCPR2Re1xGzj/KUXzAhYfEUovy1/5Cvv
ih228DaFAJrMdAtt0R5l9WmSKAdH/Jy+Jy0GH1d9Ai5uL3MtewagNtVeDjVlkMPG
+E7nVcAiSyOsLNuoz2gq2sOoYSrw7yyQ9aKs5wEYXafxIlSn5ScP3nZeMvv9+zO1
76iTPW3ge29z1OE2hpqI1Lw2neN0Mm3j9LV4yUTodkCNPUbarx8rbt1NOKrYWKa6
YqnXzVpKnTWNSXT1HsnXVeb2YFEEv7gF6ietqSLwEAv+fCl5aXSm9k2RMmGuv1aU
NUsogMz/CEYnzHt4+tpe0MMPCUMHbCTVSw2Ewvkudj+axXouN658789eXfUW+aE+
SJIUaCkCPKF/5Isd/4nencxbanstX1lA2vsL3GJLlW13m6RENhZT8Rv0ECj8/Bsf
YhlFpvZGwxRE63jYp6YuJRrUuJtpb/ENiMbxq0CNmCiQsWFti+wjQ8CkqFbMoYzI
igUaA9li382ps01DgTGR3HwJtnkygWH9aR/j0l00SFVhr+OuhODS3oxRhj1ipye3
K6qOYeJ0SnWcCjBbQmQDG8v04f2QlrY5nGEMAgV8kd+9WFUlGwJZQwXMhemqJM9N
QyQGqHMblxBeVm3k2+tJSAayJL9Pt2iHl3rG+Z289eLrZrRLLVD/nT1G3MZCa5Pr
iJOaLki3D2W6D9F1uEwnZfhOL6envl+HdJvRawHpfkE2cCUR7br+hNesmeEkweLL
N/DNVdO9ir2INwSPojBhCvLFETdxMMKfhrpnKyS2Lo6lAVvRE+p1iuGPVe76ivDe
vp9u3Qvktm+jivQuKiH7eyAmhknojWDNcd9G3+vVmzIlgPL4O2mTeeCTb6HK1b4M
Fw6SpfYW3wDzoFVsER2WMWcBCKKHN12Kk2IETPgIhcWj59btS1HLZaBxps9meGZ5
pnvt3xm2Xp0to56QHRqdAQbzl2467ZCRQc91bPlax3LYDD9dTizLAbof3Q/HGFi3
s9mq6wNrnsjIC+jeg8hgx7KQWOPzY/+wOy6tqXLm30AtJRO+pYwFp6iykt7ZAdeI
h3X8MoZNEzvDN9h2jKSFmKA4j0oTYXSpsrh3kuj1Ba2PoSUxN/zvxSyygNMNE3Az
Sw/R4TX/KT2MVDufYlrcEJTzqMVDFyJ+7gmIsIKs3lTTtewQmIGqJOwG3hjSipiG
JhwAhtr+ykzGduvx9+PKcCCUOQNHm8wUBURKnfAtV6u32W/3JpeJ4dNy3j+IQqs7
5qM4mQulX0Q6wEppy24OSYRU8hz2AvgxwfueYI9ytrjPgMWFOP0cj/RayhOfnlbJ
so7UT6jjx3Q0aWzm0+WCCqnzpbGmbpXks7aR80JZQ8ZM69M75tFwgjSplZIHedwW
7zolDffMWP4n2M+yaqz60kUV/gGnHsvkIbRoD367YgBn6HnnQ6lVvT4IAvTsv508
5D1rUC5F8jQd0bCz3V40sVysIIf2gAvMMYpoWYGydWl1rjV+2ZMcczTJCOr7gSLz
ReHdIU7wKHO1HH+OJniraW6Rd8+hbs4acKxmciEYYFvDtE+lCVDTCQTfXLhhaRc8
x9Sz4jbM+Nl5qGMPMOqWqwZjtbIioFNe++zjiMwmv1QXLgBULj2bmcjLPg7B5d2q
ASxGAP8R6PmiiZhrH29W/xcjJ3pZsvbMjr441ZLJ79k3j9LB/+7703MATY8LH/XC
99RNCRnhncSrixyVgmfFNDCNT0DXWQEWXl20zqTav6QkpdnC0u8rHVg9CtMN0M0m
gspypwuuOwU6zPTe0CGTTSL5tz1eyi7Jg7sWQm4AR80RHgyUF3ILO/KydLX8Q4SL
Ctj/6EEv/qFodmjC3ILYmKichrCxrBNBzZpWb7FF+6C0fZmMQX9EvK7PALEC+sdy
M9MKPetVo+wuxt9W1ViKSXGpe7JdsjBj42nk3dSsuLGsotfmoks6jsOqvCGY+HDd
kyTsP5oOhaqbGnyL6J543uFQopp0qOFbxOGeVv+OyJgIT2UfUGS1hER2VlzxaVhj
GtC7zulju13sApzwZitxe99gBNyZmvC3G6H2xBeA8YrYAI/qN6puwvRTsZsn4I1W
7b5q9h/pNJGzzIyw1eb8722hAUNFu4gGZHdfYQqr0m8mLzeWwsWmnbzwot83xlWl
R5I1IyYY8uTcgb4Uv+6nvDeuYD/5ob+0jsP6xAeepeGoFouDoElHLW/CNksL+LLM
rEux8AYJfCjb84COsCkeylhDsxuA7MOPiEfDu6oNz+KPHCMtjmCtd4ibSKOhg5gz
MRDdEQccAb3frYMMKAUUPhVFxJ9fIJZActhpYOJbDGPIgYJzrPfY/LTZZYMr7xNY
Qi3Ncxln8l07RVaohLeBG9dHRsqB5xi1rOq7dwz69xP0f3QkTMkznKgD0GTjax0v
E+AS0zP/zedRFe8T7qPf56JB58NQHvonfBbUekAOh44UtZt1Ie/TbONKGwqw05wh
zN5+CTIVZnwGEb5Ff4K5SUrRCaOWcQUhdV3Wy92jJfa8MbHXUPC9OqcBcc48JqIi
SWWeWsC6z/EZFGh0Ot9BrJWwMW2Zv375uzaiQQEp+b3l2gecMKFQWjepxf7vUkB6
HQHWNMDH7fm/QKovX3HZVzlIV3dj3HLm/ZYUNemmnUUg6duU8mvRwlqcUs0Itsrx
OZUf1JTVCw0aB4FdnVL7NhjoUrLkHiypWN1ym56FDQ7Vuv9Lb3XE0iaZp5nC56bn
ZJd+fuiUclEdZdIRxVoWUizz4yHz2Dog5qSVtbT275Rs0xJLLWdac/a+5csa0+SZ
9u0lF+IZzys1St+5W/xV2lKIESZodS5B2Wl/vVd/TOu8xbSk6541XYCpBwdrtKme
Am2jlFLF48Aua/SAToFLqT6tLpq2Iy+kejmy8Ai4Wktd2dyjQ6fTvkzc+uhXcHW5
PGKYK8BElHlgL6ecwSrFovtTnu34JxeRZrSanw5QyrNfuy89cjkubh18zqpx0BjD
L0GcnIXVIJHUHUQlFumTDF0VoXBFbQGyIBoG0oweOkrjbPvxQk4qKCfgxEYwFU5N
WfM8bn2xZ8YRK1UXnBiOr+lKrldbgvG8+ByISCpYtEIn2eKB937lAzA0fc2fqxSU
V84tlYvqk8w6sGLgEgC6CnoO3yHWXgH2Z6C+da0EEsQgvAeV3yPlFhTT6fgQ0cum
mq96X5ALSq3GKc2+P8AZ4xiuoN9IWVpspqKjSU5CHlePt5XnlCOyVguCQbk8wFLK
D184l0A42BUH1Dxft/A22aHN/ESEk4c2IGpaccDu18F35gxIEG6EBhHko1bagXPq
uDVjx2R3A93Bd4+EL9ub0Hh9xKCW8w+20kSla1RRFXVGdbR5SNVnYf3ioozJtgyV
xWqqGxXcw8IdC7gzNabF781Yk3c+wrTIqOYWViW/KSAwBZ5rTt0anfagy6BttlvV
OIsf1+e5kLp6cXc1LgsipLsb+9dGf+7dzlAifXJBufDrsn9GzZ4HHJAfVGskSp0q
2gBdxAlql8mnc/J/golHO0P25v4P6fQ0jPAMTEDHu8nAil+EY22tob64yqrJ6k4X
A8kjlOr2/EK+FrRc74Qa1OuweoK3UF5VZqwu+gw8B4m8x6rnA49DSI+pwOg1sh7P
HC/ZtJSzy48GCfxy8YrgbdyEnTe/MfcKvOTQb0PKM6tf8H8dRTDqGyPrHAbRqjbP
GUByQdc5DbyAp6lTe5CzxfpUQLfKlHt2yktPNuzs7HbuorL4VTrLMcfAtkomohQ5
ZQiNotS7KpAjLyXM21rvPb/Ygxzbxug9KMWe88oqlq85gYdCfXpcBwdmVpXR5hal
FIrNjZreO9PAyxUUjrW6RG7hQzMAO56yqU8703R1k1/UbJxuemIkIOAD4FRj10QS
tZiV753gKRnbtfXc41MSfbOA0kJGLFuHS3bVcbq2YrZKheevO2wGqfgt3SsRm36C
R9qmWnjJC/urh7AsD9Spr2KvfzdKI3oIYud32iF8+GO75j3r+CFH7BvF5C0Kupus
kwRrcffaugz5Zf2A+1F/WYphtho2U+KL28a03QOMCSgmKUPTqcrJ/q8/CFWAU2QF
BhPFhdwk/QxS7ewerNiryA/IbUKYZM/tVQW8D9csv8lzeDzOdJZS5Ltd7IYQyWjl
NK/ASCN+hOjUl5iPN47BEk5HC2LWe9n2qC8KdbzAdlMzpOBxPohlasjgqDS3GM8H
a1ZvCmaJUxpAeebsMQfDoZ4KGzLJRQIWZjGbjVdPXvoDA2M5OfJFY7E1GpBYzIaH
2kbGdZw4wuqrSdQfqygwOdb+FkQt5hKOHAJ+YD2lM5IoZWqBoKLJnTsHEdEaQ7Ki
wvfigS9C6eSCJjPSNqFHBGc0saSdH00dZ8edaQS1ckk5j/LloCNNQ3S5BvipW+Ro
jrdxwhTj3LNh1WLh4aYVP2rv/f+c+x+hUHLpYy77+2aX6+U5pcPb+LPRNU+K92e5
26JHg2e5swo7RDXwzXNuGfSB5l4NF0gPgPjl60mNHnOR8KJBm+w413AuYhynwWBJ
/qjHG+RmuVBiX64FjwhpcQK9jZwLKfx9Y3OHyqU8HRcDq5uU2EuLR8F8libN3y3G
uEwK9rK40tgEU1CgP3UFhByeF+JCjWogHRrPxmtYilYJDx5DR8eAKpxlhtPs0pfc
SMKe7fhxVB7Ru6fRi6eHMeKPL26u3zW4KJRn6WZnV+yBoceQAtyT/mM46NMCwlhz
ale78a/DLsMy5RuDJH85bQ7NAOSoIg86xYG1S8LDmXBY3B3Ce6Q6JQec3p3yvPIw
BncDoqYqT7YdAKzAQX8XFlr8VFnlnl66De5lBXE3Gjf2AY0yDnCLnqvjV21fCh7p
6lgClWQbM09XDOPD0/UxX2JdABxtZ3hc0TRlZrDBVaccc5J7cFbkNGixWI7QN0wQ
uU1uye8IZCvgu+hHshwr9bDUJUoSjuSN5sKU5eX7Oa2OwDIyIGaI5k7kEkmdj/3x
sqvUYTiehpv3KvdT2/O+0lGmZceINjaNAg20MqCcJKiGSXhT/ialskYZcyXfflxw
BEMvIZFw6TlFdjsy7eHxfHNJa3xo/JSF5YRnRfkJfgFD4x3Jk3pJrdSrKk5xxypI
96TKB6pdL4fRzD8wYIr8Q0O6r+9Ok4ia83JTKrVzWU2I5C3jh+ZrKs2p7wUVNELx
Fo+53ddA+CBix0mIVkTiU4QPImEtFinqJUf3xMECJOOb3QRS+aK6LVaBlIKhirrd
3Wq/FztAxIKhHgRO6RtCXIDl2wuL7gDbNCJRxGaEnJw1QHfyY+dIK/MyzBHQHRVg
37p9sAPKvAUITguVk3wMA3+nA6YiGzo9p9qd8b5DfVwS1dKjTTRt1M1d4dIQOJne
GUK1zsBGEYyWiSApQS/0WA2twqczvIQG4Xz91j/p4BBk00Myy1Mg8/PtIOcppHbe
KD8YLNFTuD4Lv/4ygT4uRxzP0Ve2N5/aB72+gsY1ZJnzfK+KQBUcJNmlkc/tRDUs
cXyFK7I4767OFneWdbJdbDnAqfChZKyjqmdkr3aC1Zx4lhp0E65mAAjC4CZiKqDY
clHZTP5PZ2hWeaawwfBnGZOZ5+tTQOkQVfxUHEdfDvTIN/ftPkxvHAWRxW7QjKb5
BejKphVakAumSPMwGRX8IxshE3cYASyV88ln6LkQyf4Yu9zCjw/6crNAkXz8sh7H
0WC2XmeqV/Zlqcf7jx6u2dt5mh9ncBqhMI21VXSDQ9xj3jYVH/+ayZgJnlWawU6b
NHEdpN95DqG7vp9Ybrqb+i/k7QGnOehEj1DuAaRK86lyHUHyap1fPPC46l4+SBiA
qsdD5XJ+6dKVNH/7H1ieQFhI9OUth4x9IGKY8+qNUtPbhucmcmzSZ8E7mYf9LGz8
XaA0u4+7CLbpRmlDUKHmmBDfb++s11Z+Rj9y+qbe5KKf52nLKl8ijlQj0q1zjG+W
8EmZYMdMBljVWoiLVMlqx42yzddHc5MdURcuSr8zH1q2SbYdsVBYNGZ9hGiozYPP
nhspuhR8bZRrAtUe/IPWGJfvWUATnDoRO+L27QIycw3Z/hUZwzyVBq9ntx2cpELU
WD3qwu5wFn4lOh8e/w6J5IX9mPRh9MZhSkI/4MlvayTy4rFld15Riwyslc8KTwob
vlR1D3ynbv3eqwcNI5NxFm7H04cTC19CjxEMeczey7th3jyEwrfR6REIOswynKhg
nmwelEaeEiR8h2HyBA3vmDsmfEPZtTLYpLmUnids4WIRgJ3RnzKdzS39aPK0mdrA
+YA1mZYjiEh5tWkm0ILvPXFtYgpWDFZOF/ijTMCGokHLSMPDGFC4XVBT/D1CSx0K
uujPT7qGzk2xmndfSmebQvyjW65Y6yRn8/pjp1Drkq3en7lDjr8/TZSGkcHNfsSD
tyMTmx+GqI+yVhDGGlRlH6LDEuAeW54tWeHHIhx2xsggKGHfa9hV1yfMRp3Q7e03
KdKWv77cktufpgNF3gtH/iH2Rdp8OhfD1yMf+/K2bN68v5T2LXil3/TWk6+qDril
8nog6+SoDMQkjFg0bglbU/5usx3JIYMrLqy3TRqY+jf+Kup9YMOe3Q7qHOgrHfQf
kv1517Af4mfDInsVBPthhqkasmHAtGX4dRiM4JZsYNpy0RIsY62hlSdFFqkd25fp
GqV7TzCom4LHcn60UWwiUHnMDs18aULihkhUNhk2XemCf/v7u+43pa5gYuAApDi4
/aGkAw4GLZS93KLOfvTqDMun4nsIGnpmbzLnsA0wtxv+tYPnBQTlLQ0Yeq95x7cN
XvYyeXFGBil8E6eGmE/bpjTjFxBIb9wrVAtGT/LPOhUj87aK8eFhyvxT3ji/5jYa
TYEnCdTpFMPgbdD1sTbnNZVqculZ32LVeEgYd/87w7zdrY/86qKbfICI6QsPkiAc
uhyLHkUyYD5gSZP61XMYXxn/va+HTk85gb4z0l5KhCalaBYyWDXy9fjPDSPPTZIH
lcBg66n9qQ+cWX03rzhc8tjdbm1BCdajGVcGzVtwbUYL7YWKH3TLVVG28ZG9/g5e
Z+cWBqCUQMes8Mk21qdivmIT/v7P+xxsgE/Cwtex1HCoUYTJWKgTowamTklzUNbm
8eN/6A/Bizvv7hozf+ZA8WpVzmWJgWgGXqF6ZKDMUNR34w09zA1wcfNHhGlu3OMr
ULJK3G7qqSvoXpW0N1nrBm6AeEbu2DOakvauLfFjcKms4xNU8jL3wNu4KTBdFmc/
KEqOKeHyURyE+oNUIApji/C1GRyDi+0rp/xzxA8OHFxxto9W63i4WImLlOb4GH4e
a2Nbj8lnnzO7L9Nxvv19KmdzBEbB/yx/vyemFgYZBgeDWrLrgJKPMssUhRTQaR/D
hFG4aVF3plgp+Sc+W+W4ZeDPyYbFZfgAX3lAOyJ2GiNEie66PUD1affRUbPkHL4q
pB73K5yv3ndUZz/MoDs0q9OWoBbRywbj20ts3jPC7vh0CvMIuRpZ6SS50+PfhzkB
1/z1HNkRIJ66TeUWfVHtiNSP4xYzXShfZRVnpEuP1TgV7kpQIbHtGpgqj7off8sq
DqrqPX0bxKi8qmN5e9xZyDgioPwCEFft4bfJ93EqPRvwr9IAZX1Dxem4rH+xACBm
IGndJDgPiyEm03mObV/39SQoeZjO6n2Ho1vtLrQF2eCCI4eIyNTpKshpewnxtMYi
2XFhQQCWSHdI40zDHrffH9NsLJddVy7Ax7x1DNYpPFG2AsaT5QDclA2xG/bjJl4D
KtGyyhheOe6+On3G74ESG5cI7X8oxcPIFipaQ2qb45t2/Iu7bsHChIwe5sUSgeDH
RJm3XwUPxL92PUC+gnhBfdBDDtcC9paurhuxtI2AXj7gQyZaGa0oCbVPOLvDcDJq
nKF5p5KER3+sDH0lIXF2sIm5PHPYJ0CpU8CIVgQhqCD+NXBbOZtm2DDzm+EaEsNS
RDNGYjsXQCYNC9yurz2YSFCaiOFUfZpbNeusVWxrDsZQ4ai/WQzgSrCxUMi9ga4z
mN2i68XVevE31/62XgqR00rMPez6yrCCqeafcG6p8aOXUKbMEHWfF1Y6k2XHMP1i
bLMCI1Ek92hryXpF7Ee/PcIatqJMZ5G6LCDIL4toGPPLtLUKVdQJWVNuG81mOhAn
U96goJTwJk0wLMGy14xYy0u1dlSkCEaEsPybD9z/hfEXbVdzoL7B+whASDDAUK6l
TRJCyTIQt0Y1q8ya6Ksrp0/mKUdLvRTkKyWwXNQa/tnMQm1Qg1toibYqE7xG3Iwl
QkHSyv53zCKdcrkq15SW3oNxzIguxlsFBZ5F93KY5C6zPTkwbR1OBa8er//3FgKa
EYdzFkiaFh+S0xtBWGbFSybD0pM90lc9PzsDAoh6PN0Z7FTsLd54lXSJFwD/m6RC
35qNWWadkQ0bT0VCyjo+u7yyHcp7rV1+0O4+CASzVX/0lHfUAQrprWT04/08whZE
nHrqDu8TvQNTdzFI3y8qlAbNybzAWNWdsKIvQFR3WIgJqjlKIU87kMCoogR6rcxU
C2F5Fez1WQoAw+g6xom/jnan7llKPZB0JlPznoNX458GFhuOvk4+lRF2mehVF9Yx
Ensmfa1080P7XxmpKbNz65qQkimhKHhH365FOdUBNLtRBXN/DWSv63YJfEV7Mbiu
0LbAegco09kaDyN9ht+Rm3vE0MCyN58FNBhLTDBx16DPBzRQF9IEGrUf/Rfj4FjD
ERke7EtPARdkFbLtRsfNE0vE6C98n5MpAbzwr5rktIYtevyGxFVPzpq1t+Htce/w
YajsBQUT9P2ByUy2oiRGsPxd8ItMTtZ7J9ycfP6F5PovSovSKU9+mzd6bbfdnlui
f5ze0zhkU6NJajPz8T2RrCtXYziyQd3bhNpTzDuv8XeofxS5FMmjICucxOOZv59t
/ZTABlbcg4Mo8Dh3c52k/nT4ZPosO63Ww/UdyXjcZmYfv5QWY421tF42n8vbbrnE
KoNI5EpHPOpM0Vtp6akno/5I6rrvjv6ihVH1IR4mZ4oZlVihGPs4ooRUCuKwaXbr
LHO8iJwTWuk+oIB5hqbOzqbVn6AXPOE9M8GPLHxPQ7Gpz0ds7SxW1f3vJjx53sTh
guCLj6QvO5x8zIs8QgXSQVP9RAF4EcUoXLQ8HfO4z7ivM9kg0rLbdQfhlGfk29pP
JRPx8BSY5ZqjPhCCo0CWjllPaIlarabbK/v9JdH/YpN4IPB26Tu2MnQ3U2YGG4Yh
MiPrwygj2xfIkSGpfwvDBRQBbKX5LKn3am+JlJOeQAsPGZvOYZIuXOfSpGxPvUI5
zXsmX5m1TPVVSfqP/9mgHNyVw2SxbrZqVWNyk+rxtGh3AAfCx55EVhxA5Inhg58E
eN38pAHVBWVmqpTgwfyTz6A2QcsI5gGHqoKiiHX5Po9UgCP6ytkFMDZg0gNbJIEi
nAHyD0ZvYUqwNbPq/bz58b+LoCZqkZft7h2g0j9IBe2pXw9JAXNEP7aXK24JqR3f
7GLS7ioeRdpep3EY54xIrWZlCBhoFAL3Tl5FwluXI9ipXFJcoJNiUjlwRjL80ZpH
1iPCKpam+hcbcY2oWyWJMieTL6/DbYyPYXYfa60ZW06rpSF09FEgdWqMLpOVox/0
DVvigNOx0RoQs7ooJKR4f4EA7dLmXLFRdqqojREAQtpDJ2MIuok9ViGgfUkzR1A7
CrdAG0wi7TffXLWjxAmSUUA4Rji5sjnlsR72y27hDsBn5yzo7opqDALXdgZVyrTS
VGfH/jxcnqg6XNMXQtoPuV5kgqpuFHwcvI5+nbGWRt0csInqp0sOfL77/hSP8Aq4
O6L2WcXKCZtv+gBab1zXN23Oz1xC77UPByeWurcL3lP89efgckT6XeU4fDy5yW2H
PL+2Uktp7VHXAt+4/EEBpSzg2SiQ4EYq1UgtYaRJBrlPMPtbykM15kg0a/5KBWYT
lyYUhjAbdKBmfIO9t3G/J9uCNAKzZciWzo52jX4FXmRyPnejLK/4PAdCfEV8qqL0
CRamJ/cQUOMWk+0i2b//N5REt1nJ8q3PFf2tEYLGVBeWdIe2GaFxsiGbBuDwRxhM
ZEFLNKThkiKI0JXaC7wwNai6GZjLZWucCjF8bipoeHSJG1A5gQhBRYSR0E/4m/wq
tEd/Saho29ywFfa1SSlv4XWjwFtBVUDWYwCC2dKtDtGAn1IKZ8e4oS5uiAH76CY6
mCwWnmwff7/fDIVT5WwvFcyP10QckvK/+rbfjbXu+Lgf18zF9X7ufEbTSy7lCRX7
PQlhQc3o4IZKP69upVOIiVWVyiait0Iu4ArKFUpWlRec2GVkl0L0hbHCCyiqIbd5
3oq8irIzRGDEJyf14irGJwxsOuiE0VshsoIRFPKacCAXZGEk2fc49t5kktEeDhpK
mFAm9PRk7uWHykVbt0uUG2XHUL+BM7LpYs4v+XkkzmOqco+55gkuQLklabCiA+B5
YfsFucivrQQQN7AbLplverWhOYLsxaqBR2h4tTAutT6k2wJEmz594D1EMy/Id69v
FaMPRojcauY0n/LCTUl+6LZ/dfDfGlyslEw8orjOOJTtOIBRN147W4p/ik8sC+N3
EETGKXbYc/b3mmzlQS5eaoNxuzX+TH1QT+RRMnO2VM6vM02ctlC3k4HkF5wIHWYQ
/2vCQNO9FwkYb6I4v4dTAxZhS09JKmqf/o+SUKZHYEK36A57Gz/WIVXn4XAlKp6w
mfZ38SN+I7Xu4Q/1dXRgsCha8NkVHvwrmcQx4W0+122biez7FUEz8hAgwVpbER9Y
C1LFNAzTLUtifR2NQaty2GVnAxkHdqvkYutZWQPHFOEpzhy5qhBGLtQ7qDfSJMi1
/jTVL7z0sobLOPQqJpg/wgA2MSVZQi3kbBFBI2V7mBNJHL0EuXiCOubGv8Soktxr
zlD0rJzKB4RWkvMrEPgQyV/HmG9/yBe3FrQMNPzVnzCTe+QOUMAyvRHsP7hktL+n
a/oPFyppfVYqf/bsOcmClpKBHzRPshIktDB3N15uRGjDfnbM4bG7LgTmz4qBpq0m
gkACSyH9YLSEa2Y+lnnj98o/v3m6TEmT21orH5id29L+dqTnVdyxZTJS6cP81khL
wE3ozOgzPnImiOCobVytlJAZdHoo//K6wR8JAaVYcSFGBYoe4vXzvcDiLatK6k8X
tDcTH4GFOUfXC53aJHAdCJL/IWOGADvoCYJPA7ZkSIRWuMcIpzj7NQCntFzobph5
2UNrOT1xir03sbiahYvEDLr8y0f9tLummYJbpoWSK1gvD4BvzvdFChgpPmUxuzgi
0VASQ66SGBJsPPzPZQeDAQalJdC6hyitQ/8z06wlYJIbNZ8JvlFm1jmarWFmMqCp
iHKaOCFVSQ5vcDWlpLHI0KekAT5BDHXi6lf2aB1GxoHBIiOSciluMZ0VU3sWgDpf
vN0WH62ufJ/ix+4X2P/jqGHMV6pvEerfPMc8M+K2H2b/YobubQdvUMSVv2+vWTip
nXIZTSGdVL2hoYPrNiOwfpEqMZYOv1Eqm2dL+KTnOy9rOesIXvaZicyVXvF0xhJQ
tRkFQUj5oioM6+7tte82FSWC/uEyUZltudLo6hpmwjHzPmHvDmVKSH0sgTkZGAcq
6l+Mhr3BJ6Od4o3B6eo0QnQcbaSrUtuqUTux3OJ5t8bSFkQQUuKUdoxL6Ntzoyzy
wCoIq+ih1JAj1CFcBIXsbZ3Ro8cxFqrhafVvBOdFkF7mRZvJST3/tKIfb/RQitaK
S7NBghoHVM2T9znNVBzAbN0KtIVMk5wgXkuZCN6Uggr7jIYr4ZoCQTfGgafC9Reh
z9+ev7afHVraSis16uVZIAg/7hranR6SB73ogl4zCu1gF3Mx1IKiUugyZhPqfCOM
GIK/UczM3NBDzB/PBZol1GQ+h5tU2R35zC/1rsoFow5bW5fXYk4bwqmPC9zkwVdv
YgZ7yBHgii+FmWjNKlNmf/WH1B6N/Wc/hfQW/93g23ohYcYrzRWYNwrjBaOyZ9m0
8MsGo/WkVJcqCpY4DJ7CTNMLn383SGzOP3lTLKKZvrnv6V8D2BeTGJhN0+WmJZu6
vRDin31FPZq4vtBKe6v68yKhStxFjOfHf70j94fjoSBRQnVRA5MA6szdpC0QFTDw
kxWRT9lENpXx4i9vEWNZ2p0JWPSNsjLSw17zkxq/VOWGKXdLwqB9uBhaGtLRYi50
DzYVLJaMZU1TtCPt2+Ov4GPUk9o6e6hAbTpK+4Jpxsg5NQTG75olp5ZINdhi7tKj
dpVQ8W28sLbN2cEMy2jQNm4AlM2EvN6Qz1mjfHYCs/SZHwO3HpSENY+O85mBs70y
mojVHm438WMKlFnQZX06W1mQM2TZanU/qSyTeTx0fJASoMdhrdvQXbe7ZfqibkpX
4QGqgHm2MB0gzqSVpckgt2PbXvG3ZRkz2vW8bSmXsSA=
`protect END_PROTECTED
