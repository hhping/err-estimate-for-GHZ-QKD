`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkK9Lp4iMbtTEmwfpPjvmVv5qsNIyrd4CX6IFxFywNIBrioHtT/Ed7ScovNSUus+
iLNXQk78rGCBeBdqdyLmeb38uhL05PEbIFDNtolry0wn9LdwhY1jzmNQqIwOLIUL
JqEAxBXF2hiUTdO03D/6X97LGN3BotOzyNbKl8KJs1YY5XS+OL78HvJYWX/9sQKl
oZmQyiTHhe3GnNuzq/4eXCX1cMe4YYhRmZ6fvwaxy2WDnllCh2XcAMPYjseZvzXe
CPW6wkx4TBFKB+Am6m9HxcqD0K9YLUvMHyZgEbTZo0NNFMvRvUFO8BgsyT082Nlm
dgQi3LDxaSaGUChtj7eMI9uOhcoQd+/7T1aCVmtDEOjROx+JcEYGZb6C3q0Zfxbm
R7+XbMoEB8qN3Xkr9kZ+5nGAzE779aADVymAfOphK5Nn/EEdzNgVZZNBH0VAALJJ
zZHCMuZpVU7mMBaIci36nljLJDHCJAwNMBK/P2aOZ2HYFnB6Oyz+ExbXOagfcuZ1
Z9MxNHtM4CdIA9Xky92E9FV/LVXZiNT2Uxf7EamFqLYqoFfUq2WgsDTc5JgTMcJA
awaU0RkqX3BBoVkg+hlV/FkhbNVYDLkcK9zeorC4iDqYaymx8O5h3NyilLLBwFzL
4QjHP3qk4oxgQrDoLuxg+n9+WQIraDKAl4YPnAMw4IkKm3FpY5uEbERUicE2OCXO
irHCiG6sBeAyHQ8N9MnhdyacmaR18KaFh9vWD+cPNND7l9xowAN4N232jtYHmsZJ
Zi6nGqC3DhUIfyJusJtDue+EdF8ISGkY3nplUA07lFUT9SkykrLjfIvud65s12zO
Q7RqsLAMnzoRNH6CWPayD6eDTy+uo2i4WkWYKoLUjrrw/TJu3T0s7p3vjeka9Z6A
bgLOb8NRo6kUqFNFqMx4cWbsjxmBYRPsQ7zjpbmbhpR8V1XeQhPf/k/tZQ6aJOD5
uM3vkQnjDbnPaib6Rr9ThMIwSqO8p6i1OMY0cpKzsf6CdS1T1azv9kndmmqy+747
cb6VPJBVe3mPYqyZ0hhNaGSLFktm5c/u3kJ401Itjcf+1Hj0cz2hzhzSDzoppnkZ
`protect END_PROTECTED
