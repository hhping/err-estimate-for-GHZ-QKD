`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpvATK+vV82x5BSeXewvABa5+QGJfYvtYdrK9bddyh/mP+WMZleSkyZFgyn80FA3
5m1pE50vxgi06EFrG7SwTM+Bb+moz6WwZ/+loCUaYdUxbBryZCbLfxSCFdtC+oSU
lQwfT1SkPUqae8tUE7Wla0YEX/O8XvCp0F1iOdqxeNofBjrluro5QiTbaoyymlp8
SjSP637naKL2QorUE5mzPC8XixzZn7CzKU9liS2E1ELdoRPuboKFMTPz6B386YGA
GoFc8Zp9wiE80mpfaxO/5Zj+VF+EkQbB+qVjQJnnpvZZEOg4G/HeQNiuTURO5Ilb
ChTYMNdTA6R97/q4MEIIcqKAt9F4JGifJbbaTJlRyVRAlLH8dWZ9vZqVrlAqpN7j
`protect END_PROTECTED
