`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwTowKmJowlucqz8iHNjNn3Eno9JpMjx/LdW62VaTEZxVE+dQIQpF5iKg8c93mv2
cXDyaT38dUN2uDBpvHRL3XVVHMM9IBBqH/2TyEk+Fg2NJIBF19Yr2J4ywc5iBm/1
2+XYbB6YKRn7++PL5smKEtgjrB3lVo7hfDYhWv+593VLXhxPqwkU9FEyfwmEbvUm
m3McqTNqY2cT5i2Tw2wNlUGtu+N66v7KdomRAdOZ98aWKZprgIFGy/ny/aZSea+B
wR50n88uNmmypOfzNwXvTZIdQzF99MXJuAs1qOzWRMO06QOzAUYwweRB/Z8ryO5O
ATnfRIjFQVZOYW1RTh+diHrvpqdUD2Tx5MwXNG/YEw6g/zw6HsNgBl+YGeboJzqT
VpxLS4zojfmPgivyyByBD8bsSpNUOc0MTOn1N8kkswMT7bmRw6PMnO3DxMBZpYpU
PiBlPisMLY6Rl0TZHUf5uuQyTWJ6ZCE0nfTPB6DjxjiHSjMuapXdsKFIW5UCILQQ
U+q9pj1XygTn5p8s9qSpwD4enerzsBJtchY5WSf9wSr/27E12CwsHl4K0GmO7rwx
yp00ez65NZlZl/ebx6NmYnVVNWV1PcUFw2vewFMYzPYZ1eNWhneB+k7qIv3CDmzu
+aSz9t09aFX2yl0YocWGoK1b8ueFNKW5tUmZaF0+96Ikd3Q85w/Yva4xBRrzeXnC
ndE8akHUnQHxx8Kd3aMly1yn/9eGgIZpN3SthNSnOI12ESd81mE/T54VwMPRRzAz
xi+BwQ7v7NFXWpkYzuWAASG+lfYZBVyOeyBtwaPe9lFiUXEz0+DpawP2ytIWLmXi
rwxUzwma4pZs7FcNY9uFDqKsUQS74q7rFYhEmyE1IcBWbiCGIAAm1eQho3f1tjuS
ROoNjhdI7mNw1DxzSaqwinDvK+ofA6JH5oCgrr1ujAge9KOWpXHB7EBGKBIUm1X2
YBMb5uyD6yh34uIW1bNTdEeDXAtO6uUXB6UVDjsVmX4YmVY/aYp20pPtG5EZYHvB
AG03toEZlgIHWINiH17Dn8I+6/JyMp46GfumjcvpnzRhqoYOB51Kqp6kPjB2jBII
v+5rI4WB0w2+RGBAvfrnaA==
`protect END_PROTECTED
