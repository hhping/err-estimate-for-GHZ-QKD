`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hJVXZSPuhseizX+wYPBfFo0sCbVh7NOqgjQpFBZMm6DqPXggZQ8V8lQkuErRYIN
SzXYbhhL3n5bjb0tTM6mGNBf6jg4fLIIhI+Je6vCiZqiBHaYtvHorh5NDlMcl6mU
oPJLO5u8tougu5Xz0WKtJdYx5FgeKQyF/LxRx3eXS7b00am1IYH3R9ks4fzXm/fF
k+Hmc5m71ev8fDoJ2sE1/+xYMBSH95SsurCTs70oGNRjeaZbbefYWbsruFqijx7m
DqbJmm+8tXh6U9Wx/pMWpzrDxnP14VjoihEYBCRpI0g3vK/rJCJJGCblOp3D/tL1
8NJ/LZ0uLgH8/bWgqNSyf9KiVLuLplQFpRTKMWpq9Ke5CP8Nso2WWgNS7a+SpC6W
Repdf9dLe8/QLudAeIZsHE2dgco6QCBcf83NphvoF9+RJaQsAhqte9mmr6HAndS2
lmQjU8b5DquYIxws6kIK/avIsgRRzkmtvrbQsvb3QGXXZczzO604CIGdw0NDSbzi
3pQJJ/rajusfaKFjc9qtNmSDiYB4QmqRkb6lbC/M4VqPjfYHPnNX9+QGlWIGLXgY
u5LfkCNiurcqsRS3j9fcy9GLVc0NlQdvuIQ0XgeVxaJdrZide0zfYLsJCwvzkh7L
txWgRCx+ReKKtkQHDkM58FOn+mVLHKLCgWoJy5D+nFqWZbdJ7/xZSepWZJCscV23
DqAP5ntMM/ybspuOQk2x4BWAkuRxhoWhylJMR42KDYIBcRfF7LMxaBWxPBGxPfK2
djcgQVaoKmGb1aGnrw23K2eDuuSM5aOKDt8Dv6PNN99V84D7gNZTlPEgBv5ikXJA
hHqBuEKBnK4Y6Q99ZYKPuUUekhPseb1MiJfMtBREz5i6nO6H2A2GqHono8HTOHRv
+fGaWd1vd6yyRJDAiuNmCcUAJmXKPZ4ZcRgBeTjt7JYGVBx9WcOwGmKiF+5/tT9G
Bgs2764uDJe3WfRw165gqfhUB7OfWAneZ8fCjtRe/YHRN8j/wiKkX2k4CqYbJZd6
a0KDuS1g3oWu/ZUWXnlfniRSlhvXJtk2Ru6JNQIREpRxYcL+OqPMVj4+YvVBDFgo
bOpUfdcbqUHlHgAlzJACc2nIFjNVlrKY4XNogaprhfw2koPQI8BBsLs+MyMRqr3x
eP8JXdeoulrby+zrB6gVpag6stoBGo/7MZrWcfq2Asa0M6XJ/wzdBFJ1fVsanNEN
QasgM4yU3OF2W8LKlPlXZ84H8oKllADwW8oHrWwhfVqF2dhk2dLPhTXu0e5KqoUz
BD/vRA2zFhKpUJZlCSTimZX0J5JsdX1psCzx39uHvdZddNAzqWqsaDs/7XGYnQ4R
b1IS7CkxWVJFit8712er/25rd0D3KV1pAPubNHpVQ2aPvuI2gMG7vzAUrRcejpl4
jATMWt7g1uPmT8zsM+QTQP6ZxM3WUz8rjGTs7bIJRQRRn0SGIRI1vWt0Q4hXGOxy
V1qcDu9pB3HH9PJ025BQB4S7VKaFZ+9RkT1NnQOM6zCVBq86ALvLN3WaQ7kgO1jJ
w6M4xX8g9NJ/aOgHgDZwOw==
`protect END_PROTECTED
