`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bEHgXaokWZNezJKjeUAyNg0h1iiD0SgMXUeTh01MDqWE2dDZ4NJlXtbIsPWXQ7go
4XoCRHnOQ48iEecD1ImQUSxMBeJ0lZf2Bz6T3ctdgXE4903LfySheC9OMJOsIgiN
CTG1VkTDUWtRxsPOi+FW0nG69+LwqOpWWu5IkI6hI/FYDgO9atEzqfaexHAZu1R3
IUkGKeWP3ECjMbl7WMqW+0hEHuEvLMq09LCWvsZRL8F3VuvIfwWnR6ax0Y07lTF9
92kvDx2b0xdUPJSuEct4Imla/j2DrpOcQDAaAEv9MHGDk1xhT19ElCQs4lrPa7z6
cY+QcFO9Y7iyieSsn6vnyCafe6tRnQhrtYl7chjDPlTwMihY8r+7GIga87sfWq0H
wavu/mII54IOm9sXeVTWedZx1t06zDQlY1eDUBtqARw3yutPldVP0R0YvtDCWHNq
Dk71CO54N9Eq/OXvSQug8DLMTUgarNp2/rNoljb2wdnfS6hm1M95cE7uYMogI2Sf
dqHhv5/Ie737Pj4egUphsOchNv+T7Ts44yK7+pPu0Gi4+jee7y+viAL7DsqImdO0
sf1M457DpcEjpWnIt5oZgJRe3iiEPZ7k8YQuCNNnO3GTazNyDacf4AeLOJebcmCI
5FhWkBHWXkcHR1q//bXeI12WANxxlwr/VGHpX03wmVCf8fm284TUfFzxNbQKvGOJ
f3XKYBdjr0m3qxeebhC3DT3pFeVQyOOUahRZEL4rLDRs3uH6WQ5mJN/hyB1i4OjB
NtZ8aShDhsQcIxj/jq4CsCYC4sunahHZxRlZyGmbzLE8W9MeQvqDVWWL9lXi80Zj
4AYuTOryiZKktiR5ymQJ/XPvKO+0Cn3+U2YS38yDLYQghyiM2jja8brC1VQyXuH8
yPi47la1wyti+rdeLl15txDM/jjpcSDzfRZNuOGl18wwvhYbXl0lRGTNt9o8APKa
uxw8Z0v/IHjBOWCw4UgX1WDfxtlw0jz2m+4pZ4nQLNS8+P4zVH2FfhHQibF0aoLF
6gsaQ8qVVrswXhoZ8Qi8rL//D2jCV/n0RTEBYUyXApECf226pn0q2Y1X7oIE9Jax
Q67FHTITnMMAUh5Ekas7jREclHoQRgdLTSaMkuFsQ46FaLbXEcLa0ihSf9kdDgsL
ZWWPBm99A3TMaODihguck+vfOvf0k8s7DwYLMD9FvGPoakxVa/RtrUAlDd6/lpIy
B2EZ2b4odgUqzmnru0LXP6TZpOYK01AIcTI5T6CQlZ2UFKOyBW2mvDsa0rS6mJGD
B3m4QhhU3NZKd+Buc13u3GPfrbhowqJ+1mXsRDgcHKGi9sHlMWohKusOXnEij7mx
QODTq+dDpVPdpqG66BauurvF2Ipi13X7h8YCFuEi8sTmigjsijUyh/mTuFTHVPYB
G+13foJ09mIdM480qQm3qPzjTR/HQaiUMuyXxxKrkLeRLYjg/vT4RnCjw3uQYBC8
sr3NyLqZzJuHfNS9T4t03c2SKjqgywcgelvPyxb567buN6lIaA8uohEzHWJAz40m
yOqpa8nTII6v/qzqNBXG6GWFv1NFzKI0pej5u4CGUjc1KwAHzISVT65cLJVdfWJg
RalUwe1OyWRVPLoF4h68l5P9rN8ilqLkb3aVAZONUNkJKuJk6bRmbd1LacARWZuW
5ZqQY8PpmDd8PKfVijp6qjdFmU00dj3Q9GwbAW8JF7Sfj1ikJGBIMQDk6JcLo4jb
R01HJVi8mSP/vUzw4fmStXSUU0LqgfuLEU6GpdqkiN7r0ivH/1yi/Mojzp++tkK9
TEiQxrIiP5Ai9Hn9ytuz84eDb1OmcEo28bCCpX8hhobNNuw6FNldgW2nyHiG7x9Q
W2AjwGkPvPXJLUsak1Lb65xWIeNjjNOu+Jos7FaJBp3BB6yg9FWt8XTqb97hfIpn
4n6bEk76Pa+2WC7jEdoiXDxA/JYYSDur2MdKGOffFkWrpm3ypKW7jGt6gXO5fZmY
v5bbHOfB3S9sGXzRfVgdEgHsiwcdchrkhLn94R3knUrEHYp7IQcB+FDRMINMB2Kg
INPwolzAP/BCdh1FZS4CevTiBu3QOqryL/neeDQhKCHmCdbhT9WtpWrQWrU6tZuw
ej+E+9IRclZsxZ6zSorytbTvGEp3yCPLWu6nS2nKskLH21LaNrcpt4h0D9VSUR0W
/mSejuB27xxcr4txkm0jFlCA7GlRZ1rWD6xDj9aeWWIbXsEKddbRhFs9onQgzGUk
fjQWCfWePJjHdK7au7b+YzaKozq6BXfoR8w+ZxO79mxVn0ml3kc0t9Nvi9YOMPit
Tqedfpn5pvQoz/HPq9O+Jpimi7sZbCqp/PkZX1IJS0BAzRmjqbfz9rQ7TCu+775t
pQHl47xHO8I4je28OvXqHOtdfsgMOi3PGkMsLIs0353s5+fmh++IjemBiRV744/j
mDAxvG/D2QjrAti86fnh2hpU2SV7wAnlcsweFXpw3eneK0QoxbI6WBo3bzKeNl72
AhG9M1NTNmYeDMMnjzMWVzTWtzTOTylFwiL6iZJ42x14ZusqV9Isb+egVkh99ccT
b2giP9ljEWM+jdqIqLqPRtBCkny9+Yr1fOf/dbx/GjN/culqNBFxoetVJns8SaOe
gm4labpb8Kl4rYZSq5yrF7PK1xjDqVcjwdzsOoN7FljkOTMveIZdZb5JHHQMB8p7
fs8YAPqslhEqycxV2x+XI51L+W0lW3bliRxLP/Hig52Rcph6pDs5WKMmPZGxV/BK
c11HKbPRszGAKRonWOHFgh55L0iybo0PQTs4t+vq58WQVZhvlZlJs/h74tlCqWQm
OMs41STn06FVB2VOOrF9yVHH7cfwnsgqWrHjId+grsyKtnS18apKwrbdb/QT7p4b
jPEhI3nIWWW8kgb7QLsFwi16yNBPFWF62Ij3NDzowMg30heOYuXUUU1zLrOnxmWP
2dC7LN4kTGZRIpKkKGmH9XahBED6QWZqEWpJ+qCVNQkx6xneV3sfjGdt66jX/ZQ0
rqQFusMBP+XSizXCLHQ7nNQIg8P9unhKs+sT5qE7OHabE1sg/JbKBcuep0Xldmjl
Dlvfu5NpwOEPBB/nvl9xLvGaAHv612Lh+R19g6/+6Lc+2UODUbo9PHn/0P6/VwTc
GzseqSIXJrKFxlhI6vhO08jiDsNS1bFtZZ5GR/AXwiTOm8ZKf4GLRfVv1BwwTabx
o1/OyXw68DhHIpB08V3tjXsjvAJbF07tkhUR/6MkjeMhj09FT0YVV/muWM2Tjjxr
ubI5qcvsVnR7zGox35TdRp1nTLUNyUDlnhJAyEw8IpewQB5YrjPkztUsSfKIwiCq
mAyiJBGgJQtOx9QfsXpNb+42c7GLbFPzJir1L4tj+zwl6zfritojrbq2hceEj1Xb
kYDPBDrMw35HTrSWUyjskh7nZUss3nuieVGnwh8NApxMGza8qtsck4VjQIJqKqXP
QHfY1GgSo6bbDbcvxCyEGwFj7uOu9j85lj3BwIF8iGco0QfWRX7sHLtvpmJLmyvB
gvJklnkoe+VcE+pGp/ETG+6PtF2fObuDtiJIk8ciDp1syGsBTwmLvomvDEBDSAFn
Etj36wW4xufLe6whnYdITabNysuacdojWkw4K6M5CyM7jHVBquyALJCrdoEir+FU
ZwbINpJlQnaMnq6ITqxmqhFbrZ3NcVf1+emWF+B0dyTnLbxCx2TRs3j8juE3+mHg
w18XCxIowb3Cy+uMMS6wEP166I5JOs4Cp2GX654NqnAj5YQoOFYbiQtnd6MlGOIh
Lu17/cDepqcufuUV5gU7WKWlChWw25UNoWLCcRuX+9IZmAI86e3o3Fd24xA8YW/S
u7cZu/wHkiC7pBsI2JaosJgWq8MHvst8AJeznqv8P1tS+wfKJCpFHTLqYiTDsu2U
R/sZLBiGUW+lCN4XdFIesy3XZ/I/ma1N7yXxUFO0GbQ27KIy/H9QkDaWgvWs75FG
0SNc0bMrXIVY+f5tRAyviFrfrRzGogVaEa0UrXgwCZEB7f8V63uIQCnuzYa/zn/K
cA5aoYBWdRlCjrWJ+iOZbemP4yl4qYZNhKlCpq8tfDhf64zX0U5fzXrDn9HIj938
xVSm+05erI2xPy886Ls8xEAYUZPFplmhzev4ZWtJfcX05URCtGOW4mR9g8tqYdgi
e1lr86b4tcTj4yMIqgdBrQz8plgzDDCpIdnox10U2dCpDEFsarsNQ0K1lzQSdEJb
pahGH8rAwHMW9cIpE6hEgfAm2RMEf1vW/lGNhF88ffpQd9K1f0qKNkTJZJDKhmJ9
Iod54GFUVAfLSsftKyuiZ4oSdMNRaYSpK6eCzSxfpSgxhyNcLxaXZmyKfjZncYbK
VJTcZeN8SDp1stuQPUCzupLfPqu12UeslqCwJQGa+3FMcaFs4fBzx5xQ1CDInyS8
vHjVhuqqvL93YFnTjMytSZpag/uQLaH82Rdjp+RDtkjRBt3NqMJOEe1L7FrpYwMt
o++6x4bnfbyIHAUBeWYZkhYAdGwifXnBmaJSGsbP8DXSz+QJNS5D+Bryav/KN8Wu
JEzhC8kno3vjkW0KA8hglWtGbZOp3nwPg+IOESiLKKSMHYDy+Ah3WcBiVtLV25jP
FJZYqRwB7VIOOV+liydh0370pdgDkttygUlQnN6FiPoZxbz3/M3/P00m+lArG13n
27tyvIntQRzuyTR8XwLiUJjL+WrRwFHvv94ZT70bw+Gs6UgA1Wj+BfjGOEkZM5Ye
wuuPClUhZCwPUK66XlWHJo07kZCpWlUSqR78iUQU/Tuj66t5ZB01vSmHwbX8/+05
M7qCtXrty8q+Bo2qF4nG6BzhZfEsGRMCzX4rCIUxrbQQMkcw4+743QO/fwELPROS
nhKcgH7lLfxtFqXaajJyHRrgk1QXAQEA2mlXsbmcvNruxRrnMcPcTpZvzbXmjPt1
iU7bn5Ie0XGutAnfB70eyo/N9PBb+SJ7C/LzUvERR2jQqQ4BLa5XNtE6A46xAKLt
ol8TQU6CD8KXcnMn0mFOHplmS3DeK8y6zgBBS/gLnAvAeO58iKdvyKFsN5pW+y7l
NcgFoGGV37veC1ZW07UCX41f9SXWhwUmlU+ZCTR0W7160obPU2/8UdaWeew1OMS3
L7suvNgO1yE176TnwZgurHOllZtAx6+JPZ/dsxnPxa99y+SuSYJpbMqO/Yg7nnfe
+V7HlMdF+8mI4Yaebw0nVV7opBVO/IuAEFJ3Vws/iZ1Vl2MgLzFWYAOGtnBHWoBz
s8hmzOTs0+RUiotPJF/7RhfbH/xnE7GsBsuco8blyw/bnYXetp5A0DKfs1yM/YAF
BXGm16OXy+gmwX0Z39kiR9IRLKCFzy/gz7OdS1lOiDG2GmqgTrTIzFoLNuJLgET3
d3lh36yCm4YLOrbFj6rtME3OPsESoWCn3PavVkPjXqnIEzTVSvx3Ed+tMFzEJypW
PLWgtFu5+rAuw/xvXvrAvkOdj23AaTUPEDbEOjum1rReKe3PDsJvIQZho0Ixg1+9
kmd/64KdbhaioBk+8RV0Lwm4Fw69zR/8eMiDyY7Pmcacb/CTEUIPAklwtKvZPn3R
MTCl7GtDJXRIG9u0rkrqX1N18ir17czK23uh1OhHKygzSV+0NTfTc6KFESiC7gXc
AwD2Vgl8wHaigjphHHFqb7MoA/bB764jaEc1FYKXDFFFBdpzZuY5reEN7R2udJBO
M1+c/FBXTlQGG6ZEFQDSZdDAxwJvzaqXemXyBO/ZDetfzC8oG9jEdrO1KgpYb3TX
nTT0lTcraQI8yh2XsFRTujjfoCqVhCk/LLWar0vLagsbQ9ozK/zybE9av3nNgAXQ
zXrkCF2CMGqUlojGP5xMbrd5ZKc1fYt4mYtHFAjD+BhhGgal02ewE7h4utyf87Gi
OYwtUnuP6BH1uJOB1JmUY97olNhoU1Wg6HTjdIMRL1CWyk0oNQhzbAh7iqEF6MHp
DfSro028u/XvmQXrU1CZuwsWR5QxYvr30xG96NBhA8JhUmmnrwXcj2GDp/QGyC9m
p/FPkUW8NOQelCYCEnLuLNc900SPLEcsSX4zXninELAXhZbLLxnPLe7GZ/jNVhhP
h8bgKcLNLbgIz/F4ixMvqp0tBy2fK1nX646adcj85Zb1IqpX5mvpkroHIf+503QP
y8z/r5p7zEv6KMZUl+W8CHPFJl9jk//1Hio/fyShXKdv/SiQjBCHNgdftJyHABnM
v4oIwdeVSlBQMrIC8qrKvlEyBvIewMXeLeb9dp1rX/vvSff/Y2JuOeCnIf9m3e+v
5b0EJnaMjNApAqlb9fS1S451jaG/Fj4YO5rt1eEUbkXMj2qjzVi84UjeFL6y4eW4
m4yj087IpucGa8mD/cnfddsphxpUhkmzhQnQcuHtnJ93RZThbQUnOPQWb+glhPic
Al71oVIsWU9ANGiSnWbZK5oEzkjCI2AcrLefxzP/VgQyIHEuZ45+swWK7Bm3IY45
MzoSP1rIVzPqlsEuJnIfaQ004WEn3tJT867qMU/Z3eK4WMRXx688y1p7oqADJaqJ
MLwI/Hh3QBlw6mYAQ/A9le993GKRMCHZdZNkB1ETHboJUYy96zZDuaM27sUbl3w1
2dwA49kOlxbn14ONcE7dTztnkz/wcyKpnwuh6kVYJWiZpBjo2GZkdAiOH6PAgxnm
fiIBJKUhV+YXlksDPf1stiVjRIk8tfCHSqH4ZjkPNVNWMLfbD4aCPb4mrfoKw213
S0O7kBmMBbiwAScu1uruxEq/4O7f7S3GhZwdffA8PK1x6VRowD75YBF5uwvPa08s
m2AFy6ZfzQelW9g8kOYfdexZ/aavRoKRrFaRtdGffeBzctyDTMmLgYHWR03EqLAR
Rxr1HVrfSWKuNWBMWYktigfN0cC/rUZzCGv2P+zH1wCtw0NWASQTfA5rYvYKgAZp
AGk2JfinfilQ7H5m1azlDEqDlV55evt2/kwZmYtdfPbwT40IYTwy3KQ+47ajZ3Aq
p5Kwg2isQxsORLENTZ6tvcS2+Nc9qw13kO0Tmgerm2bpi1z5EulEK8vn0MDfMcI/
US+YjdPFfpTfDPRhikReiXdkzIc8mC9OGm9GLnQdaMbhvzkeb4WrXeuZDjJB7cmv
tHhHLZ8f1SPZMkuTuz22Fp4VD+WY2XnO2s2jnqN4r9bI9HDb9llx6anCKldG3mZE
9E/36/A4QOjHaMGP4eWRuWq5Q7q0OikX+pNICSF+PMuS5hERcza3vGJAOd1Ydxua
Mz23Dkp9MBUf8oK44So4qSdQ8T62M+6UykGmkpp4st2QCwYAozd2kzayesQc0huP
4krhv+SU+ttrTaSlF9mHW/dyRLJhBliHdJt95IFM4SeyR3DZD3OI4kFJjZFnx96W
amTeL89hX+QnAR7PqNsu2Jck98e3IPTV5e1bCdEoWyYQLtelqwiQMFssz9xOmQxh
jVEByEDHKbkKzUT32U+spAX/Nu28RSC3GxUChPzlvAEmj0oIWfXQ4tcNcSXuJvKg
dAeaSCvpip7SQkWANUjqfni8eSlpOH2uoIM9e4uLTjrpDxkBW7KJ24mJJ7Od//pM
svNoZXUawb7uGFjq6gcPcG7yrwEuP8pZmqmkPF8m4lyT5j6UTzI00tE5kGcqfd5s
w2S53nvnlm+rzqeqIF1E09dtGetR3ZwVcsxff4ybr9ovD5xNDv8jV6nRCjMHGIz/
sIhl2QmkcNQ89uYL0vkvJ0DZsxi1/0CYWKBPpNbT8lWV2dcDOfWlxe+ZYkbaP0Wr
WBabD/IJ7hoiyuEBXCYME9uanLxJZHWbJxEfGNKf8rHv5UHGLfHbPeTxiuMbfvKt
KwIzBPWgd9MDYu1TYKXdes/WE3ZqNS0o0bkG6HW2dLK1Wn3L/Xt4yEnWLSdzMK4h
9b5TWGRbGMfZPq5Zfbu9g6mRg+9A0hojhMlDygAn4kidCIbDSoqmAML1MkfT1Ioo
aPQwUw+Kf09To85xPnMdkXYwzsonMuQ/E1RgzeVfasVFQMdJm8EgYtWZTppugJXC
Wmtp5jMNmE5Ln/VmOgmauRPz/bYgp+zBc2qzUfLiKys0RQraFJhwDXvBV2Jfma6M
af8xfwU3TI0QYAO22QA42vdBg3WEuwMBpMwcDb9wEph1bOymk9r2tLwQG9e2A23n
jj4vcv3ppTicEKoBno+yHkhO89Uq37/pEqF0DwYdeBRptmbgGk9IFh2TzaGCORQf
dqUx227GLr9qKxexBYzXGCNFyMY/FXpIshBP9cZ0BAxsO+zmoLH1y7sjeZs3VMPa
56V/O7CzAzac8AbpwG17pO0X+HtcGCCqVRl9pga7xFRwKw1lcB4SZur2L1Z3swKA
jG9NKgWulXt6F8M0SkmwSNOe6bEe8rqFGm71GgOeLWHqQzPA4ZdFoiwB7IG5fiFn
CGML/S7oOpSuOa0N4ksPtj+s+IOrZ0KzV7zofA3Z9sZiehc0z3zv9hLHHc/EGjWO
bVwfTa5EASZ1ezVwUE34gHXt4Kg1hwebLcLatPJBJrqWrwvnxHdIrPv2TRdA06fz
8ozAHCy6+FsUC71uaDdVp5BterRPiXQD73ETiFc9ptaZAeHjdQ4ONXPTUaKvZG5+
TRZ6SDvOaVZxis4ZIaltdrpHfCyKn0NfreiV4MjLan+Gce4MGK2HQY4w1/Bwy+K2
ziywzFwc9Xh4nY3Hpmf/BE9naJdexzexvhH9THsbuGLp6a+R6WGxKHjnzj9PB0W4
WpHTKnmSMWQehoOLOaTsbtI3LLNRL93Prn+lJMtvufBJbGjxKjFLBXrT+BhrZ0Xv
dEMYyTZdx2gCTf888/C5ISBSsGRTsR88t5SgW6/Mc3louU6kegkqC0xEvXFJe4NR
wVTxaP9cvwmd8pZP065RlAGjx+3/dMqGp452+JFyFLb+0mqCxtoj8ZBBy+G2zbuR
81f7pDTqowvuPTAuprEt+A/m5YPxnO/De2XHfwuSsRMKvFrZ9xnqAD7NU8suJ8jE
WAihdCTLqKC6ds98DIAhMPbXU5G9I7PeAAE0PXsnqt8VWl3pfoqkmm/ETnVSQmG+
WodTEB2nf+oUxP7RcK5V+esZdtPC3a0vUpLdTJw34T/hhYPrVLAo2ssTmTFkB8lW
JjaG8XnLxgROLhycO7nOQuimLiK5AnVM8FLRl+8uHa6usLmcTBWw0GJeW0VI3Q9r
FA56WJaVnWwVaXbe7B+bK8V2+MXl5eNU08Ii2c02cTof7XBt3+/lDZI0xaGScNg/
PF019bHJjKtw6AbCGSCADFbNZoysYfInN3VG31M8p4NqDuWALfWElpyxAp9saQ99
jbC+DM4T/bDqyT/ZvtfPvD75EaPPSbDS6O7ULB16Tq68k65UVioPkmv9t/imxz7z
gaPi8vWiAMBsj5ugAPm3/BL1u/29GQwRSgh6rM3V/HGPW8At1W+m16sVEJ0YKsiq
poXeVqh6ceK9J2XWAPQdZ4XGoKjM/KyaQ0ZA12drQXV5VpAU2m6bkncQJMf7iqsY
AHSHfytjledsZP7rXodedL8JNVqouwJ1ga1dGKY/SYHik/1ueo4XHhaqCKE2kxEa
lLks2y7G3LVVGgkMlvLEkYNJ8vhCVbgNVCIHIMqlXZ3EsiKUBXcr0LPz58SSlk/m
jSjgyVbPNWA8tBsfg4pXzSRf07jWk13UXlj9iE7IIt520kJF5Y2rWdmqxfSLQd0A
9kA7zI69YYrrjD7XT//AKTe9DQdS7u5m5bdILIuDhY/qQMJFXKMCgZbAZ3IMe2wV
t6SMUY6hdo+CZe+huucaDiNkzUwB4M95IyJLvC3YsVokVKWQVknWzRbSiSbgAA2K
89kwRJ7RSUzGFr4dEI23Y8Vt4aS6ITztIcLR3IUUwMut7JP/kuKSqVq22frVpa7h
9DPDVgnBffRTPUJhX6Mv55jkj5ubfz8q0WQWq+NJtz4Zb3zBIzq54pCPKmDFyV38
RstHVzDk+SL3j+KXEWkra3i+Unh709Hi0/yP7DE9INjkXBlpoZybfHWhdZcN249h
rOMwuFwQ8YNfMKdb9t6/6vH1EKD7ar6k8PklaobuL+rTLsaDNzNcX+vFTubPZwVk
J0AUz0LnGIxhAksUi1RjZf9wDycRVSKFsJChiRkxKq4CgJdXDzakGFgTVKkQY/TL
1lBwaBvVVEEsFr8vceNh3xsMsBFTPdZcyXTe8q2AA10UbQwSw0W2dF3X8dy9Txcq
yDhM3+l4FI/rQhf10nDD6/R7lMQGXpUYjEvlG2kOWNddjDF3+pDj7FKBRffPHwqE
l1SoHjCeWxnruhkYFd7mN9nfuXEZpwqodEEC2+yUCvwqLZNC1apvgcLzLaMIDEA1
UdIxITsshoKKzadPSwo3XGm4CHY9nlil1g+TZgRZEF+n5caiMspyiMc0lN65aQju
o2g0yQ5zJxPkr8XmPcWfM8nrEwBnqjlR71iRE6jTAzrjgM2NPZC6T8HFWh6ortnv
swbTAsFiKogtzgsXiAQbdrQPhYQczeefx+BKjS0saiWoNlmpNX5lr0J6xUychH2D
m5XodmUwUuminMJ74VUHXTJHilHoBArCIoe/zSbZst7ppCfX/WIXKlciwMpS7QLC
NW7z194SqxgpJIwMX93+gNubd9tg7DjpAxgkd9vEN9pI4QwtQsi+ELjxrpLx0pCx
DvdfvePpycsZGThhAYapVXfjSEeZiYOiN9wIBYQl5GvmwSBWNYREz/Q3YoWRAHUo
pm4MGC4UqYT/jYBeqdCrKJFiLYAmh2olH+9qFJFRbzX483Fsy2DcikHOcwppLedp
N6YrmMdmf100Jga10OcQIhKteVaXKY9YhUjHbRX3DFTqWaXkqdz1N+zELd0cz5RL
cXgn9fl5xRG+NIuieftTJSx3wvkzoBzzXm9qRvtXqbszbbp7HaDtsITSsJ9i/zm8
R3kDbSoZqXWna92EYsWtepeMfOVdb2XZIhIRDh2oXpf30IJTkKCBTbrMGCF9gUwW
aP6VqBg2aaSUheeOfmexuqHw+Ac+lCq43dD01j8278aBaykl7+qX4ZngJAjkDqt/
V0dBUjVJCrGSrM0g6FI3Zi1LO2Nd8KrStcvCXfirc7ilU0H6cIpszoa/+bk+hoFF
z2oYuOZU4AW5Kr+Zz6Tlp3mdDJL32cjaqpuGynA1U8ToXnL3l1wDL1ioVUn/kdKo
qYjQ0E1IHTjmp/CX5DxYl9MOziM3nwskKuQJo4mNshVSvrv6lQQu+wDAJgG4gnrH
1AkJ/ThI/umd4g+mMSaaoZ8Gy0WyENsmbip2J9mjkD1uYFugd/2rp2ifg2qTQFQ8
68+fJrhliKI/jJ8HozKDiuEK2U28ASLxoSZVBc1g/cbSffJukm+eQjQjkH1OOQ5+
g+HbkSmGaCC65vmvch3GnCg3PnHgHLA8WHKKJNuAXXFp9FTCqcdzryno7PPpC2/G
SLSm8oqKT9e8OumoAdH9yro6+HIb+iHgsOeM2k/KOGfHxPkMzmRaJFZJRn6wxUGs
K7DOH+KT2s2xu/HsbZREc+W5A5VbYtODkZNrbzAM4dUNSiZ8hZLWuCguPLxCEqcG
9QLfJSUaZ53Vhv2jNvYpWcLkexBjnczcru+jwGL298w8HCSMKlH21Q+pqqXbstDj
FKfIn+TOkYUeUdSXn7AjHw8ELMuBTlIckEEXosojBaF3Oc1HAL9TeCMkrZBWE9oA
l+rnSzSSNOu8vhy7XDDea0iNfgY1uHPZVQtJ8DYZ7DiXWqPRS6QwlJYX+EvBgC4v
2ITMLhVhir75K9NaDdQ/OE1/kCcbwWZtFjr5NNq90LBQcU67Vo3I7h42UD251mU5
IWA5xeiJMsDtPbU8qrjvjrGXA1vHkB04F9xOc5zfwibiqBESNhXbWRaF8Z2XEzTF
rcjzpPlAir4P5vmjTurR9Oq7HGS2xvafoK+j89MWZ2bAucT7oeHSePOWJesDx0f0
8c4AycHm9agVJMmo8zS20kknn2UxIbltsP3fjaWxb7laSWfzgiO3Pcu8j71fz7yn
gVTL2eudFqPKFWQcSTiWunMl1KqCE1Ve6UtxmYqKUKTxDlh7gt9j3pQWFR3/N66I
bnlnkzhqO3s7lHmWqwo66FtODCgaIdkl3xKKVvdyN64F6G8CkgqpJH6E2zE0wxM5
fKCfbxGpb0lVCNtEW780uqOYr6dwkwLJlD66WMGzIfcXTxXiea9RjBvLm2Us3AF2
/T7NvP23RlbhGueXN3mia53jpziZBc+3MbG2Cu2TSuFNIdaDSlsWAjq+jQJtCV5p
qbX0C7frbwtpqu+kF/nun5+OIi1nm/fw1xoqPjmZWL/BKpKZk3gYsynMgLpOnvPn
K6z3QjGVYwoQqTau8VL83dEIxa4zHO6lm1mlDVV+V33BycE9eAS5YDDhHWPi6KZ2
WfWB6ngSaKf+KqnhELJgfxLFJg0rEcGubXefu0ztHFBiN9phduTuBVLLGVHUkt4F
UeeMXpvsVSNbvoDuUKvmuQK6utqmkKtY/4preUCTAoEAPljuFEcnb9IHxw8UbIR1
mu7q7VqWWsB6cqPTR3X1AYgyL5N7frWW5CJbJxHoXfqnogALWHutNlSlpS2Np0QX
VBfxMABjapXnfUw5eUUPL/TwfdERb9WTHW91Ergr9+KKsnkH89Va1cITPUw4OyLM
36Oolj63BiPxyT8Y09Hw/cbD1H9TcY2AM36FWZVx4cdTNFhz16vn+X3/lnPP/PM+
5ggB0g+L3N2d0WZcxCA3gOuHjcus1nQ/5Z+IE36eUxHvr6xlnWBynrhzahHNEstH
nsiqSrGYmjq36/9e9uV4d9jvLQHqceAhZtvlFpfoWqovR2b+PpBbpEY5qeUUE6kX
rRYlb8PJMlkkmavH+Ww4gVErAQflNg1ToPvouNPR/85VsvC6tTfhlN6Tv84+Yrkf
vaXs68DVQnke/bZyey1B7xEpoCgtTQm4vt9DQo1lrZzBYeffQEKSV3b+/tBl6XOo
njAu1TVg/x+KSELkw4wmyymImNPikUfCFUNqotqV/jqCBPT/Vx6TeJgq807i/djT
hQChjcDPuL2I4jLOuhzuawuZN32hGAAtgOznnKGVUr2h6GRqJZ97owCL2TI2/QTS
7ecxZyVCWdegLgk84pQ7Uu8D4TuqIrdgp0eJzv+9OEsty3X4dQaKeKuJ9MF7E5ln
jgkC4W6Gj/2ZxMfupeP4M7y0P7F7BWvGEOe08mo67jdXUlbPO4nZYSrsxImHSlSY
djLzXVW+TFThnLjOnz8oujtcJGLbobZ6A3f5e9wCNHFo+6X8HVj1m+zh3Gfewz73
mQeTTN09fuUT05Wbasu9ObztKbqhGMK4TJColzSqosj2zJUj2ml51niXsX/xGViz
BZR/4BhjnskFDp5CfOH1d05WItJJ3mkJlT9lrQqxjKhET9oxJCTF1NjDMWZSD2cp
dbbTlTeC4LXi4AC0ZX/dAUdWcV3I/uQEm+jHXyItkNj+7++ZTiQ9wffeq9bdGNnH
DUKmvjeyv5G2i3Ho2mLhxX7YKgaXDp/pucIt1kuK/ndASH2oU/MZ39KgPjlf0KRk
YnRwOup97zSUFcn/FkRhohjJOFZtKWMQJ73paLj/hc35NF9WwNtmSt/Ro2G1jxO0
JvQnvWq6sW4PD66TehLwPCez3/QIW78F7a5IpTIlvyGfd+oaUYEpmk+t0VRQLnkx
8rZ1wJarZ9DE8BDye1FPUmx0FOeSnZXElPGXK/Wb39MkDDFgLgAH+m2qDaqNQwuP
`protect END_PROTECTED
