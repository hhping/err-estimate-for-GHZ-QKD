`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTV/Ycpe4AO7Hamsfh92lYX3dd4i6aNjC3Hffaco675fhWkLR39wjAUAOc+yezT7
CaciwwzH5iguGSaYJjhgMUB4QDjRGndhnob89hMquLvn4uOq5ZcU3hRp20B9Jkfx
Lr85Mx0jc0nuTk2ABHssZffHq/eTsd3voMMuahsHBNPRO1dk/h8LygdEdfb1uMS3
oLLJRPzPt+xcZN7zIxUkrOEmdXf2H/5iVpwyaUVaP76pcSYykgw+o28h4bDjC1b5
RhIATHTcHCnxfFBtAdw4Pa1HHtwDlLLKFbqdKfw/MA6tp6eNVXvqpnmRLWBlCed/
WOGFsKwRpB/ED0Il8dW3IMqX9TaLaVJ0I69lIdJLaM2NimpZFmjf3h+0bKOyD3R8
dxbaWIhQ97TPLDkTXzcsu2p4JnNkNLznEpk7QVBp0pGeWdXm1rl0cmAJ2gNSGYjE
PtMuPULii0qR0BfglhanBDrUgkmdFbj87ftsXEXeAC0MDcB48yiBJMcpzvOHHe99
jIZzOsKlEFvsdfHgGjmIKZ6JOfj/Tn9fbm+MHu8OIOa7FIp8WrFimTwoKUPYAmab
GIRy8hMq8Ccm8uRU+uTjgAe0KCoObKV8mVcRWjWHUyZYaya8iqMRV/r37gatbcak
D+neBJ1Q5wONCfxr2YV1hU+3Bpkog53WWbiAVUKLB7ZOB5W22onSc90YWhbAQ0t7
iyjq2bkt0ocnKxOfVIlESc2fllv9R6H70Mr/EqDCbC/yz3DpMATaXgRsXF+sqFj8
6uhkkYrvrypIUBmwVca7iQAY/3ERMu2+ten4QWoSSw5rw/0OfCcaSEeqZv0oStTb
gO49TxldggHm81hngGYuyAG3vUyihAdqalDimfo10pvYcfwxRz+rgt0KNME73dHn
v+O1ZmN8aAiSbfME7XNc3FvsRT0Lf+XHvSFIpWRZIK8eVezOJ4hpe4rrjn+OnJXQ
apn0dL7+iDYlNqOzHrjvS1U4cXXySMiLxKmi5AW7MK9nBc0GmDnlh3qNwn2/GPrW
C3fXD8QLWPxX3YRb9fFyqEa0IJY3Ci1UVPbscLVraPXScpZPOLdHYy6HsEzghAUR
82WvwGRr8WZVGr79jvfWmb7GLxQpzg75Pwm4+pctMaTgeYKOu8GG9KRcaqX8Df9d
`protect END_PROTECTED
