`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdns9o/eIDFC/oQoj7LfhUOmtPdLrH7gpF0dRgerJGKp0JPwzlQMVfrenKjBUbGj
xaFVvyZJL7i7JpLflZY+0tGlpCqx8WXKn7MJYtnOvthK4FKEc8rZnm6B72p+VwKJ
we4G/gd7wi2ujrlYazP/+9m41QQsjMO9mBURm2CTFtxg8f/QjeCAXTRm+x8wW0IH
Wvi8PacERVDqrnFm4ZipDPjKqixOzC21kbg5iZ9v6x/lhBYZS9c0KCDAKqqSKynX
3dqNex+OGxopOAhhbvh+ks3UCVcbHY50B8TsaA0Hntk88CbAynzJSx3eVcl5VIQL
kLGxvK2wCw0idDgNBG1Eb9MNUYL5nnya6El6i5MuBJE/U416VISv30lflMvhB/ey
oLStD66xnqnY+Lup3YjrVazQRn3p+R7PBEGTvO00Eo/qVBFpp9gPIBij70RLuT3U
GqX/kwv1kEiJ14ryCPG5dSgj5R7I/waEclf/Ez615MsfW9n9WwoDJ4B/uzKk5VuO
QBDV5+aJxuwk9C8Wg06LGL2Lh4t1I+eHoDq7/l18Xp25zibcfWSKdxc/2XU3cKiL
VjXpJROCkulRRKBGuKQ0R6Ycc+zYqrbymdVPuYQgKuTRZKUgKqRdE/WWwCW5IBan
tpqnrtdQAsaQg7WshmvLIJYxOBLEoupLHhJpqFiEGdbFhp0QzsvMIUWIn56tXN81
7HQjMOromSeHNj49qzLAG4Sn4OnEp9iNQ9+h71msl0kNC9kRcQrG1RmsrpyF2v3j
`protect END_PROTECTED
