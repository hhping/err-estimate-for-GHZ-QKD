`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICmNEU2JYqsIuaqKeIWoCK0ZEs0By9nMwf+aAvSwW/s/bnHoESIMzaxm/GqmPIFX
zoQYRABqlPp2IkoBH3esHrD07JQZAsY34EfpbcoRpHSOQSFn97Uiwm99KXrGlVUq
5s3YKKhPVaNKgFQ/81LyEmgzb9T2eseMKQCpdSvX+5aB/AiroRDyto1zIatEoamG
wcb6OPUPs+Qh/lsCdm/w05soWyFciVZn0bFBYLauyhUAiMO1RH7JFrjH1GaNNJcM
Kt81Y6UIyzcCvQlq1+sdzT3I+XxbA1RJNy7BIJqjtZ+QsK9m5pONBZQUF6JFo72P
lMFIjHc0FLYK1/b1heDSMYEcKjgV5jCk1zqXzyoVaTlIa4HMRIBqTuK5gveGOMmz
MBZ9IUmgYNCSz/FBGsIS2itCi1o2bkhQ2z0A7O1L0Z/iYVtO70YlZpPQeYpSKmtZ
LODZZrWiQAUTozj4cmpi9CO83++mV4y4x2ZlfHhtU9W87trQv6I5GvT5pcWH4bmv
VAqRRtxT6Z8yeDNaLTH1d3myB21i2U7dHu7fdIchoVrmqIIZBQsMVOg22l8tF09t
d8nexMsXnwBtKpMMK0PyowtplUQ0fNvuSs4EWLSF2EuqUfXE0GegVuAPOT2AWn5u
l2QoNQgi/v+LeOYhIU/ZjSaRc/CeCHvzEP80fvUumKW8TDsPFJAumobR0hzEJWY/
ydZhUKFGLf4Jh3bcbqM8bZJcFidB7cNTQ80e23zHvW7+orDaTbRXyRYUbK4uu5zg
APW051njh5/g5qXrx4r1GeLDWQNvxRZLTTkjiQmlePXYypqd86r6peHo8B+s29IL
rxmhi4KTds2o9icsECdceMmpirNtt06bTiH6ksgF+ZIjtWS/qAdxJ4qy5VV52ZSZ
OqSsb7KMUPXtmzFXxscJ+nvZLfmgLJ19p2YY/IOUO7QToDJIvGyWFRobOKmyNEay
`protect END_PROTECTED
