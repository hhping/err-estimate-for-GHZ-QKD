`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4GooCqxMDCK7fquPN6oBqIEq4Tf1xoYYZjlLzHSC9fNhIenzw6WH97TisICUS9Z
orxKYQLbU2vjUJNkCk9JVHfLo4Cm8chl03DBCslp1blZqIL25Wy76V5EYbR04VXD
hAXszqXsOYGFf0V9bVMai/wEXd9cfM+7SEHFgKcTgf22A3mF9xoiIfHVeKxwIsr7
j0DW+UJa+gOgPX9k0wFoQDr0cQ4fkhQiW9BY9U+wFI3QS/8OOHhnxHE7EUgksENz
lD9IltQgD3JK5kami1oToboJoaOj/8dCAR4POcJqIevt5g3q8O3qADCOkMZb1MJn
BTV6hmF30Esux91cZwXh04ysY4GSuf+zcalWL4OQLFqBdolQuzW+zAKez5OA6hZf
8wrGg6hAB47Yimd52INDbPj4wwPkr7apNnW5X/MfC882RUvbKv8drvW6XfYnzFKj
mpSPBlx/vtMmXH+VXVX7+A==
`protect END_PROTECTED
