`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VlqsxW1lw9U3OLvaEdRyz2InpY79nSVMlBTX3/LvMy0du4Q9Z1O414tHt8vjLlvy
BEPK/hxNo9mvZo1z2fgHmp6x1CJAJeFac9s8Kc3awF8AVrXEdOtFHg1RfP9vXRdB
69iV/9vHTRXzmm5VYRG+k67hk5WP396OzR/nLofeuEJDYLI4G0khJSO30Il2CARM
n6FT6jTlTIdqsSrNl95JKRR2+2xafEydCkSLxKhQPkakXQxzAlPkZ+BXgqSc6/Xf
d1BbEJGhXUD4QpiU/TcpsAehJiyr4TEHaxTswyAEbFYIj8xs7Z8lWCCH1G4odR40
URrj+nDwzoJMXNdkpvaWoazZbLg1UmwJpNMd6IDkKnk5EWznI4fziaWiZ2QY0cIr
4QfHpESAHPY8cJV1+fF850T5DatqBwt6yLWcvium73kccIYY2KSB4PNMwGnhxAXT
iTkgKOA8dvgSrIAldJJ2vUi8VtGQremA8HjdOLRKg7SoZH31VM3v2gbICpAKe87t
3P04i4bm0WHZPSRQN1VxaCS/sWK9OVFxr9XL8pRHYgEfzEvg/5BN/di4W35TsVd5
fRhD3PfH6HSRy7th2vC6nf3TlNjsI43+ceQnbrbgHdCdVmivnt6NDbMn0+bKPyY9
AdNFYYfrCB+S1ergzeJLlA2TxmPLdkT97HQVO0oCQhtQZe48bsKegotlr++4VT/A
NuxcCrwmdfR5LJDKK0aZk94NFo5AnU3arxSD3B4AQOTxaNSqKi19Ss9gqg6+Nlf8
bUxdqeUQg4pJGbW3VayDHP8AQDoIGLtejW2g1WagxlHirKpQu5D/Wd2bJUCOj+tm
E+5Kt99o3mADzG80qKYiM4zBuX+ULqIUseqPovr/KheSxzMoevO0lMUEAi9LKcE1
tljYsVJrLWIlzpClmoQGN9MDzLR4kG7Yp1oz/mXs8DZ5/QbIaNGE9FQwwW7buvWL
BpHAYAHpnJ184n20B+bU98Ts2mCMSe9ozGjxJ9cUesbLyZfuoWcJ6MwNHa03RDtB
1rclFfjB6ljeMmgjxOeIs8c8+CnmRiOdeBUGaIgJZCdrYLx5nWBCWdTsPw62talq
KseDZWLLMdmFp9a9evxQ9sF/ao8WJiLbcU6Et+4tU86uNmSQ8pzNZujjwKDlF/fU
0zZ1mb0K9VwKs9Aug6tc1WZTx7/63kT07+tfwOZhV2biSioctnRyxg/je7I3fEn4
s6CucNkljnscNWVNLDDwSxFqwaMzn74UQiE2TzkePrvBSTmLe/9oLpJ1UlrN2HHG
o0lXojwpGxUAallLtpbkW6i7RJN8UpM7MpL8rv3paqO3V/hz1mJM4xh5mrKY5Ws/
/o13tV7FnTFtuBsUcVURqKP/MUjAE/8HIkZDX3y8AtpkLXdCIqZ2xioiOvhR2edq
UYuXp1Kcrx5tJZy+PuDs7qe/pHLsMrMjDoNSwXApHgTIx+zv/xbK4KJVFsyVK7lV
oOKxDkl/Bj8aL7a6pV72jJBVQFsMnQ7+sl4VrwxIC0TsmUMhKbc2t6/+dTCL2PK1
BAMIei8iumkHQQsMVYuHVWBq1v/MbITwoGWxdKz1mz4f8DAEIN/qW/Nh3mE+ujyd
JpWFjKjSdjVHY2TLwMRKg+g2rBL8laStP8md+UHrvOEu9jsw92Y4EBho3kNKVdQw
7XUCt2KbQTOeSN99LgVT5k7u+6EPihNUXS5P0REP1HIq5YhiqPOAX0sxZ+V5EUY4
YryXrnVJyDIpZdAQNLyLhjLyUa68q/RYJA9UA3jJRN7ZVSiPJ3qev5ftlr78SsM5
/+5sk27q76/osqRnTvoQjMMppUujdVIvapM46juu9NGI/a7jGJcMEnsy04AMHFks
3Duetvq5ZtACJqujmmRiPXIuNEmlUgkszhVUyZV0MmqsiVykHz2RiFRWTWCZCPlE
vchtOKO8wZtY1ATyEM1dFd3CsS5Xsxb4CfvYVT/0tEqMCuaEV0jJJ1tYAEmMWHlO
iumRg4qrZ2G7NfAhnLlBOSTYJx77/a/Tkf3xqjUN3lCIlJ6FUn7I4LFXGBZyXtWM
eogN7GoRVQArL2cbOgNJh+3hqo4tzoBJM6E5RXbXMeHA1HbwC65viJ/wb36BIeDy
LG/bZKi6UDsJkCzt39CPS7bPMgjFjqSh/0/Hjh1DXU6QEvDnjtcEo1hYqEr8AbIA
VFPPm2bXfy8vkl+z40BIA6HRFevE5m1NtiFYml+l2up9qap4vbx9kFA6Tt5SszdT
EG8i4b3697UE7Edr5MMLttLDQaUrVZPoeGcIkr6rwsaY0kOLGQpUmu/BxIp8etjJ
20+xCMUHGwzCtVhe0q1P73ARUlO4w3+/kwmJWVT3PI54lpB/AynGB9dpf2ZqgvR0
c1sSKnxd/zhvyauOO/ez4tWuoFu4WYgMy+Yp3/0YCQGZ7jubk0YrJbvdWslVy3zp
T8ckvJd5WFWcjyz4SjT0jW3lCf55TP0uL/232xTP/dniUOartpoDHdWCLAzgWSXf
fTT1kXM46odWMSfsgeWMDBBX3jau8Myg/+6LJB5Q9d0bIWCrPMWC1iyempW2MIcf
S1fwQnML507XWLMiXRn5ORYSqN4NPmCA2sgRlt5CPZ8wqHKlSjeAPAVLec/WKjiE
aIFL2QkJ3ttfO6guKzJRJ/Esk5es9rFtadXUau7fH0tcHt9ymj1WJtYIC6o6CZaz
jhpT3pR327cfom9PXlIRP46jCUDYfJERH3N5GLnBXbS1k52lz8F0RSppHcK7hizo
6g9u5XSpOY5TOvqyK63PnG7bxa0cvthR9rMpZqzsgQwgCm6kdKoyq7uvT9eAlLFR
g3mBuOjOklnIuggV7kuA7jfSnIDPGSHFPEwd/pWSDk18rpSzKjAhDbv5LciDDHRg
fGkvWWLxp0ryRPp4B5WKQx4bveKGHirR+uUcC9g5ob4TZkggj2Dl51wTi8wwPRIG
kwfE0D/QDIZVSbdjUddax2xnQDAtok/QtwGtuaQW1QVv8eYNJjG5oDKuNFBMvoGG
H9C1HejL3M2wRHPtLk1m2SJZ+BSdCIGv8hv2TsI3WeDpY35HnNAnzwpBeNXL5U3n
8eYrGZmy2WLGD11WppHz4g==
`protect END_PROTECTED
