`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcr5OAtNxHRfJvQLWchqiirZ6QioPxJIYgj41gCCsvsj7gBcKMBpr/YWamONS/yN
C2BjROjaLZQUnvZbsEklAPWe5X1yk8G8NlVggQiSdMu+EP4wj+Fial/OrqVNxvu3
V7sSiopH4erx5eh17Zmrtq61BXdZZK3TjArV7WmLJLovd8LferAEX5AENdqHDzuj
0KqYZLo8v8yT5tySRE12rWIiTycpNQjAXKTS+YReWBazY/Nf7uc++MC2PWE4/ibW
AzxmzOHyMOkLtcPTilHWLOEvRcptVyIvBmBXwmSg7HQxGAd93a93qm1PNFF/HxQj
ZPscUubLjw3kjQcI0TDeVHTtq8XTIGDtJmagEVlB8i3nHdUcDYY22LX1dAbMjRtI
jPYac4QIW/tWwOPxGHnL1EqKvgC+f+sMNG0/aDWSRpGOcxZjJlYwDsB6UmvfJ/7i
9R90MNjfr/5XBBdad7ER5D1a4ygQQ2eE/FiFErY/N5I63gE4MrLAgWwBUeGfe2JM
`protect END_PROTECTED
