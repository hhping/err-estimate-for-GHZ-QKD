`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cr++yewHCsRRKeO48Go7YcSw5QWPWac5w0XZamdTUDaTwBr962LKRkRRpFG0bSQQ
9jqXQDYdnSx1mnEhRTGkyHmjgy5GZqGqQ8qaplMives1v9TpQAfk8zF712JDCSaM
xWdzFIoqvZrw/eUUCEF35iP5WQak1WK34+dfSZ3GnktzgiImhayrOd0V5ogsHdBX
F2Tvd4ffblRCoMJUuTGKXJO/3yYReYkV9KgandpbKq3tkMT3yC5scP98mvx+qH9J
4fL4qC9vn0igxlcYBJKtBtvsyBJX0AyEC8D/RKx39GSo3lfUBiG9o4MDTU95heeH
Dsx8Jb27m6J7MBK/1y0dsIRPzcHCUUUuErdGRWUm0YsiGs//N2HOJVW/tfStSkRH
AqrCOokxg0HOcPc7luqd/aOqhL1p0OCWtdGETn3n+0QyxWeUdbQMkkjq87POIua9
I6nh55XMris56l892lzjxMkOoghwB4qgRx4tLnAECD6pB6lh1EPZHFQokuxmLZyv
mxx/qdf2DyT/AibIpk+MdjF8jQk5DRSoFUfQe5FwPpruriXTIPwiEXSFirbHxx/a
almQBUBWPDWkOrA6P7X2P2oByGDl1BjVLcIJQDg7DDqTrEVS48PBEivVVl8/GeH+
0p5p/xMEbiKO0nkIrsFkf5rTIXvF+eBW/bUwCDWpXtv7gS79allRk1iHPS3957dA
RWOw1FN3uV6u8nhuGNj6ECvd70ayk5kzpBeD+WKq8DXJK3OVjeISqTRlym5j0gWv
lCjRTLLfof+Chsb66hKVZqydAxWahkbT32d/7KCXyxeSIUj6VWf6K4HnOFDr4UmW
YvSfO0VMIcdNwPlgx1kiie7fMa5HLQxHUmwfhUBrOY58Kj6JwOx4eEDBN0yVoy9U
`protect END_PROTECTED
