`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNk9E8RJqJBh5UpOePGgpk46SipBLYE1ykp4Wz95l6imHIeiC4CKbSgfHwS7K4Gg
2E9Uqtw5wr/MTQeLWNvco2fFN3KzqLCcRqQhEMZCDIkQhjA1sKdj8fBMXbgn8AoS
po+Fe/+1+QX90+SxyH2oyOTVyS+TeiiBqZGV99ocdo1c+yg/JgbGyi5wAdZutfCK
XkDLblQz3XH5x8UtI68tE9PYz/PkF9cpjoTOEbuThEbmq/uEvl0sdgvHSO9j5dRA
WWN12lM8uK0EaUNAU4ZxExq6npnAwtaIu1gjneMCXzwi5yY2lVfDe4yDDTa0CZDr
dg34KGyVV74T1PyEv3bPDSnYpTlumrEpOc3OYAEoAKZ+lriqUgp20I8Qg3csjbcT
78XS8ZriECgTlHJoDlijXPWuliTSMu74aCSGCE6KkC9pe53j13WTU9FPK0ZlQYm3
EL+8t2Z5PHGtbZ/C8HYl96xK13FipJvQheZc2RBFmwhslT4a5JjOXSmD55WiZU0I
GHfvgPuApiN+vHI5yb9zKk1FKBA+51WecyaBBUOwJTuryKi/qH1uTTrBq6lWvzMw
d+1idwDqOy6b+q3QKokVhrUyZ2QyxFEu8W530fafTfXM+20nYvZj93WGEUaLdHkr
6j0Eo/jkOWRkQc6ro6190hUAXPWpHQ0EleqfIqRKt6ZydI1kDQWizzoVgubeZ7x4
TaNeEseLHFrzPLq7+AqCskVbmO19Kn3zHC1rvCMvG9l1mgZa85wGh5QB2xcfK2Eo
5aQL6vqTcynYnlj+Ja6ZcYNaJJ4RluT4hJZ8rrpZ50B5G7zEi9jkNhiKnB6btaZS
oD5pUYww2SRLTlfkxaNbJg6X6sfRo1MvbAMaMjF3v2v0W1uWSCU9J5w8iumPXUND
3x9V+yiWajWWdc5YXseVdXjWWKeKLXg/+EArvJIjUY0t5KdZgGqEOkZJ7bLFBRrD
SU4aA+61/CHT115AWuia3jhb/+Y/7Yk7EY/xEYr908aPyJKACRmfT3lPLWL5a5lo
6t5NdePagGYz2Ns2h316Wb+fv2UO8EMqVuCKQhfPkH/w3YYfHrSwNkxUlNALmZTP
DLQIyIPf/Seq+6l8ow+WCrCLE1zwkhLeoWPDHlb/P3Q=
`protect END_PROTECTED
