`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/O2KnJRr/nmxf/EoA9z+K/mpCLBvNEC7VBPTGkJv5Tk19VWaBJSU0NWXOAJ7gFv
8b83XDQu7kKsA+KixNdD0NOZauXQSGfiOCgGPY4D394Wzv7mYaITJ23H7UvNZZTt
Wo7auM8U7rVeKnNZOCe2O14vVmHjXpDKESLn8x7GVyZH5YyU4czuzoIJpQGIT/B4
e4QC7sC6QI4oXJ2++5WTsgRTIsL5j1uqWDaiDXiO1jpyoMiPzE7GxW8W8ouHEG97
+AD/83Vopcx3RlX4oX1S5vlz1HW5K+X1JJcuCbkHEi7bbt2TG3yqmHUIavmDP3LN
mNxCuYd98xCYdOTRgs95NMx4xcJT7XU5RDWWysmuhBinmcF1nRyAX5Ix1qkNPpQM
q+j+Q6cMhxfILVQHFe7wjDWEZFJsuRkOGYsQ01au3EfPSwh5wcuO8UkqULmPEiIl
QwAR0IEUYJZA5uprtJyKN2AecL2RjaufW5PTFqOfdg2IjUzWqYYaGiL5ICkLaPoI
YtQfGl5qQvWSCqiNwsQ1lFyKAKs2dXAVQlBAu31qfEMU4PlUQqoPivx1kgWnDikW
QMrQpObhOnzQ3Bejz4Wdk68iPAlZQ5j0SLgYnrFhBfFFWuiQiSbgtY+aNbOHStN5
ksBEkHQ33lHIyFCutqiNJE4LfQ8sKRTx3ZyYsjjtz1XY6VtCE+1ALs6Vv1SWMk8x
2F3n7vkQxjc5Z3ZQIVD1Oi0mrIj/rtDmlIFkztFDlCVMjuXvAevwXsQgzwuEfgHq
XI81O4xfRfrGvMJhWdzDGMaWPXt+7MwePv/cfbWW87Ixp00Ui9Q3UoIwJObsjO/+
NU26cjQfuP5UcxYNZ8wA8glsSEny9Jqiq54G8SJ3dH2i2buuunC/O6VhDi33wApH
QXv9uEYvdFswHD7krBotFtoyBHUSAw9Spvk6Fltv3d1StFKk/pze2YoBJAMfJQu+
9IMy9fFuQdEmGHm4cPoSzeOBkWwhvFMoL/3e45LBdDtXm1yW0tl+8SO69TrOM8ZY
Q5pJ58o6zXhUobpC5w21xM5YGP+qcl8DTGGWA4mpUkxpOghvfwhYd1C5FYdDFAP3
oEooLsuKxacXdjHUWJl2o9Pj7ERmltyww+sBuKq/AjC39FjN/p3KCw3CMAwpX+BF
wc+qB0H5bSBASDTeRkY15hmefSDedmu8CZtUQRu/6ivtR2phLHFhMQCktbfbjb5O
zs4YSipD1kSx5tb0klgJEMQLF6SFnlLFBRwDkWKbTFT9ugbnULwezd7190T3cnLG
x+pvB5TGAZ3cL/hPa8hwCM5CQnJdi+1GakO2ZFCDXyeoTix9yQWJctHZWi+h7un3
YA5nmOaAAaNdXsAljnZr9e/jaXSkaGH1ILCxXos+JULbSt43JDhzswVbl7uEUr1i
6pjV/iMhrf2FY0WnBBergixZli5UvaRJ+/mzy5QrmFMuwB1ByIsIo0h/164x61zu
UwgBSVKrETE29QOu8tUHlL7lL3EoG5bCGGgN23Es/ohFhuRSN2SUvtuQf3iIKCme
XRqAS7Aj+enwSFriIdUR0qwtsA0jL4iYxEHTijKuNLqVZLykKK5eVsrVnNlggWKK
`protect END_PROTECTED
