`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iwo6LTIvX7gVXHlRKH1E1aQobpc2KxzWLKeng8f1bWWCzJ+zTTE38xvyRVqLvhCe
guj5awJfTCcmoVreMzEa8BxKMSsMrrJrtGzsAlXlGYypWkWbWvDaZ0AH/PKkEQfD
S+GyDUuZxGujLCez212zI+/321/eQ65s6W3O7WQBqDioLmfxcTp/t6nPgYUuJ67E
3jDcNTrX43UcI1kjmKXR5xMcYf4Gv7duCCfUob2YA2trWgXfROc7CSdce+J6mC47
h9vQSbqZBV2pGIrrodf83cm3JTui8L3/j2cbSM7KAzFXNy1fg0FsV44sam9+hs5W
KGXZBxyZ0zWHvcCziD8q/xvPkoGHEAO9yTeCKGgYeMcubkWQCZLA7pmtPfFbctK9
LFQt7c7CiQvAQWA2xq2KhQE6kbGMj7RE2dy46SmVI12iiq4pDryU2epS42wkI5b8
BoBLlkgmkr1K/L+LGu6+kI77fhC+kOdT4KeUijuG+BJEP1LtZ965inJDlbfJ8U1i
TzHu1b+KT3YxARqnffIrrfa1dtFNpt2g9Bk1SG2Vx/jfWOHYUvhzj8MVutk+LpTI
KUJYZrE7c5Io85uXK+eCniDRxnBO1P+ka4VILyX8Jfz0W8VSIs5potLG31Fegd7c
EOBnF00X/RmMGeyFW/m1gG+1/UjIzth/RyPaIKdq6Phcj5815nj7Ifd8w6z8lXlM
hmK2Pt4SpBQpFVmY6Sx6cWeI9QkY3GyUoP1jDUkTVX8t5TmLiPSP4pPjz3jiGs30
xON8n/LZGsEMiRaTw9qVl4NjWvzzW871f6RexoF4pLTpvVSIZwwkazu7QzUd5/SQ
2XzOANb//Y6H/ZELnHyIPRyAeonLuw8Ub+u6HHkXn70=
`protect END_PROTECTED
