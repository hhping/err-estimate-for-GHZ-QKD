`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meDJaIzvE0pJE4NxWDrcDU73DTpUYR8ElU4VuyVbO8qNt6OhUZ9uDPeD0HDCkMfB
W7f51n+Oy25u5S0UAo04PFEpOswidt28Y9ZDPoT6aarOfv5Foe0o+WIihOWg0Y6Y
k98qAm+seJCRAkzF7+b9QsFjg982evYlfB3y85ZSYwUqGk4pnNJP/cFhoScfJwwR
5eEzy8bJbktlS6xFo7Y4j0Q7pHT1Nk8Asf8VOfgfsnku0WRUPYx2l8o/Iyx7d+Ej
6d9QdsTH57ZB1XCiOi/DSFb8qlqZEyJPTi6Ubx5Z/YHKvtQPXw+MhrOKlEG7nt4S
wOWDvG1ftakke/oF6S1pGr/KQ6wRYRVLmcKnwWYjIYBTKFefeD5PeqHXKpwTQLxY
QzFhIER4ablInp/2JpvYRvjpThpDe1akY8rr9EcnPX+Fxzl6QVw8yxQhm0DNOO86
TL7X8oW72L7mrNV17nrAyOxBkWN0TKmaUQdOQpZn7HPnJo2mt2AddLGMSFpM3WMw
sGQZA74j8zCNIIuO5au1WSLgcKQt/Io/HeBEFXQZY5GuCSmBC79MQ+CeV/R+zFFx
edC1FBUtGIGTuEH//ddbqtvSYxyz4v0qP5eZjAgNgnp3nzt9tmkc335VqZi1VK25
BdJOZi/+7Il1VZPuQAE/GM25APeZueR0de2x+R021OkEVh2/B012WlS5l9tdavqa
IKIC2r7WggWInj0gXSE7DU4Kf4nMQqmLrhYk1OONHdqi3TslDT7mpO+kbTPdJMQK
oJH+6oHyf5WZ3atYHgsIp7zfBE5QIB100rLEEwg4GmVe2oY+Jzep5VTBncVuy+re
6zgDbTWzBHUNcZFS5PEyxh9wn0sO0AXZQq/sQkB30itGdWMhuKHRUC/lIIdtriGo
hz9sK1sL/kbuEJGgxO5EEQStH1eKUFT4OwZq8kTb7i4sGul8s3DHnDDwluG+/7XU
c9QaxJarpNRzw+vXWGOJt8Gpy9brjtic6PY+4cHoF5FYTak11/nURnxW8gISwKmL
jYmj7Bcn4GjhBOK5RLtnqOh2bhVNY/H/npUmv2WKzvt8oVWp90y2E/cD5gToCZxW
HtQfX3cg7vQGlgPdsjYRjX9mJiFHcKQlw8Z1qcJzp0VtyXr9/+hw8H6ShQdL0cmG
lBYaV5WK24r1fTACegvRdFlJtRhKt6Lnm837UVNTiX3vTLDP5hKYPkOYXZJn+DrC
ZVrGVrf1e5LRoLJjEkU2ECgv0Ajst49MIf/a920dUIVNpkLoa+xFqzofMwAqjIXC
ycJ420GCaD4b9oJEj3OUxLdcObpdD0bzgqhzhbTxUzhsVByude7owNp1zEGphGzO
ZYrbJiLRAjtzB1JurMKKJ6+QB7VS44Zo+3VGSqtCNWKPCo1X8LTo1S8Y9C07fxtZ
1tmfXR1JNCUwE/yGzKR6tr4jf6TpljWxgAkff1TkjSnxdHrsRtd7d/8ypTSgOmui
dw3riqszpWOm3CeuSuMYCmvzDSjMA2yCFHNsKRDijq5+DBhoMaJTWgpMKfBQkD36
D/aKjMsyY1mFtKK73xVb8piv27iEGUiCbq7sYQtC210Evzxk+jaIIvHrw3jzO7dQ
kL4zXHRBpm3uqC/F0+mF+P9iucFkRxi0SzNEV54aMxvsZgoTkNOvJidBpT2wT+Du
SMpzadZ5nVTcE0E+kCb8KmYVe8ZRvQ6+s5ElpYWlWI782wLrlAKfVaL+rgZbO2CL
bWu9n160EvbNTySOzQuzLvt/+x7HL/XXNQJq0P9sr5Q4O57YVmGcCIsvJEkwWq6d
lHeBsL7c+1UYXJGCHRv9SA==
`protect END_PROTECTED
