`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/bexEvGdUwif1bAYhDKTkDRQeY8uGF4nG5rjZ/aEle2X5WgPFUagJZbb3tdgC/7
U4yOIYYriKcDwlns2Uc0ImnLdxAPuVf9g4g3QLo3u1zlTg4CwktOIY2J0sSg6WXn
33iESknXtkWJ1bN5X0I9rW/irWu0hQn3KgK/TXqZtqqz8Y5UsV89JDn21IHo/bLV
0+2vWbdfMuVu4Fi7ljzt8nZ6qfmtmG65oSpp6fIDV/XS+ENHS9GiyzzwWUQQOz9+
cKxGu8drifYC5KQvyNgXAAcf5jJ6YJ4sYvfx/KFCkUvshZuisaGOIKK2UdkfDAeE
UQ7sfjeZU15Q2hvnkF6JqiqLkWuXDkzOsaiSOb1N6DzO8OVvM5z+g4jxWL6pFB2L
RRVUN3t1W5ZvEHiellQRGlESwAqFC/8mpdo23Hs45NWGAj81AgavSLCID3fWC9+4
Iw6e3XfnctZpDK6uLARyB1vFAhrfnQJQokr1ogwH+ej/NEDgiM4/RxliUNV97968
la0OByrBeOKptqXPGCghCCQkMaX6gplRXc232NKMeHzJL5lv528nI64JF032Fmi/
HGh8sTzcKPAbO34BYiANGLrFWQ8WrkWRFveLEGqyCbhiNHP1QIWC9POpfr/TcesC
5NEGa9Lej0do4Si17F3rpJQhWFSg+fgSn3776436lSPMh9asPHXj+rd56HFyizTb
ZxIY1sHo9/wn0Obs73iriQxJIB5RI9j2MgfEH7/COST1efQfomlN1ckQAqgNNrmw
uh+bbaWWGiEAiZPmzFF52wv59AjspYGmkwo8++tKBJVMFJBOoyBQ/y+egWFGXsVW
TiwCijuAaPFMUsSq0eJQrMcenV9IhOGViQDCgxEa1ejxLY/Q/H58YZpxi1wPrjGS
2tW2pu9FQSmUzsSLF9U/qua2GSSH5uoB0yCVW6mbeDFLtgP1/PrN+8neZFXeltuE
vZ/efDANGsoWi3nz4w0Dh2loy0Ysxf9nsSaMUrNcjc6dSCmp+4WN5VZ09YATpGhM
HNWrAfzM89avXj8FQ7jQcbQkGtGSVe/HZOTJXvBQo7NWPxGGPg88cmxSline31TX
zkCr1I9UnSOJwrAuR7qf5/IA3PdQmO3hca28v7NM/xSgNDiLmqrz2bffRB6Rhy33
WBI57W/bT03wvb7NSLLkVNQSKnZ6opWFCT5xPht3LyvykqW9z4it6T2FSG+8Agp7
6Wh0Jlw3l1C1L/CVzoTyxGfNALyCYWCCFVTuYCzBH7OLKch0Le/rEvE6lSVRZSuM
CbKRZvI6bvL2VNt6zUa4CabawrcPpmU/4EhwWcxQGiSNOv5zoGVjNKXAsmf9oqpt
T8Mp0Ds3Fya0qYjNSn80y3sJ90LkZn2kzvG0+g76xzEKpGwKg1GDG4Fe54zNAs87
vOl6M1bkq6Rupv8QGx2o9eNPu3BPradU80X8FudPLOrKJniI6vC0erZO0KNcW4Fv
7GBdBwrJcP/pi/vCS1Z6XexxGc8o2vfEq9vx9RHcOIQqfwDC6UusQ6603AjrLmdy
YLz8pSJVYO8L9lSiMqR+rjyxZ6n2jEakkDy5JnMDL1mhMleF6YSZtIQwVfYK0rfv
s14jiUdSaHaNnvIUhF7kenS45/XkKnVEGZBWXEBx1Tz9IjQOvhUCyvDE4mlD5A/v
6eyKBr2xwa4Eb8GJT067eSJj7DzFxINJU1AUBa7uDPwFc1ZJzKIROZYGkPqTtT1X
rUHpau8h+BPtFKdKpRmBP23YmfmeeucgZVyw9jm3DJAS49diz6Du+5WB/tdAo43S
4uS+KXdyUwm7Tmr4JJWOsPO5OUPT6dKovbX1COy6XD37QTrG8Tu5ZM0IUQ7d2uZL
y9ulZt3BtUyn0ODXkKaOwPxL6CDcmtKD2piHDvAOJiVwek+WuUAJNvGTCRZD/CHM
nM6DkJF5nF29eByilsASvpe3EgnYotC805iFuso+JeODUR8gTi+Pnz4xDqJVJ9Dz
VtGwcr3D0Yy7skcXNxiweDWXwVeNzhVWDK7tW1him+aKejZF/CWBph+kh+3b7NSs
IjqITUfompJz3fI2rQvL3xbE4qfGPvG4QpV3iMljASJ5yT6b2ZV7pdELLGrHg7tg
QrkBif5iY07bs9hrjXoH2ikw0GtGdVtAlWs4Bd5B238q4J7nM/1QLKE4xkRAsU4L
iOGj7FE87qB8fs9LxafHtkViwslmyC9XNmYp4tp1vyaNiQDJdXPfiAU6BOtjv6eu
1ZvXBRqDeDfTb0BSqFaoucjaDXcfdO+p8SUP5szrjH57P06N3PRAkwbnNX3Ylwwk
VSGczjgn/LH31tLxRa3o+97qurgFECVKVYrwgujUMAgMf3WjJATP332cduyzWLiD
y+jojJPSJXFole3O/ax8uHp6RI37zyex9f5OrAsQQ5A7Tfts9+fIeCNk7+V/MLKH
4kwmV3fESOmse8gvIV0ELQC2e8hojD4Ssu6t1FZ3WTD5B5p0w6IaBMs23Lv1fCzS
1rZTL81BbkAs6YHG8ewm+NQO5v3baFlgypE4jaDLPUVkn88bwPekpeNrp5dU5JSG
cHtIVkyjREd1YCJzg6cirXvCVfQ3ardH12HumO8c88Of6WzU8it8HOMmtCtJylpt
dClzt8s5ybHieq+3n84ewxRCcQ61swC56+zDKSefxbAzrUlzF/fHZdj7tddRXvkk
REgS79XCKQn+fyzOvBv7bcYUh1MYIFUufJNuDtf7q09R9tjEuXOSA6JSs+oSAro6
Naev0bfBuQWxFTPjSUX5NAda+85x6Xk68MSEP6Zv5sG4vL7Ix3UhOS1omqEHObHX
jW8wRCemAg71pS6S55csjUknpPlmCN+XZ7/jFA4waUj6+2WLeRnRE+uLsCk3VozQ
XQ2pokfQLe9dklRVCci83nLgqnn1uXri6u8LIyF/Tkg//EEfyYTrhKKVrPu2dwkE
SQwPbKZmUZp9PnSCmvus++lRFu92jarE3B263303Uxik78xV/eWIZ+2Jnm0S4YZS
TWcfwb+OhvuXdTAhVsDJQ1eFReD35DMPTOF7QkFM+OwXdNZe3Bs7YUlcL2SiXHyt
upuz7WIp8XqXGfNIqVCebW1E1T5ttBvT7Np6NPYp/On6w/tteU3x2bgh86A+jmOv
Zr9JBZ+IREon+3dwSonnxAMSIwtZ9bGorcxSzBlAVBWo9DnHIEU2kLS/Ey/6nhdT
pMbxwfKlPIG9C+IHwO0Mw7Hm1hXS1mrZnk+y0T0mxAa5LiFL/winemw+MIg7lLiH
OPaBmXmKYNsbkXalLo/kTM3Bo2o8sYcRRL/K5sqcW2y4qkEKFiesg/nsVaxEVd64
cHecTIa1bfy6zFJftb8JS+VyJxjpCejb1hASVX6qpIJGcZ8ZYOz2/TuMfPuMjfCT
h8ND+TpMkpVjc43IMqzuifYdleFjvW1JSXkNAWOJgOoUH0YWzPOKjKA9Z0B6SOQD
7SymMRLJ3y20cyblAt4pjibXau9n2qNiP8sy/GXA/P870yiGgW+8qZW0rQxRYvMo
UcW8ByrgrHC3iz/BrVMW2jV5BteZ/56HKZ7Rg8OjC2tNUi+OI13GdaCwmc3pRq7O
YLg6VpyH63/UaahMPD1rSpt3Bo7gKuwconf8WiJkJATmOee+egq9LXen/65m3UIN
64eQ5j6PZPJYCBvOgX07pEQBNMrw+DrdmcPahC1FL0/07likyavnLgFHDTcvbsK9
e2xHK591tIlE2EEFwcc2nB+o9b1aAUPhCRJMc2ik5pe1nuIYkuk4X36so5feuKaf
wqObsyULdc6j8gME1Li6Qw8Pm3JeT9uxMG4VcBwLj8HXXOKgMgpTRuaJgy/agv42
YQ2VcehiprT7Mre53FxdPx+jrShnm+qj8XWHnHVW4DZS72iv80iq0uOoZMaECJvM
79yqSMA15onRBwkmipdVt2dy/5trq3Tz3yBh6kHXGeOyGjpLXOo+akvQ8sbFPYjC
wSxonoWSL/57tY77YJ7dbAAN9xC3ExL2kRnc5jiQ1OFkZRDenS8roO/uvlQMR9EP
dXu3uG1anVA+nvJrYmLCome1A/21hAWW5kzxTxSym+kTDmVHntgr/qR/eII11K5z
SqX7bppWsZUhCL2+aZtLySWwL4xE1/1pAgbHmdwNDYk6ejv0duAx1Ide5FRGfTpF
20AeNk5DWgycFEm3IEk68o9NvdRjDLzPAA13DqQE0N6aruIwQLXD7h1O4sSPL08/
KWoxQ+eR0L9WZRLSFFS4Q8iHB3+PNK0SMZ1ZnepBJi3stiy3YSvqwp0UXu20KYoD
/sYd2kzHYhT/O4qWRT4ce1cToVGmygtfX63mEjh0g1eWO4Xp2bmIp4DOen1zprF3
ZdXakijwG7QCvAz0MENqr1DYrw48BAy8Bk4n7ysG/VSMYnHb6N3zSjG8B043/3Y8
ddMsmUcAp3VgBGUMxtClnURaJBJknMsS6TsDFP21pJ5e29cY0+LPXo1ZEr3rYiZI
47Kc03o1FTqqIttsrG7nX3qI1iXL8TO/khaVvLYADQriN/jlKlS2ntPTjeZaznKb
uiCVE8EqruT/0BDyzhIL+X71hN90E9jo+cJzF2Lgv/hgSraHamdvEncF11lteEa/
maSBQzw7EDBirwSeVGLeFURMdN7wvmTBsKoU+82YN4OZbppVBtIEQ5Ro4dycSLG2
0Zmm7OXysf9i/KEDTDID/9nLB4dMW6vEU2PNU6lDr04FYM9CnMjxoNLmfVlDUzjf
88ZjfFjtxxhgKsFS6wYsqvwbK7fEd8tqRe4A16Vbh8wGSiuoqCs1PG5PA60HHnpa
Vs6qBn+GJ6s5XQZvDY69LHDohOZ+JZEwgg3yOgTMLQY6KdK+6FpBuyHMVHGUlb9W
Lf7rLToZ1dsHMuZFNYTziqJCxOID8e1Bzwk8vQTYszXcHc6VKl7tcxvps7kPlgvW
AH7PziAHV67CPPes/THH4JvIjfoNKGNtzvg5vc3g7DmX3hEbqCrfsxFUnW1CUj9F
jUosUhENVNFTW/sqCqdImKMazho5UNiQSP0uKW2NLDqR2tseBd9Cqnfg0ILk+6H9
UKcsZWfdJX7D7lGGiPrTbm2NkOYbVrhQ/P+y/lSBQZq/Bsky7dUIRxYQBOw9M8NP
yxJiNJawnTGS846e3C5V7BQLxaG53N1N895a8lJrHdBn7NHxGK5GOOcc1SmWImIF
m4t/47AUdz/PArakQj7K0SGt+khyAZR4XjNqetwh+NMzzgcOWvSw3/Uin9xu8Ifg
zU0UCgHXsquSB7VDz7w4gNXUbJWgYNZhoyCl+RlZlGJvBnxuoHCG+7fd1PufvqHq
n3rAvCoskNFY04IuYUt28UD8nRyeXuzDlI3fnZuKzRH4Im6RWETmGV0yCsPupFrc
YRpstzD4e7Jun6PO+80Ju4L0W6lQCImZCMqD7OoQmoRxbp5lKBT8RYIgp3cfa1ES
GensxVKb8Ol9aAA8qUgLtgA+s6Bhlv9s1W1cGKopiGlvCRHGef0sqc1BLxC1vK3u
1rD4pgQkPFWy+h6G1BFHlbAXYpE9F0Azyk/TgLhhppNYfrsNAultbiFVifL0xfEs
WQqFqzJUKsZa63onT2Pf+JIlDYesrzUd6dRUghkLR6LJYD5D3x6vYSChzzOl2HPr
Oeo5Dc8lChz4eiZIa5RDpPiucbMQL4n6NuWm4ETtgGJkoaE3ABxFsIsbV3A1oyLv
25B0GdTMaIZFcTgRsv8SsgSQOPiKEHzc50y9GysMbYBZj4MRDQN4xNBgh7q/CPrF
TCxVg7mlQtgUQY807y1ryWvChpuCK8GeAjPIW+iZmWjYIAsCvdF8qNn58Fj98ol1
PvqJ2FgEL6e8r/xmG9dE4qLPC6jkJ0Luz/tLQr5/OKwwbUmY9VA6KquYuwRfpa0t
JQKVtt588q8Q7LSAHjywNJiS/AVcSJXabZT7y9pwnbhZ62VhVtaY6pKPEgxwXAGm
r8FuuwQMW3Ca0GVsfTGlKj7vDklnQuY7vvyX6rXDNyEfVnj85FQf2WiPKcKiBwMO
e7InyZv1B8fpvDDWJz8cNdtlNRuuxByV7+JYwjEAP+Oo2AkGwfav8QdWpzeHgTU3
w2yiwfFVEYfIXVRYqxnJ2I7tWAwyijl+AmPvQnq+MCS5Bo2B/f0dHfdbjNvijHM5
xen5CerlLl19PUZZcE7AgP1g88oyQ77gwPThlXwP9hxFVZ3Zlw2+DoCuhCbHUiZQ
0E/oC+PNbYb4tBkW57n2hDbWsQyJ6uMXV4uO1DVRVyKTHSm2HRz2YqSe8oRHGPEU
0yYc74r2wR4V0K5f54x9J0b/CMRnkCxf+7dBFgx4i1M3p+Rnh9VW8lJ5H1rTF3MU
XDCm3SZp48fN11lh1CeMeoETBCd50W3/1cKXrmvRypCLk0WB8nQvyAszd9vg0+dZ
7JoOm2OcuerK4wR59Xikc6kyi3b6PCFNZsxRfk+c7UID1Ist+jaKBazAIXd7yhv0
/pqBbm+RICHMyIjVdxsyEG5mkWt0KEya/zUYtUKRt6mj85kcKwpASKcTFJkGya85
8CUIAKdAsX5aJSMF6D+lXEITftcE6+88X54qxeUnB+oroVSzZFt2iA6jMlPczsfL
7r/65G8vgg1XesUXxX+DCOZK5mkYwxN3NANmmeQCmRvKDc98dyuDlw1I2glCVvWQ
LdghVbcnkI1In546qXGTtuo9NwHf24JJThfGFdQ8Wyk5fkdnIKpinBJnGpGfnvHZ
/AnRNvYeUN6IXTG/4Z0Ng1Vw/Fe9zeXt37PvP62STT1T/HICNnTXb35aUd/76ECm
5heueOnYLXvFGA/7BcKLViNXpEft2L+HGBjj1Vr4htX6n+o5H1TcN2aFZdRdDggT
ejAxjqnkPgDCDlCkNs/yj2n1TjTIL8XOhIczyCsFa4Wjyocxko7L/V9CQTNl3VWk
0zqErPhh5sjqQ7X89cOycDz+C9t9uOWP+ysJMQ23sYXlgm94vh4FFlKlGc4FfVjk
W8AsRajZYFvYYKUrQogSPiLF44MsjYUoD/9TEIb5pUStEb1/F2rJXxR9K440Y3AF
7EMByFnnaQg2ClLLo5cI94PFTRCqSz2bDV3Vz5b2/6zKQF3WYVXQ3RW7ahgF4/M6
gRmulCUMP0usyOvRzCXRMyngedUab/JVzdjyvXjw1NSERGcQ3tVtgS6vO/7am9bA
4l1lmO/cPOyinoyHKRACvh1dcJw6S82l1YUmc8COPhCGN+8MZonNAo9kvnynSKnB
5G3FTPYBfnIaHJ8TiFo8huf0FuZl1ajEIkk0d3NTOymSBa2mjZf5qq1yN7fnb7fM
FOAoiXbHmY7KG1rKkhjLZMzMtkJy3qD+rblHD0hxnG43Hn3ve2EXZD5NDVo51275
iDqc+G9n69UhkSf/vKEkuldleEDVRT0gMHpjCAEVrJrp1r3BS6XAO9h455pbsF+u
NnzSdyZLJnN055SY671R2jTBdfvrXK2b0d9FijWio98T3RPDHgbIntusm+NY+vYF
/iTcRdVlFIv9Z/EYzudd5z7sJrT9JaWGhq45u0u7FAdNihGtbYbOKn5FZjx2wuBW
4DKvRzNhGvTvNkE5EhrV8riMggDel6gKKKNgfHR1XGDfcFfjp7yzBgy5SMrmqj7a
xxYRI/ik13XYsr12zdeTwrbCnIdr6O3w3Ue08k3ith0lGkfr7F1QSUHC72jZRnW0
stUx9G5N0BjeR72wOKDHNVnfWDBABDlda1pV/U9DVERCYdwUymGEwLcGiRWsWr6I
Iy8iwvCai2BJHDs52hcVLM+rUiL5szMJM4K1aEbzwFmoOl44WCwHEwVKJDFxdZjP
HHb2ZI2PbBdslCu38qCskOrIatL6Go7w4PvTMFxCiiJMIV1ANjXmuvQEDJbeTxGr
5HdvSQxxqJq2KVjZwFVRFwHULTDJqLKKAJkjEGChIducthoLYfWhrCtzc1ja5n3k
mhopP9DD2bQGZC5MNjs2gQ==
`protect END_PROTECTED
