`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXa1X+reMOJ6TM1grFv/rMBhfIvChWg19oRXujf0gk0+K7iXqG6TgSgHJLA+EEuV
h4rmGs52ZR5t7T/lClNWX+/MD3KQqYhbZEWQfV1T3iODwAOqYJBfOs02lvANTjZI
BpOgSm3OF/bKezRDuvridTVGjsEMv0nJau+QovSNmRmnUFT+taW9jX4iUOKVe3pq
HQtqAi6tT+lK36v3lHgSMbjOLyP6ZXV8508b1FpNK4YR21m31WkrBx5qOMKKlZY+
mjr2kt4dCw6a5w6vlvkLmtiLxj7GEvsRXruSpwtVaOucBwB+j5wjnEghec1gNpno
VTKzJ827dp8QdxrAkuJ1zMduQMVPUQi0+CfKVTRuUUW/GOmibtdVgL5NEdW9JD2n
EDtbLkXuX2nzKA5jkjx6VelVEw9QEw6Zj18QqB6/+6n0RzJwu9HW5h0qWtek9xls
xSsXzcMSVDBRNglPDIAg6XMK3Ewg2phuGS7y8KlWhTF31Sy4zixTl1YCwcr/NBGq
4Xu7LLfvzXWn9BHaC+RJWoseMvpB4YEjGoJADd4pyxpf+sq9jezwWQiA589AXqIS
ChE6e1ivMmaqf3SrP8wKQA4LzJMbc1BdgI9FwnhwQKoC5iQckrc4YXzKaSUlS0pG
Stk5yKl04qvKVwCyi+KSXgx68or02U9gAmUOtR7gDmtTHsgW3S8ye5kZ51oedLZR
t/JZxvZ8o53m7L9c3JD3EI/hRaMh5jEAEIZ5zqLngPxYcucvi/2RkYVkVUvCirZl
8NWyY7lTnM+PX4+MJdNAaiEYrLJJK5D8iVQzn0aLIZ/F5YsEgf117APbnqDCoV7M
WWHQiOIZOC1dpDxbq31jVxXkIOqhgs7jHq9TVtWipqIo/dqbMZ3d+26+jNjP0tIB
/wTvudqD1oFjDMSN9jwEby8SQbTFuB8eiMPEDfxTCTvWYeVcZ2L9eV1h3TAoSsvK
bXoUOacXhuvU7vvMqjowESgBPU50F+StvfPOx1iacPLzhg5+bShes7lSAXAfAlr0
wmbB6RbJDI9ZrolBAzzO21Py5qWdkzgVxXQgHYjMDbdxM1jPKF1ije/KTjaWsgc+
Vo8XWrayMUwo7ud5hdxuhuZJ81bL2t+hFrWKZUV1Gu7KgfGmVoPRl1qJpa6ZmaUv
PfGOQtXXjAySKODTBk/SJwPS5ePSumxE2czu3k5f7OaSMPMCaAfhKy/FBwKdETLh
VEgTr/Jbki0GHPQPs42BHZ1nIcv4/vVSkyF9HyNfMCAPgUKklEgwTI86OUsYnYxU
bSz550DO5mkGWgsFqm6HGIMHN7pGIQPgeCz2TEnDMlF2vSwgbPqPRK52rDavfbLv
muomgmFCxgzejdmpEv6yCFvDpgXKwyMluhobAYngdUlcWVjdm2Rr98Jjk5rCY+xH
YwROVjWsyh9G8TxFikjyObx08Wi8CmZQFhvCuuOCjmh2jpbbTV7VKOqWxk6VgEQw
9b9qksUVzIfE+CRnHtL9j33S+1vTXYClh785tdf3HjEwpNViOxhzUZYGFCbFnKSX
BQ8bzXpqGgA5eHORlUN2WGT/yt/EM8P1scwJF99vzB4eCU99DAfCSnMhIxwSKwFm
OJOAyNNY7on7IFW4rzhn1UvIoWmMnHjt7uyA0OPE9eJHv1QjPyZlcRDp4H6jkaCS
swv07krfPBy9CDrt9G6tjs9UD13RrG/PbxcZZzho16iXMaQibWpqU/4teVvexsnx
wwO4IZfvi/YAhS9ITidFdiy1u4RSybP/KUphhVB9dzPMYod8x1yChtKfJzShKSlg
7zxkoCAc66YqLFIHqdyPFQMEdJ2eQgbu5MONMUDlfIR3JihRtggtyW9lx5JQ1wJr
lyDvf4NcPSRWIAw9vPciX8WhnEEc5VILvNueNldn3BTZfe5JpFroOraI7TL1UgA0
Rl8NDyFsiTnes5NDuOwlyA==
`protect END_PROTECTED
