`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1O6EhQmtWJj3I0w6sXDkKKWj04hBQFNGNokmD/2dIHdxrLBaRj+uo3132p6s+lwz
cDRZjSMQ7v5ntkVDtG+jvz1Q/nlTNgiycoWkUnBE5G63e/Vvp4eeYRjsYgsdM1Xy
fNShD4uhqDzQ11whACpG7QfMjmtRszdoJ6CTe13vALnFWo7zY95fDXV0LRLonL5k
9H+x8xuia0rxKsaE9ZaVxZumGR98LXvp6XnZUqZxUMSXD+epzOCwgRClAV08BM/t
GM0xbcIyb70YrAOiWrXDfEMiiMRGNjhJdqns62SbPc+BTwBBoZckuT98frvGyOSp
4WlpIgaKEgivO1rfcEzaayD2LupDicl96cIhm7tj//dre+1DrGHxFXyVj2qLjNfP
7l7ri5TXGJmJB0tmPzOTHaIfJEe0c2p7OhGdHlFMLDY9xABL3EzVNbmW0lPV17Yk
Eq/wPQ2YTQPQbdHEwhAPl5uEB3m2J44/a6HRPyRWEw+7GIg/IKavmp2XBMnnu2b/
CeEtg2E7559YwU0lTtC1eDuCw8WJ073DqEkKkGSQv5qj2BUQbRounfAcNhSg+9l9
p1FkgFEzoRo9NQSX6xCGy/Z+wGdrGy6arM44nB7F6mLVjZEgJFKvVB+b3aY+dLyY
52IE45/Cgqq7SnvRBgYp3PBKkd/2g/Dhab1MoZnuTsqBGyvI8JK1b8tOSDixd0oo
bVUNOxgyW6hJPQRS2clP6j8MTWGKfr+DMZl0SgVxHZl0sGh9vnewgJwbs8COytLr
dmA16tG3Tw22c5QkRpwodhynLm/uUFUBwp6gvLbqLIldUo3bjseDVF/gccJ5uQlI
rE1PNU9fW4JcMPR1d17JvpT90MX7wHKFWBZ+n66sp7ioa09HUEFLDnlNYg9B6D2p
z3vixTR1dV1osLVITQkfSxV8XDxgyoQLMVM1wD4PUStfDEHo2Rmh2b7l5e5CbdLP
KbXMRYFda+kiH0bBnCPbzRhG33yvAoZ2msWBNj52ykSsNdf1vRwRYpCkRTj9G04v
ZtJZmp8ejzVbkd5B2bNgXCeAYpMxtB9ojHCbRWBfOAaWFgUbmEzaFqWenmFFXtQt
2ivheAE9o7hGfCfxqhujz1GY8/GS0E3DLB+08bHxkJEcUe8/8+7y5XE3A90j8Tpl
IIWc7NErm9K407bGTDLir3SRLziE2f0n2eZVkNKrGazOVoF5TaqGuAEcjD+CZuHJ
zhHpV5bAld8WHL/u7nYoUTvV0jCUZIDuMwEEOudyCnKmXtQKkb4kRssznav5Xxn2
ycAYWZc1QKT/1s5AKc0CCFiP/1DwrOXBJwmYKFr3+bVazahL129tzLKL6Ap6Zvxm
2dKR3ooCOgVEPrApMfv7A8StvGEcpxAWh79PVnfthzHL2+nP/+v+nKf2oG4Fr8Zr
p9UOeqeMCDDQvK2/M7sEB40/zdB1kSK8FQ00ApuoBkQ=
`protect END_PROTECTED
