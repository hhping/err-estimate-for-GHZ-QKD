`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TdhZ4kB4f+Hi10a6V++yjuzIApNty47FR7bjO+HbaKm/u31bNV2+bVOKkwrOlTZu
YTBFIMdwVfS3j5mxcYRg9UWb24CbKP6OrrEv7Zc2qvmACf8haR4dVNtEyqE1TnmQ
RsA2ViKNkEk+Tusei767fyLkfTM8oyw05aVKNB+fu5eM+lM4HOL4lF9DCj9FNpha
fOOPEsPDwpTXdXYDZiXXDJdOhi7TTu5kq2t5rByB2pK/7D86B1EFyc7PtL3Dvjai
UT5WkkZj/FQuka20vZeJuPtAaGArSP76m2w/2hNvQZ2MS0DpiUfJA3wUWxNrNC24
r9wk4FZHSetACG55GvOxgc8Pe2JP89oDvkYbmN/50cb6hrH744KqyWcwyTk970N7
Zl6PcR4sF2zjHqOMttKOBwTkdZ/IzfjUJ2nerq+b7vT980LHICzjBqqEWngvLQGD
VTKZg2XHiRuCwTXQ1TplCL1sAsDDAGFpSLCAY79h0cNBrivMFtjoWQWrxxGRqTzR
65oQxr+gye4r9pFGunr3vW4aIIXO/5u0ABl3fBrmG91niqNn4ac/vCucvj1BVKeS
Giuh4V3iXyiXedKft1Jk3MFdVrGoNFJLFmvbeSGnGlriaHNOF52Er4JWDYcpnmvo
nkhMLrCZoI52Wc6iJdfkiRPFTQhmqQBGG6NpXFHZqQ7BnNon6jfhArys2b8nMQ+S
2eKBmOCGSSmdSz2IW52OfuhR4Kimyjz+Ef/6shE1fMUwEQfFqFeAmLrGUnqCwgk+
UefHrArY8PaSKnBFPmdoq6R4ix2gdIwqiyMpoCtJUyZLNT6SRoiP/ZfSX8IneggE
NfCLMbDyZKEymo0slRcNlXHQfZgMn+0Ckg3PF36Kunhvr2F8ZCSNf2YzF4+mQdAo
FeJp2CiVT2kNL6I6zrruAEKSVEWSP5SfAeb1ie/MsDBTDhGoSuUu/rdpYZ019eM/
xAS1X4yigO2xOhf9FLXyQzApxESDKbbkw37VC5ueH2pJLYMFEZTa7tfhv7cio84D
Esssw1pyVBo0Q90SheoLZtQgcvmZTt1tquAUP1+q/JEBEpApvuas006iPSwPNFAs
GuKwBsOjJ9dHaUOqWJqyYjbhL2AgEPkEQlwRY+U7ZyMVpW8s3RE5QSaVuklR+5yx
WLVbwhwYRf/UPtUjteONt2zSwh9+ao99aWhZ0LSZGkvz2mHZr556wd8bstJTDgCD
xTs2e1I8R++p+/zpe2dGfVjD7gLQGXq5EoJ5gkUO13q0UlmBMZ/u6shMzYO272DV
ct56v6YgwAJKY0sVfz3LUf4eu0b2Pj0SuztauY0fwEe5BIqMXyi5VPwn/8wcp+Up
THtb4qiHmMygAYpEV6NA9EtH/SNi0EUY0ejgBnO2dgHCCSLQags3rSZ1KYuiAmt7
/6nRArtmljNEQEF+WVFOhCN9QqJOddRbXHBCY+Xw3suIYDl9OeDuxtTM7utMO9si
gUrS3TI38ruz57KlVudyEH3b+j3LlaMZwCEvKcV+PuTdHaGGLiIKBFU6xtBxJmWO
76gfeyzhkr1yviNa3+wA41OMoQK/9RQT3xAWw6KpNris1JRTLpPXVe5wY8I7QzNt
8cbtGRpHu9q7mssxagULitI9gln+HVnQTlpI26pnHkVva20ccEhxnJksAgwBUmr/
SDLpXjv7jRIv8VoCn+KqOysRO76hQSR46sfcB2s107sIlKes3JNqhYzGmwvYAcNn
6SURZkVY82xcUqYx1D4kzA0GWvB6saxMaKAzGcg5LJyPrCZK529BpMmOFy4xJ0kl
z9OuCEwTt8jK1u/ttTKEbMoId94I6Dqphe0I1F2N02Y=
`protect END_PROTECTED
