`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKK91vUiF078oI/K0Ymub9d2/81wPkp9XP7u3/i1WtRv9aniG2m2vL13ER0pD5YA
k0sYwYrk9ATEjZoZJr+g+vAoti+lfbyRqiFGj9OnBGtsAbPYvbVeii6C1avzvsPz
PncXN98yPSBtxz8VmcccCrBos12bn9S/VV+N5/4HXmXxw0WkHaQDnt+vEEVCOcz8
/ZtxsW5DVI0o4vtBmhkjyYiz2OgWrmO7dWdD2FvgfJ68YTQgugZalNeo1Vh+8Dux
lZPipjff9cd73xMN71OEAwj0OQIyXtw+SEV9tx/QTyGGq+4gdGQBDdA0lnirOH5V
3ZkP2vI0YYnkf5RKv/Q2TRx3JtQ20YwvONO67ElQuOlGoVpueuXP0uzJrwpJdiyE
XC3+0AvFIBLYOF2gFTO6Afrr3W1FStqRwRgCfxBas6XVjI0q4YszhO/yU4rhYsyB
mAH8LkCl17u0QGOuHBW9FrKYQLiS+G9VuZBYsp3CdUU7+bymOs4eNAMarsED6vyu
XGHLI0YtGzve8jzfa9m/876qO7zEA2jhaER6ltEe2kqdD5hUgmSa7bRqZdIvPQCg
3pIM8scxvVJBNa79TTQL1M0AvrfnUQHoWNQ4zl5mJz6QocVLWIghRCMRXp+KmSHD
R8qRULWpY1ES7pGXtOHOcgyBQSPi+sbTp1usBDCjyJEgpr/hXRR/SiBo+99m9Bva
Ub0SK4HKyF5RY/3mZ7yln7Afk1fnnDLMyEp19M92ZlQclGEwAiq9JYQaJr9byFfh
KOy3QYD384u4nM4Kt5yxWCx++g+R0HwDP9Why1kuSiU3VrLLhiqo1bgJ2OZWcXGC
DewldCwt+YadY9J5jsPgtsh8VDTyy/5E6MxvkIMjG+JH7ikj1y7gIq7cw/Gzp7/I
YCgVDWEH8P01JiZ31dU7JYHxXQB0j9LJ6NOpM0JnNlU=
`protect END_PROTECTED
