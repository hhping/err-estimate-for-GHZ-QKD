library verilog;
use verilog.vl_types.all;
entity fourteennm_altera_iopll is
    generic(
        reference_clock_frequency: string  := "0 ps";
        pll_type        : string  := "General";
        pll_subtype     : string  := "General";
        number_of_clocks: integer := 1;
        operation_mode  : string  := "internal feedback";
        output_clock_frequency0: string  := "0 ps";
        phase_shift0    : string  := "0 ps";
        duty_cycle0     : integer := 50;
        output_clock_frequency1: string  := "0 ps";
        phase_shift1    : string  := "0 ps";
        duty_cycle1     : integer := 50;
        output_clock_frequency2: string  := "0 ps";
        phase_shift2    : string  := "0 ps";
        duty_cycle2     : integer := 50;
        output_clock_frequency3: string  := "0 ps";
        phase_shift3    : string  := "0 ps";
        duty_cycle3     : integer := 50;
        output_clock_frequency4: string  := "0 ps";
        phase_shift4    : string  := "0 ps";
        duty_cycle4     : integer := 50;
        output_clock_frequency5: string  := "0 ps";
        phase_shift5    : string  := "0 ps";
        duty_cycle5     : integer := 50;
        output_clock_frequency6: string  := "0 ps";
        phase_shift6    : string  := "0 ps";
        duty_cycle6     : integer := 50;
        output_clock_frequency7: string  := "0 ps";
        phase_shift7    : string  := "0 ps";
        duty_cycle7     : integer := 50;
        output_clock_frequency8: string  := "0 ps";
        phase_shift8    : string  := "0 ps";
        duty_cycle8     : integer := 50;
        clock_name_0    : string  := "";
        clock_name_1    : string  := "";
        clock_name_2    : string  := "";
        clock_name_3    : string  := "";
        clock_name_4    : string  := "";
        clock_name_5    : string  := "";
        clock_name_6    : string  := "";
        clock_name_7    : string  := "";
        clock_name_8    : string  := "";
        clock_name_global_0: string  := "false";
        clock_name_global_1: string  := "false";
        clock_name_global_2: string  := "false";
        clock_name_global_3: string  := "false";
        clock_name_global_4: string  := "false";
        clock_name_global_5: string  := "false";
        clock_name_global_6: string  := "false";
        clock_name_global_7: string  := "false";
        clock_name_global_8: string  := "false";
        m_cnt_hi_div    : integer := 1;
        m_cnt_lo_div    : integer := 1;
        m_cnt_bypass_en : string  := "false";
        m_cnt_odd_div_duty_en: string  := "false";
        n_cnt_hi_div    : integer := 1;
        n_cnt_lo_div    : integer := 1;
        n_cnt_bypass_en : string  := "false";
        n_cnt_odd_div_duty_en: string  := "false";
        c_cnt_hi_div0   : integer := 1;
        c_cnt_lo_div0   : integer := 1;
        c_cnt_bypass_en0: string  := "false";
        c_cnt_in_src0   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en0: string  := "false";
        c_cnt_prst0     : integer := 1;
        c_cnt_ph_mux_prst0: integer := 0;
        c_cnt_hi_div1   : integer := 1;
        c_cnt_lo_div1   : integer := 1;
        c_cnt_bypass_en1: string  := "false";
        c_cnt_in_src1   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en1: string  := "false";
        c_cnt_prst1     : integer := 1;
        c_cnt_ph_mux_prst1: integer := 0;
        c_cnt_hi_div2   : integer := 1;
        c_cnt_lo_div2   : integer := 1;
        c_cnt_bypass_en2: string  := "false";
        c_cnt_in_src2   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en2: string  := "false";
        c_cnt_prst2     : integer := 1;
        c_cnt_ph_mux_prst2: integer := 0;
        c_cnt_hi_div3   : integer := 1;
        c_cnt_lo_div3   : integer := 1;
        c_cnt_bypass_en3: string  := "false";
        c_cnt_in_src3   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en3: string  := "false";
        c_cnt_prst3     : integer := 1;
        c_cnt_ph_mux_prst3: integer := 0;
        c_cnt_hi_div4   : integer := 1;
        c_cnt_lo_div4   : integer := 1;
        c_cnt_bypass_en4: string  := "false";
        c_cnt_in_src4   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en4: string  := "false";
        c_cnt_prst4     : integer := 1;
        c_cnt_ph_mux_prst4: integer := 0;
        c_cnt_hi_div5   : integer := 1;
        c_cnt_lo_div5   : integer := 1;
        c_cnt_bypass_en5: string  := "false";
        c_cnt_in_src5   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en5: string  := "false";
        c_cnt_prst5     : integer := 1;
        c_cnt_ph_mux_prst5: integer := 0;
        c_cnt_hi_div6   : integer := 1;
        c_cnt_lo_div6   : integer := 1;
        c_cnt_bypass_en6: string  := "false";
        c_cnt_in_src6   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en6: string  := "false";
        c_cnt_prst6     : integer := 1;
        c_cnt_ph_mux_prst6: integer := 0;
        c_cnt_hi_div7   : integer := 1;
        c_cnt_lo_div7   : integer := 1;
        c_cnt_bypass_en7: string  := "false";
        c_cnt_in_src7   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en7: string  := "false";
        c_cnt_prst7     : integer := 1;
        c_cnt_ph_mux_prst7: integer := 0;
        c_cnt_hi_div8   : integer := 1;
        c_cnt_lo_div8   : integer := 1;
        c_cnt_bypass_en8: string  := "false";
        c_cnt_in_src8   : string  := "c_m_cnt_in_src_ph_mux_clk";
        c_cnt_odd_div_duty_en8: string  := "false";
        c_cnt_prst8     : integer := 1;
        c_cnt_ph_mux_prst8: integer := 0;
        pll_bw_sel      : string  := "low";
        clock_to_compensate: integer := 0;
        merging_permitted: string  := "false";
        pll_slf_rst     : string  := "false";
        pll_output_clk_frequency: string  := "0 MHz";
        pll_cp_current  : string  := "pll_cp_setting0";
        pll_bwctrl      : string  := "pll_bw_res_setting0";
        pll_fbclk_mux_1 : string  := "pll_fbclk_mux_1_glb";
        pll_fbclk_mux_2 : string  := "pll_fbclk_mux_2_fb_1";
        pll_m_cnt_in_src: string  := "c_m_cnt_in_src_ph_mux_clk";
        pll_clkin_0_src : string  := "clk_0";
        pll_clkin_1_src : string  := "clk_0";
        pll_clk_loss_sw_en: string  := "false";
        pll_auto_clk_sw_en: string  := "false";
        pll_manu_clk_sw_en: string  := "false";
        pll_clk_sw_dly  : integer := 0;
        pll_extclk_0_cnt_src: string  := "pll_extclk_cnt_src_vss";
        pll_extclk_1_cnt_src: string  := "pll_extclk_cnt_src_vss";
        pll_lock_fltr_cfg: integer := 25;
        pll_unlock_fltr_cfg: integer := 2;
        refclk1_frequency: string  := "0 MHz"
    );
    port(
        refclk          : in     vl_logic;
        refclk1         : in     vl_logic;
        fbclk           : in     vl_logic;
        rst             : in     vl_logic;
        phase_en        : in     vl_logic;
        updn            : in     vl_logic;
        num_phase_shifts: in     vl_logic_vector(2 downto 0);
        scanclk         : in     vl_logic;
        cntsel          : in     vl_logic_vector(3 downto 0);
        reconfig_to_pll : in     vl_logic_vector(63 downto 0);
        extswitch       : in     vl_logic;
        adjpllin        : in     vl_logic;
        outclk          : out    vl_logic_vector;
        fboutclk        : out    vl_logic;
        locked          : out    vl_logic;
        phase_done      : out    vl_logic;
        reconfig_from_pll: out    vl_logic_vector(9 downto 0);
        activeclk       : out    vl_logic;
        clkbad          : out    vl_logic_vector(1 downto 0);
        phout           : out    vl_logic_vector(7 downto 0);
        lvds_clk        : out    vl_logic_vector(1 downto 0);
        loaden          : out    vl_logic_vector(1 downto 0);
        extclk_out      : out    vl_logic_vector(1 downto 0);
        cascade_out     : out    vl_logic;
        zdbfbclk        : inout  vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of reference_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of pll_type : constant is 1;
    attribute mti_svvh_generic_type of pll_subtype : constant is 1;
    attribute mti_svvh_generic_type of number_of_clocks : constant is 1;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency0 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift0 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle0 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency1 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift1 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle1 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency2 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift2 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle2 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency3 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift3 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle3 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency4 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift4 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle4 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency5 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift5 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle5 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency6 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift6 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle6 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency7 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift7 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle7 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency8 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift8 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle8 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_0 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_1 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_2 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_3 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_4 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_5 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_6 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_7 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_8 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_0 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_1 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_2 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_3 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_4 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_5 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_6 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_7 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_8 : constant is 1;
    attribute mti_svvh_generic_type of m_cnt_hi_div : constant is 1;
    attribute mti_svvh_generic_type of m_cnt_lo_div : constant is 1;
    attribute mti_svvh_generic_type of m_cnt_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of m_cnt_odd_div_duty_en : constant is 1;
    attribute mti_svvh_generic_type of n_cnt_hi_div : constant is 1;
    attribute mti_svvh_generic_type of n_cnt_lo_div : constant is 1;
    attribute mti_svvh_generic_type of n_cnt_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of n_cnt_odd_div_duty_en : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst0 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst1 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst2 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst3 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst4 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst5 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst6 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst7 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_hi_div8 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_lo_div8 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_bypass_en8 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_in_src8 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_odd_div_duty_en8 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_prst8 : constant is 1;
    attribute mti_svvh_generic_type of c_cnt_ph_mux_prst8 : constant is 1;
    attribute mti_svvh_generic_type of pll_bw_sel : constant is 1;
    attribute mti_svvh_generic_type of clock_to_compensate : constant is 1;
    attribute mti_svvh_generic_type of merging_permitted : constant is 1;
    attribute mti_svvh_generic_type of pll_slf_rst : constant is 1;
    attribute mti_svvh_generic_type of pll_output_clk_frequency : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_current : constant is 1;
    attribute mti_svvh_generic_type of pll_bwctrl : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_loss_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_auto_clk_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_manu_clk_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_sw_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_0_cnt_src : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_1_cnt_src : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_unlock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of refclk1_frequency : constant is 1;
end fourteennm_altera_iopll;
