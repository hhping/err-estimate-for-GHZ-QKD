`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+t71nAQ6jqfAkYuuUj+zWeYynAOtMnbDV4kdNJjm9evnT7BoUyqYYl9SigGwvuv5
I1M63EWTvYNOYBULa6gahBA2Ui1EraeBEgj8lq1zNch0f+aPuYnGEyTDkhmBtywJ
zNaokkHlcp7Ji7JcgB3y6BRJ/O90ocLa0O1iklmwWMJtech7eitPLu76HM/NlgpC
HBQIrSxsO59HOEuFQedPl9pZzBrMthFnYuu1+zQJb9/Cd5/qK2m8ld0scPChoNXc
hlx5Ybu1hxk/QvFjezYcyRwSWFziKHC4dhtxhizOR+dv0sw5tcwdbw9h/AoQQww3
jLpUuRTLJcrfbcsAT8aSXgaAfsjtK8h/Xd3LmG+z6Y24zepK1vowmexVhbfUukq+
5UqePihSJotX2cA5cv62kp8piFLvPRhpTxX0SmivqOsJmAGxQfKPi5zBnkmPtJrw
Qt9bjfjmmwL4CD2JFZb3gj/v/iw0CWuUZXvVYb+arFt81rCFRangz41zRYwJJ6x0
XdKIrdd/t1NH+9qcKBTpPQf+IWHAWoLk4TTbJqlSqcqiJ6eE+f6ZUDmIDRSVruiy
THd5fp4BoLzjJeaoNs+ZinEtzzEWibor3AmnejjkVCQVbYmevKRs1RbH8jXRpz23
XcWdRBeAaH1A42JyZVeghFtfXkWU7yCzY+RBxvQ5gPCaM0nnmvKs4jWzd3ed7j/c
2WxGW2ZUQ2VVS5ilj0i5mLMNjpC5TehLUlJx/3o1yfy20UzEkz5j7JyUs6migUeP
IBg6tkOeWImubpwzd4yX4Yaq6XrTun/nzbnbJp5e0OfB4S4YFC2DDjsT111pGy+8
+bXW03zSVPX6o3bxO3CIhFZupfykWeWseTeYtA7Onut8UjZjheepl0bdnr8mhepv
Ok24OKFFxKAkukem7e/9SCtOaaW5AeQx+pq2X63HxdXz+5bI7ylknfU9cs7jKo+K
XoBoymd9isjLfDSypVHMGHn7+fgGHWsdQYzhlYqQz9fsuRGYee+HLga0bumQph14
hNgiX408+z0UEubyjwdfi19EDFD5Dxya1umv2pD96sX2B94hQaKPn872WCVROceY
bF/KzL04DRJAkoje7JoLCdqk3sjT6yw2o6AyhX/KpBqjXcQTOLlDP7TXZ05mvQpo
ZK7aBubMW/r5k9ln/dIu5XVVZMSk/6532bHFbFng/hKQngpxH86fYNuHhkpV/JLO
a8RTxVW7ZFIBwFDI6NOm/MVoL3DW9B0mzqT+iBXNvNBBHO0hhny/fVHJdku/841T
SKre3TTwrW6+XFw/bbwK9VPkbo6IJGYNoEbn39M+NXPETyAJWoC+WdHA19v+QzCC
8yIt5Qna77/6mqw7MrPVgjYprB20bYIjn/z9+5kVXdJDQBBLszT2tFvAQtVpS4Yi
jD01YahAcYmPX/3NFjdtQe9ZFS4XEyQtmWKNtdUFl5UKMPW5YhYqyaSMEspaJJFr
jaZ8wmJrYzfma3Nny4RQRnaxm+3DYjqg5CdMpi0S5POYxGQVE3RVZcYwl38NJB7W
/YieWVliNajEUthAPKFRpyMuot6bR31vn8ydCt3M9oyzH0l2DgRcPBlq8n9PcfK0
LQhmkTaApKpINnfHwhKUI44IPEJd+QG9WQY6DOV1UQLpBpdqRBRdthyQPLD7lDAa
+gS2xaQeWom24D4de88k6cvP7aID9Nn5BLoyOG2aLr6A5p/XtqZeumB6f/3PILhr
KtNbZu0FJT2HHE5yO3Kud41MuQbf4OTKEmknJxZ5mDzMqnS7OGqvl+NDqc7T5fz2
XYwiJZgxfGEavmRRc6WtVO8M1oRDAXPoH+D8WbaxRn+ZPtrT51P/I5XGONTg/Cz8
6qa50GpXdVbPmBe9x4x1PK1MdaixExYCrgyKmlrBSDMhas5JOy+n4hbYMW7p1+tZ
gDNVReJzILUsLxBAe3kIZOl6LjViYaMcQ3912SFEA0e3vZqBNqS9ffkru552hx6t
3Q4AYA5CdKmLJnuj9Rj2UBjLTQ9yAOPuKXyVeqPPGaBbs2nOX4Ct6wqv3xZkBFzz
awRaTJUa4r5cuosaYETmVvROHXnFYRF3AU6WsCeghLhJ9ABw+fGZzl1HlGUQP0cE
qFRvSGvOg142y/VhdHrD+IyfPD5EFEgKvKX11xsMDteXExATuphGljJdEg89RBFR
huTBeSecRbjLvy6kZdMzNMfcesgFSDNSXcuOWqzpaZuTzNBNwFg2tyngB1UTSLB9
4skR8Cy1jr+jx1/qHpxt8yCmsDX4QJGf7S7w5Tzb6vQQuquH/8Ep0Fby9Qb0Uvzh
b3fXJC9ZMi+V/MvNYn2IQaHB2iaG3ettbN5I9NGGNU+5uBMIcZoQ69BfPynPRQxm
Y9mm8i7mkAYR/+IeOacTklQYYUGAaE4hQh2FnkGMygs+UfU85yfYEgcoq567N4IY
AUcLk9P8SDo2SYZC5RRd2cUDI9tdHBoRxRiua7hMSCwj45YCuvM7098zSLVhWudS
DQ0nzsaEUZmmA2Ci5DRDMOhkml8QdhAn0kdzB6JCiDXIf22p+lcysKxuJD6sFaBr
XzzuM2uCzo1NgBzY170At9gdmSw2RkTJolpwi2jaGfsO0M49j9I/DTggdZE2Uoi/
1/gu9cReSMgVnwOxC4pnjSVtyor8JaFV2uyfY1GhOV8Ig7PjgG6Z/8u/XXso96nI
ZpwSzg0+tlfNy2nVulm0qwyNTRR0kE95y06PjHVZ5WbhEegjkbRsEaugqzxLRYgz
N2YpCcSUKNfUijf9dL9y8nViZI8EtBF1rArfil1KmZtvI+XGmv54kFEg1ub4F5As
Do6FkuBlEv3wg0YMWb3NqjKnvMe6JaJRHoD3pLQJCeo3WycbVtmQoKqcBM5TTpnx
sR/X3UQoMenxHuGI8GsTF6BdS72k6FX1+EUDlZk+O7TlSekkc5pUAXRrhYlj5Lgf
uLIoUJ4k6q6McORj3j52OiEUHNhFqXsqxzygqnO7kzC0QV26NoqmG4vJyjbXAhAs
QkXUu6U1naLNTcgZtADfXcZAQQoe9Cfm1VubZ9c0maFYlJRB16/sYbEjgo+GG05m
Grxw2+YoP3tPNQoDQ3jyib5eSggrdPI75e+ol+bAca5YpmzDwJRhLKbWy5kBDz3T
Q21LMQuXlaYTJyZ1N24jN/NuJ8i3qXog7SRDuEzuFqMNsSKAjTWYRF064++Twf0w
YhRBDmLcKR5Vacgxb0XdWAHVEHM5zE0zgKv7BaijPVCP3yyZk98TNHNFMN0ec1/G
lQR3mjsF7Q2PPw+F7VAMhtDjnPvYZrtoG594PanUD77fyZqltPorIzjvbO3AARPT
9LifyirQP75M6igFyR/2fgeDqzzSNnXXmEQ9aO8DwNiEv4VuUgz9VtiikmfmSkpN
OVf6yg/hQhUnVyocUxZqw+QfjJAticbkrk4Jk1iNFj3/aVikS+3m0H9c9LCsOmtZ
igciDma9EzgdNUn44KFDqXvCUlpRo2kUfsKCFGt0ZEuPB1VLGfYsTFGCj+8RBAdB
gbwStmxfLLIRvpDrWOQBiiKvU8+8q/sfQe8R37KmJ4GZRCYsVMcBBsm9PXdRCNMP
mYBR7mMoFad9YD7Cle8+4Q5H5qdKQzIfS5a7Et2dT4DSDpMDf1EQIYgyGBuPc1iX
P3yIMsePzk0g7kbwt6YAsJLpw8JuQ5FF2TMpqazEIYhCpDdhqCJt3begaUOYoGgS
ngcFm/MjOoVVqmZfDoLiH7hajEebk88j8ahTabJlZ3XSGyv90fPoXP+28/hHhlUc
kBKNyRBT4/AMWwD6msk2O1b6riiunYA4YOFg0dAJ0a54CfQF2bmIwj+Ev+3LV8cC
haS9idfOF60LOtzyDCeRsSeQWx1DcsmOVD4QsMRRv8pGK8jy9bG4A0+fgaxdUdGI
QY+gZ/U4PtMrJpYaUw+2NF5+YY4kQDcgcVZ1XFYkXDw+HLS5K2kFnyW35BdtwNlS
pSDuqkbqhN3ZYenZQj2MVVSE3uVPTrpsI51H7DwVJ4KqT+OSIXZVK938nrGvYevT
YzoE3SVbQGqkpPSdsWRDOrrknDPgZGcjS5BYo+0SiT6DzLz1PVn+kmPtu30hrhrL
CFUnC1XrgNWNOxWyGkwv6/9kSdWoBU0lgnuwnh9QngwrArfh+wTpNTEFciMfd6vS
fmIilWu2jS3ee421u5nLvDNUVgrY9TayVP8QFrPaZ0se08rJ7MRD3ys6zwX3PjA5
6Z7uo+04kAUH7Y2aao0e7jVTJPCrKGR5l2xiqUJoTKtirkn7PYLiwR5Oa7NytQtG
64/DeVKsihRcbG0PBkHyxggTUFTI8GiEafp5adnj0vud9vp+9iKLtgdx67MRR8Xc
88hlHja2/tXvlVMQWmTSDczg6/WK2qTS9Oal/UykLiPDMMtX7MhbpmAdVvNd2KnL
YJu/29feItb9J5laiIO+QhB9RXCRUB/yBwe68HDl3xA0ASjCSamRT78Fx88Xj7rC
XlGmO/WDH4WkPHeZtT0M8k/7s6fwS8EEKOPxB/+qriE6ESw5oFcBtDdd4REsfeEe
6fU+brU8oTaplH0t6dbeBg5a2a8pOaOguQW8r9h+Ur6PR6tpAUtclv3+PKX8vxjE
X1r5+lgnVt53Jg9ECwdaz0jbq6qYS5hV0i1TPX+RAyRUTg26RUKtbmP0jfVEyucz
0vuNv7NyEL/aO/rbiOd3AZAhKjC1J204vmVJMSfAvXkATfS+d4dB4tAOFPPB7hSs
232YmyRRgcQ7yYzwDFKku4kKJ16Syq1wjJFRIwhqmU/iF2Lj+j2gkt7dOk/VwgJQ
prfQfL89i9+rAputUrXDnlfUZq+E3gW2raD+xb5a7E0ClURZ7h6G3Msm2Zq4UqjJ
29mA1gI4hcXIOWPPXPR2zPFcMDIH1bemouwPBXtTVfN8MV2ZxMPmro4Pi1Ruxcdg
+wgjB90iWMulcQWMsIWtZUr9Pv7dpUPbKG1MRjF6BQtjh//9NBPipYn/+zB8Fgka
/OIMwWTBTaLKelHPbrYTZu7fNAcI29YelFYQuFp9xRqnsfZ8s0rBDmfbYhyZ/8ks
YgfVJJty69QV0tPt+Asr7+DCVrH8L8y4ktAcO7SU5ewSfDc1Dr+KXTg3Z/GsjqbO
TKIynozFHamMKBMRelVNH6K8UST5IOX+qGjLWcLH6wc2YtKRZH/MgZeaAQbvGrDU
UpyRaQUqlfaV4Ylr7jkNq60RTRWldSyJMdyo9ICf8TeEBGwvt9LBQOHagGPqdAAV
4UPYVkmQwpZngnVC/EVGrBBdtMIW/z5Uvugd2oKfgcRjrozx29bbVergTJ4fTFSK
plDZA5/flEQ5zCqScMdzPqxqAymx67OUTw6eL4CIvX1TnnZdF/bbY92UGoAW/Nz5
wCtH4ZJa2l5pK3Imur3OonDeorvgdpOelIwe4ZRpUg6Hq/Z8P9rLDKkoLP/GlRpv
UrrwZctY5SY3/bgDBEF5aHMdtuKLO29CigCz+y+lSXlcZxRLXYX4fOrGmU+SGofc
tSMq9ZIM5zR6Wk5qDGQJhq8KLWTko9o06Bvw64k/k1N5WxIUw3wWvEmKYiKejcxy
Uw4icRRUTOYjpLReLA3+xCPCqmeFiBRDDGujcI/G2eKECoGXF4F7qhocaCnJmVbT
YFSV3XGqEUvbA5TImBPEIP+IVH6+5a/Hu7ds9OqNSLLZ3Dvibs7CUS8zAE3BcrFk
Ix2f6oWMN8jOXJWDafZ8BC+tyw2wyofj5nhLKsRm+vNLaQNrZhI7sq/pasjYmgYO
WMYfWJUQfi8otpvP9dAsoTFJn93liUmEWASkkovNRTxe/Kwl7KTU7DTJUUIKaHxv
loCVf7OX72Mw4mVTD9OX69e2gsLPYfeFdGtqNfvlLz6IgURStnxgEeMHBmosrErI
/QCVuFbDeZAfF+4ti8LMHfmJ4gEPdGV+gQuel0rm8PuuU9209ygpTZZNOi5qz24D
JzP/Z1KLr7eNumjI40ZsDwNYV2ErV5pR0PWJO39N02gbGt+2ScFXsK5k2rc35uGy
ionaCe6TYglflsJyCJEmj2ND/5cggIuovsmtbzWC+hXDmj0x6p+Y4WvUODRGMEXJ
PtXx1io4+AonRSuo7D1Tbi/zLLLsX5D38n5lXSxZe+1dZ6HOVc79KDqvrsyv0Whd
eqc7fCIGBamagu9rKLAJzfDhamRSrjZb1pjBD8BEba7jJgOMyAYtBilsxNjNFHHQ
9Fd8/sT+QCSEbHNMC0UPmBzf4fsetLtgmCInokyrJF7cHeaIO0Z6jKLrqw5+2kie
gl+roqCVVmMwirAhPEuAuau0q6ZnT5NB12045ta47nv0NZy6MjaImItAAhJhMnWF
Z0KAIWxxmmyuEk8Cuk1wwZScL1zvO4O78lrVBfcejGWrF/cezdcRFA7HkLsTxBEg
DJ4yzoJrX2XWCjJQFwkzQPItc3Fq5aOk9ADqQqKkP++4VMhp6zQleKv+XpsKIPkw
dgLO9LhMw7uXrtPvna2yrnglO1/W+QzFMGFxsAZJMHl9I/dBnP7oGeQjE9NwU32Z
UPrLIbYquV+L2NCK4n2rpvLSU1gYIZoFjkWFLn+8lLEZQYHkfKPRZcKzaWLeB/9E
T8fz+ZjnQKvXyaNRY7YMGu71jWVwL502tqlOtfJgnDX8nBygtZLn/KiFivSp2u4E
Pw1oecPagqqCvZITbTATM3dsRl26F9fj5i9rWsvfXY8ri1m7Ew3CHxp1ewfOKpsE
CIgdbE3MhIPzTP5rnxmBTh7zLNduX28RsMPpGy9gs3iAcGPVISy0Xg+PgepwYQmy
nMbLRb8LyuJbivS76S8UAeMatunHK9TANdIenI3oG/S8kp+YKCerE/m2WCYnqJS3
1ERIc3w8XNoZr5i/hfCjY/gzsM0CDiRYYQqA/oDRMlPIV42yGgckIJBmd9/l1c8Q
EnW6/m6Q6l1OJfXqkE7wnLd83bR7nE6Ubjq5ES8K2EuerDHPiuclohEKYvBwS700
YrY3LOWqAtE9x7W9Tf3hm3W41OpYxkrEXoIA3KqWROqEqdL8D++a9t3n+VqBXbc3
owtRAVdyENHHSoa4Be5tMwbf9ZVYZItC2XzHXR6jfBKwok+iNOz39Ln4UWh0OfDl
AQ3o9kwq4eeIoi7gzqsjqQaFLRW3bvuIpwXrYGTPovutmfs88HEUbDDjAEzd42A9
kbKrzW8HoeOaS90hkF01MQYih8fCVM3tNVFdMrMkhcUNPm+1lwm9c9ntHM9il9Yk
TfzbaR4bTmJnjIAv94Up+5Xcb+QOMKK6HLVtKFlDOzwJVG1dr1jjfdxsX6/9kqqe
UoXf39krVnJfjo/SO0sOIKFKGrUfnTs12PTS8mz0pHt9khfoUpizRnIxtzPjf4ot
zmTpj1uCP0HJh6t9Dr58xVyZ9AMngB7Xbk4rT063HqXY+QH73vsaCGe+kH83bODY
EVqoCsG27B0OKcMWjKwOuuPuO5/JjWp/DJ/d4uDMy40b99S7HEO87OFxCz+X056z
cBtZXYIxK7n/a3jfPaAup8pcKFsaX4Nfd6i8hMz+41mKVwdnmDHjuRYWWnvQtAgj
NCtOGaytgyUt5F/QJZb7H6z/FSsup8bCgGcfBN1FQdq5y8CR4IyT95naMKjy3jgG
t0lJ/ELJ1R2TaPUqAwJNiK4k1GgrqPPqVFccLWfo96f79NUkAlYn71Yl9Mb3DQqn
eJ3ghXogXabDjE6vHwhIAAAfcbV3KEpqxc6scm6FGN7bHXC1d2Hl9cLXbjG+UFPq
+ODRM+e8xu2AoND/Yc9/ImFAmlPN8Qm71kwwu4p2v10/DUq8fZc7G2lMMT2kMkoR
sDjEIcSUwrCuBXwdQgwSzxPqp1culqdR+1PKd6KZhDABUnMd1Qu/qO3oryY5c+MV
HE2Db4j2x5YiSqUC0idXfHQ5Nse49iDWsXwRLI3AfAk6Xwn+zs1nuofMiDj9dSa6
JOb/yYFRYvdoGskbm0obptAC6LFI9csnyH6UfQVi8UsaYabO1Jg+llduLw2eNnb2
zodAqh8heHF0xWtqfFX5bgrcVrhEPoqGewVoMWbZ03sDw3eyFVQZszd80nELMpnr
kKzm/OOmUpl1ZOHbArIfsbqK/K18ZLQIXtpsBCsD3E/LAyGOf6Txs5HS7VF7Yet1
pum7miheUe0JgCK0ORTVPiHxRUZ5DRECANKrRNL9FYh60/23pjYyZgnSoZfWCscP
pbnUhbhcDrVy31OAUaHtBV1NrVKtTkmSeMBcEe4OBHwqFijgYYe9Dibe4l2Aa8US
AJHx+78MEygJPckBvMn4Wk7VJKiPTgwWMqCWjyjcXHTwYfwJMtavQxRrKmAL1ofw
LSNbDdv55kFqg866FsHKbU9spJyXna7fV5JCF8Szh6ySh1Dk5Fk2ZyLJ9aJpBTxl
wS/DD6Q9OWxMKdFy0J08KWmQsQ9xTMZk561bAPiBgGpQwgdDoo5I1/1gPIemUimh
3cDasgShK1INwnrinIhsV1ozQblDUM/Oq+ZGYBVPUwAjT0y8bKhrwdSDrPaD6teS
stBJbLmku3zcobD5VBJyyjyeZeJuVMdCdK1gLqCGOvY8tdBxstVqbFS9pwtsZTtl
2xF8a7VFIv8BWtwx+NFmyE2wt7D69gu+dUe+3q9Gnq6Fts9w5ElpdQnX+g+b31+t
l3T+8sAoqusH0PHv4mEdnzP8FsMK8cR9YnzRoobIuXFzH4y4Yi4yPQsE5bmXfCLN
Y9+R1oxjUQg0UZradkxNhFsOoX6flEAo0CdPEKyRo6e2OO2qJZyHTkMe/QRIurtD
BTh95YfY5mBTrJgXYZ24eX7V/AJvGwbgnL5q0W24k8Pbltkz16TH6W5PcQO2rWoc
fb+GHhwUbMD7Xyh06T155EMGrOHxSLDWNgkktMRRsiXXriOmfOjjaOyR9+9tlbal
jR8WoyulWNVnMVbHjuwY/gPjRg0pXxkXdw+Bf0VZvQmDVYUictKMxRplmRmo+nmv
TPreWsJCpkuG545oBmwndHEW6JgdZi3WMvVx72uy1ZWjecDz2sXYMelp5GPT70/3
A77YrqqAfxOyndbixkam5IaU81J/9CnzwqQtm3UieEPIYzux1mN4IgvNLpXIcWd1
FoH60LFlZtiRkSLEGqmAVgX5mGeVmxSZR4HRzQQkjM6STOuDqPrgMtu1PrZFHs25
Ai27vsHwWQO8rAv+eqk72TLtoUtHa1P3H8igGSiQwfMf2gsXtpRm2a5hfRpwHd93
F1rWxlDuq4yFDTL0T+A6157LqR1V0DqueiLlLBbdB44vxLk33JNpJV8BcLvc9Yoa
+iUpuU7vtV1Y9Sefu9FWOk+dssbvO+Kk1KAqQ8y1AAAYBlaf7Avcr1BlI+w5Gpge
uz9D5moqBMRzYgt5LHnrhkbYqelOfTkPnCKB0YZhMBoD3Yr/cj8oMxmofju2SF/+
3zLCzhi1OIeQ1ngGU51qvMgXEhQM1rAvh3z3/xo/P324hxXp6JJP2939ClBdAHLv
gHxu2vGtPbyyL+FOueEcW9jTf2WRW5j2QrHzNbeYI54Wya5fsxZi+WCrLB9ZbWq0
qXzmJQmXzUz/IY+/UWpgNA+u7zCZhSPE2HSyKOkS0OVOhQuHzL00uBKukF/FAsIn
EFEfnAImo/WA3cB0O6iqyA2Kyl7BfYBi+al3Gxax70FqrsrtV+yWBD0oO3nNQxT3
/bu54Sd73Z+kEvSFZWQDtLMFwdDoR51q5Gaiys7q9UCIfCm0FphTGa+b321alhhq
xDKHOINMkNVO1nxHAouIbskvrI5JtkWSu0LQIqjOuXAwvIaoykg92xsrzNmUQEvY
277FN6h8QLunmF3hd1AD0puNzRmo1F3QX9g7qVElF2IrGvGI1IYo3iWxIl8/xEhX
bXMMIzU4aCM+5Gb27QFtCHIfrslmQ3IR/SsAxioXS6r+dsMZ52H/ID51lUbBtAPO
ateF1DMhRMfOUIaF0NAZoVG20xGv3GCN4apGdM+a7cWUpS22SK0xcX+91XxaHOQf
TJGNrqUc7YkFVFzE+OR8KmBWroDt3GcaiAEPxkSYWYCn0QmK1hoyQAqIodfCTSOU
3sHWk189i+z+V0asfjhabFK71hOpe0Crw21eNI6/cfSrqqBD80/4SIljue2K8c28
KU0HR0TtGON9OYDTLA9q5ERsISUpELfp8uPL+FFu7rYpjOklJowoGdvqOIVUZO1r
t31kb0zJsNgaJwfHly7DEC90T2M3REKryy8MANycNCbdf06b6zr6PlKYJD/ahr5l
uilfkHiifZLmIw8yocfJcn0k2ADlhdudYFgEkR6t7bodECvs9BLn1eQrItMBuzRh
ZJxbxUfyOdMlUztquP/KEn9eDVAmd5mSybjxUCgL0a3aVlZryrgdCmlmcv1aht49
a2lMYGLuLWZhSfC7TWSHZdrafUfBYRm8x/y1NfiFcz2++nHbtgwKjzcLZh8UOeKe
I5SdOH3jjZVX1GqePBeJGK2wQXwZAOJMgY32FVaVy5Kdv9dE3bYvgyYCXkIgXahM
i5Hp9tu+mkBtgzoqMVeOtB8VdYVfUDR6XnsHjowJvqETDGnk2IdutzqPzVQvoUM9
cOzgFkcLMW0utRlsj6Q9hSdxjNBycca6rKpQg7iqw2taSjKRMBuZ1BkurvLO4OeY
NlH+ndUTgnpt5uAjQ6/VhY87tLw5otbeQj9XOYIn4NJ0zTzWxr+yyju3z/Kr0pcn
mfGMkiFXqOmW3PskrYOcDIsjeDwgmmtmt/aFwt6IYTcTt9ZJBLhDW01aurCkQaXc
JG+ibVZdyEkFouUSF/zHUsPIUufGy8+8XO2yKM+9atMuyDDefbH1Lx+jG6l4N6De
ZCPhDutgyZ7+MWKonWx3lHm1A/lG4S6iPJiIG2gQQyfaF90IwzMoWLd77U/Wtqdb
oLRZHhHW3dZVwzDj++zN60H9qflRmGfNweGp/Ifx08UhIxyMgCiABifsm+fHtz0Q
wr0jKQlVexaHtFST4dgIfVmgonIFQ8sEtwnStZvlznPVJxQ32DlUN+2dbzvceKs+
U9qe1sJJehObyAJ652nRbuQDxi8xWXXf/idnogGmLLx7XGYH3947+AVnla3ubQnC
nVWgaixysKMrSVrt1ZKI7Uidr3vlKjljLlPs+O7B1Pc7XL6mevCcuZmJInwGDPtV
tf373t1+4u8hVChLCDpLHrVVT/dtUciji8/MlyDVuTqQarlpKGq+DDerjVC3wQZX
P0gvBm1BvBKtOeV8SOz4BOm7abxbM/wLdsHoOYV17ZVUU1PcFcEdpfZZPB3G91xk
4r7lOJ0011wLG0Xq/uHyBdva6B20K5gPencgDUE/l2Vnj0AButjh8/bSl/gy8KAj
A0WmYkXJemt0Lhq2coXS3sHZZKze79z2vMJA9Jcodm8U+Hc2d4Ut4Jo5TwXsze8P
DSwebQ/3XQ8+k3/vDGB5i7JevTb7Uvf21VJmsYzWt1uk4NFWjucRSNdPUdQvgF4I
5qwRkPiYMs2J0jyVVdGcCiCC517byC0qcuHeUnzTdNwDJqvGAOWsPM/0BsV1Dtsa
93uxRITXsQCrQYPTQtjDl/v8a76l+Sf5HVWIIfiCpiRPIyeDjnrZZHrKI1a9QKOa
vGEKPzQbzikirHPfo6IFDpmENkreDm8dLs0xJUyR6Eep6RPK5DQUd6lwNHijerZE
UW475WgCf6vKkZfJZZkmqQZJ4y71meu51nQ09xf7WLnm9fp6ihiOdneWS87lrz3M
dA1tFoSidAPTzTUAlmUHJ4uC1fw80UB1PMPSrXkxkP4FZIop6/01bi14CyIPwbKK
LKH2jwlIDHsIUmIuTwoNq0TwYGKKdO49j/QZZSXM5xXRqjGTQV8kh5r86Dx+P9n9
IFYQc7NkFSTpBNUFNPrTjqcAQFPEvlOnLAovX6LUOfh8QAP17pbLUoxN3TELkZ2s
JqBx/8pt39OGKBGoY2cXVTqPmQcwAOC0Sp2mL6/S/ngSzAwP9bZpTfO0qOVa0I7Z
cScHp7DDiOhc6dksbVnO2ZfQabPuE3mb560ZFPZ2gW++mpXf0vQigXJgKxjj2YTJ
VjmGcJQ53L4LxisorlyiT16YVsRfa9UDulKoEZFlnMwA2n6d+mGeDJQe4WyFXQYG
VvzHuF+3ehuZGBEJPPYkeoUMJxilwJUaHi5OP6v4Vu2Ssd2iYci2MwuV102m8zV6
2+w7f6PY4C0mb5Vn4nscwiiHeN6lKvd3L7ne6wbD6tbqm3j1MOKXxWke5qWK2MrM
Zv2d0KB6njDQ7fY8rlslOnFk66fM6I4hwFtABxlCXpr6RUsfCr6m8V7wJGFyVSuN
IHdzbZi8LRrRnYTsYIgvpV62sEx1GZObrHVaBSjwxPGgjQStV8oRLKoEJaqzluPi
RM3Kh9hAuWRT6g+BWO8fryetCYtuow+HB6Ag3fBD2xffyo+OAe7SsL+UQW6yHuWs
Cjm3xHMC9pTyXiEfrCHM39M48HjatI1HT5S0B30ZYKtiAYhlZBEWJz/A6h9vA6bM
/FYvIMENMALe6iyTtpzNMvLvs/0vaJ8ICX8b8NWiYYfPswPzcl+pA7e/l/rIFQCC
RCDku7QHhSRmWkkwCyrXZMjdiWYRD3agbRxUUheZTICwgkr41LWZ5bTkqlWUNyDP
PSAq+a0vlkMmFEseEynKksJFMCrlAz/fiexERqZ/lKciHXz954qJPfJbaonrXn2s
aYLk3tfgOtyVEWpByruWsJ+gq5j1UsMOAbR71cmwrKsd57+8AI7YU4z15UigvKTC
EKd+smHmzphJn1VzJqeSNMZFYSPkSdz0hDzhjkJjMgNy4uXyaCjTg7wqYdCEn4pS
nPWC84fsNxDDfaUH/SRbngmJCdY/ImZ51Jhj0CteM4MkYlKfESQKQIDnbaOf7BGB
XnQk0rjw7wdDa5MUUjfR6+pOmpIqRwSG2lHVTPVijS0seh4sjK7esQhAWJx1BA8t
t3UYg39Ug4h3zUeRyT1B85asQ0WoUuasVOxuSNGsujxYLsWEXc0Dxay1H/3FmUsq
ws338SohoJFFrsdrtAYc+td5PbfJwgj7e0HK6pEzCweiZvLcoIETPlRRLfBPKP5b
DlSwkWzhPwLvJOHSq2KsFfj5by21Q0pH8/Q8+wNd/YflaiCXSEWGrq2cTeJorI93
KIc6h08A5KV0n2UVTMJ/B6OFUHcB6h9Lirm5bBXl6fki2IaGIb7Yc9M7ZM47xthR
8ASc9BMGHodzHBaRTKN8Tk/EHWDwRuwRrR5kPEZ8GV0Z1LhD2lSEq9Xribng6+21
dQwFmQqk1eHPKaUq80xpUDCpdFT2Whc2y+8oHuylgBZ7DQH0Qg4+HFCaUpgu9TTu
jQHxORu1l7fNbJxUKdvCn134yNkZeNjZangNYqfWwqXzI/fe01SzrEMfOSV8xfDa
U9FXnr3aGMrmCGqjrxnCPHSzAZPc3T1IJOM41gpUdLxPmbyFKAWDpP9wjij0MRYP
riG2u4wY8RDLZgLp+7lj/V44n4sbBrW3nevtcKwmbSwszBMvrxtAxLAnGHWSa4d4
buuxd/zKY8CCSbacybyBePgj98yDUqCUn59IjGeJ4Bm+uU7Ccken/SV0lPQUSDBL
9fVWG4Mh+F06MrV9QsBu+LvD67HwfO+QfT8QskQxkfmvBOum+ueg4dcX5Avgf6ql
SSHUZBjVPMBQPRa9wfUUvYgZyJr45yrTh7Flc8VVgfHxhb9m4jdYpuoyinw2Xvt/
WYNfue4Vg0jBZ7VflCcL1Wr4S33gz14zVFMeBosuTO0MVpu/UN5tsysY2yBrIAbr
iEfdrVadAS+/yFeXQ4i7qBVUynqCePCrOjDhXWBKB1EuNUTWiRFvUmYjIF7v1DXx
hTWgbvd44LTg1vRGTDX93uz1+kleo8X0CstDM/0x5EbC7LZu39BPh5nEhsAtSWoI
GuLV8kTs9e+AgL+Pec5uffyM61G1S+RwgDf3T31dVC4wvhO3rdqByNLKyURhCrIe
E/5vVNP13kEFV2FCk/HPLhpoa5cWugl7JnrfnsomiOjxGhIHi9UUHLbYl2mR2bpz
pCOY5/DyClyNtaISUIIJlV2vkzdPjVGem7bRmLWz+7Pj1tkMoMM9q8ADBbc5Fooo
jF51bg7cPJF6FCh7EDxuR7M/E0hFtVjDQE076KFwCu1UFqVCcT8ce/OdrcFwxf1g
eg2oKbTpDlxuWs0UZGJqWNN17/SZN8uxwSKNKZ16P0KcCZZsId1Dzk9WrOqaTQhV
cUrmiiD0qw08RE7mWkKns7WePQSFl5mYiXqz/Eq8Uv+ptLwK8r7YqbewUrYYRYOq
X44P21q+0ppRrcmwLwjomzXWVmOuO2JyauWkBY+NLhOv0zSBxfoVe8SSEoMC4bZE
y+2A4s7DTR9Rxb90h7RWWS9ADfQ0tyMlIUdvSSWN6kw7n0SQatWROGVPXkS0GSV6
ZpY3buIM8s7fG++l4ngeiO3fWNi6vt+VRCRAx6pQ2qkQESLxTuPmVg+B70IOWZw5
o7RpjrKbx613h3YX1TQU6ySVEdRwMUYgIh/svLAWfWqkAuz9jl+qiETaGd1F0nEq
5AMCqFZ+VxgqAqg9uA+QcWyXn/AuxCo46HcZWr27u3XepsPZ64i4r+lAXiKujmU7
Rxgn1+vdTacMab+rqD4D/cwHXrZXqpJdlbvbEzOXego+EUvyPLlGa2LCKG9pumXW
jQdBgaaA6srcXkl6HOMonI9WxBUqmCjz3IZ1zV1vwU9Vl7dL8/SOR+ibcKwrXw7H
EqeimNDiACUOsSxqERnlbE+YbZ8pmsXPsLqQv7MpiKKpQ8s3uS9E1hJiDCBDdQp2
fT8mEY6SEO/zlUCxZfZPaiqgXA0ww5aUbBgjNEfyopd4N7tHQBJwTt6dzQ03s8SA
VsGpg+1OG27pd1eCoPLCCszM4lEEIIRlDnwHdItyn0hWFF0ch4PPVsug0yaF4Rli
Vg958Bc0sM75x0uLAt6v6sTb7mr5d8L5vwXT3g8ojAlSBRbfD0F4xdVJv6Wl/rwi
Ee46pmWzoN3ZMps2ZWlTWQwuk2eKeWBSBwJti4HWvh9GOz4OFzoE2wzmF1NkHHhR
25XlTzR3SRnpN0ATl3FXDHu891TlHobQ68LOdGb2aoVUzoo97xghzXu0XNvHQ9fN
NPOARLPe+dJ9BwK/MhbbNeNi4WxLgMxudNySvnmVBiNCG6znvfjOc8Zh6CaLN8st
wN6/mrsonmuS5h9fp0gyf/v3dB6rMNGe/sFj7ZQWq3ptDYtGZ9NMQYYfAee2lx1x
Y4rExboovKTNodTKvxLWV+O3CqVX3alR3Tk/EmFWgbXVtP8YBozCQ+GlPU0zeRV2
0okw2kZtHfGZdXd2h0K7NHOF0AnCsiAObW1KM5FaXipUvu6NCy4czDuSMa6BLB2W
uOhBrsF6k6nksBsOjIpz5MYHcbjNMclOdBSCa+Y/P0qYybSNyGbLl62MOrFFrgHW
4ieD5XCZVvmqcWb69/YdEsB1PgbfFAS7dvOby3bBD6LMUZ2jXP1KINedaDkdVtqI
JcHio+zdWXLh2RKeoTBtdpxvEbmLiCeFlciKtsdltCNC8R5+0FXZfiJBiILOjLuW
Anue87LXPiQTu9T/bmUaCojw36dbeM5rjD6D3N+OZyD1XUmq8yHeyPDSy5EZXsy5
wxsRz/dtGDPppQv6YBkDud9DhSHQ5yAdIg0GLjQfZl7/u9yLEqgOy+ScVIUNIEx2
JgTEtsDU0AznP+iv7qtSK8NjZHn9EefVVS3blPykkYqZ8iUous/1RQpqLl2R78NX
6jDY+Mrgax0OK01mlXQBfBcusbkEVmG/o3pFsMI8oCiQHtqEYKdCljjNkuDJYn/e
bnbFqN360ps+9m2uwmH/zBNDhKGRs0xIJuIXLgTHPot+HJFHnCpG/yajCzWWSdIk
aUvikaPI6Uo54tTszi51keP7DEcqs7gd+DvGKhy72h2kYUyYflOZDW//HCNlHGhu
+RZTjAKRpUiyp3Tg1H7u41L2OjVWa74ME/+Pwv1JuNcYYPnLIOu0KXFoHz2gZ9IR
acPt4B8XNMdQQnov+OJgC2gyjwiyNslinF4EPIrXFdmEIZLOc18cpvXiaWIsL1FO
u3BmL8Csqbxk5SG7u3+RxMqGqcGw5CEAA+RdrHKfxgkpaCkK2p9BpVUKwMlt0UzO
BjSxcyPgKmH8f+7ZBKkFtXdvvplsoyZayicyWSDVX+XebbGlU2NXhLxCX8tsoJo4
qb6poyzxKhrhiBkp5oOTKIVTxWbzM2ZxTVyb3kEE13Wl7L7hoRje0EupSw1ViOjR
QhdsWBxfKPceGThyQ5V2fBs91ylVBVYA1rANXXWr29ChXKrvEWV5F38vxScJMLwv
pqM8wiwDexDexknlqzhCQjwdk4JY/Ud6vfOFwTI+A9dkkqAMhLagOrBVLLbXiR68
+tqmwO8Td4YbCBr98T5NeuIyc0Opk3ynqIQ8w5bW3FvWHMqx8uphfx4ZkVOdei8T
TdTsW0E/kQTtb52dI7T6VY5EQwh4rBd0nzjiChfFGibLxPBRPsC2rungTBQUxz+a
e7YhoGSiHtimAIUE+iw3D9ub1Qh/kD7J3d0YgwYqRIXSX55k2+HaW0ioWI2aAEqJ
c7x01Rd0TP/jayn/AKcQk1SBZOTdAU9Pd9vIg16ZVsNhRzEehzeY2tUo9goKHH2j
o14ytrEM+h+h62Po2ZbE0EndYJRA/TXqr9nJ2JR6+t1Qes7wpS47JlwMN3VhxBgY
EoX2iSQrTrRoVGGTdYNFx7aBkGjmX5/ZcntVeQW76XG5/5odbiqxzhVnubkmakx+
4ZqltTXIMGXS3j4jCp3p/sXvbihUw/+wplwCXY+nRILqvMCFHKoj1XB7zwm+vem2
Z1oQFvnKurJvdJa1Iwdmh3AVTikScvpYA/bTUtbVM6XRFYuGOyN+p6xYt97dYItQ
7oWuZJ8ky/sTyymn979lE2JHsEwbXf5QLXw4Jpy9oOF5ZjmPM7NfsqJi6W/HYh1b
8eKRcONsJOOSUiEShZ/Mq5wy9CWu6XE9FzbbcVxo+paNshRno2oRBWCa/lz816mz
wm/HIZYwgdzwmX2K2Z6irkePIhvDIHBa6Ig9E5PwBayUMAOL0659O/bdO7lO8AwW
ArdTy7AVT8o9I94ZXBHzFRQw5ctJawQ3I0gO5Fszy4us6jtxBra/+ZbujRyestwD
qteBpXuppFudaJ/KaLDn20TS8JlGGL+aZsQoi7AFPr3Bzi3BnUL/Yy5I7q+UOhZJ
tN0K8tjVosAjEZUTaISeW05uaXlEPBqGAOBIeYSyp7kmRxKQdBcuYDdKMROmhlJm
9JhcHP6OsNbxw+TdFatm5jDpfsikQCSyWjBX87rc1KLirR/HytzQJWbbanENeEJ0
eCrNBXBmfkRz+ESX5IhJMW7pexdp2/g9wLV2dp8HM15RrcpSLQTWrkAOyBJzHb3o
mB0x4GTaW7NQFcrH5KzAxnOwPLKyR9X9sXEXjxd3YSv/NtGmaEt7cusYVYm5iUkw
KebI0Zj4aASxST5yNr+O+E7oDkXHLXoy7710O5nNT1l9pBUecp7TeYlK/8y+gzTT
kjkucIQdKQQzv1JV4PD8n90QVS/78RBOEwygDkSoLTV2/3Q5NVF4w5n9poD9rmNj
AqolJxC7Z83j6PX2OebTxOm5EleFzRdUMOZCy0yLaGFyMqD7g5uGyovpyrpTY5FC
Da2mZRx+2Zt8orVDfFGOk1SWt0Uh0u1DGh30qOzUqGacD8iQY6z8CtvxZ5bjp6LJ
gbOF6YMSAOD9rfPPfQehxd38kzqu21oRwnGEUmvrIvtheC9y5la+odBvrZ0Y84z8
m1xE3OkqdcQUUK4VA52mnVd0ePA8FgPngLdKx6IsjVVxWKGuu3G5o/Y1p28fnF6T
rqnWdGm9v6RX0/pzmfnQ23o/25IE+yXyF3wUPIq0YxYYRwBCuW7wGPGyAQ8fWg/5
h2+iq4bIhHP70IvSNrcRpbgcC2jR/ey95VeDYwMe+PpTnFyEcfseiZ8SmqEGImtz
ZS69SStw3XIr3cqJhTf34Z5OYt5v1CBmXEK/xtd6ZwNxI8J65wuS6JBHJS7kOuj/
v/85zPZbPHQn6lF6UNCQyK7BnWl0KzpzzYPoRwc/SLTuIQAopzR1uJWOowJ7FKmY
5HBh5aLJAF0r83JZekrI6GtM/pKC7ryfWxTJEoLKKjHohcHXl93IlCDiMUq0Bk4c
R20MzAGaTdtEgFCXCnVhlhYOa0z4MNHI+GxZfx+UzvZ1F4mfpqMU1wme91UlaW6i
QVYicOfjgpoYRvbq8g185Owl4UMTT8ul0IRic77UkIr6e8PYhgq8Pa4EYVCiC3hX
iWnNLBYOWtr10tPTtBi3Krk2HdjVfCf3N5wR+6oWx1TfhnYWJnyF8TfNdUqg5yvt
ftgdwlfvE66lS7b9bgsVh62AAc2AKVtIPhCPZAtRKCeAtPEYr1hFAwiIrEjWql8K
W1e30Tk+io3eX5UF5XbIUCutceq3YsA6+/8/7JbLwqYEij8XGsNgeSxQ+U29ZIwn
KP7xInpKOLhxTbA+v7hVekvDNEfOoGjciIF3252aA+OdwHFBuXT7U/iMyLJBLpJG
o5McX3Ii1KT9CwhQiRA1uUZbX31muL5VYFdlsFHLQIXpldFAp/GUgmJCMpcFb21Q
u04SOYDj9JRMdiN6i3SvoicYvxldJBPVyPiI146ja8EqBZgtfRqYrFQ1zeU2TNXM
nqaQ7jM2+0zeln4BCXaZbuEqRwmtUkibqQdIRdcumUNCPwDQT5zOUXBymhvJ0C64
SNN9s4aC9CSsdVyVu67Fi8RV9jyyvKXYi5tbz6sZZWHy7ASPQoVlMlC2+scCqnak
8hgjPw33ALuttPCW4uxoCBhvVzfOdMFM+Xgrvr1XR8JWcssHR3B472lPf6T5CR/v
QkzwHwEtYBkz7QblPKpvwL2LIJ0e8aK0NaAGn/UHRjjGBsqm9YEL+To4lr5ta5BM
tC6K7+NMedE4co+/jc9TPUuO2+SZrPJonTsPbwi4lkwF0slx+BbSn/IGqRtNo5LF
Y4zo0u2/jcrliV7BjBmKn35fHKMDP1nsbQGoI3c+Nc4Q6nde0m4l+CR1m4w8wbtE
xixspjC4/ChK5aqnFLkWzGeuDJhsQh1vYkKhqy3dlZnsm1dbPTkhstC8AvGxCa0D
COwM1cidNkVLNgvki1U5NtYf0q9jkxEJiO3XKI9COEEL1BkI6+BPW+qHAtH6fAh1
XE3sX7Gc2Wk5b7NT/1xOEfi/88EOFZks2aqWDIFBNYN6/VMyGAqJEdzBgnmV45GF
TjM1ZjrnoTAU/EazQisu/kOrPsoufDY5+J5b92ckyLd17ZQo3kgrboS5JNuXSpNz
Va15spuztBVsDraQE9KBuSwql+oOc3utageUKg9psP0qjGZsAjdccFT/lFcUzSiO
cHK9Kt3yVB6/l9geAOcUKUCHvScBDmbNbzs2ziNY5jxDQEnTKztDL32f/MT38t0Z
2F/ZIdJX2emaW4pzBb7x2pawn1FeqZhUmXW1S0AjsuqKU4+Zuqr+v0GKARQcVYWn
zkf8OP0Jm415DD54SGfA3X8un3B62GKaoyCB9R6w7SCveuT6cFd/JWZ5orAHnZzc
B2d9yumXdrDXHH3k8Jxdn5jUPSTiBRBbzHLBhysJdbPc4moxdQ9sDQH6Jvg7Zb6C
oOWpcvYnkERHEEMWfCjbnC7ZqyZrCoyQmpo+INkFMc6qCYlGVMyvsQk0SgEVp3+B
p1RKanC2L6PFvDvjlWS7V5qwgv6gLRLd8QoGB9SNMLQh7ZI1bXHy7lBXGEY99Q/Y
l3kYQQ0tbjfYRvBFyfyn0+vfw1hA5vD0F4nyJg8GwOfZ9HLuGTosd07AMuHxmUo/
s0QPRcTeMn+qVyKC6hGDF6VMnW2rqAS+AsQdKpM0AvsV01Rh+tftEXd3DWUMpOi/
/R7KPP8qiikALQvF7BhqmHunfAxyCgMW6E/lXi0Uv3lhggjVDc4S/SLPwEoo+OMd
dCJCbYhAT1WXDIdyWgMUqAKmu74u0tpEq8G15fRJW/PjmOiyfLsfin1C5FYpHGV3
VZG18ZnultDxp3eCgkI1+l1rRTWZN3MDq5zS2H82L6O6oBvYpA/ElE/anLUq5XRx
yaGaQZJ1gaywCjoA+ptw9PP8ihV9IjcvPU0Zid/Mjrb05JNSyAzmDL+EWFfVhV4q
IENsEMHr93Ey8lQIjDgaygg3/Rf0ArvPzNylEZg3BMUeteNV5l3JTT10iNzJW0iu
vtIOq8BRzBB57vPoSLE/vy2N6NjE1CIa4JyZYA+ROIQcgAXMiPsE/xLMtE38iKin
exhg70qPDa7hxUO3bLhlyeJj25q9CtHt7iNQKzl/FDAVFhXemiT0qxfayHAztzhm
cfTdJ/NWWZt2tFrbuSVQPwwgjTDwS7EgDzFQsl74cSckaAOGZr9up2RsQeedBoot
DTGFK+UR1YHz6UojnQExJNPVAFWcrQQhb65sBauR7VshL5mzpGesSP2ozt6lD1id
z45fD720UMZqLvDFwD/LnON64i9P4tZuHd5ycJyPvZG4gSo72F3CnSzf7tVpmBU1
qQNz1adNpiHL8H4b3uGq60Ug4e9lS+FzugqCrAC4Ge8lAsCxCFhZRay9aWDhh5j4
xKF6B383GHfpsYBp2yg+QLpilDjReJJygi/CO+Ilcw73aNXJsuWF/HJbBsDZ55D+
RS6/pg2W4MHUjKnAUMRwWrEJzYHsz16n6y84woRO0afgu38jsMdPlvwbDfEEbybY
5uk7yOlRrCORsWyzyZR4D2aDRy1wUgG4ARHJRB5Z4U6DatTIH9i8bF7wF2RZxlni
2Hmti11saBfO8UO0YvQUg0V9RNzgsHSEWopxUZlhGy2SKq0sahQyIu4cuDwCX2uf
CzwnCJUASgEyPQJDigT7PSFaK+k6iKtqFUcz33C8M4mhcpuoLWCwNf7jnacSX/gq
lq/CJGdCyF9uJ71WtGEmDd25rieSJhfn702ZXNMVho4G4RKXGVkrk6wwdNirDo+b
+CCGXqJKR2NTriYmUFm1pvQWFsl3cx/t9AF2Lq6ChM8aogra/XPo5HiZoFTuz5MG
mKRmjuZUR4/ngX5CyZ4nTMxQ2RlpzxZiAc4rlO263Fbi4CMbrrz91rrKdwAqr/cY
fmP/LozGpp2rTofLlSeYnYTAR/rM9dzG6yFuhuXt9/XQSXP04Ma1Gn2dXlRFChXD
1jZ8TE4GVOpeK6LoBEMXp37ka39Sd6fDJf8n1PVf1mnTaJkMUTF+W5saXGpzu+Hm
fPH3iq+3gClps3KEOCWSudX4c62ETly+zHFS3VU2uyk9P/PEMhOIapd5ldMVhRt7
qHkvoRORhnluQkjQWpybt4ND9c+oJyz8x/Xkt958OIvWirUzCMqqf1ngcNwnEW3K
c7OWJ7tlECFbYrkv9Z6/TjXRIpy4MLEjWE6utydQ/j2fNa6OhwAftFAtuQQelCUw
ZNxJA8oRXNGavfJv7++QJ8o/gfq/DOqhub4ajESxZHG9JXVYnaW9tdvG0wt7JC1n
CmN8Vh0AjGmhSY8x9K78xxJ6KRrqOmzZokHfYKiiScmt7arTFHNL7nD2CNjAXN80
EAUqGBj5/7BYeN37ou1GdmFg4My3or2UFrHqUQafiuSHz5yUjIcYyRlvZV7MeN5x
w1Xm2odOVYOrmb6F/NhugA4tLuZHScwYsSmkZK1bkjF5KhhCQDGFI3fmiO+8Xc9P
DzI2CPJt9nKUHctRqpY90PaO/Y3iiPUIP5gQbxVIrB0eTL5RF/kXkMkMUrdRyi//
mVBwFRjbK5g7fvcRkUMG6NssfJdIUnLEC1mCV3aLVAJ2X3j8rTvdpxK2vGXcDRIS
HtlM/nKfqpeOai7kg7ScqpmqwrDwfqyvRrxpQHeiuzws4InGtJKGd8qfdfbgiOvQ
GzzUih7SWzRCZdJMkuT12fE1RugGswfcMXLFPTYUEVkMByWcLUGvTRQRZe9Fvg0I
cNkzmyOQ5coRrojFJEyGqmM/j62VFGtEggslKPpfwWA0egbOTLl9a0XYJVQ3ezJo
wcX4YmOu6PawUhLrZZzYYtsE1h92ApbjF8GfF4aNyQkJafbIEbVSynBajXqeRKtQ
GV3eiXx61vp7x4f/mpfEhBDlnztMSYGu0rNA3vlIP7ZYZFfPFRQoidk3qiRomTfb
aUX0PkJs86ZITrnJIcuUZ/yym+Ds7XRcfemA3n47gd+tI6piOMd9R95QBoQQIyQ+
Pudpf1SpMv50apAq/OH/dhfAJJbFjNo7iyCo74LXnsWH6ngF8yXI9YK+JrU+n4Uy
UgtNiP2Xhy4eoA7MJxs1Vz6h4poT7TdXqqv3zlvNVJVtfPsB/pY0a0hRBeccE7Ol
lJ8N0JYJnE3fQS4cSA2aEe6tK3bZPWH4Wt3141NPdgMboO4FDRYkruo0sa9Kz+JT
9J5Ze53hsKPIt0gfGAurijeKXettXxhjK/QjDYn0UrVMLAehZdQiWDa7deO4FpQe
QilFtqyfkDQ4W6AURNPTGMb0qyCOGNwooyDn+5vA6RZJmsBFdhbbCpE3TrRUdIdo
1GTvJDmKxAiBv6Qi/+dr/bbZJiyOgtb3g1cr//VUimSSjR2KscGI84AFVVYCb7ch
n8HpWSPHaAqLl4YJW8F4f5EdXtIJpStdzdaTi7em4jpKleWQDOVdE5x+1NqfWnN9
VdqZii11Hy0tPO5QrkVWpwjIe53Dd/0McNsiBVGxeyq4vc84824ywO0GtYjlxqvh
X0J+OpGoB6IEeg5xufC1+wcHIe8t31ui0m+BMt/pVcXGvp4tYH9Gb9kP+DM3Yh09
On1BMgOnzhXv4Hwsz/eevD5s0biyk/g6Y11H1Hsv3NPbb6J4WjE0v3MtkcjqPtlT
BRTfxV7sCO/WufxxwAd1w1F3veyRIiCHb0DzdHaT8V07dfUsoL0xgR5X0ZUCwcnb
B8jC6wR68OKP15455DNullnkMUEGcFnhMWq3QlVcDZZ6OpbWqrRxD21YseMKffpE
o2gDwnErxBz9ptKFWwGYb7ygbw0mqWZx+qIJ2fRosYLR1BIsJDZbEmz1MUkBuLha
YLgAQh1aTQ8yzzymHDkATS4KkYr14L3tWD0ksaoqKHdUWRJrMpvQehpf1DWsSyX7
DawS/FOG/+E8+vIaVXc6xdyqrHTzv8MZqlLr6vEtcNLY/FAimYLH0eXsOMC0tuiJ
IRcFdENFR+/4n1N7GrRSlU1TwBtrKQPvMElBrsQl2VykbNAjt79W0r2lVqoTtkbw
Tx0EV+Xs1mZoBk4erkeptL0RehZMZOI5EuUW9PPQMqG97UPNeKf7SzfrmvrgwPxY
jfgT2m5v7Qv6rXeLtPxQlkkFhFNKGuLhnFJnD0CfUoRSAVmupCcvN2at0GpMVv2y
BaOHkfFB+TjXBv35kn/i/rpQpQ4pbO84K3fBrG6oySVz2EeeA3D3DRdb3XyrZpqb
AoBrIeS4DPTxDNqFUnmOPEQRWNvdoCdlzFcfRh5U4DLDu32N/WnN5cCPZSKd4k0f
v7/AiQnW2lPZ20+EqKdYR8MYUEDGzJjyNOLiePEH+1PBej6DHa8ygBtaIlVfamF+
Q3FuMuFB0Scin2ERfHFwk7lXa4zzkPXZBiCq45EgxfK4qOoTGCUiuqOKQII+VKxN
vNKFCk9XLMfYP/wlj+C7p3hGGq/hSi7YJn8TqsjW0z4aoz1lLRd3Fv6WyDzJfxPR
JXaHVV2J7/WFW6xqo1qBiU9+sDHFlDZt9pzH1fGNWwW+kEDqsiICU8eh7NI+ngAR
LhEpg2usoIMowBAEh6aG8k6va9VFEbwf46sm+5OAPw73Yo7xTctNos1/7vzrxLNe
47Wt1anASEqSRG9aYo9ikXADbT6Gc+WrDe+5JvjuaVVdCZuC40WTaLeU4DWX9pRO
qXTGC7B+PKkAiYynl26MXAV4bTyQ70Ys127VxQdsmhDUhxqShImESrzcvjTTeesD
FMsv80iRxNEPRgjY3Nd0iWCsFWr22CJ7gWSif4nit+ekB3y8PIurfhyB9fT5xw5N
s8lICzRPDgiSgrdnAcF4XbnMjWCvVqs9pbxVAeyYMf/d55X8WFICxeOLZ0XJFVop
k3tJrZF0wtexUCamR/j+BbQI/BpambHYnHGQy4RXSQe12W/+EEZ0PkauNi5VBrfC
9QhZJVU03vYdLoFREHVBLbhx5GAvq7AOlOiOAfD5b8JTZ7b32nmrw1kxy47TJk/U
9xUrQrLA96b1QVkP/mJAXklHJCplsFYoV5La+CB9t6YJqU1uKxdXNG7ZvZpxXfmg
0RopmXgud9xodVIkl+4X8D57RCLpbxTiNrtLRAMYhiXdSA8mWXQGrYIy02lEalES
tC2wi4/lgKcQPWeoT+W7YYikSHdVM7xqT37DrQRcblqG4NFeBp25bF17xAEEe8vy
fYjjrsxo3OEIkkRVx1ASiFTL3mMBWLpUJwij42hN7SkQlHUKlImsIwzgx4UoHIcu
3zk6pgrBAnx67z6KNHdiOuiW+5H6/oDAEq+htLJVTmcyO4d1A2QUwZV1DsaocyLc
3FLPi1EpUuO0dNmHh6sGV/G4a22DaNSR4WYDDV24aenyWjwNFIvcwU9TEJj+4tjW
L1RPhK8uuK/6zdhpTIldl/9LPZmHC+Z8gw83HhSSD5KlYyDdCU07SnJ3sqrRIK96
//FO5DERDkk7pMd+3RhbBwkHMg1St/n1eL9pNBeM3oD0gPEXKgU9wfQyowN+GCIi
wMOufQ3jPXNwEaAISGszSotO87RCBd+aSar7zMKFqANoKkzvK9stGSqDdKUvL/Bt
BNaS8i+zNuCU6M+OiayyWivJc7TZm6XIKEUsSZG2oA0ZV+eOtebIz07IQg8NNEuX
Y+oSHQWfG6mm4j9j/4hIUqM0s8oFOkcdAtZDnE3qx4BpKylFyWlOSpVFDHxUPMAY
Wl/eWJKjPAavPJWcT14T8HhWs8nRobYLh8sko3Y6NT+yWAs6/21tM1/5d3Xdz2B2
5PFF2+V34qq3/41Kt5+rtw/32VDZhBQfVAsCCEXtAz/Q2U9SUIOelUnVhKQjA5Yp
M7LGnTdkOwANhB4VISqoL7k4oM/VX0+m/0Ngyk2bORE9Dcyid1nq+S4gujweNBx7
8noOwokiEHhZZCfVnHqyGSbBLi07rnQwmtwvcRpmHeFKwWLjFElAzQSAO2nR2l3g
wGFsOWPcVVGNFt39bG8jHBF7dOgwrf60TbX7OfT1SvHdqa5xpx42yTKOToY7i5kz
dmQi5nLF9DmdWvnb/m8wnlHl1b7rIvlegXN6aNbME4aEqbgeZDhh4jxMKPE1N0uf
xQDS8TNBZ5KEZ0JLRoOdwmpWYGdnTfWuQHqve59w9HlCEAN7G0QF95/J7LYQIXJb
8FOAtNB6Cphg82CVQzlY/7hNcGmInZ/UyhVdp0AqqYKbe50iyHg5qfEtm34XfcGv
5p1uI9FOcPM16bsPN/ge1kPCvO9uooBlhzU8TYxDmSfBl2AtuhH66JdgNbkexmv5
R7834kQTNvZjDDT/g7Rxll4ZJ8IKTovRPjJWzUljUoVUMDCZRpqqOJWrUzZJC8mu
4Q/qJZqf/i3/zCZMM0iLEMilMWOmGAcpFGmT+jZFpD5BvRiqG0Ia7gyXAweNvtll
eVcD8S8vJUTkOEvjAmn0cH2w7UQ8OaiMXnNAn1IULFtzGxaQlmxd7aFQTXf5eNW7
c19TQluVm9VD0fAPWZvooFdEyRx4HLKTVvrNJdjBu34+vphZumBNb20yUaC3JRni
BdRVu6ilfVs2O8paF5tEoww4O/xrziQ0uO8q6w2I3ZzIBkK8q7Ytn/+MGv1XuGnV
KAsuy+/ebkxA5iNiDcxKpyZadX7JI27kiBDcZe3BLIP/6aJl7ftA4o3iDKUHI/xb
ubpoYjynOoVNxBIW4whQ2TeJLnT0jkvA6RXlobpDWDrnKoGJS5z1tzDO8wBvDgLh
7/k/MiQGZJ0HJNVyOnZr2RNZrUwEDe98TGMOJg4urxZKekIFHeN+OBCRKQaB8tmt
DaOhn61rIJz6/EXE9jo2MRIJK5Y9S0ZK8qbpgajDI2O9sxyV3DSk7RKBgWB3aM9V
6KxMzTyxVrY4jahvaYeCMULEsiUOw2CYMjfpTGaRDHsdlK56eOzgBw+KqtaQnigL
dzC1J8wlgHdUaI8j+IeAmvBTY44w4xFr+OG0d0X6HBkU8mCBuGCHtcfUjmVJg2Ft
GhKiynaJFsadMc++qMq+XXwvA7LDQaUQeTdGU7w1+9b5nVh0b9fTrN8oCi94im+j
CiHzTJQ/ngo4FD7C1zMLckmuc0Ki3gX8eVTRsHObCwU6168uWT7p2NH1PsWvFGsF
PdH2kWdHZs/0TQbSzz4j/k7U/NuKD8mAsinI0SEshRa30L6OK4JBmTf8uO9B3/mX
3SblLqBKzMQqCzWzLhGuIKaMx5xiFHJdcgQJHJuIqtCduGF5pmfrzk3116rwvgDS
tyTAkEtrsu1gUaRJyaznQoA8upqg+Yfe/qav5xzCEDAlRQiuFVwNN8qylMcLG5dH
VkxjBm7wFTvv+bJTeHxc9199e2CymbDXMWDddwTsHUbukbII+Msg33S17ynfHqOC
Jzwpuy3R0RZ/Dtxf9MKHOlpdmN6n6RMU9Ct0WunjZZcDXurJuRXDQdJsgEOKR4Ub
YuSIADQMCIltxtwOtxzI8zj5CjVQyUE1PxWSeQaUbkctyqxmbFyr7QrI6FCcQ7CM
9xFp0vnl+sK8KcFMOQ6TaJKwME8dURm199VCtONutagg044R2N/RvwD2YRcQ6JSn
IeVvWp61d7oZt0orlRSKXk/dDg/MNZylqrfDbsxNrRDJvt8xsFrdtaBTp4PaGxzg
SB18u7kiCYMXmxNmgVTrcxs3Qy0I/89Vjhfjw9jX4Mw4zZZo6UTRSuEDM/CR1Bhm
rUjchoLP0WwOEZZcjKEsW2jfS5WFRZN/AD/HTORiMcsftI9tq/ClEL/Y48N6H6Tt
BX+PLbTzhDETR0yoEB2Nn5ay8avvcZSYQMWRarVqtLgphzJTFf6wMs8O3jzBydOc
3seyYGb4foIyt3VnEVJZAFTj6eUKSvKa1/V82ethE3eCji0E+vxM1zW0ipyv/6fC
wrdRqoYHfC7OWwfiJeZVRwkW1/EWfKmyGWqHf29zmzW9rhHstcQdGnAfUpBKOjv5
A1Ynw3wzxUSJzlKz5zANFOSiol4TpHaCWaVFlIrzuJYXQhp2vFWeT3vBjMpraTtB
F/+AVVr6S1370eIwaAreDriqSBdAgqwY1vAiCnDQ3eFexJRcf/7ouNQfgDzSXf/2
OUnxq894uEMR0fdbu5k+9HavLpl1VFOrKtV6nUfZFjDHjhhMylaXmqoWzzqpketb
LCQn9nfY+5sB9xP4MQuv1kjzwS5I+PTVBIUcxngoyI6DgmNmrRNRCDfgwUEyFd8t
iHg8yGWyvQtxf53uZTYv6LK+wzVmA8DjH2gfKLEsh0NHg9gLkml0O/a2A0OGbMKx
IREVfSATf+J+1llVKAwJneyFs2aWVKULEirqzi650AtQhxN55PmYO6naajEdhHUh
BFZy54SVkxzHn0Z/x9P9AcDrkWH+mdD8mWJF3yt632gR4sjzS04EGRbSZJpPX3/m
+tTVqB2P/g6qUy79W41Rce6+nE6YcOqMDL5VTKA4eEkCqvXaaVpSWd+u8qbDgoZD
W8UxrVhxWWoIL7RhEs6OtFIp0jPptC4XH7pvBzgWIlTYMd5lMctHwVFLAEP+WlPG
Q0WZ5Wi9KhFgcG13bbx9ni3DYdJDEDHenCpNs1QYJtEj9zZDVputTzmKuEonZAl9
SenIRfGd48RbSGVT2jmETBtzCPK70nfzn3ZXpYU4rbl25f+h562uwnyvhAjVsRnF
fsjxLt0L/+9a21A3ZaDLAmmJWVsllJEyMtrew0Yb/i+wyfOtnq0NWYVoJPSHRlaW
lbx8IbArzNRAqE0QpFEg/CXN7Y/fTs5/e8yh343hdzdmTOSp/sHOSz5hNDqGAS46
J2D503G+Mn0B+1Yf8g6aOUJD4GNuXAgk3Jp+boViDksgkj5xgpEoTZP66+v/fpwU
ovpkm8oUr1gYU6GbJruUddcOQ2HFG+z88urrSctdedT50zC3hfm11JVhBSRgjuv9
eXiEEKB2IjTzq1Gkhd2frReC1/XaE91VDWhUOzJ+NYP0aA1qC+e6frP2g/7yBZ6a
srUOmrvXXGZUgBga3iZJBhR+KLTyVZdxg5r5rmcmwQR9SGsndcUbXGOLxUS5ksZx
ci6flzVjGzXWEC9Q/1D08qMAwTBZbztJH5XWjDoZYRz3Ne6Y0ASDxOCwcWQNFdVk
8v9tRz27PmjaMt/2lcR0Ke8L+W/kBq0s948zMZMcgpKRs4InRtEm8+N/0T9Ty6rM
J4Vl+Kc+kQPD+iU4p1/bbUrLyHzJ75POBEu4gw7rKTrTGD8z7Mopot1VhM57TkEO
Lrjc1fzCrMa0fJrGMsrAONHAL3bafLOh5hll/MLXQWlNLX2regNpoZvcZjm02GXU
HIcgmoTNSw9+yju46dVM6DrRJgrY2lsZ7q6xCKq0W83lbMbpY+myuC/DN8hkKyxD
8JGc/qy8hnjIpizOjVZRsaSmUrzxGQKSJmYuvgw07DvDXIbvpSZy8elOagsbn7i1
+zHR2yRtMO3/NPtbQ7vII9jq9H8u8iZqjByT43LAOp/vT9kk5wBD18WpTO0Iq9Xb
FlVWcb1XUi0b7kKNCbWijDL4nwEbmamuoU2OOOTY1vwHo3Yaff/RA758c13lSnyS
86v17ok3V1TVwl4adj8x5ap/kNTCTp0Nj2Ixb5VJAVPkET22St9zS0crLJtcxRQc
E/NysgqU9syZIUiDrqgu2b9Dof9fRX8fxtbYRwCKd1l42KfVuRgu0fTDxsMW0FnH
7RafTvQUQEcU0VrT2fj7toz/ty3y+fa/rI/kW/CAgW/ZvwvkCCk09G12QF9Z4t3L
CDgbZPT7t5jjgTvm9ak/Q8aVatNUBe0JFzrQDxOmzlpfGRbP0CZYU5IaqlPJyQ7E
L/xqRyuZycVvtu53cxceh5sFHvTK0t4jD+cJWu1KPON+U76lqBkXxFkMT2Cv0IKL
a1KAglZzU3JXxQU826SyNHVat4aFPWiHmD0n7Q5JNiAqSoVAYYRCGgvkLXcmJl6A
fXSGQVeiBYy31Y9gYAKqDVd5N8Ku3Nim7NhBffO23CCHCRsXGgJBi6tw7c/qI0Xa
NQEQgigy8PK2TmridU4NMYbzKRtWHuuyrIGJl2FkbjynHPHCQHY559HTwc0sBAI9
hx5gdgnWvMVsK/coXJahGfquy1lML4Yae4NA/7gsh2LsmXrDo2TD6TXVMte+hUn6
WR4+1M65qTVZ2AeS4o5R7mjTDkROWOYscpLvzVS2H02Ey7Ke8rd92lxkIrURJDZ9
/wgBf4zqkF7bUk77I49a3lOIKYqbdjRSX0UuWgDMOgjT23u+LOdNrF9USMgrj5OB
UDUclWyPJ+bkvMpy7I1v6L3j54wKpJpq5W0rA8adKq/IKk0yY7+XlDgLpyN6FcgW
hZ4XpNe43y7XgOeu8889ENHYgX/G+Ax4hc0BzdVkxW3WiRj9I/t0R20fIUWINwXw
YKR/UpYrfyR6byWuu4Eg+oatbzuYRWtmXN/Yf/T8UjxNqMP3x1JdBnnOfiK0WsYR
vscIB5RBaetmUdisXb7zGBIwN6Np0NUf8jZG9g7Bw2ojNzhOVquAVFw1KV1ngU6Q
DI5xZ4yXZq56dqv7QlcjP6EmXk5U8Pysi368pBNayIcZH590sT8koZtfkirka+8T
ydBqrRiK4B1uBFRPMgUr4VN+FYmd64Y4ON11Di+DChK824r+BY+9pfQ69g6FvdI8
JVQU6nhFwvZgulFD1OfzTZRrJg+gDcUpKZqZzadGwd3RiQSydVb84H0bynGO7PEH
mLUoWVqBqko/iI1vcsL0MtZawn9tYEWZLxychwBA4pHVQTsVuDfomKGT5xxipkVY
CWMjFVhVPIYen8XHl5cHZdVF4IzHfy3mkZpv2Ps8UWXbmdobF0bHXDtxWxnxiCX9
/Xa+4GuTWG5sMrG/fDrZEMSerzYMxX4kT4iVypzPdg7IIuuNDT2wIEzHzhSnAYKp
8gNT45HSjWVz1+l66OuWr/HfYZIuGN50jbNTjJENiDHjXjXPtkdrKxrGuZQQ39HV
RNBqNMBAFJBkjOt/sddqRUuIjiyGOAGPHh06/QFKEQlbDQQ3k05VXkhMn5Df7o88
parZJ1iMgCBhBVv51Mlxa/AmFt1SCWEF6MEc0+PMQfd8EPun0pNPKQvT1p65Aph7
zkeo5kVHIdU/D/QQIPULwDWOGczvMa2omen8U4VV4D7SI/sdVkncAfoN/8FAm52j
3YPTmIIM40VxVd42jdw1oWtk1fUGnTpA9Hihv5pJNbQASVc0A2racr3PGDDLjRK6
7qpUDCmimWg68OkawPEk3p7mCV72yb7sSlqCuw0IjSt1Tgm1BXyjqRsPn+BNVmsQ
lPP8uAdqRYcpOr2tI+h33mprlY1mnzWhh8oK2s3T8sPpSijwOvr0e8DtXgjBK4Vy
VEM1mV4SH0hUOJjI1iEVSe+ayw2NkGrb29GMdWQLUG1plTGHSUtgttVW9aKwcQPV
mqwW1tv+m1VI9Gkd6pl2dD5iKI8qu19gVOEpXTVscFTvPH0P4U4t7+qBXve6pa5u
Gy/xT1+Z+pzN2TMtuGbH5R3pUbzm2Z7ga029jOHFMITOTpox+3XlthXIOMyn7IMK
ilT+URrSx/ealKpjc5677G/z5rPr5fi9xeU1PTtJhH01Bw7zxY0o9PIp9GbPq310
vY1FWIr7tHl3Ukv/fYTe0nfH8PptWLObxhru4rjEkP0fkb9bzY+Q4SJufVmoyc5B
T9WSiQriRnC1XRSsYAMCZ9SuuFHD4NKbEkKo5eEHg09WtK+0B3rqSelhpTQ2xMYT
6zIUNRXJ95quqwuzGph6sIWSsVKfcwgK7ZSBZRsYdvrZncQGOfX+cW0zrdVzYz/N
JLv4GCU55rFq8kOWgihb+IVJ2xvO+uQAzG99Is0PODiEB9EPAj06IZkBcbMavYS2
0V1lKkh6K7IArmqEx9nkmxNg74KNafhtwjlL7uey3EJLihjzWBDLWGvuYnyxpXvc
Tnq6xkEgfd87WSTLbE535EDNCHpi39bUgknhFBQkANXSA0fpWzUyoR/cdDDpzcDn
lwabwZutOFc667RfSF6Ce0cG7jslisxcIG7PJBmSYf0g5AgSzxvuQyAqGF0IcV2/
SLhW0vA9VrXcyYkT8mFC2Sit3jwbh7+cm6wLr9/DGcY59hGRuxl0Q99jgeAHIk8s
3jRH6YRRHMOLZa6t3/4S8JfMyDxTjyC74PLI5HW1OPcWeHcTtucJOmNtHg56/koE
2EjCPw24kC/TwwCFQIRcq7fHJVRjkTTrkBjnF2c4VjXMds7K6Rdb9rOYN1TKUaJI
dLfrPYQjtTUAin3EqSKckm6dVqB1zfNvnLzKddR/XWQLe3DcJNY9bx9VUw81yN09
djz7Oyg/z0DCaw57E3nwR1Dme/cfv+xPB7q9Eseo77U1BKg4d6NP4Ih6cGNHWReh
8Lt6/kmMhKs4YPH0EeuUGOBRc+y6+XhsriM1dRmFKTsE/brhfoHHXbil8vfMaAFP
Ntxm9XOAcnxw0A4KDwt7c2vxDLB8jsGBCckxc22tSEwYmy/i7t9lvalmM3sLmWYe
Z/hZNz/I0kH+8sfHMQf7Sn+g7lTDYX7dWXM/UYRQWCNRMCuXflYCPCXXMQA0a3Mb
EnYMkIuAXw5OUxbCLn7ikg98hBQvAL08dBz6jCC2JWwGju7lO/1yTfR0QejhguTE
bZvpF04GTu8VRKbZZyN8xd9Ed+yUDuE6EHNN4BmSEgiXJSWCbD/hqbDn9RZsGmq8
a3+se0WvsLq+8Q6QIcdzkV9mr4Da8OmVTavN2LGobPIrsgUrlvlFpRdBTJaCalO2
Gx0/2OxcRpf5syzXsf47RX/E5+XJFv+wZYUjLD74KeMW86rbmMQZPjpGZ4wUctGJ
FrTpn8iYkbK6cpyoTQBF54oLNnt+8D99gj/+TMPL+T3na5zy56+y+WSZuMxESZsg
/DBAcI0bOOzQcjthsIG6DSD0BcFqq5rEPesvl35I8l9q4ODdFZZGFzzDIqzPUOIG
z1dFMeFE9syFTCe5ZRTNHq1E0Gny+uZKDS9gIzSDU9f4MxJaqT05MboPbt19BlCr
I6Gqpyc9652AFP8BXaTD2NjvqyKcMqSNCWx218s1VHP5Ive8VbqC6r/Ph+LuDHQf
v21MncwweN7S87ekHGlKzuJHHwk90K3KXeCgveb6xJNMREK2hFkryJMAilSzbGjy
vlE0arre+0QTa3f+LkLWegHYg57kg3ReyIfaO7kMC0cea4+QEn3ig45SCoDrJSx8
RgZfacWjN0DajVx1wHzQGGoPMskCKnh8Ytd2wztToPl6pQeXCwZuRzmtogwJgXJf
E03UWwonYW5NHMLpeIj8wwJeUGJ7r5bmEKvgxNKgCUZVX//WAWRyNyaDjJFOXW32
dq0UKMa6Y3k5EII+2xmoX6yOUD49BnYk3Q0zk9ZtC+rAGoUW6+grKsbW0kVsVIRa
4IYW1E5P9Ak4rgiwCqm/U/iuuHK98STOh81nYrh522SlG1t77NE1Muyogd3kttyj
9QK7965uzFlXe3QhbbI5E/s8DdjAIksrXN0XQnTI7P02v38dV//2l3/rMWgLSjxp
v3x03M0djOu1VwczW3w5EygZi7vLJJ6lIEz7+wGfpTc17dWfyVznHsA7BaTdE5t9
ZmpjpqhnMv5+U+9nbfB94jyHm4kZ25lI8j434ybBzAqC2/VzKddwvQQl1enqYInW
Kz6h/Gf90gYwEn26DNcgtXJ/XpXrvC9OWTGWvqDZftJOgiSgNUU1aG/1hUmRMilz
KZWt2s4y9d2yt8JvKLxpUv8Yb82mq9O4Y1bG50SM4Zv9aGTvPUcUhD3OKWQVP2TG
nWOftvdRUgtVg8RbhKR/u6LOMTFE1c/Jwk7j2WoQ9m0eecmrUcjQtnzr/Op9LO+l
gUtN7KPAovZmNelDG5dy7JeO/7tETX+akHsujhLXdz697Gi8hAtNyArGK9GslA+0
Guv6CySE7DzXPTHjb3daCrOBKzeds4xh43LQ82mILl7irLsrx3+Z7li5efSP68zh
e4ELZxWob6L2wTG+hVB0YFj3ItlLiQ2HZJ6Kc5/qxvQuW78w6GEw+MmrMtgrdN2Q
Z36IqSt90ymI6zUrjL8zmVe73cVgEN43ZK7otF3N0EmlI1ZH4Y3ME5rDe800O8sX
8wrJxDLMvZ41KH/t6nJNpJBnV0yGQMwSOZX1fc+rskLvH/i/2KNL/N6mdkcaiTgW
4fs96RMHgTzgCwF3UDuLFDv307zLOaKZSkY0DG7Yjp251a/FF1UbDS2Dq76fZjV3
RzhhI//wa58Su17RkeIE/A/z3Ps/GGfsOFV4VIOZy6qIYMRVlAcyZN9q01Q85H2W
v9kuDgMlBUHTj2Uodk0eO6ODAtZxasuBmp3rERvlGNGAhW1BXaQ7HKUyHheGk0Hf
YiU7GMTZXJBDWTdnbIdwIw3ozwkWFObapy82AGoSnij2Fz5cO/k/PjnWosZ1bLgK
TWRqNnrJueZaIxzqny5gUWIPgoEfMbYSRaffpGZhiwkYhs+fvr5Crs9Q8rgcO/mm
sevMgzdLdB3kOJ0+Cr/szXYkPegF/rfRzpHENUSwn2lRm48O741+4NtMaFEiRjpY
KchuETal2uXwNMbSw1tq082EgEOs7DG075Jr5VCTd5cQiu6EbOt90PCVEuAqgPvr
7P/tCfvYGAgqMFGr/T3ToisRJWb1M5qEIXoBH2sySVDCyo8mkBZta8LkQ/wk44Ix
JjmggYdzZsbPWZkcb1WcQn028uXMlfkFc9+RlSpR0xsGgSJ58kWjB6OrZ0URDKSU
fuEZ7pUVHjTErU2CBKr5uJVUlY5tacUI//76CW4UL5Y7R/T+alF7XXsMWF5hE/Us
d7jPp6m4j8FYEqY6lQPjXDy/mvu9X6QCGf8FjbSmUdK5QKHVfxTnE+DQ5al24eiO
XH3omebSnOkdhsZubOjEkNYM8hGyOS091Ur4jTgfFafFk6oRkTHcZMi+29Yd47dV
sV9lmTVsAeOkAY4Vk4yEzrXu4miPGW9asQL2Y2pz7KLQLtLGvXW2f+6CvFk2PTxg
oBxbSUGRuhwm6xUY1qfbEcRJO/8zKFx/HChW2RFDu+K5NObLCmnJD/e5Bm+xP5Lo
NFxTUZUi+at0Q2ms92yQMZoWbqUBUMjq1GfNhxlkkO1G8bVJg4Lrjf9cIQNheAZV
FOSBnbbnanryWjVSqkWPUG/QH6Or9l4mZeEiTIH0XX59O9KY1gVjVxXo0QmeIUqe
wFeGDkvXtaAMMo7vFxPw5gJMK9BkFvojkALdxRZFEXcuWALIKZFEIKUuJ/wIWJvf
HdHjsRfEK98GrQICnNErRjyUurxu2W5HtSLme2m2YabxU8YHHE+5u3NgcJ5fvTIM
c4kdoEojVlsLPS1cTfc0WCdcvv1/9OVR16AOEwhuGTymYBZlchV1bbxQhNQfHVxg
tR+j+MgeaOVa4w+blrvX8KijUH4jzrZGQwT1OT30qL1uMP52AeL8hlLkNbiYZhr4
r+PKNnOzjXw+C4SIsg6LD63neYjozVOwpBh0c1XtBCCFuRrELyY3C9cLCxBJaCXu
sJFjem13aDIJ6HwOi6+bVbcJlJDASLMA5QbjaUA6Cl0aVErkB4bSmEWTaEeoKssw
jUun9si17XHquFLUrrhNcJUiuyOFQQNkY1yFZI8S+y0mPvSSwQ/JtIRVQ6o3pwcE
LUQUf55jSxhO2ZZR6gjKsU4pu9gzt6YgYdDCiqxa7q5yF1si7HZsjNknDo9Zw8Ej
Eos2LOgQPg1hHRmh9Ex1B6YEirYFDDV83P+ZPsVukuiIu1mI1Bgz/Ci44sOSqEM0
5gNujLgSBGsnhduNy7CyJ/QXq7hXUbVctsWlx54boRKn1m6jYbIML1TLIruNzaxC
kqH7vKkQmJzLrsS/sLP+wyNd6TojWMeWMKy2QH2NM6o1HQaTp/lTqTTD9g8IcSlT
zQLGg9HhwuO/cT0zF0kfJNF+8L2igR66s47Xi9g7zPCtTiZfuNxY5CFlJy4NH13t
NvudpHgMrqeFLKBJMe2DXm3rpLhqGWuxl7flvQO+5UGQd2zBulo3xCdnzWWwI8Gp
LRCerk4vlWg+1GWESRXO5Op6aT+VC/Qi6ODui9a3OUJpwnzMixEjEL/gc8YA2J9g
bu/r4KFHIWENQRZPI/mldY6GM0Z6pxxHAhJg1Buo6s4SXtGUzoQEAWYCJWUXl//I
G+BKnJTDxOiZDULWJg2tXdqmQksaITJtA+QkCnVrxPOEMAraoCqvdkXNMNJ0rJr4
2Kfo/4UqvVHIPUY6spdDaQsM1QG9enh2znttlNXjj8B+9dykB6kpdSAoDAkAcMT0
ycvYGsYVkNoleJgONMxawctfKRWijoqTFVReplZ/8fYDTRrZ1R9YZCJQQPE7z6qn
gVfqIdrmOjOEGa4HGrytKAnQA7q5Tfe89HhLNN/6/Bt0cQ3sSXm3YdK9c/Ncsb44
JsYbBp/b1B4VzyvHxeJhFbQXr9abtyOM+O/1mzDlp/MWMDhdalrZVhc6Od0oCsHY
qFpYXBH3cfm6EqEfYE7ivXsj1B+l+sTMSwlIuGYZFqLDXlLlCk0/XoCwp0166DAo
c42EM5LYwPcr26t9Kk54gmOcqYb2oFsXdv4eheiujIfp72ortEAuIHhBSWQVVJSV
V0obraAyJgYYj7Mzuv4U0h9Q7loYD6lEuxJdJEye/P/bZhz2vvmzOTHDAgLXF24W
VDde8qDF6mM23DwTsYaHQwCw6mevaux/jc1kjKoSoycGse9OtCGO3KmViIIVw2Ge
JJGzRdW9U8kGiFGXe45opC6nBIu4zI7S/eWeqSrgvNIu/pqSR4eIOdiEwTK7793B
chapgnSmeX6MWg9GvLZEIjOezYBaKYPEK02xbKPnjJJTu5EdhVyGRWcnqYHbPG1R
oM+KYEay9NrM9aho+1i2EOZD08xWRhBvdEkFi4uWuQT9QuBYxXfYjezaSpqcOosi
Jbli8nkkW/2otonvrlsetSsMu3cXQTedKNEngZZB2DKIuq5htphJ0JnYJ727Twsa
ySbBUjXtId/P8dFnARqBEH4x8QigPWgDFt/Zni4li/Y6Yr41OyFbGMWyQkplJicw
MnEEXvRXCgCA8xj3R11mzbW+zv2QhTSoOjm+ePJQKZZvWFGhN+rQhQZHSAhlGegy
W36qpx5Qq1uZ1pTLjE1mYge88qDB+C7ZHG25oVdo6s/GWawr2VB6M+siql/7uDiM
Mh1tlAKNcq50wlYNJGVY5LAIVEFndbixJ8ytEjBJSeA8RaFmgaZf4lW69HNvklv+
gHskXthiHVCDQ7nPiodv1D5bAgqCtXfrQXqmC46vOINmXnM6114CYYSE7TYE4yxV
gyy9o4x6cwcJDPjykCRhfOV4bL4sNtGDIc2sty0I0jSu886QAYarO+vnYyIXsxuG
Lli6dFywjtIV8KDeXWasn0spbdqOvrv7gCQLYotKs17okaXvXYtgJQmTBvdWB2tn
lHJ7IHyuLvhQLo54i8ugqMrYAn0ab+DWd2LSxz6/LyPTdOK4bWhjejWNC2p5xNf6
Mddh9SUM2DnVYWX38ETt+TU6vPqyDaXx70j5EkkYR+J3cvzo1yYdewo/oV7zLXlt
NjzFGh611M9JwXkFwfTUih2NUSRXR0y0PfIGi8VsqAgWolu20U91/b5qrlM2jtMi
+QVchZoHTR4VmTwdOa9zxT6OFBvMVUTvboI/CJMC2ThBFTBnYOr1LDIVMhtr1qtH
OalMuI0ufcZjg6eCYJNPyYfzfPRGzE06B+gLLcp+DNvrwIFgxKej+EUdrtt4Q0pO
E8RukE+EuTx1gh/kGoCcBcBV7zBiwI7ue1qV3K0XoK+canJBk/YdoQCKvBeJpH9O
oq3Hy53veQsyREgGeoS3ldBbRmjWOw+Fzr7ZkMDCCyCOuTI8Fq5Ar8b+HlpzLJzi
+hCxdoueCBFk4GsT6s7/rRu0tKHaCq7/R6atUcfnPPwiYGQDEvnjgIQVWCgl0ytS
tMKLnRDP3hviKYX5kyxHjdxl5OUWt9pLFst0RTu/oJDtBcOC47QARBhq/LvOhJfD
SWFCV10ygPleH0oKq9zETr6Y5YhioxZPpiujms/nYyYIXVx0csHZ3tcaNifgKjyq
RDSbXq2OpEm051bbT20XB0SQVGnPpoU+ln/ue1Q6d5Oz5KhhNJUfel4n4kN/SVFD
0EpfTTQR0WyfufYU2HmRVe2ib599zC23MK3Ii16cjrQkrjskxFjq3NHX2idtIt6j
KdzDiQhL/kXi0wlywzsYSCyx2mX7IZPTaaHxL6/HQ9I1jzb+oIELkUWZFYqQ6ooh
xBHax9Ap++I+eKFDa1zgAI+pk82XmJKqbCtUIGcPdRfwqvgLGSekpdknvDHcJQC/
AwaQDQ+m+25jv6Vntp61XxZf9/6QcEUocJle9RAXi2rMht5XPpt2/oqw//UJQIDO
iVlOK5cB5lfrB19uS+0YhBuzM7xC6lhSJ0PfzTqz2eQPF3/Gk4w5A/oXqIJZBOgt
D00/6x6sfMi/R06ZvuUM1GSWIK65vGZ+1ewfmyn8BN4Dxc7bg7nGiPB3nj6OUfm5
C2t25RgHmV75l53E078a83va2qHgRkb99ARaXRmgZVnAvFTIpnfdZqFDtCxiyzzG
xYovWSk50V9HY9dnaWXuhSC2XRwzlD8fvkYYD4HjfHi3ug9llyD/eQ17RRYss8iY
11/Nl159XAYDilVT4nJbvYHfy3AUXirZmT7cHaXCr+bFAGhO2DGBiUyVvhGF9Pxr
Mfx9l7rQzFPGUNcQ7sV21nGT/TIjT8tjAQt5cKgOH/ErByUSTSJpRyhPuY8EFuGD
oUFZZo/+DNFq7LZChqyBWdqSNTna7T7cNFaJDlZAK7/xn6f+5oLRHHALtcehCX7a
E2aFUPsUIomCuTjJxL9xp/l3VU7qo4Ul7EIKBawiac44vvckmwGofVQKVXmiksCR
LibMSruDTdQlcepQg2F7geqbdnORiwWnu2PiWcykBfE2TpimcYIZ1TVzR3ZBw3UO
UDSEk9meKn9wTwDaBmBHtuHyPioKpYsnBsFnWuWBJJQ6PSwupS8n/47WekCIIJNj
QjcXPd1WCjw08wS1AzlztwtgdCIxLIBlqS43wAIAAxNxWSDDOgEPMYSXpsQOunuo
mCRTy+w0h2QEkwan9g1Y6lyTp0qdQ4jLhZ24Jl7W65/eYrs11HFPIfJpKYoA/GeF
HCB2hdjpsPHiPjcHU5LGYsO+C6Ef3H6U8xlDEQSTKk9kpnsWJdq5XC+HbDfVpRdq
+inGJ4850moOy4sRhT2IC6Vw6JPn3qO4qqpuY2mh7P6p7IGP6ZlzP7u6jTMM/rjC
X1kYDnmaP897ADv/u8fI1NE5WKURZ2WH0sOl8PIP+PI6QFX8XyMgHPqed3zWkdv7
QFSKOyaP34P9TtY3g4WKfVqCs/FUbbdk2ik3g3ID7o1ZqWMNDy7nJCoRH8bhrBoI
7hwYr5n/B74ziaMsbfzWvCbnZr8kHBJ1lt6bpNpXETPk8br82vuPJCUacOpR0xKH
f319Knu7GceXgTLBwZ8UZtn13Mn23IiZl+BwgrhMuHKaWybR2wgj5b14tyMVFbDh
fnhjEW+Uj8fNR9eE8WMSYWp1tEryf8eeNUV4HI2rb6eTw14ZNZv7QxgLjHohu6xK
pHbCrbIydJpeU9eZhRJj88GsoMRMokdylM/fumxvfgk5/Am74OYXbf+g5/xkBIBL
hEJf6YTzl6ag6M10skkkWBC3KZqkZsQ5RLBtBRmnpiBmEeXB6Dzs2aTDcGkmEjqB
mmqvPm5mbjG4uOaho5udUzkOoZeWvXLz+pvCZbxGqmesK0jA/Eh5fweXBNXrPeTT
QI7+AukUApK4u/JTXGyb9f+jpoxbn45f42yACWPHwVmURSr0U2JrtFxRCVlOKCtJ
TOHIFmdLWUZ7/tk87ACcKmkvef6CguLfoSC/AHWQm7fJF1jB/f1Z8fYXqiao6f5u
7PvOnY9n08OP2gyBBBm+x5gjUCzSNcFFQdBSqo7KOGkJ0rjHaNAyVKc7rhfhjg97
Fvmm5yZrov9932nQDLWLkOL3RuZd6Z8gJN50Z4k7V6Zz9mjQ5iyD3aq3l+gdIQpy
xP8isB/mWNNjNKB0aPXDPaghcVd11WRWsnhB+fX0cUp1k6iyih8Lm/16OTGa3VVZ
fq6FANfaBsnFjy2c9XaXKHunjfmNR/fLFTDUyMHDKj22WJhwHe0VhVJnPamHJYJy
cT1JiC83JZ80k8E9WKUSSY4WXf8GkjD0S/Wc5rDcx9/Ks5FVoafFzt5R2u+k9Srd
0SoKGzXdxgKyghnaTJWuctpHRBGkMxZSYlInczkXwTaEdpsPUU5AMFK1caicp4JH
kHvPKgCbeGK2BeHza2n//YZve7HcBoZDjmqB0+6I0rajRA9oVHJHtBvUz/CYoUfo
DW7Rn7qXvkKuRHDpU4zNjvc6m38AfPiWNywdt48CVJhNyWwu9Xce/1aBP0Px+zVT
Fj3GG/1OkdYsO/B/rYlz59/SYXg6wD0rDLD52mpfvcG4UA1+KlJggjVkI/hrO/Ny
FXu9zkS2foDzfokTJsHivZi/Lk9ntQIJyV9cZcnAObec5bd2ie3D+cYV7okEsMYW
pfjzfWRqoT4YtoCsFcvqhq7o43LEEFm3UHxLZ5x/6keMBJju8Tr5Y1XxZT+JpIlE
3msEHALMOkiuopyYV3UmPl4bPQJB6JriO2h/0555XjX/iCyySqFb6F+vBeOxmjNc
rn3aKYs+p5GbO2316NT7nylusRAh7K+pvJ9SOaYKDW+eoD5QXE2z+VjjB5UnbhUx
DrFYlVGykbeDhmOmMi0ymZ5e3Ir8lnMa0eM5Y6wGbfGrFyrqrNmOqTd+j0OH64kf
zU4FvVZDGn6k2zULzoTCRLi8Ms4hgGZy/Wq7TwgYzIriHE47Lg55uS3Lu7IoocOm
r2XNzMCF1xxYXYNgKsXVBPLElhCIk5ZS3nxjai9kuM24GfKCs3nNl+HvAMy1iOXq
3xrB4mIRk02dbF121JvUY7+OcxPDX2b/iHbhMr5eTZH1nMqeX9rQUYigVd6kc9Ut
Hzp9whwm4GFXqmDIMOJIfSTesZW2mQcBdoWkV0zz4EZPsHcUqtMki2aPxC89kjlX
ITQWBduYanxzyMbGA75aDpXki5bsHEOSPXrbptL5W83XJd2o/V9jAtkt4aaKqGrG
vkEvDzNSQT8H1BW2VRrxDjReP2Pc78E6CHeu6d9u3lDSNdSihn3NX41lxPqijr1V
0WQAY94U6CPKAn4OnYnhq2GeBShxGRZ26f1FmyecZEDlBoSLdcLvF9OwG/t8+PzH
3ZhJh5nsLx4ZK+9sWUHE1ooIoGPT5xWYNQ9v74qNXWZ/t+PB0aoSzRVaDtxy6aRz
xA3iYIeA8m1N1InwIdogN0UGM19/2iNv5Dd/CS6x53sHSbrNmD654s5JGODtOthM
a+yI2KJLauQtxFZJ7lnqCYTECVX5ALF1ZfDnu+32FufMePmjUSfA471uje3LVcCj
tE6G4zibtfWc65asqLyD0n2VLF8fQoVtbBjGJ+Z/25y5p0NCNH1G3ZMZgFDH9RXc
GoacSOp6tSeL4X9qSJbAQaxl44YZ2ukWLqc7StVuHcSO+EHJODOoB3sgSKw6rLFM
UetP2IcpvITUEqs9m7pF4RMKooc+Awh/ila4/s5rTEWmJrX1p6/Amz6/9bAEod9Q
KQtlwRpt3Jt6uRmL4FplXP67CNVJzVD6YRl8DNn5vQlfy1BifMUsLNYeVuGEGF+N
1Y7CfHZeFKUBEIqOjwjxIkVPyI2czfuGrb+wml63BA9k6eAgOMZAGK3HwuNriwGP
+gbO/NOhVU1nG0BUMJkXNE3LTzYq2GaczBoYAbMKU0EhtEcOq4IjVYJAe7nH6mm8
tfmybg4ViKbUS/+lqDL1F2DpYZJhIZwFeEENeBU3fDnMnrTmDtO+Fw7kT4WG8YH1
36+CR0EKDsSMxr9t7tDaOBHqlRf+iJ6eNbeahMUuz4Ewn7dgIDB+JGcl83PF8esK
dpnd7k/UctjB9kI8OQLDHWWircM0L2VJPzRBsUHPrH285rhYzpcHHd1qNV8+2Jg4
kskf5fcClEI79iekpPunKolKFGJCR5FG5MYIHTJHhMqv3R5CH9f4X4yiIjPMsiua
s0aRV7LJ46ThysdMVcH92WVlMBJcj5eLlJxTYHEDvveY60MCVC48cBtHSxK5Njke
tjll++GleacG/nGwb153s0BNWr3xrJCde1sVaWLr/Mw6HsxAuO7b3Or5nH8sd9TD
NoarpL9BdUXS65gqtFKrQBziP15b/dDrNP7+m0liUXfu4gxl8cGAB0id5UuCrI9/
Adj/5dtXBSesrmWjCJpddWZnC8AWA5yc7YapJA741tsj3r18Bt42Jz5aja6tI73m
qIOtBE7COGnyeOqf3oWgO1UOfWzTr6lyuNzhxQdoAs31At5QcwxbQr/zdTRFajF+
ulvGC/t3czTQFRM8H9hvW9aej1j4gNtVsJvmHneyBi5bcuycYfoffu30mG/G+e1y
BtKfD9NM5Ln4ECGGxyrEupJeqSokA9XO9fgrk4qZXAvVOPdCIkONZJtzPDs5dR/O
Jj1AAFYoUY50ZllsglDyxQcNw8deB6ucTxaH5DgJhNAUaca7KLSIRm1T+qJrKRVl
Ecgj/573FiefGnp4vUlVvhXMn6+T2SGHeSPeOGfg0dV/LVGRcpXrJTHbDVXgW8fP
1XxcZk1r3+TIUcbe/zM+P8toHURHyd3esGTZ2daQv3UfZwPNDU+9Rk8xxzFs99bs
kLnTxYz0EnSiH7W4Z993dSFVWfh5fhqp4xVJNsLrteOesqGphbSvCauvaQL7PzNn
mQI/uGZ3CnSD1PUirfO9QkY5Xl5n3dlxBBOdLHmLSCvypqDMsYSaokbbD8QpYITp
jr6fvPi98aIsz0Qt10M+xXcSVYArgmf0+t2BoEsiXw7+P/y1HDvPaU1c3qA5Y8aF
CUYsK5gsl6oyJV4dAEOkoktF0lobZEslS/4PT6X4SwLh9SyXzxc4/MSTbsQgtlHs
cxiQ7D4+TyhPcjI/xQbkKNmlTdy1lRX7dbpfetmAkCyU+H8iZx0AcUMiNq6u0cl8
3/Z8Lwjb5n7Z5QQ0E3hms/5ArLxZQPVOhImhqxy97TffcWzKaHafS3G6Ipw1JBqw
R2I80ELtolOKKHQjIVYnuw224bzwliWwG401jgU+7kxMO3lebkqwWfX/XglaUBeo
F69CSo595gbMIFTkvIZXdxMtLzv5lr3eq1kM/4P9ARHSXFnYEEHkC81v6Sl75cAV
nDp89iW40U2mAAkzDChP+iiqwly0Al99vGrWEs1LU4x3kiYeBatjwenZay+UYW3k
np018EevtQWiw0gj81PUFelHw1vCs5ZVyHjOeSlxQy9WXBasfWvJ+pnle5pVVy7n
hvFM3k3cMbQyxvgpi2o02u7GEO+0+9xGNB53x5w9W/jpIKefq+ZUGceM5acy3v+X
Bcdh3Mr5qbVEmhUNddee3xpb0LXvL21NZ20X/Okr9XEno2SEShhA5wCv2tP6TD/r
nsfLYVowEw2anJVX6DgykCVWZzaep3kZDqdpG676CoDQZN9ZNBX2bRrnUrwUW0/Q
45XMJ5ycAyu2nFynO7zXUWR6tsK1YiXmsWIRGXDYiwnMT2+72xZ4sCu6/zAT1jYZ
ppwuHex9T6ndFly3HLsiDBmMdKuN7v1XgfIgTHdzH4rjCAWbcWjoM5x+zGNQftQP
T4ohAzg/3jslpQ5uBW4u1CndjlG6G87BsAalT6fFSjK+3EV/jZ3iIWpY1vCLo5ZJ
l6E0MfjpbkyzN1ITLdEBlkyLuioGo30Jp2ELkkb/RH3xGRCvxsX7yYiNwM6USczf
cPaOLxKvsx0wmSAeJc16R4QZMGFvqxc3DvNKiMvYep7GLQplo6gbnPbb9BA/o8g0
HuSF8Yuh34KaZsd1y7KSDI3fMcpD2Es9vRSxlig/QTpG0r0fHSGpuNf6/t+3Gby9
hLaJd8Q6SEcNMumAtwkCohlIDqwYumRGAHBH3C/GhTPQCYiI3IyDH0CfCD2iP0A9
bRFlDa+nHbmcAoYiUMeALISvtdpnjZwF/SFqZOjAzMe0uYD6iv4f9JCU+b5jTvW9
b5VHmZPRlorUp0jzCgDdeqHwaVGIjo5Prwb62GTjj6SyzfUhhvsTCHsd97xu2BCA
Xl45gdE3+SpYmNFp1a65pWL2s5A8ydVqkvnyoLUtZW2Ja0LVwMlAqHOBzHFq+BH9
c+gOYwIf5nCGJIJXXjlPLvxyAki+/zIF3TOYWuSIa7U4Nx7dFltjAvixJrDIJVWb
ZkwyrRph01BTkiZ1MFGVF2eP2L0gUf++p99aktMgPXv9Iv2zjujzTkKpCo3PMoGH
uLWUveq4n8wm5GhrxLNu9REzdtdla8lASAvEhkmziHVvK4Ihn1ZfaCkZaNDpmPGk
6BVJFDzkTtAQsLwHdcEr4u/0yLWLmIvs7gyyJ20QqOlQ78JOQZ6Ctrp9AY4JUjCW
lhgbspTtRuHlg0cIfnG1zY735+9/Jee2bSoe1ehHwLGwi7y9iTLjRk0Lwv6Jwajd
EmceSfum/Cu/tzXtEEZ0o5Tc4PlpG+505YR4/gsbTitjamP0y7gz4fuOqs92I5gh
HpmtMvYfXKYiE85c9O7GTiNv9ckJlS3kqdR/743DqtPIthcTnpHS1smlmhmgGMF9
D0v734CfCHyHx8szFWuNtcoZaPfGJU6yz1lNF452L1igZSnWvUquw4EIZtIyp0UK
vgXFNXYl3QvRT+xh/Z48s5/lbXp/TCyMy0ctbQCK/0gCoiYbLKn2m4DybLNAuZcs
ImxN0jrXh8fj1+4Q9HegF10zFf0/h0h6k4WipHB68MjyZV52UD3bziPn0K/QX4TJ
KGlDrHusp6vSbBEAt/5HIfzr3Vs8bNxOBIqtJgQZgwaBbt2YiyMRZHZNJRdYRJyp
v7O4eCUu0R1aUUnefQ1m3tx1nABqFjS6/mC6jzMZgjc6BFJlUs/h6Zu70dlIW5JD
MTFAtAuwZxLOUilhS9s538w4phghaeRFe+w1sr1T+gXpWZbclWwDMEgR3vXaPqmm
su/axU96cH58+6vl7IHSOh/7LHOJq8samra9aODmC+ng6fDVR08melmYfdBCqqAo
2bnGNLG9YM44LZZhNm+0ID9IAOuFBdxvSVE94vtLmlmIA6h2KU9MlvvoDs2Lcvol
5TRkLkVNLH8dwPlu6bCS6DjJJiE0tyFw0WFn8HCt2PjK1ys1k15RZQMYDnIHZiOf
dTrrF0TyqRgjjdcms+zR7sDKEa7GZPTLH6PSQ80jrZfIMKuISkxPNoe3lRqSNG2D
YA07yciMTv207Xa32nKh/X+KN0oi5QY4fkUx7ENjm8oUkR/2VyXzIb+0Z992aJYi
HdLrsB7qRx7bslWRzM3ZLP16B6JNqHGFHz68rI6TvCUxfUmMalOLnASVGSJUuJTv
9Pu6NLF3zwydqhgxbBVGvbosV9oLqG6G2lVQ234K8JPvMJfA2vqF1k3s2T9gt3Uc
yfJmrASx2nZB++IA/DO+GDUS6uxQFYEI1oV4fd6SvhGgiSHJLeW2gan2yJY5SPaw
ejFyfk7mMSY28YT9Bl+6Pub4WqtFTHAU8EqRHMKsvXuEvFzhcozgd+HVvSD7Axln
LtTVCes3+SEiaqJvQWaJ5HwTsfZb8mCaWy3Zy3e2ybvVKSuTtUWUG9UpSUDF5Q56
f10z9aoBl36Td7C9bm1mjqgSlud+OXvvE23cBcSw5l5KPlbni1XUTuYs04aYBqIQ
PwvHtdSC3Bg9huMPmLb9Bl0zlfZuuaqr/yB4mAZj6Df89eosJX50/mk6LoTiGuYb
yFURUBNwxk3LHXzOEA0lk/bfwyrGVEqza5X7Si3KCP/tOrYMzWpH1g7uvJuWAZ5F
f4n/gVpXGfQphlL1hkPeBabGcain303E7R9bS6guEc6kCBSy3GoGrUXXi5Xn4Qfc
Ayu/cU6ksAhui5JRoJtprC3ABaSD72t7OnZdbKq4sPtm2sllPuhQTjpjpr2+7KwA
1wa0zvdmfJ8BIdYTalq0bq9nZgjHGZUigsz8NWTw4mxDRgtQb/JB0B54AxUuvk9U
J5ZRXkLbCu5mYIU9aXcEhJTbwMklTIC5/toZu4+okSCObNMs+MAzFaMTfWEoEpDm
iP8KKLyI2tpjsB83dA7vvHgs7fX2GycJ9Fg8fMKdpf5TA/8wxIctAWb3kPeX3KG0
FPQjULYWhP8+TR8H24SxPAm3Z6asTpJRefxEAfjqcEhUvg2CcaS0xVxvqe79oup5
s6oKFu4B7mS/vbC+I7xHEZCpLNIHw5tXLqrEKri05Y6NKZMkZ8r0EZdAA9/rgSTt
2jptST3lHE5r6gnkOteUgWvWBd2x7VUSRvMt/wHrDkcN8vLYsau73xvu7JTUmnPK
giw9G1KEqqewa3SN7D/uQ9w8APubvwoQJDxXduDFx3eAPafCJoqMhJfd+tHY57fN
nkzsWGIKGkIGflIJsanSI3JahllxbV5xVYlzicISoBgWs67D2ycKZgPY86Z6Bxiv
/L12i//Sm3BUcfYLuowfH6dRRafo4TN6AOqpMfRajiD1JEONxHZD4fdq1za4olzD
Cvl7mB2miAGPNt5eQxS1CYDhdmF0pBPdUXjy6keUBJmpwLN099Jrf85Ez+qg4gHB
gGxFKuGB6+Fhrs8q66rHy435D1Vab14+8POQsalznkrVGL8v5xqP9BuSlbeC41pV
R/egSSZNLBnF0UbJcrvypRlO8lrPT5DGViCXnqYvU0L+lCr4dCb0XatAieNnWAkG
kNsWvU/lSE/yDBF4FK4Tx9EU9bPX6Tqd2bBzn0Uygaa3XvWnAvLWIhi7oWmoKw7E
1VZ91NtfHy1C8y0DaqiYc320lfMaAWFSyqpmSLA+4tKrqnAGMfWs9VYcdO1fI4gx
1kBgh6xCdce3fF1lnmRxeP+LMrv2DiuSgZF2cqrFdqUfs4D52HfotR9MuIY/qfTn
74ZwUbbl++gHilmuoRMZfC5zoI+lzWkFEG/KbDWxM/xQ/3c3uzctJxrGuaE7RddC
WdoZmurfYopNbd+lj+3+xb9mJz5AmRl9rhnvSisdG/axffS5hyeTwrs2IVJSc3/+
anECiu8UgLEG3so2yhBbQKdF6LDC2ioB5T0/vtVac0htFsoH+NDugHYFYaJ9nZXQ
YMxEO30XlLuJeUve5BJiFLtNOd1g1zjnNCanE6QHkh6t2jGrdl170Mgh8cqXhmIO
nHAAvFcznxyGZ12b8JlRXFdfHCEWpu5hbYJ7a4xt98UGV1cCASq6el1RDMgMg2UQ
OS5dTK6YTsokdmEx/xNALYkFZuxzEB6U4N6WkP9v34DBIBr3u1mMVqpOkEiGWhwE
uPZw1o5L7rRtLdcjTNpsxvOp8nHJQdgLn0rO3bD51YwSMotPuCtiTsV6DnpY9PV5
n45ZVG7Yxpv3RFWVdnx0DlRzFKK1Ia5viymaAmjl7eOr5Y/7WcDr/T6z7dkN3xLo
wHCWd/0BjqVoUo5TxQjdSFYv9oWXTtKFkgvBga/JrR13PdCoNNACPeOZjzM5bp7u
vJnIhmSowe0Pb/3m1JVPSbXCT4ars72WJ6UTl0xUJ7Ucru1uaAHEo5JhY/tiCZyl
FOOcfqXSkMC0/xfUp6irefh9uBlJmDCLMd4QqIlw4mL0VvgZyah6mBjNknOci+vB
gUtTahDJiv2Xlk8cp0HHl+4+yzTsPWZYJ/VA6cBptMcE671o6CbQJJbrU6I8PvuG
Dt9tSVWe5+vJtm31b+Xv4dfiEZqJfDsym4quCuEO0qs4Qvp8CbdcruHpttil5gSr
uY7rMBMyvw53V4ahfOelXYiQfIBhEa053tI2CvFWNjju3SuTxhr9LDh2WklVqVQv
oM8ex4weitJ5i0Rhmwlz/kUxlq3Zt6yEQcdV1p/rfNySiKnsVVqVnX8S6gallt03
GFzAVA6SWujcbpqOWRgAcMN3m2m8DT1wOspxuK/oRNXFUpyvx3JirQt/1tG+y9Yv
cUhMgFun4AElCU4K+LRlY//aSfyWc6LMYecsAuAjn6hVOGgDMRXQ51nHsF0WX7GL
UEJyxQM/Uk5MpUKfGtikOKud6AyLBGcL2+BHm0wtSnA8xc7vM4Rd+juwOdlFOA0Q
rmnI5B4QjL3CB19qx5AWacYalrRGkDhGE8SEnnkkYHhmyD/YUKEMDSr5goBMPUVm
1j1HZsXDOtQvoqBAFM8CtIJSi2GRXXJsf+GQK8xoPuGlqZ3N4gnNSpLzzkn/J6Xh
GtFl83AfJ3q2rO0RdGi2AF57OV/nkto4hAja2qhddWZz0WHtWkedTv4svVGOQg0h
aKQ1oW64rYVIW4P6iksL4B54feqgqNOPNYJsYnES9B2bAIojzwf0SfqHsL9tZmWJ
JUttba0mjtcK/ELRAkTXyQvwDEPV7aZTYJ9VdtXIs4lz5mBsCmHcjGF9ImmG99rU
PM5g7a70+1md9YFNjRNGXEWiRhAxQnNmSFMxXMxT+oq+u0ArU7bCgoVZyw4BoAA2
y/j43Iee/zXPyWN8Lqf6OFhHpgDhsdoCMZv/abXVUjmO9hdmNoewhDs4k/k7IeEs
ZOtVJDYKNx581Ly61/TEYG847gVm/rja4oqyMW6v5y2pb4YyksLt1ZPqPcvwFglL
LDAeZSInBH1lmolwYujQEkH6EJ4Bpw1G6ckXgI65FnJ2386mtmr/9dBtii3/k2xB
v92cuYEv+DrUXIiqg7DAzLGHgTtrHPVXkbKY3Lo8z/10/iFBblHSJ+Wji7IO0wfl
2KJMwkjxk9zYKplVPZxhkS6MqFBhEAh/ijcozL1MxVBqy+UjS+iZkdykvRD8ps1f
Tkh9szxga4yXiDJvsF75Be8ECUo8GtT9DZo3QqSMxjV60acLTelYLpWgc5uVHxbX
ctu1bJae9zEj7PZjpP7cSvwXAzdyLvbUK+XVPdwMByIhzmIwZswdwFZSMfUL0CaP
x/aQniEF7+hN4kCzGkA0OOqYzg4JA+EIg5XO09lTDlSNqh4AxeKPg6kxyB1MPihJ
+ZOPaiPSd/lTSEWOgJ+hPULop86HhwMxOXrEZ1qSkk9skGqdSMEdrRlA/Kcz0tzW
O1xe0uak8qL83mNVKkF7gIKHM0omIVzOex4o2/UumTQXwTrSXIo0P5OpTn7iaccX
pOfOxjBxxqbKAXnYSr+zvyBrVDouHtQ5TByVhExbIrYzad/6xXvMEnRxn8L3YrWP
caUWqErfb7pZo4tNlRjz/3qz/9a8f4xtVSInz/JNoXhX1uV04chS9+gvaRpvBuw2
u1DTH0L8KWfWCzQDeYBILqmPZ4YKcTpoRf7Lhpi08Ha9lz6BAo2agkEQEahd4pfN
cLnKlFRDcBXU35YuZ5Cn40y9WNeXcKaGVm0awInVJw+VU6+lPfXrbVl6fWaY8Fzp
Ec1m7jsiFuG5qEmVMJOE0toMygynlz+JpoWYOQLE8PvuIKJB5wYmcjACNdHIffN2
rq4GpbNKinQHeeYXa0H4ZHYyjJD8myOUpbp7XGR5U6vffjdcryLQjLIOccDQ2GBK
+ajmntK4c/MNtsmbQQL+leeXp+8ZU7rIE4pkYWqel34xIXu6IioZdxLq9rqLXr9O
Mp0SWCIuI7+fQBY1ShIB5R5lfC7izk2IiNnYG32fpgf2VyPZuotafGvj69D26BOn
w64+3ivV1khw9hDTiY3sNCltd0nkSaRYjz2bGdRIV1kVwfAqz2TADn70mM3n6TSB
mqKHEKJ/vK33pKEdL9qPTGlnKEtag2HdzmSEVewLb/wd7eoFfGJ8cwPQaSWpvewe
1Q9cb3TaUH0eKx0kFpjIm7zbYkrOA3XqQ4bYekrvB0Q17JANOFsVbour4kqQaO+V
tx3V5PNl5IkMz17d4RungXN8QY9hXTEeeCWHc5XGnCe8YcisN0VQJ++M9Kv1mVRJ
3SLznSgqK+6WoarcNCXh7sM8tOiO2zso4J+BRcJDuc5tLl+Jp4UDbehoexTJuTQv
Y9iYTZjBieRPFU5b2p0GWCoM52gMEjJ5Jw9cIPdO3jSnS1O9GVvFPo/1ATlLazhX
G6I0S4mcb4dSeQ7kJKiVOnjyXw/IDN1PQ2TXhLHYx6y7n/IhRnrWXSzG26MLik6l
d7qG/avzeKweW8AwsoR2gkx6w7zD7oF9v7YcZ2+n4lZMBQofDC/y+L8tV/rVG9M0
6mv3xT3Fsdf+x+E+IUJfaVPkz1udGbk+OEdQROqDDQrZeKmTp8orEdYK/YDFTrov
bLZltiFDiA1sMxiaYKyAjRjNfOH0HJJcZT2Jybym+GTxZtXf1JQnnQpDrUMG4nIZ
ffkYnfiA738F2o95hSHYkPjBTZHKiq+JenwhCKAXwmm6gliM5efDUJ4TpT4T8uzT
AVGRgBYU0loN3gYoOCACYeoeIcZWj2PC0Svsgb88vvjvfcqngtgUEl4p+8B9MdIv
XCFZ+a6omQ9kz0deZ9dMcOS9IQ5x7M0o9EbvVT7hFzYnlVVkdG/d//rLi4+fIPy2
f+L1BbMMPHeEMgTtiNzUPmreHoiWmYZKANW228LME2i77jrfr4MFzns9jzfH57N4
wWxxl66DZtuVdub1UaiYC8QN8qBi15MQ+roJ2UWII1BLrvKxQCGniynfOrD5Xshr
ZmfobgZ7KYkwABOBpZvxWtCUp+XYfaW3RJB6EtzbvqEZGU++gsbLSl7mAGHKl++i
p5jgeA2fMK7EPpRv2DWOQqhHC4pT2/92PfVTaG/4tRmdq1a8Gb93Fa1RgQoLmy5C
s3s+71c7Zn9mRb7wLrtsbk/ljMB9oNjkt8cP8mHXFQ3Zjil/KzT4hMF+OZLa2ir0
rdQZsQUcgNWI0Xcs37osk7mytMZi4lEQIOksft0rBIUHBGyPaPxZOrCHCscDf96t
EV5XZc+TMrM7lhNZOjhXQMC6VAw5eVWgu41uTxwFPwQ2RInnH+MwOn9KmGSxYxLo
3kY0sAPBCY2mWtxl25kZb6DER5ozDbimJFoxqSchlXskMRW5w0DboRGLwg990lQS
CGDEQIgLq4f/cdWSdv/Ml5jaEQjN8k7q+h/07Dzu5qC7YRIglq6mQgusnOSMkpeW
jxqnWRQEPZrbPJ8AoeulqqHa3jZJjLaYuzDlh6EJXdRUNBNDsdlAxgYDBG3WttCu
wllN2ZTxePVUiJ3F53N3v97LqglD3RByI6QQzeix7G6RqNvPRPAgCQSyXEQseWX3
Ms4UJHfgM3elEoUwft3P5eq8M0BGjeL/iMIZUrCRyJUkRH3d1ia8gWSpB0v2c6k6
gwFU2/7Folz74GrDhGLJuJ7F2hhX0bT9EXoiulBjh2uWpKbg68Ognd5AEJaDZ+TG
bH1nPNIdcLO8dg6MHStG2e/EK6wWwJYaY2qtuIW9fYdK0Mbno5eTB2jmYSjlKRbe
CM+nS0DZ2JKypVqsDyMQElbthb3Q+BWufGu0agKnjGgjBNQhaM9YgmomVUJAEFsH
hVsTqf0Ox2BTY5CX82tbG8dpEC/d1UIG98S2xQB/4g/T0abmSNP0Jc3EKLo2o7VP
ZLwss8yY28+O2ZzQMCGTJR3nxKHl2I06/hWGJiQj9BoZuoqWNdE44BiyVWjRE45u
AZKv2/TGMhqFgOdUal9nPIj6ZrqiUdI73CyewpeAyFRo+thqlizr1G8AbsLRAkDi
p1eKLQpCM6q5ujQzPwSdT7Uqk7iztLF7BcXMN2Fxj8d/6Oo1xJcjw5fCnbuU1aEr
n+1xiaBqsrEZzKSuUDswUQqcKKVbrpHrXsHGV8g/jK1qgSfxNjZaH9mvT3C06Vud
lVKGadweUSui1xeoABFwtU5Hcfyzv+sGDw66+lwrWpzTyk6x/gZKE1KRZZOnh3jV
m/kp8q8dWByzsdGb0/fR1TQbE/s0hEQ5H1TcJHLKxrYbhw3sTPsLMR46x9bNSNW2
MJbI0yksJ2w/Sd2WuFAh8l6h5ttLDNQWKBOLMbuNxqvrH0xVnlzIWSPxM9twhpzt
bLin6IMeDEjgsIibtGdR2S+2C9AH8sHXt6d5FrkMUzQBnqAisWqEyvn0i6i4K94c
3GQrc4Z5w7wu8KUKYKhN4mF5n2RlmrDtC2FjvGdFw48rs4lkXlRzIuvalqNKhCyl
51Lbe31u5pm3yxkRhI8AjV61FHBVauf/WbKBfcAgZqXFp10iL8nDHctVqUBPUdk7
UlkXNfOcU+tdhOtZOckxZ+aLe/Ov+3HZDzHp3rR3PorVmkj3Qp4TAtHu6u4+W8u6
d3LTavKGHJmo2Hy14LpWJRRK0TwOgX+lOcXhR7s84lmGBwt+Q2tX1B2+zd4A0z7i
Ltpmj2JqRlSciAXY45I3iWx7WxjSDdxpgppk9jq5ilcZayM28z+gjI5PwD2jSYgW
8D7ss9Uw0Inad4lR7obKS0nVTK2JrzIclsjKiSqIw8OLWolPoymjgVK+CgVgBoHn
DhKc0SN3ppLPrujLwzf6pQ5oA4dEJG23HH8l0C2tMMmRqLYeELa2nwrmwKR7o9TP
Bsi6dKR6uoj/WG9nS0mSoe+vjwesSqLCkMRQVh32K5MKK4zGGtKhDgNmw9sK2Uc4
CXTCgtNfLocBG2A7TTrTBtFB7qOsmixyAkSaH4BqQCEHHZNoVWcxL/DH6zLBgBCg
DoO+njxhD5kp5c+y6WhbWau+ZiP7RVNrGyCJrVebds/GNWbtnzRcFRA85v2N55r6
slfJHCpnOiO2w3UGcGkyB/BAxdGlnglDyEvg+a7xU4P0n0JYRGIaQ9fV0H6rsP/W
njJemSwuw/xuVSuqovIAqmyd1K5kyTucgTm8/myQwv9TH8hxjnyu5RnW0Ry2cjp0
vvmoOgp3vP0NCE8kaUcwekWCFKnkY+/by1wXRiAAaYxHSKgBNH+soHsXZF6o1sT2
us3A5iQTW239kJvr5BoPjA467OyANolqnIGRHcp7UKhULyr2dkLVcxth6iS46Zqv
1ypK78ebVuRGrHfI24T+jFzRsIpxXINTEf3D1zlvaQ5vzCccp4KZbtUVygbTAMfW
qhqnrUO3NIGlWWuKSvbSfgScXRuUCi5yXtdECNt7ukA0gdx5mEJhOIpryjdyEADx
cCzCB5GutkD49j58xzFWBgPlOEh98bHTeMJr9STAt0hXqDbPrE8aQbnBXTyLSnho
0+qm35VxKFaG5Lw6UxrKbiQnvkyiovYJiEOc+2Z92+FMsYjAcZh0kTi1AxWQ4uCI
GTuKnuEGQA0A++foyZ6GTapIK2pRnJnBkQucPagPfTPfgXTI/Jg81Tr6QJM3R6HN
kZg/nxUA0RbdCO7+rrsJebUlyHq/WV9lYEJP4UT+w22hP19neL6J0BHKVSlBSYKy
OqoFel/OytX57Pyp3l2y1Njj3rB5I/Aiwbv2lPX8H5JRmHeTHxfEgVLCPvIAYNpW
eYNUDnt6FZrzxWTjjYqHK5XdXmMVDaWSEAPXgK/S3smSSamGRF+H8Bfw17Vc6I+1
KFUnq4VIJXmw4mCePu/5abbOPympcZj2uONY9tjAk6t7URf2klLISDwrcrsy9d7K
ERsJhXMuGCwBPJ02+immIqc3hQeMIbnsB9g2xRLDm/k85PUYxPiH4m+dA33+Jq1v
+PCZ31vKZDR1a+MP59U5TuggFx1F/dlY6Ez3zp3vNApNiWOY28RgLY0iVbP1pY4X
hhMaEq9YcEYm+uUMuvTRgEuUrYgeYQ1te3pP27DvYRHuYk1EXNYSkzEnk3QqTbq1
UplMtq2jriUIfFREwF5YjYnbZoJLWf4QnzMja70bpkyi96Kwc+P/TZA1onuvxfe3
1AM4Kh9R+Iy8fnZfRtn+YV2mwkdfBuAuC1/PXaP3/ijs5V79Two/uDubB2QzZD3o
8DlaJ6shU7dEqpF6gxoAoxVggt+gAww1FsYeW9YJEDvrR8uyXYjSIOVtGD5PuP9G
Ti6PGHsOTnC/+s/m59xo0rnTO3sGXGj8JrnJMI22cNPVcuI51XW5z+LdvvRJBCNS
jVSMwmA1CTSnJ9QWIdhtctXXpLNwLqlrJTtRt2H/tJGoHUNeuhTaZUg0Ks9d4kez
ghJiDtrYYO/O5NZXS0Q/Y9GvyEoczu8b1/L8Aa4vdA1wUdGTancK4vf2/t4KiI9y
HMbXW4HBERl9NcvfHFp48SOyN892gbd71Kgr1iuRjaWiK57segEszPbr9kFoNwCC
UcG8hr6ns1TPXZx6My0ryh3bHaLiSUHazVkxq9xX7kIwwrPCRpcYjJKx48lvGxVF
tvhUDM0lUa2x+QKHoAgRjqryxcj3w9RV5rdJs03j6GRoFv+vFBA0ux3/aKxtRY1c
DkemFzKs9co2GN9b7s/iojTJg6cEJCxWRiAAjhXrPhTijXtZjGCO+/+PN7E7RKTj
Xw/7HCXn462xXvGNNJvzlx+wvOxK91HzBF/eA+ceM4ZhyJQG+b+fIjnEHb2LTVia
SkLN0HmStCRrQFyKOQOuKGOHZuQukSQpMlFvuZTuvXnlYGQ+Zb0Nzgj7bLw1GUI3
Pst73Fp2Whi5lVtxFhtzMCC71WBURarGwuTJDTK9vTgGiw1D2ozNdwkCfVE4valr
SNN6WNs4ly35qGyQHcN1xsuibP6ug10aCOBEZ1JAdaUaFfxZgxXA3NC4OmneXku5
uSDHSBgqWVb9HDmBw/Cs55bK9xOnXp6pBNi9fW46eX7Hffk10nqugu9AcjCXHoYc
DGeXe+FqZHvy0rOB2CKUxEMJXQb3n1AD1MUSt6GlcLX/sRLJ/AlTQXwAJ7HQsPdx
Ye+iaL7zS7DdCj4XDSh4bAD4yBTQC9mqezN4HOz7IKwbFf2avsleY5PpvVvBly1c
0JIoCFYSYrfUa1wBUBHjOcpblrz671xs99VQyK3kyCLFRGyITc/O0OshAlm3L1F5
SK5AxXzQHMJ//az2DbSnu+6teaRHJBzz/zveyzOWbJoNpuDkFanwCYJwRrUEsKOP
vHKJAwBRT3c4zxJpShizwNK6EgiRMWX5ibnTyZgv7RBysFdXGshDffyEQ0tfhyYs
6RZI9GdOqK39bmka+SwXlewdLKm99JhQduq/IN6I+XJg2Y8HIIoZYzIlblqd4JBj
GaHbwK7t7giLhVBefeFhGr5MBKDrob2OpBQmx8YPppwgudrY2WQln+FgwmQDN1k7
yb1OqIrvO66GU6QgYszaWhhNRxlF+UfhiKg6M5lRWe11r1CuWDWWn0MD+C4itWHF
8mzoZgXDil44QCV2wUydOLnk6q7xWtidon/t731EPpnYGbUV4+FBwD40+ufvR5L7
yBKEvac7dRk4VK9blSb5YPbXOFeDWZ8Gcasj5ErClVNSvrOIwtrcZH3ksHA0x8mg
5P5xuvxPgY4R9zUqoqi94nFHbcrWCaLUkz/mLHoiMHIfjYa6NpjRBOJAj+2vRDh6
6rhA6i/d+qwnvZ9XbMQkWVjSm+sEpPqTaoaHYiTTeC3JRLHP/IMI0epUXFQJPo+9
2+lev3+q0GjnT4iMzrtLSVIQkMmEJ0t0lbjnQUDw9d0AE8m+ng5KmLEjsj0KbPAF
geByQS6zgX6HC335j57qaTIAzPWtFPb+YH1I5sca+17Qpmz2Oyr10n2oGgotPTnJ
DR/TftN0haxnWZHk2IZlsGmXaAp0R4Dtnqx1y5OrmfMnVUCfMWrG9nMhozjHPSUI
wplXjIcr0dXu0f9XTDM3Cr2rHo0rwS6FLAsGZRhEZ2GkJqsMr/XkdHUx062VxtnD
MXZ/QC0yOb2EgYkVWbSoZupu3NBVZQKDVXC89eSN1Rvenlbfl6Li/xppf+laaOlF
4y6pNTAzYjy9R1Jy0+UlVmxf+zMLaJ7hZw75Zb9MhRNAlUFyg2YDhDvJD/hgkay9
TLzmQp1ZhPHausbFr2zXOJstRBwuw+ga61uS5CDEuIR95Qmshi3dqoCshAjWjaXD
/MACoJJMLaCc7/8XIXztdGHUPYVbXpCPycedw/35uHk/DlXpF1Vs89sgzoCxiuQN
6MecOf/M+z9KYcw/47HvclgZd9dQ/AwaqQPjVQl/O5gDPaK02F2OX/D8jKVNA0u9
bebeoLtWn8XCAaABkNjRXdCPYmS3skjVIGj/+aMPaRMFDnwqzFSn1Byv85jNylzy
mSeMvkIqmmIUABIYmKivQ3+FGj6lQ3kYl1ovTDwOQEY6RNrgGGaX6QTnTnL0h5kc
5wcjEY6ytIGMTMcFFCH01Z4D7+d7B6pHa1WIrZfp13yqIoS5VdXVNUQ0aSkyoUWP
ll85ekv/OHUoKBK0hhSjyyD14KJsdbAnX17Cw6RrSd9y4PyZby0CyOWtNm5uUM9w
CsxbkHesmSC44e1Px+cCHwczQHPPG4K1rE6dxUO2W+7jHqxzVPPGyRc+ECdacQTF
S+m2kv522C1axj5ZhnEKMCtfE4MGwPW4iSrkQlvhj66Tz9iQxV8oqu5PMniEGuko
ajSLo+IVPPo8dJUIZDoPcpHlLNQqzBaXZ4+hRdr6t+T8fKBPCDTWxwQvC5zZuOzp
nQvHxHqEgQcpzZEyfbBXl+LW6RHSY43a/GVvEn0N8yBli7wift+e/zDF2wj5knci
c0pib+jSWiceZbRPol+c311bUFFH0gie6c1xcxM3DAkKRbG4FPbI8BrSiHCmVEGv
gA7YrKyvrPbH0f9xJEoXoJEyvkR+0o4RMOLuyGOdAGrjgqCnH6kgB5VYBcO7KCvp
0TwGxZkP3j5NVMA7gE7zpCN7LRZXSsWjvGVNUSmrJZY2guG2Y2f9tQOJ7XLMbpUC
C9AeyHurnLk2rkXnzxjC6jyc/fs8WNzBHRcZCNWfVoTBQWnbEtgYKWqJUKaw79nY
/v4qxnneCaIn1uUfOR+xQVfzS8DyQoR6KTfruQDyYSbIfn6MTrypMU3J1muDu9/T
onmDPguyGCxusTaNSU38ytbbW+c9xK4c1ivjy5JBkzv8eQe56LBGYBJ+TFY6aPTU
jj6rJnEqL3DW2ZtJqyP0NFYOabk+4EfgKlN9e+OcCr11zxq2Im3HTUuTXYyrHMye
ZQgBlewyYS3q2ii41V1TP26KgQlZxFibOhccCg8GaP+Ky8g/M3NZyMH/2Msy8ywF
qeHjUuyPn7QLobu+KrgtKdXS/Euh5tjEY9Zqhj/0edveZLmZ1LgKGmKO4/fIFzw7
VfWtopJ2GPJbK6O0tQ+pxXOAO7h3+lOXQCbQwC2Oz6ruSq/uKwcl1JM6PTHVW0Wl
QmtRrGalLxgMOKKsUK/FX/LoyNVxpGwsO1XeCmca1SfwBNx3R//Dd019q+aE4UTT
5tzBAMZahAGlC3tKA4k+Y7jzoJsrQ2b5/IczkC7f5VqwkhnsZPCJ69H76EBYh9fT
Zmfgy89RkxJ5UEEnACDlGqwNxB8Qz/fJD7+10yh9BkfTDTaylUE6imzfzSHTaTwZ
qyRu0hnLp9eBpevzEjmUtIdjKB2SBDP36JS66Vnx82QaEvF2GaUK0eKGkKV0O7AC
aKnXrB6zmK/411JMcCWF4IIGruup7tUi6lMUq2LhtOZF3Brjy0HkIYdUQpn6d2Dy
SzMeh0RbB5DXy/swWyg8EqKe+tP5cUsw0/b5NCP77Sv6ZNfW8rWaA7ca8iWzq03H
drduHmjp5Z1j3Hkc80Nq0LV09iwSnoAaME/pcD/i4Ryc7oLZZWmCmiEYm6s4mR49
9CetUVpwRtydP+2QuJQnDmkgABHB/EXmTufqDEb1sQOvDvKMgnghgd+qqTpw+7Zg
NYGdghUmQK0rlVPtMkEGo6wLqyuBWVRF+q//ALhfVLMAsSjM5MSDCzvRIgZGUz87
fcuK+5VhpmIZ/+U8kA/2ocByLHDOYU9pISbiHf3Kiyneowq8h0xXubnudBCYG8lR
5GKhAPXLSY+2PKGKjquR95tsPxVyaLi2eA/NmHkL7m/P6D5oIdaj+yXiKx5lcofr
MyqpzlBKYkRcLq1NUSmAAvO+XY9LjoBjSv7QdGC6Y04diXDe2NGkkyLpzbVPopqf
S4lO3mi+4vBaSAfSWerEUpePEhal2fQF39jBGtpbFhRtMmvF1vgdDM1oaw1n5wRL
Eoh4vi+VqBqdzJngF2RWVyxn20KlwivmoXJ87tS7fjxgEk8VwiHmKw6upO9HvlWr
HY9rCoxN3lJLbgfFNf4tKZ2NME3vI5vyuA3UgXo8XC75n4z/h4yyxfWHiXXTJ63z
wrju7a6aBSgh6+h9VFKue7hbD5sw5q+xKJJvg9mGSylinI7D9m/tkvIg6sop9LNK
BA/zpAjhWin3hlPMR3Ih1llkGQ2+QWk9kPAYYrpTeepP5nlZ/ISloak3aJTzGekD
ja9FqKAQ9KjASGPhvExelmzfNG40bycbw+2S1DSWApXL0VRB2nzWtRzkMkqFOY6r
T3BQ2asFhbUafy+/E89oxPHNPRJKA+TqdOOzoCpjXabZ5QMhWBWogQcmmE4Cn4KK
4hVaX1xpQWCH66mQYvNV0gEWHokNuAdOXTE7+iBiz+LCMvRuwTYiyOvq6eJsTRuP
y5NXMST4kbwFSL/VSuGFT8/5RW0uG+RVJff76O3VXRxPbJ3Kn6VDRUHI0sCCFCsa
CES4GKesp/BAhBCVzCN7JZwxTq7vt1mzU/e3d1t1/ceaoTN0VSGZDvHtlXrGF4D/
9k5zqc38JIoOhnpuy9asLbXwDiEM/fVyQGBCRDQQ/kAT3lPwKSI5MNEdCrYjSL1r
YPkrXgfslaOnK9Vgc561jJ0SQLi9hC3mMNAfmK5a8qjqSl+eExnmquTXxEwYnL5p
tRK5oU+cbHiUDIMycd+Op35kQV7Me8q+pS84uyRF8X9jU5ZHMopyeiC68GJ3FuVN
3qM3OI8Jez7Y2nC5infYZpQzMd564IxtyPWe6O+F2DhWz5YkP6u6QDVXcpERqrQf
QhYFndsZiOfdYIeO9+tBJ6Vq7kRWAymUXKP3suE+WRQAW8Dbeym7FGJ+CbNaOOdc
dEf7VZIMi3VbDqCSVrzZmQvqysrUx18zDs7wFU6xcR6ZFVjt7a3gEwdZewgKA6Rm
bsP6PzIOlHVKufdpcxvU9li38BJZGSCMEA71J/yBNuTCxiCtjt7CkcWSPjliTTvy
Dz6msqdN9zvPSYQ3YKTQBQ==
`protect END_PROTECTED
