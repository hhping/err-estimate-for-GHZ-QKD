`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLTkVE/QmEllMQRduPZVeGZrJpMitiNq9Em0/UsbfCupTqjsA67yOxo+uYM3SAsW
8w5cPEU4/SMEZMuqlWlobiCnEFu1BpZTanaupltCVsV16mSwdj1ub28hOtMvcc36
voHniC3eZjiadJNp7gzzN4nWE8EylD+KlWBf/9qyilHGa/ilwhtbasEhLcz60jRG
8BlboccyBwzKwcEvyDRoHeVqhZXAggoGqFnlsbdrn8hnE7aqBf7I/1q3u7uzwGNC
pLABwMC/Uu9gsQeYd5LgPVeTMA2OVqgIXx+I60J/Gkj2K+qjtMZzWJyIm4y9wzrP
2D3tVXn96fxZCLG/YvFCyD6XLlmLfZPCHI4Y48ZFypbKsqLs48F5jTg9YC3X4xHt
hX59xGHI+VC+UpNdGCwhuNSUvixLVGBofUsIy6fzL76YLYGDhpnMP8GttoKQIhxi
D6F4bawJYwqFR6K+ictxxWJBaUW275AbFrxLFWZyd0p/R2iZoolLCoymnVHKhwtI
ue1HjWLUimlqIsLTrRkgPqAswI+Yx7UVIepToQfhrlR1Y8vX1KC72tEs9a1FUodu
`protect END_PROTECTED
