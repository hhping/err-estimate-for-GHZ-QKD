`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umw5vOhoIBqfZK6XwTsf/YazGSKUyzGHicrapDVn86dHD3O6ShoNwcsh3fTRXs/0
wtfNnJ9XXK812QnHHSGhs2CsG+EF6YnqrlDROLSzp5n92EUbsSYGCqhLSQTYIkb2
qFdnsHPzZlIW293k24rFeSilu+ThkMJxX6vA7zsKw953gqGyDcVI2WN6SMo6BEPK
6TgQbRg5YKSd1w86CA20DusYpE2NtZrzOg9niD+6SdcG9tN8mKkEDUSnLh1ffX2W
UqiNGGYp9+AdCuu+AHq8Iw7HYr6a5FLdmmCeGSTnyEP2sxCsEI0/k6xhF6e6bbI+
yZdWC1jjAlua86DK3MyxSSYU/XiIysRYvD0ppos+fD0mW0vpbz3wQdkMMR31xh+c
1t8q1DzG6nhBcWJZl0TVadxyNvslNHIoW3K5Hs8M6qOOPjoh/YkPyNJKrw/Vl9Og
VyzwvJH9ky/ieKExAh6wsspaoxWUw9jW3NP7mcK/XxJa+6qbR1IcydqG/CNerD7+
BXwEjfI0llWT/CShNVmZb0buKI0QYx3d9DYP7NmfDxpaxdMzHAh06VJ8+YVvWQrx
8U37NcoQgkBdqdVkEgRFSTp7+RnwMpG86lZJKDzgOSKCuyb9JIi2TTnnbnoN0/CR
5fIni342gIQbiwKTLJQCzA==
`protect END_PROTECTED
