`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ec6I5uk4fWfmGJfbVina8HydIU4D1oKJbC4RFuEFG1OqHF1YJwpT79j4tyfDN5JU
1Z435PRbx64pc5BM+sbye/VoSXTr21jsg7JI/Oqusz+piNa0xYYLakoNquJ6+VTP
m0vGFXN5dpnDrCZXvlq2d6Qcw/YmCTJTHvmaXVy6I5GYaSDCcETr/Vy5Ftzk+wON
10Hjdm5z+SnYTaKUsDLZL/6Jtuky2K1wDyUvsfm2i77WPNDSzYV+b6xf5yt/edDt
pML46OXCK1ibH8yVJHNgFfAQv6iQ1GTX90mXfj0e0yR7Cq2ymC8E63fbcJvqSG0g
tAt7M+3jXeonk7ccwpKBx4OX9avhQC4OH6yuLPxB+ffNILlL9PF5jJ/b80Iu/llc
Upkmeb8GgFYfykaaE2TE087gt0/iOORMlC2Wj4SpTQrIipWqWEl1HEwErT5k0HBk
fN6ktsufoDMxgeGIJZzXqnhY8otQDZIO+aJ8DRt/NhYnuh01zEe8VCQcplDYoiqR
6mW///RDN/mj7H9+iIoN+TDPjnP5VehPdLD3Zzh2Qc0nV3N0htY9w2ayZhmoPtBc
DpvNXoWiZUfrEJVKXN+TOHecPdLbCnNnfIhMX3Y/6S1Kwuthe93L1lxmzz6OsoFs
U47epdkbEBHGOSjqelQ+neRRpNk9xB0TPfiLsG7V0Qk1kDw27+5emDLdkowYKAGj
lMEqVw7B5jg0hI7wmxp6Fw==
`protect END_PROTECTED
