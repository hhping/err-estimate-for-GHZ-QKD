`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2oc4fxZno73BFzfdbJJgw2bwwwF6uO/iKFqCB644l4YQHuTguooI61M/jgPAGK6Y
9ybdyDszFLHmqPpOWUrvRqyzn5nBYeXUgpg3TgxLf484ScsliZAguvT5qv2V/Yil
+iYad2TmIQbhwEVMsgTFB5qZVe9zcYWBAEH2yydetFFvr/oK+NY5A+zDjdeoofln
2u98rYrfbcmUvJ832C7liwfBITYE3bn0XMkKvz5b2t4Zzp8mnfy4B6TMQ6ZRHclM
k48FI+XjzsoOabKweOR7Xdy7OY4CTYqaumDyFr1FawDWR1SblnU/FmENlfMmbBb4
fYSlZLxO+0kV8+DUoEb1pfbGjhCce3yDiWu9qUBLwsrdQXFciPsd3jraqGJTqHTC
3a6GnREfuVcZbQxURAgHuqQ4lguqMr4XC1uM5kkW0SFzO3FnJzoh1NE0YSMR7LEU
5DaAbWd2QjpJ1ZcDJZvXHl6uMPYYeBuJoePOgOCow/GRcj7aKCE3WB5O98J9dTDk
XbdY/eEsE4G2LRvcwgdFePKhJhA1Gb+U4ruNneuDHIkQ900hFF+sSy+VWH0lH3jE
/pFIOxZ9/Vxj+o+aQKzQE0PB+zF1Nie57iqB+7ZgzLE=
`protect END_PROTECTED
