`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gIecLckJkgpJy//CApwEqTbhchun6Piwncui0w2ZSRIdBnznq/kmTnJ+6oFcIzM
YrJWOY4SlL1vVg2Oo/rqFEABtcjWcfBjg6kptmX7KugZVYnlOb6eclAsJE9XDxIh
nv3bo+hC+CnduypoZYtnuRQHI7Xq6GwKTy/4+qHd+iSk9Fo7dVe7TpevLEMQ9RHm
mCF/KU2tOA7jL0CqwaF5SrW+o7wkwytVBOP8w36J/FZJcQnGmgywZdlgJ0iMQiQN
8ftOMaSCUCcQSPYj/MTeaEDCN3rDa+S09811FMM9nPRZ5k0yJ/+am/lLb/yvJeO2
cQh1DT5T41wZrmovYPoX0i5FCIFvQyHnmlPS5GGsFuMZPSmjMc7VSaUNRcU1gXoE
GkpMsPLFE/cVwBLJyhByD0FhfRBxhG5qjLB7JC0yHv/CVOYvZgCs+dKLtOGDyPkQ
HDBHo8lMVhY8F9/NAz57X4OkW/Mf1sp6KVuh2w030hEGzLV6oB7AIwRhZwsJDJtu
IinIjZ5g54zybCU2vX/LrCqqed+ydD1bRKlFwl3Bzst+a3vSwYxAgteiOVyng8pm
a476LXHTRUrPYHc3h6OjnePcwCQ7baFmcPsLuf+ZAsUAX3K6YKr39cH8wwInrYJJ
7utz6w1LwQl1ajI9rq+/exHbXqCG1NRJ5LrZin6Gn5w=
`protect END_PROTECTED
