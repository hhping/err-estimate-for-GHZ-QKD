`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82bHh8rx/EitHbn0WWb8y4R7YpEGiJDMqgW08Q8+8bE+zutL/NJAC8QnCBnn6a8Z
PjnVoxZYVOvIGDJ26fgNr6wcKGxIPKbr1i8K7piTh9HjjPbzLi63cs4b6z2QaPog
2KPjQKKff5kNi6zWxhawvesjyVTbQ5E/7oCCi0hrbqM011wHUajJzxhG+tAQwrI/
wF7PBOkhHnK+dHyj57ttOf/VLhf9pS2Q4jZdCqmGVvVm4zZ3Vm8nme7+DyCMQ+Sq
dZRZ91zxshq85Kn1Tcte73yG7dE7vJYw5rpZg55MrCYX/kiNbfKhybU84jDw2eKu
yS6wsOLGwt0JUr2+NhzcTD2bacmDxxslKoSUZx5MUJ06TsAOOoDQDhg7QJNgbKiy
sHHi02bJ6yTE/oEhlKYznuKdapI24pkdqUnbA1VR3VkSlIUKskh4dzjrp9rJTnjz
Rl2r4DDKLDfUhqWDq2SpaSrNPX2EavkXL/pwdJpeIFUt2j7yDUTv17HfmyRTM4h1
9/RqpLMneudu9xdGyd7LklUW8/xDo4ZP28DlwJhvyyZP5IQePNh+bzjQjt9Q6Gmh
0m9RTLpGS/IMni+xgcotXi/E8nlS3n5+DNGj+AogeOcXJXxf0mLq1U6aOtQh5x10
okoNtIHhLdXu145ImVW0HJ5njSWEKMZNsXNJg8c5/Me2LG74Gvvc44AC+Xnd6J42
CQQsdV7IZumunq2OppJTbMKOH4m+f03lPbsEJ2sgotyrP2JndNAONpahEZl//TUT
DvYtn5o9tecdsexsLRQBbB3zlR9YpcfiNpAS3YE5eo5tel5BvDJL6tHNCDHnrHN+
TOxjEmIZfEeHjs6wHRdCRLhYLAopCjdlL94/dbzuzkOVCXsfJ3GtmXcV7rdY0bFv
kkkGgvYLittIYSXDJwuao9Fa7xxJ8llD1yy5Lv55WFWGJxAN2y0XPE9p2Rph4wKO
Q4AORTHnbzrt2/+4i64aoTZWU83aTrBcwgWTzuViUEUbmvxghjArMfgulUQAL2j/
kU5+/gzDyEv78j7JqDWXCqNLSGPxzQIp8JZ6WwRqUcFWXke7bXRkZWzrGYef5eY6
7cqqxT1+XUDUkoKc14qeMfNFRyldHoMVeJ+4Wygb00oUnsodyu4VKmv2Uc5lUeuY
wZMkWR3TdlXvJ5Z+p3WvfbljczzRclRPmzuYlY+lhnU5JO3BDFF1StSuSXI6MNbF
Ej7PkOpmJ+HZycAshbj5ulldOpDA0oHgJswHs59PxyCV+yXRe9knx/9BlIm1sz1y
CJ4KHD0oNknz67Gw7fc3S5/orgZgTiDKlnXPDitgkizk0y4DeHESDt2Fv4t5c5Rm
`protect END_PROTECTED
