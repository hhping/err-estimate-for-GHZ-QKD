`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pODBZ5UsTK9/EYauWJWJlDajKmPzFySCzbOs7YMQqrgOUzAFrBteWr8WzNPjfFNM
g7BYaw33iJqm2sxi9YKBVt3za7iu4S37m2OQBe50Bqt2h3LJXHgOv3izBbopv6rI
CGRuciGCJ7aJeqYKqI/VKzMMcfw0dtuX4FnN3w9U1K1Zs1BosqEhcsHwwpb9mO0Q
lAyBdJJprTSeY2pFrb5LaWHNDawvA0rcCivCDokJ+4S1RWSKLTymSUHJouGvjehS
034w63SlkyhPAgYeUAZElDDijZ0m664OK1kQQlzoduywMJVkmI9WLfUJ2pDHbi6r
COUvT0vTZDYE1HK5SkhX/gHBeSIiIyqnFJpsHLpn+nseKCoVekBr+3X5WS/SDzqm
v+hC0oaCv/ZcKTbJH/yPM89eh83kTkKKAm+team+qQUZcVd2Uxfplr17Cu8SxJ7R
hMqSqnjPrCOBVGovCDx+CoDnqn6MDL/LOKPyqU5JXNiSZwjydrL2/AnDq1jcGuXn
Ed/5hcirFhV8ODAU96FJ0ttYcwQUEf1j7xRzMBvTKjhgM/TuOUmaR+SCzW/PisM9
yHxy6rOxESIWEe8tgiCMQsOu/010kFee9C1c6sLka2mCbRSoBUXtxvW6zNLCokUI
7ZrKYExLqgkl8v5IxjxSnnn6R85uVXzstqbdcUHbDlo+n1/LPwidmMBl4sJGNGVr
TnSyAInZWMVcXEw0jFVSnXvh1L5xdiM73Sgr609zn2hIlUpyMyJWGzONgap2FydV
HV2JhHUN3EW1GVNzmKfbcATVIxgK4Q7i+m4WPAJwKUQV5xHHyyzdmkI6bpTOX9Pm
ujeA9qZJqjDTvV5k5uen9jZy75uC/1IkPmOzCXS75ksD6rJgYcUqcCVEEEEFUExt
5J/nL0Ut+MCze7eLIayhE0luu9qHUGvIeSkbjIc3xEu9f5/zAD7M6jXMQ7TkoUyU
arY2g83VKMWhCH9LNLvDUAR6M5JUEGXFdMvubRCKxHMAH0lmWNM5hubMRv0eJY//
+fU57RaUKPQBczeS/2+6q57ec6jAAlJW5/EPcQK30q9OzBBPevBFRqqCj89vQ15s
L8ykvb9SEK0jjMCg4GaW7SeF1iLomH21jGSMR/U49EAYVRUta+SJK21+rvBh8wxH
YOCbVLq2nFQuskyp0A9gFQKWGRzcq+3UC6yCmE9AkrU86i3cH+G4aTE34QwTxwdr
djtEEEyc113tq7ITzqk71F2vLg5ddTyFu8lokXhnSHEq7k9mq111LwOP3f98NlP2
BQc/RySp7ilqpunQXW0Yj8vqT5sBL9iVEkv/q84aTZ7FwJeXY5Zka49CBcKZ6Joy
zjdlyz2nAVX+VdkStj/SvH5U+NnbBhZZZkBn+O7c9jwmQBpHKFAuVtMlnAvRfehu
RL3vutVySNFUzBnC7IuU2DEYDchYChfk6ub8HBy3uBDiKWttdOwUpFvM1zWUKt2l
4zPjtjQSDKFKlccofLLe6CLjgvWNxRhXQHm2axP1yIgxILZeUgLMHGGWdebu8jui
0pI4xGfD6ozyvd4eOwsKcQ5h5ARQHLSkqGmrcQFjm76PqfVPCcmLKTMFr6QlaYXH
Zj/yY4H4XrE1OBktQL1P8j1bs/1hpfPSXmf5wgg9wXdPqvsLNa/asBTB9XRlTB7V
jk9RIYVfmMmCWiC72RSSNBGddmK5y5Xe/6cM+3M+YISeOtdwxmakHMCGCdIAIdix
gj8ZeWMeNNpJOgs6e+f3FG+wPDssOnRsTndVu5MoZBVCcGwM1klNVzPRe2rKm2le
qHPb3AsMwyFrtHJ/c1KvBh2IEXum2p3Ia5Z7xBdx9se6XS6f/68MpgXKeFWYeZEi
l7x2SBiPcM1Ap6U9e36i8unoUq9VtAy53ZRILLzS1043Gyi23JBlv7sUe6hg5f/c
3lS5SCAuj7RPgPTph+LOJXO3aiMPYIRQD/a/jPuJw3/ZsS/Oe67l+KtV3fvfe8e9
oJCFCstwbHxvvqSGilxW5CCnCrnMDrjFiWS8lhnx2PKpJD2rR4fBZHr8zpxuu2H4
VbxBHHFS345liVM7VHOczt5W21dh2R0F92ODY9YNNFBrbBHPx2nqWfAhVuKo48Ry
2b+Vdkz25pPAq15mZpkHsXG03cHl/pnT1KeWqCvEoUfB8nChhqjVp4c79G9JAGLl
WYYNISE+ap922/n96bH5QbgEDpixUkpngh+4E2OCwYZe85cvFWqAo+wlb3yygFxc
317fDGwUz04wb9ts9lM9ZwW4wF1aqNaWCqJLRa5/bSce/0IPDMrcs7Z1oToAqm4G
4pxysPW7ObopDJx8qkKl9kaXqXhrmFzPr2p7PRr7pqtyQPB57ames3O86EW6pAIj
fedzX463U4JMU/LO/7ULu6TcAVThWKDbv3TdqAFZ7QNZrqgStXxdspz9KAUyff7L
DRr+TdSsGS9kQ3E0xtXLtqqw63+niDppoKYEUfjSuL+5pRGzB55A1oM/8rT1JLxj
x6JXY5Rw8gtG0oNxJeLp7TXyg7QIztBKw1Rig6svm23A2lINwqJZs7W2IxeUTOpl
Ke5JIQyW+2uO+2DsEGqg1bfS9w+p/LklQWrZ0vw/eiuKX1lRnJG4q94I3qDj8156
9aLqmEwvKbUFJJlfj61shT5FX4b/NBkYdyDBdULXLP+mCSIdm0lJf+KJHtSWJ8ey
GNvlMz5563EFD09Ze5uOjWEM5SKGAnl2xyRqvuaTcI5lExkrW1A6xOPXJwppERWT
tu4PhICj+paVp4BmXCJIyOq0Z0k7CCC4g98vQwGnIPjazVkoNwrD6m4vmr3YNAmc
sSShxGs7otWtbqS7nakS+F0n5N4a+ZKomxMQI7XVpTAK8cpnJg3/fmygwtlmqYXE
DkDDfYpwemRpGTxvYZcg3TxgSDwVa1jesJFsxlzP1sDz4bWPE0qFcuI943WrPljt
fEJLxXcLPIDFAxXl/8Sj4Xo9svW9wpqkLhGI/xV0CjgAzMIlZhdJ3t12tFpRQfFG
XMqa8iPmU4uCJR/SHcbVYFG+DmMON6wgIhyDthjQYGE+v8W/YFtfVPz2Okz16N8z
hKuVI1E4dlxfmlnqiqURV327RQQxpiQCcNyCBNrJk8annZJWABOR00/TPtmW2SSv
8iODnTxPSLsjEYbCJiNhVZfBHmVvY2Acd3a4IrUeLSeWv4GFpcjSxx8aCBEaZLOV
nfBqIXkbFGAIy9nTWgusToxf8DiHNdmsR2Gswm0rsAF+L4F+BX4v/KVUT1scVk+Q
XC78qO34ynD+GhV4NCBHhc5L2QKtX7r7gHjhMJdpHT/fgJKkRSfJpCVIN4inedFz
U6bJTsr2XsTxaXkRdY/RZyWwWpTXNyfaAtKQB7CayN81m/cMyPpPYNS9Xjtz6fx5
VNjZsonrzARmgx1kOIUv3GkkT4CHt5j6B23gfEN3Ta4l3lSuJADjH8m22xnHH2bt
hEMESky8txQji/aI/VnONFKPAUho0lw8aKDn5Q3yD537dm0ni7TV6+qju7XK2qdd
dd+xnUE7fiqBjbLui5gj2bL9pYn/gPF0GV81dAOwMch0xCuFs9BK0my+B41LO5Tu
8Dxx/gUxlkuyf7HCQoEDQXK4ef/XL6W5KOG1IF+A4dAii2iIRb1UwXKd77M2EseO
5O3yRItuwkE4uQMDkm2PMNXag/uw1Y8bPUI/jsNOUkQNbPcok2O3dyjARk9m7GJL
G20MapairGmguzcjUhcnaOP9+8vYoGl+3/nkqLeZrDfUC9eURD9fz6P/ZjTcQgQg
AloSd4AmoWQcvR5fYa/cIn6Y62KORfooyy3j0gDPhmLfd0QueR1hJ5N/GUEHkdaC
HtnN54HctF9jfIjqfASAieg4Og1yRBKjvy0Lh33hfjNiQGI28pld84XV8IT9zAkM
sTWVNFreJJIceK1kgFNMZAbxGAs6cIWvg6HarCkZQfdfY3vyB/e9A3vHbrotFUFb
tvOb9ybjuxRZQYZGZ7weC69qqmHoRH53uC+cM0TS7e0afKHl86gD08Xm5JSY/Xq6
0LsVsz/Do+auC0UBX+qyfabfAt3PqOu8xGxVi9VtB+OWY65JD6JAMjPeH8qK460q
p5bS7DJNV+3vg00LbIdnIDNAzyzBpAwXjwoJnZRK4jfYkZ/+dHgq+RTwagStDFQH
5P1rNZR70ALiVc+bTBpFNYvq1nXRtAUOBOYDREjGzeCLh6UqvWRVp6aK4/gD4UTy
x58WNz9QeRdRHamj6eDGPabkF6prSjpt+my9P/8E/+xF6rXWTtB8Jtl3aW4xOsAm
Po9CWduMErayrBsakpfwaao2moQPMQwXlHwG/B0MfdIkdg4zkgQ3mZzuK83lwIsY
yHVC+rWMenLr6P/QMfMiifLUjMMDs3qGO8JfuF+/XafOp9kFZ/wEF1sCnQ2C5LId
vEms/dr509IunC4btYaOlACY6OO6BmqwaFJmPbd1JCvfX27Wn8tcgJXdcEzU0T/1
y/+Op0W7xMwEEuIWEwEBe+REqZXuAzUrusQedf1MafRvEl80JXcL/2yXo6YdPIPT
/j5UTCsU8ZyCNDnILqbVoXtkDAjO9+ggr1EHjsXv2KV5ipMPBtBcrEb3ZjskcVSN
2NTdu3G+GpwwljtsPBYRzxtEaIYt9vQrZYIB+WtXpAMyQ5h5JByQzGq3DvIJ2i0y
1spMthcgDgyEDnhyCFM9RXf6cW0XJIMDMzDLfEm4qhhs93RW+pld0HrBGeaDMq0X
B+EbZOJ/JUwA3hW+xULZsc9J3/NyFrqZDfrH7LNKXG3jURj20FzXTwywCVdNjT4N
4Wd1MU+FlVV7nOChIwkVVDrufG2ee9xnHXGggHl0Y2Fp699R+AKrkvfiBoYMx8um
S89SP7qWmLwOpLnBOhmblHq75aPOuHKgt3uJLEdCO5jkZvKE2hEq1IGdpXz6zNTB
01UjSM4HYCU3YrD3UZhdyEhsOkB68W2eLaGvroxRqnuTg1y4KWFXPR16EomoeP33
kz9dt29EQpsFXk/oAvFuTNy32N0X4R9KOJWnni8nIbCIhKpgloq+wZpCFllP/O0k
RpuXWdnHWUxzlJljdppYopu122CVCxwwep5qIG9XJ011l+ChpGGDU7kKgU+fBcIE
RmukLs5L19EQrkULXMfX1HQBrtyuVxeFrQrhsNEKBy+HCBNkpvdvvfwdkxLD9xEb
q82lH56zSs2k6CWXpWC5hC9gYTYkE+VEL24Dj0f0IR9ux00uwcciJSpM/JBaleb4
CEjvnKk3KSO42tgtMUhleQ/uUSFerVKm16MYGfjCmUBKPGGRQ+fyzmYaGNKEopvo
E+c7k4+V2jE4kkDLAUO5RGFYF8nNXMfuCZ1O0xkm0knpctwt8DSWa1AKfczNDcdx
2qidtSwTjZ/XwYCYQbq8Yz1yA28ZKyzPBueVz0N600tcUcjOfBqqgrB5U1JaG6Wm
0kHqqTB05h1j9GvX6VndVfmaT0KAx0jNPjQ7e75ZCK/3zzf7mc59a6Z1f8tsPBJx
S4IkrjWqQ/eNDuZZW67gc2RmE7ERjMEK10k7QbjsPkyQthhT2Wtcv/rEeehYhNgX
oSXtqge8vP0mNe6/37vYixCxtdFhRtRAiCcoXCMiomamz0a7QX+7tViYzhgYC1ZO
0QDZIiGAEwJ74u2SRnsBlP9KBflrtx4KTnP1Go8fxqpU5PYuH8/kqoyY4zphtXlU
UaZWXEZwgmPXjShjkqEizNP8Y59kOs4PmC6I5JrWfqu1Ik1icQKCl+9vxVxyZ/qo
okNZE/7v90eH44Cmj15JUJu4GFQRsHi9s5Gbjh376h3JzprSUvZM7/gKWTcRCVzM
xu+sIiLLQewpgr3XEHeF9FVdZrasCVbuxhcu0QsvxuyMIOmfm9Ni7qYqZLBzHHVr
WpexmVQchvkzilje7Egm5tFuDhxEC1NEUkT/9D82OIS98pPMLAhmSvSSRkKA7I7L
DWr/SBjpGYRlJiMDcN/lvmNOn8xGMvluGjLh1ZwW1RQi7rNn0PJBVxtb+6w0YfGg
cpzEEOUoxKPbUclQ7ITwjbFv/HQvcilICXKKG/+XMAOoSTqvNyU1AC4CTdjjZr/p
+pJeXcnv8ZGmWKkdeG395kwx6K3I/RseW9736EY89/lGOCl+F7Z8FctY0tKsSNfN
o0qDMJcG50e2wgqpZ8p6Aef+wO0NYk2+ak51aoU2w/6uVkkjyyKeSEyZIvSepCtP
u24iHU1T3lKpgnxVih89LoYmnDRmyBTrJn+u8IcmDLyOXnN64m5C0c5c0n8iT7FX
kTwLQCR2VudQKkP3nghhRL5igzt3iQ8uKbBTJns2rafDcPzo5ldRQzxsrKxeUwyt
0aOo9gThMqC8niFjJ9/gbA0Oz6o6DBOpszhzaJ4pYWUSubKePPz3tLSpV9z7wIoA
Fc/Y6hdrirbcaIol0YxhefPXYJTp8s6zD0SjqRCqSfnR14FSKBoczjdSnwplrySh
HdOUH09rzKKeAHqa+aAQ/I+6pltfHCpytM72Ph6mkgbk/8QCt8v7vbQ2MVWNBfCu
A9rdmrcET2UNo4W0eSqgTQUUcsMI6yVYElLYIkckOOu9eVu9fGJOyt7bj7v/a1sd
JEc6iywstGV5npFyYW1xKdp2CisOVsZ+koGM6WaYhiRveg6VHMiqR3Pw2NITt2sj
nm3YqLKAm2ZSSRoHRi50vIGUiWFNjmwK+WibNdx8DyOaZMO/hDFjylUGwqYWL89V
QXqwunLcN9QTaSCOfahvh2shgH6whBusgM+V9EUoDbuINDJXnxHOt4KTT5YGX/iq
YMo0kI15HYT3Oh9/9sh12F+xmi5TMetiMGJViSf0bWbyrgwhV0ByDBAmtN4/rSoU
t1jqTK6Z2F2+UUWjTJ4QAmGc6RmyVgULjUdAIX8R2YgaC//59XwDCo/N5X+ZpdKt
ETdpzr1iFu1XfopvhlO+D2heIP2PuKrRP9lJ7At3aVyJ7DFTXN/RcO1DnSvNdpVe
gfmcCW7PiO7Pppm0QBU69cLzWucjNo4lQhCqn41cMkI56Qpm92RWpFtbSOev7P/t
nfaZkZvRo4a1Fq4NO3XpBT6FYIofe4yCeZByFwHR3oCtUeHwnyD2Dh/juBGImdm+
9JXjMmsOIFt79aKWcNsb1eyqYQKjwdKz6hiV4w2n+Jfy1yX20WQW/fe2jfXv7QSS
O9iwaNjUcsVYmaMg4aghD9/IBtDaCtM9kcZ1EnG/BZDFIsMUbDhep2voR9EUxD9h
o2Mi27dYLk0QBuOLCXDUfuE+bTdOTERo3ESIVEwFcaIjDaqWFMRQh8V+ta6FNQZl
oGhAva8/kBmjwTOqAkFioU3oCIDXYMqmz7poLGttXdyxDDkkXzFdwL+OKSIDLS3P
hqcleFw4207go4okyXLn98IN63zzRD5lJW2w9j8CP9HABLyJuzSkxqgX9MdWjiVR
H5xJpAes6wTVvxN5dTh1AEDamS5LevGPJ1lNQu1ghg+f6j5d8Q6SMi8pZALA4+MB
8m4xF9+/5BoCI31DWeMNjcnahplS7cQoLFUF8nDt78I7ch5aCI8SHWYv4kkszdNJ
N7dTbCf+DW+xvvP+WUIW71QeFdiApRoLyyeSH9sePfyGPZy9i75OdqzDuLjpx7Mx
1NKVZIK5lUO9r75//3nuKjuENzHTBtjvqK5RhLw8tmkLufOQYSnh2tRcoVL0Itts
p+Mirop4MfZ3TxVwNKJQAeuC3YmWZwbu6IVqkkLDQSEzh8RzGF5yOyIQR9mc6PL0
4xvMW0r0Y1hbs4+b8R6qmsPR4D5hT0l0g1SfgWDSr58Jsh3Q6TY/UufEbP2uac1T
O/H/U6+bYj7sHrzBDJfLR9sbjqkb1aL5c3YykkeD8kq0xpWo7KnrhzRySQ634mL3
48+aSnLMnTZ8hLs48rljPiEH7slP661R00/zC3y/c0PtIhH7RUfYjS8Uv7KQhlIC
UlTtVq2CSUjdyrGtGtHZ+EfdHBdkXC1rznsU9KyjMyeuP/CXtnXuUDo1+u5gjrPT
twVDkoP5E9GaJtBVV343d3bV8c26WbV6ypU1PegRmDJkQ7qyrM7BGQEk1/LU5ak+
YUQrCrSZPceTnTPHFBeueHwoCuw0vrV6p7WZ8Bv9/2Ht0JayQJoC0rahIZPELB0J
xLBv10r0AFLZPUqxZknm8+uRroGvUKgHYQ7tdgA2RPmhRChRz6MGU4pFRHvyGBk+
EPiRhWJcs4k/Pg49Jl0Eese8t8M5Bknvjh9vTZE0ns60lOD/qA8C8yIDp7pzy/Xy
MNZf1XdldHyTewjoWw7d3GnmVuSPcEZlqUPfujv+2lod6vWJ2X4fM4iwCY0NRNUR
XC19Tt/xh4yvL77pQ5Fh3eGEWSk9I1pfV83zY1uLFzvYRUPBeuF8OZDWa+3tru2A
aSgHcJGKEHU/HJtLqda3b9ED/ef4HDnRpTimSa6SSPXnbLpYx15LEPbvpQf97URg
1QS3kOu9N0I3e1/s9t3JeG0DLQEBY6+IA5SerKVnvdBujCsB54Z2tO0YEp3Gqk6K
eSIUNtJV0KuB7bqUNIz+ZcoACSFJszDnJbyo6BMTxm+UX0TVLt0V5fpWBdj8hEY5
Q7Cjuq9cp0nTWvZisBFxa0FG5FJlzlg35tScAse+e1QiRgato0rXnJJu2aRGBlo/
1JAVqT+MfxoIV/TCuWOAPZzl4Lu34kZ10dcOX1wza9AW0IYmWK/OUqMkVgYh1nJv
HvsE7zJ9DKWY/rMX7Fp2RDwvbZbYisTOLoSy1wVncB3qUpclfsfSwKIi5YBSdcUs
QCPfZ4maQPNjkOzDLlWKslqFLkHEOXoOHfK5Saylbcq7VgeNetILHSn9IDvSrgXu
yclcQ1a2e/tRupVDXMC13c5DiMjy7DNWpMjCirqdSEdJvklW+D1W3QCSx+R3wlGX
a+v/NZfbVyohaS6MqY6fHknw6YJRpBhVKe+Tuc6wl4xOKmKIMG36xKQ5HovYU6YF
sV0EKv5FqUa75phwyVtV5L6LTkYF16LqSqSxga6SlERy5ai9JndQrSTmilBfqvp6
wHcpiFGpr8/4Vxm+qQHk0ZjvJRU5UmYiHWWHDl8KQ50VK4x8bPjXRBlFKlCj7GwR
pXlerJ9ZstopwDnQbGql7H/J4HeReC07Cy2zvjnmeQzLdl+B1sKwFnPE6DvdcpA8
NIxJSPPMcq4roCG8IPpVHcj5Al9DhHYj1p+6wBXTeZQBSCVKvx2boJnjWrTGHEPG
6TBKIg2/nT6n1SzvKeBMwMV3zcX5SosuSVGt2ETePK5S3vjdMiVCdb5w0ZLGU+yR
dSQxodIIVHPbLNWE6E47n6TzPrUdVfHGEWUYAfxB64Gd1NNT8D6SHsL6HTFnOjQh
fOTfuxNqt3ol8VtIt2HCe3AQcvdX40n8AkucBar2BEftat8R+3UNVUm+obQ3VGS8
eEzRfe5sgUfc5ve+VO4KKW63WbMuF4rffsTTvmHLHlttQWMMIYqih1rmVkbq4D+Z
HczhUMVSej+ds/e1PjaL1zu/P+zll3dH7r7mwg1YUMckRkMKkc7/CcCZ5XYVbP8O
CAJ/8zMs+ha2ETZ1yEmKvNBVkCVat4O9qV4RCeqlSmLBPAc/aPLIJCHjj9LdRp2j
wz2fjeuNvJodElDFxKlr8cNWRAme4vGzyO1rkDFp6Qt9R2rSXDPLPdweKLbT6hV1
pQSyrsewhQh2rP7TuB8b02oIbYX1ZFHB2iosTOmkOT/zr2dZzO9B/80FN5+Ud/S2
tP4WNnUyxbPV69M4P9ljZQZinuzHCKhdcKv/YiiUZTmNGFHPuu1I81vIUhWjptv/
yA/Tw4AeWLUe73HVYEM7u/f/4Cf7MQS/e5AHn6YUnwYAKYhEhxioE7xidDbYfwmL
MToW0i1I5ZW2sfR7439XpP7YQRFxVzjTieUJtCWC8QyXhJ2X6CB9SUH3ippGE0KG
gG7a96zNfw64CGckeQzupl8kS3U1MumW4Z3kRhoSrOEQjQda/EzDt5DdwZ3Z0i9D
FWAl+K+ZqO6IsULJx8VuMDB++h3kwJmAgnYEpoRyBWue6RroolXRbCoN5NN5fCra
N+kElpQAPATD0I9s2rBARQRoA9c2rjnvqicYjCVdOUadRy0LrmuC5p5dRfqNriJI
0bfQjqQK4g6ecH0s7Q6MBJXEn6/9qJ7vDvfBCzD4PlMrAyrbHU/JXwbwnjjpbLHY
gEtj+1SCkq9IlDDQ38SBnJUfiIj7XMeYWjNsXhJGVQbMr0Z4ZLYROrgqGBYyqRUL
wJTqNnx/41iY/z2IaBOyfGyOh7zZuIv4nRP1fG7S8/Mr7yPZpsp/l9OJ1kddr3dz
mLZH2LDArnAI37PE5EBHt58i5OslZODKh4LopqfAfmHNHzSkQZnyT8pncQ1lFyIi
Z2a2iwqJXmUTk0r/T03HhUJFM/swLwmaVLfEmMZbHNXeU78h85239MHn0GcPZ/cy
S2bMCyhg1thiaMmL6yNU9Pw3DwB8DM4fi/V10nC410idmBbt63dHyXV2FToBwfN1
W4CuybmBI6SA24WyWJaToc/4s89KVZTuKJhn3KPPC+VhqlqJbzYEA25egTvzXo3v
a7NuMjYfIO2Xj8guwezrHglhqsrlvZQL6B2kS/Njbtu708aBPNyE2GWyEdEU3w3T
dwqJ7oT34qsx3W5abGm9GkW3usPbR/FBVkiSsjmhVB4uqOKe/k4aCqFNnRl+spfF
IAsCOlSewEAoOnY4WyZ3mY192Tu/8spvs2cJXfdv2Z8+ofdF0CO+DNSltb8PZ4cJ
p0FaD2d8YERz1UE9mx1CUkW2y5rTBbNQdSZuNv2GXvqXtZI30UVQ4MdwEvwdQjx+
15KtDO5aDHwbAilFsb+75YRZXxUDjSLGdBPvHczgEi0BvrdKI6bGdcDRCf4lgaZw
z80WFKYCDyg4ErazICyGIsLSsVEyhU29pkAKX6y3zm6oGYEPxkvkdpbqAcWEOeEL
WBh0UCj2n4h1dPXirWIjVLbpp5zV7mCNyIr02YGN+F1SU0uEnxXaqW5jgz04xySe
NHrD8WRdeuU7MkqcUBI903oOjhxy0+Ygw5W1FBWKUuMjy5SefY8+67Liewfi+e24
bsZ/sZF+gt2zBajzc3Nr95XXT6e+o9Lz01DhvnKiayD1dOejJSGmFxfzriK9vpuk
YBNypm2si6khuiFFL/8Yu6vnA9yxyGchdf0QSwbrG64+XqtjInZ9QOVwudcRUXOI
gpxkd+Nm3BtGBoeXEz0rlBoTX3S3m9WrmW+zOOognyNF9vKFB0QI/9ob/xVEeu4q
fgGkQe5KN8a68zp82XD1cLNAtPScAJi3OHoKF+22o/WybxeWVyFlT/I6Q4ZckHVR
KItI03ZuqG9QooBzzqKFPRi9bjdPsQinvVoSOgym6KTTRQ75NGAOUdD65Lr4MM/j
9aPt/vQ+Ane8qZHWeeKGr93veIkAsb9VHBZOVqwVhajnSZSo8QVxXpP3Q9Xf4a0I
hdHk4krK9/JKVEf3oWwEZtV187spYXE8cTUyAC4mwQulUfB3LsCrXaWYK0TDvPDN
daTYXeHmDB5+V3UHl0thcXsNy8S+RxVke6O9UJm6H124X/xylsIx9R0P4zSR0SE4
ABbTERziDeLptkwAYl1e0fHLH1iBQZSzPJENpEf1oj7JDgW8H5N8ZPx9Z6yQvhxa
tUgnFP5EpoPzJ8jdzgbTGGKE9pUzBLR0HxNkvXVwey7tkW4HkUrAHrVSb9lAFMoM
+i1qlBkVBAujfkK6QcB87kFkVmv4T8Oc5Tqtnj3py/TDjdUghFd7T7Nn7l9Iis61
e3ERpiVIITGbA72w/SQhlCg/p6qM/mTBoY9xg+spSLaJjwxWjGxR+Mt0vDSh/6VH
UEh7Q/xv3GUJ+dhCQuiE8aEIAGkkVy2aWF5eC2uy4EKF1EevNLu1d6XeGVpBM2iF
J1+Pco3fhhmQILtUzwAs4TdXOq6Ka2ntkB2iQKkmnlb2y1YvItBtWOa7tIvl/xYF
FDPIX/FoSJT1hIpEZ8zE/irXIjlO7OI/wgZD/7tOKBvVPsEwXW91GN+uFsfQmhSS
AGeV0RGV0SCMZmHpaI+zF1a6Ta0AUAKsDd4Tv+LuSk3r672cMrukOixBaPQm8KSU
2bvvy0/47EfE1Dw0nmrmazzsWCGvov+kiOe3eDvuWFRVuIvBeJyI4VcIioR9ufDJ
bGnpXPgpVXwWYlNlaNow3NJdLEzycnZh4EPtzNvnFIX1aQWtH9U4Z2yY9nlNr85x
gCE6GhpOov/JcwIsMQnueAzH3K1bm17Tm2FRll6X6Ss3U+OsND3ER7l0PWF2sdRC
CCHeHrBhXpbfoKWmYfk2/bBw6qmF+w13mowqcTG2xy6hxHpWvzdcXhsLL8Dx3eqT
b8Bdq4a00Q3JBD3I19f8fMEAtnYiQVqRsS7Nw3k7iIp2n4pkvV/qu7JbF1JqbO3j
nDyVvy1zahJAgjq02ONtYunDqr6l7atxUluZ7JCLCbGNxmr+soaZH8Slv7BT40ZM
btUfGQzOqJLmXTDMcO/4UYXc7cr3IzogpN4c6KDtCnHw/68PxUR/Woxq6WFkxROr
SPHsY/tpnLMIDDFTRvButq6tQcPiTgZoRVmH3fqWBCrL1VVAsnox63xumllCa3PT
b39TfDESs640UaFhf/JoCx+lE5AHynUH5K9ycuT7BwMgsqCkSjixErzpeLhAgz1D
N0mGORfSuFwM1J2e9zaTFpiN/+VXCpjJPR6oEMhZ3zz3AymVhe9UYxSvTt0ycxGv
YiFTTuCqE2mca5y4EnSOG4zfHOU/HERJv74wZ8B0Dp+o568SBdBKy2tDZBwhw6PD
J2CpymRanTsLJhH2OL7hjmAoE+ShTtiBZYwjWoG/oNbwN37aRK4GFxR6sPFNRbgb
8vib+05gQ88VIe0N0cRrD+gYSD5taG1B/OSvW5i9HxR8gRZ/ImhhtsPLszJ5zpbm
S2OXViBXVlXq9j+yHedz5uy56Zisjmx8SvUPWVmvMcibbhKZMst1Iz86A2UV1q0v
hqAVr7aIit0aWnTnp8RjnvJare/oE00PvqibeM5CoWypvrwkX8lLJ5TzB4SGE0xA
0CjYBj83dy2OCK4oDSSiQfNwG2htcbBdDrRvL+HZs0FEUcdOuxjo+qK7XhkccuGN
rdngjk1dcM2qlb8kF7ic7XgNrmy4zMOkGwGUpfcKxEgITqWr4/6f5ucMGisaT+V1
arPKpXhv6F4tQLTNj4AgTnGCedAl5vrr9flvMFayVOQf+RWi1FAd5ls5B/h1EKB5
BuHiL1f+3Bz7paeGz1vtkFfj64ibHsAK1xPd5jTsIK/NalUyYVuNnW2omvbRTX9R
ESyT9YJ9jTJcaYxw2h2vT0NJF3rUOAWj1+3pHGuWEgCUX95/pxkGu8sUDfUTy/a7
jXnWobP4UFi4rGe9NhnEw5+NgSU4FURjmDqtMYnjvmLmN8UWACgJM6FAWREV6XDv
/RP2sSvjCamaL5ZZrZ9/yWqDEdBsuH6ME0OyMj4hOqPNIxbx39nHC7b2xhA5JTjU
L+HBOpF2vxBPo12eFu/bpUMtCqO96IpTPXlaPvegHxMrvee5dHzCFpSWVznS46jv
JAMRJERSjI3lH/O3wrF4H7WAXkllMCsY1KPTY9ePmEAeI2mRqh7oW3qLagOy+AsV
J2LSWCrJEhZr4Z4iKIB25rOLjdybRZ45sN3Ko3Ir7q/ZHvZGM70iTdozh6dUFyHE
HOgGwh+BdVsTZpTX5D1btGmnRuoLNiUiOTFWwpRtqbczgXMenXyCM8OeUnoro8mj
uBCRYqztF7Uci9w8Q3MiY7BelvFBDThatv41rg+4JnlZEDeSDnHM7PluZ2yE/0XH
4OLDGDIce73pzJxSGa9qUYTnox6pzw9gU//iBDTbjhdHvJBuHtBA0oxDVoqvFBjO
c8PrNjR7GQ90m5mzq6iDnc6XZAB4/3TFH/Q5ZyI8vBP7oNI7oci1NQeyDtzKqXIx
hSHnJlNcfIxeA3FUA2bsTAG1Yirgz0cblokniohB980MUQEtJdNxQhydegKOXtZE
QgR2RIvpLkkLnm78ciErblsmlDb6gsXOTJUjUxiPJp+GYz7oFWjcO//zC+fsZeMZ
1PjAkiN246ow5esI9e7Alg09+U4qry3bzAVlGTVcc5xS9j2yvUBmzwjUSVy6A9j6
lWgpsGjX6x/jPTOtVK5q/+BIWLXBpeWZlBSzFU22IuUQnf/FPAM4SiY2Qv58dyN2
YjFywk20cIOk8b6LrPyD4d700gCy3zGVmZgxCl/xKtkcX+Ry7E9tKVDfS/tMhBrz
qVOY92xJnFzHyZ8nAM2EqhR5LnnWqVb6eqnh9w6jrojrw9RHlAQdvEdfQT6uBT/5
JoE7kJfrsVhvJvppna6VQhbvCsm0KuHEEADqPJ6oWvhR9MM4tNRvPyhIFSdTfY9o
FIBMZuAJcV7F2Cbfra4COpieEaLO8DuMAAd8yYN41h/T2NAdfOMKZa1upJ/BABz3
gwGyPTjmJzkfjWmokLbppmWfMfB6YkWEDVhW2awqUGt//RUmuOsUUB3B8l/+Lgjk
qrbDP/Yl+TvCKlOu6GgUQzaHef6rgqzttE6JGRw7ey2NuI3DfbVTqcnuLPuEJj45
ZXDYHv4VuZEKK5ZrmHjOTr6ciyaWXSrsEbuWdTG3bHDjH4nSA2FD5il/Mg3QuBSO
cEwKbdBpSrOuaoGpBn+ID7s0kuB0/FgAKmaTbrTHB+d6tFXbqUWJRu22YKhWNsfv
iFNadMSTA2q5k7XzJkyfHV0BltyZKg0mQ784XHuiLfY6zQZkoMM9Vd9v5xrQ6CKD
nuVt6GJ16Um3Bds3tHhi1+4hq/xtQYRsA/62WV+kWHUnkpQqXbp+qcz4EoL9zAsM
JfH9MhuQLVUY6cnmP47KpzhcRMmjIDpYPxLM/iJng4VZYNW/qoH8JBT+IDlnzW9+
NArsmpp1sfi4aG7E9XWSZcXu6KZGLsyjZN6HW5rlSZz2g0w69GOoe9I/SbT6vIKu
VGA9ox49x4gY6WxGDy4kUb4Y+dfLHZHclrKXvZB0SE2lJQdHNNVfhVLQN7T658PJ
uic6dyB5F2PZPhOw1yDRoYT8gjHEhyIEnXxHcFkr9XBSDTmzWRaawqRYFFS8EnAP
YCTrMKRujw80P3mqvwQUhp+I+KIyCxDIHTX0OkuuKP/I5QCWVEPu7HqR5cD0/2WY
nL/akuvkJBqY2SqQh3dc68ElT4KRe3jUzjES1ASDb7+GLeDXwulllrGWfGMpdr0W
OK3qZ3RXEISp3JXrBTLNZ64DL4iN1RyF+k5V3iE0Kvkwq7Dbul3OPLTSqL9B4LCq
hM66H9MQvtsqkdw5uOd3jhpZOso9DKPMA0Zy4+HgTNZPLswWW5EB0Zf/4Uj4nT7W
/BU1d3k+DwaIijYObVN0jxcQoRUMiK5DXsLacadpKeeLgpKyMgVRJkJdfpKG+Pyh
PdJ2Sej24i+fkQFGZnKBgGTLrTt34+2M05yjhseJtdF3Z4VH49bioHx9AUPrnC5i
c/XdHr5I8XLqACfHDCGBvRGjFkQmZep4YLgeHfGbr96fecykcPsIvsv2kZcwgfcr
GlLmT5+PQCf9mDDJwsR8wcCJqLFqouEcShYVNeXf8fEUtSFVqmyTzf1xe/DaB0Jq
AwisUjqF7SL60sqoefLkR4e3P46tf8D3ZkoYjkQ2goSmbT0myHygSWSD9bv8BhDv
HCG+S2RQjlKfBt+futBVdie6eAwr16r8H1i9YbqEr/KvdO3AIG1pC1R9Ig5oDqAj
XqHU7Q3o7Ec4HAnJydVyxeAz797umo7Y4HWyhv4UCtlDnQghYhyIOgmNvLQB5QPO
WhdYJiUeGJ+ms9R+t6CHpXDOIIPtMbSk/jtQ1tcG+6HMhfjUTwYQ2sDb5mW0GxHK
voUo7UK8pfDMdLoeQKSLuUc4/qB4ptGlWVhfWs8JHZQGUuqOxKDkiBChGN1LCv2g
P+GcFoCh1WYAPwbfyAHL2Vw1Ssmv1NxwFSf7ZUCZl7lyHv4NSWEdKoe7MXLHZugz
Noej2cOiSkYXszk9j9efrWyT7U2y1duSYabNmycrCuANB6NNxcRnjDHz5/zdOw7c
Z8EKMdko97+AL+iGZcjXamvzE3RLmEp+Yl/iTF96pipivJxtvZIRB0POEPvzKVPd
lF5MdJH1tooXgczjKyuCgmUdz1oELxqedR4rhWzIUWQ7K4IT7ILCr8qP2n+N7YiU
bQG5QlwoxTsSNuS/JR5drA4ZjDJY5pmi/BqPHtyJaoBlMETH0BriYo9iyfBRFAb5
U3q5Vruwlwt+C1vXbghK7g9EeZX+dGFkA8y9mKGa+EQzYhfECKdKC/yM8XA5JLi0
eeNKhUkkVEL8GqHrC82hhmLXe1tBAOUY4HkpSfHJjuCmlyJWJHj9dvF/9ZD2L8Zi
mdT3DghIT6xB/OEaCyP9dAu3xDpDGal+F7hiWpUnUgN7PaC1Zy/HhQ/rcqtsuXWk
e7uUUVRreU9VB/sm949ZKBiTAhXGNXupubJqMxs54Z6osybUknYCDbkdilOIb6ME
vW0IvmJTIe990A9B+DFN2O2FFY5dG3ROm4EqLFb0NrzpRMcrpoDZLNS0kC1/TD1X
Ewzq71CIU8SZlK9jyMyBvmojscdbllwZfMXJIyBp5HMvhQaPM19vrfFYSDkiupbo
yVkPyHorEaul8QXAt99Z/avUfYqaziq4nYwK7BATrbGYHP4zc8UvXitF/3OqCPb5
tnoP6Z3ZzELUTDqT94La3JgvwsXdd92kCHpxRs1Zyae7G3KiuZ908T7yRLTGyMe/
iqmFE3KGC7ou59iNMBzz4WLRKZ3aEouC5kBYblwsqKwwz4ELi+NrVwbCIDkPdzKy
LntfyDrChEgPXesquNcx9bG10kEzyml1NalOMLo/gCMivuw0oOCk9GvJrIhy5dl1
dWzXbi2ZyucFlwQgyOfKXFu6nLLbzqWD/6p16sb9dxnYZnYL96vpEIB+J0MH2q9Z
vyus7j/YY6ixCN6WmO1uVbrFMun3D0ayUCGoeGi+YuWBT07KrZVbQX/BmOiMVi8B
+7JY97Yi5Np2VpsM4YLsnTiHJTMktNo6kAW7/1ZFQr7nKmCx41b6sgGv/WbfECx1
zBASZIMs7wO8TsvXg3LKHhbtnkb//hD2bgmE7m5MlykNEcbHN8Fu88DiGHJap4eF
GfUnhn2JJMwZSCoA5roP+prApoEKVBvATr0jUOtthYQC5AZ/oPagHcRqx914PMgr
0qnOFlR0WvdQjRBHmrR9bfpc1nDa4d2AaUCkPUHqRTp0uOkDbbzAdrzsLu38P5kd
KZIyTJKPd/JcpNsS7M8OJH7PY5h14Y+NL27aiFna4J+A4M+ZQnW8D0Bcauch+h98
kaFvaHxAHKqHaafAgPpWeod4NOHZBu+kbxQcdXw6VWdadWyhZzWP/h7zQgIGmNXb
dGw4C5ABoJd0qbDRkc5ydSsCH0dclTMsn22wHrd4s9Bma9zIODdUqTiM1SHUxcmf
ZQesMXX4EypBv+XhhiSPpkRGg6qGehO7B20TJKt4vtuufa12MpxY8WSWgzkEQsnc
uPsS/VAsuVnrvBPx1nXN8/vhlNc97fuGWFn+wOVZfLHpjCgJSwBRFbEPgyWFjBfC
LRMls2lFzZojbSWsE6zSoRTp0wYyfdR/J+1sXf3el8FzeXuaf63lQj1Wv12/L9wi
Z7RmPqDD8eX7PFCsG2ia5jELUI66LtjcP0ss9nEgtyQa+5QKIeiYCUiGe/GoX2Af
3T00P7+QbkNyXaNvJhbdLW3coFzVmlWt9AmA5KEWMZAnnnUtAzekBVSyihaB6jTN
zFW++y9gPfQA3bFFxIQQdaGalb73urJ/H/l7+zZIejZW+/Kb9DaFjco6ouHvHdXG
1+kCjk/kIH7wfWOLk5iepeTLHynmI242Ci+NCHqu4zyqdtRsAlfq3Z2lOjFZhDij
rlNbEXGD1BlnsN8s5m74hXis2jES4ZH+KhDzmonFGoqjsJXdgJ+r6P+Avcc887G+
AO/7iqf/AYfU5kJdQT0NK2zuqTZrokancUQjgM/TKmruUUnZSZbKnrj9OISLvlcK
J02MqJPfQScd7QtSyMn5DRTSLaiAOdBLaBsDFUr0bSKB+0GmeQFXl9I8RM4eRaO5
lFn6+j9PUhcJ8eK/VZq8LjhtXuYbeKcdIRxlwGSElaD4KIx5tKHu3Bj0EFWwnkMD
gAs0kipRV2astkaESN/D8j23kmK0/QSupOTTyFJBkGoMS3vTgguDntJ5Wu7Ij8q4
pd6yBcyiUXBbM3nd+i/QnSrl0hwJeK0o7YwhGPMDn58shq77KeIdFCyTtLQEZBG0
iZNsbDxfXrxkn83BxA3gGqau4L4Wid+MAseJqcLMLxbcxmxJzn9v1FN79y5bj4Aw
0mE6b/FLmaqllnbADetQHu41B5zt6WLIF2BHyjMd3IBGNhdzdOADdEJQdPfc1Cj5
EaqSrSBekyAv3wcIGga8zy+juXASHKcvzroE9lfgC3q71uH7y8Yo8EiHF5KTCRr0
mlKSKhlXczABCHwEGqdY328Dat4GIcFqsAXwsbSv87ttsZaYNZjDTRAEy9mlLA6A
+O0WJYjtM/g1Y1cvC59WXLeYYyUgYDQVRFy1Lv6zzD6NM6Uj22oBPIwMQ/ngbj7+
WUA3z/hK79advZbYqi+NuKSEKME9gDOXP4u0ML/U67aiMwbAJQxn+xbiJzi8MY9j
a4sKkpzx5B2AAw8qVklgUv2jhKydFKIcvC7Ujg9BaSzcjpDV9cnJNglI2tVw5eYx
gXT6/4QAdNcwMmXm08ngQTNk/yPwZfc6uYCZOA+jeR4By1fI0po+Oc4REQN/VHAq
czV56TnWNlZowtfSAa0PCrnqbbMsODEGcYU4HO9XjXoY532R2A68omwfR7YoUZtx
GA+GgBo6fQRtVXjK6PH2QTSZxupzA3AzoI1EQ3m8zq4vcVYdnG8uCkWelYQhhF4R
a2fbkqkmyxYNlSAQgmdz/aooiLazmWSrU49W+V7eUhWE3P6q9KRHd5eTDajUNxYR
gEffEeyOWMWQ+PPIYvCa2qGDZPAkKeL5Ku0hv+HACB3ENOEZ7zetqXdXZ8tPS3UB
26BFrjbzBc61AoGTwFijDptTfhm2iRVqssZ+5+AzcVkfguIRNhcV8XhHDloIvfEZ
gLD0yvJd7MrUEQ760TIUN9TJ7Be0fdYd/nYSo+5p6ocB+yINycxHOBy6IdUHbm+u
pQiLggAecgL8NY4tPJ5fOWyDHIkOS9rLN1N2WLzQcloXwVYQgUx6KnlDwJaLKjxX
0tXYQdRBW5FO7WJy+vDSCJfNr6M+B6/QaQI/nTxIyj3VM+MLfddLzPpTVoWHmIMy
uYFufNJ6nlfTU91a3eZgHT3bW2s2kI47tFE4gVzbPcTZNeQAMs0a+IeqQexFsRhH
Tn6xXD1qKpgKrpBRPq8YsnC9Bz+L6dBDE0zYpmyevHoJvNj1ttUOh8qMgLX56kkd
ZCK6iTPaqJcJyfy+YuLjEY+/5C7sD1QA2lKXVfVvrFEzxpYGyjANGuNSMPGc3405
b/RPRuNvi5tPcVOtOsA3SznRSHB3z4CY2qAOKTXGlYjK4Xo4bvvMpOlEg4QwmW48
b6s7fJfZszKjFXcx+lCP39UN2fbBqHUOMhhJ24DvBTWeU5LdwJcRvk2BbKNcE4sP
qkdOmBquMXoHzA2A5oltZUZiibmShoCtqTkxVysjuHvJTyeWaXsaHUkGurU/mEpf
G0pQXSpjaINOF7SP5GiWFGKqqfGqpWLtvMAtrATQsMaNG/sXG3bPkwg1o+rWiVWv
8YFwbQaBRmV2i+Ll6oz2F2ccQncS9IrvAe7TfxDQZ6JB3qNQRkKE1rgK0G/7CYPL
5luDOIa0k6/AFcfNe9U9tk74btOouqiCLlWmhyW9qCOutOwLNeHkugCeC2us7dXi
205hqKYsnvIpmiL88QsmTsYXsezMClptOUH7HN8TDiTI5uj0wWN6oCEgKXYmCAt8
EnGmfcGyJ2pZ6RK7914gBzJpv1y1dThQCqjaN9sBuiO3A/mhB3DX0gWsmQ7EwQ9h
LueO05Za3g9L/12Fq79gbZRU/GySvTnW5+AYgTEwDq1makeyqP/B12q4MUJxpfZe
ArPJnFf7/UZiw9l9EIBhp/DidAhfjAC2fM7femMCR2ujzUzeBmmZEM611w+f23eG
b1AKnQpuexJB1xWdvf6UqijcrB5a+zr+rEmJhDLUUYVEIxx5f1imUHysS26HkEcA
boMtrtAyZ0gMkDNVrFPD23xaoE9v5Y7rYWibOjGtvG0Tn4Fjg7AU7bcD298m/3SR
BMbC+Ql9/00pei56t0qb8sDNX4ewDiLwaAM50r642aSLsQ1iE4lgEa6VazIQkzUV
ftkuPJKHde/u649Y2NzPhOueAuw+VkSg3uIZ2a7JVik6oHV87CEVDgC+URNO3mfs
pG0a9H6G9bU8O8NSzR1uxgeBGx+tuxogvuJn56vXvbjHuMimB+Dphusa/AruQfCs
cMZgaLvIqq2xOSqGE8Fz2plxoiafn2r4rwFF0VycTyWXAwj9254HWre9Gz6JSkgX
xmvhKkXwMNWcpFdzyFj7cm43bBhLvJ8FVUe7X0vCjBbrg4bHRHmX8dLVstFKs0xQ
qrOctSNOGEhvQbu5osbfdJ/RyXQFhpq0YRmbytHmzK8xm6DUXxN8ZxrKP5Pgyghv
BCrv8vJyN+oLd+udg9KmXLhZhD0hBuwac99lzmtcfJ92oS/xD+lhEt8oWRYFmGWK
oSR9pDdB/7vZ6JHqoGuIJdIPzW2Cr+ODh9CV8ypTBBNK0xu+mVECvccn5nJTUgnp
e+V77bFunb3YjoOYoPafV0PB+idJcd53t3LysnhNH/MlkZqI7COnXVpHWnklNqEP
6jPO40ZK9+/39hHrfSRAOZKzxXvTwIWAgZ5Ebr1Of45A0ylT22PZLSY02VYGFDE5
gpkSuBsTOZLOGuNya0Cu+GU0dopZqxiZwi1TyXXHEFnKUnOwuyl2vS5YJ/ShEtGB
M8+IXIpyygzG+oNQVERMrchlPu3zVbLZdY/uNgISk24mzDghyV6Z8C+hKMyG1V1g
mmIcp1hOjusoiVRt7WQGYAlStqvs3msZd690bFcQDp3yaw6ncbbcp41i3uDicruu
xXskH6lzuKHzJKmyeczdu5zLIiLUz8JKe+pfOyN4wI+ksSpxvuEf7KVzDxaJQfxO
4QoxremgGrt87CUk5McjzAWKcfsaQnSrd7Bclad0PiGnua+N9/KMMXQ0Khl9k3ak
jrfNEzhY/U6o6NK6S6/jDasJiwglAqQgH+SZbYQK5/X56WmEkogKxDDlu4U5G1vE
VTrsfhm0d97J09q5cHQBR5UNGO6eLioET4vJRi9y+sllDdli4gCd3eak7R0Q5Oi8
1FGNxoXyi7q0K1tOR3eKg0efnJG7Jh9ukXGOTm47NkxNNw60KwV7ezs1HMVlTAXC
jEphBs0/BV4tlNyJprDCgg+f1oFo1/c15zodYWHmncI7YLawljRztekXzcun6ciW
S8Gd+bJZzdP+RH5z6t6mfkgwZWArpBxE97GttEeM7VGVHgVMPY6EJ2gUEr+YP/i3
mKjJHeoJE3r/XSNF3wS2YbJKFelkq51jtKnlw32cnRyQPnpc/ofE1CA/GyesSZtX
+ffOZpq4Oeb4rsmH/GMqc2VPtArSeK1Qlfv3SOAXyijQHV7MghBXC26yG4TBlc4R
ygdeIO+ONwPEsk3LxuOoh4MXFtj8XkpPfbL3T0JEadUeK5cYGNwzIA4efF/b+Ork
pKBXDbH0n7APGSWBqekp1BoTbI/DLnAv5re4g6Ua1FTnGcjo28wAYrDyHOJzbtPR
TRWTo4n/rpbNqjvwkPg2Up5tCYAVY9BQUZ56H7ZdnN0btuifoMG8rEfNHKQP5bEk
ySbfE2LXrZiBpNSABvVqQA904px4FjLSOc/+GSKLiDheS6QtNNzfUzmnC/Stj7UL
qDYjqahXYwiG+RdKc4HJOmTZaGnd0wngBEFkfYQYNJVXgjDzBTy3mf+Pfs01txr8
MegSl1JGbNK6A2G1tiUUp2HntUVNGbNn7kJrS6wjRdXcZTwpCtoSglu88VFR1afV
PlYKkG7+aGXAiOwaoiHdWxtEHB4Uh4FgwWK3AuXVSw4HjuUlRBHZojdkOjKMxSGV
87Uqzs7URHC9cdZO871JyT52pYgG/CsVJsaMKbqtuwsffsezA3+BI2ZREp0mRrAI
l5X8V20dlb1GsgyCSjCE8oU5mhnEcy2GOa7bic+wvHYMMtIzxiK+ktaDlyzVZFGZ
IvCW6i7kU5WsDxOz/G0CrMgEGgZBvrkTT80WDauiJ2em39XAatlP24RKYPYzYAl3
Y+zP1Thm/wJhUnuorTnJ8E76LyTLuRGUEoVNa6aKNCKyWZpGXmJjnjkPKAU72WCI
iZV/nNTUvQxN6OGLjEp8XJxzqCtq0pGoWtqGj+mielbQcGGy6wxBOPoYNvRNYJCF
lW7WVs3+80VyM5e8BlvRtyzHlgNX4kwd1E+MrRDneIgFyvUbieXI3IppDnaIpvqg
cXJ22BnCFF8gyFDhdCW91CubP8i1wdI6Ggycv4l8Fv2QiBDWsAqBf+QEEyY+gHzD
ttehdcJO3pQvO25YAqJ1eGIbbExXPcFkvUp8NW6jvWHSho0BnR4yhh0B5/UKavv0
3iz8tZFVul2graW0rt80vLaLY7Ox+yts/zJkxt92lGqwwCNbba7KqfI1YQVpGExT
J3up43zlw7C9ftEzU3G75PHtHKtgrtgyaru/Esug3G8+ODC1PmFETpm79n40/zGg
wHsJHnBkzAT+Mxr6yNppAmBkzB+bytis/2pl9pg1XHQe8QbceI46+3+EdDMCmOZd
QNdeaedYU4P6yx0qAk8M6kEs63eVVB4uD9mnPfBXk6m7iP/JIT8OgeIUWNKy9rtN
lR5IUmjT/4Q2prc78qE/vZgt4ykJ4RnpETkSBhDCuMATY1WGBgufs7QjeDCWUQtV
0n06fgG174Bq0gHVedVVj6Qem0uPBMCKj65h9oCOrgppt5pFYYdFHNZsObBg2z0S
9td6b67HltZrTlncV6NoR25BBJMGH7VNQa1m3IpMYn+LMLzaNLdTl/aACYGvVVIh
2l4TLFlQsqtlstgwT8B58uJMGTg0GjiVPHbgF02yFVcUgR00/0J7+r1eqUdSm8LF
63VXUSpuyxEdinWHZ8T2jY9RqLd3DkOS99EyvptkNNtcbyW95RiAsbVKhb//9GMW
IpzB0/SvskxfQ9b/7E4UmbBKrr1qzQRUX6Kkz66nRfs5u7e81OkMMK1slJ4p5LuP
nxbdLikvQ+xk+TOwDfzVcZ1c5RJW/0FYd0ZW3/YtMzduSuDkA3ekLvmCWf2Zs0fo
nYMpoVg2CJVKDMfllD89U4om2R5a5jHm0D7kf1KxVlH00gRWbD1t6LSwvUvaGZoF
1KL6R6RSqglLHSfUYcNhi6uXV54yecF8f1WbA9yBQScEmV6R5pdlUfuCCtd3w8dN
SXMl37rBtcANyBNgdkOjWekHI79Vbc0GMuRkRBjYZ1yRJHctZlTYmFTBWb+o7zJ+
xOZVgg+ZArWW6rI/oZF0a3hNeuLJHW2p2mjVsC6fMby4IIQqAAjGfvvL/UeJy9VG
s0KaCVx3Ph2JJN9kqfR+9Oz+vTLB9k+ULO3WEP4+kZuzk3LBqMdH6hEmlOMuXurU
1kIIu/IzL0Jc6QJu1u6OHj4GlZdK0bhllEo4NiLQeWDC8kLT4lcAK8e6EHfupOu4
YbPJLwaTwTWrzpqo13DXgm/HmvSvGZdPRSi8LXNzUgzOZ+OoCuYlZoakXCtGicM5
6wPFshflt5ZP2NrFBUdYpufwfMAT9XCa7L7KnyJK6442+/ET3lOk/+PRkOOc4w8H
70hwV2uYbByIN/WtxnZIMvKEZ9kyyN0qDJ9T2Haa4ynQ8HQGtQbWEEKJ6CoERrjk
M363ze0nBgOaDvlWCaSQp1SnnoPJKHzHh66g9QFPqjGEOQRwF8nzJMf5GhqNlJ2t
Lj7TLb0fJwdbBw7qfZGA4cK5d61dEbG18/eFz18CcpohX5W/wlsg5pUt90hLF8V/
tmr8Y0wA/VrSi/Mktpl+duRBh6OOs66R+5awVNSqhZ6a8oRZiGMw/k3lLyVOgOxk
d6n7eTi7RJvANGpuGh3/A656zF4D+TpBuxQ78y3CfurbkIWU+5wAc734ffJewgzs
mUuuWA0dIngYQyPNJCUFw1TbZ598QwbmMGMH+f88GtYTSlKnx69JrbAGhYVej66r
Xew3HoYKSIFFpqUcHZZ3HKdO8MJb0OfBy/Ik5GRi9CaQKkqnefHsJMgFTvZlA4BL
4M65Rk9wZwUcqOu7WYIc19oDTth5Cm90yA4t5GiQdBGtRX8o3D+9XhIk5ckN5y5B
QWgQWVvsmJ/YtCQpK5u67fTsUpT9PRfx24q17IbqP7K2Gpf5MaBETqUCSw/LDCc9
qnQAwJ5YeCZA7vXeO8vT9ReJJI2Ysdu8WERxZPMGQ85GixEOGzRgd4K5Kkjzefqv
ktpPhVsGfSm/xdfk0FCh9yUM5SLz081j+hNkzOWVe4z4iJxlIO6rYZX1RtW6xjvS
KCVhdB9KhrJ2kQVc0U3JZ/wR/xZhj2E5HnICoKVDF6ZgYwKZCuH8YCN43szlvpsc
lqlF8KPMUbFxkOr9w+9FV1ccB6M3R7RIW9HuM/EKoRXHoApKAdd6tbsf+bzQqTtw
OaKRsCfm2+r9AbLUE7r03UWBAJsQBA74Sj7VQJaYURgUePxx+nouJUZlRVJDe7nd
OqqTrMM+lpmdjYWdkKoR2t7L4e0kG5ZP+G2WecdppGKrHJtZtVlxESggpL7xU8gg
rcfhLpjqlBR18IgC+RUXggv9Tu1HeKVOsoQDxmC04an6r7OeS0Iuzm/CnF1F+a1t
hNrj8ZR+zJBMgF/U6NMf/rXdRL4ZG325qmJlDWdXUDe4HJRPR5ywBTtDFis8Lh62
mHzGN73fN3O0o/KiXhgzwcsjq2cJZQKXKi4N8F/sKhCDvqjOEUEx8+HLAKdnft1W
QC2rL3Ub6Fs4mw1J3k4RYlaXbKPcnkDQWAlQxZU4g/lkw5QHsNMgYfYryOw2AH+t
tb0NLEmQmYy66zWeL7H7KLrv/dFxkxp9IZgChWtHZrh9SP3KAuZn4jjKJaP7C2nP
62lSPluyaGXOQl9Tb6aYcVxOm8FH5Btl18PDLDcme6bw7jz8lhpSH9SZWCVbcTGq
olnLwz0ntNqRjjvr8j4g9piqnLk1QcTEN14lIG50mPtlUSuTQaoeSVJSdETS7p2f
ldYmouCh3DyPQr7qAVSEdr+7aJNUQfzpwYo/VgybxivHcsCXpIb0pbsZhKjCwOKP
rqmBD/v/UPbILh/qHH9SEhEEcgemLM5DYjVSVq8PQkFuk7lWlNilxq3yJ6FXVhOd
z84aI1LTzRcpI8bHbAtJBnRkyjq6iscQG7m6ymvpsUoCPOp6RZa8fPjlIyHEmN8b
84/yrGXODTmuflhGSajkZRAQDtwwBW1f7cqq5Di7glezdUWdIu214lPVmRbhfdIX
wCsENEtaxGnxHI2eFnhAOzr/Pm115kKZXCFNpmVhtrms2xuiqyTmJPamZ+4FeK8v
ZpfaRTdgBMNnUxQCuE+CNErW5t8wyk6XM9UJorqUn+ukHOouXSOgELgtDSLnfrrp
0fo038QHuq6c/9sq0112lROY36XnwMVdSf1XDZKufKbHqEK6O5WSXD/mI2/iEreG
SoYKyfSAgSSaCz4kQuTZqrPHMHmlm66h0BcUdJkslnwSmTzzEdARF0t6S7iAombk
f0SXjZK9zOcLUWaM9qkGEhNs4D9wWscDUkiG8sDlqe4cP5TuPtpWx46Be/Wv312n
obckeqN1wLHGc3117LEXzdLkyZxvzlJ6Iy8Ji6jchP+Vjs4eZZgJcCks8Pd5Pugl
F94e5WciG7RsTmkqEiWgTLNsddRVhNAfwMaL/ud6+sEzvOzvtqDO+97y3KmHxzRt
pCw2w+CRbXAfILdL319qDkd3DPvRlgIGQuA1RgDYGzPZfXgrElftN3eFVExQL5v4
7+T4D3uqtvhtjHMtQtPSFnqS/jFY4njVgTGDLHOAT5l8pdwGEowsljWofUEiKcxI
336kppdbejRuagDeaYms0yypUmt0MdVqYpFSPGMe7WfPxdFwwynpsCIviM+JCsRA
nFWEGKEPcSX1sLTmOTtJDUW+iNM+7CthV/VkRaYJYYO/ZdxJ/uGS9eb3l2BWeFsC
yWWTACTX/KMEJMyZ+Y0k5LdqbQzKIQqQ3YvxV4EblEnUIuOWnfXstKCUNktSj5Ih
lrE8MdwTPY+5rtJlNT8OTAr808WNQaH9E06G2+mTSFHYyYW0Wilx1v8v/jksqJQX
T2nF7ym/2Slixh6tpgPRiXGaMmXEnsTzMhffG4+4GQCwV1Ihayit0F6qujOXWb+F
1PBQmYeorEObEBIQOV5058y+fzGlGs4qzwC8lsjs14+aAqlmDLTf0fzFZw5r6H2u
wF0cUfQ1oZbZrUdmCEp6/rakpgGsMhjbFcsDswwfuuR/sMKQm76WBpHixJmDvVoI
RuVcxX9hjScpjHKwJqrUaL/aiR1bFGAqlDlNYuEnGZz8KcZhQbO+CZXddAH3HbpP
d9wfQrZa5l7Wkbne9PDsaBj1NyBZ4AfR0DHQx41q+U8jFHy1ctmgh2HHI6ZBfP4J
TeZfey6KxuYhSPKr9HV3d47uJiXeHvJb2/oZw76+C9kbNDt6e6G3ljcUmObLlOsi
JKvRECYLDt5lcsWzEINIha8VH9GK/iA7m83akJJ739onfCCnBz6JKaufj7/8AfUM
dmSGyPfhWnF83ixtAI8ut5GPfXNklNIACKyWb6IbItMsUKy3FhsZV+5QENbcxkK4
YQ+rOFA4mIYm8S389hHDlh3l7zKLv7A5G6pnvU0SlauctAxZO8W0FwAiX0gHe8Ik
Xib7ns53SahUj+33vicfpwV5ZuvJYVJpfPYUMSkVGQhII8td3l3XgZM1Glw3rD7Y
Ve9xLBaFBaYfKfLaNvE+VvcoMTFPmySo+jQOQXX0OQx8fmTkYmcymqht32i1QVbs
hwESo13GpFX7UcS++upQdKlXSbFVooWKZaq5JkSFIZT8/DFTv4Rt3vJk2Nx6qGs/
zFiKwoJ0wrakjiJDbPKmzdMNcwWmddOLFZlP3DF1Kdk/9Q+nR346qaz6C1PlqCae
5mOx+1u+cIL42yc0wHV1W8BATcM3AQ5GoeA/8/l6CFUs2qKsV/mGpbAcf4tw1XnC
vS+OPAV4MmZxCYEAsAym0bTyls8xXkVk15UN6IBdJyEhQYT6ztPXlB71WNZuIru9
m4uEr9YWgEGzyblhb9EoAvufV8UKGX5CzSlWLCSlqWRMj2CSJKpfU0QXK1UMETjy
04fvXTktx6VjO9BC7HOLNQ8IZ48Gd7cvU1xDO/Zm21vWd5laWhkqwLbJO9bhPPwA
C7l6egTajzXv6rbdcG+7jR3SF1vpoOnuo5YpCzpQjBben7rIg6ZYRnEmDPE4RVDM
LoxEumK4/YM0Rpl5vyPeXRUfG5QSRBP45tzEq2u9IGHD7nyhTz3bn+9aVK9cNROF
YRyZe0CMNKCOF8aws5F1WaprCE0R7AXpxcGl2q/cdQoDX72kOIbGWV//m+9sYwkB
1OftT7ACQuurIjf5s+zS8Vus/lUoGgMV6GWVMHZ65/A2gA2YiPOSVKSlzT4phTy3
uBdJnteIAo13EcaXAU4g6BhPkPEXelh+vwAul7UUz5G1M0rkLep1VEnNVXE0F8FW
DMBhu+smEXyQb0hR4UUYzM1BpEXDd9Efkkbf6YKKrCBu1rcTZsVH7Z4J6hQxcc8q
grQGIJtD4SKFO7fxpfi0tWM1OiwL2uQLSoJiNNHzboGVMQhSQlke6FGCAKdBkYzp
0k0TDStJiHGXrf51xZCJJk6dATdXjwl8HsA1JVIC6wo2SJ9zmKjZ4jgkMnpkHX8R
L36kw3vEuoDd2boMwY1LjY2Eze/PUngJoOxgg7xLfKZIl/8oPukjR6186K8tA1n5
PczzwMER/hNyppClB46ttC8E6X33rH1t3pP2zdJv1t/T5gyuIL0h2jgiNFMYoFzk
Ty8ARDWDHyaq4jiGH0UEQR8uSNOxyxuXjIyykj435yYuJt4lWmYlM+Xx87YAeSqf
DD4pUkgTEY7FgbOsRvacm9Y3zL7yZJhvtZMNSvsmQ0xjZyRsmFNWzIDXjJnteTj7
w9LketEh7olu2kkuvEeGUF72xvEADhErDyCz6eHL2FRCHfr7fgQgdtfWEZKRHKdp
D4mo4HPxbqJNz1sAVRz9W/UQ0JMPQjUPqX4UxxfsVn/HbgLKW3FsV350mA6tuHh4
kCFw83yaLfa27LYaUKypUi8qvBatn67BTmSTmIzqDDgrj8rmL2gJFDZBlZL3bw9N
H618eb59V5y7jCaFbklH1uHkPjiqbebJKA7BVz0pipvgBwtR0HbuF0khOCBBPEDL
wfvk/FUuU6l0KaNKg2NTqB155qMpVA33FsPTR6VoAgqXA5u5oJktxheLJI2MASFt
cNnTLtyPdaA30P2VGgNKJ+eJCx++RcuMivchEyS093TxDk/Fi8h4gVQyEOHXjs0V
Y+cUX9PuzOnAgsnR0SrI9Fntg35bU0vnw8z+JB7dXUWOHXmehj5NVcdU/XD8A62g
cEuCgPk1BNAWObWQDcKGwZYu4FLhUCcQ7EzH/l44WIXgcvTJm7gnzhyd8pNTBpxW
zNGbWMrI0gz65KS++6yVlkni4WntRj+mH+pyPY7kUmseOcOAGIGUzg5KJtGRYgw3
ymf3umN7JHmfHY4z+dLtkvQ54wJHDCPl4+KpuM/34uYnD03O1WmY2dBkF/1hDfcZ
IPioRFYHeNF7yHQZEx7CRjyCE117rxoqBCGBlO8Dv0M4yZYghq1usSr+vQd7EaT/
z/TqTP4cfK6z0a9PO51qlZDOnFKuSrWV+yOBRkk6j7qBYkaoMNYy1evSkzlEoJhe
y6tTfauyhGAI+iER265JC0W0AOx6phl2ESuFhM2q7UN0sa6w/ohwCmr6inczLeew
XUqL0syd951jFruHZV+GeEeDhuokdf/0H9ClgYnGkwJ3rh365y/aexS65EZMdbIQ
A0I4WZMhR0O3fy0PPnMSBVu/AaaqGixCQd3x1BFDbngx90ieMUSvwOtrtgH5AQ+/
FrSe2PERL+0D3EVBSgrGkV7W+opEcAgL44Dp4hHcBldZ12L2gA1qPExTAThoBNBc
JKfbHfre1NsAiqsFicKennUZR0NESyJ7YqIDdpGP77iJkmB3akg5PsTiViPauasR
HfpIVLeDWdUDQoe5ZX/zJNkvDO+6jLMrnKDRvaNX9KSlL9G6j+zbhjtWYJBsyrYi
70YMeUOM6xAaVs9TW+bz5rEfC9GnGy0T1pxv1Sn5F5ZFdVTvkICbMps/fCGKzRxf
Q99Kl9JkcsxxAK3R9RpPAFM1wOAyX+2bVmZDge1cKIyjSerj4HVgu3Lu2srYErxB
vYZ0YEGGT7tXO/4AFezDvHFfRL9XdTKVWNz1tjo9iHpsWdXw7qLNJclERjL+cD+V
fSGNQLZJS+olJYY5nO0qpRe+DgO0PvP7ip4y0KnEfC8qtFiYL1WeMjhHzuGRFJhC
eVqI4y/p31tT5P025ERqS7wjq2I5Nfm71RKAfd8JqxObIVr3Ee9ZO9zF4DnxR7w6
WTKFFIwqO0kXzBAYLXsC45XDM9NvO3wKYGFr0iukH9FsqHf73FAPdo7SzICpw2Ef
czzP05kr82KclIIurNr+aot843N/jjcxikMARfG4vmse3PnbdPt3xx2lozJcuS//
yGb/8UKaZfoMG6Q8yuPcOERgRQAyx/NuHPE3uZKTdms71NORKuWjj7xT5e+R8YQh
YtweZhhNpGMlGcLHk5QE9M6FpHZknDY9RvFefbtDZ+VFTjzi7N3YSc7S6Lwj+1Ws
x4RpQ3z/+7b0ZS1HT07E/Te6nAK5iLbge1rtWMR2aVGtS+Q2lTCGOBRr12qls+4S
X0kPGPGyrphUKmY85a+pqAIAxlW1vq/XRWagiY2S0J5S0rmS54QG9FwyAtQA8Ayp
fTiKFqdaUKxKXK3FQyDp+/rF679jLnlcrbOVPaYW0Ji8fP31meeX5hoQX0EtVUSa
QicjjgAgXc5TbKKR0C3Ulmw8MvadR+KVlTMx++67T0av1kfhelZ9JBLVS/Zy2FON
VqsAxo8Ghcegi2kVBfXL3yFn37TCFIEl9CzD7gfHaafO1WzXt2NNtiYf6t8hQSPY
NvgmHrkrE38TunT3YXjdzfKKKW+xSCtKNU4fO5lZcdWxumFoXhx3CIruteUQfbri
z7WcbK0HUXPkzHeUcb1kPo8jyEXs220J1WshZ2hWn5G2nXa0phmLL95oe8NgGRyZ
e2ChQVx8Dcy0poeAPCFsuy9WOExtNb09Dfw7HPp3WabtRzW6Qh5v5Bhig7luoa/9
XWWGNp8V7gM2lV4GMoF4tHf6luP2qF7GJCasEOUKSq6xB5A82jiGNonif3/iWfNv
HRSy819/wNcbS3kGuISfiwVtxlOzIaECkxTXF9+hh2rO0eAMnW+3Aiun1vz5x8aU
qRds1YprGKt+TsGqXYQ5GDAFxJZiHXNlp6VtOT4/sFclkrFtW/bJPlKcZYgYgpQR
p+TxS4Pct+LxYlLR1lIq+fI1v9SXMQhZGmJDYDj2ApvSfV+uM/s5FvtZ6xblLRWi
fDEiJ6+vAhPDnw9v+BgEXJ1FSuT4EO6unSY9Xu723l22mhiwA3d9vSTTvS6RMpyg
qXlzKVIPDgb9C4aT7sBUjFOPvJM/AkOQMpYZZvDZLeniNVHregBgOYei5AJ2zaou
cLWsmR0+FdwKgHdvTMBxuXuXPusSWLdAh+ISr1lHXGPkgYOYWaTZEYb/rxDTaABh
5ZXYWe3qmdWIyZQmUghxApZ6OzwzcQJr+bxewL9BBjkezl7RvRW8mkyBDycIYlQJ
KodwM4UolBact8Fr8LEncnJiG91wFMl4xLGSiHla4unMo9yMU+fHgBNGkT2SYrC2
EP/9kFAU9Q4iyzctJdZXw8zN0/+57gGlWg++xDM5Hcj7XE7B0kPrT6t5mSckGtlc
vx/RBBRL4Kl7filvwUom/WDuOdWHbRjQhKqz0QbDtzvkXJwBLSAeK8PkmM50T61N
lhQIZSfqWVZ+nPRPamT7bS8czdgbFhQNpMJGcHxxpMinFWg8qU8kvL5b3axp5plv
f7LBEQXHXNFrMvCEd7lCPCWzR6n1ysgMTKtv3aGDb0MbAtnKGQCzJszIDGXuLHQ7
LF8a03FSLNFhlgaE4fF8zGoCgU9bZVsl5Xw5LS3AiYL00mkqIl3JXAwnS9iYn7u0
uq8qpRwmdL0YkNtfIQrkKggkAEr7KvFuxsGYYuMmZXpy8g55cyMO8oETp4ie7Zw2
OKli/GYAoyEXtbWdvP3ja5/ghaRV+q2ZdkBsAB+HAvD1c2NhiylTJnC/Q9i6ye2o
mWC8kf7gBlvAbEsICS+Ib40uBQAIFtDJG/uNrfTxTD8Yo9rqmRyH7kqUAmO426g5
IHx2OiP2ygijgWuDW8XlcOsH9hfcKeCq9qFRsy/h9vupDVJVYBixCuuudwdTLJnS
TLrdSexWrfuJn2trJTgFSfs2lGH3YhCrYPG18fbZztBXNwIub86TWUu1Gj+XYaw3
hq4LXgjJf8WatPM0fSn7hFBtlWPEl/YO7oANBJJtdknEHnSQS6AXirvJLf+OLVUq
EABDNQ/rPdp3+j2V0Z9ztFHiVfw1Y5qZG/WmavO/N+n+m6yjP9sO/DNU/gOVIN2N
WiY4QyqKdSXyVS2Ac9yjw7rUUOxXyU7mLVQbkZ8I03ekmdPftgq39Y9t5m/21Z9x
5TLRDPbQQhXbOucG2vTjZwmNDBvf1g86Hx1o6Q05PfaDN0wDuz4IZyqtFqPnTFK1
VEdPKLJWjRiJK4XKfh5kyEW/0OuRMh8UAKB5zWE3UQs8ruApTBrLjP/PaCh9hpN5
me6S1MaQVssIVM4l3XqM1rgpxe9LBNp9mOGf/CN/3MeuOkrGqVBtJko9Cqu2Rmo8
qov06NZQMNL2vbbE8jcCLNKrr39sQbiSYqzyIDP0iF87W353UmZipiaH22FWqS46
xxNx11uISx7/tXTeWSvzmSKv+r5jmD3Yg7off2dLxDOfaL4Y2iQ/S3uq2pbwqrCJ
XfENigBFJ1e36a+3Nislq3b+bjxlLVkkGo711HkpV3D3fj+icx5F9DwpApr6qfEh
otNTkA6EWOcv6ud5HC14tQy2mzydIAGnWDF6pohh8Gyodd8dsG7fiG7KTIcXt1gT
LTH17fpDhDDGEusPJfPKB5bNCdeHB7JsP1LkGUaOFxJMuZRN6Ccd7bmM0QbM99Bw
gyMxMaphXuMOZKU3oHe8MLmCjQAJXjYDv3wE+qfUxGXZVcmBqnAJ9oUisK885XYj
00MYiLPx3mU9MQeKhnOzWgsmPSvdnqJXwN3JPBwMnm7LYnZDoVnJ+ZlmThk1JbUl
9ImnuJpwgdDFP3a1YHzBzm8DuDfaiIeppP1Z/GXMcekQFn+8aOa2en+l/l6i/6Wb
3+ECCjSo8+ihQCrGeKGHUymWmtjXYcZMTYeQnTQK1+JFoeHBDk+j/vR7CDWFmevY
Jj8zRfCAmdauaGl4lNP0Iq7UydpT8cZWqneQea23V+DDcXT/G4DEZTp2dlDE9+XA
IsRXbnBbqHYK1sWcrauczn7i74vHGnjJ8FaRbnj4VmHu6in24dzuThHNKlNQ0+f3
Ws+8oJAdiGW9yb5BALi6dFjH7gJLMZ+iIUe3pTklXlHy/ScM32pRRvwc5NoLXaXy
/UhAPWa90eLvS71UUX3PaLlVDpPL8t9XTkOJorQJaxg3d84VkCzq+azl+tDiN5UN
vkoPUKVMxe/fpItX4CTq8NSojV5Qu0DDBNRoRpx7bDmXmRVTJchbZYMjCU2QUE/N
wP6ni2n6jcHEtVuM4FnzSn7JLUwYC8ZmllztcTYSgoHK4cS4jii8dwRQQrmqCais
X7cxLUE0BcR/MnDVDul627YRRMhUnmzqRWnJw8q9Up9neAVmLc9EF6AWG+oZmSQd
uTIUPuN3OksgbKGg33X9wlcjYJ19dFGL9MyDK3TuMunluyXSjb2hujbYB8VV5eD1
82XTICRSrgJhSMPdMm7J+jqThYUo15BMzmLm1IK4oiXKDgiHY1tMTdjtvKZROG+9
32PfmahmqzL+C4KjTntJtAR0Ndvf1tSZm8212UWbL0vfloh4BR2y6UOC6e6TxV0R
/uuD/z+VSPQI0oFUniHhl3fMIus5xotZKmXzIhfPm0JaEUT+X3O5loxfmPHMhoSO
T2ohpMPB62nXtBq34ud00pUQ+P7gpje9foF6uCaSYTkSB4UE8WaVY26GrCNUvR8S
4pl2EhR7wUl5Doqd3ySJOt3rWNJwicHESn9IBOvcjBH7yrFAk0DsKEqK3IQEjo5I
X+67wd0Q2jzeh40KsxpRTDqpABQtQEYFnIBhqBYPMcE//af3sUwgRJW9oILr3wRa
di20WGL8Ju2xkPxqKBpNcygXFnSertOfNwSyF5AUQZHyawnjwgemxfdFDrDx3hzQ
4EQc14ldU6w+KZjY0fZgjWUv1x8Tet1Tlntz9ehuoqRskzxPARZ/Nh0XxrBnYdyh
BBZGcel6V5fmR1nDR2vXDODPfq0sPQYCApdXPtf/RrMXZBagtMMOJBO7bYn8WuFB
EWtKkXVw2Jt55b34KwhTXWfSMAQxBOJpbA/Cou7Ica289vpRH5jmeZwYpTdTLuqU
FKVrlN6umLM9t0RYJw88yc/VIx/X1zetHqMYZWXfU0gOgYA4LBVuiOukzIXp7OtO
BGof/gispIXKv0PGT8wTftN9caKueOF+yE/Vl2MOXGWM1lOYORexiC/LbUsNmZg+
5aZSGgz+4JHimNFFT+e7P7vVCo8wTZVBWQG5WdF+WI6+Du+Lij57S1GE15hktcIn
/ohdX7qIGRWaDU2J+VW2gG2Ez12XusmcegFRnReWi2wReoNNTOUfaNnnOXnExmKi
7G48dqfpSnL87GlIeQV4Wp2EfaS47ZMZcpVVzOJHaBw4JOyEdMjabQvO/ii/yARl
5QAk+VZGieQqk+EBaC6RogeVxdnz0E2BzNa3oZmI7S4fnFbDj8IzVuZ1UoASTT1q
hucoT6L3kLBHGH2DBPXfaXslHHkge29DYH80YQSkmdjj4QbfdT1NX8wkmDXwr/NY
ambkpLN6G/oxNOe5s40Nlq/QCbPcYwBwSni8ifJX0HvuyejCC5Pm+pU/UbNnpmsU
+6c3ZyuPOhqjLotjMj3MSrt9PzKUqzc8+7h9JIel9p0iCoDT4jZrVmKwzT8UFH/u
k6XLfyw3PCzsxnguU2fEI1HR48sjAl9/3JhSNciZ2lVAxjSCbWRx93DL5EChddFC
YjRsHii2Xve9SH4BqEK6e5sjiu8/LOnh4RLKPndSanao1dNkVfE7kuu3jkMlWRpG
DlnzMmdKR5awAmwvwenK066ZeQymfupbZGZ4EpK1VZuzwVghok1+g1IN2W76Zrpp
IF9tkpf63OdkQNDn2P+LHdYO1iU5ZzUXyYIpkuj/bqx463XLOSi8MmTI/1yHXkUp
LolZEbCg22fsgM9TZ26BjRZ2OK+zQJLgRuImXKVUqurRhwPTwKRe2/Gp707XQqVo
JG2sUSZ4pfhUqUxxhdlKA/pMOrjnSxOX/GWHbM+Orlwqye79mmvmzb0hTWGJ302S
CqJS/WpQ35ucl7ey7apQwbWYWrSbRMIXXK7+H58YseLb7I/ERzgNW8FMkC1LkxN9
EZd6/V6QNof4fWuA3F8P4d2SlvRaBjVh7+Rc6dABE30ShN1YsH8dfYUzhD0LXpDe
P9sPO0Ry/b4+2UZyk2bqVmcGYCiG9hNMWVgyZD3OYlBS8cXkyHbORkZBEiSdYHj4
gNBDL1m+SXbf8v3OF98EcBBDEeZhOqAOkTPvSbd4ZY8EKenEnGI4MBWwQQf3832m
TzacL8tjTxuBGaL68wbP0bXRUWJH30ctuEd1CseVV4DDWd+BPU+q1JreLig8Ikkg
4fv5dvQRvWDzxWNoinkZPJ1BOaVtCAA6hJJBaNiSSoTSO5N+MZQuxtgJ8+ZmO0vU
zUOCGVsNrEZ5H3+1MBgCIlD4/+3LwXEiNK4RZH8ivLbzMPnJFI+6+jnQ5fsvEMCl
V8KCTENhaxkPt0XCVjllMUzphj8XV52TZScE2sj5fO/yXMvhWr252H4j/Zw+i6/N
OwBEjjtvBmV//Om6Ruz5iMIjXJ2M1Fde6H4pd+3mjYOWE+vcNIR7ob0iXcjGmTXZ
IGICIfAeFnLWL6TkTwPCETBHaMjs+gV8gGluIYOTeAJsCDtr/eeVVykPUcH2K+Iy
mQcctrLCRIhGdCVafwPVQBmkFodgXxG8MaJUsHH3hEDnVdVWlANob2n+eHPxmHIa
RuR5DPZwRr8Q2mWS9aoEiUnAL+5j2faElq3KvINZdF8FMkmgxKvQ1MEt8eifOjMu
oMVKgz94mtiLMkJXraT2+pABaeCtQ+2Y9tvLv61M/Iz2uIg1OHnwOKUDv+YSW3/N
blbaBxLHhoqDoHT9fEzRoQpvsJZLh4r8gZApr5WrHrQ0BS7l2gQ1SoXiwneJVsNg
T3zZ1FaNU4w5wOPII0cfRGfJ32CiwqV92KoGH0KVO1B+NrpIkn5C8hdHNWgKifM0
/OipZ7O4SrypGjjibo3RqJ9t6QCQIsy/gGFeDSZ/ImLErOQ41CrUeyRFHkzNP6Jp
YHcN5Els5ccn5dsKWNQ5F9a6/BRoSW+C1Qg4d7QQ/T2yl6VIN01vUAjoxLBFeV3s
aP1MDzKB0b3C6EE0dLtq7SjMlNKqdSedMdpUrtWKWP619lJxBjp2p8euczmv2H1w
o1DIdZg5aOFgW3QC2BfPqxo71wrlGBu/tOPkZoJzFhsZLYUhiUz8xwFZzY5f5czo
MJMqK8Ocwoqw5298h2ZYtBSRyEthFsC97Ule2hSlBz6MeddLtR3Noep7Gtc0WFm+
P1M4oC478CeePA/qP+gwGVJhw2tQw0X//RG2eAtjhS/BQKAge2XeqBb62Q4NK02W
KXAYSih1vAAdCLPkTpL9NWphNwbGJthCX6cfWTkBQwWKoziy1C1UiYQ43CHuUa3B
98n0+1ffhn5ABebd3jELI7VZOJFZD1I+i6tMnmScLNz8OInyWuzkFL+Y+6hHB25f
uuPgO2l4khvnb+6OtCmWtyONi9U8CCnM6M4cK0D3FmPUUDmSHTlWcY25Zdf8KsAa
XDxyr1DRLRSD5Duy44iqhYzpwrT5I3OKITnI+sRk4zppYnmva5hl7KhN6UGO4/px
+6MImBiUrxydL6dtNBeFsWmIYTKoe1iDpBh+qeUEQx0RgUJ6imHxYOBE8tdFBfKM
HR6C0UMiUFJxuIP3L3NZWiK0JeXU73PTcYozdeFmWPzy8YCrGvE5mADJrzkoapV1
X5tfd/yZ0NO03XX2/KR4Nolqxo4u79iYundyA4AgTP9HOrwrC4E2j8rP2FGVbBMr
5QzsOV8Ro4TuiwRXRnZyapfbHf1hr7qcJYOxUOlqoB2tU7QNMHo5Ugs8piFecLCh
rdT7DJO08W7l9W9DhZnVbx7anK/HjLNiRFwuEcinmmxoBHVElxk2oLsvYdlAoqCW
zfH3+yGZddhEIE34w38j/iaM/j05VRDHySefFp+iaVpyJ1Vuqzhbz94pTDSno43v
3dCmup0sJqi9ilx/5GS0f0RKG12frvuz393j+FMgf6ut/tWHltNgdhCVvF3NyIK5
kQjblLzn+ONNIJwDNt+LO1dtHUqMKd8TzZETCJ6YyNEF01nHDhBs3kR/BfxDg5Nz
wzj4Yfldop2P1w0CIUAxb0pwBDeXhzMZ82HITVC5SodGA9Emm67q9xZqHRjgZVKf
tQBFfUJutkQGstYwc9zYVXLyGffOZ/Kjqqqqoz4VMyKaMbI+6pfh7pqkhtcoGlYr
5h2LLHBnTVSvbrsHYGtSaRQOmZIbgY8opcUB16T4Uk7iF7EAvdyUUfwi3SyKTKjG
2nMI6C3hQeMsGzuuKQ1uYwNFeqR9/zVMQDJR7tOmNcVQPmqeAyd0x+PIdhewUnVD
TyEbAN/8TfdtvRa2qPZSud7C5BncPd2JtYUx1CdCxcoId1S4AXTXOMhojjZX9xqB
N3DVl50kRf4jm/XFL0MA49huYWSXDvG+cCA1UZWnPeTgZ9n+kmSHXlB6smLjqxwa
cAx05hKm2Ma2hKn02j3YGGAgdTQ+TwcKXk0qyUPigx5gZiwd3gFTdd+k8umJEH/r
ROv6xPCgDhE4I7w24Qmn/0D5wp58ubHBu4hkvtxPOP8mtrlretves4/ZRWkwlzmF
Th5dnfXueE5iCad1e1H0jXbSMRMh2lM29HeQGzrpJ586eOodvaD97zMPPUdrBYbp
+QWVdxdYCPlWYFV3ALLVfMdpFxYjUnaBZWfYv2hFw3NAJ3vxNrHzVz7TjTws+Cgq
8COVpZP7uDjxZdgCXsz2ykfOQFIrKEaxN7yHbUrkZdWeypeFg/16sCh/PKpLO23v
UvAfJjOyPQzdqwA299Py8NPU6q/Qk+xY7/0gmB1oT8DIJemyJwUJWKlVR73gQlDk
13A5drgwJZjWz+kVXoTyVHDK33jfmPQn/EJk0TeDJ1LpMT1e7sx84ol5dMOu4RAS
0aeC02nEKSca6Qen04uQrxLNHFu8wCAZJTviq6gZST3WC46t0PEzcwyj9qiRGoEH
s6Tf5H5tv2CKW8ZKK1zRSfZGCDaR32MT8tjF3uLFA0jRmEOsat5qKMfnwVaozbT9
5yyLhV00OqL3K8GZvlXyJPNtQ0fNPim4hW8V/McJFPhJJMRq4AGKb0jxcguv6aWI
tOgNbRpFMRPMIqQ7FpSfU2/OL4hcIhGzINCh/EoK1dUXPHu8D31YM7tsM5Dliw7w
EW/Ca6N5N6TgTJfWcD26DG8c4B8yg7FC8uqojUFlPYavO19CtxU8puNkrtPMEwR2
n8Ap/NeMXNLgo5JkYrXd/qJrKXm04BzH2u5cmdVZG/ZZP1/KifLCf5HIP6hDOEru
3zw0VNI5f2HsimyOoYHVUrRJnCeZUzZ+uVhz9HI3eJ2ApZjFFJ05Y+cWZbmhtT3R
RFouxVjVnG4lynK9y+PUjmPXnAESOQrDrwTtXE3AVM2FVpbwllqBPJiBLxoOv/Jz
8Lzj7kpwCqbiF9oiZLHvb/7gCsb6gGWP0CmDxU1XRvdaQZi69xMlkQ2blVyiUyB4
Yc2AYYhTH6ocoda5dxFTa2SO3o+ksOCaKWZqJEuIhItKLdhaYfkzSHOSq8DbEOWy
CnFP4rHt6bv7JAeXV2we8JCmiKY3ODBWACHFfKhfHS9a1eIcbV0EeurC5DZWkU+U
xjizPywg0TLfq8iAzILwYfol0guAjVxmXNmA2lD69emqvuivNQgnsCbhulrKYi/s
BrKIxmTCtf7yqf2yLoByOflBmv8Yd/HSo7JXiw1NnEy7sjRoR4VCnbSu9U1LM+Nt
b38Vd3tFTpLBRF9+F/Jf2A/keWyeTWKKfO721+0ZOLBv7Kyp6ULzSd7B0HiIhpws
XAZFLvq5ejcpU8y6iQ3rHjB0NEPElDLoyRie8YJGJwAIT/9TunzYTaNp5/FwPGoJ
t65qjJzHBF0B6KOA4DNc39gI5HyfzSRM/MnPt0L4p41uTd8jbr8I4txWqm99/SBM
beUSR7wmoAeEgVKgkgD3cMaELoRNYwkhZhm1I/qYf8Wb81Cip3D1Qf/bUs48L8iG
hNo1+07CFmWbF3IMxH13SKcCodKi0Dxyz6YV7d1yShrDvhVDPB4GAVeI+q66PcS0
XPKgPvAEEHVfZyrOdx7QCiP3cy578AaeS3g2tzoxIi/7sWo0uU9ypRjlQtfSybml
+NuyMOJHrYq+9dTKXGhZjRdKuaDnj1xfiz/B+1u2WhLPJsGL0qeE4HiVHo5kfQH4
W6+IFobrIfYJ7LLP0NcaU4rhIMlZNY2eLogMIfscQDSmPNCAXd+yLVLie8sIs9fa
wkyDWi3t587DYFjCkTZr6o0iqWwltyCEXiGzd6UBejmjJpHTGm9CkqKcmb+In7jt
1hwvsBwWh5+joz1BFcwC/3rIB04IAJ9RxMkMf7aRPTKSt0FwElPDL6XSvDHxAL2+
oLloFjuD/SxREH60B4MX/ZmWwX6hI5n4r7IO1Qh/L5/KuHbwS0dkAutOFj+94ZTk
SfTxz1lSe6RnxQ+8Eb1IsgkpV3x/P5xp94Du/9JO8Bd4NSn2GMjfDIaIB1Gn5EEc
RLLNmj5EHQ4qsRJNK2/W2mXe8Y+DnFib6xvVcAiL+bS4AWDRQd+33JNSLnNhH2Pw
ENlM+EohS6lgV+DOLiG7m/35kBG236/CUyIs5QV0qGSexXFHpPNZ9t2d1MBnWgot
YbNp+eSW5o80ZpkTcpmzLALHEbT+XlynEZQt4cHzKDFzIfuezs5tVkJ4jYtC/1rh
RA98j2Gqb/Oz2eUW5KMjEl822rk58Y/F7c0tNBOut1qiR9v4cF/v+ir/ERZ3vOBK
9gJxm4TNBiQWi87Lb8xUOuluw7xk3sXQBFvqWBbyGllPjIvFTytjoe8Qq5POqsft
FEbA1ucfYYfjLY6KktF3X/PBztmlOHFNSfegcth4uAem9Q5HJJQzAJWnXtKeVHrA
oZ+el/GwRNJ/QHQ351FJ4cSoZfDSZrQq0mokHEv235BonITe/lt1iD6A4pFldWx2
rHaNWWB65RCDONuf5Jp1ItZ4mry/661Lap9XPf2HikVzWXIFjSnSt8bB7FhMIjQh
XCBJT8BxvhZgMOcggoqgfn0NyctoPlxmDRCP2NK6nf/wBcGCLUiiN4vtV8NQk5Jd
z5H2UaMijYti3iRikavK0Raa6hoHsxCZ898Ntqq7ae+pSdoGsXQOJfmPMVGvyCp4
GmyHy7OF1qZsKVpcwnYjAvyR/Ied4bllue7ZrYyybFfP9ruxOUa4GbckoRKbkCvt
UihP3MgPQD2C9Zxx3reNwE4hM1SbrrD72TMpSFfIzaXWE886AHn/+bLjp6vCygMb
nod7N9gNLO34SABNxWSDP3qUq2jyN/bn4CiUjyS+wKISrhIN4z/CdOl15T5KvaDY
iE725P33HAYHQ9lYCM9ap7Fe8ihcQqmwyREFFkYDpIgr9QgPLpSkk0AwtnRFGItR
UFHKglLx/xEXHHiVSCD0VYzm1ZrYMQZLKBHunIMB7rvzzSf3x3drVtpGjycHiN35
qVOaKb9VsrQGn6m/tOOlXHPg8zFpFDpKE0aoCtsVJUn6fQghpJTGUOmphXLyhs4I
/k8c3gutCk2d7PTa35MdsJCScDlA96FR0ERXtCqq8z7aaFIfBX8xSekXh0HW1WFH
fDNDgEUW1V2WTVR7vj3rQaVaSOxL7PxZZ4isZZXqrYlekUudFy2hDfE2IJ47cVtb
n9eDI7AE9nHOTNv6FmzRxGPoK0NtKnEs0pzqdP+zCSGP8PWbIDzJIOJNNTBMvTEk
dOxH5oBI8Rl4s03r9CS56viD5YzRXkyF3mfO7fRL52qpX/TFL0G9TyK43CwlHFPy
vxJIELxwiwJy7IpxWX/aUKPVDPc7qCV2nMTkDnlir/6joPtv+FiyU2O0BWkhvoQR
uR7MafHCnrLKAkXCm24yG2aJTwzzOJb0zDuMhYjFbPWZHRyuAgiY1EQ3d3o5E8/O
C1kOZwxrdlT4jJxBlGq6q1xKnqLCO9tgBL+QW1p4V8+Aaee8/GO2HD4rOIp6gJRz
ZLF9YLjDcGI22eV9s/w8lZEfjD4oBCZ2CIstroD33Sd3tiOiKgt8mfiVVrvS3VeA
sefu1OoEckPVx7iWvZLSxafhcaJS9x2gvZIVw8gHIomczm0wu05225b7kqsvC9Es
e0Q9SCU+8AUidqiyCFwii4XphuHt5eXBZmK5EUpKq5f/F21tgqqcduCK+FeKtlWu
GFeLtesckR9u0St11/0Vid4UWoiaQcT4IS1Y2nCQDxawexm2HvG8CVOSkP5ccodz
kv2vtR2fJwShP5PItK0grGNHmMzIGL5Hm/CMt0cSwXmWLVb7ANzGKp3e4GJx/8tY
eXpZd4lqyPvODU4SKC2s30E6M9WvLNL6iJfW2V8FSHPl0Kzt4cIzJiXvzOhJFll9
zbzX1/lrSBU7cGqtCPlv8TLBx0Xvee+uEjJoVeuNJH8x2lmDAKNb++8NyLe/rF6m
xL09QqQTSVmzvX3ANFZYG4dm9wh6fS595vwXNo0SYLJkuEOlaEK8iD5hIhA3Xjvy
MokSr+iUpH3LyC34EECqkC0wtWbjH6b0R+GwjUH3BJrOy79dh4oziMudHVRC34QM
hveAF2w197GS4OfWxrOEQqaH8uOaI/cOgaOsxio3d2LapqNXWwjUm0aQF9Rr4gzJ
OYdmxkVA91OtzE4euusMH4uyOuSIYnyMa2IvFdrtj78jS37/l6xRAvbggzPYxiqY
UQ33J2SXlfBLgAF99ZeJdPP1gg8isKySuy04f70/5Tq6ZEm5khwR7W4TNHKJmBeG
UbhsvF6zguVGUfgVNCRGyA3E1M+qYS2mwlUZiGWHg7xTmnoMNm5GJRb6FQAxxTks
VeDOV6gNc8SrqbgdparIiqm1zSj9hlfdLwyg+o2xM7yluvw3b96rjPvArDibsuzP
R5PwPkjb5WyxkYxqCoL9/ttOi5/XVicFaeCmMdLVEqtA0UCvIz+31Jnowahzes5F
AQe6eKqOaNSNOsJGPr2ZKzRiGUYHpbPzCXVHFi4BaM5CsfMbOpGfPDrcBazVUHU+
qiAhwVctTt9PwbjLL8uM/auehvdZxwC8rsOt6F91Kr+rkIpoMUZSBKiC+v0C0ElJ
WFghgDZUi5xeFA6BimW/wocNhc6ncy4fmLi0JiPqQ/GtB+LwsDS2SiPfpIpii4me
6debhy/wvtGGqO3mkmTiBCzlOXr6XOQxIb7FM6iS2QOR/0p2zChIsUzm5ibYpar6
xGyZTxWiy3C88hupljZPqrzcVAfXQznphwsf6+pvryCtBpGzxj63KVHquuJ/3uZ+
vu2PKcPiRXa3DWmtZZtSYIV3v0SbBok0epkvso4YC85wtT3xMT38pF8K+p1Upglq
k/z+FtP6OY01sTyf49Wjv07+mtd6KCMLcCv7FIVquZ4GEQ8LDx83uXv4UBY9U9fF
ZdYynXrmn6nR32GhAHSWkr0K4/x4V12k7+fy3HiSrn2QDuZmf7iCec3CsrUduA11
+F3w3yPuieohKEAcA3WR3z56RpWirWmOYdro6HVtZqPWGi06ylkqcPrYTduVO/KW
8B8NpBGM6mf3W4FG3f51sYqFhnryeUkJnY/OQ4b5q1bNjXTax2dzque8BG1/zlbA
FPcxV2DQgYxxZRgPHtpBg9/2QceQiMK2C08iEYqrhxSqvG4MiFKO4cKVB5gqjm3G
xe8+Tyvv0wqD5re7oDKwbo6uBMIloB5kd0JQT+oDj/LwTop6mso4T8KBaJBRuoMi
HzqtwoKAltKWjzu7riT2lOUR3yeGhvUBXJGlhqVrFrhS6JDCpLp49VOe9K/MzqJ3
0sCwD4tl9rkXFjkcwgqduzxqeGLqL38aZfor+4pHg+BxgqhfwomwA7Hngfw2QjhC
WzPnx4qIm6i1fP9F7+LKiCUNcgpwsl6rQNEaCHqQ+GYpILdbbrEndIm1alEFRg0+
XfTxOLr2rbsK50utkKwEUteDwuAYGzl3kUVidqkvCQgMY6o7P4DuToOInLK/Pz1X
5aMM8KG8eNIee5BAEl/wQdB08BppNCp8D8jTO5KgRXThwd3kSG45LsU+8saiFxnq
mfsRvjfIwed1mFUWvXfkwC+mnqSSVICPX7hGaxKESDk0TjLrkQeZBHVJ+uwQaiPQ
7gaplp6kyzB4jzuiHsYatHwAVnqH2eoMe8CtXYkApTN48HsWK113PMKiMGRfyIu+
lLKUN0H8MSLLQnfoZWt0Ga/HpXzkv1GMp+Bn5fAJ/QPanRt3B03hoffwSTAxZ2AA
P400LVssefbn/5lH0uBnJ2ttsYyA22VhfUnvCBL5ltN8NzlLAd5gXZWzuQztSbDp
e4ktr6xqKmiQRX4TE0IZVJhmCybkOl0RQZbePDm/NllLvg8WJ01r/u8wOwqsRCMI
FZXujaMIy5rEjrtT6yPqd/Xig0oU2absUC7dP+bPRPZfqNTcYp9W8nuTdJNValqH
gHSpxhdhDNpR9wmDwKS+7GZ1eSmwpzDkfy7kxGDZe95cco482NY+1AhY5WWQp3XE
YXr/rTbsDeLBxoTNCQL2vmCbcgb+3WFO65Xx7BRA23wHwN0HhEk0MQLtSQeOcXll
B/qydUWiLihHCqM5AclbNOi6CgRwBrGj689b7MoHa/xvacPdm6SNDgHS4yYZC++O
jU5c9NjP2nj2xphfQVp/hFQrR9UIYjYp+vbcVvftwI0plFnItOR0Rqy4nxO8hvs1
g0eavok3wVs9oRfCjiQnrBGZyreDuDz+rLV2WQM+VQuw6ugt8kzpDXFHblqADerc
n8Cq0XhrDyu53Lmq1nhAwcqngupc5vQHpEA9YEDgh1HVrcLdHIsmZkVnCuyLqeMT
pmi8FONaLJ9ZlfTUr06HAFCs/CrLFjx7eUJmtTxVj0kfnGsoK+Q0u6JeSrDHjiRH
oungl3ZDFvvTVg8MoINWvzfBOwr40TAwX+jlMi8qlqlIxbM7MHa2fGf7c3Kbnari
Ma8vHjXUGkAv44FE3Wd0LYh1AD2qBKD21Fu8ItQ5FffUW6TGe58+d6cTdWGNCMWl
fc1O2ethB4gIRWFszXFr1/6ph5Xt3GUuqCso8k7sj30TrrSP0nfL8Wm4geYOENzc
cdHjkEzSDM+39+CmnmZEOx3dMRQ1c3fq/OGBhipVe1EaReuMXg0tWnXb/NMrm0yc
vURwR2RLY11kUw3p4ptyYGQi24XS1YJlpGnpCWCUYz3p04WGdDznl68cHib5b8qx
7DQO8LnHJn5Ehvps53hjjcsN7kheU5K2RdnrSp7zTd+6SFQ/NWNuKjjQj3DVNV8G
kIa6vPEp2i0aztSq9QgjbGh0wsKkKuLk4sfw9u8SMAMmxA/d5Fxaj1BwkzQXfbzF
xq1phoozkpxypJkXMGRuLntQjhNRFaBjk1Fio5ZF9jQ1OT6iWMMDVYAGv1EVC5VE
FQnw6n7fQZ85TRYRpZgZ+N0iL507vsOWsOQzqtShQxciW+LKFjFTV+A4ubIv6ikB
EH/wF6s4aCPGONKf0qwKC8D4hX/fI4RdziYnpeuYjtKe1nxOnEnPK7GaDOD9dQce
pinZ1n0IVN4T10CwgC7cVHTXQu4z52AcRb7vK63azQ7/Eszhm9v2znX2fCvid0TQ
2Xx7hmtufFfL7guAvQwldoZ/lT8jneDlNlHPsCkHWLmnwFu2iMWOuSBMC8Q68xkj
/sN6cWEV/1TW4NXDLYQAcaIKf1QEITdVF9jQ5wRtQc2W/+IaWz9wGJYzkdv197wb
DSJXv3BjH1fffR6zAlhTc9r0E+u8akCem7rDjfk2SvAFP/HRPrOWdmzs0vmu+sK8
KV+1Jm8DLwh6jOzfxjxrJVV7i8VYn38Y3h49RYaPAZTgdmRsTrwSNE2O3/wm4tJq
ST3gyu0LbygBNoxAq92FHhCvDmb2u6iLJSdMWyNfHxoXKM1W5ukRyh8hSUdethuE
bxNoaJbEUpYDJCNXzMdCpY+RBPS4S5rys+LzXybLo0KuIupkZ61erPI/QtBsJlPW
I5w50PvUoaoERYnfnYS0yqtUhyAKBp/Jj+pGtjToZFPB3S+GXZZIR5A4hNJhIdHt
LEthTkB1di6rjNCm1S0SJ23/DOkJdGKHbSM5qWhdn14hA6TX+7hjQw81XJaKBH3l
KlJXrQxNRiCZygrucBakvylIINEJRz45D0tN5iN+2oAnYKF1oCmMgHRrIxo0NHqD
62jBv70O1t4c+X0YwLbgr4m28E//mJhAQCriYWDN0gFIQqZEua54VJdC9dGVbW6c
k7/3px90DWQP3B3X+lisOX8Nzng9wXPWFiVgg9vL8IXAy88VGBmwmFFjjxnfaqEt
KqCXYw2+P3ar3oysggcbXXFv6EH2W467kHAdfFZB9J1Htb2wJHJMkLPb0CS+d625
/vnYTm1ofoU/psr5gALfPn76VmgDeIRMZCDf399/qqfUngiHCUufXJaEH/8j1bm/
cfoR84j+VeUlksx0ynyVYvvI38QaPdVi97Se7vmfASK7h4BZghzD2EKYBZKWA+rn
qqiz6hzSrhr4T06so2/hyU/PtCwy+iD/+iAJ2R2Czz4wxcHx6+s/Z6WN+MobW9v9
t/r7zCm8l4kuQbthuLO4E1izDcoPLPlzAsF2NR4MhkffjKWB2AXi0BMtMPVo1Qk+
i3qo4ESd1GJ7KOrgjH/c5gjSur7i/N4Vco9POTxAOyf2z/mTT26PW95Kg4KwAB82
MYCkcPn95aA143GnLzk/lf26bc1oA51j33TMNiNwrz8uPMkTuL15qe1QGAf29rYp
QeW9x0YXHSZiTTVWDI6VC9KP0H8Vc8iRCvXvj64XBL4Wtxnwx2zhJaubU4XMcXFc
rAozvf2prpnYb4rx+Lh3wzdiRyVbu8c1k0XgULrbwuQ2vj0Wn+kwGZX57Dm3Ts8H
V6MuTy6wwHaijWQ7hp9L8RghOMr/2Moz7qeLJoc7LT7OcG5m0Avrdy5sqv42sX7M
S4cUZ7IwzCR2lSG8/u2v/2yeHtSzWyjbovah4CacoLJwA2pl/6+dh3m0biM6OUYw
LzGbd23WUpjIp3EsY7QZF3U9UOdwbxVb5XGiW4WECmTZQZNwLWxGL5aBAsTROupF
ekDVvU+LSJvKSUtzo97meFIEk8VXjFfAZjfRYs5HL05aJEDTIL+EwjFQg34Y5PQV
8dMYnKxK2WCdxDhl7r6KmXXTAC1YuYwwPwE+7jtwSRZ8YzIKXUPVNJbabQuoAdif
eXghwywIWaXlvzE2HJA6ka/cohhxzYz3PEgbzS5CnJFd37728U97q+2e75vCWNSp
yILSFZUweKbiebMo8U8hNGhRJADDkrk4uR+VFX4FKpILHV4N6gYKE/fdKm6+5G0f
H7LbPZh34RAvJoKTPTCAScJnxTRYnfw6q5FY1FQMYgYpn4JGCCSbx2S9Z830nDbP
fBw/BsJ4yUHOT/+3VDdMGD+ezeyXTMg7TjSTeMB6boCNkpZuObDqtIvaWXT9p8ET
m7C+szJo3JC2MJw1Jp/RUrzimY3Buwdx0xKE/MXnJMcavp46LUxMvo7z4a1+SaF2
+5WmO0MKXFs8APdAXPvNHVKd/yaIOn8n7ZqScPJ5WOzDrfCggHcx2ZpXef8t5B+h
zP5o4qx/hTHepj6SdnKxTPQn5gIvcsD/QlUpTa41ouClD4sGHQR+gI+fSR2EeviC
l1zJq6fNSV2zj4eqe/f1gv4SAYV9Y8pE/yUrrCSoFoa/E7V7+ieLa55yz+zorhEx
HAj0lI1wVNmkVFdaOhKLumFW1sqrg3Icn2oy6yKyh9SOQPcjF/gfPMIdl0sPTBpi
m0BAheYHSbNlQHeBah18vMWNqb85RgYmFMMA+/eyywXREJVciJxfoOaGfLyC92OX
lPRnganGm6y1gf+w/26V6Io2YdKqPS+UtGhFy8/IqUaeFgJeKOPlSpnQrOItdEsH
rWbFBRZV5ncvtMhpzSsyTryVlvLs0W4SMh3SiykYjyRzonMiArmM5bCTOWcuiXZ9
8mlASAP923+z7Gc6oSgQ4UL4mYCvrwTzef0FbLRAdpP5oLed/t2AjRCm6ZRKDbl/
tWVjWCMI38kq+lPuvujPf/U7z2XrILqapg3GY5QD//dlPtylHf0BJwfsKy0FHzt+
pGNlY2qATT2cBjd+jOWn95r4abq8t7HUuRSWsGH1Rn0/4LibLV/WUvHAxYpRaFrd
GXKWnA590KcjcT3NudU7i/Dp9Y5/NHtlMNEl5IzLk4ovLANILSmKHci+tu01DTQf
Omu+FybkEorVYh0qi8fTUlKBTw+yyDJso3c/JzmIvJEJNKKx4RGjaLuB7D5SUr2I
GNB7xOcF8CFaqBeITiu94LhtNoVQbt1qSqrR7yL+Ts85iVDO2hw1b5+rCGgodWbV
T4Tmc57WydTa9mngNOEfQ4smD3/x/CD+TUJ370y5DoA8bSGWAAmu91E0mtxU6Ycs
FA+KCD12STkIcnJ8Xrq7KQI0HecprIkOjrx8RAguTmAjcvItU4JRW6AlepipmhOu
/4+6fo1jBMjYHWCCmiRW+bc1r9c1odBX4dA8LMAVfF3z9Ut6IKAvQsj4iNkabrj6
W19O3OSKAagoo048q9AlD3uKo3cwd2ARcoPMWfrjNpQlE1gWnQKwf8v9vbRBdA+B
ZFkl70RUBBKTCPXlwvsQ9sZwDYEuugMHdJjMzxIZeo33RyfVvjV+WfcMLetzWQ4e
136+GxgHxWJoLCey78MyqJSct+rGRKKYVcu1b+L1lZ2GwiQt1imGYh4LlRw4Q+16
iCVM0O3SoGp9PY6odyO6m9ELz9CyjWCrZ3QhZBfbvzNzz8g7rKDfC8p1Pr85qItJ
BWQn5z5kFLPKZfLDB8JU97BWcVHaKXN8FxsHrRhJh6BE1qFgUatSDSYuX/VjhuXE
KtTIKkr7SYA//zbjPQ5/Enjk3/L6axSQC278gzFENxVJxGex96ITWJSTTbKiA7ig
URo8L7fLhNDV5SdXdE/k0CpWFZdpGS/48Olwg5+QoTYEukDH9rRR1k1GhhAg8MkC
bp0wufWPYPmk/EpQNK6haYG04agUhnHmPjM1xPyEkV9TWftLVq+lfZn2Q822ZoV/
SJJEp3S/N9AToJ9i+6WDs78FeiN477SJZghYngUDcMtFqyf7P5WlzuP8HrfDMOeJ
6x2QucuYfnc2xA8zq1fwABhn8XL+GWxOcl7GBtJSQ3sYRWyQz++cZNIaTCJRH+C+
EKK1CvNVkUn7Kobrs19lM0R7xwdZlJD//pWdcfPuVttT0tWFWBpfgk8rLLdtIv7v
bOxvoRaEU4Y5AI5iOs1kcRK93yxS6UMxhSPtXNv1iQfcrn0coubEXO9W2QxosfLD
CDX60izrU4sESs32nwW+r7ZQqIW3CAGPAl5XiiqHkjZvRORZgr6ABnPcZOLyUW0E
JOoEU5jQIkKQvRF8nWCpFBA/mjMUfRA6/BJ9pAqxcRoyzNC8CTsHE8TyqZBsqfUY
LF23QTioGpbCHInNes96mk4dzAYKGFaR327a9BDdXjmmhQiG5xsp7M6Wf3JHLLhk
WlhsbImJ7GsoHuaov1OTVvZhluWn3uqVdiQ8tf7+Otlw/bZ489ldkyFvCkf3nNO3
tgX29ah9Kz6GmDnG5Jm5cfwXk0uS253zXR4DuIXPg5lozMtx90x43otBIUJj0m55
RbPrp9YX9RbSLG0UfznB2QJ8JPpSwx1GWPnY1ymItV0zAK+JRtTEis4XEz5HIqtj
kpT+8cgpCCeYNkkyOH+wt0EfTrXLu0Qn1ffgj70P7bD1jJbyHDYrm7/BA0Bi8n88
UrtlyyIm1EditmCP+QqbdqFz3Vqrcm7b25RA4GO9rVoAGF/k7v4dPtzr1TKL+Zbz
n1hb8X4Stt2RqQmlfDABWhBjsLcpU7O1igMkZjXjTtIu30NXJHEOYfqxVBRniAPY
h5leBYYseZJ30n8fC53izyckg7jbCF6kyG2oKPvT2uVW6jQPLV8A1/lsVqzeTrss
xW3XrCFjojmN0T3QsCMTFcY3UQ6TKdnvGDf5ESzRzIIZXtbIs7o21lM/qglT/3Ko
wtO4NtGsNKXYj8EauM/IxSRVS8Rx+gTU807hza0t8PbWGHCjNauo6FzztvFK+gDf
SMECbRFkGQdkxUE+8iUY2xLREQTZB+9WDAcuxd1AlE/8PsKsJe2GPSgDJhCpUQPq
/83LDHm6EO1/9oVzXHdARdgzSai4iFJzn98MIOeO7tSgpzdJaZrxX8iqzNVqap2l
jXix2UIzsWAbPYG+wtp49PpG7dMsKc6UvCuWjeUEM+C8lLok47VWzxnxaAJOWLCx
jxDd5S3aouuCxownRpgV0xGryZCL6+F6OhwAnLgMm+fcPDcS+JZY9lgOlzLsyH+M
lvqDW+O49qFj7AWA5D8cST01qFCEMBJAwvD7zc04g+IUit1/GeWlWvgtZ9u8scwf
bVuj/SkuuW3OXZ2fjDgSLChEKwdw12aGD5HbrF8PNyuwtq+cwHudregy7IrPxfqV
2QMuF+ejUMDMGyuH3XOI3Efv19SqytECaXPAO2bsLg951iRvL3XHuu6ZjVeHBgwl
xhagPPTm4bTZXPh0/32mNv5ibjyfiG+VodCpvufFOIMIeQ9RFni6xwq0hhm36ns8
iymcnIqT6PC+gi02bp5VnxdtHaaQpE490MuKk7MoIXzB1XbX2CYl1AbajGVclRFO
jdO2nKCzekwvCRZJ5htfQFWO+pUSiBTEM3X/8izVwQkHdXieVFeEx40ju9zZXbcp
oQr7Xuy4LQzM7CYcuGowTf/Bpfu2dADBlvN1IcQqG4BVFhy3n0lqSq6aFuKUo40D
fOoJemMNNJas3c+XbaXSWff3RdKywIY8QrfzNlt6VYRxEj17i4phBaYWAD7q6qgC
LU/gVAoAg13V9jcPZf0Ohr6nCmFBSoAGtdVyPdLiP+N4W2v6YjnEWJi95pKqVQsQ
se/4QZmcCP/eCLcYdz3J+i7PZmppTOXwptA+nAoLOld7Qgf6dAX+N4kUp73dES19
w1NIEmhUl195QOz7gdpfiYFCzF6+4LPHjueTsHp77KF51FsPbA+DUO8UvNH/ysht
ZcyCL0/99hanIzKTHSONRfozcDm2PixLu1kARymvvzLQm+GgDCJrdfNdIjhQ6zQK
F2y49VcJrLbIsvBGpbr0dScpQ3AAdt2lWE2yPPrHbPsEz8ZbEu15huI4tkgfLwdg
tInLwxXE+BupHsW4FuEbQ0SAODQmUFDvY5t0nuMmSX1HR3LTNuU3/K44CaEog3/s
W4vpps7lmz5SxZ8tGT8YKHFQ6vL0oElbDLBCI2z1LSEF9MA+8ph8AinxJ/V0vZIo
CPL8V1VvbQiq+tLGl3vQbjoW/qn1/bpfbm3CNUJq4Lbcb4u31qyfWDgUsTC5Tmdt
xF7Zm1ThBxBiYbKtZQ3gc8ToYLdAL9F5VC78Cu1uJPY/zV1Y31LHkptrkQlwpRgq
p7HeJnrEFYDJxHVu4hO4ltiQSvtRSL+99jzxQshfMSM19vqz7IQkXnmyqMFRx7dl
sBQAxHdkZFmP1CCIbzSoEXwY6e4n5Xxwd5ltlM1SaFXG3MwM9k6fX1XEhhSQtHMU
QtZmnmeJPZlgGjT2inbNvx2qzITTjPfrSfmEs2Cl1BLnFqSBht/Ygg2/8DuFKPpd
wZK1RqcPGBij67NHYidJha9PCg5nj+JDtPyaC/jH7MfY+HXEGF+v5fvaLYNZ/Cws
WyCuE0CvPhCwks6GJBJ1FlFPUFVW8N5wT8lrBBsyQAhK0PiimVTyooBdqZUzgxcI
kd25kWRqhJsKt5CRO3xGj2F7AW6Tj0/Hs45kRcDf1b38JVJp50Jkiela4z7okRfo
15y0eNAuH48gk/gO8/pzMpTkMV80uJrQPxcpLG2I2Z2sdv7pgOerIGOSqT9oG7cY
alStg4qSqlxKw2elGRi/h7/67+hoal/DwoIY+ScJhtKO1MWpgABue0LXCYwkKs77
y9F6tocHfefFjTV2qzkv/l2V/YvFmmn1pKfepTwvqVgYNdbqRRVFYfFDsdmKW5Tj
aj4EidW3bc7cMX23zLkfFZUrLs2EOlvHVplShIW2CTLe9gPs4vPOH7+usCrMBU1s
yypjLkrRx0x911H+i938aFjCcUCXqYYrz6bGufY42aSdX93/f8WO6NllkSTNPPe3
zSrk2UDSrbV/RPKgrpFoJReV+7M/TfsGkLYq0Sm5Fa6b+fEsEoDzj/uFmeEcHHdK
T5I43x5yX8A2pID6QYhZIxzxjYfEYN8SKBvz2p0K5kH+kTpEn0JRme26/SrVXh/d
k0QGsWDRinDGm81IOoZCbxnoc8c5k44e64qhZ3VcrO5Q/rsyXe7Gi5NEZMOGlgFC
YTuM2/La7wSV7Mv5bIdD8AWSwp0kuJp+QB0HfbuJuCBFyrlCjkMa9C5PGOBZO9Xd
Z5lvqm0RL5QgUjCjp4o0wH9raD04qN09QcuoKcp/Grv02L0v7VjGxZAWRAyQgf35
2DbEnwd1uxv+96I3ZKWjc+BHbrI2MXLWHgoKOMeowH9KN8PP3ZjHOd88sXKQmfSv
e4sJ4PJIliWyMq4MdPPnrJ2Bmw+lh9B2UWA3jOrDV2wB/955qNfKN2pWj9u5Vf86
JoixS627TPPctZtReoDHq586szxwMvq4tiJColoHnLmmkIlBPWY4zJmroikGnq22
71K1YlrOf/mUCzk0UtQOmIgAUUc9Lctfq/jcXwb9k4bcwOGVCAA4nJUEHk5Bf2kj
8vIviOdG7oyaa45nZ1zZuPy5QPWo9mf/41kDjHYI3flCVsk/JrZwiKt7dB/9ZzIi
pBwt+8docjQICh3+Q1NLe+YQIQG+colVIvQ8ZEHW9VyGVHiTZdz2diyV4OKni/Zf
qsnlq5ew1higOr/cS/ghzheWDDq+4dKuqqDsGfK3WGQxF3MDb+YxI0UmSQihlSG8
B3IK9v7X6xteJKWiuIWHEdNcAjnTpstlooupzc3IA8/lIY3n7lwcOhyNrZ7MPPOz
jsrzO16ewyeFQMLOFWKfLuqpplcQ7GEJfw5hK/QrDpTvlWsdgvkgXGBw93xvCUgc
7tHHebg03lcEYXG0WiqRjyzYjQcMyMn/26OvQZJ0IJgpXDIM0aClqVoE+6w6mJG4
z8Mzfkj5ytRaxF0CQCrbjgD+olM8pFoIH3DKREtt9IU67UXyzjr1jSsC+wcu9Hin
NT3XKk3V2ADVjLPx3E2C66y5dfcLYyW9Bjn342HvLEqzOm/ap/GMBcDxZrdilgct
zDaeIo54XiAxCfTWSdViHQNILDNkwATa9vvLZelX584GxWpErif7Lrqat6jh0xKM
ngMZ5I1/jXTs/sOOs9oMc9d3iUdbfWAPJilrYZV1VqzAwDFhz64GzABZlROxsgjK
4ID4n7/GQn3oPnvgMZDUnAnEPIBYjyKlRXYIVOG/5vq37ltH71vyDhXpug9oKUpp
Yq3sSRnR2WXgh2JYqL03bJI804w17B7R4EEmIFI/vHy3bCIM+qSQ+hMP6fQ0rUF4
bP98TiXpINmpOqr/S1vfO3x6hS+MRlKgKs9ldl4xVTXiYB2WuGK5GpjZjSKMAqrg
/Tm5cqWOKnr2mZ8vfXrXu9Poa+morJ6rjJ+KyHSo9XvLj0t9DVaDwo20XZjR+fyW
2Hf0TxE8Cm6YNUFzT2pi+2V+MbvSoxuEXINPaIIA8H+VrkX1gMwvfj5estIYQHFT
nnNvDt67UOATSgb1n+IhprX7k3s/j1xZHUMTmmZ9VpwsKK0LNWg5MMMSHGsgiqsD
kNVGTGl5deM0lTlC6h92D084x4WBX6Oqwbmv9A7LyxiQcRGcrmyT9TVgIw6KZXfm
V/j9lSOekyV3x6bMD1fWyDuYIVd46Ki4M0xFOA1lY+EdqshpTwj8CE41K14g1NLq
nOr876lIafNAvhKrPu7sqlYbSwTNrnrVGxmyIXe2Hi2IoyqNHI1nBB4bj3o1Fngj
8wUaXuVgOWPAlp0h2TFD7BP08ddznbdVkB1Y+i4C/TwPQKDO4ruqvvV7F/ngXhFt
XXtOWdpf+8V+IYQ4rz4FSVZIVnUdE7DpuzOFZAKDtl+qUZCrs8t7tXnWekuZqIW5
+LB5b+Ftux/Ya/FGuWGK3ciA/kNOvzdyM1cMu+9AIfXJXsJUukCJTesMZ6WG1t9x
x6RHJrW+K8DV4lRbiSEuihB6jBzEdZmRy30elt3BDIo8JSSzoVl2cqImy/hElRFH
1cMn55Wx4t6A13QWLoNzAgfZsOq6PqZTMq8z+Thx5uggKUau9UXoqXYtljy8XwlN
BfsiYOE5IJHslCYRJh9m17gMs8RvNDjM5cLie/pzXG3YuRUbuDbacxI9qVU4Otdi
8O7u3k+i/xak+L8wvUuCxZT/4HPeBYLa09K5GvqM+yc57PViPrQ/ZqEuJyC+cV/5
YBS0qNvsOhK5VGdvx6s1NImELcAtgtTwQ1fy4K6jv7rXNOBeYK2IhtGPB2KISSF4
DI7E7ahOvKyq7DzkoE0D7yZMWgSnu8xZQDevJhH5xKKRvqttlULK8B3feDH9Ok26
0uW1tpIsFrLIg+VcFDkJrZUsxEvY168Poxf8ZmhD3S7vUj90//x2pCKu7Kyg5Okf
jeVio4CjQakMDNw2n6ic0B1LZ7yn3ReQfbWfRCXO90qgmIxtPuK/Tp+kpgu3+GK1
WeMRnEH2G5862FVCX3wyPif6a10guyiNvOvtnfhTyJaWr51RXAYqucrv44ZD8mJz
uUFNPe5KRVk5ynnAr15LBVTgq+0DKvOKcR2d/6tJap+QG7ai9XyJu/0ccNi9QbYp
W0RYgneS9pcQHO9AU5mqRGIezrkIQ3OXPJlyr/mYSnm1+ZTXxk51D5XMAL7ioYT9
8DHGor7aux+9WK/Mp4gGhdoQLTB/1XKTPmty2S0ULDktCX+0t3PBG5iRoPct/xNm
WqgMf6ptPl8ZUJX3MWL9NikMfS+ggAI+r+euVyQuOtGAPofEf/pS5qepzz9jxWeI
sabtuZalAEBeNU7MN3cUIxQ52jplG09HTd2pHfjMsDgNr6wb9l3QHywaA42y0462
Vz7n28a0biP17x68Lu1bJrjKIrAjDCMlDwnNm0wsIuOj3t9oxYipELA+Ezpbgpu1
UJwldRPiWhNcjZPUqcwpgZDk9XSjzx4pEtCpCeIJuFHAZ0l2lDGMYzq1S6EYvRFi
a0O74KUP58DPTG0y4Pjb+nnHk/gHK9BhamtiWHORVwlnDgQ7qQFgwf3CXMKxZvjh
usZr2SNpod+O1YvNObQNoK1iLTfgNmgMTNKMOlSq80/yyMWLDGiaKsQ+igQY9v1J
o2tBS0ueAy5tB62EOnzEdFDMWpsNVTvnSgVCrPieNXItvs700Sn8WHHFM/CqYMdX
Uo1mNvfWwP2ZmgpucehRe7gzB9aN06fx3iI8r228ijGO9lqOHRciTj+f4CRbiZAl
BHRfPKqVYmnOaycV5H+mIqJ/U1I71CTt0Ts4CWMyFtcD8BZfwbOoB8epDv32RRV4
Rxn2qanKGGEgKKhhbvgB19FVGnvYo2y5IGY9a4b2xQ6mHql2Qr7GAN/+PoYohMQf
bW+E55Lr4mSVM3j7MGVEXbz7GicjJB4Og6V1ofqH/PAPWwf2WYLj8Q5BMJoAKGXp
me4ujkwrLi8BLHOA03G5NxjZMHlNxueTALpmLuGq9C6MhJgp2YQMcYe44rG/5DSR
oXXnmgf3V+vpQR3QHZS+5B693fdY9J4u810o+CHAwaowJpI4LYr0FSegjxyLy65i
+ldGHC5+c+4sz1bUX1bBXETNtgexRA1DpX9AeLf5Qtp5CuBFcP8SeYtfY+0zDiL8
VE7cMixiPPXva40hGE79q8ohtLRlOq3PtnD7w4oKbjkibfAMOz12N8YKcvpFUuid
HU+6A4ErS+z+G7oDL5jucs2UBEXP8trb9olHdpL7IIOqiE6tjNWLy/MFI/ITVHNc
lKOZmq/uf/WPNLTYbfHw0BwhnDmFqvmMHuOSGFiE9mBmn5YOCMy5isG0ySbRENBv
esxQ46QUexbCm7HOpF6Lk3OiIO8jpecAQnQFMHAOWeDU6LtZDZUkyWI6Ca5YgAbt
qljXkcIxMRU7vTlsjmM0QyMsD4Lc0yGkdDjpvSI6j2WqkFQWtowM/LZgwmPyWnkK
k0NG5ja27wAJ2zMxnxTN7xrDO1yPDTDX1EsZsXqxXFNiQM8tQv1TszPKV1dno91A
ZUtAPpTF3iTOLBelpRcKSlyRs03vnZi/Srt3OX7y0BcquGig8/hK7WkJXknyH/O+
NYNFJNa/raY43XfOIRAkh9TwkzvUDGqYaPW5PAUlEhrILW94JCr9UM7FYrtMlDlH
j9Y0nEsVOY44qwUWTvoGIeg2ORVy+1clZMXrtPjTOrLZuvJI6nc7dBxKgujrXpx5
DhRYVNEkvmUpgfkWkZXwMWDZSaEg/yMxa5VUGyj/EzG+SS4oa8W0+WvoKaArJdlM
cMrzqmk1aczZtcRbPCd2V2TOvNoSNfim5GJ/y8jf41cwcD+FECS8gtdGxgT+LWg3
BdOVdI1zplbPbMQiXsYcHyLqo8ESxSmCIgbsgOPX2d/EnTnkds6rkf519F+Jj+io
fworGcxeQs/Wyb9FOvGQPCwSJp1zX2pultUDE8neovx553yGJ/F9z4yYMaijAmnP
BHPtlDtkxfjP2bteNFDJnifY9Pjb+AqDDoLMViit8w95PR2yyuDUmbvgSj8vRqcV
0FT5Qg8MPgCYJeCo2cU42uuK+gnKAGijej3mgzkTvPsLLS0A/G49/6eHttqJDSqS
TyH7CT7jXj8xPl9Xx4Zo9eMN6/t+0dQQvWlqvbO2zRIdsGtQw6nB7+k4oFU5C58n
kkICNru7AtUFCUpPjddwFL6H+DXp71ble05yagmNDoK7m9J1MARmkMHNvCRPyi2x
D6OrsouHkH3wM00GxROskpLo1GMoYyaZ41UBcmAjs15f5Eacn3jI4vQeVR6zvhgi
RhHtb4Kwb6B+BL/gor9fgW88NGfYdU+PaiQDSSIYorzyCRqLCix+HVE2boeAkM4F
CPJwsJYVmz9AAiFESco3AGacFsb7uUZZdSfqCSfB+Txcnl55zd4SMd/3AmHiInJv
SPacwQspUdt/Svlng3oVdiGOerDkLZQRU42qJjMs2TQ4pGZkDGBYwS3TwyfDvL1e
Yji2YlKdSmmI25K29Stlykhp+K9lNkYV3ovx5AcbWGYpfevz9j6lDR7ZzuA66nBi
r2X/jO88ned6CYqNpVXqwrGuLGFMtCmaU2Cz0u3z2G3Gt5vxEp9+k235OSkUukcV
o41iGv/8qlAR66X9Pog9YxGcxKS6E9OvUY7Iq5fgucIyfyC6uvcg//TTcGqSAMmX
WMBB41o2nIzaJmec+wRtwkzO9hhbP388BqYzsVu05ofIqsr3LxWfnz+Qn/xLtokb
yPBz957jvOz6kcby9VYfkwq2W5ooWN7+xrgrzBJgEWhxRqRcNcQA+U5hcciBocmR
cU5oxE+FLjxhHHP7cHk+3TcAzuufjMPej4BTxtHdQQpoBoUZm+LLOGLQ/ZeLhcqP
+m04JuCtVV/zpRv+5cWG4dGgQQ1GGF7l05ant7lQa/qbB7ZB/2Olh0KDwbQhMuaG
tfOZjaIzwpE1Ri5A6CjmwwYX4Y+6b4FmOKYOIrhBVRUajmOtBOZDUifTgwBkA2fP
Zom3XuoPdfktBlasg/YijJZSq53bjWs3CWVUzqHBt7HCvLn8kuR8HRBZX2UxrnBG
+QoQtglsAF+Xz6PevbfnrxZ+R5/jizKEWI2J0eBVgUQfV83A3UeDgRFGwxWiYqV4
eVZhOnLFpDZYItv505QPrIIW6Js3XaQUco4Ojpex02QtebKtnCeWotxhW4SIUvJg
NMJDb5JXir3cOpgvnLF7y0zNcdaKT0nNAeHr7WcPCdTixhl6wTt4BCixjpRlXqG9
kvNNnG4WZnrt2wmArmNRc4v46fq9kZ8bg0S8izmiJU4cBZVecvAT3g2kwRPKimUe
rRAeVFvBsA21JmP1p0hmBTZtsPVBd8KSgOmlNmgk/u4CJMohRfqshEToS3R5XGW5
nhx4C4vNU/VWXpdlgphuPmDCoB21HO/Y6TJUJ45dWz6px/PcW8AXWivI5UbF+XF3
ZwGQh0nHbgelHRn4uml3hWQoy+hHhHXQcE69p2eeGfFXFOcAXMkrpHbHRpc60AYW
Kt4CuoYS9PzvqUf887Denkm9HOAqCCtQ7e0rxPdXgYgJw/3Px0glwIuj33kVn3bO
cmowv2tB5rUPcF1UHvb2tkPVoMdBPIJmFlcJuAm/qxD0d8ac9OiiAnmRgEAbQ2yu
74QoSQe6JySgUjyqBsvQS5hl/AjZcE6qFXhyKKowvr4V3AH4iglI+988iik7ODde
8vObt9r1fr5g9M4pTQ+9Ro0PHhQwp3u+Fgt4GouKNEx+YIbUUSZBhFMldjTjINMV
g1UZmCLyfIoU46XQzTb64JSBnZvao8lWQSXNf4Vz1O/vrAh3kEd3hU7hLRFthsz9
ZwuYbkJNLEncrbQaJ/joYCadpQ34PLsVXyObAR4w3imffvDEH/fUIDB2R0bLSIhl
fk1WxqTxrV6cSsifudTHSil9XTQx92LN/V9nULsb95oeI6VRH9943BrKU7sYpg+4
07Yv+TWyKW+2nZcYnN6LUaHl2Xuw/TN8vMxKl9kIEn33rPP6EHXp5AeW46i4wLTU
/N5tmQTTtRDRG5lHknSPaoAVHvXy31T4Vm13WVYBAzQY+JgbEJkEGgQQXtCAux5r
93MqTQPutSwzAhRgesKNcp871um3HYc5dcHLQKV5qIqf4ZVFTbdmigzNVUKtXYoR
mCQMxQzLEHW7VzqP6kZAIGyeS9DrIXzcsxk28iLIQBgMKpiSGSUwK5O4HidHzaNT
7DadbMXn8qgORA7+Si+ma+fUxpDyNZmg/ajVcP8NaBFWfJl+YS5LmoVJuzJMsG8F
xb44zU3DJRWgtllbinXh7++zYp8iv0m6aIlvJbzqzVE=
`protect END_PROTECTED
