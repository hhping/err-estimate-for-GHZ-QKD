`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bf+TenTYADNEW6hg8Wms6AbJkyiBgB8pD2oQypqxgY7eGyR3Urz/zkhi0vwNlDYW
T8ePNONG79toD65inYbch336YpBBJSGnn9oWLNpnSyTHLzjhfAcjrDrcIZ+hiYix
WfWyxxlUwUlnnbwWrCsyQycivd6CF4wtLWs6gIUOucLHTI5MCYhvVauehGbo8Vs2
V3uif+J3lFxeufII1Zy8Ty+Q+NgNGe2gkjwd9XQCaQBXQszfVG+so1XSEe3cYRdb
i8zz4cACMiDAjkqrMfxM7L6B+x288SjfnIPKcYsJE5eRKzMV6biekPV0vmoyk3D/
60fpFhk7OIjYKCNNT7xdJhdyPE0as9IXQ53hzZ+MnhWOUuwRNIDX3Md9kpKatRV1
fCD5yW+Uvtewf/rcu5u22uV0r6tC6ExN06oQZUrg3yeOuvEyrPVnMnREf7/kR1pW
RDPX+g9JjMIkkgfG2QuMU/KwWM50aCnG2taKU+lNNv/bDycxR4wzHVi7GqTMuNc4
CoOhsGhcw8V0+g6fherqafI+p7X6xOoJNGdqggSo/tXM5oXk1O7t5vnpdpQHicBc
gbU0GfycH8ZU076jjHXMebVXdsZgkjPH6gofSy+N1RPjwoLL/aSpNbxE9mVzT0ox
4YhCiPEw/vafCN9mSWAbF5AptngI30k0y7UNbMVf7gKOUsYzCjObQpJGFNc2jGBn
`protect END_PROTECTED
