`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLvPK9bPGRVka1tJG37Uf7/LASd1bqKMtTd7dP+5BkiLki6omhPoaLy0jswYNsWv
5oXCz5ZbUDTzdVTSqNNuxPunT4u2kw90bLj1QWDxw/0D65DI21AOQ/FJ1dYAS3Bf
EH4rDIV2g1D2lezrWu4xDTsnAJ0twy5uqJzF3akZraqpIzhAAnuTLFHkz93i7vhg
GnH4b4Rwq9hFm3Yuw3KYUBC/AM2HU/ZoL12U9BAFx1DIsyevrc2H0L8TTSlS5RWK
cRt+9QtS4ISivrs1RCQU+ueCL+ZcF0thz9Qw+DJO7HN8QNG8iPf//xjcesX6DvET
3qCkN+RKKmw4Hye60F+A+zcnxl8Q1UbhDu7jZqo0Fu4DpsdqhCJMlSVMld2UqGsL
vuWsVTMauDHZlxtRLK6J+HAxkoZwfq24lK0hSG/TrOXUq9vB2fMJG4m4JzLNX6Zn
iELtNcgjbwYzvL9lD9oaG+viTGRmH0m5vFN8hXDOtIlHmDBUm+J4IuFVt5gpDuTc
ThOSlGFwVcPzt4tu1qplCVM1DbPMLrciSrm9W6kF02Mo+NJiP3O/wwlLZraKp2LG
`protect END_PROTECTED
