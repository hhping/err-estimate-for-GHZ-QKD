`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CssUx1kG307U1k+qcweMKnx7BZ7Vl7Z5OniDAFv9HoTEL9tzNnfeOBFROyZEtua
WCqz0e6+SEZj822IesFpo/PwiPpsUV9iCn0iOB8CQW8UhlZH16E5fOaeON7bLuwq
nSt7bizrxnLgoVY7uVpqaDxVx8T3JyJgfSybudjS5wQGTFhLHnaKqvk/zUjoAPfc
M+tOLQfOxBH+1V6/Y+IOoYvinvQVQoSAi+e5faRS7+HQpXiMvEAU/4tLsLuJUC0b
LzG1dxDkPbES4V5c0ve0jn71e29/240B/uB7KL6BJ6Mfrx7ASbsYf1v2p6wP3TYS
qSvq2woqxLRyZePYlzLdo2JWd3Bru83e5AtievYCBBKzX3sl+bMsvPaySJ6DIArs
9gwnL/qRNLTV1Dx8oitS2Dj4SDU3l9oNX0FFd5ufNKqg31YcZQFQvoNnSfDbtGst
+/878SzkcghVtgpWyfVWIB4FHnQIlYv4d7v10yJpGpwrkeVg9IhJ/o4DyS34H37h
kyecIzJMfjgpw0DqEsRDRg==
`protect END_PROTECTED
