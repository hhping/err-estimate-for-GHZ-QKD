`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/biZF0mIPN2UqKDQ9aAgM1EaJp6ePhXBNiHWNvoDUVT7UIl+L6StmXc3vkAgaQc
6xItOrVt2/eVhDFTHnvNJhpDXcORpQLMhollAwrnOVDAV6XrY+2HjYL5MQG16RrM
oYki6R85WxwWG+z4ddvGAF+69iGpsIJhTkXYaLavieVZ+GVZClv36K2z08KZ/HG4
HhR5dwGDRnVZsMwFANytW5cRVBkd8iTKIcTDs8OEso11S54EfE0Z8HUaG5wTuWCx
+3rePyxsu2C0sQ/WO+Md8G3Nq9pPp+4fyaX4md5W4F+NmcFotHLwWoziU/kLxr/v
Sf4YJa4sqaLkJpn+FWgMDn4z9SFHiCiOcub5ks0lbYWQlRWuSy9FAgSuaCyep0V8
v9NU84jh2nucMbxY10hSAqXiHCx2aK6HnEDu0qf8quwEuJFzvDGdQbuO6oI+NeTY
GGwOMTb1Zge/NzM6QnJg1RLZ0kwMiRBLRoQoNrZCiyFunRoAYGnrR2wLe5oQvUqI
OHpkwnHbccRrTjHt04tF2uSAhCPuK2nFBSNSsTIEh4u5fbKXzqGmE1q9mGkouZ6E
QRSva3fSGSXCMzwzRfVPV7wDk5wzmGH7Ob6fWSPlBC86Z8Ds9D4c1hsuMJr8yYYu
AE+oDn7jhQM56Blk8obsH/C+JnZz/2bc/XdpoiBZVERbaiSkZZAAUhWZ5CnTa1CQ
t1yJ/vNK6zbJLkVDc2aZf0ozb0cFdrMxIHim3Lgn4PaK7Il8d4uJdlFdbayFeg4t
WDx93Gtfv5fwxgUYrG217oQdpX9CU86LG9s+aMzybcw=
`protect END_PROTECTED
