`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XTF6LnMrdUmxjwrzSV7SEj/eFd1njNKsA0gOUQrZF1wnd5u7mBpadahxbJi8EUst
VIw6oEM14xDdwec9x1un+C8+2bldCE0whumlcWEJAu9WteaZk78jcGzlApRATd3x
AAk9j39IIv+6MMYd/nStVAZim+pcEaCzJuifjlU3wiiKTEeKCcNHk4jFxurwPV/X
6duyBBK4iosaLL6nMm9QdVrarucuDeS4YhBA/jpcYDfVZee59hTxULoSEc8704RH
r196+a8xhWfkWIL/UgWygPeXlr8XHWqPeCRvjaJnGLWHmbA3++K2ImPnYu8E8pbs
hclOVbmOr6hcAktf+OkPMwqdVvQ3rMaHTzzjOreifwXomybkDoLC/Hxj4sXT4zsN
CXr9F/kJ9zp1xP8LUgcRLx3uBJhHdyVHbtbKeDyNyT63TW1jXql+m9fQdoezMYu5
iwu5aTjn7/xwQa6c1++nJr6HK0RlEft7BNIjYiGnkl5XDRVDNV8OwoMqBtfhhOdg
TxXWsVjqKHZCta3P9c7JwA7EXn1Rh6rF/wZIhxOz5QK1+55vANiKf+Q2REt+Kt1d
1S51bhJ08549r3+k62bo5zt5UrekdeXxaub23kqyy+0IKrb2a+XAKu8kq2zTVkNK
x5JwSj6wYAKeIs5CzWctKSxOsV0fZNsFrPQ3FIaSt3M2aADazx0UGKDsjAOd2Akl
UDS8dvPuXD9tMfg0Vhej9MEj/vayG1k7XMGoDOTlNYwVEatBALXtpuGqTwV1+8Hu
Jy5DD1DlR/9iAXhF+WcJk+rEHt9SnZd/Dy0gQ7780U63o01ZkjZlXDXLEoHYd5BP
M6GdjW/ghaNQTK2n/0z0PFzfkX+ecTnJhYgvUDT90WvEKv0dpwfgndetztkLemnu
8FPuuilu/8nwH8AF8YF/1kYMfVnU8dEor0fUNRCa0sab7htQazSQ+ZMvCcIGxbep
Ya8Zd8ZAlhoLBJpH1snNiCl3fS+bptG/ydF3kcYziczrzxQynTqYtiMsZW1Zm6ea
8WqhS9CxyAcmc7ltq1qjlM7wL8iEXl+e2etV7Bz0sOMxxvHepaeRkoeolzDfEErk
Eh8+qPEc2h+cIAmtvcWu5g6KQfSb1g6yEdxgn7Z/lF35GinONWpAhtyTer+V41jA
8JCQAJEGmZa9IEJsMFoIhCK+oOeKGxz0SGWu2Fy+Bc58qszc++Z6YQfEUUopzahh
bM6jjb3N7FKKU9JzqkdGs1kepRtLoOVq1qaNCZP4hqWgZFGh0wPR5F1x+MgKc4FZ
epNsSP9BgVM/ZCzcpmS+ySHhdA9E/8/NoHDCtWTS5MjZ4iKJZQQJcSSkSGSG49W3
21GTyzKGIVBmnJ8ZxS1FwGKGeKTVUUga74b8v/l3AHyz6xAHzeb8UrvIejNa7xiL
4ORYD+vPU1MonEr6QMGR+ci6B4P55zFe2Hbl4XASNGUJBtyKO0yjrZVyCsPkKKtX
FVXSiBSIgA5vnbkUMG56lx0uNwC81u9PXq9W3Ssb7ZrEU5LbuOIKh6ehcApep1sq
PCWFZOWFzBEE4dG4zjhC4Bu9B+TqFgd13rBC2rCHrI3sWBrQzNXEO+GzT5LNak7p
sMGB6t0hYPxhFpTXyI1MULDTKh9nAJC/Lt9wuaZFnf8o2ZAXtNBPaHQmmpZs9Dyi
Qvy5zRBl5BeZny0IcEQbpUaKWZmgeJe5U5/BWWkyBK2LcLV2TqUy7DnqXPHOu2/E
kR1E82sTvGLLldGxCekk/uUTZYIp2y/M/b5UaKC0G3hUr/kxod/XvSmg1eqkEWfZ
PYHtiB9/zqUveOrQMelGwNpIiWzzcYIGlnuiNn0/27tSDPQmHAHMPOKHr5RMLxao
XvNCQz1+Dbw8SzxIzIoJAoRN8Iib8BwIZyBMoQVAnLnQJtHp3atjePAvuTvQt55w
STmtw8bj/5veFfgXlGkMH9DEQ8gWn9CMmEC3h4gTmIfsw5TUJe8j3KPrMDm5yttv
QX1X65wCEx1MnEQD/o7sB4UlnV+gZMwQG/Z7lP3h5zV0l43ob9VvXmvlHHRUTrtD
U5My3WEvaj/up6oz9wMsx3yNZuM2gHuaqfDdiPVEp+FIUWTeJi0X325l7O/qKMWE
tsHvW426q/yi/oJBmSgdPaNH/Jv/9vqkLOWICrnPaC2T0GtDxn+kyZlj8TZw+rPK
IRRYOueQsGxD/rN1KT3BuSbpsyxwfPkqVhB2Pv9ZhRNiy9G2vahLByBDPnIMJ7oF
JzNOSh0spwQ4gz+JwIl8COgrUXcNQLPhhOEfOSRPqn6cC8sJeGTkdP8dA9I030Jo
wLkx/i6taljSegnv7AVIm+u40hfffsd2GYMtkW2rCfUor7TK9Wi6yeJsCQqeyD1v
IGpKWmwT8gUGqHKelnk2g3mvfC8KM0tFseKG79Qsm6YdwXHH8LC1df7QNnVcGxdt
ZtZ/CG/PoehpPbDKNFGZPpZmusqRjrek9sIIM5G4xg1DUiI/1YMYzLCcHb0nlp55
OiIn80l4shERD10DojwGBUtgrU5oh0i7O6LQ15o361KGGZiLxArAWv3Lq9g/xPfv
TD4lphs/vJEi0ktvQMIscaPyWW5F61Ki1mT9kylWit7ygprht3ifiZ4TzRrZSZJP
vm2vlfxEkVgSAl6hvRTd3VZKuxaRt4bCt7Ow9IErNpM=
`protect END_PROTECTED
