`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tMq5MWWxdtftm/q8+F9Z/d7FvE/252yLXjLgSL8DjbTrNfNeNyCFQeu6ztQ504S7
V4szzOGVQMEcq+3GTMCp7u1MyuJaSaZEnuYPfVFrEE0NAG1gAtAVWdUPQRjsGuUj
/+p/vPbVMovTKd7uGGw5qWtNXMTKAvEE0kRVuk7bZ7PgBk7bJlK+sctbbKhw/ZOQ
N5wzMLj9cIFlybD+Q6pem2gTl86KMEpZXMz5ZMiZoBwqSj2NsiirAf8yBM95/RVQ
P//XeJ/+9qylARs5NDIuX1ZYse06wtpGvxrDYZ96hqbuQKaPnvVPJV3848YluFzw
Fnz8ZYY+XJT7TLjzrvc+gLIOy59CrLC8fPId9x4JsVvPr+3hDYrIVmbf1S15eomg
gigdOsrgFclO/xfa47Apj+JX9igXQ+roC4iILoeoxLZmpe9K5bVXAemB4IhJ5OJc
9z33NTuu29+WXPhZ48F0RFUDPjlR7OvX65WadkWi7JwbSJId5qqn+Soe5Lv0IQSA
lBMVMkrdsa4TANNkkZPM2Q==
`protect END_PROTECTED
