`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MEyjMVCD2vOolti21TVTJeFKlZ1+4JWhm7lLthDgn4MCdtdT8oXZ71fqxcdd54h
XD8glJZWXbXxwfHi5d8fZZKvq8svcUI/M03j7itW1i4iWzRh1nVkJMZNeWDVOm+T
mnOOheaUJNBjcCgIIfpqhyOex6CzTZLd9Gv6/XeEir/Yb2fmsK6QtbCYudY4z7zj
cmgHgkcpZ/xZT3znkisexkERFAIhTk0vEZumccu0hkYjRwTfujoaaXV0qdnkLnlM
RoRZ0bWaOvazjMXsxj8l6hujo4bRlujhTnfO5Fwy/j6zRMcI2nprSzlzEdxJgJmz
yLhXsFw2732e+hXR/28anNzPP6Mtb9llKykpA6qIQlWR6Jsz1zldvTmNnGEqrQgU
/POigNPaDVVRtqq+bYUnE6fnlWgLPo8eJmJAgXpl1PRxHOokQqW/ClyL1jz2D+CE
qe8cQlvK9cXttJQyEdQMBg5Xq7WJX+HxnAKzQtDBJANJxjtpUXjTXZHDOzB6J+5f
CRoOHXL0jcQr0tRtAAUkPqI8nNvubj3bryib03LBEaDRwRcY5bEzuNs4uiG9unfp
+hFKzzZ7IuLeiK0u4HAoYBgXH4TGRHJFWNY6jITN34TFHVS25xWZJpZr+TAiJazK
xTR2TtHyW7HNL0jZVTO6KMPSnq3GVNvWiN7JsmTvndZkbPBsaH50Ew19dG+gRpN1
5vsOjDGPibGOkqpBqdfn7a3o89JV6FC0/Dqt/iDwBn1qTrAGJzjt9ch3ISLpBZxr
invPEYtjSgeagW/U9+hV2OKwpgsEMtaHMmK4sS2z9Kc6dpN9P1Y/aO5IEQRS3sra
OZXGSsd9JRTHBgPO/ig1Prps7fSIZcRHFZYIW/SDzSZrBBO7jKogKYenRSr+gVcf
ocy3KWQiO+8vWO8PknxWKaX2JmRAXbWIKM1mHeXgzuGeyffjIrl+ZBynWZoL0cDR
WIbR0sIQ5NMCPhYdCazQeZ7MeQF6P4QocooOZKLHW3SgukTNB3j31hA1Rqie1rUr
AviYBP4fkMBm5TKLkwFwj9f347ic01u3sDe+zQe7sqpiqkmMxK7PkyUmjjjIapWV
x/hwBDQXi9Hwpz17sowb0Abi6JFNVZ8oH5IyDan9w7y/7TJCvZa/mUcBPKymPvru
`protect END_PROTECTED
