`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6kXcHhpNYA9sfS0973xrsJKfIGdlewMk4UucKoT6XDfiC9GWQ74R9l19KbeEEXb
1hBvvSJUvwT1XxDE8FH+SToQkHQKpQaKeqnIvZymvoyBB9QGsKqyIF3mq5TxYqtb
IpUHzeJjYcyyigQb0fsdjs87Fn0utyrF1G7in7Fs5G/ygpTuanqvqwgyx84ts6fM
VzzhKki796nlT6kRh7cE7BN0xM0Nx7iOn/eWIRL0PHShOR7IidDusDUEQ5zNmRmH
0yUKuicBLgYyuBJIl7fl7pIeDujY3cnzyIHcnO79u23YGXiw3/EeLzeLDMv0W+ZX
cG+U688OGsysXRkU7GT5yaDUe/eoPPh4g/01gCBAAk333xrGa/iPJmIil5+Bqf4m
/kjHQ2LzzgGG9PTnvO5YxJK4E4OS4xi9GQyRy1phPfzTNxIX6uBeAV0Ts0ApLS+G
wiVKm3muDwqLm0Az92a1CZEmAD/LOUh2cu3gymd1v5ksMJI6KD8W/n8dhhYnNAuR
XlLpLTZAEFvVp3dDlxK0wBhR3e5zV7oSOJPNUvWutwKyhtE9RpPNsR0ayq/bFZwc
8y4jHqQd2i042C7+vRljl5ST861zgQ+3QfLCPcJ3Yp2emYkcxo30CNUtSHcaGX2K
dU5bhgRQfprLzm6EPJTGbfnucm5TK4T3AgpnFcXGj8ITnVxI1sMFpjaDCFCCTRe5
yMZXCCfCG8WVZGKJLJaFsHAsn4qlSYjxZHydrc4J5cRsHqxoIZyOIAQMTmqp2X+T
nDpncH1RVl7JItZSti+Muyq1TopDLGe5ztAOVtaek4tOSenqArVNUj7ayvY5Q37S
uAgsNdjzLsbHDQS38lEg8Kivad0LMtjsX3QnhWrdzf2Jm/vA8T/iHjmAK2PZKSt0
R45O61hw/uCemO6dFcYYio+FmMBfzaIDkhMK4qbyB1g1clklowijzXXW2VJlZ/Sf
+/0pZQbJnx/1bjhBkrzpOGsQHh+yq2/m8TJpwWAe8TrWDL882ApaJQOdoEC+0++W
vnsB68uqCQ6sNnOgqCtODnGgvhbYG4FWjCOfj1c/izdTL7CUTHf4QIXd0WvoFZwh
+DHXLrGPweU9E2CdE6avlreeXg1IwuT7Suoa2pur/AI325pfgHJ0vNnoBMmHyY2z
HqLTOoTcp/Hm20BPG0Z6B2zEgRBL/xAA4ly7gl8bLdBM2FvIPWUduGCEwK3K6Gfk
Hgh87i1YbQB2xo2zUsNPQqgzEfRcTxrv1GxNgI+vECdRPJKc2mNPWdrhAm9OTAW+
039pr0VC0qvcgBABEF4S0oS4/XVAjyoLynLllhM8IrHSeAO1BL/SS5Xr+aOyK3AX
oTMwv4a2IwZigrrdEfqY/vQ/m68xsgmwopkM02zv4TyodkMFIcv2wJifYJmbvR/Y
ahjfqnwpWdfAZHIcP72TwzTVjlZLHbVXyZonqogO3mCMSTZ2SvPjyTRNs9ECUdbP
giAN3MLGvBHNulDmmLwvJFpUFx33Z8z+tY28BPGXYRDr5ETh2U/5DS7V1jbOR5vI
2aoJhfMNXlBoMi318qDwDWindkbdL04H0ZQijdl//sXzpIZDrmdtFeBTCm6MSWWs
z74lgWbG1uxQ1McjTyv1ivF0aBGYjrPpUm8DADuyCP9zYGRTmPUEEnXea/O317U3
9cVNp7xr8gwndMG18Bc0oD3aYRlB2DXo7GjhHhhOcaX5bgKhxfcBrsXl7WyDLC9i
sax9eXvUo3j2B8TMXo4YhcnhOOQN9/WSwKNaWCberHqEShSyvuIaMbbWlsMLIU6A
yxmycPRs5RkaA/jHUl33QtcijJH238WuPoTfwhxm7phe75kPwkmef61YXkBqPwa6
hM/RtP44R2699Fb4/lg7MJo9T9pUPrUDJFbGuz4AxxR9cMkGENH/eIRJ2thAaLzU
NI+L/Ku+9IUUT48MNIIjci+/9XrYUmCzjpV9jnBZcbk=
`protect END_PROTECTED
