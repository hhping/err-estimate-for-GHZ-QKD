`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9aGuba9/E/2XBGiGlT67CEc4twlmWxeoWxJvrTocf0ApDz+mT48GOsMaXd/k2Ed
A/QW5eMI3FO9jRn65FT+Gr7Kky264ifNU1oATphEdCc0zidp1fD57cKq4ReYa7NE
PPmFzrkbNkXe4mEcV5z0bljBb+68zW06mVqAieNZKgCEm383cE6VX+/WBquVhcO5
5OGDEvBngO3qeSo7xTgJTR37Lk0JdkYQ+3pGH7398FqNtaVrlEDHJFhb0+Qfx3Jb
bxb/mvy85TXlTqMLF58StfKaSGaVir1c3OU9h50E2pBc1cNV8OGOtNYPskeGlZed
KIfF4U6DmHf3UYQkddwYJ34UyKPSWDD9T+DfggqfVHHaFQ1Vn7PF+64bZ0sB4Cwe
HBIXdVrd4Ly+YvS4Qxb4CKcoa/MnerPm/FsbSO99IjSnvNs6n7uSf7r4eeh31KWi
UAtVZ9UcPy2rafr43wvc39vNXRCTsLS504r/mRWIjIK2RNRZDgNyh+GDhJADNXqH
5CbgyahBfQvs55c1ZEsVkMsUzsZHKVRJ3o2GFEBqCKynRSiiwXdnZZMu4kjF/CVn
/40hTP8HR061NaM4xBsYgfFaPDd3vVTcfUZpD5B545BwGLah8SZDlZjBKH2QEuYS
8vYkR6KC+yDKKc3A+xWXkciaHePDX7T5N+KM7SJaoCULT1goNYZE8r7GMdFzH0ck
as4NlRTZWjl6+rpsG1IhA0uDMG5xbb+yrWl+Wmc5bGvKlnprThzEHiUrfGLbX3iy
3NRAU2jRdhyqY+SIdwtyGViJrvq630v43Nje/9OVYVQWZKg1yTqSbvK4NRJHIAHn
`protect END_PROTECTED
