`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIJs5LE0c2p5j0eP24cuxoIxvj2ftzuDcmFzjIbGhbBvexu5/CEBgC63ZOYGDplt
uqgUoCkdbZq106csJDx6g/c6jiEoEDGJSAtnMEntOmUwcb2c+DVVAOWtDK/tdjlC
NaUBcSSE5LkAdDmv/R/hrJzu2qjP+5xHJmRBI0T9uVqEIU66/dmTSsjh4SJBBs+n
ZGw6EkkrzhAhaUArW9JoFMoU0H5pHJmsT6Csam2CdOOWsZMGhmpaqHicZRFdOcGT
fRdFe7fYvKPU0sh4ZFYvYZGQhz6HLKy00CfCVWyhRE8P3EhliO6vLkWbmsFCW2Qk
B4p774igDSNlS3yff43WLnci4CpLNKmwZUVc11kKiEDC+z+5DhNtni2SvDsT3e4M
l/bHyTbOHjnkYZOmAlYNXW1aMOuVGRN5m4zp4gPalHfUQei5O1RsjNjdhoZYRtV1
+32KsJuudVIy+By4rWcCRIStiP1hO17QonGnhZw7I4Qc+jaBTmFH04Mdq3qLti07
JHaurEIrv1lDeAB/SZFxpkmtvYzfclf/40gEx8+VsiI=
`protect END_PROTECTED
