`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3w0GEYfFw/OOK6Mioi8/4uOQPOdSQzHzGT2GEPpXMjlnrAXJumcjk+DkIb+cspY+
33jwiC3D49mQfmn71LeerdLHj8wm7wH3XWkv4svN53oTP+2z1GoJH9pyS3gJonpd
MJaagzaikRtfjZJnk37dzpHL445d3oY1209cduKbnsfaL28joeMwz9bbg+eK8crr
HXkHPscIQ/rPfaxXpd3BQBaG+qtyVPoZD+ze7aKe67pPKphHMJdP2hR/cf+hn2B3
/G0d3YD/YOIwxR7BeMIfRiu0Ye0oAVK8AyrNnR8v+0b1jPF5krh4UjgkdaW506NP
jwSYrigZfA3kt7HIYRUH9bS6bBuftM1dBhQjGUeaG14Wc4xASis/mU0jdH+7HGEc
cRqgNLaTuQiRkawmt47duXkaZupGvsrlcCBrQKjhCcAydO7q/7qK8rzonP4tw+sy
c77ajP2WvPuDwH2GjF0POQ2iE2RvLtpVPzppV5U7OBSsVyuH4anv/iMD2+jJuLKH
6PqDGYjiJ9EgL3k2rC2EUGTl8214LLKfcV5NAXOuFd589+nSvejmQl/T8+7YG08X
9My3xQ417CptrXuBRqdrqjPEqgia1IGWLwAb/iBvKdr9D7Uz2YW7oJSGbp5xpYD9
qw/mX//bstT8hUKOeevsEMf2O27nTX8Pj4DHeZi0vop7SeoexY4NcKWAB3vZmKmm
JPZnuUxs9PKYImeBU3w2nWx+3eSq5ubTelI3Dq187e4=
`protect END_PROTECTED
