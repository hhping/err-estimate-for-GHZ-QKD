`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOFXuVQ/RHRV+rAKvYg+3Fls4GBE79J/y2+N1SLFYA2Dsy6WR+UndZ2nMy/0ut0X
Fd1mnURRpN/TI8hDRIXt+20c6FgqPlly20Rxeodmf5tdkf4gtOGzKTbMnZMyP0js
FsbzUeLPfp10fJIOVfLSQXYLOm8ohPUhQx/vRmdHUGEH3R56JU51PsiG79odjS/p
igYI8rYQuD4ZShIU9G5aMYhWcY+Bff+61u4o2Lfs+vM+QUQgrgtVRyTF5T84nXxl
ApH2yBXZEflLNAGdW5HQFPR2Vn9pSseSwnpVAF6CERH7qjKZfETxaX/hFu4DLHBD
5QNZEx+sYl/paIYPCal3dmy0OULyyUrQmz6mcxZM9fMXM8xK2rIVlp2B2wcq8Twv
jOnH5tcTeJj0Sh4IyeJsdQ9fGDfAPFEqRGmb2vl2rtKR0dcTumm/e75I+6iYZXWZ
pvWMcqMk4QHjY0ZgQ4v9/0DmrkHqi+sSdJtwAe24PhA3mZV9jf4Oj0T72QmfTPiL
HDdaRuh5ou46xpJDaOcrTgwdWxIAVlqBzfWzUBNB5gmsJ2AG0f7kiJm3b45UFKZo
ns5mc1eYsamZcYMjCDQrmB4pNFUzY6nVqyffcG64Zv+9ytk3uDjCrtSktO6yJeyb
X40KafB9tib1RjPYfbM7BAquvbhSzr4Hj83xzLbriTJys1uepht2XHs5C2No7jOW
BJ8ic1NbkK/SLOaiJF5gbViLtgreyy3ToavaoK3RDKYf8Jq5jKscWRXc5l9djf05
wXCYh0Gli4y6ez+Y3fSWCS5Mj/GMj9Xe4wwhfGFcHPJLGXVB7ipkf7bSQcnlQbaf
MuUL1RTp8hOFEwZaJi+s8xTSxtfgCqTl9KWS9SFz5JApCGKKM+JIV+45L6vFr0ye
KgCeBxDozezRCyCPj6KCC965HR9V5TKHA09IOH2lVrO/fP8rmhFhh/1Rwv9Pyy5h
4ZF3eawgI0zl13oc6rCk+KwlXxp7P0GokjaliYx4yw3L8ma4KPVcZQVI5wx/iV6t
pZHzV69X8+Id9iGMA1z5ntOEULVuv27gB7IEFd+e0IwGNf9gDNKZpHR0Qajaipw6
Gi/Mug8i307IWmPBMVrOMdep9cO5/2wKw3zaHYkNLzGF45lq+D0XNCR7bTEOBVNa
L9ofUNOApVGbw5RTqZxlOhZ9NBCng2hIr/mh7KZqUQSJ5AWC6+rxsko+CxZTlO2o
B6lZCKb6AYAstBO+OBALofTjKHpiK0EKQroa17atyLcFmqhFYbHLO6XRweNrn4cx
2Pfqg+3HW/1b6rzswinvP53VAsdvcTtvIwHcPT2E7iNm6BUuTpmUHLJ07kcTYvoy
p7xlGv6bsHMgZGfYov5EFSLXsQ5ZGMPTnwJoKlamcDwmpcQooSvMOROUl/7SnxnD
x0llhv+8t2Kjp6GJK6bhw4gyYx2PDdN+KWivF+nWuXrLRJQiYzz+RDvmK1aPMDeW
WYslsplUbaBi+eejJAjJf4beAnl2ANByHDiImNrlijWmrdvFdzkOS5X+P24FUylp
MSSP6fiKUZ28IImriIdMGEGL5iwNgCYXkHoAKDGF8YcZPDyHSvencLE/vByGEZbz
fQXEFxlcaaQqN2nNWiOaQO4rRgKqjHX0VX4gYvVltYWxnEdabjwj3RXi5XWl0U4z
n1zMwdlHUgeS1c3otBDKFEnxNWgqkEqwUIuEN4mPu9TmntnnleEm9rAtFHc3iln5
8q2VEon0ftSi1I5rivvBZ0OiJsRevFREID0Vr4GWjejHzTsWQdxywpeHy3uBqtOI
erETLOPJPxhDRauMZQQz8UHb8btpQlIFAMvcUeim0ARp1CbWn2wSPwe9brlPaEEu
KthT797SmA7/mXZoI4+ZjXo2nrWjSkKUUCzkFCRlMs/VFB6Y90P0vBm3aod/2Y42
1TX0H/gsyP1QKMDYDQEQhXWmruPq1AZ9CAFvtmmO4LM4pEpj4jpRgHtUPXHIbNlK
jKChDhwyvHsJKzVe6Eo6DOhslyA+i6VxSy71I+j9wpVdbc1nSLxB8v8KwRG3j/li
HjnvBRiA/miQNk42MS5eMDR2voNK7CjA1vj7Kk0GeM3NZeny1uI/U2T5Vi+m3xZR
IKdwgSW25mDQt1Cm7MLrTpntTAlywXAv4vnh1Vp+YvVw81ZVcXcU+Si0VqtN5cR6
gCTp4y65/LS3AI+VbWDkW3Q9L7WPMtgA5G6p3rDs4+DdGeLCRZnQp92Yp++ISwEO
bfNyip3jE9FSu4k3+mRq8furQPw9uPMfxGiiCfcAzQSKSUpcMrzhMsZJ3CY/IcLp
7Dwf8lzqRpoiYk3iV3WWjQqKR+3nBTysc2gk3/c2e34tvMriuaBhXbJ8bpPBs1zk
EfsIshiwiwe0KcY/dw5JW+WENcPvadUFXpp1uxgZVQ5bwnBXYC7JEWtpDudpI2yS
BCbDnm4/4wzbz/FrKNtB6ZkabnfiE90whjUUEl50dzP18G9rc1iPyMnlpZL1YEtp
CoMGfctow2lfPqxO4f4qv5TBLYmYmlSy4/ifvfftm71foZgEDZhm4ZbcxyheOOzY
a9manyl5xKq+5sebn8MxFoj10+v7tVkLSW2b5hZRW+QtKGCXzRwgs+tCFtvmJedw
ACVHeXKju5CGU+B/0ybGEC3+eV01bwYD9clcYXsWhxAl+zZs1q6/lLrlrfGSCGVM
RWAJ1ThzFG2yBQ/YATxTngrYtDRYILTvwFOuNEMG/Gti5JqFtk8/bsmr87ovnT57
ulte2KlQXHWz5HJlQHmRh8P8iSzvBiJD+gH6H3xJHC2zU0k58EHXAx4xChJRklfR
WMgWKVAhCfqa9DyXXwjynnssr8UFVDVnkci44K5JU0p9msjnMXwaJ9Gw/9eWyXY7
HJPJHuQaGf2DgIJwaY6tRFaAwjmBv5MqJrnKRbpJN9evkTC2cMHUbtefPy22Epka
7fuoa6NgvZzvqJNI6VNL1SUQDaWlfCd7ZpetbVJeSx+VLxA6jgARv60PTqRA9F5G
rvkhl4PPs14A+r4e0bVMGFkD4LcJvXmsvnPhz/C0bPu61BH1SQMHYxXZcsKwX57S
GEPANFJAQGk7pEFwqKfimuCY0SySvc5/cpNKEnvNMy3yGxxIMyuc2kMozGQZ4Ukm
J8mK/lKtzo2DoIauPRL1Kjcm/pwiGQOdXwqZCDSPzuRC/Qb4s3PQMPKxbWfE9xU8
`protect END_PROTECTED
