`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gulSW+DR4M2r3oW5FbGvNx+xSomAvKWctm+Jd2zqF1F0lSCzP/18T3k4yI5chwk0
Z9Q1rHHLxoEBsznXTp9bGxgQw2V+z1iU/Sr5uPUyddfwk3EJCipNKBN3j9Bb28mf
wGtVfG55rLu3ySzHtaB8RbKPjDekFwFhUCaCBZBS8vKnHBvGv2qmn9pLmvMpmbbI
cgRLERo0rKan8f83cPfFk0KJM35CsLLSEUbo/fW1dbGrRsS3GGuUGDl2Bdxaz7y1
mEZVqPtb38b487+ujGOGgakrtlk0YaNEOmWSJEuMC35WdqRKbLdlhjG+rK90vlv6
5Z/fwbXZD7F9XoTYT8+5uTIFCBpd8UXMRhiDYXLVsJkSU8xR6cXvz3TrsWWlmwIt
bWPPjnhA2GMbYd3KFP6hdh4Bmrg5BqAE87+m9sHB1diXPNpYXbBtK0z8zK5MP3a2
dXRySwQvozZZHk8GStrWHuAibeTLkjot2JI84S2wR71j0WmPyGLDdEn51r6Z8BCT
GR/CGWSnwqpAbDrJMnox4znKDt+UOhMy0i/JjOKaMbKFcyn5fNqjly3QSZ7zexiI
vvSOXsr6ZpyKUKjBarzWQc1o1XbSp9l3iJqejJtwl2l/+B+LrrI/7oaeQhsquuH2
ISZI4vTtVZfxKV0kVvUng1vYDj/vsmnEo8i77oe6WGP1LO/ZGmrRJV1+2savSnQC
zp397HGqf193cum3PH9/47p1Xy6DD8AhTEPS46B0pxzc0yeEVRYn5R+Sv1MNLc/h
lzr3Fs8YmNQFPePHkfYFYp4wQIpozLYe+q3v6ytK/61jbQ1mpnfnjQ4jzuRalbOV
BKd/dG9exDZzP95hJL0A48tNHRCWjTgvw/v7gVyVoSd6v6bZ90z2c7nijoNzp3fG
BpoAOIsW5Vn1vDMu6F3WD8RjeNuXhEosSpXjgR4gtfqJpEC9h1JsLogJ4RbVqmn5
OqYp9Yjrp1ontpASKqK30H60P0fzJTqzkg839yOEWHZQYfknlf7LOPw0qISg5BeM
jwzzMwREXcROdWjI8FqWcLuNdA3BTo9HTt27v9qTHsxiIqYGUD//VlnQGVGas6u9
kBprPERCUcrMq6fGJCcFDnziSy77XL1wGCGdpmQPU3HulIpERXdFmkyZ4JC9oYdo
eQun9C5MENKeZsgALjNFf2xd7Wamj3TffGJ8T+WpbiEIb2zY2rGtrS9lZU1+HHr/
NygS2WMHgg+9gGyrtSRkte1DzWYgCm/PAOWrRF1QZ9LDvipyJXDoRHrvW0mFb0lf
H+AMiEt540M4vFwU92mWVeLN3OMnSYsP548K6MGlHeqI6BPRuCxwmQ7UooTQn5XS
v3kWBEpzZ+UkxXflr+l6+Z9Mk+nGW/0pP6mAd9CLZCI55wxLOjw2TshQ46w612Gb
KrY4X5NrWyZuiT+Nvso2tTsIW7lxUliDqCULMepY2D3+YGTDogJ/80Li5kjh75BP
Iya2JyzJ9auH6OFBmUzoAshzGIIlLcXfB3oYls90stab9U61AK6TNs7p6PO4JjsN
vAwPw/KpkoeWm8mQYwW/TsAk2Mj5jy4Rmb3sRJwN2QAXHecE091Nnbgo2hj3Dg8T
PIREg75q3gnIRG83CEAZCBG1CJtJQma7TnrG9DWsEZwUO+tzvpS91iRP42LYobHQ
jxS9geCIBf0OUoyzTwCFrw==
`protect END_PROTECTED
