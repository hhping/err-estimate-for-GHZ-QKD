`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5DGdIiRfoduOSmGgFDhsEcOK7k3xeMYeY4ZDjXtoG9NjOCCXqzrz/Svl/CwNaOQ
3FTSy4w7S5ucB234n2mYSnX6MWMdcEEhNwbNYkTfsN0Jkxxd59SwMMZ/+GrnwBBm
dwpJvQFYxUyZuPd0mcimOQCr4gqq4HtZwDZxBPyCnFy3LdU8nlvis8IzBkkBSBc9
6RxEZzWUuh5vzOeeiRJV2ga4ncTERwjJsQThmnraaHQaPWwKh65sz6JoWLtY+vEB
dYhSR4Ezg5FHZpULE4dEWYvzs63jDu36mhFQKeUcHcxn4ZdFDJzvzv2w/4asXYQC
5yXKcX3Ts2ntn7dF/vfnP/PwUg748ueRAzQRSLxWhUA6c6NFi35pj6XxRa4tXR1L
Mt1roZKi5J9AFbapL7RMiRQina4AMeMJcOQ1EAST5D5JqePyNQWOrRlxQHkNDr0f
Sx6W/KAKQ0yA07OC1IMJUS+ldT2ZR4N8t0debaZ2PBTCqPOixh4gAdmabAVxPRgb
isrPK4Q0mjF+sBpnoKDw7f1tgRXMzefMtd3CDXBymN1mIXAJgvmv6cmspA0vRaNY
Iu4AGTz17HRgITp7zroY/sMk1aKun4KaJzw4RXDrKjFUO/lW3L7OoLvMqrhfHRTO
1Z65QCZBMpfMmahPPFhrsoEzhxiRlBRvOsFoyAbqF/XiSR3lyNJULAk6WuVYm+rR
pl44eWUoZE+45Xvvg5VcNpR1pzy/9xTUXX76ThMuNGqbVWN2snheCwQYAOduNqbC
1+nOpg6w5fbp31dPDySSVBykYzUSQc1mCsaYOz7VpIacwhfe5cjl7s60kHvXvQCV
otLAVYn+BXdnzTJpAlaWIpGJGYK+ZrvV5T+FYR9DN03tEvGEFKIx0NrFug8QrMHV
ijUZtWZm+j4LVkNe2n27P+CANSr1imMzFq/xcqvLncSzAU9+Fb/gB2n1FI+8Yx23
3HHIzhQhS4a6sb7okxapCFDwmfD+jklIsVgpswIeD9I8mb+WhguaP0vQ/40K45dA
rt9R/fS4KWZWjUVRy36nTNe4gIa3oppAyyHOFLZ4ygTskvmXbRyHoblRwo64g51r
PLIMYM41TaLYK7JMexB/eWMFYTMRuw/1JeD8g/+PuLQHiEbMBh62vHhxLrDfPVod
K/PRSrzfb5AWur+G3z2jcOi35S5eLQtkvpQVSeaE/T8RSJC10O84HotPzr+Jh46B
G7pQqmOw4+2a7eOgG6Ahs7IUOndksIr99T+jA7tH0h3mwFeemo7+exxnv3i6rNqG
lp1z9onEyTy3BrnBVYElVP8aBtDp816Bd4EWj4Q/GkvRA9lEyCmckh6L7KFLyWst
`protect END_PROTECTED
