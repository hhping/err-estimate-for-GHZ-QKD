`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRDClZpGaX4MfaBLRmlY+xKLBaqke1qimZlSu/J+bYVSE7vEKnp7UAkJTqm7ZzN+
ZpqHDF3tSWRm82Jpjoc/pCVi64cZFEBADIcoQsxYmsqnJFus4yYovZrYnoRpk4gY
9AgPeXfzcMbu+M6q7CCKrbTMlXK2V38syp8BaYikxdenip9vJOTAJnBQhvDphZMz
0PFHE+kgdnDFWpUKaplrCk07O1XMQhhiOMJrxOWKqKfWb6rSYV4wMfQRDi/Ey5Mc
IVOcit/bOIlBbCH2zLHqzjPR4h0CUu9JE6DRv0uHcR4YCj54+oI1qO1Omc7OAvzl
oHguFF0qkM6Pd4o7TYpTNTEbikd2lhiMGcnzHgV2Efo/CqjMtsvTnpVudouEpnnx
iSMyamWS5+TLZTfn6ErIzcd689nLZWyZhSPx4b3I1eg9S2knR1LkuXHM6siDQ1bh
O5K4Dob2ydvPbQxz2vXwgoljhUd1lZBrN5CerOogSl43SEGOMCwE8z9+V9GyZDuN
DQzW54i9oLhEkY3eu1GR5Mee+QdTuoh1+1aj8GN/jk9toFMcTAYFNvcllRjTMC5V
GcfZGFtR5/vs9ps4d6lG3MwQ+S812gvn9WAKP8d+lZz5uQZZQXbDtQQQIEN5AsdN
LvpEI5qMvSDfkLhLdD0G9wfJ0BURThsGJKXNDydLy5atuW/6G7NJrilpMPJDbUsG
yP8CqoEjOZ62Pj/F016cWQhzVhrzz5ygppRrsNd1YkYRt39s6l5HrGRZpJB22k2/
ZHghoaJ+anV5roCRwIur3KaTCeHLGgJsK4GQJqaakb6zX+xGtzk2BvMjjJQhBXLW
PmGEqPQMWMzf22XxF0WziCNlGJHQny17DsvAVwCxOk7BydOHhpL1MhF+z4C3RE4/
oIMFf7f+pY/1QNkIwJTKT95iWdPRwNMMXfgJP4QINqpxQLD8qV/ssRZolxfqhbZ+
VV2X4I9vyDDQ/Ne45YMRnjd8rZ2w1hBfm+nWSaPUM0gdU/YJy7juEhR4lNVx+zmr
TtddgrLtYKg4bi5ShzwWfDue7Ifm4FO2RjHBF9Zm3n/atjapeJzJx3csKcfyvYdq
Nz2bwEfO/qzPtb4x7pu/2PWUyUkBhl5zyi/5KnkqMUuRl1YN7FY0EkoPNx9RuRpN
tH6DC7NAVzNdoAR9X/0MkRH+q7nyDkCrJICZJFB0/WGhepoMDYWp5889jIvl8LXI
S4aFIdLb8q1Zz26hlUbiWooyB5+4l7scdGzYj2J15WdZYO4AFfmcT+ilj/meiWH/
A7BHyNUZ0ktStDHDTzyl97HnYIgTy6/eCv7dQ6r3nqdUlWv+y13/2FtNKMeciZSw
YemA6eF3GAJH9bNv7ekx/i+46y8snsdF+214ynb8pwTWM7kpAaUwvEOqfwUAmHtZ
AWuqLqRYCw8XLzOzqPQihksbjeUIWa33BJFzlV9o+xeWa8emOK7LAboqmmy9g1Z5
VbG9dqgws1EOf7nfOFN3YdUdJgJTYlJHFADSKX5dtNbsIxTDycHB/ivZX8QO70QX
d+JOxXxXfJ/T7EE5zo488b/gwFiOQ4lUsM0nEPBHNl+H/kz9temM8QKg9kRVlbxA
GZmwaWGwL4tmGqK/iJZ9GY8JvffdXRfRzAu3Es/NmTX9Nepc94mK+JYOZVCwUoZj
IdTC6N2KAoSqvmkN3xYt+8nM7xGsng00jMMFPPeKCwamkolYIfCeZ3wpgzzHp7yF
4+q5N55PUo63tBcOSotXo/5e6dxfO1QHMM28IxQJWl2O8/ndzYFJgPzE4pbS3c/f
t0A7lX+C/Al+Jj0Ngjekz9ki6lX9wkqOdhJwPRIbNnabRImpPsac/4t/TMpCSn2v
gAyGCOGADSSbyTymB+cGSdbtdoKDqJIOWmX4BRDrJfYioXJLW1ZOGEzFJCXPUjhT
J3qUjE1LgmJPb2nuGm3EUka0Z4UrWoqHStY9XlSbHn4XiBmy5zXU6NCXOF+goxJp
+MqrzKULPQc+yPX94S7hcHDFbkbAkWAo9BwpDR/IjuRhirNVXKqc7zZ1fukWl1Wh
U3EFRzjvczfiJYxQ0lPi2hWgFn5phlLe39MrbYZkNjf6Z/s3ntNDspcSijMKfPNp
QmsQSDN431Rh1lb0S9bY7SsU4AyZfNvM2aiE24m9KVpf7YyoCY77NXfkc0zq1w3j
9UYZ18uYNz2UqBwomBDD3UWRwBNvTrfjoTQjdHAyf3gdTasXMNSdVfR2qf5WP8N7
JSVMkEH/tLAitiNH6Cy0lroYOfe0//RqD7vXh/yOFUOW8mI2ai8KBxyf+3AokOM8
wZ5ShpkQZgtOhRFnzFeQgX4q6lyS7nMoj+TBiDQN53zHTScgLjGJQK0ObVvnLJmi
6CIrTrnDppQz+1RHsBIVMQIhPp5j1W4airYQ9gChzVcD9pVc4WKP1wrx/4Cr6SrQ
4lSzPX+CxEggd6ip0ZdtXDF/uw4TXZGdfcMBO2jyoBSVMERvYXYgYkBM1W2Lq8kh
ruN0u8Y8AXVHfCPHFuUp9NAmODasYn/NX5vaos3qrCnOwdsQjV+IvVsxITgCTQE2
8rNHn7/cRAiqUP4Bs2sFY2zXDpkAiOq5Un7sUUE9QDsUOKMRU6hzyD+OtTX1NO9t
pPZhcFS8a9OQPcGOGYTHETrz0RqGoyd1fLGeKXwUO2CkbTYVAu9WmThm0y4fO1/j
6kEvtLuxkbC7y2yzzO7yNZ94uIqJKOMcc2EyBv6bnJ2f5djoGpThwsOWlWJy4Kon
pGcujeNS2M7ZWw7XcsIeKdqECmcXyULHK8EIYeNpOWu2eRICAwIlFh5yHHHxzmzf
FIswL2fzMG39MPx0IMtsytRxeU4aYmz1nxnxPj2uDpuKgsfS2f72On0d+sGDtMF6
37Mjzp1YwVzh8TYp0uJoXiynGpX7S8Vz9Fq2HDA0fKWRctiyYBaHh1ppHIHQxoji
buyFrkosrvOGNE3r5T9mnuuurRgiap1KBKkx7pbve1SKMAQk6yHpuQYqBbpYQgAv
7bKG/0ddR9T3KbG7tn3WNBhB7L/DQvvi+7eY/Uql6etqr3HZOxqTfy2BkMlCrzZ1
PtNki6csIM6b7crPPv15NOlbqUsU9JYr4C0NHo1Aq/MzZ2xXcojICUlon0keB2Ji
sfs7iYFJ8iqk3oK6g7Ui6VenQBdAqydcjNoxQnurxTReZn28ZYCoOsDM/83lSvqm
Sxir1tNaa7nWoq7clpMUk/iOicBRdOwgPXNftELJYPttsBFDld604r/8fbradDMx
+bl/QWL2YF1p8Xs4hhEYn9UWobNL5d8BAlwgsmFlvbNoMcEBiIAuZQm9dRPqJJOl
2QIA4/++usWSK7b7zj0Y8JKQDD5IU5d45HAEE/TXiGDlMvB5fxGdvupYE2O5E383
ejdmw9/c5ISEMmVrZ4Tc3uDTRGIAarREAGFKR8OiFUpjmuAqBe5GBsEqFKoynCf8
cKyN+qkh2ny7zJQySMwt/rAr+OajyPgFKxwyO0W2m4MDWo8Tod1t90ayHbgcv71t
knmAb1zKhBSV6pe4TdjnCIXHZnX+I0IB3MsepnpqMRyOeFPyaE1RMYtHJjSHT1n2
xebWOhaI5wDdq1/yfz/fH7MIjS7M40boEgN/zdRF/xlZhUWiW5rZx/3lu0fxgqwb
PaG39tNk84aaRLPBlbPC6dcydHd1hE95sgX4ZMEpFE27FMwbuhQTajWnJDJ6jgYD
qFeWUvGLLiiwz4ECPsALUcOHGsXfzySern9Wp713vOn8Z5LGGd95KZJ7v5m/wtQa
4ZU+OpeXvrklJRxkBLjjfv5WfosmfwQQ9BjsnWEDHoHXN9spLXTnyac+y34zTREs
Y322Vmx7h16w2nkFn2xsf414E4EtME/UWKh94CyxKpk9imaogQXQfHtlVN9X0Izj
HDK07Z4TltC/9NGvo3U6A9GraBkZxxzO0TH3sGFMMS7LSP1Fm1qUy3PazkCYDV/W
I12sSWg2fHbu+0pOZEo2UzuF9/6Yhacpr0Q1bYXWDg8XmwJj5X8Ved9vhLxdFonJ
WHKSUgA2BcZmdgCHqRjbWQbB9TBrH5m71a4Dnvzw5fIWEVq3AXF9NVK30U5sKT25
+hMLAiye2dH+v23EtTqGI2vu7Gw1Ft6AQEUcAKi0FdFKWw9dHDYmeeocQojNYigC
bnP0Psiu0O55pgFaxDIMnFyi+uR2LHQTNTzOQTJKPCACXU9yxzU+DluMGHWF/8AO
RV8QYvghfe79iuj9BJUc4XLhgT69n5SbZDEriSDBZhxw/vlF0qx3uWu8lo1VGZXp
GKuQgZSCkfgLGT10ddrlPgbu21chsr+hlLbfav6QuYwqoYYR2Jx4YSonWBOzPhc9
VCqItcKdCZZN1Ar/EyW5MZ80uY4CA+B0zu25JMo5715EV0GroaxzRchk0X89nzE7
Og2KW8do12MsSGP2xsxpVZyTE317pMZkbIMpX3oSPofo/dKmuEeX5XzcsKAhHyDM
eYF3c4eQ+hd8O3t6D0B5pO8Bigk6N4nzlonn7Q5jWBbSBzqpQb/NjTeRaCZsUmUv
z4pfUAmi3YGEYHTJ5SbYaYU36n58RaxsKWkmSAPSvtoWgxJcXjHaRXf/UaWr47yQ
phZf4Z8WZnCeMRAigiLDMfqC8G/MNCrs7bDzhwT7EzChQRkQ82Ki+qJ7+9h12qmF
3xd9VIYpz/G4P6YleRBe9LxH9ErMK75/+RaAi7N1nnGwAMqlwsQGu0/d3VlJxyoT
l1JxwSaAkt/WLeEKqxG8v7GL4U960Kmo8lDM06SH1zbxTwPn6OdoCz38EonhC7y+
ynpqkxCTj19KQ+6/cufzbsBjcyPjzpJ8PNjntDfJbMAZ0go1COOfQ7qk0o72T2S2
vpV//M8bdDJg6vmE3m495Y/a6QPoHYeOGX4ZA/q/aSBe0L0r2v3VNCd2N9Tk5C8g
YNy5oZPRG1z5o2WY1n7wGUvmBfe7SCax7B+o0TqOwaTbiRhp2fculuKIsUrJwOKO
IYuJ15ZHeNX50M8a++msFrgHN5U6MzsSMnRJAolPZXuqm+KqWoyK7feYmS3ty4gw
92xZmzICvkdJNRQn4ne2Cv7H5Enj/FY4evwNWM58I26rrAEtXvkz03IFu3J0CP/+
PmRYxLyiEPYTVhow8kG6gZstWoEVRow/p/0MLUK5CrE/Lx7nnDEgagO2CcrA+RWd
FV/F4ap3PJ8w9prtx1y1UowG0UhtRWIS2WtqYegING9aVSDilk42eVFY2d6HHWxI
gpr1f561pLH3+KYegYNhi17zxgmsWJ/D4Las87uLN5zP31MfCZWbiOKs4IvjfFxa
2ZRn9/+CLQ4zYHEtyaZLjH4BE1LUjCNY820DrGX5rqOPIc0aauZLC7wMT3zxVGPa
ds/8ujg1yWsmus0g90dijuxcccRKJbKVPc9G7E99GCTAwWnjC2myitROTSHc837g
6DqMhrkLBMMQR6YVSUc6slAr3MtrCKYHGwY7oG6EEMRDK+HiOZmg2BymwmRvgFpY
74hz2CQWxlrmwatmCCxpB/0HjnfdRA4NtuBiPn6+ygOxt1apapG8n9v2QSs2MToD
1nvyK52jSG50n5jvwsS13RGRIVEfs/vqUflNPpDpS+2+0gH/Krf5ZoEMMpbabAYm
2BAafX9vZSgI2m7Ab6gixNuHjDaLu5GB+WOcd8pdPKPkQ6vh8ZQKPz7OTLf3dd77
nAia4ObLf0S9GoXGUr0iMb0h0bAjhL335CVz5FetLbLPZNPGMmXvg2ogc4CGzEfP
j/MQCdi/LF9fTEQ+/NSIN3SewDg8k7fY0QB1S5ZGIusBdKcZBoK/Pr9d9F2NsJYd
nAymjK1VdTjG6PXrVKsxhlP0zrP+gY7t1MUo/GAndN9nWvMYzl48nUgbqSZvoGqV
orZWz1Mx8+JHEUVYpMpFAQjvQ7/lDuDIJTZ2FcCoGwNjraeJhvLZXaBXon94ufFK
rqbwyPOMJDVWVWOq0XMW4abm/DOD7L52TouWFYy+y+C7gbRFpoWRqTYq5ktvzxfS
1oPTm7Ikmw5WT0zLrNRbrrQxgIMgL63hJ4CA8fzFoSjrdwloK7gSCiltIT8BNyCG
FsrC8YPADwm/Z+R07F9KU11fuVc4/K8h8v/kjh8KgfHtEVMGGAGi4yCv6s6L/MsG
39PgI85/tVgdjeMs9Rlhy8PkzLWoyM5O7AL3HzKUFKNVK3fDG1jBP7W1hOUas58c
cqYogWZOYx30jheMmx30XPOJ2P+iK45X+Pi6yBaN8SC+b+VdqmxoaeSaZDWyWp5W
DY6j8E1O8lFegxlsx7GAjKLFF0QkrxQuii/kOnJ7Xy+VJk7A6YC8WIXAvm2XjTMv
fgApLy9pDwLTpXi3H3jctuFO9na/6dMkm3s7++f0IpVU1sspE3fjdU2v3p7e7+bI
Stdw6lXzMxV8ee/3S7aEa9VXBA4qj70lI7fLnTEs87TkXn/EsmflB9dCmdWA0oRM
9JDF+ytzMoigmenkT+1THpKjyzIMwSOKt7C1B1U7pPDqJLledgW5pf0lY+ZCgiIx
DVSAmxxiPoeEbBg61H8sa1jByUGDA2nQanCFRE+S5oWXHkJa29HkhmdOKr4cM3DU
oMo5QjrfRoiC18eTqAysLePehUNov91KbRyjcYjsf5MxJvtzIbYvYl99EvAsDwKU
VJVNUxMIWkUy/6Sirezo1SDuVhsfRmtcCdexSRJAoDrpht6CQ/g+OJAIWD+gLGDM
+7BtqcwFwdMhlfe+voaMQgc4ihwg5Z5dYOeTtElItCWYADpFgmlUCEmPWKVR63w+
Q+t6dZcbHfUYU4Ov40ndZibqcbvZv1hEybSff1P/jeMZ5zWy40LqM+xvgWoNxa5g
S40hXL4Cu6dQEIulOvGtzitoUIPSrU4k8gQq6XAFbsvda4l4+7RWYdTWF59YXHld
XznbSezkxs2YGpdeLw3RB3Ezt0wl5ucqHgi++Ca9PgvqkDU5nOP9egQqmLXuGOv9
hd9k2lJa4BSagZF6Q9JKuPSM3nrn4g0nWCYauiwX4O2CBqMq7Q6mrWEqCIctgwTX
9NJ5aEN+5grfn62T0NRoiCnzk0dMtYkuoGW/kkFWuOa2j3bP+NJPfBrnV1phgLyX
s4+JQuGHthuyrWJOzDVVH4QEW31UkdFTulu5DXh/CiivbOhQnZ/IufS/mTukxdob
ZsFkVbGj0/Y4pV5DZ7PgILeKoqgcQKF/yhMiGGjz958oqqqAFym+WQ8x62qf38e8
TAae0sPhbLrlmWUWRv0xQMEkuG/8vEsu1mEnKxOfk5N0fvkcVWshdURnIKK+Z36l
2tLOfm7Rf35NXhIAW+hmvyWfNCtGx+8p0jXVaCJKuArVN+i//aw8E/zOGanUlg7U
DCEGiAgp4sZ5tAf8Z91HFfpdk7Ssd5umYXgMT6RDhGWtSr+60Jnc3p15Laekd/Dm
09bkvXKRxktCSXjrKcuiBsQype+OwbP/PqXFyimyl6Q9CDksnzg5pVnqDrTM+HL5
1/M9hw0OeH5xRHQYtXIXn5z88cmmC6odxsbeO9BVuF9IfVpwa5Tr7eIbaextSuWA
mJin57FsFb4rl2yBmOuV5t1cc9pIfC8p8gtyn/cdoS6k5cpkvO4K8pTS8Ve+2vvR
F3Y/o9Z9l50FXsXNJrM7ort28YISAJYKO4r6ca8Ldv0g7gNZ30KKHqQEV1NXQpLQ
E09J+ur0Cj+51gcnXPKhtr39Upo6bGv+L34spyUm++TYlWEMikx+6zn3IZ6hW2aZ
6N8fqF39htdNGbMsdhbT68lAFcvxVHna9nU6beUVg+q4DshlPNK7j8N9lw0PxpYN
GmpYb6b2R/cPMfi6xmR8R82/Y4uLvdfXZoMhHp7pnH38nA0ZjLFn6vzk9UFJHLVW
CcNk091sjHkzpnRHVbQClx+CY0nfAXP6NPTpAsQp6JvNk1XKOv8wZgPHFHqqvsFd
gWLzaRP3uSV4WSEwW3kJugxHCbZG3giSW/RS7ibUOG0uDnxr3NlacuVjAieDhv5I
ha32C2CfpuKpgsM8U+lr8vzqY68WWFNDFF2Q1zL1+bVHjOtmlGz1Lrza29cZI1IE
RevQSf5Vxqkp6E9+2eeOwrMrTdq8Ydvo5W+gcK6jxsWSoHddF/guMUvR6XavGgek
u83LFOuBTn82yd4alOkLgGPBLjogh6FlkT6dmYLEu5fZFOYPMKEZ4+3G1qqlLPYt
qCW3atVeuVLaSzWtfJn6wGWe+sBg7PE4DHmF/XFpzH0JlrRFHwKIjt+WY+UiuX+g
ICzwy9Bm/8pSTkg3u6TGtwOUbxyxMGbonzqOJ7ptqRh9sYuQlu8z3yk3ppPzkWpG
VXhQxw16oZdooO2JPYTWrGU8UQH9rbpAlH9kbCVo+NQzk5cgvMRLZAuCm78Q6tYd
nwqnh3aqrpUbSeWKB/pgIDG2DGCQHBO1Qsjll2utPE7ZG7pYUyCXrqoFAqK8a7Xu
3iPs1vi9KP3nJrdiJ4xLvMWioxhEOZ1LY8o4CThpP4QlT8+rb3O18yw/+Em+HUuX
UQ2iaKa3fmYLJZQ8rDZlnSChIHU47KqDUNhdcsa2FaZKKoTHUjciWlWUxHhkfe2t
Gj6UN8NG6lt0MYOrVSb7A0qazFJC+u0ftGFLYpMfEifMA+c9I1Trka1yA826AxZe
XYMcBcJqZBf3g8dQKwCET1wX6cgqK6OXYYPZ5RUy1woUfvKYo2xJVznB9aZPs6hr
sqE56i8i7FQbrM2sdhvsvw4w7aNN3FKIySHVt4sUogYz5vvMxU02gtph8RpLygCE
pjLqMlr+edYlh8ZLhtdLxvYJ024g9Kn+3VXerk82SEuqa8CzVhlnSaVPpQ47+4x9
QXQZrMiymQ7VzjhMdm1yAMyaK8cOVn+eQbAmsOPqsRRM5lYV4/Zv6e64nkNM1dwV
0XEAkHfujxyjDejht7dGqMHOHoCvCjU6L0yKwM5r6ZdB2FYYVFI18Xymz3pqiO2C
cs67oPUM2kN+h2s0fY+HOyB7vWDuKLYzWRafnVYgr5T+2o12FGLMfEHqwngsT23V
1QnQmDU9swUM8MoEiM/JjG3Ez7esi7gJcpXVTq7h4KHLdfxojKNj6OuH6afXMH/3
c++rCmS9hvpEWHJ3Ynp8J3TINfH1p/5BacDxxODRj0jK1bzp1WEavcopNMg/SGwo
k/PMQWv7uiaadqhkbMLNC8zppLmrr6DvNDDOqCk42Kew5FMnHXK2qb4Be3JCQ7a2
B5KkOlFjAV61e9GG/M52pduST9rW8jZ/E9967U/64wxdB1hqXhkmcPfVuP73TTX8
LCvnaTrj8d1FGXv5VGsxHquR0Zss0saFFPOI7o7srNRGCCMaBk+CJwWqUnh/1gOX
sS9W9Dg8caFWNUKQr7PUKi4Lv6LukdknlTKS811AHEgYJeOHIVS2oK5xjBwFAS5D
zlgpACp7Y1CBHHnD4NwLZt2yXvulZONa8WUUM9RBtyp+rF++apB+RJ9O2P64MGS0
htUkC9dsqWEfEWWmHs6cm5lxjAlSt2+LBBOL/RbtmcsyhOZQ4o6UvGiIoEFf8IL/
SQaIxPkanJYJLjq3pl/kM9ldRp6K1het2e85e2h96hpXMt4QWNj3KskU7lGeA0YM
kLzXYUBbLlBreCskOGa2tti58oQMwHT6VcsHW2F8RbnrZDWQ3oWkFL9qDz/RSDYY
I7OUlsWFFj7mkUW69EzM4BvXYiTsZ6yBTcivD5tNuaJT74pRAfknkrO7q2IiIO2c
hFNmS1Paj/BZOgWWHgCLwBmxScD662ysLww+tLcwnfmxzZd0PUMW6tfwkrCOL2++
I02Qhk69WokWwcDh/qTXeK1we5BSU90j175OJtQf+kxxgBYTbzQgr5cRzNM6TwmT
onFQoTDrQXzmHXt6oo9TRBTAyd8JYHlntDt8HoOpQkZRrzIiZrp/20yTSPukQsmz
HmEMeIgq5fGgvLYCOpJxj5MmSkIWstf9vsLOpV7qqU8hh7RTlY05KKBDY9luvpj0
NV0n1XXEKFRnzS42EV6xZFUHeJxotSJcwgLo5kyrrvLlpZndko0l6vLTpr4a1nVI
8VmgxDqOO9zY58YaWia7eREFUGM/IFXrMvYEWcI53ZgDf1hqGwYGFLo42WU9swC0
3Cj7iO2K1peCNwQ88h7SBD+CB4tEtT8WRQxYN2XHX8TOOWLq714dKikJxVv5iNBr
Nfwbqtfn9JXz4GVMH56RXjgkd0/WQXhZWO/msXYd7sxWE3UrnWj9z7u0c0AleWAO
UWRxBg0QgYNriJkrDpyaA/SLaJznjy7K8MwnSrSWaAqGFdWXS+vXo/RWV+iPFOuf
26AeAWAjdi2ziEJOxQLcnMAweqjKSqKRbbHhIcrnX9hxdCJ0POyco/M9W/KjGnzx
cd3U/7EXXn4DyCWXbeq03jfMxvsxcw3zp4XsY5aqL1T49tmBcQOB4a0bXkfunkln
3Lw/RcGXpwv659hBX51GD31mlIq/Qyfvp9OAOJtT00+a/75+6snXdClw+duFLbzL
JCDRsXmvLA6rTm+1FRGnpq/xPvouHTUDJX23zlIB8l0ybqgHoK/f2ddZiyCwKF/X
S2AFKAzl6BaqaQ/O50KG+IHKnMxHxd65yr2GWNUG7Br249UgwsSFqk2mxAelOxLn
ZCh4CZYrl8i6ZKmYmVQA6hxBw6+dTKy3SyordurwdpddTq9AG6F74NVElGHMkqqQ
bfe/50IP3tJMo+JHOJyU+sW+Ved7RCyFbUYnCFlE8ZO/7LUKiEW1kLiQ9NQp9aFf
z0Kj2KYFB0tKpeaYeFsYlv97w4ReqVI+fUmtCsoerMmTCp/HLZT9ggE0hIerwN+Z
pX5XjlW+27u5jl3BkmjQ/91OJ6HTZfj91b8bJiSr8i6dXNZ29Tr+hX9Y5IGE0jhh
aqSDNtC4RMz05VbZ9tE+Y/FgtbVnU4QQiRshlB7F24aAIi/IF87QEXHXptoEfUEc
HgrtJk9AOnL9XpuI2vzBwP2gmBXY9y6XqW6FmZNXvJWigsq99nox9p/JpukucT5f
KKPb2VE0D3cOcrpky8UNJjqFWfUw/d/O3rD+0cq2bO3D6m34I628/BkkBdTQU4RY
QE+e/N6zVaT2GblfgoKkHYfqsXkl1FlP5z+p7A6D1x9J6w1fJrtBchZL6O6bsxI0
OsDA4h8CONQEPyg4S51XMiWbd61Z/fzUW1r83nOM/94ckTKE+COS0SS48YH0Rcen
bRakZKpicSUY//VQEMKr7bCRQuSHnZGuGKVb6epafuwxc+j0tBP9NU7fKljTbfRV
uB4o89XPC6kGHCKToZFRZjd0xE5SWXLWlW636UVndtSGp9NFXuXomYoNkVxrqleZ
rGss3WUm2/U0AEpW5280GJTOelfJyZLiW5kB+WMEbBtDpkZ2emRUW3dkq3EO4SN8
uzToyyPaKRk+VtQuXhSPk6dCR6YY4HhfOtuzDSY0TO8pLfVzfXMXQ1xRgh0MeEDl
NA8CCCjtJoA0L/EUCBPeN5W+pZnfZhW2ymig0VFOS0RKulrhWOMY+lUKG33yD7N3
nfo8EAki+gKJjI790QefAL8i63C76QfX1BIRd3KZlRgMHQeRjcF9bjopHKUxl2Pg
+11fzi8fLyIFPMxU9J/d8poV0ZM9lf5x1W/RYOa1Mb/5zgZqLDBm3A2bignNT5ZH
9aW7/PlTUOL2nmQWMQTbJiPf2amjgYNegcOGDYWMrf0LpzcNPsSvaMsfJPE9mPqR
PlFgADUsj1cLMe6IalF3RsgSJbL2hE3PsJEmrkEEhqY1HTX8OG0K2vdbZbdkffYx
IRCTen/2yNdRIkAzY3nZe52L4hpKdUA2UpSyKq4CCTTgu6N+XHH84EzSCf0XUsiY
y4IhMV9c/MqvyDoyjgYqkHDx+U7YQVIBqj1vVTU2AIFMm5He4Isk4o36kKOhC2sG
+Z6iCraon+Mq+4MxOpjMzxTLCvB2sqhrTpRKTHNDWMTe3UePIOv/SR/t6qClgj7i
mq90cwKyaTbWCDsNwtYbKfbIQ63EZBqmvSgMcj7QlS3Ppzjf9CJozYyhSExdqccB
k0IhWvH6TDJHhLVyBPS3Caj+jkEkGsxjxj1Lc85ELhFM+Z6LyZFK2gRuONMFwm/7
7vqkuUynXnYKspSQUgmBVpbProH7+9ofoyIkBx7iet1ggr5QA1uDxtu5Sy9vkTpo
mTIdjXGlt8fzIhL9VYfze5NJo37ST95H05vBZgpPD2MRmDMmMlhPs/SGyXo5dZBg
T4g2uWDjq2k48w5ET9zPN+peyzHKNTiczj+kr4h9PiIjs01lbzyEj7p1sXTRvIyA
DUN96yqRM42lTHBXBdQnGTAHhjP+/sfg6QAcLX0NRfGDYFxkDc0rKjqZBKlkS6+F
0hHCnJKp8OWJP3GIcHxe5/CpEDV6c1+NuEND+RrN2YUgDdw2e4sZjomGOm9bHQbq
iBeWH05W/NqvEsiI3gOCUAHWroWSKjOxHkwQhWk0CbOfhXEN3ifL4Za1a/EkThCH
WdIMXt5CdEsaZHVmECcdrqmzZ1gjnADnwpeHMMAiz5iDaO6cckAhDvyukIQaFh5m
42eV7eBZpwPR1nQahUMb2uU7JHCMjC1ERJP0NkcRl3HZrQujcqWC6OQJIEj0hBfd
z0FFo8qoJisF/nbAJQSxIbyAnZ+5gg7M84aMe7/tbzJBvDJlYjijctQ1rCLVPrgu
PNuP1JtvEUmP31Y3iQiNQ4M5nWZhRNRI7OQWuEsbh1vcVhFvuBYuJEY3f/m0u0FH
kFb8Ntk+965T/PdXYbQQxPmL030JCPP36/QmYa5xQxM5+hrAYelVwLF5btSFmAdl
YXXK1TxzrdOjtc/MKJvrdx8u96y/B2MrKpAO8FnaiwABN+DkrAp/C+X/wQApOnx7
cSa545o35gJEBq8ksSZ4m/ujIa7Ku8DkvbiOIUMWqjjSH3mM7Cjck8T5fI0QHA4C
nrzgpEnSqZyIKW5cEEFSZeMqJi+27qfJTqolrF+wJaU24fIHJilmes6/YUl/HksM
EGtgQv1MpO6ovdSJbQtnejwSkgb9ciRYyRqiyrJLxeFV7SlF/2eIxa97xFwBsD+L
rGO/yrTJlgB5tLsrIt8BLjUd8vMPRcTPgOx+gNCI56Jg2hrmbLzHg1TjwH80l+oM
7+Z15PDZaqsfckegwnLRhY5z67kGPeLoOyBvhFkoVLLrBo2D+rj2ANSRThxjZ+or
hx1AtC9mR89s4+EtL/+Vf8ZnmFzxzUXQxGkHgAPnl2XN4eTReJU9U0fCMOsWLBkG
f5c1GO3j4bmdt8JvojBnPDkcZop2kYZXNmmWfcyLLlWOYOg8AcAnrozgQCmxdgNy
06MeM3qAivvy+hfxkPsHdW1cNOYdKDvAL2Ga5TvPr8MeiENlHFFxyv8iaKNo5Y+w
CMSLWuQV1RAyCBl5gHCbO0uaCI+MrX96YnBOiNRkGyfsU4t90SdvluPMPDYof5sk
+qSqQoA3g+HSnwpg2ufDBQmMHfPRol+UbnnlCpkFkLGYsl+e2GtgOLFv5bb970HU
+CSHVpQRjbtlhq3ynkt14G1pq7wMHklwXOjlBWn8M6bD+M0bjYP4KxSGzVaUTl5Q
0CqfKkiR46zmm15vOe+W2n5q0pLgthx2Zz3gJ0Y1g9VYwlvcYMuKu4QUpROM+v2T
dZqfzYqqhXbuE0YLUowSvB4ywIpFaluVgDQZZKi//BjNf/9S41Qa7c6BuW3+Na5E
/w8HgYumWlbfvQUS5ZVZTU+JIpPDIGfYSOqe+Lsy6xOSKSQBkVZezupYumnQmbr7
H0XhYEjU+dZEUVKR63YyjazAtjvFp4CpZyYAlLI53l91hFZTua0j0AqeVl3XGUSs
m46wtxKzIgN65kkL2XsNfqv2m9lfSRi6vkYzzwjuF8ziWuhyBG2JdnimxEGjfj/N
7ziFyWw0Y2J7NYXek+JtutqGAZT3eTeytvebTC0bj87ch63V3Z2UNMxB031NORD1
XJzJQF/mNCDFN/oSN4Uw+50FejKgH2jxOvlTyrOPbOSI094uyQRb642/C3DAm/ha
zXqizvra1Te+wFeLqhAraitNMRFSSrwzPVFSVMBt1ICaX6x0vdkkdnj/WX81xZGz
cooxA7aiDyORVnxaha238WK8vm5++aooy8z57jcacc0ZA3aZx8n4RbVpklIAj06M
M/4tvlnN/pkvlTlWhsWMIMna9mlhhhp5+Z12CCXZ/DRtiXDSKu2YaYXEOzPyAqy+
0HK4RPR0H9tqbwezJ0ajFL2gGI6sIycIq8f6IVDcNTmqX/RBIsppSh7QamyIoQz0
0PXNe2pAtA4b65pbTTtjVSEq8QXVTxZv5ljvQMvlhsySdM51ZZmcb1Ab4psGSuqg
VJw7aLlUWz32FlFVeR0OUTLElnB5Wk7JUjXrJ0D9iNWkLGgQ2QqdPvaCF/ttVyBi
c9xnVfhMhPdDjeR54mNNm5hRI2auUa+cVbnq3jdhScgghoZDww67D7kpk6mTj0Uv
FwioMsLl8rQrr4o6DfmYCmhlvkBCpwhKMhAS/ms6/u6JB5RDs9XgyWuyCb8k3wJP
5KyNQ7XZVdyEhUEDGl07cNEG2ervl1Y4XUQctxQoPM5s/ubSE5YF9XjVHJuKScfh
zbcEvN2EJDrp2nGZlBYO+mAbd4kVg0jhY3Jsjh7VumW8BweCO1UApBP3d7PVGb6b
YqTRXXhAPEMWjl6Kk3Sr7gNlko1r9bOf8OvlpgTkPUUU+EyCrxY8afSO9tQQAyxc
EJb3Q8XuoiEATAvS5R3avcZpo41ATZneNVWCFjydPmfV05b/l3AcqDULtlqJ83c8
l7uI4Rxo44ZD6YdG9pEX336/LBL9D+wKDHAPSPx8xOhknhSfN6eCcyXNt6CKs5yM
SFWhr9x3aSys/TSEgAnp/3zTnRq6nK7CyDF2z9DJP0lzcoOJXD7B3N196BF2JtRG
GB2vesOS4ViiB75akleMsnuRuFQ0RRWWDWoitgnGa9ZPRn5VUnsiqQ7IJ0pVUF1N
cK+wq9rFiGEUtXblR0fQ57yHi6QUera7mafLcr/YAnNeEXj+nH1A9JcqE0qNzU0O
Q3s2gnH4GosEro+jQcsSQAGsLB1XWi2gGMQN6eoJgayjiCaxQ9N+iFzEcfSwcgJj
TRb3jyPJ+vR8+tPmEzM3dNeUjFr8YrZLsRhnxwIiiXw5xrY4OTzC5wPFXrO+dD/U
GdIwLsN5ezG42S1kQIruOuRpBpeU6ylz2/1Vevu/gN2JChNvlXt/NwayEaQiFXtW
pvB2Y8sKIfnvoV3sasSeIFrM/9rNEJ/lYYyB+bdxyytRVL69KtlQr8wPickIY1De
NkcN0WEWrQZidrgId4lmJ8Tqd5VJrTDx3FOQkTouGxfBkuuzSsOa0fZPTHHkRGBy
g/2ri5YyJoVKY8awZ+gkEwjl6aTUkRn2ZqZEmglhESdHlcCi4fID8+MddNERZogD
SZQnxz2GFY7LqxsStDY3cNFeLg9JUB5L+bZ53Pgp2MRRLDztyX8T3n2pK5NHwnk7
K7/qzIVRDMfKFUOKWJ5vxcjSqgBGcJXTkV8D4Y648tvC+NLCoHhBkUQRyQ2oSWih
worM8l7Wd3+DA+HibC6Bd3HSzOb/zE52WxKP8wp42kJpOROsvphLPeqgkDu0NUUF
J4MOXkfuUjKMON05oxNj5FV147mYCJuGSB/WsRRcI4he5o36kB9WUU4Ur9IveM6a
DhsB/c6sj+h7irOz5IWRwoGeCQwJMSNJlwsV3e8FFiBxNAScbXrsZ7wARiyYQBgW
jGpVPOxn2UR/2S02E9/wiQJc9HajFQcAlYd5QOzFE0eIg4SxLnAmTRUmBmEzENyS
fBpBJpxXOCvCco5zfw0lTh0RVMYFQ+mLo2+SG+Q02AvEY0NMlQLPt1R8tmuSC7U8
V65SBqud1fJ41lDzHUxg/Js8LjSAbOFZskNP92paVNDQJKVWKet592VnRm3D8Ilt
axh+Z54MpWka5OyXioLCMthzoVNJxUGMWHqXEPR6c3g89j4oKBjESo9PT5OMaJ2e
0C+JQvHkzgHa6qhTIriIHcFFdCa1Vm81wdYdJDzonFPcfXz20oRnLmPBcOn2eoo8
jLxJUlQViCY/AAelViwO1p2x6j9uhFDUNVeS+V3pkwXTffueSsopApNAOxMx9vQY
VKxwSqFtLj9QeTGWBl2DFGD2iiuuZ++0nC64iauwtXDWhLgw6tAIaEeBKFDo5hc6
/fpyFEUXTPJ1O8WjhkiWHrSP1djSwyzl26Z9386kzCntTbZiscZkH2Wjde3fnzu4
aysdTEqH9JKYjud445vrFHmhYsJhM6pazLsgtinNNhvqzNPEnrfJivxiC5MiPjrj
QhNDpzIct17daROQNeBjdKJ6FPcxk5XIYEEbqpGqcpGfVSTVrJWzmSdX+tzvel29
f3PN122vH0Q0qVpdU8EX1LV7i8+qHgwSKIc5Rr+YUz5WpiCs4ZaHpJOfvWh7wObZ
bmybXwdoQ7CtXZbKsFx7CwXFYZeI1y4OMTCzvkVXAmnaQ2Z9jPAC43fMYzRo8O/l
jWryIKEy+oThVksFwoL8QL0kvYcl8UnUrb1nUJA28yl4PN/aNPQdiV8Ho5NIuG6r
iWFpUloecsrSAQbN20hTg/iQc9K2uFttHz7zWd3LkjObV7OZ2QjixDqDpEG0iptb
8DxZtAEuoa5LlUhHI3dwRnYVCYchyodF0TT5E5dq4/BIyu3ssnxQGieUbbJ3zupb
Q4k4+PKZOpt+RY0CNqzjAhndbP8DNnGaNp/+Fn0F7T785ObxoolQdwvK9Qrq/XLY
Me9oC9/YvBCm5H/MUY4rt0N8rM8ef+yMPxL6+SkZyAMg2/mKtLfjxIp5sBxTlKue
4n2Zav+2tTxWqox6UrngYZv7aKr6OTfXBKabmY5hoDQF4GqkylbW6O+coeXicEtl
2cd7iULkr62NDNRqZExUrFrWGQry81kBy575lgYpNlOuzGw2hauqmP/URMfXGGfZ
f4uLQ3wlE+ug5w7q4xGlgpurSUcy8E0jbcpaG+ERHE6kPvDbwloZb+r9DjZgb6vS
SDunVcMIx7RUuYUT2VFHnBDTkZctKaKAM6ZIMm6vv9rZfEfZcYfgAl5jC0QknV0o
LJXKG02N/7nwdihI39JCSuuT0a7mMuk40+PsvHxxMVyK9LqJDKMXP0jbJiLa7i5d
E9hbDo6FHKUoHI+7UjVxPhI6BbAhnd7AZQ39f06olWRfVj+W9EW6VfLYv01kCldk
Qkbby7Zx00m6YVnihFhB1AuaKwZg+f+AB5ZqSUv6yN5m67nq+sTcxnDenZia64Ke
LawW2SubilA50kI5QnvV1rXL2Dk7InmzrGOVm95Uf2E0CJ/9S/sUziapPPy5Ty5g
7umhS/GwqOimTtnodudV8iWtaVOPhF81RiFkK+MGdKJv5XbBhibM/qxyoNrPLhUf
xZz7rCKXze0gUlsQ7MjqUBBxSO2PFb273xRuyQQN+xqOzs6kC1zZd/sbrYgmCQZ8
4/htaDOALRuW4za4cup3GR3J2oTfznJiYnwOnyDcycDIGMa5d5Tn3t6NdDqg3dWx
5V4FKChOgia1lN2pXwLA7BWGdTuslmoV8KC8+IW5Y2plwkgBmS1gflBrQmM/Go2G
5XXZ8pD6FiGfefLf1ymH3cSBjmpBu/L84/mknOXxR1f4EvITx6nRkyjdcEA0n4Ob
++XQG/DicrnGgkKQ0p8GcdVafOs6b61XatfHbycckOk/3ssB4RlD90QSJwwpG1uo
VHOLO3ce/3XEsR1FWFpXieGGdjS5OU0QDfXFLw8SiGchESKmMA7GsFI4+kHCSiCf
GggUTMtgzhE3sBdWibaPe95HnhyGBtgsfjT4yCJvSNOj1FqEMp3VZEtMBCSw0anq
ELL+mzclu9cPqJRRxwbM6kEBIbVHQH7qtIKCzbhg19nIfnmB3MiC9d4Xa4qh7fYF
3rMIWGAKD+BMn/T5qMBvOyvNgopaJ9lAlF3Lgpc8kdFTVHRIBb3dHwwLERmNU2HP
MdG+tx5UuTHZ5Dgyx4dLkn7J2ARS2JSXE6WAy5yswhifOQTDN4be1QBqNiKJ+S83
V3CRgfdZezenxbQQzg6aehxO0LYDwP19WajvphQEp+bQVKx0pVDp4hpwj8fjIy2p
CeeBtwoduCNVLdzCITGeYIPq6+xrWyp9Q/HUFLI0V637BdvGRSeiE7eKAQU3oafs
548x5mDJZNLrbuosM6m7XfFG88U/o4D3kytBu0VewQ73LpHNhW4HVeMipmMGe4Bc
Im/ilhlYqS9Vm6uhC8SqPb5BiB8wInXLRYpDr9k48jITRsFW1JjnUsI52qeYu7OR
jpsIYr4aNUUV7hbOSPZwn3h3oYadKoHr9QXMSqiFlapOe0CVgDd3EDjE/vbBp+RP
RRzbHfS5v7GgiNRAPBbrOgtse6irEyJ/tTg16yeAuYjTllhjn+mAgXGZ6Hsd5XCg
KB/reWsFYdMXgYrDF7wh68nVz5PwbTEunDSEWVDW6OUOy3UluVbAv6pZ7KXFabjU
KjXXtRiDUse4pEJ8Zyyx6AZu39G2UHEEXwhP2aKb9SB4XzHpE8PgfI3NP1luSgln
j/Hl/zhwpcO3an95ev3DUdRzEG7E4/iZvQWVnYZqPsi9LwTUZXwQ9DM8JXYs7dN+
iqEgEB8gp7LV57F1vySxva2n22TEGppU4uUOJOf84h8dBJfsp37pCu0fyZqOgqh0
QzvGuYjPw038o8AL6l4qzMvuUGTaunRI3cH6WZKLdqTw/qPvj4Ry8G2WMdyrSa1H
odgg6n0yJ2SroDUMqnuEEsJKtTSD9fE5qsmaOyNcA5dlI4RNw+MNvM+wpUVxt0TN
tSYTxzBy2ZI2sg1viOTgoq18uvpP4SjcBoPQJ75xD+MBH8T56jq79VDOS0ho93FS
XZrnvNvvOehPmpqivFGdWi5OfP2d9fTyvy36Cw+8GxhXy1QDEs0JAjom8+LZy8dz
DfbsS/73zxYdC2axx5L2t3K738acUoGI6k8I6J9j+MsthMpCVF6UaaxtCKlFnIWC
7B6eOv3rjYXfCJv7tcjOSko9ncRI9KeJs+KlQVTXMZtmjkEbOWw4CA0ypugkce27
KOIktVXRWTpapUkVZnB0gAIzJmNaZPfLSRJ6IReONVOdXMOTzwkU3zB9OOZOYhuk
SjsXvsOZ0SVcvdqWA6iyjpuVOhCOWQfeU5Vuh63q2oD4B35ZEclA9UcojpPKihZW
VxZU1fFduchJtUHzSQAd5H2JuplT43Mgj/kQwRbO1VpiZU5FqXuxwqDABDBr1nAn
gBHibPLXFeMhDkuM7rr7rn9D7tjj57OCCz1xyhGZyCpM3SrJ6B+Ime+6O/NhUpc3
RP14Y91GZuYd6VbDmU9ZalfOF0ryEsvYMhO0aXl0Kop6uxLqcGIvmEv5JvNmguHg
RBsiBUaaKsN88sRNJYw8xuTaG8Xh/TaW/X42t+M819iGA6mE7sDEUcZfq7S++YwH
qhF5VPnMvRQIGMtaCZsA53hBNsUH2PTKUJY3AROJxHr6Qe33YsNAramzIWUeZG/n
TxXmIQI3NCOzOrNGHjI9Rq6rqVbYlfBxqO8Lu5gMl7MC3JRNDVz4PzhoLol4XKrq
bP5FHD3JG8UOnQ+iGB4Zx2LiYk4cMixTiUfOff5/PPZy7WSbkQ9JyF+LPE/jlhAX
y1ywfWZfS0TbblrPDDxhQeLBsERQ89TVC4D8y+CDnKui/PQbLiJ7qr807j04M28V
KL/7gAvynHqrNKb6y34qb0D3rwtsITX2X2IV9mtVgqb/qIVenmzOqJQDsO0snzTp
GtLSuD+1FtEu/3IBPBMazkaGH4a35jlqH2yenD0EaYx9gI8kmduGllylGlbqlcPz
VsOPQgp+IQONEk5L16lxJJdsxE61i3TxPAs2zfauTEdHuH/nN+E70imnomm6vxBT
6W2wSEjIj6CFMLGe7KEhsJdrimvigv50VKLDDwFveJpBR7AQ3Hw+oIIkor5D9yy3
x7thBnt5I8mW3X6ay47JIvvTZiZnFcRAJYYTEgV1a14PLcf5a9564avjt6sNjBFQ
fJMwvGKNAE6sUtIOGA6eqLUQ+2fMcTkMUY3GX4HPqEt4fpfvRzjRcVTFxGNH+KYd
bWXhelviimhXKIB5Pm/wZN6hvPRMUDv6LLIBbNXYEKco/ukBCIigKZQPY8emKX5y
vyqlhbZ2InuRsM7mMGebKZa8UPJk1qit3dQ1zqKpp/iZCburvdJ3aT/05rHUdVU1
V7oveTMyV5Cfi/KF1Ccdjj8/+Z1+CXk7uVe8weayGE3VuhiYnDF2Wvd9rCPkxxIT
s0gcRi7rYNkuJUJdbLee9BT0jiz++HrHwEUysbkLJKkRslHjtOpBFk4oqxVHaBpL
TSdhyNGPiFiCvFf3AUF1CKwX90Yl8Qwg0Zu/fIKJadRhJ+tb6Y2dNg/nX1qUWlHR
42djEtGxQqJG5C6/yZvnAUkU4xu3wZWZJ9i0VDZSHlgCSH+FXo/kOVjApw9Y+Czf
0VnQAko6gBRGrYqTp4CrTg+cNUnl4jQHLueuRMIRMMUfF1KfWG9k21bQiXBOqKnh
HNI3gqiRrI187Y6NDVXeTCibvgP1tPdB8bgNDn9mDOYNVO0IiDr2P+XsuFdfiwRA
vkmN55U62IX/nGZKbTt4cU/eB6Ug3Xg6hHALIHR9GMktxHOJH+ZPmaLPg/i7h3CN
Cs14K8Vjo/NhuENSi55dnjG4ee4pw+Dj2E1jmzXo/uo/e/mov1EpaVMVjZZ1TJum
HQuYdXg1jlmjxiM02+nGJVd4U0eGlK7JOFRGcwGc2nbMz6unX6tltctBpFVpgR/X
vFWOjteg12moH6krImtoNiWBzrkg3QJ3Op/FZ5jpD2ME/o/9S0oTpu3WpDfJnaOr
I1v6FRs4KHZSE0AkudnHHV6PE2e4KdexDhSbFkEaBeRf2aebSjlXVWOEqLXOUl+P
JbLMoC81bNECO93UBZJeeFOsyKYvy3rbxP2kTeUQkxGDxmCHnHwXKrTuVrfJsKD7
PBe48vSHH4TE9Qrl412ooL6mp0ULwMO8aDn8180ZNeEcCyQ1bPF07eIl7nSi5TnS
fszNZ17tQBqtiQOExtzc6fl9u34wAQG+wtCdWjE/3i2usCF4TQF8b/goZItl/ne7
r2tA3qh9ytwA2e7SU73ZfIMStEHZWCBHNTgI5LoZZsLnHq2GTsTvv4F6ChKZeAGV
t9Tww/psR1FPitHRdRr7FtSFZpD1gkVVEXpj/cNNFYveGpAtwgUpNuiW+0mhPJEi
2C8dG30iqBLEdLiB5KBCSuntJ23qDJsybayUR544JTUoA3/qgPPDcwU4iO8/EPzR
a8hojTwEIN2V+cp4by5CDFR3M4pr9neTjsbucs6ozbBysPFjreQsVhJctKbyCD4t
U8552/ThopM7LQhFmgUd7lJ+iAqjYlCsSpihk/Diq/ul7pakktae0EuuSIhhU6CS
NxQREC//05CWrxvTgTZ1BRJtFjfk8M/vbA9YLS362IITg4vhvBLagWRM0QWuxr5p
y7sZC3JiBvckreMZCyn3vZ+MG2zZ4Zn/7kNPaUJx3VmuRsZd0iwLDUYwPpvjQjyD
dDeCuNqDt9vW7kdaznUQmQ0P5AgpWByoI7TogGp/WvPvKpEJuFwzIMPU2R+ur5ox
eBDw55v5PdALEdinXnzcm5MaMXZ9DqoA6bnhYbBDDb+e/Giu5RTg/yrB5pGr/cVx
qxyXILON5KzbIG7Feio0oGmB/T+kQB5Ohd2rc4NYn3HfUyI4cgZwijdjJdVtwKBT
VLkOQ5qJQBeM0mW2noOqrYXcwUl7js8XlfG8IFmicta16V+WJ4ifEtzV22qEel94
pnfFqtrHEQPffLzZT6bUb/DGxOdnMhPKYmKun4mEN1vWisFA/Y/B6o2U1rZp7qoV
kuCRy//a0Ye9rZsn1qCCowrioDX88P/ERuIjDe5TIgg6+QLwzTa0hmjxYQPHE2c2
7BUJxfJdNeRstEeftUlO1M6EMl8uy2hfqUA9/5g5sE0yc+MfY+IMhTz0okVlPXMe
I+A/XZZaJ4z78cpqcJ6SxJM22yA3ulMAVmzWkSTi+WGF9WvRg0dMI9xgScaTPeFs
ZWMEDVCAFW9jSezB1As75dXCMZNRSv/UIHNWxdv0qJCkrSy0ngHSFqKVCc+OLP3r
lknj+ZsHTfrps/HX78kX0tO9yVeFAI/MEZoPAGzTlmacmgdIkZBDX+0ujbdfa65h
QKRGKBpZjwbEEr9t3hs8EQw4EPiLT3AvzXdLpjIoGPRAMMlou3jSlGaJByn4eP9W
fg2/00kgT2xgq1diqZp0UMacpCCjonTWtL3CYWCeakcf6p8S9Mctj2DhjBztbIzm
pAsMbQrNHryeiMSJYl4GNdzxJyC0FlogLEeykWfsRulPNp6MGiTDGBMqI2Ic5DGs
A6kqURdSSEX7R8nx34JHxeGkWLhYREHCw6xl6NQJVQ5JppmHgk/cuF9s14PFWO4Q
0O4AzzazZlSZt33s6NktTXT5qVXNR3i5fLOs6ynxZHQxO9KCh8P6ZZ/U+N5tgzfW
bc5TC/u1mtkAXkynfe0QI4acu8zNZChvL+X7QDV3AyYBEQhec4toez3ENQhSElQB
4VxKo2PVNqXiF2yv2D/trd34gdAPr83/HAT18SxvW+ZaVA8YP2mN6S64YHiwnlKl
JL5DoYq0Wx0f0v4R/gnS2e/6vcwwZQ/wm2IxVFjIUk5QfEH3zkNxibv6u8qVYqm1
U5tsd2dkH3TrG1eE8i0tpnwBejQU/0T/CdS+iHuSc6ezjphIteZ/wjLgs31919vu
8LUPI8jbpW42to3pBIL0Ete6hn5uJE1cBTicSlsz1pE8BKVtzqmXsV/uxqCz4dTB
GrYBlPiioZxZ1nEYrSiWDeWDdXYCndfmLxFxzVbIHvS5SMnD5/oqwdjaADPM6j+r
OzpoPC4ssQPU2LtroW8y5FfygwqB3sFKJf4iPuvCKOtYENx7Ui5l2zZL9XuZqioT
mLus6Wg+KCKRkCC6LxrN7koeim29AZzGz7v5vj31IX9eDYPi5bRf/2DBdc5XG4Ym
WcNoFxMV/2QTW85aN2wG7LAi0ikS5CvQCdo87lsTgFco1zjRYD8OIJvXQDAS8tsL
+2meVrDoBX0tACbAJMR5bxg+awgJwIAH1n9o+d5XtIFHA5x0ZqRA+pN218mRgYHE
WKnH1o5nz4vyW2kbFEUX3xVJ/2kwEB4ZLx6twQbtE7ntL5l/FnpCsgFTPDyOSRbt
Zdf7i03oPdmEmyucjI7v+C5qsnH7gEC6cT9O2QfhLEYJN5MPmCAlGac/4BZyq8m8
3t+WQ0jeV8n7CDKRo4JGMKYN+Zv3o6kkE66NCe8BB+7bLHv9iOg4RK2KeXJL1Q/v
shuEVaMWiLUKasDOfebjrc7Z9zV+WKaih6OjtWEDWNfClJUeRcYdepPZ8nyW6zAy
73TNS/sefst4+7WeQAnoC8OkYF0qGaa4fvkBXW+HNLYxnBvBPitGYKl8+bGs5fqz
u/sN2IxEv4xX+1/I7kJ7Hsvm3pTJi8cV58kJg5KeXxCIJXU5lGbyBlkONz9/wRNo
kyZwBdoESLQW/8q0bM4pI+mAqqeEKwii4/BaC27XYWE78Ecb+VPwNt4Q4PvmMhfY
wUaf/VST9yZk6Gn0Btr0s2DNDYn3X7shZE+PQVkLwZxmS5mgpBREIjWc9iPEmFoS
qbY1AdZYptewKOBupTfRskbGcJl1zTEY7bMbp1PGs6Jh4Z+CpC8zqteHrmuTzda5
Y3lJVvK7J164CS5yyyKZEHdondOmjUp5HsCQtTAor+d846JfyNIwckJtwYu18wEX
yrA9c2VH79oXohGJJl/6XC4Fnv03ZTuux3vrthXZvBAThDuvUX4tAOBONxkpZYBB
ZoILAK96YzVfWW4pRYpSz2ivmwMeHMmZ8IyhHqbWSvhT4oLgKJ83KQYT7t8fpP87
oUdpgsG+58T9YZhUzQGg0u3bWkpFwh2KohQkxFyJHEOjwzEd1SkKbN/MWBcS+l+M
yFf7TDf+/Ov6/Vt2HMrY/d2GnOy/jTqM2w2nBaEjeD/TYIjNmwpZk4IvHweagzqW
EbpQXzGX2HKB44IhAJMAFxIirmlVn7XQBpnRVsKOy16P6H7PXUbRAl9b8cbs1XDE
4ct1+E8Yf6A83SwNqvVo/q4fJi37YyynCw4JB0z/5SEgH+OA2RgjDbwWn9GqR7Tz
tNH+0aXoRnmb3pLm9DXOkAFUVwOrFf170okG/lA3N7esCvxCgK2DBZ2oj+8xTjwI
ynegLhU+CB1w9F7thw+L9KTdZutviOYcl1lsciiIMSWyu2NOGRQ5hU0yVfgeHQu7
+cAFjypb2UjxUYc2gTCDj5eYoVnnr8kUmFXk205nYn0AZIOlC6KqWijwKjBCb5nJ
0T81pUgcUu3tF2QrQhQqJcXqjA7g2XhhxbwnRXVS+/modje+loYSLLoWE5fTYClC
ZwFdn7j6Kbo2yUaJQjF5ThkiCUPmGs2YogaGiFhWHYXi4dZ5KCt1swVu69vgOXDO
THlnArMoOPnyJJZSGVErKNxeq+i3C3iwLznnYqFQophRIjyePowY7T/YRz4iQsca
wX2+loEXA39c3DTp9CIS7T2QKjRevCk/licfRIx0ljOzW7CzhbhGKDbOkooDmen9
1YehJvm3Zgs8Vpvw/7pia1XGnSzmqThjMKxu5UjmO79pRGWuE+w/t3oGzndjq5Td
hkoeresTkCjogxAxdW0tJle9yT1Xt1UjhiE1BmmtKCTrLQfk7ROf2PnQ2OF7MDbP
rusIcTQ2WCNMFTbOkkVlmuzZybe9ZD7Yb0is91gOCTI6WedJLfmeuoPajvp5B93H
KJvUZw2YUDJYwBVM4wUCexVMYgaDe9QOKJebx2WAHjqyLFtlyOTqREdAjttTvSZ9
7ZaYm7maRn3Uimi0gz5eaAv0HBdBUu03GtM4r+A6MRKBW8RGSQSs9Z1GUYAof2rh
PXeBc1bxXKekQBXTeAvu2p/VHNXb0FtnIDPX8SSf0qNs+syMgb8AtCb+Xgcsf7Bk
KLlhjRIqVu8GN/gbomJJBJgNNvnth/j5QZOBeZaDIF4AICqsGkO97hzL6XRoQNrN
8kUipAWPq/HSuXJ5d7pemNXwE/lJDXoDnjYCaJU2YtWmZ6jKBKUoYy5PDoU9SDyE
8hOIqgs7EoG7UFnJCfZUUYCsUqhuUovnracSprYw5XIyGd/H8KK0H+CFwRojIwbA
/Vtg3Y7FB8D75xLoHt7pmvgbFCwMKsdXNurmPdjaPhiWxpmKGzCSSEouq6BS6PiR
xqRY/X5YmkIhyj+ODP9BqKFi2QBhrOoJtqdvFHvaWuH3g8iRINzq6+DOIEwMnV4q
CZuald9XLnnWhyepfwMV8rIGH2D9B5zbxMGd8zqZ6mE/oLOHk4mWuP3TSoZ0vIvr
a+yVgJkLCRW1iD2ew+0TJO37SzNt/2QK6XiSGfRhcy7uneDm1koyy260gBwG6PTZ
Ebvxymk6Fy86rllOQh8DSbiT4N1BdvPN16i5imsws+OpOAoKeR0XN6NObxn4XNbL
yHePZ+rRiUaNs93P7s8CgIH0ETFgzrB7kBXICedm/NQ+MJw05CHKw0FQ6RAH/c69
yN9iR/ELDpmyIF7pv6++UfMtBhtGTTwLYCQHNZADAWrdw83EI2N9cfccKBWqbjNQ
YJ1jVjDxD2tteVD1x4BioDOEpt/XzTETSxwxAWx1DBigBprUkQC52aBAVzB8S6uI
ChUj5GUhKG8tQByjifPCqyfNmeTCRptSZppLE/6z3QWIKqKgontLInmiMCCgbMHj
9j7BzUQwQPcezcQOI9QBokMmgC+Zzi1vj/QzHPOwQVHlXflZEFKIAQyKDXtmeWDA
zN/aVFdNtqasxlbs8XIlwgiPc99PQS90eMMiyhjoJDXd5syrx4GWRajARsFn11Ov
eNMkkfnFJVBWVYbGlQ1FTg1tTVsoFcrGFwzDBxm36726at2wJzP0OqSeNtyHpjkM
jHSf4Dm0ZQ5iWg2pvU8omq5f4xEYHm7fg5QHB6lUm60=
`protect END_PROTECTED
