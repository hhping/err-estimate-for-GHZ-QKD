`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXcsD9Yugy1ekgnXMm8JaJG4/28ELjSY5R0jQ0GBl7EZKrkwNwqlGujLzKnqrogO
gWfDb80+J6vKrqCR6I6w3QaVc/JqWwbruKlASZfwfCevNzfmbnA8UVGxJyJVKLts
4DXpkfqe8AhnJpECQtxIDE06dZJTgq6FH0qsdojiAFcP9ygJqFaqbqTBqFMEAGHh
wD01L7SlJKYoodVUCsN1aPwqgZT95KODT6KvL1Y4VnQMlEHQHk6mk/V6BdjeA4si
s8NBi6t7/uSe8SmrP56olDQwPnHjnSe/eMRjAFJqL9iLJ2pVdF84noPq6U0iaG1+
lH7WwcRapUgmA38J1TNH2BEvX+hlT7fn2oIBFYj0b5XBjIBVmIQB/Z+DDBwthmrL
AOOl1SU7Qoe649GSqX5j7Pe02YKKbHv1EjEfdDNK37LREoxSb+mtrNCC+TigfZsT
T94S2ZmJvsF49lYtyeHcGCNn3rQpcAW7zepDY2qx/1IGM1os+mLNoe+/EZK2DhL7
dpIK4kGBlFHAdOPvqr20DjHOn4+3LP7jqe4KL2fcMf0v+ecW1w/JfiGkcIkAU15O
hxGgNJ9oDW27gag0k0lUntUiuK31nOuH2BnojH+/s6tmdAOg/WHKgXtFbDQCH/aj
rhLQhd2+LHpv+0WFfdB6nLL7Ehzper1oJhyTjXvW9vpSm1PfDifSrXB5z5BoUI9W
086eJxbbxCt0rqN6EITlDnRsCXvNlFrOGqdf+c6ZBXg=
`protect END_PROTECTED
