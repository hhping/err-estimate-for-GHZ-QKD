`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6eE7xaf5ENZuG3lSyW5g2OG862FtIMjxzqa9iZ8K9pXweRRyxDS+R8/IWIbnRH7
Fsydaaapql90aOjUMpBg6/hjqgOOgljnHw7miFnU/q5wqJycyRYARQe8LHPQrlKY
Z25yCoci+4OeVND638Fh6lH+LIXCtyibYgE93YzwXz+h/MPNJRUz4xHmXj1oKusY
X7ebQW5/zflUHluDJ5MzESdb9eupThs5q8UnMpmipCNvwmqf5KxpQBA7VkM0fAM2
2pQiV8UqlZNtIPgfuoCN6B7YW+/EOTmlDEj1kzFtPORdpIc9AOS8LHYm/NQjIYWD
fW0/bpT77fSV/uo3WPY8zXHWlBvzhw1sncMQpwZzeFS1lkdN2e45S3GoCk4okVR9
0FIceQ8jKwtpY1jxU9OjywehRQQaum3Ij0m3wU0VnsnNEVYbRPA1Uhbjm05VJEG+
ZFgH4jrJd5JxQomY437xWvHC/FZt4PjUw9l6t5pL49F6WbPMbQKhmkJx51PqEjpJ
ZMP5e3Ek7Tq++QWGHj43ERXHOS7CpHuyaE9pek6lkMRbpTLK9E+8snTxNzcn6v5r
1FkovksBA7jWG2Dikgj3+6cd8CByBCC0jEX0Tv8T7pNQ1EWXW15F/fUwT41n8Nc+
MzFk6fOg3727Anr+6VCA3YBrtoZUGpahtarxUDJG5jdXNmwvWPwbH8RdkuH6XDGZ
xsVfdM2vPEtmzO/dux5Noc9mJvrSOlPdRYzEkZivLICo6TQzoJO1DnhJhTZGkHkH
su5Rfer4ARGGU7E8UXSxoaeQ0cmpd9BDNepwj2U2ancJX0DkOExFe81a+gUqvBaD
uVe2htkwWf5cnDMQdk/sVrv0k6WypQKLUY4xKFUbqc2sQKO6jakzQpkQc/1QVtrL
jjzDmEjnSs/WpmTEYWOn8wo1s0SOVyMFSdvWysehyx7Sjw6fj83giGceC813hdHN
RkE+36aNrNfyaQ4V5ywC6ZIQknc84wUNYvQRXOOCR7AmhDkIu8gQbFLDtwBnIMEG
DuMm6Wg5VpdDfPJ42G12cufofIbzq7k6EVM1CT0RWsk=
`protect END_PROTECTED
