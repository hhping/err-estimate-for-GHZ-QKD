`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4fdFwsJpz1kOkORbJtcntsaZsszi1t0aXciJfYZ6kZOiTcjig/YUHphhyN2myXb
S0JNBiNxJrcV1j8kVvjWtAsu08n26OTA6k7TtSyLh6CNtt7QrRB55QExAcz8sQIX
VegrOOjpt6GRZHkJX+JEtQLvDOdO1YvBvUfQhiDf+1SejnwVFmqyY7dUZVFKGmPR
L8+0c5CoUSU05uZmf1CVs6bdbGHU63i9K1dDnmnkcAM2b7Zx51DfedWUpWCsst2f
BOF6F08o3OnqKjWTQv7MGlW0KZXU4s8zJI8mXR//ut1AkAN6kfV95+PKE/hzCbxl
e2UUC2pH3Wm3mGo6dH81Y1gglTiKcvt0P+eJNX0NDeksl/SnYb0DyyMiTIFPjNPd
VWhGMKYsCV9nT9t3ISqPRjlSoqdlFSdkRfkXw5+q4t3KGq7lO176BA6AF50F9Ek+
AwFqMuY+1BnkWOm6Fx1pg85K3h5yzkvAo1YCMg53I/9K8tgjOa/2uG67IVq5H+54
74qsNRl9oz/Pr20n7K/Wbq/9rYblhLZjEi27bShRekq8fddt7sGJchBfGNiDtvuH
pbgWF5W0dPTnIC3frTFAE72NxggipBnweysR6qA+2Y62yhyntb8kjwebQysr1h/b
/hACGRFZElRSzTv0i5vuGHc5sfoTeceU2gv403RCUuq9ZcPNWrsBBI0MNOiVrFmX
0jgjxw2bpnuodW4dJl8ILl+zIUNkd2GRwV/g0t3SGxGet6IKC8+tCHQCXDihDl+Y
Gmjp1p8PI16hxf90lINsYO6jnuUAtko5AIpr8hHna/NOFwgN8vGj2F9lDj5I1Zkv
OR1t4rX542scd0DMmQTgJlD3wPrXaEpVYnqOpX8bM+ncy9WeY6EbAWXQFmZr04EP
aVEYWmjx+IOFVReZDmTz3RBE5DPXUQhKm8Uz9Jpdx7cgIDYibpnd9nl5BCTRLJTG
tnLq0tP3ia8sNp/npF0UNNm2woMv3G/S9dG9LaWx69Cp2GSum+xU9DwAwWPemfPc
c843qMPrduWTklf9H3faejEwEF4Yo9A8KyPs4zPwWUnKOPdx9WZseA145Oqqn85t
RuhtM+mqNf0GkGKxiq8hKQ==
`protect END_PROTECTED
