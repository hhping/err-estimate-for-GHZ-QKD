`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxuMnpUjDvgOVqKh1xzVt8ybGmw7KND+f9yr20Ttbz3udO0BKghDJ0XeSzv8zCVH
OGfhw+iZdpRCPYpdQiB8eTKO+Lg9I8kiEYLuF/Oiq1KQdHY5tUxYbcbK2ldB6KJd
fm4nTOBKNpCekB+4MFxaVwZ/T6RhbgksdfzRnT7DNGwXYC4FbrOWD3u+6cAFN+qv
CajO0e+NiVYRfcN2aUehc/5/ih5vwUucF+qmEWSBGXABIBqbQRCI/EjGvgS9PaKf
6yPKHuJnj/4GXJHBBUcKeridHVh4XBw/y85VbDf8k9aNhM/xk3Rznjd/wJUHb86b
ptJi/3Pb6liANhYbxqHllGeDwV4XN+Z+MG+/kmCdEJVTXBZsct8b2fNJGecoEekk
k1C9hflZ1qlvUM6/H+kd0wahp7WWO3YvDER6JdkfBKmSuY4IhT44XSdDJKBy8Hz3
B0IffnPA4ZSFK4+PtxH3zgSLqRxA3bU1COhKg2uZKOxrP8KU4uDjqeYmqUz47jyQ
GEjYYhL0XHU8c5ooMDs1tFjWffon2fRurBiXIvWFf8X0U8c1bgucP3O6F2wa3Zme
UOFVK8WE3r/0zYUOloS5HrGJZm/c7TwLZQ8NDmAOZzLuTaq8n67+g2oKs2vvDTP+
AcB4Vl/wLQUpKkDwK32U1UzqL1ns/eRcPIO3EgNmE8u4rOWkbyDUWRLWxePz4Ud/
z8wrBBBbBS+Hg6WAxzbs0HR5/Py3vcIJDCmQNVo89FkRQ0hGCvvmsrsNi/J5YkRw
izoUKnDD+/j8iqNifuqM7nYU86SJM1KhVQX4Ase/7miZvOn/bjfbgo93fh+yAOAB
J9OgTLbhjG4KXgJ6JAp7roo5kEt5ErTM33mZFPTpwAoKWsTR7jMcp8WI8S1kKjjd
VueU15iiAHwuiI9p8Cn2hsoguTZ9XgcR+rv1aHvJIBP+3jHw0KNdc7kAMfd/T+4r
YPyjAu29k5sM1InyTSF6tZrgIhHPodIVcrHkt/DCNA8GzMcJu2AwcosaEfA9zerj
eyEF+LT2e22Y2PekIrgLqmIYlPs4FFzr8xYM7EUQ1Gh4H9yIvTu7l3E8okMph2tP
yj3hlqd+Fwh+YVisamSn0OU3NlwoZYsYzdHPZvE2zZzUfKWH0o4gcHIODZ7O6XMw
m3SLXVjkjIZ1yuV5l2mU9vORQPHeNJ+Ipi3lTAhTPNsD7Aawhga0EqKY3O292D9Q
CEG72+JI5rb41B9z0s3tQTUxnZAhwGSiktLv7OJaDWIq1Wx+8jtkyg+cNtzew2Gi
wXDnND/MvCMOhRMYBn1tc1Mcuk/xb1LjjA2BIqRF0cbFBCBdg0CbCjhKPezs3t8O
dGKGkqGiPsZCZKDuZD7HL4IaAphB+BGD6M4ht2KHPtjFpL6T+q004xITofRqkLBd
YSxu3vxp5JX0x283qTSOzqLSA0yoSbvwSsfU2W+TzBkStT+ALJQptYGbQ/c3+bFg
E2EMDKvyv/3ZxBeFkQ9/UDAdcIrTmMuwjb2zjIZF67UUbehws6FRHktJMeBDEqFh
PnRUpvhWmYeIvULGfcjF2/yWBSQsEB36VfFO+u7vA+M48wEH49wKcSp2TK6ufKCE
e1urk6AcdGd+FPYokgTn5sTz+6Ls/XzTNeZfFScdhTnQqxiKWsPkKOO2qF/wQ2j2
ohBIpsRwvsHot/Pkodlvdd77+ZdPKPDWSH6ylBZw3gRAHvxxxYWPNrsFHN3PntFe
QARmQBjWpLSYNoWwV0RfyrqtZexmB2BC2BRbAmF8PKCaJir6xMIEGgThqYSpZJFQ
GBORNHkMQjY6knId7xJpBb66MNRBy9O/07nNadMRCvA5Ee+TFRJU7D3lQPUTTgQK
9j3o9TeJkmt04Bo4zDu/tQyi3lgzg19jwWfn4WByBDmBW9GailqYx7bzc799r8Wi
Nsj3W/q7h0Njd2VqFScK1jCqe6YSb1LHpkQw6cl914HiTgQOMMX41J1rqkgts0Hd
Q736i07YNh1r4v6+XMq3Fc2XeDPWE5BMg/Z3JHMnQJK/LJqzQC1rV2fF5h+Wd/9+
Z3+ydw2CswlCayRshnh9SXbAhgrMesmpl3dxuoAG/KlRcQEGVZt8WmJ0+lnpMLB3
5Gjqa9JLDr+5UFVpiNlVgWSl871A1TTr4X4TISOWNYpnuTuRNlfD7xMGyiZc4yO6
nUB/5E/JRdH0OKdtOF8NK7m4effsGkSKCdwHSNv1BFKgoRSyyBDieLPBINKC49/C
TEAjTzfNnXBkumO2M2zw4acf5SWVSC7o2lM5XS3DVIPtyUgGodeWqGCAG66iAlLY
hbXyMVwhF58kzQeC8nUcSwS5XtxxflRDMFE7swOBc/dWAk7D7FRoZjkaKawGQ6JM
t4ivk49aQ/V23ls6VVhp6lFlTiBlbmAR6qK0+sZJ03O7ZewH+U0iRU1vJ1Mnt8QI
aAKlATm7Pm6+uCPReGu0UIPVdD6i5AhJJqWAMNTueZV5iaLVTJ3zXU4UcRWgS6oS
xNd6C1XRjN48IQ8UxL9+Hc7OUXKnjqYT5X3zeS1iTCAe9Jsu86bZ1NAftUrqHOUe
hcDJc3PGT3tphAqH4xfCLNciXRl0QJt73lo2QolynU+WMBm1UFXP2+niLUkGbaYV
uGEumxpBlu++J1hg5DZEE35PhcCSt8BrhHvvCy/FmpsfdAPgD2z8RrkfN3im3q3b
hV/OVLCo1seVXgcinyOLY+cIlAtkVrLKsUg97sfnI71xvlpBoMR/OJT+Puzw5wV9
VsEeqF1FcRFb5y+jstMbEG6T+HaN3M/IImdKGiWGj2BKYVTXtLUeQygXR45pE+D+
aS4kCyBarMbr8v6aG64qbRkK7LvaEemTk1BvV3PJLcv9TlFqaa4TkYkb5wbUBR3M
ihXYgnsJ5uQbkCEkebtult17x+7nXzc5cgpoto1ExbTAhgx2c6JL/SJsFe5wep57
ep9XBiKQLn71nyCmsCWnIfgmin8Gj7/IscFHFSB/Xs9OliTGKnHj70xG7jIOPUAt
2jkJKQiNCwVPeHncGvAl4IfIQ651zIvzEVZ4LAbPYacllnguVcbN4pvKCpNaj92o
35wixH599Mf74bIGHmfGXRyEVYEcukqYbLiM/01626K0k8zZLuwEPzgZuSZiOwx9
SIA5nGzsrgik+da1BKR7GLyQ6/sNehD5WUHMQRMhb+Ip53Wxk0vDg0nmCk3euW/L
o+96mtGd4vZ1trd2Yd9Ou7HCvQl8MTWnTslalSM4q3XC1Rgn3j7YNH2+WXiMLbOp
zOmMX/7CyjtuxY9aA3tZREhMbglxvW7W6JuzE26Urfy8kYHh0Mk9JIIL+PvZUBHz
7UPZ47nLiu2P+OTD2iOH8fY9feDOrd3U4wdlRWRERTiZCrT/77LMhHsPf0IglsfI
ph4K+SG9nMUoT743ye69O0a3GHIr2omXZvrrB9O84vp9zSOSTD8sUEODHJnJKQGT
NzWAqszGsKx9bz9y6grMUI4XfR7MmUbEBHSTM+DsHbnbKECM0S6GeqLu1ohpXVm2
q8/G2pb3Zhf74Lj4wrOwKI2F+qCofoF/biqj1ZJTrTHnG/KmRQzdgw4+xckghRDA
r9ZTMJA+I4TxIeVOUcDGfCtQ06vYKiwoCd//3HD2Rcji6hENDNCGEigbo4DSHzjA
3h4CvRCC25n5amF6Lbuoz+4DtqT7m0T9O+GerpujnTrHsXm9XQt2ipa88lclCs8N
wZOklAfslB+YsWnCNK5EnjdjLZjLz5B/Viy8fy8Dq79tFUGP0AJZBE0/HC+yeNRY
4A15PI2T942gd5GAJ1kYiEJJfoT1GjCyMhbAwW3r8HHKaFKECV2x/81FyTTdtfFj
zAnTg3GkDKchmRNcNOsqb84uToKHqSPawdkKNG7040vlT5xJnKPzuVcN7rR+pg1+
BLTbBxMdA2PqUq8luaQ6Hk9Cz7M7J/qLFDYEoUniCcsMvN6q+cNRHycnXQ9tNczW
9xhm0uuyCA5OOKyF2rCFA0BGKx6KlYO4DDc0Un5SjRY8qbEUgXj+IOExR8Qo8+hu
Z9sd8vkLyhMDDzq5oQT+HRcIwwJXWfwRlaCDgjsDlUTCiUHPmttSyn4pFidh/V/Y
H5PRlQdmiw1xtIEi8VRT6omrUhFGR+sqdrvaGuZPsIPC0bQziPXpymgUqmSZaeIc
Q6Tb2PmCRGmG6Dy2+Pl4jsDIwNZfkOckLuk34YDhk0r/8emQxq0VmMisFR2eJZ5r
B3lbhFKqajJ0x7xvcZwtmam4wvbGb7ruQxvgh5eU9+uvFgpXqJ8pjTFoveP+hApZ
hh4HIL3gTNB9nnJ1FdhhN5QDN8Jfo9AiNEIUzfLOt3ws154inPzOQ99QafEeGDfP
fvqE3m3r1iEZm+9S/KsCpDZgtBNokEq7E/hlJ+Ik4vTIevjQOOKXWeS6GWeYsm5T
kJ0M07cTqoSl+bK1OmvnEc3TFbzVOpcORk1Lmm/XNo+QbKWzHiagvWgSfX5D/BIe
830uPFgNIuU5nTQcLyMcZJuqTmR42WZLN3L5+PzriOOTDODzPySAX9aoRcjqjzSg
+usNqKAZuxbPOhZlYt6dlUY+tciteZwAtMG//BjSUEydh7G3oEhvG/DJoa+JMQyk
MyK64x+6IL9ZrDyDDLYPgATMWjOxWBs2uVzvaJPPlrKR54HdSgGrWbOAAKbEha7s
gShOt6SBDc7JrA83cM2i4dOSqoNKDRQzCzXpQIDLP1gtm+fj0zQNIpfIKyDVIcDu
rYXmOtTuIEWuVOMyha9VYhxwoQIyG6HTkvfGR9IUGqnTgWK8Jocbi5nhE3qbRM7L
8YFA3dCGXNhBAkJ2ceDVMBZcayVTMagi4MZcIm9NGkOgbVQo76hSO1LZWoSN4jfI
PBqDeNs8ohU170EkqQ23NKn1bQnYyevMupUR4nsllqcE8eyom5KnvfYV632bAFBi
XH7G+BrUayxkZuocXEPI6hl9rKfDNlggNdDPjjZ3A38+tOTmr682ueNhWKhETlBx
JPI/WxkCbD9Nr5Vd7XEgLnVHWXLIJc85mygi7fbThQ5XeOKiH9qmPR5Ss47HrSYt
AFcF8iZKDQ1JKUMln6IsobPYKxwlGJZJjoz7Vg5XPTtXS4R7MkMIubZttCr1lHYm
wxO587vAP9UGoSSglf3Y6hyqndFNGxuh2xO7Ie/uECshpw/Rl6d9gSmjg/D/DNmd
R2mYZQOq3e+F/xxxyx371/lal/lHmwQUsCC7kxndDsG5Rqz+fw3VMN0h1DXesk+1
cPIqUQ4yjnBRjjrUhGC62awNJGIL9pSmwqcS8xc+wfEW6b9AX0ct8WqR3DV16BE5
+X+zx7Wkyd9wVGVH6KAvqDPRyDXmxZ77mP5uUphIEdeLwrnhtfpb41ONVeBHCRyy
skDLcDVpe1BUZT8KgUlQLDpvMyq6jeC9FYCelzIEmQNSQBWB+pM5nY65wYakJaJD
60JEPVQDKGDKL6z9uyFLjwRU45LSNJvautUloo0xEln9BNpVBbwMvRREErxhq/Tu
w3sM09MxqUif1Pm9MwlfBrnxCFGVhEBR+sMorAKO/MZ8dYfKtLJou76wglo5qZ4O
EEQq23Nd0I3FsoVEo2UHM3KjjYXLOzvfvrkQEQxHo5yG/Bj8O2XjG97J5BGIud/z
xE59f7nvzc861YuyXW9MHGiaYz1exnU2Z5gH3tx/jfpQXUAWT/Bmqgdv8jldoG/+
XJyKets/mSWbBbVEAulD1gY9F4R6mkt078Mqw+8iVFwZiItUEyhbkWRPhY3inw/L
xJhrq4N72vCCyfhLbJzAQW4PR60Rqg72VR801OCTwWDLndluKYPVp7EriEq/J4RK
qAA8ZfesDjOvQIjAPm0q+qjGtUQaZlC7SSvM58SiGQNvTtw2uy51aj1aLJ68DnbS
yTC2BIuu9GOV00Sgzme+WKL7w2Ah/P2IwdJE2aMM1TjM13NuKAt62JLphrM03+0J
s4fOgHt3H4olXZw2O19glO+qD0Etc7CAzFnWHXC7/EHCQqA+CUw2umoElWNmNz63
tLMIZ+sgfzJzfuQmD4QPVzn2/fb+DKZzGSCywIqtbam0U2UbzQ7N6YYq5GQC9Cj0
EKEFvyN2vnCqF+pX8ldI4v+RezIT5PNpKZ1C4qgguYyXnipf5ldBeGxYvfVX+LVq
DkM+PcbOez25XB8cz4TCFdX0uyT3VpaafEeKMs0TmEmxzVssIb/Smxl4kVar6iNw
mGwfiE29Si21Z3KobVvzhCA3ITZdss5J5J5H4jNEPJa906JZQzXXei+f8Hry+5db
VWj4Y7zT5+7vwr/qppmAu7CfpsdRdqbgI8fuDt4CO6yGHkmP0WZrdxH2srCcUXXS
VA6rVKuAXbNpveq+IMMEKVLjuTkr4Aviv+MGIKKWiF7ofEGg70feENMMIdT4eDQT
bDSTLMSzN74H04U7xMKJIdOewvfVP6adcxlnmi3YOcQB9BpWjc1OsV3xYOf9YKgl
njF8VRJx/wMOflAJOoPdUewd+/o+8SIvZZZmZw9v5qdkWPE5qQpi+Ul6PQQQif9S
QCqKevsX7FQOYDVxy92nrCeUvVezOQ1qhs7RT2uw4nxzl4vczZFeRYYRXpSn/8kA
KB9jYT9tD7X/mLVPd0SVJeEg0o0hzOD69UwtKALSCWHNojPfe0OvhCSqvwlcpZok
zrnVx0+CJl0wdLVP6Nb+2Ccw52kWQDfGT9eGaxxdu5Q6mqQGDS+JMz2Mtrmqe9eo
8ncx6U0vffzctjytEV+vM7jjMOTYPH0TANanKZ1rVewbD2jOUKQH/wCGgppU8UK8
GlwA44taqNs9sdVgGcfwDjC7i93/zWcFlGMjF174G5de2ASR1ZRUGwPeM7Pjz127
W99Sa01f7foXlrUHTsZvR5YjiuslW2QTGznkENNoA/HMPpVArJG/RMAI/cTNd0U1
IrwCZKdVmowcwJ6+MNlcsc2BlE9t9zW6TZdzQ6FkslUhs6F4mmTMJGdfuYUgjxjx
itlWt8sxrTMdoHPNtxAvOZQFzwsu7I+P+ntPy0g/mnhMUG4bjVvsVPyGTwxC1WmD
kRC2r0sOM5W1PazFZAZuS055Zq94lKQDBviJtkSZiJE0D0m1VkpZBz7LquHJFc+N
UQ/33fgLME3sK/tbMm4kzUepLlE8ue05ITZNxe+kvDS2EYwBfFbJ8FGCb6mofGGb
ezBDhGEE0IOTEBblahOjC7heQxdQkuvsK2jd67nYlObFEEriIsyqyYniZMXxNjIX
ZGweCr0Vh201yCyejeNweNucbAAMDZ5KtINjzx8Xi5/CSkWsiRBr4DkEAIAK/N4+
GaAQ8kYsK9Q8/5oeO93lpzOgP9ABtR+GoMWcEdk4ksFvEkIL/IhyY9f3yS/fhHkk
ebldvt7mLuVtoLrmV5VZOueoiRP8ClR1QmhUtfps+EojJ+KMj/ux4VKSIljLDYr/
+HIpTmT+GAQMOsw2xOkgylVi+Ei6siVp8ilUACmqIOc1y5pc7H0m0dnQCFkFE3K1
2FNobnHpRplLUSN/06YZK1dr/l0XDa4mo+pvtHOeiRjqC4DfDsh4L8tQzIBj6Kxr
USCzlE2w2P9+CJYmgv5tbhsjw8lFmjqRyiT2w1bt0nPklpTvNC/uQpCq5RKLqUj1
740gtFHTYjr3esSPeuo9lR4MuPTaA6OFDmOIvP4u9JMooGy5n/kMOwC0a/UUEmZR
ItbEN8ZqqQR8tCGNTTBcVPYK5y9P46381s1ZIDcRoN4xol1U3DqgHNz8GN9vnzf4
eZJUepxmjbmnv2+kpZVN0zo7jn63qjghdhM5KykrgsYzvrDDYdjAxHKR7IgwF6dR
lQMwi6r5OmUlJieIbAtxy8kqwqd2Ze7877RnXupQOEtQBPuAK2jqWDj6tJxdYAsq
ZLKhv95+F2G55oBrL9VKO6jLk0ZYcS4m72+gce/T/VGuynUEBlBgE4Iz8yL6BCvq
adYWyu+iwWDJR5L8xMRpwiAxSZx4G66CpgJ3x1/+D5aNTMCFJOzoSFUl5EE7tNZ5
K6RMtB9YpH7LQxfChZ5J2jRar8QnBjnf1kRVEkMBRKm777JEj2jy+02BHRK9SBfm
NoXEIh7WiHKuNRituHXrl8PzutYXjfhLH3JzeYX9MIZjWrTR6ZdHlghN4/Txo0iy
LOxHdjkcAflaY2Nop0iu/FU/h1d2wpjFS7MhCLiFUssXT2YOz6oXmo8ozTedOKsL
odhdt4IlvZgS5/0oqYEjajXyHox7visuHXQ0Y+8g+nWP8yYx0jndZoJuQHgKdR02
4SENSr7j3SZtWtBw5APkfvGzyRmi6EH6uXowRDH1rNkqkhpBLRMnj+mAIp8MWaac
NwyE/sS2tE0V19BQnCh33+XaKqZs2RypfS9I2dd0GejPhTDffYpmNkvMNcA5fs2e
SINO2Z5ZgJ+HJmxILPNHbSeI0ps2LIx/fucWHjOFTSAobGYw5ZdeQFE1zCT5d49I
Xx7eq6nXB1V4w2lcey4cpwzyf2Ss5cT632pjax2UllpHoBdeQKYBGEnCWvZv+9o5
pKyvVqP9tTGfHefRI+WGtGtSs0zv89jypHNTTIAMPCYolmaYZpL/dKEcfn0iffES
eGslrEKRZpNet7GFSCbHMmugFb0W+LEeuScVJ3EHgmgtKUMt0346zZn006bRy6dR
Bo/MnXYx1hqS3i1tc7wsoMlx2wIh8003aZsYHElx88XZNcvXXLJEYjr3ON7P4g3z
OZwg1MEyB4N0YvULxRFJPa1zBYg5dHC4Qtu/b/Ff2OA/sVMvbcmcF+61EwHszCvZ
y/AVDrDZrW1wz+gmrl3VyUgUFINDrENj5TiBvYN5Pxh8zCUs6f7NY4a/V3BfPtu5
2GgPFaF5aMluMRSBkEi8FxPvw1hbe7a4O3MCRTH/rWFpRFXBLyie6EZFQBempeRI
0sw2L0ciegG2XgT56kCigseV3zCxGyZMziJmShjft4B5c5etw+cY6sZUsP4o3VzP
kqOW7V4Ly5CpYlfGJNyqgYwlAJ2XjTyHufNFf9HFJ/FcgJEkNN1244vrSVpI3CGL
ek1mC+DZNlwiCiqMvxru56EjdCCv3VkrbOCHIWo6KownrDJY9diUwbr35F7mo6Y+
CfPhR+56Kls7LOxb0dzpum99j0y8oKOO8IAt6ocoPJQ6YcZX2qmsUOoQKaBGrSdC
9naVUvRpyzb+QqsjCrKBgh9YCzm8ExjCBzIZzc+l3DERYNyoB6fzT/HAVTmvB7Rs
kJm5Fcs1Y1SEXhxBmlDEgleFjcPuCBcgde2HDp0mzNUAVEIxfV4qpvkZziDPDo7m
2ZaoEchx0Hcs0L3ddVMpJCQDcT3L1n24OEEdMeE0t+Ne8FgJwQ5IVz+yS4nMAozN
I3NCpTubWiCs/hzZcBcxf871XESsvqh+2ZBBJ/swIZxkNuvyYuxu4avDb58rZoIL
zGIAzQQHa8MQJGOEqrCxI7WGxG3+aWE6GfBp1wL3w8melwLYLBsxgmb4UdxvqS0d
/AkePirTdZkHNkxhE5vWbVE6CIFEpoG8eG4WD3/+wvJ+bdp/Mk97/zNhyxvrcFlB
zlB42RQIYWa91wPbjaKiIIpm2N/ea9XInjxfqAFPIHghX65UQz0zj80FiROMIMzr
JAoKMTxMH4btygMRdSFlXjRUHMrkeZFRCVx9enB4sNWc+U7TL5tfTOILRcDH8DFw
XMsZljm0VEpKRT0LShsy9XHaMLHmuxTQyq4ZMLbFmSrlnRQovCrVvy1Zi75EowJp
s+BTKHOngwUolfWwO3EcDjToXGSPVtZXDA7YDEcIXYvbi4CvXUzD7lVAB7WfDuos
sBCws3Qoi5cCk7G+iITgiJf0xK/bvsbJWzOY/RwSn5jOU/HZlqzMHAZgTcl2vtu3
zHmajoRMUy1+jjanceQkw30SoSlG8oLHOw9vtnJPM98RFvYjmU1xDcL0kJPRoqvG
LdeqZHzOCyqwY6iXnu32/bv3cCuwR7/jS/KhEt4JUFxARmSXJZ6KMWOLU+DJU4KW
3L+8Uy6XNb3sPGpGEJOt2ddwk8anJeFAttq2cpi2UiFy3hQNvpRi35hKx5Dpvhbq
NxnU0+QTcNkv5ilwDjZ+OecabyZ+hqECebUBo6een9ugVMjNp2ARr0OZu7XijR9i
noPSeOGCM5XWj1ne2+KtFip2TK8a82Et9QkErJjfpHBlxySeZut3tLqqhk5AdIer
gvtPXkFsIyPM73yFRNpF0Ot/AFYdRP6MiApbqgcbEHR1qQZoUBls6d3ftMrq4HZB
7adrDmW+Js9VkiFkR/AF0+M+S0dK9NTfZxBXYyIX/fcQ/L0avLwDpo8WrvLaDxXe
U5X0g+6ZS+JjK4v7uGO+jMCA/Vy7lU/3AYStvWq8vVwghnTCroTvI4oJph5105lR
fYgrLHym9xXBE2OgeJfFqmmIdz1WfsrFPyIesQt/TmqTl94zlf1EiT5Le+M2TpU2
Z6e1Fx00cN8j4Mcls8auPNlsFESS2a/oq9uupllM65PzUB6XMZxg9wSg60bVuMr7
DfD0tKFxwuIYAdI1kEQ68qYEhl0bdtue6PfEnYzv1QTpGbnHDcy6OIVtXLpYDoxB
sr+HGpRhEgT4N7iztcNls+at2OvcF/sKhNtQlkWeCqyMPsBbQUttJETj8pp/8rff
wDR29QITvyUyZMKxmPrKRlKImxH70na/tFD4Hyl1gCsCntt8bROw6nMnIo2JfZ6S
3B1VDqmKf9ZpQ80VCJ1LoFK4jj9IaMTFsTkuF1BfXv1JXOtWFXKQuMa5M4iakWsW
meJa/hbgwK0aAkCCopso8FcgfeF9cLWpgSggglSuYQHznzhBGlhWZsxqX02m8HIA
UsPo+5f5jxHgwPHu/VsEAeOjpMiYCg0PBUJykM60yPNGUWLLE3mmIuWCj9DQiZjK
JMOKaCnl5sP7gLLKeB4wKrYIvdrokHl6c4zDZHl0uMG8ATQ6pR46kA7VlXM7WIN+
SbdGfQwl5EREMZRUp633CwAZ6kr0+NZdimbn/idxZSWQVXJgxVDjkiS5f+7LvsFk
XaAZWpPcmAflOmJ9vPyCnw5CUxFY8bx6WO9cn2KbyYbmcNjjTvIGmvFP+oW1W2uD
/mv8Qb9YSB3YMx9pjnS6VBXRuKgLJ1fr8xE325C9mFQslMZERupTcKxoshBieUko
h9m3PNGpct3l+pty5SMgqZktMU0ut5pJN5PivVS85IU3/tJrP+QxvFs344MK1Riq
Gk4kKHdx2bFBoOaETTvQYxBdiWnsL3WGd/iKu4ragY2WCKxu9ZqcK0loB3d7oa2d
7Fodzs7+mTl5TLpnCaP2HXvruiVCn8tQrx11V4Zp38YMp25FCSWozWk5Ct2ATPb4
dKtsVYtT+GedgzXwapa5iEzCvXtDoG/GpziZy5x0xia2RBXxOx2z9hRLdslGMk4Q
QB/QVigqBT6fNOgv3aseSBYttW4H/rksbVIGlK41ReQp/84xepuQCnwFcuE8jD4O
Q7DNyuvO6G4fvkIsuKnQ5QP104OZoXhvDjavaMaZUcdWZKE5wQwxuSlzIyp9mOVm
vx80pLhpv9TrCA3LK4/GIlSZEuqD/RpwVqIWDTRd2Zn456zaPd94QwD9dMUgIRV4
9PhNOEUXLNe/gFZpH0W2HGxe2SCBwtMUJsXHvbeKUaQcF+bjjHdUQou6JQp9rH7F
I0TkSfmZM2ofJfC3lyEy9A2ODFVkEXVYqp6PzJ/27kPHhFqg7MmkN5eti62kxsV8
qcV1vlwsm8rQyFoqO2aSJuhtwdTpY3dAlWwPdckXtr9GWrN+lLFWNKw7wZ/gedbd
+wdCQgNXNAVi9R0izwCEmkFtp/nCxgYGthwLnnoJPktttmxyanupfATCEjjV7M5N
tuqvyY6ouzfq/7AbVGkSrGlUocfeGHzSBhorRVtxGzwDDlGHp0zdxaBSYaQro64J
pk5pMpma04NbCuHCH2VkbVw6CYejQV8OfUFhR40sxk2rk3MVeaSm/0tc9uBk+soX
42Mw8EyAZJJbB8PbHNNDFxeVsJ3kbSSxUoNTObry/gdj7vdZMl2YFe7GT1u6p4U8
Taydkd4gONgrc3SxZgMNR6YmAVXVLKysv+YRWtKplS+Sh2Jsut+YRMZyOFfCZ9TX
6SOKMFfanvRtEzKs10EetLia6VxOBHfUe05HJEN3w8ZAvYOTLUlsIXhit6vpDTC8
bz+tZnYG4RWsjoPW48BY2O9IFkx06okhyfabaZY+NllBJJVF2WK9hVT3B2fw3Cs2
gPFxFB7oS1A7G6WNbs8/PGUsT4jJs/HaVU/67oQTXKM1b51ymspma7jO+f3tpUbL
6huRuaROzapr30nbZJRCCJEl5oBUxpUBfufLG1+UjgzjhPGCoxX6SI7wJw3kEJLp
Ssld/WlrLwIvAkqR6ew04k4HvoI+wHsmAI5FjqpR/9FlBVc6AXP4nC/PGr9npVP/
wWV20pgw8oS6u+58e7vvlDOpC+n0dCDAQKsTEDSIhD/JTwKMx56BeZBHOquqOtAm
zt/B0srRQVkFuRrJOWOQ883C3GEqQLN89L6fNu7xrU8obP3SMD0XQx8uxHIK6RS6
CNQsmV6p8HOTXMLHZNMYd5F+pBIos8lrvDEP/cS4VnkeMPkTne5oFx2jH5p9PrSg
Q9Esh2/2tCQyy/m2Kx/7vKjJhzo5o+KvN0bvL5SnDROhJ5IsX7AAl4jjhD7gb42C
I/OcoXlGxq+dHg53XusBqydhAJb6x9SuGdeP69gKfZWMPxARmGGTI+iBaAaBD5E5
6dH7NJPs8y2PkL+bHHVb5g4FrQLVpX8rhxgZIPnItVjiuwYk8oKRK63RdY7KcfgF
AQHr7SFU1DRCdwf8eqfY0J1rKOgvDPDYEqLuH6mvlvwFvdjg7s4SYc478DNVMAyb
Z8xgnxxgUt0+MPbwqdZzOqF02+iKF7joOG/fweSivfWzyaePmqKgnZxq4a2JK+YO
ZLaE69Qrn5ii64XIKeQzlbLnx/8/W7KOm93bGutWolHMWglmKXZ7LmCXuT1omfM9
38BRAIJHGv+IF/r6RPU387j2a0tWYU0LEqXdnVGbzrWQ+FuXqDmaa86IZWvp6uqB
2qBgwf08qFhHHya9yUjOkDp8nSZa7aEJCy1kFyVx4K+SeJI5qTryPf+7bFRxRw0N
RGji22PvGaL6BtiPyyyxTTbvhnvuRd7zRnqShk2vt7+TNrkFZSI+EJVX2qUCMmwC
WjE3WImG+WoLyagCmN9t2Hg+HSmnYoGurL3Ovl0eIEMe1XPFvPNyIPnT69tMdFIK
U/YqIc1tXgvtbXHCVjT9nSfb26OlnrBnDDR/vk1W81rZOOkGr1qOjbQ5i4fdMo+d
r+D4EZQgiLxYY1tFJDjxSgCezI9j5g3gBWL1qyV6bq7EHOlNm+HwwSfAvWEB8lGX
CRVHvmV868YHxLtUPUpTljvicHLyG3B5TfxRkKxaq0ZEg4o43dw4OOdTuinUWd4U
omihg7LJAlUGyIv8RSUILAvK10BvtFmGyVbodzJHm5n1wUxeqGMRp9sTnLca/QGZ
mBzowIUTautsEBtnUM5pzKH8SvsWGvo36KjVgGAMN+hFksmQvx/jVnud/KJ/6MKC
NZ0Maoitk4HvYfXlE+41pC4FOFps/LWWztqq13NfaXM7trxI/2rhO8VwtcymgZvQ
M+VA+R4KXW1131lVstRX1kwZcIoDvsN6bqHyeD3Zzj1Oh/JJy02wWUx782UWSfO0
IIrjRS00tShRLOF3l3JyI0FC31SWgPIxuRyrJG7CiTS2CDrVb4v5hha7qaMivzF9
wli5tLiTPf2UM9YFcEdb62mVt4Qx0Ms+lS0GotkABNsiQeDTp/QCfaIYHgTwCnE7
XJAlWlQ8/Cxp9ceMGobZj8jVKtUufOihFo4s1aupqcBGYLrG8fbwUF1NPOWglRl2
jskAPAwlgze9g0jB0kL/3GnqHI3PoKVTOITzASJcv+zCxNOaQHXej8LuwQSZaM7H
OYRM/I3BfPJdoIMCJP4yXKLfd/m+5VkUAXB8u5wGHCQqWpEPygOaLO2eYsNg9224
LMU1TaJeBSKC3DAkYg8exVmNK4lJzibMddKqnD2hsfWRKmU0BiNiDNCuclbEo/C6
n66ktA+qUUS/+10a+GhWfhr9PsK1AgxGAX+QmNh0Zu3hPkBkdAO+KScHOLry+hCK
xwp+dksa1/JEOPClzButrnyK2souFntUsGbFRMMsXE/ZZq/h9EthNF1wA1k8xzDt
/j99IH3sijoBgeeUb2GSwqfprJcMLAOkTcnNjVFpQ4dI4DOCxQWb1BwwKNOX0Rcc
tOrdYgJ/rN/J70qX4EJd6apGgdZbbubqus6JLpxXAJBg6F9xX1XE4TBL3HJZnpap
+LJeZcNdgbU1Q4xpSQKoBlUdvl/dyiVa1WU01B5Z7kRCG9HJu6VXokeWstruJKZj
yrOyAV2f7KwKyfWpwGcHvsVV2c6XZxO92BmJWi5zC4DfN05v3pbjr5xfzXxavR/7
ODajcNRlSj2vrdmwFQvZ/gtiOtBdKUYCod6s0LrMdJ9DLi8m88w5ipApgt/xvLWs
xAaPIoUXcSaYex8xyS2zvCo5ZdjGVi/2ltTukpvLkyy8u96eR4hSOIqHhUQWmOMO
oq8V/0Qdv6FK8MJlB4A2gWWvZEnEBenFpwkqwR25AnadpOSQhBhKFP2NRlPqnZAM
1FBVXa5neZGRFYZ6tIrs9d9zRN2IUw4If5OEfHSl+fT5Z3wAjx97LPI/ulCEEvN0
O3aMnT3V1tVpaHPIQ1G8tWAztyoqaw6oezVuPtujZFP2OztSCwbdczPJH+xTDkqG
WdPpS+Du4yZImYNHnaVfw6fQFdAwf2hh9N7GczfTYRp5sOY/xEPvBo6VGcOoDWRV
5dDvqh6sg6Z3Nt0L+ohlYnDYqX8FjsXEPozQCMb0i7ITQVsdN1Xsxr7COQQYpfl8
GcSRzKgad6P1Z85ChVbuyaFyAPny+SaendJPtFtymMtN6napv89j2ajb3XNp7371
bLZdv4/zRfFSZbvyAUDe3x/DD8pv0giuyZkMBpK1DcAbQ/xMGmpqgVfrJHyCXDag
6s/+qBDmFnrEh1X1wdmqrI1P5j1muphmfi1mnn9H/eKVeTFVcuCfD7hbibzezIgn
nnXWk56zKWNOOYjgJIOPsvKTmnK17FXnoqPLONTD3P+envYc3RPEWsqGrV+K+/M8
+y0nlDycH3G2qiREE4NVNRmZou44McoqVu1JmoN94jN3jgG60tYM/QeKAt/F4jNB
SuMHp4piuojX967l74hUPaaoNd++4TRlIjIqONcCHqkcjrRwdck3p1fBiWl3qQeA
3h1dFALj4x/6yWbnQG/oI4S0Bo057Dr/A8h9LMbpBknLRucen3wN313TeqbAmtwn
pGAvlyhhLYtHgkdwhDCxczGlqVf/Wotae5WTsi1hNnf6EEcQQk4IgIInswpiL6O0
EqSu3vmdgjindpifVxK+I/NaFCc3VPGVrjp78QYv6u80IZEfgjZ2e1SGsKDe2J4f
t8jmCzEwLLopa8BZRx1pHrSeGxsBR4ua3qDxLrbBSCY90dbSUNu+/srH3yi9jEvx
f6wMA+Sg1KDUx93rCOo1k3CNkPGGbZOG7Mjvd0rHow5M+9JNmiZS+aBcJBo2pnjY
ifZm96L0iLlBjR7P1Wfo/a/kr3SXbeTQufmocPzuIYbGRco9DmXxR8xGMRFa4m9m
/Ltt6ddOHzBMpviQ1zvC6iJRuF+Vi6KgKIq3KT+vXeJCkL69bPC3L9Qwuv8l6Xj4
C/2KAEUfltCCDI+QGOAkQzzprRbQY2lMC/Kkgh7VQeYB7d8pMh4cku6t1LwmQT6f
S4RTFxWdFn606PheOepFdna1OmKbLgefIfMZKbs7MrYZKdulYTAOutbqPE2wXVWK
u/IcZlEIabITaNN/UKhug78S3ClnrgNjrxgVjuHLtM/L6GBx5DVXOZwczxcJydU6
ky01iI9irNV4RHL12eGWVIDprc3Vs50HVxWTjE65lVP5BPz5h0op4/MH7AUoRyn7
9lUj4PfVZjg0px4xyQdi8H3sGATybyj7CQfQojadXVCzlPQlCXYMuSGt80VBUdGO
jeLJFPzfytFT/esuqbV22RwF4c/pEOfSgKTwE1O53eFP2198D7h7RQ93IEzb2n9Z
Act1N5J+Gf6yLF5jMG3OezH6IFhC2riPg7628M1LFEJlmBZX4xL3hmLLsziau+ku
PVwknkEN/4JtJgYcoKm65KQVxFgxD1jlh8DamulwszHhnp85o3SvGccpAoiXxJmP
ypijmtFYeeAvXEppYht5fRv+hhnYHz81sCknlpijBkHud2EsmLwfm9ay8F76U5mc
Ofnn8Avq0sb8Nil8m9FMd3R/AY7OrVZFZsdJDDb8G5U7TNPM88WuTM95iRc4L0QJ
RrYWui7utRgHW4NGfwZfWZPh7XlnXXFpg3VRjPIKtslozolRAer+iY622Ti2g9/r
vu8gAlpBQ73iNgOte586kxg9SjZG//663zm8LmAzcQe2rPwZ0+UjVqocQJrW7zcp
rhB9BUv/2f+tlhDWNBacwwoGDluKVnTAsab1eoW28Md5MzSZSx/BXz/Vb5MCLK0Q
9vfCvD9+sKZGzXSSkxDyKrnN3Nazy9jCs/YbzDBVWvELvi3w7n8rQvtz0zDYO8ht
jvFLyqnXguvQsbdf3JRyxqesyC0BzfOZ1eEsBicm6n5bW+b+IwYYJTq2mAmdo/DP
G9nJY2n3QfYP/n7Qtb/9ldmUFlDj232trLae/WcCMIZi6uM2qppJhygySYa3Vh9g
JelRuWYbx0TvEZQpnGp08xvl95ysU3iKL7k2b70fm+tEXK0RAnk16PWTfwIOOTFp
EilwAsysMnrfcmZXicMlZ2CWSxXzJPueUntVvf1d1C0hJpNxdjSgEhub+FYHa5ZO
jLq0kvpYV5nxdmlPWRMVhKgmE7puvfwqDv5IGv6vG8qsPyyiiGjQRkn8R2VZZ8pN
zKQUCLV23yPBX9QxMCHYOOP1Foen26ETBOl/y4rH705QSysvm38c8Wr9iZz1PLcN
rirvZDb3A6raNHiJRevLZYfeaMq3fyBiADfE0Z6d4EMhvB70yatcajM8a03H3Zwm
U6uFaOMKW7Er1+ccx69nH7GIwlvjQWqof6kX84gfV1LkSk7WrUDwA8eb2RUJJ2Fa
VNAOpi5tHQQ95prMq26YEipNEwBwgUms84TAdMcHEFEHlwIWRHkBLtLEYewgC4hU
m/EIweeOLnabRrKN8mI/t6GaqmrLKiAavd+N9XwR3GStllDhkvL5THpfgQpgmVTT
Msv0tiPq5fAqzitdMfmA+UEKK0eS6bH7aDg8h53xbF6dOTN4P7ifbQJ6ncEYjnID
lhMm95iG5d11GzndwxnyNe40fANu8oVqPb/EoI0T8oxEh7EYFFpO0RLKO04lGQD8
aDy++J41C01jVeeIHCPCeOBj9gYdpqj2DPb/BekjrWTZOPJmdpTxQf+b/0xzyNgW
Q9OeM8XFjqBqkzAeGgJQwdxpSTCEAbXoui8aTlmU7Oo34m1X5O/0RMUuDhTwstlV
RFOabCIsJYaQ9e9LvS7rOqwmdDfgOdExUZHjYaSiNZ/TW7YIgh9Lq9oCQ1G0G1pS
ygFvXa/IhqJD8cOdz/1N47mtxzhG/b2qrIwzq1wh1Qxf+9vmvpjfY3dlvRfGWX+C
AixCn74npEDK27bAjs46H/fOjwJU5BTOXhZp5HO0yGk55o9h9C1148pmqGkXO46o
FfgQdo3O7tu/2/pSMxqOBsMHfY80INA8KYeDO7LVcxANqGgaO9WpWpRe9xrKdKbY
5gOjGx4ubYb/OaKEpeq5S1a1T6M+Ug5VC/egQjlufSIO6NfKJnii+/S/Ew43mPDW
p2rVpKjvyisWSwXF6JlPpz7PVQCSAg5OebKd3n0nsKhFIhNAyKQTPox2XCnEk9Kc
TIhVkm3PG4FFNbbgw2U3MXQEooFnVV7rQEeb4eS3XdATcjQblTUXFCxxetXSa6un
np9uHXA+toHvIUu4sQ2bQDh4Q34F8pSyrsGRJ9cyiX8BiisaYWAIo/YEMI5o2Mtj
J0pujr3vGl1vny8OdryqWCTnXHAfQDDqxnt+XLRIknDgndaEi/NqwqH94LLhaFcS
Jok4kBTtvsejsD1aruQeRQxf7b1hJ/cZJHLYe+noosEaLa51j30IPp05a2yvvbW1
UGVpkmN/MyPjUJcD5UqmCN5Azer7p9N/p2jjDLWKLk7t9gcrkY4sa4TydPWSfuJZ
5jLqScGxHYncc0P0mBlx7KQlDPNU4+/I07wDLMz5U1Zb9B5fENqEGelaq8v0RNXb
E8gpK2aPp+UAaYgvGF6moA0OmVU5h0PBNcOg2xTT1+S0mToMES/ii9UJbiVEhbWS
5CkBNsRJtUXLO7oi0UdGvABl6OD01NszbVCJiYMvhnrMEryOPGpUFOpl+ICtCv0s
w/wayoO8FfJTuNQUWhslZsQH39hEAP5qaxam9CHkJsNr4G+I4BpvObVMriJwhjjb
GNJFmONvl1f0BzlJAOEN4Zokq4CjI2S+U2otn9rcc5vYyyXAOKyHfL3SAdvNSn3F
5VYvsTWrZrx2W+lHoU8KqSDkS9EaJrDqwSMB+mSG0f2+WTyPufrxzcnRY7rX05i0
n/8X1wLU8c+zSRU5gDFgd7zP5dEwJ25tBVoiFAP6P0ZP6fJlYfzjDALutKahOrlf
6rRADaS1HVh5SQxMKa1qj/HcK/EoGLqkkSL3h+7tq5Zm467VXnHXQhIflvZnHP/n
MRkYmlPMbAGKj0oaiR1c89uMX1h5uXpqUo5UJJ1Im9EGJXpXvhMSp/HFOFS+ijuG
W8fn/4yBsDmHcms7qxp14vsrZaN2zsHmU8C6je8En5+lDfXycpgbNQ2TfWRPQ4ul
nJd7YZE1iWuEkVbj7lgmPSy4L+MWhne8X8O7735S0OOUDAGhxP5yTmP5Z79t7yWL
pFWlbSPaXiSPvHFPBJN6fYH253aobwXP8MFdr+UQSP966wDGjDZyCjMavGeVFaeh
o5USKBihAQQscL12QCQpQpU1Ml2Qj3YXWNQ9Q7bkRd7p3+Mx8Kdfk+h4GchFRs9b
kajU0R+HhJasxY2plpfJHqCPLASyUY5O17PI8uD/AfWFpsl2cIV9u+ayjRZw90V/
+Uodbtq+6LC5JJlfwtCNah2HmiM8kXbmOpMqfCx9OQR+m3s3vts+uJOZWdcLDEl+
F8CevJNWRo96mUUfb8tUKWXUywykjiwjONAaghF+xvavY0yatozfrta10ly0EpVW
k870E7f/g9T1UBecr/i0EhzOTSPo/vKgSK07ujrm20K/Y88iz4Nx8RuMpLk4TJ6d
Z2o5rplrUnyTjWAdjTvwW+2U1f9MuiMD3irll8xQXJRe2yngLvXuDteuZ22klpOa
nPAhEnRdTSM2OylZwVlT5q/uMqyWmnxw/avHbORaTAIHIFz16tK97ULQnudNakwG
6t+f+zl/cauwmI0lITAw1/0S+peOz2pNFVqGoFUYmFHylbzdSJ2KkUf8uJLPdEp6
0iBcczrFpPF2x/iZEDRXkBvBaICIwrmxPgNX5+vt3/OOakY4CMs5QUcO9FoE34tk
SkM1WHNTkXzLcUZ1flMgR+eQBC3ghz1eFny0ktbnzkgKFMEh0O3xfxtHqxn0DJ4A
iiN4Y4USi4cI3jB1p3OKFxBmKMvcwrkOQaj1Ayyo86GtayqlkinmMUocFeIXERWI
FX+i1yRnGKmfka2piBlR+j/82BEr/ayuYIUtjKHY+jfCCrVpeODouJZpqarMnUgb
lm6ZAbbqbTwmCYjJfZfhBU3szyMeaiJZ3dBfQHtjiG2zLdvWw5qGNfWwjFRIMAvT
CpyTls1IhCKYVOVU3KSMg1Bi022HGc7EMgyD/lIDG29B1aCVtLkDZ0FuB7tsLopj
iEEiGMxOo47bMO/Z4IhilmPUzDiVPs8lq+vrAfjBStE6WRwDvMtiP2ZPZ8HJ99Qd
BoiMFtBMR/V6fuJmvHPZc6xgyoz6aGuXS5M0JP2ES6t4JdESSWFWimOEg0NqwVoP
N8MuWVXByfBaUZTRFr+in5t3kWiAGST+04Ik2Rfb550XYlcoBo6Mvs6JCCsGwPKQ
0Iuz6v2EBN/dx6xXwCWI30+b5bNXJSJKygsU+fuyoVdEq554D383BQF9v5UhJjCc
hfIYleTG2Y7r9iBpAyJBRbM49fbW7wfxIi9RhQvAt7cmO40zIO7AQkoKu+wF8Oq8
qEtTzreQZL14+zQzIV5TDlQ6GGZzGB1F22sxFPcF7wm/MCC4CLw5bWrZC078RZ6K
Zj3WddD2eftNaC4xBHHbrSBVdO7kyi++YxLCqnQtfGaZKCrf42z6kFkaYnskpTI1
tD2XKeMNASANJNTc5IfEsjlX6xG5U3LtHjvSGg3zhqrU3gavjLJF7JKNJKjjlmFZ
54mO0UBvioTvmZ5QM0IClJL0t26KGbe7lW71nP4UIY2aXlHqgduYaIzuO9aB/8+T
uQLHDYG6gyfRmCPUY4X+WXStEwysRZvP6EXkmqTKFJe3d5IRlz7ninAGG5aUu1vq
0I/xlK8xBps5+7CI9znJRVhzuGzyXVn6wKqDZtWlRTzbKc6NenWhniv6HDDmqG9x
3QYILqDweIeS8hOmKwcgYprQvuXudatM2x1M9ToRTLSJbxI49GD4gtfjGN8ufSkU
EBtKvIkB9nrlm4F7KwqXCE3ePTDXRsxxd97TP42RU/0U7grLdC28CiGLI9zuvGqY
JU4HW42rU+busNxOkxWY0/WFxSSIgH25Cm07A3ieR+NVXCckNKFEquJfKCdHnfOO
vEgWKSlmUlUwY/7URrDR6mJF55AxucuDld4ymk7SNTHseHgOb6waxWn4Vl9CnDeR
w7CX9VNkz220ffvHjB496g3ib+yOcR2U8q9RMPR1IqnJ86B2sflpVCvTIVEJW84H
e7kUK+EY0Y7wDHw5ItxNkZtOxui/XvQ6aaTpzUHrOiS0LOz5fFurMrjLhFldaCJu
ssF4hztYyN+HIvmZ9wqUYgPgpeTHorF/PKt/zJow2LDcwb5zSpg8UQiGGvfuZLMF
OKbfRs6abU5YkaQCHUD40pkpn6HBR6NTZbbTYWTPOe/fluxMLGzazh4YFk3tSBOp
+JD+1zYGjPVdmEz7wC4fu8RK++ovVJN6mtCMKpZUz0Duywdz0JnNFdPrJauIijpv
drrVZP0UQbCpwURFQysb9sy8NVQjoLne1Qybjxdaf5t26bde3Bv/Kf0YEy51v5Id
HKJmMdzJfoBTuvMBGzJL3UDF1LlRGg8H7WDE8D16z+n7uTbzSRoCtMZV/6bzdUdb
7eaR8yoz9M0nhi1pIwoklvxuGnfoJxNpSsr2qoi1c8tyYd6WpTP1g2mtIkB4kB+k
ERn027Bc3fvEuC9nF6EpnAmQX9JFyC3o7GL2FtR7odVH3pMl/bgJoCriSyNmsq9X
tW6QatJrGzoNWpsxQaY4sEKko+dH9UO9Qq/9nuU5Ieq4fEVE5hK9V8SsFI8UAOX3
RT0zX+zagPYVKJSZPBEvKZAfSiZR2eAHGMVicojLaT12qWxVRWDOuOhLkio+IGdV
cIly+NkTUKL73nWSfYqndUbiEVlfAQAdE0x99qB96vKB5g/xfizDyLl3jNHOes4A
gTISf9KrXePRmWfP0V+kUODkzOLjnpGoxUhVgslMHkgyRJI9s6EewrV5MLEJyuKl
X1eVwa4uDHGjxlnu6z07qFD8cZ8KO+BrxFhtv4BVUI31gISwje9GWOKky46kfuC4
Vavpnq/eUw6J1EqQE7javmaZgRKgc1XegPqym7jaFNFnD4ENCRvyAm/4ktUIoVU6
FRpdbguPOAneFVXQd7+tsmrCXILpJoENCDFdd7bMktf5Tp415RU1GRCzrdpbPOoS
d6fujvE3uY4vbez5cqdqUHz7mkH2dP7XN9lbm5iIlUHxfY/JYNvJO0FUyEOZgFFg
I9Vz2lebzppsR/j0EQb7GheHY/mcIgtb14sONBM4mxvXNHdw4MlO8PF7agyD7amu
XgZtAt8BdapBrHM0XPeCS4UlpkQUWLSc82zUNA0jJX3PHBJiT34wXhWUSrosGrN0
nXympOYqdzoN01aV1yT/ZQys/UZpsYFJDi6LOEVDBk4c1/VQzX/CGuJDqXOObUdG
HBj2PqPMV1ihhyUuG3vtIWPoOMet6NSomqpNENNMWeSXjK240Lmsqmzn2I2AdQs2
unuCkyKMyd5pD74IiHr3cUXzjrxhxL+G76hdruQmfDWbFE8V3GR2j7FgnaqsL9/i
T6mEiyY0gDZAXGigGhdEOnfPIghceFL1fgwEg29uZ9r48kZngDa/V55fHk0GzKo6
C21ws6cwjxxWyHpOFdvvlbkvc8qNl53DfLmTOrqUr8dI8j2AQ2nXen2CEri/+Vf3
IX6nuIq2ClImJgmfKIBsHCWDoPM0WMye8ubCxHgh+Gnky6KQcfXIEbcJ81RcxbHE
YkjVD+J7tF7zsWSJjIF4Li0ZaeqlyNtaBVQaakYk5PIg/E2vSEfRZ4NUzbaGFEeY
zZ4EK0h+JKj2io9h4/NhUL5yTystxHqSud3W8kGhY3wBXbUcfEAv/Po1TinncdGB
kMzwNyEo4gHjAA2LsGMBTRjXRPZ+1dIYOu4E0UnJ6z2M0QoprWeTnuJaxaf0zinl
2B2+ROI2DMaiRRwgz+5DNBm5Qi5PbhEoeXEtwcvxTYJ4cGpkRhszJuh2Gih7FRtp
13iVS/wt3FO9X4KOUx6JSIiTl0UuCdl+7S5DTR4LRC8q/H1sDbd3NV1Hu+QGCsDF
xCVzT6CeeimhTBmJLQQDmlffm0D/bltarBHJzcjS9C6ibzobGhlhJAarqXN+8f+z
UAa5T4wYPdnoEfu37eRDYF/lp3QsEs+nDpYocBnK1xxRa9SM3qtoJtRzqWQsYBuh
uuxJKgM/IgTggZwTegNmNgfBCkcCLnPsHoSHptvm7PQi6XG44TDJgjLgKIwYBbxQ
4lxL1FvWKiceyk5AaLdC8melLH1I5PlWluJIhzuBsn2OFvNdbr+yd9kYThO+8gjh
4D7g5gWMyhclAY90F4If24wkEL+TR1CcJjV451sflpwM9dAfE2XC8PgvdkzV/JVY
98ES4fXcHizz3OXTpcsh4vFuF11+Z7jF67vCOZqTfA7b/0F4Rmg5SoNzo7ZLm2oS
it1a4OyAA4Ot4N9oOHLyEHcevlinf/0ADOc135H7G6W+wiKr/GJ7sQgijH5ibQBg
m0kbVvovlreRody8RWBizEnsu8HFH6+ONiGQGgPRl5KJeevvE+Js1HAbp0TA7xe/
C3Wguy3EdY3fZ7qtrmDqpirWUi54Q9qx0bThaafiZ2GCfhpAdxDp6vGIg9ofyZqZ
lTv5kPU/NSf7YUGSoevnj9ajPXuXmITTBy4jqd8qcfOoHkNfxfzQS6SeskPuDuYw
F4cU4GbdBBzA+sHI7+A2zaC8GWxabAGy08Fs4kLIGFjo7y0LI3/KIi+Ib2o5PuKX
ac/eSDTAR2fc6ZEcirI2zCT/9vS+nKEzSIvLXpwPv6Tv+UOMzNVdsJHD6wOYRdGe
kbxj4PXDphdLFSGiEnGyb/l9mYBqSrX1RwDklglGvsNHWFRwSba3JGT8EUCZ4+Qy
u0Vt8qV49v7Q4+SRF9EplPW5+MLPRjYZ8GTeVnGc4c4HFZg6EK69kCGcy+YaBZI3
KIu4hdGb1DWKVJSu+Lgjts/7Gqe1NLmEertpO/l1KbnjH8E2QS/2i5kgs0gNsl/y
QoGNHrr+RUE0bHeOLO3WSOLD3mM66g2Le5vvda8OQGrvsOzZ5XHPWdigwOida+3C
Bco5iFY1y04jqc85YqOxu9sucbOn4GboR0uU5B5uf18k2rTSX5SOq4Q1imRqYm3v
lIawUy1I4199QJsEqbk98psCeCKIdmzPpjTJa1SdFTcC40iYeLtcr/3NXnK7Qruy
cGPxy8j8QBuar/neJtGcQY2xOoQ5OIKdWBJv4BDbrzVL1qGsiCx1aaRZSQxkSKRo
TFOdlUoSG8X5+AsC09Q1+wnY/mPZnTiuWoIL6LkofdXJItw6YCAN6LhRycW4x6AI
S11J0glisFX1DTCYM4fBeIptG/o9he/ANeUgDv5grKw7yDczqTpgDqfsjgNLaHmI
5hYpMUEgmzvT98m5HxgEdCbK2HV41AtGq41meQBPOxvvQ7VA5y/AGri1QQ0RGz4E
5+LH6066iAOMdfIaXqwcmyGwQ8HwTJb2u4m9fOZgj1xzp/u1gXWt7/brOWK8LwhB
9INNLnxz+wpdeUYm1z7hrXipeJFmEF2TSmQKHmv9GfSzbvPYDVyy66m9zSv0oQGu
LRr0t6lZahkCbfP/231DbRfCMoqwENBjSvmI5e3do3H5axBjcJPSumsDW7tseRd0
9Zt/swnF4xinwXzmOUZUPWt18F/m8Tu4Laa7JAR9SGjCWTzZMTt9uuQJ2Sb8J/ap
Qlvgzz+uGtrSAuGH393R2reKI9icN/+7GtIF5bjPiaUzOdzhfZhbS54y7QwcwHCx
PhXyk+KSUWEIb1BuFpTfTuBTM5SB8uFARA/d9b3Z0YIST71xC7ZEsgpuB1K5LJ1S
kv9N2kYTL2V41/YMHtb01+HOYr7F9/WQ9GIl26Tvmw4f86exEscKTDulFjos3zJi
C7YBLC7gbqSIeGKi+/3UyryMF5m/nfZh3HvGZJrpbVy9rKwaPYs0IJd+q91hewQS
xGn25sDM2QaKiDJc5lCfaZYdzL8c7mss6gpnRdM6N0w4JXVjZPzwa2BDlP42dPid
jIkOIFwuSvUUFcq0gaQJWRx5sPl3t1ir+iA+KzW79gi+atXJ2DMfqDipHgT7Odnn
Ta2BQdqrjR0nviGaonrhy6D7j2ckfGczenVBfams/sXXfoNcfcvsfDpdYDmnD7qO
G7edd0PhwSDSDkZS2E0W4gxU9hCts3D1iXji4zBIvXBKDeWs9xKiozwYbI04CUfI
p9+8hYR39qfb62dIF9H6N/VtcnULwwqYJM0ro1B90LFeeLKBlJz8/iCx7JGDdMCm
jMkMaQfEIuh3RlpdmMK+B4ON8mrRs36OlUpbt3CdzatKAprPaemgeUwoqxptNSer
QVTAN+PXonqMCQGwnszjXlfYZXYUFNmr95NCtfZDPtz2O4qNgjlU0OXzWX9f25bI
P1cq3R0nhH87rOMf2FFL0Hkj51TpioMEhxbUfbZaoiG5Mgz6V27A0qifMoQBw/Vi
DPLC4uhm6T6O144AcooWjFEY2Lt69zTdiYhmBdgMufqxDy59be3MjjNFhjgyMaz1
sREHBZvpCadNJiFcru5ZFxua14fgcXhZWnhNUZI4zaya8C83WPsp9qFJ2EakeXnI
XR0a0Pm7BMdQhk+OC5TNB85lHrqcwBZOPYJvu3sIAuqaIblOc1sLR0tKNVMMrufd
Y/ygk2eoFR5YoL6xpubGJmurhdLJHRNDMlwexkuYC/l3DQdeKai2ZAtF0xoVDr6E
n/RY1nytz7D+1MY5kyuvnqQqxwh3U7p4Qj40KOgPAILZDRHH+M/on3TO4MGizcAO
3Kw/jwxbkFtlQJ/hCnmDWu7bn8xpHsiiAtZFYo1MNJZWpSYeTEPmsCPLloc+tya6
wevnfMgLtNkHBjjplTnnrNB2a1GD2fiBjzJU9vGIIlCqyx9Xc3ZhULCJdSSujnso
BOKCr/tfmxRJXNcvb/kQCF/+Dvzbmg5QDRllnSelCAHBKmVPfc6ky5uQOKLsNbc5
9OWohV5lNnrVN2Vcx5JvAP8e1O4r5lxV9GAtuqcqKxgiHPP64OlJN3pNQduPlrMN
kYToKQaU1Cx5SxSeq0UDvHqzIztOuKCXIX55iL505t2o1vxtXYbkm/Vhw34RDzOz
vwXEY23JZ2xV1pmRplXe9uvHkhpMXASiiXQNWHQYLJ6m5geBB5u9PDY4ylnxzXkX
ZOE23t47NirBMfkkBj6HheBjoiXqwMMF5Me/d4isnRZAr8Gru6hiMUV65LS8+Qqe
N+XYQe3ST1c+rOcWDN8xQZYdZgXZq8A8zIkMHFSWXwmG6nrxjixozG43t1pnrP6h
J1LugMx/ywCBG4YoCPXfauRKg49gDRTi7ZbfIf0SxPEuxoQIvCegqhARKSvVtnRQ
DGN3LTqM4V0C5dcCvad290aMbLSaXX1COjG54mfeQp0h4JwrY5m5mn8Z66iqmu8h
E8lRq3QCcbPjfsVWrOepo/So1sl6qUTxMKcC8yhFMFBes8GchKCtmzaTUKJdaKRH
dfQ5bGf5Vh+R/H2h1RYNx+EY//SZlgqS5TV4HD/ZQY0EXhzmg9HiZvzwHIhPmyc4
kjOWEmj4ihvYPsDZP5Ojm4LhkuF9IAVwi9zG/tUq6Aiss6cdEn8gKXMhaR4IJx2g
L/77GfhAee6mCOsWj+UVbCHn+0OMAZns5L00ZvWq8CH7m4YzCWnuipweDs8qqLbi
eDTRXd0LgmZbJ2KVTxRSRl3IN6e69OCnA1DcK14TIbqLeaUfXgNEshjxrigjFIGd
v9mPqCBGVh0EUPc7HAhBaiW7J3oOS9mmnh6Vml2oDmHmwwxNlZjCp3ypptpp4McK
31benvnnQLdXRwv5DN8wvqW8tQXHTcLXGNzAfLiDQuYN5dp7gGHbgJc4dLCo6wpo
YmvXWK/9vi17L1uLXlCFTYrJyi8FD4FkfCSVvRKfjUWBoXAhBr8JcU3Yg/LYmGoR
hSIyo/NAkxWYpaNL7LQpF707Y8Xm1oFPwPoVfDP0+F3Cb7gbpwA54MQ/a/67cWVN
edG/M6V8sVtfjTQJmu1n6EHWSWQGlSCS0JzQWj/5GrVs7+5yz8RDnkhCP1aDHEoE
y76qvo/Lh5fvgXQKogIhmPLb0xoVHabjMlQSVbGUNFjpKZNsv+sd8UGCzk1IF3fp
fo3t90fOcmSsDJz245XDx0QVYbUZlEF+7zWlGa1NFsU5pkEqp8J62RkCz8rOcPEe
bZxUj6+gTXEINCfYa5tr89evQNU3DNY658Kagj6DlM6IyXJoVUD+kWTW0yUV/yxy
B3Tx+M/PU70HgHCE/w1SN936ibaYVhBTB0VZB1Cq+a36/NZii0AzCqW+8824k8mT
0mHYmDl9dSdjDX9pJMqnOkFY6WCBsn42Jkj7jmzOpWzTf0KGw/m2X5ifkldlOtqR
EE7m+bFrYXM7UTx/emKkWKJ53K1NlNmXD4ajvFqTOb6U4PyDJQZGGGiv0x5r8NNX
RZpHN4wRfspR1m7tQgPrnpBjSpRb4GLJRr93cv5e5kkdy5ZegMWnuZJGiFqABhHT
0ohViGtGnSGOp7CePqLJdNCGIUC7aDjR2e4q8eVzU6DwgaL/P5G9jGOoWTnpHlp2
rIAKHW3xtjhCrkwmRK/qR+d3jFiO5m5sykcCrCrCAO9xILl2q8TC6h1b7gB1GkMW
8fQJyGKmqZrtLyMsrAEYmZlYjsTtNuMrw3syXWIZaFfzYnudNRYHAU8Ww5LuhAcL
aMS0MyyV5+mf4ybGaPzrJoo+2Stt6j8GnXPqnAEaUGLTFeWAsIJ4HDqg807obsEC
dFZP72GSHDFc1f0Zk3eq+ne8JeYoTLNbNCqIloUcQcR4LUhNWVf/C2wgOzd8ycxN
ubw5fk0MQn39W1Icsfh6Nf9HUGXPtaugXedGCN7beUDIlgu2mrZK+pFrolkb2nGf
9PZB8aJ7boXCAunMQMy+LIm+jAS7dpuQ/FVokVPIP8VPoU2EB4ED00pC0heg2eZI
NXrJyWRP7LaWgyxtyKy6Ym6sg44kTcn3mh2rpVAE45v2vPb/LKYlIYHqcLnn3X5N
SstEQJ6x4H6ludmB3bV5NEvOSyj66Qx5QYjAgaOSXQsz92SImL+x8frS61C2R0ZG
sw8HJ17dLYhObFSCGYbUUD4c6KzPHyjTnQAm/ru6ubtgmV1IiK/WKCzFaZkXEuFE
9JViShE2giH83/cNmFZSYnc84/fDPWqTAgBZ965/rEUhgzc1hf202Jc9fOmFkH5f
/e0lQfh1ludkbu3hC/hS8DffYhJE3P+7eUJpFFaASJyW4wnVCv2sar6mEq0n4GRv
uK4OBQwHA/kFkuj8WMZbQj+HVrXzNhy/GCzYv00PILgnI3mbg/e1jxYtOui+L4Qf
pYyyDEMefaIYkt06yXreU7XhV4AgBXIAbRpGwT3jPJEvSg9KsNHj+dR59euQrzp2
MmMEi4ENxZrOjhX0B39h9lrAJeim8rwVjmFdVy/9TiKYmGBqtwqYyHS0DXDabzub
ciRta6SuOzg8E+rm6MxERVEWtkq0YGH03p8NxQMqQ1rVipaewZQHn+8dGbFmFdo6
QKjN8V4sbxiopuEtNasqcbFGPjNgTWZa2iqQ5f5Htibt0qbWIIxZG1g5fnDHhQ4i
3lEzigatOTsXbU13WCWorCzreWgwXVEPKeXeQeWwD9ktIl7Bsm0A50+2FgoWeDyr
4gbVAmshAEsJIBlC9pB12Spy0i2mIO6ov4Vu5BYmLHH1HgN6c6gA3PZth9UYXKBE
5j55lGCoHzplEf88T+ju8EJv+9RIZDnKrgbrK/i6c27zRR9KpRL+nCAV9blF/aMB
9vGIuWjmkPQ7McKj5cff1/7Kq8AhJGJFwnwAh4nRREd/PMGKPbRy8LPS4FeqguMN
9ZkBNafjlFx3YFJ7r6L6A/SBspd3TFdpCPAGsaaZcvnyXLFZcbjroXjWQ9F1G+V6
+FU+JUhkeFTudnb8lYb6F5cF+wRfxw93oyHLtitXH9PRDmVLUZFBWxVcziq45GEh
gG7TpgVXfxdGPSQ4wr2UxdtaQ7DEGaGx2sjal4G5+NGr0QDY70gRAutSk/2kihiV
c75viipM52jNUmlw+WCYZVb+b0Ia6eLz1KiXUAMiSNonGrYNfy8icWtjKF3tQu61
TDbnzJ12hex6O3mPGKdHVTuJxA6+Ac/lFsEJEnEGZavZXVf283hEujXYlbVH95z0
jcUJ7T+Q5AttZ2KP+vVsTB9GPJrwUROSJSurOuIcYfSJ1WrjQwNqig4JxT+YMN+u
rF83Q2A0+bnpTg+di3fZmwiuInzpFFZZHGNWycXIHKw4x/JFu713RZ7lDK1J69iW
OYu66bAmiAwf9pOJcSf7DUZvfe6waEk8UJPx7Djg4dcVKFpdNpBZGopjNrVhf/xm
IbwCO/XyW+CfhzXnvIPZgvZa92Knp28LGLb9uQ3nW/9MGPe2Oo1Pp2KhUsCOjH6t
Qh71KrA+MU5HLPchEcSzyNrPmByXJbM/JJFzNFvYj2x2VbEPAi+CWNao0vMfUsu3
bIZwu71PYBX/r7dSDy4dhuiUA2aK9Heq5pUSz5ofNVorxzKiTw6JiQN/hwC+Oetz
/k3xUu08KlIRTI0ibQaI52Ft6Js87JfZHuH7m4SsGHucRI0B05d/slOq40PGGcnr
JXwWcAqbH1o6lkpqdtwsJXFRATrOt3tJr6ATV6KJmUGXaxCuTmucyMBQP+54Y6lG
KmOfmvj4iSs6x7UatlghsfzGGf1Fs1i00Ss6DiSgKyF0kC4Awfuo9OcavfIILMkJ
f5toiZXeancBK7Gk8i2BpUZfmGBDitdHwE85EfOioWgK3zMjcb8+LN+tBjo8aV2X
SE+4+7jqkxdFdwlM2kTfAtN7KcTviifm6fb7iN+KOmi/75ocH4cEVCgJLmegIcGN
OgvhKgW408G2TOsA4ec+sLs++258tK4z3P4q99etmazvWPzBKteBEIvj0yFjW+PE
+Lcek0l0KwNBHIGaRGa5NyB0d1GwhA0Ffkq9OiqYXeo8cH76YLtcLW9bLMlc1egM
IvF8SJLvIOVnYcFW5To95GRiDLG6PTgejh4aQe5ug3mdQFN0+FlJpmZKuL6bUwOh
Dfl7I3ASjR4q9c/0LXt3aJoc123jg2/TcJ7Z3zoGekiIH6TZ2ulKcoDJILiekKsx
CtEXm2jP5eY3pwK6UlIuZzhKSVkZsnp9ZsbCToKpiUYBEiA1GOXi7r3b5zaz0BrF
ubRA0246vZjwdbEo8t6lk/K1+ptoX+RXq2lfQKlyRTuJeijpSb2ajUSJbAvbNqlM
5cwlDVvlxmHHwMjNv2cw6LAoMJh53sB/vEWat6bspbWRzWITRwIRpkpnyrQVc391
vN4sqSdaovyahd2G8PTxvNIV5WGciQTmIwIFNP/8gjCnErMuX2cT1txvWXn6Fntp
8bZE3jNzib16uZthKh4XAgbYwjVeyxOgTFpqQO8a6CxJrcrRvP2f+UjgBfsvXPEw
zoLNgkgM5MYm/VLxuHVpHEjmx2si2U74kOSTsGto0FgIVUatruWyF0Fnr5LbB9FL
hUJovQHtKVDGyFMJe4iRWNOflUf9IRcIuK4Q4lAk+rDlSnLqJnVQ5ZFg2flmvp+Z
v/BwXG+13kLCztLWFdqljPLRGS4dNEUWAUIYodr4hRxnCtA5n0L+EwKsQ+Lc9Cgg
2w19Sff81y4C1YIVTLk61RX+by5WPTffxtIe1OdHtCUssRAkxvi4ToGZ2Vqrpmez
MJGZPjIwZI3yUgEzfMSa/eLFALwX36w4nz3whYMT4+X8uuFIBWfpkJjq9KNdmtO9
pvG8mRe1Rx/5I5YPi++0wZ1QOAKQRvFlp0iwkh7kKOBbTiESx8GqjRYfQsDb0Wqc
4c6ftmK/l9LgyKWkd/drCk6IywbMlZmq9Oh03PmWRCfbwWaQRivKZXr44ESW9tkG
DgZfbXxW4Tu5lyaHC6FS8AJgmcdSJxZr+Fvf3gyRj+6fsckTym0T94Ic7Q7hKseg
q/yxxafxczmMS7HXciAvVjB1S1R2rB9VYk903nlLuFBybvmYN6lkuX0A2d1SOFif
ms8Wn5SCEXDVXR3qOSInUIvc5KCxIl/2npjPW6xPLtGd0pAcmGfDHKTHW52rs/59
3kKkjdR0I94TsTkFQhKEpLzOQyy6zw7lnOCtL6nerzNn0StxMLsQAG/6JIq9bJ3/
FyFMH2Z9NC5aYc8qr0CZ6lx/uBzT4E/5g/tQeTO4wRS3BoqmB4Dzfh+NbaNQSqdD
BMOm2tN9GJeX/MZyV6xyySwF42/D52JrWgY+R9ippgLhuGwNVVDLzDKxDOnz8mjP
t6GlLFsJkJ+xjDOXioOSL48DdS6VApDuUd6aypvvnL1iqKJiBD7T4DiIiRNLUc5y
N27JlOkCSfyfYuSW7s+8fBOoRcfhZLvHyaszvxQ0QwBlu6xAwFXY5AI2MW8LiL6z
ivOeWNSBkh+BfBy4Bubm12Z4NzT0RwIc0Qgtk/JmH6Cat5cJpSJs+o578QF3ZSuh
1bZqacEKVOoZSa1fUwF/pSJDHdjyWsQ7ej1LqFZ1/Z1iWjaR5Qu83CLmPUF/IOW/
94gDABW0z8xzZDAMupNSSex1qqQXPy5uZLFdoxHhMKz0yWS/8q9HOCSzCf8Ahe5J
bON4mCpaqeXrLOMVwUWiCtzNToP3ExMIvo4Ex2LMP7zFZf5OTBE5nM9FAMUou1AQ
uYJ7BUG8dWXmNh+eocfCg7Tm6XrI7NTmMyltcPvm0LDMQHJOXHkI0Jq8Hhzm3Wvc
v37wPf9cPXCaF9vxp6SpfLIB+9eOwRNLFVS6YfCy341FzSath2uX/VaYpE3liz14
wd1s9ARS9H4H2HtUuEkODjF6noDmmOTYCJmOOOz36k4TEMCoeJACllTIKBkJ56fF
ebZZRoB6UNxcixKxkDjA141xuNXO1twEdZqDuWF3I0bGiY0q52jOzf973QkwY2DK
2/AaA4y/BtlVZUbA+31iTRH9ypvhDkARnOqBeMM9sZ9aQHQLyXguC+2EFE4OROAo
BEinmYPfB+WTpE38+s2Mjj1sEIH14HdLmS9G8HIj1RPeL8zzMstrTQ+xAdZ/KWEX
KkrrGyZ/ZW86MZt1qVsbiDn1dkSEOA14TQt0sA44r/QQbkzhXEy3Kn7wfgDhj13A
e8ZuzW37fKAdYu2fDrfasqCT3qvOXmWn+Q6YSUFYVoixI7KkvmMGN5bZkOaw8itO
Yqt2yZTRdEez72iVw0a/XtmDYMEcgxWEz5jggZZ++ixyzyArC4ee+8WhZSoB8WjC
s/2K2Ii7dh2JPf10mNpLZik0VuxrBGhmvq1+18w1BjE7zlFlQvC2OOd2/uNWSWpc
hk6kBBFn8bhk7ZQDi6qDIJ71IojkgPXk71q520itLKKo5oV2Etu5MFyY4Gj2Mhix
4yW7uxnQfdnUQUicbjqEoNnpCdLdcjseI01RSeJ52Iso54RIbuqg4CFT6JoLJUET
pD5scnFUOQhjBWMkTQHuF4LcW/tThfoCOtH47S/dDEB+Tm9KNkEFeljeo2MQhkYX
TvgYkhEVMRECoXHqtwzNTFlC4SAwxJm2HhZbDlNbVWNzh9QtfaYo0Hyx62VTR1xl
6w+G8VMUyIptGOSOIedA75FxzQGA8TgS5BmTTjSrAA6nkjSzin2BSANGSXwRa5QJ
GKO+EWxbOYVAJMff/aBpoJM0Tiqbfqacwv13l3fPAcQ05FfXj4eMzJZeKkUvENHC
Ik+/Hp2i11UPmDsUilkuF7mwcrPudNYvxaPSRVm87KIcr8xBEfKZsh5QL2y+iLPe
xIGDVdnK1S4AAft6rbxvikxX8aBh5jxTdBgtaQaWTWHkue8hFUZ+U3XqgKJWGgfR
6RS0nOgqSZj9tcrQXGTeG6WubXQai+Jc+vnuCiweFGHTN5nBe9XSXXdNCQSGBjcG
IVT7yrqCRIftNVWmf0gcYodNyKl4Hcpd8YVWCi6OI0XW/21qJN8QNa5ed6QNqIL3
/dH7cZOcVcpDuQowjFn+gQjqWrRCRxTRco28Cqu2+h53g70Gl9uB6Ib45gSW8658
ax5u/ftB8bpDeROQukyY6AcjjGOED5D47pUqTiLrIQSl6QII71z/L7c4Kip5P8Qz
8Ghh8G17bpUulaQoDfozaUH9oUZsfOlQkmax8+mXAHUsfrQ8vE/6aHo5akiqoi5O
yQKKDS3VwwUiUKTLNYM/YHb0qn5ytGeIvQmiNn2+W6FJDJAA2J2EmcLTBz0ElJ5k
PmD+Dfw6NvacBsFuo4LDz1h5krZz8CC07jwJQEUBSwZ5pdqwNHtpmE9M6M55YUQd
O4uJPCSu5mepYO6wR7C5oNgozsSIaJgvaijX6KO6zfOtm3Tjc5OK6ycaA2Pp98us
oKpvmK456FKBAzrJTWt1Q3ljduUMvW05+lycT2NRQOZ9srJBP+XXSVnT4YjHKCUk
GcnF2yW/uYUUkbLHnym+L2W9opE7EPolkFi2eCkn5weRqTHYu8JUnLnXyjknyrYq
+l8gcm5biYIvJVojBHF9aYX7Gb54fluPFQTOe/L1Ai9eUKzD6zzUFZbyS+hT1OQ6
isqeJZdba7dEIX/AECJ44XwLQc5rJrnHb/RqB2Ija3uapzDaN2c6gZ44zKj6lUJt
otSy+wNyA2lON898yc84FmDLCk4uDBrMBKLn5h/QLbgn8E0XteDQLUnPhq9T1Tw4
CiIR+v0ClNz+B3AeH9OpRz/lgwUvnVERf0vGMcsyxAFIlAWvlkfg9O4MEO63lslv
0KlZVyK4+hFKuMKcIk6SX2vj+Xd3xBwrj1XcFCXsbAPgYa0MvSjBiYSALWhoPCuL
QS90jNY/9NAzoRimiIKZfq1HCi/o4nkDEmDLqku4AFtXNmw1MA+pHZoAI6++30rC
oTRwmkmBJjt8gvaYJ7ipazpRW8M7+0E0B0X65/QjCBylCCTzT/6p2gddBsolTmrs
RZgJa/9zvJ5OtcHCceNO7lx9E7cFTNOnkXBKwDCqflOxS5bIHbrFM7E6rsli4uR/
Pg2IYhf11Z2Tdturhto38rM0mUVSlApV4RvghCy6mFftv5cfdVx/muZfDEhHXTPt
auK0BOQnXGSG2bfWT0S5osDs8nDvEoDjqk8v8E7C/rBnfxVXikayaBGiAeqzJlcj
fdsnXhu9yMXAe3L5ExSKIeHc0HVwlwKwp1vY+RAheK5mluSLNomr2MOSgm/8Lb2k
cm+y9eM70FlEn+598iv6prAOzgDiUFyJNuce14XpFtSqMWBrddmXZuPJlP/+iGBH
D9T+cG0Vsc8ejiJo64tw/2aYiwiz4fPeiggr/kyp66+jHcf4oFuBBikHTgAKKiH7
xGsSXvzBV8XeYLkxJLSbPj4xY2bRTqJimGKaYXqMF6iz/M1BZc6AbHXSGUNpX8lN
uVNHWr12xL6u2ykuAyUgs8xtSVcPIWO3K3XoB3kmwC01EXjOcr7BvvrLjMnQv3IS
RTz9DqHjqs7vlrwCXK9He0s3mbC/v2Iz1ovd/lIIJiaXqG830VupSOSVp2Xtq044
ksyeiIivsyGJKUr/mWWkJLmSXMCJvteTkG7El9GrbKltwfqpZicrfHwt4eNOvZg6
6oGhaeL6yq6ms3DvrFL25Kv/oPi83s+peOlzlIa9g6vOuW4WiNHCYYXLRFnTyhGg
agBcoeURL1ZhbiGrEpJCD7bRevCfw0XBZaQ6xPEW16drc5hI/XsrXtJlu/eHOd2v
D1k35vvQMPJFziPwRWHlRMUjF6VI4HZDepl11i0F/Skw6YZxasrh9F6vHvKRCLOp
lPJx7v0xINiTs6U+jpvb46WPTFe+TBmqB1jSGndqavrZRx42PlZ4W0pzA4neZZhN
FxHmguS7rdUgQHWJdrlDXDCdFNsd/jhKv2Px4VYI7GS7oP+tBkN/+vkG04e0r2u0
ZSxKwpQdD3YsZ19HiPrStsddvKaMdyrVQel3qdqDJlMnO3wHjnvt8vLZJhejm6hC
oaEqRAobKwL9d3dLOCZ3wt2ghB4P/DNZ51Bn00/4QYYwlIud1S3+mCqfpHncXHLE
ySTAvGWI2z4dhgxjZMJkM8DhcdwFT21LXfrmv31WHNcFzZlN86z1avR/LVKp4JHG
CBg2nvwGUQv8OqkpRbGt5gPvMMgH2LWLA362xQt8Img2wZKLI6m99S27iVkIUnlE
5MltM0y5t/0HZhiAEgValxkx00EntBQm7A03rBV2omqYNqQomxbRtdHyU3MdrKR4
V4DNyOcZHUjAdlW4j7wqSlzgCqvvghRgXXq/2TmECNGj6VltJ2GQxZdNL7mYns/L
xPXp5qJrjNLVKQexCpFAQ2fbJnbeWUvWqehBua37bl/CW9W5zdesYt26WYCoQxlz
96kjGl/6PFB6a8TE7E0tPy7W76GkS0BGYSX1vhhwrt3YX8Oiho3Re6YYTMdv8osC
NUkCC0HiSxmoiHZSTAfUY94jodiyYz9pY3PaQ+agV0kiVWZDMtCAiQPlNHpa5qeM
feF/mRKRlfQKeYoG0PAE69hChQrAHwSbReSmaR544Z3iTLCjxB3D4ByAs3BEYLVc
EfEf+LwQ6dNxQ3P/3C7s6UZMwjs6XdTVP7CM6Nu51yXdBHjjapVNPRZgPLKlrpKJ
LNIHtRryWKyK0WuV/qluFBKNkEpEv78WYVXtfOino+msbGjgegTAkEzpntj9f+2/
lnDmpiBuSaZJiDlLNPSJD0VXpEnxuQpWojBYbMb1nmyeCcvQ9neopu9oC4VUlYdG
wqzgvv1Da8DF3KMF+ZlhqwgDnpPkDKUbb8wjw7BN/NmYOi1ngR75OMAFCjFfdpHF
F8qvJr+rbkWJF1iZD8/GQKgaBYlwiOtCwpsaGfSjPKXUay6cDiPrWotQcRvbu7XJ
lmo/doTZ6CPSuGNGbLaFv02JCVeP3Vuo/ehKCMNpwWHXgQVMjmra5lmfFi6pUeVc
N8KDI13tRCEdIpfXArpEwLM32E5HqRqGcZVhinSgQY+LWp5oF8Te+/LZC14MpleF
e2J27DeCWqtQqSsMLYV0eX/Z46QAnb/SQvUq4+bQPo9crE2YbnHvOl4iiUluQpgR
vzvc0dFuyQ9xtPAv2P1dleyhwRqnwfhdGwkL7q2dWGnKthgsUJy9eDtaTgQFd8cO
USxSLWaKTKBqSygP3dwU943tYB2HC2Aw+vXmLzb83skqI5t1RZAmej9foOv2Vk0T
Z8/tRY+SfORlvhkVfF36hymEuHkAJKTLpHZYt6CksdNHjiW2elAUsUmvORsghvOH
vuJbRzKy0bpIgR38uLKx3soWhIY03F1t+VgS2XZCZEpIU+n+r16z2Q02LOXcfDYK
y9OI4yCcKT7HVaM8zcBmR6O7JEJ4gOvi4kg761viJ6ZFaTk0avbJWqWfOBmDEe58
YaK2LOaXbqrqr3oN5RusAFHghE39IwHUZkVDEEMwW/HeyJXZUyUTOSXgX2Q3M42d
zmsEAMe2VaXhK0Kj7Nuo3oFJze0xhokJMq3HoHFUrxQS3KqUbjmGNu+Bd/RORgYK
3eB4BZvkRjnYyyhoz5nGg55Yptor8cpiyuvwGyiNp0Pa5Y6ezuEnraxKjkBwOs7x
7NhpaqTjSnEQGZ/Pj7TWokN8zekfmvyvFiZgchi6djkdy7nGGGWICTXCJChrF2Kb
Ugxaz5yTY/PkffDDNEqn9Jguc7d+Ad64uFpKbHs6kh9i2TcdaMEUGnt+3IYzM6rc
OODUlCsC5jp7Bh0fl95jXtIzX+incKejTnCpxRXWDMS/rYP1cREib64mLiLyHbeZ
Cyoo01C00EWd3wDEfA6Xa6cA3XH0glPZt0bRVma5CnzEU+rc0XHhEHgHJgDmvnAE
OW3J7roo6A5WyXALHtkMwu5xPNKn2GGoukhdYbpVC59wj2mJDil9r4rFPrvRRxex
5+aZVrjenpAzYb3umJqedyfBAxxF4a+HntIC6hKUKSdhIotpC5fADcNmZYC0TIV4
sADKPMgn3mW0bkcsdFTvx7DpQex2LPyGJieagvGGtTqgCXzpo63KelqwAXJe7/a+
6+9+Jh5xxYvS9DasOEOf5MkTnHg4qieX2+ecYPe6pmgNXkxQVMqTuWZcREfFS/cu
eRCJJDWgzglucfNRiQcymImsjs7KX4Q1hVHc4A3Bv8CcPfjqNTbVwWqc4ZYOI1EY
o2EFqGY4pqIgOPJgRKr4ZndhNTKPwiSawAbRDEGPF4GA0GMh+V2QhVasLhefsUm5
g9hqs/HdAqcsqrdZ/fi/RNLm9+LzypgOivjl4cGF/X08DlSG2YqIJrbHskUhuY4j
ZmRpSddi4q2JYN1RRbHAI7XcGsDa79UhqQ8mYKBtQN0RVrzsi5LVMYzqnSKSLwWl
DMRik6pEolXdSdcIbCE+HYafDSCXd9ZXa/CsQh4ZLH2krD0a5Kl2tP0kc80sWxZg
HSPp6dO2qW2D0rIZ/RQkqTpSGh8JTslC6+5sZxQtPuJgaGMYrp1+l1SnwXB+RwiA
eoEL6ZFp9rGThaPRgatEjDD/Nyd5aJhvFU1xrXm4c+B7dpQx/JIGgXWW+iTTDLt7
LOg3dYiSHA//Q3CRA9EkY0yR/bervL6mbEkLjpK78GqM5vvxJocBcRiS/GGdFs8z
NhIvjrUAXov4L08RHF+HGvt0XUlxOgIAnuwimh5kQdeIr+UB906FUvBxSiyWj6wA
v8xHXpK+Q2dEMVWTEptdoOquScZcnrUrnlxizo/cFR2mEf/DfIp+m/MD7WBXg8+3
lsmX9FLfhF2KFfaV9MuoMUTx5/i9CCibY2zSu0GMaX0EBX0OcMtdNG42aWQDcmVJ
hbVcbH12FB8cmW+ENBQbHvMRqWjghhsGhLhEZz+Gis2q09gGyH0efg0eAbhi1G9w
mPAllgslHCrpVXTUcSQ4AxzWQepd9bww6qK9YWvLF0Q+6jL9s4Ue/H7L8zljXLm/
jOikwjSEivWIDdYAfzifcLKXLz87ZzBHv8/EH4k4jXseFQgLoQ6sPnW09uEn0CY4
mhchcjJ7JjlwBHe14nKD/zX0H32BJX3PdZuihPQ46rOKOeyPNP/A8lnAYwYAIBed
qtV6GFUJhpuFRgCKCDxKGhfwO5cf5y6PZt71BuNaPMKeFalrYrH5usuh35WM3/LL
oW6JYXCGi6Xbr8hn27X2KfCDRb3SN3DhqgiamV61xBoh/N+SWkAnlfXobrHnPBT2
XnVUWpwjqxO/OT1XB6M+ZN1S5VY1+3qjFLT9hlvwaCNh5vIMD8ordXadoYDgc80A
/0XFD5x7bPKr1vf1rataoq5U69eDApPsvnQsVGYs9PjjCuibXWFRJjFNVJ5vQluX
07B9UojEa85ZNZzcaBMJUfCk9q0Gmp/grtBagHYirpqRzPNjjJO2MwY+Koon9O7X
nTKgBYjHbybl8/TMXudxfC9Rj6YiTb5w1UArHc9Xh7LTL7+4UgSudeG1t1im2Pqz
3TpgqrEz714yo+1he24lsuCdywAu5MS02+72Csht7In0Wj45oQHCdqKhpb7y8erg
P6r23yCbEHjpv+OTewB9xmy7rCRL6xL0uX0Lv2caQ6Bv3PhF3klnckcWq4HfpKSn
eed4pXvS7majbeqydG10XPdx9ejYzkCSONWzSNF4Uc5Jsbz/TsIWmi6zExEkKp2z
g3spBHQHbrKJYxCtYHpNRwmqiUjV9eJej//UKHvJ/d80M1gMdLwwTEobTkXe8LZ6
X8YnCu5sgdVbQQv1MZ9iJElAkGxiwB8metI1weyPTDQzuUFTeBNpJqx5rKzc6wws
rVKOoNq/9ahaEQ6dGFTCJDOwTgKi7DEMU0k6NsVs4kkqeWkma4QOAvkFVU0H7cpf
a88/7Oj5U/qV3bvvinjx98oJa28XJrZuxpGfq6JJbu94zwSd3qvDYacc1KmxAIoI
nPpoxt2PEARS2fbgNY4p0KmKOVkK5fbzfte/Y9LtbqJnES8ZSXCfWt8MDdivSPWi
achwDKfAnAZoY+CHc7OLX1b/1JDov7y8UpFvUTpxrV146razoXTv0YI1ZJ17pTl1
6lmpWef5YFfmzJ2imn6E4vOqRLaVqQtHd6jUPgN21Q4vUwGZd1sY4owqc8OH1qje
+ntr9Cm+x2nmtLKFiQkzWMXkqTq2dGcsq1LB5H0PIZP5CxDYfKtm/HV6U3rhpMPZ
5uaKzyveY9kvgNK9uS0cx9F6olci3gt6m40vqQsMMnxytC/7OpBrBf1hDrQuIWh+
bbgqppK0/K9Isv51OfnfzaoD84rioCHl4LeKdv+THJT7wxpMxDOrguJoaA2xy4jn
Vd2zAQSvh+hQXsxi68rbVRrvUwPq6XopWOZn074VxUazn+fPEWj8klrk0XAQbgF7
LGahRdBQ8SeV+K5ghoywB9/YKsTf12LF6zjAy45Ly+WPUL/gg4mvrUaX9T809+mH
9xirQO4D5bx+YR+IeSOYZRBFmOZmtcKR2YTXwLKuI0F+xYzkFOfjleOA0GeuqyFR
J/6v4A+Odb4vJEkDMgfDMtfwTD+P+kJa6EbRLSYOA6hjIf63kVSeXWzCYQx9DshK
4C+h5IxFevc/sN3RPUmTvCRgoo5jIFobknx0AMPeaKyL+Bc5Ix1qsH0/D4DG3Xlt
VFo06cL55IU8wVfIRA54xv5P3Jrhz1gw6wHo1+cW26aRDyqXCXXrJYu1n8wSeS3Q
v0Ma1KYxrIExn76PyWHDCkMVchXpQrpVGFSo4F9ynvMYtbwfHC77LDriI7Z0zWhS
qZ5IHO5eQgjM2Xz2ZXH669zem/v1w74Z+X9kD8qgHvJnjeaCQrDdgRrqhV1rdFzI
Oe72wKu41VaZJvF2ZlksKZ0BbNDpRzMQG5nB5Y/pUWn98QdiHOnEMsEHMU0+8ht9
3s5PHPXZM2zu0g+wMDtQvbyo4TD8GtnOGo/jke5sKBEMMX0BaRJkoxKS3FP19iRB
yZWj5aPlw6gLflW2ozZsuBIBt787Bvfzc+VlwPYiY8bqjHMhiRK/ov1yEhj97rZP
Pb6LrADfgDJbvkvAPJzVHVBmwajM9b8SKZUSh+IpqtlUJ8Gg1BmhtM40HbVJpKGW
QUYhJ/h10Yman0+yuRn7394LzO8BnJV5ZtYHihM2YgACPaleYXznC5seRLhf4Rfh
dJPKQ1vGLWKRmHzioaZO0qoX9mO5+MHEo5cNx7nYjGeabDaU4e6u+TPltDdszfFY
OCEIeKnHiUaGF/csZTaE7d/qJZyyeBZmIVLlxcg7hmwyeutMz73qmIZzKYOg9J6+
lYrvnZryuWbjQ3kGerfVrVPDQV8hIv4L7STce9a9SwwbmlE7tnWZB228EK56RqyU
m9eXKey5JhD92ZqGLDUIP1EB5hLvXjtKz+aA9jOj93aVcKzv/SWLZY8msr7hv2XP
okpk29gqOxnALSvAmjDQi8bQCbWjiyfEdI5d0ilSAI2t3dm+m7j+paNp5JRQYJXO
Oyq3GI4rIp+5JXpTNTV9wPjraCcDe0SakmLxjM6tBrnYPzQHeVp7m+m4Kx0rWP+r
HdncTa5c6VWrekOh6/o1Vl0PZAdBv7NHFFuv631bKagq2GG09QtS1opivNZXWCsj
aVvNC7ZD/xb/dPUzvt8Q7FoL/JUD59362401mXw4QOOqZAOwytubYSJPzyLBtVpp
bg+ROowSrPiCTohMLLf97/gIfE5nujWA26KVvQYYsT/xvekbTD+swuV3ILM2PYj+
gemy5zzMUbK8NTjNQlx3qGM2fT3cfN2JpRoEJLrWKSok0UgtTZHbTuMYY4BSp8aS
ovr4pEnsmlsBJskRpbDsjQXB5LOgQ863BCXM5SFjENQkbfAy/kMif/qsOQkUw+Qi
8zb0ZLopkSD4/qVFe1pcQ0Zi/6J+FiMFv/+BEuj6yitSxYzZq5vcoWCBnBWsH8/Q
xArs9nk29opmxDS6XW4GV52ih3iXA+OrullqAcNdwwvaqEYRtlWdclmxkpk+pEVP
SifVxYEZ/l5LODLs0lsMBb7KwcDi3ss/E0+ToSTUus1EiGcIG1k9hQ43iF2+6HJy
N8wwHL/KH2HnECuHb8orUvrfvUBC8eo7tTsHfS5ZaaBMAc81B+eeuR+PjSXbeETv
lDhBlL5bw6sFi/a313uAOTJAZgPQIqZNnZDcohSa2bjKo3No7Ki+aVqdrlXDT38m
Wk24y0hZ8R5JVsUGJtRb2XU0owLm6IMMu6SBLoeAqVyoOtpSMQufeC/BddETIxcG
PCN97ZVI4slkU3acc414dqYPg/BhVtN+6hcifxJ+wlFVViY2hv1L+mSSF9ez+uVn
CaaxnE6DoRbSpv8HkTgGpPD/DQQk/Js9Ge3hfY6CD/jELdH8nZw1jWKv4jYsDCYS
ZkRsOpeR5Fjusx9C3cjmRtfF0dwmNcT/NqPNjpADfyjyaj8/kYC1CoIJcRUVHqAv
p2d24c+e5tMaUVGC5Kd+W5mNwvsl3QGVxdJHJYi01bR33fEC7Ipi8WVP0elQ2uBp
EnTffkJbBb/IbLi5DePKPywB44+fZg9wdQ9ABI6XJcD4W5adhE3IXlccTFLXuptv
xBTd9rYsxEnawKVY5KF6msGXBWdovsYSMi9QXCIpeSCqSgUFlH9c2bFNQBUfh2zW
szEBS059TwdrlPn2eNj9+Y6yeF/1YuhWUifrpAAAYTy2LxaqXgylk7ipiTaWfHhf
VZZvlZbBjLBSJa4WpuAdSaPwKt5/XcYxo//f7uudjcFcyHDDb8cXigk8cAde4YHR
zDewd8OOXWsExVHqIxTyKHVbgS57YrJ1eVcSzUjSC0cwBHOiDmV9rZqRxDzS2UgC
JP0+vDOj+zZQcoGy8AS/MWoMzjNb3ss4EpNTz0Zv7Kq4hJd0uT18x26/rTNc56Cc
heAsj8Yp7BJM+YUw0VbIQNe5UZ3HcTMRhUBmlKPDa0UjaFkYorqCX3iyzl22Q3+C
VKVPokciiqGUVpP1xNgqLn1HXA3b1JEXGHDStmahOWK1CZZUisD4uPecGVz4Fs28
eocRgL5c3ON7DSEI7qwMaodvDj46Bd9BtTtDJ/Z9u/V1BH65yUDr3wVs4YfC9NP5
/41DnH7SwdngAdiAsL5WE+YmJKx56Ecf2zvWEFmV4IB9Yted3WR8AOVtDKbjp0Vb
7ISYdElrW++OH8q6dbkJk3PY1fvyGua5vm4s9LJdlzSHhop6UYO0hTxeDLBzKl9T
x2u0JBiAUrUWsBw8ALjuua6fDtsFp59Nxe2dJL+IebHCtq6bmQ6JsgxlL0CbDZYU
qwmY1PXfyzeGsCqHI+bszudfZC2fsbMW2BRofJo0DVEPAbG7JAHPcBvLFmPTAXQD
m8bIKCkWphZ1Qca47fSGh/CvrUSny2sUDEe/x639hMSBptVm1DBm0w3Np4xUVwux
Ofg/qfMVTH+oQqI/CbCnDHVnXB3h0Zq4FW+Xrv4mvVIfbTtI7z/uygQ4z8ng5oAf
HAxveeOvrKFfcUkp6tK92N9L+qC8lBMOZzqIiWCjKzVUKotBOIYzif0b1rujK/f7
WeJuM0cBxKYZJQV7StUqG4qZejDi7MgcFUlUyhUqCiXJ2yCDVVrPVTJs075E9Hjg
Gow5CP48nRWJQg5fzYsLIBFoCIzdSgM5x64+xcJVrPbiLCKDRbTDsvrRN30jBlEW
kTTQVaQtDo9ItJnyr4LiXmawLt/PCDaiMROtDxGahKmfdwcOsn3WVFJ4isAQ5MTO
7Pid1wWSA+kEtESvrK8YTKCIRlrqSCxfvhJFIh9JNHkDD6XPj+N0zKY/13iIYeiN
bxcWW1J8zxeNG/SywjWcHMf4wmwTAwv7prrnL/xas9v2XubZMXbMMp7lQ2/hpya4
wLWQmtBIKIi5h/j07XGZVcUfBzzsYKI4rEqKvS3Ofo0Ph47OHunM9hqBhPb54ym7
F0IavQQ1vRllJwSCrlsgxqIl+s+PDZMnPDGfjiqYYh6kHW9yFpDCiZ82J2/fYzKH
dYL2Zg/pHoSQV0h3lCH7F9E2hmCUYbD2Jkz6L8zvdwavd63glUcji45SSDMDWnHf
Kyf8SWxvFnr5Kwx18j8MdcM5IYufTyOLw3CBpsOiLQufSfvtyrvh8EL50GBXl00U
i+Ox+zROXw+RkeaK2wTj6eXEc2dyOVWqPS1SBrjhYjzLICd1sq6fe/JpkH9DsA6H
N+lu2iyog/8ze6VvB8JjTqUaqE/+us+Ynt+iGBjCEoaIIpQ5JVir8p04pUHzzqfE
0SGSiptuCoNAWycJ0fG/ZxpLGMh/btRW+6qvlkesuAvig/RRvbiXunpYP60N81Zn
tCWe+Mq6s4tofIEt7lecpO98RUXrXorXYOC+V9Z8HS/TsyZ3+sVkR6gRLZNcfjg0
5fB4PQiYmpu+6Ho8r0UrB0m7J4CD7rF9bZMD/lMPVP8JuHNrKMLOoPSy4o87f41M
MW8uBLlotjyD/9PKpvUoykQqWZ9h5jNhKurXwdnKIygl1qhwvVJO+9i17Byr5phr
KuK18yoIrVGdJthUNSTomnEiu3h1gHRSVTexAfgXWOMnYwf6+pvszLzilLqr7bZI
EyKuIGdoYVVHjk8zOJ+T24cJdyGOJqu5Brj1C81JeJK+lOo9JSVAsoTf0BHVravU
VihnNhgnU+eyiF3fecR4nP/TjUYc6T4TAVyHUn4ZpNaR+4CsbVq3ZGJwFbwRek3x
YEvxl0sfxqqvDxBlONwDkn2ZKOq+O3UQTezMZ/OP9irXmD2HEdn6NZp3bvEMwjZ2
HkAb84WUqhH5dpaJExhtOLwtsXLj82V5YptqHLuUzfopmu9ivwea0BAzw0ob12d0
APH5CiDKz4o4+w7RUAsOJGAKsWxakZ9xpRWHrqNOxhi7SyrwyOxdTwc6WdsrPI2z
vCySJmY3l9IGVNZbibxjjqal5Z3FU7OScp31K2hXMqo9EGcttGqkmi0ymbpgLmWz
+5e0KW33O31uZ5IuNJZZNEFyDytonfxr1zHFFEKp7IHXaGhiAAW70D5QVkWqrFw+
ZIkmMcGhuziUQZRbhdjcou077TuEIrOcd/a/DCjJHOySHzDpTPcGBrI5FD3cXU6b
JdcEhaLWk4WurLo0MPpqW4IjSXK0aCNhMzSqzdmNCOPzxi5bV2p3QPxKXSAUvNLi
lY4a0uDE8tojWPED4ltqVxmIDTHpMNfmVH3FBix3FoQvQXX/v3R6zPOhAvJldIa7
YgFEP0ubTeLq5iyDkgi6pa9pbOmC1aMgn3VTwTSnvp6X4coMnw9+tjh+OX/8Pkno
aKtjANwtn5KAa2sRJLTWVHLm0q3S+Sun3TZDnI60W6ch6ykkRFzCMqCcPmHkqEpJ
2NoBdQkmJ4lbNH6Ds6NVAJw/cv8opnxchOMuF1SK8DYHW7NPvIZcn8ni8EaH4yDF
dRMpIHRiR+Q6n331yOeLgyqa21/kD3oUIm2skvu3tOiXWSFK+NZJ1AJe2De2l5wE
KcyPkXuKeaJv+b2Y0U4FJ5358raeBmjXbP+/TvwETEk3C3x7IcQaPN9UlgZxFjrM
CInoZY0quI33c8EePZ1yC+xomd4kDCgSdLzLV9i/rlM2Z4to2CZH63MgVODU0IZT
+kUoM8GRoYDHpzXjaYFXoYiI4qNzffeQ6kRIqM0dO4blaEYN+P8Yjpw6B3xoEo3u
wU/ALsMisXcWVMUJphr2MUWi4RQvhfCvRyYill1Hlm5MjrZdmDdffGwVGEj7CBDy
xAQf7qRy3CJSVZIdGeWKPi6g6Jlz+QSwJ4x8j8KcK8dxRHCl24blc4FOVNOTdMqJ
G7La3OkwFc2VR6PZai+S9Hp916e0UUWUJTDT2JCPgCqxDFMY1E8O5y5ky1mz0V9U
9b7nEcOjDDkHQe5fHG+vQ0MhHp3lNXEQD/b4QAhBoIPWqfc7ZaRUpkTUhC0N6FvV
QhAxJsEZ8FY+o4ruF/KlJ+L2j9QwdNukTFJ1d+zNch88ptRmf7+ELiIEMRecmmqk
d/9aXO6fLwZeH7srkITp4YozH2vmTCU65cOCeu1yhC+VD6ITrAKhbJKJdnjjYpYP
UUliXHs/bLvSompdAhuwKq2zj6Vy7LvDVNe9C42Q84vDllHEi2vgOukjU/wGdY6W
U0wmyKn6ulVBe+iW//PKSMrjEcFt3YSNiRivVkCaus/2qGgXHFVw/jXa1SyIADxF
0C/ztmdKVwkVAmJ4WuG0vfuwaeO8W0tuBN2uJ9Izvs27mtUPHmlG5is1SPDt9auq
TqHSXLVDnYaibRLJolwX+u+rF39TwwI8ysa4M40wqtYJ4KczJQV4bpYHckOcLT9G
r882DpEPSazoeqvguq6KeYTC5muk41Kzc6mWR0B0lXAKikWnvMCcVLsxYUO8JTTe
V4hc6HBLy38LVQqhwrQjjW5pyvMk8Nw7rTXugW0Gk4eWUt9xX+dClEGel9iTi7k7
n/kDk3zwFanISHuRrKedNCf34fBaxn1dzioe8EeBnPUr37+jHbslacwJpWRPr5QL
qUkyOYUjpt/Ax9/4Ho9P+hUd1Lz7DJ91bGMBQbfNsuIPT/nw9gsA+YcUIkBpMEM2
5CfDHoxFQtkiue6zhntv9JATjBwzztTifw4UZFsF0z1yPCTP7ZF0lFlAIn8S30iW
VgxbmiFjYxBP8OpFBaVYYlIVOBYqJR2lUjVxqR7m5wIprlJfTwN7rITSKbVtSuQ6
TknLZnrlZqnS4nYzxF/6/MunGNIGc/gwweI3992+MQfAuGytMNNemb7AZSFDe+v4
4Voo4zXKYoqIO3DkCUb9x6e3dTAnLCmF8jg0NhYmniD0VOau11THqZrbVTimcHBf
uC4R4BQPlV6TJml0hr01zrHOoB38nnhcpuNnoZWtXGDoBCDoho6dnNVZuQHjagPV
mRR86cd9aQOJJZKHq1uar5oeIgI38YSK9+1Z4v77xwnxi46YbwA+rd7SvfTJy2ep
uqWbCOgZCV6DDRPQF18+lVzq+66q967VBHT96R22UjfRRommdTk7deXCrsHZZkB8
6TIsBRTVY8x3zj7iKmHziCu7FUJZsDoysPxC2xJf9BlCDcsOKGFQevVDveD5Cwvk
uHF8xvtIA/fAzBgunLf9Zx4Jf9GOKevRTh9aiRBsLXE7fJ8jMvLh3wqrVbfbAx1u
aQss6mgL1LYUq7fYYTobej89Bdo4z9RJBdqbdFQzQOoqotyohe1bheHweMBtxch3
aaYogfJk25Q8vyCLlBLrs6hUco/7Wyn8/uRdeGa1o/e6fv+yKJ9CQjMEkAucfzGA
TAtvZtNE+43NMzrN7XhL6ZxwUB+TYfiNSsQoH2q7dQx9fdctfY/GxSczhSKOPtrd
i+jH9lJYVIw6l69WYwZNORYLaMmicgVtkQTQxx3yJX/0fhD/mdzQDHd2Kqmw1gYX
4IL6xxRnHjZpKnSBtNREFfjk7UODQcskAU15ONy8S0MrMpv//2gPAo/eFH4CkozE
rFtKy5gHPnE6fTyIHuqYHjJvgZ9M8taBorPt9tuFw3SqlPu67P6d9a8NgHVT8IFG
A+m0e/BsgIauG7g9qvvtDogU6cv14XdFqimE3nTEG0sMBZYvRCdSyjBKvRHKnGPj
94QVvLqCYaooITdzOxUEhccHACI5jRhC8pX2vxBnR1wTaUr+QKOo4IDmG7DpjFLT
Tv0fR40rzv+69WDGe6YOzL0r254xJM3cmpZ+wfQ3VwsyB7wgOnMNzcDwBIciLzHu
GI7dqnzUjAbl7wJAASkkRZTI1X1LO6r8hJiWj8YWh2e71hcKUgFcUZ4FI+V1bpnm
co6ckHekqQHrZMAIhHpN8nWBr2B79L3KcPMmtrkFUsrFOyYhNVjEuqUzMUjbLriF
WLvjfDnLFrBOsOXfUp+PkcgIiCraPI5pOu5l3EHtOg93rvv9QiBl2CWcBUAHyLqs
NUWE0P3ojdTUA6xsGm7DUaq5iHU8mZs7b6ZCDeWaRqMKV7xlyprreOPqs08Omki7
L67lfECC3B8tbXhDxfDfDf3Ahq5MImbxZaPNG8y58PECfMVziZZV0WkHYJJal+Yw
q8sla9edpSX81yI+djWJ1B0Q5t18ckVTjrLmy4uikxPnZtce3L5GxL1PTaTMYN5f
o+/u0c8jI5Yg8R3B2/Wmko9At11IjkKQ3FxBR7MV0OuR2rsW2ffq9wmGPNg+9nYr
PXIsNHz886qfXajDsuqDCwnhMJ31kHzCs2a4uVeuY6bxyAUDxVCg9sHE9jV8oSho
gEdq+33Na6ElFjbkr6YD+yv+b2okltthE0HH7M1GxB1JHAlnbncAHpEM2bzKvNtg
qUWu21KRRHQV10zZOC4pMKYoXlBdIbpriT6E5gy2o1uDbmGwtZlSPrJGklqJP0rT
xJeg4cyajrB3T6mGdmSIVJzpXei2QI2/IQ5bu2LDeM1MA9svD8upgVtnga8NKWWk
6GkPT6hiXFxdSNA5DVf9zpEETbY0SpauIumPJVBEX7kPJUHw8Y0H+k5BToQWmqiT
1Cxr30x4ePnOLJihFFspj6QOW5N7k5Kd2F2EwW0jrwKCP6ROJkGEt2eE05G0JlqT
yy0QDZJ0ahRI2s8ctely+4lTZiQjA/zG2H4x4t4qcvoYYeZc2z7tq147xvL0mWnZ
VmEuj8phcH64jiM+k5a2ZWNUOegTOR3Wc3jR228WFEqNkaujH9G8nP1Nwp5pUsBQ
UHXsgsf4pUt40dJWXo5U95VLpQKHQO+ZahZu0D0RVVqnMCjaZX4th8tPwPaUuPwb
Z5ryQ5j/HgX+6e3WKWs9K3faV0EUjBlMo0a2agE/HL0jyOH3FxVIkgOurrsyj5kK
qqPbCY87MYag2VpWBQnf1GFwMnwV1aoDh1bpEpxT7qplIr/gUdztoKvWqqB4GepR
vdGPI6icMFfUN8UbwtLwkIOAG1XFFm6+KNErSjRfoopxRlkw7F10sWGdyNUv01AR
nZ8h87jivQrvJnQExPrz+vBXqeOpn1Xkwkn3CBC0iABIKsh1Ofcj3K3OdZeuAVhp
JIzbaM6H1fx/t8ncbqlsZZ8ccEhQNIuPd9LvMN4NLr62NOzbjJq8les6rPpmclvF
Mr9scoYWjidIPvsB5qTRX5oHF/AxwtqJ3efU8ugEJCRfUDH9V1kW+gpPd+YrwSzr
R/HmZEzvKc+OQ/+7DJuJYBn9m/tystcrGQdUVC9qdR/gdiLD51yS93nvL3YK2hKV
sTbD0s/AUGVv5Bru2Uqo5DqbYsoqKmYVQDr6Z5KNwoDSfatl0H4CPSFI7bKyBWa0
h/wk6rJSmH87Y1dI3yInkE5IvH6Zu3aDmb5DcPl3ayPT/9QejDx6jhZD8gSY+Raf
OClSuMGVPmoliq/8wsmsa6a6Z4zPqrsT8QPny9UXqPxuAFznxajIes8yfQl0FunM
5XXCl2GHPIn24FmJz3mJH0kDvx9LR4ryYRIYE7hRtFVt7hVVaXAPS+8A9/JlOS4B
O61+Pa0xd0Mk+BAniKmoYxpu1m0x/QbVTeYMGiJBmn8405KV3nL6/+MlcVShIawH
XeiGszdHEnDQKe/DiI5mLuS8cESwqhEVoSospf4LYCe/x1999t8sweten068YHuj
4XS4NTnK/RTOBheknBTWNSxTHVS0Ss+NOvIuQ8wBvl+cQmbzrdjiEQUgb3Ks5k/S
eK30sRHCL5mCO+Z9Xg1SMLBhjxDgW5OqeJU5vWP4SWa16PM0glbXUlIm2+g0Z3Cz
WZmTwGOmr9BAgpSNAPlhqdttTR4CyMh8Std1gDpFh7e7g7MmnBl6QJYg/aWgIcv7
E9jmuH/ri4Wg8ckrk/yseelRJxTOSVSOOec3JVbzOmh40OIqfSJhlRx9I0inFyIj
Dd3kJMrU88rAwdpP9/VQYjRHBYljzfpLKYVSRJ6Qs+Wkl1L8YiF00u09Bh5fZD1b
YRFNpuCL4s/g/U5ui1VnbX12/Rz3jgOe2jjIcMp1te56ACnrwJWi4Q+7AVdACWTq
g8Uy/1BJ0QwP+xu/nMx5RJLRDW7RYmlk90MGDubff3pqw4Ue4gS3AEBl5AXF3FkY
HxXC7JFT3eLW6wSfqRt0jM7xdYVqhvedXNgMNuUBjAw5fM24BNl9AjGvZK8ohy3M
DareCyzAq1cd4ZrXrOtv23BVN3fnfbe9LGbcDK9LvIzcg8qvojEWj80TJV/chpjJ
Ped2nQ/Xce/Wk8cckQtjXkIetrap74wMExrFGf4l8FSQjGEG/+dsl1m0G2AsAyBa
HX/XjpAc1VtmGw9iLU4J/D/i4CcJ8kCr/BM6oZ40BvPnw0zerFvgRLSpn2f6RarH
SuZ3o/eGlaXMG0EUx2QrEcRgzzO+j47wZQ4Hk0nLLbZybHLsXuSrR543tm5uqh+Q
iN+DXhS8LroPfVgTBJA2mK6T+1qsoNmUeOd45SjL7YsBFgoiGW9tnmNp3gZyArKg
/YtGs5m1NgRCzY8UC4QF2WzFYH/Q71Wbr4I69/ZhV3i0/VcNg28CJ3nDKarAcuq7
7p2jalGDmpwmg0Fm8LLWxjw25vNplpq5JDufqkQVuALzImpZbhi6sCAZliX9UFyq
sGdIPhZGrt20FIPQXKng7aEq9OODmwarF4+ktdVJgiB635Ff7V0qc76LdYC2Jgiy
n7kYjAE16MqERbiuzOzxhsswhJvPPkdzQHSGx+RcrHm1rpiC6gLkTbcmC5sDwcmI
TxIenASz+TeidJjKiG/iH+/4vZ1dbz7H8oJhnT9w2710q4nuUDwhFhAAxX1IQaoI
3yYRSTFf7r86MyjRoso4a50XB9++xMQUzcpB64x7u6zBNI2I7TONvWxB9iOoCBeW
e3JScX20bZmWUWT8xPi65haR5GaX9n0RKi3WNz65mdHoYmjcAIP5L3TZRnFfpTOr
0NftR+lWn/1IaIcQUmWCDIApBtGmK/+UaEqQ+oArMLI4utce50ZzfRsHtvQxRCBH
oFjIhBRZvYgo5Z6ZM8wQnXRbC9zMepscGrP3m9dXCVA//INYB7Wxn7ihZZw/je9U
r1hODQDPSErsEl4Zm5EaynZ6QQ9cjuTKIfzaK7G5BN6jTi6qxlNbPfxGDgBxer2w
Thaz9ROKT3mVfNXPHoJPbmUOY+EIjxwQuySbrsLahwQmLEdMRcxRiDUkwnSnZsgx
e+sFs4ePoq8BZ4wDbQiHtmGanV9+DorDoEhy1m3L/A+RwPSpuOyPhGVYgZM+gkqp
P82x6KZwGgdfJbRUTdKb26Z227JNvrtKxCwGflrBm4fLvskC2x4sHv8y340KtfHG
GHmuZENCF44Op8ehcz5hZpd8SQrT9mem+dyaYr+aStT7LkbE4xL5oIE65j3jHuAM
3zqFeDLl/9NftTXYtROR/mXjlMFYcxcm9PlZ8y6ZGwfqi6+vTiW9RqLWhg+Xppka
7XsMmFUt0Nag0i8IWV7hH6wwUt4sU1hwJIBGu8aXlHAO7h5xI+3gjlCQh0Q6Qexw
GydDAE/tTFR67aTMD9IU6pwbnFke0N/JP0dmhLqR+5WEZDWUFW3eKatiW22TMpp1
PbVvywk0XF8g5JUNC5JOJhqL/sLgzSAhwpjhgliCqLEFIvaDunmd4bJ7Rlm1eqY8
N7tbIMjahEl40buLUFi/0pEB2r7+SFl72XX2HGSPpCdt6eI7A1l+1V3czeSe4rnq
nOlJUayOMYLYHhcaHicnag1B73nW2gqVVXH6VmnrS07dHv46mf0oIeQkgWCJ4a2T
Ui6cxxh9VGSqg6jxT5IOM+/rtLLbeTKAA1OiBfYOQffYjnQM5weBe/7uNX2Fnymi
OnX2vIbUhL7kpuvmTVncq4/5w2N+sF3zCxneFIdlC6IamOUUdXj+gPHG5zlt1V0L
ekWkX6+Rf7g30XpFTx92k/yW9/VhUQ0ERLnTmzkH4K7r5XB2uXmEs06GxOkvbbJX
e/JAbEtachJSjxYZ1/0+qDt55wFrTnZB14LRX+IwwSt7wWM5dL9cpRC0fVYHlvBl
qoAfShVjgUYr8fYUuACaCpAEW1jrzXCzGYO6wjgYQgZQ4SOyDjj4CbsVJuM3lSTa
ZnT4xQrgoNn9ku5OmwZ1r6Mg/Pmbo+yWV4leSC4UHmm60WXxRQ2+//MwlsqD6y8I
5oT31XPNk5Kl/gRFBkxHaitrYzZ5GlP0akFw4QrRVpUhSjsvzEBmEnkPji+p2MGA
SkzNIzw+mqWEa0AQPISz1ccWQteqgAfLoJo80B0xNNUIJuA6edlNtca4YrnrAxQ7
p9Q2quCGDbBkIPUEDTVMzOqL2syeWiYZz6V8LjOPsg1Bse6Xh4fITU45HwdVbODW
1B1eJuLKNCSn9zSZCWa+52XiWklnBZ9VO/1klLwtrsKLuEoKbYcwHZ48I5arRsec
PdY+aO/pvN2IG9ZScF7DqPqCf+EZuQOeCCSE9bSp6gUVWWJ75Ie3zLtyeJC1E2Dm
NbyjaIZ8jVrOq71lc2bSwWbnddOJsaaKk08cfI+C4WR425VRlXHgH0t8OjJQHIy5
z+wp+fKZNuOReeH8o7WZ3bouxxxCb/dffUB0v78DgyIvJL7qiO73Twbe9Br8zq52
+K2F31H2+bQzi+asoVKuXqM+qnQpFAvPH4+PIxk8tec1g98hUXTT9tYRA0z2R7Sb
3pegRUuE8fQsnHiZh+vF6DiUafsLsIQhM4sxIPcxODhP2o/Q2xAuCi8z4Km4FGae
e9lyuNyAb12AWo6i/wVTmR1kM/7XFDhUqVpbQj9e8ItJh3PhgmUIinF6x/7aRIUA
qnluxketxpN3YRM2AhUD88qrz36wtRmDFDyiWx2ad9xBuahCAHKVr7HQgrEESuvj
qzzZ6pUrJf2U+KFLQpuCj2VFky1s8yMEwkV+d5bJK48zKXgoV+YrxvJC5iuslfIe
ZrIg62AVBElC9pOEV91v94FSk9j1w+PBcckRoNiID2v6GpZgXf5lpxcpt8Djx2fV
CBmXyq9nNzVRfMpHB5BtLqXunsTTX+u52Or1I8SkXln5C5jonr+OySMb76Mi/N6c
8woysgLuhVQRaZT8KtbsZ0qgGZ0Q/vc30vXvlOx2MhJ3eFwJSuE3ZtapUMuvC/I6
d3aVvnqBaI4E+7PZYVjI7hMoWPb2kkt+39uJ5OE72hdxNUnuBt+A4wBikf7cLHAL
/zPDx/99KedKXozgCXsXnMsfVxPdKESKepAyJSDPa9CRfvRB+pP0jY99fJwxzDNQ
DOAbECW+tgT9qmNHsKvzg1bTV5aBpT1jJaM6D2SXF192WISOibKf1rQNABhX3mfK
Ty/IkILvTkyH3z/WGIEtJmtOmemoXxFjzY48eQQrD3P2eNC712/omgKAUi/1J1rU
twebvwEEhSm/bBjDcumVe+RiqZRFI00f3XEFJEiap7c3G55aYcU6CaJuR5J35OJa
re6PBaT4tnVnvEPG8LhwpwIaEAHHw4snEnUbhDnfAsxvPnNnS1+2g4mwlni3d+3K
hfCzctGe7H3F1hKacnWZoVhnoGjTKKuheFDQ0R0vsVGd7LeW+LvD070EYHb//1qg
8zScy/8Cl8TqZq3rg3/j8orsWV8NY/jlNKJ9qSFfkhkZr6oHHD3H81EMpq97CiUu
i0W1dwoY+/kXMbcPWeASprDwe17PuYQtwDOefksuez2b3Xg8ZOVYs7d0693066ni
QOiPeize8MZUwtD9qPwJJQOiw1Pt5DhfW56ErkEsLuOLTK4cIsvgY5kHT37qn4V7
pLWErem37DGlyOelEjdTgv/YlzAAQtx8ylLaCCJGdrlC+RoGgpfzXLP2kvATNrlx
GstnVDlaeLE5HN8/SOC3R5PSBsSnZr/acxQ7mNmCN73gt2oWvbXx7K94AMAq9iVH
+mTWnvliq8IUx/IXdfh/dSy0ptSk5vhfmGJiQ5IS6P41cg1tvf8RqKD5cbOn7k7C
4HMNkVLrxFuphWrwpQcNrl55Lk0EyDjqG+5AoDw/XznAJddVZtGx5FI/clmjRp74
6UhmztnVRz96wq+5RudX5j9CUTBrIXLvPipvk8YhYHhs+9M7+GGPR9yncSLWeUVU
mjRAgXCMa//gpltKZ/LmFKz8xVdvgnCzSsjYSBTzYmKo2ZwSG/M2G+ivRhC5ovNF
56gy8y3N5UnAs2reqpY49txm1bgKrP2WW9QGI+N0lTFhZjVHcXwbM1Lc6MJv2J5D
r+THyxfYCJjt4PcFdcik2bQ23QggOddnuwET1VgG/U+0rHgvHzeD9Kx9Hs6dsOJo
+vTlWmQgb2BB8+qnerd+DJjMmmxQGhTzQ9l1DKRLrLvWJ84lz93RgmLL/8kismcT
Y5N7BOL2nHzt8UlqD9xsB84h+DTikXm+066dDp3fPuMfyRUGLAZxorulLYUuAX/w
AMF6btQN7QHJb6HAxqHhPDylpWqpMYkwIvPblW+QK45FPBEEAWZzg3rU/lDQ7Guk
uZFcjvADT8jqrU4bysgM20xp8cbGqHwX5T7Ccrw8wFYwyowvlJjK9nK3+rVrYk2r
qx9umBGd6lCJgtZKmcB4wbrSU95qTJsJ83m9T1TGQMoVDr/HaXk1w41EzYUBh998
gZW7HTxO6FFZEMj1u++IMyiiM/mN2onSEVC6tdkY95eUCgsXTNoxJnc2YzsguWAI
0hJp2H5YS2+BojR39sRoh6QBLweDijIhyVoSA3DbVtPuPxCPc0A1Dq7/pPJnX2XA
xyUG7MRnKxyFrHfOwclHIcq15ts+6bl84zDSKq0b90T/tmBFA9G+US53wZndGJZv
oeP5DRlv2TjBb8IlGgjhVCCnx1Kh7/LhI8AbjOpZ4lzejy/T0VKr3SJ5JTaEC+Sx
W9rFSm0qIwIOTLCPK8GF6l/nT1feaARizbn8cEyv4E+OnIrGi3oFXWfXaGOBbbyr
7W2LzZp1gSsvHZkQqKWIIwrHZJhQvYGyZlAl+Wo8AXOaZsAt2RsQGFU6Avh1qzcA
0shu+MX2ZYEFAHINdzWoeW1secZjivJ/rxSGBcP8QB4OPyWWIOrnsyMX4t8QtV1g
FUyZCzQqy4zzSn4NXxQv0Ksaiuu7mFig6k4hZzsa1LvOy/IKIZDuALakxTbVfcWv
pttGhFZj9cS2rBR3LPsvHHygEGaD2bqheAGNWuU5d8Pi1mNC8HbHE1qP8YxeZajk
UuqMG7mF0DusFD6WtXVXCZGi/M9gu7ypnf99X1EcO9tu5Qz8guVwbLgsdqEDodSH
Hf3xQ31yxSI3gD3jtIT6iK2+eP8DkxYmH9s1b8aCstpaclTDDO2r3N7pMrB2X+q3
HFNY+0co1SLnSAFyaZmPpXotqzL+uDo7zsnuWl1RMXoxds8f2958S03HSZSeo4fz
/H2eJDjm1aIPb3aWX+EdY5qZkbGoaigP2bAvgACdIeNo8ZeMtgTU52kf97kOd4A4
tjnpe96ZssFnD5DVgEINn2GXJG/2Lv+dmk7qSsvX++m+fF7RqCQovUvfNrEBpKGy
yeI6TzSnpBspH0V8+uP5AlgCaJKlfExLTfgCaWH5xuv23iP+MAlEkenkc+V+Ygx+
0wPBIzmVjS0eSVoKaAS+5aHrzewi7a7VBEvqkPSS7ycrzZDafPxNR5I46RkyV2Ah
9m3xOFbFkWnmEU3PvGllFq6eWpWNgcHwvqR/ByTnCWcbzEjiHLcl4iVlZVljmW6h
5DC/sfDZZ52crv3/bf9gKrvZK6LkfU3oT75UG62RMVtzS07BEa0vXSy/pfJTagFs
REA9j/G9Rkq2j0zyswLqmi3BSUAHpEjgAjlWh71oqxdX0jY2cTpzv+Y5VOd87kxD
oOPqI6/8iW6/6g8qWGgD76MsARhe4rSqU74+BFl+RQgbMg8P4I5Jjx5vEfBW8bZh
UWtdvtEq1sJSW1BgXahQqJUX0AkK7/F/hbRc6DDpNCLyNSFKtM3rF5mdCwyReNiU
lqj8+S3rOUnce9b2JVseQ0gkyLhL+JZLlnxyTalGVQxCf3Zy77NSoQhhpqs0sQHq
ESUfvG7GaPdyc7H/YkEqQjm32Y9uwjt889KQsQT3qP5e+cgg74ziTNN5AZKOHbbO
r9dh9ED6hlDekEak7p95ezEG5dgQGojlzTZ1efNj7AX9da28M0syar40b4OsIHvm
O2Kcu7489LmM6DVaNbS6pqQbZQQQ1j0BhbuLlAO0aK6lRqjrTyPcCYfwnz8cEofz
DtUG5qkDUlCRfUn3fcV88XyGORdHIhpNxEHuy3Bj41WnMZVXLACjXS4qbuyVjP+X
wh4qura24PRFFQUW6/NtBliQPoW3z+R+BAkw9cCJBR/8FzKY3aMZtddLYibxiI9C
t4VY76Tx2qLTJfgoBsdAFT/MHpxvO7biC+owVk30p3ywjVfpCjvE8BwkhPjv1qm1
AeFljjKRraKCmdGOwTdYH3wedS5PdLWOUcue7kMa+ltOg5Giks73gQj0iTKb32YT
3NnUcA34IkWjnRxXuSOnaUJDNoRkrWXToBJZGgN/gcp+bKTuMWgn9efvXh/EAyCc
OtgSztxN+heEHcJJGqS+QhJ9x+p0eZtlmZAYPNJrrFr99O5U8p9ho+nTsLlkV6LY
5Gk4XrEfoKL5BhveovuWHfvjoDZF6C6K/cLuc1pnHm2V5YEpg86pzZQ7FQD0h1jF
g9LsyJ1UWrKznGvv//0hSIMTs0Ah4E3veNYXfBW6TWTfZ+13Uly/eez9lgrk4H+E
H9P2SdZgqUQe4lq0nTk9GKvJCDFkSf9UCk2RXU2EIsMc7Yodo7zIc1fR5lYWu+RE
ltmFz5sr2NKJwCYBbmo25kHyNgo5n9x4MlkDc4mNkPd9UGU4RZ+PmELCrKtLXWlA
TQjyAk3rx03+f5dOKebbGLXuLEFthQqLtshgD7ed2rZSQ3HXTnYl/WOL0qYcqGaB
KF5Y/a/ywI+3QDSKS9jOgbcmu2awuRDz6HHCfP6YTiyEUaabqLuM35iIY3LtK8lw
iRExRSrD8Niw1lgXrWDM0MVS7keU3fKRO6rWA/rry2gIOxlLBEewfyk/Qa9KqIxs
Kn0zI2ptZEeuNad79zw+miaiUToHMKdHzsjc8caXlgKY2Pbn3M2X9G7EGbo6lG7/
e/Vx5C2908FzePYbCHox7PFmfBmkQvam/Iwz1ZG4Phtv+GQagRQY9jyKQqLAE7sW
dBa+PtdO+9eeMruClp+0KaWcu/Z3SLarqyierkSOMQEo+f9lNc+evXHta2IF36uZ
AucZkL1u1Y6MhS5a+ARJZG4peKYQaM48GRhNxFZquMFcUJzhOuTfV9ldo7/tQg8+
A30URTCQFUPMn51496zWFQ4oibLM/lE73rc/MBISYYAZguh2YVQdAfF2AjpK9oXA
skYqW/bTJUoSfR3uNROZ5+y3Mi/q7xyjQRerMjSPGgKAYXXz67TAHOcnH1HwQw0n
kkaGG/15UA8k5ORyo3G6Le+tvKX/nyaWszXKJbxPUbj/eUvy7BOS3U3RKHA/Uys4
i+qSc4LPeYGEBq06oglGbBMm5BGIEooVKq8/hcpVQij6SC97WprI4qLbbcFxOSLM
VnWpVkl4cmwR0M2iUFU/hb1Qo9ucs6mKaCiOEBBM2zBHSFcEQUKSDHf9VylBZOng
gi0GVa895uAs+BXj0RhthjRTUBmx6ihQoTPUfLNG0KRuS4im2YMcPOj/aEDpSc0H
CqVtS+XkXiTFE1pYxMLCEhpwbnSNS8XifRx4XsFvvCJ5wQHi0EShg91AIcjaY78A
97GBeLFclX4lb7TEI7ccHHqI2ubM0raB1gK1hHx7Om01LXKbRvURk1OGv2ZrzoEF
DWaJ2OC5XHnMJDlGQRm/VxM8Jj8jnUAZdke7TBPT36FXE89HPqbtbSEg4B25i1fH
BXnNrqu0MSj821H7tZuiQgkKLxBFvw1LjQBjBInxqgTByNW9MVIXlQ2NH+ESLi/V
/kJB8vPWxrh2AEQ8RBoguuVrgScC2yhq/VdI1KlXEL+eb6be0OGdMmrFTOEgUUWg
GLi6iogaW4Kt7dkN9/43SxSkhxuXIIrFh1l1mEOIaXcGeFN6T1NG4SxipAf/JIMR
9/zIs0v0FHz0cuWcRmGij2wykQJx9Gfhtb5HTFDDDoKcqd4NsDp03eFytICmz+Ql
36tdRPi7as5SDb5SS7u37Ad7eJ31upCllJgNABxk/RNF2UGzwcgJiWGzZGVJFiG7
KNXWiGdmYqpeYucQthxaiT2wyUWCD7z5LKHKWaACE5HVDxp9lqkJttAnioSq4ADb
zdOqFTTqIQzV/ZWjwZCcJG1Zy4LJMB14BmnLwEWhn79/p7hCAdSaKhApu5VBkYdN
QXv5jzHRJFPyTCBiC3KXZL+DqoOJPYcvIpFqcN1pwunDMSNLGdipqsZdYJ9/G1My
ETCJSajq14VvWvM8t4DQe/7CO5AWf9tM325mwfyg8NhPXFjgVQT2bykJj4g37fkN
GGNHX3WIc4bIod3YOHjLLCLeW3rAcGqQJKm201X3EX1FAkLtZKT8mfJ6LhrbyIC8
YOX8uh7UXaHPjmVhghIsWtPBQvyGr6r2dWL2Xf2m0fFx1xAVDJologC/xlUq8X2f
M4Mn0Co1LbU1JsRgPZ5B06htcX1pgCcOo+tL+gNB7E03KIX63tOLzDW5qUx+qIk/
f95GNFK9fJDJKURaLpVC59xSqqLLnCwS2fw76IHG4puIFkNJ1T89uzuDx2CJBOwT
VUuS9cET/2Z9cHr1Z/jhx952m6QB14BpYvuRP9RTxmWm07j3Z1kfivSwSadURh7m
z4AStNuhKHxXEux4o4YSaYa1B5SswLFdaSXhlWC5t13KG5w9yOEF4in8GPb2bqyv
/hAhEfhV3pfky/o1i786odT682CMZ+AN5zLE4OAq/pivcyJ7H3U5IIbKQ/6l6rV2
J+YZmUNspwrxNdUcI2LavdlThYuI6t/YrpnfPKzV9Nx11xynlBoFJr8aGjjXMnVQ
ZH823iCiOLJKc7fVtu3+b9Fy1PBT96kShcWQhb4vbvNX4FMOX9DgerG/0XWtkCXk
7z9hsEuVxkdZRjeoYfNXlu6A70UmMTQwd62k/aXOOllcILjjbPR+3qdxCeukCUZv
dIlpKxBB+dGjSMrw3GA+n8GD72uhk+BZ86rgiVSBPKuiBjOTFqajqxktDb/kXO5h
dV7KDrjYlcgX0x2XoWMg4sGqcOWqDI0qN7ICNHyxGSOUvo1DCHKRHzkqI3WmgYH0
T9tTjlRwJtkQNF6iCWnRjsI3zh3ioOHAySgi6A//Yt0wCQdTIolRMWnKpfrMWVuh
tq+LikvSDLQbdmSedIJH0ZAYzS6WSBX9Nm0kliIrDlFQNBlICQaG14CqlbIcP/Px
AZLbi3rHIy8hHV/WQ09fJUf5ZoQ1rIIqgOYiMOhw/cCN17ILMY1X5oEBq76fl80I
cwFmbEzlxyw1QcYTLswpw0A0rmVw37D+vz8AKDl0KqxiKWRpBvZ6vfaA2kPalE9b
fU8Jr3XpF83Jj4DhvGDyPITLqy1VbUYAeqm5Ay+u+FgsS54RGUCvmTsBGLyGSvqf
rRKwo7ooy2vksCz/nHZwYjF0DwLFGAdcCk4Y/HRay1MG2gENOD2lleDkuY/JviWr
ewW9rge7hZXmscfC7QZEsexZcAkOx8cT66Su4SWv4WITXvLbK5M6dKoMRlPrxd8v
Afpx/VoVWEKvDagX4usoqNRdC+f7duPSllS3LZBLz7vhW8Smv+RLkW4caX8zqRdm
0qfovjjZc5oUG066EJsPtuM2q2YXKI6pvrj8JkcKb0aMzBL/VxS64QPDa3PYKtGX
gShfCqLIUPGt1FTM699NckhCxzV0JNpLWJjdjxZ32ecgWrmFvmfLrn9MWoEPJBCZ
/Y6+Ky9v4uI2pKXC63UWpRUz2KBo5Z/AGgvGQwoe8GQwQEizKB0mdWtrSNuQ3Rfd
MJ/CAt9rB/jy9bALxwL9nLJsEcqXNHpgG/hFu3e9Er//rPz2d0bWNi8of8xL45cC
C+87HVSgqYNKjsZ3lnWg/s9gKqsxhKqB6ATVskob4auvamWrxJV4aOK0pP986YDT
vj915rySiABtM0dJhxeKUCk9P8EbL7cVWNv5phCk3l68oUm5USiGuNTc0bu/vv8X
Bt33bPNrAra1kwOoZViLBClzUbetKots9owf+TMkKA8TGldMqTnAZcbMQoVXBfO+
QNK4Po0IoAwTbZcrKYm6y9J2oMqIlnjz2qE9SzQfapt12Y3leXSa5AcsktUfWbCD
yX/fjnHjtBKMpP2UTq6IVzTAj7SfNmr0vrHxgkMuPn2f+wVo9TQjkrpMXaEL+9kV
xlIEIPaByLbg6I1tIe1f9VobThOyKe1GWXmdyzEcOD83m5k5htpVpBfFxLnouyOg
QHYwcWxOBfbxzX+Rdf9qBb9T6dDaroi9lFrWjlD9QnCWkqz38gdZpKtAcR6mKA02
3dKaqMzxjauJNKR2ugHi5/k7t1hx5QeZEuYCGVkgO8u2zoQTFLJtjP6Ldi9ikC4J
35GcwaSUa089jgbSKMNPuddu4jA5igipKOXfqtLMD6Q2rXhdlFo+e4Wzglw0Js0O
M5KP0yqOU2cKV7KYHCmxmK2JTwZ6Tky2XV8tYVX25idxbd3XBAIIojyUhC+T4prK
XDyqNouxZ5ktPSfTDQ0WghNuGkX0VOKCnJk6A2Qtz5/D0tRSX5EeidQxS2z9EuZv
yF6gb58nDkyKbeDNdPJDE7/mKX3T2kOKV1zubIwLA37B6jSVy2UBHpRK/SwcCz0z
usi8MAG/etgsWGTOSkEIO5cBPudWOvS6hJbgQWinqyWUCdpLay37HTvGhnd9nTOJ
HFGTNEdJt+kITPe4UbwWheriJgdr/ij9F2ANiw0Su2puBV12TyFIuiAS32fxGLK6
QmY+2GAyOj5jGNQNfpQto9phohPi09vJuCdAAy9O7PIJuDTUl5nIetDzbvjmMS7W
icBtkkg/2jhrz+iZWrH+1pVMztQgUY/UOVFCxaRogG5MV5iPyF9NmuPp5JD/kBE4
qiTdU8ZmwSc0oO1Qid3YDCvX0wRBpFeeJThIm7sG8bxOw34REvMpOJiIM3unqh4n
mZrTy56m7vkalBbaq4fXQkVzytxW1cumYNNwamyDIieknjiWeMsHQPJ/cP4gwToX
6qUrW2NAmlctGK4Agab721AQYRjAQdu1kw4KjWQtN9c5/NPi+4BKrGTqU8N0TV67
R+MkTDv0Dxoo7VSxmqr6lu4dAzW2uQe9Yn4PfEkL+RihfvhNW/lLaNfiagYz53fX
I1478YzHWSyQy+5vRyBCD6Lg8/y3UGKSDoBLUaU2JxDb69asQFK6Ctl3QBqJAsTb
lm5HJeUABt76cBB4Ut7UCQFUy/IRGoegS/CkYMCKlN0zucE0nn+076Ufsvr/op1h
hvSeLZhIbHDccAnqYPx93D+tJTtkjvKUkXiHamE+C4faBvGQgpd69BxD8/0Iy1ZK
vU+1uRGRW6M8zZDOHC6/esEd43KFTuXZf4gsfTDfLi3a2GslzGAbZJhpUTOYnmoG
eaeT82Ag6eA7NHMCOz5XawRVoojaDiOg7hhqKfdhmCf0dNO7cKkm3UM9+w8KLi8T
NUf4zZnLGawI6IFZKVdNWuBUuQnkrXbvHY/iFxQ4CC5CIags74C07sL7627bxTNz
Ojqv+3o2q0xBWg9jDITG6JXKzDzO91E9N+V7ld2M7t59qxFgZUq4GaE/gXeHoiJH
YR+aC5F7VTUgXCzv/EyFjbd/gneN7vBPZ1Wvamkg5jsq0ezjGQ3d/OdnjNB7qAdb
0V2J5fK5TlVaZDdpFRLCBvixVUoFB1ldBffvnqIE4c1TAKwDFO99Wwy+kqQU5EN9
idQgeu/WgqH7uh3hRV577M4C2Qe3G/fP2RBY8TMAhQ88rujt9g1tHv0zeE+s8/pe
PTe1YcogYtmDi9hxuanXl2wF/qkJAZrcwdQ+pMBY4NiP7a+8DWp6m6gW3z4KEyee
eu7xilBPpFWBkfVyz0bMQp057VtxxYYZ1cCS9AhWyJzj+nH7fvlSvvP0fWIQljID
blEUqDdFPVhGpHBnBkJdQ8tL5Shxw0+V5N7yPHz/I5wUei84A/Y4atEQWfx5ocIR
1Zw05xcgA8hcA+u1gaIIvQ+4FQbinMpHcc9ouDi+9kJ5bCxETmSerHK+9EmqFkEx
hT+VrAonyxiqLj8JYlwzOVVnDYnYUbqiwQzBJciXM7nzqqqVRl+WLmPnXauupP1j
PgdHI0APGnjgiRZYIYexLEUqOMZpRUibCbojy3G6cSFwQ0cXRK0jRJmf8BtIhS1p
fQ9F2XDWBA2s++eoNCwTXujILB1rXBSbWOYr4MF/mzjeAF3H+TAyHdJVJAimsDgx
v0a2GLLafvn56/hz5fhXj6Xiz5vYsKc9AdrpfeOXeJrq/wWjm2fFMqKpE13UCeNS
pGg75wxnRjans6Dn4XA0h2axWPotNhRSjeKEgj1yKhJv14HA/a4UKkL+KjSc1AdL
0iwSaopZkpffRkooZ38gqgb+e3Es2T4x53pUheko/IjJipndC9j2RrFeTieN9Srw
vrQreFSDBbiwYgoWuzmlu/xSxPhdsZk4cCH2BOpTyd6YHJYJXLQM1nAHe7Ppq3u4
CnH7gOpqefB4EG1DZ2nLz6nsQXuQtt/39nDEdsgX8k3abBdFJRrdIrhGMNbQ8AYt
nTd9ZH2yMlTVm3KErJEYWMwx3OUZ8CSC+VNaY/D01nTQbokgaAbfydF7Dd8Sb1th
n3zJ3dIrmsBmwKDNynRyLPfmz9J3jqrDsSaKL9QZcnwIRSyHHnzJhbUPHrhx1EGK
pGTLJ/X2awNx1+DGCvHgOwDYUExbuMj4VEpBZgtZusZhN6S0g3edz8NQYw1FCwIw
b6vmvqmbSr9TCVMdl4W6/FWjygq/HM/WOlu4bMSEpWfNLEiU0d2/xof/BfPxx+9W
9roy1aQFdqrJt/UgTUPOFBwnrm4dUoeKiikLqN7PR2AZCUA8LLgoSC+rCsdlelf1
4PwB8HDWUnfK9LrqUf8EVz7EzCzFsi/bI8O3wgvcptSLmXGgArqoDqBHpHPJBHF4
ofSuZF8es/3AATQWdFJbciYT69fw3kAMeMGSBDGtnRK3gBlvVO0+1c4GmwfcSbqu
2NhgsQ6fpKzN9BC7c+o5zLN81eDtPC/G8tLE7ZzI27DoaVJAw4UsTVKD2N5RNpCJ
Kwo+qXy4syuWANyloMwrH6haBbVTnpzJnVuvk2B6v9jBxqtmWgFLDCWZk9A3VKQY
P4Yf1C1ca98oqucmkL2ntYOTzq82SRxXNt+l/ZxKGaQ6gZNjjISMC6VxYPMyjDWQ
XKCM+HAEiWkeSkyLU9Jj5mW5QwZBWeyG7kBIheiPgMiyUrvP0VY2nzJwi3AoHSvC
nfZkNCPILN+NEqOJpQMeB8j8Nkwn4hlamo5McChaDxUzgjGI+BYPhb2Vr4dUMfOI
TjZCwpF04gqAmiUgnoR5jL+7MyfMCmb7yt3i/g3atC5LsxC2Q0NZIb9XP+K3fR+t
nKtDuGhFe/ZFbEtSkEcvEXq0E++y+fsiqcRVTRUzvz6pVI43eiwDwGwDm+evte5f
tGBZXiq7PdbthmTL5M6wWgRyflLfr7joQOhjS8eQLbSV5KYwK3thVOtkcPerpH3b
9j4tKCyy5UanqkS13+v7HA01LCcIuOoUAdmgb5nw1a1jhEuyzoEBOysajgBlXHse
qZAwDsurE1Dbo78Td66Z59AKVxm7Vd0ACZt3YGQ8Vyniw6wdq9XYsA9RFY091zyU
J70mSIDWHlFswXt/3M2M3sdeOApabCG4LN0ptpsOQeqGiz4ffnDIMX0JvO58zhsy
zVz06SkK8kdWshAmF0Rb7XzRH0FA/JJtmbC7ZT8+5ybVPs8aRcktyA0o/jhK4rrj
SPu10G14DDT56wFxGIxh7IU+RINEaJqgnfdkKDVvsmKTiB8V9qH6dBy0VXXVwrtC
4TB2Mkj4ZkYNRiTIYlBkY2YhWJGccJReOCKiOdLiTSFxysIoBBt+wpiy38ney9qa
AnfQBzAWGjVWc1KHZbZ9S35oFleR23FcXe2Xt2o7IHKMj21un5FX5oGE52GVjjZe
IPNNN4xeIrRxatnH4Eiw8HLkuCZtT8r2ReKbZu+jiqYuTlcV+OEJCueuAQwmMX21
f6RwIkFOfTbYQMxtvc0ami9miafrZ3leqaM3S2xwSXDK1zvIH7dCvC32FvnS+3zm
jWXytolotrAZxXGufWvVx9mbDGn0JpzEO0rr1Ma/w50flxSL3wgrdgFy7HQ8Xl2M
eYNuR9P/5yuKAORlPakEv6efaE9kd3+xBxovH7AEgN4P3rhSMgcxcbAsO2Pw44i7
O/CivDpl33KekJGgl7erkVIiM5ztaZsFakM6b/u+FloF1u4DsMz6HtGiu3N3RW2K
1naok/xu8Lsxe2hQFgA1hISmNmrW7JU6hhsol9RT4PffaasF3KoxLrUlWnr9KO2J
cz4ze8u+fKcoRndYF6UGuvsOSLRS/crIU0GteFA3uPetGu00tF/hibteZxtMHBfv
zpkMGC3acUnIxH964YydnhMGYRX1MXBTC4M95gdBBtdSBDV03biCShr7AzXOCZQo
UeUfmhyLA2OwOVVbv8U7pcy3vvO+vS3cXw+0XpUFry8jEV3SGP3RzBXrOqmhOwm3
OmnRiOAGfQQp36Ag6FO4uVo2nfkmi5Nt6w+CsEceNn+S+T9sfO3+SuBqYkHCNSme
lxnk7Fawf+gBa/kqv8yGDjFcnWP3vNPqvocJHYN0DjDy/mBRoiBUTATZgPQ9l/gv
zPeHpktp2spziCyNGlhWc8iGurV4kTltEG+2IuVCa6APyOVQ/OBixmGsDZj7uSPf
Vd4QvPZFKVCi/4sK7UM9nQZGf7xMH0spy7+K3sM6FCuuUAC5lDNlHZlRE0g38DLI
qJnenIX5hq+9eJbubGOMC7cGNTYqIeCJrr9sUSQCJprwXjhJWcTLNb8dcmM01wuL
L5HzNABvdkwLhJnEaWNYRjvWDn/ETs/miYr2+3LsrAABkrLBtAz6YiKOGBmjWWn+
5tvc4bEaTOcX/qkpL4TFvpzCWBsRg5vVM3oXmK92jJKF8NgnOUeJkWOMXi17PP6v
oyhnEuBJZwh1HZWSlU1x6zIDyn1radCsKYkypZfu80pV7uDps8mzi2VUwZgbvn6H
GjCg4CaFFkCL2G+AADtNra0QOD3F5IS0IzWTZuGa0oT8TbvpymPQ4TSEZAMpsOTk
t3LIhu9NYMeiv4BL0WseGjFbOUnB8obZODIFQR0jEdsnpLi02Lm7lOC/kozhH2KX
6aepAWamfrVF4ZO5G4sEGFmqLhUGXNRvwpWdSnpw1j5h8+tUOaieaK+zEXwQSHtF
BdTwsb/TKZhHQQVe1AUDbADwszSLwo+cgB1ynyKidASQ418jPIuYpZy8Sz0BGXQG
K7qvpk05dlBPqsEJ1y6N2SVqzRo5DNgRv4vXsQLol7U0M8kArbyzt4KBbzvx4hCf
i3eVJa4663j4iErD9Z2fToJT7BbpOreJ1qnnoTkx5GVMf3oR/9dbGdpa/EtLUQlW
h8Yt15INVaL33ckOMPT0e10WqPTe00nNy31+KKOWKp1HcOCMdqcWqhSVV/B8AlDR
J99ASJ2n1cLJASdVBcvqwnzckC+l2OiH+mx849+bxe2UwrR8E2KDhhUvc/+kAr+d
sUPumqGIwI92G1+ro5vJyi+uxEW9cseiZdA1+YXXlr9KFuU5Jo5aHGNzdaociz5l
Onlh0NAjnmO3EBXwPlq1A0iQ4kE5rU5HJ9e7djiTVJXNuEA0Rbg34O/fl75CGnHf
a9eFfTfWuZuwZT7l3i+FS2Oy00kYzW/jmLeYpIKKtllvB7zNey84gD1xYWByGCc+
F/G75liBFRL96BvD/xHH8bat0MfRCUPPaM+AETtQlkfJntaUiGp26o4lpBWk0Mqd
gFhjVhUXGQBiPs2cZSSj8iUL19NWxn/LkJJMVHdMe9UTtJCrKOz0fhQsdVPdkO00
LLDLtc/EmMpgCcWqphZ59BCv3mNUjg6MObeDfyU5A2XEtcVcrDHcTvKdFtCcJRwa
hbvHdFLWBg7RC4eHo2s2Q6upvKmSbExrx2UFXoW+hjG+EKfGQuQjaf7PSpR8QJEs
u0cAtMR96jHNSF+EBao3F5xv2MfJrbpTIBdLG/OnoEcJ8WjltgVrR5v/aUuBWj1D
NkQ+anRrPwoaXUKKwoGI1x0B2LhiNO9zkmsSaGfkzznDmso9aY+gDjoIW3gxl0VI
P3+zezB9svq3AoyZhHCffHVns5DVched4uxQDdp8OfLtEsBh4yyOGbtfWpanumZA
Uk3fU4nASKFBzmEQ3Ef+bDIS3z3c3VPJptey2bmtQ/CGG2VXsmMOPH9a5baPhqAC
klA7jOp+r8hbf52laq//j1m5lI2T7F+kvO+HrlbhhkscgH8eGdT9BknEAbF/Nhua
t3ZQhElQnz0IFj/AlQO4bRM9+bpxd/Z5gji7SN0/Pp2dRqf8ansFFB63U70+9aHO
KMicQp4G/mhqaVOrU6nwcKliKwsf8gyuNUkR1fo23oeC7Wf5Lff6XgfbdvZyX+iy
sU2cTjuu6VKls2AY7qA9WnAMxWlB0RYqt7G4CEVVv4l8xcBJLETqIAligqZDBEBZ
KXxN2yfuNgKL1hzkXgXCtY9Kww57xntEGJgCmlKU4D44rrPLsj9FpH0ebkpvXvHL
XCU2pGwR4cjdCNyp5FLwTEysYlj/omX9Af2q8+1xC5T4mHqHvv6sAvQg/NjhWI7X
tpQOIePX+juzt8L8smlWtPbMURXUl0Fn98x4CWGtWoPjt8Ubx2s/opU3CN/LwKkh
wQg91JrDVopBHZV2I6xpxIAMHL5HxhSTdlLmzMduK4ZWlGfpKDxivmhDKTD0W6C9
QecOI2Kv2DjGZ9IbHP1mEzEf1D5ybozVEVs3cooLxcw6VZzmgyGEDhmOWe7u9rBH
8Bcev7QXxOuYGkgFhUuVspPorS4YRrIjEP0U4Teu4VQNbNa553POjDL/MK0tqxpT
aTEMyr0q0nLPQYuwkObRl3vh5R5CypF1P8ZXJ9MGkUBVJ0WWfUcFLV2Wx8eR0ikQ
w69fbSngwsv1qN/Y0JAVHKkmxQ5u727Iyj+CLx8w7gXEncba6qBtPQrBYT8q1in3
IjatnkV63T1BgcRaAjqLFXgo84nOo5Hpv+8ye+yIx+aRWkZh3j40iTtF9EPaE6n8
Sfe9SVqK5Sm2Ony0u793SvSTK2pEVuykjo75OEiKaw0CTiOx6jDe23enxtRfMWQv
dgOMHdlBQ7YQBLRWlxWoRkpFg0xvifAoJ257/4akLHwhZctShy6X0fMYpsRDlIvL
giSqBp9GL0b7n0bACvU/7pPC0JzVnXqVrkJEx1xD1ERWXPS/iJvzHjE7xYB/nDux
guIAbLBmD4Fe8kMfED21+mMnF9Q/PFTNR5DGVEghp+bVo4Vbuch5LhTO9LEySSDz
+QgnwusyeCCKa9vFqVaTYNGA08I4X+QOIi/VBgfkxyq2h5kIiYt5u8460DObe0AL
msFy0yjHWxNRy0HHTKUQoIsGKJFZj1m1MswJRMJ5b+f1t4N7Tr7c50SUydfWJeGt
OEobwLuRZhHS+2HQ50W9sXx3U7U7LG1vBsC5n1FNyQ0YRtuvp8sG40T7R+0nm/13
PKgVMsyZtbUuqyr8ZYO4IKdqV3F7XqRVex9DHoa+0NQVLUTgJMmDogZEFvA7UXL7
unofwMpqNfFH4xtXgquKLIJWaip45TXRsT12/EOf5Ye3+hBVsTZbEdycke5nDpQP
1Dl0OhXxn1xVBJbCNWTUN97Fr4otKd3AzVfERMTiwWQ9sha0AT6FMjA4kN2NGDoJ
sN3R7s1MUpC/lHcFuXUZIEqH8xU+hIjXWENuVKfTHGZBeQAZSibL1hZIKeBM5A4G
MuA5nPuCjW6IZ2K5qPJWaC2spF7ikUgBrQ1PQBVXO0jlLkNwHhQNQ5LQdT60e04s
tIWTM3wK38AzPFjDl+vRVi4sYeR2N14T59YMGMtbRDWLmmvVsOf5lPp2nafVjIjb
NVZqkMVW7F4mDr4Bw4QRf/CwyYvJtUMTVArUNuWB+TjIIwIDtCkm3nXi7i2M3ZEr
hKZSpIVqNjoyCWzVpw9CTyIvhZNv2L7ieWgYBnCbfwU/qaoWiYawLQ9Q1ZHzAyAu
xl8KsSPT3W2dk+r+LXBpvvpEun3z2QPMAryzHROfZXa/BbT6IIG7S9rEHrR+kmhK
MCzlZrasK+HS1qVwF7DwIXVI6VPTwh/3gxann1uqrGr0WRT4sgD2EWb0MJQsqNeh
UkE6nZZ9MocRYyhHqLHsLs4zT2IToA+CxXjq5WyFq277w3aIecqJew4q2wtQ4hAA
MDus2H7nhrzRcXkWqy70cQ4OJ3z+mjMlAfxeh025YLW7x57UM1AggEi6A1ChZ8Up
4IBrS+/zj6qv6UaLn54n0GbEK6b/xyWT48sHQrdUVP/C0nwUWxg2xrFWqClBlmwv
PcTpUwzCY/vj3L9vY6rYjXmvyKt9Cqy0dGpsxFnlWxkWugg0u7DsR8yfGXsRGII+
OaYGT/imClighEu9rhoqF5lkdmZfP0XK+lVXNWIVTo3CuXgIjZG8kt8iD2zyMIQt
13ZRwA7eJKdUYHznt5JD5ddeiAdP3TI+/RL3GbFSZSNjZMp+2rXZEnQJrFMwByxP
Ay3Gg/0v/4o+0IhAKEXN9OMT5NBIc4Unns/3eNCV7pl7KvrRUA6j3zz+nObNeB6/
5RXlcl5/ImSC2r6e6L99Iptx7cQsjls91QoLAbHxYFMnLFA1SsWclz6/y38V+xXn
oVqIwzl1G4VTGUOWu7k159G60nJMKCG/QHnC2cfcuCsRCVIKQZr9asnGnMSFnQ0G
2JcvV19mfk5inT4u+7HChwpmQipQxJEq5VYMWPcmq4c1XYAyyf8Z+fAlO2gyCmBs
+g8CTomryGuANelmyb6Y36q7tVjN6U0iJSsrpTILEFCSOJzhXQObYi6vJeP5zwWM
wGHkmWaAwmsN+QgPi3sY3oP1xsutuBFCE3RFQ1p+ou7ZhsP29CMh4Wr8h0TukcBg
Lx8J5sohb5GQgWoxYdJj7XLmqn/hqBZfzldlXuw29wtDFTy0qG/tomVLB0RJ8zFs
DlIBXYcNN1u/6tYgc7E2NiElgpFxXKHAh03+gymInuJvdt8/qwgjNcxtqMTxF9Kp
XFJS79BP5iI5z0s2e50vL8i1BjhniyyfG9yBkpf6VNUV7KwvklumFDuv67Qd8+2b
qn7R+AbUUNLWVXMptcTtacbjCtPs6h/AcRrcZO4QyE/38KLxksMToue87FegIkSO
zV9vTH+tVnjYgihfr1hxYcJSiETgsprq2uO451u6aizX9kddSzM65YjbrOyp+7CM
pGcTf5apwyIkgP0HT6lMPESBwB8bZ29ujj0xugBFfRHXc9oOGNoRM8brbT+PCAmG
6HQQxsyseFW6pjBzR51O9O6VUO59+AlGEKKnFZlw3ZMlH+f/gwnGDVZxIudkcav4
wc//5oLUKh3aCXvS3Jzsts2qUV704fBux9ayvhvheBftd7MMwXqkpzwBD4iMQKTQ
e+kUNnIhARnQ9QZWtANTK0EGnKyKOkR9b3wDRWUqrTdJEDUW30AGxwLnmeNPziF+
KcUMID6fze5arZ9j2FtbZON4fDO1s9Yw7jzNhRd5VRtlCvRTYqbDOj1hHTzPXLhY
qbsZ/8SfuTacByVG660rwf9yF1CA7qErHeNPJudy/taETDrLOR6TjM6WL+bpoK3x
RV3PayjIHImfm2SUba2V4PrBLvPoi8w07C5IEoPyrjs=
`protect END_PROTECTED
