`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YdsiWHajv5U7aAfKIpWcVZDruskhjEfZdKlxKBYPSmjreD3bbr/QXHjhsNLTvDCS
eGUQTuq0Lwgs32HYTHseoyaMscg9x4pg3x+bR8u2qogQ5qBYrp1n0Yx67taclJgx
1lI+KS86szJFV2DlQhKIa/288HPb9AICWbAji2d0yJ9X4bpowrxSdPSRlrP2p/P4
nBEoHLZSy4ea1bn44iDq7f0tax0heF3Nlzh7QKifRUckmk3rAEqZbPsW6ZaOCnMH
idVj20euBL56gh1UzWCO4x8BY2v+nzHjpmepdNemBtTydwa3wpIB6dvOf0Ko+ZKo
1D7CxnMEywVYQUvS8ygNoxCJJvuUZNsE3Ve7lpVwRRdgW0Bp7Kw1Vj29PGxdoKz/
37ribbjWqQyhMGM+nv8gyKt+5nXUxf8oxv8Grl/7imcbyUUQdfLcoSd/qkIvgZsE
fPV57CatQrPt636PBjFeHzvmdi6686zyx5DwqVKhk1tG3gUv7zaU/GkDXKiwzgZM
Xbice2GMvXTQSvptOedxetES84QG40nIWrJkKo+TfePn0yoglYJEOlZz7Yo44198
uCP2CbR1EgBToWtCc2kye41eL6NWGnLtANKAEHvj0aCquqsitt2u7olWMH490yg8
51QehcH95A2JluaTI6aflZuXGq8smjT8lWFQDHIiuUKvjXYI6aUI//J9V3z+RIWF
f0zUvGr2Cgm9bj4t6H8/b9/dreHCv/oTRfc3a+fjlw43tTyPo2Tiqxl4lJQ6I6Uh
x9VUsEl1e0SVal9DY+VSbVX8IfiAorc2GMDiDnx0EFIsSreHPcV8O6PyD4V5JEK1
4skGvahevOjXrYxyKIO2feilnlepZeJ1jTjdVmK2UT8cJVao4W2dDd8MihS9k5cq
YJM6fBz6nTy+FAvip9/eB4abdyYrtgM6v3jd4t+nllQl7udJoetPVlTpG2Yy262H
`protect END_PROTECTED
