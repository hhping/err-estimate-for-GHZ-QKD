`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29N+GA4bqkU1FqHzbfmZqUu4KeloFRHQI9Kn7OLQ3Bn2hUMYphToHQEoB7SHY0hg
C4/l+VLoQj/p+/A0+YXq6nRobsNzUwuZBeeQWk+CafbtwrlJJmU9esFPEp1fEVye
lxR23TnKkHzsemqYiSUrRWkccOMtfCxwwe5oDAbdwVr5oS+4MNfvFzfOvSzI2W7c
5W1VVQqHCJnJABDzadQgUYqlGm8a2YP4T+RDpCSrdgVAW7A3ugxFM8qNuEVpbKmw
T/lIC6iJedjCC5kcz3YSxaAKj1xVS/lqG0T0EMJkmreklRlmEQDDJn6FQbef8eOV
SNT8/lDk2BQEVGj82ONxV8wkB5XwDdXKo71j3ahHyAsScLZ9gKNUlCWF4amaTgfA
N/rEik7xpFBwL+lhCcXeZ1X2Oz5r02ff1MPrAcYdsulPE3Qrc0aAc+qjHAWPmS6Y
cZ9pweKfSI4vqL7zyxz3r8O4JEFjvRqQK72yG14s1GUXRuivL6CqdZQY9EpZ1rvM
DQP/TLbnVLetXquduKuD2ppBl6gwWgbhtyd7j7pyiO4vDJac7Mu/pbdXvaJlfd7j
/76EHRvntql1tUY5jqEYHQSNxLLZF3S+29H5cuBNf1SitNEj2KpQScj7FId/bMm6
lePLcjqF0LLEXF283W3qq/1Pdg9tX6F3rxdNtNuGZP88G2xF4DbvpOjkXU26p340
vCGI5Scwkyr/833Q5/THXjXimoLj0GLDCNYgwQtiv62TBzxWnsVQduQCAgUSNV8T
8aA+j2DyyHlZS0vcMVyhU8q6SXMPsere/8KL17QssmjXdOQib9GSiU3N8Ht02jQ2
JWqb834ZEgmjH/xkSjAVvlqe0fEtIEKrxo4kE8UYyrS4V3ZPLoi4VlxWwez8LyFD
DIbGribnglSd0E3Oyva/U0dOB5HL75O8HVoGaPB38iGw3wEt+TlBgBWDqs6w70VN
aG9RSMwoj+EZMuokexRGf4dffU1Sp87BdcfO3KEGXCrMfftQnYBIHYv1t7NUxz3q
3IRW2O+RODCCJVZoDMOwZQeH5gmXvs8uM//X72OFxMbex5pQKAsbwwT4VeM+Iczi
tQUrsgf8ZF+KnCV/eU+CMiyF6dPmoN80pInWAGdgGaCIRyeawUqHcYcGiKTfToCV
a4IHSQWwdTDM+mQ5O89iwQkHXIHQDs8A8lqLYYXifUTXie3Go0VBTH5yEdMaKx9V
H3S1ws/QiG3FWBP4H9v8Ib+BY383sh4ekmPJrnf9QLffYZNzrxKZH9JE4jUogT2H
1CWn0BVzaOXuES9mp16bVw0rdevkd7cAsOHNZbKcd0tWV4MD+xGfNNThyf4Wsm4k
mZGAAomZs7cl8v/Gjf9eafWBGL/B0mhRUvUMtGaKcCTtBl3Je5GWeUCd13NsPF76
zHNtc0N0IuTeebw3qfbYTEpQWTR2DzK3l8qTwfUFy810AHfF57+9+gei9voNfi3r
GmTWae5oVYcoZprplosS67QN9sWZc6vDHWB+9a7amGggqN7mR1grkunlaHmEinlV
TN3ZZEw+12/TcaweFOgkgsmMIIaQlQJJaJZrBrAjfdvFE3nzSifm2tHGwRMX/H/G
/hg07IIIhoO3iFJyhZXB3sT7aQHIShpZSBuQ3xE4k0Tb5UzWzDt/4VqqHrVRa8w+
5cjXQukpNOScF582EOb7aeHcapVxO8CN97ZzlDY0LnkxAHFqhRkMJtepOramHzxd
C9D3F/xeDio9jBBWzSZcp92Ycyp9lih9kW5PyFx0yY+5tEoKt61qwg72vowGSp8s
MpdX23Qf6Kl9bbV0d/UYto+shIJtyqZcAhIigzpPUThx4pP5FmTc5oWC6jpo4Q9K
dVuv+ICyLc9Yrsu0Inkwu7RetW/tzVIRzs+LKg/8gJtcN41+LU70CwLNagRN8lCH
1ZYPLeDHc8SaOvwrrO3wL1BONU1SaTWSPkgNRG+DYQ8yW09CUQPaBp7KyMxWeChH
31RY2byjFbdXHBw6s6GDdIHtBkVNr3eO8ATNjT2/5TXiY7VNNLsfUmSWpHtfKWaZ
I3HFHOdAvj32vlA1BqLrs/E5SInNieGZIkNep3VvPeMVmKLkeAcZ3NhMDvcFClbR
g20yX41/XKr7ab+oKQBO5tujEzpgkjnAKmhXIBjj37t0fvws0V7YPzSL3WORUl/w
XH7mz+HGc4zXkyzVF+8uDwG5CfPYhv8ADg6wX527cJjDYIjLdcA768VLg8z3UKNd
nucgIVRCeXpDVCOKIboLbkGm/ZaYpUFpdYvUr880JUDTy+JOLBD7HJib06HT3kev
ddDgWc1meLpTaQWivW72AB1WaYslqPBsz+R5VLmYUHDWKCxSwFQXCHyalPrZMp1t
ZAdpMF0hX/FvZh12+zT6z94CaGn+FNts6SvjPP+givaVdwhS/DvoMGdDZXsa4Bng
nhgwCBntMND+7qxvx9dPJyH0pWam51vNIvZ1WuOI5NqG/8kg0/rPD0YmsEFFFOnn
C908lYgjUxUNQhdu8nqgrfAbDef91q4DQ8sf7BaAixsBMvfjeDtr5EzqNC8pJ9DB
btjygnJ2NE8N9OEB2EH5ZGxj4u9Pi/Ck6wtTTiBZ6brJysrho17g4r1ccHAPXCeA
izkTa6IrmBZiEk//RsNRPwBv4TvvVrIZk+Z8oSgPkWrxYoa2AmN1rOw4831CpxK2
kPswoyxubcDbg02WSfh5Hf258T0TgciyknCrLiu0fJ4xjHxbsFWYZvig1RUtB70Z
tYdRCF3/b0Cz3rVM0jIwkoBVUKDQqiiicmF9hhtKXCrkAlxkxXqc3BTqG8VDpr7N
jynyaKNDG4sVJSdOy8DVW8PvvKnkAYRtESlL2OAYkwWsjB3qVXZ4GFUVTmnaa1g1
lNyypxK2EaNnS6BuBk9A8MCBJ2TT3XOfPxOUNA8iK7/MJ7o8j8wK9WOofnZGYFuL
EiecQ7VkJ4nkpZD6PNaH7yEo00wpdN936UahfR7AxU8oX/lp1oGFQeDguemhosb6
t1wzQL2JGhTveBgpZV/LXiabRsLw0M4FMpJ7VNIC7A0cezf8lRF14+Zm0vs2KeSU
TPgmg0dyvIYdTZyL7LlbnZkZhXJlo27b1z1x9dLawmMS3Z2DHrKUSN4fHjYshkko
iUgB8jK0OyvEjDBNdaCR1bIkiDpA8pzUxW8fnArmtiQ+PDbbGMdIbJh8LMqgkV3H
S1J82ya1abXgj3b4SfwsOcURaP47JTAAQ6N0MNPwZXbkpui3Ub6dG7Nu7yHSUwur
pyJorSNfkGavgaXJBhzOOnp04hhD6Sf4y+udW8eG99SM9EZwZYVjbKXQkljeqhDd
wHhTW4sG/QKbXoUvFxKHRPip4iQ+c/ldyzlTG2S3vgLdm4keYNOxjDdtsyWWi2vH
`protect END_PROTECTED
