`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cedqgynZOMljTXvE0WluIczCqo+v5mz9rxa0RcNopXMJdvESnMccdrAfI/hrEvhW
PKJmihhAPTKyqhmxCrE0pWGyAUX8VmX1PfgJBdj6P0lLw3eenGVifmGdBu0UPljI
ilNpFPVL22c0qCbaYlV1Mxejt0XWSYe13OFSqsfyDGNOE+MSs6WdklOoWXE2w4aC
lpCT550gLwVVyp5tO4X/gebuY0NuwPBy5D0A5lT7P6yjtwO4DF96kGBmQs5oaNux
B1CJ9PlRXJrU0XJq4M4moa5ZyEO7eihODblc5J24zBCNWEAEGcPAYMjzBaxcqaim
RE7iyCjRYE8bKLAJB42fA/THqNCXw2srydZ2wCqu3vlIO4znPBng23FN1S58WnmY
juLBhOas4x1LLl56sDRDw6Y4DESD5iatrhSh31ScReZaASgrdSSbTFmHrVAHQkTx
HBnPFfcDca4Aatajn9bq9JVRIRgd3NRSl5EvzTxDt8YhvSOa0enC6L9IGO0+xpXN
7NCyur54OQRJgJ0vqurv0ncEHHyUBdmuqtE7pt4QyYa68vPkEiVN/uKNbM7Axg2T
1SI8EE6TDFi6QWIOmSccY7vo92A0WjwHrL2qBAEuHir9K6n2y5VMaZ7qy1sEuELi
GtTm4LWdDC0bYG1zXecQk43Ec0vxFgL5xb4D9s+Oz2w5vWOpNiI7PqXyzVz6Lep3
uNoGPBnCpvtAJdPrmJmy/wcsA/gRoqgFzAHmh6GYGv1ww8FrWtQXm/0g+RtQlXaq
cdfqnX+IYnz7vIb3Kj9pJsUYiVOPGQzlM+jR2TpxoMEFpQp9uU4dSDyzCEzQb+MK
F3fpFfNRNpL/4uie8Waj9g==
`protect END_PROTECTED
