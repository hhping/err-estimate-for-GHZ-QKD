`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmFZyRT2nd6WGzJ4UNr3g8yFahEWqPM4YA9JT+O4iyJbjvJCdWyQn/t22RGQ94Ee
NukNQUzCMPqgq5HhydaYIsNQzf2VvH0rpkqpVLc13jaXTdp0DdMo8jM3aEhutrGT
Xctbk5CKYP036XFdo8q9K+H6WOhETQlhRq2Zz7ddMVx5CsJwTSNnqcEqOyl81KEL
cDOCCXOIClsWoiPryexdhgAtFfT2oIMsdPDuhfG/faK46JMqdkCOYqOEyqdvioVz
C9lofFY8iEi2hAtT+8okMzSf67QUaQYmISKRL3v5ooENUKRWebm0q9vbHmemE3+h
/RkmySleMWMeD2WnPLgcI07eXDbfzaepIgP+xYHB1dKc7DsGccsNIDLLZbKOfG3u
JZTLZI/8DbKiZMmqwzOY8Rldh10GPOqcyyvb8y1es1Agi2K4v65DHSqlHC5Yjug2
F/xWLQ11pdqUp0U4R2R0HjY2F/u7lwgjmQXhQX2ZYCuYMevzPM4dEu3ZvteTzvQY
jrwLFiq7Pt6JtHJgA3uIrQOuKKvRl2QjV9f9z/f4IwZuhSXWpuVNFUB9sJ3maceq
vuxr/dNZqOnd+X6SpfZRzX2ovemEbvKzK/vZQbIaqK1qqZF4USX+95yEez1oSbgT
ZjkvwFVnrKTyLKn4peoY45yzrAECyKoF1lx8vnLzXy+EiYdv9NNnxRUzmNVLd+2l
YAa/jIvwSWr1FW/cXyrbnO0O4d8aAFJ3K1qo1bEeJSGHyAdQvo1ESL2ivAYerAkY
OqI3fdXQUr/fRlma1PPnRkavKZJBGsPDXo9dCf2WWLOw6G15MjmXFF66H0cLdC2B
fdcn9akDIj4Shy9/gUadWzWmcbsb1XvaJvpCdWFopJJcEohzTjeC2i4EDACZ5Tpy
n54lPbUIPTVyMdVH91fezcltrr4BfTexWQlV0VyH7LsYrCRnLV99AzlKZu/H1GnL
UJBws7lh1D228BvJaG7AoxDYFvw9JVgCqUbKd1GZ/knpO9VOknBjT0u7S4D/kPNG
1G7MG96mDa2UTgYK5SJ87Yrd/l5y48xwwjIHHFQF85cAN+zOdIiMPnPdMGsCzDjS
`protect END_PROTECTED
