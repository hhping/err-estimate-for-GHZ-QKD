`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qLXP6pdqAEIzfFBbKuj/kRTMNa459Hiemss7gOe5g3q2iS7H2ZvmU6lzKxWmdV6
d/PWbrVNLYgApsmNz88lFsH1dmUEAJQR4b7DVAKwNGRlyNvuF802iMuV1K1F3SSo
eqkVl3c1NZtVEdb2Tf3XitF+Mf16eKQe1/A2xsFp6dGb9r65J0Q2Rof50QSogOCh
lVQu6j5z1kGo3iRUc+qWgYH221mpieClHLCbMssbDSv9JqVY6UvTdaDPWGuftXeD
hynUEWJPHVZRVtJsrtSvmNTkRSHlgKI5ors0tLPVr2ETZnLJdaOXw/C762nc4VR7
NdFOnGpXmIb6VLw6lU/HooD2efrek/7qO1J10Z+Vg7qTqD0VbsuI8IrjDJ30NNPn
PQgzFdjX59NmoEVpmWVeuKjlPM4FtoUbE5oWjRlKqbU+/JR3AzeM6exT5XdrE4eV
vkyJc8F3bEdE2r6IEPAPLngiHvfy4jqyC/cGgPRHKROTTIFDWe3/rzpJqtNKuGk7
YBshzG5UBK1soI3l2iDGfPRKtPkkTq+E/LeD81GfU6uh3CJg7NIY6ER2dvNEw0qv
gQ67JKV/3VWhopSH6fQth/CbwiXzqY1m+86W3jtw5Nbj+f0/s424u5cjndLltfAO
zmPsaGEagUBPE6wdAnmje9p/HIgzn2ypMrbX1CgiwsCg188K1lVXGklkAtLxt4j2
VD7E2LY3A9U8vF2O02ZBmvmfq57NmP/MaMC04s0rxJbpDgr+WXxtPRgZOAzAZX/X
VtgtXOlR8hpL64BtIIQGS0LAjiaV1YOegF8Tl8eFwrS5w20w4I2d+yayk4t+ICYJ
OLYF6LcjfDwXJfQ3vFi4fKZk1xhRNTPu5xNl4nH1UYudGZRQJyGkpk8aM3fE1TOj
wq2W+xmgd/2CDWsaSxs9lofoqF4taExrn3ZhsikCfaQ7VlmYtc1eTQ8LUo9quzq1
fRl69y+Jk1rNx1/D08cacNytGXFV9M0xOad4S/B59iQKjGb+dXkfWELikICl6RTU
vFUEcp0ozomBgue3wDIt9haOA362f61L4AieTj8403aLfK1sNohN3lDOIHcTAs2k
T9GmnUjBkRcKx1YHYN8ebMa1oXQ1KNBoLUtj60Nikx8KsP/U2eDG6InI5zVIWyDH
GFLlbIiq89qgBSwjw9OTZMazBIMDB6zO2KYBh853Zalirl1M+rVzDgUuchF/+7fS
T1KdS4sP874fnS+sH++RHXl0y9b4sFlM6S2DjT6ijSxZZJmf7z/SO+GY76RWGI7t
5OJgYPQ6E+ZpETpUEHtfNhyy3oYsiexjbwEM5vohAIEtQWKlUUt2dxZSMoNRHTZi
zX7SdL5PSprBinAJmaiS9XOm4jt9lcia1uK+dLaQu/PnHroGsvx38QUdWdpnwQBs
HPdEhV6qPurT74F2aCjHwsqgaEJlEkXsLrfAlje6riv6kzkWksw0r97yqA3uhM0c
oUx7E7vsdd0/6CfcaI3Up2KC1RiJRm8RXMTDbMCbjluMzXgYsvNGmLzOl/4AsWJe
WBN51QQnorLpkn0Ym6AdO5KMQR9Di5Lhu44RDBiuus3qmzGMvlXug+27ARq8OSxI
qo8t6Nskhf75ng8nQiV4Q+FjJ/5hIqOfjtkQu2xVyxir6Qim/77R3nNMTFM3x1gC
QPR4yhuFkcDa90ENJ57R+dpXvTlSRdnlNBwK1yHXrbCg4k3wyVr6z8xC8H2v4+Ms
wxyij5yvf6n2EaJ26oylWlbya2kWB4tfvlykxfanFrbZOBHYgmyOoO7NaVmdCAAz
DCrtmFCC3SmWetaMW4LsnqTXV/5pYkjdrDdkGf6qDJ1a7cEVBKsVPWm5qlu5Sfvu
6tvbuYmO35XPHG67DUmivsSCgEpeGOJrnil8FuY5VlwoyPI2Y1tIbv7GoaKjETas
i3rLY1SCb7djeI7JjpvBzZYPinKuIGZYYNTbyWGhE1p8x7IQwlrxgm7KxwAQ+08s
rF9dJhwkh0i8ZCxagInj/2nChLSaGqyjTsbkcqdT+N1NJFPXY9WG/YhEDSXwPygy
pMsQmxYL0iiy2gHrmXrI+18WVL8NGkz44fpv26+UmMFo+2vpR13v7liJ58E7tu10
SqTCD03yi7iC55AcuhmiEUHVJYE4LQJlsZDg6LQ6L8krKfMa0AWKe4Zp+UzLZb3s
6UfKl6Fmzqk9p5C38QT55IxfQCCFWAb3J4+TRMcTAfSHwO4n3CC82d8mT+ikds60
LwTI1RzUwrCbtf0PSLMrD2EMMwNrXVgksr/Tk6/7Xl1ErjA0cSVwHxPzYrvQYqbN
95HUurrYrCBAFHqW8VZMMjehzFxpm+oZuAawJgkyg0oZr1Gxfc+kzmym70R1WDzw
09Vm6/fj1bPo0nKy9ulxsUMj6wSQ1wX79nK/kfEp04r2gist+SVPHvEx5GUDpjod
Wf4ooHGUGihsgfAA8LqoYRxMo7adnQ5hLVlNjt4B+Tf0L1yAVQ/cBhEzSOQUlMvq
12zQLHwjtf0DVd8e4VFddEpShBiuqT9cinlrezlDhmZ6Rd6H7MZyJBz6xNfKHZBb
Ofn9ROOiuWAE2p7al7hsAmLkqvRvImaqhubfkOxz/PDOuBeOj8WZqzq5GQZmZkjj
ZZ4mtsSbvJFHHjAkOg3bcB3aevX+UCw4wrImS8rKe3tcJ71FV57GA1s8doRVeEhS
P5Qw3lKEJzT1Z+vivddCkHZkUMNahWFcBJidPGfwoZMVX0OmcLtjBCMHARrX7ZdR
0YLzTtDfHxxQj9Bkp1dBg3wqVzme24mL7YQ2HzdlHQvYJW6U7+7IBVbkQP284pvN
1VpmALr86/vwwHyFFg3kR8D4Uagge1x+xZkQzAdTQtTDKCFHUIt+OuvoaSNoiXZv
AdYZ06o8dNmw7f6U0hoLQWqloHzToIxHgLAoea9gcyZEIaL/u7mEo9PXXU1/Lp8P
2Ju45b5xsmbj/G3fHuJHdpXpC+qwIlFvRSyBBqoXAnyEQJ4UMABajA1RslD89sz7
8LmqnjN14K6Uu3mn92S87b+1keICopFpYrTz8y8Sida+uDKV/aHGnaLNxkGrXQAL
oJ6Dfzl+NrQ1JvpZpsN6JvOHv2DdYr1+v+vHU+wfe5Tpfi+Hy3BGv5ULRPdtdQMW
QftDetYAlsjUQgEuV/rJol8f7dDxIDcQNuQt5pN5/q98+n2aM7T0PkRNpAW/jEzL
wduIHG9+hl1jVftNIcVmR422XfDvdRUWd/WsfpDyyH37ELO24UmnwFDS0SpJkNng
9ajNxz11tOKbcoUGX85kxiVz+ThV1fuB2vnNf/80w0cQrFHvSmHlmCFRkzZpmxyk
5V7tyD+Vlko9FfPqacTz6EeZg8Exb4ydML4C3qFb+Y9eXrFZ7pTMPxijtlW2+9Xc
Pslx7WI5cgGv27THiKq6iH2P7X1JORNlCs2x+3/DMbHK7d5aZvA+FB/a69MebTB/
NxkOuac+Qt2BKBYfT7aD9KsVirUKp+Zlz2cj/E+S7LOhCA8nMyyXvdV/kWThxoaq
4/CYQPWCa2G3ST6riRGaOq3EVgyOd8wwNZCB9XFOm2t+tLJ6rj7UwGdnGylWQDND
D5+5iNuh878ZE0/ScgB4wj+9BmY69BHVCeI2HaW1EOP463vfKPScfQRuPMoe2RTU
eRRSeluVUZjcfgt/asc3cK0x1B1RdQp04bpAStfld1yDRnASzELEmP7v6XUBn1Zc
GLL/NHPlu4z5noKYwRURl9hXLV8i7KvIFBRyz+FDyC4oj+gwwvXONnZNRkfHOzfX
5jgbmd8Dtarsd0QmOraIIJqlbVsPEK458lDxVPs70YHE8sqLjjM1Hw+a2hC80arf
T3t45U4LILVTEQl0t2rKhya8wEUtQOa4slKU6EIVsLdWu1gnLezFVESp4GgJ663R
7Jn3NdIIHjFt9W36mphk6cs8M4B3mNpEthrQIaDPJ249jQutOoxE33s6md8FX2jF
`protect END_PROTECTED
