`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgFp5dRjCYC6pPMbz119gUFgdI5MADB/Xw7F6j95ZEkdMTYH6fwXG0J3JAOlU/gl
DU+JrhQchMHqpasLhzLqPitjjqzzfunWgXogGtC1+Y4slN9rXDiRXU/BbzhpJuJQ
kPoXNLO0DHgfRNOw3oc6qUNhbFDa6wqf5ElGdkdlEDRlsFdgP5b0vSlL5ZiJGRtt
JRgt4iXjyg0nQfAmPuDF1CaCf3ZN/hI8pojbmtwiXUaBsAC6rCgELRZrAgGiQejW
Ph4s5s0KPBs0Cw4Gjq9FqM6R7tSh/SPo7EetAgA0cf9rgNoWm8FpO6+w9uyxFME1
JWJIWy+ohyc2owULEJvQVSME2ZfYckc7IQ0YVvXl8fTSBbyTPJho1XMSBHYV0bTk
pCcCOGV36qEbz8BMzmsIadhgCA93+bTD1Cqr34/5ZA+GfS51z8nWIvjLytt9AOLl
h9bT2lIlSRRt7021IwZdyRrtPOtHLmNvQM2UV0OHZVhS72BFWNjklzTKB44nFAIR
LFEl0pMwPJvEk+LR6GzvNrSDZdA26ecNkdi+EvZ9VKTEwz7EqAb7YsT5Byk+gBzR
z4WFkQLkQpw43l+mgBktzGJEhHofGKefJ1oXB6y9NYHb/WqATIP9ovxvBtSfSMVW
8tFbfXViM54EIL9+EJfPl/yJPNEtBSrcQcnbaodpeOxkeszDCXuHEH/J9JFVQyb8
So592Q24DB7/TYB7GEekBwWBjYeVVqGJu9QeUS4b//3r9SLOIqSScvTJ5Zv3ZvlT
3ZjBVYbU3ajMOemhq4ezZfb180hFBRPY8AuhIjjghYcXqS7gxoD5fj0ZA9GmuyLp
W8VAVBd3TSibw0jxCb0zj+3HsLvx4eL5sIdDgKp3KQffKUaR4urEwkImyP6Fpeb/
Q3bTwMzeee734MszQayTsJ4WCslxstaxiuuDoYli34Uz3rKOEadhEDyxKuHJphQ3
qY8CfQsd13E4PC285GA5UJxPaV4gwsQEdQfSbmgp6NIgl4AmWFDMPSn9wiLV8UOm
dIErW4YpdrcVD+T8RaY9qBdnyyYyap6OSL1t/uiW1JBBELSWjATD17x7aDj8zzcB
JuiXbuXYyOIQCuASP8c4VX4dTop4QmmkxBxfNKFq2ZWJ/a1esRz+bjNnaUXrKVdX
yvELjOiRF0zvBfLPrUkJYCVZb6hSaJn6EmwlaDWAn0YPdTAuYdZHrmS4T+HGo6+H
q1b0CPmS10cyIttSgbyo9YS4idrDUWBmwEu8HMPXOFvVLUY6eSCitcFdVj43UfxC
Agux0XbZrYADlbmuvNFXbgCKEfIBnJhIhhwyDa8hcYOxYyp9UhbqQM7sPU9LXemE
kcHz+3ifqjgO0RLfNo1rhwEF0a0udTB/7ytDoxqtjHYn57CnikK0kMW4W16vVw4a
MXzqWlgV9YRqu8vk0D50nDJx1hl+iY6Rvio75AV1/t8xpgLGR/i6k3Af+ZQ23Z6f
mZjs25BKbJp7xi4Rf474vO/qRkdt/N86VuWmpeZ2JavgpwkkV+dHWTI00bNji8l+
TCkWK2YtFyxaWX0jGy9GLmLWfHUm913PY1ESILrRaqiP/wVzbSB9HEwzTzXo6lh2
YD3TGYya0CTzaA/Q8njSh0qVEiWdKOqnTAwtBCT1iiNhsw48GWsOaYL6ZKhvHJ7Y
`protect END_PROTECTED
