`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UqguHK5diKptfQktwj6Bqr4NAem6thP0UQ7PsquLlzXtj4JJcuXd9iR+WJMuNug4
OML7KnFrX6fmnYax7ij+gKI4D/aEGXtYFKW3ESIQYA1Nu+MqZ65muYSXfjh9xJLh
mnF0JVEpJVvgosjOTRMXm+2ZQh3Iu59jFeisLrEwSyfRQfEIAKhks/nTPhaLlH71
VX+S/8Olho2j4Si/hu1RESVS1fRYaCK0Aua1pY4/0Lz62snIh/Kj1tvR1bAoDVn7
S7xO5wfnpIdPyS/LF14nBc61fs9Z6EHQDlhgEe2CmCTsMUoH3DiA+OWd2kOXyNV9
1gryja+4AG3tBecXxJSSvuOgXu+JPz2AzX5VxFYPdDrz0OMwrW0Z2u9ostMrRi58
fvUdAfymWiEdjV/Jz+ydmVqguY2KXBZ03jGIWCe4o5tEWU27jLLldLCXOuoB6DaA
McZzNtfMLzo/7PjWmBx9NzjzbM37I9QPTv3A9b9+exXv6p91nI4c6JkDAfsTrYkU
q29928pRLNwNoS11HXTsWN0z6vROQW1jwB+lHp3IK1YKqSrrvzP1ByxnEk/GPZ2o
W4IlzsqY6AwFlDMRBWnxLR0uk73gCpARed4zq0WDjUoAEdcDBi3OrVGNNGVNmOM4
gLgaOOHK56420u5w+8+jmjNT/H/JtK/aI14ZWE/e75E=
`protect END_PROTECTED
