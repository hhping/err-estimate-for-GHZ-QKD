`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/NsdVNGRuU7EeKCHzkfqZDD1Tc6FQJSxrwQdIZ9oNs0yaHyxvNIz45mf68AlpkR
vSxrc1npywx2aNMHBD0k1/wHNuFuVwkvTHKq13WsJglCw+XIxoQp57B6Moa88hdV
RYxbkC2Iz+X9PirElq91Ue70+SzPwcTn87jN14Is+Jizf1XoEpe7kZAIDW375eBI
IkcuG73wZj1agSgythsHv61yMpCX2zPCflvl1iaVYYu4KLBVbDffIzAJsJU2YhTo
FEOJfVWsYsoCXfnuYDu19nTDjO1gqANlcIBJX2ELpgdsbzPMEw3cjzOPM4uDKKtw
DXoVIsskm45B8C5KlUMiq45BLuu1Ga/E/aW2cWLN8PgeSlVO5jZE7SzdHJuBwHQM
9+5YZxOwD0XH/kyGuGPq5mShTJ6DEcQMgC7ikJhBeamRft04LF/Ks0mWS3BFcQON
MpQJuyFN3KqgKIsX38bN6qniIlJk1MRfU1NMhZ/2u+0Im6gm30zuLuZLunQJk+6m
xzz7Zoh1s5aeKTDOaMfSa1wcWohJI0U+96qLmR8VxQw=
`protect END_PROTECTED
