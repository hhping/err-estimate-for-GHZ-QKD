`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3GMo9zlIsGU/uRuR5A961pCM8HP6wVeQUscTtesxHhhIePyJVGmLb6qqQfkNJtjL
xMeyZAUAFRWl/NkKAmP/yDfmImc0j8LJ7QFr1JGEN/YTWxwJB7oNF8x14KVHXTl7
w+JvKYKPAweVzhiGrsKzqbZv0a59QF4nvJoOn21BIglnl1BeftkSYjDSfOb9URMY
gLbCGu8OFMOChFbkeCllYdC+D1kPc2+gs/XOEKlAlEwlCxaGQX5U0sfUMWYsP7mc
IP5SCIRwx5a5yuQULnD1cS7iNmKDsStEZ0RRCGq39WnBIBlzLWypUudQcnoRFN07
Zy8SCCOW8ylGMQpjDPuL9h3aly61yJFpLTFBngiZebPqMhi0xrrdS3Ldhe1ItTZY
VM+zqs4HU+iH0G839TmyF0vHSFATzHVjX8LpQEOgTGtez1Cbfc3F0694Y0wN7/D+
ygjrH0TERjUaHRFLxJo4Qu38U70Te6m20LhE7O5LhP4pdl6ZVMBXA+G9ESLsLpL2
OvnuyVPvLKCJfHi3Aqvp79UQWmDgTV827jsAWLt0aksfmtgcuNBzzC8cbrc1yHdR
q8djkg6vcBJtp5ADJ+yFKuDAZro3HCBKtDM0ON70Lku6VYtkA+m2N1JEKMsCijhU
bMCPDUX83ECeh2SrHPM8aBeArgoBIymRe6EASWPV7DwbuiyPEHR9OgDbx3rrJGil
GcV4poWLPduqQNBJEHD5ZQ==
`protect END_PROTECTED
