`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuqnbxWwyrG6xwrA9I34OLbiXXqR+hiAiLF3xum6RBiAhkiRV6ACPQgTLF9VbXbI
wUnt/hvd9oc9fCzCy57Af3Jl8E9xxu/JLlFGQWveVBJ9HZYbtxp9nEju6dBCBM7q
iQPtZ1pchn7DAud/Q/TfJzk+BnsZ8I/iQY+ZWkvIfHnUN7Whri+R1JMExeNuqYlu
Hqg//f3/M08iZHycmyjfG9P4dMWFlZbkUYz+GgV971IWftAEVhBXOh4ZmctLoc9I
CAE1VHsi2v5TYAhpG8KfuwPJloEfyLJLYSt4O8yrMNb3FljPCgk7SmEvBa6W9AJ4
MeD8PylIppWQlxtSGz0c/iquK/WqDoiwt8De03EEtGsc8Fny5lE8raayiH3PsWc+
sqPEVVlzhKtBSTn2ymQsbaWb39JCuQUSHc5x0F21z+vJYzp0jAVUVuhiEMmDGknY
h238RtV37ev4npBenQhKrpJSZwkcNhjtS62V06oEZYBABYrOOKvQ+pPgO932N6Ar
sUI5g9wSsfY8maF4PE5ISJgI2/pB+X9lHZA0gqr1cYn3L6O3f06MFxHogyiUMf11
GFp6Olq+PIJpKiCjb3zA7ow7cJNLE5KQ5pjIExacW33rsx8SOclAJXeDf5IrpkER
Dbl2ayE6pHubXSHv6W7zxrjzg4vsZpAEhWqQbXWZICJx6IWlqw/mdMVVycm/WnPC
2f/Anocdk8NzCVGas1KpL92k2uvujG2sVszCzra8Spa3gcwO2T+q3I0/u0lLJk2j
mXnOFuaO9LDiLhZIV4F2qw==
`protect END_PROTECTED
