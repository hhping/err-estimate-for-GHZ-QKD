`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DeSKyfe3eWtPR5WXmMq7BFR/e3vJvGN8Z8Yq8Nmc1Cdzn17xhkHawY5eP0YnJYp2
UosT/xPTKzXeUKygE7aeikCvpn4sQsOTFSh4opu+lYdXt/T1VRhcCnjnt1yya5ZS
i6U7aDpu8FYWwDW4tqFfk82UhFBDm1NbP0nGS5AFzyZMlIHwRG1i/vbD/WLxxQQV
0ATM4L+eCXpnemM00tMiwbQSe7h51uzF0Rx1/Wb4tWLDdBg1CS8lelTVHFMvWXXS
O2xlWQB4fBrRd4xDoPsu3BgTpjQcFc4YNCP6rt1IGDn4gupDcJTYWy1OI/hmrGau
J5lGxFCUfGPPuRc5S+rahS9GlJatyDbYVd7MLu8UPl3NQpXBJLVMpmRkuWsyazbC
tkm0qbY98wp1F7PJd9JCZZYSOvc2nQQ4kp2848g8XvRpwO2Q8tzNrQbW7/S5cIAP
TiBYFc6O3WphGrquB2b+HPcHI67TWmcpzd2kClcCOKeiKgx9MWQa2EWb3E8VihP/
jN820r9+McL/wXjteuelq3GhImtlN7p1WJTeDTV6osio1qvHYomnOdmLBqcml1OX
gYiR8xlRlxTws03jix/T1gLV9eQbiNq3UUgYp42pilQTM2aYxRovsVvxISV/kVX2
85fbisZKfJie5HzPPHs5PIEznuCGuz/tyAc19bFL4lpgqhcs/GfDlWUwWSyAwsPz
49zLA/dkgONXGYIlRLYctBe+nr2MWSfgqfLmESBnNAZKpRMYbkcdH++cyn7V6LAO
dMtimwJL93zVIzamKL/KHhvIRA5VDJfw4m4U/arBdH4KfyvhYvxjl8p3k7WGWadf
BcF+dKoTll6hTHEh5XJR3vYnG3GjwLnVkOf22GOLPZR2Li1iw1gG5C48UDWEPbts
HoTNq9crBverLvZ/4DSGoHK/C2A+DNwttksBDrdnW7nVhDVmicPd7kPH7hL07EWQ
KXwCce/4F8Wqm8wkH4CDk79nYLlg6ByvC8HMunuLx6edjXCfz5cytBUAUkd2pfiX
E8WgfSOwMge5uFBiSRIUalVnXfpu48NcMeEc+Z71mD2SXt/BWHQsqgm1Q39e41r6
W0SKXU/LIib8r40caJKyB0D9ZY7tHQybCtuVfzTXGNBcKyE/sMsDYIkDIK5L9DVo
IoZjoFBfYOnV2XSGtiSVli3E1J7fo4RUigfhFT7UnRpJdFGdgLzIaRIWhiDep0cR
tXekl9Y+8JdH8t4i4bHgtDW3S6ZRE7I568dSJJzqKxdeJoTC4l7lJN2b8HCLF1xJ
GVm9GK8T6vm6FEndSIhk0ptdaccZJJsDkba+8x4a7W/1Q1Xiuw9/03KA9dvFyVrj
/r55HqZ2symCYHsKOQbsx32BwDJvPEiaxsjkuscIkLXpc7Mp4mm8BII7cYIULwJt
pTcc2U/HLr+Su3R448VsD5kWyJ9UlCQ105/SiQl6DCGfpmKBrDq4BcofAyPTNrz0
ysdTpg7EmjcBnPwPl04I2jdRJSoFuzZ4EnCCcraO5Oor8MfmtiEOzG6ARSKmYwev
IBR8e0uCFMkpNXV19ci8THHqnqhPUdbHAB4ZbKgdzS61QPV78p80KlMfQrCmRGWq
TePcKNy/1bXyeMfD+YpemcGDC3TdhgN8/aDseQCULSPBhqYzKjK+wqGOJpj0BoK8
5Hj9Y6aLW0bTnA422G2LH3zviMj/Ib0FTC/bBH0IYX5wvGXFUQh/G++Bbxko20YH
yvdsozB8Ky8DDJ05I/vdtG2+78TtGL6E8CvRvEOezc+/A8BOOFc/gevIazavXJAj
2fCEoUxhI/ZWO4ue78/kK2mWYDiCbCyLLfDdEHV5xcPt+q/3u8E1lmZJ9VDciO6Y
CXs9sZsuLVvesikw8SbeDKkK8tXV7yjMtkUAMNqhrw6l3Eiy1SNPmGODUyhxkccX
c70KDrwPZTc8E6/lFd69hdbtInKUUWt5J26HRi+717s1zYemtJN36TD5kpkMmsoC
/hqdMIXBWP/syoH+rk/EVcDCLEWKhQx9cX5gnGdOBm9gsYFozG1Co6n975e9bLr9
7/ZkVJ9t4jEEJgoCNcZzvViydAckMrdwdim9+S8D4RhHduOxQ3YLOtr8jKOmEMAW
v5afI792sS/1daGqK9KnRXfIiQRvOSVD5B8l2nOiXqXv/7tkkpkWCN5fHYnJ9D0g
osSg5NmyFEn0xj+zjT4Y/LaLK+4C3qcJEAHbM9/FbumEPP12GmVQrY97U1wuyYEC
N8xF4nr+X0y/SnoMDZthdBVoiM0pz5TYldyhcTIiu5d5AnXcfNLXqgybdRSX6nlA
4lcud6WxBZYJGOfIrtJYiExjTswr6Pg6RnhQmPMXgrAKhGAS4BpPnFctSb5NIR7m
hE/lkajt+mCavANsdKSzTm30x9RFj9l1XChsCyZtRlT8f5GYT9sQyc3XtfBRfKO3
0gCMlPeWpBeGq+hAW27S8OMEiYWVlgVNjS+MEcqF8phxfh2/MGfRgr45gAIcHZAC
TZWaddAN3l7K5GO16fVIZuuTPsyY6oNq+PhKNyRadz03NJeXIOULT1O92KRAj5jP
xqRJqXaXKrTJl4KhkNkLiCzNWetWTYk1lmyr0uho7T5xBLlT8QB/WMWi2ftye6Wj
ErANUXt64KLD1QYQm09HdDFE15Np/Dry0VOWcNStkW1cc3RLlp0nFevb8F3QFQm1
O8ST4PNxqfgzDNlGkDshVn9Mqx3WiMYWRIA2z1zq2K0=
`protect END_PROTECTED
