`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vBtWExciKwOfT3XR95sWOQg5obtQ4N/TiFsM/UyqytSuaj61NoGqFmFM4xcwsVj
V319v5d1EzREZ9tuLpUJDPG4LmiYTpqJ+mbE4FeUyXSNqByvWITNom0JlB+TSd72
sG3o1AA6BIzjyHDbLuCA06uJ+BYeN6abFh8aKtpNORj+Tp4KcqIaKiEeOxgahPUs
4HFVWAZXOqa5R1Iig9LLmgpRyedUGg2fiNVZvOmjQOQl3Vy39JenIXdUT6FO96b3
Fvl68iS7QYauQJM+7HYwHYsyuZrQj2fjv9recUrF9qXeNv9t7ORJfBB2hnsbyYNx
owbhRkV6E1OSUcKLuEStHBCJtn/lPKXUQQzNIuCvL4k7renxfdZy9oDIsmyfM+is
eXRsv7GlL1yCrzmUUOmU0fJCF69JDbEMTLyMEgNs/TotHqc9WPVi+Vr9o7u8vNA/
BkntNfdF4gtYFYPf9RGCLR35kjWpdo/AXISWFl2U5Q/iFmvcpWWG/wJcTLZFrKWe
ZFCG8rnFeW+KntR7ahJkzoMW+BO3uf2EHyS3UFVVwXrWPUlBgsOpA2GBkJ6s82UN
lHKGWydsoYizfPlCefGpRpLX+cTyzNl2FgGXo34r9/LtSZK2A0honJhG4arKYog2
+8ddm6awHk4VAsi3UEhcoZrDQq1t9WQojiSPIHrxPL+zzlYifyh7CkMP5F7/M14O
0VZthEm2i3V0mgDIfPzPMqadNUl8WssAtjM4nrxge2zzLjYi7UoKObL6By/3la58
GxgfnDejnBQhuyENccaaJ8US/s+5SvvYVoojhmP9JZdICf9XE/c8GrimJqVXLR2G
2rBiBSQM7jhfJ863R1u4w6oF5ksUP1cMTJLILoHqjdZYqnR3sVACH/9z18j4xCyL
vRaySElAqh6qum1cGPnPEg==
`protect END_PROTECTED
