`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqXtp4L/UtRrVa1DgmFltOPSwC3cKY0l9qgWtqTjOOB+rHk1qoRzTGQbnCEtelCf
juaPBvJjfGQ8HTU2pIgz9kbFDDjqPBCo+JzIPKlk/fvk/jQnF7nctkS93/wP248z
mqcyulolZp+cNXV26WjX7XHw1LNuTdvKMfoNpZ1e93JKX3Pz9wTwSU8J+CEtHDFo
vNLzditN2Cw4Wk5hvbxJjIAa/Ub4ynV1cirNinOahN+CP33WSjABiiweIShZSM8U
oqBXZDqrK5Vs116pFO5EyZoq8U/3eduyz1j/dLcufCisjhgEL06cqCYq0NIeYfxm
BMd2drCsJQe87iw1ioG6i22w/V2x03A/0nGR8MphAzqmcFceiNERvv7zXtlNMlFt
15sN/5dRDdKZdpcwvvtgVUtU8IF094K+INHChJI7SF3wVvftuojCd2T89OR4lLQN
788XZTKhb6Khli4oWBedm+zRn0W4b1v9HYX0nAZJi+d2KIivZhz2GVzOFMsuPR5U
uJHowVji0ZsnQNQTHAGe3tLlkCaC/OC9bQoj1RyVCeAaNVn/ApNebR0z5FboKRy8
MJuwAhX392J4ZqHQPw0pVufKLk4PLf245VUdwHr6VSbpjOdpajDoukNjDKW1s8PY
etJYAil286GRTRkJJ6Ir5F4QDgbY5v/YjIhuvm3k+yxuIkwpUFyaINj+kLm+eWj5
r0PV1gE9Yak5EpjojBcJkXzMkJVqhY/BjjqCbg+TmCsmgSPSKNLyWRTXP1/DjPEB
LVuQnU2ffb3xdX5kkIuFNl2GrwiBHd3WYRSu1TlM+QmDtJ81CiDrZFA+vEAJNYYc
qbu+D5c6oq1Hy8yWutclmtBBJfgeIlUdT2TZpMp3ITA70nfU7qLnRhkxtrGyXUau
sCF49rZQoZdKMA+MrsjmOYA2gt35T7e1ot55FPRmDkSDOemlWHnOKTbfLU3WvWKy
7vHNqebUllUb3NCaNd0DxFaheUB1hyTDG4F5jPoRMK+pawYrqdcxp+7L0dwABnnK
XY5UWyrpN39KHC1TE7h5IPao6AqC7ukzrurL4SDgkPRYVUONONLWvWbSva841OqZ
i/YnDXzHaMLVqNqkKRFS09AbaT8ICCS+C9/bWpGtATj6SWeeH4uiox6XQ6MbjcEO
ZszJm1LePheaqd3CmvN20jSsRfdbg9xy/ANY9V+RvpJwZqvYe8Rz8azmpPbMB+47
SnK84c8cWWCoiMJbO/gcElbQ4HXjYtYsBawFABVPGwhpHd0fAul/+LC8lRR42gYD
f6lDCJc2q9aiQAYeWlw1ll7d5Okd038GhFmd/9gM2jMYsNIcxPR5JsE9F4v4YK46
jadikMzfkP3aAy92yGD0hhespkR7LmE594WX+jbDjX6LdAdjGHhYFAb9hVBE1jKa
kekWX4+ScLnP243WuSptK6hgdW3YH4K1C4jlH4UE+naT3m3rXm/HdfkGx+kacASu
W+tsbR4SDx7FYaTpXnTBBDvWc+vFg8Cw3S+R5nKFMxr4TscgTVg0F6e84pBaC6kO
ISjfdoiKUWU1w82O668WE+cBAAQTNCamns/G3bymw8lCxIAfzp/fybkg7DwdUrsr
zMXmxYWxAwJafswG3awv7gFQMsFzsDpjMLv8OmwnKLwJ2lAZYSCX/pJDSrr7pyl+
iMw4eURu3V7oKGEpUjtXatoiZcs1vNYGs134sdn9ckIlcIq+uqThN7f1TPH9sA+Q
NcjQnQcK8aj1BHf+bd2hD/TumxgiM6Vm2gZ9xE/UFfY8MZfHj4AzzsHXiLvNo0to
ZUSewqH0GelNcBp+ZaKqo9wOdiJZDLuw00aOTLxQwR23yzhttA4oPIcL0nYKS5ag
vYe3DcJ4OBMr53pWR0d+2VdaxPC8BvAaEjWCaJfOL65/qZ/5bfZm9hHJpWSZWR5+
g9iCHpX+wR9elEh64T8DkKD4qIf30Z3ZDv0bEcOXZHLMvpiv+jsu5bkKrFSxcluX
P5t29GhHptna3rV7VBx8+cDWhOUGrX2hNg/yM+qAA+y54g2KE01EwsUHuP58jqIS
4jeUoZ7YfYt1jcWMbVMk868b8GBgDaOfqn7bcsumsbXvzjJEUSckMxUKY3TuiCLT
lOt+/sFd/dSlNpgXhZSrgq3wFIrUSLQAZIdF6W9FAZe2Wjk147ITWGr4UNuLqoy7
i7lGw+MiVt9OWPVgREp1tMy5bItK8bf4dYy2Ulb1dy/yi8OZJ/8eKuNchr7bQlUB
LSb0ME2LTYeRcfr8E7WsFWTXCwvlHzNnz2USI43ku9VG7vvprF+ytGcLw6dDqciW
vW0ZysY7PW1Y0jT9zehk9nJv0k9Bs+FGO3oOBI9GIQMVcJYLLHFYJ06QqtCnWOel
t4MamWS+7P5b4U2QdFeXLgmaApo3Bk6biDbgM7tHFnG2D9IX9+Ok+GvfmHRcIZmR
xiBa5ycV6Jv/VPucdHyJ7yRXd0caexxyroVC7LfoRZajUV8JA57MOCyL7x1+xMKT
dKLr6eAXRv5M5fUMQYXAL/Q6MS5PlUl/BRjvJbZCZs0k7omBulhr5sl8mBuGDGWc
iLNQOAjiX71ocDoiVkTB82yM97rCotTKOznlsKwz93at8hmc3BePUa+V0LgbQeAp
O3TxkmExxLnZi0G6v9eh40Q7vwg2MhSIWPZRhmAlIWKnb5OWCtRJhGIU4YS6HWLS
5gn9OVIexE69N0PFVYaJtCaXmBd9b2cO9PH/AYnlkDMfGATwymJNwEnovBTcJRG1
2vp0mc+6giwu1qZZK3YiS5MpARYbr/Drb+/Vwnk07H8zIhhhwp/Cvm733+teHIuK
P6YVNvgo8Dp/Q+zWBAQDeLhsr3iT7r7KSLeIYsw7OVGN+z7/v3nQWoheLoh3+Nbh
ymasUGaN/CBHJJVklK41ZafbPyP9499QwkvedTMmBFSn/y+kxs89If0SclmcQAt5
notW23yTLW6wmItwcqzZU1Q3rLmhRsJiu30r2j/JilirEpMub0wznMthwSgy/Md2
ZoNcs3t+rxGg/8hA2BjzN51xtX4f4D7K7kMzc2XXlXKwULBJvTBd2urqRlcvRxw5
oJUrA7hHOnK3ySTT8tPivXup/JFF6i7L489J9mG/VmMpKFSYpfz42ujSUzFzV9Ag
KYU8NNDBJtrq9ThoTmbwiXjQ63DGmvwngWSct+L2KRiSurtWG9dbefWYqj7iV+IT
ZpRedMzW3ID+qZQxJ0/2TnLdnhuk2mff1H7Gh0lTh5ayg/pkkBge/W4fpTS+fqy+
XZqmzYTFYbDy/xa1+jw8wYoBaX19Ri+VcMxGRX6Y+An+OWSVkCkuKtqgo+pWFsov
2tZHA924eknKSwWoHylUjzEiyP4LW/I4KpxvxIsuQre7aWT3A77Kceg8PJY7fJ/h
JyCZ7GeApEPihfMFlRhazfZDYmSwed6FudJmGQKnRWlbRod4tL5OwhnKGAC30OGl
DAD8jtWpckPCv5Bv1HgMBDof8jC55rgmyVHISOmHVEDjsCJVFd29anDy00v1ASzK
wAuX5NHzq2eYZMjhEJw1/Bq9j3WYIrHe0qoyWr6fZk6FB6B8NUZcH4rwT+JPCndG
yHeaZedy7+MDvfAd0q9p2HDre5DHq0P5L30xKNu2kbypK+vDjw4dL/6QocSsufmI
EsCZztV4g2J1QCV6P9rtVRoDGOYyHL8Oe0DgZHnN13qIoa/8wO0iFRWhHNGoO+p8
PftOqo6IbQE4jcFAN7kkQ2/OwGSixhaBGE/C60YRU8/4Dgl72Is3Z4UhKVA3OPy9
z8IbT5TuLytEO19qE/jUtyPliw8TJ3tvsCrgCWQd30SXMq0cjLnF7HHJZf8HWBUW
3gDr/f9zqZ6OBQEH4naRTICpAZsyayQOHQpiIsRsGzNvmTzz6PABltE/9flAHsHV
ggwWRcMLZdmY/mWmmT1+94c3hLdH/c2ztBxA173d93zT5a3Wsf59H03/pydPALB6
fSFHVwhR8L0nmvAU2q5Cy3b9oNZdLOjkWu+XnO1+end6V8ePgeICvCII9tM+qlmY
qgOxwQvaZW919ZX5MJ3b/SGDPO4DZU9IaO++35YoE1wCp/ZwzkJqu39a0ZxbR7gU
gIT6HvJKyJfFWW8gT41y8gN+OJCH2pFl7ow33TJaKNOxAMYrjcW10C1SShcwi8LT
PAKsKtRRCPGMF7/mQgyHV+LYzL90zefnK+TryXC9UQUBbqEsh4Ibz50ABbaOZCRN
mwdMWars/ZP8CqksF9NgokPbe9RIke4xq4T6qJV+FxGurHrCFYNJ0ss1JTwwHzcD
0QHHXlFk2MP4aKqWdgukmfxZhMEXwxgTCbx3D3ZX22E25AkfPCXhsi6i1Q97uq7+
u76i0Vjap+iFILApNKghjgMsYdCdUUl4J4HQ1dbHXal0AD5H2aRAa/XxyTkrN4bM
G//Cbxv7eS7NKNA+znGT7aX3BMGMLin7Qi8ecu0mKNfSKv9bGmGzIFBV2FrkHYXR
Il4SdnvXflTwHtsYGvuiMeqR3oFYvecVgy0lyarLFu+407DgsSaeTUkEHLHjGXU1
8kQKIIu8hOENd3o9kWKAgUjF9/U8FWzPC48kxRHdN7ETYt6vWwMYEOB8FwTNy5uw
dQa7Qx6RlCxEVhu5SxB8CkndETxbPUzE40X5YOzGgMZSzcdK1v4/gpxTB2yKAz0W
T9++8JVTlKK5UflpslXFQQRX7WOVCV+wD+c+YWzV82HuGx4t180xA6+SsteIg7Yu
XI51PKIYlQQJd8vgDE+gxXNx46XL2JWgbQDVH5LznmZgYHOLRUGirwZk2fdgKIN8
KCW5SLBxAL+3Ooy8dGuJ+P/cM1tavuRktW6AeKhT/QD16brLSCRa4gyZLfg2x+yL
XXFZE6+5LBjiZRIDy7x0XGH3mxLDN5Drf6cp+dOyaEoc4jATpOYzg2GJwtxkZIj+
0uWqYdVSxwlvDntniCgxNfBTO8SFYDDSYpIVcpexEhoDurjFoA3Wji7J+xnL9aDY
xlQ0jq300XPnKlbd/rKxAvatjON73KDma2nSTEv/T1+jlXGIs0OvfdDJX4m5Rs3R
j4/PM080Nj/3+qa75L9v+TbJ0L6vl7e7Zkp2ZAC2OirIkzj8WITDGiwHCjeG2XAb
OBSrSnwdw0lgVO6dtjwHf12anEgoOcuOUj7WsRhnqn5c5SBOiIYKEITeqUcH9DK+
FiAPcdBN8UV206dAPMYyKa32UxEb/ZFJSSrOF8jP7pp03v03FVtvaJh2ToXlLFt4
3K8OR9UCcnfgjKq1SETiqK/2d/sUoU6ssxtbxTqQ9kXXWk9tUo27oY1rG20+HbJk
L9pkg1nQ9jXYuoZ4oJWen3/1Pf0IorBGt0ftAkMbY7u6BSLsuCi3YP1gRZcqILzT
vClmbpZv26Zmi5oF+U+l1C4nWKksykAjc+WX7DnPdkYaxQd4EcLtXfNiBuBrcbdk
JSPsEwfJWf3l8nnwWulmdkcW0glpiEkTNC/gEq1+l7HWH1ymbOuSPbhnLC1M+xc/
qBMmG7SExOb6uwQZnGOFk6h8nTVxIsd2fgsiU0XbZtfiBNlljROyWIZgKZYZxlG2
Icig8vmWJYUwW+sdioNsvt/7ZO6zwiZz1sbVbZW5r1rDBpceHKs2dhbwi0VRSg9B
XogzNl2Epv8m31fvOFIFAonMQoQy3D9lS7o4HIa1+N42tyvyrAQaukd3kdqc+Vj8
YWBafXS6yCeh+U/cmBs9xsuhHwl9Te00wYWtL119DLcrPo4QX1W26fPUs/lNjrWY
1zYk0/vv2655oKdPW3XxGI2vM+QnDJudH7WuFpsiDydqfCdnO7z9kkNUubpAnhZI
8DvNlyjjm/kXIlapUge7CMYas3WvGH8H6B9DPP/PrDPt7RuPBde+6OoaNBV5jNXo
E8HUif9w0yOXiPt8GxdZwQX1Hd4aRJKV2YwKiQKgSUkykfcmQypsRg4N3VXlv708
mb62oKrwna8Vm54mTgIiToV3HSfjK3KAq5C5i57K9oUokZrhV2x43KXwbjXV/FWd
DmU/OKXZNucrz2WhmL7bzrm9/+kaBSEgMft03xo9NUPM3jf8nvup/3j5ZtWZQkwS
y+VHWmR2Ps/58Ll+6W+BN8RL95ZC0wyOZFE3pzs/MuOUFnbBY1LRHg8MXIW7qr8o
wKRBRjhVsSkiLQ3HGMEhl597we9PBYHTP3PZNQrC5YC8ChDo2I+FA9afSUh+pZCx
Uct9KNyRL3KibNM9ZBSzuknCSCoorC6z1a9kfL6nMxkL2bCbizaOpQMbUfUqbfIT
Wt/kqn61mjRxsCrbaVokACuMN4yqdtuQkOf0jjBUp2nbXu+VFdezWdm8tTuhjVe1
P5YLNuIGmi1kKSsl9mU9ETMmfargRAkg8VJL4xTjhGZ2cB1mPjDBNEmepg6vSHiG
KrRKgrKmdCr7na+xujQH1ABNU6w7V+H1PhbYw/vOkcMCoHqYeZ6g8SLQDBHE3jj2
jM+9R/rhGTZF4Znvt6no50B3v6ZjXJf/LNo7nJSxZpPJisW8YhLzQ4keCenGtxsn
HXyrDMeDrAZluiNMar68TGuTVzXio+DiXAENLgpV7eDwaWh+upUKN9MOviqNNASB
qmaBuo7vPaNTuabV8uJphdcXXvz/u01HD5Kez8sKlPpZarwuQFlV/5k5J0XxKfbY
5Tq7/NijvHAlwiVsWwPxLblLSQLhL0VF5bwT+3zOKwXEjeZ4gNHEOmzL+sh9pQCw
oOMzvsW0Whs4D6GVDx9TyvVwBRW5b7NBY3Yqjob6zwOZhjdPoyFi3NLREdhtnxnY
bkzCuBxWSPYpwHIosCnT5ilZ2NI7TQ5+xZJwHFo8UX+MH0GJQsgSsI0StJKB8Vgz
7PluHCgvHRrwksI6IRn0QpdDlo3ylMgVy7Rz4gACghS+R0sqMdldL24tYcZaOLRI
1tGj4Oz8xYEqJHY949YjiX6UMMYbPGSYiI5S0SPlftmraaXTlp0L8acmK9eyRDsz
+CPmOxVc+BRc7Ryv0yYrMguav2VfR16IJKIzOcnX+8p5UgChIkkthrQL4WI9W+uc
qLixBiQ33XCt2gcf6oHl78teYRV+/bL7qBCGjipHtT8ZUohStX76EIhsShXtvW/C
NONLX8xB91lp5yy8+R4ZAo7tdb7wXH+kLUkCT6px2Z1vSjWo488Y9hz3yBXmTv5N
OuPvvG4dxBdVtW+SFN8XSGnirUtU8VuMS3qzyXkOneNoU5CzxtAgZvW2ndh3EmKZ
IoGx8m3U2Jx/Px3DRfXPprPrQEIEOHn14WAd5v5CPQrJGJi4rhl9t/l0p+T8qHLp
aYOLIB6hEowAGgv5oOLc+wtmeAoOGl3pVPx9dh98U/uA819CEFPbggNJDPIjNUu0
AAeZI6vuqeZyIboOLzl5e8EbYsiQ+iNsl6LUUyxq2L6eOMtH51KxTm6lQINOhfnA
aWr1PeKjgtun7wZOCzEkKtiREN9m8pTKA9WStpUnL1kFN2ECvFsZv6u7HHf8y4BS
A+bF3FqnRIFUtQp9X5K8A0ay+kHtL0ABT5OfIYqLYZNZciX6NgusKCaPdsJR43My
wpRXbne5GWTDn/1r4YPQ7fV28ikTJ6a9waszAeqI3HN+IWWI2YjYtqg7Krf+lmqN
hOcp4KLSzwdNE3Q3GQ2ORk3iZRqHQyDc/0A4NG0cw9/4VrzXD99yhF88hZnY4VHF
SlqbLd2zQVJ79M2m126cDM4bbq2cRflywz/bv3j6UZsIopp3rAAgsqRLHqAG48lV
kBwQKLrns49yT9ND2/k7IJN3h27YnXCgTPUCpDTWizh/mFCBqZD+4qfN5/nILJwd
oKrNOM3/3neC8Yf3HwzaBcgfroVYx5b8jLgLkV4MkZzRcC7vslae9O6XydgFsds4
5nzOMYvAjBG/FX9cDOn8cZwjmjAKVukb2WXLP2qb7RhynYZcGGJie8BLAuLK0NHP
mHOmDwGwoorMxK3MPp5XRB8VfxKJWcliqb7D9NCdoIMd9IhQhMpi4vJobZtoXDZO
JPwzMrJB7HbO+NDXcFaAizbFAxdXyY7hh2jHFCorH5vJ4i+Ft2teZnHebOdXTxph
DSJFL7vWuqJRHEO36BrlaLYMTqcuB6pD7m9AEKSu/yhp1fSWMPI9BA/SrLmo2PYa
oDcWmIioo3JpbODJdVV1ye2QcKZfQLlUg1es7HsGbQrnFjgzkCMRe0K5E6OOf2aB
OuWms81YS2Swt2+f1dU4HnIKy1MM9FPl6LYLbnijQC3f/8mJPIlTE5gSJlRoEekQ
+GG6DATMTfIhnAkEI8GzK84xoJv5Yl5ODNOmlAx6QZ+lNCUwx+v9yivzXt1JugS8
rD+2lFuCyWqzA2NiOuGSrYfKaG+0SaDEY2OZ6ZstxXlYGZAwNX0m0C37TtS2D2sk
g0veqHx9muLdjLJkQ5Blu4bdhM/CpgWqm9wvkViqGIBFfzVYFRihEoTHLgCBrEgE
aZTaw1dVzsXv0yKPyt0vr6yMPwCDzwXyTmM9JxLTUCvTz9U16J0Q1Lb9w/VXlJmT
gWnZ5dsZ3o7H8FKIpRBO6Jngd37ut/5idxkaEwJocLyqWlrHsYJegiAXEHLAiEi4
dyoiNwuW2U9ggzH709wjPTack1B2VMNLY1/kyMJGUDSyVN3RB3l+llnT0ujnDEMU
XRHxYZEmFPCoobKGE54WL1mck2SNg6pLPWyS3qjRQagaCj58teMCw/Wm7AEFn8/2
hCkMX4tSdqpWpMRO4GAWA/Oc9nW8xCPGqJ5HcHVqQ4H4TLKhkxFpqw/t4ptvcqF5
7AnraotGrDso9IGaWoRXCPo6WZgcIiKGbbgLWPi8yB6TfPFn8zEwmxRju9EnLDAh
I7nSJQTjLc7uxHJuMUNprKsYHWD+tukiX9SgA0m3JdOotZBWOvs1HRghbcf40ys8
ao0oOjl2wJE/v1Cn+8r1gMNpPiYh5ZVFJG2153QIgLFszIFTsihRrgSIJ/EjYe+b
8d6sHMp2Ho6vB/0YCpIXhaHk6Kk0u+7DaMdjRp4vGUp2Npov/rilHLqRWRjXU91o
vbZvLNV5DknoBo48XS0InZI4qV4eNdoWqcvjRHE6efeYSz9cknyEy0Gyzpw27hA1
wjrb5R8kLUcilIFAZ0uTamUzutN+WEcsafxOCRy0NtMccK5P+4wAWhlCW6adVkak
GOoYHxy1qdjE0vIerg+/gopz81cwYNSI3ML05/k7O6E4Xqg7NJk/kbFG2DC1hK2m
hMTZWWrE7/4IQQgd6VEzy6o+xxjSstX0lpv0BUZ8jogqB6B8z7+YHXN7LWHGZQgl
kks6y5WI/I4hZIPQHw16u9leXoQB1iwn+EA2hjQU0PiWRsmJ3L8C3t4OQ7y+EZKS
zyEQ5gsOs2TBDe5hQHNrSiiianRX8KUadAAHq2Bf1Xnpb1r5F58f3XoIjCQjf8uv
+dljy2HZEZhoKfpM6WZ7J7KsIPEJddUoKRBO8qAR2lJAZVh/D0qWAM9Mjqcubelq
ViXdKSUXXCWwApjkoRYKWGeU6Iq7IqFwDhoDDjd6CWBWdn6odUzSWKV1Y1MfEc3k
je9llvdw9AJsTP4Zt1B4h1wUzE2gfwqT0XC1eI9R8i+7l1wGmpKRDVlUS9UiivZj
TPxiy3nXhFB7dT7KZlok3zdNhp64dwpM0BdbytEoYm5Krp6J6nYMAL5XwuBudpN6
gR55Zi1H8pKsvTNpOA9jADeFF6dX9GIM1NG8NBiJEWlzbTDzUltv3LosYIGhm+p2
2HyUMYHKIYMEA1LElbns2Fiu0movx9c3e3MiWxn1NdoOKCYqKOmgsHORbFoLGyGa
wya2CxYP6iS71uF0maoOJtW8sXzxO2BRMcNZAzZC1KCU3Ts+woZ5lwLPvjgpcnFg
SCLvTcx8CN9XmQpvIfmKWN/gBlaHpopxQ1UoOSOBaw1s/uYiF1d+dolePCWdchA4
FjofFMEjI9mOrbGIE+BZ7XQvwnlEixuDu1AW9F48G8uS4cOTZTlhYSg3hssklT+J
KmCc1i8zZR1u9PZ5kEq0RTJLkEbgNEiwQ7v0zpPZjvOSx6CckaTI7s6QaY33Rg5f
opaLkZfbPAWiyP9JxM9OWuKoJLs7PTzPO1/0pjRyV0xPVH2oJ6p01A+mWUIMd76S
8I5bannytFJjTlOQn2VOe0PLvRzvW0yp3JbwJharHAdhnb3xuLbotNIhKulwBuQ3
eqOZyvxCxTisMOBQA2nBoNgo4GBc9xHYNyGg8RhH7QkMuSDbG2TWLoJa6pt+rhfT
4asvGnlaFbxySjVnUWYgYkuSGKNTFAsSGZashwRtYnY84oHKHtIm4l00u6nSiHKB
cPJJpfSF8F4LZ5qFheud8iy/f7WBVMc+PNypx3azAYcPvAtwSLrtkOzYHjzU1A6O
4r/CfCAzgEJrprPIJzAE3O4VuKWCLe8MXatC6pOnwCGVpTYMPibP9aAE3vdjnOiV
51+7EOOwiXuJfW7b3AowMnoUOlG3x//OAoBnNi6hXlCE+9zWpcS3C1Sc8lxu9Qx+
qDPqquSPnYoNCbLVNA5uaVCpjo8GWHoNnkpml7lMX9expSk0xefouhRA+lbNTUk5
ewMciuLVV+mRW2pra52dgFsiGtN5eqld/VtL90zI9/FfCvQ4+CV5kFpb3rlY2crs
Qg4vM4fZ9lNIrUe2OGH06l7wPZrQMWK2zf74MI7NDBPoG5ASktzPgyXSJfWhQEoC
fQL3zfVFJso72AWFKssa9FnY+ZyhmsISnssANOd3cAkugd3fJRo0jbs1TIrmq2ze
D/Sns85QHuiWDNufVq6v1lqvVYwh2+Ih30gUXpsIoXTPqfX5q0urmHcQNVGi4Bwx
Jh1M6h3nDdYi2SBcvQK39JsEBnkwWlk7Rc8CVc6Ic7tS9qLnteoMo5ygZi6k9QkS
vsvAEdFRRgEn9fItGsMmwLpdM9sTsjqj/P4CQTzoYdf1nA6VKN3RCaHwKKh7euuR
rGnJuEKvufGBFU23PyZAXOyumzzBGgn/1sFlr0zMUkCN8BwHtvcdOY5FmGVwQc6V
JPaS2f1idbfZPZrElldl2RB4vaRzODn6GPFP/GD1ewy5er2zndOSZqWbirCHVSD2
sgM4Dvc/P+xCrwP7j452fLpkjvPEH20tS2wTixB+syHVShhuGX+VLbCpd0P5I0An
dnhPjYM3nZ3BOnZj2unJGYBADA3x0mJEBvW/kDchgW5xsFlefS21EIo/eRBbo+TB
LAa/VQDZl9HyK+S+JZzejTzT0WtS1m8spAlKHJqSYI5gNrvT0NnT0Nt0R11gNF79
2Kq/T2owye4Mn1nN6i4SIKi4Zazvbq107kY7hCJlCcGg2ToYSHesN6DwEXXNJUlr
m8+6JYq8UYik3VQzWtIzztid0hrASoGskX2Cr8YwOgCd5Gf2RlB4qW9VkRu3l/wz
+emX4qvpOxTLJuyGUirDstfR6PEslF44DOOVt3TCl2/reWUTqZOaO+HY26C0RjAC
SjBG39A0nVb5DUEUJIl8ptu76gG3TKJklo1dQCcOUwScb0oV7qTYtReAv2wT1Rye
BqAtxTB3/Uv9uX06Tnf34I5IuRaLOo/UCn8a3gEv+pTx+9SS26taKfmhgPpEfrCo
E6jM8mnB8cbKD3ezTe736jPdNw/f9FW574WXZe4UAV/TEqOmQEkAwR9/aCglZL39
SoutGtYGg2M4XzmEcx3SiRN9m8MdcDnipyfE+5noy1si9LyTJq4/wiUmEPjiWANe
6ncDC6ENfFyL9+lpAe4BRzxcYGVJ7lJdL1Va4FqYEpN9xWK0e9anQUhTBKR7n29W
WDpe1W3y7KCeG7483mT1dNxNFZdwJ1gHPgsxMrXr+3sgs4EaI3/Qc6vMeCxndfHn
ALWYM24vRJBJuBDMpcRPUiYBpfxGZ3B5iUXnVTBU20Gyq0GTjpvtA7hX0dIcQcr7
qAyzycaFrTjpv9YgH+oLpRfNEHSAdkIEU9vfXNF85I3EzSlHJ1Iq6gBU5lpNenMB
RR3BpsJfG6wUpeBZApv1I7TiBoBH7hfjoeejjSd8kdSVDuiU7HRKDzTvzFDEvWKI
RQQl9IQmv5ZvzPoPyhfuWLgrpj/P+TumUH4wDMdqdm8hfYMkmGrhiA8d31ePY8UI
1+XWIekrErtEh+wsnDwUloyDxcJAFP+Lt5JqrTmxk9V6fMNwx8/1OksKtSGqscpZ
zl3wwYyxACPQHv6J+5rUWh27uJk0nYBtYfOPis+D17IzuoPPpMmNZ2Eq4dTuah7z
ofxSsc9uRP5HFm7IU7LqArm2AkRh/3SrRPONEmPEv53ZuP70kl69sCrkppZBVBYR
xx6OBK4faAuJiYeiCenm8HFzO6fjJ+Psgpn/jqsxFDZi+lNGVym6mD3hxTs8+oar
32bmxLlJuIo5x80IUdxugKq4LFY7lU4HLVAA9ITMkUGKXN1bwKDro6nC/IS6V3qB
Po8HMLnOlCGwMhC1VWQhYvXjQ+iGV64ZaUEWFLYggkjht9STCzLR/9RG4jZ/37P6
mD5xLu6LbqJzta9Sig/CvbOOXPxJdsPLCoHfVCDR+BWVZ9XN/Ayrsxck2nWbEGTT
uiSaenfOMgHRtR2vmH3LvyffB8tCPRBTL5UATbHQSZFMROHSK8kQm6pjdOF9Ycf9
GqOM8M3G+1oelglvg6yN2Q5kF+kJUMNJVvHvp6PnHTSBAVct8+uuMaZVEQ5GFeqb
ishfBwCA1MfJojDnU4kNT0HG6ary15D3ldSz0+zHI6VV2rtC6dTjR5LtDyy76uWj
RsNQY7z7xtuZ8rg8Uer/mEhbH9bD3wIf+G6QirnCovoC4rkuMl629yoxfkTahPZM
j1lZkGH+R0/LGAcG/fzHFHYnmqGOudwmxJI966DyljKTlpZtAV2KuTZpnSENLRKY
z13oPmTkOmCbIjG3S9uuRdFgyXn6TfOAs4v5OUiwJydpqwyHCoBkai+dUwwJ3aTJ
aQ7BmYnPpcbnA8SKKhhoAIk0PX8JjDILxgDUvnmBFxWb1KdSbUOZBZELXwd0Ir3C
AO7XT9OzOii02d2oH9msZ/NWnp0SqijwG5wRztCMwBURpEIv/gyLBvUB6QYzRsKx
wIwB8VZKgNgQzYkvVPzJzTSMSodTgkKE4LHiAScKPxXnjBbyd2ZfSUUeFTtKpEOL
DkHOaPaFvo1CUQHdjI+1fMGs3ulIrps2TOqudfClPepMNnvI/bNUMNXNmWYJBoSr
BtC9h28dbt0YPNhOLBjTH1l0JDl2DYIfFvgNrbInivwkjOtIZ9SLbZm3nI40NCtP
xLckQbG0mD7LrxmWdguoCscxSSYoofDflUVqYtf3fhuwYtJZrPrUYOZWS4VVSaLr
BN1ueWzxtPzDkRBaihprNOb6VWrBSNfH5CV8OFvXONeodbT2dN1fG8vafSbXVUG/
YgleLpW5FQnncJaPGIbBIreqtVX6avEBJYdsF6ocuore0s4VKkno1riBEHXj/Vfr
9rQCZHIFC4DZpt9s1KcRymMM0jRHiJ2/wT8tJpR8vUU57ATgV0XTPZrQbTzcRzVn
DzkEbpoKVI+5SWaMoHiN37QuuopWSjAGIkM0ySgXXKLmvPo6EfGctnG4VbDcnLea
BNr2tQ8U5YrosTGzBo8TR61KPXvTzBy6oaPUj5CgJ64NUqiV3MfH8ZO2GUDXrpD/
z8lFpqL1G+D0yzgh4K5hYxO5//pIT1Ot5tA+0Uqa5/WsXAxMvc5zlRwaIqdegjOO
q1oFrcCqu2yb0DlDZZ++LY7D9VxXcyzK2BFEjwd82g2CPcwLcmZA2G/NwkgRxqP0
aAfM87gcyetd1aaA4rJeyTpGBr8ETG+Vb6DPoN6uIIptQdZClcTh5IWCcA1iADk0
d5G0FsyT6coJwSCHurjExQ9Peo9OnVe60tMURoNM54l+RFD7R7VR4hZ3OfBgGK4e
grhxVHtsC8Jp6Krc/YCKi5kKSlmzpyhhQ92RO9Oi7epptDruWpbk69aMmgSa2Ekc
BjQOcCNXS+I9dQN0OObXJzY6QzmFqH7hLjFPiELAZlfQQoBVPu6RR9pqCKphEo39
RbvgmzQx1PcS3obAN2Gs7DclpiL30m3zs5sCWGqrOCBdFQ0dBzR7YFSrQU6sendo
oudJyoLgQ8ykYrXoFp2LNm3krs9VpN3i7Pg0Tv7Pt+wKtkbVZZn+asGrmaOlwrJE
uQxfzuDUiERjvJ8JaWGTAsHJKf2Bh/4FuDxyGh+DDPHouGtY/7b6Lhj1dh0qBpiD
EVLb3OZOJxneshIn4hQ8uD+L/kUshKIlvRppcmweXWQy4JaT1l9yiUfDkhNOdXxr
VyiMDdCdmiHB9ZEgmjpRKh3rNSm72ti8G3sasAPGwHh+CHu2lxiZ0552sbfdOK9V
tAUS/JAq9IYrH+T12RzoVIXPn0FouGKpgT/YeeJQdfQW0SyFPA+u3kFCKi4CCDYo
omlwpEDlJNw+IbiuEHX5r5X70TvxbJ0LrrFYJN1dtGnTzPlN3816yUkhrWXJ2Rcx
DLJzkV8wa5uv06w7fxtQ1rp3rNFwgmVH9W7/K8vLAqV6/XnvEwp9RliO2LkvEeEj
J+eA3XufKq2nKjfJxCk6qPXGqWmBBO8yiuewm3DgL+u94NdNgwh9qunI8B1NVw3a
q9GGQTLCe0ivjSzckUSZYcCuqG7JMqQSBehG2MBv3ov+0RoM0Ngztctt4qOkx3tb
byh0bxZOnCq+nt6MADlALieO8z1B1aBVppXf7M26hmarfnSl4qsdl7wiDi4Hs361
ik6vYx5Tjy/YsQNw9Me4SlSKKM0CseR97n1EOeolapo5C2lDNBjPRZMJJp6cmLcg
nH31Y8tsYgO8y2kTkmUzerEKlz6r0pAdyOvA+afpTKA1JDz3/pdlI60o+D0puKhp
zE5dtLoHjvoCAoRSn+JrWv4VwjRV1DmO/cEXYKrwlGFVAOL3GELatzu7jDa0wvTv
0nnAh6+deW1VXmXXrSDIWR5H8mQjBdqkcgkx6IjuHkO94oK6FbeCkE7HrnDQL53K
7vBRg7wAqcz6QV2EndlnmpbtAxOQp3LHi1iHJ68G7XNk1piu6k/mSL9ojANbSgWg
vyjwj0NLLYtMQW2duyRV/zdCT8OtT4gjvgQ4eemM3WloT0qxTNN7Jf00bbqyZz1e
YNDrGyNMC5api7tc3Mm25w8q7pC3AfFZwoxpv4oNZFDaDOyfj+cudjQzHi1HsByJ
fCs7y5cEUFsvqbTxz1IPYVF5DefiSqDNZQfLuJU98xS2aJ7c0ncyV8BVgfM6wQ0X
dmtrYMRgI3gMaB/m+f+6kBMoYbW1B7sfJnZU+wus7e9k8mx3zNrdLNJqA3VvJYjP
xv7JRiLQ9SKfvjw3dzvINZLx068Bg9F7hi4MCEpMFnjDiwKVgMswNh2ECPJMzXEO
pJOqIuNKtSunEW901O7r6Hf36v0FCO8+d6xUhnSKwKDTE1RU0YW/saQ4rcJGa6o/
gcgQCaxdjMjv0XnuCDkcOrw+Fy2xOEDGTSm3PxcVyy2N7age9Rim35VOra3ONb/t
eBVw810a0uJyJ9sfod/FNXQw05TR04NTpIcK/DE4poRBBP1/tqrEoOp51tSVCzFe
QHs9p/KTi/sldwhui7ZX7L9Rl38G1AMEpx27XBx2O/djR4LvjAmEvkc9CsMfnPNr
VwODaewBXjAv1z2uiZ8rk6/BeUdZxq24owqjMV4Tf8wUWb3UrHA0xwpk3w9FhZA6
v19FdwZtwXuxTcxSnr43V2Iqjc7yejaeVq5Sk9o9JebJ4YIF+6MPVvMlqTPt039B
VhDMpCqxvkH2T4F/QxErkebyKUSuxLpg75LIiKBPPw3UL7lb0dRiZ0rrOE3UYIfO
68hs93+z44RMqzgovYY4GUMOU4R9SQ8zEd1jSD0TUsGX06wtddbhivAIZwRDjg+Z
RKoKYH71pz0QY6pI8vQJCJWVk58JfpFFrHMyDor5GuM3uJU6+360rA0MJE72rqAu
uAkJSNdMXNegodUegqaO2nYSD7pw0eblnNBP4oQTlAn31zj26LBf/6YP0LHvVmv3
o7MlZQvN34CaDefF7s2nGFFV4JmEEKlAVMJ0fTiLY16fsZPf1x0OrA5agSF73shD
rh8iEcpPTIEKNeiearthrJDMdpqcymE63JWIxukb42SC2Vz7Mqy7266xcs8wxdkq
+AlQxh4rq594LnfdfRh0YFfihhlZA+TnBOaDAoZwFuE/mf9iHMRnf/wRTROAvvCH
U19AhgIAVbuC4DTf3QF44w3X6vLAJH3lpM+AbgKELJbcjWabkyVGcyxbVb46uOem
4rUmNWpGf5FyoQGgWdaE7CLADVsVt6aPfphvQSvICRIWKIn5YRDXPIcAnQaduNgb
w9GNYgM5yGr2MjtGHhr9azyF32O2JT0CRnNoflCoI5Pv5LJydnvkQXxL3j6wOFFK
k/f+CEVuALGbvwC0C58+jbwMEw803q8LDQFNZdoU/Ly4nZi6goPdZX8xDFumiRG+
FX853R1UVweXmFL7zJLhcXd7QAtwbiE5xhbMdsKwewMryyPbcPJplMRnGOr3ete9
l5F/sW+GbkVi4cODqGYfhL4PrD52fKGBc7dTJS30XhJPEAKLVRPi8zn/aODnerBh
g3GCJb/DsFBRWHP5NYybaf9fFukg6Yra7M5B6zgw+uUgWQElb+EWd9IopCBL3nnw
O9QyQII/DqT+sT1rxSnHhATAZL9Md3hAByxFmJKH895fC4Uwv6n8NBoED8aSr81F
RfxHuoHnoDtYKmZk7tzoL42wIB7dsQf/IVXETTp7nBXCtRZ4zktLAYPKGcAgPXRk
MLKbTeO2un1b1yK8DZ2RfwPgpcrBpdt6tO8mBcj9Wwp0Wj+CIM7R1MjL4HkFbsO9
CMsQqUeyJsZ8F/8ccmjo9FE9UhCUa/lwOJ0fWBmuaEjYZuDqGjCCXbZnZMV0QCuE
GhPsw9piyrHOoTJDET+l3L0z8HK8anFxwoEzqE58imCwKj5K/ELcEUSzDs9k/otb
uAJe06hYO2JnLc7UkdBbY6Fik06twOnASCSrIvAO5bvowBr0qNAcchik4zWgps/S
pQzRqHYogk/PtlAysfY9eExLBpeWJa4QqQOvrr0OeWqt2a7egXs2CTZ6xh9jPmHC
a+v5C/hd8gwB+mKctNX7wI8EgjZfY33q/Fc5W27AUr6t+DY9e6WNW8T0KnBZCNuX
+CTri0G4NMhSZHAp71RAUKwp67yLpageexXzfUiQOV5ncHYzTk9TojQGwftgxbbx
ObELWMA6s8FVoNyIqEuwvC31EWiNNt0MlxqYXn2yhu2Z6HYzic06SD6MIu/lhgAy
zQ1OVNpOq+MT/+jkXjSRnrmV8PM3YInmTVYKPdN77nIV+fBQteVc6v68vhwwjbNV
Yn6RtSiMnV433QAWWL+QuCONBTAtabYgcq4eXr7CYp050PVGxYtgmk5SNboiJuz5
Dpbr6jkOdWpagJpeIgkRgQAKK1KqUrt7zBgJk1qFyRJMZARnYWNtu7R4w6F5TR2d
bi7DU6TdhUgDYNJcuLR5nYm3ZKbnJah6x4CtkT5jIyxFzuL6m9LF9/h0Dy0HZCBL
c3zQMcQCae4wa1t59/okVx82Se+vaCUVHMy/UpSfgQlLG9VhSQMIkIRauozgVAgG
6RKmwbI4QQOc9ZimnQDYREijZfn/Ywr5Itg2pNrV2YuUI9etTVtQEx8T5jtYdnNI
SZXkuuLF9U+kPGXpdl+stR3holLCa9vAkAR1/DxPwI80ltZpmNjXDZPN1LH/3uQp
bhia/xaEVCc4rwqhdIfPWN/Sd5GXByOEfKAvPeB3xGCrgP1ZLT4eK/BKoV/YKg2C
7EpaOZEn/64PnTJfv7ahJxlCBfO37LnTkXHzhSNZSZbiVISr0r49/v0E23YQokMm
odEjSFt34B2+8dQetBqLZg8zc2HVQznK2r3kqgqVRGi9NdGvfVyr4wfK2CMVlpOQ
IQjvK3N5eB5c8Ly+5qaeRAP/8xYjfXz7RMpSaKbExeG3dddDhRf5jqVB3RuueKYL
GRr0OPRvSsZSNNcjcbw8RUhizmX2SXjeFq+9W5Gr8Ffj6+tc3lA0I8n1cVfNzff1
lXrvFM3GfRlFtlYobaSUHvdxt7hynzZhNsdvkeEVCAuUXV3fB/WxEn4HHWQmlnAf
qn0iD6AdCj0nftC8sQ8gn8RivdDh4NeNKKsjeZBSVNijLB0bPVAXkj0k00oeJ4HV
yX4xHSgf2/dW9AwWdrbp0iNwvK126Uymo/i0y4rQ80bEPiaU1t/yRhEd+iHoIYC3
RNh4+QtqhCLxRdXBoOkV+1SL/2amSNX/Qx6ysJWqMB9Dm+qjyixdw8V6NkEFa1gv
SqUquaz4zMzvz1nUbMIW/q7MeZ/1fDsif4SGM0JwnmorF5mhW0c1t0awhZiJoVMN
j9+mqOoqw5+VpJpqDqcQjvMIcjzPgWTXFGr8lPFq1LJO8N45rHMyaT7oDFg5bBO3
4n3rab3oFwp1jwvPdqWOO+UeLfn2tiEsAhiywoXDpiJMM++1/5Ml9w0AuSgxBib/
6cuje+PLAVMtfxBpY6+4+dK2Ia21TBMFd9upU1Jm3CU0xPjS6ugVrkwu+rH1MFZy
fe5Xr2V+rT1INzkB5TfCEiV18p6gJldQLt0QszlJYmyKCeU/72YQw8NeGFNWa7ZH
8eTqs4j3cz3kCRkH8wbZnOJl4jIvbrQyomqADT1Kry0K+JG8y0oYGXhgYhsPingg
ePzUJRH0WIcq8vEbOy250dWd2sKB1LZISV2fOBYPoWKdteFn5wUFcBSwmaRSh5fC
JRsBruuVwDrF5spWx0VPcXBZ4M/BE/H4FP5i0Bnbh+PmmeDhaac8MTqz34zBzQcZ
Zi1smmlN2twtFIcubH7GR7w3uEdl1RfUtS+JmB/+2JI3Bd5osG/Zm6MRTtJa4Bj1
Tvu/tJRFIAGUAcMNxO7Y7wALzsts/JYDGaYT++UB7Csl7oD8085kFddU47J8C8EA
+B5m3sRoO9mP4boAwZj30vvYa26YZgfBS7ElvoDOsVKFkFVfe+MtPXk1OY2AFjzi
ZBtdB4pqQPsz/YleE0l0Weik4LGVwRwn/E4ysoj3ATzD3so40aLAht6WJfEk5TU4
xklgsrdk3AuO+E7eH1Ps9l6vsfFKI6UOaflQUdU0xG31uptbMG61ShBWruDO9Z5i
aOrcC2jlGe2Zq80c9EUzaUrXefeBkgw+bw3yJ2f6IaLi7AwxMO4t8Uv+IFbDEhFw
8nzysfFDHtH3L6PZy/rPhOKZciEW+sFl85coYVOxfdL/o93JYiRfy8KScKxzghZ6
tkfNfDkohpeuByDqoSb9jE63+q9UhVNuF8iuD5TN2OjaKyaI9MborvK8kb8i1e6D
1VfBMcTbyRBnjULelzkbaYiXKfEWFbpk/ycMDRzheF2lXzIBYjSJFYRRnt0PiYJp
85/IWFt2sV2u4kl8ct1j4Qrc1X4rkAGob7L8qa9FeE8Y+WeMXISSt4wZ40p1gtwR
HHUDdpirwUHiFFRyj0BoF/ZSuloYFqGTLo0vkPxH/9a4qo/dsjdGICNFX76G1uIk
6B5SHpYiO8VISbMeeNTibKeVhcVtX04XPuapv1UeQ1m3YZuUGWZ2n8IxaFzvQODr
PFAVRt6ay3sIxvdpn4bRn1m6nMSOYLupD0sL/eaMt1AbmkfeFwTvPZKbJopSqRlY
018sqViqkmi/BT4wX359OYtDntZDt8vNpjZgLvtQi8OJKfQGKkldZNa8H5FrkLmj
ohBHQ2u+VhBJSGlVJcPmntSN38/MWIzYiWfb3ubrhWUWdk7/72ZPX2XZ1WbWeBc2
GQq8ohZAddttbCJaSknrkxxGJytQeXA7LOKjlMZRH2rkmvVA482XdOToCr06d+0e
ccFJvZzEquc98baJAjsT0fL5A0ppPkdRNwHJfzZSoHmgKDbu2K3DfiUKOpejxj/y
g2kzbYaQDZgHvae2qLqSmGcP3DQZEai+4IKlvHjR9Xc9xXymMP74SaxorjyqRbx4
sQ39rjwUpqAH47rjb68VfqnRuq1pm90v/87WU9lrcWlZwDML1X42ibgLArRH6eZ5
3SJkjFsfFyCYHJiw2tpO669F1fh5G5T3cea4GGnrS1R31mKFKV6dCoOvWVZdoH5o
sC1src1mfeCn/7HvMZREVN6lplUnVjg7T6sjcvACcIsXfFbHMZpvg+gd/JC+xIvU
VP5xqmI9AeLJUk4lAGy5w+MAwC+yxy2ryOjuaPpPHmIhNd8kpemljVy5XmGe2M3s
dgEdeBiiiwIkBsnky2dejc3jEONJZ2DVUN47oms8SHXuoGhiTm/l0xVTP9RCDafv
L2eMO7UY1sdw9UNG0hxKp0ibwUmjPvxtYMsijc1azc9qR3cVYjU1ArXq2hXrYl4d
kbACgqj7Vw+i6j04Mx6v5svGOb2eNQnHsqSMoG8L3ksqOppdN3Fj4KZFalDg2h7q
D5nxVr7aUuemzjO9tXhonzJERYr/9e6HSFBbhsynWAWy8IEs7e2/uXPlC6lybL7u
ykw6shqaE1yKyHcGPrvpP5PIS0K+nXaseeAoFSLHxhzx2Ht56o9Yc0wl1CvBoSp7
//uHdZA7bmgnpIK3yjXL9Hc1m2x5kjOuuX0LII/9IaZC3wm6ToxPQLT86SFp2bWA
eETdumG8XMDmeTGpHLIoKMgMLO8DeM6Yy0eg53CuP8SyX8jSYhZguMHrT5a7yEDB
YVtV98iV2e9mWv+ZADb7SQxTcq8xMeSUNo1P4M62qtpE8XTk/k3cSDxXp6GehfFU
oVRpdeNQ91KERRSTEePFp4xfi8zu3hSrz6uU0QZlP7STTs35mjemSO22DYJYtD4z
5L7uY4uXPorQmO1eWxhav7P6hv/Zg4nQ2VshLQivoz2RPucomUP3mdPv9Nh6wWCY
n5DMT/WFqFRUFFIvwETQ1px/Mn5bGohzWu+x5t5Txt7iiIadbKWNxBeQ9xHGxDyU
VkjPxYQx4VMe+bMur8v2F66HVUd8nwfe5y3+kps2IPBJoNYGdhBnoqqnEO3H0+qV
qT/BKkwEher80d+Bx9HJavt4tZxpmBup8yD/33LPv+ehZejD6o4EzmEMjx49rYU/
3jT4evMOkbQCWLCTP2J7YPDHLLKOQJme7qfJQ7i1kjiE2DHT67sTiF0TMvwSrYcP
Dsw8DxISYhvr2R2wua9HMU7QlfhULVZUDUYCGn+4gaaodSw6kiquBMCFjOe88cGQ
dHPUGN9sZmJJfccWBpWj2MEDjp1uf4XxrQHOGsuMSxcNVXvXvRRW0v/q9IJUTtjj
JT16LT7CorYHuKr9nFQTv3JnUJRKn4VmeJszcGkJbiUY6Dr7wf8JawfrYtexRcur
GAfnOync1xy9q85yb7h6RwoLHorgkMZQGzCHRBc9C9ZlbUWKPbQuBgIIHx1nYegW
bwvkeySeHWeTm3D0/JGCC2x49u/5zoh+m30DFLXS0oh40X01TM/OC8xBIgSSvx4e
B+SzLDZX5MlzPQFF9zivPcBZpz4wQ/ti0/YqpshHFooHAWrWdFBhlSWFjcLW87LK
bEHTSfEeWeb8gZN8fwZX2XffNS+kDH1SOT5UtFNjRQZWufoOFRzfs9gRUDILglHm
bWDzrCZJoHN7UA5wEjJd70FDzLY7NsK1Es3KNFqJXDO8s0xp9xzMZAcbI91rkkUV
JuH2K1HuKuEpp7PxlUPzc8iAFTZRov5ffCkIAlZKRPIIpQgfpuSg+R+tDdGDh5Eq
PAPHXq5F30xwRIB+fBT3VsnK3lj1x7a22rZJnSpx7mydFgGoVxBl1Y+AeUeX0FCO
XJcwNG2+GfvwMVY+vv2P/P8Alp1P5sgKsyiWyyXfUcCKueKzG2LqKaVdgaKD4xyF
a7ZXz8yIbHFBWMl3ppZmx+a934XQ8NroZO1dh+PpfZWHFLtQvzOotfcS8uDbuKzQ
jZQejuItVlGtC7lix4RlQu3R/1YvTaG7I0IWa3PHMibDgSWtg28mEj4XrbkwQ6MM
DvjfgZRBPCf8fwUY95onESxJDJrGf18SD6N6RIg878lqQH6wbaXjUlVfoPWt8d0w
uhdxGzr/eq+fAe5cbEWO767w739+o4jnkahfM7gAQn/uVSlYJw4hdDX9aZgMEDAI
gHmrwZ8V/Y4z2m62loNE/GP98KEiih1+wLRLADQMDoL86psIK7kacVzqhSMptBHs
Gvzl+78vDO6CGgjJeM5fmFyNENGBhHG6GRdBWoBZYnTVppK+QUMP1ASpYm9dXlmq
LWidzFsv7PNC2X//q1c9xlxGi1/IWPubs+K81J3XIRONdAQ3SVjwRFKyQQGibmpc
rcXQQOvnVKmfUXGhSIBQTJSLD4HB3KbW/1bINBEEXL9JZQx0AYtEg4KoTFSxmeym
m4i3u7eYZQDT0I1hHGmSWOWgASB5ctmBJj6mWA4hO6ryu82xP3VoiXXP2DxDhoRx
kzh2jKGU0bLQykunqMVPPXf2x3OEqzfgkDjSLfODHhz/W/6HskGnD0RZIwpNGqe7
2I8GShcam9CpI46xI0xabjCoaNvVNe7DNXf2F130Wtghak3BMw5nZQE8hAePYxZA
nNcLqwmejS1ebdV8NTvvTfCECCR0fkPMNhjm9etBzUfElrfP37DB69LZDPrY1xGT
WTfSi+huSCvOHRRw99HtCAAguyKFTlFTqu2tCpdpnJM4bwAIfr8x+tsvY2OtZHbL
lxrB0OTecjhN9LLxrq7bes5ha6TU9FAo/chryWOdtO7Lb49hqSc3zHoq7JRmAt+Q
0OEO9x0UmVmqZ+snjN8yyZIgJ/x01vGJgts1hssg6O9AFfGZaxYmb0pMVPK+8TLx
dJfmSvZ2M9gLD92Fzma7JIoomdTJTl+HMGzUtAruC+eSL8NsoPo/3a5hozVK7Wby
mU6ni96QUlsbMGWrPg9pm/9xHnkhb12N/EIZhyqwRfScaDcBsdOqBdNaH/n+30M+
pnZi5PV+dagLvCriNzM1gSSONj6oCF4KgkHesFNd/RAgW/WiAmVrWkOXGeh++oNU
c/1AwVlkw32WODjXSiJ9LMTnivvyTrL2gMdYKpC09BoFh2XQZdcouNNQLMptz6bQ
sZoSudgO6KT1KNIzgtymhH8GthaAuK6PDVglsuHDYjm08aoNyItQdQttUZQXpIPt
mpCHb40PJxMf4R6FNHwUMFN5b7K4nsjpvuQEA6/Mbqf9z5jOqiqVg1ZSN5GzXlOC
nNFITUgsLB5unNvIRxyaP/U11mXliYRwEnoV/u9vcjUkdxdsGplHBXBY5MLtam9B
BhHmQxBPXgedwOcfXUaCF8Lz9olZzaJLK7vPeYx00i+WjI/Mnrrpb/nq5omkIOjU
dDC66GAiHvKfFpvrAr6Qptpia2kTp5hfovduUROieI29RejMTjs4ugZXjLDh5WTo
/aAUVQHnebkwbQNmsJVgwdQiiwLEWsULaPkA/ru6hw2n2pqm2urIyfEGib0Tc5lc
K2b3zOQvdgl/NG4zPLdaZlaZRtkYf3McI537KK4zy22ZamN4/akcg2+5JifAhvSL
TY0lfHrhrXH2LOjD7OYGl/i3HY1tI3CK+Ytj40mBPcbQuj6Kokw5SarH2Kg60zoD
loEUosPl1QxkBKLXcp6UBbcbyL59R9LcEdjW6Ub2jbv/8yxL9N7ZhBTF2VB9NXzN
7bjcEfCA1OS0tKn0vppnP+RzxWyA++vb2ym018rDjOHaRGvKsPvambIp+oT9V0ag
nFNJ8vj7/dzzvv+u4MGZnklVaP896SJghjtGypiY6oVjlaFWX/vpFGkZ7FOyVaDf
xY4gOnq+p0uQ6K5EpKwQtgZcNKbF5PV4IAW80+rxZCHKph0loiQonKlWDD0gQXtl
DoEGWs/YrOtkCqHHBVZJdMGJjMIhor8cbHhTxLcqI25g1wwr+Fy3aFF333sGiHQ8
H4hnPyabfzJCm+NIblRdwSQb53PXvlbBdQZX6W0zoreadztFUR9uUESpR21qW6Pg
K2mzgn1REwt5yy6sxn+ecp6rKY5XjSPWvzOrXABI07hGFNWePHQCqgN1ViEtAJt7
Vx8Y5uzH4zhriivN5dBAvzE8MukbVALZ94S6fAYXN0tDRV1x2HWzZW1InKYYWhWc
DblgVMTSYYTcPCKBy9HblvpVgMNYKVlhCtDe6Y6URvhnFQXqr+xnlYj8O0AIyqZA
3mEFAtROLHr8QoO0bUsB0l1RMk++2Pso2VZfT417aPR5s1IgoRLo7yI9P1jbTDSx
92cd/+uzMqx1JbMqzgK4v+crk+jJLq2tf++mHKoftOpO4rJTwFZ4WPSdljE+R7NS
oJxZQSl3Um9QyFNf9vLHF5651zU2d7ow3Ukyd27wbuGK4cpcg/WW3059kwXzSwgS
9q4ZJ7QsaCY7KU2n5W1Gmi0RUmazUQZVnXaAktaBoReViX6zO8fOctTEZoDi23Gq
ftqXf05n/8cVXxyKVdlKoHUzWwNE6/HkyafQ2/kXThFWgHAxpbjtg2MgCihCCAOt
K+pUw9UrHyFomvd5b3X0Jf1ynqiTKDRt3vZWs2vhLgL0GJOj5g5KUxpUH+lmA9YU
LtPbvQ25Z04GKH27sjBsd/aJj6Ro5ouVMAMWWL61S6d/NXwoVFoi+ZxIOctXIXY9
/DRtWmpUkJEkgETmCZJQvB/kjCRDodUziF7UWoFcp5+BGOBogirUpUx5zDyc2Q+9
TmELv7RI7uuV29q60xFH6lZ9S72WjFRz3s9q9XjuVGOUeP1jvhVYP1AT8ewB+pCE
MkJYv5KphqSEjFl/NdPISeTJFPWCt9c2RSeyq2HNGKDcldH2LKKVwZVQChsICVO3
2Q/xKcUnourwd/MW0Y45/wNbKX9/a3GFqERjZJHsAI8wHwB3Enk4EfT3ru7fRmR4
xl9Q+BFLNtw7zl9p3dIzBq1jsg2eRGdjC/hnHud/Ms00+OSjTeG9hoYVR68mtltu
+vtzMAnhfxhsjaokWqm4AsxmJFwYxVVIVzC9/ofBfpa3s3qk6VvUuZxbs9dVM/X5
e2iTZBjHy9cBJUe7fhcItkSWZCPJNAkMNFQ87dLNODS3YHkdbhYGAoCqp+MULKQ2
RgGuUOKY5IXEybsZzW1CsM9eRL5zZocLdRDK9JHzSjir0Rm013uP+HwAhWuCfozq
kBVRHeX2J6mh9gq+zRLlOIBWnBsWUddjVg4AekL/NX/CvTm3eVznM78ZrH8PptVC
9XBwVCSggLlLwE9r2jUARf/1S59SiF9DCZOD98U9C7Qg/ESjnEZODBlif7cO1TRC
0uYval8LC2CTA4ZE373T8hI5nhCNjvT4p8uZDIxf3Xze9N0l55pgXOCNtNgcBQND
BOcFy7adrsRJSgCiVswXribfo7NdMEBQJgrjy6JrcIHID6QWZWbiQgOaddVEwGIT
YjrnvE2yLXBmPl5A3mDgnR9I3m2VkBhzdYLbjJrzxdzRGXvgj2m+qigKx2B4J9/q
OI3JqRPtJlauoxDU6jPDdgiHZefTCB8sCTqiOdc+kt61Go+TbtwsME3TG9Or1KLT
LZo4YbvwNZUYfCFbr9lY1jn+r493lRwsojfZYFaV8xLko3DwUUh1N935nqd3oX20
1nZlRW5YvdL9wsnhmjX/B33pxTqn3RBmDwwQ8r4j/WF07itSVhPc+jiCfbbz2sqs
mR/jPLqUkPG7elRBYjOkCXgmpQCfj1LRi1XTDCAOJ2M2WeVBrbX+fXGOjnOYPl1V
M+QoYKFArTnXjl4FBY5WaTT081THyqAPvmF1NXbb1i2PNz71za7j0OLhFZCrq8Yo
rxG+WukhQfxhxefkGXStnJL85r/uiX5Uv5xrQaJBY5wckNyn/Ew2ld03VQeXXP5D
iTigoQi8m/JoHx2RMuYzzaQ6CzL/30TVyyS3ZniPaJx0jYR8UNKLLrfSUwlDAbgD
c3UHdpPYtfCJWTdSIISsqZQdr96OW0yemlGm+3rKAWgufU8yfBnEMZ36+n/PwNQM
iWLgDuGvZtHCD9y/YwKGZ4tNlJbWERJWnmWyKO7XyWHlX0pPKEr/eOJjl4ms4x9x
56frN1Vau+LbykP+iza71zJeSwPmE2knBhjskAYr/TYAS9yMtEcRaKXafEskRgQv
Qn98RnfFeFB35InH2AobLRqpDrbQiBFh29NLmpZU9FirKtIoHxty8auqVhrQyS1X
GD41g195HU6azmH0FB+KYIdDizWGu8xFgN0vDr8uTkfjDpIErpbbLZNYUs8ROAAH
wvSGuZnMGrWIzjeVr8jXmahowhqDjYO287TnKG3UhCf/xlyo1HyYgOyqceXzmzjU
gQVNs2UUU3TJ/I+yvjscVz/jXoaV1FTje002VHGlzCxhcoA4URzJ2TVz0CRS+LbA
8mSfa80yiV8HO6IpBwdEJGQNfYCSxMpIXFPMHBDQ1SCZUqRTsVlgRtOuKy/jD6Q3
ezj9uZwFoiRE2AtSiLBAo9lM0an3YhZ8ZkeF2smbxKzjt7r3YZ0D9hhh/PvilAla
8qJRwnYkoUKm3ErX8kirTsfu5TiUl9ZH6gfr6evz5TAyyOfT89oU9FUGTbjSq4Ci
+IQlpGD4RH1o19DZ5aAPppmobGmOdvU6fqTi3ppDH/ybzLVzSxwy0X2Is825K3ed
X/C7i1/UNufBsc7kuCNxlOXBMY2+ElrQgUCFC0wk/5xhWENcap9HtfQJpJtqyvro
XQuQsZyi0xQvfOe9Yqx1KL6nGboHvq1Bs+o4AyQhOI5IxFgqESHVnhmg+Ljlm6oq
WYhBV8W6ojKFlPoQjM8vPCMt/tmV23xLo0kjbeTZqmKttlMXTo7To+PfLQoRSDD3
rSyibA+N35LbSGsUGOYShbCDb7QCcUvW8weLI4miDvVvWTwR7oF+H3zm21KmtS4g
C7qj6jtRlnoMKtxnC3+E1rKW19AU4sYKCYqYaj1f8jVEEMA2+5zuSmczC9xfanFH
hJiYI1kyePHv23YN341gJmSc0Nw7NZN4Qn3G/LyrbkJr/kIQck/hAwO4qhqMTRDy
lSWtdTi8uEllQXRNqEV3Z54GjhwQfGihzd4npM+N2Zq+q3x73ClzyvWF1m+u0jsV
r8mhwph8WDMHFQvRxyqz8J3OrAMh2zRyds+IGGdw8Z0dX6UNVjr442udgj8a9g3i
IhceArWwtT7JdhjwcrxEikOuMBweJ4JCPcPtRSwjZKR+gy+RMXO+GURByG3qoGtv
DhabGFR5DjSKU1W2tvrGLSzghGuwkmFPbUvK34HJ8H41oksyz4E4xtW8QbkW+0V+
jFGhNkXPO/NoX6miAm3sT8Wi0ivCdASH+/j8qTsaUafjqhhtUx1U3wGzJgW3pmR9
lL3aCwUcCeCNVrZCs2/XnAuDd0AmmcR5HvxVbr8sp+vZAFzt4ent+sPQU/xfpLAl
l1eD/jV2426LOq7uVj4yHuCSgpaZFXhD5nddqPTEkoL3y7yWk3BkYmn7IMtKKRcq
q/Pcznrm1mLiSryVnS5e+RfNj0jBh0odeRAHHwCL9XSUuP31RxTO06xpawHmcnUT
cvZB3NMF4qnKRgXdx58ZYkF6gG6zCr+lNFd4k+Q0FrKoxQJepvNv639ABUovslXq
aTCLekF5Xa5zhP85qqA5fiZXpoaVl4QTREFnKxZC9nDdjW+Zjyzhes1ZgkXcl3Sl
uepmV7CPSxH3VhpT3/n2RQZLlGGJHjwoSwmHS6WQimwl2pragTfp+lwZJ6DcqDv1
auuICkbTLVzULOZ4bBckTfE2i1KYeDo7oG+ZlmDa2Abn2WWW8kKH8j/wL0XQX+tG
6cEq4c85gr4YwV66hqNC/VGFd3n7f4xZUSqDgKHaO6SZ1RBZ8v2YHdwGPOyvt8zW
109GDOEVXJvJeRnmHVtW33xzl0092QK6ApX6CI9nUlLvkNULgF58UFhup9imuTF0
1Q1/77KEUMNOGuw+36UX/LFvJknG3KX02Dgz/XxJi5A59I2KoCi3MgjK6trq8EZj
lW9V0sI/y//aiiNUvZMNF5zbPqxjP61BmXyhkl1GMNmgVuD2FrCHWqdhOulT2m7e
9pigGpCR84s96pPrskWdnUzY2LnYcFBll4bmn3n56QLC2IPQb6c8eLPX41ukiRbK
05D/jk2QDwz75Hll1q21EfpYY/4GzYvjeKJiyafqJ8XMbPB5C5G4MhmS4gDZ4nc8
7+HdqFLDeQdqqHA+hr+38vtyLnMQ6kRjsLHhfH8wEcGRWlBrcBBBrkmAuOCHm4RE
I4Kdkglan98EMskFeVZquaRumetYFrvfQQABasUGGThCUh7+u6m+ty3RWe6htZRS
Ey/G7w2M0bbHMRscgkaSSmSeUELJDbm8tvzmeHfw97AoOVWNbrvvrBsq2oZhmo2U
/YlO1BG8QLccBzkm+O7AOPOD0KrMOViIvP8mWMYs5aVG8XSWNq0AJDnME4quzYsF
2IkAmi8mnA7CWJ6Hx/O2i2xbD6coDV5NVSJJwy/l0/r/5qNFL8PBWvvtdijWCfYU
5fx/tttGI6vdNEgFZwgxNWYcevITf6VQ1ws6sq3iHOHvTMEBhgvpyT0NQ2WDa/7U
UpFAJfsMsY8dU83nnHSdllv9wZyFHLFfjY5oXCFo66FOlTPV0dB0R80NlrhLjs9z
gZ3k0kjwQ+qttxThWtZXp9uIncaUS+V0bdhWDZw72+A3t6g5S4gQyoA/ZwHxBLoy
3a72yFBYvjlnsK9RulGIMQDX2bg8FvyMccEAqmo1/UzKYPuf+T8JH8OYm8uZr0Sr
4iUKn5FsO4WklOI2hE0yH/Bnnn0XjWeQQ7Nm4OVrno/khLQ3JGgKjjlV2wOuykmw
47UQmOaqCC91SGlpmPGcZOjUytlRdooTAoyltBAU9z3gqLzNFPws9B4j5juFY7/j
YVZL4RHUWmB3Of0Z+ITSuJ9pfqlFsbkU5XQ5czbJfxTlx2FOZgVd8i6Prc0DR7Ly
zUOTnziigjo5oHzGB3pddKnPNYlZNbZ6qawpYRF3bVUuriH0AeefDWht8LGHqxHu
p5XUoe4DlngUmAMk7NffufJIUpNCR81xIfh4xQIr7K9snzEG80Pt5CthBRFxtvFl
MyGjwDB2ibIbWmO6bbz+QpuR5Z76/qZJyWn5OLCw5pk1iirSsbMQ00Nw/SY9q8EF
p2dKQFpD/FjZOiH8l/Y6ogKKz4o8U5uYUYYdDrpZrqm1eh8IrC0eCbwMVD7S2PWn
tikGJrmuCUHSsCBxoAy8NLtpK2zYbdbn0PBSaJZWDzwC0Px5XXLFO54Om1DWOlRf
mu2K1j+XD8HcCgh9WISvgjwTxECPusE4OR/O8Z3Ep8HJa4QKybgaY0w4hKHC5eCS
KuPZ4JTD8ZLtUp7PmNAJ/4Qdflv53wBa+G/gANIDjuLGsuaEOYyfLr3YC0uBMKH6
VGLOFxMoNlngeGMAYzegm9KV1WLL2BX6bVIGHtCu48gip4T4wcp7IzOUkpfkioXW
VjAB2GMMkVm4iLHt9BM5B7Fk2Op04gfpon2NS4A47UPIfZbAovVRBwSylNMlBY7d
XLWGJPENq5s+3F7LwLEQtQSab2twDkLP1wYvpE488zp5qjq5RtPlOb4+aZrdoD0Z
VTtCIrwY0HeHRh8GD4SV48ZwBvQMKMV+MV7aOzOrtHDWOwNYp47QDAkkIGB8UC19
Gp/iqcuDqLnwFyc2odEoGKofJcSUOZSxrQctQsLKShqTXKo4tRWNkztkDzNihREy
NFyu8KebyUGZpKlGanVRsML5bSVClNxgE5N5xgIw9WsiS/WL1WorfigPifC1yCg6
GVx0pLOavv+Oit5Aeho8MFjfwESXu1HhTp4YdYGyUaLMgo4P89P82Ppx+alzug3l
i3ZxoptgewsTuEPMPdFQq/ej382leyN2mb2lhRMt3nvt9BKlA/aGTC86bSfx44SY
zAqrkV/CJU/rNaQrSRhQX8PGEpLBMddA/BthwZBRsWar511fKwpEo4SWJJ89o6u9
Y04vjPm//pTOsXHbVkeSPbbkwuagM6mx+QX/jVqB32G101k1Y40v4IOuQd4Tzh5p
cZvPoCOF13pAuD3h8ejLVKM0yy2LmMF7fhxCXERqO7/a7JxeNY3zdtCuoO3n5/pQ
d7A6uluMmeIL1Ilwt6FDHihng9sdL9vomYuIZC4LIxqhZfEuQpGM3Buyumale/hF
L+tboVJFEjj8++pQ+PHIZ8t5SkoUrY7Ab44+fjgORrG2s0vgA+X6rbx47Ludq1hP
lweFXuT6ZYo0MK2KOrlA74sPNIqz0aYvv0+CnjoxuZdipXsOtLrEhsWKaeC7e147
H+TrVDuFdl48i75j1pUBIjx5VxRTIO5EJhKgJeJ9QdV+DHfmnDgBSaInuXqQ6UHN
gcACFyf6PoN5yFGGjVQMIsQP4ti/m5wXZCaGNXnwUd8PVFGmX4Pm2NvJZqwoGV5Q
zQwIZHT1jOScEtsIHP7o0UjsbGNg3AKmTNw7jU+0deMg7z3nETPSfXylN0Hu3OfI
9w3d8owCt9TQ6ThlrRF7R8cffBd3mfnpXtztRp+qe5AGUVRwQ5o9nusufxRSb+Ti
oFYzw6akSs7yOWflVp2fN4B4f++6XAfUl4HBGzJTEVZdiyGM1n9ZQ0ZVhXaJ3DsD
j0gzEOIpaGIdtVJOgvOERq1bwsrcJ8zoo6eUREMQ2OG/abHPVNkZRIq7p86wVbgW
iHIowQ0+vVB0kG6oAGtAFECynqtCy1Bh0rEHGeu74vEZh4TcAWBzR29aMmvjk+CX
da1Uf1F/YFOIQ8Xn4VbR6aEAnk8n+Qu1qCkLge5NKvrt5pDxItZA2E3ymkPCtSlZ
G8W4uuUJtCNZwi9QZwq3qT+WBNQgRMJy6+vewwFpFgV92Kl3tPvahFlqmwbEirz7
kA31n60dxxjkgK+Yn5AbgBYXsY9Lilv8cbfgCL8nll0dYc7Px783BOvJpAWy3MLQ
7lq09vHz0nMNrpb+aWSazt+PfyPaLOYa3jVUJFs6sACu7PCheZz6H9gs2E2gG/mm
+KGFZHBaRMFWvs5X5FR2t5e2Eo/yKRnI8z53j5ysix05F5CeYNDi15Mt15ORj9Qt
8CbPuSX4VkefoN2+QU949ScSu2HYo/zPC5q5P15n39nayl8fhuu0KOZAkKPWGtRy
7Z3/+sH/KfmkHh1XufjodIa+nsHLJTX9vQ9F1qk82Eik75j5JqgrkeRtgptvCwNn
2xUIQB5n3bp+rcHwCc9nzXnuPBBIr4a47TD0r0kx1bC/oq0Lh4IpbuNU9TpRKc0f
iXayhdXiE74avAxv7fCEdKDoHT0LB9hkdD5eNa9J+mi1uUYbzeAquihMUQ74zSUk
sVHCbV65UvuAfR4rB4yF9oV6+ykDd0VeGk2/COc/KMiU0/2DTKh1WIqaL70TWx4W
7G78rIEf4ykwTHah0CJnAC4ICosAySO/YlHqh7eqLTvSrKvpK/0clx79lVUfjTb1
LjV5V22SVX1azmewNQ9so501BL9phTFHpQJBRc+k1tNrbWuncX/o2aLT5l5wW+sv
n34e2+nPeU9+uqGqFUM74ERLrVmk/HLICx+1GWMdFrVNEIrBvShB6qQeNUJK/Ylh
yNNcQefnTCi6+PZG3NBjQT44b8KL61EGpNc20UgiZwYRgiszlkv0nNPrSApW7Tqv
ObvqwNXiP4f6oUur5OsT8akj2OXagAIJlDGRtZ2ST9I1Dzbx77Mpc+CiFad44tFW
zy0liCUhLrblnXeChLsFCaEV3T/AEK28Civ9KyqOdu8ojMzuWE+DqLJFB4PByzgc
HYCscPZxeKN+VeWpOmVbkUlm0lyoxbMD5ofRi0c5pbMffFpY0kuNZK8mU/2k+Hzr
rMoavP2xgTLT4TqCA7+2y5dqXek9gSjsB3MRpi1kq7jTHMQE352+2qs/ixFxZVBN
LK0EqEKGsWMJ+jyfex6z8BIJc1UpmYC5K5r+NBd/pu1kz/OCNHM5CN1/A02dcEsO
ETbezOd/ZS/DfpKicg2dBcLnxT8WAz7s+v29FTu3VhWmIHHSdjjbCBfJfSH06kfO
Ptwac8EeIozYvNjB2Mq2PgW0s/2geo3ptSvVQtOWKeOtMXjMllb4J126ZAoB6nKc
DqItkd7VUm+9rWPPTN6uIn37eK0qLjX2E8L+rDfeOBSgqAohrbnliX4mrTc0i/Zh
3FhA3pc/WFzVlu1O64Tf26JT/9T64SGKh8Xl6G/t5F+rBXwkTa+b2EyC/Xxb4g9W
wwhmPjzPwF3oDMW/ZOfNv6EV3KsIAZLSDjTy8zy4OK0BWKpk73FqmZjTxCLMGW9j
+R7zZLBF80CDp6Rr6XVJ1Kx8d2U7blSBVc8d2aUZDjV7UmSTwo/EwtrkbPP/LDra
24L+YpwfWRHk8QV68nVMWicE1xJupkUnlGGmj+cIIMCTvyP6GxoxzU4GIS3IL0m/
x92++0rk50jsZFdIyFVGof4XRT/F6spLSKC8VQAiGZTXRdX17RegJNFEmwbNWlzz
3Hp0NoiFAUd3X5H6+C+rSOhkgv62xV6j4F2kwxq6D1EVZLaAxmCCnjDzK304intg
h04/2pG4Pk6ZjikNTFyGUpxyL8RvhWMsBhS2jO7tQ6aKS0utkBXO6eN+DZxXDD8X
1t7rA/Zd1afJfywZzODmDtcEMDzxP8lquaFfBT9GJOSfD4d9CyAmF4mWPwPLU6RC
AogtMfkpuLvObfKKNKSybK8XKiVz9w3ubx+QnWdnJjFQsHOu5ukk3aATg+wyU0Sc
tnCsiktnRbOhLvyG9erbAySqeW9hlF/zj1Sqk+ikdCQY5oo3DqEm0gqCobh8uY3D
KVOPGGz1+u4uAevbY2/EuLCsVz8Pc/TJ7+vudc3tEAnhjlg/lqNueZwwD4aciC1X
Jl+zA9rOYWwoy6QPpuDlTtegAqxDxoPK5ngQhNCKhsK8p4cktncLnUId7mZx9is2
+OYBMqw3HKzkp/13NPjmLoFxUqIUu75dUcmmbksg3hnFPO2YylTOqMjkylpkdfaF
wb/2QYr1ack4O+ef021LMfyNI9GbDpjHKTXYORTUnzYie1uPNsDE3f15Bz1gV08E
YMtpmDx2g2ePWT6mSLJIgBqrv2MbDdM26yq0grFRtni4vvl95X2LC7u16FBMJvVi
yl7vZCLr7rGuX+IYHMx0QzdTzi8fp9QZWTdGT/w2T/cgPaazjHUwuuuG/QxbfoLi
/3rFXudJ9zdzOqgQ55My/wBOM8dXFT8xr3ThAzKlACFjgXmLRFQizxijXh4Iy1E8
WKJS/IO5eNRE7mF7ZvDMCuF8ceRysCEbc7ZWaS+lzyz9X9TfICp4EM0cg876yBll
K078/QAHYI9/szFdymZA0uqkSOIGNyQ/OkxXbkxvhEbovRHjepGGusy68D3DW7kB
O+HYqMU/jSaAoIxhBFIo188eciD78OG7bfB/JpQpZYwPkwVpVn8+lgr9r5OyMHUH
ndnZjvne/fXVxhjCzRnmL/fzYW9Tu+Zcx1TmcJGeEqYPEU82I4PCqtXJDrXwCAs5
EGkctgR3fUK0u41cN8ryAoU3xJcfoma0Bj/5fhCTnF7noCOWm8Hmu9H6d10YViLT
EWqzCoinNgxhb4tYpdYJCofZGuFdEMaosJZZZyW0cheu+x+aNT4grKJ6S1pI5fg9
aphHGFoQO/X0I2IYWFwjRPYHb1UucQHTlIGs8oxLZuSiHEgqkvQZHCxSzXE5vA9Q
PoW9Xn7GYGwCLFKnkGPzkzE9JKcOKF2NLLxlW3mLP+wlkOP4SScgHXXiuFf2KvEd
KFhqiRTCdRg1s2Ss7BrqoVXAo5fWU3B88DcC6JDImpuYLJ3bU0VWM6w1rwrVJs2H
zfmURd7i7PtUIDIK2rQql19+hPN1sK73O9gugQAU9+gom7RstO0V7+RxEzBH/CBP
Qw9VLG4C/4UhPMQRg66zyJRy1iPkeEYOZK24pTr7QGa94V7/YIvX/6/66pX3oXzZ
oQx878Mey5QgfNXZF2agTOVEldrSPMWCy7KLqkbJCY64KZ9c75am6JqJHqATMKKV
GCgOKgkdfpWP8gS+52BcELobGGfEMTxWkpXuTnhlWuG17LTA7p/45/xBElglL9Pp
dJ+EJOLItAVjf1dQ5y7zkwHGrlFjEKQ+M0EYCrNb4T5vADHLUGZWAY/vPDsgdd89
mu7JKIQLPY+LTKA47DU6PpZfy9tOFvXkGDUSbFbkZTwHrlm8ZThMxnSgnrJbtAFa
XT1ifM46UcVinxxkVChYSbQjGSNDrAaLIqNRqQF3GGjj7+yUgdmmUPPLrJuPm/kW
87EmUVlPDU7rnvCtjecSuf8GBR18/4ZZ/wzr/7I284NcGnpDQpMe4uyyUBHNAZ35
P+7U66YmMc8iaJ7yYMkzf5sCgNXTBQfK3OsGfyAKKz6i8CBUas+lBeEQojS0TTzf
7ioKK6RQnBWTG27FYEoOq6hJH4tUBZK5BBjTsrbuQMp7urGeMSEwXAPnXdpXMT5l
SCOrLsxvrqZEg37QQYdXZWvJo6hsf2tUHO9so+bP3Kjt+9/OhQBNj/ryGHwICtIW
7cACeo6tkx1BOEZv/lb4bJZkqZKEemBwax5Qwg7rBQqf2nMnp1LMYxctbKXSegM4
8mrxeF4jZtzHQcYeC6hOwqgRMGsI09fpoYJ1lMpRJnnqm2EOylEVehF81dMwL5Lh
oJYNjcmi+67b+bOej4f+KiyWbbkGzdyuMHxi7MomZ61bFhnnBOBw1mfTP1PTbQcj
u5wfGtdruOB2EoLhSqgC0R7VfOYR4WG1q94H+D48fZLy05OoUXGUr1SIXA0mG8iO
8c2MEIiLv8fDKhtsC6LjGnzkWDUChgGa9jIsrwQmwlldYtoDohISf++00fW4HdNA
q0a6JCgEs2w29UU9yvFDnSDeMMj2X28bYSNKNPg6sRw6kjnTs2FeFL1Jc8vZjdSR
BIBRelacx5ffTrioK+IKAxOMu2RG54nllmlHS4Q5W6cWhGBp/q00f7kBD7bOlcBe
IxrgaLvBDz4r24h+EN4nnHOmUiUSM6mKZ1ADOKTRwjKLcXzi6OE7nbIZf6mnIDD8
wPK6bEeiwg67sLyUATFHsup5tQaeK7fw9kJRMwKR1ZFIKTMN2ymIQdhK8vFwBoBK
wh7q9sz4VeJOSOQM1ij6zbT3h2bSrGe6OG/dBfSEBMAnscum25t3l5EpCF2yi23R
j5THtxMyzNE1Zsq8eqcP8F9SD/u5ajKfLB5op0KXd+calvFhzgqFpnExVczYfSNl
fY9YJnmmqhWQpRX2Pba2vt7c3nd5mkLdpImNC2rI7COCPWx6VNK1WsA1/wRbDvbs
0xqRCuZ1UgNR/G59RAcXKqQ2Fs3/t1toMT020x5ZwgbovNbDbg2MTE9cObwErsC0
iPd2RSrqWTV76juEJMm9rRXjfZTOpEoXDdAKRI5m/dtcVDRAfSQtyqCUHeM1QK6b
vS92X44Ui4LQlsEWcVrdRCbqJEwh3X3QdPqze/X5rANKChUzBMr+8+3Wp42wN+8s
kFGfjlHWqYsp4WUZp7B8xkgN4Gk4x0Ti9oI4OdIA76DpcDI+ubDuD4+DswAqAemR
Z+4JIHLmB9bpbNl97e1SAbuzHp6Y0X4RxuB0VRrblpwrJqUlug0iss9IzLoSmbPb
2XiOmjsEOwEmNLdZz8V6tUQG1IC+yZmwEPJ6MBh+DAOsA6a3zqAJoWqZOTCDefQY
WySDaAsAjTIno6vlL98pSmTsgmrq+CwKcjGhC6Hsf7CYRHHztOzUmcoMZKlL32pA
mmRUHfxXsJ1R1Quqj2U3KsNKS62iPxilIKWEdPEXBr/pqs5Vy70/7F8oc2CmOzJ8
Geu8kuUiyulyW9jfFyaYYZL5JYL+299sUkGQidU2GXF4dVoIAy8YWuXeuw16rCfY
OMw8MhTaWb35xZoiroiSAJfnWwlNcbyEi5cHI4FG62LWnvv2SPVpB7zXsATwmHFk
2EZhjH+uDrq9tnLw5GmtFO/2dfU4Mw2Cp5TAzAv51Rx7AxolGMztyiqJZ15GYV31
oJ3pD+Oq2Qeo7BjEHeYKL/XzGynXWU4eeGkDSJ8lonROa4NAP3+ZIR++kt5s+l1d
Z6/KmeNWX/RipzlES+pjHNd6Wbke1z/S3C4JQNs7+EwU9QmH7Yvf+FFcBwVHvvoa
sb7iFLn2BRlsAO0EiY9MVeFURR0N7pGLP8I+JHQK4YdWft02J0KKMIdHtt0vCiNN
XKFFWNRHDyLLruP6jbdlLcP9pITEdRXoKq/FttcU4G1/RQe1OTgWhODRWm+S0c34
n9aGZjCq50ljO6eG3JoxdGpRQ9dBmY9fZySbLPcy6HnAOICdanVfN6+RYnVRa75+
8boa8CS33XG7CJRxQj5ST8WxWcw2LmGnTtnwaVyXw7qQ3w90QazbOZfhxVvhYQCP
34XgAVgNR6T43SzxBwBbOzRNhc9IoF1eC22ZbcSpGS+xN+2l5gYT7yW+TVPxLi71
VFO89P4iieuTC16V5ZC4UBIieUCNScy1jkH8opAmTupHPss8NjYP1KIx7PB43F3b
oPh0AGcNg/L2uudjdOKFtnCKVsWdYQH1l6LXDOZ1IeBEgbwAIvGxFZlRxJ0sbQtf
OXJspEKkUYOWceQwF0MxXGg2GRTrlC1Yve4aiYbwO9yZfVZQY38fFvmyvG8Um/Zu
MBmBLFj/7IIzVE7zVnKbxTYETD+NbHzvdRv3zCv7Usk3de1dl78JPOS2Ojqpy5cu
Bllqzb0LXNjrr7Exp14Ad2mi7BL28TolcEmmx2KxMafxjUeAP7EmirG4+RSXP75h
8s8jeRgqqq5PxwPVf+Be0QM8kAdki2WJw6y9mhJmoH9XVOBHh/l4siOsLGoGcYid
qCuvMAlJx+XliYpiFoABYVldvgOtVMRz+vtC3aG4FIQSHNMCEGjnEDpVFIk8DH2D
WrzvDrLqNaHw4NIvRB7IGLmVIZp0tN6Eeikbw5BHVcrEmSGj4d/g6Zk47gSde5qg
7qQSTeUUUXLJLFNbr5hnaifd1wA4KWIhq1yKolDMaV9Ys9DLuPWxumCR8wy/olWw
zEUYUO7FeWxOTQF2ADAPXyPLH5smf2UDhxbKbWdQq/iTwX/YvuardbXjZ75GZgyz
BBGi8CJioOmJZrG4uxHzqAtT9HIz4Y7RmTQ50huPLvmqSqxKR8r6uNaIAOjj9mA4
2oU18JnCU1d2BIg5z0sk3JD6xI5vOtdQy6WPcZ0OTwVw4n1+DjlmElMGc4nHtztc
Rj3es+SIr6hXwSCvZSWspOtdpmOJwU9HesoF/gtv0ZnP7hs9PaPNtUcpW1rUGxzT
jTmTxRiNgkxjounnVY1gMDvSHS2AK8KIoQOQp4T9+5EFtlWmLccFWk6X4WE3LUFU
RnoU62iYM7ZRXxtcoeegKxvmr6Kzz/Qb5seHjGLXBLOLgXInkgiYqxkTFWcKrBKt
T6+A3p2ewPVNLCvWDTk05qY1qorZqPXnQBOI9j5XS/HhgCqkD60Da3gowqZnvwgf
h15WU+u+rzd96TXxyVBvW/o3dqBgpavHeCZbobd6EzvQwKayjmjeq2MYH2j79kQR
byOUDCLU6tN7tChnr2wRpHq8/lWebX2+BwWCGqzyr7r+85hYLd8ENh+QN10Ba4na
ppeFZFwCJbe16okVee+m9+OizVK6iRLoME8hHohra6IDh2Fk/2+YPLzLxRU/hBGW
THSOHYd54dVves9OZbQXMYvV44J1rrXhy4PX/7lDMn/54cixvs248Za08FBVtJ9t
s3WKZAABEER0ZpwtuCzIW5jFlGhXq7GCvcoFJEB4XliVKYLg2RzurCTP6mXnZL6X
DoLcGTNNJqx0cirPllqg3uVwpLANHP3m7dqtQA2C5uqu1BLCfgHqinqvXd3mYuaK
K/W9yvk2fq72Qr5pF0zU910eZHKuEEzGiGcHklIBtqGjr6ZqZPkDJvmVo41M+w8j
75LpX9usPIF5nOHIjQvCuj3l5lSegHVeTloy9IR6n4XJwo6pC1/8oCg7Gagt7ZFn
ZS3eaeYQRBARnJWVxC5T1BlWKe6cMcoDfsacT+ReV7r0JMQh3ulNMqsZnIq6z0Ty
VIcxPer4SWzE9DfRWM3lJvExSj3zGIfr1mdnDGxZ6Qey6ngY017rW98GM4xf1XT3
GYCwcNEOMFTM5zXkXesOnVBvtvRrvUK6SEs704vrwSHRvHLcGitXUPX6fKupH3rB
mV+3tOcmSQ5dHWRIjqO1t20kfDTED2NfY6ZxDNxulgn6n7XaevoPAWYG7kOXrsM6
0gSO1RR5jKEvAMm99fOWbPOdKckh57f22BTr1fbCjPO8HucFtFDYQUDAm0VaUQEo
mYIADFwOdhZBo715LhEU++x+8DVwzwRqMgpzp4U1o7vCaGaLioHY3KJ8SEP4Kd0L
MQ6vZkBTXkVBo7i0VPcdOfPXpiuZK1Nilysp0v/5BzQ83QwiCnDwRT+QU5tUscud
GQL3cpq9t3iZF8gSnhU6xnrpD7tN5BGmzvIs8q/6cnV0ypnE40CQCq+MtPkKExv3
tS8hpjNDfmyeWsrhZx9Jy/hlhNAmcD9eeBG/x73iOx2JjRDDOENma6CS1d0Z101K
DsR0NMPrTM3zJI5VMPW0p9qrchqlPoJ1iqrQyt3XNk1bP7tL5IY/HvFIe79gB6uH
usvLTI75hje20PLlZAM/TRBDHe6586U3npM2/mhnCeQh/bRUEYMbXDL2NxW8I6gd
pz39c0O8Nrr8ytZSZJTx6T3k3FK9j8lQONa4B+uY/4JmqwFHt6q1TywVZlte4goS
HZJ5K82Jjxs89rAEBx1295ZQbprIHzPU9KtPD+8J5QXxOO/2YC74nHJRAOuxa3YP
oaCI1xN7SvAUEU0u2v1UOXmOTKg/6LvSinHQaLKiq86F9zKRZxzmdyXuWwsvRmsC
nXMPGE0lWNecFnkIjLiPj3kd+qbwSXIAlEIutVUPcihaZkyjypPo/vgVdwCkOmqI
aEgkPDeo6aH/MtbG2ZXB8KgNWBX13ACFuuhmRtYPU61rMzzSbfm6bfkZ93ZaZvcb
ZBjvsQzmgqEU6qHungOU74QTbhDrH+fu/jZAPtLbfb55+dulnaraqK+gcksebvzM
kDSXR+E3rVJeaiqG6vbg6wVJ+kkl5j3ElyxNUsy6yRaq1cC39BQmDdjvXJhMyGDo
VqkZtfRwnuQVPy+joi8OFw544eFOjgUH2OH6H2Db6ZN5RrWkUzYIIEGfmjij9Ow9
6S25hIJ+SQMN56DnN28uFT8I6bQyTd3r3JkT0tG3htWCc9UoSo2HHfuzOtNdGKkJ
Fjj21Gic5H/OK8xleX0we+P2brgSMRg34B+5hirfVuNtLZ103GMYP1QiBs6PLvhd
WSlcXFzkxEyj506xOyh+IDoGnDLbP1U5qCLnkiMBCIzTRREr7kO2I51pTM/3Z4Fm
HvvK5+n+bfmlUendclyJBNBev9GB18nZbRJZ4/sDWpr356dA51au+5kbCQqjJ4D4
Ls/z1Si4RoYBorWYI0yqRe2U65Ms3leWx94h1ySTs6bV30ESCdW4ll213KCE5Qs5
qh379qQ5kP661RjkXr6r9g6Jvot2phq5U1V0EDr9I6m1CgIVbjQuH9nJtNtzqdxW
JX9o8trKWeAAMeuIPw0tlwzTP2KqdS51qUMnDXP0/MBzA0RHoo6WK0LjMmFm92c8
hT7avAVu2jFR6zCZ8M/xmyYO9F6WFGVGoU3LLwprtsGBW7pYeZ6zZ6sKQr7hz3pv
ZbHk1My49SORxclo7M/fVNcPCTcjTTZXJCjS5OflhGewBwsyO1EBYiF8XiTRc8ev
v/rCH39QNcXAdDW8sraIoO2YHAi4aq9V1qLya8HlSpOK0iQH9L+B+uhKKaBf7U2q
bwjDYqop0k586WKUY9RaoUEIx/0BG40xj6DE2HPYWm7svfzac5xtZr5nex8PMHM7
GdkxJR37RFi76+BIOTC0OhZr4mN1NAVg5MzJh/NUH2qBQdsGdnNfENVvjNuDlzOQ
QqEuOZ469tq4rEcXV02Vn2m9apWn4d/PiylrMWpCxzZa4BHwqlsTb6Stfgg/M1Iv
Lpu9OCopzDO5kDyfzZhwjZ1ILAxn8qhrp29yHudu6uvGHi9EAY232AcEf3UrTnP+
/y7tO3uaKMUA9RwOL0pXamxuNnKzTzNReYyAK25jZYn+OkfVF+VJY7/8plNxoe3Z
6EdeYCLTRoyIxYjOreaAssCq+WwDhVYdXzungJqRQY5Fux/6uVJZsEFGdMebmjBk
KguSwC2DbBiE8C/LtUXzs9VCQH4DPA2tbrS6B3qcPItoa8u1jHGhegB+K9jcwk3t
H4Dj3iGCaAcRtfgSmLSV97ws1sSheh+pEyw7yWMYgA3MgkI9uDuBzTI7NalyY/wI
Av5wO+a8hWnSEAph1fuI3r15gUxILPe0gMHBXd0f9GmlxfyVe+dWony8P6r2jsWw
2KZiHliHi8OiqA+FCAzUVCwSzNWchQf4XlGNiYULAU7szFKwe1R6sGdeyTVvCEqH
VdANVqlAcItu4PMRNk4YD3ZtUBHMyQo5cH0+1Q5PxlgkRPPWN+OrNjlzhuO6nozH
WUdjgl2OJHUdMvxO3AW67uOlM34TTViV5irPKTQLuOKd5FF5okChM2E6YB8JbhzK
sUv30QUzZ9ZlUc20aFmM+gcEzP0vXG3jOGMdwqWNtag+cXFusxJFqhEGguaNG6rS
pd244sEY43ua85kNFXCiq4b2iLWPuiE6WdAYiD8atB5KYE3guRQppjfDoGRie+f6
hNl1nf1I2tgo6FnTNkl7wnwONyak0S09iUQMzVnP0dtv7Z0beQDKFTAs8F7zqfoh
U3kNUlkMZZQvwTXThGqedC10prSl7cN/qOpuEV8OPX66JKsQS3LMhuA0Y0eIw4fh
XXT/Aku4o5xtkZ2w+AOITDOEEL+DuWM/F6uMu+gQ/FLlddaFMhTOm358/D9ZrQZ8
KMmcXF+/4zgtj5/KWGsLf+UU9jrezIcy8hM7YJFqm4nKcQ3LMYyu2OjAnkHnYkxv
rgctoMEEOC5+ytwy2+njjnrdrvIiFV7Kvt2I62s5qnSEsgFbwSI5GYXfoqRObUrR
NTHq0p6sIxFRQ3gj3WG4OBoyo2xgmtwbVUd1owbtQrBK9Qm2sAs7WUinS6OBc8fA
KKfrUHq+FnTweNFd4opstgghbiGXIFr1gItLDAudtHgOMWFN+wdUeo+73j6bOD3u
3PEZellNS1vGcHsOwVt8qeK0GWghYrHwFHATmBid7S8amZAqcKrD1zXzAiOdfgfD
/cZyAZ9mKbvSJLxvM0E457Z6Y0Rx1EdBc9DTlI6wKUl9FA3V3WRgQTkcqDydUBQ5
HazQyLOmUhIwGS4Nb9Xky5fN0agPBmb0+2DOcuOgmk4rEZriexRC7H4J1ZBNf2zS
PcITeHlrESTMRYDJMzoHYh/4OdBSORQMUVcrjsjfLGrX2zy1iU/xCG/wxHzh7Uep
bau1cvSJLHWhNHYlKCbxDH19b81JkuQKZBneMSLTgXorI63SIBF3TA5BJwglmCwd
zpF345UOdN7Ugen8yxohR1Naz9DV2jQX3lcgQUmtBbMmRd+GuC7xeFq30xkfhYIi
aS3Gbk0tDkHTyoFA5+ofwQXsYq6H0fag6ipcpp84ixy4kuh7OCD6tnXD6sS3OLmy
EGyHfbpKuXk/kbCjw+W8PLOqY9sBSzeRFBKmRWiPm27RsPvLlRndp1HmVgArkp5a
Co/bROoUwZ8y0IoUtcNGmtjosNZtNmh+2UMojUFmhVr5Hx2Sh0SAks5KZMUFrOHZ
RNabIzGzR35Wc/BMD0Jv4X/qdL/uA5nUXgUf6bgt55LOMc7KSd8Cg0SVaTpFD8gy
zS/gkjFp9uF1DHeczVgzIarnGN98Cu0GaoYlnvtrig2nYM+Z998RU+5N7e7cuDL/
FGMvJkHBx+0rN4Y9MLQ6lYO1mSzKF1m/MdUuwZDi0+CcTTV9HYmKGUOBmCE+KhSe
8KbivoXU1UlOhILkcTY/M8SQUkKFqcYmc+gSwUUwOwcf8VMi0KVMp8givGrcPamW
5m9Ol7p6EfVcVcj6hdP2gP3TSLRjjTIUMVAPSkBlT6q8TSGwHadIWjGY4KwUMLQp
hdO9ejm5+GWaRfTHX+1H70hhL3a76UAPdZUCAHmrRTff35R2F2q06/1FNdjTwcpU
jNTDf5cIdP6e0lt8ws/kOw4hAx3ZfVttxYDFSyhMAlYj7eoMHPZhmu6oDyts/VSj
8vMxDbsDbg69ZBRYHrESQ60icug4f+UJ/EJbQz3pBl1G5GQ8iZnorZ10I0GnK3+p
JEeQCR4I1yupTWm1MJSTYmCozwsSxnGEJpEfH2Hrpk9Pgmh//o3hO68qeorGO8eH
/D1Oa+0bRjzF4vYJxh+hfRasr+v6wTUZFtNhfaep/cnYRRfzxvMU/cMs9kQFhUUh
vxyFHaaFAz7i55M3yON9hNCQatarFzwEocmDYc1u95aaR/NN3bj8Cvm/ei+h7z4l
jUoAOvBj3iPi9SF28CBLC0wVJBj/qu3zzHBtHfJdBYO4Em/yyf4VfyWQs9Ub0qvD
oBYDfDcYId/DvlB7VLVdnsMya4mta+R3CS3EaaGvmkCQrkeSusSoiWb205OTaSJe
LOG8G5wRdTE454S1LaXDsVM3HEWKuTBlGUNtTBNySnO9eI20Y2hKDYdfZVqsdmTF
h6+v55Y0kjHbh4zCVaoP+VuIW8GlXbYgeKdERfkitEahdbH/NWvWVL2OZ82lHrjH
j7HTuRemiOv4PT0qiOAuxVu3QhH5mX8QAoD+o9hVnNXBAlUd5kYts5oETIxYRTIg
qtovICH/PFBbKTohWPbqPPhxuDW0UTR0YOZ7y93PTy8zBLH4Wb2MK15lh+ZzOweV
CfU4gVJjjTMCy7e32oTmikDNq/v1FxQ0wL07qc6FyvVkKr6F9a1daFCPjibnR786
MScAi/8yMoukFZALGyswvdD2RYH8a8+6e2olVArk1blHtDgOGqnTmqdOsl6565C4
5z89Tzs7SyiJd1dqhuDOUA+FeSukBwGJ5u+5sU9kxLs3aK1nNX0LUriVQ50JjoSo
UDlLwDLTRkuxA+sOYjfaJxOzj+uIaIiVCl7jTjNdSuwLrD+RNxiSTqc7Kz491R6S
yGZp+N/kHJeNgqJUQKAbwAXNo0xp3YIfv3T0BxgkrgyacspfXTSjQ1+Q7n8a7/4h
R//MouigxnjJDpDniKGeLeFeEpM7lRMWE9XxKD12Ske5yiBahXNtCq3q+LQv8wqC
YfyEf0mDijUbSjtmrT7GPq9BB/7mSpd6T8hyZyD+JpusGWpvwrUvZyVW0nnoTi2m
kgRdK7T6Net1d6tu02e6EZNnP+swdvzdJc0E/eWG/0Ndb9YkBUmEw/AjA0NKbWvn
qWzGP9yjiSokuUMI92V53zlVC0TqqD0+qUJM8knBzi7+tXnc6eypOSt1JC8PQNDM
E4a1TKuCW/IB/J1w5M+WXmlxbdVdxE6AVVuBhvtj9omqBrcUJ+5mwTXlRIroB6oD
xA/Y9zfljVsoEWQzxG8aQM9g8lpWfyPP/81Q9wBkmJys6SC4Xl+Uf4XtAXr03stf
L8a+JfC5uXJPv/ezlx465FiITBj8DZmDQ+7bsvbbixxpyvZ8e69z04v6Pu6sRfd8
ck1YTXZL0J984DFo3eEwgTwzIUXvp8z2EKs8ZddlOfQSWW9ZquGJdiaoYVuiAEk/
86T6DGrUo7kWewV552T32jUdDij8VONMx6RCHJheaZ++WOnGIyUEJUOSJAHaU+go
INcvQDQSQDVF6Bhp50WnZGAOe5C563s0dvXTBc6kgfp7oa5jr4psldOVAxgaD0fn
IFeBtq5S1hr/w3KUKdaCSdu832MATV0cB9ChUXfDsH6Qz9IhTDLWVTgHmIcYdi4Y
kCtzSl4/r9UAHv9ZiHxT/Mzo0RZGyeSaf05YZzfqcoh+mCBL5jDTBSpYz5+MvIgI
C1WUQlg/bIlwrYfZst4CQSZpcWcyqNHR9th4j0QGGDHFTFydNlDKl+GzLyASRhz5
hu09oEb5f8QmhP5Xq9EGBI6QZhZuh60/fbQtqhlRV7X4bQylKKR6gb17wyXprjRm
Ijz1HXJXJiYzkKTUxM/s8wWRHuesxooz5T8aZigvd3sx7y7QbezYnRx0ivm5GNZ3
KP8q48ISq+8L5M3/FqLLkQCEuQSMgKfk0G1xcdlnts7pW+oT3FuWTxlT9N/mvTpY
C0Ly3tKhlCi9pWthyC3Kx5gHECWq6S0hFbkIPyb5bywrK1FafSEcHU9y4vL5Pe13
UfWYcVJlFyLgEdnvdaFrJOSG/afGDYlitAEW2Re9VYK74Sy9xUzhminjYKnoJPTw
LFMAZG3vL3C03zHsAXGOi6vRYKDPN2xPDtJ15SuizqPlYoUS2gtFgg4dajVhQtYf
jhqG5OGINvBgJhsCepTvGsMsgPJPxSvrDIqSUUr6E0ZNeSyZB5ZR/hRtryXrsNZV
q+qP/0sPxAF6lRVEqltmdvSXrzZNGQLsy9sLFK164RUBgcT9ydVlgRh/ocE4VcMq
/MfxnMfUXml10X9AtJjh2tl6lyRyAKhtFgzMoLzZU+Gpw3we2KyCdGCxU2uoxVxr
erXpYjqYkP8M1KEwIaTk2mrHMwQsr+VJGPYWmeserZNYU5sqSyzK5VffDw9yL2b7
utKlRpZUkWmIOXv7/nCWuIKCAFVDgXKXVXMB4MPQxy60eawPLuuJUW6fCiPrCeP3
6SUBj+Dfd7M/0+s14E7GmEJvb/GpG3yYTENF+FbwGHd6ZQ2SWmOy+AV22Y0xuz8F
wemcicQ39w8CVx2j6j79BAbOfMM58HxFW1nO+8XJRY8MB4bphFT22gnxja/Tudfi
aI+T5suENbD2tn1LK2eo1zEHQrGVxLyF5SsxAILAO+uRoGahJZ7AJqrkgpBZwlAC
VMiOtFs6sjKnC6KQ5y08AFiZ63Dv3xJSygMF2AKH7ZZst+i9ZDO3QBG006FD/e2Q
RCXg6G+gsxzveev0oBbw+d8cW3qAwgMhO/RiEH+wIzRPdzj2OhRC0sLTQBfTz9md
2KzL6ulxHIujmrOc07X+QR/UWblwfF4OXZ8hYJdyusP8BuEzuFvHBeyk5HEi26jc
i3nam3YhdWgibaCDUHndGnI4Q9YclzDU+CJ97TBXQRrUON+ceAsxgu/955p9kszB
+kyzEBysKE24SxrKgHEjTCAZEBmkYagkhq7ZEr8gA4+9Cop1GjEPKrZUUOu3bE7U
48l35mrFtXwLZwuLLcIqyy/MOy5bphef6mykZKK+i+vtASGCYH+iVkmP9ncdGhJk
kjkqi8fT77LiAnDVknpQsrYdSNq5lEDadGlfu9tIKdnV1v8E4azE6GT2hWBQTIuG
d2HX1b0SgcM2tBzfRqi0olNu4g6LsM60W3ZyLEzbpevK/zaLVuFKCKPd7bZdMAEI
cFWp53cA18jZFJSa82Kq3+gg8114NT38B6oH6nkHByxzBDR+wluz5RkgeNAaiKNP
bN2ceJLvUnz7sH2wO4hCGVdEPBBlgBcVZPuOeNFUFbf++zWepEljFmaOAVEzqvY3
APzifSXL9VyS6TYB+JW/4zEsnJkfYlta1hNZVd0BTgSDeXmsjJvBItl/1KzuMrVx
EkgxVG8VhCdFr2prRzMTsAZGGVgQA9fqUMQlg2AGbYB9BVIGdXlWjW1ZW4CiC8ky
OCVfKgi9g8XqZcuHfTXaQoXbn9E2J6REoMY129bIWRqLjcarpYYFUjnURLWguGzz
BMuvB6BpELZLb7sWVOWD7duzLJh5RD2WKZ2iDgEhtGhgrOWz7PwAB5BX47dtrpHN
7AWdPJ9Dd9Vmnx2D9dVZ9jdcTfvVU49ChYvidSuslbc0Bfvl+05LLJ6iJwv8CzeB
IXCgRu0a1eEUdPZcda24UBatw6MlqzbX3q+5pCRX4GB/YcW3pRqd8zxb2XajObvN
k9QHQye96tiR9z/lOGyD37anlwO5eyiuu/4w/BvzhpfAjNxKI3/WkXqsRdbtwMv1
NrDEfCEMsRm/XBynHjMOzYMBN7eSrjjgQoJOjUncJY/xRSeBIO7It9JIdlQWwJR8
3uhCTWhr7SXYdOh33HTB+uaUEvyndJlVI26i9o8t0slky7BsCG3cGnt9sd2zemqQ
F8XGqpAwdrezT/gLIRcvwxkvXm9HHZw8DPLC7hDyKJu5r32yHwGROGhMIakFKrTA
jb2FKHg0Z584OBQmk/SiJ7Hmm+1LRniEj9s9v8J9XZHxKhibxiMQBMNpoiovyQsU
G9OyLtjHGbS1XCqaTFu2krttF49R2XB1el/CcPT+80DIXbHRPJKcTWD9wZHW+j3j
g6Re3U7KBh/RUlza+k3J5L4f3+q6SrwxOnfCMsGOT1ag6d0YWKgTdCmw6fYCNOSX
8WjqYMUQKLvveE46QH+jvT0/SYtQvMe4cHGQoGM6oMzxJeuJQSvwP8WpQjyk7mgC
nvzaeTSjzIgcds+Swcz/UJWOIhlDjrB5DUaxMjtTvxCK7Ezx0sbAKXCu4Z/lhUs9
Fx3ucfwqbwxSbnu+x3Gg1m7JQlk9k8Q+JXOXv8syrKmtY0IPQh62dyIWKS7EUXlJ
9hA2PqR985trKDE/cEfHP9H3eEwrJSocOX/qKkBXa8qhUvP0Zrg2ZlfO3WUomwjH
eTqkcq64+rwILhUKjnZd+BXXGMXKx3Rp8DIUAf/m/HFE2byFDXbcNYSAjxNNA8qd
h0I6ZgMXfMRpISJPsqjtOM0WY73/1GN0TyWSgGUHlaxss73LRA2yaTsp5tM7RafO
nM2JbKWquO/UWwB0hOg8CjGdXl/k3Jz38BG6mZarjOlm6hxdJVoYnM9u7jhOJBsY
ut/E+Qd2DtxtrpN0leEKXY5CX0BYiaAkSGLFszq/3FJbomwy/B9cZzHXMmS/wt++
D/66iaV1snZxbxp3cVYi9vmcvnI5MFcIlP7zzlRGPXDdh4vw/0ZHexFxAH6R6cle
MeCPN7mU9iy7SFBTVw0JmtVREXOG3E1cTzhzjtvI3t4VO3huzza6yo2y97TlIQFn
BbA/1uekHQ451lRWLSgF4YfLPxUNQhNn57qHaUErAfpWKVqMgFV6PZpYhozXdbO9
4Vg6R9A7nyzksygwX+7YlC3HYjArnQzHYgBKLRafJY3fNI6l8nNFmCqnM+A3SdjI
aDaN3Vdl06GtXy4gceVJThR/QFhDy/9VLbLhHDkPLJ9QzU3FGmJy/3ISaBKXeNFm
oS2O3ib+bkG1VewZjtDcp/4CHl6k3o1cG5JGmx3LoEeyKjFDKpjlCY0bFsjbG47Z
JBr5KkAlQNx3P6WmPiJI/Ar/TvTiEId0TrNpjCLqhYTpsUTz223NkPnCni4zHaoD
uACIbN4DKA0GB8YRoWHTcc2omUgufyWAiUA4msbQH+arFOiMrnoX30/+dvMr5VY2
9RtNlk9HFOmDMZz6j2Q23QIGN6Kzn2JzOFKUA9pb3oC1F8GVfGF9V01gRMiGrfF2
UOKPkMwdMbmLAafk6iwfh/Y4exRjR8S+xQGjqboIa3Fa/gAo7OUKeYMKxzN8Z+dY
GkFSx29/t7O/UrtTczdfS0ehXckwNqekreByswMPmUF3YEoprhINvuKP7xOdSBww
qtXDW4r5Iqd+ne6j2oBZ6o87DLJLxstiHFWwGQMrHpVCKZVrOdjKjBUt6gEvkq9r
fJUapMKe2n53EB+VXiKwkvpwP3WKuXNKbfsfXyOSO+IwaggygCPl+oMU+Y8rO6si
MBhVYmpigrOOPYVRApXW3E+UMnibdg+Tx+lDR/iquAH21cOput3TJhhdcE+wmg7x
da0ELnYX9eX0gbp3FNImV5WXRGVBY9/qRuMY9TwJVmXriHbFEN9LcnnrnILRh+yI
nsVjHOJ5EJqbSQYNHAMQrCz+kF19h0liH5NtyT7pJCesmDFyz5yv4S2+joEs9/ar
XfXD6oVifiANMgQZ1b9Xa51B1szN/Nck/92UhuDwczlf5ytxd2zpf/H+V3JeMxP6
RbnqEiTWm5I89olBGCxVQPPfXn9uErvqcwtobnQvDaiKYI+tmQ0dhHpuU5fPvRKs
uWt/iTxGFVsE1pe4EmkjGi+x0ECENNR5mMzM/I5Ajm1emozhknikvqGk0dl7qabe
v+sGIHk9qdcsC2isahGDhUk9+0cC/ohSZX1vjeArLT16lgaXiFJFHzVPQkrK9gXy
Y3eWo6lWFwg4gVdS39v9hbrOwRiKtxlxEmw/cZPzC9VInmAbcQJ1sLoqzc4EN6LK
z7YEM7mzx4dXTnqP9rs3RxLgNvEv/OUg2AcehCLdsay4KuRC7JTIuczmOMuPzoEQ
I8hiJm0DWO3v3/0soU2xki0JQBxdGv3dXlyeHsvQ9E0p+qvPsHNbk838+4dQC8Sr
g0dCAtVfa7cW6Quqa6EaHbc4EsggCVMgTXyvHLFkRg6dnAMF6nuv2sTaehGClkmc
DlEcV578OMaYQ/DulW+hwvZZ85ctRfBghvqWusj3xeTkOngAbm6t48FVcw/QmNB+
X7NajyAwQduy2Fg4O3LOoDA4ZmNkpmmY27emMpaMLWcI10AoKd8r+qBo925Ttmoz
W4P6BCAC3+iVUUKVvoiBpjYwtD4L2SiKLdNWani60fbbLrvv2uASE49OS8lrfRoe
egdXtkQKEsAtMzHrHUy7FiGKIcAJV3BSlyXUHn6eEs7Q+9PoclzpqC+tzPWD8gHV
gml7Yk0Aw63c9KV8lAGWb+D4pUi0oV8z+MFy27kvZc9afnly3+0kvxfEdMoqW2Af
fvSlDshP3/bDJ17zlyJ1lUXj2qZihLKAGFlBXqc9wT3sLrws/B7eT8FF5SW78IA3
jpx1a3WmO1THl6NhR2s4Z1R3HyIL0nXjiNQMe/dCP02lQeLcDRhkZgzwEKeFXDUh
Y1AMGNb3ldt6O4/Lc2cfC+hHZATMxjdVx6kXypRm8VsmOhdRuMtAHRx1qxHiryBY
O44GpMQrxx6sWLlPRWnWCyFXkvN0frlCNe3BF9lpi27FC+AKSRmU3fRpZrbKw9Br
Ff3jXRwJADHYHt+KVeFtNTdPH/ni+K8oXt1e1IS4OunGI+fI8fssFnpbF4V+bIHo
Gao+Kvm4IXTSglqpS4NC0XDDazZKdJMDQJsluy+k7ps43V4M0El8SdUi8wayEmOP
TQ6SwXp+ia8a3XsFG4P2Rdnr/7Jqa99nGM/YYUQhYxRkSdYvNsj5gvZOVLWtXHGw
ck0wTz6QbfFLWFqDo5yEx18u/UrtWxRxUqcWPr54iz69W2LRXrjhJufV5MWpCe+5
uDP4kfOCAxcjWbPMVjihbW4OM2WyDwqWosdIjq0eiehqD0CVy1KYNwI7OKnZkzso
2ju7XM9TVll7l2J8S/EIxsBdNN79RoodGm/+wqa8JQJTDKa7qMSXM/5L01iBmLms
itqIqV9qgAZ1gIkEOB4ErvFE/qfO0q6fMXtqBZfGR1TVWwt7gGQZwgeW+/C8UAW7
2F5+N4tJKDka2ejSTO0z9AQ8P+ds1RNzjFB1v0tMYNlCKRgxzzJ0oWiy9ufJGZb/
Darzoq/FZxEwAIrW0hlrK3ayNisCFSIYnrjBgq7Asgax0nEKNVgAad27VhTOeFY6
8yVcEBHaWodIlZr1ze5D2qP/xKx/Ghs46hnF7+Hm2pVSeepapzznMGWwwtU3sqDH
wm3JAO351BquBZCMGUIKe0n8FpZa2ffHLZPXcYaDEpup3FJBC8xzProYS3FMOuSz
trbWiblE5TG9sjViFeNNR2Y4+0e2lKkD/s3zRqWrTGVieWWSZ0OqU6CKWoe78T7J
mayTSQZFUK/oOkUwZpLzAP7KJnYTqImwvv6dTyqNDLaJi2W65URN+8qa3tUy9t0A
ufTHJWJrXaYeqlgD36h5X9BmRFol3QXsrWZWiMF0TEK+UZHX7n9N2O0VID+E9ywT
PIqHcOAFXKwWh4LOinXDZNJbvU6mZFwDBGxVEgCCKrDWgXpH2/DtAqgWcddu6yQe
2GGw3EvlAV6anLX3ErEx+o+9K2O6D/jLCygyvj3RzzA4/8G0diUxZkUk7AABiTIG
N11plyoBrC08e0s+rOB0fC4iB60V4V1K728Y8ioYVIeYvQLXOvFqoYYBceoBw7bx
yZ7BFjgDUz+9u8TFXdPP2VserpRHvpJv2/Sd36R06WHB3SOJNueeHIO5K0X8nMGS
7IS/yAanPuJBaLUSs2X5yyp/MnnXbJNvTn+U89SLAuc2wpFE4WuBPI7YgVZ93n2m
//jicdVtX/1cIDvRs4UJFuIp0Q4N9UT3AL88YDssDqwS6fXYALr7s6IcGOjgEwrR
Fkzd8ikAUej0NtrtRUNY40mCQwqyXHGHdbusU4svZU/TE2CPhYlsh6EzirRKzPx5
ezS0i5gqOvt3kGwoMed9xQdRqHaF3txJ0B7KiAm8hP4VWxob0fUt+MzsaySsADyc
n4JjvMWwFY6zxGixZmKVQ776nLJGMPZce1Hz9eF1wqcbZcL2ATzDSMr7hJzWMMIR
FGJMwkw4be078lq/8n4IxFfjpG5XPgXJscxvutrtzoexYeG6b3Cl1QiQJ8reMDfF
WfLYMRJe9O74EGGCbhuvcGLIPsKD8e688kzJesMyP4umuVJ3xwKV91uoEZxuP4gm
ReuhWllFnbY3TBUz0VvZg6q0a2rm8Dd2is7jW+CuyUUIgfY1zNGZGS1DWOOhj6MV
EZ4kNRAGb16ECvx3PYPn0Eg5T3SCJ0BuCsa0MD7neUlD9BH3doUxpNYIPAIO6jUd
A3UEbl2R+rDQnrp8IfYIEOFhyRFkZ4ohTJUrLMRdQ42wUxWkaaxgrn3A7mHvxE92
2orNlXCQP0pdFhjYL+kqu1DDn0DDn6QwO1LaSm2dXEPKNNDw7zdHnjDus8dYOvrq
Iqi6wPr79pK2SfhziA0xjrAphAewMQ02PUJfAHeZhhrd5dYy5NDludmeobH0kp0Q
7694XcURB5ETcuLBiJYDXV8rFL2zxKE8szXW48QRHfABc5bWWWKRtdJLGUVNG6kd
gae8KCHp6Gq2j7YRclkPMJJRgsO9av0IlqH7X5+Op55fiODIZJHzerT077d46H8z
dBFJmixDrFHyOd3ZgN2OiZfHv5fLeb71pZNBsh7hPieMENFEihHeFtlCZVLsdeQS
9Glg5kB1EPJxVyWz9YXYBKomob2wWAZ2gKD1HrZJB1Ew1V27yQCVoqMuK21aBNJB
gQj6sbBe9nk5CIjQSMKbDaqCbD6hvVHRa+KExve4eOTs2i8Dpeg/NQk0qNy+FWZC
7Ms4cjWehpT1DJLfqqVRM/La2+hF/keUvqe72MN0LqwPvBOMPxPoY/CnPflbVNuz
PKpyN0l38sjiWC4KwXZuSPgDfeHcj8z4aVJDgF925y2545VB5Rhl1L9de+IK88MO
yiDm3up42SiSv7tPEbDNaX0tch/fxzevwGeA7ZsjRmYoOiHGG6wW5Vf2Xuj/DZXj
Fr8l5xMJKREYNJvvRpLNdPVWVogkT2H7M5WO0w5xPDdjL7e99LoHvN2bJrHNap4C
bLiRZvbtvEZsoIFyOhDIE3SrJG97amfcBuGrGRFWNFi5vcnPyGRBnc55j/96NsEd
RNZCuXu7bKT/lUtzC5wZd+FgTFywBaJXw8jNqSXgkd26K9Rf5P4vYgX/+8RpHKgw
TTE8dsojG4FR7aur2D6JGZtawxS+N0OmgN8H7kTm0GqGeglqWDiI/7inuqaxDqjQ
fnyc5BofjrOVghe0aCT+KHgzyO9RlkIQnwnbMcQVQTJiCzPpDKXN5HEeTqiBjMVj
BuUrQxXZfoRZBTP+ZZ0BsxhQnHsLQh3bsbz0n6Q0BQNiJW5Xtbkk3HGdidGjTmXa
ASAjPmUMaFz/1IimRXK3CMD0YYRXX4IR4v3rCBxKndnUjwgEN94qdmwLw2azflx4
ebWob0pCPkqC77Emwo84CszfPiwxeqt14dzRRSGUtLRaKE7h6ADTh1VnO+gG+EOo
NE2Dw3NfXVWwGUiu486s+0oXfWpO7qhveiaGdHl8N8TW9mTOqQzRQBROJuidr6gF
1NcZkpXXXSU0rAOEy8jG6W2W/IduG2b3wZu8y+KYHsUjZm+71xQoLTlpCrvcg0/o
cx/NcAEZhXRnymIgCq9SZtbFkCwqhJT2HHhpXD/9IMIBwE20szESRdn7hiK6iBlm
cVMjkSoMmSOvel38vrFe8TEGfFwgHADkQaOpcO2evyW4dSZWyh//IT/6RcAqE0l1
5dmO5e9cCaCkZs4nGbt2GNa++nc2TxoaVpUbxUqxs4iKyrieXyJYClWEsAfpA3Ph
RqWnxzqTA9Qw0FWsCzVfJQFWQ/iHhYyTFP0J1CdZZlxfKw2YQBwt/nouoxo17QoB
wh31cgWREz789xe+e/6f5hPIi3gmoSL4YEWJjDEMDO/D68KBCvyyrCRzxjeQgkv/
LpVsnwe51XvtgUnwlCsOImJhHa06sGr3+S1hwL/tRIsimsFCEJV9eSj6nSmmS6Jk
9nZ8vDi6L/r522nsi0e3IGJ5qQLDpkhsG0QDt4d7Xsn7i37ifzRh2sjQyR/qg0dJ
c9TDNCdR+aCUo7w6SKykE5POHA82KCrzEjW/4sxBydz+HyWCbu/yoj/J17lRi5vc
uK/GWkLSzKDNJeN5ntVDnby4bTvMCJtnPc0rcRTcaYaSUsgoIifgNC/jiq6eWV0E
O7WuSMv3d+8GEilzVvMKfRGmtt32MCRsE4AX3vhgs/4/IJ5kx/eTlbKKjmJ5I247
3Wrsu0sYuDd8IxKksbEciHUJ3maeKnBGGtc7QUKFbfFqrFOTadgInAsu/RWrkcVa
BKnv/sdnEfydweQIA6OEnbSF9s1EwyZCOzP6biGt5sW8qSuCfO/h3BF2Bs45Virb
nNtRBY4xywy3gI48W7rBEo2UzscTzds24AE/TrQNF3JL67jo7KtRREcmQtj/aPZA
8XqghCAMWxizeScr5CheYlrnw97PEJT5WaCU/AmkoMSDX2CCd5y83GhUAxkug3oe
kqFu5Wzhdghodi0cCxRqmB26PByoxpxRIwlmri+7bZMHgbMWFNYLriDAF+SH9PR5
vnyXVc/tel6BveP653B8QCx2YbeVz3Tx3OJyRvWgeecSIiEDu6GQs4PznkX3LJpY
k/JYSpk/DnSbsaBA7JTQOrXrpN36xRiQDNHEywEBhk8z5dToBFvsIVS+1Y7ra8mY
3ERnwDD628yvy5yieokx3qi7mCUwQ0SkzGEdTFWKWXIcmLy1o9DODubnoPDPJO9F
5T/6MTw9m1jVGM9vrP56ew4m0Z7mNaS3wbtz30jZdSwDCs3xGYMaj1VWzssLpXK3
04ptdkw0KULmBAMcNL4DrSrs389ZuAIvafRCH82p5APrG7Mvczp+QFk6ByKUrJdy
dVEsWiwiqb50ooYqDz2tq4p1sTBniPie+7s9tlIaG8nj7lFK8lk68Of6WoAcAWXW
6uWP/HQqp7YNEyXcQ5WS8Q+c1n0sjBp5OXPfiDQbebfbP4XNsPboOvz+WUk+a5xh
TxuL70gepyiIUWvpy+DL8Yea+DtLa8UrkctU1aLnCBm7HylXQgprLtgYqjpJXk/k
QHQzPkM+D9IuA+3J8idGvLM6Anrv8tHuBrgA3aqvjPN8zJOiLbLSbIZ+20Nj6KIC
Gh8+PFUQqdjT7Y70tMWy/pGUUoc6MKXOC56SWSfTHMP6Cf5LTWrFbEEEzx0nA1R2
dLQ4JB7dPVT17xBD4nttxMrMsBmcMaYQal2xChtKuriK54DwxKgMu9vRWpojCEHw
DOniR8jbQZv6h730BERjHx2v49FZ5F9q2yyy8tYKUO/qPf5TZtx8gvK1E4SDmmED
/IH12vkZKM5Dpn4kzGP5SjcKHaghWpiftUquBrG+GTxGsWg+LXJXxTn2wq2f7Zuc
i1lH9Q9RPQ0XSmZDwRFCfkZcss2A8wNkLK9dLUcmgmUMl8PJl+zfvOcHjpdOO6cN
Yd/rGnOYsnOeP4FNwEQMd9f2iZ7mtsG6AqyRmrYpM4choqbPXHajX8tCnn8KsDDM
VXjsAHF6hbufr/I3KHUVv3ww1ZoAxeAWDB9BHQK2osBGptUyQwc9LwDp225+LkwJ
LabjzNPdDST/uoS5IM+EJsoDeMsMcpVU8v1oiWep8EWZCP+3Nd4F3T5tTjV1nyTO
olPYLMlEx4ixXO2+7K9TxaBlQHAUiHe1ElZSJM6L9KtfswFnxiOSGtRveQs+670Z
gb8D2sTu1rawcZn01erWnlZyb3KyxExcC5btUjy7cdTjQTQpkCSOz1qg/XHy8ltk
cph9MWwwwxGROuqVK+7OGxRHNDlY+9FcUZsQ+Xrrcl6dxQrYYwXIr9WGpS+yqVs2
By8DquCPLe+fNUWn9iJaV1iZtTwCcuKpxh7AJ5st1xbJSmDDtmGFgL4oUM/tDxYz
Dvrgk+UIB6nd7H9D0+iJjIaPbrVb8jyuavL1bwl1u66FBiVMVrQtLoH72bp+B0oG
t6y9X3ysXo7fV5sUxw0b7VbuapKNi3HnVuND1N+w1XHIHYnoEOuRjrDchlMXih7C
0ArklyiR17gv3S0A7DrQH3xRZtBdQNnHg1LHSCcFChvJQ3c+HN5oSGlLIgToq9iF
WujRihNmNDUlySvxyx+WCnPyD347s7e5biLyEBvCblNuOsANOqYLWG5DU0bucbeZ
O0NcpcIT95Rj7MnIXafk26t+hTjT4CbZJpUCU7rpQ/LRJiE3S7rKGszSNYqag9GX
UXq74+P6latbWpiMZmfQVeaiYwKCMEzpjvss/iLKw9V9i/xgeSYBlEVTMfiEEB4d
Bg9zpSCbk+HQY2PNJj+BKNjTo0gSxW7E/FRM9PDwqwEzf34AtKr4cp0Go2bQ2VOo
PAb8xINgsa775EHS7hkkrxbcvbbhCF9yuYETP53Od5BsfX1PAFIUSrDY2UO53sfg
wLUaTVnpRMwuBz2kNBH8Hgl/jkec3U1sYgW1S2x03VhyyxpMqt5PejHUpAFx5W3h
lcpIcRrh3i1LqCXRlO77Smv96EaqPUlGFtzGBaz6b1CnwuRxGiDX3U2xibs6hrG/
047gg6hWjmQu1j+gJsRWFzaGR+b9f1lTkOHNnfihFt4oDgNCaM8leJvYr16jkjcW
pshcaSInmxmTRJdl4CBb/MOC0jW968XFKZaHajSPKrlIfyZT6lUuukqVuGVXzCcD
pk+CoWrA8epq5CBsMYyZrHwiifCZ4sdo8KQAa1sE92yR5uznyg51Sabty+kXI9wP
/3gxylftYCynNaf4ESFlQfwi1k5PKg8jSLSwShRNsfTRoiA9jYR+9/V24IoaZQ9p
HGrtBNFHjL5dyO0JV9b3/M1szoN12/nGki0yNjXIf9KyZUJ1CsUdiQd3LH6SY3xa
L/W8nAzlvgRerzXXI9YFGm9i49QT8O6083I3InG/ClRuJfH64D73EB+jZHR3rZtK
nhnvRgsCty9yIF41hXZLRzrxjkQKCKknef8OZrk5lkZlVdpROYpS5pX8DWgFvRIj
tw5j+Dp7GNO29FDLlfeRrFEYewzwnzRlETc76sUe1IMmdymGPzEuPq8F5OnZJKkk
KCAeLbfOAeP0XuQ7hbieMWLlLzccR7tG0EquNkVRozSV6ib+h+J+rq0h6czPI8N8
fjJKL8ksp4uzv9VL3pUSFZOn68lQh9InZrqEbIJ6GzDcPcp3qI2dri60yfjs8A4T
eIgOAyIum9c7QdIri+OXIT9Bdvb5tfWwznHyiTSovaL3XPns+q7058ArHhs5rCF/
igcdq0+9pPItvztBFzejw501vGmZJtohe9X/ndkMw8xR6uoYjO0FnID2uW+k4F+H
PxOmWmzt7Vu3e1pyHGwwLhdoU6yPfjwHfqLHONj5dpvLjs0e0TKiardn4OKFkAr5
m6tVdzLiOQnZXAlNn8BonaQieTB6IEqGoqNY8UdgXtiChZeZDX4dBWbfry7AMN05
pX3ryu/XAesNEwTDgJB/DCvd1rXmIis/NM9hSfxwyd5RkMD4otMAVNyRv3qzEq5k
sh4PvslyUu9hvS5ZPJlR4pz9uYBDohzReQSZ3nDqtIzIaGGj2PNJnaZ4mWzh6VeC
s0HR/XSEpWWAI4oS1CIMqkPF75BFYo5/ZEsviHSdbrTxdlFt1S3R4cWjCjJmw0pq
vshjUjsJRAEfI9HpRB35SxFmf2EsbJLWdEB9AdSIfFOtSvMWDU6mW7bxbLFgbkQ2
Of0h5RJharJvTMbQzv7rLxvGTMkGYjTmTrS+2N72H8WpSsy0QYiXrgTleqoloKnc
1TQKHIbkQhqxCZyxQpoMZhFSmYHd5uopZNovhsQ8xurMqjgRFGoA2wjS6+pSHKGb
mW5QpOwPj+h2B5qpuGVo7bQM2OnoqkBHSK8+lOoOKP2hP9C7edvh7FwyWZtAeIuR
/CtoiOYO4MjY5E7dNyJq3IuRBDzx7kOL4ch2B56hfLlyCmmcGt6L5V+PjvYwgx19
aujoLjnBlD5Spofp4KJungAmtpsalZEKbW8V6VsPec8a0eGsCMhQ9L0+yQEFgid6
4lxXJys3j2lykknq25VVXC60YHvH3bcG3ppnkZ5uLYnai9ZKqh3JN5yH/97HGcTb
m/3J6PBg2wjMbnMjtv1XAf3WURcPz3ql+j5+4gFRfThSDGr4GlwAmROQq9y1nxPE
PgUFNLrIOW2UO0t/jcv+dRGmCBJuVkBemUn8CFziraqzqA2vaCOK7+gHXfHwKkfO
KwsWRiNmIFN+7wEtyh5QpXJ0iQoUBuRmonjV7AIpgrjnHefIbvjHgyXuC0z3JZvW
H6AyRE8jBBNnnAcnbqvDJeDHnY1n9oArW7L0Dxum3qrkYoDW8MlqVjKju1VB8Ai3
u7EZbGQyOrPAmpqQFe3ZW1YFoP5u+aszlPjHdrfDnQjtvbZSg8WQG0I0UFL3TURX
gr+kyn0W4iTSUC0mQutpT7dsObUSxH8vH3npFplW/s91bH8dYITHum/1pEJljcze
QgwnXpmWqJXBOc3+BhJGVh1AuC47aRktE49TOqPkk2NNUDQQ13+6vAt/8eRHHXPF
uHQq9jpBWH77rHf9W9dyXCc4UE/8CyRclpGWl+NGewOt9A3IX38UogHslG1YJlxG
Q5lTYjQWZjrK/UUnDU/bfxMbF2nKB2dpahemthThYyLH+sOmVHpKvCGt7Ck1IUbS
zqwJblwrsvXu5U5bid6FOmgp89mq1gB5cC9DRIdC5YKs1YFcerB7YFeDXjJvTejT
0YLhWcCIwzj8V7K1iIRsIBnSlZKaTG4DY/OCSW9oFTrD8BcsXbQEAOCcao1IHQcC
F1J1RXtvoMvqEH8XgiXBOzJeSGWul4YcLgYS6KQu9kBi/10gvWLTixgPjdR2ZAw9
3ln9gPlPNzMqaaNqCK4FMWMDNduCP+i17jlxrVF5r89h22V4dA5WgUOgVLUsdSBt
tFD0pamqpnPRiPAk7LolMtbCaLPNfz+Pb0FTmUzEmShyifmlOxkOBYadK52N7jfZ
TsGHVcoEj0xNUHzqCFUehqCVJv8gJs/00vaEBxwbgeUr0mhnM7yHribpGvkLBRja
DMOomaUYG21TvgRCVQOtnMG/Opr18z4x0SchGgKkIZNOIMV7oxOJ6hsGxQs7y6BC
LG+e3hg+ldhylwSyAPT6YQ2bF/PQx8lXuCC9hxD/A46P+Vs9Roq9j3dlmFfUMbI8
9TUFa6pNCt3QMJpn5oPILnMbZjd6VpBeW0f+Eeu81vRF/Z1XGqgy2y1nzTJFfcGL
rL6Lq5AeDOYfBcFQA0yVvToxrHUSU+9qqM3S599QGi+pUNnsr8wZy3tdfmILppqt
D25LmxahjsXEZFHRwYfiyyphirk9K2h8qlPf4S+UJDh49cizA1bkh+FtGsNEZOc5
9H0b7+EqgfZKKqSanIDhr8lSZSCuQu47mSG0cxaptX9d9hlHQM0E1TiMQK3tk9nz
QHbTIazfX6hmPywj+aPfLb6Zfp5XcCq6PgDxCahdYzmZsGI8X98E7MDH9KYWUpW4
TJ7kk7LtJDIzsZ4bNlRuSbvozUh82Oo0LvHe/vDs0qNF0gQm2M/Q01F8Yi4ndGRs
g3Aazf4Nhqh+/PezorthMgtZwWIgP1xR4rWbgYYAPOhnc69XzmEqs1g3HBG3mnAJ
K7+SpulnqXf4mh+LcUGuDGNoAF2x0CWvDGidiBpzHA3z2iyn3k1Gmrhn9e5a2Kts
wegXsyR7Z4lOBF8wnWkR5fIr+kcaCsa8VpWVwBTz7ZP1f/n3WntxY0vP7p+5+Isr
bcfJ2sf6S7AZrwC9AGn7FUwOB6bMnOzE/0Un/AhbP6Jxj0NBmirVSnGOA0wfjEDP
0CtlKBGJx1lp/Z8y16lKu2E6PHY6WLifk9V+S6YDvk+P8cHLcmvnjp7E68L3AiSh
8RTi6vpLtezze4xEvjJkSw7xSrhDDjDTrFiekZpv6zHfHWqpgto/le32v1qxqNqX
16jglw63Yj4LBsHn1BTsZ6ZrpAQBApz1BokbADTseIZe3WECIoZoUN9zLp1+9nOy
ieWzdq+Imf3+ACnz2VjsiMPABlz9yNEtOAVQ0f3Wi/3tfRzXwfxtInX1UpDoQO2M
b3S8fdMkLC5m73B40rriwPSjEDumL+4BLGtJnUyrG4yZ+lOCzKWDVR1izAVTWU9E
s/6b6yAzQyN0OJMiKNGOlsSgV+FHGLOl+Fpm8dNbKaP3HDd34gujvujTrMZo7PFb
EmJZ0LYoxDmItDjtzcOh2q1/EIv8AoSNA0B+Kmsgo4eaBTjnCwATOd0ZfdC2OcGt
dq7ZiOVtDpD7rHlI9fytywA+VJFZxnJStGGn9C7eyombiXPUdWysa0C5BSnKIR7l
hf6rKc7W5JyvRzVPHenQcL7rm7+gkK2cKdvubsYQeQCcbGxle8NmQfLnJuBOxlPA
V3kZnHWNvUt50AQLd2ymWk8/ZsPL5z+L7w4Z9cTmvHtOwuzqO9wuWTNBBLWlBBZm
+iFgdGLgBIkcTTtn6spiL5jj7g/2JzXqAohTVyaMMBJ/1VX3H/oQEOaZthe8LaRR
7xdBKxNWTb1YHXOLGHFC/K1xM+bFBPRiorDnJ9rjQQInPWZ4aY7NSPMa6t7BI+eg
y/E1emAfz1ohyaryn7utrpKaoLa3vRwC/raxRoUetCgqL8tftOjJZQnb6zjV8uhN
wwznFQm+koWMXK6v27yrEaB0wuflr+XLXQjdQo1K3RYO+dF1o+oUhZuL6mGAP6hE
E7VCnKTbHnVf3ssSg9RMbEEyNF5qWGToiaMTuiJir4U1H/FeIUq3x7HvmvoE/MPR
BtYSol5DCn8yFDbbvfbq6yQtvecVaarKceruKWlkmSS+++8mbRvHJ1G3gcBR5uxP
Xy7MKcHR0ES2gIEFvmx+2tn0psy+SFqZmFHKCioGm+etJOG3IaKCyM05Dl9YExjl
qa8YKx6mALCQu5grGFxw1yy71Uh3UVMISF7VJeQKEgX1V7+ZT+xjD3mKV3u+AgiD
5BfDIe7tfevX+QvJIYyURqaj0Ux+zdTy128HwuC3FAHhLipcjzHwFbdd/ImzesU3
gwwiYCCsPGXAXMk+ikCEX2cGIpJfNDTlVNu5DgLADPwYiqeheBSbhXh7pX+QhNWO
1TArEhBQ4VpQ89fWUeq65/FpIO3F1YWT4RIaVXx3phhF9sVGRumDiBInhqSr9sPB
vJML4qXPG6hzXSgO6BWRmCr1mZgZwUYciAWsUcP+TOBdWhxPWw3sfKHMbxO5VEZ0
RbN+qPbSt0QnuL1M6z3AmZTEpI8eKufchMjTJUORm0xNvWTB7hIUXgPyHL3IKR0q
5Np9wvJS9jMekMOtJDh1zFdjpbyxfOa8xoAkggjOe7lqkKl/3SYJsgBUNU7B2Q8m
SZg0Xj92SQ4svBN1ttfzLPmYUWgInrEYdgyN9bSVHITkl0PKWrfqpC0Ghi1vz7Br
ETbWv7U0EEipPMIagxRKTF+Al2cuMkThKpbwZMtn9Cto4mzlPs62kxHLV0olKNcu
kNgzazmAUQwBBg6FV6rjZcKVx0GWMBZirgZdzO51kVuFcqbkAdaIPOul5SmXfMVx
cSVW9hE1aaPdnh01niCen+NdRfh0hB5VVS4UBcVS94GeTAT86hZ8+Lzs4L8KRGyw
/mpBy9ISCnHSqeDXYqppDpEB2Sp3bvuu4QYh/mKGcnmPWXnnbtIHn3EnTHKO9dEA
KzfXZmsQmMw9hp2sGUA1PYdRQrinSeH1EfRRF6xm1JDmrkgNtLnb2utbwN6Emaec
VquwUX67eCdY2EkGvn6XGtC+dYGXdCKNRdKZczwhLHCDfWgJtOUpVESj4GmV+nOa
jMXbEs7eWsrNrlgVpSChg/A4aYjq/sl4gRsrMEzqHzhMoXezciEppcsa7qy5BkBy
oQ3XiSuHquwf692AbbHG+oGzRu0yS2qlgpnMcV4Vw0c+jhYtIV+YwmcMK5iGc0Lx
KROGl668esZSDj/vgBfmYHcJuE7WSQ+DPLpTH31o0BfRvHyxFU4a/Gtm4NN15mBs
I1Hp6x5WCANSGFWee2OArlELeEy8BmGpHg64FaXWR5oR+Ts96ZT8OKxx7oOedV2L
TVSZCRq0C9PNeyY/GtzEgTaxVncHv2qItWo54M4l0NHuUbMAXjA8qjUrRaf0Y/Pl
AL5YR+8DGpsg5MICASM7axuqZ1nXab2RzQja2axabSVlD94H1mlMRfaw3E2t2+g3
sdBjn5/s5V/tiOLUNVaPQB2izKJNlRVphiLrS7GGgLWydP/I3MIH7A0GFrw5Cm7Q
xkxrP6KnUSGy9TtvoO+1ZEYrJ4fMFqwNcaloZN1z0Lemy9Ix+wPwmpLmho9LsTgB
DPgNMG1jmTPWQH+YMsbsWqwr6vciq55SLAZQK5GnxWk9g8D0ByYvSrSupwDMAw4A
ydpBfmumBAxJP1btIA0BRfBjdix0WKVRga7lf0DOTGHDBvprBO7HHyaJgfitKZED
hn+WaILqZdLbbMpUi1LXn3c7evMVGLCJQsbgLpOoIyeKmlMgCYLket6vgLCM4A0r
iJytrpnX0cckcidYjokEju6Txu98qf1+UBTUvTyA4X/mz3skaSaB+EUGP9zb5/9q
SNVTGqLcO1ASZI2U4B7lGS5NR/YGcOdE152FcwcVfykZnsMT2dlS5m6kOqu1JqHG
tIb6ZcpcqJZHMSneyvYzrNoVxCkD7l1CZQpPpsqOLsF5xzxqUH01jISyDVEp3KMb
r5VB0rYJGkomJ4s92AA/v53gLNUSOYDa5ssjF/uAcvfNJhnLZTMmSD48ZZKskEi5
9tT/ZfoTzrKZtL9H2Yo5oIV8K7SjtNskG+X2vkdpbEyRm0pnd+kyOCPqW8kEf/Ik
M7ShVI/L+1Trl/Ko6QlslVJQiyeEOooQ3Hhg/rc1pFgXeKK/jJNbUDQS/Dj13wGu
Ia9tc0IHz6bQs8Y9+8duekabVzvSrLPgZtvKY/mPVnGcLfq9wY3ios7Szpk1rBAZ
KoekeGXSUXe6094hwZx3Fl7llBi3AP9+iHf4/+TE/doWtSDXSmnhQSxj7zIYJP+2
JswzWFSr0MVpxvzIR5vJWvP7xB/QRqyiV60RmoM+dypQMM/+g7e+y5FtR+DDkrYV
cWrOGW/o9nRWdf4x6IorCUaX/W9NIYgYdoX1pPGTzS09F8QmRqH3L2TGstUFNth1
hWOUQRWw1A4g5huDKALP/CUkHiO0KPOaFMB3TdgWuQkSFkNpvWrCE32jO0z+QZev
Q8jZgX+Y7cz2C669+e8aYCsNubpC5U45d1b7lPmsD1zTKoSewrt589c0D5Gz5C+n
Vo1GLukwLazEiStFrulVOD9A4sC8bD6Cs4YP2QhLKSl6vtC/PendkHADTBHe3Xc2
E7Xl21xON8fwbbWHKEXgRe+QQA5QuzAqUriqyb+AtsTwNBllV7TC+L9WTAeRXw3b
sdLc22WB7BL3n99QrkTiiGWjmd/LVp1y3NOT4dwGEpm1CJm1ELJWpIm+kdAinNoc
5cR6ge77Dh+rSUYtjMO5sl0fjQbzYbRkc6i4krF90ajJZOmm2eaZC5oH98dTqFNc
O5/tOmYcdsSHacR42Rp2ZCi1w+nVu7JF0OBtQzesekxW/HmGlLxSkPiIpbu7Os8y
0WQwa9ddi61gqoz+HWp2v9Dd9jJmoqPCfEvMwbQPFQca9NOcvi9zVXJxw2ftfPm3
B4KMQXuW0XeBbtqyoCMSG+Zodoi2EpZYgMKHhnMg+PrQURTBYapPXpIy9vw2UqA9
NWhdIjN3tJJp+wPFI3cKgx8lQ39KM1TpXeSST1yvjNiWgc837vrIy6pPaigsR9Rm
tKjp+GZZkLUlyX5FB4cr4z5IiodoK0KfaVNVBqQJ1NDWEjYO9zfPjbfP05Ry8z0e
2YFv6AkcvvQq9PtvvTLS4FW+lFmABLVlPYQ893a8fb7bqdggUZsLxoGDtdvPZ4Fp
rRKwn9a7BD/jwjdMk0Ex9zp01TjayO+M+TED9RYK7ICKxY+NTkNgLNkMfQqdTT0i
/r+hsDXDH0sVaj/LLIyRaEQKxBrcmDrk0f2ACXRyqXcipnKcohxACo51k9VGBafg
48VA9y4lcCLFkv94JUTK1Q==
`protect END_PROTECTED
