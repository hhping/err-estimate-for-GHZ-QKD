`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mR3HaYm8bcFH8y7IjHuwxOev3SC9OzTmhj5vT8t4ufQ6Yb8627EInftZ2SPt7LP9
vtHLzhXEIuVFsjPwuW1zrQ/QGuHWdwJRqimyRkZue5r3s/M+HdwQNVWqsuXnkrBn
Bq5hkPD0uNgHIjA/DIw6d256Y28YUsRAYGKAXfeR0Tmcz1WWCcIz2ncs+Ex26iXD
m2L+ESFNK9X6ZChPud6hH4EOfw/QPGrGyHV/6wCO5lQ7cj/yQ3VrcKtCa10FSuLk
sTcNSMJF5yZL/6ciEGjUnshsYZhARs3KB5M+1TRzrotv94PcOHID0XTRzB4p/ckV
oL4iWlCyIKa6hil6UDF0eCFpPHBMRIjUBBmqjiWeBkJGle1Ji5jq83S5fzKU+uOW
LwbaGTC7ejxl2JvHOl0Dz/GR/IwLLf1vTSyYU99mse+CKYisUvek7qptmpnEoop8
ciCEcP0QSddqxAK+c3ORP/cpNO5rt/evBKapKI6QUwNK1yWjzC1Ni5FFwuc839pG
2mcfsdQVvZWJOXmsg5gMSGBd0BbfNZhzG3TFUYQHD+004TQiEPPxbMqSw2YgH8aQ
uhdz7ERY1DoCYZf7MqMIk13uXL/RpcyCRvQq9bxHnYGIzmz1Z6exMdyJp3A4dArj
dh6v09laZ7jznmpJJmVBIrdb4V68tbr3sMYItnNFA3DhWwk4buNzASMzEXNIrkSm
gXe77MU2GXP826Lx1eZofulbt7hQW9mDhlsYsVBY2r4Ib/OUtVHDc8BIMGzyGtc3
MbzG2rA33wEMUsKaeKYfLtqV2HWisMFtPaG8ENlx9c2v4OryChJe7SuXXfAedTJy
9WSotMPCID9jtaay9Ng2lGuExCqGQWedEkYdiaRfK9Br6XUp4Jx3yoeJ/xQ875fL
5uzv6cYmi4mgAa8rbsHzWI1dDX3reqdTox+rFxn7Fy0Mv2hz1G/X+wEX3XxIaxoo
jHQ0hmqUMCgJa7+1gC45iRSDRsRiY8o3/9Rtt4QZbugEogBSpTN/3q1uj3fJ6iBC
VxTa9j5kurOdmOZqcNxSdD7kuwwaLpGNoQo/3LiZycE54zfK2E/4cb63YUffcB5m
LuRXTD0/Ft+ZZvoKWgsb5SJhCABuVBUC8lygWFrq2/02yesC1VAv8cjCnzT50dME
hME9F1c4Qlx2EOasJUiTm8gHbZnj9Ce92NYS5deywqg/K7dLm8tXJCRtMXXrBzZn
9izn1t8QdvCYfFGNinbepkxcLz0Z6K5stGk+SW4YBLpriKgKCkHz7UY+HW8B/tgb
Wu9+IdRiOL3bBx7hiHg2AbNioq0md0/vUVUQpO+wXU677LhXP+hdV+cvhdUB9tDB
vLljEQuCnjydGqVpBbCLIa3BJHP4BHebg+u1rAZHmMuANXavxZWAV/sTIEz/okpq
JBNxFCt7MbyYnHCnbBUK4SDhGLSoi8A339ApeOQlvH4zTV4E4DNh96iY9fnKvnYb
rM+ruDzTREJnwt/ogvupxfIN2D1AGq6vpwo9PUMUBzCkRSr0vvgPAm3mHj99qTd+
/FF6sOvpJOCDacHyexLrRnhoAeQ5xY2PLYLlTpAhG8hwPaw4nwnjuccUpVGjMoFO
R3z2VnNilHjK0MzaI5uImAvNyNMA1m+SFsiWBV3I85UH5TBsBj7uV8aG8PfRibrz
9Fqx+R3Xa71ctpvbLHRDMe+BBY49wmWpwe8Ycjot6YkzlCWtR/Yk7J8FBm39Y369
94LxYIfJcuqshYlIyx6ZN5Wm6O58BYf64wytJqwzYJ5r0mDYWSip2Vdr1IDVSQj1
7WQNY1hqGxuA1e1Mh8Mqy8o3YUjo1eK09jyeHS1gI3e39rlem4tiU9cgwiVkeUTd
F8oy0ELX6071QTeETMGmeE3bAHHDxr/hOTKejWbUYTrVA+3FeTsxQLOogt6HXZqa
uy6TvpfcEA9yQaJWY1owauFjRqeiTfrGONxBP7dSh4QfwroLVVA8UG+KaMXEte2v
AbOEjEIHXzCmHE7AtteAnuYg62TQ+CEvxtUZRawJruNG6y3vKf5Ze6dvrDcg9AIz
C6klnqkwFxv6YQ5eeLj3PQAfaArHe3V4JIFbXRQSwtzoIxqcT+dB4xKz9Z9Lidez
YS5f5tEd5cgYPAoJ0nJW+WGsWdat08R1RgxI6ANDXRM3XWThEFIkwWctox+Lh393
LD49iSAQf85luW9J3/4mySchgZwfJNKOuwgT4qWfpQezKphaENSy5zlfr1TA8mOw
glq5SXVFsCuR5Onh2lKDRufvH1lnWqzJFIszzzhuIQl/K21YSaREuWlVGKCHGcKy
6rRfLTNTUQAUJ+OyBugibajzico//DMd3nbDeKBpo6bT0Ydin0C0RoMLFhi8uj6V
fUs6xHuZIUL87eyPLG7i/HQ7WMn5Ww5BQgfIuPZerlVvVw1InJo12uc/Wr/uLo0r
wW481Dv3Y5f4yeGQxpIf10d4MSzwrISkwwF47Cnf9+vE/OCMbw1IylXvzLxTkv43
LauuqvihOXPhNhU8xVhNMDDsPmRfFWbo2wOihslocc+PurZX8P0dSA8kafQz82Og
Qsv6PtJ5dmoQJB2hUgV3BXg8GxgHf8JCZ7N6E2M4BpC9Nm/KbJ4RQJQBr3c+To8c
jsbyGfvZRZiTjZqDHTjMZu3TodJxTHjRjhnCXLeFPfkyoWLm0JLjF9C2X7MmGGBq
UWX4TIGu2szAO45VcuH85rniub46LSavZ+vWxIarPDP4qVDqzyqHgdSODp1ToBxz
EzmJg1aAI+yM27kToSmj+DYEhcJuxMmk4IK/4MqAfynjEeLSDvYhbqjaOWta7ak8
3z8bksE3u9aTARx2iToB1qMn4Ir9n1W+jHQf2Bx+nNvWc3IcPd8fdcppGRVOfweq
Cyw7YUxP4ei4n9hBO8P+mGqnOaA5VkFA4yQDvDwUvdGsSenByE7Fjeqd2Eyt9Vjg
se+1eyNb2mZDcDJWhq1L5DdKMxJq6NSWnU1eoYWaBeEhN4skR2Mrs2O0mSY7vZi3
A2zGijspWqvO6vQsDBFLnYn/eoaJEQWcrQQ2hSyuPv15iBZl6rCdBTBOM7qEyhKv
R12lt/Oj2Ch0bR+4Teo+LA8SSc4Y7AYRR1ZcDc7vFIRa8VyzZY5GFG8ZZNFFZKPJ
HoVzgWFBzUmfMTrFimRecoWS0AO8iBfTFHY0Ql0rIbva1wke414S8Yj0n4PmMUyE
P3JSM8kksUbfGNa7ec5RstWa0UMcegbgeXumcjdreL8Fum27JkFmCyO46VsYaspv
Wov/LrKOnUXCTOkgZITJFCKYnH5za1BzcbOLeGmRRFOti1l8zsM1EFWPHcD0oOoX
U/jzZi8H2gFMrD69Z9otdQugnD+IFfDPhFi/AgziCquL/qpRqew8uKvUReZmBRLx
6Z2wat7UFuSuTKTN/qUmmOL1104JKjL1akxVfXQQSL84oU3cJPHzpS0x2Ly081ig
2LAc6wUaH4el8H7oLsLq/6C8zF3n9dFHThL2zYa9pDXiAHWv4UsjjhIqVPjkNNX2
MPOsHzljFleWMfnayrU70He/OgIGQ0g2owg2HW8hveiIzM7RskU3+/1IZr+ap3ub
aPpMixZO+bATS89w22S1NsaKW9Lkh1uB2V6eWdXvvvN+t3GqDKD/L9dTWTSJDfCJ
nlMICXVXsIy/7QuaFDFaYVBpbDfD2HclXxcUiPX4goB2Cp4u+FfJD7nN9K/vSLwu
7FUomyyXET1FZGs590t1SxjyvfmkCEklP8Kmo6/oagZcb2EHBRk8dCEvFAz34a8X
3DsNw4OcZFZGdp9TJoejSeqm6iH2ATKh+aVbWNC9ITjheGLi8Va+k5X/xbhGWRLz
uUfbE9CNrcrFteHOeK3W6FmbqT5QLnphkNgvayW8S+IfS90CeDIDnG8Q+1pJGg+G
TxmuQqGno74EXi1Xa3b3/jki/yetv/vgYfAZrAFnJheseuhLwh+wcuybKoQgV3gX
JKTUQmLe6H4maDHfuKNJW0Iu6JBD74LAlZQ7i/aCGFesxuxwm0vAD9hHtfsWbG/L
i+EneYnlnlrWPufbFMgN4lI5Hca/hSHXu2f4s1tLDPQHHF6qqmaDPRYWIktsgbwH
mVNwlXUEv6o8mHfRTvjbjIQD5ZxtgXedju/Byrxs1d0tRhMQtKD7L2pVrtRiSQ4Q
nEtcGmdDNGtRGlKJ/rIqXooOfTmBBguHqHQLqsLNxPqDrgxdLGg6E/VJoPxeSpjO
7OBKmu/SY6qAxtSKsynI8apX/DWIKkjzesxb3kJgUeChVTBthM4laJzAAzHEf3dW
MVGi3Iy3ZOe02xWdrr9J3oAYl0/51dceJLweaLG+5lI/r7L+53faL4TykVC9k5LL
vgtucfJjTF+/iNQKaMuGbata9G8El0/w880eUFHOLfvdNOz10w27lOgaM28rtBzh
Z5IEwmU8wfxm6Tm4QfmsXBYXXDQ0SLszfc7NJ3RFk7MGNJ1SFTRlgWKkvjqm5wuk
/bTFrfUKZUfR8lso+6jLIkwMMohjrcJ96ffQet2N4S/9prQyGZ9o3uUbf/T/MljC
iYXs0ImA8tXP25Bt7MQZbVcY9rRqFneqsb9kAlFho0plylFvOpRxUfpVj1oV1TF0
jIozgihjr7nxEc3uZK5ulxZ+wYOhDQu96p9SAS01b0oXTLxX7D1o6zqFWPNteyCW
ginNJWuww+/PIOWGMxxv68ltH5WMQZxU7kLlVgI0Xqy5ST87SGhwlqf61ucVbxNd
ru3I75QIDnKBBZjZ69EfhKbkItyTDZWIxzUQK/JozX+bKci18wFAn3qWmdvZa2rE
j6+S/ftrrOpjyrnIiuXziUTdNT4w1GNPbwOXSiWJtCtzNfAzt6zckJ5mib95Ea6h
jAkx84HVn4nuPGTn8HqM5Qf6L6dp+Q0EONK8OhKTLexhEMXxOxuSFeJaHMzgZjMY
SZdFp81SorO/DOzQUYzYiUGFaR4YapXFaKYPUFrXwEolrc4KpvlWER3u2BfYLfv1
uFaFNeqyOYHbb5ODCXK/mQ/NczPK9lH8XczGSY/ekszS8K0xVcOhb/030TX4n1a8
4NdMQfvmUYIa7Eb3WJWQGAUpAGQ2/w6kLWyirf1qAxSFxLKoUkYgMhhOoq6jj8bb
ccssAjlBSSRSHfPSF4C/oa0pgjNBKHec5pkN0gXvc3/yYrngmXYOMTUmerQmFtFA
XLl1WT2VQY0IOj8MLbshMKlK+LG2HlUptezjE9OTDKiA8gurUHdH7+IzzjU7+1MQ
rBrmTkWoUzb8Cia22w9i87OmZWhu1kmdWFuaKEAvvd/nCNnEanFcXSxZoDsabuqW
m9g0wGnJFJiZ5z19WObOzzS7mgZ/5QP/vc/Rqep/TDqvS7fyCpRMbpDxwr6UIhY8
o9FX3yHoRRjHCxuMfSSDfa5d4vnNcXfOX86gX3Qa1p9vHnsAx/BU+Oj3TEnAr13D
P4K8qcT1fZN4F5yI6B3E2tyoFvK5sDXuMhGk7OCeeWNdqWUgVdW5friDuajfO5Ju
RZRuAczFFGNrfSbBS6//2++qyEk7l1AwX8AiyVdXrhp60+anQeoXeAhuuRmuSwKO
hafl/N8wVeNW1U7DHYxvmC4jpvYjgLGV2uNYMOKcxZF33ZC8PFVOPAsuLj6ALAFT
h58JxRoHHWMis31wVhmR2WuqBoBoIXKmxS9wM9ctcJ7Um37IGDMt4skXP8gANput
XKpGxxlAhjNH7heOc+uFkkwfBc4ZBZ+rT9SHixyjoRkRIQ+QXZKWEba7UYBcZHoh
Nl45FDmyUpWnyLTkSwrb2VD64lmAozm/6JpePJPrmOBtFwfZnwC7/HoBerIkj++C
eiRdp5G9zkN3imnfyM3fTllwBrFoo//FeN3BRXA/120/qnpRXDSUPKiiSiQk4OQO
ELVizZYHPIQjPrtlh4NFfCfy0rHeBh20kzNieMvI3ySh+RCuFnnuqnJWAUxkmDRN
s7iXecY3A9cQ2KZNQri0GDJwcwAntFhWHMwS4mY1IYuFCFhX658vd3UytgklUjOe
PJMyUHMoAPItuOF6D9vK6lH6d9IjBdnvoxhl8Wjzt9evrl/jiLrAhgBr2VEDRKzj
4i+Js/m4HkzzPBIDZhTaOt4zNxsbzi+RIwsu8zVE/1R66N923FywZP+M6QXhuFxg
gCwY/ycutQwplxD7YhZrBJIV9iiT4HN8cSlV5HKd84CwxAmQZrICyO4rtNlvCjQv
pphrCXoonwlwBYS7cnd4PGSngKz35FU3Y9+tE373PWsoWVCHkUhqxUqIKk/gUEDa
+KS7Tw149dh6zNHLo0z+VtbSHTMHRxJECk8vNH1N+RVo69fPNG+wEUoG0zUnxEfX
8+XmjmqLNnHTLy/ThEyfuUPQBjoQtO3ICvW2S/EaJWHTpvvCveMuICasmjpmSP28
5T81M549F6m8TyiQ4gWFTEsD8Ce+GyJrz9Kuvvn8aN8KcGWbtme8sdym0VCfF9Jz
PJVk1WkUiZp+s6a87jFy9tK2pfZFjEwKaSFNih2cTSqivLJ5LM3oDnM3GdhVY3dl
LbHBxJu3ZeCg1LfnlNKsdDHkusR/0yAcX0OqMlrc6yz6Mo8WAXPttKA+SY7liej4
1HEP4X1CGQH1PF2zlU9igW1trLrrxRHgW0YUiHjmlIgJk50D/fP9XaIu4r94V82d
WRyuoFj2uRuOTSvsKxz2GLjkjaNiAOAfJnonEp9beKTk75D43Z2Sj3hQZygT5piD
b0xv1u2nWKPICk9BMH9KLJhOk4l/8OojdoYKn7vejr7EqqZk3c+WwZWr51bZpfnD
pYUIql7NDWZV1Nf74vuDNFwbsN/bIclCpBuOzXgnf7AUErOl8NZZjg/oInTMGN6U
zkbHVMUeZzMpHnetK+wZEvxBEnSTRDIcN4Fl3mXRhv2WWPXle0mnBkQM2pTy00BU
CUB1mt4Ik9SC7ztwZZhX7hxEIzTiniN/0Fb9zfSrVJiHbGAnvaXvfovnZYTwcwJR
by+P3YbkCdCCqHIbUoqTN5Q8B0eT92thH/2SX9bw4vVyeIibDGP2WB+8CNS5KwAZ
zuPgu6VhWTG9FZtowcrTrRM7fgSjddQR8euq9G9yyTOe3J320SaiD3ZAPn+HQJjC
2S0A0ssgid2ynRWS/apGEgTf29d0yi3yU+sw8Z7b2NZGW1aQ4XNNWoStSesaQtQV
+GyPP/Duy5+k26tQU88VfsuLh4nb5+Fss6mwottEdNs5sKDDO9ab3tQHCpZVUIef
/GNn0QjPxQGBEkjWxKuhAxX2sHLY2Io5rxrGVboBh7KphP7FzG/DIC+1dQIDMhPG
7+QDwLr0MfhCHu37FS6LGopAW3l5omC8VNQ1Qw0F3R4WgOfA0nhVE6orcmT10A4O
lOs1OQNOfscKCGWSbBWRWbtkR209kAQM1sV8MCGnSAeuvf3jZPktmaImil6570oa
UzDbuX7ocNJ8mTHPXs1MIP10DPb23U/JmzLA08+JKE/mXSmu8pEe+1SgTC/QfZC9
mdlKwt8dAVr9wdjwV0SoBQWgR+tJecDT844dcEt9BjQmDsyM2daHZqYudTvHFukx
v5PB3rGZDDADwzU6/8e/mHmqRA0by2o6pi+w4a4IroZilnlqJ3AnytjhW+fyUk28
77F8WAYoXQ85vx+R1E441LbBZ7IxOP6dcaI4d8wczokcSoMTV47u0YXKb9kbDLbV
hiHshsYp9/LhdUv0YRwuN4DfChT37cT3OWnEl7uPhpBBJz7h+BrLZC3fZUjDy3fI
u126SnWWeN7An50xfcyOop1JGnpE9jNyxAb4Urkjeysippb6He3SaVEDwbXj0Zv0
8T8PcSRicXQtqA93ZfwPzHpsCj3ApvSoTkVcUzNKmHIok68n3wlTzadSLALheFcv
Xy+qV3CEeFhHPjOWB3WJxhM93VE/JEJyR7GCQXzca6HqoOFisCQeTY4W5s8LCswf
RgMlYImpUvzfNbvQgXJbUIsAf6VbM54hJvMswBdHk3HWCkYOeF06kxDwkVNUDiQq
cLcjQ8SJe9JY2SoO8YluQGJQukV/EwRz1NXk9qGChWRkX0hkvIxieYETi+fiTehB
8ib4CAGCo4MQcdye9lMWpVSiBoCIJNaZ9bwtLXwV3RU11ipMZT6sVhE+j2znyWvM
nh0KzzqQd2YgbcpgmMFDlPi+G7ZGJKrAQLwFAY21iwjNCDJfFWVk1IGnz0rC8Wqg
gFsPl0hwlcTqFV5fYZxqnCFdg0E5N2J5AqzOM5GSB22aU1KZNS8KOEDPDTok4OIA
J9ENkr5z3Ai4YUUGD4kovSEdvhqJZNWQ22kiAoJLnhPDapHKa8rcU5wpv11nj4HL
QQNbbWDgit/yLo77EdG+4Dt6jynxYmw2063sW77tFoX4NqLNg891EjgM4syoSZDZ
1aw+sK4yhP98jNiXGBVnpSgfcFw48MxFbXJV4En2CWi3pI3BWugHsXZXF8Rm3n70
8pm4p5RHmEgUHFiTMLlpNSRft/zV8cWncBu728+lLXZLiuMfm3tYzPiqIfmsTJha
DCQo8Jqt0E1gmEoIXlVODnHRCbz0VSTq2oNyQ6A0B1RgX3GPCaw19b9fx0peH++a
vlB2bo5BnMDE3VyTFp0dR3LEAWYBAt6la6OmwHnZ8TOsmxpjAJ5avCv+ZTrXBxef
6sW33If4DcwfGWWhlbkPmYHaK5vHbnZIFUGoyhL9dRG4/u/3o7stDW/6QDLt8Ttz
bYiIaBhbZrDDArMzmKOCtVmJWi+skHesHvK27x1QyoODZeewc0d25lcm13GpU0Um
hVjXTFEC9g8PKWKzxPW9OUKa+DTeJi+nxNEpceb13icj0dmRkBrq7HWhusMYkiE6
7bTFxYRcmDqKUh+NKxyGVEkJSui5G8c4gmh7SQDRdXaL6+3jqLKXxZRXC6K5nCbP
JHTz0+aW4G7Or8wRRfuR3nsmtgvrfyzbNrNaES5T2sp/hXI1QTmVFEsiWHJrbi5A
CONzUnpK8233eLwNWFWXxMCV2ZQBseXmaZikSKAjfh00lmr484cLjK3cJgLaDjKx
o5QrS+YZJcmLHnsWRTsvrlhftLFTLeAHDxeOpxO3vLYBc29/ZfbUdkVivC2peKyi
wQaljlJvzQygZkLBJo2MnyDilqXU+W13n2U+hSzPe3uuT4S5G/L74Ib1Ff1qoa60
+MwRho15Ov1YtqHi9QB5eB/hvc/UhwVEjsyinF6fFMPFK0SkfpL6n37BJ8Dlw6vA
wH0gMG4bLDxMb5GJ2Ft3sLatv3hcwiSss6Zj/rlWystxZWy2lvk5ymUC6yKiaQh8
KNqm2oh05xwis69Bguez+gTieOP2xetbR1sh8aiVx1cXST+RhDOzjb9TNgHtHZ6a
SuDPwKR9EkdLBslmayAFOqeQ9NA3o0PmAjWdKfWEM/5LNjzKtR1f/Hz68YNlGCa2
D1AVRdTTucPADpq/tigX5Mw7uRwsErVWy9XO7nJ+0q4XGVPdibJ2kSfZXMONeBv3
PgoaT6kisrmvonos4qrePI5BxX3v9skhZe4ftzYmeB7fY/9rKWCo96DFCnoI1SB8
NtPdbJdPGUSdtcToWZisYPLmLQKAJUDgBdd1Vs+5ry/K2gAQFPwJTpCSLAaTqkWZ
36Wkm34v3zyhtlnQ6dbRJ+5Go4jmGDOfZ3ncq7pEuzwTm3bQvaCim+xtFfmS6E24
qRwUyyKD7vAAatA7ZNtsqmAvpyAYmC4bbcWHhU9YJyS1CAXiQ7L5Vng09D0dZtxz
YuLL/G5qem77xBEyzCmIxsJTrAL50dFvLTuk3zzkPdAWfrEhXmJzsJXMJWdYv2/H
dwkSbr226KQ1vf/U4K/853pBWO0FjIFkss/Mqz+HMFVZAqCyDKPBXFa5hoAODPvI
CNQXXRCfLe60Wll6yMI6Y1CA8DGd+Ue3962KD7+0nNSGOqbz2EdrOg4snhm9A+8s
2qM1EsW19ibd5TCPNsfWTvDqdeQpjjyTOKGxZxnD5+Sj6oSjb2FlijQyh3kBtGeQ
Im881Kf7P67C6shTc8j+i/E0uUMKETYsmpWVibNWOl6iHofsKzhHe+DK3zV7+vMj
cgV6vDuIXSAqjjPhCQz3Sf1CvsX/4NdvARWa4IYynbCGVGH7frbTl6LKVTeqcBk0
bHx2s4P/jUkjIpSY/GimaMvCMuar3PqTJEkVEr3zVQ/nx8pqbIxB6k3gjpOGD9ka
rJJO3ufVIGbGJ+AF6mcoDWRA1Zz9MTeC+9PluZRGvTQM9tv3gnXwWeQhnaI+CNNQ
g0tgtD5hzUKcGwLm3oKPQEZnTb3KNXN5fMxriB7beNGGTJvm4nNbZ/E181R7z04w
Dq4BRK+G2Au1K+ErWkOahcRiLmoz86GkXxCrJCpVYu7OHl+nUTU2Hr9jCSXBl+Ly
QXC5U1uEuZYCiNu5Ib9hRmRUyJUBpKtB/34wdpVVMj/ZprB7wf53qqsAI1kuPkZr
/Mo2j2yEzz3mYIaM9qLZrbPjHikjqfPwJd4hIfzjH2lgB0DcvytkgwKX9QS2O373
3uu0RlVo8uE8BSk8kw5+x+z2J280xF5zzc8upS55wl3TvpJ3U/P+dtgXSgPvDIRf
Zxi90UCyf7SkFHg8ywhbIYN24hMpLH09JzzB9/QoVpeWy3txXv09DWGlPAevsYzx
zp5E04V95oaTEax64J8pkzqe65c1oR2Chzd9Rs1vPeyLAvqxqbEhi0KoVA0udqbZ
eUQNu7sRYpn0yVVtfp4QfAe/VS8OIvlmcRP68MD4ASI++wmyIVJCcINDwUTmsQ/0
XpE9uUfomGATfYD2q69Kr0P6QKYq/m5IpbCgwPLMKWzPehqSOyU1kmAPKxUCPiA7
An0qo/tvFh5HV5bWIKeSPl1tu7r3d+iVT2gyP2Rhcqonv6vsJJR620Ge0Q4dX3Lj
rXbGs3/5OosbWVfqCr5ZrPnM7gedvDOLQnLzDhPQiP3F6t5WOFWV7vhSTyVTOOLC
Z+iHB2BHzun6i6yz3WJo6IK58MObrdPIYbcw2iThkKk5v45tzKjXFZ9KRuT6/qrf
xMvpLdZ3sFEenmmU1NC4+cyEjvSUotItYodZz1xNoRy7KcL3q5RWoULBS3L9L16d
eBRD7OrwbbOxCwK/FBP44T/tzUP3X7r9p4wlyTrfduYaX4V/0rGP0Eo0JfpflPJE
nuaRJEa1E2eQybWVpTSWxWqcztzKUpRRZtiZL2jHhEiMwnz61qocNiii+l8Z3BdP
sDrVQI/N4IZziG5YifqtosKj8nbVRjHjj1nY5dulx/ML6ONC5b74+64E5x38/H/4
ehbXhEndZ2c/pt/+CieYVhdfLj+2qsxeERqTGqGvcyP9PyelcXtg5l0c4qzp5tWa
evhMIrsxsd4izCSMpAyg2UIT+aSXOB8O8zSZZ4k5HOelSEohAgz9OkblalrOwstH
kuPaSkgbn+FjwGuJN14zGi0OrdQCwrDnTotIvKNe1gOdOhH2U/vSj/8k3QDglYxX
ZJWeZ5TBgMIYO7kt6hwrjyM4T2OJ4Qolz2Gc5UUWfCJ4+3qtPmrZGapoDn7aBlSF
wOAdI863CQrnue6tO30JX840FzXiNr8NMk+QUUG5+uY2ATYhcT4QVqHIp/ZJboYJ
mChQmOdfib31LgshcrvUMPOkbluTnkMEQjoaGUgBBDapyj3dZ8Gb37zlQvv6LwGB
D2R9prDatTrqUQ3Fs2nCOrbleHd2E7k8a6YQ4opofdtRnTtPc/UxSa1/a6+RuTyj
r/MWD0cF9nCVOr/gxMFfPEp89EuONE7e3LrMJkd/AkCGC8zT73asUUEdBRXZDN4f
NXfXf4/AyFWjLt7+LqrWFhhdG21tvQtSt4XmhO8/RrKF5Cxhg5lnOcWxhTuT4xSL
c27jNFDXzIGjIS3XXyQFPyQ4bDdlQ5Ureo4BmP7fAaMYc3fdSsbo4nQB/4FDWdD3
J3TnPwNmEDhU6p/OTF9ncMTFSWhuVzrjbSdqrajqkYZ4HlHTvyvph0fjUuZQdtH+
S5sphJaRgOevtMX2L/+2O0JLHduMTlrhZciNeBbnPZ5qRO240H1NMGyf4CFIig1k
ugL8UP5uoOGN+AMRYlwpWTNrcvWXH3xSohPoRwu5C+UuUzPpvuVzBDyz5poOmWUG
Mij161gCcFyg9IdoGXwrDbbBpRAdhqDji+PUYgh7PSGZo6vqLmdWRrFn3VkQTF2i
dJpG/0GK00XyepJW04cQ82WKOMQ7f7GhXO5Pdg1I9jpwB5PKJwz++OWrNBMYZJmg
RdypwL1Ds7/azeN1WW/9k/JsmXiQ7nV1n3syjpjb3N4dy2UPewQQCKUlZvNi5unQ
daKmRKPJMgZbDGr6PyaqUpxmWUbIyipmwnnq8sBH4mYVKCFpDCfXrQgOnNaqj/Pa
t9/aNqZKCwF6U/0dxtXw0tDFHCD1vrcnzky9Igj/okiCDzxJYQI8oUXSOjeZ+MPi
PvisKd3FfBaUzNzPUatensFlMF+nxlCiiZ2XGhswvKc8DrFq8rG+y0B+4TNIHSUM
37ECdD/NgH684j1C2QxYKh49ahAk7BkLCvXcrDwa3X0VYayRNz8ivzV0JqwmLwil
SGWoY0TS15RtffNXc5U+jNbhc/YsncE8vZBHNi0+PpGRFju0Tjnzoo3o8qdydZxM
mm7WCs+xhipLO7FQe6Lop6JeQZg+sMLJRHRNvsHWexX58tRKJZFyPJW3HuX8rdKV
O4cDJqhPRpWxY2LHmWh2AwxZlP3uH7DBwLiyxpIybYahxvhl1C+XFj75ehZvgPuc
tAS4Yo95WjytnedQkXxwX9HNzngNdur3DTZo3Xm/j5i1+dTwDod6VQNWFYedLFit
FNSVAJdATfPaZLqDI83c144NsE/t8tx3niM4lPudaXHrD/OIOzMTGKVkZzwFVRyM
6C9TlD3pdl2y9SFBwS1IpJ4wzsrn117fPh5LEWMX3XNWLEuInR8MzXdQaCfo4I3X
ZVAz7VYkqmhqrd6wPKM/c52itDkSuAkv8laWcYacb19JfvQbSzZpBhV/2jkyagrJ
ChLNjG4Q4Js0gBSmk7m+VHccV+Pvrwrqia6BchXhPYZUp2/5rMW0W7X2o0rvN91x
BqjGexUmTD+FE67T1Do/wDHFu/B8jaoWs6HFxvk9oiCLL1eOjrNP4BUHr6v8KmEG
mJIXHrRxPN3RaaAQelOJwbS12mrprKnzTx9G+kuLvtotiyFCwItWIl02WYijnuAq
VJmc+VhEw5qBDKSbxAe49uam/YUgUguky8mBc6zFsTZ6N4kNyUBaTKhCzTKXE36E
O27HorB5BEnwkVpiZI37zHMCLfol1bS5XoRUMy1dEmvHI6wjeajyEWhbqoY/H+vV
a8gtLtgL281Oiu7pvSTOPnS3QcVmXor6efkL6v8W52MVtcm/LDRPz7QdjnTKtwGI
xtql4YTlP2ebeDcFP/fIskvF9KgjBRxU3SB8SROsoQ9adMLt8V2251VQQGUOLzZI
VZDuIHj+vvFMrKZp7N+BQnBHiB6JQH1GLmpMO+M958Bv2omv+o/TwLawM8SiPsB3
z3zk3CBAaxY5FJlGmInJM2iJrEPZWoNI6ebPG0eGDXdW7cFHf5aUsA+yIon6NoRw
ytJmBh6LMFEokIOwNL+/WJSy0cmiFlEENQD6p7AlkXo3/V8BWfT4g6kNrW7434mi
3o1xL6Nbf1oJBXdHRZKO43Yl9qQMn+AU71lvFkMeS0ZAX8dAlrb0GSs3EdOWdWcn
Rtyy7XI8dRcvAecFcYOGdnSx2JoAyp2/gItSytSu9xm0cshnlhGaNpfKp3efljGT
7Zif2+cTdZ894nDfwurNHD8bkaLMufW1LwBMWa2Eni8sLgqSblxd2SEktL1rlaFa
xKZMlG3tUs1V6oGVPlFCO4IKEoChosL5fOFs8T2nu8XSZmPd+2l3QrTel0O2bG/s
0UInKhKbaA4Q0X0+St/OOBLDvtcTa52Dgd2YOXzPn/9hQGVhHUBBimraiWMOYc85
hgJoZBaKZRjp+UAM73vdk3xIRV7/HGWUT8YbQBXau/68VejAtboQ4dpji6/yUZ3u
m5IS34mkSvcy74/5LFZWSJ6vEaDBg/wcDAcb8r67IgECAs4g9L8SZbGUJKssZAf3
RCqjwCzqzsfAAlpV/prkLwLnmC3f8SLkhxhIkIo/hoxIxR3j/ZPNJsk5Ur5xfQbV
Szg3b/mSjlSdfTfRzfJ3NBU4re7D01CsLqW0oaQYD1JjHm8U+LkY32eVxdgnoB0x
oIsSoSXXVLj2F31vWotOM1u6znfLJr6Dc30VMbxsteJw5k9zLvhkZ5+bDtckLnJm
/nZJ0XSW8SR1VJcN0fIwrgzUgKRwS3KNR4ZAqtQ/FkOg40wfo/Ryz/uu0ef0cqvB
rsUM5aCKk4ZzrHC/G/dsgm1TVbYjm3MmAa98yjT7wuWM1CZiI32OWmT0FYxiUYY3
btUHM9YWTX8KIqUohCDYwsxqqpMXk9hen5ELLC1LDvPs3WsxiRz9qnE1fMSdfXPg
YieEATgAnApSPIuQHJRfhsAfIv//bLyX3SeJUz3fRJblPNL23N0Ektr+n+PeVNpG
ZCFd/1ez+UBzlEYy0dKBwzHJj5MZQ7s+JOzlr9YccFVIBYtMNpb/lwzXfATwNZ1K
m8FTeTvnZHcg3H+acFM3bEG2jkeayJF0lWgxK69SWobyUw/SCrEwJDNT2/flGqdP
NRDb76IY8+ov6IKwGLdAG/FQ1NVd+kmc3wuVNcCS2K0eYHqo0PrjMspbfISTsswv
GFy86Q+xGMkjSYGkdB7QlBM3Sp/n6TsNDsLwn1mf7kz/1hj+XB3az3gxIEPDiqtW
XBmihCDSdBULCBJtWxyudJsIniMUOD5DHXjbcDl/6i+gJSylRScgxp10REg65Bp9
XnPKnRhmRov7/dnkIolvFLXso/ZaC3s6QzbU0PFjBCHVjwhZF43bhBlzJmkNfApD
WxO0vFzQyK02SFAUczqCOX56JIaBtqukFBx7yfCzh8rxafwo0XyEWniUHxzBM0Gk
+u/+rNl7rMxZBAKXmj2Kf4qJc1A+JONHy5QJ5r7mceqZIosN0pM/u+rfCEQDRN7Y
qbOVhM9h6fcc2wL8BKK7J6H9OpD7deMHdSV8MfeYyI6rkDjw2qykAkHRpJA5oplS
KrUvBSLfaMBzcurxV9ti5J0fCeZoh7GvXydcd2UQqegaiftqyat5Hht9ZPL7K+AB
+qIqM1F3VlWElKWw9EVgSc6JeGa243g1vGJ/NCtjx3R0y4h9Ql57vSptVxrentZQ
rUwiWIJqdYV9U0vuo+kxe7tSm46HN82/ig0qJN+mJm2KcuJqyeW0BcxHErc0D42U
WN3O2A7ohZuN+vypk9AbvkMAzEWKD0Akce1L3ZWSoL9bnKAMVfyXXQi090H2Bv3G
0eUf2rrT0J7v/DY+QxJq1jN/4V/n4VcEuCq240Ft0n6RGlP4B1w+bN665db0wBPc
b0fkKqHyonHZ4UoIMy+uniA0Ft1A0wFDYbQ03MJUCIcVRIspM/ntyV2XE3qFKugz
fc6e88yVRZpLZMWev3/ITI4O6+anZHG6GtptWCOoLsS/PvK1jyIaOHHDdkAZM0F+
UO3NHlS3xTEgWqSWc3tageAc6kOT42ysI9AxEiPzmTYWLrukXLIdPLNIisnGmk+x
xy0VAJs7i9npn/k8Sjy2gPuaXWQ4ZcfdWtHmghv81/OOvWNTGSMIs6JwlJKiW696
3PcxmOfVB63w6kRPtaYzugDANYSGOmdyBSb8CPmrRjM+qEbL4zOVR8c5fYORu9aJ
1fV1asM8unNqXj9FB0O/kOUae1SdZV7803f8eCUQnJhBIf3XVgXI8iYQJkzV/DdA
Ta2MnXx0WFK9/qsmv6yef3DoU+qUR2xPqp5Zne8TueBbZKdSSdBnNs7LSLP6g79a
TnWybY4MYWOvMUJWpi6ZeWEElsIsedSo9H2zHWRM89/xQ50DQKgm6fY8fy/82ezp
4WrbrqTm43JM3M3Appo0Kvdn1qpU9+U8WHVJpou4nRyKp+9Ex+5Rd3ENtlh3N77C
Rp3XqIRVP/RkZQKcF41+ASHrtO+mREMCLNX5j7oIAqPbPf7BG4uXRQuGTk2n4UDY
jPpifovyFQX+DMyWAQ49QoEUQtfWtp4cEJCcVrsj3Ra6btKWL7CjyxUGKFRsk1w1
+IOEQegM2S1dHvO8DPBHSTGasAW/fBvkzRuKV2DAo7zBuILqQOPhvPA94C0XICeT
83dEuftW1kc70VL/vdFywnEOBsS6xx24NkWGqJv9r/yKg7apNl+rUoXW2fQKhT/V
wcHzoqJzRLLbl09ChNLBC+qBENI1ZPcCOs4uE3QKcmu14esdh6UVQFkzT2pmwNvi
LRcHZeG9/+wfjUre+SCq1YxYJHRVIO0NSYDCM2IL1PmtqCe1EZuFc+Lp9m67jTBu
8nEm6/ofx6QRXRWYWFQhJQ9rLG9c85HGjobpONlmve0k9B0BXbswyJcAf8Qn6imu
B6psHppHOKaGQBNBRJ76gLQkv1G1J4A15ALNEwVDWpAtgAEp4D4cJk4SJ65zFt92
Ri5UOXxuy9n2vc8TANUnValKRUcQlrZVqkpvaL8YBGc4X6qEjft4wMLxmTqIUsMS
UP/UFLjGUeUBLMl4SKl1Xj0bOKjw5wC/2f5lR1NCExC7wAWT1SM+EiYtqrngMTEn
FfBmWWMlsUT/PB0ncN41cR++MzmW5htzxMTm1owntbY62QD83gdd9C6pFMjleNnq
7bdQfeozDIPh7io+EWxzuyV5kDVNdR72Xf1PO1DdKbU9DDKrNfcGuruP/P53lHvx
GK3iGjtyWAR1GvGVu6mkYmIOZNoQlFwXOxb25TpmndLejqOecIbxuDd2PRHZAum9
0UvNZIDNo9w8eZ1zfwiCWpLptD+KTjFuZaRrLAw/Ywy0GZlwFcOYZcMBC9BF+clA
hl3QxxKZV+T4a4mzTnGn8DESOzhZX4CKT8cJPZ1JHd5QabWwo2WhZdaxKZHjzPLq
uU9Yiy7RINdFTzaXU9jAsui9d8jhqAN6zn37zCu/WFB9u4NKOYykH/f4xcd05vIG
lSSPbl3tW2SXeZNQNotGU3PWWo4V8RcMwiDmE6FBG1/XcQrgA1Vf+A+Qiasg3hWR
3pOBmQgkAMAlz01UX0hpY3OrPjq2jIhpfadogcNoFhX/PzQIkHsbjMSpssWm0o97
UOduS0F4/Au1JEmzdi6be3+85NGiZ6tCn5WZ9dwNyStK0Ymt4foEuCnLrVGG0+wF
N/LsOtOEx8jatz8/P2nEtjMvj+I4+7FL8kY4ZQ9IrTXCBQYzZDL+bjLSVMVrrGfd
i/DSSg7vr0ARgTbzQ1ft4DTh0RTWlhUSq7CX48Iv8JcD94HdDTQCJU+5Qr8QGrc4
NBxb2ti+DCZOhVTijU89w7lth1mL7+fJzH2AjXIlaQHPgXjauzSXwuGxEwz+5fD8
V983AzbN8aST7X4kfsZ2jxOr2pPG8/V7+38mojr72RM6Gi3Jst2nt2utkok/2gK9
XvyTVcr2gNdBLNXNKT3Ff/xop1AVxORityetS73KvsUlJ6Y9D4qd2x2yC5lQHCQG
YjUe8vlqs8jJ+Twxkm9Q47cu6foSraRYZLfnZ3lbYriJOHmQ2ZLkOejIWJyQhzvv
A2PIh+B2G49Xzs+Hf1fQChzsHLHtqFmDnvR8BbmfE+pZtD1mYawsm+zrCilJyzYr
GU7OSPeIh97OzXea2ktQ6YNPD6OtLAQ6CG63Kd8AovEAolXK6BrUgitc+ZTKTk+X
eDfEb1/RKE/34ErnhDiIrWyTAIjFuvckNvZ2yhu9IWM9iD13oj/Daxw4zavl6hNo
MLfTbs/aN1FozNOYHOnEeQYFKPPjMC82sbAPGTh1HWKSZq1uqqCIOhLO4r7m+x9C
511QFcmHuJ8nT6ksybCupZeczhad1pOHKgiSY1kDyO/V03O4KfXz188Fu0dFjO3R
mQWTrRmE9TGivAW1fx7fnTBf+QEQRSLp1Amku5ES0Nag7uc4snqgMzVduEx3zZMe
/gNP3O51SHY7i8Yzk2z0j2wLY2Gc7/3VdH4J8yk6FZYHthl4iXFwgZDWJi9QWpdr
SCh0yWRO64G7lc+tjJTJ0bwwmvl86Ou2OWCosuemFVl2hOu6WutVLvABMiDeMoT0
tDrPDNGcFII9nnzGLAs0p0KOtPvBRfDNbAFwjRNEMlYWRlxsQRNzUWINgR7yBF0G
1Ufc4Bs1hCxzuCVAtz5MO+GKWJqIjlEwwYf8LV5EW4YUcOW8QKbYihLl0Ku2SN/Y
FcBJvBLKG8JX9+lQgDxosDXNppxcSARiUrdvONfGc3o/GNSW469K6+j6o1vWKx69
TB0EyUUQiu7s1b4MV67+IL8d4UPH/W9MkfP+Lkp9+GCx/ZyVWTPR/Cuxje/7OCbQ
APnsjtimytXq5KmXWl8mSfE99vrE4pGa3DYldJfAmP9lPp+cZWYl2oLVwlQSKpVH
DIKgDfAZpkPg6Q88OO2xTSBcbL4V8BIv1NAp7uQVrqd/iCrYeMLLYOP4/r5y/92h
yOzHglRE6uDfMGkLb3J0qE2k5A1HrCDWCWK5W6ExxFsjvue5zJ+D1vkh13oBOqYE
uE32/VbMJrAcYfBNMJfb5hZQ6inGNH88c7vpBpjEh+c9T8MuYiMocMzITHM6AluC
xsElNzb9XcoSGbmzl7jbsJ+40AKmPzorbwVVM1BiIWVCwniOcgd5kh/efWB6ZKIQ
J4G1dRy0Wnv1+qN/Y+ZxLZ/G43zX2bMkLuIe73oY4IL/Fg4wTFa0zhiD06W8NdkE
vH9l8x6kpVdcq5BkV0A2qCFBVtjSa6YFTGj3SdzQpYNLk9xOq8PRzy6d30/hZvKU
FwcV1roEMCXPpogl+bxgn63s7FR0ngSqR2dp2RHBRHPPnAXR9guLGg+/KJqPwFTL
`protect END_PROTECTED
