`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ux+fIjSD+OTFqgA6rC0Mc5m5khGG0YOLgMXboWSEgLjERQtHJfNpKz6uzCFjUbQh
CDWXN7Poi8rzK2cObtYzkdsK3BbMPTQX0zYx+eP9XNW1XkOGPkhi9+BxYkdxomNv
UnjKVfOIF+BWUFUgxo+dqTr6XCKOI/q6SzM0smXC1ZIxVJVPY++Cf0Puzhnn6zXc
RhN3+PqBXP8g4ND8cxZMT8wVzkUSQjaWH5eKuQtwE77hEWqF+mGsYfmGMyyqQt40
eyI7y7mj4Dv8AZMqpQSjrEzrW+dgw3ljojhQZKTSsyQ=
`protect END_PROTECTED
