`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTdwslOT9x/FOyh86RuqukASEGS0Hu3kMlcJBMM6zdbDZwQgEAnEBWFZnRuGbnoG
bogGJRfYMbfBMtrFQTmFJBhebvfA0PZ78/s5+9uJQWiuFLc4pTxCjPc2o83Bl1wg
Cm777pITjlZBASYxMDvbBiy4nRmGn2SdGTEXWVmFpRRm9tsj0zwnC+y9tedOhWch
CXNsqOx4WwDp0REBaCOV/0ingUOf9LHAw2suKtAetrq+5e8dGLnYnx0BSlZKC/UZ
L0fV6m3Y7SyxE55kgYjvlw7XDpviwEuLq3teAKUpWT5JD4t+WLo93XXKTwHPF0GL
ZloXGAtfaMlccswoCAR6NrF8RVZvwyAhiJuFFeKGszBnRgCHkPvitn4hADbMAbly
XYVZqdrDx6qsYUM6ySZYPuMuKlKp7gImJlrwuqeqdl91uelwd30n3Ejc/Ccp11cy
Z1jC3+lI7kqPyN7ABnK8+TMqkGEgW76ht0eC4czspZd89CvPUTFP/kMvJkLpTpE7
QHu25/1obmliOHu0aYREFFPuHXR1P2OIi4cy5Ye6mn316Q+H9t8Fv64Vi5UqVee+
Jc/aru4T2pIMKsEIREPDRiZ1Dt1dY8RZKTzUIOqBu8KB/obW7E9TK1/p/LL/FfKZ
xKM7RMSMQColfjg7NgOKlN5KDnKJ45BlBt68hCHPfhrDpk8vwmPa++gnBbK2L4Nz
mL8diRXyy857vQtCKrJK8zMWKBe63KcYxzCIF5BLxufyu0rT5Tc3TDRJa3OAdxcu
Hgb7zvRIKnwDzLJc5mnb8kZDVxv66IgHAuBISWGD3oyJT8XVvzy1qBO94ndh3XTi
R87gZLFq/+rfAwUnspCQpDXrorktoGYamp5N8QNEkaG7uj4nJ/Gvp4EdXYIoPHok
x+SURY/tYeadyrq7DSKF77JxYBzVOdqHsqUPUw/+35mpDR32LduM0mZIS/Hy8Di2
E4QQUywDQoZfTaS4WKxj+skt2zVeB+wXSOnJjL+3IeAC6Ve0aVJRGsdNxfcGenBe
lRUJQb6tP43llqe0YaI+mUBbq8UVYIK1EGLx4Dd33PztKrNrrwCktJR83ym/yaqW
AF/b240ll4SVi/DvEz8M1KxefwbGhwXbxoOZEeleZL1jLvllNkiUois7PKJIF1XY
xnwG+z77qtLlo21aylCW/yDI5LQuVjCvhkEu+FB/hDQfBx5lV3vglR7Ixb3YhFzJ
0MxuKgZnuD6FUWXUUTIFR2c/rJCgVGJsLuZY8OcyAbvcuCXUkDm1Iz2q2D25FLCq
Huds+kF0J7b6mQopXQXXxM5R/XYGb8+ykWIwkS5JFBhdSa/EkVFGFx3A6BEWbf60
`protect END_PROTECTED
