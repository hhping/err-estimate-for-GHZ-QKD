`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ixnd/GMoO3OUgnWaYDNEudaKFuFdtUAbntaw5NLkur6Cck1rpjeDxKf7ZLrbEPDa
uZvm+3c3+ce8vi3G+Qx2vtJ/6f3y73UnrIoSn63vq3sg33sHuHy4bmCYBqRamaOM
dmQtzLCUoW8EOeIr+f//3QtiYZaI7CY4aLeD1pM/FfTXFLdb6FzGE7baS6tZMfRE
ZhLar03+ahZZqxd9NMd0zIChZG/ohLxqwp8JZtBPqpkb4m0TaC3msSTwihZIOeZG
TTq2YtjHDD7DxuPt6xZY+w9uarfrMiK4o5n2Q/iLSuAwsNsmBbQNWtbivZCptGYi
0+3IrnXwJQa970cWXo1MeSUgSrI0kifbPud8MbGo1XgwOtsDY+YwWS/BemlVTeZF
1f8Uo2SoYPB8tToanl22+shL7rXx870mx4o+rOa9V8dvPypzKPU+9A8LUUEqXwfq
yy3FAyhTkOeqH4pJXtx1L0/Ksn2irkZHo7fYvoYr6O0lRw4ry76jbNw+cGLEAIg6
8YHcvwB5z6XQJQ0IpcUXCGcJ+ig8W3k6EVIFqjrVE3PCBka8+R3ntOjAhwSu6brq
I3Dlc6UzNyYtxwsjMONc6Ihn/YJMjoqWE9/YWGMwAHe06f2IeobWgJWVkWk7Vk0L
d7jZZznlq+ymKK2goVl6tX6VmGEebmOa25BZjOSfyYIU3FE87E7S+39B1j6Gks8q
omSBfMT9STDYe02LcpfZdnwSwnHSZ0MOkc+Wzj9SBbAdyuPtXZPr5gXS1h8/ig1C
id6rRAkJT3meT9eALSNvkFn/Io9GqYqRwmk5ijWHzL1GIAOP2Lp0Asbc26zorIJ9
/hf7WJJtSfwEAUovx9IQAIvPAtE2iKHMP9e13iNXf9CWwf+6l8gckZeagW26OFw3
VK+GLxJLaMZ6cyGykmDNyFfdWG4xvEOvBiDeaw0Hiew/QCEYInlxsYbibVX0z9IE
rjh3Qyd9qGF5EXux4VuU0FUqBLcCUGqquHqAmv5hXdhpKjNEEAT0zhLgrONRtSnH
Q+BvTuXXeAbrgcVdeWmhmiYHkNhQJqcFQfL2BDsAvPS/1EGrllU2QBc21p6zMzM5
95GbDPdCJ82Mzo1EUfZMQWik0cgYmV9WvTM9VJ/miO1BuUPvTVqxuxn1NbAo89R5
8bbZ4A6we+5tuYqjuu4BO5r4/VpPfmJDuDio3XBEPAlJZsPhNt4GPCGf/Y+P+aPv
l82GTapHORCJ824HRzBsPAWrGeOkXltmbPcLj3JV0o9TL/HaDQ9M9/IQjylUgT1d
nlFI+QyATFskxtMtz/AZ3jkblF8ScPaS58S0F15Zk2B8gQ+Vkq/ZXANZ29G0ohqZ
kQfh+z4Z3YUTy7sWWntGcBVxOAbssIlCJchZf8rK9icgHe2Fnzg1azp6rpQz2QLa
+kEEFJCLmdo4odKm03F6KcQ5oTLtA5elQjjuCRQCuQ1o+V37j5Is/rbPVrouAPze
RaLp0Gc/LHs0LUcI4J0UsJOKqx4ZAuNpsF+cGmGVJmsrmuEhDQ0lhWVG+eumWqZm
DIW6zK7Ucu6E4/aBdD8qg4hgT3e8aCN5htr5gHHtcyf88ME1n2ajsBEcbnJjL+fa
RB5bBJHfgfN6FZ7ZZIfI+wTjxHT8Fu1r53r4mYqZuRB6L4gX0FKgYHTiP7GDv5Mk
GXDKct3Qaktcl7lxhMCXohLZSgVAaXe1ijDjZM38XvLCnwLItN0bbLJqQFbMpyui
aJEeI+6MpQ0RqNFrOI+XEqH04JaONMrrrYq/GfHPLL2emnNwIJWrbKX+WztckbmV
F8iorprejJ6kPBVGV3Mmz/0ISLy9IZAmWc0Mr2zyuAA1vRVh1DpYS42FZ/WM+lBT
oLzg9XqHZn7AAHMzOht6lBAnV3F1g5MuMvPcUcJYY89e7qvWrv+7ftms9WiLUOFj
VZjA4QB9nHGEtgbCqttr195nZYZ38ublDAt74gPhom0He8TdbRPmTrUU9/SlCtDv
TqTyTWGHZEyzZaYTFMHQp8UQPnBDqCw0LzsXJNmQDcxDhs7FqxC+pt6Qy2TeJVSf
WBtVYTYIcTwGiTuPV+JwRugyNUDd2dh3lqBh2uLqScvENVn1MS0rJe5+ZgDkTRVe
HAmnNLiOSSmjk/8n0KVoo9JA8pH9WDP+0Hp23nuW/iwO3fKgqPwwr3U2+h+azHfI
yPSFn8xipz29DgfE1I23kgNJzD3RAJqp1ikffp2awJnScN3B/KnSK4M3QjlbVAat
UYAxXaIhPr61uN37PCZkggeye5C+UmG93LHSKGQZk6wvXo2OIgrx80yxs3B08oK4
7x6K/KKDHYdMDd6Y+ea1hKgxExXBtHPQkHELxfudOrehPTLOHEibn3e3wMGun6DA
+t/Fbz34epYcvLtXp/nd38pRqW3Xr+goVffphfNVE/sqlXDLR2GfUWwgbOcxBDZq
uPfIkQdqtzoodILIYR+TJlObxDrPAXmSYXUJ6VAurYQG6gDTS2HdJ5GtLntcUF/4
Z8fC/3+L/rLOaRgDQjqxKMa08dNG7AWypmCFsW8PyOrldolMZwC2N+T+eHqf9Rn3
CJStqxk4HGb3Tb8db105btfN23B1zXHnfp7echAR9z8Rn9WgGXjTNM/YvBpS9jtM
EOuZdAkwPnhuwGInHJ8sUUEZyPH5dISFFI+29wCekLGU1bWNIS8WTT9RYnC1o86/
QfdXTVpTsoJBWXB5NQnYz+W+mxfAcpqGkNuOZlG0KZBQiuBNhVZTs0I7g5hT7piN
m9Lw/YFBZEUNsu3wuVVShX/ApPLXN9miYUp56TDc5MXfv3Oe6mkFqD4dwWAbEqa2
BawXH8IwEEN73CJDFyPnuowvavo4zXEvw8uHorKlrX5J8n1WwPqfbdSsuboIiqjG
xXWUbR4B74s+Rm3YAJqyZuwyGVFXIr/exa+y8rdEe+WQ4jLc1lghm8P8gFlIOF5D
Kt1TaIh3E0T+WEPD3m9dL5ekEEG05X2ZjdCUzMcWyPj6gsBfbzCo2FeDhlUnezSQ
QTtbh8LMOYFjeltOWhPQbZMQ1JiwUAK2R6bkTdWCOH45ounMp1YmO2PgJkZDonqf
Ke4nY1E9mCPWGj4tlTZjsJte32onkaHHM3NxcW0ltdJpHE8fx1Fk1oBldrb4BZGZ
UzFm3lYd2/GdjGpWrNWjUBUpbjt0Vy+Yhf87QcVYRs1Hk9oh4P07KFuL3N596Wol
FnzBqxqhEYu2RTef2U+dPAv2Rk9AwRuInAA8tFEny2rv6S2nLXwQqxlb6xUhTKYg
KRhL8K1s67fK8XaHVUR9VBCwTXuwbb2c5vv2QLCiE0tJ5IM+izQLiawtaKDfTkju
vlIg4Xzr4N70wZWLfO5AfnHFItdTu3tiZYDhA6UURyKfnZJnikZQu16DP0HbRVf4
mdlLJD8sl5cNNL0EZjzYmku/1ElIfqkx5xcbMYNDy7W6N/eU01cOfhBOTULaZIyg
qiRoLfirgNckEDIZHopVX+hQgkLdcsLl+CEvm1QL+xbfrivIOkRLxJn62tst8Zrv
cLm5AROXyCTEGxAAcl9twUoBhKnqr6p+IP67/yrXA3kFo8N7530rtGP0plKRMJxf
50XTVgu8uyfCikrF7Yc61N4dFBy0VCBapzcZPZdPAyhuaT0L8QpTGaRVylJNzsAR
stnGaRUqC9GF2nsCnB5XwNVJKH6I6GOyi5ar+tFfQzBANFtAV6V0eaakow8CZb9b
n8kAP5F2R2YSpqKmFKDQw8hj8LPdVHmWXYJ+jgsalSrK59cxuMYJR9qiVkMwMZOX
mwd8xG4+7ylJACE4vQN9Lm2BdQsSISB6juS5Pq5zNYr6mECo95qQUWeMckCwGneA
lhOwj93vnF8qT6zVcV/u+Dn24f6Br7X1HB6eQ7wu/0ODUfzbs8jEblvoYFf+LeoG
whf4Tstv/UeEPuL/GT+a/lE+h+jKPhI4nPdJXCs+BkBF+xLnp4J8olgCSnjUqtXl
ms9YiELWCJ6AvvQQJMj1fUG982drU54THQv5E6+S9ouUJMpAR3FJGa2n5mp0T+Lk
9JTj6eXZc+naqgwONu+xk/1Xb/JlzmbqA/LE4UEu5aUCj6gD8iDnXDlp9PZGrLK2
nCAGlFrgoBMW95yjFXeCuEmUTUEPaLY/Ve0KRlNIRm6+D1ASSSpNAjc2vIm0Uquy
Q+Sj2McZjWfJhFNuNeVQnDYaesF8qwDMGfIZa3Dg5s36FUISQbp9SAbGiYcG0UKv
BF0r3ipuYP8cN0AQ+d7JdR1ntbSA9NTU+UPFyeAakcvn/GPvp5q6ZqminUXDcVRq
1MhstQXzGL5Yc+nYrRxm/2wXZ+Ybbv73lqhgX37l9Jh+l8EDAhMj9ZPGqlXceFqW
cl8kC1gVFP83elVD3RuWhMhqaDZgSSrPFnGkMUfb3+GkdCem8+WTIVGKFhFgnD/+
a+PDKKYR9sCaXax/IgpqbWPwb5L7wzgVPd2SJ4UihJodVB98KJH4KLBKx4vLai0D
zAocz6aOmp/zfnTnBaODtFE9d21TOXeEG83+7ZhKwToeUHyjF7ADpj0LqfQBYgDb
wZOPkmtI7pqNTT4t45cqKUdmbdDOSHSQuZqslcutNT34v9c+nK7/twfcv+1TBubC
Obfq9hnI+DCX4Aw2ftcXAOQwylnDBflu5jiykbWqLnlpdee5ZzNvsaWOcZUKMLch
M8dprK2NolvMl+lyTMjQsLgwrAve0A5kt/gcGboN6bdVAiyY8cDQkKoJNp2NGXLr
r1zkyYyUMAS4To8WiifHU+bxzIwot6ByMn7P/bJinCpefQQdcbPrTvsRTM/qHEO4
Od+xCjZXPBIrk/8H2MBvg67HQ3ujyPVw0EIJhsnttzGdFZQM1uTVHfQLGUbpMsX2
Ki+AmEiQpdImMXRQxFI5fYW+itab5Du6jN+ux49EdgoWo6U1i/ZUWpamcKunwUfA
ZCQgqiVuV+tiPvz/WD4WFkRvv1KvJi3qIM6SUhQEhq9rTF54ENPoaKTAKKQKYKB1
E7sPBukVZzhoi7wgn1I49bM0DvjhpSg+0IuOAuMUoKucPLD0eIZ74vewXPaJUgGv
IGajncsKkPm2vtAEMByw9/SvKaJos+UV8gM1EfBCmQBgTjZP0tjTYQ3mduOyG+/d
jGjXTs21W020M277eut0K/udu/UJ7bmj+Iqk81TqCaJZH6U4nh1ppXlRx+pSAmqr
hia/mlMo1VYlvvxeRbWvzBGEUYrpDKd9pHheBPEyQAg4Aa+TbVp9EHmqcz25kj86
u3qCrU+OunzcbZQWCAyFCbPO1kQdfA2T298puwUzkze1idZObuEtXeybNXHoQxgd
Ln2YqqJQSJBKaS7/TOGyUCFXHgahjLBe1HDmrY+kWNam5lyIHwVBJxW9NtFoJdHJ
Hb+N4lVfkq5hC3EJBU0qvkBAAz3lOpjo5B0030S99arF2Kju/aBMlGSfPn/M0mWb
kOBW/eKFb2z2WEuyjrFuW18pex1KbsWBYlM22yDH64za5d8OqI18kDHId0x22e/b
jRNoAbuwhQUU8k9SZWtibYkYuetLCfdFN5spxjADrcNySFf+KFg5pdxPEu1WD31G
F7MXHvxIJ4cmm9SC/Zj/FmICJw0PXmIXCNSGkBpJvEjywjgWWByz5/azv7sM1OhE
S8+7Edp2x4YsosQJQb92OPCpy+t4FO1StApaPXS0azQuuSYyaj/L5F88KWeTREQt
SMauD7zsW8Nqmw1Vc+uiQ+PEz26SoNvZB5lkd6kXrcP109AwBPD92pBdJY9SLHrB
9B7s2Umc6qf+ubjUYHWtSSeYBVmOY/RJhUmfhI3+u4f8JAu9sMV5E9t7xNz0Pyxn
RnhyJpqrqkHle8OjeMknxuBCVR1VexMGhmT2jcJY8PSToLtLnjbsO5cO7j0dGHd5
kCiKkBBupVHIHKRj7AvsiPaoTbSpZ6ym8ggpBxhas6sLaBHs2a2iljIGg801IqCG
tk5aPx2WVddE+3A3kMJs3NtWPbJuukku8h7D2u5JacPwFLZWChV/7cG1t21zrb6o
2SGmo2uXru9LChlHqB911L6R9Q/jp5A6WnmTJVBaIxEY2qlr03WHo2N7JSp+SVOt
jkpPsl/1F64ool7te298Ig==
`protect END_PROTECTED
