`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kObAXrVU47ux+mgjvAErtRpcGNRJLR8IXkv/qsyX+6313WO9ld+STLqeHvE/JsRh
ZlBHF9cKlJYfZYpVBgqX7Rf95wWjFc0KAHekaGlBHJHW/BVux5fh7SeYWRQa4xMH
16l0i3haTEQkuXhXC/wecMS2Te8KCoQ9jSj+ycEUOnoY7MWasK0pU12pzRkDXQTe
VhpWO+M53HKHOk7TKoLuEVu/AQJWjrMuOnf18HMQ9oAA9IeJRGVl0d161yqzMsVs
6I3INqT85l6+Y6T/2vu532B4z3yKYqFLfEgTDIR0iCJYxbDAWQyIoyekIJOZbG4T
rJz8tl/yk8MzjY83GTEL+SOPNRuHbLtQm776yLyUQpQJ8q1fWTfwSrsm6T4BVLPe
9uT1CaMsfA3sfBROSzbkJfFC2CTGYSPpgyGfrUBDOOTuMlQvDkBCyuZnBovFgjHe
3qmHkyDj8ifsG62kQprGF//TjdeARLSqEEtl/8VFAQeaWT0Vbc7XbJ60vp5zZKSY
PV37yU158JiFDtnuOL0OLtaJW1uFBv3wOqlk3kq/NDoxMsQanMG9ZzlHb+uX3z4d
vAgeiLaTqZtkOOA2h8DP5VR7g1Yq9ADhSHyQzMF1/P3pKVa6oZ8hLCH2CwvEl+Hl
4RmJCM6bpJajJGcjAWq4taowoxSx6UGHfQgpCFxOErAlmHIeGAFW5RqpjSQOyTJy
aJ+/YWAYWsdm/0/iu8pLtQTQSgytthFb3ooBPrVAd5pwx1KYbTodHBdpuTrvXh9o
u9yyrGrblZH6UTOnhpZGknYuq+QBZdWATCd+58YCWKFIxMOzv6AqTA1WtiQH97RN
79qInMDmCN8LbbqmktCj1UfPWHUgeSq5QNhbF10a6+OuMlAq8Y+rJ4aK4UX3QXOv
mYMmAjaf5Y5tXMgqaunml05m0FLlLz5NIFtTDmNFWu6/dMzGwv9CfZZxwp3pQKys
OpPAmSV9qkGbAzgiVGYRb1LfFOTL5lgpI4wBFgAbLOzdQ2aYb7HMbsuJsioXL+VB
hKa/lLHchnTLHmx2nDYkIzR62LfknBVCikW3z8GOFrsAhiNgvDC12mJ1iYNww+M8
ShPb+qzMcjPwfqyGuDtYsQ5hHxK8J7jkWZejZBYOI8JkSnfYXzdUSn6LCavhaNJb
Zp8LXRMmQremd7D5BYJuAoBCoHgWIrEKgr/ssmwxsI+MhmUAk8vWcpcexNiNsjlp
gsjZqvoFG6n23IsOu5UCZmj1zxEYzIXQg6sqnFquSjCsDxeNQdD+2SIhh4FmLUF6
yLdndaKan3cWV65b6wfTVc0YYwjGem7QltaLaqBrWTkBo8wRVPvihGlMnEoOuP/m
n9lkf8tt9bYoo3ZV56nl2fnpBvOI1NcE7lp5qh1HxKN/YdWfl/9ltWwAaSY87qH/
YY4WdD2W4ovhTRQfvrM4KgF1Uqx+iRANXTBEtI9wWvw9rtWW8fdxMkbm1nod7AnO
emhJNvmcW+JdVXQpLQiCGHPT0E0Ee05bt369ZvAXKl5Fo6TB4tuWXLtl+Lk1W0no
PoOhLP3Kcoiu77KzdxVK1wuVOPDKR8Ag4Aif+K6xoASOi/wZxKyEZM5huyZzGSI3
t3NH42IgS2sSAtMoAVM/uh8Nwvumxjz/cf/DNkrduut5V69z4+EAG+pYdmMmpc3C
pjiywI3ccMvpSFEgElq/jDVhZipOCn4Yf7Lk1CmHTW4rOrkW9HASpIARWG9YkIPM
1n1ddMPlYaOBvfqLq/piYc7Ojw1neGjMmQ5MvXQfRtv7YC18w52V34V7I2Jqidde
VA9CgP/e9wTwXS8NkqI4IOgXHXPjNzBMithvP373Hv615uDkbcibzKoNoXKAtbF0
sDVDo83iOIexN1i5vibtw5WunPwMJmF1Wd8M9/VsawY0fAf4TDG5J95ORNdKAA+I
iW5pZ/tAIAdw/PgemI4FgtFYEO1Ly4sIHSvkCYAYQWeum1eVNif7fQV2xYCwGCyK
I/iCbWOoGSP676BLBklgXGYe0OBagGtvvUCEYps9HGu0P8jK3Yh0lNw3gc3O1pXr
drrqsh1V3WNor++awE4U0FesSsEEctsnDJ2R7I13KQC5/QaXazLSE5zU8thAEuFi
nB5aeu+utCp7eH019jRIWq86o2wt5uSf4Fcy3TYBsMlN/c2iKhOoKJQYC3m4s56I
ZLb2vVUO/0x90Botc4I3noLJXAQl3F7XTqyGg+DOowDWhmk4gNsQK42dnM9X1YhU
RggDgDk2S2u9V9wPTCkESdhmDNkjccsH/dU3yUZPcMwZSPG8npODAvwTy6XvEUon
2gZuNEhJN7c8lK7zGAQJJY9lKdxFI4ecWAlwBIgvGMq0EXIz6SU95JiMgY4m3s6t
2sSnUP58a2iphppr7jfqNBs7j+zMl+Lwn0gJ3IRQsoOdCP3CXRxxh+DbNkK20hA5
MGvdJDOpb/Io60Hr4O8Ca3mCo0tz/Uv1sGHU3XBZ/qBOQL/x+/mTbSJcmFfncT6w
Zcs9dQWs4szNvOlUcwfB9odzA0VITNfRLpNLdgXczlIiomfUJGzqBzUOQrtlFGrp
QnSLoAlUDj01METiOZIOItHBWnG+Zg/aKPTVCo7gkcPsEGEe89UlltDVDlVhJsdh
uO0NAnN6eZap/znYJlK4zXZ7Q2ZglCN97RwISixW/FhLVg2lVrEB5AXd7A/khE16
`protect END_PROTECTED
