`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKIOUbKiW2Yayp4tzqVhZ2EsLZ7MKBa5kq7bqjCGUdBt+XrR7oWHPdLlAnQLBWqr
gFkMi17KLhuvbgATaMUOS+e7jtl2mqMRPbo1u+gtOiOSy3+TXLFZvbmnc3XrgO1E
ro96C1l1nDfxnfbfvEUcyI6I5OmhIsHxCYq+43DRxZYCID3vICKbuadfokR7xUvj
Ne2Xju3os2zeII2xmXW1LD28eKy70aUwwgLwEMtE9vLPae3/e7EPXsW6x8NrJ7ta
n5m2o/yrndT7QyjogKpY393Hdd9bSqvaXLVwJNPOtkqVSP6reW3vfk5RPyR13k+g
jsQXWq+9m2lvhc6NuACWHXouEEeN15dLcFlch13/S+rD88cyor4kUJMUargeuVxs
kIGqLmH4/+g8v6Q+T4iayXWo4033MhiDhZm0ZezptMraklFKRWKHMcQ0WDQKtAOy
HYV4fe+5wRZLbHlIJ1K+kdA31i2Nzpd7NQh7QKS21Gg2VQGyspMlmpauOM4o09LG
kOwJD+R8Obh5ZDBIkRQ3jewZLAsSKV5LCynTC1okkCVQOSoZ7mwU4XEhfTjKkMPQ
oc+ui4UTSHs6m6JxYA+UEVvyrWrIh1yyhH1Dmz1V+JPPWHA9YjixbzKFSAkBNYc9
`protect END_PROTECTED
