`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDn9hSVyXYAzCsVXXhbaePHI/xLJXUVVHMmm5VJYXjrf610r634KjHv+auVGf0eD
aRC3eEzPCvybdpaidgDMSsk0ra88v52mTHtF1D+QuGFimFRauD6bF4IiBYrjHrN6
M7/8Grd+WEM4aK3l6xuDlM4TQQ+q79PWEfrNkCLt+yoMyQaRzDRHy9SLKiyprhxE
QjaFdbdQDoPU/1DslcFDE94P+Ro9PKR9q8jY1DThlwljEAKq7EmWalSFQV/rxHFL
swrZKxHsW15CJhcb8Kjg3Z8tD131p+ea7lidtRGsNskAQZ/GvzJO3nUuL6neg1Bi
pewPw9nt0P0em69vngEJQ/zrO5sSFE6U+/RNa/uJWtbBg3Rbun08fjO9leEwYkEY
BQLOIMDwPtnkWoKclOw1L0F949ZKLFiiIeVxUlrVxYcAOhRyQZC8bqo8IsfWUSSb
M0oZota/vtDDpfxXgDsU2ijOImN9c8G0eUDMgnrc+sxydEo+6cCAswEQQBhZnKQ+
V4UD+J+oYB0nIP+r1M1iN3H8VCmXoqsClq4DzNo+cn+5bGM0cqyshovksha3Z6vj
sc6Eh+puU4gn6Tu+qj8iQAYfvN3Iaomwy77FS05UZy+/Wu0QnmsKLoj8Z7kDxywQ
vCF/1ptVQDBB0jTg0krbH5ucRXkZB51hui7YLmdi4hhnP0zcUbLDJrqkA5j9Br26
86OXR1eseFCOaMyofzg5mUQe8jPGeQWVp+445rKHPBLbHKU1CmYEASsJOOvQNwEP
puNye81vYqT6NQiu78Ie7gHnO5TPRMO/ctXXZdIGS0kKptHersD4xVeg5SHAPWD+
oWoJIwJ4MLbeXiQTlSnzSQIkqSHjbfvJZ2HiwYn1nZMzGUzz/pxO1ke7BDgQOD7D
agkRtTCOFvsn1vlhCp/LkFNhSd7Rh4dHxyzxiOoVwJr7VfAs6XbWq1FvzoseQyxM
9Nmpj5ZvRNDuk4kGlat2g6uKNUfoLuOhmOoiGI5NN+lIdobSL6Pg0sKacStOOsCX
hkkWT47tWebwoMSq2NX++WPysRxNw6vSVcPZm5ZpLuoanolr7NI8aEIIJx9k2vFQ
KrASmn+gDFUcDDS2traQ7fOt6acLn0Bz0PD7oqXQMOA9E75t5JyJ2wYwOqJeWNQO
kUjOhyzyeAkKfTIdTHbKMMMXIbN6hejrQCGMmTAQ/vgCjmxrxMiwZVca1x8RXKbN
//QgFnLV3UtsYKO/dj7HZP7hpPSZAxAH8yutpMd5U9R2THLYgyvnGv9eJ7t3vjn5
Os858HUXgdsOB53rY315VI5NfFBN5cu7+1ljveRnfcSQXaFpR6KKeD/GKMjm9dUm
JXl4+t68/r+uNuCtmidNl0Btr7yvtvb5ulo2Ylu2OnEYG1gPf7Z9BraDyq6lTyU+
Be93g9Qxg7efeFGTEyWfrAiMsHx7/ETeo90JsYSCVssob1YAr50A2nZFfWrlDtdI
6DUxxo6MmhBXestB4CL6IQ==
`protect END_PROTECTED
