`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVAw9TZvvqvmB9W7A97nG2e2+VehGLB0q/3Kau/ICAVTd1Y4Ad3w0IytvSTGP4zx
uoyh4GW08Rea1OJhahgw8fbCwD+/BPo96E63oz5x3Bh8D4b9KhRQ41b9JT/cXNa/
OF53nEG1DhxaDXckKW+EhzQU5YEsO9hDCHpHwr900qlCke8Cpb0022rZT3wfQ3UP
MzzQXJFUNMgQZc+68VINAFaVazlSsaAchRTXP1If2wnJczm6cpWBU+KZ0ic6F8ir
q8ebWicvAvk+4v1ws9bZuBb9j9TZI+2twwDzxppiD8QA75/gJo1YJMowLvV+xRR7
oXOyh2EQkEq4owxykq3bJNSGDN3Wy16tDIGdmxJIUQ/xUWdtaJiumYWgaPxztv/c
qap2UZURskOzgFdKLQSOKEmM7vMSiQCSXEvmJp4idc6R3cTIynH/CFZytB+ZzOce
YmnwjK5T8pCjaSObMHDS7iqsZBUSvw2RtO+waMcayuQZ+b70/Xl5a9usJiTTj32x
dO/xfgcMZ8vhb6ff04R/V2vcEkDb81tt8zovbpwiCEBCi/DZwTBMMqbkTgGeD6x+
MD552h5ynGJzsRULuYSg0Wr5wLppNGCCpQC4z469CbIwxU93tuOT4oyiKl1WhSFw
buG7de4gREf3gMLG1qdTSFv2Ydr3dVHBaju6XBp/3GVV50c5V1e8BijXTckac1NU
Ed6Wr+Ny4iRSLegjd3xT/9gjFWjZo9/oKZujXVNIKPml6Kf03lSif9kL1m3URLxR
wh/CTlCAgcQ7rdD85Ur7EnJPifdqxLRxxKGFXgYkWC0=
`protect END_PROTECTED
