`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pNGSl3XRpk8hiEqtfhp8v2Y9mCR8kZWDmkVMLwNr9Hd5qjFomCTvBtel5EXYKt0c
UQPpv3lAENoWzJUZuBFDzvBTBirEAgawhNLe2wxuykZDDUzKHH8C+JfNSRNupYWT
WPnWX1Pw76Pa5xV8rCEoK9Uud1QNtHOi7/fpUHu4i4orO+CfOd0aJ3y96mQNk8Jb
OrijTSklqo/FVTaCuDtmkK2pR5UGewR0kbvhysUtJU/CvY8cdv4PqMfKJZ3YNgkz
npartmQMAp0AVVP4mJ39qpulBDmmVpoAd+8mjwfBnsI/Fj9oChsPPbscgYgOe2pu
0nvQh1wAahgmQQqS1lETtLUG0F68ybHSRZKFTS+L/jFNYbYQjmAXan+i3VxKnBSx
5E3H99iyQAStt4xISWotRe7CQ0+hIdPs68GUWmcws+HwA8kVal2pHwaJtVtLRTGm
Q+UauJ1B9gBiF9fD46PVjfSCn4YvHzthX95KJx9rdnhJML4Fb4kZ4FKJnV1voP+f
hxZZ2sXHnknEYo6auPTMC5aCxe+D6iztrMkCYOj87HSyoxBRHUvEOOoZDX9+PnR5
mJC/uGpuQMfnWQHlFn9HJIQnwLa9VUFFB7Ar0fCs6BW/dmmJp68W9F2yONl4ROH9
nPhNXULRLNE1R81t6g1gi4o01PnxTcYS7lUMpANdA7t3XfujwsLRHk928VaorpID
ztBI/jErriO88JF6SzKl67RFyWp3OLnDP8a49vxNIsbUbduwKuVaR4Ik5AIqD1+d
/OlFx956ukSY5JByJ8aK4jH6OCyt7PA9l7AtnW51YonM+t0kMtIJ0Wzh/S/3bmwZ
69eGvMcx25lmnmnur2pOneuoWhTuioeieRpCVgxndykAlpR37ccwIL8QPf1FJlDD
dI9/XAUeyuEDY0DF+CsPl0Lncku8IUlE5Voyf+Pcl274RjCyaiTtmbzy9H0CVmXO
0uxYP/+zAk7Mnzx25DvrLJFgBiNRmrGFMMpRQYLoHv90Ie1JZ4mY5VDI6AM/G4Re
8dyqtfEF1yIqPrDCAsQZGlxNbBsmZmfo7BfdaB5Yj6epDDjhk5gRF79NRp4KyHSu
nuYZ+b/MPw3EtCUuOtENv5ZjGVaYD9o03FmWp06FT9MKkvAtHnXRfy91bDym2KNa
RDcUwrpkgjeksGYi6ikhKlgxIfbTCMG2hTUl2uJFgifLANUOzI8exhsb2an76qb0
E/pvxLjZU8KkAUJyxqChHPz+rTo8ptjrt+jd9dwMLj4PSxe/uz2HB1rSZR3ro/h0
99+G9zfTk2CFPL+H8t1mOZPbubXfhDWvpwr/U8P1B+Vc9E/ugs1kjOh+9cJUzN+q
Z4ISqoedItC5edwcrVNnRMZO+hEDB/zjy3CKondAs3wgHxreZeEPedzDo62esICi
YEJlciZCmSDPQF/nObuBDyGrE72qr0KjgC9m4C4jUvEtoxDT/E6ncwsMwlnRrJ9T
mVet5mowggJky8XKJq/bITNiB5dGwiggbnbzuuJ4vUTOxTSPkbblh+QV1flpxFi1
D14RkPGHipVVao/zmuYx2smlCiRSinHipvS2zEe42Ds=
`protect END_PROTECTED
