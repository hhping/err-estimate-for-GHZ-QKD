`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnCrqOM3FH8omK/xUHfJo5nHAOXwsU8wDMbMDiGrnV9nNQnaaTBXEKDkHuEdDr3m
OUfmWzqa0U33qHStBVo2goq1OThSrsjofrK6Q2ujAIn31hBMMSsgRLfcCxxu0gVn
QmRuopyTYJkTSGexDIrnqU87KWK14g2isuNMSNpLe7UCPHPKb+yJ/s0gb0b/dIRZ
pkXd8PEctyIj7Tgfy4u35kIZBnGSqt9CavNlhI0ylNKlXz2QVxl8+MkcLtswOTUx
2khnFyoCB7X1uHUK5D3v5Pweenq0ntKe/NdtqEOwVCP1tqzwUW5Bs506wOLMGFG9
LQOJBjUh9hQXSccG3mT4LwJUT+SvNNXb4d44oLzbBEmQL2sU61PbuD+WObLWeO08
VfiSWNHUQ1olIb+LLPwW/uAiU/SzSx+2Een7h9GBiBfJO5Z2vOPg4lETNvalIk1O
HGjThRfRc4JyTYTRPffGQKB2OVP4r0RzoqpBwK+UadxqkFY1y633KE9Q80JQpAa8
/fhsMTY8EmQroAxWp5DYdzcIpkqiYVkA2E1DRHaLTzyxx9N6mhh2CEOhL8uL5DSO
G04JT54i/WMWZDv4yc28o1KFFCrTm0Sy4UuU7R7kl1rn7WQC+IRBnn5jt5VyFKiN
W9TOMR9EorE4XnOY5VL72g==
`protect END_PROTECTED
