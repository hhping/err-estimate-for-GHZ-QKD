`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAXPbsWX+rNuXeigWUXv6MUCLztiw/qSJLWdxbVpNOqgYO0ouH5o6haQrKTvBoqh
xQGoFOQmAH4DQswvnhqkMUFaRhTFKnXGg95hKPhLDXc1snnH3BBV4mLHxhoJ6Ckk
gwPKhUgLnzSqwBwEmb/8zH1GgtHfMqyc9U35N+nv5tdYdJh8LA06ttntglcD+CwY
qrkDl10/271545Mw5KaIPHagZ9ZFvanFImGTdcKbgO558sB7hGuNZHIJWbO+FhEK
SV09VyV66+xZU6+lKBNVZ4mw2xOqAg8jbcu3sVP2XVeSiqszxahtlqPE447gEoeW
GZ9XXEVkp03w7J31VT/ajCQcmVYjOfl7Vv/8/UrDIrMQ971bM1pg8cvdHSHH91uR
ZpqhNdisIwPVw30CatxooA9H/ZqC1hz8abaL7Qd+PwNAUMKYEWwa5hdcpCApBnSc
wZF7BaLOd1TbywhHQHRqco9RKl/vKIaUFqapqQGT2gQqmD3MUxSnUvd1AM5AJUZ7
HqD0rps1Qfd/hfmVmWF6g/Ac8vZWZYUimhr7SwLgBKIVyYHmFR+e0ChigT5uLMNV
vtatdPedCzqeF+onGOK25Z8UDu5LQQRNo4dtCRtOPXQsoNGXVyVzeKgTCTXpjlfb
tJOKWPsaBve32WIjl7Y937MjPitBCBB5LOfGzRumbjD2Ci1/lmXbuFuvljvlpiUZ
sB1Fe1+40nFBzel8puZ4kxFEGzFxNf34elWxS15nIZgT25V/BUVncoPTJp9cUsno
72utSjijxDzp9fmpU8YgRPu8NGo9py/zv6Ij2ZXAYoZh57HAZLmuS+HjnlSZAXBR
TOP9cBAOj0onFDGoGpreJye87hRVK2mZJnx0bDDNbb3IAQoYxATkmmt+w7rwqbTX
E6fcos+jEVtB85Kr0/c5sfh4NmXhGzeslvLumElL5FDDkXFWKAil4FxSn5zG/8vj
zDkmxxE+GvEvuo6cC+yzZXR7aD7cYClXmJWUH2KohC+euz8X2Zu5V8dbcyhU4Y1s
RnWEdGuqBt6CMvd1yIQ7S6mkwVfBwykKkbVnoKge1JerTFu1rqbeOHY2auf23GUd
tlwZ/Q8Gmkn9nLFn3yaelMtOvhl122z9cRtoJKfIpdxaoKTU+r0GuqzsEXG3lL1H
dsW5a7pWTZa1CO3gxngbXpinVsjt5UZwUx4/K8GHSBhJMiNUw18I9P+40t/S8L0p
Jm6RhqQagn99Mxf2sresaw==
`protect END_PROTECTED
