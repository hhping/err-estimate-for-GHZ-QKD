`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4FoFCvZpgv9ZcWI/y30qg7zZPyfxm7mJNL6nZkSAP/aKo43GKT4iJ9lNGBlMR99
RBzCdjvg0mbB2/WlmCRN4SFT+l7WGTSqXUdhPiVeTs07yB9LsnKmYP7QxjoKeGsv
N1rIvUvQ10hVEeSqjJ56js/bS8A0r4wRQB0jn8SWN5ABdtFn4VSBDLXwIlyOcjk1
q78iX1IP5SxDriKhgClaWGLRLkq24u3wZVKufXO2LBe7H0IFWH6/LxVDtm2p1nvm
dH6g6R6ZU2rQy2dMv8fW4ytWI1am4u+/msytBMyxolF82WOd9EP4bChp1RT/8dp+
mRWPD8/V2V5abFBU+CngIpR4m5I//ttOWsk+fx20v0+TbBN0Vg78gF4G9PYMhkRc
HC8XwjzWnVKi9t8HWBH7U0HBzFWxacKnCXKdyw/kz9uAVAO3+uxXD/ukRVYETBVD
CrSM5VPbSqs4Xa+3eWYOWBaTUxY5Y0mAFFF6HUIlrI/yVJZiHw783SZnBkXfJxVv
ROCqrJCvTyqFP7s7LBw5VQ/J2KBPGVSzUY13EjxDloUi1fiDcjHaZFj83e/A757i
yo298fLH1zN0bop2VlmCZqffA3XsfloCNjz+LlydMIPsrg7gu65ZX5xlPHkjWNFd
xdBwmq9wOg+C3d4Tyh415tJLNtN58v5Io065/aV70pkxoLimhowGhm3kLUYbXZL0
V9M/3CiXZzt5nhkAq4xQHGH0Rra5gUINpSJVhAyj+TFjyj2aqbYsFhS+OFzwVVKB
XeTO1l3vnMcZmxfdkfuBwul+SX7uedmzFIRYDDcKDFQ2NoD7dZ0fnVtdRmg2TNET
JtEWm2KoYNpIrxKFgoD6hPSp9RKHXp5vCZEY6MGcOaDtXW7Q2LRJ+WuHDSJxvgkh
pfVXARcDOMzGkJNHe4D85qCxqOdRplp42P/1fbQcDWku0XN+4Mb78QAZKdQZTqVd
bStbxDXt5cTmf9TwFOa+Zw9F9UklifSutRKGvGNMBXFi0vKAolA/NVBx6+E7i7yo
w3o7DCVgz2Y6YgvVplqedVJ+av/8pi2Ew+/DN+ghgQOefhiaHpoTXGJ6GyQ1zfEO
hDZiuU7qNsgyITWglzebZ+puQM5W8rakaG1EvRv0rKApWL2B7d4Cfi+XYWdXgDcr
wIVrsDhPUm9GFKvfLS+CuKQJ+GQBR98v9hDzFgAWqt0LcAcSBzV9dW1+hs9tUVUN
eG4X3m+KxRvC0M2/jE9UP8Y5fLto1g7qzg6Acgxav8+5ENXOfykzFGl/ot3WG7i9
hABuopR0YNoI8lvak5ch+7cy7mY3cEmZ43Kf73ZYPGH3ckFnyx95ruh2/wMjIh4J
YwekKB3+ys/1oNuQmbyeFN7Z2oSJzTtShrwJ0WCh9RRqpBhkJUK5maUpIdLkVLmL
eRSAcu3cW8/Adb4nrmYutvA7gM31ouJOk+MCGKM80+xd2X1w0f3kxVGJ08ms9Ars
08DP3F4wb0p5lvchIgFHFByt+4hPBMdaxpmv3sgbWT92EwCnPFq2EZdKH2JqzTFE
zpjLFHzUHc8Xw/UivxpW5qsWeY+jmMzbtHPUm3MCY7WTWQM16nqdYuRiz8UKyEGX
bCUaAFv471dqVl5i2XUItTap2I6d5XF2AeGhDiRAM+uHkQwpfYaclkPBiFMTHqoJ
JJu8nlPgdFSb9wT7elATp5lU20/HpTJlqFWHNuYkV89QiH+jkr21sc+WgnvUwg9C
ObdgJ/ey2uZpkYwTqtVOv17YFbKM3Oodl7K0h2lsQe+fqZHIFo7TnhpWXdXd7Wdg
y4GN+YGQvDdexoCvK9qEJSpAEP9WuDH8ryFl57e/iPjUtktLVjnjdYFGDR6LPlmi
UVvhCouKwcLJAb9WHnvFK499s0/c8N1y2RyE23zXAjE+K8wujlZdh8IPVMDzDimA
87fKmxa7wmC2pVO3gjnCWIICGRl5+WOHHfbyzV+PHVmOHnL3Gk1jBfcKVBpTrjdX
t2jz2j842Q/WXkKVFcCXRVk5y2gLJ+PP75bV49s9MNb7uVk8EUdVADyejhTJS4KP
ntgvmQdk918wLgTLvR5/ZWZlsstL4zAjesPhu/V3UMa9ebdTfF0n4k+9itV6P9MV
Mn4rq/bYtIN+I/J/5qwaByyfeghBrQuSWuGxee+i9gQ6CSvG319VOT8HBCsq3tsL
AKeEVQAXe9TeuveXfcEmntk1iXh79PrrbtL6f26kLfa0tL5dSbJ8kCBaIpKPrSjB
+U6+ksfh4u1k20EgVzIyaJ1enz0K+nLkkEgVKIjfJIGfsseaCSbAfl/ohkeBZOFH
oRrhNvhAc+Us7E4kXYpQdXHkrc8ypmfC4onOpWhu0DSe4oEjMhDjandSdazERwi1
K+db2c39XSpm8RvbAXqHloTJKXAiJbtf8K25wfnT8vxyseqn+AuCXqn3OVy1z4CL
YLX6AM5Kf0o2ubm5dqFE9TVhExEA6Qj6fwHBhPPxQsV09emp3ZtSvMlsjRHIOrdX
XQTvlUEQtJFPLz7ZqU3IhG1T06wr1anpvbcOktwdBFtlbHoe6LyU2MjajjhR0FI8
wzOdSP5DU8sqy0xv1WsLpBCWDL/V/5OmrAqatc4i8Lswp3ECzzhPHnOYH+H5/gE4
kEcjyxDqdMKGvJDojiUaByD9V+aJXAfh1LEPPY7M/EMpW0W1JWJ5cEDx4n3/DUQh
ku2FZJS4XGV5qACO7JtRnGcBoR5Y90NiCY9cl4uoY9CqGYdREEfFHR+caJHVJNIp
e+NBp/Hcv67hiJ1wSjrsu7VYLMaf6H6tToE3NiJI3xNTnBjwtSC3Kr5N2xaq3Q9/
C+xk5EiXaqzzOUUAPcOB1D2GeC+F3UupPRnhcai/N7gnJIwVS78AUf/KlEq/vHiX
+ClIcHUFvYHRx9/KOvaK3D19fRe3h9cKjLJd3fE6kuI7k8swXKcZfA8WnJe+lscU
mEzw4c6ZFuUeKRjpOSUDbt8GvrvVq+rhR+Yc2DkZu3nPks29gDkp21VdzMn7C+C5
n258A3nxq8sT0YCEG79yAwBpahvKey3DstGdD0IoFz/XcJBNKX/1m3h/1HZRmKHu
NZ7u1k/BgMqR4tk4eM8INvG7rhYSpKcEMqJ503yehT6LF/UeCtzvYY5nfwJHXsL3
xn49tkFdtj1YmSKCP5GTR04sPRZOmjU8f1jZxUToBb+JSOa5tMlZez5fFdWcNPRN
izP0H4fk6u2LLk24dhdaIKNlWcCeA+XGi2qj96Bv8rj7WchDSrestvpoRqI2/5in
4/76c8xbSlLwro9yEehBfKBWRfq19XNCF3CxVtHx3CeSNBTrcrLT1XjDEqayN145
R6YsJwaS7w9dF5/0QckOB1lk01N81R5kWsSHhqqRvd1rT5KcnnB6urfrsMKsXnDd
HdwGVY/Ml7hi68awqb4bZArVm4IqN3cST070rCvbNcuVo0XUh5i6aMW+9U1zHzMn
w8tIpCf+poaBMbUprmUDR96aSJCmJM+H1Tds8PisU8EFNCB0kfdW2d1DGF1N6Occ
CoIONPRbALafBVL3EAQueQPRPPBtmmKhw/bzGXk1LOgakpC51/djNfeNrVsUADpo
ryT7KETc0flU1Nf5zS0pJA+OzFILJSXdROKzHANsQ/rlTwTiUIVPpMsW6tISCSjj
G5QGHGLtUVuO2LfTznCyc0a1F9tPKq/cU06V0Blbb6QC9HbFyOBIbXINWQ2MyFab
OVLxFlTgWisiYD839VkkYURzRwQbZ93N2E9yhDsq1RwE71VW7Cx+9+zDfQJi3nFp
yQwNfa+ytAipRcBwwJQlwB9uMawvrClfby3Hae9Kv3RKeE+IpTqxbGkaKB+o3yeP
4mzQYJRbrYp70RUwR3/G3KJjKUYJuapMam4l5GWCWqqdRkPY0hAcGcM/iNmh8gkI
xC93F4MiK1qZwMzCCLZQLViOgcuWNczPsqHDykxHiD/EUuVLl8mZre0HIznPuQzq
1glwMW6kDXIopBQGwaLjs0tIg1x30t7oy7lMLklfYioXd8H0CKHLo1ksdVql0ltO
HP0qJ3ZhmbhwJFHtdARh/n1/A/EDPfxfIKjF7483xJtqbqwbMKpDf422YOfQvIuf
vpndkZTZLMZwkrBe9EvGTzLVE6lSf3sFzeQwzzmmcczWbhjhT3DX4/+DnfUmfrKz
Khl0J/BMyM15+u8+Nb2LbEcYGE+6XVYh9IguLcKX0//ruUmfo8nUxeckTjCAFJ2j
hc1ygGoUYVlvPZOylfh45sAahLRfu8af3sDMlzANb3ZdYVrSkxaSLh8essexiVzn
65xbp0eI/LO7kziGBCaDZOTrasoKOc72uz3b9IOz4g6U+68Wb3O9Og9bYUYk1SlU
8nNT4kCdNlNh2tq7/49tO6EVx0h8okGjBEjNbiZ4n+x2eMy/c+l1JK/hxxOGU6ud
fyXeqUjJxBhWvuF5liXYeKWpz6DKdwfJkq/Yl9YstPkaRgr75zM/DiyBElfR1WIr
gNLeUEQtQfzwKEYSEkLv77LGqXdeo5/pZ/tgt6g+4rQtt36ftVoSn6EF+V8HDB7U
8LAdoNL17ajRZ0pXGJbZFS0oWsaiaAdXRlEKPdOPZcmDgU6F8mRgurq+tb6IsD+q
`protect END_PROTECTED
