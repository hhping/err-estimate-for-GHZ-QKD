`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMMWVThvbmLM+zVIBmiJOwtxmthcrnYD6+nBbEYORm+n8vesFdv4nJ/PSkigc01m
qrbzILi01omDkYnXVP2SconRI9LZng7sGUtBfJDJVJxhKmJ0Eo5dsQc6iMZgZnx+
qar4TD84G9wuRrVJJsd0Xh3WjgUaW122wztfztdhE6rZ9EhcKMSDsEn5KUrkCwX6
DpAhe9mf54/dyUzEF0l8tLZLfpftWIzXdOrNL4imPJDVBe4GJNmFShfyyZjmdzqx
2k0xi3Z3RoTnVTBponXhjYGRBK3Ld4Pr+fxwALL046QCr1ojUac9SueTRw6eQfBx
lcFQFcGaTtmhWEiMbG5I+92S83DJRDUcKO/HdONF6jsAeOyz8R9uqFcnZ71BAKVf
zA909qfim78qd3cUR9i4V68nq6GbFtv1Kpoh5QaSQVecmeTBXG7bODFpCSdF5W4C
V+26ruefhoID2MG2l6u/5KWXb+dEMRjX9K5D71EM8l6O1SqNnPYbYQyoLvPgpgBP
X6r0ai/3+Je2PQBrpOMy4HcZeQRDKGUuJR3mqKK8sd9ak5pcmDTbtXu6LjmVfSAB
3sicIQF8ibv0aJdfjRHs9XIDtuaMEPBnnXaFNjxkhl0/GnphPSoiaNez1RKiwOlh
yinjlIrJSAU2aiG5S9asBf9G10FMBuOfDlY+607W3d9OpVv6dIcTpjp22BB8oeAZ
pfSmqQrOMYxaq8gF+dy2ZydprkvPbK48pKc6xiI9Fjlb3IantNMXoR2GWW49GTrC
9759DCpItBhZgRfE0ZVvK4SsvP5ooO6sVMvySw0Vf3EfXyjX/LgE6r05Xzqot1JN
L+Qp+0DRkLoXt7PAgAVQNwFRnuyO8axiiZmwDGvKdkArYmiF6UqdnzcxdbimQUob
VTQ/F9GtqIgH/POl18RDUw==
`protect END_PROTECTED
