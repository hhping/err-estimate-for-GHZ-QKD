`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W25QJIj+nGQkUwA61TKgkWIS652euNArZu6q1DsCUw1ANCfqhlWp1n+Ks/CVKMiC
qFmWbdUFjyCuzimDbo4psbepjKiQijeUrQBnsC1DHaMvxq5MNzMXn8KM/6jAZbY3
8f8cVJUeEZzu1XAa0qI6mw59d3i2JOuItEc5U804rfxy4w0mVSP4mV4VmUPte/2K
4moYRkmycFAsDaAKhnlXQxGyrV7Wxk1FXtFI8B9C/TNWlga4V17RZILCxMTnReqa
mKiAKBXERMPMye2WML1pSe7+jKYdGAAwuPhUDhwuz0o9wUdolW+XghJuMBPV+Wc9
L4SeKdm3uLUmzjalLTIboFEDL99StRWRs6gauYxwwldHo5XRZXx9KA3H4b7IxA82
bQ3rt+d+xrEpleV7oVUJ4WbS4CTqw6GGc5temHf+vJ4BH6xTOiXdkXjT680/SlNs
1S9oRV6yscfe6O1ayEE19Mrjz17s8BfyGTFrBM4BoYxuS+qXqPE0Usv9tn6CQ5s5
khXaDxCMHY1amQzMBwRCN/up5uoJzYAhTMhTpwqflUKH9fzWy5LJ6cv3I9Tsxtjr
1MeODPhrYfFPWYCPOk9EpKoKB4+l2WFlS1BVKyyDPj2YE+PdgJvkG9O7GZCylxOZ
kaebjwRbEujo/TltbdGqBQHteSYwi2cqxnQqJIoh2uKjZqdvfSdFWV3ztMo2HkTV
ukERt9DH6bIiCuOksIZcOx1XIpt7+2bfRkQGw3gAIiKJ/u1PouSuTbEfxeaipw8f
pcN9k/3s3XXlzkaO7KepNviA2pr6xEhlfVT8fYyHkjblP+4hHd3+mFSrW37lkQpe
nbUTJ7xzXyj1NNRBUpZXfCMUHkVjBky+LtcKV/yai2qJc0KIUaC2OOP0Mo2tKBQz
KCQxn5797nfPWpEmQ4Sz8zF9O9YM/T5+ZiUUKuGStKjpCSKk9UI3v4wCPk/n3dPL
cBXlbyKsKkRultc7maoa2VPWlg5bJZvrxtDr0COLozfSnTeHcH2vs5gA/DavxfQV
UtnKqya2KWhaj1mkAfEKqWgONXMKqLb/k/n50Aw4x9FDsF3MHz7O+RNGvgCxI9ca
9fkZCnhvSHkLQcDHjzGA7anP7I0CommG/2FRgniURKcT3X4riiRbiWSCaWog5lOK
V4yROJYa18GyuBuIbNAN2QQ6xoZFV82bdQq73nkp1beEVJ1J85sYhvb9n3Zrw572
JkwrkBtH+IAMX+aRo/+iiRM77glivIopJQwNJrCOsbM5ZSfxHCvmRfUFQWh5qgxo
mxrXUwJ67o9wjyvgZqq3sige+v2+jCTbqQV5xQOVqIUYjkhgY25QC9ZKZYs3V73V
gb1qMWSp7XVxhIuRQyjyK+Sd1CaYxMOXZ583PgDcbXjrrcfEeOmlR3XKJTeCA5pb
93ukFTrhzZTYMgKkuR6gkV+qqqGdlq/cHL0lir7qAnjgeZY+sABe8HRUC20IwBCp
5Wy42Rk0/SettJmclgq4rdlatkUrpFn46hAgRR22rkXDFWDX/RghGajXBDf0jQxP
mUzcYCDexa13KQBTVZrJWnmJCgbhQU9mx4G1FOQkeDksDIhW7e7cqA5CrKB07D3h
piPWtBU6hGyylv2bNFFXsZrNnNDeMDJvA5P9158JFaWxW1kWXmEEVaxx1SFN7TmH
36qOUYJQwStGX0Tw9KWiHYQ07bIHI9v2O2BNqrh8Qd/2/lyWan2/kS2riWHrWyAJ
U10f1dTJo2x6ARGPgpD02H+OMkJZ4z1I24HfRarYmP0=
`protect END_PROTECTED
