`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcyQ+b5zlj8eeotaYZ6tyUtecRm4m07CcqlTIQG3zm5ZFQSbGCyop01Ewsns0Fcf
kaw2H5Fp3UscUuVBC3eH5qXxzzZBYm6EuB7iTFs0l0CPAiCn8vRxCNaoHsE33Emz
W8l4BD+rQMgtd8fUCXucIGhoUcD7TZSju5wCo69LXOXTW+/MEkoylf35ChUrF48p
UD+UYYd8LzXyRCeW3KZgKha3Cz6XquJ+PmmY0jhOFyo6ujQcbk3c1w1QccE7xCE7
WDGdHlsCy6cL+0ssAudo+2wnDrDt4Ngy3R6XDZ+iMJJ1AgYnwr5jupq9SWy0dVTa
HN/TFtDS0k/QNQe7YW9uSPHFvwycJEZDx8ygm8Qulqo9mqCtHbHF6yMstQQsRNaE
NIEpp+7HG8MF04/2pTc3c/AjJ6B3ftxMnv/VWK6Kl/xyg9ra5o97smsFo4TuVrvl
jH49nszqtwBWMQ4l58nq0dpGYscnMDn7sl39Cuzy07cVxdwQTzitBksJXq+Pz06S
YToV9IA8XFfSQUZmNx1bVV/0MGjdETbBnEUcZKdgpiFGUm+l/vhlbYV5Fpcyrt6v
RVGfBghnh/VcbPLg7+bKlxF/zu/IyKnJGMeLfpNbBuUzzsd/3oA1Cc+pkO+b1zYS
QyCkjHNigIiqK0N49hi6vWpvZRasHSVkxcEMYXcuupA=
`protect END_PROTECTED
