`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36HXxXhjrm9ct7Erb0CEi14madl+9fINDtHTXH42VA27cfc5bf9XFVcDtO6myOUy
u6Y4/JvlIYi30GXNYNEiTv1NCGHKvDhGvDqtzVM4sgutHGLt0TZtcdfqrylWWWVw
PBxW5/aVrko399/6EwvtxtIgXvqE1/So8fLQcCIvnQsQtK1n4zY2mkVwpcHaOmCC
zjrJYEcCosbw/o1r4o9s/9ae3a7dg8nG9wVQ1Tp0fmP5HgtD1gP0gk3Fhv/TBgrG
IMVOmlAAaYXi7wp/yeNNMmHEPhMP/1EwGiQF2GtImTzCdr30T96kMqE5nqLD+IXh
rcO3BWuykiQexoKCAM/LNezZkmmotyJ6tW8IPhd5MzUXpyrTAlpyaWqzyeUno+ci
19E3ZgYcKn98XXsgxgSd8A==
`protect END_PROTECTED
