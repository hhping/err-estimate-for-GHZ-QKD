`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52nwviloKJQf/T7lVBmCxw4ulOb1xmqA5KuKiE4g4LijFnuNX0+GHd4mMN17FDSt
APO5LgbCzYkVcRcy99jOvGBh7W0jAoXFOH8BVE/46mklG6FG+aKofrz8dIV5fnxW
HKeZO98WPI+UsxxShMFZIq1Wyl1Bp8Beac0LqtY+S0ltazvAFK5Q45mEpNSBTw3Y
enztp0VTYSRiXv+juNUFPYomYbp3dyhF6whNElQkSmZBPrePaSAwC/PJowlu7MuK
tEgnMam4vN3QTRWL8bPA3New2RGgqnYrmzU4yHgJ+rcsCwtPG3M+Z4XK+0x2Uki/
UvT7Ut+Cmul/RYhfg1DgcSg7+8cgT2jLZS9W4It3h0G6D0BkWaUSMw3NJTXp/HD5
iZV/0tigCuXDI5yDcQpAu0eN9VHXsHa3rK2OjtPJs5m/IqZcvMRWyczSX8rLcGjz
vxNc6ePAEHfQecBvfv9F7QPIXXq7Ao1wP/C4kKURClXCecVbIgusalLDwp1/+qHY
GOmvE4nWP7AD/BQQ7XRbZWamvcptdcjfbqL07+mL8oyCtnm43K1Nv5wOFtuFwwuy
5ySAAoEj51iclDF7I3Lfn4Q/QnqsxRLjCBstIk9QJyxVV8rVFplWQ2BHECMEDehr
zqS0QjvpHtplvZlUENFwN9kL/Mrb6JYjoyaxvkASyzs=
`protect END_PROTECTED
