`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
77QQtRyfrz9sihf/ck2fzj52PiNlrTq2bKCP//Mk1hSGfPyz6S7rquAF0/1SIzzp
2qYao0cnU5m8usW41EB/hlp5p7qdxPl5xTXHTIIgImXGAcmJaYCIzKFa5D/6JlGH
0f6lID9zPJcE39rqdmxF4tHpuT53dDSMQRp/zBAQNPLEInB7DWxMIRP9MO9yBNyY
85AD/ltX7M6LaznBgv3lAkmv0G3N3i3Alpc+dJQ3gjvbpwdjv5ttHYU/TTjQeNy1
Kd6iaREN9VsMzTMkPVVtlqznPxP/It13+sCR4MO4aXEKW7q/JGBzQICQQTXQ9nbB
2SHYwKPgYvW0H3NAQq1NAV0kTEgw68aFtgxBMJ2jhsDI6Eq5h565BI7VbcogvfUP
OeM91I6vvevsvxxjmir2CXJJE3qpP++H1I561RJhR87eX3gy8Q5WDXjNrBXGSAhx
CJQkUeHlZdISI0VbtHhenEjBVYyupUau8wue0dtCLtpRxJrkDkSV4MeApE3QRufm
P7EQkgFcmtmxVxSQPohOOx/H2f620otw1gALa9sQuxAE9V5SKiDO8o46sqaogM1C
q/MpToBzX3zyiczhz+4gFspxdoe3X+77yE0AIziwuz8f6C913E3UseAwM57bZrqa
9vpXM+/YGdr3zLvmJsQx/w==
`protect END_PROTECTED
