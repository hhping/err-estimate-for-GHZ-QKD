`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ES4ukIQFKzgOFfOFJT4oJ9ql3gjZArIorY0MD+efISJH1IUkntdfPy2qPM0xLSpt
2Wg/FQNi8rSNIB8NEhTs0iGjPqTkWfdVoVjiSQyK33gKVUTqHW4KJHngAMCd7adl
I8VSJN660zPWxVUfRnue7MjH5mxZY/89T1KjarLkrDEHpgknd1U/BOMI7YM/HZPC
5Y/oP80Mw55GK/sWemMn7FGa1CTuPeEm3TtiJLzgSTO4aLNJ8Y+Ui2eEc0AEPkEj
nk4GcBn7sRMrkopxeL5FVxNDmgUbdXcXDtEpGerO8N6Wvi0ksfIlY/cJzn9ZlXNK
zFtFqLG89IR1YPOigVdkboR0ZgiR6avTzQwzrVzIbzrUgimLRu3aoOTrNc7ix+jo
ud/Scvu6uWpWc2kpViFmbbIFNaOioEarIPG2ICyICLXYoYD/M6DITY4K3hTl2DNy
oD52Th8xjUAIWiavSgNNFLs45ta77a6ViexWR2DfTIixsJvVivaj0NmwhN5EX6sx
M6hldqyQYF0veAJLmYF2GTYPmUfcmYt4TJJXMtVr7tqlL1kVWP/ZNkG8CJKcY8/B
a2rwSmdCIoZryb1OBx6k9KbpxmMioHlOyv3+lkbDeCdJK9bc9+sAYeyHb9jTlm8s
Rbj8nDZuIgr+ZRhjYr0IblYoumquVFluK0clsW7vHvny26ARy8M+SWu+ukTXXTOi
mrx5u4D70ykB9My9lVIMevDv3k3wZovu4Kckb3V3wWHhiWSX56xtmn4s/8veE8Xn
iruSZBwL1b4dRI9680b6wAsK5lvMvew1hUQCk3iFNgye/zwcqEPzH/8TExDHx1ED
N6b3/pje8Js4GS87QS9Ii49OLLvt8nmrQUC2lx0Xace571lKMHcYk60g1JFPryGW
IpOz8Zlw0rZhvjJtzYE/VZWqiOqgbMaGt6nC46QHKM2iJxEpwrs/HmUlI9rGHKk/
OY++KemmTLWx0e84m9NhYj/7idKRfddcPP2k/02DDKRjEPRk6EyW+iz9GIJ6noyr
i2cYOKq+XdlhU2SmM/046A5Vurts+/KuNfoRP4uEri9+2/WhhTGpLIhvWKedAbB2
YXpQju/PJ6S3tHRu1iWWfVMvqB4BE30I6mHgyvSQpDsd4dQ8ITkQiNQaahV7Vl0m
AT8T6zaufj1TX7BASeegZNHNozOXUnOF2QMlEDVYDl5rhkQeCUgMp0jXAo/byADi
NB+bpr+NrAsF0rNGmRwJIHgG5fz+wNXCWs98csA1EAqk1YM9+zUJayegAGhXWkIS
cOPAkuKSW10J8Hkv13rBmsBoJRxmbRbdoaYFXlEMcr1ea/8HBgJrZN8lVe7iaEYN
baLczdMf0pdnkKaPi4zxcaf8GnVea8cdv+LKALfVdEC4LAWr5X2wWmHLQvxonCNd
3j7MzONNss/l852XQEm4hmNsYrBFqASbVNGNUMnHjYRD88bfZNiihXKkZ7Og9CW7
c3b7cSq4A5f3ZL+rffsfXg0KXl+XFaVezZsjGMVvORUQNV1FhlYWqS+JPu86RQgS
LZAZaeTADJfN7Fdzqpxnb//zurRriI0sra5/O+E3Zd2CUnfEToup6p9ambqZcUDI
Lm55AinZFE4Ywhzr5r4RA/d8baInF24yWbL66NTYh9/aCSnTQ7bBT//36esd1bLZ
5OaabrNkpRuMZzekSsy5UsWI/hljIoGwojPWmlLKZNRB6QdRt3pmy2UYnVJHukOM
g6chNOS+fMj8OTZN69/PjzRgpTKHr+9VrWbZv7CQBqelwspHmbbv3PB60S6Jc5DX
XmUpOh8sLdJnM6RjNIcQz2GNn+qu5VBliPFd52JJqrAn7VKzq9Pa0T5YRaqsiEun
LsE4HrucdY+9Os9SeiG7hvTIiAM0hQ5RkYjUis3PW71X3Aqd2g3/btgq4jQIhAu1
gs+2zdrUXa0O6V+FQwWq67mz7CbOId84aj5Q+Lvh1q2zx32a0UJEDALT27kDwbpE
ijMezFA48KLJxe0g3lYn6oKCNEfh6ItlgU0/1xDoc/POphI3JQ+eKqe/8NyPzPLg
svw8ZSXNInpfVcou5JwHeOnt+jxrp8k43Q6c9rmdizr55vg9HrM3nVOUlhKmHslq
OsVLsYN5o+XcACQDfyQg41/9G4oY/sMGkhgoPZ3lryMnmcjbeOg5sTsHBa/gnavJ
8N45GPrTHjGKNXjp13Ofz+F4MdXOJpYXgJZs2BKm7vBcxYv/DNY76D5noYNYVZCx
GNdZOlr03/n+SjjOsTyMdLIsQp/zLM8RM4+Z8NUqOtSN3lzH46xeGywUMRXJQsBj
inZ0jAd1qUveA9CiKqVZWQ==
`protect END_PROTECTED
