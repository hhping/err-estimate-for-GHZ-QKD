`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5n633/bR4ajApIfurVvune42LOdrqOaKUkmBQF8CubjqpEzPYfQEXEXRaPnVSxLi
jWmhcqF2SGBJdeO+0Ex9xNfwn/uDQjDnFy6il05ZxDfdoDgSN4N5eEpxJXpYpLWe
tdtkkGflFvV/D/MVo2LQjgEjauc3HJm1DZeaNkqJDCN4umoi7fbeHoU+3P/lJFBr
5AnykRtI8gDuU/tqGQIKUPCOdnGU/hHY6F/g59ok8oRrczds7kO2JdMOg6Ympq6t
/m7bWob5W1Wfn26JFuT4j+et/8BB28nvgo7RMZUQZoFPGSAzfwI6wvjWy4gaFAIB
HPohXpTlzXrl+JLYKqnv+m6/oyGwSI4LUvl6WIhGqiTjLI14iJQkfciO7LrvUoIR
f9RcH2TYM7Gyp5ZsgxgN8R0FNUpWPHQ4i6cXmhpjWu4rJ7EPEd3B69QqkvGoUcyx
WhscSX734dCI1GNjcgx+z3OxaNZR99J47iNAfuTwjYEiE9wfOTSGCPvlZ5SuB7bu
sxxgufgWwfFds1XgzpoHHGDMqLiThD4yaLhYR4IUrL4hhXrL2RhRzuT/caLw/0Ew
PNd9af+Lntq3Xv1IvKEz/eAvhnkU6873d5wPW/1XrGbAEi8i43bVhEhhc22vKRNB
4aQhaZDPXcWyZvAkKXTAQmt2P4j8ShpSYkqkvCwJDJCY0fLrw2Tx2Czl2PVaEIi6
3ecjPye6L5qtB5EcMCPQ5Wj7rIM1m7bM2v/WXrieUd5opOTxCLstYBodRXbqGMrk
/83VaGom2udjB/15pBLXhjwzB7qIcxI5AoeJt60sAbjBhdFnnCk4d/QUbdHguR0J
Q0gYeTdDye1OhmxiTSbBFcMQv98u9Sv9lX/i9qxO2VRYU/1awmYrStDmsY6ncVj3
FP5k6OYMaj2hluX6GK1gU3Wmw/V0uqBXeQOC8G8szy3tMP15GeAi9l+2JgNJ7zMC
7dPRBBfGhJ2cGyZmfjmyRwotKn03R7udthtVCJuOr8kvcSF/0ua5qBlnmGKZh0qv
CPQN+a6l9vK4gZrEzCtlsa2ta530Ik2QR/Xo7+SrpLogz5CXKUMJDFGPOquo6/AX
/rwwqVm0v9vFmDddzgPEaCyzhc8JzFAP8ufY6Z9+wUJl9iR4UMqlyfuJz+8Q15lz
jNz3Nv7WBDOLdwEE575Kjwze/ZsEPbJ3oEFCW8l8zxGyOBuCPWRenATdQV0Zct2i
`protect END_PROTECTED
