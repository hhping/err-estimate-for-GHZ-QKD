`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFkC6+P1Rsf4xfLVFg9PVpmquSgHFK63YP6+mCEjb0rmUl2KHSJTLGjrGRFesHE3
y55Dts2DXNmNCOI+14KajI3Q7w+Eujp9WufK4xXsbtFoVYsavAIsi6RJw5G1NvvW
a9FJjsJoip5rvi7o9LQybr+shiq5ll2g/Yvwng513NKg1WOBepBBmzzFQx38EmTZ
pU2LcEkRCKBJqrAfhElZga+L6JW2RTrxrcI+DM5IuXrd9H6nSI+SScDvJm+xXkzo
PRflIAs/Xsk0l4s82yDokrnmRR3BFKf2hPj9c9kJ1McaSN9R+9EU8HbeIyDfKj8I
p09EYKQWpqErlMeyyyjqtVfD6ctsFNTGvFckGRYi4t5L3deAQpLWLXJdDXt65y1F
4ciAKMUSRjnielwBV7T8Pu7H4yp5XruZWP/GYP9SOKrqjrroOMDQqNSRYIUYqBk7
fg3Q3vNLkrLmAdFCmF2UTWdF62zQdBzYIPaeF3U6u2cHMNM0mQrm5+SxcCe4b6Ol
z0cKEellOO3NFD3fZLO+fzbqJfgaODNB3DZY4kNM0wkE8+GQjGi/n3In0oar4k3V
Dl8xBVWJTWU+uBKEukoh/o2KbXGWA1cRKDfUU1T4NfBHYoB8jAm3V3Ehl+a8RigL
5eiKigoPhb9qlS7Ss4GSDbi4c+kyzLBgfALTi0pkgGh/KryxRUFs3yZ89xRtKwKh
MtLIdyuhhfLV8hMZ1pQmXqVeqte2Kp/fC6p5XyaMS1aBsv71nAAf10zyB5C9rQh9
PYe287DCTRBtu6bJOF9fHagnz2OAGUkIw6/yjQz9GAp9MhfCFEmzLUVr4MjLDenP
bApAAr1UACHPjCfu4/rcvg==
`protect END_PROTECTED
