`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F+RG/5UP6P+sCFY0wAux/U/gljeYgSYxmXeFJrL6uYPXrQaRZk2+bYVrRE6VT9Yp
r2RBNoxHfm+MunhbQAU0Q3gp/AQqYxK6BHpHb9pUS3QGhfxraCbD9ZJC4sYlMKEI
BG/AkOrqqwZeZK+Ud/bgfRWiT6kJL9b3+G57r758RKI=
`protect END_PROTECTED
