`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4Fv0y/wvke0azuVsBVPrY591QhlQZDDIaANwLvQWYKEFJJlIQjlhi3XGdCoMavm
nZDwB5kPVVzYn0xq868V47mRYNAnfeo2kX6zj98XmMAJ9yrcTJBNWf1drhxuYkAb
yOFYyCCuvkR5tmSRD1jhrsIcJRpgOnXOMAVa0Ib0skLGHlWN7h0eQCOxqA9ooro6
V8WyV6aLm8Nt2DCuE8XUD8o9fEr8Dnwvp/vGZkw9Pi4eBgK7ls1OCX4UHJkUIHXT
zgJDchNEwmWAoceBs9LET6fxJoJIb3bMmz12026XVWpDlh+6cCF05QEbjtcq1Yi/
GxjCGR2K/6xvSUR6lsOiGM48Hju41dOA9a6xJlZ424jWShZHXxCg2pWgy+dhYjzk
hgvTCCTkNC2P6DaWysl8cNhp5+tLv2EiORN4HAzeRg/EKBF9jnM3ArpER9Rv1dlH
YBaVhGPay8+n2nZjN/UMK9hAQKFyBVkITu5KuISJdwaGJ8yZRj4cbaNS3qj260iJ
ubP6KhB9yv8y/zrQqvxoDbm7e9IsJX9EL23sg3gyflHEB4nmHFLxG1LiNCVnvA1k
250X8HQ3m7tLHkQFerv352gRsKoBSeSqBX5j+dwRord+h7+WwCwoAy0xUAya4OzY
EhHwgjxuoeQBUJTYwkZDcteA5SsyIdEMoCxRpcXCq5czOd/So2e1iBnq5YO9v5vp
5+9ACdC6V+QXH/7AFL9Ui/nyxHf74y+uzD2BqFewxQNl9QM1qeGnJs+17HxuGG0G
Iu6CEe5lTKp/eufwqB/VALF1a9Ch7nQWvWwLpmzDdDMY+SBydWIVJUCXRTtHNNl8
6TQAWydJ2ijWDvlM0CGdncd+Ew8YVPQnuur+BuGnqrjxwGnBYBErv7EitE1p0bZ0
EYHsuwevDZgPAlFlK8JCl5cjc1GGZKbnuq8vsTKH87sp/eRwLC2lxcAAeq9I/UVY
97uhZ/eV0WvTs7gdv3KDyfOAu6bU7ObwYhWtR/ETxGJUkh6wwgDcSfjNtNt+H8c3
WUqv0lAaHRfxn5sj4KfDhudkaUsnLVUPb0XVsFBbscyqnt+7K+U1TF2AZ+OQ1IXp
RFxXf6HNPsejePvYC9F6DhpdfP/qgFBMe0XZdEju7l2QDjO63C9YVoJHbdT83ivI
F9mV7wbtmU3sTeRAj6AhLeYMQqqaw5NCJPW/hAn3h04r7d70Qa0WCnyBHcwbd6lr
7/+4tIJn1eJuz2kNdT8X6WHzEKXEvXS5Ay68jofQS8iOQ9gkIbatZZLxY+K++Y8r
xMcue2qLdlZcd9Ban2Rvbs8kWvkaaVU4iOcBmawmutTvcdkR91AA6LYlmIWOSEII
6u8Bydf27Rmk9SgHvZbF1B5qct3tjmM2jAm+OV/B1S4qg8j8hIRzpafr1xVp2iGy
53dpYCgU3PhQcHrkieLWUh2NZSm7b4dLClob3EA+l2ivlVEngaSne4ncQfsGFs6n
pSGUAhGxvR0f7v02P5tdXAlOAJJscd7HnRpgBEjld2cktoEOiThNLZj5ZhnpSmB8
fihMe+lz/7epxdvIo3iEgSNmIr89iJt45yo0tzWJ+unUy11e9V0rRgxHh92+pjSY
LQzzHQpI+dYZ2Ltu3LxkbiyIADGp4AULbGI7hzthRG4H2hXRWD8tTuE0DpL0kI+q
bpMiVXoIxtvo3GJXTWgXQLQkAHXWPzrQ4CZoiYgORLAQ+4+GQwPssOeRXfvPSFyX
u+xZ6PzqKGy9TQ4hjuv8R2HKUgBaXJYiS4rk7SssZSG/KSK20EoB6to7Pt74F/Ve
PDQ3dnwJW+qz4/mhmsYTcOtjeCmluzIoyInA4OkDERBDIlToMSNBGJOsV1AFmbH9
KkZCQo/sZ5Gdytb/A9blBPHASy5ZZx2672xu4smtLTVP4TqAcrxKlDL+1LdQd0Lw
1HDO0RY4waLhhLQltuMARdtxBJ/q70GI1SoHT1NUBrlvor6uCedWmEP0AFNDB9QT
HXLuI464uKjc3eXtafPymcoEXoglRyQ5Ebbs/LesNWXvxrDf1vU2oRQt7tasCKox
kutViopVX+XVYM4hwiroGUf3GrqFo1LxIU3VNQXd1Pc11shi3NDF2jo1zQYSv/yI
vB8VB2k5aMIvZ+AugeXKoFWmtS680ny776OuzMiiRrlCu9w1PHIiikFa+E4v1SdG
eT93Ujpjs5c9ucR8g/n7SitwEnTk6MhDSHwFCSod4k8hZhZrQnn9n2xY7n+I/G3n
czlDgTwkCsJsXJ3aGm+Qxswp0QmDJsQlT7uJyrLboriJ1td8nmFTWk33b5LcTE/r
Hrvzi243mFvew/uqlRtpRTilXacK3Nvy2jyAysN0qvVySNO5JwSvyhaL82O9gbZ+
DWAVyIaDQQa+psRMrRo1xO+nw1LUywTDc+n9AqCL01tqP/0GSiZQ/8D5vFH9OtpM
`protect END_PROTECTED
