`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qS8hITPp82ueyMOHWn/kjxbIRIwa7ZtCMkkq/1Jo+dMk1I36+XBER/pa0LPpweDl
Z1BojeKOLQ4B0a7dC5ovhp2Q03NKliR0vRDwraoykyyh/O08yjD57C2/+rbWn2xY
8afXeKFCNw7x09aNF4l8/v03SlnJ96GiHR/x0UNMc6LrB914J7MUJLkf9x5X2GdR
d3rmwn5A9hPRLssiWsrJUFbHOIWwWY/tdklOIPIY58GYqybuux9Wg9ps9ON9mOaw
lOfFpmrzuj0579CCx3QELEMVQwCXHjpgFLq97GCDE3PTPI/uLAfBDqM1EtXfGh+Q
lq1zAu0bGcjcY6IbAxgcmgzi0kc/NRrnGIpp8QsxZHutrjpsKb5HGj6KpRKZjvqe
f+mH/gRbVYY9T09MmASMRm0U749BnzbC5/x68uXmbQhmGGVNrwo4YJa06zS2ZlXu
BAtxmRGzskkTa2xD1nkiYbFKUDVvaIhDdNnphePtIt573+3Q+6FSvZOZ7+/nMM2c
gpTihZ5MaGF3fozAq6dcOIS4UoYPILOfj/SLcakj9mIm7HqgN3uxRIzG4JOm7n5A
ZLw2KxHQclt1TlZqpbgFrWVudBRq613MnhtJmD/pMCF6zWuP5YMaqi0i+2lDu9VD
MZiGk+5wkwYe+jH9U2n3JNNQnRtq6oyF6CbcuzBtDLt9DKisWR5yPLR2dmm39svP
QfqXEponHyibM5Ksdbbmkyog94U/FLMWftCBzk0UZ2icVnekIUsTW5QlgDVTP+Jn
STMvcdZegkw1yAxVmBCgyFMCPn+BK35QLkYIiyiCqvruQ5OmTOF4wjQ5J0Mhma67
lybSTeRgi43sNrYy/7/N/ftDoJ1kmYiBjo2NIV+M/Pn5GJ8L1iNFLMT5BKsHXkpV
7jll2hzsk7jTtkGB8EWeepzUg9PtMkJvYWP8t4PAQ/2jc3Gw7TrLZQywboYrrH1G
tpFu+23tx9R25TrpoDykyhrextHDZSJFpX3ZW6EH9WETFtfK4gEpEG3tygAFBF+y
4ePpcKtTOn8hvp2KmVDL2OI5fo0S2LuU3juqf4vk4Uq/7yElazfGLDi3//LzOanp
EmeaxQXu7+aYNAM6vCNNNHXVKpLqGuDEnWLKtsDQ1oOhlXh0tZcbtsQeu4+qYa/A
M2a6ckRu/jyjQxs5qEV7vrdyv3GxVIeuIDByZ47DLtt6gkob2hWPQWagELbNsqyO
/rcspodGMZveHdxY8Oh0y4WekjLV7FgPTD2uPFHSHwAuhjZRKlIE9czkOPHh55Bo
8RoOjFEuo+9JcSotklfBL5Z5g961+Px08wf02LkAThIhRfq8xYPKueELjRrZzfE1
GqLIQQ2oxk/+tfZQJ4Qw1jGlg/YcseEUBQJNqKkR+gwqmL3GPrEPeNIIbMerfvBY
3OJ705a0JRwodaoT8bIHrx7SZabemw4AdoMB464YdkTj+epJtyVvSt/dkzZ2aRjI
lQ6f2WPW2OJfRJ/Yo+eqrOEUrhPasYAL2xkt5tnnS/TZ9bDTUvdvrXCGFsf3ijnh
s2hHdQMTERpui53IvQd5x9NR62fNHeNlXZ/cnxLMt9HbqUZl9Xxdj/Kj2Lp4J26v
+LPgKjHz6HNcJ376DU92YHmJ4e+1I3b9pL2L7ntiJ6W9N9QqhkaHlUmQsfPA30mR
52T1TCoStHs3YBFd97TvHo6TrwP4qUT75jPH30pmQ7zL9OcNK3iEpGT6tASnwDwz
5iHO/dYJAfC2etqoopHoCEnCKYBFoIh0OhRyyNKIyHvSfB8drP/jeFjHQ8taGQll
UDAvl6VN7IyYfL7C/B/c/TMf7vv7dG/PFfWC8Q7ZG7aJLcblm8QyqrcFxgGzIPVh
mKjhB3VciIeopeaZcgWH0mma9rkkgAp+fR8NeLchKJu88xNP0N1/+sN6o+RA2JVs
DxevRcJ5Ktpw0MHlcgjhgYn8WD2MLCmzWB87FV3F+tvEPe1ulb1JiTz7nqQgzP9x
gtpDc2jmDkKYz0AGW3b64ou8TBcYAaxB36j/dBDpXt/gMT+XX6CMm5ewwvDau93b
pL/bwyNr2a1RcqUcQraNBQUZKdkscStSipYojYou1gEqBhMIQSDgn8WS1GhrHYRk
XSU/uS4VEG+1U2fCWY2f+8nIQUv5zBzePI5o/PAm2DbuEbe5l4ynJCAB5FXmwR3h
S6dFSftng2Mx2jQz9/EKbbShZ63smERdWl/kvkqA6fIwidlel92NkTLtoYEBOnJX
IMWSoYw7TmoYaQ/LDGqQ63XhgdsvZKvltn83gRSd1LF/5uLPeGqE+4s4v2PZ7gw9
ykNQm1gHGHdM/OlcM2JRTSkoFyv12+Qbq2H5lku3KFdQkJF3Ute0PQh/GKFCrT6o
8C4tJCKLDepSyxZ3FMKjIcQq+KI2Z+kRpnSDUoYoAmv7hd4kQuoYjLksWdSmknnm
kk2rLP0DYa93DhaZBbVz6UOeoQcucpYs5A996Yk8dR0LILYMansQEOHQsprinEjj
jZCFMxNulqPLVyI7Db8wTwVzkyugO68XGJEhjBrVGov95+ihK9CQgu0VUJsW/v6T
9tGHdVnmx6XwpwZ+CA/aS35vq4x+u7Q6ujZI71ArWnbBhpI5RSmz8XOnVnXmghGO
TmKV4UI7lSkx+e7VlNY3YpFFI31AZPr0EuIU30HodyfHGmS4BxaH/Ko9mKlMB3se
zNUJhQ1h6zr/XVj9/4ds0sgo1xpAN2VAizl1yLYIb+uqSJ6rEyCmJLOSrARn4peS
`protect END_PROTECTED
