`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdT09OKPHVHvoYpS5UydX9jt0DHI/MZI8EXVyST3gzZWD9y13ziBsjpeJbs3eMxU
sGD9i+CS/osmPX3Psd98xkFXdCmTxlWJJyGHX4VM1LLeFMwRDvtk4SbUYO4acAFI
otMCVoZ8v1U/SYjFNONZ92//ANgzhPxFEV+JoA8CAqhN04HK/NsSpgBH8YXPH/xv
PXMBhMYU4Vj7yuJhtm5lNhw8YDgY2J42G+Ns5vWSYvRIp8PAjmwqwV02MB5b2Sgc
EMyz/Ib2fS5Wvj7YTLyEtU+2ICsRZ5ZEcmpMHP285ZRY8q/ZPrZHW0nHpZUL01+Q
mBoVROzi6h0dMC8VAB1f8FsZdvbo0i68h7cOh+l1bD5fgU79zJYquSbG1KABOCpW
4iL8TOn6bSLXQDtSxuWtKg9Sh0+f0+tbWfLs9cINM3jAickk0AwSDyB5q/+uK6ex
mVS3zr5nggCJtl1JnT5w388Z9ioIqFJiLrz+lgh/5t2n6jQuMzNBiLhDHLi3HGH0
ncBo6+A3w5Ihy5t0SPznre/wbQDA1O/WQkT5TyHo8tv476Tmda1jPk75ARoXeRKB
oGZII8r9dbiaFhA/GfoxgiNW+eGnVHKSzfGwfGlV+H64PwL8gHyLLkNjt0NXNkN5
hci+MZeLw4++6hKXMPoda4VJ2T/0e+sZnxCC7/ZqdoLfZRuPwBrlzALSxezgOOlL
s5TTIIh8kaU7nJfGpxKPuVtIGHWTiqoyBVt//PnNkMwuL5oHtumm9G65A9HIUNIF
aSWUny3gv6hFvfUaYclUCWm4VNNBgVQOH3eJrhodqmpB2XwRKyRXw6pPJpaWA8dW
ul5WUDWhP2L6kw33rKorNRm1x8pimOMolaKe4OZbCts/lZpjTFne0/Tsx94rZCB0
fuG5j4tpPqh5K2y9iUCkyRtnct+pF6kKgLBAdWhAo/9bK0ILb9LfZ0NNTq2A8Fhw
A1HdwTtZaIVniE0F35oha28PdG3sSgWrrT4coGNa7cB58ur/44vDdMTInx3unmOR
tW8AxCioZpXaR+FiujbvOZQT0lAUVsctr3pp77rki5ZnoWbQ77kXRLsHOaIZfh9W
Tb8b8JI5VuAgPC6Xe4wBlxqpBS3amaWJy/QavvRq8HBcaU4A5SXJPSa8yxxf8Dyp
Yv3RVu6ZIOkODFfiW4IIuJgJlw/sL4ykqBv2QVIVPRzyj9HlrVp5OLfJc3RUpLNa
qFA6oNydbPSMj8c6xqPjuJc6wQvzUVpKfQ0XoXM7A7+Vm27+HR3k+60scdi4E4+y
Fzb1TkGPvIKi4zQeyBRY7EadhCCLoIWtPwyuI/kH0uFkm/v9jb+gt0yJlQJ+HrzX
tMw91WsjAJlufu7BSqcpbW3BCnHu9eavCetX7D+OLS01B4hPaplaNDiwcmnOKtxS
lAP7t+r44rEaSmZR7YdU71yQjknriko8CIZegQePVKa0nZt3J7ykIGyI2EQ/VVFc
YuAQAbTATXinSNOiKye+SXjAPiTqzI7LF23+wTdAcyteF85+GM5c5lRu3kchV1oJ
fa5bI5OLxy4IQUBmsZ9+oBhA70KKIiO1P0WSS9nF7zvPbepTbDTbIKeCBOhD4U/c
UTq3XI9ezMJk3uWJfcyTQWIiUn4p417gJeRAVqIKuEHzKCx8FSeco3iLfjTyPV8h
Iw+oRgV1MxSdCK5ZX8C4x7huxyaz+L259ogJT7+FXttXbBmCM0v8My42BKzemjam
Ej83L429SQvENibP8GaYskQZ7m9WZCx2qwqMqkYIgB7Xdo0d8hxXsgyi2lOFuhQB
znC/m0NiK9EvkZNWL4u3n85eZWmAJrgsXDWVbsnjJg2p80Gm0yS4rFxoVag3kDzQ
zHv/zWY5t6E1OqdOAlA6scXdRkuV53uxLnlvBRXgfr3bhkktNSKZSTOaWKhv83tA
33xjY1Gz88a7fpx+SDWI7nKYz8ZoXJuQBW4tN6VYMRy9Wx5SoYr5p4xMoL5z4HmA
HiE3cvIeeS+eZld3LLSkfJlSSfI5sR5mCwmFWDxe5lMKVsfl4tMWDmb2lAgBmw/H
rSq6XY+dtQIiHsBkhYiKuG9uigUV4rXzc/m+FWaqA8/Op6Ue0iSHaWwHE8s6N2Ll
E9DHgwYlYR3AcsV66ex3F+l6P5BLD/J6iUTKYbl2G+QxMaJ/CEmg5BhATLfBrKL+
m5SdefIOnG30wBGFaZSU55+r1lX4+i5DMKxK+i/DY1QTN5jmBOvj2/OExVE7MN9x
ApKXS7OUp+AuP4xTvj14td9myavQSKs3KCO63dVNIOY=
`protect END_PROTECTED
