`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7IbSv64ZT7LfMNhjyqQmbRv1SjssU2IxYAMOOIpiYdCK+V9TPn+CXzJ0IWifSsK2
rmflDvuXQOlT3qY2z6Ws5Xw9M8NhabSCH5GbH6GNvTOAkaOerm1Xe/d1dsFnFr8Q
kH+AnuDPY/IJHogdWAjZ6eXVQ/yixm7Zm+xlYeV90Z2+pJZ8TyDC9vSbGQbV1yAC
2a7Vpij9mVDr+zpvQU4aAvgWi1G0LNls8xuSURd0GOgf1lKI9vCL8FMm1Eh2eIKi
dLDJzm/q7gw4nxlJ78hEobNvBEuO/nxFg88MUoGQ95wDXF+IcWw0OZpDCNGcGinq
j7Xamy9ykmBH5tyTIiHk4k3Uv5ebQMw8zVsRdgkDcTwUqaawJDz7a4E71HiB6SRI
UeNrhJypzD/e4t5nvVhdH6lSGwbKUOr6fEsf4eeYXMfPJFgIR6ppJ7e2BcQO6i/i
nkKEl97YYpajtudGctFiASehYarBnfwfAYA5RxBMO8gIRLVQSaWr4NLoDswmtpzw
cjSBp/gtcM9jvVFaTeO019DS0Y52PWTOwZKS5ga8k1PJNiHXZTrP0OEPgHkz0Xeb
fk/p8KpfEWduYjoi0bqYiAMr8f3qQHFaVksQuBR3NcgtzEuhD2Bm51oxOtfUz+r3
KyEQWguBR+SpuG555QVynYGTG/HZB9WVAbVg5tZbFP0kOc3fbvJNP9AEiCEJKG0A
hKzZmgCLadR6BJLYnI99RH2EZCtUtwaRUTiFIVWMakloTKniog4EJXVXvKRjnRHd
mGjx45lac8IYX9iiw1NI45mmCa+R0MkG0s7DZOE359Oi1eYaKmH3lpnrhEd8a99p
KU5grPXGc/iyXDOwEL672A==
`protect END_PROTECTED
