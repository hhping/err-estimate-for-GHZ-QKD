`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oikPlfGbA9jOVqhhOw38wL/C3AXahSR+sLNSC8wLSmsyGyUS7ZTup7KPji9e13El
3h592bN397ixZEvAviKbyHqHixM5tZh4zTb2U2xKi/I2WgY5MHQor5rLEI+4gvKV
gz4+fLzJx18C2DiQujC8rZY2+awJ45GlKYzQxjGApzwX0fGvuru/kcKl5H5e+nIf
YZ5RsJDE434CHrwk86+FZloXT1HVtyV2U5WDOrObdgmdF6KRY+YXovveZuifBvYY
WKuKC1tARdJ/41oDRok7035mzuFvBJTjThSDCX04k2mfuIOOq9FENV1BJHY/31qP
SYlLlSTJoHc1sYQHznhFubplPLCS8fC2s0KjGJIj21XcCN4vUp/Ul/S2AKjBmxvx
1Zt9xtG1h99ccGqt5Nm2KQbDEpFSiV1X1xkSUicrZ0F4pOn0ev66yTqW1bTVlH2n
lED1r5r5yFzTp4ohWto3WVR9CRfCRJhdGqL29UDvFUVXIIJBBoG3zuq6fERe/z+5
Ox3XCo4lxF8dG2il7X6b42hGaTy3RyYfVdcGUwZUPLk9Z7Xyiev5tOby8qgXwFzn
SMJdnvmENXLPmNbhMzIrQ0gZqHsT4ywNzdq5GBYmQjyyyWKh5Wkv+RlwxtNissXr
VCCVbKY7yKxuMhZ1VojqfOjievFrnqfr3Zc/9zEXMrEQEofeoMJ51F94lzF9tcFy
K1MCsfD5T1JR1BBh2DbKu3d48Y0+nzc/TkSziCfZCMEAgO0Mke+k7knseBt9E3u6
GsYS1oM29tS2NSBxzlhSiwzv01X2cSbU0SrOYq5OBsREgSQ4i5JRHBGTBnrTrAOs
Usm9wKHMouSmc8EwNPUQ2EyuLj5aqwnHwgsP1kycuczGlghy2RiVE2Bo59ZqP+TR
kN/80wCLMiZXiPWdm5nJBfMZz/+S1JhV1BtZibQMRKa2lWM34vyGm3Iqfrv95wW5
5qAisr+l3Qt66wtAK58wN37oLqfpbJLJCg97tb5TWvDvDbJIZHzCKF5Owcq2O80T
h7My7Lt1uwZPezRU0mw9eruQwF5PoyO0gqOhFULYipw1YoShjp2bxdPalL6Yl4Jg
NiOktVlpEpMJBq88A5HrTOF7nU3PUxskOHl6IMNudkSahyGbnOJ9fZJR52hlJNop
322XlfyoA7DO31T2ZUYrmJ29paueckLQ6Ez4wsJQYHgApEKU7aYYhjgB6UzTvoAC
ZJcAYpX2kS74zg9fvHzyzzzfPMUWmfms71tIBbdLx97EdjmfrynG3ua87iHzHY6p
7+sGsL554xA5YWUV4Qshg4qVGnjm2g+q3AFNB0bcoYBAr6l2FvbwrdV6YdPNTbsd
B7SQoUJHsPlWdrq9ZlIAzbCqcd0+B3X3o3QgOoFNzddGYjE7Q45ABMPR6+9cHXKN
KZ1HfS0A54ZO5hCvgDp982gZs4GTIvF+mKxv02fwHrEMJBXSX7u+qEDp2mOha+kO
6oClJyU//DnUfRB5zcmHQOUDOuOGQKeUqt3rFRvmtgo8kQGzi1NT4uu3rhIbu/HJ
IXJo6sbBRbhqEabRNBHYTNqVAaMoIWf6u2/cOCLHN4ha0O8zVmFaaC0gxzlt39ZG
hoaAItOkkzA8RAuya1+IEagdmTA4PQOOpLxRn/bwSBqGFjmqJWPrGooxjQrxgwf6
o+xhrNIgLM4yEFczDAKykLuGyoaTEBwVfh7kYfgkPC21fkug9hO7YLaSwvBC2TtK
OnR6IMsBp3L5/FHxifXwBB5R13Pp7f+jJfLFbRSxFWoEFHu0y0qS/IsrqsAXNhS9
ur0au16ov0vZmleBooxBKfud1HDhjR04gucgwuybHKhC/8YACvDbrK8e1PwsQkZ4
rXDifZl6Io1vqrdcwWOgkbtijQKs4EZwVOIDH3j3OA7mtT8sWiYghFxm393tfXrb
gJTfDA5lxZTbqYgSgdqnM39GMmL6VaYNUTEBlzosmlwHNN8cMbcaJsIoyeMcb7Hu
5ocv1vOpc+qZZM6Xdrq1aKBAmbgS0c4LWxkSr1BJLmucRw3QN0xMxJ1oDAhnuXfM
SKkAVDhCXXxerKBW6+XpIpd1V6C+DrQWwaMMfySWA9kdttxMEczSFFWH2hCQ0INM
6UINyubgPwdaNdvVadYIL1PlHZEFU2b3YFz5nW7NU6tJMdQQ22u50HwEpLHdfknH
`protect END_PROTECTED
