`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRirfcEeu8ZOUsx/SrUsp5/L+txdtbi21AWsgcixOdkoLUSES6jpQgmc0KUVIHsY
+GvA57z88GAQe4DvszTXCgLghijwhOEbRhyfAplpOp2H1u+zvric21Vd6SPrNNXl
CQl8/RaKcw0tYi/gY8QgITYqbHFv4Odx9epR0r20ziY=
`protect END_PROTECTED
