`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzjrr8wAlye3RoI0AgxOct20bEesiHLEqlIdJ488KdNPKvkJ8kQcS6D8Iy046thw
+N3AFkOIgMG0LuvsjZlVB1VOXZCHbb8B/kRDeu5JBwtJPMNY0Usm+himf6RzVVrQ
XZpdS+V+KbbIayfySn+saydc/IFnDiw6yap6cWxrFzl/xtHkm9JdL3tQ4mU9juJu
TF4o85wlb3iRm8Q+a6mWno22ykt44ZxWi7lEzvD+KkPZ/O72r5UnZ3HAF+PAvTIS
Axt6MoBnRUovVnmAbSejXj28iapCbA6pAK4xQuqCUFHvpnqVoTlEukROxEiP1eK6
PobaYQ8fSAnLSrSSJgo/5zo3G9oQ3p15JZQstQwr26oQjMtA5xw980Te8TQ2EGhH
B8xhRwTtyIXMG6ViE4VwO3Qr3/fbp7BY7d8nXsM89IO5xXhgZ6cyQsZl0CgNqODL
niC7vTSHaaVfnT0GqM+Se/nnbiEiUk+/fB9KRlV8XJKYUMmy+A5B7Jvb0pS9KF/C
/7rsALR8RUzUPo4q/x/GXA45UgdNscF2+p4m8Gnad+mcQML0u0rijiEI4Sptq6ub
Q5Onm9KMPEkmkyIfI4aRO+II1nBrimcfzVsxtkyto42NCCkvGy6wryi/NCcvjMiF
PI65WF9K3ePcQX8zAbueulwAALY/Z8pT4ICwm+swkp93t0QS7m1atFC9klWu5c5i
Tmf/z4Yee5v0znC4UnwgjnfQHZbGaW1pJWrseTZIX5YzuwkvK9Rj4P8Sj5ckC5Uu
m440yfoNLVV0UyYyQNgThDCLkkVEu7iWDQpUZZQg3nvXZYO5ghZJrTWtL1Y9H7Dt
n+eliY0xwDtvZojBkw3C7hz0xRqawLppXfyztodOw5shsdTRBRio4lhT7vRifJn0
RBtJZa3LngU+dXOmcGR7e2o5rSqTpQz9MZ1N11wQQddeJ9e/oiNezX4I+DRidwd4
2TYPEvjB92My1Axv7vJNfOxijQl18QxstKhg+Iv8iB3v+7zG3kbmpW53uftINgKp
Woma/4f9ye+77VCKoQCopljJB0WD5sk9t5EcfQnvid6DTJ9Zp+ubHVMeySL1H7aQ
Ek13B+KVfJzlT8OmaER/vLSTXOxwduXX6RZ5AGNE66FgFb2W1jOe+QICFinx2F+y
Hgq0fQj/Hw3DISqna1wRBa4myYh2K88RNL7JhgbbIbtoJLSzprBDYv9oWRc14rRa
jYwsL/1EckTpOjqp+9g4laso+ZoxPOX+nte554ddmuGBhKVAEUpTEwPF43yg2Ad2
MskUSJnRB66RE6HI0iNy1mbvmjICvJBU6ILAAUSP53UGlxQsV94wtuooBzMNsapL
yRjVAblWqCo45E5MjSRrm92rye3MHIFHpjVrBvdsU99tJ+kj42XOGZciAvZGLstY
FF9/e8eLKxxnLxHjLgokvXzmr/a1kzDgMrLms4lJ1SwuZ21IYvnYDBC6DOMKuFkW
kC1VJ2+YZ+sil3K/NvGlChWgoAVsLelv8BQwbrShgRtL++OB2aev3i5ly4yuuBZZ
rUjOurC76JW0zZB6v43QusgSPVxN8FaHnVAc4Jr33hec98vcnAAQ4uIBmFoGZ035
aqVU1Viseh0qdIhdw3h1LdHo9l2eBAbLu+akBVEFCgb2Crk81H+WIxnXj0Xp4sJ1
0nBYz2MOMbZbXJNgSN70alyrSBSyIOEkQ6DE9vj/8HLjaILR08TlH5lPghs2ozK6
pbZi5cPN3n1EnmR6NZinX869s2NeqJ9M5kSXRHgY2B1jZDs1mGCtbN6pYvMSh+Si
5c8njm5SRHfG4m1hDTCWwpbQEr3MMVxwlRskxRJKiWcODmmlRtwEfQmSS0abl0/U
BlYMxeJ7x8bNOyMYiQyq+yFY//kIq+0M1yAhbDC+KoIxBPYL90dLOCs4txLdavX4
OtvoHXMMVHjw6+wi9ZUKEh4AfjOYqExL1gHJhA0Uxm9Hu0FT6tf1r8TJJIw0FFWs
dCdBCOe3nBPtydMvCpk/ZGTn3v7bnyj/wBH9KTZxb282NWNtw40F7FdBTueRDpgk
OZ/H16PE9cy0auiLycTwD+7aJ5xfKfeJz749IANy7b9GJ2MmGrkOUeq0CINmwsGC
VbvYtEjW/g37Kzy08W6AkE6L2r6VY5SEIcSGUDndpXEor11k6RMyrVVvy9hQEt8p
GCEQgNDG5ExIXwAfFxcvP5gGA8bgPBPnoH8Bdy5JBzwSNj5oVqxbLA3rkpLoUVAx
Acsazw1gnZiGqWyFsPouz+O4ZoOSIIMDbNWHWKv1IZmv/W8Dz4fP/SRGgyF/Iy7p
7HvphgxCZlpQsLi6SwaVkJkDmKEplx1HyvB/lxr4X/2JBgBcBIAWxohJzVcnBQjA
jysESyOlXZsg30jg3vEEjdpo9bM7A/spaU9rn0fHu7c7aHgarEYaXyCeRYoqqrpX
TRbDZMtGjT5z9zTWK46lsemnH5J897LeyMiaNzumn2xGSWy8E8d0qUG0pAHk5mEp
3KmOW9hRKPOeD0mMjcTCMMOzeO9bRLKMpSsoMn2htbsRXoOdSPNIP2DxceV+6Aij
Zv4eV82nGN67Lg98jTO4P6SV/g/I/I6tfK8tU4Z7V3H3gLY68ijM897AQ+e4JWAn
xZ5h794vOAm3lccFQkYCwAdJKrFRbeU2GZuggafPuM1iLF3AcBfLnbfOz83aIdvj
zdnu8F75VywOy4YIqZGmC/3i0HH71C3t5/A1jlNYovVUCN6lkSGB7hgQ3xZx1WJd
g/2espddQj6TyF9cwpx2c8tXBVLXHgO5sAusSw4vTqszszFSXj59F47Susms/09K
nSn074NhGB0YD/RlKnxqK0hrsG0gFhhV2SZNl6mDu+sa2iBct/rEnBi2YndSHNTi
Gtjf9AbAE983CRzZYmrEdHykFXjkSJr4paGeg6R5c9TwBU5O0tCSW8h6BHMnoDyG
yX8A9d6LHweMHp4rpSYpQFiSnRTUlTy2o9SNN4pRxljwwnJTaCJOJzQSProx2sng
vTAsyzYvxyMMYm8Ph0ezVPuDaY8YtEOoI/tQBFhznPXYsjQUPLv6Fo8tGclAuPUm
TJS0FWRUJHn3FthQkREH0H/uy4yHTEkuR2CdiRtfoRAVkE64MWn5TejZD2LLK+XZ
fp9Xbsu+ELIVYI/17mBTwh4XLyL1WSIdfti60oQDm3Uk6zmcLypZFW0kuB4FkvHg
kRo0zHSJmTKEI4v4sm07CDSrSifYIBGi/x58rlawpm7AIXEpApmgvUX/2/6QEy+m
CipYxp/SDrnBp1WEEEQtBLmzkdgmbcfFAeJcmc+AyhfwoAhjUIC5g+Xi0mStRxXR
5BPkeMPg2X5vC3v0vJpsQkTEuTjGQG5Jtw4NKV53ZIING2PLvnhGJ+4wQKVDcHMi
pubWAMIr2JadcO2qXXRDXCtGCrbdbsmY80WmASYubrjsLOsXjn2tP4T2XvFEA5y9
sd2mJSMdqnnspHTlfOimP/jD2fr7syaOJEMH3xXvL3wUZqF5CzGcQKHkfGmdecC7
3Lva6dVNjZjqA+phJQ9PbE+3sT21Wt5O2OQjXk2PODtLh8UEA3EtcGAmLIx++lsw
0quEB/ppIO5zSgN11TRo9dvkNVOeB6gymjeaDsdHZ0dTLQlOUZAjDOzoiMnsk6jl
5/Gjf6NfEvs2gcKuBEduLpp/lzdAofkmabcUMUo26vhd9HYAph2ZCuuc/yP1uEFz
TfztlKXNzYykQKLYu/rwDHL4qIsGaRV5xAGS7EAe+ZGrN+XRCoMsHjgzx3NJd4ev
bx+AwE/pRr1HQZNr6PTjiYWrhflbtDJv9CpIwbZmLWXPR8JQBAIgKFCrOyWL1MRT
MS9adNIJ67oIBg+86xqZTEBUmTtSjgjYhQmK8soB1CUtMObP0BE9U2iAtwkirAp8
ef4JhdBoi37RVNbuWTP6bya2/qiIVp/AYVk6LdoqvFXzULBT+SkugLISHwOv7U5h
brH6QZyDTfbY2pSk0mtP5rON81AudZD7HzI3ihS1/WwwjwhS7/FTesOrYOW8wkZE
K/D3Hu/I6b24242O5UUVwN9nn5HfBYEPmYJSbB7ynj7dep2f1KWTt8vZeJ6vGPuM
nRcFcQFc6bQ5kFQHlj7y/0lj9tQ7ClBjDCCqCTsYzOM1MbQNbEtxQ7SqlxAqBDQb
18NvjLrzLg/QQd1+f8P6QrFZo2Je70DBMeQtLKguobChkq7o8d8Dkl7qWIjRUK68
UaAZhEcQzzYBYw3Cbex/gw4XIAbSsdkccMB5YUDbnY5QtboHIjU1c3SitUm1athO
0CJZpSniQSI36xa64bs68JXbgvpDzRH+EI617yyKdoHPGuJomm3ASExh0K8TRnt8
zuEiTNwqFohaSJqg1DON8XRgkszFR6dnQ0ALw1+2ji6mSwEar4LGRAnpUrWCvzdz
c6YCb4IAK50IXzAh4DFJ8wQykufC4ju4KGAi93/lwYrx6nYKTRixgCg2fi6qvVVf
/1ME4wC2JaIZYEMDuewdtakzvK7Z5tFqDTzaMyNw+73ZVK/MxjJuvBlZukFSq6IA
IFNvCg+xHDCgtoCqZJy9p4vPfuCAq9ztlsiC7jdkJXJ2/5UwMJbQvG44vFzdMnXv
WCkl9YgYA9qHCTtEC/yIoz81qWwEhMlBFbWWKa+Ko90ej4UlhOzc1DpoHMZcH7FU
a6vMH/uM9HpE73deVJQzbr3uf5QIrRIicsO7vvU/Vk8TqUSfBtBlgf2jNoB8RLq2
E0i5HBZ4c8JO5uwTaKPqDRPxYkPqh3/2YIOCR1kiNv/wXfA6QgROYWi8gs+7QPVe
nePTNS3sLDqz95F0+EJEJwLLp0GkaGG1NC3BHJN+UWVUE7HL63/6VLSuopKSIZsI
WlM76cR4n4BKfkIwBP4AKu0j3MCGaTMwjvw78WpiO/f0QxGP3e0kdqGgczGLf1UH
9yH+iwH2NiMoMktvUZOljfhXFjWpPyVpAP0ogj7/Mcr8RVTNKmwEK+oN2beJBiWo
y9dJOEQydMNbn4s7qg6c/x02BAJw5TEVqzlMmz199SMTZLyY/MIhGeu8nsOBpqUm
uVijrhUmcYgqFJ1CE+DeoCznKZI67lJHHM/dqZA2IEG1pyC8NG5T1bWbTgMJdclR
a1bJRnLtaDvTkEZ6WmmHnVG9Kf/P7D6HESEmuvAwgzbst8QORgz4l2uha13wCj1p
b130heuTnIiinLYvjYoSqqnWJRt+B8hdEU2ZtEuNq3UJ31sKTCj1zPCIGRj2Tv7M
iea03YSVcK90Ehp8umDX+RXOhfIGg14BRFDKui+sZMHnQRi4nmrQVZu0iY1fR7nM
pKzUIYtBMysxb6NEe7UD3uIMlCtNv9etE/4REeTO8ar+rwUnRyqK7jSZtEDRoTTl
s4regwtRaNoHd/vh2BmjSo1BC9iY9fQIV3UkjVI8CO2QpqhiiBV+0FYkNTlHDLuj
iaVJtFCge4nWNPYrhNEeUiXAAH75/wZb5z0esbLJkrNxjI0nkKqbq6Qeangc9BmD
LdzbNSAZetKoWIKKxWxedm/DyRmqXqtddNeNHfVgSibIQw7jKqU/hIMDGIMXVvY0
Yyif9P58ydOIK1nafjlvxw2hAZoAKYb5jtk+zFPCCVYNmPgNXZeYNuPDjS11VNC+
qtA27qGx1YfRETJ0/q1z2JCB+qEwxU1iRgRqhJtU/BHDdCUQ+Oo7DtfRQewhoyRR
YlZa3HGaBQY7DpPSYbcIrOeGKGEBVjkmtLDCorilvgsLiYNa9flPkjTYpA4LGw3Q
88RlYfoUkRCeYVVXJIjIx9ug1JYvuOVzYC/kiS32vsD6XqTrP+/VMnriFfBbcdtI
MU1GqtPl5Ua4EqQu/HILpO9nkfpaOzeqHoznDd3s08raISByuRW3lotUSqMPF9f+
P+79ZE/d0BVP0qHttaZlTN48RX1MT3XlD645ye+Qd7XayT9p7A9CnjWZnfjsx2y3
hvGaV6Eem1RmG0egsDjwLtVLPvR+CW/dM0ROFnGnQ/7VNCCvQFru+L5ucd2iEGZ9
Dl/922zBKsGczo7fxEYdZwh6HCMHKB5xXTW9Ks62txIbaZUxtz22tAGx3YiGt4np
Yr5j+edEU7AWXlR8EWrKRy+p86BeoUBwetPoAVouGKHIcPXhMa584bgblgEH1QOz
W4O5FE4P+Fn9V+YDeOwOJI39AiRoCXHtx5P0el8hZSsF+J7zHq0jCXHU9DdxrDhN
9f7vLWpYn7E+qCHhNeEHQr/5T04K//gwXacMzBPau6ri+0bzZbbJHN1h6c2AaqYx
uXYy2r+DOy323/SBgKtFJZ0xUykFsuoIMXz1DrBctVK7KxytCevhC+cXAWnxyGlA
HgoEqbBEXM88OrxPBQZ09Xi9qO7A6aqEuKLwLYwNIIiKyPCrNvDgB3TXy00ZizCM
naxIDDTBHU9ZWj83Rl2WTHVjDYCohuaizoMMue/QQbs4fj9WKuI8/7kB/NvWOhrq
JnE2eTi4am0xRv28WLNTBdRNu/Oet9LkRAX4tsCxEqGmNBDpdzaTCKkanXHx/SzO
rh2t72o2srQXknEnDPQ0n7o/t/++O20t4RCEYXReFDb/hX5XOKzgM9o5nMbtNKB9
hmZmrLvY66ZubqihIe4JFBZzkx0yOtqXNQtvI8TS9WEtuvT+JEmNuHvLYe9RJIKf
FHCjkXf7qHSL67tuoSigFn5rl+MdIxf5bSu99g7jbjF7ZLJbEmMWHTq+HWzbc9LV
6MVgWgf/qFy3spLw60wGpMoRPY6jbRzdhvYjPRjx3xnYxFUIE+uO91sjSByH5XdG
K6dbntguitfOmtUve0CKA+BDKv1+zKEau5bIdUVlVJr/fIFBJNPRFwhIzIWgFZVV
QzhVpjzvkPof3FFRIaKnOwE8GAOuz6oiIM4pCjsjyHaDumhLfijS3yjUU8wGR8wh
eACIHgg1mrQtvrwpPkPQtOCmi6ZTA+taYiKMxl9Qa0GJSrwseEWDQOd63LYmMJXY
exPnn1CuXAaAdTGWg1Qv8le/T2/vOLZb0VW41VoL/YssyatsN3ytnSyoJIvVlPDe
ZsKhFyTowOPH/bG5HaBcwpFgOvKEpPlg1LnQEQbSVF3/i7HN7NYaQbqu+GjUDOkO
GEoMldZoQ1P5585TWHf3i7DcIngPxFGKzaDqoEBUS0PMaXwiWSIhRsh47BrtEZS/
kHlqPIDFr0sDtJJYz37F7aqYYRP91ia0vjJcmKuDuWFK+5EWar8Kis3pWYtTBep0
V2RBe8aY4N+xy/nnpnJsBY/+bIfMA7lQdi/kMcjHW8oTOywzszwMx7KTeaRF3D8F
xNTvPKXS9WFJ4WfQioN02y1OUWCNhCH/wy/PJcV8YAjkPQWEDz/N20aQtlhmbIxM
4/oKbCKfQ122U+DsmH82B6WxQpnLWdIl1IvdWxSQSj34Rpl56SGe5l+fQheI9nPx
D4jvfyx31vkigUOOTf03H0LK2fqr+psMMQXVooaqSjIOTQFxs7wIBODJ+1QH8mxQ
k/F0r+PV6sPZh05Ozp2LSfmT9dm9MQbVcYh/kmhsaUR9Uy8iz7srRpSY6ifIBd/h
scEm7tLRxdys/wt5cAZlIR702VYiJg2VJMZr6fYFphuyziuuRn7JQSnI1uIs01zF
WKmFKKkVfDPnRw4998f3Vz+Qk2Vvwev6diXo9xjsOHuYZxuwX4vErkfrkhXZtY4i
zpfnLu1jGneFp5506ZDissOKTKGAey3EUohkH8WHUm2YWioEJbJ0Qg+X0ee7QBrd
Mswi+DhiZIYnAzh/msz06Oa9ieR0U3qnimDuhLj43IK+xTAegyoGn2CVYuhp86qg
R7s5sxp17LwLVZW8EyZZbQ5dmWm6mbiL4Wru7lV1HAN7vIhg8DvP89JipycWfS8X
luvyUNdj6muzK+53yocdxecLx0+oAxqciaHPMraru/0f1tNPpse32DPDoNLHuubG
szd9NAijpRVOlNQxOkw4hsKOGktC85omwZV6X37RBfnUGh/rYzjwTQ/mPjCCDzpx
wH/ApBs26jZaWzao/2IoYgMAVlBTGcfr/gyGT1hDT0zBCt4VHFz8kVxuQsr/k9Dl
H3nKlfiFBidLiYK1L51CpnrVg76QGcE6AWfOI5f/DEjjXoDzZa9Ph0bsDsgne2ef
tHFmWDUihI3PT3R3kXfAYinHqOsGugA26G0VttEDzwQbVwLTZum9FNHa3Ob1694w
Fzb0XKECfmPgbB87TVdB8EW5bXVBjeEQ/btzGi68rvRXhz4ubfW8QLMf6EDLwn+H
llEPkkFRnGn24HzQyk+OCkX/Ah5Lr5mvWXaa9Id7M5ve+38TA41xHac/FP7OPNxJ
+gRbxKJDpkOB7l6IGFGpdLKPSVCgGryYeBFX/dhUfPS8Vf5RqSwAyQFpKoTn4YsM
sZlPvEetoJonWgqIxF5GcyAetXhCC78fidOckakvovzl6GPgo13BlwkiOXRzcnpq
sa5sxj1VQnQfkvXokMrJvYUJVsvnkSrazeHF207fDHw59MdYL4ruOZXXJ5S9KoOr
92iLcD8WggkCR5O8GzUowHY1qpPdOswFRpRYpToqflhwQlL44ztiwKRFK1pqOfXq
dZPajp+AZBw59jG40iipdRVqwx92adbQKEu3ocXYDdpv+jHmft/KWBs78p05e11Z
AadxVp0wl6nHKlwUgWWo2IXb7RijtF8I9YI9WgqiaiJRhuhEPz5EQJIox2H7vG4P
4EXq3ke43Dt+l5HUyHiUJ+++rVTEqkjYD5FB+x89kMzvOfJW8dE56vymdAUVjs5r
7gXQJRZfYCtZoE8OVuLbBnxJHmm1JnODdWWlefbH6r82evmqbYFrJN1l0Byqt9SO
c+B8YYeSho/377D2B/aRiZeIlGVmLF8PmpwHm8VSnW8M43PS7J0mAzInjA6pJXu2
nxPvTGi7w/k8dzRa2LZu7oeBJXLVxLb6+bvLx3YrWWZwXW1NA2Yk8+RICWQ2coXN
66VfDv9DxabQQD3j4e/64ltfr88I/AtnJROn9jOYU7qz2J4svcfEIcKaZ2IUDRND
snYNGKIAIXKynlJVVHOH0Ls9x80jQ6D6npYpQYJ4oUJtp4qXwX8Ul5N//2dc7sFU
AYG3CKZNCLod0vIZX3HNDieNVDL3ALOSAKIeRVqDbFlx/ITB2dirF8LNlLXvVW7b
0zXWyekEe8e+7bVfVYqbFcUfQU72Sbbxj43lS7AiNQ4pV01xMEMs3rb/8ruitWd9
oKpubyBwDCQHKLRaprgBZgNu7lIOn6SMQemOxRxL0GOUWJ+efd+uAkJmMwWXIBfX
ahYNYxCNh2/sSdjExFFQr806I7CQbzJBjP/zETvvYpY6pKYfv+yYbpbPp3JhQJof
NpAGZ/e98OrUqkdnpV2x681e0/rBbh++67HOT17Ixn+Un+zudJiH0EbFeZagpglr
TiO6eGlDDLjT8rvFCoH/iDOdTt/d2l8HPulAsAYCxC94/eTQbyPTdGuU93Jg8Z0N
loEO4P8WoUaKE1EjGztBKrZN8ZOeUNpy4Qv1NPnHEqhkmiKiTBQAOnqijus8VkXF
WBOtIg6/IeQmke99MpDg7dhBNU/25FIODuCAZ+Fekp36F7sCGiG0wHkx1WRlWxSt
uNJndvzbuGVqLKOaqe0xVo4t1300skWVJ1yMafFw3fRb3/F5m5QoxCzkME4Gycc7
xozGgFdzNrn2mK3a2lXicE/Lz0cyNbNgLB05uolrsZrHsa51VvLPKYqgOqjQVFXt
mYQOLA0dGj/cVbnHPXX++Y/5FXojLUd4WyiqntLhE4hVlQGVbJZT++x/EjFAU4ws
UWxlr3GU2j9o9kQwygL4gXhCM0/DYnhRlGHnCU/ccjrr3lEdvyPQQfYdkWzgeTBj
swk/TgsU91RGEQlMei5ZrOPO9yGUKWgPC8fF8ty0Kanq0QoDZvaq5BYz6gvjZSwE
bPaVRq2hM911zM+f40U177kyvtr3VfmogH5Bu/8f/4fNFkfshozbc4e3e5Oe0Syz
gO8Lbha2XU9qW8tgECmb13YO76ngzMbtR5iR/UTpxdjGJe8Gt2XUidvpeyhGTPb/
zmRdwcApm9M+rxR3z/cxT2I35scJ/HOedsTIZyX1v9xscXugYYs1ajk3t9g6oe5i
Ok3zlDGj/jfZtNc3bQeHXfpsRa5EZffjwYxIOfWnjbhJZ7p62NmbZ3q+C/tL4XWx
rtFpNlt+TWenxiMEZw3QIHbguFYGfjV81a6j9Kr3sR2KaSjzOV8q/WxVIPWZYUHs
h3qCb4Ou2FhwK0CiPHgv8GsYP+FjBHKXBOFrRrxrUnjxFDsUXrvA1YArHGrAbl+Y
iCceVlpcFRsddOBNwb9QnHx7o2KuOrQ109GVZ/oQsYxCKvV/lQ0XeT+DJIvNs5sK
INv8dDU/TR/+z3s4ANJB476KHy0w0gGbg2qovFmUwQ6gcfW4jXOwmb2R9R9FrPqO
8rH6dC6JOCrgkzJ9VY19meT+LKi6Vi9h7fb/VQCqKIWGGeVz8SYE18pcI5Xe9om5
g9qyAiz4+7f1OJtxKIHKoLfA8n07Y6bOtIHsjRQaKG8hNnHvHAKUEduvvbTZABaX
33uGY+JBwJplcuRclIZFolGQhq+l5aDXuqYm4bBczTxRBywhzAwwSQHAHzF6oUkL
KJL9Qm2s1ywavVsUSAc7CllkpT7rWXCvixRMS7aPXJcjNMh5DSjx30OeIN5uEEMC
B5RVF/d1LxGLZKdZ2yPrEwU6EzDiBqHazcHtiggvCIWb9wwUjkIWZXE6nLi/BBfm
Gg4pH4t/mruEuALaCO/X2WSB29Bj5xIe3NyGYMLOniXPe2SJfYA9AkIUzVa9bc+R
YK/8S9YLrtYfDlTnNpxIYE7MyZ1V/ymommRY0RBnREBlZjZ2eqjZJHy1PftZKcN0
KEN/wK2vbVtXyMP8/UBFrRGuhtRR/u30ACkt7G+IZUY2jSl6OUqQw+8VWRqi+Mwa
AkkVG8Sxi9W0r6upsNvX+qwOBX1H9PcXoN5tge6iEMNKuLUx8YUmEB7VCmvVF5Zx
SU+/QY8xoW5t7AF77xN+ylzQcIoBm7xA0mxls2LgqJcB+jX6HYhDaTNOTDyJ0x8/
gGgg89uuB6eO/tZKPbs2Ew1/7cP1Sb5nksbXZMVV29c7wzVltyTw/kJ8mCCi0Hwb
BY48y4o4n7BUTW9i2iAD4MEVfJLSd17UU5YbIMxlTtM61VnPq+uDGQPqt+vr2Buf
JnrnwhrUFRec1H7KCPbBJvcTXTH22WKXNR5Cmwb+djZzOZuRfWztDRzT4zALPK54
hCXekV0neuT1yHlhEytwO4mFtxqJ0GHaxHJS9jH7yghNQHTf1Qs6iewuLJeRtEch
KT174ow2ZfjX6B2j/jKAsQC09VdlYOrhTraVi6P2kIPRPyPMP64rsJV9lEed31vs
U40UDuXC3IT6dhSrQ1FlSKg6ZRw5bTSNA41SrATzVx9LEisreqHEf2DQAH75qqIU
wHVhMR5VqdCDy2AR5CDKpYwZkfB+ERkZOm4FLaEm/VfV44ht0UFzXd1gn1/Po259
APUeSRZ1QiqcO2qWkm1AT9CyNxp9zIDnBrrpamBEr2LyyRtOftSXXrwX0fZmOVIh
95k5wj7s/7FElgOWswNsgrLZW67JUokraSBne0Jqvw8AGtA/ccee/ragg33ZSff2
ca+qjSBAS/trp6P/+21VhBmHSE/w9W6w59jmB7+wlEE1r2yBeBkIBhI8nMbXyvcc
Pilndg1C8U8sjhNXaP1sy6nX9/08vqpzrbuY73e958sT37dJJyOfz9acGuKxamz9
B26RUx9Uq7g4PgQooxfh66JR6qsOALm2pnwXNDfv5QW1jZBBcbzWW2wdiT6MLzUm
9dTu/HEfMk2G5xYqvazH/DuyF1tNjYIIe+47D7QHpspESFca9Mlj7ej84RKniNom
dL4rJeGDxMVcvaEdnKnJjYTLQSQH9E5YgKpotPIBSrQJzddoiGCCmML0oPUbsC49
urjKknZDWt8Ftq70FtCZpvTNuvFwfyT4I0NqfhqDnfGhSCWraoBhjWKzx/87//oR
oavxkYiNPQEDmElEEHQpnpe6xnfvEQ6X6NGzH4ouFfvI1sqP2vDcOYSx9g+r3uBo
3Z77P5cA1dnQC5JOGFaFTdrmsr8BK6iWT7uiW25b6Zn/HutR/DIeONVyHZ0QZTir
VKue2C4G/atzaFJ3pbaUw5J4E6LsgyOCkKIOueRMV+sE71U1m8Dqcy+3XHWERv9o
vyjSRLlysQlGPsXjtI9INUD9zmG0nuMwEtXp3JJBox8WRmH4f4FyJMBRLP80U7WQ
yJ6KVFX4ci4570zRijRfhipOCOwIFGDe06RuJoY1jLDBIPWpfXdIfr6d51VJtoor
MEh2KxHLLBOwZCmuLNF909UYYa1XQ3FFjlwUAoCl2I7ZJFbqCnqFvHfH8lTU9GCP
BNFAAAMiuhqX2uG4rlTwziOSpOp5/XWtuYkitwyQe5xaNfi8OMEE0x1YVeDx2WEu
hHJ82Fw1VU9Fymlb0p5bvj3lombZ3Dt192QdLTyHsOr/wcytNMoHIEcPiWMex5Mk
hwHRaS/X3yqIQT39V+J1fUFMBuXXRy/pDNvoBajLowl5LMFEIx8r9T9REoizpc0e
Ra5vjVSo8qHDYNs7Vb5/zmc9F44wf8SPFIfIMRN5aogaqy59sD6/YtZwBC7LUDqL
CugtC9htDKCn+eQizaTOnTml7r8sBSm/IssY0TwHl6cmcr9VwUaUDzXUBcLxyygf
2cVKr9Db6v5bvYqiTo7Y0elPv7Qr/NGVVn61xbDDv08l1cO4KHo51qlNmyXJEl1v
H32JOBmNZbay4OWhBGYzXx/50Zk+ogX/fEBtW17BJkQcvwAU/J3H2zROJFhbQurO
LeuGlpH8KpKXTJ02irtzITsfcxDozMsOftplfT5R232/raS6rKhOdgZHgfiYQgnD
SAEBMyg9++mMDiR0jiyHn4TrSyH1oqoFCugoUTRdxeJIueAFLicvbQynZ8FYKD4F
QvbK3xLbquQfl/A60van7s7rQHzAdVoaEspRn2pH2iJvOhi+D/iN5BapkeGXjxfS
ST+lrUcFtpd14PVeXPD1BCvQnG2IrfGZrRm6OOzGYiIM7WXfw1UWZzmTED9JxWZl
ZtVGh9AvqZzGvUyPMM87QvKXQKwNksgHmNZQEmxfvGa6MhkDIN6x5AaDG0GGnv9F
ETFTb8uv8/PJzozIzj1lbUAeKpXmW8wP5GlX16Bq6D71rVTpU5zvb+Bw28KjhKuT
riC/IQKi30t3k+OMRo2V5GYfI4eDECYkXgcoVJgRKuZ1pLt3NYY5Qk9VF9eN8YH2
ocR7Av8yHDavlMlg6w5tZ0lQ8k9dyW3iZNgMdoHwN2MWmadf3CPXkjrblJqcq3RC
coJgGdMDZ1K2Lqv+Fse6iWW9O2IJ4k0S30njdAXC0Us6PYdKifXfAmra9KUEOlwj
137NBh7+HZ89N9yDrQ9dAGK1bwZBAIEWz2h4a4EZd020HlsDNmkfuyEeiOwqzn5u
RLR9UHMBx9wCHpcEPIk8N4C4UQacBy/Iz7zFKIWjwXdjhntX5Fr0ANPL0p3mkcrX
dLOOY8IzYGz8vNCKt45TbxKheLtofl+wE5C+JpZd1TdKb+g/Lr1Z6q6Yysv9rygj
DebRpHXvauQyfvU8qyrvV470mBUFyxsR4X+xbdg7+u8/qA6uGl9POQ/xjQ6KfQj8
WyhpDCJ+KSvFfY2UzWQMJJqBcU6FMsOpM53OjwVEhCFmol5yJX1MH4rUnTM/5The
hIBQGxZq5YiHbYHMJk2p5o1WfE4rO/PpIH6ajXE7+Go0maFRUNIY7td9vGNeB9Dx
Xcn0KPCoPp/+S9b+g5AQdpxAq5xeFI5Zu3rL1xE+Cx6Wj+0uv12TKq3sxZhNjYUJ
su1C7/Ny3coe6s7RrnLVe0wzVJbHS2IIkjHDqSoOTtWctUF0GLOv4R0r8RGaFSQz
c22+SiVV7zd+c70DzJ3+rfKXbDio4duoSEfv2bDFG8XPxXU6K5t4n2NYwL4hnp+9
IWdiHgHiWCZ7QzR4cUo/luZRCYyFfFbl191eq/Hnhs2a89VzmnjQar58rIjGM8PZ
olkKqiWq1tduHMHA/ajjHt078Pj1pPc1qDQFKp49EZnT8bsXyKuUCkhozHO28NOw
FxXitb7oQoR51OInr8a28H+w/Q/If8Q8Zz9ErpzvPO9mFPDewBayueFh0gnWIURf
R3QJYmAbfWjtQtwgMxtDYg6Ke7ZdXsXwZGTmHAiaEkkzynFRj1AF8IqSxAduCWAK
FpZMBNf87h/GWyVO6jgXZTLEh6vexjHQaj81yvD1bQjrBsFJ1mWLcsCQGF+3zpUK
IDhu++TuEDDR8zCbiEfATVwJJ/ksVPqdwCLtXHUWYBEFGWfrh0BYpX193N2um30Q
RtaUR1hyviDclEYRu4eWP4IcslanbzaPmxX58dDBc8lfw2cIRk7dpzA7CYShXMH/
Sx9O/nJ8DSbM1R7HcZWO8lA/xOubqCMcq9o229qb6MxlH4pV0wMQ7MZqscfQT+VR
+4rD0EPGtxBAOOPdSS9E3gY89QavF+jcPNUml4QwxME6C+qWEFLMLxjvaUcl3ABB
6/bp4aSj+iSf+H+ZEhxNof60SdCU8/pfwiZsOPUkOsQaCBY1pK4dorRTvn64ULUS
f3PQH45ThJKmvC7qnIexEcWNcmNCMfwkn9eN82WP8DyFg6yc6Dd3Ib455K0U3XFg
cvDZemop2jn2SlSpm2lMmsgVkAw86vyMHfBuBupVyKSoQjEs9JDX/flATanwgMYw
+oL62jyWGMDGPOV4Ex024CDhXn/bkjKdp4GPxZ/2hyhf8A2o740ySX9oGoNwZsc5
nq7HJYwEpXjdvrNFwNaCkRApGQNaLw5qnNBFv2yulsuRphb9mjyhaYphh+QD13QM
XnRQtBn2rB4So/MaFdFJAgM2JQUD9vGR/k0gG49/LZp5sx/q1YKHHO3r42U4jpVe
E1EeCKkzW0wEU8MohlSkrZuNzWrJb21zlgonoWBThwZ0Ingm1aFWgr6h+YaHjsn1
0AmatAY4OKXW84s7KnkwCOQ+yaf0rt7ZQwX0qee+muBh42dYLZZYDDWqOBYZzGTe
MG5enWJ1W0y9Sn0jYBBioV+8WYaz7YpZh8keI6g7QjKeZT9zs1JWQj+LhQyzGAwV
+Ub2AjmvkgqupYeWWu6zGN2nBZNfjWoycsvPkYUGEUz4VjWPS221ynI7DeLtV3JU
Dob34jM9AqvWIYrO3eSK6MmeWb9fK3MTP04QbTtMNFYBX70M+0wK/xJRG1kTR/+M
yTg0k+GG+PUTkD1nsZwJcx8eUBGv2MLs8BWVWudJcHFhthX+KQKjiklJxE7jDIlG
05aPOXswgTn7OMyuma0BGtb2VO7F+KroBAScpPQ49pSM04JtTWesHkwhcjwmJ+kW
bxC4KCyKWfJqHUqBP9xoQPbCmwMfgZ4EY5nQy66LiuEPi4vbXpJRiGSBLqoEY5b1
GG9WUz1QHPDbpXlz4tdpotXnSI2xlvpYfbo0m0LpXI6jglNRH4mSDDqdqPIWVEGv
bW6H++lBc13MdtEtSsXNwRSqKr9mAbIlSBuw7QgK/0Q/TlK0C8DsBH9miMKkom0J
eMmo66G6D5tTxpH/K201yH99lbImAK1qwZDXrrEHcPBMAlaZKFBCUKpLpt1cY2kD
iEqRvUxlqTmdO79LFIthL/jB4PbluKEwfJoIZ+m2F9+ePlneQSQam2rbLSKEraPH
SK5Lf9QG1MbQQ72JjaiE8YJg6VF+KNnw5WJUAowyomjtBHsA3Cz70rHz0ls0lKQ1
zaY+QMwfvgTzXten5ty9Fx8qOf1cCyE91Zjahx2PWHI2OgAFcsQl08CY3vhsV5iy
lmF0OmXPMgKjnK9noxkcYfBW/e3ASoEovELjM3c8mRvuUQChIUwbjBVV8fBg+kkO
WddvGQ41d31oTuiCNa8e9uLVvDMkPfP6CxEV5bmHa3EY5918oSaCFfAVxeCZfuQR
f89m4Hp5nWCw9bxByBVuDQuhIxjjcR8UaWBhfY4OFIR9Ovua9huFuEePW3yTYMGJ
DXB8+twys+nq4ly8rww7JfBCgJt39R50M5w+HygOm9vd8tLqKgDyicOmWHYHFZnc
Y09Rc2KL7MuJ326AuIdJZjMkdOwax6+Acks2Cp1yXn4qYXSTKtIZqg9iPxbXhjN8
k0HX0xBXwyN5B30/61QomyP0AhQYhQ9Z9tBoWOXL0DwpV9HNLQMBASMMwiEkpyUf
rsQJ5mPiCFTucRf8RTyt/vlMS0Y4UiwQtBAOZjlmCJFgoyqyzHTOYKlqCz6LA/s0
u/r/N8yEZiD1SSD+MbqcDUY6c7sEHuqxeGsDfuwEND3YXasFaV2YmzUj33AdP0Z6
jMmJL6QPYbVOhkbXA+PM3AGP8WhblnH4cbe+WsJ4SXYc8p3jGQRmit5OexXqukPh
iwy4bnWgAxGTDi5mKbt4IXY04zQ/i3IqJg9gLgmaZgroAC2/XEHzMTjel0k3bNxH
TI11aaYq8quGvL2ysuN9FIviWGw4O7MPJuisqBvifc/RI0rOjz02MJTptGTnA7Qx
mhCHOSARfQJNfCPQhB/6I+S8ly/gJm3Y+FKmc0t64HjK4IVbHsfMJ02Z9SsiCSf2
OAHR5MF4yrO04TWWE6a0YwgSG1+v8BBF4+hzbTNt4Q6qhWTidn1Id3JkL58DRcAL
kAAw3Wmtl2KBz007wKsi24rZ4sFoXSKLgw1Y1YpwAh5um9ho0Shoc3AoGzXjRSB0
NoMcz5UxET1wfUEW8oz7UspscFpG7z6wrVyHAgZxm/GX+nHUwqUd/u1ZTaJnsKof
sn9e4QD1/j5skwnwg+ZpSDgECUVR7FYeqMZdR5Hrw1qAZ+dmWDzj3d9ABvytYxF3
aYAeN3ZR3I37e+n69eaWpjX6/oBEWbG4FJdJVzjoh0oYVkVP/IuLNzl4oYSstIfz
mmOR/RUmJesLGYLhOa42wGIYW106QhX37kWrnpDxT2j94o+sBw7WLCq15cRQb9MH
Womg7xTPLC4ek6QehwfA3THbYGLAWmBjcADn3ntLZpKxRptl/hsHO5GMUdQ7YtpI
iVT5zmJAKoRjnoxmgdX35hmOB7V27suCNtOUoEEivBKK1H1qUP8tFWM9vNGCDjn9
IPUQfTllNIpyFgaAjTRVhL/lcx4DCHLQwF4WuZjWefvYvwuBHPsZ9QMiNrQhcXVU
khpOPhGhULJBpaqVfuTusBhsw0h8yGBzPNFbFBGoRB67t8jyGmWX6MPP8zBWE2kx
HdaCUgj7LXWpjil3lRd1enMf4bFDgTYWRPE5ymg+b8hG+Gc+5dImqPhb1JaMo1Yg
VtYvSQxwv+Hs8Wonc7bqNIhzyI2DUc3k5xc+Fx5JGsAzBynrUPkhz5jo2VIbhIjV
MlcfIxw8LakcqYBBYzZNEJMgOWA4i3Gx+V+ghmqeEcDI9ZwYsudJAenkN47Bq+4F
UQ4Iw+tUkiyjYkLJOJg+RIbi1y2z2ha5bzwAV+9uFsgt+fIwx6GWNVOmvcl0JsxA
5ZDy7YPqz5MhUUYrmmf2WwePjSNYRa8+E9dfRgNziKsj36C7xKvp6nK79EJqOruE
wzOHEkwT01wbvYH0cKOye0FqZC60i1pHc00EE6dcr9KGUCEsw6iIT/5rGwyJWAG8
nuJNfe1dpIp0REY3c4NUaj7+gUB9bF5LhxjX3BQDEGWHHUxBmq6DtL//n1umkXhE
baQ00OA/MRMDGOrAUFjrGrUW0w3Ewy7a6BFW+0BlxOjT+hD7Cn79TZEWMwz1DCMh
dskAz7N2WbqhHI+rjEEhje3D2DN3G32UWqXqV/RNGq0ZfQi4XeuyGv//4EQ8zMBY
bOttd4iZcbC6fB6FKmqF6IwzcpRK6y6ONrYci2Pys+i+aD3CpnJWjVM63yoAPMY9
7ENIMfgDRZ8vTLJOYGCiQEtYPnu/o+uKGD4HXeVBExuls/FwcnOe5qdKOGLpmL+0
sHyavxWJ3OPTP3wZLuJsEBUFO3PLMk10ZdbNtqR0PY4I9zR58vtz2wBCZC3Fclgk
0xSgEtDTO9ewUJDEmP+nU8MtYiiozoCsa9YMepiKIPH4QSPsOcgvkc1vSX8EQ+xT
LsPzv2srSlC74gr3+bu7OOgx+CQ54KgBT4fSvAa7r9OScZvswI7qnYx8BV+gUThX
Z5eTFBxiMCWsc8ZGNLe6E8UiVQzq9o788g019xafeotntqB19FBQEfPxH4PzzhSu
cx9w0Vol85EmADm6We5FkIDRtG8EHukjF7mK+HG2TDjTnBlqCPuobsMFVHX/gdKB
O1eay0zoENlDmzAv9HHJ2hwpy26dXfuUKX98a89QMHxRLnDAQYeJ8/nGatvhEn2m
FYhnygvYiX8XFy+MDHz8BnVOV75N2mEX2gcNCvd7KDnyChSGe6dfddjlBTUVdeE4
YwmFDveV67lK9SU0FK8qMTd+8rQN8zgne31VmS+XXxM3SNQokETK0P0W/vsGYrIJ
/nSaKI4a2DbKIVpuaTRWK8sdB/kZlnGDWsDgtg2WGbnpi0oN621X5s8yzfkDgGfi
aqr1HFypGeBkOAhMN6mTk5s55bFgn2TukY5+6zeqQ1UsQfgWDFJr+jBdLev77FkR
w/0ZViNmv60iQnNtAMTiP2ze2XeD/7yVaZk6zVD6rjm84C499yRKRYqhirgk8hlq
w3PsurCWV4pkeuJH6Q7MMn3cvft4hAjtQfeY7zM3/JJjetTq6dcJr7zrtAVyiZGF
LAf/kkLIeL4ybIwESd5YWrBZ9v3uuFZRorrBFh0i7wT8xqZgm8oCVxEfkkeSAetp
KxxIR+J9PXIgfPsZiyhOyc6W6s96niB55EV+XeqzuAVKBKYS9hhPtWW2b1Beh1uM
bsBNnKac1gK9WVDRk+4bOFXI63DE4/GfUNoBX4UGY/tAKlch5vOAxSAMRC9DtnjS
K7265YOoVrbYm9ramQRGgEW8rtzsMdRCieITBBVo7SnK89CetKXbX8lAJ0tMq4hB
MDlujcQl048EMOOYy4ucwYAcOZG3jSkqlapO7+6NRQdQWdTm2WXCcJM/C3khNvIq
jSAmRdRkrKWfTXNHYP6kfaq12f/++lXMXvWpJQb3Dkfo55xu/LxEL7JRXfo8+yXh
obd0+oJbYB+wIJ3i85zL9mEYrSCKlEx02emPFeFZT6VFmBRhq6oqMFLAznSRsuAA
uYkNQvLF5/aTaMda00v+I50Qm/IjAqgjt22F1Wmel9BpPiXkMaiZhEsBY0//LeHq
KpNtGdH/l0ChKjX/+2JZAVZNC/IL+4Apd1GWJVyEGpaL7RafBmz+hO259eajFnmg
e8GeGRfS+3hmwEFjHpNnBvlTlqI3EkqZO0Ir9gtF1beWE9aovHVjJI3n6qRDHS7j
DQpSKIwEvnKs6hK1jHJGK44Qo00oRLn/x2qLnPA7v1l2OnQwJ+L7DyvFvRSfCXSG
+DklXHreJ1CotD++8WTK7GYrhan53tAi3E5dr111nZ8VsyKksGBrdAAyktQ5GkHk
U7saM5xexNC8XT4ztSoA8POQneAVExddZpfO807whnlh/0S7Hm8QL6KJ9i0GxmHN
4n01DeMkZrW4YEBOqrtJinCfv1mfhQxk8YWVuTz1n5Iuz1fPSRsl/2+ocjvmd7dD
GxEFbJvIeiqOBg7M7BLwOugg1zS9Lmb+HixG+ePjM3yZ+DYF7gWtyvSJgMR61NlD
mstAz35o5/PowYCDV4OYEaTw5gnBLBI/16atAhBMUNJ0RpVrKWfCwC7wubAhpFgV
ZbPJxfaJHPJo1HDqPkYmxvOlMbiVFGLsMcwNDe/m2EH/c26Dhw20qdLdPyEdOiMq
61LO6Q/7s9ug9GoEdkEsheWyWeRy+r70cDutcnRrEPYI1YsqYZnRO+BZKCa2l2O9
1R3NcpL7YLpaiXe9pVah28ope8DwLy+UTI1AqNLvGJcxjrmoRygbYdxzLM5I/pI+
e/3VzskqBxe8Likrvv5KJB4Q0kgdj9F2kNTq0xYjHY2LS2E0Du4cZxOiT/rPbn1P
X3F54ovRyyRQ/76LZXPaNlCi78lczQWjklbc4tKO78KK65liPiNjVPGwWivX9kkx
H+ZXUp+7+Zw+clENzxklpz94y+u/ezGLk4+oTlZ1a3paRb8tm1K/N+oYr9WPS2es
S/q6j4RguK1zcWVDvf/PwDsVG31MO4zQNrX7ePAz0LVZ8M0s8rkCts8AbvyGzyWX
e4/FNY3LpUj0CHkdx9C0JS6DjpVusqVin0WX/c4XjCALok1cjEM/Vdk/fiD4a0XD
oClZuuwZ+Siko9Th8YtDuji8Wcex78W+Ce+DUrxaYUivwY7FMs+mLwbdem6s72E4
XTOtSOkvscyt23Rz/set0GtGq7Thy63CScc/kGaxv2aPEaSliiP+5HH309AHeERM
SH3bTLzY8Kw1Gypr50a2Xu+FGtjERKCFXENPKdLr/CtA86JBPoqbdshLIUyQBGyR
bI3VV7hi5xK6gApo6kO3TbQ0hmxJbUUbNvdvRh0CCPHt9zhOmZeC022RzpymFkqU
aUSxvomCo8CdUdHmlRjQNG1WNUyMDNH03kkCQZVk5KfqlsUhcjgVZUZKUQDAVPT2
WTroELeLdYu/YelkWGZ22zVsXBfhGARnZyk6LpIcSzAEmJJ1Q2e7A4ut3Ok+9Nhk
6LiLI+IPGv43EL2tdD36wKVomLXaYIc3f0CQ5V3fxQMtceJeAR5PQeQJSxkAee/B
saQGl81kQDYK16EmmXhH3utBsERjagyDSkkURR9cMHVWHSypgYzuWAGJbMaeQqpx
vinRsfFeNzh75rpS6RoIBLKXWTUxZ4ssMIEBh5GQ5Epg/ebBh9nAdnjdsRanlr62
NjF/hbqOIgyeFGvwimz33Nj9hhSlg+dbMc7jxm/rtZoiKpyC70+xa7kCrwYOKuh9
zQ37+u7cVmaTzR7I0kzCkEayZE/oFYphwDs4cpxmUvAz2lRoWIgUfQr3Bhaoxrb+
wqc0GyrAavepldiwskAGvf/uLCIU/hvA/lqh/o5qyyfC43bblD6q/l+Ta86YWU1z
UFpUG/j4hKKZdkEZTVCi5dxXIWqZVA0V1WSbB3veUy/2swqH7Y/9WHA0jL0KzAvL
UZYAKpnN63rOZisRwAGt5tTQsdp+aUqvsJQD6x0OEfRR+rwSg/JhXM2mCg/uFqcs
o2eDOlzhby7FzddxsiK3j7hWEKAJwtTT2wsK6Mg6RXiTBMzbpNMGytfX/ZI5Pmnf
b+u3Lir+LoqcEAMHFeRKgi3vxGidV7aWgTmi1jdnShgJtRe8ZB44dGFuzWdkaWFR
S6HhGj6tgg+GnC4mK+2BcmvKqwEUpyacmqC6sHDRX00qZzOVFxFiphOpRaodbqoR
fN3GzvLkOzEp9FZ5Os9UUyn0AKkc7kg3ishYd8dVAZS75iRLQYyul6o+DlBp5Ay1
0rDdbkRqVSn78DRjqcq9ZRkyoo0CWTqKolofziX7OQTSaAdMp9CPJAsWD9iMemip
25XaGs0b5mtDqKAzSjHUid9IGkrO9Ijv2m8XhITyWIwEIWDAeTGAKCRxZ/kaJxp8
b700Ljp07Wpr7Lu5Zi5ce/nqzvIHErFH+H4lAV/I/HUzJyBWXvwuTLYXuAa/RQm9
9Yhcl6yCTCwhiV9ag6U1SzyqFbxBukx22yuwzEoTc8P3pnOxdy1veYt1TksZ9XRJ
EfNEZORi1e9D99jUm1qtAtBW54cVzg9du1b9UwEjDjqDVSzNBWkuVQqvHlnHzTBa
DOYNyzc0OBXBJRzyoKa4FMM4J5AAmi6URju5lpYiIU42o1WOd101P+m2i876100Z
/QgESI5s3fSejoDBF+hO4JViRPov3n20tsc1qvvnoCj0xahsucYP41U1nlFTZclg
I6MdUL+/dAP4hWutr0OpfF4Dq9+MEeqAyff4NDj0mZzCs5UwbvDn0dbwzdq8PHSa
6uNY0dihltSTFmMMbWaIM1YwR9o/0i5IS0/w3sLBhmA+nXRZ0vVym6lniafGfonJ
hUXD2GDXopyXDk2yHx4byMAT29D2Zk+zYs/Vz5nTtElKUQdnqDaxK9omBs434J6X
Oi8fRaWTvB6QmZ8u/wd+/v53ssnw60SctUo0UFSfWbVgZqrimrtf1M0HZ9d6UW9y
sjE9IgHxtCLxW2P0uiLatrcxO9nRuLimNo+9WsEewWv6qeEV2+ErcCWbr6JC7CZW
lALqjEbmgwNrS1B40UjNEHgcIQePx3kkaieVR1qXCZffhYOycKyu3hz5xy0fCaLp
kqTZYgSOupHzx4+09HQHFjaf1i5Kt4qHUS8VsFiTCW1+U0wwjIRXUeScC5snXAdD
hdTEvsFz0EuWOrfqTD1QZTaB0mzOWXJlbfY9QnAzZtD5L7ALOGhhpQeINJ7UvaFe
Cn9TStUS+s8KDY5xbBNnQ9XNFnv66GdT5+moNm3s6eESuNI7vIEoUqVyFsuowbhL
QDuNbjHNAd/bdmrFgfl1KNkswap0bI1f0V8bazeTc4qULzk2lJ79zzAuaos/Un3L
cPEIoDIzvsAlF2eK59UDZkW41Aic//5PAVuWkETZN3AmK8Fszos7EIElZzHVnbzV
bABrfVlIF+E40LVXyVpSAP7WmpoTRk8E337k0vwUiilA2APBGrFE6EL13zhBQOSL
M58EVT1GIWZ61FLL4H9jzT7afHkEgDfwi/nC2Cf9PlXgVy4KMpx/C38ux4ZdQ6UM
v+AhSiwrtV9AcBTp4Kl8oUxKfUYNAB2kmQGZiTWDTYGrH1+wIbMXMVCCHLM22X64
jnVqqiPSuttzrzw+qgpmx3I/GThZI+XSlczsX41JpyH2trX6bteW1nK3xXRgedNs
skqB3nkRNQYSsqNDmgmtNlquYCdMu3DtXPG1LWbSPVIu+UhseajL+8EkbM1joP7q
y9TeNjHBawFo3EafpxbhyPDTAiZZKauVHPydEjAnMcwuAdTSAUhkGSyHcaIeKzBl
psAg8AJVhOy57ZlPwfl5yJ97ujA5LCbt99FABOy4LC1DAprUhefYxUO97MNY460U
pJ/iSoBVZoTO7aKrEkJAXW3cJyO7oX8LiMVBmYW++FFbaUfIIHTPyJO6OmjBN1ue
KA/dOsRMwQ2V45QJl3QZJTsPOQVoj7DDCs8biDvZh+5j30wkzQgcrwQThhGo6ahB
4wcD8ErZBYasv97jtMpC1QChV4QGBq6pDwkWErz3m3pUF6dzVT2gryO64w4UhiOh
0f1QIG0xC03Z8+KzR0KVU0VijnEvii7XgXuJy9mJR1TfcmmdSMErJPOdggsFrXwZ
pLcnmCTWpoMAHM7jd94KxXXu6Ek3IzZ9md6CRCsn5wHcXcWsQpabNxN9zkN6ZcHV
CqmEDA5STlBi9r8WtQfPIPTKZSY2Gh8ZbFdnwDQdQ+DwSD91sx93e7ax4+aDFgZC
rB5X/hdAvq1cn/VevnbVNpsz6JdvZuKx03b+4ej8qgBnAhDAoxdCh8/e2BuU+P5Q
srzVotu6PM7hV3MGiosSvRDjWQgCjjMdHE/lHzy8hlgu8jzcNtLKH32x12eca0kX
5cs01oTUityCFI8vOtLN+P+qMHCe7wXHHN9Gfnc/Ly+3yFCch/nGrC5SESfspLf3
k00oPW25S77/1OW/4qrYPY5wd631pXXyWDxBILC+D/AnYED3BW2Cz9Ak2kFtCELU
TgqXzUe8SINhHv7K9RKZWzy3sgokrdjpSsvy2r6EvNCzUUh+l9KnlU8JgLzCxMsR
yB/JDwEJjB2/B1nyXlDnYmtTxbQU30npCSgvU9m2Sp7kjLXUkDUJsdc1UC9Ic3LN
WD6s9fWoOzR65lk4Q5pz1cX5/yL4zW1EGbUpXj6QlGv/TfmKnnWZ2j6jRmIQ1zE/
LM+Mgx73Qkhenoc5YFzcIPE2WMohrXjSbp0ucKXXiW3XmVNQ4EN7Ajd+uOVaxLuU
aMZ8p/sC4hYlHZjxpC0nubbvwyNWS3296fxdWkOZ6WNJehTswJxyr7Hlpw5YBomG
EiHGaI9IGbXHH9pKFzgtel6FlMnMzsjolJTJ/w45oiq1YeRe7Uacs4bU7xuNPY1j
442F48Ak3AbNxj/LU5NxzmVLkKo6Pf4YI3hqyPy6M2m59HXPywOAZh9wyF42ssU8
6zLgLAAQmpSkjhZPadLc+hz/TqWinmEpX7Khe00pTwj6QOsbq2h6tXhPzC8Pl1HU
PbMcDzPdLYk3A8H22/EUldS0Bp47UOAu1Tbg6QnVqGIlE5sWaLqqAnPRWoa28egy
/RatC08Dx5PWjy/dqr5OPSmmCteUP3669sHieDbCiy9+Cz6r3PuRdskT2EgAy5nk
T9lK5A80cP468BfkCrPWeaq4YZNFl+PWLvmZapo9fWwN09bSLxKrhsfiDPv3sgt8
gK90a9Z0ooeajZseFpz2Q+SS8Qmd8cI9vcjd9NyXTOW0UiODsuTni0/RZvqMurgC
iYIAfy1dd3ELj773BDRZzktnhQNMTqAhsnn1lNf9vrpeCQ95x+N6/x5zFpJyRIoh
uS6temlPAGsuKGmyNN/P9bS5/yxMv63R12bwby7iiIl7D0VtaMNj0D7m9DdqdQgj
oo78e3erkTQZCvdyNcy1h2NY2X8tynjMXe0rstZmZ0xuqQE51V6kGj7nCpcrPbST
sTpDf3zXvBZqMiQkZxQaYNGToPF/gHmkf06sw0Zw3npxti5ZYqGzJs2DN+3lgxVH
cyNPiCemGEII5xM7EJbKz9pw3YhJNKOziTWWEH8llPKy+D2/rjnLZEhMyOlB1jwf
Cch9YIU5nisjVbItbaGYDxLXwbFgGZ3lFqPv0PvVLnBz3sI7Wnkyye4K7SFt8g2W
tq+YfM542+kIb8qfpQFjWe2sLrBT2DPo3BIHR29oMnNyc7q6OnogOqNEvebpRsSs
VxiO6hvE4+fMTVNdhqFdIDdm8gXDuct4rQN3P1PtbWfhcJ332oMbIsl3AO5yrYU0
Y3YHiJDeeOKnJZec+DUcFl9eUa6WAWvMecjZ1Fdf+Uzgf2Gaw6PYreK5VEdK9FNL
p7yV/L0RTWhVvHKZBLFfNr6WvbnaUk/LLiBNd4U122K6vTh3vHWvo7EtZRwnWzdQ
V+PsG9lMN+x6F3GyWpAHGJ3L/VEBsbiyXsP+m7cRn5YxY8Z9W7tl++ulq6zOPPdO
uw0twFVk4+AUgt8s7qTwU18d3DOlhTvIN5mtpbjRWOJjg5s5m9cto2N7cKOB6WUv
VgzPGZGQsstCn1Q+CGLOJIpwIWVhb8BWYKf0DT+qL+qp++yRhF1fOb9x/I+1fFLr
oMHvygbkIYc2XPry1cDsZXb4UalfMEbQsmYJo5Xrme9sq1Fst+kbPMnpm+5RGcZP
g7UBOkLXZwxumVlRaHyCL39w+O3Wr9WohUoQtzxA7Kk=
`protect END_PROTECTED
