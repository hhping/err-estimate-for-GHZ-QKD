`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJy7W8gm4hW/YptcOVjUlyS9LQ0EfPeLzoq6uZ1+x3+ghzjh5/EDYNFdXM/EjnuF
2/nkvurbjUEmidFRzTyG7tEXoRYu3GUO1vka9vobpkAtwBQl/ToedLm5sp6X0jrN
PAv2HX60iArpxCO9g4p3l6rPzp8KeqEiAUMKtqFyUHujxQe6t2+7VDz0lkmLnQoR
pTfYQFRSaeJsoKBJzz2CNZemHBHqQ8355X6qW0WEs3gKlvVx22M3dBQgBLyUQ8xL
3NJxdSV0xNh1dsemY1jQed86OpqcyyT55r6cg9PJkuRiyJvnGN+GqZrYWUZQAqby
sDUbPLJw21HAO8/E1snylXc9ioe28Dp3bGjFQmCDLh9pUfpBtZMFm22rpwhN62kz
N6w7ndKXXNF65jQKPVwo4hphsPhLtr8y8XfJ3LtCESHcVMCGfs0QZdv+owSxHQtY
Yxi6ycCgsZTkaQ7jmNexXu1FMmhwOnUT+9VY6OK08Yb0CEafsvMcusyFvWiDXrW0
Gv4L+iW8pt/ssRNyU4PYXYyzFTLxeRwqgbGliWlnVuFeiVZdX5fFV8EC5gAOWUBI
YcYvb20RKWyhesTGr7duc3ghKioc83TFDY7QXhXHpasx/G4+Vzc57WMPaqbfVTh5
GLOukIHAnZYijiLCul1rDD2h1yxtXifqtjfpkKl8bWhwP3W4hyjqvq/ylwt2Lf1P
QWzaXGVZuGCCCZlOlYpQGl4Wdar+ngWQekH1EMB3hac56/K6NrEyKpUBbnuMHq1j
4Jy0dZ81H1u8WAkeW6tQ3aJC9dvY/UuO3gyn2Z86npP6GPvMjYBsVq8TM680bbUe
H007R4Oi+hfBBalFIwRe4ASmDhUU7/ZzplPtgmwLl8p11dwkvV2CdfQcstRQynIv
oju/uzjHouQQX+72HkAmb/3Z2c/7LvNvC8JUpMBDqY5375WcAqzybTv90tXEfip9
nU2+HmtnqZhQwLGEFSFGPJJvSvPh3m83nidu4ep87JxsOFG87c5lGz9deHh4cO7j
X5wwFcSxRtok4lNWKEGdBCBT0hhIvAKKt5sVmLxLhSZtq9PXZ4nyOFM9PG5ftp5f
WmM640LlThuJy27AXPOGBaPe9af4APdwDUs0eaHaxVC9N8/Kt/BLyWqY28u1Ho9M
kyOokDeDqE4/CaAf0Ss9BUoibOv38IGrFjVqB0ysgEfYvTCG4S/a//wsve6JkyH4
m2CV6te+5xqgRt5zARAUTEZxsXM+kCzzO25zS5F8kV8jhvuSs0Si0wZ0wFlUU5PJ
tNhGmE/cMzurSTanu4swEwa4grUZ50ugeZzEx1edeejQlcixtIqUFYtDx5mW0hLm
qmtKDi7y1q15jYpouTy1a4/ZyVej7wRr1BdssGhx7s8sinje7EEVIH7YGY0MXG4E
iWo5yuhMyUKd1CMdQtyWfhtH+luR+MbBh1whK0NlepIlPdgPbOc2kR2iduL2GnJw
ESUxSSzKam+xuMwD0Yxs4DArKvjqn8ze/wMo8Y5/J0UkFM/+i4tUPb9llF7mHlU4
VCBGbOcZq7dL8dRyyp3JrgJEAryN8fAC9NjBaXibbxBb2lYqxI3saWbfb8nFnyiA
TsmkmRwnS+Isvvgg6sAHAcmG3Z9LfNDZF/2JVv2ym+qdO1yLwfLFbuXoVVZRNIhh
peYUr2KTaJ0fpfrleDO3ZvvGjmWnopppCNjOEcwuSOh/8OdVwDKeOxR+ds2Kajgc
klItw1IG+2CXJSrGPoS7kIim5DYg9w8C6ykE8dRn0nUA6ogcUhFMYPDh155A9jE6
73qtaZ39k5qSYvNzIXP8xwHJlYScf2Dhc86oL8S6+N3BrKwme/gWpIJjLIWhTIhR
H2lNyasVm7BRKdyPcWgl40OB2qM6IntiSEA5ZQWjFeQ2pqaIL4OSmQ7ZIFwhCOiT
NFtq5RkqH4exTBlWrdaykMf3R6IY/ghDehVcKvRSIA+MgBsox23ZCifF7A9n4ssx
ly80+H2xcmJTXD0dbiKwMH9pJ93fjewT/Z7ImnGRM/JlRGzKjLbaaLuT7TqmiyGr
FCu0GFuOlwvR/OEVOV5Rx9fmARpHaQKM0PabHltFYdmN/pRpDsZGkE1cZy8C6Xez
AdXtn+cJ6EaQLGefa+FDF7Srd2In2y0u9kTh1rgskpZW2Y0pYyHmHwd5rH895kjr
pKWdo8c4kAMTwpnF6aqDfcHV5WRNqMkQNWTu0TE0iKXGy2KlpA3JpwUnlusNDtaz
cWKrJ5B5PntsX0geO3iYxIuqoGZOt+oxAmt3d9i5H8Rkabp7D8zFYyO6fyyDZMiU
ba9gPu/UIt9TqEOi1/5aJo2tKLVRxPB/P8QSXP91lyj1OxYYvhW0E63oySuIDGTN
qwx2/5EITiZCRkp/qTlSWgukjg15kqPKLadxDKJN9JWgwagzf3VFe1AlHPuAufEw
dJelItMI+XaNKdWVKhCm2WWzkeGwgw60WSewF1HcQpkel/GlwL8z2ou7fH65quFq
s/mKCfQMgdZErz9tCIXnM/i0ynibT0oGjk7QUQVxZgJr6lDZ4XYqlENd/B1nzEcE
2LPkEQ5atcgUBEo1vtcV6E3Uj3nrYXEciT8DjS8ZcUcBUSfRnv39yamxrPbeDe5H
neBBNpZCGoYF7VM3HS6vx6SRqhicIcAUBIop5kZuXacwMs/qz5X2E09gQtHu1o6d
ykBGVOgA8fq8ijtyTQISvB09qaelwuNnY7x/nzJ8b8mN/0cCgkdLsweAidASUFqd
9diRaNFV2m7qUImX5CdmIlG1kGidu0gUzTPkLl/fdCyjG/nmqvrMB420cogkC0XJ
/AVtGQ5aXM2dyMQeIiLvaItzPWIGkVScG60mVS32lMXTpm1aJXF+0q8B8m4RBpta
HopzfClgftRCY46iPsqUwKlB3RfZ+OVuEHL78Padu/lwUWJnJ2eL0/tYs8179S/P
PIWozBkPX6b8qw/Z3qTITJ0KZcRf+bH1sTXD+ZrXDtqM9RmfT72LHE5o7A89pz6H
lHsYJcJBja8CrXMOe/cDw6nqmwkkaXZ213tQejoMwTk9Z5gtAvYkF9rFFaBpb/pZ
RZ3MZSCOW7U5KnEqdsjRBgc+7kPtBjtHoKsMGrx3tI1ReKH5cCid8QbuWZ8ob5M9
OFWUH1NkX3M2za/nHsyMWE8fMM2Q+22AHF9D0AKC4B3qqJv8rMpd84HcBNEBlN+l
M++ADI5jduItFgmm2j6zCHSlegofoTBcy5yKAg/S/stffBb/LOKwu+1m6KkPosOX
N1xaWg8gL/+IV99ldx1kZPLLkeqWsPsGhkzch4M5o1mGiOVRuPUvaVhuCyKxmL1M
jsYNPLo1w0tyjmWAH3rnur/a1yh2mkL8XiWOT4qOwjBaNMxlsx8W0hWZ8VJTaVSO
81drqBgAFHEQwad3MEhWMf2p5a3idjjoyL8gV8rkjqWIAjvSsUGEp7fwiUDIpfzA
skWdJWIRI3eGVJimAYmKu7x75SNqvsuiqIh57o2BxLsSWRElsiJaviVlItQ/JkX4
ZC8qHB3jQbN2Wl72KeI25KAbi4G02Rd29Uhc9N3dZrdAT5phFWLf3jbl/5OgmiyA
cBE7HZA8F7HKjurePbe79uGn9nXQPwyU1w6DLL/h9bh2DrATmyQEihAmglZmQc30
1hMO2Jxtn9BV5NrhfgZ2+j+Fi2NhtUs3PtiHHjVUbRMtuKUN0+jIwy/EmIpCCE+4
3IUOqRKfM2qOSuIaFsD4A8IYxuWNyWF+7yRURdmpKdqkXU0syWedTOSNxpTKhiVH
VszrBCMc+MdTXOawZ607HwDF8M//M4Ey8tU7qFDTFt9mn2cZvNXDHGTEfKW2bzsz
ZBBdFvYtHHtk7Orj1s6Ou7twgTEQN73ZwyAH3IVWUrsq3ucJFgLBq0GGmc9Sx3Bb
uCB2CdK+3skiKiGW6bCMmJMHZGWXhTJ5g0+d2Ejr41QiMFFtRZMdlTW6uUJDJbKX
8mYa7Ik52xikyNgr1icr1jkzbT0u7oPvFeeSLpqZ+PzBVpUbr0Asw8sJcsrBDj3p
GvejryKH0HbKjgCp5ShGW6yVuv6TZRSkSqqu0bMyGCHtpTDJP+IKMUDiZHrZpSyK
jf7Mf199wS0zS8PEkIl1vGUQNEfk+PB3kbkgtSWguyEoK+u/tFDLDVLReiwBv4hi
0sGoWfeG9gkpAP6ZTQywJOEfyhRjjPb2wTBWisAX0Oia6VLUZdaIkbe4VPbxnOcW
Xbx4MVBkE9iYfFuUSwOJVNLH4KFo7nuH1hycC9UP8Xff4B0OuKq8d58lfn297dWX
/S+fvWvcFCwERXYzaNVNV1ocFzv0qKNmYrNgYl0S6LpnRytonqtBICiqNeLg2aY1
TWSi5skNJ2PKlUWHNF3DrjH15ZtB/SAclCVGQCNAk8EPmjmeNAzJW5SYdvoYtpTb
`protect END_PROTECTED
