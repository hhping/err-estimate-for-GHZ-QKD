`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUJYtI5PrONqzH70FtTiDUQ6TkdA98YZ1qEQ4pm6cA/V8laWiDtaObl6gr6YLr8h
uKvEwsJgSO5sCKqF8UTv5IBHXo82VXme0LokkEJksmstPmaTH5HRvAoDw4CUSsQf
d98I2i9GMVpsIUEQQwgtfSS7r9Dc0GudjIXT3APP0a4Ay+K+Df5mXGoeEGCd2dDt
VLKXllBJHwsCm+awJkVdL14+llfR9wZF1H2lfU1218q9HFyIHjLQFfi3MtrVwpnx
0eNz5e+KJjIo3UkxQKJYp4kiqY3LoaXLMgN3J+DQGpXMT6ESIW7vjIpvu/FyY1Xu
hmgPObqOdKjGLMI5AAfh66UY2Ch3XAQoA2Muc++wwUI5AT9lbkBpm8++j4AoUOJ5
yXyaKDdRjyAhvvTJjGux1AwbHMp0nbmyXQ4zh9psscF7ecbX/ifFWUPf25O539SN
Vc1GibZddrYUNGmYOh2R5jT552lOYy0k7EWVcZC2BzmvY7I3uvsvPuurnb7u3Mq0
u4dl6ROJBf8fZcDWKbbOgw==
`protect END_PROTECTED
