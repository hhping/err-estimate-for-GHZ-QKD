`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kUMzeHAleYuspAAfZ9F1nS6RXaMIQFcIwliE0YPOU8Dq9tAgxbBdDR4PF81BxU4J
y1nwjsBuOvS0YqORQV1Fgw3FovDxwbxXBgzM/nbNmPqbjoD7xL1y/DGUOMDwbipv
6BAmz7l3uMrFMEuFfoYRPSFh/2UywD5aUKPUZSZKaRpUMIRq/TkaQkq6ZjJH/BcC
hN9tcD0J2uFdAn/D7gDzh3C8RMAmZXbPvZzN/0xMQcNy/ZC1nfIETS4pEdAy3wWs
CTGanSHAa9CG16duepoi/6VSd9QTLLBX80l/m51+V3WlBh5rwg4Vr/wNHdnX364c
BnBIhd/a92Y1hF+7KztP0b5nDJFwcDAipSrSKsfdxerDKLN6Am+lJzkvPrD9I2J3
ZfZQs0Ql+OBjX9BIAPKcx3u4EuFmXUrDKNJP4FUkXajR2TIGvIUiK0vkwOAuEEKI
SGPlNxpy/kBoFUB+nCa30UpE26CC13e2T/L6Pu8dofhtOcqKpJaI1SKh4NSwAKsV
UI2umsbGQDh9UwC6VJYXzVyNm6Mwv6gVdcMfPq9Y/Es+yZjapXvgQB3TiAwWy63v
QEcLc69DpXRnyaLLcK8w7kyPIsrExg4iY0x2ps9w2bX6BuJ3mZQmmrxtK5PJ5Ozp
fMzBkmAavAHMCMBef1tsXCJSiDqFrmY4/5eRzQcVbIFqF+NiAqsaYCtt7MSkCri2
AGlnftSUkVvFu2D4JZa0+3Pp2euq1RoCeRu6FXkpj7WlJA7L9yyxJtHFnO/jrszq
jUXXn2x5+IB5YSgIUqU+XuDTQlnV7+g9o35XVGAAIeShL0ECkO8cqVsSNzwB+xVD
7iPQ2dFjsONDRAMNwCBLGeAYNecqE1M1FjxPyI8FG5Mu0/tIyKQ0+07CRZ92HNiD
ak/FYv7suVf71LeG7UlyfS+F7PbwKqyOgUpULFTSG2z9Mc/xdNOR6g4qVM24UTgH
HlRiezJYGLOtn7EQCvDl0eyyi0I3yr+8owwFj0P0XdGj0K426PyD3og+yw2GRwvi
uaerxQ5xzVIKDD1zBZkcF/FwmTbuaqKgdB4wGuZkrFMjW+AhCY69bNLvQNrCYYuH
P3jMvCLIUJVxRcIb2ZcLk5FPSOZjcWaBr22basoj/840Odr25wdrHYjIwb2e9Lfh
17p57MoC0GCuIDlRV5S4wzU8j6Hj/6lNQ2HwhIchckeKQ2ZlaEBPXA5J7PlhqnZG
s9QWUMhs3ncqBSasI5HmXEsZgdPqKsPL26qQ8CUnRsE8GheHwrgtlZlrwJ67wJiZ
MbjpE8dkJ93P5knDE2rsD2Bj1g/k3yWy6QqkgAdL3lsB7s0No3/f7im8HFfXxheJ
q2qKNV6jIgDcTm3kwlQfy5Msc0WszlQs+S5/aU7Ypv36v2WpIo4Cq/iWYQ6zfTi9
e2P5zzoVu7GjjqAAWkIvfNh2CdDPuIYNCmMa37rbdKpXlT+qweWSbLEkgKgZzoiP
3UkJpc9S4/Oyjd3FZEt46oH2BKfE3/nEsfqRmXoSLiNfILjbFGUzTzlYP9TCEW1B
RYNb5EBhNAWpW2dNpX3SiyZtP7+2pviHYx7HmIyz9tEIznOE1NlpfzjUP92kvATA
dV5/xg6H4G5TgWwhQ2O06R0WCqDee7KNI+iCMMg1lGEjXO7BIheK8U8NUZmtsTjC
exD0MYGuMv14BULvV/XIBk0geOG5VQAi5kBhjqwFVWjbhdKqq2wv1oINg0NZ5YhJ
o7Bwkq4w4Sw52EYY5jYr53hTiaGLsZnQf81dOnXsAV8/72bWTqwvtF6WURyAsFO6
+Yks0nZ+6vJC4Bse0QKgVJR45w0MeHCKkStT8Mn3U2QwvcYX6atiPsA8k3oyHRiM
la6KBgox5JeN5rQOP2CL+G09EghKpRLJHHyljcz1BirQc/wNKhDvh/Ugb8N51gg+
hQ7fQ6Z9uB6oi4JMS77utqAGmf/Fnn7DxpZsuApzf+pqCjfdAZalDaHLCipoudGt
ex5zKt/yM0L+hRS3IxG74oAR0MFRPT5JfcjYnjjrr3+nrUr9FL/dcszsyihFUg7O
r3u+qG5JF4PBi6Mu0ObNd5eH8eprhgVKralRvbVRPmuK287ogZuQ16XsmJGMlleD
8edU+bzG3PjrbwqMWQDU84XucIObY+hMsIGBnmwmLGcp+e7AqsTvfjnp1YiA4D/d
DKMsvWFc/Rh0SgGFlZu1hcfvWYyNFJ5VGMtj2lIfMTnBVNFPmEtPi/laoUphsVk/
H7ASsDQ2tn/7DaywTecOFnlN5DsXYqDIKry6gdz4Q8zjrTsD5b5yM14/x7r1GmGP
kkImtvOZsNr6c11XKsGnLXFGvde4dCCFWDX33F9WnMm6FcuI9TPZzCmhFkpViOUg
LP5zYfPB83LfS7GQL6s+zvfQ7ecL5gnwoOXvYA3JObXzleJXcPiymFwAiZnOt9NN
GVccyL8OMQ25ARcjbGRQwUVIm4YIgH11+rkzgVSQfbjUuGFkHxGrfHTahT51l87D
36jtWbBEJQHYZBJ3+NY60i0V0wGB37PY8skOWRG+99KgsoUs3sxt1jULcdnKjNuo
t7eWBDT1u32Xow9NUY8RP0dQlH7eXotADpSmJp+je6Ezx2vjrIXsSmm6sqqKk4Fk
mYJkgWtU/FzAp39g5udQJGN13IW2ZAI2DOUs4h3ly4zlAmK0OrdwxdcrE6ZPDy2z
K9O6bcZ0ZUg7IIojEeGMLC4yBdAFc8v/FuaSSgjpDPLVQJr9JdcqRI5ugLn9LEiZ
bT4Ue1iLqrbKCTAPfJ3arjIHyh3yxOJvS7rKPT0F0NSBKkP0kxeJJj7o2bJuvrj4
PVENbjAMaymHI2r2+TDuHMAYIU8RMXl4qlUtF5VV2scFqhX9Cd8drw5NyMuem0jd
xy9s2l7ZvAmYGFGTxqfbJli0LKQCCY6UvUFBm9qNc0Sx5pHLcuvOEwuHR7P3UROf
fnQP1c1HlvKWBvY9MA/O2XqeCv7F13NDJB70IQg8wdwkv6gyBy1gIM0cA1YCmqA3
OWGNFjWzT01/vICWcvKG92YpLlF4kVo2O24k8a6duhc1avV3Smxr9bYouWCm+ot+
NEuRsMgUU738s8Xgr3WUs/2cGKlTY70JZ2foWsQM/b/woxdS8M5X5rDoM+t16yke
+mLG31UEMVhR6dmr8fiM6h6U69GD6RJxBNW5KOamFcPqUvW4pR5MHyegSl3Ppjvy
T4yI5u0CfXXILFtq1Dq9L7pb+mm+cCrjNy40ovhFYqY71U4UAf1/WYT5jY5enJ/1
FhXbeg+dRriCZlPQgXFmJisKXRiNepyD1JpbGri/AyoOxyfELAV4C2SCpjRbxty7
YXapdv5EORZPIw0+Z/7Qynp8srSQfSxgj8p/ASjQW6EF8D2/ecQ55xneXAiXBJSt
6slcgJep3fbjYkl2miRDIphlVihW0+FZ1IxgNV0oyjlsNJ4dRxiH2ZAJXslPCgHI
vjsSvXWepacVm0S0uzeEYo09BwwhDt85ClMMgNOf9uR23zeU8/EpFnPIDF71ItWb
Zhc68qbQqMKSBHoWoBPjHcb47YCjY+Kw/m9Qou5OQ8fzxfBB636rrcwyYbDAHtDh
FGWzvPuFKA4Z75UgBNzwntJGnQBvpL+3Fje+XwPkDRkNUDlzY8BkztX03hTBlrm7
LraddNaLaJgjGb1Clw5zPnx5BasYMyVSIsvXMa2GXJ5RV4GKVD5d2vk1nXrJuOEP
5FA3kp8AVL1XXdMGh/LaRwoAcqCoZbYauNReBVfmpvOlozHVoWtdvyMbXevSb0fL
SbHAdFAFZGOvFPFpgjpffoA78n5oqeqEzAWo1W8yGN6KCWn2t2tMSQNxtQ1snif4
ZmsttEOt5fccsQZw00NTh82WnSiCOHnhaJiLi9d1KKYCBcLJZc7lsP9ruaQaOOoz
77QzrPj50b9iSZFfcWZDgHXbe2PtMR1he+FV7f48kz1O+jcwsXEg62cKy9B29N6v
4j9BJVoR8XFJ9eg6HxekKyKxhNtB3oUsLucP3NHeHRS8PSY/tfStzB+PMHb9h4TM
v1Mr1xqlnnTDkva1IdD6wcBToQfy0PxSfuE2qjs75uoVWuVkvTdlIxSIgmJFLGTK
2uQ1dCfCIGCOWO9G5LOZyrAP4r/UUvtOjCStiUMoFhzI/uKhQ78pFBdHNa0gcB5r
7th7WPk8jNm+8NN9oEDR4ETdJAFmvt1hL68y44p2Tcnjd/ky2jeEpEPl0ZaBXcFT
6pmeHeTGFwejwSVQrXN7Sg8TAa9kRs5QdL2MWCK8fpC84Aieb9uVnfjbtwNc1e2F
X+ksY64SOr/Mc7d2lb4dQUVlH6+9P0Kdvj0oB4VXGvC4tXj0GrEiClZIFMIHhx9M
NbVCGNzxHau9EWHMlQxbslpxt+AHf/bVd+/pPwN01gEwNlT1JivAHhtdGmZQh4Vk
LmH3xuxWWKixoJweheRhuV7AwA5gW1IyEKMpE8GU1ExPOml9piPjVeTkoHNMUI+H
/jsyQjJek/SEMdUuVsTmat1ZkIN3CEvN9UONen72hQHYkBaAAG1SI0jnk1Ftgefg
RvrX5KUeYKdhsbw8A1aGLIoSOLvPIHdoydmdq0YYZWXCH6fHcYExACiZQFPHU5AV
QjAVXpnXV90Osx05fW5hVnpF3NcTUtC4UeBFFOw2hRStLxFnCbMMNZWnsJyZGr/8
Wi9kLN+nDnkgwVtaLeM2e3uR8iUik02AiJ03pAGZgTnxgKkjBiSfX9j2JePgygd5
9tUxpfczTiGu8H5xlNINZLGjOOI0s/ko2J+b45k1bOgFnEFn2iweiFuNAP7nKdaR
jE2Nb0RxJpS9WLmlVuR2YLNdFUvywZXMYipXvNsMVC7vR7NNnusxWas/POFifOex
aw4qtpvbJVCLgHR2qlK+g9VqbLc4OAQWO93vQhRnlGLtkFQqWmIRoSkvT2+y1E/z
wUXqYXK4JqC8UTWRsj82yfzSchUPQrUDtorfaINOStBvdIiEf7zhB/2rAC7sZNU9
5+UOdJWyhpmXLwVsvltC7aAH4sOdhoWCexvGEppVs8pvFe4GKvjH+GZgmYBmnsXx
UC9SzAGSkjzqdJZoDTZ4hAiEyiCcmbNspy3UgnHdhY54NbZN0TEqijJmbRxg75wd
q9MtW8u+70JGSLuPPRBGF4XpGFQxCUehkl0bCgc25otGUXg+Rwg2SULN5J3pxqZF
VPKy//pNpXF3f3bpBQgCAxA1Iz9w2rrYVDhI4Zx3wCxL/QM1hjIbLagdd3qu9kdA
FnSRCPlmEwuRQlfnA1MAgPt4kFjnffeo5QyLw2uL2Nm7mfUdhDjOE+XAe3FSz9u7
49Xw+IEThg4+58+iSplZKX1QJDxaCw6+f8bUutOYpuVo8FL+/pVCdxO7mpA/yKpc
8LqI1vN+5yaU//kZF8fqysH2a4twCsIJo5Q2qSWCKYaExzcw7NY4yW508GD/vQJU
k6ybMdzZ7sudRyTMrHNPBrkpNNXlLECH3GjwMnN+34VVSeURrMyE3bMIvnUTTXtG
f9E4EJkTxN6SpjNcidJ3FeEBlFZgUSv2z2bvkETgaASiaFwuXAqiRcgGvW0yojzA
qYLk5y+2EPz6jq/ifL4/p0L40DP7/p3dkTi6ufZYlbgyvx51gti/MsSQChCK7QE1
Msk/HzGkf5uT6WRwu1pGllfoEYqvRv57rjRb7S3eZYzEx+nEEbhC/LA6OlvCmbw6
14fW7TUHT8lk8AKJbR7HGfs1/mauhZXn0pUJg4Q3kEbn9zr6C85wKrDzs6zuyRi7
4yVI7xR9Fi/tCBKedlhbcsTdQ8LFlZwHENwJm8wwdHd/f953EHWcq47Q9L+qft9b
p9hA0lnPA5UP54udxVXTc1ukb0efW3nWC29URMfy1JooR9bou8hYoSiBo1I2vGUX
Xgq497856+e/NVnQCKpcCX2IMFQf1ei7Qp0NdohRZu/vbBvoiB4IF+T1hR9szNHU
xriCBx2sG+QxxiGtV9SqUCdw0TdedH7FEriAY/UHRH0ANTslDAnAkvJwW5BaJq5w
x6KOFCjEMO2mtEnzCXnIw4iDk9eVmACvVJ6Y0gpz52tMgXnWd2GfIeh9LsQyqjgc
XbKSntKDLge5T1HZBbQdJ5sOiAwHDb8J+lCsLBnU66ljqZ5WFY6853kCz2q9sjty
exSgEEWUVLyPZGmjKtNoTMLUxq6BQXR7D9VDPNaVnU3ZLmTRFKs/ZNe6aqylfvxe
2NoANJvSvR4YGz03viqnGhir/4zgILWo/KbQOqGz0lijA+EHD6PPg7cI9PiFRDQh
sEb2WC3uCI9m+KwqND36bsIoWE9NwSH+68X95sAr/nteB+au4iZIIPmzbcBey/AO
+eIQqzmiyFmCjWcjwPjauLm/hVV7E/Bak8Ow4A4xAJIbVpdeOWwnrn4/Jy+8nAC5
giJvHedx4ciNley/tJGcO9nxhOzStjgsvrjtSzZKYKegwC7l963DYQF5LvMjJ3oK
4divX0A2DHGjOw8ObxCUhkM7N8t22wjxBwlIYfFitYiqS/3PfCTKxi+9v9X5yz+2
17DdclP8bH2+sjEGjkATMD2se2jWgJ7q83DPtDQbn3WyjAFftZ7k/wxdKoPZkOaB
Z/Cx2AD8JRti23xRqs4pNsKhEpK1Ti4+xkcPsn9y5h4tsRohJix0tUpzWNUc4uL9
sPWDEYckEZUzc075Osb08kVfcZs1M4eRafwKfCdnh/Uj7hEZamVnsJBiJah+nnfE
XAD1/xQjqiFwD7gi0K93i62LqiO69Zd+R/6dEgphY0CIH90L8OewKQKzvA1qQ4sf
feHAFDeAuZrfQS5D/0zrkN4hujeeCv8hgAPnS+KNnfKTRiRemtJuswaOkgo5ebmg
2X6pUA7keF0NnbUPaDqDC7aRAhmcIyNVvbOhiLfeC6Iaf/q/jHQ/j7/X+JX+NLCf
1Fy5kxeqx2aPrI7jGSKWL5/vXf9ZXkbeiQ76V6ppgKJrzyH7oAOvhV43Uttoqqks
gUm32PMHTS0QW8LnpymtyvKlhs+qd+mWvO8yQVHn8+RhCIPgCnZSxQozlE+vzFYx
mQHBja+PMrNsHKMaxpGukJIK2f059/3c0o/52MXpECp1DYssB/IixFDVaPmWO2d/
AfZ+Xk8/lKAjuEhf1zMadsRZ0lwL5l9mzjHWhG2qdfFE5HSWyLsXx0cDum7nZZZx
FC9XtJZ9u2MpLawii7sCVSHv/hfSTMXkT+stJoaCxoGg8HygIZvsSf58nECmBMlr
/mMe8IwOUP+waZ2aZ4lSHUddPvvZIgxC7AUT97bWTL1H04MONKo5v6Pxyj5xLd0W
H9g1L7YcklZmWJlGTDbRkwDQ3YQ2IQqZg7AuwEPkLlkxVqc1hoMKik/gqSPQ3HkL
ux6abYks6RacGj7JfGGjY+kSTnORYRZwgu0f45O178bmKTAP7BBAcSSuwoSUBvPy
pzd3f9pYIV1wKK2FwQFfzxjZJgUP1zW6v9G8CpmnQ8OctXaFFU1hsQcaVPbK9bjD
2XBLmgAxRhg0NR2YyIkdphgWykQ1dSd24ZJLN1eZ640KoLZWt/RjpH+/nNyN5yAN
Apa3TvikNaEaMIOsVxubqI0PsU+Uu3BvztgKXcRMfsIfMg/ae4s3mEBnmDZnnUl3
L3EA3GDtzv/ap8vyIvIJt+yiU+icd9gFJy5a8eYIsCkQy3iaZZqUiFlRGDDpAP63
VrH2MGs0emogPHENJk69hHx2jtDH0mbhG27KzQGhv+bgOy2428rgwVwVA32FKDjU
D5LzFGlI69RdAkqvatDbYTRZGHBJt17AyeWs1RJKwd+v3cn20Zj+FFYRTovZl51I
3rUUweJTPccSNm9IAGcON6Af8/tQtYFNGMjXeYFDAF0kS5iLumzMRIShr7XYwqsq
7EcGl9U6nbyl9mvjWLvgMq74x5LF7AWsb7rdK7fskWK2QzghkrXa8bghRC21oYKX
eZFiaG6w8stE4/Fx/jERTs9m/cdDB5vfXzOEUr4zsMMgTKGFPxvy4ZrrOGSJD+HL
innBrJxR9ahio/63QB+dKLPCfInNboY2DGoGPx6EjDguUj8p2aWahrhfRsxgNzly
5/yVp5XJ2yIWn/BGft2T92OD2kBHXw/ETHVqVIWWk6uFyMlu1ySMsJ2r8s6XKSe2
Y5pFXkIijM1LcZyZ1fWCzYyJG82ZRZ5UpyO0EdTJBhGuEMOoKXKvdlNl51DqCyRp
1fk65QGkt/4o0nCElx84UdAIJwZbl9FsX3wFzdtVrNnXUXuBR/EvdOOv0ItufpUG
ZwqiW4ZnWRWynvAD5ixIYkzWxCGQ9wWesfcQHpiBxSh3I0w+bnivqB6WCwO+Zkc5
pLq4N7jiDPAVZzxejrkbv0p+Zuy1ZSuXA9X6InUWHcp/5w4QPDqCCDM3fF0K14iL
iFEqtSGAkW5H+Abi5wE9rt4k0WJc0PDntSjg4GuXl7+R2nTyyh0h2wj3etpc4Cl4
BM5U83eC3ufI5piXYcV0cAp7PgQjJLn9iACGgT+RrCfweJ5BsDQhp4YiLylWTFKm
sJIsPL/E+P5A+KhppmFzmKVgoikb6ZYP3G6DUS46m+xeXAyHAM398m8RzD72/k2s
r9vLMeyctZD2lQnfs1LYxllgseTOC9lTbJ0nbtgQgzeCb5pSvBcahLri7zcEnYnx
UkyrUV5rRqHlhYz/PjV9YI//L5p5vcYhGJvAnql+vaGVVJ/up8UszrRzllUbwO6i
5T0hN/hQ27r09GJ//zTO0K6Xp5LWpVZGzv+NDG/VuOEG3KN5BnJSrHKsr8st+vO5
OeaJNK9IcA0owuRHii107d7laRKo4y4JAtUNyX1isfWEWKL0XzztniZjS/070A/T
k0E+ODwGgVopuGThY/XkfGvILo5wbJ5tdrEmbTdPBN/roVF5q7s9frbW+lACXs/N
+Q4slaOcNOIEFgaU0BDTrqU1BSYo1pUrGx+vIkJz3rnEIBRj/oSD/YUwOUVltipu
q5K+mlcJNIgLHU27P9G4gl9DGTqEJvd79dwj/2hwhjksuQXrDI+PZbPTjZS2n8j1
yS+MWymFLGpA+/NFlhRhByyEONP2Jo+CumlOoTFw1WenN1Bs1ZUWvUKSBp19tIJr
ctAUXj7hcP88H893g7RP0+jx4qmuwbu40OQk90RPyV6r1Yul+tzA3fH7G6pQzVUB
Kxr2SW5rdwZFJEn+AHcCjZtwxKbBMNdUYXmxqGvgm3WKOe/R/GA5K7TUkvtNZpoY
JJ8KGxA+KE82AcjuCBdri6ovWHBhi7UUQ7LI5DePkIZ1UsshSuv0iObDoCKLRc0W
X2ncbtCHVJw6CbhhlRRNUWs8uBRcIi17pLP3N3PmGs9Pb9QfdmpZHt1nHeAtM0s5
slrNxnGnfeKEcJnZoSfsb5BHYcaEKEHYRJ9iGtcCrrMI83ilXrdUBVurYqDU/pUz
5sRDdFeVOEEZlw2SfWJ9RCZq9AWqKpFJBzQMjUaqkmnAnppSAPWYyFLaEByUBFPW
UbkahcfWM06AJv++Ew8YaprQ5l7iXFrngzNXBnNVFzY3u5tes+GsWNajKoiQaPMt
FsP/Tks7hJFC/3u2GwGkt5nFyrA+j9/hfsSSyfCi27p4aAPi/66ktc189QgDwwZ9
P/oCtVDcq6UNvo8/OOW2fIfjS82COC2ipf1t4/jGuLhy/zLkh7YzbIHoFiqNsZMX
TWtTCSTi0g7S2rUrz0GPTgqkMg+5LMnzktB41zZmluuQ4qQYF95bmzeYk8OePV6y
sHbXtgkPw85eRwtomO6ybtv2mDcaIRikf0kl/UsAMmiBk7IbGqXpFBm5bfPnMBCn
UL125YSkfnvgl3Zjt90dmMrHWhByFFNSXvH7mPTxHWObmye9kkcrVVl/IEKLWGSk
XeNhfce3wz1adilBhI2y5z9gW5MD3aKLGasBS8lQcZFxfJppOjonopMG5lwT1E9E
7E+ld4t2/YX3urFr1w0NsVfI2ovHTZF/t3BTcOtprLYnUq8EZqccGvxJ26h3fOzM
mU3scFmsVWsCQSLuTUzIXb9SuBNrB2BFhjtl/8SkZEWquH9JAvX4Oms9bc8Xnuqr
ONSe/dkcZ+v2xw4peSPSQFX33D0UNYPIFdSO8Knu8s3P0cdllYrRzuPPiZwjwz7u
MxQ6S+/MeZk6Ac+zDg4lu9Y1XipIDxt22Ih/dj/f9UqU7HF1c7O2Uy1HQFx6mRLb
kG4hMyEmjPpt/R0lFq0s0PdnRreiyTgfT294J78QpqZjzoREv0ZyPOfhVG40EVrz
TNPurJSl0N4wigvfBGNTfdsOcxGiRcyRhH4cUf2cqZ23lzCDLiQJsoU3puwvRnpD
9YrQVAtRtYK8Uxgjmma3gKG68wKF4c9MQZopZrp6IE39R+8XZVHNwVetmJQqKSzU
LI+5FUWsVg0W5FHPqZyBs19oiKPpa9Hxj9RhduTszdZ0HEy7dcMgjlz2Wq0KWnFv
N+gA/Pm8kXTru97f7po4poWg31rz2mca0dXqda7QT2JOB9w5mPozlhkErCDG+2LN
Op99rMsfnXISnKcgGYdsfzQDGBg/7UsTDDpg/YIO/rLcn/RB6YO+Kx8hhEVNeH42
wvPuyroF4nt8cjm0Pd8hxdfGlCMzzFyKaSFvwRb/z25+sHBmQlzfT/Hgbe02vo+V
7Mak40/ql+CWIuiESzuFw3P31+tfTIuocIMOi7f5Tdp46oHwOoJ0NdhWmBfsdqEJ
ny3TZpkyWpVWEsWMU4YEG3PNnxgSMZqZdHlOp6pGO4s1a0xN8+9T2rkLp9zTt65b
hPa/HO4REGKAXR4drhF4LSeVfEQBCX2gIBE+2EfNTuu6uizGAdDoFc7E+c48lr3Q
hQFR9sVs1XrstjKUPfmqUfm7X9ObD6z1KaoMGHKPc+uv/4RBhzeWQKdoniQvb2Bz
6GzLC8vIrr8xLZRpAezT3xmYhYuvBTPg29Qbmy2QkOuL0hPaMkx5FX+sVTkYCxg/
5NvMN5fdDsUmv+VujpZ+O+sdOasj8Q0wnBF0vVEndgzk4oVoAicxDqO2FZkz9stD
J6vyhZvujYdYhch/G2OZwESKrVcIAvpnBopIw/5hZKure6Pg0d+jDSoiALHTwkjS
MjZjnkyk9QGMyBKfGxtMF2SHlyUBkYDutfDH0qHMaJXFONuVXc+/9/Imre7RUXGk
hRGviyQertZ1sFpmxMP+rb/s0o9FNCYAREE566yBijIULcT0T3nRNQn8hva07rtW
Ws/7P2Zv3iFMUYOftRBtPz6xDdYndNH7qxp0zK4mcU8Rqi9i1cEdT7H2ZlrkXo1T
WhwoX6j5XxCCTic/Z2jSyioVQPfZ1cANXwtdkLo5W9VN1HKa14Tbzxsxq3t1QYZy
yB5sySd51UPI0xM5e5dD/mQXaMw5rj1nvq6D3lC9O4awEkXn7PBY2LPOkNvtgAzP
WYrbdIRxEFVISfeeLRhtzcJUqez2vXGWHydUMaT16FdxJ6gyx5K1OfPynO5N2Irz
WHrRpMbeTNzCcrucfs0BBsT9QzbO3kSou/4RS49poUNiFyQnGCq3ue2r9T+RsRzt
o3/NTqcy7kh3JaAQY96RxuXa+IUJljGxMoK3a+P1w2s+dMiMDOxD30Yynf837RMy
RDbkuT503TkOvd1ck9fgFBcn0dnZOAC9tDOuLfoWTzkKQR/GhxG9MeR7AiLjY9EX
++pIqoh/g1eBn0HfpXhh3i5TdQbKLnf/OPstOfadyOasCP2bz15F0oqQRFNbxp8d
Kv3yFgmH1SOQyIWwTdnESBK2WJw1GNLfD5tWliTmMo2fVwDBGBhp7Zn6k5uvUk/C
XN8HlyUGK0fe8/DlAfKwzxJhtDoTsu50ryRq48KZ5Z0hvhdA7b/UimXhBu83tUfi
1oZx4ZtfVHivZHEdD3aSSx9mnoZlCGYON+VbT2OBGMF6f3bZ2a8is8injYhdP5YO
gJO+8ZcIM4NKS83D5UMJIZ+bGauFWcMixOsmOLRIBhCsxq9BVutkWFKpFmMMSsoD
1+ycG8/qV8HT1lgZ8gkvIoexghBoQ9DiBOToJdRdX6kz3C5CBRn3QT+dopGI5jTi
hULJFWGn178Cdf0ISUEzCKNxjZ0wt111zFdPRGdIyqik+n/GJGMuHyzALEtxnj+9
5F7binuMJVWyZ+9s97SZH8qN+hHX1C5YmKo7nMEHbPBu2TQqfU7FP6acO0qdxR3M
E+zv0DU8sUzlv3TLJd1tiU9NjP/oBBIAQw0Q9QujoN5WcebMqItUaTY7GNmRLn0M
0EmvG5V9GXxcRgfkMtAw5lR4Eo7SnOsZGc4Icu04cYOWgmYfm08tytDxUuJzblAq
Mh63UwaekZK4Ofc5ary7JE+0FK1vfd5dnWsmidAEke4Ja3ukK9R0rC9fqs9BbmTW
t16T86X38/it2ybOkMMY/Uipgiev3TfVIm+ZxTMtN33Ds4cvbFs4QbuK25IcRm3Y
BGyEe5uAvnB2bDs35Mo5UJylPFL/yNenXs59gBcDglnL5+tdKlkx81X7osoIqvS+
Z4wtRCLQ/fokzAb+p32e8jTXpQ462hOCng+5UQ1IHkgHyvXzFDcl5OtsBwjf2agn
Msev/eHnSGlDf2++OsrO7/GNP3QlXwY9yJr3bprkJKxyuSm4FgfmRloGT9Ou4CFO
yINmmINRLSighhsnMeoeyVqmkzdGllt3HHesdQ1fpZLBIlcAQIWPeYW1MBXePZ7y
lvOH1fq3Uqd/HLPyHV1JEsJD6xGFYpZxsYbEXKIPMOzheQlCOKhvTiTHDYjY/qH2
vokTydXDaA4CBK3eTLoATMRBEqG4k0x3zonWwEuseRy135vzKOGBPRZwQfDdAzzo
YRIWjQ962pkvNxlcQd0m4vVACbeyfaapZcTZeVquzmiOWpslMbu47eky3l0m2nMt
5gVAu3xkURSjFGkH0SEPIi+Z6uy8xLQ9R0+ahRy1zMJFU6emW4vs96HMGfxHV3AT
v3UDD5bjK50BKJNx9LxO8pz+HMEXjDID+Lc+6SdmzJZg2QqJpyNmRWPGNz9u5Yy+
5L7FH3SLHf/ds3h7kofvq/b2PBfDRqy77TOITwo8+48F/QFX3pyGGMPW2VhWBrYS
Ix2Y011x+JpbeSnFGhdQWFUR8gUzEcFBc6LFACYbKnDRYsE+zQbw35aCWTON18di
GDVe8N5qIp3G9P0SYD/Wm4j4mSwcT2SyUajbUtNlzXC72k+hFfGU7ZWRdqoO5R2I
J5qNnMdJr3/fmvLCUUMKKsnWS8hfo/NYA0nqkYymppbsboPQ+AG6oVagH6GY4goA
3/hmhSNljzIl0FwmnO88fNHPZyikiAbcYxE5XOhI+HdEWG8WKf1pk5soWIG7GYwF
YwkhY4vH1GnZQGffegc+AjBvR5mkSFoK5uRhUvT7N7fGQ1i4Z7X4Ns3IbHxvDjSI
YlNev4EP9852HzexeGuhEFvBCf/nNqEyKHiYJEF3TZoVPxTFyD0ad72Mil1RSqzY
bMAcOV7j91QcaSZ3fpTgeHsFlYfRmV9AYv3floOHfQI+N1o44nkJQu7VaaOX1vJP
RTLn9C3hSpZKZEKqMTQvysavfRp1MRrUayubEeTVFjmjKgs2ukBEBktZZsI8Otzg
Kv0nFrSGm+WxlXSzKQHmWHZdOGEyW7vDv2ehgMjBOu8+WpeDBrZj+0Iv8xGXqu5s
DcT6QW2CignXO6W7rJHpMRMihGwPOJYjzO5TaNJI09n+GVxvOB4850OKxtqy+Kwz
ka/7AkknNnc0duDTwERVvRwbZ9DhtbKcI7sW5oSFRqNHJD+xWyzhd/yZIiVWtkI0
5HLJTgv7NjAhyIFSPEe2hYkSFXrWpDXbbXtmn6M8+aVSsZXedrhDnDfTp/ETls5d
UaYpOtMzDjkqQ9hieKwbenO1WsM9B6SLOJMHvnKFz2zF5ATR0eW4pe4ODSFo+S98
fonusKedXzvXsUm0s57yzNiolUwu0aWu9QlGA/TRRYkHy3OAvAV7jk62ElBAl0eH
H+SFckcC0iTxSlBuMupmPmeILyaSm3YeM6GYJPF7/snVoxJylcoIngXaU1g3L3B8
xn63BdcKW/RBH0jUbXFhj4shDu1EGpQ5hEvEhrl6RpxCFmp482dxm6fECxdV24va
ua5nw+UmvDALXi8tq5cl8+E/lx3CY0NFAWeQ0Y9gS3kTD70pTN0KT0fnViw8Ctn5
9Wu7/FUdplJMLNGVcPuhSOIYrzoAVAXBu+bTcX+RhC8uqOr42Uu5N/Xkr+lmXRBh
fFO5VTuNFzEwHuzdP3dUnUPPPuoCsiEyXJnS/eBwBsWelTNURI1l9k3ZZYJZQfrt
/Nzjx28vDcX6n+uk1iazmVxFLcx5PFZbJtFCh02XQar/U3D/4/Akh3hHy0ZbOCTF
J4hX22O41MPw5nXzzDdNe0dfpsm0OH16Qb0V/m7/ZOajMkkd3GEWHUBLnUIkA1dy
YYkaVQn4dsHxZ4aDsdNTngX2bXtFVNWsWdttjUvSECnT2TgugaxVjCWTa8onZmQf
oD6K9PkCOt6FbldQ6MlUlQYB3xv6W6lEtS+ysNIZ+wsk4d82VnrBMRtJZTVxpjLj
DzG3A9rz5u6VcigC2kNEFRQ0A/7gsIf5Z+OivtUnVZxpTK5AvRCG+uovRQ2Ecx7i
7LbE4vP8k0/NPQKKfUTYAWUC5ZfG8JXVDNpMRkz0jyaggquL9mX+iHtQ7CyPbQ+f
37ce8a84OUV+Yh1FcnjvJFpyzCYei578aHUfNnqZXB/S2vzXEIjs37iTZ91rcsDb
vxuUh+MgGInyBK6js6O5gYGMXjSF1YmkvlLq/fhGgJqmic8mB6DcilqlgpnHA9py
8s6um1GFA50ybvUDizbEN38s+pPokv0/HsxZq2Yf5+1IEiRGTyK5MzPklzCYwUr4
McsIxfJZFYB6Mk/IFF0nkj+ue4ISr6psG0IwcQ28L61iJsE/zrgiuwGvhuk8HmV2
wM16OiElP0i4Ny2QT17adfK7CmaEOuDVprL80T/rumna5fj7xxpQ9rMaoQSAAqfX
eqIVuj15lYIeTrpmOaQrtvTWjxnbtUNSei7cxu3naVjRfcWMvudgPrSKvlXviv7f
7A2hDwfrep9/U89vNueeLkBZtLYcnmULJmcfql9hatink4vufAnrDzT+VoEB0HAr
LgXVxnWy7UMtzbgnrZB2q44qHdnMsNmK2wBluk033WYw/iGbNAr+wTrQ0FFxdy5G
WuFgEvmdiCFH8PsUaK1IZOtYFz8+jynjQC3shUZq0YqjMMxbYmZyeB0ckF7zP1eS
ENgOgyj6EPPvEUDCSVmOoenYJ8v2H+3cyy4gQOK4AvI1N0rk03cREb8LNivanFEU
Pxkbv/bwQNgPuoIZm882dGFOZ8tjG4oWj93wrPRhc+prFdZQ44mGmhZ5ry5GlHz2
BixkG5JXtRmaUU6Hcp87ozXQ5tqAmUsk1gGQVdLazYDwGwU589sUqgnEBbg4ATFA
IKFVU4SlB16p9S8cOPG41tqNYeewz2DCYfE0WpvRdkL4LS5uIuqWmfYlGhgZLHBH
GT6QbUXQdAPU3wghk+KY/dWh39N/jSbaH9QtQPhgcmXtLlh2HCNbMIF58zNZ+1PC
j4AFy2a2H/j1wPauT4e+46fGlQc0n6K3PGZduyFTf/0l4Xn9RjIL1AsGdgouzApj
RY/erFv233yOLxHorCRat3dbUl94XtS2Jk9ukQKZOpHJCvJFgboXMlMDkyzeDn1l
uTY2cPAVUNzSTT9PXkwR88jMh6YW1504yuGGy7lECaxksbqX6L7CZmo0njYvbHFa
De1/FSMrC/weD9QHC50F1gckbJbd3DD6ZBlZ0GB2RiauKUU51w/epmuwb6wJrR1q
Cms98wfXZ42lf3Z4SpkX461frHGk0Tyxoz6uchwJ1lMnH0/C/dxi8Hq2q8UjaXvp
vwAM+Q66eedLh9440TpElGq5Z9zbGVtB7Gmze6QLXQhBThZ6ZHUleXq9wkzPop01
bJf9D08zZBp9CqK6YY+7JvT+Ahp1S/6wxqY7nAteq+QOlzyywE9jocTXwAIaPkxR
0TCMM5OSLd6okj/t5rkHV/6goywjokjIKVtHsK/fdEVVEihdCIf1RxL968k81IoY
FidREIqD34eVjqJck7Y+S6+GCFps9EOTCz5rTX7AelgU29JbKAqxbKshDkVdcgAg
sNLv/rMODaIe7wL8YyHcUZOsKpxHoZbovvIfdnFtImsqB9KnaJXP85hHpNTQNi5V
AP/s03ObYzZb/OfXdto2/qNP54GXuc5/tc9Nh5s6Dqk/N4svVQ/ImfwH5aH6fiJO
jnz9DI0JvmxNexNkfwrNkvY9GR8wCOgPE4ILzXnJ1iCYYsdBsu8z6Jq7du+avsi5
us54rvJOY24Pc3gwC83TXsQo2WhOCE15TRFM0KE59yV1fxrguvJnoPDj4OXUpNmL
Hm5wqpVUYu7KhqKgVacpLXOkEcAIUP/MPDlLtjJL7qvLkxMBswMqKhcqJaWJQ2qR
h3lF8W8tjY7ohxxOD1pInxJRhUgBakUSFFFg4+Dy2xNacU/9zERlv9XDq0+t6+TV
ezM2JxqqjbnGIDlDwtyt3nn/KWXmBf70uwVg+7q7Qr+2gaJEgVNqXgHM0DnF6AR4
YqbNJ/v/EivAdx+tyN0dzddV4HriUdFnZU2CDge0Lg9eZEY9mS57N6im6yueu65F
Hf4tMsW6URa1/EkIwtpBerOc2qBFeF7R4chLYOmCVsv87aFHm4wfReYWpZwBIpfD
C7fWJTrFSnDgk0pE3HyULpBU7cyak0UO7r2wparyoU/NJH1Bho0JC1B91Daj3x/o
vd+X0lDINbeXkrgyfmmqCQC3BBGTGKVcuE0MAEK+uMNmzsGlUfLcou8RGxfid5iQ
Ync9Bt5Oo3dmXtWo48qV854uiyDBhXVlhKEKovyT8P66yLrk3tAGhfyvLj8/y2YH
x5g1nxfRjeruibM0y7oPuypj9KE0RJIwZzDe/KWl+k5VuDJAYyMdFL6yc2vSZdF/
5if1nc+QXjN3uvTJB8Wqan0trxufYG1awvW8I8quw9HXZLA+QF9E39iOlbTBRE93
q7KrTn4MaS8GnqUGierieBuVbptBVgae6fJ8Se4zDGg6/tUNtLVguWZPOoXVtwoe
VFZQ6PqHpbbH7iJUKRuM6/zo2x4lNds6+QnQtACaWqF6wr37C0R7Vrc419iRSvzu
1WlfhLcDemRxFfK3PYTaihlJ2ryxh/hm/8vzXLlmStfCbSpPCPGfqBvE7AIJB6Mw
h2b1ya8pYOio5FcFmKmgnnXC0SEuu8inpXLKKLu+m3Epdh/zUAKIGnTZgliOp04k
Vxd9hb5lVXcqedKEZnp+d4j5QTFOaawBAvDbNjmmdI109tY0JXhXB1ZkGgg9KJOe
lykfpvbsB/CI7oK1qPVND/LXREe5ZBrb8uZqhKeDGkRjr9ojRJDqkbRXp4LYsPJG
d/tVLuqB/2saZpft6KLhAAlRqvZN5IxNcbPJjM7ekt9FlaHAIYddX+aaO47AHAoG
gQhdJoE1lKidaJgfpXmlVn8dYzLSiZIvF+KXggmj7mB1FYNj76FwW8KLxQZtu/D4
D2tbRLG7q7EwwMKKDZiTgkn64gDr961aD5E8k/hjDVDYyt+FBGbQzprNfqdejL+5
bjQxhmXETiM2vLtcnn2TfKD3joFD2Hwq8tU2W4seChM0ZayJU5/URHM+eVzMb8oJ
khByydSCQTosBowOoTDJ2esNQMpEPR65NGTTm9UnKyNqUuItOA9kbTg1Rzk7t3Ep
wdwxM9fXcR+6U7xK4XOCSYs6kh3/iXbiFr3DA1y8CW/5LxllqpdoxITTt8+Fd18S
FsQvVAg1puUak0ZIWGtu3mJRPH6BhI1ZJGO2qB4htA7PbHZvDPLZFaJAXU6dxPGF
tESjoqBvmQJ6v8Ac6+WKIR2HbT0cwLhJwJOfSPUkfakUhB5lekHZMXd+ETB+APN1
1MECL0ubazio7iQauaCoZ2GvMpqwJSSyq48q3U0kHN0EnAcPtAkU5qZ31TR5F/0c
aucxvB8vYo162ngNQECd+2Wp+7paYBhUWiLGvALfx6bdlhfzyq9b2Wm8C7IdBnSz
SW8fScSbzPPxPXA+23JycqgpwbCPdsGkb7hrwy0nL0R3dgKKnbEw2S7m9ieS8b6V
HY85p4Y4SLjOlAFNHMYTI96aLNcVjBc9DOFw0toAObBxvXeAzJOjmqYIpXgQIo8g
/Mm8KCHHUv8ceARJ2gkn1/l/XGijK97lIpLa7BLwvbi2hr3qaATMdQrPr12FDtqc
jPIcT5d/w1t2hu5cb9vt4km2oLaPhun6RhWr8HhRp/TBPs3dtiv8C8PujgbiZgiB
0/sK4s0W/8oD30+mXnbDudnWeFEbIpAYywuMUFdphwFkoPl6yS1GjEI4p2fsMX9M
vuw+FaGY6AKFaMwlHSKHfGmnlgKobgVgul0nxoHpVIul4GSTsUVCC4njolZii2rE
p4rgjYZVRQeZ4rBqXf6f85g4rtqbuPPxT4HIfKp1Ay4z78i+XUtWloAFqRkahigU
uwD1uN7LXIDiv5YtcblvO4G81L13bL7uYWMc7qTeBxBufvbYjMrZ0oiPaUy5cphk
T1psTocGKA8nQRKmivtUgJG2Nlb+2lt7lvnILKC2kimI/BvszQw0tEPzzpgyqFeG
DffesyUNWsLOlTXuPPHzLeKILughPeAA0JDwk/W5f6ezcUROPB9CWyfncr+em0Du
0DYhfthcHe7OwQPL7M/TtHAsEuFtLLYu6G5AXYxMTxqhB+NG+RL2sZmwEFImVlrA
BSDHvo1bm2XlC79JxW2XVg12qJGZBqphqnYNIb583RXFYGTvdta7hpKDgWBSgLCC
LNU3lzdPJ5biDP78rmLU2/DeM/Ig7NvAMSwqq+QTGSQ/Me3xrl9SIuFM72wSan43
1dCmnOY7irlunUs1oapHAbNiSLh3FUpJ611tgchLkQuoMNwQ/2d/iEGorZgIpKcz
VHL1jZO4RzY3nxFmS38Qf5LPGzijpbml3KXQnBwwK5ZN9YV7EZtUdLxCwBGCh5SQ
cGnoQ/rMCLdPC3o24/2HB/lQ2a4dsnjtNIhu30DTttnvAfSGl3mDjkSKcBSys7+Z
5V6wNfUK1TSD3u+beqiCkI5TtHUUNhEuAzU3MIc8Vy4cPU3w8tmmQNHxQYqmta4M
K73/pnY9F3R07AT1uXf2YAgZXWF48ts5Oa6XgMrlMR/6Uq2Tvwn1W0VpTBEPOLHs
mqulj/xQBAcrnBn2eQPT+B1VCdr3KIxHQ0HHj0dVGzNreINYpQCHq22SwanDdYLb
O4RcHIqYdpJ0g22vjxSmxl9jfqyOn5vwaNVav8aPKTMGUeXvUbQmueST4OMf7+Aj
UiOc9phcykcBoGD9923ahENME9mLgmJp4aPDAk121TkfZq+TuK67J6IoxrjeEKiG
6PEAkG4lPrr/3Uoeu0Q5q1KTpKNzLnpJoU8OpuIUpnD8YqJbdLbeWjtKFfF/MRRt
Rt8aBrSy2pch2U2X8JB5ktZ62E1eN8vvGQW845xlP1uItEjsv/7X93mC7JYTmhXb
ZHZKweBSsdWFwM6SfQDUrGv/GDWQrn1yJ5j9qUQ0Avor56rruV2N3XL+EuBmFkAr
RRBIhcrKPP5lq0V1d/Q4pIqCl8TrI6tLwGCaXECRcs0+hA9+tZmQz6YsLSb6sEfp
uMA2tZuEPinbUJtV2gXASlkiKwxdXw8zIhe4PUUI4UwuUy3NqImWp4wc2JI2Vsql
yL6mVTY12ubFKw4rKSn6geT/PgbztPG6KwhINCdTIFNEFis7koXY32Z4/6/UjDyX
1xMbVC91smrVSxtwZsrbYDIgqZErjmsBFQoNHaUVYq79JVz6qbvcaTGlSYzWv6fS
GU8pA5g0Q+FuVRQFbXsd24Q7fPs+xo+NU6reKv9aKcB5XczS4zkciEedJMQwv25J
UdQobsmBE9EaahMOyTuNmA01kjAeQzzuQINzd+o8co8/vTaHfrE6B0jMfKKxZhvM
EXSByTkIgesUslohgUYD7UjHdfvxQzmaXrBJjSfZ3qijvK0VpGJDxM+MwX/6zGx5
/YEe0NcXZbkGq0VLwGAQDRp+UZoKZ+B3HPdfDNJ5BVMqx2UE7Ckixw5NqwmBUQiG
wgBSd+79MOu4SsQ3ODHwQ/9pcMQHJPEIPZQpmJxV2fmhl8IRr9AqFDX4HfH3jzFY
n46dSzUbgrYCmqAcaUH2+lLet1AeHqR7/EVaQJwKsp8YU78ob/IF+DPdWepWllq+
qg+C8kspv8ArU3zyNxCW9B9uHHJeE0ILasjfrDdcHveRXnKJJaeYJCaIbwqiF++6
jK3Q7ran72aMwG0tOfy/QpcrELyIu2prdi+w69MwjWtxV1cO7LBCUN1Vg2s9IL3k
FXtRmEIe56GEL288UFMW2PkgnsgH/aNGdrFHaDARP4eHgQjBi9PN6bFvFxoKMH3D
DAv49irzv8ujpQNUeA0a88TQ9mOswvrQvcciWfS0/odusrvBts57sQuX6J9u6iwV
rQObVCI3L1d9SwSobzibYJA0TasPyjrZRDN77LuS4sWkYhngj+6TRq8xqRduOIg4
RkvePcY2Tr+utlZXE7lwvEXAsKmdO8bSMu0g9O3/omBOHjJyUi0H98tQIScktDa0
+xku/cKF7v+rVhwimg78k9MY+1jO48Y5W0Zn8d/75FLepKVNd0AdOA/FqtfnsPk2
2MxbICwmhbYNl1EAIeqHz3Q6hYmGOdV7LLyuMgtME6oP7DsVwHJ22c6pbOMwr9hD
myJEo27l96hGQCquFqB909gV3u07cM3nRdht3LIjy6HgtNQjIJmJ/bt6giAX9U5l
zWloAJunZo2BqZqV+CUhQE+Z6+Xa44zteqOdv3/XpDRgVAiyj6B/YcStI/6p/2sp
r+CTa1iFY3Ko83Bb0aZUfIWLRc3FKUFyzjihpQarCG+U8mHvAe3c0C0c9Ed1j+c/
BY055u39QD7Og4N+YGN0vMMp6Yehk8iuaJbWmSPuPZMgxEGTXSqnM+sdP/uPSw5r
caonCQIyHfGkCMTm+KqWSCpQymGJXeqeMGPN6NH/sK3OrCkqshUtf70YkZiJWAhP
4xC4lV18LOyZpqdFwKnbuTD9XZx7ana+GD/25w4RCNyH/LyEsjPrtN0sxeGEhAGx
cRnpewSaFF4r7VMZojK3FGB1unSuhf///Sqdr06A8i9o5KE8KfbdfCUspEVSz512
1eHgrKVlI4BtuAAPE+OgF3SaJRLw/KMOlZY0cFLa1OJcvlqK7ZguYwb8wM8JkOKS
61sxkdt4N17/yuU96dQ4U/J+1jtqCZNC1ef+ykEsigWf7vaer3wecSDPHkCljkFl
5CnT17SUtBHJaw9oi9Lem3ul6mNuf/rXNNqE4bgWyrH+NMaQn91nM0ypzih2a7U0
bxGUPZBq8Lt1ARfBQn673jC90ggpD81X2Q9Qt5CopkgUsF9Q+vjro29d0/2PcSJS
F6XVFSZaLhLODwrRCMPSg9facDRa5oO84GWzGC+v/rX77o57WV7SR58ApntXSk3w
Y/DsNn4AoaMfNGBnbbQocw+GmB073XoX9q49pTARoEwkRmcFcp1GJ8gbYS7C9jei
qcyxkC/kx4cpytBSpZcmuri7LmPeP7lITgqp0uJagj4NSF9cr3tq/yk1QpkMVpb6
1W6UBzCj+VFnF8cUeL6jOnwfc3KTe8XymoaLBA6pgODwxWEZjLV8Kv4GsqNIl7uF
IDRfictzfWqHJTLCBvoVgdeXLrWKw1FUwdq7UtfkzVwpfTO/qoZfjncVvOvQIXmE
PteC82MSiQRHxi60EFv7/mWJ9oEaQmIQSPrLRl134a6pYvVlgPQAQ86R3L//z8VZ
9mf7W/eKVXQkXgDM3M5VP7qkep1BiJdDbc+R0MQZhuhdb5PNg2N9pjm1dWFT7Tc4
/rvCbg2p6G4EbVJ9/mZs7tyNVEIZSwI/Qo0BLUraFsEwpGDhkCnO9+muOOEwfMEg
vCwHfbqKjPRo3jnuoRvM2rg9TbFdFZEwuxJYA3ogrT3isbwvc+hHBc6LUYd0wbrn
cg6xDYehL4jXreG3Gy3tV8H02/yvPNJPDbeTf9AVqrH+mcLpyxmCffNM9ZbBTFSK
ef7uVCM5nsWgrL4qfZEcJzgtD2CLaXi3suwBh+gaEg+Rr8D4RKNoS1vCe1Myz0eq
hrFjB63PDdO9/99KHNJUn4SPfwPjnaMYuBRydHTrQUsrO3sKxCm+eCNkB+kGCt0r
JY0L/POdeKMasOenZSMqKaarzReZhufgLTJn3NKR75k4dsPzW7ZBxMwjh4l14mmG
BZ5jKuoJrhlpby22UPWzWUKuMzLwVCLEShOIzQfpYUG3NnBO2L1hoUhugOjJDgz1
vEykqTthbnpPc2rld3sumUCNoOfPQGq5XE2vA65j65QHI064kRB0v8Mk2Ku/Y4yq
4nwKzZOJtxjvYwwUy0v5aerk+jsKOyL3Ugq4qa5IEFeRF8Mpjm2M/yE7GbINhbeg
UaNMUSF6B45nj7m/3bTdF9BSJ9//AFt4K5XqlkWCPgvtx1bRaCZHYSAV8o9gCkli
vEB+Wmj68YA6oCyQs0Rxyt2Sxvn6MaXGualrZmkO3g0oqOyHLRBHkPx5RVfIi7gF
pPeDlTEkNstq0fRgFcI4e34LqJTzGznmHpgZ9R+u8aJubIYQL+0C7jipjRy5jCx7
4XGg4/e9bO42xkjj3Jf2HuUMndwW2i+Kh7IjA1zGKZbe+W2UJjuSWwhhpmmA12jK
CZiIikOBvdX/bt7nxPF1CYjgD6ZKWTXosTamfBYrxOrX9haXVXL49ESupH9Y7gd+
RR/ldt7WSNxiQONRUlAQEfE6IOnXq2pyNpfG9kJ6keqbPKwvmIYWjOSqPl/sWTH7
JHGSHrm6qcvLPBCI06hXi2bhKfpvrJEfUEoPsgSPng5uaZe++hEpbOuluweSCz2t
QGS9U+1NIQRUrbs9DHqVHhZrj1/xnvp2FJCnkiIKoZw/aYaeyD1X41MjpxtaVVpC
InNRGEjMhqRllbixdJmoojacHEBWHEK6iGqE02pzRYQ0xL9cEdY1zCTICDuhMjf2
Kh4UpC9g0m3iwA2lJFVwEElM9HieauciKs+2AOYHBbnzacITZtcb8t1mOnNGlN12
Kn9Cf6kg6iFg7hHOPq7luvOfFodhQMHdZvQ/SqaXLzkdVaE8P7ym8yQXay4FdRxg
mOpHVA6GlbNMD0j4/BpMi9AjoWPAqsOIVFI8Jm2cM8CMAHe4sGpkpHWAb2pGx0UF
ceC2C7uZYiMJJSv+itpJza/XbaT46iCbI+YPpmgHKkzIwC451Ga6cB8CsQvy3O4+
aGxSl28eaJ9cbjxpKUr4I4AehSaRehO4OA181QCg45iIhxE0qLEXjl4sLCme93Co
ag1CShk3SmWXjjravOyfn6f0RIJdWZQyxOqEmszK9/fu4vfpTXKlOa0siebVcJca
D1u9qcouJ4JEyyiKz5Da+AofNaOVdjw3XhTBOT35OYEkYXPJLCY+nXkKGgcpFTsF
0jiKC5MbKXv+E6FOvXR+E5R6aRjXHTxIUrsNg755UJ7AyUk1c2BMJNmGkKBtLVLT
Y7gDH3T7AWa8adEkmJtJeT5Rq2dNHz0TEzDtT/0HRmkdxlqs03LjQGk0IWKGTKrG
N7g2M9XwJCt1sL/aXqp331Wvg1aMZoQSP8D7MG3xSBICEEtHr++YGqmD9yMV4B6R
XeJqgo6rMv/JaNaBMdgXJz8J0JD3k7exoKYaahhKIvID8httLcVRBOQogdDhAnoQ
v9+OjmmJnr7zDqqZXLqsmJYXf5rEfZ+hnkDOVzdzd7fIpXahAp3iA1qENd8qzQBg
aZ16Jt9QQnYywVEWi2KZhcE692xgIJwaFzZy187pE47BMLrN9oSK55PUc6B0sRZ8
fBiwoXAX1ATBYG1mxRdNEnA5VqNWX7a++deGawYNPIsiHAxgACc6wnYFRNrA2suz
Hu8rOZlL5midOU+UK4M8XNLE64Hk77LaBNGeTHYk8/PKDhu3aFfLrkG64dEX3DFo
p5dkl6lZbYiauB0eyYXBrGRGR+FGW3v44xy3g3v6OBzXLW5UL1ZBum4vtkhrJMRR
Ehxy56aFSmZA969M4Py6a+uzk3BiNK8KTvWKoBCJvAyYoZAZ7nmuonmd9qXS78EY
AHw32w4RNUO+/oPaEgCdoidmHt5Iy1G6cpwPPIRd/p3BA3RRPn5dlx6gWo1VL+uU
ydvMAXzN4Lsm+9Oujs7ksU1zsIdUE3Aqh9VsY5RWVUN+irSsfhRb4DhQL3RkA5hy
0vx4XgDDyn02z024M/iDHPw5HRnCPGDFCd8/4MuPh+ggXS/z3vxs+efdhOZHcujg
q8/1V80r4YHcPe3wMLR2LQSvjLN0OIaOJJs/kEo+h2s9NH9xv/B8Xx9c5SWSh0gy
xp8eG/gadw62kpHUdIAGApANuuLlC9qPPm/kWXlgWgpLf2vRbYKMAbQwbbxxMhJ5
6szAPuVnUbsJBQaPbLDGDN5BZ6ZtUl6AMJ9v9S76cWXTsXQihAKQWMA8tdzcQifQ
Tv8tbodm8V4Y2i42Y43gGw2ZGGmnOdMyU4ptzC0JYikyRbBJQ7k0WKOfwT7UCh98
M3St0HJ2xFCXY6vzk8Paqry1atds4+FLgFYbc3oVDiCdJHhoqAqgpcOZU3W6mq2Y
i2bj6WJztP2Vm9GOtLlaHtrrOoYOiszKY8yaEJawOKCAmxpwHaoOzYiQCuwP5JzB
M3Q49bAVuRepm8cWeFYirfz0FEWBYEMsp/erxQ/Ngw7p95X2wpTdTN7SJFTYTU6V
YiuJcfDjDwm8mDVpdtabDByEomdj9o56Untr0BJwF8818fjPZsyJm8sQlgBkt7UT
qIg2MZKrr2rfesvSuKj7eXC6C2nbmxP+a5INNceK48JqPq5aYWqZVLStT8UwXLGi
Ym3WrIiN9pZkCpUPVkcwRslw89w6ub9EEEFEJPeLyzLsq4Db+UOjAeMzllGrE3YZ
Ti8Qp4/FhksXFaribFBRJGH27xDgz0jCh+z/CE9XL3lbrQij7rXVsM0k64ZK8B9u
Zx46pypd5qw+U7yr5II0yjY4IrN2IrG/MZ0XgZnI5W6TLdzTc7Nq8+MfG+932jxv
K1T03pmVICgCwbHNuerJKztADb2NPi6AGbfvbnDFw2I5wWlXbMEQh7QMXbPoWzeV
r0zm31g2y7S66FfZB78PV3pyuSTPXaBx+j9WSkBPIk+7i2GsvbuBCTAH8EgRZZTK
+tpAv8PwqFVB4tA5t9I1zDERX7czpNVaC++q5Z78MX7KyAiGj4rLZjRRI8L0L8RE
xRMKyPnKGggNvGRgfhhnOQnkSd65srLedfcuK4EmCQhdBGluPPvm9apO1eZ4yoa6
t10MqLuOv/ZzD73ctJ/2uu0aVO7jkddGOoXAxhtyHnITcsZudi+mts0YMX1YVNrb
+LuhHR7HUUpTQGbubsPWASUKxFGeekORsswxTkDeSjo/u4tIA0/si20MgRiQY4Yk
xl3y/7lmXdew7Y7hmyL3WssePkN9CJhF3yN+qi52+pNW3p1wkTzhlWRUMWqqk7rY
9C8UDrQGGSaJMYKrLU5gSwaIxyLSyYV0aqDiYK50umXoamk5NEonOYhjTmMgKZBf
8rEyW4sgJ8y0m+qVMRZzVKF5q8+MkdgkmKVawIfd0WNlJK572k2jgbt16bMVaRzU
h7VNbfNz1AO9HuQBBNFG2ltoWstWXLalicIItcfiXPOi0Dv1Cmil71FPfL6BXyxp
1cpL2P7L4C9a3+3Jip8cJgmySxg03oLuQWsI0q7FOyLr+mW1pluccoX/82etD8uV
Ea5JFn2/v0Qhc2+urMNwX7imsy+r+ZuIYABWNo2pUmZ7CMqnFEjBPGPuc+0RAAXa
/Ky7UZzcTdb7AeQJOafKazAEfFQo5t6eL4+41VPG8bail+miU/i158e1ZUz4FX+S
CRnsv09BIFfpB7xiiuIwQPoGErCYGx3XZdjReY/8z8lbDAKK7osdOYmF0W6ZMS+X
OrDbnJj1Z0erJyJbthpkZFymgvoy+5i5TyvePLKzGMDofj2G/rVKK4PFWsNMZ0jB
bRmbTLkIN2eSZF8WRkrUyRq1Z7Nnhfnyg1Qe3B9iruZtl5IZoUoW45tyhQRlVvzW
UojzbdTYpavf4++vh+bkb8x66ySsLU9S27i14cxEa04JJn0FRpmb+h4sYf16R/bx
sJkXxYLOMarSleF5yajVHuczL42QszvoSeXY6CZ32lIq/lY6NvM1Pe/dMjKutw9M
bGpT24yxN5RvXPmWn3WWXYQuIX4Fz4ANuFWlJlHcYBjTrsZsg379d4Ta9Yb9F7fP
h7hjgkrSfZXvyEjcz9BNQ5jb0XTmz/O0Is+Pv8fBpr7Vutvyt/DigWv77tHgOt7e
lYUbofha1eYnkaSMb2Fs1ysxfwHxZX592caVIyTaw3uYwKT4Fh79MHW48HyxZ9YY
fBMBWgjWlgBDeY8YvWaQr/BcX0J9d9PdZ3RJ943v7IOf1lMBxDyKFMO4tBrOinGa
v4j97OA/H4eGDKLxwiPtd1VeeZo+MIXGop2zIje/r6yHUV8MoOCXWelBkjCLQcDO
+S22s4GpgPybvXe/HhBfRaUln75c1uAygo2uotlXidx29qgJDdfgMunKMW+b44sg
u191MWcyj+V310/5TGq1pOBhY1BITxG+k29qCxj8TYiCYxB5F8/484ONBONmwsyd
sucxyZeu4ndnOMOBhbQKtHi3kOJBGLvwSp9cGh0UO9nojyTDwXkd94ZmIb1od8QB
SOdKHqtRo9aITlyHm+TIkLVAFqMg12w0KNfTn2z1WtSuVq3zu37RcJqziDrBImST
W2iS6MTSPly9GYUq0jVZIVAu8CgLcgJ5sfGE9tFq7gFmXTUyrXmeFZluVQehGjs5
Lo+gkgGD4D+3qiOhuY5onZkHT1tqmlcui1ScKqcqrMwYaYF3/HFrm60LUQ6rJDUQ
SbwhrdKr6MAF3eJO+9P98S1zFQexFHTefzlnI6Dgio9R2NJyYM2p0jgpvs4iiZRM
aWLsB5ogPqzHA3RBJOpptw1GlkQwjKusxKW1vkdeVtQxuX69cn4VzpHmoAIczR9P
pz5Zq8dFznYLU8phXrVM583yRA6NsTgW1FQTX2drx7M/8wWdrgPFGLyivaIGKkOM
fhYpD5wP+5j6O9RaIvB3YViSCjjKMSNUJTiymK7UE+YmBbpoMB0IaiEvZAaxiQKR
Fo+InhrgAxu04wzYBAbVcF8HL1HPiH1+NWIXldiRmcN8AvKwYPPyqx+8r3sd0WBm
qk6emKj0+MTwvf/a3kXdbRzV3qHPPHgSQXQa4ibpFs6MuguUcra1hHTcBjpsvlsK
0/isS7ngm4z5Vl6L0A+c12S6OKqMVuXsqyDnUEu/3P6OQXuNYYeP2HQJX2VuI4sO
BKiYIGp7rWoR9zCNkslCyxEb7Qjl+tvW52KM/G3VrgUj0i3J3Q2822fuXJxGsx2o
ARsA/QU1XaicK1H4tQi/bKQ+xMKsSbPIJSWZChxuJw+dFEDZrVkMUtrSs3wi9BNm
YWq5YiaB1gTd8mGTnW7mD79DkqYmADN5sY9TnAxWfVWC2Jfy7hH+rqswXO4+mHE6
qRQyyjJipzV0eoB5XUZheGzBXlA/9qRinfYruiZqrqaNnwOeMwn8eHfycKA1aJgf
qGG0In93w4Z12C7v8mKmAB8gLZAcVIZsfpmiRHVnvzM4V33dGs9K5X3ojXlppPdV
cxZBXVlfngbdHHFPZoUZ93/AjY9rJBMcG5k6qptVCL3CboBDCbKYXeEh3rMVTD7k
FUgq60tpG++IbEuvm/lY7bHqPMC5dQWx41ICl4pFN+tHH96Hb0NGYKBKzn7ejbyn
gifGVy7osIxVCxkRRZhHjRVNrUjcDigmVxBYquQkguwPncnU3jSJ0b3KkVO+77i9
E/UmW2laBpCgniWPC5vW0tDG6fPSOfnZx4Vdcoedx9SEUQC24Lkj3opqexEM+pPV
NBCPhv4zicFXh0W4E10l9hlgldfnUt1M8ncvTLcEd1zHS80Prg6v5WvE7l918t40
A/aHq7WE7dXLvUm90Lkcin51TNfTufW9VVoll52k1jQpPt8XyqD5Uf2fVSopCute
qIGgFSmwO0IotDOBDIOymTUnvL5LhdVA9ILtieUVFjqkMdfyim8PzIMksOqakhzP
Wk1RxjAwhJhR+Tbm/x8reX92HThJ3cPCdQ7lmQvv0EjhPPTVNalAlM6049Unf82U
9uMJUa33VlZbj/oyE3ALUp3Qw4mPc4W955F9wu2WcRs6I3zeWKa/nYCTksQMJ/pm
NhxKf3Uk4Eb0i2k3Bs7htbpAMZvDDiTux4+Hv6mLEe3q1KZczhIvEyUhVJtuaiVg
DAwCdmv9Phr6tv41KgbVSkK6K39t6tBnKaGNFAivLDNjwD/Rs3Y3I3QC1W3J08Hp
2pIsRhrD9yX3d1a76goz1Kemwr6jIKT60IIupqKNpPzbgPmXF+MD6hvTV41ehQnY
dLaPInOxBkVPDX9AU/7TriZjXmNOAvt7nIPv56W+IcX1GjNUJgZ+5GbPt/+oWpHb
j+Y8nAw3TuwKbwsdCuTjYKmJaaS8o/qSN4c/tNCwARdiiezSudDshR8GEiSjU3AS
K0gBQxsFp2xMZT4TVXj3TnxT1Sx52p2exm6+Wf9gzQxjw2GP6tvwhdTt5QhMFe+G
7FARdONDI12LmfQ3xTCLTP0LIJ62yKmyDiI7GySFBb4E8m0dVVgQovwBeLhwW+0i
scEljvs/eNEbqQnqw9wKXbj7XL3QepRhVndCCd/p/UgPafeoglLN0zIqYgvlkhwj
ir7171ICrL8Tx4ASJ+mwrmUf7KQyLFbd+Ft/j7UPdRlJRSiYCfeDM/DBhq+OuKxK
HiN8QkKUslQyXySQowwUAMyv7Dq7bBsPYMLzey/ssKRP+I7RL1JZ11y+PqUSfqtw
3opXetXTQMdeR5Z/4YghDcZJtAb0RUfS3ixz3optG0g8ouwjuKctpYvftY94j24i
V9SdPG5OR9aP+W1cHyEbiQATt1swR3iv+ESsQ8EDGl07LGafwukUz1CpNKFculbj
pFU8HQseHsYsKtatxO5ZwLS1bWuKKzNir51tm89jf6+b53UYe346mC6IG4NP+yjz
Re+KI+9fOvmaHFmrScvLHMYCVQSd/4VFgBM7fDpqtRBp40Cf6DT0WYUdPEwJlgTb
Ez+rZIrqh31lZUBD7WilP/5zfKs8rxB8vu3O/lwohPQzHVOoH97Ddg2znyCFRuzH
Knszd2JYXKKOP4JqALrDAk4v3IU5sVKpvqqKja2oaha9tJe/Y1TEOyjltjyC90O9
dQ+/QaVvJ+ag+8L4jqWsalBuVc+1JL8Q5m9HOmRqfgCQq79MnRv138Pwc49T2ryO
ukqKMmWSXdgX7IUa1mF8w1OzInO8GRUdrMbLb/gJExCkXwJpWQQyoIxe4uGObABo
30EgZlwn+UKkEf7b0ZCpoOkWC6HxSQuHEHg8KmF56xZpTnpdHWN4RYdi1mf8wg9d
bB97RomEaBMNTdfaP2Rr8eeJO3fuKGfBeqhTfH807mbEI/7fD2P4R7i/gfzB/4iZ
czF/uzqBiemZmxiPiHhNbFt8kuGXCipDDhnVBgM0dhfRX3McG79j/halTDewjjDC
xGJS4hhm5yCwUSic7XSn5Uit8RG4QfR2EhXnLl0a66vVbPIl2Hsg54VrtNj1pTMv
HFF3XabzIUKASvbMg35gSjhJsy2dG6LXcY+kHVSsoV7cEHipvfXXxX6UDucOrHBi
bRis9zmJTPdh6Js5aYLZHr0oHsruNXqktWNPHBtOsh/kpZxBLpDOFhMxvln2pJum
mdknRq24HvavlvqDONMoS+ryNs/xUnXGDdsbsVEJoYw6KmbphV+Q949BSVkEoEHM
Ulf5Cx6NDQxwH+m+iFC4ap2PXMTzMFaomEzHXhzPop1HNv/ZOcFZToSVtklhtL/k
3QTEfIZywk1jrj/dsInek44dcEr+TcbXlbxXya3KgDjVq7LLOx9fz7pwZoNiv8Yd
v9DYiG4Mnc/jT+27KPTlgpAdISGpEt/1heJbk/FonCBtQMUEWBfdJP6VjMvy/8Dg
5FH46oPp6xH5MFoVnpNag3dDQvi7KNS8AC1fmVAIYcYKs2enVaYO883kfkh+R86F
v5Y734TGi7RJy0mhU7Izva8fjIW6DpZzNDPZKUBnQ1HN1XKMec3CNbW4PPPKgCpX
GWbFFobOWoH/HIK21ulJkqbceKTOyJj+hjmtiOcpuVeyKl/doxl36C0dkwdXvFt3
9G1i+UneTtTNmMXWHeE3fgSYjaYJSKr4nY1GW9GDXwTOXO1D+OXuwCxx+iIx+0/R
snUMjIqJlsIYpfPO+DMHechTqNEh/S6puGo3QNQuinfMvGWZB5SiYwzl+zS5rtzY
OjHrO2XMsjdjoE4ipFzaK2Sb/KjoUAoKfCiSoY/Lzmzlfvn62rtUH0SVTmsUJ8gg
IbmgMHZ58mUY7EbW2qHydQwWhDopDkeAzgmWpQXZuOKytrPD7LnhbbbX4krfVtWX
4hSZvuNu8fZEORvC0tPPaHSkV2MEn04NghEimsk2P4qz4L35/85k1bsyx0P6rye/
M6z9HZJBAdZN/Cn6Xg1t8jcD+ZFSpLM0/oXEXJkIjs9RpeF7a3PXFc9HUQ4nTmnT
mqoAbgDZ6VPZgPJIF6yQaC7XchPeDFDCpxv2tOWv5BFBXPFxCyFvCa8T2ACUAlpi
omRDNYW+LasCaDgTTmXxkMcb0BrTT7ip7l20I7NCci7J89SjLpmf3dIEO9waG8+c
Nik6uBBi9zzgf6aDRLJrVhxixeseuyua+ToIeD1hcv+DIou6BkeLsY9KVbBkW7D4
6YUH6jBRhReWUBiOEV5dunYN0xeTiretarTSlpuY6FXWtrDDJLXfuMBMebd4Fs43
la+mC7uA866vftYnQVIyFUqF4668xtzOWtSzU6NpW05yXiuVXEf5cuvAwHbwO3Cr
iU7jwPOcLBvwJdPqf77bkkbKl2l8iSN0PmXAOv4WGF4kea7I1SHQLqnwhTQXgcZt
LhKPJ1Z72jkRbDqVlyHGgxUg5pTNduICpQKzXLBUEtxQGviEv6i7tE6Yb4hXukBb
URwBivQEAbCASf3XGkfHZixBZfFy7Ew9Lp3TTU9zdVf5cYEE59y3Dho+6UdX/TpU
KADmlAhw1KIyrrLmMtoEXa1zDlDEPZdh7GPZEUvkW9kHSlrkAqyebwYvLyHP7X28
vmfJwJQ1yGNnzl6vST4+Tj9Pm6EbiOyHDsC6SBHgvaEvR40a9TVsbGbsYPv7gyw4
MklVT+uUFhP0kaqsbBjVIbk02UEt2EKvPur0q+6yjr4nOKRg8c9EQy1HM7I51KJl
8bx2OWWRZujoQhG0Y1LplfLlyqjAhgr14JompL43JVuA8o+3Ow2mKdOEoZaxT3Eh
eI2QcvQuGJ4G7UEGGQ2k6+FRD9v5qInjCGerQ5fTzVlulz4xDS7wroTz3/lfR82R
qna3dkzGc5UtrjcFzB1wB2rqeJkKb4KD9sLOLozqhYEuMbM80Tk/TPcvByB6xw/w
u6RUrLpEU9M/uWvXtw1VkFS0oK8zxQGwuaxqMHo+LFxD4j45Nc5dDUTfLX/mq5xY
pFS1ukY8dBp1gkC+HB0qvZam9IotIMzeh7MqZuYyS+HI6x1F1R0zEjyDC0UwdEsj
1qEgU6+626NHAvz0PTRfE/+ywQXZHseykPi4AMaomFP42NY0rRiuVvoiGUpBCuQh
swH+x0X9NnEUIYfVxWwr+SL8mWzI8dQzWyMF8LuWy3C1tzvSeI/P2K+dj6fP4QXz
Zc8Z8Hxtnlxs/rg5rEz7dcoy+2TvvSVsnAmqJ0K3Ai7IMpvZDp/oynzGS+AXcSAg
jmX01mJZytuLpIOKq5SpUVvIw91M0ZQ/JGCmaww5Irx7I9DCfKDLM+p7o8hTYhgQ
ZM0+iLBLBrtnNhNv0K0CjmfOIWuxFcvaeCic6Y+vepGpLFCmBlEdcMiZ7a5te+Su
65zASU2spU15EjvzUXeL1+tdZX2pKZwxa6fqTFb+w3kZjqbb8QEPh3dePQkTnkcc
HMFSAhiHu3mOL+k+A/OlDnncggUQZZ2/f8R+27deOKAmX8PwMXMgdhUSS64wVwWS
ZkyNzPdTZb0JoKKmgMiVI/VUOrch+S+dZqyizm05yKcSqPPJubhMBT3Ms3wsVS0Y
B8b9i5xkJiNUXdtZXc6mUfxQaPdhiS8yTJ61Qd7T3SxA5Z2S3qhzf+fK0iz4KcSs
k/E0hCnOts81gOOwmBkZD1hy69Mk9ZOiYrmU6whKwaFAmitlIJ9Kth8bFCAgZLIf
qVuoxXFfmCRA5Vl5p2PpcJ2Cpp3r+opRNCCPd/g7iy1imTcPnMsTvI3SVodUU8p+
FTARtIrLXQzVmyJCgKhRez0HSmcYHiDUUN5sCUkn8udIBd9GgkHgUzhiTQFWluBt
ujXxX4WcRp754iLPZDRG1pHAn9SskUhVbPZjhwxnt+cSNIncuNv5qk7as46hNXDv
DpWEB1qkWnLgBlFlCxc31q0RwQsyhyVDB4IBAiN3IPamGZ4IQjYoy209l1gLlHlb
S50n995dwydtUB5Aw76J7+5n1jVjGMdmmqe5ih5RAO3cufcQJjizP+vJOFSMVumq
I2C+IcI+TgqMLeNg/3yi+lyqEzknrr0dD3vBQJZGVnMBRaQZqEVkQPYzig+SF5Ur
YzL58OaHdrQI6r8sDLStIJnAgmiy7fZ2UigOQKhdJSamR+ISLXN4VG6Nk/UZAKrO
XsrQQJl/4VVsnHql5rFQIm3kDoLEPrahJvP37fOR63W2dXNxnv59A1z9zdsShk+Y
gfDoQy9gua0wyhto7q29kl8LAGonHpv4Tf3QMzwbJ+7ZWOPoSKcakRLzuMPDvbmb
OfGYKAyC3jgkoumDcNwA0on1ZqMauc+99IXqcT+pyq+zQPL0U6tmeNopY9cDm4tA
hc4oh5k/EaQ9rPKtjY/aUnKEeU4nt2EXZegbq5HQFspxRLRFji67kpFRoIeyj2xV
zSSWULn5+phi954K3e3nva5B8RDxAfgoiVpLcivWGIW0h5aD0mFDM9+atRDKgnv2
C0rsEO9WUam2iBmpUtyrMQLxDAJXioqi+RZla07Eiy8MuP3ol2ecjU/c/BzL13oY
AC4rEwLezrGNurdXsd52YkVf8Ag4w1ZwqeOaYQePrmbqf7Kt01BaQXSOgZWDlIhZ
wu7Q8FVPgftxwId8pJ4d5KMrJtIJ77SsG+kgAVnwSPL4C0ZtB2RDAB9UKghReKvo
AHGdEpTwS7JYUDcm9BHvAxjSCfdqctkRRN2tSEXhBeNB65Bpzgvn9GNhlxWPSpVy
Xb8/uasVWR646eo9alEopLowimO3eIDWcSB29YxilzI++IWwuavq692+pnDkvOUL
xUOtHvKTEAI9mkevwhLqV86WgvFPGXjjl6nVeTEtpI2konloBGja59/xrS16p3Uw
RXErY70s2IJ5n7fkBXQdLoEoexb300k+IizvYtFi+aRnok6/0B1UxTB2RzQCzOM3
A3rczlFlqZgigkqXrZ3bMn4fUblB9VnUbiQqQQpfDXD/aMEcGFR+2UI8CJiPlvMG
oiSvyQ8nKi93HUzoHCtbYvUmwVr3LqSSdJyb/qxQbImPd3LIS7hVVclpXJeS2u3n
P0OLy12GEfcBt7bcW5EEkx187XALuvbeYifmVviHbbnZ07lTdk46RMsJ36OBlqFE
ye0R9WbCYVA7RixrLVVnEFgcODvs4b74kpUrAlFfiVV6sc8F5+1b66CKYBf4CmHH
49AKlQI02aktalHQKKOVVHK/3Vi7kn9IVTV6CFD9ogq4ZhYh22lLPjP9846cpv26
AdBS6tKqRsRGfeQeD2wBEJLYcROLHouP9XOH9rCY8KgnHuLjuDwoOM8Ik8B2yrTJ
lkiGxyG+1UWjt6U3Z0WJifdXV/btO645q3Lu7eKvq5Ye1sb6mAJ3qV0qxiJzN2F9
Y7I2ynkFXhuIo4FC2/Ivw+6V+e9mX7x7VuLWCp7WbNzgTS94ZC/eCV3Nb1kOhzQm
jBVNBEpP8SohXdiYOgutvN/WhpWbuWnV1MQWnTcKDQPEayZIYYMCSlvUiHPuDxxL
RE/1v5sq6bc03mWrIZewldYVjRkW5ZncKdy7jV3+YaWc6djITrpzez3wlrFm50TV
v0/u36e6i4YNoKRbzrlBgvV0S19YqSzT+zc7VAH+z5sXQ36uiTALnoPWhECHmdP9
KWTm+qbN055hKm3d03kP6Bmu9oyPNxcGsAH2mI0gq1Jj97HTAdXVyNs/fK3hcPXE
4s3NB6BcbSzZPu0u0xNtNJqyyY/sG/VbHQwImtt5qEdz5LNkNc/NeRLnxbVCq4VO
YaRjKOEtk7cArg+PgJJVVkWI8EdyqH1ehcNcHsJUDmzqrCHwJ4dXInxbi09kytpo
fFhDXe+kthu1sLywMct5jtWLAKwwabKhRLT7A4T2RuogCoZLBKJbgfamgKLBZN4I
enziIXmBOvvss5fUOYiEYjyq9y0gdRksTNS6s3KRbHuKYdDGCQyyl9xZ0as/2Hyo
5TEpsMjxtUxiqHBLoFZ8SOK4Y+c0Ia8OCA6VRBlGFxvGApsp8G9X+t1bTcho7VNM
hJoMoSt4leRYrGsFdKHwh3jw7H1wQZ09JG5vjZu1oy1YXWpSrDkFkUFB85SEizpY
ff89nOe6Z2/STTNBUmpqo9Q0SQH4LYUV1ZVQsNJADfcjyD852HRFihS03cVljqt6
axGcvY0fiQeEo9dTb5j4GVt6KDH4aEFLHJu0w7nSxTnwsktsw41dGCGp2mXcHO3y
O+vsuoswv2ZgEGjPUsisB0tT/2YwQBKojR/1yda/1FXt+PsnvICI1ggnr9BOByPd
bH3KflBRZT+I/TSguZU5+xurKGVGqgVzqVcqblD37HPZfr3hTInyvQI5RTHbcK5Q
1G6P6HntLv5Bxi4tNIwpF1Wa3TTJHJWQ6biLwP8IiMzq8nEwRhP+zm0awOEI0Mb6
5M8uJtSUOO89Z0M3obeMS8aQGX/Rd5E5PhzwbBBFczXbOjiO2EEcjhvrC71c+9gT
aMJKvKGYSNxm2BfF4wqgolvMG+gE8TCn9qr0HJsVvvTQtKXNK2JgRmuFt6vrs2ou
3Nfhjuxe2XTcBE9QN6CiCvGSiutEFU5Jyni8yN5TZt+fpO+SnYE0M4SbUafWKhCY
AULP2+7Z8cCDWGdcL8XSsqTl1bTlsoYhPLzlP4l0He/SSKr0+mjMQwoQSUZAja9W
F8fjL3P9eRxoUHhHaiq5uv+l0W+sNRMnVPUsuMQT7zAquCUe59Nk5GZC2pVPRtkA
nezqp+n5/Xyda5tYGvlNjDZ3/9tR14OdeWPkjS+kdT733gh/yUIsPS1gUtCJAddJ
gpCPynXUQJbsQ9YEB1o7n8NH+NnujuUlkeAcaKK3OcNFRZsssuieRrRVy5O+Fyzq
SABbbWpnwEXeH3v1XxW7//CsYaA5Kb9xV5oGNRU8JpyfKWnioNxRRMVCCgY4c0jU
O0uMXmuSIv4qHpuzdnYeos/QX290UMASQJFGxm131WFhOUpVuHGoA2ET7dYhr1Fe
3W/JkGE+NQbtYwwRELb8Gyp9zlXFDW5NGM22A2FtxOs/K9805w4IhrQnbTZ1Ng1W
WI8+rraGWJ/EKDpJTOm0KVaDutsP2T8X7tz7z18XHMeHc6k6t2+Ksb2HwnJGnVyf
X1Sru41h1slrT/+0+wFLdYcneSpsAZzFn21X//ejfTMaX+DzsekxMAkkT1kMNAmB
wZNlWMm9EPq8rbJrCiHPlUTNq0/L2VuGoD5erkn4IqTbwgBKwO5IrTgneymmo3VB
LJhBQGv/sE1ZJgX/12SAakVM2Ee/VHh2R3Npfva2WbYjg76gotKHc8zlyn/GDWbj
6pXIHlZvn4VzsgZPi+iEtKNhWqsjqR+hILD02E1XiHbIAiNtnhoDjZIR/39p00x5
LMDd+0Has5xmO/d78ST4rg2IJOGDVZVZci+KIdZnGzfQRxhP6bJHqON/hiK0tpNW
KB/OsM0mipxwkLb1qgfCQoTZME6O7Po2ZQfF20uFDIN9A2Xs0mkQd13z7qOZPk5C
giSKxr1KEvrDz6GPStTKq6ZJkX9B0Mz3BQs/2Z0q4e53966HukIDnE+1cf6QtGlr
RjyYqmPot4Eo8XopUIDN63B6GCq2d+VPb91d3D0+lLKzhYVuLgPQyrQ9w7hdcsHl
b/o5a3HsbkIGsWCM5pjgeEep1yft1OOeikauZWywDtzVES3b7OwHYCrgaRJCdR6l
Iws58o4QeWP2+MGyGy+mC2qfDQ8kiklGCuVyb/Su0S1yW+PE7wfsvArvLSYKStiX
I9jkko6cNpHFf8xmnk3z/aPbaOOxj9LzJ7ihTszyDgy5VXPn+uVy1rnpeIma/EJ8
jbbi6rbv0XDoxOmmnzEOyWOgEL6O9uDPjSY23We2NIcw8oGjRtslvHONF+tWE1cl
wvTAVvnuAyd3OKX0IwtWNeL3bHK71n44uLQoZx2ifZjf2f9Rcrfj+6JMYVKyfOfE
7CuvCDJT/jXtqEUFCfrqD8rbPwXNUFxyzOFh4Crfh9g2jSAomxvd/Iy+2KBWPmDJ
mf034AapXpShAl3Es1M4POlWLcduM/gNO6b1FFgmYUnD7CFlYfeKIHOgA9mg3Q4d
vQqZN77xTzKhNuSCZdD2jvGRTgnXgkRFS/eCnOvbCAGYly71IsHIkNT76/8mchJP
IjiVuqZmsBoDbeu0on8FVD/OIh1nRKG4QMDd7JIEjBcxO4hEmKCODKsqG+nC3XBK
Nu/pK4XXtKNIQ4VCDwTuNpO4FxWJXxuk31PWwTwJKyKD5fFkBAdFAaB09qPsu4Ju
0UWsYwQD/ugqxZzINNWzmpny9FfSuge9oE/3E9fnSf2hcRvCdSUX8JzWrffZlOtq
a5YwVIWeNSrHYNnGrwzrvOMUYaAjY6lpiGaDlmrD8szHMpZ4Yg9orYE2o+msIEBb
wr+Tzx8yyL5LlDeJY2g9+cIQ7uXNwMIYegMRpgBaWEvSXlx3Z7K7v2QqUbhZf9j/
yc5IruIbdkjRGIlohbpXBxXcFuSHSDzBQY2F5yipO0wSXL+oSNW+Ps+P+KUJzy3p
fcx0+gqt50ZyKjYYHyOlJIABCzHlSJgNWZFd+cABwDME6LEm8jpsC7z9ay4tr40X
NPAuGHr2hu0cxzNEMAQ+uw/MFK7pARsyPSpizCxNdrpweDfQYTI9wg2TbFz9c5S5
ziEYRUlTmCH+XsDI2Uao6j1LeQBaGrYZ7RBYbRIltBVSZ3FGj8CifkolgI9R8ueI
v+pQJeLlRarSpl0tUqSsDLSvGSYhXXq4hoYobGeZlBLO+32o7t/BbcXFYqC18aNO
Zhw2srqM5taJkgz4DHGX4dH0bMxRaXNspXWI5VLqaDGwmhe9lf+Fj0hN2EQiFy6k
35JIKwV0PjcPKVkYXg9v5zLEvBES0WavsK6nmuZCAdaUIEnreJIWbR9hSp+y3BZU
2UMFW/IASI2HCmR0kBSLoXLrlIRPaVIBQao88A8KkjGmnRURXZoca98+QJliqj6E
arqLo3G1CRwIvWLsbwFDxAtRFvT97QcDjG8eh53QaoiIHqBR4jH2rpwG/9qTpRGg
me6JtWVJrjrT7BYt+5J+vT1TAP0ZzMv48y3MpRkZLA/kvjXjucR57uu37X+qjnBN
UT3HnRFjuCbCZNT1ENLZ1wweeet7UCKu2ANhiMrbf33eOEZ2QkxjG93FONl8S+cj
3xHt5xbdB7UHqNVJwS6rfCO0TE/INqCMW2oPkWTi1Nx1lyAbhbuF9hIQrReRggTD
b68GPae7Du1QykxtH7EWq0C1PuCkcGz6zcItZvW7JAB47R7CPsHt36fhLf3BEYD5
mdGTQlJljQGx3n9MbLYrsHFYiDGxWx6M2VTfYTDgD+yPwvuCwAMxIODV1XeFHxMT
vpihI1hZrkRxgjkEqKv6qVsdOMaWLDZJNfhC3BfdULi774cSVhIvsjIv49ogK2uG
bJEQHA0NnYhFBYu6cNPHjtloiJXhyvTLT7cRJoies2KtuuOx/rCj3dPTAaUhrq8t
sr1Dp0nBoeHQWQulsU3TgH+DRsbQepMxKumsWB8xIXplDIrzRN1owcTX09fh426G
9yXrusyCHhxMg2vqWTNBM7ZHSfcFT8W/hhQ1BZYZGrn+L/gLxDKPpMTQkV32vrDT
62kVyGqaZZYN723XyZWXynWFuVfY4yTu1KwuDs8n/n0Dd4hcxCf7TYo0k4sdu5GG
1KRWIs75xcPfbFjMG4vrYGhtEjzMQqOppwSNf9GGN/Hq9ERNXIFt+D6nf0dWl9RQ
modQxJ32bP0NfqBObcAkFtWUcXBh9YjdUSpPXRerFn4B5oHayL6stQqFgparAGdp
q8MxzEtxB23JPnA4iIZ8hxwbLE/CoVwPoUxF+3GblCvWsDe2Hqb1SmWVz4JUQuyX
Pg42vMMHj3nccT8FuM7e29zf5I3nDx4f2/ydX/yZIAvPr3puzG1u9gKxvupS/yTT
PrJ9odFYYkG/jYHSvcL5YQBhKj0ha3NYlxAJHyyXqv9q0Y8vd7ITKT0YevFNnV8+
FaI3FKXFOPS5QDWqo3sV8VUTxq8151lhrdrH7m6D4YmZUxzVjCZuxa5XrM0ZS/dX
hs8je35K//fxAGMpG/JfJW/PN0BwIduwYZNKwjju/+o+I+xE8le++XYmQy0OSgC4
O27TPmVrgz9oVU0kSScrs9csG2GFYvRv3nHnL9vWS7967+xRJEMa6Da4ObzvX3WA
nTebR2KId6wjGxh/BaRoH12MLgKMKTqoWDCeZWRmqHzZFzCBx6eDJVPzylhuHwGw
W4iDwYv4QazIaBwbN2BDpxssE4Ts2oE1sIoj1e7LajUvXCBpn+xe0GTdMJQ0zkbV
Jz33ENeR83bOkFXAWfkL49bhVoV811QACu7NrVPQTBaLNFgK9LT6nnH5Ps/7Abe9
mj1/JFFHncOvFRDGpjPLDUw+EAeg5SbRiCLz/JAbsYfDSXDu7O0k/hmOt6QEGFyR
lQL4r/sKUQ8D83GZ3x/B1IIsMK7Plj7Eig6dTkJRrp9TLboRW0fk4kAvi0QDLHeA
GYgTqAFC/KBc3S8hw/7EG/GhVDGhzzPNwKqrbXmLIOAhR4A6sWaIgNiCF/uqOR6q
TWXEfLAXeImam14w9Vboj1GW+rrzdCTv0klZx7/iltfw16A1OoNe32ZQvHykWF1/
Y732juvc476YNmf63aYDscLFY+gxCr415DsF40TUPfr/5ujTNmyMhXsSzkgdNFfl
3O+cyBKdD1PSLyddjOK7uQXkNtN6/ERrDg4yB12Bbl2Qaf+qBmEWRAMWg+bVXRcK
zpob1HXmcRfE40jXKQR16F0/i4T4LIklUW5N2zdAZeUZJ/ALbPS3C6WlmH2NHCJU
LhiTK4q97aIr52Kqphyltcxqv6SX2TgWz65Hrg0ZmOUHA7rGSlixQxwj3eg6JxFJ
ofigtbUSERo+jMwfzt3RtuRwiapB3WA9ymsD/stsjBGJz3JpsOG3/sAp7wa5nQUA
OApfcqAdp8wQrJeT1kvtcwodZT8pQ/GRaMDjKFpjyetlPBRozb0JqFWZTtKdNFMl
geAG5mcWzAw3jTXdqU5UCKMJO04kuRhs0hafl6b8zzRT8mVZ2XeztJpYm+dbvyYJ
pAdEP4sP6WrYSvkCrtF2Nt+GU++70K8SL3NxUqD/PFpQLDOEIjjoch5QdAg7ZC9G
6Jm7uThtbN9oJ1J3dfdJU2rUbByeMiSOOinSg8h0E78+cmfQ7uyG97NpYouFVjTs
pEKvDi1Vu4AzdH3AI6zHY1zIec/AQurAWV7Ph7J+P24JxQMyToSpGk47k1XuL6t0
ABC+aH1q+aGu8FkrDL4SmiIeBch94CaNqONEoF57T2aiXnmlNvF2TR60UHDp5usu
PhRrnibDuZ1gMl3+peJ+7KD20+MNXGvOSpK90qyvfMATF2Fhl79KLNdBuhF21Cyp
mEBmQo0oktjUD5M4vW8KatCVvVjhh2ZLlu/O++0R4JP3d1aydSD6OxPBe+TrN8w+
w5Bq//6Y9MWtLZrlLlPyBFlZC0M4WCro3HUYKP+xU1GjmUmq8iD2xOYkG1oztOrR
zL8WAoBKDAHfOoWPHXf3BBJpjhy+Tc+tDzLy8wYphHBBBFvsH5q/Rd7lyLiNuQY2
/mjYhVP/63b2kxYII2oJ9rumDnR1AdKqoWUlbKowhIW8VFZONTEpWBdbVjLIWmmB
I98S71/LtX0tn2/rlksOXQ3FDVvQwsqfG09xtGfdaSyelwOWadCP78rTsdUbaddT
NxXMijrDco4Ym1R3evf9xEkLkdCXst8sK4zS8A7QyPsuevK/3QA5T8SQX6Hena6x
srPFDq8foiMyP1I7frx+ssA2rbFFOSkn17Wtt+a9qL/WYTcQOfnA1iQKK3LA+E7N
UK/ol3/AjV8yocF2bE++NubeTh9/V//ZESHYtGCygkpfQUEPC0h3qM/HzKwrpyvw
7+ubTwKvqT4s0r1h/zWyxNyobvn5zXuaO+G2i5IYzgUTDvqS8em054zKv+IvH4wa
iIxqq0pJFZtLy3j0rW5q6NgNy+HKC3jfK9YQS4Y/5/LjdR6Zhrp6hNCQLRBJ66S1
ShSmjYZKU7p/AiUQoLtO6CpWAQJ19bUvtNTqS6zzmKbVdjodFu/iLF5DKkvHRf1D
NZg6+SDMSeGIBgDkiFGcgn2Ag/LXmPAtFRhVh49RDIn5F5eg69yDJWW+hXDVbLt8
RA3fmebB0ZqYVFmzYK4L1IXioT+WPK/LZyuzLhfurxjEKxdYjjc3h13BYedmrGT2
e+gjU2F80tzHtbNQlZ89lrbLnSd2NPzWvf+eQzwEGG4PL7+RLOIs7FZY+FEPWUD4
XLQ5dcMW3rfSDBDbL+eczbSy9BTdJxPnCjKMfLhUa56RaPMxmn+KObNUtof98ELJ
lusJIwtYFzfbjXdG1McqW15NzoD6MI8ziw1bESGYEbQisW9Mpgl+aSgQql8dp0eq
3HhGmyKQclKguYtleJJWwIK0Po4YRuidRGKR4KjWkdgVzW8BriE3jPKwu+LtBAw/
3vvdgQUZozWsSiAC9c6Kwvg/qf1lzTn8M2x59mHZMSNLzM4mSqc8pTb0DwhVabSX
wAKUbGSeCFCo/zfqkC9YYmLzrPF8xRB1FxZGmfnzPmioNwWB9sMCZeRMEQQchecr
/UMjL5xL40Cg2evkpKAXdNl6o38V8350bFH31BQznpfBiXyVzVPDBJ6TmTwnsmnX
8xb54/wGpstzwOzuiwxC9cYmA+sha1gbsY33F7vJ2cwjTpM5VJeAfkEf/qJZSo1X
yxsenouHOgPzpu/UI8SoEQXt/5qHMqSoGSD0EbTpG34miKEZofHs7mtYxswB9TuS
dsOLbcIC3Vs4a4j4bo3vnx1wMo+D2KFiJ7/ib7tsAHLDJiz6FzpfSPLF7hNm/JcZ
J8tqS3PAN8kFN6wUSKOOoIa2j8KiVcjXcse8Wb5cFeNSYNIb4De02N3zRpeeXPHM
QP/bid8DRebOuT8yZLLhY58X874bMaWfoC7iOQhujortRaF5vB2AxvZjmZmsEwaU
ibnzByyMM0cSfLAHU9TYu+W3+3wixf3yAOKCNECpepJKv5RpJJrhxgXpgAILDReN
zjhOgHGuIGtJfso5YnyQzDnFh1KHMaSDc61NPvke0KBkBepjW673ZJ1w2CMNUYQ6
xkM/Iv8RxBEcAr6TNc1TeyKWcgJ646+rmcU1sD9hEKOWp+mE16LCYAhH2bs97JHE
6I4cP8WYEWvdJ1aQOhSYBr4HoyThNvDw/zn5oXmj5DN5NX47wGUNe4hgsaW6elX4
Jpk++4cNRcYHTjAlzk7v9E6ErbzwKCzbQcS9xU1ufhGdNkmOnN8Kh4xMYwSyqxmL
2bXjKx1unsLWsxYMXy4gDZrzB7WRI7czYCf36atZwkM5EONweKuGN95qsc3/mP0I
vbyOI9r6qNBfqsNSo/db0U8MnXmmvOdxlc73RZW38BxFiMw57Nl8WXUpQG4DZuai
EaUqpqDpVjFYupI9UMKTFiLPnkM5IadFGBUO4uITrjMUEb5UghDU1Le6w0NgZiHu
MJIwq0EHNo8+/AQIi5D3suRLBFVxIXdbE9Gzp3UgeU/xgomnGgLjqiUKf42Yk6nb
P9C4XeD0Zf+K1gV8RperDWdZJYGKJRpdT4wfR3GBC5Eb2sxU61VkertUBxkziILI
+AZEMKQ2oStDUsUHKtho1QKAitl6sOlx3TT1vq5t8fLua+m9qjJT+Jp3XX4kWW9l
4O+KeN93f8nULVYUFwXonSqhyZIces1+/9yEKZmxAtG/jL55CvEWd+Epj+NiJYRX
BzRo36pr7sJfLZlavY4YbwIgUBi2o7J/G+j7O5egSf9rGoxEPD8lAp9Fls88/0UA
sKTR3PxEyGLtsqjWXMdiHlrGq2a5UenfI/beU1q5GGxYZiK1NP+/i2QZFOQvehhP
og+DJrORUZr+bdSQ4L1tp1iaVq0s8bpxaRTKwS7q8Yv2FLrRm+8YdHxUTvUbsGV7
Il/EeeJYZC707Zb1eDrafWMfo6iNWOyrjssgYOLMcBpUgUFYcwXtFqJ5RvvMh9TX
Jwqe28mUoNHEHUdfhN0l4AfDAS47eAQSTDVp/dt0DgRdC8osfomkbL/70tYLbyKj
l7Dt3VtQE+FYmW1mHR5Hvn6FKFuqBaoQOJMq+S4KYaOtDySBr4QZlJxGyf3yHHt/
l/fZW23B+yj44NOL2uvZXFnKZ/gKzA7igsQ00ct138LSNfL5iC/dByOfhBLMkU5B
N6nXbuEyNQxytIfVVwz2swEnU8tMutR/cKrvFwbcVtFVliuIF7vgEq4wCnrWf4hO
sqhXj3pVa4DU9V6DCcMBudI2RpvQVqtjIH4KxWQ4cDsKGHJkSF51/2s0Dqt94D+P
z7IRoSyR/j47c+JkOrlh4+BVMgbNu7fzfDwFghajm95ph9ZZ6ot60iFpByxUomI+
MtnjtVl/nzxmtZim9xB0uOZ7IYBR8jqke5qOuxzAZJx63RdVkdVvkiHodhjkR9xt
FKY3tKRwzXV9RubPqUxqCpqK4uYkg2SF2j5RYv2Q1WPE+uQNIIWKYmCJEmz74R/W
F0c8CL1kvfSx4g/1dNcssbbFguWFFaFa364qjhIuBuyNSPmX9eVu8sqOvHT8uziD
RHkLy/GoY52LLmNm0+yYJI6iLumsHuwI19fq70nDWpifSMBeTs5fVg3rdEXK8NIS
yVgBDvmex/vKmK7bR1RMlwBJL8N5/rk2iLDNUwKn/1G3BCYQLvAk8ASfDwzIaJVB
i7lQXaQQWF5u2ABZ1XoKMlBpraA58dg1UHhv/kJJMUnEkUmlS2aT457MIOxbfS3s
2r+E2CCaS9IGgxPcbwf9//+LgCHDV3FQ46Nfuz0CMd6RpY2g1cSEhpTHh3HKEdvu
tPQgILNyKX/WyelMJIfZR2kQpIzr4E0ZZlHRpABaXWFTFXtIU1TfX0OUjw//7Hd9
PJ8G+u4LrkmlBe6ii21t4P+tmIeYMMLGWgloNA6ODQuLvNRNRvZPQUoFWDs2ygVG
wmeAh0dymeSfWzEB65j9ba3nn2LODdnnSCld9DH3NhGVaKugEgqOmpoAlm0fyADC
OctPGK/Z/tEPqK+RkAqE/89udJz52/Ufj1QxcQNTvp4h8xzayHWWZI0d/gZd+LuB
finbm9A5HAeMme4RWxjdPEp50SolZADMZBn8pvuTumJglg7SNJ3OhDhRWlX9gZ1o
Pz7ABvT3lZi246qJ+fXexVKzODgDjJWjUG1npzqZQmRCob+sX+H3sMdhLwnEe/XF
Q4Sci9Ru1sRQlaYM0R6lHZbQQV0ufXJ14ON6NyYiEI5NPPTHHRv5uUDDZ5Nt29u4
v6opGRK6ZSqy+UrgICdGYGCTrP7IM2qYyKvopC9NEzVA6Xy1tdD0QibOY8Wu4ziF
gtW0jSYelqdC2LY2wghjfoKa7HVhtQr32IIRpvMdjMAmkLyV+MUZh8kxnNYvAhQF
Tq7uId6YFR3PeRQngCs3gSnhKFqvcdVeL/T5VZXNEiDndGhUiG1pAcq8Ge+Esd/b
phtcBmf3B3318HCf8JlA0gi6CuIEuOaI9mG9aBeKkjPWPv/zRASUFiFBIJ3+H7Io
0j5G6xj0w9HdcqWykbXmJ15XzrgNPcIsnLNhWpCXOcT1ec2b5Q1BD/hxX/5+hmm2
ztXG572oxlygADCKxZkkIoQb8bJrv4lkvYxf+XRfQZldjIceEMtZGKOwK2I2/Ek2
ZOln+FtQIP3MCIxC5bzkZkJ3NZBqOtFGVIOjBCSNDU2HyX0Qn30lnY9jaXO/0Uq2
zEVNNy7YifEi8ZEeHNuQmF0acCacq40BZEUNtAaHYdx913hJed4yYQecP3nsFe97
DfPACwwrGLHYYflXYipO9KVvr79erNLACJgn2bZty/B4M7w05aMrcWlsqE5OgVvn
F/l8Jqg23l65dzs4jhyyNSEsYoi2rzuVSsHpTG5knhcruN2xrogjl0dXeZvwmWkk
kcQ/qkc3Vji9q6tEtEST0SS40PkietHvUK+SjnnnReompODrgHwDxs50qEKNyDJO
1BRtp3h3xLMiy54iROPX3OdBqAcaULDc8aVcP2w2jnnbQGyIe4e3kIhYvp7m8/P/
Yv6rjTvm0/vlyn5KsFosX7kEKFsF85Rv4w/faz9wFzSWQUirwoOnIIHVayakQc3f
G8YQn6vA8OLI2CHobZpdzXP7X9QGEmBFsUsBNgFBrOAUx7Q5J+QacBXOjL7df9eL
bY72oq+gMbY6S7J1q8EaNvcQsXt6QsnMSDUnNCCfwNWFjH0nS3AgNMIPigbEabO2
I7gS8/Mko06rKd6qJNRklOi7OPJenSnJoAXuHJT3+5mK/py8jrn0pOR/rHtvYIGa
/QO2hUABYEnCIW8UMp0fcxvT0wXhG3oUAVsoKl9CjTCFrQYE8h6Udp2/UpTAJowF
sB7t024vuba04/bzOdU3UXEha/I0fJtm6Z8Ad7tkZcHceA7vD8QQsjbjdoaGbIWd
WMYAECqMZJHAukNqG7jiqTxiFrI6rmNOXc5tb6NM9iUmEpCUJ1cMX7bGq9J97LO2
g6csURGjh25y0IF5DxRMseQG7jWgKH6SC4ZCVlRPs6REwykiS2exR3EvcoWuFZZQ
arfSaF9KrQb0DLsqmWkYzLjz8iIAPMRaKhQ7RzzjMVSnyx7u8pxwn+3GGxhsxKj5
egS0cABJsl21NjcJGfHJK1qlfoNWit0AcF9vXwOzeosVwbOp284ipTszTWwHlxMu
JzIpjixR4XHauI1eZX4D7MNf+Rln9+lYxM4Yo0VYDkVaobktwf35ii7mCGNNcsRq
spOnqLNP7ccG+qWrvytrtio/JARZzqQpErj0uSLnc2h/7Ys7UZDOzrludisUbuv1
4MPHdrHUpajtjYcwVOhLRPmTxHJieGCBHZCZZ+LJuB59HxPvGnjsw9e8fIndW78S
ENSo3dN1YkFucGj4imYWsfGRVqL/psuFW83Jsx8F8bE9hK2EvqMsL9jxMQz4xdgW
pxSOfP9ivlDbtN1874mSY1kf1u7QIoEZ9twpNH7dpaMrYqo/blLD2u2utkCZjwfS
Vjcl70Zr0HdEAXsOfwZIxEN5WznVT439E8LzcseAJDelzreV4bogKWYiCHsR6bca
YQrf+2rqiJA7D8lukQjldvStfC5NG61MJrg9mzqtldV4aOKuxVA2cEbYY++g2yki
jYXUsfStf5sRmvSGaauqBJLgcBO4v55fpL5tX4N+EI+dGTevgrv7zN/FpJvsdZ2K
FvqQM0yeHZRVJDEVj6GEhC0xu0b39edyJ6EO8ru86DvkiIvc4HwCWbI/QjSag834
7mAaSZguHduVgGi3igaZ90b1o9TbWA5Zzqn42Le5pj3e44OBnsOcSX3vbpYCztQq
KUiwDcOrZoWQVEEg4j6Pp/gUlZDsitqqNO8jdngQGiVcp+voVpy/VFCIvY+QEy/m
PLhSvX2cuzPgBtv8CynKaQN1lk67i5QN8lFiaMUtxf1ZdxTJBwotteXuAAHduEhd
tZpwMUfvxwFgI9IgKAKgV8fDq2u4AHCA3Php/DlS2KCVNtu5Rl6mCq1VYPAx8XNE
tZVsaJeZOUuShWQY7YctoiiLN4n71E0v5h0G1lafnaAcE2wz75Qe73r43f9GwMiZ
tNkWgq/Ddofyf3y4VhAfPMw+0Gqvo+xoK1tLGpntMzCwn739VlvSD+jt1G3E//HN
g4TxrnjfE2GQ6vYkfuU1ZA3HbiibQRJFwe3i0RMRCjmkWliPOLLf3xv0lkczPpyJ
7QarCKsXtsdRYUDOa4FLfChntLLZN0KoAeSrrKCRubm34pNrdjQ8nuEwO4B+zI8h
4vCjZ1zakP/HjzGStMjobFA8HAXCDPNmO2d2/QqHYvaRvKXGYaNclSXFwHDQVf8r
Xz1hn4om6Mp2ZleVDicXTWUvCbA41f7AfgV+/u54djMJ1JLE20vxod977ZfaBtjF
LeV4H86aDHJGnNPw13ikk4FgDRg8OfshfNucW+AluKbL1Ysm0qJh+G2iPEIRywCC
lUgh92zWlMs8yzKXtNvRAEIkcWuCz6j/+9uMelL/lcPOMNqJgjl1PCP6ahAPM5Um
QPcLvG8qIPUdQCJsgeuC/HKrAazTWs9Luv6AcXDRuNHvdLBuo8alVwdsPCMFUks6
dNrF2yEelkRGL9oQ9JaHPBWuoqH2qFiMYmwLsVl78WHucG98iWN7UgPlFb4rfF8f
FieD9kpN5uwUfU2Kx7WaKbXn/j3s/YHIkB2NVWlJgnvZoX0vlGpwzXyUmaM8ZdFD
qN3muxpyP1UHUGcNTCWRSJsem6ugRLMbf/rcbEEbyjEd6xwPAvM0OJ06qFqjfAYf
tl7cDg5HPL16xd46aW1a8jDsDF4nuWlX3Px7AXrrqZDsbKYJeyJupbzvR5E5QbQ7
9cDaY03Wrjt1P23w0PFeP81oW9k1bpxMwTVJoBNfVUlJhqlDc8ya3XUzmkPUr5nO
uUobzQAksZJwnj52XHMm5RVyjGG2jo/VhNXfjq2RpqE7oXc1Fa1Sx49jsrsGgSS0
5Qyd1fBXAVFd5FgB4HVsXsW5kIMSDTor1Kxi5YDW0tGKr9niAIAh88zodnoCPOmN
EnzqwnTOnO8oLZeoClo37JLQuRcrhkGmLiYrd5Uik+kRiT5BA50Glh3PMMMScBot
2EUIueCyX/ygEK/A7fPj2aunz9va6fiEoxMw31DZbovW83fIIAcqYqxOnHUjKCy2
JkA1nCNqQ1ePteX2taOzHDxHWEgX82mJcT8zYeOG5dQkMaSDXRJEYfw6nQaI5WKX
nOlIox9NL/OF8LBrHx84BZZMzm6DKEhzU23gNjaimpLjwophraZcR00yEgflXV3r
4SPewHAC8LJ/btCLjb3t698zxA5tCc3/AWg97hfcoPR/Eybf5DP1BioMbMwvf5j8
Gj/0IjIoxGFIkTnoCtKJu0rbYNMVEr4WYktT7XjBDtWuxKdI6sOAr7u3fwVrIeZy
pV7IrLV6gpBSI2kZqcrDy+WZJzSlE6LCGtQNN3yc9sMU874El+z+tlRy8I43Gvzn
lLbaXSGyxgQO0ILNa5yDVoPQCxeA+c8shqH7j99NFaGcaKTGn1f9QN9IdWHjmmR5
wy4ixNjhlgAXMuqjeUSUdffQ4rzVV94IDJChO4zZgUhxxGn9PdvlvfKneYsNVdoR
8ZZZ9HKZ6azB11ZpMbPEj+bXSgALJb9auwzqxP7McZf541UM2bZ3ASNbw6Q43kga
rYN3rm3jFAWiQeHa1NEeNpEGfn1tU1o7HSjmRensXJLiS6cWUzL3xAeV0ktTn3Kf
RdFDHrMvWxD/QoRCV7Olu72lPn378n5GI114f5H77a9Ik125QvOzLAsbfptibJMI
zshCRG4lASBLrK/7sB4JN7Ov7GDDR0k9zflraJNctSeL1qg/Skk4QKWEMLHN3ne3
R8wsUOPeN742Vn7kEGoASvEZ0PMAqlh/TikZ4tuofylnF2AptS9Sg5ceTZHsrsc/
uEsT/tLYAMQU31FirlolMh+m+op8hnqtiuhHwqKSlztIsCFj+8riEYa07Dqfrc5d
mb/WHS9ymG0fOw6h/Xkm1jFb/MLnbnrfrp5yP4FW19vrl5ao6mTaHYqJUrYrz5TN
98OT74jiytmvUr0ckpXEKcvSjNOlQlN+717b0n6TjQMmOJsqemLjmobJDjccT0B1
xZrnY2eaZByVmhMTm8aLhlr8p6ynX67W4ZfPg/D6Q6Tkk9U/awSmXKNmcMgECkFK
8/AuRdVPpNzj/GwXfw+reY9FPTxGJcCHODgWAM3DzKBECC/9HUf3A2l5KXtjZ+vB
qud8DzOKNarzjNxyPyFRu1lW0ymAAa62ob847p26nN945L7ekpkD2BXkWanjvq7N
XKg1+hkb1+JoQCblktFwqp4UUZE+3E31K3fWe6NpjhOu+BPHTUynq/VXBe9Ci7T2
MpfJZUytpOmm/2M5Y9uW/1PcMSBI2c8MHecEd361eMoVeDhYaeGYZjzcXLceidsl
JNrpcgakJUwkyS2lRLaEJLJ4AwyID+kjTegc92WpkMMsdQ2K0b/Y0CV4hQSZuI6G
NqH5U0VJ/Cl3jwVBDEAjN6S8Gx7EE4mGEVcuHSD12kqBq28ktLeseFhZGHadkN+F
ysQCosMsG1JLLIzX/o8ZVSrN+Q912aGbCg7nib2+dURt+p44WBjvqO16cx3kq1tQ
1YgDHlY6G2hV0IdDUsE4RNQDEBDOZo9Q+GcEo9GMs+JtJjbGZzAAW5oVwsWaDyYn
4rP1/1wE3N237Vdp7e/8qRRLz+Kp+V7Rs3hB8DUhczQUNgDuM+h79htRHyl/f9S9
qYAgvbx2nNAMvryLK5lH3m87PCHIkHs37WLfzLJCapeWAEJN28i+HdERBM4W/qkU
oc77FDdH8WA0VjzxbAvYewfKZmrBttHDbZdWI3VL+E0+vi00ad1vAQi13g4JfpNy
cN3keZWP2zNR/1RPAP9XViZJ8DeoUcUPJEh2XXTEASkVNKXKmzE9Z4PpuECWgIpP
trTiqWqzOibIn99PqgkXGcBW2/eXi7romEmgTd+7TpmZTPnMoHtU129KKCsr+JwT
3q/y5grnDEMCHl4W0tGWmGFFKK0Ew11C/u5fChLVWn4E2ZJ0yKrejkwH9aTOXJfs
qFGj4o92rM6qrAKjKSBCbHazpcRa50nLxCELfBsVVm5WKEfoKL197VeQ66Pp62iS
Dc8pX1a7p/HR5mwBRoa37M7322HNSg1i/hUbUrlP6aXyPgBlhbmeIb+0Msqc2tti
X1q17XdhzF5a7Y1DAP9kf4qODaPP8tcpXO+75wtBP7SgzHo8GYP6boL/o4V6wURz
iZciK7fyB04TxIA9gaaaZqXKZdG20gPLUZJuiy0WUyP39AhN4OUIwVzRxV7BlWO5
qxpQ435q9AtNBOhpu4c1do6ZDolcmxUZmhdJ1//X9HFnTS30Yt/Sc9K45+o/yess
wy4Wm+5UXEVl2Q5kgd6s2g5I5zrxMIN2Qe3Mqq1aCtgG6KH7LCp74/FQFANAnnhp
x6WJe58Fc9eC4FkEduhajIEpMNHQ4Yt7VO9kZWfFIP9BmFWWM17VcFcYTnvWC0sV
rzAP2P4ILQTGRnvnmzvI5V+E3XUASzOHFCXXVkDmghC6ZEA6r165Z1fdMdRg6H1p
PXwFFbpeVzDFL4LuJWIx0nLd/ISzJO9jvtuuvl6231ufTL584xxuKNGTzX16HZ7M
SCut2o4L+zVy5Prte+PxjNZfK9Im8YARRKf/ibxqLd3dNnqa9NePRVsJHUOjrS9N
6Yv19JttiW1UBJ7SNnLqYfaqAIrHKetP4ovY3OWysRRYxuLYhof9cVIo6G91s0dV
cSt4PkLziZlV+HEl31VxcdvBAKLlAJfDO+UoL91UNwI7RFsbX1txmoQE6GS1k9ze
5dmt7FFo5GpMAu1I2seACp5MasGD3jWnVKAN0I/fNo/pGS6h8jGpzxVVeinYoeZJ
B0IQUw4Cx3dbrxK72hBtF+DaYWOPsSYZBMXyK9rUypSV9gJvh/x7TKCv+vFUmrHM
Ikfq9lymMjIvCYE8OMt4Edv5gvrB6FKBx/H360jv/ToyPulxtB6SwcyNVl9rLK62
bMiU5iApp160qcPzMZnSwJs5+rchxgWRG760alg6a8klkFQlbyKXdtRn99RWEDSK
ii9qcjy4GyXiKXQ07vhC6rWqqMeB23fNQUIK6HfwX3pFM7EWx/5qwKbWtEJFkgsU
fzPI370bSsLZFA6QguCy728ZkrVCL9j22KSkPQFIMld6ZjpKiBEF7PKXZNG3u1kR
jv9KBB5JiDLvQFoVvGtgSsiQrCkKUMIfgj5nAq+2OnkCGAAeWzX8WZd+4j+d16X2
MdEegNVcPMkhJM9O7sBjBuEMQm/bPzzKLL6HT99mgrhQkS8kaJt8Gql17zyYtphE
gm5TvESE68LIx/P8w2E3Ya/l/wrDzGNh6/hnC/hdlCC/3cw0RfjyPUIGiTNMLcch
noCKsadPLoPmsKyTvMT3uXTr8p9m74w8eK+lhhpklb4+2mJxfbhDDOznVrLBNbEa
lpHLkd/cc0GBtVIoHR8jzqKs0b0PQ+HOPE5J+tyEMQUCTM9T1Gu3IWw3H/AxLgK6
2AX6zg8dM1i8mXu8LepH+FXwO+laaJNu/QQeMP9u4VwxKFWsUehdJbpNRKxp4ers
flyaXC5cRpU5JCSoAa2ZK7Rzv++VMwbWafDlmvyw0Srs6w66H2Ije+XwidYY/N6t
MiwTePK3doEiM3jCUTtijs5a10GZr8FVrKJosh97okKuf8JUJlnUvMRmpvHIt4hk
/8mIPWN493vxm4nwSiz5YAgmRf0EZGDGTsTIOp61E2NlSGdToL92h0bwAY+ubJbP
SK6L+5/ZqwfTUYopaJpXd1uQSOWxDmiwlxEa0sL/vroV0Yyu1RdQPa1GkPWQWk5b
OGyNaMbGPgNUASLtlQNz7WyVcUkWMgjLo/TYZnGwh9qMRaWV+m167FeQ6X9WEz5C
lqxmyBAeFpN3LwbbAcC7cpUwqto+rFCrtS2nQ9lsCk9q0NnNxGqROa1A9limamuq
Lm9wIzonbTTtTkhDv1F46+px3gDr8niAem+fHVFKFqk1mi7yaLIcKkPRSyNEr8a1
1N5NEvNbf2AuZt+453SeBb00zW2za/w8rHAqHY3/oh+/gnL1DriCtJekvuTyxG7+
Az2CdK8lLspE7d4pL7tADDHXGaVflx99Ti9O/fmHKDuxyq+INjEQCDjekgLedR6x
QSAXWNUeRXDALdmBMUP1kVGZCPkMEq6cg/lGNSOnZ3htdDdnDvtzv5TH/nljIQOy
71naPwXBBgV7PIzJv0cUcw08KEVovurOQlfryEaAIqSinasduvAWe38A0SjYlKXa
0Jz30NnWQVt2LJnKPFKGXFI7uVcKaBvsgb89zqcrf4knkChUktLYPavccaGGgZRL
meZ2xr3HLtLlr2eEf7TRC4MdHZ0dta5c+hTsep04PL/u3Yz2KcKgsvfDtGN/7v2O
mvVKA6QiMnOt/cFKwVC1HnzNuz3XrpBDXcKq/akm5xj6nbH2w+RkmhIF0ofzASWt
QFaMm++IJJUhfd4+1mQiNtTM6F/B2BU1jE7qb2PgXcqEegydGnbdauk61G3cuxkH
ykf2mABmtkBdJ7iikvo2oAEYSGkfAiOBwVpnDD6XM9auIBQljlWsl1eCPy/pt6ZF
s7i6+Rmnoc3pTRPUnFi0j2nBnq4GB2+u3yiESU51jD9jopmV1gHi8BHqP3U030Fx
sQY6odjX3nExsph4Ucb4ZB/0TdBgg852hKTeFQWLs1qDXH/2/fT6HnqJy0RDNJLH
18tedK/7AD+oEaUtO93+Ffjdm/MdC/4mYCi2kz+rQPMff8S0I5tg61ih93IWH6p6
j5tOIifnAfR/hK4HstlCz3P3THQLqmopVUKpbfWrvvDEtRWH5yGGlOxtbjqZ7pHY
gBGAQp1xNIf0yzfiIYN/Vb0s1nLdTpeHAaROpl2Pz6HGSXhXqrqjYGUHYKo1u8eS
I949Wal0Vex5HThbFFw9+Sz0OIap2wyGFo6pFSrtEHRg366Hkdzp/bxRSCaF4+Nb
9FjHB6aF4Gdu5BYlT4rbBw==
`protect END_PROTECTED
