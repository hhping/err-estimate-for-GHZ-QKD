`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
McBa7VmdXB6qsbrkx6nUALBsDVRpbYipMChHL/LwHFg2Yy87f+n6KLW88iFUN375
nq/OJV7vzTLj5DX+Whp/ejsW7DiR4PNuDoF83cbJFoX3uMzyy/7MbHVky/rxisay
Qb0tydOisPJxCNx+oQA7gog3+fUjYK5X5t6tHFakoGJqjHrCIppvnFKuByyVOVji
LXDPwDczxeu+4UfeoNF1dMZV8vtaEdtjRlRrdxf8gLacwkNu+PP7KFMz1HzDV9+D
cHcyFPDTeB8lhAk4NjevsanbWWaB1/B+ibjHdZWA/7jBskMOLAey5FoG4KH/Pzxu
N5SccGZyp2AOQ0zMjxjhvuIiig0pHDqLjtVNYzpaZOpELevSH05yZzhMiLbGZIrO
OOBeDFaF6gTS0gbDy+U0DAKtPYm70JZORphJdX/GA7Nq7ZpZ/WsVi0CsMwC6GS0B
weEYLo4iYL9mrBnhZHCsK6pfDbskq/DPe6ctNsQLR/X1zGW0h2ahOhm7RSFtSR/W
jNNv6rXIXXIAZEhTTLzSf9PAzkNCK1+/1z0QkYC8vDApUIuJ04LsAUmmn9ODWR8D
C0AuppRBQdMR2/t5KJCCrGcRSYnBMc/wEPHRi6fb3PxHDER8XVhQLEOkCqi6kUXi
X4cveiJ9aT691T7Hbhq7IKbpmDsooog4/0akunX7EX33zNRjQs8v0E+RGpC82lyi
fMKpTykVrqshj8VYLnBs0h0ANWnnO42YKSsIJn4OgWvQYyWW4yKpignr4uLFnY5D
wduvzpLGw+q4S3KVgy3ln9Z+42giJUgG/Ki8b0epz8MWc9PZle0vS6y2RCqc1wOW
/hxABNSwiT2JmVwQmDE2l56osPx60y2HbUS1W8Cu02LhXohRPYc1HoE8foyYmlTi
IEfJQ65QAUuQKiFImLcTlXFIRPZLJdLJItCoVbXu+PF3DwcZcr4FlgLwNzscKjrk
A/XUzSBY8F4OHzZKzp7cj4+ayl2VobpkZZZmUjx2BDj3tWpQiQTHyr2Vl2/Oudwc
dsHVmAzHY3A7O/OeBGzFAQJF0MXy+WMmb8SeL4c6Am+MOZlB147s6W4/9yIFzo84
cSr/o69zcsUyNfVl0hDVu0BPGOzdrHmOzlMu8I/d0cjd8k0bTmhrqJ4qDQ2JEdXS
ZrjDM1HRTcxLK1+IirjhG54X8vO7jA2jLay/LF3lQfruw69VEP/x/1m7+iP6EQ2v
i8KmjkPEGoULruDlxXif96KAaJTDuYo+1PPjBv4A7fHEJZUc8OPc0+YAftXcEaan
vXeMdduBOiuETQO4dZ5NiZgZ/8xvrYsX8Sw6J0eU2u5F4ESUkuAPsgr4LS/sCHqt
onGSNFgt7I5/0xxSCsA2sdwelYjiiHQrx5b6uV07/BnIARmdSveyr8eY23UnVZ61
yGsJ9QDufPXTOXBnoZKI03Wc1XWnTFuNYG02vDvkJhKbOZ6K5d27GmiD+JE1aNhV
kptFewRlZlRgS2L9fjlXu1v6O3UMb0GEAdMNGDb3NThsTSHCkEb20DJoopdLS36X
wobm/66NN6PpTQIhMmX4Mo+qO+9uvDY62OkR+qPMLTqZUSBQJydYSeNvT2GR3EFQ
5g/6Cfo4CL0/DEC8qTlhrffg/CLcVTdJEMIq78IXVoadAwN9FXWPQMOHK+fGsbVk
mRgQ53NEbFN4RQ/yGIHbosOf5ReJ848dj884ulYsC0qW1cqGmKuELYIw3dKNvUJ1
XjQLojN0uKD3HXgff1Lz6vYAYunWpudBehp94k6TUbt9QBv1yHZAM5M4FQYAOnCB
eydb/hU/wgEhee2AprDVbcspbnRf57TBEnxR/R8Ztyimk4aGxwxHT0q2FOFa/6uS
ePWoKPo2JjqvR/X2kFh46/0t6L6ZqtebfIHjDl4i4qQF7Ij2zu5ppSX4stq/N+s2
yGYr836FIxcT5a/LYuM8vAalRDVa60onbjzd/FtgsdQOlLDXpwaVoo05803R1GFL
23MFtTs9THEH8PseRP79vEKyy3hoNa8SbDBM/uYi8ZWuvu41GgEfnGbavHoKW0Ej
rAy7gbc61BjBIH7S5KT0OLmWMUFzII3S8lu6phrUPu6JLUbTsQyKrkiFIW4MrCd/
bAvVK+0Dnx9duEhQf5ZOFabAANKIEyN1MYc0hp0eFtC3hs8NAs+Vvl69N9NI06e/
NwWny0Ejnco+NtJaGb2AxazWMRym0/+Dd8I3LJjobxisrEotgBbY64gORZl+iZ3f
+DfC/aaisrEDyS6xt+fd69jpfAqjBdEy7HU1hAtEOvysfnIik0yQjW+aqxMQfFlt
hJKRHnpWvMTevwecaAYIwGaTv0RU6N6kNM7KP4Lw/RwyPLwL+mir5jvERnBY+jB1
fneQoDyCsIx3rS+OKfpEvGADswjmgkVz/I2WnBxhlmAFP7u3ASpuT7DsWJ5KDTyj
NblDTGCv5V3m3eweMF6FKcDIKEs8Gyo1S+rzhm8VplTNqFdlk3wveMpSPcfv0HJN
Pc0t9zLzPUMkkMuvq6RILZbd06EXfXT5SHVpAph8t/8TAQOoqU/mJZyohqFdURpv
8bHMc5GmsulsO8PiBv/+ehPX7qYgGk3oE4StvNo7WJ7VhzjS6qfJKypKeiPjKMzr
lgPiFqdelWx47CMPC4S3nBPLVCYYFa8/VaIGmiYIXEgRT2LbNZCEkNNB3lerpj8u
d/k7oFCwReNk0tI7bvNJCVi4FO+DabqZAAHaDeX86cR6KzvT4EjVzpswPKGJ5KB2
G3g/RnN/PmvzaWovJAZ8E8MJf2Ti8BT/753Ay7rADZqMzKLB51rQ8avCvowALRei
3a4cmJGqmHDu0B0afckY/15QcmIAQkTIA9obsnWujslrtSYGh6nPCxt9SY1G6Ddy
OZQDH8HjMxTWIg7PO5NEjabzK4lQBVPxFOypMkkW8gOsqktRUo6GDgR2Pw14EgWn
08K3AggM2TXrzO1pAaOujG+79oXz7YGCmCfykUTUknWlft/WNoxbGbfNMb3miG/o
noOda/06P/2SrQhH5fdrjrVQOdiIDDcwxFQcxYt40euCNaYya6lrlKJEIK+OsJrn
hChC+mXVaKZrQrH/lmXyoIO0cJIX3SPvUQiq6w04Awi8z61mA1Mu7mNfN6ymINkW
q0EAGcAzH3RSc5qq/c22seSJXeVmsrbuac1FWvUdBbuYaOKkyRFUwZw0ZBQDlhSe
YeYLiCyyUCFApLUZ/IeeBbvRdN3uaw50CFqipYmFBPqZZ2Q+km56+90MC5HX1A6z
I35OCpRssfWn24dNDpoOFL1HfibOjtM4KUhl+I4N2pZEJnBR7qEDHtRz88G0MGoj
WS9AnRLoWJixIktkKEvyH2M94zJKK870zLFlewF655Nj7eHcag1qy7LU8LT1bYu2
JN0/CquwnhmnIE2WkDnJDrioEmvkhSttdOg9euiVXOaMjx4HP+tUzRhd5kcsSAfx
JXilVD6284nfEzhxo8ZK/yAvr6nXUeDnx4oD+IIPwbS8vrOW1n7YJD9hMjG323gs
lWycqTlHLXG3SbSgkMbcWthG23eWPioJJIdZkzb8B7wIw6UaZ1WE9gshdtJB74IB
GkSP/lxnRsnWPsuqQDmpSimvoHswpE5TLnp0vcrnjoHJQsM+J8QA7bspWTNsVrm3
D9lyAv6pCk56QI03nfMuj/CN73Lj4sYtGow/OC/O/hflTKFkarnj0HQnfxttNYwj
rFbfPEw5tF4uIYIuKMlwpSCMwAbatH3maOiDG9F3Enx+JNWuMPp34UK91f78DZ7E
dQrQJxukRUA7JcxfzKxIKeEZEDR66+flsGMftGJrtr9f0AmeOd3xojEgb+S3lqSH
gLIP2SqOFGR+VIUttk0dMwtpJfRgCGIwnanjL47wrkhB5YNsfErTY0jdyPwimJHb
DR8alhWkSnkVFr+V1rZgNyPR5eKLWt6aXMADtVWEYuG2QjWJKsuJNpQ1GY8wMh9K
lIulNLY+sHtmqzNjz+O17FR607vVC1r0T/H+fzunH1SrwsIcGqU3jScE6sQ9NH19
rJmm3drFJX3AsGFP2wYMlk3tTDZZdPVZOI1LHRbwDptzmo0ayn8OGtxPsdUvqmNj
dPNmnAx/KFZP+670dFABbco4pHVpDh8mkaCfZsDxkY/TxhxuSO9wDCWGWwLXFWQS
fH8C1EvILR3KZCnNLNBc646FXx4zpZ9rCkjJn5qw3fjy2tJbl8bZev5wunGocab9
HxjD3cRZcCTVV4q2tUmRGQ==
`protect END_PROTECTED
