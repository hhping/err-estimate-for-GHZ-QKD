`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wK02Up6LTvM3hW+UsS9FzPihtnVsVCPPMpnCCiig4TF6wOXfG12ibl//dJ6VoeB2
3WqKQ8zkyAS5wbQZhFYgkxycFtVMLOWH1aNuI3ciPbWq4hHGmHS+aNwkjDathtmS
wAFuvvzOAxEesp7Gv237gQ5YqoqlDCpcs1ljc6AKym/6WcrJGlWbQPXdx4xIHDuH
xy9jfC8Rr18DPqpJ4ToGffOBBFRiEyWGvWWWW3fRfk4pJkGvPb8vAvH1Ur32i1xq
wfReg3nqiECldXcnHI6ebyGE/CVDPGURY702WgXJqb+opg6btKBbqI4zgNb9s8BX
yYrvAx5F8wzXKmAaEfv6EYqEThIFdFvcv2aJYnIYXyjpWmh/V6QBQZJUbjS/babN
u2GKLUEIe9nQ7Ne5YTDbPxYjH60YOQyl389rl4dsEQpqUqEUgiAk0oUaXpFAdMc6
HbXoSxsApq0XVTznCVLejSj8vv3+33e9kLixeIGBlQcG/fIi1Q7RIm+vh41iDx+i
0A7XQ8eGcDrOdq214zOZaskNpYpfGajBOocSZxp2RykyuFzHn+dnGp7N+IA2OrEC
fD+gZQcPHBrY8gVfPEqDkTvG0XJ6FzwmOi7oyUND6xlcUgxDyU+2ymA2nqAW37Xh
1amVUxyW8n3gX7cmMMqJ/J2D9TU8bKJMX+nIuFsIcwT5/3U8zximx7E5fdhYJmLK
UywMXuSVAPp5GUK83/GvbnXUq+IEHjVG0h6One3IV9FVwabcbYjBjA+S25m5vKZZ
w5lq+rYP/pUrGrPaWd98WhcJMfZCA/qUJofJ9Dkmeob2WIXb2LZpK/04rIruQTSK
qtBJdcG7qDKeeX+rMPXet7SFK6fUNTdvsnrhQLIa8CymDN23V33PxKM/C41U2CS7
pklY5FrS61y2liqZDrTYoN+Ued2jsUD1grx5emCK83lc8ug0dyTD7cQQtVSY6io4
mGvB2nj3l/DEqsmddWCG4HbNJFMHndNoeoOEmyZE6NKgi0SD4I7RH5DrQ8ZJSROF
don0df2BpDCCQ5AS/uBT4bw1+JVWXTA9/+QB7R5RwCRaXHIwWeN7lBfTB5cadSup
UxACK0G4zcawN1xfUguCbLgafa58ba3sUAlg/I+If4FaFunsc718eg4fqis7NDDb
mxy7f+rYFUna+aT4jv/2J+Il+vfoAb9wabezuLq0ID7S5LtZGb5sBExpQttxuVId
PAjrkUMWobCC+cUwA38i2sUtmGmU09BRoqvystJbZNMx/cJwny3K619niQvfetzi
KfqytN5a3I96tVimAtN5wOdsLdCSXjJNXGx+1Y4cZAB3AYb+5kMGvz0CzUgIn6VE
C0vrI0v5KEkM6AX5njo4ZDFZ1qiR3agEApyGHU8qgPlhJoiXLI5bLDAoYAFzyI52
W+X4a3c4wF0BoO9qFFZpsNpG8k04QhexZfW4gpwO5acnGZeOazzsjJR0OozAWWVZ
q9Wr6njo836DxGEDjBP5f/RoE8fTzzE0Ls5CNKmofitk46vgFS1z9R75XJyPwq1n
iu3v+S1Ql8/LiIk29lJS5qyU4XYsZjYKP+cGHx/qQhbfVxezC8D5tmH2jNcmDEND
arM1F3Zx1ARaXYCqvt5wo5ZvN7mmbWm9nR8F2oSDZysvyDJA8IF9NZk/WM2QQDF1
94qUF34WqXcK6BujS4ARgKyYO+lk0w4/7s6DYbvAzYA+ViFzv29b4i1sXggvxsq2
lAKCyEwyxWHEbXglFan4RpFk3iK8jwgnX2vIuUsW03BvESNVac/mPGJJrVXUu7c6
B34kdPIJ2cWHt3/W2HdPLLhpfcW7qQL+sJrG/vCMmQGz2rfYh4T1WOBdCA4UCTeT
GJejat9OSppcFfFpbnNfqNEgsIbjzdsnoMa/e1j2+7mePIXr+yVuZ/HlpH2YOpAx
xxCU06fOm9sOCN+Z4ypYKr3Dab/dAbF9+MjRC3lK8CUDHKMqN915dU0EgvBK3tv5
2mVzTkwlZRraTT2GU5Wt5wJi3kPL6sPEEQqAVdmXmcCF88LMeQxaVbXVTQj1o1U+
2DdRIKhH4xDtjC9bBgJUvFMCxSn+40SzsBVkhywxjiEHQlSPLd5Y92vj7cUtoZol
rAtjIukG+R+uvCCg30iKIVB499V2Ne7trkQIKB2iGsT0/p/KGJAQjf5valUyzKgj
lX97A7VhiXh51WA5UDFf3j89UycwQnUsjzCpIv1h2Yoy6M8UZitTjWmdTcrtJuBa
B2wJzQHSJ49wC4c/W+epuEl1j/HYP7R0/k79QJvJz2hsAbW2p3iYAiqmRoCGC0zl
5wAyLIQps7q+5d4lWfy+FVY3YFJxUkBQjtd5I6OSnWV/MjiUuJvF4N6kHa3MsE7j
CfPcTjHOBcdAiiov5WrMq5rYbVuxGi/Wk9M8XGBzgk67Bo7lgHzf9jtBrk4+24+o
4SFATS1H0Qw9z61Gci7a1o9pLQD/rDR88FOBggKMT8GXC4lYh72ukagU6FUu6P03
DjJr/6aflceAHxVKtKEtzxdLVItG9rzYDa8M+jOsX+P1Tv8AM+ukTBVF6Yc60EQi
wRR3KP4VxFwWDrENlalmNTB543ercq5BWfrOEWeuwTP+35oFLYkEuTtNj5qkky4o
tkaZBD/vzngdPObk39NGSto+RS6UKO5gPsEOKQ1EHTusFs8Y/SUQ83q3vlEB/8Kv
Kdj/sQLDDB+6iYVudiLmxATuXtDb+oJnb14YPFXjb4YVhuwme8f9SjdVyUvL7UvP
MkRj+IVF0I1HpGzbPV67t4XuuVd77EW/yp8J1r5MdjYiqRAgN0WbbxufA3ZfmKAQ
1imREgxzbl0J3HL4rWwyK7q934DetA888OuB8IBE10YGSS6pqgtcTaXSO/hQNrFJ
vmnpXRoBbZvldfNdljFYuLxSakxZbVWDmXEFuE4BUK6aRJaLZq+eptqWeRDMJ+iR
y/9jaqijXC3G+CDEqG/w0rJpnImw7UF9LEb1Ihn+TUx46f2/3XB3l0doJu/FDZBB
zQbPhxr6TCR/p912RiL1toUPbPeAWK5kLxdQV4+nj3JleWtsiEOTSoVdfbsSLvUP
3unqBIRv47BhfY79guNTSO7gv3i5HTASREQV6KsLpOZkCZsGUACw5vZJ/OW+JB1t
iuOrGurHPbuZTXdyxLi7xWTcB2UMULkL/UMOCcwVHdlbrqsHtWlE7uHuwfzOp+ew
CPoVbrj29dwYP7k3KtAVwvGy8Xvhf91p5i+7MQdLdz7tiRoharUeWhCxxGssaSG0
d87ZeKbqMRRGm3LIeUlprXHElAgDtHC8r2HBuV40btko0LirGr1sc2nLuhEk1EgJ
Fv/kGdLDMQkDfBLMPbvWQ+oNQkliV/RpauiMq36Jg6cEb+0cLMGdkEh+7+PB2DrV
vA+SLTVyqxxiAP2VyvNbU28AQP7//ElyDQ7/IaL1Wv/oATLz93OdEkLbMDoyFPNm
2kMzZCNtRUh5T8F1ti3N+/+zW6AuRz7aHmF5fJsqd2V1yHGBQH2KclLk8rwosYC9
eNqKEMaP84ONVTzMNdymJYgXEJPEx438akYTptIXanjTNDWfl6khogvsMwMpivWz
kuFFChEdKa1Qqx93aKTH9pyP6PT04248Mof9SuNThmiUe2LJOOi7qYoI4jenOpqz
lMgp2NZh4qgrw8p79sXbAmbXL1OfGAgLVQlixrtTtryGgSePxWMwRhSrbrvqRc5z
WECJr2+KwNBLRjC5jpROo7q0+Ubf7QIw38RjBsuDqtsHlLEqB1Im7B6K2jAZBHMA
Jp6XT4TbdXrijlXnlm0ZEKj0AMPDYv58xwkFCGD4r7IIGxMeHkZL7KspQ88FEj4H
nAHFLgnkv/kBwxkiOTN9za5+Cf9I3EnFtFRTeYSxfnLNWy2egyqz/wBGQC3SsO+P
88RORAr7YmF1+wKcVo5UQySh6Cmaa44GyPtNDYaxEgAgLGA8odwAJEDWcQMJrhSP
BVmqiBWI8ymB0rqGewtKpiE9rP4FLWf6AH6c7cxk7dQ2w7HlZfNAAPbUAHtCrbsk
ZKujGpQaujqM089Xexq3q8aDAcq/iMDuHAgq7ZSBr/MeRtzTM3wG0QM4CPF+mSXr
n+OmMi6Ce8r/owmyQDkO7Gl/iYSrNoxpX0qTmBzzCL8i3gMh37dhplHxK/CVYArS
k3FVUbFoppErdV2P2Qh5dhi4C+TFAEpiAC7GDiYKUt3A4Rv9n/Wn/yKOkweGZ061
kaU3OIuUlyAUD9yVNj7Yiz7wjs5ATWkolTnIzHQmE/3bGAZv8qWaMM0sqggDYZc4
mxarX6jhzt0WE4g+BwfEm0v+bXNGEM3h/KSCINtkod5xMrgS2N35Gin0FeZU/5l4
8Skatm5Xe26+FBo7AyTKgXbu5JrfPSQrzvL3nnz7cq/LDjc702iLO6ZzyvK9svRx
YRf7mHxzEnvCIOumYvyX6GxK4FpZhkAE9Uv/0f+dQGRHcUzUVo4oVVIiP+nx4HdG
eQ8Qwbipb1EajD8S9vhG4cic7ZCnUnlj5B7zwTc9eJcq5N7wWEeDLvPS+pcRLxk3
ColqEirNQAg4EkPLOooc0wTK8gRIAsFmKR4ya2MRxl5rLzc9yQ3WpvukSuN7Aneo
u4j1c/mjdCkVjchtv9Dl93IJMakrQ8SGLPzbUyjxDuraJKRz/mPjlY72ntpD+/0e
9o6LCowoQ3Hff8dAHxu8U1T0o5Kb4tYvsyMtmUHe8pdldEroYL30Tjuk4qfyxQpc
Xdz6Jc4IwtjTDr2bjyow9cBIXmsDOC2t7SdiTuoPmUya7YqFDQi/e0ZSRfh+ZYyi
hqStUX9/xE6EOfLVTBo41fOdiZXHeAhzu5Vqw7MT7BjY5B63zFFKB1MCH5lSKtJs
PxjPmgoUU64xzkzeh2UJ9eiTOPMxxLjy8OO3jpvQTw3gaVe2nsQVRAXcXkI4djwi
k8OF/gXZFUV1i6gKyII/eRqoCyflScXZcuhmyJ46mV2txI8r/3Ysn9n+0Ujltgt4
UgPg9hAyz/5kJ4rPaz9L7wmdDz5DgaAPlli9Ulv/qhlOuXNjnbnRHHVP5NZTdjvw
UM7Zb918tCIWvkX0RxaWWQhjDpAMecGhOpm6s3qRWK050F8HXXSaXEW5kbB7Xq0R
hFDAXb2G6yzhoJ+BDM3xMZse8SVz2M/van6luXh1HLVVjbxIJVuHI5SMRYsrXimL
8dStMAkRCBDLJRlBqgNZC2YAJaWCNMCN9zJy0yU2xug3QpQBBfquOJk4ubN9A93c
NBK5j62fJCo1zbYhoEExD36zOQZKFVELNW+afsmCJNvRJS+L4q/VXnAyuNKuOCwU
vVTju4V1SFFrwSy4eoHNcTOAqnW5Kncdt1ZXuYZg/yW7C7QGkRONqkfCyge9tQYo
pmUsRRcdfTx4ZEf+AGknBT8Jv0C+F5romNXjO1sai1miUHLRyX2WoeZ3sk1BThQN
10//4EpqHO+LAaNYSm7aNURjwHqJD4KXJkjApIh1OwZ6iztVOIg1OmxfsyS6k99D
/x1js6kdJQzrprNxJVyckqXY3p3XIagv+3+ovUsc29KDKsCautblksilVHXT9UKy
SvLqvzpyhW00TC473aPUKlxk4G4aZY0Suhhg75QI3zltCL1eH4dJ/JOEO1gEOMGD
4sJmTJaov6dq1qbfOKh8gHYZrOE8euF3dt5z82BesDX4MLfTEW2ojSJGYGXe2zur
cF1OjSAqmkSLHndiKGBQ8h1B1n0jqk9UWqi3pBefsUhKEnZleVyQ9Wutg3QbrqCZ
5JOBnsTW7ek/VcRMW0CXh7jyCG04dd+gB4OzwzDf/0jYZttM3vqqSiYNhsO/C8zs
ZP1AdVkxRjQXGKHfur/qdBA9FlfaAzln4JRFWuTD7k6LfBX+Ekr02I+lOkQsfZCR
D2UrnUxnEa+mzxhsTSMBnn5Gr69TmGqMLYDNDx4g8NnRYS4E9SPR7a3R80xJDEUQ
sgkV7WCMjcJeCg2SoIgr/67JmRRFgwPtz+mewB8eEPdeU5/J6gFgYgpb8ECSP6qZ
n4IAD3h7zG8fVtcob5XtRroZ44PR/rJy+KS4bp2aMk7EGEEEzGqB/y9/wfM+4cn9
ztbCRd3MUUR+uxNUXiq2JN+/c+kfE5CC0LuTJ38fX6eEuRDmFangjYtQ0gSTSYOZ
SkcsK/lw8QTsD4bknRlFDiR+yvPb95wpUzUFjzj4UmX/wnWoiaufzwZsGs4mlQjw
vq5BbWCudEsb2zgG0GTqm1G2CD0V1gTgZAH1VJruJTynjusTXjDAdaxSWPeelxph
DFBcBnunbAk9y1UMwR8lwWvVcwx4Fw0/Wd/ytA+DAbj/mbbawmUitZC+acJOtpRT
klPdzAfq9Jngk7tAh1U539diHDE+eWVM0Yz4Wj8r8VIoS0703MINphTv/GugGkna
He55FlSoHiq2ozbePPowvpFSX3oCeKgBFRPCntw0XykRUOwtg3s5MJAiQLdFyEj1
lkeIhJ2ao3AfpxKZrZJRe2m3YY07r47uuhpwCeHnBhxnDwDyiVWEgwXzMYATLnCf
sT8BqNqKky30l2dJi2D4HXfJJ0aQ3HLfndbQRucbxfa+jTY4ENxDeOYLbvvJ4J5f
eeML3BKeXeUgmxKtLhoe55vdpOJx7DBDUBetRt5C+Evl+v6vKo8A5X9nc8lwLPJ1
ZcSg0cEBv/q9W/KSHah6J6Vjxbw9ZxL4ZOgP85YfZw2TK8c6pYD1Nd5kcq+jKM7T
BLULz+sU+xfAA088pu0bgarxi7+wxPun0CuLa08sYQ7FoOwt0bk9iSNsv7P9Upis
Q4bw3DQpag+DvDPSRwieMtWuypt5yPCxcL5WXkiBpIwNGdZvV3OM59vu0/OQrYQ6
rFji7CiIxHvXoxR402hCfEa8w7wrvqivKbLCuOSYT4tb2xcZw1H8RYh4wRZWFmZS
2xJ22an1Wx6Kmu7qK9PHLFceJAkp5fHbJriMNVX5eywxfPpmr4tAWPH/JcSsjEs9
KyQyXvPMGc8Qskbcql4/lmay6Tfgn2ddJPadO12roicW6oaROXQTN74fZfRNUG9M
vK9OKufE+D3pDVOGXPspOhOtAmPdSJKhfkndCWwds6WeU/0PI4wZGNyo4Jwc3ANv
9+cD8WIgeTUNfnLpK3/aPXpufhJGvNhLCyaT9cx22Sk8orciwhJCA6bdKQDd4DUw
GNm1lK0Igr1Mqu8cKXGQ0sNPp+hYS3yYSuNVUaK7nYdYfjfN77xP9shjCY+ESbQL
VvlUSmfwt5iJGGkAx5x9m8bdJ5IvvYu+gTmODkjCJSjSRn8Bcila0iGeo/Kw5iXc
h+NRA5cF8/6eui6xo4NfpnsmQQCgmpxQwHbi8A3+vnu9wHW+vQTRa3fIj8Ij6V7k
gjgoRHtXBtk8BWwrJl9/WUirYtNwbdh1Wo9XhE8eKof2oM9fe6Oyy1PWlmgGG1Xe
j82KhStF5SDZSSOp2x3PUCsiEwZzNXYqnv2PDd4UyUJyeMyJJSSbNij6jQBCnJqp
ycXb0xFVwVyNWXiW0FK5eLAHOMWmaWzMFfa8zeZFwb28X74EvJL+tALq9v/iUxgB
I0lGS3AZ6Gd9wziZDYqIFucfBiNbDkmDEgb91rn2buG9tw+fmGMyQuaUBh7bKMua
SN2D7t+5tSqTdhmThdlzU1O9b4i3dAWbEopFOloCA6YiNPyqGYgiY3VFhPB7EfuW
LQ9xMZnisWm1DFTe9l4r8dR9sk6Y2no2UScxH8u8cxiEb/S7tqCC5X5MeawgdPCM
OAnEQs7AoLXrq4UBtCmp3LLwzUV6xfMQ2k5rSiEr5TnRDI2qqKI7XxSwNIsArnm9
WOv1C5OlEldrC+5+cLaVH5VwCuh7NpkfDUg4YWZ0KH46+DJVWNr+Uy6k4wGX1IVP
eoJBNrG3lcYMxIHtRErB7FUPg8/8XBejgyAnMiqLIbL0s1OnVdFZvbysoz8Nph/j
ao/9wwDm8mYp3RDYQj6siGCIwYwVEa2RZioK+3LQOg7heQYjsl2CLDC9CK0LUXnu
YdtY/yCNNOGufNtI4H26W6zBXcuqqV2d3i+2mAVPTgha0cMwI2+Cisp/j2g/NJEx
rUnxgZDr7PIY0chUtRgCh9tr1gp8uUt12RdHAMCa8uq9jM3cIxiZjzfJmOyk5DMk
RRBEnHT+oSILuota9bPraDsJEZdZWPbRrT82A8lNq5SQQy/wBxborTPkVKv0vdO8
kT21J/xRwnPTvoyvsdU4wrljbYR5tf/051uypWwyj40XdPFID5J+4UcRnYhGg9vX
8HDiQCyTpva517+Yws7M02SWpNR/gebz1p30fcsALBH406E5oMmWnox+RiW34Er0
/pAN1XhK5wPd4usaZ4O7jbrvTreV9si0jRj7YIcCMuzPh77VkqcHJiUNyosruzJD
XkKE0JuYz5I9PrqKHvpKlGnZrNzGOP4flEnqLYBVWTikDIRVh+AAM3z/O285PvWX
bUtUacDz8kl4xzhIbZdXGFTtnq157vzDoD9qtS7yVg4Ip+YgVrecANc+GxfkB12y
X3sGSnT1tLRp9kFX5M7xI8eVd/0t61QLwalUvItJuUU1Vc4Q0B4Azm81t2C/mdeP
58BfCLu7sru0B4uzCnIjcoVfdUS5qnuZgHAeiF9McT5ZeL2iNnczg4dreOW1/JeC
YvNwUU11iKjc4wwveTqs97Ymz5iHb79PvbTdVmVElKf4lm3CHp2Zy4hhPL3E93E/
3RTygkfikTNmQZcdo5g7QGfpBsRInj+6DVXJSEHQboRTS2s/guG+cjVSwwIBe5cS
BXoNgRyvQWrxhLfnBkUFuQZNI9EPrNcxRMwutXNja7pXYDLY33Cm1kmpxrg60oj4
9MSDeBL0aUhiirRg5BzBEPSow71E0vCOgBXQgUMBtzJdPEdBydF+qJuAsO0p9lIH
GCEWycPByHzCBpnLG5L4oUzcgpYfGF2XVk7/dKrDWXitOEzuOvQZDjWiWHOpK5Lj
Ra2fEOSao4FgwNsA0YVlI9SuJtpvxmuJYaSWK+EUMlvwzNPMC0PIQ8caYJLQHh47
PX7amfI9ExVu7HE+5VHzPQ==
`protect END_PROTECTED
