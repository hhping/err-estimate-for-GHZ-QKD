`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QH7IpxICo07LdOzbdQ/QBRvwCb6nT7bDIQltQ+1uENJ7BMpWB2wjUMOr/5EIJjs
JWkTBPPL0O893fAgLUPmonkaDJkhMkDkgRXix5e36Fuu85eIv/e5rLXESpeWTdup
cCXvmp3E97WCHPQb2hpj5h1I72u0ILSzB7rXS+EsrIJRkC902ZzEMt8igYkPjura
ztM8YF60HruJEMXQdL8suWw1gYnccbqUwYDMg2MmSvsb7j9CMTZdhqsgcB5EvH1x
1KDX3IBpxz7kBbC+A9xuEizoJdI2wmbKjbOmi0jLq8CkgYD/e4PNGGSXN4OJgL3z
51Rjhhxb4yOBHumO9eNsARqC/X76gl8qKxK9E59ZqzNzIlxF4j/ER4SaT00u76ht
Ll6AuZGN9BiFiR5qxhtQ/2JtZnfBkfa+aAroRHSxOcCY3QwXQPp/qpJvW6K154+I
dxGYdgJMOEXDtbH7RIrWWPhhgIUV8IfkuL3VyRQuRiGLQC5pJRZUkM+uFFHxRvT6
uM7jKODpX1d7DRStsk4UHtR2V5XesOQHChZRhUXSh6OKhIYb2EYrGX2BRyHYRiIt
yhFCD6vtZI85skSVtZOx3w==
`protect END_PROTECTED
