`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0qojhrMc04vtqBS2RuwoAyUaTzb9jTS42osf3Agv6tz8YGZf62j3WroodGaea1K
a/jCGI5KF5akkQaPWRYkANq9QLaUBdHinohxGEgwFj9UZOFXpgGwUYsHWLzX0lJz
wUaQVp2CdVrMNKXlncEkGU3yZsRSH33V/tykmfrvu3spexlRT1B2acGiebD8HBwa
REifNPYV5ePxPQqya5vaP0EGHigL9+n8H3mjeKdaeFh4YPNKpUmZQh1w/nzcniUV
p30YlZv71I9TMDGtcAvAyzSQ0RSIi1sZI3iLwy1inS0/wyvW8aOomyH8ObzCbD4w
NQl1P1BWC7K71DayQiSsMhqCdPqePcvnKClXaLwp7L6sICylNUXAg1LJMkrdUjX9
IYoUtw5U0kv9SvDiCWsV0f6F+KnGLgk8oVrezNQz5ILZhvdUKsN9bgoz1OeLVPpI
/LRUQ41P/NRUlkZnKif0dG7ajHH+/59/oNvBZGa90gvzIH4HPMkgh+Kr1LZfdUhv
fi8t0Edi6OB0SzII+JV8Eq6k5JNhhRFuMDYfbg25fOIJnztXWa99i6OE5RXbxmqT
yn4e/0gcnPYwdEp19XCfUXEMBVL74R73EvpiKRpwFuKbCEwYu4Wy9dxlKb/HzsFB
VJDluZFTut2AiR0lCINe5H2HiM9PXsH7tBJvxO4qFyXuGEyeRXG+YOnxDtPr2Twp
`protect END_PROTECTED
