`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DYyoZ4EOm+XzvBtw4SR7wikOBH1BnnFSKFRumgdAuZO//F4kzE6Gh89T/MaCSa8Z
s//VoPAgydgNVOvcLSc4Be/jaBwDVkzwTe2YYi4GD0LgDtgh0Pr2UG4rNsO4oG1F
tfw8JrFULwQXmG9CrWuELaEkqLVkyUeweeGymsLgQlmTxaUKntou82cCwHP/zSkz
vuquMHT21ReoyJ3pPMKNXgIXwkgAxFwMyPlqUs4wEnFhS3n3/6sXKomDHz74PLmG
C/0TVpW9biH2MFlVtxIROZxncut4xCv1RA66Xo2hZtPwtm/AI2AJbfpEnIHz6HCC
2l5CCOf/NhCyuwuAar0uaOwxxms7viL1PCCEkYB9+3d9dz3ghPHxcoDsE+Aunf9e
68YaLpi2ASBWqbk0HzkzAN0/+UlHif7G+7UZQvNDex+NxGOnk0Rqz+47yNIM9X90
qbu7o3tG2D711xvndWzJ3P2xPC6OU00zqRAG/L/R1bS07GUlxrGGR7TwwaFTK233
YSXXQWuxuNHqesjHgzcQxIV2w+/cFGosGeuTmQVngrlweOHHjE1irjcU8b4Zi14y
igdSvT1Bf9XxYNzWjAOFkM12iEh3z8UTWCIdBRfpFJaauADR1t+jF5/5YUGHA6iN
7CNUSDoKGxD0/q/dw8vEsxSJpeDQY+h+cVMG+5VMm71y/57xidjU2qtPWSv0b+9G
30kE2LwwGBkwMuWB/WFobzEYQlALYxhco84RGBWRYms4d09YdrVGsi8UkRQY3571
2QGcIsGQJnjisrnsCNNJl+lRRvhb8XnF64ujJ411KigecQ0W/QYfe2DT9dpihM+4
pdu9X5br0EBTA0O0Y0dk3IOk4+2Gj4T6fquO9ZXOGwBYZ7mec+G6tblKyhFLwP2J
P5BHTp6OfM3p/CU4GhAP36jWXD46MOQ3AIYfZlRwdGoiHLg+9Bhn9eKLnAypFcSY
/fGjdZyOJOhP/BHgGEmV19GgK+MW97a8Oyiud395wI1JRNNfYNscfU/w0q3LwXxw
Xf9bg1cd0dj1sqDeBRoMX/W8VTpDZncV83CpHNKrRjcakCryHVt71kU9BEC00KK2
Adjooi7/3DTe8e/EhbY3T3mv5KyV4atv2nTxmkl5v2TEgV13L1Lf4yecycx5C/6j
0ZTKuL7e5oCXFxre3zsK0qchG/FcRvgurxJ9vRtBPiVORhBMK0org3aG6QJyyWas
Yh/DWyoc/r9kvxjsQao44lfKS4I14UGsqZ0bBNiunKSDSLZT5NE/88bhAwDpEyr6
CCrmM9WNJ67YSmfJWtvYKD6MxoHxXRo/1PkTr/l4ev9EHrLgPDsojvJL19b+Z0eY
AOGfnmnsBW2WoqeBY6ejqJBSqLC900zBe/elqmtrj99u8nhOYu9Np3PwpPlGzzFP
9HdSvp7OmRxjQVUaE6n4zThudgRI38GaGt0CD2pxLS1lRmyu/r9WCYx5wtK1WdpG
uZj2Dh4EhJKbR+vAneWywbaoNkmJr6OIJwXldoTDH7rXsoFXn+Azxx+r6uCcIeo7
KfgrvnpQcS76/6egfwGrS3YZMJa33ogSk4FPMKFep6zP7qUz7zDc0VNpzR+vc+T7
ncoj+Kayl5E7UoFR9+u2uACuIdRjKrkD4i12upTsr9rdFBJ15wVQMq8sfZj5Od3c
5YNPy9+HImS/k0EJxuaPPREGffDZFm/GUD2vh2tKM7KUGDI19Zvpw3LteIcFGh6g
wYpaNcNzgAn/cspaEYbRXLNFu7MYVv7hfjGBCTV84BhIROBerseo8cnbGG8zz1qh
nDMWaDKzIcYL3HAhb68BAUObGBflJZbfES1MoiKw4bS1q22lSpDos87yGkww/cM1
mJ9NDgta1u69WMb4s5AkOyP/JJ2Ywm0Y3PdJ7NfcaIA8KkQfQ+JFXusbuy0u389C
B+329jcUQ0OegljD3K+zrXXh8jMV8s1qWsyPsaHvw6LbZT9JsHLh/15irCMux2vF
MwzGv3b2E/z2kQaBycjIIDqVF62XJPkRwvd1SEbtl8j/tYwO74+CNzV/N838VE74
C+nDn5k9SNosmt53GGqXvQGrde2Hq3/PazDFhBCtviba7YsXiCN279rNNfiAwN19
DEZ529txrgnW48c0vgNdNxlI1GpYzNTPMsYhrR7wcPDMkd92b5MXc+VNZNKuPYFQ
2rWSqvGLJifeBF3O3lTot6fySnZyktXRxv3kxvIiSxbRpC32fmvRCUiOryG/TQQv
ojrAWBawHxBgl5c6CGX03OhmbuAxQhcIN/Rz8TtGD1pVCECc0CM8dF2Dve7/U+6Z
ZgTeqYJTPPiWcBFYyx4SuxMq2qZ6e0L/JO9jC3wbhfWdueAB3Xg+53cm6TXxqL44
8hcDUdOWlBCw2XG9HH6YwqXp7+Qbz1CuKXMyd6OY995nubDKZl6nc+7tlHYQO/FJ
NPFdpPRCaPQ1ThKINAzf41tHX1y8hXeeOKvP/ZNT5Fze56xokwMKjtgaG6+wVcEt
wApbaN/GvfIEWEtf86s1E6MFhf6NYPb9LM9/xoWIURwUo6cryszumgMl7pK/6B8V
NEeRgHQckN0hiC7ofTGEHHib0GRgCEFqGklKYpySMFBMI5j0QcLNtCJ7pQBBZgVA
qVq9Q3rA2DNS9V4oJucR7jlKgkijxEQ9zbBIL0CN72YIxT7eFdVKlRPwQv4XqXe5
BAAyfjcYInzHoSAcHx625vT/PeYQYeSz1FNe7jP97scNdIH3QHMfHWDJG6cw4Xhn
tAIqlP7oooUhi9xHL2P82CtyI7SMiIQbMyY7dlozUVG0ewUKy4JNkEYbitEJ47TV
AQM3nE1Kh0aRNY1sx8l35oyfBmDotB4VVBQA3dDl+lpWQ4R9V3xyhj2+RDfI/7F9
XZeEfMQb79UxJ4DT09n3yMmBCjoVVbwUYJ3TOLDKVPEy8S8akeGKriRia0/Kgj8p
nF+x4FFAnOm3Sv95F3bglr90oXLNTDQKhifHC1ltRHL9zhuVs4mNeDqxxKj6/wmV
4xXGhcZFfGjE598zqg8Yyg8rITTfPqOoHZSjEuEql3aFW4IQ+dAC7BY6S8dzbs2j
G6GEiLIyVbwiGKY7j2i+CwCWnrv7ydw7gvdHBy1NL4kkzFFB7HlVcQPYov0MHtF8
+Z48w/wASnmHVrFElyOSDTinWvSAn+khQ+WMBpjnP47L0DxeuqhIZWwzWGL0O4zt
OXdMUBuY5iKC0fSpt7Sv0Z1mZcPYc8UD04/rBb/sN/ZpHpleWlfyvLO6vq3xBFO6
NvXGDWS9Ul6MSEaF+bghdyxNFArp+ao+TehcMLTQhVVVWvy79eWnY16nokrkr+mz
tHL3h5FpweNYu6MpduVc3Byg3sa/TG81wMaP81KtYvm4onargqCZTO8FEnolbr9+
sZ4W8/QOmKvWbklayd5qmZjJUmkE3LKG8qhhHBhrmXWqwXpWutWxRAa18iubXmaU
VjxNj5Z7uRN+IG8zcBPBMQ7G6HWU2ob+1A69qzpu0bbUsCFY92KGODpHKztfHHdv
TQPVRfTnV5nuYimEeeJRstgmGyKNG+JxRSMlDh/0aQeIqp3KRk166cG3pnSKccEf
L4RVyAfK7CYwlZcP9prfPS6eLIC00YH8yeCZ4VWPu7aq/rot/fFewCSBPoxS1/hk
zjZHLIYkges8n9RHIi4GnE7XXk0L1hUTY7Mndl6VShwH1F8C0KbQdPP831puyq8f
xk+uTrx7B8s0NAVoTumG9mrlcTAR6BUdWwyCGYb6Z3C4mIHiHnx8aiFqo+EHm9fm
hk2SrMuCiCuOoBK/bZAA2MQb68a5l042LMSvpuBTqom0fGHcTh4LMbKmNyQBQupq
6BlxtOqHcAYWn2K8gqESFcW29NDcU4UB2AFczB7kecKcCPWcihlTPLmD4+a8J/9L
SBvPcJUFKE+9ZEeFYgJxccb/MB/02CbKQAcDKLaINXacOB0KMYRa5tof3Igt9Xrn
+ZpwjUs0QRAARyTP8bbTbiQ1fiN+VeK43XRswxDufAHCE1EUgdcyzphPcyjb1msE
2osTGxkqghbYlg2lFOhQhnN3PCZG/WMqbJxNaOEIn0oPOgL6ZKZwz7VWjnWgovOJ
UIPlVpJomEZZApANi2ZiaJ9EnrsG2fPCJ8nkOe78z24YhqR/w1Kbwza/gGl9usSu
/V4lgQ2QZCN5huwsCgjaTJXASlm03B7/YofKHHrndIkA6uDsT2peIdU0e+NM/sfj
wMhhD4f/9xuLG8by8dH2wM8YND29DBDHVj30VCSrOMyVWaVqBXBVSlreVUBl744F
pmC+Fvng3w0pFgDrGbQNrwTfCy7A+ua7wuJSbTHZXL8pyZrzCJUdqbTQstY2h6TJ
ev1+rMZaepnsA1mnWb9Xdtzb1lRH4NS5VMHUSxjWJIuBS4lnaj/obfhANu8oZVbE
Xlt9jROvqGhvqCKAZurcN/asVDFyOk5pq1l73LmbjH1WcLxRWZrvaGOmBkJAotkY
gB9+ZCQtw44GYgkv57y8p89gZzrDhkYoA9lPrYfr/GD0Ib8f2AVko6H/ngQ2w0aA
QLOMYo66jRlbNH/PPid+1LTqVazWfoo0bWUDHRbHTsvKi6/yKP/EILJZV+Uka5F/
QLoULiQcqkg8WGfcTZzmky1O/RUIwEzWn80yULZAd4/C0bDgSenHhq8BdCYyIxqE
CGvxFrkB9h/MgrjFanLNlQ4xlny7tc4PNhaAFXYsfsNorMNNSig+C8pTxjsLMP09
XHiThVBO+AE/1FZ2hg+tJhA5ePMvzi8dDIuKuLbaWnSAU6hQ+tS0QwGbKLJgZaai
LcEYGka5USe0HLR8sJP/554vdE11J0VTopDU3Em2LyZs3aSx2of+/8e4XpzyJXi9
ExawwnsUXsWagWTg+/L7x3/ciugmjm2rnpSOxEuB4Vd6JcPIyKYoWCJmFBPR8Pkz
GgqkgG2J5oOYFRHa2Jh7gHimxjfKVs/xZIbT6XUCES+tAFh2lHmRHQQulgoEL1DY
CmlK2aNPI06Fpo3t9OMfAfIx6pUIYNzQVk/vU7iMJm8a8dbCM9NmlJ+hLB5/OXfl
aGk3l2MLWmALl+U2k7N30m+2k5vqrCl8ln4Ix0DDrmc2Fp6KkQSs4+fGgWd+nreh
yTzb5EnhAv+ppvfRX4SE67vnDxvmHgojZVnmat46zTlQKQJ+TaIZCguvbVJaUHh7
ex2kzJZwEHGskn2WcmiYlDfFe4Mc29ZbeJo8YllKYrD5bJsf83wHsWqI8YMdPJOy
YmpxJzl2yjYoikNGP0jeqgb/6lNjKGu7nihKKruCdi8UkLjcEDSG2aDRY7bU/Fmz
VrC2Dltr4sJqz/AuYu/mrz0GwiT8XHLlUTZmSBWvTtEUFMmiruEmiWWbj9mgeNKR
jUDes8haLe25i7pkcvD1AEeQisJ349ZfqKBBF0roYz5R0wvOBrnkBa/RbOaeD1fN
sxSG4EdvFtKrhGk+bmD7sWGJTJVV2vwiMc+GQMQE0r+EUGJHhaJt9HJ2Q5ldkoUc
E5vsAV4MN+DmXMahGd3mq8zk2PYvd+Jn4TtdiDWBbxMXkzJLyoUYGIN0QVphF+8q
zW3ji3B5l57laS34FQULESSDyGAvwjPV4EpGLRtO+FyR6MdF2TKsgopm1TcY/hfG
wxsIcYmAy4V2HEIVhZ2TteDbZ8hmQ6oJa+de+ZaIaQn9uUE7+p7+MRd2TaxRCLXk
fRQ3rpM9XRzmWEq7vJX/iPCWN2BWGZbBhBMVWc+KnmZmOzghHZ1jNmpemBbZ9AUg
Edaal4Rmt9nE7aU5NAHzxz5DYgRt3Qeukiq3qddXemOulyQ+H+dN6hr2OqfCGNFG
oG5g8bFRjk65aHsVsuLEEhGDAq6OZ89J/P3skxq0KsgjhXG4SZ4DAlBzM7aVG2NI
rmCU3VLg30Z86PCNaRL47l5J7X7P7C2vpbjCMWP+eKCp42TNGjnyYPs8MZUg882P
jaaWcri4oLvKeTbM1LwX6ZmS/pPxCaJ0yf13Y3gz6zcWRoEr2ftwHtuRC8ycb/MX
gyYrb5h68DyEmkEBOfO7AnsNO1a3Md6ERXMwHyJfaL0X8fjMBNQUP1PqKkjBDM1G
uMaBPBcn/5vrFhY8ne9EYm72+afsOwfrPTA+A6CaYWun2OA/OfPTClISdzLncb06
Ee5unlBFlIOmcmwMHbpymJ/vKkhuFdx0BmGMeKq4JotdWDmRlCL9LSSR3wf59PuG
co24+jyOkl/xHjQvnis44uGVdDELjaZxE/kYXCQOJDZhOEiVzvjVvcVhfmRGiHB+
huOKcmupy8seicenOhNrDJmEYz1g77ARtGLlYH9KS7uqarCm4au+Uq5HkA5RAA2D
R1n1t/bbFAdWIsXdVlPKIWhBmszIoDmT9a9x/AybcrMsyKFiZOclUjS9EFRBKaVP
HG7GVqsZoFo89LO7o1Mn4mc4x0XRQ7MYskxXTtwN4zbpgtwpqbx/4KddCq3/iwji
pfAvZ2IxIaKObUKxIjzyYGjCbv8kqrB+ONxIZKi8jAqmgwNNIXTfnV9YzdvKSgE0
Wg8xYBDVgoDKXxp1YTyIPjeViBaE5AWSWtmAXTqxgg5LGB0EVT9EEu1B1yeh+D0t
yKGFIc78gNbpx4vQ0nbMiPknEGqEESlhQ3frZMfO3Lbh33BVKZCmxvV8YH5ZnTGe
1O/ox49XLUMG+3MqVlC9krL9j57+WZRaf8+pf8wy98CUOq7+jJknKzsYWkzztFQY
vDX82t8/hfck1fX76im1GE8X2Go+x5WCuNWBcV4B/pZukGwceMc0mZno0aeZEhHa
TM0c0ELkbc945pO1S+7OxYJi8Dit+qgRdg4qEH3bP2tUZ21NmnGLl13LU3c9Cpf/
jQy0CmlRxMMWv/PrYz0V/hEzMjvmAEqOY4QNskNXOk0LiBpia7qG26YK5ZdssPWP
n3pzY5K81K1IoBkWIFvH6npVwzk+Sh/BHLEBbwzL1FDUby9HU9q/UKNyhRZ3sG/5
4jhE50o/jRqPql4K3IvIkQHAS8t7kmeS8urVsZju3mfEZp2Ts8BUzOwF1keqoUYH
WiNFN4F57nDTSX8PuRQS4kSAmDH7SPcaKBCrpeQZOGLLPnD2IkWXYRr4llUWsa4t
kFDg+/zxAzNQexvlojWuk1CdKSPqsHIf3ildmnnmdgEdniCIKrXIkK1FewjgXwaX
Wg+oaG7OlTjil60n9NJIwR3DajWk7gmPCdDiX3LXHvVnBS5JY5cLP0wNnjrXc5qS
LIFsxo47ij4NiAHELN8iF61CW96HYREu5n++Nj5vK3wy8hIE4ZES1eEg8cLNXcHq
IYYAyTw1udht2QKrjOUa/DVj3bcm9a5wnwNVZx1yN5mYwCF5z0wTthmO9vAqljh3
AaixE+t63fH9BSwtVrFPdi1dmS63Luhj34QIRRf5Kf4VCAiEdWx2RzOSYieSH1M7
WSlzF7ZEShWbsfB4XaR80QzP4dUpAjKMoXBfod6cHuvvRSfYrIpzOJdE2To7dtWg
3G95wWZwzisnsjd5hVHTbe2ttINeFMfn7xv8UBO4mo3iOEBW8WYfy7uG/OKK9DHF
TudfaUSHyT+ItOZ/y7X2QCSZpStTPflhvUJNOQ2Ez4aMLLmCBYoBspRhJoWRTI6U
+f5siKEs1iSVyfIREWHA2p5ms1BCMAti18Q373WSYSWxd4HjM4Nn39kOh99iT5CV
utgDu3gQVAiMY6xKB2rzaRGrsVdDTYMffIofWHPu000Ob0ZH2JccTLlmNVSjCm8H
uEE90I5aNvHOdXd/gBihnjS9wdnf/qXnMY4ci1F9iy4zwilqNdndmT9rTZCR3cg3
nV6bLUKudJ7k0IMeenWrkjqklySAGMT5GqZsB5loLVe+r/6+4BtEDpGT8wFHGaK5
jpo78jm/yv+YXaX6XcL0WOsu6je3Fc395wcke0Qvc5fofTxjSPwiHBYbrn0lwESB
vZFSXChIF0hgRQBtgv1BvxRfou+l2xHzQ31RI6vk0LBJ3V8SWUop0Lr2CHC8ussr
3FsBr4rudhtZtiqJie652fHxevzHSvf/5BQY023tjzxeHdXcfcXK9pS94X0KVs31
NfKdjGszDvx67VXJEaP1Kgj78ezjYriakPinWl9rvQefwIi+GQipzczKgNMUK8xD
iuVxcfWMVpLvbX2Rp4SwZjwYh/xICvy4ez6SN6vC8Z3T81Q8qtTzPR12+RGyDSyM
yrkmTJLjMnF1NNk3yLwtxVcMv8n344aDjWITAaMQds359f/E/dVdFuNXDSMo5+xA
jI5twXiFttX81rsJWU3OZfLN6tBsxsKMVkowm25acvKdCL/uuII/2Dzr3iz7x6Jg
VmGPWa5vBvIJIQQDhCskW3LYoWp3K0Dgts9aUnytBQciwoV6hn8mpHiHC+m1/QHD
GAs1VmNCe8pLJwxbJolsa33D5h1PEtVSGtOfsa26daQ+dm4oA5gOBHBVs2GeU1nZ
7dTne+5N8zCVju+xrgv0LUwiabWhY/ZgWc8zrz41rvH1yjqzYxPpQ6+TxTdTqbjJ
WsJzfribqu/CkWOztRMtH4YDTursJlEahMjYyLnsGLc+zsKeB0ufe+XnkvQK2zgP
9UUzGk/AKEcKyYPhti+autRL0RUKNspMjugTrk9+JGqwncACiTBKwN+NANI+RRa2
aSa8+1N6ipaRsBdVuJjC+0p7h0af4w6+X+9lcBSkxoo3VBL6a8XaPNcCSUknsnNe
kjNDMObcmdX+UXMuZRmybuAlnii0Jm6yqllaDv3O8Z9uL8H2j1k4ZtDGHZd6J7jC
+L00Osoxnv0BPK4dv/jQ8uJm/ZGNyogj8Q7jWAIfiQqtQV1HSfk1L+/gZDHzMLnO
j8qi4sRY4eEF8qtkRzXZ0LNyaTC9eu7G70n95VnpPCePJ02hLDyH5d/sZfdvbFXn
tLK+I6gp+y606Y2dnIJCmqBfPJl49B0mQcKP4M9SPG5QjcO9FfM/g1WqDlVVujOq
hSDcfAKyKfMbFpzXsys82pEefsXs0DtwzWll0YOG36LgmYdfVNereQFlvilsoUGe
4MhIR/7xREqUTox0IGMZcCTI82IIy+KUr8w61p9043QayvxlWYfM25X6fUz2MOrA
u0vF4Bocg7cX8WQDOZVrWSRGImVjH2cWvq5scA7c5RYsvviuCDgy6/tnazXoLVVi
QuQhzwmnoc3UdJeB/3OHjmJYOD0H++SzSVyUiGL1C0zNkvL2MoFSsH4D9GnvoalO
hW5GPbLuabMnjpBojjQBJOx6eF8uluL8oE2cBxoA25NQb4UXdEZWKZp+n898EDnz
kcK1M3YwIGKrB5p/m/fw8pNZ8yVLLGTnZVETJzK7t5k7g1kMY5tLlAJA729s7DqH
EtkZpnacxHSylGglFQvoac/wEg+jW/5J3OM3b0YIa2jW29ZIwyxjXY5N0QNl4zUc
zfK2N/88xeHQGrt2IeODSKHhrw6dHfkhh6RqSrsWrZWIST8R1EUgIMtryfJURUcu
B7w8PYr4Bok8IvLGGCzdz5vjynEM/70zcSz4hcP5asPL26X/T26r8xF1l+nseRWe
3oL3hyPFMOOgnBde/yC2h58rcQJ/pI+6/FeN3pOwBe+HBveatDfoFvloKSpi7u3K
eG3vzqwr65bRt6CEsAb//7PeDG9luHCsUXlLgj5DpchdiFWmmLwgaHFvXRQvUV6G
cj9zyyqPJB/iMsXn8tg/QLucdsGPALpN71YUK6vpqHTtp5yAbNm0ArcLBmGLCx/c
NGsYAT/w31+9bkdOeVxkTIMabRyuCq0TRB/RbEqI8ZfehNkaNvKDiMpv8zZizBXd
m+K2h4SqicvN+oeQzf9n1argDSjKKrSU6dJs9/Te9cJoIakQXx00JiHAF3MTquWV
o5ou5RbdIYLur0+P2VGfyVtXAqe5L66mfseANFgpTYIDXKLAjuHaLNcdPa5Hjwi+
oWF8SjotOBBuMWeKZhdjw/R2gXxZXi0UzACnpmq1I1O+/SmJycsFUax5wBrESoRw
/Tihj/EJZaD7LMwtwAydJpEPOdjgikiKoNphe9GrNi8akJ6oUw9mDVfN5cPU1/z8
234NozzsioEopLcvXV5B5Jjsr7p5tO4AarqIsh7qTjwvyKI3AcTe4fvL4u+WVXk8
IWogvh2ryEKKCz59mq9eHJWA3/Z05Rscok4MU+Na1AXgdy5GOFR0d72u9QDS9GjA
P+3q/l/xH1xdphs5Gpre66sFj1ZmAAKylIqiXtPTZ4aH3+HksykAXZZVe+PBEzV6
ehDO2ZoBlQqNrFy86jMHEFPNy8xQ770gzioCv58mUrW7BSwjWW/FJIubSZfX+7sG
sT791eE7xKnbo8VKdMkOmKmZhITyvrguvd6ffLOZOcMnx9ydauaA/iY+aRLGnhxn
bARR84ugL0uwJXUUd5u+PM2YVxl14CSbSQ3XF2KncHpg5ykjQSlraZLtDtzThdOZ
Gwpzst+EdRVuU4/ijSDxMPsADFm8rIqGYNUYPpw906a3HaaHhBtWmFNJ1lthi2ob
88uys8Aw8sjeVhjNgBpHJJMAu5ixJ0XsP5ebSwunWQ2P/onMH3wNYjAYsLUdiH5f
FzN2sZglTpQEcAZ5cwEYqQH3QA1RbdhaL0g7wgLclVCqlvh4tKVeg+dlXbx0gZ/4
JY1PzwZSGFBRIvPXW8cZbuH/FgPg9QtOtPDg1wBRlbcA2lp1MlRKF0AwkRfMeFx7
JWqLQLR6RF5GTScPgLqztGYwPIn4tpRont7b3t8YlmZfQk2Ifs87qWPpwESokGw2
F8mUbbeE8T0qs/BHyKfAQYN03jgURJQaaK0b3KACPYCLfEaUhZW6OfIUm3AiSUhg
T6/PXo/4LnJRlS2DqpUVQrn6ExrwvX7up9o+bWkhY7Ju63gZ2zWVJ8wc+H9CbOv9
SCjRRU+C1+wmg2Q9+zTqDMwPYarkM8CL+vjyrtVnZ62X5m6sH4/dwbHo8JGtWIET
9vG+4EJp+pQ/c5/1DvbRM8H8SUnoK8USjREoAlh0frpA0ylfQGzZq2FOyjOeRLz3
y45TmlBYiZnrXQuNiSd23LzNbR4AHR+ND6mpC5K/ZGmwlBMcAvcugeGN4sKIuUEu
QtN+bMcM01fph2G2lXEI1ucwhIUaWqMpYE3vs21A+/uCpwdslN6PqSHHhWLJ/6Sd
HLmJy8DtIsjgKj63BpVbKa8oVVpzk85uFvXZzTtc9eI1/D389ypS0AxeLX/d6Pkh
gyg2JWUlyDyce8IpwT/ZHvloAV4Je/yBFRTMdHQ/9MU8IP/hjT8uNqCLmILeDVdZ
mt3snubv6mdZmOJOXQLFVAnZdQ2E02bPbEigOT7rzgYXy0xNWcLn8/3aIYgqoZJd
/HarWr1+XSaU9j8+4Cp7Bqc/EROiLqJ2lJt/qmSYyypbV85/nhsGvzPQClB+vfeu
QPQxu08VJ2FxsagXpPMTqEcdGx2zkaLbYkkTJ1sRpP4MSy/UbvvObQfO58t6fG/9
8rlUPHszfnqaaRws9+fJ18jd2BpIKUHffrJ/2WmMxtAtpYDOVeXzBomwv/rzL7ab
Vv3ieXjDVDFekZi0ACjU14Y+PmREBxWNpQ7SlSPYQPFG9CXtBaOu1GQh+nf6d+LV
zmA+R60wpShk7vPCg05vCH2ENB0zA209SZuhBNc/cwK0jZArAkMniDF/UM4cPyri
BJlTaMSCOx1b4GGtM5FRh3Tno76pX9DjF5IYPZZ2mOOsgZrrdI3Fim2ckPJApbJr
RoTrcL5aNtzSZcvMrG4kpwpkiL8qO+3+Dtf2pqVo2aC1JD8liJ6AZok5BUdOcaFv
+TU4ybLu92oLo/DgEMHKgizbitOOsR7C5Ytw+J2vzEcRJI7V+1sNWRRqAkLsxarG
EB3D6AqW/5NlRQiVMn7q1YMGLOI+usz0rl3lmxoBIp0NBQcl5Cmk+I/z/5AcCeNJ
RNIRSvR+dkNjxZEYK7SSb3T8lz4F7WdBxYoB7h4z/hXs4mM3f/RRfanesqMso/Ao
40JtGMBakoAZBPKm1c8zN6VFEsUqemb963xSJIw470DY8TC1a1ssw1qqnw8RybIK
8ZRAhr0L6YxpPOx5fj5T2vu1IYIdp3wJB0lLMX7IiO+ocvnUlOOzWLP0QWl3xaEJ
0w/QSiSxHgjkNNjrN7yGAxZuBiN6GddZN/1yEBh+LNK+SYkhOn0DZQ4fAE7TUVx8
RkDaB25iGGzSaKxTsb76SERTBnWVGDFrlvVmRhFagAggagd725aQdPVyExH9oV2e
cnTbcO+jUK/kXM5ge+TfnGI58HMFPk3KpDsO0BpQV3nzL2Uv9MF/G7aWxpp4EF8w
qZTkq/tnvzeu8XAZUF1TTe46mtQh5QmW79vaFVrRLxIWwRc/406DlssTKJgUtyt4
9ahf8N9wKgA+/3+QtDLSMFt+ioAoxx+fzC6HeDY+IZ0aZ9hWKCnap4YMOSchBk+7
rYnJGOvY50eFla6yRPPP7fsSVoHwq8XJZKbTXeUQZA7tCLwCSlK7Ot9oWkKdNVUD
ZG7a/cjt4kmw9TdMuGdh9F/BkUgsvG5oMfK3gxXY4hDISI5zeh27mAfCfKJHjTmt
f4sDEwZKa+5KwbTwT/rgG8m/S0kMt62pug7Fb0gCSxPxGwW/dpjoZIDiRc2t/baq
DPK0nS0NhGqNfBs0fx9/Q9fCSL33P+kYxMr27PhqQLpwPLhbz+SJCqMT14tiMnt4
BQT9gq215LzUFKKJ0Vo0Z4TOcQ090IUXNbTHbNzJ3AMEqkRmMSrOLPesBUuyWU1i
fApQyQ8r1H6yrceNwyVjsXEsXCiJ6HV4re67vfSjItwWQSszRc4mfWZQzElF81lQ
MMURRMUE2mzE3kV2xrpLq/C2WUjFumEWZ9tBVpNU6ot+WVdRkaqGhxoSytoBSeoI
HDKq32b/sXous/VRCGyu2FyF1dTaScDr4cSojrqFu9dQdmAuBkTxwaoeoRj59VLv
jmgtd8hxfgytgiauVDL3+sRTJH6VtmNVrUU6fHvgSUsL5J0OWFJbtzcKXrSYL157
OvSakV+3xdMrbiRxfO/AH3pAlgwzF0PhUQrB6IA7DO75epVjSqxmD0GNTYQzeHS7
o11Md69nPYTFr6I0LgYMO2RS4mIPcbEGZHwyToOPRVQv7nKmwv0CMBy2e1jNUebi
Jd79Oa86uJvIzJlflPvOgARNJrDRvM3pavfLPn2/IR2LvhcIhoUE9xJRNqsgCLx3
JAEqQP7x7wfleGHRQkZptB6S6D0uvcS9iG3SK4WwUFgwU1612n+1TEwZaRKOMPdj
z/nRaBQjspsaTg18+N/OXIHuJIdOnJvGbcnQ2r3rxCxkU7k59RkFUElWfwWhZO4Q
c/qt1NHhcx/0biJjQVxrzAVAZS0ZDKc+2GcxQyl8aJecOBDnionaYZEZ1eUofGIz
eZ71HvZ0xoT7vsyAD7oeKTM283hVlcYakMVGmqrmgJJLguHzEZtp43m4s+McLqaj
QiK/YPAabcQkPD6n9KqYqclxFNgGpQi/tO2Y9F6FbzzCEX46BNJzstJ6Haugp78x
S8btgB/q5IeRsJYOZxIXbDLocsvJxqztBlXlbWw6P3Z+G7AQp/LgngDGa9DJzDxC
K2LOaT5eB3l8mv1IN/hWUIb7PuASnBmernTRL3tcxZWQyNSX3RFkmFnuwm0KJ8+F
n5NtbzEHlv6flOpYirbH3yXrdKcShhulByyh5hlIF80lktDE64jAvxbruoKweahB
lzWtkjYRPtCgriPoKFkW1VDRksJQtjQOXl1BSxjpQ3ZxZL7qs3MICIxhVfv5PWxc
Xe63ms8hBV5GCjCekfZStVShsZN9Ose71PJpT2ZG5702Dw2rnCcsk5g0s9t72ecM
n4lCI/Te1mVugsSLS0fiBDTNCJCHb/hI0HCK98yGzZ9mMBS+wD4MfYB+H6VGzyGB
UgIFxaOQOukq36hmbUE5+1cnzjb3lG87CxuAiLMuGpMSf41qSVvEmoRLUfRGkU7u
9Qn3F4LdS9BaZEfK+Jj9KzZWM7U4kT8jszdaWBlBpXZ7Wpimza+JC1HhIcO0CDMS
Xx4p424h7a9SRUSRTu1Ug86U2djMucfgrZ/MlfyVDlSdtYSoh/OXmWrkMv+oJajF
Y4oo8zvSCiZJDCxZNGCsnyzvoLauQdR/5SZRd96+xeDAQEbXnQ+lMp3AIFOm4TR+
1xfhBcgnyToJQO4+krLT43owoPB0PwHdO6dl81cj+hDhSUAqxnJ3PA3otiQZGqX3
ZQXRvxrZvdIHY0dhmrRUPzyGYF2wUaObPhaZloTCc1iZC40BdJjhmwE6JYspW1FW
jivfCszpqcW59bNxAmD5a2QfmrotMJ0Eu8SrDOA2YJXSrRgySxP/1Zn9JKfrajy6
jHwnHCJJPqIi3w9ozUUrbgymrw6oYtvbfu5Zmg7+Z/duAqkvRjs9fLBOFOZIcY6D
/LvATPuDFj5pQYFo9SxrpycL/UpLcNSo0D2UTKJniF3jpg1z9SD+rCao4hmdRO1w
wXnU8ElyGpMoKb+XBiSKf7FMiHj/mT1hNap9L5lalZNm6r3fHVCPSbA84SVigLE+
MRnlQeRd7KPqX7Yusm02ROef1WSfz05ZvCBpjl1tvyWKa/fBDqxOvqrKaVNeHG4a
EHkHUcsBOKuFueXhoqtZfOAEgLtX6iI7xf2y5G6iQ1MGECYL5zJuK/jlreshhCtD
4rtC2fStAeDhBGYQlC0Td3p2XYk+fy9Ime3MTp79n0f7G6NYXVMvykTD5PhQXkzf
Q/ka/FxLYe032aifPl7MB68M60WV/M5MsrHZ/I954yEzck53ORu5DpldYeTu0f3N
hOGsv9ayE5mioFffEDZlJn1Zv2FDlXmnnTLioxNwbCUCAGKfMHPbundVxLSYGBod
1J+4sHHqqzfUHHevwZ4IB2bQvTgNGnySKLzKuNs6NLVSS+BAA3bjEWjH3tX0xAI0
mPj2TEDAZZv9KXQOl1B8dyAOh2s8dB1XfF6WNHWd/j59xNFjkNII3msJ01iw/3lV
20CN+JLgoM8qEYFrVFOGYNt6s7hxxiA9n3wfnOMF3f41JymtbrZoFY6DtOd9hlzU
U9B2UU6PZHhHynTMjq9NirA1OmSCuoKszSWHAjcAzSYKzJhQy+5ZtZEEN3MGONcD
9BK0Gdrk5hRzUf0HTi5hcZEeBFGnRUkzOVaZcxxoAyiAi56is0ydebqGdo6T5lRN
kyF5W/NxFbS4/AgvROravn8DSgz25PxepudUB8/xdbKTMq8xkkEreeMV1gWQ0PEu
CSU3Ldu1GSzl/3wNzJvsR4Fnyzm79czDzq7QavGoKf0MnOML9X0ovjGSlFy/8xim
tKjITRkAPh4IjXl1HJiDk/b6OqU1xXwyF1yNJiabDYaLX5Mh8idmKPRieeUFHl4L
NjtEcbABZMI3TsZcGuwiYkVjseYMYGnK2X/TdreSkRe53qpbt/rEYY9TSLtMIauR
vju3IktBtwAnwsQVmhjsSEGmg8PHRKjK7pPzb8/yJK5CWg3X/M3ISn2Pxoqx+yWH
YdEoUyFnarqYz8gm9xE2vIObrp0NVQMSrxQsKCyXmDuNSd5IZJRMwbMvlgP4feAS
ZJau0mnFXM8z5FG2RJQrqhpV7kRKIU29+lIrL2goMmfo2vRjS42ee9hStZDyQu7t
5i7Vhg7GbhCZ2rqhWTvR0LvFRHHx7DwviJ0F9XX58K0Mo/zK4DRVw9qgAJRyDYoD
GTWoUONW7jjwirUybb0oDD3XopG1J++yKuxnNbSvTY3yE2EEluCH93NHVXS4EVNi
I3mc6WQRZrcUQFJVlmJBv8HoAIzTklYB8FA7UDQB+h4Vrg59Jr9k1j2+np67dgD3
Sg39ZhvsNqK6HwsbhLqOyxDxpo0ya1ood0KZwWCiBcjbOueUNkC/mwlV1mhDjgRu
iKKG/OnFONNvjFCBgbtm79JGw36EjTW57XEUEcLVgoGnHiInI/apjpt9vV3PBlPO
lrzGb5m0Q3qOFv/LQeiNnRkli/a9kgtC6BiyIZrYz+5b3ZEhouF3/lWH9jdUX+Ze
K3TIEbXT5bdg2OWH0TuVHlcoGbHf9o29TDFELeQXBeEO2dXRDTf/OJIuJcgTDjn1
ABrhO/JVts3OT8x60mBOc9vurosvR4PUHF1pJuPhrJk0rmeq//TFW0xv0ehAXZ1T
2Zr9/BmyTP00zR0JZF654wi7HTA8iaEwOhHMyLuz+GSVNi1U6PhB8ZZ3wFpjWwAQ
gIv4LJk+LObR4GKL3AbYTll/1GgTL+HI5t9eHh5iPdWvzWuCijvTANALheaeCxXO
MJBawdNOO7ebRf1AQaR8DhL0oIqQFNmmhNmEs5U8sluf9p0eL83ILtVKlCVFI9r1
8tazBPWqtkkckVpWijsq3LazmWAO0z+4To3xKW5Y4tG3gteWMX3dS63YqbfZu3pZ
MUpfFMWSLdh15thNBbYZfjzOu47qH+tt4GaYgEC8fQFaXS7cuwVttxvgQP6xULOw
weXN2MpBnjSLI5eLE0oahDPUdQ5p9aJG8K7zs4TbvFbPDU3HkjLgFySiLNb1MEVs
f2aKcb2CxAQMA/6GoKVHSM4rBiELyp2eeNMdefK1UihMJbnWkR1/mqB/MemNuLOW
Zk0ra2W7e8Nv8ZbrHXNXVUtXySf9ZV0kdGoqCTTFItPizXkZkCsnVKOeRZOcmpaJ
mHCA8v7a82EZkRlC3BwzB3vrjaDy1vz3ybUk8UXJXz/Um8PrUkM85I9igHzviSnK
fvumzeES8135jIZ67c21wg2rdV+ansrWTUq/Zpui82amDVjzJSRr/bYqSm+U+vx5
Ae22QL2zYq0yMQxYQHqUbzSp/pvXj1fpAYIkCO8NFXHWp5BMCS/3X8yhgemIhd3X
dc4xY/49Z9DUSdq2ay2geJp2NJOocNnhAR5tBE3ybfo9UCzlEaZwlysCgzCptjUo
5Zdc7f1SvLK9wetNc8hikRRdtqm7WiG8QJS5bK68eONk8/K9qqfwYq/TQReKvq0s
x3neTDG7VTl98SAsWBCvPMoq9QuLvVIPYQoWwbDMf6BA3reOQU19ldUSMAWxP2zp
FK6MyF5XChXFOwcXSH78iArX1DR5URhd1ydyxL8s8rPMECMvQHsJhy+VG7nZNFor
fKeuoR1bG2QoHKw4idnrSRUJ47jT5Tj+tGNwFXEq2MCMAEBMTNrr6rrVO2g7bjLa
G/Rc2r1X4tOQhO5M+6D8W0EuO0OnaqnSKGq2Iy+Mg0E6cy/LCH7fbju3d8p+qnXI
tndFFwj1ntXc9HSaGoSJkmq+/bvULDxouSsyQ1UGeJaF1OGXZj3KzPyeRR2TX4bi
637NeDj0uPVmK5BqJynARwOIevRe2NQDKt3nRrktN5/oJ+972Sc5F/JDxEheDvb0
JNVzFu07zeRE/QhOGZOl8uHpuYz+XgKucKcr9LcyCW67CvyiQJFNbyJFKUCrGB1f
8iCPwpKKC7nkIDLTBNeiRVWEIhQRt1DYKd6yMyYZyZuwTu07CRB0bbPZapk4bJ1Q
yGs0Cramhyu3KS6s7FuBC3j0/ncT5kHtLRMxO9GWnurdxplT3jzN12jCZ528ZUn/
LHAUpdx/P1Kk6TuEfOZI+2eYatDgv5dR4tU17nad4jJD0FsHtgtTPjB4THQI9Aq5
axNWBGTT2TT0vPEJkJl61Wr78/EeLccnr833DP6HxeiUtwcRIKtGDuz4ERQIYBC0
p77UUtg1L9nZma17QfwDqcdv7GyRclFSg4mQyfzSpVJAUBcxfjrg+7Yulecs6KUe
QtaxotWyP0Lq/y/TEIpoJXmGQ1gktOMr5oHIXcewywSsJzeTGVHV0WnsjeUFbzNx
MVt5EM+ZEv6zebsMNw1Z1HfU1xY+tk/lTFHhcTHgLQGpdaNvpiqzdhIWRkNhNHmL
7j3+5RxyOSw2k3FmsffXomT83KvVMLR7BoyXcc+OAnl1uyTwcbNJkyy+odq9xlWX
YNxq5rI1YgTTLm36bNelQB21W83Gu0jN4s3dUbsFAiuVjdD8SGQ2EwAntW6toQSv
NLPQDulgTGYcmm3tQz4LYCV09teN2GSGh7vbxlo8+gQybPXCr6bE5pkZe2uByYxR
q1aXJWn65RiCA1le8bashxMpmVOGf+lGjV1kd3DaBgDYQ3oBjlTO1Z8+pb4g7IP0
CeoUC2EDwn+13ODAI3t+LNY6L2qQVVgBFJ8aMypYZVPwOJCRAtRbCJSFNHvY5KCa
k7pRXx78UPgQ7m/bupoKnvMVoi3hOOH/EGmJPizoedNjwGSLmz6YpGyHEiCiar4U
5/pCGopzBSONr0Rclur0iGtuchAhd/oByTSCmrqvQ/TvX258wV0bDVDYJ6vZ1xcE
sn/osEz+LyFvwXsusQO0CAW/gYIoSrExr54gw31A2lZdUn0+oVtz4wxJtLPs8Bp2
rcfwRSmNX1se6y4SfyuMfeuQHaua0yd/a/a6h7BctmAOeokBl55SH32ieRUEyaUF
rqOKtlvdBzvPy6KiK4v7HOpss4wpJ93zcX9Lf75C/kJoHNpgKu53dM1rkNAxGwzb
2rATLwyIIqBYP1C8buXxBGJnK20GZivqoZzVAEYPjqIs4kujOMAK5plfz+Mcfopw
YqCCpVuuPr4tBTbX8zrB7ztpqoitsjX38H7m1wq4SmGm/3GPx1mg41dpycfPZMKf
VoV+8M4O2AB+D2+vyGFt0HRgTGHx00XaaCYop12diHEkpy37GNC25pyinROxKz/r
GQmkQmg+haI6MBEaSjscqn5UwVYPl2KEyV5moKPt3GHeC1AGGLsv+NT0Hts3PUHz
w7lzEnFGjfvsMLS2IW6ljn6Ny9k6BCG4rQqcaOpq8YgKYu+3ApG7Tx+4f4dYsvRo
8ThtAHH95vQGxxb0KSKZyVx3P9X8+GVn1/shV173Q7meHuEa6CoY6GRAs3yw8kNe
t+mdFMpZXz2UGin5ouY6TtxIXeiWsp9VrZ4h1reLwBzCqchoNsYujBS15D9KyZBh
5cS+lRoGu+qX1hoj7ztFLr7rmmOdooiymPsi0CTwytUBrRGTZAHrCiuCCJwkvij8
qf+Hs9/bvZP2qEMS8rUHyKlLFsIwNWUIxg01S6fBSnSEzsJ4c7xZja6S/EVoDiE9
Dv945NO2Bdi1NwVb508tOh+tz8OJfb+lVHQRPI///HIyITSmVsIADIIbGih8aJCH
//s6UaPcQYThoMTQirIXt05KrFNcNQ1JuHKyeHD830CegYLEKK0tPax1UORulyou
CCRweYdGh6xgDcuU813dRC1NHDuowGVM6GLrXgh0z9D0ywmapm5K7lc3qGYTkWW5
DOmJbXCHJW3WFCMVGWnRwQ/7HrvfsoC4TCPpiNlwhVIgjECsXFeVeSpETv6Q4O3O
FxTTc9lqanjFEeRoCkcOhDlz1xJnAf5+3hwY5pQw5+XC3uHjAiQhxEm8Q6NrNyqx
ZWb54zQ7cdDFe0QEQqZtxCz0Ff7b/JxvbnLawQjGi29SadB7cNvsFsquJlv8qTB8
CjndtJeMpIADixmSuTHVM5qX5XEXHRd0/ccSyRwJksdVQsYk7keOX/Xom9W66Yyc
6DoY9RlicFmmeBvyACwgdO8sCYGtvd2/LoRBOmKzSSpENx4bhZ/GtBpCh829VuPk
x2m+d+2dN/6t5WIjCnPol5L4rjUBatVqKmbJjOvxHHyv+nNpRzXxhuTJEaMP/eEy
poXNYndfr7ZcWwnNRDPtNnQwC4PT+B04y0/JIEepNKiDjbnIj9/4LD4JbGQ5I1od
joBhxhTAe2ky5iVu6/Y8HPW7G/JWBcPQ81qnWueiBg/1fep3apGjvAgWNyUodvDU
vKXKZuBwoXADPC/xepiQnkqQEgPUr/hi+sxPsSe09xAPPfjq/sOXo9355/wBd4e8
Hs0C0EqS06XcpQOrT2XhabI7qEU7Jr4okDPUFYSVtZrCvoGo/P6ZLL2mnFd6NMsl
UK7c2XsvzyZVU9KTUOMIdNv9WLL+oQbNtv+y7fU6AigvL2b01CRq6CF1osjUeGiZ
6EkTyg5Q/1oHfvaL//AMxXvNX1i4QPx8g6JrLyRUJ4NDFlPRLn/GwRMWjvo446Gw
0lNi2gZCT04NGifPCe8ILUuGJYQkV92dZRfYDBLm41qC0SnnTMjoRpN8hlX4JSea
RvQ+W7S/ZYAgimuUMiUBH3RbQptezeFJXjidrcsb5H3u8h5v2xLhtkkmtaPve3bv
8u7TXCKFz9eLFlpkT0t3CQb7f2aDGjwl4ZdFnpPDunlOgmYV4EAtR2UuU2W+Z5hO
jIi8ZTKEc8G1mK8YlSB4C3RP8lNdfYWO6MuAS97VhmbiXVmzqqyRgCbCHTjZxBdJ
/Aia4dF/4IQ3TOP/jkdyw0QhlOCYIPOvDIBkdw6Qy/F0mDyhbxpLsexiX03K8MUW
iNVvC+FVs/Ey19luO7KKu4nFC1vv9/AadNKXm8lBo9+cJT3Rfv4TvxbbbS24l1Fo
fOje0ThYXEx8ElE/9qsfVCDhmBGenMPWfbSmuFt8r2NdiPP5oaRJ5GoL91jyt1Ji
bhsaHqb+AO4EGpJloX/WqxSfPGdIEMXtqK4oiL50GdqDNNhstDCi9ppI5AozDPAi
s/RhaMa672KY4wFtnMwKJZCBRxJoF3FHt+epMnLGw1P2hkxcOZWjFjthVz6o+vMn
knbaSBH9JhtgkjUy+iqYrcpBQre0DLLJDkwv//Ea3RDqXYpvjkslTiNyr4mtPR3+
enYAzwpYWizRk0CdOjmu6X3gipZGtWCAChCZE6bMmUVI0O3JYmtCHgXvwSudgLpK
QbffRF7UgAeTzg0InuUSKUEfGeBDqsgPj9xAN5GjhRxDVSbEfyXtDGbtX2Ss9jVy
2WxkxTRDTdSv7pyOkG1jteBCCbtSTvbw/PLp3d0aKSYdiky4h/Q1RRNKG6KMYU3r
n42Ru1LX2T0F8IPaAN9jGJtat0tcWtNAXupodDtS2mPEn2bVgGbGf/kRJy6qDWdD
R+C4gUi/2qi6icU+YhOUSXlxMTPZhWBu2kjNqHQRMbiR8IVwlXZQZXmi7VkaunoW
jUqsBOmkudPj5rW+LVJh54hzc1kL/FF0/at/QnBgFsdO9IsiL7j+ZEycsRtaav38
WXzK9HgI0he2PYlIo+sfel5zFMkW3s2T2MPJrH8eImomkaJyicvLRnCMTz0oGyOB
Lakv8pl0+YnrSfTB0XRUscScorYn9enZyDMpkA0dGRfPCRcPpJ44aMHZdZs0fMbf
T3agM5bDYOzbBasn0fTqfc0x34T1R2ZotQMb756q8tqbcfgwn8zXvBjbzVhIuEEM
GNy5J8QT/R/uafYeKAaI7/icXbLbqBCxQei5uiUImLk2QkJwQie/L1W6pKAlPmGl
GmoxaoUBxWNkvOnEBV+Jwr0NuCo3ZCpzJ5jPAMXUmokGrgD106062/dbcTeZCL5y
B8+aQDQUhHp/1207S/ZxmuNvvKaFs9ygkWLUwr/lrqnNBEtuhLVBR2KzKhQ55d5k
cMjJFtfXu1EgWvSkkzgkrjLlSAxgN6Rzoyra1NPTXYu4WrDAdfNvM4YT4/JsCpR+
za/GTGoQ2ypMxwknTVRXBAKcVe+xGJSvqD5REDxskRA0lepHUQGV0HNnd3cQ1OvC
9eHwb67N8iCEltKzuqapL8FfyqwDeVKvtT1yz4AQ7pIeNsgmrVXbsgKqOnEXIAAL
b1VYb/+HkYhB++KrD+q1mpchlRE2njtOd00BIalRK/hnWprgdFxwxkikEE50RuR0
rL5BSRVyeE/HYr24+kT/gRV8zklN5o35blmHnxzNikwiwAhbUUKVIWUtxv2QO3NG
cLrRklVWkurdSEJho7g/oYd1WlzT+Dhgpd/uOab6K/ff/kECHOypCctXEqSgVX1a
iRcX2jO+EeF5qWneYqVi8cXKBOMwvUmbFQdt9XcLI693XviE69J8UXrMAxs/ghx+
hidbX/HYJdSncXpz/TIkiLWhfIW48ICvk06uIimyIA/xHWP/6zP/+VtFBc1JYiIX
ubIe3J5oxeJGN44K2mfLrBKayvo/kUJdOuEFz94kmJUgWmZLzPAdMl0xJOz3A7iz
t9V4c9Y91GKwyXk9muUXH02ay7xTIUcgwcgzHY0+g/HhiC29UBv8XHILrc5y733U
+QjdScQPYBenKS+x9J8Kp20aTr/RCFAXYSHpSYkPA10QbjgOLLd6vvoqT9JgR/cX
fq9qKKc8l9Y2xInE3pm7DnRfbBzCjO0PkUoc3JrrRUr8R36NNR8D7RjPk/5kzOEW
In3Nnl71xdzpgbAHHPalGWf7T9QQFVoglIk7AUITnNrJsIp8jmYq1Cb0O3CiMYXe
XFIZy8yNvu7XAqL/dhq0gg6DSkFAO8o3TZLik8EuWvO/s9HtKnb4GYO4NK3N3NLi
LUfGYhT7aVnyePYbiU+BqAFuquB8DECTFTQDtvkHxZMCiDhpO2MzAAMfoxo5Z8i5
CCMi+kHuNYNRI5XV/DcnHu5QYr2Y5zeBvfJoGncRWUvwtxFRDp0Ne6DcGDwnNDP+
DybJLcVkuUBBIZsSkMxVnxCD4VO3ZH3i980xqgt3FwSlDgbtEZ/6R/563zgSMHfN
N875mdyxE7B2C9S1O73QJuZ6c/aoTRt4+ubi4+PJxECa9CKSGeK/9yJSX3MLpD5E
addcJw5B/9uB6+o5yyM+26TDluGk7v2wKg+E19gH5EPcW96b8Z2ZiFSkbO8hEuDv
y2G1WjOBlsV8+IflXEWT5j8SwCPvGzppgqtCLlVlO0F23OB6TslFIb5+qrUp0y3F
Urr/qhkrGzm5a3NfLAjMtptoqd237LszrjigMpwbUxC7AxWTjyuVU71L3BxAXkmM
eVvI3JbHBcnEwRr9Ko8TeAVje3sP/+YNkUdYeTBmdZs3BN688MUxCzFUYNHS2ZEl
681fGdcAXs18G5EHouSnme+oxPjw9gj1b74o+zRIERhepNUZPNWrVegAkKI6ikzw
KH5IOYRdf96E7MBLuq2tiGQeD3EkOV/VgcHmrasKN4qT3hNPmEWIZKzGLRpjNz+d
3N9WP5cUh2Uo2bs3Ay4RMEq0bpm0SL6ZGCBK2ypXqFusySgXiQO/iY97RjwlJWx9
DJimx5kBpMRBCz84ubhwt9v8hg3hcH8MdN1gERO2fsU2rSh0TcmCsgsRJe5corwc
RuDIM3iP3lvjh4PGQmZWfHrSSrs2HPR6yLiIyCF0XSkdZ/Mb65TUW5j94ZZCH3PJ
hCgsdw2AXOqHaABpPWWkzOGS8g0T+wAxV5tAtDTL5GKEXhynhySQs/AihdCY27Gm
XJ466mjunsYIq9MHvUUdOFKm5glz2EJxs4bWdMYLhA97qFwxbagLdgi7KQggBtWG
e7glQvx8Ea5CFPeYrAqLa7LskuVP0AbOxnfOgo1OMWF18yjOIhJtPUPU6M4OtjVs
XtmQb2L9GcRTthUvWm61LE7VGukcE8x6bm0h7fS3JMNIvP0S+n354o9Yy3EN7U5o
CR2Vu4SY/PNxtUhqHc1KOO7ZSjJmCZyIjEO71ftgE/W31eXbPunxSiwYz7W45/jE
BfIxX+Xoz6CeM+B6RZaN/V7vYLORrCTWo1YAe2fGiip+I62xcyyYRdGmTwkQ37FL
rvYd0Zr7dj91KwaaVJCB5jVdMMi6rv0pDvEIUEfQjyf7J1YlCbWSYNpjhdHCNYvy
uw7TULYd1c+RjYmSOUKs4txFTRi+gFJt71MmR4QrJr5UWB6To0DR0HuV8WMe0bOt
ya8l1mZ6wEywnHuNy8Q1iZ0+YVvcqNuOVIltE2bbj7FXfbBgxdOaAT+P0p69b7Qg
1nz1xHXhpyAfiMsq2jvFr0akYkzsepp/x6fzprcFHt5ibwwRa4xThhEQbjKcZBzA
aSSBGtkcvVtohux8n6wnhQEw/wiEC1/g9M46LVDEJcSlwQYqHJAEcn+hEU3psSK0
y3roaa+gPoheWq7tlcwKI6S/oq3yO+warQdjsBA5CasoWAP5d3z1sPiNBt5flaXY
IdSf3s77Nic9tP4LJ+FUK5vbjQrZ56BRF7umi9MyGaqQVov1o6khoomqEuq17x8d
KUSVgEVQJaaoMWFRadaLPLN36XOH4wSo93NrBTcK1a+0q3K5LVinuS30X2/3LLXY
fnT5PLIVTX/Nbf3tGbo4O4mlnw/7BK4nnpIyjk4lDGO7+9OhTrhYynJMNQPUWYBB
XvOWtl82uifYO35c53pZp3Ss1zymV+NbJaF32cYgVf0doSJZWUCrBH6IyJRF9AmO
gRE9g9U7ArrPcQEn1k8uJoHEEmFfRtZsbRUfqZ06fSAm6jcUNurlolSmPMozr0+7
lZkBy2DO1FWuYBQoDN6j/GXh1alGVQVnLG0GGreDupLOA6736UuECZc96ezwEUWj
wBaiGHibXJAKYhifjg10Ughew24EMn+beDr79XCkkYlKCSHFcFZ7B0S2eXAF8YGE
mIyai6B2/FiuwkTf5BnzswAdjGKXW728IJzj6CPDzOgvIOz0smBnOgHPHtpcj22/
kiCCqUJ7KrWVXZ8FZDR0Umqh0LMAMXS8Q7Iut7E0XkE5xn6Nq9kdg0Lv95dGednB
xIuNGON6TPPR7xKRrMcpRXA0U5XL9nI0JiMkC3sDMmWUJkB3eUNrXSWSIg7UZ01g
tmmsdNluklG+UVViwxcuiAPqlWe4YvxXK2oMi+MjGJKTU7JIq8d6mF1NmQ7ESqo8
Q7AhW38Xu+q4t6NqFyXEBgmee2jruvjOD0b070IaEYsD3DrVIQ5Tzi+2tK0BwkE9
oOCMefozuoYjhsBebURyM28APxRprDcTgu8v5CmfpYvJS6VzPdJF4JnKZJQrAtO3
fAISPOVfri8xCyzc9LSqo6eejYkyrsa6YE9sJOsYt/UysLU+GqSX31kTT5Zjutyy
UVdGGEz//aZdB55oIBjvEBROU3vf/1bZcPlL1LxTVPPVv/mDXBCCUp/LntN/en4S
eU1kUVhHbBYvLLHeYBD4nvMgM1l2x8YH5WwrgXacrrMGlKYOFQ+cQIO3gxbrKMCl
3s7fJKOpdNspcakYvVDUqDOP8hrQIcnsmT6ksMN57XSBFRL1HsqEy93qMmk3U8O8
Nx310GdMzZpR33GyGeZ+B4ikFEeeht4AIXeIeZwoxcVs14gv+NaNbaME5IWEGpZ/
/yzSDEE12n7MUQzvrJkC6xSg1q5KodYCSRYx1ES+Z2R1N+b8LxxxnZmtShtBmL6U
w/aetIrGbKa30+LttqhHAwdKuhcDp4ORgMHnxx8+pzc3vrAuIYB0ff8zF/Hd8bhE
yIwxe/qP6PwGqLmsVlS7tFyipQWupaQirl8tkeyvyZHKSKhVbLFWORExhR6Wvmtw
JzLk6qbJcZr1lFsbRjMoAWXrIfIGZxsuhYPJowd+1CpG+zXD4O6gjzfJV8li4OHs
LcDkGqKq7IA5Mb5+BlOkyK+3DFeeESD25LIp99c5SIWBkjhbFXLbvWP1OMifbDDw
Xg53J2VnaCDCj0Yk2gyFRfJD3VMXv/1BPYvhX8a4hVPHf/L8M909NKstIDvAxk6I
Icdn/zdZu5IBIs7zwGRQMtvTyQCa83lV3snjWDzwAqA4E8hC7MqvS9EsSa//Gy/s
urXItcVgNvv1jgT7dTwBptFDb+Ezw4vBO2Z6Vn4Vy4nyU+8Rsahb3i5Vj3Kk0P1L
cyJly9N9KeC2v5Rghibu0F8EpCUnIB6x6iav/Vc8noESZlXjFXQ168ItvOyKL01P
DRYi0n8NnfGlmhoQz/JfjanHgamrHltMR7NVnheul+sVEd5u/AbNFqvTnxftIWIz
smM2X4eeeWLUTCpkRJ1xUpLFXx5CIFSSGuRObqYeAyloVMvnExBBLeDcqdUGq2Zu
8K3v/idGp1ODKpBYyk0X2B2ik2TJ0QD9UI2cbIxxGO8ciBZbRQOg9mscpRq4vKYY
qOBCivD51FztwkXUaaBEDAxlDr9i/34N8shuIIsta8p99sxc2fxSwpyCLDuhfB9m
16rQx6vBiswVltam4WZNrXjkouogM5o6dU3dVH1XjBEXABut8rhFt158tKiUPl5y
B4Okt0up0yXQe881xutQFGFopo6PzkHOg81klw3jbDIqrFcPDQYCnK9H5/UVxIsy
z1r/X8lmiOYWzvgxCZMFkSRoaolAI+8CLE5XGPU9/kP7G2SaHB0Sm7AQAPXoKwHE
zOgCaW7sWJgjACnP0QpU2XU5uLaUupajAh24YQWMlSpLl4vbl5sM0S8+Jisg5Haa
SNwqIlQMh+Gb1YvAwy19u85+X9iprUQOCitIBIbhSnuo4ymdULQ8l8vHz65SjZsA
s0ysXvY22Zh9kx4q55hhq6Qeuk82qBlZXZNXQHiMW4mq5qXnsqtzGlYy4ZiLzuJT
dcH+mDtY/kWpT56RjbyIZJURNlrcu3eAYPPBUngZqxIEWTd7oKHl6j9jsHAI1U03
6OdTk5BTSW04jxWOtYhngGkMRo3x5SbwavL4SENrzPV03AAeuxuuKkbyslgowS2/
m+DgbBFJ/jO9Y/HYMuQtS5DLA3zhe4MhLM1rs8e7hZfTVkf6lzh62FZNVz27Z/7y
XsI19orQiSR27rnbVhcykaBsuyetCldaixTU+12mnBGBlgk9lNnhNUixfuJXQeAz
lcSuh14h26apQIZ9c9Xr7hGkxF43hHauPQO/KkOa8L4EvDFcd61zWpdFr6cOlq9U
61FModjXh/pTp7i++s8jxIC+ZHl7qODvSVJK2L3ijlRvWAkPKCLs3KQN+MTaGSkO
gftVlfuu2AJx3CKYWn9ZtgTdM/zJ/y1huk9mHWe5MbE2VLAGJ1IHQB2d+rPI5pg8
YNTu1YeB2wNcn+FCr+y1O7bHbTQwkQYXVRcYbOdWTw0Aw/lX6X91suULy3vRQMhN
p6o3Fek6KbIROjc3RdxoR1QFCNORq5Y8/aNshvO8vv3gwwDa4C5IqqCaR9QDk/XZ
RMQOC2lFxfAHo5+Gp4Pl0z+W3AxCfg5T0lSZlgvduxrwQPw8c9nUv46gZH/FUsg5
FfcNsrWpHrz/5Q++6bDE3axn0pCdnm/lXzWgF0uIWVH8UlqMKWhSyZgakYNcpTNq
1LS/uqBSahuho+NPOoF0bn/g7GZmJW0bBJkmHYdjGdzWTLYe3+DVqH36eMZ2h7+m
euyHfha+a0KtWMmITXNNvmfpKWEZGSKtyggwc8An2zkgTTv+Lx7gK7GDG9tOz2wJ
Za6ZptfGyAHH7YocB12Cvnmdesi/AEF0Ghx4Y5fjC/MCU7XQ+6rTgG6AJEQs+SQg
mzHv1Anp3HjREntSkLPBF0N0VYachtsitPArdJQmrrathxWYk2f/ezmJf+kqaflM
u8orvFjB8cAlMsdfLgLoMmLdQ5sHC1Ug9y2eMqfTfbkWs1xtmL9NN3218y6QGyeB
Pn0dKqheY+ghEnM4grRQ8g6j9zAls8hRw6H/VlZ7RPQ5OrUN4Q6Vt4yQK7Sta9kE
tFCmeU7PBB0y2nAud1s72ZGRQ0JlM8oDrJxaWx1EnnZPZypwrdi/+NfPQmlHoyTU
X/cPKHrb5p/oT45Odlch8dwnLQNBia8XhOkQzrR5PjsG4zFRebadM73nionpCIaO
qgAcSSHdFskBX43ckPXEr7gMc4q6bW5qRtuojSWDhqIcQ9tk9atGo6U7H4/+D5yP
K/CxmdQDY1ilAu8dPgWGV9wQoW6xpRylRiuCRAijuu2X6TQUzx9SPlyGU3cWdqzj
txkyBocLiQD7McBDd8MV9GYmYViHpB42w8eZU/M+JREBNqGL5LtBX8R2sEQpKfsB
MKQw4t7TDuDtS1XQTIj65auykrwyKigAZwftnx1LwiCtBbohpXZgZ6UHw46J2dv9
bSwxbeqqRQQeYxQ3+Ny0gWqM6n++yuVDhKbz74QSPjIiOZecjDVLUFu9V6BCkoZ1
9nSuQA/gzOpn9mPVAt37XK+qC8LTVnQuFk9WNYUtfkcrDWNiahhMLwS9/F4Jv5XN
SozQvazPNGElQ4fKfaKkKNQGQsxEtOBe0HvNgZapv9Dz1FgCFLt/9akb8WA1KbEp
ZQ5kEjvDkckzZktoDBngH6ic3yHHozyywUO6hU4srHWYsv7MMkmqQyMoHb9Rw0W8
SgUCemhCzCVtKxB87Fy8UQqr1B3Nhtnz/xK4/JYHk4EvlVT4s/YIP6hts668gLw9
gxvjWzP9BhqnTTYOnDjr48MZtU3zxkG1HgDZ1hM4icRKA9pyLS+gPn8l3i6M0cZO
6JI/7WmwRSISFThSwHNx5gYKrv1TJLFlTItJ7ViVpCC1wkq8Np/dqYkUYARtCkHH
0MDciCgdYKp+ctoddhs5u45eTQnCbm+vYC1XeQjnyi0QDRh6q2C8aamIXv4SbA1c
dTsKRk/8IvqgyZOAf+CFDOGPsME9shvgamJgnT2UhtmUAEqopLffGD+tTm85xszl
Hy6D4ITWpUFMwxm6OInycJFeWd/Kb0Hr1NheisLUTQE6ktuBxE/CbGvxWS1saeBg
IiGLXUa7KezXniSOxH5mJ1GaIsp+b27ibio6l+LQz5zzL8MXDTXt4Krs5VKKN5U6
KBiVMv5PKO5hlMMHNRzt6Itt9ZQmW8C85D4vd/mlvf5XBZPj5dsYzv7lAB+CxmnJ
iyYnl7u/NTaL7LnhOCIR4zh4XtUPEPuHkjWujeh56MrxgwwvxabT1q3zXr93QriH
BU4H23kwunptAh3FXf1uVsRTs4daPgNHynqHF402inowaS7tf+xvRBOVfbZ0ehWb
t6iup03pwIO/Obqk/sdUFDi50a2lVf0J0owsoEngikRLnmHa7s4NiEJIOPXxnw59
+JlssCUFQUSdYapKs4DEF7siaSlJymuuknhXckX8LngHoK5XzBdgwUsm/JTOmufO
Aq9Tst/CLdCY1yUNZuxR9yXuOZxQuJ/OHJA/jMj++n0WGYjTxw+UKOeorKYayxqQ
AXxNzrLoKzKVx9iepk5NSGOq2CqOiIQNX1qfn2Xoecva5QuZm8rmmj8MZifplE6B
5eL9+gtGwd0GK7EpvN5FJhvhy1r6VIYM++s9whjw5PZZxGHtVnxkO9ihlKbr2Kyz
HZVHeHGBwaba80EefnZZmhxYwUeY1F5QLG3fqUTXo2giXU3PEbmyrCbdgeFXsi4X
eHSJrtWsYVI5ucqhjkxR2KjV/6iaYONzUB7z5EPKNv8+fUXL2K4G1HZq/5v3SjHJ
0FGkTaloF0PgiGOtt1xArDVw+q+lY0+iM5J6hzQBkYZkpHJlTTuedEuo30e8z0FH
jPEP6Y9IeMKjAHNynBB7jQDj5IXag6YwQC0/vX9QcIWcJxmOd3mcjDNq/WyfCTLl
MM55DFoQV/1NQCRF1/8+/DUH7y3mbZT6JocnSRzL5/raPy4Plygi8qUI3xEu0D4D
f9DlyuFIyD5VRw6HmiNKjdcRTSW+iMSIoB4CfnbS6irx4P+CS6Jx413Caqnd6AkS
QFJfe+thVWV5IbXdEvLTVmN5FISQUWarwu5iIjj14YRbWBLYOwkxj/rVReVyeLhZ
X1GLZNYPhdYPB12CpdZ703SWEpH4FAx2cNtZYtyWCNVvYmQVsLHex7WmjL1uvI6S
o9a5rj9turwON4t3DyhF2A+zzixBCMXF6IlZPglLscCCInwg85fmZ12WjmbnkFc2
lfUfdWxnfMdK03hpGeEa+SPCAcRGAA5u4mg3pXBPmDLYQ1dTOFbPmDgiYGHNqD7x
Gjzg8ExdCIbDIlgiK31P515xirvJcsxvJ6DlguZr3bZvd6YPmxRkuk6GzhIH9/eW
MQzQ4jTyv5txW/lH1hKMcFC9sBAtq84ZmlWTx0zzz3E4pN9w6so28FLlNLIWU9eS
33H7taoT2v7uw6MP00Qf3w9fiwn6/W95r3conboFWj3HiS8N/uc7RpirFaeSAnLF
l1WBmsfDPy4NQjap8Q/EJd1eOMwRRAD2R1ufpXiAYzRFke0QFhuBIRCX5w0XTbHM
CSYmyiebCfMTypggrg4imil8XLcmcEHm5aEos0V9M6LNcDqlJA8Jl3xkHdVyafVZ
/STiVJ81Sk4OQSxYzJpstpe2LbGw7G01a4243DHki3cHwvGSEvar2YLL4s4Y9Ugy
a/kM+spTqvqldBU2B9cJGTRHYC4UDZK0Xc5a+dipJ4bu5/uqZqI6fJwSgircXNQK
Hc9kcfNpjQN0f//jvkwla155T7SBfvo0CP2gZUWLqATgUcgYXff0ErbQCHEuR7kj
wbzYhWxVDERJ13K1otqAT6XKng1hpVxLj8IlSwLxUKxGoHhPHw1Ii+WoX1zQft8U
i3htgY84jbERoq9aouif9Pxk4qOSi/AdefBBuo79Gkjatk07oFARypPig0iHidf2
g2YAhf2M5bo0tOsx6rVkJSNfdKyfo1egFKg0LnL6LzZY86eF31OOdx7VJrux34wE
YDpiqGAQmc4FhI/9xwSBo9ciahaLu+dsubxRSncXCq5ooQEVWpDwcaUqcJZjv5kz
YXmP7OdiDY6k5VwpPKxpe/jGIHZlbWfDh7fKaW+uuZKVvnDkIeX9/xnWkwgVCL9U
I3r4+41F1yBeXIzv9pE+NKUayGRWhi4nBs4Tmsh/Csh23wAHu/5sNNh1DCi+9c7R
Pb3T5fIIerlDWtdnrQcE/nzVBwXMggj4+K06tGlVSKs8bw2ReBSqNamCxxTigd2D
+15wS87T6N8PwAjVheoL6hYj47Ngj3jqN3Sj67sZVx8iJSW6N/qdPAKXFebnoW6W
xk8bUDIWVvYcqxroUo1h9uFPHEzbwCPfcwB4SCZdD4PEkO1NyuLG2TsbhUxXnxIh
rBK/oletxL1xeMTTm3g16NEfJRSvuPJIDgxpfC5xp7N1UniMCOD/482W9q5ssWcQ
fphGhicIMS/m19RHP5umYqTrConeu+hwskE33zOTz42AlQsTDK3ONvDg425mPhJm
nUFYSmSj3DAG6qGQsYON8+oubinbnXV7MpRZDotNKXge3v+d+RLQdWK1r6IiTu9R
BR4AZ4FYbMxbNrv2lm4DRhq5rp6SmMz5H4sCXRWZLbVuwSlGR0/rsFyvN6HYgG0B
WwY4EKP1L1rk7JlKxmh86127Oal5o5hqmlYHKH2KFGP5aTQd9xeJg1qLI+NhrJwL
YBNuYVgZQGeYRu9Khoi+mk1/A5W1H5n0ti/ZsCZiDfFYtZYgm2BHepiNNnS+FCBs
NHRIanqnfYXM3/UZNorx5n11WbN0y67Xfl/PfJNhIxM8YXKq6YkTWQxyJVYZM+hq
OIr9XF+Ds6UsE5KrkAEF7OpBZkXn3NjGcvHmWtqDyUCfnqsdXMD1Mq1LLTaMglLJ
jHfLNaNHjLbrGTUVrxWmySgN0eu8HhaqXwuKlvlQZvqGxvRU8EArpEiliJViSLZ/
CxqsFV6Qo14uJV1lMMdUV5YYYV2jPMywkJ7LsgaKVdO6XbcgcJaNH7hVKZkGzI2n
pNZd5Z6wzBCCLoDU2dxJV8N2lTpkBMGdIuE0BLFj/oecndQgkE9OXXqi3JW8+2vr
VmVJRJL235YYrJSQY0XNbQOcu0vMbpkH6g48snHjmVH6CsnszaL4FSYFhGEKBGl/
R+y5Z023iJg0MEz/U8smiDAg43hS39gszy0HopGvO068zk2X/+JHgUfDrvF/dwkR
vhJ5EUGO3rU2zCodS9IrX+bqe6NZ7IOGCVyhot6yh1f/Q68PB91pNhBhass9lys3
NAlsmWf1XNP+h8hstWQR+kAA/KzGurDwYkRSg1YJhm1XeFpWPENJpO0ycZF+uhVD
Ej3Op5G9qJTlFX0ErLRBXavu7MdxSb29hqilic+fqwFtY9kbZEPAqSzxZYFupZnG
dHLdds2893aPap4q+0t+txHBrh4pHvzGJ4GIWs3M/Bnw/qBZTBkhtMpKYFXA2XKb
Jc5Js29SpbexxRYF6pHsVluEk90yaJcpUevQZxCoIsYme9m1eT2apJ4uS4sp41Cc
V6TarP6hPp6mNHVUY9e7ZtgRT+LLnEqiwLxjqo6DZaGehI1Snznz3QHu9wXL+zDr
YPW9phgZmK7a+s7Qr0cXGfZcPVxoCJzv/Vjrm70C6aLXz7aBOys8kKb60eJarOz1
9voFFXNi0nXtCDNYwLtKUNtp8k5JbWK3afjNK9XP40P1le3kX/jGcv04B4vQAG+P
t7+yeW+Fi1HSdOCUaz8PpuT6E0GmZxnyTv1ULwgogU3V2V3EmRarcKMbjNVMysEf
W0yYigwEWb0n5nIMwEnquclnwD0p+67uKhSZySeIiz97VydpdPBjFihQhwK+1SkD
7gOpB/f2D8wNnRm3qYr0rg1gs7PcZrWIpK5MdBESgZjCaRZbpM0KjRZdD9sVuiG3
GxU53tMTGzOdzIIwNc9wjntMsTeJkRwJAAowxXrrAW3ZBk+mJXOfaz+uXOZTr0e5
93K3rCmrK6YtcVK41Bk5f8ayZIp9mXccIpp+z4RImdJsy4Y7R5XFkk6s0Va5vz3W
+fk0dJ9peVgjrpcW3YHTSuU0/XS/d5f3aROTK+oFN+qJV1a4RtxwI+SAXAnh/5LN
6kvN8cEOMng3LF93z1MeKt31hfCE285t5MeCb0kes/7VsOS1YVrw/95mS218LDF8
5fMUupnpYR2B/303kAKbs2c+zQ4CnAx/GxQfpXzYemSwQlro14KbGQc5f1M/c3qi
qCBLo9olopkUQZJ0aZ9NHQukJyixXLsIM6MTjCdKMMzS1N7/tRVTyGW2b/CkjKT2
QC0jp4cc7uTyCsddoWUJoEccPGuOP2+P7Uo1fy5fxws7pFOua8ChsbhxaThoKtrb
N37uSBOOHO8W/SdbLadAJpjOKwCscOv8Jl7x2BURzY/+M3moC2TrMWWywY3VKNOS
OJjvL3kiUu8ivi9cn9HDGGiExl+geAsZl+xb7/Z7XEw7GPXI7GHKBlbNZxEITlnj
v/iWsU4G8+a3qW1BwfcFssXzJqQ/DfKAwRb1Oh9ajE6Jx9plyuHW4aCOBpVUfpRi
IVz/N2hkB2rXL84mBAjZ+Aaw7gZtISl1iYY75KTrPcFU+mTWQghTYe2/Rg37Gwm4
Y3romncajE9VJAJLv3aYZz3ixfAQppERKllcZJcaJto6v066G2WvqA6aVF87n0jP
AUTqkzfUWAyqAzRkijyDavU1ekFKsS+0ERq6E6w7poh4pC7NjIVdp7ukMzZoTl1k
czAiSKFUxsM6eJrkO6t/2zbtaQ5xM+1lG4TuolJuV7zbJFUK/N+IlKFXAB/+JqzY
ksIf+WzgBs4iAfOqVROKmRob8VI82/Q2w96+N189yr2gxU8231fH78Yc7gg+xS3x
djpNRQMk9QnB0e/sp91H18316fOn4g9cJDO8iv48Ddp3ZhlC5Nas3+9esTV3Ir3D
KrOoeMMoXiryQQFlSyJhFphqIlPwZcK7joAajPazIZBRWxTZDjgE5tHhrwuJo0h2
txfNnwbOuMsCU3Vhw/8Idlol3p7j8IrTFlsYENNDZnHrZlDg11SaL+t+xvFUCh93
tRT36jKYRkJzn1Fv6/dJIo0ZoYPF4KN2UAR4gyv1EkXMghtv6C2+aEJNPwkmmJGv
Z9eslDPPAGMyvnoMVZk5TlD76tOcvTL0hzdz5m/NiIqE+I7HAJ+1cBHbplGRcPGg
1wu0YHlgvicqkdjT9I3b2blhRy0yt7As07kjMBdyvx8B4a8aZaVq05N6JOGBigLr
DgUlyZjrIvbjQ6b4//uGLfJWw3sEM9DTFJxpNuSCK1xTgNGM0HOAjGabRpVTk9Wh
NLSxiML4JnOOnXDcoe1gcyY9qJFHVG9NZA1PcaMYEHvAU9HE7IVH3zug0BioEAzz
rHF+hDjt6vkkX8kTfUm2zof5i7Qt2OZ5vhw9pkEN33QtB8dzilrPJVcyCDc/wmGu
9fnVIj+WHsQPR/qqBLI0FCk9fTivretXNAf5YSoEeh3ZOAvnoUYjEOHaLuVwfOjI
PXA0PwLuQHDL2YEwtFFAadXD7xFPYwGrX+KshNOXfsyF6NCzSaSZd4P4j57xRmMM
uQezT3Ki25CPERnD07bl4hRRBwsApOJ76zOVs/UMEYudKYwsDKL9oovfpd5nuIU0
fkbCTyfUv5566iCA9AzKQLAjnxhfh84V9mlDrY9mAo02jMN8r9DhTeLtZrA/qbQ2
DZ+1utkt+ogwjZGvVtz+PPxrIuV2BxFf0N2vW9/pQYaNy7ulbgd6E5Vyufg1qVsU
NEtm+EwzOml4TFCBzZXBYADuxh4642lRScflpIDInRPzPPRnvt9c4i73iBE69nAc
00KE4eiwTF4qtQJGZDBEoymuM/SMIxAFDr2q77BJc7s+ez5iygwsxKuyjBSM8HAn
4uMG5Y0alnW9sfDsANs9AVQ/fPCFpQkillhzbCjtJUXbB7fIoDhKtsNWCadcwQ9B
qv5rDHauFHoMGLUcMW6tYAeqM4zXOFM0d0Agu0n+14StG0BcQy+3PK1BpSffLsSv
LKlSLPU3PDGxGF7XPFrCSBlecfUX7bRsFzeuFrX77OiTY70XMqdVeH1vLl+BO874
AqTlmuLBZstXgb7VIeHYmPTfAfjZShYJa++eDvKh3AVSG6RRQcM155JhSivBCM85
Kb4RBzG9B623TbmS+HvABcZuROQyTyZ02kxlthC/FCBEFn+bhbwWfU72h66ou7yG
3H53KVvwB2QfzVSbW+BTerWWr8c6JAr2NOW/SwfVC0xWB8S/J6J6lAm8MTSL0yUp
TbV0OF7rXxDYViQSNKoEFL2B17wAUSjv1cgfDwF9fevwJ5zTQlQnCfknLnFol/yr
6uf+q/XiXFMbgghvvrcaMyDKgQgQUl1cB6CIAR3FaDmWgxCofxF8LbCjjavOrtoJ
cHFh6PjUgKs3aMkCaMIogvxF+k8V9RjJMLzsQZKsS3WDKMGGTIDIPfkcMBQWgwV2
J3cUN1lq3cCbliTYlktqWW9G4Vz3fgdjxTnAnQe+6zN6LgzGTLex6zoXJXCiIIHK
Me+yh5aSFaPBvyMEX5tT2KmtVqCpJIqC1zNavmjQ2uOKISt81qoh1+HemhJOCbwy
CAd3s5RP2qxZj7XKUVAOAh7+2dPmGZoKN++oYjMRaMOq+Ap6hId3wolMS4BxQ7Ih
Ve+vi/5JI25+yeLbJCHpZJUXw+abhOlckVyXhI07uN2dJAtxqgw4qyz4e/A18QD2
11D5AhkW0/8G+2zFDB+zfEbSlsvT0cLFhv6rICGzJ2rYgEhPVQUVfC6HnXzhQs1i
ZJSeP+z+VvoOxlttEEih0YdBwEctZZKZxkYv4Wp+VHptc+6flxgRHdiuO0TLqSNe
JbFMxqKd3dMwly0H0ge4dM+pqSn1eJMKMx6A/WMkztEN2DPvIwfqTAd7MfWiom1T
TRQ6aTiO+8/TG4di5nKk6UxZ2suvQeyoV+D1KCrD7valTaVRjogPEYuzryjuzRFi
c8WhfG8rRcI92vW+vinv+KfoMJv1vEX7xIm6n5FjJu0+1hQODw0r7qXfoeRhqaLV
DrtKee2mzGvE2+zhmblo25f143ztlUUb9AXyIgwPhJu8lUHl1VbKwQ/dV1eMSAmp
DzmgrK94YMXWlGgob045Uc7Z5KkDO5s5PWuCRSA2iPZBWNvJH5DtEKznFBP97JtK
rXvpfLbLcrtqPNPTmEYtAp+KFTCpN+dqTrEIrF2O3Lll+fQjnKTOWmS4kosvOiBg
i8UGpU2Z/o4KEu/u5atHdwZz4C2D4cQ1XFIPMRSrRWdn9zrCm8HDi4UWk98h0mFV
ultoRIUoX03t0/MoOg/axJL4lvzAuHmBr2gtsnj7II45s3Ut3Y+lOvrXF1ZfyyRr
739nE3dv3oorOX0zX7snV502f7OTLp5g0x6bsxsvEmHSPr19HVb33RoQcbc8ElQX
VC60bnRVTwC/X+gLIxw8jjw0OfJzkn379BxURorNQnOACRDBhk67DcUGViaQrxtw
srSE/8Y25Ta6bng15gSfah5H47L6AgmXZtO8xbm8EFfFtbVVypoFHb4IZO8oiPlw
wMvjC1W9x/6wkiq9wuDuZmPMjwFBQPXclxlMjPV6TGF49y/lRNXABKpWeEOfkhJ0
NotdnmSyjTo6+tX1xJVIVd4J6nu0iwiyBrVhQ/0aw+RHqlYtU6ZxLoUv33He2UND
wz+D3rCp9btTGbRa1u+BYZ6wTE3G723YJ4Fca2ca2sNq2oow9KXjZ4tKH/pj8bXq
AMm7qbcz6OnS31jhB+w7yZEU0DOwjlfiKyrB+fsMypfiHx3UDDwcrrVdNClDCMY/
QWPhqHwmWcfzUCYEDfdVspcY3/cLytJ5mQcRTYndZFQOJGoqjeZuZ7s4eSHZjVRt
f+2oK7zBqe9wgDU7qfjbhuOuns/2/TqXwpE/+jA5ddK0Da7EdQTOMNWeQCmDvLAu
FEWm/CQJ8Wl+NxzixV3F3/Kj8kngYCRcQzWNHxoSItBVh6jdd5IKmmMz/pyWAKj0
fcAXx/LaTpxKbtCg1x2AecDe9a+QkYWsUvdSLWdLkhz4Q9X3/zRPcyLu/cls3E6z
lUblIAjA7JHmI5MlFgddEYRu3XnmQTKuVq0OJU3mxtkJBd4i4an638BUlDbf8Ypa
KcHe7k8e+Q2IGnJcmgKlvYf1OxDGTpe5yMivRyfDlAMeDMIrPS4OcSOZ9H2uLyy6
3QRlFJg7VO/sC5r7xr7FfHPdaV5xjxHjPCKUSLWvbV10mY6itIa/7weXNLLjctIu
jUN7/ZUtREW05hQc1W2T6+/mCrDIiupghA1f3O7UejWNUn9vhg47S12gzP3UcCKG
gqV4nU+4inmN9JIxkz+qVGlvGV2ozsxYlDaVRcrr0A501v4tyA1uOaXakgaDB/yg
xJj8gGi9wxqTLxAPsAaGeRUIAo+CjqLenNuE7a2QFj60k/SzjBpvUQiqz3qblyb8
ZH0mr6GrITbuCX5m9eYgpMnGYeZGRyN9raTtkfHKNu/F1RoibJopc1iMuekNce0u
qFl7TGsmh4sWf81rnlqqutO9o6VMzn9xtHXZBA84q1m31/yTPHj5n+WX1KY34nY+
mE6z02D7V9kjRp7drlhFkOfVGL6XLKOr/Ee3jl1BzQ6aC76aM843yxwOA/k6xYcF
11SCzpwnbZQ84hpjDL9Ze4Edqz8p0XVn9+ursdsayP20g/2Gas4yDzNpsakNmDmk
7I6c5uEAFKvgpEjc72NaiMh8ZRXghFPKhlt9/tebn8BN+cQam7BQA6kwoz1cxYnI
qS5Xv5hcvym6GlZp3YKDOhBci6rTRJr26whbLmIyMiDWiep9gYGD/wv/aNPRsZIi
tYftbREzyFIfDF3m5sn61KgRnaSvA3o59oDj75nlX16HEKgBiT9J8qBTpAC34gRW
NegDY2e+afATcBK44t4ZVNU9s0dhjrzmm46F7yx1XPHvUke+BVkaWg52PfBRRcvw
chxbt/PcJ1nMeAbjXOlGl9lqWqNwIuSHzCRY4fmcWo+cv/nqE4olwdU6NeHSkevO
eja5XWxXB9kUOwUbhYfBeiRqJQGoE+LpNfaLufAERlSMcypQ1i7426yFcmLePmAd
iHbztYle8dOaHd/+JwYYupNiBnbYfBmSCrBRDCsGIzQjXaCcOcK4zj3eYSx7MWQ0
i1Ndlwc3djuq0pjXOlz7BFFmxu40Wde05ipfKOSVpPnEm3Y9E6ZotadxJeftQ7sv
A8yw99SVO6llTyb50PhcjKA4XWr+/l5RgejubbKSMDVm1vLio0JHwOLejC6fQdC6
11emNuXs+iOARvgLRYX5OPt9urfo8ELJPxr84f2Q4mxJ0TiLt8prUE+z1cQvm8U+
s1qhz0GQOqDeOhAuQoqB9ezIK2JLdcD8pLP0vj1dPImKITqd7QBiFOxNLVXEEGHV
R9W49op8PjROZzwXrLdRCH6pklQsgvmxajQboN2BFGAAIaiqGiwoEzzG32pOIhfY
7syWBo2F3cCMENH7cT5h/S0Z35TUd3Atdd0Qsz2vXnEVH1H64B4Xj9CDKRGmMPIc
APaVdKQRAf3t8wH55Hm9WtBaXaQGP9UCzMV767cHxkPi0KlobYe7z0AdKbW21PBg
ZVZM1iD42HK9eehkYIKsreLEVtIVDNstl2sr8yZXS91JHs1Efs74CcZYrdsMbU70
fEXGAJqlO0e30cVlZtJXmTQ+jm1SsFzZHgCtfC/LZchD69cjR0XyoSoVeRlvSjR9
gXu6vda7zkqLCH8u6U648XjhOYfxRQunzwzRGJAYMUK2k7WvfzhqVOXxYsvibUgO
ZYgkzkkxemPJbHxCs6b9hQMjC+KSZschuIaU8yy5bVZdUHaN6aa6syXNY5y9NscJ
iVp6A9gOEGv+xnZK0VIm5BVKNr1SXQG/9wjFWHTR56uyGSLYaFzKgIQHUTemCv2X
63b8/KUZg8ouT48jt+ED0ABMYh/kG+DZsJc/oFsqSZstkWe0LqueaOaBKwRXUfX5
iNPo+qAhYXFUHUYGp/pQmS2ijC04MvzcFYMW4b/gM6ZV2Afs6aXsFndymWfNXCtT
8JRpa/Wy4GYp7Bdr+o5JE0t1jnFubd3evco+TEabDLebz4TbjFKCmq9V43jrGcic
D2nNabcDWWiz/8xtiO+j30Bi3vaKR0w3uYxmVPPeWNCCLSZ0nniBek5Ig85eUUIS
c0bA0dhCZl9NHYxs+I3fnxzk8SJ1jZ50S7Zxsg/KZZtTajv6CZggAw30OEUWra5Q
+TVTwkaejygeFvdgQ0VhRARxk6xaxlSCY/VrHiRDEBLbfmf0d4DRYr2mKXiuIsip
6+2dLz2AJ5cx3fWiYSjv1e7gvQGH5r7sohHzwbKiiovVb8lxz2n8275HY1iIPiW0
ihvkWJVCDACH/5+smI0csEAO+L5n/kqwLcgKwFaPfyoFZKWmqTNapEtmRgSw4B7i
Rrr9zCNuenD0XNMIkiRT2CnUcL52HQ/fv9nHxAsemE9GlpBZfy9neMg9juYDpK7D
7vtJwGqkDakI9P9i0aDXOoGXDupyHsp6VhF1raZx2LZasS6hk6HSXLlYVg9uX902
urAUU72manyfiLbv2Rs4ABeCPdz0qHIVp8cc5PEdB2CBj9SMirbu9YSBM9/7TQt8
KCyZSarZjTMKD+GTP2pSuSIqP0clK+QGTDcyWC8iNztTW+ZVSrNSPmL4Rjpf+OaH
VX7VrmHe1grsWW+yNvcK/epVZUCNqm95dUBq/pmKUWLMOd7Gsr5lF468sJEVDhZT
y9KRFh92XxFfU2PVA8p3IPiu0aWdx4Qe+zSeRM2oNGqgkqvkw6M+5eAFZg75vblp
XBVi2Cs44TCSIa/h+KP1l/FA83c5Cn5ZKblUA5c8PU+un/iRckppMSZQeDj0nXlu
MSQoeRgMx0m2xxWdTgmtx8q345cRsHEXmRFK6vs+7rg5Wn39WFXpa3k3a8/MFvha
MjCEbAdKHHHGGosxMr4QVfh+CF1Xb5hGFjQHQb4Ab4jKhfwwZK1Zp7MQQLNH7RI5
T2yrVTfh4UeWTDHdsdTTLC/aX1DVvpDz1DhNkIS+KwNhCJIEUuFUbXvTKls5ONbU
kUoAf5qVOIkUP2VCPMKDU8STasEytO2swGVHpXZHJWQ/ECPguwB/pMTZfdObtJHB
MT2nCiTe4XLcyNFaTMMHxgMwmAiSVhFCURqLJ8BMXMrHh32Ly+l+RNbYfiiFd1Lu
YtXsYtL+YBSol3c6iovXuCG1RKiKVh3pJ00HJHY/ecFvRO57vZUYd7tFjJa1bgSf
eGqCyHCrwzMD3VcZya2dQQWxx7OI+7whn/232D0k8e5gGXjXoXYjmxZYd9vNp7jT
izC+A8l0FyZkkH1Sn6HxaAwsQP+GvLIzUjGOrj5uFnumqAwKegaeqECrh2otffUJ
8jlnoHj8BnVGdqSzWv7qIVUvqIG8VKYn0o9j3nPQYAOfV1mT5e1X16e3WU0YiYNG
tJgbWHTy5DiUnYuBWrc+AxFbU68ogPTYqfTiBwzxrc5RI06x46HFzuRfuCSLWv42
NVhLu/M/3v2ExvSO42SFViFVSjkK/AIkUMgE3xTqKjdGrxtGxBmieH0XuNI93tRF
ZOXLzq+cwEv6d2N1oTl6rPg7mcOx7R7jjaUBlsfn4NC46aJyYLS0j8Y/zs+WLbeK
jL4ERd+S4IX7GLokdRHTyJ4gCopurClYzk7POvT2lZTaEklRX5+Yvtg5pTpq1D3s
NMPT/ypd82XmFXvio3eSA+WUzQC5Y/nAbbQQ0RnUHzuVkbmg7etsPLmWHoeCGJ3L
QzBXFNZyyZKq3f8JftBqKOEmUztRFhqf7D1rvzV76ADjh3NhhDWa1sn3GJC9pmw1
Vh7O9bbz7vcH7cmwbUcxDbf381R7UhrUiN8q4aPsDZ+sm0Tx4zjTTqlEuhc2rl6H
WjvM8rijT1khhYR9fC+i/cKugn/6yrq0q5Rm/RpwV5mujZEDG3bjiMoCwELmMhzj
PyLm3AYK71h/jT7V8i/pfbwUmXKOdWQmH8cX5OCVBwc0QZDo5PL9UZIyInjsdO9N
u9BZ6uxEZnQC/bSGk25HslDkdxz7R0p6i7Py778r59hqWf72kz/Y65WvK3gLydq3
xxwVzs/W6QcL/tXdAccDb7HBE/+P2vPh+SSeAjBSn7TBF9rPMSgaan/bu3bobb99
XnwunesZGXMhbCS/9avXlzgG6MFjSKMuJ/ft3wIMY/jJI9iBusgAtHL0uvOtbEX+
5Y1zFgBQwps+WvjJp8wGREVQU1kug9l4SniDxIWH282PWXCQlX9n6wXLuiTT63ui
pP3HWi6Nyj3CnX5Wpkt2No9VuHxLfsYWp9kg83E9C64nBB7bT/G5QjA6egZiQeCt
ZH0rbBobc74spJGRPdlZRO5zrdCMctThzo7Hgw7kah2gcLDqzVFio+9RModHwcLI
USKfj1lqpZidcv5+VDTKq4yjlqkULR/FDfbxbWmoQ76Silr2zMj+KodJN6dTfJVA
x9tfuW5Ie4HQME15gqkRuyjCiZwZx+EWTUgz1yiENNxuBeSPpt78rZLONG3T6k8X
55AEiBkS0Ux161vnwg4OalnkqEtx08KX559KJdJLwK3j3mwX3oc2vHMw38He+5Yj
Duxebebf83ze0folSlpsLDiG+M6iKAOks8S9H4tTb6ihUHHEf+Fxhb/Ol6aK1/37
bYSzFudEtHAvQPXrExJPrDioETdI0dPQSINtSOOB+a9FjSXkf1LavpAUawLajmmE
KWebaqF3D7MEDwDsLWk6nIHtO0RqiqQqQZaDBF2vezVeFnib0nJoYjWTETyUJlw4
ei6Bm2IllO8qW00rJeVqD0XzI5/ytAEuFx4NPRKrgNB11yDGcYVwMVe3ihV/+Hvp
imEmYmGG79mqF78C48lctwniUnzUVv9bvZxs25PWlAlcmI357R8U7VBXh+eTkxOi
tEvXgWhabdMfdCkoAF7CpetLR9CDhlkYkyAjwLC1axbDa/0Zi2HRISKRzoPBmN9I
+NXMxHbODsUdZxc0EJP91ZOgxd5bzoXTcVRzF3YLjlhgEdVrXzp7TxlKgmFHiKZW
iVdKF+LVU8LveheeigfkA+K+wdK6Sr+DUg8Pv/CdLC1tUNJOVKrJWIM2BRBravQ5
4yw0T7zeuOwLYKBkMHpiIynk4DEsMwj7ntnsscNqMJ1LmKewdcklf/HMHkv7mVGC
x/0HHvc5CaX7Ymu4QqciN58L9oNl/gF/KRxlAPfmUdbmrsJspaN2mef/eFcSirOc
9LbAugPrB7hCpWCl9UR47hlYc+ewtW5xealm/L9E4g3neQAYZpw5qM41prPMx4ri
VFzGGVVgpsbr9rt4k1yTyj0snhRZIbn4r5TOMsocPy9tqxrcD0QBisHjdNPU8Bn6
wFhgL7dXN7Ekv7pmM/N/12GZTfc/+GH3rXIBZW+aRKLBjyrS57cgbP5ZRTRo+TvE
tQZ9FdNUpKCq1Fqxyqat/A0lakQIRjQtHZYogMBmZyCrNpO7an2AzPEPzQE28KsK
sDJmuc3oGJR/lqQz9FUIWXkmwbbRsTFYnhlaSL8r50WFWPzva8ZA4hiljPqSjTEd
XPgY/i7wJ/cSr6xk7UiWV+lOw6tRhP44C/JOXR0zDC68P1VLDYGy7V6eXhduj502
+poR1DyrNLP4t+CYqPHdBtHaM1RfUpgj9APiHHiMDY1VlF2bGjEVlPr4QbM51HYg
ckI72pUrCdUswJJVgAVtUsBGN+2WruxAOJNgTq6HIl4ehzF9/Lq8wUvsQeCMc3SC
DFl2X3xahxmDU666YA8QK3527qqgnMttDlAYU8+PThZVBE09jR2SsogV4MaQNtti
a2xMvQMYk+SETn0s38qWE1px14sGr1mKzYfM7JQWrgowr/WF29RtuCW9gf2w2R4N
QLev7l7ASTkmm4yGnJM3BwAul3yL3qWKlTJm3EQZm1+TV2/O5ojZlAdYZ+HAKAEJ
zWI5oVVN2gpEoxHyA17XCfaZquwJRbIRkCZ/B7YBsr/3D7JFjTslRtHhjnNe2i8N
wL5YCK76KSmrrm+jUkh7SQ+OOX36l/Idn90kg7BSP9sLihkXshndCx+CYhNUzgZm
JDLgf+uvSvBe5ygLU+nIVzGL0dhAMjYcEHGBJyZ2uPueVYmMSXCzd+Kohqto71/r
K1K8YJr2XcbRXjDPv8J9ZWVqGj/YbfBWYQHkN8oB798+8ibm9HuFtyS1gNoTunFM
v1jUgvi6GAxfjypG+j+CFxu9RKW2PNjq1cPmCdOzd4uD2NNX5DfrqIxb8OHFP+6u
uaa6zdl9ijyTkU1XqCu4KS4P2IFjhliKTmqpy/bVvPWW55rxppTZHiMSBTWqfUIr
2ywLjOBFWE1ua+NPs6KRd7wyMs2dJY7bw18pwxH4Gkhxtmk8B+NuXSERF6gP343f
phVvutcJt2sMkormSMWMqvE1VIV5GtaeTO8+V9ZTT2r3mB60ByZRaFoiUR5qRH9s
bEKk0AMSiK/3QQrB0VI++z570XmlKi4bB0YIw/QTqfDNZ4Ex/HBoaoFnNI2EWu4X
R8+1KjY7sHBySNHD/7Epo8TGUhjuN1lwspDlIGh0hNGMBKU+9wmnex0dgFE4j5vE
KFuzQL2U0sbCCzdFnSQOhrHHO7jJckFRGPwMksfUXeQev2o2jdIVqfUDQA/a2Va3
4XQEYlXb5rkqIrDMDKcBUG01e0CiALgM+mcqGPIxl4kNtF4QxpjvhHQguaejHxoT
XPeg10yGYbCnZHPopx3bcLNHbHo2qBIuwjtwA0jYesRWrNSV0/iHZXxJvHBDSU7x
JMqHWyecV/DiWBwwf/RCf9XedAU/Ndy4pV2+1GvbK1JEVWKS2xdN0++0t4cof51X
j3wVEI7cdRdXaaERKieZQNuC7ZRC0aFqQJNcoeYGHgOakPCtQKpTAMfcrk4cVFrB
mCaMxbhTOCphQA3zLkyb/Fb9AS0sWRIXcoqWpyVWQRDKiJG4tYCRKI7CTIIsFuT2
AgMIE8GTNf9DQTlt56rSHQZtGPNB3GhbSrbjU/6BBW6FV1lw/KA7a+1WfWsfRGwL
rJdPSNx8CKm8qfjQ5vtD2hIePHIkQgtWlNe8B//SyM4wxxG+xMb/R/AirogTh/e3
RdCIdl/ecPPC5Hk2iWoA+YEfHGzuwPpRXELz+m4Rn4MVYaRJICILef3QyIy74G32
5V2TfsIaXsnr6P5SO+SdifvutmAoY9eudVxrqmpEnNuHX4slGeN6AouV7BlqetIZ
DTSYfYRwGN93g0DmmSOTiLHVBoe9Y00lQ+14cx55mep72ayC+B1iv+p7x9Yh/I3N
PspTxSlZ3H/DcwGBVUTvg/bQUIRnuC9jK7/LUGks81PDnHKR4qJZ+jTmcFR0Tb5e
90sij8qqMyOszIb+mqtHhs38qOjCFHspGA+mPgWazPHyWgSiWKT9RVY+KDgUS7rG
kKD1mJug1/NPJ5gex131bBc+W7044Yj4KKx7idgeZHcmAYcTMcY/+9HmDPpMvKEq
PUAbTnNFx//CGk/9gFv1SfdXJUP2OUMs+GR4a3GmXGKvFiRhXy+pHiq6qsHrpVL0
rmEnEpccEXnh8ow8ZtZ98CTqGCxRW6E03Wjns1E86vkNUkvZwsG0cqQNF5nAOkgk
QzPpIbZMyer9O5/aQOsEgHeqawYdpXNQh2PaELNK5QhAAJUIP8Nz8EbvY75x1Pb4
3jec62sHBlTMhrz5WBfA0Ei+1xz4Ckxgtz3KUlwNfJ1Bd2JymNgGmQTyO5npCC3S
w9nbtDXlZ9S+47ZD8CMaxP9xpckX1epps6Qqj9qYsG8tm4MvCgZsYkbVw40U4m7n
Ma/d1LrYtqHDxte39ELioLe03nfn5C3vDBpABLa1ZklgQ9ZvtshrulxXotnkskVZ
iTbmZT5VS01WLduXlCVEi7bXD0caNlkpVFUJ8z1k5nb51ShBGa6EnashceRF+a8m
Q4pXhGzKinEoWzBkzE2gncIquxfC6hiAeHYBYTrL4//Y2MXIvYcn5lKQkM6eqq2W
V/KzTYHTfZ10HH8vw7sBfxNJcx9J29scrKTw1IjUQp6t4AODBwiv7+oFaUHIhrSl
e+IVXcp5TO3MS7hSlNKnkRZq9KVJM40BN7D7tQ/XyswZh6MpztkgrgyqVpxXW9JE
IRcjxLV/D2g+4Fq+Uj5C2CkeNhWXsgNJ7DB4R2aPmXAbJwwFKyrum/m62/kVN5F+
HcScJNiuTgFlIcXqYMDqaoiVIn43CRnOrvQliqWWh68OOJjWaNM7unma4kmji/9p
Q6+nHxoS5ul9vJIdwH3zqZGcHQ6LEbWcsyh10A1OwRSqgKf1k1qAInUepolDJ0WY
8hZufPfQsGYIM3RE4r1IdPwHzHiMBzQBCjoNQ7dHrj3EeMffZ7pfKr6aXXsxAl6d
cHDdXMBdzC1ExtKsR926VZTEb3WKb9+fx4tMeJ3Ax8q7G25nngazpY1N+mFtgDl+
nEw0AYEDoXj8Cw6Ad6LJAfjNia/p1TWWkSq5BvIIH9zCfdv3Ag8jfRgUKaTulzVP
idZZRRWwozegXm5CuOttbeSRBctkXTXi+Jn9/+lALGqy9MoD7pOyuruNdoxZl882
8XzH8W9/yC9GVtnIKvM+9NPybD/6p5otOaeovz9I8nFVmCTYb4kS6fLiJX/mxeK7
0fW8B2c1XHSno7WeT7pAaxK5hdj5krTbUfVSyQ+C9ArmB8UYfObYklcu179dp/es
3Ka9fZ8PL+SozWxJ6Vij+lvTzCu2ngdpfq+tdV99VNmQhz8ZFtoqEgQYs+hoz/bX
T1LWTV55Pxzz2CGY9q0Geeiq0EZ1hoV/raDIooqRpAqytFZd31RGbE2/BySc3x8x
3TjGJAuYgkPfPS58LmrGwVcI4AO8LynG48yDrsggMGpNeQVN8E5L83LGokI+KMr1
`protect END_PROTECTED
