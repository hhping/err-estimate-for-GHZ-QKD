`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPKaDh5XP/l7FKGoMz2CwU7IoTSjlovU6nibXzBAwtDZgz9LoL2FX4tA8Sb6GY9G
nqW4VIqYsgyc1qEVD7hTEE/85iufkefMpq1YmCWd9uH8TlTu+5fv5V5VnMPrCp1H
Ub06ZVV094MW/ouBkSVdeNGN9/qOOT9wVlSx6G8DOE4q0cqUI3/nmojtpM1vx2Bh
nrHdYpyjaRRMCgqon8CrKWY9H/Gx5Etm0FVJvofx2ZqJc5kgauXowJCIGh8XXMUK
JG4wdSTZf22tkemM5SdjSIFbYJGERnJjtZRNapdtlC2D+XVTflc87VU6d6jO9m7x
fzm1+Yr0dOMN7orL8g50McRTLgFWo4QsbCmScCXMA1f1TWlPZzdPu/m8z8NPTSY/
8af+aIP+Vf1LhdtkhTW4R7caYV8DrATzg9czdevBInxhgeah/BgyrMZA1GJKQaDE
FSIKmbl7AhkDxmM3iIuTTGEY5VtqZdA7IUyM190/chOL3D607GQ+RWEcTOfj957Q
i4FXYwKcNAtgXdFaOS6KwpOZ/aMuk9EZppyYRE4GI9PgDmQTEo+oA/d9aDUYhZy/
vPau+0ejAnV6rEVGlhB7f5gOfyKj0xrtG0XSMzcVGNazS6JANcZWdn6yJdJyvi90
xbgHNk/bvlS3l6aCQGyp1braQgwjcB3o8mdvBQkkl/f/BfHdAzEcqiNBUR0+eoGY
iQAmXCT4CLQD/irJ3yxUKV9sM2KhRXWRvEdDcABhJZaCeL8UAMgl6IT8jreP4tmz
Y7m33m2laljArhClayA5gbThctn6TjCePaCxHcYJ9IbydrcRdfl6AN0lACDv+ENM
9n5XW09MTCg5bQHYU6wIFojogal03AuC0zhzzMHF24tXMJk0xRwPP8/kNID9r6wQ
3SatTspQE9ZuzhXO3fkC8dMfIedIE2T+MzeSSOrA3jadZdnDezfd+cM4hl4qyCpS
jrS9/hMeguMzNX+5jbpAq9uNb5f0SJcSN0RVO0bnu3UfusWhbpdbGHaj+bvyDUav
MwgW4XQFU1QnTPcU1PvppcuGtsdn51eVEicj2bF+sT8iCqbT112bCForfF4wgQmM
ifVIYuHyezfRElUmfpHmK8DpkNPXhY56EsQEdhOyRftgdzBZuVOxa9XcizVBpZbq
hNUIOd6hpk4plHYN+4PPsAnUpFjAY9kmdu1kpL3m2gMSGeLs8/nsuW9d6h66ee5n
HwnoG09Ho+oDY7OH3WkTJrcbA4aidBKtk6nTaeuraSCm5Dz24UahzYE2cubB252w
1OVAaoFJ/Qswy1tzCgYCIilxlp/xp/tdQzpEsDrVAMg=
`protect END_PROTECTED
