`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eyeyP+lcPzSkPGUvakBSFp8rG+DTeCPlRiehOeT19s/D6HxZvUa7eTWpQyItlzf6
YjUFAHfFS1W3Hg2mdwoXBRaK6xIg+IAOiaeNX3NfXU/9km14wkHq8Bba7Fr8dlfG
NShUlZ1hdxCELNgA/PAKG4cgixQg5VsK9JQWJgGFNupboACqdOgfWBbko+BGSRzY
++msphXEEF1pmtuf/0GNn/t+CzRr4E3Cw2Pu4fNq/opGGagUBk2lP+iXwYDALRbg
EU9OmKSEe0BAG0PbyWK9IOzYkHEa4EXDQxQesUPCX3vP61IDcH590WnetxFHNgbY
jPDzSKPdyPgHjlDLlZBEnWPq0TLmXVb94IL3W9OMreCS2pzCO7bxdcSmiSoHtb7k
ONthyAbl6axxScBESPwe4gkJayM7iC2cxn1e+9PucqnpH0XzUSSOVms52k9ZLELs
xK6X2kcVieNmeJx/PzsmrW1K0WRStj3dPpPzBX83IzfcDoHk9/MiEFtCHZTFeq+R
b/uXf0DFmaCX2N3VX7kKpOBCIvp4GzOb8T1O/SZ/aGbWnEKSIGVezPiTLe10XJga
idHsG62K8dpYaSixcLkExgFM6om0K/2e0oa9UAjcn4xkFG7/NgFIfbdgp29gmBJC
+OpjXVQHufWSjfvQu7M31uFowOf0fpsnFVXv95hQSiIzkb76EBhzDjpvfIaQSqFZ
4XeUASpny0FWqaaacZnA/ByY59as6FgbvJmvTAPm1v5iCxaS8MEsLhQ5P28p9Ygr
iQ69Wzq3ajoQRV5yfn7z2kuFX+qMGmY+xZqnAygTE8NnNsP7a8sZF7a0Cq0DNpgT
ZX7QPIJ0ZJYSiaNq1Lp5/3++cGhaSRWBgMLx1YGVDSASa9fBmFXX/ThmdQsOUeg1
X6vhTiAkq8iEgwgShpyyCq7Pp9x/zzruYQVhSNHtdSeW8mOJRu3SBF2pq0unwEKw
e/qYlxxJDymvLwRrHuZRpQ==
`protect END_PROTECTED
