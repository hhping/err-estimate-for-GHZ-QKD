`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtxQAk6lzC9gaczZ2/3XZOo1o8LUCjFJz59Prq4qk3hn1KEwIDAYH8AhxltJ7mVW
DkEJZneTsiE1QKB1/Zl6pZSWYFlydmmwP2BRcGoaFeLpHSRkCqEZUdTorsGwXrMj
NjuW9ubYX2My8Vq9OLbKd2cGj5VNUirUfvxJCWLcxLJZWBMoo5Yno4c1x3Y1TSEr
MCqaAqYUhC3Zgz0HN0gMct7JMq6UXIez3ebybEebme0xD1i0zzA8AjMa8gM2e+6s
JUXMNE8CM4zDIRicJI0BTnMDoxWnL8pFSKsUDjc/y7cd/jTTHuz0iHyxvISBJJwr
HbUYArls3NJtuDMH8Fyr5vexl25T8Khv5++p7IFK5BU2Ysevhix0u9pS7P6Vn4XM
CVc3sBnZaAo1QLo+30JJx1a6ivfaeWZuS6KDrF4IzNZwNqskFX7G1bHm5arXhtW9
EEVhSMxK6reBrCthleLoiV0A0lqn/gWFhInUVzmbZY+LPgv7+BvIgUSJeCTxYAzr
uayDAUu7cETBzJKRxPebp3M29noQgyj9qJpzJ05OOAONUzNBeMwfQOo2FgMsjSJz
2ZLy73MD7q+osvVHu84MmNYL2pVtKtOjebMnd7WjjvJh+jnmwxyhnXW1JHNnxx6p
gayd6UsJww9ZsM77Z8RSmbIy3OGv92vNw9KuYrlqeqYwUXiXjW4oULTObnLth+f8
yvLwkyv2HK5lS70FSizsZjPsGHUXcQW3vGTsmzWQuPeggdMW5ldbPgNwoBKPCKXj
o8343B8Qh3Yx9WocbEFckndsD4BruIdP5WXFQtjQ215mDgWsQahG/N5J2RfAGQe2
UY/QRP8sxqKSWmf7suRgU1FvsBdMzr4tt3gru2G+jJf+p9PuwCs2CD+fEiJRwUNd
6W7jR83kWFsBdkWVO3Z95oPXJhcY7VnErkFG710QnZuPEi0nS6JZKie75zakUq5s
inyiwNC6+xK++aJUVXcbugyOrxUyodnNll/PLIQtm8dNdzRT1bbkzi6+gafi8Llk
V8/uVUgSja+z4/mgX6HSB3iG8Zqz8f9wjp7dnvRpl3uMKYsz/YjR+IoPgRCbh+I5
r0Mjrqs19YS6VrkNlIelEYg0k9LEWUOhZlbxbyqJtWkJ466n62a50tvP6GDOXtAb
gUASuMEVX5ISLlTzmhDTqCAPHm0M6BUpewEKVZiqWmFIdUHIzyOxR8Yh3FVfVBfo
zyiQJczshkm8LRthkSZFg0BtNETb2Ih66m1827bJrwJiZ5A410kvytna6kSL/3OS
PYdnU9QZdwhywkfAWWFzewSU7AoBelpGjb5mRsq5k34yg6dX79ZXdBhDdeOxsVsn
jftXvHC5oBPo4ESkLQIc6D8YIgdAY7t8z5mZEiqBSdVoIP9Sj3GfPFZnIAc4D5BH
J9+KudgEoSxwDOKXSQqvqNjrj0loEL28W9ywGhFpNDvWwG4JabxkULlve/1L8qOd
IdrWRZNFiSVpMi4Lpzk9Kk2se3piGUY01U7cqFi4+lMlIyRaNS4gDAk0h8N5vDtQ
DPmv9d/BQG17amwkvZA9QdDRz226G0iLJNMnChsHR3SeAvZdTDNMVOOJwr2Jv2ka
udqgXAAZHQyap7DA8Vav5j/v+sw6qgRFSxhSeZidzHa2pWzwWkSL8ek0LXu/BnJ5
OJqxdyBY+0rpCf3eVQGwnc7/Y892ogU0cjqCfrYsld335LdR/6lLVOJyzdTJalB6
GBkHZsrZgxYGWDfH1dWIK41RuB6Mba4YvrKZYm5vXtiltwCDVJbXHrss5sopqXSf
qsRq8Piqh0NVcLMCXrMMVVP8vqq1fnhfgNN2FjdhaHNP9bNM09xVJLSA5aSPW5e7
Mlu9alyG55cxZBzpcr3LldlOIHHgJc2xIBlo/fEqhNy57BVG8AsfRm1z02nI6xUJ
Lfm+qJhMFiEl6ylBDVpjPDXlO7LgoWtprDOE9D5mzU/K/kCPLw2fAxZ0fP0jhs2b
gyxhCtTcVTNWiJXOVMUv1Tgg3m+HJo8UBG0xHqZ/V2QIoRUv47eHjPgwTJTbbzd4
/6zxLadTyoLYNDXqlJEBoc5uXkTGJqSpfpQMf4xHD8NjaOACysGgSIE4t+F1RS07
d+99AUrR+udfXnEqE0mkjq+iENKisssSJvEmPnKy/r4SSnquNHWaQrq0bmXNZuW3
i2nZU4EQRoeJpmdwTCUO1RFhbrL8beSOwSnjvhdEVgYY0vCq9MPvoNWI0tfPRuOw
606GdK3uj0tVVbh7/0yAs25YsORCcgnc4758pX7GwoV/wRXYtkARL6rvMiPdtAhF
+9sI8F+rLtq/42/KZgW75NfsjjiGlO8DlWbeJwBGmkUeKhMwxS4fYSWuQgR4sN7L
9lMbbi6EPwOqwibnpV5S0qzMwHMjMWS1qb7bxlHVufVTlgBWBObBpefQ5YRR3mO6
CtJ9AHaJ7jKmk+MUcT/bcPd/DNwNbP9op75MHiG6j2PYjP7iR/DVZJCpp5eeG3m2
lWjUY+qJezeV90ZlSiqx2sxjromMkTxLo3ADNi9PN/mvQ2ilxA9npjBot2a9iwxe
DOZak5+XEQdoHTBtQxGLQT6gPXWW2h9otl+bX4bvmObNo0K03/L/qUQMnxjHe+7v
nw1OI/GIkR9ark260+I1kwIxMGDgO7RAnDGhuyYxnledwTCfE5kwQ1ovczQYVSRR
ATMBs6YIyEnYPmcdU/CvdBbCYS6SWdFWYQaVdRkvhVmkY7nXOniIklrrk9nfeVCp
urmUpc0Pj+nkTp91tlMJSSsSEQ/y2qubx6QxhCQRdME8zZsXAdAiISw8ZVKxSNXB
a79L9jO5FqgXgTIbxnTvEy2L6lxLs3ewMVZSRazzM6UODCpnuTkCARrA00Ijfzk+
uPn24YMS11p5hF7DEUQkYs1WAK5k20qp4Vl1YpPH70PMiJl7mWlZ0qZCRfSHfNjf
ooLkMsIsE+9mzVmuzQwWvSacg45KNAxibN5+T7wM48bII7Hny3vhpIrwnLU8cM0B
4Na2FpGAVDLVdgwSnUYJgnisRESVLSS89gq6hPdjFtp4wMM4LM+0fRznLsgAeBfx
SM88TJ5BVsN+SWIcGbnyckxMrwlN+mrO5q24GHnFdOo=
`protect END_PROTECTED
