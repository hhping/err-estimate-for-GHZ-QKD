`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwapfvOTeuoIcwO+29PQanVNH0BPL/IM41c1F2dTTjz20G2FmkE2xzQXGE93FKic
J6dY0XKKsCBFXoCF9qnupg1eBTc8FTUt3bqjqeg1DTNCP1A5rz0AbDg+Zspt6dTi
YVw1nWj6OazvXA0YThdl+OFbctBGb5NwlszuA75L3uNdUmNcI5wNg/McKvVczUjY
r6DSVZlquj/sdwqWPRKe0oMpehtq/iyapiylzuqysgxhz9yFKa583I2bG/Ihonz3
OR8XSAlk/eZhMi1zY13YhNcmEyOUK1Rlkxf01wWOlMQo2Ee30ei4y54JdTW7K6Sm
WVNux7r8kDUSkIBbP1u/U8wFP3iDTS1CpWuQyOH9wxRw992CI2bovErOaPJtvau0
NiDuNm8MOa8sXGK53N8qa9TdPScBFs6CkP2f4yji5stdHHldIzWt8k3pnZVHXHn1
P52Y+urcu1xqmpWa0O7tDCG5kFBkxCoR7bq3KO/UyoP2q2OCuZHckQE+5woVYV9W
GPqO26V1WB0nb280yCOzOWq8KIjrwjSaETdUE2VFKG98w1oSsi1qtMb6lbR0xpCV
pbPGb23k9+dVutkJTRH4jVjF2QHmFV53xA0hoCC6lvc+1zPgR7mXhdvM2e+HDjmO
3RCtLbnVzS/QDiPUsjXYOPrUmvUXofwp9p7G4qUN3AvwYr46Wvw903RUfDP7w2cU
Yrnu1gk5bwIDTyBOD9x8A/+iSdOg23KzlvpFr9A3ErQ+ZRSI4Qd4Pd9PIa3D3qZF
tB1NxdYhoSlXMilWJ0qCvIGmz4GsS4RKs7DPCgUlG696KT7G3/gp4uPLcEvyLdg7
X/CXuvtBZLbc2sD595l7/gLva/vDdCy4dbMHYIFrpIqrIxP+UHEeZq7ImDNv7sxn
lKWXGRvVIyrWIEnnTunr6E5QhxnMh8mdg1WkKTICBC6h5YmL/ftX6TRQSD/G0YTV
L3HO4qbOSEkW4+p5/ox/GCY0802aQYV2Aj7uBH0ozmNAACx4mEsf7pNFjFpONomE
Tm0rWmpua/2Op3/lSV0YBsomg8gTsZn1U6jtkYThVrA5fWz+q6dN7w47sbGwp1D3
qCjldUEtzaounYaPX2zqA/3GyjBlybbVIDoZY19OPuM9UDnsGGsZzKOAJScxqBD9
W9fCwV9c+Zg8Y4pbxCJtpw8YLc+bfxJMCWxMS6x3CBaadg9i1+fWeTmyt2d3Hkji
9QqbhcWCCHjYy+5rU5wlej83z+H6YpROPurmUrdnbS+OcbRwrpfw0L4Ds0uNw3j3
Ym0ceqWY4BfQfGWmuyMUhMrAtoqyTn7VoxLmOasMRg/UA+lmPZ+YbxeFfTCW6Z7v
yJ/uHnI7W8zsLINWokCNdkwKq7Og9fJ3XcLBp9uDvWa8EZFLwZhISiWGyRhN/T5/
yY6BSYuZTYbORCtMNjvc7rwQjmKgupm+S7lYo52GOahGLd9WbIgb6ziQNoAmtRiC
15xobYUA54Yw7rnPImLV6if+FV6lBrDwkiqZOjl30+4a/ZSzkvbgxVZlHbUnAXzj
lWWT40Qr7WRzGb6OPVMLkhRHYmjP/8rVe2FvCR2fjdagZ6jSclyME6hpcXCkvBfL
xf+1oW1VysLdK7wjJYt4Ib0yl6NqWhJ0EzxJU1ih5BJ6Bl5vyF/X3S3t3xgNqKbu
X0TCa5MilhvVERo6pIzUPGScXUyYP7ZTUlS8flgkJ1LjnHcrXY22HAutVjxgyy6g
XKNOFD7uEAJbVucLpGlluCqDPCEuyVVOeeTJGlTPbuSvYFoC926S5jfug0bkLc25
s/EpLYBSN0csyhLAddpd3mzjkB9UWzJ/sCBLqzlcKanO2HhR+pbpZ4AQogObwNoO
`protect END_PROTECTED
