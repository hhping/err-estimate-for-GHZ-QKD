`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egehF5/BFsm8w6Bm5OS40Lc8acoyuWy8ZpQOVseRmWTk9Z+PwG7/EIdVj+fvEAIS
e6aaeYhp5ZRwVIiJPP3/D1QhzwNt2q7AcrS645pp7DB9dAoHlWqKMZheJNnru/6O
e0yH/z/xwNQBBB5YYxRWqHm7c5UdQfVxjaapjKHiwHHJV2MzKQBsViXtTaQ+ExFs
+Kc3ZK0vgxaPNWGx4DQCY8fPX0hL0ogCq5e+l+Dp+Saels57BmzfpojOD+RIZT9O
aMrw2rxjJJ9yXoFIUS9PZrMo4WgROna91gmJaZ2d7kVJx2bFBtLst+LRRPeVH1ky
l6BaPVhvJMz1XRhiq1k31Pmy3V7qDuSWNbyWyv2/NyeMPnwTvWGZFK7wkLCpghUB
3ECZZqDXBBY8gNHkjoUD7SLqLAO+Qt7vALiSU/bAUPdBANBlCo5+RLp03G6z+dkE
sW3v0ODl1dJRrkignOETEKKumk9iekRAEKhOorCX2lmbKRXGsUHuvkVNXKSN1m1c
`protect END_PROTECTED
