`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uSvKY+6QGu58zJ78REdFcm9vhZqAgR9iU3DDvn26pvz2RK8VAmOAuTsQZloyQnL
JopRW7xHgomX2K6Fn0Y+EBK80iRVxhi42nVTlSR57NOte6lSiB2vl6W5YafxVOzS
LTgSCJHboIkaVffhAs2nHHmco1rfWHZH3BMD/I+xGu1CecgCh/BJxrOkUdNMsrY/
zY4fvTgus7M9mVYOsA3+JLR7EFlua+fr89f7vN9XzTFX7f/3N2blQkZTilhHCv5S
2AJaq1DF4OWKs6rYa6cvjPWnIwl11f3fDC8IKFSefoUU+J7X8vqdwsyfsSOC5G4U
rb21EGre2Kb0dLT79hh5HJxgipXKE5m7d3IgfWysOO3QZTBOS7+SgMmiqo7+AwRv
HX/h2haTZyWGBWM4mR5J5+bdfpXU2GX5dWyg2anuRtRyDA5WlJJ8XUBnZzQ/ncRX
Xwgkd3/wiTYsedC4E7cg8BWjzL1+ahUGI3CCh74A5MuXxsdYmVDpd0ZM2Qk2pdSu
oJIKtiFL//v1KMedNCqW+nPJMbQOjF9tHQRm4xCRy2g=
`protect END_PROTECTED
