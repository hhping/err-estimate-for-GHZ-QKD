`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQFpy2bHbL+pHfroIB9E0T+RcHDCzMkxaqz+oKUEDDL26RmnMzmUXFIAIBNcAwPI
Ci5jc2z9XYV29hDRWhaMMxcs5LhpcsGl2wCg3adqDMVe7uQcCyoYAwj32K5R7C17
dUOmmlqxjuGlmKJr095X7Hf6KxHfRUKDtlKB810GwuJK2/NO67cwOgIsO95ZLNBP
hEeMmZeh0Vh9Wz+zmOeZ0SUxwJrE+1RRY/gAQJK126FN+D35A3nCbfM4B0is4yAg
d+PEGa7AD6a8muDA9nX4s7FgeudBYspgIcWDBcc83Cc1/2WUQFkCmhsPPYKf8zhg
IsRCls93UkEn4n7D/MuSDw1JrdvFU+B8yXwntjAtVtPRsIC7IYut8mFp2cPowpwD
RJuhyaXYFORFOt7Pt4TogRMLKz4CmxyITLaToTdTPVYnsE5aCvY3pfoHiD18geWH
a648NYYDrICGn/nUBMr1Aqv3zryJu8pyrEGvoyk4WjIhlgcpnOG2ZiBL9T88q8z5
vUPacdkuxPreS4npYIgNVoSnCnavIMTlGbWCxu1C9sIeDP89kIgnxSHeZ4xg81/2
s8jwB2QyTHR2sdcYpJqlqw1QTK78XsciwgOJ82ks+T2kHB1LuCW8e+EmB4eJmCGD
mQi+CSQ61/BH41cPwZMIck0BTj4Ll8L0zZQV89gMDL9sYtdgWEv8Gx31QAtrl7F0
KRrYr1y9eNUpYACBJLH4pQ==
`protect END_PROTECTED
