`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J59mttgmtPX+bM0kQVXWj1EjVvuuvIZ7lTIqGxjkKyA1tAyQXnashD+A8tmu9mL8
JYFpUFwpsxwk44ZJiwsWk7OgdV+DQrgdtNRy+9QXXFlSio/DSpP9YHMLtTiUnITq
OHmj9q2YIindXKfxUs6q7gdcH+WIfhRlIyICO/C3nS6GumQWIMz8Okw5pgoOFg4I
qbkZbyCL3DtvatDZJrM/g6MXwosPwSACUwmnYiC+HVSgrKTkTiAA/oyA0wDxoEhD
u5QwlAuUiUkUSkPMaB0p8pY6LSpS2OUOLlzeG9cxCRKKirk0TTNbVvPuMCnW/95A
Toy7GBuJFGT5JquQxdaYpTNE5KU+Y1ufYRGjtVYZPLIbAhOPT7UO+vPyHV8W9l60
eRV9hvcFTvgJNtqyXtbd3xwMJjoNeEKSJFXk8Gl9xphbKdNLdniAnPY5T0P0rJPj
XdOCPErmRaYLhDIj6DjI2wXOUoYVcXZBDXWs9M4723dN08ZQU/8QGMtt115wR7hR
O3uXnn+vaT5uodDWqSgKQHiyb9W/I4+a33XFNIMisCR0R3e9kmWGhMbCz3tIdvZg
/u+S8gF02pqafCCoA4i8og54taMVgoGgVgtxx9JZr3Ht6AonG7uAdQtpemw8/km0
lXUzaiY7fSilOlUgLXD+wc7nR5w9Q28CYcJDR0Lew+4znmhfZ8Cvlk91kIpP24Tq
sqPfOtH0EFPuUlEZlXnpuA3IvnGxahSXrtMnMed/nYWYwAHGlejw8dMfx8B3PTY1
M3tdAzKxtI6oNAW+GHA6mNxrCvXVN5GMdDFnL/Ff3KUFYMemw+ifI4J/FJXmiSsm
2AzG0WcIOLgliN0X95YCKPok2IUCzJ4FhllBF/IBQ16C8O9GnvOazJMDz12LstmK
Ru1SLZ76SH6n6ESPf4i24Apr3MMFxyqr+TueN2L196mUQ+dqgkXKPAGsv7WMFVnp
IER+t7K8EDBnJKbkGrShZNlRmkZIbnU9xDjN6REEDd0xSivxh7RywTFrTEsqOwI/
ZQrKarQQGKfhHjb5CVvowbAA1kzW6vzn9cUNKOmp744aqslFaG58RU7ftaRYJQX1
fKmBRjBrSO0k0dGpAqJ5nKOU/XZ27yPA+7C1D/c0t4cNi6DXvuFmZwOtWEZSRl9c
rC2TDZ/Ud0+Bu8xu09RV+SQ2aejKepg23+lCTwCIZG4K8PBeK2t4708JnAOMfOJj
HASW17pexaDYVk9wksXXmOhumEswe+kVch9m9udP5f159w4Wpn+buNYZSDuh4E5B
zsCVJklp0APqfaNWZz4ZSnyRK+zSss4gZkepmQQSB8B7G/suXvi2b3NJhSgmJhqE
ag9tEom3Ev4o7odHwEtpPA==
`protect END_PROTECTED
