`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9oYQnjPxgI9ojrsL6gBncWy1b9oHs3OJub8+MVO0sR1R11tOkRniUqDX9kFQpqjK
GNIyiXNcmYr9SGZWloYUeN09WlwVudEpWdF3+Htx5hrU2HfAjrcJzBvD4YVB+bz0
fvXwiyI0esQ3Mk05xXqx/28SFaABLOd+mOk8BWIfWwVQsugDsr8UeonxoYWibi+Y
MCON4z3lO8Qt7ilaffzU9fQHixkBqlhnXQS3Riyq6cNxk89EAF2ai4dhMP1L7mv+
6Dn2xAxzH4yBDNt5cRUPZ61t58/It4RxTmh0sK30vbkGRbzHdrcXDly15jRexx93
Smf8E8v9LTrBRaH9ay/GWY0CJtwMsuV8fZndCLnIcyeqPPguDBZOLZP4g8BaXgwm
03J15DUIG9TiUGy0jMgtjIocZnCNrGO+0HVBB7vcr2b1tyIN1owgRFVibTdsUAhY
Nw+vmJ/C011hhYUJtJtFSFZab+UEK1LuNkKtXlod0jCnO8c1nCx/ODL6fnjovbPG
SfBwi3x/uJ9bxckGrZE3grmc98w9KsFpam6mVcb3EosdV47MiwYk9Pv0/ezBSdQt
VKQqNgMPpDBiZDHx9Z93T6AiujQnRhyCTEdimGUdxqPz/1nEGrKafxsPVx2B0q2O
+AcSDwxyV5npqRGdg0YhPNKhnh1qxsZb91dg5oHEzi66TAPs8ySo4bzDAHuPKYaV
61b9JWhAdk+W8LXNnBMnAj3mW3NgDG3zV1RIhDAa2sM=
`protect END_PROTECTED
