`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xd9NKDcG7N7fTuzF2TsNBXaT4R7BGha4yQBgiag0uVLLZcFRAcXo9oRKKlXUMQxM
uhaUFWD76+nI4jtMjqa6znwFNNb5a07coqTzNPPSnmkbN1/PilS6moAiTx0B2Ghh
mFoVk/quOJVMbScaOtgoMIYmYGensMSjSilIGKlnpQS62Rh667CXKy72Pz8r+Hr2
Y9raY4iBTuos8mMKOO0J7gEl1w92jWH8wjz70I9fLRnwm990gTU/Fxsr+tO/sQ9+
jFKYjgztbJBgeEoFaRzPwOSzQaXiplNDVurwt7V8yl9BqiPMAp/8Bep0EbCIoXu7
XhZoFzdMun38UAKsbHv6jznKgXLwdetNPGXzZJEJ4HPoSCakPvM169pwkn9KsMGI
yoLGBu9PtCtEJQ+fzjsb9jlyd/JTQhdWqjoVjW9wXClTww2XEvRNSaDRIlkK8WB/
wHXIpSTcxIzv1bQn58Wlig==
`protect END_PROTECTED
