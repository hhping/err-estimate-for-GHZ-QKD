`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SM14hDCChzXTjRBD0gAJSXDJ2zlXPMR2zaBC9Yq//IN/qX1GKOms9gqd/LjSM45s
vg1yLg8WWeVM/xt59MPblvn9uEVLQkbwdThANcDqdybvFiCDzX0iWTDwmCDtTc3J
6BI41QDav8RhoBPlk/QOdFTOoL1i1oDpyQLyHu9TpMPQOJ3yf5c9V5+b8/t2USJ4
eJrDskuu/ZSmAc5AUzHXc++39TOEVX4A16KCGZEuH99gnizJc2zlD4t5ohhQwDA8
YtJCg3Yl+Y0RC+nM+lBS90KpDRlknRHXulIyjVp1SccpzhKZPTE1jPy3GM6Bu9ls
9vqhQycHPDvU/5Y00FI3c/XbZc2VJ15Z/QLLwT3rD4M8MR4iZAJGytuCOIkyQ3Um
WldSaZmZYER5cdWWnp48DLYLQwq0neJTD+MIYMCk+JaUUtMOAdsQiSk4E33h3JaH
fV3GWhEaNZKOfLYkG8DM/Ic5iNQHbAaBXMJOEQHgUXWz5wSczZyZLCbKER37LIdt
Cu3z1nPRyaYXFCqt6MvYCTqs2wWjzNVZyoWK/VsAnvjMiBRWRw2v2JlVQwtjFnY5
zoY2mzjVLkIYoPLUmj/O/fPkdfKdpU/AlCiw7QjYzcwpDWDshTzCKFeDQaEN+yhy
jZfmPRBIbpRH6pfe0/x6c8evuUiQtmzojF2eBuZ8QqAuKmYElFzt0ql2J1YUoDeO
UH+fjedmSgp2/vrLH69x601nhP+C+Kqxer3HNeTNGI/6RyikmuEozfbUynsX6UWP
enMWNiDFmLLKJHrwMvzw0uTk948+OKRcqDZYGWSggsC1/r4hYJKFdxHO4OMzORkl
iyHPQWMq5pVk3o+S5ei5xCEov1KMr4YTu3vRdaephbm5Kg3zaQwYov/knxiP7VU/
qDsUeO1rDXe/kRefaCODpzu+bTbn2cwyK1pOKmY2gvsQ2sDmXiGQ+toOdnf+zIeG
Xr+zbaAQ6ISUn2Sft87AaJtW9Ndd4DgXxDeFOmBykYdzlypKR5fd35NG2aqNY3sm
o++gl3/ZUjmn5wZMB9Jskry2EDJfzC2vZnb005ydPB1fsFfQSMT+JPysjctvhUTq
IleNAIB7CUXUiKg/qqXIEUuJRuWfuOazXLFRgCU/A7zEmTca7XssjpgniDlXz7w5
DiVuZm+ZOUOu4xxPSQsGPv0r1XVomEJ39cSQDK86to4r6+Ldba19TUGw3jSE/3PK
69F7Ex0A+dtGTsVPeZJ2CZRLkE4RO5lIibikZlyFoaUYq+QDkE6+yFKHNb2tUhDQ
fj9B75mn6LHJUEYCzlV7c8eJJuWwQkCOX3xMxqcHXKXqwojrU/pMzq+yaaFK1g9+
dUmEjMUDEhwb3BBMeXuK+qtlx9xL8tL1ybmKh8TZ3YayR+IEKGHmGT68BNOpfLJ9
LX8Dc0wMKSA56Nvm35MBMeV/lRgvt67EL+ZNQ1K0vFCZjT1c0XqJMTgXBrGz+vwu
ukf6tAn7cdvbLe44Th3olD0nX3WovdONtv0Q6c9yBWWKXrQrAmRbfkhaeXZ0dQzL
mVF29Zz5QJeIsmmnZHtgBoAIPnZshrMGan3MB9WBQs+1z6C11q92fmtw757EagE0
ES7dDFWcdNkvwC/t+N9zynpfDuCp6uR2oEqTxAj89dnIWz3cceGo0O0TqNlM32EK
VfuuL/hx15yV6pINHasFa6DAy0pSqx6d+yestR/1SperYeVp+0poshV+zROaZ3Pk
8H8m9lxlrDNrlvhtrGeSacewSxxCwSR3ZsAAc9T+oj8bEDnyiTzLUb8lhmtVleiq
9nWzSRwJA9vGNhuE66wRui6PF+sumu6QZIqbKTb9tJ0DwdpeRsQklQrXNSj6lQ76
cR9Bb/8sUvIMiCFgXpBMVZ7qhBReyi6YzGsgvGP3BiixlQ4sMEjHa+VS1eGbHOKM
a99I3ohWWRUjbw9VerZJTC6effj6GHyncSs/KBUCm08=
`protect END_PROTECTED
