`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7FYtaIx/nl29H0vPEeDUjFV8pQZgtkwrWkrBCdmAkxHE04BtCT1SNfexiPP8BYx
06r/DMUlaNj9uZgcbWIHQVphuWWAsSCp57l4xILb5oPSjy5p4Y5uAC7M7t5vpPlI
VhY9ojYZ4YnkNOSFTLvCy2zNvz01i7d6w2Qd5x90Zo1bja/hRIejPVAabYCRoxH4
pij8lkAleAxCdHp21v1zxGxg3t8KhZpYUVCOzkfzvUyaOeGIP/wA37xC2D1gd+Wj
P5D3TEXXLY/rv7iq565riSgDGs5iuG+ijZRcnBg4bDCoVZn5JBG57erWkwCOh86/
VIRyP2OkTiv/zC7SGRjwc+M2sjbgrD/pfOHnsywgrOiOhPjWbW4TEFjEQOeEP/UW
upMJPPE7PnC5mwgKP2sPZzeIJlVFJabmDad7lp/rp7hD2whVeunNO9nrvUcLs6TP
9dtkSxkFVe2bmML1Rv3BgN5ITWP4dalYZrurGVyOeiijCQ9d5yoTw1Qkvwsqloz/
h1cFaBcCMATiR4R0BswaOXNiAbC27Rmgu9Twpx3jFlRzrns13g6aAppeRyFCdrL3
SDRxapv4GnJ70xzZh6dS6GAIdl1DH1lM/f3ggsgVbcW2vwnkW6kKqfgxpj5o9Ren
`protect END_PROTECTED
