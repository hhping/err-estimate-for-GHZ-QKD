`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ib6/yduh10hl6qj6sJOKYvdQin1MMJiYVt86k3cVhIImXuxI6dHAzw7HHWPUS5ed
ZZG9eZ61BaGlrw7p4Sx0vqkhL0J2kafjNXKk0nHsIi8N3zZ4euGLWq//jYr8ovc0
l3wGyxcGV+c5rPglpTxvJdJ+toO9jP6G/68lGSjBbpHFlhwSbp8Rsb9TnZC1xbh5
E34VUz5Z+qSV1yuog7YRq2jOyUO/lQsNg2muaZ8czX6Yrkim7YseKvQmch6RJfiK
kaHkfSsZf6vMUsOcVWenXDZ/RfWH1hjk8c2wiLWM4/bYtKWnNrehcDAwlGiIJOv3
ZDjdOhhdYlDWRN6vPJIcrVC0AkcDyA3DQbVKsYRoVBp9Q5B3tlEEzONqxCh/MBKl
xGOlpTFvpZpXq8wS5d7zZuV1L2jSzoBa3TNYmTscrGByh/szey3GBq9Jz6zeWiv6
eYTgA/UtTXIT+NRaIWbuzsS5W7HsYpCjOdccoKmtePwf78d3H/SPlwYvKURdWNQa
bPZZxcw37HNPtxW2V4lRCOsK2qewD0zvkuBETqDCtzf8s+/f2R/FSTrRyUbl9tM9
+Hum4uvC60UXu5oxFdwC6qsgxv64tSNSjE/rQE5DTyUBa76wqcVk8WHMUcvhgZ9D
zr+7H2Q12/k5L8+xOADvkNH2YGTA7eh6NazvzXlnCBNEhbOyqaIUhN6otkiyjjtu
3zY12lXz8VgnWD4pM3s1WFkv75/SYhho2e3uzdbwBQOBX6VLtfxIKOM50DH4o/4C
gnhck+k7wSCaQwmLhl36e4Euznu1jxgUDzwC5fcHjG24ANztRkLBQ9cpc3PSYnS2
At2D8nBr+v4ngAfWhzxV5Q0nAwU5mzXl6tLTh0rZXeqZzehAcf3rLX1Y4rkd09tv
hBhX/qja9RgFBSmAb4Bvo77j1P7d3nSZjmjo2UBrbFYGim+fEwTbs+rUpScI38++
y1yy5Nee5kCqmt6+K5RbWw7ZxVv9i8K/eZ/9nrOe0hfsHGF60ukvqCjCmwcMHqfi
P3LRMvjadrBjMtfKdPYHz46H3VIpgMmfxWnt625iGSeFItXyI+s5/ED11qLYV2JK
nZtxXLgHHwjdjp8el3U/KzOiPCY6acmNQxRbsv7zQY5HqRcX/wgHst2ByN3HAOs8
vpU73M6wIKAR72kKyq4lMUuMhkzs1nK990oRBgtzrUM930RxTZls9fVObUiMPQ4t
NfPEb7Uin5cKOpOcG94cA4cFn9nncGeol+5pj/xU5GG9/X0scIMozdM3TIEwAjd3
YXbVLqO6fxGMJD4gNLdDNaAZDuCWqUp8KlJkCQYqpIAyGBqoeS3rFxk6/qsSbGWQ
wqd4vrCR55YecwpvHJ0ZoWB+/dPMNOre/ZkCSBrAohzQreX5JhuTi4g8B7Yy/UwG
1wbxVHC+ze6X3C8HDc5mkl8gPexB+PLNo03D5yaEFE3H9JbogGNDlGu2ljsOCRqc
nEZxaidhVGnakR7fuQkMWTFJO+Veglvz9h6m43mEeOzdtRCrqzlTYAibEA47oCTX
NI9wR/a+ie5GEhyIery4E/I2Dqo619tYU++DGC1AX/MMWZHV9zOn5cXEnG3e9Wwq
1NxmctLJZySPgcFmgtv5MrHogAU7VlgA7utMFJ0b7SRuSIBedIkNUCwERFtqu9Sm
ma/5j76eecjCfg3Tbl6wxQ==
`protect END_PROTECTED
