`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvHRwCZNIARjPuwsYjW/9O+y0JT5m98nroadqR0LloHKTUA2bSRBNwegA6BJaw0X
DiQY2qIxqeBNVOEYPrer26ymbbSlIXlPmc+yafvOMplUkNsgvS92GY0LVvNeExKc
+92oLRrSvvq2NTE98ijkda7E2NQQ0EaxUsK3iJ/sHUpnVJt83NqcvtTZYCL/RWzt
VPoekFIFISgEkrVj76Fobixnzmrb3g8bYRxz7Iz4ggdehHIAWo5SVWxCv9ssoTpR
9FgYeNDy3OfHk0l4luX0x/Wr/eRy9wVfzeB11pFTD9aTkh7P01Ap2n4gH/QonnTb
PKC1AKz6M1GRAeTZtZ7c7U+jcsp+6OcJ1+IWXEAAhpF0FOx226Nbw9G6AXdFuw8U
ASUmVvyI5ht6RZKcv2y/eV03lktWfkmY4wOeUM8Td0TO0nvekjquAT7Xr15Y1w9s
6mZ3WJ0sYzXBP42zGf4IurJXBZP6+uRG+hEpjRSOH1J+h95JD0AwwzyndUD13Abx
971xhkHU2aaARxJy+kGy0LU6mOAKz+6TwjbqxM16Ad5Kd5FwF4znjdGlY+tro9Jo
VjIOC1lg9Vedx6+xev/ItP3GH3kYAfSvcH38RMO9Y3fvP8IVM1RWBTBt+CLb/pJ+
+eAaAAZnFohF5wyjsxcgVlELRz1zhDULXdKwsBZ0LRK8arPKSki41FFQIKzcx//6
4EPwUOb5KQwTek6YWS8VO1xt78/5Y8f/OfAEPenmcPePc+6O5inT5LW31AOGxGt3
Z+aEnxtGVSt/UV+ykij36Q==
`protect END_PROTECTED
