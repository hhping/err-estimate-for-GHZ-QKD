`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KP/k+2E/Lu2PuPoSCYX394QikC3gF9AFmXDlOvOtaZ3+R9Qiy2hscXh0OuKQPhuW
yo4e6oxtUMWlbMDzZKBojHE2Gs6gMisf+d3wZMr/o1oL7Zke/aeqSQ8HvXmsrMDo
kliasmQpafEoBAB002QaSczzEP6VyuIKyr1pGmPEaaTdclJhQ80NGl+Zubzj7agk
S/wUz2gc3Me7eRKstLlBVtl3mSBf338FNOBfkTutvVF20GiCeYoSXdOLd5jtGSPv
AQGWmhmgyNuRZ9Zn1sMdBt3tPHXbMKLZlfRnsS6OwQ0aitbRDRhODE+sEAvIzdNz
ZHp3s5UQkrqBwZgTRtU/XdpMW3My4H4XasuJ7+83cOJZIlvCygnn/vhLZaKE+YTW
QHK6tSq3i8KwOYgUPtTKCfdsruHe3euj7vUetWS5IlBG6Hq65SjTndKGjp0ARX6/
y2aI0H2Cph5eGeNHZ/olLGqh5tu1moqlUb6PSzTHfkqAAEqm3nglWlTihKDhYQuF
JvkLjGhdV7KyvENr+Z23qRhZb/b3v4TfepmH6PVYR9AfEk7BBGzXflEKcIacJ8Ry
XcxCYbugEpi7qb+YRx4hepBt3DQ5Z6k3VpkMOH1qvUNXXhlSdr3PoatqwZ4B0HHK
jvJ2j+D/F4Y7oIXmp7b3C/BiwodIvYTIxYyhvcFLDbZquhZus5cnk1/AWmgtV5Ek
nSZnMJxDTkQVTAr2B09q3eL9Tt6qlgEM6PvyBhTBT1PmBHo/ZhxBKu3OTdaapGOG
`protect END_PROTECTED
