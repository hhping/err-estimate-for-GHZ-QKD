`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+u8LlI4K92lfwXJqMwkVYKfuYTSYxO3Ipoe/qJb+hPoFuMr29hx9PSMi4kLEdBl
RMNVEv9kMqW54RvTiaP4PS+k8VKg0D5AxRJ+rgFYDQMnHkk/ikkd+qpJKJ8BpY6B
2bUF0DCpDTyzc5mML9Ed/bQA1j6CS+6VNpjmp7AqpFPxflrpVZASoxG5DTv3dIpF
bGo2SNDkskMi55slZQCyf6BHTrFLW9yLf+anxGLF+v7WXBKMg1O8Db/IQtnQO/a3
xJXFYcCsifZr2rK9k9HJqo/Wiavv6SDOo4cJDC8OcEUEypfkGUyk/2NrKyAIcaHC
BagXBLiRpl610vmyGUyyjln/CUFnPG0H7G8qUDf54SW5ZvTvrPvloHdlkp/3Lpr3
fnvV04GipfJSFMyUg2aa+1YSsLQCxzZWFh6huUn0nzn6izc13xvgOKJ2+57dfSz0
FK6ZkAlhbD44EKvYPnFHIZOHuc9VhzF9cuUQlS3MY4LzgKDKoHFoMgcNAeVUYUNz
kLgPTETCA2mtQDBKcXRRMgQiCxxl9cFl/+WxXuhWu2K0uFdc41FxpOY5P8s7j01D
ZGvBsnJpjyD0tyMLv6GlbNwRG9HU4u2eMZoq4J6sL/5pUucDMAwGVBEpyI4J2A/Q
HcZOu5XYb78CD9pI3qEZqta3uYd0tWVI6r2VHJpFrN0/FHdWvPg6MF3pXkEYDsQ8
hzw+DMKwyKIKEGoCKtIoXkJASVnuaFrp4u4hf57TMxCdSdyXfX89aXJGg+ykHGXi
W9yVvRmKw8kVhpC3yOcQ2o5dRiRbVhRyovkXFAuzAF/rlfLF2kojWlxrNVdS1y8/
jOYeTrG7dOYLYMJ46tEsB2r2jMlqW48uTVYTe7POsaf6U2ydl6Ofanr9HBQcxVI4
i8bfSV+5RgIqO63HxYltgriC7R69CR8gMka28oWB8pqT0sfGI7yKHEPIwYDQBWCA
Mrv3cmF5dq0mmNIXqQAYPw==
`protect END_PROTECTED
