`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oE3drEODKKXteMIDsbkPj1xNN+YoDabiE72EB99ZnBSIDxTWJKkzSQINNqrM5Pow
ab/Cm5VKrC/SiGWOMLTvC7xS/6Tz2HEtnvyXqI5to0fBpz/1oZ8HAnmVkfrzf2Pl
oKVmo6ZBmI5EF4EoA1s7TSJ5cA0t/TUNhn4WxJ++p0XZLpuPocqKK6cG0K/ncTof
EAjLbrYXbwyP1k8TPLR1uyhy/11V8wMjM8/dMj2T1gJwMkaNkP9hc8fCCX1U4mkF
OtsGkgFgs80GVHzJ7sEOWW1VcDlVRpgPTbKVQFoL7DarmgRyhQRNijZFnzbCNnRL
G1odTkOOM74mmKpdBnHtBW+hIA5+6p7eXTViMt7ZYzC6HHdAXtTchLSvzPXNx/Ic
5QS0c3SWmLm8pb+mxH5u5PNu1cGoBC/rCazB/q4Y5qoj9wm3Qw5eQoSaXJaVjiH7
Cs2GDwlf3q89mf/8TyRnp6+5mPiT62LiSBidYXAw0bI=
`protect END_PROTECTED
