`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRbr0LvmoZ7mqBvCCP4TySTe3NlsDj5Wm+2kXTT/hlEFj8uxrMe9OMPs9jml8LkD
g70/oLaWvStVrxVPxW3fu4vD+YPlI4y3Lxg3OsFZAPI1a7IolgmYJ1qQva2+6EDT
O1WH0OOXM+tDunllkVzt4gpy0U52lvUsbj+Ei0Z6rcr8zbIZKxRj/L6a4YwNwool
gag81fRoaxJFA7DJpakTcB0G/WKwPi1YT0n+DY2xNfD3lyisjOHFYy1cbmcjgDXd
Z68gkzU0WEt5Hzz+iXImJ6MrSFk2TMyqwyYxXbpS/4Zatvpn8EBW6z6FUHAqnDVR
H9D8mNRKbSsvn9IkhOknUjbL5M2Zl+L4lBmXL14dCPP0sRBpFFZSmv/2UXYWzDZO
uBejtLWfX929ArTMq9qjp3QoNkEYwltojlhCDvMoM6Ud2pcigdgSU2ww87PXn/O9
nU6ny10Pyj7umpRaaCSdr4m837r7JsHEaVO1bGCV5YrNwce6xMcoYtpkqPRvVYIO
A26OhL5FpHHwpinvj1Nm7jx4pPKFRzNjOhQ/D9+vFEoSL3BhnmWFSurGPpbSOLOm
gcPFIGajngcKF+hgWdodajh4RPhsFqSQvDo7w8uey71v23fOLFEG20OaHfSWBhKL
pwh3D796F9rpGmpKu8SIW2NyIft+R8MT/gOhHdUEgYYvd5ikv9yhknIvPNiNWPte
qG5o8+iCfJkCFCc9dtFGP9dqOff/1IizlnKHLaRG/HyL67Sy8JILwwcMl/sPFdIz
X2HjtYcA6O0/S8JmOYJ6Gg==
`protect END_PROTECTED
