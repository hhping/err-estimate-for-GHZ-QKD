`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GhS0BCN93baVMYtvOuiKE+NyCxO7JigbwJKnd4j7VxK5eTOImIHTud5a/wnFvAiT
MyUETIAJ+mTM7kk72hmWKHlHuqUaOycwvngbol2hKst4GuWcag2c20kIL6sQcPh2
T0JAdi+R+4uKqggf9azSixYmj68rfo9F8rYTcIMZJEcaaVWs2TgQpeB/es6VB0NJ
9ZrcsDvAxdYMXQyKSGuTSK/mXwpX9fboiXa5ijZbw7zZ6+MjVU03JvWE5Ioi1Kj8
3DQAEprK4i7bBz9S0eU1T/qWBLBAX6tGLldU37Phd/qYoSEWF0Ag16en4BlikVm8
q5r2PeIcxvqyI7YjkWsy7hvH5FRHcFn2eB2BNdG3G2et0AF5jCeYs6XyXNIMG4yZ
geuk+JZTwS/mf4pJNBREAyuwkgeFzP3vx8C8RIkKdJNosblD4RZKPClsHNI3/KZP
aSqfESUhjVwuSWerLNa29j8Oz8l+J7gIE1UPlfqyKYj4EiRPpvULk8HzLnh4I2Ml
oh/d+QzpMqLO7W5+lw2eohUqLqL26cgYCCRMROX9j03enSUypZ9AYZUhBZRCxwJk
ubZw2nIJhbMirSILg2hYfELoAw2bxm1ly4Yk/JbLoVs3QwheNpf+taVfjC/h/2vt
pmP/PNbflYxhyIGEAxgN5v/Uxs5doFfVWPtFJhmn3UwlQ/XJsRRVREmko4DZuvUI
N4DkxklBky19SAIvFzxTZKHTpWlvmtyoTkwOeAIa4+63h/d0CSuT3faZjuCCufVs
rZalgm/0e2jR9IGqcqzpw7MMrVCYo1svwoZKDcCbwGKYjoORPVjzxAkonc18Vd9k
OBAp+btvaiRJrd9e24sUrp4Q9lTPskVCNJXuJO4jTVlnoF4mqVtkj0fYfP/hMyox
xHOKDJZ12Nnu4elwpZgHSXx0CVwcPkZ6D9ma9/iGqO6tNpzDitlp6aX9hVgVjcPk
AA7jWdRmdviCsNQ9UXnQWNiIBCQIV5pyha+tzlR1no3ZNozu7X4UAWhEZp4FRydu
o1pEBNJFV/tQhmBqwyd4PtOS6n8Gsei7sljfjPm0skfyUi167kGjOVTh96UQb9IU
KbCfCm8nz+mIxXnQEYmzQj9eBwabD9eTI67J+YiuzZKnQk9+Em8DVxtqgnkRwR8M
UM9K2gTCgDw9Sy4I6MlqRJfRPCpdzo5ajcU4Sfg3gfgcD26IS6uxUoB5z3trKL/J
lbWPv/3lOm/H8sFEihrTnTCls9LDesjU7X6sKmPqfT5BYmwEFyg3X/vdZibl7hnZ
lUq6KatWx5C6UGXrmLquOVrc9sGmbYcLKFGbr9Q3ZSu7IOXXv91GhYcP9R28BNhf
ibLJwwNSHW6/YLGTwx8zL6X9njt4S+U3gm28n1L5I1Eo8l7qgUOJwSTfqZ8CSePk
hbXjw8f4H0dxsV5dTmOv9xhSWLBTN8WqAjQPMIC6t0W9qaf8CaPzBbG2lWlup+OI
gyrPiCe2SRRolfoJkRAR88hyb35seJfUCyaJkT+7wPxrxyk/rf1R+5UpjhGo2zbW
gsp5ATQeAW7/rTrySExdhIEwXd6xwVxcivYLjOkr09gdFgNGp3nnq6KbKpChLfTq
95WiOlfORscMfkktrBVdgM6jma2WlEke8cLnr1420xaITEvTDG6GME009FJjnen3
TW9t6W1QkcuD/zqzEOyrOI4cGY1rbR84GRc4TgSosoU8UMDLJkAsb+I3hOob4Bp8
/sbQkx6jFY9rp4xb7woRYVKQpI82W3d0XkkbMy6C/NVrdR8NkfP/T0zSc6SLNrQG
qAutJLFohQNLSzsYlQSBb7z4ZC3fMgsPOS/L9MqIEUJ5SjX+PKl1yJ9zZOQM5YZ5
cLVwRlYWz8z0IO92dH8qsuJLFYX+N2XyOQVCIekL9dC05684Xyse+aPhNgZcmiWE
klNrX72eTDAN38zLLN1qc6AZXYmRKFR8ssYnzUnGAvttscM5K6IiAlOIhikiXtQQ
LfB3wwSRK2CMoNXiuZJZKRPJB0X+ae6Q15+Vs2IrCgdCl2u+RhqMatp17u2iiMk7
SxNbtgQziJkzhE8Zcd5dsDg0boexKYfGcNV9gMmVbUa1UNO1vPfA5I0yOyORcbGM
n3g6VZ5ix+f6d9bmrxb3O3xQkv5dUzdBgmCVcUlhYuty57UI827VR84V6mOW06Wz
XcQJE/4B4ST8JivEK9nuDAzo0j8J1JSA4Y/PaRnJB/ZElNb90cm6EiCuCyISWgGk
suxcxLdL0L+BvDftuNId1FLhwOaM5Q80z0uBC/YyafX22OkpdfFXkwEPfwIgiiDV
zVg/65ibE04YQQHSuTRTzNo7A0w5/YEeBeGSfIwi7MEV40W22UpphzyzQFAzBHhw
ZoMReD18M37cGNhku9pnRlbdf5ZiFS4o0iOuZ06ZcL3lbqEKWhfojN59oLML7wHf
LhI2/Fyw+Mj9kuV+KFM2Qp/mYMtTICFv+UWptqGpL019HUDPrUAKfprDPuUsl0Dz
p2sEPqJHfoqB9qRuCTv8sBejKlCYT86I3bBn3383h0u/qnxpC65Wv3szGpzHd1yA
ntHWBzyxDVh3JnS78LkjCkINx7/cD+y9OUG1VOprlkVQ5us55Vj1Z72Bi4cXHrrK
4Q5tohvqihjT7QcBfsjhgvwWvU1/zfAICGVbeYIb0drboSdcqiL04RUitBa6JvIg
rsbNihAA2qI9rF4Gj9y926PLOz9lZBco5VARuW2WMhYtrex06F5qnd8VBBaYgBC+
+gBVPSWjg6sS3UnC5javWn0kjulIikZ9xDZix8om3QqokemNhjW6Fk0eZKeVC5fF
VY6Qv0RpFX4hurJCvO9Vmxdx33Ec++dkUYSwVLyco+jjPLfucVjVDfe+WOr/ry5H
v/bO5o7K/8NAsbeSirCkm64v+dFL26mnQ6UTDKv3QSRq9Apq4Grya11cb1tiwZn+
awtCs1EXYbwvqCzadzC88+HrW+0PRuEd4+o6WvZvYvUSxHJ+WY0vtLu7rrYW/zb8
alA8eI6sguzQTzflxWi5dBHFmXeAH42hVaKdVSclznUD34EKwJCb0dVy3QzHTlsR
jIYXh/+hmq7yVzsO0D/FAneXFhK5pSSjrQdwfMxLqSGVXwbZRSO177E5ioOeMKB2
knXdsC2SQAKsfouAhcSamAdi/FKAUSdTkNFSInoa+1TVD7V28DpIGg0DWrvaEAOs
LW0cDpjBUNHrt9LlbSxP0di7Lu3Y+dStcHufTqGeS7f4s0raRuxO9Bpan1rwjtKf
lqqeHyf0NpLYw94Psx24UCwbiyAWoH/6lU95nAbrAvjiPpK8Qf93Qi9l7ABHBPrg
zxTyDxJdbM/1a0Nb5VzsikMVjJ7r0JotkEgYnHAC7FA16atY83unLt/LufftKPCX
4VLYMD7WQfmxgQbxqoGmFiTBYWSaWq8RvbffWm85cRmPggAASBCjlxuHqzJbQ8py
FurLiCOywH+SxxcbZBrQUvKxMckUoinvIsgFpzc94x9kZzfBmE1ww7/KL2FVM1BX
9VYVfxJqKLQMj/5YiYQRPFroxTKc+WXVuWwYIJMtKS5w6fuLzkqvVQGVDix7Fa3X
gXLCThpPKoIOwc0wRAyAmT3lYsbK1e+Pn0p117ybGaravmFgVKsbfCJIWYiK+H2Y
Aa2uDt1Ew06Xqr7bLJVLKNLQWMOZJrpn1atY8Pne+xovLIO98qBaOpWHfyxbfCug
wSgWv1gj0p5X6XwMUJJ0ZzHWUNndYzYphTMgR38BWZRneLfjCIb0w2sGaq6YwxPG
l7DTlPRzDM61nWHVBxc/hXeKggjAqcn9eiYV/Wc49g2nJ15US6B0z94SnlD1s0Gx
FgIMIUlTLCeVtkEu2EJBPS8LCpVxqN560kpCZrIsDg6uxEUqA/OBGextLse92hn3
+uFnuEsiJnuqnZxLklRA0zqnEnCb0hNlf9A3fLcaLwRhKzfTpEajp1vHUiL/HLTz
ZhOQGHo7eUJYf5/ZiFGcozYZ7ns7XKDHhGJyoDrgbN382qX5jpu6gpuSrNmzB/ik
xHnmPznihDvbMVKtie1Kx9RfyDR4cQ+ES/uoEjDR4YMADlLkd6ZDGW0m1tuVu1ax
5ccqf+R/Z3qm5h7CChDYEhhL3+nB++F4NhmCmVs6hW6AkaW4FEUmBZiV6VIbd+0d
RdmmZiDPFW4JEJkdhWmwUu90iFTwmdi1zWpz1JzQykhqjcDjV1hjXlbUU5UpNbu4
NM8ZPekA58TY5J02N+HLPzqyN0ps8IM1x1bz3DbX+1JMR0rKA7MQpCLhAwGdBPGW
F5tDIMdwhxIycXu0GE4UsZj6y70VKM9AieYaguvQED99+bcJJ+eL7I0nuTqfKW6d
jCXVCvVPxJjlzosVzhktyWTT4kKA3DBZBgsKA2/TQ4LBJk/hG+u+PVjLKV2xNfPA
eUiraTc7bKbhFS6GzCy7rO/QSvH/c+7q5sG7FLoWJZw69OwepDVgxFzoP8vci2wW
jNXdu5sD/GnW/8xTBDerne+qPoZf9G+9/IIFUOpq22RKklEEM3fsImPXEfRmg7h1
jhH9WYZIR0wBQfDP4iEVntzNQRrwu8PPLChRQJ6GMItPhumOcnwC4ghm2YEM2e8K
0XGPKOnWXhH9xpznLxmaIYVcGtierrv6XdbYIXLuYJWkhR6F8ivA557KJrNvx17h
Ms9nT2hGSPkW0dmJRMs+wdaicyie+LULaLlR9EGswFIA4qhaKmbhWI1BO6qImy+Q
vw/DEJoy4cZFYW/86ZC4q2S+nylx5NLGYkfi6TP/BvZ2wRVGJWvAq4BvYdAjI60g
xRiMDPPa+yCkfDJTyqOQnadlcC6MYW0hR5SC+2lkfsA4FAvPRaaCuZjWstxfEGoz
LmBfGVYMlksSMNHqSvTQMXsX+g1LmcZb2TolcK48L0xVaeR6dIh+YnDBNXdhpET9
726Y2D+vz4Er/RljvxOYs/AWSQ6j0a8ZnK8CpKTnsM4yZTPaStEljeoad+2VTAqk
6eN1WuT2BwmTKHFvzkApfg+6AE6dhS7evT53FCqrAgAPCw33AcIGJ3FjT8jD/8Na
PutKpaA3BaRkGnJSR/7S8riNUFBWWhBeGY1RcQXK2OZgML5S2xvM7Jtu9UDrnO8+
d5T5LBUnW7sy7r54GoO1K2upqlQPwzWOoBOmm8FFKEU34X1qNBExt4grOTrNW58r
RKQPLrx4NN4srqPbdlQHVjejI56++itxtFvLI4SAPj7ZTksDyXzKFV3JHKlD+A+U
QzYh0gGY07zHpyY6iy6cjb0OBCnYOlFcbmT0Nf9NlrmK7FQqv6Ur1DHMmn+zSu7x
+RSK8xjMEUxF6bZ3JaZSWwwlEnNNDYnVE7gdFsKUMaP+FhINtIFBz5F3IYTkSGpw
E7uaztf0tdvOVrQm5Tx1R4UzV/MW+r4P+OJgphHBawsQSHkaNR1MYtSDvoHfwJjv
uzysmYdlpNp9a0TVjLtgvHTMSW6q6nwU+kvSnmsG87UiW2h1F9LgQgBVbe5iYrHh
22zsbNHhs4LG31U0kAH/4+wfwErRFpCBaYzmb5HNft/yYcgqxPIHYOTqSXyUUNRk
8ZexoJ4K3Vi8SAPFpAOezmbQAT6NSOSyf9QXHworH6OZwd6ilufUERetcdT+oxkv
03sz9itkj0dBn8tsZr0/TJCv/EfEhnrEQd7vDAK5jVWU9kFhKUstoEETU5cTpUNc
QeDsvAlh4KmTZvZlPcTPODQZQjuh0WF0h/ceAKEkgfIRQ5ndIo3sLfbNBhrXK/kY
hw+sYFRunFQrJyDiT1Svtrm13S/MxnbjXMH6PNbDZWlRVO1dVT2fq6MxqXCFcgzr
gCYzLHLTFsej6/FGNPg712mmPuqan8rTqfgEZwMsT9g0Xosnb3uQ3gsOegnrQcQd
+C1XhIM+d55kMtJiX1kB8TL0QM4TQtxqOc/KzOBDBb5gkmNtboKQez3OWaDl7Rti
NZpnSpya3MgzMt4Rf3UwOu2sZ/bGUgiXdzxX4N3919nFMUYitvhF2EsyMadwGDYw
RDg9S8O/3rfQnnWAkBIUw/AnSN8NhetY690d/U4lnmZA+WOKbC27Y6WEf8km2usK
DoU2d6TKkf+FR1x4kKGgNovmlYVcR4t2De60iHdHHvucUPLULndJTUDCW2vl7mFI
s/mwUqnyR/htmjTi+k/VdunTtH2obe9ZvnmJI5UrRA/RH/461Bh23Nd8PaERL18B
UxhQ0qEA3ESOlnFR02CQJri6NNpm1evDqkOTGa7u3419bWAypMeaAnC4Rqw/3TBh
tKYeiUCTbZbfimkXTETtrtcQdEt2sWVyr0VF5jUG2xDGplS5j/ZZvfmpbOQPVMgF
2dqjrBCslhdRFEXQPme+9DPyIePqXMJuhd4oEivG5tsJjyDaeBcgZgdJJ/90tXBG
gplJ6PWeLyGT/oncML7IEW+F4IhAO8n8NL2pSD8CeeHAT71EPahynbQyARfsQ15Q
4wns3FObZdU3wykdPPoWxkXGNaBqg4ptiZfINkuoV/w8fqpzhzHBGF7aMspMML11
GQ87mV7zx7nG0kNsNKWZbSAPuPCCVhwPhIAv4pDPT1Zlq+fWiTCZJzXZCnBRVxgk
dlzMxn6VnOOFcmD69jd/j8x/Ab1du3NFPLqTrJqaGJKy4RiCpKVBtUpFddtCFRCz
+hcwVJF/kp3YRXOrHV5MHJRHCYZ0bsdrioCcpEEhzUuHDw8+l3wfIZNVHenHE+Cy
MZk7hqzicgxs72TjLMymbWGpQwN7ne8Z5fZBQs5vfx56wD40j7n/+PYHA3hyVgaC
8gh5k/4H0tSZfC1S1xzLd0/SIgNRF/axzyr4VpVmSsEkf63N1Zndmf+NFk5jdYWy
vvrflCr7RFTmUnwHx9diMFoMaGnr3rbCCTZf/KlLxd7j3k219vkknEEbWXTNej0m
5j2k40d8OmwXvIEYJoGbwx5xuH6NtuIyliFLj7HiqwTsZc054VVKQU0zno9cz663
zuKA+NoqkwLnbRMw8neJ0404kPOEj49hW4B3c9EsYkCM0ARrI8XC1BhZ9hhlpe6G
5s6k+3SbR+wGP7ZMNf9TbFW8DMa6ROwTxYFQwBGqjk5PtE66RApbdmrzHC7Vxz8Y
MW4zNerw2S/TA/Ma3yz/OOVF6w+Rjr9D50NgsudNK1GvU6hbApz4iw2gY7Fyhx2N
tfiFWZcwdPH8iFW/2lZO5KgWbb5HknX6BqXpByoVZU1ry8/RsHc/jna4harYi74o
zWjCHAt/voxn9eN4H5xVzROoPABSFnDM0ewVGPLtj3SoYeakF14plEhhxJqbGdCL
J1aPGfbn4osnwY0q6Vm9LBPZAid2nOQF9BNZradhxjfyTdCk+m1o6xgOHjbiGlSp
hbxThMt2xtoGmueXHEFlUGpdhKJelC18C39OIOGcCgvVIC4LY0U8tTx1uiyt45qN
0AmqQQXZ6pc26LBdV3QzCECNppyxvuibb1ZjEM2pGckuZSySZe5XwJIlpGsYuhPn
EmAb2ZgDKCKcLjaVjrIZABWReBApU7Q5M7hW9jGvsnTVvjDNozzx2J+alp/lGgUF
WcPLzEX4XSEw16g7hK7lxgaq+Rd0/lNMUigxiE5aX8A6Be5xBHs9VqUgj2eyYRi7
PeRpF/0pVGeaAsSMTJ3BcLz/eBFgGwBq1+ak/BFwdH7IJyQ5YnVRNgsizBHcqESc
zVb5lMUc9Uxd5HKa0wpRyCW4c+fMH7mMKXbOjAwd2lCVnhjDit8dz4fxKsUy0ta6
wkdfvqCTgmb3m7PJMRNS/PwTVd7Nob4dWltLeT+0xgHy7ubIeAtewxHPEVav/Ult
aPdlRVKh+TvI+oJVlm2wwW1QfAcDzrm/TnCfCLMILAcV49+yQIl3MyLEs4b4FfKr
jBmPYIRigILADF/2C9pPdA9T142x1Y+FBZT0iLbw8DgA7PdjLPtyOYw+SA65BT1+
tuww3+Dozl1RMczDTiKrR8Y1BOlr1x+Nurx8VDqUC4MOJSnfgS3KLzRU05S9LqUN
3HLKb8xk2pOEtceBOCqM1kncW7cKxtoNkjtzd8L+Ehzpw4y5Fx5Vsykhh+c6h7EK
IiVmaLzlBUhSfJhVvhtyKNA5ZxsvXmn9AueacXuY5RY=
`protect END_PROTECTED
