`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFGNQH5xjy3ym5+Rd1rLrSYiiyft3XqTkOKo/kZO1w2fwgNoSOgj8Nl3ahtVxeEo
2iS0qvwB3Z89+LJ4sfm7TCcWYwRB7q64NthbvXchxlshZjZFIc0Y1JNamN/J6Ujc
lTICqcdo5O9MG3FXgfBU/qurpixRvxuOMy/kRNn563YuVkoRBhy36R7IhJjyoIkF
P/sO1iDTi8pkoE4bHhrqXIL4wK8t10BUb60ur9d9SRc9NIfLR/K/juRHv1uQlC7f
GC/KVLpz4Zz2xEDn9eJT93ySo9JH7TQMmdA0KjXo7PG/I+R6l7LQGfZHlZqRQDAU
v0qFOc6Kv5sI/ftCnVTowWLlNy5/I8vHgdXxM3Bqwd7M+iXfL4C9d18H97Ki5J20
3dD3dNX3wNt2wZjuFsalcN/6tKDMJPBAvXI0yRU23+rrvoo2qNw1q+TrgbY9KAAt
xP6ALqTMOLJxkbYhGQ2FUoBUUj8ChSmtb9LNtpb+5jBnhIQMws7JvmlKYqckPeLd
we4lAHqbLGBlbfqU2J4E1bZPp/hmmYLIse4SeR8tcjNifG7h3xrkwFt85wVgNR/u
h3CjGsNxi19M01ThZcYc0KNjp/loR+dJrbE81S+ZOgvSkoCv8WTn8kkMnMAaGTAD
dv5M6taKgOURMsovgrl5Bg8ffCHjICtFveoEy86QTiq5U4KfmR5DxgrEBQ0Hg+V5
4f4Eq3Wnc28nJe1xTXFoL2k5UoULBx8zPVqgc6NkrwWloPlQvZyPgZltlXYGYRNW
`protect END_PROTECTED
