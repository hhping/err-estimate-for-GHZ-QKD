`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mom9UgFTn3LaiquSEI9kOuPcxbycxGnr8XmC2TM31LJQvPmnoXz6eJVazW4anTZB
vp772LfYSmfFIn1gIEvnveCGMPlsFmMV1jOOBEsOTa/u0GGlVdr9Hdom+LvQbU1/
2WiNVpQ9YQIJeb1sTpZlA8lifrc3jjyDUbeeL1qSo2l13LrCFst5U0VycI3sl3cg
G//j8yHfWLZDBxSu1SbysbIzSYdtXUR/qAPDTECC7RsMsp4lQQwErjGBQLSGDgN0
a/xk3KTwMEVcWB278eXuYSFQ2n4rQFKKWohWH2+E8BHDQEo+vhbUdtQblmQwnsQX
QrqDPnaY1J42vzQ7TsGYGTaptUZiWGFjJaUHgNXFHZxYeOIlBQsLMTmySzY0tB20
OcdoNZxfih7bEyXJNp4LI+plHwX29Mqbo8hYNIBP7HJQK+8Ew5FtP6N5lKF1/3EF
DG+EmKVsV6RIzYqa/KId6+2IMS/eaJF3Z3hg/ydlvoiln/KGp0JBT93IRwU2M+qM
dGlaD1uaorcclpCTuvrVKcgMYjMuW9a/18o69/ZboGWdOsyGxNusztqFQReilg5o
DKqbEt4EpdxKdowUbJOGc6FjCO6yLddJ8Ck4LLEuBzWmNP1ZgNjzWjBGSpQHZni2
/6nTvMZcaKuBjwDSIW/jEeBzohFE0yekZohkLFFoxNLBpE5GZEVoOdOmyNBUo2og
K1bjWkj06CPuqsQEBfwdwJgwa86xR06jln6KuF67y9RJHL995O+wUn/m/dk7yrvF
eDmWwPrcZfY/zERvOWJRkJc/Fl6T3cS/JAVJbgpmv2A=
`protect END_PROTECTED
