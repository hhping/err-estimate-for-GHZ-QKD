`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLsrqf4uOtM4W3BEWbl/NDIBjoRSnMNd9FTmoJ+4j61tiZ5MLgRoS7IzWp8M9vvu
KJ0xIalUN9pFPJ2fmGK14z2UXjYnw1Ym2AFu1Fl4k7thYSmaCwKCf7sRa3GEY3C1
/lDNMNEcyvHd32HkU92FhWyPM1522d0jxg9j76iWepER4Okna3vasNnoCjorwk1I
hnnFPe/tzzfhRJJdr5OwQr4UQW2qLJWSFqbGujZiYrjcbYT0dH2b8wXn7srvQOIJ
2AXSiUFj3A3hQI8Uj/V9Q1trw/+zyBbl0UxxLhCtH03BYSYlVupwUU7a0J14nMLt
yjzLovYjWjzbYxzlajfLjw9gfYQv95b+NTtp2d8mwUKboFl/y8CsLLMeoDI6MwZH
boOObf6Kz2X7UX8J7UutP8VtFmIvOl72lQDhv+tBpEeQ4DHEggtTAfyy/kEXMxcP
iKCJhM0xlEhOYiNXPpSeM1XcbGPzz4+p+kQnJNKycw28q/pI+Mtb83dPoW45viog
VWd9Fcm/oZWcLx5YkKcQyJmDK+3/EB2IntVXeI6pus43xA3bA6nSFqhx6oxMStdb
y38oIQd5tL/foB/YFndL6HV8Y3oD+tAc7bGYqkK/1CYxPvbcXwOs2WqGy44pQjKc
SDclQXBZZrI1P09vSpeZ3+80iXucRwDjPA8Otf7Vl0ApfTwYWE3QYQw82+BUH9hN
IwTy7AYV+5GllQz/IiovbczwXmCoeorkKfFRaMWmtj7vOyQtSlTjkx6OG18znKRx
8OZ4vN38Hm1d8Tw5ZGvECZz+kLStzKoh87+Oy2qXw5hy+qFbteD7YP5wpcp083DC
+zmTaH5EzVlzuMMTB456r7AFw8wRFihSdVzZQa/VqXd1uiO/6jQTHL1rM3USZA2x
KsFlIa8G6Qf7H2+1d6Uq8qYgwUVNRyInfyOwyHBoN6iUleqKgdSNCiErmpgOQDKV
Qkui0IsucRQy0q9y75NiJ/GdFaDwaTTyiaa0QdhjjUaRrIQpa0JTCBFaIL9k5LkM
qHZyTrDdygLm+pY3l2DQbAwheb89+i9GgzE9rbygFuzjupEL7HiU9EK4b/S2+yP3
onZG8dsy4WSe2dH8C7NoJJDqIagCn5uUjjsp7ICLjr8c/sdfH08nqgIoqcWugCzU
0TrIlkleN+Un3FA6loF1NK26+HOD4WG6n43yGiWhJTPE0MAQj7wGr5mpcHII3ABN
2gpohZerh3KvDS9Y9+iuI86ReYXK4xnA/JEV2Qu2H+rRA3nyuCoS+arAY+L3xjmA
WIMO4Yp3HaqTU0E3JVlSV+EK+OrmS+BBulCMkbIViufAYS0zWXPJfG0/YdQ+tb0Y
6ZAhmSYshFdV7jwMieDl577zuz12dzI+jtpGhJJSJ8/Nef5+Zi56LnzGe5STMfOt
MNzqJD+YHLNklU2SXA+LkWWcNpXu/vydKkSgqobJOybPiA0+Cp+bV80YXqsS43np
2deSgnVCeWPE3/JEn8mqZ+hZOoorNSs1Etk+SDlCSilmS8J86Jjee65erAnH2kNW
mEiIXjcmSc85AOX5Wg6t2oqoawB5eYzCZHFDcMgVkpbXu9mIJmqkQHnOz9TyjZ00
VSXg4m+TH+FGSoHhPcU0zwrrD3+ZaYDtdlI4nqvba8dCCvVhEut+np/2HPHkGmaF
cVQWQaVo5Sj76zG0cBNqho5PnNgWnSCsy6EN8Vpn6wlQUqmVusaA+2N6iGAtYrwN
g2vRCL7ZC4gnGw0i72PckLpAcrD+W9xHjzxU1Min9HV4UUxe+fdJ9Ofh3iezi98Y
WBFr3U4Jk5FsADLlIxlMuxFQJ5l0EQ3V7yX+S1L7ACj2IGlr1wO3/xRx4PaEt8eX
a8/heedfXfjDXLS9fyRjcSln6J6q6qFe4eHvdpE0mSNbCy0Cm9fxWt6GebhH1EAp
oJMr+ODRMv6mTTBcYzzrRyXSWaXeQUZjDX3YQaVuD0ujfM23ugtvnKyhw1Mlm9pq
4rCoz+GTibBuU4vfNXFXH6VKX8uequs8h4V+nJ+4AT7Kr+TxgA59TiSamJAyhHQH
n0mLw2ZkE49aCDGb/neIaMh1hE2ay0xB14I54/8Y1wvqAZJVXNU2PCRIDhR/bAyp
y6+l0I58Y1yD08QxHB7fd9Car9fLaaeUx8aVLpsuxmFptWl4extub/KQgMKjbt+2
KBAHNT7Y3y8uCaj7OX+MJ1FOgHxCV+EQhlmp38K7pN9+XqK7N79Lwb8MSDAciA1I
ND3SODb47Xff+Dp18losEt0BaTPVDVQGQjmDhfAa5ED8x8Et1LVX61P5SxhDFaKR
UXgfNUmdG5QmrBiSfeiw1Hlg0a9CcuQHx5FsRJAgmsokFQYVyinvxOYuSgFQ6F3Z
vjdXrJmbLoN4qlCA/T0rLlwKqdQVz8wDlmX0346v2Wn8y00qphto3WUIx75r6pIR
ZXhLkUhEYFcLNVUPX2k+BdeIg8AytxU9p+GbCIqfL8c8OqICEfa7IqxS9X/8m+0d
MQm/r11up949MWBN9Qylf2bgqBNgh9ZQPiS2bn8dH/Jq/Jyx/VX715/U8pwYAdbF
OgOf2K47smLb8WNZDAhBOMgOnm9RUOLnN7tFn7shJxF2d9brxbsR45d7Dudkyamm
jgfe/9dFole6DFEiTdpImM7Oc2fzsDn3/Z6IezRPgRD85wHCPNIOC4khABFrBPVw
LkS29wb2M/n1WSI6pZdxFXaBorWtRbHHLsY+nZlxuup3gdKycyrWKOoyQpZTnJ0d
d/ZLLCXVy9aBCaZEZD8OhbLZ+FamP/acz+nStdfT6P0gAmQzJXOK4UMJibK+02Pb
n93rF93yORBus/iw61Q2iFUvh22OVMBIU/ZLPAN97k/KD6WXcV89PcwMAadbWFdf
wqw5S5xK45vDbaYwJ0YTKbLRjCrpsqWRPr9BrTjVk6uyXb/JdQJ3FRLrZl1UzWNR
+KOef3qjkkXwGMgxqRwUq+b2D9LHQfY0jrX029E9uv5La75v7IlMAPqsxeA43BBv
Jm4L5N1IrZ3wnh6EqFXMkifDFDpzL1G5VkVEkIsQj9j7qVXAxZL0CbKuM+0vHBIj
zga58UQDJvwJSqiATrTuqHdFrRgRG+FSDD1mpVcaYX6wusVXk9s++DYdLeif2A6b
7JWslNJ9JDckqqf/WvPb3zrygiPE0OfW8rTbtKeIGVhZS5Mp8ZrkGUlLcpl75q//
YTAWkD1CgNl+x3XMmBVeVI20D6DQ21P/J+TmW+JCAER/4qugb97Z7CYyhBZk4lWX
Q70/zYbZrj8ofnp1yh8WVKhHXL75u54R5uuap+s8mri9WbRGszI+bk+5qkosClZn
ykaHCkS1eLA1pl1UsgQP7MKPikUSiMAnYiYuS6LSNITPRudeVnzNLszaXIl5RUYg
WPfmv8/lWxuYOQwUYzauVFbHHvAqZgMK2db4g/MiRnhg8NVOpB0xwbt6ToIq5ufq
rH5opWhRBkbnSv2glCFdh2sSzUVplD28b04FGXdIybONV8zTdu3YkSKN+1KAYJVX
DJtLVbxVniPYXT0dI7wg61Elc40BnQwvaA1IdchZ5HxLhmgYWBGfRHeN1WJwGspC
UGUnZBtrszt96oBjB7NAiS9tS30N5G0SH7ucTm9qk7/bhOVrSaoao4LsweFYuDY8
V8cfFpxXrMF8akPBTJQwFdtjE7bqUKIbwo+mY2vr4aseUhhbkNsKxjsw53ZnPKQe
aImYPBetmhnGbGQJHDXaEGOKPy8Wnie/L8smxsGcKZlTP/3nJ1CdhKx1SJhQ5haX
RrpdAzyJVlHSLqKyER8b/5D7m2wXcIvltPiDKiGOx4X+W3QLzKgC1FcQXg8h8Xns
OihVzLdqQMMf7pzOV0BNTPEGIHahgqcbnpyRI0sFVaJ6zfU5c24YpRr9V1S+j3rE
wjbXeD9KVuU0f3nTuq9RpyLly1iQswomPB1kNIZp9+sTUPtQnWVIQFvfgfZ7urcQ
ZcuSKauiIeGP7wmxA0QdFjU27jxCjtHdmee1LaQIBLLR4MW+SooyQu0jYWR48mzB
LVC/vJuAuC5IEpPJybYABby8JVOL8AGTzJ3/csJ9b9EnuJIGWgtYP81TUNN+L/3x
906DO3hMbD/YykpraC7UggwQamD9xWyv5axZ1M1dURIWSzZyWTr6z4Du+v41kjA3
6CKh65aR7qydQDMtHA2blCfsJqEy9JekXDNWxAngxntcP9eKHeLDapTmWZZ6FX5F
seHLLK/DCaujMLI3XrK/B+LUYxhpT66Uxvz+qfTuvcfm+836mCNSAkw7kqYoHKrZ
+XpIUE2xey8GILB/SNftAYaQUTc51Js6ISDD/VblBr+P7zmZNU1VWXxR/9PzKmD3
k5w1X6Tsv1JqXVzU4SReoabFnxEDuRurg6GZiI8OtyieFLFgBgYkKiArvfR3tVOM
2Tzov6MYhiY2gESRp+LMnhmfglbDGeUq0HinBjnrEE07ehJei72wH3BOf9vCSRmq
FlPUhwIRyIJFIAjHDDd8SN0JGm8WorDEii5hCkDc4IYHPtGffQ/9AW7+95bjKTsy
Ze6wPe6rv3AFrbT5Xi3W/IbiNi8nyfrb2m0l5KP4Jeb2snd6INldqpA0N7TMSG8w
7DZZRCriSvJdMDqqmpXcJa5ZDb+04IIymVrV2l0u1YG3A+aAc+yVIn0p+IiupkzM
HNqv2z3eE8nNfiUReT8kmLA5oTLq+vhRkMdEsftM22u7obytJloonEznQxvBa0qX
4hRO7Oa8KiiPI+bwwk1CkCV4PSrjnkhvpbv0ndRxwvjEKV/kObSHo2xG0sf8s9K4
JWIeIYlUHWh3VXNjlx4U+/eji2yGTd0xLd1ZcoBRL7B3GGzdFKppeeDJWhhg4J/k
RMemqce/vj+XbxwasE4yFMdVcG6SjjcEz1QjqJZ+vCZlr1wTQVGQesg7IBp8f3l1
r4luSa+aKWPXAejuXJs/c36Ad93jG6qeaPSBLMQCGAgpjBNES8SaLJu+FzqAow8D
J1letKSiTJRzXgtf4QvxnolEwaXWxp4RC4LO83YTNXG2E+mu1+9HNarPp/wLefEv
vE0Mc6J3m5rIJ4KHAkKDQAin6j81qawMRn/woQ78l7YZsVWmN2r9gC1F43S7fIMv
lPjeqASW5J5lL2JSaxnRHPMVBNRqoXrHfaaqU9+JSWvLhEvFDfo1znjFgHaryRs1
SKBTfNpc95vSr3mCDjiCWsTpGXcNbtO9O2TkaG9kQ3+0fae2iBIxBTQ7CckE3+B1
Pt2gjpx09mbzZs7fCo3E/3KG49UR2skZTXwvTjn7YMPa6AwU0igAp+QISbLiaMRS
LwRUOM28JAqIH+3ET2moYO6ud/Pq2xXStD27ciku0+Ia5u6Qfjgxm+BykhHc3sE9
Z2kwi/EWf3zy1x9Gqtu3T2w6F3VxnJjvSe0UL1cLlV6OyAx4XSkuxfbzuy9xUtWV
08t/6xxBKaqrLl4c2A1gBceno2CR9GjyWIwzHLpLHIWG2f56f+I7FfbU5Fm8KeQS
+ZpUPzA8gel2copap1r0c3a3lHPix9WCSPFmdpcgAjaL2zWfjgdvHXuSlGD4e9o8
NeICfx6W2SDwERkH1sNGOyj1a7s7DDYd4p6Hw6ljaU52kUKKyIb93T6o8vI96FJ3
qPA85Mk3A6IxNI5EP6ZrEyu/mHAoqnkpA2L+NSc3JMMMBpJ83siXgMNfhyoNvf/d
0OCTPp83HbIYNx/2GeSJ4XKmGKmtrh5ni387kJNWYHz2KTQMNsfE49ogg3GMJOTS
pzVWh+eBuT+f/odQGaUXhEBhkE0qmJW5myQJYwQmhdvvVu1FnChiKfH3n85sjHsg
BTp2YygBl0TYSof3M6veKcTpSyRzWFBSyxkbKb0CChLKuT40N3662t91rzkg8kDx
Dn9Cj6JyAgtRkuKCe364RZxr3i32pp2cdj9xr9L59gIfJ9DFc9hOQREhfLjmwPig
h69V58l3e/A6sFScwPUQllY3mYkl8yvc4Jfdhaa3pYeyPSvQwxvom0RqE3qgt5De
3HwUph1BBeNPAqlj5iGAObPBpOhyx+16zfJNVB4ZIaFpBQlFaPc49K/1/u6yBQF6
ZA8J9g5orjo9Had8TUR5oSF2IvPBDgkbp5mo0b7+Nw/xKThnTiMl/ahSYR01takS
BqdI/usgeld4NeZX37xEkOi9kQmzpsMhl3/TNGG2eCJUhCBDGQ60xUII3nPy/LA+
lT9jauQIrBbrD1/Oh6yi8Xv5MhExAjf56CeuohkBAr6i7eGIjieF7JJSey+wHasR
V4dIrtyVxuKh4LEmb4VRL8DtdEdDo9S/PEig2R65I5QEXbxCDiKMqp5IdRhP8rVc
esmRD3UdbLZbQepzOu0C5tr+0z/RCZY+KkegJH6OPuVg+FqUajP/xhU7LBPLgNLf
ZqsxdEPBvPy6F8kwuYdIk/Ua3MJvZOutKa5fXAPhAf+TM207nVhhsRtdugTZTm+j
MZWRezMDuKHlH+052d7sBsMykV5HkoHboEcj/0ILZ4eEqtt28R6BzCtpsv4+1kXP
ruW2O5J7Kzi+QQ45Rxk2q/GWPngXWAhzfdeXz0yi6NR8ncqXzSt+uw4AJqJRMjhP
pqY0ySXo6/MdV85XjDrs1xk0btYhidHctiNy9zEdaBFh8uOIMN+x7l7GgjXRnRwh
99U84V7Ecg2eLpOUyAjGAtjsb2FzTF+f9P8xylW+fiQ86T08tlu6QHG7qCJpR3Dr
y3n72N3nDQlLeUzEgyY+2NvuA04rdAhEV8gXf/esBiALHTMwHpcGCS5XcD12SjVN
G5zn6bHfwOYys9pZ0gs0ln/XcNs3Z9ZoxQ3HOvLGd8bxVfYC1Sqr6mBS+P4McLtr
vLLzcWqUUBh2WD83OIB4jSLMEyb4rr+m1sfm6SiURqhylz2PpfzU7tFcbUoErdsO
V1Edepnuan3c+LxB/cTOkR43AwDnFtjFmN0TBWuFlpzewhrPoaJ/Yld5Wt9ZIqJL
CjLuovVjLDDNgcLsFUlVgXNWhmjECOJBGPDPQajOPdvb26CB+WYqHmMMUwU7MeFZ
pyE1UXivskilytV25FmzmeUweOF/Myb44eAg8yjPkWrqXWtxfRyxvbzInJkBMk3/
rCTEW+k6QWCp8tlCQB4T03e+nnn6rj/BgH2anrbrzoDcBRSUFs87N7px9PdRyzmK
NK9zuQZbgI/+W1Atz6YhzIqZ65hlFNo2GtBZy4v7CSLLNpEaj7grnkQD4Tww0V0C
dKeUin3v6YTrCq77QlM0B14XGyfz35iLyQe97NajXtbmyJZxFsb/X+gwFQ5wZ2je
JdA2a+g8t9VYUmjz4ygHYcLmstkMc/tYdwMHPUI4kaM=
`protect END_PROTECTED
