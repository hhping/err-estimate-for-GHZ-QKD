`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCjG5f4+B9YGlZwdzLqzClds6Phg+TAohL27i4uHepVEoMrz5yrxEDyjMXWdoRef
k4ObkZ8rtPs5YbGRkLdjrj2izgGyIBuzVCwUl15Vi7F73d5/d6dQk51CAIGgEUxL
j7dnDu8vrWMxWy48LajaoW1Yd8touYqG/KJGPBl/g7DjtaY1ocRWUiRXIm2fFDV+
6hqp8sBvAWYzR/ryQjsyMRtKFJLimpm8L4TQE7nv7si0XR3tMwU+VYAPx70XXRNt
ZCTu6YR3owCt9WVK3n/bANprTbcnw6+/HnAnOAOeINjfEC+EjxqWaLt8T5A/Fgdh
anIbrlCVIEm0fpxiE4EmxUQMCk/N9zZgb4kPBB3tyoIv8bODtNqm3F1T4Sy/TSPw
B6Odn4nVrnINpPuVg4Qy9FmO9UzavdWdJqFTlXstSueY1mC/ND4Fzdy9CwR4ucsM
ERt4ZVEj/iTpaDJIOW6/bGzhwOmjcrHnS2aCXGjLnkQzx35OfENAkVnrZM/p3Jxt
0EQ32TNy3TfrppKdkxa+rwS9zZMS86p4jswlfiNmIGYj6DFa0AxzBOVlxaY6rDVX
2csBAsu/YxwPthW01TVbEFpPKMbFJvdAeeHpHJvWmCrUCSbdunJsQsqeGFolLCrK
9InsRtYPyZb3cnpS4Vt7gJedaccazwxGQihHIYF7RnMlJivbiv70tRp5zK8OruxU
0YdJqamdy9h1Y9Rye1BKqTMpfjbQsFpelvZhOBqq25uLizoDHPk8Hd5xVQK2HhIW
P0okxMQLIQT3wIr934qKWQ==
`protect END_PROTECTED
