`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdgigC+RtjGK5T8iCh6B/j/+ai0NNJznaAv9IS1yV6KnzeJ/fJ5iUjPJVDSHndGD
CB0oLfPkU3fGo8er83Lu/4eMbTSwouwP7lJZrslDQZxlyyPK1Z01mKKJyNWD0FTd
K/KEN9TRIBKioqIUgqPq8GSHeYYLrrXhRw8C8tm6bvuF8rllo7DMdbVBPRGANLTj
8NtMQd3HfoYQxhq3OKwXKu4F0g0z7FmBFhxuSV1sELT0LYs53CN7hNbg7g0OS6tW
2kZoVk99sGAVaqj70EZ4cU4r9wsMTXN9hllgTldl59pk3OjhLLEIT2TeGzCnhsZo
OmVnrblh8VWjbUDLW12Q/w29vbycdz4POt50vyeyM2RplXY+dmera60ZYUtWAX+a
I1Ufbq5yAAamMfcuHW9tyyFB6P0F0hH5wJicHi3EWDHSYVH+Y9CzUToiLTClAdS4
yxWZ1nOQOawpeOTcsbqA3L92xNm/MEFYksiOYQez3j2zp8CVDQTZB9cnP6EhvWzQ
ZS4+b+wiYet4UdxwGGEmJC1kOCuwBMa8TcMTh968nqn9waLduJZGaqKiNDEmBGrn
IonR4srbwUQjnJ264Rb6hoeXyZUl6rRknPLhoagLLRMguEj8zU/hjGeoufgQKblz
1NcVdHFFNotlugEmzvjBHbBu/uT7+RfiyLc/skFOUZTN6rr++sO8sDEVeKVAaQce
DgJQOPp74aNtWLv79Svb61h0dfGXFbXmkIecXh0MoHzGWyqhNeX+FQmeyAtbBkKv
kxHGtwhQaVKi/wN+Ni1ZZJ/pCR2SCyoAvzmDs+x+QEzbokoik8GrbZHksU3dU1j0
9nG7+2DGgj7Wepqh3b2v+Gf0H2kfr1su1wKfImFWahM=
`protect END_PROTECTED
