`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2W3A+Nr843Vq+kP2iKYdDojBhmfNKcBLnFHG79FlLr5CPzk0OLdPEyhHKXONwcZ
Wx+JGX8h3QWHlauIFFnL2+MSHDA6wV9rWg6ty5pY2Ki1oGfe4udSzdiDe2y8wC9s
L6SFtESoYNqNb7azKDhK+MbmBW0VRVyETx0xhMLtkZeZ077XIVdfTB8YcX3R8NFm
ULkJizUKFREr4wEzK+zM7oUGgRBeSM0s/tV6p89v2NxQ9Wj35X5SjUU7KWKt2tjh
HwRebvIpaeV8j7HrS2CWEF1RKZiId+UREOdgsNawDWgGo+UHZqaRkiyXQfr9TpRT
LNGac8aD1Elf01d9hQGV+kciadZSfIAoEZvjSrlE/d50Tjt6b+xFN8a6+KwGnwY/
xujGfN8Hjx16x96iCxohi4JXihe8W0Q43rALl+O4Vptuyb/7/jbj2UYcnu+/tPxL
vfaY1KeT+tXsAOUdAHRARhxBvY5vkk//tkIeZZc8UifXdo5+dF8rE+ZCpiZZe6RI
AeK0O9r2Upr4Tjw56lbQ0f5sQHm7hGUsoDxslyILVpXzLjnTJC/k7+VMdR+hnKqc
WoLp2IQbg/vbYfAzX2/vzJmvK2rSpCHVDSTh1pAgWyjZRF9xqRo49X0NFoPoaVQB
UKtLC4m5GSvSZb55kf7Lbfov4EwtQJARj8YA4chZOVJjtaLbflP1sJr41OJuFhPp
g2LLB2t9tP19PRrQYHR67u4BEYdZVlakD8zo+Hu708acLY6QSb42hoZQfrvNO7gp
HwAEW9KSS9gAyUXuloI29xgvYE4AyuxVmXPd/jR6KFykE/1l5XWYvRAmTH4IRDbG
/tlq1I8WAt0Cw3v+GKWe0pJNFEP0eopmBETy9dq3pcdXtAz4ijJUWZg9Ol5Wpsf5
n/CVOLkTUAjMh7Ke9PNda++gadxVihg6vztrTbrTgXzb3c63wji45T9Idk/fhcbg
SRVn49NOZC5GTCvrCw+jm6C4gDBH7AZuzCZUr/WaUFIt2o5DMntjgWyC94ESLJoN
XVW76DLuLb2p9/PFBTv3MDnjMnzmC3nNJSbwTTfnzWV0d+RDF/zSNcDkwoyxsZ2z
PLoRrBGaQPYJ5iil2GTYPwe+X4Tvj4Sw812QHOQmjP9Aixt3DseTvbhhN8vve6x1
AhB5FAcQVRLMT0i7KkwMAzVPNCePZolBIOyWxxb3i9bl3aYUHhjbuwHM62bxhQhr
ZaQjSxOxCVO+p4AkpuCm+T6bcWkaGWH0p3j9X1JGrgb4UAU6Ar22yacSWkTmgNZR
B/lrbgvxgq5wAS0M50EE9/+sN7UpMikEe1w+3PVfxlUAhH77T+KIuNe14fmDpb8m
eWx0Lcz8iETXKEIGwF0p+q0KwpwE9XQT3Ok+Kb+XNVzO0gjJmDcdlfPZrsbkbyFK
Ikdgm/6+VOU8mBe2p6sUgrHwvcIRyAWW9ZqZFY6QF+kizEo2E5Loa24q+YOaUNqT
F6M2PnbSx4PcjqAb+fAPk+6tX1DT+k5Du4I4hOWA6Tk6dcs6vb37QJhJgF99yEdE
YtecI1wgG2kuDxdGp4ml32CYzkrY1f9LDvrdUw/dhKn/5eLraLiwkyohJcERsBiE
Zsy1nCwFD0z8vvIoQ7NG9JumJDy8ck+7pPOdStB2j4AmH9n4CqcAXU32t5Wf+Lkt
Fe+ajnWh0l9IrQCRuDBGWQ==
`protect END_PROTECTED
