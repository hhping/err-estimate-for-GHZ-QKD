`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpa6ymV/gVzEBcEOfskyGtSCSCJ7ML7VRDpwE9NsY/NdU+WWhVqtQql2wNTT58Nu
n7/biMezwz0KcaxBNiwvLIT5aLFgLkjqlyBP34B7mkXNdoLIzBeRj0w5BhsOMEh9
KwORX0ONEFpDxRsmo6HRkDvJht3vpnA/FZiljpjNYjiKDiisadu61vMcyqxdy20G
CCyWEO0l/sZjR4FDJ6XgMiZreW3FwpPbYqvITOoSrs23imcgueulMaXi/aQ4JzK7
l6z4FjTDuLYg5LVPv/6m7nSXjrWO7bcKWZZGvZHSwPSMhMxovykz6oOI87yaTFKa
RhK+6SIoUbUPNJ0IefKZxGNZp7PqY3AE4JmY9NY5XrE35ptexioJdcCaTxPnbMZI
0ULoKRIgmctyMIC4PCjiFhtMaVXzT+lQAXqqKPUgDmFhBEY00ryRA+ZYwyjsQdds
yA02gpHUYB7q1FlSEURZcudK5kSX3gyHp0x+opjyhC3PzPW6rV/ee8RUssUJ/JMq
GmsrUs0w7hk+XEbai5GX3YaM0vBk0y5jyQkZv3f9iKUxaK+wGUYZvtddpGrvM6cy
eC3dXPd//TNbgdG2FmZZWmhbBdgICFZ0p+Y5rU1jVySHI8MSSlJi2gKJs5wOwV20
BwpSo+kQZxHtgklc4T0gPr9dy3e0BGxnrxhf8Ydsgccw16q8L1ckcdNo4khrOHOE
BNNZpcGJinzINe63QUdAvRcIbhFwUEle/JkXVcbhAwYlS2WCiUNSnBoOZwRhpNqw
xftNbT6+k25foph947kbM+mJk8qf8dvntuyCD6aDqXJ2npFMvhrdQY/CaPjOg1Vw
l9fqLfZmY7lkvzeVlHQSIapOEVpJNlpcF8ArwWsYdoXYeVzEd51Cfo91iwTXgQg3
srX02lpB8j6RLCFRPATc1bot1JnTgQjtkIV/AL42fuU3kJQARLMqYPRxN2MOWwIQ
41HWa20oofru7zK2rsRkaf2H84M2dWMFB0snAylyFEHNJclXAbNgTzaTkHg9W61w
Cj3tpFkb2CR1PwpwSaY8mUFsIDU1wufaZfTdPAepRe+jQOPKtGo3cTvC15UlL+O7
44RiIoLgO1SCaM6815jQXtfzupK/fbcgyXLpNe1gGyE+y3hRPT21E613lRWLQkyv
HLgtSFnzateqzatxpZPED+4Oh86ON1GpiFpasbMI6y4wZq+C4DkGYtzYKDFmq4Km
KQWyUsoQwv5qIC/v+VbPmVtKrEvz+VRKRB62fwOHTV3Zsprgi8zYRanrD0R6ZrYP
lcplM/Yq9MJmC1r90eP7zgTshtB76PDckd7vSQuMkog7NzxPGkeUKVEHgtBvvMqw
gAJLCF9++EoJA1wrarmE1evcDs9CdXGenU9MeteG77zCdA/w5HVCQxDu7DgLGC7c
aIrNWWFgrxNTToMtsIMJ13S5dM5PZywW6rvREehQYC5cvQ52HsqkwRJH4Ra2sEQR
t4vCRbCZO102nLt+r6m+wsPbnsFJ0Y5woBKDtYTPCj2yaGUVil5TXg2Vm/KHmz4Y
MDE0EMUXgCwCAkrLjghbbIUlTq4kDtHgBAPepwyKW5XX+1fJox1zZsQ4doQZSiBN
s6pDr+W5biHugPdgcsdMt5QAfY0g+U0+oh4rcsmL+eMSZPG+kPc/sdlDnu4TgO5h
2CI2RC2e/lO5qpYRm7R/WGdaMIH+0ugIgowwp5gFsGL6H2nG9tDPgmPryYf08yqe
6EJgbdM4lq9OL+lMtFjxnnBe5CBlIEHoh6Izg8oPkLuW+r0lqj+lMO0GwU2Z7Xka
KipDKTg8sxIvqwrSpS0vYWLfoanFCHFlsqpxIxXaTp2UgGyAxRORPoIYdq+YeNBU
GoB/CGdApFf5CVudXxx8jUkh6BBghFAtCACPMsblmIUB+esnciEk7MzomvTx/opj
m15qnYcEHeG4/OSo0bxP/yOB1evxgMp4FjwY2WT7PbODql8zyi3ajqspoC+co5Xg
2BUuAeoRENoeJtAgtbM1sftZpUxUm2hzLPqjC7yZb/bY93RbM5OQCMdHaDxRVJsT
s2qybKlM0F5alyQ3d+R3eMWu+9iT/uM9uVlA3Zxx5LHX0ab4JdXcq7YRPgqEVwlS
aNAyBNe+pquL/NltQcOoxuqQyFcl15F7zYD2Epjzfa0dRSOkLSDTS6IqYNVvUSje
MEcrl8CF41YmAzz4ArTQ4WXx2fcdiclrMi00iNzvLrKrNeFLWFmhwo0I4iCXV7yZ
2zWfUCH/8GS0nSrv/Q7bP4EMumg9FHnPgrG3kIEUzO4w4mo9l5C37QC5wkS4MB+R
w5dE3EBq8jz8XBX8as/kVvOc5SnUTmihDPNQR5Fm96mjwZV49NnwlClJeB0zD8sG
gcpeYK+NJHgNAKCKfK3kq3gskxYtdsfckdiB6cuftpHyYzwfXtrr/llWARH1rS7W
ADucHnqgkH+is3nr7kLTeV2UiUeBhKWFB9lKasiOSNW47/IHmR9fbwOqX4AOUias
dE6rvFSqU2eDeW9kwJrdk6J3deBOIY3ebejhg0UeC0KfWKEn3Q7I8NX+1wz4g1xg
SY+kZhRbpQbdGWCc6NoGMd78xCAnRlVIGfmh4QrDR34IYKGsQSqAlcWXLLW2f+He
G7K6YOSA0DKuSzwV8CP6NUieHmZ9n32lN5nyXJDJg49+4YVBPFVTIxnC4vNZKepp
EpLTb1nnDdEV69MJT9raJ3BbMpTWQUQM4bQrTpaU1tyKJBGmN/RMkZQkp10G009Y
JmIeCMwD8SfceSkCvoqqP4xUsaIJLJ8vM0W5AdwIBz+5M8X+UC4NTHr688hgxqvb
XEPBJwgJdvAw0txSHyzggkBQIn1En7qLZhdOXM9M0G+3eKsuv6S+3LVWigU2BqVf
LeaUuoUDc31ZHVjVrQwgeHFbptcqVXT9UA1pJdv9jymsEtTsiDeqVJ0vOHnHjOtu
QXCqPLjJAzyUMYj13HWetYczmKRZ1gD3NwG875kpYsD/0t76qEUVuXnbvaijz0sU
C3st5qJmGlQ0izO/zzc9X99HbMk1aYgJK1NGilA+s7Kcm1EhqQpZkMeYfbb5G+4a
RhJntp+pjQ3K0SYBkovd9jo00jsFyXy8PoaHn71WiOSP4kUQjvrzWQULk5JM+6lc
GsN5VkQFGb4qLrl3z4uDsNTeWDzSlQ+Vh876xPDvOSNSv9+WN55VibHK8ekGRr5m
B4QsQRDPipN7wlL0oEmWnxQ/36c7R5DSjd/IRjNVhlqq8wEKgJcungLEilpIKWiV
GRMjXqs9iyiM7YqFRUVXK2vxTIbzaYvoVEbyxmoZZSU64It6mZHSHU/vPGxRgX6y
RYo4/Ko9ZRNelvC7jDC4Dma+rqLqY+ND/QowF4kXfrF16lgsuIYd+F5B4vUUiU8A
zrqFNrxCtls9q2BYjluyUWal6VOIvKuYHm4H3ajKY32dTUfK25V1TxuP2hYUZmMl
Zd8wAJDBqSIhLVRjx+FpYYzdA8Su5Z0g1XAGUQPR73WEyLHPCGayuN8yGyhU7QV+
qD+dr2pFRTSSSZ1DNKmwGZ3GjF+YUHOppqzFfbReG1sv4bcfboyMOUBwQXVXareq
NzMLOpZ93IQWZTMmRglx5Mhv7g1SaE6/2OK0xd7Zxj453wRJV92+CIXNWdCPNHzs
5A7K8e3NbC3s19JonjkKjiEAEFgX9/qfoOEN0mlVX5eUpVVAsk3dvW8zcQ/7ZmRD
+LXmg8C50wyK87t+6UgnyGv+2ROWOMAYi9+pa+ju1oqBUtLLhHpiVZ8Pvux2aeiB
o56icpBWdwFNM1cYBNolW3V7oQQsEfQJCX7J+0yqnKRn5E/59xLIEXovAIOCIOYn
zQ2/rmqsMHYNrjVUoUIQJp29/akF72+0kcU/OLsjDRmBlLFVcMKSjgUGupeX7CSf
pB/MsBXIPTCH2pYXy+TEfyr9+t6PaS1IzYCMcMUhCKmlFk+SKNc2EKJhTOioSsYy
qF+CRYap9YN/UtelwWXzFuE+z8l5XX5f1MfEguFBxZOmPdak7Q8WHoGqQnbKpVgm
539n8/bxmYeD0pLjUgQgl/mBwW+GcUIuRC/ZTuCBpaTKOmUY+txxoGeBR2ARPZra
rSKXkykzarrkCKoYz2m+XHobL8VnvhfxxyJH5LHt2PqnaeW9+gHoltGqQhiLJ3ng
PmrJ+abL60nw7T0XIjpYXqWbtAmfSTyxwXhPbs0oTt1Ps5TWZNZ6eaujRj2/uQJt
k+TmCVSF6L+dB2BYna+2N9cZyxTdQ37q0nCZzaZj8dg38lFKcCuhzzP02gcoRpHx
EnaWRDUqYR3QJfYBnHrk3SK6V4RIbFs/1CizW//frYnCliTZmgyGIs0jLA6keVeI
7xkqEijF1QQJr6sOtfBa9la1GAlzJo+EhCXeQTmRrUKa0PAI9Srzk28Xyij2Q1GW
JQq4KAz8hQ2kowjyER2YRSCMIZSoyM9sSBnWCW8P5xBaPFK72JF/XfSK83dvh2ND
alkhecl6dXFURaijMxdKE63S8377NmWdW5StqqwGOTBwaadLSf5wqTyZupn8i0uH
qdek59dl6TJ85JMwVy1TY05nOQCCaFBdYtEOBv83bmujE6tav7YFiWKL669MaMSN
/gBGcF9yEM3iGfqsUdU42uLSXoPWdJR23FK2QeQI1HvvjrBkgtZ2CUvZ6QQgS6TU
w63+tQRT0XeQDCK3jdvJZpleXp73TmNRJAv8+fInhrU6Sw9HHM2QOgCN1OI1u8Dc
Xv+DWJlJtzaCRcIh6NLz8H75UhIIvD50goHPM/rH+ais2Qwv6qLLzbqfuTJ3kFEY
hzOsX9MpKctB5YsgsCsogAbUY0FBrZvGaZZ/XXYUWWgyFtFlFmZGFyUFQRn0a9sI
Hfrej3RcC2iDqn4fxK/LqkEsSCHBT4xPDODZS599rWEiv0E/npH6MKaahKLdinCx
iILwi94dmFLwh8lBkdiBxJXj0f4zzawqwaM3PAV4ZQKEuMwCfIqCq3DhSkbb8A8S
hYvqpvUvs/Qk7vct8sxrnvH3Qjg5Jnfaq/NbLsiBYBrVoRuM/8yhpWP+gxb92sN8
jBm3dSP3FwiVnRxuy/mdzLnAJHE7DuhMSRAYTumvn4lKJabWT9eAC6FWAQg5NRmR
uxtUGktmOh1NpV/8Dqc7/UOVIbsHBr/qNNbf1zypYwLxZV5SaFIjsGvKFyuG52Jx
DYHffr9Rcf1G49oxBACp8F+mJtsU8ZgvDX8PwXuZMN/N7IfeAnjvgoGpXKXunDXF
slvxK7m2VfTm2FZEsZ99eFWA0CO135kZ0gDtCsmox5vhiJKAm+8OpIxqojZ+T51a
ywrYc/gt9Q2Vv+wBgs2HmlIMpHPJRE93SXvFwzKXc9OYk4VBpMSIrUJJIWCmL4tF
lXSc9VhuJ9VaJzfe0ATeH6yMl8VY9ff0gb4ggB4UQYcyW931KDpkUqomtnWiC7Gh
/9jL0bu87cZ3+ZtWVqmf8SYP9Oh65mQK0HVjKnTWNO5Hfnj7kFv4OqD6hJ6sSmIT
d7ZagqTHmwwx8/WA28i25i1iwiCrzvJYnJBRVvHBfd/m1DijFz8nn+394uFb7Mpw
fs1M+eSA/yU41F58hcNbOluwXbQ8xswDLW8tUFC4Xrh55xR3etvxf+KweS6CNwuU
FvS5JnUF52F4927mH5jj0SNwM0gEyht+cvODStBSUVCNPEKmHExWYLsD0Jk8yC2o
5hw0p+St6LmU2bUSUnda1XLMAx8sbQjhV/tBNFc0q0z23LdpyxqhEM4mZsHxBMhK
kZNYJJUr3QfjFYZWG/lj0NksBZghqPuRYaN4IjyqM/cbvrcMmXrgsTYyNnQWSdy0
rdnphkQrBLnx9SfxgGI8ilRrLZm9eHo0uhlIZ8PxN4/sHp3K06Xq4Rm1C8E1QAj9
Q2B/PiAFDRKuFfGnrwQxMLQpHV6Yh3TnBwNjwwaZC/3DhWZf5o9nIEPDO4+pziFC
HlTQGd6gpv1ipyQCvTuPabmMPUbjFiGTEg8S2ZbCZQBcpVmrfQOHRs0+xPbRCk8C
miz7xezi3ch7WdA28StvO1r2bS2KT5SbQrXV3UBXk9uNnJC/Q+3yOUokcJNVW27e
QQ/87PolrbOt69VfDJgn55FwSLYoDifLv2/B0T0f58uhIXmJYJSm6Fr8SQEabUIB
WLKlrKvT4Pf/Rg9NxOS0oM6ByineSbUMaW7HZgIaRHHvkVB7n+YaTGytU0a43CBt
fEYIhtLisBpvW0E7g/kyBeSITYLj4/vlGm1KVFz0pJe5ZEKDY+TJfrBlx0DmqsPN
TTEZ3reTcOaN980Yrr4TlgXixiw8YMzg4yThrtWWwBrVko7CxTlP/4KcaPK+x/mo
pGjHnGwzcUGcYI6suZ8t9+gIiAGuUX0tx2PtpSyz/dBNowKDcFT2cLLe1XKdYb2W
bKkPGWkMQgG2h7XCW9qrezZZqXAQ1VQ5o49x2Q3JZKGuY7zkzMROBgkPGhhX3nTL
CrAjvzq0hbH6Ol9OC17uQ5sfPnMbHKkNCbsjm0ZO4saRu4XR/9Zg0R0BPp42lIYu
38lbcvLs2pin4OucbJ15bV/DdjzquQB//y0oISD4x2GL/iIRLk1OJ3jbhjKBZpjW
2A1q2mWpx+diLM+Mit86REgOwrB+9sYcDJm1YEqsEwgCSK2v/ExSk/+XthFiu75d
H/FH8lBjNwvjbryjGTDfbgOQi50zz8ih22O/9bPPc6BSc9v0vfSZT0P6epX4Bdi9
ME9wVTSdTPLp0vzOrUzl4gyHMmj+RtvgDvNd5/QubghsPL7mAgsUq7XVPGculXyY
DfDM5X4Nn9aulDLy31tFok4ETt9qu1SyToh/Z8U12RQ1QCZjeOl9UaOlbpz+YPX1
g9UpxSwdnTV6A2aNUF6N5fZJAelzPzCuml3e3U1XohEYrW5PmHTfbX1eRj9ZwJ2S
FzAuFFqwYXXZJF6MHR+VS2suAok5xsgwaWTRwq9bckfPAtsySreYXNd8tHObNRp7
8J75JvZvkFJ1m8KQhc8+gW17jxPEv8iW02lPmzaI9mM6QpagfCyKdgvKzx5YvEVE
XfouBA8tapDQsw/NzwCDn5kZtDRkaCMJf/LrYeorNp+iis6vdJzBeXLMdhGD8j2m
CIkQkX+k6y5ffq6OjIV4+vHaeeYEJ9ViQnPXW6mCI0yTJfIBmSktWSX1D2jLX2Tx
M53Zzzbj+VEukiVsR5datnG/1EaAqMB/O9Zpxm74wM2dMmbS7Thv3YPxPBCDVJ5e
XSfJVGBd9+BmpAZ4KEFw2/v7+E2aunOgTtLXZO4/mMPgdBV1jhj+HfFtBlmeHhz6
HPapaUAoQXrY2AJqirsCAW3dYBdeOmeihoX3YEvoQRYKpwqVpcGIl66jC9a+IceG
wKpqxn/obsk7cRRR9FqW19qyLE3H7ETU11Y7GGmhTR3kmdmVqKVR7yoOJTc1KKE/
b96pIZYi5Bzq1Vx2568TSqENKg9EEQdlrG6kE1CKeT6wvcP3kySJC/BUVVK5xbP/
o8SPwX2cZ+gRVZdMX9fm3LZAT2zhsG1+F99ZU3vSMwCuIRTszFpBblN5/6jAcu2K
c8avLLE0sUlbAi1DphRt/W5VwsqsPvCDay5tDLxdLZjo2DND5KAHQIpF7r99v+hU
qnR9e+rNJx+BKgwrG8Ov1MLMjEgAoiDyPjETZvnVK5HqZwijdriGNJyiGJL6Zl/k
dctizklwRVm/yOzsnvLO0jQar3tleAwWd3pF9kZo+SctwY01ysXXxZgUi3S9CqQ5
SNuNJgG7wnCOOsa+MIfQYvYvR4oadT5CbbQcjSPbJBpMu+hp3HztLClXyhXIrgMd
TRZH4J3gfpb6kc+gjne8ve2JmTpAMKZl8P9vf5nMsaVUXb8yncJ6Q/h7BQes1hGY
SsQ2z5vJQ/KtQAxZliRwb5pomDihowfBZdRQugM3U6eqkRe4EpcBQMsRTwb0o04c
58b7G8PrZZgYOLL/X9e8/0m7VxSP1xwxHfLnuj9byTW8rESCjpKYStcRAf/QwXMA
pYN7RZK7GJ48FQVE0acNL2rx6FCmbB22dd+PlnISJF6OxdK5Bnc9bWYJcDHYeo5Q
jbDKmO6OLqcRIjM1mzngYUZQQesJgVkEDehuuzH5hA4WF/Ja7ViMJK1baE94qhjM
EJMwBKo2j07hztwo17iRLZM7xCmIsf9cPwompPhO7JxVimyrlEJqqJw18BXL31NN
RRPEAgtuB6UFLWo4S7DKjIIqb809IuGl+xZxQ13ClvlvVTdA66nq4lxeA7fXCVp2
Gbn+7tZCudRFDFKX00SBxjO0wVLjind1+WKHbcoCzlrBx3gHLJvXRSTiqy6yyi3A
HWBSJZ7uiZtjTBwJVIWLvcJtEd8YOv/k2ZLdQQoZZvDToT2bc5TX0g5N6OhyF+TS
9iZKAI/wE9PO9X3Up6i8BKFSDVfRW9LC7zHRebwEcu57hrp8YXFm2MzKW0pYUS7k
cS35XleB0UvZWDqo90lsVu3BTLVCd75MuCbXWek2Fw+Xmb5vt/9KvQstKyX2UXso
yl7RieEJKVgpdLtNDXNHAtUIaulX03COQIBoFuQ+x+2wDUBe3cpr7o0qShMezs44
jcch6PuPR3Ma0TNwrObLy+fBhwmYTzEgg0OJAS6geRbWITHZmMw8+Jf67OW73329
HUSdeblGRG6zJfe+0BhRahFl+rK99a5RP69/46rzFKL2rYZzAldzBc45M9YqeiCL
iPjK4CNGr2qQGivy6ms+T2lJry2XHIjqNx08SGLkphI3EevY70AJHGMyQMDxtK67
wc+4dP0vxxvqAmk1kaBjLt4mYCzmlJy8cDPJXOVcCN4rmsiZ6KLVcGrab4IE0frI
nUA0DW0QnhMhYn14RE+ZHr/pvDTDNKi5ZWLOyYMWjAdTNGzAbw5VW6dYP5YmsqFR
MN4ms9kI/hPliXCvkR8CfDvKCXMFWUNCxlMZ1luPU87m9HiuNdkYrzU4oqLmrfF4
42yPVJcXuBUvMAwd2j50eLtAK8zWHQFQq6Icj149egkWm9f86qapteU2ID7cfZ+H
vkTwxe5dY6kfmHVAE7gyxPh5QF0v1k2H/1dPv6DnZWErbEfXT83rgeKw4cxBknT/
EEzFaXXQZh89ThZL6c0Tbv4UMLVLK8Uy78wk0iPoN/zpSGlWk01amB9NlHYOCRtx
N2ze+UDA4ao6Tjo/KEiP9QyqTGMBCG0qoHNXJBIU9m7BYSebo7A+gvKxHPL/IOpz
LSPttFLL4yixywdz0MaCRn+028wPsYx5LegtstpXDZsoNK0eNC69dugEWxa++OMY
Sk64tSyPHqkG7R4BW5pH1I0faWpJyGHUYzrIFvJ5YMRoQ/HLJUuxZa1RU0j4q2IA
afu64Hn257g1D/0qBPy/eljWi+gNAKIvbyGnvFFsHPYsfTerqFIpgq8zJ04VTZo8
g4mI8Xe3inwfB/oJ9ieJdWpalbS/WHENy5Z5rU94mgRrdrapyBjvLBnAcpcTVFV/
O29ig5wVxAxQhNg3wDSx4lFopfr60cG3fFNKaCECYFeNCzW7CL19cwk9u82h2pZm
psv0JkrP9NuKz42cFanYEvD8jerfyKZzjg4YowHBUiVY6LHKYAovH7OcuZrnqRKX
0CJlVWyUMIWyCfbIca1mYV/+nHAbC0Ic8dtvsg5tQXn62FXaXQ/1JvFAApNixwHS
a0bj6if2443PyqzgFa6nTka9nP6mc1ZKy3UHqMueLAvE96ogKucQ0qI5CFvXyt4W
+ou2ArAkvlsEvwgc4uzEptzS+9OaKluAsrXRu7ZpEmQweIVFIIqMS8U2bXRRkt8C
WWANzmIKFvB12WVLqRZzLWrzYDEykdtLw+kX0EJqhZCojaQGprw088+gjxpyKpAn
mo0WkcUP3v4xz4FRIjsaQfo+QY/DFdrDtuArKE99LshW/G7ca/DzOAMmdi1sGkVK
5D1xPq0xx0zVGmBpsPdWGMVdLdDHgKNQ0s5T82gvgVLggDH2hRwXh0gBJ+KDvAOl
Vzaekg4/ff46jVGWhUolmHXfurF8lZFI6cevEqSmguESFHjIIT5IknwL9W1UCpzz
ijIC2quNd+2Kr3sDEL5O20Uwe+hl/aOvTiA5/NSk4WTE04+hT39joJSBNWiX5r4x
j96GHCx8Kv2cZCM0YrGij2Mc96NZHMnt9nXXPj61c5ulXL10t6uYlf5yyQtErg87
LdwdZI/wgTok2ku9SMb9NL0tg2u9Y7OPjWoN7vSRazn5vLebRHJS65DfCd/xIsSL
pScd+JdvI3YkcYa1Nh9GJuyKw0gO3MwjktuQQrA+pNKF97ARqzMwy5hKhGAS2Mxa
t62OngblorcDMXORrfhGSPpI6umywqJpF6wDbSqmJOdIqDcALKVDx20ZDC3WT4xF
ScgwgtyF3r93vPiwJwppuZ1GUqhgQQVf3UYIngvWDGPEKndE8vufyO0KGBRWrHxV
C56m+3KIj2FXuiLRRSErveVevDz6sgSKv468+quprFdwneklLcXMjpVwJiLc7B9P
FlPjxc2z7+VE88fQ6x+XuXGy07pqLDcN3zFMyKFpK2dI+7yalLkUUt6kZO0C6Q02
pfE1jmL1zzSsEtHT3Ybwb1ZyaXxEw9aWSZheGpTnjfn5Ee8QGnaVFbiTpPN1WUIi
/CkrcJJX+hfJgUCYjCmfrV25sm3wpPc9ZFOepT91HYd+d5mIE6Be0ydz8wL8o+ca
Qm68HEyWgaP8Py6qzpdkgsc+mdNBXIkx7ktwt165Bt1sgbHn0g42smGtwog7OcOM
l+s/p4zbTf7i5+o1ByS+RaaiB7U+ve9SrKWpeGaGq1Psp49Cq+GdyZZsYnNfbn0j
VsJnKWGQtZo2B1zGzPtI1eUHtVTp+RH8EBhsTEXO8iiSgcbUllqncuLa5r8Twspe
Mcbc8RN870X11vIGnfe9+ipkU1r1c0JIjgaEjUpy0RYAPpQVtJclklrhYbsVERjh
lTvrQ8/b7HFlbnf9nxAlHDSTj4zusF376jYRm/KXO4HnlVqbVwA890pDRjeY4aLK
WuqZCcXDgoT8iLmz0bFRTiwyl68zQrI7hW47RcHPM4UZEfLDsLNQj+/HOph/wMUP
FeJGA39xCU9kfmqrzXQSHVVQby+FgZ1k8tAskdbxWemAORhLTVa44iRCUCJmhH59
ywFTyICe6kDK0fmJqjS/ieF7evoVs1DCwiMuJk+NRYLmNyTPyZCW09vLCNJiPs6A
d+iRT6jd074HfH5tqdqGISeX5uYTRjKR//Gr25PB6lEy0o0H3m4YWw9IPY1tt/ov
8PS1Q9myr/XKveKf0UKiB1awFpgfP0wlVcInvdgjjiQ3rK8EmXvJTb1KoPjejXnm
KVWv32Fim9v8ReooTO6M2hI4LKMK0siMJqsuOn1t2opW2TclMnnRfEdhha5wgqNd
SS8stS05IHxdvBsCXtoIsmSrPV3O5jLHt3PcZ5B2xAkH2LQ8+xmgn8EJmEGmIGV+
1drBvF/+64bFlsjjXcVDRB0fTt/oF709m3c9KbAbNfzGxuWjjZLTpw4ChFtVO+ZA
jdcYamVQnKPzGA4g5oB08Wmt4sgnVOCnzrPhVWfZfgm3uHyBSgevMY5d3t3+LKt7
bOwEy0J2mdN1mYXy7b6q3pzemwdj0rFXWnOreo4YD6Rt8NpV5K2l0eup1yLm82cp
o1DmPqcQKGVEQB39W1dMMDAipKHxBpzRwO87p4s38zZxdwBCMnVv6ZbcOy89Vnqb
vMdSvKGCHGM5XHRfuJptg0nCOKQnmvoGcigHG+ORPlbOlRH4+h7ZMihMBh71cBqA
wBfvnxTx7WxaDok5UJmtagkrt6G1jjnAeEn+wl3gZOgdHh98Y+lfmTV9EH1rhGW4
ot4eNya/JsrdunE5NAYhMokwJqy4gF3HpTKOyPs6BPB7Modekl2SwWFM8YILTWUe
Gv+3s/POuyJPrTAG/K2TcRfRcwbSYQWazuqEvnOIqenkNVAlkWGtkoVJ6Ei/v+CZ
PP6wh6mwA40097bb+AyOgTITC31ztMkriaRtxyQccPH6pS5kPc3nE6ls3EQ1nYEq
xf7/dpRhM9/Vd1lnQymCFEgzxO4wNpOpHxkoefuhN+w8R/PaDiZ8snWBJVGzQCRy
zN+0xw+ZZ3PpW1/Qyc3xZiOtQJI49u2Woe00X+oN8Kbo87Kc31PZydKzTWSYOCO6
fGDY4mkXdktNM2u4PLzv9AhDu11LQWwp+jOgIo3T+0BYBpjxojfERz4zrL1SjjLE
FXO1YJ7gMJsRBrMP05iujfoYVqg5XbiPIiPBf9/ETGU6ns/xyBj4Coyxo+SFErPZ
c0N15SzjQ6wuJm3KkHh2iCT8L35+/kKc+sanaITikaQqi16ms0nvsM5REovhDGHr
Y/0H9lYTz+sL2hsoEd5RnD4/+JHdi/7zCoI7zaMj1ESUEIYnOi5LUAhUfvATOwNu
ROg3BG8/gxM9g81x1Vnj6DwdPo/9tDwz7+hmCc/piVmjqP0hMbzi+jNBKtomGeDG
NrKUGcNtieuko+/ni7M8vGIwTqoBGdzXnG1+UhpmcFjQqu7Z542yTY0crOAB5bE1
+DBy2JZyNbWgPjE4wT0R23xijeASfseG0V2PmtoRVCqg36PdsJgGX17GBTwLnLFi
8bB4pROU54RSyP8T/1g5+7679dc+4IGfeL88fcd4Y5x+IpMGqdcz5CplgZcGITgg
AFmgyNdWs8oHDRkzeYXKfP0hRcYPD1oyu3ydVxP50WMMCMJt8zp0XPtkEFK08HHU
gq6ZL8FfxTczeBW72zCd3VKZKBFY0gVVsRPbrjFHGznGbTbrwInS04+iAcXTNlbj
bS8aM1YzIkDOmueHi0MZDSDTwK4+mtrHS/+Y8Rok2Wwy5IdEQFoSFvyDi+DePEpY
il7kb+4wVzp02AWP5ixnzB/SJ4ptbRGjONqQ5gNIH+JYSoVl3v1agsRU45emf08B
AOuHgEa3fcffSU6Qiyf6c00ylXVaWgoy//f55M82mmgbCeiIaHZPVR+HMltcKKRs
I2EpwQHkixWu0dehjlS5Fcwml+p+hZg/dQXTpkGh5tg1Og9qJ9fVl/vvMZsl7glA
bYR9nhWBQqTDpLdatrDm6Gd+RGxb3DY4l7nWeR5RfeEDvqp+sNJO62q2T6OJVV75
HoLLqMIo0JtNubM2gxpxwK0tpAj6ATPIL/+Y6NQHqZ408r/Xi8ZKTe3shDahsfCB
ESUDNUAKWhogtqiUfv720vRnsaDyy7UISO+oq7fl6TsZNMv3jW4JK0pBwDzvO72F
s+kw5FDIKYE9cLfLElNReEx9vNapXzuc5v/4/D+C4QXgpybSrK3N0HBM/GH/fdF0
hZ0+LhpYpVqchpWwwU61efq6zxn7Zcb5BR/XRGtf2o1giTT1FYrI7H2dtfLWPMNp
eYLAtLfPv4JMaWTZja24wU6GDTuCNFzehhpu/ngW/iUWApCqlN6sXp3iWKr25pwL
4V39C9TU6GDVtyEN/SzHHHS4PrHJG09P9QIzVjVCEOTfmVnsSnN8VOKs5YZoT3YC
UcraXhwGgWFkWQ+eYgkUl+KhP4Eg8hc7thQn/78cXZjwVt16CDZ+DSCUJC0JtcyH
Fk6PPuKxNw7qPoubRiASSFNQC2WgnOgVJeWbXxgddEiaCPaekrc3luA5cVr24A+R
4UPwoC89uhyMPKU3Y9sPeFOIlTuOA8HMkenDN2Bk6d8vSnkLa1tcXamqSL/DGBkK
bFv3Nq4dlBPGz9djRsBpdmyA+yQajfGFwS+0eWk/3USE8jTOaL8Wk+qFUR98Md9M
YWHR7o4OA5uXFRQq4dSsnPK8gf74fgmSmmU5y0zcJQI/lM0Gg3Y9YCfpS759QPgW
+66/h3uHAlQu2FJAVLhNNNjxJQVg9iTEJPz2VG+xNACwclxRUH7g62rd6K1NNIDh
`protect END_PROTECTED
