`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3REybm++Obs826659Gi2QMve9RH1kXU8gNEJpHcoVDToesopoOgGy9rffqqVZPEF
KQ42Igu1aCjhDGQDHoM+03LM9qCgicNGqp/PrOBXMSVhkej0M1D4+1td6lrTqdfp
KlTR0xnSl5ow1lYkS9zkag4+Jdf5xnTzCgV+BagvxJvDnq4fj9vLxqvcFyXeAamx
kXIxgt3U7jwUHSIFZ128S0Kt8JTaMCpnMMcDlH11lKdKA/aCBTVKBtRTTSQIDksg
jYwpt2c8XrCveFCaGMcGqd9jFyQNIIL14WC3x61Qiof/cNUcGG/+sZi7plizHLsd
d8Nv8haEE9Lfaqi6MsLfkaiwOjncdNl0kIiRMZy/n3J5q4XukrrweFhXi9VE2ek/
/ZEigyh94QwO84HWXcKd1/s1UIzyBxVPjCcdON67aDOnSUDe4soMp5QUO9Oip6Ty
kPLRlZ3nckmhdjPQFzfyF0t9Rc6p/nOzCQz6agh+7FTWhMIG25Oo7vbv2alg0HcS
q3XiH86vEjEVwsV5dMqMgUSKwOi5Us10iFQ6uhzOLj3d6LlcTH+nm8pFnicdTO7I
u4icxI/QCYX2dmgcMZ+KZFb5++Ff5Ba8e24F1DVvY43kzbwVA2bEqHVsedSneo2k
BmwEsXa3QrBdL/hRQiTl1DLvb0Hrdg+xxgcb7XUWjj8vs0aip8F5m6tX0V9cyM+1
HG5nwQheTUkR0qyBXlKo2ViInlaKXvjxEjnNkEtbI6xOV55iiTkcwdJHe0Y2EGhM
aE2vq9b0nfrT+YZHVUn5yQZBbMXkCbVkRmPSyxWR72SGt4XiLXeyEuftJS7ffZFm
nG2WE4oEtq3bPuXyCP5JVOsVksbjawCgr0ftlppF7w5OCtH+baEUFCbZcLHOcPkV
B8/DvSWphSEwgE+jKTrT9e2rv/XBS+3ro3L2bl0E4mG1BVkWA/b9+4ICts2AQPlO
oQTm9xL20PvOJlklSVMXCFKM0NULDfjDJfWmE43mgt7c2lR0TZDAy8x2INha8eqN
HfqIUo79H4NsMirLo9szVg/goaLdbQgZFSzQTBH5QyD33IYcZzTr20oI42w2/oL0
liPi0CASkm/KUrdfqBWeELBO1EaNSXZF+UgrFyHu+ohnBTz4sEcATjqUp94m1NUZ
sckECVsd1amS2kLqYNPixLnNX2yaGsjfNsVKYCadWBjdZx0VO18WcR8rrsBPLJ/T
9ryMgSLnmbz4D23BHfmU45U+zZaZaCOaG9z2a3or9ybbBm+CuVDD9oxyIqNGu1uV
d+il2myWFcw5A4T3emKt7y2p2v6Bq+tF6Oj4ogPXkbcq7ZZE2rBe6E3lqcv7sIle
P7/UZjLQF/oCmaeHlUHN/YzulpuxN/mBKfKWd2A2vtEcI3US9HgAxijjdUJJESFP
H3o3mV2nM569g0NY4pIlfHQRu1WYQERTqtqtNnm6Vp4nMwFClnSN32hNH25/ONSI
VY67qI+LuzIUYuEkq7c34dDmYU5OQBicj3ADrj2IRRZ46B7jyYDePnMk2j/+r34Q
Apj9YvVEh2chxk1GpPMsS+oIcMqAhvovKvVzj9bT5vcdbupAy5+JTCQP93kc0GYB
RAYrzOkGCSFshU+FenegGESSAMK/fLtOaTntklK3IWXaS9sLgdwRZkkWHfbRa+Cm
SmNFOC3k7pm1L18tNs3PS0lx8Uk5O0ddxlaK2uKGhAhmPsHxhut+7oEtFrQZEWRQ
Z02utPFqQy6CAGHikBDcEvcC2sq1QAb1BFpyUMgPgMSgMgFnCjzdc9hwWWLm/99k
3atkVLDgujeWMYg4lPDs/M8gbI2/bBQBJaogzt8tGVGrxZqaWm65T7chcivVBW5e
D7Ds3xeaFtCzqFaNPPRwVmNqRTGuM1r/toKfhsWh3sp5IJkjhow7JWo0iayodvoV
Z+GTCQAO/t2ty6QphVCjqR/lm9RgG56Ky2aAiTZRKImWntw1RuZkvAzNhpbA6VT1
LBfkd6+eI+TuC2xcwAZUaW9tEc16wtgRAmy/Gr+XAf4yhJvjEpQF2HL8+vY5izhh
6A+cKY1Vjh6SN/vbOBSqUoLkIFZ1sEgHYeuRyV9Vno2fBMR+fO4ItgUFh6pCX+D0
pPQ3qGyyLV1mzmUAQkA3sCZnRMTd8uLuE84diJSW9L2vEs0DP1/s8xxzB1bH0mr4
bfdu9fhOefvoalgD9UU7J+Q2MAPt0WmtmIe9Skg1xD/K5LnALU61SaB3MCg0DO2P
70p06EX6S1jD2rJHiHzhIQNvGhM30B1wyMKFXz0ql3uJSfyLeJhdqhdH1ME9GVVV
cZ9ENRYct1wzsBCtn7pTe0WLmPpP0+DRYVnHlhM0YpzLqDeMdckVTivZwh9HRkJ0
6R7BrA6uQgqzKlDiGXTK9mvdv3pTU5nWUKv7ApD2HwBOCUzXsResTKd3FMn41JMV
0vZ5LeOAA4zK9F+urpV6lswJf6bAvks0JTEYL0gQzBPLemVgdS9uidJVT8A1YEO7
cWBPQD2ySS1AsbCf/HHAElFyzvRcypgzRsrkA4Rw42YqFCkqalO4UYD+qZ20C6h1
YbzKpHElq7TvcKuexpLD/Jy5hubTpWNslYxIwvFgSaX/OEuuRYX1OnD089Xm49rB
jKbGriTXiIcJ57kH3C+woI1r81Q/Tp0juj4TMQ+eydzEnYNiOta0jzzIHcMx09GJ
zPO0FuW87izdm0Gvm7Cp/PQN4IhsfLfE0Lls9kxsAUeqC+CWHA8vtjKhq+WmD3Ep
tlfaA8eKIrbKjnwyZJ2YDsAD4SfEBUogKrSythnKm6TR9C4alBTi6/PHuNRJO+WN
gxgXHHes3YwBsowDdIdDn4JWh9oxAgfQ7f0AxvKkO/mtfOZy21PsI6jaUYMrzJ5l
0sHYv21W+khFyIOaOwGkWJzFBdhya1KGst9mbxd61Q6OgWMr6WqCvllSbPEzv6pT
VRSABW+cbDqgpayiskStfYWt3RUZI1ZdMyUqhzXfyLjA3pEpp1cL6JDR+uLy51TO
TBSUHYfZBGburXULUZzKOGD79OZmm7/SS6dRwiAqkS490BQM1G9nzx+YMHl8J89n
U9QPM/RlIbm9Oi4y1jghVGc5FoDPjot8cvedzbCk35QG4HodInhxxU4carAjTIw8
ixXvIM/czWRT2sFRaP+6jx5E7ZfO38cIZ81goWwnVbh4pNn2R/N/NCKwyeXJYqEs
2+/S195CTTf7K27T9vLF7LEiRWzKI8N370VUJpnJOVFAAJemLrL0pQUY05mptvWG
Pu1+w5cqubsZiKBLNrJN0svgBMcIR+HDsqEVqqZeDvPwJsNMC4unstGxIPciINSV
TNwioTPeF0y0yqRwyciOprgMjDdvPE2JrrR3xZqLFlFtZDpHLijqt9Fb0IzhwntR
IRKdKyHp+J7/bPKBPBzxff+KiZdJXw/ysouztRl6BkMgcR71fDfoachBWuW0mb2z
Z3PaHCPTOBmtRmvee3pKM3Wmy5tKyWnpdpamIGvezMIWCn6sLK5VQQV9dhkfLRT0
q0HHZObCVFMa1MlLfY+6dJNW82+Ykr4yGCdgxAg9Aqp/PMjoWviaBKdgYE76qsGR
FwrRXUOZANN1qSb9FljtxB3RftjXgTHmcYCMws5vZBvJkW3HnfXgG/rQnIMPhW7d
XGr6dyheeE/KNTJAJyVPS9iv3Xub+8Vvxr5CMiR9T6HcCTTTuLMt1iY2v2Q0zXzY
dW6u62hHS2ifiTqJ6HGs3QpvT1VbgqG0WIUr+6CP1iJhPJ5KCmYGc1fE0P95CtTT
Gs6qs/fZFzJPjm23hCFBVm/tts7gl95cUi/2A6aIHPaVs3mzyPkn6cmzrw4dimDG
9eTqTVuvMEgkBFVgYZc5+u16/1n7wS/BWi5J90PotkRuaYbGV61uK/Wtl8K1mhZt
GtRSbvGGru1oTVO/0dgB+WhJwn08pPgdwFhD2IV00E2Swmr5aoe1CCSgwQ9CIt+e
98W1Vo7/dC2m3KNwNNnirto/yAIOfJOupJhYx0lZLtBdOL1spqoNMKJlweSp8Pe0
szKs4UEpC+3riy1KIhocUMI8XKIfDhtIdlbJ5bSPNe58HVAmnlNR8d9nc8UY8jXs
CWmuYJ6Kqc5YeUx40AsBkgSCPGVMKL/AFs5jdCMpGO1lPe1oW3fHUjaWK0eLO8jS
hP8Mqa8wqE17pXKFZWGt5XZeFVYNMlnM+XpXt/0iPyj26B63e7Ea+nOvZceY5Tzs
temlYDH5ObqBh6u04XrpNsdXVtgJPsE0Vk1Yu5cRBwBjfbpnUvAd6lMFU1Dy/1Fv
p7jgigKpgekXhAaV/MrHtECEhyT9/6eW0Irqa+0BCh+7I8a8lJ3H2LL58agP94ik
jqpJ3j4ar6xlUpekyLnFmNf/7THJDiA6448JfJlIPf19+Tusa0N2Y9rMghp9jKge
4Inr5GR3UaEg3z5sBb7YG151T/JkAHkoq8VAA5tIsu0mhpGtsO65G9J1OxZSMwzy
hf5YQRzPKOB9whmMkXeMkt4eU0m72bK9N6Hhma2l4PgyfKTVsT00FD2XECXrCz2h
EgtZm5J8UO5+eTpwIt35ZU4CA+DOP41K3rVq/4qFV3hDsvFqkkbI4Lc/TeMb5Mvn
86FIzyE/Sgq73e68kG5L2tacyIc07+1u6ghqA9ZsmdIqStmpKAYLbHilaKkTFj+V
aJvgb9+NqijHptoDZ+c1THsuWxlNS1V6/G5SXO60Ox9G0mAt/bi+gtIrlwp9ytZW
1ZzHNgJ255XELKnrz8TO3iipQWBQcPQWId5oFdG7nZdXmjDcZdWMfr9dRqbpsA6z
bvm8lrojbVzOC3W1iLvnV5FNxHTNTCxsxgB3XtldpzL/o+gcfRvjr0IlNOHq9h+C
2Pu324nn0+/pYwV4j9ZXdNaK9/GHs44UGpnPpdWOd+ucT5NFcmevWPHGrf4l4157
8fg7ZBMWnHnai7TBcs1cjM7/dp3fwhEoNC+cOQnFZ5+2l48ecAenASUpX2ZYuLKS
c0vkAGofeUUbkQuflwYrzaJuhS4WEyvLSW1hsCqZ0aNbHkbDTjysVwjpbxWiUjOL
oQGa8XgPwfawMHor+ioBfpy7E+bcKpCK0WIhyj0SjpnAwWE2ggHOjAyBhJ3qztAY
MD8WaJZL5exunh9OUtji4oKQ2PG41BzvxFTlsIWbISybKhMLoD5cZ1nX9YWycvNp
A06S+Ktk9EVcR9SZFlKIauhMrMCbbKRb9FYTzCayXTFuF+6SOMjMzIRCimX9IjkX
B6OVO9iIBJmkFAwr/v+iVli1jfGq+x7Rlz2XBNPuVcGHbx3kGm0R17aMO8WQ7ITq
hFUO7UjM2ZHJwghWgP0weZoD/aLjz+Uo7PkZ3HblUsNNVEkdQl2YXQ6L96vApSAZ
hsaYhRttqP8q+nIchENHQ2Ech9XJwMSvEX3Tb5am3kr2mcUtFYrkZGJBJEENld6S
RZuF6zxSeNU2GHuvnRWd2gxg6NGyAxaG2iTxbINBDPJ2jaDI3b5h5A8KaBX3SE/p
cxxd8Z1N+zJIZ0S3BqpUXT6hc+u10zYZf6um1D2R+ZMzqaGYVwolZXK416edeiop
k5v5bGx7PmpMh/tx9+OwcMWFx+rUenVZI/9JnjleLyFe4P1fAT0SIZhvGuXUGd3F
M0qK6nryyvBR07WSXxDh11h8PdFZFavVxRGVnGcZAg3AE6Ds/fO9bY7sI9KbTclr
YlkjGVVunQ0FTJpAJWJKv50quXq+jGgCy4Be0+PzgAKQ00I4JwKEBq1hV5SNsO2J
5czKibI/aVdlHEYmDza0+cNv93q7FwhXR22X4ctqAAC0C068ox4VhYXWlfmL+hAH
r9h3h4l1i2K/W/KghoCjmCyQjkYPin820woAcP4y21BhKcJOuGq6swjNF9VNlniw
V8V0hdFKT26XdGp7T/5VqN6tHmPfA/rbrdl5Nf1LutCbcgPKIWt9C6fCSOP0fL5G
pZXaL+vUBU2QYD6q2hzFnp8clL3epgSpYkWdsKKPp0nvWYTEhvU3ev22WudSTvb6
N/Qu9WZj2Rk3jJGNdWmI5hP5goUXEB0e+NRHYnP1/GkfiCYIyHhS/UNOpRZQxWQu
nZoNlk/TgDDsNBvXeOCAYTvEDQhQWa9vbwyk2AmZPq6/AzlfRVkQBylwhertV03O
/25SPQFpMKZx1UtmBlWpYxyczbkDk2HhkpusXcUae4ptK3KKZwF7C5XANahUXTDT
9gBeBjs56yftrS4cJPzvTAVNGegjLMZa3NYpTio4XvMpt6z3MRszGgZnV4kPMfji
HIxlXTzKf9tkASJ4blOsD3FUZjjRr2+mzF7iKUZ3xSFiB6/RSGKI2X52ajG1FlaA
uzMoL5Km+HCTrMZBrAZM+Rgetnexeb8Kiiuf+l/N/CGj+428oZjRu/DfxKcbr3KA
wGt93tvanwfyLAytMsz9l7S+4imuYXAALU8jfS27NuKBCqNAIhopcckUfbphNOeG
oP1M1ZXpHoKr7+Se+RQYdjgMBMS1bzSr9RT0Z02X5axSxQZB6HatpTcEEytxc6iv
IbuyPVlGreJ0hlj1cAOP0L7MIaiKikzBCMBUnjC4ba7pFQwi12FK3JqhX557kZ5m
cyAmYZx/AxNRFzkvzhRQbPfPC8SyMCex/K58pkoETP/efZZtsYqJoIq0RypuOXQ8
x1f+l7CbtwXdmwmx1E67QI2ZveADf0HrIpHwvAJ+P8eQnWm9cEglv57sKJ1m+gOu
9ugz5g57PovTHm1S3ACyYSsFByAQIm3d3VQdMi9c4DOPJGfN2rYnI5aa96X6x5UD
TrKPj2zTamBHyk8IC5KCOr0z80GnvpAfRUE+MQDCGpk+efPdh42bJedv8bvjoaf0
JyH9uz4IeQGd3A0F26tIOXpEANv5ixHrZF+4xhNaRiavUr4X0vEktMsSy/ZzvneE
ff1apWW2OvlYUn7E4FukboaHhqYlxuF2SrJSxbYdZGD4L5Wuk0xQxJn2VtgQbkbs
8um7oBWbfBNiT3DLkW1zBYYKvoFFlvi9fwjvNTm2ludrzEL6Qb1VYAV/vd+djgs2
ddJ1mZAxdGxFJNZZAA4navZcThw1BMCGF7MD6TUzDRm6R+wf9EdkoWsVSdhnDepv
KAeoarxKu7/F/hytQ4TO/y+jHX4thWpFnwx56rc1Ky9/1Y5mVpgoqJDN6Is2axKs
/9FWHdb2d2qW1q0Jsc8Pflw4jNYN2Y+pZ0IsDJO1oi/hUXm+BiuFuFEN7tciQzx0
xjffHAEhkhAHm7ymCACMG00hLecnv73JmyizlZQ5ydsJKK3KFIkT2BEG44RXMGs9
ofykv2tnJK9y2TQqug88wNpAVMlnm4p2bxbiRrgh2ojMBcguXmasncpRyIWEykJx
2/hg/pxsBWgrvpCgTC3QZ4HX4S6VdiXHcsj0+yrmqshvYoRuH1HS0nXhUyg+6SsH
DARQ4tNA5hP3hHgp5rNEAmkWSo5hAXUAmcKmuNGfkf4NCJzPE3h94oCm5WwU0dGH
xOdV3+T7jqmkdBrn5Hzl04Yb8VmQfFTSoY80ufX3LxpgASj1jIbhXDc5GCNN4UVW
YXvwdwwwrgn27jSTGZZctjLc5OuMERXvqeKpTEqMl2YPf0ORaE21eKa0sBILJKQv
NARkuJzZPnFhCiPCtY0/kAYevXSIr3D8YYOxhtC+vaBoDuPNi3RAqetiTa7YhYZd
MgqzEE3V/fjthI85Wze8/NgmpZaH6Tvmucj1DP6CAMcCHOInaAaufRqiP5HuygKS
8Npwa7PJebDa9eRx2kI/Ti+UQ77CnZkxg6etbyArfDcsBSyyX1uqpSIe4aEfWtSq
oyZqVKWx9dM68pF+ZoVC8SaTuc7931URza7uGHgg/lpNubDLgEQgmrN8EaIiqVRb
W+jTuqpIRKoQO+3EzzKb682McyCjWxtuVC6WQUrLEpt1bS0zDFO48WlIYZ8u6k41
F4vU4rt74HQWrjLsnsHhqTshsv1fa8Ghv/hPbPoYFn8wC6KglCiDZeFHh71T+sUW
/wb80Ng1F8jT/97NtwrKBTk096EoBw/wusxrWkTvGUirQxQ+WyOU3wKwhQAK/9vH
MU3JOt61ruUQXTEM6jDJb3GMw/5viqiyEt6COLZBueC8KtAgYejX+LiixUAz831s
JLxvRs8fMzONI4Cp0n07s/jj64nkdHyvj0xTBCbXkAmzfI6ysdqMxP3quAsjNphS
FHnQws3J7IRHGHsiDBiMzeiFLsVu7G6iU3b6oLs5h89zt2SnDYEK6w6PYPCDOKe0
oeK4pJfEnAVR62iRv8ift42pjyFVEUBSXbeOPpbDluaHo0FVev+2F1RKLdcj0rWF
075S8tjahfDP5bwUvXRcG2yJN+85xaEG/MSWH7UamURW0hFJlpLHGXXZ1eUoZcWu
Z/7kYnpvvsUcJ9Ipt7iyiTLKwJ3wK+wfoc4TVoz0/F8SbKUI6sSPYvN73gSa223h
TwJHbV2uDJxnW9oqzmYF18JKavbVZsvl7BYUk0NiGPoGKoVA5JvIIibyIizhtGXD
SkPvy7dHyr2K7kXfWHOk88ZV14/d4qobhVZzWoJ3qBDYOWk8erCnnGkjNHhs6dGE
bj9+F8ffRFu+fvtpLmBnsBxG0nT1YeURNnF/pJdio2QoCrByu20SvvR51K6AM52M
E9KHs0F/uKtiH10eJA9CchICbme1iPr8Fi+qPk9WFVvBgNfL5Ge5pvk5JQbkkyGm
GQBmnVnysyho+M3APrwshumCZWTyyqCI4ua2c15CT10gISs0h7UUB98gvKuCnUwA
GJPSASzEknFQP72W5K5sBLD6c0OijhaLVn/cNKIEgmsGNnyAzIpvEyMGzlxAlypd
go06dD6ZjNsuR9TFUudvsQOgTVjrqC7gx+foFrt5c3osqB1rQwI0cnN+FJn0ZFGX
QCSrG+nJiEcMP1e+hCSZWh1u+23oKUby9nqrmJlx2VpIxl+u25MGPabYn13kr3pI
N0Fz6+qL/zeZGVUxK94qKXUg+M5BSRckD+F2rv9Ta1/kSGLwk4VRCmULgSmBGK7S
x6e7YMeJOR5FdJQiWBR8LYvZOTaw1exKHnfdYMtAK9WfyZgF+8pyTIKHuGOh8coB
67qjQ6WdVMdRaVsxIiwoM5AFEUsOCvpPFDw6BPfvcRsWE5VcG19xisqyZuPzCBDA
JjaakSSrBiwzi/LZQrDKrb8MAhclsOgre2WVzWN7P4SdkyiYQi4GEWmN8tTL812H
Xlvs70sb1mJvu7nWfFKuQkuwabfIDVQNNwGHx0NTyj0e+cO5tNRQxDLDgIMuBqhX
Mzc8MuORUjkDjufj8PZgmq1nRKOdqLWZRMxuUTDb1qsWHYyyGSLHOTBLuXjZ0tnI
B73Fp1btAg5jM9hs/XfosuWOC53vye45tnKL+hwiKBFcGLwZCaY6zFvZCcowGkV9
2FN2VRqsEncWJlzcvbEyeuAO3FYSgd5NhDh0qKpQ9TYLNmyszhS/xHmCMYqx41+C
NwgTG6QdAZwwHin4p/47lzkwqVdF6cW2cJiJ5txTMYBNfsTMir+C3O6Lk72Yxi0f
A6oSfXv9rLk8D3PDzAdf4UVWZZbm/DrdXB8m1I9E2IvFuarZO+q52U3JWSjlazal
T00K1lBRQuob/sXP0tqWTkV3jtK8Wn3RYLTL0DVbtVu1ME2MYOR0fz7nIbNGg+KJ
KupugNk+UMGqwYReIU8A28dnJUcVE/rGaB7i/9Fos7Chd5jaosGOdO6qDf1VKAUZ
YMDYQiKB4kdUUOkWvxc7D4wCZ/XfgEVB5HzSfhnTCXYCy7UxnpFuPc7Ffdf6FVR6
kE+KPd8s1UzYYP1erZypRJoEyhAGS6iO5abJULNOVHgXmo8MHhIzIEH/L5pn6/mP
vrwirmmc89RwFdFP4AHkPkL53u1K1n8yZ9WaddCN7+2y2peBd0WyHK7X3MdIbn4+
tLTWnP3mrMpnIKH5o/3MeUcKACG9mb6bXsbkOlV6J2dAHvmFSxNACNasE6qcD2/a
zMezE5Iz8U4bGbTASowgg1IKv6yiUlcOqpro92ctBSABBsaYCaELal6C/FXijy24
xnGq6LynBXsbCJq7KO0q6XdIimzGUxUfd4oRhEtw+ChQsZatrVdqEKeMfq7vg3eo
sl22RTAYn8GM6erEHRs6zlEys81BS5sZL9SWfhPJq3CyLjU58r5YwGdSO15HEDwp
C/aTsYwbBCuy1nKaMOh7jS9HCiacpRGRO3rOmcF/9KWHoI5lc0KfoVOY4UfMZRpu
NWj7AlQuhUlTWmDag/3W0KoX3J1M6Kewg+FRJtTpVkaialZS5FGGv/1OETMaqvwS
XWHizGXs8qyM+a4ekOiKaj1KoKiM38FU5GuybIHWJto46G2Gqa0baNiFDKvDeUH8
udw+jv87AgLPrT7OaXlvuEvhtOfUx4PQvpLlVuYwSNpzrhBZ991GuwRidjGdwidR
R5EQqF25UTz4WU0lC1o7Y0+0vcTdYsd/QJKOIZemM43s0wBbB75uZMon2+8hocgh
WyZtjZeyqMOL8HC/mBlYzaklQGccmi3F6coaAGjqqayzDWxJuseI6UWo5XMI+zoe
tgRifxoqF+7Nu0/iRSZdXegDu74r/8abIiR2mST+O+0JJOgnpiT6XkPm8z5o+5Zf
W8GMRqWoC6ra5PgftJ/O298DHVKbMjNO4whHxducczuEE8wd9H/n56wX2GpCdAaN
3IEIM8J7gDgXFb2ie3ksELX+4O4t5Obsbq1zsQUJp1rl+sSCHm0RtGoNXrrOT22B
lK+uOlUn457ZEamQE6e4qkejJsxkIY+D29Oj1GooRJ7fjg+LT9JeBpXb1I1uMRd3
uQebR+hWDAVyWzBK20FztkiJvYLMT59JsNt+0U5yRxeRHUGwGH9a/q7RjGRp67wT
nEhUN6MkhgSQsHpzlti/sMjSSls9BsYl1kRt0znMqfQGVbZo5YkfaXwl1jGt2jHD
fNXz/hmJBJHHWx7Da0awrlb237qSjrYmLyl+uZIOLauQpsSGB6UPHCYAgf6OAfuL
f7qkVTjO3KxWK+eFDkL/6UHsN42vEY9CdHkqtqF9QoxsPLasYaWnvJAU/W4P0Kpo
AwDYw3puBd2A0uiQLFd+NHVci/kOX3JC6iRM/4u28EAtllqqwBL1r+iwBdQe7+p/
0bL/rPOmKhIAKNwxYdgeoEYIWTOxW76JeAe1wEuWyeOYGHJ8foWw1wIWxln6vjNW
xaqhkDqkpvxlFeQ4FCn2r3HyBz3hCjP8l5FGOM7u5+Sbk5vhNoL/1E3g/4c5GJNT
UlO6chOlgu2gzRWuZIKcHpe5UoXGIOaUjttNiPdlcgMZXcNzz0tp07cxhIiyGSNx
H9N/UDdC5yUAQYhB8VGsmsWmPC16hnRmfGt8rFhLGIosy4qFkhaMSA7bJyExcgA4
ihzc+mBtHm7iXKQ1GxjIB3HkkfOsic+mYuEuEvF6IR1y0Ht2ZiuAntuuuJg3RZll
HQxtw9d92dpDIu71F0VFJsjIxyt1w+zMrA0znO25OTdaNWdVnX8j2Eyo2L1wsEUt
yh8yMthksMB1R6L0LFVaprB3ldonc6YCMip14Ae5ZVr3By3vTPLUTT67kUmp4Ofb
Myf+lh90yL/5fvVn0mmbXLslyudbUWwBRBAmQDZt6o4Susdy1S/buqmuDdrrk65E
HIpy0fThFRX4Z3mfkoMOGXvPt6nJUSDWD2cEUoLINnlOjP0HnX4TRqxBFkfaJk25
TFiySK20Lk2I3WMn4NfKGuBoF/1oe0+C39W7BGEWCFYZ2PbhEURxjLHTpT2iRlEQ
PW2vuAGAiZdrXvP9Nx53CiMV5pbwbcP5xI6NwFMAJJTRw7Bi5c1QzMhNElGqXgH4
Kjdl1Gkaijnayw0g14Zs7XfINr9bdgPfllucVBNyzNG4qfwSqnz17EDN75lFs0BZ
+e9e0opmmTPFpc1sMjzG+ej/x9tFY4/m9DWmNJf6LnEwj5/rGvgyHxRbvE3V51Bq
he2tVyszKvjfw6HhXzVx52RRJymoiS/Kej8l5EiuyTuYqZFcZQ+vVctffgNoevcl
7+uzBKNhCc1R8B/hgQi2KTzqRNq+HMttiov1p7wyKtj2HPn+AqzjKCmY+NdKTLSc
UCglPcy9XVXTe3xLZAt07v/Jse99+M/V4zgxpoObQ1+yX1k/JZV9HqAQTDfq3ozH
ptxjmI1MdnGQvhtJjUiXIxlznaUGEnJs5SHpJYOlmE+pu7IkiT0gh6rQqKOVtjo1
U6lZxOiJBQ9PcddynpSPNodbNiuTn4s5dhSEfWrf3StxxBe+FJdQsb9Fz9DHARDP
1pRymm+TGb1ZwxlALD/TRkslVccY648/28TzQUTNIkJWuGWgt8gXLNBS1BDxacc6
hzRxqSJp8CWqDJKvwj1kfCW4eSWCCADAgoQT4W01qsz0eMosg1VqOKGeNyd6OEel
wydbfSEL9eR/meawZncD7H6yLv605NyPMkkoelHvdxQX52ysM7qsLrJr3cSo2Euj
zWoHBYX+karwmNPGsMtwCTCsLYdg1YG6YlzKllNF58gdui1eU6xzJGT7BbmGEo0i
1ee4oNkyEuazwgz7hGhcNzmp3AbpwAWqhSAhNR3xLG4NKdyMIinppVi7CyVZWYUK
K83b1B2FTTQsC3O9CCS66ioW+4cujbHmNxbQsczRse3GzwFJHQ4A218G6LHqFNNC
goVJmIV02YyUIWQ19X9UfEqd4BymWn82eUaANvk8pThbj7PsaBQ2tbVJwYbh+l6n
kCE7cW1NnoxeinR9dJ4kPncN0TxIwy/LRRA1SXLTG08PITBvcyKfuqJX/fVou7TX
CJ0KOviL2yubR2Cf1TVcqaOnPKJGO/UGOpF6xbXFjTv/DgTV9EGUeC6c99xg0qMW
KV3NauFkVtP5qACCJxeE+8WZNPt0qHmIxQfXMvYA8ILG+K4ojNFi4F5qwyT32D2y
LPq++/ZTAAEs7FDRzHlEVnsKCgZzX2p+HnpEX97/tWwDzc40cTo+kfc0jgpypJoX
ilFg/qGkDlbROAw9ifSPxED0rjIWQ6sWiRW6npm7KBo4yfWL+Nf/YzxWglzpfWOz
SLmizo0b/BP43pkZkreWRKde89H6hCPPWK98fabE7hbmX/ccPAL/+S0hwP69wV60
43kW0mU0t4e70IIzndRwAFCHa5jfz+zE7MhSjM1ugMZv2Ohczqxyplb+N37Ra22B
d+STh+pl/VKSToTCbjfPa/kNowTt/SqFVHnfiEw8eEatP1YfDizhx5fzYujaYmxO
f2hLD95tl4FGi4jnnhLblp1lRNusMMfrKsOHTT6EVyXmi4riaxrD50fiEgccIAgc
BDIwg+6OTwd/YaN9lTdHzlg1RSZ0mj/U5DRlhHElBav5EzM6YYqIKML5CGKrZARg
9Pojkb6Ruli6yEIvbcW/TIAY4g7YjqBZNyrRuyS+vqFFJlr+tYAuYcOFGH3Xge8f
wnucxGYulVciI5TEupSxoj1G7TqaQXORZLw+kyAueK8FXbwJnXr+frBXGlOczDk3
+SjGbWjzESW9MY9ZCV4KQQ0ZGltVEgiF6G+4xioPZsnWTkH29cN7M53KQ7ELTSBi
UmAnEV7G8uMbZNvedOhwKNEeSvO0J7TMlvYYv0jQzM/xeyjuP23iF1UxhKP7jb0o
egZMGnMCDabaXJ9sY6Xyqkdxc3QGZXxZarUnB+XP2k326eHSilPz5YzrYixndnR+
wIhueUaf6LPkr9M1WntF3SGP20kpFeU15N+pp3tgzkFB5g5GnCW3QJmVoVaOoYAK
fjCOImKJWvg0kMBLMyjb9j48rbWCvXrZpnMnRFBoodeCmOxuxCeBFMMWsjuGhN0L
MBfajGN1tB9v+dA5dXPP4XdBstc3Y229Olcxsau9fS5o33WUQNqJs+dE0lqyEgdq
JPq2d6DnpwPoTVSIhv1iqptp3KAsYVf5xxFLyam/1mrA0SNCAtwWmCOgEDOnDGo6
dFkxoI6tmP1JJEzW+wZFbR/QzhwfCnG0+/lmzqCVacVTqrm+mDe4/sv1XmSJ8pY4
OuWa6b7MLPE8g3Ysrzh0ge9ofIeTWyMoUI+aU3INumIwS4R97gEMnC+ZG2VjFW2I
9TRlSWfuLC4eo0gm4Pz5CKKI+VOh/OF7Zp1dbisWGy8tQHFl72Lc9rfDJOqXm/6q
zeFyYQnL3fI3Eu8FihuwdlKgpzXXf8RmDSvuDmlqNVDUvmLbcCyq0UF5pQ6ouIPb
lhNEmxRZOzAphts56Fa+GNr5Y8W+3Z5kJ6dyYlIMFoLuGRQqCkx6XK68EMQ43ep5
JHKb8C3KcieDfTFUPbnPBIhZwHr2DHOq9IyxuKoZZKOXo+3Ttmly6HgjwYp/UbnA
LSQEEtbU8CNfv9cGMRi4LEBMTo7AhlOCKwi7NNuM3UpctcWd7fob0SR8rEbjn285
6CvqSzKKheqPnppuKgcdh1Y3Kf/uHMrRlfvYTCIjaYSrG4tmuAEY8bTgq5OjyPoj
wNBrZZEKI9wdfBDnsEqX+kV2Urbkaz46UbAw5bG0H2yWjGgtF/Q8LNUNlPwA9Tqw
lgr0/IouuzhAPvCwup78Qx7MQh5reIFmZps4Qk89T2pGIDX+mPotA+oJl2qd49CR
MPhzA3TsEwqW31gpTyhtBILT2qMJ4+u+QpdQZNtsc/LzkeVvGymaunpmXNLkv619
/F0aSz/nFusPFRx+/RA9BXYSjj58gz3dTkv1aT8BfbHhz24R1Kyj+kV4wRqCwgkU
ani2g31riX94QBDjUs0e5bOEsCwCyelFV1WzY4d9guELqGAuId1n+jOHNaRKtVDs
pnPuQNgDkoP/CFy1TeFYtW+Y4jk6VcQaorNfXrltqguMScPFe6gUPfz3fFakWU0Y
MfGntXmfecbrZIk9y/szUC4C00b7mdpIMMnX/75smMDtr6ECu8YamSvTjcjr8xiv
o3YBMjetdMSmCfXICYFnhOpQLtwvm05atCLNw+TufBXC0tkFWE0KiV+T/xLo7Sjr
zZlQhYdTnvxQh8vD/UE0ocTH2CGDdf7KsWFddo0jhtTDaJcXEP0PHC4ejKL0XjDK
75/4LrhcNYlgy+hHRtatqazdyC0mIKwX5dVHBrx8sFv6FQR9B4X+jWzX/EQjLDxJ
E7mjhmjxe8GnAuCjr9GTeDh/7GENi2ye0yiPX4jitJaAEBmdiFuXVcARzNBnjrYE
hVSs2NPfHFpFClOg4mYV5Us6JFyo6mYHCfNhBiI2VJo5V61LbMUsMDdP8vw+R0aZ
NovIVlFKdA0VtrYUOS0PeeJHEcJMeXahn3A8iZYZw+/cqkPrPezfApXikHUDXVCq
B1Ksm8Vw2h9YoAl4gBqCOAqlVtzEWPLHJb+koytbqahRzB6a77eXTf+XjlZtqNpZ
neY/oxWvyoaRAvxbixjETDtqQwP7GtfCyuA1UDm90L0OFXc5poMUVXs9LoQPr1RY
uU9c7OgTsphZB5gr4ZoQWwjDSN+UsmHtd6DHU/+dZ4CFJ2t80c0ix1YfQ/8AmYtS
KeJqxBfj8d1wFL82ice515vM+PFh46ysgapQjBaWPTvMN2lK6aj/KJ+6mDBhp06x
J0wD2wv4QBQ1i1bFFbikqzNnzGI5wWsr8u72COr6wmUY/ylFKV9bCuEQG2UHSVgF
nyMeKPIUKPWjFkrNdilfg1u6bb3xfs4XlzmE5KWl//o0CUH2NgR+OpAp7d4Wd7SV
YDPm0pR0d3s+rn54jsWzMIMbyyZbD/NbFZkIEw9V9NxSm1GNrm+kdiiB8Ebvb6tz
PQwM43+jHmfyjboIbhIHw4uCc+vyCEiIUHEKDdfYi7ayP2ajXBLtlL7trI1icCvP
OCoxXehY/HPwxHyoYFWxHudcQh0rnGIhLqURiPeQvIj+N51b3YJzXV5xDtmiwS6w
585EV8OqnfIPN8RTGRJHcxo0HYKlIkZxP0+/+ntIpj28U9UbPPpAuYqDk9Nm2asX
ca+4wTEPh2p0jLTUWJE+fFHmfgGNV1m6efOrUIrvbc5isB1RrAQtVs6ee83PcAbw
6a9o+qLqsX2Sy3+v3nPm80NKudjFSmIjwmPbGxk6xNWnfyvXGcxDQj+KSrbyz1TZ
6hZXPAzXzjuBnTI5cxeQAqrVMaogUddhuflbOZSkwVxlX8S7GrqkA85nRNJxAH0w
CBUqZYn3Ue/Vryxc/RgytwjHj3hIGmM7QGhsAuOjEmuhugHnojphVdxbbvkLVQXS
SkinKZiysUz9F4DFfEUyxSd92I7dxr+DWo/tfJTvWIvzf5dquAtfxJho1N1ecLkp
vZ7BPLTyoKNcdZLTlESa16UCuR1dROxt7yTBtX+ZMbZcCpVucD8yiusOOvA6rRnb
2XERDby/LHzpQ5wLxqYIv3vCJqNaa4n2YW35Fp8y8mQt0rvw3uyuuavYQR4K9HFX
1/so0Q4HMCnPPoFpO0/Ak4NPaTqs0tr3GewT0GE5lPEg6m8QX5mmy+rMDx+Huc3N
Z8s0FbQNNviovy0rfy9aSA/6BaL+aTBJB+ssS+49ywI1wNoVdqHs61+krYwmNcgF
fzcCO9rgRWN9gvseijCN1mAZEOC6DlJdaAGzRpKBpCII6/YOkW9INFcSLQAxeUoH
lfuN4dOcB2TIdLcRoANHtxXmcuesbq6RCbqNlMzZdGHxJKrgdfjZvhJc/Zrm+yNQ
idDqBu+WoAET3RUbJLyzX68OMMrvBNbbesKFIO5e3j++B4hvTOya4qmhNBtLWfR4
iNANpPnSYjMoIU8YlAy/64ooVlk84d42nPkcYQBfxXdHUydoh4CZoAYcxuMBbY/G
1AmHp4FWYJtvQcrU6WPDk6/yFdPhHJgOLE6NlhM/sEOoA42Lu4KYU+Y1WUOF4pcC
d12eAO77aEiLWEA5WHUexfHDxAry0HvarNvGXusInEMOfnXlDLg5sS4GkDEE8oca
F1zX4ITFGcSkN6zLRzdbHD2co2+mL3fkpKXvFYY7oz14ICz1h5cIgcYO8r79b5EW
6rpCmyAlfK3Y0RqsHeFY98pOJ7a/s3rWgtPhOM5k5JGyQUjpidzLgDK/9QrqrJU4
Pfo+kWU7++coh1mGyYMsff8C1dgFDkBMH3OwpzGdrcOQU5uY4ezenye7K40/kPQm
9eEjbOyR95EeH5jUARp+QAhmHfBVFuyWMkCVcrEAoV/iBZVOFj8cC9oy+oGvcY8Z
0+3jQiM6N/1gv2M4mO1xONM3V51adMk/QYZLccdipZ13G9MabjwTO/MlgvDkMGdm
e7eqR/pqarndhrtpgbjy4UymuDPnjOPuQjkD79TtCqrtAo6M9wrN0QQFj+z6k8Fb
i4Ee4NdPNfetoDbg9GQRukfjHGSLxobBaBqh8OwsCnpqBJdatHEMPOW0baouFfXf
wnbL6qapuE4OfxC/HE+VJ0AQaSO143KPtEfsfTg9J5NeqiesAIFbPDiuIEOO5LqN
Y79B4/eQ65Uts0n2cqewshJJOq7rLO/+CIxyysf9pBjnpvqvqH1oOWNRjr7fentu
+dIWSa+4eGuSmJaXBXbWMGQdolwHePXnRksU+Zu7//hfANsuQiN0BHfulrFJ5tV2
zlUQIB3wIyri1hbTNA4tK6xGEEyj0JP1c4i4CRjOImiKR+qsnJ52vHzCIdfymxvm
ynWb/iDwp1hRK8y0b/du/BiTFAdeBq54P50N5K+Ti6XUrFt7/KiY+KsBv816/H++
wapdp3XrMiwBUzg+Dqe4QHIjmYo4aSe1V3jEZpnZJClvdb3J61oI9vIt/coHiOHk
39pUztsZnJ5RSQ6hNq0MTHYRx+/dM7GX33x8PCX46/hWkL/3IBYe4GTi29Vjzy5K
tdVfq0Yt1vGuLz2jlI0QWoNH5G+Lq3u4i4EvATE7m/2+PhkuHJTVELdq3jP7f1da
WlN+z82uOWegQJeOp2hjLLJdp+irJ3/0VvUJnDom3Y1gleRbMuey75RGULn453As
m0MAiCdK1Ed3ybOdO8OvalAoI6sAtoUi37qR7IM70CPALD7hJ1Z3NrF/cxEUFWJD
7jMReODmBuyMiHGbhF2eiHpuoTyPsX7yalr7lTPYm0HxGkLVoBxBpBxUTAUorwFq
tO1rLGvFecj6b8CQ/plh+x1j/ZZLfodzmB7U7C+cjcmgja2cCvgmhc4qEXrKw6RG
H1IZNvu9pWyNpbx8q37EykaWhHWPSDalC3UM60AchSOlleYmxG/Z2tRqOLzEvm7d
G7U3jv25/aXac8+7r+vXeKfHEG2H+UaL/nAESbvXlE/P60iWo6XHwk8mZZ7kVEr/
MsVPWd6FmzWEvJSpefLhUPcie/YYVuZn2jRRHuaEQXkX1ivtvs36Uk/Y43uWu1k0
yW96bH9hip8iwJeiayi+4XsvLbU3g/LLVwg06YLm7jDpHOCwL5wtkMbqdd5iAb2Z
9kRvLViR/RkdsSGDFwO1XaCfy2Z5yieYrcCxdRui86EasJmD2Yp52O8Qs7sJle7E
5JI/7H3ricGi1ZIqwZCk1ayULUggclWLpZYRwhROU42OOElP7xriFzkPdggW4XDZ
G/BOV1D8L3VWM938ytgfMACPA0h+Swebqtb/m2L000BLCq6rD/56DXkVZNZCRx1O
y2wcGfS1xgLr3vuWEY40kKztrPoPjMqCic8ByjqUwXJyOSiL1nnA+WViQzMYGPoi
GQu1HwddUf5+lBOhznNGmnJDP3u+Gr9aqa2XjvLCTnm1CyeeW8PsSSRgNcjKtJUT
y5PwkALdX2RacCj3X0X2x54R8i31SVjXEugxcosYb9Bq9OZSbGav2ZNTuAWLxh3S
ZVuV55FFTcRBQopGvYnlekzAEQgCVrZbFp06TnmjeOpAFBHbuEDmlRAlSs39BTNE
HPER6U0MVwCv1KR279iGPHHV6i9+gOVVzdGQVNsYEc70VMNwE7pAxbF5rhPK6Lst
NiHIsQV2q/ezeYzhiAk8Ev6cAedjorUoeb0mLn8+3vfiJv7UAswV1nNO+K+QufoP
MKevu/4ot84oO30fI8q50qTkkJCvQTx3Y4oTtDfPCJJ7wpydVUFx/6I1qVTHNQ5r
QWknmgtZnsqQVLdfYK2zqJnivOF1n4SrQYi+9toMLHy+wIOEM7NEGSO/tvj+YVip
NbxQDPJ8zuHpBoq5zQKU9Mwv7L8sKbAx8+8GXLS++FbgPtdIhxvwh5agyEjO7zea
x8TPrBH/jXhkeAi8cCVm3skwlqSGibghr5GBoDrGm6gmaif4wCoZR4zJfQ3C3VAk
YavtN4Cvul5WlwhZn+YXE2DFPSQpMctFBrpLWMrM7S6XlYb6fyZ8wX19wVBATgLt
rxab+mOAzqRsCPD5oYOPhKgjrZS6rqpLBOXGMVuIvh39tsQBDNZembZnQ6JKhieQ
TZi/vU2/N5QVggtDYoAp94P5PYnYA8RFbWVq+d0SWLS1hrmZIeQR/jNLYz4gFF/L
EzJTo75vBZHR5AurRNbb3FVkaEnEshl6zsCURuLCvnok9dWU3eg5qNis2jQO2epY
LYljIc+ei9d6K8JXDChHUCCsqXYDqi/BxSQqcTbaOx8vkJ56Q9r7Wq24dTyroru6
ag/tGnc9w2c+D+8rpOvjfrHcJS8sizb2UhBNPqSi3qs6iFiUBzfYLh1UtoY+g3OP
zDHCMn7+FYArwMYLpgf7gUgd5AL+gIlT40R+cb90LRWXtWGdgGvsTV4/VKdKkqvp
izrmZpRhSWAQNW24cyc02MzhM+BK/Kn7++F8LFzJnCKQ9uAcmRMS/5i2u6H6gFaK
cB5YkU1zjlt1iGDydyIneWQfRywvecvqyeey56kP5pRPPMCvU5BpOp1byvqA+4uY
2xze6VRJKbWXF2DrYLVGw7kiWGJEkWaTIgPcDH4niOP2w+hocdNhSFaBeB43Dfk/
a9hSG0Qvpxq6LIJWgf7nkjsQEQ1C1S/r5VAKRyvuV2Lnb3CNL2H+MMaFcKVoQwVT
1fdFIVb7EkBn7PSH4O+IgBKCV2WNsDBM73tpsCOh8/bHluGwC0xRmS3XWn1FwWIz
nCbV/JiH+JI2qfOAUfE6ZwBxFh1Hkrnt7X1t2wYVDCnv6Zn34XNlYf5nK/YYHxyK
oBJWmJ+lWnEGGlyKSXGGzMh8W8/3WzSfOxkZ+fAxQWz3+BkCKu0q+eS/xGhAUfVH
giW51UEqJjriUlyoB6gFivZ7pa5WHlvuN+/Wny0F9XQME+1qs7zSSyKcjZfRLka8
E1H76WU+yBTdKUANsMkkkYzzeRxAvW0sZIgOMN8WgvtSxMbAwpYdV6DcIsjcY9f+
gPy9lAvZCAdoB7y2/KhA7YEn5idHxAlJYL0P78M1CTCb3ncTz/lXjyEMQIaMPzYR
3v3Yo7e0cMGUXZe3FcC3zyiVQ6qNbcM2aja8d1C2zLnEZwYsQcGOBfnbBtoloYax
pA+aCHb1oRoSvsy+mg+67BtGf6QZN309R3mU65PL5eWyyy6BuCXYdtqoYHkZ6nzf
tB8vfvKURXvw37MRBEtYbUFAzMh3lRwM5OBi42FywAEY9CXYY7fEaQ96/ZilBHCb
o6yHGmdTfXyTzqGR5QrmflMV4Hq4qhh8NmKSB3/rGaSRvPj+kINuqJPwy8g+/SOZ
MnMbPsMvNFMcl+P2fXssoxgYcmPc0z0jzLEr/hfecr783MlZdNSd99vHzUa1tl3Y
9ZIwODfRTB4n0Zg0NMZfSE3OmxneWPUKAzuEkrDUT8Aq0l0/eTbooeIs+yeSa2W6
5x2nVW30FBP5dga2DnbMX5KImweJdv8L6JQGkBZagBI0Eh1Qv77ZNWvAb+O0Ow3V
WlrFONxarGEuiuUMhBFj/ZR2vGlyAtmf9hUD/3ULoNlScCv2EpD7O0vUp6Hup7qR
+hrQ9TbN+8HxgGyDY11YuFpGWRgKMknuuGYmabSOhTQw44on7srF1GFQZ31l19lR
NX2uhcsyb0b21cfN3RBbIihnOrj8svEuZC9oo2E614AuiU24iXJ+/2htCS/bLFB0
VuaZucTScBWwJKVlG2f5OcwIuL5IXkOE3BajTJUZyC/pFGg+JEZyYh6I7CeAQnFb
at5IhX0ZqUMXBgnMDCBM8I3n+XfPbmwjDcCjPJCrV0Sc7RoIE0Lm55sDhL2uPXsH
KQJqXhsFLrByfeZ95z9IO1N7DUvnPJ01F21qIhYpMGZmTlVZlf2rRQ4R9/xjF7EP
msfUGsUzSBiyLnZfLrrZuXbEv6XBtzgeoA/eZiBLHI8rVND9EkjtgRofbl0SpIOv
p9NSYeBF4K6zr0KouT36SL7XCLBlIR/e/LKlnsJl9jeCLx5ruElcYJZTTC9E2oSW
HXb7uiBtyD3dHWHAjY4jom/4E45Xd2IG954atJIJhbZWTlS2AZ5FsW1T0CtH2iFw
Wiyi6vBHgghkN6iWhemFWtUAExQoQ6PUm4PBveOMGXSjT2gfFghPSXcl005smsH4
dTW0++gUCemD4zX8o0dwGlHtFLlj5LBUuiRv8VpY7YmQgo7VzY5gm0o3JG9hRiPQ
rC/u2QfwXPUf5KtJ5kTX9LtkKblTcjhEoq1T3+3dZx0C/GHBn3gNChYEOOdPDrTr
QDJS9n4QPvE66TAXOglZZeNjQ9RYrEaTb1ldLC59rSQvi5KbAQ82lnspTNA3k9QI
zgEnq/WDG+YK2djafY/BO6kYZ1427D0FVTQG4q5WQsyqy7QEYx1aJLY1fy881H8z
Mh0Pmqfc9an+LgMDq9JNcnv70wnKBZLHXeJYqEtjStm9pbKB4DG7iUFadTSTzVZA
X4ADiSf8lEfnULGSqqpB2b6H+Q/wiA4VYsBrgETDtPQs/JW4sgvOzfeazClPbIQd
e+u+avpoPSiiY6uH/Re+uPqL1k+QfuObDKSKHJm63d1VnyVblSxilC/MPn+X4mCY
IutiyNimpljXwWMDoDkcYutpJ8R+Dy1nXo3as/Jn07JAJhxB1D+PumtJ8oRQmgfT
aD0XqtgdU1sya9ojqfVqm6gl2AmW4mqhOmF5gc7yvje96nKJb4aglFEN7Dw6T8xp
JhoTU62Gqn/JkQwldPli2vEoz1C4zBBxe0DC8plAlq88TdgB9sfOvZ+Y+72GW0qT
5kKSGMJUoo57iQg79itP4TftZl8NCM09Vx0wXP8FVvLDJ8covMeYSqDdiZqM56fL
DkFEzrY6fEm4wLP4FxkhKbKxYM3iyQn3/hRIqgGlxzbT1NyGc7NOalblekoBhxNv
ovUyv3tCsNlKyIv+PHB9mOIwqClyYroZ9UJgd5ucabhqEi2G7sd+HFykUmtoovmv
CV5mJv0WW6Jrwm7z4JbeMUWhCZyL308i5omEhQRxDEQFBZ0EQcrpcX4KaV8/VfV8
Jzy3STcaUnmp71qd1Khffocmp+vVVHMjS8MWTkYCHHlu/Mypn5PlHR1cqY046UZs
70GkHIm+kgU4cbjf2hulYQ+aVwe4LZ6FZgmSAZNSBxjUneSn8VsEV2s6uv01DipB
y+zi0LO35XNbgBBgpMej1VW3eCkzxiS5ZvaiCbhxr822r2r2HJpe7jIrKGgHwzY2
jOH1HMgzIC58h/0I/waUHHVHpY3vmrsFJrEHN8OwrWvQJLkd4UqnyxnR+GCbqRws
ep8B/AjCAKkoHBl6t/DqQJinibbL3ZFWkNuoZLKnurKQB+c1Rn6tp+r5oeKlGqzY
3jg6BcOIumVj3C+wbF8t/gAx7V15PZmAlSNjJjbrZP1VsODCLiClazYJcoMrYR+b
JeX3uwdQl7cm4w+Ji+qnFZeVbXvo/IlIyR4TJpWS53IVh8JzI2S7WlgnmhSBNfsS
nNQ6vmPHRFk4So+Kvhjneoj4qtI8uQNERXaWwnQSm/yNhVZ7EiiVkFmmdP8ty5kw
iWaDPXPggsaYPXqo6eTjsiwe3DTwz3F9Z9wAG7ZyvSEjGJYurjugJvnwujxLfmHp
p60qYoPl8SJafnJhr7VO1UClCIgzdgAoYXJYqf0Jd9mlfe8y4inrZd7/ecckCirh
7CiDo7Zd8mOoArqzFEuVOj61Otx/mxZT/WiOMdI5hhWW0N52cArmdfShEYEmsxDM
HxrUJI52/Mn3do8ebh1ahn9qjzaY4cvkWepjWftICCWTMLb4M3QNOaC0vWVRIBy1
nsaEiQP0xMjz5H1biwLS8T+bhSmxKjcBkJ36jZVpdSTDWbWJRZU3HFdMwj6iWuoC
c2/3WU7Fn2qTC/iBuZ/AhrTXLgP0JxGkcuTELKSapXzyG1nmqiLo+zdniQ4PXyyy
l0ecqWFhbUCi1QbOzpSGkE7W3qpt6CE4xtNCeDP72v36DleA83cQABNl09fjo3DU
skgimg5EsAxQvNfWkGLplO7JoPc0XXFtuxWaKdkj85hZ0L1X/J3NawBqHDf9dyGV
wuJ/rINH9pKUCT9g7rCdBqbLwu/xBYf3mQwvXMNhw9lfK2pQgVft7049gX05wyAY
U6iSjoJE6Of54QS5EA5GWbi/c4Wp5+hsn87PUdv2cbaBTLQihFwt47jVy/iIMQ/W
60LYqv2UbgptxrSSqYWWvTyVRSf+qODZcsjHSCjQQVTEb0cRYB9sk9SquROj3niQ
NrpPlHQbeqsmZqobKQm1L+Gz0KhN0ko9sEku3BcuqngQErs8F+gkWHIbqJFqKLDs
rzRr+ukb0uIQLyOLIhbJhXYlESzjM3eSPOfuKTdoNfAnuhk0hRVrG1Y2JSpMvYYz
AmUPymsD45iD+Z+dr3HxkI4ID6QMx0Zm86OH+cFTjS2hx7sj6ES5jPOV56x1Vzoh
aHPEfvlbN4HsqqyhMasU4yVaj3lGOHczD3lH47uPCdkhodjrchfYZDnUq89aGAo6
PKq7Y73Bv2Oft5Vas33ffT53RY5Ln5WMV1a5NVomD+V4JOxmKsXsD0gGnB/J0HYF
63XGxVlfwLYq6sNWJcoY0XWgM4dl+z39tEhW+6nE5CBvgdyMltC66Ht1opJQa3AH
iJWVkh3GdHPCWq8x0RGMS8N/iV3VqagQWqsEcKMN2WpGYYkdfU3JhkxFoRfoQPNJ
wZ1ZYRlWBTPlyBA0Gi5V5R+wOiB1dSBoW3toHpzOXJo0V23S/0lAFzZkZvIH7HP7
IYag9eQbyz4WLQ8kXDJQLBiqRZygHxz0lF4hEkj+iN6hvhOPTo3CPrca+R7nBSmt
y7o/3QydADxU1wII0+r7pL4YBByT1SDjKGnNl7IwvOrFW8NMhx0BN4P2CCOJDV/5
CpgZZjIOcaXK2WfMUg5222AvolqE+G7ryw50U1TY6Dw1qs9yYb9RUnBYGeaNkpEO
tgVaQpBaGxSqyYlY45mOpZE5su+xrSH27Edh7Z70sh12BW361fH2GngrjfGj48Ar
Ys7HaxMQfcCzR9GibvrNckAwRbWCwY5k4hP2SDqmE18QzSWuyxcUWuTgXJ5Y/40i
mUBqhoeImRbv3HI9qkeVWWHu4wJFYpFIteLixH/rN1W7bucnuG/+x+Wo2nnLvtha
bAg8wFvRz0ipGGvrSoUSCPtXtz9WIneOMAqsJNb1pMBcQPlo6wO5nA3u5O7Q3XPu
FFGPbXmiiD5BY9JjiD3f2tG89bDC59g1a6cy30Gn5gnXHzF8etyR94ZC8w9E5BN+
DzhwiaC9yNasnCa/sB9gVoDSLkZnW9CImxzTJJPYx/nfLfytTmPhh5ikJKVQkrKG
XC1/pu1yRwCg6Ka6+itp4X0ZVXO6aptkYlzMDT+tV684Qr4afmH34aA+0dtHbmCV
b4D8wpkeNiJnYmpMAZ7imFkx1M/raSzHWSg6KhCJYH+Fu5AGIHp9gcqUfDUSvcBL
ki2IvuB5TOABkvyA7jyQLTx5PyR2tBCznYJuDVD40YIhT9ZyuUUV2blGKCe5zS1g
DP+I8Z9WW3oaantPHsL1SgbwUiI1kHzjYNOtiKAfOUUrSPaNCCIthD8PLOWCDBXl
T3mzd1CCdRDbdYSTl0d8YrZTIRaFQSwpmPInPIyxZQiXItvNPRQBxG/XvIPhr+9h
CdOTMzoz6CW/1O1gMA7ITsn02Iwkaa7jWWOPSPQAVSJuwCIzAJGxPcYG/ZWMQpPw
edjUjDtFvZpvnG61c8ZPHweHvoXoEk4Jb5fTx7lMy/+QQb0qFlDP/aqzH+Ebh4bM
8edEUJK0yAlxnce/sVrd8ck08ijaTAynZ1efKxYQyMf6UzjWZ9fmAIUT0Vg49RCl
m7qYdL0ff0su20gOgU0v6FRj4ZyS9mjToDs1DJW7l9zR5LN0WeppaL2lu2M1mB0H
EYMCG50v9UbrRqfy37AOAVUrz16jva6/zWn/u4fvH+2p+noOrqBhauYzejmBq7iv
WS0Gs16thR63C/XQLHP8HoLUEOk0AUZjFFHJNayAVvHtBe4WF3XUki+P+LbPako0
X63/PAy3IwDlY7fI6XiW+3p14TxSKvrVp+XKQ/fRC9lcrItQ1k4RoDPeqRTRwuSz
YIH3n5VhPwHzTAv3NJH3boVbm5mHEbRqjxaVJ25U1RCL7UEvAhnvbzJQGvaKkuex
5yxg1yPs+0CIV6uY4Ehl39mVqlCOUf9KlH5cqS4vCcLD6en5TT5cVzkoMHvBOA51
7gupg4G2pTS7uuvpod6w20EdXLSRkiP6ZqhwUhUITfz0l5mRp/r1yxMD92QY7t1M
zlCgAPnnpta8UW9ihOdhi0FclMEziufrXDUBFek0AE5I/qzvaiyslO/b1tY+lQHh
tGImzMzifWztQbzC2snX0r+ug67J0kRShGWwEdvUphrNoWxYf7ccvEMv6grFMJ1Z
YETsU2bku8qcd5Kz0HCJZ4Il+aznlLYJHR9bDvcob5CZaalMt/b9jOvVOBR2EMY4
lC7bLWM7fRsWorsGjuJm3lQivR81bODeDWIOawn0XLxoNjGwlS94WU4G4uTo2y7m
/TWdZCqMBHCF0mpIggK2lOGubyPDv7TEQuyL40VJWpg3M+RZFyuUjv2okjAUXLpl
RAqLdjI1bnROlbzTZvl+JnIM61SpGCgjF078V96VQVwHQRVR/zCK0oyI3ny2sEfE
vhE5frIBWfqG4qA6wZ01eVoEALUEc/2g7CnuN+34rnoX4rDpxUGj6g8Ye7F7V8+s
VR4M2lsIXkhUAzVSUoYwlv0EUlGtBzBuC4MPLbzhu3Usqj8mUzXU9+txZRWhXZED
F0lXKwFQXejOdgDq9bon3+llXry0QF1TSsavD3Ew6Q3iVpGm3Cfy8TRLcfkEWheP
XzG4Vf1l8kAKSJc25VKHmj0Dn/0LIFk1Eup+G7NLVBl2Xd37sBJZs83TmYTT8/8z
Ditmai15XehFpItu7S89TZueTmG17+/V813X7zfRRij5TkuZjDck6BV/q/TUDQYs
Qxrr928KiZFA9DRTLApelNx6Fbmog+wtDXLQymtVjXk03VqkzitLWg12J9oyQAS4
fiRDixy8ObdYMl8VFvXXfQVEkoiDAlF+hlYRyBP42yTiiczgv2FUzoDrPzOnPara
EP5cG9nicIpchiq9E3Y/m6yrLSzvgBAoIfXmdJhIGgAvGSQ8tcLfzRtqiochNmz9
oJhUS4fG/+vpt9avhJ22c7wr4x2/gEPgtpLWbGpf/7PKcBI7XnDipphFE2Jcb2FJ
mHoMtImu5IQ+iVV4qzU1hUjtb7KiD/hJhC/b2Xb8aKM9xWNFRZKoF+1q2mOrCJsV
lA4aanUXCisAUaczCvmFdzBcLG6Hq5PT687AyPypzvVDxBzT4370CKmsMJrth4hC
ep8GNjefgEu6HYMeokLBq2vS2Uryq2qHzJF93gEuATtoB04LvLa/56ihiW872NWv
sQC++7S79tckPZo5aoz6pTNrnaVzPo+8opBz8dgj12CGgCyBfpKB6KG8jBLNu5DI
W0AXlFJ+CT4Nh3AFsul/Sbi++lvqX86eP+XI3ipek1YcjOC++1qgueRuJaTBuSuP
Ei1vO3Zi8qVKgp4ir9Oe7oQ03LeFPwxREa2Y1MAMqU7ansmVw07Nv9OsXFaBbYpF
hkroV5qVq+KRt+Vsj824Ml/DSIUvk8DFLH35cIp8+0klz9qOEw2YSxbB3Tg6rvMl
Y/RfBWm3IYSRbkm4MmMU6pXWs9CAHUiow3bn3F2CeZV9F1zbqLl+VJhq3mjkgcKr
WTGFo1klZWeTJ4tS7YWVQoelON3p4/KserDUScVWE8kI00mmmG1UclK4Vf9Qk5Id
GvyIRqQnEdF0ixCW3C/f9BiD31pWFKRREaTaEC+uWNUNJYAeMtAt8zOS460GebJl
VJS2U5BUqYiXgd74gxBdwNO3YTgnxd3U5Xu0M/71FZ/mDEK96mWX2/j/fQNGxTti
t2kHB8ViFGnkIJOyQ5pLb7hYaro1JiDISR7nskE4Oq4dfLRe2zlgAzpwWR59Yxom
cvu/ti7o2Jlw2EY+4bolecADlJp+a8v+I4ITv4JPc07EltzEI7W7NeSjnZetNMZG
aaKNJgeCqUt7gJLpxcBxyAWY17vjIMjyunApr2ACumhpDMM2gmbpaf4gujnEdi2S
1Hsu6GgGDyOw17K5+pxilV8mBQkyYrRlbwcQTkczGyB5zt/RKOTZIsVG8ordnxpG
sposbskVzy4d5vS9FSJPapHuJgIhiRachXF4xOeATlIgXuSyPWborDGYVekeT4RP
ui+qGvCtnWGi3Vu/Ga/pbvqEPudPgIwN5vk+VHGbf1UpQIQcxnTxxLqBzpbNcI1n
5CS2lR3BXGKBT0YZ50vHlcH3T2rzCQxUUP5V+B7u2E3Six3Yq+QAsGYHklUTUTJs
V/kzjeUpkOL9Cuc+EwCOuws852NjmkkfVTjJb7byk/5Cz7Vn/J3hxaeD2aBlRdty
5jnzlJi9OOnZmqRtp12b5cKNVGu3bsgRkyAWJsuocJb8K91vabW822qHIjxlIdfc
Es+deWyF91BSV9ixMpHU5coVaePP1BAUchsnt20D21w1/ue0cHGDwuC74Ojuyh+G
lPNcuKPILCk4mSUZlFa2TnKAbvui3Kkchupyxp47KoxQc828Efp5STuEDEwp/6xe
BO5RZE60mwCKttPe6RPKYoCX+udgLnjmB7KaL/NefK9xe/um9N3/JgIg/ePW2+1/
CudIzLx8ZkB7uM0IqmUkfpJZo7mPdAff+HA6eK+mf5HdEfCX8nfcNGk/ywKaa2k/
d1dvlGcA802CzptHvMu7TpKXFVqXOLmRN53Dn/12MZEhsVq0ySjK4VFIeKSHevvz
HLEF6jYCLzrwSA3BTEyAwMWYgmfXMGLCj7cfqu7W5V79aDgWY1el3X3rB0ism5H2
RMkwmgdRTvxY5f3NyCv3u8y7vr/Z1qU6pTbfCEYEYSgCiMvAj8Y2env5lDP+YUe1
lWA4+iNbFN9AUU9mCCwKVrjZJ0n/fuzmBex+Ahx0aF01noLKKpSz7O5Sk+lJE7rX
izI+pER3ygaNkB7JYTQIY0DQXfPCsG1Ko2y3rkkzZmlOkw7K9FIly0HKjXAT4bma
2shmp4830EQbw6oReqRuDKL4XcpRqIwwaji025FLhJVXDITZJxaKn3V9iENkCZL4
K0FtciyLYy/DZF85/USvEjdqlAgpKVF8f0JFUfjtY9pbFCyDPFwfM2eMmjsSK/pI
AhWAAsOlkeVqXd0qLPKCI4O6UJP5Wl08VBFZIzawKpMIk4HUhXHoe3q1ziju+Oph
ms3wMCmPfqdV0QrCqOoxu+tVmDzIZB6Grug3rtlwyVwFvSJGuL0q++LPL2TTFvIp
b6OW6RijF1OHPZ5pyYrAsitVOQDcNFCXD4lTTCqF35gBWgQTT90idsaNU6ZnJfQ5
o9Telr5s0A3UHQwD6mzkhFCK3zBtjSMNHDnELsC0M/JKSBaU5ayXEcvPS+RM2/3A
Q+D/TWRG/qFkDvxiucIGtg0ulKXGvl5bJ8Q+TXzndO1lEI+gFJQjItFLUAL4Zb/D
VZJ5znMshUR0nW3XXSSX0Esc2Mf1YOacrh6unIBgJg6DGLHKULqInbJuE8WXXsl/
mRIRD/gRC05GKDuE5f/al6O2eP154yQXA8Deai/YRA5xAy3dc9pyWcK629d1s/Iy
9MotlIjd/IM/hRzLCqJuFqGL3UuX2Pv6hMOidlMw7oa2IRNVfCv8NnMORRONL6Wa
6G2WguaORj+/6bhsRpKND6ANgT/sZ4GRYd6a/BLbgyR+qcpFH6Ax2bLfh3l0/602
pAeUaiak55g4p60rTTHxFstxreCM6cDorSouWIe9RU/ojYf3ajDUKk45LWTEflno
7v1M7CHTqH2R/iV/MIQfRRRUG2lfKSnI87iJ5i2Rqz5lEmQpmpbYnsGc2BfhTDxl
Ev28OGdG2bUUkfdKn8yZazXiMVv+uAZZ96B0LOFl3fPLGFFdrk87SLFMt8JrjIwQ
xGc4rElRld8HCqCa3dEwwfIsZ+EKqDdj4JcFQW5MB+bsy7xiL2bEAvy98p1V/Ue/
QuPgrIPtPdChvDqkicJpJlcIztXhcyv3xK5GS5U1QJBDUIkgtXIBVkoM9FTqLyzv
Emm2mHykQGqvZOoNNbvZ+LaYbiOYMmwjoBXbNu1+2nUEKtYfptWT8K9O2hkJUCR6
Ifgu9hcVAEei+VdrnuV3XmH7yjCBSE4C3cuU/3ZlFLci/CbSx4SBqKQiq5ch648f
EXiV+5PIOgNR7yMuFUlSj/WGYWaYFsuEGgxZX2l7zB167Wj3JWSp8I3GnkS4F809
tCE2L3XEEks6AR3/N5Yfz8uawFLtiVfcmUAKX57RsN/HqnZRlzUT4RJM4jPF2VWK
JMtlO8F6y/YEBNT7tHxe9i5YRUGGOa552I4Rd32NTtswLPJBZyTXVt0UzSsT2O2+
J3irXi0u3eQYR/K//i0Lr/Xlk1cjKA5eW59Z8HhmBtncxZAAcN2rE9x+S5tQMIAo
KM6m77SZKJxBQ073y53O2CMPbTRMooPm7YFtPdXn5SjcJxjJDJpJHz/YVmikYaL3
1KWdwRoGCUV4zhmv5/6pLT5wZ6vmRCeCzeUvwWKV+J+7XPe/mAech79xAJl/q5ge
lepAiVALjv7sqFMbKb4RAM3BorwKVQzG3gGkdt4HIVeaESg7MTj/BPlqDn7IeZUm
zafTl9bJzKgMUGweJr5CmhO+1iwW0HLTQGZMbUwSEetKVwpTHzUgpaeSvgkNno0j
GsbtAuTxNjKdX/j9LVdQz11U5EYmV96nVtoWUGi7wKgNmFiUB+Bd1ahf4db9SvEY
tE9RmrqJpJn0frb5L4Qurc3KoGCHm1gFw6krYsCfaWhq5gcOYQygtd0mDVT69sT8
2mvu6x3RMSoAoPuis3xxNvaTBQZ7NT5hjixjQSdZueAU1Zmg35SS1JbZ5Yi/1aQo
Oh+ZSWVcJV2z+MkFAIvswk86bk8q9YGJ0Wr84VAq7A/LzytlIyuD4F2az4I7ci1J
n+nsqb2EBHir66CI5KoMMSd4BwRjoJYGCHKBMHhN1VmmQRcDzC7XkHA+yI/ZtRxU
UeCQKj0zD+rdyMxS8oA4Emz4ySPX0eNtXFlJMHzXVMAC9XpCLkTCqwHaxGyYyfBa
kcJDYVOVIHwOAPgc7TYE1iL/JcsNs3g2f2u24cV/phpqMIm+gD3mfQtsM4Yn9NJM
39KcZ+YWQe0YW9z07pjbnZzA2SzL/IP2wHYZKEAY0/0nqaifxKNFsHeAHDTvueAd
czJ3bbaS53eIAXx1MoYdsp7srmUuUVTi1bbbCMAQLYTF/d9817xNri8PNWjYuQwN
0C0exZ6sV4HWVct+gYGiIF+UUIgQkxMPPhAVdisBXVK2GovU6Zdq028hu/riK1c4
uDg2F15lgv+qCmPKeBltyNVMWLVJYXdTjlVTPE+mzzzlIhFXajR11/yp61izcwZG
Gi7UqnFEXMjGF7K8gyqjeVTZ9tfe9IsQTh2D/U9b5EUetL8W4m4q+ssmy1mWG3Td
o3TEvtYTB6pnpkDJrANlPmvTs1SBz8C7wg+kK3Y1qxbMCvP8/ACnIXpAxhx6MUQA
nw3Q9jcZrPQNZYfCGb1jk//oUEhIwCyXLTcDywpd2pbVpvFOu0Hd95eAg3YNx5CM
flQ1IJxrJC/YKR123rsIEajvkyT4nQfrTzuY2A8HplpBd4Vwv2lc3bGnFLJ3c5SM
LiIZZS2bH/3S8JVTkKA2snT/BfQKAk53zc6GRYGoG4+Fdiw1ggys+sIaPdG2o+Dc
3l6LFmIOd7upW+fTWLP6mL13KLBdxhCNtT0SqVpqhwpFmQC578DRbeI0Hnbopowt
vMbIzjIuDF+xtTmB6w2dA5foSFN0oKq0U/v8GULMMtONoDHx/+KgU7hzycx/vYg6
UpkCNYeR0aAQ46lIdrzgfeApB0QewPghoV0a6nvBBSHI/EDoHjvNjq88+iiY55vq
NO0GURkcbbXNV7qyEUPxSkqsUEyoimHsvykCLS2sGQdO4ws9/HA1XYhnEDDTXlTj
hXJt/jKHDEvA4T8M5iSADNIlJXjwcZ5ocfROwegYJOzGaHRgZ4YWqV4X7Vs2U+SE
WX/aJYWpJKaNhvuB+s3/yijDlCZHWk7kZucMjGkvaIADMStoSP5vQByOyXBN7isB
0Vq0aGsy5WnfGHb1PchZNpUbpTYt8qlKzJ6lCoiSk93ICoqr3LwRvnnJCfyXnJIS
bf60XXVGou+mIRVNDOAKwbP85GocW5l1BwW7p3rtudrQv3NsKHKsQ+tLfEu9Jt1S
W0oHoC9k47+0PXLSoV87zQZ9EVoDmGYk/xP0/WyvEQQPVg4S0yj0YN9LZt3UnfAw
LuN7WBvNpjELMccZVFhDdfLfeLhPrwqO4kf61zJjc9VbHX5tSd6ezXERGaP5b4mC
pWOAeOnG6kzdUgY7KIvXSSZFbodnASDgZHbHJDnQaQuiXihdDEyKW8dds6u39RHR
rVh1533YH/dAdCJJhUa8enorXP2ct9NQmsJreL9dBX98bcFPvMuO25HoKIWhbmJA
tK14H8zNzxHKtplhQQQmhbKzGtQMCtKUTiPVmHLNXjHH5dapjcUXjr6V7HO78Z1o
ZsPQYa01ayLPFICZvGbV6lUw5taZhPKGiGS1ElBPe9vTXtovrtjiSlWdBaHbhGiZ
nGXbWUlBG8fOl0ptqJmaeqjqVbqtZJpcLG0uVBQaUIrH6KrIkRpw1TRWBburhikQ
h5zKgLoqh914vg3W6uWSRKF2OZxi+ScBbFKUFdsmgcz7KWAQDE3Z7VNY4xyoBVMq
jXJNa2FW54eLdIwFgt+gSs+Ob/0qmVkX/cmazQ4BFZgKG4acTEVrqfu3ykamEbeh
b98k4f0lq27NVtiw4Kwlx2T2HoLqPNwH/DchgIWQObnj4WBqf0QKPLSN6z9GP6cW
JjrRN4v3j8QVsuLJcPIKMj3ERQ+1DOCsCW8IzqVKLRpxx0LctUwfk1c35cgeJbTR
fTWrxpavNfEaW2oRlIKQInH+3uR/V/6qp7AsSYjhM1VYQryR4q3215KAabLUOXBL
J6ktibF/SvXaPy3N/AOhOkAE9rVi5QQQC4LGG5XLPlSy8wd4iEpM6AYELHl1TDeZ
fnojqSlzJ3NXqcbCfHj8Us/abax4Kveli45R99ma9kYvsG118za2sFrlwVNd9YXx
a/9s20gST9jLVN3cwQO62gQQVoRXKJms6RZIvdyjJN4XpIn2CiyM5yF5LnpLj5OM
0hH71IqrDAqmc3fFGyMP0A8pTFjChEUl20Vhsy3DuOLbxEbgkjS1NvaJ2mH8k8jK
LMn6miMtyKwAU6wapB7K+DC1x688tE8IszD0OZi/GC8MqRA756wPiKgi8zilICvd
1vL4pyX2keM/M0mVQqub1iUi2BG4zVvMKPZVkb2m7trW4okbBDiJ/Gr2O4D/oNzy
RMcdsY8WQASpKP3yN9VR+OvQdqy8kJ3CyvupfV/lf+k8+8S0wtAyUdU3XwEjpI4p
MQRWa9PPBFtc7KbNgdDsaFI/I7d/Zt6Ea0JJmSo4dY2VAqQc++imhMLoNYF8vEgy
gIDa6+TTS5yHg/KJ1CBlSFRtgQWY8bZKQ43b67ha/L2v0Niv80jLYGpXD/W55XL7
XWWICczweQxk1xS6D/h4MZ/yh80vXuiF8Tqje6fIC9QFxa38tJ30D2XCnJAt5SuL
1CAVKZZUAr1Gnpkf5/2QsWrqm9yE3klKvKSUQs0z1LCb8kljxeirL4nz4kThaA4c
YBZWvKERsQbSoG78hXVzPAOdzpdC9MC9cpfW5dMjLS44aH6YzL+2tRqK9DUB1zfR
jCWm/pZCp3aJO5sod1AeRPyFuBkUYhlBSCzJPdKDyVROki2jTR8oXXhF2qoQMmkx
CA/lcU/y04tKSl1q3Kfq5coVcY3+h4yCUJgJzR/1AJKiP8J2tf29eRiphsyWQmmH
8BWcTnpo+OVaR+d1lAvDUDmKOGR9OpmzIUFg/ZwXPl5JNEF5tbG/lnIOaM+cNP6L
hndiJXqDYGMhudAUj3bVyZvBqgS1iK/b2MTtkU++sSJFLC6qKtJEyI57PFqZ0WJJ
L/EoQITnFKxh0/EuQ894N81wXZ6Myy7i4xWV18T+rlLqKLkyiBy17U6FW/4G31bn
e69sdFWiczuIhoine8MXicIbynC6QGfiFsXyeOcBCxq5YYGXmZpr0o0KpbjP9Ntk
DH2jN0myAtcNZ6erJP4HW7xyaFaU5tw5EqeQ+P8wP1W6lm3qmdnZdMu1I+MCvnqA
iCQ7cW61GdoUM0gbBFbz3o9sepoMTWa73Z8VJgReRt+5jYoNXGoFVMSU3HVYsxH/
V3jsnpuSPL4gQzmEYi1nXolx3BhHXZDdKQBqCoK7t7M30Hf4I8TtwoHhzlujp0D3
nGT3GikFtVArRtFW/40DV3EQZtrMYXnzmAJX7PKVBOMVsmHzjEHdiVEGG9QrtD3Q
tnl6Y7qk5sdVphmGn5dVYCvmLugoBzB0TQNLRDa+N8EG7mEFF48mRxuXuhD3WDLS
xU0/Iepgn5iKtqVCqorWurd8dtbLmKdyXyy6c1OdWm/IdTNmWjKg6mlaCwJb2dsL
Qqa9wCKuJyEm6GVm3LDIWH/eJ2fKHszH0T3b8nNh8NWj7G8f3mSHayJhAke3Gxm7
3AzExE2T62VB7hw0k0zf7O8t/KxV8Zs2YDxRvJlzfa+c+eRhqOrWJwdIM8pDfVE9
SCqpuLBWrP/J+1tWThTQCYts6Ye2LBY/l8u1IKuP6MjGUDiUAejLQiq0QR7OLAum
MnEBGo4wpeodDY/7lQTlmCNsphgZUoi6JJ1u0g38M0PKPvXb2bvp2vGvZdas8piS
8OrK7jwc5JsZ3cqBL0qlu/+AweP5agftZWveuPTpsfOfsWYAKSKssWAiw94wakfZ
K+OVUlmWr+C3C0ArEMmvFIs1y+ATDDse+2cnbUgf6+HPo5/2g1GyA262Ndo4YNa5
ZZG7VtMJYu1SrWCE8RWPhCkWZDosZkGwETQp2egYP76X2WqhDY0PrNeaixZp99ze
GIdJQKbil2UmvCMAUOxTKIbbdCgfGpRCCOqgnvTGB79AcqH3sumyMlHMxJqcckTW
fkCzdGulikrR9N7lsbcsroFMEAg6NuK3reuuSsw+H14kfxV7KSTripdNTreZpbHX
nr6OpZsvMYIt2WGV7tat22Sp1H1p3GXFAsCWpvibfp1Z2ygUJrzlOVNLBxhGJ4M4
/m3F0rRwosZAICywok8YvCp7ixl+rXGlPNetOrHjWEpFn7TkDRYb8MFSvWoawFMh
Atdt0f434qnFst5/QIxpVs0+fXY5g8Ib1VUxk5V5jd6R/C1ac79u5GBjl6l4Ow/K
/krn+7C6L/d+fZrj3OEn10oIBF5Cmq1gY71lc9r0+CwYUL/TCdiZCd488bdI5BL1
8X9Oibaj81PsbwFVvH9tJLCBs82fte2+/02uueLr1WBS0JrFWx3HVHtV/mkqhuIg
PKfmjjYwpnFySwFf2y8Lr5ro8SzT7qWToQa+AQWmdrhVQsIOS3/6LDrlSHPPCoJg
OvEPYTZz2wNOHlIMzwwW3gZGst8o1ZC+mV152fIGWhzyTe0gb3UynNEnF8ejanAw
1DiLKByfVx1eCE7yGU19eEOV7lbYyb2tJK9g/33X0xfSZ1nZogkDnLjgrrlLglFm
ZhEii379m5M/KHEreMSU6oCGQ3K5m6mBY5VVet6Qjzm5qPjScpe86bxAZub/HuIg
tp3QEXCODW1VbQQMVjHCZ7ZNNmZFZo8tyVMWlZCCW+xe+BrUb1A4TbdWJeMFkYzW
b1eoH5TgaJBhdNnn7fZRCnAogLvI/UStNuZfnPP9dsHGz4cxjmbNkdkB2nKvKLXU
eafPjZUPXESrVJUGkoWIsHZbRvFtXGNSoL1tPIYw4PdZijqKxC06WTpzkoky3qdE
w21gJC0h/SPru1yQKriLXFPN5ySQUsckHfBWsjvGLwUHHdx3Flxv6JS967lnNjVC
Yxkq6LGu4R2Tg/iIUOB+QcSsaUOQTFJnwW6QvH0mGRKHX9JZh51aI1pLqYtfVE8E
LGDUOKqYHH68LZRAdiwqwr+sgFbcT7Lvl/SIY7sPO/TEg3l1iUWl5iC28dibF/YI
OgpYfGOu8/4ZFHDR9dnUM0ww6xKVopcAsGIZD452W5vgorwqbJFQ9Nkq0/4jygOa
MQW+rnlu1ZhCBxL+1XbdQRglUXF1fHYPBB2iBYiuyEaW47qXuZo8lsgMiEdOH02n
Koa4OuifA3oQfHUaoK72Vm7Alej1xts/T+mqYVcOgSbfcSpNKHVKTF1sQfa5O6UP
hOD0jXoVz78lRFxtx78WXjDXxQtNN1JtcveJX1wOeoXXZxnqPoQVMPJ+1b6lZ6gi
vdC9AwAhi6C5U0/KqR0pb4635nGfOTGEgNgw1iPbhBoUwmmoepD7iFtpVvZnciNJ
B1sXJTXlrxX0CIVvx8sol95O3d5ZlprfVrwrLlm6301dcRCIrfiZ0BkfMX/83HzG
FA2gJgUj4VZPC2+uEFMLkVaRRLzMGHA2d0NNOqi4ZOTjPtSU1aMP+9LJBPnozhfn
MXYeCrFIR90SoUHHhW0x8+9r/fm+K8ilRs8I/MurUwkkzA3fWC/HYbwWjjvN9fmS
aDOAUFSmpgYbh6vI/UX1fwRjxA5wAqGrQCCMq8AeKepoXRYfGd5+AeSG/aGjHYhP
ruejsn4EwQIW2Va4NllUcXsszfOMU/U62rPayp36Ru4+wgQijtEdc6M3gtt9+Ter
0XgYIehN13nFaz9MIyghxbMIBnvl2Z4t5/xP51K51ASdMn0DMiqHJ9pmJ2NQgAQ+
0ZKrCWTy/9q5hFlnLPk50ymzWvLy0UBSWRLxalaUDeav5ZUOeWHPceokcA1dMEZ5
kZnYUe3x85FWHu3dAbem+Z0RF3HsFOqSS082OwWMtMm0Wufit/MaehSDJlcIdpyO
PKCOmJsXQ9ADRGJOfPZiNxvi+7wPwWMcmwPvqIP/axSG22O9KdYHaoTgnq9BGwPc
eZDSg7UejYCyG7JP2Dw1hmE4VT58W5asAB0TpwO8sEaOXKDxWAuM8GGmVsOjnSap
h1dOe93mJjehefGTfbF++54OVgtU+0A3SO2QCgnaFCkARuZ86B16dPb3mAC6f71/
E89FtKsdxe5PplNP6Dy1wJf/zg5AhaZHWGGJyqt/zb6oulJz3cmaKzjqLP0osU5Q
OjtuKaoDtSv/4vw8FtprbwJQFdoUipN54m+g0lqauTXyHHu0g/0kbhqrsOkUaStP
P03g3TvCKQroYiIdL2J4yE/hGVn5D9hsy9NhgOv0q6HRl+efu2NgTLA27Wx6lceJ
VvMLBA6+JjsOQtJN2TESPKy75n7jlN2J/7SeA5CO4qpjRazTJv67FXYMSf8YYzmj
bBo9XosSLZsbIfdIJW1Txq34qRT6BURGxXz+WZdKqIJbfb5nzzBewceyPc49Xw8o
5W8MWEnX5hQzKFuRAWqpGVFTQd+DDOH5OneEhFnKHuTCCqkGKX+9UtXJFbLuKKIW
OIeeDebqQISUfiHYdi6peF09r4CAWUrPNdKW7CzixqQQgovA9DfpF8eoOdczCRMJ
vIoLDDpKObPj/f2RfLYp0cMF1A9mqvWuCbYLyZPxcxx7Wqsk9kHBPRfeAHNm8N8o
RhAhC0kxrnIvHd9WcSR5+J4ESFRrt31+hl7cPAMB8SH06CP4nNfqKKy40rBhWcKx
FOJDhOQpwk7fTLfQix9hIcgr4vroXZlwhwoimGHPnC/aduDy5Ng9AeYTOjNnkGmm
rvUBBPq6orA6BAE78R1djV4qm4Y4fP1M9leGMa8h61vrNhjcSTvxasdQAYCDgwAU
RAx8MagEeExNxq2J2Tu0AuoduNzVVAp5n9AeuurNzQrowCbk3+Nze9nwydIBQLjV
+wmj+w1wGvADWgWXhrNi90DcyBbJvPbAv7lVF+MWVt4pnYG8v+0KZlUdrPjPCM9K
C4vBaaAxKWLAEYE/pRjOgS31uQVTZci62D0fHytQyp2RMAFLhhJV2AKlfajexALQ
HU6STxnl5zVhRA9IExs8YudFP5PnzK6Dr/3myKbFBPgAZU1qIDIkFTkWk113mHit
jaFsccsldMt0mXZqciDKtsN/ODjck42RSlOUsMfW1AZ+Pd/IZ3kZzxM+Blap4RPv
oYwvXJAfiJ3m+W5KV7mpF5oZ9j4fJjRYqizCsMJuEqN43W0dlG8VT6aK75uGBsXJ
l+LhC3ihuN2fWRf6u64rJ8uSSeR9A1A00rO+t4tjrtgjQVq3G8/E7p0a7W33ydmQ
DPy35BpweugDDcZp3DA0e92Y1Xu51NH3HI7zb7GFDzIB8zg9oYu2TwrPEjXVS0j2
pH8QGFe2sA7bdKr60AhE20Fh3vQoqEADqrqX8Sw1upiQxQhHxtnHl8jCzHmZvzUN
0ti/+k079j6EYO4uMy7SBl4N7KU3U7pc7nol+OoyPd1vdrXFnPzbof2KZTsMusZX
0fFXG9OSPJRMmHcFSIqh6dFJwOJQ2pHnLNzmWkAki1zPPavm7HGue3zs1RaMAXtx
WFzYcIAsnZourH5Ld0RzaQbVad4vaElp2jzBxni4jZNalxD40UjK3jypPNNHBEpU
Kboiw+8hc0LGBkRds7DwZj08fK91fvZFEpBMCZF3Jc0i7qP9AxX1oKYSyvy1PIp1
5eM65p9Qwy70tq9QwLC4cgaaMHSvD79J9vcaoWzBufUcgV3U8SdTDbkHkxX7+Ths
N4fxAj3FQiCDfD4xTQbbYuOHhUbaezbNKgoZbu5m8BlmYcXdFTVr+gLBmewjw/Pw
8lxCOm2eZaPx2pz/GQRd+zGj9HSUAE9rOT7H8EH19XIZ85AkyeQA1arz2vi+Y0jM
/JTlV9O9K2Mv2wPJXgx87rVvWhcCkQ24uR2Ccw/loatc5ymhhU6ByJ36nHnOOQnY
MLyjRJ+qdwTahqFbywt0smfSVAC8iGzdt4t9dSGIMYsFV1GlbIEyoRuOT/72lzw4
T+lYGdvhCt2LYUQa+eB9ZntYkuFaeowS5jsNaDVpgwUKMopWjm2PKmnnLKXo7wzG
6eXyboGxnHJOy44ItbqmSBJpTToHPybQiHs4ZEwOQRfLJr4m7Zfkl20h3VdBgFdE
ZtGUH+lQge0Dv6eDBk0aRh+SGq8J4zvfSNKVEdPDc5NhsCfJWIyLqdRN9t8MSlUd
4BhwKW/OVyfa/Rxt0fe0hy+nYMiVDST3f/bcCR7kXCtLtyNpu5dChUoIMTJbEYBC
4ImPUMDgE8cEyT2Sr+NdsLDi7ArgVH0421EYikPSrVlftV+NrKZSBeUH+f2qkBsH
NotWAW72Y2L3kMfzlrIoreC1ouI34DfEOe9Q1QSD3GUVP7E+56t+jYJft3/gBsih
vkxN7xH7/GH9sRHEOSyhdDdiXKgti1GlM+ZnAM88dihQtSkIc80yhnu2Qx8DiuVo
V3Rd44yM+ZWMelieHO4MeSj8cbhLZd/zdmmeznDxNTnbEKLTJ9HcXbdmjlShY65+
zIEQl181eI6TzErDQo05dPWz/x92k84YRL/AMGsSkbRNaSf//pvHcWng0F+zInDE
yTkBXLLNm03QbErUqseJSj7PdTJOT66N9SrNksHIT7P6Huqi6I8Ly3HyE4Z6B8m7
fAplh0begK153DweXk4/dDEwpBERpNSYkAj0BjqS8DSCF6PzPSIm56F40t5E99VA
KVcdzrbK0PqpfhSMNbVpqweuRDQg1uj7bBdzuzJ4wE+b862xpMYJHTAqKr61qHXx
/i/hc1ofN/+wMGYDnA47FHYIDhUgG5RFqaa4YUPlSQ9EGoJ6Ge5NNICtCK9+yNVI
RLCmQQztrtkLtfMA009eZ/a4Egzzv7uefXHZV/d0w9JJubImB4Gt+kSA3lMXWMA1
vZ1z7Tn3D4hRp1nSabTg2SE0Z5AyxS2WbBKkk3VMGpEvxZMrTuZiquX4AmbHVWX7
f3kDNYV7DsNc3g0AYBLW/whnkxqexmpt6dfOe14S3dvxTpgcj2MnwB9LmFs8+Awr
/2CrEZ3m6IWx0WAesUL9twpTX6zcVaQtkhjpzSQtkd3lrK6uiF2eIQL7e2JUFO92
e+qcx3dWW572ODUtKC7t1gLANWg/IgBDShYHsYnIrdqHNzLjShHx9E4QXOelTbhI
6C60J5E3cV0IFUmt33rP5z4mNtvT8biouVps6HwoaDSJ2kAubbl4zYCgcqKJltOZ
kCqvZ4AadY3ZaolRvbYEuABMQPQMIlwBDw+DnsBB8ylKYCVCSZ6s6r+usZDxdoYk
CnSBZ2phSRcAskCnMa4mO/6Z4YbQkQ3MFABpJCKhkfckIlmif7ZakRMcmq/vO0Zv
l5qAbYk0vNuM0pG8Lmq8SzwdzDIVdjlSzo3fEhZCtRw6WT0D6WpR7Mql00Y004MR
czZbijBIYaNTw95Qzg52a/2+7j7gIxKNL5yK2bxo3DRKb9zWnDmYk6haRN/t+hSo
Ji2p7XsYxm2xXCNdQIT6UeAyjgDhKdRerqR5EGWPkmBUsGBfLweD9pmWmw+++MR7
Gf4JI9dzfOY0lRy2z3Jxm/P1VjPHMU0pdaB/FVKq0Vq+SsE7oVWVfnmpXGn+iP1b
Uvd3/Tdwp6rJbT5vCyjYmvgUsUExPtihw8inY0mrb/XnCgcGpceG8pJjSfZsowM3
07tg+2d/9WT4uesaaLd+Nd/Ha+84dIbsEIJWic6i9qtj95i63sjTn7ZwZz9YpzF9
FGmjgGwn1egDXMa3MN/Msv1EWTEZdYleuRm56BgoPHMU67ALFHzkSBEnGZmqjH2N
X9/JZBDvOYcSvKbrueM8m+vMmVHP7jwkeBGCDI7JHB2vy/VS0weWvYywO37EX3VZ
PX7WhYjSimDQJXYVLBgxBBUS8KZkr1CRAOSDwiUgIfFWtVlQNhsq4SpxZG1Lz0z8
smiXW6VaeqiGnwKFhQljQWvxavg7C6nvdNDH+1Ew0BZEEQp3lBh2yuB9Jdg74aPE
GjdGkxfY/2RCwM2Otk9gR1vEl5ymWrEXpcrygW4UBhCgQk4ksLl3R5fYvLvNByV8
qM6m6Ob15JDXwifzm2WiIocHGVdzi2hl5YDzIxZnvbperhS/xPd6rPPn+gjrabR2
y+dkaoqi8EhkaVMp/ocyMIxIpUS5gxyUE9w+Tyd+ijVBm9iDgHBSipTRY7YDVtzP
x0Q7F6FlIM+Z7FIuYKH29z5yjZHn7SOIoUxLVnng5VEemm6jh9mLjYN20PPfZVeA
uUJKQWaLC7GD/3HhZbMDCCKALBCXxf0264ZltC83pey2z6/BwkPfXAvYLiICQBPF
Q7MdhQLjRhHwEPywszlXcssM5KuVX4LOWZyAXWHri1yLzPz4HEjZ8LmZLzYyI3Ne
dbG0gK/Mjdt+gJohrwKLR5iuWp4y6Ttx37R9Y9E03CdGSzA0yCDvcyGkVG3D0Oin
3KIBXZWR2OEyYXEjMjdJdRvQWTyFQeVQBtDUzaqTw8hQAYX1GL1Ixf/yZ/cflw1g
04C3l58Fa0xicDBYjw+eHvYfHx/5OKRWyA29msICsdQnolPDMrhG/K6fEp43wlH5
O26UQpZOi6tReFp2krm+2orqCLSVZq7kg2ZFBa3f91S+NBwmEoJmZz1/3bYTbmVL
GGCqgvQSoEkKm8Tk9pF7ZYGny6BUCqTDLGs4qsrwPJOczm2N/VGgWL8UXJ7UB4ij
FDIraD87uCqd0Nh1u0ZSp6BsKy9NM00K5omsX5LmUBIK3nWuRrM/jZ3CMyay7Gqt
Sn3kmkNiDAwUy4Odp0gkZdvbwm7GH7YPJg5jIee71yNuealVMjybZasPqNS2BfVA
LJpnqRMrQecpRBu0cobH7lBBztKZsBkw2RSuoTDEiZoqjsAeSchBhVjyMuPOwWZB
ZgNvJcaZoJrntpaNBIi0GbneSoBAGpYrNFWTu7fQYE13JlktvJbOl9HJ80oD0w+c
jeKSBUUUrcRkpk9QPobwi9aT/lZ2mxfkgTr8MIT73uR0JY6qgtPmU8Ue//3LYgGS
k3CZsoKMPy4Ojro0Yl0Bno7cFiyXCvGoSoRdZHLlkcyJ+a1PKHqsWxrfKAm1UjmA
p//5fcCgWD0imZuKE5fHy5rYFdOLJOBOM2fDGwM34l6VVEyZgiQjPkW99OdT7YZi
IhzjQCdgYcwQnb3TNFg0ShwaQstx1XMaNzxJ9iqbjBgUhqG8XTWUwksN14AXjuFz
Cf9Q70GNINwVqG88Z5ivqGDLzef/qT191pNdOVETQ1bsKo5ABpcYFUgBrejUlcxx
VDm2Gi5IYs5or0H1OCiPhjK7sGpzlZlcb7AgsZxFn16ROomWDzKukAUMWMXgMEW5
Khz3gXB5GiDlIqdIQKrtNdhwQmq757kc56lRzfqww3rZQPeuOdEPkPAyRP4wLp5E
DzXm27vFtU0QYxouq1DogQYBaKRMpg3dQK2CD65pG2QOnWHAv4j+yJf9hxqzucjW
/CudG9/WSk9O/xlZG62LqAwTRnAgJmKHYBmtlGkrVY0jOq0xZahwcLdT63Lo4e99
4ALQI2f9dXoe1Se1gRMRv/5p6o7gUSYzbx/iETceJp+J/n6Uy0b78nyXvpdhQefD
POsHPtSdgB0wdr4dN62dEm49uKeDWUph3zfFvE48SR6BtjAdNI+GLorQra2XZNAk
VueuYb64xok6t3a95wv09Ukp2ERwUNiRmkBKZZV+H6cSbIPslRfQMxe8oedl5jRI
o4tyAdxGsqbm1196vNTRL0AXL/gKuRnVXT+8DcRUmhlYg2MQzMpm2UKzbERCgQlt
KxZgDfIN+iFkQFrEPl2PNQh5Wuw1tgX9eNiqYCPoqDL14Zc4KusutQTwcoO8sc82
IiU37CEQkcdwH3nP5opFSnaySltn7jbRIjF8OveytzNJER9g+RQpCzbU0Y2bJ+Ru
Q9TzQ/lc7jvZL9RS+2En/xWxlp9WlZjFw+3/sbOAE48U4lcr75RrYUTzquvKP7Bh
Fdb71C8BNmuLxdtYuAQ77rwxCu7tBYeLI60ydQ/4qJbYeD2Y4aBWVUqhnnfapgZx
LyrlZj8wuWr4bgJONz8pHf+BKZM6amKpcP9qZIOA0IzLX/P7m8GLNvqyFgxKtnkf
FJTsb9Y/W8AK+OXgQE0N6DftP4RfyIOi3MnbrrUaMHzGbvV0xr6IsnBiq0rnwaL/
uNKUxrLjQ2Xtg8sspfKYi3DjsgEdcahHyFq+YHTZhJp8gi1rZHVQBzdBSzwuduk3
kzS5DKZhtzZrgcK+0MDqofsH3vaaKgHx9yYvSUv9ccO5mrUGt0CQ87jbuRgf7YlE
QHluRFrit6cxH0lJWcjksQLwZtdNeAtRatOURWda2exikGWBNeNYNp5d7hMLNLdt
e2mj7NxBdcK+KJO4mI6OEDIySErhdJQt3iT9gyisWln4xpm87fsv1lLcaFg3Cmpu
KTZv0sdEclGkr/+/6dCfYSgHj5LHbIookjOJcbX6IzjN+UkDFOuHytsY5xB7Q4np
vavnEqCoiSm69sRgqh0+sqa6xZtRnY5vL0rIiFrG4hdV0LMbeu3M/L3hbfo61Y4Y
Yqwg8OuI3sJezI7wIENbe/mpEvfO8ViL5RNo/MClHr7QlCBNt3TIch4DCGz0az1c
+p6rJ3LDiKWUSt0M9mWwT2JgVgC+t3G+9VT4cVmwOMhQwLo4xW7K73X5vNuMqYvC
TLi2c2ZslJb5tKhWk6U7MJUKpn8wYTFKILrxlR8XkhG/n3yzOamIm2Smv1q7r1LU
Nq6+dQ//gN95MqJufPqSi+8icyepZ6xB3QcAYdJ5Stoa5yof/QGfHWnobRe+GUIP
X98Uri1KUiiP4RtFtlCr+pEtkZknLWTEgI5k94rBTZdfUd2pGMYFv1uVTOs/oFXL
mwV5BVDqmTroMAkFjin7rpfbdXeHsCUrULnSodVCDIc5w82D7ksDts6oEmybuKkM
Z8LGWsJ3NlhXOzY+EtdvHhmI2vUnbkQw2bSz1z5fpf089pdC4/C7+0W+3KyvWhlX
9ow83oW27lN1s9QW3c8LeMyrfPu7d8OYDSeqgWt9UvDf6mY6M0JTWDiSuZODgsEq
aBfL6D3Ib4T7UUmj4c0iSCsUZa15WpwHW6/GaU4vdmncA5ykdimDchyUxrVACegj
S+d3+3tCa+Sw4Tx24R+SA63V6AuMBJ2qC7KDNr4DbYQ0T07NTXbNppmm00JL0OPu
iJ97G1gB4+RCPd1f8XMfbz+BgV4MdVDH2QCaPvZEVSuGGLZ0YsEMAd8CzZJy0X5F
Jcp5jCyZNrqGU78E70ua1QIR5rUM7TvYcHJ7fGkqRI/zMaj7d9KHYc/cMD/1C0Ej
hQqqZ+d36bx3QmduWn3bg/GPcumRva62Zs7j9hw2zLgdOgvKhRsa1dM0ZwBmqS9M
Po4i1G5UKew3FN48TBwj7bi59wKpOJSXwSJe6NQsyitLSmrtThKqTtmuAtfxxsaU
vH9XpN1qjfg4ZPwqJygFvLJehImZ+Ltb/ZI7Pw31vDwYM22lIV5/+deQFG9clA3l
ZcQaUR4kcDWgwsODjvFDOOpzLnmWc7vMht1Fzxa8CP4rxe3iX6Q/YCV7CfV63MkD
Xz0qnVlaECM4CWk4S29hqnqWHGuLfdoUDbYHrtKcUtRUKqv1qW8zdaUqZ67+r4K3
Amn58vDeGcui42quwBkLkhTVVeDc3MT5/b8xJJmVqnK9wZVj7LO0YcpORs/emIz0
Kcumgu9fJ64d9red6poICPCvvljXN8scYOuRzMUUEpD5TZfsI3fo5+E+Hcn2aPUe
R7mGsoMi9sFAsFDvsFvnpbau6KXX0Awh59IlqZYfcpbGZd0d/TzV5rtp557qVHjB
TN/5/CHM8VjerYWUC3JFWPfIl4mMIszyAKq1R6y+BblsFdFSpBBWOt2IUwh4f16u
DF/4qfHQoo1xuy0jzO/j+sxv5g437sXRtAXOtX0zkZyZd7Sa8/Xm0HRthdt39FrV
a5Q8i4mI/4gRgiA8ltl4MtP3C7XXaKCxIxFalVVZRw+43IBu6MT1d7T5quH4qhNV
PeIZR3xpoGCl+v2Ie5J5ZetjmT4JSuSlL7+oFQ/uTfLQK+vx122GPE/e7f2IkWB9
pXJoMa5G0b0OqwuQZUtxO/OsEQpjC6UJHNqXbuPfszBR+wmh+AsVCbu/ftcUdXU4
7fvYZemSk2UdP9dzifgcISv9cl4d0Yry+PP0BBmNy+owolSjRWuS+LLlNG214W4w
n2h+pBf8zDTYppABZbpZYd9EpW4GhgzK3DWY/O58Uq6KKSxqGfkhGCcHYieypn3m
3kPVFCEeXgE7uwf+HceHbnS2VOgSANp2483ev0cSZqeiar+z6/p+4KEjTOFyw917
e9kTqSnIe4tA/izFZXVkbAfFi5yJrpZPZCL2TTyt1CaqhtbTXG1GxGplTqABn1yr
MEX/AsBDABxUoi+aA+RpnBx8kPn2eUgGvvtDMVwNrPEuizhLZziGoiSAxGndN9La
vlhnCMPwsmZ5YFg/3bMyHGyv09tAtHFlOSa2GRnDFgaxT6oTc9ueQiZD4vJcn36x
oT2GnODBLgx/ndVgbq7GLrEXRlCHud5LFiJ7u1PPLu/IXMQUPLnWWQUa5xcc57lK
dIDVJKQsHPv63PLzA1evK32s3rhskDsryhMwq2tCk1Bmd23yMkn2yeD3Zoknyyk0
GncHloABVwKpW1eyC9yLCpPJ4HEaobs60pFTWLNfsTb1COrrINd08dcCV16jn3JL
h65VUSnwU6G3CweFnZSjjMfC+2Bw8Eb4P5KSOM6JEQUc2GE0Y8ObTxaZCMmwlWCn
PifBqxOBEpmSmf4yqTtkyLHQjWATv3Ug52UmXWtg7gFMOeXKJolcrNDSr+O2RUjr
WX7YtLdPavhEs3aKcjR3F8dnfaURauNPSiqvck7DIwUEvchTJX68+ATC2NPBa7jN
PbBW7BXqla/BkrVpuMIJlCF6BzfFjYU8J6DEKo5EGop9h2Q+2TVn40I6HQRlN7gD
fINIZNABbJOWh1ddI976gurYd5zxeSxO0nZtWX1LoYrhcPvmEnnDr+sToq8Pg62o
1ckL0dOANZ0EBw/oo9Hm57tLjaNKWbNt28cERUWkaOSkYku+vITjUI+/4+EuuNXs
OwEQ5ySWZK39obUFUw+e0E/+2oKFAuGTLLPCye1uKDM7qsoW4cxfHy+dOvp/wgV5
QHoB0uM76aMtLKsBIlPam0Gh+OBS1abk7Br7yaOzhgGKyGEoQXof7poy9IyG3TjZ
tuuA001Ypdx7QVTazvGzZOsyIdYB+VC6UHppLHwkJAk3H9uKW0u9gZbyX6UGYoeA
jt0COj68HK+I9LLlvQgOuZGwurms9tB7Fv1tComKaH83bp9tGYFapnywhabHCUGp
Qy/EGy5jRkjkS0rqf0zpTJ1NR2ycmU7y4tPWlumU/jnvNwJKhHknpCbvIsBuYRIC
q3NQWYAbcZQ9SH4JKIqEPhvHXzui4F9XRWAG0I2vG9Auu8jX7MwL1cIs6qt1AE7S
qiya53/DQVNQwcuPTLdCiGMAvs0t6xWXAx4qb3RKDTfBuSZueD5ruFAeFAgiWGG9
80Bki0JrZI8T2iTqCn8iNwp8RLpZkf/KM8qmb+7tNV1FoT81Q3QJmZ7GBf5gN25o
CITq+z5FYCrrk4kI0gpx7A2gmwPmWGYeGK3tGExqYp1YHb5lqsa+EYzdx2Xnd0Ua
HSiwSMSqRkpdZcHL1omEPOuEFPhDfbMLrnCm7EU137A9B2JoIIOBfShL+YPP2g2O
QAsBH+ZI+rbjgYQnCKQdYNyaooVbBUJ1aEtvWNtYTiq5kETanJdcTauF0oEg+wgt
UF417fSbmwoibjZMqlhiBO7A55nlHEPNQ30L9J31GI+fU73a0SMx7UWFXV2hxmC8
OfYfqJaeSWL3W8OD6uWLh8q/29wjaStxwrP1x8gFRWV7QKOUzHTz6vteR0imvNfO
HZCztji8dxj3GszALwQQduO4mPRYqkLrDF/WxtpzYgvacvxoHKJbwid+Sdq99fvw
c+vTE9QMKoPvU0eN3JHOGZim1x4u3NtPfwsO1STfff4GD+/aTIK3BI3lehzsZyjK
XkTi+bt+hdFaZgur+H39u+KjGqtDxFJlCSy8hXUmXFjTwTVLGTAd6h1YTS0NFmHJ
7LBIl15K0tt77YIE7IySlehKN+QQuyi+4kYad4f7wcf7seb9KKn1Ll59MhcHjfiB
esmNVnCXJ7BFZ6Hk5iVA18NcvITMg6rd0FVCwhXgVHjrYCUWJrDAavDaS+Z2FECk
qjcHa06M2W376LQUP2mjBi//BDRazQuNDVC9vHI0COnDZ7tk74k59YF0HChCtMMo
Qv9RtQ51oTZAc3AdUb2lFGxIX8SdjZCHJPlC3lHVpU8TvCZwHSROniJInYIozIge
F7wNbE8iLPhNJhlrXghSHZAfSdtFCHjBkYAL8dJV6S9N0bMzkIdsAcHLbrOezU7K
x1HVVHBGOLj/9O8UPJwnMa3Ip/fAqEl8cWRQdr+kfFBt4aiV5fIjYqsf94iZ/8Tb
LM1FSkUc7dEUoO4HQV+6e8nlOzkw3IoNYPtskY3WRiSVSB4G53ycq7D3ZXRD5ATR
8wj44chdFJnp4r8wnSmhYE7+KWE2JnvH/fL1uIY+p0OuECiKG04wb2mkCURHZhcA
0mKpbtox7CHb3g7/RAN/yHK9784gTdap3XPBtcdlD2VlhoDSHJ1hM29Xcj8isRJN
73k1O5QPYXN1L/ziFVjQ6T8SmwmYHtALKSEavcA1XEF6wgcdecVCu70hstd/JxgS
76C3K4gU0TfJESAH+7dtS4+c38yfuT0cvhSYOWMt0ieAKGQxwz0fNjhmg9tfBwp6
miB+gxuS7iYnRR2OdvUXZqfo1GYyhHvTBpcRL1PKlHU9tYOgTDRvF1Y7+OEwg55R
vOoyamH8i8Cr/3GFGBoVs4B2BIfXnPwr7X9GTJjfRWKBwNjA41sZvpduQJm/UgQ8
5i30y6tN5/tJrdpI6+QPQxvt7+fwVuI4amQc/NBP06RILIYEpWbX/HavhXGS55Xv
alqD60CNavjAjm69vClAe1m/iCO8ENvXKC3HO7/A6f3eod3pg7Y3pjnnBtorTcGJ
Bmhlu8B0tdm/ul0fRfm5BVPYu2Vj+e33OnIEpPgJSrGDZ+V2ZnQZG3vkbWREaghW
lZGbcZbLem33QOQbh5FA+2qNPe2MpRuDFzCJNRqygWm1VN3eOHXACnRUtbEMhHtZ
zMggy1ikAHJaVz9Lp6kV5iuiiz3SKFV3yB7py4HlfWkDhqeAYQBDRKCwxchxni7i
W3unZ3igo4Q2A9byCWCaGHua3MTgGGM657qiio0YAhDEmcCGPr9ptj7tUlo0ZVAK
JmWZIQ8ZK5ty+u5BAzimLRfiBGsZe/gJOo4MaT2d8bAY3IEZyCkeYTotFAgj13uu
ZOSBq9gGbtOeeQJHiw2oYIHVkNbaLkNJXoaIkMLcC4+7/u7UfH3LAijBdUBJoGsL
IHI9ZgklD5y04C4KKp3FhNgofBkXW2mGrVs9qtEMDLU4JgjMx81GT76raqLKzrDB
j6nBUUYtiIBjkRNOSzGK/tvf+hXhfPJpFx0fisoK9kraISAakBfUbfNYLgf+CSnK
R72kqIXK20UW/uwCi2cFr03NYant+NUHejD5vG7rKMSACMG9YicsVFkjKKkcDPRk
qmsp0C52ogjDjkpYEWBuTujZ+F3rNKfRdCe5bwP0h+ylpCLMuEWmSTKADNulBCot
v838EZx377gdIaJKMZuqelSPZXV+pml2QVLXTgaJfVdzRClm0z6c2GwW9q/whsOJ
Qx94otgdccgNzPv5+ttqOMtb6ME9gEpyFAW2oFk54jMc0o/4XqQV0wOqwLNxlQBO
FtDHSvlzz1Davs0FTZJZgsX3pqgg4cdWI4/sbGGWPDUAoe8rUFhqtzWj0VSJZpdP
qpzm948M46k7RK7CzkRxdmIyBEo9BJ3SLyt/gkkrLJgtbVR1hz+pqqAw9A5oNlLM
Uop4Rnl1iRC2VBQiNSI4FSlJos/2cUaknEju5bkCqyLWHG4W9Hi2tW6pKjC3GCV4
r2Tto/8UHj0jh9jmloy2EdWlsqxV7zHKSOM13X+l/me5r6B7NTDlEglXo56eB2kQ
3Q57lR5w9o0zWOb1n2V/ICiR/Msg9TWkWYCpsoGAxyxssLuSh54DOdLFGWv/gisq
b9cSO6Y97lRbCsreZeBAm6SzpvJhqDVMEg9adUVZJOp+pUs2D+OCfXSaI3vpK+0E
WnjpGjTLR/y7NVRaG/FA7ppMwJuNHbwOw1OXMOBrjNXWOzBHHfXw9Vdx2lNwvVo2
esrscjkb2AcSRptlWJkwQcPcHwyaTd15C//m6l5SAOkcCVOfid4gRAZnxdOb8KsE
vQHAOVRjMtPQXNbYTEnjuL5fnrXAeHZvKrOOBv90ThVgCpbDc7TFdVgNqlMuCLfS
MDYiuRvPtQkhtlLAatco7vu392WPDuVsfdMhBj5kaXO3NBAiUX8U8cdeO7DtC/PW
vgsjpao1t5x3uLEoncIYDMKod41r8YP4Pj3voa3aPsUa6esOkp5He6uo49RwJdhx
rdVdqW3IW6qq85xnUefpHT4zMm+O+gL0V0nt7HkDBW7rumSfYkUpA6Xt/pPOgNJ6
DYz8m5SR1eDhTvraLrgUxcpceIoeb+ED6ea+D55MXoTy39Qkml0trGYfTbO/cxMd
8k15pCsWtca++ikmg7kcQbI8pCNW3KxPtSmdefk7A14Kz7owNBmsjeHOwc6Vy2mC
0Sojz8m5TzlEv664umosXs2fp4yQG6gn1Ib0BOLoz01C5Ac1f9VANKkKPt0FbK+e
kpDXNQbdENZm9ZawqZThE9h71FVDbkhtX832iq0GsIYuN0AyPuG7GqwXJXShiby8
lYLvrXk/8S24r4VctJomtQwVhbpZXl5fp9ovjqbFwrQUvj2/Z24pgWJTjHpQ5pRK
5lXnyD3oYf7z0a7/44tWTioMzDBNhxhS6rpoTPZWa9MIzp/6/4zsVpp25Wi0YkYc
BRmBRHrcZWVhka/5A6cID25fRjkw/G2NOAhsyv8+EnLXX+vM04I0CC+Ax2rlqsmi
gpZOdG/rYgeVDcYL4ambE+Po6YwBjZq5u4GkU6abhHRiUIpGTRBu8SEiAYaNP9we
dhFDecfRFitV0kUwzw4X7DX+CMesQ1hFmGwxDyrTZYi2P+slAn2Qz24a29IHh0/k
lQZYIIE1ZpBpzlHOLa3diB7SOF1lrmpX8PVgNSyfMDR3uYmgB/ilSU/2IIYI0l9T
G75/awlkvahnD6XDTj40Fprp+QwaUDG6Z+4iORqHktJAceHDq3AwG95TjmjHwd/x
Y41hZegJANdMbkHtB//qluupodmrW6H9SvzxKqSP6Cy1CaDOwkrRdKDydabCuqWf
Le0ckPCHDvq63zopBfWsrb9FZ1HtO5jQRdDWMeMErTXxGxttpR9DY7aAo3m4ADJZ
xrcbPR8nXABWZugn41LgYg+Yoz4JzstidODjoOP4XuNux5zsQTFI6OSHXf/R+pDX
mxvhworBaskdTEr5/v+roM1h0/ssPWByMFc4pwR6pH1QSulia1zsZhNLgnWAsWQy
7DJwZ3oAC3y3hX9HGeDWCSgvngs5WHsiwPpGYu2J9g304TqLDJqWEx8uIn3Y5Hpf
mxTItMMmtm06yJ/ZKi7GJijg+lbxlFMAXNe87XycmGEN8o5/Nw8GLFll+POaur/k
4iVQJ5mZlD/5WgpISX1nnt2DWCfKzthGyc5zSAcsbKYfmRapLzGrDd4xbfXwYeGl
N1Zs/ZqvZkx/wqcnFjqRtD+ATdedtPsfHwgOl3nUNVNwJXKhn367DLtV6KPGPe8h
jmlhKF4nYi1wsxd1rB1knaY9yFiXkcdiW2WJReEwKm98Ff45o2u3qJhZv6KcMLsX
aR1bB+eqP+ZyVhaGjPOQw1Ch90TYHruNFdq2Fzsu2UbDMDFroyJoJmcr9FJrTmSR
rxdJHJ10ZU3Ux2DMBmS3TLFzEGuUIUahBU6sIL8QSJ07Jt5Ktj1TAiIjWwUNIwon
vfVDnN7fs9imtm9OrxhXAMghaLw87AgeooYhDbCd4VNspH2JFMr/thbnnU51ktwm
/+zr6O5idZP5zAq39Witud5j18495mCvHwAS1qnlHHQNEfwSwtNAHOaIWdHBJ84B
8CyburdNXG4piPIb4FKgDMGOgj3P8UifTubwnWWR1fDpQW1sn+MtVbgo0UrAf1ld
+TIqy7UiRT34fVaM5AKeNNTa9uqWcE+VPAarfxqae7JXLSOhK4ruzGIdYAfmIqiq
wObsjnXCt+roqJUt2+lZBzm9KSJOkSrz+RxdYYEXjy9SqWSQx3xzFSqgkJlHo7h5
OqFzbt3sZyZhIfbf4y0XfyLY7i8yLnuP2GHVWe3TzIG6iQRW86u7WdezG+mDR+1l
+9SdDu1rHDoFxseTtfcaYFz3Wm51BYfiVNlNHlrfUEtuYk8Z3wKFzKL1kwA5Yb2F
MpUpsOWjehYfRftaPsFaGriwsBTkQaFbIBMTrufRycxy05A26Y+/PsNfWSbe+ULq
jBgzSmRHBhcSpO6IJbWkr69Zn9djnp6FyX2S5yUn84qqLpWpigeXNvePr9K8P80P
6orRXMHhTLtHRzmrWDuXv62owA8VXyAY2zMXvGg3DKWw+uJmMe+lbWofEtc4fTh4
CkFBKGNVZR/64/AsKQ+C2z6enZsqBPGeAHNapFVwXy/Wp1Aai4IF5aI7aVcZyMm4
RyaS985SVwZYOoUvyodRD4shNqQ7XLZcvFK0lhO73tONtGCJ0Mmn4QU+ewbUItlw
EYH7HgEX6kn5Q+BJWuB5pVbSfe4JShDQwbRo+glcux2EGeRPvN5YmvRXLmThRDmj
15WhnSGxqaJQJq1/9lbs/QNjHCiCBUvZcVeqiat26gE0eSircvl4mhau+8dxj60q
O8N3oZQ9QZa73uUdWxAxGaBH324wiO0caCJE08r2CPuVhiX9eShlmRm+Z7wz2LU9
LtnDaADVGctB834UDenUeHwqzkMLMny2YA//d2wQ8Q5psE3W+J5M6/WIivPbEsPL
j+05RY6VrlRyaJ1s7JgiGgHzyDPawCIKZ9WEhBd8WB48b5l8/9RsbBJkUnzKTRmp
5HO68f55lwr9KmZdFUcgRqBcHbUBSZrstBj/iJzEXgS+Y6JK/LAsv0ZUROmwDPXO
Z+9QzRvXoscrECY7aBV6esYHG3q/fE7PFakbcb3D3rSsS1jL8dza61bcQezHLVpO
ADkRUZWfIln/zR4BXz3vp7C3fo47jWhUQx29prmITgvoXv/QfeDUEyqVMkXjcFdn
boNJb3tzqGOqWuHAODc3tUY1rlqgeKWGg7e0Vl2w2CIrbToweBhKBARecNrSHPH2
hPGp1UtZhTHmB/HzN3RMY5aufQ9sejaONu9nL2vfOzTDv6F2+Jlq8PXEHrR+9SsA
ZKz6rp9qJ6viHJJ1zRqBrMBfHoePKpyt7UPGCp/66a7sYLBBUM/96I8xiOCPM++7
x1Ti6u1Wk5t0vKjTRovtUHH7wrqUIzCBb43656mc+oaXyD4NKpEDxMJR049LEaeU
BvUvZXNhk95/1UaUjfChyJIeojz9WAKUNVHMCI6D6Ifh67lnzr6c2pPfG/ZpyLjM
QVoLKe303BKYzyuBkP3V+21ygUFIiAi7vbpupjUMrSS6izYi3aRPQVL6OKyprd9I
q/7H5OqbHC3W4ORPysV/u6q6KwlG0+a6W2e87ihpn3EZ7cQNCZYuSskfTqjjk693
ikaUS8eOpGlEdqwVgZSJPdtENsr57P9xM4l5Vcqw81rR2ivWoL16hkaPpn/Jw//I
QqUMFbDJgrEgZFenLoaW0/aIqDNlQwAJPJTONGKYntFCAQQZgU0fiC9M3Iu0Cs/g
H5Yb2LNGF/mVcogA/1LvVImy4TdZzPlYb54Dd0cc7HrlF08uHUSrEImu7CsTHgel
7phJBumy4ulKNl6z2U3pwKcCdeMtRGTqHXkLa+DaU0xjrRhXs3iAo5lFcUCW57LM
HSyzgynFaltycR/9BiFQurzMOaxtI7o+FEMbgPQKiShqXsbw+BsmBa22G6bcjPlh
ag1Uli4CidmviHkUKMq9Ubfq5wUYxjmtkrbMtzAkPFfmVjSS6GFJ0mCi/y8m6cWW
FYkhcHmPMxGO3k7aCmAmSzx4TF2+uu/xMHl/bT6i6bCiZoNnFlzyogCjPA30gk9p
VAqzunte39uHQjJQUmLg4VrBPQs7pBf9UP44McvuDHQE5H+tQSSg9CLKQD9XIEGE
PTErioD0TTfqrMH9pQxPQzVjfRyFmeEc/QLlcndZBTyEpJYvR1HSofGzaPxX2bxk
N52twhATnzd8bfxTm0CRTjWrQftnTsCFsUA48ZgAYlRcq5Z9erCxtHc8Q13VMUDW
2Cn+QWElf5UHnBsnpeVSzvvmJ4Ht0gV7s3iPBx86twJ75Sco2zEEjMyd3LRimx5w
uSnKKa7X9acpWZKKTrq3WsrH9wctBBGMtBYTbTW/l/l4ZETyiVYn2aEOM7qq13Dj
S8CGLxg71egjKZ7Ehsw1vNUyX8Id4V4YbmT7bMD4Di2zPDb10VWKZ12INT/33oYi
WTo5hAGmt6GiW3S3OEZbW+KX4whpIkBnpFep7JA02/Qsr0EwGV2pJGZk0SrDWCLb
MVi0TfetedbAa3jYMK5AMwrIsj04IIpHi6Q9pJpmVELeCs50roY6bF378Hi/KHb7
USZ1duzYd1IgREoQJ/Y7YC1xqvS12Cq1bkMwGNp3kS+Xqh1Q8d/X1h38xfWNBfO/
zXOYONYErsGA15so3xiJxJl5mpQ2mLb4rHUK+gYCXeQv7nJIybvUFcjOaNisq9zE
ypB3dhcYgeYbfQQXnlKFBFBYJQ5SkL3ZBCDFBqHgFDtdnudjHvdH7veKMMrCP/3R
ddB3rYSdl0Kg2TPReDD7+Am1NdpCluWwWNfdm/foMLu0NPsg8PjgYJoBo5uc6vWf
7LR96pMBsg9Jf/QiTdQ1zBC6QA73it4H3l7b0u+x/00QLBza3eDgBNmOTKLsJXWP
vAMeDPf4/O7gHAqN/5RcWImU2TE0CExI0oh3nxLgDKc/NqIHR6llmVe/lmDuhIbN
3EVy8Bgq/wxYYDt+3FGmCDlMDh1HZkCQg3MWls6zxVqo9JDJWpC2ZOCX+2DHhSq1
wQlPu5MKk7ctX7w27F9piENcRAnbXrnYGeFq9pNScbtE9tQK9SYvaUg8oDieguPl
nX9tLZwz4IFs5kSplzQmfd2NU217YbScil5DHXYlekZejp0/gWg22CV6oiB/822O
GXxow/FRB+fx6hHxaQIaTvCavtC3Nax4xQ/2GfFV5RWTCflf6T02dWLAYxkLP8pD
GPNDaxAcW5Xe308XzzvvhmjCgwa5u3LpKObO7WtweJMWoB4rnh0BTeBVPhikUcNO
LA246IkPzypTJ08YN3uIHWpNtn1DcPCMUoe3x/0+mnWwRCXeJNCYdbt6Radc/wNx
PTM0H585nEHCxqy1NfI3ZnrqVePIfqRfmWTWocpOfi5i0y3Q9i9GjDUJ0j1bLLio
d84h3NhfGErdzHPI715c7nX8dA5pNU/whRTO1k1qfNmOXPe/ZlblWEwX+PbqlTrw
K4HO3uh2yHo/+mPM698WA1FpWfO5jkTVPkYyeLDFFPeTcbx08m5J1HiPEU1bLma7
b1s3CSrUr6AuHddz2hSy8UcPA0pav/v6hPfKv4dmH4wC6LJMF5qtCakMWtRkdPOS
z9AtJOgHyPLZZI8/GkIJ1BAL/eYozEWRHm5qFU7fAcb4SQpuU5nahu1CkWjA3cpb
GySHtyCFekLUPFA50kWXNZxR+0eU5q1GdUP2iNLrWiGn/iowsgpcXvl9Hk8q/JG0
YlpVrBI/YKs+3qr19/U72KrXIi5erVxXN/R73OlK1bLMruEwPjyncIAoOrsOODOz
Gzk2jkUTdPhpNSqiKq0gX7uyCpzXIGUjoRioE0VkMSrHuuDJLokU2DuWYq4cLMW+
llHQPPojC3OaNmSxZjAITwQ8MogQ24WLGUw+3d7gVsvOzDTcSMomIWdZsV+7cZvH
VKWljoU97t9Oshpo1+hEFNCtbrIX0IHxAqKiR0ps/7eXLavSypjwtmYuny16xSWS
rf2Kk8na0IQaXP5VsQctnB3nW9mfjY+UUNfPVQMp5oDTBnw6s5tVHwz9p+rtmPxB
GN9ruQlH34HqrzN5zcqrNgyYr4LQRsPd8noY9OZlJe4gWXxyyNxDQXB/4cQNo3F+
b4Hhc2SfStqBZ2AttVdqiwiK3EP1cDOwxjhe6JT/sikrlGM/NIqT3fHziyOFihG6
spM6JRN5WEzHTC4uIxKWfN2t5vFtdg6kUA0nCTX1brIDhMFwwYKC1kc6EmMHpk25
zTEG1v2mX8rIDC/tjJ/gJN+ErGwIfg5myvus7a7j8EsFfPuM6OcZgESRlx2yFOAN
Tax7CnYNy9OeShO69M5HfmdPxR+8zbV2WFrpPGlKs6mvbuIHqA/MmaNokkI9PUIe
38bKCE/9tRR2xQYCa2AqZJFxVHBn7MwmlWrfQJmPOgHdRAYbbAxHdrVKM1IqFmGs
u/GztiDKaHdnhKpnN0NhYDzKhGOtoHNZgX01Z6jqA2uIDzSTUVof/pj+9vdaQqjm
tiYO6UxQxIJUJuBUjCUsBEdiGoTdAnDHJ1FbRdGgB+249javPVGqurjfprjgHxQT
v5ihPkSwBeLFN7WcqLzA5Nl4CuDfhcSeNIYU/3eVdlElWk9e5jtcz5uK0KBdtdIu
AokQO+MmxcXPw1oShvKDANsAM8JxZq6nOo6Ni0sMECPlhBeqi++Q7Z0vkV/EOM4h
KmZ+M+bddx4a1qwaQqReHJr8b3xo3Wj0ao5oXIR3wJubN4uIG5FMEyLiigKTjqz8
/DlbHJONyHkVO09R+E7gDF83gFgS1eI9bpT40exRi+Ke/A/iKAobZjS6llrvyWuF
239MPWqGqp+/TH4gxBNLnL3z6s/Yl78rDNM4TNvjIvhTvioFLzZpPSZBf864YBGh
nE3joueUR+meY00Ke+IOl7rb53j8G6BVm+cwb2KtqZLNpEFjh5eTTmguxe69AVvH
rRyCeqknG8kg79d3K19QtPA5pVQ6sgy0DEczl17tv6qoqxbYOD8susyuY/0Sq6Ko
lTKzRVQ+r6DPuNgd17XvNK+ES3/oEdlbp9x9s8NINVHmwOeRCliA8pjRT8rN2SVk
YhByd+4DZRc4ISP3uU6AegxkFc6c3u78WBEi3uGYXCVFXdtKtwYuRiYBvp51oEnr
prAvhegML9wrvc4BGjmczdinhJx3K7ANOQK3KGaTkbdKdqzCHIiq/Bfv66bBmWRs
xE7uJoMEzil+c4KlN4ImoPHhirsJEt594aRJIqBt+aRFZDxVXhqN3sPf2UbYAbX6
mIYZ49wToWNg/mod4nnj3CNx8Mh369T1VkVkUg3QSnF2bTPH85VaxNRjP2ykMRjc
0lCHTdGTcNCa2uQnx1kF1cwq0FaB9x7Q7jaH/k94iwjZHcnr1wIpMCZX6qphd5Sz
gGVpyG9CgXpB4WiLJQ44cNGspw2G7vzOf+tM7MkcdjzCOoMoKhMxMwPmYRMy4j3Z
uZyZfhbzYMNyoFT7zivlHDfrMKZ22wO8zLp/ScIUVXzjsMPhk/bBv5+PM4kQH5nE
Fg/7PVzXQ8kd9XBWayPBstSkAnNCdwd2L204BbhCpUTgTHa0Vys6uPW46UXDkANW
Ahmamz9j84S9y3F9bJ8we5qBHKxGaGfdn2Gjib9HAsr8WFwmvwGwDRptU7cOWLpm
HJEea7d1mxsGRq7e++I3WQZ0Bi/MjWth2ixd4rqQt9YOnVcNhZgJy1UW4tpvloZy
zwyHIBwRxhtw2hKiHrJBOGDI8pPHWOC3hrpYtBI+5H7CxuQfRbY8lefPVuM7pfzA
DFfr178PVDbaIWc4yy8xhw6JcAOY/2WPq8jIZFOLdpcu8uuMYXocDjZg+gZfF4+B
rfXQrVwYEK9RZpTRSOHU7vcyft/izekqDcKh8p1ehMYlSMPLKu3ROouSZoo5nGL0
tIuvOWEI4TbXwWjF4rExE+OnBAHlAfmzV2B3RR5b1EaZ1Vsjedme8BsNXUKwlLcR
v8CdGvmRVG4tvD2GJPlpNYRDlRn+APD+i04oD7dWW5AUIPydKlPO6vc33GXrK2Q4
ZYu8aRdJStnvYjcVcUrt307dBVhN5UWA2JT1LW8cyAjOYcmddtY73sZsdPEblZkX
Tf/s0Wzj2IP214yU4VL51QGvAE5s4SNMam+W+cWO7RWwXWMUlQvLRmuEikXXT4yj
AaD2PkLkC0OJW6PmrnRVtLkalh8OlhxegTgMC1d7YWhLtdWJIMtYXbTUSQMIpR0j
yyLzEpUUyXNYIYfUaGMBYH4fGCCauMiHAJ5LmnqZq6Q9FG01tWvMqJdbd0ZyNNMP
9yY7z6/Kv9btxjRfSXJ6fd40ifXEoR872Epe9AqwejhlXqrM/R/VW1Lqjz5yQmyE
bjLrb8jQY+bopIxkxitWYt4CoSYFXvYqICTQSj1vefeMDzZsjOjB4NJGVxNUuM83
I8pUYurpcOV4sGtaHS6Y6qSCuBz7qO+oTzQjXjc+r6IrfvT0cwICcSR9RYdMwcQd
vUEdFOfC+7VJWx9T871ImDVervq8YeD+VCDDcHd6L05kpcXAtT2YAgHOxBd31hfh
wDe78gYl68L18VOn7R7hU+A+JNgcgz+Scph9/j4WJw7rG0lZWvqCSD03sUOj+X24
IndkREJzMRwFwNhC3pOzG3KvvcdoUyMg1cC/w9EBjp3cuMblyoE3EYnuFBhgqnuf
RKudeQFjM2lkXmSrDzsNfQKItKAM2gCwrOSGY42rfe3lzykLmLkI5oEcKIzqv/La
6g+Qt4aX0Ha9sxxUhiBUK3YRCrbuNpuefTDSxdDQBHma446sa0lyJtu1y7aMwNSB
`protect END_PROTECTED
