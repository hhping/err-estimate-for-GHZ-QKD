`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4CZdxpsTsLSRZI2F4bRHV/Z1OLr61mv/vw55f2AYnbn9tezyDL0+UwNNTWBfRNG/
2Kp8jh/FI7KSqtBOVsbG2g+jVCSajOqapAFkBcZQfjRDgyCs2gBoogD0R7J28iRA
w8qm/icd/shnhanoPZek/tfRvIsLBDhs6bn3dEC4vuuWDfJVYudXC1xdcqygYAK2
fk06MY6XiltJGi5c54pD+fCWpoKPN9pSdqARLdwp+/TCnEAd17ESkFVGorExP9Is
AwAtBcEMx///DLNlqLbqBUd8bVm1P1xRzQMkQxhd7pUSqjbhLWCeHiO9jkwIX0fd
S5sqkja7smMCzUCdCp/q1UCZh/HJ+jH1KqrEyX1WkS05FFy3IRoXzaly29yrSy1h
vNwPyimScU6NBLrV/CRywG27e4VB69mklBbLue/tZNqJG2RR8KTW1uLQSQ0OqEWh
aX/jkEJJCf5WY86weyYVZCJBvqo3myjhTXRL8vynBA4yCskwr9biYsU9hXfcqIZP
IPDtzdV8K/B+dmy0oCIwcawvXbU6kEAqcsmqWxFBgd5RI3/BzIMVdMkp1vT5QdER
jvttJ+AVaa9Sbe/ABs8SHEI1jtlI1Jek4rVgfsA8CKRrdnsj2wcbOv7qhQA26CwL
PeAeMB2A3/OGHG9cVaHrv211R5OefwDlGReNAbdplRB+HN/769US36SLfeQX1+S2
l6t04LbTav87d9RGLTPYk3dp/OI1eqvYceCM4M6HzvuUEbtmRIEsIDp82/wsqHTD
2MnD8RPyE8OMHK4FbSy4r+9QvrCZecdkeGg4EOtgSKbFUHjjzQq6n6qoRxXbRJWD
rzUDalrEdPUfAOZkBAUgkZp8IDT81MJQuJUPUwP7XYgSFcaVfwWn8crUg8uEmTCi
qL9sDMu0qDrNCU15ItR4/z2sG9D7yQHH1B79/zvqUp9MoDsQWSPJO/nEsebQCDLF
6cCNzetS4vUl2se2kQpjr7BV/xUqKP5wQwvn2mktiwf5280yYbV/88bUHEZvaGSG
hq3j/AbcLf3qegKq/xHmRVZT6DJc0E2ZnQPzdMZMuEd+TqJfzoq/2xn0KM1meUwF
xXshEd3zkEm2gB8Vh8WFBAUeZwBtwQpT11CWYRNBtam9oiV+EhLors9EaqTaVX3u
pBy/8uqToJDMdivyvY7ESKzxB44JY2Dc55kSHik8oGsZhebt1NzHT68B9QViLqrd
y6nc/gtjZQs9xUJMxcq2BoDylNQWQDvnaUEAv2EP9nhWWDbZx+hje83KlKRcgQ8u
GwyebHAk3mg1/5cIuuEGn6oE2IiGFkcSwNQZE7IcieLysp49IYIieV84Ks9VmV2U
lxs6ok1ggkbbC0jygq32hZs3X+gaJlc4GCdfFNllR3L5c+EdexuTYgwe+LDfYjII
VvnkJL1sVmlMeA2QNEEoE68pSm+POgL4YzedN0S9runIKm1CjZdr5NL7J/ZRYDbJ
FrsfG9FUrkoKO4uovQ5o2Wqp3KBeeURyUtYfCX4lCGfnGSaAchGk6zR2A1klxJ6L
`protect END_PROTECTED
