`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POKmD1G9vIr5boMElvGJv8DWPW1bUxQCliPcYvqI4vB5t8jSJTRTb2mgqYyYNCr6
RV6Hqa5jv7ue+IobUJOssDKlVUSeb96Ip7lIibkA2AouwlPmswsm2fC4i9fIxUKL
dIBrYqclpzMlkF0vR2BT5GPNfGQtEjpLNLcIq4fRg0RZxKWGIcUVjNWhFFwLrbrG
TrK9oBbWs47qIRRXkRkHgpaBA4fl/+skfhfBihpMfSkEvFk1bV5TJLx5bddg1ra3
bMDoj0xVtmRz89u++a/3rfAsW3n04X4HcRLAC+GfOqZj7yX62fc8dndRZ6U9ht5n
i3YpSrpdTBrixrjCp4q2n/mksYB6UevUCmL8QjrHHX14+tRHaESwf2c8UzgpcQYZ
PoPmTy9fjcUhpubOTRVHuasUt6Li1eYydpEVJUnJRB94oyEc9mB4afHmZkgrwovC
uik5l9Lz0ndM/HRhzXdEtw==
`protect END_PROTECTED
