`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QTJDCl7i7Ub00P3FQjtQrjaAB0yMomiTnpxPDxTdeJ98vlmEYlZPNRl6NFkRcNxT
CSSGawVM1rabro6VTe7rNx9GU3iYhOXQuIEGEtPF5UqO80TNA2lFpWE+KSFPHid5
mtGjwNQniFoFhniqXudSqpopBkE0Nr8Ok857to6LSEJC4fNl0Wet8eQsmn5ERDs1
K2K2BMnDxDcPDJsa7//++DPAzSqOCJulh4P3le6HDG+b8Iuk2WRqAk+EsXwz1F8U
wf1XmyYBzH0mdIXOZnfVw9iGk0itX+K5oRWannJcVQ+32WASVc5jcB7uFA/UteZ6
eyK8J5JGWrVByXoq0L/tcjPXBRC43zR1dDaVJ7JgsCyX/NOWbWLbiwwRLdy9c5Nu
Hxo4mMDOi5m1WEFI6BR1TD8a+38An1w/GNl/t+L+AK8+YK6reWRmADjLFTKakiBf
yxMeFH5o5gCRQB7tIayxNqFNvyn4H2JYKD2O7nriZDHx9GrKerJonWTtA2h+Q4VO
B4uXMtzURx8UG1Qk54kit36yXW/9RT1QiVG6cX9QgCs9jwAnxpZJTKY5TOTv4QmB
24ycIip3icuZD8zLkeQkNH0XptKLl6lRXYoAc/+9lA5JS9Yf+YJoINJp0a5ER2JO
gZvdg0vbJS/oXU3Dqd7YVaRMqeinsCQfGPOLmaG2pgOL9SBi8Xsj5y9avKYThUuX
lYVo7t4zTn/Bfyah7P9IA8BCNCcKCcN2VNoQ42nI18sfVkZpIwEOUV9JtmPu9HUl
H9CVWEPHENNbi5eHfex6Pe//Nyv+7O7pVAzXGAEK/bb5WccuAArPqOBcy0EW0+pF
bLxA7gfLO/89aU7cGIjGWHFsT7o7Wp3HUSUc43Oenram6e4//YLXy4DpvNgcnky2
920x3DWsjXoiJLsV/OgCjyRon5/KXPbr1XQMxPDMV6tC5UiFwiqU3C1qtzlLzmdk
Ao5pw0dBzM/VSnt6ERe937y7Xguy2hLmvoVBCDdk2hfY8wRjyLDDBrrspf/ijlEY
s+utjLRz1/U/wrWGUbbolyHhZ7qZIqOhxcGgmXwEUXKiC78ldBD5Ikww4Ua/njLE
n40riqsxcadjKwrdbqK0JVCnnKSFQLy1TW9Mz9bqytEXRrWLnE5PnjZqKfE+wuQl
8OtblIuoL2FbX6jP2CWrM47olTxifgq+nK4GSFsacxCLYxdqnH1xa2/imasRaG+L
/w5sRo1ULdm72DqRYfz+oUGzO7fraMZ1jrIU/UqEiHTNeX1uJrODaULseUgWiFvy
pvLFMLPlUv6RSLB9qYopo6TWIxRer2BPr8uRB9k/oewJdWdppH3cNb8MWSAAAHUc
+fTlYT1f8BrLHK9LTbFiHVXPBNK47RGu2q1jD1J0A/tdxSbFHRRwYkXd5EQx6/lZ
nAHzGj5Ry3kLMsK8X8rfLQlC8C3fIwN3PapjPegeAwU1SU5Q4D1zb8olYvSMEBDv
oKcGz9LBgL/xi5iGTA/OSqfNRUq/y79L/T7fykMnc+za9LyDIHTsuaHJwZJPwKTb
zYf7sGaxySOdqTCyv+iWocMsmO35U1DARI2xsihkITJGdYfpZD7IMR/tyDL11Fhm
vNImsoRmK75HzdhIwIOTLm3VncELThv5I2QuFxUJ68gYKjr5uYGjsDBVvft2Wpd8
LfhQZq88H2FrR1VZbnL7qYa0DZyJug4Vh0PYpeY5pyEl542CulKSN43I54FkB75p
LhHaZZnwuDdBzVko4RAKGdWdsZQ16XKqRLClkzJMPBHfAzuKY1AxD+eHr3ciNc1D
yynVDIEu1zkUd+SIYGSwcN4gQ2llDuPtt6m4xr8m1iD+ZDsxhrD+BPZiO3GiRhGi
0UqkyOcwAyWQXXZh9dh1QqgbLguiS2nmiH+Ath80T1hleuanq5mImt1LHixTrGfa
`protect END_PROTECTED
