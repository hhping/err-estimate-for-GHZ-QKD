`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXo68uz3TJNVs4i/k6YVBvIbSftssOinoELLj5r44gE5Xps29tVQUdAQDWkO/3ud
uSh3W686rIgijKPRW4ygVMUe3XlT6dkWQ2SRAJtxWu7MleEPiVFmm6BAXGWQRJKT
Irbx0dLJ5P0GKjR89XyZrfRdN/2ENm6CX4CmWC21SI/yZGgk5v9m15ZE2Q3YsWAT
RShn4Sz+asxyPMOOayHePdg/3hqP9j+2hIPuOr7sSaneSmy/UK37qauG3GJJ3WSy
7FubfQj2Brz8TqJQYfAtZxn6lKMcnZyxKLfi7pHOGODFl7H7Rg+s3jR4RRN35Z0H
Q23km6ngDwEaK9aPkkqfkTzh3QMHRG0gRjVNv5pVoXQ=
`protect END_PROTECTED
