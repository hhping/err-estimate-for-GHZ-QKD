`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWmGWfi/NHuNiN+ecSY+v3kfNoeIA+/z8a0+7oxbyvV7FSh8HNLVeyHqqLZbYxS0
Irirjq9xoZzwGrs9AhY4UMRdhcK6yR6bri5XTnB4BVozpWZEbtoNZQaXpjLPK34D
OA3t8mdETnDU4g0xGMHlIrI66pKlKC7hr0YlkgA5tieqCRvwKoh5WgLybChSlmCl
JJmLUCMTaXMvebxb2xZnaR09RBpryy157h8680iTOdJKpynXM/sQsgMTKjel8jK7
3zWYfUgdJ0sAC0Jcd31dnAGjw6voL+kOtqkQh6xCtVqKLVL8sd9V+HtrRgIFw03C
Jij3xo37WH4LeL7LY7v8aRluVpLHJ7XhOA6t4K7w1IVjC7+ZZhYDGDoaaeHXz3vL
4gvK0mHU+pz6HFGb2wQS+KjRRZV1ebbbDoGLjzzeX7n+J67uhdKUQTTP1jVvLsUW
1Z0/OjTYMDHMyimSwiShNva09jKe1uu+yDt2C0DqyWRAQguZmmBmlBUIrlF+GA30
Qu3XDBFE0mMmzs6/vccFpCOYqh0DJoJefE7frXXY/INQvhyWN9KtYEwTOtGA/3DG
/BGJuX9isNN6v9D3Lj/kaXnM5rCymSkh+x8f72VYUQI9VPZ/R6BFM91jp280YMGp
uikPkowk1cVxDsOpwe3x3SZpw/oVKb16h6sqHL8oZkZogYgth1L8KTCdaxcilnjn
mP0LfMW0Bb9pOjnrGyhsl5SWXshQNbg4sG1ZB4rfErhvMikDrJdfHet+UCGxdPRJ
HjY8B0ear5H/xeyxllwZDLtj6ySpCMyr953QhqjJrU1Q791Au+1914u8eEBWXUC8
aHIu3+3VIJ8OvPamHVE7VOpfB7LtQ5Fq5QUPK8SvHQ2yoy3G0jQ3OWDrVtgd4Yz4
Hi+v+7xi4dRs5pXHSwVp+aH6v/X2egzsSeuvpVg0poPGc+Px45f6JhmgG4cucWJB
Rh+rpZ7kWM+HEjTdIEz7igqISrsirz2ZDawG4cIo2DO7PQgvpY1xKjphAOFt+soe
AI7jwEABj2C3VJINiTCwf+q27/ZY9zVs/w/Kg91lvpV+xq/+9KWaXa+D64t4OVoY
j0LDpgs66kzT1YTzOAsEiQhX8adqF5AfO4rMTJvqt3oHzAaksgCxOII573giiyDL
ShbLU2IkGftp790ewrebESf69ThVllzuOqIT4doqjH7W8amHC6RmVKtnfZ8pt063
F7cRxXV2n7Qc3gxeH58+Z4CZhd6uTYB12cmyVTuP6TBfMZhl29XHWLWkSK6snp7P
OGEU2z7ryOQjv4Hfj2fxkOXyu8ndmMvArP9ymPXzSCgOMHGCeR7pUOKqLmbyWQ/S
jvGSLk8R4ptxH07MYFstz4bMsiq6KRwR2fjDzEP0UBX0F3dl87s9oNOxd4G7XkAr
uHR+ZI/935B6n7n7Eqoo9dMdYnH93vXw6aifTcfoNnmGpvXfOvzQh4eZJHz7v4SL
6Gb8UEe2HKuLahs3v6eMDy3BZTJNZ/gqC3fGyADRNSnRvPzpcIHzyuf1wTzW4izb
mm8VstjT9KcrNrqZDcM49Nrnyyb3GutgewjzKZAMAdKhBXzM8PDgL1JY65znjAWs
OEsUFdhAHjUypkQkeRjcSeUn0b1ix+HjQFv4XfxQ+ICaWJW8dkgqDwQCMtLResMF
VE9RJs37BA3W/sPuiuGku20qFkH9dSSKfJ6uh90nJBlrUXmQiIRJyFiMW/3/cPsh
i7Qv3meo1LTUDRfCJc+qNOqFsGzbh6lks5TlSGC4fQ9fhDy4Fic+gt0CHCN3VJ2k
wD0GKsSWHZTD6xcnfRdlHxjvVtlDnX+is5Ncyro+ymocK4pxUBGbONOfrLGtL4ee
2lhXLa7+ThEuZXwp4NAZYv3GEPmmHelUzYhyR4O4JJtkhGvhTo5jgWQezO/PLBAa
jX+/HakmL+2YzACATucAkQVhSuJGpJkoY/YtYdfJbF15bm/uvSYNjbLfUrJNygIM
x3rhtXQJD72L048pTOVBDjBNdI2QDJH4Gws3wrJ+3hXbOgTZ5vrcglqTQ25AdQAT
O8cIIGt93irPMH82X98nO7n7coYPzKprDfunqyW2jK5rSVqdQGZ7Si6g9rfG2Hgr
/VZN7hw/4qHsYdy81u8v1oGf+kPoNxkPBltJLTNQBC9MeQDqXfU5/JUQIEQP/f63
SiSFxZVJDWP2qXn2vV3Bx1xCqm5XBx0kYmswhFNHYmYJz/vu32Zp8rTc86MnNLKV
hPq2IABJXM5ZLV/RBEipdk04y9xp3VYatP4t8wvrLJiqisOVM7zK23q3Vwd4hiiL
9/y6h1NpUukzuJ9RtPg5aCKlVnWszg8dugVQ13ZbwXNwD/9+dl5qoszBiA2u6W0R
Wm4/LWZjiOeCjEBpmlx4e06rY2PrBJ4cxaFxO8nG44tH0Vrt43WMcVMHvBj9TeK3
vh+35gdqw/eU8oOAFjdmSJy9NXeU4UWQ+wq8zwkG+n2T4zugRFzepueGxInDJMBc
`protect END_PROTECTED
