`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7IT83IGjt2Pi4uB4Jx4ZORd5oLKbT6w9LSBFL/YqI42IVo2cZMTqwDoskW81+mq
II4E1hHLuoaBPlvVEZAiIsMDoV90Ly4tFKSnxzIgTza57WQs+aUMkbgI+z/qKyqW
aDO74KwqLQjsU6v3rEu3PHRbSmxXawnBXS61xKqXDYVR55Wzv8zaHdeVl/P+I7gw
rQgNbfdJ/DCKrCgyHe8/nXRwWdaxWq404gHlYHya3qwV+1VB745neQXlpGOLuPaV
QH25kbvOm4yXpkfzMK46kAWoXwaJGw2WvZgrqE60QhLBHrAzW6V4jQJJP6Kdbcp/
U+yj/cCa4hSXHrv3I+tEPGG19REQNIDDRwQfGA3zs4Lf6pOraB7XXIDdpf9CvLSz
C+S2FW8/hgR+g8cc+pnaVsFgoKeH7oeC0ZX87nrd/aWr7IcJ+XlPxzAYK0C6ZUUZ
hogZkJgh5cE2jY1XTuUPEnfVEg/i+z3D3NpmFdWXWydzDNDlgIP7f1/xd555WE/7
NzK8vkV7mZBS2BpoU1xWFAn3mSqVDDbzb3VSuSTxG2Y9qwg1Aw3szqFoIFhXWang
wKdvTDnG20HSsVT9geRiIQscPDRrXyBljgK1Xmp2A7adxckS8HMDpo1jrCUasBru
/8rJ9ogg+wUFW10f8egW9THnsqRsjvcny/FrFvmaPJKpciM9wVIiBpsJduVU9z2F
bPSmbckN8M0GzXdEjjWdYdOYrH++BYj3YX7+hdPidbgsftcP8YxbTVSxYl0Nlyww
QpGIZuwMD4zxxQTl0d3BsLrpmJmvvvlonCvQV5bVwBVndbItARUaFwSmiAQCzCh2
38vU32m0M7/1Xfh4cBCo4B01nb0alY9TMqZxX1cRYqtViDlS5WByvlFWJnPi7N4B
UVhdlzV6h5Fom5W6pViyszVIfheFEJrYG0UVyLIzh3E/vOXQW9KzCXtNnUU9whhD
v1LMJK46wFJOh+OprfYm5whyXBk42oRlaSsgPSDM2YDsor5euZpSE1AXs/AZVe+I
3D0owc5eCOESvLXUsEF3v9PHL4xULUun5doPuOUVKUvQkaDmPxD0v2/txtZunHIS
bn389Ec/ytOrINPrysS65QWGlvmopWXhFw6RmZKnoHcwhI0O2/fa4HMAKZu7FnNv
S6C0EcpJc0HDSQMPA3oybM+MIIxC24dbc4oVHUZMrvFTsQ1QntKuEINnuPiNB32V
Tn5Ga2optuC2CjoqiyJHK6HpDbNQv0TQg3TxlYSa5Z35T7XbAp/Kmk0ClJIyxl90
1o9P0U0HoySaTAGKfkfrUA==
`protect END_PROTECTED
