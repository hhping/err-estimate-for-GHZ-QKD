`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiuq3w+o8fijGcJOlmy8Cwxg4GgcdAN9VvEzRNNGFrx1jI0LOz04SZZ8/burVUnf
J4/13WIwirH+PxcRkmSbdymYNdp7AyREp7wU2IfNAe7h1DZBKSpEUo+EsssnqN5n
WX7offSX0ywpe95bvaBOz6KrA/vCChEf0oYC3YW+EnUMBc9fJH8QajWpYBAl+5Td
pRhW2YJRT7OUAAppu6gYHLsqhWHvdI+D1NW60ZIcs58TDRMd02QIP1Ku6J/KMoyc
H+l1g+1hEZ4TLc0YrDvNiUvUhGhjyP9YB3IXaoAOzIe/n5z9ivPLS/FzM/buvKQi
g955pz7svdqFQnR/k5ev81GeE+lBMrG9WxNAI8AbpDqAMehsaVm7bZg7qnCa/ppI
6LfLwsnD5PIygXS5vej9++HthFBrCc7Srh9O9qnOKmWnm/BrzD/MnnBjOX3QG3JC
Uhk7MihFgG7o+h+E51rrS2pqcpw0EAIQKsOIAUKN4ceYcjiNlY6RD9tStccnmrKg
MSjxtXz1NDnEFh3gPpxoMADnFy3jOEpbpESUwXG/2Sy/jMn+da5trsQeJok9rKPY
HSKGFzIlytLyHKBx5JGak9q5dauC2NiycOSWR9kLdlgqpSGHEttyO/9eK6DYbTQ7
yXHnM3EXhpv0K5QiOfGsY/qsCWB8g2zOgJeyZtELufsLLjHN1ZTILwgT9ii87+7p
oju9AhgBtWEZPwFX786YC+iOzN87z20dMC3F8q8t1bQFBIA7I0Yemopd7raBxJzp
laVsp6FV14LAYOao0h1zcAJ1v4sDiz+JnHqFQN4xjx/KQWPDQMMILXywSKoVjCjb
I5HEeeblqQqNxFVVPSw1zQj8x2ZYC6q7PFAtHng3FtVEzbK5SVS/UxrEUOoHhqxA
2xVa+Witt36mjuhwiLRRbgJUP1Meisr0bYYHQqaaFDCVwL9FIyl5cNbou4A5DJDU
+JjWp1B9YGYIvId5FFU2NuJ4UIGT9fBpCReku3N3d1SQD4HoohE6syy9wvHn+5/H
6fVvwA9bYeDOtSDLZxLTmzxbwoz8du/cLfpkAQEl6RlSNBS1doNijA6yVjn1MQuB
J8SkgKz8QqBPv/V5kfGTnp+9MNzFZRkRzT7h2ZvT7iBU8Y7XY01bAE3A/nkOUrk6
D+QED2PFdHmoqvpoyydm1El3O7tXx36qsty7h9f35AUMQ8gsiYdf81OqeT8iCbV1
0R3zs95usEmhG+Gr/c4771+T/uMC+HnFy3CONr6F5Efc4Be/e6JYuFFyrYUcW1Eh
RFTyCp6CIQbVPTCbVkxTlfKGXJoco4dBoxXIRDGFNmITbKZzjWSgi4JbJXOgdxE1
RU/jWUpXUeTRI1j1tbsi7FwPhMKDmWxM7RAhr0IRlc3MZgv8be/f0o20nbSi6ugx
Kqz+hjlNXkMhtM5jf0JX4gOZ47MGjm381/A5U5/nZ+gS2YWwHxLTGGwT6Gr2AOnq
rWTR11br8hNAN+M2xAGlEH1hVugJCAdWl6LT5/M2BflZbvA/n4vY2t05rKO+Q+Lq
Mklyfs0q6pYZCDPEhAF9mry0G9L7iawtIrDj69fjNHpLflQVw602p2qBIVq7I+tW
JaJK8DMpLWNcZOpr8+tKgdNcP3YSfy7CD6XX1JkMiJFUj6l+tiw+q0RVXhljfQgk
I0UF9lkx+sWh70iBIjqCZQlxF0cS+XG2Mv2pUZT+Xmu95SjKc55JrmzsQZ6JTKqJ
s6Gi2Sxc5vpj/70QpZ97OMVL0rn88EGIkL5pU+sAZELTvk5z8jxVSMcepYfmnEv0
3kWueZFVxUn2iZUcP2H2rodUjNy+RR2OIDhu65lvLQ9ebd54g+8C8HZvViJy8tN1
zA7sY3RGQ/FdXVaoS+CunW0kPe/aGu2WAlek+y3iJO+IqdslfJzewiIAj+IkpSdN
YAO9SW0bLXHH+i7tJE7VS3dkVJL1ajvFV9DbxSs17PYIAx1h81zEwaihJnlAW1gr
/TTrDLU8COHlvMjgdbhMF86FeMQ1SLAgxqkuyu7nTjEIEzMuOjQwMkQ35vWKN6Yj
HzTvr6I2+y988PDokZzT9zclQM1O3KIHutXy6u2WZDUsZJL9ksW+Nb/VrPAW1Enx
qntLNJvRBx5gW9MTPhMUi+NucPHUCltTRHxo0hg+3by7RZOkMHE59x0i7qcuhDnz
53TBZqjxepqZ11Kl8c9/8nAyDjQhzhKvS6DKO6bLfBLKPO1Lbqf+TwoZ54Uqttti
poNTX0QElpCvDvo0mL6baE0QQHhhblIKjJcqN+jHJDnb5iDU4zpgrhA07gssa8Zh
nu6N8gWznIAVzFftVBMpp4ekk4fjSnvsT8KC7iYc6lZDrx/bRdgHgqQx67o1QGM2
wDVewtKq7ATItOReVuO5gnNWMVgCvPUtB+IDd/wMHFQog/I7zDyfLuVA73icDPV+
R4GuzAi6IapIeeVaTpnSmm6LVLoob+lOeJxvhrSAUtK25Yy6GRXRTwXT1sIJ1hQI
8vFaQW9Xo1bmsBBBCeYjexJ7Wj4qOfWlRm38TMFOz1o8jWwWCU0uebcWVH9lbBZw
qZH92PxujX9CayVHfO5n3BiKVdePqQXcgt5iViKNqFq3dbj298JDN4lCcvjzmr20
lvQPIuIhTj+3VYUdbU+eFRgr/zClcePZxgwQAesj4A2Q/JOSbIXeVAFpz+T8DXQi
bkqjltfhWQt1FLol6USZ2kxmY+myMN+qzxQjp8fr+/rIOqgsgApGci9cR/sNT/QM
PzRrSx47eLFTvD7qZJIWeuqLPgou2+l/R1rxHMU2mNt7L8oAt8aTEzieuJgQDI9/
eW97FppUs7bp+Txl5DOaDbPYU+AxqVtUhAbkZRJiqZbW2TQVgwlAGwvbCHAOLslQ
7zBF3OGiiinxjacfF45N/eFSA+7LO6cFY2ulLYjEjqLMYBjPv6uVKehFXWlJb/8k
3OLQZh6MPvMniS3CpIgaNg5T2MDdWHl4ns3uZVR6f7v1+Y+iK1XgSmO9dt7juY1Y
DZvOdFl8mE3cKp/jzctSWws+tiyXucbdeZK+A9yIcj/PzqyNzeIqHhnU06fpE0BO
5gaHJ5VV8+pEGjP4R/xOrSijmk9yFu35gQ0yQ8WNcJrcFVxWOdaSHHzWmN+JG5ek
gmZ7EpK9e50/+4bWDIiWEBQl/R766kwsjKAxdUlwVN6syPCMk+52BIORWcj5bFqv
zT5r4qIV28n2G5M9zDIG7JD6eCcHtjPvW1AMsrsvJzC5VtPhIZC8H7k53kX8yD+/
aeAiCbMGUzX4kMLC8ZcA9aldxCQrhrey/IfMkccQdI6bh1lFpIiA24jO+thItvCa
quv1UA2dCmchXpL9kFsvncpIbFyUy14VlfLgOSaG69/IcGyIEhwH8ijacdCbFvTf
8BIaqtLAL/rjBpGLj5e9zLBCJl4XrcjVuYU0xUyggffp4w6pg0LYvsnienSez80a
V3uCWKYql9SxjQyuspAQqpPogeUTVv4hTD/xWjQvoopzowOsNnUXjqvxVngnt6RJ
4qKs3QK4af9+b3Q70fL5TjTAfRLvBHY7ft3hzVnwxEwJ5FWftVp4DgmY9TNpBOP4
sC0h1JbUWKbySXsSWUcc6+CLRixgjgrtHr59qRlepO3nrsiEqTmt1DKugPDPUUa8
uesLXuoJLHdKPuvpQ6ukVG6uw1K74C+UuL1cjAXmQu4rjfaZaD5CBM8XXLGW8zaz
Gx7pgOvbHJLClfJ4k2oSsQR7FeZV1Mb7NMiC4GYsKrNT2vh35sqAkTQDeyzfprsR
VEfaQZSq5Wy9KzIqpZVvM6WTLKq20vMw4p6R5CFYMHlB8G0T/904Sx8zSo25b+UJ
`protect END_PROTECTED
