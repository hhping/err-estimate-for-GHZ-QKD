`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omcn/Mwqth5TKCC4EUmQ/NzyCc4Y1FkMFio+HmvZVzo4/dnif1mkqZcNqANri+at
El4WdrrAc1canNGFtBz9U2YVPKVRwqBG4OlyA/neC3jE5UEn2xqsGereMIQalQh/
gostTxULZkLiEWsLxSuzQsPWAf0gmWSixqLqGJp7zDBk3lhGfXfTONCXl8gJGlpe
ZRS/KOO7Rf8GNgnSLYdLahmgc3JLRh+nOMIcFwu+UDxGhSaLNlFhYJKOXdvfIdBU
NZO2SKFMR/X2gWuP0O7unxwH3NDWugjDvKIlwEFNKnFY8UU+uZZH3NogUBtS/MHk
vkV0QT3JwKr8dS/xA/5ijlnmwVvBjEJ2eTIm2TADbv9JGqceMjvErKiEse95sEzR
1V7Er1SqGrhJr9We0nq8Zzi+o8IVi4q1NRnQr9xCQGToZWdA+Ls1HrsqAw3FC+Nl
xCUZqshyr7DDExkq1fMmyTh0PPgcdiyQbs4FVMq4bWpB/uY6dCHU5uQTQ3SKayYg
CQeH8Fgot2VvHhDEPha8MaIZ3x76NB5uorDuDPGfalxTZtFSxz9ff51ugSd2aCVi
HH/Bq5aYDv88LWyqNE2wSdiSGaYoDz3Y5EVvYw0Rvr1EUzj9OUwBxfgRp9Shnu5o
6pUx+PmTaVo6jeoHhszi+gjAwLefiC9/TSYGjlDtR3AwwTRG08Oczl2WhItAYTlZ
PRHNo03ff0S+sQukMQ9OcqLtxUIQMbU+86pd4YSdKsZQ6tiNDDl6/kIqNqLqudFx
eAfGN6ZAtaZcLVv3VUPAYrPS5CtSjBGPcosAkE35Ybc2ADI7EYjMY+lY/7kDWst6
aqBxGYPuyzm4I/97Kpc7L+6qYJGTAYpsMk5Hi+QE5//DlUUGplmjeR0GEunlrd8F
i5TdklbIzqio375rd/+CREiSXmFyVdjXcInp8clkCyGPKQ1sCNLiPqclvQx26Lld
sq5BTUkJp17GOwbTqrfCpEslHya1mHcxeWfwDqhkCrzW3tzCJi+4DxGTHGFS+MR6
4uI7a74Z6WeaVGrTbFfIKVJQ7CD249JPAL3JgPHdPmkhwyBKIVJkiL9+BBU3Goqc
LIPZi+BIAIy2rZXdHFD7uzck1c3fFTAzyv5ZIKMuJ3CQ4zkPieQDkCl5UCXs2jV5
rrIIHNFMpiUcWE0hEVUoV9Ngt9kmZSHDp70m0j7OKaGwMu3nVnbVkUM+w5Q/v6nm
E1dtkHq5dsJXZlamd1hYlvrBoQIg6lHO0Qx0/BPbcp99s+vxJ3xG7RW6ZBeosPK0
`protect END_PROTECTED
