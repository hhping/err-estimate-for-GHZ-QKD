`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YvGpmDxgnmYvyBSg2Muza+mVolF6FTxF61P6cw9XWoZyjLFWJB8e+oZuPOkD0Uhc
2Kyxe9baJpVdepoITG21xxWzQBKODL8260PS583ubWsqAs3urCTDBool7ZRVSEDy
gxMyl0yXp5DXncgBeuwBqdz2nzxrAmdBxQkqy172/9/MTSEu9HvVqNgdpV+Je1tK
3jrnJiDdFY/zhOOM90lgsUgvpgNqIPB/9+oa8+UxNyOOVJWDZOmc6i20jh7tp/fg
2P0h3yIWUwVwf/HMQzRH8yZHHx1yCDJoKL/wEKXQrjYK674MIEH2DQ6WKpXhuIn+
CU9Frjk6q31bTcLzLB6384B4kOJ1FA2tosd/X9bu+SNBqzZrVuRP8C1ZwkmdWxt+
fo+TX+e9AnjabsqW7habXgTnaeuAtJ9nzcuwesrzwe68t4nNHbjexCRjgysYfSrU
qTTNLkkcz35e6E3HlT6oJCjp0LxNukGwFw3RoL2w5v4=
`protect END_PROTECTED
