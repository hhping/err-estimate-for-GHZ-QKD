`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Up2VC68Mu6DdKm5iU22QRW7o2mFH7/5tHAgOv7X3piKv5Kt9YXLasH56s7O4YY9c
xusuuh8oPlFUGg4z/uGk8Ozp7lJRp7hvKFZP00XXSgAt32LFJWY57JOmobVum40P
aymGkq5dGqSvHEvKjEoox6yXRSL3RV6IMOw+wY+5idYaY9iy84Hkr86h6hfy55NN
IBc3WYI+8yY1jpKKlTi2NNqzVgg+b5QqrTsjwwmJ3Vtg5foWXc42rWXXOmPupZoZ
9P9aTbDRrU3xK0K6nlrfbXdcoPvGd1V1zgDzKqzsdcuxZKMbrY8riCf2TLBL8Am5
3J9GZARAf5tr52v3v9f76/L/tMKV3U2HGfIVPMrZy/rBX7oHZoSmA59TfxwQzydf
jNV+Z5OfcfS2PTJ1fqcqg1AG0Cc6RZ24MMKdaaNvD/uNu0Yq1VXOwA4d8Nk0mNTh
PbjYHjBzaJkNaaU4y5RTjhzOGG+/ZpmaQVhNZC3AXd/XxQTZeI1NtAM1NiDEBc2N
vylFFG47Uj7fjkDlN8PuHg8SQyVetAWl3e9EwfmsMKphLSiwGiTXUs8ZNCxcmYju
opzKUqLrOBAN5tLkKYBwvKxC96JCSoaGPdMIJnGJOk6719Dpa/uHa1FJD6iDKFbw
6NAmqouDKzy3jUy9WUj6ocTc/U34Xrmbb0nsKpV/OkLWNgoyYQS/35o5sXmszDKa
7IRGF+cOxpgiWG6kirkZZRzNuFvwfgbeJoxXOoPw8UN+MwyQsgasGkp2gbNY7Sd8
4V/LsfnPnoA2aAqpJrDCRB7qZcKtEy8HCoH51USHlFYCXPk+M0NL/1pghmBbI5aa
xjHMsoE7iUWK4HehFe/H7riWSvi4baMPVjunMBKVuqTV15K4ksde5Q9BSMBUIn/H
fRSxT0aLtvnrQuUGAFKWCvyDg5DD7Jw2rOL5qpFZhnY8Gh7xYBPAPRYu0aT6KW3H
57xVY3xQuHYgk2NPBT35yMWKUQIIPYGl0jF9Khe8EIJbB60ty39R3Vs/LBWHfUfq
EoZVtxBJdv9T5JLk1MC8vsvUsR78VLeESz4nFyYpVYTHo10cOx1Wpef9FO6Jx6b2
`protect END_PROTECTED
