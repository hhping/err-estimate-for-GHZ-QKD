`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOhPRq36vNUuZSwP6h65cK/Oqtj13WDtXJYZaiQpvfDRCxGBajbeGm9VBpHg9RnL
19XUMo6rHk7cXlNqU1ctD9FOIL8hJZH0u+Q4ok8s9nttQlr1eh9J9xwrgpBMxVxx
bqm3fRq+VETNVcV+b8J1ThbIL3LxVu5ZxLoy4UeWVOUblP51BPiLxUyL7dnhuBg5
9ycsc6pPhANLZYbTOrWhqw5hYZqiZvzdZJosVZw/2veQet786+q780Digj3E5I7r
lLLi+StiqDwAVENGHD2TmOBV6/sL9iMit1v53mHp7JkrV2hJd3vqKlA639QMEggn
GW21LCiPBZuX+p154yFHYbMaOXrbYhBjWyb7A7hnoelH3ZAi+CVhL25+bxpiBfYJ
Q+CeB9VkIJZ4sGxukavTiJKuIIi0UD2Hj0cMniHqiIN4JqwWrYUxWFM2TFrDxgs5
qj/zrSXOyE8uOsuKVHKyRRFCPRJBzU7kEqYjRxutDc2LKlYgThB0RjNI1AIVgQaB
H8TeRspDcgLPqWl2g0svp9JIZLvnWIhgeHS+lKZFxi4YAUgm+zR4nSE3WRmy7So1
+iz9FTO3TC4lZ+RcwdTvCxS0kyOP2xGCxQEdIJXRZzu2O/eVgY+Di0JUWsPh25M+
9lDjmwb3nPlaTQtph4LJKDEPd1pOKKI2i+OLirHy/x1ridCLF3PzsvVIHILp8wLw
V1ykgfqQFc6Dz5oY0CXJTgu13BVhzSMUTZTQPI2cbLhGIVRk9eiNgTsoCCHCfgHe
x8tngzD1TNBWYvADFqfEXm+5bGG50RiARgLZW7NEOxjRQ5visvIz/p74xrMIL65l
`protect END_PROTECTED
