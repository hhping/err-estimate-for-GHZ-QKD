`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BQlU/1BlRR17Paywc9x6ucfeDxtZKelr2xmTdXZKXxZMbLRORh95eDNfWDG/Hly
kKfhzW0i1g3AiTD3gIQ6QKu4dAoONTjqbKp+Gz3R9265m0RO2Ni8VoAiTj/2E6El
WqUjAh3N6LpHJ4VlWn3f927yuOopz84iNOrXD9MmC1owb/d1qevwCSosKnMWo+w4
d5Rj7Xp7bjWa3G595Y4uPbYGqNJwYEjSqgIFOXnLeXbINpILPOSC0qavQX6dqUKx
gJcSFA0+C0Xr2XJmaUXys1CpaefZGMNhLaUCJbn1JRxxftrEgo9t17MUQ9u/Q/5E
/D+WCTgPtvvVZtn1MF+9hwQT6mkKgtn64HZ7PuGH9UHuOiggutpAfpB3GUXaQCZm
MNn2eNxkglLrHKWiOBUVuDG5WHMgmX7W8T7Ww860U+OeWh9NM+tuf+BVzvwtDQNl
75xr4yGAPF8u4FmLAwwkykEEpyrAl0H6fnnu0yq5IiFenkTP5MQj8/QgvBbM/dwi
R+ywlQ/icg990BJNi53YbrSyAW2mzxS7iLiDXIROXz5oXmVDFVdRLXG19XBdTzza
Q0kMMP/y+ske2F+pHi5AcNcZ7jCuEpjfestQsuzBzzNFme7mdOPTkGUQ1JTOydqP
7dvaCPj4HISOkIAw1RoaHzJ0fe7piamw6uOFv8xlyTOk7yHbpChaa0duhi06PK/s
58glbGPdgAaeAZ2EepVi4PAU+SMsKY9HYxZHLWek88+vghF9/HSWwPa0LPe9GeSZ
8nh/N5gwV7VqjUIwBj5Wfy/TyPnXc79tBmWFYKBPJQjsDG4rIfzIkXYA4eR3Kcn8
vc7Z+qZYjrN6NXpfRWP/aDjzVA5Mu47njorCEfzmAn4hCyJhTdWhAIRg/7oCPeoK
sEidBf3brCrDKv7DJLXoCl+3Whqz+pbhEAp2TDcNk1IWIcYzpxt5u4D0QEjn5fkH
fOCiGQ1IvtUJUYKrkv8Morq3Z2fU9Lx/9SGlV/WzqtejDnQNy4SfYZ8DDc8uZHtX
9VoJpqAi6PtEkHQHfHuBwT2CHy/fcnwOuSY7nvzVHUbpC4o4Rgs4IPZ22poUxGw+
n16aIEf3r2489xVKwVoG0Egl9COxV1P58x7/aiO7bhPsMadEYHNxlTplpxYspR9d
7DXgEXC3AHu5LMZjkvyYkiPs+QX+oUbpgXRPprlD43Vnt97WJlHc9QTLv0Yf0qqE
77KI5Z/DSSzeEj95sYJvct6MgJbLjiFP/ncdsj3boAyGIVOQnPtwukucKQRU395Z
6Okpy8MwJXCypbu3tHlDf2IpP9D7640EsxgRJi2Ax+IJanC1JLYsdckPWRL2SXPh
AZgV/+yq0ag8kW9Pw0nE8uPwqgCMo5hcKy4jdixUBPWMDQ0/v5rtBVi3I4lOoUFO
ixkrYmr6s7ZCB9ihEo+yZP18T6YXn2rBXB5j+nkbIoccp8fsxzXjpuugQyj5jx7Z
igCIYTldvaXNn2Gs0pOZfBlHKGUo5RVcVt96xYrjAMSMrU2aGe1SEzn9Qx4Cj/GD
+XMgtD2jLZVAMpdp2gI0Dsp+/C4+PF8/2Ij85ww1XorL0DyMOG30YYQ5M0nSGdpQ
xJseHDJqjwDX2ZHONboglB5oi8S+rYzlXfiF57ji0cEleJH9aZENIcfzekz7sex1
B93jHOZsIkQmrHhn05SL9A3zGXOUR38z3NvLG4fSKMEaiO18eLJT8HlZeE02PLe6
3Ff3SSVMEYQ89rco6S+y90aLBcxfrmKk2Y4Hvx5Isg7SG/QZkaRYp8BqOYkG+Lms
kzbNmJ34Ii6+V4C0NTb25KWjnyn1kYt/fBKffAGo4gZVKsG4EkzX9/bwIrDGTAsx
XRdIU3M60diF8gjgH0MgObla+W0GnTkWcUvGn//8cdoreApYudzuvIgGmabFWLNu
sKPBSegS/oYBLAmT3/aPs81sXdBoW6eRJeQeG6zI/73bVxiU40uwQamkpGVWjtgZ
d+7XPfmGwdz8Xsoi/788aDqkj7jkVol99W/sws1v+2h5nb8YcMQlAsTxQsKunu01
wjpLrMz5JOPL9FlyafEkaLX4dkJyZWGxp+ZIBXv6dfIIGbDAhubr8IWzkVhrIaC6
OG8qxpMCjIAW8Rhc/SRWP22gx2WamTepKIVlRlTcQsAw8/oSBK7ZnasJGFicf75t
i80VHlLv16MJQXQLLmVMqLZxmVTPKsw32kmclWepactrG/J2G9e0Kgr86vgarUGv
BWYNP7hUojOZdhLNlhjV8beEShqH26aXrzh4pHizsQ9EgwL5/8iq9OwWy5rHQkKu
dBbqeUZr8h8B/MGEVPjjLN1/5iTHEFNAzQqEQIJVoP9DkhJOZnkz88SEdW2FkRJ2
RNSHrZVhQEe7RxwOamg3q4bhK2tq27c+w7ApeFw5P81DZvg60yxTQBOPQD9J+oYF
mYiWdtDeJ6whAdcZhy2CxaMudIV1sfHLzhw/gmEVH/gTrYovlyrauwGEhg/iQYDu
ZhVqw9Y3xrl9MLEue6pigNHdlFGxLV4Z+mE6GqHRTDzquRF9/IaJtgXZm+BJHDwp
0XVREF0UPr9lDa6/bQTyJ52/uwDc7JvBDqNIBXKdFwafGShOuPq0hQzpee4+lrgK
aFLibzHlu/ZdvwAoNGI6R5o7dmmDeFG4dSFih3kzbzysqRVJzmPgjA0VOu8b/K2X
C8ElczBwHmKG9xeOwRSNZSve+zNXSUzTnPDuzHqp3f25FNDSRlcuNLF2WL6V+4PF
yvX+j+GIQsbQjZsyW2LTmAT6Js0hf8CfMvhXFLHYUFQpIVSRoLoWJCyoWeptvER0
uYP5p41rJCY952MxfQ6BWqjHuMMcpe7h/WiRgL1C92PicJ52rcbtARi2BZzXM4++
0D2UjY3bXh5H8kQIuI5wBGn37TeWzY8ZWGZRxIWz6XMOhkcsD7/li8Lo0Ad3/Lfm
UR4/LFmzZO68AT3g7QdAIPTNiV7DXgTgGDaLliz7ugmbnVpHm1McqiELBv/PAWm0
I4yn1FaGMPjJbxH99GRW4Sgi52JNOY5gWg+nhTV4VJ1d6MGt425Y1hoWkbHNztGX
6TS1VOidC2Ra2bqd8WCeYg5bdL1Owh+Ctsx8Y66m8wvwTVMUWFf0cacTttg8ZZWd
AFge8a+cd0ucM2+txf6x9eYFEoTFKYaewkLZUCHj78JUPEdwBTaheM1PdDN5FS1S
7xaThi+pjuphtsmL+xqL3l+rrDYhT1Ee1xCeo3cF1qj9xw2wrCkkvF14t5rOh6qC
R1FzaKnwmmCWJuuDrb8Sms/vnHZmFiWJZnX1IgVXRqTq6J7cHGHwBoMfJ8x8lvrz
XHFrfkJM3lN+zHFZlyMM7mjB3n09RtMcESEmZ2h+il7Cdi7NIJU5TioGDspr7JVX
O5LWO+tP1Mj/MfTge9p/WQWToCgXJ1WwP0Zh3XYjkE+g3ZF+50mLm1VJQAWnP3ZW
LWHoif+LGXrwZTZi/IomxVDZQqXBCaa0FaDW5H1K/OB2Hcog05uIl3BlvUbPsCoV
R8W3oFwM1iRIOc/V45/GBuh2BW8tLr2X/UvcIMd9RVxBZfxQQ3oN3R6C++ItnEk2
fQIt+kRr2SDggTm6+2XD3XgrU/psyicre2rRRHJnOE59KtH4i0F4ouxrYcnk96Lm
jxLeghGZCK9A7dyEY2mhZ9Oxs0fhSOSlK6K8ylE/JcHAhv9aaC/eIhvmUJC4dkcI
HCsK3BLZcUcFF7nZmGnt4rtrS8mCl4JXv/4sj8NZLSKdH0R5sb8lLyA4XCfl6UXv
mcj5jX4zCFXiYorytlHia1F+5cDMczpb1ggcGBGbj3zRotu9fq5z3MRTHQzRZumO
OJuB7cWB+AHL2bZ25vrTqEaWOtusWFWUE/bC6zzPDCVUngx+ItzHm6Winj+vTt1F
6/ynerjdecWEIr2eILNiuvFXxCorbTijiIUgFSfmSQ/TYDvKy3RwkU6FjiY6uXVA
rI+sPrKfZ8QioZ1jx5//K2ZAIeyzDwgPA3uF+si90eu5F1p5uyFk9oZ0jwcSQdkN
lP2kU5JCyWLXHR6hGKXRxl3Ug4ELrKX2y7Zf5IhvgRdB+aZtJUVnc8sdPALsGo31
DotStErBYwxwD2mepaAyRXha07a4yG6hI4hYntZetgnPMHyMDsdGMd/tipA+77c2
ZhE5ALppmRHeI8ctgpN/ADwwQCXRUGhOcZm+2ADgAavq8nj3jihosgRRfj3zWzG5
9N/4D6ijlFfegxGqf3Mr5SMKHgmVQO0qF3t61vPPpv+BhDtJHdztzIjRhqE1t1bn
MMywRT9UAnESPPJIXfoF6uuhPV8Uuh0V4TPTCI2jbzzMpyvO7TXaprRK7WgIjqKl
x4u0nMqCcnQpr25Senuiug8/YjtMwQ2+GtFyJ5lRy4Exgy1OkruT1qsux3rZ13H/
dlUB+WuJu8abaP9emcHlFkawjiB0e9GEWM1NauLqpcyEuCbP8Utb7pT8DkcKXYmg
pzvQMvuczikOoyEy10vQDzknmltV6uKK2ebzPCIzjtoDP4zSH0ukHJR8qvNBQtvH
HYro8fRVeweGFnBbPy+7vs8aJkpr6s0WRKpRfZW2seK4iiDXe658Nm7miPWUD5Bt
zrbjhS3fSpeYi3FKuSSbcrAw4gEc9G6tF4wQXOke8uNo8/6fokQlYuEI72XOYU34
RnOP2MiE77tBRypTLJbU3g355Pkar+mrwKI5w5jjteRr5IIuHuw6mnP/jBITf8xL
cfZqq960omiiqhk/UHszOxvWEalq/pv/7pio0CQ0GF4siQvWbomxOAAIwXLAZfMM
oDFKBJuk4HDaYRrgK9LdNXa9iIaLJr8jWNaAZ6ZC3An49YR/Jan1A3GHAKeUCFwb
c+At/F89IYozhKoNyjucmXhzEx6FmUdn9JdbJvVF5BFcc1UAQPL0DvTswqtRrefH
wH51bWmmWd0zBAs+2Tqx4nPDV/cBhlSBBiYKfD/IdzbW73+E8cK3vlZt3sfHlH41
K/Q4ww8ho8SCITJqtvtmNsXfYJVwWrxUAu2bYfmdT+IPFY5v1kZ0weThc9bLEKOL
0AsXWGZNUeF32khlw/33HBF4+8rlW5qm8vDP5Y02I/zv6ozqhcmYzL8ksbpmkLoN
0pm/hjKk4sYj3r+SfGR/zxEupzhIYhgVSYLq2g60lwkvFnqQK5aecQxZfBAAAeOL
sCBO6ipUlcCTlEb0KkOMkEMnrkFQY/PSKzNrO02yx1BPDQIuZqQiSd9Fd4EmPs0j
y11Bvu15qwv44gtD5w+RNKLs7fdg4QcruL5GVXCL3+pfFXKVlg3Havlqot4HOsmJ
i7+Yaiz9Ed4tUHJq+tOPe9RV3FbgOpGX1jsl5gzxmqx3jGBa9NYBd87BKr04ORbb
+i717udlPKLVa/OSJZWGfkt1a6HVCjc7XjfMGa7iS+745Z4ivkcSf366eDjmGSR0
+BByAL9LZbd2E2STWkRh2yjmoL1npSW1oi9JsN2wuNFQvo3Sg2Kr4DcdoCcmvMIp
FmwSRKKrsWI4US6ZHQEnijQnJo0E5shWj+0ZTu82JsNDOCEEhNNNGxOfBOHS7BSH
Qfv6hhZovk9EEt2jh5GugZKxvyQQaZEESju1Xid6nZV2xDHReO7TXkeHE+pVz8hC
pr56jC1uJ3o4/JHOGSV4hVGbOa2S61ckIEN9xMiqhbxL2zy+lIGcM69b6b1Gy5uJ
e7gc6b4pBVbNA93G3CVMSb1WfavumoYg/nJ+eBrM71y8jgwrPgAC712Aa/Bk82K+
dAmJx3g1L5u0yF8YXmR2Q/+B9I1K8vIws9YbVhZYLeTy60ViDOOHE19F9COO4Rwu
I1gxGgDaVV8SlFBrHXvB7pH8WNxnByw1PKCvFH+EzZ2Ki6Vf9biy23dqFHXXlowS
TEnIHSubwZiOKDPZZnjnxvaP1UrZMPn3bTKRsbjmv6W5IJh8VbLeIBRIjrcQM/IG
O2EiXtcgeK7d82XcQGganK+BdZYrAEDDe5ruRIOlCLDtfQK5yJU6/uJTTNIeWngg
u35iW5j+wsVHZcPQyVhKasWQK6dFRK2fqJiGJgTNgEzz5oaweeLo1XELBKX3RB8X
Ueinwc028IgrwdOSHy+GtAxEQrMfr1NYHewRSHfR8tg+ox4sQz69N8Z2aQA/7S5V
97aTaX2UHkDH3P6T77weOCFQo6lakvqd4sG0o22lDWupTpQNxowmH6K749aZSKoq
uaki2H2yWAdY/WEjI20+4lerek4gLmCTBpcsJ54NMOQ3B1tSOfIkvzM/+Wvk00Y0
nQDHuep3c0s3hjmc1FS4gLpiHILm6r0r8xcrBCoIHxvYAYWw4HOoh3n3xgsbtPJ8
4g2Ln5/+Xoc3sd5BQxzupgG6msTurmIeLcaUULR5Gfc2pg3DLEIzEwOrDrWoJi19
Z1cexL++o7qaVGTTfLL6qX6u6dVZG8gL3kn5sX7d8A12HxR+7SaJfEpR/hS77tbz
+Mk1oSOROE8BoULR1d1o6k552EVBDKbLWwU6up63cpLpyiQKuUVW6gusPT7A8Ri7
geT9DfvYnrAR95ILMKDjkK3b3IJ8aeKVjl8svBPk5V0njsAS+sYyIYPsEzKimHP5
V9kHxiM79nJrhJlda24c1kG+UDD7gxNlIU4z764mAN0ZQbPHTFJd83YhTkR4WLPt
IAiC7DoJp5u9VicY945IjgTm97fqMnZ7RLnxSYNhKQRo3yYAYacB4BlVHVQ1Z89x
R7LCmfaTOlnXRt7uARW0VKeuXFWwoBLQ6mDKLKaLTlG1V1JBEcQS4cM/+ACGvlXu
pS4rUlbpUP9DbP2cwq+s0NNBfyx5e+eztRhlKMgI9dY9A9wSN+MglFo0CZsA+L4U
iGoAVYpH6c7MYdva9Rd/4+oU0lM82pKXd2WnzQlfd8id7JcDT+2H+tu+q8lvwk/Y
gmv7rHyBqqyIKMlD5HIn14HT7YvkRxLYGSh9n0yCu94vhFMXcMSSSIVdE8n7a+gb
wIURickRKT9RSIk10b3yrio+NlNQcqHeG7xPwQPlWwYjlnLC0lJGnxJCHqTFerB2
/n7GpiLivYW9sgNSqv3KWNZARf+ZpkbU7aCxCyhZCEEhz7iAxh0HV0kn603V9cf8
blVDYP+Pjn37cFoB6j0R9gby2PuuDCcnbQr4gfk5O/9rUti1yOZQSYGkO9LGGHi4
Or85MxhXGLLUJ6cIjCs2xuCCrY7t62bHdmUxDdwbclbUMfI+HRKjFDco3Lx84v21
0b42/rS7Vd8s2epWgKoF9Oc7O/C0pT7q58fixGv60yRCi6KnqxdAZ2Tu8dZjYSq6
K3S3L2UgzxBEPd0qwp8WMccg5RQaQDHAkt+FTOAYi+/eJmjv71jdTmtrfYsW/GUS
jnDDGJtCHe8K1AYK+R2nIzugrcNf7XN1QcrGbrMEaKFJizXK1g5bQPREKEdOe84W
GjJF7RMN1OZqlRCGOxJHyJaH1ZoJBb9zUJVHM9Dp38POjWj6/ME1s5g2So+B4NwH
hil5OmFFtO2LidbRdDjiQgRr+sWz3Z81c4yxFRihaDVODhWC9P3qT0fte2XQmwnp
JCjlgzFKyvIXgy2+4SHJawBgIsBr+PEUtivD8t5dXyZt+e08JfOZz8NOyCcga6Ez
LbyDgFErA0uESdj8Gg9j9teL2/sw4Y4DBz3lhE1Il6dA/cLiyck8H2zPPu7xjEyU
AE32BFwTxdg8d3ZXNuTM7lz+tMXPUNDFT/XQAaKW3BkukLXp1wrdO66aDEztDd6M
ohuqJrVv6BEuAdRNQz5JF2OoPdVyiUoqLyYMKDwuVlDXJKdYC6M3xcN8VKHVKt4l
KeLAr/9AxngrqNGahsYQSFGyZVKmUninDYq0MIkR7xSkAngYjTU6zU63w2aBUC62
Xy5f24WJvvJnfXKnW/T5KyzvegFp1uH1VAzyvbAOnwjnJ4zPfDp76uMhaYFy9RWp
hWL/GJd/nYzsoJlVtPUYP4qIn6CX0oxIOyf/2GdscYMuou8jE5FuVA7NQiPen/sS
lWWMUliJcITvb6pNrYw9eNXuKuATqhmsA8qwwaOJEAErzF3dnC3i8QXCaMti9BzA
UsmLekhXipCgu5Lsi3V0jlRcfyHGsoZevUKoeug7uFhIQVFo0zjta15KrGW8MN1e
DcJaUnHn+fSSQZoWmRgY1FH8g0/S1L9eebete5xLrXPT5epWtwaczjm/CaPBmKC2
4rHcMHqTyVBO+NvI2xCcJNgMVy992ArSBn9bPlql4eIrofhnXDqgEoLb13hRnWo9
58YFyA6Aoy1Z6LqZZpqjIbrFv0qdVXNM46QHjTlvJb0zaloAhOn5lrFOWhy8XX+i
G84iKhp3FiYlQLzbaMAdh21BM8hWhJ50sv2XPYm2BplbXjS+LgDwY56pOKUFwXeE
wdR9J0uf6XJ2fCQq3REjPNqZuXVL0JpDPw8vqAqRU4IpfCrJ4fweqf1leyKaNQ2M
OS/9D3f1IK9moJY5J/gIBDb05PG0J33j1JVxC+2sLISHsqvj0YNsF+cxqw9RQhDY
T38fsrnxEhcffMdrrRtepISnetfzRhcsVYQd+hDz9zB+IQfQePK3Da4DkVApuK+A
a4zDSDd8E3SDJSpM/H6SHr71DeLcJZSpqXLMySoA2pwmg/s4O/lj26fjI2K+WKiq
oHUHOFpjskFB8JlNudrzP78+qgvvztD/ThWiAQulLO2yddBRmnlwenwv5MA9RQ4A
9Pw4LmLk3ljLCn/64s11rRIMbj1DMCLAP+RKbkiNmj/5r0YXZyMS+MpTby/xae1U
ieAz1dbGPN+PHfae/QJ3KEoNTtyhgvaC2QqrqJdhobkrnbmmxkUTYbmMrL2ue9lP
LsQVgL8qDYlnIQxr8bwvpdsJlpLSlvTJdrxIbjKBhcwWKk32IKpHWF3FeZfdRZQe
3xHxuf606XzjpDbRatmZQnCIUZjOQX/KSuek5RBe9oHoCu8RxZjDgApdcAfyt5aS
itxAdmM+zlAMLL3ksQdLTwxEBoakGRfxvnsqIyIwpkHiC5Fwdqu/yKKwrjIiR2Pe
XoyvvFvgItAHy5f4z2Fy8Z5gcVwIaSucBD3cREeWh7B22zx7sHIqM/R0Gg+3xFc6
WaTum2h5D7LYIuCSmd7/yQb5aROt8jQVAs/U63B0Dq4s3iWT6K2L7ggsmPSteLGQ
4nPqQtq5LsdvEJW0vgbwcQ0aHaMXqk/SG08bSTJ1ykZetsohJHVW0VZUY5dTJ7HR
FLNrh+4R4i85fUvKQnpgFRhD0mONqqwMxmSZ8mo9TOHd/X5aX2+JGD/e+QBBAh9B
AGxTv2x4pEmFwCfdLFYCGwtexP8o/GjaRErCYMbjq7h0S55rocy6oZBbLmtrepX+
UCZqp7FPOidWnSjlyMRkCn5C/la3Vu6Yqen5jbAUBIYExwpvugvB0jsKG4xOhKiz
810LfFkn3Z6S9wDCi7LrpyDcrDnB/eyw9ddZp7apdh0UYB8j3YKruOl0xC6Vw7s6
tCugi5U2LK23dZHpbTiBf6F+pUXFi+RCczUniVoznhlha+6aRrhfRofpzR0iWpnn
yRjOlvdLSPcJ2vAqAapVUpchaoIh4okOY3fh0IMsH7FU9az3HjogyuO3DLhM9eo/
A3S/ns9q0zcuhCDzkEGulx9JkaIV/K60mAo9PcDida1PE97LTsITwNHxPgPQyMCw
EVY2q7TLitn22RIJvkqjKMs9/jlL80W/QIlsDIfCSLcbMxpDB1oWFLSU/PWk2JOC
NVhH+2hPfgQF6vhHVsas1g5g4+4LfEipkLRPg2THkuXxyh2kiMuoBwJcapcEk5rg
6K+twdeu4oW8qLQe71ImWHLJltOkf5vG18gjtf0HCUuzr2DI+bOFPCcPs62d5o7D
/1N1XHb5d8B7g59qx6rkEn7BXDOYCVPAAVxGeVDwAE2FdCeU5OilZSg6QvOiYFjR
gduBM7eEdc+sGQWPDVVKsr32Ap4sCMQXPqV3Ed+4SAuQjL7Orb8U9CkooYmmFBEi
nBfW+wl4Q+MVKjvcvDLVDHA0dJwM1EYnvJQGDHe4NQvSfj59Vo7P4Jh2yoh9IBW9
lu4ViLAwhsWFC8cdtHNRzyjHXvH+UiwyjgRUV12FclRIL2WfuySHXFrfuJVaGz4Y
sSwblgJqNg9VgV/8Phpca6Ri+QKhlcFFE+mNE+rV2pIZI6Kozx7Vf4rmmfF+XBfe
ktIly651r2xziaDoybDA4INO3GaZEvXiovA1oCMut2FjZ5Zw9vgJCnCAJ8nKMjCh
UexN24mSLsw5kXznsxHUA4wFUeoKJhpCl+Yl6ztktaGnUr+v18tr8P+5sql4DSFV
T/qoXob+Y972w2HuKCSo/jQvTa29sHOOBYz7vPHBsZ4keOLHn6jl6sN4mbxvGf65
ppF+9oDGEmnaytkKxKNVqcN0subOBU6+IFPgxzfrq+8rdaQDChXVu5+QujHWoq+7
QPlVp6dcT9Zska1tOzjCn+7MUPrAPWBbLBqWeUw/7cV4LOnAhJ+95GSU4mEOYxiB
2J/5xNBsBUvFFQyaIahtb81LZWRR0BzIBxtT1MoKlJnaC4Iz120gq2fslQLa86dT
hVkekfQW8vCmUmdo5pcHRa+C9cM3Jp0e31FQln6uEB1kvmb52iv+mZx2eUNFH2yS
M3QUGHDR10bCExkdZPjnazKDX1onD3fbPrG4tBO6h7Un/HSfCTZH1xVSTRdZjDzi
YLPX0tSvrxT0t4pAlV8XflJib6gPtTnuWsiOXX/pTXXaUfdam214TOWPCMoqxmsJ
aMLum8ROLIDCaR8nKbf1EbT9pZau9sPLRqi0pZ5AblDdb9Oeke9JEdKs22qfJ2a8
04RnJedulw1HMQMmMTILz4P5kV48ySs7ZkUYwhV2b4GdY4GPDf0vU+yUpvWOnRKz
fWLIsTpwilu1Rd/OLKJI+7IOob2nTbD6UWFsB6oxLm4R7Y2oSgVexaFNQEX6sbDr
lmIzUzJdPGJ+Og0U3mjuMUk3FTmAPU8Tv5n76uFzQxJkEhnoFNvBEit1jDAs3lUw
3cEDfyoGXJcIZD8gBGlRTJfZrowJZx9qClt2wh8c7qtMwNTaqf/1Nzq5poK1i4Pb
+eLtC83MtFEqiiqpX5D+Bf39Ypu7OBLXVrCPDzSfofdvtupesPHkiGOMpWS8PZ+k
OIrDrgplA/15NM8x760OawXdOm3t9EijABtcBZVW6dm96QwzFDjT0QZ7CH8VdfnP
BfKepGhMLvQciGY7Jzo9RXiDD0NIvwKSGa3ATpCf3HdKnEa6jIxqcPRsCcxkkGQz
+Jh4KZ1nzkc3FfN3biJ0tRaXlgFxeRDx32lNRTvH+uBgT3dr3x37ri4kffkAzLu6
6eAmTrnQe1dt9wh7tJ0zasl6zqYLe6dhJUxen1zugrRuGzsGgsx65wBma2xDSZsH
TcpKKD05TvtLtHNl29H4Q2SU+lRxuTFn7Axpp48zv/hL3g2SaTHudfyNV2sWjLdn
7647qAAugqwAYx8QrvA3PV94JO6L5HULTybXprM3OjTBdY+dXsZmfjVZ1W9qjOrj
`protect END_PROTECTED
