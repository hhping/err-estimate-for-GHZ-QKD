`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5g8C8ps6ZG6cMU4ClVJ17PV+sy5MeVj8kFVHqhS3qVsczcpwLDVcAix2YtM5jBs
N8u1AOA7tpQuEc8jrDwJzhlD41k+LJp2rK+IDWRpo5PPhw45zVr8xNNmf+ks6Bft
gKb+VeDeIZAXUOF7+q7PUmhSctIdgxJocx4XcWbZJIFQMVRgX2qYO8iI5l78Xivm
wI47AYxvXGtpfQT+Swyia/v0VrACjHO7coXLzN/96kxUqJpXytgHWmZNi/I5FVgY
ITpBaqVU1ZRIw46UWX0pDdIkYHMddN6BPF6HDTYcwJFlKP0DoseKjty7aVg4dH6o
khkwu1d8YDy6S9RLuYSLB/mw08KM8YjMjmZCRYqwDy9Ow0xe65kaXGyPgLo/9LdV
Hq8IIMhl6swLdPfh6BU9Ukp2HhYJPfv0sdZ1seRMkMEfz8QajdgQGZUOfCgP1JAj
ZNCQKsIamZG693bULAcw7xvrDSoItabZ3d78+/ckQX6FYQDpYUiE6UY9XWFpptpZ
7qwbNtUkehsjjL6HthUTv5/ONu/0u7d9/E1bEAyh5w08ndOJrMcYbeXrfoL/2cOD
oezDBsDl2UIqhibGZZtB0NJYb9vwgqBUunHI+yLfXLuue+vFoGbb9O44CObBAUl0
c/RQbZgarTsx/5LI2kV6pusnp4Hwt+QvjJP776FOueXA6CkjXC48tvd98bgX2JdX
FrTATxZtmFFItB+iXKSDsMGeos6UnOqHy/xD+t7lfU5vCxbUI93HDxASIhUAcnBq
HSY/VXfer2XAku7KCtSkiAHqve9vKAJRjNM1DHgxavNNrbqDvN9aeowB+E1Xjum2
flD6MFwLGKsYS+LaOfe56sAuzqzXOqRea3m0plbJkKHE8bcHrLRzIkSQf44KUtR2
SEi8W5adP7iM8bclT8Uq2vopqe5UZzUBz+h6RKqEEIfkc6+ZX2RKSut1caU+qQ3k
2Vr4XtTDf+6W1x8Kts0fOIjsoOvlurbhYhJcHnQThbVE9Uk+qfIgc10t49gGl+RL
V6M1tPFd1xCWLNijgB81Dbif74+EAjyEoyr+yeLSRltBiNJtiN9rHdzBxxkOCG1v
6/JmBk+Eyffl+tmRxYO/xcmrKT3Ur5jkiLvW2I9B7TNwLNQacdBVNKUDlI0NzmVZ
nfhjQtI0pxmomXE1OLNAZw/dsq4+SRhY3YVK9U1InvGGkQFi2wq+kIC8VvVRfXeA
gpGEHGvCcSoE3TPiU7CL8nKRZwMy6YdnWw7LLPwzCqI6ujbfSbzkMw8Cr7wcMMk5
s4IrdHVvWLJXwRMvGPFq7tyo8xu4EMf/oqQl68iIwSOxAFYWmpvyinQ2UPCnLfQ/
mN6d/j2gU8oMEz50b+op4KUVGyaf2ov2I1U8eNI34Cln6JsWgKmfxl9H4KhxsVFM
BnxEiTC79oWBr0jux/9oIIC+TAd9wB4Fc1ryFCrwE5LLsLaZieCzfGLB92SxEZc+
/7h/aRLids6fwVX8sOKqc5rZEGYeoqCKhYc5HE5Vhf8UPu23a/P7AbXTeZg3TGh3
zlYcA8lkyMldi1b9j4+RSChr6XPjtHrNwT7e1nAMeqpmwVmr31tdvNTEZ1ZPq+Yt
Xq9NgizSjZfKXs5DtXghownjt9EZR6hZVAWMam1rUQkqJzfcJAFj+bYslpJDmTbY
tM7mWa9iTSy39eGi+qViYHnh0KxY6RJA+T5dQT5A/WpCZHMn/vfJcmIFeqn9lljw
jaWPvYUGeOsywJ/WILf3wDXCMahU83Je/9zUCH/IbbKnmvccDd9zpfZcmEiUiGcg
oLoPcA+uBNnX/X4K9ViGmCY8mU0axnZpitpu9tI7YczG9sVBBBbM7gJ7ua5zThT4
G1xpFiyCiXp133w5Sf+lFTjZMyfK3zOTzP8QkrBaKB1E6baLFlemOvShdCbTBbyS
8EPcTGmSpSJD5FNfex7RWXTL/73+fKa/e3nM1s7hdkjf3NEFRkSO/a75KmKUK+Fa
T2ciTU3fljp0/w51wzwGxaALYJO2mLUgCPfhWRyFMr0INmNlDKsn/jbjAPT9hA5U
wIGakGQA+CQpDCFYu3bJ/GSy0AoyXv09efXR4xjzrfPWiUq8a/Ep/1sxdUIzKZf8
XIDWAciZcfFjUN/79oLXLDo11Ui18UXn2X1WIXLP/jRctnzxfP7KURuJv+9t16Ni
F5J+yo2lnolqENEp0yMZTEzw5jeavAx4ZHpWjZk/R3v00nvsJU4Qg86iUyZ/0mIL
Y6fDrV+qq4X2YxE04Cp3EnCYF3yCz5LhcV/U5IQ0G7dzARYb/pAu1rGOju8SaQk3
cF0xUbrQWVyTidm4ksq9ITiee4nEkOMSWQzio0r9ZnnkmzSebDQjeKPRc1oTy7dp
t1+oJ0wAKwBJ6LyS5oY/5TFRH44BpxCRVLksyRShIxsOXmR6wxBeEJDN2c88Im9k
5/0q7YR8dA0mj/t3N/G4791/l1pbEtj4C2NxXy9s5gJMHqU3+TDvmdy8b1xvzcxt
J9+LkiUzY4MDJ0uWJvxjdKUCZ4HfptjWxS1pTF4xVfi+NuxuNtwtpeiwvSXrxkdp
nBlr5NrBBmStB9awTOdZ0xl6Fh99X9/dcLlYtceRp6MlhgbuvjNOb+b8dWaHzQjK
28JE+Nb4gJNmM6+gf2YPkmc7TDRCnSgg59pL/4qa36ctGzNqLPioDLY9QsUAiyXv
x+gsAw7vrIH3oYEEU/4s2/vN+o3bDIIyZPQXDFv2ML9D+E5BoxqvOoW0bDeeoQ9M
Jux+FWBp+3mSetYYmVt31ZgHxRkGApKJbufEInrR5xLs4pHk/Wi9mDsoooH9eUVo
j4iGAXysyhBFV6sVwVCabak/eGSP1F7huMLqsCeAOfhyz6sHe/taRIIonre6SFz2
IM2fvZe19VWYZmnjYnv33Hnep6H7krJ0Bjke9SQSTgDYkiaoqjdwdeXeWFbvrOnz
XbTv35M/GEdZ2q+2kmjbDRQwhiJcTE+QJ7CrFHzmETgZwIJDgVsO+aCM2iXE5LBD
WFRUCscG9ezoPAGifAV26HB0ZCl1M1sEMdBIM/1pF7M/7x5KYoWW+6Qhk1rWC7Gc
sOBHrBa+NYBb/hmKMNoN4WUNndQTZIYqjZfItGHq/QuQMoW8FO+nudX2n4UkAGGr
bSp//ADha2zNhIMfMG+JyfRhU3xBnGRmASOmmQxedPPHMgLMPQztEM1fUY0sGBzt
xSQ4QQ6/Tovxqw15AEvIj+qpRTkrdQYLAJUI89wzEN61C2yQ1o+KBbv0bk5kkGQ+
lBDhZPxyUhoLJsVL3O/4+1dUzJKRGVXiIs3hj8HQC/op6nBc/6A68TMQnSlx2l02
DLsEGkS3pFcYH3okjkjEyG5u35UmDOy84ikXGD77DlSyTIF0Yo8yes/5jFZSKrei
XayH4PHDu4dXwG44fkraoZlRYXJyJQlmdM6dIL+iM4+e6bCfEnCz7Jwf41fFblVs
7OV2wI0XThaYGTf5SxWCXqQ0kJDX0NBRnMWJv/6bIrC/L8afi6LmNyWtuy6lfaC7
8U/NwvQklTBR2ukR155VzJeY7wf137z48iXCopGiX1ke5NyfzvgohfGfxIlnYZJc
xjts0j1OqHelozTIlcz8de3XutEro0sNHMTsnVHhobRk0ANKu4D7ahv8heMD3dUs
dUO3g+zuI2v4ASknyuQ1hiLcfmWQMXxaltv/GU8wbq+YuDR1P/EFb2s5NRo8Lqhw
SrySEKiU2H1M0+auHZIe1K6OxKLSQUOlqd4Og8JtqzRrGEWSfvygDi80wG6CKUy6
2ypbyiN8pjVgJSHyHQKHWFMxSvcLcYQuPEbzAkmIretEcCLkUMigKklownSAaaMo
oY3jFkd+NH1SVI7TkDq/imV0pbY5/lmFT7Nl2GOOy1iTqjJuemYPeSNT5lfANFcG
JXbjf2HrZ+T3TZ+agR5SWYuJhFnFlZrJEvoCh5ndaDCryqQGeAmUSCfLfrpxr2pe
RqcgzN+yK/gxI57uaNzeOEKEMReoSfw4kqX4mh9xc7sh3ooyDwpTx+E8ypyGKLnp
2P9wZ5WTssb/Auj3iVAkY2xhlxRFXvHooTqRWKRjFoSJ7FBMoCSjghd7TEYPB8H2
8APyqoEIPnS9qQ+n8B5sfhEAoTsbq0YwCphYXzvx94bOdcpNAfcEdMLrqHQGq1l7
EWU3Y5vX65AxAK/jZXx+UOcT4AwR5ccXkkHFlNhnlqJ8Gs+Y3gS2AdaTXhl2vPn3
Q1IZdtTZfx9lYTTyxVkNP/Ho6qFUMl3AuGQTjUjizTFNeQtuJqqF3Gs/mAlrVXa+
mI+H9Y2YhP0qqfyVLPHz3obr8YvAbPNIBdwWvTx8fRNPL5r5hrn6axw7f28bhYXZ
U7ODiZZo2PUd3uYdjCKHz8hMYZwRTkiH7d1G5Nmvn2Xk7P5R95hZWBCqXvm5IaCS
Hj9auhVeA7rHdqB1r8nD2iwurTa2KwjgIvnORHGFi0PK+um4qEaKjY6ddiUZjp82
NQc/ieJsthKQskEWLu/USRQWh/vaU/ahgpzuI/YYS6R/Cotkm2VpuJ0+i4LLrbRF
DCBPcmiYUldKX4VaS7w2RMqBldNaMU0xs9JfL23J2GWOHn6mfFJ8g9lMoTl37oFI
EBO4yw0i+UkreoHjQGOZnmKPSSJBZcBln4Bt1jikh1sCMUm3shM1pfSL5Rar3/ma
z/DtfHuUfM0qw9KeXG6Or3VF8f99Y3L1AjXcpsOMkFuVv2tML2B5nGP1fsYKpltl
JmJYfFwcwsqbbyD3EU8ijlcvP1CN1AN2KdHFC6HkK6pyYDoEuIE+5hcocCzEyRYs
QhgHNmfkZpFpxfuf+P0cPNA5Xdcrw6xjhNVQ5wTdYyieMfkbVbKzDtlL7Sx9YyCg
Oha1p5aI1D+Zu33Nr0S0Vbi1xhMDDVH+PE2XtFBHjlSQ3utGb1/J8PDsDIbAinJv
OgVGBpfl7+04Qh7RATow8/dVpsiqwgnfFRfmlfm7z1ouJGFBJpP84bj5c97vxBWt
hwVuYmTjsl/fp+boHDvK4H7Gga5bLSacS1oQfN7A4mcem+zDaEpSZ/8Q6OdIYmtP
sF1nWykdGQvSWR+8anKSDjV5rQZ72De0H4sOcR29r80EDD+QD70yj4Y1ur3Db0Nc
eVdQ6wPnMppJQaDPhb4LUBsN/6zcFsEUVPYHh8lobzpk1Q8pLqA6t3DGX2p1kEP1
DCHQUywDZfP+X+19FaPFhJO9x7ENCBGzNAb7MRSsbRG9JUVrZhs26VO35Eow/rr5
JJZGRXJ9cXAm0SXuVTj2QPbwmIj6RVT/CjD1285/Zfbsqp9bEqC6pWTLRyLi2aMi
/gjGU7CorI5vXJRrROWughNjCqImlk18lTxjBpZ989I2T8UpX2TbACPXPyGxiXZ4
ZklNt0LKD8jRIqMkPG6EYM89D4Hsx36nqZSTmR05gUuF5CXt00ule57uMvVwypRw
m1mlfqYeeJb675Wzmg6EqHkX/iQ+nqAgm1Tvl5f/ly5Wsh+/4V+y1hdDMIBQFnHh
g1WuZfv16roGJG0VmsUpWMtLOQPAsdJlOTpgdIl7dacvCmEbUQRYOnbHE72Um7oy
EW1gJtK0mFdsQJemZfeEsZhBn24sVtHpcNn4IKAHax/VeqtVXnY2VVeUK7gHBfPJ
sZ/KOazJVKShln4pel3rlzmgndFOSSNQ7igTYKv8TMip44t1P5Q7SvZJKwlnDaug
9XR2ORt1THTHmBzBJjtYuj+3oc+j4tSGMcE/OIumICZIXJ4w/M+hIv4O6hQLf94S
LaXb3WHrhbruvTSlNRwg8OxGr4QuYItiFelic2ECUnBSzZM8WnJAMc71Fu1zpyq6
fjJhzpE/gUM09zXF70YsvtpTbfxACI53GHgWajxoJzms+dVrfo+qZP96hMp/GPnY
/xYHRZyUOOHRnkLY8jTCXDa1xotd28wx5wCUgFoQSl4G+MVOGkQXvFUPJLw9UBJo
ugp5XLNRXwpmbRpK0NWVy6QOZIDqpttZsbPeAJ7aGWU9EgAx+2SjE/7z/yji5go5
zgqv5hz9CzWOdsKnu1CP8DqrhF/la2qb1naQyF1Y8jY7F2ZpPZcW3Fw6oGocUZFP
OJjn75/YVzEimCJQW8/pd41WeDPVgBiJ1Yhg2KKl+UYsOcJAU7CTpYyrjalfZAmB
OEpZd1RCStlDFO4TTQckfloSccMceD1lNJrq3aaIGstsuRR/X1Q9UUEfhORxsTD+
RXiSNZ2qNvJD3krHPQmrP+fFQQOH1Rzm/UmvYBMM2x31p9b/miQngaGptBBC0QSf
6x3x739Y4c5Rd7qDDOAMjVU+NZRXC8S/PQvBivOrZn+Y0uMJmNZakDam1VuzuFs5
dG+s+9lKfiq0EDhfHxvOKgLh0m39mvMThwwPB5T3UtPfm6il7AQLh+CEYxPO1s7V
Ke8I3/jBpjA07ymaW488aHuXenqDhmx0sZeDgYUTV+YUfUlvhEJmfQ84/bMBQDYo
OAjxP8OGkDbOlL0P7sAxjHBPFx32O3iRoWwl/fSJ+qzg6cPsu+gVqV2olOXyG0Zk
/0jsEjrSA7WfnhfU0Xyptg==
`protect END_PROTECTED
