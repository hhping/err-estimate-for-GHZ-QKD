`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TVd1QUOz5iURsU0OZUXpRrqhW2bOUu2lxDQEONKpB7YkutSS/LcdLWygUXULQNI
01mZBSiVZHYTX8kVvk6IpLoJ79aZj60G5dWSEdkEY7xdtJcWecMxclB8KbEniRT1
z1SKKAbFTVG2IcstVkprIXB0mjkznruqt7LzY7UEvWWU5bUmye+MtAk8L43oMKdG
rccNRS+yaJ5Ejl4QOtQefZjH02ejdfPJ9h+wea3WjAkW5i+ODMpIu4MSy7jX0ZSV
YL9uZx4o12ClK8A2iyxZ7CwiHTlapKKEMM9x4lQe6qYtYHcD6Np+irSHklEDWl1R
N9tv+12aQRd48+PwM9Hs4ahd6DJDOZb2dB0ny8gRMbwfVmcqgZ1o9FlYrlQ4MElf
3iyaSBo9/WaKu/VECW5whVwMIBSCcHgzoGGc5mptTlx6dhka6B+dMlgMHebVtWAe
0z5nQzD4jzfyTbhY+8oYQEd8UGHZVwpTDOq3C39ne9KmVmmkQxmx6xGM0m2V82ww
8bVJ2j+qy0PLQyoTJ/jllMbd7/n1bbdqKqa+99rRDTC/RdJUQHyqX1Au3n1K+sej
EquZrN3g3bE207xJuBj7QTSXtQMfD1ZeHSuwHda4ns78I6MBJJZwdPZ9lqWZLgru
XV6L/9GdLT/dhIxcZFVgIx1wRXguuIH7si2uYJ46mxbRg8Uw1YtbZfu5zs8VoGH6
D4U24rYr5/8jnrIF2K2Q0P0hMsV3rdFC+1H8U6G0JgM61GY9Ro+8cvQy9ct9pESQ
3INOU/p/M2r9nVzJbXIyTpAcg1wE+2rq8jtAaUlBKLVSQb2PqySfBNFs7P7Mc8MI
Gr9OWPZtgb5fiu6zd9PO6shbJ/kguMwsLIFvU2XUZf9ArVFXzkgu/JN0PykK/mp3
2qa8XGXA2okekXixPYu7CrB774Itar2ajGhG0DwcR+53rMBHJ9bGu/Y1NVm6s+P9
EVKOx8AQ/KehPomBBo5kt1xwzJ9yr0veA2BCaLwQ0p3wGKrltFLb+/VVGVzZiFyR
JkpukEV3UltdvX4U5xeVHW1xw/FWNVr0xmusI8gPmIy9OyURm/CoyPiuLxIfAUt8
uGtVmblLbFI4omv/XR0m/D3GySi5ccuKsLNT/B/YGo8rHKFcSMZjb7UCl0t4FgCw
LaKgroZSHGbgF/tJZnj9BXPi1/4Tm+dYi62mQo374k7iG4aNuDQefD8KkYLT3Z2E
ehVb9XuHkgTD7gV4Xz9s5GZJ0/YBHtc712KYIebJBabCsYn8HDasSDi/Lxzz0MXR
z2cz+TPTKTV+LDTGb0s/koRDDNt9VZR/24tanyGMmQu2wq+5gU3f5gDGMyLNyFxI
8WFTl1Zjq3F6dfqvWEefE94dq4XBWVDeaU8fPPEVvHEKU6c803Htds8fCNrrHFd5
ERBGmvheDjqUAjI6wJJGxFfjQQZfL4vd0Pi+rA8WLAGtIGtPnoiRrOnW28AYgdMh
GZkvCZeXEyvpjddWp2BDODfR3/3tbfbSvIKOay2+7YajlyvqhiPXRVdVJ1JR1SjD
XnmKVlkqKaLGAdFgsKpStZOAh/EfC2BGyxVzhr241LaJljeOAFtVsx8nV1n2qxnJ
Q3CmQKRh5sdaHK7gMPz5AuEga5qVZQuul0lZyEoUYdP6lALPaDUnovhFBPw+n1uT
85v2nM1WUKWrX7lUxY+TDnOL387Ns7yGFkG0WK5C8eZwWfAp2SMQEMmsG70G1eDn
IuuMoxRvYpewaX24r8EUCgcAcMP/QhhhHcE30FcEo6DVGZDRX4pA4TWYa9eN8jyL
Tu137KHQ0CcRoFMverEBwXQ7IncI83G3j80XwgSiuQfPXt5XyxvLzQ+B4xE595Cv
aI8JGBXsjLmTOrsf03JvsJzCBRcwTGBivz18eBh8Ejkyx0pBpdKA7WQ/ZM+oOtjj
l+ccQvrwk+LK0KuT/b8tBUly+if2D04jHqfvyXdG2CZOO3eJPGGv8BL0xLdb7XTj
e6lvyPXLaqo/tv/BHsY41+IOjnq7qPFdbk5tPBs23p/lVgeIgG5jW++jjntzFeBa
0mGb8YmwlA1FWeC9ro/rOEyw2FIIe8rG4uAiwkYnsiYdxhPJ/bgHxlEIwSOYc8za
sOMSPmDl5WyEbKF9/rLvd2jWglqFRbgUuLGbeMFkQ0LCiLi0Vf6+W3WeN3fxEGnm
RE2nNusq37M5w4dDjNsEfrRQpjetRR2TEuv7chlouUFq8tmY+P0RyAvuR10r/1Oz
j05CIVpSV1ox7pqrlQEEHP6tVvMujKOv6eH4jAIFLNqbt1gbcBfy8l246FYxlk+x
xn9ftg0Djki3Mp3Ksmv6ELhxyw40YClneW+1fVcBbaVnMeuOPmUVFuPJdV5dZ8L9
rNvsgfVvmhw0VJwasfXXCzLIM9UFlpyA1btnAVh0bFP4RXf/nd32xGsDAGbv4JQw
aKeHJYIwpG4HGquiPCJXGoLEGu7p0B7H+ABQUAhyiYbbdvpzz4hd78nK4BUrgYPo
7mooxJtgMf5HfBtFKTiqrDRcFkgstq2oM/4azGp8CJPHw7HgkDVQVVKxsosKWVOv
qMK8cbJ5nhm9Eoz9CnbTMZRw/0S8n1/dsy86COaVAlljs0SFc14Lmo+fS2dc8fWk
uQ4jG+6R9Y7OTcip+ZJAPfaQDQAySxra/1ZAacgsy5GO+ZA7mWKev4/l7SQRM31O
Dx685UFcZ0ikBMG7n5O5CQfbu1p2x0ZxQBiuZriToL4DJDRC0eUMNzrYupls9rai
RLS37blqkBiPi+2HQbcDFiWmBrbrLZf3pcOKG3zLEubroMSHFZJHh8DEfSAT0XAo
DMDSY5At0HG9em1Ei/hn3U5KGc66Q7HUgYHpL6vATGqRiImPrlfW1rDq0a3jKjJ8
i2bZGQnGTImDTKT/FAvd6u0N2WYgh8x6F5K7aHjdAW/pjZ89STQvZweRmlZewQ1C
allMTuFdlUTu9tiK6Xq23jN7L0xD0c01dTyaIXBBO8r+xV+p/VaHOBvGvuLyfNQ5
5rUvdOYTWgqqnY7KFYZttdRxiLUVKWVF9hP/B09yddqo/90QYUo+Ga7dU4EudhL3
70gnGVlaZKzKp5tDTtBoWWXlRFl310zna6L58IqHk4/xVnZyh9f93sq2CPEUgdO+
bbIJMsEh3mmKwFiZx9xu6uw5UAt6ZcxHDpKPSX/URlbM+aSgaTS9W6/Dx5fVwO3/
q+5Uw860caz35xnpdiPyWeMqeSDxVmAqCoCKJQpkh9EX4rzAxXdseaLGCdS9qDhF
J8HJBadNNsS6PrFqtsg5RPEB1LUVxApkl0MvCdFiCcHxh9oIun2TH3bAOVRfiVkI
LNSsQsuIJPLC/R2HnoVnehnt0fGmc3sjv5c0DCS7EqWYpL8e6pVCtPvhtEbRm4Xd
o5tycyrD3VyfNd0YscMjbfPA25fyDaDJ/KfaL/LZ+iQze5MaHUbdEzZmUrAOyW2Z
ZMRDYsj00U+Yxsh1tvQ4Kl0ZFbdnBuLdSFtnG6qsrIoAOg6tgIaT6XNAv9VgxYpx
VMlCiGvRJ2k9dmVrQegAW/CTtGEF75Ydf2t47QISAlELZNvS3wpx3vzWUrwJIKtr
1ckCMe3S2JJvNyF5VocI7ctpaqdEY3hPIS4QXPkhO8rY5Yg9Q9iiWRaubMdPV5GE
lL7CHDj5Y9jheh15UsO952n/P0nWDI+DbA6MJpQNBQl85+wL/l0lvfYuFRRsg74D
PxM5So4TDxTLvwkFQZkl4Qlk0CmATH+eM3aJQ0yv908OirEAnxaVLIr9pxB1K8je
RIzBtLF0eREo2edcG8zmwelD6UeAOL1c1EpkP458BDoeQjCRLgcP6U2txQvbn2QT
uhWMeCKJiFcYVXkhUMvkzrZBfd7qqNXti4yzk6ep8ubSVX2jnFV/UmGhKGp3ps0j
eNM82KtctnzfIxI3WS9edIz08Bg0cYsN3/nFiuDliWuxFnwc9V0N4/4wZrAUO3Cs
OM35+y1u4PsTLNGx180P1WbERiXMzvimyxuG84hR5US7YvrpkYScYeVpfIB0eb11
Nh+G99nwaqrxwVSjo6zFDXKKeNLtLpt916pjLgHnca7EegzM9is61ULe0NDdE0kO
lIYt0o2HWu/Eix9mU2nPWsq2INHGvNzFGoVYkS6VuqqdbThxc7OhDb0BCOQBYEvi
b1eHPQLrGJZ8Kv+fMMyWTTVBSe+W1pi/EVXfX5eUawjC/Yp3q1INJhtSO5GW38D4
9gS4l/q5oWMWURRTJEVnAepvYDOdEkFzlXrUhrTa9tBoM0hzuX1qf2GUfrafAJ0G
y2BIgr3bRlg6sEbqwlkON9EC2GqvLYbyL+WT8/1kLEJkiLyjbYtiqjweeEsPkQto
JL89wbxePspsckslgJvvPY4jSPc6NPJm3mPNlEzkfzcpXwM77Tx6ooQdS7SH4b38
QyPQX6FfsUDZ7WKXIPEtc569q5h8gvliNYg4DsGkAc9K+PSFc8SNouuCozbepOnT
kPA0wcRkiAxKuvH0++SC7mb04FDjqN+3w8+l4fRQV3q5dA2/HDhNnzlT/ntHyYtF
BCHU2sbaA2wcIWfB9IK/aywZLrHlL4TSt/3rD6b2eo/6HQPRb4JLkK19fq8ZwAgH
Ln0sR3l+5mznAeIWjVnj2IgU3c5NB43W7++4m0xeq17Ah6VnRakseewqhOssAI8J
NUN5/gp6ntaJiRK3eanjb56kht0hQaI7AswL+vmeu3BchZgQhHP71nVcOxTlq2Bx
mKvFhJ3dFw3myo1AviAXo4+rGSDLn9vM+y6ZHH+gXu1V1ucTtGFDPDMHIak61QJh
ApzsRDZzcDnwLCxV9agTYRdvVNWBC/H1iNUY4D2l6cJ71MdVAXowKMuOkDiLV1Vc
UXt2djrD/P3OQRtX0YxaN/pYA5O6CnEBFTYy7Rokif5JIdd0AfHUC6GFbahjZite
MZk3lDCITd1Ezh5eVluZHs41ypJSGALAcFwXOGQ2eDLZQNInO/hyRvGh8zr49Ghz
z5rj5pBh7Cp21W22kM2xEpU+Nm7sq6oOoZ2fv9SvZf0clexXiYEQrgZgfyx0vs6Y
tzHBtTOAXCWG+2eUxoLo65QMC9gQkP7MmKAaNmNIMOyu+1RaICWq+Rd1t2P2guRi
UOLCV17hqQXPTNb7hzQenAfExtS/0VGZ5IlAmbA3v07ccCmyE2Ln89bR5FVsuJ+K
aGNZtpCSKUuWkmzbN9cemTF9ZKbGZftA1j81PVWpD/w/gYMDnA3V5NFPaE9chbYP
3szcDnoTzDuTQJBsFc2bmxXt0SX3Lxs0cb57n+jE1yDhF+7uuI7dnlwCyTbwgkWO
xcz8oIeYIIZ23WYgYssDG2IMLs8EQKWfVdsFCCXBl/wpE/meL61xAyoewrpgsdi5
u/SfQ6qVpyA/a8VTB5Dn9HGkPmH9jotDJTupiu9/5u05bk2jUOmOH+gGJv0BYa6b
56JH5PkMcbcTbTetjezHF1YL6kBf47delIUyD5yuwWz/s/LMB+szFPehNWNs5niU
wbsPnoicZpIbO2g54OdNzo0CDPasuvEAzKVgRgUT7300wFYmmpwN7w9hCH2DBz7A
1TJn5MNQfH+qWMAuRwi9gjWkdjWcijYHkPQjL4oPk6DJ0NYUO63w2FJJbFAq2okE
kMAPjDZd7PGyKDNgBLvvE/nNnIHoj8K4b6pNWrMObcNw406hDtQEm6hFB2BEC7Ei
KvTTywzJI8Qwcgrw4KLddbwoZFXQl3tWVOlZjYmcsTLRUwhW4FNyPr2yNpFCZyyz
kelqRkiz4cJZ4KbAa7waNL8Z8jAYclLWFs3yNwTN8vDtT6XwF7bSkl3n8h0oSEcH
41rHV4t0GWX77Uo5q73qjNz6w4UAiEVLft75raKt9sx6jajyI3QrJasG1s7QVmlG
yZoktnwvsuBVNIO7HvmfuoIPu9EAvOumyWxFWVB9hIvTfs/QRRwClHxB6glhQJf6
nlqAUv7WLaa4t/NEDuypoYqhCU/2nJIpoUbJ3AlgpCwOyi4Sq7wBDwjy2dd57zJi
Rx8voNiaPmkLccOadPmxJQR2zy0w2Xe4cHBmS24UXibLsfVex6aInjQE7GlWepgr
iUCOdPOXErovq86hGe7DPQL1umVVGLAC5jly4FtjUob1ZjYugGQyaHvr75Klwlcb
rPa89zH0suWHp1kdNdt1PYBLEZA+TELSLH7YlCrzzcrnBYLw6/wdTERrASOTGBjp
phcGKywmTonRKCVjXUH7wlIddNLtddS++yryjg24Rkpu/zwVG/sNw5LBtb5aqHhh
nPVBUPweLXbfKE5JkMu3zBAQti4/0T290Dti9929NG2xhvlvTIJjYxAfOnedRIuh
J7f2pt+swGX6FUwjbjGna+KT5PWhVWIViGzGeiq/YeMksgDgzhKc76h4U2jBc/Ek
y+ctjn7Qab1otALvXZxngxjzfyDadxAN0KqHjrUH47cusl6myQgh8MdciqZkeqSQ
ZIyTz7UCwN7K2p/vIvoqEwSA846U8IQqRcB/yIgUS9Yadsc3wMsQ0AMIs7thFenB
7cnnu8JCr6FWELKSyJsqY8oDMSpB9qQ/2/qQU51vKDdxZLYNzyXGKvrk3tebDqN3
fpVHldYbz2ytiCS5Q3ulpYpkHnaFuZYVJQ3Ctkg4Uin1PWgS+e3OkvAg8K6tgDjC
VHw2AXcWzO3lz44pLKhCLpjCvU38xhO0v0EGzmI2AHD+FidkK0HA3vgb2YBUcvDx
wuyneKj6dOhncgtM64VZYs74BOWmH2pcBlpPq0Qm32Y4TnSSH3uYSj4fVjlp79Rg
Ve+GDe8A3jL9j62S8iAyVPM1Be3a0hFGk8PEPRP/v0OaRZtinx580sAc6Vp2ylNJ
FtJh73L5+QlM3ly95ZG0VoOFQjNx0RjbaNwJm85DRw+u51WDr6L7cfwio3G+2U3T
ElEiL0Cozq33yUSN38Z6tGtxkrR9+LA4SG1rvt5x4GxbViFLz4+FRmsAPPN4dx4y
HEg+XK5nhmsDV13S2afVPaAv79zLqaDL3AG6D8+QF/Z+uRSVCqIyDn/f7v0jL6UK
l38PKLJwEHGvgnt4Q9euCwFTZQyqob/wJXpNlhBLG53Ho0PMcuXcqqh1+hAO6J+6
2KHnl3GJqC7vTGCct4ibrYBBggpCXcG0Gb39QjS2t2UIZvnmq5/ljUHJ6419AAtT
GsD3C0ufMozUUp+idnKZ5sl0u3W8Mq9gb5r9vqBspEwRueHGifrMmiDEkBVsSDTu
EG0tm5TXJRW9/YJAPBT3kolyToqYeAok01KTi3fgq7r5IpX+lzGnKUIHvNnAdygQ
naSEIasiNKLCTCCLGVHYXbvVnn0GEFAX8/ybj2ngqrzTu5Epk5DDC72l+LAJvtzY
eJQOp5SUf72hnD5vtiZ8edn+VKPXaQM1KzTeZLNEwyx5Nnnpcl6ZuZ4Jras9FK6E
j6qWOtb0GwT2KTMlAxTKUbL5ojjGiBkP2bThMwcyibaeGJ10Zj1J5EpIa9yNhWwE
PS6ZTm2CpAhvw39GkT4/+nVwkMx8S3IdK/wlH+5HjsKSZY+INYFC1yquatGd1JrO
faAIAK85eQ8P+04B1IInqNY0vxXHenrAmo/DCSp1iPGLUEebNiR7/IrpBNlwhnCf
E15/dOBvA6mcXQ01jWU0k5agyi5AD8FGrOOswNx4bDXrsCJMLb92GHENC/zzULV9
UC/wywJHk8Ixax33lloEHVaJztxrDIPszv+0N485EvIM3YWg5OZVqrwvH/NtGHO5
CfQIl9MjKVxqbNRCpr8D6iKYautISE+3NjheBltWat/AoJ2OdiRa62CdhCuJM6ny
uge2e97gqZCf9ezRLIPWTqo17bbHf1jPo3uiSz+Oah+YOFwYz0dVh/A/bj2sNpk3
oBMaFc7t7Axh3kiv6jDLHyGpn9I70XJ0TtCKyVwBT7YvplgtPXqFQnR/0lOhC++0
m5PGoCCDasHan2cbupyTAaJW1qdWWjixWM7aQkFrCDJvXp50R8m8JAgCbom3t97+
qPyhm79vmwPUhiqveqzZxjl8w8Ospb5rJ6mZNBnNApX+VR3A2hZKqyargL2w8WkT
3auYeNBo0hsWOBmxuZcyrIFLff3EQXPJtPP56NeshqDPytOC06PNcCUUjY76Ime0
LHCFVMkgeJwi6cdQ5W65Xoel1jxnItQ9rG1U5ZfXKutPt0kgehe72/3bsK+8Vi/a
WTPN8v1kJAxTys6KIPERyvy8mXmmwH6Mi1kLwNzp2qAHNxl0RSyuK+5WJNsP55tf
PolbpU22SJ3nXLoWf3/7m8ANOYktqErmR42MmBStYV8n4DyGEdQ4ki3b8egRmh3L
ubR33ndZ8zAgCmH+r3loZIuTPYAVkzMaTq8ioOmWEfVY8F88rZfMjPHs9+mRj8vu
fHSMrSkvgxJ7Pu0oZl0l21f8hc70QpTtOMpl6ZOdP2+gk3n7WIwfb3IC/cRf9eHA
6iJUaRk91QmXKvNc3VS8NnX2bjgoYtntc1tc5eL5uN9Qs7nyC3m9aJUMC1nLWZtp
c06ub1rY0f4xfmZ7rFB6bwpwyQAi9hjZRb2D6kX+LSeyETEYAVV6y0Xc8R08yuFY
jbFCC32BwBsrLaVgVDhSlZC1QOwloNkL3HzVSxgRbUXXh81gn5w23rIA82HUHtbm
Ops9tEW+6J5HGAxVoWgEOBG4wrXt2mnf55ahIpKbb3oWn/a3Ii2p8gUHSJ0qHwhz
19XbI8lP6lh9S7ef+8R9d5YvCZn77LfcrnElDQgCx4q/LELtwzGhqclDyCl4zhRG
n3ZtBA9l/b+zcjVUnm15w5/pDCUfhfWhk9XOzWGUpAWHsW6V68bwhKN89v3a+G/a
B37U2UVbvA7/d9gA8zFJYabSx0toKvRorsiMkvO5XEhxWzhu/xVwNl5/151Ts2Yy
fihWWhmCljnfziyolRzI92ZQyuJPnVh6F0tr/8UQWVcjPfO7U9LpAfNahZAdMeRj
3WzJ5GZXrq0XqIMtLKkgakEyCqfeT24o+ycXufLgKovKptZBjVmy9wrmRvZ74zs7
t3/0DDw0QABlBRTNu56zjT47pbJkr/vGjPkSX1eG2uIDKvUNc0/5DId9Lcf1xa8k
O9V2VhSbz9GwE+Qg245UDz24S4ynk0MeFkScuzBi53jGNAeu+4sZg6rPHVQzKd2B
Igcw4SXBhPNSDU9WsZiaumajleFNAdaudZ1rDNx0yA7D4hlHqBN1d/JPHNnp1zuF
PMyNvXw66Q3WHk9I2HGFDDsMkWWJeiakPWv34WwbCwxmcgAiX7uPX1dZZFZyYD7q
5UvGiRZoiYry1l/QkBZgcPDW9Eh+FnZjDAGT2Fl3Xr0gUcQHyZyu+i+1T2JqYbzh
n9Uyr+t1exjZ79VT+M/HHCI6rBr9cgst2Td8pkPulY0iiyEkNJj49T3UBVgfyGqz
eBYE27sNFHtQmdxT4WGpb/Vn0kG22qSH7yoHyARODx1vWKeblJ6Isy0tPCkP+e4d
exG+fpz2qeSwxVxEkQVjJhpF5UJyg/XwKMjeQxeA3iy7nbHH48TA8z+h5JuiV3a1
dfOmJHtuRzsgsu7V/Erkx5+XPLp2TxK2d3srfGIDGLJtxAm1b9M+OinTOVS89Yt0
3jvwXxCzug2QICZLefiMWXxkCVrnVf0l9vRaDznuYUkupacd8+dVjolWP8JigOnt
SWC8VIPYt8PKgTrf1s8HgJRBOqVcrBZBvYwdviGO1Id7M4lF3UEXLqGJSnW4Ok6t
stJS1idsfI1MyNLBqfDExpw5tFEqLkeRDMtEtZ2QcsoaKL1Qs2Fajn00HwVkQBDh
hzscfce/ryygtvQFjxoj7xn30MTubha8rCb/yfaHBFmYDYa/hD8jRMAtRYCUbUjy
2NoBj5FEaQWG+dChM5js9x0kGIHQIkqoyfGuFa20q2v+ZImpEyGZBbTMKoWnb9aK
dTSavS29+01BVu4fqqFdZRPRRTBkYFMN3jBYzS2zH/7QXCaQSlfEQdPZ1ctbgMc3
0gOj5OJUT71GG9KFMFe68bLBIP9Yw/LgpHBgiZ6VRERaMi4iAKk2mciwDIgLElH6
Y0I8Yytui9wFlJZGKVfDLMaz6LyaoGUPNjbkIZhh0E7viVwey8M7H3NtCLbxLbr9
BUs08Y8oimfGhuTfIGdZwpd9KZxaWtL+sYLj6D+TzHPSQYYMcfhOewoSoLoqDICd
DLiEFQeE0NlWWfQNpdKOazksLy21SGR9E+wwEyWv6JEV7WqU+j3xS/2XyV7R7MIy
BB2N44M0rHQUABUXPsXN8+5hPTsPGZU4uIU+Btb6HbjMzJ6dW+156N+SfJ9FCIch
YTFZTq/2okDAKOymemI8YmBq0BY98WZpuFbnueZ+jdgjj+wAU67yf6IM1d0gayaF
Gc2ixg3Yn7SXwuEqLcD7iEVsvrra7fCXx0uNu31dey+9xCNf1O1UeeWCgLGHMA5R
EHoHCnb+Nh10kdMBZ84nDWZQ1lxmivTYRkILP+pa0QLCZd7M9GvEUgGW57CmbvFZ
yTzDcI0mPwl5IIzvXbFP6l3eGtssZKOBihwyoEMiyXTOQQwwxVLma1194jCzCCMG
jB/eYlPrkqPzwDmAdf8Yu4xoePlaZcdQQzENEwCauyF3AghNmPVtNL+L7Wdxq9RT
Gw8jMmJY+tXlvSnL1IvzulXhZKmj8ffFpuZsKA8Am5VNaK/ZSdPYy2AkoelQ2uH+
aNW7jn1H4M1CQ6rg4Wcc67fr7aXJNl9jlOsZ5M7ZywLpGujNND91R+OXNxHQU9ng
Hrk6LINCrCit9XLsZ0gwAMyMwOwB0APbSX0g+V3OFug4e2ew+GmMqFsLeecqpTiD
1sUK7uVDUiOjVWbIund2itjcy48eB8vkaefVKdswusG/XNanSFlbR8QzxV3tsDhh
kC6mFMnlc1LFE+4halphFiTKy+c4ab1kQQt88vxjPZIPChPd4ah5VR8ZbM+ABThG
KSJ+TgCi0ylrLpebbmttpuEiWVdYp2S4XenUGN/7G1ZEldXHgp07j1MP6bIPxFnn
eu2wgRBejpNf/RygTnkOuCH9/kFb9bPLMxX0WdEZ5XrmJ6CX9FwlTYJxbgT1ZhRh
FG98f3PNEU+gozx7fr326UNDwzht7sKHwd2XUsAkDVU/ZlsKl4FpvxxlKdSnd5/e
dusLpc4PoQLa384lOZQJN/8fNWvcpXaBtEsC1IljWfA1FBWEcEpSgmC9N79q1kXF
ZvzYHCj+VDMNraEEqLYSKlq6lk7VMicG2Da7RqGhKo+tBr52qz3ZpSEqWIakU8Hb
9WUbnVazaKf0gbfjyMnfEbRDfws4t+gpUMZRRgcM7VC0IKni1BfY/tnalKye4WRP
wMyIjsf2AvgRItEoilQ4fHXfDcwyZdXb/35LWxit8Uv8r/nOWOD4beUftKURoTEF
6qEUF6jQWXCq7CkY9Ribapue8ii27tdxZtH2CSszH8+P5Oyqq6FVxJ7rw64TyMFN
`protect END_PROTECTED
