`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVPu+VwXaV9Vhx8gka7FxBNxxdPZ9dbSSsshyvLPcK2/8jIZHgBMnTB+NKV5zRZH
rQVGRdjg7vWxGgF/Rgj3Bdn42wDcPQktJU3Y14pD0nJOB4vA1TVhxWQG+tIBO2+i
9ZccOT5zB8F6cY6ekr34qRj72i+NDlDgKXU5Gef5uomkQUUyvosZaTirn09pBtZu
mdJSV8cQ4musYyIvHOvjUtzU76Qc21ZbaLEA3jYiFv/yO9FB1yoq39iAvfj+St5M
RqOk0msm2eida2sfkLQk7jJgBUS0MvYa9K3bnMtEFuz5dM+bicpMTUedgdUra/T9
HOaUGNueVYnfbJeqUcNnaEpvmOTNKi3F/cAZC97iblwaOau2LGlXSWWkSgJhRXQi
ueYGBYH/+wdjn8aRJV2LE//ZnGOU5lRlNuiD2MeEvWCeef5gn2Bn+tW1faMjmM7a
VX/wanf+YPml3rSnsZpPaZKBZy2uS3fVc3sOeSsP81GxoiBr6+yQUBKV2LaZOGQL
IyPhm02rvJ0+pSz6DP8OgeGEaBdJRr+0SX0mT/3Agr9un2ohEqheknA7VCe5FTMy
DCwRxvR3Df4dCbVH0+dh9CdxsglVQd45FqbRONvQk+Nt2oOtF7mRuFU5Ae1FferE
R1K0QAoQ4UOJm2Vztky2vEMxC3GJWw/Qi+AcmHE6H09RGRZtiDOg4IPrCymrYJzu
+Hs6QlonOVv0KQ5Zdsr4qzHCO/nf9gwsFhzZP4Dwx/nXp1VNCCiFEQdx661gWjvK
CwQMbU/ciOC7jXz9swyEt9cdyHwHvPUWBiw2c+YIJYraoCJERa4z/P6AB51Upb04
e+LC9roCa6repalkY3qm/LI+Rz3h5EyAFqZlV82MTViMqvI0F63qDv5DgquUJQTk
SdoW6TSTgo2ZZ7/B1z8CTgHTlIQgOCFUFjpa3lo9l/TBVqu2AnLDJ6u3BvQVx0PD
JeFi0tBgtmOoxp8ULHW2GZtwi7uCMR5iq+0VkMBnk9/ZUUKLomW1NX+b1ikIjqqn
VrmkqW7n3jNwhnoeTLKriQ/O1moqdtJgyk6/fNafbYuo2Be2gN4dWWnYkcZkdt8s
wIF4U/K4gblyz6iLkWTVnSHTZfRQ3fZNJIYTrJ+VoqPu4gvxUrvv4ksA3ee59+cY
sPvLA+UNcbH/QbC/Yw6iHWgcq+L4tzzirZY7y6gBGS7aUazTqLB0nEmsQGK/Q0ZM
UJbZrtk5uHmIXXrY8u+q101NXOxm4tPhvpDXBlI1s2XVVJAC2xQM9Y082gXGxl7i
NXPkXMrqVh+AYOx7fBIinQylVpc/sfTARo4CwUawlFL9wtEJuo5usx8svhnyJfuR
1QwzIt8DhPyyzAKn6txL33KM3TTT2NHR2poiuiQjVMQSHufZ6tuAdaYWYSHH45uh
SwRxInZwSMnV9zMVeafzrg==
`protect END_PROTECTED
