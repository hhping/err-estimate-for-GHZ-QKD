`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i2mblVbpoXR+BAVUGelwe9GZ9PWFMxLuZxN5EDE5weC2rsRLCKWnDnUVSBKVKCK/
i87gB2L0hauyrLTLyg5R/RjBZ/BxcDkvHFq3lMETftTq+d2won1HTxoc8pZJhR9P
I/Tv8biMfYBaePJjLR7mEl94Ptv+i1Ad5vLjGrZ4NJssu3o5lLO8U9XbTjUXV8tv
QaK/Pbood7WU9cmAHdbmeyGdjrj6plrAEe0MTEiq5wVFATJdh8BlA7/jQq+iyoNE
53F8pwTPyLwYG19C9I2XjHDYwUxTJPV7OQLIhfWHse392qDiRiWOaufJymMJIJKL
LOkJxbL9JqlNd66cAthAZQWaDIjLjwXzL6JM80ZRHk8NGTAptN9hwEX9wTEDKNri
//+uyvlG6awpW3JsLv5lZ04rjAaeY1jrBKkwJ3YA/RzgnJs8bXW8UdxoPa7ALsoh
dnvRU8qZTk0nHCmDFz6pYZh90hJKNpir5vXZz9pSpYbop6A/zCtuVVi9fcgj+fSu
Vpi07mt9wbOqsE6W9NDZhi48DMDzMjQ5GobE2dTYGl04ZMa+0UEPKzCbn+dJlAK9
tygzDrC3ZpZvf9vXE9yAsKpYBjE8c+1T9IBYiIb83M+fmcfNnYP2RKvehbA+HC9i
8B9axKLPnowMHIjq4blxf6HVBERNFjjJ1dfqLuE3wtBbsgKOzzGYm04uTJpYss8l
`protect END_PROTECTED
