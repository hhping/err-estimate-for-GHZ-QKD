`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcUpPDsT0SjMwk2+JoNkIsJhA4XRppOhM3lnpVmcZR+jdFTqX1BanSTRdXQInLxW
0sf5zuWKYXyrHEmk2P2QDpy+sehYkXpzKn1LNAifjRGIb8u4Mi+h8+SEbtoQ6Uxr
G7d1QAhoL6apKrKJM4Thq+bIR1mV2KYb8lDS1D+UHsK2IkwSTJjGAclrOQjqISHD
7yQ6UOpugiZOy+o51hIWnIQJmjskP5bQ2GKi/z9sSDCTv0pEZeAkScpiHL4Xy2OD
KHZRs6+YH5YB7W8qXeDHr/8PT2ctK2KaD057XdmABnrlE3ZlELxnqMgzrRopD5VE
syT2/OjYOQZStxiCTFJb8mkvU2cBDaoIzK1EvXVkV0AdYavGvZmVO9iVuxE4i+IF
cFuyom9tdq4NqivRnipZe/Nf6bRfdBgj9nmWfDmjwmUm93X/v/1l3GXbBvtHsPrh
puMUnrp2yTJMlpB6LW1vVm7i9uKEZTzEEA2qZLGibasBeR6NRcGzWGTuTw7uOloS
en2w5ko5WqDtqbXar9VumLUMyZC6i4P+B8PPGdx7sLLTWHnjrxnCyK8JE5Bajskz
nLm7ioMCH680LZhDsqyg3154apykuhkT2dR5jH/Wo6Trr+145XuNnDT35hmBmiTa
YLcUcmyaW1NzGURXUJB4jbBM2/L1IqdoSnGdqptBLHxpKTpkKnB8h7UhiR5qGgXT
mSeXka0kiintcAB3w3J9BtI+Lrd4+YjOEOvOi4oBL4Q7PhGsJw075b0q1b+i4GS0
XT/LonJPoEnbeZxt1kWH6CGyrR0Ah37qvE8zcQmQY4MxVhAmNet1in9byWq73fhg
FIFlQXBhhaxFn5lXS+FKZgo6daexon74NI5L+kbKLU17z0CcSwvCJc+FMjXBfwao
JcaOcnymFjKz42aMAMHMZUUFlEtlrGSMFljiGyMX24IheGBtuPuuUgMkz2jDMXbV
aBzzkHKwZcQbKhQERQ4HVP5BR/FYLlm8vGkg0UlRukKvqviRJqvBW3J5Lsj394R/
eISbDyCixcDww7+E0fX6xEi5qsdFS4jbIzFVBvCAKmjWqyS/lq0VC0zezKSSBRpM
L56sMdYkinWHUdIMqMhU2stblEEZRWuxr4rHxSNvpO6SC99MDhtIQzrJ1dKTfZ6m
dao5/2I1yf8u16s2PVLQ/Q0aqzIPkr8pjcqZQxSOaVcbwoEuSwEak2DiOZro1xAt
fTdG+8KX7TbzFSVrpTKuHc5vED1CxOLMn59eZQvuvKuVtDnwV0o7zCQJcfL/59uU
zh6R5IaUyEw1L4skP5npVpK74xqwGyYpAdaREMxSnOc1EuCFNXkRU6XjSk9BV7ii
Pc5Xnyj9Xl44qQg7xeFT3B7vXr74waBeOwDZNAJnA3mkedcOpJN1FkbNlVYbKM5i
D/iMnMMiZ9apWJbbYm7/YaHuhabS0C4Zf/Mbk4wnw0AWXb5fpopkMM1C54H0jyt3
6J8tdkPjIdKcOt1k9/QXzgLPdaa64P05G87wYjS7lh0HoCTf1Slzr4LvNMhnSIYV
SR+XvRjG58Ms69fsUA/yNVMqqeRqX64olI39ADMM5x+WwpSupzJ3PvjWhdo6ALzz
L8M7cmHlqXJJU67GNqnym1HuScwZuv0h6skf1mwj2klNUeh0o4nAt5e9tztCyrTf
5Bskrc7CcF+44SW+w+g1FQCQ/aFYBckdUlT6fXFx8maknChnvtJuTB8GGuFWUaAh
M3hZ41tzKGuxUiLV9S/fJ4VuAHEadXkakOgErOzpYqOjVdQHzvgMqnfrl3AIlXSA
jR+P+/uztufWAMqCoz2EXz2JsqKCAmfh7cgUgqZiEePairQmUQpxgTOPrk6TvrAF
MdPq61CxoVFuaUlQ4m3PVH8g8yKIBlMsG6LVyaQ2OC0Mk6K10wsInfTDNuN0pK5T
ObAdZQ6MSDhydbBGJQ89K/I17zKTxQuXUgAHcmgf4k5B25QL3cy3BQD7lyRNgT46
rrlt32YmEx/Pt6Ed7AvRqtkpwhowjJJQ9crui/3BP4jCvFl3gB5hiCrDsSyrVciB
fsCKu17JqoUEWCpgr15enHCU0oSvMKyHB0wK/bfncN3SfmZu2ONypsQzOp8IcV5u
5fttDpj2D1ymi+RIYSJcrC3MWrCGlQLExm3gMbZEzGTZFI+CcPwVNNQM93OoE8mn
4KbuWl8Q0lcePfyS1BVVsS9kbW6+dvTu4Qh9KP7MaPedsUtrRnjVbX9S2KlLDHQ4
Xid6uzCpxxPg4EHS7XlN+NKEHboHtgfjYk0XkwPYlbLCPKW+YxGj1Ox3lAGJFQei
7uViFZmnPg8FKmvN4lI53c5j/3kgFY22/TZFs18Q/+gyzjiWi1rZt/O26JkUQUG3
26mRmMzY+LYhhF3tngw4zJ4vmE3S/Wlm0N4kLMg/rkTAYHvTPP+W5CP/dGIerWjs
TBeAcvCfspK8Uct01jLh+t5A90i947mXLFE9PTgS5tdzkQ0YKi5o1EpNYz74dXG0
hEsQFlePpytq1frMrvPfVkJiiVGU20Ozw+J5B1vtFcWamyiQ46rcdCT4jbi883MK
TyzNRCJX6I+dwepEPXoXSu0NQePLYptMmMFM3hykrm79Njyp2PI7IxFRaCDla1O2
CkReJObfPipziH/O9ijUAkE8H3EiAegu//AIASkRF+kT7f4EA98N6iOdWYX64t4v
t2SRwahXa44E6bSeX+ThvIQUjg1FNK5aO4quNzqO14Yw5SwyJJJ1uVt+LBnHIeZm
DV9HT9LtuRuGjhuklIFO1scxGRn1eEwCzjO4HTOY2wmYGDHKpjo5tYXWbHNj0wAn
rUg3os9I5U1oJp/YXYtSq+mE8IJ/PGqojZoVg2vVenxVPqyVYQBZ79vPlnbuZw9x
lYhu17b+Rtvqbpmugdg0WXObicNF8XiPK0vvv2xI3oNzi8XdPXobL9ttSnb3npBx
yosAygF/oI6z2IQlY1KmC6orX/xikKPazbwAgIY+zwByMkPvApcq3HfJeTCDsd5s
`protect END_PROTECTED
