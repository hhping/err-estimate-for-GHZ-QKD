`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BPi1949Pjk6N8jRX5pdWOPay7QwV0djK1EIg4T6JWpLKmc5HDLgCKrF6y22wJxbu
Wc+VztpQPKazMe6lU86u7sf5/nfklaCBORaBmGBs4m45UD1X94fHaZ1xGMk6oe8v
S+HZDMgnObf/P8tFCh7sEZ9uLIrE+woJF7JwsvszP9wa1tfBuJXno9zToKj886UJ
h+5r0HbO3HHCpHs+76OXCwKqLgGaqguZF39bIrl1R3GvOvLxwpVfZa5yZqellNsL
5eI7kIjTM6FFHiRrB4/mEWW/BP9Ozstej71aG77N5afuUXApyIO008Xzs18++wwt
u1nSOM0dSitdyFybj7X8MjHu7vRtCOVde4/qElbbOCjMX2fnlzEIgtnyVriGKKAg
H3w0uFvPV8l1ZaMBxYfxXVOPxLy1gLBOFaC5SAisQhLygnXa3105C/r9lZ3Mj0xR
OP+c/7lndWQ7hVXyE+HZoGMpAu9EUxUdZAF3vievfzyEHNO7Ve+es2V/IV6W6b4E
4+fJElct5V1Vh1p5hTvcvdLaiyHaxCwo4prcF/zFd7qBHjNR1VQveYDsJUEhYUsu
FEiQUDJn8rmsXn30IHt/ENGyvN+rSni62G6t/fnoZlIjAI0ErP3OaivT6fXdLHSI
5b+tB575abSV+crS+LcxOQ==
`protect END_PROTECTED
