`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YcWK5kvrJ00FtjtMlUAmG+sx0nFOvQis8r0fvIvzxPvI/SmZ8WxsJFI0jz5VnTGj
gA5ZA9HvRMlVGol4SVQudQpFHj5lU0ECgzl98zA+OO1hyR+09proo9u3ZM3MmpOc
E4MnA4lnPh2vKelL/yY/7PuN/g3m31w7MQRmjoDkJztRWvtT16oSoOqZR0ZQs+rS
cnoLNl2UkgqPoFWlhGb1DDxSbkUwPOmTTnWKES9SmXLwSprvTUXXFNdT9IjFSyGf
pRXil9f4OxoZ4cJig6D5odriZ7Ftt12GE6WXCkUWa+fEf3y6d8eF90/6RXopIN91
eTlxeY7kfZxT6IGEIYwX6MNKCmrx4ngE69mUrFLgSyHBG/USIjs//bHqxr+uFd/D
aZEHPaJAO5rYjLOJsN2PFX5gect7BBjXHrBuyFDl7Rqw+szezwPfbVcSvOe1JmIT
qaqgQAsBav4HeCxb0AttbpN1D51cgEvYfzVGq1ppfKdjgsz7Ekfj9P4stywraEyF
bmI+I2DGF0nZaL23996bbb7hKWrpVEBLhWSVdLFGu0QjrEVgNsdNFH/SMBYtHCVC
1zFOkkCDkrhy/HnvrS0zdAoP/WKFWRY9djzZv997KACuoqyts4a72OWgUVDzxRtU
PkN1Zx3GmZKXu+C8ApQ8w25+kZolruyNuzA8TLilumg=
`protect END_PROTECTED
