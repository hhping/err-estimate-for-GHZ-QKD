`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6FprWsPp0XJ2dsWioPFjChZyZtqeGm7MAMe7fl9IzX3WGB38bPZfXBn3I7G974i
vDA6RGbamyLn1qcZMVlIlNJ2+mmVqUk50YHtmQreI7vhfogi01IWwISWmy7NC2WD
c2nO2MnDxlz5kgK4C38QzaFZvysmUc+6qdxXt9NedKuCfazS7cMUPd3y8OEkQmJm
hNQagijYq49IPtXsIhOWpYcjVllsj5uVRlYtFxSLir2TPRpiu2HUm53UVCgxg30f
/5WgS05Jf+sxtSrHmUAcn+biLA1NM2DXvTnsYeDi3xvxEUiO+n+uFrlw+6viWNSX
c6sCg2ACI37FEETSjd+wFC7EaCQDTYZ0VSVeKpCm48d3Fru9Vf2NrRsPW4/c61a/
DrCi64cxiShInnADkhyn8SLqvdAm+2RyCrhEkFqceBXQ7B+6TVEsWIvFlnKjxvIt
DdCM7hGJq/KxPxZSvttHJ15X+tguAGryni0Ej4s2sKOea88dRBTgPFW0I7i9j1fi
VNEGIl9LRo7DYTX4GlMrO/Y3+M9GSl1PVlbNWdt3Qz7p0DNmmIRqi0vuhL8F+dat
UW58vweUmnGNIvJR7p7tngIzvXQogCq1j3ZN+qixN/GMJbRtJWetM6awZW5qKDDG
8hbBMSgyppko0fcLNYbXFrNo1w+58E246Br1HOWvEvxP+oNsL2+7AgcPiW29mijX
k1i0VIKDDbT04HcGuIuDvjtblmJZh76yGuCume/ubf09vnHZM7L1RLkgOVSNQk12
gN2D2+1qCjSHEPcBEkJ/AINTG5bHemBqAATKRlY/iPrYjpsh50csoHpHHkxXQCm4
r91UN5Fy0+mN41hQhQmRW7LLFKrAbXwx6WqaixsVqWtbgY2MQNhxIjZ5Q5TkfxM3
pttKeGPLZwrH1tK3t1i4KPhVbhurKEoYLibeFJrk4+IpyIOMlOU+p86bNh6yt1sQ
kRzLN/PNOTJnPtxfA1OI2XKRHbd9C8zAQTiBPr+rjohFVDz8NOHr+jTPLdoadWxR
csV0GxHe626F2JmqvR/dlBeBnbilAZ0Y3qlPKQN0PgkySUyvNkiczPEHZ4dU4jSh
5ETXucCDkaPuaYNDE3XfSP4UD9LkHZvLXJkLW9LDe7ztDu0XHVe8AZCWuZRF+Kb8
nN0NSdUdMuTExu5a61PYHPfuC+4jEWBSnc3PJHl/jbHaHexYYCo3gv9QRGEylaMu
ZpQqXnKWVeTlqyByNOFkQ40ohaY1QSk1Jnf9X3J5aW375cD2M5FoMJSd80XmKvE4
31uM4UxpX71we1GyxDByq92Na+hs1EGQNaPA+4M2zS5OanXI3puc3sswryJD0Na5
2c2z7wy02Qg30LZzPZSwmXL4OImNdM+kc5oNP1lft9qRAKXybvkkCxo+F2Cln3Uv
Rebn7b4VWLIpemC9je+//50+UeqwD5A4RyW2TJvWFLJ4lZXpfGpOv6XCCUmeFVlo
KZWxA6TmryV51yupT8u2XD45f4finZkoUnlgMfS0rJ0OGQo6zerJZQBF9nyPUH3i
Rt+CCmAEyAnqjmRUN3w5wGD8gzGoQh59We61GfDab9TPsXcJ3AW0thONU4UU++oF
F9t+Kx5eQ/a18KNCV95rMziLlCpbsO4rw4ofXGQtxQtCuzHQFqmfLQctb6oVa9zq
BTxjS/ubfxoGnEZwMmq5sGgkv8ZauLaJPAuLnT4URuRUWktqZU2sgzlWs45UV9Kg
ZUaYN5WxjLQou+UDLohnKL6MhY4Uj0Cb8Usvaqxr4sFiB4FeIxiepD0wVDhnoAE/
3r6utHPSTLLEVeedwrh10zab8oyJf1hE6+3MhB3qLtkbDAArfQ4iUtwtjCeNJO/G
gLgBFNF/W38f1ezvqjLnaAQz6EPGwjusOcJZd3Kz2iG+kEbDJtF3aPbJHFtSNGoe
NvYKHJ4EifLlB+7wx2NspN+T7rqaKj1+5gqPjUR0hW4hpDR9CaBBz1VnFPxedN2U
Pt+6lyBfyO8LTtjxNPXYFlz5VR8v7g/AseVJgw6jpBUUnGTMwYriIpmkrP/eo8PY
EHMJyM7SWxIGJhu/5bDNhI8c8d6xVMZB/I7APsejDTbKrt5uXX6N9X3P9sN+Ugd3
euO5WEUpK4ToPlSsNhGhU952fpTLDb24gXSnxd0/KbxOohlwOJT0T3mmjUQ63PGO
/qAOtcwmXDSte6YlCrmNYJlK+MFVDAfcfzo/KvY9W4Ag9f4tFCZ1hZ7BSjB5q2YB
NvizvHJ0gmKxABbCjtU0ez96MOQzoKcVD1IPpBBxaWxDxdP931NLTtWWsoJtHFWl
iu+usI+Lr7qIYjpjtUuzLVXusOx5b8Zk0BTaOJ7KqCpPPeULZY1l2nbrOFGO8mZJ
YwbfieiPBFSC3G00BuQTUz/r0fmKI2JYAnoJCBWVAW2jEtgDZmnmfmu1K6hd8Z5/
/I7pDQNPz4epPxbl4s6E3+i3EXfOpmcJ80JFm365kRqN3c2Fw+ChmDZoow77Lz1C
1tIraLkAUfqbCYCK1nO1uwhA03fRIvKcFgIESSji3VU=
`protect END_PROTECTED
