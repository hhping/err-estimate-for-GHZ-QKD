`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4FOGTk28ds0W9dF+FFM0nAwr89MKqWcshI87YrKLVNG3hb5coG1Y6rhU85KFn/u
J/IrwxCs2ERLHRKLjvMcEASu1QkYh2xBov4YUlL1tQZh/4pzVjWI707h1l0DBtmG
b+JHTM7g4Xfz6DbZb2ygDSDmvW0fDlN4TuzfB0Sp0rLrTjxuOA4k4WukgAXi9Wv7
t6M/M9taPyfVPaLenBXhzjqL8YQyFvdwRuutpT8A0EYVcFfSEUMKyL5mIHxh9Uk+
1iah7tDvRScqRFYAl92ZxTPwktFCBQRYIxX496ZyofnRnL7K5W+7+9rRi41ukmA5
3RMtmWQBe32WMwLFG2MuVoy8MTkN7B/RW7zLqVwTc8Zby9868+OKIU+erRnpVtS+
AE7/BgF+fckQPMKSB15PD1EWREtK8IqxG8pPu5x05fU8atSZxO+FIIem5b1Rwk+O
UwqUc2AZipx1nn7QBq2AgqT6R/rGzyVse9pLXNuIzBfjNQwwerw/+I/VMqaYtfaP
hPEAuvUJDDLZoUkbbKTVZ8+W/pU0sf3i1SusFQ2FVrDpT8bIfT+rlXiyJHjKKVSW
IpK/MR+RZPDYSSdz1cNUcJB0XIFM4NowhXEeYwSbU2YlsfZlkfBYwBhHQb6pkPrp
qvUnlS6Pw0y0AZBGlh2iDiRgyum1Khs5a3Uwqxmwjy23bhyIx1V32JK/mB94Wii4
AuNZ5acwSFaik36nfSfScX392b7iCp+pNqrzKGac7ZdKmK0BJ9xi7Pps1NCgdPsY
1P1h4nGbiyuo4Px7ppqk3MrbfEo01RZC4+tdm9kwBm1LFIYrCxOTlBOcj8xuAl9a
ltZvekJ6o7PL4xKNKQfV5ui4JNzjRy2A6TG0IpZB5UUtT26ubaHE5ZEepI3Q9GNN
cG7gUgyBrJRd5AVCxbCkad9MXeIlCfhKFReCvpxuMWHkAFuUJjfsDKlWZiuzA91h
Q6Qiix48UediQ32i6bb1mDi63E8uu5RmPbeAoK/PliVkYfoThKpInv6hIHjfsRhC
xiVns634AR0Cn+5Y5iI3wWic0vmlDepadW2FoL5wVOnGUmXXUElDe1iV5fY2YxT8
6N6SRauDrhBvilsPkDHSP/3/9TFgd/sb8Gwp04hceudK6ajDSN0XYZ/ze23kMpzS
u9eHGDwiI/rmxPstKlEbVgL0tbgI1ZDO4XU0RzEIGKA5dNtQQqYjT7fjWRgqUUR6
yayDV4yIZ/IolmtYshLviMfpkrslEOrJQ0KdIakHLgRun3cezaQkLTrjZuanJfxH
vCoj7GZa9ztvtUVlDaDc+AGIA7UPy/zZ6ndj7yQ+pSQ4TlSHgAlmFveeqKK1d8XZ
KurUCK4O++yQbzgFVx5QvCNJSANd6d2HOIfsC85raAmT+igq60gihBHpDHhT4dFN
2f9aWZQ0s/uAWA8K2xM8ctSJeOkWpElPxps9jHmbumaS97rO6gWaahHXYWgmNm/U
LemagC4HHL6xqYujB9/C1t5XEmU0mwBpcADroIgx/dyecZX1AhMNUz8RGs3tWord
FI++up80SuCAX727AVyz39Ixe77nZ3a3B+KrDCyGp7XZtWznmbdpPWdxAu5oFjD/
B/Kx8at4PkTLE9v2qKnunxyasuSmPXMamrW840nnNi4XiDaX2ubXAxYEplPG3YQK
ressFPM0AWlhZoLTr6zdRYtQfLaKvSCWiFlJtrg4yJW0g84tp1vpYolDpa1LdGxI
AhQlJQKh31TWqrYBOspcCxUeT9QrpxHKKlFqINna7dlqEciWAQbBlA7K+ce9JUjR
ldV5zcrsfrz9IhH6XCd+wNwAp7Jwal3s9ivozv3oUZHMnRhElAvlOb4mf97wDno4
UdeZU5yr4egQR0IlUyVA6oLMvDOM0LIr7v9JTUGgjowBbv8lXJaGx1/xDWlZHYBk
ofWklRmxMC2lbX5tMsaFpmCceV8oGqAep31K9J1ZbIth0l82EzIIcNF+IsrRavZ6
J5yaWURB724YndiomDDNauwRujvoAHFwXw9x/Rdfy8vySgMfN8ODoijD48r3N4xh
0SujgL7O9MPX74ZyHKx1IwswiNqSL26DOybOezh4Fh8X/rAlCCEA6sLt5RVKxlvM
lA8jVo1jWE6gnN8i9PNDfbaPHRrp1U/vUZnFnZfOyNmAQrqQgb2c6jNjrekPABLr
rqMb3evE/jRPYTb+OkQhuvhUjEiu8LDIpe79so4TodW5axG5CbLYVGXKUy/FKbMg
PyooptkQDNvs8dL78Yj1fknfWkMLMa7EFqHr7ZDTakbapr48A2Ic7Q6dUUjLiuwM
oTFDT1IzLWvzee4OuKP3oV9S4Db/S4/aPs20AmyNOCoH29yPeWfcDtzkcq4TvacL
Z42YVxxaJFcDRBISi/vGQ5DECZ1j1GC7O4ozpvupgdvjOe/qUA457QB8BVVRNBWp
+QaGmdrAp0BzxlxdejruHLQl/3O2njV7ALp0ozjyVbaWOkoplTzbBMWJNBb9cYEJ
wBMbwYO+SxZ0a4bWxqMl13/OECZQ7pAmRh2d25givYXPVgZWfNWAZF8+LtE05FGL
Hm/2Dzqzmi+qz3SxVEc7zOEt+NIenV7/TtW+hi7PR7kWmCF+ILvhKjqNDx7lI6G2
uIoD/lmallrubWXCM/qxWpMBfHya7dCrAk/eQXxEIKxZ0tb85EdiIifo5CfrBBYK
913c1MCKrd6FFRJo/MYfErK0PVNWYQ+oaevyCwSaK66UEDN73gsTo789QXM6DcK2
SePbd8uOqtx27KZwzw5iXamj2Jf/6G5nSNK6Zz2FqhlhYD/QvPPAGye/1NoA3YdZ
ZIRai6ehsrDEVZRhpvHdG7tdNrmBKQfQ6d2LW+qxI8qOvOkPuvVKwfTJLTLA1WML
23OpUUBHT0+3tLhriEg9IFDxNiWmP8YdsNGRzWAQqezZBHefQ80ZxyIO61mI3t/y
7pxKFj7N7PAp4JqKtJBgTJs8AK80vfrBJOO+QHZjxf9T9yKpze0NNT3xb/I1Jvi/
gmevVy7teiktJT6QqwWGQ2wDUTjbQLpEsS5sI8rH+qA0MhZXuES0Vtp/DKAd/elS
JluMuwgcTKGJPP8xXpX2Aq+ahbPeWoJgx3vkwIAhO03yFJDSQ7Au5Zm5byLjvFiU
RTZliLMoAX6fNuRTK5Gorlb7RTKdi1qk/WvxnHtipoCZEwhj98Dru6uCzVDdAsVN
+jQjLEH4JBh/KYSIwBnjiK1NyQ/9W3fv6JGv6e03GZoh4X1FuQObuVuKyOGtQFXN
sj7i4U2v4zbJk6L9fg3jItNjSN6iXZ7YnvrA1IK0yp2mH6BoBr7mKC1mWfE2/Rvl
C2e53TvWb6Gu6exZoJFo20tZrl/Kx7VcMMZmaeGu559MV08orEwHWQZ3tZqM22D0
u4m+iwcMLo96OeJmeitVz9Ken7RVih4NrPQa6/1fVLwFjgb9gMfE4xlDaENZjW2T
GKrJ/33MRUut9stgrUDdGzm4Hi2MT/a9ij1UKJ5dmbWSiWQniAKjGbwtdDMYVSbl
2W1hKaleRHQqTqHZRiiavA==
`protect END_PROTECTED
