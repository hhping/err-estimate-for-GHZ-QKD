`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAqQoN0a/0ejlFGYfE1WWk3kDyTVm3KcL+VERERe3HePsOSAUT05mBIBMj5w+dR2
Tgctpp6+qVOYXtPN5+6X8J1beXkGKR3psIexlGvNwa+bxXd++iyxD9Wz4USF+yC0
YMrHexoHHiN0AVOjErCePEsT7/3Ttk6HRAeZhrzst+qQghMeLaAfLOoIeyk+JA02
rmgYUSNetuGkXc/+6r1ecE9+RmoEjhAbItI84vNVtAifH21Vm7QrD9yn+l0L1xRh
lhQpi4APrrmxd/5GoBmKFkNJRS/D88PivnG5cioCZ3UQ88gcQIBQOcpgluumqr/0
2enJCmX2SDkMeJi4vKpllGyWw0htT+Yqv5ROwiBQy5nQ00mbgACpvknX7a2KwRar
xU2NGhG+ZY8znUhz30MVPg==
`protect END_PROTECTED
