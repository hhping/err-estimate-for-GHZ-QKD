`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkZ4ihiArQ7IBsNXhx8IXoVXEREV1+aXpQQeXYTnbUnuf02kH/85WSHk8I0tbsx1
X0uz8EdWV9+cJGfEOQCKdYd8ckjCx0w3VJRSS+K25LzT+N8Auml4tmrCMbV+jCAI
7EfcAbXmoNsRdxeuGzg2QYmE0QP2MjGuKe0X9SDyImkNFGi78t4jOXOu7IL7/OSe
ltw7pA/jE4FJdIYuyjOdayL6erS2zddu0TpTrkCIjrhDh8nsxaku2xEiCJ6DizEM
Y6Kuyx8ntiV+ZK05w4rcihLtz5Y1dOlmS0yTKz7s8a0FtHbr1wlZ8h1gwz5y8kNa
fACjkfCyovcy5ZF3qEZfHZJpvBV52NHvHcJ990DG4ystJaer44gawKdZT2RZ+PQw
9sF5KR5w7H6FoqsdpeGjc2BmKt+qWU1ogxpt1jGmaxS1Q8ePsYsTxgK3gYkRETzR
Pyh5U132zCTB5Z2oOfnOGOwDzjZafgFQNNMll6CGJRse1B5Mb+045rVosfOL55Gw
`protect END_PROTECTED
