`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w46wnKmXdiMZBEcwJiFi+MJPZztWoNdxRl2X4aZzd13e6y4YsBZ4WV5tNA/urHzg
zmSh1JX9i4jk3ZE1C3R3wRdPItS8TnX3aT8oUx5KBHctXaPOA2Mpx9e8ej0MQWKE
JQOJC8bsvAmhyBx/0Q+TR1tKfuYAKCXY1oi2Lv2R3ZoBFWlyPae2KzBjxEBaQYx+
hbNaMe7rgnEDreTDkfrfo3WyQY/qvi2qLSPfsBxF93r6rYJfNcwqoMt2EFm4BURs
DJO/B18SsicYl2gRKskwOkhcykYBwnkfpJYm79w81PAcWUQHA/iojZuHGYlvACxU
LYv//vwFLykX3t1qONjEGr8pg4cCT8oXvxcHpem3rsSW6QXvMVJTuyXbRh0ndpL5
xElosKTilpXNvqbbibiLf9fTBHjgvMXT2nU72r8oP+WKPNvoPzHif2Lrsvw6Ems5
S9Pb5VHB5CLU3XN7zfL/ipPx1A3X16zTm8w834qN6pNRcivkOAy+orc0Y/FUmR9R
ed7Y/tMrbrh0sfdHfhNzaBPTHLLgbDrl1yRihIUGWFTV4k04mM/GHLusjeq8FYN/
dQGcVPT1KeMuOIkCpEl6+KfasCfCNuo8B881sGQ6LqFbbprXEaNGxZiALJXfbxSF
dMZyQ7cGATvimSU+kU+VwKi3honjmv5YR7VqNfNAT+i0zTVnJl/jNG3rxvBp0Sgn
CzmZ7BsPqI7JqBPrWaQF2r3dzvdg6cAO05Z8Y6y8m07DmXVFyzbVZCepN0kj/03T
76FT0wlxqNNYjCruUWltF5Wb23vyo/UDli0OhZkDU3rayGDQRDwP87sn7m+L/o8z
lCyYA/H1dMWpSvYtNpLxbgHridJfwLJ+WYUAjqOk2f0IX0FcFt0WBYoW9ovEPcOp
0lanqRoJ5FLMOLN/0kojn+0UNkWG1EE12HjYbCts02rvlh+pgWIb226lT1OGGKvA
49gb3hndvyFTI536EWmY4XYbEYZGTexmNXCd1Bwwnw4HizuP9A6DCL8H+ThSgyeb
JWyFtkkAONYHqfxGFuXLG5xjE362oDHomStiM68CK3C0zItPp6w/77el33dYBZY2
fzxlzdDGeFYuyMUA1+ELNf8LaQS+ycjkbwzY6PSe8veQTJ/KkUdlWhuiLI+5TnSG
t4cJjZwoUviYyCM4y/hFA2R7iioMSVvu86+nHa6PP9sNWp3rdozgTEWX1RQDjRoJ
G7ZZeZ5YCdij6CRW9F8hi195qEzD2A0ODg5to2EKSG6tYaLBo9FbvhiE47TgPc3F
epsOuMLuJPm0ipESO3py7eet4TIbWxzWy8Q+1Xrcb3GFF/q+LvMrmY8DG/XjKbpw
d/1Rs+K2lQj4pUOHMO8vdetjWZVD3I8O0fPUnjZJZwjH2YBM/twU3Ahy458jNPqL
M4h/gfjl7VEaANKc0/EdVD4MEcJGnNK+KLqjEgtuM96wnDj7LQE1oEg9DYvGkqu7
d3yR6pkmNxUI/dBh2DBA9f8xGW9o/1WgUxREFHuRIsZlwULIZLS3i8iglpqBISgv
xdBMtJPZIdqV5VUHev5qCdHxNdyn5DQh/6QhXOS3upTIZksqbRvGLk9VsjMGHHmO
f7Jtq8cT+V/I97o7nr0Q10Mu0Vz7Eq5hBoJSRSmz58gbm/AlQHIoqzQqSv9yHHws
GF3Ne1ONITADf9EW/SNNoYJLbzDMjyJgE8GqTlBAOjmxsFv66EA/J5Ja14ic+Kif
aP1w1t+gAVXDXy7LGAUhDE+oF5t9mev+cMYFw+oosyS+KRLyrcWCMwA0f6FX4Vvx
yQvZKY/Nt+HXtnnyyzZ1vGSvN7+BVJnGedb7qhHQtpGzBxttF7jBE4oSCTkkBkwS
UqYugmctcdaaSO4cCRP/wYgptSmLTSsTooyykBwQ3EYUurDY755945joHAc+r7Ao
zJnXLNmVgV96llh29zD2JG88HZxFP+iSFqoS7cTmu6Xk/C//RITUkSSDCCJYGfsZ
WodXpVnvrlmCjjtOtaNc0ktY3ky0IplxPqLLjHLCld5Wscnh2XzGPpSRUbo+q4OB
ljGR8iJ2QuVWjV1kzxI+jVMoSj1ZRXmO9dAV6fjw/NR6z/RIFN8a+DYJaDmSgsbk
wyDg0Ryxro/Ml3cZpDAVHYePnZP0qOrIN6vjoq8CaJiNlrYp/HyHF435H2tEuesb
A6jRLmOpqcOlqTpK4HtS5Q57WSOx211V2SuF4cYdsMwD0HFrmkbxcz3QmozgGe5B
airyhM/lSPG86TjQtyNBokAYlZcZSN7oGY0/L6r6hMhiCjESloFkXEJKFCdOEgWV
/RbOK7RrpX4fvJtw/StcXqONSbjM4D2HbGZTh4ezXbcxxjR4lXM+1hHwPPloqjEM
+NF3+baAiyxDLm1EVcnuS4ReW9a+onfl1TgmEtnGXlxK7JjAn16MWaoP3GXPlffx
y4t0A4c/GsaFqweLQAl8lnnmtUKe0MEpYkVsr3LLPb3efu16hDnp/XiII/yM51K0
Bb7ly1ZYVr6RlAnTriDerhM7fVNZW+fvb+cqhH1onTLKxS9b7d2VOLbM7n1xk8VB
1mR3pJwbUBIVYuSo6Mcw8+uGuXKufY2IurpQ89dmwCGYJ7CEKxtjGxBdQVuW+xLw
Ed/oGRnwNUq8PXLDdV6oT5dKVQ1BpQ5KNOy9baLz5t9Ma9rxUfZYqUt7YbQq449X
w1s4wiLMJNuxBjG+wbVB6cIjO2stJLkiuJDSKkuGKgP5vuBCbzQ0UZesgpDX7qzv
A9nzEL+S5MwdWmqqeKcLN9j7zfRBWeTM/z4z5AmNLG8PuJH4TnfYItLXUH4iavX3
x1PNBTZ3hv8fmnSeUVHBwwfMCzedtZoKBh98pH5YWI0Xz4lwkiU7yAWbN4DiuVPC
9ysUFLGovxgzZrt8q5tzjSkxY89nNmn6KudsVYVM4merZeSpkeiJ4mgoCjCv1nBH
39taacv46BWTyoXM1PA3fsW+O0M0C1sRGoqA8DEw+wbDuJp0vmwMVZYk76GdxDpk
+8h9SJv/shLFxSoE2fNrgC/uOFI0rcUmyRnqaKcKE4IPw5V2D6xOWx3rz1msoQel
tfDDQTTwvwWRUlK0qb38jdndRJbXmQTANhVYMMajNjz2lASQtPBz9ckzChExSLFS
ma4M4w5qtvKchPKTuukYM1L+kqMVFawyS7aThbh13hTix6JyADzfrUrIEVYT3rHh
dR3OrrM1ivbbwxF065FRWfTDBBG5ewNRIhl7chaeece6orR4TX29Wte/g3S1laOg
YDOC9W73OlrPbmSlxrQjIVGU/oSsQrzmFIQFEnxt4aXLUYytiuCoh86bXu+S3RyB
49Fd/kocRUO4hMCU0gSzubATwP1a7L8e1S59CT9EJ/0UX5c80iBC5CDpaqOAz7xl
Xf5J/vVIvgmKWlMbKkBQ/lckJpS2ON9ThlH/GLHeoSnKYLvFMTT1xbG4H7SDPM3x
MrpJGCSDutSP+NF37RQ8zUI64Cto7bZorMPGkekQVzuJky1ShsqS93/Kh94wLxWq
nwVJYFlGFf6I8zxAPZYQuV7unXrbq1ZgI94Y9/4ZodD8TSRmVMZUGMyVg1wOMkt9
F1Q2B6SQ58m87nzeE54lutv3yGFt3pp5cQSXNZfxraaUZb60s+tukMOdR7vQs3PF
xcBfB8jJjS24ojW0OehpMd9m56ofKKSC4aAglctuHnEnA7N6+gHW5Uxh03a3cTdT
04Zc4xu1P7Qgs2WoZTZ81UMH8wW9rzRLiY3O4rAU7RXuDpBVZiEoX0d96hnj+yL+
Ssouxlk8P/W8/LhZl3Uo8TLHh39NzEDWl+0EHwgqsJIzTxad7K1K91MFpEdzM/7U
j5tFUT6zTttdBSkoysd4tgYjDEvZIZfiiDuy+k3vVK3z1WR3Eg38XN5cgvA+tnem
UEq/ICsNCLG0pUbzuVu1yft1z0nlXpO4Wa23y+XM+bhpIgugqLxroCevbriVMJID
B4mtKfmK6I12qa3lYgOHmnNMPbWeH0+PNpj/PR3gHdE6iZEzOVPCLLMt/ahrGWzF
hWGgRfADZk84loMsXub+KN/upgrQunLm67m+07/FYaC20UiUJCjgyFK6Ht1gUwYe
tZHMdOCszsmq0vZ93bYMuy9nw/FgkDhgvfwUbMToqTTiyok8dsF8uTalbtP5Ncwn
NTWvjTfoBiz3N3mXIk51/c3hBf5Y9wf9OsAR7CrCZh3cLuaYpBbjq1BTPVFQkfeS
JBWzFVSFeB+52kZtsoKgxZpT1/+FHweUoC7FyYJ6N2324HVz6qFsa8F+6YiHsTwq
GfYkuIsiWrFxW7Ukn/9kAb0JJsywW6vIRvplVuDMwA4wbOqtuvo+gpResnP9Qbqv
jM4i4JBYH1itdt7diLwh3PkGeGyPrTpzDz+FXwsJjdiSqqInarqdshcWuxrqrepN
OLoEoAydDiLSEl5wsx3vJb2uNS1zxSYzv65ny7+25FxZjCa5M2lYtXZxDUtr+6C/
0/NVMBKV14ER37AVSCdC8yw0Vdt/TkMYBZt9kGrjMN2g3G0ilogWQwmcwsNrZogP
YsmXERPz72w2mhMVEFQpp59IPlaqqYwU4GcOaHe8ZjRukalrrgOcYvUw6Wvom31F
QZkpURNe6rxsKasjED77qJYXC+0ceMs+OhWzV2X+pDUnASValv8X1qLFu/AfV8+Y
Woez4dUGlabZkIf9kKtUIwopl5hHpd6iXUjpxkdhPKEn48LCnI8Biifqh6xNxeB7
jVLbW0PepPcuzDfhTrZE09WPjlG1AmWTH0Fb8h4oDGdFkXd7Xmbza/5NsYAc2QXl
+zOo00BkSCp0Sr7arbsMPBupaQFie3iC/LGHEu4fSdt/UNaYpfXW5ru5D+lfTTaY
5B+RIbAjHwQXVkq9JcPl+47v0l21o+KIKX8uK/Q8v5O0yUvsWd9jP7LnViONiyA/
wnvrY+YwFGDNDRpILiUZQlXFsDYoehI0w5YGBGbX7ggmSNqHI+YX3cXDosvrXf/w
icDN4PwLHKLCByDKudG6oT2nOMSDT0uTQqP0SXllbBZnO/ISnyelO3047Dk50MGn
gcjFIDSV2yzFgWEWEi9rkheJXjkxaq16M50yo66PJ3h/ls9q87ZPKicOiNIhadJ3
2Rl/geRNFLmB1eXKWIhdRmmp5v9Dg9siKDoSPfS5d5og6Z73pB0e5nJPjuAlDxjU
ViuJ8abOGv6pBZUUEfdNJ8uZT4jDHPeG7qfp5EWYy2omk9NjP2+Eg9IN+TfTv2ys
0w8hp9x8/XD85mQAdJsi+mkwGwmXeRqg1CN86kn85QLwcrwYrENQrcVvJSKBPPov
Cm8Fxq6tZYvla1F5cPJxuEhpjA6z/K8szLyVZxZCy54XvYSa5np8CsZFUmTy3et2
DIKlUhJ4d9K7Ixnmb7EtqPHvDj8Z6u+dwdaBYTYgBTrVVm7AYwW553e0kkU5C8DG
MYYXHNeh8/o5GgwLBVxkIDPjdauLq6PH5HHT8gOVpurGXjwLBuzN2xkyBqwtwCCS
6pBj3oaQPv3S1LZ70FXqleKqfeqt9BDjygf3GXE+DZY1zoPxJXNQTFrhO+XzK4tY
NBCUIg+9UHmWqfjbmrjdThJU9kcMRwIFvoTVi08FhEHoYPt2WBEILZBFyGT1NtXQ
4GLWzIejSVI/5q55YF3FeAagzmePnFGg+uZZ0Rg+1UVkGjKNFtleCDQAyxLZxmhB
srnJ1x0HE0Ptwa8tlobqeeoowmisS+I2PPnaoYmdZiUkijJQr0tqj02vs3AXpFez
QsBBqyL/Wb4LuiPs1mUndqXxxaUp2D5w3jpG8xWXHxKt/o1bFWU6Ix62RHHQIdPp
bPpjgwokEjLWwXbVaSq1gNya44XfsFyTbDNynZiQy/FKtB519psy47LFyMi3QDSo
gkoyz6iE5InGVCQVi7Es/nuJ0tWmEKuUKhqf/tR18D7yk0aRkUglr2f6Y0CADXDG
rtf+1h9RSefQYqWmudpHm25h8LQWaSTwqhcyMwttOb8gL5epD+Qyy8PmUiznY1Qu
ww0HVSVGAqVAHNCCXd9U92AIpLgYOZ0e5oO0pYLs9DsjAmHhKOBz99JbvqMAR/t6
e/0GOC7MxxPiya7A86qm86vuSv62vE+6ffwaT+bfWn4SipH1uZzaH3FT0YCxmcct
iNX2oUk0nR/W3V+CKo1Aqn6ubphK9wHgWr6PTiBvjZjcubD52YwnewSIKUKYAiOP
JjVoMiXhYqBAFazIf5jdnyyY4XEIiywI6HNCpBKFWRVyhD3REEzKtDABkR1oO/CA
54ZpVTYmbi235BIX5QIT54o36vEvWcc6QMQHOhwQDMVQgZQKXvoi+tRavHUvNVgE
wn9K2W896UtMkkRvJye7gL8BmeiFdZE3SOltEjippVV8mpxonanMyduMgEtL3ljV
R2k6nrIbNRCS7LD8w8kK/xyT7BNyRDJSeDXo+y0Uiuj78bvLEWhhGrJdvmjGP5K+
Uxgg/ZNit3DNXMiHXF403V6fEN/vQ6x1LA6lFwcD6ZKnAcpMn96yDDDgb7d4PuAY
C9TKjRb9a5Et03b6EPo0Q0DvNkfAKIu7VUb4IrlVNKcsSKb+8290Dfg2PPUl5UGx
fpRVmcIGX32KCExUx39vYyPi8IzTs148hZ6y9IOn/WSj48tSEITeuxclA+dbGM0e
o6bNlBaA5SJz8sdg287YHzkqzLMFGBQS1wEBA3O17ldCbyxrK6MrKyXwSVhGWC4y
epU84oV3EvV0J5zj4adYqxyBPE6gt4T7WqnrxDGlp/oE4OVp4q6r4tmupafmBm40
1ERaPT3d5HJ9D/LZXeW3gTKt9ctreVMdmO22N8sX9lU+HCmhtykardbEmlVyfwsP
WVeJEw1dY8xFFvpT7NGHpeeqGdHu1KPHwwtjGH5VgLVqw8HuAcOhd1kDM/mZUbCC
uDx/V+Hv/04EzwSoiGCmd69uGzwdQHwkap6wHbMUPxuL4eVutq1F4uuHdWwkb3mx
xOUiGCSfNOyjsIspkRsLoI/PomcM1Qk60i3fQzsc599LXYcK/yXdKoAIiC2ufmjd
iTSUVa2IO+tBz4gcx31TtZwA6KqtQG1CeJIsoq5/lrN9rZnnbN59GaHongTqXzdd
ZjFpNi6tZdrdJCl+dyUO4BmTK385x2d+CzIRTof7jVrhtCHy2mZWjR0bpPn51soO
Ybyr9iBJFOYI5giA1V+EidxPfDXOL0Mu6y8B/u2X9WVVj09ZJ0UDpPQ1hVYVWCBf
Bj5VEsc3okJLPEuNztoO/Qs8rddpVxjrnMvHMSljxUV4eDUR5eQv6Qyv7qYrAX04
n1fOgxkrSbaD6zcN5nRmGa1AnxtoGuEEeSniSDbc8w/XhqxxoTGq7u0Fmisxnmcj
aZJ80B6fw0fAEc0itXBX4n614/4reNdgXqgsKKazvej9/JmG2mEKMqrRWtOxDr9g
DXErXntQSf3k2NJFCU1oOWWWByHGf8IUk2PWdZMKdJx40du7SawRY64jHVDjicqR
Iy7fcY7UiXi1us7Wn4PX9G7LHfOEp1jh6fe+JPvC4Y14CHXHQbU+dEMy8kfqh8Ia
fLYMD5+tAigr+azk9r6u7WpAdhREdDUNq+yQM4kTeDF8trSrBJTcWYX946Rs9WgG
kzgoUTHs4BZI3YVnU46wHh2CVvXnrLS9wbGco+xlpUaaT5SfQCYyQxJaZbedyxaF
czLwoc9qUlDJBQiMVvWM/mqKdfSjzNnA5unVjKG9ibPzCQ2h+2f7dopdw6LWMB8m
pFw93aVb+ddH+y0M+1De1ZbsDOV547l/5kwSVN7O2Qir7nuhtmf0+YxxIjLzOQbF
mXm9bWcSZhwBBpo7OERA4dRbtNkB0KPbT2mkMRKWbIrQ9QvQCEx9azPfz7FbXTAK
ETDkPz2fOrmVMbs59JO3YIUWQQ4Y0McIklAxX9fIMwiP3PsEt+SNSVKlKeq4+3bZ
KK/FUhSQHx8/ta1DzhVg0ZLpj17YkZOgGsCCM2MOS3a3GWMoi++tWvLPcwlRBm9A
OmuaHZuDvd6wLEIkgP0jTr+mG04HCl1i2gszWUqZitU6VKK5kvgHEjv6V0FPQdjA
laHTYEwl0+m46mmOO30tfWE4bN/uV+JrLuhwiNERec1rBMPBewMTWbqUECjiFIEm
kzPTrbz6pRib76M8Qh756Q4346g3woPu3q9Wiqq6ajybanphXIN6iYnsNkL3afJZ
PNi1T9cKNVlkZcUWuOJHzKybDMFuE3FT8qw2jGW0HvhXnlZ+ewgz5gZzl8qj78Hv
rHy4DZ1DqvyjyLI0/Rg6JU1dhdr9eNPuVe2nlJR/BM5d7Dehj4O7xqq3nG9N8iVI
v+Wff18HtRzUYixGzqWwSWQRHZyNw54Bbj1hcyT/B3qw0k0AvbOWa7Tc/Xv4UdGK
/KbYeCgXdBjQn7mnL2Raj6zLKXoGg7O/hSh9wEtdNI3ZQcRUOF9QYrjNOIUeIY8b
wI7DENLf16xCjI43sMkAN23x6kMt+MF18bQ4OX+td2uUEotfgk0q1VxI/Jfs21Hr
wIFrgSSRA17+s+w4E4SwJpIxtxXBslxplbajhECrrmNZL9x763wVvw3prLWH/rwh
W5WrtrfOgiWB2IWCJWBEsScagGhoUxyNXNv4/YV3rWEG5F/1CDTP9DP70AhsL9KU
iVJZ7PrGwhUGRlku+xdD0Jikj0ExeYEX8VmdEXp21h9QxOdHSp8t+RK4i3tLOXrb
AjIArWyCsuQOHDIyt5Ggyfw4+X84yXAAb13fq+SoVNJABCSpgE4mW4codraRiTg2
F+LdFXoo0DCWZ8/RXa1d9wfrZLJL3C5wWXonNV+Lk3qv5SpEreU9Hmr08bqVf1aM
/NTE+4Qv7lfXMwmb+cto4tRhgK8BLmogpmKpFbyhLjrKM/512DATe+sX8/6ikK4X
NDa5hxL5ybmpEECkSPDg7HyrunPvJhZNKML6xhNJjvHdN50OUQxheUSerIBWMW7f
d3yKIv/UeLM2PXM019bts69GIMOQJM37j5ysbohsn1NzsMbSov6sMh1T0zUspd8o
9Nk07nBFRm2kJoi/q9tyiYZ9f8WY/rsb/1AuP9SOnYiY5T6eIegO9bwqemDiRJPi
lX3X7WHZ893yjQNTt4OOrPGbv7oKPT6dTRDuO2Nw+Y+JUAzLNm5SgUvN6jLmYssF
wc6YOQUh7EuUDQ/BIRIvr+PB4my7uHWO/jIMd8pNX5gZ3JGV7nRRoMbfVhBWNyGZ
NWUMwwjItUaLBQ+/2r9xL9L7OQjtdySCx8/6gq+S0mfXjHPFj8RUAxBCmp9tQ143
KxBKMZw9qBIlm3+8uMTfrftfQ+uevlc8mYoCsaGwSh+QnIJuZB+oBEWr6ioh1Bnj
r/SYCcwrM/zE0vWnnxyGuD3HKF7ci0OalxS0GI+7LbDGlQ+lHnOu4rmfdY1KXwvm
drd4R5in6Z2bTwTZX4LjSHGjusxKWlLxckA1OOpSKOyZiwkibREFK2/M+xHSSSXX
/ZEixeOZ5ESX6lEqfQVv69bRbsRaQyizYQvYXOLEp9K1NjNhX3ODRu0S1WprmLaI
TSZnNDbphr0wtJDqG7Vdw72uVefprBNKo9iCwuVd7gG/JtWNLGterLBmf/VQDKey
Fv7GDtZPirmp1tcSvBBSjTzAkwD67fhh+G9/lpMarBPXfDQ6NE6oWnoG3RxfN+SV
BAPikX1WAp0ORPbCqVEMtFvyfst5FLCDSJx1ITsXeaI1QHRuV67TmfDlZHDDzXn1
/dygqjIIW56w8FpBJ+Y4207sEk/5qXTE8f5BQ1mGgy9miCLOPd4B1xMvc0XC1npA
W4Jel5hO6aM++QkvyzVVCiAdoR2+uepaxWRIWCNk45IiEHJFhvZhkDn/9r//xt3F
1kffztX64f3nhCW2gx8d29ip1sirOPG0+95liO1ooBV3tnWjW/0H+/1sAj9QTxbY
KOJI932fFlR+y/kcCWy507nvv735rRBfq5ZnWeeb7zn0FJMJ2aSRBATQlIu2Cwm8
x0MyYL+XrtaUP4litaDXhczdso1k38D2dFPywV1hNhB+qc4DKbT3IeB/vXbGWMf1
j8yIdw9cocpL9oBvjk5SfB6QigO+GW+/t6Pi1idCKDDapZsQtOek/sZ89GzZ/mgH
pnNKRmavmDHAHycHrAofLUu/ztsjz9klFYd9qThY5rMzhS6Btk4v+NnN+rpMI9GU
B+64fdYpli4ytZXBFAK7hWKqVLB0FrnsIEQAQVSI2UUjtRNrbM2rtFuN0UlDCqNy
im1OcYaffmyRPni5PyWujBgyIkN6oe/aFMk1dahskLiBCJyt8+qDVA9iZRpuEI1D
kbH70cya8FkmTPytAhaWBOWSvp1u50Hf120f5yUjEHNaJ+Itj++oJcWxnZ4+nJRa
37KrsaiAe4I5nLkvkk8GBIAeFl1ZpkYd1uWMgUrnqRKNnvQoxL4BJO2dEDpCcTi3
VRd8jDyyMu41stcHLbgHnsV2mW8xOyL8kukoHSC8oidqbGPeM4bQFvenJV2Hw2V/
v7x9guB4LWy4Rrid3APQ9kacPxuEaUZX672wF/CwffBeriqpNfMLD4hb34sI02pS
vKcFD6aSZPxsdaHIWMsO4noEkcEv4uKvnrzqNu9X2mgJZJn6r0oqQ6Kc/miEI8IL
UCFhxDwWc8FXXcjTWAGfnZ+L6dKL265YCInKUcykzUe45avPSV0V8KO6eFoVYXqG
tkSRvlfpDWt0ah6dV6kqSbCQjA0GByCbGFaEEFRSYVKwf43SZHjTw5/cfx9n9IUP
x+zuudMFBSefmi95X6Yg1RO1xtjn8ho+qVGfJuuxSDSXpaKVU18tUCJ0aKcOL6pC
jYGOGuFLrpm91duPtt+alWvjstRD0M6o95tBNyu24zqy+yVHLWRHXqoYozFbs3in
/oBlFZmPKkWOu3jHVRFwte5EqKWtIcd4saBVMZ7kFcFXeP/ECxmAKNAnmsXdX/hP
ghRq668KSZJwXDWZ+6P0KoLSO0iFnrdiVxnzzXHOgEiWQwTxxAni8eMemS+NNEV0
nOkqEr0zHzAah/Ir9/imqVhMErbXwMyhOq/CstDxt/WU2JDtPGOH5BvTICthM8x9
eELYUCnU8ym/XmQIBZA4s4M8hD0gbjBO+QVj5oGB9Zzly08DpDm/S1U15bL3y359
gOPmHttctsFL9erbZejFGeCN9P/+N7ql6g6HFwKY1TQHaJauIaGBe65y22MLcYuf
42/c72GEONlw3tJMUibXd8ZxozBSdAAj5R0zSFC/EwuEYN+mwl/8wyLr9GuBEUdp
drEdU7zargzbJ75KdtiAsAnUbTMgDsYcNizB7zw5uN7elx9ZKbFlo6r3OhGNEra5
Ds0M+wsh++VuZvCtpNvsX7v0PKMhf28qd/Yvp1qhGOvTve8mb2e9p41nCpf5r070
hK6Gb4xlAW8chZUrNOzzeBKbpwmTX44BmqMRyqaE5vs8kzgZEqUZQIyAOsjr/9lu
`protect END_PROTECTED
