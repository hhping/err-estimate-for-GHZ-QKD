`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9q3SBOn5gh9KkpSWIIoYYlKXdJLU+WBMSOI0KWkUUbbN8DRkiRePTUk3XrC8ieN
73f1CnnGz30GcZzBTjzelt9ATFVFOkIHehKlie0dvAw2LJ0rMl1gILnSncpFHCt1
Fn9yohgxQ824b9cGzVzUHJHnJuzL4uV25q6FhjBpiOSm3JgDn5Y+nXGLCdKCbs6r
USKge4FXcSVddJqzy6ak7xnUzzGB8Pg2zYaLEi2/ze0BNcloO2ZMg2LZLniS/M5g
PluR2revsnty51xbHuGfNwVRcgfGFR/44O/lM79vydzcEhjyw/+umns9Nn5hm7k9
4VaeQCqKNympMnpiVYIgqqlX5IcrQXTgjHB+sBBf0fiEWyo21LHtvTlZd97p5uUE
PUWZ8gCN7zHo9XvPJv4wyNUI8ti8BtELhJvu0w4ywlePOQ+MuhLHLNij8UPbhend
FmurojqROC/vIcYYCFCLUjMoyGg2UYInXGph07DO0A6YvV+8GMHQT472k2vLvlfZ
t+7nGtdM6vhFhjstY9vGXqcg1ksSlxH7vX6ugRqhOiRlPpDHasNoEkO44gghOEE1
U8CD7M90Fhj6D2phfzD42+7cgr2AamHJrddSJ2l412gnAq2oG2+Xysl3SPWkmUTY
OnofT3+gGa6RbgaNeUozDMrPtB3uWQBAP/L39g/HHSS+5BcsY9yYzjiIvToLqTa0
FhFBRVk2lgcFLDnnCC+n5wnUxufL8w4BG2kupfJz8Gi+w7YCjfbBJa4vBLVkZAgS
KQ62DPx0Dfx4CriqhngFrWSd6GtzDS7S3DkPezEXMVtA3wEG4Eb0eMkdtiBoDD2n
mm0R4FG3mERvQz8i1/mrnWSbHypYH2RjKl/HJCl4K3N+Ksv+xmMiUgBV1kA7wqFG
J/JZEVH9Y52gAwFhQ+2R4sh3HAN5c3aH3+VzEMS/9nBNCMST5mJrT0J6W6jn0p9r
xTOmWWzmsu+2SmKnp50CDnvcCCeNLSvKYj+cydDotIGaFkk6PstEXWdtOyKEXRVP
1lv8ovVrAoMlM8IoUxmTNKRXtAEmLtIeLxuv2ry7NI8GSCSel/9LVqv7JcoMSsxD
ImRKYDo1Vb7W4AA4jQIApLrKbmqg5fVqYfWk1CH6iSl4FNUiKHCLQPiBRxDmNPIc
vUeIXEFOn0a8cEVyRWOgZ2TLelR+UP+qkj6Iv6fE8pAIBq89EXesGDbVkilrCXWE
FZ34M1kRTfhsdyEJ5rUE9lv35YFFvoqNFvjsCShd0cSJ1rj5M3iQuCMHOAySH9z6
w8BCoJa8S6dWWaLxILZiz7fjCJBwDI3S3GWd8y/o6seMBd49VvvDmffTv+W0NSri
c5F3zULE3t0RQQzonIAeqZ8XxyNo2BlLPuq9KQbGlWIsaB+lJK7dE8xeD74cQ9T9
L9qHNrQ7G4RLmKa+CXHtgLIHRkhTRT88WKyYGG+mx3tlkln+oW1XkebJiAQwyUiI
iQJXQfuh8gXbmtI7kYAHypUuiYnarIs0lYSurYGeZsi93E7XvT2JrNbC3oquMkHg
uX5izx9mvYpxCry5Eq9xGsOF8aZ5tkY9FDhJVQuUm+uXrGPAC+ERAaa2fNXMRLJB
70P2sJrid4EWeVT/hA8St1l7667bXoQVH1M5XwcCWuA5Bei1kVuvBm5UD7ao71bN
oSNqqHlWAwVK9FZxmXHTegNOlkSxLXw8rM17vJVIoLis3NWEo8spS443RFp4BJ00
HAa+CqN9arfzX3nWGFYysMXJYhkEZnamZQO4FZ5Xtd12Dc34+/F/TZhBqZQJSM06
/QCH/tk+0CT5iJZDMJ3k9/SfVy6kKTnlGn/+Rn3JiGtC0asG+AARjC0hF6Qa920D
IHufV2oKqISQ8yuZ/uF+eoY06CROJYJmi7M4FjX5Qebbk2QkYxrJgiO60YS1lItK
GDntVVMqXoA9AUJMADz6G/lNuH6C8z7+yBB1CUvHuzlv312SVpktGpP99VGk3yWx
R5FpF0t6baok85dXJmBo8uTSI3iSdePAEBAuyU0Q6oD0FcKsq7ZBTn18yseDwdTo
k7FiG6Tviv2/OJnCI/AXmZNGOaW7Hozq/H54BCxDn1XYUy8Xzd4nHzZC3Nlo91jK
uYrLrYXfm0MfyThrtBbJElv9q1YPFqIrFM+FA/EwgaNtob6wP87TSA2+vy2IONd1
h7JJN63u0dCzsJfqpt/Nxwq6LXY6zFWlhgjmi1O/CqLjxCzgsdtO3AL4Xdpxx/0v
P1i3SimX0IjYWfQ5CGs3eggG4oRbRXM4RV73DhCII4+th032CUsnwr9tU1fhlBPi
dWTk+CcD6uk6mtEJd8kQXEKIe3tLQwLau8jakd4J7HBIYroJSvrtE4zdgliWVbSi
vEAx1I/BEvAJkqUnlKPsADy9Xx03shjto6xn8eprXHb6jUXvoqQuYvFSn65v/jX0
Nf4qhXbm9imyaq8cK52Bh9L5l8HKzUCDxQrEhQN6JjuDP+XUgEoz2dEAeQuBjH5Y
+B7lbyV0f4RvAZePg3MsNQ==
`protect END_PROTECTED
