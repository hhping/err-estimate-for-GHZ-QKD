`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
np1zrEsGdCbcKpHw/FXnuIxfjyvBqQ0JW59BuODn6gNLGe9jaHay98wl0PhzA4Mw
Rf/27wNeqnxw/VqZ0PaRfAtbP4lJyMBiw82wNb/jazeawT6bwOnUmPTD0oC071wS
7JRP1Xu01+IV0vf223Cp/PiB8BfAVVMV0HwcuwQjAa3jT9exsXasaB9qRrN0rSCd
cYtrJkHPL+MvK5hSyp3dmHNanFNKMm9QDa0qfwX5F6G0nbFXjssVB0rWI4AwvYE/
k3cagTR38sCElZ5koLrHnsyb/Uq87qZYDoMlXEVnXfyXF5lEyiK+vU59ovqV6r/E
JNIlazXBIYm03yQ8WfmTlfXk/vyAk3QH2xBpyydPdgx+ubee0rrOiEFe9mQc1k0R
dsktbW2A624qFAdfqdxliLOjEoYxAcMZlj8hv5ivi8pRZog6alJgvzTgFaRPWkIP
zaxdcfgdSVyJ1Jv0smaAgD0eD/XDn0QuBoq/V9LjYaIhw5wkZyjiy0X5RV1i9sBu
oBDvrEIkYsqBritXLwh3Lrmwl5LgffhRfEy+Q4UKQMtmkFGnpahAiL6u50ggGz7K
vcxHk2WWDCzN4N/JPr6L/7DoZVW3GAQzxPiuahUOQFdObJcX/wxkdsbf7LbUVjZs
Vr3ardkmyBuE3cu7NZ1f/iVbh5iiYfaEEwGUmtSOcqnxySE0kKzDPHGTMhPtiKry
XWC5c4qLPtH5YMzNHG6/nPUhA8hstkSM6irJsI/d2hTZrZ7WVRyAe8ZQSma1B8Br
rzyvK606h96jp88Yq2q/Bos4Yxs0IdK6dZomabWc1Nl2tbt7zNqzo7g7GjEFQRvS
0/HazJZdaDu50QNiaXV+eqBB2xlgvKC0UTOMkN6imAYdz3eXP12sLBeu6lcpDY43
Vy2EIzNZaj4vQlpWEORgW9RO4mZ8GTLEysBzwAHWXNtdBuFMISZRZVS+EyhQ8fpd
WVb8/mpyF6oTlPNpyXNWaKVk1Y2oBjT5F9sq+2GAeJHr2BQF0oXuLkI+xbuJWPMy
KFhNSCehTFl00xiyJlx+1PlHXSIw+32JyBJyPlqRx1e7ExDvreCFRU1nIEIoGlOO
/hQlR4XWZD3d0h0soxkwfqWACRiS/rTqNkHhHvkfggzL8DruRJf2rhMBzEuJEWwm
rkJXGo7WlD4ueRzz0AZrTYu+ytVYJ5Qgc5n1Ic6L+S5Odq5WRA8mfCahnxty1Kpf
5tjm011Yxd54Nh+xJC07GeENSyoJGG/sA6lKTdbNC515tVI4wrfEkIbyD0Xda3D+
WV/BkocbVHViyt19PRLMMo7O5uLuW8cNpd3gSOODBmX7ER44qZLk8KVBGkxyXodT
KoMhSQsRARrgFUP3kqGay1BqTkmb57IUL50FD0lVB33q2uCfo4h3hnCo4u3byi9W
GrGfuKd6q5aCSvIQxqUXId745e3lMfamI4ytdCr3Q6cMxu32Vy98ahax8wxXHh+n
DQpj5IkVypF3quEONcCAopm1iTqPJaK9qcehDxrq9IB6qYazcUYesiKu2RIkjG+7
5rYCLH5SQknIb+sa7socrU1bdwH5m6+Cn+4kakqLIbmkjyCSOMS7BLwNq28YwC9D
9+nv9+gsCXNbisriABbYGTs4yA59E1f+9ZQQgjpEsQ1vLcbdv2Vzva2ZCyW/6KMt
l+JXe86aEIiHLecgJFDMfqQiJCWytxNWmVXmqlyDSYSAyf0+ahMCEFqGVDnM9QTp
jzu8Xz4OnAb1AI6CH1bQAtuknWeS+6DnFJ2Wno/j2y4JcsLNxuTRBHpZ50fcByRg
BIbTvL24Rq50ecwgKuASd/Rl5jbXhnZ9F8lTFGznHDZMEc6XSGlE1nqclFfW3oQf
7LvOoOXBwrPZ725ZGwzmUGF7Bpar98pn192388yGfC712LnFfGqegrRgQ9It2NNj
6Zh5sOJ+sIUR5yMueJUCpn06JfVWD8zFl6Ax8Q+AzNDyeQx8zd1t7IXlS1ZUp/5d
hNDcUAgUb0oLbWsGQ3Lfr8ZKxmd6l61Do2hwQ9LuCfJuKujfS7iBDlnH2XRiqUa7
2yCN5nCN698qhe4Pj9ProOy2Te1jX8rKraTdEubbsuzoMLJM5bTvJGB/4ulkhhG2
WuZMldiTaJXMwhAcvo1/3fnG3MWUAy5oi4WMurk0hz93flHHqh2DS0tsv5VZL284
EpwszJ+eC+53D2+yDkTDk1mk1h1hhnnfE1vWgV9u/SYI8y6sd0lhNCIpJ8Hgi62F
928az39QyOZwUnNaZREaMR2oCldRk8WefyHDMfPlMlMV9l41RgEpKf85plJ+hXyv
bUOuEckYhGLllW3Rc4hc9D+Cm6p/AyqY/aPnZKTpmewG7BBI147GECCrynm1lPVi
5rhwCdYy5RW7Ewea+X9AnTWzKROAmIs558+hbfR0vVDCyEi05LbAf2s5UTUYUI5L
Q5wpR549dnvPOgbTk//rUIdB1x35sUF/NVHMl8ISkthvx6PG1r7Mn/Xwu2j29gWT
nU0DS1pRGcKfWxMyq8IRMK/rlaTs2JordOTW9gVYqE9T9Elo0n4r53EaZyEZa9dr
+gQV6OLuZhzok/kCMT9LRDPgLmTkMMTaXZUn5RxA8VePpucRKwTq8CTRdzt72DHn
0drwQ0EgwvSp4CfALLLZvcha91DGnmswVI522cUu2ioD3/8WzM+Z2GwniNAMQA30
paU308eHqaGp9mjdnCTOhlDt9QI1qvd/1rj62lSbRTh0cUiQoeQfDslZItwzwjDD
i/DXtvS6LnNXM2GPIBXD9UenkXXv3Z8wWV3SJMTWxD1y3/JLGRtfGxO/WPPcm+YQ
6G/ZX5WEYAnSXHiUEimwlCV0kA84FNpFoS9j/aZFVf9kPtQ9Qmv4hh2Emf7BhfEF
GAJdDmE9MrEEzF0E8H4NZmrIpRN7MDBMblJ5CM+DtRwuG/KXZbAkISbfI9M6Bw1S
R8IH+rbkth6d8XAv1hrp4Lwa9Ki1+hPBz0+qcKAl9rZsd/vguJSGtq3q6SvntMEN
gfg2ulkv//rngSjWRvy9300c09Y/G1N86mr8ZF26hwXIOpAr8ahCpRTMucqLxApK
FRpTIhzj9ry6ZxFz/1UzL7p8lByLLFpTPo+v+rw6H+xr8wE9itKOstIfTrQzgxOd
had+XKwOzi1UbQ1rrslxsVTMY6senK5D+w9enpXqYUrAbGEK7OiMk806l6/aMQFX
X3NMeZM5ju940cN6wn2M4mnJcTe38Sz+pp4Nm5Ic7fvdTK/2nygkyhxl3iJmzSbo
y/X/X1sUEM65Wzw/0xMS0Dm/IBHucx9O9MZzAzXGVWKItkUr3y4DRuqtr5btyNVD
Cbw0JuyDGPgAOn38HO1e1puuFQyxwrklariUAZjtRjiXfK51aAaFWJ6jMgqXjlKG
VFyaQKqrz2afueGs6YgrOopP6E9SQWJkBNJZuZwnswkz0y0Jx/CGNvqQqd57LorI
dnt13oLnvv/S6NqY9qcFZsSVrRw+1gHxoIM/0vPGZ6cUS6XH+QK+SYpG0tbrwADn
EiEGILpwaeffp9G9aOTEx47ePpADHtNDJwddY3V2rnNQpbKBgQzeDLcq+W2f65Dk
8AXO9ctrULbnPqboKzhOTmte+fOjJRJsMST7cMJ98Vk2ayg56XhMjt2xCMYIO/EB
VhFaurR++98DA6wvwhFAzr8wqAbjv+J/RylyG125JZhpZrWYblisk2Hj9g7qLY7l
`protect END_PROTECTED
