`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6Ze7orDngFtNxylk2fsTovfmOcQiehFSE5ScF1F+Jfrm55U/fCToITKuzEYMh8o
ui3E2Xqvl5BfeUUaeNgdFZB6+OerFvQzESgeiJMs1QcAy9ZU4LbZ8DJha8ncU7yG
2QLR7rsl4estixP/lzaDfXFQKDl1iekTkablfVUOBJuBj+PkreejLGIBparzcGpn
3VtXxtjlKAkCPPS0m2Vh+TJr2VhqsYwE068sXxrSAoqz494k1fMeCwYTQvqnCfvw
IZ9NEk1CAVEJoFBk1izpLBigD0vNeSb3Th6hF0TPoZ2V/JmjqMrDqAqmJys+r2xN
rAwmbZ77WH6llUut+ATyPt+fsU7AizKIyWzNHdKrfLnSbKRC+gkWeOe1Htrexiok
/5O072ThTk5nz8IlRCbzdRWQgDzG6ESTFVIKWCPmPJAW4LMLtpM6L1wi+kViZ3eH
t4MlQu7DLGuZectGJn2Lid2xEKCdqYodQjggZyCQSoHmAAQ7XUgnwAPZYTxeCkus
Ewjsh0I9riXRhS1USme4EATAwFXxg7gDG0vJppjXQuxgw0vHX+uGyLAn3BhS+Stu
v6Y+Ga9DQnPMf7+Nqm/dDQ62z+DCayzxcol42ccwieKEo1vqcIkX5R+t9iMEWxd4
ZAYziywzc47EnTeA3yI+mMPcJvMtV+tAwD52v7dUtgM3f5dMWvrbQXY8hN5JnW8F
5uX/Mt6IR1JbZOqLHThMMxxmb234k0cbKDGrrWYQbECaZF5aTqUOaERKY8WKCXSD
anCOOk64rfzbYoBSA+GdTZslyFD8KIpmjIQdN3tm1ysg5PcpPWBF8eMR+i7PIzpc
3ktQ91foZg6IbNt5qO87tC7XQqfc7y1ehYpFl9Xa+ILXFgEQBIfLsi/QlaogWwgh
syCzyAxPoFIPbq6ZF963n2St86oao4/DnnuxiVBBfW/XSuLLGCAs1HgeJUukpiRi
i3BNRdddfmH4jKEnWGf/LzoMPwANEO4cIXcRZDmiFto=
`protect END_PROTECTED
