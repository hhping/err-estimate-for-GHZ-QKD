`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+To1ppsujl/1YajSdOV3taY7AQepNtyhTsi8qKJ8anitj9/EYpCEeElndayNzbQD
ELoXSa6qaPbCauDmQbfjuU/TQUyUwGB0mTGzVCb9xjhISreTqJWFn/GUvStWfmPE
JKbXJ8Y2DxBuMO5urhtGW1i67IONrcfZNdOm3Cz4tExgCDRF6LrSWrVRN6/ayzwo
lQCcFbXW62Mi2BietxPGGqP6OSp7Rzd2r554V0GKsExwkm2aOD6VWs7rEMINF3uw
cKKeVVfYUX1tzZpOanKwwyeq55pcyB0HLHUvlSNqQNSRRmW71dcPlcbGGx4fptAp
fca6LMvntrR9cUuKr4yObH7v5PRuGEJr1dxI8qtkPpG/3bnDbyYWNBcu7i0xqUXF
ykCrT4xaPYFYXHH9IW1O9/hqfp/t+eftQmN2CxnET4crNi1ekRBelLDq3G4OTHrM
ZN8DXHfSEf8pvo/ljAd0i0QpBgeTM/Hdg+DlD0FTXtNYJFlhIM+RC0IzysnPaJrT
ui3GpedkIFOdxBRM0WDq4cBChCNGS6UIj/X7cdizcjQgJuZ0O255nyg9/FiC4xUe
`protect END_PROTECTED
