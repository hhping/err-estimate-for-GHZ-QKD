`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YUSPyXi+C/hz/G9shLbvuSoFDiqrw+uv8ocuDr0CYy2415JGG2JxHjgRUvtybC/K
CxZSVGYNcFujRrTJuyhUDID/S5TXhdZ4o3XwoBbTu8HRDfAx7CpvLDni87T8FFuV
2xC/Aa60muxhTelKZn3SBEO3sVnHKRIJB+4mA+3vZu1I1EhMGNhlAMRV8pdyzirv
6Uok2rdofTFPAs2ejsi1DK9vBMgFD8IXklZyKXox0Ss/vSnsWdkRw+kZ4xQ3gu6V
wDtdtBYu+FAr05nJDNef1jEZI6SwLk1GwsCtSoEN4TLrex29ouFEgNCyayivN6Qe
NguY0c9vRUqZqDCvSjYrJ59LsS+FlMNu52jHqzAFScyitlljCFfc6H26xI7Nxvqe
pP+BmpQj95Kxtib75W9E/hNIvYulD4errYyCkd3p6prICRhPOOuad0OytWcomxX8
/hoVOiLoBLwFuRw3SzcoKvVVd+C2+Q3dFidBlmAAgcWL7Fkb0/KlAWNiIfXVJ6Qg
g1LEGXrZkoZXTXbVRWTi/psvSGOpYWdnW4XO0SP/eHrNnpTWy64THn9vWg/50sza
`protect END_PROTECTED
