`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
465zu4qrHZbme/lYacJFrcBFqYQvrju4GPU77yYKn+53u4zNv8U8kzZ+tKJ+kvWQ
5/fOgYZQMFKEpN3f23BZkVNk8cEW0UErO7lJ2MGdca7BRz8MqiSVioW5EK2OBhOS
94J2X5N1Nb9edUbfKroy9wmnKLTzOJSlsjxNEggQQE26nQhfMjKLBo06XiVRBK0Y
sFPeWpSAJWTpJx72y4AngOMZCEveGLc2tmYHvznQpDu/JwH7RuWx1qRPgwagErSm
GKCO0YIlXKUdPumBSpsepqZI1ygFWfc03ENU2QVDGZR9Mgsg/jioqMRTPa+7N8ws
Mru0Ns+aGMx7l7udBH0c9LndkB+PPCHApDX70HTMBcB/gmtw/qzhD5MG2jhFcQrq
4KJtR3VoD2iO9vs31ipnWK8oJlviGAJYhXV07xjaLALTp1w6Ao2a0WxraKcj7IfH
9Pwp5fXyH18oSPkTtNmkqI4wTkfmZ09DUoBMf9OYmYdkEcCirXRLfFyGQi+xRgct
sj+yq5nf4waijAPvv2RCmgxFS01m0F7XCRE/RKi8dMylshxgJJph+UOZzLN0crGe
l25VZMMZTkuKffzD5yT7cgndTxBy1cLTRozGOBiiaffkjOsXGsMqESz//cirDs+Z
Fzt1LtwnXspDYAAuDKtx+tZmdf3UGM60mktoACUP14tj7LvOAcOIy27jnZmG+R/E
YnxJX8Ka6/QIH0tHhFLiWKmGazS6QQPW0ubkjxFivD8CmH/F+pEYa3bE2vswYmFA
MssmJNM5IreKYbnyAsYXaT4U12lwDIbnuI691QuGC4J2zfhIhe7fiUHY87nRepgR
xePAjp/0QvQl7qu0nIcq0SzzC8AH1/fmhidIZnkBi6mY5p1n47VaOG7aOrS5eiLc
x0C+mHzdeWIVpJve1PKE4Q6MLohqzeyWkRs9sFvHqIinrGCXBthNhYcPt7U4Dfjr
YoLcrcyLHaWDjlKexWct4g==
`protect END_PROTECTED
