`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OCEN7DN5HdkOkaI9xLxJPv4p6Wuz29Cx+OvQN55p95SmlVzr/8W5POQfiFHvTS6
Pg1p+pmzxAE8x+B6dHDGx8+bUfs4OXCzzXGFAqlnuE9C5vR0Sl8FptXwqGdMVQo8
QU1Gp2U8mhiZpwA2BNqrP05hVyy0yVUEfIDnn3rjjy4SJd4rXf1J1SEDYIu/6yhm
6fe9H6xwAjUDR0Uz9AdqFA1pJNTVgKyaAzzaaCymHD4ctHoPgCIPlgP0U+4/zcEE
XgeUhef5a+ZKDbwtDN0N0Vd2xtNczVWAylyVKR4/OINP/vFKXyJ550hz0icCusPY
amFBjxJbW9UFBIRjQ1OPIPHDuU+IhaDjVFRTQVswTK+PgDROHhgkh8Vb59GbNx0l
LRsEkwPNsnACE+A1IwGCLBoFOkF2gzebFOHE3Ayh3gaqG+BKpUt0QC5ZUIj3/HS9
TLaGFNA1keZquCspVVe6/C/ZRWn3ohsuTHD2F/n3z5fMfB//MasNDNVvCfxpbxDS
VbEKOSS/3aOAUybzTw09zA==
`protect END_PROTECTED
