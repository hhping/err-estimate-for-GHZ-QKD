`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WR3A5PNxtSKY2sBrZQ1oNWWDUrNjUGeNevKyrAomF1W7OCV7aKF92rLBI/liE1xW
ccEJ4cZnLIM5C7GwKqhpdBZgYOMpwv9GCCag7ox7VaERQmou88gDytNObL59JqUW
2gzJpOZMOPSAV9bwnoAnQxOFxn4KSv1a9utbmTJXU5qLIej4XKY/yqqm0G5jy5IZ
awAPfcqj9QHbAnG9JaMVDsd11a5T1C+FIlWnvlNy6hZ1rbLNjTm0XZqX6Zhlqxms
qkA0YbEr8sUaKVsK/eaeaQ7WijLhvc0WQqaSFVsiCEnKQJAjrfENAS8WfUqMKx6d
OnUpRfpvnpXoCEbEulkm9cewabFo7pDIcxIl2XiEI8fXgCRytX0G4KqeUKplpXVb
l3X8P9x1zjO/0oGD6E4hZ6X0rlV/6oQe6Q09W77mWbZOcy7wRPu1U4tUTQlh6XPv
5x5kPHODQ3d3/w4cjEAsulWo72mmnLG3gH/vJBAdiTq17pRmpEFhJZ6VGNmr6+zO
CGHFXHfvbT3Ng+LJpKdZbC4Qy/ps2slXNEFOJI6oufzwRm/DX548q53TquJLX5I/
r4dDTAXQlxbmYoDJjtQtgbJrJDWsai7yDenEuGQRcCBLgGqSQMnXx28edQip4uIm
puN35kRxxNDoI2Q+WWJiJvV3lgASFeSLgS7wShCnx0X/D/e2vjtJC4L6GOEBRCsZ
B7ctoT9UHA3BZlJMDE8o8YStFd4Vjii0HoW1oCnlRK04q1+ya/YvSYq9ne0lTQAc
`protect END_PROTECTED
