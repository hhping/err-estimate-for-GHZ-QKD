`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lvLr0KxFCkDahJatnZqX5w7SDdx8PQiFkMJmCYNLTL1yzoJVSGdtE/BK1ccLov9E
6Zi+L59LtRNj5P9MlGjcoyk+DWIqnZqB8MJhUMHeMdFEttyD3dYlrwP36eWH0j8F
mvsgCFOiiok0ARGfOdYTC1yOLvEDxMrXeWIgclYwn86IobeIjoj8B3d6hjQ5FHRH
ZuVVYTGuOwTnFVyHBePDuulafw1qUlZBTmV0ekkGSvSYW/S/QTq4t3lVKyfJXy9X
ewOXjdthrIWCEKJz4nxAcoYgjhsqCM4p+OLIWn+cP8F82MJQUagPm7suyzFExbab
OsIIHw57MfY69h3MIISzD8FpjVAAvHtI7eWyIsSVMwGSPfS4jM7luE9hoQ9Rc5E0
2j+k9pirnCBT2hRuWhggc0HAmR8Y/wmvDRAuGpbFCVqsuf8nHxfKoJoWeqUd8X3V
Z8bx0b7SXsjnVAB9T3igFGBmAGV85CvjmWYq6pQByeM3IGr7pkLONOzrOL25KkpE
rvnkbrawSVHWfCxwrfYu1J24w9Z3SNXJPdxvZJcDi63OICzKoR7wYzmPClL0ZcRl
3vrpa1dlslEXXZD6unTy06j3I5JUUKarclIEEZ2KBOdkZCPKbCORCp/naBrigJQo
/8T+xKG4M1cTrmA09RzFNieFOVy0sR5K9DCcA8g3nTaKjVq0XzfKzMJzQnWGzkzx
VyJGCYen8t1TbpuHPkXATrYcaqIyMpQiTQU8kzalvKWWM23R4ngh9rVAH0/v8iB/
RZoQZn4l/txAOayA3wd6Ne8ezhX0UpZdN1W/+5uOFpIsVzwD+fAEaU2NKlkrDoYN
9+FZeJjXtxAcnKuHbCHizJ4Y9k0+c5c8IVhiRY6Ov/JNk3c2adIqbhjNa8c4Sli6
ke/qMgA5Ai/KA5EofJj74KDs61caojbP5KbxuHF/vHtbZsFRC8Y3NHHNllnv9XCo
6qHSMIOSaCTLNNQQrrrpDonkuzieK3Npa1NpfXGO5K9tPNp/leY/qsrP2fqgFVFJ
VDDaWisUPdVhx5gnfsw7Z7knie9UiMeWSK0HUUdBJET93HdEedMfZziryhXjcF3E
xZi/mn74Y2+LnDRSKIkxW00jaPqcdrvzjMhvMirSa2s8d7CMQdGLX2OVMQNKnnWs
gRoL3TQRwBvK/XQ8TN8QPCiwnMhVzDpmaE26KdjpNto5ATOimZkl7dda+nWlQza+
+lEpwcCndLKN5ax//mnOir0sR3J4vcgUkux4VkxKCHQvXsiyDRwrqXoOSbQW1ZfA
QqGpDxb1DART4gYmE8cYtBl944DhxvHK2N2dZqIWRpFTITt47keSvl/7mFR/k5QJ
vin4WvpSbMK8S11KloazfGR4Zsn0ywEHQRx6F+3xpSz24A4VHjc0iU2QTgXzEs5Z
PcqadcUCj9Xnmoq0gQB9W9rgWES353UGPeupxrMWtKkIGvVJSJFNB4ZKdJZf+8sV
boguizFzFgfUZazWDMqpPxw+bjjKfsHTmL+h2HXJiUlwABE6aSRkE1OjAK0wTtNw
kUKwQxwfP22JN8zZcv9NSoJk+jW1AxzlpRTyFnoUBHoHqK5kn5EIV6db/dYiZdxG
Mwynp0Rb/ZmXcVAeQtuG/S6oJFb3OKV1Yatf11SHme4ZV7jy2IkqzDmtdTLgUXCc
SJXivDTXO+4xIOaYaRbusrM633rcCocvFVex5kc3Sl2ISB/x713tHcRIbskdM5z5
34sE51cFwV+PxfNrRELA6y6dj5fETURjN8LAK3JIiIdJ7xuyNCVIV7KxVSQ/G/pX
J8DbaKw1pafIgU2zcMQaqz71OUfgeisWIPmeWiNG3o8A5wU4Nlz1s2Yq5UAhP4kL
5W68rZ9Q9c1N6AcOfIM22lKnk1qQpVj5zLfOwy2KJZwm1YvWwSVlvdz0xTAD1A/a
GNAFYQeWy7dNWJry51KLVlRGk2lts7eHDEqzA3ettanPJNjIcIrjv8IBSSBRAK90
31YqgyIs5KqZ1G9rxHw++v7fMwxAGcnBmEpB2S5qFhxKbm7eLPp9pk7A/POvpks5
A57vyAd9/O+MZEPm6SwCGorvUDlVz/7OloHVJPWxFyM0z7PJ90Ax1lkvSe886gYe
sfJXABnrwHcyxgkgA2N6wRXu/jRO69omfXnvhMEvGdLW8wUKa9sRfZ8K8YWUT3QM
ynks7/fF9iKIWxAVJsB/LHLIFanekTSV6ZzmeSeEXx1n963OzpOY4/dEgHaZofCu
P5nh7cB8VcayeiTfvySVkct9L9zZXbm5R9JY5OsuVQ1yTPc+zH4TyzZb/7DJ5U4W
Fp0fLu5k3juG4nBvkU+yudaVu/WToiykn2kjpt4H7q7cY2OD6S4qbDYH3Bc186lJ
OFv7jNhUFZDfNg0MG5cZCYHq3IPN93LqLpfD/UfO2JfLSQ2vWa/xNJGgm3GQhfkK
2z7jIa80DPZF0n9Q83wYcEqvXrIbhvMBM9Sb/LhlbgKKX8xaz4sgpkb3Dc3HaCrB
uMrwB5cFc/nklr7Hpwb/RVFpNS6Q29FfZBp/FF5wlPqSfosRoJ3dYHx9IDhDTR4J
hU2IEK/2B/XByFp0P220vXIBnkz5OadbjS8VQM2bi1jlKKTSEezfBmrHigMZKNLo
3pwGSFwWhTjMXmKQT27WHmSqCeu7HQTxWE/QUITF/uqQCD6sjDCEBSF4ZjoqnoqN
tz7R/NdOvAsddqZuKzqxqhmF+kCbduKJ+SvJS0F9EIB16kg8KV5xZVg6W/vw9r6L
`protect END_PROTECTED
