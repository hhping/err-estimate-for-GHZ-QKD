`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riERj75uc/5ZBy5xOCMzfVLUqcNvvFY+vPn1rjBEmHp7Wdl8T24cv0xC1981g4Wo
eVERDvJrpkJ3OxIhP7X8kwTuKn9W+LtmXKbpXKb22jF+rJdK33g0pS6LaKCdqTxY
hIHz85pHH3R9cgl/WlF9jMTvrMtotLV5HvfRKqR836SS0SEi8F1IKnK+b+3JdFAW
ULivnpNtetbPF2evbpCfCPgpVo1R+eoMWTfYPsvoiByRgWZZjRWJb/AXpBqtSk7h
7aXDM3qUelTk1LPSKtPx/cp9/AOsvXevwCmuaRZBvp3gjqn6mAXD/vPyVpK9ISDT
BcTvnrYkmkZdX6HbGphzt4vF/aFeQ/wKzrdrSen4dWhAkURej6hrOIbpOVeR2W3A
hkC2pnmu7LFWY54aE2Qq7VabnpNghA4UoQOzvIuJlHfLiCCwBF3ImKKAS5rN6GrS
vhDc+bA2wgDY42BnoFFhPe+HDZxbDq5E9BlBakmi43VhMoc6tabZDcKjsqQxB75Z
7bmmVfg9h0moQWM6RtnRaS8iMYLhKKiSNTCnn3rLZHV9VrzGPIQcTXfegMZikH1/
goR4hnpHtvxtaIBojCM90OktZ7RhfEk7Qa8Lf/NDfC9HCJiv6ccdnCSndB0D8AqQ
iF20pAx5UxzV27Qp+FVe/26onI5EyaNrVr/QEJ8xu1sL7J6zmX63DfyxlUbt7RGz
OWuXnsNdxmkT9vsY58juYB7sEAKzTUWqYDlDCC+yMzHYbjC3kj0SAMsTOeXDTcXw
raLmdZX9erpwWPrRI1nuiulIPZLzyZlVq2qV5xct3NzZ+uUbIIjjMcEKZimEhypL
C4cnyhfhwKOVFMZF5byIBvvJLKLOm1zwnQkpm38V4eLxidsrCdLplVyczMRYbtgR
W8OTW+Yx/D2IOWinG2iCZmAB8BVmY7TRzZcxzN4ft3qX7cecDFoHCchS4s53oZjF
dToV1Hefix61IA77OwNR8ceJaBfSOnIfo5cRLiL5XlvHJQWerJfqpebgUc1cToA7
bG6mFAdtj2x9PoeDGJj76CHaCcEmm7sUKor2K2T1hTVdvksLHx15fGn3thLQhYRz
jOS1UfB+hNvofGzTjNq82WyrDvMSPxPX/Fsyk0XkAygTpVs4+2dT23pxi3rmqvaZ
xRJpMnKFSVsJW9kzFGDvGjj1iHphmSCxq59iT4TOL0h8vfkQqWQCii2559M9ud3S
KnaMMVf27nT6/gewiN7spjj8j+3AX5HCoMJdtNYms3ySTwHKWXgLx6NROTR8SnOF
S0Ub3MujFToPrVRuLN5+vmx7NSELUIlKEMMYLmh7SPNpzMwa+L2cqtxcVU/6ctRE
`protect END_PROTECTED
