`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7yoF0SFc6sGKUUDVcx3YtDHPGNxv9FgIbONAN8D/U2kGJM2tVe8/wa+C8SxoL3m
U0IqCdIPS58oFUN1fSZDbWgl2NDe452A/6ChkOgZ32HGJTMY+k/xMefuArq3x6/s
mL6VTAB7Z8f4jvlk8KzJ42P0MRroKCiDqG1oIoJuTSZAMJ/o+4mhReBHX/+zKQe0
aJvBJb4K7asx4TQEnHRJwUe3EO/pGFWMhfg6DyEOBiLaCVhz3puZL9529LEL8my0
Bp4golIvebVYNNdg46lWFQdsxoyhS2dVGZolAEDXMYGfT6LiMasE2f6+IhWXyfxe
6sxTS7ymn7wPldyN79PvzDULI7BD8K7q+lkFUEatjOwSMC/JOgFjeUN3xiuzMXnz
EUj+aP23O8lxsTs1qeUhDA4lX0VGota/M3V/tP8OIjdYIcAaw7m9NbqzDJ2MjFbR
I1JbaAQxG9Uai3ctcMWrmIaRH/ZN63QGRflK1ag8N26AuH3b/lbxsWlJjK4Bdpje
b+0H7OjlHDJrq6/EbCnX/sA0pqO9AVVwvT9+2vHP+ImVyCRC7XVckqj1KB0I2kS1
7OZr4HHH7BhgYO7SzL9/G6lw6kMEfvYZYdPBQFkloK4DYrSvpEFle/tptxE9J56n
Jxt8KGURE2J86SEKTW1eyCOU/tl0W2ftVi95vfecLeJVUyegB/iORAN37649w2PG
lw5zCyvEdVKVadYC3vCaPAQYfLpe67WRKtZkcR/JXqFQvOW124O4zEDW7M8beseE
YPo3kIPkcPdZ/8G50s0jBcqVaH0G7wdDid0+A5qydZX9zmRW/7fbykiZqvA37FmN
1LqKG4ttQ7Zti0PNaFnkhxZNs94tusRb9zZojQd57p2KX99E+W/3joAKneNtE0II
OD0UezrwsnJbyOxVQpT5KufihMRLCTqJozIPnv7ZxFPx5PdKrI1kflJo5w3Tnqkn
`protect END_PROTECTED
