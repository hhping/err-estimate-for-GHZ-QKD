`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zv8/ttWGDg6rYbqCzR8ToSw47eCHQpuMYOIgIvlHTe0pjIghaZWO0HWgLY4YF1KS
CXecLDJn//oJRzoMehCg3lcHevPata9eOE3SwvEqomzClGPxa1iBIG901/Y2UvXD
Hh6N1DO1bJLegpyW99yUU6uzcfTXcKs7Rzob8SDClm2kCdelaUBhplThEbhJ5JGg
fBQjBfmHhWumdinlEoztRPtwXMmqPjhpc2eEDc3QX1ttmFQJ69dZDl0ipcNEuBkO
KAqzrJh7rgJ7IdkanHxCJoMhIHUrsBo/GNJorhUdtkZrU9t7tgYtJe2ZE+M5AMRY
/O7LSPoCPnFXXomV7mnCjubxPyyI7D+V16lBlROGdHsV8rZ0P5diXMIoGT/8mp0s
00e1ZYbmFdI/ZjZmu0Zqey3O/EFdAPBMUBfD3dZhzVSItaAliH3CgJL13fxHwkgV
eEpEZTaMbnSE5UVos5lojbmvzhzJznoACB4CiAR/PGbUeworwGVhKRt6UC0rqMHY
QrM+nIE0LN/BDP+dZsmDqSJuovsdXq5+LMLyArWNWwxb4B4eO1hQjsC/rtae93da
802frjmBvyPqZ/JA92x8qUPwg1t5kbM2u/32iWja6TS0Ehl3xR2olJVLVHUbaNWt
QGdCtMRiJg8qZLdKEGrvQeX9zKv4PFjUc59DYfNjUWJTBJkRAuVueSq8i0NcWGL9
Sp04nCGdLMPNIXazcqFDm6O94J7ssSaIMQrIFxrXhMFDHg6SFpmOzBtHG80SLr+a
0tF9FiWrqmK2yYctrd5cYL7W8V8bVYE0+QMx5JI4PB2NgWqPk2oBOWutPtjbFIbE
`protect END_PROTECTED
