`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqAI60VxuuUZ64RyAXEulqC9KJyJXrbSlCw6Z1kbIeOsH+dhv7Y+3bLPNdW6wBtR
FOM4Y4S5R4WxZgE41eA9rpW0S5cAXzl1IRK6eVpPuQaNP7oIVbn8sBCHEXVCKro2
XyeNZqJzeNlwzPQMWe3bjgEqaNaEk8CaC/8+IgyM2lDM6JKzNrXT6IKSMIfCaURA
TV+4ibF4TCYLQc2jys/fJYQgIbR+vR3A9AaXnks7QzhBkN+M8xwfq4fsYeMw6Ksv
JwelZdwCIrxniJpMgSXNLIBt3MQ40GR1sM01TC7GZ9ORnZ/Bhtnorid4xfCldLU8
R0jXv2wQ4J3YmkuihiIAsfy9Mg1WCnbjFJEnWqD0PU2pSrFNUsughrFiVgiP3fja
BQrUO21kLJHy2+uLRPku+sjExA8uH7p6jO15HaQ/0gZRj2IzuJb49UBB5efc7ux+
7Jnywuo5Gq7fazxXgorhaL+WoAlKT4ZLnrhuI+VZ6Pve/lSKlKRzAkhifrXEQFMc
CHKGcPblF1ArooBPXn332NyyuOZ4BJDAcm0KBoJeh8noFDfEubhxH9tctWiNwX0G
I+mep/2Q5F9OEpmrFg7I7fthDOry3STQqQv5gFKH00+Uuntou8a2ozTfetvns73U
Puz76yWO/X4ErmfLHnNAaYXhttqsuVIwFk66KeYUGO7PJhk/Dlt/5SDWh1OFQqwM
`protect END_PROTECTED
