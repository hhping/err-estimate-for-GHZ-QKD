`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeeOuftLSDSTr8AuYbG2Ph0egpTyBqNMhvG6v1vt8DXRseSTFLI0Sycmalhm9GAL
sr1U/YWSx3xoa7G0rZZmE0Kq62tsE4V8e73v36S0u0HI+5LZtulVdelen1flbj5r
DU6/nNtTpz658Llnnb3sE7jpMIM2OQBs/F9U+kjGOh8vdJFs5mg1LPiqrHc0dlq9
3joKXouc6WKyTnnussJ8DFria71jeROBYDBTr8EGkkDKMmSl+celCp7faTdTBhIB
kyHwkTlBL2666jzeizRotoEto1oNDWqAyxWw6yq/qw+kdqZCG7I0l5QJS96h4IIo
XJvvmAeHob2U25V6L1f4uthN1OS+hWUnkmu6HjJ5fseVI+7XlBpaGNjjsGssrbk2
mA6zgaNUZYG9a5x6FUgSX7+bbMwMoDrXw2KQXIMVFVxwMtUCkhFLJP7g6yuyPZMF
xFIPIFn1t1jT2LznEJEWKxwxhz3F4deQb5z/Cf4cRzqtZwARvh1YK+xShOvcOfiy
u3j/DticWTchr8iDv77VDjkW7E3qafcVkvmg9J+QJw3gEhHc0oGbDPtbl2/jH78S
CZXOot8BK135lvXdm2tflqoNrwPwZHr0CVTUWhQbPnHAJoVaE6xtWrOVK77vN6lV
R0VTibM/CpidhjXdmjm5my3eQXKlwvZl2XVhDBirTa0KY/Vnux+3Kcn6DF6txx6y
TZDES/x/jacZbQqBkq0/T0UPGk1gIGpq2BlMcKXSItLMqW5N1UpfyD5Q9KMwn/dV
Y3YI2lznAQCmLzNU1JVVXOoX+fBv7hiX5XQpim+v88PGNo4D8+/D73VYomybhTV7
ODkb0wif4/Roi8sCI7jOvd0aDBvxE2bwuYaTCCE3XDXZCK+Jg6bw05k6WFTm/z16
ZlYixe+dW6behuqiquU4XiyqLEuN6oxgyRT2gxl5uL0QHuRCMlD5OKR1lBpx3sGO
8vpp54sbUHu2Z7DR83L7Q9jynu0HK2wWo6Qpk/Yh0BXuZhJG3NxAHJ0JKMrznfCZ
vR+3PFt86fAp30/+ksjjr/aPfHv2oz25zc1W5rCFwOg6jBrS2GZyPCzmOc3ZV/tl
f7leVY3AnNwxtud3sVWH4zDU4E+UTVu8s1YLAkr5gf5AoX5Pr0YE0ss4KtnHE0n9
y/ee3kewDUydLMtIrwCWI93aQ+TWDmeThSwwgHwGg85Yq0om/z2cf+SF/bTflKLH
WxtP2xcgXGnKa3OTYl7YA0uqkQee/O7WL4fjwmWKvk918yqR83GobTONuCr3KPQ3
6s8a4IPsf41UVMLuqMkdONkkofHeNABejJ9gXcqur2AGY1ga7XyX+R1mptd6G9AA
LDPFmSmq2lNF01dq9Vf2MtWIQFU+7dzIiZg9QPbccdwlr7Wt8DBxG2X5i1I1wf0w
4MGeXCrmPdkoFpKNvb4eqnxtNKLbJe47NAQyTHNSTrRKgjkNDBE4tMIiMPaK+rgz
wQzTW/ljFcTSHAFtHTMopVEPRbiRByEu0lTsXXqvu0LxtajuU7A8+2XILtR76vlP
/Bg0wpVSaF+IcbvfhtLBIWZDgxM+lGWx7lqG/HpZOZ/ESNUC1T4zVm6v6h7FNGQh
DcylTqaMBX4BvLwCR6aIzl9WFBZ025nsVVzUD4LNuojFzC78L86vwk0VMcM240WY
siZ9QyGmpPyoBYYBOXxBM+AgYERbwdEWKCcciR/YLgJaaMXePd1EnSqNwuilhE21
iYjegIG7mS3Jf2r2s7BmvrCh8PQ9plgGj614O4FXYAlEWXZjTtpbB6+ZDchHm7sZ
Sy5hIeX+t14d5DjOvNJqp95ams5WmM5N9a4qI6wu/Ud53pSkc07uVnsecRrsxfFV
wXFHQOEStyYNzNHgkZkzt7uGNiy0Hi3hmKgyy9t5gp/G19plEM3cMDffcnkTGuWI
M/8/FmRr+ccNCv5shaqw1EUqXVbmIP4nq+D77YAjq/MzPL0XVddTvCePiJYDTuoE
ITGLYM9klSYTQZGQmwgd6NalC3Xr8xmmg+sTtHAZr3oeXEZ44OACf/hafqgV5xQd
XmqqnoLDevIFLus56Oi43oCrDB47ALtw3H1sDdzgy+AYu1WNWOP8Qjvh5UCg0sz2
G/yo1hbixzNQXTUwuhL7EmZevBIlt05i0zAs1uX27EI9Y1crzmnqgaNbdMf/A3tS
db42nVhylejgdS/BkNPdgUYkZ9aaS30dCWvxHew7w7kHUGydFRA48A7LJ7j8Zi0u
dQVFGssYgFMCix6W/C2YTkpSEWPRTgUJFU9zvGEvojC854DpA/29Af3uLl2KRRyf
7AHUdNarjHMWjbTIS5Sy1CPGzd1hxr29vhM9cPV/Pbjl2vW1rTn3TyYZWPOY9843
WzxUTzDY96uv+7HG7nBMsjRLKvnnBvU39xyRz7yyyxTnej7ZJ/Q0EZgPtO0ATZVJ
Yaxr5bLxS6K/YlWbCISliuxEZkdxFkb48UWoHX3zucVVo0cUwf5vNby7kv4TlpSV
257HzTiKpuv2hL3ijtY7gOt/xJxz6UUWkel2z99UTB2JaLY+r6KQCgjpBvAsxv1+
5Ks2OWhdakr8I7x7VcxdtLD2MBZpMx09ck1e33lV0B8+wj/vCbRAZNBtry7mrktd
ALxD09a3TmeEZQ8BsNTLnCLveTof3aqUXNB26lYYkVyUc5a7Jtvi8pnhVvoYi4gk
tktCXJaFGZXJ+lD4B5w+Z53cDDjOGJCryB3NFL1utZV7rzaPoZ+MG2RWlYtXn1Hw
UWtRhbNgxQ21Q44GiNeTGgU25JFLmUkCw2cjS/4+eRLEKx5qxB20cQ1iri0SsiLi
lw3kcLgoj3nBIQ+qcoCYuyXPrBk4/K8wkmssCYuzETgWja79eqzeqc0+21RunM+w
VljWkv+dugJEcBtX0Jbg2n/1q8ojtXFWzmyiXviwC/FHGpgEW8iiyRipvrnUxFim
cl8U89yckS8zCoRu/CM2P2YGKDGgklAZ4l4pD04x+3efBMYrJh+VcGBEId6J2PVO
8NugfBWt0DWv2RHA+js4Y1am+UtEMMKy3oFF2wmQB/q8QH3KHyMisVvheg9kHRsL
Ffti/TV52DZm9W878x95MCHLDlE4TfMtXpaJdoJdzctO4nrE+wOSjO6HU/ohJJo3
65wba81qWpG/fMtQTHv7jNGavmg/ZKljdCLtkZgjycg9JGo/9dS+qX/8dUtUCEyb
gtCvIDxa6pDz2wZUB3Ytf31L2BwKKm2PRT9VA2+vEQKRc9C7/EGEMMU/PC3RjIq5
`protect END_PROTECTED
