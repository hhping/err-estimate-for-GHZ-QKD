`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1xEJCw8Bk17hkPLaeSciH0Qb4MifPPvOvvXq/G/x2NIF8I7RzRRGtjL502wbID0
1JYbzbsxPSWOqw7icpPZ7k6i9YuE3wVpH7swZ3bXWRdd1KTo53B4oWv2psFcAMNp
MTXXnRfHh6FFuuiNyD3HOe5LIekQr1llyenvC4MTTxiPDO+ZxewE3FSafqumlnZn
K7QLN2Nygc+O13WGmLGfsf2bGepcg9yRI68XSSU4p1efipk7iJ+pYOnivliZFk63
Pktw0joDYKopJIeyYAMA1I/a8RFsAQE6TSi5AsFHCdSQq+xXrCnSvcnOBfKyYVIB
xaJypGss63OrJ9uY2Z17MOlRtxKpUD95P64K9iW0ae3sWABxVPOl2DkY0e1SYOPc
rKAdfEACKFy6A5nq5/RU75UroLz4/88oV+uyIVY2bEoKJjAgaYXYtmZDC2ItpqF8
BEPrjox0Py45scZbbmiKOdfhR0x+7pf0lsl/m5r2p86ygSzGbPeY21M/DhCZ7Ocu
60VrjlU4SZs8gKD5gaNhHVVhX9SO3wnCKdjIY6lYYFQ5mZxCdWiImZSoc0iZ2t3N
6teAYojRjjPSZ22XtZze+0I/8IfhGYfDat9uNvl1YngWIGkN3oTwNTPDAnnyvlcu
zpatsydGTTrMQNdAoDlhw8UhPVRbw5cGIKhs5jotyCE=
`protect END_PROTECTED
