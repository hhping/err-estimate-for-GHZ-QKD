`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGDVjtqlH3wM7KR51emvpWf2Xxh7evIENVSDw4KTkhbiZCiNf10yWbeNTlKAUFaf
PcdZ9pk/2LR+Go86evpp6wKgfFigkMEBN5aOEAOUvaaKZ03juD0lV+DpoqkLTatZ
2ofTgeT7NoIwJ7ckFowr5ye1Rn11CSH4DG0b2q2UT7aJYisbOZ4iMBb1P1IRf8To
INnVL4ftWprlQEH2grz44b8fRyl6IXlyGVPvMiSKNWHmSGaOEHmlW0Y6T2GnRNnf
/+ufLHf97GPQ+YgmtrIkjOoDmxuAvUCtLVZoOnkE3D9A0ViC4nPHYhn+6jCGynZn
cQcjv6e5GiOQgWbkehw8jBSTKmqhvB+nB0KksCB7D3Z4HwPzujz2Z/hFnUsZTNYi
MS2XC7B0NNmOBNKwqWXv3W00uiF3EGxeJQW08NWeXXl6vg7yfvJC1YgXDhSakl8B
rk2JE9xYyFXfrQM1sDgEGv7V+9vSKMFeVg4IvpsazTajb45LXx1cOjXUJ8Ff7ODu
z9f8IQnBqEium3eE+dqgBWE79jSzW4a6NZaBwnQrrPZUU8fXFQnVNeRE0PI2DEnq
qBwfMVcoPrfWulXHkXjA+9WH5Py2zmAn0mYx3t0odROyaGAElMnyieLz2S2KoPJ/
wAaxmxQ0gbJcnqOUMwMClfZ8zBtOAH+CVMFoImTNVAdKcdutanuUTtqPErHHQO8n
vDIkvP0tGjhKEu49HW1eqXFYNA3JMTn9E+W1ESAgmtyQn594GI7ubyGt8YnqcBby
k6Fi7KvLLPWDm52wn51C1esN3fcuZ+0DeWOenvelDBpGSvjn0gZIKxL0mSYKuZOh
sABv3gnMSrH9t+yVu4/ad/dS7y3TkizKn7Oz0M3II9suZEJXoMrkrdq0SaYQpG1N
4z6ctwFsERU9qLEWgREgXkqh6RCZB4jRk35KjjY9PcTs7z888+ADYRdZMvDVZji4
SvJI9x2RfiOHVwvr3cXwaUw67vXB41aqPghXni0SQDS64j4IR7GMBUR2qHgPaW+C
OTkgkiEEJ+UbFMMA1v5IgFb2WaBgJdV+mVDvzUsAFM3+/UsqDwJFkVUyW9dSTm+9
NPNfjUj6Z+QFqj7IRVoYFJ5tEuV4Eb3KT51RbTzYB6YIDj5NYXB+OS6Aaihm1OFQ
5x6TuOHPENV1q02nr6JTTKYugyc86wonP8dl8VI7pmij8v7CSZW131eqHT/54Bb+
doe6P/U7f5kA/ARP3qQ7nnlOzd4bK4bgwI8w7++4AtXSYskqQslszuA4dIn/VEUi
p4NfRpZOaI5Ps9EshOIk0syZbZMYfBGaV6+TUw72Yo/p6JsDyeIW70zWloKxpVdv
CwgbBYPy1Jzmg0oGox6y47Ly3Wp+kuSZHci3QAlmJPhAtTGKFlbB4ISjA79xXcY0
zzH3rImo/mKQBbZukuIk8UxO63N6vTTxt3bQyG1y2V6cJelfPdEPhQk3qTOLbRgu
5xAYYagu04RDxmEgoVAMMd9JDHlsxWMOdWjiTbfpEwcpHtlyH+IBIjZUXQjlp05z
6GeFnrvkfdYTKetZxFmQLDwJZzeJXUe2SgVP2+zxViFs6vu+cgyYNdfnCOw8o2Ev
nzL3jpHiGO3Jwl8lp1x1d2uGq31+HjU4UG5/8On+VBG4dOUPWp+SYQ0Vq6PdJg+u
`protect END_PROTECTED
