`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l3C7mhPEymwA2pLNx/7sqFzeL/oRfvyKJia0/yqbwzreWen0hSReflXNrK9zGN57
PFPTjRd9fXj7YpbaF1igWFEu1eZHH46uzHwp97rXg4pTNjgjt6zGCI8f6n7K9+Wp
30C2xlp2LwUzeYT/y5ZWwWZK9k8+8PXRTZAhAoNgJxKyC/I7JAC+akKgXD6nxUe/
yF327imerzdBR25xJvcWeynZN3K3Fk3x2cdTEGLCPSATA+YKi8XPzdhm+MqEugMJ
si6MGJ+mCy+1mVFySz5LjHjiXwAhBqhAuwrbllnGSzE7zb4qsr6GGkCQQLuc6223
TEsrUbiduWKoBG/vGyUl1tvWUu1+alDNNeL38AzEsx/Q5j/tCOOeYKdMMXcwuOEP
qMajVEW/2eZsO+MuhOt8F6pbuFJMem7/r5pVYp62e6HXksJU7ssS5PdcH4fMFvZ8
pNSN3Kx7kri38qRNoholNEqah0kgggHboEATkUH1Sfm+QKqBgr+yU7WJKn6XDOnk
9Nz3PbyQyN1PcqotasAyNecKzslS/ZBUUNd7BWCcLIWMV21XPkeKmp2hrew1WnFs
RKHJ3YCNmtK5+paQcQtuD3+t4r3P6dLJkbatRjryHi8Gk9xxE1pOnaPm0F4dJgsB
5lCxBTNkhq5/qq1bb9ZlsDztx/Mx4SkpDP9HGkUr5HxPQOjBtNL+zNE0xYbSKour
pMQ5j0YlvPTpT5HONYnSAy0le54I6nuLt8iC+N8XxhJTiMVzkpCm4KzPHRAno4o5
b+IsO67w7cQAVIXXTd+Oa4lBzXL+D6fGIWQEakyt7frjzC37wx9H46ExcLFYOQHR
uU+LeKTCKAHzNEcE8zEFVPGUY74SZ+JLOaDzYNqaI/aomiSraK63/iu2hCS8Adxy
CF3X/TvY5iDkqJcSPnHkJWOBa7QRr1N4lYftI4IVDRu6oZ1nutl0fyUUpN5e4llb
dkWYXw+/JnC6tThFBtCP/NfH2oqrd5kKp/1VWg/ofHejmJEMeLHz1w8sgd5zwCH+
g0ZmIx+zPTuT9lRQmm+RlHhT2T6WpJn8bboLT8rbrXbqwApF0dwOHW5hqL5HiG9f
olp+RmajHYv9jG7njF9rHVTqNkuvPAt/sJkSLdPRgMLkytDivcHy9NspTBs7vD5o
I9kczK19knmI3LtZl7hCwA9bQVVVKXZqk6/z2PPsjeSG9kUiiSMyQa+X07Cw7uWk
1sT9oKxQvrK7EOKE3qsqmWop8IyOfl+xczMA8yb9bmACdWh51eJW2z04CjnLaAei
G7hwox7XU41oKdOjG4UspWN9TnuhNQ0M2QICl80lfuzImao7Xk/JSrFPdvlrfb07
cnQzMlHb3yo944AmqOsXAmV1FZKXbOPHFFDaWFN30yt5Il39bfWf0NCylwPYiU9N
qxcKbwsaSPiZYIc5AZ1E18zmkKpuAhIAeJDz+H/5uvcahQ4uoPb+fPufq6D83sPo
UI/vSIkbo6wl9oVR0zUEjdPla/3fpJl5B4VTM27b8cQM8cp8F4re4pZwgIsFXaaE
SwBjROmV1k0vhzXW5HQrVLlYT2iP//wrOosGg0M1yE3SVrx8TsAmI4C1WJlgrIy7
9ASa0O1SEFDsDTdahAhhZgK4JguGcYnQewuP8ye0j0iCVQhxpOBlNbLqOJZLpREH
gsFRjvRcG9QudZwZsfSGY701rgExyqWKH+VYy4v95bkdfL0ETAoGk5RhJ42m3dFG
J5q6j7mV3Yoh/I8j6dJnCQlfmIogbqyhVkw6ICxhAupIFte2Af4L048mlVrr16M0
p9dQ9ieaZ9eWBOoD3XEDIZ1Pcu98IEEJ79yxmpJqaqdJygwl3E6xqBgk1kew+Yu3
hAEhR3xCn7jxRECLUK2gzM7HygIoG3bXXQ/XlvC6Gkwq4JCyuyiQQqb5xs8xm7Qq
+EG/1uaqbe7I9DZjhkYJZY7J6BYds7rucQahjYBJ+1SCw06VHOuw+Yt07AFKQ8cD
iu8Wv93oL/M5cwCoOBqiXkHhmPoneq6YSqrymz3ywDkjvmSHZ9IoLJ4OEAGNvS17
ZHfq79yiL+rQmpl/9GlubyZ+DxGtGMqwmCXZ4B2GyEYZ1NBQ/pvDG6uqIi7Ezq2s
i6hQfW+nx1ul2N2sfIKN6eSSeZjdJMkeRLOFdXMbQq29x8qDAY3AkkTVKzAK6GRY
GHzKI6ZXmXZmSm3dcIZmqyAGmHlyVFVkgS+mHGE+mUcT5PSIcYy2Ua7+bqcGHpkN
rsjkVEOSr7oWkaeMpZFooqIB24TbPCvXP4XyfNTH3Iq26HTWURwTTLVrAlMcBQXq
6fEobIDj99DYEFpwsJZq3VgzAklQPsUBFjNNIOQ/vzrR37ityFJ+3QqEgYSRIBHz
D9uWthh5di3PIkOKf+AvAKUQKMyDCcRuXVzKxf50dTwsGkzVPQgTJT+Ga8R4afud
7jICRW1GBiWbcaJqULgbNeLw0kt/qgckO0yB+apWjeo7zSSMiCeAjTMfRYnFQu6w
kv42fk8AIXR4TbyGOZ0A/jhYvUHZSZPoGGHe7HFhcR3J8ClgZcQXIIXxGunFXulT
S70clODIXOat6rjRso0xdsFbMPefjtv8m2G8AzYTGdJk2IbH9psr9wHaA7WyWMRw
JaH6OW1Rhrns66Stfsmv35CeCa/+0z9O11m6wPJzzLGwqtVorUtn8L8ZTxoRS+Ac
NbNBTY4x5Xo3GHaTj96lzHn2tbig37f3zqm0sjBHAzQjPNC7qio5AIbFhipM2R1I
a8V7DSuj0ZGLqljoUa0EQnNO+CQKnY0GJi4QoL07IKqk6WAJuyznP4hfEIxXWemu
dnU+IFzTiCcvzKm6GBUHU0mgZjz+zHk3FARowSn/iW4LS2/xpH7VprWFKYbdkKK1
yvjvju/cEe8aPFlAXWF1687dXpILFVATGbWSrQPoBSJfKdcoSc3FfWgPV1fuGMRx
5GGVMBOeI2V0TR5My8Q7WD/dP5/OXvXU3rc6tC/XW5XQ7L1tjkpyZGLibeuBFut2
Z5lZex04A9XS2UUEwoQo53boweJl7+jW0iDtWTgWlnlzU+kD6d4GZzRfj+HgX5py
QjkMKi4plV33bhl2h9LgMOfFRTt2960clV4SAy2QDFih147fZhfsBHXkj7qsZJj/
ZFhnN2ez+yAjlxnyDdonb6/DnA+OCEuV1GTDqABxj5BRRMrUn5oWdxTia4QnVxhq
m/f+inxfodhqnYElW1UHrpTMlIt7z0xEXo66EDlwgvyXyiDYbL0PtqigQYxcbj9e
s15vlNrWDOuUkGv43QGa7gzD8i4mWxQHte7EeF0rBOq9eFrGtVnSWW9QK7cm6Z23
TepCETpTFOwYFr2uh79h2GcaCe21P6isebbCRM+ajGrOpdfDJSAVlISIPFW5C6LC
0TVcKEYyxM7Hco699aXgs4/dQ8Yo/Qt9MUM5X4Cybs3eyq/BbXuUEXab7YD+UjHc
rq2Kx1VtVwudxrrejgZW5bZNWOmx7Li+x+UBg7f7AuYtcEfZO8hoJQYLEFaav04g
zbSUW0DpX6Myw0bWmy0KWJReBlw6ccjmx03Ut27DGCiYS55oCZ3Q+ltuyGUiTHbU
vlpxd3e0fnGMCZS+dX2p8AlNd2KBjeMndmjZ6NLYVTcX9e6G7+eR6PjRXn3fhZSq
WKiW79iZr8fzWlHGdfYYKwVmnenoCa969hYmY5XerlGJfkWDJfDhPUis5nS/j0I4
26RxsTon/FAO4B/BhAS0ReJ66fvHgIjz1V6b38al2iYemmRLhjwCsZfRzeRu5wxs
zH7xayhS3FcRkoSp630KKNZ7rhKOG8XOOmHLnF9acoJtaxT05QzPb9DhJseBQ+n/
Sx5dCpLWQXuM+WbMDSSeRr8bIv9cT7ia8Spz+T4F1QKLQYlRR3PdO0KN1/PUl7K3
Yz0rJ+XvwgPCt4tu+ESRxR76j5dWueZmJKRHQCPxuJnfTCA1xntHF09BXVBqud9H
BbgrdK8/13P9GX+mPIB0/EZ9Ss0j8UY7pE007CG94NiisWN+IpKTKNwBrkFQIINZ
JHpqkT+SUO6HBJSv6H1YOSNieu+9YKxZ6fcI7tBi5ae3oXv9DLYeYMPMYjRG0fFQ
8OV6CC6sJ7fQcR7nodEemfhA8//4KAjAUWxWOUx5qMPjSNNrSIhtM457DBlnYj73
zjMqayVYNh70gdGpOrsQpaGKtu/z4tIbK3U4DoSWl8JUGADrWin0snQ/L19lP4nH
RrRbxApPggu+C1GCLUE3XNmRHFG2OkFbXIhbavNX15Wxa75NLp582m9AgWXUVUSW
ktkhHCrl94lv+0qVpskMb6oLD5sUmn0EqSsaMJK6GmBcFsw4+4PLq0u8mvTM537G
6fGlVZr+VaqyQ9A1XRDB/ndywpyHSL9CxQsjNotz+ceFStOl/MlV/WODjydneFrl
wCt4B1vAyshzR/QNXICcGnynkGF8Retap4zBy32mSzIpcdHmhPUtQqK5Dfsa+nLD
lDGGmFU2bbsnkTfoFq7z9xT4ZgPgrJ0ShkMzEQJTieDJu1XPwbvoI1UdYHPl2Dcc
sgiCwcWH6HTH005lOJ/KGN4HJ6ZKXACwiPNsu1h75ejVGKSFBrsZsGyM97wj0uID
HfoxiFWmMlr8te0WFCewPO5yPm0co+oIfxqUsphNlCKz/SbeRy74ZQ1j00KLUQ0C
/2AVVQoY8APxhH9lN6IBTJVFX3tqK6w8Zv4a+IQLAasOauxJix/rF1WcDskzRXnU
FK0YSJsskY6+ATi1vBMKVCTqOLnX1+Eh2b+yAk/BurUJfUvHH6SYlOAVR4W7Ars6
i3XWSiuvOvrxs9FeiAmzunYj/hxDjoX3vB5wXCvDc/o9/YBRvgzzWDO3uLwyRlnc
Qxn7X9v0dYJpX2Pof6PV29dxP0xUufu/tLq0oRbJs3cqQrhXqfz9EXNG8RXNZF00
jwkgAiuUbyiyKKj739GvBxMm9daCmJcYYYJhTH2DyiUWQJi40SBjphv+EFUdyv76
RRYY9kzxRbCpZeghdKU1Sd418ZSzp0zCuQc37UfUXtHRH2/kO7JdVK4CiKAY/d0S
YgtGyeDfk1V6m0uLDJp4eVBn7YIB6EmNdyMDeNSiDyfjBYOooMH2SErfXUgqxP+H
cym/HXrNnBkcD6vtemxLUzwbEovjcKiD+YbiAkm47t+RYtjX9w6Xcd/vslGNsYsF
yYkw3Fc61Hz/AgJAz20Ppk+dtbDgBKifgvEUKaIgguK/ovHBA+NOHQ1wudibalFC
NsU3dLH+S+FE8bLH6HOe6JPs/u7XMkOUxwAlRL+q0JwDHSt/Sb1O8IJ4T691bgOJ
07cU0L8HDwNJfbohCULnalfshUixQJ/r+eCKu6RJgUr1nE5BiY5bYWUUlr8W3d9C
qltSwLImNnoDX7i6YdZhqQjenWkLmsM8BSv/X01DnSshGUFN0GAwmUCGY4Pm4M6m
Wr4Y2B0LokFmXqOvzgy+r2amDV5GioQtXAO7JhrSXNRz42bLdzxzWxpsYYObX2Jx
TSbKgu9Q/APdMLoqacyGkx8V2nweGRgUlYGwMM3qHS5fXkkV6IwNKXbt1WNci8EC
AYjyL2+selhQP8dnt7wTc9fql2FfvnmdQk0uTN6aXXDL7/FJ/1yk6YyE8kRaHpUf
O+cM41Io4VFsBMMGCS0RuaPSgvIrgOXNckgkYShyAWsYC64pVRn0cDdCKIJwZ6e0
LApEC38gGlMN9uwqGMPGxC2DG9MbKpxom6h1sDk3Wg7/dj9v3vNKe3pw80pCDLsO
oH9dnUy/IGOCzmbRJ5yIeZ5Tbx+v6cN5j1KUjTWQPj2TG3aiNIRfjrbOH1P1XTYp
SkZHN5i3pmHRl5PZAw8XR1iZ8aTKOSZOXYbLwar74C8epSvBW1Huyb1TdMS07nQp
RlRJy858NQRA1ZLqMQfDnv3/QMGfAG0WZUyGeKW4MguVtMjq9vGk9KHnvrVR+tAB
1X2rWnmWYLgGGrVRzasYaUv5pSifHjtbpIZIQ8bUS/1piUOMZfl3hZcpkW25bPB/
ZpQcPr8yTFZOn8LXAn7B/zeuibJ2j2aXwSAf87R5awk/lW1cXLRSjXBGsscMSmj4
RSEAjyk77NFqX8zgHz1EuA7JpHGN0NElcnF+xocvPVUhA4E2UDDySpTN5ddvLpnu
5x5pNzPP2FdkTDRPCkoBd585QkBt9YqhAS5VACX4/e0uUeeh48hKvC5CKBdqsUPE
YVqoisG9V87PUhHIJ186kNWhA7KXA0XsgGchD0hpQlhM+1SyZJfQOAe0ED6/OvRQ
5n21A51RUF4dIdwUAXK/nRvY30Z95RklT7jJ5MZsE3IRgqBfnwMekLG6YgDDycjJ
unaNqHV3a0WS9e4ht1xbChFoufTxiFpEws2guaff2LU4Sgzh9g+pXGLUaA5bFsQS
hmoG9XsNjHsEuG2UduWI2m98ynXHiaSAF7nxLPGibjiHCjzw3+e+MDUJiV3gwVNf
7tPRQ0AQl6H9mewFJ2g+1tHtgQoQsv4zYHwnR2ALGUf80zpsm0WzvlgyrqRhLlaF
QPCfJQN/gIyTjoDfiLdvNgdeNWtaYKubJAPmQ1Dg+ck3O++XGIMalKPFs+9IlCu4
u0ckdV5h8wAIHEyGzdsz4gXuRkk5LVyLDEC4/R/Wumc1bdrnvG0EUBDnuIEJbyha
Z9qGLtPKAFbaRmNq0eOWycRL6eh4DlIe6zYPxnveHaMkXO2RO7pFFhFm7wmRtMyx
HBWZqJSkPuZ5MDdQ/JyZLQt+NvjlDK2Py52zQPoswByqYogOViQwloE726l0AWCe
M3AE423eurKDPwf580f9C+BwOw25JzzObFArRT4kInQbYy/rHgwfkSsV22BbbeFc
hs4uv4Uvz2A9OR+9X5ETL+p/kktNaFKcM1gmsv2ayTQxdxAkc7mD2t0niT6lO65i
c9Ui0mDLnLxJWZ8TKN2uHpxgUwyJirO71sUfHzMhFamKcXt6qO8I6YcHAYAc8iUT
ZLIod584V+Q+jwh+hhuHBt547Ya9etmuuzQKN1tYmGgAENx4xmERONetDt8MOaTd
h62CnUHJdshNyW7FvrYze/OLA7wNCIZ5h6bE/x5lXs3bPXde05gODbQRzFNlDSPV
4u3uq12YrTJt8sLkx57cto4S4uHdL775Mj19u6QJDryyqHSjp7OPhCQDpw+pd1XT
8cD2uAfOM2xIsUPV2ZMQfr5jbaQXYnI1v/+jn6kVEDNzH0lI95kvaw/CEYqAutF6
pPQUmA0aMWQh6hREAKblmpoCHQ0CqjY6mFD7y8oXLXTR1d5CzkqV69eJkfIurtnu
Ir9ENV93wFVbDLHzmAAevGmzlQXxk+zJSE8mOhn/T/Lej9INt9FfICzPErx2jotA
w+QhWieyQx8LEzTG098GQzMKHYRdSSxuioheq7574Jk0eR/pRnZ16reU8Bp9WuOD
ti0Wd0/YiO4bEfCfImvGkERoTJOl/DhKwLY2wnGVR3gEnaGiICTo0VoMyLH/lVH+
0zA71BiEqRSxgdu5ajWgQ4EeY5GmKpoAdu6Cq7HVA0vyMokrF2OEq9tow82A1DDx
Gx7Jdfxg5itW/Gwa/C2/hegd92ay9OWtf6oOHpU65rUGq/APE5TQ4JxzEC6NEz+p
qwupmCKm7PqcClXlHFSaLl6HDOASa5JRfbiHdB0zjjsvSFrJH0O1sDRrYRYop4OJ
AYDk+S+6Jtlb0MiZLbwoRcZTUbOFWozuOQDFvN8EFwWKeHSiMTUfWV/QWDdmsOfP
foEVWQjyi5ua+M6r2FHMpRUbFqsW3TVRtRQqn2kuTJIt0Cxvdj9D4dnN5H4x5tDi
Pr8AMLc1RpY069I8RxVk8l0GKKJ+eUEdPoCeUgagauts5AslmE2y9EuqZiWr8E47
rVbMuw+f43UMmctOZg5Hn/rV5sv2rErdAI7vs+DC18zBO6RaMzNH3/SmGeAXTZTz
qu1C02tRRj3WkzkwEsdMX9QQbLFH/21hVTvxXIBAssQor5svkprOAaWPwWqyphlU
0O+o+AKEE631CAYTnAVQtVpbPfEKDMvqcHiVdRfhO9pJhOggOXJW348fzAhvPoy5
+P19Lx7N6WqaTB7eDfyIjZvl5yWVXJvLNjCHdVAIPwHML8WaGCgeZe89jhDKsYK9
chjrcd55UtnVfxL8vWJyUnqTiZYvctEU2Ymd6MiHf0ZR8k3K9seRdZdE3evmbPFm
/GBnyW8lIdZ0oU0E1AbGWlQ5kzRrDYHKFMkIpcKhvRU0xjA6sAEukGi6nKScGHcg
0Y82iqC6MFl0v8sEfC3euEmuBpX3rYNxXtIFzYtoJBjuAgnODmZgSe9sGPUBi/Zl
SNqikTAtAx6J3SG1IPPGdfodQ89LNLIkUES5bYpd7NC2M9pq7MlMfcS/dTBO2xEi
rDKtVNcwcXx08uEhAiLYcx6KwfSNlmSke3x1SYiRhPDb3WxN+COD3+hQbnUxA7BC
YuzvAsV9sAClWo4VDo6REZdgEIDrWDCfJM7d9514oC8EXr2/qy6FIXU3JpS+bAZa
piR9CVJzHrkUlWp93Z5IeQVbLX7E7egz6jWbul+oiMhP2an0cpTApIcdhzQmNW6U
SYpxYAGOUKxOQtkw23EhbAXNt0Shr85tyYYC2jOHwlpyne8u8c01rJIkFIXeJ/kR
YpuU7N8zmkdFjqm68xe4dOyf/fMJ/QUdsKMZ0jbUXQN85QGM8thWoxQ3+X2/cPkU
TFvIiLyCrx9A9Rmzt6PKVduRvHHEg9zRCCni0SJ7uWw71wlQeuN2HPENoWERHivl
QDVn7SHnm2aQ1+SHFOU7ppNBirdW+YNnxp9eKGM6VCSEcmrYiNapiQcfRSMY2NF2
Hh+alwF9mZNjH3CrvWZXIliY4j5XbGEu7f8IM/sPtDTKJHo5e057t9Pt4PT4Bro5
kitXUTx+r4cfMfdox+Xwg+vAEpp1fSPZLO9+GRj/yHo61R6zUv1425SI4eacW94w
kWD7+SUTV7V7HNOB2hZ4tO7W3uw5q5UzFtATZ0iS8bpXlcao/b1Lkax9r5iA37gh
K5Xgf+D6OYnXXvvx9bG0GmXelwgI7x3fPfeqeiycGU7RrAgA8EU7tw49e1LoBPyO
ZtcxPIEiBHPn90xkKWkwPU3MssYtJy8XBN2XrwKyavaIy0Q1QRItaoeJfARiOq5c
RSDU4VpZsq/qK/Mk7DJj/a/9lSTISFzmSddiLVCuVuvwqzBVVqxMyS2cSKEQn9nQ
HEtJ15Ex3WPk3zqCl2CTw2RblPrCu8bBvKtmaT7I/NCCOesKOOgrsw7SJeOxcUsu
e16dKsF0/7eI6hIs3+UPjVYhZLF2kiSj87ZqeNcdbw9251W14tspNuaQeFEOojoq
2+1C7JMBUigAf4emmUOf36QTAkojQTCgpMNJ84w3pmmIclL/17DDRhx1466ELFTx
UE6di9L0/hzydc+NoatRZ6cIWrFIzglXKcnQVDHlmuvVyXm+FPeuIazCTpZ76Wqe
ZyoHKmCS+p4TK/TEihFwxlA4Se8P5laOkW2rD6pdUz/8LaWGxq6ETgRoET7NXdOu
4KKOzubXj+YBro08iv2HYGL+CiohDmsv41TrloXQke/7DLHByb+AB9xBBVUbHmZd
shkpUylUiGAIN3AGGX8cMhMANus4ifsbjPjTglv2VC90WkkeXEqPOOjSlDI7jwt+
1Z2q3Rr4MCeIBVsqm8vR7NiEQTB17+/tnHCRRhi5hm4aCDtAz46YELEah9+BqYtu
d/OsutRbN3tKNLvzoCn/D43QQfTA0VQXUJ6TRHQF9Dd6t4dWeGYRJjgKDOK+ORay
ZuJuxm2gd9rt6X/w4ChkJFrHVOpZVSxt7Vz3gWkK4RGVMWCQzF+qcmgfO5zw+Pz+
sY3HO31B/UwskA/2w4KHxUIU6uzj0E1fc+gPUBHTQcnwOl1B3g9ahKbodH4XaIHO
D1ffoGH1BwhK7pxnNA+62tJbb+vlkVyO2hJribPjQvRDTloGgQKatlwMC4CXAq2b
J8ZF1r5i6c0ffQhtGIax34gQMBE1CbEdo6d6rm4ddqBcRpLC+UHo6Qn5hVAazviu
BordIu4freyKVOmS4OT/zkCucfDLA2gMlFyyXV7e0e879j0GGVd+VHAUjKZcPeD8
SDc3vggaZEnmu3YT+6d8dCTvBTu2DReO+SlfoFaz6pOzIrJIO6uIq1YivDg4WxC6
nzoOUVD+WAhErA16G4nzdU4I4aWGEPHZmZ2KzBJ+AdLnsYGhhOOB7x19CveUfWBc
Ult+DlVvnIePI5Y767vLWDIG3yLhnIOyIFexLmiV6G1a7d48xaIk4A2zH7BNiIAg
Lq7ke8e+mNYcjS11vc5BUBl3PgANDnrI3aNzlDxyAJhLKUiDaKShS37NqbtfK/BK
TaSRpwWKJ/nCWOwXAbyoVtig/5cpCJn5A0t53Eth8pZX9bXWc6J3c572zedB2C8F
UCQpmnS6OL8RauLQ8mKJHP+8fHJhdy6BZl9QPVk1+CkWazIuGI7kp6eHnVKZQvRG
gS2Kp1FOyI15a1ww2QDdNowMt0S8spO5hVIxO83PmFxsT0IIV/hWq4cv780eJZjq
t544U7UMIKvGRJu2CuBaTyGyfElwwvqY87Zjvzh0xzNaNWQqEZ4K0q+3c1Z7qJ9Z
OmAuOxM3lhIWaCZ1VxJSAacCqt+tHNMlCxzmbJxTtspp31qkbsmYzutWLypolan1
cHDmIX5m/BGuewjadfNkLzgCVUmk0mIkN/BDEDgtuTEU8hsrq0ozNecMWJP8xW2I
4W0ZE0g1YKLoLV2ZbyeGye4wkU9InymdALYx9qM//+cO3nQZIxKcTnUyuamz8OBw
nJGRkZESYBo932ztx30g8GkjMJQUhfVcdqXUiDlJ3tKogJgwUZ/UdeKf9oAEk0Oh
glEdZH2SDcGuZuTyDf9cusxM06U119JH9JQEeWyoE23lZQcTr4qlMThKi8S/9Pfw
roT/KH1salO2ZWCMTkXmUHz/VPai7AIFvWw/cJMDJdEQcnipC0uXma/tCrGmtt7o
eUdHlrFt79CHWxzPiCXaAdc29stYenILfm6XENhzJ9p4Im7F2ZD+ylXoLqgkQkYj
zzM8k7NReW3tyySMOoFsDd1xyWL3/2vNkYZTqSqqmDTTJITC/v8aZisc0XRKP0IB
3tlWyubXcfs8bU4RETnyKt6HCXoZ3q86oIrQaIevcAE4l2U7pfIzCvx6+oRBjORm
h7rLUx/ohW9Gu5EIrU5DcKHRJSi0rqbBZdkZDGa/2yYpsF6gi4+1T4duc0Y6OOks
8sbxkCEm4ZkSeqox9TXb413fW/k0RlxZbra0aWZyR+sPTcUjJYYbKBgRDayg0nVo
4WP73YXzTspcC5shHW1X6cH82GAZK3ABuRSF8zFVJtshdJ0ZEVzNI17hnN2DR+wX
tgRqGXP6SE/YuGwvb9KTV/8YVDRdHDTV4PTQ7WE3/4S8UeSOUBcbEfwoWUzH7Izi
rAyhvPDMc5HmN6huYZHHSqDI6VB/h6GFm4I0iUtGka+FvqzceAvFGDVfOIhVTh6+
/O1CjTbxTOcFQXkz/i9i7ezp83oUM9MaGoMbwu6d/EWKGWoqdV6jLEXm3a3cwZ//
3FJTZK4TzXQFALYsRlVofQYmNaEyiz6zNLfshfDPjSjlkZETbQ8z6u99UgAa1P+1
wzdHpVzU2pOKFPZcBTkvyai83InmgLbl3IIiIx0yWqGromEQgPtk58jilrkx7p2S
DXCyyjtqESE1dggNnBZhyHZKQBDmYrCwDYRqQqrV5F7FPa1WL2oY+yYEBTJmrSlu
tP12Pl9TrqWWC1s7jCma/KdcRRGyboo62/H4CJORa6VvmngUmD0ZcV71BZGjH8K2
zy/A371e+20sK6WxTgxZCBQffrP7sYis7XHUNBpLDIL0XgSvUiN1TzCboCJjS/jS
jBbdA+NF0erJgLiut7U6va+DtUpi9TvVY2CZrmjR/HB5HpvHcCs+Izw06z/b8JK0
PrAkH3ODYD0LMrUXk8xBq9U8N7Fcy4pqZmYZ/EyeR96DJijB4twcOFQqHM7gOolj
4w1QvgkZOS5mfolhbMr/GGWv1Ye7rW35e6ZspLIsrHTfyhQ+Khg9+Ur8CtyWlzgM
Wvnok0+qht0eTquccVygTIwmh+7sCPFRK8KOHHBW/tPXHenih+vJn0hyjnG7/NGu
S6lrKAfxnG1bYRNw373LrtzKIKezSPTIsShEUMbtgMFpjaqlSuWTGZ83e0AB/tPl
9ysSvyml0W1HYESCwq+P8mmyFLAswc+TFpYcxWmzNkPUcwid/s8WRabLqqqTPChW
VvGRk5JoCcig4g8avmS/J4S6+t/kVoNzVt5gmJg1URn7l0e8nlZcN8MrkNAXY6/B
az0FXpuzPRqC4IkuZUSFqa+1wfQUHL0NASfVmONTTZqjprDh7caNim4ewvbAsEY+
4gOe76yUVNKEoSTq+8XIlcxH2whbw3DDFNnfwIftfbHgdvxzMRsIUoHKGEn2fSOP
pHFfmOb69tnRAspGHF4eJQbEpvouacOm6zKw3WT/sPbXGsP3+iKMvCPw1+T7/Vud
im3EvBk+/bQJ+UsNf2X5L4/M3LwQBKHpTzIZkqztcg3cYZRyP1rpUXT+fa5ss8df
SPYO84EEI8MBKcEmKMXsePj+eGEaBIftLauPnd1ur16E+BT7OPBO4jDgxFNoBTCZ
9EOBZ1JePW6nWIaRA2xk9Bqiabe04PB3CRsUo2l7AYcCuU/q2XTE3Jo2moRww//T
K3yNwroR3n+Dmcg4RhYUTmjaqw2yQjRkWZBkTVXJeJDyMRY/ysto0YrWWiHkEXpO
ruDZHN/L63aAJzCXNhxScKqmxQlnhYifa/5M0H1jFL0QjKkYboXAEJLJCEXosgId
807QU9OO5AemOzI90U5+d1UWny3TXHjDdDpY8cj27xn3675/qS/u4P/EODvXj1M1
EM6HKCe+R3F8mTnqbD53s6iadu3Kt0LlVNX7wIoJeBV6ZsFpIU2mM25unXYCoJtU
p60kA3a1uDx5Emh6CCqzamj6Kokl1iEQpwel+QJsxgTb6o0EsY7DusXZR90dEb6l
ZiSaalHXcf60pRC8IhfJxKsbVRFQBCF/+luQ19AolgfRmMoH4twevLnzcf4zxDIO
HoEDN3GDJr0WVdXuoFeFCv1ccwjJMazUf5mCRjf8u6EAku7gYM44MDjLTFboHC8k
2KSl9xEHrnAZhQGFpH+d0WlCRJL1bMlIfycEwWRJonk5S1YnFax1HgCjiUVWYLWm
IxcyznX9x46zC/awItvEOx8Pjuz/KdRpvFTgnJY/4g33NoU2EFVJJ7Mbjpb+AHXD
aO49hHK2XVIn4PxRLo6K7UfDFkHs7doLYMVNFqUflQUYJD/UAdSiSqNAEip6HVdr
jTOfM9PQK1bzmvQtLRjnWwR4G2UKp0bboeE9VRC0pl1/ST31OYAGMrRCP4BaHIpz
xE7gf6hP+sF+WVO1mRYU+NyX/dqvqRIxn98DnKaKFo5RZziwtXEmHSLY8FNDDWfW
i3y4wMW34GC74gRhGuOqBfA4kFHegeKJZUhVFaOPkZqpd9PoegwSue6IXSKMFa/h
rAjFNqpi3rjXI85wp53cNjgA2bJDIMyjhA3Xj6H+XG2esk7uN0Phl+gApY9fpKUe
zEAEhKmB23zwWIGoYt506d0Bq9i9+1ayP8ARVNLzQsYihiHEwDTcYZL+ielf1JBY
xYRc/BjzrvacCBMoODdg6SQmH0qtqFVB4fI6UrbudUSuObiQsVQ3ZZ95vIqk0Bx5
em50iJFiwVmwqgCDu5vFbAf3DBEV3pCcphQTtJ1KeYnKkH/EfUOg7F0NfP9sJ2hc
EIDx//sx6znbJ0klEbynWPVHblFsFdUIjyG/7cYnmGfNhW0e19WSo57FscYFmsza
XFsJr1r/83D3683+7Ub16ATPR3EvyaQWb2bgtyQpYeVK//mCYkMLbTdhoVZH7SQT
UXtw2QJ5sNxSCHBpUl0F1tNzfAInpOd2mJtRFy6h0jXF3RkpoFg27gFAO9xC7plR
h19ipIZ3HEjp7KZIklhvmwrMjBsD0TzHwyoNNg19J7qhWukeiXE9ZBaHVEWXJpAU
t2MR3zE6j+SSgQLjBRusbjGCi9aQpqIuvmASwb71uWf+n7WQD9+YdR+Ip1giJv3t
fHHNEhyW3yiuwophaGXldlPyjk0Lg7xljHjN8Pj1V5AiqiMKRoR59u2wfkw8rO6P
Hpsb5/prrgDCe/lADKFUZM8zIobBOxISDNpmKBH0Cn5Ba9CdLfJ7wwFxzN2/GgzM
v5roChfv3fKhXkQNDqwcwL4u7FSl3fFdYozJzas4HSc5jv2tqXHNcBefBMsk3pdf
ZGA0y0LQy5WpXgAVYBKxbYD094OdQRFeaB3Pl1owR8eQ5erqa88UYz+UxW6E3f6d
gyCMwE+PkIiNuTTw07ZMZpNHW7EzhUP9Q/iuKvteuebvN+INKACDMNZRH77DHMd0
laSrj9R6R3Xt0ccORtMHTJ99LA9inU8wo/j0Hxd3euPQauR+l/opdKWTjulQ7wO6
+NI9I9FxhCjn9M/S5ymbVl4fTRoRzCOrNJunsOG8g2zQjU8dFC5Z9vch4WkRfHfb
sY9vl0hqeScAr4n6E31eW22CRvPv60wboXkmdkRm8WuL/Ufd3fcWLwScxf5GRnpl
mviLl1TstrQg1DdQS1y5YzWEyLYEuQjBh5uLlA05F95K8l35FleAMAnSyVH3OPBv
HDpwngOorb7MhFh/+8eLzD7Vke3ANyxxSRyOVkuiVynZPXVZBmq2m2Me5XjGfUMH
W7Rgs0Y6WocxkHVhKhy50+W0L2S+8qPZNztSBmQhMw5/IhmKanK97dTkvRCMkQ8k
wyA80/+qa7MOKTAvCStq7oR1J6rnNdCPw/aHSf0NHoOGYtp7SJRLtWsNVIXhxOpw
5bMCO50SwuBfkxDfknq+Q6aqfcjMG9rjEFxiEQYRTC8Ct6OvgHxcYw/oEGZurwog
fJfT+ZxHHC2Jz9FN/q28aWuajjk4bHp0llBwV/bfYYzg9yzuCVnTnAyMZlCR8fEV
flLfC1Cz72kXjaA6Izuu1YIHt2sjokmuDMwqbUuUjgwuZo27Mvs9Q3U5qPz5So1O
FTAPSnpWxYgP/NMtito5u4CKjMjc058cinNKNYB2T/5zew+RGiGU8T0w5/7YLN+0
U1gY3eRJ61YmJu0Vk3Zb4o8YF59QAbsQcNCeXgKyFNLMcY7ByXwZHR05ivvZTp9s
w5iRaj6zih9R+X135u8gI3G9WW3DvDjJMZzT9ZOInxF9fzjmm3wI3RglSo43/I+O
ubIJYGKkZGHmfOVxI1eEslMy6Hd9znUVTKwWzM+eGYoQgbj2GLT86CY6+RXFQpcV
t1QhNFUXmsjycPD65rE62GuhUPQE8JCMtWHgpJtSdCqsRiyTpfYUVmwpwb9v2Myi
brQghI98xj3aPTKhOzdqnXljnD3rfe0gZUlJJJi496Hu5V2eSKzR4lSRpi2dFVS/
f8DX6gnUc0eX3ANTAy9ZdrkdEFdarVARLyXYGO2NGOj3JVD+FTN/4CMgUS886l7H
UdbqZi8reBneb0rqrFA8A0j+EK8nnylidbWToF0EAg593uLEvEOh8ugBXD3iCGcx
RNrjnli99fDwYehsM4To/52/YNBs8lpd4EakCjhwnuMBLz6hB/60lwYKw0qEdZhc
6hFbamSkdt9g0UEte4eIz/D5Z8+bHMbk5uZGE5eoCZwtme16WzSSZpKtlTd/MxQw
NV9aT9BJ+H+KLwlPZnhbL8O9+V3yPlF33EZShVowTXPY6HBiXWfs7EfrDjROItBY
OccqtZpat2yqhfVFmubmnKeu6DFeBjG3upOSNp5GqYZ5TEzGPvGBf5/0dVGDVJK7
y6KP9apr+CrYwmRlYUoeonruBHJWx7h/m2/Qv8EOGBiOwWgNl81lAFZAUWeURTWE
efa6RxTBi2szqEgLxz8OuFA3ZKZaH5JlbUwivQpfuXS3UhA/9r3rZywC9hmRflP/
QCmgmTXfi5rkxdYyx2uAFQTEvDySFUvakDTg9/t+wwc0uJwrzbUpIosWP9XjYQV5
3s7jOxy5OHuYszpCaMLSrgXCIxFdcMuIAP5m51dEbsw6mnbIFAczMkBMhXDgo2eK
rpOYpLpFF+B0UW0TROT5u1UBbhE5eRro2fTAKmVk9LzImT3SQyNKtumuvR5jSPAt
0V33nZGpF6cjgUMNq3SuTRaJlbkH98Zqezqd8iuotiJ0R52gOm/Qre/rfXu4WnVW
58+CeqLMMTxqkNWXYAR/6sLyqItj/p7rItsMkw+axWPZpAXzgLgK92UUIZ4E8Ouo
o9Cp8Pyh+gwwaDoSqu/QBL9SxbrNE/5zFddHxHS0Frzha3d/gr7bFwAiK7SehY2l
TrivJQErGMt4wuRbE66l1Z1PvNEmUKGrn9t/ATxp7vtImybPOx5wExZ00pGSWhY5
9Ij//gQu0o0WsOWhDg33If2EjTdILe230kmnoSHFIaZ4L5jHmGeFnRZVwSS5elmO
+GUa1cu+KJkCOiISeDUJ+u08ZdFAEIEKBRLkPchZAfZkcggEsvDCom8cZhDdh5Sn
XZSxyZI0gxgnPwsa8vYNHM56u7O+T59S1kBL5rJZt4+60bA1GJti/RvENaxDgSlJ
bZw7ibSl3HrCHvwggDxVO1WeOG7ZExTUkYEns3+ts1XxNxnLJ/WaKcs3g+XqI0pE
+cCcr+QiFsZHMe032zTi4bxaAtx2plJZYD0PXPYO/xmEF6a844DIAWdM6hq/rep/
M0m3HOhNmMYkPoLYSYbRK9oep5JffTETAfMxNEI7oUv27j6eVNOirsR1S3HEOuJR
zPWwoWQbOnrrWOrrxhXaLq+oxkqv2rNZ6CrlE7THL9b5LqGYfPzFBy/E20Q1lgc9
Db+GOmKTv/T9rhyXckjyUd8A7pMbTPJ5IM8KgQx1slnigjcOu8rb3wrOlOoJL3C7
Tg6eBcz6hNWHb42oZr5qhuo3GZQjvaMhD6JKVVK65zymqfns3WM1VdI2apsA7lUn
n1u1sPBoXKMHmMFSBtzDMQd728arV2o/qa3+MuZ5xeEfV7pOjMQvIhgQ9lmzseZt
JcHVHMuAkzn4YyCfrwkrS79WTI4/GvMp6T6CPrRN/xPHxBBqIXKDlNfgw73tGEvd
nnz4BCOpD68VsDpRQrYkEtGC4AKH1ZAti31qGNCYoG+zUVEtJoXxPtw/zMfbnTUM
jRsQvZPfNSmPQacijMyazM04n2spmT4ErgrHeliN52nmHPtmw9EsK6D4l+aMYoKk
5InRnwAhIxxlCn/U3nR9Pbj2Pcz8aONbXFjr6nXzb6N5ysWbZKZVHKLHy9eDNuql
3U+uf3/DagCcIT650wGD0WuyXQv3sRluEWtMKJ/5VYv+BcP2Y6gAqdX0SCp+5AkO
LVkuekv7KPtrPjVcDUQxQSfIXVH60vVeAhsolNjExJj7dn2LnkN8GW3SEFRrCrJO
ZdZl0m3DTGcHkObW8hSGrfCQ4VbtfT/5F3JdN50Etoi6dW637PQdBFyji8/oWLa1
hUJD+OnipwVO/TzZ7qM3pLVUvI4Yga/Ld9VuLmYxb16y/0llZC+Ob6GtO6cr2cSi
if+fPmjIwa73HzsawB074O3Q3Xgq1Xm9ddai3qkTs9kAX4JsclAaJnwTK+Zwvzf0
DR87emR41B/oDwmku7byyHLZd3vWJWnYjSUoOKkpKcpCvuhWC1/ATQufCa5f3EAz
+p4+p9UiNT3VLGu7wStGS7uJ/4csWCZ3Vt+jUsgRoEGMmhC5sTcm/MbBrVmnYvme
tbfJnnJu0f0FUPl1wjgvY1vhbAdBXJs/AqMBFBWrjdkU+p1uqNyxLFRNvFD64PZA
VIQZV/B1kFNUtBx8JLC+wS3Fh2Wtjrk1RS/rm1bozjb5AXR8VIipVC1ahxjvpVHD
I52mjrY+rCZTwuDsVM27Bc07IdlfOSw6dKs7Am5mt3XSN/NHb2/p0Gc2crln8b+I
UaVDhXrk8CtYMxKzRDY0huIeSuqzjJTM+qvb0MoQ5wXrEhkd7atCvJN8j5+VKaAV
DnaeF6TpvYpEiNXVsrJ9PlG5OWojU1f2IS9Z1Rl4CLFf3COB5xB2SbtAORS6zojY
elUGwxr4/UJ+jQ8CkQv66GQqZlnyqIBxA6itQcWv4ib/hsMPfw3hWPex5kLrhbu8
THfQSKyPSImtDzr10aWNveIZP1xDFDjib43bjkpRo/uysMESEl4IuZofH6KT6Y7z
NePRcjU8AI9Cmo0agKu9Lbk7Ao2+S8VSdjzMn7bFVpzSH7kuYOEdA+iKv2+jFm8p
r5L0ebtnQq3Dax5dSxwuaw9nhoOGch4gKYUpvETUFGjAbb+vy7Bgb0vy5Pz1zU2V
AeiXUQMriZ9Hb7Z3/XTpWXtUv33RGEuG4r7y5G9nwIh9YBFAUTJjVcbRr66xc+O2
QvHz8/l5nv3YMG7MIA36WEw8Y4IP6B/01NSiNEy1S4pIsHLodTUPAXLilIJ56EP4
kCtt57v24MYSzC2RRH/ec/8+3gyEF2vdqZmSumx0Ge64zbgIF8jqZ+xk6KLGNPvf
3m49iqVUvYh939S0cTqD9SMzVBdpWZ8ssbSjdFAFnqHb9S2Dv1v5aAYfBG6A2OIf
JYPOa2tnDEG0//QpWRuHbQSPS40l36463eVJyP4LQe9iqDGdAj5BtPnlQ7PzdVKx
crLzF0JlNgYI4X1XnFba40KSCF9lEx32j1tO1u2Nc3iCD1LLdOq3K8NbEM2iSK/H
H5BUJviN8U+NtDgGPMvizSrm+sNFMITqXgZhbo0PJ/p5UZf2Zven59EjQcqLZRga
iJQNka1D6uGfBwFhS1TKw7JyRHvKiEyLbd+/Lg0KPuzewAxi+vfA9caJ7mJnOmwB
B+oW6VT0FZ/Rd8Z3rSaJIzlbaINSbK6l+AmvZkiSw+GSlF8DJOqLwRXLyd0x8Sae
WmjIq34BCgd0NfRi72J6LE2RGl9kYSrfFstQCt2qjxkjw1QbBrPkaOHyYq11soU+
k3LcX0dBSV6uMfWJ0Vx3QPQ0wHBSPn7qTi8t+wXkTE5Ky56tuNCcnUxHQgkkjfvM
mYAL9EPwltw5ged2HoqIznWnkl0KUnXOwfAHkJtLBBqrVEkNa6X8mLUP0LNIzWRH
eBnIBPwYj6ajah/uER1ZSfG+QJsE9u9CsO7p+tJNbbjoFXonvVj7EG04l6XXddxb
x1iMsmxnpdbdMId6rN//pyhGfKz/6ZgHUyKFrzbiJRGLaPWFqwJa0nw0Yx97ltAF
7PqgtRVVL27AhbdzAY5ttomqUtSlf+5FhGXjlA+SQdcM/ye+xvR/T7KwDrdwCpdY
rZ3op/bxa6fJ4G1UjEPAWz6LLBE7pwvB4tIpVJDcu82abT+AzhyWpzr56nOUGzNZ
3OwRRH4KtLq8ZfzHxb7H1HzJyowVTkA+hpqxalsi9eKcB21cxL74MXW/sf3n3njv
MxcIFaS1CLd1Wq1UPYDZZGHYG9eXox7VS1VRwNEqRGywAptHn2MHCahdSBR/HafQ
UR3S/oxlfUvJoySiZqwJzsHGNNIPlXZrJ0Rxl/BdY2PYQT0xI9hVcDrPn9YqTxZQ
jnoUqtmac7zpNqaiEmvRxafgGpKvEJ23OFPuW6LT8ifbGpvtFldRZShjjdTJJ6zd
7H3A8s3x5CegOmziH9qoOdAoMSDHdBcdcnQSu40arHpWtBh8fTCplJ4NxU6djCsM
kMRaFevYjFq8816zn559JGhbwqArzoRwq0RJTDcomLcbgFqSiZuXtQFTjby5EcJW
NvGwQyVReUVMTkD1D95Kk7Dqx2IBQehrG9Gimh46D+OgwhHechwiPG+mQQ/u9oiQ
2ZJgAxlkogt9Dqjv0xqZLXtevafiz66I4CIDtUv/Qo0uGQxiJ2r0HJBmFkqhYXfc
mzmgSptLFuqXDKbHoH+tbMjKRyH83R/c0iofHMtSTRqdbMxxtNiRgRGPJAmoZBlS
Ic75uafipeiaJrbpIwwZ2FXEyKE3IujwBIHj5r++/z1EgLhrq4+Smsi2bxJbrrzw
IvOD0RmYuzyMRJ969zIZE5EKx3ay3bzyaq11PvXEMfOU95ssQeNuXTB4Hg3XGCWu
uY+05nomHrR5vVG7z0g3Svsde5OAYuEenuEBOVn2EbsAWs5Rx0FNvYR7sE3Jz55I
bo3sD0i21ks8Om5CwXYZFFh+l4SkNf3gVXIlk4V+sH6rOZkBZPdQy8G6ERpG4GHO
9l77WBivbohHmXYjf+Z1v5cBOcM728dMD7ffDIAcdC2Bd0YeNaVF9zG7LXXBYR/r
bH0FuPtiOOH07xvQ15jf7UM1nywl5ulXISdxAxO4Q7i4MPfu5RiekUhLk4NzG1O9
Es6lyND5lsvdlzaF7cYef5jLTxpxujaxgnvAXrE99AiXFDbKIWzR+SJfPhKbVhF8
zXYcV/pLSRatRd8DrHcfKkmyu2kr8+KK3hlZa8sPQkGGCAceJTFYJa6a/775cmcF
IjCROpl7S05/xt1Kux+i8Iz5XSmx+FQUu9QsA5iSfleU8pVyu6gKCsstxFQd5TV0
c6onKRfKMmdfE+HhBpy8TM9sMT3dEFPy+foKehKpXCuzXbHpaNbfSMxZVKzoay3e
qLdK5WJ1MhFx/2Au6irUgLVdY3txOx58GMRhxcSJi+sTPOe2EuIHPoh2gfr136nv
/itFbdUTbBiqNHruq2E7RX6vmTLWBbEBkgHFECa7m5DVCLKXzCd40wvYXvwEd5RW
FIWQFVGVIktaIwhFUohRMFOww6p127X8WsVkRltHW94YUX6SnvY/wzP1tHX9ZYCo
IsJ0/yd4FK/RqHpMBYjDSUGo25GXLrZdbqpPhkBkidJvQF04XYVj7z5SIL2hZQ9h
lONJywNPlReI4Rl+ZTDY4zr8IeqoDRjAX24ui7pf7BRhcht9c2f0hY1+2lBE5tlk
urglk1okU2UTAYgxNeXxXD/xA06+rPPaV/f0EKZmKQLIGd4HGYxp/7wu2YvXl5dc
hyZGXIVH2ZlmEViR5g9IBi5uBNGZVa1DgD0lfCfKrgu2jE1v9Aa3cob1NeTH2X4J
4A4/Y1XoZi3Jjdz2ewVDqqB4kxtaseKBL3GiM9P8il+ddiw7+4MN4xv/StbWn+XR
yYYLo3cQYWbc7fWA7/FrinV7gtf3lxBXWsjHfcLxTcjLEDDxZm9wG50ngDAxYRpA
RiS7+GKIh36DmeNmPQC16mOeZ83OAmA7Y7TaPW021dcVolGotVT4OO3nA5SO22ik
4ff6Q2ivilM104505Sa8PmS2KCuKv6R97s01np/TIyw0tz5Rb7SJkCJB/wCrJCZv
0UkqymFqimYQBQnKZqzIBNWNopGdxiBlhfWo2ZQAsqO+ffaBvsIAjw8iqvBdbVf4
jiYZeQsBiEht251cjdQUESS0VT7xbW5lriEZXfivO+ZC6fS5ILjC6d2Tjj2TJMt5
dJuyDKccL/wU0AIYFk1CCBE9w/z1Y0OK36i7xt5w6VLABYwU3qTs3V6G2xQy/qJ1
cl3aLsLOQ/aoMl7E+Ikehuw1Z3p20B1qIyEib6xquIwCOU/cWew3XJq1cebMRDUR
lU7mtPxZlX3tI1qfJQ8gi7i/tEnDfLpF99eaUd77ZIITcbdYncbEKTGzV9RrJbE2
wUg0sJ5xrRmvuk9nWNJThXdalucWEP2+RLwcix2rymE0aJ6r6kgit0CU09oEPovN
X1mNtEi8ckq+WQySTkZ2BEFXSoDjV4UDaxKg2Hcpre+YdB+BCMP98JUrsGYHTnK/
l7Cuzv0pIkDyvXgtnLBfqalh1VM+1p+hlsvMSj3YJHjrbUveRfWyv3p7Dn04qcUw
Py+Arm5PgdgIKW0qTnDF76d1lU9bGdv3Q9ERvP2C5djhECFjpaIrPacic05wBH4b
YWbislpN7kSzcs2b77WsKVQfxuPeoBt5xSBmhBtgLkUSdytwVXpnPWag1yrLPgcl
qYmWmq1JqPsuEiWfTV7Ps9CRRRBV5VIP3acLt1q/F5iNzWrtPBpwkl6bDsIPdf6a
khfKW9nM14/T95dPlE3OykwtT5oIt/bsrygSQR4ZsE0rOdRNfxKB05pK+vXV1vOc
3StJowpYtoNC3Zd3GCE9G+N0M9tnVxIRWD9J3Uulx0Nn8l0a+Uoc8Uf1OEQMj7aA
ZKadIrCoIllMhBvQuTvHWgN3yrNKxWFu6O6n8ipmXoZ0PCiDfY7lcZFSiXcgR4Pd
yoORjzMEnEGc04f+9kuhQVCIInUq/I2QXPEFJOi+W6l7AKxGFPcDMSw+5ojRQ/FA
23aWtihFCm3m0H4WWm9ucP841vjCV6vImNWr9BzgtDCioHQqsp62tc8WrFSPGGzF
dw+OSwbXI6jRWKtr5iicBq+yWYMIedSNxFuysKaRyEeuh7zxKiBmL7IcjjD1gJAF
MYy+SfJ33u0mAtNp2mrHbfxn6bIn1B+xT/q81qkss9OL+xWEq/l2WiE7aBE1Y5/G
qlzbXywBJZve6oh2O4iavBn3JSnQmElnAZUa0qC+jJdQDlMCHJHF4kFViy4vXSiZ
lwMrowMrhwBjnyBhbIf+qdIctVzBNIck/X7pweRdraRDGGA4WdryXfLpu+IFmkvo
l9l+wEFzXyd6d5Ek+qaXKlo586FmDnhKl7tcmdKteIzUWmjcoPiTbt8Oxv5Dv0ym
+5EwRHBWndhPtmuo5jyV/qqekXTUinTjDQ6PBzJa7QnqwPD373igbl7GSCWGvEaH
Q1KQdkneggZpB9tkVl1kwyElgLSmXfIw78hSdKBKu8+gHsfDmDyIXNgaNN6EJWJx
yGGUJv7/k2VNNt3JQ2N5YWiVgC4TQl5CvuS6Ac9ivxjEJHvdIVBYbb0JUwPRs1C7
leVtxY0Q7KPGG+9sGVDaJNOw+/ucGwRUEbbvX5qcZx7KwOI6K3q/6I3/Tlk7HqaN
gb235fAKwLY3/hjvPENgbo61l1hhSM+1pEnMIhBvwpWQxcSrl4ZZS9IBVT7zARcq
GGLOtP4EQRcAehJzhTYCG5m9rbQsnIfT0p1Ur674a1mpyR+hbuMTtnXfmtWVNCfW
KwV2DtqPiuqYKth0TXy61dB/l7l9lcrmJDZPCaOnGsD//lS377sS2gMkB7RLP5QD
1yKCNuoVokAPUOKYEI9Yh4INLZYwBX3Q6NzKRVJA0fHQhvkv1pzpkry/V8GUjxv+
TzhebngOMYI/tYhXhPdMyMQgO9dOfzqIZN98e3C2SnEdH1BRNcHMv5RsIr7V12Rl
SkNwzKVsXMtlDADcH0TU2AYhraKeMRXi2kC90nSMNoi09w3dNuLf+5r+4bcyS3R1
jhwCqhtBydbxyTlNc1dsxhgy43r6PpOTlDf12FOlrOjbgjveUF9XOoG4uuYhY62G
ohXH0s5v9+FYPVFqdIUsDTgHbJAjycZpgbx7deGMMHnAPRZxdtRf+Piko/pRhK0j
JoamQtJuQ73D/1qm4ccxaPXZpruG14LG7lqgoAxfJdUTRZxn1lPs46KbJ6rEi6DM
fEUNKDnmItZC1CUrFES+ozCunfQwT2OpIwtzgbkh1dFwePtfFr0pIo1HO7pCzAim
/tjONnCdwzJXh8jgFtaFcpYDecXR8mXKwDdpxVLKrCsHIHRgbNg7R16HO4asqJrV
MRGVoWaJAyIDrfvk3tAyjLXS0w8uWLrYz4aGHlOLByIFFmUfAAMqR1ZAvjGnzsVx
DJOweAgXq76IJXVpMdblZmK8pJEuXI0GBbRgIZvTMvLls84/bS4ALJypUbfvHq3f
s0ihk6LEu+b8+hXhTBEQGWekYfSFROkaG79wV+atSkbmcz7PYDAK/0oBcLzzH4mg
+u/hzgSaDMoa5Tt3ylJ+6jx28BQSl7miAUXsYn4Ipc5MbY8XgjtyS0wrIKfntnD4
5LsfN0/K3WkEvm4XzPca3rPjipbEIZj9q7yW2MuYUdWKLcE84U4rwaUPvrnYBYIl
n6/YyWZBCDVA01Je56c51/iVuCGDCAcPH8MfVR1o3gv67iaKG+ZvkPtXK1Vz4K5d
MBYrDFn8SqY8WXaErHNWWX2aJYTc5OUjzCdZl6YImSAaY65e45IxzINrzJrnbKZj
4RWfvDVLS6mihW5YG2PUPbmQxdJW4+/FNfw4p5nw+Z0nM5ROdBTtV0Uyhv1q9Tiy
XadE/H3mWqDk7SFkrbNV9E9Y/SFnMGH+JyD5lR5R38/aMI5NBmliLD00QVihmuW6
asCRRl/uOf23QMkADmofDTt0XZkhQAxlNFP+fKzeZ+595G3pT/NQ2I3zjNY99y20
QjXcAaOAgiprCUldACaMKftJR4cFwxXLr/bj/RItzTO4BafNkfKJnplu1M9zavUu
cynNTh1MoGa7Pjc1YGgBcKnHSiFQcmQEBvv/ZgCAh1DjPd7rSDyqiAsaXnnrvSKk
MQGDx4l8iu4ymSRjWQWtREZOjHtz5DN2YYsu7Q79z1VA9jKJkzWhGRulkgo07wIK
XU/k8+kXZYhe7epjsdrGVvVK5Ci0Sau0n8P7ZF4fLWQPDIpTrIKoawjHMZhXOEW3
Vrn5vjYkDAzyW/iw0KA8A/7BHMJzBUerxfBV6NLNSI/P21k3LYyNF1Jl+lPH/aBf
I6ttPsGqenV7Zq86y9LMmYmWgGsTqEJ1XeO5dpDyWhjLo33UOYwR5aZqpW/UcQx4
EK/pQJw6Dw/owLptkcGl2cWb138m/kYr1XSLoEXjgFo6uKyPb5nFUxYeiL5twPCn
v2XbHZVU1mk9Z1VYAvLdQVT81oBICo5W406ZYGQxHWZWTfYHfwzbzT0SmS431jfz
hklUH+9Sgj7+1GCTiaT8QXZxTliSqMbnZYN7ivxYpTKS4Hr+qzZ76Y86DDYI5GVU
B+nnrFvVqyJq7hq6VdLkBP1FL1BX8pLvv83ABUC07sRGLY1XGAf5AyXEhfXFCQTG
Pvoq32aY88CoQUKP0rp8fWrLXLdOgwN8PmxpRMBlgmE3RzJLeZpdwdloxvTaVuVp
IX4nuIMwJ++8OFpr+i1WtuwOUemqBrvLFqmP9VkQPYi9NwN01Iv7nAQc1etIqL1p
ex7qindzLUfPrHIoEJZsdkyTwfMoBEJJavkqkLvk539I9HZTcVQ8fs6oHyNLDMjV
R+phA/97tmvp00OIt9S4eZMXa+F+H2WY+L4gBgxKFp+qewCwB6cwFtaFNvpDyYuI
L69N4UkKcWeoNh2yCf7kIDZ2rgyONW1Oeyfe9piFYE0t9XhFRm+qp/Q7NRSjZEZ3
M6d2xbPGOADhsXGrWZV0GF8v2JR+6Yt/oYaZL7+Uw9W4NZjqSAAOJDjOMLf6mIIB
rfZ/PjP5RnxCqfWvzvz4giOffJ7xD7DykdF63tNmTN6EAFLj9QWqJxT7630er3gp
DyMdDMtuvH7vTY/XOQBWPGC/q27Q4vED/ySo+9C+zc0inB5tdMYV10ybOC9+NP4J
tVRzdmyzfgghX4auxeeHZ91bqg7YuzIrHWkse0dTjq+aelwCM2dhDU8b0BmwzYL8
zcaMhNPy1w5UDi8lEU51yTX56rjq4GalSYC9/GEv6styFfK0vDzKpLKMJdapeabi
mfZ18VtbRAxfZRwegqOxGi5wooM91Y2bRHnrir0fK6EQuHi3XV+aXDQmtyFrl7jL
w0LH/cN/76bTmHAKEUigmiaFj6/LDMUkV+/Hvd+L2UQDKiu5NMlFbyjHFMAeSRXu
XwOXsFzpTkz8kJ4onab2it1kuCp6AyET5B72hGNiwIyODN69cXpKizbyArB/7XXK
ybDi/rpkfi6mtVK3Bm4HKeWmQ+rZJkmCJHFXAIEuJYbvG4t0tg8FvPcolDNILFLO
OHdA12e9WP4FJ96fl6rfZ5zpqGas3mHAINrjb4jI3yfiCBUTzoGKZ0T50C2jh9Ve
/qjkKHH5x5+TgEVxIBZIqsYfQB1yhyOKpi3qZ9WL3oSVMmWbAz8ys01l25Nnu3f0
JFmk7+/vYMOvaPjBZJEb8gV8c2kAYuqKxdqj5UWdiry3OQ9vBG5BISJjbIVPU+Hn
XrlPdnTntlotx/ZbuY5ingt9MMl/0/lJUF+HK1RZ59p2KX2pp0xtxk62Alxn+/BQ
Omt8uZ6p2Be3eWRBpXqByH0rYEKv4PfbO6n4YL9I+eDlh/iQV5UbtycNfVqlRm7f
UE52yIsGu78Ei5KYLpM+zv+69kQ/J0PQabkkD9PNumK3tI0ST/WD5/LpuqfOoCwY
kzDDqr2Y9AbibgKuYjFN3YAHRVNUJ6nyRpF6mIWaIMNnCBCwU9gD8s2t1ZQ49rrv
0hDnmPlFbEd3k6sAF3AUnew5gZg5tPGu8CWE1ZN71jAo6E6Z/2mKt2/aXwxKUWZ3
8asEXckEItfI2XheArcFCPC3FPRk1BmEAWQl8g/OBTO4f6p+NXN4D0YpMChijNsD
kVvOqfscCC25BbL6TeXb9O22gzCQar4JkhicW2I9gSUD071IqacIOXUVymGseejR
8E5lfR7CCrQSAJPBabg+5abJWWezexkInKvJObHOvrWW72ZxNflxjcNYwBn2ozbH
oT3t4yNkEQ6Igdj5IcWU3Q9I3Lp4YAgwojMemL1Zg/H2xhIpNwKFKS/qsxi0bZnb
pi7UrThioJNn3P9/5ynO/KHNwjarejc3EGgP012+m3Ya/yLBe2JJIQ5yrDHNii2e
iCTU8uxR7x9BdA2hEv1ZDHMVm6q5M5yJplrWAP4i0xuZT3T0TdK84jzrTgryEpJm
GKaaWLwhZ7W7ubQSXlEmRHwzkWPi60cZR6VUWCkLwd+S25hbeZp905+Z3hd85xV3
mHeWhVGl6GWV6bD/VAwgWAIL5+AqVuXvsuAbg/YW/xWmaatRMHO3+AYvErEVz2QX
qLlYf1N3e+6uq1+0uHVYPXlCZikJH/fvyP2zsKL3MM92wDu283+JuVFWgVHl0mG5
sUtzxkDz6l6Br/YFAiTSmDP4y3RT3ET8tjakyaBaGIllqU+Y8cNAK6B1ZFbfo9d1
uk9CryHV972yInM7Pd7eSaQBb/mSdI8NkF/3vV3+Ls7v/kTeOxrD9pp65riwPvfq
arD6TQdQ/I3hMIf8/onNrmAK8JqGjja8aeSIouDxvbCtzyRzJxG7abNTfo3BuIEA
X1sNlKR6CYpiPev/bi9ti+PJvWybTILsjmmQa7vZDqb64T8K0luhUvfuQTJh+vXT
Y1uKvKbJcQ+JfD9iv0EqzqBa5DlwE0X4Vr8jp3LLuK74ByK8K44prG3oGTiwMubu
h/VQyw5uWFKyuJ51mENOND8hcsfY7+y8DtReXO9cWd6rNVYwCeoamVy4TT0S56eo
Pk6Z4Mpw7lfxYNgQXxcYrqNsvK0sVAnXxmHIYL5qu/QXNJW1+7l/SJLr4mjtNV6v
hF5z/2G94Yo8pfEd3jSuJO6bXw3kDhrTAaqzN2UJkY/ojLRqXS1LV1s4HUqRWKMt
8bLElon5b0ZW3whCVjiRtsVjS6+GNul4rdDj4WrMAHtD/8CDAF3D0uOgcRLE3baV
AtGLOIta72CePEJ7/FjqUpid68pPjQ3l6DcDMAXkfL9RvUgddGHdQZEpb3kN6mBT
x1DUPtmR2JLeXEUUlkcPum5bPvY8dI1T7vTrMV7dV4GDMiGON5io2XfKwENG8ViB
r+Uve0sqQVCDgajM0pkv9R9PeINXuRQIkyvbjC4tW2W7YZyrmvxVmERhPMzHSrwI
Hj/EpmGbzAegF1C3nLm7jSQKr3gvWzj5LoPZ6wSJtfdYpVUNjSWuyzezKotAQzFW
6yjodA7DWzJfArxGVh7BeQpENfiqOfGeGwprA+lP2SZL+E4vi+AW50a2JVaVWlLE
kyHkVNwuarF8b6ssd5wUH6JC5ZVG80hPEp/tDi5XsQUxvUohfo8+uaApx+8wFw9b
JQDFs//CSDWGVf0ZfI3TVoFTovLdNZhQrLobOCyDERsYECOSjva3w1psWVrrtKoZ
1ktD77qe+8p+DgzA4t/aKg4mdC0fO0QhiyFSLKY9rAxCO6Mug8D3DyVpXT7iK6Xq
GCN4McsYEmbJWnt9i5WzHNgVzULkLgsGWQvd8R6Bu/nrUrz4/eidr83iEoZlnqj3
dIjZ/gwUtc2kb3BYKKB+tjY/W+dL3tvH5pXm7EM+yi/yQRMHQyoaQgZrYsEV3QIM
9XK+7bUn69gEHtkbrbtPr5o4Ko+7mTd58B9OffkLlhJ02jda+tixX58HtmF9Nno7
HZ+9l5au+Nw7STUeptdYmhJya6AzOOrlPOG7lUE/vMScLIzIX3pjZT124/HJAMv6
DbFvxdK+j0diuND94AxM5l5fA7ONJJWVCVnMOimJH48ZENgDL672g7yLgR2ktx5W
PWRNjgKIiXDYuJmMG4qImXVcaRIdCuRgZY4eh61s7og5NyOaZ3Wm9Qsj+8aX2v3f
l6aq3Jb8wtjt3lyt37wJKkwTyQ7bpApA/kJ5NF8yTLRCjpaSVWZ02ivOqY75Q9S+
txNspbHPyQMtExUqV7WMno+pHtVrufPY+S7CFsTTYPkg35lJF5DVkedhLGtktMcB
btdPMRH+n2VS4xNVLNmqmAtlEgDUsIo94f3GVlI+oHak2nTi8afhEOOKE2EThcUz
fSzq9rNknYggqoonmr3RByg7q4fz1vtWNr2y8GT+vjKI2x0PirTY3tdJ9CNihxBA
TtKfExRO2dRrkbOUaCLgb5XuWxg23VgrnNivHYnMfoPSPI/ykgHyGtY6KVD2Q1Jl
utxnNd7ZdRg+1SadAtgx6/s6frXh8hDFlIabyxztNupVC2veBgNRFTkPWhr0WpEh
DlDvFzX97swnYPnirGnPcgdyou4ApU578P8pxIH731RY0kcqhOTG27BcCgWMkPYQ
TKnfYVao1NlDJA/BSjlW6SYHlC4D69OzpPEJ41UUpO+dYqo2grDtBEg5iF4k+uem
xsfSURxvq9XFXBl7RQhmkXk+WyK5AqZjtL/vSQQAETAJC7EkEknivfiQCz7RjSWX
gJCJj4U25N6Us5RkGh7Wy2w7ascy10ofsI+oKTTej856A62AgOublDZrd6avn/di
XzSbFYRf+ptbtZyPCsvgp0R0PhUYu8dvEJmBy+7GiN/X8/ykVEzK3kMuy0FLv4YS
W5W3C8tDWd3zUkT47F+z7iMRx0g7nPM7yJf93y5juT9kHbEv0HD6L5iXZ/Za9OHQ
3DiQ4LyK7zuEUdf1LTdSRw9HauTlZHtHzbrdzYoUwBQGhgAtup1eNqW3nNfG2nV9
vTvoxGs8fGQvqqwiHcPfOv6kPQTfejpEUTfJ5xCJQFEOKZiaeKVfDZXGVGGariEc
FOudoo6BlWzq22bAd/Bc5QOienc0G3ESi7Ze2v5cMw9tgT32mhdde6WBYGnZZHFO
TVOAAoOUGhvhO5474xAtWeVKdzE7sC7hrRYPb8xOkMpkffnHuL2SIUTlWvTheJ2U
t2kWxbPfdpqGPpnKvNjuNlSFb4N+9h8X0Mab25QhGqYzR1eJsN32NCVgWoaKBmMQ
uOz8fhgjFlASRTx0qd5h7Uvw1MiHL7PljU0K/OGAIyJ5NgLimld2i8+XYXDKeEuQ
D485NRD29GSzrIRJ9/zWpXogQV+e8BYBIYLQp2Xgn6WcLUn/C73keBPL6NYK0pQj
g2ozvXkNZwhnV4aqC8FuwGd/Y+wt4ljZbSZlPpXMMdqg6Dlapo6nwGaTgb/+uIfb
9euoWb21rn0bdwAhoSpsNg+rIrxgUR+lL4jOdwcH0FjGhKOyF+qBmpmAAfmMRaQ3
1K4tQu3VfSnPl3rMr8UKU7SAsDbjhtlVIfeSpnvVcDTZL2QCIGmcwPOr2ft9ChWv
LDVombi+8oAs+qJDtO/ThprgDGL1MSEzcykYWctYNAajF/SWFaGaCY52GWA/TafT
9lBIHdauNiT71js9gtsXc4u7o8BsJoXeBY0SXwnzAkzUAs9W3iAIxKQg6dMgJMzk
lio36LPNQC6+yns3+5N/+9kJjvAt84JuWByqOOWkUB7Uzvlb4DXKxlcTAeRg4Q5/
fFixSKQ2WlfPYwhoDuoN2bOoAOIig5LQ7cGxXGpc8GSEwiZ42XUlJc2Lz5gPlgoM
AcIFGqjKRFD9D8k8CB6mGeOvGOAJQ2OQPRn7qTfHPVxwQle4tLyUP6Aao65OLM1Q
OO0tXns7vyPNt0Ujgkz9BJUoQIIAps+P+ew56EUngVNZ2doPareTMmi8Xa0b2+b0
eajDPp+tXw1DxqGa08YzGQBU8C8zZz/GhEhBZFTlq2ZWDCJalQ30H+a7Bu54KX1a
6/tnSSeHq0dscOkZKXmvHbfs25Kbu9EvA92VBMCrKKRNh2X13WpbVBJC4vKm8b7N
oqyfeW1hTAlLPi6AMuL798AJ4yMAbyPMljEX4DbrU0eX63c33ehYdpWxo69sQ8E5
FnYBw3qPcEJeZdq+2Cz1giXtycgBAjbqWKnk3O0PvRdrHVGOj5odDLeFs4f0xBV1
SLpdr2EoIUks1DoUL9k4fmLe/WIlsHHi4yiucSWt1s4xGS14e9UBHzsNr+SbuAXy
LWdY4bw1QMM1hUzSD9zdlT0o5R0d/Me4muS8gz0bR1acbZCdWsAEjQ14qZI07pm4
ljrqm6ROXxKfEZbv3n67PTYbOTaF3lcn61llB398A9cuyfDbfSl4/yCWDweRALTy
ywCkJsDwV9VunN33qZQDSefhCDgI0beJVNNocCd6/IX4VnqYyveXo7VIWslc5fVn
T4GTBUXJHhCHZBbRvwM1dtHQGXrxbUhKFR88Ak/QDcxvt+pgZUMuDvdo9ape5XJb
iLRqN26gdXqi/1NrSbSFCU+iTsnbEv7HfDjSs+mkGTjBm3mlUnsbO3Q8Na5cgB4H
NkCnEcSwxT0ZB3RrXtXyo1dGvFqMlA8H1oUlpFqMnk/Wcd46gp+xzgAE0Rc7Hr2N
AQjcl4jrVpvtmywUmI/HjoyX4lZ6/b2nvvfA0qFJrvFCSEMgIuCCPY+gv5n1ThXD
9apstIQrnn4kgdjBIwVeyuMgmmLnJ6yMLo60J85Gd6x3f3yI1cZuA8sZ+R4TgTWN
+2BSo6dxyVvO6H75/A3UoMx/3Eh1fjREA40MM+4PLwo8cJ/ZpvUMq9a9D1rf7p1Y
rzVeNPEuvxtvfl1IJDBcs2p/SGCMFRXm2R92bfmwJlaQuuCcqFAm+gQwd6wwBAou
mLy0udgqXva2EExv88wahtByh3fvi3k10FPiPFe/4rxTZunkKneihoDOBWI+7OvE
B3OZdMAWZfY6dL7Y/IaOYxBszxqO1NP7/+D9jet9IvQfqCr6j6eOSmALbAGQ2mv3
jwW0CW92f1MUZF1+bnerApl2eNCZpBcLQA9Ylxl1st3ckEUixK/3WwOPqIxGicWU
L6YR1WofcH9SHIJLwv0cMCUV76BYA84W3D2/ZqxdDhsgMXTS6thT1T+t9bj1W6DD
zcVqJ5covjcFCrcPTnLbzKbkeY7seCmJxE8PayCBDLs+WUTC6QcMRYUa5histP+1
+rpuHd7TP1hF774DU7F104+lnVS5qe1BJ/eRJqODaLmEbFfhZ0OuaMM6DTsX2YN4
RmfsheO1jx8yqLyJWKvSqENoXyob0N0s3kLW2uxJme+UwcFelptnSvWoA55GHpxt
jddrayoEuwWF4N3KPbnKixuFwCye9Dnj3Q5IOv1Ge0GtdTmg2xytAWuGfElvIrt8
Bo+kBF+2JH/tEhyv+x+ZmEWBR4OhUq02jFz15uUiB8lVIVtATi6NN0mXzOEcS0Gx
3Wbsykv/FNKd2FGvImvXnqSJ34R87ASI3ItUD/F0KPZ1kNXX1q4jYGnCo0DTJD5N
/xJW2NI78jk7J04ZjHzEnNrMW5CC8QPVVDOzsmyLJt0PYHs0Y+mWrdY9HTIgf1aC
f4j7youeDtsGqCdkOKjAyD0dI8HSxY5aQRgRt4FwMc2vEAUFNzyUPfuc9srp8QwY
GvdrTc2FMH83zhCSPguTMPLy30fdOiznbcGTaQl/pX4NZeZEZglP1C77AaEUejgv
MVmU+NaMqLdry1a/GHehKn8h9g+lKKXXM1ItSwOpYmBxLtkkjVjrOKaxgiqLySpe
Rehju4E1R7/PTTMh1x3brfJaLwy9ZwbijXvgnNinm+dyRJNbEoULCTtmt6133DbX
lG7pbXGfLDKcBKmP2swt0bkczPG/3XAHXNq6PUQ2Xrf2cn3oWg/qdxGz1CtAt2Rf
rjw2SIPyRvbSjkjwBoorV6lhLXtKDdkCJtMEiEnKGz/oKbVjNeignsOq3xODrdGh
ADN3e4cgU0bNB7oHyESRkxLaSKlLkpSgDGy3VuZPfaDSfve/ZtfoHzp1uh0kd/Zf
kNjBttH1nv+K/aPKpn55XiSDuHvuUajhyg30hLYKvS0NXThDionqgumfx1yfJEPN
RZ834qEpZSd7Wy7B22nwfDFkZGuKFAbAP8FQGxBz44r1ovVo8cvnXlWDc0jPKnKa
0RcqhXNdI0KOrRj4vD1OHhZvqhyvaZY0hUG5zsYQrZsElr66cu2AKD2d+2jIg96X
yyu7bqm0QYYdHjtdGstWdvi8T/DfGXHrrx96NuTDfM6BCg7XyMu3FnG38QmzlYQJ
rHqqYTOAjcSR9KDWhC4fH6P5bgSy8FOqvahSnXfKYcJqelOP4YuLnmKc+9BmBUr9
PYwiFb9zTowOyr13xrCFRzhdCwk+D1c6x6oahJ7XDr978IPAcBJMMMpKqLU0e9ES
dx9hXbJdtNzkpqX3C32ckm6BgajxlbEKuV09APBa35ddw8hny5iBsIH9QwrlZw8i
6wbH3XLJBWkEB7Bc6IOxjWDEVehMsIDQZQ1JsEyPy0CNQyAjs8v+jxIXieZQqZYl
rvApbyrEWL1ST7oULHQEpAY1lExjlwzLmKvVu4p7lwKKyO8UqJTiGGAl9T5MEw+Y
t7gfVWj7GMUFYLwWJdC53r39LcHjJ9CvZ3Ekz6uUv9j022i9TPtzpcx4TZ6cQCX1
Nb1Q/+QE0SVcu4h20R8iGik1e9nF6AvmG3Rh1ZiBGPQ4HcirrW1/SCOp00Wy5kL6
25oaHhiRidQqXOM3RMJNqhDAwpGAl3MNm3yCUeWEZKi1LsdCNqjpAbuqZp6enNGG
gRs+enMWZPyKLuhIx3QXc+jeVla2ZQCagZxSKb0vimubR/3J1HfSYA8BC4VmJaN4
D4zcUEB4xc6F0FP6zx2eKlYSgDVQ3vU2ZBrKNll2rVumUlHObYUBFTuNc0cLO+rK
NBZOD0KhdBlHMeh2TojY0dgZkcqoHqIhp1wCN4RapP3Fcy2bac2qeSfRLNLDn8Zn
CnyXdT00GTDLBrffqB24Dieba5QhaWd9jmZfc9C6P2sTDXtB8+mI0gx8wh1sdLX4
GMOEE1i0cW17JLVTFZFqHQZxhe6FLBssF/pLKvg1PwLgFlS/x/8FU6zMZ1YS8QlR
tGmvtrCk3zTsp9gltskLLdYf9bTS1QfjKADo1FAo0kv1uwbClMwTszB/lgJI99Cl
Zb8Qt0Jsi51gAFsaAnT4MkeLS4aWAYIG8iFBJyDQ4n1GDevldTp80wmrLnv22TEP
ZhP2fSej7ssfH+HZqp6FixFsw1CS/gCySkzJ9HnRvlqo9dK8I6CJsBVLNELEJjPv
0+KJTQ1maU5GDGOdmGzY532kKl5jz9SPYO5EwbxAHT/WpsQ7G8v1hJUwKuB89CYz
3k4Y1Q/11O7iKuU9L9VH3GoAkG39+b33ihrX0PlWjMexscYZBQ6nDjBJrKio5qIq
Z6ak2A8jkGKFYn4kM0VgG55RR2h3bKKPPDl39iNxFjwMqQWm7F6AZjaoIU+mh/Ia
isu1Ge0ShoYiYA/qCHTD6J8KKmZQTpWsbxwV6mRwv4WUF6N8Aazas6Wt2+qXYu8W
z9zkTH1XQ6M91nLnBvjFLRxebY20CgfJvKe07tuJ0j6VVocDjqVeBkkr0iJt5eQ0
g6BmDmDXs/+fMl7EDClY9kCK3NbcnkSkGyvZ9cy3lK88C4f99pquaa4mMCBWYdna
QI7tGlsKgTc6RfnkJGrJqgOr/6upfJwkSZfF/72+Eq7Lpi5+DEXxPFYFyl07PLOj
gxOT1e9RXwxcX1d042xaTHfZzjG1J7k0XmnDfxES3rbcKHyQZoEhrJH5oIkWnxJ1
zp6sU85alyZ4/RToj+H/EOCsYOO4DdWiVOIOv0mvFews3u3g2GXM/pPj/1SO8vXu
EeQYUZ8HWiMnFRzelRrBQvIXaxoLtokUqO9NHeZ3oiderZsf43E1qP79kTIP5p5C
lFBJzgVec8hr/mshN0Ta/kmUdahBykE8QeypXEGGI4N3+K2S7g7A6iLxHORT04iG
muAy1fXKaQDhHzcMz8LHsObyhxheXBRPBJnENw9IaqVSUI1t3eeCWZPJkJFZzDWb
Uyx268BMZUDNN7xVPdfy0V/qxBelU46rdk1AQsQYoMvy/HruyvcvnjIYpkkTD3E8
r8TI8KDRLDTyj4plTG55jCdiJNrsBPThEqUvkPMVvokf4nJP2nKTckZyIWFjctDH
KqPZdEH5xF//c7vXiP8ua/FTHnZX6aWqqwWtxuckDK0sFot0Z6P/xSw4h5Jt7810
vaEAT5NPJjatHd/Xd+gjU+ugkD6B1hIJffgSez3En2eROdCpQyXPpQWit77Qrj5z
LlcibMNShq/8cflRXfKTHG9gpEg/Xl2D24re11ixjwCAl5FIYT3YRjJMsGJruQYt
aRMI0Sq0uQUbhzCEOHoDrNJGtgZWlKYcX+SL3AwjOYSkAfnheLEoBSgA9Od6YwCm
/tD5JgV0gYDXG41c/vCjNtWR40dcDAY/fLW+67/ZFXXK5MxC8GMLih8UKA6pYbkX
+iiaqv3rrQIEnWPeN3orP/8EcFYEDFiltFzwn9WJnXVH7FQwNWuu8bjQgurIIt65
Uje1CWu6rC5I0T+ulXxW3NSj406kmCGmqUS/iTjJ1+8arzjv8Qo4NUrI+2OCTup9
pg86/98+Vui76pFqq/kf+k/6Pe0d5gjKoFdiFA5leK36G4pvUg10Z10J6c1x9RVT
Sm+6LdTnqJtqk8ZrLxlRMMOfIFcWw6+ccO6ormEPAHQusxS5vL6GTvrdeGRFlnwV
J3sv5uLLndI9M0g9POE6pLuwAR99LUw3oMEKmSwr8TsnHb6JBsF6w0vriKBZpgyd
Iazm/HbDuuGYo6iopQCiH4VvzMyAhnSMaBUs7TsStjvEO9299xRdrE9Ic067KqGy
91aHN4205Jv3uzhoyXZSjY91pLffS1aAWhbZpp6lxuHrr6A+qmyEHiaRrfDLM2N3
xMK2CKF8a1JT4DamOWpH1UtHKpVyaIYFf1UzZJe0+VcWKDToRr2z2csHX3xCOhsz
fyntDCMzuySMkKWhZ3O4fdpynswYz9gryvNFPrAspYt3IAgw3Rqub6XDt2ko6MNM
18JvSeRSt7wCrNk0n1gGJHJ6TNtSEHrxs2FE1/T5D+n0aS4/0/DT5h60hQIMDF+U
UDwbLvqKDk4oC6Sxi1PUs9xr4ZnEGzl8ifN2gKav9aWhiii8OXLrUkc6CFqxBWQn
7cGmmf3G4NGcw6553fb8dILPxM5yahAlV9plfXpFLWHzZiozpvXeJiyNv3ykZ7UJ
tR51Vb5butqbcssiBUXBCuC4grNSN572GrA5rDZ/e6ce9dORXfAfB6jsNlsh+Tf4
Hyx0gI9Hy4YBjxl9AmnnRr4y8Q3u1B664DkgwfxH6Cy1P+NJVHXvccz4uQoqfD2U
TbpfRE+BDtzdXbCtaNtqhpRiKxpU02vSoSAuKr0Fo1jCfnNFpqktEK3T7srJYXF4
fa0KTBR3InqTE5TSijmF5bJx/G185mN9sqwAmzWQla56kNwITKyBu4mmxwbfhaiP
EaBKMOJVKIsIdRHXsdJdJLDiJ/Sejj9Up1BlmndSSBwJfggqCVCI1Kmkj0nUVbPX
iZtN0Gb1HNaejihtZbxi4the/aqkV6eX5+HgmXafd/TV/hjDkZyTtqXm6oppM6Wp
Ca2kwCdj0WC/Lg7BohzQACU9sEVamnzHwc9tTQmyuo/ujOV1tZZzN+hByQ1IyfQE
/2mB7aUjy1hUWrVIxfzi26Fg/TFypvgVW/ZRrE2ClDgnxOzpS8dmo8V22y20mS5g
r4asOZeuGw8PO8+0K7RNhtjoBinOdc3sixu2DHJXmN/t0r0w05J8Loqu/DlSB7ng
lxPEi0+/IAGRqwVQ/++s+nmB6Hmwu85GeY7HQTHjz77GKziAquqUlHNvsSRuwx8F
n3C/xxg/Lg1WqhRq+ilXvIeCgAJH2XaMztr8XyheGiuzj0vH+1ZVPggBC47hMiuv
edYaKSEuj/VIIFKrbw7VKpUD1l9xM+o5ajPwILKgTX8TjnnBjjVfpW9Wcyh4drfM
pT9gyRBEJZMmQ1C8zriVRALnlpdflcU3LaU0/+SWg0tR7EWoG8rvWwBFib+Kw3Mz
VUcJP1FFn+jRSzf9Z0L4ZwIo2TOvSkMP3FC2glMaSx+iWp9jZ8eZzxrJDMgf3hMX
Lb7MwYY1EWGfazuBcurZka0BLB5Sd/wdvEYLn8IFTpwOjrt0P+fy/N/cFOVuAQnR
kdRj7EFEElYHRA6lWpR/CL9ssyRo9IhdhVcSkLMHstLA9vz76ROANjAJ+FugXYei
/D3Ds8ZtWBYgi5pRV20Z4GFuISUAzxHwltqLXLVZxAYlFp7/pITQcufdbmW3SYRN
1hR/rwMQJ8/1Q8FrOlxujlJtskGGNoKoq4arznNKeiLx1knexvOq9A0h4XetInJa
5XM9mVikTECQOtdolB1lcuKjyp0ttc2MNKbVc3ohZn8MHxKQqz2cCDjysMV2zson
9KTQ3reHbsMQG1JdfCqoj4P7rWxhyjMi2wpGXFWxQpnCPMo3vChAj1ouyQM1R9O2
vsA0ZzwelDIfwX6jY7+lQKhQunqz1wEWTollSi3R02wdG46eXMQv9LiUcoCkKNUO
BTkFm77E1Is45zvmnNFik1bqdEQUP9LBVlimPLJWRv6wZLysY+pzyGLVdlkL4eL2
v2Cou6W/NyTaHKI5z1shw32zzV2eHeIoPwX0ddjcEfI/zsdXeO2WjzLXp5yd/FyT
RQzqYSGxWdOM4b/8k9nzZbHWugUHfJMm5ZzC2jjqo09n0IDNaY7lHsPqhKPETcwU
CxoJ9ruLmKaOebHCkRlB6U3ETFCFzWET4O4J09lbpLRr2da0fejpMx2nhAJEFSWB
jzCglqHak5/JejKc5tpANEZqAYUT3AeS2p9ONF14I7k+op1hCkTYGSXKWNUzVNhT
KBK0XQ9Owk1Hwe6u7qXnf3h1nKMnSqpCgmSfbAUHL0D5zms24oYo2q0TaeurY019
Rq+AmNo9bE9/EVWb4qzN62j6Xhq43ikRoMPck+FYW7l3WnTW0/Xo6akMKdfWhqFu
lpeizGxqoZTjTAiAwxOak9dJXG68C2Ph1NLnZmiRDGVUznFrNVgTyrTcVDX1T5gK
1KMyfXCZVmJCqyCFSthl2uU7al+hKjDeGPrKyes2loPwYE5/yfhJXrDIZ9Wa2hGy
eqKIjopv0c/PylXX0A7hvXGOOVlhqjE1F1m9jUHdnzKVmwj4DvbMbit7qj9F2uKj
rh4Nuw2ms3F+jCIXkfm7uNgGWx8SAdShzvfuF/ZI/UAH1bip+fP5ff2i+7T0XKRT
ydQN8+SedPfMxzZ5pBTXzD8Hh+OBbwGkikVMfXlBuXxytuGTCKidnOT1t6QkaILj
8ORqRsFf1gLF7KsUvbXLL7PTHqiP66VspZ6ffit+cpcHfYA8Z3Z2Ae4W/vjPK+tl
F4qzwSqC/Ks6lkDrgJJ8RC/f7pvyU5mMnIB7+r/Pl8Z8pCcAKxq56bTEKY9JGk0i
cRNgmQDQj04oLdcMRFQ9SUmcWTSXMy9vEmfV/ZiaIhoqf/9EmwJ0bF0rgnU5phXW
0k9k8+kTDzU0+e9XgYmmz6zYGEO9UXFkk2UyExNXjVFfb7d/ZnX7Qw9MURHbFv+f
LZ3LMNxwa30oQKBKef7sCBTk+pMmuT+h7764VahfLZCMWvTcvpEJa2IVSOsrl90I
EWGnq/4c/rmTuGPMlFdgJNIu+xdtX4/oAOLWY7YvcHiRbA2y3Ik4gUV3p9IUC6ro
ZYUX6VjaLPb+NoVl0EDGbvOq21eVVtBWRuZlqJLhfZvhXlwfN5jSbwKqIGeUbQPZ
AFDp/akg3RHZD7sET00VuxL+AGvd3DqwDunNuziq9vnWG8N6DFqMdV1j7sLBPLzC
Fv6r2N+FJyzrsrgcpRePz9V8gl+pZBg91i8Um0WLMsIhNuVRjoFd8nujKA1GP9Pc
J+1rl6/TmCX2ekLLWyMM0IHXhlhpT3EcMCrPfVF0/98WNoObrhEqkkBk1QUGPaDi
iw7bHL4psxHsZTpbhbNjUQxcLuJD6ToCeo7zbe3wzB0L8V8CzYx4iXapzMIHVqRH
2EXh/h4euCNOdQoxVmhAHjiciQwHoK7HCNsOJ5RwDgmMG9cVukmmoAu00PrvueVn
tRzUpLslw9ZBcLMo3QSBLdD7ALNy6jDwFDDXjhhytc5mIZSG7ZALl5BTdC6/gHIU
Rai7aMsdO7Oofy0mv5fB562LIhDxz/wFWbY/74EnD2BUj+75NpSEYw91qI3uk5rp
DaOxbtC+zv8TYXfJtLTtHx6FSNB9RK0Ezzao9zcr68KQEmlYvsgGRgdnFKXIwiW0
HKOS7DIPmHfG2vGt+ie9f+SHwoGFCP8+T+N9fqfcnsxZ+pCbUU1T92f5U8gtyjbI
4NYMbZvZpryAKiUjipeYJhUObrbo0iI9mgmWNI4Y+Exr0QxD2P0r1MwGlG/CU7A1
s3IlsNt4FwrhGoqPAVVSI5zi9mfxp255SEeZ+P6hTrqqcd6JYs4FhxZZgZzbIEJ4
VFl2Ig4zwbo7JWPWIzXvsRBc0yXKv5cuYyAbJUCa8PdYSaB+9j9FjCUXP41cKuIK
+q8uAbhMcFL6/hW7aSa42+14oSFejvgWxmzdGGWIye/OnMfss2I1FJ70EuTe8mzb
iYaBK1nDfBrs88bfO1j3xpuwwj2GjaoYosa0aRwWzG3Z5vRUjtdaV+rjn8Tv0bX6
8Htywwje5xc8x+zOzRkkKHHkCKbQU8uEQMb2wcrS+L6CllTuaYJ4bYbldvuGbDn9
FqGYa4QAjfjCzR9mrwPrmkkZeiJ8Ueqc2Vy9rcYI7EMQh9li5bhYjBmOE81a7uam
qzThAw2p6QZOXFctK/nP95Wa0ms8cBAedCIrP8XAtpK2yJsRho5aeiqqHFuoaJ1E
XbYFjLLAIRt6KhvvgIBXYcxCfmQx9tfUcLW5RD4EbXxP7AGcg1a7p5CAg2832MDm
TmxbeUyKmeFTuqmE+sY2AHs3Op6eMcySDtTbg+yStIKqCPk6QjR1EFeAMKXrxhbB
idtiAUQTs3r4CV7RDi0YUlF2vF+XDJShmXySLR2bZxqpWAqA/IbWQ2ri1KfT5+uE
c5Nve9757Drc942PkU5BhAKrM6Npm1reebIhIWKp6MBvjCePmFxkcV7FkrcBCquc
+E8Ri6DXA8E89EaZFSb7sjbTztZNEfuNOQQJ5dcqp9hR5lqnmN83RW2kKku4DFll
4iiztQXVf4ikWiZf4tN3kLOVuFHVqc9DVYzyh0XmMPo3IB5P6lBD84mG8Zw1i+6o
DLUSeIzLjTuONMVh1/qZhXA5Y6gJCbl9E1YAp+RHUOsIY3M9djXDdNYpMbygb2z0
Nh9piaYpGO3lireopkwBGJM4/7PTyMX57It9gmsplnU2V2bWluQdlUoXgU+kA2UC
xpIM5eOg1Osd+tnp7g7Q3VC8OYXrdLPvTUP+KQfBRRDEy6vPfdqpgV5mJhZyRrMy
QC2b9EnSNlcf5U4xu12kiKQGFUHp56fT0NjjgF8Hmvz+8DTKTJPqbMllFD+RIol0
vSrOb6Cs2j6oJv6f1IjkIASYe48LYXH0jWmQTolMVhM8yJ2Qe4Th75qaKlpoUyRi
BUe+Adydygp5CdIz29l7hpxZcrLT/X2WuG0NXnSJfPi9P3oz+rZQ4qbsW22vRF4K
7z6v2dHSWXjEzCbsaxyXA8CvZOl/oFwJestAtK/Xggw6QatkylrxbA3+GTeMngBv
PkBmweZ3CjZPFHjmbHiy9A5NrRNtA4lt1RUAIVRhrj1ykvknPUZbay26YgL5O3B0
+AwZb9F1q0fuEMNz/OyCvzvO/Ull6d0hjbG8AXXSCSby7r4re74IF5zo4MHUl8MT
Aofyk8T+l9BryhZVX9t/D8eggvHpybNM5uShyvpTEmkZ63QBwAxUk7111TtkpvGv
kbCXH9jhYwFhdoYFuIUxrE+9ES4eCizi7+Z+6CvWNE73p9EfOj1S3E8ZVTgtbheR
cFg/k0uU+8JLQ7ftxn+0SEu+Bzv7aMPuTlLFXrxesuLd3Tr+NjsUuUg30gj5gkAM
pkl72LuETxPYg94HSlweoEisBxmkf/nFVcCpVOmPvpB6N777MrWHKPU16g8+erdH
kSWzTG/TpaMjtC9pvSxJzIrsrMawViTQDDKG6/tOAmx7t40N/7Je72uPvqz8wKq9
aTdg6ONaOxowlRZhwrNomHKjnuDbVS+9IROdIajMWO/iPXvCt8BnGW35saVnntk6
dOfKWAbta8EW7AW5B1+XnCBXIDwu1UsSB5CPckk+uz0z0dTzkrOIGFo17kOgenCM
U7cz5Okv1G8wQ6XVpFh8a2srZJS6fx76M0KX3n3BqN8lE7wUKQfk0Z26dA5DKBeo
qgn/uFKcRNj1oCJd7jsQ2X+iQkOZk/o7MJnfHQk5j1uml71OCludOddMBoOpWQnT
gdCUOMYxP1J3wb4EnvbmJcZ9a8fHIP5hc8F5u0J1PUPxc9hpq+0sfNdd3KtxBipF
I5UZfdRo9fbeRkBHvMCpFmCGG0ckaQlsIbFvThiiDpWDpAWNKzp40i/MTHXsV4hN
aGglSCqDCIcb5hL0IiCQ4HSX2692JBzD1aqwIzPNyKG3383m+LAuItAb/b0qBoEv
Tt8h5dp8L1ufuBKYZtOxZePHtTMIKA1vW1v4Mr9X9nRQtwFmieKEXuE92U6mmnvm
9kj0wI9vHxZF6n45lD722WthIQg/PqFwo1x1NPYIiH/HxMGF7y2vAA8Z8f83Qn79
+xC/OnJncTtmjLe5gKEe9LdfjIjZeEpt+ZKSu7bWTYi2Vs09INxPhjoFUl0Ox0Pu
3nBFNgZf2QEHzF0M7lAzrV08D2/vDBANUZzrvE2AVx9y6lAxIuiYuHVtMHDKc2xz
urmJGR0gvakQisW19fdL9Am1NfIzqQ00RVWW5AujRnYEZYQ05rulJJl/o53unler
Kr+U1y2vhsmXC/1boLH0z/MY+PbWnsbjqqpZ1rQv0doz2HfrhyuA3GhPDbtBDG/e
5JQ7cReyAviLoXVCrbGpFxCSsLqukQdS78gkGsq6UDsKdvV2zKsOev3i0Ybu6Bi1
x559q7mWyTZ6PQ+5UwLfilxIe/Bnvb/i7CvdP8l5fGiGjTflZPfap4jwnbx1feig
ZYdSB139WiVD3zWeUYWwo1w3UMwf0nmQ6eyvKVMzpnXSzzAECLlg760YQlkLKerV
OrgZxNhwuPEU8oLtvonWarRxXdmYVGVIiwOsEKgI4A5v8vwDM7jTOts9Nd+U4FLb
RGIlMyPV1fzsxKqJ58vhDj3P5XtY1DghpxjMG3kBbcCLlP1kXYIbugDZpulteLRu
zeEZFbgyAuMZxlOVgr8AATIc9kQP6USwoGIthSDRmOmE3eufnIk07UbHr5toyycN
jHcHMl5S5F6Z34dW2rkpoKGNSbJP9CWb4hcwvqvNm9JGJ5FEAbB7giCwCchMJaRM
qLULd2H/Im+kz4VzRp8IR/6j2hjOZ0UmPEulWyGvQGzBK2jstsNQ8tYC7HRN7HJu
kD5b6bizmAPb/TJBebb7TzuuAMKFk9ljl2ZIU0YGhbwlobgoDS2l2NlhfIV0niSd
D4zCy71HAk3kh/yq1oCGLN8ilS/qKvWW/y7hlxexO+v8ft/XgRxHqrxONdc5Adw3
WEimL1WmbZ/63jJDmWzUaVzAgeLJgbbFZuI3le0rA9H3ZV0tJqZKeY9/pB1srWe4
jLPfzFHoxDwUCfwGbMtYowPnMEsq0TSsnWm4s2DGu2iaet5FOeymBrBWEbYmoQCe
IQD3CnC7p4OmSU0cvLWKE5HcaNV69yOkT0MjRw04qlVxe9feozwUjGybVH6lINKx
62EXfIt8dcePrEHr/nMe8bXuGKhfN8wR4WemTG37eWjXkWDgo+0LxE0qOt6lVJh7
bg8lfLLcoY60AUvb3/JunFIkKPauVic3LGjANrydGikJWVot8zE+Fop+G13G352L
BlJXXSr4hO0GPpxJAqGGAFOWiWjPrXb+Rf3iadv11FGEgxdecE2ccis3HmP0ts73
z6L/rqPLdAj6f10PBuofeRl9HPoAI5l69e2XsIws0HsVNU2uJePNo1sAm1PnkOZo
mmeCq3LhaAlPDG+aT1H7FvDEKu9OgWnEqIofnikHo5SkAlIKqeLpQZfGe2dx/cYJ
Z+27A8wUKjQot+mjp/Bosk9mOrx+S3U09ocJgCa/AAiwkpY5SzZQ7XAuRjJKV0ju
5e1HOGDkQnpy7FGpBsnbJDYw5SaxMhB2Vj8DJIRBncgQCfSeWZL/eOl5b9Gbs8y+
amZvpj14+ZGXo9nU4XNmdO2Q09FD6ii4p1jQHl5K/I+hR7U2VnKeWsYwnm7vn0Wz
DVVE1qQt4MylK624iKyXZ9JTbi1ZdguPsgendJVZNXwWx8pEOBzvEaxRvVtHD3iC
xHKyMnLRUk4FZwCEpFb/ktR3hBEPE2Gf3ocOaN+CQtRKfhum4aTwS/Om7yqlaq4e
889ufHtZWVuaAdTc3FvHy2v59lHwntIyCYCCVVqMP894FHTUZwCaPPdOdjhRlJkF
Vzsfw1fCd9JrjpKRv634NvVUN5qavMo2ZgK//6Tiokzvn3Ho2mORHbnZTAfEPYjv
EoNfDah9+P44M6pbdRT5jnzUddyVcoBXwxwV0bsPPyfHd/AmmJzmYiFDggdDAxvn
Xk7AllpaB93AkrQGAqLil2VvkPgxyB8rh04z9t6DwWU4CB32pTwKT8VdduSAhGOM
beGAvsVQYLSX997v7E/fvJuow+F0p98PZ9tjAGjttyPmXfSAzfVdzianGFMHqfSW
e0ZIQ5EWbkQwbTkpkiGGWf90or31aUsstzohKxyw5vABEU9mMA1cmqqSw3H/Yz5z
5OP87+cgIVbPTlhdVw3jb+50dVa3Q2Oz2eSnGSYiFic4UhEdxYAvsvoR+d3IUiP4
mUvvQNxmVBXioPlvn22srzPZpnz8NEdpSvJV4hawBsJ0bdIOckvyV2N5n8lDwnvq
lzUzs5ID9NxTANMv539zBsGJAO5pyECGXJKV0vbEHWj5DabqvA053zD0GqC8ur1t
CQgojOdq5wXZheTePk3EKHg9fHiyNdgDbMg2yxPun6b40oaqCah2Wem3/sTjK/My
rJ23eGNlYqE8dIF43ThvghLD0ChGH7UHMjjxz4ijj2snnTtJ2jcKH5Q2dvUSDvrs
ISkW/gS18ibaIu6sPwTTOaLI8F1/+cIP7fLi8ZXmI9/t77IpXleR82MXpgXOu7bQ
dckCa4QQinR6O2M/K/oNPN6yEOI2EdhmvNtBrKpVZZBaUjCNSTlL/8o5Q/0Xg6o4
hjEBUxmXOCEXtByjtYQXcQdG8lgoIVEPvDv1SCauwbO08m+jXQfwEKtBPBGQIO7V
InofaRg2O0vV/Jp766lSUtsrDV8q0zkXkfhd4ALWWYfgT/FTsmlNTzBG41yf6D0v
+ywMrtoLmI4kZaBTzi+ajkoHNATtVZnyRC9kCDWYt0tM7ENkcAQzO+o/bIqiJFLN
AigDNyPri5p/rBv5nAqwlMQsEmE8ZhbE0dNHSswcDp9bv1qaVKJjhZae1kuSE/Fm
OXR+BAG2PGGsA6tmT49lX5rb394oyHeLcd2pNpGdBGgMLvtBq8ziCiPhafNfcaw5
BAySe+YPcS0cEd9i20zEzwODKJvwqJAeN4XZWDqaMpt7TRQ7JBgK0ha7OVuJQLg/
n+4aGv7m2lpPV5hZSF+R2yGOib5lDGmXnbZu1N77veBCq9bsGHm+OYJpHbvnu1rn
ufMx3e+W0hYOdviecI+KY5Kw6bKyp77XLDgHi3rS1AKE5BTwBDPfCp6rWz2WXZc6
zNoWrIx1wpH/j5mVkCNFJFtcwL6U9NXCvko3rFQ8S7Qj1VtcQWXgiXumVO/YtsHo
FiJaE+Okm/6nMJRRX6L3x55x1lHH5K/8ZcCwh9fT6t5u2uUPFe2Px3MKSXNWVDKW
Mn4tVhgKCWnJuCVLlk6JcChFat3kEpmr2S9FDpyMjPoSYDGVcOCE2OXFSfwgoh8J
82G769xkh8uoxzzly6oJAOF5XAuJ8xxki+OhwnKemqLI+LztZsH+mD3eG90E2m2K
ygADHsAViEBZiOuY7ODHwDwTeKnGLd6oj7egskCleqAWoFQuKE49aUMUBsbNZCkT
DtxYguhc4kV8Q/g/SZ90cUdLhYaftJzim1a94CC9rj2gVjtFAzwTBuUAzLcA44lC
h1L8h5nof4aQJt+82d0jJV3Ebj5t+mJKW4eEmc5QfrzxXac9QpMpcUNCwyfmVPtC
0T5WHZRR2VcFiAZ8SK6Qd5gFddVkalfH1T49+y4oT5Ovq424aK/1hSkK1CSazqqA
BOA/25lAsXQSXU6cTSNaJdYRhMqIuK5H3o+CXbGHeFGypgv/0645UN6OmzM/3MPf
cqj35RKYj3NA3rFpa3oacyvEGVC9OhFt8eUonD+7mD685P1w+SzCN1jN5c2HvMM3
zaYxBybDNx3tJnW6bmQwRlT3fmt3jCNEMwipmizRDBeWH8IDGfnH4mrEw+SSwkT6
jVMrntclgDXQKDKSRVtiGMuoYQTgKWMEF9/7nKwrcKxwb4lmWt0TGBbYNBeGp8lj
Bgz1o3sj9P2XWLu661YMgp362wQoOjCmf5chUDH+9yl4tIZs3m5pyYweErcfVLd5
6kG0nN3T4zDelZagNKArjPvEAWZ1d5JRM7U84yokvLPp7aUzOCumIMoe0Hgj3C33
A3qX+QtT2BE+bbXKvW35c0GRUvOCg6EVePU8L9GwGvgWKFmg4ZmjcN7RCBVSIYPq
C6o1rU0pSNIG/U7HbALWJS8VP2TiBQIOUNWXaUUoerQWxBd7geK031c0yCI1tKRc
Kdg+Jp0FUwVtUNfVHM1Ox9RA5c+lCOSfQMhrA3YFiyc7CeEL/4fOytokwWma9/6Z
EBOBzoYUqosDAP5jb16nB2JjQr6LS31fdnxVP4Nu1Jqt4NGLkKVGo3eZzgOyFcoL
M/n/zsH3UfPxv4RYrw22/Pg75UxPSA00kKp1YmQJKYVSEbFF+3yfxAVhUdvslI7l
blrGSihRTU1FHWmcKllpLNeDZWo74e5QWYYPwatff0anqZsc9lyGophLG15L275Z
pkUxyHFALkj48QNgAf20gk5hUX9ZKLNYe4DtYt63hE8hjI7GG5m71h4FCk20sR5P
6aDu06fZDUmxblIQsaVDw1W3ilW73nD5MSDC819aKb3KZhv1EZRnunpXzEoYesjM
p8qOEdBFihXg193WACX1CNFOw6TFXJK+32SOlHE+NI/L9vHu9c6EEjoigfhS46HR
c85Hsxw0inSpWHtUzw8L01IaTQiRkh/J3SJfmksvsVvQkjrgkeOR3dyizD6fHt7J
po0CTPFNnDvPKZO6akfNXDs/cnzhV5/CP5DhH5Fhbyz4e2nl3/ZCF6+hj64W8CI2
jVe5yMN5FhJVsMO5RcV4Ft7Bf2p2zob4ZEvVq6q9r9TR6rP+uSmxeGLIfNxSBYUG
6/IduM2hU4sBMX6zo78E25GGrzOtp590jyDATS7gCme3eqeAx/raVTiwNQpUgwYu
9j7RrhmyYdJKHrgQdlzJppkJ11KCo7zoLIHjwanw/T05Lkw822JGzeIsnern2FFO
LUWC454OcGqSbnhCdYwe+UM9FcKy8FTyJvq+CiTND4B8eAthoqqnh1kMNiNB3IP7
DEkbvjSeGVEYIChtZdNOgB38G52rdSGrs+bX4FimRI6HHRhGP7ziN92VkyrdVrTK
CfJR+KwcgLcla7mgHQ54nsBSRtXdB945TZZyyLw7hje/rCcrU17Jkd2WttzSEAxb
lZVWTW5tOu/KV46/+Fn2rl0G+0LhTXRfGFe6xDiOQm8RsOnqHH6SLEpUsKwBNs0z
oDYewQ2Juv2Ejs2asOUJQZxTEcBRzFmEWFTeX75WyDXRprvV/5ETT4lEDdeLg4ec
1//XiNjx4bT3p3U78AYotu2oKNUmSVfQaj254df8A75GsXn3uMQxBh9xqei911IM
IzmJlwpDn/oB4ikRl61t2g+jhUaFVG7CHx0gvi5W02CqlmX945MNeoDco5u2NHcq
c4Ef5nV7/lw3nYpaeld0f8AQEQJlYG500YSA+8wz4lr70JiT96oSgBfncNPult93
n4iwnb4x9pOqNZQqGZ1nXwQDCBYp1q/dfs7ymmaCZXB9iYGITREQTfFXBEs1O/0X
QvHA+X/pSNacsy3JSNazyQDZI2i1Q6/N00kHoffpTeCcUF3vdr2ZmooSdtqtUXsI
6ohfZLJENBYB33J1olc1c9V6GnAy75Dql4FWaPXG/B3IiCVSqNffpCJSwmgujmp+
jzBE4BqcBxIDsg9QBo5MQ3o1upLfaYaW2O09yKa6H+eEWMoDOhV92Y6T5SVjgoNU
whAjWt2ZX0F9m/67aoweMWry7SONH7pSHnaUDbKT3kuzDVW/Obgo//iC6OHVJxsb
F97KaoTvL5Y3fvkDQxdGyikny1EJ29MEPGNzsGzw8QOTN08T2k9dcJac0L2xP4FJ
zXV7xt0L50LQ5xvaC76k1Ul08uDCbQsEf9Y/eLC2pDVc1/Ms9G5ddEw5X1SleGRw
MvXy+ihf5q/ngHflUZdJs+NqAjkx0SYhJJ9PL/HZVyRAvdOod/jRwPOwLQPFJtLX
icMhS71Xn6PowXSIDuKSRoHHdSBbkwA8g5Hf8xYYeQRxqFcxn6lzO/UVgi3wroe/
gznXh/qW1ZfRXEs+ZZW8Y5lPGXgQHP5RmgdbSwnTPdF7FtkOjKBfkpfWvQUIA70e
K/RflxN4ryRSp+lE//nHHjIViGLyU5YFMl443KIjn8ubeGsjZl5c94GFr4acTfby
Meb6KS6iOAwnnJXB/6AT+5iXEhxFyUGupkrCQYOnwlywDd8IeH6ke3M12c1eCtmX
wNPz9cvCoLvfCiCVIz9rXpFQwjMVyTKudix8U5QeWeb5e5Vqs4tTRSbhIY+qmdZb
ghSt8ZgqbqdkCcg99GkG6X7SEjlE9tlORqx08lMju/5ihIeT5SoYsybTX05k4MYS
XnRd7J+bHdmX7vkDHT9yaHJmKDeEoiGaYYz3heajK4f+KqYDBhbIOtBfQuFBZafK
RIY58PGCishe2Pf3ed+SttL3GdFaV1cvGX1F0ZpCWN6B9GG0b6rtE6Ht+jnct5n3
D9ARP45OiFMrwXK2HcTvQmyvdbzPRgx0+TM6Jc8jmK9RS1wzALigO1hfCW7KbdbO
i9H7pCYS7623C8w7H1YtY+m733yTVU331yKBPS8RmNCkq74F/M7/PYIE36xTfkiQ
a2RRpjGAAFPAFFmVCxLGBU24JNeYlaeleKMThAJvZO9qk927vu0kfx1DCVuxK6RG
sbB7k5izBdw0kf5/A+DkYIhrA3/6UYWeu198hMtkKqYVdLs9+wIQyZuH45TTlGo2
imFsQ9Aq9RTJAALfroeQWbnVs4riEaKEyqanH4rDBZNlJMj8QW53vBh8P4b3hPQC
NZE7fTjvYX0E95Vq5niWn49E5qIufHlB6ZwI0tUYMdwYU0733ahkTu6Gxi1dhaKv
noArY3vp05hjC8RvomzMG56F4qbAnLptxDkuMsWkJbJG8rh3zZrzOute7rjpwpSZ
MCC9Edol68mv1TF1xNi6cfPXnccYB91kGHqb2RKDbeZVS1xIaSu3P8wAhLwYPfnP
ggBBDY0XEMbMxk/wurQT69P5bKyMk8rkTbP5+Bd8uS8yQtLpfsdRp+gtooxovusU
JWk6LKvhHKXn6YXkxwPdle47a1j9871iRXi9DvDGCi+qdl+pWhdKsHmjRUDY8Cnv
1+tXiBYACs1uJk7KiwjbKnswZSL2LnuxZUTzpIqbMR0LIzTybhlZJYKPAPPFYesx
4ZGq6ySlNPAbNYTVhh8SacovC41+g7+cqXo3l+bAtI4RvpEiOlewKok1qKgK0Rbr
UJn6IinAZM1aUPehDt+18Uh+5s5tBX24zUAL58MMGc9/h7lxPvMC9PYM6nTY9lK5
5ssh/IvJiljkos+Rc+zVe6IgCOrVKU5stuisx6rcAEKCjJFHU33Wt1Q6ljheviqK
kDOkG1NFVk1HWUQF2lE6dfisYv1lUG/K2D4sinevTEfU85B10KvFkFC82+6hiqx1
6cO0FGVPyOYqTLSNsv18PRTm6qm+BIKX0vADG4xQWM5rDvPVMHe1pkruobe0wjWa
i6d2nU/7erzkHroOISZlD5zKdDtPTVyR3TrFgIE947O1TFi/Xtjrxl0Ip45HUCT2
/B9X8EzqsIuca+PzaWFuFpu396S+nNj4XJfKwxKFzl+p0YLUbOhl55kFmwCzVg6j
EvtSmshogpc8ERbnMv/FufBZvP50BreizH6FVFLJNSLmoifF5EdyxdKQTYyuLrpO
zcgAHeQ+9BS0ElWZ8EEEt3+s8kKdu+CCznkabFNLlYmr7rg4wdcKJljE/qJmaPUy
UQLNi9cJ3e7cz0QbchdsnhVeV78vriA1gRUStD26nyOTuO/HxTfZdA4O+KjhnWg8
9MEFH+xx6X8jhv66sFo7L4GNRhWLLM3kubzCX6hEtu5LFjWLAHSZf7c2ITek7Jdz
W93nDrUkRdg8uWKNLuOHVpx/esFVNjN3zolW7KW213KBSvmM09eTxRpXIBr5EByy
4uWpXg6aYGbEnmbAs/wapJr2eSy5yWf/sYU2Ehnpw1+Y0LdtOkHVq/SAkQIMql0I
QsJReT3RBdJ+mVcdTm7XL0gaaADsT0wQTo7KUecTS19gOKWqshvPVJaoAGdsqnQj
dCH0kM6kI9tZe2geca6OjQVRwgjF1Z+X2CuINsrffDavox2GaUBxXxjJmTdxJ8PM
WmHKnYw2yBRA8Jbyo2ovvDRRrUSYniWcYcVsPMtoPfMNk6HRrjxDwkhuEovRRfzF
29/i34lzclZXK0jv9DxkKxDZ3oFdEX9asWlDhflQndTKeOw/t/gubC5dHR0LqlY+
gJ0GEcGUMSXlTdeJLIB76JuqtMgOj6QuzfIyStPptrhef6otf/tEME9WZz0jz6dq
yD92oUUv9zFhuTCYj2yukhgwW1bDknF/pyX3AlAnrPYaEmv5JgUI+5lGhXyfLoWX
Ilbs77ggB/NQpOJSv4T8OcXr8Tat1l3vTYR0TAfw4B2WQtegrg0Jah9DgABRVbQ1
ELKRGTw0FWYw+ucZOo8ywEgKFdMxPR3ZrMwBdDzv2ZbKqiEKqSTzfYw9b+9URqjs
c7ghBkDIQxsWkRObYFGrMOBHf/Hp+8cLLqaUxMBzgEFsRtSzf0ZRK6wDIF1aIsFa
EFM6/QibZP4xBSep8vc0sJ+aCwOgC1xD0S9//OjLZHqm3cZlxLpE60GqFjDRoF3j
gKv3O6yCBTLIVgeSlCokUBnJbB0U0GxFicsCNQkoc7Y34dosMC7ia9/Q0zC3q3Wa
voYo+nxg1v3ptOxWMpjhj4BARGwMda9IWBwBx3ktDaG2tion+bpl6ZN3WHhytEhb
b/DIMykCqCDKvYePVNTSNFuyJxMr55c/1+AnI/Jjii9312Z8S/HOtTNi5Q0Ea4LJ
7i1LpcjaQp85TtKQ5guf01HN+69dnLDFOCwdEsbe2WSqfWqkZ7qQfgb+ayZnj7Vy
YgsEIlyJEBEYY7Pjn5VsivXcmc4tMjsTtoOCqA6srN1FuR+5Rid69q4ESH9lQpU7
8DtDjrlaX90oM6GKl4hGp1+OTIriNpbHPPIeCGdy1hT4Omddttkkch6ANNIwNqL0
GkTWNut7dyA6m3GQw1QAsmLiLE0Rk5ibvhxVwgnZkF+4k1K3heoh/Bg0CWI6qy1w
MT8/t1O75SRxDoSGEPBuh6+B4UrzeqrRoGAJQu5H8YyiTDQoYjKM7XaLju7sYytn
5QMJdUDUBq1sSsDFPgSCQZFwRBhVAnwE4JIel9f97B/QeiruQDLidziQXpS1ULH0
KDgmKqyTphDQqz0qVpkqDYkSC3kdEXnh+JDP8x4mUPTahy5VDp97sToMSFdm0Y88
p7bwb/j/MQxO82L6exhH3A3qAw0FORzP3jHgZwuYfQg+K30SCd8JJVH1kZ7a7C2/
hndJeezzEF0KezNflBMi4ltvVFOn10BviNDhS4+nLP7uMkIYr/BPUlG5j/a54dEN
4vPkTeH2OeytahFA6UbJrRBOFT7eVPbdMIWgQiHx23AyN4v3u/I6odW6RofkpQD+
GfeoArnohwKA2vvHasMYYXa7ArH9fppNoyyuCJjtpA1dN5TIKs00HkI4YiLLt+Kb
vUEVIzCTgbu7XeBLc3edGnv1uuUH8VNeb8IZlg8ChA8YswBPvuBrXldmR5jRC2A7
TJKrV48X0weRPyFPxfKfzXBNgbzrvusth9pQkwUmshYzbGxGPL8Nwk/0avoL8HG4
uj0YRsUC4bpusz7SGKzTeJ1biMPWEIDue70dLPwEjA2Ckja1okOZghFWfvol7DZi
OcMM/tGG+ekdzMNbObezc4vnLYahc073BIVoFXrkLsopOEflpeu2T0gzcfgTtHsh
HgdFa2+ve4w+4hTeK3uF82U2HO0Un0VKhpFZy+YImI0uX5jI58dWlwZ6UZbVBoGB
h7LV5KnK0bfTmgUw/Pa0fStw0UFKDk9uMw51Hb6R2VxFyAf5dKapjQIoL0Ku9rJh
m2y4QdqJaocPS2FwsHOeLkZLVE+3fbPM4lOxWMDv14wGkBYLSeZnMbhvxpRvNND9
Rdr27cM1WaknSp5kywySj1VIcmviRK1zna6WzQ8s3tEtyz+aKh40hg25A63m1wGA
w//3pD2DgkS96X71LOMHFJRNcPuG1KGWpyPgEMLI5WiiXa9WUN7tHgdT2zTQsJ2e
LZS3Yr2wPNZ2ggTYPobBv2W+SQXy5Qnh1DpUcYlD+Qpa7rwxfEbcPrAEmosfRwEY
q1D2SyLmzbkCtVYso3EDNvHClNPldvFq1GRSD6JdMczfEaSkt6l9DYMRUfXQidne
1eKrKVAeCxq+nZDj2IdNJUaJhFY16Qvu/mchc34Qdg9hnPINu01f0in80zpdb5XG
PJHqAMneQEz69v8uiCI5dVX/R4k4bKtTjx7gGhtnufYtWmbhSRRuw4mgL+hG3X41
WhBPd7VK9M+u0rKuzc73GJBkzRK1x899YY2/aLN9up2YcGiWKRwNm6fHIY852Eig
xkF7frElrnfi+riFNikSjcuZhFTQZDQ0ORXKHPQ1sjEJ3+FDe39UijCL0ABPSVqe
fH1fbhA9FGpJ/N9ZSB6wsg/hd41V6zbldQVrF/ASAjaA51d1HIr/X8F/zOIl7kRF
2q+YErdiuPg6X1br82J8RnlKZDYMA47uemcE1x6XOV74I3HKE9olYF880Av5C7Sw
7VXIq/NbYcXc4i7C2imz7uLpBKTsGqL/wweTyPw620rQ6RA7eFHk51W8/HZYUtzP
X/vMizR7Z69q65kziHSiCEx2uy9JwcEjbN0xj1VQbA6PB8n6/HVWlS2+e6kDxztm
GN3YJmKcy2OGxT05P8llLTFSM8UKXL0YW2W6A7HAdx2NZWtNgDdVXrrA/UVn6Goi
isqmQVpuyi6/T1A9iefUkHd/EQixEHGIEmMQnWEuLDY+qs4mhd9B+T+OpNNsEv7C
BwdKxy9W91gzy67Zp1FLVnrR78lJzNRW5Hwm/AF1AXw0V2RLddQD9+F9FzTx9GmX
I3tAhu9IPfXEsa40gB7ci7DfjHszR4EVeOVCyR1RUUe0R5v0WAmXHQAHv5j4r1qz
34BZ7V4C4ivYMOYtSSFy8Qwd+1zSUnkdKxJm8sS/2JZ5XDOVpYMVn+pe5zixRIRE
QD1VRB+Q2iSNj74e4w9EhNoJuIyCBa2bYk7W7f66VaHZJiZfifMG9+Z3ALoBEboY
KQ+WdZFrJqB8Of31y8ErBLo9agIQudtBP3KP+WfPxrVHMr9sIOpCuHcuSlgCeWZk
2zfUmFDgUAw7h3nM6YcnBxJLVDhFTppuxN7x1NMAa/KsuWHfEKiNMD2PbMZSVQ/D
NqmZ41CbnqlzsU90pWU+pMRmBC0JtDJ0O6XPbfpYE9iRuP9f+bIIJpuAl55WzxWu
nAKd1mh8EFfTVLU3AqcfItwpAtIql/gyMz+6cWcYvscgHrvlBDOl6kkLvmQmRI2T
YgYO36bxQqGTBPCKd1wfqtZArDMETWeZxqd1TlOxVo1AJNmlcqzMZyJd2nfTJRPp
WkK6VJ/765v1jMGNG/kwU8fXzDl9mGI08TJKd4pG8GllwfFHba86rYySlyGglDLT
IKC6hbYrNZN5WC42Qs8Q/FfTpSrmE23Uodh0asCK+ueTTCbkjvgavbAF074fChkz
HdYRdIL3rI18DLoficEj87xRCJgdc4cB8avAWwcKVrfX0khvoc9aHJfebT1xJyoV
mj88rtRdXCcmjYg0O/4AZSWjIuXw4sHrpHgWfToUnY1ufwibPgp0OII0CzZGnYjW
bc4QKFCknikAH0gPMnNJvlNPjsK6VoO0V1fFChBebH4a45qytyp4t4ecT0hKiM2s
AciJw+syKKoHbUE5qCpU+VXXXX+q373OyUgTxOWJFfnp1dP8fJnmVIsapjq6epb1
M6pRViPf1mA5QgyBZBlvVJcKAucFAgufWIJ8MRBIP2BfVuvc3k54DFga2TVUvcEx
+hdFxAXogFkyGL58AzM5rWfNNAd/0ftEDwt9eONfbfoklGGJsXGGJnBC2ghJyZ29
PnhHJ2lXL4zqm6FjteJwfN6j4AdeithAFUlnrDvVDjWqGVJwFKFYEHl4dAbAFHw7
cr/QZ8yglauDYRuaEF6IB8uFX1alvHZvP8ALHuq3lTTxh3Weuu4ye00YKU/zc+y2
Z1IAybqy2imB97mI1gTOJh0XL34ZMa+tSfrxkN1eRQFlKUK3/zUeUmNLA72t9T/v
qNKeTq8HN5AGO6FgvtzWAoBgS9Comt0t0rH1+zvX6CWMvWGaOEDwLgsqZXEB8UKH
vum/Y1v8mo79M1kPoVrg3apBILO8WzoqDDobPhYmZ5JU3GjzHkXHCu7dHCD6ophA
ewUlbwM9CQ1DA2sNTQWpF8Y4JGuCK82sZjO5FeqsLwMoP4tzAqyptpxHO5ZGhFb4
Ww3e7Z4qPcJyedMBwULoRNWXdLf+np42mvsXQvXZMrxEHy+bhbaubbqQ9gO0XdsZ
mdNIXr3RpcHa6lErFCrrWuECBiO2XSKIuYuiGlUS5cCmLcLTOgm4p2wQ1U963F8+
j+K+t7hH0RY1cE9mVX1DQo2bPHwl18eX1e8qSA/zWRrBiF25VE87oJAKrtmpsApL
gmvZqekt44QvWd2XwuEzVYgp3m3vhwRgFQ6Hqhst1yZDhRK+e51D+Th+U/p7Hzma
AffHNqHxUV2TgLIIJCnBTF4QypwcShBqwouTvzFG7jnikOBSorzhEih1tjVP4y9v
e3TBpv/rhloUawRtWoT0P+vJPLMz9NgFtvECygCHBNyNBge7S/G1boYIcnjjkqeb
2g7+l3N/pECtAji8NYiW6ofzkTbkc9bG0PzPXSxv75HWdRFEObFo+EPJUSGDM13Q
zRfVQ2CILwThw+9ZbLnpHPZveBFPRvZPz3pznWSrv/tN2lwLpbvfMepgkr6AJlOR
BqZDSOTdOVTGmvmhR9lfMTFghNgrmjwxB4zDoZ/jJ7pUYPbLstGBgs7NY7v/Bmv+
ObcK+5nSqq119oBSzXX08rnjvcBx12LY2vqv9ymLDpY5RS/VDj2XytwLObzAJJy1
DYEzpxg6iGpgEfQBA4qqgq3PL5X4EQPP8Mp/dngn4vyF0RqnHNHFD3h+fNCixtWf
nHacUNs++njoapxq+ipgfL+rVi/MB1k1F6UGk0P3u75eH3LVP3oaR3zdU48iM1iy
ClSxi/kqpc37QdIBDDxOT8lJ93VXHiLLu/l0+xMlXZmbCdddgSSZSvkOBdOG0cFT
QmEflH5rQjXeL+pO1XZ9aJFYHV7gI9bmZwGP/Rn/1ykRUuGiwhO12y6ohQ699ZdO
pEhDrwH4pLbMnVS4L8+lg1HR/GMmGVj4XYtsFpYVAiZN2rJyI0JUlBp5Ec3sIWR3
1K9ezCZYhIlM2wcoU8upnZ3uvaIE53QnAydkQvUPGx5na9vz2TtvJCBM8/LfM9+l
i6DACOZnakilKX3SLKVBcALUzDrDGlQPAJbxW1zpgTxfqi5xfRys7y5Vp62cPxHn
VKyfkL5oRPg2xZnHZeMBXzQD3sVQfe2BWJ5mMmNpkv21yapFScdTltUoaRjDGXNW
OR0ZSoPTWBb84KljqphkfHfGcLoLdPM9YO8/rmH+vQY1rR4TPbMf1RdWlRfr2uY9
7Qpxi1iSOhWbOfER9+SPZZhKYcvWgMuIXuexUH3S4P5Dol8b6jCq5zlYLjit71nn
A/Za3t0QZmpb5wL9tnGVYXRNDVUlOeWlQqwVV72in3R3X4SSnCZ72XRFYlFiNzhy
cXU1czF9erJY3EBpplUpX9Vm7VhRMysVsoUxt2jP307my2ZSQIk0eBwAhbSmf/ZN
I+mNK4EKdfo4l/p9ykjpfndr8dQDIo0awrdyHQMDI7BwKgKJa0AKsoQfpxBI0b4U
Dw5vceO42U9OaxujWwBocOsR1YgSLnRr05/jA4tv2zvPRyFP84975sBnEqQ5tRB1
wfI75UavfuVYWPDmFwSbTojqZZ+dZ7RUX0HuiQ69kjBrhXVddgz8zYBchuGWKdQh
OFtAOfbzLbEM2NWrJ8CMpGfYkSxZMJSQVmZHmUidC8mijcGIMe0IprjRPpEoMm2m
RNjt6x+Hzi6l/ZbaCkYWmzL3HrN6OnMo1z2RlCvbEaquhzvS8g64al0O07mr01Iw
d61QQzp2iqJESjYJ78b5WlEeVrtv6zuiAqy9ANFdAYHjZi0HFB8eDaYluqxOHHWq
f2Y79RcIIvmIwOveJx8ennXJorRmhYGjUJtf1Gy/ib7f2MNgnAYPlS+Nu19Uh9R1
giLtENW08oNIE2B0O4jZRdGjvzZtVbgRy3DI0uDCCmpt4QSv1kewbK6J3tHTxzsB
8m4zVZedtOR7f36ys3prTBIdZtnbJAuHx/2yDd1jnO7fcO+mNJlXWmIUFkp0762i
Y64r7Kx5eBc4rNBd06iSpq3b8VKYj3/DlsOuT5WsTQtEndvalgUQ3J5NAXJ/R58q
0/a7A9UBei7NYmNed+ds9df3S1tg0Sn3FqJRd3v4PQn3+MHaSK6kdxybgCbFsG6I
j8xgvWlWkRtoTvdbkrf5bXCzL9ud6/McFKZI65I49vuSpLdZXggUtZ9qJQ0gy4Yh
1Hk86h8lKyTZj4poWHR0TX35GRqqh6j6JMQrCFirQAyB4Qa0tXrvFeng91uDP3mf
xrqX8sHWF/1rIbQBYWl4jzROP/tBjbamsA30GOIJakHEe9KkNrPNIOpvsm/zlI5M
7da/kHGHd+gkvh4itbMkHN73Sqb4WRn8ZsYQEbuOg9Fm/d8tSa9qlx2K15pqYDJ2
yi5BexR0y07g0Bb98UIYm+gRkEgJG2BNwbnq6lwWuaBgSp6nO2VOyO1piiUJogwa
jJJooI4MGh0WUOWUFRq82+eB59vp8FCC3xZFl91IyPRvS/BigeG5UgX020Sv7Vtx
49Yaso5A7wkSoq15QuOjgkcJRFUYU/TL7nxGsrYRlUwSuJ1QPXWVIrkTkM4mPH7y
tepK9nug8we+qrUEMwyCsChUFwmnfIF2cDuQ4rAbmIQvjvszUOxD7bSLZcAnubsi
/W950i87+vGrOe8c0ukdLWwlwRgOz8JzmL/mp4wTEkS5Df/TkFf84wFkVcak+ZtU
PKQEmY2sDwUCcgtMQOTMkyo6iQV7f8zAn7oSgB4YJM/z9vu4iM4DPqxgJ9Zk7u26
CUE7qi6Chq/wLuR7c0V/bpo0JFLkNly1AXIQWIgi+25ByGwmv389CfnOQqGpuuVr
8XC6NK3FAHOIxxEnIn1yzBqheIbSglzJknQ5bQZoYMKg8GJG+LhLHQpROzbiG7n5
Py2YXGvdBONgRT+7D4fWxgD7pNdi+NkLd30qUWDPVE0zFNXoz+3eMCAdnbDiDBbA
xWhhA53dP8Uml0saAKqHkH0AnKcPWP7EjWXGPoFYeMKht6R2TzeV4HnBV0V5wTco
2ItqHcZvHc/pvR3VxMzWCpA1mF3SekQ9dTiofsO29gdXxTH773Esn2GT0dvupTu/
V0hUGMbO8nQA/v4LK/vtfihooAELfIFavRfEi65jS9CsziqQ8esS2RFI24omUaLP
bQkktqoTIvNddKjnqx+RQytkVxc5VnY1XjRTocIhaJZbcMs4ICrYGfamtp0GUd8m
sRIDTrWvqXN+BWimvKbge+4v5ZouaAIZxjkEkVZNIEEoudRtRat0io/Q0dnQ7cR1
iukZKq3SlgtGaviwzQiQz4GxvhsAZv+jS32PRMjerMoPsglWWaDJbO8hgDbtsRHz
LXWyayOorbUNTytqh2Yoj9RqTsM+J2e6S2v6jnycuahqHA2VfpgUjL5UlgGml8XP
FihuwheXXTirmGrIs465Ba83Z1S1qa/aWvA3iJuO/+sgjy940asQQ9imCG3hkdBP
7n/hTkMYLBNv7nGWOl69yGR6u1b9xT/R0TlSjpc6pb63mAsR5oDwdVFrHKY2W5Qs
ugifJNv8aHa6z9IIyk208KUVrCIcngueC0AVsbeVEuU/t8wn16K4CHd8sOejXYKl
dq+sYMeHhwVXJr8mCAaa5m+aGBxmJcLc6ooBbexIiehhUzUDCb0OlRprL6X0Gsi4
Y37nhG76pVElf/66H0KvMZmTlE88sSq/6cODOE6lCRktT4nvhUVEXhdGlVBzsIQ+
71JdP+fb5BAwD/6YK/NBlmHLWtFo56q9Wk0IihCdFmPhR3Tr6jvLCdh2SiX26+Nc
BdX2OMYEEJ8egZM0lsXH7isvqSyxZYEsoFGsqvoQ8NU9L0jY8BC+BrEk5iNY9i/O
3ac9O9xXKTkyBtKcRaJ7XcarFhM9RX4kwND3qYjh2M6KZkwdj4E0wvca4PeRAmmP
feWAHCxSTqxg728JMR9L5ldm6sDyBMdBdNezmud4RpUmyJnvZJd1nnbP/3JIrskL
p8zn3EQnK5bzdlTnwGXb+tNokKS5ZDQjW7o0Zxq+PHXM/XauRiTVVRxxQ34p9NEC
5tRLncmw+eFCxW32Uf+ts99dSufCwlDXNDq5FoEijzTNg8cDX3FbvyAR47M7Qvg5
thSZ7Od17PefxvR9j6bFbVU0FHWHfJEErY29il6kV/81fj4A8u7f4vUEGfvGHO4r
ROyFqiLasEyV2PneDsB5xd9FYVNgieP8Ff/1Cpu2ZMr02GZIhMUfjquYIwziBCAu
QYjlGlRFlvyF4FRDtFCsFRCr0dksarxNwR9rYRkJ3BdMqqjjY6yxwbtva5RMS6w5
AwnV3qct6cMopOGSETIpG9ctF3ORJSfkNyH0h69tXLuhM7pOIPoCfv5etcFzz9io
uiPTnyHuLNwGr3gKwbJvAt3/409oCCkFLPlV95fAmLDmCSfg0cdgNvyg16xjRRQF
JwgV83cGPgGrGOXuoPIvtZiN4ea0lXcLTWOlz962d17Np4XexcFcWXK5nC1CkpU3
8KSVwvFgnn4b++8SDqFG7s8yJK97MZ1WPcq/7VZkLapHFJDLjOZE9bjOO2XdALCC
P7ygIN9aTwji/8TJA6zrXVSsGmWWKPZXpYz/JQHxft8WWODYF+HcRi3Uqb8pOH+d
aHxtVvLJ2wnYpteSlN8rpINy9Dv8KSWz7lTX/5KLRzbhFkgp3g18DQfpmObgVd/V
0RBpRo8SHNdKN/9m+f4x6M67SOEZMqj4spf36mn/+ROmExF/jbvPMYH+PVuktxfB
5dxicuVcV4bzQSiNKtepdA5wpAPFCXTSsbPJcKS4+1qOsPPvq8fIpWfl3oALRb+C
Vtvq63XrFP86XR52uBnH9EZ9nNYgnfAni+luHXqvRcOl01SCHa5HSTzdvTuuONXt
4YkKHlMVD5mx13Icm79XNM/UiV7NYCFl73hdj2HoIsrm+coQeuKAYBEYFrYLl5D6
Y0KFPus6Cjzgwoc+g4mFlwf9Jzv//KTNtfthe0bpE/lmv4//PG3Yjj//kZHt219K
u+XVr1GEuuU5vMrYZU12DZnz2W1EMbQ7YxXOlfzUPTEE6YftsJSVtrCqPalQV9tK
I9NBKFf8Xl56Lt87uEGP3Ql+g7DSSCTwik/rEpLB3q2ySv2aznXvgSGG08Qorc6Z
xQy4EWY1LRMyCT8dfrdV37IWoS8wKkIoRDX5KCIqx1JRAvhhEldg9APGC3fV5rci
wP16SPwA1kjsmKDtZxgJP36r1I689hRfYpOECsCHG7rQA0eTAQEnmiH4mU9NsRSs
cR9+jgYLkwp+N3eyBYVrh1rgaahYmKgj9wriBbGSWji70adMn3KE93neZ2HNTsfd
8vk/gK5QwJ+/qowmVAsu/kQ62jfcHN+XRdHp5bzrirwjSZN6RM0d8YosUzpxrjAv
U9wRyftIubRAnLHoCEbfi1r9lSrDQrnBHJSGjsLlWCp+7iRKVbcBVPAQxFte7TNa
GB7wqHe3IvLeM9j/RiYbP7HN/Es9RD3f6r9m+W2jYhpClDMaS7QW2gct071fFM/n
r3t1ENsSkhfBjXhcdQh0mzlEdHdIDOtUzRC60AEMnRy4IV13OAXXJx2qW9+iv933
GPXuWQTmMeD8lR1TbT/CJf8IFitBUDoGq/NHns4ZNcKGwb017McnBOP8NUQ53JbE
ijm1Z3koCRPGRcvLlLITB3v0e47pApHmZT8Mq0UPq1OuflXmJCa9RMhqN13HkH7J
GY/OzK/+W/strAQ6h7kvfDGYbBdXDc00GOpm75aBdirc4dwAN6a8kXiSPyJ1Wt2Q
QoGxoQjPHjeVR2X7yTye+1hd8RECaddYgljfSXArP174TnqfXUDmgAMMEd8KwKdc
3PGz9NfoVQ84nEhbj1W3l1FzUqiMSgsmeM9mpPZZ8ASNhdOC16FuGTXHi0PiQctR
rek2mja5f7UX6s5qsZeyups1UjxdpP0WcfYrFi4NEzRjX7+2i3yLprnIT8uJDrez
6v8zATDmnBO/VHmhL7GkcTtP9ce1MXEvWUBbce4l1ilEFRjKc9uhMjjgUwr/KOPj
l+huc/oMyNZQCyMQ6DKdpSCvsXFTGRyGQpDxBjEJztFWmKB6LcBQbF0xhb0ARq6I
rf6O8NPzuEAWtJnDpiUgaoV9aV7WCd0HmWoaeeClycaVfgAE9cOG/CGVpcxFBBv8
dJiGZIJuegapK8NRxaAWVxu3HkJ75n/5UxFj8JvnfyMOSL0Mbsm/uZSXReTEyzHE
wD5UoZP7RjFRhPWF8CHjysMtrn+Uhudg/ok8pDc7VSRpZZNwDSR3PBxJvbd0tDuu
leYearp8rGryUbFh2P/z11+4HA08E+pQG5tZDo6y3oD6VEwa1XX3hJw1tmdCwLQe
9JzIls8U3qp4vS9MIqM5hAUsj+mifZuhVHOFWbraAJHnS2i+P9yCRD3R8IjFBEvu
8dA8p4TDQl670RxqUqt8dTYbSk/S9Rjll14tvKtorwKXbAp7RdQFk6J5xaJZZsea
2KCDc1wjK3oTY9LHK3H69eOnim4qVOetM6S9cX3ZLtOM06mcGt3bu6NlCF9er4IK
MnFunu0JntPNBxrm1pLFB7ALJw/y+OSncYwuwUe/k9/gHVm46oWDADNCwG1QF1EC
R1S27Ki572eUSU/uJaykTO3fRkAqOuP2PjiFOneHl7hAvCWj7cgL44FEMChaK1m1
tN89HikJmL7SyY4rCdWs7XDXlmdoVaQ/Buoyb02DSgGkvD8U7aT5DDBsLOB+PSZe
OwXc/+r5GJCdnAzoUM3nwcXNs6FlnejHROxqJLgjfgHwtEZj3l96h3QXsv5ySPES
OirLIFBocma38wZu66xC4E+pO3d7PpSZrlYLQzRVbI3+pUsSRpmJuUtWOAGcRw3t
qT7qYfATPT9FlUfgjGTNWIANWdnDfL49r8hOdKNJeu6kVp6d400JvCwRG6ZphDTQ
60d5OIUzxIxnYWkWcqLnME8XuNcWm90UuOm4jNHebV3U7qI/xGS4w2PMD5rU5liG
tSfcOH/+KRM1RZn9zM9+DzYuiRwZWuLHaUvjue2lc2uO6BrSol7u4Cmbld4LGVKB
AF3xGyFk/vA/QuICbQCpMQ3x6lD2uT8k3/Cc6+pVknDgYp0VH8UTrZqQuSU2moQc
+GRB73Z/6bqggV3nhHXBLtUccE1zK7truTRhEbDUrIMlMEyLUbXi6sdF7T10FZWO
2ozt0y1YcN6vtH1TLsDqusdf0DdMSR50LaSdMDNzOsasF0FFmvdVhEJTCWLwY8kY
TgrmhCz8WtxN5KW9Lu9eWDlnTad8+BHBUl7W1nSBCClWuFC4UBp6hxzd0lneYLAK
YZUmo84T7/8SNkb2bqSrL1uUMwq6WPwWsMoS3x4GRzhaTXMjkmq6r36bhohQqfVo
h6/9KxbpYsPrVS9hNc6aepjkqaFMi0/74uxOsqvlDPiQwUYvFvv+JDEC8UhJ66Lx
dYc6Mz5zHHUgnUd54xsAWKLC3y7HOhluh5aAL7dyWFuauW51jClQIUIDT/MBSg92
pYlCgRCqrKP3Kpx/gM8EV7gwC6lyEjMUgT7jtBhauHCMcSKRcujXuxiQYFAJ9zwv
G+mLGIAG+PcZA+LnqxQZsXISq6PplyNX6o7Bx7Qp9IhPk+DaFtYZjlT8QJLSaswx
QLyZWcPN4ncNEJ7TN3OOiTG0fE11ICwTsLxaw0JdejgVLoO45pK5inrOfZropQML
mG8fmjuRjI/uoHfDowCe7mVTBvj5HtvlbXM3RSAzwi1zr74x5ILpuz/Snp9GcOTy
TPgZdRo9A/nKpT9/meZcnII2EUkiydNaN8ck6l2Ey6FQ1DnC32+zVfMwrEW8QPeY
u0BK+2X6xjNJR8c124Bn5BblajSXOF+7mbVP+oXiaX6CbKNoNh6uI//zuF3lbAyU
MDnK3kIJA0g5QoB4sFtYjUfWCzZDjKh2jq9HCi55XdakqsHMQNWiskdas57RpMII
3MrRqpZSfuEFMhzFIt1UAA2W7N8vu2WWyvRYGFt12QEfO1PnYgPsMSeW1ef+K3P+
zcqkFCVUfxlIQdJkq3ci1fnCAu1GrfQvhENRpe8W1d7VDz420En0wYZ0gDyRx/pG
KbH5iXxo1pexfzl2Yf8Mg3hDqRF8omV7D0bwovOwrOEWPUYsepXw/FnA/Hi6GN3K
4FXAKX1wgtPSjVBLeEYQUBrz0MmbySac/A7IUrMSYua5+p22/7YaA76NeWHCFd1T
rXXu0RQz9rNYsX7eb3H74FdWTmtfhIs1QdiuhgL66FwcsS1N29S3siOqj0f/TRKZ
mOMP2IM0cMX78La5SQbQ2tsyFyGbMFOAK/dW2OCFh0/iCvn44V2Y0TtZH20fdGrB
xsmhknmjwlZv3MKqncY4EQ5oxBWr+mkOGHQBN2Zmub2wVyoa+tfyOrRfFFDimLOK
MK7zeiZSZcPxLvYRSjpcxDG1iYmmV2L9beerAUKmyIgpzz3Dbmd/QMfvgwlbnyzt
3fSEsKhISe1qWiP9Tc9BuVMAW7fHtaPs353yT3oexU+RMPta9Ij0UOUrbelW6Qc2
IdcPADusOANAaVx/6wxUAXdOlW3mjk1NqUaDrqgTqVNS/wjoKNlNZlvrksF+vsqT
ZTS+ohqn7Ebq9gqxZgY1kM9gB0z9L1Uixm3swnkB1jEajENewivg6jBsvctUmZHA
Yz4F4pfEAwZpWRHxk8t2SsytchGCvNuqQBLIV03zeUDy39RQAyCyBYju960Gb1BV
tx64GQFkKMJj60WtT1t577cNMsTmQccJsD2JjrpVFgF81Fz+HbWnmODFHoLCtf+7
tpqSOzYp3RVT4czOlR8xBPCSiklh7XbJq1DChRyL7FmZyqeFUzZO18RKNYC+Rof4
Lp0N2KzLSe2oTGhuPF3KBT6pOoIPi2osHqa+dty4cINOb6reqUkFN4SCqWt/XNVp
YhxUJ7H6tkZxQ2pkC86YM/2oMQpM93IL1RIjQt6OQ2k/kzOc26Iqz834hACPVWWz
PbUVNLb+9jTur3xNoU/sRKhXBdhJwBu53jxiS9SSBIsdr8lCZnZwBHnH5+0PA0lf
mcG8kZfZaHKT1HZth8NRQIaG5V69EJ++qtI3D+yPqUtW5xNMAw0HWXOuU5+10NVr
IX+BdTRFhFy48VLbwfP+B32bzEP4LvcHX7jzxN3tR3lBO+2zF8Hz9SDj+x+/gtmO
tuAxS0ydMEOZA75R9EXCRLH6eeFT94x1uI5riTeCXg3IgHarZgb0OOuxmYzXS6Gf
/tYuwejETkpquBhC44MrLnHMpwJZ4hkL4RNL4PRvkK7NNfwgsJXEDW60u5iQJeGA
VV9K4++EW+6QB59rEQvUPE0LW6NFSGsLmYh/gClD532k/n7F4mqVbx/74qG7zWi3
B8WsZTCFN2izH7dgGpUlGcYK1w5whnzFCO1vzv6KZHygfMSEBrqQZklDdQNQmmQK
MHInIAcBdQvNfvPklSoX+uNHai9ChciPF2B8FiBViHvPEzm6Kv8tufVlqlwUpMHn
G5uymwFQ5KdsWN57opySoa9oiwiWtOiNtuYNjihhaUAAmp9xP4zif5wmKH0GNGCA
hE6kle6zb62YvPEpwGEOtjbSkZoOA7WeUqoT8DHJ1+zCRN09Rpr5Azz5IDQZC4Zd
r+V9mcBjNB40CHWkwozjBPcSSyzMFGC4Rwq0Fi66pdbA3m0CfTxBagi9auxM/iDs
xrBb9eoDfHs8oD4w2tXuWpwppVlsaeuyTmbRigYbCh3ke5nKvcaiFWmJAdRWJ29B
AVQGZvIxjzkt04vI3S+UgbCtZhOyc9IjQ3G/biYhlhE+ZDxGAHjisyuXpfWO4pzb
5hl8KIqCdaLN66rVURa0G78J8w+uWEZHOOAzrDHWWrGyDbcbr5+P31aJ2GPcG1SU
bjx1IH3cnC7Y5pedk0ei+NTWFc9/67njIpbfX18UL0lQmelOPEedO1DaChTmZiyK
IL+OxwfWq7Nuq0tP7/czGCAGP6v4LsWQ9/Z0Q0j+ld3TzJJHDTQQ1YYApCurNV3C
3csTrjz/SrnF6pueruwqMwLPq9iK9YLj1hnU6FDo21qOpSuLDDreVmw2S7nZ8Ejt
LRF56KBoxOc6zTkPcyucY4igakKkFjFsCHpTyO0Z4xgxQRJmNP9J8mRdq/SKHFMK
4qsstPHvdGwYsnGnOxMIZO9TicB0f0sPlO02mEeMtRjoPxvy4HKKen2E4L6BdZo/
f7L665E28Thp2CYNsNA8QonfC6+6NIH1ZcLfXpvDhiptR1FuiY+7GqIexGBuGK60
lf2RypF6KVPJaLpf3navjnPo+dCmABMacgKfAxReeKj5+BuuwoxTfl6W6oSjalOx
R3s8x+TnPa2c6JgulIq1zD4qc4LN9E0YpOtgjcOH0rQ/Kcyt/MNGYtbnL+Q37eBV
I82JkRbXLcrCvJkTsO5sGtPBKYRlujxVLZis0I6oNdsyA8S9wo4Kf/KCzLbIUSxP
NbQGZJUW2MediTijDzV69uEV7Nw9ArC1U/AvYlGPqponM6QCJsZ73nU2VTWEP/oU
lzpEOeC6MXper8q3iPrKuoaAor7lM1jZ3FO0MzXHfeEmLu4GwKrPcHsfcedP2TyR
VWNM6pX9D18wA08+Ub8wpoAOwUd4sOXgf5t2cLCAh9jvZUHClSGKwf+ipkQCS1oc
aazfaaulZX04cjlwkeF2l1Wm4TlPcgmtItUoo8YJKYJcpIy4hjL/QMfQjvreJG2F
PP35tGTnbQoNjSgVn5fpZTc1/zbIHjzk5QA6KdDwRpTY6Q8cJaJMBgqb2pS3dhFO
AYDSSeWT/pspH2bxR70MGOPNTF+MWP6w0QX5PHL5500K6smDGK5lzFAjTT+L5CMr
xKJpzizKeNPwvwlKRjX/COTqqCoqzfrI7urVomTgFc7HhEyDI4geK31n1uJufhni
/fBIV6OrkOjHw2/40ILn82cHlbgrVAwbh4rnFId5UTbBnIPTn+io8mExZuZI40+i
zM7PL2UuiDQ9oYhDbSMWD6kIwKA1PF7HYxxYgYPXJIzxpEpNeswqEemi4zIVuecY
QaCjuyQ8/SQSElYj5IM+1cWuN3DJyTIWw5ZOtYtfy7vVMXEiuG2wHO4puwOkY6be
EmkfiUmUH/5ujpDQtvEZTUhwTkAczNUgVUzasKyUTVY3Q2J8QMvxYXEtylIyj/oy
UI8h5LNQ5ZsZ781jFssccsu2IKeQ1tXbpqobaL/vguo/prpS4L5Ux6RZ/S2meQrw
feWS76i3baNAcrkIYohplu7bJD0mdzLIVDkCuK9ysCZUzYfc9zCOqfmD+Ga76VkO
2j3ehkwUDYiNYnqDm6z1Y0BWH5dTVqT5iTkvTpUMX/npOgYKqa60ivAOuSCMbvBq
umREsTtV1afB7PhEIjDbvJD22n8KY1zEygH09+nwGoG6g0ZMEYpUaRMRuSpC/BDE
fMqYh0crxCGaXyL+cLQ7gGDocwObEivQJ6CDeEbWhMOYBgm7t72Lc44vtMs0Pqgq
hD+1qtGWtRfHOwjTml9PauWFpknXZYGqppj+OAdyVMWDTjojoiWvX/1X8A3ZXTZE
DttgWO7YYpSR+XeY5jY/k/F+atddn/A/Tkm4z+ZNhxoZoPz6s5ifmhR/rztPv4Ev
PbD8GVjE2I0702+PnRfKZyWNgBb2z8eImHeCAdQLmsrqSURztSGTRZpqSQQSP+NL
5MkvAXWURzHMQY3pwAPnpaOsE/0y20NwKC7X4qdYQy+GPyeBjOoFUo+x5t4NyG5N
ZkhAwW9boxhgukY1vN9aZZyP66Wed9TyW8glGkn8J/9vi68ag29CRBQW9XO80pXo
FIqvDMhZOwKD9KWKYMediTnpbsEwqivHm0iu+ex3g3ss6x7jDL7kpnLC20/U0Ozw
0pvyLBE60GGVPawBDGZlG75u/0tz16RkqWPP8tivI7xU3NEO8zdRxfXQ8g8vyA0Y
LE4aHbho0aoaMI7l40STeeZoUJrXH2mEllkt/2GTYqtTAbh5o60dg/NPqjryj60s
pX2X/+SWI3Xi+7s04uN8CzEPR0lNHe8K714HIX1nI30DCa6eyE4F5G8oSp7Q7yA9
UjCoB9zThQKMsqE1LD7PGb5FrpMxft1Ep089gHeS4XAkCjULXq//rNEnL4vpdOd3
7f0HhNmo9wt2Jutgla7VGiGLXKmYN0YRLsuze5Gf7oo2LsdOGa3pPJ/XfXbYhWUo
row6iZfCZhQzKY8ZEUrygfx7FVetGx02jE50UHfUk85eSMBW/k690vlLFZyfAO9Q
FQSa+b/xorssEzdqgvjqEWhfBLg2fkoq6wBz6ajRL/Lwn/grXAS/jHAFYwUa1fh1
wfoiJwyNCNerzZY0h4iqc4gGCqtBoaoh+vIg68zwXzljvLAPXpjVbJWiI+7HUC1w
I9Kyh630FS62I6Wv+VCP9yEwX2r400JXo6P8OEm2T4y572D5cXGAqZhSNJtbjeBZ
qD2CL66FhSpVTR2gg8AYh6D+4MBgIqMmAy1PSOImma3wWSTpvsrP+0L3sgaZemm/
oeAcILQepHgv55rSv/MQ6PyowsIMdg9WJl9gU8Fh4hTXhInNu7a/XjtjacS8nNjI
g3o31GVpfY0Xj4wrIkYCNn/7h+tSibxv7jUZ+yjdkjCUPHrAW5uAj+5VsOOzmGfi
jQBSazh0yoPY2pWVY/re1n3hT+cGcMAIlu2tdCE/+/u3n8VusuZVuPvAb2HMIIxE
YSN3JHRAh84eXHG135HIHwvCTe/oZ8+XzoLywk0CvfSwhAQuB1PD2a0H1MFq9NuH
2bm5MDKrpH8Bt1+iqBw18SHXqjcPIQT+H9RIGF2HWayOEzRuETs5J1zQ48NG2IYu
WJ3xdNiypuN+jxTJWJi/ibCxXPsSVIOQz4k580mEXt+5FB3GlZUIbGI/zPu8Ux4U
zMIcWqsfXVvktGSAlMuFzX2u3lXA3twp++hDc9SLeuKLW8I5cDCKWEQTHB0m0PFc
23YOSPeIpP94tn68ub3YqbzV6dUtzQMqSUeCNh2235Py1VF/dNX2ObCGXJXCb4im
GMab/Oa9gsbZ0Kx8yZdR6nM8/2Zs4K3Q0+RXT6wbDFvYUUJ1tEeq7k7oJ9Wt6+xS
jBz8gmOPS0P/k4ntCuJbqLNRUkkjwrruHlyB90olJUOeoGKY4keQEBT/m6fgdyH4
RhHKxHcH6dbROIFdPDMsPcRDFAmagWinDeoRvsdMoslv9FSoiGt7RWk5eLZkKrWG
6cvSnBbx0+h+zX5Awn1b2dg395v0RWRPH5iUwC4m7cuPJDXIAk9J2OOguRYiRlW2
onueGSEk4xNryaj4ip2dmQWTV0XtWkR5A97hMcb4nB93C5qVA40QwbMhh5z58eji
r9ogPaOLMI+BAx5XHDV0wSdhB8Xlz6snwsltGwKAZ1XPiPHiJUvGrrCJDMOWKssl
u7vCet+oE04czPdBFlmu3xdNUNg+zQ2/brBwN24+sXYWzSNvNLjEtV/AAxskpOs9
fTQMPlXlECIEmY3VJzu79uVSqjPva7gUMXQjaA0fpe2ieICnt9MAx0ehC4jyak9a
pQTT1kOZ2ZMvpPN0cn0QIDqe8zUqWaNo8SrGMP2FR/HibnJCHerruWsZj1HKDXYq
CeD13jNYoh71T6Is3Vd1D4r3sRpaiZ8J2vLVLarKYnP/xzkK+yBUevGZWDyt6cab
j8CL+BgSZfVtS1paNuWQTFGhx+9+iI/P1DCy2YIGWNL5uW3Wee6J+2cFQhPROZzb
58ewsVEvLHk4HkCGeb/LVtclQUQVI3NgX46S0vmwl4bsjSQLLyFvhr5U558whod8
4BYAYDfqqHRtdaQ9YQtur7EAoJeJHzXGnxc4wI3hFH4ybAenAyjPsw/EO1JHHFwK
g5cZ8JRxwvaAZkqlXX6U/un2y7TLZNutl0ZN0DFKFN5C2awN+JCusgXtue30F0I7
cPu9YHXZJWS/2vxi9il5Nh2kzaqnlwmhwpXfp+zP9BKhpu+XDftUcvwO2eCQK6qv
xResY0T8DcnFuyj10ngndisBStIcdg1SBSQc/kvWMXLc5IcLf8g6KZdvoWuD7CUY
NU/IanKjo0pBV8cDzCcioYbjD1hynGjDcdmad7RWGJdSaD6ngbvZ6ru6mKRKxUXX
b0ymrVxkWlqNZNgOm7xIT6SIx1GZKD3kEvkKig6GwbkgBUUIuEh3h/QPbuztOZJE
efp8izQdzuCCkxgpYBDdYittVW6TeE+s66G1NlFMMyV/SJR/FRpTlppjl+4sM/HL
UPx+XS1D5gVvPlaIRttub7nlT4+QZX/tcMJN+PcWogN4uioAUd2xVj13hEtN10CR
ihopAJ3MUfNoIxk7U/DaohltTwK0jt3e9ISYva4dgUFkoOUfrn19qWQQPUMo3F85
Ydgzmb2bbXPYttTjAdxp5zUu42Yb6grqzUvyF8Z7gsPUYn6U5EBrnpm0SuG1LLZJ
S0+tyVhzXXOGfbxkItIA3J7agTTez7XJE6Tuye3qWbwhlTTDyPHm4UaffA1FUwIR
BW4qHnPTVr01E0OoMvH1bVT3G/LP9nkFpl4hMbX22XUFTTceuc/xQ65oyJdbc+fY
JQL4X3zyLyxzdBLBgVva31YC+CPbyHeLJVG+5KQ+2rycxqvQuk9SxUd2Aj/Ad57L
f/ACM5tUrNdIgsaGgzBPtSaMl9JDF+ymnS2F7xUjeetLRyrswWoHxhomXEE/hHpz
6ljI0BX9jy8Mu0+0oj6f+5ypuQoLENENaW/uqtkwgyAalxhBphqbMevlWs/HST/F
+TDijwTimcF7US9hRGxxKh8MmYgMkuby1yF2NxGXyOKIOaIdXLc7WN8LtasSYwwM
/EPvJVV89136R6LWdj0fozevc7kUlDr8iGJBX99InwWDC4DBBUThVPdPfxZYbLzs
5UQ6Yht00HckHURrKyMQbeIabukI12RwsFjgl7TULRE9vEysGpMJaQj9Z0/N3qgr
lrkyeMGNJtRcPRHuRF5hqSgsYMZqGg/c+Loa2iyUbywprWti1lovnPAmiBCh+vXW
830gzGtgtD1zQh0TPoAoWAwQ5aktVJHujBgFlif5XF1yc/lXY7MXKcmFCfsw9lbe
5m93J9o/1OKku/1SDBN7ebItWbt1nrVnU+35iUP1EsjJhjWoAiDn5kxaeOK2YAvs
ngdMj2ntzAYyvsMm+28P5JSk3O0RcmyfruYZ+dUHNh9ugkx5P6WWqK5LfFPpiork
+WxgMBOJJdyffd0hpxwDCk0xpTU+UyxRBAa/s2fK7/VWqK470wfbAeUY1F6ptNRv
pJAasQ3ClmjI6mK0q23No1Ij1dRswvim45kHrRK0aWCBef7UtMqBqxq5Ex7tGw0Z
eQAyl1IIVcmdZFb/ksarS5A6C01zLXn1gQHu471uMQTfpiMpu0Q65ibahKA2DPyP
J+ry2OH0OYmYokCJiEvzIEDND4rNLZbljxl6BkbI8LHR48kafb0LvwpbyI/Xi12f
UyPn9F/rLEwrSqvXSHgSSl3hOcEDPyNQfu7ar54aSfEN/NFd4jw5onbBT28Ekf58
DwMJfeKKNukUsVx8t+o2jbSPPqOf4kyRV4bzPrPsxT1ak+W869DFwi/kVxrTLV5o
ZkUxkzlud37OS/XWpDnp7IR7WnQCcJ6Vw+WhnTn0rmwTDRM+cuc1tx9kvQflH7vr
QFln/ImQPbAgwO8gZZcbqRJtLCAaXxr++OxFjQb5ZdDiRLQ/floXC7fQZF8wPSzt
Qsl+v1A1onBSE1+haeR50uGN7SyMUryzRkxxJXF3LyLxPIl2CZo1tZhTgQRRD7hh
lroQmph8stvOQb1eb+vuV4bUy4OifOF/sKdn7rXc9brfLtK5nOblUtaSIlWuh/zE
xKqbQRgVCA36UoKgAYgK8evAVQT5rzx/P7+TDtx6jkZAsjdpYWOaJrW7S+V1RhCu
i5kDSsg7tIWrenOWFbFEjiaChgcWH80GIeHRMl+TamuPh/j3cGQeI190F86FH99N
SzC/OG17y1xUkdley7pNr1lxPBUmX5jiVWu+fmb61nND2MqZFJgnj8IAkCogSBYY
nZxnCzUQ8CdGhd8Zae58HisjHeaGvX1LMvRh/65ppRXLHuZWq1u0yI/eK8MWqfDV
1NFjdWocjw+Fe1OGO1vwtq20Z+d1aO6QUkfDKHNPg/IrZciy8tbAk9gLlJuJa3Js
zLTryXVQO4gyzZErozQabenyk85hicCZj3GShRdS9tyjcvgFzR3Uj0sFzsme0ZA/
D2RrsocXVE4acJ3KGGMHjNfxxqkmmIJDbp27jck3bPpGUFKXM/cfxxcHvtdfw417
XMZIPyzvj4LVhKtU+s5oe8lr/ty7agc6GCWKsR54HGvtWdKhbC/WLnEKKJLEME50
YecYV/e+8F6Ed0R3M+vsRz1UESlnP2eTtJGAlGlC9+SEpRj39h+Zi/1Rx/fP4Eiz
/+L5BPYFM2ZDGnOxNazgiqfaXKEo5gBQlmzFlBIIAgTr+XItU+xhfUr8zAygM//+
imR1Sd2l7eOuS94pnhjdYBXMmzcA+g1XuHxzFKZFS3Iz+hfRuw5iJpfSiMuMYBno
UZLHIvatXviUFhUmYBjyGbqX2aZuQay4XPvuUFlAo/VEtL7mllel8OA19jxCUu7q
gysuxdePaKiRYyllheIwrPiltaW2wBAVdhaLCxdcFmKQ0kpOZdVYQvtH7wGaDueE
S0SyYkRAlMsd13jE2rmT+B0iJ2sQcflSBkmcxFO4Vs/V9oRVpWleXbvyDTZEUgwb
G0Q+WqXmPHgqN/OGQenKTHvjVYJ+k1mJDlCv9N7J+Tw1HtbI95clwQeS1rjIRbq+
/24fkV+gTYjP7ZrY5JuU17WeMZPRdP1LM/yqZ8/F+JZyxEbDhjE+fVkgtPe5py+i
BJAV2pVit/RUUW9StHdzKU/zHZ4TSApfY+KioJjRmdEnufidd3GUwaWLYnDFZ+Gn
C9B8Ia/TH704uxqS8MkneCpflvPl7PuCq28yU2LYp9n75aMMSF1gQm54bjIXDNX9
Et+ncK93mnMWx5kIr+elVbkR13VB6FpGCU8WyCOVY9NQoHU0Z5saXX43BVDQmJ3r
Lv333HuRsSE/d1H5hm4wyhTL86V3K8b4NQ5ZHahrUPKwfXF6gD2CX5zutZ4RN9dx
RNvOkV0jhraoqScUcJvK185j8h2rDLzgZjRdyVJsoJeuyeGGQnhqpDSJDjGMiNzR
uXlLxwiJDAIq3dGHC8yNAAJkyhn9bPoZYs4U/JMPh9ieEOFghuJmLZ3QJQIS2cmv
113qqtHOnhbddTabUdJSIAdV/8MtLVx9U6ry79oG95wNyYInZ8Fz8DivmNbYdKMg
SaGyecIk8wipqYNnTDJEdSdyBfNq17Lhw4Y9lHjWuZ1ASIAW8JXT5/iwRcwGr6Y9
oqTQTSz8AWeJQYShfVFMu2DgjmeW0ERczG2z5CvrbSjgvjXUuD/n4N/UObhHnrVQ
3akcKXsHa0KpkCiZ+uMHmQyRA0IcJKx6A9AG8IqPULDWzPZ7G2FpAqk6bC1yz3lG
8J4aHOM+w+prys1gi0r8a0Nf1a5BNxzPNHLSRg3MMqDYu50L1vij9w6l4cKdVPGM
s35dVUeiS5k5yfW8GVziI1zwITzU9YbIh74wuSGvsu69boFQ+Pt7lpKIRW79K8x0
EBfJaarTRS5TQr8bkNQ+zJPikCls3QFUkPdPh5JC0BYrkSRR6cO0fALtxSWD7ma0
kXhBVlk7xlG8WWWMCvfJv4n6cQ4vxPAGDwUc5Yq4eG+kZE+7f00ZdViEufcGmPF1
3we5W8p/N8u60eYJTH7eI2f2/UKql8k4H4SvgvGwebqTyJTjsnnLBgFHXRtTXoO3
HZ50bZk8Rx9yeq+rrfMVAj+/zDU1tmrlPkLf58VA6LEw0HDg5NU197VEgXC2jyBA
vN/PHN9y2AAeqcG6FOfAJE/HWJgxQ3JLs9XfHMqhvJg/u0i0Zx3HTfwCuTJNqMiV
tt66tW3gr9dFcTdx1L4I6M6XFUXO0zU0sDxLQf8Kj36+fNmAaymoCh2SWzE5fs5V
Uz6wPNi29IkY0HpRvcEFY8IlJYJFT0ahwKXT0i9I175xtneSz6QjgvwtZj7TIaF0
DG/6ZbgQqtVtL8HvT5lv5dpR91PTszdZz79xPDYBAJ1RNAZONHSZdBc9b8cryb1w
HTRMfjcMxuHfBtVjZ1bjwhNULmgUd6SGlng1V9NNcUieuahEDlnPL19PuxVDcEib
Xv5Qm5nm0HnFZ2RjRCuwXNyFTgmqCeE5Vqvpc06Zc+8UiKeMCULsVkdXpD9YgkIH
SDNMop7B5Ew+2bt5Mwsw5PiTyd5ua6jMhX/qB7v26p+frdqI7zfHyx9UhQ8qmSg6
D5qC/vwbkh2ki0yC5Sv0akEenbyGRzTk8p7Z7Nq23leIdqkmab4hmRhiSXEXjjt0
r2WX8KQrBbE9QrdOlY9n4s/vio8L52PyKsti4t7dW490pU2n+GBNBidNj7lEF4W/
q4m12+GexBn9sAitJaH2Yvpsf4DJ44UY4zTZ+WRS75XHqJF9agZvFVbGJ7Sx/4I/
9JsuoHl5IbZMEKAEpn5frrVi4aIJ2sP/Ls/cu9LTD4mK5e7PFY1RNXHIU1Ga57XF
9/rsJyh8L7uY1EKlf5TOywGc/eJuTJ2syHxiuU3de5aaRftC5g20/0F9dzgvp1jw
tfgZuWW9JDSfAWcCuuwX84sbrwODvbvdXeYdSbw7hAympanEVyETmyc5VwxEn1c4
ioQ/mLThV4KwB6d3aTVAKwnIC4Uk3PKuRRj0SLuYItQNgxWc/80EjCN2PmSRIBKF
TzeQkBrqhNrAuLLU2AYWcKBIzLmriMlMXMz3qHl7MAHWV3xpxjOo95EEFAOTt75I
GHTxvZsb8pLI5FPBiUMI9sEtzjN+KHp3lcsXHCOuOZYEn7s9hF/Sr3vHL8qf1DfT
lTYE/SiWrdzaZ7pWWjnfjCvJSY1ueWlkBai/5vkgnnk5ClfyL1NkyhsyOVPbVxev
ZJHWMS7tFvSZ8eSXO/YDgCqHkNsT1EjcmAdiqxM3KFM9icb6UgaDj+gAbRDRXn8g
YjtLNfmOFM1C/WigpAtGBQLp10UsJLw2Qp6+woE2qnzzrLY1B96itSsyLhgx+r6l
Fljnc9usE80F3FMJErkaPSq/Subt2QX4eY0DS5pMLoUQZrT4w978XAVKBYgmt+s8
gdNmcCKXubExLmKPO9Xdc90G1dl8QgR+WLYutLX1cUBzTKrJqJ7cHdzqxQKU34pX
MZD/WRxJLmUyJAXHtHDXj2dsJVcX/+yAsrQxWzcjT58MZjdElLgi0zCnwV9Q09QZ
GL4fP7rRzyOn+QvCy/QovTqfMIPt1FCkiLASsI4/du9mBMPFqGD2z0OPu6dMJ/Nj
BhM1g0a+/PsBEnnV4i87nBbvj7tA7VV62hL491MVZvo89QrP5vuP4ZPqWPHIK3tw
9TRAFftXMa/ZzizlbGC4D1WfQLkjtvV5V7Q1fIC6hh1wVfW1c/diacweYfLQ+QR1
15GuQF0yX/qgs1ghZm66Uk1WNwxxrBmoBFKMQi2XBIOHE24ZpLeZYvkfzbFRo9QF
c3hREi742kJKQIs3lXzTRqyiHk9ErPspsfmi4sMbIvEbJhL4SPuS6IaIffo3ChnY
cbfdlvwrOvJIj/L1gCkVeh3BQkmjvNlG0AKtAcBdrWnuXtNZvVUwpSfb/X98UlrU
nGx9mxk0w99IJoAaRquycxtFX/zGKRqFrKrzlmslaZ6ldMzBXbG66kBclv7wL19n
LW6y2OfSINS8sBGGrC8UYJiLaLYXtt2LqMHiU9xjSyrC6u7/d4PCDZdDdUh7c5Iy
f7GosL1ImiFcBGcoLR/ZopRFL3yfT0TffWgm2h7vPc6Yq/Qu8DOMULW8dp+tRXD/
yjdtRd7StTRfCU1QTJ6Yfu01W60aSNafubqDwADwP1TUhaQrexQiejwsZ4ARYjex
iiVldyNZ50N4Q96DdPxuV0UuJhXOhxn63v03MipQKbqWxVSR4I6BtQIFEhSCwRr1
CO9NW2STedJSwhUi0Bw5/4IzLF6lsDFkZ6CCTuLjDJPCu9ZsNFH7I3o595SpuW5m
IEB/BbcGIgrVuilUEyly9G7kHDWYIvTF2CUw7W8ZPc3M79juppwrieR4H2r/awt7
jlwnogVHtTCsmyJdqAS7/vrzQcxP5EVXBS0ataGbnQlKF4gEdbfmlvYk5dfrYl7n
+gNFtemE++5k6wLQM3rX7DkBsQI9DZktrENSgk7zBQti4aRHtk5uTmh1ZMLGQ5C1
tjuB0vGrAtTnIIZTOokJGlgFHZFw2Qk/M2OFpKV+rdm/h5IT1Yz7ElZ388jjqbn6
BU0in/6kHSTG6G8KvpmcPyIKlYKLlCf7tkWRYGkdGpgqNFr1QBx0/W29+uPCMAPe
ClMZtDAj1EY0L58dAE5kerO6fH2GEKqjthC4ffHBFt3MDBPTLd/h7PJ5y6uYydKz
TQpmHDhqlk+outfh/qlT66InjRikV1nsD8cb8KLREYMkig2QKY8koQTXZUAF2SZl
RBIK8BaRSTcLrpvuhKg4n40Qy5JDzd9aPeXi2uAqIjWOc+0SUXzGbF/LTMTV/733
1W7fsgVTOM1BpiIkGeNF/lDwk1X0MPCBheyBPFW1XMpQF2B4S9pLooULX6BkCtRH
7OSnirkEOGH8t7X+fdNGSgoJLerRjjpwt5spj9whcI4ASq+TwaE+MXkkRnZTlpI7
vO3DRIK5tDh8KiTFaKtptEpG49Ph2w6NTrGdec4ppBt7HSlq1mxTHc2ONR8un+W4
VjgNig5PD0Xxs+T58hpXlVKaHs9aHQknht4L4iSikehAl50UwfnVVYd+FH2ZLVql
8URdiLMCV9i23PYdJUnDR/BuDKZbzhZja4fH1l02/nXkgEFt5s9JXuVM1DiCGIlr
3m+K/OnQ6fLXAMsj/yrft08dpv8qAlNneVkp3M0/noi1jOlQHqZ6S4UtT2Ot4lfZ
m0647clMwjJfFuhI6JGywqHwEN7B2JtOuU6ASXC1U10aAquwheLnBRkbBWrSgEiR
5hI4oMi9TP2Itc6Z8AR84cZ95PuI6+kG3502jE2wsRcMjWvRO7Osz+lPcb0CTrik
T1L3JKNGMCTy/VR23eyNZxMBI5a20JFXHvDIz1E+7J8yzssM8c6KUrkgeeC14rQE
/QPS/e1I2xqnIH/x4HOLp6WCxON077lK02hKqwf/o4Wqfwh4CEEAy9Iffh3TGfbi
N8+dYM2of52YVzT1044xCj3TId/2Vc1QG3U5p/dzigNRj6R/nEubmA696RRsYMNi
+5mGMDOg4cwpofTAuWG9ryQI5bf1+OviBoa3MOzjVtDJ+JO+VPtVDPbu4fpgX9sL
Ha7lf/0uOAMlTeSa7KiZG6KKsoe7+PSJVS7L96cLrlcHKJx1/wBBOUcjU11mCCC4
J5KZJMmg0W+VagtlxowN9Utdd9CHXwEg7xRoPxVk+1gLW1fLi0moEtSa5m2kZZpM
IfBpOSU6rFlLdT80RUdx9z3UcORU64dNm0cyMSHcnycgf1cvLuAAAuk+r4Ejcegs
ae1A9dWRmHzoBXg2/2rIVeCvgLbH6M9CScNDnNGJ+U4HtoxQ84HLQSmg5bQBNqMH
Jy93xhh6RuNsxw0nioWh8LNa7LkNqgZm+79y8pRMYBx0dNHFKBPcIfZZ9D1KD6AW
HuQopegMLd6c/D/tM40kZ4kENSvdBKAhgYANSgi7pf1ALkKBIZs5U64f+XtpejOy
S4DLsvkQNrxNV0iVyy9vDxdeGyhHA8ltNhf0HFgpChC5F5Q0F7SOQ5P9VD74QB5k
fNgQDz0b2z5Ds18ZgiZu3oG/QAg69U/QMc96O9cc3ZBI7/iu3h/nUecso8qNI1wM
BIBxj48IRHwue9bdGnsEYkUv/56zf6nc9KCoafLf1LnyRtfdtHP1d8toRWxyjYiP
YpYV/TmVBzh+i+e/Ahu7aPeRyBp5mOoJ9vQ9C5WKl+M=
`protect END_PROTECTED
