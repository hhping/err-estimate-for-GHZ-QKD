`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zf2//ipw0yoqxW0foAVimfKdlemWj5KDc2y0EOVOWki/j1vGqr5oFqC0P9mZy0to
ZxLYjWd1y+b+kT+rucydIKjVx06dZKyuo5MLg+rZz3oP2Krq04M0BqbjBlZHZKXw
QSkx2fAl1pLzC5/CuT6RgrfiRy96nPtQAiG7zDqJGwDEgBhlkkEuY8PNUcCABbeu
LBg21Vp7xJMuaM9ndMM2Ys+MoS+Fl4pEIeamXpM24+iFp3QoiY2Ajr/X70r4D31S
917cT1x5o0ycECDgBX5TeXxl7yilM061clvgCSVgS8QUAshs1HiZP9GvD88SNW3u
ep+uTa4pd3uXdp/b6Yc5TPgNGNaEl2XvEsCF2pUJ8JJX3SpHZqNVHbMJoCp8gVg/
yQ9eyPtQCb6Ox3bbg5tUzhp6a7EKM3ids2Y811DvgNu7kzTBEQJE+noHeNtcp4cf
f4BB8M//lVk80e43H1T/oVpSLI51ed9skpLhMqk5/9BpZJKjHClhNqC5ymN3yO50
G4Pe8ukjbGrp2u9M4AEFF7xqoMF2+07Kk4LZ5UKl/p6kFQoh4exgm8N44yZ3nrnX
yXcRAf2MROJUTC3uF0l4pdawBACRcuaGGuKtL0Csxi2gxqv81iR9xt3MCb0ZamO7
6yFpuCTsmUGOOBYprHAB+jEFLmXyAtStD6R5LAdCklQlD+3oND8kUisIbF5UY4mH
dnAAEDb29EfSCJBFeTEfMQz/0gOWZkNBXFwmIszKXxsVE8wB4TBq2coVvSE/upom
LkF3BXri/ec7OkZQEUbKHVC/WSaI9x4o/g7yK3UldQvf6DWu6hpIGvwHfWCKQxMa
9QeSieEhPGAXpomg1c7izWvQnztMlHjfj6iyTE/rgK5J/hJOpkLNAt3i8tU1xMgp
PAw/nqgmNZGNdRHXrUFHSUjhz2OzfOWkUwKngVLw62L/sZliI4vnUY3oeO6COKj5
u65b/qiUgFox0vbPCOLxWLRB/0C2j/7WaYeJDtP3ixc=
`protect END_PROTECTED
