`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTckh1prJpWmXHu14d76c/9kFyZ9Yy/eLT+V/0zV63oRXP30WaVOT9JuojWmNp27
rdP1Elxlhkis9qv5s3gjlzcpHk00X/40Kg5/Kk8sVZ6226ipoY+1aM8QGjVy13vI
r1oT2Xs8CWur+XHW1agZXkepQD3FCvk20RI4gNwFKtAyOWyY19w5ln+aNoVcahj8
xNlh/a1aCdbvukjJplYHslyTB6VR8fEH4phG03q3FV86YF0a9qoEJBgAaYzRYv0D
opAD06gSm5u++W6q7+LJzQvr8PHYnBEyUhmkIfX44jQf5xJmUJCr1Mxr5gCFsUaQ
bB0KEHB15xJ+uw8SbYdfB8KuWc0oEy/quxw5R0bjjDtWTyW1pIeTvhmlxLiAUyeO
2Q/Ay8ReNPFW/maMNVeGNdcfM4amULISAz8qx7vipBCSxYLawlPCs8YbmfdqaFCY
h4tsnarxjf0n8Jm5jrkUFaNgSychpqlbZ2+cBs1t74C4Y03JE13Mx7iF6UdeoJPy
MUHxDSfHsElh2mCl2crB6P8Sb31VNXAYgv2eOq5gA821a0D0+rtLvPRTU1jeS0E6
wTK9CFCju7EpGJNyU8Pq4+enCvKGljqkFd/jHVFDE3Zf4ZudOviyIzdiiadl/zJX
errNdPvPGt/tYP8OMLS+S6CSwHTYnPRKindi2aawvjqcHT6ofhyOH8GjkgI2nqPf
ZGxKYf+LlwU8go08k56uKEO+RDA76Cg5WHWSy/b+19V+O4GxsMWaAbt4KNbVyb9P
MAZxvZZp6CqxVWNV9oOijSNo9JFXyXp209b1wM5VzucaL/5NEkXvBi5M0cKtZkVs
OcD0KoqC0h4VD5RKATAiJ/6IETZIvOKoeqe6WKJFX4CcX/VEvWosad+Qv6Fz1JU7
fAyNKiIysBJ4xH/v/xU5N7hW0QPbbd7gPQkJVy+70bG1Ktjxwx0cCmf92+ndggpb
Z1Um8qsgWzxy7A408D6E1AO6EcpwdPN8T9yabJSMT8IU3lHjPE6zNgAmPubI6fxB
`protect END_PROTECTED
