`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BqseT7+keUVyxnd3J59BjR+F8Yfqjs+Uf+gFYfHq0uZ4tU4KXH6cdSDMoSmY+nEm
wqPtDQfqzcDozgqXp/w91By6LwDENsltysi1pqviZzYcq+EnUBrcOdVbNJns9Zt8
yQQOhuHdEMki0DIaUjxsiwuPd6yt4AanpOXSe7g2VUEJ7LXZ50w9QeDGzhQ9dTS8
5SDwmoj9gPAs47uVrORjMxP7VuexXuGd87ZSr8i9SGHniE+qzVsP/W2OsauLTBFj
tWlRyzXo4hRRDJmHl7MBsIAe8lmZeNlCDLHxfRn0qvXXAKtLjvFGdta04BzDuvyn
YNrV0OymCQDU0YKeonfbWXZjnAlUJ3CoUfS2rcDmDkAQ/crOMtGmeTx+gL9uyrjo
j8f3qGGAG3XH4vdcQtzMAOdm25T6UOM6AYsU80a98fIk848J/g+IdZzMQX3an7DU
9UDzOcSlRBywSBNhi9Tltj5DCRHq9JR+vMdn1D5XDUUEyscOiyITyaWlyuiY5ZCV
ETKoGsW69doq+kXk5tymXJ+UbJTD/hQbGVQGmVQp+108j5TZs5LKCsW705wcCYZv
PICZ9XxI+MJjnkstvLcPf0b1a+TWGMF6x3YEaLdn3Q0Rlu0s/IZ+9fIsh8M9PUyH
SvMqCNjk4gWCOdAwiWGg+leVcqITgECSCiCzFUnK2aNPwL11yq3U3WIOHHhEv0r+
GDUz9khBU4ScfRuSyQ1XTdqsdIQPYNfOKZbMeCo5lOl0p3N3PPLR8pI1tecEGpVO
VKp/6WyPdBnL3VUVHK3pSKHyzbolZABVcLRPLx55II3slf48f0mf7AYqkRORP7tX
Qv1ElwbNyCJ7B0pVSnVLrA0qcDvR5vlpytL0ZVOZecXDj9R2zDoQjYr+UJPyWL2T
mmSIaES1mG6Gv48QIie88tmOZsTgQkybST6fOQ0Q3pS+ljY/6AslclGOTjBqiq9c
bEAB6V7Oav0czyhU/KhNoPFdws8PkDIoHZEuGbPm6qzJ08DLOF1JkOLoOTbMX9WC
KInru9xOlWOYpLhjB21mlksjU0SxT5A2ORqMbV+dTU/izG8JI8ovYvU4Nw3DCvvH
wXX2h67SkqR35bJDus48KYcrgqt0lh85Ji/hSgGeSFdOKopNTyHKyr2DXtlmDWD2
pfFP+6IanNEtMqDnSoo5QikQwurkC3kivG1zgn1a8l1ivhNep5NHIozP+MLjYQgg
S7s4AmokjbBEMECSlK3Ejg3kuwWrBFrytmWykf9xsg6iVRK8lCP9zCjkCs9ZuI0S
bWvSbHbVYLdSqEmwJzDmKCkIWcnZmBy3gvyqvNyMc7bK0KzRNWOZasecunTlVySU
z01gcKN5HXZsXaK+Hu7OB0Gi3Ci0Ivj7FwqpzSaeZQI99vfuwFuUttpekhx/1tN1
4dSQ2D4XqC4Ri2G6nYWIFepiBpJqP2QOgx81qtnVc9YGbkfpGd/8Nb2mO5pfQMO+
Muy6RLwwWqA5cMaXnHeLj0E2qiLTfBjXIPS/RlOrXGvQ/HpLYzgJuxrSr1EUIslG
AEm9DNVRT79Vxa8x8PALZMjqwGLl8O0wg9GJZlVGXjWnhK1CCeJ8Ed9cFsmIZcip
Cr81QZgbhgur9LNhEELQvQ==
`protect END_PROTECTED
