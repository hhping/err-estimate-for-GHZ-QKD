`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0MOTcNSf/5wuNHPvuka+Ppr5LNhSzqTtG/Cjj8blB9CALFOlbX9luMxAe27Zhmb
5vL76prsG2dH/RRv4p51IUvR6kFEHdyCGQczP55sKD4UjBsoybenigS6q6KBgQ3b
pjnmHKU8zri4nWTwRi1V5Zv3xfhAtwP91PPRQOPdtrQLX/FKRIX126+uRVhJYwIo
NTqOfzwsqvgSrB02VI1etyqUEZWo32jzdx9SIYcYR+TUhqK3XyaWJkPwG9E/puQI
54+rxSSEga2IgqFGxKfh1WUuD0vDxRYAPygTQjhImAxncUYZiHq0emTaMQvYKgmh
IUkpiUmTQYQ7ZZ7HQH9REF3bluqOy0ooKezshcvxfAaPdsvV+JRryqQBH8awQtNP
sOaj86TlbtpUn4RaIMRP44wce84WClWvHYzpTldsFqgik4KRM3pGSHChx8vd3YpG
k2mMb4C2S6xSslG6Vu+6hBotXPBFl747cHXKJhuE/nPIpwJWAa1kwizUtciHWTC+
yjc2mkG6kOSomaJIBubQsM8rFumtXdLhbCkRLyJzD8xqbIwpUT58MHe1klQp7D6k
n+7vqES997YTWFWzftAjOaTSe3H/p2+RCLiiVUgXr1DcfWwhH2cxYgqqmMyX4p0p
ssQVE871LxF5wUYoBSWWDWnAGxRUQvugbtFns8nG/HelY3GtOoBZ1CUiOkdyGQz+
`protect END_PROTECTED
