`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJLT5tkH2oMQb0tKN7cT+Zihn+2RXM1+UWm948sokFhh7yCA1E4o8soP+4rO70ZW
TiGuFLQ+FoBXkQzYU846GbSjkgRVDAAXpXMyz5UEJB1HXoB708Tmb5ndZm+oOCsn
PwxOl7RP03lXFtWHfGJX7wmEzjx9m/YSskES85DFZfSTjynSNGLBLXQp4fsUCqfH
wZti1q8+1mEANLT3DSWYfbdONYTAr/GMtFhIJZOcZQK7RI56qDvMMD1PdDF854tt
f24d4GnaVECIBSyRqQm2tAogOFq1RXgPQv8CkUt0uymUdbXDYXWOQ/DCcXk3lHK+
E7CUbJfJpIH9Ko+cHYw7K6TOGJ/4WD3NrqXULBjMLtOMFLwoaiIXtx8089kmA6TA
NbAp9loiEP5oxIas1x0yEwvA1AFcS7PgXCyee5u4Pwp3uyn1b/xv6j0vFe7EibGj
7W3EfWSNeGgeH8Fxpi5sVE5K8mqh8NgVwkZfD6Xu9N/jmA/kyRYMSu3IrKpwAeje
`protect END_PROTECTED
