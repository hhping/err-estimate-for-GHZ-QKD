`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1iDFrrYy+Oxg8ZWuVvb0tVYOJ3dq/e1fi4j/ASjkNBtOyijG+5PDdW/Ubl1a297
YBye1vCy3VAikqciz3YkFAVOSLiURDxmeKZIAZj8oZ/33wF0GOrkuDbY6ynkbJ8e
iy5KtKvsDDRPE8JdaPzwdH37IGQLqkAceZ0glpgcHIfrcdGVIsrCGXUhfysDw9bY
FG1/2Bb6NwkIb+5akRHGRaYo4FX5v6AoHur22JJzdNPSwfH9RlDS/jylFgmbirL6
mMORr85IQxaXjVdYWFqFnh9bofQvHRWTAXmqGOTLav8KmP6W/BBt3r3uPxqJyTg+
ey36FmneB2w2/hDpFfTk6qI8V6FrAQWHSZykQguxwYXF6EVU2oTGHiYNwQIk3HSZ
LREEB1Pc1FiQuR7z52OdtacaHBYsLu+HFeKbZZRDdgobTq7eSlV82wYLpbS+jXqx
eI0D/Z1UuutIQnm8rhHIVzNd3NglDwDgZpeemaDA4XEwcZifsrruhjv8AkJX0CCw
D+ULQebvjhdTfZZPMrPOE62TtGTvQ3TFc8uu2lIuBc3x0PzrUCLJZbTIpz7OjJSL
kDkDLuK15fw4eyMrOz4GQxw+GmwDknBYAsps0nlhyqllZwm5wm15g3lCo97ErfA5
VEGe319UqICt/MSTTeIy8KcEp6iktZf5gcm0CHXad+Z1hllwQ0WVzRbsrRYYjWnz
DCBbCOJ+BSk3NjcPaEyd944Nj4KrHPfjoJG/zIe7q+WQW5kbQPbQ4JHxIq6bl964
VRxHUa85fHWMadcs73jr8u4o1BE7GS80n4HES5R5SGeRQcGxIDO0wrXY3u0OZUwo
VKMO6GZy/AP/OEMXbsKvz4fB7uAEFN8wkDIO7YthCFJaZyFxYzCK740abq1aFNmD
13W9TA5rK2SyqnvLGO+HkXKuJsbM2qbbDslvNi/SwAp78uRZokDYHqSDPxWab63G
c3TWAY+NFFmYl2mOczKIF+C5zwriZ4TKsHjUU5qTrmEpt01jNzure2AdvZL3rzxn
X0Si1JCuvkLz/xKkT4gcqxCfcjk9wTFSEg9pkccuvREDDGFYyNjDpZoRUgRFUP+C
1mWH/+uI7UFQcmrCBeuzOsfiFGx560g4dttAYC0cX4h2xsbi0o0Fk6X09KPZkyZp
Q+5ZlOUhtNeigse4jBAvNxk2x9VjGzXaB9HQWJ1xeW0biuSZo7TvOe0Yra8+Zlhz
lWGAVzMsdFrNahkuvX9NEsST4CWPYu1LNb2uLouQv4HiQ2EV2lqIAjef71ZkfcIB
FAQnMVTObkVNjyGitNcPmp+9hFPkeDoeX4TWGT8M50I=
`protect END_PROTECTED
