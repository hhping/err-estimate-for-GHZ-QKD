`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RHqoIFT60Wwl949BAUNEP1mgb8eaJy3qZu9wpRQgEscUG5Gie9vcGIFqksDif9Me
BW3wObAAtai/NMQd0xoypkYUc+LRiRi/MLv9uf3+Bn7xbhKcHMSJfGaNDx85myc6
rwxohHq6hRfsKa0gevTq7S1WeJB7/zbiNC03v58Jw4JEyJR4TOlH79MKDTaDNmlL
7e9DiweAmmkHZtABGyHGe0WMAZETcMDL4960gII0GIip4IkcbLpU9qzdUL2ih16V
rt8kpmhBp4wrrtNN8PcDXciQvO+YjQJJyQMGvRpdTkrYGkebpb87Q+Mcp1mTRGlN
O9igYncvqbqge9Tfa/j2vUKijK04nuic3dH1QC6y1xoB3UM5TYjWQ4rWRW07QE68
hxpd0lkOfRuLQJCQA831jxG4z4CXFcVWmb8uUsGJYysqmROQ1WGPxX1bVabuE44F
JXJkXLiE5AjqTUyl0VBjVmiilnm5J1f48f1NyRYPBbqGRjJkt5r/MXJfBhHrwMKU
s35W2/zBtHr+VHfvfmTu+3nw9xqZbgpq5Pg8V3S+W7NUheVkiVqnWBxQD+H+Q3qB
A38Y7NMV2yZpKl8OZsP/Mcv0WaJMfd4gWtwcoU+0AjSy+n/cA6f12EEupILK0Kjd
5IQiNkIUkXkb4oX64+uGNs4Exhs3qVHiGRFXwfv5GCjcl5IUCIPCNsp3Z/63CiA4
z8T/I4C1m2ar5Q2rnAjhSiM7swmDIiYAz14Gw5lwVWGSPviKOqXK1BGdTxb6Ai+r
Y6CjzPsB25kyLarNxqy9VTNPTUKUR/aFYffqu84Uatq4JX0Om4dUrUbv1j5Wdm6c
hCUdnU0AUG8BNUmgjFOYh3XrZRnOEHwTITJ4Byn2h9MXWBKzmUR4ciMthrS2HjPj
F4WKslvn6clEGhwjTVEe5VNpdwmWCpen74XncbLzOlp700gWinMVUcw0V7Siz82G
aDLKdLG0mrNhZ1RiEyCgNTacHDnvb566J58Th7tuMZ3+FAcAIZ8KCprYIpvIZjJ1
hcN7ZNRw2Xwu/rdNoz29EsGIKDIpioC1ZKPirKtEvf+/pVRueWUio0enhyQHNEuN
BBT0aPcPIfu8dTm3GDLrxCK7LLzGPNtDbIyMBqXw7DDsbeWndxbGvyr8STOwfN0j
qE53I3So2B4RnbUoIXUVWagtL62PbH11suRjXp5xfZuU+/CDFY/xPoutzBs6/Jjj
yvGZk8puCm/v4vzrUEUm7I0fDOSLj4M6sIxPwtdGyITuV377kWjJXjZhBbcCb2Vs
Btw/5wGv1S3nLntup5+094w+ws7c2kGjZ0fLy84qwUzNRCn3ZBnqSz4KwJuV/xe4
G2pxl2whBRhdOPIBeFIUIhOf5gTo02cR3fRQ/5zziqJpgwQXxggq89qn0YeyoKuy
tZS10JW0pnNBwW2vhN0GKVEu1teJGAXwVet1JrZ4u6npXGmAEewEdu4eFswpbIbj
B0mz80u0Fpb/00auurdhr2QWTe9HhzKjMqXPtbPjsA9AdY0LDrBrTJShsW6bDji3
gsaZygbEd2SNyZOuNuYJu1FuX8KCuREFFb7EXYjoTu0iUPFkGe8CwxifCZ2xN6CA
v0SjnKYFvro9VHFxukgIp6mr2W12fhMVQ3+GbY6r5UzDmMTOrDFNUXcpZj4VS4lw
48rf3W5hsmJ/wvanUJTeDxuFZMMHGjb1eXBYosNpDWrEpWvbUR5MIIhEOQrfLGxD
MsmBgcStKHLJiD1IT4Ri4iFAaQCqHYQkCedsHnkFKP+6rPB0nF5oj+r72w3bHmb3
ah59Z3v4eL2wKQwq77x3lbdvXomHpCmGJEwg6WZzDD+XTzXsXrBURoPM9oubOm7q
IVR4M+iULlPElCgu1xPo8atLmvZvDQlOsE8pY29BM1WXEuO2IK7Y7AkFp1nRGhSZ
EhtYEACLRlCddB141UyWM5/O4JbsoQTD8b/O44i0oPHJgd7SGk7D+Y7AOZRWAQou
qJAFHaQ3QArvU+7Nyf4FFIzTOIB/5t1K0DqK0WIGez4ItYoIoMfF/yduVs6ZtWPI
6zcNELqmoVg/uiTICorfEofOfmDBCMTaJn81xKLcbkvUlpVXsLUKPXDXWLZzeniw
A5EYPmUOD74gyCXhWaAqPdZiRQ/JrJriWKvAiXwLeLwqgCg6VgFwpiTNv+AsY1KS
MPo0gIBkjgVjHb2vDKAwdSwZ3eKuMZBs7Wt7QC5ghR/AVnSqS5wQoi9xCoZ+8Syx
OOk/ZGLzi7gwqnYiZGUip7vm2D4M/IjgsdwHqpI/RugDmRFSZwYpyUcPyL2QegG4
nC8rqMeilOUjCDjHw6HMJCrAZiEHPVunFxNv3Z9WAF0pdylGSBeCCQrs3eQPWYRD
vDgnZdD+xVY0hRrWovTTFi/rlqOt+KUq8F4kGPN+MeppEUE1FTHVpJAx2puOHcjt
77wsbwcnqrv4y4WCFBVZld2Ofvp/PX5/nqMcX3Iw9G9rfbTt7WJ1s8hG8mgP3Vh1
Bzf3M663R2lzFwRBArr8OlFgS1UmTRtu0w9496BhAU3HrgZ/vr68v3ROZh21ymT9
pwGWw1Sji1+PbReroqWE8Cp4zRV6/aYm+Lk4S6qyYJm1LW6xBLnuYk0D/1C6Jx3t
SW2y0SdxXqPEJ5E3J+Uz3snp24SF2bYYbn6raWGPkHWxUtQoxn+rKsY3sINsCDna
AqvY+4hkprWAmsl1uPTMvEl+dH5FsZZSDGiP78F2F+l2XPIw14kxZCpjYwzHjUWh
cDhIYdslwiAEUF0NY/i6SIH02h4oTuU1rsX0L6HI1JGvLHZ2/moPC9zCy4/GVtVq
OdBSY974PEk7cDTcB5Wn6/ndOCXBOmPMWB7Xn6EfzTlrnC2fGuODh+Do6U4UiIUb
2YftqFuBO4fDRQdvVsDrPiTY4Iyk5pCsv/DBnGo5Fncl5Jc1UMhXlKNY6GTPTOEN
lyJFfYx/iXdF7HSSqHK4PXD9i2dejZBOfiLFnwkjido=
`protect END_PROTECTED
