`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9Biq7SnYPjBUUjSRGtYBrwolORyTDBJd5ihOKmujUTeSYtFyjc7uythKYdtDnGJ
AgJU3ywXSs09HCllfPZ3W+Kq6bBLebXR2NSiCzNP12O4rCC5u2SAHrpyVegUrbEw
DeqhPpAdKAu7H32VolQZXJY1CK4ZMMsn2E1FwO4GXsW9WH0LynEH2mqfdD5UZW+k
j4q3ty8/Dkrs+2gdC+COyVi9AXNfST/8Nmg/ZngoX3CKfAXYfW3YyIqMkVazHAS7
/rCwk3t9tfVvrkA5JNmBLsvOlyEol5HUtakA0kUGxyq22QlXn4W81wMpITJnsdOJ
qn5Sjgat/UgT0PuSPWoLdDnVpQM1Y9DBf4jarX4YtKxGEqTy2RyVqRD3oP+ecewI
hzbluJ0YttOcCQy7aQk7ddQGGD8aaEDaHQfAPQ3kO982CrLis16MWQK0p6Et1A+u
jmTzsCm0pIawgStlMP98Lc+RyOTnpctEmX1v/6YPYPdCPTobCa6YKf96/tYI7zzp
WanxKK4BCODhME4Z8EdMIbpGrZCpjvh3GZkzaJiYzXAPuQe9O6EZPReUdApbYHm9
HbzNGMP0A3tZy4ih+W0pXZMgIavnW92dAFNez8tdnSPA5pvcwdDux5zSupnvI9jb
anFCE0LqhlT6B9umP1Cyo7fwy9JeEs1W4+V2Mjd6pyRJA2PJ6RPhdX22BqiPc0OU
uudvZugmiNM1/GHwHQNzQ3y1lBkichKNQiP4bjZ59BAl138un5/6F/87XmUOlIxO
h9Ds1HqOahezNBn+8zHLfsDaz14AK87pQxK8d4iXlOdTVX9iUPSKazyiqM6/ZGJy
JhndkqD5p1YGfCyomB9xyVP6NjOjWUXlFYrxLF+iwUnFMBJ4WC0bx0nPppqF1oga
fkozAhcL6KjY1NAtuK5cPw==
`protect END_PROTECTED
