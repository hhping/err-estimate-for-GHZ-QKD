`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YbpsBDrEqwBF6a3DGTmzA62FeNMDiW+dHwKSrAiWgcNE3gha0H1y90fy2h96qhF/
OOQAL5GvmDIHUuaqxGsPQ0oiNlx8DNhSH6QCQnDJ7od0N4CM9os7iyY41i0Yn6h/
70HfXwHTYe+HdvAwyHt1IyIudkurUYEjYjQ0l8tsLNDMukASzQTEHeBIrDd6Z39d
iudklwlWukQ82U2yzWssNq5b0sH8vQayQMYgJtUGoydplVro9B7JAuxXTk3/Bs8p
hwFeXWKq55eCu6ssmGQVjrztZNpqyoThUhoy1vQdMdKpucvwRIidlQwbd7rTn8cd
7acf1rs/FlOal8jGv/ZCdcJIAu3sP3L8CMbPRNWJggH1Cb8TwRdR3oBpgPzm/TQq
7twqOQopGh9EIZ3J8+t3YxfSLyb7TVZaQ4NIFwxuTZQfqLLbspQvSFgs2hl+8Bm4
7K/2bhFzgdnOWRzHLpxSIAvdS3ARGIS4FBQUPXBq17TzoGFb5/6MpiMqhA31FZsT
1GGlM0oXT5QQOrqWJAg6jP/+/lOcfz5sHJHnSC46nvstvYBLz5oeLDzTm/0b+Aie
xJ7nYPiVcSaf6w2efBRrM68YNZW31HCP6aICNjmf1e21+fRvskqmF3B213rbfQVc
NBkXAQG/u4Cv30SkCfdOMTarfKP1z84WiYylgx1MgRghwZKQE+5G3pP1oRkZBWi5
SmdZv8hQ0D0xvQ5zpt+Pw2cFYYIFQHsef3rG9AFHkEjYUyQ07IWhrKyDf1CNiAH9
fQUEqPOwjZpgrgTB+U8BFHawA3Zkq7q/mSWDBQ9k4KkqALQAZ5q4BYYB5sIv6pxV
s7x6upt/eGc/jRLyVxYx9JeW3nSHgRB3jGzaYcb+EGLmWGRS3vUyVEIh4Uq/7sQZ
jbZ2+bj7GlYRlfP2P+oh1Wpl2D1OzjBNHAOeJTQ6KgLHw8iboxkOV/CXoycInUZ+
rO8QqL+cf4hWmFqhgr+zBudFmzDZv2rnadwTFo8AfwCTCHgl2bY8feAZGsSY0yh2
VuvXbFmwjpv0gHEZmOYd2eYlSPWZt/TmKog8HAsBGhp5Av+XQ5BGAKHeK3AC3Pra
xkO4aSq0h5P1ijsLSTBlfy5qjfLN01LNJ5Q10jIlSWk159c8/NBkt1JVoZxI0o+H
TVzr15N3wakN6aXhOImiGjNFTKS72RkAFJ9LvDBvra+WS9aXOxNBeQzxXp7SrJsE
1iyqS7yNkVfIdc4F107qjR5XX1+y4WecGIKI5EPab0R45IDcyQK4NwlngUPKVLEJ
KNiOqEh60esOAuaaX4sN90YPFLnPkb9FpP7sPa6QYDeDagKPIU8QWTiwI55LJZHD
Y7lM6Lb7AKDg64wzvNC/BGAjChtjUMunvukyMZTlnPXlKrvqL8dU/Q6kPsZ8/OQX
gZWWhZIe0W8w61CYuR39o2cdMVNN5oZAWcRpI5+HViLvp97QxWJmV7RzPTS+QaMK
cMzKfH6/RfAtstJTQez8dT1hGzDp7dDn4bGRPrBEjm30nIlngovtH8TfjDxb73+J
Rnuwe3ZOjY4lYnwoKEsNYLnj8HvOZCtxqAKDofekhy1LsdVV5+bALKayLyjkH598
ToIK7jAg8m8TxRjvffM9mqC3q7RAHMvBpCgc/e7BsTtVZsjK3TmQQpNiD1kIsuMs
E413IDChZY06n6hNg3eiq6LB7gkDHZLAiOxbFplKqwRch90SE7s5gBNX3lZupQQK
D8g7NnU+wneDQLGqWbUI/D3p4meUB1Zpvh5FZuCvjC1EW5suu6y+9VCUZVTVyMCe
IoE0/36DLAmIXj/l8Gc8xid5JN6ZdyQjvolaNMJPJxtkR8gclKhn7Jev7orqOhJL
HtLdFHkQWWSuf5Bj1Qj6eRrfUyAZ+iNNO7OfO9NFzFRE/CmqeyrqfPJgjtPfHELX
xFzFf+04d4DoccFgbny5Ugeh1aqsl2OTowtLWZ+HHoKyM0OqAac9lSYk0BxJL7Ww
rUq+DuiwgrKEYNGOlFEGiEPrvRTko8hSCV7bx/cA+z3KxAGXL1qmGjfL/UKdbV73
tbACiiPuETT98EixkASHt0VlnKD36WqnW0p/K4FE35/Gl4cdqXsId0i3ZuIyDOio
H9tpY8oUNDdNly4Wt1P5d/xbcL+eSE63hZAxRceS8ctqos9rrQ97SFCLgw4sb11M
20C0i1WlxuIZysqiak11DjzQ0ja7JjhE/DH34wIUdDoe/chlS203g9q+Rl3vy8cj
NsvMKtRBTdBK90g2OXKcoG94d6i2MpEC6FFMmtEseCEUUZV8bEtKEfd5m7G9Mg/3
VS7kFyNueYCQAlRoDc+QpG2xScV6uPx/zELLWAYGu7jcabZoxbNv9K/Okg9vza96
5R9cAtpBdCbAcao7KRj5yY3xLZQtIZ1W5VSfGT5IuNIYwzZs9U8Sfpg7ftzxnpnT
kWFU0vGcYhXWisHYtPFfsYVpOGQyFbcgB8jw0Iv6rK5vPyR2ZfMM8bAYIQfhtasD
m+gtAA4cWbOVll8nIiurjTfKdnF1y8ccYfxxvBckhoZTPDYHJp/IucJrMY6CsLA/
B/MV94A+BFCALUEvcDF/U3YUARQGM8c3cgRbHCVzkd4vtr1pRtBtbrJcgoqhQNor
G6U1d2iego+WXTJ7u2miscKHKbQ+aMhJfn0vpuxFWZga2kXg7W6HmSTibwtYoNSp
t4XEXeQBx14Ipt7pLQ325UKYUObazD3OHeOqI81YM0h1bcT+tKmFhIMXYHLWDAO/
bsWcB0p70XaDVk8mL49HhLgs7XnKnC17uo2mLSWHgte9URxUGIqLZtRziIZbIS+S
dcvAsCEnaf6PdT+9Ec7NoQ6BybkjofBwqgiTc7fXjH8XqLM0+A1LaJjIYQLFhceF
0uDbyzBJQzqNcFD94siEuM8exeSAJAVNvKOCUynff3Ybl/DghWL7mUvo/9AkCbqP
jcgMOqfAzYeRLqPgqyRAoANdjHPsOzwoJ15KvOuETEKYp9M9CTbYq63MJ2wFIrar
/poaWWwjrNRt8qfnCfC0DWD/0sVtV+RDHJ7yC5jrUAJTyoCkQcjlHuOlLcVvfp1U
SJD50+0oJtU94aGYWec5Ze/FzbgyQqhzvlJskWZdZQNawS01LK2AeKrEeSe3/XwX
i7AVlhpx/Qhd3LVZ4/ZixLFdwuHMMJWwCZ5NiZ21P77SEAsT6aBd/P4pE1Hpp+Jk
/yFR1MlOxE6j+CjsNXRURIcuk20zqlCraCf19e3aARtFrarad+2Ev+ikggLAzTRj
c43aIsgmMisu89sAQR6hN5+rYlOdoSRxyNLN9kAZls51pD2T1Dy/2DEkIQyHcGOa
e9xBoHleu8NCLeQXOKJMpbzOIcyxEPWFTdqnm/NbK7C4F63Tj3TiTT2yVC8aAsM7
M+EhhVa1RooBV6lZtZZ7stuco4RWAnpO3XieyrI80bfTL7ln2/6ccIuaqNcWQuBB
LnKs4Ffara9jEYY9UY3AbpSqWq+pwMlVi/EJHTh7ZE3RYrgIc/FQldLcGvwEkrR4
WSzZ9wg+SvkwVHE/fFacgii3jhuTfttqAwhtmJ+h5jotXszpJpCKBw1fNwY9Kvdv
V3c6tZ5ujbpU2f3IY4qgCF5J3X43L0Bir+ACEI5LO7im3FzZgaJCuBRnJ568sNTi
RVrWYI3MEr3QzN4os40dHOQRbBSnlgj+ljhrkwQwM/wa1wb5wf4iHBWCCPJWx7tO
KTlE9IM/br7n6kGxc8uuQdAoIJ8UyRDaqPmMCKsMH9BlwuWkhVJvTplxUt2jbVMh
cg84Dr0F2q65OOLa9qkKSV0vHHZheGTwogc8c9WvjyqgR317I6/DwkVnyYr6gY3x
VI1t91GFUKd0ldzfWplCRuAeN+4zoj2G+DhZUypoqI4ZmnPg+KOl9BHspe3o8XUm
I4PAL9wV3A6Z3OKH7y3bieWJK+OIWED9uOI5tT9BwbpyViUIqn3CJTl8+fIdbmd4
lqmtrwDntbMAlWbIeiKI8+W2c04YKPBekXF3xoWmUspgZ0pN/ctMVV1FjC1l8NAg
n4ViQMEsVGt0lCbxhqhVcYcO230aHA1MM8bHDu4hfdiCa7E4xoUTSP3D3xYYY/89
XSRhoR7v2HMRFFCCWSRa/KY3n95ZKm5ryjcLfez5///DXKYGao/TcgmHMF5PjjKK
/ZVoeOXTJlSqK8YyF9w4twly85bGaSC+LX74ZUYpAnnV4StFEN0RL2Y1B8F2dwzI
+RpGegN0t92ecCaGof93o7gVRbBt/3N9z3Yh5egsCyhx86a5H/8LBPgJCg6aTjpd
wP5N3gpOHYRu5rNTnvyB0Qd56vgxlInnHmy8BJpBYgh+JNm0uCHOXUYthoWqarJb
MuQNWlHgCryK3aST1a4I7GKCt6Dw4bu78LmbgAa8xdBgXH9pfzlNVzHBklS39CR5
n9jbDwJyJFO1p0YPyIntFUU8EngN2KLvgHoRIZKPTRxUvu7RQbfhd3dlOZi7Cdsp
dccqUXl75cQ/xs3Hoa8YTwyd9pWCHMOwqreE1OmRONq/chytdhyQFZW6IWGAZTcd
I25ZokhVBIGDookYtVHtL3KLDTxhG7UBeqY0IMaywkdqMdA0tkI58YiDGyHnmRDN
RzQVPWxvhKi3DdAet10zR6ILgjZKKuah7UYPSKFxQXn/RwB0rpqujeYxo0edSbtE
pKp+Ng4gU2bKPH7k2cZKsa5/MSowwx42uwokXexQhhEdzn66ZBV2Mv9myV0AY0Yr
uZDYSoMlvBy2FRYkBOUQRi7xE2GAa4M9vCaZ1hh0O45MSpcZK/1pIZ/HHnxQkFil
q1zXxrjfRhEeMAOsMoFLrFoaeKg7NFuL/aDkY5Oyi4zXCkI1VUg05cx439g94zAW
8Dqh0Ba6cKxMaThk3yrJkU/t4Dj48ka8e5z/tP45E+pftXk3RkMBtMZvZuUqj5En
5jgVae/bvaBa8dlf9UQma7jCRy9dog/eL0yERz8Zgd+uvrhRErmcrDs4MqupmNdr
tr6lJGphg8hnqUP16HRvrdpWrH+iPgZ9PQWhXy5856rEeokPXo627M6WXUN3ccN3
yBUsxMGobOD43Js9YJ83raWiCGn4xubjgCs+0FWCqv71tlFLz6jFvo/SD6cei5/4
85Q/APQ7eWrmbp1V7hjRdjy5zlhoL9swDauqbvTFT2zthlNsfSi+P76sEiuqtiY9
L/gK35XPVG2b/3uRNvDvDfWKl4if66MoG2s9jG0jZQAZCTq0So6FxKDII3PXFxSH
`protect END_PROTECTED
