`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZVsfWBAvocuOltsHElC32x3fgqO8mxVSBCDvI4ZtryBuxy8KFFi1ls7Z0vGvBW0D
alIGpGTqdlrhOf5U34hmmEw+Ov5dTTM6eTRwfqUgyi6QvURKJNjwHosOhHmnTb4J
nKAmA0JmIhVgf2rOqrKqOvHmqw1CX5ZyVEpyPEo8yo37P9NPTv+2ud/ienBcUpsr
nnhBwxaqNGBhOocs513Mm1h7+ru46XLuTtsPO2JyoPLu3OTyWDkd4mB4NQl2mxqk
p8I8iNNw1Ai4uycOPyaBWP21VwMKYEi4dQ2+fgIYsyWuNnu3dMXnSYOw8M9eo6cV
/Clm36nCT9ys8r7DLCXeRyrQ7Mudpyfd4ewuicD89qc8XlGp33CM2mPJ+HheU69U
ZqQDhmoO6HLKAyY3j1M2EiU7rZgsGkX1ue5hLcI33rB8MeEXw/IZr5nsIUVF3qUh
voWja94Wc+LHbOqSsAqNEg==
`protect END_PROTECTED
