`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viiM7yP4F0JBN8BYrsinknpA3JutLTjxArNv/g/xctrvvIOIb2bWB1FDHxhemhBN
qbMXpCpIIwS46nlHip7ymw54bLvONqBNqTqFkR13tvpmqg2mZg15X9zRcRpZP/Kk
qD+EJ49RbVh0bSWlk17XK7/1K8Yz5USlOcEfWZTqQUw6n2QXLfdJuhdyF7g+z2vL
NOKnUQhM7JFPpfeN+Z8cU36fNdl0pT4N33l4Yj/S58N+Iwsbo1hp6OfRCfE8f8VT
+T2Ko9G7lTohmoBX4vFUMFMsyrZu5yfx3Cojw2l7SsXaz0cgti2TIXFcZHGBBskW
2AzS1K1OT4tBmLQEaySfTPVNQiBoXYjUFB48qSdNjUs45aDODPM6kqNlnWvWRcTr
VPQRwKyt2V+KQUMjPnZHK5LuG5tMDa1lKZQOB57XmBqxePCfTPPZW0BJjcMbo/ww
x9YeD9Fcpp470Ob1ydF1vkjMGZlMRQB1Y0XIxfFn0kwfH987C7nu4AR73xmJYwxD
gHu6bt24Cx0tjFANXHFac6p1cBRYhZnMLiMYgATpoiVrm2y5U/+Lquxy1MiibQOL
gbAM06lA3qKLJ2kTs4mfYcE+vMdJCi6ZsDYa5FftxNL+WZEPYOlimIYKWl+u9rbw
F+SL40N+655Bv/UlQpUlIXg2KTRhPvNDcy5y80G32PesIMNRgBSVCdmzR3T3BKNZ
CmBZ6JV8Ix9JUcwDfGwiuu5hNGptkLp6Syy9V9U2jUAw1sg+SQtyZNOGZu5buXfo
BV1AkvwQavU+P88CJUEqDNtQlBgH8ua2t4flxigirbL1H4iOUiyyqtF2TluKH9aZ
BluH/4oHagRUMhn11YX7ycqQJUf2pzKla7SptYHAOdk9dU10eDZe74Li3omV0lYv
CCxQLNMM/aebx24gl/pVXdSmWQbvCji3xkrWKOt/YNI4WO3vzVk1srEgYMZVaY+7
SOqO2p2wuxwJZ1rtsjXKQGqpziPrtzxdR5mvSuVDnnlN7pLB/CQgS9d9LAf/gzr9
xtFmPiaJ/OPcsPmbzGOksyRfOIhx3/BQAAGFEgBewbN56UZ+wuPmAVpdccW6DUx5
0p6VoV21tIxY/Xi4gZ+tnxlE6MkAcKCxeA70PfKW5RjhulLt3h2TgnzZIggj1yX0
DfthO3fUCFjzdlkNAgBumS+OpyfctP4XNdVCQWr1WrjSM7+Ye+JGkM2F2LE22I9n
98jJfp167Z+FXO5q+GiKdw75dPEdx8tLmHnlXvuvaWbFM72wV0UBw2uwI1rCdWby
ZqfRIGHhoarQP+0r4r9JYudJaOabdAYjdlWLtcjeFr7oRdtznl/Ei1PrW5KwgIiS
7xff+SmF2sxmH9yrzCJTQERhSIuzVF2NtcTa56hd9yKK6L8ODas6Un0KJLIqXjkL
hypL/snzHmoL7b90NlJGC24q+vomBzeTwxBD+/MUdlh40Mh5Ibuupsqdt4olVDcT
Hq+ySIqa92q3rhEz5HTRjeq52JjyfrYYtvzrSdP2piI9cHUBLi/ka2Wimlj5MDu5
dI1i4pZfUVjG9hH3W2AG21Is9LOQGvEHPGvSOh5C4g4a3JJag8er8ONSXbNsg7vn
cmFrtcFV1AKHSX3iIeg14g==
`protect END_PROTECTED
