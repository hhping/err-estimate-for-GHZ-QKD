`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldOnX7RsDclQfHbib5MCIFInwwyZFa94TvYu9uCcKdVpZvCHwtht81884sN5/edn
JyV0luT5Kx8AaFvvtNBmnWftVnUG+VUvyznWL5FZU3zL5+K15zgLeJrZqHZqUV5Q
7rCyTGBmMUV0co3sUaa9qVjQ1k9AC3GUd3ZnbO9/2VrG8Z+EoK9SKTdBlZHN0xrA
ImgQxIeFNmA4VsBv6QznDg==
`protect END_PROTECTED
