`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+VUDVJW2U9aTwc+qzVz8WRZC0uJ2C0L4QVbGydUJcoR96qpMyP8O4xMtDocqfRw
GrVg7RfFoPWa5gpExzZ7w+D6brBzQfyXa2hXVVx7wfBobe+q9ONtSgnZXrUVDodl
x20Oxnhaj21gQZiPv0ZuKrJ3HuawVwFbZ8wU6ar56+7qiTH/6AC/Fui2eoM10Rq3
upap43LG4QFzr6e5S6b8h5gRlBQRL8Y8ERru0XLuIDmPWfhEattUgD4RV5nOSJtl
RmedunyWsi8Ac0F/ao1nZSaThzHTpa/wPq0Bd28xgYjaGca3nWfPqsjpFOcWlUfz
cGIYm8TxGSipvNTysQjIrUV+s/UG0brWMWAZgmw0BsmhN0TDWWddrFf+b/VcyCYh
FbxEFFtMQaL853hS+S4mKw2K0xsFmeqfZx8oNeyCseF8mr65YQBk21Rro6OPLS6h
I77fpzZw8ujDOvti4ztyiyUv3owH2hbqdgwu1ZyN6ds4+HroF2mrGpchELIpg6hL
oVqfnv7HFbsZ5MNgkrMvTS61YmgGjtXtIqGuX4RQfjTzu7T0wcPlCE53x5in3JnS
0GmwcvHp4zdNx3Wuoy8eug==
`protect END_PROTECTED
