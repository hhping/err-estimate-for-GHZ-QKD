`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WaEmyBVozvrBQwBwZXgnWhZIoIgVNqZCyVjycuWf+eTRbIOEXJ4lpvBZrCfMdIp5
HWDceyWepgZHuWGY8XK86DVT/fyDVqrXBUBf9l//crUwD4NH3Ga8M7W8w2TRvW0I
tvS4A0OasJ4gooiVpiX/qHDbLManPq6ArdsT8Q7u1J1QXxb8omkDAnwgSIRB7+DE
at0CqvaDWi1YWvBwAZMgMajJL2JHUUqTjqwrHfI+okqsRRSIUZC1WsquGbuPYCCY
2CV51W586aD8QjKqK4IeXUOGVISUGh2NTkvTmO4F7++PuZCkTeLp58T76kqXaMiK
rygymTlr7dgSo4yMgf7gIdr0ttl/8xlQWao01KQVOGy/qqdr4XkXeltXjUUo29aj
ZM00MWqB+rzmp432rSDsv6sZgoN2HfV8/2KYavFH7XlaBx43jkZScFrMRdzMR2MN
bw1RS/s+awmmLG6yKBfrRitqZzyt8xQ2tlMtmVmWs7RPqSWYOOmg7k63ZIbPWKJQ
Odp05IFBWg5JJYUAshdpdIKocxlObQSwD/EJfgD5IWmbYRU9NCPrbZT1vyRE3Q0d
KKUJvLoeRKbm36CwzTjZRdUdjsJ3BxdtuhVGFezEKysMNr4FIcX98JsiJG6/g1w8
zzdSHHx/YYtpM0NGFvO1EA1IR59A+CTiO2f9K4hnLpgPYCHXzpSMwCVBk6s9ghD/
lR7yo9mEYoV43afv05Q317+ack2LVkS3G6qEo/YsG0qWpmzYdg8Dxv8kPa+fN90g
gl7648l15zwvsAWgvVx64xbDD6hHHioMl7dlNxqwRlA6+k70XedpsVrORjxbuELY
`protect END_PROTECTED
