`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iKTU44IwrR6UEIcyJOnPHN05DZkjDlSpwztiw+5uyIfOJ3uB/WspslyvSVPaRr6P
0TzvEKyMVkdFErOt6SeCzl4H+1h4UPCYi4M1Ma7kFFbyJ4hnvBebSpTSS8nwzuaI
iydFPJWLmNvTRj5qtAW+L4E0qsddQkPTQvyt33OUEi/bY3j4ax6n2NmG46eEntpM
TthFW1eNpPWC3RgFPVDjC7r87SzlHcWGRXtguzY72ROPDRTPSkd9KhqNU1S0dwoy
uUcg3DUjB2etcHVo6zbpx1DDpkBbBMKZ5E75pS2Nt1qGZ1w4p8u9mHGJ1MRckJoa
XsUUsv4Ipc3mjMMjTRcfLvy52HaWZtNnVArSG9Pnj/c4wnkIj5ZceX0qjN1hASsj
2NUHUV+hZT/6H0buLbMIwrnEd+C94Iiw6OEIvcDfDifIk+ZAq22+MOtIbjIUCWC0
tnHcxbmydcniDu07Iiyp/CSn4rkle73sIxFUro8BMWzYI/iy2YMKtyI4jJT1IVAw
eTWvXdLBnKluIabGy4uQ061ASWG1ewbpoVWrZPGTGV4iV+E1GUVcMrembqgZcPsH
lIeorJDNzhM6CJ5PegkbJl5AOishcle2t84FYfMRnujHDEozgfHfcRpWvOwH1I9i
10sWg/lj0IMuDLHKRXrFE7Q2SzIGC0Pbc5IUjWbGUq9v4y9eDc1EQ/q1+RIfEVsM
hioJwRSSmthvq0AYs92zxvI7WZBzrHlTGzyIjhDxJls02Xp3HtcIUW2tnOrx8HJC
dwQIs7hEbE8xTJGIhVJc90WFID9iRxp/eDlW6BNql4xFTTokCRPkcQo1ye4EDTy4
sST755Wz6ecqeHlKHDeUNcRoKE6bF5GWtuJC22yRmbqUlcF2OKgNLLpSA9rZfluc
sACl1UMSz8l50cNtFSAqj0iSYfVA9Bxds+LawkE7AezX+21xnJkWnlOappminFnO
qvaEBGuEg3x+bvqyUxDiKvg+G9bhJr3Pe40Vn/6TaK4H52/0oEQXQcras2Q8vEAl
Q7iT1aV4AZSIZtU1+uNmR90hqfo0HV18FC+dhNzsiy/oLjVN32L3ZpyMc6hGgoxp
0aVUKau+wb6mPn6NMWoW6iAoN3Kl+IgupY7UuU8YBzRrE/jWPaKue1LGseB1YkRW
TU/+sFm2nAPJ1zIcXt1/ZZQYp56n+fWKACjmMbq5k0/1mPs2Bqiq90zQ9WqgU2j7
ptW7ISbbgY2sUgm48ydagAMDXJ1P0AHnCGZONGhxnFWFPNupx2RY3gSd9CL7w4t/
23NpcownghtPAIVVDqH/PL69yKzn3mdajlp1MLGuVtfLUzGXIf5M+KGAFm4TYfCi
aD5441Z7pMhukuxXAkGTK95QseOvDBm7zussAk8S7M1BfUGiQeCMHAGzoOyAXajh
POigmvg4/z5JUby+1/G5MROb2J/vOFAW3kdvolkqWkpRrCweW6IX7N75bSx/7XKw
CHb99BsFAfg6uAQJi1zG46nMnvQxX6JVTcpUMSVYbB3jpFHB3cHd5N3Y9ve9tBIU
Xmwzdjoz2oS2KWvaRW2zbyEW+MuFYVVTRgggpigAsRDz/HOdFWqqkqMz6Rze8O+8
l8rMaBbVxK7cOeCwYLBzQQew3k33YO0NnwkAdJpsapfJ6LnIQXp9/ydsDvCuzYRD
r09IOzn7OTPEGJurKnqmli8Sp6i0bbWauzfAJQRv7HFSEvtz9Irx6c61Zc+K8i9r
5U92YhXeG5WZ9N/qjTWAUgcfuLkYfPF9uFd2zlC/1JOJCjmN83jiZZjxmpvnaEDy
xPvu33wMpsnmkl/I7OhECkHH5Bweh7G/3+1IiY4hNq6crmmvjwl6+JxUmlu4XK/L
`protect END_PROTECTED
