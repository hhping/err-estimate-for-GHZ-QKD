`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MsL0N6uf/w6cHZhHRrXelofr7Gp/d6w+BNfioSZGa/EsIEoR0Q5cG5iXHoBTx2Tg
BE74YJbZhN0H70vqGEIG36YPLloqYHQ0oXG5rLSrL9ihu99MITwwAlFkE7z/fQHP
Z1K3b24fb/0s+XgTi1NrmJJu9c8NyapZ0qmxFv1lvkWq8vc9kQXKsN8Rf9RYqvgw
e/KfKQuIhrBCduWXkND24SfHBtjVGFAmT7zF0SGWNQ4ycvssohoKjt8EGafBKWl/
cvd8A9jJBlZc0vofFwC780gyiubLPwuLSgDCIzqrcTo5+uWr0fRdwN+EF7fAi/pE
AKTf0veNl/ziifnYXLyg21w90kvJ3DWVu04G+PUcGE8=
`protect END_PROTECTED
