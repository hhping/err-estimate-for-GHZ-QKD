`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5osPEWSKyuaxubpoIf+ii0hABJszeA6ENH+V8H5EDVD5AyiOzMC40QGwMX2m1mZV
Lwx06hStbaxg1OYqRuCPdVyvQD0e9RqDXvUs8v1fje+oReoiPfZBOxq43j6qEhE8
k6UEJIVHtf2PrkK6/9YSxySt88CfN7JAhnz9wnIIqVCMU0h96SKc9KLQS+Ic8Krv
rM8/WiCUChO3TJ/kQvJIQQim4+KxGfmlh7rsPo4MfDOXMJa1OfIIHMdu15cpq3+e
ubqwA+dnDxAFd98pS61KqUA4bQA+tSwQaDofqIZUkXQxA09UnwSosa02oEgxtAkU
7PsmLbH3kYQ29T8f+3HBDFdwBSEd2ygQbvbuS4an+N3J6eby1RogXV2+9v7ZibIw
XCdE6qh097qiPaaoSaUxYLoJniGbTEbiRF1mNzbsjYle+V+/ba4Pky/5gdDUFEiu
wCcWoAilhoc1k+v4/ID85nKp7wICab0pVrzTIjkDOcocSchDjL4oIaGZXTQ0yBSr
1OOcJkMvFBTeJ2Yr8G3x3osRTKZn908FLEb+TJsAIgoAk4hHIhEZZC77QahZv0sV
HBjUye8Vbb3dOcERx/0T1FJ0DpfsyLAFk0Ta6oHYUZ6fgSo0Udawmp10uN9yHM3S
Jvx0NZfpi20Jk1vLVOA4V6sM1YQFPqzXWGR+da7vtjSPGutodOvazh15E69vm8sY
LiMKb8XgzVaox2EK1RtxKGiZcZbHvc3A/iMuY6auf67PUtBUjDLxJqqEeVD00fQf
HpFwaOTg1/DKIc5S7TNfYIKDejlyWh2K6dlH35ZMWPq2vQJQoN4cfWl4DIO9MNeD
yTqMnPKDR54DQdtxtTIGKDLPCOqggbUunRpHrJk1GM1ZMyeZAu/UKbk1QTH8pPfV
Xw1w86HztY9V10SKAR21VZDZZtBVkH38LqEeQ2Sqxs9weIJxJ15wtH6wvccOxn5h
0sEx7H3DuyoLqirQ7mz+TDeLrIpAjE0xvUtkkQ8R4RlbIHBBdERQzEGgN/Il78Sh
aKtEfJn6bC1/wy5l3QwBTAViBrO9YM5sHYJClzfQOpgOGhq5ijsdNBtRr0cUmrtf
5dapSdNESBqh0yanehMmkEHJrTzxSzp8na/D9UtvZ86jLhu2P+HTQPIv4AnncobZ
CzXf6cQe7Qhga4zGEDIaoRIFzTzQsrsNS/oLK+x4JATVJIbN5vFQS6wwTa24XO74
OYWwwMaIStwHsXNbDYOcb/KI/83unJ6HI0RD5fnvKFJjDOGjN5gVjFnvLaA9gYIL
bbxh8Ul8JwkAZuvfMSIFw75TYdQ6sKN2lUPteMAKiUHwMpG9pQXtSPPWjRvqwsjv
swR2uJ+q3E0aeO8E06DVTl53Y1Y6H+IkEZ3Hijp685FXo9ZGgq2stpXUDCqLhKJt
zXH82glIJL/L9sfJem+CFwi3oCDb8Eq8ZVcBmXuolEKzBYtpp3BRnE9fPwDljCDE
SpbxR2HGRU+3ckmPE0iY9fvetpeMoGf1Hy2rRE8Y2coRE7aYdr1n/xVdbYYFRZSe
RsFsEYbgV3adKsiNT9gwRb+4GvVNKg1SL8eM8lkcwzwZSAVpLGVcGnJhSe0B4L09
AAfC3kTu5t8AvYyAb2/pAWOAJNkEpRQz8eCGqTQbDAZQfHJMLVyRt+J3d7Uc5FC7
OOKiUBJbpNEcpWt0mfwvt7EzbnSrYp+RSNg83Rg+OGtzxDDhvv3sioRMTozw86lQ
irDhpCF1CwrNXMbFOY8VOUeMfD9bi1TCibuxzE3XMZWlQ+0vp/hiz/1vBV1l6CWc
w0u1J9ABTwngOC+YlO5J7zKPfGicVfB2kZF1Zau89/LTAOcMSr0BDo1O8xhrHJXR
Sby/UWMbsMEEm9MMq/2u5scDK9OvTlGPoy99gMCX8FmdTYv1TQg+HMMXIB6JNsFA
pVFwumENmAWzhOnppabDCd60I/wa46iZPd+SWlUcdaZzU22iL+Fp7c2cNdm6rU6u
LxtijHlc7n92KR60Y+FUiLhlmXtTCCNhDyLX3HpHNjUdHMRYMxC5focq38KQwaKF
drpQDR8HN6ZPQo1lICtVKMvwPL/jhKwy05Rl9mzuvD5bWILFhku55MJVgbdIOznp
t3YgEZbIx+BuOc6iFZmlw65CxrXaizJWjvk696/3Gmng6IewvfRFcLVouPUQbQdV
0x8D59csPfnm5haE6TcCk/QzEiwWatsFF6whJ+bP5ZYDM39HTtS8E/ToHLULKdhd
zerL5RhU3o80PuQAxQb03o0S5TmrCwMpJfEPAIAWdgoSHFc02pOBz+0i+GsTl/Qg
ANCWcKDWpEoHBXAzBibmR3W2iMcmrQkFSXg53pkCUXRxolysw00A6ecvOcLNB5wB
4v9mgIJJ/6rXaakt6tzdTU3di+3YjMjb3TsSoo+kHNuGDhmEzbogoTrBaqUank+S
P0fGQzn/kmjxERS1a2C8K+glYAlqnFIyioYBedUjalx2+wPz+/J6tgkz6+zOO5er
KZwRQIYi7dSvTKKesDp6ZXTcvjN4m71+QfMUdFJ62+/S8HFyLF5D3adwQ+UXOTyY
Iuqo6I7EPygfEHySv29mdECGURdMb5qgb7FoLUlfpyMdNySe64fCs1HMtbgb5Qz/
rZEidDKxMOiSgVFQzHMr3pBbitp1wqgA8UpEr7UxYvbVQRFJLg2u/5AFxtbQLnJt
lW7heYtw+4Tuu1I7cBHaSAsRvbMnBm+aYCdOR70diAQ5zU+A312yUGHsPDCC4yPd
UIYwU5bQGN3o8EkahdBOoEABhMe/nisLI/ww0ETQYAErUZ7pTuETAI38OObiAOR/
SWC3dsCeVNyq1N02NkPk7iiTWlEzEJyeLk6lpAYkgtRbrMSd703QHh1pbFgOL+sb
/vT7UZ2i6ZI2sZqogL+z3/H9z7ZtWpOShxPYeIyC00OhFeyUES3QqtMh0xkhKKrV
QjDDBKeLZoO3WlRy3Gi9uSXqwe/xm8FhKzXD7Psi33cxlHeo2Q9G9KrXZY8ag9aY
Q63a6GqqD+Jy8QLKYW69G1J1+UInrpKqjwqC8P/XeMjYJLQ1C6oo+agCd9CnTcNz
NCs85NltlnmCduifxq1xuexgTECjr7WaePFaMcXhdCz3WxLe9kOydN9LNYsNlG3R
dAlar3/ieZHvNbK5lyzGy4aAspG8SruFVMCvtth0MXnHMzJbvcG1ICHpvmTe8qgV
btqEx4wO4/2I+Pcc6cL3peDTMsv5HLshkV7JsU039EHVW4trC2GvpuMusrMtebbd
Ygz0xl4prl0g8vpMvoKoPDVyytY/6fshLkjCMtTaqezDDX4POamIjWw8C8rlNNPY
9b4PGhCY/ocotmIB31vCZwOHVpWu27qpkFqd2C/1P24ImpWgo5uBIT+xoLU3Yt/j
TqF8jrQF4wC/bLQzFLSQ6PpljNnU4rjSr+fvVaoy3SF+gnM51lviRoxXsIS1Kbbg
NAVJ19gwmFFd4VWdUzEREZZ2JoAwiBty/inluw1HhijDqh2PZzkRzlKOeLosFUzA
H02QPz7S6etXuxkWy6TGzR5g7x4eQpvUIIXQBS9Atj7yQrwJBdAmhC3SrGsuuuPF
Frnhog56FkuNCCXVtpVmeKcZsv1dfyuPPQnhYlT5f36jBanu7zQQ26ri8grn544Q
Dnn8aNUHOg+caFb6sCYwwZmgbF2zUdt4/Xhkt9zYOu4SXZUZUBeleIvMaWUyDDPm
Ntx9lii3Ox0tz+AXcco3a/oIzGR1A9BvtkMG6PkrW5gu2vh9S61h2Ru1yg88iPjx
bDepdQBEFsD13b16LN1j3OyUsc9KnlxEEH59rEez16F3Ufdsc9B5p+2wZ/nDsHhv
DavdY0IpSzc9lz9WBFQOxlJkKBt/E1kBVCuvaHOFnC9Xy+/PbuBHjISjzAY+F5Qh
BTf3sTjEmIrvpIAIJ/oOmrXBcsvGy36N6v2OucxYBB4TDbjKPv/BFXFy8UrEOUkC
WYJtCvw5fOLUqFp9eoUB0moNgiGewYWzwnFiNnRIkUPU/fXJxvRA6d0IOB4qBdNN
Edc6RK1IHX9iKf6rTLdPCuEoWBnQVNzxpiPQtICaeOLDmz+Q9MzCidd3meNsvVb1
PZjRwpJKgkLtzv3Vruvsvf8lPwT+XIxC6TyXNqRKsI/7ryGwgi8Dxqwpi2h9beOG
6UKQRnHa1ZjFACNrqCh8unU7SIfjadBeLfNq0nciBa9w3/d+/f3ya5+yM+PitGLM
4nSdsoyaPGBbu+BNG1UfQE8gxO355i2Gsbptnwp+vRDSJHPH+YtjJ9AwkW+1/X1d
4K40bZsK2w7IGPW1dYL1vvAQwS8xEcXuifyBTKlMqT2UPx9JaIS4VACRxe/AqK0D
sVxOlPMgJEUZa3IBl0YhvTxflvGjE0VKZry48wsW9hltL1dG1nqudN0f7PJdqO53
Tv8F9ckKkjF5KkRJL8GmYc2kAnGVKWk/LtI2WzfYBXu3xXwurZBO5Ikenf1IFgXZ
Ps6KhabKgBD9NOJWdnBeJNvnvgWH9wVP6KBq6CKjb+1HPp9WKeyMSk9H1+Eqh+OQ
vOiTs8IxG8FxoW954Ak1mvknD9cm17D4cK2lD+majtLeYtEuC3RZYyi+LS7lyLkI
22/TATeAWfij+5wANm3BenMrMVSSTgbgE4YXqxt4u2aXktHVnMTzvDnV3DKmartT
NDNr1xQ7gjBISGw5+GdfohUBc/J6qyNI8ib98AReLan3Tes1bhcdicHuB2L1QFOI
eP22BtFh3H7ticVlt36yEP4NZInEN10jVjNzUo4LEUH6QbVGIKgqSrouv42A8BW8
Uv7jwLIDPbbUdMg2LqcwFsOvg4Bh1o1PetOC5c1cuCKKkEP4AC9lxEtczAtYVgse
5VikKCMKD/MfNdGDv+wElLOH6D6frI3ucBT1QsQAzJn/avMYH08bcccotJfEHPyI
fXkfM/lz9XDdbRHGFxy41PSDCRzHuUK75GFybhdfKQPtIjLug+jV++ZwBBaWdKfk
YQQVW9ubTNz5d2A9g/sIRFHXa66J6DEyLVgcmNXven3KUiWv89J+uXghVCDu3/wP
dr7H6ZDGWUfRdcRCwLj7xnOOVlKX9KMoCQ8Gjb8nUUqnPf0E+vZVmLu8J5x1DlqJ
jdA75tdx9Nbgaw5rp26IQPclsqId5kIJD3QUTIA+BaW2Y/bFkAXGc0yYzK/ZhYbu
n6WSOxHLvl6OrAfl27VbYXh+i8TPYPNo4PRo5WkpPTXh39tikleLAYFSihNQLNTh
7bHT6McjoZK3v2RPxiCx4QGTFyXqEfSGRQQ4cURp1GFiKyAYhiR7UNPSWTIT5sSO
cr7pYD+yW6UNnAYkjErPeNv+hZhgllPTXOXEjvX4G0EJOEqHhnWPR5+c3AeB/roR
+8kJFP3spHuyQa8kCqLct3WK8RemE+3UEhx3eYP7AMeKJPTtskmg95WD6S+O4nHS
w9/SXM5kPdvoBxkNau0P5RzsI/UArexw+3ISOnmD1vxWyGmyTMIFsAyRMiATnERS
S92z8F89YZIT1KhA63MPsqE8s6c0QR0h4rOQ2PDEU2AfxTrdtwlQMQ1gpzhQnHtn
DjSfNJG5CA2320iZQNny0FxsZkMG8R30nvYJWoPC+XjEL/sK9K/dwtFxAG6tdk/Y
HqJCEdCjzQxcgi1AeedybONu5NVlNEVDxT473eAPwbacakUg213HMFmakUneEGn+
WlGgj7Kq/QmHmqgca0L7UKPnSStLad006INZJEV5abo4zE8nsObN2KAsEMn8IZYH
LDU0ph0KD2qW+wEzeVRC9eqhHrbmLjOgkXXsFfDhMUYRPrVrmaG6fW28TRDtbbow
VkvRbsb9emdKy1EsUeTzr9yQtTCHGQv8jfIJt15QNfFRucC0hJzonPCb0j6r0qOb
m497GkhS0BsitY1Ej2bP+GTZ1TmFEwvPYUI3ZaaskBVLSye8vOxYYTl+hcyQzlym
5OdmAo8fPOOyIldViKUEGACWiaLbOSJo2w6Fu7dXUPnOYO7K4KG9ax0CLDY7fh0r
z0+Z0ZNMtUnefGaL/Qf1eyzRkhSlsXmq9cx54fdFwe+lfVzoFwz79R2PjN/MKfkQ
bnC6gZbGietNKReGWQWyH0dZdAIroO8wYLXCutHgi9UFu/PlV5NxnsXJIkWqqA3E
vD4I2yuAUIezujG19Fyurnz25oOM09gexX6lviwfva7kmGka0Uv1k8V65wvRjtqM
z1H2L3nPy03R3smso5wqy9ceOHFhvcAyytQhPGR3QS008KSmrvQO5utm8CycSldB
+p/yybOD+fmShxoq7iAKGzK/C8jokiZyz0E0U1zrMgJFe/oQgScHFS2IE1IRjgpE
6zV8U8qcHZoBJUmjOmE7hhdjYN5KvSMqV/lP4YqTpalCiyad9V0apndli9rWVxO1
9o9465SZHNfbUQM56YHwRIGzGo+K8shAAS61IvPHJTn0zNXruY+1e0fvcJDuoHjm
2WLacRSE/fEPZkIasxA6BxECSg2t4maanRttapsENQorCNgL4sBUIOfcPIV5JgLt
0mrgzvNpzd4qnAbB00cOLdygq10wQ68QbkAj0BvnB85SWLlAFZmCwhw6q6mhrgSU
kaUQq56s+x6c/gSUcg2bgAEWXtTR/zxqKwi/lo+yho8NwppebwBRtDnct4YyduBT
RfKxsqeZ+xB8JBYdwyuVIkFPng8POkBzqEDLW5mz4wkL4NUu1iDZSaNuNh37q5V6
wOXjSwotrqA83yDVh1zkFGz1FNorEWe/QgyP09CRmnn96V1OGtwDZE5b1ylwnmzu
wa6sx4gKAGetruEjZAOHqyI09l3k5EgSb9pTF+vhYIA9wDWgh8rDa5F+7ehzZ0D8
04t++H5SwZYVaTQUssyuBjnFHdrlr2RnJqMWeBROylHgaZRpmmZ+bZueYNDmkVDj
d2OVb9mPaWhWnmP68V6F6lWX2TrXqTOz0VAMyY+XY8EGpFkPXVAJOrZHIP0riP0/
dN/PYnL96/PLtBN2s5pqj3VemFrAG2BAFSBTXJxlT8uPpVmEkykdePnpQTAvdfAC
TjKGmvtZwvcG/JyY98mGnuLzzeHSZuyv1QDMmEb6tRkcne0S7r3hCJn2Dw73yG8R
zGOALv2bRnghQqG9iO9sSswtflqJSG491Q8r2R4UGVFG85iHNQrb4w8IXh/YtVxJ
Ez5qBVn65VSelMgSVgygAr2NAll/JXFlx8ml5vcZOaRGL/pIOYtAE0flft42M47F
/aWt047z/3UVrA+ht9uhYhnJJ5QYhT3rkDcnjEUXha0gY3Olngd1OMuffNIkJEU8
Q7479cIn+se4nB4YVEZjZTxKFkpXmRol6TQoeR/LSMW5lfD0uPqepyU3Rj2s4OXZ
OvcVeeYvsOyVbZIS0gM5KOoA9dS9+/aw+JfVMLzu2NBjjvuKcbsAOflCBwzEFCHz
ViuzaQ/vVNwDJyHT9h5OmYM/0hZXbFLzE8no4Llz8CZLDsf2W/NZgvhhFmRiJ6IB
8szr59RmDZWc1LHmJPveSl6r5xe3J8tu1n+4kAh4X3JDC5fbCHq+p5sKJBv00X9j
qO3oXB5f+/+bjHob11vNpJgr4LI4av0ddpUyaewWSYjC7Fpyj4WrksWKExaWFkEE
0JSoJ3jbln6yc1UyFwkcz0pN0O5hI/tSocLDrwAjoWLjo1Ou8WC6/2zOEtyuAL55
fv0Cm8jtoXwUZ9ywwK1k9n134Ui8T94A960E3mVlIzny8TzlfduEhLa+DfFI1oO3
g2oFbe9H5YCjGd4qalc7yjnN7OLUHtrhSBLDGUY3wwJQER3ZCj55w3pPsRJrjfdc
qyZQmwXnnliaDt+rqysJMc0jUNJ7gHbzg0WvqgjVnff8QeP2Ac79XVgwYazONTqy
makgvtfGH8QjhACU2VBw9tQLdUnWr2DFQbYzmGmiI4E2rHGUQOEz7iqvQ3dQzX+a
2zDgyvsAlsikDYtfGJOAskbCwh/KgeL7NUuo0lafi8c9n2FWk2AiKBEL53bzKTmK
xNg9uR4zdLqVfWsnec0JZN+9uuyxiNaGywfE7cf0DwyGMB4N88ZUcEVaieu1afMz
wnvY3Y8VsTVbb7nJJP9QEJUt7q/jzNaw33nwGs1NMITfPmm6bO6khGXYksEpKzKx
pcuXw2TTvuci+BawRDx4OQLN6eFnu+YBqM7Se3laFWNE+bW33d/zRBu7W5od0ESi
SPjfIqvh0Sdek4JaY89GDdvUj7yN4iSiFqFZEvCHqctrv850qsirNpKsrFw8NAX1
`protect END_PROTECTED
