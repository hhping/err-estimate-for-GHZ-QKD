`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dZxrR80NqIslA8MP4JPGlPkzzfavX+HymQuE3A94xvuU0NDdS8m789bw2+PXdcbB
pY0tda/InvkZqhs6UbG8QsVGcIQP6DhXox7fKBJqAj4Uj5M8HZnIslWfs7nRbWpF
k/T2I/9LXYkxHGmJdJp/wNYaoje1UBtBbq2sxGo2Qw3VlnogjnrPepG6sVpR6sV6
XPhAAikc3+qf4J4lwIhqamnjvtVksdzR6D9zNzSgQXW+78ykDTVr2SBt2bFJvkkf
DXzE6VYd18bycumLO6peRN9h7rJ2wwtLr7e3/9cVmsEPBkTvm8a7QX1ohIezuyFo
0ARwRHC4vPkPpQ8b624yul4VaBguymo38kHIQtbBR26G1eVz9FEosogt93MuWLO0
amDz955PZY4emHCqUPCaz6wWJvebPoIjchP0DBD7NnjQUKkdD+u1HcnVcQGeGm3y
h95TxEAMdIlg7OfW0AdZqHa3yUsgMBRyZDSZ1UFvv/QxNrPi9M4WbfV0AkMSFDbS
pBDr39dUpQ2vVa4ssVnWYuZRR4CkHYe8H67e9ATPdzn9ei8Bt2ppqV8zC7mMmv3o
Bpb9edC0r7xOqTYaD4MjvKYP88DrUlyMvr1sTAmhvJcs3fcSrYH9x8WEgfBFgnkl
kpKwu5/RJ5Yttl/QN11OuXpXs3IAJask1X9waO/ZnOqiwO4S+ABeyAPI0k7kP/Jp
OBTdXQarvGFvW81Ce6FZfgcxgL1AZwXqHWguM0qZI/fXQeGOdpwAz973MJE+Eumw
tFkMq6c/arCTL30xahiffktHSXwcEUTbssTk41s9x1f7VB90+3TvBoywS74Mu7Jf
tpawJiS6HFz8XAZclFqxGwhkcKZ02DydNaTaWydyUMElJVbv6C0ffzkkDskJp/CT
YLBmg0uKovJm2y07zS5lgpRu4USX6So+z/p/ZccMgP/yLWRdB/w5fxZTtnrdYyQK
QqvoxKBwyLumPgn4AXBke+7ZkwQYsjIJEE5RZW6RLbVWbx2NhuNf5OfLvdxcUf2a
3FfhvN7b3dR0jT02tJoNaZOAVAfIXgG9zIS1Z7SKbNG3vgCSp3kSkq3aKONjr+hN
R4ywj0j/1na8Cdb+BXYvhCndg18GEpqkGcbUewQzB74LeTatbJeOENGW50tVPr35
bple9NS8653DIgoLsJrtLh1kyvMR/u/t5nOJzlpv4hyDDPFv14knDr6k4fNDY7+G
9DPNHd0mTprs07mwYGWE8XhE3L+//aaoPSdCvIC75SRUZuierjmSOkVmjBBwBP9T
`protect END_PROTECTED
