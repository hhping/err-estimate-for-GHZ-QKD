`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a/9Kx0wv4sWoYIBGWFUBufHNd+kHDugUfHoGXoEONSrgOR4FhMLb3EWfpr2xlFNC
7PA8SNB/wi8x53q1Mftl+X1nnt3lAn3HDpwQBmOk+Stedx6U7iyHOQoQhXwIcqAh
bC9r+wQ3oqL71sF242u4C0v+YRkHYx5qUjGaZ/CkSZKYGeyAz93T/JKBpXYEbbh2
ZHH2PlVjpY0fJGtZsw322FsDTP2nYinIO0zFQSa1OGfhSaNsRdPrv76GObt45k4Y
fUq5sr4J335P60Gtg/o9NxGY9WL5UOZH8A0qCYJX0Yp0G2SNliHbvefmkXuBfXLr
mKAqYXuFYhQX3IIBeZk2L5yD56JTBRsZj6/gJJxWKEOfaL1bpMMYTOQtdjeCPPK7
YAsp6cWiD4SDU0FzR86PrRGSFWxKSTCplo8Ll/05q7psy6WtzUIp3/9CmjxvBrQv
piRfUsENTkeoJ+wwkEe+O+xY4G2H4LoJsf+/Ykqt5BON/bcRxN5VxvXce7Zdj1Hj
C64vlS3RW9JXOhAFL7Oovr6Tdc+naexJurk2Z+3BRRbxrjG0JrBXH65iP9skVCMX
XJZqlbSZ2kqGGmSZk9gJSA==
`protect END_PROTECTED
