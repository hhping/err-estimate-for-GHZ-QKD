`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twUJTv5piDEY1LWHS5NsbBsdwN2zzd3BYuMVwFJUTU13zFg2U/yrTYG3Qqz9TodA
IEOtJRGu6eDQmaDaXtUSwGwOKqgXdR97LC1plPF+7LmHZjoWqNkhTGFv7P25GM26
kZ9KtK6O5JNw4lZw54XJr/fBW/RTuzk6eXltXh7dqusTHEM3d02HPa9zMI2QP/3i
5EZ14KA10WV2ybF9Dsgb1j05ZIojaDsPKJR9lJObIJpNj2UoMWKqCHVXUsaP3QWU
DN1T1JIU9PjHjMv2XW57U3WOzJK6BkduSkRqSOqLtoIcht/OO3QwRhEgY+YbuEUa
qgKi6odxV0fIHmoMrhEo+HHSlt64mN25W3gsIe5XlZ/7cNxZhKmJsUdZLalMl6VB
V2PTNXE1Yvke5Qza5wOWduh/MQqBrwBYr4QQvVFFa7bkgB064wGPHZquMNHbCLJG
Pj6qeFklUbjB0yhRxDy9yUY7LsAN720lP5gNZ0ORwDXca6K55ByuXLiTpNi3NOI9
K9tFvmlvc50KENFoQOY1Nll9/ov0791uVJsj1hsoNZViHOs7Xykvl4XiEP3268Qs
fqNmVyPXIeubD3x9ZzrwA7uW+gb5Y0Fypdafj6ySAwH1yHm2bBC4h27DUULahaba
pQPS519nrn9jl2NceFQwoST/ixHnEvlqIVuYxOVHypQN/w4jIlbcrfD6lhjCvrQi
ZPO9I4jHblCe/59vKrk0sM9fMkkYbK+Zwi8xc3v1RgxAD3F6wZNZnv1vIj9oyrgs
U1b/8K5hhddOHSM6cES+x6dILOUSQuZ2ZYjh6feXPZk=
`protect END_PROTECTED
