`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6MUckTAP9TOUEB+Y3DiIsxwyv67uuAuW/eTfvQQ1X/YSHBL9X2umXP8HyaO9xkE
6QKF/N7nu4+PQHHLQ/q3UhML92t9P/QoUi7LH5RwszmqGrSssDl0DQHIbEmk7I/X
N2XYGrRsQnLqX5qjtLWwkNO8JoC/Agl1K4D3GRpvW7kdjkiVYh2zcAeqxhTj6meq
i4XvIUkG72V3ZzjYV6UAqFmHcSxy4W9HtIrH/oupHJDJkwLulPR4ecVoazO7Kew6
knsK/fnTVx8BCEKi2nlRtDnrfzxsWHFwyjbx+haW86eZB3atcDyL5TkrFP+9TUsQ
dKQmvNKTtPNTDsMfKvtJFYr+ACyG8zCEIlDdbQSxOiyDTr6AGMXtIWduDs0fLkrB
hjbQv/NBejZBxBHMJfJTx2dgr2beG/Luab32XU4EiAUPsms3dFgw73LPsIwNbZuS
VTyVMAk2FCGo5a3M2w34deh7BmqqjQomEL0+LOyiRo2pObuAJVuUV1v0YCyS0fct
uA0A1EUGdlcwEBcmS+UUiecinP4pYZNr2xyi9MPcXGTgMWRUoPoHuK2OtcWgoGa4
ABe1+8p4OnkmkMWMBxYTPbAf2uVS4e6kcn5pbPUN5Z1SfDay05v4N7e2gYAMi+/f
tABgpNJFJQw2Vz74K+q+KrtykXm9dD6dSd9wForjktDk8dKGVu2Cp/jWUq5riJ0m
VKqzQFW50g7I9bQ7dFt2wjGv5RuhHf9m0mBM2MJ2fGWFP7DYApT4dRpwt0O/GS+c
cysYs4UuZfWH/75SPC6xDUAxXV24AcuU94DH+q2TnxsaytKIIiJ4Wg9D7gONuNDA
Fw7zS91T4mxRrHL+Bauetg3LWwUIIi2Ie7tNBjnfv9JsdY9sNPSD0atoIZGF9zzb
5BVZdhi42gC7rK0mEGKDhu5jLxjO9Yy/TgM8cKooc9CISjwSH47OvMUOKQ2doobE
oT5k1DtB8VvHVKdYcZ4a7BpmHl7smH0ElbMAiCCtoZggg7s+rW0qsRTnJPAKikZz
2XqbZC8tzkHZtPnNBLAIrPE5l/j0gWWDZMydyQW0QCBpGj/lklg7tWY9/9rWp41y
kSDNtFMJIiencnbgSAVoXlonM5MSeSLxoBWoHYmN7XncaGKt8ItmRQdAqL7KdQJS
5xNQJhDVmA6HXH0ucofaqsivAo2MhI+uxufFY9DKL/TaV6cT0USec81HZml9cV7C
kvgRovBdeC63IuN0tFsIDHp+9Y+ZYoHiBXrMWjaqbdBhX2iUvyldNcPE6vZ+Y3eF
s58fQ38da7d8MqOptH2bAUs1peAzQ4rfr8Aha96+kU69JtNBtOEZdepN+yvgkSgY
ZwQZfA9O2kbdsfkZDvkpNfLENJjo7ni6oSWL9iVwPHEt6ZkH8DPNz5NDl4G9RhSh
mNJiBrYIReJr+Rhvbm6QcN+Oe83hAK02b103LKJIIKEytcNoOtFMiOT7l/8SklgV
WnR44QgqIbCL4KOF9DsFC9u2ik2W69KzWW/XuJPNuJGr3ZSMBOLbR8OvavWHKWc4
aBdvSyrrPZAZkVfqfM1N4GYfehx1fyBZaJ87Zw4q97X2Nt4a/l9poMAE3MsN3AP+
tZhNdEpvsOp1TuCZ7shOFFlwFONDCqKc6IVdXa8AHfg7uILFurhkHuroKh+Dt+xn
yqyOp+jsyAtm5VqUa4oPDTCmDZ+hLphWVM3a0/TeIzUXztTnWL+ablWPZl0TzMXc
0kXPbGN1wuYoBeclpyQqeZR3wSxPM+dwK6uaF8wDp/u46UcLERUIayD5QyuBMT7H
leVC5iiE7F4Og3PnRyIc4pINFio+6JqXAnoeQswimEvOiHuN2rKEGL9+CzndXUnB
C1EgsBkcDAo3w4QGdbLeOqv2sjS9Z4817IkQ1mLewPesQrtP6Yo5zRZK5QmSMY/r
w5jnVRwGR9YoMj09UVvEXCjVRwwh9y/ML6jz0RYON2LTfIborCn7V9mx0ae2MWKr
MtuUHurJhhOM6NcHdpjXq2PSJeGlugP1/gcUkzgj+leXPPse22MEF0UlcK1L8MIW
8U24C4/9p5c4l9ADT5EAiKbb5BAL3IULCliMTCoXXVp/CeJ2/3AfYbjtX++tiQys
jkJlTKuFWPRNLHq7P+SL61hHxDkKYo3jtBN0yNy9Q1DSUI2DsGQj/zZZVtvfEMia
TvOmK5DSvX9RmpCgbHDZG2rL1Upo6k8f5uge7bDqg4519sW5I1z5UEi1pfaSww6T
Ithw+qA9c71sEK6sYHgfc8qIESWykNGH8O9wBD/eEsfcOIaefgBoZTGbf/RJgV2m
tFg6zAPqC1lL03e8OKJBQH27kJR3rZQQUvWNQj6pZmW+WiGIlo/aTKIeRZchdIbV
INScC/iHvrqgD6Ioe+GqHCB1U7B7E/ASmFw0/P7Yap7VzW48n+Tmj69DAkX1ZOuh
8MyMYEvXOeb4YgSwffBKykDkYlsLG2Tl1Gv8WT+lv3/TqiOdQ+8esC+b/t45Lvcz
WCHDxDxLvbZc+cn0mlrP6eJyS9DTpoFFUYGJycW+vjhmZ5Lk041M0P41cCxLBMB8
iNN9pZptwscAxuTqzIh2Ix6kzOC9wLejzgRVP7YwWgTX4xqUmrSrgqQakqaQLmR1
/qJvcrNaTW3ky4cWxLrJrusNfqYIKix+NsHFVXc58jRr4In3uFJDqG4vnLq8o6KC
LBz2o5JcQU+DzNN42SnfV3CRWzYUxM/HbWsEsrdY3g7i3guZgPF/717XBElXOKub
DYxisPWuUFsjfYprUSnrhULVu/H2PfkjIBim4dgNsUjYLTDyS+ibswvVmfeZYA5A
PMfptr1vVAph3a+dzyq5uROijIiEbRb42RnnjB3mLPJki9s54eA4FntkRIlz9pex
FLGs+fkM1iS6gLwWi/XiIEwQadrtNxxgomIXq6zUW7whG3auZnAfLqqzgh0vbMDh
mOnwrmJUblAYtsb7qsDwUSflcd4VCIkH1seL13eY4va9waeAF0whRNizR4BGaUPR
FRgUUq6YvA/gSqxuWbMJOALW/8TokRaxHQgzXigmDvyp5zqMlDm7vBT23eaOzvZ3
H94+IV06S6+PcU1WwwKT5pVBqy4XTGyaLb9NMlmFnWaNipNh0S6q3kDCsqis3B5E
VP4PGm4ZZRaZqYNOx/gY4AQRhOuc2yzecKcJb1SOgER8TjmfjzYAuRvJW5Iir7kD
8zpUNN75r+MCapHMoXOcAnGZcFH0adjckhuhxnaJju8u4Z/x2ELHZGHEIUetWxV/
vxYzqPRMQWY5sDZdDIOXyWOrJGsAIEOLgCc2wanxRDuXUrkkh+X6pTPyEcmVMjlk
5rC9c8uajkDgJpKM5S+hpPA4I2NCnehNZTKse9IPwUPqWbh329HzGBOdovX2WRC5
8E/+mHmT+e34rPJxh+X3uZHJt3mfKdIZ30oEijdvVE0NDtgko4VQ0t91WwQneRQU
3oVvuqQW4jiwz5x5Azq4iinjrWMwqJUg3PKy9wQpgM+suDLcXe1JGn1301+zvX6k
g4z9seWo9dv069DGJNlGpNT2qdCUJZnf6fLAyP9GDOKKW26BxZDA0ObeOuvbCu4B
YsfNS8I0ZNGHZTijtdIw65tinNGWtRvRvGBXJMW3X+1tsJvfXdCZw1llF00He5z7
V+OnXGQCMuyGauwLkw1WRaOO2FCc3r6LqpLKU4yyKMQ+dDYQU44sPIdEZjmCev9l
itIOvijX8IB3u13PKIVyyDRl4/+5i/pJgIaHLbvwT3nVk5OQK0DcHxgc/HXY1Na0
O2FOdH9u6h3XLbdQ5M85hr4hJVfCWtCcFc9pQ8xWiWRzzhYcby0tvmposY+T0KKY
WuP052gx9RQKs8VvWTYosSzbbEv3DiB3nSQx830ZX3Ni13sWQiXX56A107FcO+xp
wXqLA7l+RbXrd286nkaaKbZBGi7361vD0VGY/Fe54CK3GKWg4GPeNBhOMqOxM3fN
FOTgbcsOftkDNgEvQ51WBlWIS5YFJw2KTJyfkfkiZ/C3VKEiQ/XlQrorsrre3XQG
tZSBn9u3wZdQRqsmmrqeNDO6WCKGUXX+7YB7MeL/+Z2iVr7mJMllDQGSDAZWhNnQ
669dSBcAkqgJotH/6In6cULEK5+/RovFPLOJ6phpDAJZLbxvTHBxLIsu9RByjeto
M9KizO1fc9s/KrCOqhf7wVckzWlZwxse2MI/3jWu6susnJQJ8Nd6S0VfePHgHpMB
aIW0L8eDT1BZhLTV4RBm76zSVXW9H7o4b1BIE7PyBrgXLwswOjpc4j4YzSfJMYg/
kMH8GGGKSiTHQ4rY9D2r+Ju3m2dtmzDW3lR982q88r/gdc1bcJjK0IqG3zR6AzxN
d7XAxxzbK1SS/K2DIpwSIm0WSYTVsf1xAJkEgwr5CThspCE0vTrMDrlJ9tq+kY1l
01p9mYFO/T+n7IXVdZ05QqoIRtAC5rQm/zB/EKbTk4yYR0xPkTiUnsjbhsPkLMSh
bLbFgqkIURuYB3BQ3pf5UHhdptPyIkXDpLMyU53eHKzfOdNOotxQlP2S2I2k+yyy
urmHPzJAdQs0fvRpLda+U0hIDjkG3bveIiO15jLGgB+g/l4OST4S0IN23IF49O7U
evyEIKFRoy4utol97CtlS7CPcjl70/+zw/ZomEMDvJpAoCi39KYFO89+Q18n4/Fx
RsXuN83bBbEqEBXYriP28MlU242f+dlnkXKx6p9+HEDL3jO8uKCO1urrpKHd7icu
ygV7KdFPy1cuYBJ47LaO8wJ3C/L5hqR6QZ2WkOCc8P0IJtd28sUhto9WeY+6cnEA
8AIv4EH0HXe4UdLOK8D/3+ciuxA2xKCoCgL8wPi7V5ihLyRbjA6r6Ifl0wAH1Jng
ty++5blbUPssHa61DaWVU+Gx1ylfb/ZRL+1VzdglALCN69fnVqS0ANa346BvlsNc
E4Q6xh1tYYART6hy6Z7IxX8XNlq07fcOsde+6+vaGJnyR4aLtlN7RtSAbN6pYgFt
QmfnrTA6zhal5l5zTXAmms6clmqk4BB/PO1r6Y8vCMm2b39So7pP0fGfTXUtZVaV
HrfF7yS9WatwuEFeF6FUVz/TS8G9c3Yoi/T7+5bDw/ADwOY9brNi7yQJk4r6/7A9
nnUag4W0virxwtbfaj0XY/A9zdSboeQzPdg8xXgL2CDgYAnwIpTs8m3eGeTZccd0
naPA5cjVMLLmMIHLuuzxvkM/JZuJUn6Zoln5qc2ZYcqKu4I8ifphWtBkLs8g4anW
vDia/bhbuKdedX9NT6VyoK/bqRlCHeBt2+9c83/8y/q6lxzoH3OyajArE760WUiH
eke40nxJyjP6qc7a2chei8vCMLFzPHmkeX5J7+07oTfunsOBOjvgUqLIMCIjfiR4
5b/RdPd6SQYNJJpzASRGX6yO0CflmqvaaUeUNVP7DAHRvx8lG24i1Yr/sd+DZp8/
Z1zQ/nauNwmJcJzwgLHLyHVx/eABXkIKMUr2GGy9wsmM4+LV71mGpOxT/KEcu/cz
QfnEpxir+ZHc0X9jUXb3Si+mL9Mpqn73ERsaKU/AVCEyR6b9Im6D1QGh252GyiHx
NRD7hJi1qq4UW0tAWO8ZeggHeT1uWbfoveRJ+e711hs1+o/o6cXEf3S8pd3+6Pyp
5QA0ACmquCkIJ7AmCnG6pQxRi2MC/8JhZG0rhkMQIm8aLSg69yaZPQtq6oLAakOS
rOcGEtx/m+zb1E2K9XGb+jVFH7bZwddEAf52KXZ3Vm4eFICUIaolGQsKBz8FQTmR
vAoY0jtdutatpJYeMWjn2Ti7oeQktBDL6lEEMzNVKJGm9/fnjAk2yUssr312bV77
gWtBhyi5bKBrButmTgr6883k1tylbogTi84aMvUmK5fKdBKCJPzUmRnakn+CDf8r
VV7k/yn5R6L/pq2Ey8fMWrsjxzLKIebwds4Hfb9V0dA=
`protect END_PROTECTED
