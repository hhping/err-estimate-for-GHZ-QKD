`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+EobQ9oLutHwzUF6lDmvKw7dX9hk+ZUiEgsm0RrJ+DlXF+7yXQM/7HpQDogp1G/
rLILnJ1iUlDl24WXL/zIvikQdMAVJO1eLsZycCP9swJabnmj7ivH1ni4JvphfjL4
c420RdfbSXA56mwIDC4umnwwWwmWWgqI30Nud9orPh/LQ+Gq/TrKKh5Vs/llIfHE
xmvgM5v50ChCfuhEYCogjojciMVvIM1iGv4+WgIW6/rHnQJk/83bn62SjdzvHtIE
wm37o3i+yRVm40CsUR1MXxA08B+op1pu5/zCwKMsLp7cTXNpQg3c6g1mLpJmsmnt
u+0Dtv62J4baFoougEGLVac3RDGj6GEPRxhCwb8GEg3SD1cX/Z75Ie1X/6J7W0CX
xjh/23C7WZZq3WtELcJeWeU5mBkmF9ByJARUk4XpCIQGcTF5oiNWsQ1IUJqG0ZPT
+8Q/8nZ4R2gMYxgt9r8NRBFhNKQN4fPKnfkIvSaCfWzHsVTMQDQ/baAQKKCM5T7l
yK59juUF1RJpKKx7J5sxECJybp4Yx34jX32ciq0kCDEF3QWg2vyapD3e3AIGep7G
u9JESUSiYjLoJJQ18n2jL7VBDzXn0H7S/yuwbp9L/KQ=
`protect END_PROTECTED
