`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0rLgOC/QYyvo5ZJlFh8hxDwWCLlGmjHbi+ne925TXy8pOqL8poD0ZWadLAaM/lz
Tvmaq9NrB7HfxbXKgeoF3kScoXJ//EWcK6Rq2/Q9vw7TQKzP2vxY/VlhZkqEMp/s
ekffC/2hJar99vkWI58ZRDInJ2YpVyplj+q4HsaEdRCm3hi9TDmLoO1UgmgVkxzp
l9M7d5522Y92RdKvqmPZszQdDfPkqmEZ+V1bc0aZcWoW4MFmONcAYQ4UJXaO2RpU
7LLgcSgtF1LL5gZnZyfEssSFj2BqTimS2Ww6tuG5X/UoR3DFabrUt1ySWkvxkxBs
v5X7VRlGkgxvH8CdX8xwnOycc/YjFGjAxTZxbQ6FZU2I94tGIMDkzY+LxVrBImYZ
M1D3qTS1snRUD/0oB7btIAD7lWFcdvB6HpQNgbyfHHdDVyR5346rZJKqgu20FGWK
i/kDs2BEhAtovVYZ0OZSggGfOt9q17OdZpjkTCsDx9XRePlwoJYBCHOiple6nDSb
dCgCqgE0gcDow8AI/LYbEmU67nSGYE5cG3+mO2H/pFfEMhdKfIrvEfQl0rZR4hHc
Na+5l1nQmQiA02BBnm63mKR21YuDG3orUyFGusNfiWgjxBwLo98NchdmE0dS8GQx
p0xm1sYSLcv9RwrJ7Ga4W/nV8xl1Y+Jy5pWPukHIrVNa3LP0zQcdec6Tp7G53mg1
aNEwu1oq45Phz+KaU6upGWD7su4ZOipgtu3CTNn3vVU3ZxO5MdTW2GpXZ23FFVYb
Gulhnn1W67a8+DyOpGa2DoTQKewS5cZPhY3PC4mK0Rz12+gDUFncMjKs0GpF6HnO
ej8nowLD7uVfRmbsfYNI3lBdEMe4Wbv71iOKfW4WEOk/AHUOe6Db4t9erHAiJPId
QRqEaWqt3froJ1vdxRMHVRA1RANIZy5WTLcBjnc7bvx1WVc3NfYIVSeDzhLn2YuD
BofRGlMwEFZWXrBTPjzjJFkskD1tPcjqVk+HTic7MxUJyjkpjbFRKiGP10U7uvFc
qgX82F4Jm9DYV1QB2b6r0K74d1k0ywPYCIHh/S1/Ner5hZNa5LsGHAk18B68P1oE
PoNy3KtblrhUgP2VrfGqFoNIynWuHE/WpogCAvTechIuHVOWoNf1RixshijmiSw5
JKrdm2wFAy1eusZ+7VmtaMy2Be7UGzeZAxM94EcwhijzrbE1ZH0akYVcgdbSeGY2
jIaJVgk42lLgKHo8/VXqwYoeD40MYMgLMzkKELe5gQM16IoZHybYLnhfDKqmKuWO
Xww9/dWtUR2EDMZnCElnfR76k4NmtUjy84MW1ry3Z3PJCJPUKcAdX4WTCKrEEpky
RYfJdtjTx2xETckf+z3uB34iMOIyr6PX666N1Oi04cZZ6UAWLa9IugqgOq0a2keE
YmtiEm+emHU0jSCxFqJ1bDsVnxmvbGYFE85t4/o/JHkQAT4Ngvw6Q222xkAVA4l7
C9HhPmKJ0x39xj55nsG28wJZg7cK4+rXNO1M2ehDbqUKePnQYZeOEDzsuXNMGDMm
EOMQGW36BxtzMXgEFONvP/Jd7iS7+fjcSDOYjJBDkZtp2Fud1655UrkUXgPORT+e
W448QygwQMt2VMgfMCfOlsa/6BUH6F4C2S1lRks0xAHcyUofaSRewOgZFtVp49E/
4ik1JnQUn8foBB2IKnNzr/eZPHHD5j6Y7e9O/7Ze9PoAQGdzLT0kiLhmhynEg3FA
KNOBrjYpi/Uno5yXRpT1b20s7lOMwve2Vh1HgtMGDBfWrggSiUmewKBRdaRRumSz
WSmEkprASexJ7oXn0U3l3akdeDeJekRD/AKTYJ1FMEQzQn05iEkF4W1urH3a465W
LztTMXamxjrNlIq+QaDPt5s4Pg2SjRp4y4CjJymHjx7ehdHBSzHn4SFm3D3wtvZ2
fx/kCmWbZ+O1qa0J2AmhAuOnjNmclklKW4MpQeLTGSX1UTcJF2Mw0hX7icTq2Z0x
Aje8NJbOGrYiyu9RJWfXnRHNrCm/JZk3tT/Cz4xPQgPAzrY5IdGb1B6bH/rJSAJq
n0WdFwLJPfgRrfkP4C+Y+QHaMU3fBgMl2Dq4GzGSgmZM0lx0oh9ZpYe3TQ2IiLXE
`protect END_PROTECTED
