`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2wBawz6ihSmWWwSWlqPAp2SimjddQAFns5OLZftPIW0K6g/aKg2AUvesQ/uv1w/
pUU4cEdpIfXjUN58pHJkpdUgUUonVbsq6dMaGXEU8hJbOqD5qqEEK+x6fQ+ytyN1
zDZZYfXDHVmWzGwYiStTmuPusi9CAl8g6J5764e30v5rODcakSd9RbArYjUeUeGU
U0yagL4RMRK75FbIh+d/9+kDDztbJTOFrP+6ZXLktlRCugpgA70UqkhkeqixSKhp
5+FQa56Jsct/VFl5PlXdeoGPhLW5QVMuYkZRECeztFq+kTSIWjXBdvokStyMAil4
8rU/87Nhz8IBG1/JBIKdvw8Ew+ewOx+0D8lKEXT4/+YiG6p/wBXGeGku1PCQEjfQ
J9e7PGtI/GEyxRjNRZnIetYdRy2/2ZtXa1zXLGupH50aFx9llv+Pr4GxfISARxTZ
IFtSK2vhu99Puy02vJgrCOcIEp7S2XjZEumcoWTkins9YhG61/coaXB3aLUqRphJ
6Klde3PWFdu+mxRDN8T2iK6uQlfNx6ZMJ/mUGvn4Tc08VvWTKPumELduFkT4bM2C
B/vUIr/RdXaDK4aOXk/y7MbCkd9KidKdLDmz9uDnSLY5tLJrNLuF9x275UcOgRiC
/4hFyMxHA/Dh5q2X3iCOYricAFBC3PSCo+N224VKYxEJoHcjIWAl4NhbpfDFhhBV
AfbtzFLhpk++pFAlKQLim7SVL1q7HcqWce1aRDjQSielxupRGmjPahc63hfACPbu
4o6gsF1GVE8rgbEhJV8OefKS/pYcWQunlcJx6h48CDAdih8gX9x94PY8GhBHQnSt
J1gq5mq0VeuHtEZ55yHf+QetBWfoWAqPSKhlJcABjrnv84KDtksOlkK2gF7y7KXu
EhAJR4gQrklbkI2q40B9VUXMZ/Cm6J8G5Mbn7TqScdPu23Z+N7XcEpi6WFlW3UH8
xfiF+0o1o+RydHA4xxB/lnu6a2X19b+Q5PT+yxqFmaVE8VHAT7KqcqYVxEYKJvjC
+CTEReAop/9DfgWYX4yUJHquku7LK9/zNvxSZXYyGlmStTxEBXrLRsCwEOjdi7EW
kUlfDmkKBZRt9rT3bylKipT43h2UBqFSlYhEkCNgf0CKFjhibc7WkCIV/mnHUudm
95zZuDKTt+lCfeAQlJEsX0Qnw0OSWlEJM6Z1Nmansng3zfyImaAUqD8A2ePdRpCi
0OcyRYG9PhzeGcmLcl8tZAKhUY2n9m5oRKgQEMIY7Bk1LnootNg2TnXViszAHb3+
h00gxIfU6rFBSwRK3dFQeEPW/qmbv5QIAdcbiLMrG2JnR9jwWWLFCXn8ZhYRLiTS
deQbWoYrYkNM/v/7u2f8bq4TaQa/4Z1kCPizrXDybfFoB6B6L/MZqvs7T86YNiBz
3DdcKQznrpMBopvQ10KOpwip8NCLQo7cM9b4Nh7E5AFqfHXvsSnA6XX6d4nDQgHe
/c4pnoijiMpfbIUApQNLj2njJvfB5wRlpSMaXd5wqWp9+PzpRRNF6K5B5SG3FcJl
6YOdQEpN3kZOXb1k2RWHE/sz9h6tjZkioAi0boGJcADOxGkNN3//0YP/zxxk9tGy
Ud9uL3uxPYyaiM4IBL/2Mt3aRSKQh8boeYfeZO1mz2A7MCTVrKlv+jtkwILgt7ZL
Fk98JH6thlad2Oy0YgVQa7UzKKUcoASxMrVvEF1wxOameMpLE3R+HhRIaEGnZzh5
eIgzLw3Zvs382TTzDNPu+Pnyg2tmrFaRFyMzA/XAWQz5QcACPu4fCUyKwdzKsFBO
YFE/QvDghiwE0ab0p1tYG/Jphii4nP0S58nSdPoV4Hx0Kl99Vxz2gPghUYl8+6e3
A5mkpBnYEvuwk2RWVND76cO6OVrt2ZfHC5NPSvJuveoiboDALHaxwO7D57Ke/1nc
GtQnDvugtLkzjcM81Ii2lA==
`protect END_PROTECTED
