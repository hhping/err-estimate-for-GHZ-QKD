`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PZiJRjrn/I4voeHxzL4O5u3MhJVhOxJ4Ed8BB3mjtw+FYVC3MmS6Nv1XF618O4y
/Yw5AtXdlHE3Zs+BN2dWxDAScU+BPfI8oXb53kiKOZBzo6ueDVefYz4j3Dup00Ob
M3f4i9XatFDFzLiSpp9u+DgmybxRnWZyQ9qycLyIVGplDcf9joKXZhDFLpHdNoBt
5g4qnTduPxOURjOQPD5RpeQ09i3UxfEUTts0v6dC30eOE4sdeFwwZTNZP9ZKFMaU
kqI/S5vuazXtSsswNxm753vl4MT+r08HFw0ZCwUdUwuVKU4i72uLZ1lrEfl7gDgS
nsh/clofXaWKbPov1yaCkaMCDhcH/MIl6ev5m+x5qEQAcGRH95Wm5ybvvC37lwu7
dSG1A3LWyomgSilbLx8AZWb5Nuc04cLARkcKk1PRqf+mOt7EX7dxH1lxrno2RRBW
fsVvleZ3usDQfcWo53LI8CbiLZG0cVbhUMbO+lHu3z935lxxZc7SBwlGGO7cJye3
`protect END_PROTECTED
