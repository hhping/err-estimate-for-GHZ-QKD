`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Gy5iM1zvzaCriWO82CkZtioPzXbuG9yrKzrAyCNXnXtbjK+NT2EETXnw8B+Qqjs
3rnTGI7C5qX0buCECR+CFw8az9FV7sZPmEKSTO9VlcHBhv2DtJ1fxwxMSLN3C23k
PWbMqeX1HJBW7ofR5FTwKuA76aojVq05xOkf4h0jnbhwNUwJ3hsJkyBvJGpmYVsV
cykkFxBCwbLnkcqWqoO9HLV8bq3pOI4wbbi47sc3gNBXJLFeRmMJ59oM8rxmnfvT
NaiSMD/+t3D/Sv38AaGA6SeSoG6KpgL9ObT7LtMXYrYQg7172EeGVo7ugeioIFVg
jf85mZM637oPAI9VPnz++EtOtwOvZupmifQ5NABHksYq5iF5vTnIecbnvsu2ddCe
GQ7xAYiI5KNavD3Mq93SbR/fEpKnovFM3rA2h/UQDFA/HRjF1cPHLUzOWEQG9LUZ
kD/69/f2KQEnHzzdTt7HdRJieEgm/R60PL07FGZzgLyKVM7FGS9DbjOvePNMVdx0
3RV8PM0yyRFg9vxUUzAfOb+PdurVt5k2EF7IfxEPKYC84RQ8uyQkDiNSyGJc7GVL
sdUW2I20Am44MFzxGydwvg==
`protect END_PROTECTED
