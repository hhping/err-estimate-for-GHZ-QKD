`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UekMrAnxNq4jHyq0ChdSnblAdFOpyN6vG9VFKqUPX9zmaiOG2xuzryk8+I/FN2/T
g/WSVStS8kBQivW2X/jFUdOFtyx/rH2jWWJGP1AI7OpaBJ4PV6awmJFYo4hYn95Z
63rQBi+iKsuaFHI1A+Quy6k2uzcR+0wI5pNxGcXrwWoRx4hq67yYSJhRgAIK0GBk
zihdUE2molPalEw+mWHnIXNGYuVeXSPttNXtBhvYUB9Nm1+PAki7QHQ0Fts7yImV
tnx0AKiTTyuTe3hy+p1rIVOdWbVOvCXXuwnO3/lePvXOO+pG1CkCuCiMrbadn3FP
i8EZT7vWjm6UM1a9CYBvYevMJesYpOoibDlZRRvgpA3ktacDywpSdFRUCoSk7nYb
p10v1y5zwdG/Auy0Vzdx+wSSimVFbu24JSugalOXc2/gJCApe3fn/+0JPdxdnz4k
Th4yj71KO94fA3iJl9SapcFmgBv8+/tnUlF8Snu+6k+fTxqnXx4iWKgV6f22lz/T
AySdyRigza/Zlrb/SSKbvUmW+XYln12nqvgFA9qCUk5E2AXoiWV8BZXto7Kyj3PN
bLklSuOyTO22mJPugPtAsZ/zK3mbZJ82p/O+eb1yH2MXdGbov/4GCAW7UmPYCOaM
f6fHbwTmDOaLsZugCXJcX4j+Z3Ht8gWODUqN61xVZKeeYTK1Y6SRL128XCj1Ug29
P2yxtFd4+P81Q8uSvMQiAD1O7UxF3gWS6f7cEPJD1GPP6tn132H6spGWAxsTniWO
FAcvKsynE/Sc4BaRuWGPseXSnzxbzXphQ1rePYHHSHe6LfLJhmiURynN1tY9htmy
iv77USnebyoENaM1MOAgfZm98RLv2HrVtUi/rTqwEm7SdC2bXYopUQjpMBJTl+aL
CNEVaWBDWR6Tnl7vNB0TF+MWbsacJBE3LMXleuIvqbvgFpgSUSa/z6gOiPQOMkOz
UBbsRJThyJb7+qPMr49gJE1TVBuVKECF3JzxyzW1plm+hAG31xm3Mshw9rrYvzec
/hVZNziR7278ORsPAOkVP1FKvMUvKflu22diNn831sV9nhVBFcfkdUARwpOtfFdz
7Mp4zK/IcnexvMIFh9XVen8bYoVQcXbKwidvorKwCYcL2Idk3mK7GZ81ZkcR8nKE
/qaQLrpea6L7fbqFMpGrq88ZVgHZNClvU8VXuP5bKj2ARF0Bc8Nm9TTQuTWyWWmF
wW35pJZlOZvHP2O+Bi+R4ayJk4XiqEAbXMFSwS5OcfalUZsFYSiZoMeS5M4gy/K1
cbjFgT98iJUKuX9fjr/XbF5OhaTSA/QNROyNCzmUaScr7JxxjgQzJfetzyAuBPU7
4zei3Fq+FPuHN3XUYlazJSEaw8QCuuvO0mbAuTXcJvXPFN+fD7q+L4BsHriZK04n
qiOOd1cVmnu/Pj7leFrPtVk+e7fwW2aEU+xRs2fgKMVHiuEWuX1YySHaLpWjifGu
4EzK0TuEw7l5no60vI6zojWprwiqAVyC92DNqRUpxVCN8X0SX5ps+1EQXG3Gu3g+
6n0xffzGU7lVVKkDmoFnsgx0iDclnvVuKBqyV0J4gm/hOle747sScY5uHqtj1Lb0
ceXJQ9BgT3jfLHmJYr4FhIwnyldxt+rrdIKa/t/1gVcp395SQVba01vDPYggYYez
ieBGRf2KN5bZFcgr7fnug7WuD+PXPkWb0uPDAuaOQ25XOWJ9ET3F/2yo+DbCf+xz
HfjTccSElO8PYdGDhN4b3m0p7+p3tK2zQKAjQ/vvj7Anz4tlw+KtA2CS0yPnLLc+
dQRXNro+Ex+Pbd75At1P4hrUKpCe0k2IbuuJvcdOO1tFNpVyMr+Wl9hZsK6YWO+w
sZ3S8VDxtRALUTH+iR+8Pacvefr16SzxgwfPwLIy3Ec3kdCcMeAuAxZW7LfKd/iW
zUHW4TZzUfG9vXjQai2tRkmbvNZ8LNayiPHRwbK64K8Qbvbv4x12MrkPNtDMnyAl
nG0NHFItWDbUC1/ZTOWp35Ywo4puB3VdGsyi4Js0vFUmNdLstX+W4PMQSic+nVz8
dobBPAEuQiPUnzN0DqZN+0Qj4a3tNvRxYSF4VFp7zHCOn4hTMfGU9jLeedoaSaRZ
qTcef/o/x2MX+wT3pIRHhJ9YVSeprdA66KQsqsgG9Wmreud7vSzeQ/YppKBmPQZc
RqjPfjd5GZqM241jrJHKX/dOdb/aZWmZ5b2FUMHLPeRdPbGABW9+FF8xb+8DsZbg
puhABGHpHZRJtwRE3J7OkAr3CmJGjjykiPJy3PnpMHCCHyJBNuibdo4mcuvvkoT5
+QWUM24dtI1DLzmnibCUBLy4WZg81cXcwLAwLKiA5m5opPpptWfLef9FgT7QdAuA
eUSEZN5I0n4OHxmsX7klfsdRVm2yzLfZqumUD0XgoOPTKec0VDtSqAP4SUmwSCjQ
g/lY+XKydFc9X0o8HclCNIwqEe+b0LMh3vnywNGk68qEVt0iJej2S1RjlAv0c1HL
fD4n33lEuZ9WRo3TmbZzKrU4NpCu1RlooMvDR8nWacxwRMtsA6F0qA34LX59HiUk
32MlABOneQizST6QY4vksaTVNdilJaepwT4IVeecsmt90RGAhRDT4I75MUpNjWK9
mjmXFfTxKJdyy1dEpCEbee0/BWnYhbuAOHnZya2zHn4bNXOvjWstdPLfraBeFQQZ
pzMaPPWrYzMHS6R7rdDe8zkTbP6G9rVbhKztTpwdChjA1PSkheQOseHPjBVHsMFy
hSFU89OlgdHvkihYOBvaY4aUJwzZLsZJle7axz4VNyA3KQHt8vSEgN21v0UEcNSB
jadeKbt743j4MR56eA0ytptjqY0mjFVwFwiylsN7iwBrRFBWibUvDFXWOMghQE2i
8KKCe3H3dlGd0DDKVQQvQTFNctJSGgQclU0FhS2dySTbJE6FPCj2dxQbiZ3U2gsp
csKgr0/bsixSJVQ3ppLY+46M+MHcLyi36nn1bMa6LZvbH9CkyzOkIik3Dw3ZCDy5
MHlS/QcpKWzQeKpzOmIR5BIHFyKfYwuBPs9uNsk5/3H7dY41G1QsryJY7jVfJTYb
KJgr5cygYUApL5yBeXKnGFqRRO/sywAmRydmwR+iDVxYv9582kgbzYq8d0r7ycPB
dETrnFBFglfF2ltQagFdY1FvQbY0UFx7YKHiUNf4J4LyrQek8EUBsx3liZyNg6Zm
+XI8D5FbUHMdVc4jttTkG0UzIuaE9XeOPi6bJAIyZTNI8sFnpjKD07RiygSjGzuM
VB1qXjqfil+hNiJLSbGw0Y+EryFKiDW0DQtfb6M7P+4qY+QmF+25+rgNhfuA6pLR
oHpMd6q4CC3jYJ0O0o4TJI6fSkUEuTw+KvSuswmD8GkMURU+COVJXJq7UWVrXu2f
M69M69Z2SUSc3NKMTHhl8yR83R/OYL4WgVrybu9PB81ViO0hTlcAeeL2goRFbe0G
YxtUV5LCQKS/qgQPXL4bkkFc5YM342rAmvjztgbPCrXpupQHuEGr/tVtbCTUoqCJ
J5WbNVpPbX9CGapNVFy54yz7+EAmfnDyyw4bxjib3DLyY0di7Sx6NN8knPQbSbF3
2MscjVbuKaD6Qmc9TLf/GAYBA5aHHgnamhUa/5bRSMRxZ5k+NlFppqdbwSBk720/
gPPp8YywGfD4jCWOJf4EQii4iAmpj0NNUinJuIOownFVQtnFukMiiMXWpas6MeNx
/aaEOAHyBu3isgnKrmHRe3FUB+v7ZOTKDCbJWB9EO5ej4nObWuuKjeT/ytnoRAUA
gxkZMF2ZgzevWe4h/F87Yned63OzYzLdO/l3vm9dhLGl6LX6JFDGQpCaie4Y+4oo
I0Y4V6aGOceOzKY/iCOOEnx/1J0/eZCmRESB+9zApPtCDE8Kn2yYdMj2VENirs/Z
+onj/QhDqHi4fjXWscaOXcvthZFLR6SM5fDcag765gQYoDtvynDvqfyU75szFFo6
nRzivLFiGLilhRHhjHGTD44EzSF2yxGhBHN3/KjmSamIAw/SoFEudyw+jEnATLoq
yMysjbH0h6hz5P6UaOFd/Zi251p/FPIgHBc3CA9rXNfqoXBSoAuuGkW9QGjWprK6
rdUeQq5Dn9zXHIh/KcAUHd8CQFMsEQLsfnoi5WiQtzrEeRenfHC9BbbY/mHLV5HM
139Af/tJzvesKU1kNAHf2XiPoIDJmYvJD0RuZFblRxU4N4siQBdEA6FMe+k7DTtE
dWGuIbR6ev8w0f0oaakGwB6K4R4H1FoRvz7nO0epTDc/bjwVCio1TnlGTvhtkgwh
icVo49cM/TazEm0DDpeHnn+YRIdCdzC/G3EsoRA0WX3He3mL6Up5wBSNEu8z/NeQ
ax16JBxlImROzO8E24sW+79gi7Fn2Jrto8RwUnsX2ECg00r/Hw9if7t7YqeWIbGN
fa0sty0UPWhd+ZXY3lQx7diSbuVj3rhkTgHQpPv5+MWlByR0hFm/jBce/eCLFtsj
h3rzDTk2W6HuzOr5eXJnNT7GFbXQPgQ0ocoVmP4HDIn4kdBi5+BdK6cPlVxB+h0/
JaL98vNcu5ANXCe+PNeAzt76XStg0RsprR8+5rf9SupgifHFYpE8kXcueU+Boypc
rOH4M0qXa4ucvCNgLviJuQrA6K3t6P7eWdHfD4fPunFsTgnEh7BpfMVa3JWbb0Ve
e+o8tk1UVGUY+1ruFlHx6l9iwA6l3UCpGLHmERvNGAHTMeNsb864Z72wCF3aebgB
26Omi+yek7U9wztKyFFJXhG/RvVGvlvbLlf4+pEJBEShYyDtGoaOe8fjIrc+JsAE
gAhqbw3nW8lneESiduguJ1vu0s/ScMtyN/inlDvETrwGJFghhDsZPsD2JsAp9hwi
MfX89rVhBMdznL6Yjuupx5VJZaq+FE5eMBNebgTBoW/63I+JJ8cN+4UgIWhlFs1p
eV3TgtQWNF/zOT1sUErCTHJHS1Sm75mPJg2mBQfsWm0cQwNZQX6dDr7AoQu6sIph
RB5SQlQ1ZLjGKlfVD5c+E9qiriPRC1NDkz/w5r3FBAy7t66nurOvMvw8mKlCRiCY
foyX1nNclBCybvqd7E9w8iGjXNOWpg0ACrIQi/BzRKEqQrJsPu+H583tmizXVJG8
3vovpwD0Av2uvXq+Lq0h+yNCr7p/c7HJUG2FnpHapsP9i1i/Uo6mMCnXdm3uPIEv
GkxzlVN6JPc2T6I3XbKqboiVsOYfo/4XUNHSRn0iRpL5kWIdABMBsn5Wm2a9Pc2H
E7EDbM113NLxDCrgYNXu0mI3DgqxBvi1+H4oOYZHlpcaLfFv6tFbEtn2QEw380+a
9jljd7zS3GRp7Vv54lYdwnwPhHszKpw8yB/9sxGX3SBprYdvP1hVILg8Dj8yZbui
UCLs60KZ/f0Ye6K8ZwSrJbdORVF1OSXtqQcm+ocl5hOA7n39z3dBNXaqH3uFLOSt
JY0BcilsNefo6C0pg1LDyIDqREyNVEMDX2a+ZcbLdMJXTOTMDS3onWgLmmpIvNld
3CuHkIbXxzsi/A5BqbZa2nUVRaJgNqRU1w+2C+955C3RFBphcufllHU87uBu5Cl8
0/7p2EXUTJXSsOUGxJKR3/n1XKL3srWSDuM0tJlBacG5juojJo7MOFKkHarIdSNf
QTeHV+YhmaY3dD1d2EI2jrtOjav78Civ3aulR8aXWd/aCMlK5l8enZptjFsssDx2
P8RUt9NvNQPk1rgQmTJOQ5SUUjbg1RKtG4gJ+w2RVM2DJbXqxaTuCtED45dzN9ac
MvplxzuRJjOGb5c2nhkSV7lXC2YF+oaFhKtIgX5XDJEfvZNBVICBx95ihKwK7WKi
sF9hil6tgTrrt473avjUO+7F06koev55vk3VrksJQyJgVkQOIm3XQr11xO9HdRph
P6Ub4OsXc3ArgQHb/1V3x5oG9o3255+jqBRarTKmZ8pm3ZzZU8HEUUYct5BiXtyJ
DmLB+m4MEzuP9veWp51is9rzjl5+YGqVw+MdSuONMtJfonxLgXA1D8o7PI98JZQZ
rFP7src7ZIXOePwZyK7Jyti1qyTRzx4ngFlPghT7rR9hhcwe+fUh6A93dBIDPPvM
JygkpLEOWlh2O6owGFuaNAz0tUKhUda2x4rS8rftACsHhje4EBAe7fsDZSFqU9Cs
fCq58BqHclWUctLLDLVrhUd/BjWA8kuThch6z3W51I1CYp1KDblpW2supfuEc/r7
BqR3Z0mRK7HcagNh191eboas2xTuKSQrL2oWetg8FKxMtz3LGtgOvXVkBSLWSbub
crzmPktOx9ZWPQ5ZmoxPx9WumgEkp6HWcOU546dg5VjyAtdXA7pfiUCO7m2ERX3Q
7T1quwg4ExxjO5/bTMwD/QL/rvBhFcs/bs4D5zyAJJVwER69m07gnSdIB/W+ftRa
5ZFOtZD3+O7fR/gCd1+0qeJx62DlOPfMe+q0Po8W6SFw6Av7MJFRyKs0TMA9Uk5l
601PT3c8SiwSugscaTJ2MiY15McIrOSGaBitqdZ1Ayhd98lFnloomlhEW4+atpmI
2xZUky/hpKivRz7wEObeeZ/63vNtrg6RmqZxNDpy7ikUf8uiB8CcpJmsCwsB/TwU
na3zCxmwSgYhAATW60pgHM+hHwKKchOhzaRXMaRvU5/2GFqyy8kU/r8EnYQqMdpf
mMRg0FX7s0e1KSCvBM6HJQWCGKEAGNOJ5yilAAJ5/vJS3M56Z+iUaZTQJMv9nOv5
37LPSaaaCcbC7g8LXj6jYD2LSLk4oDsjf3MLQsqFCNEQ5jrkMFljb/LzVSRV2Ja8
MjeSewWVnPVV4oWa7bSibIj3QG4oxZpQCrDghLZrYFUUqg8L4mG1fsBPnX3TV03g
QcbTedgwRqCUw6QRfufE9YebiyTf/F7ItPysnFKBI3lekQrhOQG48mXPb/d8zgrw
6pAeek7e+ImGlZC4Gp9Sqk8V8b9cYUBDrQ4qK5nL5S81Jw1C0Q3t6U8TdnWtkS57
QbuEhAvIJ4/S8BqV2JlE5lyRAoSY/Zc6kWD+Ge4IE09ZdjAodsuA+lNmy7mLv8Oz
8wrXE6NGTxbd4emOlPpdYHiy0IoRDTdXvw/Xrgrzjjp4lm6OFyKx3H1E9Da32orb
Qv8uFGYE7aEWOe600pmjjd6yu5XtrAFQNDps7lnOdKKyN37AgLuA2wa7xp3dXA2U
Bq1cBgzuli0s4mRRHqBX3woiqnBgK4bfh8GBlEcAjFZ5vxfHrvq0/35NdKYphLCC
AH0MYLNC08zbOwhGp26dzyb1fyYUGZgX+c/d+0X0XSENiS6CY6NqhWu+YupHg8IA
h2JQiLF6A1f4AyO6kL4IynootJ7ejccijU783qf1sz5FqWGa+l94hZ7Hl1xZTLUG
/GnVV36sZcsamBpChuaude2J29J5AiKiF+ZtFLfkpzFh5nywQhHmOgcjOnlColMp
5r/0AkeEWVA1iQymdEJcMf2WyMkfhe0ux85wIQSLxw4yz/ZMyqQhQA6bWkHyGp4e
q+6fM/OeHbo9DN75cHNryxJ3m+Wi/WahYDjdjLPhm8raOGh3r7hAWH61YTRyLrid
PGyQH8Wajg5Q9Bj1MU+j9DYNdClHIbZ+8oF3VPJm/yqxI6DE281tedvGyMYl7v9d
cjHv6FEmntC1eauxjQuH5XiDwtkfgPDZgJ+u4bpm2QeR7R35lb9TGzhqTq5KPGGG
GOuJKMYlN/M8QY8g14+Ue5YHFh8rEKFFNPmYCD6k/W7bbunXHLupi2Fo7ntk2owE
BgHGaBGJLASGQfNlRMZCXhW8zO03MEXNAGY/ke5WMQwlbzJO4+90fIbC0QH7RWZH
9MrQ2r/xtoxp/ur81bN94RvdKXuC8P3Kfv44NbW0LyW3dH8gCeTo74bk6uBMyaT3
CrQf8W3rbq6fNxvfL6cBIdh2gfqVBE9RsZMxVjOK0/gOsAht3zKubNopyE+gg9nO
05vPLmqICJDvSaWvPklo+H0moAoDbOe/3gvcDvVMVu4k3x/RnrKjVLZrJWM+ImMp
uV+fxH7/6gbJNA3G9LZitGUchPKYbna2YIVTuFyy63WX5IogatCu96+ZIWGVDVfr
5mEzQYnXHa1JMsod4/09V2+WnGpa/1+GstuWB2/M8ByvFi5PEZM6T3aAqQzssatI
ArCkMQqtIxjbaOZswdXjcOJQ7zO/N72jJQq9QJzRddFmZZR6cDh8mzo8LsTJNVZH
KvUBcVN1lq1rc8zk7DDr14LbTq6pGNccVpVG4byRBqV4SjGTibUqFAPLHJizm/T1
vl5Kknq79XV/U9Tz6Hb6wRYw8j+3/dtYnC+ayGSepmrBFq9WM3/C0WTodhHYM0eB
7Xp7qb3Wzy113zEiS7/Z5OiZ4PnoMYyuXy2b8Uav7LZnoUBMMmZZJXdW11KAYHY3
OjWXt2t4oR74Nc078nUh2vMJuLTIfS2akhdcCVgdA4CiYxDLKjHsiTwxoF6jfj5L
wffzy8yxK+TUYBZYOJWUm+1phnFCiI0WhMQ8yQJoVQP79gKHVvkr1/JrnzbSCu6J
RmgsYD4pDDnhveOlIuwDPq3Djcfx92bnNshUZ3AAztChoNiEDYOSbYtrw7wZtybK
aORkxYaNRUEqY8LSvLraJHb1vSYTIJGfmwuc+kPy4x7lwdNk4haCFXM/HW5GmrtR
FKMnZRDOkYXKPzsyAiHkn+vajWLUEfpJOFnJW5kxNfSVAShrlMA/OCIGlPmgVkxv
wLTcsWJtb2wcP7dFIYdlCA4swkQKZnmW5XCbllH58MkQhRGPXqgvnZ4dauRh7DiI
pI2DDer+Dd6Hf1M3PU82jSSzd0JUmO8DShXelLdIrmfmd3eRViwrBCDvHZ9A5ENl
IuDlHTKDpQiUjFBNQD9f5XrRMVgBO6N4kUY6d+yTX4GQbYxijdqfDLGalIWupCnj
UULSjyhKFqiY4bn99oiiRFJ2fSNyg86e+H7qWuyFWYSqQH1PfLyljXFJoHBxQRwn
onR8kPcmWkqp9L2O2Dz+gRKrsd1yjRIHyVdIANS19oNbFrXVw/dVzoKfSqo1DfCJ
Pd7wuvHKsivEUZsq91lCsH/5yT2PvD4HuqQ+2zAMzDCKC8nAoRKxh0rJnYZ1lifQ
Kg7jHvoZqRoENlot48Il+7Q4UoOlrhltY7ttWCGzMVxjd8iSGlEAzzHUQ2rRLhjP
c6sPjbVoaW5h+e6gShlckPpqsGc10DCSDsi57Q1Lbf2ptLjNmCMhFEgN3GkgmSqC
kMXtVWsKAmwhXqtUQzvJFTWMc5C4tfLl4TPWZ0s0AdPRLbfTL5Zoly2tWXoO5mZb
Bxl9CQBetMyrMrStU/h7HhlxDTNQV+CLXzA85E3ZglQ3Y4u4OtRF/gavKZUc5kUL
Ic5y7dXgkBVkkyXjvxPwO4DUf5Q61uqEO8dOCfwIyW1Un2ArDHz1GKW/Wx18BZE9
9E9rKCKcFg4fQDNjNnVOPzrH0s/SkLwgFZ6uMLhFBmhWsvhkI9VqDHdD6p3btfQb
f0RMjUKfKGHUxK8yCzo63w1x3nAJZSPt9lE+AXNXlrC93P5vRVTAjzUB6YqZO4c9
0DW8H+9AK/l+YVnrAcD3RJlgwDZkzZkeAaEZijtbEt2j3LU1SZwFtYRFDB8tbLxi
FxvQWLfOuunobGR25K6Wy9f4s3VJE4v/rGVYq5F/aCFK44d2EmA16ecbBLBMPWVE
T9m1lC5QZJhEZ4+nR+iMYuIG6CjsA1XueARFoHmb0UNwvbzdIEPFl5bapIU/v9DR
5Wvs7ape6bs4mI6S3KvQ6WZidYpZf5Oi1XZTjt/JkirzyzfRKPwSJFDFy0ve8swi
dSRRlIbNNLXInVIXWU2rebsIWOBM1ugPE38tmwAhJ+2h3cph1dLpDSt8tydVmCyy
E/NLT1YwbT4OEjsMtnS7RxfX/W7I068tT7ucUeJrG0N/BsgKZTF+S5MBTSORKywM
NQWyGMMj1f8CiwP4pdqK1+/yqABUEJkAOegJyW/haDIIu5yvIVDiV1dMuVooHQ33
JVyXK1WpQ9BdUYDK0PFmQWYKIUzhQoIstYeXioOMXIGfswrzDxnzNPBAIZLPkb5J
iYrHB5juBEU86j/iCmsmCsnM7iSwY/l4LO3YMyaDnU8D0qeRiD6z9xBRAXUGqhOp
mkFQ1US9aA3oI5/BdxKyZCwK/2+naIohhEhrKNz6lKHIdbpEtz+g+JsiZmbFkWJk
GZWDkKQFcaKeeIRpY6IdmWRDv8UooTBKgeziCNXUPTtitHCIjMS2VT6pzip3HypV
O/+nOtiqs0yu29KKFNlrfEz/8YnYqp2oAiK57fzS+ELELpuinarr7JUjOi44cHLa
wsk1XppTn3Mthxbe5hLwYCrWhtrYbqvvKcgA5nCVqJYFAaGl7c/aBBRnzeBYiFXl
Q1CDhqZtZgfUdsBk5orpEHCmaX2YYiystwbw2ZfX5KiijIa8ZZl2RZs0JEzaX9LB
t+nKUWncMx6QnHeEQH2cbmpXEEbkCr4MapOTrK0elS70m21mEtPt+l5sl6O6xKj5
RLQihEp4RUwN8UtYGc3stYZEMwfqr/P2YYskzVn3LEzsKIWOe0GXIvrdZS+rMGvF
2jL5u7qcM8kmxQoDKSLcoK9OP+3csL03MltEfxixQfssk/MmcK23CqAc77o8hXyr
sh12AlZhoya9yWbGz8Vcc3aqv6+pc5rD87taVnyTG3pVpO3pClHQjh4/VHCYMNry
BR7cpDKVTkR1nkkaY87ujh6/BUapk7vY4dkZa0+a3wmlyPVTRWpKRtQz8JtUp1r6
WOow8Ya3gewdMC0+MQCSX26YxBiKE/QoeFsLktjbT0NEXdtBsdhxXaTQQGlkutNx
Bbn9bEhSE1mEDhAeOrf/mYLw6LRHkBDtdoD8Oi8XOUV8K6scy0oQgi4ixI9PMujM
IaV2M0x/uTSZCFi6sG8q6TOmuAAFJAvdtf4GcMjWoMHITdK9cgmJ3Xcs/pp75Bpj
4Vsijl6fQnHBK8ph9QqkdNoIebqU/3acsCKckLct88Aef0eENXTQyK0dszQcGtM1
6ezLqWyOqfiUB5BiyiEThbMSun6kd7jUQrq7Uv05IJtY55+jj9BekEVi+gMT8/Cb
dZNFVcpSJ/madjbHBuVooJtSJlvTyFZ5AOp2+cO71BLAObYas62A6uTzjAPIdz7o
9NgKFAnA1/mS9xpFimdjFefNHIFeM69uYOxL11wLEiyocl1MGaChgLuavC1IBpU3
PyqYXaFyszXzUo6m9k4UVeJazAJ5pGdqHQ3p227Ue+wjw6xHZQzLGto5MCR3Lea4
aJ6SppdPcLPmdTmYRInYvL6O0HUM1AwnQ7THBdQwy0UNlzI5NMe3q5W3HNrLXLNT
sDW/4HKLBTEa64YFXiQY8xVYhk8s7DIbHqia6HP62zGrPDrd9DYO1LfbUv29b7Mi
UyiKQ9cKchtV+Im9udgXRhVUHhtKSMtn+SnKF/VLpQvDJZDgLtVhwQ2ebcNU02ba
3+trrQNx6+48GVS4QdxrRXzsyyWLUM5bLT/hyqTtSjfgyVDFcHXJJ+4l2g+Lqk5G
U8kVJPN4h2KVYk5DyoEOviIQQjdYLX/SdVX5Pxvcc1+Tmee+bvElFU9zeYgMRCXe
7voKCUtqW0jlXBmT7DQAneLqb9RmzmI5q6Picf6RfRyM3OLzVEdb0F36SlA/kS3l
tU5dZfVW8ctQhwkSi4RG0yF2jUCGO2LMSd6kVoiw0XRy1RE/5rfve3ArLOHF5cJd
fw9Naz3qoaEztPyD8shg4fBmJ9yjJB2Mgd8sNBBD+KTM/djshuHvjqhZ1fRnGTpX
zBingiKrsJK1de2HGXa0Up0Gje0HbABscpFn73RfkdWqYYs4bcIhvTPrnd/Yt259
dNXu4Kzi/GbD63itMsyniQZf+DHNrlmVwIolNRON677GWZUIgLH8bmMejSHRMsm+
+NABFNqABy7GSxMmdkH8QbVcWAudTfdInTbwnp7IY/W4UDdolQ/Far1An5BTk4iA
aZWbzQo+u/IbpiGRW5ZGqszuItxy2eMdExyHIEuV/Uvmydu8M+iD0CTlFTCKhLXi
YLyNhcOIuf61/ZfJC3VcHzSblPgMdG33F0aWta6wY/9IdOwbOFHPTQdJ09LbobnJ
Hu0gqLGJH1qouOsGuUYkwIt2u8+kK9Id9rD9WArRhX5x4wqU10TYyYkx7i4FHFO+
CzlyhdPAB7rnzrSkMsPbGR+cjfNBIVny1UNSb9G1VP2J6zCTAdciyAP0ZKeAS3/N
4G1RIbusnR5siaOj8Ihlk5on1cJmk1DulAwdIL5ZMW1WK0Uutxe2jtVwySKIt3Mn
s+YdkiCxzDUowbKWBjLR2s5GOr089UfQEOZ7rgd7NDPM3FSt87YXd3/b2vfDR0nG
6scgpZOj5fULud4uxgCUebV+CW6E9XzVvIe4eWzb44ugV/2BHxhGQDkayYVT8seH
5evN2VXWcWqCEaNL7UHymqGSfhyGaQbuzMkJ/ncxqd5MV+hfPDBzgUdhGNULWBZO
oqeiDXM66C5K71BnGg2o9SQaJlrnj+RAanr6KgL6d79Bw6gDsw7IM4/tcPVkk97I
EijT+urHOXCdgAEbUB7SV+WRfBIDAXVB9E47xuDakravU5Sm3uK5NalQlJQJhAil
Dw8rYTekWaLwA31hpE1OcQ==
`protect END_PROTECTED
