`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndrmZQ8Z48INVkpqZSpa1Lm2Z+3gwhqQcyU/r/xCf7AHe3VAros5+jNowfMCNLRu
3H7d9cv6CafxTlzThYWyBc6GXWPGadHp9XJD9iiv80C0VWTa/V5YAghGj6VPjVOO
5tLKqnQY0AGCwFihXFnxGTsUFIdlWjqpDovLHxltb9KJtMsjJrnRwOXgUKLQS0C9
0ZiJn505NeVmfXcywoDWHM8CN98uYDuYH8+aymoiQ86E8SQDDn6z8FGUfGX/bOrq
3b6N4KWuEp8AccktzjdEDSkCyKdzGb3inpMqErw5vOJcIYGKgzMqhyB06gxves4p
QmfPOCIPxyevUlkdkkUEvna5g7zdD5GMwJeYpxF3FRuSXIP/M3SkyWvtodENuMQt
t6ySoznFxnlEMY8Ge8Lq9hCcj+VRoKgq4PAAN701NoXlO9g0kS0bpttkT/AokbT5
F5tAWAb6DRWsJTYjJkbUOwZyKtxyuFjIumT8A3nkgetSaEKMzA3Lh32gv0v2HhJd
p3VnkHGGT5A/8VkNeS0Kn7N45YIG3piAu96SGkihhDyhDk6Y6+qpb7krVb0OBpbr
zy6yB0sfeEah+tWkfFaEsPgBdt6GBOOeGoNVVyV4XrlKuZiwWZrrR6ANr58UXKbA
splaXlipNzyuxFtcCvBsDTffaSFx+JOibU2f63/TOk6uYKvzlUjRLMt0osA9cY1v
atf73RHuglRtVRIocTWcLwLpb17kgkGpT49uL+aM/nGWeuVBBOffTsCLdLTFyFJL
6XSexh8aYhp0C/jz406OrnBpsF4XCtSJTVmu/cu+sdvnTi9CvXEBXdw0CiYljUd+
TtrBmw3An1FRNDFEY7PFjsH2yRfRCTYoz3xU+hFhs0SG1YEX1PsBpzXqGWymPqbY
YZzV5+sHRyNvOcwU5R0tS+7+XO005QOpsdZBUgkzhGE18oyBOI96V/f8WW59Tyg1
Fx+3zs1/No351TtXsvFDNwamm1+GokgbYJLbTRyW0Zvrg6SNdapAUO/iwUU+ELCE
CH1eBzhn0lxWkDO0g2xcVDCKm/08dno0hibiYTez/hhr9m2J2z9OVdEdzlgzIO1o
qogjShhBhtTbXEHyscZqA0p+ha+0YuIFeiI/XufIQ6nXDud5YXA9w50Bqg6aIo7e
nOaGl6i/r8zBKHmcLfa0JmkkbYCwFxtO4RuTgS1Cg4VXUr2Iw38vRLcei+9tIClt
sYmnFwL6i5fixH1UtggmMHVscpD2k4FSMwdyRllZj213Y08BBMyHHefT90Rt2EC0
3S2CllrRjDqwzyNYjAuHRZR/F0FEbKLJPDnpX3MOkE5zuRN8v9e/1BbikDBef9vA
h4CPEml1kTo5av6cMnDFbbDyvOS91AcfZLAj4QvFe7uicYWcveLBbbn68BAqa8ss
CLws3wsP9SE8c1nXiGGEgHidQedmW7PGCS88eoqCV0z0nH/lVp/9GITihvf5XQNS
URq8UIRQTUMHXPYWnpDlPgYGREU+XuoF6pUVBnNarTEQR6b6MZHZLGNjS1R7+kc3
OUy6SVmBS/EfEyqun83xQD7dPdcWW8aNP6X+egmt7mDvScNkbChe8RlZAba1r7L3
2LEtciP5zmx2B4AgprlDwCxol6AKrQmcfKau0pW6+Sa4yCBbox0ctpybJHxgKRjn
/TZZ2CdQHDpYgy27ZB6XV0KxiOfiFTGfXJDLhNVTLq/4/6Vipc9qZGngOX6k80te
Iv6CP5I6Z7enun9o3wrtU1KX4hqbWXcrvV1rPfLTmCiOO+vr13IiwnHPXquZ6rEN
3Ba7edJDK8KG8SIypgCSQ9H3kFD2LMyMxpj5fYSxO+yGBZKUczgsErK82oFyGQvF
K9CAIznvH2SOOw9tO7JbfRq9Hoft3NAohzhLh31b3oymTpoq4x2Oh7supY1N8iZM
3IBpD8NomFqHx1nCtC7L0z/vSe8bRzLuYlScgquGwttw9HcmagH+19ROHQZTz5Uo
8VbhoM9cy5Xzxbi4TwAz58U7Fo5Q83gVPGwHGbtd2g2VaIwhQoxYFyjcWxrFkWR3
d0jK41/Z0CQCpamqkb3A/hNWu09p7tnCTwB3kBH+6fHVVe8/D6KJgq0QylpCfjot
aZGTkCLZ2mw6nZkQfJBdqqdcw5PyrDxHtKkynxJSgHgrDsoNrYavLeWUilrF4oKq
HiJsXCUOjqH5rwsRbFOvdxUkTLmLBAAMRyHFfey33R9k+doFmOXul/fXq+t5+HwG
R/p76bqzx2ILbM3wfvkiYD/y3wdDBTbyKg3uIxlBcbOtkXyQwqfJbD4EL3a6+8UR
eqhdV/SKNxcwKpxdSKnpxRaqlUQXjLoLLhWwanRJy9PKC+STW7Of+XTF2R5lf8Fl
VZjJkTH/hO0aPXdrFX18tH8m1mLeaMPSSDVGVayNlAOuCLPkEbQdeq4pAoLHJbOn
+1rXK/JVkVwjEPl0HLcQjcC+CrxYo9D3EHk2ukcAC9aBEXUeAukktX+woxrFuhoS
PPOh3VMwAUBFb5AIMu9v0XzO/9zvT1rJC8cJdRBmK4iVWtBDt+9hotgJjDGWZJP6
MxjA/xjlIU76i7NCN1Y3BGIMmCy8KW/NAdWKS8MvOfOFEqk8E7n5QTGi1j+2bh5T
/iB6BofWyG/46XRNoateNY46qMwMfRM1k+0rSDhceaO14fnvibNgj4GspNehbvzJ
ZgdZWVk7z4Fqa4qlchVRx+011A6+oSCKxIh7GqY26SL4ZZgYzfslY4VgzoeLrLc1
plgCZgzWfhSghKRQRYx4WZkKvbaHcgJDbgBseTU32aoklRzgq3d8gJN0p9Tj+dh2
6CB7S2WnOugi9zt2bMd45gv1jCaOPwVyvB56/2aO/HmJu1NbOoYKPG6LYTWalXOD
4NM2rSI6/YjxJLFR3HMNIIbdXR1Ctwpas7xCAGPKC03LIyTNb9i/0gBBsE0Or2SP
CmnpDCEUtuiYkxlKTpQ9pMme7Q4S4zkTClA++/NRC7hbxDLv0u3pFynAXqQYvqbk
p2rPS0gVHpkn7FDtWxvbysAUACmlkTJbaUsM9PXSt+o9qlNyvMr/igPXvLM19dm5
LSCdGm24BKMWi0MViKdlwQ==
`protect END_PROTECTED
