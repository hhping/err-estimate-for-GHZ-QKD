`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzDGeGsGjyWbqyQ7lN9kr8OqvUa4hTLoheK37auVVRVKmOO4RqE5hVdi1jNEo9C0
bBmcIiz+zPp+I7v3UXe0kogauZ6NMTnXiFdUg5gHjuhDzVbEtGc+Awutmvs5gy+o
3RhYkI5WK5k4eO9w94W0wSvWaX6vsOe7X828/LUmkqYIc0RaP6hgJcNpBr1v5sgo
YTM04MLTZddvniuQ/2vOWNL2GXvNMicY5wDa5xRPKO2K7t6xGFx8EAnvVD6tUxr2
cF6cbX/sUVgvT5i+Q2plYfzFOylIMkt35vBrPCwqLlvvFJsQZqQ83uTyIgEx/oMu
T0a1OvGtXHuteEGBsq2gO34IVD5fYeNunapU3jpx1I0fsm0rx3AJHoFEqQG/0nHd
GF7uwC4vCe7kaXdJeyvptTXxl/VMydAYl23Z4mAMk6Vzbun871tUnAEtnWazefaI
bDL4kkB9zlT35xFBnZbX7Y5xfbOFf0lELmTT8eWJjit1qvaGpDxpgRdinHS2FkRx
gO5GK1JjJeE6URvO8LQIp9fucGB8B/MIMtYOxepRPcOILZ5SQzO/+U7GKQJa31Tz
qekErFwDILul3XASm+rKrFOhOgiu7C3X1nSXjlidvf9hTV5tCYEWjGYgynJ+eTnH
m5xXnbkHHkZGc3UuX9EnuKLr4B89VIN218G9uKVFoV6YYP1ErmzP0rs4sJbrwznE
YsMALSLWe8aq22p9yYSASzFRFdiBwf2YmxPhbWGUQ3I27NZ94mA5nAiw1GTIULON
aAvNTAc+gD0htF+U644Pwg==
`protect END_PROTECTED
