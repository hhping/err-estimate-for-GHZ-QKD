`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzBEh+jHKnQl6dM6KcUuRWY2V/n3D5BTsUdUi/IdKef00cNDmASFBddrZZEJS6X/
lIs8wHVr67C1sI8TO1As4EEGZpiYzJrRjMkEF3FQaqpAbWy+LNxNgW2xNwg4Jw0k
KSvRr8Pp2fen+dglTt2XSOxXot13+LmsGxAS4ClzX4pjq77aMAx/gBgd9hQZRJ0H
a6Qcddt8z6BQ9BEASVH7H4a3Q5U2JR1c1K8hV9aK+338/v6RDEDmbnt54ttnThNV
PiKhRvZKY3Vn3PnNbKCIY5Ynu+q7eLSxlqCKEXbQb5BVInj+fHii144iQPsMiks0
fCxKiduqs7glehDVVb6iB3KDEKZ86D0xwGZY/1vgVYa8PUAJckZ4DJhhVrjclQkA
7SJ35vC2HbeqRhMnuo4Ig0CMd3eE8yBjaH5FTO6YA/xfo1GToaCb5Fc80k8ZFGzA
0QdvQbSO3s4qputF4zwgxE4dRJpKP7FoGccWqx+rafBBkcWcO41OGD2CZ/LJfB0W
CcC3E8uy2d4cDTBtH5VAZDWSD4mVMQoreMy3uO1H4kXRzjp1AcAH1WN2uBxfaYK4
SIRNCn2MbUOJS3bXEv0b8j+WpfbNototMvx825K8q/n9PEzhBCmcca+irH1S3TLU
ImF3RZWgON9PV9cZRf7Nf3UBbTtankccYDGdBEcf0rrSiSwejoMoTKicNExXSNG2
mx2VnFlJNQDjcnA/YbFSGSGcefyG4SnNf+1EIkEkwkzxamKRqH1JMzTJJX+0eQgd
YfEFGdEah4CR7ekpsyi2DdKhXhruP0YrOpmbL2VeS4w7xUUv8uKRCEp9gAKDQSu9
UekVDP0y31qkDo4/UiL/X1q8BjXPhG9mvhxqYQ9iOwQoVtH545C2K5Eli9ELD9CR
SGhZQicqX3c906TrDyDqaxq04gR60idPnmzpMsth38075u0PbfoWb+5Yd/3wJ1FD
7GLKoKl2W3Eh7aGQJZxDECe1YI3o8nS+Z0UZuFW/fXL/SP0mO8ec46HabLgoAjah
M9HcCvOuOo+OA8y8STE3ke8RAjcaWs8t+xRey7eRXWqXJCXIjG7amPvUzYEOMZ6n
LA/qE8LGVul1fa3TVb6yZTfVTdfVsdDRV22hqsypZDJUpVUadPRqF7PDY23GhiPT
Gwn/oqjsThOCCDbzOgLXpkkSlSm1wFpkTV0ZzgQhu5R85yMdDttOWMdK3fouyjFL
IPjCNuvn0Zzj02gXj6KLZ9pwsWHehd5v4TOLcnYCvV5J75Q4v+/+LJP0Cb3JXZ4d
Z1Gi79BEEgvKILMLt3YwwJKepFQGyyZOyrN0SYBYK8zomIEwiTQ+D8j+rCO3eNhx
k/yVzQCNMd5Sl062UUy0ofeNGHrE+tK3YQxFcju5hEPuniMqAFepVwvUil1c7BWJ
AN02zCETal+Z4R/cAPyDSGttiwRg76/yN/K5oFODgYGDV4ZNOkENSfDUEfIuk9br
lSSO42VhIPtonlIiUUa9aVRkJ3rz1X2Fs80kMJlGQyWw3ecnNbWYHok2JPKFUIKY
IzqcIrKA8o6OJ4YTrshjWlNZ3DNg/LWFpil5I7MRxyelZqFeVhjRkwgu08a5eyg4
kFeB10ch45FTl0RQ2IWWtT7Xuwcd7MWkTbufuC9FFm2NKG5GZutvWc7ZSZSVoedm
Gtt6ZtZ+76pS319XQ296cbxaT3EVjMg7z4S2LC68ul+soDrDib4hwW9+KZ7kde2r
3669TrbMHx3ZdhO7eTw5+tz4VdMIvTNrgiv25XJu4SZRvhNGw6VFxwabf4+Wt7cp
LzprDmz+/c6YWfvEex4Mj17wCC1ijx+ahr2DmIQGMpxjc430QLDOFYD7DbVsnHdx
l3erkZAackfbv3KNob0mz+BwzNRh5P8DpmvYlo1Ar7bQ1hFJ72mVMYXclBI04om5
nsVjcezMkVY4kykYPrByRjp3vi3HBmBw9o77kuPJvDTzfSpb5JT3fzG0Iqet3NzM
QxPV0T3HgSbZauo56cyMdwv1/+0U+ZyOrAE0gjAcy6JFNcgdjUp9/WXgTRnfdVwU
BfjPGB0BmdKeHAtILXAQhEW0uzNbY9ECOCA+AAQbzHHhEU701VuepTFS+IcIkbUC
lzkLRwZcQ6h5BM2zxsH998yJ1ilK+dexjf7PTlK5jWn8TXXqfwARNrVAdbIGTwa7
gotafDlSNeV5rY8dEZH0cy4gF9oZK2QkizkwXTHxe9fqY3u8j7HxQR/096wjp+h8
zmK+xEEfNKrGPEC3kuAfZd1Be+cKl9FMECgxx7VRN1lFSZMtmqWdf/2UsARFaBQd
cf/hcgnFV1/j9AJkGwmmji/tAfuTmDrRSGXCgceu6TRXUQ2KAZrQAIgszYzK+atn
HTCNvC23NfkatWqQMThjsLc74uDNjH5oyu16O7iQn2LZM7dArWBOI07e83PGzI/i
d7BWh8D6dlrXMC50NZSzMbhUhJ7VYvP5I2kOfAbpTSPdTzjNdeUeehx9SBzsB7lG
BZXbQ3XU7FxvLdssNSKJtw7KSyTOE5nR+Wpw4ADe1GGVj8ofXyyg7gDKtpirxTww
EgnLvYPlHaHCrDKhdjTJfpDkK8Qg7a57aFT9p/iNgPJHDuU48J7BnWNApOr8sEuu
fhDwC6zNIJMzXzRwyCfl+kMMnVjYtO/0F+lso28n41Ph5cWlwL9Eh4mVmRn/AdFU
cIGbxzxY6MOupldk+1UbsRvhxSgBVJ9WSK9ten3hczctcCGStYw4G1anKB89ZsJe
Fh6c1JcOTD5iP8v6iXRSH3BuqzfcQrS36F1AnS+sI2WLyvWCulF426dPjrzuzCki
NxnUy8AvcdNdiMSTAbZs/NkUlwXkVn02ciHgcVayR8wBd9iesUi4jTdedrgNv0hm
kIlIRuLUrsBX7WEe8UK6pGVke+rtNHpNyYtNyufXW60Wr0Vy8HiM1yOGLYQtqUwy
zuUsVwMPMM33DGvY3gOSoi28Z7SZGDG6JW9qZPuMAm7yoL9Qqupb2oWtf8CYZrV2
XIzFmeDdw3/0h6ujpPQ0Uh2kibQv0zQ0yMKJqMwk6yiAdm5Nms9NrvptGhJ7UKCp
LdLcazJeA+P9Sah+rX8u0iQ4lsaeTHo0VLBTSMt814b0RXrtkF2XKiDtXCKIuYjN
rGFltkTrMx/R+IoupXuLnwkvRX7H0xGVeufqtpAgWTxTuhU7Nr2bfXid2mc1rVxq
4WBTPkz7fKwEkELpZ/UFUgqITA+xzihYDaNg0WO7SowU7fxXkEz0g/EcJfrP1b8D
IlbN7rtwYjx0YAZsAvGiFydnWCPHn4OT0z9Hsz3gmyqcrREV1yPOQ8xh8atShmiS
ojAA0lxzlDco3TRx9/CegYhG3claqMfvXlW4a4Ozi4gNUc9wNpkScrEVy2CXa21z
x5ohLk07063mNTA7zrXVSFlkV5fuI+hUAo09n6/AFLcCfSib+oVE2lkgrBdwoxQH
MXFWTpm6v7rOm3RbeNUrfyZIz8MWS2eSKziVq7uxRCviynAr2ETPj23sPGgn3uxx
jZlk4dE2Cer8Sj5/NkuB9NYDjPyHwf9DQUKe99D8QRiHrzQGlzWEN+UyyrKEvIAR
HgN1jetAE4wZqZQMnawhfKkiwSZXzhvxj2937ypjIafLL6l3M7TGimlA4IGtL15B
ZoQ/HKgQ3BFCCgSMA0eefUJUIbjYVEG0odRIgyNCinEtHAqoQ/JBjpk0PINJDxJO
V5/omcrBak1FyAxs2XcZ7hoH4fhpYYVyWpYuts0QJSI4Wz33Pf/z/Ni3srd50f1g
307ARhE2qWQhwQqeb/kIVLcZFugae/mb4SDU+uXZ9Aanb6v87rtRMRFmS+oVoRVN
rdaRQsl6gHWzHLjue/cbtRqXNhd30dERqVu95QJJyLZtFhmnNxIBMl+GKcCSKAph
mIteWFBfU/NZUMKowL4lzM8sTjXGZ21d6bG3Pp7J019rdu2xJKBg/gR3dYwdoBP7
0CdQbUzG88MS8XJwl9Mmj+/M/+Q7K8gVAfDuN+ulf3U4+dgwa0kyJrQoeRrxI3Ru
jRPnkyQh/maCzYNe9K/eBkKFNqCrwnpb3VescqBpS3Fq5c/SNvUVURtv/+4VKc12
rcEu1izCWHQCrvJqYPWRsuXiMwYBlVX5sUHxTNF3+DGdwKXr/aiB7UAQCN/ikpXg
vBLL9gi0akeRHNFJeMzm1BxD5514hZNLgBZw0Ia2dHH1s9Ag9g+meJXXFtvzl3ow
wmXAintRPPM1sDZ6wV+XokG8zA+AyZLMq6G3pV1d5vJe6JJDHbACZbIiG1ZcXIu4
cm4uQwV+vsKLJG0otdo2mViuioTejGXPrDMw3TsWbbYAI45eChf4PbDnFOni8JPR
a52cvLHft4qygV8KkOyVn4xonfa5og13lVf4oJCxGd/ImvPsTOGzNrBLpH4w2Akz
u5kGtRfBSyI5s2NAzbJlst80MfkT/otcuoyDQ+TiYYDLBvL6n995RgphMTAHcCdu
dpFKkOYbaCWXFCZHAQ4jdnAQbEQ99KEhOtr4hVjoRERuPQnWOlzwHa9ch0k/DCuR
Pb1/mo4kYMFWKOQyyQVU/4BPYMt3udz9RD7bjgBSTG2g4Owi4toMTk/23aozFSNW
ya+9r+UaBNm2NVIhIebNDWdaFaTWjF11+swaQBBdBwAkN29Ji1Z4vGDKD/yc8CAI
DloPnkxq1TvZR8wu9239QdO780BK7tlmhZU95Nrim+4ZVBeZa8/D1hyqQ4BcamHZ
3a9mS6nW5wWUGRZjU+0+nWadWpYJU9LIbfGSe17sNA+5gFTHW/stDzLQw9QHX4Sm
LBN1sDyKokMWxpnzhvwlHD7srIl19pfJ5644b34KADCtalAh3QusjeNt87jNEbAW
WiDR9nNXwO9lCPmqCKsZ/rMenzrZz/OkajeUY9nxMRCOKvKBOvw63sFPsRzN+Ed4
z+2anL9qoTdcMahu1Asso9PHLjfvrdMMgjKD7vgkql4XSYPDgapim7ibPordpKE9
HaP9Y6tVpArwrB5oDEx/ip35A/vvggc8IYRLSg2TcvuFGVgPux25nCuKV9d+7KPu
5njmY+CbAJwQreT8oVDa+fvvORUkvAaXARu3giUX2y9EedWy/4QH+X0DJcLE8rGf
mcpi5sJmEpTgHh+nOjGNSyiB5j2+Utt4f0pQAHbQIceHCo799ttraYCeF8Qxkaag
SjOduzUG8O9/sMYUBG50YNdOnWarEZdQ52ybEmJNZu+WntBNLLJlyWVNFte1lcUY
wTTi9tA0IPLHWdI4k21ESOyp5CRwrO1Z5z+bu5UeLKxnkugbIScnOdjE1Z/voMUn
yTp6npDAGYyI14ZJ6oFKghhF0QzaI3kVivAqMCYQyG9RMekfy75HofsLW19DE8Yq
rH3LpInbhQeCzwcSdDKgk8YlBdocnstQNXYl15dvEy0NrHrRIy2xde65QkYH8JtR
P0gJz8vCRv5R8EQNCpjNu2CREWOim0dYTuIJ34CpjliA4XMMO8kr0wgBW8tnQBNu
cwQraT/H4B+Yvp6oOZFGhukO28tLYIdwAHNrmC7BTbSY/gXNGVZld500R7aIH+Tu
ZI+7CHxHm6FS4d3IqTuYZdwa02xz7xFjC/Dhx6YQbVUDT5pZzf4j8MK5oflEb9yA
JoUwxNuaGwAhgu2eJaOY4WVnKoGl1rFhE2lG2N/kDK+rGD/11CEScoZs5ADRbX4C
pxpVLDp/p37jDGluGjk2hKw37ena9h15XpaYmPgtVHV4CTEcagOyiRZ49NZGcsNU
4zAt7QkL7K2vhVezkFIakID0ezChQVERUxHxtZVTrE30YfdJRNnUsyZXauWhEygI
b5TN78fJRDqz8w9Jd1CqZnPmZmhHyGZRpeV3S5Z+bOibNkeuXgsbfr+nY3dx/RWZ
hu0d+JU3kAceQIM1Xi4GNl1U+YIgatmesU0dSAShV0+5LqaTfu0GEcO+oobgCMKx
/Y/QkKADP6R1a9SGSCF9wwJNiQuTOr51UDerV26TlnrS+tpIoBNEn6WYwiJex0hg
BzbtwTUfKBXEUcSasJs8XgINT2eLmgGnl5iViK1fuG2OnDLP/KDNPfry98Ob5n06
7TI95W0569ko2BJn/Lv9oLSaI8UZxu0jVj+aFV/CCNh83ZHEICUnUeRAcIc9DLCP
0tD0bhKIlvB+VLoKlPTUisJD1Wcc21bHAANp1YXngJ+aKk4vdQctNA4duDrdpCmb
Rt0YhOY5VX6zpr5Iq/GDLvZIK10WPCGBmDSmu4EsVoEsppyrj0O4x9y+IwMNC8kR
h8O9W6xnWmiTzKSoo/O2Z6VS4dTDv1bTkZlUH9MctShZjwdBx2eLpiD2YMGuNsxx
qMKxapcIxUD8uCMLuP37NH7zespY9S4pbwunvCzVU7qyD1jhxHeEST6g2y9o5qdP
atE2muH5WVFd/JgofckFn3+Z2BJSWKCqG31m458suuQqDA8gkavTadNUE2s+jut8
IOJ6JSv3DWmuw28WVrvasvRMcUTxlb9ljBhef3joptg3TGfVgG0SXsOvl8Aq14L+
g11TZSxYz6hVwUQ4bbVZqkB1U1OiP3sMK2yFNq5/aosSxCmwg7y3aXKN1y35Bbwz
1lFzbUO2JDjS7o7rdnEc7BJt7YSQWmm76l24DBuuQ2vvKl8HqgqQLr+4THVHAteA
GMaKobWQeheTvko33nhauYLtBrqipdFU2vnRyv+TuGLjLuh+ZhZuAy9pVmGiRacW
vaBlaHWTNHXuCJZMTzDLR/yt7ryowcirPQh3X52p9uxnB2neoE5QQjK6tsc5eJbn
0EDFlmrkRQOzj4pquv5KmjXrbu+eUUjeIQ3dVA6J+182PBvXF0ltes+11q9yo2RG
d7XhABmiOlpOlvAyfjWWH6bVRLMXjpLTJ/8aDPN4b1aTlq6VKleIyukbJU0rtTuq
cawGcZ64lqa5963xiOzVkjpvNeUg0eL4O4GxoU8K245Uko3iJYaKLx1z8xYYgzC9
MB/6D3fLyJiFXUFGS118mMkwtZZgRbQB2Fdc69JWVGFhgMaCs3sC9X8Qj0okNUEY
bXSat49ZNyg7vgQVj8mfS7g65rQqRN6Pb5VVFYKpu1cfRBsBwR9kCP65ISlgvj9H
TgN4Mh1abaHH+mOID1OlMaIf+U4qaPcSRKfw1f6bX9qaH8OKobVpi6HU6cFAMkLP
67KAKEAC3bMZ6UiqM7EegE+xI7FeHMtNLAgdOyB2mkf+XG+dN37JfLLtCErn6az3
bbG7TByIpe/WOoqJ8F8W6JtAYYCMrCE5t7lXjJGXK4NnrtAHSmqM5JVB3BMgeMLv
srcsVUI6kOFScsScpD6mnARmuMXJzTnJsm7ZoWSocWbVhD3HfYVRCSRuK8QsoQ1a
YOd5AjXrGJE7v33CdsKsbtoEMYO1ePNNzbliqcuDleQyip5klEJRp+QCAgXO2BOC
haHVars6+q3oeT5HLag+2j4cG8FQFEfH8gCeUPDt6urJ1Y2k80Ogz6M/GvyMW5aH
HnnbreEUkHsORmZ0+Eyr56BKCTLRL3kxFk9Vd5XzLNHixoJAiZJKGjfvbdS/Gitt
NxZiuTCfYe9jWjs7tkfVJzveypF3G4BZ67GuIKc8kEscQiLwqYWpmacx1QBVMAFp
fKaOHMZxQJNWS0I+KpWNOCh2O+q/QwSvfUr0rvpbQwN6vCdZkAVjZ0x3iL0mDxZI
+5/k/LJ2yqFibi6q+MoRG+T+HaEl02X+3QgxFiARQuXr2+iE4O5zYGK85DT9dcmB
ZqN/iD/7KCHm1qw/IBJEV129euLFNLRPaTqMOf3l+tNZlEcPGHBaHdTH5zoutqE8
obAw+fZqVH4W08wVaRdCeYMY6fPhYQHtP39XOGaZ40//IiQ91nf6IgEDGEFxjsEH
J9L0aaoUcp7+bvDfAqpqAyOcayqMVTVVo/4RRWHSkCDyVpQeOtZ9NppZ65JxBv9W
78KZvR6/ulCHqH/Lr+ThQfvccvpTaUsdT/4LrgE4fcvkGARhR4LGWo4GltSABN47
ESdv9sLsH8Xp8a41+6FyZDQ/PCVMmt+g56L/MzlC6bA6cnIEI5CuA7eGfb/WdE0L
hLmB+B8fDAhPCqoSYnf5Cq9JGUdwt44bAMFSuJ+2uypGtmC/Vd+Tj9qhGLRnIGmM
vNmmb/YlHkKHt0gSPSNcthacJsisrkXhbuCT2oadKHXRAiKRhsmhXnrGAqFgF+zu
aWP2yr4gk6CIutmCSdfRYk24rtkVFIlY2YzEe9afGDWnggF6BXIgqxr2YWGuRaj0
E+tn0AvvfooA3G1f888Rqm5+TGfXHw/tX8OXLpcwLuny5Jo+mYOdxQe9wEPBQHjt
emorXuu/Y3nGq8rZP3n1JmBhhCAk8HmdpsJDkKUtck/Gf/YfDV5d4U0qrsh0cwNU
h3sTNZo3VbTybpgOj2nCCSxkMI3yUmYv4zGGzOo7v3ym1Pe/Xci1CeKXBoNz0KCC
ksF8Nh+ao37CgwXw3kUkwhJXGGgAYgRzJ6wELOfmNA1hQhzI3n0/u3SrtblJMQqq
fmEH6iTaLlihj3Ek9hfrqxlox6REZ2R3hIoFEpdYvanJkmDstIqixtI5A6iQduXN
W5GqglUZuwc9TxB72vc0Y6VCSthxVxRtkkZq/V+O2gQx+1uBbO9Up7/7E5xjxIwx
IXPfZa2X4c7LMANB68C0vZU/Ei3DympRE2xES5lFsrgrk/IJBT/45vUNQM5Itm4I
qPW+7d2NCWGkIwYopr0Hzt4foAZMEK7I3OALa0vi503Ouu7skx4e4H2iUlhSeCU9
thxz3iwyBIO2aDB6akeh0cRQ031rIjlpi00UW2piCl3C5VefZ6Xpdo6tFb+cLh8P
nbMm/o2KFGHtaTbKkYTbV9+c7RkPhktvtVl/HkVg2gUYkz1hY4laMFgnM/5NLkYu
IQxzF+hz4WQvpdTdP7nh24MZ+Cw2XEDksVuNGeZzvb9t0W/aOukBfmNP10I8TRiK
tgkRAdzE0+W0acM3a1BfarAKpl5x27RLGdqLjSZV5ePpMBUVjZW77o5eyMK2Pxoe
cNNpyuUAixwqcm9uAFEfBP81Uco40ZfU4/amyC4IzOrmiUngVtN+p/+TaCAJOLwX
j0viyUJBN6p59eCrnaKF0gRChE5dDKrdijmpjkdSzndPJ9OtAUYXdSbs88N7CNwM
BW3dkIWLMy2+hFQMt2ongPe1YWSQB/ciZ9Dhdqp4V5lEVG0qWm6oc/clt0i6G290
NXsOACv26nt9KPV0XB2g0bbg4aoJjMKWaTgEE36BQ+Uu5CqNaPV3wXMhpnfcz3P/
9UrWggVJpKywcpVHpCt98q6qFhRSFQv4F2sCoT1QLKSQwdPiSKepil4INGraLMvN
dbshsQ3VBrOCw2djtPgWjXjXxp852stOacQ40YSTX6RnrXiKUUuqkslFsrQZNXNc
lTdTpWrTeqYM0gwCsz8j0b3MugqS4vEYCFaAfPcsfe5DkDPgSDPOZyGpvzG0Vvvy
kjHJ825M+5qcYasfc2unznmkURthBcxwFKsuH5BBO5CnNpQqdTnEhD923s3r4IaC
JSeOLujz9fZVOGHxuoHjQWqHtm5+IrwOlqkc+uronrZYnI8uioD3NCf0Y6bTXbeV
pmgdHWaLTm4CX3E9EsG50jdKZzKrflnixk8TeS+B4yAmqSmyIAABlyLwPpvyU3fq
/A0KE6dgPVoaZeWZOSjVg0gilntCYBeE3yR5YxCOl5gGL3C6hhPqhk3/sscA5EtV
8nsxThJGamn51WcqxFzrQ/zhmr+xiTj2mLGjIlzeqUAOv7fBVi4CX3ucy8PgIGfe
mZpiAGUlOGEqc8Rbfr+8dqeqNhhWfE+xSSiowKF6difPALaFNpXK9OFXYIUrr1AY
UEN4zmFoMra2sw/i8zblz9jIVuodmZ3vJmzo4dkeJBTkq9bZfLw5VHTV7AfC8S0b
up6BwI1nfozU+D2AuiWt4C7qGuN+HOzvyQ+4T/hiaeUVM/SrlkqzNl1ZthZzEc6P
V3OYVXApFoz+4WIMaynF5MXjtcwjvAKNqbdazh5H4/zrLq79fT1ERh1kneIKW9sx
nuEV4Gy7zgLrtqtyeWCnP1tRH89ae4tcuY8i+f1qQvnEZRCfG/Aa280Aj8W3UfCy
GdKPuGc4+hDcK1YZwOfAfXxwenqCzgr0xwKUvY2Hw3yuXCBsp1JCCRZKiAx81O/N
qhp3L2rvndAXskcWOhiMXAXg60pJcPbEYbH0betdRRiZoxMJYM1YpRLN4ZIP2bh5
drv3DtV/m7nxUg5Q9DEQ3w2KptnGgJowokrnqq/bG8+xdgE0NlnNNmvMum1HnLQ3
4Tc1Mqk0ZHdT8HcRkFox4jfgAEFLRrsiwFqYdCoXiWMNRVgkVcQjQ1fySu8QjHTM
lwYMgj1rk1RVHutKCHlYwkF9k9L0Bfx2+xCQZhf72VJuui1A3W4cEmTj7aZvLTQH
R3VIc3Btb0J0kxJvFP39brxcZtaQ4sm2iSGSJRwHtQ0moYSqu3RZ67l7EJqB0YKa
mwS2hPhGLCNx/cswWWuPcjxW0/zDprdqSgoQ09oBw6rQzYnNnDR2Ste4sgtFF/K5
uJCai/+c1uAJFFPDv7lmQd/Ia28ItDuEyiB8rRDrhzj3qhpApD5ncSeI1g7sc+U3
rDVRUSGEw1c/LSjALRqXWwNS/r+np3TiwSLS92vFyhv2+4wovZBWboHJUIRZ1L2L
X9sjAHZKXXI3yOKgcS1fmxTmqV8mdXV9K6zvgurKc31nZqBhcdLmCaWYT+oGuaDJ
YJ1eMUzAi5JS0P4nU1cfzTHkMAR3KgBe/pvyTz/Dg7oQhPkaIFW/Qun6OopdeNrv
eHB0z65fYio6TzQiKCwAMExYmwzwyyj6X0NqCLPED19V07SQEozkyqum4/YS5/Cb
YP0ljXGjppkW5ehOWOlURDGvuFYIOLfDUIfbDUOGQwPMNWS9v4PPkM+V2BlTSbYR
AN1Ej3r6KwCLBkHZuLD3TJStUEhij30sYgRyF7obK/1FApPAyyGJEv3lvsPeMMgJ
bgUgUMz+s7vhDggJ/a3e2lAPcQHrtw7fZy3Tvzz7NjJLHi2MD1ueZ8hvAFcMqiva
PIzmurDtEUhUGmMPT6Byok0eVWm3X+h6T2KGetM0jTBn1SVWYT9L8EyRQ7U0Dlmk
dvT6HGRfI6ozhaApsOfOvtJjFP7DVaEXIg4NBh1AOmUzB58DB3oJuCn5SA6eHZz0
raoa6RQ0mCNoqab+Zojp+Z0vBS/iLJ70iDgIE30zSxLU/XwjKwr+lhXzZHl0zOtN
GGmxw43SD1NvEnLmd2ikfd++KWz+Gm8dHCxqzM/JxcHUHEo7KyEnIY0ARIz+YsnB
wGf9DeE9+6f8gLA+l8PlWVydDMM8KE76/NEknE6CX9dVQYCRsGXYzxXUlqGWPBVq
h9SdiQ6aorct+XwcGcGZeya3BTTUZkGMRnS68VJIItLDZW7ApDMNTptRRkZ4IN5G
qBPqYhFpJrH0aehavYUzDkfJ0zIofSU7/BT+kWKWU2RMsPUAII1rzpVpxCsIQnaW
vYzHygsh1CO5kcD/7hAsgw1qlBYKW10cVKrL6LJYnRB/u53sYd80j5WOpcd1OA+W
c0xnsz2RAm9IRWtGH7vY3i80g48uNHqwJ5Yo7nrhQx45QG8TsgrJ/DGSR3HxKsr9
gOvY6y/PeOsEkICdedr9j+BSoe2+Q44RtP3W3u++yn8G/KKQTGU03ayjR6IK0Rhk
SlaiGLsWQrkGTyi+pL0W5dYFLE+DHdr1JxXaUHdmTjTehUtZd/mIbK+hQ2p1LKD4
Qhpiaz5HF8acSqTzpW3TmQhg8SjB8TMfguPAatCDcLrw2RrMmJ3OiRXkTTLbmndE
3sSKvMZLb0Ee6kACAQyGohM2K3iTh6hO3s2Mkz8KB0eywPBwko/sq3hCx+gN2HsC
XHR6XrlM0xa7DZtzjiSVCX7j33EpnlcD78VZfVy5Q92/vuHN2xKeGfe9oeV8Lv/G
Tj3672/5lnjo5WdoZDO5dz+j4wtV/rv2TOpKh+KOh8EF9J9vhNr3NbJPTiJcpZ1S
hyCoaGzTsFP+7fVjGijmyz/AoRXkT6tIrlUG7++p0xugMjU+Lz2ZPa+7ilt2UUcX
a4LZJsuNt204F5+y+RsrvKsnwKIMGmxAL7JLtaMRxzIilG0ZnXRdl8Y231cJgNll
vW3ncJxJhesxNENBtL2BvfxFXav5qaIp9NfJcKNJVFktvFUzvSCRZ6/l8TPKWoaQ
xpprdk8N2GIbgmxQyH2OuNKYN1WumzzsI8tYAd3k4DgBkEip9e9vM6OTmZcO7tOJ
fGkkFZ0qo6xoEsmUS18F7kXTiPIKESnk6U/RiIfoGqiu8m8B5nuEjTNal8b9CB3a
Gh8Gzccc/uTHC68zWiv/NHdZJoflFNogUj0bWZcH76I4ARDMIiWmacnhYqjOACOs
lCrOCSKYLSLVBwk1vB13LY384+wgrTbN7JQQLpLmxW0oFicBX97w8Ptozoq73Ty6
aefx3zs9QpWkcvdtcTcMo5FoHgF3TMcQWta+pr2W5uyqI8wYwmmS2TkTjB8dwiZ8
ZLR90AVPMbv1fsBmCmQ1AO/rUsZJFPKkj6/QopGaPiHLOWsjeMnuikhDSr9cy9bH
siVtVqvWe7NMED+vHjWExqyF0IMWc+Bqog9roXARmLo4/2TYUNRiCZJdIer3Leo0
MmIm6g8fmPW/4pi4BP84DdnPNKLCS+d1ngrr/nnCqLdvNQYeyvkMFpisQI4O4neU
AEVx/dyNP6XdcYuFu2nKu8j9baDgV9ph3sNAJOTJ7lBYyNuW+/rIhzTg3bq7ERUz
CItM25AVmCFxBGFDoVQmE5i8mV/1odOpTX/SXfo82P9q2hA0OpH3JLf27H4So7rS
m0dzctI1ARN+HVRZlRTjnmBYqY83UTtrFsZ2Q9do3dKScSY0CP9XaupXRZvRXKCK
sHmJnRt9Of72Knyi2O3FHgFhpPJbkIorJ832goKrSRlbmvhO8uj8p7nRHajC+buT
MkHVdEUxRK//fTaLRaqDP6KKmUB15uROXRFu9kaF+tTq8497qqZPG/XokMQm8tfd
0EmLRRbH9AwlHbRYSW0xpoAr6iRXIiqzItR4XTtyVx6poQWA+QZropZ4CWEsCYZj
uDQzw0r2qtANtZq6ntBumb0iUXBlJlFLvwDvfL8TMXzyHuBElawmwed+Dqm8qWtz
7FCuH93h7UqzGqd52Na+HDqZvE+8nXLEQtO7Kh/wflO41oTJIV5amgCt4oP3QikU
X/Inb5ZWVA/pM4M1OhlDSyRYaGEOgSJ9XpunR0swRzcnawhKTVP8/RuRWJ0zJZrD
Af6fMclrHF6NnOL+tak5StfDbabIEDAgnepYdXyQ7dzHQ8NTSHS1C65F629+UkLt
WJTrC3qHf+ZkAMdmcN1NINrOdK+FNaGRAWW7KNQtHCE7yZRJPiBaaNSxEolDszz4
33zAIGtIxmHrps+qAJUuxMGBKHgLd5Ta5G3upk5BQh7Kzz+/BzYTQ/b7RXuq1xoE
titXtWlf44EqmWrTN/vR1HHJYEDvujrs3NQG06amEZjfKK7sP1Ao8DrkI6Rvgae9
r1oJyNm7mbqChE2vAefga/IgoWyy6+WZehXVg+rvh97pgMmrQUY3XSFJTKtPSZwk
6Vdrh9QoCY+M0yUlHmQkBfCuBhuLCcOOJ1GuFZtc9LfyaUh0TNAjnF5vtlPQLcn1
kG4bRNwLrGig2UrU2BZEqNH0fSaAE+n99kjkTFyCxMm1YN9F5Qh2LVhymrQWDf/E
lJKiw4LfDHuKAMNtUJrBp0VzkBaK9zUAln6IJBvTX9IN7w95QHGTT2zUCgt3tatk
Yn5YJwQoQfrkN4lSXmZ3ewEVOl5xNT7pNhQo3O6Va38l1W1vF9G1xqfRP9z1xFVg
PPSP4MzTj7fpto1hqgZIEq097aFMjRc5fqOIT10KKHZhWYXXs1tzrn2oMcAX38Jh
wJHf1HHMJSm0eKsSff0PY5Tx5MRBOUH0HdOjETv+EM+SzsvelvQ+2eM2zP4SatVv
wr8Yxp+gOQ8+9ztV3b3HNM6223xL6lkxCK3lDPYdHtKCOudOniBzzFE3CjzvWqf4
RpuePV9MEv1TL+i6jbOreNgwCdfmPMJ3KwmZU2h2jdG9c7PqR9Aa9zLHFB5gfUgU
tMdWUSVxK3Fmrf3Rqx8FLJ3e5MRdWk0ERDI45CHIvVwKNUUSGhbdJM0lYURPnK5T
znsj66cTBhBMXbjVnSBTj1x0sCqiOpQFyUjYhrRt/G4mV/8G2oyVDjSmYESy8HeJ
+S7w+acLg2kPs71EN7uSzKEFehyxxFWZCRti7JhmwPB8BwMr73Hb11BK885utZZI
b7C7IGQkBGM09BHV0ap/V9B+DAESAaQS8+AjEuxyaeYsgzxnXj7DvG+2+vEtQ+Vx
s7yIhG2SsMnz28tOT5mra1LqDz+dk5VEchLzkLr5RrKD8l/NfMKqr6mD3hVU4eiq
aiJCUuSvatlGfCG5yS5EfK9MdxMzJnb0PMcCOWvmyltFf+Ucs4X8p1sb392GPj/J
OjzlQjRVUa5u32guX9lGL/ZaHLpuzXCZVgVsvA7gLy9Qi9KIx9k61yJrgal2Vk4f
XkzanplP/FGcz53mCZVrAn/qobdZVdHOfnFGP9IG37ELZLCeYIsdPaCguJSvibqL
eSHn6ZIjmyUmxfGCSntT1WbSRZzPkijd5c/KptMClRIW8OGNStbrEEKD2KUSqwCc
oagK5f5EePGjQUTz3Yxd7WvFZqxxC/+fFHPlZ93jo0l/uQ7mTYbf+RSSH7t3c+Iv
ScQt1dRgnIR0VuXMHxXTTH1exlBSoID6+/Xfls4g+YRRjNDckxkW1oWcqhcz/74B
ZnZbwp/RD5Xcn3khP4JRNhxavLHI4EeKrO/HeDhpcbRGutwPgFyeOVNmfq9PVAgr
R/LSYQDF6BVyHWwEgpuia6VpN0MqUL8caD4j+tfnBRzy/Yfv6RaqQ0AF4ROuh6tN
fn7vMaBdi5E7Z+ipgxxQ1eKKkxNsr2ocB2yitJslXUjwfRfW8Uyg/Fqy2HpQ8yQm
7IdrUE+rKZ7QogPLJ1kWRpcvSjzTL93v28Rq2q5X22rEAM4uxV6mBzqf9iTvNv2V
aOM0ji57giNha2SVzjN+ZKudP11XzsBYxKqOcDOz/lbL4jObYsabJwE8o4jkQIVA
tmmkGDwZF6U/QKGl4j61p290Xz5oLHHHVSkOwoLnyh637yPGBGq3CG86083PlCo7
c9zOZgSnXzeT2jXOM3/a/KCyBLDEHxTMiIhHiLus2MRlkyhxQWLRfl8a654fFRfP
rLAIi+keUmyFw2uEURj0M/OFwu3z+eN6b2+BcHk5PDP8qFkMeORDrcnu78iUe27E
xzHf0TVKmgIUaEM1RBAo2lQsIIaIqnKIoCGiQuOg7YuNyG8o4KB5XX23jEyUVzkc
5AfqMMF3amrinq2BZ0eyzqIUPtAtCVEmB29StWJY+Km017jZU4ilhEsT1JjuYC7x
R1ny5VACIBEwvRkmJ6B+lyc0oXDs4Nyd8m+iMXek/O99AgDNd/yFOvAjPJ6IgVbo
C/jw6pmlpqYzzVsR6H/xRcK/T2m3Xcfwtg4AB/7YDV2MJwSgYTLq4nKqrJaXB1tE
eXpk+f58OUntxDbENtYkqzMgiNw37STGgU76rvNC7BtbXjLutZVq0bO2xhJC+ph9
HRpJYwk5D0rAze+HDhWj/cPonwUza0dEG5zYY6fYahiIX0EmGjMvYtQgkaPHV4kp
uSRCsjbF/NZJ3RCD/HJ/mpXaWjZemruZsjXwseBRJlAysQQKzD4Ar7zO9CYrioGS
feyJelonffZyzMg5ibOqSuXHuu4QUvCyNZ294XMEfbaZXl/Zzj6LM+w8uFukoL2K
/ho9bgMx2eNexa+wMwudZokRkgACs0vwFXyGhaorpo1kV7P0GPGAAl4KQ60oMExM
6ndCnzlpX95nl7TFrvMSXbzvRZIt9ZXcIKkxaHpUQt+p1qNTRAEHXL+qq7TqZ9nw
uiLaafqvX07brmfwZAnRoaph8p6OogJyFSyCRLUoq33/UZF0SLkUCX65F72JN4aH
f05TJmyvs2ThrV1GPutOj/FnGp/E0gMy0kkrxTLwpmXDKzA37VEoaZLiA27TEqlH
VzfO3m54klyAmjJ892lZFztRR6uhIeM918SmmS7ojECmTszM8h52Tk7TTEOCo1M4
lP0qJkCqWSRIEpejZCBafo01c480M8KEGViBx5dGtsCP5VmLMArcjqLV/I42VupA
EZq5IP3XQfCjELgYxnfQ/5jSRf7EL8UrewIrlQITZMAHfxxjMGIta6fZmdhgGQiM
UnLkhsYZ3r54dlWeqOBnRm9xjQPQ8kaEtgRZx5/7zhamDKHw+mLPBdD+IUS1owg6
MKs8tyRd8cfe4few/4HHz3qEO6baRJn84B+g8l+msBK0j+ZAmwD87d7ykDN9bVVk
A7zsUxMU9F7rU6rt9IQ2I8U39pMzDMSaXB6ytrdrUk88OpLwIZH2iPt/Ys5d10Kh
AL0Of/rd8vQiN/1iyix/YKhcOjf/c2FuJnpBR9ehV3dojUWIpYLJ8AfBCPSbOHkj
H+9976g/UnLWT6sP28DnhHZk6zrXo/x5zpDjk2TykAtOgg/OHMWZGPR4Q3xfVs8j
JjV3no3TSFdnfDN5znOzIwsYoAH/1JmZgiPsIiqyK82k7r0IbuUMkq9heoWyeW88
MxkDLMw3x0u71J0C8uOy87q8ObqChfGgZ+izMTl8lO4HAIS4rorMw20CY/EOvgIg
EyiwDSSRWa4xti+FjNMwY7AMZ5ikkZ7UcpWDVZ+mgWYkUoxEkjk3K9J/xFz8XdLK
fW4uPaC7YcYVrBBzgIV8Xp5gv5N2GTfCGYV4lum63WonBfnBpJaezSaYoWwLSQ4X
TXJixMTVLuAvRD4fJwZqQW6WNvEVBqySwb1hHmDJ5pAemo63JXjN1Rq2AbQ8pR+h
+c0KN/LuNQA75paagwnUuv0VJaF8h7na8TbPwCw4jPRzHnh1sCEPMy3dslwTwzjO
XJDi4D7SWjyJNW6ZKH0jPme35FUXEOOWOgJneyZNubshC6pmN9MvPrNvJYGJS/QP
Uz1LBKnDif4F1TZ06Pn6dkzjwnM1EZwmQVbPb0tsbmq9pB4R6sdI6Dgu6QHmB/gv
jgxnKRieZFHvHPyo2T0UoFpf9WkKbyXLu2F8T4vkhHZhavDRKIba95Aa03+nlIAN
4W9qwzj2VbwZaZFOJ+fGMK/Rmk7bfppsDdGgFa1Ie3+YpdXmrbN7xg3IIIuJgaZY
Vs25CYr2NqVD7o+VMlHzL4Hf+e3flI6JazXaeV1zl8h9wUfCg2/bvWpqw5QIg/4N
Ws/I6axXB/NqSBhNt0DidvPOiXw3OrsP0z2hsQUKfnEX6thMyhsqdyJKROrsfpYO
iu360cIagT5jWTLDCvbRayRwK71TuAXnxXxkbqVTC4C0ujmd4VN7/gj+XZYffI/R
WVoPpH7vdO7R/nJAkZdYHOagzN/goPLBXB7PzCKcSMC/Sb7QlfiSEqIppyie/nBA
qqsAQF7JUVCXbxG/gS2474XaU6IoP/7SBQhbVy/vsy68pfvhuQVuw9rdiN3Nc6LL
iQ7oT+NK1O2ZGRq4q/zMDVHSqd5S+emreQ5nErHpGnaB0u75xNzeEhzLqHYpxf2W
WoaW6Ot4BMlzqbIraJ7qjy3ooqtYcZ194IGUgWNcqONt5ekcYi5RvALgUmWOQxsg
wLvQIAB8Y9hBtzJNRV2gDiUZ6Xq8evRDcticEuizWcClRKlskzkv41NCLXQgkBZ+
cXIA/PhznTG5Vbbl5UUjzFXBNzmtWR5QGp0+/mhzAdI=
`protect END_PROTECTED
