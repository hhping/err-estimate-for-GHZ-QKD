`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ea+uRCcoherJUCqDaVoIPTx8qzVbMaeNSPRxURHigkvnOn3b1fYL22oBuVpVKVGQ
QPheQGCeIevIYE5gJ42sa8IrPOV9Wqg0a9fMmdT6OeZFBq17kGNPe8/wCdi+O9zF
9fCp1Aio/o9zslk8VJcLlQJQDNV5DnoVmH9DiNdGlF66m4o7PUbkmppl3Gd2lvHS
yqppKHvIYMOzVu7C2T8eLnnE0kGpMlguZoMxNsnVF2qKU8xH91kIsuU9GdOz287w
NHlIz/WVl4OJ0J1N0Oyh8vsSe2l0DujgjWg+cDuaqwOu/Kq4audGqIGe3kM9mFxn
dT6YZzLh/y/QOe10EPuSU8pIzPPUZvtDYpCPWqJN3f2jwjtl2WeFCZFx18Blb/86
vkKKnIe/UaDZxpmqg1oiOT9sWEC127hfnNwkHiUxiquRCaVsZVn07qbEryMvTdVk
Z1s9PRAvxFG4t/am9dxEWH+gDvGgzypX6S1T+1HLUJBRxEQWnBC6TSRi10MWJaV0
jP9Uw3wcQWnRdyzkn/ilO6VITocVcxaGYdDWcOBgf4nYTfmy3WNxcef9ASDV6Q4Z
jkTaCSKF1FepdW7Vj1RQyblGgEfFCYj1cDT+0ejfgPnjqiqWRz5KbU96vLpRzy/3
qBrvEKs1yBhLc7BSMnZNQvBCjbNWMgO46cBepo36ntfOn7tWf8G6tpK8269bE9V8
G6+mfyMbxztZP1mWoQbwIQ==
`protect END_PROTECTED
