`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/US8/Q/JCXYiBlgM2wBmLwwZ+IbGZZ7am9CQSnXTtHp3U6sHD/XByN4w8m/iOrtH
XsDGuS0dRGKOig7X+sXGqr/qgcnLpew3qzpn8FLVcbt2cvq2LntTmsjgdNlo5iYM
QCjz1XLaODGIK8LPnicDn2gObErorrjLI3swp8DBHQ1ih8utfn5ZW87YIibGZxQx
1Us/AEdXGjB77uE3zA9xZLPEM6oxdNKTriTfzxEtDvQ4xq5wK96oXcRwUarpyd+P
urAfG5qLHU+i0R8XBv9sDcLDzdUn9Aj5WBSjYQ1o/0sT80JTulejd0xejD89H32n
Q1NjtP2REL2te8kYSwRtu8Zzr0DSX4w6/jhq+i6P4UlGUA6wEydRF/PWSyu2K7Th
VFDFWVeSaAEXPZXc12UorQhP+3fwqCIXNThM5miE6HQOYNUcQ3dsG5gsoz8Q285m
3HUXfRYI8HRZ4RGWmmf77PqjJMw6FwolHa9cPtSKpRfGcJQdYGjL5C+ZugGylYDp
Z7G9sLHRnoS7ejFmgKFQvla9e4bP8HlKjd6ITEZ2u3LDoSGBs72E4SXdHbhVF9jI
l6Zf0b8OgnBbi4jqeqOml4QSTxRUtPARwneofgBApR27w2e7duXkqGr57fM29hi4
Ir6dVvkxHzW3+rErQ231/Bpb9jqtW6x8qZcIGZ8gfw0=
`protect END_PROTECTED
