`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0LTqzVJFoSQyS56jK1JtYihXacejce61U7IQ8urBl+1QEMX1uOHLfbjU+UcdfM7
xQZuIVfOw6ZUr/sZ4ewW7zr1x00YYfqayfm4URybORyuxMIqY4e2aiFZbeQmhSdn
zG+L6yEy3O8hHN+HLzRqsAzBHvT+184SFMX/1YUVtlh62ARqWvKfPAZGEtc6hU3M
ntLDzUjiiLAhj88XLqjQLRrrBGGsjxFfqT1IppDFYBW+1Gx0Jtf0Qg5btce+QJZK
3CucR5v2tz2aD/c+mRSCYtWHZ3B6AWCNFnpH2D/ZvvB4o1qNYN/6UrqVwuOK50qC
HZpBwQtt01WIkhyRc4bEHvZkohtMfp087TWzI911I+R7/MppqZYqxDzR8x+R395S
`protect END_PROTECTED
