`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pr846sn9XVNjWhctwKIRUrUiix2+c54dnPtwt4no2TjwW++DjewwSCVYhshJ+sig
ODnBFqusokDtdra0BmUFpcjQiVK4XOcFwfpUJKArHt7aBWDqPIiAx3IbrqyyDJ3l
X3G0gS4VpVWM2utWpB6j9gf46zpVB9ftrwKc1ChMVEFH9xB+0SmxF5NDzLmuimGh
F7ZvGjy+hdJOPXm2cxiupdARsVfjCBnhgtjtiJ/bLrwgPV2/U8p5eDJB5kkCGuGB
SxI0kxcCt34WZiOTOTHG46Mn2Ka0W8X0F7UP4/AGemW3YF5eRC8+OM64LRwl0q8e
kdKztmLUABylaQpNChmCTzzS5BEST+6cuKf9RFQEcRxMECRJWY0upC1bQAJs1NxO
WQ4qVWM20SVxcP1zK7s9jlfamstcToCCjHx1YV3qBOMum97GroHmLDalzqBso/NB
3IJsny/JgTTIVuqvPVCWJVGthg9jpeE9twz6D12AvusAFEn6bBGOH2vgHSziaEec
Aj2PjfpXIr2KzfaqT5IR51Za6bHkNNT/UngedclntV5gucqzqO43cOayNfcn9+uZ
qpKqpqVzRDnd1SvmpTaFQLMrBUI0Ikvoi/971MAJxNoP3TMulRmQoFifIfJH2Nf0
LQP4hYq/UD7FhqSFDycWxTU6xGybNMUV3+0Tv6A1+BgYWpODKrFizwZPUA8LE2Q/
mlqXh+n5cQaRICpZWuQDAieuBFwBzcPijg9klnSmiIT+Vokzb2KeuC40vbuGT7Du
q7mXtOCYwfHJIAfo3KqiAz4mNftAx4swKQWXrdI+2lZS+jw+3kr6Gn1jEknFb01Y
owh3RMGMbldOUAPAFYnyJt0tvYnjW9HbOb2eXT+rfZ4URiN+ASOKv/20JhQB2LHF
UXXHrt+i9E1frYpYMMmBMOMOT2NfOaxmClxXtkGK9dK84b6JQoJvtiPB23E1Q37n
70RyYBEcSj/+a9IC3zisxvtNa8JnvUBIUUwrK7wkaLkhHyVkq3D2KzcMgMz+wo4l
DFiRHoJEBMh9Kqn2gIbSg64SDYw41DrOE8smirVOaa16Ly9Q7bWxXu7wnolj7lfi
S2WMS0e667U0elfnux5iKu04Aeo3w8oXq31vt3UfkQ8/Fze+peMdhW/T1YkC3q3B
GoqqfgKshZt/FCI3YHTcBy49rJSMwTcnSriBSRC2lhZSbyNkSzISEiZdyyo3PiLN
DgIigXgCaHwBgx1QjXv8BM2sUbOOMhhXyPtuUah/ffoh+ha0T4L7RvLIPOVMGPAW
KyoGOM5VpIpuXvEai4YM2w8tlOKj/HXfb58GP2U3/Q8+/+qSchr7iWYhtkWzvuGX
S8x9SxiiKfc0sUShIvMMmzjKYpIGvXw3wEhD0Lk5IaEvIaq6yLd6JqYZKJg+Y5M9
y7QZ3OeR/SkFiNYyxvXzU8XiqMKXvEiqEp1vVf5d1YebsbVRskzP4OhL9u8zYtH1
RAsMEc8gYg0S1t/gyQDbb5EiuqWCxtij4IPq3fMRpaO/y6qCWwOYDfoeaYaZg09i
aYTnvWQ4Nd6iZLoc1g/sg/LbrPZ11oc30HXoYEHkx0IPgTnyi4BEYM8JWJk7jHwz
C9Y0Rb6P0D+X95YIDPU1VbI/Q7nmbqbdT0f0I64L+edY2Q7DLUU5OWBlzPU4/bL/
EExV6wgSMHhT0OEfXtN7cVvmDYrcjAeMpVhHISZD3iPE+MAdonHUCt3cn28k44My
42xQqLUrCWl29Ruqy18+P/HwwHEIgDdi1gUMeR0SxHAMECg6IBwRCN5WC7zOjniX
wkqEpsS6Gr7RSSS2UQX4UYyoOi+U0aoLEYrk+fSAOiQ38hYK/uK/Cgzak6nbKOWJ
3adefZx4nweDCilhtmYQgx9uWKFRARAxxammXv7n0Z+xGrdOLzUzUEpd6TrC8Zvk
Pc4mogHwyRe+QsqCqcB2iRepyXnsWQJoIyN9DotnQJqTFVcCYWlLO6fzFxU7F+Si
opnpzLCLS09CCRZN6RdWlXMyOW1BNGtCnatgIN5jr3CTi3kN0wGUm4A+Vy4JAfUO
1LR8L6G2YftSYPKMQm7fSqBy4RHKkdNQ1iA5RUWpoFirM4IDMAlmahMakuCsH6g+
hwaGK4h+Vr6YEX9xbXz4cJMJZXs9TfSCYK6qTB2Pw2t60CiEHgfaT/q4I25aRLDs
GTYTN180+ZYRybxmYk8qNRZECWOk9ckrE3YiXfwyxOG51wQl9d4pQ2fBB02IaFWv
cECopWDUzJ1CxeV73O1wQfcqYvWi6ZImUFk0NVGidOyCIfQTMnJ6JaU5VY1R8ECi
mGGosx3jeQtCbJLPqhGELUVrkkT2xrggTDMUrdZ6OHRs6mx4SnYNDlx2hzHtQgo0
Gv1O6KMkHMcmoI4IlN/IDdh2F7gSEWGqulxITL5QQwcXInvecMypowfT5PoBkYBd
2ur02IMf8U2qs0yim4A7MsSKYMiuN/ie8aWbghY74jEmjGODH9pnKVTuCzBfQTxz
nP69D6pUF4zArz64lDE8HZx2TMQJoS2diOWROsYPR8Ic/12x8eh/nZ+YDzetSfWO
Ej5LyVMmH6ApEs/MowJylhs7FKYjHNGblSsUl96cpaaJ7zLdIBKYiZI1Jwadd+fx
Fm8vsi6kqXjOebdjphF+7iQvipjFU/8YCTzrpKMf5eNLTMf5e8CKwCIwYjErLtct
VodHixb/2lfS/wNhjgMBWVMNJP47IN1Xq0X6bGBU9UAXhu7Ss7BP0ZK6MlY8FOcg
8mk/FoSMvBd0B9TWversd4MyHLvssYRma+3BgLmkUHdMpfGpEsGat68PV1WX08W7
O0r/YyaIwcGsEiUqwJdH3reHbGwhuOvaBx4ZNQ6LRV4DPEAlzta4AUf9YvIobZkp
t8hi1Q1yK9qqdWHrM5LpHvx8O4eSxVSsqMAyvg6bxRkJwnoiYs9DprCvY8RiFIPa
WfdXISb8grigJg94fskCUlHVx2+rcVvxdzfc6TKSGV8seA/a7urUOSUS8LeNZE07
kI3Zppz92xtw0ces/UTozCwyy9cgQa7ycYmhcdvcESsFZqIWFyBVHbqUyQCX3MrJ
DBJ3DdPS67XDkSI/+YqiFZKFJrgddM9H/Pxag5hDMQjkzcxPRYqeMso5VOn4ZmOv
fufSwZo1tjLOrr7E61GnJL5HeuMYtsgXe2nAtG6kFJYPLqTm/TTaPv9d3QId0Z/u
jo8PcLEh45uIjxcKh43PAGQX5cZu9pHlJQoO9MhjNT0ETE7XcVr1Dt6q7EdNSwBs
oCQfsdejrC+HW/dyoFxlh3ZBd/+nJbuM8/u1+/jAkiHT8SWU4YFtTYtyUIexbrBh
i3tOGX2yV4odv2ATNbxxDEXj4qEPlxmHqpUZ1GP9eJFKD5eETO/RzaygBLMvM/YY
2wwYT0aEgd6TNhdDR2yX+Q==
`protect END_PROTECTED
