`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B7ZIQ5XMo/Ldo3mWx6ZCjCoM/2ECrAAWXv6WlO9H/IVgupaU2fLunKPhMeJpk9B+
2fpMS1HQ0EJIdQlxBGyet8j/dSn6uoNBFFBh7y3ID00auHXrNf7cPLH5RsfdHE78
o5DXuGseRlrZg0LNDoDvzU96Kz4CA6QjJTvLa24dIXCVC0J4v/El8CpOOTYaQ4NJ
db2s17h4KhbIvrRiG6yLEnQ4v0kc0rhsCzSLg1Fk3T1OECpkSGCO/GpNGXWjZJmT
FUZtX6slhHmOFH5C0AD0Z5/f3RaENVLXJ4dcwoz0m5cjOWaLBZ6d8DtiwfqebSTo
t90xjVr3BpAbD07lIGY+RNqLRBgduXAqjpVy8KuxDKogmJMtZyIaFeWhLwZo9/sp
npRVx7QPiYyO0XqaU5ifCq9t7nQ6i0fIZx5yo5vVRryobBoevgBdQHGjnJeALI2c
lyHCUwuTC5SXfPICJg9SxgJ8Yf2hxX4UX2z3qF2YVW94tUYkB9jHktu5YYPGbCpf
c+BZT1zJm4oysGoAhvxFoWag9N9F12E1FsJfAchihXJHG9O9t60AhYqss9625TMl
GJruHFMIlriYDXH3bcWnUlNfZRokTbbiwuRz0woNlwVgl7rXs4adudUchZ/nZPK4
wfzmcXgmiarymxxfjRljaAaJeg7ynNQduso3gRtQ4D6j+NyGBo8P/6UwYYw5Jc7e
7CcvUzzuGXHYK6A0vSiCYTgWvo6WZhpPXOqZsA3yT1xX9jJ+aAPiztmjn39JttT7
V+M4qDItTXNFN7jck0X2jCrAe9rol2Ng+rLComYG3cG39kjMWgEOCT8uedUtDIlL
HSvi8GWwo7Y4+qhs1Vi9/hgpjQmwwl5Yx7Yiq2dsZvQxbOVrgsgtuX9vteYD2rme
egv24JsY4aM4UlsACnbpLM37NrjC/IWBCeDPn8+zAshV6y5n07xPe3wEBKk8qhTo
Y4FZWo6csuaMZljXW3WcdgQxy3GiKI1XLXOsWhgavjodH9UEh4ftAmfoe5MDUSco
fSJGfVhMxHTcMTiFTaDWPcQd/jQoolnD4MpTRsL5EksQtz7GMABbeMzWK4HzSq5m
TA+qYBaL93tbS4tUq818rjM9W/OfBjNyud/9T1dFHFSFfZeqWGg5afE05LErU1e2
BPZsLYVDpigsl58rLo4HnoV9G8hMfyM+osDWG0kdLl6hB5+JqetQy4c4n8PwFyrf
FlmvavB8gClyA4A7K7djnJe/+q2PAQ9GNr01EPB2Yq25g/pwsEr7uAHshx+8WlIv
/pqwj26DqeB8g3xwBlLwma6OviuWsz9CEVpR9GVcHxrTC02Mvkf0sHuYKqvBDIBe
iXxiP3jCpdb/w9Rw5gWAWdERj1GoGXUBRzwqK8BG3e1mfnl/RFYvJR9KYhQ1+0HK
ucTW5Cubafx52Q93dtyz/O+KjscZAXkfzerT14aXHZ9CpJq4caPIR6PM4D5jbYsR
4FSz3Qy17vRlXQ5BXPye/50z8x1psLKOONrNE+JxkgZ7dDY8jFThHu6A3SQzCndy
58F8MjRTvCO21wSWJJwk9QxsA44bL1QbkPjxQWUBQEQJaBz84ZwuzCYHw3TONOOT
xnrtKU6skkJfNq7Cve05Z2ZVgte0zZXd2u4DvbWecQ8rwjc/2L14XTqjm+qYg+Cb
XI3Pn27ITd9L6PnB7Es6XNG9sZ9iKCa0b/8vGQXA8ToF10JC2HVzHUc8xZy/Lzq2
F13xEZ7pwdkbKxrUXu2FG6xS3Yy99RulQhotICScnvi1LMnoxDioE2sRbBE9/7OL
QDrK77iBAUWhxQNfclYSJrUt1gMD/pjIC30mTECIa0pNRIhbxgIFNbXhHop3TvDm
Can6NiNclSHQL3E1BTJO+DXKL1NUxVUaxFyQqaEAiiAyCG3GvcQJTHQ4PlH/e7/4
zEaN8q5tGkLhKuWUiIGZcVzkK2rf7mZKct3xmhXKJOxA0dK+hD8jOb8tbAK6d2E0
Zhu7mpal1gHk3nFyA/sUS5KKTeFoxAKv2WIKbRrAMMwJwZGvWdjetfvanwuQsk53
r08hpHqm0pahvpPaME27EFFl4lFFnxME/YELkU3Dg5KX0Sfg15e/jSgJvzmBKb8X
L+gpBW/s/6Cf4aX1aVY0g6dnZOnO17YrSrVgWp0mEOJCxz4HdDdvZ5Sw1Coh0BnI
Qk88ES/XCU3iOUc0hTMeb2+3TRzFy5jst0Xg7TA1xNjpvMwiLY5vblUZNwwHLPbv
SANvt7PUg+Pbkge97a204FbfDmYyVdZ/S2IEXIlRaQCHb35+7dJcKg5TZNK32Pou
ICU6jpGoEQidXpo5/3XdT5ZbFfQTTm5Fxn0lm6+A5FE+1SZKKBUZnGoqp1vIvt48
Q9is1Hhu2TIfmPj6IaS3q4GGlGxzUd76LKVFk+pD372FXJLBxiNzHInRieiOq5cU
YybjJBcfi9ZX9Cdy/2kXufN1pAX9tzMYHwAFZV6drbsNVFEO3NCiYpZxKzxUYZs3
hzRJ3eJETG5n0X7BnDtSn2PLkwPiCeAZppWSkBD0/3u4FpOjkQ2XkJkmff4pZGuF
uunQlEV+I/MZKq8yNSl8umcUlPpiINHGH+yrY5Il98TBUvz8LSGhTFAGjfwlXTTk
mnqQxrOHlKOEho4OiHKjJ8VRdjIX9l4dApZLXY2A5I/V83Clw7Te779OVFurG5Rp
2gTA8U5G0g0B5cSLKmNcGaOUh5FOWzyAD/C93tUunWYqBYlGBXFlW0eCOPmojDHM
SoSS6RqzHyXj20C20t68Y6xVRk5atjw2ywV5IlT0kBUeoB5nKkqD3GhJn3KQwqd1
`protect END_PROTECTED
