`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
COvgIwIL1iUmX7x4H9tVnftj2FUV/mGwTSOUZg7XZsDxQiJy4aSjnYPS2Na+cdCH
grC6j1xWHaEEYZyn5ffAqR8E+cpIgtbf+H27NQhluRBt7SgOyKJ31uF3hKmVqB7s
onVIurT8Ci6UTLmKRT+QEZte7OrWmQ45g7lXyU4pvLS87b8WsNOrIBMa1q6mpzZ2
pJtjA8q/0crkA7w1Odu/taFNTTijZpEbeioHiZGgXqnT96R9w2CByTIAfOSS5N/b
yheACJP4eX6PR3b5+Y4aYHTXvCI884wEUO6HIjKO/F2WbRWQnCD63ZvAUmuMqcHT
YG0VZPXfo9jzGaAyLo60Jb+JGIYXOHHZJTdPVLXOg53yigSfELPlndwm1F0u+Fja
nRD1XMd7C0MVByOJrRH/U1CIJsZAb7rAVaEVaPT/tVW+jtlCtPv1IUcIrllc/zxg
9vqHsqEk1Wf+h4aA0p7XTODgK3F25El85YvJDCYdcn6JaUAAU6GTMFLW04TcoODC
1YmrkfowAYF36pfJGs6Xd6JmAeJcJqhdShamlwl6UjURYT/Uf3075qvWPj46TN7D
8vTcAEMCEpg4yIxiQvoV9rgkclevMAPldqb3tBFTT+7j4YJXgTcsbDT2zcG7kTQO
nNcMjwNcd023B9Ur3vhs4YA7tIuBFgZNtTkt98ixlS5poWVek8WLYqrfOQ+hXgMM
eu3KamF7EYpXwUMo4GazUYkuYiswLbqYW/ZnGYUbpc7qXwj5i/qXG+II/E/m0Lh9
O9rwReoq0fDBm70Ugwkw4eYegRqUJhT9Zx2EGfapEuwPbqf81DgLiL0vkTrmedZI
1COQnNdgJQ7KTY72MIzzWjY/lJZQ4dQFuNlVs7O1hCnfXRcJ1ONgkSqLPEfZcbhm
c3NX37Hacv5BOUfVEBqsrw==
`protect END_PROTECTED
