`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ePutPiGw84oSJDOnLy8FGuZ8fVK1iA3ZumGgV3BavYLB8n4Dp5WIh+UvNG/CV0yj
MlqipNigEW3Zu4vnyJQRlg6LQqtw9j7IFvF62zcsJ2lcpDW3aRkyC3q5B4J72cqZ
GIJxVTDjQckD8vWx1hVTUyEgi/ao6ttCDIqee6KQtKxExcllv5QBcH24zbuL/drf
yPXoUo+cge3/3otD0x8JY8hOzisaOJT/MA7edvt9npSn3I2urfFTV9pBKE19o6WQ
rYl78AoR8jJceBx/qlArSuNnBmuXjY6AcTVaL2+Bc7pSDg3KvBaUjnfkr/Oqrap0
jkSVjfe4AOwQIIWv+7GzS3d3X/V/H0vf06yg9GBbHzjjb8dkIjcjApW4diIHZik7
P9cOqQktob3f1y0X7rpH9CndOij/yvi6lrzbgPWxW/xappAAO6AZM3FEm1hia17E
HRBm5VOEjeDeZzTCMEvmHtHTSqBQl98ZNZBSNye5zcFI+rJVLnkP3onk6ykyCmSM
edMV9M+XYaB4ch/SPfl5dslBOBGoEy/e61N+oSlklFJg5mQlHE/M4sPs+bZ4RXpY
r8EtH6L2udtl7CiJa5aal4EjqtBOetI/eWf0h8Jc5grk34rn6O7nyKc3YxSBm0mF
+T7FsawPxJPlOgaqkXdnlyx/JsHpe4EPC+15sDzTd+lcMpOCqwvYzc62v2QevJzx
ZQYVlSiEHNqpoPQrHxsU2Sj2oI05z9VGtyOaatpZpCKbIPeUmpLx0FM8yx/gAKQo
tRYy9dcLO4gyqnqRBrLZpreTPyWiZ/068i38xRxIFO7uSsMaqkw4RKe9OaTtw68e
mAJR/KpTa3Ha2T6BafnPDpt+XCjfZqivw1Hq66NSP5TPo2yS4qoifc9DNNvgmWj9
XeIUIwTzGAACe3a9i7+OxkFRVWb6NanvIC51Ae4VRsz25qb6t5KH+OFsjOZXnpoA
SOIjbCMc8TQhYKJdTspVbWpQ2ibDUCryld7ClNDGWBuOMobdnbp1ldi1WvJ22mHu
5GLrierDpDTADLlCfXembB/gZZYfa94vicaipOc1mOR4GbpcoVXIBF1HOkqOIHyQ
KFb00Hhrn31/V5ozYYu9OujXS2gBlKWAC+4d/aoGMWsYGLmFHW/y08Nc5BE5gM5h
o7W3xi/+8GqMwAY12XRrtX0mPOyAxYNLroWZP8ZcT83ZtochygNZKT/Lc05a0zt7
LjowuzfiPa0wnKlP9G0KCzQjpmnhmzbXPpsxlro3mY139KlQt9LXga9cu+lSKHzQ
gyGal+zBIt3JETvOjZ5uOIUp/6sNUkUtEFs1v9JBP65XZIPD9UXryt+1uXRBXETW
wZE79yXRb99990HRVp1Qb2BjZ5/NhR8WWzj4jdtMk6yC3qMl5zPaxvbWngy3SlYI
PAFWYxOZqCv5HUF4OnuBM3qgI2FlB+WitNkAbhEoC/P9iKnOrAKvP6hTcegqmkrc
3e880dFAmOqSPGiTjNoo25zN/1E2aFFCbWuODfs+xv7O5TF8On8PlgD9bxJoB7Xd
kNp6XLW8QWea35GG2ID+P1p+qw3QIqNERBS439F77rldnP1XL0YB1QkSrrVzJ/9M
cXkWibX5UWPvmpN4B3Av5btxM1c5IaHdYh+LtDRH5gQsUQVdXSfrSCd4PjOxzIMH
WGee6HF0d1JAV8cQsIxkC9/iQJCWbYEYUsuVE5n5b1/fNCrLPOncySaC6ny8ECw8
6Vfma35VouQBbm22RO+M8R+ivdHakVutiqf20TAouLQY0eGLcaDuQsmGqNVmqNqB
XW+L7J5TxCXBOLcN0xquH4E4urU75TljfLdb7er2YVmpmusWaKpxKeS8/Lzb3b10
A9oRYdO0RTFvYtiJZZX/mA2k23tRwuxsT3DpEqueDGohjSGV/C2gctzmAOgg7tzv
YdBPCuejga7JqfE+F5LnZAyrDN+Nxx6FN0kgdSd2P6G1cjehNUMze0KDmrvVxB3m
tjlXaZI1xXWuHt2BewM0kIGIpCG0ijutbRpltOLUT6D49s0nTsMeuP93B657kfRG
P1ZPz2fN0m8Gwe2iitXva6pNJjV2GbYvVzECxy8bzzYOCO4fRqu72yxSfqFbvqBF
49GLUTlU8pMMKNwImCGZQxIbNMLpKAODToPdDfjBfiG9bF48FULkr1wDUHePiHAo
8ABoOqTswUZbCmZlsq0UGk2psLVmvePcRbk6fm/Fdg71r6df1HwVdhWpMEwGKqnA
ADAU00Cze7TU3ITJjRB7vp5V6NCwYv9e+WGo9UfQUoHWt8hgHH02+EFVEPbyDtb3
rkaZl/83+ul/nJcEewWujhIc+FRco4EoJGb68BFFZTRnzffZFvzRKLKtPLdRydSG
D5B2JuD4pvHGaRHPy/xU+t6crtT5ZbP6MA0XRioCBztmlPyWDbp8UspppgsqsyOa
k9psg6IBop/iPfMnpEUR8AGDjnrR/X4z/Eh4leqeqIs=
`protect END_PROTECTED
