`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHq2PKDw/ae0rhRxTHiJS7DKOedFeIc+TKYC/vV873HYNsWotaDhBZpVYTyC2SKb
77T8ToBhJmRIlSNc/L3kD0JidNDo13fd4RKbjXFAYdxc7hw/loOgYOqTfr4YQHlt
28bXO6UTzdVMRDOIzbek5yD5hNr9L0SJ3WnmE6WwDB3OtoV4/vhXqAI6bebnNinm
4npFbdDTX/gJSU4VHID+MBnGGH4GVzuxyW+W8mEv5Ac=
`protect END_PROTECTED
