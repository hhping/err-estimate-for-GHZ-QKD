`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJXs0y5JwqtPFxtcVcgoCGjeUtz3h7XJ1S+Lvt5FFfz+AGlNmSyogbw1em+fF5Br
fZkwcyaDVu+SakQbkAXKRW4RDB0mS+5kXB7b79KIBVxzW5bosyKHjyNYr/I43+FH
zA2I3689IOxLnv8SEr4JbjoSX77wH8arJy3Ech6kk1OjUavPZLcK+c7BolD1rWGt
B5fP2159VwZqKZejazYoRgUtG/8BziXonjiETer8jwZbjJdhWVbmad7MaRdre6x0
gvVWoeABHBktjAE6UNNwg79uM5nOrEm0WmcMM+pGv2+cDt3xIgXjEf0beS1sg3tO
g1haVWBRx4yxF4i3nahtBdHgzgqpqpP1z8DDcdPCbnYJzZZJ6OkHQDeQtblg6s3Q
wq3yy6wvF1c469JB8w49PR7Hqm89ua9X1h2vuSNqOrxmZseyyjAn8BNuUnm/XS04
WVLAQJis3dzwdGAyzIWTt81XISjxmPdOwR0aAsYwShsOECOVHaWmaWfpQjqBoUMf
gcqOzRjtf2x950G0IZYMU2Z9CUg4dQKdBauMGvcJtopkaaTDP8R0AAT/0pSXpKpo
y/vY9pJYwcwCgnSFBXpH4mlttW+OcH4LEaufMgOEIFRDLY0jK1Oxw0F0baNNNTGW
zpBxpjquzqr7D3MW8RZ0VS/UDdy5/VG94lLrJb0SaMgYW0tHhY/dIkxyIuJqrEMK
57wOcbyZ8Kry0w3XlQNdqp3gcb+D4lVmFSYtsaCuoUs0YxbXd3opuXatbZs5Iphy
weNCLYmnZNNHOynByxuKJbMy4TLFT3g4WfWp14aMsVSS6zEudqXMSFUooEHiuSW4
9uW4w28XB/z36C5TkvDipo1CsGtSdHE8y1+6K7nqa1ORRnkp4JbzENUfLS3DHD1d
J2IYbXcuU2v2Xuulrl0eeS8yEt0oc7EzCWe3qLMqfP7RwaHqwxkzIozLOgT6NYWx
aCxetWhlyZlnbOPVR6ZxviMz6T821lu5Ml4lpa5socBfm/xUWnp6+nns6WoqmXvu
ANLw+xuBZXjCEbt1NchBR6XEllfhncRNKgB61TDcnqE=
`protect END_PROTECTED
