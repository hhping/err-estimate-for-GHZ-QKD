`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8nt6YLZSVj4mXNCNLlIThFS503/Ep+K1uhvipVFMEmYdS8u1fRg0peBKMK/DJW9
IhQkpZcwARB/MJvIdJxzmf/tKQ0TwUAcw+wlfJSFl9Sl0mnjTEZY64abTypYHEAD
jFCAGoUldnxOXWUvGrrKrnH1n52IbhV2yevqpMvaJwUZloX6TBZ6AF5mwVYgy0ux
5injl+9yXsQdGf8lJk2mJFd9+gf9n4zWH2Mo2m79bP+Ef7kgQhGuFP1AbVSFPhb1
0z69xoH6BxFdgN6+VlUKWkIxp1J9B6oRgc0uDuH6jXKnNa0mjiPYyWoHU2zvqE71
tVZZ522Qy5WWX4U2+hNvO2THB2IDqHsnQ7p83Jwv7ukVehl7Ar3Lkrd+cCSgqh+q
Tdr+bk4LgLFxF0jkNfFQm4fUo2Es2CI/4vyDq4MHQmrKwtkwPgoCqAgovlbsnwuZ
S/3aGdHQqkkxIAJaI7fr8+jaBkEr9fiAxGkPTXxcd3kOaMw7cMreXtFD8jXTucRD
65MX1oUaS0k4+Poi00a4H+e85/QkNV45jbO+9Z8fsb4CHTolEWi1SvZzshl5WfL+
gwx7TDRWqVDUC+dNcHe2XVlwkGms/X2yPQTgJhcT7Br0HfbbS+HGqhIeFEAHPE7k
HDHXVt46H3o+Tb5NjXuIkCxpDbfzLE8/FKRVdPKIU5PiYkENf56F20NPCLYqBStt
3oejKZMgzcnI24mFEXIDzznfeB3cG1oltE8kRKiJqEnAN//kzsBMS6YIvJj1cWq4
9OGjeh+5HIPLnsXr2WeiYlMwIX0tr/Yadc4mfjW/ctn6hzAncmgY/LXvpLPNggTg
Ann6gTQdZgC8XxgYuQ/aO7YnxFQEr9iZiLXF+xwkgS+XfcnSYWYWgDc5qbKST4OT
lHip614fxmP58XWgiQ4tVz/a8iiaZE6zFmvD2Mq1COjBaP+7b1OA1hTu0ZMAXcHk
D/4UErUkfedjFAseYTjKndVMNI4Ykr/anlIm4EeguuSfQMDWwYVm2gZOKm6Ol8Pk
rZNKb2zSSY3Tq7ECYyqwKr621JVnmzKRK9J0xwxogEqNjF8RKJRZZQmj2693L7D5
C4qcTPGAJUoiIIHeLXXKNUkxOz4Tz1cOTP89MejZseeU94JHkz2osLTyoQQ5rubR
6WrAG48xdBLz38/Fer1FrWtocONJ9Z04cVC+ej881rKhblNILdeP6IyavStKCDui
9juziN0xtKI9tzeYQfzK6bq0mnm7gzac9P9M3R5NV9X/rchy6LNhFRB+C69xdP6F
FLPHYNlWFNP/ii93b8ABLxxl2fDjssYIci8HtredLFGq0lRo9l3uhnJ56mlWcW+g
GLXmM1ecCwK5bk3+1wkFLacQB2IUrvtMFJhr+pbLCbgNm/oQT8QIhZRrFgmcWZFr
T5Lswvu3z8MtzmXyN7JWygaQ/qr9kU8OO1vJf4J+TsZjDXgAj8bOVc69Cp2lZnDH
gp03REcDPlZEVZWr/lvylkH6ECwlSXo6ru93nsSsL21yR5Yr6CdxJE86Q/T7n5D6
rZBG5e11185+7LyGjb7qnI0QSukJ6dpyOjYpMBdo22b6KMBUneajag/K9uQqPXKo
BYBuVKh3xX5oQG5uc412QngikRXhtli5yPjB82jfNsbW35pP4/kfeGgGYxb+dUlV
8Sp6/vzwSQcAeX8ldord62IXLgFYX3Gcr9YX7ilEbMI3XLsWwEeMfoGT2k4Zb/PR
0VVmuBkevYtH5W416YdCZotxM6lwsdzXdNmLusIjJJ27sXJiVp2dgKM7SOz6+DhI
r0qs6YFNRDH5bDOl7TVyU2ENlCAk4s+t5E5pWz1iBtH5UZl69wJQILlRWhwKG5q6
gHzfyrUekXmZUL+AFP3f/e4Tc4ATEpPYFSoGENUs4n1wFqdaOA2p05//dMiAEqWB
O0HtX5I78AKQBOFh94VdThZnM05ktcwX3jJhbanzdxWa+zVywV1C0Mou3/yBVtwB
`protect END_PROTECTED
