`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5n3XtGjMx7DsubIGMRRJ65kn+U/PgQLF18J3R+EicBOZOdwbgpRakln1rDNokyd
rKF+V2decwfq9CQ3eNANEMCMHgnZs7hSPw7SFC1y4ogRtGNzmFxTSBOJ9jjLytYq
Jpt43Itppb3lYu8JVQ+jhIlibUsSdJoDgqoiJxohGVVLCPeXkqXa90YVOh9hhLtO
hl3nD/SQGFAmSyv/olVe7tdbMOQYeqVx2OYsapAprCRBSNnDXGdhOieQat6tlSfI
PfZER3hbcYtX0bKOjsNQizby/BxKoadumcK5jXiAAfIfxH+lUL25NgJZx72Mgqag
if1rac10088IzhxMlwvrQKUvyMsTtyHFLlk6jXumONWyGL1RTteumAeQb2bOe9Sg
iIMDcBQ/Lq3xiSQs4n/qmukZhbwJuMVHN+NCug1eZcUozp5jwJ8PakBfl5o6pmWC
abOgkuTHMJ4kbvf/aKDk5SxDLGfEFFWEtNHZWaO2tkABVob8hPVw+GFePvQ5PbgB
ekO8YYslHKqZFmucrl7y9y6cFuJx/OSQJkchXePq4rjHTUhvhi3oIpvM71l+8TVh
NyA/Wd9mTxA69fR9dGbJl+c8BK/YwjubREOvZASiGbzwwI8kRZADd28H/0ipXhdJ
W1GSSqsN4vq1zClQUipsvfiSVTTNE5vG6a1Tp4d3imDfWmOEU59HHu4M4Kr/RiZ0
X19onREyLiH1oxZB+BAPRVL3JGOs5pKAPQlsFnVZ+MsQXfK6lGlnFoYQO1qU3dX1
tENAc03XOeDgSH6H3I41EToA6LlvOhg4/Bc2Pahl35gKaJxAxLvK4Rx+ihfCKJye
wqfVRZNxDxB+Hvkwaqv9BsfemJpebVSM49xRbTUSYw4uY4C1nL8fR8DWJp6tZT4p
bYVD1up9HluU4vb3VCUtBoa+oAaB/Rt5Y7+8H0qpK7xig58nTFBP9zojEm3IYKLr
R8gHrR0WdpZLSuURoc7LKMWgKDs8GeelpYKCwvWkWntBi3AOw7yYcIYGdijrFLMT
xVV0W5p/Hu7XakIyzalMifOG9aKUC88Dku4Bt3JjSzb1b2Wb7DO1uuFFRkpvG+OB
rPLWQVqdKGsG67YEs7fore4W9goMmNaANpAc2Wspgh7EAQC59bLLgokIxWoxeFUd
Vz/Hkl2kv8OS7NPgSVoVLd6TbsRmnpD4JDISw8w2k+qpcFsqRwYUEVtjqrXSFx2m
5bthN+jZyMSmn5UR4lMjkyzjA5SfH3KJ7BK5mr9pBj2zV3XY+NMLoEdDJzIElB+S
RlDyvGDcGoXhuzltw+2OlXpy0WgA3LM+YkjCZ48AhEIxnLcqMCmDfhcYiJ51rGHB
967dWRuJ8S31mMqwFOPUQSJRI/LMQoE/ADCsP806ZMxUpJ2jLYe+kBGsKXcOwi4H
QrMVLgr2xy5Dh12ekw1Bjw==
`protect END_PROTECTED
