`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
At2CQbVMVhVpo+j08P1+OoYJyzlKvenFPX/ZNdxsabnNZ9LdMHGwtgtM3m1JTqBA
8omS1sOTKjTJaAJY4s6iAHaDwDqOHSJMxlR+dYy+05P9gIZcc32Y4FpbDrGB1XfF
9avnc3JHBR08RYwUCyyQejGMw1b8EBZSJDbTXhE6rfTHBUXfYWIfDxm276vYYlNI
3jZ9nBQwPNOj5g09kncWrkMTJ4KMs4IWKl6GVxkBX1QfNyl4D0uF+zdUh0X6hUoT
Bw/xd0PobIEKnQf7xNkbjVGdZIbitemVH8bsX3oaZqVe1sTwOV7GH8y9W/Wqmjyx
vxgIcZzq02rDicLTdmU6mTw+jrcPzuBq/i9qY35pKQXUNt1hzbsPRxr3iY79jlMm
IougtK29BQBS4/AugZgAtOjeaDTF0CQcyx8TXaBzy6M8PT4ZZJRewqzT5tkSITQx
deeWZheQhdaart1q2nKnmRh31JHtg1C5edgSbjaVTfL9IPIggHuqgkPzBecuQ/V0
Fx3Eoivc8wFBisblxuzGGPfAlyyMBC3fIYpyA+eDuA9Bgr5gUaXqReSFF9Y8je+q
jacI3VujMzxtCcr+UyEm9LCjn4KNyC0EsV0nvms8CFNIOx4cN+xOtQoert+2chxf
e1NZKNGEJxcNPzZcATrQSWTF2fKWchqmLFZuLCU8tssmITFxzWKKEkzAaBy3OkMc
R032/6gUrH4/VepDP4wpRz4TBQWYZKFhp2i3Xof3mP5Ys26SlAUUJtMFu5CIlpPw
osBWflOVQATJXBc/cvnfhBR0QHi+uuLEMTmKLmpo+Tl1bi2Wvg4T3/Zvtel/7S9l
R+HrYOF80NlljOc0P8qZqfH0QN9yPDbtKwmrdG/3GoYrKNory5s21nKn4J9xHIaa
pBHZbfLSWTNbuE9ElcQefc7Mq+TReCY0VLEHjxqjWUXnZ205AXz8XvmZGRZ1byIU
1YKAx59vGpoR2jq44qY57J/OsEp+scmNVlcoayPKi5X5XQVeOxvDF0WcVzBww5Y1
UgbxkoQ0s0h9TREpJOLKT0b94++JC9DY1qss4uooX2AQY4uKE0Qe40e/Ogl45REI
Q2nd1racfSPGUjSOScd3WpBFk+XAJ0dXAJF9eRsp4uSuuGBBsHr+nbJYM86IdBnb
`protect END_PROTECTED
