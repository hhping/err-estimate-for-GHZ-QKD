`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZImDuPP8+a0sPl1MaE8Q2QVxlv5Fv6YgLSL4uU1hBKTh/aUJGxTCFNqcHXqZE2v
2oCyWkUloZSBR+TGim/4+ilCiNqG4XzYijKpvmQZEsmuAsGwMZFPSYMQ9MYt3jYJ
FQKMXWDPT7mDH09b+rPdgnZnNVhH+YURD6zd1SJNeXkSUkK3bpy7nD2OpMnjCfG5
9IfF9x72574SbDbe+iseKHhj7D+8uQumd2ajA0ieOO7EW3SRsV/dl19pCDAFGG2G
/NATEduh34LethWldQTOsJP/FrgRt0QwOBAc4bwD8lTdsFg//nzG3KhoBypbAPNA
OZ2Qwjey5OcL12RY+bLz+eGOb+bydLg6AVmKOwTVytG8aoXlFHSiQvOyEseOMQDf
mFTs34LLU7FHOk9DjcYDfw==
`protect END_PROTECTED
