`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
szRNZarQyy6srgKAxyVDHdXFjNVy9FZjp4e77Rg8Pgb30w/i8WYBdkmqLQsB44z5
sR9FPCvApVvzc/zwXcqPvO33H6XDW8BN2RJPEudVOoZ79hjRfLv415j1Xfpd02a4
NdasMCztQiXjfAVVIqGFjMYj0cjDrZ1UNj/YIvo9FZC+4BCSFzA7r91KtYENYHB6
jxzZR0U+BYApGcCYbkdFE1z4tcjnGLCBkYL10KB5DiP3t/qnPMXL/zdIgT+1MdvF
H4uxmQUGmbdYCJ82NMAHj+46yJwx6dUs0lxfWpcAWB2OKCGpcp7gVUHFYoBuo/7x
9PhDxoytWz7Ef4QRRtMBWsYPJWzu3K7I4zReOaGWaxrIG4UyT58QiLWybPW3rHuP
4DSAqmVG0+kZ7KOW0UCWt7QuXUQF0TtMsg4En7+cxyRVxmR20YY8GrgmzHAhznEu
cBHUaRVj7GQZ0PXOiJVZNXBhhsvN8NHqzR5ZhlNJINTyOJKnSo05d0W5xa5csVF6
2UGBuJMp6m1ZBhez0iSbhzjWw4HLuIzKxufmeIyKwFpQGyKEBZ8O6/17H9xb8Ivi
4fA4IlLZPSlPFy5Ow5457a/kfNlTPT2BJ5M78gn7PyPdS8NrX7dDV5iK+AZo58oy
C0gN9tHSDlrVhq6rI2vgTNKgxRmq3Wa972OnxQmr0AgtemyzHf5HQ4o69GsiqkdR
Dt5JlRBipkY1wildONUgHzdpu7aH4ljfLgNYRRzWXGknLeq+039UPHTCLT5r3jLb
Oy/5Y5AJVj40+6MxsaEpgXDc8Ag6An2W4jMRVeHQM8zIjj/h20+zDKRvgdmEEB9X
0vE76Sup1LfjqVTost+/aeIKHkDUc5OP1aTMCAzcjPNvN+foVjU8562lRG+RbzuB
nKlFVJycFzmg24l0b4ztLYCxJfpZaZNgrEno2IyIwkpJeeGlhr1igoEy0Uf9zjNN
RipyN9SeoChA1unZxzr/DnUMMof7LszX7I2KmKHkldXJUMuBOFJaQJZ+5YJCVu4E
djof9nxi2GPgeQllFN1kE0rF2i+xj+cfA6kgQd79Q3Hksafhm3USa4gRdj2L6P+i
lDNgMjfq5DpzqptXbScTmWNdog1ApEJ2RVlohQ2xbDTRSnB+4qdNmisKYdNE6W9U
2aMZ+oxq0gYP2GkFBH6NslVELezffzveMRhf7WSHodxR0vepkkEet3AmHKO1XvYM
E3GbPVnNkSofUt5LbLfbn9CrhKUuKXoQi/8ARcZPvZ+wbcva7XIgwBSouT0QWnBv
741gGlsuYr+vF3Zp+ESmimUhL2ov/9t5iXn+s0nOmfmFQ2Af+CXeo1CzoBoYbdhJ
bF6bZeiFrjeGM311ldx3MewYP/HVEOfkdqXKlDyDu/IVcnh0WzmDyKx95h9l9PXT
Zo+5+4xHvFFnEPSkw0dK9Mf0svsXUkwYPMBsPsud1AzlyfEA1+gJq+4HmAE6sJtN
eg2NIt42zyAKGFWHqv6cn/N7xvo4yspMYk0nziS/Ow2mctP+r15L/eI9t0Lh3Ohb
4m3qL9Ea2utqKeSBk68p4LSmM6ZZ9hS7SqmyR3eab/FHsT/yAMU4ZSi3uhin720D
7BOpKirFb61cCjv0nVNQ5BoEzbjXpXeLWuKfnvd99Jw1/nw2Pr9HWubVf4L3dEPa
8+746rvfLkF1tdxd+h+1E2ZPLhCRtCfoxOoB+JqKk5sJOKQpoLhLPIxO2x8YoVut
Gy4Tmt027SqjndSkYBTnSGqDojaaBHBmq28YkwzIhzPsCxgzLAMsXmA2Szr/0NoV
1RO5IJGW65idknEXV0oMIRnnVWsO8I6aP8ctKwFk5H9FisekiMLf+RZIc++lz4T1
eb8mLiS29ThxZmwW5doWCAQkSIvofA+hA6e4CiO1j24xRIHbLyEAHnjJxqf9Wh6q
`protect END_PROTECTED
