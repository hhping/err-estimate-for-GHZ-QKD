`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l38bdgRhzSpF3TZhPpc0wEMzO0uK5CT1TC6sac0lojEzKqNF71r3humL96P9Lqz3
ENA8RweqkyEAjMSz2TtvGH9IoxYcjWwuGOcxpI8LB5K3TXnb8k4qBnUjvq+XidvL
Sb+qTAaQD4S3fwDDICfsAqU8+dPwSl6ZNfyfr0ssJGUuWJfr5GhIXhvrwFhqwUPD
+cUoFVVaUQXzo6/oGOAmU+Q9LAdDK5HapLy/1PoULeDsXG8Lk2rlnpvDf8C4xg5E
dtAtrU0gKDfJD6Yw1qztoYlU8+U3oomYkcU55xPZTM2/SfHgDztnAFeqFqah7/Fn
IjSBI1ZUJDFjSqycRkDWTT/PSL8F3R7ZQZQDhuzlElvlw0oX7eoIU9erEZKpIN5n
hLlV5it5v2zGdAoMxJe4p5uTI2eQoV2+W0ucihu/reVFQNyvEFHGafpgKVkp4o/V
8kbKHHOdm6VoIDkFntPVBC0OJpkMJJ7lLrXpoOb2a9HqBu3YyZ3OLBI6NT12BiI7
TObagCPUquDBN2CS6vH1xpZkEqU6KkVmrDeYE135fd07yp/jqgnBpxlkSWuI0jL0
1oGnCajXPnI0r7z/iupp3i04f+XyC2aZ5KwQsmMLX+S0FCczrjEVkvLq47P+DzCi
QXpo6wdYeaZQvCRgd7MKrZEzxhUpjcROtkKp0tht9Be4h8qWHBUI5oQfpZs3/7CQ
HOEiJ9qkNPBHCwZUquccaDiWr8AE2gKX6SDrNuMcwu7GVmELMnCSzIHfcW6oH0HY
V7Q6plbqCSCtgeDkEu3AmEm2BsAFJqqIUjHgJVhc+e4=
`protect END_PROTECTED
