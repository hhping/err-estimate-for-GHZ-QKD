`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V03qXK9o8WmNDriW/nGfABWIxqdy3LS0ToaXS9CSIoG3yUb4XjvkIFCL6l+7SYNn
rAtcpUKcePUlXfWIwI1lw0JDbbx42hg17oU79IBb1P/lQpgbvHzep7/v58l6VbXa
KOM2Q/tq4y72HutRbU5CGnlkEwM+oAhFq1IlmOc0yD23RV8x6mnTJjIzhN0eSUpy
sklatCiNjEtmbJDQ5Yk3ODIGfUlc79wZxb6uswMS34w7I+AerQGb3iKNLVi+Pwyt
fRPvvQddNPxApSyhbTwk+lQgd3XTsYUJxKFBVoXHY07/KpCLXMUyP2ttU005phk5
q5sBz5G2c/576kuMtr57Q1SEo9V/Y8zd+z2+PTT/VYAnL+cwhUFeTWHqFSqH46vV
fxXLJr92Ze3/FS8WTh9mcvw12KNAp4wQW3Vw10bBWFz0JHIdK1ckjIbOlr4/xwmK
Z2GmvAR/Vkxy3HLA/LjOMaeEKXRAkRO4Aws60Jl3auA59wTSQH4moIs4pff/uVjm
mr6N1NCBnTxDl32ES6BSq7ts5a2Nh9T3JMdGiFkxQpFYGi+T2+oN4LuVp/qVwgo1
ZUhYwKbqvAaeifvZzwTx3Z8iBFZkznHVXlwDVEKKt0yoQ2VVsGkaU+bKDTN5E2/0
81lAlOMYT0IvcCthmhXVhkJt80UBc4qwOCG5yCjANlRDKSAbkKCZz7A1mJXW0lvX
I6W0JdwQn0z97Q18u1S+qPp0crAkFtr1t4PC06TNXnulDx9zNs/P1RiRDG1FoJbP
3Ul11LEq8akUtisxMHLEjOB8zWTmlSJ/nl2aY2n+EHlUh7dU4C0bfwnEoUs9Y+5c
UQEDFgcODsXZy8DT13QmAWWvOZpE9lTqbvKII6Ri9AmdjiGNyYX7W3CT+7RfLikU
R1wxCIL8K32dazxXTVqqmCVRX4BcEQ1aJdrYo74nzDw9WKo1/IH8bsfklC03NgfY
1vfzEeraAIArC6c2SX+Of2EBlTLGn/LisgX0N/XCcRnzU80khq0DS1UbkHBoMsgO
xaXSnadtsyKwqvxFD3O4cDG9bljAdHxWNSzErpp4wVGGCBiqu7dhq/1ARQtNhGOQ
FsVUjwQdo0llsnQ8DIUdqzUz54/yiC7gGcFfgZk7AwCL021E4W7P++z0iNnQoM6B
MpU9Q8V6W3907ZDXvj/TCPZyVSXefknT2Wc+wEfGUC1x79PbKiCnfx7z8tR0JrJJ
tmdYIOBbz4HjAqx5RGWIFowlzlRKNgGlhRySp97gYd9q6GmDOeiw75WZ61vj2+0I
Te39R0TMUCBEMS5U9/bWPugZTpjAPgLZvp/+nfSPUJaxoXW1AOn8daxH14XTPuNa
8kw4G2gxlhjSgZuHIVqqnJQQtjdtBMBIYFZ4g3QFAud4iBeY7shG5EzbX1PROl4f
IXbM0FvkVODjvGi2gegkeL3WHKkXItCa+rPeTZxnrK/HjvSv9rzGSLUIwsN4dA+2
`protect END_PROTECTED
