`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gi3RauVVGoBVKn9Jrkmcv6BVnFHA21m1AhG46id4acZjvpVnpCGEWK04XDA8AcV5
4YnvLPwOKxw9+yVupvU3iF+3pj+dap73igNtBzXN5oBKElRD3vinuQaoFTWRmkdL
ukg2e02vn6S7SVFxK9mNrecTiW75ZyM1GrEtOrKa8wEszuR9cWnwL2lgkwjo0BJW
l7p6cDJD0dWx+YI03oypTHSiESfJqKXd1QchI1JoYrZ2GJumH8LAB0oQMBCOKf7y
k2xxeXyPBziypeDupOK8NtCqAmbdkhMKbA7LXAjFhxrIV4zFTlnP+UCNYtuOJ0S5
bZ9lZikep87yDxeseAy/WHwx/hRjtFn7JHvon7zfmlOjN+EYluFUMGY0KMPEYl5H
jXImWmzvFBTfGk8mqE7mkeQwP0hHQ/W4lclzrAhuACnIVRA+q1Q00Mr8823jm8wS
c6x4CClaoWpKiO3cyUjiCo0VweQ0vtVjr1nD3slw9cwHW8C9pLk17GE+1U63JDOg
ULhf9wRS5T2yyc8G0ibg56vy6QuNDufrgFgyn9FBM30ZNinxuFEZP5K8LKUvvd41
X7R0EWITgxUA7CoINj7N9t6KV2m8IqB1OSJES7aBfC+mzfhB1AAWwAD7sGs+6E9l
gB55dMVKFkwibcJFk6axfvklt0FAdQBGs3xQ6ZbZcLo5/dNCu5+xRFClv8KpBaG+
kWoEY5ShiqZpFlyqiXnmZojQ0TUzfeDRHVquWKiLqDpaqKctLkDytn64SPR7ZSU2
MO7afnGKSJqE96iEabfXLJQjo5fAQ0gKd6M3Vv1tEpvGnpeFpU4ZURgNIsE/q3re
UQmyeZzYxV/veJcq6jyEqbFSCpoNYgggp/1xmZ1JAuPp3SxPhgun+evTKoAIxEmZ
JdbXp2U2Mpw+kjPxmesPFx6iBGhcOm0sW0nZDl48wwUcI6dmNjpi5aNpQjW7YPUs
xESh1x+SMjNC9q+h4apnsNfTzVQejyMT+OKga96BEPYqchzXYH5Pyk1nTEn1aX/l
LyAAvgVM4uNrbgXE+9d3Dpz5kxVtHibKJWzG+D0/0CLp/qfOJzkBRQzYDS7WPa6m
C64RiRzT75J504LkTP7DrS6l6R9sPkU85BEiNeWW9DHrlpQSFn/RLTiLHDQxGCvG
D98zfqkxlquvWM3s0Cu/1aecMDzjzhCx+ejljRLfuav9HPGTTrd2xuSZV8ILMyvb
TkTmcUScUuQsriIZ5jHp89eI8vt8YMwO1mH93sG3/xNhB4Cel6+arC/JCe/od5ih
uN/J58TJe30wkWX2WG7wm/T2aTe5+FGFzZIyjMLZM0lQMZvbjukAR79BbZ81rwiE
eUtdWCChIG7C24hqpvJi1c9aBApfUXtFLFbM6O9rupcMo+xYo0UAY6b32AgCXnmT
vMw//xgLzLL0i5X5uZH4QmIyv2uFJJKHOU+xdRMGCMdb2XIubL4xUmQ6KERa5KRP
QTeDYD0ewaPp/S4GMQ6972cnqPiv2eCMX+E3TIUGhje8qVdWItac3WDBSi2GA7ZM
va339lsTL+eIq/zg6LgCbezbepuGC5Zz2jv5iB9T0xiZvBBgUMifJDcFEpyTI/w8
dcjz7cSpsvW9Ddt4pREdesoQK+50p74tRVQ2omq4EF0TSRnITol2ikFCQDiZSG53
4oRQ154q6D0UB1jDbhN5G4s5+mFmOf3aR3Emowj5Ry8G5kSVSd6xhYZ8/h6EfsL0
UzQP+7aXypbckXCJCNIzLmAB8f46p7WjQzgLX/IfmiutsZ8aWhD4hRwotcRbVNG1
f7UA2a1efsFEsop5y+CvL5ddphmOTtwAV5qGNVDO/L7Et+RNwmDVR/8T82QaZv2n
AYzG8R/wutlatVaU1MRydu5Sq48JhF8hiQ9PvIdvR0jc3CCUksXahmAnRS5Byvo+
p0wnaemGzcWBEMfaoSIGO0S58Q+sNE1fmRtCwxjgvM2e6fKVDjTgROxN5WAwzL+h
FRTTSgZoAilBafzSl2FJDIdOQUQsaJOIk/6F8hswkQ34AljyUvDdyF/cfZ4hiFHA
LVcIr3NIvvSMMXASxwqeS8ESX2VBi8LVW10Fthi8mfBImF+j+d0RvR0LK2V0Ez/c
BWuhHi9FraaW9XkC0cOqgbttGyX5+hqT/gUIjhZAAANVbtoO33NEgj63wwsrzGXf
+Bhjo6pQhHfYxJy+FjCuY2KmTR46MMXI828bNJCblFJHHpgvszCEW1exc8b9k2Jv
4YMq0gOmhTWkY2/hH36PtDEoTUlJoWC1ekK27iw5TWPH3hEJ6M17vlEEZG7jZSXJ
wYTgugBlFSwcVVK9lHRlAwPlxwGjoBK1QpocBozPgs00/Rv9kZnlk8M7cUFAoD4R
LT9GQ477Cu2YlFjS5Xowz9YEoDd5sHd8c9MUilyidS+mHEiIjY+W3OgRN2fhQtTi
Xmzs2o9yofxcZeelcpG3GAK2/TK807dxZTs57+2ef2gStx1Kl6OVJlGBU66mT8WF
A6kwIuBGmGAv3LvDys8s/+nj0UW3TuMQ1THbqBj7Kt0azza1/C63iN3p84tHwu3i
vGQx2wMZS2gte+r03Pc3pyZyrGe4UMYnbYahdtxOZBj6t0onEq5RYxQ3v0gDTW6X
EtRLniPjb8KFVSBazpzO0bqGlF7eGcCFtvWVaTanqWDRXLAD4XdRXas0iSrpLI2K
pIdQtqWBNfolI/oMckhgFVf1Zij9O8r/IZo5hnsf06FwyfnfZRgy3o9rq45uEyak
bXIWt8aHsdopHHZ4MZRGGjV6SZjrG/Fu5TEs3tlamkptn5zPVu/9mFfgcV/0uaPl
dFb1fM+EWmf5OqQJ9l+wygTr8ZkbfIpJiJS6IV8LCHJgqBS7NOksAAx0tvS62yvB
rI/ZeT8BjylO1et/UC8o7z8PMKfTrBjnQZB+D6BqjiaSqHTh572DzQlu7IWd34L4
UoZBiLKvW9WwOvDbRC9ews3WpKKVLTi4xXBPlEno7+NpZdTqZ5bDAsvXbJVF6FRM
xYoDJNHVtP0EvQNn+kyWFOhuHSul9W2Rbc+9nbh8QGpK8o/EQrjjPtEhjgjznVTb
piF8Bwxw3+FyVMgGR/EV0TkGznZwIOEaV9RKnOdxRayAnWIPaDe1RzLIBoMJ+2DX
fl9j7LptmR2cAvTYynli8vlTg3kiXvbcQSRd/ct3/J0ipneM7cjWuDbh96zYgR+f
2Em7bbli2D0KYjJ64sy+CHGGSMQgDYJCcDpD3KT10QzhzSP2Qx+7vWF5y7Jmlx9S
i4rve8o4yfW2JY5rEuTPDvn3gx4BYIaY++35ODZ7iUkAYMX3scUIzk5orpX7Xone
OgB6fUswh0kjAXA9zS3VwQ5eekKvyIy6fpNWtLKc1lYd1p+vY6bIkPNDmjsespvU
RDO1ktgxXAnCyoJdD6GJhOZhOSzR/D5ytjsdbzj093SWO7tFNteh5UaAD+ukGcro
+bbDWrAoeynHmlaW1iJnmJM0uYcWqPopf0ORfgcMPu6pVvYFzXRtqveSkFgVvXqJ
yyZBYcBmozTHN3lBWD7W8E7CtJWlAvm81hTeTYGfzrzyt9Owz4PSCAyEA7hKE2vb
0Rm0Klo+MJbeLAorVRziRSkKefUkbRT+j0gWywZZoEagHOAqr6KqrCtKU+1zFGdB
04aDFpgO5A9FR1gnOQYc7hjjCMDxEvTgeIJpSEY9uEbLhgXCTcg69071oN+6x4tf
DsYB/WR7RO9SvV2Joqh8K8fZF1lSh8JSSb6+4bbc8JSFXhUYPBB+mdNkn+2FU70h
zdTip9tLxHLBI2iWUcbOFyRm162EddjcibxVB4iEOqOvFyNpdsygeY8bUjuih3j3
DXw+lCcjNl5msiINllTpyc5k1wUWvbGFlsJnqcQr0wJrKkX3ZJeYzX0mL+eo1MH3
iGUZKjvcB5FBsyIrnJ9IdSvpw2Bw8NsULhnE9fuO8UdXv4NLBMYSsKaiHUfulTE0
CNP9zaTIh9iQzzihuG9JSX0DFymWu4jLWmIz8MOcq1YGQHMSFSxtAd/nYHC1O/aM
qcJjOLnCmfvchqL1xN3c+U9Ba4m2rL7puFLubHpUyvcIV6+ZiZkPo9BQK06XxRkb
QHNHWJMooXBZW53bz0eqHiPjRZfCYRUZ88mdZxzq05J1d//DyrWK6Jn3m8Vzn9e0
wPMOVlnrw4kFv1Ny6RBlOtrssfmSB9GKBHMtJTji4kt7Rj6jo6xOnU04EYE+NNdc
L889T0Wd4auJrt3HTICNPPL6NEdhKfDbDXbhH6NiwxA0xTjKDHtg41XILhnchRBl
lyezllgjv61Qw44feG4B/014agrXYC5hTPuCcBWYNBX+WuCKMbHjhbYQ2DbxBBID
hALxV+88LbjPqoVxeJeAIx9IwAemGk2CbAG4JHLEGTAOg4nYaN2ejflh/PxDUMZI
bfV24YnyEKBPRy+Hh7YD8mZ/BG3UCDFvEV6rVrB5dQjW2vSt104wGAlDA1EjxEj0
xlfQcXvNLBKeuE6QK8+s+2Q4f7Smqr6ZR9lssRdB3bXw7oALcOXjYDusStpZ0+s1
fg941d61xU7t39tgDioKNTD6aYWVsF/oZVNJ19hHyAwcPwv9IfmJiBnqwftNCpch
C/8DzROaZ94YwzfLBJdV4KAa1JMQGlZP0XUsXgmQM3MveLMNg7Lbd9mSIY4glzZ2
mX8kkY/D+I9avgok/mwIwt0f+Pf8yIw2wuwXDOKwIj11FtGynbMmNgZef4U8lBfG
54e5REQibmp8mFol/u+hljdLwN8XzMylGGbYTvvDCTqGjbGeuIPGF4dgl/Rjbe+P
kbM3YVVGJA9zUpZ7TABzSMx0lKKsDY4MBCLrK/9zQGlL3xk+zN5eA1rzreW9yp6P
lnixS+UwUn5mjnCBM7W47ObL4ILCzuEgfOHVz4Guy12vnmRgORUy8zlib4ZzIUGF
bzljDmcuho8Fl03D7A8Scdy6WKWDtp1SVs6u21nDtCoQDhfrWUHGKJTn7376ffc3
cV7tNtsla2NNjuJhoOvsZWqFS2Xi4zuiXrLr2qB1aAbFXhfa1cKEnI3D/PjBJHR0
ZIaWiUXekAjVW/NpFtH+JBXSlcHm+hUEplf8G509KhnnLBSPy2A3G6ARViU72/Q9
lD3lxU4gtMGyNfBfz86RV/f484FG+J1zNnSxx8Uk81A+82Q4yZo7a9Vz0rOnk/Nx
W1JnkLJmTTx/DjjO/6TRsu+HEp7QFFQ6sICdmFb83IO/ol7jGtAmt4Ngi0RN5rnC
HeXt3NuITnc7coeIbRVDxJdjHVhxY7WeKdnsX5SKAp/2BPlhfZTH4HmLnS6prPsN
OdAPziMTtHCOBY09e+ZPInkH8jV+jZqqlWn50cIqVFZmHQX3FHM76HTZsqh+OUyX
ex4h0v7Vp/4QHCT8AU0CaeJTVRTBykzKxTAuqC3NRkDgw6UHSPUBFuhZFBH08nNe
BeRyAz5Al1wzw/LYG3UG2SmqTg+s+A8DVIe0KKK1YpkQryZys8FMWsSAW+ur6Xdd
vLwa9Vwm/klzzDQdmK6zR9ReVwNvo5NBaJ9YphzAGcGgAF2DmDOoph35r15QEaGE
bGgOx5Jftfk0ksslye4ajcCly6oKhc3TNd/2maodF9XCIZx2Tvknnic+VwgsQlDz
JLvZd374b2J50zAGfOa7MyVp6IwnUfkwqfTbh9BpSsWkHRF3ZMj+x2UkNPFuYa8o
Sh70ygaLJqD9oe50fOmVsixYSz3VbfPiQxaJHE/m2atgWZ19VK3iiU/mXrJsN5jm
aDNj8hr08rKbw0XA7nFLfzIzQBu1VEdkHBttsw2Ap7q8mwNoW/LicB+aBWDIjv7M
ND8n3hMZvMQjKR6e1YTScvBTotTCA12vV9+M0TX250zAmZKDXoPKzL5pztS6B6xS
7BkTdWHIZiFVjdOVzi0ANtmz9zbJC/jgr+dtIG+bYehB/v0WpZ2qNoVYcNjBDiHs
kJ7iSEs0PLJDc49EyQPuK5HMSmLl2rLBmn7dXf75bIohbSAvW7vyfl9a1EZRgRV+
Qjj/rFQIhDqlg0oPkcMPqsgYvZy3QLM4Qx772zM4SidSZAato0ViJYofS0I+Uqbp
Q6XMtku1HnM5uiprGzzIpw1ppUmEzIdop980FU37raqnUV+bPvFspkSPooU+gi9c
vEdiLTKRKGooyzh19G/n1CWoflIMPu1kipwPtsGdXdaTm+peBOQGExlpSeWBTS3T
97reqpvb5gNn00BKrhND6Nt6vDQOzq9VMmENYiqeomccEdz+7Nlad4p3teUugEgE
hXq1YKETH6yOiH6iWVs8uf1oH7oAF5zda0crZrM8/NYfTjFqC3tIEWxXGdeGQN03
bC/BkZh9Om/liMHZ729Ii5JUf9J1C8+Xg2Ks0So+CFhc27uAU3bHIvukFj0vavsQ
Z66YcZ4Brf1aD7KQ0TNS3kzSHEdM2DfHoYsIdcsEUJ87f+0hn9xERxNtW47xSPGq
9ZFL6NidV8C8917uIe20OPhAyBc9JGemsA56SwCxK9fLsa+eVQq/QQplPotswdu7
VXfxL8p7IbJbhPBv1n4dDU/o9he3LcmB2yaP2S8Ghzjht/0WcN48gMhQ6cxZWHJy
g5MPk+J8XRH1mjw7hKO7sy9X+o0PXtXZaybcsu6IgA+nZZ7I0RY78cQxptyXIvVq
2SNzZJvuHP6rimEQK6rA3LSKuMdcGRvlwtkk4csQjcOfmJL+5xNG4XuhaUQ25EHb
6Mc+2IdGwL5iukytsu4EeXG4DnTK2F0N7yyezr7kQzodFtimIS+pLUkFNLUNV6B5
zKnADJA5aOpdNZ2DqFleZ2NJZ+WQ4qp8CIuZf16QX5xuKrbHs2A2K1ypQr0p5JxP
/QdlsJ5fe1UFhT2oMPD76Lvaoah7rD043wFeTw91TkgFKq0D1I4hZD2QczvYXRSs
NxFuAJQgFmq08XEIMe/ATZjLdZc2D3KOhgs1E9yttv7d+xZX3CBMOAXsHlsXhloZ
HcZUnVOajjxeDSA7rO39whgz+3ckbjN9rluMsZywBVmcUPBvcRHq1jHvwexeMyAu
BFSPZQL7XEBFvTtfc0i9sfgUraF30SDCYB94Lnf5vRC/nIBcQ2/8yFe1ox5mlzgn
+u0MpeErdobAIwuiDxFT9FIpT1nN2SJS3oyTa+UMYDOREAP1dxlHU9v/bGSgBK/a
k/gVGarK/+levIlIIaVmXBJkNXFdxlijJ6GTQX5ZKNggXod36pR9Y3S/PVq36DsR
O8N7NqYkQ0YAKgjVMEr+dAGpGPUrw5k5R+4qNdYfdiWnbVdbSL9vPStgAX8otBli
bM44ZsUpvZ0g9GRru2H4tzepgEy1/xtzISqY4Ezk742TB4nb0Ou9sgxuk0z0E3Jx
m47refQFrpLfysGOJAohXjGQs5qh0GFKvBdfkrHyo0ICars5CN40/N6pKQXv29yz
m6T40aaVWr+tgRMLWZrXyp0sGRXJSWyLVS29Ayh34tzPwSCSmAQ35of2N2IrcwgY
16ENcl0jo4R6j1IUZkKDJ/2xxxlatVeLC6s+Mei3SeFwR4EjSfmiuonb9u5cfaBN
RJIIdAsJw+eJcvXVFc+qKmFJEbpmb8i8z/UVOm3fnFy04gIZB66oa4Iwinz6dgZA
7c/J+vjFb9eeclvW5aKnilAiTCGzT2BRz2nrqSNWH/1fYynSzrXxTf0gV527+xMd
qfPWfZPdh+tSME8VWKmh2MTQjKkqoA15SkLF20ye5azWY5Q6OoSbi1OdTSqJ03nv
OYDcC6ooshqBr0eNI7OloydK5rm0aRyqlgR3cwLO1NfDltX0fRsSB3d9a0RjhN9i
6ZhYA/xqjfGBkCrUy1AyNjDtxzNRn6pyMpq1Yj8NZZ3OkfVBl7jnbdsL9RbpOK/k
T5hdajNJOHaZkHh7Ki3NEcOqgmSUhrkq3QdZtzwMGLcmap1kV1xhbQf019SU6hZK
OREW50JOvscXmO1USZzf8ppCFm+m3g6z8eDPEuAsyvqnPFkiVXV+I8zsMTYQH8nr
9IOx7+36yghfMpCOUvLS2jctqm+qwq0uSBMZo+WRw/nMRO86Vn+vAKiKrdu4dW2h
XQUVc/2RRgLNVkX684M23Qu3Sn0Gu68nE5rU83e+KNqxedhJ4RzqeSdl5nHA8gwH
nue44DSiyH992A2xQi5Ohm3GLHYDzaKV6ZpfSsDQh30pvsE3XGa+4ezvpHdaJ0n1
13cABEktMUGjuGd0cVDmrIK4LoobvN4zLAspDVJIUX7uAxC8hl9pMUEXwyMAAoSa
tvaO2FttwqePJWk6up9BBRpPDJZxQutZu5mFs2e/qQbjeJETkIps8b1mjO/QW9js
kAjDS+y+sZZX0Ef8vXlJvA0NtbrTTvnXjJZZXhRvk7UVHT6174uR3EvDeXVgJHRW
nzKy38NbRFRZasLdQGlAYimF0wHBP0KUlLUWiom3OB1Vw/CHZwNcr2gU01vj7L0m
t7LTcP7sQhDGgwPc9PDCzVaoUsd5MK51ggcswDEwTXfc4xHdLkoIlraJO0Hu27UX
TAK2CMHjjw+o5D1tJimr9qOwl5bmzo7HtqdvrCZMnxt4dmHsMXlA9Sr0HZUFwH2u
HdAvFgh+d7WceKIeSN7kqwlQRmpp05AlsXgHoVy4aa1cCReZrdUBOqzsMFQxEfY+
jxPLQpg4OnOu/xpNKf7ptRUVQ1iaIdaOEGJzQs8sumTjKO64c2jqs+n5PSRqycU6
F69D84EUd5qa3l1De6Zp+Acyshyh85VxBgTvtj3R5iDQPwVqilSRuTtuUbV1jhao
SfnL2okCaXwZVtIghyps3tUl1AIJJcOe6QbfYjr5Y7QhEcY5uE13KFfpYdjQ4DJy
f8saYI2gEK4AjqZdhoZBCv9ayrT7Um7kyJuR5vvRNS3eBe46vssxzphPGolFSeHx
i/ANjZVwqPvYP2t1eJdFkgKqCR4VrbC1zWBeDk8o1JU84O5CrmAqlnNt9mRRPYzq
UFdQdT45+z4l8CkUr0rIc9eLdD0aty1oNlDOvCkIyAq3tUtzuXjjAdvG9avg2mLD
WBVOBKXvWQk0VcNzBgVoQF55PdZzDzMWrCgQuRq/6XDVn4OCrmWazqSx6zlb98G0
8zXKd6toLYyQSfgjkT+CAnOA8meO7QfwxKX3f+0XWTbe6se3WiRF0argFB+bXSfN
oiETHaPg2EQlXaNChdoGp7jsDdewATUAlrljVo1grOKoAoJHUz91fenqwSX4JjrP
hE13gjQAupm3G/8muBiCs6q1JbHfGzRBltMS9xcmmZRyq4GBnLbU9LMAommkGvKz
7KDfXQH9fg3G8guCSHzLb+ugAsCoek4bYa2eUONhJux39UwxHYnq3rz5K/8/nqMf
Ef550YPtSON9MTrAxGsjH/Rcr0H6t5OhTdyNoFQ534m9KSPGVCO8injBHheYSC73
wnNdOPQhOrAgm1wfZEeqIABqqrMs8tMrBra3OUutLT3UD5Hl7klZiWTdRsICemBm
H2739ioF0BAT9GMqPc8IHiJKhAwn4VBEZ1SBsgA9/o/727QaZLbBDIGnuLG/DFML
SzznxLfKsYWXMbDdmJOvVWGg0UklZL3PLg86dtA9lRzhIu3y2MLeXvrsKYKavOHu
cvJ95tIHOE6tT79Si3Xpv4CPBNvZcu3dFS2306fpJA0WRryxZSH4uir0T6YLyrj1
6kHC71m+rCLgBANkn8p9VwTN6gWG9G42tnwmo6AkAIvz4CL+OPLv3Xl0uRBUpHNk
aQcNhy6tqBtXH+h2/NWvdRtkgu0Kf18/BeTEnfp/C8uzEBy0Ya5dw/yeq96B6Zah
84iHjGReYMdGOIwr3LEnrI2W5nsbF1yzvjKaM91HWPeighmFm7YLMEoRnoCbGywh
j3zK55X8yjqt2ZgKecmuEOE2wFQijmTK4U+yPcImf3p0+gJbQbrSYRB8ZdPZ/N1t
hZmUGrQbAglZcwhY0zkhEq/g3YIzcFmuTOCiN9jyYIZ12jrV9jtaqK7doA9vUhJd
zmfBzvnleQAogsxmFo1HN494rkrv4w9UmwsFWKp3Zctggnmfcwl8FRt6TlP8u5Nz
sz9KjLNvHiW8SWrJfLHsHaqH3DvD6jkT4svulGkS2esao/Zp7GpkHSoXTr9tkIYU
TpgoA7CgrJPtxPklwUuSrVW+e2pV734euo+TQ87XbtqomN32d2uDKZWc2UMjCOxp
xw3l218W0gOpzJLU0p7k+f1gPK6PM7WHaSyBtHoHM6qeQjAc9pXAYXnSlLlqa4eR
acbcldJd4cqfBjv3QFwrGiLgBsUDPSmMTsse8sPqJSlSy4+rAnBddHikR8XdJoVs
cgTtLnyGPTb03XPOF+j7AkM15tmSoqwaDyqarItiqysbA2AxKVouxsTQBgSc/pgl
XzKn/LuXOk7uJFqY2SS11Mmx1iGR2OiV2MCxXmJvjqfEEX6Dg/EYw5V6igSTQQE6
sTvjUMWgGLg+q8wvRKckMHVJO0kUyvwQyozzc4eGAQmw8c7oDmSLwXkjrjv1qPeg
UZDJX6PcKSWWAFl4DCVSvy7lU/wUK5grIJQW8Qtm/PDFgWMhK2/LDYxmfpw51G1q
b0kRAp+bpZVhC06dutp5cy8WX+NPAQD1YuLIpOXwaNRH4itm6ji68p0xa7WzIb4v
O7OYpemUMQrs6hF7PGGeCMw8mt64Yejib0RxH7K0SchlcAKrzOEmL9HzAnHTZlFP
fYh55KodYPU+ZK193yS0ygWNShM3uJT9ftCuCIofmQIP/IjcEyI0HqdMVW1jZCsI
PZ14jkoWRulEbPTUGdMWGjxFVdoVxOlgADJ/9mNXa9EvzTjr2tOB9qb6RI3DHcGh
695Tqk/HznPenEhnHtVWWFCgjO/JnqPzXedNIJ9gvYK/mhkOfazLYZ8SkzhdhRrX
r+LQypeyTj5F3B0sUmSk3O8ZKKgpkPrOjKjB/lcJ0TI14OX3UbP98vUa6K8ir0Gm
xbTaXlW7M3BzAQN83pm6fqZsL9ICGopSa3JQcy4f72sau1PF+i6cmOk3ySpGph5P
ers7ANvW4UItFvaW4in/pumrdWZPnrstwvUbCssm1ZX/gpMq88RtuSjrKaZh/Vr9
siq7AIrebvI5zNXl0B6jcNnAg3/wmapu8ScbY2BNJU0/9uGsakp8Urgn1FkrlfZZ
rr6ACfQnisWkP4IOJD3Ls26HwK1Jhud/QFEUFTmYOLADcPaszNaxYhwc4KXLVypA
LqzFNpueHa9lZmvyIyPc/qsaMmMy2hSBz2H9m6Hu5lBgeaDH93PT3OQG3wWleKYx
fhzC0t8iWNZZQGqTbakqpIWEtV/C5IY8L0x6tgE99IyTLRiGzUPUYgy0oOA9wz9Y
GzE2qAymIidQnRZlQgKhBf4ONY+VWC36wo80aH4uf9IdmqaT5QJfgBRRCunYvsyV
QGo5FBt518P/pshP+7VW7UOemPI6fSoXs58T9pE10Vrim4m2dNo5ceuvwCojs7Rv
Vwi3KLyWWmTVZ5sQx9svfHj0rl48qC5+WcCy2UGUNqzKVxDlROjRq+oaxew4x4+n
OkGE3cPdh/O+CGK2aCga3SUo6PWLiklCs4Uj1iAc4914bRS8Nh1v//PLmcvctHFn
9YuGD9CHSJod4TA4KTpxGnt7unSmmkYPXM80QxwAzF72Vl96UUMIP36eSozL5KJ+
K4yvr5GjCmimChm6HBIUgfGQWJISi4wH3qd2UfdZ6RnWZ9M24iDnHGx83/qd+FYp
RAP/sfspYn3eC6yKhW3OW8X8Gc/8PXi3QzaX4mgEN6Aq4Ob8CnkPTxqsU1ZpfhGV
xHPCIMYLOML+TwRZlrkGWr9/jc59zb7ce960xOb9ToWkB7bCTfCiynEyt9N1Tco0
uAoyiVC559484rWiHUiP8C0LoRInfaG9HpBRFN9w9aSSrTM/W+xoX+XE7Osdz6Z9
14kTVZCehLoLRK6zb2Lh2Y9UsGa4r1SGQdYgutiZwy6BbPkGdE4KxU1D5Qr6k71N
RIecvDKvfj6QTWE8UE8M54752xKs//H7s+R/oxA3ufxluOz34eD4SgK9Kva5mwjT
pTZa4xju+EKgbBqsb7hrFlxWWQPpnOWEi0In127qqPB4/lcceFw32Oc+QOZRjM5U
WMmissC5bjK6sMH3esprxHNq2Jy9OxDvxRIrkIUCJIqrLSz4BhGcJE7TtPJnTcS7
/9frJUz7Cmg4bx2ZKZham9++aQOTzjQKveZiL+zh43itXkWvwnZXkK+sydyGJNbF
v8xd9gyijzdAqp54V+fFwJhGhqSGiwb/mvdZszJczdFLkEeLCfXocWqnhWUgzNND
8M8klsbgmFv68mMj/upOuoseTi86kxgr1KjhGMPg+rn5wNLr37xWgSFzJdkPl+nS
QXVMI3v1uleTesUP/9eeLhtupGwHJ+8tAQuI0wcxpM+XThon6BiX1BRCmRnRsH4m
p71BWomhTR2bwEJ+DD2mb4bIALDaeX+L4qi9vNxUKLtOXAIV5/h1XLqYbn5jjeo+
CUj063hy+JrKaJ0G20BFw/Au0stuF4Ql01L6WsH47zbAMSs55OchW37yHpLijqjI
uuGv6wZwAjAxn+XpppGa3ScIqQtrPgZmGXTQbWkMPDI9c0Lq64JiQOGiKbPYxEJ1
kvqJpsB5AUpEEE7asF46oAFCwzeiR0HqA6sTQ94HeyiW4RbE90nym0FDPwa92wt6
wqND8zYrnAYXe6Prl/XNkBfBtjslctE/Hxc5x07rdv7G9oIKowrBxTkD+nFZPCM4
ZyVXUXkKGcerY2R6JuGEcRL1T6Crd9QcpdZYiqZLXyFlg4loYgo/+3Tb0SEEaDB2
yUj1f078MpkeISCuz2hQWSf7xppzf7W216a7Zf6lfN3ueGOiThxPSaJFejXaRNsu
ubK3oCJDMpd5TZ0cuBKYY44em/WvlAsi/I7KnGJJW0Qa+G47HSF6mXJtuGDhqxZb
xYVmCvr5HtEQlU1gQyPq2klZvCU+J5siaT+HUPcduxy/IzIVvH763rkJ+nmvQKo8
S8F3eRlZ+IBxsTSPynD0KQX2DS1QcR5b0RCjd6t9QlvYd6C0uyv/jXin3jhhHYWk
EuZh/vg/GHTwwTy69H4iwmnMQ1rzb9ZUVgouqpeg1VIL6lEnSLH+v1zbCY3wJy+a
dfWbLfQMw5L+ME8KcTa8bph0BTXxWnJ7XtDhgAy+uOfqtNq+gDawo6eoWp0MWNCP
UAQzBq0/bVXh0EmLuJmoLx4vk6N/RSaWlqHtl6axiiZ3XH1hjORWGpmz0+mUrHqz
OQMIlKV0qhWOswyaGvQCRNtzW2IVUg0tZd2WoUZfjKLnzB9aFTZgNBZaR0vb8nlz
F15E36WulOaDURaK+rY+HDHZn8dmDiPQxdQhvN7ehlihjSSgdLHimhJp4O+a8/EM
rg+QLvBIT89ggykGNoYQQv0HRoZh6nO2Y0onhh/iQkSZQm/dZbBWUIOuXZLWcPnQ
lSIWam73YHBvGmNNGXgT5Tz33KDl5ckrz9bKEDghApKq+5t/TleVK+6rg0aff4Df
6E7lPWTvoWE9WpeJhIHO8U9OEqklDwzeodS8a4dPAdBVmvJj3cxVAvyG6yEQeC9T
mExXlUZqp0BWCEqN5Y9Nn1/v+k9QrCj2/mvHZgkko+Ou7HxsNBv4tfILI+M5OBhs
/hR4oSX0l1qpqDyKaxQoWQpj7aRijG8t56/LuHAelIFgSPxvxZcf3IiRsnHHsO1T
4FuQTXUAapXyHxCW7suECCN889/m/BlA1ukO4+OLNWOfjHSX5HaTLeH5zy3e4rgm
q/ovohjmrQh+bwe0+VCeyARBKnSrnJ1uKbt+YUp89SqgH6b2NmtJTm0bB4chcFfa
7DLxsng+y5A2GuaN0JOiqOrEz9AfpQIXFX9hjRnD3vaNiHQu7s8l1SkXI92ywthd
cANRkX4Itfk0+2ju/zhqoa/0HdkWLsGbnjhYO2bovDpOl8O+/xciVZMvhP08RIfM
UtX1myjALgoFhWVU4xN3LzZVMAu1mNcfQ7nDbvYniLFCKX1P1B6TEAhlchbWoyUJ
yc2cCRCEkeNg9DsXrLP5IrrwGREBrvBgHqM2lbljDg3R71eZ+EE0ZzzEssJ6JZs6
BGML+3/9bMsybhm+eoFAi9mTMl1Udo3GIuHx6ALHLN8YMpX8KOuNIpHj1Vcw+Fde
bBzgFhF2TwAFDzAJltF4L4fve11tg3Q+oiVOesPu811uu69BCNqK7a4seJUaWwnc
wA9MOzDjCkL5CfalgFPs2cf8fXckxditCDjWBTWvK0jf7um/voOrLa+0nUWM5Wic
ghliZanZm7xYd7WJkquHrrKpyJ0KS+Pn+3nG1otNzc+dxzB/12qdN/g0L7bUvvIc
dACwYl7uYt+RbUWeY1flsrIPmrVSMEMpuROWVNHKVnPf0/X0DV2plgZqtNppA02V
VjLaTIU1NJ0FJWpU546F59xUoRjtylnwdOQ/8n7QythWErBamcYso9nG6QiTbgna
s4/NhWZo7gi+1DaaDmdPmtXj131Apqm0vShE9F4Tx1KC0XO/g4hewz3pV/Vp9JTO
nRwD1M7+zqedXJPC1jcUNLCiqlv9RT9WS+bhxk5W8YH5ZUacLJgMRyBawpSQ9Qfv
kwuLvMz48FeuWFdwjPbpkOinMX9BrTMNpZfyXSgBR2oZYV30dHIgckX53JGG8rx8
qmhnkqPtgC1UGi3zs9GOxeCeyfpQCZxk8hktGZ5aJxFi5vbB4j0IpZ12Nmy2L9kN
z85Ya9h5AblKEu5HvvG5p+x4NGMPgOGpAPWEy3aPZ6+Zo/mI4OlpHGsLzDM+08+e
17+ZOgC/Xnv8pZlzwyKl01kNkqWD090fdEpzteR6nkcZMSlhLrFBHzrgQgLhgALS
+fdc1eRj47ROwasq65EDIztFTtnbUYAM5+FeiXTPjnq8xFfXBheTzJjka4L258LS
bExmtIfona3iX5mso9h75QbeNOuNslxienyrORDeARhLQBzwuYpM5631IlX5sOMn
pVkKVNX8YT4hyaU5swZpWR1OntDGdiUSzCRx8Lg0rO4ghOCnzDVcSb/HcPk+CSjx
3FXp0K4K1MbtFccSLVoG6SoI83x2guzwkYt7eg4TeDP+XQYe2gyplPBiZwMVXP4S
Vb+jjJCV4Ggb98MOCXgifiZ/y+VzeUkaxUp/Rd1cwL0Xif4m8PnD3cARTxcFQoBS
QOIztaeCKZv43a8jHewbAmOdIZ/fxwTC/KO4Bv9riVbG3mWukQCp4q9k3+2jyZb+
J3wBpTUucc8dKC4o1N6H/tWeUuShi1qkq6M0FUEzxx17PhGU5D+ZcIM3umOmQ/cA
xcxBmGfHtaiuw1w1QGi6vT0iY5OXMl0/uB0igpwl/EhWQIwIDh6LDH5tCN2Be7Tv
rAiSGX9Yn6VZOzioGonQYiOx/5ERut4BLlE6bgjaDWXd3vL7qua21f8LnjumXq4x
17bndEZSYHy2ibDP9cliiYsoRPp7Du5x1DIlTl6TAwx+PaflmfBc1bv+zu2H5eZx
tkeOwxWWtmxCZLOLt8PN0b65HDBadpWAKPorvO+IK3pTAbeCHtAheo1hJAfiOZRM
hvQZgBm9dPeqUqQsQmaYRFKwVf14uLEvq8LyW0q9hUpGfba4JjVZj+Vd8ZfKD+m3
H80JvjTMBlcdabzUlk5ZKB5GVP6UMztSGSBAMLJL1ZHf5b45K2Jn2BZ7BFabULaO
zqPB2l7xCYaPzxyUiADb4twx9zEHGSEFvPUGd8RRMHYQHoYKvM21YbjXPIaT+cE3
BuyZR9GqyvwbQxe6jxRk8kPr5JJ9Txk603Ef9xBP8XZYPVCHLvfhLbH49bNkUiUh
V91jgJTvo4f2QdVdCKg7aMFOPqjsUz/3o7BVRfj9bUbXNL0fbXry5KCwo6g8BFmt
9BHVwc11oFlsNVx186u/WvxGT34djCs0VUjjK9l/kgcY70uDTgBIc+igZT4yZbhI
JucKXXKtlm9pbceNp7I47l5QfkFchqjQ7kSzafD3iRUjDTHVGyzxE/swGXTlS4Af
zzG+o6QXQCgeZwhiBgmbLED/aJ7Fbidc7VZ30CRarEIffEaDMwY+Hw0taiJhv7xr
n+oU4y4y02afI9hT970bf5n7KBiDb4aogx8FlszRimZnuYtc5tLo17OsrDaZISYU
u4uL7wYwBTej0xRSuBdfq7v+Qu9wfsPJqHDfuyNq4RipiGLRx7CZetCLvQnp6xQ7
ubVcHuQqahG3VspjH4l1Gc9/g442JWCh2X4mQTRv0IShyM3mqUor0vsi+GpsdT+e
cozk82wmlmaclq7HphBJ6k84FpKL6pAsU27G8Y8T+chSIylqctfenCQouW2GD6Nc
Rbgq7Ymo9XiY2Hcpupwroe2/LFSjnSe0kO1BJHedXtoR6lhqQvibTwvnLruW5AuF
GOtBlEIBO/rs0fsPEiTjwHLwnQ/n1cdrX+uib3Nm/5q8ePMA5k7fXJMlfwAgA83Q
3nRFoRAHzVgQ2e//BtxQUxRMvMSjH1zKZ9N7qf/yi2rm6TGwldt9Nx08aXkO0tKu
9Rb8Pd6GeP5inVq02PxiTpAzc7aXrecWyVRZCcBvqKyq9WaZmhCOYNoVnj4QF8Gf
RKQweXWph/562Eezz+ktRZ1WwL0XiXpbgp/movLPSGEQmLDQcQnda6qcJRYpBlBD
DIAiOnqGvj7cLNmOgiBPDaSMsi8g49ZXGkBzMeu8rk8H6FPdbiH76iqvZxTUByuK
FlXvkjSn1+vnUipSqz3jqtMxLQ78vM+FydvSuVCB1yfzh5MYQ2+3eQdG/wJ5h5ac
4Y3Bdj5aXPV4hR1+KbLT7s9qqlPqmslh2OfmUhuQSMAXyapmHa7YSr5pSTOOjfIU
OWWglzbnh89yy2rhMZ7Z+PaI8JOV1Ypb5G6F/XiD4B6XcjLBJCZnNEQuFQEciAD1
HGLXps0UWMwOpFnM252fi7mM98VO5REbOYY8utl8Yp+rCUtEsIsQUn+hUh1MKise
E5TZkiynhhWe2U/r9LlHyXrUIdnFMyZYpgcw+WgaUOrD8QRFfI4GgGUoKVt+b7F1
ChQU9Qi2hvw4/bZ2/Zr9cfEirW74SI8C4GLwjGS1AOmRNju0QnpTtBVTxuTN55us
PwrAXTOo4+aIhkomGQYf6cQEUVZyll/bPtzmYBSikaDY96RxUkFLUkUsHGxauvql
DNHMOs359TkgI8FdyUfjqQctX1wq7tGHyVsAlBsTWrDHqmAmi/qeVBXqPUGfyCU3
eDtM0j7JSkZVKPMwjf/hAl8mP7VfulDyL8Ofp57YI49yTBGdXMheGky5WDCO8BPm
F81tMrX/WAuV8XQcPYiJtlGuSnaylcmx8+Rjm53QOeCIze5WG6vsFQt/+gdydn3q
7PsbWYIWiZFyspzIjaewM1GkIII+n299Co7Ay9Zz67oVqP28WPthoOOR0iO8e8EX
fMwZrwBjo2u91CsBmNbABwxqhs+L5MmhEX2yzFEmVGyW7qfW8PaN/kiPQWKF7iBn
4g9GlBQixqZCvzyckKZ6ossExaKU2pSzdYqi0lMx6NR+JiGpKXjNV+UFIZGsut/L
Q9pReUfw3wHYhD0M55znLgtKVTw+PtLc4eychD5rXxQ8NEDY5S/T82JjEc/1STce
NNuIYV9S+lY3jGlq+HwLi2TYtO+Pe8D5xNdRtTRS9STF1gxTIIY+w4ukArZKXDcm
uRdLg7f5I25bBeoensPqk61W295UhyID+bM+w1xzMUjVAm6AQTUzdqNrwcNUtd9+
24nEiDFRJBSgILbGvJS2sy3fMgVuLDQNA+GnJEQ7qPXqYtH43HxjcURuIxYmOT6j
FRkjWxMfn79JuwihIpFkQJCvUH3GE4Sq2dqkm3tcK+qlX9vqaMICvALs0mpgIgcJ
Uj8/SD5qgJA7TKGzeeZxovvNzxNeQt5zWH9mayv1skg7sJgNApBZaAh8arw+hlwy
ROIfaNxuEP4OeWOytovCeA7blbc4YTA1JW1DlA1ctYEIHMKN/tpV50bDcZWt41LX
bCI/XhfL9BBXx0/j8/T+P4drUufIJNEgrlnY7z08NCy53dNuSRzcNQkKl+AUNOEu
Y3AxSaYHaXjq3uiNywezuaKUx8jj7zk+jIe4RManSkscHpd2Fr9eSMNEZxMDkZu7
VJrgyZunl0QFYl+bDSOzaRVUlF+ejZTRW0PO0+lS5fgQaO5rxsDhVr1icmNQtq/r
GlPD1us4uMUDHm+Rlyfq0qTwykxIPRBAMBHX3Z+pjcYH24szPZaYO69XA4JW61oi
yHH16EnO8Xqapo50FGZS8/e19OAaAsLnNSlOHPw9eIQF37/ZjkHXnrUb2vC3JM6G
Ep0XPKBFBbRfrc+kK79UNM8OYF0YI7r18ZN5LR+fPU2igvaoo4dKIqYElFk43NsH
HsR/5IakCroCW2F6H8EMClgI7HayKv9x9qlqMS61HDiBz8J9Fp1qxU4Omug2DHbv
Wnt16Sh1VywePpkX0XmdKa96BMqqiguOkoGxYs+dFBaygqFlbb3XYk4NgKTfKIJo
F+k4jGl4xdqfrYWk+6qCDG/LWTOPjO/87TaO9TbCZ7IE8f77wqkQJd2eEx+UDnwP
53l3L5998nH/l3kXTIFGAbzj5w2gktfeitAJmtdNIiB8ktbGnhHypIju+UU0rr/C
GSAQvxfrZ87or0PcbOMnVoEUi9XXrKW3bJ2yexAsVJarTLGRRncbJMumkWlPVXf2
z6dAlCspdWroNpIbc8xihQOxxdfllSHGPGZ9DgLnyFm6nxLCNCGpfxfGorKb1e7v
p1jgKFKVN2gmk8vH9nL7oKPHOvN5cKu2yP5C4lrH/HDYGQx6ea1DwWsK/COrUEx2
HOyblMPLzh0UZbDooF12zezd3QmbfJ84vswrMtlX92VD/7+rKdjCDtZThR73fdP4
AkGRdM4D8QHTzzzAzXxCcUT/2IRWQdUXi+sH7306GePYVcMcNcfhx7x5v+trIYEp
BnckiJ2zjbb/wgG2JPqXXsI0PdoxebT87PIdN+EuG0IOwl9iBfn/ytaMjJSAK7Zw
BXOd79YxpXU5aj2295IIr5PCIBZItbLibsKfM4//Jmae+ly87YrQ4/zuuNU75jNM
hSYtmMgWczJi/ciDtyqJKy0Lm2gdMJpQMAOBQmkc2/bMUAhu1G5VbHXqALQ5rWOw
sf5U84sKd5IPrMIojJp9zC3YmTjPynrI4799JF9FxGomjz0Pe3aHrTjOCTB1lMxh
K5O3Zn4LKJdUM6jDh/QjOKM5alU91KVJhMUuvdkk3R7oTE1m4mYONjHs5LYdwjtx
FDkznlZTw+makP53ZpGR/X+wb5aRqZ3TTU7GswSDM56TTdNrKoFSapX+YEXjUDxR
lmqh+dOL+fSxrLRj/OvCsodsndlJccGI/bpO6L5B328/9/xEnbxY8ySHKvtHA7f+
zxEZon36xuL4K69MS+eISSwmOUvyFmZW+H+OMdCUmuMGvB5mb58ISXNnCNCYvb0w
JhHYUg9id1n3CeJaq2A9Aw9xyExgwH374E4Kzk0E9NUw/5zH7NYRgSiP5duRBcSk
3zhGaLQDRtF+8oD2VuCrPt/W5sYwFjglPVIWU7UgINtCqjZvnFMsKvw8zdfTi6lj
cEOiHGFk/8qeJ0ZVCJnYQHTyhl2hjc/l+2LD3VUBZEiSbA5I7gO3Q9zkVZZ8RuJM
r+4pUGLWf2YeMHH12RD3Y8ZDO4KIDLINpJ3X+1rqxR2qa6+5HcElowgGdjX60+Dq
wlBI6s6IEsdBcJ/7xKshpohH/imJ7FvRRZlpUpSZBbp7OM82J+p67D89yvprYcEJ
usyI4LpG+lkz+Ay3TOx3uo0L9gJgaBV2SQW2WG7ik/kfoR604EIGzNCkF8gEeKtm
RM8GaYqZK6Fk2zwL/1j9QVa5UvMatRD7L5OOb38x7XVONxdklBC0uNFt7OVnpnOL
G/NbIUW79HwnPFvSpiiqjqfNAmsyHis3nzQ8f0Vgl43JZ7Ue969ZDjtMEfv5qFl1
dc88NiXILy13mAyIryqq6EX28DYNIMA7TDINRadcToffDunvymLPxEud2B++vQJT
gnB6az8HMUU5eMTU7exmyWl0owABPYYCJOU5mYqPrhJ/SrH9mDednsPbvGLAfid3
7UXBVpSCEfjNxpBPTCo5mTs86oIZqjb8RLm6IuiMgG9Glv8tmXFOu7nYsP+SOD+V
P8nXavRIGmVfwulM84vKT2MuDa2mbGCAcgqKgZ6weiKvXBMGH5vT8SE8IUa59s2b
s0dmMOOsGYwpt6Ha38YWcqjr2JT7Qp41qpFFp02ptA8C4sUE9S/Vp9eUW7vRzPjZ
Js4PXRu7QiOXu4CF0C035BheWeoHa9m1XE/e5eJeAugfNXkI+Jr4EXAEbKMJ9Rak
Oknv3n/dw59hyMmRbPVVercRsqheDJap9Wyn0yUVWb9FIh5BsUUXm3kGHVHwCLOD
n+zCFwwbJ/SXUoQg+s5t726bRjXCU7NqPH1k5XyF47jhitO9RPsBk3527ZWo9I2q
xlG14Wa1NjN0/FwOK6UG5ETWR4ME+7kFpbZdwuFXW0DgurQ+azHjUkyTfZ7rB5qG
2rREYFpTRPQugiPsAFudbsW0rjYdfx2mLuaIUmML1jAdbukQfjiPDOsEONAGFGTb
9wdV+w37vLvv1CbL9OMVX1uSqCT857ECMbWeJvQEnGO7x33zAqyTJbQeV3LvlqNz
VtneUbw9E3nNNiDKdkAWn0VFlO1iDWH0ElIKX2e28ZeljjvWaVkE47OkInUFuDJU
qGsrXHzoME+TqxV2NQ50/VHepjtANU0ZA40ed1fyR9lWgttxHvZCtw/5gOxtopGV
BYW54WCbOF54bZZ8cjVpUz4lMc8KbkJvAmjcrdvEBcu0c4apajbe5buvSE6wN8BW
rPcy/AnbePhidJNqAm1ASFjHnWDOToXawbJoIz9E0bEqan6QG/u6o9zrZtNCQfMY
tA981dEpc9R7h+EKAiIkEclYIw4R1LH5RV2bmRtuCFKduTx1oDF9mzbaUFo0ailY
dUW/Urcm2jHGIzXzxpFKx+npsG9FntS4pZaefpZ0ATQL3b6ATF4POvDxJRfXBq1X
Y57OkJ3kBjRHzmEfM5PjSC3qkem0cf67/pzysvn/kTYDQXR7hsHbGxY8uCz2xHi2
dRbfNop5YK7PHHBM5E1a88GuMLew3DpE38pQuSAWVz7wo+q9V8RBgYEutTYUjnPB
uHXFtEmFH/Vv5Q717FI2Ru8T6cvKJWV219XtUNPl6j9i8Ud6Yj7WPso56k9u0UPY
Qu3p7HU9PsMiTJJH+e/xm0aYrfmeASwW8hqZRI6N8E5mhFZZjDZMvI8+JAUoylam
hbSUDwqGc4unOGaSm4pV7AWxHzeZrMjnbw4KirHbRxctcnMB+zPBtwGcEmv+MEU5
IWBcruY3YCteXvEJ3VMsWk9dEVKVeF0ufQrxWCPjuohkYOTMy/DKUm3m9TO8ZV43
CMTBYUj1/rntqs13ilEM8rhX3naYW1LkdXyzhxSYk3oaBb1Hk+tNJiu3D/gRmhhi
2C8H1Gi04PG2Q9oSIpKB99kdfBUxdGRKfp1aBbqCkOei16zor/+TfgjP4jf8GF7q
5zseiq8R2n8XbHMZm2C9GvoMoamWvFrgaEOUUmojLVYuaSGPpDSA3ZJzt2yuLNYx
Soqwb5O7DYa0fP/GL7NOEcUY0DKTIwMGurKQvIillaNssuKZNaDtMNZX/XLT1HjP
EaQiA+LvFJpX0CFzKE0MGAi/Puhx1Ru9K7u6NoiLoDhI8v+1fmNTzarOs+dnqYXc
zNmr0JPCkYTb1ukfWPJ94KMBVnr5z+gY+LmU9vhchkZ4Jo4PMfFzCugHP8euOwk5
PXv1ghTBPN3MwoEE5izNNJ6hX+BJez9bKkpnmvdt1W8ebLoq9tCPz/qKzGOlRW+G
jWEbRoKUvGGc/MaBw060GHm09/ikwTwDO2QqttXEO8xu20bnPOwKnJhlUcgQKUTb
EY4jvuwb8QbQzkpjb6AO7ORMvFxII/bK0ahkv7KuZN9jQzoRYmUqVWaU4o59zr7b
veIq4vPaqO+jgevHBNI1xWbZxK0MTI3sN3RBW/niVgDhBy8gCwUglfv4GWGl6cOi
g+KuA2lg7K1jhkg2Mx+KB6Ua5/+PuioOVh9GtZJcNl75PvL1vVg/rV4XaWDamJ89
/BI2NfJ/yqZxOtz3PjIHvCn4M/nhRv1ib4HYr3rK415QKzL8BqUX/0sJO2Gr1KnA
WkXvMeJV9rb0481a+n52kqdWoq7uhW1PpOMdRlW3fWgs8oNNWqWoaLBAt7E+z/fc
LawpPzM82ExSS40n/SoneiCsoMVAIuse3dEblIrfEVQphoeYF4e8BesPTx5Ef81V
jRzpKxWLegNsAYGhNfhnyhOnDi3Hs3bzXDXtqFp2KzDen/DJmsj1+cRaKZt1nLrx
ihI7ji6zP4KkSCT5OGd9ueLKxRcpYcKcd1fpaw24Av2pfMNX73ezQiUeaiG6ace/
cTRs4ZWmqIuCKdQWdR4KS/kQr/Ot1/3nwdl+uEO0DUk8BnHJEa/gx9UjJbZLs/DT
bUV+m9pObrbKMqi/Qjz04ox4/A8hS8VkoTgxk9Otnmog4nrHz1rBnpeMlmAqeK3w
SKXO4NviY4ZKSE61ako7eK9/jyahavT5/7pJsBSR9Q2lILyZBvoWTGHBq69B5+0Q
1RWsfGgWEAEw24jn7npF5zszu9dfpNwn9Nx2ieQswL4hKdzW62L9lTKyLGbY3gyo
2Mte6tVMwMBQY0JiCa04INCMM4y7BtMfBEHjPUXe8ziKjeA76Y9z5U0883o2JSKX
lM0FoD7M+8ZXgwLri7iRBoDcFnbUhShDbLq86iRiX5gjPxXgb8jKLtOCyAa1MTWI
ZgDy8gZBz5eVcfe+No+XJrfWmONzzDJSLm8I9DC9lHRggXiLA+/f+Av5gCis8XdG
KnycCHgf5d7LpD4b6PdAMDgUlT8zjeKBdDSsq5jGAFkb8XDitdtB2HpfH98wbczQ
OrgvTLDQ8Vtp9L/HTM5O0pBLmfqnm+dwOhYhVufAppVUU9e0Ke9NDUu2661fKiW0
lgt8TNiObOyEt79YKgIdaD1cHZvXh89VW5P29tq7VwyHw91ufF3rOvWEN6+8fiO2
42dJGk6joZngbBrWLotuD0/C9HjRFyHcB2t+gxI6siidnrGzhKiez99na0ubXkXl
aEcfGubeTDYDsNcwI3zOfRoOhGQ08k1401RHEKKhMBt/rrVDRljtTJDUoXYIduGS
0FI4O9WuQBRP7IT8DIyiHFwnH8v4FGvBgU7zfwZmqkEBzw9XRwlCvc9gHy3ZgdBm
dl8HCe3AD53pRF3fRi7FRpUtuEC8kViXp6PuNMQIUaeFm6wL8FF4YX/JvgwMkr+U
oGgjaUKB2eQCZCdYeeCr5wNeCbH70D9DkOd6wENZBkkASRMhbFZtOJY8YaBCe97e
MpPxdcgYq1v/slPt09EeJY4GOXnV3s1PJtmE59V8b9fhmNoNySCVLG6zpwSYIZ6u
+i195MuWFRwizc1Z0LHhsedGsWlIS+WQnOEUNXrgUxSsvvgHMk/arzhKfV2cBDr8
zXniJqgrEFeAY8PlV3fZnPUpGCt+QLg/rPgQbry7ATr9e6JubObwV3LChMgSM97H
SysRq9vBtDfy9EEBTDRCojT52Mogav5azeehb6RHAwNv+e72RFztJwuDgXLIaQke
H4h/Feq1BRiQ7tU+cSu/GIy/qhUslKUFYyZVpRXMEk1JcjILqymQbe1iGAre/HeY
bOrFCvaYQQ+ZtSpeKB+4iMPPHftve+EYT6iF7h6k94bEb91MUpdRIt7Cd1Mv2oNV
na6jUM3iwzTpAcGdcLqmKRujmwVEn3FmvXag+TEUfObbmF1ugaeM/NIHyNMtUYpb
ojSdRnyKvV76cGdO5+orQY/0h13IoqKHTOHB2zSwNd/keqlLdVllxaY/Z+pI/i5q
unVh6GNx8XRsSc3gDgx0XEI3MEbGCkv1gcfT5GXkyx7fMJh66Fu1wMO6qDT3FpG7
zSR4L6MKp58N3w1tNqfY9SYLAlRBwjZwrrU7Zo0sUDYdasTQe3VDIWID40BDIBpg
8rHZIH12tQ3QpJuSRsGBPl8OF35AR23GUSaP0O9f/tzSYV/4RZ/WNjzvd4wQzG0C
WvBJ9nDm4v91aow/1EYaADhDWUYTlyU+lS93wMPuSUxiXt+K0shAeMmS3MGHl+6x
9WD+sWbJNu/J0YM/adaWAM3sk8yaXu5By48Mk8sqMEGu1C+q6JVrswM233oikr5M
LMySE+AetE+hQvzswS4HeBkSd+/ApBay3U5F9sG5antZR2Bksm2eLO+Di5phFRp3
ONtg5IMWjR/qToqa08yRDARK+7Jq5SFd2LE/F7o/Cs/MxjB/fYmM/tnRWSQRLZtB
ED3sW1FRu1uuvcsZh6GLQ5ZeEsHXMScOB+EBOmmyaB8AYk85WYF9rCOk4b3+cvG1
xjVfqbYiAkO9dKqMDE+BxVVM6hfEwb+WFYMVvaNzzcbf0BmEAfoSclick/c6mk2D
EcIvgdSr8V0s8INTLz2bYagV1vOlgbSVOU3ZE1zrHMvtzt52C8DcxfRpuHawsDv3
Qri5aNAHnMhYZZgVPqik/N/BLHS6E6yGdouJfjDNGazmxYYDBlTkamaWvBpJYdxm
4W1nNQhnYklfadZjNfjJyCVRLE2VtfrkiOmKub1E/Ku0yD0zZkJq7FAJAS5OWavv
tCxx0sw1nijCfkUldQ+uXSivmJMMeqLaSwxS2QXe7C/urc6AVKONM8LUq0xOSqvW
Tfh6jkALYCRBfeFl16cYnL7cwM6ikXhjdbW8CHF/Byd4tC0JlXgOwsP2gkpS9EvU
agmrJrhayCt/2ZPsj8tHXMOvxLo0rGapspSq+YBYSbZp/m9XAQUM7KgWojaunqgW
qh/CdILI8r+h64D0JHfRHLtI1RhHdSE7rWIPGkCBZo/Mx0zxeqvXypw0iZB8HGOB
XByouJ7D05zJV6Yl0/htVlU9aPU5aOYMGKzmMGngX+NU3H6WSH2ijlSSD4FiTzpL
FsVRVGxAaRa06JvYtme601CnzfNYXH6R0oaMKCEP2ZwpJem7vgGppWbNTmUSFINk
yIQQQv/QulvXxaNCjPVbIKzyY6LwP9kFFkoumvWM553tHC1rQ1O6wtu+LHWeags4
h9nxUHDeY4qXcx4xdQycFJG+9J+2AmB0iMlVwXvHgeZaOsZ5kb7Cb72HJojm4bNh
yKWTejfHA5cMRP4kf7LO8WlqvAetqasq79elf/FbuQJ+i6Jv6I+XCfVC+Es344U8
Ir7Rkb2vmxXAfwG3MIfJmJhz28vjYeHo3DvhkVLkh960Qr4hzIhNnVrzeqJD/4x2
QQ8FYNbs+JP5IlchTGYPPuA4Psg3jqNLH8VgOoWQLRRcaiJGge9lMSmoBElV8RPY
f5G6MP07Le3LoBCUmiAe5+g5ZQb5DBFEuWIFy9T/AkTTByE9EYVJzsSQHC7f64Lh
LaYuzYFNFQ9kJi05oJwQOzvKpykd4wM68WModsXmo+yVGpJRTPo6EuFaf2+xk++g
9mLhC6GOh8aPrelzsf6kTZH5UQHqJW5uGXqEiTYaTn2SAACz04lzzUDPfWPxkPHj
fbYhN0R+3Qw1OTwpSv6HgRRYMvh8bJuFIhxggNsohjrZ2QAAr0i/kGQ4p58ufTUI
ovDDR+hr6Tgk95yh+0Q6FyAVWFurbIaTAmnNFb8Mpj8knXwaqj7t7sFJ5e9Mu1ZU
WzgLr9YREye3OmgyH/7yvLMTR6HjVEqoZrEE3mBm/0iSPV3USqgV644fYaXDKgFP
ieL/aRnuhoyWnLlI7qlDWdi5m2QoutTopGWnJt/gjzj89nh9JZs4agMEjFDoo6PK
50QRac8PQU09nTcD2q4WfDtzuVr0Zxv0kH1xFj4wNchZnEkOeU04Ga1dlnuCKkLZ
9f36wK74o1ZVFAQOubz/qjYpkk6s4APVOTY570sc1f8Ug69xkiFfCdtaMinD7VZz
TkvN63t7NZ6LbCYsD56mQ0piGSqnkXteyKOKM8NyiX4Sd5PzjYf6EFusDfV9GrFl
YsTl+p7W8FN5ATf3MR40B3gKcWnOreDA1N4SMLFc9v2AUO8PFh8ujGZXhFdlCUCr
nbHvllp3k+My2ha4DHtOyWYfoLGvAKbHLayzqmqz4ocxfczvt3aQb44p8hyNyVW/
jP5jC8GZ+ti1oMcvHLD+WkUr3BbfF2c4mS6RLUiT0555W9gNh4//SUyLpM+Ywm9u
Dja7P7LlelEYdxnVOJBOcIEXzcCmnl3DZm+AEqQKhaJeB6TWyTFwNI1Za1HW/klg
lytfcN4QdSZiLlhMAo8kSC0NdONcp8MO/gCtOZ+ZNb/ygjtcA25bO5Hcei9l1Nvx
ekDfkJoqvBy2qBRod2XrMN1hw6xFL6zZZCBcMcDQtGefPkaUBKGP6oJ4lNptJvGY
B7C6jrI57tZghIzSnjBGe7FtgxAWPZxV5inv23idfkA47zw/Qc4YM91n143hBBKC
ZH0D3JM9lrwSsGRkM+OCTDoqjY0zD3zPDNKIl5RpPcE2HPjsjLfaoBBq/uuqxAuv
jkYf/R/OFBEITjBRV7DVsWGtW/GWoNoiSlIWlEn11ACaMydKgZyUuIWRxZhe/G+3
G7Y7smvqanaypEQVvdB0nbkaBpw+8G+CEW1ClH2rwIoPDoC9PEHh8nF5Y4gj10v0
fkoG4ej07GNSNeadASkDLyXg/Xb3MDG8Tej/rLt2UrRixRZ+/+Mxy1MhHNMVLEOc
iuRRU/AyuhO7Q0SNDe3rVrQ123/gjwMrU8dB9icV+rTCwpAwMeEDyRCA9/nXdYF7
A3wv5UxxRDVOSgPPoi4PT3wC6+4AXkUwx+wYzNFsJ/XrbDUCKvFW+U1HuMVfNu8h
IqVSz/x+leAGNsCGdwZhrDprWpC9CoDY6O/m1PegzoLZiPA552kHnstn9qa38rMI
sABiA+hCvOUi5hFeT5hwZnEX3tM72RevJGDqWkpshzk/ERrgm2zwkdlpL1qojdRj
8S2KgpUZRU4iLNc0nUkxGDJzlPDwiek3WdgNFA1rbiJPsGmr4RZ6UT9syAh+HKWW
DpUtNQI18lbnTGA7gk7KFzE0hBB0s7Vaca+KuOp/4NX0jiv81+tBVxbkKvcAKeDj
If65RibqIN8GmJk8cjtmOmuF89F0F3Bf3n2hiYFiQPYjiLyh3wnr2osSMqaxFX3O
qmXFrZSNgbkpvfL+vJwLKMeF3GXv/vVRgLxTjHRBLFmovHpwOJTbh0w3rsH2a9e5
W8EX+4SNOLdvesFhY/LFKkiiZJL9c9VQKYQjCxvSGxOSzkm8O9tvtfzNMovzVmER
hkmTyZfItIWBeJTRTcUYnkynj1N44M3e7OtYqxIYH/3pvChiyop8ytBaLErlUe03
tN3u+5QhH5AMnlYbeSKBByAEii4ZdpUNmX6JG50fqhmyUuPngP4WzSB5vVU47X40
KJkLO9coYgFIO3gKIfESIDzaV9tiiWaUCaCF4u8MpFDm3VS2NewqXAJWEDiaI/sy
/H5rtP9OeHUW3xwGTZ5jdAFSs+LGk5Xv41eWFmisWXH8a0ba4nKv1XaPN4bMfnbL
DsJtBmblk+vnyTi5O/iDo3hty4zf/jEysSVROSJGlpVPpe20IQ9Kr6q7Yd3d0FSD
8Kw3Y6VA5KUStEdoj6vQ4xTXaavLZ1o+/qqyTKMSbKlA3SjucBLWL3SH+ygo2He0
3tfOk6cDjawWlasSvqPoDXn7NqwCv71/G/Qp5RxiRuML9UZfSkXgIKJSdocSCvlZ
xiO6Fb/Tros5WvvoFcV2cyLRyqqGibL09YmeM++xOFyY4078UHFb7DlENeyogu4V
PoGGHg6OkumLiuW3WVYp9J4CXW9olMVilisq9AyGIKHMFE0kE+ol/jsrGay77Edx
3MKTwnFlfGJGObUHRlhmBHFMAHnWAVtuG4BbkqZQne3klGqhIv/3JWCJozY+hZP0
jfyiqbOuoag7UW8lTqc67uMfOMei4OBQkkP4sHX+lGNmjd0uDhW3G539K6CuBgBv
h93AXCzELk/7+MDpqxXGWehvnvA+yA6qu3HO2thSLQXCBH6vsVhZnaOjWmslcIcF
dE3bplCj6AndrMFMHAMTkCDxOWEjzOWksZ5l3lF3TOPohv5IcEefI9915yvV1jJG
LCCJ+iR2qcRzZRFNrgK72tArAqjU3wX/qK/T4Vz2+JrR7AhE6XOBKh3JKsDZXvPp
tvdpdWM79BLiUxYbhEACFvcLyfjlp4KTYATwSE3wEJ+DnSH6kPLx4O6g+G95yC/O
C5uiQU2SBf9cdQVCffd40ZSHIkeushvk0QxWKWPhZcFuVRhKA0raf1HfKwDMYxq+
S4lPfcFixUeikTWU8KZBB/M70usjJ8WAC96DdreVTesMMVB6qSG+Db+jTUZwuQ0e
ENw7x+hGu8TjRn6s21DmYxp2rmgCec+oavd7j45mwuZhxIE+d/ZxrICz3PqEeyF/
LWPINW5gXvUuFwTcsQjkGKVWEJ7Gmmnxf4n6mRDjaPTDsCrGVMW1Qm09MhoBvFc7
VKQdvI9WLuxafdVu+5cowJH3VjkVAoDTLjbq7MBSBUzEig7LQIvQnhmd1AD/uBg2
XNU0wbThwu8raJTdvTKEo3Pykl/n+vHrO8tiunc+peNAal4Og+ByPUJjbe+bJ7KB
pHozCpJ1P6gbls7rqgQF09Zx3CXr9ANPjUbFt3HRLhspH9qq/A6qbFykp/HRG7wC
cOiyXYSBOK5vP63gaBriG6+y2WfTVu4LxDojbbmsUbOoAKaJ68pkO531elRZDqSZ
rLXkPW9VcTN6PgT34WX0+w8QPr/mfKg1Tikv9VPHFbqJ/XJLR196aMHcq2os69nc
Q31AHdTB9xJ01/+JbPOYMN9ZaQx/ZNEyI3sjZ1hQRq5zgJpRg1yvCkEhHhGh3KAM
zAdAy3WhPmJXcsMjCNQAV7br3czCxm7fTS7IuOywVT2apSuHJodeFj/oIvEZDvTx
3I3HPoqYebsqXGvQebb1FIR9YmUuWuXHPV3QaCTbbOOmAZ/A6Rqv6zPfQ7oFuN49
NkmeqfruvRgC5j6+S4P4k54J11hu0j0m3Sw1Uyn5G/6IiXfflDDsU0ARekm5VOOX
9l3ZaBRmKkgdG9Kvy+4sYqbQy9tDAmd4QlvyEaGftx62jl9t3bRYD2YK8pknoTa6
k76F90voumTN6kKsc5VVzPul2WbRtjIIxIiWypSwrRNwW/ud8ZmcD9Jv2/ki6uWR
3cttG/rfZx6Oychrwo0laVPBu3Dyv96CSMRBN44tZyBfDYTXy1q1dGBnnI7YH+4a
E9OlPTvB91ca+ZTCx7qxwjcdqbcc58T5vXZzWQm8YYKk6yGJT5HniRLl6tcfIR1B
jaSdkbaxNjQm5ZDKNHoctPtua2OgELBYmn2hnzO9D+lV0H+g50DHrKwWO5Xr9foI
ZFfvOaLs2oyCseWKrDZe9GAIxxDQ+bsBdz7+d3CbKwO0rYvNaazCeYvEcU+V4OLE
TAR6gy6Ua/nmfO5De6ns5PwzrsyguGDhqvsCu/XKxPl1lI0bNu4iLxHV7HxfSbbW
XkIGnv8FfhIiR/Jty+Z1ifkiCpyw60nygHthkcfaE2ebH7yTeVejqvhvXvXeUKXM
EeYbrU2Bc5Am1n7tQB9gERvoQ3YqsZUnwO/jXwy83cmKWseSdELhBuIzOtBxfYQF
s0OPcbDuzYCKqUohoYs7iKY6Z6ppbR5qlMOjIKqAXEZuRqc04UwPLVNzh1Asr+AF
/HByoSt1mbJKFmu/S5MUvmqq5ZfNOOt8NKQIhJt4BSEUAejLX3EYPrf0u+mijBlo
uoDVf3suxfj3MZltFdRwhUZp+5algKsdXkQX+6B+dBiWVMzJoleAcs921Vf5TTrQ
uXdG39kr4oP8fECq7FoggVtnOzPiUiXM935rW6sjuhWUMXbQUG8UFcqurqi99K2T
TvDOHI6/CgzOhDRHkexTJtJvmWgwUmBvU3jNmJHSogiNtuFeXCzFBx5AmlQVRSNA
Y7gFjoxWeENJCAVOgOVNzAHCMre9kaWJ148pQPfqYjxZZ+U0FOmF4NeG4znc9njP
gLaFdBSqPVha/aZBzQD1mgkGLZSwRJn3BOQTP0RlwqVIVvtZfjNymdElvRUE8+sH
pYsnJfg8XwsFTt9iY/eEJiF7N5yitiwUnko2xc+S7t7S+L4+g5vDEsyVYIE3QQAJ
BDunGQgfqWDl8mn7AmkSeVZvxzLAQjFZf0eCC9o7/MUnzTONmET9St3w1FyA04kp
aLc5mctPJN2S0ObQ13UwA+MOK68bFqvfW42uW3GIb59GWxZxbDADRm0afhIRaoL1
gTVA7uvsQfvPuj1rRbZqFgEKxKOdu7lnfC5zfmXlcWE/UdP1Vcmatkue7/hd/3WY
dgKPwPGaB4miZ6tMPPyoeUFLbNN88VHtbVNrjfXsG1L1/sGYjy7tHY0wuVK85ENX
xZQPk1ySZVvnle989wDxmhj26811bn8A+7+5ORcmUabpNLGgR9QZNQE8cASLjfT9
sL1AcVo4DugOnYSIpq/U7MAjvijjc12lici796dkwWm334c4RLPyAQm+bCtvWKng
N+qdGjjb1JWIL6IkXry6t0P8VrMkvYgU1ijJbiGS0rhU2S0waWIEZuwAfbh6TLHs
g3A500FlQSZN/JuZmJLari7y4O0ZqWyCjeCvRPmd/0ceODuxwfy16L4VNGcMK+QD
9Xqc7JPQCOYinka2BWvcl8z+/gjNVWKS6NJSBCBwgg9kBXic3QvFbGqszivNeoj5
6PyuW6NlfycBTzdEFBv3M/bdsC56IS+OX4HiIZFNfopi5VfWf8MzB3DDGGnnQX1W
NZ1KnPjKpzSIryGQsdFw+x6d2HFY8ksxFPJSyqNmyj6orUm/cRSOY34KFLx5FFZw
/BhSn+KxBtrL9hrJ2mZG1Nk9c1uXCkqbl8aYJBH3HUKe6A9k5PDRXbovV3tDSqm0
z+1qqtLew0WOt0QlDludsBC5E8NTP7dapqnabMdk6xoieZi2NoZ4oRzhO5j3Z5a/
sZcOuaCsc1BWi+U+PCLS64iSthiFkpRBanj0pSXMN0KXlKh05CSC0XyU0cg5KP3f
TODtRAScgLjax7us4tfcJZc3A0EBX9Aor3ORjYkwdNcICKSG2URY7q9V9p43oGbB
yF2YVYh48vPAZCbVB4A3Dk5Q9CoG0cOiFqaY1lXQJJkVWZJiAwR3mgM8jHPaehGs
65FCc50Ec82MXjgHyAMts5kp0+dLXq288Zc+0OcoM6ahXQFr4yvghIrtN5KHOp9u
u8lsjZfMp4tak21xIGMf5a3veJWIuP6LJJLSRiu6t4fObXvAVHYHjjH7Hi9tF8BJ
McJVTNxH9uLn/iWw7F6lBV56ltLC+OOIKU2Hl/I3GE8hWXU8t/pNXJi3zZtQTc9w
FXtoV/S3ZHgrPk7fOmrfddNcIAgSXepTkdseOiEmB/48MRyBfYyLjmYj2pFz4orQ
NFJjigKgwOyJxKGYtYBmAPhhihsWv4K9pa0WuLDApHeX4CXwBGQZ0UhJiTJ1CwWY
ueNEQl6GFXFEYGCzSzy3sv+d4XisdW0u161wMpf6rGezWW2E3cncCZCJb2/nkmR4
ltaCFGtLUpkhokncRbOIbtXXKTPbEfe0BGWKgET3NVbc4EYziU+/WEp9AdWXrG/Y
apE/1/KjsbTh9a9VFIOSUatrPTnV1kbU9crvT0IViNq1txa2NBkHBJxvDB5wzppI
EwIkgy2qhwUufzxsM5V8lOE3D5Ntvy3N2jhdno20Ud39CUv0o5qA0kDA3Cer6Vj6
ifsTOXpL5nadeFUSSdjZ1Y/T+9lFaFq+ET4ZhUi31qpHp23MSrs2AyqsBj+SdJqV
bwI4QuYVawDNMVplL4LYqFLpIPqw3nVTvpE2f2VzNtOzu349XD/NI1zYlWw3jc7X
KHEufUO7gd10tDwixiiMY6eyYfDa0WJqXHeq4zGUK6PZ8KIxCh8Y8iEJieuNb6u3
fxJlNMOq3284Bo8DDZkTyBVxBDgwK6MvpQNKYISPZoF1iTQdye8unO6I46WzU1Zq
JTSZqJNHSSHlKN+NX1BPYtUS9fhS/23z77WQuSQp4xQPOeSy7kC5pVwpCjSXRrnW
ozvbQ+aLdqiT1XyABzZbwmCfXPphOAO40hDAyzitlXsfzLVnYMfJ+3c7fqvov2rG
LPlzf0+zJIJ/7btywQ4h4vLwOxTn95RbZziBldXJvB401ltcK4SSnY02yPFowxyT
G5N89Qb28LKFehF7jza4jMrNaLsOuG9+vGR7/eE/3T4Kls2YvNzjURj6YCd3zgN9
fdqWSl4GYl/jXEfURSyPfqW7l9rdZJtD5k0EpKfZ0QS+0Yo3PRVHsfIZtEQJtCNk
NycQTx++yVpVWcxoI9MdSTrfD/s+awmHh7l6Q7H9CfDKrCHb1rTdbo7S+hIH2EPt
RNfcLjKFhczVoFwrEkGsNjRiBnE+sWO2gpB379KIFxl2d8juQ/alUrNYJP6ST6H7
kVGBOrtxNeAdnlHNkLIy51y51oTJh4BvmOCQNo/V9MKQG48htbtSgwA5C0WIyWbT
OWXC6VYTJdsER1N677SwgOTVrf3rDGJupMm6OoMnTEPqZEE1KUFuhlpwtHadsX/d
dQBIqksxdtKfL27+w3f9wATazV4BizymLMros3qSXk7rKhaFbWBOni0Irv1t92rZ
wTvz8n/ZcAw75lIF9H/e760QUhX+ez66flUJMI4k4Zl8aaGhxQO6QdQYQJftAzxT
iQC0L/u7FWCAQF7ncUxfvO6sOW2nuwYXdRiUxfuOvAUVLdyG8gzAJJunv76Alw0L
vsneoTTkLtxOk/gfTj9/Efu7Zxj+VvfJ4NTDjbDaWT4+5E+yMEA+m/AHsGZHfQW7
a0uGu2kHkcP5mZHHOVUMkUc3Z9o9t+ASTX3o4U2f7Ygad7JqnWVTn+kCwTFFvTwE
zst3hDyHkqXeouSLGgwRqLP1mEcXpqUaTwwyX2epCLcxWmN4G2DYJNBZntSOdD9U
45UBmEXpFx/T09vmCJlv+ZRGPXetLTcg65ZUUI8SSAbUTg733hSsUU9nRYpZ9Ga0
BuZ61B0ySkdoFC9FjCpH30+v8EJ7xzlIx9PtPhYCBEbDecmJcVfxajZSxAJeNyRg
RQMzsk30mgxzjgaqwpYyph3IdZX9G/Bw7jBBlIIPjaZqDst0u78yfzTmCwOhUQJd
5X+Du/13FSVP/NvfZNRhkIp0i59k5PbevXgCBowymAzFPTENold2qjY2FuSfvXNf
I+cBsK50ulv6AIK0YsvQy8czZ3A/qtDrQZMfVkV7McRBFVDJLTkxWq1EAkZhQqfb
kt114yiC75IaDvuHZZjncCjNoBVq9sfTyoxNuef14+TBtWw7vNpUGr0KyOz8M7uf
Uls6OX88CBoCCumQoChrMLGAyhy8kFD+cDI1Tv8ym8kemVQ1BM5l1Du2XjMgUV9f
+RfiHaU2VtJ6az+4m4PRv+skPCTY/9pl5OZu6i+i33xBhVZ/xeGr3WjZXvZNN+89
yU9A0YRwWfjHZTY9N1kh+FkjmGhUQzKNWm6YHyhAZg1EHyi/bWfn/T1dCC8xVag7
oVjTT4gGLVRl8paZBzCYoiKc7idgmWvHHfwLyTwptC32uVSZT9McKbjQnPX1c7rg
U13XKMobDOslGJ88dqDLtdrRmicGkc4q377pV9kc7FpejzhgfG9sWWbApaZ6ziB4
+XCv5ndfi0GIYY/1fmW7hw6HEQglIntGJ0C8m3swfPkXa1tJDj1+RtGbgPsFMP1i
N1YTGduTxlJrwb/LXSASLw0/hZR8YXLnSdS74qLmzV+Ta59wDejyHeBZBiyNITbV
dkMNVw/1OHYS/H+1GgKYJTVxoWUqn3EQ9/J9m29CM1W67QAYUTJT+8eaLsEN+mvd
vXkPT22RlyaX7DOFGorw0Gu7IKHTUFuOUzGG7E5aUPiRx1ySIfVsG15d+uvbI5Pq
WT74R/NZpzCjBnizyTbsY2bZypAiINTnefcOa4dLYyMFx4NabygMO5cKQdgrnHwJ
SSnSBZEvz0tmrfUsojfkx7LkF350qdqEWMeHjqzy1ZGLMthMn4KDsmbRu7FCwLyP
qmR2nC61xG+wbND8/DT5EX5bJ34+moRnllob3h5hgg643+LNYg60PUVAeLqkqZVP
cV+JLe6gMMayAlrjnIZadeKIy+tQw9JNE1VBLWb/Cqj9HjL4XQ0B5LSsE1IK1GuF
KTvbkPxQntdhE/jfUATdkjAI8lxH2piZVpkj8fCi7CwGr2DI43BnjPK+fB9JEGEy
CNOpRgfxDwauvT4fZYUX7Bh+MycIUxV2RObcDD8zU2sXWFYBO5HVmtWPkplRBXJ2
kj4bhzEG9CoCXv4g3RyrNUrAP/KLpp8yzmt8qHS3hdgZ7QVdLEY3ftNtpu1Vcm0o
RtiJXo59js19EXlafX7OKAWTQagWTWa+Wzt33dZRbivOUfUpMI6x6M+NF/ZB10uR
0I2k6qnwlnPFKEG1sDKTnxKiarsUvDHcJqdpnqiU83CmowgT+KXW/rWPlx4MWS53
nLQB9gypQZfuMftyM1i9HTC4Z69FRhXwQNPrf5kTM43Mld91rXZgnzyLwRUp7rg8
ZzkErGUiieM0maJuqKjSerQK4o0FyECq9zTloo+OuhaUYjK5eUx/bG0dcQd0F6Lx
qZevYtbbXvnZozjmYO5X7OsxEFLBQgw0PyoR6Z09zaBm+VqJJvAOlY+bLDb9SBwr
QZg0HK+BOfSk+r7hBOhp6fF+aIGLPCmCmlWWTsGP9sVN0Ok4fIcj8Q/8OFjwmXNP
J0juob11h5SKkNRanbnnyMAm9zK2O1l87tESGexrgb/lcDssm5oLTm7we5V9DN4d
aL9aAUT9Y3CAIBr4SOtTNG8OODgm3AorQ7kVLrV88PBJApfSg+V5M+OnuG0sn1Y1
dXh0TAMqB6RrWAAdPlPtlYgscIuThi2NTN1rQ0V0+rCTK9tMUq3ru+MWHm+cOpXO
p5Df71Jz2PkMDnWD7NzcGsbeonc2V4SmwLAShTksFODpCDg6XRAroGe7g42ckcaE
rBsQvhIycgswOBowGe1gCSOeHqsJZOvErlPePz8PnsriCApDoSYhxBm0DjMNaw1K
GJf6U2GTXu6VW9kDzIvuDnd2xTt9VyJKEa5eIygL4wQB/GYDq+755edmMCild946
fssb5+OA6gnfMWyXbYCvczsOEasLoW56BVYikVPIXcf0fsZWfkr2YkAhkFzmkFge
E/wXzBzArLYvvijYJIEpD07wYU/DMTBPAB19VUvP5gV0B7RSE1fzxkuuSSeif0oE
Adq6I1ejVbQ6wQj7HVtXTBdkW4HCAOldyBeCEjbzMLsGAKvN6Ss4M50FLf6wdb3u
iXVmoWEYhWlwx3UCzqTttO8FP4Ch5+HqbBY3Ii5MI+XVQuZQZJH9PqEsYlbrMcPe
DMxn7hJQkLhy8la9Kiea86bVcelSDBF0gOM7AcHiB2h2VGgAO2GYUUUXmDtplRul
SURNY59AOatZIlXHLz1uSQy9sharZ+3AN+s59cQNJjTZ+cetmFxG4tXqW3YEhc6f
Htwm2Wt+eK7RA90tiM1xy1VdYqKnSol/T17h0bUQHPoeO+3UFZHjhQ14fjMb7DFI
ZhkVwL1J3eEY+wJ2/OZDfdEdMtxSMtF6LSXe/HhS6SMOzbUI6sNM3/HIqNqYjVuY
R0n97S6hzTvBFUZGcvp4w1sZFh6S0+GmJ/s54aTRHuT/XiNuJUi+Kqo+4UmLwWxm
vcfPMcKhIewExgTzNtSlJnnxHjZWJ15KnZLUhs4+M35uvij+hRYPqouSMR18QdWW
vBSJ0BReytD+7UsN3da7QkleseiNOLBC6FzwdWOCeurqEuJeN8AdvDHngmqlu0XH
lj9QalOipW16eAmaiTnAsk4MzZC1X2Mpg7MDnfrvD1tnoJKI8d7TBup+3DIimV3M
2P9JdZHtT5+LdPwVjj3UWljG35VXJd6znkJAmJGQ8pZ7PA54dlJ5WvEZECZTQwH2
H14OmsYJQRtaPIkbkPBNgynwG491Z0275pBTx/dWff3lU1bcu3SFQidsErmsmqno
TShvMkuWwScqE2VTFZw3DOt7gtYFP1X9NW6OGWnCY1drAmsoC2NGNAuM+b829Uxo
vRvHjSRS4kHmTQsLgZt/evmE38GJxMpZeaQcUpsB9NYpCHaZq122emarNZ8wWwG3
fwchv6OxvT84Vo6gQJF9ArpM5W08/XyVlvPhd9M6BYy1zOrLkBB1Acu5b6JmU5+A
FM4VCN9VrDeCyl+imxFs8gR5Aii79N60LS3QoNF7BsXzVFxchMKA8Jui7wRARvHq
lrepGGTztZxaVq6WckYGptmuaAV5c6jbq6rm/fGtuHzVI8npt33Poc8l/509Uucc
jcMpmWu71wr5tcf4jpnVJMQ8LWEkZfwMk3jUQxL8PrL+ked91JdZcS+fuNxyTTnM
1SjOkspy5Ih/plNGGxHecpGtEYtzDyKeK+4rLAOGTUAKX+h+VMzoTE79YSuepBTx
pVdVMqgT2HOxP7Gav0mNDj35SnySzCQyUfHv7HsltHws3huNarm8EK4N8V5DxmGq
+V2F6vk67cqm8WYN+npN/6BR0ONy1Y+Z9vtP+3AXJLs0rWhQvjPnw6VDghhmFlQX
xgdmhyDVV6P+s1zOODne7BnZSddVPOmbsYBmzKO2OI8zT8NpkUaUitNVcjKiiUGf
vFFBR+wgJytH4QGmw1kYX/V+Fy2lMm5nrMNDE8gRc581jNqXSVI/JoheezPpPRtb
LZlL6V6mXqkUr+bpXDoQNA8j0bz8InzDDjJxV9Qg0TxPfrZJ7wiQ2zBrXMd6NXGM
XbkDCV+IfgYF+5NZiGFtg8KTG2hzOAK9Y58B4nzAGo1MOVZ83YqLzzyHbkmLgVqs
4rzpA6IMd0SkJbNQHjAPkCnuAUEjlsXj5vxOrbmDAYXMv06nwPfRlVHB8JtVv9b9
RZIVtDTsPHP1AYkb8uqe8R1KKywgT1W1prEnEA9T6xiltXLI+BFv8f5zlRvsznoO
I5mD98rYrHsXlPqNYckIDETZsh6XYE4AxGvdmj705NCn7mOgSFuHZCinhUo+GFrT
nyjAANqRNbLnPpqWKHnUPL1fOVmgswZfRTJU/45FT01l2DHKRnHIf4VqpI/EPGls
VH2lLNKhaU7Lja1HQW0H0EHfMSLKPkYZ10dPAmvx1NKlibqz029OQbnLyPrcCig1
n19r0x9NbCEpxcd/A8oLXqj3bLNmbahnU0SAttxokjEJMFzU8/zmuxXhFQeqrzSV
WHlYaDQVVFkszsRbaqFtsrgIfiEXtbdrvTOL0v6c3ACfkYw5vLPKgP4yreXJx2gc
2ZzaejS9KPICa4M+qHFr9BHOtklV0ljqFwABhluJ3M8e3ko30tQnO8hzgs1pK31k
+WrQyw0qH5sL9RTriJkk3rvq5Rxzk7UNmfVt1zKKvGdmFLY2qnCaEyhuPQEJoQpr
N+CnNeNaCr6FKyv4hW56+6eCTRRCd6BTl7eTdfKalwtK4LJ7llT1PqCW8itlMysX
CIveZ2jeh59JBt6BVNHQAQ1yvSzYhwnNLW+YSV34U+6i7fjQhcAyoPOJHkapbbUr
OZgNtKEn/u1z4rxZnWvHXEnKn2VxTcEuD8IPLzYL2MUar6pDQlYadyNng2+YcxDP
UTVMytPMfYUujX5cE213JYII5HwZxB4ETOSLExxLc2kH7dZ/iFafLL4O3E7i96Lx
CsglFrMzHGPp4290O0OVgcG9nfC3vwoWMyw/GQA36aXj9AbspVqxbJ4C2pZC7aYt
E6mjUJqGx6TV6aeSdBhSqpUVIM8P9ApoMvycC66vi7XQrrQDsbEhCRAFxXwaklxv
r77+3Tkz7ZKlUfU20opM7/tapTblDTJbjOs3ua5jx5R/fSfladMzwbNjwltNdSbK
lnuN2cKm0vPacZcNsxWEy8d3xj7ejKBS4gnlQ6Yf9BHW6a8+erZuxb5mdxw6+icY
z33dS+r3ZzJPZS9ziqqOYw2dm1EPDyNekj1eaZMcYnrLUMT5x6iYo+QteBLDqI7k
sjnl+mYwyZw02p0BtJ7H98pwJB02MFMkAGkDDq+9dlZCL2A5SByCMFERNa5fv39y
JKBC4JbpazMx/fzE6IwHhHvlLKmVal/sCVpWxapHrooR13mAbC0KU+B2nSzh+0Um
5B51mnHIcaf3EXQq+XRWybJmrkV44xsnXAx4XXndIFNiBuXq+2t3/CKG6SpO0OAv
NJqVSsGSKxeWzrUcp1cH2bFlEJitmFSDoxh7gfNJ0+3Rlv0lUYMWjePM4L2iPEqQ
dkvp6L24coJXGv4CvBNXjiIobEbwVDc3ond39uzjO0wKNPgEyvxj2Sq4JJHmvAQ+
U8ReYfIooMP+RUzwX1p16fGUeEzosNEzTz5y82ZDYIlUUie21C8zhWJxk3UzyfYl
REcNw32CW4zTM7X9iqZD6e8mz9dFUkeqsqrdG0vGFHCFOq38zQ/pLDGCMYx1g8Dd
L3XEx+CiWXwhO1V/t5MGXZzuJHVVLD4V01XMl0UMD4mOoCwi8NuxkOvF79fyZg5o
j3uE2WqmvcchD9HPoFWv65uzfARzglviS6fN1LZo+6YyrjG4dx/ehSF5nTb3yIuT
f9liz1NNFhoH2yLaVJ+mU00ebiM043rbgxTH1QRYhjqdAI/D0jPrlZ4cxcDZnYeO
XctjwaLGGM76qQ4zM7sB8roNaI2DX7xuzgCO0alIze6+4ZcuRW+dtMeFTnMpqCRr
jUfkZe/gQE/0Ub4H34mg1Xesj7xqfQJk7+RXjDyNKgxlXIous5rKnseV+yCeKxph
/Z4DnN+gNtZDppafVE0qr2YJDmie+RMV1cJvEj0BO0mg/QEaoWjgnhKwkAwZ+6wW
WfVJpvv7jsVnb5HS6ib4yUUbJTcripQcT1H4PpfaHRKQjVlTZDUS+h//D3XM5ve0
0zy5bvWpxG4VE6p/gN8GGioVAEh/dHHrTy/YKDsgTLn3ABpekIAmObTDMbhB1Q0B
XPOI3Nnpfn0HTpa35sR0njPZV0cfkn6mJQQU8ZefT3mUztRzvHX6KLRo2Zt3S/b8
JKv42oUsun24jX1uoaIkinXt0TtlrHwmBRU2XN2T+501XaRo9IpTpe76C0rLzjAN
o4pJMD0AhRtNgt7KJkYZ1e49ZIgHCnxAbWVj1R3mKfHgI1eS3XGdxrOVl7a0s+xP
v8CYOu5Y17eee5R+epVbHpnOW2CCYYhYA6VJ+VE7cO6AwMFx3DoNUx/U8xarqrDv
dEKmy5hUF3vBRdE9Nu98GhJxYbyPkk38FIivINo05qYRYa87v3l6LN1k1gAq0KSW
zS9RNlJDZIpX1SuB6zSoYr2cusNCXn2pGuF6fFOMz5TDKHLJGEF5iSi0sBm9LNDw
IUl6yA9dRPAabHQ5vZo1AeFg+feT+hmWPPcDDNf7aR/NkQYgVshu158WkKnliahy
ypFT5OAyPuIQKTiFzHTFvBd4rVqnXR1+l2429DP3ZcAX31HOi+HD1BV3xcC1YAGJ
mGP9MiHl63tfHxU3jQQq3PuFV9xzVRSttcxVj+9fcRZh0zO6c4ayBGVLW2//Wu09
0PnSaHjMKGq5ZrGTOoWbFJOmqU54ZnZmdJrSwqZUeyGfQV8MRq+itw/rHex92F/t
pjfBSOl4PiQiaXeai5xf4Fe3CwIuiewBWVPWQifXXkbP8yvUtl6ViOKr2HUVQIhr
02Pz97MhWXg0D2mLMre1pPsMJbyO9U3peAI9TVB80ylt0ACiLoGhHr3yMXG0WHF3
+9pnRxFbiEgFwdAt/MkEV3CGmfeYvl0E05CZsWraknKB/WemmuaCNkeso+a6VNHu
TDeiwigO3EwB09+nF1AZqdhDbA/xsw2vDUTgcK5IvdkdH09e9pqO1+UvUEKhjot+
mDUXuNAocbXDg8/8NDJUBn4FH24xnCLZwlAvnEHYotWR6GEGb1EMuAVEMJDn5bo4
lfWEo+lITJTCtSUlELM0ixicuigJ11kOdvMpqNjeOiqQiu6HsyUz3UGYKEfx6cnx
lwGHt5J2YMacbGXv80AqqeFNnSX6Ykfoc1KE00UZOZLyHtA9ZWwwgnXCpsTvDHzV
+0P8E8fYjsRy6E6FGVOlBwLDqJuRRCsWkNi1XDHam7z0cnuHILdEZXSLO7pbWotc
w5+W6o56+Vpq7dadUUijNeOgLPb+e/AUvAb5ZnFzlCAJfM4+k0PNmHi6JuFgyv50
wOEWM/Io3vxU4gXPWX/T8rsZ3DyFX+niCsViK65hHVf0z0XXXcY/fSGoM1cwppYY
VgOGXMBqmYwHs9ec3j25gmJ1/7ZhiexSntBPq768pUKXVIctdzRzVTk3jCoE30rA
JWoUio1Cy59+tvhwpOT8PBKeG2cQO5W+WpeQeVHvB6nlUaaaO0Ql/v9bRdurseGS
GJqLInzERIflT0uGW0ZIE4SQpf/t10A59nSOhrL6H23sig59QDFiDZaV+cMjK+2m
qaVmrvvXJN3RyAxv/dNLDPTeN4nqXNhg/RIrPwvGYugGsFQ2vo3z19QRXlE/7C9e
Fk0U00QR1CifsCne+Sc+VmkCKbEjmfn1dYTtuXTL7wkJie5yVo3+yaYio58HcNFQ
j0tvmkfAnp+/jBTMdoRRxzCPl4hLWzL92qaWzNZiwEohIsXb/KQQdKINGwXZMp8K
jp48xeGqPAGmT5Eg5sPLxQhKYUVrmnarxkrTXqVpbG5+Y1tqQKxFj5XtXIas4J2Q
jDPgFyAl8XT5DaGOj7O7bta6fscY1d1SNMYp5LEnYw2C+xHWCny7yTNFKBFQDlWo
8FbDLEzDgNCvszKhjDap5yGApKpyG3BzSoY9kUxrsGbhTddozJpY4cvigzJwysth
fSpiNW9y0Jbwgm4x+xtzZedcJwvh3LED77a35PqfGiNY4TMHUSH/bpz+Vl22GCP4
1lrc/K+z91nAoANGz3zf1ARu0Vh7Rr9P683sDRxnHH6shIvDX1ok5d7Ku4AKx+eC
4jtLgMYtkW1u5p0nV/ACsNG5gZNeX62VePLdQSRqdtNkkGgRiS6VD/ByjyNu8F5l
nf2QrRXlcAIAJkHYRFwH9fmX8qNPBnCGjnGWIxau+EUvIV3FMLi80CWYekq4UVwX
1GFDj0hHKG8qEl3d7ZWD7WfYFYDlEmtMml9BDZWBUOezP4dxVw7dGKZtPVg+TSl1
TbnG39SSx2icx9r5jnxBAH6viy4sm5uidyvI0nJse/b7JqRqFwN6nH4T3UC2pHxI
K+pjKaZSGvFNUW/gUJ1fFg8vjp1t35wAVg2PFwEsPqXRlPuB7X12GhfXleSaQ7LK
5iR5xm6fyv6L9whcIA+PWx0Id8Az9PfBg4onf8mHNaazQcuGtMumjegkRgW7Bild
MeyE97UWnS8OfyV4ABCO5Z2eR78nSFHr3pYlcYW7UDioVze6DvgaXqe6IJrd9yDV
1qGPPKj894hWK+SsJsUh91iv+sCZlGrEHYA6BxiMdttMU3+AD2Phcy0Dmkc6t6Zs
sInxLcfWEAjis3TAd7EyljP1vnfQU7/5RC1+mxQRLNWttD1QocHtYvUAksYWsXn0
M1rmgAX1LXOkHMrk3SPgcUKQRVPUhU38bwfIVO4UxeCkackgwF8zPhPupAwS9ZSh
TyLW85RbD/+3eXWJDizGn3bNpmBDof7ltWhGnhbJh0i928TikaThhN4Rqh8pQwUv
S1GQBf6N+YrBIrsd2Ijh0v5/ljgmWWbJzB+tT4BUul/g2zmLScq9G6ErX2bOqWTI
md+gfmWQ0mf/Mvo7AAhjV/EMKMsIER6D1dqZtJGYhwExfnSLpG2O6BVWmZTbiYD2
JbXOG5xy0+zeLr1VA+f0IV//EIwV7WZOaIKxEUCAFaielU3VDqT2Wjq9sZCDczqx
FG+1/fZZKE944sxcOsSicuJvl1GUkcmSeiEg5sei0yOWugpaR5OOgVn/3PKWhf4I
AMxajjpP7NBNAkrJRjpmlYBaU7fP5YiQk1ow/ARlG6p2g798h+lk6JAdpasRTAlw
iMvxH14/SR0rKtKM8xIWEVrXGHaS80JiDAw+2tPi122lvzcIUVxG+bcK3m/uBPdq
qkQBkmfcqLGDMvgIe1FqdflLdsAMdF9OPc01TTU2ta/mU3w57UvkGB4gTm1FNE5z
cq9cPFtG3qdcaNmeXZ9RCTDgUDKcqxZDpwhFc5LnlLA0o9KwhkxOI5JyGaltUHcF
27lTrw0F1Y1WcSVxByYpjhI0yxPvHSJey50sVIsdmkQ7Vx+dCfD6jRPks25xOPP7
/mKY6p7eTAUA+eNWGrDq29BAvEkYoU+SaNEHrAZprIvQAeCYG2c/+OFtbceH0VAh
dMCv/3YnwxPWX0PRAREjUcBd93P1AX1zPqBrWzBfGsWhdHbPOLp5q3BQOKzc6ihp
wlhYLiJIfsnknU/9iOV10fDpyeZos9f05wY+CqfKWJcVDRsaskuJ+SHbTqRzETNd
F48BUZO/0hTgdftTxoKQYfuxPAmguhlJ/FIJW/rqGMdPxn79rRhYnzySxc5RbemT
wKIsq7Yz1KRMEbLbTKvs5zILntvSGj8RVv41vqITniYt36NeWhLO3KwK9u3YZIOY
wx2mV+m7vLYnzQT20wdJCFM809OT4GxabAHIj44zch0mnRHaw5YX8hM+5nTkh8VU
EAira+5HUt05NxDA1bE9PsioIpvx0bl69tKcwOCZW1es0t2/ljskIGpQK04ecNJX
ARiYVQYpNuIS9Qt3+wW53Ncfj1S9cq4C3ZH7qXPRfl9Sy3DWzALj9LvITYP3AGMF
XizK0NwmcBN2Uw82jR9DTHpFon28AtDdklCm6oX8ulHOP2MZbNwKbIiyqQYmlwoZ
IYtjv3MTbe7HyJhWzFZfSqH16WPH8PCb88QoTlF8pYJZi3hnzeql9BXW9U5rKnri
bxWDhykrJ0lR6VYvmfms6aF2LNz05/xq0YMZVv1hJgwfcKcD51G3RjbYk0midsAz
j6KDLnZV27hpEBzGHiGyv04EliQbBtOnfSnA+w1udCnxoQcuknOS24eQ0P6kQ2o/
tZkJhzt4ZuLy1GLqwp+eOaiMsOZnOErTqiRU5MhcYdiGLclKQZ7ZnP+Eua/O/I+m
SPn9J3gYA8A4e5OybKpiYWtaIktlP2k1oaInLZI83LqwJ6bTsr/H1CchdJP+8WM7
bkGKAj5mCxTlKe6rdsbvglydbkX3wKiPsAYW5o7N9aluSiYTY2iYQ/M3flGIQy7U
lNj1K9V9QkntFcDXpiIbOe5XF9nST/7oxF1hpFu/ZRxH/bTCq1eAYzfIGX911+pl
yTjAdoqnMGxmpgM/9/yve/ueQqTzW6fBL8HAT9B2z1Tlg62PufzubYzSS/Glnftc
UNpZqnC2goPhzR6pF0ZM2zqlNAVUnHzzybUug0LA7jzkc7svpRDaNGHADnTgzJXH
J/eeM63GhBasopUEAA7RMfVpPDbSmezgswxAWld4B2b8On+I1IIT1WUU9Uqf3kbu
1sKIC3iHC+x6+e/oTliVUWvJfkQUghlGofPVNjnzOhfOYtCuuOP2I8jVqB5SVynL
VOUGLjj5ksns2lpxpCO6MTUOa6IAdmTp75XKrqGtJgpdqMTL5xzqs0HG8rAkut7C
Vy7+5+ito7wwekORw67NUEfbwB38S8BU0WdalN+b5rn7ZG7k8RnnmrY9B0QZDt80
Oh6Fed/7yFxKNpMwz0wf4fYb81TmFDxVfE+01kApoqkuFd7G/G3wOaSvnjHtSB65
QFy4MEBfYlo8VlBKsK/rWY5VmnAoLlDWze9CwDyXIkoVaH4iK61Z1ijgzC7JUwvF
/w1ctD/zEyAKzA6TRKK5HBCvURYRB2FxAJXdmNskChyNwptMhE1Vvocj3mVGWKKo
fhcRehFPRslnpvQ4Z324j8LX3bWDV3UBJkOj/mwrHTDf6pSge/0pRw6+Ysti4xmK
aRrMGiuqT9Su0zyV9y/IevY9PPg9zMnvXsjpi/esoNm5wFw4X1AtYP4uJpBED+46
tF75Ra1lrsS+yiFyIOdOo5so3sMhsz2/7b9h5SAtdzicnt/MrCjGvDEViHm71yvx
PDNoUp8VXit/yxsuJ5OcIb6nI2c9PkLoNQ6TwmPrl9dxRj5tn0ZdgXVhUx1CB9hV
9kIvfKI4gT2XtZBuKHx/nFGiY/OynQCbn24kCKx5o8uvMNfnie1TlDGIQR6uqCsd
36ivksUWEp/8IgKjJDyzuaG/AiqcVAV0B/HPtu0nov1Q9z1SjFovzAuZPTgfc1q/
Ukop6K5m9m8DUG9Ck2/xaulYr9QzEaUllUw8xBsSE9gOIgpBxt0m5ms95PSkF+OV
+p/GXaUki7a31SNhEfXn55bGl/zpe7v0LKQ6uWM4jTVrLPyeaxdN5ADTRHPskl8A
GzohB4HIGelNItk4AYh6Jhk88kXWxbhEeA6qQMQbI/iVP8DX0gSSAxesrQEtIlXj
JNozO0AiTeZ6cGNLiVm1i6FaFX9FcMPbpsGwDA0+23cEqPDJdoWoa/W9O3/ifX/C
Qyp+MLrjtlFB9SkRV/6j7u2bbUotwPp1HX4lkZXODX9pzOfiDqvrPCZIl7G1j5Kj
p22HoC0plO4gj3Rv85lXUfsqxlgTs4yycC61toG0H02cDm3eT5I46nsKsxyP9Vez
gOI9/vDq4m++Nom3i1T/O/OJ+C3Y9il0EHjq29vsegM5mcpL2Nqh9K67V89qjfX8
LwcbQjWBx478Ubm4WW1V6Fe7I0lVR4uabTkdRDoaiHEAwImSBxcORQ78D3ulW1ZH
BoI1euFKtLmAc5LM2bViKGL0jVNvGUYWeEhv4ju9/va/xRQOQpTNlof4RYVzMTci
rIcVPTI+BVGZ8cgxmqFSLJxCrmGH4x3EQ8da8RKkGl4jPw+sASOtmoCGOtNZ4W6D
4Q0AjduDCrDCxMQfquY8dfr1GKbvt6Mg8HYvAfnJ/4whe8upYjjKnIt1QTD0y1IJ
R6JUUiJ5qEltZaxUSY9AnI0YdhvWo0+pJTW5wq3H6qs/nraZwLljZ1ZFaQoT+PSE
RichUzpfZwPRJxe+v9WXbUbVkuK7ASxqWE50QIDI/Xbj4NW56LAaXwhxYUAIomUp
34YiwjoI9yWY/SKNTfcK//GWKZUnkrxc1MXx+aYEA1MtEiOufQdqdzqsIWbZEbsO
GsulUmdhClkphzXap4wGckQsrU+F07mUdGwXyhnBqNSVX2+kfo60+erWyS0FLu+q
gbotwSZlnTTaBhYMdgMCISBBpPbQQxsWUnlJPuAn/0he/ixShVxC/Xs74QfageED
YaM/1O+JxeJoNVnJ/NWA914SYOhnlxCdJKr4eSD4dpNNpNq5+p8x19qA43nHeQ4J
7yTYmeAdv8Ycp1gjLQ6U8YOUJT22yobsBtMSrTFRhlm2aq6qJIZGaQzUOmaCiQMN
Be/1lf59h8zFVKu9fl8a5LDOEUpt3slfAgppNV8fe7Vb2vqoQxMQdHc+BAbbxy1L
BG6qNVqu5XNrHsLmcpMIIgoG5G/dVVGLss4THXWI13SbdSpXN6rsH0v1iO1xffBl
Jz9TlQYbQwMXf0Coj59zROFVlOE3mniQVjQ8LLFqSLQf1AnHwrZoSFa58rf75e16
whYE4Vy7XYhWx+A92ZW9kRyK2IEKENjW0twHUtbuzyQgWgcTbpCCgnVOH5Fj6zVV
BC287tuu7fiI7SHaZtuf0yTpwNfrAYB89dfzaRlycC/8Sd7d6sld9d13IIdAx5Ab
dAMYgsSs6W4roJ5bVip6S4HKXibALSpE5wO+z6ooD2PD9RxbhqoScY6A96HbgaXn
WXFshg3Ep4x28ZjVzYwYVQy+JTkLoFsjbmAw604AO2RQMJuKgIzn1kKImQRLDkTJ
If/IdSeOV3d3Kmjr52vHmtmkLuEvEbyN0s5+Do/R/wR1SEqzCJJraj/BkRcv7BdI
tNNa/exgX1bK8MxN6ugc5G1hYLt//YfnfaxMAspeQCu/ZXuwaFDyD3/wtLenCLtM
phLWvXvTxso73zJCdx4st0rXhQ+Y+dfrEAQTfG7bqYhNNeY5zVeEZ7FbtLxAUE5t
lQC3c6rFfUGGnBbVgWLwtXa1XRaTuf0KpdDYJVfAsh3PkdzaDdYv51wHMdaw4aoF
J4aDx+hWd9Xr8b/wjddcGY2ENV6LtPDEFxOSlF4N5gN7UIkF48W9DdRbbBZzczT6
t972kYtOmpeVhpzsyW9A/2+td/SYaFkVwF9gBlX16Z24nuwnME7yvHnsLmadeey5
UyTI5IyI8GtXp8tqdXrKUm5wsIo1VtZzfE3peW0VOkQKXHvyWo2QBWWTLkss8bky
G1PJFlgjk3hh5sPEH714x2CLP61mR4erzdqnswtb+Bfg0vMebjBKIjpaprh3AnJF
aEWnJ6BsQ8dtX1n8bBlJ82r+FctQ2zqFmBwVc+MfQmxsAfaZZrjg6/Ol8eJrJq4r
Zhc7JBW2U0iLQc+xVmuCXOWd13q+YtVDu3vdeK7+0y5OGg65Gfj+diIR99BmCvky
oVOh9InB2Ccu7rJX+A2yzDY7utAYzMydGfFk0v5IE0fL4UShzaPvddZNWBC0lrLX
xzyXg3bhkwwst7t+lL5hZb8jS//noZDSXYUZT+YrfS4X0BDgSYdtcLUw2OaZLChc
MiIXCsdPOS+YFJWOCAmB7u7ICNP4cY33QkMt9eUkMQaNnOGq38BYMerfDXpR2RqS
c+KLXs5nfHOe6jCxguFlDv3thaNopqPo+JACHsiXWiNF2k4CylSXRttg4ZaVHQNi
DhXaEPtm2Bhv5J1w0Qwbc2uGb3weGTgdZ+btIKSMISMU5i5KxI1TJfiCy+cT4cH+
7wDwNV2k+ZNbltLIlH4ZIVGC24FeQ20VKeAehCXJLEIKxk9+LAyIaMs33BBEft0g
zdCOK+U0wpxusdhHC3wTWgzeQ7ef/vSv3Vl0yj5YR7HOELXD7hp0Z9akFK1QnX/A
g36B8MEcluM+c/wcp364XXMPHiuRg165Tck3jq2I+3c87om+M8DBDtZAthRbFNYz
hhpjL/x3+tUQlN/q8PH/X2yjnfM7LSh1M5bud3qDdfpUaQD6pd7FwNXBnV/ct53V
nRqnzjIXy5h959NRi3Vkkld6mIhE/O2gWpH0phDAm3Qr4COAPrQSZ9R/KjxxHHux
UUiFpdkX2+ftsQlZeKivo5beSm88s/xMzAMRq7IBdQpsW4d+PkmrDJfd3p8/3aqq
w1yzARBPN6VwMWRtBwqBkkDLysQVKcPiBuFJy28xkc3WOScJPa1CkmETyHmCdPHM
9L2iWcqVXBahQtMyW8cRy+ziqHR/nIFra0zgSA6Kd6Kg0x1dxnKEzplXVdT3ktyo
kkYcrFZmtrdz870EBqmWOUV05ZGNKDBGHhKbNILPHK9Un+3hgXK2HRclegBR6p/J
kM9qYSVtyos4EkydSlU6tgQGPcL5OooJevHTiwR8a7rbx7r/zslMVloT0VvtoIIu
+sYLoQhHE/fuRPZDc4A6gtWHwD8u69kiVp8QOUng20ZzECc9Pl97o0LTo6ljUfmp
YNnJWx9oKjHQgy0eTqGDTz5UepLBRRhYgu2JktMMJODnEk/NNP5a4xasCzvArwD8
Zy5WwMiIKqYkrQB82zAUXyGzNDEyDZM5G0DgjK7dKuXhJFg8xfnDknCH0173qjBI
TvN3TuaoKaSZeK+Cz+m9Mf6z1GB1xf8jnYw85iHPVDri1/Nui4ST6Ai54tUhSCqF
3VqJusB3dJ7p+bbz1smBp7qbvD8YuZ2RTPUkCRuARdyIM0EXsSOc8TYvwV//Z+c4
ToNFsrr8Co8jq5DvG6yWETKSnhvQdWHT+TIrypQ5AcYGv7v/G5k12yMJMzeZjfMi
Xh4Lop03VE2MACbmllFZVBsI/xY81zucu67igphSKvjxsleUT/zi90zrUcIjm4WW
jr3698/j1dQ/qGbuA8A0uQv5ProNE1r+ZmtTyrA4yEurGp+nxU8kCv3GM4GvcP3R
gwcJsuIjv17QVu8g4IW1T2lk7zl48Zmu2wznnODdb35HQDLDb4fwiSpZfpW6IaQq
o8I/Qtdu2IvYmx5jVof06PaFmuIGJUgF6J20e5Q5Wz35rpIiKEtyrnbRF0Bv1oMZ
ULISDLtk1d0HA8Owsr5tZjlej/9hakaDUIj6+lytlAY9bNFKyqxLkpwEwIMPYqog
YFpjKZCGRJWb7KV1maGcDV25chNXzSlHRtCWsQinNN58lsiH66aKMnGAMjbr4zj7
D43Qje2kdP8r4dxHLabAL4bySx7UFyDnHvGRnkdwLQOBxF5+2P2cAwLyUSZRkiet
8Xv0bwVQqXHHhnJPdhQvu4ZAyvM0KYOPsuGlELBqvDVbLAxJuRFio85yvSXGwV7Y
ETD+W6RKErkigd77kf+EzjiCWp08EHCgr4sIcjTp+/EfTt5XwHNmoK9Qh+4WEiof
B4HSOmbXWMErwcWJFQkbAxROYREWPjzb58WdgMvSrq90gTr1toybmgEkEXUDOgUE
kidI/ZEyTV70yFEuLU6uoppy9n5TUDdHFxCxvqj1pdZxlSF0EwXoY9hRjGiSpfkO
1xhwLApYHEAa8hsRNA/LG6Tn5DiUtTJckrJ6njQMXeC2+NWFI4QJ0573XxgL0465
MYkRxIy+kUFipOXCaD8ev/bQVlBZktjKcnEiQrSupwSAl7Cmj4ZKZMMfP/wytLAp
ExYk2l1KCaJAEbXrcPwOo4cf5k0F1HLPTgnIsQ819hldTU0iQtfnzKv+R1TNYjeh
7lGgcG48gVHz9kaBUxTeARRTv6PoYVkNVToDv2sJuBRcWGKhdVdj/b0i1zmPGJd6
V1NfYOrym7519NieiUXYjyY430RDjeoZT9kJWoewCt+DKh7DEK6HBOdrpcULTp7A
6pA1kbrH9QCnaejl1xanmE1lj6XFdTLLTqkgFB07pLihpxgFfBs1jkh/46UegPPJ
VgdiECA7wnhoMfkKNNEN4NO82AWMMBdhmVZwVv4UZWsGKsjNBsCBHgoPGHzhMtP8
tQWSzqXaJ9gtKETOuiaOIAKLGQ81D2cNV/22MD0jjWUHESyuQoX56IGyimDpyLKf
nA5v2xatkZOgjY+8Fg+IJszIzvFU1eDXdlBiIJRT/1AfkmJTm53LYJc160cJdbzR
vKULhOoxZ7c+w73pUTut0Fh2W1Zplt809eh2a5sTdDFBEj1pGVykwGa0g0ZNm+PI
r8Muj8heJRpdjB0Wp1A3C3InFuu/GA39daefMPLl9ldGCiqSGocHsd9iqZQfxHka
DTmawUjfwWR0LZ3YDOMNLC+PDJwl5w3HUZeNox3jehbquwDpL5waWSC24m4A3f00
KSRz+IYU+iBATgETzXYjIS6t4q2nc9YVCYpiIEUMs7Junq09JgmdIOMyLvwbx7jO
Fnc+3HR/f8kch6jmwAZkGZ3RYFYmPIYx5KsFGORXdgm3wg1tlLaThkElxck/PuFl
3h+w586/Z6xdNVbYp9MgQVloulqHDixnN5WRq+iApOvh2+FtxMWGmMcq+DYMQ3cP
PVkv9JPHSTaP7DBdRQK2fTBHcvm7sUrWdex3LPPRnUHsv1iEWjgGH9iD3rN5pSuU
dV0trQC1H7tDDaBTm8xaTR6Koc7FT5B0eGJxQWnEvktCvQ9xivNL4FpIOoR+dvY/
PoUMK8UvrXGnQeOwp4akPiruSFxLuq7NHfXtmGhUqjIK6NOOUlSiaK85aSDFGjh0
4Hl78UBJs9/KCRtrzITzdLmSOvDJyd4zksfWwmBRL5NZxx+AV3SBJlhRINg9Ni5m
VCjXRMvxpQXYO6u+QxNWpDDuJxgFwwufl8Lzrkfj3JLNxeFhnsNyLHaWFRZudrvP
tFBXJ9FMdhXbR7L1JPdimN1j1Ho9wzSHvMIdlCROFAD/RYPQQEPDGzGQjumU9hDq
ia1PQj1mtPOUcUJapvYx7v2/VD0RQPTrktrHHvNQcVNoWgnrtBsP7LXVugWLtgYl
hVRNss4TJTEph6xoIDtin8Wq8xznWE3wkDGxRrQsdX/zFCWuqlxralWuNTsSTqhA
Qjs1qg0f+aEkRy0sHTQmDOsa+pGo3LjKZGQo/4CIjEjU+fkN2Zs2/XsA8dFR4l1C
R0HULISsu+rKUlsTrS+9ipEAGbWXfniri4BlqhJZpLLTxTx34R9KBCuDk1I7ur8w
npdMxq/dOsQToaqOTWI+r/z3Y6xoWPBA638KSnXmLu7xB0dGdefxngHVN7Q2Q1t5
LW9Ork1ITO59ECj8YtWSB2VFepljkK87ehrCAVAhC2waXUlAIDf9TijgFV+CRZ1B
94lzM8pMh7whk20RsEzvO8Tahg3TafFbZwYiTEsZpMXGKq8zV12HQ6vfD4tV/ewl
+gH3GUIjVn1KwKyn67apMehn7zaZy9otjrqCGbpGP2J+EW/V0vQekFOYGCmqtH29
RnTxLL/N43nUHjgF9aG7sbGaJjNBGP1Szknl3zbWElcrGV9VEXG5RzxWUiE1xMEr
FjFd51/QucJUBcghg3I6C9Sb2W5mGCcfsxJRkTLqXD74ocgr5QHF6E0BzHcLycXK
mfUDMlU2GCXd9jBdBLxgDnTMVo6Uf6RBMgL9ovt9IvZeHDtjJLbJf6pDmeU3Dgkv
66CRmXFeIKlCYdeA+L6ZVfaK1tDMzd44+y/uvmgPzNCiVtlJCW2gbIdvphKawHyW
jZpttX1/YI9/lZYYRC5hFLTxglEThChCGAezsiXRPLGdHIfflc/BUwt5kSaNSSBm
dmnIaFNyeLongQ5PylFVxUrwUZe+IwDZtt7H0X4JJDJaTvJfToJMHuYf6e1zoTMH
hSRWRwgWYlYUvOgEhXWxUwsKzZtMrvABbqe0LDzNctkzqU7C+27Bs2W2u6p0QBsV
P+IUb3xL754u4n3beuvZMUcxBpt6W2hOi3d25LWAuQO1xPjSZMgidemex3v2QOwK
MEAepZDnGXV1nZdnLbqz7i+HIbFcr6hJJyMmsIFUG6TLoSdTZoW5l9X7niy4ZMfC
c0Z7NRubCvSPPw4O8CuEPeakS7Q+wLbtvw2UGW6p464YXCTYJ5lhKJfD6lt9uRG2
p/X5TXHmvPzxTI4f/IF+ah0yjuM6JLHpBbbUw+rUfDxnoDdrOv3PQ63SpiPwU3Rj
gHsGxKKYV7bDIxmGsC8VEbVz1exGd3H9JsaC2pNZ6QlhSldvOou1ihegBtMN+g6c
G6sp/11y8/KS3XfF6jAXvnq86BO2NeauU05atVrAWNC7fzmcVIcmoFlGx1T9Ex4p
nA5oYHnMTXSnXZY5vu2UxHQGwh4lib/9yTEwFTNm6llawcqc8l2SDiMH6GUdXk08
Qs4YxEMJYWBka8YqYnW+xqhF/+jGqWZ1pPU35VnkZ9ByjrU88ftV5sqtACJaf8xv
G8uBEqa1hGhO9mb1cYPTS/ahKO2xTnbdDxuCrhe/yk5ITvYkPuLGXvIuMVCIQWiZ
mv2me3IiUKw4xO4Vlcy+dYwxYwwwpva7A+44zF5C43kHHX99iBxm+YiQ1j1/RU1b
iN8gp5XFtv1z1A3co/nHsW0lY/ZwRRL2ViziZDidPnuqXI9UJVrMpJCYUthCJutp
cLvUaglOexcsp0jwccvnTtcWgY6q7+5NnfcJ0QFo8xKRYraBPc5fAO0bCmY9eAEj
sF4XRhkurV0w3VoyMXBkJf5jLnValz4vNeIeA/pG+QCEk/i5Ej6YT17XSW1PSUg6
z+g96HIXdntYFFK4vZVytKA/s7LWhn07L4hsx4B+EQVj6BmY7YLMLVjVcX1MzYRL
tL3hzWyNyRnlihcb8QugfZvbhXUkgG/XDHgIY4DjzlgKyCZopBv3nWx13gn7u9hP
/GOOpzdwz6GwL6B6J8UArKT3uOhS363oQfS8FFZ+a3ZOKSt+P2IRC6QGUH7abJzt
OvLpQjsitPK+oNr2CB8bCwiVZ3OW89DFjX1UI3+piOB4k+27/0XWDLW+8JTrW5vq
96VqBzI21zB0szqYGlAKxCTubTDewBvjxBDh5Kimrpx+qRg53OHklVv5P3P67SJh
mt6fwzUULhilQHjOHKzpwIF8ZHC1KxW8xvj7ODEYF8glTXSsGmi+sqs06W+dM5Rn
K15kEBGh4fCppnz0JIzCWAUkKYchcjkMlWdz2CtRDR77pFzDV6DjxDXxsFfHqgTc
nN9eTi2yQRC2U5irJpNo+QEcfKoiIQGKisSfFE2jK0upwVJpgyv0gOAKcdrCLLoz
T5xDeRmlCiIXbcCQg8rEYkq4UgS+TySwPtv3cLWwI78+jk2bbpKdsppgPdHzuEYh
rE4QkmA4LsqdvwdlMQVNqmMAQAsb0/CrvMHUY3XVvxjsu/4mSKMBgAOrZlvycVqs
j7VWL0XoAEfdpll4Fk9svRZZtu3dmTX3mSxdqGfFrgR/8/GwCtCYGWZq7fnefxr3
iDImdYhhTThx9qEK2pnkG2b6CrCT/DGnfzoxDvFZcN2LmSDlhPcKIQa5EdxgTj5f
cTzlxSe+hhjqHt2HPFYjgOjsxfrL94oCHfbxtqOI6nJ0VjGWw/KP19lOzzdsHk6H
0OsY+MYlwzUc1elWzXdjf0cjwJhNDwg1jNlfYPiUMGi74BSfGoxlpiCs3DCqA58a
MH0/GKodIm9IKg1QX6LtHkosfhUzPqRLKGXD/i59h5azJgnwEX+xKlOWTf/AeMty
Cv50jQlBQJD7Ky7OCqm5K8f8sMeYTYzcCiIYoiNcXs6uL6oE1pquvJXf67KkKm8+
G0VKLTuLWrPxptbPezVrKWd6556Ioqa1ewCmV4FBu9K6STmsDi+o3xLrw3zaYEXU
q1CdZJUKA0/t8hPC3nCRHrzR3hVP5W2pNIiFkOfdrGeswyh11l9U1xmLMGkkKGJE
kmBACX16e6r3pAtzCc0AXHg1AJ0XCbpFn03mbGx3qAcfhgX1pGuZ35iuzSh++qe9
cGQJgpy9WXf1Lgd2MMfrHGVwd7c54oFeRFdDwuxZ++j23RkhDzvXhYffgONv7NXo
sma2F/nD79XKhPLqprHjoHLrJLHIJ/E+GsT++OdjRmZV9jA4y06GRtw9OmyWe70a
v17leLspjc4Bpj0K0MGRaiaNfm04/IWBTV3idEmUrw4/g/2/zlTaTP1mAJGoLgk/
GzMmfSNd8on8pnHa/xHQ4voNkexNmibAothzA6WpvXo4ha8rE4CjCuL0CkTngPJF
PCIfmUfbZOHVyAdpM0YRKEBCJf44FF5MKNGCm9NXT5ZozX598SlSiKF79LA9nnia
3sWBg2AzY6/gCVw0TF1uvGsY7xvfM4iXrntWfLUXznFMiIsW/Kl1yHxXGMa8DcjU
PN9qBX26UqIm/A3CFg5x0xGU3ZSlZHMhYqxN5vW/qo3tOrP4gvF3IB/ij7MAkPYo
5pfkB6i7iwSWcOtcEHZSyenSaJv5G970+PlyFqVZCxJ99zUU9FBJ//u3pGsLznFo
oRGKDa2JTqCyeWGCD5ij8MnV//KOi4x4DoJnAxD2hHd/u/XTqk7ltgXgpPR/4fAA
1KKwvznUfHiIeZUFJXv9fgsOOhbEK4p/evcOt7uRhfs9s81dDZrZ6kK7UUU6SYOo
RAnZFU3KHBTFVM2j4CIMIpeQFCiLDeY4Xfd0qYG67A2DSV1+Zv5FofG9y6jXGYvf
g0/NOWjvKl2K/W7afdd0DF+aDsdVsV9B60pyI7EIouQXS4rpk9Vzpp5eUCUqmtWT
loM+QL9YS7T8JuEY3ENRc73F+I+xVIUWT6YwLyp5MBkE3SMDIgNbvavEUE0kRMuD
8QdgWxRAQUEPGG4JNO3lxpVY5NMvxmKW+QRSekU5H/bscM15mEbM/fyOcAiJaqKX
RWhoFsIsT8zSNhvgnNRNxvtBLQ8fZA2nEwGNvCDd8WEpX/UiNtF8K30LCCThTd0N
LLVZbViQb8hCy9whFwfahmszGjIfdayyhxW9NNXdEavG+Y58P1b1DdlaMqR/zab0
8lSJN9b/aPDiBPiDKwpGiaxXJ1BX3wgvis+AVaajZO0nObf0VkFHs6hAe6flXWGe
Sww9bDewdaOWhx6jgnxmmy8LV2uaoFdjKmVpeaEtHaYiHx62gaTV3V9g1AKhNZxz
eQG5dT8IoAF2STli9hqslwPznRjXCcowUpdpMZlvQAvio7cUtKJJekRUdLhF8rji
LaXXaxJhuLpACLfUNrjRRxh1ue9dEfhuyJx0mjXu8DoesNHoOHTN+YxOtiEWBHU5
T6XCzdd/S7uI9qRfTlA98Ap4rOz3BtN6n7iiibalwmrT04Mv5ESz+y+6C+vT/2AI
A4/V9idpYbxLQgDDDS41MO/cGtsPZZ9Jrha7KNQE/po/gaS/ejMEC75nHdDZet3A
9Yg3ZXf3YJ7P/ED3azx5flUXWPc9emvTJ5BIe/No7VU67V9kxfg1iysC0rq8+0ON
hvakn7tveBQA22mkxiaETRhn9LZDjXskSdFth+eQZnJtwjvcHD+IDEXb7/lhGt7w
E0BVmKPOeDkvifkKY+Aspvw2ZmNaaGfCX2vNAMQQfZKfT3v7Qjb+awoca9tXX8hC
9+TOuQ2P41JXNgn8MBSdjDK7WNkwFGCJrzd+LcPjGQjGqgWYSKfGWjFI6HZCZZeA
WbJFsmnxC49X7B50FUxpMEXlO/QKeMKcD3qXZ4GvSSguabSELIXa0DzMUqv0Aihf
MjMVN0aYIFMkb3GJ9uh3JjtZpvoPKgnVbrAMHHAaKD88sK6rk8UIRVJkrPzFicpQ
/mib3jNOENh2vhhGVCr13hs9EjEf8kMS+MLQIaEWiuoM/bliCjhwFzefMGEJP1tf
RcAPIGvgV9E/sKQC5iqOTiKwEKapF1s3ozQxlGUYhXA4YBdOSdu5G2ZoU+9RHDth
eErSifNBPuKQEMeGOlDq0uXdCdPHJmw4JnVJzE3tW3SGsdl4bNZPfO8ydD+8TQGq
Iwfxfj7xhWi4DcY20/YrCWtU7HhzfMavKmAAWG9MnpjXIMif4uMe7r7w/mw4LIFr
mfOcYFMlPAaJ7etm3M4HXlY7iJuW8wZ3xwyZ1r62mBExGRkydbSCTcnvesjI9/po
ehZILlcRyFT6rGqM+AjqRwzeQ6+2jnxtOR1jikdsTxqpptBMeeLh6sYY6BFT7cl2
M/8meDZuEeCXhdCdS55yxc/mx8gcIqqbTgcGW/zzcjCG8M7/pGFfBjOiBXwR11ps
paxbXPuRSS/2MnwSAgtxMNoGXefM09xxsj80MzOhYDJumg7/HGsl+cPh6s4XSv57
z5XM3VRLIFcA2HR9WfywRP84YVE6RnUCUrZR4FZuMHW4/nJpVyw89GtKVx+GGp9b
FSylRqslgqdIMGDzUMq2BAODwBJuk27+URLbnv2Cf3FrknNJt7G2AtNJjG/n8Zga
FapeoTt9ra0+EH+Ve4e2JwhmFAdi+9eSx5R8nAGV09hbnIgaJp+FJ8xtXkeYYn7g
0yXjtBx2x/wDBWrQnufzuYktKFl/U2jwMJDmLEYJiSFnStFjHOlRQISBsdiqS2Z8
T0TRi2c8hai0OR7oQ3/3QocM5WbTqh+Y0Ff5SWXxaQyud2edyRYPHD/rIFnK44Oc
UxQcC4HvBvlNyZ625TwGTIuKzNEDu9RzNGaBvp2KoHEWCwGYa5BH4k8AeI08VJAC
FRouAvZQxdO3XooQn1pr6mEBOBMzWK16hvJFlklLCJj555UtT1+eCh/R+k77tXG2
s2kAkyz3LgzJ5mapeVVdSRbn3xnJR6KGB4wdasoleOPyOtY91tD67tlou0MVm5Pm
CD74v4W6KcLIKynPGPR5LGRklcTDQ0S1OENsKETVZP15Sew7fWkhHSWfszEhWjm6
puwlPLPul4sl9VQiGtlqVG1D1WITVSqiRW7sHjd9+D98lErQn20wYbNjcdHTdk5w
h9BvT6eBupnMwNeOA1nRS1yEl9gRzf+GvJnxvLMjm1jvcfTO6op50hifA3haTH3f
9M/YtvKxRJ64plUJPH2xvc/Y3Q8RKnFvDooqjEsWmI7MhIFbVuLw/b9CWeSyxXwm
C9sfwXnGoMNSMePB+GqxATyYVRRMNJ6yvGp52nkLGATsSFqqQ2nsF7HdQzTG/ykL
0cPtzzTX4frOKu+xQrO7DubXpzFFtiX+Ivd36K9vnJTMm+7f8AS/c6NmOYThjCKl
PE1Ke1d3nY5d5zYZt1/hmr/LRo1BaFQ+D5tvPvDhPTLVthHFpuTA86sd6PpZDjXy
NQqbme8ig5aC3dbVHqaC+uAh0xW+vaOdcrARBLVBOJLHFMWiRGeDtoulw8GxjsKo
M7S7hP9xx27eZ5CaEiWVpM2ks3kDopjgl4CBcN6nCGr3LOZrHytqQlOIk1OPfZry
51ZBEn4lmh04o70Dz8SpJX+tvxy70APctFYZ2cKGMq+EpizUd0isvj1uU/Isfot/
aEHrsMkf/bMoICMmVXRfaiWaTu5Cx3lPOeNT1Vv86f1WZQW0hAQlFlP3W5xyy3VA
ZcNLvdk5Tc37KbA3i8H+Rm8GlhF+UIk9lLdLkELuTP+frYpZTxzgv7gI0W3cF3ln
mbsVg3pJDO27TfKs8Skf0WTZ8eMCzWZVxtxaSocjNwG7xzEwSpFf3WjlFddXBGkB
XoCUJPUSENvo5aMy/T98RJD4FWg76BnLabK71YXgIvwzwJgSKoXh4qLy4g+Z24hG
dMFAgz68NW6Zrr7k57o+jcmO01Hbn6SSajtMGwran4km48ESAei0/z6fEbzYlJK4
HxYTtj1M7T8RpprvonLPX929AQdoE9vp54yH3MEzv0itkUg75G91ZlQGdAZ6dqlU
BCozm3MDcTSzjTezIAM5w7J9ZLJRTW+RVckbAW6FfOmzRJPiYHwR6L4FlH2+ujTC
QQDw2CCg4WK8U0giSfWlMxXmR+asH7cviZsL+2KKXad4gNaqZswdW9KAfFel+7Yr
JPcliRTLaWNPYey7CxOEGSOta724sSyXaaH6QU7HbSZp6TcDWk2Z2DzDPWCEx8Fn
L21d0pDGSj45n3nAo6yz5/RVridyYz+h4yEYhA9U7AGIKkJH88UYYfwahHw14/i0
mSyqMlN+Opr77Mpzp+/lG8k7GcSRifoqz2WkbqF4uYO5YAImanF+r+0Qucx0nFab
yS8OLnwJE4VUwwr5l3CnUDo1Sa4GHfoZTW7SkERyOvBXBD3DUshzqXZgSqBjYRj1
AVbxB2D9ttqhPKGWVaaSIad2c/5bB3IItZMUUZwHdKKUdk5yaaVv1+4P1+mYFO0Z
J5PVbTgcGCV1hlQBVgzrNGEASj64JJNQ00saV9vOo2fe6XRWDIu3COfFqErs6wYj
BjrxYLG7DX7lky6bCan0K2c4izbOow+Eo8E8g0d9V5ACFlxjDcnl1Fw6ooxYr4Br
OUT7aKrPCCM+NpgZD4eJsFwJkNuiStzWRnYQ8iVf57vfGDBrceLr/k2rCspVUOoT
QMRa2ubwTOf3HPJYx6doAm9kRAmtI4fImbyNHQm+Z1z5efiXBM18R7KKEM5ctIZW
54Ci6094E03A2vwwp2q2n8pehtKwoUrH5zXnVPW66PufDN51E9jtlpqXv4G4/o6Z
xS/Z6Izs3MLpLtqeK68463fGy/YL7LbC/NfSeBKFnV6glC+Fk04lpTlNRhlUWAq0
vSIelW8YWNWj46oNjKtpKOd9NpBgvsJk3vRo2jj/qLxuvSzojs28zgJHNZmX8nWq
36OjURRCtYF1p4+RziJoPE9Ze5axObVKlV9Ae5Z1EKU8E3XTpKqra95JRn8kEdWL
WYvHpl4ELP5tqf09pyggzD7a6Eo8hrsSPshyYu7mvnAaUOwO89XWWLqR4dG997Vj
SfrmhjbNnKKLZct61vGbwT1RnmIpRERzcphOPeU0rX7XowqzBjjU28E5UJAcesXm
a5r9rKvulc1/VV3ZJqV4rdT2LrwMusEOZY/EUBUSIN4DMO55YSva9vpT0S8cogDR
cqzsB4lVXNsMsfbmyvcN+QU9u+Wa8tEDDiuO5YeuAxT4cXXy+bCNekuzueCO6Yq6
nVzMxBP0GHsj4ujruHub9prfa/He35sdSwvaLzsYht2PaR08wgrhDwZYswGFi/Ju
DF2pp647ReBMLoEtZjU8/T0U1BXTEC3z6+EG1+b2n/UhWwr6DjJ+1m5nvYV7K/0m
cE/qmx/Qh+u54Plko/J330+MX4Z4e6L9jUViZaLly40iIlFgdzTv+kyXCkm/VkTf
9wzHz9moFvgoHm/HuBFJ3BGpogqpN21fGLkuh0DY9AtCy0b22mWuCh+Drp4Bm1G3
PsCevwpN7gHewAsMA8XzXBlhbYm+RviOr4OgBChKhqjvESuRf13xkfk+rlAi4vyR
ZaVXdqL2p3yxfIP533/3xxFs86SBFWOD2LE9NQhlxwyr2tiY8IGCAjvHOUBXJ2xw
rmunaMMI3Fvt7bwmBZlgUC3HwisA+pRVLDA8Smxtz13pOceG3XvYexTFquLhwKy4
9N6AxmE7pCnuUaYFI0KxIbdFyYcE+VYqQM+1gl/fLh9CBiODPi65Zgow4aSEFF3U
1I4cyAGZXHmjSKvF7JCzm50iBYu2nhoj9rjmMvRfw2pBgoUdnwJiRpfHnfUPKAGi
ZkmNhcD1Z+pU4m+gpX+S+4se2E1Rmj0FDlS5T9nBcDE1QuLI5Rt+1zi7gCJF+xRx
liIkQSgzG4GB4o7eoiD3NEdX2bqzeR76p/czCZK2lTXaCH749j9csW+WgUiD5Foh
UyNrBcxww21aMPcG6QE8PZwOfOEt2vr+vxTsusVL6oEjOT9YENEoJRYAxI5SDCyY
aexqH8wEcVaE8HCO9XPvoTaeph7XG5xg5cywna0rz5tpEaa15syWx4F8xORiAdCQ
lIOSPl/9EPcjm2MA8jZlPbUXMyLpQVhIL7oKhP2zMkTc2QnjmPf1t1Lht/QkdqNf
cgcoY7rF86ocjxF2DBcLpdSnuPGNWZJ62r8P3SmukpJibAbrzp+fPSfO195QXJvm
QvzMtYtGt4tYGOW8FTa/e9WzkXGkbiDVZGMJgmy2KL9GYz6+rdOcSzzhRRUPRaCh
KIpnvADFbb2gQfR7apSq7CSXvmRFwuRhauTkXfA+D3bOYRMkc+YBndrEjFg+79AQ
JfjBJ8N+Xqdhwx+ikCSlqRUmkpFY3vVvbkU8/09zWfb7QlnWckDrbw5ITsMdTQGB
BeKCWe6AeWC8HziLT8/4BuM1JfoL+9H4UAkygcNAfi84A/BGxsbC3ZnXKvwOrUW4
xwt2YE4XOsLrfODtO9N4ZDfRdJGmk4VNQh8IJjy6Fe5OnQstVO9m3itYgVVm86fZ
D3huXPC6jWXWIhzO0IOjI8mgXGQpvTajo1jca25JchwCEejtFPU3NWdO+sIrf6AO
J8rmgKAO1/ECWvYWauORX/6c4n1vVzNtNHyyxAEF+HbL3k41W56lSrd2WeuQqD6g
Z/yogQEz4oh4I9nP9K7qUHp1LeWuJmPocl3qcGXzAoYQ7XeUMBBqCBufV9jyKTwD
aw2m2OWZoprFo3avRwjHTl6ZrI4e6idGsyJmnUjEJ0Pw8KD+fGsTiq5MoJfvFGov
Vt4vt7OXZOSESnlx1rVHBoYVL3hLwzrJ5R7xWykJpbU+CHOd0EeQEW8BEfCea6ro
uux+nAJNP28Ce7YVqaddgroJP7q1nhafMExV5MuU5sbFSUUcBhHBNv/fIuknsgh7
6O0sUDpHWH2QU+a4rcncsvXH7DgHgzfox5RV3bPj4msWp51vTZ6iqc582DleWAms
M82nd/HptfKfFVcWwV8OVfSEvyAu30EwbFMeYfGorG2sCQqAeM5olYfuteNJEvVD
qvKtaKqGXcf7GlkV1Bvggy8O9R4gkpdeEKl0qwR4KhXHXyxq9bBzoVXyXdLsM359
WmsksB521zuByOeHlKJgD7NXhzy0J1EXaqGk7BOUc3nFchoK9vvNVmfe+Fi5YC+N
Xj7cCfXlfiwk3bSeyIAW4Na2T2A2+4uvunxGJGT3pGL+fUsvczMEBHr93mAnipaR
cz16I/C2U23HxCO3K4dpLfGXhsG98t5iW8VP6h0lg/1BEyytLZOtsqBL/Pw+hSAC
1HXQb2eMB7Ar1db8IZOlTtpn89ROCRACFZQGsMMhpZXl2voQumoCAMej5I0VSWJw
Lr39uoaZUD2+5Rd8j4VzNGrATOPj8Sg98jIDqGpp6y64fsR8K6JvcUiUJYzMfjMC
eD5bo03o+qh6MMU8aYyQAfVvRtJhBeIDWEIzTzpWFk+U1cc1aG5hp0cgvxJaw2Id
RNQD6EfqOqmQeTvOqJAKri/OpZrbPdcpmsjQ8V72Y9YTu/3fsi+RGt+vSWbYBHbZ
wA/p/vDOnIw/tAExycBp4P/qEeTtMmvK/gK+ADLmrQ2cBVR+GHOFQsTvKA/OSC7q
VsbOrQleQjtqILdAIjOgIgDJP3xkFRLj0oTdOUn9q9lAa//xHDd9NRVNqnUX+Bvb
E3TWHCtf9uQVRk+BOcI2izjRsNR0+bCaJUGX9sE6w3W61sMv/9XIE2nH94tWGBhD
ULbVvQJPgiivMyf1wIKRYI+4pTkJ9JeAHB+ZF34z5THKjwg38HiG4uDRsrAbGFu3
lZ9tDmISnb9gaoHnvN7VuEaQvVFFlh5o99sKnFbxvPnneS1e/4e/KuW3w0GbyNnJ
F3ZAeIIBe8/zWa1G3EYUq8fdriuoOAN6qzCn5ZJlKtHrgKDcgelE0y+6oS8Fo8Br
QbuT60nm1MjOnbpfBLTpkbNR181OmcIEqPLbamzHFA0tYOnCGW4akMKA53X0NqSn
UUoO6ocA6slSq4DTvCXkVYD6fQwFbO2M7DexjQIBlp97uXQuWHU1XuiPwnVmwlMw
cN0RReHF8umcMC5zpUtnVS4ZzkKCni9RBLqCWdJEr+Qe2KX4FTkaEznM9ypyD+Ss
96QRM3UaK9eBa47yUM1fUFMYxIM+W93XJgRjF8W2RaZCQqMxxSyzCAduqpmqFl2U
h3qROXL3duw/vMWvUIo4qk2tLRPMejVGZ72JLyAt5lexFiLcCVZGQta+MBVv11+E
kc++IqeHn3f+zNtd874T4f/coN34K8Ki6oZACRK1y9Ov4iH6+mqGkbhQovz59vTQ
XdMGnyhOvmAlXY4cvXXNXFUuR6y7vmHFoivDG3MZP7jFMj+5I0dzfx37cBiR0TC/
NBBIFZiXay5NoHc0rat/kj+BBUN6zYRfM+QFcS/0MALZV0xNNUnup+iEOB02hcBC
3h5sii8u59gRSTYQ8ycZUL5G3+T4HRVo4rmCEGxF7JF9gv4NNlSAyo9CSgrXjufj
JTdlG0v73/NYMl0rwXKsXrSSL56NWruaK2HMUZKi9wXMACkN20gjbnVBRO8tZxqS
zocmHbgqksVIODN7LwAbUeyaT4FzkiMxidhnkcm/fQT+I/c0YvCS0SH715zITV3W
SE0WAiUQqW/hMuNsimY7h/boWWH9DG/JtNJzMrYU97U8aI3XJeBAyeDYkYhjLRMI
2rKasLvBC6LRDFkDg2Qcbbg4qSe6oZUcq2/6MBSnldhbVpEFPK7F3fx1J86PG7r2
LK2zHtu1bHaklTEPa1dwhlVWP8EeX+nipcvvY1S1i1vIuQiyexSbbxmJmbKXmqxn
GFkskUO96x0fUwoDHFVnXRF7SNKyb5TcPcSwsBlhprTsrNhJLaDsTGdnY6ipaSlp
OU8/Bnr3IYySZSmBIA3WDo5WRb9AZrbST7ct8pC3rzhlEsrPIqKuCwKEYMEurDUE
P3CfiZOZehtuuzm1VOvzSbLUv81bXpRbTWeK8y/AUKrKc+4kuF5jF36h62RwCA4U
ybKyJJrDiFm2bw9krDTGKvppFmaMXsJEB4pH7+aocuqo31RJJJjWPLQkJIhhBt92
WFb/CdX0XTxmtV4gMtMsrWYREPVVjpnVoZaAnUmvdzA5FWuUNyF5va5qQcve2em2
ZHueXyQ5X+Nmmir2+0eo3FyRgOxN7hc+BvlDQOp39zwTUAYE9CWJnI16ULbHC1LG
6D9D0m+NNkd0snwzKfq6G03xaTO8iBhtrM5Qa4XYYMx4p5QYq6wxUhoVHqyfJxp8
pUlRUVXCRydSW84zI8nSI0VHU/7oiBS1fT97CJCDxv+PxXfB2uQWt8R2XRsYcPDB
4V7HxYe3o24W2wud/G/VtTc41K9r3d59G9eBD60Bs4oLcXJPcevbm8JHbCXdfS+U
EGe/eZowD7dA34JJoT2KyNKwJvsuAWWHYF3st2obbk1jc1NEscVXFmTPnb2/AgWh
sR0cW8vDfxj1MuRUAfOtI4FkXZy6f7ZZvFuimMkOL4zehFvQ+MkHceUeZcZXkWZ2
GzCRhBCaAxl/CnD9AQU9orE+AxdrgmfV0EgpEqn0VOzY6ePPa8WZ1Tkr+I98Uc+3
MLlbwiPCcGTw1vZKiFOnaDZVP3JMoZkkJxY4rflmVeD08jZETTrMCYh1XV4GVuZO
R2JxODW0ri7eusQ5i+Z1ElwpDTr8g6uACfewGF1ck277JmKvNHwfi+GwmxOkRt8P
S+r4iMPIDt9ViNctFw/dnkpTkhylcvxMCAV2SuYATARu93SNTLBFsXCGUxn1l05B
jcsFSsta+/pUTKm8JXYpLhQll8QNGkqVxUnTW0reRYO892aMkMn1MpbbTNPAcmto
iiGUxJUPZVgboQVTtqhyKBiE77IdZrljbwRZf2TQvkpiRpavPr6ivucP2q4oFzgG
HNOAecQ+99Y8rteg0v89OIQNYH/Mlm8e+oZq2Y1G8Ox4WlGXk+482mwLY/xV9rP1
hqpLL4F47cDcnkPafaL0ngjRJrSFLfCHmuZ7MGGYy9dwMwetqon+/Y9ZYIudmHL8
dxAZ4a1glyqw7WChcgzjTYpwpVaSJU9lmnD+lKUoEIxF2kJ3yo56/cOu1X7vcZIE
z+UUHeyAgWx2HAG1PQF927wpgl6MVHNdElAPnA8qP7wHfuDpRRlb5WqE7LkVsmr1
AcVSn0P143IEccdd2IELGlV8KXo/A9azUejw6sV9VjtbKO8hopgyBxTbXORX5no+
upfYhZrFXc3M0vYByFYw0C1d0Z/od+NhY//2ZVEvwGPU4rwybRCZVJ7PEJFPDiMt
ktoOS8fNSzBJn43fKu96PgHAu+srw61LlCUCb80tMlGtFr8k57JxeTjbDvb1OnoZ
Tbu3MdWSdM1IJcG8zSEMrEhsjZyKVDJ6ySqwps7FWJdyJMP6ve03PtCP1auoBeTC
MmzWYAgcrzRS1areodeGa7PancM+Neo2uFITOHLfl76FCg1NTz7xEPtBreJyIc6P
AQmfsFnGVoe66EpCiM6uxVICjgxIr1sSZ32XejeaWhjrRmx7H6RQrnNu5z08G7Fq
dEapfP4LgfMK4FEJOgLEpdg4SsI/MEywt1+ayUULFfoCFVxeeGCaf0huI61eP9dU
V42GRl7XXsKIVud90JYj/AcwppYtGMPmUe3FNkdFeuw7GJGIVDAFQJ3OenPdnTjn
4mY7ZhLUHfIZsbX8H4dLb+MiI+Q/OWWKTcQsVA7xXNY5nJj9CETJo2aoWotf0yO2
JASa3LuW7F3OZFlw4Ly9pEwW8o+PR+pv2Uk4kFVCZ73JX+7kuglBW3RI2ja1YCW8
CmL/5rSrQnlwm9Okbr3ZuDe2bXj9YY4UR+6dbc+pv1Ccpw1EFOX6XWNrpCKxvdfJ
tyxYP+BPI3SYc7orM3uFm6m1m08JBxgXWOJRPT98I/f2Z4dLI50sEzS+vjOOXae+
R/cWxq2bEKNd8okIwD4ebWiM4e+FBEemRuqJWyUMmAcOvlDaeyrfrAzSlz/L/8wg
yaflO7EzenmFZSXmDe0nNzM8+d0eu4FumJKsAMFBUGWgI8Tn5X4kaqDXdOYZBN2e
A9opfq1/qbR8CUGyp8UtTh8odTL7BTXzkbBaav0fP2sb666vHqhkc96pVRe8/IjD
1MaoPj420Cfl+sxqcDxO/ackP71on6L3Q78m0Hf3ed0RttThl6gjv5tcY7HEQLBV
KM7rALnJbW+wVUXTY0HPZX8Oc3KFCZrRmA1IwLtVd8dNQ17ZGQqz448s4048Vnnm
gn/cHPJb3EzEwzlYiPjFTt4RIXnEXiS0IhA3IOdhZAUH+p9NRdeOsVZI8aWcvUMQ
pAMqXYnJkRC94sNzCGNhKjDtfrmt+ZDa8vOGiyrMASbmMQxUeRMMJ+/40YLMCxAX
BEXGnjidTO1Bhgyw9hajRWq9sGktTXMzwgLjBpfvwaml8vqsWaxoner4pnEd8Xl4
y3cB4anAony3vqv469OWh4yvbbSNfD+Bvt7rpO6ppXTDEpLELjzDXCo99a9KwNS+
oFt/dHtdCirs8X6NNXxj7jeFIDvWZgt9SjI1b2fM9BZpDqmHN7v/9gbEvmvWiZzE
E6Ch+G0i5chc+SlX/JafaWaacoOecXbFddCzhB6KwGkGmQdmBx8kFpOcC4RXoFaX
oJcO2Mzw7ZM1Ed8XCdlp+lfMpL2+N0NsYoKnlOvW1oMLWcCC12o7umSjuKTGFPjI
mvLYKu49NOma2PI9+nId9U6XlaBRLAvfhz5++87gWNH7qayXIl0GGq+tTKfVLcxk
gCkJdZtToC13rVrrkbiYZIVx9BRkf1hCbZVvh1cAumy/5EpHAHkfoS0rdtKu3tEm
6gyk+CLfXac1f9uKz0gF8lzQQVfXtZYN0rmhoywnygBgqoCLa/gkyoPCfWeqJ4d5
mTkvy/oMft8hH3ZKDT+3Jo41UbKyS+Tn3m0bLlpEZdYhjdMFM3bQrlEKri205vxe
Mxw/tdSK0sKwafO3NcbnLaPeoWCjs0e8yp6dyCIBWYxgHAgks0Zp8+IazKF4ubQc
1J3kkChhZ4dNfiXyTImakE/WDyhxL6rfKFbyfERJeyhOQ7PtJq5BAiksrqf4VM9H
nhZmoLjyeUUY3uwu9aj7cwUoO6r+E6dKfyYMr0I9uWk68sf778RDTRMBkq+qjBoQ
Y7ijrh9unMu/khfUd2pFGMDDw2ReOIKXQxqMupg1HGWCYSR9HtPWeNO5dXQuwR33
GfFD5k8XuHgEPtfYioVB1LzGvpuwedoaTUWdNWe7t7lMWs/z3I93QYcnWPe83ttd
40XztNmtnxJqwweCcj7lsLwcAKP7HTDoe2/ApaBD/Z1AZSalHU2zBKMBIAi1TnQG
PYiAWWHR+0Q1Yc+R7e4RU4Hp/sCAdukvQTvWy4LsbPB+l/MQG1h4gX9OE3FcMWGq
c28taKrgPa2kr5aCZcwKgg9bFLQZUe0MrQem+tYODVbyUOf0U15GI0f/RdzuNYs3
zFd0Em3wHhcnCnD7rF2sQ0HoY6IQxeS/J6zpcYgnLv18mnMs8UuhehhbDMse+EZM
mC26XHxeSEI0ov+8wOXpPYPM8EZRCvPsYXuLbaAtCYMzBqAzN9qoboF91zdsPgjM
GF6RBs/h9mR3rCS3zP4IJ2Qn2YwzFf0gxlUjbRmerT4HekIQ84ETgl0wJwtbEH4F
Pw29AnEblxGX7QfpqgHUwtVLZWinGNj+TeFPaw0pf8o/ksGz5lyLVk2v/2/bzXh9
GMb2lG/tgzQztbSYu7ISogNsbTnCuy3RNpiHpjXxMX1UyTN6e4uCFaLPNLsaLx1s
ro1ZH/QAVNwnHrfRrgYMVEez/vfq7SgZfShYla7B+/g3v4Le9yrUPvTTQSm/peA9
JB2Icf2p1hYalqnAEtkMI+9SVWgxWVuLNZVqJBLQL/E5tpzoAiyJOsDvgaoDMKJV
OffRNyWwk05nszVMDjKkCgLXJ9i1eeAYIs9h23r9DkGuOdxwU/0VzQlMZIoItyLD
Q9rHKKvVYC6OA50yNuUDN5zTC1LmCJwHnGqk11Gqy7i88J931wqju3qnj+i6UR9j
W8AhQpqqfAseuISB09bVMfv7XWAvGRsQv8dZtQ0aiZNvm3o2AIjG8IRyl3SU37nU
e0Md/XIlji4YxnafadCYrrehVlwZrNX8xWWQwq+Gva9BWDX5wRnFQFd7HfZ0n0ZB
8f0xenwTchXvatnO8pdKAv/4glhkwQ8COP42Ld6BBpGvZ58n53xlqUE6DgeYxPfv
yYkjeVcTXROVALLMOi2wsya4MtkWXpqmDc8nFJPH7eSW1VAxAZe7i2QueM29NDyd
zrRr3TLXAZ6l2insdqV+6q5owa6aXdu+cW4gWpFBppOJUKjMSJWFG+50mjtfUkjh
Zc9VU5BHOhIQckDXwg4g15aDlDJhu2RetN1LoSjvMyDpmAdo8VooVSS+QEPdzQUh
KD/ylRYKNzag669NWTKoEfCbEhRURKKXyF061Z3ouUUTkdqT9J5jAsda4XBjKEHU
F9E3OXqavS/Wn4h35+E7irKRoAWAEbJ44QwnEvv3ocrv+L5rUCwmwXkmY8gncYAu
kHgdhdRMw2FKQ5ratAoDRnufZUdZxOue7O4TAbfiACmqnIHnJzIIQjPCTyZ/zcy8
Mo70CzKbRVUlbasC4M3ALWLfVSDKJCqVHuxtZTAuUkTiYXmJrMartlkuy0mCiD2g
4gMyymyh6cZiVl7z3wq9Zzj4GmfLIrNLBimfaDeHIcURWx7ajGZ0L+ZhBILkEWA+
xKJDgd+Dm0bipP3UDiaNsLOHOB0GNnUDUormxblaSarv2dd4FB/m2tNMgGqM3J8e
f//thK/1UPeTLKsshoS2ZIkXgn7qtwHDXISOR3H4zx2wBwvSFBYvQCqwq8GhCQ0G
3FZygMC7tWQxTdgxkaA/gHbHlfIe0C/jSRj/6xR+YQcWcASq3MzGD5af83ETjpkY
VboSrC7AcCRJ8kPSXpW1UmYid6QQM/sMdrdRC6DnlIQHOLUHgOJjFUljhomaEiup
4s1jPASLjSN6iIQcGiINDQELklMxaPo1lvc9uzmN0GIBhwG0OaylS1wrgAkyaUy3
4JaNuAY6vHDUSokIA9bFT1k+Bs1bjcIeSEqHcXLvxZffaO4ENwsf/eyKL1XY/hHw
RpkxXcSGdMy3tcd6itasoPbls3Q0CGbHCs3DwveMMfdHy5/C8J7Ql+fsFNJpZL8W
jcBnpAL06nUWNH+clviXNdtemsvOmTkyC9W3uxaaZEDTE4RVLIXqchnF7vuV3FYE
gpLrfS7vPXE87LvSYTGnFSEd7YvtPnD5SlFpZA8X4O9fUC4az9+yX6WJh9zdLt3m
gQ0qUFkl/d8Z4lI3o0flmyXsSQhsRWlGR19nuGfFdzk2rbwN8dynszHI0UUWGTdo
zT51F5qrmp4GsF0fMGwHvQOF9jLCbhezqEX25Fas4VQd9FUXd4IRF3wYLu0zfNOf
Ktxg99IXxW7vXtNLlmo1PVXIFV6H8ThBktkMKaqHkK23TPoO+VL6HAFKbkwn5aIl
k7NBJQwRwE41sGsoDtIrMQXpEBLz2G/288eOjEhixwC0GpSZ+VchXJjdb4r4GDcD
gzgthVhX2lL/ILizItgegMYCYblDQI/Vw+eIRHMaqIBXp1w8IyanVwIDhlKV0i1+
8u8BQ4wN1siCit8qwRZvC/AP/DG2EPetVDxm2R5Ir/jhIbv4OEmf1PaxosUnM9+v
zZ2lAs+egJ2024XAJ69QJ8cnbRCBZO+/XPICA0RiOY7jwFMfsHdhaZc2WUKEsBfX
riNF2SOZXo2XfclqbEckBkiB0+IlqOCITcMCaf1WGg6oB+LWv472ZD15JZS4B9wY
GbyErOpMKk4dQYM6mj8ZLg4MTeWJhlV4rXOJ1thARnKDsiFvmAwcWZWkW9UZFR1S
bgT6eBsGtsO90nZzh3fWCzmrZd8C8eW9d1bdgGXLc9hIW8dmGEbdCGQx9fzbt2Xu
TUHq/kNkyaxZ4Jc7QC58mdfMuR4GymNWmq23OHrzdJFRE0m+l8l+IND1N3E7VzMg
1X/BAwANDiKjazGtN7o5R+zEx+EBo/AWvl7WpWhDyH1tfcyc+4kSG78m8QXvCn6T
4vyqzlGmNZ1TuJwXTDkBUB/xpUSe+D1ooTzMs+XLCXVZ8004Hb+8B2tcZVHoYPCQ
HUimo+T+WZznI4tK0lLqRs8lGrHNOYspz1GmICbzOFOhay+uf2FpOIo1ITmRrFyv
q+zv9oyHsa/I7jM4dLjoZ4BWCrt+kLmdECrnp8Rtv00kjVMEBJs+aTMRnQYD+kyu
kelCNREoW4VbLnn4GBycan3mT7rsq9jGqbPDQ1p87Dhb+SS9UaQbcJr4rwGX148z
wYeeTTB6zAm/WFYICyxt+juNcksMvrYOKmG6KTLYgR70C2qAQDiSbZWZ7Cae52Zu
e49hVtDeSYNniTLS5RuMd7xnQSWfe7M9PEXZcCcIbmCMk2Jv/VWvdzWLHgeuv0RJ
xT79yZEBhi4Tq9HmE55x+GJb+59XwdtiMD+8l6iZsISdTOQH1Lv4h7oxa4ITNhN5
`protect END_PROTECTED
