`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3jCSupjDihCNOzD/f0b06F9Q7U0XLsmUKQBpLNehxkq7L1Q5ixX5LMWgreRcEpQ
JCbSAzzxQyJn6UrVvd/ysyS+5WFMZD+BTHJHxpajEU2v2BwYexTquonPigDg3dH3
DLF9JuNxZR5Y3jiF9DAiHDVaEOUkxu5TLCkKRb4LzRKM+Xy1y9ZD+CYyf78hB6EW
R9tsWpgm5A1vVH2VbtZyuk4NJIC5B0B3/RweVDse49Jnfs6q4LXEDJmkRcgGox6B
SMPFbRV4BuO8L3OyWRRVDjg2QpVtSkZD+U75xX1g/cebJ0qsRZbwZR/947vNOikb
X+2gCleZV6STSKh/Sm0XrU6prWF+71giUUfQkmUwKlXR9fVViX/lWqnGXIjJaEgI
wdjQR91VSWPBMQoYqD4217WYE4RMWsVoelf4Funce3fSWn3YE0vn5iHoe0Ew3Zva
bF9VywdEnhNWZT4gq5EwFuNgJ8vb9zmOt+CE5cxfsmZgTkrVn0DfhLzaTwix4GLZ
lMZORQftjVUB2inuMcar5y8vq5akx3zbl25ImSjUHpxx8UcCN1db7puT7XzBleSI
AvRtdzH/ACqBB52t87qWUOU9k4K/+WP5t6dKSJk+gXe4YjbPN0xsFWnfW24CRsNb
0DW7HIgp3lQNnkNLb+8G0iY5JPMzPh7WBH5TiNt+faplEJoXPmOsSSUsqbruJzsn
TaYb30SgNwdDg4YPIwzDecR1kJbCVkuI6InTl3jnvUkpGnd98fV2us0ZWV6yhb/f
5TL5sozzr80HzgRPjrJTh9EihBDSDtCMbE3jpfZnw2t9utSnMkzXJNWY4KVSf5Dy
eF8eGHj7MzKG3KD+P/ET5CFL6UGs8jaUgyn92712sApIlzQ3ywc334mTFd7lhV/P
W6hw1sFoeiN0Ri92nFRcpwU6x+HW/9qV5v+Bos1bGSPbCJZ55YQeq8Wmoj6dZ43T
e899JnyZ5eJV1vSqg4Yi9QmqHDimuavC/45Z58U1WUgCrCHZf1Rw4w4jiPeMbuot
z/rdOuFeN6oEQlBI1A5Sm9qB5eh4TGU3X0K4fwgEDDtLokfrjPcZ5t+A9UcPmjEV
LJSZLsYyegW5vhRUYFFST9WCVhfxHjiwM9wln5JT7+r8cab9UipbHyhnyjs/mae8
`protect END_PROTECTED
