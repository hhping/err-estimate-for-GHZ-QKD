`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ya9JpflPlhKwIL6Cqo1mFyvxyJqnDxkJuerPUuaGeYJPXyTUmS0BN5P6BBBPoZSf
jXf0rWtjclrvgJuFhrDg7tPn7cj9QLAAAyP1IRkdXN1eKZy1uv7YwpqKcuJrptpH
2P/QUjAX+ysB4d25+e0sEROmdkiMIGgSiJfADfTNv0l4QY35avpre/tF9h1J+niS
nxS+VmG+Hk1oqmUTwN9nxjQccJ143MxTcXTI7yaT28P5MTwNad2+BWhYq+oGspH2
1cQROh4Jcv5zSp78TI6TZqeW8XUZIhh63K5WRKavKX0HE15p6wmf8sJYn+e0POVu
5iygIxRSuPYQ5wFRnV+HoLhumCav1mG+1fsC78VvZRfY4fv2kf9XilfcejZTxkoW
FhyEg2/7aRWO5tJeidA3RbkI5PO8ZEc6QOZiyLEaVUNoKKVFxIbWzzdrKC/wU/Oj
E2A9PK65XCh0QcZGQm6+hECnu2R8GNofigr5Oms2DuOgaJhGcL8i8yfAySlponrs
AwTvs0iB1TF4+2jn2MMAp7+CMy/53lQmCDiofJUuBvg66ZpW13AMv+NZVZO7WWlF
ke43kV3ftLVfiRIojRKHb6t8yc8dfSbYeA9gZKt3SR4+ud2mULoPKghYRPbRisxF
BB/M+SC73czyNIrSEerUGHK2RpFtyvPtUrfYtROByM15GwejtC8QfrgZLkkzE1kd
hd7SnBc6nYXY61TpcOpnoJArKMfkw6WRtK0B/JDOi27bUR9AsoYQ218jOiSlMz0u
LTTOerj0v/LOPBPGYWvo90F+xNFCU6quHga1xWyr0I4QOX8pd4x4MsdD4xLDF7tO
H4sWbqI3/LYuPH21hpAFNICi+M7g+HNA6UbUN4BXJPiw2f/jyDiM+0GVB1KyxeAM
TNvJe0nZSOR7k71pIpQyNMkLVvUOkVBLgrt2O4t99dC8pPoGOfRd9f6cyqJRXE2l
mdSE1mFAuJqQYOsDQCvdd4oasReuSpCup9f/0kfzoxkfcGwjUWaGHZxV3CVuV3IE
kdFUtWWQuqtiDdVG4UTtRToAkSwkKAVRUdrvhmAgHP5/30+RajEMrXwwReUr6n2s
JAYmb1HvNy+SnOcuKlYw+eyUyudPxQucYfr5Iky/tcCi4NlQtc2GbkROlgbMttR6
qw5eYgm2qMxRBqfxnjy/B2UQcX8zrRLfM2s7wbRMCVLiA44q2c9bY3uUbMnw+R3D
2zVz8gT9Vxb5AavnIhGMN53jjH+EJ16YIpHlWV5eqQIP1fHxV2piuHaJNXd50vQt
VhI5jWMRth2gADi+FAvLiAhu4TxZUeH7lJCmJ+GmoSjB9Ny2Th+VleOvG7+hZdvo
leR578vvtoJi+3Rtc/WEQonYCqiuZSImB1sdvmh7ybkYCiGikM6DZUv6S55xVNyU
vnPgfDswqmyaxU8m6CbGHAhRQRCcj6Rp/ZT3HQ4WJwXuCewyOKXZ4FZa+zSK5Vsq
TZWvBJQ3cmPY1/o39JvosYN1Eqm2RpVnDnvub5AcZ5H+2m9eElfaR7GwsekUBDSx
SUkZwe0JwyBwOtd4pO7ldSfZFgz0Gsxv1slAPXXb+ORb5sGxwttS6dffHCwcHXOz
rWIlUBGpQdQHdLnd2DwcQersGJLWGXueuQB/dEtZ7d5mAzE8ZxmydPeCGzgTcjW3
YAz/eo7Y0n5jVDyyI8w8yyZiBr8NtnVUqYIDB2+PagGCIuPNoZ4pbqkiE+5YQRAy
DfbJjeIY+TU85tztq8V1ZUEjgMhUj00Sb+kDwKxVa1DDK0CZn3OmAoD5hoqNftOg
XaDm/pLFER1kHB2AaxT/85pGXs/7+WjAN4f0lDTeaL+KveWRAXyeg+y0oTP4HIG/
nqqNlD3eWHQ5RlI4tflOQ0388AZCs5eyZXgHq4VixKY0YvBgq6qAck5xK1iTBczb
lXBrr7Ix16UBS1K3uEqc3H/HgysGZk3e/vbn/5UMJMiNt0VtnyewOQBkPAgmF/XY
OJZnxBcjRscpprDVT0dKJ5vQO4Tq/fDqH/1FUSajafWLenhWdGkizF/v5rhzNwWK
pqJv+rFljc49s00CNd0hcuA0y8bjKRtcDrZUWDupBbdlH1pI/FmBMy6kRR1xx4Wh
jPWxLMFWCveN88x6YrN+PkYP/T6+N67rtItoAfo09LG59njRvoyU6yAu1agxruOJ
mhS9VfFgbtUyIWVVLcBxvr/twP634bW/QPehbXy1Fm3XTTwj4q8R0E/25UQbD1gd
beneH3mfoha136ZeCIJSsChLFaEXg5X4FvLtuDdnpvJ8La+1dtT1Hk4vNlLjHOtB
GpuYNDn8LqT238Wai3F6sCO51IoD2jXdl8P1+1s0JlJpgKUXki4KnSuki79joyZt
qfrrucLtOXmYXO7k1K6Py3EtI/ebMmPToMI7xxQvjkfEmSVl/NBodUgorXLyZDpE
PvV/MLOYarz2puDE9dJE7EjVdeX4OC2Vt4RYhYQYBSK7qUYe+OHBLNiWGOsCZHbe
31ZRxbywgaPh1tPI7371p+iWCDsN29ff+XANc19L2gYgUVwm7kTgBz3IOKw25uZP
H7Qk//6YcZcOWVqR1JA5bfep8YzyQS2BYcVWuqLEFftlXBrfhYLh5+cWI2/Pg/tg
cZWf74cjCAGRJ1tox1umzGNCcWtigFpq3vAs6avEmu4+IX4h3N3DKhQakgYrxP5Y
wAfbstFPnIrIKea/95aq+5CedgCe4SsIf+7x7czpRkFnd+3m7fOMLuUXYLHCU0BG
EpoJIoZf0Rj+roCQvCVeUhROzQ75GnGna4oMi8XEWqRqDK5ybc08lYYIIZXqUTcI
rafyWGXyorNFHUQbeWLgf8qkumKD27/Peo5hH2OOLu38pRYS4u0ZAGul1IgfK8hS
b6Uq1EU3ygwPA+AwvzVrgqLLnbcr3JxlqWU+4Bg3oalCpnwKDDSRdpvnEDTRI/rX
9fQDhhEjcTRKf63IdYg0qu4MOp2kgIb0C9j8p+ZFxo29i73Ct372qNZrGoHn8rMx
bhtqBYQulP8S//Q6p7Vf8/rO+3T8ZfH6O30ke0iJkTELWlOQqEhwb34JWfAUYa5a
i9mWb27vi8xUN+M19ZBaWSpUbkKlahTYyxDdxfSmev5r4f1ky84/CJQ6jjjU+Sa8
Ey4y3/IkE1EoTWYbYPYldNWWSawU18QBof9Hh+lG6mmBelwE4r5bq2BOIYlNFtnr
Cde/XAHTyRSUwzjwJShSECCmj9fLrSShpSQRCrtj8QuMC/V8Hg41MyAqPLrvH5J9
2V98fvOCyxevPZ91t0tjG8UhZseRqAXCKOfD86uXwvEmP8NX6fN34K67LA7y9h8W
yxPlOs9IYgaNCngcuwmHgoR64Fmf2z2ZIRkGlXcTSTb+rrdMGodwYgA7XTwFchOI
Z3yRSAkxhdO1QfZrNTWPJcw9XLihAkKLx4Erm7D2IyDdSOJGyIvnQgbTDfgtCFO3
Tb+lweJHrE1rsYKfuqZWSKKpSAacpy41Rs2sYeGxSMuDe8CLri4LstcnQiGOutlr
CXzB9uklMlPsh/BsRBTUvwnRqGxNI8QItQx8sIUr0d/dbYuIa1PomNhBAUN4sMoK
Ujm2rPUgvCdeDJ89WBNWF4LatfWrAKmHZes8xNpOz/KA53H030OJZ3A/zw1e0rcX
ceohZknjD0hKW5EeXh5xhEMbgQNUtcS5FP126P/B8RdWjjK2PyDYrxUFv6g3Y4m8
IHSNWWOkpW/RNW37VIYhxF2HkWEcqqwCIwzslMjiR/rw1hMw0aLB3P2Dsdd+kus5
FfE38PyCqpQO2KIDF3zm779geWNdLR5Ag0JeNAtCWS0BX9DDz3av+QYmYKLE3UNK
+e4U/A1jo79y9FMKdDm+4dYr7AMcllVjbIIdswgNpqOKVS4LD37bVeqSD5hgyQAl
tgBrdgGA+WH4NAos1g2ZdZKqtmz4Vb+KPXg/knKtPBrS0G463iNOMXjIq4oicDeq
2N4ZFO8IkLPUXvfeZkG7S+QaHec4ectTYmPgPEYxuf0363BqxVJTgmj5JnSt1NkO
/2Uii95R3GP3b/OFdPH3QEjZdcFt4/3IColl0hZnCmCo9qDJ5ZCRuG8kXb94Algv
kpiAKR8KdULUAvMubN6GrrsYrN8rgq19IhIQ+Pa3vXgjr2twmUAX7J1FDB/qbToq
9K4CpPYdRsY/+5K60uIFr+Ddpp1gJ+Rvdj/vliZ2ltQ=
`protect END_PROTECTED
