`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eoprApkFzbdACYUz3/Cm0OyxpG2HUj3RRNQPY5RkEjdiJZKA1bRSDCua4cWM1tlX
xlH50dBElhPgCNXBsZ34ZBW+1PsvvQsSBtdu5ryqcgnc/C+xIyR44yTHJ/EO/zu4
wSiIUXsJkTttS3rU+jpoRAktsWforNaZV3yR/aDE2XeO/YZr8Hu1NgRlB+TDQmQW
OOQpcCW2ciwX20dArUfLc/DHo3Sug2iBLTqYRpv4EMtzcTp0aHgafHO6cFW1bunM
Nz/f+hWgBMPoaL7jnVeuwp/Ja419DUqoBYhB959Rm6TP/xQ6wvT7U14hjXmqGrTG
GiZuwVw8liFWO6K8UphJkaiL36wpr31iFMgPvwCzj1Lr8MLIBS00KRtyYaAYxIKa
v4dF9LXa++7zx3TGwFrfWA+HCGvdS/iNlv00Op6/tyEYwLtZFLp683v5Kzz4eVge
af+jX3H2L7WqhwpwMYAq6hYeBJUMhMAgP+vhwkTZRUhHBQN+RhmlcmHuTKf6zcnY
znb8WDQ94jNT0zidsm4f3XgYP92L80Zt5oJIVOhHxmcDYz9Xpt17oyS8YtbhJZ+4
W2O+RLwLEqjc6yYJKRYXgXdOMbnKoh2p5bcfBQoMrWWzPWLJeoiwYJLqYyKJvzzG
ASNiEmbUUC1pznAEajjHp8+I4dcjMN5LMSEa0DK1/mqaIQZcmANpQpD/sXFtagXw
wCGqrh1E1eXEN1FvY+mBpsbBXtV0rcz2HAKIdEGOPB6nYge9xhN10EnRZH3oHtLc
D1koVgf5c9zgYs5mBP+kZEJ8N5/ma3CcF4KACDUyAM9I8DfllQhXCgBBi78/xL9A
3uky9Srd00upO1nW+OUon+E+umCIgGaqoAyF5zgnwLe3Jb/+msKRYVjeNIGHY6xU
yDMvvd+6C/VZ078TrdFgNAQH/QLdU+EZLcJh9xx8LgPdY300Zlxl6rRdm0h5y75H
t1sMAXTZUtpcsIJSZ/OkQsDJT4ovWh0nkNkXTq25o7tulcOmnCgZBd8i5XeqHwQF
/qlrbvZT9AWWpZMIDj2VgG3Gf5TSY0YpsSt/a2GEpE+ureU9IOajby07/Hhfx++H
+Fx/aXbs8u56ieGkcXj1J511LqrXmtav+8zEcdge+4YKpdSTHtkh1xOXfDoYmepi
k7108jGCQ4t+eoTD0JaqWGDEO/q2UnddFvGzrJM1uYEuZ9XyXx26X9c9YwaoiEc3
wmLU17Gz6TdN+023rRKVX7MqPOibvQNwZ52pdF0OhVRtRNaVZiXHOdWYO4YnM89T
4yjJGrGc+SDfJjBsaWQS5DRJWxpkPl1+hqE3O3UUJsAmdSZ44vQ2kxNyISfpkhqQ
Jbb3A8eqH653ex/BI4cNM3Z8AwfFRQX1aGGIFMa0dpFvaQDmNO9IlzDLIdvXBV+1
Js7Mn136JOhMMGLZ9RIw/8NkJTFxNBGzWqMdv81bygQjdYa/GrkB/9/ODpWtYxU8
4pcEuVCZoRy3S5krYv2BXko24uubkGZb7Y94W8h3KKvBiZF1oHBU1N+B1+kOi2hg
Rt9F8et+Hwi/BiUb1U43nkG+07ooss7ty0dpxkWtkpmq0a+dW52R/ZyaH4yPKBD0
OvnLt43VQJQFznacA/t3B+M4pCT8cPW2kHeOrvQDtjU=
`protect END_PROTECTED
