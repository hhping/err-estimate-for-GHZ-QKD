`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L5XJBNMzzhDXjDL6bAa5OUTkZhA+mZ1x7RQwvmei7oc8E0/HBYohb4tYmOr6RHfh
XmAWL/do0FT8As9JZ0EUwY64LtasYTxcqxYeY3M9UOHV+TjM/e493ml2fBufJhNa
Jc609thWEbM8BtkhHpCGGDW4eOzZIY4nCvtONUZKzegXX6o40Tm/bKcOOcz+fsXg
py+284LiN/foK3bybiA1ectmDLGsiZn+s7SwQiWM8vKqovbGADdi15J09TaNfR9x
nTdchEC3DY3ZlBM11ieFX7f0DcGT62T/ZfJj/sx02yo3dZmnrcOqAXbLYkrM7aJF
EvNGEI5K3+HM4Lg/AO/Whd0P071a75crNjA7omJ7yrv24K550UHmUVCYZ8mxVmJa
kkhoEE2kh0hZqXFgmWlcJdZCG/PcOdEJNxAtKvNKvzZVuXCHin2WuLVw/OwCtlw7
u50C+CZndvNhoUlFsyy/8x9wczRqUMxLOqOalbKLm8loh37vAiTrVoNQURUdi4Jo
8jdNxXTYG+MBBP6v7ThtyvIzk8v1om2LFJbI2bHPcevDZV/XCvPVQssGqzBjjsIw
m6WNRjxZo4VUBwoff5OLeGpSZZcYII4csQnsH+rPr1ES87sFFlUw8+JjqIrw4Q7E
ZZwTgPaCe0OBCsPYHP6q++hBbwJ/5QsiJIt3M3L/jdtvORue7TlsbsFRR2ZEtW3M
gA3sYeeXyE93sLyKjtgbtA==
`protect END_PROTECTED
