`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eRIrTbvgju2dzpcMZbrDXHopdr0qz6/jHi14KjOMqipHZ2sQmexnfeaJWw70hdHT
1/XFv1Y1e/qL1MvpchYrDVrmoz32NUlNcA1rt98XMYTuoG2u0XxjbL04rGIsqpe4
Ly+E2KCOfpVCopacRv91cgWjrSSw/bjs+/tlbft0VdNHAJ6qt5iCeb+Mll8CH61o
aOQ5aezbEhbqOVY7Wg6t0QW0qGz6gle+aSnQA8GA0cb6ohPcc1ZRYn2AlbyhfvBw
jffC6eKeje9XkPzRgUCCrvTT+cxwmhGwdiK9xLj5j6po4al2H9T1wSKvRmdW9egT
it5phm/XtG4ZxUxRzrkHFJvcNjMMy7oiXiMvPGMOeWTfB9aSyot3Ho5kHQGmHoHx
rF80DTgb6m++DJwELolgWkJ1itAknSYVY8yjv0axSZvfYd8Y6BTaPBAcucvFGlL2
ERMkS3jW442bTvKCx5MZqkgToQHEoTJ/COUGhkGfxKplCYV4xSO2bCOi2aScck6I
KStA/NjXID+cJmHqJHa7MawgLi0DiY/htedRBiwijbj0rsnW4ou2VAPQfCvkRnQd
t5ktBwNAmfrQsv7/EC7x6agZZKdOEYKtAVbFmfj0fLsnbSmSd1UVNUQaJWjvQTts
fb65VVOUF2hlE64rPL0jEzIJjDBNd/m1Omun3DDiVN71mAmE05vXR9JuQ2xdLRvS
`protect END_PROTECTED
