`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3t5ZzsJ/24kxeUyHJGFfSIDYyOjIxkxjaeOpu2u5w6aDhjPl286wFdJD7K6Y8frA
LZK/BB/Fkq33bDJUax4U2aZDw1eqsYjH/QutOL4JB7FGEERQRY6dQR84H9elL8aZ
VinRZPWpmAtlNS8Re1kIGEhhUbGRGCFGs0oz70cqn0r9rNX/BGCkxTIDx8pRADiB
fyVaS5Zvf0p6gilWN8k7kXu6cCNhy+tBKz7/c/wO1/uNlRhxMtU4FFM/DjhgJwe/
UcHAcLlSS19Czev18xH+iaJP2wWJujPRzfQ0JHu2mgyrh63U719WQK102lX7/Xm8
LbSZVDKyHud3JoOmfphb88c2Lza8IU96nHNT7ULe45MwVevxUtz2a/UaH9kiFnkb
pobPXMISa58aYQuWViTARN9JMYzoEAJYniwuiExCcy86tJo1/SEviWE2jkp4e/0x
pAEDJi95kZqZ+BBUJaZFBGGuGZGviu6O6hzo8a1nCT5tuAtGLUY5gKNiO3bmZvOE
zmLOWCYAHX0FOiEq6eOZPxPIUEnWM12T4C1yQYPF4cqoBry9IvKfs515YZtG4qUS
HbBSjllhmPTO3jzR3inlAT0KhEE1GT+aQaj3VJcoUzWXJlapuUoGTI3SS79Urdct
0n7dvS2mPhxY56LRlgdRRMTPcv1fc4tBTXgeDaxhV6b+dpJcTArZqRldLUH/Qmsf
`protect END_PROTECTED
