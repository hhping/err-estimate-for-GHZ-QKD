`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bFYYkvYUWhCEl/Ce5Z6BkIDz6wdHBUhFpI3txu+DFL247U8DBRiaxJrFaY6SXwje
Bqg8AOQnIodXjBqlJ41Yc0+6vcB2dzGgSrfBhSWKYCF0XyDGM/QkagI+WPV3VxHL
DRQDcg9OOXzCiQQY6T3QGVrIGTNi9+L4bqQU64tFpOUh0kYXIYdk+XqlcXbipVEX
3K1aFP55WXE5TObiq1Bs0bAnk662pht9C1+EdCSnQB5SZNAW6H/N0A/SkwpbJOMR
PUhpva9jyb9F5GnWkS5um2DQn6uy+w0nm3nBKDUee3qdpa9OVT6B8e0prgKRo4Wz
5OBod89qgNRo2DCeTJ+aDeuSKT4E8NaufH1bI25fnUc+0feFgExnUZNj00dx3Cbo
0vlBkxN4AdcyoGFJaMlY5X3ahwRJ7gB0LNo7m7gui33Blboq1FXOejQkXMX4Ek/j
pF80MBs6XsohDxxq0znB3EcKV4E+bNw+vvPvqlgTz+rdD4+iSL5Upn8awK2Om8Kj
skXULlz6RYlcV5yQYfjzYL8QXz5Dy/qW7my42Qu747z0VeuAyUGdRsbdzG3juVYp
/wx4lSbAQq0sG2n/+IP7MXAl6wjtxIh5kHSfx5Hywi7GjZ1Jlyaf0MrC1Sh/kZUk
hH0fzP8w4TFjYZ48vltaCMJMU8bZvRRBXyZ0rfA6ciWmJ+SXHej2tjBR6moWoJ2g
iOqJlwp53O1RyjTC0k8MEo6kUblz1FUKd6UkulHOkia8vyLsyKDzzsHIIhb6R3We
i8bqmnK4x/WUiSSecxV/Cg6k6ifq/mWLpeGqmt+laYIph233MqSidWOrAxrkeZNT
C1fv5YeDkhvr9/v1ZDrFKaXYawgLKX2VRpA+az1vHRD+UTin8QtlJ6KqUdL60Th5
ZplX0wleGkhsSrfNYmiAGxTx33Dm/IqvuhAL2nwkYb8D81V+Kle5TssK7IXiMwao
elly5Tw6yhgSbXvQk1Eud2IIoeVTJRLVsuUrjNHqXPgXYlY2cOO4Sacm8Ozniv1V
1HMQeqSBO2zUiaSEvvBpFnKVgC3fPyb1KVKfOj8FFAbTcGsklUe9pFlo7ZYRcvwR
UYZ+LU367Kad1eHVikJRHS6ZI04QlYbkEB5y+9Ql6uL11AKYAY18QhusvctEJ0Hi
aWvpvBXmZg/NQ6Rdy3KOIME8Q7GFOKYsLYtuy9LC9M0sW1Lenndn2qcvCzzTH0bm
3avLoMv1C7koIJfcMms2JCK2mczrrsmKdyO0JVr+MG8W93RFT6RY5RluK62QMQ3P
JRczPZZVlPFUdzWmZux+Yk9w+f9gL32+OcdiU6nw0XheTkqcAL7KPZYBk45xTc62
kEYeoOI3Kz92NoG2tsXmD+SIO4kCEJx5xTkHY7d87FT7K+crFfXs3gx3hJ0CbXIv
1eh7igDSP27Mv/ahBTjOu2zzyjyg+nLEWHFYCxtwuO0cK3M9jSo2rQRm+JeVMoyC
TwASZG29BYebVA+iSINfMZJH5dWzrvM+dBeVPDj/lRnidrHv/Ueq2PV4oyeLH+DQ
6DPHMDNDuLtGNHdWSuG7aZzeT2AkO/3PqCWyhu74ZuuXrAGkgx9qShL2JPIHR7PQ
E7HQV+J9JUMw5djDYnPNyyaX9OwNHfo8R9H9x5zbZNe+bcRheYwDj7zMqmcZ56hy
WeoOiQpHjFMdePCWlJmadPIFXb3osPUnS2oP4RrvlmsWVBtxpFoQhJugpK0lr6es
qfNNoG1XgrCg4m8Ppphva6hW/C5uJJFkPCshicSHEvD6umV2rAtONnjMI9NKHfie
07Q7Ew4S7d3+aBdaVkQKOVz0KzM/DoiWyTxRCQRVKdJj5CdXkLx+DeGGD6PAIGBr
GTeSX6DXl3uUjZf7MUOe4epAKKkMA5I6YQnJNVVSROF97qiTIpWLqoMSHVRNWMlg
2sefMaEDtwxye8/gZp98qLf79ib8S9sl6UBWu8hkTeIDmpM+5/NmqcHCFHjOF8uY
Ax0eOJt7jrKkpdIZp63RN/klct/rlJkZyOSvbyJiiVTnjynZuctgbtwMjgbZpyki
Q4pMU8G5OLMIF3W/SXWG6qgsHbCwGHv9Vh3bGOKF1iI9g8sX9CorRw3TwYWAhDh9
GLlidt4UXARmJCjqGL49gKQdq88sH15oLEzFPYzFlRtawu5BGncfOB3ETH+qi9sX
icekFFiebPPmxLkIkd19+HEk17cuXcXbT6F5DTxMCVQTWAQC7To9pCIoOaWWHMOJ
ElM/W3bEW0tD1EXh10XAxikbAO1AR/yKcqAkSUn9MRvuYlqwrAJUeF0ducVPuLMo
`protect END_PROTECTED
