`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uSSfF9/b8yY05WUEWmJoHh11jsoEPOygxvOqfloEtC2Lo9P+BKcAUSatd4o8C0b
+ZFtfTEXyCz830kN70L2Iw5BPQQ47AbwyZuAfGj4pcgn6QzxIAVvvKiq0UrNDaFe
gDsb2XXid0CcXslmzgisaXt30YOgmtN/18nuW670iEBj/DQX2D9q17i0EasePU0l
zD8iu3fIp1D7gVHraq/0cl2Kh5lqH6dLhccj3GiWATScA9HfmkW1xLnjPhXPA7Ms
mG0R6ytSkTaM8N6tdo4N8eHbzxg69WysfXctRqdxtPnAJoezc1SFc6fTJzCdIDbI
ZyUoyPhY9XdpTrSt2qOo9wYn/kYpcd+zzfggsWRLYWtzJkw1gK5HhirHhKxh1wea
HmgbWu1UmCwDt8euqBl+E3FD77VFI7MhaW0m2u+W1MTV+vQlkNc75sI1RiUhabbR
d20+yfMJWSzaN6DHRM7e9Bm+1WxpvqGXgIrHycUQGEAaL/WpH2P+cpEHllL95Frw
8rsRgPVhQovURrmyxYBcVNTiGoQ4xB36gCh755Hj/+V968O/no3iZw737DNuIbcm
xA5GRRRKEmao+FGlQ0PEUusDzDzMzRXwK4/PkpWBr2ottbu7L6Kto+RmmCqDJGiu
qDc8g9ambGwp7ar5S+dgV0Kqa78Oqo/I7bnJuUA6dTY=
`protect END_PROTECTED
