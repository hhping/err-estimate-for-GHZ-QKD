`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KnwNlbi4uM/n3HIeBAL+pyO+nKwhkDSECtGVGo3X1+glvH0zly0CjUDKgoDlq1mj
8ouVQiVr46GJ3ntvXODzgsgg8+pcwG1ckJxO+q1rC1gTFLqVz1ILEzAQ3vOyi2f3
4JDEGFV0TEHx26XvgI8kyLxA2Lbs1jrW/O+98mY/P+bDIX7cGdL/XWyt4tSScoH3
qieGS8IjLxnXk1oSeoRaVeuqPoqC8DmakkVr7L5S1RKGJ2VwVNHoI/ah72D61GoV
GbJFcvOOjXtgaG+jgn/LIQkCxge84aTYgsfSdUGkpN2NHeBpPprLnVc5XwBZW5D5
CRGHnUAazZF24bydezBPbsLBLEKedgRe/nlvBpv6K1GbNjZLu/mToQKSIASye6DQ
SdwHJbBBJAykXI2Q967Iwfsl3Ddre1uB3aQbwPdDoPiZ8dUryxU1rNm5Sbj22Fr1
R62VPaeZNppPn4RQij9EnYDZdhoWn6mF0E/pJ+rUmsTWQBlGdBUpmbMWYn6qvxjP
gR7vo14FT+ezSfUOr/bCQGtBcZgXJx/2Da0j9USPhGdQDS7v76ZXmFR9ef9ODCyN
RdZdl5cexGaaiFQaHidyzw==
`protect END_PROTECTED
