`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ur6N7g/eDqDGyL83L7hnhP/ISespMPkzRFvzKCDcUEDFp0KA4ogUKQA0Yo7IMiOF
IR8q17w6lDcl5btbaZpVX98c0iyxsPsGhmcGKijZpiGKf6FkTB4mS+BMHw5rH3o5
pz7N5iku4aQyP5fK77ithD8R9k7absSsk6ZVLlvK3TgQtk8EepE5lR5wUF7Xn8UU
NZiHxy1UB4JnlXLHVdmlydiHU9ZTF0L5gK/k2SrKz1e7hqt/tbTd0S4MMbOhufXw
i4Lvs78ptjf/zmB1uIkexyyUsyiRdht9Gb1L3A5sETUlBTAipv/G4gEqWsjpx7MO
48NGsYoqFnbPFt4bBnX5zbOeVjLmcQIkAu4yVcgIsRA=
`protect END_PROTECTED
