`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QNuEQRf8FaBMRqegjAG2gdQjW6sAfolqDQE6f541tHcdyljuSXQ+ycBl/uJ6rM3o
oJ5zo+MoT8UqXvpOJa8l8NOG7M86cGDnrDNgmQginT2OjRJyTSdDdVr4cTwai9IP
3PDNioISHd+PkWwXviVofRIIX5Fq57upBnlmKX7Icvr4gBuOzZgpqZCLcMDrXQ7F
NwdQfVB6mvxZPXpWesJ0UuniOr9o7ZhPuquFBXU0wIhsq7Cwdp5EGCH4Yczj6Hb7
mzOObgh7jEEldf2KbsPOnoqdtUYiMQLNXLaKJiraBNRVvnrTqNaByixwCb85fPNe
Jm8vi3Lj4piHJbtQH9kWfCbpjLqEbWz5hsn8gNUwE8JLPjZHcGu8T+RODco5uPaF
0UxQaZL8oDRyBrX7jubZKhoW6azOywGYPtaenO9+adAowz0PXfb3DeYzJfhtAI6X
wm8GiK3lOVvGPNfAA1/JMR3H084Onqw/O5D79WvZfWV0i+/baOFOUE+wUrsJCjvw
75uqWOM2uxaojg6z/PFsrrKhQVjhfj/p4T1lWwm9eP1NPSmun8GyxgmTbYiRPi+Q
9Emi+LrjN2jAGtYPYjYsBZ6hp965nP35ZPl9gubbeVP/vi1VIdfCVtATQleshveb
NlOiy0mtiGPGOJ2ewSSBa2J8jR/Qt0p93/rio8Du/AOQfflha6iwzUMFyGuJeZFp
r2ZYFu7H0SiNLJv7P7MF1OMlJagXUL77oMytcmJDW9TRpH8PUOjMMuuRKY8vpx85
XnFKerRvz+Pu7sRUeLpt/9Egc3DBQUFAE5qOuUxfkmbK2a2ykjNDV8EYq+aOKbQr
kLuzHt62IIxXPGVhFWmyeNudD0LvfMD+OhlveKbFX7YZYa0Y4DPXVde8cWUgXR0T
hKP+742zzmIcOwZu5Y7QyhXrxQd33HhrHfQhl42MlloqpyLxfrTbFoydsablFGOA
+cIre/6vMdOinWlT9VPtw3SCPLMjCD3GN6iVgLrExnpSsTq2bE+uxG4aFLN5ytdg
+uTrlOBzpUXwp6XpbagboUlBqRTGCl6ldD5Z+8tgTrloU4Xpb8Adx0wc5CWV6RNO
OaE7CgmxQex6tJTVDr98UsmZW8LV6LXv5qgC879SkJbc0KCGFaS6TjZFasvgzMt3
0mfI947dD3zQrvyFtf3hMxsx3utG+5euYT+76GlU+y7LOjtzVoW2r8kjWY2tIIzd
iOqj3pi+OPaSMg+mj9XCp74ImUO4FZHsoA6FreWvV2WrWcGejr0p30jIWhR8IAVs
Vf9LqM0YpekcGvA3LglNCUrwfVO0HFVgOcqk4fewVbXXkt5r9qr0kiLAhrIbGOVA
Yf1dNcfFjYXPL2dUUeunQ3N8ABvUyEeUUQmhX3fLpzR9hk91hL0KbPb21gfhpFJa
uP5VuJchkJ3ihzr2eNwudpeXS6PIehMlJJdboAnjqyRp39uTfV1uPjFuWcAQr8IO
TK8n87HwLK+7WTy9GyQ1T1IibIvUqX0bmj6/fWyDWc4=
`protect END_PROTECTED
