`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWF8Ksl8ujKYD9BsfkgKp/WY40/CUoOr5HYtY48WubgzMjwk6qgSk3Wm6ZCd+Sb/
XAmkkzNavV+uWShaj+3guaK1eomO8+sGHAektI7jrPCj91hNTqrj26HIU+hSPdgE
T30UVvnp92IZV6oUSXKI1is+pTdXfLVCO1ibPDl+oWRGWSAJxJ6hGLbiReZt++Ie
uq5uyuMIGjPkGWLtQoyvjKLvqMc0YurVCNwhbhqkm1xYQZiKOp9AWwxEOcNqA1fs
ZgCF1UEYYoCAcPGjz7Xokgl/Krvu7KpWTVW/XPS3Xe36VfvTcC/AC3OJjqkXOr7Q
0bcdhU+Ezck1xJ8WJkj/p5+aw64rJx5Qpnm9Ytn06/odZtRDmB4eUqZvkVRhQXW+
j4Mga6aucGwGNuZPNwct2nVuu/7+8ZecvjwfK32h68L2DGERQBeTqGg40ARhquSC
gk3Oq8CXSupkEx8x89XZqTxPsi0jeZQTdiYNHQkqmk+ffLFdiJGSxta95c1CMZx8
Cpfko+zHWU7OLalPbxBHTD1bQD54lcWS1MnsB4vyvtVX2D4J0Hbe2vqG35KPvUWO
jCNKijaPt+4wrv8ILND5PPMRkIv+aWKas8tU5y96zDbogXDhNgC6/BfX7s1f77yH
bTlQQtZ2/YoR8i0V9Ya1/TKfNpNJ9o50pAifNJtyVDJYlPaDYWvzCSwr4GiV6zZg
JZc/L6Qi8AHTEr3GU8H0giZt9XBHIbf0z2YI8BisYhcnmo3W/U/YXGvwj0Pvl7SN
0P4lioraOIpJ6XUqSgJtwPdYjGDTJrIybRCrA7G14ul6RgYS3NSRP7rIeJPE6ezA
pzV/1BFnLMoVoO753ab9Zr7q/h5Co6abuDFJenZswzdb8EA56BDpcZBwnvZ42pgL
`protect END_PROTECTED
