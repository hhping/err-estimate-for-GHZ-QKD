`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWfKiVBcbwcYi74dAfb+kXCZ7kjmh6lKQomi83lHgICFwmkGdsety2sqv3CeK1cv
GosQqyB74oVgJ6W6ZvFLm5vn4LfQJY/F4SLdEem5//s77ALCnRdrRNS1vtltn/9M
Er/rlYpjpGBwGFV7/SwuLacABWRPbWUWrPIL84L37WmNjFOAj6R+by9sDqDBBtUW
T00eFZDtq+ZCd93GpCmoEI24bfRcgPlRTdAPnepdWUXAeSJ+1ctRXOAmhxI1H9q3
4RkiAxss14DDiNKV8w3ZiLZsgxCKMzZYEt415Lg+N7alUiTJOosmBCCSptlHCZsJ
nPvPgNumcA9ADvRku7SHW4ckqWqevTPZ1SnDEBXU52xba5rH6hPaTNkK9umVNaDc
03G7GpqEDwsCrRMgfq9gq7LUEvma8SjPgeQ5sG+xZKB0P43vgMyHzpaDH8AUmStO
qUM97jshVb7OJTvpExJ2oihhzR6/Ve/rtb/7tlmaWet+HTRBvVvRBcf7gu5KnhFX
ar6j3nXUdHstSoLUBt7DqLR1y2hPrPGARFysTI8ZHYJPHK9La408FbRpziIgnz7V
LjpsoxHGyhB3CA/fLFs4hP0o6RE52F/aTkmRmeTsuoi9F/Clolt+Gao2H9fQNFTx
o0SExvgDweL/vsAadr9C22bdM2PyUk1Cgum+jB5/2URxLmqWi6P653tQH7ztJEKl
xV00RehE4dthR2HDSlLW0FgaiuZfZxly5qJYTCaM7HebLe/3MRqW7H/aDB9bHyP1
qBNcT/8Ru7A8Ki2VJiaW5LGihS2k0Ho1SygQJ27IBr6MZ5cDvkRBeCvLqYP0mGhX
FjYSSUQIjZG0gKI8H5bEycxTBhQlzzqxDchwTI3iR0PkV+GS9fzAi4mv3kKK8l9z
H8vgyIB5A3u1Y3kfZNf+CFcHG0DuCgaljB3Dy/Ze5KMASn8GrCE8cl/7SqLx+ckr
jCYdq0QD6npDfDXywONJ5EvFrQIWGE6+KW8XMHH6++a+p17RC2c1BT0CYggxdlsN
cX2o4gpL+4WdkEhLrrK5IZlNHVZfZ51tCu3Gg1wv3pkJFxa7EKZxjgkuU45eq1Ot
SFSfs/YtBPxSojRkI84zJLPVGnn6jMFguiUN4ZHGo2eEc++HJ4aBy1XHwMqcnHUP
RkcE51EfQgUrVWbAkpZm2BIfX7U4cVn/fPZedM6hcfJOGTgskUaL1bmpug9HVDJU
62xt2G1xY/EbpRXVJXqW69RkwfikbobUokE21byy4uCw5lQkUuC4H5UAks/vA0af
AxfIFF2XG8T0/5s2MECoY0mfoBrEqiqvnSeb7hglKdmOEaWd27MbwSpWt2NKasHL
5hIGiwtnv87xhk74Q3kgwn050+24QDKw6NbT8ogC1ZYUpf+LrcdUDMjLU0PQDAdj
OWOGBopTkQAymygBoNP3LjcjMEEAez6/OZ0AHsgkGGaPTHB3uj0rkUj8QNZd/SGX
Zb8sUZg6quBw2+YIzsgmI7tEFrX5VEBcoOsKvfK5pnIH3gqY25caHVCrQu2O65Zc
c80EgKC8p3Srhust+TU/hDzqKKtXi9or4wEjJM6e7zbTacmgM0d8CzHXLtcq0kbx
`protect END_PROTECTED
