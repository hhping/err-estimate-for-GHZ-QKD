`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPqUIXt9787Pj1vrMMcAvfBH80rKAa+QvhjA+YvkClJG8p4zW8jnTgxa9LFCoI8D
wUaqqddSLx6N5CyTurHwWQ+5NZJTNrPjp5X96NBE5znGe1cj7Jl9z5L+dDJBBfXi
sev38sLxmQKKsocmruI8wmdmMmbZuT8L3D2UIPhOb+hAnlJpj1pLurOiVq1p7TZ3
rxviiZOJdUp9j326e9sSlHkteW9DniGvJ1Cr5m4VY3EoI/X8RuXmB37ZqTzvDVi2
tXaTRObzCUNhuQdvgPb0LEXG1gyKJWv+SU7DiQwdyGrFLZfYdlTFN+1TCdnHvQKa
u1oa0a4DASZIWPfo5PH5pxrnM1s5RhTVIO3dv3KLlTJ+i9BA5U6u7tE5mnG1tLkb
fjY5h6sLPG4oPNxGlLwVrmDP/RmKvHOSaW5OaoyQQtUSgU5XafTj+WALZlh27W91
J7DSaTnRQA40i+hWE1hJcpmuCupd82NtnAgdfAPlw0yMimyK/BsnQp/C62C173Ax
vFEcXJSiCCuGCaHxZxjZqtYbI+s8VJRmoUA1RJH/hc3a6qiHMk8cy1MdkpCiBFYP
wKvZoNR0c64wQAz5wDHPT9M6cKLxLZxkXhgb9wyh53yX/Jv4weM0IIOpb0RRuxt1
Qa+a+mBZsTsel812A1v+vRqy0+MfuSVWpl0hbiS1lFHzVY3Gw65rW9SxTDnhDGEv
uUoql8iQwpmgbPghS+mDDHp8Vr390udQuidb83mi32uF9JmsrnpzcsiodrpA4Bf1
96P7Ez+b72B6FYlrU+A5fOQ9R/hw4wM+nsAToQRO6BeG4mfeG44kIoiazI5lEhC+
vLuRTX02231Vv3Gr2u0I1UOfoVuQ0/cv3Z3FAMNvzHJe7ZKg76os8QYnqmU9EmIi
QMxhbpQjWN0qANtk9SKYHZLRtJN89O0+hGctSkhDs3KmFQ4qPhrf9Om6zqPnQ1Td
HS6b8QFDk9e1Ax0W9s6zeBtv1VHFRk6fFvKEIjhQKMH532+sxFADuyCiXH+kTnfR
dp1QDFuWmSvGXIkiAAZqj0POXiYazWE7lKYdhwsrSV4AtNELIhES5sSKkkFbpabF
ufVAYwNQD2qNRcUZp0sJpzNBdBe8DKhs8xoR4KKarxQjHIofgGFJEcp67FFNLLNO
Vuf4/WnUB//sMKtMkpO40IeWqbBHBcP8nlN5NyijvZaG9CTD1En6NNxlis5U5jro
9AjCJfy4MqvylNU8OYWmFmvzMh0kEBwAZYnlEyrZi14zCombMgVcjtamNhPOVVyI
vs/GCE+LsvFJdu5SyVgNL+XefAXx8U15/gbnYpu65fHNZ62nnBGlCIWLDPblXcn1
mmwrGk2irP3Sl92vF2iyECBIUxl8x3kaVGbkoKnsUFcvBjJPQ2EwcSVfNYdsjKxb
9/OhHtMmQ+sIk3d4iibLYv0E3VMwOLjcCpLeN3bLTGCCta/oGevhtGG8qCJmYRwn
pJ2NuJGKXZYiWl2eUQAW1PR1gDMMiO4k5jpAsmmAD+14Jwd9gv7clYxHV3gWPYfo
HxlvABzCMHujNesXVyZpJarP8xiIwlvcz6tTJthkfAg3fJHYcZervFNUgF1sxfFO
FiTqdmJTD0IY6mX2WV57412/b+5KekX0e7MZ37mPSq85JXWp6dmxaL9q2MQn3Jd6
Wpvlpm8MXF9BOgcVtvjmQ+XMQRvJR9XVi87iWfjiU/wWQVbYlmpH8hzwc2MIUP+F
0wH3Pgz1BRzIyapJo5lqSeJvsno1NxfPoGr0ux+bc/B/lELoVpWPcGELQ489O8WB
9fnpInv+M6xAnPo0MWswpUr/yvidrfDSFJpXQaB06WXkrq6ljSmTpRLhWAcUwXEz
p9sF/HlbaURaZD+GB85FeFECaTon0XDTk38P74MJ3ZOCdSv1sASbEYes7JqiJzTh
XqAgAr5HqJoOWrw3Myb7XkCyZDj088/87MRq5ph1bvLI/7YFy4XD2yHQwJe3amBb
5B6B+7V6kut1qrBmTDl2KuwdQ9sljIjKSLWksR3aPm5MzbF5FKgFs8Z17/YtQwi8
g2+3KpUL0S+FONEPo46TbX/UWZfiOVEBvoIYBnryixHRhx0+1GvTywBrz+f2k33i
IFBbETaj0ldLohCSg1AvGGtVE1wAYT1148V/jcYkCRNZk8tKQr2iioWy1SpkBlqp
hrtFtCPUC/QtZTKpsxCkmCps/aGWNKoMOcD1T0wtpn1YJ8S15QKWXf52vSunqoJ8
YbIiWqV6BD2p+eYGBglnApB48+XOEzWJK+mhdmC/fXSWAih+aOBHMzCSUZlQdzen
Z9g43cqzJ/bGWcF/Bo5QExKpPbTJ0iHJla9/935uk7eQMlSXFKhN/ACscqU/D49L
WwyLRSqUA4ZXsBu2Gv7WrR4Mm9z43sX/Z5fX5eW1QHGRGUR9dmNCjMVJWv3Ur7/u
W8lsaqcBqCH7XqoltjVLCAvSWtyXc2+1DyIktbG5vGgbRzlOuGJA9YeTOVytqVtZ
xHEbVm/1vd4+Y/+cE3OD/ousOTwbi2SFjGXzrEyUHqdHXhjINdLpnXPVHODNetAT
MLV7vtuBQozuWfycqNPXl4V4KDtEzzGwx2+OeWl+fnzFfeQMAxv2u10IE6uE6sWu
Ox6SW4VfEANhSDvmCJ9kkaCn7dJlz2zq7Ghnsd1r8LpTnxesXfIlPLT/Zof35Ti5
SSTl+thZHMMx7FKjAFUfkfA8rfr5LNPIPSg8nA0+TTwuOZw4RBxf7Ojbt32ygGKo
NITmDt7rch9wFvpLckq+hPF/43KZhA9VJgwsFcVrjexeVTS44B0TspnVrVYTly39
PZJuH8NUQ8JMNSvWueMl3ECara1qHqmZhZixDohxWvzYm+knAQ/zjd0teSeth3FV
ZGRrh7l1BDoLIr1izeLEIajv/e62I1AbzlcjkmgZWYztPJU9PeVYjMi/o3Ouj6UP
U/v0M1IT2mRWojbPjdGrsbKKIlij2sO0xh8yErYG66gQ2Dlia4YCQpHBblu0ATjz
ecHFEUUPMxTf8k/tZo0TF2GdU8KyPGlugs2kaxQ8DKn6KNqkCgKAlNTpdPAlzrPF
0xrXyDtc9Z3GrVBp8eoWxWNgCoNHPIPMG1olqhC9iJG5DU6HvlBGtOiOT4OIFJwM
RjhDVeu5KNYqp/jPtoLqq/pBnQj/Z6bW5uFEzF2zQt81PmWjKaYO1QL2vNORBeaW
uR8gmafxTBpMzZ5ZLVrsy/RP9dfbEDueHxOzihnaoy2D8IeR+jF8vKnn4PZBI9Sb
lvsKs/JnA/y/PtZrGmwnshyyl3IuZpoDt+/0M8PloqzTnbSuSPoJqsk12vBRCv4P
onb7gaMUZ93k2t6HK/KD/DpH/Q+/UIdy+SQN8MMWd8xG5frowwQvTCvrZbSz/xFx
bX68dY5l5+S9uMl7loRgUPa1vd7QWfjjImwL8EKW90dAoXNC7dQ0Jp8mNpsN2vFg
fKc0Z+2/EqZKdcYiMQlXEs5dwXa7Zi6mdqWWvdMBgqh9eGjRjC9iquRkdGCk320y
tolXpm/pGa06i/e/Z8rQFx6nDymSJ/5/1buLfJu97Lk1mPydn1cOeLsr2/XgtQsy
sF+FW5iwvtw5kmevkac3aKXeAk1yCgKN/yDevqO9G6KjFVBWzkPIggw48KBaxwqR
aPdpJLM349uxjS1e5Vd8WlZPKyXaFIsCKaxcrdlr8QIyUd8o69yKQ/fzO5UTcG99
0zvSOaRh8J8WNJK1UWAGySD2obz1A/8H2nSSSP6NRydurN8LOewzwX4tQAq++j0B
GyfpQmalpocrhdRT8fchvpbMBT0gs9vqkI9Ehyzr2+iK8MWyhFQgxBL64x8biw0K
nYK8dby4K71+1zRLzAbseciUcG1O7WAKpefiL3fAI+X8R+ZP03dWUv35nBFSMizp
ovIU4s35uDGogfvdTzNhzT5iHgZoEd3cUQD3gNSiIBfhK9fVc2pCPyHbrLZRm/bZ
rlK1BpfhpcOS/Go0FEu97g/jAKWeqM45l6RSUDlX7ZhFKw4Dli61lH9N9uFXNnHP
IdAbzArd7iuyyd3zBFCsZP7xvTO5YrQJs2dS/NEJQryJ2RyKrwwJbsxGPFhV3o2m
qU9uQqRdPUgZ21BzTd/Zi7IWOq10+CZ5qSfG3vCn7ynSQFXA+ouK169RCInBvwBf
ChWj/Qpfn/0EGOHDgLAuCzR1s0h0elZ9m6ZzctEaV60EENzgRJlz0VyNEKXgyGJ8
e2dOVQicMNJPJtDaFrsPlMI6ylGjJmSuxIlQmu4Vp/kG1iclZq7cdch7TRW2gBlK
eUQbGWze4ZZerMB3RnAXALamw9owfneZbWxR4pTzPurJLNm8kLhnSV2lzi7Dt8DU
hx8lQSy42B4hd8ej5NJ3HrV4zPWKPbnCbj7zKUiAVqtxgc1oWoanZe7FYVUiC7os
7PYWCIGzt4OnIMM4sByS+bkrn7ijQE6A0LLFGSHll66omYdEq8yIcfzTN7iWZJTw
a5/IFuDMicj+9c1h0PG539SUPy1yJpm5RcUsirz8JC3ftcTjcepRVy2bazmjm6YO
pHRq4jGiROcmF6jHYwES4gpb7rX57yVarOx2/AVe1TzedqJC5TIDbFhYMXPrtj4P
lY4jG0OIX3axo8ZU7mvazl1jqCtjzjVa9gSxFrz2Z9l4WG0oiukRAcq96FmGIZdS
lLGyl7YpqddOdWo5Zd8KPw==
`protect END_PROTECTED
