`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvWZjag5Qg4XSP5H7rR0ycFzyQ5ADmQYxIgSbH8nRUNHKum7eyztqCwwNtr770cX
S/sKpjcCRdI4cetStaDInIXW2r1a709kwnAgbPTAM/siSb3MNKcNQO3+CTj121cH
deQoq2Hm8VAjBkz7S0Vs+lNzV5566NLxZqyrp7k0JX321DYnu34zKhDRh8aw+cru
j2tkBEs5E57FbjJ814T4W9ERMQWd8Sq2i7ogJNgrD/MdClJM7L/1NwtiR0fn+qb9
VBSzqNxcn5EFELAX12rBC5Kin2fpJ/7lXZ8uZ0dqIwuMr/VF0qhFjEovF0wcKT97
kk7x+5qTijwCprzn629or6h+R4aGgL14I+G/b10CstK0uKzRi+6Pmme8o02omsX0
5iUvKHxexoOKf6Q0Ku6g38YErtDCxHE3AWMR7crZ9kGWeWJUYRnNnrp73RNtfBT7
EeoTkr/2vK6or886zEeLxidn1BfZswbKgnE9ogiI/0xiNKKbeDTu4+wzB77+R3Nk
bT9Yrlhsb7UM/VcmDlqu8t/PBRM5WZPdJcPOz4+L4fiXW2ggm4raGg97ngrAHMPA
w3X/wZLfVMVedbIpmUehhA==
`protect END_PROTECTED
