`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
krd5/Ghgmu2dXq6FqkOZ6tsDPoDFsaHYIMnlnzCD0YZpBsKbw8BGh9wYv57Ui3MW
L6pGm7KNo/iRshYLOqxmQc2/J7dYqTDt7jBSLfpfnd1Bwm+eCtpFm6badOsyxr8t
ZO/euk4Cn46h87XF99ItQgUGZ45bLtjd6T4MHDGURbR8fuF1J615wpGpa44crsdj
x4D2cKsoyGYry7uvuA+e1LFTIuUglu7dflfowTb57O2l90fxvpfTvF0lrmKILLnh
hR/52bGbx5qy+eDZfOdGxWdcWTUvLL9lqBLItO8gEf97IKkzLGAybw+rvh0KX973
bVft1tnzd39+h3B5CjYyS9DgrD8/mRKhG7/E+xQnLxP/cQYxg4/8DyV6yVEKpMdw
6/bVNMpb5r0xO7AQR63nP+NRNE8BW38xsDeFYMqZLwYm7odHeq8V9HMhmOpiR+hE
lS7BHLCpg0pAJtoneIej1QWl1ATglfZ9WVlx/yE+AJMszZadNqeK70dmMnACDIHd
4zG0SavbOqyqjgjO/VJnlhYUOVMI7nL1JDCeFCZ10gmiJ33zxZ9kBti5Mbqud0Qw
bFEc7G9zNQKobcPy4ABWUjfszqFqfJzlWtC1n0yJlFZBoJmGGhmgQaf+cRf8LMdp
Ndu3JCq+tQpuIfeEA+cVBw4Gb05CaCs0Ivgd2c/ee0PsFPiHMGjXqWBcABjeJzp2
Jxnky6B7OvdYZ8pBGTOcRijxaJt72C1WIpL+MjfeNzytHnTLB4zhe51+I1XZqUVK
URCBLeHvdyc3t/Yykt98t8pZ+b9g2HZfbIeZEuSgnmOj888L1pJHzYibOn3HZ28R
QRSpvWve+U8oLKxLIhk22Q2MX5Nf0RYfDxRIgxKpkgAE/UdLKRuRbm24QMfTfysq
Z1WYGu+p5rBy1E10FqqZ7Wv+NgYkX0aQfFVkdAA/AI15+OAkxiGG/V7WyxcEbSOX
PyQkVK4Zqzpv+R2/vifrox0yrJEds8cxF2CvszEhNXOKAG+HL/DIaNfnOjB0+Wgb
XdCSayuvHeleS1BypC8Gp4JQ0VYN0Sp/ICaNSb9tFmSdFvtWkdV7MvSmLTlTTZ5k
krNj+ZFQ3ItqbecPoYwCPvHTdIFYxGugRzjwVt9hL5TFcDYJsX4Dgf8SlkpBW46j
v4h7IGKMQWGF+Vaurlb8N7Yx4Lz7I+/9njWWJ0MdRUC2YCrkojJKiy4XErK/VtNj
j5LpH2lEsFFYfVsHNHJJ1Wv6oNkpBTKRIRJxIi0P5xA/sQgWTZBSuEuF+kK/wccn
NAOU9+6F9sUh/GgRAK3w8CjTPIGY5LrxrMmaWSxgXj7FZxd7CBxjC14Byih4j8wB
+x7VjlQb4beXLgXdj8Acr63gSDiWC2dwCazRhj4wQY/zu5l5hSXbRMe/55N4dXa6
/MscZQVjykDZA1/EheidVzWo10icEJFp3e37+ZFDBXZfdUo+KxUhN7U/Ol77CDr2
I/sXXHioLnQ7zH0f2uaLyp1hhK/B5OIyNO7tjXXvPCDJ9z1rmhjrOvKKujBxhT20
Xecggg3BRIIoehkN2Ae9urNWF5ziP1558IXw3iCjWIja28XfOSEB+J7UyttRF18F
nxLlxAfnFqL/tN+gn7a93tAHhdYv0XiYpCENFa/7qqw0taG038VtYELKV8euymOz
zqK8Mt4GBERK/DjmIS33hyVQKY31TdKlN0mqpR4Gw52dE88gnvBec9CKWZb2y0Qb
6jWK0tAXDUarv/GNbhoNNAHKOmQkepchOPU1DkRmOFn2jVKL/ptTTg1dCscqpnt3
O7rlEYGaFuhRjhvpn423HE9MKji+M8m4sqfwlgKgpVWWE3YNfNWebkNDgvjQiPXI
cRwCA8JOlx/7YYjA8MqoQ54zR6Cewbvsv4b8FlQt4qQvSCnLsY3z5S6f9rY84YkM
fu6jZB2Rt3s70GeK2/BfJ9Az9I6fdcg9N0nLU4QPh2JxigN+gXcDo2848/wQ7Xzk
BRa0KCLgrLj4+06XermiV2uG8ydGVNHQguHc56eC2iy4txpuLeFZzGivPfGPNpxN
Q548EjHSemAUkcGORR8jD39K4IjdepTtcVWIdEYclRHf8E5UqOK0b2bmy2FzZTq1
bakyZ03vd1t+N1ZUTVC7n3zxl97BwWiQdXYZRterqfjxBY7CgaJV+aKsxGulLEf8
HDL/aT57Tj2Aek/aOhC76V/KlxoCgJo+QobeyJHv0CZYLYpwStJkmE6dFFRyovvU
yg/3lPycWSuK9kJ3vaqKEvR+jvnrh+c3MiiTTC1WCZi2c2WhfxKAqh7h2mP9VnBA
dZV8Ai7qKhK1vk6pemf+DBUW8+Jjr3rKkeETh0E78dI5ILQK5I3p22/SgAUjHqm7
wssxruNDvFV58BE1ERi7s8YC6AEvcVOOYwXwTHMegKqRGyX/q1YomtBDzktLsI3f
iAcpWnJsR3iXpDYIiP2vSUVpV8rG4hMuPt7YJzS8z9//oBz5z05ZhbFglwj2Yewx
TnQsR88BaREf4gFRilTPKMGT2xMPUUhgqN1jJdCYkQcfuOTwntt7umWYTM6MZuqr
6GqMyXNfYDJiQdn59myrfbFacOKBTzC/tMXSz518HVNFuZwXYuh1DrEGJtEfMrw3
lIgGEHY8QrPzHmxeRVx7M96JnkvH9aHBBaFYPKuYpY8tVAf26tXqorGmgLCVGQsU
DGaFRSuQG2ExRd03acOnfEeOmSyvDZmn47NXXb2ycPO1RZjXSnxAn3MWuRpRvYIq
1a+EzcnuWWsxAgrEZN0agd0OqjyX/ep+Dxrxwh1KNIUXXg5tli/VlWh74YdSCbft
1TcFkES2yt8z7wdvMbE5QaRW4zAUW4psVnwCb114RAsY+M4b8AEZGcVOU7vhPa4R
invvMGzLcoD5QUys83Hw01ohWAUCLXO9shU9usDQSsk9jND2dD2RU58xz5LW2jmU
BvqkyzTPt77uwatxNpp9dIahrOYzv0JVSluch7zjmChcHMDLVFx83qTDTMOHOcfV
njndCW27LVYB84JUKvmvLlXQS/xIXyXkUBE9WXIDDS1PduF46N9XVpFkVkCmMJdS
bPAamxzfZKE/8ZKBUeIS9tnPfnZhh+68Qf48gtvXRqM+HGZfwMciWUqeK/dTGMn+
lJMTXRorQg8TVvsRf3LWPDty7mVIbHKddGowTS+3j2po6C/h6ZQD5c3cQfIf5PDn
Szt9RUu9r2+EnNfLyCjo4msJo7jrXC7dIe+CkvugG4aek2TInuZgBmLH6nN3Xf34
5V89bhV5XAQ9cdfHNEmP28EEb1QCb1Kv1HKzzrE+DPGlHWAPx9Lo1TV5a8avnKmk
QyjTR0RvL9QXLGm7/n0maKBePWv+p19W2tKxByziKlZNqCQNWfbW6Wt//W/CweT1
8RZUSodelOrxMmMXksxG/Ty4v9ZjUe0d3t1DZfejA6gLZrPKHaxiIbkD/GITMqyG
Htov5mn/rf7LqM7w3gVAktiYoafCEXpBrHjLfqDKOU8eLQ+3XQgBp17NMCdltI8T
zA81C8/fUnBR9RCPQm6P+KaAq7kx/3wI6chpM4kFhPcyR3PwChWL/bNZdHt1n7v2
psNru7U2GqRyX+4Lx5nWChDAslFeCQpkl2O51rVgbFm2aJsOst21CqzmkF+F8saF
TirzoYgzHLgFmqsuQDOJuVdh7qoJHhtEDllNS3Dx+HofebHDpahZF8Uc2dffd+/x
6e68PuXxNQOd2KHMmpvUPYISHda0fdnAJksrCvcwLNYLIo5qV0JMH8GNls6JgO8G
eD2AFVsIQ1/WpAwMwXypbciazn+C2B0mHpvACeRFD/f/3MDXAOiduQuAZCX17gCQ
UTqE6uFhq0NCA/ICN3AeRiwAcboxBpnQXuFfzXBEscpXq+6XYvLAB3bE5j2bBx34
/oFltcqAYhKd1K10QkQqbsrwZKEsTxOg9H9jfuYPygFWbE6LkJIaLjpiRKv8lFXE
QoucJgPlCj1IrVsMLy1MoFfNLWfgjS4++EgKZQ8+3IqgzQNfQojY42Q6Fl450+Ay
ZyL49DJtIsihG7h7Cs/VbmWzFY/taL575mozVyHERJfamupv/MXjXPdJFwwV6Oah
3mCeRSUlSyu6uTcufp5mBv/2ILq8vKw4i+4PSy+VvkCt3xBuy619WKRK4GCiHIhe
HhYvpPFg4uPh3urmh+YhCWMNBAf0c9z3e7hXRXF8geFjgkr1C/gokUhxIYy/vUzW
Thmr4KxCtILEq1cjxlL8Hnvai5DJM3LQ+5abEdGhhzLae96J+St3EAKWGn3zrFB6
9n6b+ax91rHL6cRqfdM/QibOYIIGZP9KrTjk5lrUywlt8EvvDyLhDf9ZcHCTm880
22IKdO50EkNr6gQ+f7Eq/F2qkx/Y3iztE1UH9LOyEgdcVLgxAA1S1TPP4PXQigu6
5l0JaLLWksmxyVVdeviMXuzRhc3OJHMCtv9CHNWOo3GWi0qY1KurVCOuL0FjGwqR
l1hME5wHs15f3hjqRIDkhrsJdcN8UUXPcn7yrLWYhUlO39HVYBCZ4corJI/gapjc
LPg7Nx3njGyXTjPJaIvFN8whSCYcic9LZJaYh58UpG/Bd3+PnTurjmfuryM+UjM0
Tw8cSEPKjZLDlAZ9HJ/ZBGvKTBNM+TePSAqtGMlqg5r5qbXD50YpaGx/KMStX5IR
xmXR9bqAqbX9A9NAlcETyEiI+cIcTKLxQ3H8d7ikxAyWC+7ElIH7avPpA92Ghqvc
Z699fabEel9fgSXIBkeR1x4qxms1T6qFSiSNVfeblJHuQ1BL1Maj82Xkr/RJHpsc
//lkWEMuM4db7sy/IsxPMH8qEzjJAs0f2V8IN6hgvSkzv4FdGM43Afy3mm+49WWe
+gkvwqf3jV1bT81/zuFEplEr0HY7tFLaIQY4PowYL1S/FDC8u6EWpKKvZ4PZpBfI
0yilMJcU5aC6cIlvsGFlyASpq0wZQbN+EJLwHGGKXAvBhKNXevqL2LBgiZWE+fVs
BVi79GtxOdWfCiWJ5Y+iY2vvqGRIasuHb/gb7aFE5bhX2e6wZ25hNZ7kqB+VMjE9
R3SJ+PMWvJqntb/XTBewB2ED/YyjxmaoOFkOYTooQN31LqVdd6nb5Jk6SFUNjj0W
aWhRmOBdF7Eseev+vIJ4SOhZdZYT/DOHFfOaUTdMoiGvjluyAJTYOD1q168Q8vfR
pcSxiostqThHdIx0StDEjdZ0NMwHsNK9D1iY0/S6UuUMaVSTd0fFMsqyBVJwe/dC
gxatpMGET5Dg3I+NkGsx9/BSj+ACBpxGlkxX2ZoM03gDk433U4ZwtUtJKwPjdb5g
UpJXmSndYv4VOib7giPeUndMd2zfF6vtop66xP0k/1VdFykHl7eaq+8xCKX2T03A
vr+xmz/doDbUzuzW2FgVw+R+e7FtzU6MlmvswJwvmZT/je6HRUymlIcdGe2cUjbD
`protect END_PROTECTED
