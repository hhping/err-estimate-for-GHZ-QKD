`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kJP3A0M5A6anEKt1p1Ek2LyTJ3GYj3gPe8nGfinD6lYxPl2zUPZfv++H8El2y0B
snF+c9ZAChMNCK+/yX1TQOhDQv0g1eLk+8xCx3QtYgPbZo5mKJZeT6gaP9vKzh23
tqOjYp2kcO/RYG+NenFlA7TMN1QkBKVZ1uqdOTHhDiP57OirNbMxkgC7weQphf7c
y+jYIF/yRsrTbDq9ZVaVW0KRAoS5ZEq1HD43SY2xQUvh/gnrW9c4ij6TKqCp6HvL
PsZM4weykZU1E5cQSPxi6bEUSqJTnal4yP1fdsdet53wllVq5xqBIyLL2ghmjkbh
S0rcl/Vyyo4HwvsIcEnCrak7N8gwldIUVdGFNhA2YJiT1R+/x4D6L7BN6706f8jS
FkFwWlc91Oq/Y9xhiECSg6oNa5WwjmNmLzYagEbEDrXCKBq4omTdu5Znrf45MVVF
qOLIufYAUY9zRnaxYFeu0HThyW9YgOr+ZOjSK+VLQ8sEGZQs1tr296HEsgHKH73W
HrEfDKyGeqbKi4Qub92xrb23Fq1lP6P6H7/ZUTDNMFgJCUORcb3SjGI2rnnKna8q
DS10S6V5r7Ji1MEDChCjUHLwke+d2CpUP78Ac1++hKKgYlcw/kTobej/ZWo8NwqY
+GQNLAXipkDI3bc5mzcrf7hHeLOZbcwATbzdqMqScBGPE0WGn7sICqDGa9MYDWiT
ufCC/vHLR/knYfNubsTeQ9+39475/hUsJwq/agWhsfjG23jC5ropZ8gmpf6s8OFi
NxtDGPbE3l5V7WPZ5QThmFOsbM/+JDbgF/YIdLAaBZdi70p6HkhCDnXm/lX1nDYL
7sF92oFXJ7diJswWvSiYiJ8tbxkWxMwV7CwmRCFGCCWzMv2/QdoWiJjsDipEINlr
7cFBdOQ+Cq7555S5qzmnubIXReJB99jrHV7ScybvMpbkXc7OUTbDCJANGoW0UuPk
r/wdWbpbu+XxW3loydrZFh9ScW9Ka0qbBJ8d+bJ9lVI1NmWYAaNzgY9JRDlIYZsT
sedlK03lJRQYsn911jNtkljGAmcTc3pX2qBj++hXlzaAU1LU3/uLZzfhx2dsjMr6
+XUN1nRMpmMRYEp0ShuEFTFIo4vuPPKSV9qq8iNHRfLC3BCYcXsZZgAzjzwMDQkM
Ztt5biNkuphQJl/CJoyuOl53sSMXYhnGiudJyHGiUJdBiiywxSlPI4tr8gowfObj
c4zmq83cR5fboXzw0lsS3jKsJhsqfBZGo/+V9RYyaqcjuzCNLlONMY3NqYS2na1/
SWpxkbDBnKf16VhhwGFKP2BsKxBAd2W7eOPOAMgP4bqqNKzSxmE8xYCYfbeOMyPV
hxxU30t3HnJtq6EprITusJ7YrkdedVxNvKlB+bLc9v4xJhPVcogt6ETMBc5fUTHr
5RzdpuUGw4FRJFs2+z/k7UllaocFeGLMhszA5h4CQs+E6N14QyJBa6ihQRfomK7K
+DGU3IpTDFhvRtgZRrcrXs9owChDcsaJXmevj8DwepjqhjkgItuEf9g/35k/TUOM
tHM1P+MGt6cCkoLoIou93yP+pbeZBuGopOdXAy+tVXs8ILNL4qBKOn02SdYiASN/
SE1/F3Cx3palFfjcBO/6qCnHG6Ju9yWlvx2li3BlJnIN9xDXUetBC1tzNNSaqiAb
wsJFzFqbIQ/NNHcObCrUsm/msb3IWYCgQEmimYPHWKWgRPNMNE7/jeFnySLGXkrV
G3cN0Ir/tuKH00ugcXzQ6uU2aQkt1lPPoHGFmeJjepv9vNs4Vy6fpebYpSUvU1Gv
cdVj1Hw48hVTEjfVr8TeFmAkb5d0d8kNQYB+w2oBMsMfYnBcL43FTEUYu+Ofy9RC
APrjWvxa+g1ke+2O/1RnO2kUmc+mAwbfSiVNDq8J4U96zW/JqB9xXyeZcvRc4jSP
vM7OZujPH3x2yMvMev6NLMOmHJvUr2ViyAoqXF/nPnL43qrr6d88pqjqpKN93jAM
so2R1YPuzoYLthQknK4t+YCfdWGuDi5LFBY0SglJlo7sknG/121ZIRqlkwOZpS47
rorg4HCgW5Na3XfUbrjf9k5qLFM1JIzlgQh2NE95Ki31hyXJ3a2Ay33SGaSv8Rsm
GKPrYDaLuxAAerXm9h1NbOxHeV8H1OJVIqArBv28gJiMqxd71hMTSCtiXnQ5pONK
JuhdDePhY0ASHex15t8grWWlGVsk0c+LIR2k11LzHHd4awfggn/wLyLIEFqUZELJ
TWGKZuYb/Xeh/fVDipjf+YWox0n57FiFxZCEY1MwpygumdX6bU7ZpS6jWhkwKM4g
8l54kFaUbtBfuMIl3zd+7ezqZqjpozkZkQ85AZXOkCrQECstZ+Zn384aGkIoJW2O
lnPBG2v5n/ZXdnUADeKJV8is5MWa8jhPsybv2GK9401aBnjqDa6+rODCVvaJBm8x
t3/YqaOX7Kf5bfVdISucvB1dJgLgs4pX0hXo98FW6Wdt31/BhNl9afP/QsN42yIe
Jy74MBXEcvvVrcQFO7YR66bk8pJ0NbLV6Lbl8PzlypeGVwlUwPNbZyxKqc3RQX5U
bzYluD1CBhoIL+4bY7zvhIK0OLkKmy/EtVY+cnreiy/jO3U6PAojHSemU5CVn/ic
6bUmdJnsY2s1Mac3BzozwqblbOETS97O6HQ2LbOlWb0FFXsGWEMylkwe+70VYRny
1Bf+pHlM5aUNASA/YHe+aB8bXtVoBFM7zx7Fh5ab6IooZ7Tn/jNPbx7WsGuH4iS6
bIVhfvQQrEr7qA+mV21zzVdj5U6VTjElPiOyhSFUsf7SZuVFCijc44jDAxnBwWni
bNThtVQqcM15TgH7wV5dZ+YeYizT5I3V5Ce2BkH6KwAdtN47IqW2osoltcKvBtfi
ci0zGu3ntRI13eHNwkCbS5VBfZQbGNCBlGj3D0WL+otpt3Masl9TYQOEDWhNT8lD
hXkerpoO7malFo61nGBhCjWX5rDkhB8x/zlXVthrTsr7JnYrgIeMmBbxbKllYmlm
T104NbAljZJItPVM0l7/iEfOO/XXtY+Z7m/YNHfY0JV7ZbHPnePD8R1asMV5Cmwq
GZm+jils+cR77fa7sBmWbV+KiAx/Nerk0pmU92FrQ0n5gi4CuQ25TeYy0v7bcaxK
lHD23w8SYpIE6JHtQJ43/fV1H0Q5QwnKmy6J1f8XpGwe5vRr+zONwV7/hzc9+5S5
sRXiWhs7qL38Bfpfy0ClcndxSCpwsN3rdCa79Id1ZnuYAndT6z32D1kXeo6hi+4g
vR1wuDpp4cEmG8Pd9lNJAB9bKF6s/QxSqvMx9px1j+ydZBUPRvxJbqqBO0o1MhJR
iVa1Gk9c7ZqEp+br2bJ1dC0vjnexCMoFJ73EEygnzC+0IcitCceZ1H8GpJnQnYTK
RfZOkN2KbrvN6HvFRRg+OJctURergmNunAL5X1MaaCe0nCRJD6cYE7Pa9HA46lfU
QxPk/CRX+ieFwGJm3zZ2zuJ4xWCU6qW/p8Erg/Cx5BiFxs/onnFRCn/nzJ+Xs2KU
koCPWnvNpTG0UrahPixDiqJYWkWYIQrAIVo/6N6WrNsLeyOPw6AN1C1DeeZ1hw0l
/VpTXtt1FKvFndywd5wBFzhtSu+LJphK3Mzx5DGmTatTEpdj0PQMebd6K0RxSIH5
wnnhJDAfabHrXihpdvOCWCqwyHbikBnwGXwKrZP0CsRkHOe1/4VFBzc/QIKVzeGa
ydy+wviBMxZxZCUtUNJfmgNt2bPlNE+laBIE/G7bqYCcrg9/FCxro2d27mtKStHn
ioi0CPGN2C+ftCOM/hr6CKc2TGHdQ9DAM3SELuG/WuOX+eEwPIG3eC6L5vV+tYpP
B7AB/MNbKXNxOUg/R1jiGm9/6CkW6asQP0uIESS8732TNjPInYO7afdQqwgC/VKK
1JDCDiIRPmQeWYRGbtF5SI0qrpN41wL1SfPv9wfoLB1QBGq3k0CAJn/pn2mFj3YV
5wpMTrvLo6JGM+RGKMR5NRsxgY0/PbzmYliX/6IfZeiWrRnTfoIEfx/ygpuKigWZ
jwe8+TxcrymgcxLoj02qDJIUxU9lJdRgdH/KaxGr3L1iJzpcN/4aIDFTV+gfR4vR
2GKmtPny0SBTHqv7gkYXtGmD9c3n7eU1GmSsdheighEVaReYqvNs4Irydhg7FfC2
lm0NDcTTMQXSzUKw4bKgXo0JAP1zuLUGZ/Z+Xg6CesH9337032hTegRmNEQGi+jp
51mRTEXvNYj+HSJ0x1cuk6hDAxUmM5WOcCAATuvaD/a3wCL0WLJ1yu0hTdQzY5zo
4gdK/PBlJCNawwhmRzTrPqP6f/Qsb2WJmDEc2fCPQy36+YZfHduRC+kLojLGyKz+
JV1WJdlxblVJcvGv3DqsnG9pnyb2+cX5ICjcrck7XI6fR38kGXJDpyiIhDLR3NOE
rcwnE8XxvLk0YLRebdpWYS33IPtvSJbDMP+aZYfdoBUahadYA/pkXnes1Yg8++7k
Q2YTNIkFBfeqAoTk6biQeO7uwT7yBzqgAfDlEHnWfXYz7lbuL4VKniLKNd6dwsU8
LUv/Mp5qpgNWdIhKxXIVTpn0PcUBFo/7k7zx39UzCDImEpj4wW4iXX4Im5H3PkZH
pQGeq1M3XiwQM9JNlRQINao6YNIYnjuL834fJ5UjpJBc5Vwqs7bGGVpuLEkrftdi
T9OVHCRNjiJ2lCdtm0wjNJs1HZ49YHZ9bRzjBCNrTii3fJroaXBA1OGAkHUtZQ2K
WDnyGu8mabvN000jtxSx6IJia50M9aGaeuhclJ2WiYbewZHBA9K/+COAFiI6yLfB
ZR7gLeXC8O24rQhbIJ+ViZ/qosZORW2MI6yG7TR9oH+tsxly5CFlmHTDmMj/21yv
2v4/2brjjQAtBQpJPMJ/NqcBbTIOGmQFVHFYK6yYGzkHI47g6SdaoRv6Pc9cZt+G
E0syYV84Xp4+ABDW7Zwvje0UaXsz67PqLvw3cgVVajQ0R7p3zfv1EeGvEd3jAYjy
DGUFM+UJZK4C+K9KKZKi55Z0ZUFn4bJTvJKp9tS/cEH/cVSb1Isf/bgmhs65sl1N
8jyWkgqw/1mNJIG8ITCvTTw9u9SiYoqGFTGkFBjO9ljvNmn/b14b78pg2xt9sylP
NqZAIUPWSpzvw6SVA0Lu2yI1EAetl4XdclZ9AxbGq/nlT8aK2bnaCOzJrqX059Jo
dpmkz6ngvn4OWsdB409J0NVmwNCcL3iJruZ22noOMC5kptbf3l6I/7nwcYurjeto
igTlxIXk3lpAl2AP2vKGkrrZBJelX9CooquKifLno9WcCIWgN6GQ20fySaFRlmv9
nHKyblmOAoVQnmss0jIqDrFCWiNWfycxqqL1n59HANR9nNGtnHAqv236hLaCOVeB
6lSOzS+z5xmOJDyOtsLfHpiFXC5PPtjdCY+lBINjew7ce5jjyjRge37ngSe+A/PU
FRPzooF/7zS0vDGdV9RUmn8eSdG0UtuSE1QVv4AGilG/ZuUj34D+KwcizumZdXgT
b5U48tvaVWfDO8yhhpveNrIUwIL/cTq/U+gxZ8flbhL1S84RUeb5teMXJVtsEN5O
1+QVUBln9WT9fMkje70I0NzP0gb/OGMrN11Sp/FIVY1wOvtMlo5GeRy3f/FhOjyb
aXZWxncCgeW/D01qXH2Y8AZlzaJ1o/m177sW+esPe3aRE2LzU0oyRwZmd5/jXamO
HrJivIKEMGUakrunsAPHUMjKlY2OVntOdvbg3WDrXCv7skPj8kFIoeDtlqzg5PyW
PYU1VlaAjhjyRh1OL07ZhqwQM2ykTA1jG3zeZrw2emGO9VJGF/LLyDVg2uWdDyoL
bp8kYQZlnavl/IWWB6r+hV7cmekdpkgkeEprS+RAg6QP0O4yVZRrVwA33yYdkZ71
vvWcF1qJoBnY/tLNg8Sy4OCllYDssasvF8ePA0VH7ACnVjHi2qcp3qzI2Z7KXUEe
oL7UjBhLChGvuD+MG0+BYNTo3By7xiWCdE+O07IKuZ+yRWq07wcWAnc9zTtoCYmX
c6GWRGy0DyysVqTgxQusHRtVmZskp2Yb/UormLEEUgR38SnPtMhx2gosY7E6UM7V
dIeC3yxrkukpNQ5E+eUNViJfsRuuC/QbnZF3DiB5c/5uY7f/0YUqEAjiOp2+TE8P
7Qqa6qnxkQhLWFobViPu1KpWCP+pf9gwsnOGuVy4CbpwlawS9UQcv0u+ctdwaaaL
3bF4NvvJ4DvgY8lXv5m8EGxez4T+TJKK/PpmFz6JAkwBOaBNKMxCPqpxyht8wvV8
8SyCaGaXblftSF0P1w0lLKWPicmWLdgUtSisqltzn5dGxN3pe8ZcQ0vgTe8wjZ+a
rygOyDO0pI8lYJhXqUwVnGttx6hA1iEA3o7adZ2o8p+8yx/fC1l6DtGuwQP+kSn7
qVMLZEX5OlFj274mNusfANqX9eDt7BfIuv1+jcuAc0O32NErYmZUuQqlPGcUoxCq
a+fVJhPe/8rvhYkoE+pjGWUQC9RHt3RDObxd3h+Gbx3McgbCuiT54S3f6o0gNRKU
jDAzQ8sfSkc59PqNikfz4APvRvkHRlgSW9FvXSWbt8kn5hjD566U1TquU1mP/PI2
TzM94ydfxdTzSzz9FEWywqnHoJigvw442Xak8RHHyDqJAnyBKJIJCF2HnputAhxl
BI+1iEF5eZMeiAWnFdzn65ssPakUmgLhTW1fqGKmNrK3zRZMq7d88SDJT1NVJ5FZ
SNgG4OWHfBuNsffIHToZp1GOUc5BsCaGjHiBYCJh/xxGtlALFfhHXBjsIgZeshJV
mEX9rRY6V2xGxf2EgdWetUplbBc7hIy3MqopH3GROYImX7Oo4LZ/cHNo4U+HzDaT
pguz7V1jKTBJyb74Zph4Y/ZSWiF/96iHUNGX5NACjld0nxtiATaZtyqk6LseY/Nk
lHB8z1wD/DznccKTfYoZJiGB8yb+20r4bn9gsB1FcJTAvzanzXhVCXogU4rdOHLi
ZopceQNIS8c+uWIw61r93ELdlNamuED+hlRFBS34GRz01OlITySbDXhGho1Xesht
/1jdg0OxxGMcsXvMucW4fhzA+kB9vH8TXEI+sIOsv6VgdvjlVw7JLiWqHj4JQc1n
z8u2NCmSLNF9IHHo9qDP2ZPaot/p4oLTu0tc34KdZwWsmAMNhKkaYMoTNHMZuMSx
FMNcL4uTfm83QIZ8AHRYpsGpxidrWT8xQ4pASG1W6VzI8MgpRYLLcRraTiQo5r1E
JSDwdB6K72ABAvMcp/BMQzgS/TnriGn1KJtchXIyqSTGIxOBOHP0lxdox6zlQQw8
AF7I5l54nGQPELD2Iu5jC46DH0BLUY14F+csP0fKfvPQv6g4X73mWBnUsJAiOcGi
4KSSx5iO8U6OjT8rb6SwPvSGTwXH9RAqfDgDc0foS6LDEmeZ9FH731a+6dxGYX43
sHIL0FGOfUf5smhVCqqpdGnMYahXZ2sWzIfmiuaXFOyMDti4SyEiJmpUDg50x/HA
KHZjRelLRQkccnCy93S3HgbLWHCZiD5es23rDVFwXWzPpTM/mCX5LBu/Bu3LZIUS
YxFi3aX7j0OKePCq0vVMFcsqjkNhRuGE36oVdWxCVpt5vId5JFIZxkPhR+UYfnH9
I1vWkpvBVhlecO7QlADnAECKqcgasmaKnjMLLOVrRBYrwqP241I/V2QPDrcB9aUz
X19FgMU0DyzbM3vTkcl/EHFlihhKckaReQvYnBvbLs+X1kJpLICCayWHf4q5CC6D
chMRQ1qo/6kpkSBVAtIg/utVTPGCAg/D7BiDdrgNbf2MRERSk+qnW4SM5IjYrNwX
yyj70YEtOc1PfXd8jnpbmw8pqlK+gSomauK2v48GwNxETZ/9waeAFSM1q8mHzqd6
khcqb3qokfbfV9DjLE92vBI08I0zNsG1s77TA2+p9i1w3Y3SXGBEk9aYLz8K2NGu
MM7s8RGnPV18m/V7fbvh5Qo2Eg4IigOSUsy6XWIrSSrsLIe/M+wTLWE8aLzwBjFB
uEPkQ5anPnRLBOprP4fB+lur9IHAEHJiQIXTxJ+hbsyZo+IpEVUJE+ZARSE2z7SX
dWn7wCHvryhdUQ+fi7AX9q+cWcWP0Ixz2qVpWL/0c+RJ5a4u/egHnIQwcLAwTDe0
ZhxFwHwKx9CPbsob7KcMHMy/Fk9JwbgGLZAVTKIsGrv3Wq8m6426hg1A6U1YxACQ
e7M1XjvLVH9anD3bxLmGMH+8sRcAScf1s5+UPf3EgwidyN7SWo4AQ23q93Bg0FpL
Cm8aOMqo91uaKpKucNpLy0euTOZUPh4aGbucvtlopV9UghtzYLt5p4JhLGS8f3vx
h7EVc6u/qZsFoNGTZ0xYSsLlQUKGW54qLev1BUjKpFHLkk35c9lSsf+6uE4Vg4aX
1HOZZFA6uzoTz0ok1gjI+bykslPfiDtkH581IfZPTKFWsQpR+kGIeDlm0WmWCz5N
Eq44TzfWWJmk6eJTAO39mw==
`protect END_PROTECTED
