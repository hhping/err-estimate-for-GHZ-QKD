`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbzpXxAvHTLH911ZkRqLrTyB8XSuUUqfXn0WiqzmKH2SO2/D1I0nqsxtg4x2++YE
DNB8GAZSdYBDyUqp2ETm0Vm0gN8ssczWkWP8KNm/a+IFnCEo9srGlRUApJubHf1r
WlfMz43U2ySJ6cDbqmeItIjF/VLvKyYffr60OyjE1KwNId4iqkJM7Ww6n93rtlDK
BdkQkgv9c92+oXDoJJf76Xw10bOzRf0rDnGBvIoX05S/NYwsSbdBNHiEhKMNZ9M3
En1plHTwEseJ3rkHqGLSqb0RjkIE00nvHs0Of5JsoPOSwwYz0rgxDeJTqe639UYO
L8Dzc9JBHnNx8HBMl4kEk+j0igvln3dDvf6xPBSaAq5Qnnsy3UucuZi7VgKXIhuY
AqtRhaNBe+PpgrwrixHDpB/koWpTvf/+oIMizxcghv4vheoTe+1KLuus0GoBWYTY
QF0Qd/nIQMiIlPnJ/Z/xxGSrVkk+hcxsAaluamxVQZVq1/WwVPbvGclBdcBvEfzT
m3F/fBtz12MoocAKAESOdfbh0L5VDliTLy5sWJwJxKQYcbcepb/fdZE8A4NImetE
9kgsQ9zN5se8YdWqzwRwZboiyz33ignbl7ntEHoFeUihyfn5/ACJB6FY2VWkSvTG
MvaRRoR524lbZxNHyJPbRC3fZy0N1DvXEyOUuJIuGH+9Q6TxQMtRNJkASIZRvYlr
Sy2pgOU4CnjTLlFm/3BBFPakGl5qAWDoWSuA3wow0OwOTqI6POZ45IN7Fwv2w/Vv
`protect END_PROTECTED
