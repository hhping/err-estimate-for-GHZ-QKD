`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CrQP0a7H5dpb9tS2RBdwvk0tLJtXpaLS02Uk0FdME2iLMeBc8sfQkrkIEoZAlPtC
UKZ4qL/P5z3gj73PNJ0yxk0oGopUqKmSBRm3H7CQoK++YP/hcfGcAsszET5hMh22
PXCufYS2vmOpZHZj1lP5qy5iX687vXAd4WE7Vscji4xs64Quz4DsuZ5+cjl4j1Gw
HHeWpGg5iexKjtcRq00rog5s4fV9FozmoHJgU2VDX5JOqOYNyiaOYhR+PpYxhWsw
+WaUjEyLyeDGTWBXe5xTbkhgPyt1lUGGKoud24kxyoZGGpQXEdR6CsBMS0EWpDN7
Kr+BmbkgD+ufsbPI+F18QJxIHJ45iOCPLz1FSGgP1aYhiFJByQwzNHxHGoAdpoqC
hn9NrrBMXWKZJ4mI8RqOgi0taLTg0ocmO7GDuf0cDvjm56YvWziFyG+KkuOoMwVm
NnxgAmlytc6ZGLDBuzmJR1IvMRRcsg6GwjQ34bbntVvdEsDnXIxDIPHdq3VDmvWO
29H9SJmWVbzpTvIZy4awy3RCTPn9ld9L+YRDcDa7I5reXA9lDXKUszAeBX7JZFpQ
HOecesK+92/dvQK2QuR8vN3fqXnXJ7c+AQHrJwob7ar2su0ku+YMlAgWkshxumuN
PSZNBNBIRcPqxsu2dvJxa9W+/rz2dijQ9vn1kcyrhNu8HjqgUwWodfTEvP2A6lwz
MLMSdxMgq2MFPVQPJ5uqgg==
`protect END_PROTECTED
