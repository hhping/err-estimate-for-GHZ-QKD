`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EibXttmw25VMuxqqIBxC3yWqCh/LIwg9PeiZ2w1fIRZaiquADwn+nhlY3y+uOULd
dmtlG5Rh5zAqAyk14mivQ2N4BBNQB2xX3/crRgkUNM6x4F+KrQUKmINXPGyxae+S
WfmlquNl6rF2zzU33L7zhO59fkRgS+kWAx2Rla6/2JKrXgwJZuevNa8neJ8/aL7T
vt9pc0Eu8lhLxbuKjn6GY96caAkI9xraz7soZaytD0dJ4sbf2cdSGZhxvHQ5O6Ex
THJ2qAG571pTYvBExEkrGiqjxLyUQZ8Un4u8nVfubfrRvllOrGLmxZGIw0udI3Lb
04bQd8qzKxqNrxWLsJT7yhSSX2o1kTR2yD0JO6ZlC/BcJXlaqfQrVndXQGsTVKix
ujETWQOOTcUa5YjQdYPEPDDy5n3aAtuCHM65oYrrPMywcdy3IKulFIp1dzkTc0mq
ZObkEWCpePYVmeL1S0lCcv4QcnCvrimdQmSHYQ3H4pBza+2vEUvqjd6830YGikA2
UBUA1dr/stWo1F4y4ZY1VFov01ZaDva5KNL8VhmkkN0rvxSxYECCVsgO6g0qFJMk
jHHc9ZpRwGZqJAQdawBaaoo384HMlWdLstWrPF0LsUtpdSZWRzYVmOJLryFN2EXY
DWdTSaTyfm7+nL0WpGdl1DVOvn6b0U3hdlSPfwriLx7i9/gKR7pzec/FNkbzyx8C
6kbcTUA4Ti/wj1H9VU1vD1T/gJZmsoyOcroPzLAZnZjNlb52GVFwSEIrsKU8o5xN
Ti3WPWS/gAqLGQgmai4Qbx68rv2C8L02hmugRkJHQ2UDhWcs2tzyPdAug3FpaLde
erknDRIBro3ue8kdlu+4QaPtl2WHUMgKy1KVcuIYSPXXWRqnpTCz21QlpaC0xhlp
BvQsN3NHVwH6kgiIBMULHP4S6BYHl0mQLZdsqWfylueD28T8DpVhyetu5Jp9SqCq
C9q78cX6QCbrbOewesrYmNlS62BY6Oyq7dNmA+BScCqZZ9hFdjonvxJZ/XD2GMbS
`protect END_PROTECTED
