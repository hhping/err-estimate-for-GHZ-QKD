`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypsBPERsp6pxDmhenynfL3RmJGdsOzn+npNMa395DzDHxqXh6hcaLLD6Y27v5fJO
+ajVp51tJLNylgYZ9auwmKuHG3eWDyeBf7/1Y2Fz94xxRTbvacS4BHCSd0OQ5qxg
HlEEkE799K017KcbyF8w5IjJd/EN0IazYa8DJDdvr8y6fqKL04t5whTFSLV3ke1f
bMKg4KtYfWcopJzpEXFOswXb8J/0OgldZ779FssEFB7TbaAv+uFP8t+MPwOehppK
qeawd7QoVCqpsK1hlaZ7D1FdxTQwz1az+3WOXPXhv2MdSDpgbD3bbNpj+CrxM6og
3yyl2WgW3iYEIfMgGV5RAl5S66SKHTD5F0uZLfXugTqg6z9M0PK5eVjaHZN3xE9g
i1zRVeXFgno9wO3WQmm3w+jAUxG1sEsjWbPTBEbdSpI9bS50dVeMNju0C5PCC7QP
g1lncJ+wS2dqsIC7av/Piu1SuchqoRh7GXeHO1s1AzoeYaj6a69O655GBlKPbxNb
Pnyp1yDqxVhgQzGMuUijNdqMUYKkKCKJvJjjxkjNTvH/y56VnFDeieyCk8bEabPl
scVDGMcdz+uRbtVnj67A3woP2Yahmw4Qy+USrZY4qdygXdxDpIuxNSVsd1WQMK/t
2HFWhazEGQ96U1XPX1lHchm/w8ljtTX32t4XxCZ5/WVp/rOgFBX0Tlj+6fDSuF5y
Qhh7R4FrCsh5U7kLmG4WPE/v+/sWmWpWaIz1xdSovI1fwL7Gs86JCy6oS2b9t5sL
q6bcXU4xOBwlXMU7qQPVai8mXCyS6VHyWzSdysBMpoTB31tD9x/In1E3gaHXX+/d
UjDnX2KA+fMbPCR5tSGOWMbbaC2dnb/Vj6Tns1XA0oa0ypwt0HzU2xwKoGgJ/XQ4
b8uSGvYa98bEong72zvHTumRJIGDGDGp4PmRDF0mONDs85Fwg/g6DDaRz32BOL81
s2XQQEb3gh/cKq4TtlRjyg+Y9UwqpiogRTze5K2zATo1OeJmQ3uvPHnP+obKOEOm
AJlx6tzCAzudUoZFvY8QhhrkLR5OXL1YL2ph+Ku+ppRlN0o3VUlJNnzouvmO1TLO
9+bWyH7sHW5a1M07Mb4NxQ1VzYsTAmCyMMk/GyykaiYJiqe/xUV4qIGbRA/MPF2M
/R8fn+sTVkNc6JxyMNmjMqlfuBkn3bW4/t6wY9KWCjH5PC7A3BroRzh0+wKgBpYh
8uDscfEVVARU3PeyX6QOlSiFvJld3pXlNboWMCO/A+2fTdT93llyyKh5frqbnsXo
FuXxqrxswFuZIgYIOqVlHYuKhTy/zw/yjgrHeT8f97TdNP4VcpdvN2o4J08KA89w
GDMEyI3HX2sHKWvXzvSKmvljmo+44iDhHdE7fHzMFx5mNCEl5pYqsTrPJp2vG1La
M/fzQ7OF1t3OxF44P2XeSA==
`protect END_PROTECTED
