`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1V82JAWZRcEM8GujeR0l3HCQW4aC7WGB6nCbH7gnQ1vQ/d0KJa2rfsK4xrhssktB
cAXTh9QlBfyJpR/alNWHbkF9aWxnFUCRY1nheNLb/RxssTL+N4YsImBtHlTahOv2
zN1Mvk4vvkPGZFgEhiP+7ROroQvLU5rA/6LvYNIoODuasN6NCyVn3WBUCHoF9+x5
kStWUJMvXjio7dbIaoTh5UD8nCv4HvOlzEAHijZxxDceJaQ8ieAfM8092+kTWrFk
UsLMox88igMF1DoRcl6N9E0TVuk1HZdbyzVu7t/m3EnEqFxY8x0YvywhoDW9iuCl
FCZjVQfUFhwmELHrdAnqROVYvAfph3oWO+yZPCMxyZXfWC900hao0b62gP8IRMD5
s31L65Tmmqz5LLEMEMBwu9Tfc2y28frtUocZb+1rhgiUChw96hWRfmaBVT1007TP
2SOUyq+1jLK37zB+uWachRT+y96WCdcHOGuASP/hEownV40Riiedr8PdLQ045HQ6
rz9raR1HCtTaZDv5pBhZ/ol0DF5WQsr1TwaEAFUuMFCD+GQHS62AsHY6IYFJWcoY
E8QDrKa+w4TWpb1nylFXxpK3CKnMDNgo4/4siUmftlpLAvY7ExFtBphTBBYqwKl7
XIMhMAArH+da4DAH3LQ06K4gWVYrTQmFENyYojuSDWqcBrJOWpZc+H62yllfAje+
DUxeaLuE4iWkf00l9Q6LgKJTs9+TuoFdtkVaE9lCHqTiqw8WZ6EuL7TNeRqtrKba
mJNgwT5ZIuiPLf4ID66MFLJShM+dzBLimCdH/jTL2F+bYopapefEmp4TDaLWpMeh
YSy9FObJtO6YbjOcV2Q4ZoAmR7pDpEiC82eG667Bo7HcSG5+isWZ9dIlD06U7msG
+ccqLuaXv1XMyXsKFS+uT5AMoUi3PM/tzY9hZZ3qI63EINJsqI2RevDYiWFMzc/j
CPw8phBdOsVAlPwV79wpk+rGT07tBd3UlDl0UqixhRKDUei+6/ENQmlqz6OnayTT
S4nZwO+JeMUMCIEIST/Fc5u0ZjB0fzVxMfQF7miTqEhIcjyuqWh9XQ3jM8wMeNns
nlWcopmuWDF19RSp+Uhz1eDjNQvqNZa8kRi40HbFrc20gcpeqSHi0ScZSWJsU7bA
VuRtv31MdBfmAxhjESX8adnsVRjtJeTB+WYEO85E8nGjF7PrEDlTu7QwToBWJnQB
6+h/iX4rqC7+fR7VYH1GbD2mgHaKQ3r/TEaM/V+emv0PdHClZlqsu9Iz8NLpXYiR
`protect END_PROTECTED
