`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJNszrsg4RilmVJdgaRlhkhDIWm7Pp7vBnB8dg9w133AntBhQvwhd4Cy3p+4OWJf
EfBn4EvgiS+N3/EFuvLw5NylmURzvo/FnZPM+e/vWUteVZUle+ku6tlr+aCQCKUb
kPkBmzQe/xug7X9AXssHizNGy1Dxqqjh81b3EKzCDwyJSTclsQe3TRptF2erniRd
iCoFCQAH+TBbAnxDr++4955mNJAPiNUiMoQ12KtWBElzuiDFnIMeO8oph/VADATT
Ukpuj+Oz8dGzXXkh4c6n0UqCr82Fvm6cD1HY2HcGA+FwccUIM+5stXvfY4sFIDSf
xOYZ7G5p5LAtVUnerqcaHswlwfPYlbceUaofvJ4lrpYYaduYa771tFqPk2GmV5BG
UggWnxVepBW4sYj7x2uJhd0OcdwAbB/zkLAwH8LWstewJsj1AHh840zrOAslcwwT
qk7QlbXsh9Fb2JAHUh/uf3wjDQjvZ9eWw9bgysMLcnPQrYnwOyhuEv3BioUzToIx
n5YL/lQQBHoBy5uM1k4JteR7Yuhv64mManpmzJ+rdybIAEJSifL02UYWOJygA6KT
zZMKAD7jrZkhgriLLggOjEUM7AgaYFOIccXa/5EQReWsV1GvzQI8r+0ERucXyMvk
sqxzB3G1LCORi0DglPytFijHCajyaPS8aSeSdY0jRrVyEB9zjnARfJcOkPWSXG4l
cQFHFYxL6SZMpBl6jontF63dBfaAOUhjKXrifHL0vzUWUYbUdZoz3EnYoPdHLzy2
sVxuUfQ1Z3boiQ2gYvl0LhNfWIRWyZIyqe3xvT69sZ/wemdxZYzSWywDQ5IwvjXq
oaxJK1Lme9kfywDjhRc5Vm4/R2MlQnrxiuVoTZk0Tp+DMthFATOYZ7aQTJ460gdn
lYz+MtKRs+f8WDQpDfwtgVyCaC8MpM5fgURAnThLbKR2n1XhDP8P0kmL4S2AScVC
YjY356ReV+xvwTh3g2uITBO4VSsSL68MMMB5wdbgqzmwPyadGg/7jkk/hUg8NDp4
isSiQnIMBcOT5zDSQyDPTApm/BgDSjLVZ08/DX6h4s0aCTec/S5poKKwhQYvYuwp
8LdMsR5Kr0rL4gwADqW4sqE8XbeHZO/CLKgN4MvjANslLUgpVJfWUsxXFKwjX0DJ
ofyuB9RQhrJrx9xoJkkQrsiXnBK1mXSdKmW0kaS+MekiEbvHeFxm9YMLJ5cs/L4o
I9DlKJunCsAhXShWD/UiBwAdq4JzI5XpN5PLliuOTa7PFbnWUy3BJZI26a/rR4qd
0VZKcl4MxphBbK+9+1/Wgigwf+1d1J4dV1nL2UfmXfI=
`protect END_PROTECTED
