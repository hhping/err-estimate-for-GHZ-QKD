`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o24z+slJ/TAtdvcjH5g8n6g3Jh893wnMvglwgYvnD5EZ3uRRn6GygZxi9Egpbzm/
Z+Aajz3jlZNbP2+B/Yutz4Rz01Zdp/COrkBB/tgw+sOENycTzMFtYQVvri+v144i
2mEuXXZ+x+PBdLdWoQ+H7lH7vf4YC7coFzvPCqWHFl1+muzxBze/Yd37cJLSqYhL
KifPc9y5ydwqOQ9+vi9Fzmjky/SrXsVmb+WIRj5jtlcocklp3XlbPdFCfvqIjrxY
H+yA+Cksr9Lh5FjjWCIGfICtJ+cjmozJ9HHbIvKrO4oPJXdazEE/CdUzbjqOjiAN
qKs8hkMlBjjYNoh2S76HSG9LG+HcvT9uEe0LiUzH5WBcvlLG0C+5YcqblX5aKFcM
lRf2J/TNmkWmzea0d8wmQILSVXrR58ZNZKNNSPITns9AIg+Mg6JwXFzmgWRrMRLH
a0F3UdyXq3GE3ywVpiLKbMpWt9D6pi9GmqaLs6VnHVD8tEC3fz+3CqSdNz4pY9MO
ItbD+J1IpSJvt9Ypi3Q2nuaasv2EYXOb6DkmC+WWk5lLK1Mq4eiqOttdxVaLooFV
mYC03/n0KwQbIimJP3QjJlPjLFR8bxyYdYOFHw2KKkzDMupU4Fv1ow8YN9eo3wr5
0jcNCQQsxxEzt1x0vEABHBtwZVHoIV3/b5uyBIE27d9EgZGdvQYINe0A4DsDdDq/
`protect END_PROTECTED
