`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDevUGxnuNr28fHac0laspSK0nFUXPMTGwwim7XOKCQJ/WpFQ94eOdiVWIS/7psv
xdMRPxrJYwtsGg+RmGL8tJzxIuBEkeodGy/mhxh0eMpHURBG61qK5pMhwt80Dkjz
szndWAsKIVQ+ceFTuJf+1UR/bfFtmMdtKawQPtFbvOqvSrMgjveCWAZnjI1Z2jn4
a/00AOacZ3gJvN2JZtvINU1XqbH0ItLrbzJCgSnSMvb2GiBd2hLgtOoKGXhY3jiY
QOUXWKq+OaHaRUatKnhreGGRxcLVnAAZHZCdh8xdun0aOI/YvZybYxaxjK35gU6a
r7bDRiHLgZFOV9EoCiXGRJ0FrM5eNtUeH1yEhb4a7lDvzHLzJllpR0LuZjRXKR9f
iQBx4I5c/I9uY2rJyc4gtLr5suyV+L0E1eRQA56nGDDez+hN+cnLDNXc34McYnQH
3R41BsaDXb2gF5dwOyOvBNYpdbMyr16Q/telKVaeiwLt4Ydw0Q4yuo5u4kieAdzs
QVngySaW9mjWEhxJ94TljMS9Pc76IQQ4w3aorTPjHFNtcH2iySUGODFv/AynxG2Q
sIslKuFziew4vTCzefNhBOw+z3yAiPdYR8ibC41m8BBKukZ0gP7gA8Cbf4d9qUwl
LPiBewaXWk3U7QSxPt9l0C1LKhTf4ngzpDYQwC9BZ5RFEr9LudkNxj+vXpdN8n5n
odj+i150bAqeAALl1TLrWAHeLUbrBlghsCwUuOOYgEKvEpin7SP7zxqMGaJldsk9
DCBKgcxEXPwGP2bPVqnOP1wIzTUZJXit1dVWjiCO9C1X3ANCht+VHho4pMq1O6Ua
cilVKv0habiSHr9NaeHw0F015fbO2YRJ42bet6LhVr8No34bhN4EkMP35HU7P8EE
m9urmLlBpUsapA1Ls+6wCP868/YWCVX08ZPO4F+5pQpOCGy0jet00kInbVHAGHgy
D5vMKdsOLGi8nBOWgjYADbApLaTgdAsOC1Ih19SlC2Vl/J54AlKT9QmMtjcEVgl8
5QMJGaERKJErQILQSSuHzajiO+JvybufNgLHv22DEsKtHuAYrv6Zi12wjTwrzdd7
YB09Ci2u6HQ3AV15bBDVq0wIuDrWt6+X6poyzwg0WYP6rWuiBqNpT8vi4/XEwBK/
fAEY2TE63+xa6QDjWBsxyP0+TN4zMfr61p3tG8li0yCiV8+p8ax4w/3CcLxfs6j/
GgtoOX/wjBGoJ66g+dEBS32UxZNx/1VSyIIllcFkIwRaipnHHb6CJ6Kz6Clpdxhf
HP7LbBKaGtHoDdncW4VlvzTBygYqdt69AqkLVOKtC1UWE1aB3GFOkCvDlxxQgvT5
I7+f8lrOMLa4enQxtl6LC2zGzrso7l7i9VIj2zK1zsbxi7DnSTt1v5FURax0wYhz
CQRrk5uK3bv1UrD56LYnXPhlPn4DmGYATU86akqfhmOWKTgKfrCz1Kpr2V4s/4Fd
cGuqQogHuR5w9v2RhNORrZw1e2CJZPbastOXT3ukwUfiGwHTQ8hbYeRWGVROncHJ
xy42liLNc/N4ILCt8M7nP6MCFzANaef0YFFQYw0VN/87XSlQvXf+J711rnVq3TZ1
oq70m2pwms9wLn16+Fs+xNs3rqBHrf/JQmwYY3nSMPQrw+8ARXCmBcO4/EaN7Xqn
G49TdmnhlHFURk360Nt1xViLPWC/IDCUijAs4pBj0s9N3JsXQolqt+ShtqiaO6Gu
Pfl1gRuge74d90PBWAwc2E52y4Rwt0Qi2Tw92bZ8F4CJSAW41Idv2P8qNE+P+aI8
+NYRNbZsUHk+dJIKEVdlqdhWwZUsFa/T9N784GRknnsBIOd0ymI5z/0xDe5017iM
/XW8emA+t2puVXOt0MBQNVB7XzsDweeR6cylSeW03WwWxxFbGnTB1X03MYi8o+RN
pYjD0UWAjaoABdHPTJIlnTouxHnxLJPJQk6VX0qAsNCocSTSlt2ARwiUzfd8d4WC
PyNoN0VMciUPh1dmMaT1MU/lFQdmisBY+rL/zu/j6+fLOXinvYHQHwQxpCISRPlE
KCMDM+rvd/9rSicskDVo4qpnrF7K0ovcoc1N7TlWndHTuLMVg17spcfQsoTgc3ry
DdIiGyGxv8iPX8tHhS51eIV4zEB92ZlufowZQ1ssklM7+5JvLWX8pllcE+Eqkjr1
bEcX7JLAj+td063Utm7500b2MNStEuMkhqhCiE+dP6F/26ThWB9d2jH/NVYjjwyA
xNufYY0kT7QNC5wBwM0KX7Sqn6f8aiqaNFAjiTVwWHa17OqDeCtCKLtO0z0JWmVK
l9ksqQiJLalYv8YDc+Imhc0i4b9Vhtl7LnMZjGNKn+fOuH50vw+fZ+FrrVeXlqSQ
tD4onSTusLSh3bbFe023toOA48hZQAZiAfNxFaq5bMWzVMnfhewXXEFGDNXcdrte
EBMnGdx0Jb8tjNqXyrMaPVWkA1K6U4q++C+8PYkr5LaJK08B19z75CmFLMo8+ZDo
mcbVQ11W8F8TjHMwbLsQwTiJD1NEuv0bEGQD/fyufLAM4dRvJjoTwaPmQ4yXI0gN
yOWnmjKXYr8EDa39Rh1eGKsftUkuYtRFVwD/gzRzdBl/Cdp+31nDvz0MZSz4t9tz
I/z3wzvRsBt81xlme6cp8lLfmF5btBtKoyNKMAAPfepvoZj37qDQSV5R0yu1ZpF3
4AWgZhl0PO7tjTcjpJDDj4xqwC0I5yhmTEefW0yNdzyVSjI46DQlFafMuUgTZH+0
Xor6KM9VI8NPdMaMEN9Iz0Zo8QkNvtcRk4fc2lXBGloZ6PR/GC1llOHuHdryDd1F
qPzeeUCatpLJK27q6gOELG8iOd3y7I5RXrGYs46QxYkRsu7ZBedwVYhvVMMWrmNs
416uT9qzv1LTElMlvkwa+WybhJKMKWHuYh9Q4ngGpxkL/unD6giOMRzAYKYIIGjr
mGpuL4BlokNNzCopy8b6N2JF+9toAnqboAsR+uxRvAciXLMeU4XHzVc+DH/T1LX0
1VVLeBPFtyyr6U6DakBsqP5wvPhsJhrvKkE50pZtgHc/LMt64Id0oYRd1ArK30wz
SOQE0TO3PnR5Hj8YSMXT/93ItlacILq6P4cVqSzqxiToz1/mnFJYULUQYgeES7YY
G0GCw45G52w5AhxWWWd26X9wcDFHWK1O1WDcgZBc2/69Qk+4LbNddpdaMVA+/3zS
BihyUL61+vZG2MLwreBFN0BS89teM7jWNJa1Zj5Ewaq/8DRrWnvOPcZoUCQOtves
K6zZCVm2ZtvVNHU7cp2EvoC9ErN7rBnUYjBgMOPodOvCbMVK9djTn7D7MEnNw2l+
SNQNWRMIrsKWUd3XZ02SD+F6DMFGQEh6Hubr75s1jJG0rJHfitIL/+aZLBB1LKzT
mw90zB5nJbh9gagts9q4DP5tNu40op4jVK7abim6Fs+kzGrsipN2BEcB/6vW+ItW
DpZ2EQFxa0ygE4flce4s6HvEs1UavO+WC+IFdTrhfWIGYuvW88HoytDvfxYFeYCW
1PdYfbfWEB65yZttapUqpdRD1zxiDGzt4q4RyI4GrfQmzhJZvToX9M3oWU+L+BYw
mdMIf2Neyfm3elH8NQ40FgGBrVEEsETrHXm0GuH/lSkCfxv2pLAlbqIKUCr25jR1
FwjNSCQ9IqsMwHCtgmpNP531n9P+xYHDwYeDamKrtVpus5qQYNUOu10v4mX7JC0Z
qh9PXi4MDK/VZk0qQaOFF1sAHApPvbqmXavdhOy3woTFGlizX5QREBZCOhO6+4yW
AApCBULn//+wuhRPHx03baeq6IqdsOUzWVp2f6Nj1w046sr34/C418Ms/YrDXIQN
EkmMeBsy3xtx/kZt4bIOi2vEblCB0HEwYvhmH45tdRV7ZZdh9gfnnSfi7/Ouk342
nJRtLqzr68HpKj8m8/i8YH18v1CDp8sz4WhI0xBk9ENAfK5VhTvcDqIN1yujxDNW
9OloXZZzbptZLK6HM0KkdO+dKTjKPmLBU3L//lspcPcL+Ku8/fAxN2Ztw9n60PyU
aRL7Ag7ahqSEyKXXBWNEpDf/0wNmfajjLhEl/nKgQDp/ypvuxbVMRAQIz6kRWdpc
O9pMGZX8MhUXFMcnd6Ty1aPVz7BYyUHnXcWcjIWMgQjUUF2bKGJDhwJvGXHFTH2A
KvdW2jjlwsRLqpvUaXk1DdlGNAVAr4ZCellNxh3oNcsp+bSI1cjYLWnUW3vB3XUv
5/sgbxOiarXn+TIKnGkdCsAFfl5qnRxiJaXmwccF3InjH7VAlKTbgi/KEzXXp9IK
AuTI28MCP2I9Wwd06eAIp5yBEivdnuHnxwBXz8hgRmQl/ZlEpLbMq5enpvkXsShz
NLMKWOhfmkAt2Jkt1rSXKWfHS/7wkNeddWjN+8ShdxCiABhb25npU/ge7g3Yejj9
MFtFHpJuQfRig6f6525+q7OWK3x8u/S5uoTmpu2jfWo=
`protect END_PROTECTED
