`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ArDn241ohERbUhMYzGbAPlG/I5ZVzi+Qg7uW2MxZiHeBNs8pp94Wfs/gY6eiZxXf
SU9tjnjp9qMV6NaE8NJCgZqYqxCdrMN0dvkwf0VTC/QtMWjx8r7pNz7JfZ39c72A
Rtn1wGUP2PNNebJcm+BlYlaCDOpLnYdkMWzdOexfyrfdWymDvoEXt2HDl+opnDSQ
QtIpIRDFJCZv5cT4X/1oTDrrlpE6Ykl2KA7yE3vpb7rqEUMagToV7NgKGgRrTNd5
pxhjVN/op/hwz4tonjN46m63l4yZ+Q9WeJgjVCFZv7aoHxMNGBf35Ek9T0ZpjXK1
/lCfualrynTk7uv33hsKP11VjKhGbKOdtViWuojHaeoRu69TIvNklPGhyl9flcbY
kiD7n/UOCM9t13/EX9Me6jRqKp7BYXEm5J6Ab7zd044k7iQ5OVTHAJ26lsS0Fn7p
vo8pIJgTAOAm2MyRF6MEubkhzM04S69PCc6wyaF+5zE7RB0l63jsKD3rXLLJyh2h
GuTIT8lRPbgu5IrFG+OQ6S4Djykf4zXyuOWwJt25X5K67AH4upMSPbvKANuIhYrJ
Jivx2HVVxdzAdm/D3DpyloVl3XVxTsMcWmETOgTBbSPcAWZzaVLw5NdKQiakumuw
XWgU33iN2ECuk0MJyOrYJEsWvlX3q9m1kghiBpM/LJwg9ylyceLbMk1vYK+AKQwK
818rYTRceXPVf+O0DTrAir25+ryYkRaDwGPeTqLxyMmglIKvnmv+WpYmXMxU1giz
2LajEyIcdUe+7+wtCgfKwEMh83FTsXerc+pPdgAmL/lf0YHgygvfyH5ffTyCyD86
mJ63MwzvTdGQ1z+nUmdAcuyKK8psrT+PKxB+XssYP8SRF782VctRJhSb+BJzv8qi
Bh/CKQIhEay4aIBt2/4rZ0ZuxOMivUqQ3LomTArcmYKd+ptCfkVZgZQbdPsrm6zr
yPduLwKr/yZTDnsmvygB6ZgrblKiBI9iQYTPhIdnTZiEX9utoF0ergWSsij0TZj3
6RjjMhd4isAusu9XV9XlDjrYCvI7PaOepGutOkGdEqlHp0gmFikJjaM+/ycgHccK
G+3nadYRNLwvuZ2Ijwhl7qd4VK9MPmnwkuBj+IkgH8OyhjHlBAumPvUrJkzIvfWm
jvfncE9zIqmz7m+A0TP7D4gUyccR89tya5Y+wO65bVrBlw8RSssUAf3rXQ5x0cJc
+rA5V9Vuo1la9CNZCXTVwt/s88juj2UmE7m1Eux11AITIZ1aT21Eh/gS1A9z1NOq
QEOm3sWj4wi0sHvS8dFg2RQ+V4QPwUX0R63+qQvcdHHWmArnoYgMB+HtLGof3Got
fUTwBYUSNFdjZuNILYpdVcF1LQDu26UzYIoJaTWj05Cfff25ZPJp5Z+5qATIAV1M
UaEHpDI97P5FQq0IKKhX29uP3+lZYc/jvtq59OWkuCu8msWuTuQDpIrpKEqow9+i
WvRuA67XhKONElSS+aoejdJhJq9XrHxC+bVOn0x282ju6fv9oY3GBac5cVgqNEBF
XapyjVKbYNbN2j/DQ+Cw/gn1D25tde678FzSAiOFpR8/wswtpD9fXAcdXz7kkG87
w8MJk5aLOe7UBnxKIQFd7GWVyvn7ysKcNcMMy8jgJ4eaVk+KDbb33nh3ZtxOYrFu
IsojiXO4ypvxGvh5OqyPCCnxZYRoNayx4E8S9X1sVfzD2TSA5ja6O7EQxjY2+kkJ
mgTJhlxnAqJ73CJkKZ1EIcewjCTPrAJPvoPQgmxJfpkc82jnlmQDd23874EZ3D5x
dN2EEyFkrfqxBiVELTts07C7IXq8p0NMOrBe/S1AJu9CbXx+PHl6TR/Zbk03FYGk
0vyYsI0d0ZUOd+ASFisqnCKp1OuuRhgN8ZclgsCn/Bc2PF/gIJvWaez8Hc/CFgNe
GihdJN0rn2aje8VKdm4LX/yYN/8NJ0uaV24PDR4hyHwjVmhYU9orwNYr7Nis5xas
9M2Fj7L9hd/q5t+Db5qe6z6btFuuvF9kpKumlIxdB654wg1FfXrHHF020mTI+D3a
0SmGks5DGZ0AkKf/tylh+bg0lyNcw/HsM79IQg7msC91FKhLendPacyU23NKzjmW
z5mWYI/t8/wBOf500VRzWLPNc6m2uLvYQwTWEw4KtEhSs8kyYpcg7siVXXIbd41K
D6H9tuGEzgagd1/yzfJEIjCXHcbV9u5givW10bJ7Sai280eGJrUMb5aaYf2k1OUU
dlHeQ8lLI3rZdjB2nKOwJMvz9ZLi3yckthq8tYfjHYLMTOxPknNGHL9Yp50ochcP
4regj3wkdawX0tIjW2HlikIRcgCM2Qu4jNzEijgRP26GSo9b2/txFQaqU4weiXLk
2H29097hHHv+s4SmER336uwKlL3LrWpwcCYUgS/+qC4to/+bvcKrmqs1jUEVcjAU
5iwiJppOa9o5T+NFd2OMS3/TR8HslsbTNWqPYGSpbilz0Z2MQu1Si3eOnyBc38WG
mhuolNwaPOaWiz+mnGV7AMg4sZ1pR4PSzEyeuZePVWPB1J1Ex1zlEy0uPNYW5YOs
1a5RUON7UDNLymaxA9TlfUpYIxArFhIfQrui4mAtsQuRlEE/yf7sfxoiNtbTqFPp
BR6NBPHF1+hYvMr62dGneCTuJqtoA5SBI2cSs8D6L9QYiLvLzhHxsaQMOjIcE4tE
UCtP9N8R/5IdoduqS6eHC/t62uTCLWabvMHsI6KoxyEiCOkOOhUUuiu8vPstdEfT
KxIVw8mwmjg4fCO5zcczHZSUgg4ZfkqcXpyaW/ABeZihJoVkkT0zW+76FujV9oD/
kpvATdiFubFdNcGiIXaRkqESR95MAjttsoUgv0WCskR33SHtzL3fZC4S71t7gumz
CR/sxpDPJDO1+JjSLytpT56JWBhnUyehRAaka87clopdD87OWCZOGvXd5fnBHho5
BK5mNbs7TKyzpePQntCLX8bQqaWAi9eSKpNY7lwzvtqmNnBlEu9eAHme2NmN9H2x
mrtgWdmn6gh9dhP1+ckNXRHxdCKlGN9fmlheBSlMq017ZkPgoEJqqXthCm8sCrui
n859dvp/51v/FJorlBddV4nIvZBSwLvtcYZl7I9Ir6CZwsyCJi03DoRG/Otw3eE/
GypJAOnIYTF2E4Ezazs63Ppw1fiI39t8ns4K2czBLGmLgwVJVbXA7+SBmI529wYY
R/A7++syvWMSWXBwQHegpSUt96RuhK9/IsZ/ecj9vFm7mUG7hRYfaI6j9oEIZfF4
Y+v0jVy2gIRvkcv8hVSryMVtmE2+dqfsXiYMA1JWLdWX9j9ABZNSP/cRTpxN1egQ
wZL94DXZuTpbtm/mWyVDsrSOFsnOt8VtE2yqApjNpfuiMB12GaE8RRpabnjj7Sxj
TV+hePo8Fc/44EU27tqJA6hTClG7k61INU2d22M3+9oSkakfm/ar8mgefpYG57fV
J6KOPMLiSIaoGRxdHJK5dWgZpnrXzCjdLpJA0dvk4JINP6Q6v+SVjykHDPpFQa10
43w74fAHCYAzug3+HI0UYTSb0ovpPn4xt1gdBahj8RsELXd9P5FM1HZUrfY962xH
er7x7wqR4tbU0ogTin0KldMcWUj8nAJSeEtCPFqCC753qlODZa58j8rqm1H5y4gu
hUarMkF1rpNn01QlJ8ObYziqjPnvDRWtHTYNv+3/AJylxIk0BvoCOEWHRQb2lVGR
W0LeHcIMitVH03JCJO/eW1wp2tNtDB9vzBMiyezeK67MNIl+d3TJIFzyWgsnN1kn
2oFgbqdHuazw0qo0BLUZCLdhUv5o2JZRjg+E6Xgb0GnSOBycAoDhajE+bh2HooAI
VzvFn/vUGFhHTQOn5QxK+Wf3lG0D2lggy1HOfkxikIgB/DSXKh0m4f5qZFsBejzO
U2Bms2Zji5CJDmA3Ebq2ZtfwPCP++VuHejmApvkF0LreGMSsUrT6uBNjVmYMYIEf
WShbS6G4yEkkPgdcSNQfnY/wK8aFhkk90XoFMo29uBoX9YDOzc7CsHOFEwcElz7b
uHgZxsYQ2aav0zBEava+TFjWyUUtuq6vKFwsvEkxOWF8yzPwZbFSZ30hSuMxDJDE
7DwiXYEue4/RaW/IFvda2AINR6dGqYQLAd+wUQ0H6dC9BfDaGFYqpSvJc2lzUm2v
gHsJHybzqLurgQfKHwVkRNy27HafHdC38ZbDZaxdB+RNszQlr2UPXA4W4jzg4d44
tR5bdD9TtOVaK21NqqAE5uumBhcfdHk69xVcAi9JGlIChibK29roWpNj0fp3Kb1q
kaB5GUeGRzwmT+DeDc0uxWbil6alvVI+4syH83reAPlYWZZ6f0PDKA1pcIUCkf0c
JrdL42DWI2Q4dcmUjL6TgkFeNNpDGaVfHR3Hpxa8B3q9xZSfNpkQxioC6PGAISC5
hNfDMg40AZrHzqLG4a0Go3YgUOmnDfcqmGYBHEESi0TFuNgXwaevHRE7deRcISop
HjucHeYfEZrdYMVEUYh+L0133s+CPsqD52IBKWinZjPtu35rQH/0W7L30b5LpmuF
ViAmS/L8JQawCtv8IQQDOVgIO50hpiP6hbf6GZIbcjWiWiFR8evSPYT4ckTHyUve
HmOnMylaJcSK6XlsXDX5UQgN9kvKpuIEZqn8FbwGELvd5B2Arl6UWjv3WR4Py5JW
spETD+t0BWwSofzJ5YW+T4bwk1XkulKsrngSX6BmAerVsCRN9TqEFFmvftMmI+Mg
WaHM9AkHoPLn6XQUInDq4rZguie7PKYcYzeauB5z1dRtV3ufZpqriZPRLfnCX3Ry
zukg7roNE7tFrg9zXvc2Hnk0Usq7YNBWAKseGJME6HCMj8LFZ8/EEOZgsphKwUe/
n6YtbQD/DosYRJ0CNnQ5vgYC1re++5C7WifT5gjtiPAI+WJbXkwyefhEJSjiHEQR
TKSmVGAgt3BSxs7oE7H1MEkdoN2EqrBkEYJe9vBjH4iuWiQK6sQ4pBDtaxanRjIp
UQMUX3ZkS4wfA5+h2SVTGlGYWrzR25XpKv8imvJJh3RYMvoqvVJD0oOf79lQLJnr
iDvSBe9RXdBBWoVfxLbDSP1VcWLnDrctYcB1SwGsrHqXTeh9Mznv+m+fglacztx/
+QgUA5B0OI5bWbo0PLI3LO36+6Q4lnDWrGzZkcczZiQI0pSCUs8u+wg2bkn0TW48
crSEc4dV66tfhTJ/MMEux7R47gP+FT6ZtD1aoOQTTEo/fZxPVMkuglsJ0OeOjD5Z
9Ke6cvjD7Hiqlv1pg3jxXfenq/cUYwwaJBwByjNvwyH+kVub3KUBDtqRhwyEt3Wt
mv5HJbKgC4I7vju7xbIY8aZtHCdSmqzFueGDqMQBb5QPv7etqf892NR8LTmlBB4W
mngYQycgYR9xsn0sdTUD8qHzZnD+V0jmMYyMQaJv97iwxURM8yD4RQsgWP2VK/3a
nSDa9+VpWxwJKnr5WvS3YQ45hb/NvJaPq43ATYPyaCdJS8Zo5XVAlW/zuojXh1qK
b31EnnO0AC7M1xpG1QkKpQ2+xQa3IN4q42HBFVSBlQxtkoreFGH24A2wE/TfphQX
zyuyQ3EdKlgxoOdniM8U4HiwnOH2KnJ+GGKUmklCAZewMSp8HHATUkqLuwos9kvW
eopj7Lp6PA4etMMUNKQoQHO3iupJjrQ481GngrdJARjBryeQxq/U0MrsYZwxT+4w
+9nbPVYgiN1OWMasf8VU8iwcrgeAnckUWnu2HpQRpTxk9mgdc1aRLfbshGHOhPtt
3k8Xy3SFgR+29DbhQS0eZLk2/zuYNI9efblNqUc0J+ABFDA1MOjpXApeiQvmTaQo
UJrugGP/oZl80RBdeTRzvj3c8qOrHmnPBjGokrsCfmFIMtp2MwAZgacachvr1x5x
OtTL4nmTYT471PC+hGT7JP/QEh3u11cXxfPVjFr1feh6edf+fowCe8QXy7NtlqZ1
MfC040Nmb9R9xLEvtdnGHxBBVApU6ohzCzwjYRLfWUPDuSLTUZZ72dUMLHnu3HGi
lZ4AHWVzUYgAuvxaJpLb+IaklKn2b3V2nNjNduwoW/+mp1FxWb/01J85ctoefcaL
XvHE4EuRLIgaRDP4DL/X7oNOc3Voxu7o30JOEGchyNNJzsdxtusKZ4PHvA2ltdqW
rtTaplMg1Kq747ipHJIaf11qeMDJKWbJc751VFVmphIN+3VmlCz271nUU3lavxOo
6Jce6EtyWBf/N6qysCuzulUJMh0T9Lrs7IbXJVu+j/yThrU3jDsPTx/12R/M4SGr
XzfyHtnPqTAgtAC6ZoSbIWV3jhGrLKHulJAdCQ2dJs0dzmocbrJscKYG+aBWuVE5
eHlGNOiNTnPdS83PYTsQuQmSJNmmLscuurgGD6jjjDDA0M6nNUS9KO9SIYMEW1+E
yS+IWgl5ynG6tP8ZqiaTqUcQV6wSjzap6R/lqn9Fo3JdHxdpdNXje89PP2Krdb+X
O0fvKPQwfPvpBBBt8EAYSNk1hySxFe8+A8zYRML6D3rZ2J+EoQGONvh0ZYPATkUF
zRax2PcJ2yGkLlKdg+xqsk8lLvPgMvZ8JmmEks52JiRO/609Ywsusl2QdHLWVcZw
4Ik/AawRKb/g9hm0Onq3Z7CzkX0tUKGUqkmcpmxCQZFOM9JcrScHSCr8Yb1avrfe
txd9UHbjKo7adE4QPH5KX9PsrffV7PrcDuagHpGaNKwPXftXYRFFHBPvDGjiJ+ne
BdQ2mnrPYLL2X8+S5ej5SykZtWIVzonm3xXCKRaFuFChRBRjxYenNLJqvElJ7jNq
LYhMj2dJvYktiT/fUUu8/ixyw9v+khd7EyxdNNVpKzgZ5P73GM1LCWNZr5Dc/rJi
xa4C1qhEG+mMQaaeUWrk0jRg+76bZgsNTYNwJdgHkBxwNWHk5vf7Vk0qo9aPigyK
e0+3yIbvbE/83koKYGQDgErCbszr722Ndi3WxzGHPtr5MUTXTaiNejsuejWm/eng
IDr2UllJvzcPn1hIQU9jN2tx8i1UoZFt1537y1CZSP0PWnBb6iZnq6RZ2+70oU9g
HdkOTW1sIGqoRSi7eB3CovoNhZrYVX3LMmkUXCSfo6bB7BteAbeVSDLIl3/LtI/E
+89IdpjIQApCXonEJycwlZZgYSew8kbhmw61Mh47dSqAPmmb1DX+v9vfeUXQXjVZ
y/VaB4+R8YHGc4ggl7+vebl5U3OLUnGLIPoFdBF79dqsOijt8KjmBAup0FLBNgD1
7YRy7HHw1d/v/osscIMJFUvUJsJZAaP91r1wD1I0xh7gC4/4TksVr3oIajsPFJpf
Zw3OYae6JK1dZMyY4Xo4UA==
`protect END_PROTECTED
