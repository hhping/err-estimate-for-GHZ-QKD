`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i56byi9f1eng143r5M6jNUW0YGwCPevNX9RXiLc6LnnEgSCm92OpOSFPyZAlZ1/w
CXqm/AzKzJV+Z/JJk1A5yh6cv1CUF7qIC4vJoJeMYwAM/xW9QQU/IJJu2BkdyfiJ
JNo4sbF1yhbE5lXIzCtWgLPS0UKU/JKuUzuIljR2htVPG78UpRTPYOOs7g5alFo1
hBwi32NvcoCDkDhK5WxDHOmlRu2ooZbYubsnwXhgNvFryKoD/BXh45cazz/Zk163
8L9sU0JLcNgOPVOWk9b36ibLc2GiVZN6QR/tdhef+55MdMLEn/m9htStiKGUvxa6
12hVnSNS/aLwIKncOo0MAsAybkPnP2Yl7HbMspYRavi1VRO47dxZhjIYQpw5ib4/
xmFMBWUNMHBk22Umm/YlFv7SGaKllqbQLFLluoy6lo3oWc142IyLPsXhQ6GyCodh
uFZHXG5m11SVOR9hCZCezGqPP/QQ7KJrDdKZ+20aLYWUkDUarcgcJn/8MjUF48XW
o4WeC5QNg7CQ10/0tW2gC4QzSU83R0QrbCsP4FCgjmt6flho7IBnbJyDAc/IZgzX
ZMEMg3h1h6Y2FopLfHpBWZjBWCJ5+VQalc5RH1fNjSWWFRTziqxz9dfihLdofFwi
o542qPboPpCCTRwz+dHixm8A/3zEDRxnyIJwFKH/jZMzxKCFWOxIF0nHhFddZWmg
yit2HH8BHg9rUQFMloXCv07nLswsly1nGw+Kv2VTQ4jZtw5PaVFlBNPsltI85zrY
mQDXqXOO8alDy1xZMEYqHpxC+7+RTvwAnCAkZrbiEWffaEzbygPLMg6UX7oOc/6c
C/EQBOJOVM6Dc2pevEwCUCDvkdmbk//mE2x6bBvYWdLLT+lQ2VtyK2MPwNINrNi8
f8HLyxnzAVgAWb+rvFvw9mWhLddhCXIQd5t8GewrX1Z6CvO4FSwbc/HytGCARxjH
3zzhMe1bUbB0cLRDocEqMi01TO03bS9YqivYskdFHJi0+Tfrt/Fr6G8anylsb3nS
oeSZaIlZF5RYhJQPbv8p0U+OYT/AyML/z+Cgxbib4eY=
`protect END_PROTECTED
