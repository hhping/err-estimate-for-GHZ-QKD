`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XXwcPU02XDLifm2tjddo9Jsz7v02Nf7cdcRB7SIMhse7utY/BqHXN/nvZuZE8H6E
bld6jUMiFzyjgUOBr3+94mprw8CWEoV8AiMidUBUMcnQFMlNj0id+P68n4X4kOGs
nOaC3PceG6U4FGIeOSxeb8Dtu3KWlyzm/Io3lecAOw8BOHTokuD2WBO3QGIVKrLK
VNBvoW8w6q6gZvUOIoO9XmrHbM33A3jOCM1CzvJza531eKuUBG4qzAZ7/CI9I33G
Rz6/kzPlSABb1qKEsI2FIWy3cSgDLns64LTVSj19RI+isojuhglwqIs1R2SPIJ37
j6aFHNDdp7sE+7sKXIFOFMDHL89VytcE6BfUTbWLEDlCfdUUirbncMDHOyHCZEFN
UQrjMEhFrglf9KC1Rk2udrQ7XW1U/7IR2Q0oXKpc2nieQKZvP46TDV6i+oW8027p
k6+q+wfSNEpmn2esHUsuAbb19AXKVRmOVBgIvnNlhacQb5MdjXVKWeeIybgH5C+Z
eJOJn7BDhxev/3fmx/Qa+kCMM98qvp6cXVlM8l3+/17IrwGUN/53QX9eys2sgP12
SO/N3do43eLj8GXJeidtpl8oG3n7bFbguKaVgO2JlEiTSkipT4sUn5Othqe8Utmb
RvERTRQHu5JT6t3FO51ohxdvoGkJ6J+ujEliQtOyBPzB0oI0lieKf4MaxNn7pGrV
zvsaWZ9Aua6QNqGHICGxGN/wyM3yQDP7T9nvUa3Ssc6za1PCOIRgk/PBzKl88VJS
kq33Oaiqf/r+tik84koSPaoa8yHY3XqKHysG+LOsRXtNmuaFIJS+iHRCZIMbGmt2
rZ4IRmj0/aTBTDsXt4bZmBoKoilTxryKbQu3ejcUCyIlN6H6bf1KkBNDD9Nk6EaJ
fqjqbks5ZMX8o2o7f1tyguB9nnXY7FGT6kh/qrs65+BZbuDyxd4W5OAmmol4D4UH
73Bc1aSqjIh6RZnztZx3U+plh1ptoDrTLLgNw6wC8i4zaqRX+y5qO1p81qXSQW0F
/Z3x5EPKZD61me0W2ElmnX2r8xjk6Zy2dlF/DFJ0ZQH0zFNfu+PFIh2hDLNyHUDY
jm599cfXC3B1RrMs9GXEZTUB4gpGTfKYTyJhE8knVGT7km76IHiqXf4zYDGkITa0
9lKzRVzp7R/hocdhFTD1loaKh1bgm07QSoQaGizzaoPmvw5kXykqCI1JTuOqQhvH
7QHS1dQw+v4qEgQjU/KA6hrrV08ofO1G8Xa4K/EaRscWqJFU7afr1wPHi6pcnV0z
CULuvb0O9fpdxvKA64PnqmLlhfRTC8yELb59KMB194f02YcSwXhy2OgjBZQDPYwk
fWMRUKWZYs8WgNV1xkTFQurW61zfFgV9vkodLyo5KxxFSFXoYWN0qVigOFWGYnei
OIjyJoRTZ1OJuQsVwZIegoh9V+ZCwqsXQhvTaI1cEDp7ctMZtbQ1IXxi5Q2Y9zZ7
T57dOoEuyOo7LPFOCjfN7eYHKfl7et1fr/DNL0RMgaIT5u6UMFVzTSy5MMlGXhHL
W7bk2ANu1pg3+YLxbZi5mMVz20oLZ8FoSalQn+ElRNFBEjHAQ8fvu3oAcieLeKe+
QCq8JTFVcBtt5+95WNHwr9qPkvmRv1+J8YDGp0cyQ+IybLwWJbajvGrT7ZZecbTf
pSkVoagi6jRXIZMnospBaM8PEey76AncDfQhzGm2pjV73j31y3f8MWkdnvoaYZTv
KFFkHYQNP/ukE8DpKw8UAYWxHcseoT938o1ASOswM60Q0AyLnIPuR5W2PHNhImJG
LuIo6hHgbC1M/tU357lzSHNsEtgiZOg9PR0S92FVbC9OD7BqnpTYlBmbydyoxzH4
97CD/maquRlOK8TDiv1rn8huc3BbuEMkOzDTdsdiB83D5Lg9SdMdvr3xxMA1/4fg
TtXCZsM6DnWUwMC8XR2zZt3v6ATA+SFfY0njKsP0oFKArsgsAkcWfjNXVt0CY51N
IRbp4MFgxqckfa8C/Son00FbrgbhI2TZ2EN3cF9ZwBllIi/SdrZlMUzMgNks4JkN
t+Oo8XS6JmDBUxZWyJQcaBecjxEmtGWKEU2dcV3lU0EuBxsac4dCLjfl4qxCcOSj
rQ2uHFGXMC/hIKYOEPNidfhpQ285D8vjLmRUW2OWnupOPJJS80NVQ7lMobLcNd2E
EUK/dt6kXNPas/eKHL6xI+5QbVIs851+ybLeTn1w7NDUe45Yxk0NE7uL4brcZ+td
ZXMNbe36mk35i7W6N8Wz5ORPB2s2JZWqStEZMRpX4T+/If5uLtwWPKOszvP7K5+M
EXZRHh36+c5KQgDVKKkYV2Fg0xcQKY20sbQWmqiPAle/IZFZH8AvFgx1kkhBcVKi
Pswc5jOroPMYJqWWjjZPwm8xEnw9xEN7NyWGeCloKHWA1IK4vXDsVKzZbAQ5s7W2
usj11iluYpEJGjHYuvf5ss/ISJFcqIwdmtEwuGtz5LvaGcZs2t3pk45j/UKpjeJh
AgQGHZayzQizPvtEGcDI5xrNTfuoMRwyKqaubEymOwV+NYkk7OirLj1FF1G/Db0w
QYzuW4aVmmsWTt2Q59tVIjHR1zCt90e8DGLQYUtJ0E6X+93GX8oqY6dpPvr5lcSM
7Q67xgAsu1LEp1vAwmO4XuBbVMvkVcK9LQI5/WKLEGpgQ/n9XWt3AoiMy9IR6sJs
iZKPM+dthWHmwllilogAUZKIXmZMujtIyJJODzZYc7kUOB+CF7NYuGO3Bzwxvvob
BkULfX6TwKqcuDfT2ZtmIaO1EIbYVqnq+bNbh+QHSDFW572wALHcQPFBys8sG5LM
xt5yEE2i5XBg4N7zyxXISmtAhXzK/7UoLQjo25F+a/U2//hduc1vYUDVLIiMd8uo
zC/rHikWhK2JMtjNtzqoqrB+fX9yL+Y7H6JaV0BCQtdndnTQ1jtq85pMv3rrqHHk
pEcqFSKGaT/TBa6OgTYDGPRP0aPx5LiIT89co8kTFr3PAn3LAiz+P4E50TvPpZtO
JqWgqr6gdEWLV0b+IrlrfGey+EUXnnzgi1eAL8p5mPyugSYstdB7O5Pi8OnxzSBJ
fL7fFhxfhMqjJAlR22ct9Iqm8Thde596XfjtOOTnMo8/aKgJ8swvuinJu9afKHAM
OcJLQs+xXyXknJ3WyCG36o3kH9pKWxttasRHO4WZkHCKdwdin7P5VlNjDe6b3kYp
v3lCNScvwXkGJv4413cJg3JaDied1Vlg7bMKbJ7PJsB7YtWeMJwu9m/TZnmyV30v
toU6/LkqNc00aFtLosRVgIFAHcqx5ynYNkYxOj9xe6eu07ybKUu08UXCvqDyuMv/
0bcCqBZjflhqsJstqNiw5Z0SzsiVwTtI1fF2eAPdbhVxnGb/MGe5acJhoWL8NNuN
rE9NCzvoo+lGy8lcpXh/TGBHMwcjFRJJyFiTW+4XrR0tno1q+lco89h0sk/mj5yJ
SyRsgiDsyjOnRs6tu62us4qrKbjGfdZ/zt8tkdoR6MTxwAXdVxvPa1oKVWasTI9c
7n0q0AKQlFfOvfTsz9NZdWPODkMB7CHtIwraKq0QJtjrffWwr3SQTU2S3fslyO40
Mf6gUkREUgQyQfwNG3vCvnKbUPoMjg3FaUyeFcvzTz/33/W2yobXnYRClBSjpfiz
sLmdeROQFjz4fngNnIf2RNWJqqh+HMJfmNF1mtKXbsq5aSm444PgcdvJY4mjgwv1
GAHmeC5bJKfxTBDhBSdJD1ICGsPQgeDh84IwAmu4wE11fShRaU2WtJ6Ceb4oMtTY
lqv0MD0z6ipdmiqnwWAhxCFuhpJ9WQed5jnsnasSrEk+Cor1PfEPC3UTD6QPyrB8
NjE+0fq7Y2MwIHK18G4DxMm7s6mJto+iu+0BZgLoBF/QqhfnIpqGlj6bvMGsHnJZ
j1Ehw3CQmYYpDm16nF1Rps6FF1SCFmaQ9+MFPbGgg5/XjZ/MCSb6pSt9N/sfIwGi
qqtRH3JChwwFQgS7iXaEZBqJwoYHyjNLwdeL6ulA6Q/rri25RW6/gVN/8gq6oM9j
ctKyP5hZYAc4sn85QvdJpknsmWqdOXLXAGxdd4inwVwXp8VLJ+9HpPhe4TS7Fbfn
jziiu1z5jJM1o81c7lKmrZ5CgR5b/tT9/8InETcBS/yVOgWjSR8IvSfnFPZ4a3T2
HWu/LK2pzvT7lSQs3p+nkKydKULDqrVjJ8iVsjzauyfXIoex4jijajhABvu3kyCK
b/rAfFSjM7yjGWbFPsk2YHFI+SCAn8WP6Ry/r7d2JkWH8scu3tQu41ySLFc1xGLQ
zkfZwrWeOHCuqjasEbGtoJdrkweF0qaHhai7WxrfDWVtoTDpq2hZ95tL/7r7qgEW
kL25kJ+VhZactYnnYYfLmaEcQxLvAjaR/5yFZXpSwrQP71hMWzQJOBgrBML7Vts+
ddGd1Q8WtnWlVB9XmhoDOb0trvMw3avRW+et/R96A32zoa3g1MiKkSKVCMfJMm3i
AzFVEe1DL6N+apHW+ZT/IeydvJ6D4h8ruDQXRl/t6QFdWM4DDJHeCZKURGLo6TGb
ey1lsiJMkmbFhMLT5DybXewsKGDqJEN28XIiePt7LE/LseG2HufL4cXiVXqi7OXo
lU3sY95Zq5P8uiUGEt6RLVEPzxZxs1Z82whXj8tH8tYe9lLd+6oz+oNsTqdk7ZPC
TNSN/rFBqXf+9NPxUZOP81eBd1Os9fqeRMPdzJBaeIKLX0LNcaPjdwj+D58BIM0o
4HcuAEJqqKY6OvR5CkF81y1eGrbgPU2NFBW/ugxtz2ZAynW8i0zpEs3q6hHiQGMT
fZHEA3mK4Q7eFyCq7urrtg==
`protect END_PROTECTED
