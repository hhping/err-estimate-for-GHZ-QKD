`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L8Yp90zHURkQWi1HSibueKKtwMTrzCAY5AmzsXA7RmxRxuxNWOYAhzuZD6oo24rc
U6xrPOn7D/GymRSNNQR9YjvxpwHkEHsZgvG5S9ZZ7blW8lC5Eu7sj7rdz9lo0WaM
x5PC29FSPPTWFCB7y2AadTMgPy5HvEN8lwhcu1QMaOPFsZ2IJp/WCzjFXyrYclJA
Js47h8UJLeUfRg2vJBrt/+1lEgpNVoqpz8U0iALQW+fCUR3xrux4eNDHyGsdz611
phH+FdzyvxjyM6OqNdHvRNavUcG0dykMN+UCL5drtQUlMXNfiggJmPFosmPJa+Za
d1OxZf2xW2SfMqN5jHDXDCCtEuuBK00zZEl8GTT2LBlGKCAIYXdm+W4R86L5jG3/
6+YNjI3CGrpVXsQ4LCqXxpEAvey/ISYF/jPzewLjYCgF7RJ80aMZv61lBp9b6YSP
kSz3b9cWaToYIdAo5vct2jN122xAq8eTRulVzSuZ378B3N1xW/dCqMRcXozp/nPd
JPjQM2M24+pO9HAyM0LB5V5JOhQ/eA8OnR5vUaN31uLy80/VNBMoq4btJnNNm0HO
hqMzxt11BQqOG9sXuiyUsnHQlTsYIyY51yRgsSYpS1TQEiS1ygv4jEgYglUlVKYh
MDiJLTFEejZEwli/AmsR7E5SymfiEuhHO4yEeMuaIxXr3rSAGOD+t3bVFyhb+qXZ
v7Vg6hGGCkXtQb/YFlWKVtyzGswtkf53h8DYxx+bXjKjYVjOJNEkkVhnOBQDSHX5
HWRtArcnYNKRzjr028vEnBDxNpMcBneVNdYZ7wWbSaC2caAu7p2vcGtHcyXXaM0o
+AeLts8VH2m2ACLBK0PC5CwygZfkezdNvyXcn51RVDQ=
`protect END_PROTECTED
