`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1BwX+qZ6oU7FnmCnDyy1upPxsgcwt4D//zQ5Lda4EFesz1xRrhrAzx4DLrT6YWW
t3Y7bQo98gzMBCK837CRzSP1MLDA+0Xe2CXa6IBFDCLF/xxMixHThDXGWAglArXS
BN3nuh198NYEyOZIqVugzI9jpH/vpkXDe0BIJ3C6jqLdds7VVstXMy4Trf8JViki
hoM0n3DtdApHmE5GZ5EbB65287t6jA6mWZbqOw5ffyNDf1XBEMUe0jBnyF2jEVkv
x2WNN83prmd5M4MUEz5FbEzjAtbGqu55uGkTbd2+MX+5fjepGfvL3MCdUx6+BMV4
8Upc/qaQNpveHbl9OamMGM6uhxxadmCt0yToxDyfl1N9d6Fwys465eaHWhLaH6oG
jdPdWtQwFSC1FRBIerqbnj/6bU9B+e8gM+g3FNSxxkxiNuTn3tp40snjThDiJAOx
LuhepXsJpbnQ4j3Nfhc//0jEVCJoVLMmQyEM1kp5/vMXNTFTiMTKtxm5ypnPiQef
64Oi0Px70eTvF6OP9Stx7bHollMDNilFId2nHVsPgB8zH5+mUJc/iTWIav00BN5I
tZShgUyaSi2NKiW1P4xASFUearVEHBH+Z20xNLvmntRivXm68R0IHX3X55RFsbO9
RsZoVTmueL4Ho6NhMok/ZgELsIFXBA748LPZ21GsfYF0bwZYVqYeDROkm3Dx1tea
eTuwvfPZbpgvapDtKJudnjN6+dZYWK6y+OT8TRTL9BWcA3a9XU0oBeUAD9NrAW+T
WN9tk+d0ao6f78cgsO7I6a5WGVuvJcANUsPnF10RaN7tltY0TrCNocFs+PMmeYTn
zS8MRdhhST3Lagy82sG202IMzsuoQoFpKdZuUG7dsWlhDfd4QK5Te0DuTNeMPyQz
LJdz9kuBTbobYvKrZrk8+WZOo0BmmvozsNmpY5UmbooV4nyxloX1NS3HBGN2UFW0
g2KLOuA1ftoDJifAoeaCN7LMMdhUto6xoxgPi5j6it2JZyKRado7z1SGBtvjs1S4
94RH1BhWjR9kOlJHPe11PtQiskpK53J3y/c0JVezvdo819ds2uA5f5UdDO91XTbb
94gohro2+FCFRm7LyVxFMNonbrVsiD54AgMy3uSJwZnzFm7m5EScb8GxvtEgYtUR
iyL31EAS0Cbjt+3ZfZdt73XObSNf1eGWMU882k5KC+XteqMQ6ZnwvyiTpOzPztLV
0Vf5s2unaL9Ce47eE0twOURXftWFtCajt/e4iuBDUdG/GP96woOHboYimdaxlBjT
6ZgbexKWGsKqlZpERfczBVnQ0xhc0TIGKXokgEzgXLF3cBUJBMsOAdmXU7CBNCFC
CynKBw3z2HcmXedDaEiBtrsX6UrE+xKp9I07162XCIJxbGshrCMxAVsImKF20O/p
L2kzFRPUf7nGAyxEbj5FYPxwHKCBVQLcZRw/ZaDcHK/QBrQ4CxZodohrn2oNQnME
KeXvLYkba/H0aXk0Kc9AaS9FgZ6O8hYViCe2jH9MqN+aTLpuvzVkWerdjx9YMIq3
aREyNK0ZQ6iS9gZJvzw92K86lpiVFDTQlV4Yevt96Q3I8TP/y/xAHSXznaE7GdRG
BMqHvDdwJ0aWX8Zerjhqw50moAbtRLSkPzd6EUtDvKTn6gpHM5wgBQ/m4hP2tZKx
2XPWGPeLiQbO5Z/n75UAx5kCE0xsmlZPYuqOiXB7hPx6WehQbtiqGJkzwYJluzPW
cF2LMO4rJBB0XCb1HUTCpCAkS5osFjLw649wjDcF43110QXk3hum97MSjyzjrSg+
`protect END_PROTECTED
