`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKZMa1D7OoxxdwvLKueUqejdgFTVGxtqPiG3GLyE/EcOOH83+QAYQgi0CKsBveoA
CXJG4kmaEvD5iM8sHbpKeVkM6M0Z3C2cNLJdQT2WBAJUJmrDKsL2GfSE1oNwPKLo
mt2pMb0Xn9Islgj01F8dwKtJesp0HU8d60wULXUWMnRDwopBo/NjCVJ6kcv5jJ1a
rv4GXuytmAK5TZi0QR2SjN5w4EAxr/UHYGcREnWpoegfHlU4cv5DmXm8Zdir1/6X
x3WLAoSIsqa9pjelCnw5jHEM4WGN0GXLxS+smxHqvfKb1QMMgSsXzJTMLBOyiqCO
E/D7ogDuNVxs6ir/t0ojSlWYSPJO73FIlmZcmnqzqJ05vT21nMXHytMl4IFEvlQF
K+twd7+qeN+owuB5C84T8l03lDo6qXBFoLrklQg04jNDPbkmpUcjuMDyd5ZS7L/n
GDEZ1fEKCM5Wns2wjfXTb57mJTG+6e7T1pgjHtKX49FqN5UPNfwfqi7hChA2/GAT
VSO/x3d/muFwZUfteiBxF0JI2yIBHGOwHFEq+uleEL5nlaEsMvV+a801O3kjfg5K
X44ewTNzINcrZtnFHdI+KxpEuKjGOUd6pvdiSHb0fjLl29mBvNEhv/hBdqfb4o9n
Gbm8nPjJmQJ/KW5Xtnb2fzA3G4rJzrX5jOq/6cAVa/qqSi0lcRvAp7zgXcqJyr3G
`protect END_PROTECTED
