`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9oMVttJR9a7TB7Ps14QYTZRky/9k3EqzX6S8tICTmqN4+8SR61SFLMXcFMMO3iZ
J6/+B65jKVqzzl2sE+YJ2JYjkoxZmOfMh0CUKEt6bBKMM9/ItgOQf/jzh5d+VLd6
/jMixmbSHoEfwXKNXS5N7JcgzYCBMQ31lRVO3lUHwE78LMmqPk4sdw3dH/m4tDN9
huQ/rw37kdPGSolgKXMDVD7fAbtYqQuZByzVJn3w1WRvrh6FqBvaVulbOHriFdj7
wYvgtwJ+KJbLIqPDTBhVB/Mu70tmR9sUZR3d6hjFu1TD3qXDDv45ERu30xZ+KwMS
nxExQeeABS7UBXe8trBg8PqdZyCXz7t3azvCMrw/lrUphfzUJBnCReeWbjK8EX43
eJeeTTyiCNXsD1Yg4gB/tbHO39lXbNDQDOmXiLTEV3pw3O99XvTXl1Q5DcAZ6mbc
c0JN+tCyHsvhJ+BgBzZIacnpgr9nSyip9nng3djBY7ofDOwmJLq0CKtBZiudgkL8
RK7B7qyEXl7p5c2i2XpW7WXBTinuoJZCDrL7/nszlTL6hA4IetOhNStq4GfFbnsG
GU1fQTkgVdhnjJfrpBL0AJx+OFks8neuRZ0t6Wu5wgzlAzg3arQegNQc8Jb7ipxH
WI6uPY+TdPIOaV0tRifMxrbmo6BlfU+PTVYPaALUOkPA17WtOHScB4QXjSEfq0+a
x5ubKiZmmqV9y/3uqtUtnld/vDQQIuRShx+p2tjJKyIIAsbZUKwpbf+X32VY4wXe
5ZCmNnZDwtB+g96Mjf8K5+kNtwC5qVnW63ioYZD3DrDJm/taN6UlV0iYuFTXrLZE
JkmEMCM7vqaWSsMbnKluPyxfEFR2nnW6jPDuYqkD9HasIajOqvjwRvBt+ulEuEUT
qPTp8NgO/GTzXZb21yxEP00Ni5kz+58jML9VUSViM0oUPf0Uc6JKcHnof1j8YxmC
O4StDllKeocRl4BOSHOpbDvt2n4faFJHDDBItCe1dmtyX3dV64LurvNoDT7mM/yZ
dck/6bqe1EBSdagXT6UzZsLff1y3lBEk/Zm/Ni9hKL6JPnT9v3qpcK9IdIQEagvt
GAKTMHKHAhGuqSzLU+yfT5H+3gdlQCZcMQ4/cvDuMV3AdzCygr2wJjzPJUw/7uyg
UiVw+cyDw6OvxNunAfY0MTAubksKNIXzHDkszFtlrws/NeTzYUTMqGX8S134fNlm
UEA9U0qvUnrprHEMOPs4THSxHZDTNLhHcsCZxx7dc0MNnHMqNaQV138LKP1ng5Th
z0kfRjNcogto9fkg5s+wKgBChbzJRWrPrZdq4MsWwspmao5fXLTGO2KKS/qwUj5n
E6/QH2qp02eU6X+yA97oaEsXfEAwgapiebcED7ZrOhG7oBgBdHzJeowoUdcpEVts
LtWFE559XJMuP63/jEMcehQRcI6Xgz6zeTVbzaDXp+W13/jb7xCtBPYXpzq91xTX
Um1JQDokA/IPnDA3VMv30wWpBZW7pk91dIF754Tj+d5c7pBKn+tnwZw+e+ZfT3b0
nqNny4pIYDd9zrjpjtZZ/Tcd+2hXfKYi/prVRDRFQo13kQMc9RfWZEX6UBNtxYql
6rGEVTfqtmNOmwWl19yitEATmqqhGK4RjnQyye6jcWxwI4y1RwLk4ePazt3zptvi
+LddipaTiuhWBaMxLsCoZEna9JOhjrCWmbdVrqc7uC0mB91jrpsxMsIxwiA+AbEO
pGlYOdoFvC8mLx4PABiacMhl4fAvTIUfYK/fBXFo44CFcoH41XlWmstkrabKEeEG
bZ3iqP+CYz+GofDaezaMdverjYDZTJd8c5fSdwFZ6Vf8kzmjagt4nCFAhbOIfGtG
79NMtP4NpFzH0GvD/wEAdi0vuuGn3NKIdzRb3tp6XTpRVfsYS4UyhSwx/84jgZtq
HH4zBqkTVVPugO/377KUG3a3pXAig+zBeGbJgdpLrT0=
`protect END_PROTECTED
