`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
alVh0ciT70PnKiYmW1sT2+4Dbq6IE9bdvaGeX8R8JA5Ms4gKzF/mn/n3FV753Cs/
EkVq+nfJcUqdLp3ITIcYOs4LkDEMtcnrlF0/KwMnx21A864uxEi/BzFGQi9K/zM9
e2ox1nu0IHN5xTmvdF14+dNaXvCkZLOAvxX1b/o8Khq2hUIajNZ1gdPKtSuK/mxY
FifnlsDI5QBAekfyou/IhGaoadGlwLhSh34TSCIbFwmnEozHFnfdvQ1zCqMZImbN
zn02eX5W4nSrvZujUujEiqVdqxnCFC2Pk/KhJ7fE5UzbkmBKxPP6K48KGCxQqNvJ
YndnhGc1pIm6uMe7owyYTWaLhvEjmoCTjaureMQ3YMaYcY5nRqZFIz9IcVp8cXD9
+7LCYkDHs4S0traY/C2xs6J+LMnEA3wP8w/znibygySt1NvFUj2loJWX4nRu62ie
GCmcCvF/6+GDrYtevx4LHAVnZvobNaqqJN1oQypn4vTqxwKR3N0+ctfkRpT5UAd1
QbwhgSy2SjuFU6MLDE74/62MtQVqUavdLT22OuL/EL8vM5QfWHwt9pVV/1Roak7Q
Y4krgGNUJ2cpgBG5wdLRX4rz89U2+nnGL+GtfIBTTRE=
`protect END_PROTECTED
