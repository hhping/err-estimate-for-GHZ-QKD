`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTiaGMc1fNNjtFbEMGku6so/LAkHvBfrdl0VxaWhQCg8VyEVrOQks3PCE1n3Gfws
lsRtZljziJcus4nt8+jOR4aZY9QOtT8Mf4SeqBBB6lFZEPbIWmwHAzhKQw//iaRI
R+Ri7vIuup1BfTfrA0GZW/KHLnnXuoaJm2sCL9zptL+8yz0cMMrSxSOh9UtaGkCd
kT6ACRWpdqEKeA7X5YUfXfZ73CfDDXXTRjSuQAL2miCrPT0YDzPU1LhiHpqRnh2e
JkE5BklWoKyf7Jo5M/lrn3ZwnURInREnbBfC0KkzJ5zSs+IKTqOkSiZeXph7kMsQ
QtSA4zS/oqWhIb8/vE6OPcuKwpmDWnLjwjtaa9o6WzfbAziV5f2O45CUuBqcKAlE
AAlJJ6Wv0yAYMBWY5Uvd0NyiZVoCLwMBYytfSrJ3twkTyi0peuBCDGDsaHUanRts
b5p0ShdOWk3rq2Lq0RGK2dYtZBjRqqyFzciU3Rx30s7YVN9IMSxaFWq2hoXxKYPQ
B0zzhbvxj9+a9V2npEdkSe9HuYdTftdlDlEs5MeHipGz+y5ne8SOGPEJfNgKuufo
`protect END_PROTECTED
