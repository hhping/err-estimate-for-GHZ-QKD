`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFIbNCf30mtBa2shnZiy++YXyxKceo/Lq7gWhlmf2ZdyDRZh22KuGwrhsw+BVvm4
U8dTpBwnp8Hzu5sGG05Lf/AWVoFcLF8S3RqFq2hsQsTvfW1cBxYQJxaDzwYwLf2z
s1ZHfbnw/HU3PZmxr8NqkA9JOk494MAGE6XasLSU58Wewk9bp0cpUvpTdX03qCrq
tGU5KTmh+YByJe6HjDznx7S/yqUCBBjIVBSVTazZPmVuTmjT9Uj6jSpXLNqOKrCz
ZbpovD3wt/e5i1AEAVeZcCYt8C/Mo+DJ6Q66w/EfuksaiMMnfDbSsxCD3E48lGGD
1mpIqirTohyJzkIvAncKjUYSyc+wdf0OIVsf7nqgs1BByWgoTSlI8wESM1ebIcIr
AqLbz+u40QB5499hSIi0eo128xeXY0CwIlzp7xRWHxvfIjSlPyMxVs00SdoNvJ0S
h6oUZcrG+neUReg1/mVl2uxYoU0vzxMpQS1JUrhhJZbEPFW8jD+RbMNSDgZlDmQg
/Xv7kEOGXJU+P9WGPMvJya7RRDZCitl5MO7DRfV41M6GpYl1ogpKNDjDx8ryQP0o
hkOF/hRQLJ+Pb6iQw4WYgMX91xggU2RXtsbC17s/ivpJRQ0SZWYh9pAeGtgYwssk
Cec5aBnvVwVU8bBJ+r9gIQfrH+flnx9U16Wh09Fs+K452NJfatbUClxTzzWek8Y9
QPTOj4cnsmOQKVeeEzVVgjgab63ZPTHXy4/k5X34C8dDLVmiXHUr8f6Bd2Mzz9ID
8exRap+j4+GqtAhRtuU2d3W2zeYduLOP5hej/WNFNi2ZLMpw13wWCDZwS25L7ih3
qPEqCzI6jdQVxcn5MSKrdC75Grz+NWuu4XB6xsqG1oGx4AysAM02ykzeRV19nLZF
jejayIHeRDrG6q4mwra+4ZztiTejcs2RUUOtFgJodGwGKoPKn6zfZ+117wOUndp3
eqinawbs5uWOyxixT0BmUnCN+ynNBAhkYRvvs9ApLmAGI2fI0Oz2uxowq1IBFdch
I6fx0XUE0UmsdhSov39IJAQB6ZMd9+OvlMJJC3bsuHg4ib+cV1vIKd35WLpwyFqZ
ptRV9MUA5uXXNrxx7Nyk/NmiMvf57WZB/1qQ41mULNy3rULr2VwFCCUwX4P86Ihs
JuB4+u+WHxAP9TJ22lA/vzzrrfSjwjaBHXJzdSdQ+hGFDf33sgh0Ngx+jgBFnNqV
F2d4gXuEKwSKhdYa5M3SCjuYbt+SVN7equ26CbpcEbunCZUfUpRmeLyJ6VfxKNn7
/JDRpTXjsZaWIMI6fgnFlSang6G2KVXufYw6j9LCGnrHvb/Jzpu89wKOrfTauhIk
Lmr3R1qLOU7yrrSXg6+9dff7e0MUryZxKvKD9XZX57wolgnzKDenhSRrjmRe2rEa
50WQg6yPElsUmDixkjl6mXwmK5AvVDwpgXu+1QTkvGI+MjxYAWCxjHX40XItiMst
q5Zt1WVEegBry6whNAXEf/La6ukTyUhj3HRn4sBpye6NETHnBgqB68rkp8ClCF4p
jyDfBTSUaPy76FMV/UmQramkkaaGjXtg2YbHjwLlAwSSTJQ+fsM2ftXwTzotBiwc
qyhxmr/8rqsoVd7JDOYJEt8J35jhRmHZYqPQgoWHNIEIldylXbkxYABxkbih6Jyd
lGKOxK/K6fOif8d/Equ2SG2CNjCwsoaOHUxzXwtG01D1Lp2+/OdBtTAUUrsrDgh9
s8Yk7yCKxjBhs1IOp7ok/MEtQkgfXQZnQI9OR6BBCRgf5zpGRK1oyvF21yqqFnBG
t2p3tpm6+2aiM0kq3ZdzWRVSPyOTQCgu15BvvdMeVFYdfr2MIw1TQmIQHaaq50vC
IqQIPo+b2BXdh57dRRoqOQ==
`protect END_PROTECTED
