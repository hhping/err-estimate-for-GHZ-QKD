`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CAmXaBgI1NEZOmBjNtIq/B3L6Hbm2OaEyrCexC0EuzFh8YPfkbsFkJkDyaiNUON8
HftsZSSVCbZvXYcXYa8RuPMSvntYdLNtoM8hEX83pFqvIu1CEcPnCU2zw9BUoDwy
LaJkGRGtkZ4hmL9fdG62TIYf8d5LPKapLeVnuZqVW5IwuGyo+/OLJ0v+y3kzt8Ik
7EPDBiaWQOAgK5zO1U9+AMGB1Eg1PtKxIr4zJ1iqglKAv2YEmpTvgvooLaZEzQYn
lrNJyTpaPC3EeClQC4Wcoh+fwTvBqA9PKkCnc/93nb1ON8W1J1q2lctlpeGPv1G9
Ttue0BQpQnJPmHtsEGJjKph5SYQvfwkqklgGehG+Kmq9iauNE92kz/xbg8FrXr03
rS+QwtU6MdAjQ4t9luP3a1Ow6g8MjsT1vf8KNvkG3zXx3hnx2Wd4Hg8lb7kXiOs1
WL2CxIPjVJkvc/4oSjDZ+eUHKFEBgWFtGSWTK36qiB2X+8EaLbor/VC2JAIFyY0p
Rb9KEILlpl5x3jRLInFbrxBIAL5LCK4NNigfHmFeuTN/P1X53W4cgMN9OZjiJS0g
eh8/v9KnMgHNNaWwZP+1E4cYSVxfy0UmRe0uDBIke/+F6n51lqERYXrYsrHwvWW4
Ju+XNqV4d5Jwv2h39+GU8dzueiZGXQVuReSbDkAglXQhk3K0FROkORFmt0y7sgm+
iQF1U7buQGg21UNsOUFeRZextJLcEPGkaNxf8hE6zyn+NmXEDXzUKek6qG/38r1Z
0+uP+0A6drZwUgykTJ7YBfPuEcbOrTgOYZzlURXOHzSeVS1+y093JSuAQNMpeRQU
Sb6jwLlbFW3wxt+kodE8Ut6liBrN5wMMOhxbmv/K3jdPJqBqH50nqkoPXjRSB/r5
t/aDJgYjZztOz+rjla+6RGxRxjnnn5BoxRqI5g2zsazEZdSzViYRpx3O+UWdA88u
yOP/kzPZWriqQxACklaV6eAOsZCZln3IGzqeZj/Zt7Y4qZH74qYxspceM+3KivvI
167J1uJg1IGaO0PeFjQ6QaUrUl2bOxVwzpM1sOu58FNp/cEXGwdbtLQgmJfdIqfP
s2Rh4BnXyzjWuH0Z4sY6o+vDMIwfKTVXHTQKRNPOQBOAfrKYvVdcKY5KyrX+7m4s
IumrHvZR7UBHuPO+cy3YVX5AM2lFt0XpdnMkj+wD1XmD9yg5YYqk5MS/N0p68KE0
JLR+sEu3oPRyFu30dFEfSm7C8XN6DBD9Aws9RxMXNEk=
`protect END_PROTECTED
