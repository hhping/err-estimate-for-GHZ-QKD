`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsGjv7xRKAaRLFNNpY80waiy6N3EryBP0tdKJpSsfWgMm+YbhZM2Y69nZbey+/6z
I7HO0Bwe0/styvMxy29R/uEcSJY6nQornnsZSAWuvVaisHBg0hUJuCfbnya2rJwb
3/XhqSsGT3ba8swHpHNwaRZXzj6i8t6eNNg0WM91/t9FLWUJ0aXUitUZIBZ0YjCS
KQb6FgbKMSLRp7CYfjhgUQgTxgmPnYKOpgbCmkMBd4Q8SM+2eGzgO4VgaztvKcQw
mILVbswTXSNpEIS2QMN7HWIKR+cLhg3XjRtmL7e60euEKmmJ5zSgBhZnqn+4eiWT
jmy1NPD9+Z8TmyGDrDWRtXf/XH5SYufDNvz/B42/XAA=
`protect END_PROTECTED
