`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WpDYO+kCH2mzyneFJ8gyGt29Wbm4HqsmO+yLfkPytjBKzhfosh5dZ2GrlGKySnul
fADcvm9qwDD8VjPbvpCYdl8sXdDW015mp60PnttXMq+vNTQzQGlDoSZGjqtI+EKV
AqJbH4ecfGKX5GkMU3jY0xBhxh/CG2GLt25AhQRRapaGYwysWtCcy7sZBMGppKRy
+d/yiEvTCRhcpwLpeAUEIZYZTQi/VAn+KF3qKB5dR9Sdu4FZFo5PR+T8sJFuI8af
rbxld3hLJYMJTedUsj6u4gBuuKUoyjRJDTHswmIjBQPYXwQjLWnx1V4AeFWgwlnK
16TjyCltNzjsRvmU7iEnLgip6XgrFadDXLnAGpVN8m679FJ/JQwOBN3k6dwkJjWX
E3JTx4K6fNnGimt4kWqy8FevKkUNlb4G1EYoUdCnfBcz25sl4Hunmke6Ok2N6W09
qvVO+5bzMpkI+VJpa0pfPcLYGVe0YkaOkk0ARKgzPw/zmOTAl6pq/JM8F5O/ZXVf
yiwN8rAwwVXYkA1qmtPX6nfd1LsNQ2jKiW9TE7/1cN+os2jT4kjdwhZV8bvJ4zKy
c//MQdJ1PofI80wLH1KgPcEyyYqGNQFzouhfCGUEGeJ74hT4Kc10Jb4PWr9KuSp2
itK8hwsRKDzylG+gY0GC2Asdn4gCOaJ54oiJiUqW9fpX3VShIBggbqLnz5DFJ22R
WEsHy1A60pQHwKr7PvWBv2ydadX4tKiNMsTSg4fyJvUZRgnkNcAnBmQoRkzITwL4
pxl84A3lBWkLu5RpOHXceaeF0IMsp9JD164IT9f/aozq7+pd00TaP0pQko3RFKYc
iv+CJ4PLYIMqVhdaHRiSxV6QqMZqAvk99S4t6UpeOIhOFa95Gq+AqgShu/9MUooO
oR/gvP1l/l7LEXs0HFWFgYmO+FR1OkYl4cogGwYWyRcHCnM1wMuYL5sSNFn2M6dj
bceILuoJt0KM8EzM9rsFveoY1DsH7AYGjsXQhw/vUei5hn9u1jq4J1p6C0sV8uVS
70bCY3VrfK0dVFGn8nurhbQQUHKusdmU/g+lgQvFtD/zVlzCKJCSlRGA4W2CPNXQ
2eKigS1L7sN2/oVa5qJlXIrHjRLe2N1LzEsQYRgKbYamdX3K3eshu7ltiutQnEFY
NWyv7qInhKAFW89FJR8w4RKclqQS2IxhlVWwnEtF8rPdA7UWDIaLH1fVy957FKio
96PnM/pZ4xzGSZbZNHZhoxAnZ23Z84X9hrNiZ+DPGH1AMcUgSirrZBj3FNj29283
CXe4e4Q8Gol+jjCdvD23cOzNk2g1ut/ngygOVmREThOr62xTBlI2124/7GtIpsMn
8E2D7g9iMRaz696VKPtdVzoU1z0E6O6VnGdt5F+437kbk1I26IdzI61Tb8NWamqZ
P0er+jGRdnDF5d6O34iTETep5IAY7z0vMilOtQ640qNg0xVvcxjhBkmOQUo0l7iE
CF4yZdMBJn3fIjOmI5XdHKLI/ZL3AzD0I7Te/RUrzqNXe7b9PU+wrEsBOOrB+8dI
drcpL/ATON7tT8kzeg5ojZ379lB4zjiGaWX02j/r6a9biWqaDPjoQk7fby9OIekT
oO9EMGp7e1KLA7dq+1ihKbxVlEIjVp7qGgf0LKV1yXBfVnmgiAqe2nhdbtIROOGN
UTlEwn7AEQYJBs0ZxAkDZiBU2wHMuj5Pp6EAs6DoYC7jLXHH8qEsxukwr13Eq9r9
ErTLHWa7TeUsaX/zmYCPEs9RcvPGbejed1M4BJbJa+BLN5BnV4rZ1wqS8K4k0TsF
fABjH4YFzs5spBNN00Qt81Cht5EjesF+EudU8XvTC65euY6lhBp8u9yiho+5W8Ez
jK1lrJ77L6eZ0K66Xkox8UXyQUJGSmLnjEbyTYKwsE1lkN4AQMFg8KsC/84UvM+J
XcgtyqyKfOdvYK9LtGWNvSJ0QHs3jJkz24C23koPhUU9BoFtxGzC8bhaTk0ZBEuQ
O+OsxgjLCAZc7SuoxIJCKqNExpiiDLjxPHRB2MoFKcEwzX88vcky3kwo7QJQFrl8
yfshZqx3GC+JSUievKkZxc08IrlX2Yu2I+ESx1B8QrQNjEI3a37BOjaR5SBadsym
6r2y6YyegZ0SdGNS90aIsGgUW2h4E4uvto8OlMqN9dpNiKN2arN0uikqKppLAG94
omiOkwKQuNc/RDDb7StkXwzym+UT5cLTsjU2/YpFaCSVGT0YUF7jEnl8i5NCPGBb
7gM8TjCcojmDVffqwgQ1ynd26gMtn4sKSbw0i2fZwJlcf2ahsZsgB93sq9VT0zSC
imVJQcQMlQf2DAXh+iJQl9jkcPhvzMbN3Uzb1KbeE5ZG8RbS8f6VuDO2ga9nVmKE
+PVdxRnsjM6MwpzoWxjxSDlNb4PcQaPXmmzCEg2fDwkCkTNBF9fP6CZPTK2Oe2PS
aKIaRwP38CnD1BvLhVVPn8PhzTe3oNuxp2kBqDNXZN6ZTl6y6HQJ7f3K5K8CjCK+
XlynPx391vVT2mEF7lBi2zLd1d7BMZwIfctaabNMNCDE30Csua72KRxX055WL+Q4
EOiYSJv513MfttMN1on9gSbyyFdkWd5blMvHbj1MPPwDJ43V2gC/IUGf7K6LYs60
dh+Bp5UKPO0N0FzM+Hv3lpzSWLgwKwxfVWNHHU2Yoq5zZstDOddFhlfEyrpzSat3
RFGreC2pZ/GwWyGzNsHyvXxuNcQjr2T4Ix4QTkqM2zJakhtMRNvYohdDR/6Vaw7W
+cR3z1xnHy8QMuumQlb+2VdhqT+kqlJMVtnuecUWhi5/Qo3K9cpUNklnpPOJWGgo
aTQBmSGIKv6nHYjrzVZiSeU4akZT8OtgBySV5PUxetBeTB/Q/0xFeXRgxurpoqw1
UMizSfQak+dylm8B6NOWTu5PLe+XlAJFrmifpuLf6hVFTDINOZ+4kvr/RrOIdRnE
BVZqrxVtY9FNyIW/eeBYs61q3Mq+f5TeXJ8JuN49jCuKI3A2A8ssAll15FzSMRa0
CYdNb1XHXlbFxs605SoPNjkqFl57JU3hUHBOCm5gSJDjsia1fVskXdDLWO6VxVJx
Daz+/G23lKAo3Y5f+HquAjJuMg0plMekHpRRKaGZPOWDwSCCMzCjAVRgBBgVcXJN
BcOT6hngpRLBQa0DixOWOqAFLpuJd2aewfNC9FLBfnHXZJPq9U4wHFhCP5lgbbFY
bYiN2VUVuI5zFvJPC61W3Dosn3fORIZlQfse/Eg21cem7lCb6Xb0Tf0rifXBooJh
96X9pcugtfby6cxdrSPC0pW4a8yHGh1C+fIFPF8OB3TBjGCGgrLrCMdtFagJh67h
9K6UQ9mqGW7asl2oKFy86U0SVQ2ZJtGux44Chps+MDK4MuR8Jl96E6KYyFZfB2S1
y6X+rFJdiS9E7rcamq4DGA==
`protect END_PROTECTED
