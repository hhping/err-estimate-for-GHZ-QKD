`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFrw+BXF5PfEI7UBRD+cNVDoedlCc+STTfUqqd6/o8oLSDETLPyLigqOVhOB8bgJ
NGJ/GyD4IhOoBdG7AefffR22y+d4JOixHivWgWEhhZXiqfKYYXQNKZUksPPIjeKf
1N0zpjzs6px31tm73BVHPBw/y+OGXrG4b6kWz1vZR4iEJFfUocN3ZGICXt5VbhJC
0WA9YfQhgw10K1UV39oFW9G1wu1kbmAVbggDq0GSjpyIZ/vRmmiSXpXQ4+rtjDNv
HwqVl9n0J66ExOULEShHH0VIXK/tSXCJp3JdvkRKnp0yFQAFWfAv2BPmaLGhem+0
zt+YbuYcJtUFc8DPjO+3JaP7EHIM+Cv6eiS5QSVIcxNpyLHo7SgSo0HxBdw/80op
ux06WqYiwRbBMYmPprZGIt6gSSuJ9eXnDWkcGjYpi8tofnycui5ol8aMdOxAHvmj
5CMRUd26DrKF+qNIz28RDyLwUuvcRigyZdWm6/vsgjO+yWT4m6K0wgkoKKyreJJ8
IYwJXtxSFMbwZyx8LuFTk3UXAmOiTVRfxttC6LeNRycVU9c+jWjyDcu4mzNUFwmA
qB6EoOx68RgUXKyp4NCiVRko+rrt8NivgBbOjEo14cY7mZU+DR1kXZyLCnExIBDB
B8bAPyCdLKrJVLEUsko0xftq+B23zGkccpIlj/COrkDililM3/o7NjzQBDDPg8Rq
pB6HrkMpPzqIqKv3Ym4V6BNIqkXg9x6I1tWafMDk4zy3uyrGqsj3ZKYSIIG6kaFY
uSfVqg/IJYkZJ/lkRihLkbCoSlOZUYoX28BD/bfHAUUBpg3Ffb8p2tMYl2XnDVMc
TFFh5ev8IfQXZEZLT/HP2jtfPMM1mJMvBg/sAC8r3QK8YI8VmUbCnsn4SEK7ZHkV
9ZUq8yzhEqDCsgpOqOjNTI9HLOx9L9f2TliRgg/aO4MCuC41EmvDm4QxZkUNiusJ
/tZmGEfaxgRYQySunOcPPRoKYZbHAYFBgeb2ocPd5dYwMdrceUpcReSnL2KXh/zh
6aBkoi0dWi7jfKA6lawBhLgA/qTaJXODmMT7Iq4U+LPXbRre7LstC1EcDMffKcaT
5kzQgn7kUVBEEVKx2XxmrjKj7ahyw+4rR2B9ZSTcPg3XZWB+zGPBDup1maotdXz8
XEkmjZ80CkPgiZo+mHR37TuGzuVAFFVchrStfI290fUQeUyTouPb/lkneu/5oa//
SUkePVDcrYJ7A8fe+Vk0pSBbQ/Kmf5p3LYaZDpzzD8YgYw7z5FPfsY2ZlRBTmc/X
NHWq96eNQNy3mx1+cJyofZ+HyuhwQiHFd+3uCH4inHS2mDjp8cJLwVEYz9tomN+Y
sPmRBOKRosUf258NCZkPntdNJwx/MhHRO9RvWsTdfRSArrCATBtKx/P0pLRiLjxv
3qSRuYIdjTYLPHEn/nS/Cg==
`protect END_PROTECTED
