`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXgyRoMSSxRmcdO1AcNyAFseTVF0RazgPOZkis60Q5pJc1uqQQD8zNrivI4Obtqn
qkkS/Rfw6lV4LCkx5KTJnNLqCHZYbLKTEt6RByymHVYPjkbY/MzztARwxqfQlnSJ
v17qXVa0m9wzarEpslgyHNWtXzxiCkuXR0nM0BnFu2mnycBP0x+BTdLzPBXcKKNH
IM0Li0PJbkppf4joh96bfkTCvit5B3rTYm8mMxSnARdO6dD3pe5jL7SfpsNwhFJ9
mXFpGbiI/Arax1e5+fuOmcrPHfJn3iPIvcKotYzjtCW6TIaTc2DlcKvWphTR+vVJ
29PpIq/jRKbmeaCxWnDQqMaRCewRkifRyCjH3qIEAIQQihvKknBrRe9GHE+c9um3
0XvdgVz2IqjgCU9YhuspNWNpdwuFvXak3MY28fub8KEMJ5gKWDKR5NCXghL+doJX
yjpYGTn54XWFdaIa+ZPgcBmTRgaPaL2ibR+/lXjSoLLcJiWdKj4EphrM/y3tIC3t
nr0tjldI6M1ub04taDwbYojqkXnSBar2kyW6BZNy/dWDXtn7f2/ZoNAggwsrO3e+
3W74WpUYzdQH7l0wdNlpb4HQvviBgFQ2L0I/V1MbqXQVqvl8lNDB18O39KUCHpmy
hDQCQwokIDmvpUm/woP/zZyc7rK9bUVpZJDAixUMzmn1Lyxa0bQyVn6Dco5j2oMq
2LT4ulGtiyLZ12bnAQSrynd1P2O50LbiTHidiP+0vIAziK9quvfw/y6fzpHulc43
kJ0Jq9pWSrfNUobU35gWBBpPhD8KmIyW7eGwvysayEXyL/Ii0hckLvigKrWAJzma
3BbO6G25snmfQ7Klh57MuamJ6feHet98o9d0DPq7R0bPYjv0FyoJki1axSWuXaZz
G6pNrO9bQSW0bLJ9nNDoJb2TWDCXp2b3WQ+DJ2Sxf3F2fiXL/zYxjfY1zEHmnv+n
rVpcjZlvUFSx02GNPTSuiNzZpGZ+gk0r8J5yiCJQOyLjoQteksHIc0jntGe8iFF4
lRcBZJEyQtKx6y1C2ttJfaKLdO8IiU97tDcsZpEqy5ESaU2HTmPe+0t6arhvouJt
yjX9+7wyd3mLfQsEH3Bh1Dn7uXXqRmnnjJuffdr0YN1aoEsqGrNgMzd7O26monoH
h/OU0+60jV9wHR7xA6oPJ6za6yvhwHGD4abSMrJEFG+ns6Kwt3NaU1JYLeN8Cia1
BvMB6LKcyQn1UnhvrcBiadsW9huYQlgWGKZ1F/R7JLJ1VYLHHd+jG+Z7MRQ5rtMh
d3OcIBgJ8RFYFXX4SJN1ZQIiIg4pQkN5RWeMKnYJ+Wkwhb7AyzTu/zVbue81yGit
On8fmvGhMQyXBCxO1J+w0wrt2uZa5P5qalKbNOo5FbySp/P6JtP8RLLMkqEnYwLe
RR1juRMVakcG9p98RnvN5jCMULy3WKvGqOLW2vgsJlE+bIKu1lXeH/Jo9GP47SEJ
MOgPLYsb6xWXPY312bmOrDgC1vSVPUmL8iLzi/sZPMmxKW3rPXlwnHNTdap7C9zD
u9GUl7kQAX1f7B/PM3XpxYcJRj4YWWlHkwF+/6tAmNUMoMbVt3uG5VsioIOGtlLT
nXcP5PBculSy0m8jLqyH4qzaSe8dZ7FuqlBcSjUJymBzCnpaW6Twb2gd80ub3HvA
yPPo8p/F3ptVfz/YrJmJGsKFqUsjHEmlAoV5e/XKO4lRnGVABqztz3WOvO8lfSOb
MI6I/lXBA/VLDv/mUQEELMwJQJocoR9m2u2bPejbHgvCzflDULam6N2sw++B8iSs
0FtSg5XOlOoPuDJQ+7VW5f+2Yp/W6pfrx3c7Fvy8uPcSD+3cVo6amMgjTyu1rb6b
9rlT8HM8ePQ7TgMXOXoxA8Lvki7QlmWsr7w4ehw8R4AjQXlg41O5OdYGCM/w17R4
N2ArWyKzSXRStbIxcTblZNy3tEyuRJMxK7AwCvVn8eYJTSME6r/+CSOgHB3MfeIa
avqUiDKwohJUV6vQqHn5Fg8WZ95fGc2MVO9xl7+fG74IWa075WjYMFLyejfSMUoY
V/cpMNluzKN5jZSp7x5D/PF+m0EYNDePG95THWa9FHZvni5fCnbW1u/ey5iq89TU
+p3MYm1N3n1OD7Q+hf9dqlu2rNW5xzgpg5OrBo3L8Z8alnX8o3KZieEzNV2BDTbn
7Pze7qs70zTCif1a5DkLPSKeTjJXSf+KJT2JzjiZyJdhbStHft0AS18YwDK5WNO8
6slkxona7KgYA0SQ4v0nWB0aw2gb7P5PQ9cRqZoGJ8XngtsYT1cVJ1JrA+rnNUmt
LCjHnG9KiXn9Df2b/tfhSOPkc6wbnKWAor/FRe3REBGCQvwSpVvjQDTnHkB/9WTq
L3YvLB92JfHDaXE2MbRmJIOkzskh8/f75FwGGMEh5ufy6KpAb9GF8jbPYR5t3iEn
HQ7D272Gdinh/W4ggWySvoq3n3/gmxar5klOv6Qoh5S1YMbk28BmmhO0vVghjL4S
SJxT5i8pvsHgefiw7Wrsq6WhJHbcqjIdE+Vfbzh2WdHPxdpMeeNpvgwJAr7DO3E1
dU5U3LPrWviXCgcYtTLaraUPKViCKmT/xjJj8vUg+zTsNChDuPeqGwfu8gPDXp7L
l+f+VBA8kRzdLp3Q999SjBfw0EvqaKMhH/b0zFwgifmFXyMo6gI53Oe99mzdC7jp
jSzLUZRjgW50Tvoixwq+z0jVinGhMMjBu0ZX3UW09eJJanfmH6ogA0ZrSSh9RKHc
dSytjJrY32CuR6cmcjq4TmguKtS6HWWG+595cvbGYJ8DVlzF5DMqQUdw2plzLIqC
SljkcBtqwG7LSsUdxWpB/MfCHz5hDDqDDqyisDkB+kISecsjjvzWBr6uzaeTzbwG
DS1NX6776eVK94tQtHrp+BUQ1OEAzrpTQm0Qe6ehqQGQ/UHT2Gl/0UZruBgjUY4w
m/ikJ1rrj1jh7oEH469EJiFyO6opyEbt73QQu4f5XH1FSbxBFlQatt1UFpTEUhqG
bkv/zNRx5AH0t11uPWazasuNQxIN8hUkpIeDYRwaA1VaeMXBMrlPJ/26/9o9K6kT
VRsSyI2BLweX46IsOkgNAhy278r0cd94gi76kl0sA394YbgMBMCjlXorM3kPEqq1
kA/LMnd/U1LLM/3+Lnd1Nf4y7QgdExQh/ysHrLZOHiWzNPD/NvguYLLx0Z9jx0HN
uZVge78H6+hYd8b6HVdzUHiC94SkBkpb9heFUuCAMtZ56GCnd/q1+rI1dr4rYxsm
XpTb1xYIVbZZzu5my99v+VPaCaZE4XZmTh9DUB9p60ew3KPmYASPhrpXS68BRF9J
yVL/Tdx2WIFP6/p0zIiXu/1beP1n1UiUguluwX7fblo0nINZQ6UbVMtxOdVBpjKc
rcy7oLY/R/2lvS5anquUTkLMJbJs4sRFSb8PeKjZFX6hgiL44z+jdNL3e9HdB5Ec
/XDDp3QugkPZD1gb9iW4fF1S6pXx8C+BWiKhOqYAWSbA/R/VtThyA5dwTPxEBZ88
T8bpt1hfGdbFTiwPGe5kg06sOV/clQh2ewS8aqCLYD9+MBEviKUK6DAkvSObxL2R
88RfJ6aqFLbg8FiDgbLxNSek8HJIZuhrM9TrIg7KXfWjmnI9g1iiicFDmH41fPKH
hz3uGpJ+1f5yZwfyXecPHr43uSTmYyt1U6TDYFowVj21X6PyOMRCGdjCIiL2ocHW
hv9N1qybSGXWj/LwV20NfloWkpjqa75OLFztyLAOhnzAUTBU5nDiNAETAUmBcK+o
dGepzVYNa8cqdDrkSJ9LGlLkto0Ec8uN0RZ0N+eY0zWbT5K8rf1l6CtFPxe+xwuf
WXh1D4+xkEVGYy7ZU5Xz1eYjJtUUQb5NUC1Xeehk33FKemeTRmWG8h7Dnv6UGtSm
1DiycBHFaflee/6NZydGCU3GDIIICQ1MsyvZkP4kPxfeL/lNrFK87t5gJSKCYxVi
gReo6ZqlxJryeOy888fZGxBbBh5kbtUaop8qm2NrpgQPygIBZZ9kVlik9hweP3QU
qEIM4fN5BGnug0cXIxr7Dn2YNiUYRzpCw5awGhb56vlGHqjQ8cCY6Nl84flVzJUx
1oeKOZnoowlrN0YxYeqNgCyQabdTQSMOaxBifwwJ4SZrZIjTFgHsBrXyVK2JlN1z
bLLfC0CdTd9xNr1TCC7vg1ZoMk0ngiLGyOhp5W9cK8qzZj09m49n/OrOl1Crq2RG
KAkoQEd0F3mGkL0W/zknAMnqXD7KBbDCpCES/QWGf+MFwxvTb0AAPE+90xkP/Kcs
723QgctsOBMwjKft4bdaQBgmr9tg+qsoXFrTtjULB1E5ei8nyr0/TqYfQZGioVx/
QUYZo/UAdHT6ONeoyOHYtb2EdIOzIQsUD8XShU+gTg6jqStkOBAGBz/aovszNtoC
mfpZ9y8HXtRIwmV4c9HpoYm3fr2Ppya+5HcgI+SeQfzpX6al89fQ4CX7sHtQMm5c
ipeLW1mja8ytU7iIM649Uu7XjuBcPlnMt6Bf0YMA0DbtyCwart8cvkWPN6+9lFop
O1wSlvDD09GRW8tob3g/Jb8Gpk6yYt5LkAR45X4ePxOoIVMJh+j217Iz6UblvwKv
I7O/u7R5tgO0El0T7d+ai1m8YTVcwk5eprDYxW3kIEopWL20sEhCpmfIkcjmZUCb
lTxDln35OmMskcraRj3AvrpMzVTGJb/m1x3hWhvnZjZw1mbHBzGOYUm2ZTQnkNZ2
LMidECPdWlmCIso8+PvtvUJpmcLR6hne5BCl/C02nkILlCC5PUJDyLUnFuN0ML/D
hZ5XoaxVVbT7uQIH5h8sHw5gAPA4aUG4pjokVsLnDQvXAQbkQVS4dl9A9fEWoRtV
uya6deYhd1N4lY34D8eByQaeAsO3NF9Xc76FpWBr/2jOSpGUuTMu5fHnP4IQfNQL
+uv3nvjIYeuKEfy/PNHefCN4V0Hl3reiey8ly9l0C9V0K//LPOspvecOwj14K9xu
ALibRD6qi34QqAzVWPJLzDZTYLUULFUr17RZaaU8RoAQ/Jzw6isY1HaUma/c1Yv+
/zSa3O8pJC6UTxpcGLIY40HeqAHYWMHamp/pwcJbWPPW25cUnfbP2TkbSZ1A2Zj8
328RVY7sJ0hqFmPGAcTWr4F5GXlOn0HS+zJI8DpFvg04SwQIJS6kE+0PmOEcZPXR
Ktcb61JPSvs9bZmy86LBPfW/Mw+5y0qr76P4DXp/gTbxYUS29lvl/U/r73UWcxC6
at+baNv86PEMGlxZ6+FZH7nqd+Xx1VOWIehKRurss5YQ5FZUzGZy2NZ1e945+iBu
z+3/2o12RF3x4kHx5ZjONdZ3oldjVQPH4bkTqMcmqRk4p/GRF4U9uj57Jt2XOhbi
0WVI2+rMHWmBqf34MKDjcRZKmp3/Bq6+4TdnsP81QIoiBOq5pGBpjf+wCwTa48pB
58yWlDZuRpkH9jmuLUPgtC3cDAM/0PFhaz+ebDYUbFkzTE8iF8b3xfhgkBj9pEhh
KMUQ4IybNQfSiokT+6lzuP8U8J9R4p/5WudInC7Vdvxo9MlAz6mXMqDWRwkxGe3l
1hGer9Mnihw8ymjSado1NNFJetxcW7wHh8zRk7nul2fVcJBwY03XLJy33xnWTCpP
vJxWWkWkAIhKd2PEYFO1Gw==
`protect END_PROTECTED
