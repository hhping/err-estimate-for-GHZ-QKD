`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wt+XgKtXmGs4I1JJkzKS2R0rdVIRvDPBgMSC04UAlsRSVGFh0PPhyguykWFwFHtw
wIbK+Kik61Rj8wo9Gt9c8fjxCQ3wS5/q3OevYS4i5hID1zEQ3defN+2wc61jyDYE
assPGkHm2rsQPV6iCK2hWmyrjdoHFhYvdIL2dMW48YHqx4Eal7uAJwLS+qQTwdt9
oWsP1jg31NCsSmfq21TP/sS0sFTBRADNLssK8j2vh4agMq4kxs4z2qu8lAFAwVrM
yZHJj84dNb8x+4tYjlXZvlChLNbBsKgCX4zM9Y3j13b0vfYY1Psm0r4kL/8Kn6wq
IAjhzrX9kv5RdGbUuu5SSMd5M1RC5arodCd6SJoM41wiTjyUsJOYcVSXCl+d2+pw
Zfy2kPgY07Q8Bl/7ROQLD/sp6bav2yAhdfo4xmV0Ah1WpN2jHbnYGo0aR0mae4V5
5wYJUs4OT/GS4LyMfQzEjWySYmG3MJAkLytZHGEUNpPc6Zko23vcqcbRFQrDKkWn
ayD2GyhPTq4X6a9zc1vXd/Ztn9dOQ/q1oQQFUf3sXuEO1w8ekpmLghbwWasr9qfo
JlgZUwNvlZIS2I2dOSPzEcIZO8uq2SgP1PLnndE24pB2QB6HuhdpnFlC4G185bn9
Die7b9ttNamPCc1juAYYjopEMGDm6AmEHf5eILEuestYt1tqJsLeSjU5JYFRd47s
2NRhwqyrueWW0lsa6IzxCods1rgtQvUL4NEZE6FqxsWzFWza0JJHSjGRkNz88lLO
H3mOwU4Wu+I+qbATGXn6tA8p5Qw9Eel9M2/nz/gSvgBHP52vlnWTCwPh4qKuec/T
tzEFHFRj9VdBwaGOHgsGpEAT7EVwm8G+Z67v2lxguYm7OkJdNVgkhDdKQSzLxtV2
a7P31LK+wevig8ohw0fz20tNrbyYHFIv9Tc0AKPMNtsQb+ZrIrhFRaXoT8ahD/rv
oX4kkHHQGVx2nVEOJ8bBmEZDQl6D+rqQq1gkYwywLPY+ZAIxRjTp35jRrf667FWa
OxqxU5yNEG5Lvc/pehWvdhAAaZuxyrex0fdMVR24XqJee0qebQo0qTew2RsCLDq1
j06jDlCYfe1/VEJLvKGkewXuxgEuWPMYa300xUFEGpM=
`protect END_PROTECTED
