`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ix38Knt9yvQSpK+U6sq8t0XWNIm04wy/qgEY6nwS7dkJWkI/s0A4txb1FyPwv2O
Qim/LvH7frhdVZa7K1+ZhD6IzG1SsX9ucXKkDEinC5ftpOkPqcIbmG4tsI6lUt1R
8TaoHZ9o8LMHasXm/tPO1tJAqCvVc2rKoHDGUjksy2Nnc3Pco8hhl0gfYxGuf+s0
C4p97HlLdIkGZKn7BXlx+QRncF0utnqjUhagiLgt/FSrcijLGKJHxmDbxosDHY94
QJz3Li8Fn54yT2uwLgGCR3pSPPrFk3c4yPHQeJ35usbDCJVMK2y8Uw7VDoSqFpJU
oHbMaDlB7Q0bWUnwbMKfF4GBrrzZXEsksPHwwOcu3V+RrsP6h7vw2Pn0pwr2uYDg
gPnD2hD9Pnn1k+bgwtn5XpVbZIU9dK8rqiYzZuRnj154Qiw7PvkvyMsBk5OAVC3m
SeOK2wPLr4P8NE0qr6YPuGsIkd8X5AoMvcpC1lCnvySd9eTNdk2N/+CC1QMPijnH
OLERWbmj5owNvK13DFWVnbuRNJ5H1NuEJCHIas6k9YgkIuaQblMDaz/IcCdjQYAd
oJfK4i+u4q/7q3aWpycua9JHpdDCEyfBO2etNmFwSvHcbHTQjs6ODUIXu1T9vO6G
JMtf56X2KjrC08J8HJTa9hEBMSj6J58mc9fAXcbgGwyih07/ObWRaNtHMaAewISN
+3i+wDCE5VN/l1MYLbFYvLgryGQtAT9o5rTQSmfbStMF+SrvKKMx6bq+S2nFxfAN
`protect END_PROTECTED
