`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+lNRsIzeZYqr8Gf4r0C4NPK6Yiy37NT41eRcIjUW2NET7NKHUpG8gWHnRG0ol8d
DVFvaAzCHBqARzp/9J/P4wcFOlJFaK1ANbZ5o6OcAHCgnfgmj+6HcAyL/2u9V6Dx
FuFvzB+OtnWzNQIB0JUmvUG7yan9wC+PXl29Hl5SyFI/pEyiAY4d5MJIFWUD5P74
lIihaZkFknW9ZOyPMd8Op/ZdV0h43rFsVi9YyaWKN3QVisQid7IjjgtBuTYvuQBv
ofLutqGLjtrQyu2ISZ9kK9/NkO61lmAXLpBZVGIGH3Zh92g2AaL9hEJcOp6BcOoH
tP0riW4LVV0lMxNNSzFfn8Fb7bqaOuAJzvEjlsL2OpQfL3tR4UjD+kd2eFQtY6v6
zLdnIwG9z2GdMw/yEjJAXtjMi4wXTDownik9wqunyR42NJidsUGFkqadiKIXVz9m
XurTAudEgDytYRMtufWTIhP9t3cctCXDvD3MpucvCNz+L+qNlyjlXF+WMNBr5bly
exb4QXPbVEJnnRgqGNkiXGEbQs8tKx+CMGQzxn3HF3su0M8m/sk++ZfOOuy/7Upd
SGco74ionR7WzBS6/1baF04XyF+yTLGu6aQ38E4ppYtS59fVeprkXCdD1tJoPX0D
4BTcR8B/ohWLSWQCr+fZcBTlv98ArKCNlhpXRyx9cyHFJz7vQrFGM0W4SCeWZXZ/
xPWdkSn7MsWtTUxYR1BOBZs6TZ7+T7IaXVUa+CVXPaizgUcoreqTPeGAoL0Z8OFj
SROiEY9mqHho70iH7WHTsW2dEI8K/xpwNQCjtOeiMPaEt2AKaIWPa5szZiTy8NqF
i2+6Yeqa0/55/zO7Dqw8z4gQXhbxhd06DAtwaC4utaI7wV/2vVML3P/UUQF2zibv
c4q6aMFnyTOY/qQsJ3K461iGXVS0wptRR13c3gJZ4rLnmnQKaR9DRxq4+pz2U9wl
XRuu/BHF3xTmZIB8mRzweBaGZ/pfPZ+blIsX4loi+qxmyK79r8hfOH5tasJTskSn
CPMfnOKvH/8mE7nlPg/WlCUd4rbTT4iG1kr94rrCjMEpPTcHFZqWH8qeS/KjmtDD
Vbxc5EZRyB3CmpPKmhgi65BSH8fSIK15dQBh0EX2Q2ExDcoRHPjR7ZfG5HMl9UgC
w7nXZ7w2n74DNtNTv9mJ6a+0eMwi5xdp6RO3PzQI7jvpn+ob8lb7O3nSmvWGaFvI
eUz6pKOfvOXWZjQNaXZUumq8sheRDpa/8dqLOuRUPKjdw34gOnINvYwlNj0Mf3KF
QpHUdGvHrtBB4pQ3G55zJcF04l5xNWpIefPdQZFt7Uw5mDcKoPjtHBkFclGGBq8s
UJdyGMzifP9eHoJrEaNbPFa04rpz41pHnJe4hPPiVZqUv5O25TGvMuJ7MWudTPkI
gf44cDqWQw2gQX+A3Sb55rhxyMtAtSuTquAp9E3/swpRsX2to+T7xloW7aq31zAe
JdVe6/530kYGnt2gzL1y0VI7LzNbQpzXLYj5xyTaC1x1ZtXrZFsm6FH9HB/4tsCo
Sr/dzAsJ4U8IITrTdAUN00E/LhojWTtThVc26ZbKeeh/MT43poz8DE7234Gwg5EM
w4NW5pIBlhWvuCnx0i/nWrJIeeA4Z06oWW3tf8JLnsJ7iLAuKJVzASud1BbFOEK0
qlSLLkrQbDjv7fL53BJsNfbQFol94ADT2JvhhaJXHxH7wEui6QOGTbXUOqzKLN9O
A3IhwONyvdaIyE2Vz6XVXoFpnzuBpZn4HykjlWjByRGONU4M9gLj3t2WvyQUFMY5
9O5LGuLHGUzUxXLkC0uTyf732Dx1P+9nIrsfJnnWCTbaoVwcz/Zj5PTi4GErOhvY
Mt3nX5XAhybauhmCCL+jFuKssn4FT/3+a80QnUJWt/zRvb1Dz1HT0zbEjmrVANGZ
HKe9JyiYjwQrTJS6+WwdzO62sywDZ+AXN0paCHUhx4oswn2d65zEs+k8wVVS2xC4
nVynQREOXmlCNFqo2AZyJ/XxsciDacirmnXXjlnHhNBycGiFMyLD0gC3VYQUxlsE
lN9FOZjCnU2xfiNKhcWqMJ2mh7vK/s+ECbL1NiEGs0Ut8ywXIQ+oSbYAmmm6/hSP
b28KBBUHgT2ea1WKcYqtlxignOKOv4SPlXJnDZwiDIg+nUsBIpBcwFkw9Oe5WVO7
m6PhMxR3SWN89Tl6x/cbDPJQ+84pRKnmC9P+P4PtREofcAr/NChfcazAQsdD7Z0m
fj9DGuRSi98PnIAXGNZXsw5mMFovwFsUreoU6TmovhTMv+nNSYKb+/jtaLWfdYTp
Zu0AT8UpNo1UpLiHmtX2LP0TgD+OaGmD4GwHwusl5tyBxviqxZvXe39xNH5GBBux
tbGdLb1m4Uv9SI5deQH7dHRcH+zk3vOPWqWDO+gci4CtJr9Ru9UAEwDwUUDOPwHA
FmzwCAx6NNTxAgcg7UsLu9cgMXH7I4gaCKPRHXiNhnDnPphdRzkeMhplIRMRM2bA
3yTg83HbAbBBP65nqZ6wpsNtRjM9YGNRWndOAOFCnJ59FHsD832BpL0vQ+RWT4Zx
VWOZmEReoGbYVvyuNH8b9jLB84u+wdP2Oni+KZ8qTWz4bTMv9h4i897IfZhNtdaP
Ma7+XfuYuw3/ZGqzyGSWNEMn34T89L3bu9gIJT4ZyGCElxyxqASdmmI/6cLG54s0
Z0PM5mAKCiyw8T7KgqjuyWwicvza4MresPNF5b58G/DXk7xYm1lPaFGZqYWiLWkV
kz+sqa8cYimX4QaOe7nL8FsBe+C1v85kzMd7HF+gwqo=
`protect END_PROTECTED
