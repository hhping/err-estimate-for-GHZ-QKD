`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+Eeet3wISi0x5tC+bs540+UkGRFXIfAxouUmXNG3Hz6qUnMoyWFOGdn0JFDJqdc
xlOZq1sgmi7kZRld+D+8ugrpOyk6OoX/EkTn9sLZDOq3pquaz9TUImLR3KhvLaZc
qbpg750H/yiOxbyfngnT7Ixol7bDmddF5LpAgeeFGuFGnb+pKiMLKUvpkOTCLuRn
u0gtXXOo0CJhDWVImq2PafQ7ruHOuPtBF/oZxBjpS8j7SX1XFsU7Wmbc6S06lBZx
qfEWTkz/oqB+v3Ig1342bIUBuZZCSkuDxoRbUcAHOHPzv5lTS6IOri8uV5cvc7E4
VykZtmZBfOkmdx2WL8lcGzJW56M1Azf+qqRROm98Kn/WXp6sllFZmxQQqRTTzEq0
9b4tsucwjwQsNMmW0dMcHwrPnjXrhnHJgClOhKh1Q1cH6G/6Q6Ilh7jLv/vWpGdo
0YyZy/JYLmlKPld+e0l1VNEgl0ARWLDeudfZz9VkfMqgd3JpA2m3S/QCMfTFTNmx
OFHxsP/wnJ86eHdB20Qri6qWGMWjj++gaReZ36ZjBPoY07zLAHUyl6291EeJ6mdF
D/dRXRYL6lnfNK12j5i0pHI5+TcamH7tk8ra63ATOiHUrb4bbUVwhPxNYCBXOEww
XqgvDRlrCrYoMkSNofbdZqxSKVBayDUJafCqCByXr1fP0BPV4ILyvYz1KOiI3KYB
bV6xE6ZiTohI79tjJEBYN20F0bm+0nKMrYg7Ql9vRDbEwtSnulR5irh+OQlVKXFF
`protect END_PROTECTED
