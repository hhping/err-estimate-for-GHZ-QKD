`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eb2OPw/RmBnKUjEnrJ1qPfxVzo+vAeO8ZoGNlltOjwNtvmAnfblgS1L4ms59HrUh
LH8LRsLfp352XWiP+9MAqlui7aJTJu9/kRfxKToCRMjTeWW/hQ4+yYnXyjU8p9jG
O+N9AsTqXeeVlqpn96d4gaZMQAEuE5hI3cr9jWKF7P90zsc1AZ1nAXESz21A7Iig
fCrtJEZdAsR6Ffnv1m4FiQy4GdiGf+I/5alZIVHt2cml+Hj4o3rmaiVmgNL/Nb7a
31R/Fci2Ti8m+Xoqf2UchvCIpSg2cbqJe+82IYFyha3SiovzDA2ya1fchmfvQD3d
t9eIZ+dJkxQYGARIh/mIu/OQO8LjS5LdLvgfvqEKIpMFdNosDkZ6pGl61Ov6M7Bd
Srtu9hp+b8mHcHHKd/FAUccjgj8JWv8YXgAPviCKQXaCzIeINOahz0P2Vv4Mn/t5
DYGlGv8RfR/cwtWT+LgFdg==
`protect END_PROTECTED
