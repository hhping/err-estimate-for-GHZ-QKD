`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ttzN8sBiCZHMP3BgLoh+oCyaXwwEL5jO4eJG++GJer7eptca7JD61zoHkTsJ8+7L
fpheQRFnqSp4Ywg2C6utBd9GgJS8ECoVhL1MAhrO77x/ZM4pPOut/dqzuJl2jkPi
PNgulTsp8Lv4B+xnmQeorXWG0N+KAHfsTu/xTd88UUhBmGhF6REFDgTk6PPERpZ9
MaLjRo604p3keW6IvFeUJgFBX7PDqYcROT08GNwN6/DocjuhkpE79Xq8mqXgGmg5
laU/WBR6VL7t+5b99gLYnSO+yiVLzaO2JfUUU8Qk/tLX3osJrOK0aP6ttPNYE0CM
7m8pUHDUBm50jADf98b2sTL2wXppBnJrwizG0nDIScg=
`protect END_PROTECTED
