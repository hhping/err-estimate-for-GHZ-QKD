`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gkMzcBgWOIvNzJW/e2/FdtDYsYNQgRTSxjxeiMg1wj18EKmV96ho0NYXPvshD8+B
Dhe/ihFAGkdBVspWGuF2PCPl129kiUYCrPyWzlO5BFd3+oIb18du02AG69RsIRMe
iQMLPpcJkuj2nx8I6jSCr86OHjErPmpr2l7Wcqetam0miDBra/4XEIZydFKmcS+w
PGFg8S9Or+EsJq+H4EtL2qSFgU6ajJSHnmxoGYdw+WocpdItX+mmaFjZuSOgI2Nt
aQ6Lk3whJuJhhV4EU9KCZiZfsXApn1LdKB2cowKvWreGFOdE7fop/4DLOjRg9nVp
5k/D7G01DgvbhiTR0rIC3fnBLXg8u5ZihlkHaWJiGLJq2RYlpkjVNKbuwlo3qMiw
2OUVf75PPsaACJhKWifarx/eRiXobTSOrzAuwgbqDIf5mF30jTYBjZoxW4BAK7xN
yJTbLQjH9dDLqJntaWfEt6Y2aKR2cCwmozuKMTUGnxeEAaJ3LHYOMNNTdBY/tGRj
/ESE+KrCaFmGJBt5JzE0vh4Ylo3hgaV8U9xNYtmKy2hr8iIkIuTUaGzySZO1J7ag
mf7Roy3HaLmCSC6NnOplUoV9s/6fewZIfI3AdEFU7w2H0YTV8zuSvolMfh+8IPYD
LUaDO3Mb0eKWQ/OyVGIVXl40dLWl0DJt4JUAyxAp95JcebcPdqn7mv7xlmP8Ftmw
rmD39OeuRXe3slpeHcAxAL0Q7ELREKDYiCNgqRSLQQNo1ZozuU3RW3jC84j+MUq/
2uWqHOlM7PiVyCQ2AzmTjSKTYXLoxDU0R6hyxFXLDjY=
`protect END_PROTECTED
