`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gnFJTm2mszWrwld9tsMZJcydMQoRjjyFtQ0mgcEhlbUWiF/FkDP6C8Qsdywoj+Ie
N/bHoRsK/4xAJq5kvCCdQtc1pNFTuhodxQ4sOFgUOAWQra0IAMZG5zG0YUsQAIn6
Ig75tmm51nQi7Qz3eBAcHKKYsrPSWqhbUKKpEi+0Oh/PNcipFzgcyJVHx0r7JK3a
pVahpsoxinUOdqL8FH+yebxYb7q0hETFfiI5RikywkgnVql3DebC620doIDtvmaf
TBlejmC+/Slkv5NTS8QP+Xrbc1vLXbwysQp79bEUS5NHmXUTdTm7MVlt6Qgrsy0n
QlqLHqUDYmWIBuOF0x4LnmKyIW2azAwvCw6iZGxAJuDOIEagc1e2WXWrMj+1hgnS
bwVu9Rw98m8alPvTmg7DIK8gHx0B65KjXjcnbyxmvCGhuRcVAh04BdemY3A6OFxz
7cfHUExCB+7akuUKULd5jioCItXjocIwF30HJxnxJfVkw7Eg15+4cER+Uhr3J6Ez
1kYCd9CDwk5FIlKAc4/LghZQHyQC70WhM1YnqCeS4c0dLQyj3k7BAWl8gIEncMJu
qW9var3Yn95sK+XtnsjVbhX+SEd1sccKW7RG8AI8+DWJfwJbL7Z61NwGk2yqmXfj
2ybnvzL0O2G6JiyGMUON/y986FQstHjf4+qoHXDNGLGykeFWmuLq38MD4gYIUW3E
WQgTJEGr9bi09wlzLLGavnQxV+b67K27Tvb2K8NKcaAKcj/mVY8k7UMvseV9thLG
BV/IiBzVrRp281lwuiNYxySDvwPgs1gp8ce+Y7C7Ny3YEgcn2anKgB2tZwzxHSt7
8xzGQGt+7lSwjWJK/XmiLZKN3BxS+XqlevCWzoQMla1P686T/UuOWxsak8pKl4lN
oGBSh/qzz3Fjdc1VQENMWGfnwJ1SjuD3xaIxgUO71OAfj7utCNzZU5XQDUVt7Plk
bUwXrI36tq2OTwmOC6Fdg2BQuyc6BKle/2VLxg4ohBXio0+/M4DXYmbaYsO+mMHY
xaT7gUpn4eNOr5gKH3g0PIJQTM4OA8EADYXx5wMe5I6jKIBHwBq1DtD0yAgyeFoU
gdqtjneehHDVllWF+t0cvHI5lv2lZw2KKb6kGa4/oAsvz8/I6Pd77SL0KVMocAFX
6lCPqiGH0Rc108fS3KXyqpd2qShFHfoIEQbxCcPoQIuQZDo6UJ4qIKWT46uN9zZC
V8mrAIHBn9cT6ds3f9jFXqF66cRiA0QdawZhEt5PenNzIwcgIjhXOXxQ0etGJwh0
q8KHyHdE6zXHF0uJZg0urYHg8g6BTdfdReutRqA2TYpI6o4oOc1x/XSnHDpvAgLj
ifE55jcodjZxk39OE9W4h3SWviF4xOs6+OJNYdyiw8A8cW21Mbob7g0Swn9Ly7Eg
nYEEOEPR8XH+OcwDMuf6n4empSl405xCILLfkXfAGwv1/pdoXgehV83lRthMq8Wa
OWyMpT1j7/YkjdGL6mPt6p8qL7vDUzDrV4xdSbB4BIk6pRvdeyD0gdIg+JsJZA+8
UTQCursBrS3nTlgoQ4KijDwZvgnMCxe77NbymkwcfVqx8OICbClYMsihwOCEkr5M
p9G1d6UPdSuBg9WowNrGBrcianrrYHLTuExI2o6kj/rVZWn4Mya18qt0vnvCGRNB
OQNdKA+5LWt5hJO+Du0c9v15qHrX8IufZJTacXTchHiz0jOgQtvRLjcKFzHhy1m+
rFgM2DT4KnmL6TCrO1k/DStezPrJsY3cv4lp3w73uwB79SOE++Bq8z8CnWFffxUY
CyOQCBA/80VGrTFip6416wB5u97JHkiRCTuU/+JXfuLdy1VRKgsk5WxW16UDM7it
8Rqb/tTtKq0oQu7Ble/pnT20msR0LFqF8HIn4W+Xl/GsR1POjCKeH+WVKTkRvNFv
pJ4n+WcNzvKSewnrahNVq4EOeQDxQ65NGAveGRPqiAY31EUt0facRR8BnZui3JMm
f1Xgt0aqWGqiSWjej6pwLl0XYMN0Pvy9bRAynVDCL49X/6nq/JEVuUj8WzEvMwt9
MS7Da64q0VVT+g7XMn5gnV2wzP5QYiq+BfQOp6w0/xQiE6xySfYPUdbkwOYN+ijE
SdLEWPJAXKEantVBOt3GBEcfUeOpMfcs1Eq/lediuZ3GOWsrNnNcZomUBry5028O
M235bF7e/LXps0gO+H78T85kByBiNgKpd1ISFep0s5IpUcE3bZm63VG8eUf95VRM
AVjm3kNsTx/DVahfjQ15uooi0fKRfnW/uYX13Nc/gripAreuEZlqvaSeI0hjFGNN
0vO7FElRAutiCAgjdSLjDtPMrDUfBdwDwmyfcQEaD+SakWQoNAwAoGwFIYvqYDVn
UQiaW/GiX++SB9HXOzVaSm4bo6Rk3GqxS0n30I6xncLio0qr5SdpiNjWvqXppzPe
hZ5/1UHuXjfgv3HXAHO4ZR+r/GH4k+3biLLgPnrJNo/fBYLrcuAS7+NBr7D2eSJd
TqclUhQ0DajhRo+iBTeHWNIFGBRfSzvTFK/0J1CDPEzndMYuuqcrvMlJQ0QzohmO
7xnkexIIE1of+vvQ3vzsv3e1ISIZArwnD7Me2dDa3FM+64cf5/b5LgBIhjYhFo+r
Dzeleqm4AL1zrkkmF3Tnpfmsz5X6+iREEU34fdTOu8kbweT2UFElhCq2mMR1C3y1
myEr5GCuFsZms60XDXZBvaPPeYebK9zC/JUGoGX3TcNKSDdArr62uE9KAJLns+2l
hRHNOwzGqLLq9ErCqvlBSvFIIrk4R+QUGLL1y9ZrtF04SA5nO53aEaLhuTOc2qwd
Em/FHybtyPYPzse2c4Bvvli3znHASvQl+7F3eNE1FD/30CT5WOrloWJbvwPTtB06
jujmzQ5ExMsOamVjsQRSmcDplTZeGzggX1Hp+6GDZhWpOjKZimNze2mblJEoeawb
fhrmsVakkYOB/PAXUSfqHs1YgKphF/44wTwzS6mwkhwGBQVW2Fkm8Dlb1tpL/5i8
feOctlvxbQPnOOGJQp6gyhKmi7eIVY4imuFwkEAzYmRl9YKZHC0UIoWXedAdiNq4
F9RUECNV3Ry0l6ygTVHmE+Ft/ClePdBeU2yA4AxLDHWuCqjlDL8MRURxQtbZi39g
/ae8pI8n6DFOzUL5KIVuzw6NJ5KgMrj2Eees2XbjruoWDj+tAhUkvL8T+Pv/45Kk
OLHtY/Oldx+/NyuTRiSZLmkiFOhhus3HhFf8X7ek0/byuB1D1/C5wbJ4oMBlBZxg
uRO4HsEiQkHZl5dNTPy+hbK/9LX7yKfU9HQJGmdmeoP42F3eyn+UQk4PatsrvT4t
jzl3M+SvD+ZRValiTh5A845Lm7SRHcOikQKXITZFKUDb8/aaHWK1AQCYOF4EvN2j
QwfMIkVyFgR4Tv6VgjgNezJ0G4mUum8D7yG+N6mFWeUYhLiZaykpZWIZgilQK/BM
Ig4yECYSaPx5uBapLQ6Ru3LT2zizfwMwivJfmiMd/xU4be8v+TJD4Yc/ix3RtO86
ftFSP/Cqosh27/rhqAHv7oX1Mur+7VG8ckgSvI8lh5SDl/Y3A15POkdcTGVU225s
udg0IxkzbPLYg5h7hCmWAehKJLeuRswoqVfaNDeMja3ssXq8NCKodEvrr7qcrV2S
ZQKsV8nVe5wrFKC6z3SbvKyAVVzOh6tybsBBdPZHTWqRlqLX5LVtATCwL4LpHCuh
T20VUjQLapo4N29Ckph5m/Lc4TXqZ2bF5SwiEDUeQjwNBQ4uZIoVF8poDBZLA8IK
Dm4FeamUu1GxmJAeA0f4xJhfWJ6+S+OsaNGV6N2h4RApMkqAQ3YEhxxb4H1Z4GfQ
Zu/zzKdQkvgvHPwi+rk6KiwrCU8xDxHCb7BZlCQXA+pzpoOk1j7ORYSjskVH3WHR
pEspn/hpL04hJXAAaW7vOs2/WPgCyPblpjWvGr7/B20WepL6OIDdIDcnQiL5BEK1
4tzfrpBhwIO0wMpKJ2R8XhHim0m1Sj4HPGRDgYuAl3hNIHRboiCTAA6WoQ1CfPQ+
TjAQryDORh1o2LncI82QtZBMYGsConI+PPqoFH5nge+ExzvuGjpoMzYQcBfbnbqP
OPyvTEtSihGEdp7lwu/CyTWkJy/etgxF/bx/LMILXCcLIJSYbhaejIfJAi7ZYfaK
9ZyG4q7fsKZJHeG7X40Dr/QweryzZ1a4vs9gwNl+TznwVvNQGvM7ufKB3gcLkePV
fOYX3CCWZUaWsyEkwlM9UrxqkxWnncbA6NupIkQsW3jcDhi/nQryD/lmMcVq26td
ALSlgZ+pAtJNV/bL5XERgpEWN47GaqR0cnZcwFhuqb2xxaZK/mptUMuuS9lWA72R
K0HHTfjHTuFIZqfh0TbQOzQwHk58v8y5HrFlLsYQKPmXsZ36X69Tk1GLbf+4Xkjz
58ulB8JBB/BSJ2C/oKj/NTcVnOneFoheyNl36Ot7mCYYPiX8bX1V7dzHaNwAKfMf
etNPrOoOX1piQXD8JmhDgOPe2LWuDTuLcCQuAnd5r4OKTcZK0jiwu9tMMe9PCGhn
BHlsTsnrDB/h2//csXae6626QHE35a/n4H7U9DDvVjqWQGf6oSLqa4BgRrAXAikt
FNlQbwXbn4T+cSHNnH/JYc3ScgfvwTZ3VsbJSK60eAoUk8R4LBtFHnN0F5d1gdd6
MdzcbrX0htn3Emf8ahW1Rd55G5P1Tyq63JHkf3kv1EiEGTwEFuVdU6BiPPnYGOAr
dFR+VSi+AVmU85/XW0tmmLVkfydwCaHF14c3Uyeyh/kAycqnDqZAxd69shyA6PTR
dneiG9sCJD4DxYp0JQS8n03vTEe5SRqntKX8ALmKp9Iy1n9jfoVq8ISyxVZVJTub
qDnUPXos7N0Vjh7M7DHGtL+qwBsndZXDOa95plc+9fSsdjDZWg14unfOKL6Zy/rv
LrckFHdHiD7fXRgwO3pPgXSBaWT09mtxGRye1eb9qcMnw9mmWkzF+dBhm2o2nT9s
CnUlhtXd2y6thO1+mgrvJ0FHddWc7XmBQzuug21IyAKV2qrP1Enzuw4+I5SRUQUS
7c+l7X0xmmOJ/Khb2JJ7AHJrNcwKNYCFvTUAPNQmNhF8hxj61SOlNmEV1Mlw23LU
sHMy/5x0eI511oOsOdyQMehYvAhl4d2nsbDtizQZTYQESvGFOaoAgFBbiTVLXfDO
E3UfaiJ0kZWzs1gmGNKb7OrYGuES9nyba3L03maIjFGm8CS4TT95fi0TgPvXVoa8
PkIjzDQ/nzb4S9ZKGwiTUiArlRsiqCAD7zeWC8mToghXyBkUoWWER0VwdWw8tA2g
+rUx8NJEBOo8Q2jiTZWcOOBVgRNbqBJDYpT/YK1eJI3UZN0X+Xq2UhzTttXzTFGB
vVx2XaF63mG5PZ1SgLha5f1yIjyavUuiaoDeHaT/ggeq2iKcurYto1RFZ7cONKrU
Q1Ro7OHJheRMVuMd+tgswHodF6XBlr+VCgbSFeJXDyVAbcTNbYgIlK35gh0vXTHQ
xOAUvi2ouJDopVswH/VfAQT6eCWGXo/HX0snGKiMUBJph9Qqzp+IW89M1Ko/C1bj
pZcuQkAsNpzwb4YTwCrkZ7/op/Ojdz2lyTWvYkAVeAypb+h9DUolngoiXjKdKt/a
HkavFGaIDMBK3dEkD1h+17BPtOp3aZXbVPpVSxIw9CMucs7EmG2/pLETPt9wvkox
2RIBHMLcRbzq/L9G7DVj0aqAlOiz/lqgn2jDg1M6BYS8JpNQhZpvyVGmLqfOh57C
+PkpZVQYK3Xf850rKDYlFlV66VV2xBx8l0EPUAijoWaaBUjRdRmZa6Wb+JluLTrl
kwKEwBaxkYL97LfRRVO6gg4GAV/FWgsJ3GfixK1BEOaJDHd9ovEKXXkZBR82Lxgk
tWW61m9yFPbT4EC+ls5nqvYwE5lNBLbbWVJ2bzqpwCmIvfTuoc41UWCC9ilteu4x
Tcrf6pm04CTiB8m4EINPxXP+65/lcob3IhgUpNbF3orz4+z2/vVIcRWvM5AORUJA
YII2IkhHBLcJ5t1ukMRpTE52XtHwrpg2N7ykatIjhEtuBJ9+g5vBt0AzQ+utg4+N
FGTP/8F389ILjaaG++AVDW2J272vprYATqRokFOoscOufFm/+KuHfR9KBfCA+yn6
z5eQovCajQ4P4n9a5GOADSKmDqMSDRQnYwrcUmX/aDQtx8GemKqxtXDRJ4BoDFnv
fJfHCAchFKocJI8gpPscuQOBYJiqXjSKkgrSl1CEZeloLrWs0oUxk30B3b8BBj7Q
FCoDoahPT2e0WICo9XWjqqOO9L5F9lidemusRz+TY4cfFxCfqiB8gugWrlr7FGQY
HNJ7h1K2cfq5DFFBYxvSNUJdLDjGlq2rXfEWa38mNH2q9hd7DSX6/KxZ6SY4zp4J
URj8CVmUZ9uQsLmZUArmmGvaHZts9cDa8aGifpPI6oGKy7bQTK9DIflbGyb8Ajkp
RhnDCLNUCBeaXOrrtnHwBLWMWpkOFWiBX4t1Yj+Hg0j5PmO3X9ecmNRMbEVwNMqP
brDRo5IUe9AG6r5sbzvAekvl/A6LF8F2cRGCu81mBm+jqpoRX85HkhzUjmPxV0Op
8/2eMgTjI/aJzywjqt3sSicfXuRWGDKot2cNn0q8sqMyICFhy1qF526YL0Ic/5vY
4REgtSte9D8THj1RW+7qEF70kDAyU7r4y7mt1DT5ceSl2P+i5AbaxxYHQSopTi8I
RIJfiskyIgpxNg5bOYbvrxehgmUYOxZHGEiPJHHSU3LdZOkFlAZL6cmXLYAZez0G
VuM1H8E0xuQCvVzclIwbp+1Gvxcj9XZ2cbwjZalknjqfyf3cS8u0lDkDxCKXqgTt
alM2aRt0bUkvvYGd+I35zW/AT1e8TfbQAwpg4U11H/oQvnKhc8nVhmFAptb1l1Z9
BOfPopuc+6J5+hHISH69jknPXdOds5KKW+i+qy7p4iBlSBTMdOO7kp2L/HCjT+zF
M99cFcRCUKOdfD3JG0fcGQwSgqM4zHD7gUQVGnO6Kq3CPZPxoKavL94exYIB60FM
NLue1Ypqw68zNGTK5S4WHh6eLXNkwngq4JB9QAASMC2ZthS68jL0Akt4nZT+gAMR
m+aiVb0Psl0chbuhMVB8hzcp5Nz9I/r1RH4edtWRQdiUqds3kIqjaGhNBw0IgR5Q
yOcry/zFYBiuS2qYP1taCok8kzsi/YI6aKY7kLmqgJaSPeEEmiQYbrJOAdj7wyOz
JUUugq/8C0HYNZ+dCFtRjXzgKarXAaAG2kNwdGAqmhuZSkNda8n/nXPyJs3hbY+i
0Dy5iXTycVP5LXrEvpjGZmK7+uL2WsRZqzg8sfmfS1JSyrEzEmkjbh6ot0GCBx2i
EGgeSeUMbIlW0YWOH7c71A==
`protect END_PROTECTED
