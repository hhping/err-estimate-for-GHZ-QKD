`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfYB3uH7gS32vTRzaMlYxofkBnx9xG2IJMACiFzLOKgvK/7+sMOKeTla8rSlGjTK
zYMBlckVwTjcG3xswI9DXYjzXh8H9/ObGOyF4laGnUs8ZibGBGC+7veEt+dL4kp9
qt4MiX1FHDWM0BNBLGTKFzPX2h5J7qOYJ1KTGKhxb9KzLGz1d3cQttDkN/3SDXcy
BYuBgWZswrxzPLXNvw/sLV4QCWFHeoF1FwZ/xhSGO8oaJhF36DFXDYBFWe3muLcU
FIyWGy/T3+CJ7gTihogrNMV87+QxhyA6eJLLX0CAqVqjyoRqpwFxenExkWmCZhFD
Eu07I/rILkB2LIvKNKmv6zaq4jlLq/m05+EsHDpnvToBn+wCz3CEF3PAip5JwqZF
CYJ9fEBj3ndB5Sh6pbmpPsv60ZebfMFdEkgzEFJyHZe1R/JLKeDY/2kqcYdJFouc
fJwmFncFaJT209OD34xkHypAdRNRjM91ebPqVpOVkAvQ6bPb5ALKZD5R99l/d6pi
oJ6SMgSxlBOpYsLhEzZkUDLYN15Ji3Vk9DZb0h6uk40X+0j0LNrwUngzbmFUE9h3
8Q7VznmxVQDBZk2Viv2rBj100uw73INoWAFmPaKqaEVIuq2CwQ1ZCjcYYKihV9UC
OVPGwOMa9Y34J+iT2vXhYC2XS5HtiR7T1zwX0Ipbef+fctEOCFo3nBC7ib+QwxSe
X6mU91vp/xys3VChTov3s422vu4q4BLTWpF0aWJeCVSh4c6+SKlpAscFQoC+vL5n
5aXee4Xtjzzg5rcDxO+x+BnwjGGcIC3LCU93LA0kZEKv+UP8cdJt8KBo/JQjWixU
4QfkTBFiazlK8kfcick+Yu1P6xQlL4HqL6rRdFiRfKL9yx32LBwdaUvzBKMYCYfj
DGzr4DzCzj1eQh1k6HKMmQKqG2YlLTBIVcRTeG+1zCIQQ9WWOpDWs5dK/fe7RYzG
tCQhMwyawqZgvUUvQw4E+yDkf6a4fYzktuB7eToW9s9BNutyT7MY1VZNjqGrx5+N
utjEVHgn1xX/Kp/ImbfqhLwQQwxCTK6Wmb4DwW5V0nzGN5x4L4MsgdXebMkZavJ5
KhdT902vqWXWmQAqghpxHdvq92Y8ykF5YCSPt8kAnQZcIQBC4aSHLwwhkih3xO1C
kW9LddCw6vBLPenhwOS5ZScx0XoLcDh5uEIsdNMK6rMTsidjZPcKNM0M3YuJ/4DS
7IcAsQBcz/eJbYZq5i/TltEZAqUTGDijRlx7bylkVzmrvIIKlPa+e9ptWCM3sJm8
JcQyMpcDczbq3F5m9gfy6SeqChpPiAOCrZT6Jf+ApB9kyUkHlTG4xGAGqMOeMoIB
sf/ze3VLLHOvxSiEymVfricTz2cLNmgP4IiDzsYynBnT9f55RsIQmYy7atLOHtUG
4+WKO/T+JBX5i52FGMrys5l5319FXcSLGDTeQwVrI8O59S0Zfc41oD8Zp9uqpMSd
beJ1XZURIiln1mNAP6ia5vU5wx9uab4DHf8ay8FGd93mncSAf11Y2wO3DQB3WDYd
ONEuR0ccE3FXFQ5bdo4q1wQX+LGZr0GTHJBxCm/8HwHnoGJxClAQjexQvOzggsiZ
JIcICOdjXwAwfktBusNGxeGXbmlq1NcIQ3YN9JHUvOcLGhM1LqOz2h8Z926WOZ/0
S9FU8AWV51a2RH+bhv4vlSYmAk86owUzju0v75LdFR5W76aepqSXEqR8tKAUvGrI
7Tg7c+Ocvnx5UQwBat/RfpfDRtYOd0jXiwrzjLi3mi5gjRSr4mT+GgzOwYfVabwT
+1utwtPONRg1ng+hywPVX/do270axQ/3cOh4CqPQDah+Vj4RNHBz7MGBhlpQCC8C
nrpvylRojNXV/Pfk9InEDtxVduwRYKt1F2Ng85rTXBOgUdoFHglZ1eTcjzoFw7bl
AFo1K3QhtqHLlZjuoHdAPvzETa1uc6FKM76bDDA64gVEQWsPUJ5e85LT+rFoDE9V
ng8iYh+yBjLN1InMO4kVjp4SJe2toqOoA5j6E+UaFmJyIfvoAge3EU7QSVskVgLL
IibRAGGXuDVea46o4hs4LuaQV1reIF9s50SrRyWGGVYaNTREuXzgTLdxGQGxhr1Q
3BvO67XYdAKp3y9Mk/3xH79YN7vDFWTXGP+g4ufHzZdETMgUZEeUrp0qgP9PDbtI
K7+TOreEfUcNRmmDyWK4qCh5ws5USrgguWa7omFSO945wHls12juGt6SyRwD9QCH
bQMpa1if9rxXbJaIuV5wMW/Jee9NtQQnT0oNnWyJ+OTm37k7Tl4zKXQs4bbsFfUY
y7y53PchYcRpvNNMIAlTZOBYeoxuBlyMNZWrt1zqCza2cCLnSQgr57SEIhxpSsmJ
PRURNr+ZrZ0tLEmkLKuAntpMc3xiWSFZtM0NAZqKQFblAyC3pqaUeoxdlR8m5dhw
ZRMkPWIPSfksjkCv1kHeNR5CPgXdE6RasP1o9DDdCIl7emlWs+J4TcNUfT+tH3Wr
CicZMF12tzo2l3VemPuugdh6VLcYsfyZWKwh8jDTw3Tk3L3KhMlEAZDL+EJ4VEre
SlcOVMwd/2DVFLeyqzUyQJV2ZGPCcn9bF0b9urkH8qw3vZPl+pQuapXolFWXCvl/
D0A6xk23qLsHfVZs6oSGxUtlvTXDipfiYIkl3vppNnsD708q8Wpyim+VklPq/oRG
`protect END_PROTECTED
