`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPW4lmzIeURy66NgFUkPTCqI9GtbDfNg1nVQqqV8aF+XJpDjl1vq77AQmDIZgZnv
hiBpKkGcOsgBerrHGo/0/HFBRHIoT6CVZPsvcsIy/SYLU2YdWFrELXanS4hvTUNS
Kna7givhyAggF7AtpgtI4xH0i1Z5KckGhnoY7HIayse1OquWHuvaVu5m94gpNzlQ
flYU6o5omKr8t2QsS42X0IZB4Gdan8VmgNeXWsfn9F26M8U54sdXCB43+2WRG0AT
TLy46Y9EZ/ceLp7qgLL+Evzhb3XEQOrr7ZOFJYikL79yt2samTUH87zxmsZLeRM9
+8tdxGnvr9/EfrfdpFAsm9odyfmW0JcJsVpQ8gshiawK0nvYemYL09UAZIg0rXCV
2HzdUK/5jmvIjrPUzBdQXZaKVaE2cykpMtGQROLTJulDAaeYgyvar60CAYPjZJsJ
fPYyD9yF4s1eQ54JTgvdps9tRj9xwTsBRkFz86weOfMIP1g/Q8ai9KWZkyyxUcbW
YDKBrZ6ehLBmTwKg9m5yWTqd2rwn8GPk5p+GTZQijzyYhM/zHRbtYPsFK9sWJEOI
8V7I9YkNi3Uy/W80NKTFitIibUa5Zmz+sMXjWISFF0WffADTpKZXrqvt0G4WTEah
twPZ5whGOmq9GDhkkt3eKOTm9IQx+ctJSQkA5yWo/pk4xUqOs52gvT1MuynAtYkQ
aEadPjyyqHtSv8wYzJGC2aPRDX8XDV9sxxkNAjrH4Xi8kgckz3t6LHTCsLOwutrd
2SJJXdz/FvBZGkbQKF474ueZ6QrDsV/NGWZCxPN8kS1KXxxrAJ28eKqFIbwLk0Pk
66KfXdP8+F2lmnzmZRv5ARA6fiMmbaPDWd2zNFe1ZL8E3VOsZyR5WHRdJPYrpM1R
69wfawXNZyMcX2QihyNglMUzTlkhzhAbZA4qoI2RTNOYQqRGGr7HzekzoNy7ssoU
mo4ijq0cy8XK4/uXwbk8W5xcjgbN1qMZZPlGCKBY55CSm4vdOzY7f8pW8/esP93S
Gdmp321m93UJgfX9BpU4MHlmM8OWcRplfvbM7ZTYo8YbtuaA19dYqdockVbZ5zei
LYPbaFX/Fu7b+q7GmOYPCoqI9umbJr7MYrQiY6kv/FvjGlBO8WKXDQasmIYG0j5t
8z7pgpFk+Kf1x30zc9aMHM8VgMsISUjKIXcF2RRN3NPcUh/GO+j3w4VTt8ojTBKW
ZW8DLPdbtsm8W2/C4ewcS/grWjQFEgcaf+B8PeHYBPfLrzACqwbfecO98T5FiPu3
+nc0wrlo1VkDdDGOJBBKnHFeQ8lSqAUJkvE8d9wOifFpC50AEPQtCSEcL/WSfl87
t7ErzDg6gVouvPQ02je6qCQrfy3wLk1XVcw7N9pVKRNBTsN72das6T1L5WJg+/LU
vXuqVtdje8y2ef7mSJhSiAuRD4VVs6cEmFdcVmhGg7UNfVKxwKYW9wdmeWBV1a9j
Tb4Our2GifLt+0Cyj4czhGmCs10zvp+cYMjWqi3I1aS2dFkNaCU+80chwRCF4tSj
mbcUfxB0SP+/A7XIBmGf+OYYHEAFr797QZhGz2/Zeu14m4LByNbS81hZberhSwG3
6jKWONeTxY5V629Ap0hoRMmWuU7xFHI2xZrudk5ojj2N6ZaIvNL6VDm0S63mrRSS
4YCYUBTln3Nx2rlFDRbC7WmefkynsbqaFreGi+rX3j+531aIkQTToMD931k4OhVh
+j0kQKdN0LpCkcLGIMp/Z2PJfGWTjPSUGs43SSGSveNSKHLoqU4S00rW9vjHco8w
ZsVxrZy5XdLwtDfDga1u42bAIhG0OWFYMq41hcKtJrFp54kzR7bDm+z1nY06qT4o
/jdTGdJsleUzXLmfdGWDzvlSQ8RaOB8irR+aRpF3ooMwcGCusV3jAp2wrrwCNm65
/oBgcc6xF24/tUSyUev3Nh2ooBdAAJJlk9JBeXunDf3SfTvPMadGFrHeBehbmg4h
Bew94URsp52u3aXLIV7sKctd5cCCATm2Hz2hKCUhj6SdRahpRRRuvITCoBcZf1Ke
TMc6QJQApCVoJfZUGYtOyXmn1X0ZQlHB4vpiTGqPd7c=
`protect END_PROTECTED
