`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0KPsfcOXr9WAkBjkaViHaTaztvBwFDiISyi54vBJevZcY9A3CT3MIl59SyHDCQJ
Byv6hU68JXd0tKIWCphlycuSrf1VDaTadzB20+0DJ4cnwnhG8A/Rw7dy7SeSho2g
pU7f6LJak1xwa7kBYbMil7q9zbn42oo2eG4cjGmHk8ui3mvqMsU6DFeZS+kewgMA
+C9YgJZ23pJhsUMxZGifqzaRMHPV1bD54TsAD8FXV8I+YteuzIvo7x2u/CV6I1B+
bmgmAjbuRlyNxALeIoKGAPy/xTDgMnsrwwHdzz6MgmJ26wBQeLeRYKKm3VLlCHXW
JMHerCgNDUllVFmu0G/vdTrlUD4mztHpGxgIpxFiLR8jszG8/zDKqzK7rLnoDs7C
boYYAF58AdpivuGC8J3ZCE215aNB27yS9q4TDLPXcD83creHWJm0+8RGYYm5fqr4
cWWdTPr+icz5nRc0zVsreQ==
`protect END_PROTECTED
