`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhVa17VCRXqgg4oM6tC9A93ncbpITrhG+Bap6fk4+u/sCmbv3BvloiHlZ5BsRt05
jiNydjaKPNxNezx7lU5QGqA8ZMAzOzasxGbnzhWJNIUtQcs0l44XR1lz1o/c1+7Q
I1O59n+xOq+1ATYkmhGcz7gcSb5SuufZ8hxoMIyTZekFFkvJjcS+ntT9lLe7gHUP
ME33XIoVA8MovJyFSn3nt0Eb6M1R1YXwaKgjXvRuRlZtLxxRTV7U8o1IyhBzLc0R
z1HfcTOl/Wb+oERiq60v3j8xFDLHcNXrXxaHhbyx2X3QiLBOr0Dma7h5WoMDdhQB
p+uD9r4AJWTj9OGR7OdIPOYehWp7Q8VqBfGyAoDvHKSF6Ku6UYfIq8yFLp4qTQd+
H0rIQxVUnLxhXETqkF1JkJuPRIAV59uS6/cao5mENl5DUzqHPwsMaAf2f0etVQls
1cLWbSLgUnTmxtkt2fbHpZPrBrQ7AvCV+U27lAAEyo3lXwRYYHbC54NiKOfyqmZm
xMEfwVYLsnJ6bEhsHZ5J1v0UMHYiiCxelKZ9a5mTJFtHde4URvTTnKpGB8l2SBgH
EatHaU+pxSakPVZv/KYDcjuS/QLdzNOQ/tJaG2Gmj6LhF3lRsQjLAt+2xzYpv9jX
i9p2uHzcUuf76H42DeqUvG5CubqrY+4OKLfuyzIk0jrC904h2lFHHmy3bkFHFUHM
TesDTf98A+9pVXMMTBMmFf/J8j0rf+F5tjDVc1yT4mccybfZ5M0WM2Ts9mahesRz
7qAs4KjklgDKUAjzHkKbj5dsKhFtk4Y532ZQm9z9KDzLacUFJVgN65LqDCxdy7dQ
LTKA5WKwChyToEHEXGm4bQkxdk544tPej39gtRClpkLskOwXTnRwN0iHkTZ38n0e
3HRfM1VX6dWOopKAE12w/pm1mnnaxf+J/ptIFzSqbqv04gnkIzaXXVM8808FZDc6
7pws/7OFiwZkBVUToVELejBKFIO8EPv0atHpXtrhYKU3fU+anlon+CdltILTYGG5
YV7ej7U2ZbrTpYARcTo2Ln6QYSL5oLfnd8aM5dIEmb82RrR9K7mlRMkCnkky/YFF
K0ccJhtPG4AX4XXN5HbYc56+eeWzDVD2PKUeC/5NyXC5jyBrqsqNmQKtWECNorwY
U9VY0pXotEJUS04DjJ02CiK+LvausmQKIRh93A0deSh1PoiBpj59/Vn7wi6ywGLb
p592WHTnCv748v+WXETzVg==
`protect END_PROTECTED
