`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRv910a6v+5qfRr/uijZ5EkR8LccJP6oxXcO9YV0XOO6xK238bXcxXSyKpcARjXN
mdrETyCRRKlJ2itLqggnxvDUTAjU1UbQHdUbIE92gTLh1a9rOhkgeOidpQguNK0l
TltV1XRrkUKjlvhENlHcR2juQw2Osxu4M8etyjOmbjLHnDd1PLWLxBEA4etm19aI
7Q/5yrmzxepa15ZoIEa1HufxyS6wvBBaOA0fGNLlipKAtdzem67zmOowW0DpVd8o
MSuw17nWHVVDx5EGMefIJNxfIzE6sPZNbPIIgDoIDWMc0nDnHiO1HiGMMOrvbcoo
n4r5zEJHBFnGJFshgFjDCJJf94QU4AbEeeYmnAt/z8nUa0cm9/RFnOj1STwIF7IM
J9197JuPTVW7nhUAkYN5nmiMUZsdM93KWmwnQLSysIqC2AJ9wIjKpORACuVk8Pfk
actgX22vzp+1+xBwRzZNwmTsDPrBBxN1UapwwnhL6LvuvasSXSL73XCzAho3KZ8C
F/bOYm+HvFOAJTtZRd7cI2lEHIJKAsZdF5GrcvE/Z9bLkvrcLaEcnfe75YiJ3m5F
30+8OYWfUbQ3AzEJrpAO+5A7+xOK55L0UkeR6kfgOLp0Pmv3vuVFZ2fzz7zc6sjX
nDZrZb2jtwOzjbs9beO31OWeW9M6MnUCGjYypUVJGLf33fhBypNC1kha7pX/+nMJ
UfJ5uHoDP8htm4IXcX0LdkwH+lQGYISqxmjilv6eTonhUDqxHOVRt8sLLzj5O4IH
6RCOVuq/cEuuaHKGcsW8Pgj2i2R4AEK3T822Vg0XazCDFjV7UCPC4rYJooe62I+r
2QXb7P3o5LEYAqEYdoINEdQJOhpjsT9sJLX1KJBFN+fU0bN3DU9BZmHNQRAedy7A
kGQYLbLXm5eNpZRBB/gEI3vSZ8Gp9qrcJSW/440R4P+GBbu8hGX23QmpwmXh5Fv2
htAQZO5wlt9GJhYv28Nuc2P/+dwBXztEXSkMyI4ANfC8fyq7GeJ4gTDM7a/Q2MnL
zTYE4lnnEAvnjckD0TxZEAhW4dpJUmJ5+PgVKZ1FtsceDEbDBV2DaGtUb4bA/3SX
P6VL4yisBxzKKfnSdWRvqlTM+fkfmEuf45z/xiqhIP0F8L5mNMYmIGRZO+ltoaq/
iVADNcY9dEotNrnaXlD9oUwH6B8D6SeYhRBolVPDPfxaz6iwPkcZazpjlq0rb3MH
frlnwQsVlSvdo///mOaV5lTT0TXEXdM7U0y307NWWGUyRnj0z2lwWAm/BN8pNcp7
M+xdmKydJu6LGz24wig304rS4hHuK6h4YBFvdEwAMIQzbBimM+T9waTp6bvZ4iWH
W1LC2CjlHiQDvOH3gufNep3fiz5Kc1WDywpEw8bfQFZCiESrKs9PHbXiWhxDqJZh
iys1Vxqs8SK95UwahhtvgfCWzCl9EcVIxrSRJ48q+ZLCXocv2HMz0lZm8pXVlC6r
4H+sDjz8CzkhHkcdLyvWb9GJ7PRD7z7dXra1sz0618oHZ9su7im5u+5AMrl36DSG
klvJbRZ7qpih8EfMKkxzI0Wdg+t2ht0+x7EcWD3ZZYEe+VRYz577HbbGW+DcZEL5
5jaDWlCCf1ySbHL0kCFeTGUCj/gkfbLuj015eiChIYm9vTvPCR8IUSHy/PEpzz7b
v+wef1MErUrneP16M7mI6t6pcRoS+6ivbRg9xK4tejH78MbQiKcjlTFNgMUt0d4Y
qBDD0gIWJrfjuQSGpLDnr0nthWyoL6YoPDnklVMPjUbZhZD3b5c2x4JwfP8BhTd/
3iwZmxJoxDDPZX+P8wiIAEEk5tk6IPWQhgd+9G4wwFtAR1D2D+/8npx3ikTUANJY
DSIa2wpW+CdDyU1Rr10zN05DFIdNkNLbsxuk2evz09i91bY0ktdlCNm7a7HR8okp
469s9DCiVbnvSW9lIklF/EO+gbNEEaAiPcNc0ZFDlOXUtIinLUIKPRXH2xaHeXZp
tYdVY3p7o0SEMhbVjmFSGOcBnh+QILoesp4tKInVQzQgBpWFGzKjPQLCIPqL/3Hj
MUHKVnPoUPgu2/F8gIMcDMjk5wKMU+eix2dVNQYsCqUYSh2NrZDe1KaBndb1/Ddn
iTAmyJ8D35mSVtCFTMQxHwV9PyL/XHy7ZCZZq4069bbzPs9fQGB8Z5nXkfIx2mNh
LY0fdmHpwzXphzvNE7EtZvVlIRReddI9x2LpLr6ai56SfajJ0pV1Hv655rYkFrky
/B0vCSRMn8xJJHLXdSD/pOP4eqJyPWSuXmvNDaPobFg3Exq6n65IrECb+iSCuuhv
O2QYYOLX0ZJrrTfKNbXJB167KKO8zbXEvxfLqewciagYGnBspFCSTUzANtsdy3uE
4lEvsJrnRuFuzkVBYFn27jDjCr2iR5aimMY1C4SndaxumFT0/ikDqDIwF56BG0bK
4T7k4KXi15WCH4g4jntOHEnGHdsH0vj+JUr8bTHKCRtCqGQW3Cqdk510ic9OUsdW
U4Ro/qdtN91cTanoV6W6yfpga9GiM3wY6YoPcdMwZX3AcERsA0koTiQyBc1Ph5ji
nnQA/j8uZ8GtEhF0NDbLuIlqh8G6AMIsloxRdijH4Ww3GW94/1ANbK8iD6a5cw4h
5fYdnYsFnKQis62jjkpLhB0RcwQA1WDy7dGTIv1tTkaeC9GWkVJdWQSpKUufHkgK
OEJZc5UwguArzZKVz4aSVTMNFmNSujOKZTtWhSGkUEHy6wDQV1knSQEz1vrY/Lqh
LQETgOUDFvLnkcSfXY6vWh9nF1eJXo2cLWgm6XioPJRfoUEdCQMT9WgRM2rHHzSn
lxkErEFUihd3PAX77kBnm1BwYyoCgzBkYAQNExYjej085CqaDzUz5W6+ig6yXcEb
jNMWLVfHpf3HGf0TmCfVoe5vQPU0GhCWF9hDhdiGSBOJ5TH4TBzYmQfCh47uvx7q
cuVdlEZXoDF5QKpY/Xe8RM1cXFdyPH+vMYAkBZigfB6XM1RTu5WuF8m00JQOsxRi
1ZTDW0tg3WnhVBoER7oNB1PmhJSnJH6K2MYYeM+EKkXwh6NcOOX8vdjLDRfnwenH
M8kJw5oJL/EEGUQHjU1t6BL4OThWPirP3UvSCZBVe/qfNIeiVqVj5vHY/awP3P0h
nwTVsFqamoB+9jGBeCstp6ltZ5Jn8eIxjHw+fUrGWtOt1CjcY96P7fPHcvZJQ9xp
k6MwMcFdDyjkKgTUOA5unbI551r0QlAmZ05mEy/GToiTO3F/YgHiVf3N+GMUzjfM
5LKI54dhuqwIG0qh5NoZzUUKnxUGM7S/g3pLpi8iveU=
`protect END_PROTECTED
