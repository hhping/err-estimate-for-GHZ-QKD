`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
guNihufJQEyDN4i7C5ltME01wAA2sNpJP3NeRXgaVjoR570U0tQuIw2PZxjFUkyu
4NQu5Wum86KniEflPHuTEKOkJ4mtlc9nUXwGdAtC6ozo9qoosv0hfSy6YepwAXJ7
jg2IAkY9qXGJkWN7fpBiX8dyVRpHhPSDcMrR9AfqoBq9UNEx3ebvpMVztarmmkSF
qILH3T89S+sdhcgJt1Ln8VI/bGR8DWEdvWjbw7MNrL9vxUy7KHG47tPaaTEhUALa
FM51TYyZogC91sc7dzesl4KzT6RlehYRLtw6v2v56F2PrAgbK0p5XVWkAPgLGNdv
dqsFgfvsbQOEzrQ3jlbgJIE3bFPRhQ2JcxFcdHQNOIravu5/1uG/Xz82hPGnozNw
1XZVQMW5VgW/8HYr/SbAxuFC90uZgYKVH63oUDIY9rY/9mByMwI28aV/LgQWTK50
64UXb0Ed4BfV9NqH6VPE7f1YVdEcl5uFJMXeErmJfY69ANd3kfpuVD+x/hVix7j9
6Dn85LtyEuo4mb07NNB8CFUX63nw4uL2vKh1wMWxra4ty+OPL4koBenLrK4rnde5
/yNHdkbwSn9ClX0TXX6jkrhOhOYJuFgNr6pt3itPr7UOoNir02CNSiXVSr+zQ9UL
vht0pBD0rQlNsf2FGzHBlsaNL8Y8JOtCDaHjl48bUIlgqV3PpBrYKLKBnZfyh6X7
zE1r9R+pnrMcXS6fGJAT4oP8U7cf//hOPVLY7PUOFULmBlx28Fwd5KRw1SlQvQzD
/LI6I19ewbnDTKZURs5I3uL0A0J/s3D/mbOEITVKNBdo8WZ6ieS83700NCMZx4u5
qYuxUFxKVg9SGR+qOBTFZxtqiWPEsqU5Ybw9035cTKp62OxBn9osf4r9gIyggQ7b
Ni6pMKp3o7F8uTeZmcmoN5PbVdnXCMf1zDRcjOPyAQUePgbcfxagGGVA93hICuIH
KNb5SMTkmE8li2K3HYHupcHPS+9uNCLQfFnWrzsQX++tjSIC5SPWMfQ6BteLFjhG
+DLSx9oB9DWHH76Qq4sWAmgO7mK4cMMoLIPSvCZrraof7HycvkDun/DyDLNStb8r
fa0ggv9AnT15BxSS8w+6rFazWlUDVGDgkbOSU2SFTvQUZ7yv+QeEJ1oj/E6lYaOq
txwR/+jXgDJ4LkDgX0frQMuF1c0Y9L0V4VaDsZxG11JXqFxxLZorUhYm3Ylp1eBZ
3T5BlZ1aQN3bwEAf2UCqWZ4DJKC6i9yxrC6V7WxJ6Z/C6SJ4tEzkwpxTnb8WKb1v
49GvZ6t5fm7Pwmp5uB9I3TOy27qO8teG7YvhJDrhyMdJz3ZYRj3WXZl/BBdVDDkV
gTtXqz105hmJ32pbGkpp3GlaUcHORrUa+h4yQ5m5B3d8YmxffUwsGJKwdJFgxcKL
QfNDqCrXLQ0KUqfsdYv/2m2MXae3CFbZO6D8QXl/2GfhIhs+hXtlO/T9BVe6xfAY
kuabWNRn84WVtzoeoexRjywQ0T1BLatpIaIgPZzBE1NnN+dlquFkRnhxm8ofK50i
TJvpo0oztJKHcREyyd9HYLL01GRZwt1ZwVBY4VKAnwhNaAwoBdtBVwWHlAdoIRYg
8a7wmXdj/Qj17CxE7GyIcN2olOLPjapzMb87civNlkeqtBZN7hohF5CXKejyv9A5
a9eG8RjH4UL0Z328xARfaygUO7gTUuesPtsSVW5WU6NS9xqCx6pRZOJYbDRsxEeK
nkAvXlHX6jjVT7eAW12F+5NS80DFeV8BE7xGSrQwtU5t8X+wRPUJWHYd5idkXItc
1IlYbuWDamniVSwkl34aDR6j1/yeOm2na+xdCDy8d+KonL08BRre3wQD4S8I/f3y
UDHOtqbMaVDk5NpjG6FsE95UZnfjwyd+E4bRVabPLFlRVWkPsyiYufZLlJykurf4
CTmZ2Kkk426huLXgn+sTbQHOjY3uGwg0fe0/DMeNclPn5f3OPywCBdEwJ7tBGx7o
yJj+VCR0OBcKh3ccv5ySIHqq5C6kV5lg7N+dhSpJ2g5R+Xer2viLSABTSQvcZO1N
YDXqSPqGyvdejjgfMjj1MXkp4UgFwBgNcuJ01/2WNd+LVKNYv5C0xQM4yisntGmJ
GQb7Ml+L/vuqoo7tzU7GgPSWs0ylpJFHn3yMv5jE3Jio4WbMlPCBTVbtv0DHtir5
3tXK14gJaPH4Lih0jP1+HaVuI6ro2JcwtxcXyyt7hNuf2GVgIiK5WqAlnAw+/A+v
PS/1q2WkZSeT/Cz/bU5VZS1wqmPy3D3DpUuQP6kmz5kCub2ko51xDUg73z+ZncfC
q/qTRtOXsNeBtDGEbEYATL40/47kPjO40n7PoI5AB5C5EDDslEbOMLY0jUzSUWKJ
8l2Rhr92OpDi4isVJ3vbf3OqfDgmQJsXopdLUJZCQHIA6J1IYnbBvqQCfqSfYy1w
xMij7KsNoXcPShCH4IQ7BFt+CSE74A/jZ5U4U1CzFcq9xacl/OAGGeBZx32Ajaqi
HwwTKFIh3mu8hpOpRo+qIYqZQ1D/RjodkW/lvzg2P1JFfkCNUSM5dnK15MRYBwRb
Ee2fOi8Om8+y3QkCNmYS8dfnVS5SdIkOCDdffEJmi/0Eag9JmrlSYlVXM6tKhfmI
htuk1U8NC+Ox/o4GgpBxVV6QcrMDkkD7Q5f+sYmECSZe9qTlGq7+1iIdGxPiKcrT
UJfWTvn/PdRePpr2eyA3yt2kRCuqIEk4bQ/JDFpwcseu0MDH94n9xkCCiaR97ZCl
NaFyvfs1wivMCd4VhFNLfQ4O0AGbuTfs8Zr74FfG55vmriHtZEKinwf8bpXzakWv
Gcv0SoMF3m5emcNjSlwKAi91nMVaaQ8/zuvTGXDuj4Hnoe/n33WU/ytXhk69OVrq
N/Qaz87LbVkxQilLOA0hwi+q5q0GBsDNyVIQgJ65EZvAbAdKW/AWRiQT5ezIfqf1
j360CtmsBKiXm1HLwzOFTou6g3dQoGctzOIle1IQgyf9970q9WcyBRd8aA1YgJHO
ngWyEUywIaLkoQn2jgcEyBHsDRCw1uzswTVneNbH/UOo5lj2EgJmAQWLZ5rd8a9z
l3erZdzdRhR8DgelewWspMva+wSvnIKZ+1KmDd2IjojMjfisnDN6JI4kRqV56OfF
c96UqUvCqW8gwia+hCbamUjnw3eDhbcthKkKEchY+XNbiHvJir1atGiwXbPbhX69
YHqjpbJF69Me2143MqxRQ8RNeVWLa//vPLGJFudjctLwlVS/j0AWyYopA6ZmL0cO
4RWgpgmYuldvRquV/0X78FLkulrgUr/NfDyi1mgwwmS+FT8Su1tvO/Vnw4rh5sVU
h0Oo17wC8nx2yYFCIuZMRfAuQWd3eZmZ3kifixQgk40qEuDVwSBBRSd4509yThvV
QlQFHsTS/hXL4Tdic9fvAPkXsGQoc8L4rBOdEGpnmyamDIhqqiheLPnf0nm9JYa2
3xX1MY7Q7ef/cLE3t9B/+fbSYRnL4i6Y2JR/uISDDr1Rcb95yC8Os0BqhszFpE5l
rekzC90/fHc/3771bnbS7Mnt9UoU7VFtUaAacF/A6xH/qIhMTKtuK4CjNqutcAEv
5116FrQspHL9BwVocAIqNrsmNxHrgoO0+astVs8inqtl8ZGoVk5qAxO02SL2q7vA
ISDXAwQ9FKCCgLIAwvlfo2c06rWR6h2HK0DldloLxZQHap30YrS/89by85QkO+FV
/Agux6rb3ZwHMZg6qGDE3gqHwrwBn3skRhZQ30PBXBE9CdS07hcW3LTaVZVXAjSF
H9zKQAZsGqaAChcaIE3vQHWrZ1IxobbSrBJRnf7CwqaVi3+aq5wg6YRI7GOt9Faf
9W2SCXeVET3d9h+gmE5JgRtI6idMF1ve6K3/4nlWZbs0pIC29omdfmpOhIhMyxTb
epVsC8Y2nDBCzVALqYNaX2MtNS6scqWf2SfA8Jr2Zr/ugGq6viBuPXmkWfxj/8ga
lID3x410TQeAP/kOWMNpVKZKZzFDjoh2FUTdKWHyVJom2fPYBaGELweqf03b9mVH
HHrqt3RcxDU8IxhhDeCN9gu5OUxLK5nCPgSwvwfcl3MLFUZ6ajPsC2ynIKLY9gNT
imBWUdnVZFkhUYst4BD91CdWYQ7sKxsd2rcfVi1lu5JF8kl8LoNLfOc0iNCQg4zi
ldvr1nC6r//ZUFytHKYKh8EdXicMYPkpEL0Qc6umlSRYQhyp2Mahrle7L7OjGAtT
0YB+BQqvWk4IYH9B2J/pFamEr/UfzoUmvvecZw7Oo+Tfh9ZcleHCeyxcAYa6g37G
aTgpRV+ariZSFdnJAgpehsgmH4GNklmk/92GqzAYC7RQO+D7zzYffLMO5hmUIrQL
LkB+wwIpdJQiS3WriYzRgf313U7hzzTjSCH7LzhXf5zDM4MVBXyQgVI2yYLP6Dp1
9w8+WYBBlC2gKoZYdHzdfUFk4GdWg0xaQe0gdfPN4hrIL1JJo6ls/RHGijVItyEw
0wT7oZgtVXCdR87qermCMXseVQAfVj4lUmMBv/F3BSchL9c+7wJh7oz5yMMLLG9+
XGRwRb4TOpjb8NBjrAhPNMyFNlivfY9l/WKmYot1qUqB1de6n/Xgk32f6lG/mgNZ
e4rgkGfVsF8ipEohTXfTADU3A0jqFIX8iBf+R9QEhCu43P3uexBM8sL7HaHKtzVG
GW0FGqd1G59PejN1SnoiZIjiw42aQO71X4w7QxeJ5UUCWFvqlxUybPOjYzlX4vwx
KY6XwJTfiuTq8uIH3eIxjCoueW/cU7i/7VnD8NA72J/0DXc0DVN83Wj9+56ytkk/
EgT/Fe6YZVRkvjwStNrj4gEBunrh52FS81qI3cfrxsDwTV4Dsl0/Z8l/+k/NVsVf
GwUJpJBr2Gdi1U50aIU/2bvgAqaxgND9+pbr+I7gP8Nmv2l4ecTc3iTCsaAzI/60
fpaVJzyWfbMz3V5mhlxfQgVkn2ELiQ4aI9TAbJwmUBoQyeHzpf1OK9Ix4Mg23SzI
OEXGEGNbDGH0wHBKMCLZVWM0Y9Lqz83HGAKOpZDXubBSmlW2HLQSfuHqt8YNnC3N
J7rqmFsR/yVjI+wN/v9anhAlYN6cBDag3AJBbKyqy4EYIQUJaLujDOhYsJCfnbis
MTiDYMgH0lcSTsKCdpbrgnMSmlBxAKH22Hzjmk0b8q+pkfNx7UkEk/b1rdb2eh7c
obwl7vqFlEQcy2DZjhxGY2oSgTs5UJJgM/k/MsMUBLnl8LUkYynIpL7kWTmrkDFl
UrPKf8jYiJvX/3xqYBowsrG3d0Z7cbrW3KSheX2w5m/Fj/lK1w9YzD3UV16Nj49B
TYMMHCXmJsyc+TIZcgIk+UKPixvO6DEfpCXMWfBgfI0u/jdOBSftF3SHa0mEvgpV
+lwkBS2/DoCUIJKdVAWCUUUA47ioUnPOA7KdyKoG8wo0bRPZThQnobeiZiSWQ9Dg
qYmRxJtu9P8Fgz/r7+Rvoccvy3jOm3BwM9xfCwyh10YCmPbP9Dt+8khnOmkJ1q0a
9dZpRHIo6Jbhltp0ghVWysj8b/cg3yN4bElYrZkrfMpRcmyprqXQ6tXp0S5F07HG
s/zbb38VFh6LY6V9cbYGj7Y039v+ysNy2TnIE7e46j0=
`protect END_PROTECTED
