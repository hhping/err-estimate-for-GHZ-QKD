`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQdlzgGx0WWiaRQp6sJ6jk4CF7ucUZ3Vo8F1WRwTcZSU5dGpl1/jgLUB5RPU0u9M
AXxNBcCXVarYzhLEj/9RxlN1YwaoaLyMb4NLjdx7d61rpu7r+u0hr0rE5SyQcPGx
0u+F1SFcGYXgATn7Nmq3Vu2qlcs6cscQo0dD0j4gXXuvJwOA62ErMvHX1GZ91Qwh
7TxG8f6ZM+aO3pmC7JYACDsgwWSJ4mxV8USMHBsb88hGk85Rsn5fDmdli7ew6H1r
0D8jRnBRPmlmNYdFBib7xHKKXIW3QGLaJsSvvKnElQGSUpUSU/EjKJpNGBdosyNz
9J/cxrzKr3/fbuKA1TqoUR5UfJVVQc7LaeiDmOIIUFfnaUvrdsjQr8gOMF6pfc8F
5zBjh+FBrXTFauFNn9mva6YoB+UlPAd91vjxCOYM4BIETHAXv59DXT5/5gNUNvlu
zEMPuKG51UZYNoFwaIO9vn22ujrGb9nnP+wFHo1iAB9/6f4pb/EoOFPNerwZPiRI
wyHkNCQ/9K8X3yD/r2yQbVusBXg5Yx/I/oUYU3orO/L4U9CYVOgxaK2/KZnSXOSz
zRAE3ul76+4ULKt9GCLMLNAUIkihh6c7Wkv9iyqab6kBzT58xr7YycsX6aNwtzxM
I7MR49ajuHCeoFZv2bxan9A5koKwkvdJqUsZdnuEaziVwRIPE+rG3tDIg4TDemFC
6JNVRFlYD6g4dwgc8QkFCsywUlNJDj6lL8jWNDEtY5SJMcP13fj2Zf1fFU7ysZLv
+eWTZndSof7W4B+MZVW0NiMA/UskGNhyXwlendneZftNOTcbGzZBXxqQPrXwwTe2
7z2Gm+YxJlU6Zub7SeQ5s4XHVEzXsSmJE05Jl77900pQMRV33qcg3OwV4KL9s3K4
7jPVUVxm5iITgi8NLyM7sqyLjCP1kYWDXDwCj0eH5WckPjUOKBb2/yIZzsvMUYpV
hDyP+r877uJauWpaA+QSvR1dpoVHWOZ22Y8y0kV0kUphcS209si8buiPzU/X3KOY
DcQtv530BODwgmd0DiC3GBV4kEw7DTuIvCzMFAWRg1gxz9+B7pkcqnwgPJzs/EoG
pjH22+gW5EK+WGRH3aJXdeBkK1ftfaAfVo6yLBvvtwzJkSt+YuUoSaoT8+NJ28f8
TKLQvKM+GVmVlPDc53sC0+AXlWconbSytHtCCGBWpa/ag5JwTKB1b8ICNz1V2OkY
X/HIhYCEPW7yjfaZtp4h4oM4PVJJNKX4YsFAY1cauiHkpxHnydky6jveP99YesZV
YMi3smqcVENkMw2jbLmVokGVA3WY90G9+On6WW5DExLVSRtUIdfndvFIe/fkF7qK
xUEXN7QCgkNdwcyXKjYKT2aqf9Gl3MS2wXOoDmp0MF4=
`protect END_PROTECTED
