`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TR/Mdk9lnR0L9Dd3Lurl+0EsoWTMprzjfIi2hnsDASMVlV+vNkThIV6vIPzRnSWI
uIDHv8FquKDK7ZjcShTLdurJOjlNsfcxCyvOP0wKB5Mf7qgGYYEz0jwIaAQEG3wB
Auh+o3qf9haQqLQ+Mkd+QpmMcODFqQbUkgVm/h1tqbP0IYjH00OEVen5nXxsi6qO
Bt7cbJJgFo5jT8QWOf3y5Dfvgs8OzFosuDnBSx0hkmgN2ue9UnPoDZf4FPYjAfdy
rTrBXgMSgdCwl0E/PbPoucpVHf1czDKE1RiHnTGOjNCE7ZSrdSswzrp2HnlfB1dQ
agWAp4GCjU/V9fjgJ9zXJ9y2Yk5PBFJTJxnj1sAClSTxDvpeedZ6WFYoqQVWz9l0
1lrH0JlOVAcAqid6x13cGkPC9oLb9qGrR3TlUz01GaTa9IpdBwxCiO9UhQAyvoDh
qbsYfQS+CyBiQ8n11/WTABxOWcXvvhnOhCF2plMmp4DzRHaxBRnWMPi0g4ekOjMK
u6S20ap3gw0RPMqy7E+24hxYi54XsACtmxRdgUBECrhL9a7oXJJuz29+eiaA2Vor
aKBdTXiHINTxqjLlo2MxYv+2zrb86TolY3+Th2xSybrUCIbDwZX7hMQSAa44l7MX
JXjf7Jk39M8AoLsHSafTUAMVLiaNVuC9K6uVx+Oj6AvKf5Bk0qBc9gD2Co+c5BH+
DTRUgQwMklogiEMqtZhVFnc63v7WhvaIvAMQHcyorxOonqEJjfFzpXCEEdYEboYf
mh6r1Qg/slywJag58NDmYSzWi9pORs5onVLIQI0hwYG2tnTL24t0UnmSoIiEfIPh
bhZ7djROWfnvlWB552K/2E478OQMPZacJhfTIhr0ZUV6dA7kB+K2eZG2K8CEbGrW
ls9h5XmRSfSLafxj3ix63WbrIU7Bl4/+ihXFTygpFQSgYZtYo025W19xcqHQtU9B
GzrbUMWoKBj0MJ5A/UdOqFDtcyn7raFvf1t7IYZWLOi8whpxluhXGVqgrj5XAxPf
6Ni3dgxiyEny3rm3bt8zeb0J8Wp6DbkOD2pHTK2vd532yBbEap1LvzNsKbep2aPx
snYED4tAezViV97TsHbzqBpnk7Wsevid+ZuKegZbnnBYAHAmmanvDnG/aLlPNH7h
c4K+4sBU4rvlZbxDaNO/rW/Ua4V1n21epGehOQpzqAdvJARf83xZM6aLdO0UznHt
WUniHFYu+E5C15mcANnxlaS0dRmG3xRMwRHKiNlxmA6AKYSfx6Hv1dTfoslvBlay
haOzcUzCLIuAM2V55muaKpAkhIsZvyb4swvBuVjyX1Qj5tbLjP964UCgvmjzwSJq
LawS75+is2skGVCvoALzIZk2kkujt2CBqpkzUmoXYKNQyPaIIntC7MuhFRD91pt0
8STWNLf2JGo3QFcRH0ux92pX/tohAGfXpkHzZbiA8+wZ1GfZYOMzhE00rrj8WpUk
pf4rNzwqQRB+l8DeW6y129lBXro/2z7sJgKGpNJSKdRsIQ63bBSmfJsKbXIWFc3u
XoeO7OK21wECZOGvQthsL0wwhvKCnZ2QPY+ZYU9hvogEL6K0F0KD+Orda1dddpED
02q+wVABqNzm/R1AhWjPXNBBXPl/+wCwjP2gLP5mIkud5PRFm97TqGVIuIE92UKr
LzKl7OW3sFal3/isTPRF8rACHkc4vJOO/Gw/apOGNYaO/NF8grvrWxdsQbjIEl9d
oKGMcrmMlKdGw2pF0LWkhluIWZBqJ86KzWc4tA/ajNC7W1qJyjsf9gDUEQt7sBcE
gFaucPCJH6ouLDl71RI8p+0loc2c7KWo/47akgmoklpyvENJ0ZIw1w/DWfHvMYNC
O0Tmm1cCNvHN6R4rZc+2kTQ8VYedpVH9Ce0YkNfYz/4vtCIfuxRfQD7KjNfzMe/I
DSK2HdpzJ0XAFYNN/B+8eSb7COlJxSqXKEAP1o0VHDb9ZQ14JUzROdpMniAk5H2b
UJFqa8XRlqA0GSzU6oMhgjN3qUgI6w5VeIuJzFw5WUBFcGj4kB1dKLX7u9UHxTfg
p2TsLByzmZbLnqqe5PcnrO244ofzeVa9xIHynd65nyvqfpXpwEKO5CBmQxaTFdrv
eNJNQECGsX2rnnI8qA2YXKy0upHKNwqfe3ldozHoXaE/NOUPV9Pj/iedJ8fGH/g0
dKzdRzrNQHHrfM4OG+ZUohkNKt1kaaE4MHDyfYhrtTP7rfequ/bawHDXp0zA8TVy
nXkfq/1OupVLOOXlY8OqEPrapnzhhI2O/GnpEV/B7suRHVRuGZwlXgQAkdmgLVho
sSnrrzSWg/cUJ2KIVh33JBw5ncy4HRNuDdkDvmFsuKpLR0APHkHYNrBHoavrKJIy
ZellMi4hj7RRRXzKB9VeZMdkBMF8R6RWbu4gVhGi2fNAZ4OQQmm7Y4W26AJYQHU8
LV3CAhDcKhwsdQUlCzWBO0xSNDR16DFhuY0kPY7iB242En+fA93YMZsmv85w5T+r
FJzLu8/ZPQWaIrN+Ehgy4GbW1UeMpYz70M/EQ7OwVSrkWj/6F4B35Yu2yuRp9FZ5
xQlmejb/jVuZBXmiZoN2UsGdVal3E5YV92Lxl5nBqN2Fzvc8dMTC9mk5xlrnm/AP
nRir23FlMeUGB6ws5kRpWJbTyyb1ylSywWMdZpMzoldeyWpOCglmQL0TFZDF4UFA
0ZnJwB9lw0/qmCK6MQ6nXukzC1/Exl49ElBwMJkINFnoB1Qy3V8Okmk15PnuqY3S
er6t5fFaddcd/5vH6snvtWG3ZO/gtqczedk03KL5e5I8WjmNfAAtV3FG+2TgEPcx
I+w8OCU9GB0l9gqvxKa1Q3oNJSpT81WC5q97SVKE2oekbJOADxlG1it6XG1OQCme
82Fndb7WlVsQv+izdwoiZU/B+aXv5PrMUD33y0SBt2DNmzOEwO1hYrwQ+tgJAPos
4I6D/UusWgrlN3Lv49ojbNDnrUcUAFydx/HdyE8VIWR17MiahpOQtotWg773YfTq
wPqs6EosjtOgEqIxv8yRAKSukK7nKeQ6UZQmT7dMoFdOYuV3shAxuPwSJ1YMP72W
XyVrnj2wVZLShShSg8a5ab89SfbDIBAzSMdGWrC4BrQK1guoRIQdgaaXYiXyjbFr
pb6ieFNGeb8RPIkQaShigbM11qfuDs1sZrEUSRCL2g/yxXB4WdFr12z/uy+H1GWN
vc3PhtP5zhyRmLW+2A5IbWEa16cwY7TjoxiUGg0/2jPLJ36QPccqonTkiTW6vREz
ugJijo/Q8xzb0gnWv/jyMu7Xl5THuwgcjKEOUkhhm8qZHQGhjsymehnTKlH7EJVG
ADyDCTFaBcTKDZ3igjib1oLaSCkFcfqbx5av1po83GQIxJTQ8jcU3qdbWifo0ZDi
hCrVE71hERAWMACtdCNW4un2u/RkGv43pUbBxFC8DUy+NTQbJa2Wn9w8m+W0AyJ/
vmZfNld2M+5eiEbz8eqgKySKT8VueqSK6B1CRxzLMxCB+uFViK5nGruExZFg52qu
pdGk/1o6EM7w9JGK9CdgJ2Y7FSuNdIUtVQXXZ6bGH4zBV1cRLilv+AAuGYX2FdFb
Wo0+E7XL69O4Fyw1TNEkC0DBakF/PZCPPak8KYo0aNyMD+MAViYpPdYBpRP0w1wD
9eVqm7IJOW4gR4RU5SKx/lfWMPmFn8IK+wLBq657y6Cq7w6mvkR6W/pQjfMsdCK9
mKBbZv5pkpHG11eAAOJg2w4rJovo8zXuqH9RKdAZWLU6mPRGZGHuNP5Vb5jJLcZa
xHo3sORfYjnY7s6kOUXRupcvM0Ex0dTXdYjxaoGwc5m8iTWluFV74OdmL8zIBijr
vgQPwQEc9+hrW88oQVmnzPzVdCQV51DV1bheMrOKwMItKlJjcTLOOCe8B6khXJCA
hELUZgrBbGZGdkssVxumiW3DZMnKQ5/MC0m54cCVZHsJcFCXkbs3soHHucRtkd59
n1ANhsixhGGVqxoCxMiSaR4tBGG+2YkHlw/srC0MQvX06iZ89ZDaWa5yA0PRdq0B
Z6GWSHZxlFiK0U2LH1HKTETq5N8MfTnUzweBQoNyKgXjPDSUoL/ZWTA0xi7Xp5pX
ErR92ZNrb+6NqSMy6G13AyzpNQ41+6WsyUsdMsuVrTl+X1PPXRegefgQhHysMYN7
AKt/wu1a0VmnXhZQuKIApns5LuNjx0aCIGwwO/Fx9WMS4Bd+3oPNLILnGBGUBvvh
t3ixOVQgTEVgLk2gWJm6FSZnwqmw+IJzZ9+PYk86yZVPoTgmHmCR+F9z8flmIxxt
dZJB+/9oWr39pDqHrqG5k+tPI+go9fCT+HnfjSE1fwFw1Fxtu05v8xhWm7dXe3NA
OzzprN3SRYVDL0i9oUeD+ixmnsABZlDjy3i6UR3aJbDPV5TQOXQt/t89ZTJiKyp6
Vwp9R1Kfl1yGyrVCTfr58qBh7tkcJTTW2sbM2bTZKNVnCsrZLQc1vlsAUo8sVeOH
goWU17i91EnDQk5r4fROuR6jNBfW7hwW3MOhHGUu8CtobWb1cWF+5ibMmbUx+JQl
AqPN6+/E4ETostbOwnAKz1gO6GSktPmFEuq9+TAEm9EC7jWKx1ip7AeLPKdSoVzH
NScpH4/Rf3hR+5NnCVph/kIRcKz8hfixFaNMGac2+MnSHKhy6Rhe20EYfCZM+AYP
tJebCgoPg8zVgehJlxqwWc4g8yOsTk1oEixeBUVZXWFGmSSLox1PhGt+TgPl0Ej5
Yjd31AEuDMANPrqudjfh6Nyv33BU2mo3RJDASWPiE6q5ATymC8wuDsFcHBABVD3J
wC/qQIXZjofSbiu2CHgmyUnsbcWe2cezym7/G3UzLAniOuFxLdKO2LbdJ1W7u1Ti
qeLe/Tlodadx6mS2mBvC+MopIdC2DtH4CWqvMxh4tqt7xU9KjSzaOaWADrViwbQF
vOZDF3tfWhYilOfNT/rAP5JQTRN3G559U1hfMY14rfhsv4oNk3sV/D7U5mr6fK7t
zJJa7RjHZC8bqWA1UnPGZX1+qfiARnA2I14/dolQKK8+KFj6psITYv5dRGwNrxSJ
xoRgX7rb6+Agv653JLl58rOQJrWXu9jKoUTUx+n/fmeoknEoJJ7wqW3/LbP3snwo
4lu99HOXQ+tjB2peh+wrHUUur1iFz6lVW+gq020J4EkXMGhc+eRy0rZb+AvFSoeb
HrLdCjHweDgbMcrh2+QcBoc8Q0ekNTtnxV6vaVE8RN8tmgA8XemgQpx9K99aORQt
ZEyZmwLlvq1sGdlr6huav6bSTMO1yEinxHXWB0bP7RzTKJ06vIrzs4qhvfROeiqJ
mqig/RsLxh7sIWnN2B3iyjadKEv98AXKfJHNHmv4K9o124ZKORqMMO4y09KgXYyd
alXsHh6hT7E3Zcd2EsHysAQz+0B2uia5iZrJarVQH4dMlGQa5qd/6u9yLSFl9H57
i3qLvxm3iHbgq4vimYwRIB1USrNeVa/DazQ2+B5up4KMdbSK2h7iZ4zKgZiPudov
zPKpdzw9inGBpNuN1FQEz4T7N/c8X+V7T03iidLcUmbrnUlHQg8lVA0eVwmegKM/
Ybpv/QH5Ig330eKf+D8RsuenmtIUnx6NJynYVWWROZjrry+/Ui8dHasPCQQ1+vC0
mNZXfVHma/QsyskJocl2z5bjZBRXWwrOPq//tIHj7SkzPZhDVdZsCs3s35q9F+rb
DdbBDyL8Atgysr+95oC3xoyzOEunYqiyaWqx+0iTft/WYnROBN4hQ3vKarTeiD2w
MM+3ZiTA5GEz8yUjMIeIpEWvixbNwLPRnbBdfqm2JiqRvpmPd2J9aVcKsninfGqK
OywFkPr77Mg1REZbh0CNTR9JL+dLbvoLLXZq1X7mHsWhpd5J4rCDQrHmh/FaaEPB
cGLBYNEdb6ElyqUZjxh+MfTal09j2W735jenhKWcbYujUvPfrpDtGQXFZaDi5rlc
WWAw8IUKLwrRlHJ8NFmGjz9HZiwqRsFbiEtHmLgwQag0nyBy1VyUrpfY6UNER0eT
FWStea6hrVER9cC2IYgONDw6lYSJHZ5WJE+EIgfFdOmX48IiZupBemxrCKwoaeX7
zF1QQX1GhAPxg81WlFdYKerotmRRU98V/YzNJb2XIMD+0aG8tdDkoNIRmjJHLn6R
sJRNuT/9KPkIRcgV4EEX3//TPDNLbmID1XtfqFS15MTQS6uO5phdCOR1Zw8Lw6wM
FVYgHN/Czt3Z7lq1pCZl+p8nCq+yR85lvDK4Y7j6J5FVhLw6+j4xieUv6kVH7jcr
b6/2gmVp2hqZMZHC5boBFRzIK84avpmIz0Kal/YPAs8JUHqqO0aeBkC9ZyYHrL28
UPAGiahtR4bmlRSEmyhzCEC8bVVFt5zkJ/wE2jZIyTZULtrxYAjsw18PXHo+juCn
77TzrT1TGpSJIaEg4nmdYJy0p2qmEmkk9i1fDV0QzWFZaQty31gFG/fxnaHZmuSk
qful05NQueZyyr7f3V7uArv9T2Q2b25ME0Ogous6Mf+lpu08gTbBEMoX0oEL/X1N
zsqz2k8Hb27QFJso/Ccqgr12t+k0jxvSD1VyJIIFR37K334wU7aHrA/5nSh3vUWB
D8jscpCgpwgW0UustSUVZxSynh+u8mzmrUMU7Iq16WbibwdIos6DHRoXDFElMBKd
iTyyMEOj4keVOUBTl404fmXcJ7MvauULmp66t/B06544na2n7xkGN7QE8CzYFIfx
3FAbtCUJtdY3WRkRbWPndHDL5ZPCjFVCt1TDuxQ1OoAzFyhLqjVVXrcdl1lSnEN6
Ubidjb8u2gDBNiSgLFA+/N3BkzTdb77q3fCpGGlqkXBF2x8p6zhs8UNCOphpOlzM
HsATw+iKfrXshfw5cjmvoISBv2nwCRWar5te6ka7JsHZHLDHceWPvKCq6hEJkmtj
Zpb+iATQc9yoZEdc/CFs4w0xiAfoNDuWvf/52QQ0+zW+Nha8xHcBi2VdlDsrpwhW
VEo5gjTZ3HAGCrskaFYZz1vEiUWL2N8kbAtcLwFAD5HcmW4ZWyys2ks55PGk4jyo
GuRD2iMfEa53XGr6Lt8W/FsJ77ovNKm8I6VZk6lUbdUwvCN1XEcrRU2bjK23EEr1
/8hb2H0BxHnHfCVD/RODjnt7kyhfWyEJlimpScvOmDepyDi6bLUkDXPbFgvyrUHj
/iw5A4wrx2caRNV19SQ8Lgz1QyCW7NRYtFaJ8VMmmMUyiOZIrblttIVjC1uNJLIV
L9QUK+r9E2hmy3Az8KtTe1SOoCkhX0W+qRG79wU5X8Z9iUZPgldOuM/0sh2BpQVW
jtuCCRT17y6FcsVqI+k4bANRVgA6V/58YGcVJjPb1VIrMFGPKFXatkAIIDb2eGqW
RZrOfASvF4Yq2ENKUDiGTBRPQ9EvQfGEf2uxSXB6/3XEWeYnNwvY7zlpHqqH5dZw
6//id0zvlHEsb6fv6DQ5Ylp1myzuVHQ/s2rB6j6IOMeW23OKZJSvhOd2jtSPCG6/
ODhC16IC27YHY/AZz2++9k8EuRwxViq9sOtr0kzDXGVbrRlxktDVltOeMyWClFO1
eBrBXoWZN1KOxYweslXtiybGPfMwtYh/tjb0iONZH3Ga6xeAVN9uUmIXP0x3gwRQ
QLj0uHZ3dg53LYsN4/ciPYbxWiSQHdnLfjpdQB6bBF+k7KVilcjdq4YxqPb6hQrK
S9FAsxRzeo/cr3DZzCfuwyUooJcjEae+OeGvVXMnd81yMH8uZXujk95VTAh5jHh3
LGJujV2yUrShve2k6golHwN+ggNanNhq9T/3i4ruesaJf6e1O+Gih1BLvN9ZSRUC
XPh7dVjWkSkdKURoJsa/VEkouVmuBQJDj2Jxrduu/6K/z2u7/AwWNyee8w2w1qi4
/StdeNEFewylWj5ydrtK1wLy2SS8VlLeJc4e+DkUKYr3g6p4oAhSJ52X16I/b1Z+
PZSS1ii2BMkx+DmxE7mVGc34MXn1iBaZmuFP7UCdmBC65FVR6wwXEJrCK7wFS2He
LV97sr9mheUolkwGpRK99tD0GHuua0zU9lXcGdGox1o8wogekfRUyOyFYfkwOJO7
dnLeghlMqLoFlsNsdAGNghyh3UvOpLBcQyvn5RtjGALW/FcmcriKSOJ8eXtLvkjs
1i9WPIqodfpTnePa7dZ87kJMEaDsBsWaoHTud8DzYFgd59Y0oafKNT6llzDu/SnG
/X1qNmtwRpic5PBoJxjBOIetlRmx7H06JclGTDECK0tAuJRovvnXkJ08VKqy8YHS
T5prXXFot67nrs6BsxYgnusoT5JLyKqM/2ZGRxVgudqv921GHcRq16tSmONXZrij
oAgkH9Gtl66/ECL1M28YqzrAFkyEjg4arnJMbLntbIIXkSKWu0QW7ViTndHpEjq/
2kL3C8lGFP2b/a8mKxZ+dMt+OiaDES72JZVdYNDQF6W0opjWTAOQ83INmCUsPj1T
q09uCrEihRA7hzSnUXtTsKlpsamZEo7/WZH+HC7bmRLSy6nV5VAX1YzRNv9F93Rk
EszHUgaLL66REXO99B/jYnRh1ZtDZnYr7WwV9GeFXn9xU5a1XHRYM1VCzZri5DJA
usGxU7vM6GG4rs1hXm9O/V27NWvOTQA3Uv6Ic7dS6UOAVGP1NoL/3SrIUb4Jt4/B
C6sWfVo+EySgbEPQLsSwS6wuXYkKZwEARWgeI42KX8i27cEBnwg9jM1AdoZeK9bY
tFA+YPd4QYCLYkPMew1ePTp1ohbe09QluVxG5kaCbIv3crx2bWZ81u/AEdij8CjR
9AgnDgcAFNRWS3TScIx0gzo49yccugWb+v5D253CL3UyHAAiBvt7AOcRxleFft7a
X6mCed3uRoYuedvPUn7OdIosnqcnL1ahf+PcifxniIptAS2H63c8AG3xZCWaNs/Q
vV4/mVYDQyRZyHZbOUqoy8zQM4dJX5iM444A+PUt0QvhU5OqPqEMn+cx5vv5/MqV
BCHdszCFNp21HKiT7AKVk2XZ8aoppjXcx6cERDjoGBG3WuZWKF0kVPnOpAZLoGbA
XLsFQByy6VuPxGvMo9C2ypXTGBhcy1uFDhi0vQQeTT2dZDZyGo807g3BIHt+rSkn
J6czBjHpWNFluNqmaVKlnbSSh19KlO08zo3ssIUhUhgY1oYK3mifmJRLUn/ObHnL
1sWEQfNI5aQtYsnMnzEk0JUPCcGo7t0Tcc/XyjqGLx04uLvmGr+M3jOPPsdpbo+A
zMqtuxWc+rUsei3Rschluf0N8rUFZQzUw41i+i0SVU4bXA88TrfqeUaJ1oXolO0X
Px8/T48DvU2a7VjRdpoeMk1bQGZdbN6tSwmaNm9uiDECeyZtUWK/PSZRcT4jogjE
qKdwMyreRNzsv8z6lzCbEmOX11jb/tjARblAd3NbVfYK3c7rDC90Crx0Q4ZVWObG
Kqn+GrEQcndnR+w2OrqoW6p4vRFwbQAIPPVLlD0IkR4l7oMVl7iyteRu222TMb+i
Q0gzu8bioZeDQg9PXyFkZ4VCA1PyzSSjIqC45R5otlqzLvWUZGX4IRwzXYgoI1BC
gLX8VX6H4OIO81sMrXliTdq+eskbNBuauPpEmBkJrsnpPdGuCwXXcVHBjgUfUVsG
1Esd5xT+thuD0EX5UCrbeTbtt893vce7WK0x8ITll3YptUfLU/PNPebTzc9ngPHw
MrpcUJmJzQ62t+mKK6mFppDFL8EpythGT7LfW8FjD/Wv6Gp9EnEYa9lKYDhhqu0k
DhClUENJrwUOjBk6EAS5aXpanTTnRzPJqHi/sH/DNKfXONdEvTfPlwBGplFagkgH
sugJy7DgLk+D//q9eACv3rmM19Xq9lxEU42QM5er7uzWzNpqr+pnkIPLdKbQEsSx
hE7NC77WeHlU+B3i8DMgCd8SVWEw8Z4yN6LDizxriteAOsGsDvSse8FbeJohbSQc
JOu9WshcSvP+0Z2McWNgL2B4NsMCF8zU5yVY9fqPPHFwn8fiY6aootr2iyofOkaW
qTNM60mzW1GovtvrmDe4li41InIE4AS29m+jI51Vp8wnGRRt2qci8M/5CVWrKQ6E
lLecEvFT0ZJsxFCvIjA6YPdhv61neMounWiDlqs3dgmAZQsZSqt60i9WeAco0IDW
rAo3fKPPLa3CDphKf5/SozMDuiXOCDpD1x18iRNzMfSv+k3cIMPYXwV0H0wret3r
j/LKNBczT7NFAzj2+HevFY6egwpnuCywJ4GwiUNVIU6/h4/FLRZxCueH0qvMHTzB
rxcUvggqwdN6QRhOheLOmgCoE+0j58SRtqoOi93R5pBfLUDMWOq9jvOmVFedFE+z
vyLYx26w+QbIoyB3rDs42zpzZk7xlnoSlCItp4hlZ1EOhuWT/8IANHdCcw0IPPSl
W+4ZVIa6KVfXNeeEa+wThVmdxBLWplwpIBP/kvqMyi40ix2d4Mz4GembO8X6UGy0
3ezzJ7lq6ib/fLNZLb5D+pyJswR/XmF2N85liRLPP3sY44Q6sWNcMmGxFtvq0t80
CHlVB1FicI6p8dP0y4C4lBQC0fOLupJm/0qlt5ZwqUgruLTwF3kzAXtfMBTX1uPN
oq7rkx+PBye9Zs6ipV115VdlBUnzUOE82DvJSadkBMO6Xmx33sKFItIXP0AayWoY
m1KB24RbOCsqyC6cdDK7XaTw8hzMH5Zpa1zRsq5Co/dZaaL+j5Bh62kywK544x0k
knneIuGeUN6PP5Y1qqWeLkTuearXOJZh7yw75khAIex2e6cX8a8pFDJCjk1lk5lC
fqu4qFDbrS9YNzXXWwvIxAAUvwfaZTAGcND4TMLtINb3/O4arbgnotlHWz2G2Lmj
6ayBSHTfaV6JJOIwszWZUsNWYTlOzgil+M3JMNiw04eHMeS4stGskzwfeH2nkpxZ
RxrBAphog1zuDyWEBDATNc9Of4F+EQUINgdGuhZ/5cp14+Nsgfccetkk3yN5+CUt
ttT++k8hWJlrBbnnm4xu8OPjv9CqEMuR9+ogpwQhdKQKh/wGOUTpAL0ldiQ+KJRS
z1sLPKz2jqzIuki/bkzLSc22ujG1KJLwAwvVUPwPKeJIjBNCJLA1zVhEUb/+nRxM
nJQRAZe0UFkZSk0v1W59M0bAOEHUTlkW54jIWvsSUVEIG5WtwX9pB0yzCjVw1QIF
2t6pRKASyKmKpwBOmNV6o/Y9hyftAW2sBmSDtfKrzSWNsmiwgSkB3nYCboRJdIF/
f5G83C44zaspU4OoYFVrtdsY7c2YeTm7XNwj2dYNA8f7MRIKo0/ZrXayEE3np7zY
xCKRowe9p83+etD7WL2LOmYJMKFapxJIBMD1lzk4eqILgNXeIjNZAC52qAd7p3Hg
TCzSDj8EzTV7VmK1wS0HTh3PyXC17VblKqJCDTo20VpHCbNBv0aNieoH1ogiUPaU
ZfNQsgYQqpdAXTogvgiFfMRP5JoSSRIWewN3SGB2Q1R/zCxboFkrfa5gTE8tLTyp
qyP/mAupyT7pVPqQJQGRb4g3Y+HFL84LpQakM4VqO6w3z1kLimOHhXs03Ll9net/
31DmiGL4YcyB6jGK53eU7w96zierrfcbXGfyD/zvZBGjiIpjE9uRYgl6Vvh5bJOT
YwFKEHVAr4ImBGaUuLkrowBGQ+LMnm2xyXvntiVtJZ5Gnvh4rn+zdVWfCtqyDhdJ
JQwiTbthmQdQiNYQdbUjQJLlj+byg0HU+rsUXMa8/K/XJizYvudkW0A258njUx8w
tOo/hOeTweNW2NKKZRqlVzd6r3NLUzEx2MUJ0GdGGxJjEdsGnDXjYCOpi8ZF+tv/
psLJUmmbHbT+ofkml4vFsXsIzJa3uutV5dFzH1y6e5rcH9Rhkrx0fE6aX321hsoD
ImoVdS6fcjFk57fE6YovzsmhWa3rEJhBVa2dWzqiPG2HR/0VRWEO66I8O8FtTkPr
Dg13wWrKDl1IborsepYuPpEPf7TZvQX/WkoQuYtkmAnmqQA+egvNiQGrpPAO3atR
kjf8eX6E49Yw0mhdiOWH4rMbxwux+HYVBMX8AWjVEpuNGZsmKUte8WC2e9MxUFjV
UwjpQ0wVTk24AgrcQpPPrLavg9+Gsxqd8q1zQzBhcrhbqCoB1zh98NqYwH+Uj7Nk
BtiR0QB245n8K47jdj5rbHiH0wcEfFI6CHmBGjj2Vy8KPUmZhwX2VXfRbENAYZHb
ZumKxxX+g03QiGOG6j1vRqf1Q4syPrYkXC9VLqTc+ovXX1hU06fh5qVc3XHFPmRu
QjdkGulRvb35HQIcL5LP6b2eXS0Njv53ROCGbCJI6BMTRmWAPIJwq5Y4j5rjGEFZ
3Z0MqOHHathgaDO6h751CqOO9VifTz/Fqh2gJbXcnT+uejC9xCRXWfXEkRw/ZXUl
D6thmBpN9fwpTx0jtFPNflfUatP6XFSOQ3tgqsU6KFNqQc2JruTRPMZHQoGvB49/
ZVt7egS04812ITha9EPUFba2UxgDselAH9WOykOHSJrYse+tW0ir62mfMVCQsuYu
JMMX60cCEjy0+9GqGB8zrTOLASulmAyKNA+wGXsfKr8x05xFYilKF9DOg9uxARRn
hM3xI0EzdQjvBMcGWi4VGY6YSdjmv0rrViWxCiIuK2DDkju5gRxOJ3cvgTUc40Gs
azJi//blhYnCOicc6PPEKvwesr1+1r/WYhtHq7SswRRqYRvPaloi+NHs7bMRV/0w
chAtgVdr84jV46lEj2cGxG10n66V7zikyv3R+ko7UMprucHmoz3KE90A0jvXoDIb
OFTBAs0xJ18EEqhgkFBGL+iab81agzFqbyl9sBE7zM2hbpF06GIvus6WBvK2VjA+
suIGa56i3hILoPvrHyICsl21ukxAjD+9tnrYyQxJn25k3dSNcy71oMz9ByIZ9vUz
6Iz6yvPO1VadVYBRbMwgFhO/PlJkj0rQLAzQB4rpaBvuMV5v6aKxQbpCHSd/phMi
pMF4z5g1xybbaQqvO7d6jYx6epGUjjwG6sYdd8TpvjWgmJZHRw5tKlYKlhFTpV/l
jAKS3GOQzLVM205PUlxyfrx46NWLvafnusxHXNTHgc0p0I2vpJEh1ffRGD90n4X7
Z4apMmQCPSn8KA22uFhMPbMjpfhsR2IyySiG7SkIOrKB4JqP7BPL+vaEIIXlYzd3
wo89L7vsuNX2hBtpeRJXo5HFGqL8JCNSFE4LOx677QTT+WwA8Mgo5t/RB0btuKk0
PlmWub0jhbJVHh2x+05FTgLtKh2RmhjpzIk7wzeGo1qzNrowwLiQaUs/gHQRKGYD
zvF2WYoBTkWdquChptwXm9GUoxb7a7eArSZn3KQjEnp/Z6GasBFAp5BaHQbfDqf0
9VoMGYg3KobmdUGwKS+15ThA3+YaI9TQKFCjo+l6fL8CqjWD5r8aIrNV4T8r13SR
+NrepK3zquB/R0yWXVffcMVchnZBldz26IYWcb4Y9iymRc5FihAsqFnbd5ugoWM/
oCSce6gYhwzra65nHUclXAYM42qGlD+M/xb2xE5oSnYbXEsdqgfH4edLM1WW7oVI
0vsY6jvsMrGc6jVIQwCwNxD3zmA3BUzPLcYv96wxCkdO9TKIyrIcPU6b9h1QOuNZ
loWpK9HspIwukyi7BZuYJ9PDPBhxh+59QnGtImgnmD2mtnlsgswJdold7FJaunXz
idgChFrSaul57aiKClVTh6qRPwfl6KBxpA59lDQiPFXa+IMoqwXRMdcf1/OmcWvV
WbpsRbJRLqKkZaOFkScAMuZiXXrMZO+DnnUICRLC5K8gCuu9ShmyNDj0E2WYQnu9
WgwbohOJRapgVNKZX74gwvwE9fOqMlOMW8ElT02PdBqHlM7DP6UpIgU3XvEZpZrg
0x5sBQMzvIvzbIewAWVfdq0nP6Wzu/sdsLeB5J3JXiOZUowVjY8jxJxbyEX+R6AV
RUnfGVYBrn+1ozhVGP2Gh1ZU/nYo2JQ3Ou9vK03Djtq0NAjxccB9GdD0B90qdcj6
SbV0ZIYpJVDMCcfqKEK3Ou0sMlcF7v5Isc1QH5hFE5TFG3yiQ0YiAgxFr57gpPHS
2PMJbNIwcSoeXIRDXqWUou2YOVg+BZu/5csXGrXJ7nKm3tUSth3//maJ6NBPcpvA
2BqjB44u6v88UACpVyIGXpRR+t/ZzgRDuP1do5SXRvl2RMdkRolAiEQ0tA7DUdq2
uZ/8C5ie85yfL26Rfel42s+j7F3vbYzgiwp3cE6ZGfyXE9DOshxEwTOXNCC25Qlu
R5tL+tZiAAIyoWtwg0aICs+qHFhdQiwkKLFhNClyuGnEUIwPO9waI8vWRwOvDwzM
Gb4uPmhvBKlEypC9XeNh1DK23ynKi9uzcfryQjU3NiGVqB1ZYPhsiyEKRk6qKdlH
lS1XWsdlkNZGSssdnev+qvIeaXem/d1CZpwGlLcRfiHjIUCWgdIEW/9Pcdl91Uoz
RNumDiXYvOwx88szsuoHAbXEEirHK7GLW9kaMyCxceQ/IgcPrsTpujqas3u7KsIQ
nYNaiPP0Qo63iHaOo3N4N/ncbOM7h4/29w2kZdll8hd/uWLRwV4VgCxfsbuufkeV
aYjbAigA5/+962lnF5x98NqFpzQ9kneSIWRz5j0SKnACUqbqAxeALzrvehPApsH2
PWoKl0gQQB+TUfH7JEaklVWUHVz5S/rua0HEUUxnpQXHFXXRRZlkXvlJKSD66amv
QunClvk5PAcg7w62QSMSq0Je+t024LvmTz+yjn+/EDUZFcTrhdZ8+aa0gwVx05Gr
UKVKvEhQGUg74Me1hFcFDayzutVLtAKXkyXxPVlk3sBeNu0gd+s0jgj2fVHRg/WD
EAOEUshBWeuxMYgQUOQwjP8xFqo69aOSKlcYD3K7HWei7jpPNKS3NC9W7mgiUGsj
YXn3PVOLjWzpdVLgShOYwJk6KDSMyPq71UmufXR42LqNhx/8Kd0k3HCICtHvGRo+
+reEGaCjcghx3Q/Z4e7Q+kKpsxnXhLU/j3/4HRF+4NZncdreskTzqlTVWijyLLrp
x1hjPCweeJMumPE9b11bzH1xV+kk6YMLCtvRH39D6UUQtaos9FmZcz9bbZNim+N9
Rywg/X9+ZGOMQhYmM9TBVVb8evZCWsDmTmDwqDnWlWEjw96svgvK8qvJ1Tjl88EF
uejtToxyuajS0Zm0xW78Pb9IEr00YOcWQY2VsoSpf5uFHHWOS3j8E5RalTVyCXhU
bysL2XQFSjv5V/rz+qxHBKAWACAamSbJiwSHFeLa2vqA6kAntTVNgSW0ICtKhFTe
fG5Jq9ejUUe3MPnUY7MaiSd9ONkjF9Lvrb1AprZ3qRW47frCiDIeuOwK8bDpWZex
Tu8J+5hTgGoFnka/4E0WXonyxZUas6e87eTMHqhuPycXJu+QuYhe+z3OOS1Qzx2m
huqo+9PM+RAGrsbT0QDqhpz+Op6tewXQcLhhYg7bYjdUag8MGogPvSM85kFZh0HH
0qB2EVIVhUk4nupyM0rmvrPgaBfTIjU1akHlGNBqYqXwIdL8o6X4RboFOgoOnZsg
1gLOItwK8uE54yV0dKx0rznMvRHCPh+mITXU0r6oNnYP/KxT5htWzzr6AShjLNuj
wUDVhagYk8iPfFfN/VmyDj00eD/VFq1bpudBWnbhB26yulmOy8tZGQ4X3h+X0Qrc
ldjimVaL91LBufcDNMQtzXHcrwsyzage7IGhX7TSyNBKDtUUuOwz515VReADiyLx
4umcHYFvBwG869+ha+dDLqes3jJDU0g/T50d5tNdqMyHjpfUcDJrBnIbS9MTQqui
2zLNFaoYlqxgYWQFb1H5V+gGHFbW3X3FhHRoiOj87kJdqaF+x2AHURlTyf6cc/J0
zK9K8LXYekDCl3FngzwHLdDb2VMJhoS8e7Y1jUWU1pXU2gYvAUknpM7Kknf6E3BZ
LmzjH8kOX/OAYQtUle/2/dWcbwCrOTVSavChZiuKecTns2FLLQqboqTMnvwpS6fO
z2WljhpUuBoRg7xmjFhumbOMDnDLG60LKbD/hQWEghsG0GrDuKNxYCxUe8FPkIjw
0OKKVAL89/YX5fZIqnCrEEYdQp6JxGeXYcS9rw5cF0ah0llClXWOIofgomE5lgeB
MiOHAzm25Lb/4nuLRFbqdxPmSt0tk1qE6bbolqmjiJqP7lWWwBX+cTfHFGKl7yvW
IXt4a0vKiUyKdYtL7O+3u0hoTa0nCOIcOKFTR/ab+EexTbLmYeHnw2zFmD+/MDt2
XL/UVpSFTq4bnZ/Q2BrrohwJsezrR1ZxTHe7gxVc2Po7rpruQlkJU0dSVF6g/EY6
KqZ3uWirXQLeTcHQ+Sd7PH0QOf5vpkefS4yS+3/Ci0T+Hv7edDdLgd9ttbJcZmnc
ZYA6vGP2eIrTsuc8KAIHJ4ZcklFZg5ujdaTjW60AAMvYQrIbOaWo70RE5/W/+KHw
IlZjrqgo15TVYiG/vKmBZgpXubqmTLMve12pmCG6cOiR7lPQ/ZHUEEjTy1FDI+Mo
ZgFazZ+JWsEmhmZxW91tnsfiI0JgsFciRs1VBcogOYT7Q/1g1QuXJKYk3HDQsUws
JrSkpfOxo1vZs5QzdLOCUUg9zEMfR8KwkySWD/vbXIsYL41MiPCaWYt0n5J2nQC1
6wmvyPprcMijVZtq+xmpIqv6Cq7hYuW94rU5Wykf4LqtR4RqCWDKSSvjNB+p7xE8
FcPGMOxn0Ty9kGxxzyNCKumIfmZ6Rc5+AKMUbagPoxwnXqhNxZF5Ib++uAfLBtY0
pRhHUshnY0G6AdhURBxjqrXfrsVw3hCLNfgpC+H+JMrNIYQQUytkwJP2rmOi3xzx
u4JLH6cE4Ij7po83DUXMIuBeKdOgp/LEiQHkiPmtGHuEXEtSBXOoeCoMCR8SCcec
qE/StP+8tUkra92MsQV45W8jF6tSUOs7P3cSLzGXIryYZfrzjIv1U1gNlUzA2xCd
wDC1fAQpZr3V1K5py2JEcugkVl7oqxSymfdpYHrTxaJsklOrLyIQnDmaqmoWufYp
iWQ/CsMLVUztddFydhj4JbqRICdpL+Xdi5N0tZMgM/5QMnsiq0kMel7LiSGYgfhz
Jt6JSEecIVujmovLYGkfFPAsBGIMb7AoBeTfIPhbSPThlniByhUVg8XvRMmRLkxb
yOKtc5kGlFYQznhB1FhWedPmBs8a1OI2wr8rGcaPFtrb1HWOhk04B7XBVE0ht10c
2Ry9geG5klNrCLi44x2ozPVi+GkjZ8gD2UKKQTZ9Y0FiM6Pf+aqrkHHesR8NCiNg
qCJs/dtWCsfNZR58GnaDrUijQMIAw5E7o7FY5HnA+VedwWHCNujnjvo8niXLlZik
tcfhM4bm+tQ9u970T6rnsYzXW39drQ1Zx4uTg9U1tylUWh4a4A2URnN2XMtmQc4J
3D8tAUO8sjCDhDNQfekS50nWN2uUFI/vCZZdrxiM7ddJcX4At1fW5PmWzUh77a+5
nuzP++A9M2XF+wmL/7Subj8vpXZTruMs+BT80xBTLD+sG2mCGmdMBEXMuq1PDKFA
zGKxp5Zf4fbAr1PSANJ0yJT8Eir74gdCLxWqZkYPGwGmEB7NPrTpZ1cQjksRaNXT
UYQcXZ4aEN3uywKlx+CAS773k3Fg/SVoornDjCQ/POLqm+H4IK4TSdf2fCvaGxZn
jmBXGIaXWn2Pqp/OwDc0SpQx+NIC/mE7HfXyotjhXAccBPCMv7LSG3kjrwQIsa68
XemyFuZU4I9ea2MPssbBZ6Y/aaD0JnJYOnr4ymygex7jGuZwP16RJ8NwQm84bZgW
xEVOV4Ik1b2RiDMcQhhq6hcXpFqA+m3Zx2olmxMCD98nGCKTansqSk7kei+BThHy
Z9f6QpnsqK49YdERW9lXb3ALtg53NS74KzSEjVU9j8FdXhHO41HzapbmSeCcJy/1
6F9u96VSvebugvcORk/CIio8cXrLsmImc33reLkHmiAUBoUADAMQt/jd6zIVv6cz
QEEHxksV4JoKNGWL9bYFZM7tic3XDgsDyAVaySsxm4cjZs8ySXnRTKTXC+0Cd/YF
gD88852ajNamQaqxqLvcR2Xsp0mf51+SJ3/7Y1z3L/EAKsgzZtrF1sTx1QTm7uMS
DI2wD5TpwTlYIeaiR3cXdSVb3ApO4KW3YHO6y9ddF+aaByUD6ZWkWVOYB8+qa6nT
KCGLyxScuxeHLqhzr6R0mUFdZ+gKfy4Kyt0AWMeS2cE64vzbTnu0SWx07bWOrOnK
LlNmBTwuZ8kNVOJf+lMEszwzLYKpr5cQ1Fcy01zGAsT+I6U6bEd9ul8n7KyYOsJJ
vVctGa1cW+iPgNDKAeGrATfswsPURH85knzaTyTWIpE3WGWTj/+OCXRqhUldM+Rx
fEr/CL8kJ5gKBPjjDs2Fc08fBjPI7W1Ku5+O6ais4MsfVKiC6YI00w6OFQnivNzy
6ewJQ69V6MIpRXQ0J3z+PaKKTYjhKkFFdDXLTv++kv2HxTpkpbicWSLClXtODVuM
EnUsLiDnZjZRwxy+6ShAqCqB+qOazUnc5zxSrKghytDOM4dWhe6Hw7U4qivdzs/9
GI1eQCuJSKWctvjGFYIV/J39xeOn0DGv9fOOKtIPDuBs3Jw257kfOBx7dfs0UAWh
j5aKhWCv1/5Yi2jQo8bNT5jVyypAGyeGdYGmMb6dSED2hNc3PX9f66B33fpH9jdt
8W+WzF09BZHP9q/BRgWF2JVVA7wG0x2/lLQ1UtH8vKHTdN2ft2t8CfIc3HfKpnFo
EC92c1C8jPTklTQWbClqOm5GY3BL2VIAoJUKGdkT7eCtTD7uWzPLK3P/AqxlJr/B
mRY858RSpl+2NsHLwTlP6dMdDT3+J/kF3YUQoLHgrq6civLus0Q8GahAmZmjTxPO
qzwGi5pp32DL3iXt3RDgk04URcw5s58FD8+wiGWJThRchTbw1GEtp9Ly0OCoDD3u
+Jc9+tenCu1/aajihyyvIsOHASaqIJc1scseRLhIG8Wg8R8+kO2FpXJ7sk5+2wTB
XgybcuWsZhuAWmvGFPN4MeT6Yl2ftDrqETghEytahwZ5UJ0OOoPStXVeZwqx8gQ+
Zx0Hw+w+bMDId74nMmXtDasqyapqIuPVYQ5pV82z01wJ8BHHwtYf+QBSsVyPkg0P
pF+IUKDSz/pp/Zkulb5GemdNBZYCSH9v+VoYZ9K1ZN9zns4zWSnMwaFInQp8w8ws
wxP/KvjaNvyNGcsE8j82hws8S7JnHySrbWssRRje7Gtvbd1DoN1204sRApOqtIdv
OmDasHLK054UPepIXJZvF0r/jMVOQQqSoRc9bUJAgWHwK7GczQAutRLDtqT/PHHi
epcdND613kRV447H0JIe8rA56l7JdZbSYpLw+e6VLOr864takySobFH7+qq0+31d
Ti/0bYj3XczyUUr//6/uHUvBBZFWgGTrWQf0Q8uFwiVNQcrAFNJhyvboiYhC8m2E
7wyseeLRGtUKHCBrp7trsA36RsiUfshuq/ygEr9nWNnr5jzvdim4cIaWSKPPXFxJ
rNpJlyaYJkU65DNvRCKehdeAaS8xDFDFkXFg+kbuxshJWbEdr07rjF+Ml6wu40xr
GvMXI7j42+tRKF21VOcsppI8IUfKo8y/RAwHajN5GZjpjpt34jkTTTCu7k05jMzU
lMaHqKO2gcUnXnJP7hElOozN9yrWDIoCUz7LtU9hCdCm3w7CA92fcy5nUmL1jxUB
wZWJd5rq+rjXAnhfn4NJs3+3EFVCSuMsnlt4DHz/pIYAgXYhXW/kZEe1MTgU/TPu
HfPDAarCjzJww9JdNAFN9EJjDgJlenQEI9+ZAZgM1uKx0WzVai+73atsUVfB5QTi
EQi4Y2uOzXlNnFf8SbsQSvWt0wA7VAgwqcQ5gN5PgeUlP2XIiWK9GHpAPC3cKmSx
RO/h/4NCvgGSULj3R0EyVpYVhmnHivAG95EfL+RJBAE2Wk6SFMSKARJjo2AWTZQU
hIb8GchOwFe8+rmLcJELcearWOO8F1DYHg/H2V/6HUGi2/6U90S+Ojj7WhQO9/Kw
h40Mc7j2NWoHU0KPEsT+WYN+ixZAmHbhux9oupNLnNrkfRMQML8KYKukXXz4CDZ7
G5FcUjaRd+NGiJNKjWQA7puZhf4HOzhHzOzUcapAoHkYsk8CjIAPpE98rhjNCvFA
6PDP8ZhuGSXD1myWB8Ck2s/pAnsONe6WQGnVH5kdUrw2jV4kw5gwNy/jIMA3OGLQ
7GM8b+aoU5vrKo0LxkoKOthFEgmWRLiUEZLK+OAlGc6s4fx8gfY7M0tNIYxIPEH8
epvmXEG/F8ECwGtAf7GGqDFG0nbA2RomPUcGUYMCqJkrK8WbIwxszk4FCKcsxIPn
3jjtRHx14+Y0xAEzIMx8TCLFtpI2MfZwOz0gml0BFGqw4oVrkBMeQj0vT3slUVF/
WQSwAzzxRvw2jR5g4J8yBFpFRfssl9DpIwuiGyLZsgfEI6MlEkhqxTgXs/jkc6aI
uWBUTP4oN1pYRIRSz8tXT3MeDFRbUzNxmkCQut+Oi7mylHvCdNYlYvX25G89SyWC
rMKvBVcxt/W5l6baHHLFj9TBd0mAK1q7T5PbIdZYBJbgqpvkirCHfwpnRwhXaqt2
cNOIfT6WKWrRFHbOdo+DO5RfNwd8YxJ1AOivkzhKmaFMR+Ok7JmSyCbC8TCH0b+U
mRn1yUGBQYzfDUq+Y6EyukPkL3LoTd4KnKU/I7Hm7beTfNfQp7F3XBPNNxEvIRQ1
8frBsqVGufGINkBP+GxwekgDfTNJreetF3MTT7RvK7NqLcsd1yship6oQxPAJ0ch
L3qRN3fStwsb5PDq3RXo9CTr994L7+5ERX6eNv6NkeVJT3dmSpLRoVm8FE6uU9vQ
hl/8YHGmVqWE95Uobhg/iLuc4BDijnSJBkzvC0Mg+BdV5s0FsH84I2R0c/AToLc1
pb7rofs2Z6K9vCViIelxB860NfQIOnMvgLE9Ad0eJmTJb3sRZZZ3BaiCNFcOfSSa
qEZc+fPx7MAJwHCveLxoRxdARxUA05JjoPzmnXSL/wSkSd7GeY53+DNIJQZATexR
8Uh4iO0nBkHlQJQ5EnaOQAeU3e3+3h4DwSmdwEDMNPKoqiYzn/FUHpsQPqto0+ae
7MynispTkdErrDRAYdDoz5oyGFtgdfkGu2YZDC+EJkfk2t6dKhv/SqV3K4lWjthU
9elDHA4oGkm/O67JWxIcY1z4TsQatMH85fr5JiNVlY3x2EJZ3RrtQEIhF8VG4DB+
PwdhpkRuvtDkh5HAlBzAe7w9Ap1hBGMgYZPizgn5uHSFV2dTZE2BlAdjHcFjddeg
trf7MtCg8rpalOci+VH4XKJI728iDfOGSyeFGKtC/px9elTJh7xbuHdoDhp/Oyqx
K4TnWH4hqAuMsgtAs3LTBU1hJRzlmCKrI9mac8DTQt0waFrDn+Sx8Thu7sCz9MfE
/w0ZAvpVWr9kkclSsgZhkchuW3ICVgP7pAfT/fErAEQF5XJ4heoNo2Ny54NFRwM/
/sVGxxp1VLXsVsWdYMIG8sItu1PX2pDcr4tDFPbzLGf+f1Isisb47cRrI0b3FWWe
gBhdtyFCAFQ4Et/ZcBxvcUEcN3YOAWy61zcaeWYBtnyK7SppqGIBuQa/Ta/YnTK+
Iqt58pURNqkfd7qqeZhDEDLjrkuRhCsmyFZUdQFvAnjq7Kpg8o5IYxw/cT61dZ19
PJN0TNm7HSNiKlZ53GBEdJ/tq4MNlQDwbNjsar+JCMxEPEwCXO3SQreKRzTvfyJw
dJeIMSwCEiDzaBALFOjeWjcMn8TKDgl1av0KvIEZFwSYzcPiYUnqzUEdbie5nFxs
C6KEQK9X3rDTLGtYTFbqpBuucp3pi0jZ7pU7AsS6fOngK1xK9X7KgH/V+pTeQvbW
/9dhzZemiXoKdfSVKm0VeTsJBFA4ZmJAopIEYkpberyXMrtoAr283DF8H/+SdXJt
9b1//d0XKR7FUjSGJ+OOviwg/RaZXC/UmTQGpFgC5o5I85MHQj/kKVCRHTNg39m9
fnqxoBGMZs5iiAQ/mYKRNbjEaiWpbkPEFWBepgVT554auWBbaDjGx9nd/ROCY6wa
eTREWc+/kXOsCEZ6a6pKcKiXXy14uUT//AjS/0pP2vqgQqBCPouPa+X+gJ+//vyX
kYcKwwIe8pFTqrFTrf7M8lgHsGuscQ+fpY0gKNEfWEw/ZYrnOV7cUEcHa9Oa3y6V
qPWnA80RudqTJ0OVxNJiLYsqvs6xFnVAfhLa7Ygtz2ov8eMKPqZfWUIG/iS66WyR
xRXAB1wZ7G6Sqv4SaUCnZQg2aiVc3LNriru0wpBEIWRwok87otUNsGLFIliHfapl
qp1vcD1eTyS68Cz6cXSglt4rJUCgxX+wypNsaVZAVDGqBEK/lip9BF/zGWrPrvvQ
rj2iBVWJ3gAQbkae5ge1ahve1XFg+8krJ8EOkzcYm34Hqb/W/B0vWnUE9ItftDgz
DxSAmyhob27np+YpWAOJaGa35L9PLVwIP/ygO//JmLfALNxtby3fsQesEH1/coxt
incSmjoHsd8wqh0Gt0ecAphvvhs5CoT53qih3smIOsbrTtKNxBfeOj2LAgrUEJPO
ge7tTv81CBzeWlC/pTMBrfkZuophJOEY+auvqPHYXmUlKAooH9+HsNr+pBFcSk28
n2Nf9DQSzBko/QbfJziwPFpg27NXVf10I9BCHHvRAdYvG75wO9s3BX67t60vZbA6
TJ6XhPmUqPPMenYYmJrxdNepgw5gcuNMGfebKKq4HWqABHklHUd8TvXxaePm0Tqh
aVFPcGes6jC2R/o7zdRwQoQq1fJwrB0JbYH8EwbNNmmQALNZwX2yQ7IRjUnQTgaf
eASCBoKF/Rc+YkJddR9/VmH9OajJTmjNtVmbAQLwOkCgnCILHFeT32VWV0gzBC9C
oRSqAzMmLDWQMXqpLTrUBNzY0qfOK3RsEgvQDySaB8yb/kWPioAv4Ghgjuzx8+Nf
MtnzyAmql3ZRezimk0niEnWltTJy7r1HmPuVF+aZb9XLETP0E5iM1oJdf8doSU5y
MjQ/srLvUZU0ut7Df3r/4gMKU8wVpyV0f1P8OXvqSEKVRvelfZdLmVWjDl9QhdrT
JjcC6b3DtixsH/79LvEhMuTrR5fVNX0o+B+bA1qL7uejWAM9vUUX42t0HgZ+O6f3
VgZzrD15dg+LjDVqyYBEG4p/iFQIyykXYhb8eeQvCz4ZIe6Qkrj8psPoNhqSrSgM
yTOuzGW205p5uKJ+F3yD6eHhakO5BCv+SR4NFXq+akWwp2n7kHBnmPS3yXBKVD0A
EcBg8LpSg1QMiPtMi5xk8IbdPhRUW4+xEhSjOKWbzi6+rV1Se+kpufs8WkzBqWIc
OQJEdRRydGAIrfCwB8a/scqv3Hvp3QCbdSF2vVolEOlhi9sU28e2YqMktdAox7s9
38KLoBr9xXxR3wb8Jo3Fy5EzXbvCBdQOB83rqs+PS3TacLD1svhNUc49OIcWfSUJ
50bdqrQgY1RvTdc0/zVb1Jlc2yKBSL+jgjnmEGuY+kjNdvw4hq6714l909n7lJzP
sWkzB9B71DI/jsfDm6wWjbfDkGEdMwy/buv6yVLCGi+3Fsv7drvpWYyYa1WPs5Q0
Ga3BNuJOYepZpIEvJ34zhaYD1N7TGH7DFXhI18hVcRpFJbLYK6yg3z8OR/avjVVj
+OnS81r38auSbyzE0GluPsPZEBkGoajiG8s70VCl3XwcszwtOIiu9xnksEj5Kszu
ZfW4rxC0xrJcBYmS9m5mHoum/yfPx2Ty4ZBdCx1MlPfQM5BKpA3U46e4q/rNIT2a
hG9IFDMTCaDEhRkKLh2vc78NABlymF72k7D3ArZ6ksV40sHxeoHAuzVCFXcf8GJJ
KOeA6TW/nwSC4SHcwroKCsEPxrt25Q32qZLLWzSo7NkMSap+lspkxGf8OjI137/v
IDE6scZqhe5qgDVR5uKbepRrUb7++dCyWsXzHZ+RpcwBigzjPOY2mlcp81jih07F
3JfjhVNQx7IaBSJp03z2H4hsa+CA3Z+iJ5g+xhQe/DiBdH86OnUuai64yu/V2uZC
1CX/MSnTD3TXiYVv6CvVJqCFbAOCiAilkCR9akwExjIfkuvrH6MzrwWPwZfLOyFY
zvcn/UIY7od74TUb6m8EqnM9Y2v2GbfdKRnBCzyVRP9Kzm3vu/AHwSwkZjOdkYTo
GFtatL5wF/LJbYNp1VKcF77TFC+lZot0HVj1ECf5zt46LQC3WkmjpmYTNq4XNS8t
CrOJp3yLenFddoRr2J4k/DPA7Fubjo0YIjBtVVyyvBWH+HPW4SZ/TEjmA7KTHaIO
Wm2+QPOYRPonSEqbVXWJCMdPp8E2Xan+QCmAeSFwIKx+TdgmHgEKNdy5zvRc0oAx
ndWJT+yC3CeUplJzStk3HaGdLx5owED8VFuEWdETyxq9aD97L5MLMQPg1S6jRFC3
97OD5AWBUTQk+rvU8kSpD+EEO5VqHX8k48kX7+UJw0RqmN9M04ZU3fE1dpD90ovq
zclXurAyHVSIArH7bJXNO0uhnH/yguHPQwJ/C3OuTSw9RLaEPrOUYec0hkFt7EVE
SL7PGh4YBSiZocXeHxzqx+5crVZFX17N6ReD2tfFwZKRytlD6jhgerR8naOBS5/G
g+Y5veVp3tbpGRV4lXxj/GDortx1SkydGxeTGxHZiFeqZWj7WdmJyVzT2u/6uDCA
xtwXAxdPQDxDrHGe+GwTOnqn9I5Nvx51/hB6jonyWisAQpcbceBg9+atMzU93BYE
h+qfFGIlRAJAZHvAejNfg9tOMrxifgZfoPO7YPjSpU4egnmlJa7K/RfOXX5+clar
YAkc2GuzmRItbb40nBCQsDRT3QqyIZzQG5Feaz7dkgHm1/8xPRWYj7DcxtJj1kjO
8lmym/WALwQ2TELG/mjq2UL4pPxzmNJLjFd5OjRxC5CZu1A8pUn6pfix52Jdaksv
TGLY9v1k8R/K5viG9APLyFAK7A5OpKHCvsD9bbwRmklKqZLQPqLOwh+aD+qL9vZc
IMQ18kuDZ/7PxFg3VPN1lk/UC/TFF+dUdrmrM7Hzcsm8FQMUas+E2EcSWbbm3xv0
3ZTgv7JD0gERbp5ga4Kcy7UtNcUJ7AIk3qdPX9zo79K08eGwxstpVL4+j3+Bln3S
09Q2ZBsSthf8BRWrHdqbiwjvM0ATQMWAyuCZHryRYaYpIteJ8OVF2bhIA+wofrhG
Zi07rk3d28Oz1o6x/7Jz9R11twX5TOwxHIGjttrtl435vFxxXeugisspss6rxqdo
u4vAWIDTjP2FYBsNerciUe0H3JEq0b3RLGeJWl7hgjok8WuUoBg9GBXap5sYjrrC
mVTCAnMifd7RzITmPSPjn+Q6YNWR/Uolg/e/ybhcP3cvJr76LG+9GWprRZaDv7Sc
HQgZ55qaCoSs1ask/xfOQ+j2BngF3fQEw1d3WzeogwV7abyOS52DiQQU2dF8LoOT
+y7UvYFDN0cZa83vfL4FMlbKWHXvQv4iz0pcW2F70Pei/J4/1g4lpxcn7ErEFLQQ
Jy4k41VTX9LpXO4PxYFhO/VkAI2uua4mQAAqqgQxameVk0xfJnHSN5//IexZQoam
7BMuwtcJkyt8+IPqbrqKiamBHn267DfEXv4FCB5wP5zUUrPZEnTNYQLeg9jbK8Ug
5sYbvLd5MygofZHCXb5Ajb/kyD1SjC0xmbkjHpIOPe4MSDuJ0EQ1jS21LI9y3g5a
vaAzuPRZ3P65rhbfLH2bGiCW/qdrqDcn2+nzgiRg7ALK6Bf9N0G0knchrBGrs018
3D/ImmAXnngt0oAJk4bzhO+dj8c8wtNci4iE2KNQnzn0qkKkXbnJPnawXRj0dPuy
l54L6jtzFw67mxaZ2mp+wBYq4aksO/OQGFpaNta3DnR1N5jRARJp/HV3lW3g7Prf
hGHyipD78Ji0n2md+iKi35XIyKo53YX05NAx3N/mgnvSh4Z5n/XRym1e7WlSYVMy
VvVePVNVsoZAa3+xIVIh5wluF6ColsFB/lCW0S6KSXHk86yrfE9R7HKo9hqhHUCC
sSzyIp0p/NN6WiDSWeky4zB1AKo/4JO65CJhPTs2GO3PMwcrPvtGvfG2Q8LrsNIX
sXq9dFhUhNoS0KonqGIUJV57l0qNWb36QTVJ8biquNfunadNe4zq/w+QZfgBZMeT
HUt0plMHzkOkRZmwKAmxDgg2lQmnq2EgZC+yxhTWfcduVVxohZ0phMo5RoXhhsba
DEU0hGvv+LhqlLTVYI77DELJhq1WFRWrg7qDz5u2dL2geeiXtOsbK+M9/yDmQbub
uUHdRlM7NmJfjrVPZakk/BOOr5ITIUDCBCXaE04SYdGzZmavsoN8Pw4DIJLfnt0d
2cfP3U8wEJLWwO1UdCXvx9lJWp7Us21j87SN3nU4vgfXhMbJ7R4GOg7AQWemRzUm
EIippuSZe52Adwu2l+uSoH3F0v+X9ewcvZr9pzi02Plq+Sdoxo79p129kAgqTHmM
3yOKcJULMb6BLnOyXn6iu9AzxDlpLq01os5+KA1nwfEciJPvnkQ68JErVVaIyHuP
fePumVs3ytYEz19Q955b1AxJlVfH7NDqh0bzKg7X/8N1/+W3RhNQADssPQePHO25
wf6JxTZdq5UUy0/0wX98OZD7I1nxhyPjeCMPZWKwYpievyuWTjDc1KKqVdsTIvcF
bnPnVaEPM9hNqa0vJwNF/CV5IJ6s/B6l4rlOY/QnKH+miROmsPRQWUtwPYiO7wvk
uNiSVNfiDPxg25d69AxncKqejhilWp4DEXJPXWZJAGFsan3Tf8Vy8ojw1g6oc5gA
1+uoFYcLsVp/0POIxMaza+nqhOsMRegmQBKTbV3VoHrST1i1ljMmAg4e6IKhN2F1
6AR18p26lA3oE8V0GVlMgpBgR95XoWyfKjPnbYpgXtVjeVWJOKUXNuvnfpnMBH+b
8Ge4PUTomaQ/eR2Cu4fs//H7zlBPsjqN/igvigDtcNzCfon2ErLqZchTcdCNZP6i
kAkQ8unRN/5vjvuPxmQk6n4oqHnL7JpVJ45qFW6Xx7TyozkXWrA+IXTcnbRfV3Cp
QSKsrgfj+VjNPCvILoyn9R2ex9NfOknse5P31xSenLCuhGs0AKpJO5s/RJE5DfWZ
SYLxBAratCDIkxQcVc+87WcYxGZPKBWTsDhpknp56VH4Y1JbJmoLxWSYV1+gs3cO
jqO/ylvlnNocrFJB8kLsd69ABLhoa+MhNh3RnhO45H+cqicIgu8prP7yUDIRRO36
N+TmyvJLlkv7HtYVVMu6Ke8o+zGk4jTA155rL1Gqgjjv/A8q4AwUI6mGjuTxcC+U
y/y7XC124ksRarlcHwE4mggHLYX3m30DBdiiopFBfueupAx+OX6UlPYx+weyE8DG
PUnyWBqO5R3Pc+fJutHe1wu48YAqCZXZhdWLj88Qp9QPKea9zTepAJWlMyy0lGhv
1fu/6z/8EhhZTLN9H2a6p/O1DwAmKZ8MpA4ZWD7wwPP/8fTqGZ+kO3iTt1EYYpfU
0palONFITrTE/rNtyAMe3HmpnKSFxA/mgCpAw1PWbiguZ1mHrk+RSs7WhDJCgBip
KFpbNXxj3mVBoDX2JOdfdByq4Lr2j7y0CnbvBNl31H6A1wPHVQS6NLJDMKH3vuQE
edPVlUwNixtlNRpEiOKYCLjSA2X5xC4hpj9LLlPRIEoyyd78dFpcLivdq+3dcuZw
PtkuSb2PmB962Pk7dTbXJVM2ji543qoJH9i07ynML8BamXad1WEmGcCi5iCkI5gA
33fm6DtwyuMEm92h5aMS7zjPs7ab4TV5H/LIffZgZV5Eg6Wd3RV4xKRb7qn52DyG
ApYQuLy5NZkxJG7hlqf1pcQSEGC/kYxtxusG5ncPHDqL13ivaXnqFYjeMv9FSceI
8FA514sJZxbDTBmy/g/6FL4wdkZeM+Dk3yHhTYlVV7Lih+1IT4gyoIzmYLBk/Ru8
uLPoIMhcz0qm0vWceYtaD/r41OeIvutHqT6sc43fQJLVx9FJZXVAtL8BChxC6bVu
cWm2ji7nfJE0TOPhCpuJexAjWas/S+wm8G+iiyVaryvbyPAe0w9q6SW8cSArjBTy
rFoN5uTtYyi8Iff1CX2C38Hlaw231K7fSWDmZfrTSO8R1jjLqBs4ZWpLdt2WINRn
viPxQ4zWaF7q+zVkDoWfxAAeWLidVoX2VDmAswjaBP2QnGqOZr5THnULT0SaAB00
flcAPufhwoKAnOAIaDmtzXZ08v2ZjpmRTUMf9CT6HF1dzj2vTwGtnM3yV4JUpdB8
fv/QQmyhe1d+FCr2gGkk8epCIztq61pSHKn75Revx7qFKPsEB+yBjw0W0tz3+qmj
ku4mZQQX/fUigf20DiNmE4bLSx8Gp1xy//fUdMsnHwIrH5OX4aObe/LQHNlLfH41
dc6iGdnTEPKoum15VUJh9cRia0uDlkqGSOpHHi2pFz2tly9GuC7Sr5JYTfifG7zT
VKfslcwcMNmzSRPuVZnhRU1pz1PemMtQCXSemC3LqHDLUe8JWpm219tSCGyp2gha
TRW8mivdSNwtC9CJXmfUPuxwtmi+/6EeL6/+HTF4ZAKUow37/hoRkhELPYKuiQZc
YbRF0Z4YHooLOu5M3ptgu9Taqqh61eDtByaFzzFgfV98WI9IRRJ8xSSCaOBzjG+P
6NFRuu8UDkcsAJSkGfj50DcU/wfzf1bpHKRADQ3bAYzRqSLOHA83kKYCc9q5n6MY
OvNcX53XjPkevftXq8P67lHpD6QpAtoGCT4R9fZmQxT3CiVpxlaKCF2Uli1WOEp+
ZNdTNZCpqnuBuTjH7xK1sTv/uQ0TcPGTOlSrm/IZWKCObRI80CmcSzw9QEseya6T
9iJt/q8dlKUZILL7UB+tDkV824mqi828o5rDdV72lYZlmS3J/vkMFHBoKVsk97Hv
pBi1Dcnw5rkHekQKfr91c+toExbJIbJz/YwvreZ0EBfL6YdvsmrzogaqHVWjXWf/
JchapfIXz+cjv5ZLIPeU6mVsX/tQJnbmhrlTQbIZC0NpFz/8A3mpERjvGnkQlhNV
2aOMydeBSYJ3uUIcg83zlDNNOZws1nzNlpluCWusaFaJosAnlKUTJvvdxAiBfn4h
NGcq86YoVodx5ErTJooFWsiyOfUZy98zfOUE0k5xyc0oDRUH1pVrC1pxB5ae7tpp
Sdf9Xgp1Xw7pBDQpuNMkgyQThmERUI18mjKxDaTzAk/qFtY8eOCz+CI71S5CjfvP
C3C7CldaB3vpZYkxBsv8wUmtrVCoAk4OOI2q9L8C5FUZb0mlXXxEZXWD2TTbgT6G
+AlzW4bvE/3GGeoyLZRlq4ODdZfO7f4ID3bQe+Tk1wBXVICfEWCdnNyRq28C91z0
ZrM0M/TaTOBvZ1r5jIgZpEqQYGyMhxyBlcYCbjg45NeIHsVQtdLYsF8LG6xRvfGN
3ljyZ3bv9rnRlFPdhEs4lU5LJK6zyOQA3xoPGu7oXs93ZlaPvQuZ8xStKx0Z5U9b
T3Wzk1joanYhG2M14H6JxNfQ+iaAJxc2SLSDC4qB6NlaN7zGo8mMPE5L8RBlzbh9
f8+EQPOM7l8bilQLWH3RA7bAAQfznagZefzCdRR1sVN8tVKnHNozKleAXWMNtLEf
fyy8BxFu+GbrRD2otuZdinuao2FlKPyJVfJI3QhrqjmwqvUT6Q5HUyRzCA1EWCKz
NyPwbutlXCwDbD9O54Mi4EqOsdpsWUgjBXyIXzasv5Nm8Rzlwt1ADDP1XwAIChE3
zkTINNZiTvs+HHLn5Q3JnxJUMT0sU3FFizdtXoREtsIvjYDTq7KMaaIyeIubgzc+
g07zvW+31YB0p/zwGK/6bhTFevpjn30OG9Oa6FjenHZk8wajbrLG5qHvfjguW45y
WdeHeAFtptyPJq5UABIOjhApVEZT2+F+uwjpm812529rLSny1OUZnNd851+k6Ocd
Y2BLyCAuGhaxRPkeizoVUv48uNQmofMZ66qwTWP693/nojZ4uFDPbjwLo5GZk7dd
CsybWmXJXccKKmDvZIYzq1TMSUKEi4SEG/3FMjdHDifFAyASnVgLD8dIdpUcmQPx
prlCca0ztCx9SJhNnq7/KtUmnIX0lPtBu4Xgu0B0WxuCwLMh+c0/DrseRGLFGgGD
BExDP9gaAas5MeUAOyx8u40ukOShB25pw6HW1+SPz8m95B6r/eRONRlsyYa0BqNr
6Tr6yarm6HjTplQKx42ReivUGYcur+XN+epJZb2wsXQpRuwoYe0vhad9tInqB/Hh
WNKnZT/nH1qX1iQaSxa9iQ/PB5dR4Y3GH9/8/rRrJWBJWSb5LlFVhxn5YgWZKWEL
BoVrp2aZhr8qgj8rkYeWaAyW3I9l8laScYcYvII/WJflvFMmkHWVzIkObWVD0xLs
2esN6w/zLiB2XhcypeXMtZRE8UAyU6aWs701QKM73WGM8/sI8vOY3lewQBKj+a/X
CkM9DBEJDl8jS8W3uFnzx8d23LDu8AHH65D9YISBnjgHfJ2ResZsjvl7sC00hguS
WynEfhzwtpH1U8W5XTVw4twu7FeUHywR3kF2+Rj7iPBOX0d68+/jmNgFl5Q0I78z
AKocTQuQY8gL5RxJw9xV9KGnhFFTlN3BZE9PnY/qDmYtG2UkyjA3sAjwlFbFwIkh
iUQycaE3ykKKj27tidvoB4zTexn6y3j7MPgGcBCzHf8O7oApfrDoDR3fkXxctSY0
7sK8HkgCU1HQOh8QVwrYf3gelfYJiAEL+Wr8VuVlCmhmDOppnexjaow4tXiDHtTq
qKp+dqlmgIlF+9jXUP+wTAP3NvEAYJKavLUML/Tp7iRyVt6qWBjKH/K3ywDCo8/Y
5t1ieB6quzbFVUbiyCOJezbDuimdHFkrp0QxqZI3J2rJpE6tmwOVb/3w7FByTzik
C+69sKOz3DKZBX8fJ2O6DrRFdQoL/f7qzCya7v30qQX9lINTUGPnesFFdbiV0RKp
Fg95jyWB7+IfX8irsin1GB4Ui+uz+ecmA5BSr7016sg4knCiRYgYr4yj6ErVm+iw
NVB0y5euDpwpPdzHOynbbRwhyTG6zaBMkznFd3Np4pL4nFiiqKhYLpHnF8Jq0PFH
RsaPHF8CEt69IV37sgRRHT3ZB3+wiVsiLhahi1wr+ApqBJFsa3jAAikFNDC2DAYt
OjOcXAZobDPqSLNZFXJdsuTCWRCw5vp2MKkv6zwkVYpQgx7rcm7u5MQllAojIrL8
xCnRwA2n9GVxe7UKIgLJcuoRuiZXagYEeF7pQb3AsOQXt7QhlNcB8yemYkNRKy97
J3//evmonRvLNzeMHycmoJ8M52aq168CQHmVqf8oH12lqbF2v/TkQS0Inta5j3IC
0hBQYMBvS/Ucj4c6yeHSUBN5VSjtl2zTf09rIOqUzJQLVWDPtyyM5oT37WTgqURB
wmJnLBfi8dG/52XTnOggF2dmgzOG7UfXX9vTefhu0C7Z/rbZSSXkK0pEk4tNerka
7vd/8K+DtsnxFCBItRVac1RZa9X3Ljb6XJW+TGXa9PXEGxpsNFDtlUnX+KVtrnG5
tPUJm4OfBAT+jUeuIN32Y6y7DARoLQa5r2CYOqDK/kmBl8b3YP58BHNfZW9Fbp66
oY89V/qTGu9JRUulLlCBZSf8Ft1VGNMSbha0g98K2/XM02YrcQpTKyFIjxUR9NCV
NMh7eO0IzCwEYYV5itTgfxNcidCseJCSXxly9SgM/izpdbxN7dh3VY4JohksGai3
ucQCFDaWGvV1XSmGuRSc2SO6Qd6tSCDlBkYK28YLAawO8XkMhz7NB6hgwXtiYcog
FCKBGrO5BICsNVCDrT6O8ap1YlSE11SHO1tMDtwbyd4V158o9fRZOP4GREw02hfa
SOWXSgtSgUF+jFGL89fdsrr8paqP9+z5paSPrBLAG9UMzfE2itLeAVaMLaJi1hO5
pu0vWJrWZInMRbxxVUv6DmvGgnGuMdlBwi8vxZorg07kKuncZotCyO67icJOw35z
aIqdIBs/mmwb2GAwlUKlur2rHF2ewHUYyhbzY5FxuXHcdT8dMAdSUZePB0L3bIFD
XXRALtnVzsXg0+WOVhD92oY/faJ0tKnZjVrSc7Nv0tsyDrKGAyu2410zmQ6c/EGi
Qqx0eud9EvnLBkNb2+OSFfiN/0ODT9ZA/WZ8oTeR9ii+WvKBa/1Gzq5M14bOHSex
aAVT32zWctZ6FBWdlkDvXPONuiHfLQZxaKcz315cpaWRRUFNHWU0IEOqeScWBsVw
F7PqZj4lJ1A+H8s+OM6chvNC9pFI4skaObSOSwHysm/JL6CDgrC/0CsMZRxxnk/v
qvNpSVwsbVusgnao7K7ygHq5RHsLC18770/BGsqnogHdRQzpMjI0D3uYQn+2SqH2
jFTYHLRRqFpiMBaams0EoxVgKdamrD0XRcTIbHExHAKbcISZ0bPCnEILRAyUdQZc
t5ggMly6aeBcwmOPT4hfGXkiHiCNDAcqTNEY91KDRBhDdxNlJ/0bw13/3fg9p1i0
fgKcvkO3h0AgqUipRH+JBp4OnA85YpBigaQCyD+eSJGncnmP2zX73ovLi1Qg5bec
WQJeWk1TcEPe3HPqbInPeIo8SNhHmEfSwpqMCrFc4imUzHGN3ON7ZsC+SFiGiZB6
mSjSCBFKLHS+syu7DWCXL6BpjecCwqW6JrZ/bgN1eWNBsH2TT0+Vcurs6hft51ac
8p9aHJPHhfjMZ4HVT8ub0/+ZeFGVlU8myejAsLt4tzyJuGpkLHoruCGIrHue3wgb
wPbY3RYdOt2LiLvXs4JdxWry8Q7z9AAWVdX5SD6RKaLTd70zcYMbo64rA1AhVnKr
3vebkbrsju6luJGPxnzdOA+woQiCs6sQo30/wtW+Aq4lgBSyR8TNy0pPJSnVC+FP
unha1MbHk0+XdKHTQFVE4V+is/EKoxMMXia2SGJ5MqTINrPIj681jo2Qz8H8camL
sM8q7bPGyin8EliIWzj+DgWsJuFpdCZNHrdnOgDAYrekrOKmXXdoNU2ESss/CAIT
zYjS8gAyo3YDQElnROYqfuIkIkR02DigihiDLw9ua4VJ8hxPdn8lUtrMtI7b2jJn
vHTuYjN/Q5HZKfWKuIzQWdxhgJZ1r5FxbHLlfhrZk91LB+1P9KoGMtP4C75yq3C7
p6J6ToIM2hK7Obg5GaIQmsnY5CCqf3s/lCPWGtWwZuU4UFy7BURmZOFcz2UahjI7
XdSW5zqIIFc1RgCsmdFz1YtktbE4BUIKihI6oCt958DzoK/giFQXukKqHt/c2dWI
lS+T/GLnwlMVEySncb0xkgOOTh1W8rbmDwE6TIcDoSv0rA6B3o9abLsqT4watZtP
Q7qIgyOkqSE78PU+LYBHDhJgtFMJSH7B1PcChgnyL6rjpm41r1/rm3G9iMRuow9h
FeIlo/99V0Txya3lkAapqWCOfu8BqINNIzf1krO2vsxWk9zljGp8GI9VcKzz/flg
m4pJSdhcEkmtEeWmizytuY5nCDY00s2pWfm/VbRmFso1EsuayWKv4iTxeeEIT7tO
EMRXrAo11qrQyhJntdZyeo94uT54pBo8JSBdIFOdM4wEodzSA9hEMzmTaVs7qqfx
dqh79a0JZYR5rM8b71kBOfVwCVFIU3CfO7Mx+Ur7VMzzZtGlfS5y97244e5qJ0Pm
p/WjhHTjEIazf97N19bC4imu275J9gMjV239gbX/tyhUczzAqGQDJC5scii/OJWm
YyW8QyPkAmPDk+ZpffrjhsvUCVeWtl0I1enskpgQGB6IhpJWc0O/d2aVHKyIUQhI
XamUrN0QqdNVE7ffe7BfyIjAIS7yYFjEP/+0MS8XRz6QN8NU3CSir5oNqNm/OIaL
VtJkLuacbYkX994TrFDkyJB3furoEZlCxaoMvwj2bT63wPuyEMaGKkFW6zXoJ9oD
VXMt7jMjXy3PgHm7lxaaFr3mC/6z7IzeQCnFz0KwMfieD4ks7y/wPSV8n/H1RHNA
4Up3fHk4OixNudUpMeriEV0eHgSZfWtiHhgg1s7l3SV0d1nrZHOLpzssCgO6JLNs
nbrMRzjQ4CJKBguAEAtvjpI5NpVtR5uUsAtAvQMZwR0XxxP7L40E9ieHH1wObl8o
flt6Go37YKFAb+Ui1zDL29MXMEtsrbysHjYGGg9pVvrzOY0sdQskto7ylvMLpWp3
PMyTpXYbvvuBxuUwN5DoNXuI5fJHtoQH+Tf8GM2QZMgyjtgVGCbzUcjby/Cjyta4
LXajrOIPoTkWbMohWi1M7fZQElwtv+ug7hu4QV5XvpHVjlqLfoyb1olgSZpUrjF5
UCRHMDTWgGtoGJq35o0N0YEwi112HrkphWVrYofMdfU4DMo5jfJfnLOwRrVmSdmk
HCivnRJuXGzogmvVjaaB5ROgJZqgNY4gsbCYDm2JSjp0/lU8Fgla/HvSeITBqFjo
6wJuwDjyksnJ3TuPgSFIDmWeT4IsMlK/yVcVcfu6g9OxRfXKDshj2tHxea19BENK
ttTbzsu+AeB4lkE6tQ+Ymzbu9Z9Y4tWGS23Zq/etVM45gk7ocoNYVQ3muvCgMNt3
6IjEcEczWI0bk9Y19yMSBSu4lttAtQZeahlr/TG/30ILY3aay/alC5WsSAfwq+gX
UF80PKVDUdnvO3N0uOuX/rVhOGZqi3n3uYptelz0jNbt5/iWmsQ1MPxwKA/SepZj
tUEfVSM2lVmZf8aNJuEHDlKeCOkDUeb0POAS/VqMv7Oz8FXk5vtVGsoOxaEvzSN1
rBwouYjS2I6kzGj5YiEBp/XTpWrmflhOVReJUUdFV7xYgCS9b7/+cXvD736TAcZj
h9WP95OiCMVza3JXfVwwaf8Yqe0RChVCeWjVjh5hMRyaxK5MbO8UWEm2yHvyEeGM
ASCqDuayZGMms0MYAKkBD2vq7eLx+RqnDI4lcFrmyQRUkzaldUKJ/v0whZAwDSRb
qLbVaYVErIeT9itPD8ec2mMsoPVXKK2EfYlcmlEzN05wf3XGyoFAII170tH6QGOK
8cp/VvvacbyCRP2I6t7OuE4p80ignqnTZZzxJLVh0TCCSaKyNYPNi0/DiSyDkwSe
13y0EctLs12zpvqhSqfr87f5BMU/7+jUiQW/y3/pzJEhSr4eDaN8FxHFGty90Ene
pZXu/HwPHXVllihHDMhW5f23gIcG2SQZ/kIFNwKyIJJYgdnszKUYyXVLF2PY0a8B
L3Eb65ImL/4t42/bDLJDv8aTHRtb+RYQPy9W4riV60NbFt83A6DnSo3FIqrywrtp
HEyPn95aDgFJ18MYHk42RZJHqJGcvwZac329LCExPSv7z71rHxDDx32wpdf+uweO
WuWXet/kvStRnGzzbRzyjVOLiM2wwOypn0AlonmSksviULsyRGH9W9udvb9dRCHa
qXvbyf0lO04Jiq/MnC7apnlT85njGFK4ern/C1JfrQHwx8J0Pm5c7JhLyjQ2Xytz
IXe1b02m0wuemnZKo3flRMTO6DNbC5Xpp72tB8fZlWuWUj9t2EnZaxVw/yUxdc1o
3+egfsupBTUVzxTRb5HKwLi/mAk4WPnB+6z+tR/X5ZqZ3zUCKug4lvh2JBqSTNrV
s8lbvTkYevqGbPL2qDxA1Hrmg/xEdwhnhmsAicGdYD+cVuaLt/NFJdyo0JbqRXp0
PkvRJCFM6TFzeILh5xeSLn9MLbC2taQVuxVYuZyk8IsX86FROQaQtqbVJbV1RM5+
bB4JERF1KfU1jJdb1NAHGD1x5iE7h4L/V5v3HRuIh2sIJbv97ngoDXd0ciz2t3AF
xnM886M5fyIk6kDISDwrQQx9CLIdS20ld9kj77tESevlb85dw3T5tlwRec/Aoxva
uuTwyZ3uBRh9BnSU8gyMemB8JtQnnsIqe8QVT88w6zu509IiMnxjWwHYmHJo0trd
gMiz6sCmZtn8Ss4SdT2BcMKJ4xfkcsF5n2epAvPpnl3r+hVuZAqmW7SmVYjBMP77
gzItBC0dV1G+nrKh1dTulJseR0G/e6C5Cgidxpp2usMQMJc/sW5dz0Fi6qWqm1Dp
KLyu6uYb5exvzHJdPfXo6Er1Dbt0ToTRIhoBSoVocgvbYcJWdDmji8T1/kr7K17f
DDdJtUQ4e4O1NxyfF1pXxYueQma4PB1L1oxysolLhGBOgEn6hLG0qUmORPykhrND
zvwHIJfKhyLJrJJt9jhGjnwIvSXaWHTZR+elLWF8RpgP8kWjTjW9epfSGU+/iHJe
zfu4LpDlyaYDWCu3bt4GsatoGN+odm5lHm4mn7NGvYzmLVsQ+bGf4seMPcLd9dT8
YKrhRyVyNagDP4kih7ayWGNPLM5yIq4c9GUSMRTSUHkuqGNZLiafStXCDpaK0+c5
mIYDsZ6uBvA7kYxw8pSTNTh7VJO1GdNDEbd+1G3ewQuxWpVtu84ncuFytCCi7ZjX
QSHPGZXnWk5xE7iEADCkdJwVNUjgszXBVw480c+fWCMT7J0TYmj0+Rzrdqc9yJVE
Uf8DKyjXjkzvsRx2GQr29ekz9O1fsGtXf0VvsGqv4BymGeNGBkd9CupCN143UDF2
TUnl1Ma6kwfTkcMHhMXi+b1CpBS1ovj191eVV63OvOXC1dyglSIrydhC1etCik1c
1NV1+hwTa98ymhqai33IWan6Gg2cOURA4tMzA5aEACEQrn7SImwt4dwdZqRX2r4B
JKqm7Ya5CK0Jb8QX9cJqbK59UZk8NYp2oacAuL2JdVI+ZMVoXCkkvu7gxEc2fujj
3wbZa83MPc0LpxNo0KPwu76s0oxrNzX60JvxVW+OUbgnHQI8Gh8zecRU73wHOM+Q
Hep/YkQkm7dU6QBXDOwS3Oi1Pme8wJSjo4hFVMyJFoA+cA7+VbsN9dXzr+7bJe7b
ECxPa+q1wdyzeKRs02/B9WvC1fGa/hz1b0POLyBWlNCtmuQ5yRs6azc8iWbcbA/3
tG0UN7V7Qqlm62VJPnQtxxXkL1azRk0BzWdGsICtXjWUdTQfV+YdVcJ4kJ1DJGfI
V7h6rjKTQUFX67kh7J37iGCv/++el2YxOnoHIimNtsB3wL0F/2DOrfGqMWapnCOp
R7drST31+UA/reY9V++AU3KdiQWDjnzZFJZIm1r87gasXxySJ8emF0Y9yHi3Z+aa
TqBhi+xyCr4q69ktpZX9YFnAd8ukIOk/84OjJre1ian9oMV00lwmSQsTh/Yw/hX5
NS1B4WiDXKGtsK3seZaQubbyUdJitwssHQ05EEm9MroNt2jLdlaA9g12zv8gPQ/w
1D0d9mqNZdNp8LXhkciWAno8gcvTYOZ2vd97l5lVOUdeoPfJPp6YgxMdoWYJvoIM
sqUdaFHk9qwmFyctOnmQTj5AD9+8H7kmegjm+rt1fSQPlRwPWwSXpe/hIEGHOHWQ
nQNkjlVS9LOposdn3FoC2DZ9jsK4j4GKX7GnVfstakZ1AgrqI/snX4chikjL1LL8
H9+mpy9FoVwPpZnX4WbNQ7OWfs+OOC/KBu0TvT8ca9rMPVV1JKTMLJVD2p7MLwot
uEEXJ8zT9rPVE6hEjMhpf1R7NhYuY4lOQYTzUf1mSr6edzhTN0Bxy0hw0jZ1xHv/
Uhi2y8dU1vdvEGSsHUt25BNpmDqfQOI/X9N8wE0+dgdtk0v8eVHLyYewakkGhe4E
NXjC8enL++1g5ztOXMiicEKEPUcPJZj+8fjWFfavKnobJGnJgAto4/qINXxITaiN
PdBxl4342jRpJqRvTVi/UqPn6YUR8sV79c2fHJadbmn3QSLfqn+JHnrriiQPW3Bs
M1990JGDaqt+dfAU0s+gHH7RM37g+lG+AID0j7K4Mb6kYFqK7Tqc98gN0Hysrw+W
YbeEfV43Th+AcZ8dOJF69TzMLmbRlNqFkAFsaUfxR9zQ3iqStrMICwRYGdLW5O5I
QUtkFFO9Pyyq+mvLFsa7fQcOYevRL01deoYjWF2H8vxJ+RHjB1rYUQNFY17qJJBX
hChiZtM0ONiP6iLTCBBy/J39F2VnPVy71kiu0I7tWwYS6wVXQUW0V+gEjUXfvoio
XidKAbQB7slOwGrBwb1eRv0o+O9pMVxhJ3Uy0KR/OWvh/kGSywGJnezwHG1e0NY5
Y1w8TGZWvzVKjmd3TtwN+vkfdtgdwwDETQjVURU5G7jSarsj/atCef5Izdbhrt3G
QYwUw4oMNcsvCwLhLzz2nfUQ67Ik/VNpaoP0a1+hmuhlpXWWRUWVaQQ1/EO6/FF4
OKLm/kyiEaUk+iFDOzrHPrp+85XYh7tCiXqbU6ojUOYMmx18lxyElv+LDwAvEiEu
ZGsH/zopN4ChrkoZg1haDBaX3k4vnH1az6+K1IDVULkybnkN5CIb1OzYWt73x2VI
SkQe0MWFE/YEVJbqCSpLZ/TBa83XVHJhUwgutlyJPjJjp9n6GUsp450721drouSN
XN2JAvJGk6PbsPq6xx/7tpbokPX3LVJHylARzDJSIZ6b09bZyn86f7o3H/AYcabp
n4pOev/Ln/5wR4uuhr/HrggV/Xt2DAn8WrH5LY9Oaws2x/NhHPxYchyaAbbBELjq
xlUVzQP5D91Gu8NspTtiFV4iol1kC/HQlZvbPoN7fKD0ckg32Jf0WvhgG3vs9z7H
SNqeB63zEnG1FBRJBVOMOk7C21Zi0kNMVnQRVsoAUiDrndd6SVQiLN0pKnc4KjR9
wPeORIzYBe0hMSvKL3gP/uVSHZrWKa3Wg1RBYbSQaRGtxdR0Kc9blHtXKmR4BTbt
YAy1UiJ1EYBkYgnmQdhg6GCZsIW1InJfogb8G1SiM3hkbbBXGa8oyOKFdV5I7auE
y67PCjqeFMEawGuDn7PLkuJ7C9lhJpxjVT2HKxlDAFCvyACP0c6x8cVaHzsd+13E
S+TdOMRRBkjS94LhkG14L918uPCk9UHtgKYqZpSfziyoz8+zGoCafp3yG2tKoao2
w3xBaFxmor2MMDFIOqoyDSbFcROrFlXg/xfwEADNkXiJdfnGePKoDmMWQzJ0EFq9
84mNF2TkEd6HrDv5WFpHqcVin1x2qDnx/QgOLo1wyNj3HMVVal6SnvfSeX+0oNAm
sYlv2hPVB6W2PHNGSWnnoPnwA6THxBhqW+t19Gyrw5cn1mPXrCiW5hOtK63sBso/
2jDUxXwAfzGpG3UM/SpQ/HZX5deoiAvLjvPs6DO4vzRFEl+pm5lFYmJRial5KANb
/L+/D1tIDQ3lcsoSGZrZcx40g++FLxnkVCoAd+27dsdly/kDtwLHkbuQpR8rxckt
g6nKFDCX4qPul+Zet+xLBLzABcaLqvIaL9Xs5YTCY8kSAERzFsbE+OOm478ylvPp
IkR9GYpaJrsfKmlGiXcIpSmE/Lk7VrUDRb9Haa3JoRJwtPM+6KEAULDwvNY2dOYg
o6Ihia1CZsjc3yzpX9CyGfjTeoItOSLuAwAnlj5eDYUWIEtjBN0l7TkUp3aZYOws
knTKWfbSNaYcfNj+XcWHxiW6Cs4NORXllgFy81hfRrJKdOK3rq7Xs4MCZkKPWhkQ
2zBo0rT7+JB7iD1u4JOUMe6ujCD7bTfu/8Ul3Z511sLjnE1ef8DaB+p+DjntyWaA
O7rmAOl+hk1iafHMtsypCc/SI43Tjm7UIqfIOcqVy8Qt77ojqebR6aNmECQlgJvN
oIEezvc2EmpkxOWoU5zlKlxyXoaGPsDAwmetdVEz/jvJHhyZKQDBg1+CnsO12Xkp
sV5dVSug/s1WQy0rmjrH4gshSse/6fdpB2PdYmbqUqI4aNKnC8On9JkmODkSpdix
3Mz4CGI4/5eQtQXWdCt1C610hWDB6je7DX0RCDbz44r5zI98mT5r+g2uGioibBu9
qKc8hqT71kqpmhaoi+9TocmcKCt7BHlFdYp7aGd9qLrIrC7EoO/bFtXHNERhrFPC
4ZvRE7lCBKaDnvWQXYw+NAIjaPdABUIEdHfN0AJ0Uu3HpFhP1BQ3gTg9VtVd2XRJ
EtoD3BPe3UjfhWWoTwbqLuDYL80PwTWBxepG8rLyXnXlCPpPLgsAMXH8ibyddoZe
fWqLefOyeD/EBXhJNExGiEgQcqv7QoetQP059v7BSeqqBXSVzLc3hUXhmT84zXuT
n7r4ZapyYu3kGaPHETklFgrg+UpzcqPeFTfvMLH9AWRNPxvsOxe+qeCxgkKlFud2
R+SFcO4sZQJCPQYDC026QPXj2/MAoFbVsdGGiulRVRGtzMqcBO1Y0YLlPldB7w/h
Sn1nKaenyppulcY9CW183eyimUPPoieiPG3aJXy+LvmleRWC77pgXyCXbcl1SPsD
wWEHGPM7cP9mh3CM1wbdpLNKAQBCVMlz3kHfiKz5NnlzoHt7eVPGS/dlKUtraaO3
meFXGgCtKQLnRNaRscSrBaKuEwJfaPaJ1KBUneRYORjtjplYqd6D+FNnP/LXl4fl
Ouz6VNDxWRzHA+DmaLfCOf39yoICVvFEJp1yH8EUs5U/JYqLzzYqCYo11nbYckMs
QATbc85lFzumNoVbu04H8ZfSqbjzpBjhD15Gdr0hSpN1uatWrefcZqcpMUup4MJl
/QmD1ZxYJOeTXSjAQJjSDJuO+PwDmrnoItj1KfUDNFQcfoBH8SYl/rst55LFM7JW
VQXIMclLh6eZr1IcH9nvfRwtLgGurG4HyO3WgzEHDsW3vDTEY9diBrkFurjyipLq
gCR7o5osewr+hkyxCLMbOciTBBdv19jJe24BFUFkBK02b+3W8sgS1ncmvf5VIwF3
dvfrzkeVRbyvm0/2gIvneRq7oNDyUnFzHrol8qa2j6Q5PBI0/eM9qfI2OtUS2aQ9
idPJTC69jgQUNe3PrBH4sJZWEn/e1+7EB7fWUIVnpUi2u8nPXWq2rEXbhHQe0suM
ONyc3+sGrcyrYUkOdQ46coHGXZgWf1i1OVsyRo3wdDcRZkiDGPf9lgdYd2wFlDQE
bsjelTerxJDKZGe64hi54UQm7NNiB9Ku0O+hQt4SzIsphXkPlr9WWFkyUJ/pUT6I
HvGtogTeIx1tqFErDCQHZD91Sh3wM/nff/7OGTlWmgRpv4VgPGIUhDn6ngFBW+qH
x5D8G+iwzHpp1k6KdNYN8McG4uUh4flLDRlXxLqCZwxcjLmv8+FjKbi6wDX/B/hL
lVLVep2dTpQlH3MOpkrNU9NQA61BeVd8KuZx/Vr+Dz1rFYZ/byw0jvRiwRbyXemU
NIDYZESR/nPYUs2enbZNeZJ5kKc544/Rnosxt0wnsYzvI6zCEsGjoMcs2/N2fpd2
BbrGFcWAyjcnS+TFjJ+fx6aaVAhZSyeWpxG7mxAd0+kaOWjMQM4OPeM5ikdYTdh4
GdWcnBjD7zqT5sECJWcO8CmCx8kujotbe61NraeFBGl/u5sNo2Yb2tyD6DCrygtl
RHrtwiVgqrWBLu2TR31YIp2+ByFxDWqYbYFqarWEeZxFlPIkShuMJ9cV+qZBJx3y
2lyO+dNraYarXaRecJQMg9982JlhCS3h23S0T9ze/LqABEOPQiEdRhzA3YzEkUls
qkNFBHMP0TiedmLGUkp4mbZkEOaYrChdK7HccosC0VhKO8EAS680YRC81aPQwoCY
PyUCkTCXJzKLlYyWlJ9zPeNlCZeWOZPJdNz4thLOvsZdsC0ZZInczKAyG9whEGQO
L2+d8gwggMmwdWjkpyB7LQQLKYpNWIhqYsCJ8opD5vkwBqhDJ8j1EqEgSpeICoir
QBehHwvip850qx36xso+KJ/SbRCO420qKKQmuflrMcTuMzsmVydOK4rPkd8nZrdG
Z/5q/q6E3+Cwq4eIhKSmomroRDLTKDhwpdPO+RdOALC1uzGqyXSL3IapshaTm3Df
39VQC+5SgRJdj1pRE0dSzuqX/hToqsd8j9oI1wmQUX5wsc0ogIrdwBhrwOpJqRb1
eQ1IDAxgksc0IYjFbIlOFXcp3XZarbqqpBd9zwNTsZYFrw8mqrjHgfn9AMnNWqLY
vT4+KfWh1mnr3pTk5CLfFDfhRbZwycIm40R5NYvwYVITjJL402BEAjq9qmWcs1f4
xQ4MiF9tmEixr0Yd/7xyvL5LTwutf0Dn6RCYfFFIZ6S5Nnsmpkdm32QOJNx6nH1s
jc6TkZcQ39cIVAOBfdJaOLMQ01hhpCaEe8TayuoTMwM4CCFHl+OGuQci/UcotizZ
bs5jNG8MAKZBfXDBhcj+5wBflfrO6jvJT7ye7lCofQqTbNVf9CCnmT5pTWko4Qz2
kf623HqgzSLTqoX4e4GO56iWEQEoFT0slCCumWZ+G/nXmJlttQi+4tyWhS1dbyhr
zMOqXGX6hUJXQrsasDrrzBl+fDr9M6wIRLqOC8DvuJQlLltr9/D8rWrFGJiJQtpY
r64PfRDlEhp7B2g6fD98+mgcFpv3n2K2olrJfmRRgeQ/fnVY2AbrLvuH3JTpMPzO
sc5bxfXCC9RWlURdvsTOdw+DQvDRPXcQz6DCaqnhIaUfZMin6jffBjNeZ8cy+E1o
os8djwX88wmpeBXJ5QeL6Q9UuSrnBrvD9aHeZT499/pKXUL3BwslHEqHgoNc/FjS
YCezYgLMWwpzS69AgKwhqFCYkS+N4p+FOusdnDq+GSZ7cJdeGROhVXW9Jm/5Obou
eEIoJrCZ26EDnw38AlZf6881Hqj6nt2c4eci0jnTuloeF9H47L/kB1tG/MGLBh2w
5E3L+aC4zhG3xKy+LYgj8srhylfSCElSK3o/TIyCOTI0smSxyu0m21aPid1HhtD0
UsHK012SYycgnKGi8VITwjVwQ1xScCdd5TFRrlLySwcfhUq/l+UrK2Cpmdsbxgml
N6NcFchpdKaJl/aq27qaYsPSkkrepTK8MarAT5fKKsEOFheuJF+AUAT8+jLRlE1o
zoT+vPLAJ6nNf0R8kqXN7qZzBGVA4uDrl1yi4tTx5c4zeTQVtRQdRp3wr8Qfj9cK
CmEsNQk+KyZpN55hYoaVWH9ij9TnGusqoRX4qJGDfPaz42FMLKeQwV92EgkJJQVB
822us7vDHVpABeUgOIOmQU+Z2Ra+Py+Cjr4ju57JjSnXSK40ef/NFvEC7Zmh3aMc
T3mCty7NFAUNHOlvmmnK+ZKB3GKQE5I20VRxAxM/F2z1yZlumP5N3xdnk7xO+Yy8
+ETaszbxnRWyXXs6oibabu0mX36Kk4GhdtHGYTwes33eqNtWjChWAk+jIGoHp8Ho
Q9AgRr3ENoU5DZ4lyZMmkEo0SIVmeC+N9HzvgtWP9M0W9uYc5IvuINsZJncOcqPQ
2k/DwN46QrQYEXnW7Ejv7m+w8Osytj2szM6LjKcL3anbQ5Zjk+OKO+LANMsG76Iq
Ib+yCdyraTEZyR1DAdEWiqYlfY5D+DO3+vYh8m5JSs8H3gUFHMH9TBxDjBSl6AFa
XCLOXGMzWfbgy4OZmp4ccFC7XW2DzIrx2dd3l6oJwIIh6E3BNKAmAjibeGlWiHwy
6jHQXE2kz3rime4CnDuOATETHl52WgdDkUQTpOlhA1Z0NdX6sVNLRvI8odrr2Uf5
0ANOjL7MUeweIIg+I+JLlIJl+aL9kpyVSx2UeNDAfi1FbwgWl2vTF+pLA/Ig9tFt
PkxtGS/0mX7IX+49qe2PAN4HipDxrC9SPqBDDudK6kkAX4dpoHdmYNfljP09cCkY
l5qZj53JOhKf+NKwphqf0HK946r+TFBFw6kCVNoUW67MXJL3nN1uUEnieLV5j8Ux
UzXKIBthQAX7K8HZ6xdgAoajN19LPL8/IRsbhyuIeYcTAlF1iguraUE+5Y0aXJqE
yHSCLsYU2YSUoVKyg3ZKmM/k+txo+rGQjOdb5/RW9h7mlzK3CXL45XBt/pElhy2g
400KwS98eNMp7tZkYl0H1dcA5g/2ohrmHBA7342vfaqXE1kXJC1INvtQyIJwRT4B
BUsC7izqSIUlNyO+J0qJLFEtodsi3GWN9HICJWGBKF9ZgqqUcFd7eJASeiT451C9
lsN8z0njI2ATpc1/oqqZJD/QNbyqMbjCzhTfu4PuP+Iue7wUiMD1EAbHiVSjvXIo
mGgnlNbD08NUsbTbLStRYDCOm1BmkdMM6ahe+giRfbmfmGQGtDeVVRvqCSGXCdFb
vdFCy3bge6EagYJSKFFr7dG7Z+iSivFRm/q7c28ihxarE8YO5uMsf1CIVM/bV3BX
2LD5RVZV2zENiJ+3iZGBhuXATOSZA+pZ9hKwXpzpOhPe8Gor1xZSR4LVYJ4fSe7v
Cfrowuvm7ibRtB92iqnXh/bUWU0VgIiPcFnV5D34X8izwhMKx2nfFnopglb+Yw3S
suPLY48/RMijSLhc+MixWCas0AUF7Q9jU0/h5xj68hXtaI8g0v+7LW8t9+Bxt3Ay
KovC56PxaX9z2J/n3MdY7vM4S8ZSIRyvMc3y5MQ5/ISYXthV/HrLlKP4kPyBBOp/
qbxx8DpZ36i1icRe78SVyNBPRL5tX3d5s9iZo85ojn/s6+d1VuHkOFnyFmkG2qdt
Zrvl5cKTYfJEUDptpYwM6sZMfZPOJib+UFF3LT6mG1wwjRy9hVZK+OIPX25SPpyh
ILAj8SiuOxhJuc0GHevBbhBG8db1TcDG31WPMeS0J3hNzD4TcQvHFKRggTgmGXyr
MKNzC/5VfB8ExreLtlzlGnNQL/PrU5e2UUi1x4UeQ7MaB0udtKOTlCCqYSUkhYSb
UoksRZw009gruxR6f9ZDrVdo55udSk8BF5+4iq+oNoQnhmBkDqPHiJF2R8+bmkWu
7FaCHfkKgW0jQSm9NSeQBxGNFgaW4iq43WvCB6SJwnV9Ymca8u5GfouwFnfMwilz
j4bl12uSEZWODW/RmUivCV2eLyE8wEfVNhB2R9cgTbCjT9IvRS7FfCCBzHWTMP/P
4Gdo+8zU6P0pL2B87yPnJLIVAPi12JtHEQjsROss+X42cBF5/jMQL+o0n3YJ4te6
QsLPeAy510BlSvPGCe46kH7sQyJ7ZALt6b1wAdf4nPZ6Ywo2znAbuMRRqFeK48xt
Lq35kmtIw/GIO3b028NfLt3WxVXvU9bRWL6Wd0uPOR/bGgv2yi2WWyfjoLalgf5W
xJIkhjx5pEk+lAKVXE80pC7GRW7CH9lOV6m5xp1XWAYOJRC8bqPsTOhu+sNtDWdZ
mDuuGVmrl+cEsYSVHzmaXgYOH2Kb9RzgYFR38BqMHpOUVTV17SmlabiechbivbDl
0pUXiBs2qbfcpjzDss780Ql2vTmw7mBJ6qws040hCtk9gqe5fReI5JeAELnnA6LJ
fKgQS/ReXg3eC/rNGU94v1LX70yeTvgHHeUJJJrJztiChvl1tcZnqFV5IHuS9OAI
AhRNEra0FlBIYdTXOL0JEWjVdNff6sl3JsRWWws6a2/FHL6b5j/2q9DFx+wzEEB/
Hy9fZMEK/hOiHFCKPhsbIMnTjhd0YSeO/3DYVFSQ7voYEWN7u90YpGQOcITsaAOA
Cob5Qzve25XEl8ebcwrkKcyTc61fUyd9MZz6zXKVLzVtCNOvKdCZAU1q4iz5hjK8
YbCecFjDywYC7OTvGFdix0iyVB/kl8TsbSn2Jg78FwjhFpTq/N37FJs24vybmhoA
M2AYWmGzR5sXZRX7jNxIiF7R3cflggHzgSHpN509IFnEQ37TCDB04w1VTRHUQUKB
CNvPwobexPH3utv0HswkUpBk7T4k7SVQMxMG6+ElPNctmhZERr5WeHmevAbrD5Cy
6cSNMQVYz+sAunGgVetTlQNOCVJzksAffHZXXFx+zpfVy3LlcXfkwwMDGlEkmLxQ
Aa2KikEEFLJIvAhRu1ooS5n3RzspKLutTAa7rabgG0x/mLOMbcTlriRz/Q2xRNwj
1egVPi8P9M7cWiAGRfBj3ICqBUby4hy8HJr3aRHqmHbsyP1x33DMNJrK5rx3+/bG
l8gKfW9+k3/KFi/WzJDrDim3LpcpcpA2P2+t1n0KjgRZJVPfyjtgm+d7E7SuIYrO
oA5D0aquqjvGQWWGyvstavzhRKhmRGeapHkepQ64B+okoSwdNJFCUSpyjYBf2EYg
pP1LlpSImvNQdBswQCv2UV5KnQu8D7n2eUeTS0Y12EFP32q6EEjJzHlAbNCopF8c
UxGu5jP8+p9D9fhxm2QzYmwL6HbhDYal/A20V4X0qOTpLO9i5NAiX4785SRTsB+6
fu8uwOU7tw+uEq1AvnnnIqNyI9ls92zZpVckWVcEq4VCOISTqWGmXzQsud34wTel
IOWvsVY/60qYbMTFvjFGrXwCzSp7mKybWWnmC5pTjyclVb4lNjHTVOn2kGZdMcDP
tV5Prg/Zh7Tb10hg0+J0Gn4Sedon0edYarfyCiYz/u3u2WjT6LITE4fYzaA2Mw+P
/QxZ+xMFkgAZx+OrCKH9xXf8kzz1ldp7fTn37oIxxubfjRkjH6Ds6HLGHfMN7t28
IfBrueptOPdk08hX0Nk98b/5QLJj0uaBNH5VV37JmjgEmmphVqkh4Hh7VdywRLMa
8hJc7hXZf2M3J3n/PM1Q0hCmZl/v/63sfUD9zTzO4rtcdT0U0+NordGGGNWDNi0U
W3FxZktGxhCZpDEjy5F0XFt1wNGbRT8WKySDcmoxHVU5frxRCMVmg+x3jnQ0Ip7M
qFsh6nTr02XqyNZ6zPQUrDKzXMa2Qp4kb34DMZ6bc5gR23+gn9EphMdn90XviZdr
OK9SuGke6iOE0Yt4/Hn1hG1MAsEX9y+qeIsTe1NsmWppecl4VDEcgbmveUYrvDWD
pkpb4t3u0DdEz3AdB1X1qwk57hxHohptL9rLkBLeHC/0oV3M8PilttRY2WQxV2nZ
fxidEbzxgpgMir6UJy7SV6VrutP+4x04TWZ6aE70E3742vFXqbYvduw6DD6PGzVH
Zcpgz38Hv/OxTKJIPFTfkCbfzYgtE+KZz1orN+oiA9Tb+z7Rg5SqrmymCXQhSn8g
RqhydjlVvRFpC0yfEYJNDp61zfobAPQec9PhdmWq7K9TR3TMe5np+OzPVH7ZU1ox
E5FDHnIzqKhJ8QdjUsbxegWAsMXbakHje3IIW9MKpBmybU4+GCwHiYBOy0HiNSMs
NE6aw6q/eBla0srVobfxwHnEoEc78YtKtU9lFi/U0aKVHfp4nriEIqL4Ts0deZ4K
djEtQ/zDGdFDV/TktuwZEMqRc8BVlUyLqyhYZX43VLCWvAMxB/qlC42hUdciqy4t
nXvyhxk5iglAy425K7/QhkUVz+mxVHV7K46e8qyqH51Orv+BMqhZDITIkygdfziM
A4jFAU9FC4rErcU5q02eo6XC0VWnavBQescF1Af8ZMasL1ZTaZ7i9Kfp3LSaekhM
0/dEftEEVOnRAgHRfl4VeW59zrBEKeCKlZrNTxpHVhksrBSfQKUrTowowauI+gBF
lGYmdmWtIhRde2rJxqXcLvdOpelzS6rqfMApmCjYfeqv5iKJjR/Uer70EZkBYj3D
xbAHJlARgN3He6eesSnjz4l3zbbFa/xQ6l9f0dcB/hO1PqwKSXIa5yFkR7QAgRqW
HV39G24MoXnwcjiqk/HTrCNsNxaL9kke/o0QKNOATl3TX1PrgURDZC/xtRDmu9/A
0CIzYIohAfZUJtPvGUZv0GNnGH98nTrH5xO6OsFFSJt8Xgoa/J/AmpEmhXYXFiZg
IDRY6EIjjqomvtM39X4N9TuBr/Rqkx+GtqTRmOrUzWRgB/3mwMpWgkMdRnK6DaNr
qkc3pBrIEUGUeGPgKozeLa1VzpnSpYmK4p4/6H9BMr3ldgyN/dY91LkNYrblD8/V
KhbpHBh1LMcl7pN3JPFGX9PXKxhKGn6POkDlbkyFY5RP8Hwyxps+vyGaO+ASLEmp
w5Ep+0CKef4x0IR1Yxp34RleNBLsn/puSITrCcC76A9FfRjcpI4o41oSTJBrUsWL
fJ04mDgHL6VQIUh743nWbpt4PxyfDmWPGTQKw3FLw9vgjvFHzWcTTptjy4Ww4AMv
JwAoufNyuT/YH82RFvoLgLlAlqZYTJKC0UvH7ZRNgzE9KjIZbjkj4hZVK3AiKzDe
wR8fmmk0JoKgD3LiYZAu8+VBJoWMJswaUeUHdPdxzp0ZJbJ5MlplqAYMDUA5mqML
/2+hy34Gqss4wSDhU2hGYEUVkXdgHa2K8oVbPv1fDCudydyywzITrnhh5Kgf8cED
rl8n3bi9gb6kl4RGl4ye4u2zzLTPgisHkDBSsZM4UqJFxdMrQhK9cW08PBS3GOVI
o3FdbHL4f+JwLy11NAqWU5bj44uZ+/rmYhO/ljW5AtjLz//+oek+vrqBisZ+yXGU
bf/lL//JiWvLOsIptMu8zx8wCMtPOwTV/FWq2c5HjMUU8Jz/u8QDlhVjrYa7EfdK
1IYAo0eTmP+UbASZIC6bbOm4/MxqHMCtkBIjUNm9XjfRrmFpqdEUrwEUIosqBvBv
sNW4UIBrjTOaTd2pLCQ9ol/EkX2XlgaUAY6D1AFC83deqnq/bSkXiqBsqqTINvkw
Ic/lS6Qz0KwQYALhxDaBLgqnoNpdr5hZfkUmz2QW/9ncv9POwwekTUDEor5uQnWn
++4ZGrNwKb2C1ybViMLA5RUNvYuH9HzEJUzJws6FtTPtu0zTynkwS7fFoHUSsrNA
ZVOtlqLwcF/IOkU4VEG4IRR0tSxduvoibQnCcRnTWsL8SBfEoKWPExI4hklpfu8b
kIg6mDyrP5gAjv3e/vQhGyF9v5rk7jaa3E/0JdFzFGTcmRlzvtpf96M1aEvVEenM
mbdZk2FZeaHnWgJ7SGsJ8v7Ld4samNqOMMSVM12Xyb8BVi//qar5fpk62Q0tfU3a
GGk89DMr9HeRxz99DAU6KZ05ChP66OuLTa07KK9YJ+IeZNsyrUQHxpsVTOZTYn5G
/HR0hF4quf2GABAeBj7QxrAB5pk4YBoGdAQ6btiemCdirPtjhUoOqYtaO/cZrk3G
Y0Gw+Ut8dSas2JORnHwIDelk5zkbOqLbFUwgrCNSTqS0Fup9C2Ht5Hfh7zDWVvQC
2e/JlxFzwmyk9RvxSmrYS/5/S9x8zlnFEi2DaB9yBlygRdF/FDSNFv+NGgLVRQBr
hiVTzK94c2bXKFPgYFb7vrrDIk2hQszFm3gfeEM99PQxehE8kUZWQOycS/3CkKES
Q5E0CqgqsJCiIqFklp8v83WoERSeJklBD2rThgmqXxPi4399qrrBiVhCCSXllgf0
fM8o2ccUgujlYjKOucWbjBfxYjJhrUpA3QaSNMzZqV/vluBXC+o3Ce7pk+5RMLsd
5LVtxo8jrUc/slSqyOAwjyD1x8YLWE5uTai534QsfuX2PlVejCGM0E2Yxd3WXYKH
kxZF1tO948aUC+BCWAqHRSleO7pGBhJFQ3Ed2eIlmUKBvcHbOAHdWQHGxBHUYsPZ
tuXukBexp69dWtmGSKttPe5bXbAAREhhB/S16fNt8OiaiLRwf/4NSb4PGPY78GoS
zgiUcIPuVmNMWSS0fbSlxuQgoqiwvUITkeOcXRS+PY1PcPzub4CpQM7Egz6fl6Se
F5OiwPmzH3JtVcvmSze8+Yo954K5Bu37TVxmkju/A15wyMbyhD4phYp7A60j/4UQ
fyoyTIP+7m9QquvUvpTcNHlTZ+VPaEc24MO8tkuugZNqKISIF6VShk8fPM/IxkuW
R3iczxNjT0XJWkb0HtPQxslJvheUI4fJZZnGxZ4Sn3UXOofz10UKyVRQxFDnD7EB
x9zJpzeiQd6j1dsarcitQnniYg0XRl5O1CyTDGYgIrDd1hOniMUfoLsXqJ02QcJJ
iB4T5ZxjJLCTgBw/gVcRMoWpvrsbMF4kOi4R8+x8Ha2VMz/ECaonDxcpuycv61ME
s2LqUxB6FIr5FYHTffx2/bYV44eO4d3GwC/kAjik7PDmPwPq+kAOb1OlaxEERFAn
m0fEtvdesvtt5ZjyMz9IYahd5efPsnq9DklilUacXynb3BtbkkVzab5iYTVWQBYX
LzhWm+e/2WzpR5XzZxGD3ypzjzu0/h52bWxVBr2nsYZR5hWmEFXotE9qrOSWZa8W
ZQhlDoR+vcFBznaEOn7bhIs49ng0m8p3hzEdREplWgl65jKhrx/MBhtVthQUZ/mh
SyirG/lrcBn+aYF2gH1tyb+jFpYwL4nCSgtsBmhS91q4pea+Q9tW+ABbwThMHG8L
gvT2qyEwvYH1Y0/aaNSrPaBqgJJLlutiDvbNsE1y3k3OOKzqpuCpblxLSfzmS9X2
T8GIQwkVfjl7oH7pXe6vzYumgxmKRJCTA8HAhR8NUoSfZl0T9agR6GCUDOpfOXjm
1PrjOororznP+iNjp4YoWmaqdYHx5cGV/kLOLMzglaOz1iHM1Cqha0SVe8FI2Fdf
5DYfgvi+n2g203X4niB5I1PZBZGozbLFPzxcGglu5iYt3Hhm70HL2H/rITDerPhc
+lIZ9QR+auxs1oj3J9LtPQhewrQnnasSNFxjPQI6m4yCv0YgnmWI1zcnujGaZ0Nx
snwXGfnScLmpup8r0Frfo9PmyJAJ1MGwAXBCISAxZcWkRbdqGV64B8ASNvLQXpEB
wlpzAwmJS6WmtLUtHvTZAIDG+3COrUYMzzy1C53j+6U3k316ICfgmuOg1eXmgv98
f04y+UXUa7ZDMElwBxhtPJ/haa7hewcOzaONWPdoTa2G9flGZGMNVdTnhDbwBHcy
N3ifyWuu+cI2aP69z9oJVSM0jnTF8/YtxyUz/K+YAIHMUsw1zXmS7/a6t3AEkjiS
402JblAwb7GXwPlgC11mCQG4uW2H0U8NWhD5Gdc775U8UPZhXHw+2f4dis8FTsZH
kSiz9MDL2BZGBzVkfDWNihmpmo+6DlcCKlo/bA5TF0aA+qpBIrnFdcRjK8Tb9F2Y
m5ikEtCXlfFodVGN1wlntEcmtro2OECMec/bDN11b/OF7PyAlVfVOcA9umkXXbwz
tRuRkWYdY8qFQk00qRTi8AMpvYIyvyuZh/YSZOL4QJnDBCzGYej5vOGMBfcukzVZ
/fuJyJ90MmpAxUXEs/AbIbay84nM5LxixzBTPyGKquEYVmYn3h36F+C3AdQEmU2E
DPWpvFcBdVsw6SXldjMCA180Q3S0i9Iz64xZj8XL+GSBK18i67Aph3rQkeNQ5+Dz
5lMw+JKliCcHqoWEHCyuRRNUgNoFKcr1J49WwlvH0p/N6LWCCAteusLX7+QpUMoL
jHrSF1La6QCZEygPlo85PNycBWbM0r+fG7wkaQ7Z8MUB7KF8UfKumUoK/2h1Yge2
loPFQ023qHuOrB8fsLSFINTcFncWXyMfBGr8QFsBizXcIooCs/lbwgfPlGySSTOl
eUvQ6E28EFjpYub9Br7IA0+z/vsYmMAtSLLQSMexJWJg/TZvGNhQiVtsgSWHPVf/
vg2HkMvdksn3Bf2z1ZvvuBvtwvXNQJ79HcumYa8gcVgSo6/THP9lWSqwmJDbk2o9
p8yE35Upp3H3qcDCQ9j5vJSyH4oqI+uKDJgqQuvj2Jgoh04h1KLZAh2MRT83A/Cq
5H8j1e95UL6hV6X0p3xszIF4TFpdSPUpKjgLBMl5L1qQzDzKidyTu+4AWzgW9Lb2
hOK3QkU3zP5TJzhagKJit3YVxXLhGuGuOwn2vhU6t0lERG1Gr/gSaYPPYtRPsbJW
bxAnYl3DPgXqzu9DK2VF64sKpZsse2LT95nk5+DLQdz4KB5v5My+7/ZNz17+jexr
SBuM2xQzCuX2ZO+f974ECGwh/SixxHoCsc6bWc7MHXV02VKzm0ti+ZnhdZB7hEvO
9ZquGDy+c180UNdulV8+CmAz8o3y26PKLHdT7tu3zpN0lK3hsuuqZpr+WcPNrm1e
Ez+t/vrGwPXBPrC6Z/OWUdlC5To+oCd+I0s7IgLrfp0+cu76hgy2Y4ZoaC7NIGB4
K8wwX8a/Xn6EJPcvwH+UqURMe7DLpcMqPmmxfroJlmSJJu/EUzH1AdfGNkyXjhjT
pt2Kl7lmAmywxcD7gnUtlhEJCS0+RNWyy8QnQ842ZcyWjJt/ubbGj0vxFoBYZXPS
E5593xXwgqNzcxTr2EOZuQMuiGKwVJwQye149CNW/mz6F/biNDfhlWEhLnzNKBZe
wLNdSqTsCUJSf6UeqBLTtAuNqRNIw4jKYYX6I6z7w/Xn3Kb85yIhZOmZOYM25naC
sjsLxw0S53Kv5zlistrcy/zw2scRFkYyn/RHpkRS9PX31tUYfzUAPUrjdXp9PLcH
UNBgLONstqKVvQHN5IEezo2FR/aRA8f8lh5oJUv81HcVdl6npZvMD4ByQF3uPDiY
P7ieq2goWxiW7dH2ImSRhEP98okSbUixMpnOCIynMEJf43rEewr70iqaQtl2+BIS
mkHunmpW3USj92KdWJieRHwDywiCQQ5jGsOt/JUO5A5ugtCWhg6N27Ud3xPwgdkT
oqLO/JVOg2d5unWVScsIIkm2ead6G6IyX/2j4ADgKh6yBWj7oSSb9sCExQjXm7bA
fg3oMptH6/Dz2oG7BVqccsgec8MaXqAvyzbD+eBmbcFDB+XLXQlNACOKaHewR1BY
iYjwTyq2oXCkqQEZFydVEjlkIoW1ME/fwrIWrkaZ2zAVAsXJZWo9yJ0jUpCfECki
NEz41ySWHIKfId4nPVztD6mY+/IPn0g2S2zsXCVwfEesM//3Ou51IL9aAgcF6mtG
6uwFxmLbKe4a7Wl3wwl5Y+f06yDtDsuLp4t77wXRmxMQaNhOZyZYmwqfHFaaAuUG
Cy4g5zvCIHPXU9krT51Vz+o3axzx+3bD4gmVodlays8BKaOPHO9TkeFTAyU2V6jk
ofI7lp3F6S+3ao31Z7a/ywq50gad4/czfK5Orh7I5zeJgTW9s/gjkxBhRtUxf0LP
JlFVE6YgruA4GqUe1udcB/Yxfr6IYIZD5NWTXyhwc1j7/Yi1bNMPwGI/Fm1ScOp3
i0nhML/UFYwjbKbQnsgJQCUjbz9folmZR1wIT32/0PoDE48UFy//K/6zwcIuceWA
2y5CYVDnLi0AlZwzmxjJ8C4GBJIlcpgmYTs3of7fIUWXxsjNozPIqrv1eAYu9qTA
UxWhS6O//BsNCepg859zIrel4aJXOk8FKK/tG+Q4OfgIpP6x93jSPhRTXwWsZtuW
XmUmuPFHDXKLcntBBk7Bgq5N6sWu6oFpVSt9SR/AKxAUqKxbvEWKUJVWPs0AtaCM
QW4jiiNJS+Ts3QdygVjkRjY2Yy4/5/Ncy5R6yNUzYW6ERdZm//BpjTh9ZPPRrFK6
tw+OhCtBwmQrOboFVzFWPGozjj+tEEbBbo9eK5Vt3vw7tzOlkeRrrwPfFCo+y+0E
+r0nxpynS6OfmRVNPr40fF4scRX0UR1seX1rIHPB1XQWva8AKg51NJ8+piSzGUE7
ntuUoXePrjb7dVgDjMG79hQO/SjRJgLkENQLmm3PKO+7/6WOQAzo9mncZ9s8JNiw
MlGbXQ2Gm9Zr02CEDHOfN5mQoZznPqQYym2gJfNwwQY3Au0xjhA68ZXb8zCU83ea
IdyjSH09G7QWzm7uDxjcikC5eTpilTh+g3DVVocPqaMb1GUIUjno3hwQKgwJu5fm
TaquCFNGxNq/nAm18BBfNsZaRStKHV2G8OxuR/hOsm1T95ErgsjdMt0FWzYKc0x3
Hs8qOrK77CKKZDzOmWgdTonqJPbTMD0Paf5xV4zh2Rd+mF+hcG/cKzbKSQu8o4NF
duOgvuulQtZaEfVoshSQrpd96n8ZfPz9tMdhFUxGwkFdUFzupNQb2yGJrgeJOovx
6CRWA39KPiwHxcK2c2vvG4Jugnxt+W+IMsgnNFCwCstygaDibvg9v3UNl8LxQv1F
nWUzgM5jIK0rvDrd+pl8B84L4Gt4StA5S80VtSegFaj7sJ01ns1aIUQEP+VH/PKB
9mQ+6vvw0hiOtfDdZoQQWBMPO0YCTgl9aJTEjLOoGVMsA22OFk8e6IHdMAIM4zQh
dMus88sbWHVIO3U7q4HF6DJKbVUl+VAJjzQzkZ6XrCnVf8jzMNRxVAoKlfJTvlvK
MQBnWlKkjIaliEK6LEbs4CaiovbLN6EKcShNiT+896HfTBazYqxMpz0mzQNpfDA8
iv7OS6qbOBElkOaviwOSK8cZjHZx/kDlKXjVWYL3tKLOe/Wunm20MrheM9Vc8UX7
f26cbkRfiqVRvpik1xN8H3GS+0TEi+Jeb/boVtLxn5eEjS70Sn+GpPpyajOpOne/
CGSj8VTcVXxHg6JzaU7T3/fILyP71zNxsiiAxsi6xIk2fjSrlAsEQ21ZdRSxlti0
B2RuIxCxgys3Cwe7T1Uyl/bO00pg6Qnh2OkQIDPX1uorqgsNq5UH5zWF2/f3laIk
iIH9klaelLnvZn5p30l0rUn9AjyzVYab2779imJi5UinqTqJvJnw0oHccCCBVidC
be0s5oAotQzkSLwIx1CLTo6l4ibmJO4316Uf/cLv6XOkTvceTRuiSDA+4RZembcS
dVFYnpGCzyAhXjg+FtqGyBCidYByxfkmqeXbVsPxmsKvATwmv16Wax8/1v8luFvj
eEl7l68bHw3GQ8uJj0gJ0SAX3GzZMiogDO8v0OkK/ti/iu3SOe2qF6BpZHkT5US+
eNiZJdYd7ftu+c/DvTnBz9Qki2m6t4DP3xBrD5uf5QBdBzmi+NalPVvdtJOseC+w
BUL8onTajgGJXyoo8SvPYiToG7bLDjBWabyXVpSjNY+KwT5BUp6knXcy9m8V5ndo
ym62KKe3CT2YsKIGLjjOZRBn9meyEyq+AdfnqZaDvnl2mV7OcWIHqeUIVMJEYSxz
bCO0xHb4k+S4zvCia6pMqABDWDf+6zwSBD8whJnyt8a5RqpdIX1tebXiq0sGrQyV
1/sLZFhQADHVIBUvK5y5WCOF3V9i5umPVsM/d+aCr4lGfokal5i+5L57Yrs4DlSd
E8fmcgxpuE1X8wb0El2rZot9nLgYB9S7XRt33Ro+QSjFM9cezfNC6cntbaOSXSdW
kkOxCQWtn6QyTaVva9cobZ6PvOg+TwemejzE2z6AjbXQIaFbGd3jfQJmaRfPSp1H
meHAta30+TtwsnoUadqxEVwDKiFRt6NniVLlaqD9aX9mHaKARdbiUsPf5IPb6GpK
4mWFCgiOQYsXq1k4qUx/hkEdcCAc1ISijJynpxFEvSrN79fo2DlZhTz9FHK9zw8/
LjJAQfmPhO+9MHoPKXReRDRxqxOkaKs24rcowAWXxJ/1sfb/P0Ibly9IAT5hghTu
CNxocyZEyVzPcOU8Zkj4InqDGm0vI9hFa5cWfge5akaFOBZ0y4640zN7jf3510N+
xzjjkE6WhF6Fo+CVAtoAOtoPhZHxyicorERjQVvMi2v9+WLs8mDG6H74Aiu7wDBM
dWgJK0c7DjjZiMOI0Z3OI4NYgFxbK1/ZFfVkt1zoLoNbR2d5tWQZuNdSlR4EhZBy
RfqZVaXLY0SW4Yr2W2s82prkgZG09xR5zKJwSVp+6xryKLRg0MF2nFCU0XaFCDJC
n7Vxtiyi/MNzRkV7INRs3RdAIzV86s/Qk37kNa8ORVPXbv/CTYyzSbfOlUbq8hlX
CZ6S0vxmyNZ/0oiqxUs3Ab4K/kK4saRrV+3C3JgvV7K1zCsP3z9OnurFe7cYXOel
wRL+hwKxcZWsusNEIdfYulkuAuurR221i1AeKGUXbJdUk0ypnuWzTZtg6N2ZLzvP
9lKB5kSWUQf2oZtBAxXSR7BT9v2M9Y1fWF+VgNC+J7UuFyE1KnBjEd3qgkYU6vkc
kJXnJuG7jupCgiIfVfQosT+P11PU2uXvoLG1im/Ak45ttVpIgzTUgC4tgiEmwI26
mstKBR7FtTLfuPQGiHWNTw+A61v9RixG5MBCUqV48i5Qb+mGH2XpqqIvPQpO8FsE
uN8tC567fJ3JtRf+4N5gBBejDUrhaYY8TPVQoXmg6y6lQ3M8xup5YdIGZ7EpllFr
818e2A1/hg1PmdTkltFxufxzFztKJsLViAeataI4ODCpANaFBYCGx6rciIcUKRxL
FCn0N+Q2pcKoLTZ7AUkNFoNjw2LL1q0px//JVFwL5PqmDffBooTMgADeZHQu8apc
n0TaiYRWQ4t+9NXfaQi1b3zWi4iB/2WM4YTsCXOhawB7aZ0OCEQcHAF5sc4U7eHv
OPvtfh/xiUAQhGa8UMEz2m0W5hziJRBZfPm3Lip4w8HqHQUHoXIN0iqZoniWImBl
crW1ZmFSqy2vwGwdNn2dFkzqYzKdArF3076WRy7T+aryQUD8ABiAHXFJ/Jx+wMqT
d8us8pZlSKbw/5YOF3BXMY7JXufFSBRJvxtdnCn4GFK9uAWsg+fzyd3LyQmH58Gr
4U67IlAIlAyqXppSjVA3t/sE3MTefYShn/PWlOs4GEM4m2lieYIgRrpC9KwzYtpM
+Mq3b+/n+9Vu6KY96cU5qi4yWIcGxmv2bu/Vu1QAvMVVb6abTElp/JhI3FGIkFvF
6BbDIG1iZ6W0fhdOfJhcHnCPfFml6h/Qu2I1L4Zugwp5e6v9mZdNWUaOnSo8I24y
/hLpInha0eW1L6jW1kpIfMUayDgyDZLU2cgncbCK8cAT46aOG1LWjSMppthQDLhm
BFR2QbciXiyjumdNCLD8/NJTtr+fVv1R+3aFDxhzX5FY94fLlZeOuSwK/CzgZLa+
eRg73f/zXcPoAl+J9tVhOzbOzboQa+BgCx7+6hFXfBoSUi/6sdsL4Hhcy/jeyGVp
KW/YSUJbwEf2BwWRTVMwJR6zEta9OZ7yBD1t+iXCZEn4uzJcyiirtuxxsbc+PmFM
URY8/w5YzvW4/l07yNz+ydIW+V8NS1f0fYURc24VYtV+El0Q9bzkc+RM97nM12Go
3KR5JAdqrLcu3Uhe96JF7gdvL4M4CxQv+fcZbBwmi6DJjFKrpckwqgY+oFGWgvP6
8xRsXi9r++UuBVZPgs20lZBSHxrvaSJ3Tw/8Nye8bCwvsRkoDXWSkapNV+qiGsC+
/VU+zFUZT2RG1jYPnx2EltDC5N2j1Xo2sKCP+XspnjDQT99J+mCfC1GTM+JVbDWr
UCnljtKUroTjdmHkiYTSbllOh1e0ry7iJDkBJtzPGxA2gc0Km5WIWfehIMPUzVF5
F74zbUVcIIy19+bpayhe+L1qfyNJXIBiU+AJMSZanmU5FaJbfw+pz+/GsHxqj3Y7
8TitX1vfkI+LNElbBUcfNELHv3Kf/ba+NlozI3iWZ+smmfy0+5c5dwHr3Ik8JIN6
cxaVLYUyJEcHGROut3EYskpBS7rGmhu/3CG4mD6gkzBjseaw4Yv6/btukQ7INhqS
QWsGiM6r9jbR2WI8bUSu8LR9SbJ2D36opqP0EA1VepgeO55eHYAQsPPN4TtqOtDr
gzBbCN5QjMEbaqvqQEb8JpAl6/d23x+U4pVRsNSajeGTJnt8V4n/aDrzUS/AJ7uV
kZu8X0YqQhMzSlhux09EtaO87pB9j/NP0vW7drOZcYehzZNsNImUkFC2QjC9zByv
ikOhmBQsOGzFl0qIu/M77paIHJjQiyPK8M+nz1pD4q5xqwcvVtDc5oV53ew7I3mz
OhYzvpepJVy0lWMHojMrt/qD6mm3nH7oavKrWo1zW8M4cLt5KyjbVgPGJMunjIgT
qvVDWGFX6xGPbAVF/KGDjkvuWPF+vIbd+/nv1WDQ/h4gWbl/nn/YEQsNMXMYAXZk
5CX0pE8pJdUvd4Si0PL6gblLViFJ7N8kINoiXGZJg3RXTw+e2RAd3U0IivQ/2VJV
bCn7Gy3OdzmdLJhi8WqnMld3BmncIPQSD5cvSy7oUyBZS/1uePsr/RY9cuZqkGhO
vnI2p3HCUq/dqtaVOIQqf+0887jjGxsfZFHZJfwc9pBi6GNnu1YmQrw1xlgXnxxH
XZgD36NiBLUikaAS1+9rxYodHlF8l7THm979/bacwCsa0N47kLjzc9TVffSCz2v+
BaL0wFCyENNtbzzol+ilqLQxCMCaeiKhLfUNgM67syipbzfpju7S4H10F2iHerv0
FFL4JJScjQL/Y4xUk9/fUmiBxdlHNwV6dgUFEnotGa6Wvlou4RC+PwkQf3lYJeGY
qCZKA9VRvAwmMC8G8AeT/t/neCYNyJQJRrWx/N+jdrfsFVGl1Ls4+ujxBP/tMwtR
d2p1VJ5xhLs0xC9ZONO5xHRM05RSZ9rw6lRjn2y49A5k6CQ+rdVu15M7YMJ+q78Y
Ew7NcECxJZhqm/FVobBU037PsnyYaGx/GldoWfcCQ3vUFo/87x7quYKyLYDaaEjX
RSB14jozMCpFW9FgG5ADowLDSSwRCSHQGCzeZ6+jUunb62uOxhjBareRYce96P31
SHp+kZTLN6RiF5/gp+Ln93XSR3kU5WmvKqd56atFWuG4qBRsmJmDM08QUx5GTf7e
PA0LB5BgLqyb3+Dxyuoc8StzwSRzKPDJZUFnPIspRunfEi4uJp4KoQc/GDmUYVYX
5aoP6ud1KJBFyN1U/nbwuM0CVExXJK/18QChB0KQ2Mksm2xrcfh6M5nI6Q6/+rop
qXra0NA1c+onkBODs8VlF+dfdTsDXF+7JOlwpWaUoYjtED8xjc92DUt4JCQYRDU5
XA5IFuVoCPdveZKCQJ+WkTIg91JAL87YE7sMvhw5OUWj3m0sAZ+YEiaKgLuCQYzx
cWulYDPUvxmBAbF1l/ueqNFhnf4Lnl6dttKkFJUJBCBtGFACn0NVIT0F+eW2oQ0l
DDyOPiwUko7S5BZB0S6KRLbVZgXnVUa9kNcgtpBGgtOjDUFerC742bKxIx6WjHQT
z1B2dcrtqEUq4y2+imAbdQYGzq0OdaMMsrcbmciy2AT7sFX+fRo0KtwC1pe6o5U8
JvhNRyGBjPqkBfGtmiuzli675MFSKOjFQWAWmzjL8utn8GLLQxJF/3j89tB/ZeWw
3occDMYprdfsI7ZlJK+bAdSg5cie7eKAnNM6HjPvok18Mj++DfHi1dV+/gvIO1Qi
ZLCWiMCD+C35Ncr3K+F2bJ/DNAXwh2BaOFt1HO2PXL+DZxF89DGx/h8Jku/O0+IJ
voAv6DDTL80zLKKQlKCCq1JHt0m0+BrPC25XUu9pLCwY7o/xKelQUnJD3ojhrhqL
miPr0t0WrD1STTUEZN2qrNYDwk5wZ8GnioJ83O5qc9E6v7qMfGw9Ji8LIB5Il4jP
Bw3GmtPcb/mXFHPcf78VZlLGl6VI2kOmtRh/p0x1ecQYnL7LA9C/Z/tLYAXp7MWe
j2xWEKGPeaQCpuNRLajx+Tfi5SPQtSRJ5mJIvetNAMp234WzqhylWhSENAiL+Q4u
C2HLzw1w9MmaFokuYn0pGN+dZLxgldJ5JHtnzDpGoOHeVoEuDhpYchQaASsGVUw2
6tXemvLB4hWb1aOT4Gqdk5ZloshEKo7jbGomw089pYnAFjRJnVwZIR1AlRUNq+nA
np46lnvooG1+0TOkhKG4mOoYPFABLDpM2AQQ0i2Mf6ok1sQ8FiH2f1uCPKGWfod0
dR9rmDar8udlvceaAOyPS6PY9V85rE8jM5QazMMdRSVFi7Odt2RgSUXBxPVEb1Vl
lhk+dE9rWszDQhgMLCuiGIMirB/afYc3TAABG/hYJ0BuVyj6kswxWNUKmxkyOD45
0sXeoxUsPZG+fWWWQg+ZXryeeMVZ6QZbl+e48Lf1r/I5ssmQL3sZ4hxi4HYk8nWd
gTrbb93lCaC2wReh3jyeNNCgIqjhHfduoJy8EjhcJ2AsfMhCCXy7Nudloj+qVM2w
EdTMIElItE9yy7PCVzmduUVPFoHAUEr8fvdRau6c1jzN5TCTASyvsJg88zkQHF9o
1GNHQqivFh3dTepZo0ENy1kdrvmR2+NOF85NeewxSGrWtLY1cA+kRs8Nnp/A6MeD
bBp94yMQ6uKsiI3e/xxjXQVkbu6oJIDbY86UKAnpMSEhVYJQlL56CIMoc/O/Vl3K
MZOTOx0zB3GcRKT5F7x1ZUn7F8SdQwOdBhP36j6TKVe8nTpIEcB0dmndua8NgRw0
6dESAuFASjCZa+wchzUOGJw8UXfokXS1u/eeiv3Bl7mCXnwF/izd7L9hfso25sY+
6TgQfv6kbjdyOV39L72U8qH76kfEs0I+ccAtj2e8VwAt+jtUr9lkAXQvmtoNGqc0
fbx+SwdwqYPixXkxWdXpL42b6fh013XkH938ykB+AUdd8h6Oln7IgP8jYdj0+T36
8oIYGhpkReWHU+J/UuxbID+ky8eQuR/no9qwPt+Fs9qv90YUf8ClUde/c1GKGjJr
bQzWagcAnUquZA9G3Ke/cfLb+sCrCUN7B3oGfWbOgjCbOIfDSLa9obDVB73jFBSv
X1eWYmAWq7ui45LALBJL9paaBqhUSwoBjebLWz9o+gOYmWPMLRNFPXaOWeOjSpBr
bJSLPSSwoKwIrz7Nflz6Nbmhi+RNYC8/t2y/kqhsiYBolv6FinaybCpyx8nmYIcS
62/pdAzJ/ti5sjIiEAPgvXylSIqNR/g2tlsbBPJuJ/oz1By8q1nyy9IaD4FddItW
rIn7eFFdh/DNXPd3gS0HhBKaIVmI1c/d1gOkD8WAlqY2ezWjnIyrgmmSRKTvpysO
CQHrOK5n+uAWMjxXDlPbdDnmcgQzHixi6EB+/rLwaLWn83FZWPuaqowDlq35HCmL
W4KUD7AqU2E2PcjN6HyJ2Wdi6QphIU3SxBT/hJhbRD27XyuZEjjaO5ydFuYVv8hm
Qy/5uA8bwptIJhaCHepkEKc3VJGN0FZGqVEQ/p0iIygXoum55WLmrDHMR6L1dJfi
KwBo0CucJcvrvViazFUuzI7DwGUKb6JB03PyHcR6tD6N7/tGVXfWbhdyec+k/EvB
0NTHedjoGTnnEcTDeoWcoGEbHrlzyaiNL5YZt9B6rtYOi8Bj8uMogCY4cMyn4C7x
zy3PoBx+MC50vmZhiqW0Ep55Jf65rUjoTn1W9VYsBsIYSg9TrvcJSDqcOHIIMIat
OGMdgZVt3H/r3ZVsKtRTXcv2Bp08uVoznRx24J38CCvNqjA2Z/S2sptxWl5Fu6Zs
xuHdTv0QNSxkqKMvyYCG+Wx18/IHZzQW7xkrC+DExnDJar1XNNwg0Jt85XZDehwV
E7iIi30CCd5+2Ogjdk1D9pS8pjmfq1ZdzP37C3VykD7bW1Roc13j5NCkgAPJ4q5u
pwYyjAHdL+KC/MFD2bAD3gg6BO0BPk9SEZMsQZd/KkxQtqTDUS7nmsukwW50ZraE
Wa8bP4WGTPkgV7Joo4bMs1K2orDeud33r/3cLjlOEy0HpY52+qskkwRIZ3O7msQ2
D4EW/WPfnCy+q5wh31BHSjoRR9ugKuoxG9FrUArIl+BQhf/GuojZN87JW3wCA2q5
mmMRedTIIFf7eHxFjENmCY8UrSkOyUeqP/D7aUDsLIQ1omuc8HEAkgcHO4suspZJ
ko7qop9s8WiEkYo6YH7H/DUhJMdisP3DQqK2ZCVUmDRtHHAq02Red3PaJbyzbkaj
xDVrDazG2nLiLetGvlmK2Ww4R6xxFS4+ymsd1+8Wat5Wufc6bUtSA+zhhDMiqCPd
mJsgRgmtxCp5lXRAE1sVeiCcREKwp3xRKXYtLratjTmkk2lN0Pzl4cNDfHJRnb+C
JyvutywCIlGUmKsXa/JgF1a6AWB4cs+zJnVWJ/nbRK1cBemUiGFuAWWDrWYwEBKG
rYqOYYTztXag1cTpPh3uV3l68/WfJnp13xeiNdxxdoQmvBCnAgVSyNhWWIeZh0cU
N9qazv76ie8lEtFAE2VriX/5iEL7hPgB1vJdsCIipz6uD9OWkw6BC4StnqEBZxKX
QJd8TITKaQagU6WQeiw67jzmC+XNhtTXvb2sy7kwURLALucyutseFuAJ1UwYaxtu
CowkV5neH7dJCx6IgSCAANWWL+G9VK3rBkF7bnMlYXMN4Xfly/LpmYz+NjPqoga2
oCnhkKxOvRFcYRRg3FshG5yqZAWP3C+tWy9bKtf+w5cGS51S/G7nex8q6DmM3J99
97DkOFR4ErlQ0ftyHH3piXNtAeooGiI+NxwecOC9CjsZ6Bg/tKLYKBO3S8FWgYZ6
w+SSLse+FxlT0Y//C3JOrMnwUWX8v214GKiaBCVttbIhZLrUqRpE/1My6TUZG1rV
rfIv3TPB+SKlux7kKT5s/l/jhJHlorTSTE3UkaLeBVH/86h/QeKbu+vb3S6wDcpw
HeHPIUVj55qc1gUiM9woSzAakThuuY2wq82mBlfMsx/DTeeQxajF9GlC4Pi1GEn4
DUW+mvLO36KzWxfTFmvSdqUcnXFSDVVBJKBzaxPakU16dWN8nxt6mHD/ek1bm02Z
BB6Qz6wCjEN11gch0IlnJ+OwS9JeFZxVOeVySUTtv6+05+RPxN8u4MzIQXKPOhkE
4DiFMhyLZXdnvB0jhuPMAOXUzbkgZXnbsTJaNlArysLWKq5J2TIBFSyMOS5+zDU2
ClNjEIdpzKynfDHyIHOpMF65VsEI1VWv8V4RGrcwEGSxaz6IrE+bF+B4zJJwkVHK
EiIIC/WppvxKu6olCC8JlT3cOyhO6cwGs7m4t79SoWQrtr8wKFlZJDtUXdM3ADKd
jMF9C06zMmjLruYcMrs9kwSE61mLi82TpJKFhQMbW7/6+0PN3dcPIKRA+xotuf6m
/uMLV9L7L4o20m+ByjIEtVYQTdLSElNrvLJFUfrEJf6cYQ49O++vFeO2Ztjf6lRS
sBqd4X2oB9l/Qv4DrvKkJMm3bsieWqXFH21L/sbbyNU2yQCSdscrpkFqnS9gnI1+
z4aQh8o7qEZjU6DmwWR/kILr/uqVdtseUHr9EnUrH2HqDjJ6UREVAcnZBpgLKqc4
qPy7771AYs/QE5VNCwQCjSKmd1Y3MJDWWdJKgrbgygnjFjla8ThETgseaI+1U28z
EzjnlrmxsxtVGboSsp0JhvQv2zyPJO+hDPZIx/aeEEZV1dtbIosj6txMtQur9T8v
1RI4cccBirF3ZCEJT6clOh2jy4xMEukjliHHmQh1INfXeiaFSeSCm0ZW1wMeNB5H
p+6z/91G+IqoLfZZMxJAHXqVBiitkTYtsxbptCrfbo8Ab4gjd2Va7FdewEfWcVbF
iFie8WhYNnFikanOEcQoKorlRKoczVaWX2Amui8o/mjngoeUSH8vwhabeO1MghfS
WKcS84lg+6cYI8ko+d2W0iWOfPw9qn472gMr+FHEQCkkMzyrUApraqeeBAyc/RJS
OU5Q9utTaP6wIVkEeJsctRIEQpk/x12Sqi3KDAiTnKytyWK70UPcfEDYYZA5UIMB
yE32s/dozIhk9yM0xmZPVuK4W3VwiZztkpVmcdGdSD7tIRypjhU1CrFIdrSQ66Dh
HhxWcPpkQZyA4/5hm+bzh5r7L8iqqCbz69Cg3ybmfg9MyRxn1ioNAw1hkrZrbImv
TT4nTuLvvqxi4SRMrBE0tyWOqGVPk884UszQjP4skmTTR/wpPYi9Xq/IAg4BIG7+
/thY0bsBhby7xkfnx/WJudFOgrjOqaguO62aXqCCEXq5ynJOwVemTFMx+2cWUqT4
vk3APp/TNtK6XDH4+lcWD/SqDUoV81JxG4DhqwCbUNj5/bILx/Q+Swg/MeOCtIar
DtQxBNPyUE5/r85fPjxT3qM7bv4qKSgNKy3qrfxegNorkF39T1HfViAIqYX1KjIq
Vdzz/PnPQwV3tyqezoEYuSR2gRwgAnkmqscdxRN8fwtvfqPK4PbqiWiGhSXQzBrK
PgFJXQfVnJ5vlBo4e0iPHuStJbMcFo3711md3bngmFMGxR93mhTBPh8Lsssh0EQp
bhdvLxUvgbokP322ZAVsFHz6bhml9x3pBD8IL4L+JYRCAK9aD47GejVTpT60tdWZ
/KyjTj835QSrwT1P3C7p6XWkLd6ky66cHB7SbN7yRohBcZbvgpfpyvXvEniU1N7K
HFhAsbdGEKqajf363sezN5Mx4e6OKRSQjpuhiFmSSQVCE7UQGvEH5UyIOrIbppoi
KoAFjz6X3b0mmb4VkYAiY7vlN3H7yovE0oB9QGWpIGQzghD9y249k+Wx/KRe0K7q
DQW8qyDOiPwBfX5jucXpWvReVvtlVyadEKOY0XfxNA8gnc8U5//K3WiVs6/xrJam
VotUuZ1y6M/iZIG8K6aftaHFpVLTr71zBxqG9iJewcpZCIRku1GmFsVOqmWY7Z7c
KXbPDL3PnhKgvbVX3hOwbWQAjKMbeB0Z/j1dHDhK0BSUcVmpBDrhfuTQTyTlj2Xp
VfLxeTVACIuFNF1/oVNnPfHcsxfTUYb6H4TfenRTzGoZrg5pSlXFHJx+yGd0E3Ap
jqAru4lULHm77Aeh6tNjOTnijFU17tnsuoKY508z8UYn4uwCx6pquXzgw1Z5MKgH
iB9Ff8m2SGP8f71/mTXN5yv7kTtmHwaZZov5KxIsflsG5mKIiXx7UFNDT4aPIoVQ
8VOVlLCB8GUoBbRBeH8qsFXKz/l3aJ1VmruWs6xz2MHxFgbgTWzqBLB3mkvfda8v
GaIZjXmy0tCSwRrBLikARXyz9fCMThcMPtiadbJz39Ue8cpT9YICmm1579iwziFe
1Wop/OLS0+EofQvfBr9s2Y3VBtCjbnSXiePGTgaRCX0=
`protect END_PROTECTED
