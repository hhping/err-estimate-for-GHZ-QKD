`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7pPKwfOLs+sSn3CtkzaQw0VO0VLR3aGsw2I0x85N10ionO3V1DWGer8ukIteds/
QRsDCJteHwthwvW/a9YdgangeAwZeObOQgf0TalSY8zX2ERB6VgtOZ8JCoNlaIMt
IhgTIjBlonIAXoM+edHu7gRZaz/JctCn3vmfojtb5uU3CWZAAv8UjEF41TcCkC1a
zvtdntigAKe6+epuvbRO5I1GXq6v8pa4XOIRjvPkTov+9HiTZ15bowIrywhqJhfE
fhW0epySdU/vRJ7P+HEdG0oGwdMIy1tIdNWqlfx+9AXwESW1M8tot094EjLqtNZK
msbAUORk2AxB+KJ4qhiFxmFyjPx4p4VHfVL2tdBR24zvJqTBi6jJc9Ec7i7KL7Y2
6zEDmOBRKbYA2dySeFZbFPHkbs7xAox91vTfOfTAOIEwrGPeDiR931/jr2h1VnLt
5zNBmcPaGg7m6+57gon9+a0dT1tb3uIw//6j0fYaK1Lu0YJsQOF7AlvsLPUv3rQW
s5QyZ67osI7TI1lWPkWlioVmeGX17NPwUdq5DOL7QBTutLhpmEIUMwJzI26vVBTW
Gun4FbY7ZhfImHUncMQOUQp7Qm4MymQhykNH4XHz3hx5Pcu/778Vgq4OR/TvYCG1
iYUcjrA/2fgB9FX2VMSt3e+OmTxBYtSb8JcLeOe+CaYGAZJN6yqpcRlHFrBbpLyI
MDJb+OXfTZ4SAuKsmB9gcDj8Fc+sr2reXit2HJS1Gl/0jArQYMXD3uGyg0DMZG7T
Sef4Dkcow9WRegRyta63eSr/CzusOasvHH5AQKtQB3EnJJ8QQeo+pD7om8FxMEqc
+t+8/YSgPG3zvkDUmoqDZJo4Mfb5xzW9ceVg0Azxqh0DHCXvsxRLhXtZHX1ZWIDc
HJfJQP9Z9uF2nUXiDD8Wsx7gb0BtcqaXU4UOVWGwbJHTvmBs6zOtNQsshTHq8GYr
gjXu2TwsTXZRY2e6OuxNfsIGoJ+nGFQmSHhgoF5RsP5USa9q2GNAqA9doT1tgvt+
89XmblowizDVfL5tl8oc92mEM1LNl3OxQJNL4ZCPsUBZNFmxWpjYmbT4iuy0TuQg
n46LaZUYcuat5Wy51NNEoO0rNNES0HsA28lQI4BKzrZFoGUVhegPCzoZSA1SCXVP
w/z3mu2D9X6L2/Qa+Pz2rOu5AT72FmqLvLnVVRxC9Fxi4CEY8yizuqsv7btzmZ4E
PQWbtHgjxSuU/Zz46qOqS46A0UMaqDcINWdwbrNjN/WpQ0aEIqrvu+oaTMEA6Dg7
6QzbGBulSf4qm03nb7gQ0Ll7U0fGACs9G4s0ypBIVWvhLGPzKgeMf2TzESGb7FJZ
9nJS1cclHEiHhf+J4wK5B8T60Qy3e4+j+d3JacH6yq4/GSrXueTZ3bFz80R64WyA
UpJB1cshrC5VpNnS/amCb60X/zew4wZ83CVGxwSQgQeRvcUzY5D1NVyp5o02hJQy
OVkTDPO4yiI5UaV5CikiOCclHd9ikpQjL2ybigbkFHOt1LaXH4POw5B2tdHJWgJ/
i2DyNxWtGcpYvKpB7B42LT1d9WCosACUdIb8cnCJOAxuHj4w26nmRxgYl7mBX85d
Gj7DNTCiyvhOYj1s0gZXuGYrAhrusDScZtovK8sAOPuAJgBSq6Zrg8CoWJ8nQXhe
aB8YNQEK1i+yGdAycEhxbHJyZj91bKECxhpLoubF2HcB2VoB9kSIzfVpYHOkFvxq
h4PiD493HvSAXsdtNGdsJUPLcStglbTJrC8ApTIw3GQ/ZZeEw0N1BefeuaTLlMzC
WPGxxoPzMHL9c305UfWR5af/Pqmo9IQRu8lpt01JiNuyMUaC8B/QIbV1Su1dt/Wd
ubAkV8lDFkwiy8F3hc2BjQhj747Ud5uRX6cegrpO9LI7C0bOnLnAVjFHRX6Dmuan
Te5ZWA4EjFWEKMNKyCeXen7WoW3RcVcr9d0eoJbnXXxhciRDLjFVSi4Aw5QpeftA
3yycwyj7ZR632Q8YwhOCLEWOGjLj5my4W1a1erQO2UJv/OR0Oe4TDAf0rdZO480w
9trNYnHmFykk17ECZ1h4QB0f2EUBMovFyE+MFmDb7/TxBk/fZYL2jfMsvxiPFhKC
gOT1whkGMyX2sZ+ba+Yh3qBIkjc9sYDRxCSwYcbGyy/JAjYgX2OFsGN2dtV9Dy47
44jW/7jtqMW60y4LTylakzTwJ8eAl2ouxlM219rO4IJiEM2Rsj1Rq3wEjuQ+ERSc
RRYStkH/BiO9XZQpzM9Bn1ge3vUYw1HjzoTZPYDEpjNxVDB9zdHOeVun99L/c+2x
Dd6RZl1BYEhHLSDvbj6gaFa6A5JGeIaEEzdWV0h3kWaufFa7HvpmW9qAJpbmM5rT
LVDFMk3mSved6GcM4UghSJznyAreul23QawS0AbIiVQT1lBy4ZjZbqcVdlvZJPWC
XoCA8KxCpuzTJR53EH9rC+ij/uvrr8exUB/Gsksqfckvp6OHSGDndxypetM0zDkG
MB+xxUZVPeDOrOxvvPCEZC+HBfnS21D4wDGwKI33xTRMeYMzyE8Wzz+8Wdd87aYu
fFk7BGqlmzULNbWviCkbYfoT1n1+DQ5B/b6E2HvrBQol3AO/tuC/97h1QFRcAzjU
wsfKCft6rUcWEgnvNC2OwAsHHitwLTpinYYj7E8JCrZB3cC0R+Va1xmlAocN0vly
N9+EVJFdzHCf7aFPPtMx9mFp57aBF728760dkP5SQ9Iz2LElLu6Aczvew3wLOMhd
0H3Rss/RCl0qDDj2br55ms4+v51QAHXDcFBuIuY4y4Up6IbSpSzNf/qZEzJodkYr
rqrTpnR6pAc1q9Sh8IEfUeyqKsh0QblGcgak8EIWT4b1IF919GNMQ4c8L/GX6yto
DV1y788NuaDGswwLr8keem3dIxH3PKR8PQiRajCdwIz2H4CU0LDJTJcqj+L7heVj
wV+Gpk/XYjlh4KO55h/ndFS2DYNLQXRmB/UT24eySDBx0gkKBBtoLx290FiHlxt5
NpSA2WKaty6Af1GRHtw8PYipgdWLsm/SewvmDnbYjQ0/0bz2aoahlbT8GxN/g1P0
1O16GR9VyU5yxBaGME/laYxYSTvLKNBuvn9CTRiVBwAtKqq2bDa0Y4qtr7yJWUSR
HakvLtYxIi/oX8wz09RuI6nGRLjc994IGmxCVykx3xD+F9jXPmk0xdFKIS7lJtMe
MBiIbtVlBl0mdjJcsbu0Uupde8dKtLzuoPuhl70u+8wJw7jhtgQvqWwrKjY+MbJp
KaBg8XIxY5aVP8PJlmIq9WWdNkYIFElzvgCNQfnTflSBljec0fM1dNp1kTd0A+6O
LdMFnLDV4uDWOwTfyWxtYDfw0o5ZvuiWmh+1Xaipb3GmFyO4B+E0XoOm/iAx0VmA
3ZORx+WwsmSuYCq2NJuo8XR0ysuzYDF39SKZPHLAlOJv24Te21tafurTC3U44EnX
IRIZPzqL2S8m0d/DeNhwJuhUgGWlE3NiP0k5ryl94o/TUhB75u0hmr/S2UgJfv8S
8fz+TSdyB2bAYmpW9nOuLmVHDR1whVBl2SQjcyBLq9dxqCdrIDn0CgyWzg0cQ8VJ
+KNkCStmxDvtxzojMs00cGAXv9L+F2RCl/knS27aJ53RHiKfKdzKe40hi/1ilNZo
4JhtOWynv6pwIUb+BqZpqlrO22tPo4lgTTpUZmMpOU71bMu8GDOgy28dBYpTEjVp
XOmXGaoqTD3Tz9YHIO4V6R7JmKM3uebLtFvBy1DSr99hehtS2ZJwD8fPWwWDXhz2
PM6kbzNUBDdfhzG0sY7rTg/DXdLgOz0ZyicEHgQ1H/5G330MJ5i3D7ysDRy48QEO
ofPUPOg+Tavax/VIjnYta3W7Sm/M908scBVdaspWY1jz77N3VGX5JMZ7+onecyHz
+d4rM5DV7oauPLN2HSxgrUFPMsuw0EQrWyFWjPbOVX6CrrIoQPONtQAl9TR1YUxn
maQj9zQjndIfpC63ErUeGQ/+Qwxf2hIerKsjEGzOZ3L4LbDzT2xDEusYXa7PU8/g
urTB1E4aVZsQmiUmsF3jRL8X01S/cx2sxMV2LcFNmrHX46sl9RvTJwZ76JxIWH86
/eKPPKJmpWDl+OL7lVnuddsrkyJW5gT336UKOD+AEqjFlGGPiyVicacLu20pWqbc
2KH/no4fo5XqJ2IDjeS0oHawrkoSnz4d67n8PPOxZe1N1m9bzhjzWeiIOfJ5p4Je
YDgqDItWg26CkatgOSZL/TDr4oAkqKyD+IRAVEwJGLneFPJLCAMRO5mZ9LTd2MZN
rWvXwJ6Q2yMlHbOShqdOOvFEwCCIByofH5Xdx95Fg+dG7WbSe8PiZBz1olCNYFQ9
JV5OpPHyEYKukK73cH4utg9YszaDgbsGmHEKDBqOXweSSwCWIPiwe1gM3NXFdsw5
vjMjsB0izMcYHyIT8yoqGnKsYz7Dhwbme3o2aN8ij3G79y9tgE91o5jybV3NAlA/
YrZ3ULk1kskI7Ev8y8OmNH9akhEG71xAxSrwj5NkIyzBYvRiI9VKTMpSpoJpNdP4
8GbXxy5h1SPFLLCYgbPZkZQ/LAO9pU5BoBspn3xGLvnIWCpNtkFYnLOcg2DSSHV+
EtHVTfTZasiLOqG+Bm1s9i5QbSZBLbFVRv2N7nqd6NN69s5MSxpmeeUC36b0fIlI
YPipgJMtV/IriBYZ3wmkeVmfQY10J3iX2PHMSf8mwq0Y+2uAiijjEzgiH3CYJRt5
vUMq2Bhb+K7oVe+45mWg8Vzc503HdevHLJBzvsWOUfMeuaL0x/vhW11XKyLEdoeq
c96elzRM2Xcc1Q04aO+u73PZGwCmHohg6taxtPJno21KKX2wvPnJmquW2cgW+0Bc
gikVmZ+pk6wvgFmQlLozCblE6zCcM5bVSyuV4oWrcRx3uIe9eCsC0kuWCm9XD4A0
cuIbcjr+nCWHyMnZAXT9KhoO1JYfDvF4serotLtfPLp4AGMkuJLdKK15VfJ/IJFX
Gvo6YLDffhU+LE7jtfXU+rZVKPEP3xxspxhD9dOiV0OTGCPa5+BJSJS88jfNVtCR
OeBwd6SiawOrZS4pWm5SHx7Z27P0oHZ8K3zfQGhcMV7DLYpRo9NiUZPZGgiCNop/
GJO2/CJ7iP+fibwYaXLB9s95XBWIsW7jEfNYKTDEG54ld0K0DQ/5OSA/Dr/AOH9s
lzFKJPeOnWzD8uuM6vKqLOfAdxaATFydoLTfwQANnXxTh4Y1zPcyI92A4ZZ2dSHx
1j5XqWs6TZOlL6ovMmFk1SCcvTnYtLFfS5uTPiWoOFuazpaVSwtWxVn/2FksCoQB
1/WBW0QIpQIAWO02FtPxWElLaQpTSqVZF1nhCW1pwPZdWM/sGodbjDm79X6VcUzo
MJh4uCm25NcT0qi+j2gPvtLjgLH1ySZVwHQKAlH1qpaByX4n1dSUXOuzMnBTBgS/
4oWRYQRkHo4fQh5KUJtdsC20DpA1yZS4aVmAdr0vxSs30QyZrsAkGWaju8Rqcjn9
Os0/8j9VqQ9DiJt123gpa7wN1cJy0d0kfiYVo9F1bnfgfIW+BKVsSyofTbphV6CI
ADBlyABkOvDbFeT2SfSdOI/QA0PtGmaXSWkcsG9O8PlJ4JPK/sHIvY2YkKi2N5vV
+dNhq0OEZTu4gAJoC/0j5wZA76pgLxPy9Vk1yTo5RHfzvz4qWOSeD3lvsaWQYngV
c8r+z+Xl/dbcO5knlEifuAqwz9xfBdxEyeQ8UhEEkxQbfhXUxA5TzezguVL+rLJq
z5paIzrgapA7xInMPfwmYorPbd/JfzU0DLDp+KZoS5K8SHDKkD6rHQfvv+sKT1io
cdksa+AWTpU6AAgYsVdudA7GP/VDwVDLA2nnj6boFN6li7YfkRt5x3RRlHDCzJ33
tRtRhqRfmEBGBjbSMeWU/e9WXblnJxZQaEWTmcY7bOUN+9HPA0iTon5vPR8HfifU
d0C+hj9vRZm6WL/XDT1xricaf5tEC6q0mJ0cnGFssn7ptSuRoM05Aip5CCaguDEn
17uWzQs2goSr7G4fumshdgYPqanhQKIvCeEmCNFcuw/NdLyrw7DSko8uPW8ItK3g
s6i+q+YZ/1+Hljp5RsDYS30zgtQw+yOhluAqvHDjK0SXfGmUFqoSYwjwEZdje3KZ
M52rvVZYv1B/mGZ3d9TLro1NHWJ76kQsgVQw3mYy0IUO9TPzagb9qZ/YIhFqoYzq
2GPfQFq5Z//IoxWfNwsMknNA+pyoN1B+EA91tK31wm66F3GFTihJ6ngHNocb4F92
3JrtjHjBFzdIxMPh0qlPvZoioIDaL+HX16I9GS/MpIJflXpRBh5wRMtdB/wLWs+8
8h8YLH4npF2JNWbKDk+LlX0Pe2ZYQVO1OdwmCc+3gdC7EzpsPqDtzZoGzinp7Y10
DMOjMcZoqX87cTfw2+/zp86Sy+E8NNJ3n3krEtDqezcaWeqx4NtzDzsQPt3RQdSC
mbpJ26+rAG2EbIk/d1EamGeC/l6Oie61kn30cpdY5Xzz7MBx1q62dFyr8oGgrltj
/AMSqOs/ZVwTswLHQZSxNkt02mSpO94xniLVuoJxRtqF+ZezwQcUAQttD9aY7b4y
Ffybv4CTDhlK+lUfsVrQlNkQXLGoSpPMvmdCt/a6iX1XvLsVPdeTIfRsMnGXNc1j
ox0u+6gWJSta6UWV6DO1U6gfCheS96oUIDkewDxTsmcTe1AIHkj9699k+bSTYbmF
HiUXjnfm41JsWu+PjTcSw1fTsYcZ1tCV7eIqiDVyVU/FcZJy3hplHqnO7Sy1PmXX
GElLbFPaIVIjfqZ0vdt50sk8T8WWDGI8rEfdiKkGH/mgABrJXHyl8/6mupXsOWWL
Km224pGZDjE0MJBzFTHnhH4zN17Wo4NHdQDVbhoz5Ja+8MKTRP1YPPJdR0xV5Da0
rFL2rus3CdWJDAnqe5NlI+y4eqBzjYWHWcfWSE6HtGdNPpojyP93ObcaTGBZyjeE
JQlcowOVjrVKFkfzj6P+aC/0vCN5bFbCB/Doc1eYP0X5f4+dPqkYlOsXq7IrhMeW
jCJFssB/ReaHcX8IUYUdUtCti8nN7lgHXQ1Pk6XxnfQ2dyUU4Xba/Q3yT8QPVudv
l3tp4l6h27Bp66ilpHLmbM7cEtLnUdZi9aKF4aL0odPbUDt5ha0ms+kxGv779LT+
m8aNWhQuEm/4BVuB0KO8yx+9yfYCT0znsKTMUdVEQRBICOStpVTk7xdGIsaKXqkf
RoaKXIZQx5qptCPaPwakefPQwQ8ixFBD3UqoX8pkvSmjg5Npssd5guIc3z5TwZuy
6h/9QUPpyOJoUDxenXtp+yGyjm5tJOIMaSZiWz5jidc21fD11/rUPW2K+85Rbowi
gMEtHs9LLcEkW6CjziehmpkOjbZCDZX3TEzwQDJ117QLYo4p1GYfIBNKJlcTPIDh
cFYKHCEKo0cuy6KWHeBqo0E66U8MJjOggHvf6X5eOY6nwDibZBasQoLBHtU0wnzz
iEd2t9CMIujpFs0LteyPYynaRAQPmEU+YxFZM7wS4wv5ufn78zwe1h3/31Jm1JJ5
glCw7A855y1sR/k0NSa3b/g0grNVfqWq4Q8QLuzW6KDB+WNvgAEHWAisUiTuV6WJ
2n9i14f79AGT3laytjHCb2Ui3+b2W6y0AW6XvKZIxMCgCkUXzILmUo/fGSyFgYH8
4p9EJ3k3Nl5DYrKvy02qbZRcN+kBzrhuDq26diHnymL8lIg+V6iZm6b1j4M5Zz3k
F1vrjBsJfQfRob+7Xh1XSRWbSCG2JU4qgZ4Ze8gVIBgga7Lp5zNIj/9souH3wPlK
AVQEXpm87j9Tsnq66HbHgBbKOs5eobqbFSJVO7c7u0cqrLP53fMLc+Gfs9QaxvRc
Wv99Bs+Jhbi4SeNLN+mhvO89uYqLRRaREbqeKeshNZlj3q9q+v8oW2+Fh8eghSGt
f32doMQpr6D3ZTxcHWr1ATRsq3leU6WhkuhELdiX3aKTA2JuNuptgylh98VHCt2D
3e5dukmklWQTNfGkwEFJ0I74vRW/n/4/0GRB45b9ZoIiTzCAYAkmvYsaqKV2QE5P
1GfOReuuEtc+Dzb4Fd3GBKErOTNbnG1LKa/1ObqumwE8Feco2TiXKgt2rwK0i404
aiDnoUTrBCnCCUZU0jJpZ+yVGn09Sy35ulsE1XbbUOXvME8h6xD5lpDliUx6IY3Z
26LyXNDx8CBdHr6dVXk3Q0dLj3ArOh8Adm949CbQ3ZUs5fPdkq4eJSDW0xhSUNkK
szr0ddky2a/uvXb5CyJJlAL5cb+x+oikyAeH5o12SqmQh9wtpYQ9CRAgTVLzMBmE
gxIlsbRsh59esNRTM7/3UchvUJoZsqjdFHS9HpKDqnHyBhcmNBchGs9sDAcfM2Tf
kt+OLWDWHR0X5Om6/TzjVLwyb5N+xM7ck4gCPKbVV9xQnvkH6VTtTS+sfZ+kj4cY
CALA2jNTMHfhgek3DqpvoRYLJD7hbXMtZcKMqDiLhGvVAS50ko24pwbfAQq6PjtO
6c+eWFVvnNDmzRWwKguksxRG39y9k5pnvc/Vd5P60ddXUzFPZm/8vcZxDKqCDMbD
R2V5ZvAXiacZBYzG09yz44vxFfwuneFpzNnKdCcezFEgIH7CU+BiPDn7M1lLNmSp
wrRU3bb9LTMDcjzUdjlpti+ixhJal5h1ngwfTfGm/ZYxts8W4lDc5YDCYYEBjeJI
jTPCj78ZhH8lQumNV0ipIUl2vIdF/ephVIsK8E5oI1AhrzD9WjjpszGVIx7Hw12z
/mVhtZNYp89lzQP0UpcbzH7mMGQtiHqySEk0Io81FK8iMRUJXWHTgYiCc61eu87L
aIbzbTx2QjrmcYtz+DtwVHGvNonIAM8flZqxYNbqOIhg0hx0G3aD+U0A7TDPFeaU
kAzdQZkLO0YhBLYQZ/jcNI+xH9kSTp9YAOhHDjjnO0uD4LqC8dZTVWijjOwojwpH
qWaHSIiMi24qU40OWhT6DPd2lXhiFp0PfgkC+4Xj8HkT32cgzhe855eDlWvt1Ye6
14q2g6ne13EVSLC3WZtg5WVYxB5bcTWytmuRBdfVtMmCCWF3ctazZPGCLmbyZIT4
3/F7QR4Dn3sSyxcXFUo+fPvwgXi5D8JOL9vJHC9gOMNu3CAylcYyMcRqLVeDtbSr
P6EST3pCL5D7X+C6Tjp3zcf67bqIc9dkzlvwi8OTQ6QkGwDQpDFB2kUlXje+Egva
2duuEhd5hfjqBNeqGsmyarNz1ZBriv/32ed9c7fPpfR9589CWqQvZZ8oRCSd/HPc
75sv+4d0BoejN6NMT4SXiN0yy3+mVwFbB4jQX8bOF+oQVN0djW7eILelUVkyYvlm
+Cfb9Vc1oniy0R3vLTNbUtkLivewF6FwNZMkiBGp2HZBd6U0W53LnJumWeuO47Oc
dtfnqJbr16QqYg6mJ+StZgb33FmBYQ6ERuD4DMvEn/4wwHgN91deXzoVovNnEOVe
5rwG07Zw2XRf0giWBB6YUg6E3EkzF53aqj9XXUuhzjX8bVc/UKgdRqrqK2I/Ri53
zdHaaW1ISyhINtj1MnpmDCLKacBxuJlrar3hRNFCL/ua0GdTeEHaF+OCNK9SQAMd
UQ5M+4Ezsc79H4nhuLi285GzhJLimvznMUFPe9aFKfFQJd/Dnnzti9/CH3t3cCRA
QMs++gcEYEWr2/YbMt3iMODb+AxM1t1rvXzdM/AebplQG/JG6kYrZdUbJxR6I33k
MP/PXcsU03F8BcBJH2GWn+0z4jCu8Ms4sjrxpNkmN89f9F0zjUjl1muQAE14/yje
PyufHXbXmf9AMAg0++/AW/LHBke0lKfTFLDfQorhTbYgPdmNhdo2AHcjBfJ/Qhjn
ld7oFK3KBHmz4jfkQnqbcMtnag0jqVwNaqxMSn1N5+mVn/X+zqV6rdqj9r1sI0RJ
F5zagTiDHiqXpopM9jSb4qRA+nLr6+R3loexa1MBbf0y4VF27NumppcboD50ai5c
+ex94zoahOI/m4jltLCRJjU/hXIubHI1Q3zNGLXJQ07S+meYeL4g38li0LRe6N2w
SUp28clbpDzfpshUxK7JfPfSRkokqU5Dueh+YBjKI69yWeK5mFrmaWrileNoJWdV
Wyygk7b8gsXXvc0VlrNdcQfuvNFM7pDm1+Y/Ke/WLmogXtHzR4TgdqviHSoBSsdc
+PsA1gnDu6ozWU6mdazRdYHIaWBo+bUV7+u2LKMce4gR4KgCSGoJfKBzZ/YPq2m9
ZXHv7fFUcnuzBV44dU1U7+6pqmYiQFU6sH4zXk9LsA0h92mfp95ecOaP10gGDrIY
9OUXlF+Rkdrh3yUswBFKkqkhdxUCs9kEbJoW7U7AQAcjzDWDXy32km0kCP6UAn39
IJXo9NFPYznfZwH/iLmJIKvmngcRtDamFOcd8r6k4Ny3ucWGfZNePzfhLYGpO26q
x1z9d53B2JXtC3Oj0j99aux40qz4n7qjLqt6izcrdXwzOfWbEEexhqMJ5jTnuQQm
G4myBzisWV56ydcpmL5VxMY+MqRj1TFAj+wCvpLJGJg/9mXHGC/bkSxITV4YZmTw
KocKj/95xapqndsXxa3/VcCsZGdiSV9K4wgk7gN42RV5rGnKIOlUB8uTtj/I89h8
+0my91pY3qD7WJ1/l2BK/nj4Qg0s1IWCCIRh7QZvXeomnaXwnkbwxQ/2vU3Bz/WC
iKBd5i4nJewrqypgIOF6wi/KhVROgHNtN1vQa0uh+vMPT58GdsjMpxmNWZmrKePa
kgiNdHAuNfu/N7vnFDerBdqyb5TaaUt65uIDwqrx599z1cqzNix/AhfNUbCzrUqo
c9rVkbNsU2+Vwd8kUroQ/Hglqbdi9kq221gBBLY1/gG74LT8wMnLmxDjyynVbDr7
q46vEv/qFAGtSM+PxypC2T2Yitu10p0AE+VbzAnRsLEYqlAVzKLPKr6rlk6lGCIa
+iHC1Qa8Hk04m45tBRuXGmmkt3blABbm6Meq78/8k7PeiQaZpwZWNSteA3VPBkmh
wRtTKu0fA/x+NDMD/erpJQNGgKnSN2OqOObheZ/TYj3JtphFZMJi5i26tSani3YR
SZ0idzO5Hnk47cPhs9ITsQP6wHdda8GZoDa+VwiWOtyG34gF1THOi3yOkN5gQ1TZ
I9yUoGXmCuMa0tMhkWXuq96nqMnooe3L/j3A5G8Y+8ur8539r8z3PSMZt4M93YC5
CJu6/MAq/LVWK0/CkKr/VU3W9Axm1gmizS76NDROJ5zJA8IZW2JRN/eP6gE/lEPm
/yjrOeHNx+QTJnAzX7Y9dsXydo69EFCCV5gGNHEVhNRJbc/wROfXYJHXSTc67F8d
QaDubhrz5abmamQr11nSkUHTpEK6fPl7SCoTtkmiJjyI5DK2R+S0GU/VvOZaEsAa
rSPEDtrze8wsOCoSqElNppKUM8mzdeE4oe5+Xzy3CDphQym60kla2X4n230uMOYS
h8P30uzLEWTLAtCn1J02BJDoh48cEvYaRIIxAkS7R1KHhDGeOv5vOKL0tpWXGblo
lCeX5jDf2JhMhZgQZR8gAvlxTN6EaOyDiRqs0kbDk8Ffz11OXlkAQflcJgtf4EYI
XJrS0+8jUPu+RScngKFrhwr/2RuMjW3WSbLQNmkJAUGOepXZclCIEphUCScqJMuz
Xg1xYOmw9tZR8pnKWTAyUftsKml69ICXoehiC/jlI/VxJHw3/OgySz1OfFJs1YIz
IXvdZWcfzTaMsMxqEfBJufBvj+tJ3AWgfq0u1OWU9IaRPCIQalsnfw954RRz3hSz
MJuxC5XZwWjHVgGKIb3eS6WYz4NYXGOEnp+C9fUosBzTb+FWDtxJli6kvOI84+dx
HvFf7DsnbpuY19q1Sj4H0RfgQiEhXqWLRV8eoszTBnSAdd3JUZYG935f6qnqd8wA
L3v0/jvuf6sO/d3nvf5cXbxYynCxUf1tkLtLREnfJ8yjazMEb+LJ1HNOjf8nV9Cc
m+WDDF3waqIARVUittme1My1+Lkb1gK2fuWMKa2XG5HJB5WKj/+mYDMHXO9nbkGh
s41HyG4jsPkrhQWGLDjsf/ols/K1AStocD9Zs11/WDwbzKtT0PjU+sQwX2v7kjVP
psZSk9K1UEzpI9Q2Q+vBL4A0mRfQ7BlSpRf/v4Kn3R2yss4G6ke0x20l0BuUezjd
SuhvxY0TuYI5MgN2q7jk8Cg41Jd5C+VewsFS3yxE87f9rNvBqSgWjYWdJcaolYQr
4mc31BgXZSB5vTkSvkAip4gMyltxHHOTSAGPN3VvzW3HSMAF8ERb4vkWZUlLCgjI
4xR9KOM+pyUKZ40AC/qnTcx3EO9ZRBTfYk4Lzww0Zf5cPz5ohmSJcyu2oyvzhfA3
4zrfUY0tG4BJgMEHp5tPMxExsjBIZUGL2duxe2zRWVaOitXcRqD+MRc6xfcymMz/
lt6MvFwMFw+6pa24KnF8BzesTG79z+DUO5SKo6C1U09nuw3jPlxB7ZtY3K8W/F7T
L4q/IX8S9qjDD3hL0QWACC2HKi4V377V0kVpxDKWnPHQlOy0aseL6c/msLfbv+MC
I7ney3ii4b2Sobcx2lIJKFM6bxfBK9800pBGDbIvBQx4qZCHwvTrsTYA76r93qAs
rnexigd8M//ToEDPc85re6L2T6Clxabz7lLpK3zJrp8vp6/kk2vDp3faxV8UYiH7
kWY6eDIgwv9j/C3QNJ3Qzzxckww24CekgJs5rsnUQnkhcptIXMtt0+CY2FS9aI+p
mJFJ9achIvC3y2OVYpbMxqtG/q4bSTkWcO1X+NVVw2dMmBrE0fnxzTJ6jeB+ZLxb
oCk597/0AM3yfrAhYZPX1CcHg8tgzMEcO7YwNRvHC4Fz4ZmA43cFKHczozZLBn90
KWdT/NAJhtQ+uSu4HNZmbBakh9cqh9B854jALeXjlFw/TvsGI9KlHLBqnZmx9RV6
EzsDBsZZ3Yw+aldBMHxOJiz5RuFVirBI7rEZVVSyRf0AOd3iXdAXW+H4wx7QrCkI
cYc38pkl3UxNeHBrqTJfKbEdXTRBf6CJp1hEqMZ9050/7Avysh2P5M9HboFVDfkX
snlOaEppiuwNl4cLXM1SpMc2e/lQkrOv6pO26ql15Xgprcvdnl1a/UUsqYV+kGYK
KM0g4UmdTiE6e+MtEuQbbbn/zDcwGXgLWIYXTaeOQDSLRE+9YaDCvppxl8jgSkhI
cV/BVm6qo1w1AUKqYBWMJWLdE7fslfcZHjrERgWLs5XZeCAEbLzk/Yt9gw4cjRIn
IuxEp53nILfS+UbBQvGXXJVjGSvSjQLMKqA3F727H6RjY7RYhJN9SP9pqo0i7wb3
WmeSPROFkymkBfXjOw+IOA7OclcXoqV7HnZqUrTc/RIpGoiBYjestiUveLfS71Uy
oMnQNlw66+nH8dA4PQ4C+w/ycjKn4x86e2RN4xZCwa/M69vPko7MGFUr8sTmKbbI
o3dYvmmwqcycnmsKAUdrly76WzWNIbgP7P+WH3A2tcMVWctBSoAzZmo09+8TGNti
9lgNTXixOdBceFTlhQHdzvBhnsPX0vtSlrw6ouyoiiL23O1yguxhvFyMXA4l2olG
567rJtk8aAxboQ2PJf6i2EHVcW6BI6LN8w6VSEIB6vRPsX8ZAhaewMOM7t3DltJ4
DaF+4TOHh1GZZsVMoMxISvbU5sEk6QooWoRmNtKZd404xCo8GQG3jFMWq7i3elgV
/kp6mgWP04dLKod/k+POoVcqTZS6XM6fTnQmH5n39JVpSvwfDwVsDuOC+e49RwxN
XkwKZgCuF0QO37qWZKHuiFMXxPeCXNo2GvPqRXVrjeXSys9h1KkGBv2xPzUHHXNm
tXif2g7D0RnFm8NxksihtqsNyT2QyKVmeqiy27KcZE5MpwA2f9EsDJwYpM2ydUUU
M24JX77Y93PmcaLwSWOnYk1nCCv8uuogO04hL0NEJQb00zfR4AVJ4Fl+I2dRk2MZ
wuM+8nCb46IM9Rvt+rpb+CXg3sOvytydH4ODeCIQF576hL1TvcqkpnBieiAmZGXh
eskd9xkGbSMJG8puQamCl6wyC5aFRaFTcvuo3uot8GiA+1nwyh/kjnGW09bjUhIo
K0ZjzjpGfIV+cN1I5gvVSB3FIuxbxddWHzEfsBpuAsdM1/PoIktaK6laXKFbuhRj
KVBLwFhlpofgGbT+RrDTbInYjoOHOQKhZrK51DjpzMXxx0we4vt2h5sJHViCGE7a
aPdw7ACbZDB1Ozv9rYv6rXgk2wz2/6fxBH+QRNm1o87zd3W+Nb5z0pzMm1LDjjLH
y7h/eHbp+E5IODpdFooQyeTVINvUokulmpowPEoGgIS6sgwuOzC8iUn0MLM56lnW
OA5bQ9s0cBWzTz82CMKhONpmnD3fA3ZYyqj3b8KFWwXWgSSSuHkbIUcq8KM585XU
/zNC+ltJQjSthynLe8kr1/rdE2+yU3AAYdXp5sybjtu3EhT574VXE/ModEJVusny
S5ej9llm0M+WAEFCIzmYe6St90fBWQi5IkZJcMej8X+7PEAA5fAC+sXDo4DIn7lg
fRM/DZaFxV6wIuaIM5A+iI3hlgBDBfJlHgLcU7RmgShBVYs2OFs+lQebJI+fO2f4
NAhuTw69qSPRTt9vD6SIPB1C/+nBZQ13tXh1rQy/lkVkgFN7XU+bkrJHJcr9qjG6
hI5lQFvPoWs6OkjluUE/Eip6paOYA0VYrkMR1Bryxz4PAKPMiWyw/q4bLRnmNMm/
PpFhhD6Zhkj+NsP5ORKns/66XpyXXEEWwoemASuZXsiVWCcBQZ+yitmkoOwOUCqd
mxZHSQojFk4zZrHwOISLHQBrcFwW02btO9KgIbwO0IueMtfxGHKd1tVaep5H6HH1
FpIEAEb/IjO0UGzzPCoe/dzDyGBcd9GTLY1ikA5QKBXE2IngIdIRKDO/epRbGZah
zwvN9hETT9OzwshCnvn2WstpK3rY5HyLLjbeBmCQxtFp1dUIdNYjjiZnakha/P5y
OXoD3Q097Jtzq2HTIf6LhATq0CtreU4DfWpW4WGlvBiG59MiYGhDudjbDNPKgdkT
P/MKogrQ0yHDQM9F9p5ZBhDiWSqTEcXBUWkVoiqUKn8/v/1rpNE3CNPnBULv4K2l
6DvsDnTbkSC1/EC3+gVKQAS3OwvncfTGjCon9jja6U9rbg7/SUN4PUzmJXYJbchY
BdiHD5K67rFaNUH/pMp/7VMgiLx3g+0O4SQWAK9tqkt55YJKfT6yyBMa+Jb5K4Gs
nXZqr06BMqd7lA8MJMYoBOPZOF/TZLbrYDkH6edLPM892LK7h8HP3D2TnO3zcaRz
safb+9RZW08KTk3LdGeX9PMwzGzDqcFcOCGb5ZuwBqd1YW+z4TZjr/GxTzNOTePk
hkyxvQzhLm55E/Zl3hVXucwGS6E7Obw8nv3KbG+SFjT/MwmKH++EtXB0D/zmNSvB
giIj6BDFGJK6+HsUUE7WkDLbxw5YN8GtatThXqTusHeCjMkZjrGyjviZDxYCNl3P
R//bZkMznfe1RJAPISPk77sefoHFefT4hd/i3WzFn9ctxoHxV0W2T6IQ1NUyTUZw
pY4LXLHNubBVjhU3LVaMsJtBYlHBBduRSh31Oo7Dw+jS2M5DwPBOnnmbbc7PJPw9
xlqayB/KgiUmsnnl2yhwnjNRRyUiI3uzQSeiqP+7FcSTIkqanYOCa3ddkNKvIJ35
8nk013fD6jpo+tPRPlZ4npEEfxx+12rIL1jUwnRamIi7yPa0/GzXSL2jY3Vi1kp9
v1lI5rCi87gHAXe616DkGqCj/nsNEg9a7cOykau6ju9orlZHkzrsKiOM1wFucIkG
E2x8CTdX/Gk1kTCKtad9ZZ6zMxPHviFEU0kl858LmuNCoKjceCGqsxu+zoWGDVSj
egxSt5Z4ixj656N5jhkTqi2X9L9YX/vcIxG9iAHdsyO2IoOyiaAqLJ3ibywT8IgU
P83c7AB8q/ItXrciIKGWHJ/GUS5km8kZ2IjK6IDRuhX1pmr63D1yofL7SqqGU8qx
JP5yue2EuUlPLpCoskb4HanFNwhaN4oBMfWYTqROXvwLjM/3srw8Os+NRTBpY0vr
iObUDnYT1L0BIy0+nXJGgikEFg0VqS6Oy5ZrnUJN6nVjoEn0No1yV26x3H9MmLBY
U76AqhqN2Mc/Lwz7lCUH1GXEx/QQgGI+Z9LoAlozQOGwQ2nhKoH7dpE7kcbNfxAc
pHrLfWASoBvCQztiQadsK3f3x/jv9DgetOdz/xMb3VvmgOJGpxNF+0TTWd1OX/cn
E6vXHFlEFgGL9jkc68YcdpCn9EYLMiu3jIaFU2YG/26w/qczXFU0Uz5dXp4xiAAz
PxyVnhTZwxJ5W9lR5JKAk9GR4/fK+8sTiqzjq8EZ0DZEVKjLt08O0Pz9F4xc/B6P
/OHOiy8uD3lYW5h3NaOVrY0YABMj/Q+69sWA6eEr5Rg1XU+484d54SLCoGBFFIDa
lQ9XE7eIWnFMVkKJzXzO5aDLEVRtGVik1SHKZ4LY8duekcQNuWVmmXE7MO7tqxNe
HCzND/APqT4Kd0Ey8sD8wH6Jzwiezvw8HJzPU3w9ADKuGOHFoGT6hJ/KCpU5DCks
5cNQ3eH0FdylMv2dogG+rkghVPxAwhYghgXr8TjldCmcoev9uGFcHz7lwu30AfJ+
nlLtVhzBDza9uWXnUFexwERW8mdCZBSrS/oyfer6SemBGE1H41X76kxkAP1S5BJL
znzmeR4oEkJhdcdnHhuZ+4CEuPt9iaQXLnwrqyDEovu7h81IyI+D2YhFP0+lT9OL
bhVNCuvgzjnMdOif+tJCl20SR+WQRcilOdoXAhwW7HTiWJGY/i27qUaintuFqcMv
xA/IQEeoiTJE0gSRA6XNZkCsgd+jAREhdFpvUAiPGHZMvgeY4ID7RwnykHbxRKLG
uYIlACyT4rnY4kwzu6jYlnNkS6Jd1xefB/0dib6hr8UMRcs4U9GDz/tVEFyR5pCE
NSowwRLucS6a3p+78paSJdgFELuTKYIn5/oN6KghXI71xHWsbJ8vvXJQGY1WUdBU
oeLUxiMiptUCfcc/SgSo+TAdFsQFyiv7qGNTgYuHTw99mxbjGKKfGJmS2kn1O8XF
W/HW6hThTfauhR/acBzcyMtyw629qHwAE+GQqbGkPbnQ52klRQObCLDQTbQotg8S
uFR1ZySkXRCw6FnBCzfh23Gjio66d+G1jdNYsMKF7pQ4yOQaXeq4yyK8QDItmucE
oOk9UZGPXb4WOaznDBWc9NiJyeStnIAfdDKxbVwRkWUQRuY2B8RyWEtcI9UgAc0J
+/wASGq21A9CGlQPE89r2KqWQ9voZ2iZe6AjM/S8yPDGxnfIO34gmZrU+E5JJ57U
hBeYHjUAjXbyhWeeasdtEbUexb+kv7+bXeG80Xu87y95TrDAtDZs4EIH0TvuyFtz
hqwVNrkDuoF1OyAGwnOiYauTc41x4pdM+yx5AlU6MnEq7sNKJWzFp9HFzrIrQOEP
xp3hUaAeyEUdcLDnm4mMfdro1CpinIQnElzDNa7Ty90/TPdElHGn1czFYM2faQTz
6hEu/4rOKi+jOZYleiiAa7PO1e0GjKYcgSAqGFD/OxzYw0oTncogdIoZN2dEyrkj
v7u3KaHWEMmXodpebB4/TsZZc6Ngvm0fA2PhbCb1Hvef55csZlDGMAyyLZ9iJh2F
WgDeWIRL2yC4jI+LwlRjdGXhtS99fIEn0CBAxhQjX3xALUiwmzIAQtSe6p7TswSM
tI6W0+eynfT0+4Ys5JsP1LExP0y/EIVg5IqqNRnSUWwGCBbhR5SVomRbw6tQxU7K
VBfQHsoKbqiw/c1cdEp3pyUSJmShjHSAQ0B+Jb2I2OQDNx7kU+SXnp8aJuPvCeR4
hF1x7iPrpQS6LfLocvPaB6LDHL8HsglDuVScqWo3WvKP0A4GZL/eJUmX8xdkE0Tv
se55W254RhCUobD3fMcR+GQ9oMsMCDploQWG1FGeFXoHBBHCCXLymXl+QZxnCF2q
huNZ7ZS0nNosJHCFoJxbtCwowNbtoRcGNSA3vkkjyjgXuzLWzJa70xtMT48VdBvL
C45uELQOyAtfWkeMCtfBBZygGalIytJY7DMXyVmIuTD9TifKg8rZxYxgEv0NNpb1
E62m88wsrHzF8efpXg/zevm9oReCyMAgVkPDgg6Q1xYIwpFM8b4ATNfTH4xwoisq
4TRQBZfa2EnuETzkd817pZdE5j1mZ9L5aiYEAWr4W6DkL5q8YIT0umSienps/eVx
AvTEd37wogTRAWaUksl0Qc6zSpYutMq4kBcXX9jMD2RS+nurOYZRHiz06hEPF1vm
cIYii5Cng9HdJNCs6aJjKVxeHFGnUGd4Ze4Fl/2IkqBGH4fvxSglvVOdhv5On8VW
6bbZv1aFWOFH2lTj971OqlYiwUvgDUto6Ih0a3l4LrxI7IAtsa+XWD3jrW7ihBIC
RCXwv5IUG9kfeSvcevJQ345c5fjxwR+IjfINDpVs49BGnQ7FW9dcZtkeae3DFQIi
54iup5sfzfsLmazdsEWnaOoYqFkOvpUBmBZIQdEdHo8s8/fBDd8PNFdqswM2//np
IdEBzd/9tC+9FLc5+pBZczAP3HnxhkczOKK/N0+Ie2/w/z5Ib6E9Nam2HH7zpCMx
cAxhmukKD3wFFokhkdDP+3hRh+RbtCfbvp0jLsRmJlkfzAgH4pj+7XDm2oUledLN
6f2LTIjk1COCUKXv6BxKab2H49Juyk1xCYNI4DUJ6fuI7CG9rHVrEoM1OIcfbHve
idIjJjI5gffPcYm7oc5HsWIs/RI+2Y6YVK+jiMJC9419w5a/9Z5IDjEm49uV16++
KZiKzC32JTYv4bkCwZGvN3Axzt1bmR9v8Hkzg1/CSKjuhBoySKjzI95AEqevW7gr
cQd4x3gmr3AXWlUJVKMR+mhWbe7TLGhS6Qn/r29PbwT4il8oMM4oaUsjuMpYsblo
xSFfZ5KKcbUccayI6kdq1b1DWq73mPAJhMzMedYmbPo7piaTPB1Bys18Nx0xjA8E
2okMdXsZ0mPgjv8ypLBgcOdXX4M48laVWazRHihIresTAc3F3TnDmqyC5WWiJUy1
zXOQ/0TjKr4RadiEQj8UCDeIU0IuhJ7O6GTGnpy24VFbjw9LKx9qeA/aAPhdoTL9
8vnKou6QesiqfyWS9tsTrLSBXAibLikJhFVrLnjmuMaj03Yrv1jS+GZI9vNjAFyt
x10GuijJoEbPu583F/UzIY3F8L2NBA3MkKzNtSRvMFsAuW63ZUFiQ/0kCDmBdAAG
DNun3uSO5fw3819vwbGc5Hs7afuAjx6wRC8b21GBR5q87tWB9vbNyuwoHopj+6Xl
DQrZcBUc/ztc2RE+EWLtfiw09TqQtM68+xQIbd2ZFpUTBsPgJ8Z4aARmzuuwZD0k
aYM9e7RZUZBEv3eQTAG7fpE55eMHLQ0oqck561pmkQP2lh5oyxgulj5m10hFkoMO
uUWMuoEyNRxjLiXSV4nu//B1fTcnpQ1/cVD3dJsuUp18mtcWQDG0KubLyh3Mmk5h
zRam5GLjmJyNoxsOQbbiNHquonmL5ZlDBiIo366dpdPs128JOzAwf4ckpBlcRstx
5yEL9HJ/Gcvc+ZoVB4PeMuPpTK/qwIY7+FQ3EzCXMxXc5lRpqmP/i+nytIT5/3+h
NQwtSenFdOyoGS6UJWYwIycWW6u1k354cvrHu5hdBVy7hbaZ/u1hzulR9xwMlLoL
4og+iO3JnttKxxmP1Ak/r/tmfo0q+SsXt/dmv1szzTyVFN34IZ67P5pksSicsDXg
vA3RvZwxQCKFKZuqTW9dGPL0VAB6qITJyQnh/uy6OQl3ykulIQugAs0vOd6fTUvT
S8Na+aMHVG0EwN36MvJNpynhQWKLh27k+MZ27E4tLUhmFU5k3V24HJjzUqWxKUVy
oPZ50NQmO4WpKBJ8BsT1Vvl0/wnZ1/aA0yltLGwxBcFWF+ToqSHsnciWmtjy8RS9
CTta64e80S2pPihlXTiDgpp1d1sibQzNklK/2Q8VFhNbkPR9vyV8vWhnk4keZ5Xl
gvDavjM68Nza+xmFVJb5DNGARFbritDANiYDl5ywYaU8m60ckp0Hew5bXR9Tjb3h
/D65DYTYpxx/oEVH2bKhWwp96AQF8uiqnQjsB81QTnM4piuDGcmhkhcXvB/d5H+Z
wgVl1kMy4R4bhlwUSJFZNzdVXgzb9JzzQXcg4wIm0VSGSVygN6Uik0R+ndjWlv2G
rJMwVleZHI4Xqmunk07q6x7u/bIjfoi5kbr4yppUYYFMKSb9sIbgFAXhZD5MhfPs
lWSNDQ1hOC1W3Y4VVFbJq/c/W9tVKWTm8GBk9sydUusO6K2KUsjCepTJ5WMvVM4A
u0EQFcNibvB/pIzgHuiNVWXU49OSEM6QoL+iwkwOh73eR/JeNsxXLTW7etQjP4Vs
LDvf+qJ1X2ubNDKpOoJDYEtTKe+VHx0tNvSTbfZ8PzEMzJwssz6lLumM9yTI2fgU
7Az8KpIKmUYjKjlnhL103fuLnaBPEMLKzUbn9d6xnzlHyGJO/qKzfSDCLo81MX3d
cxdtdDu5QJbpRSQr8HjzokfeDMmps3ukR9AS/rwj8b5LpaviR4Xkt9YfdehryrcK
DDmt+cNgUeeCI6jOGBepDtcT03Qrd/im69C715nNUHGxWp0gJ9q/tk3MzGPmnrS5
DhSBRdh8JDM2FGEs0zPwG5b1BnljqnK3O9mZfRdN54mDOvDKN3+RWQ/+V28ym2Ox
9zF98ZZQR2X98spLfG0pBabNO2mCL8eyuTyfcDG0KqUsPbzjsJLLtAmKrk2ue/Rv
AezsZP4sn9Niw7hJnXCGLjsB/m4GC2ctK9HAT5ATHofMt3nz2Ve299Sh2Qn8i3Bk
PnICJPPAdG4S+lU6bR5sxLfFXezDcPmX+NRzPuLhO/8WyY3NFMNGiPy43aKKd+eK
cbBrkU6MaxXTgxKj5iktEp7d7Vuvt4S3ODdigQsh9Pwm5Orfy68oOn7oqCMo0Z1o
/rjc5iWDm+u4TLUV2S8jhUrD2oXCCYBw6TszGpu0UNWsqFFb0vZCq1XuNgkLRWcF
3juNA7E6neQTS+WyXKJNoH8ysXbOH/j/beGODnvU7JeZKD23ONieR2/hRYpWq2lV
rRL44b2TdFh9seiN9LF1hd0XruzVENsQGBivNeG8ewR7wRudz1yaoRKDzWUMwgjD
iXgHTZVwcleMvFR6czmwmyVNLRP4plxfJewUAKXqO4h04SW40S9dPLtl7Aa1+MgX
GvskRYak64zaC0d+73FQcWBfoe4FFRDEVYcxjmtl2ubJkrgwOJExfB2WwuBlQnIi
JyYHzG23ll2w7N0gLgEivTOerV4mp9P6jL6Apial5S7P813PRvKmSeGdQYPo7rHh
DwujCrlZO8p0pKzVJhuPEN7yUI7yrx8ap2axMr5uSBg7+arZibOuv2e+9hou3+GI
RuOtKGQvanLa2r+Oyt5PiNt8KZR70tY0b0c0cYwxdpiVQFiHJ4EZ7QQSjWy3M0sa
KagxIMqbPx7ZY8+CgqMCl2tg4Hb5vM5vIamLxqwX4HPQAxlkT5++qiHdR347g6lE
lsIfp+YuKQjjWUN0dDYds1m9FDPRl0ZKBAyKLGvYeF0CljJ9jndl2oB7oemC+QV2
EkEfYjv2Wkc5mvS+sGO4d6XgKB/SmrXmTAJdsJ3OjX8Kz1acCMmkUMiiPtANNNrw
EKfjzzIL7rs7J9cdJtqQVQHggwi669oyv1xKohk0dmuXX/MhEDIsJoKQdAGWphHW
fqpzihB7UOw8kz80+VqVt7EIKkhm5+/OcDoI6qfqJAKdiRjO+9Z/Iy/uAWU027DZ
CXqtXTWZbTLSADZiS3TEiMHJtlYxhSXwXdSq48GnJV6NDifLJoKG8W3lRjJHpzCF
V6VvinKpwvPWzgfa67TuyOyo5QhyonJc/E8e3EqwNN1htLHxCxi0+X0d6AZPLL3a
h59BP8rXzYqEZqItE1d4PhDc5gAWHKnBEWTzqPgLgkORdX8tmf4dFRENUMvX9tTE
nH7uUjwp/ptE5pdtOr3mW5V44yfJCDGiMpsiWoQyD39c17mCmZNMxTfSWiVL8Z6h
gW/FGKjOmhSui7sazlCOILCnkZB6SRAy+L8ULJ4k+xFDm5xuKqLr67mUdtSi680e
ZddDwtc6RJEcVAF30y1YXDTusu8S73ThkHT/9KlXeVs5jDfhcf5zIl1udizORUus
q229JOM/59k3QtvGuP58qObELDiZNYHMuLSqgLGk9APm4yWY5TqKffGxDulExvsf
k8bN7iU0xY1A360kzTVS9OcE36LhoF25UVjg961pd8BAeFLksaj8zkEGX94AK/EZ
QJ4pWvfx4llRsLJ4+XjBLfAsRJkbUnGBGK6O7E/QawT8PL1CIKC7hCM367qAT/Fq
nU+T+TEN/po0XxqoUeJArRTCP+R/rVB0wEFriDh/+6ZyTxMnGaDgW9rojkD729kB
KuWBLe89vlyEED5vIR/M5/N1Ms1nzyT7b+dV/KVE7GGLuKQqRhWAjO3QAO7OB3um
/RopGQa2DOr6Dxo/r/2+3Yb6R/0klRynUiFV7/MgXNvby8tuqI49iCJi9fRqDCF1
+LYfymH+XgigPm4fzN9+oiRMaz3jE0yo4/yEGLer9fZVtktQIODExzUQQqmivh62
w0HGx3sKV8Qn1IZixsxeWkA0hJpJYMv4ltvVl8PMpRHz/PTfSoATi29H/EJK2QD3
CIPgdjngMqZaEV/dqoftqJNyoFcUZcppXyqrBr8OEy6dK2+aHGX8ruPgI2a56h54
Vuhf8B4pk3EpqwEh5DMQxmyeVaeBTShNU0LDvLfAzgPzDgWCr5TjUU78uA7BwKvG
ZLxoFZ7M+tvoBb7KOAan1M4BdGSJjM8WjVRM3ETQODLa1oLZ8TA7YBK7ryIR3otu
LCDjZIE/cu37QpG+o0ziJbhufWPncMZ89qT/+p8l7GyetkiGF1DrG2q237cmCWIl
iKqZ/t0RuNq8uMvW/ol16Qv03UdKpQ4Lalq5FgB09dpv3RmuvLaPNClZkwLzSG5M
kxR5fwoLFIMj7pVdRj68Nz6v49xcdHRVGbBGNnq84FhVrN3Q5Qb+C8canLP8W5zy
+kSKkQolSoXIrTn5dWPhLkK0j5wTbNC6jU5oBuSnJq9WPoki02p9nC3C0oXZXfUC
oqeAzjQTlbR9PjQFgDTPEdbI4nCtOD77lek3gFBuW8YHoRo7kMjKio7nBb7NGS8w
YRzM3RYGrupDDkpYS/IeiqTBMDj8WIKef/T8fAiz4sK3eCCwwZ80XVNOQfucGMeZ
HmOMPrXjyVV5S83iOQkwzoD8kDHbPUhrIofwmM8ESoz96PXdy9GkNHvJ1K3JLCjD
kF2n8LdrSn4FvADAcCBICR5TfxppVpIhRUCSASwIYa9yxpMTij9hZvX08lrWDgw+
xGdMsRmg6ca66Y/Z0sG3TYYEQvjoCpKwH607DZ+tm5AcQRzW6voXAgQoZR2l6sGO
IqmGsF+DCLuUiolfQmxxj++YZeVREFHOstZD//7oPqx1OLAoKWWe7kpRqxRwvtrD
7c1vyIFj+ORu2jXjOa5Gh+h8BEeMGhDcjog2LNQi1S4vgTHN1eVe73EqpPNw5JKU
cNLC3mIRSh30wWOKiFMUV+j7LJwFldsfKfDGCA5h81OzjguHIL/lWVIp1nkJrsWX
9mZblRFEIy9KTw872s00yuofqrDIvIO3HYsOgOwi68/Hx/RChnN2l1YGprnp7Q/E
XArCdNS09odphnufwD787vtGJnU4QYa5pVMCHWF8MYFVqsQXa4kLst700VSdpBhA
MBDxw/xR76KRLFV5M9H0AxukNeG9DuNiawhb8pDXOjCpr83qnx0UBjbtscFJnMs7
QN0rwf5IXaWzvks6FkD5s+EGU/aAFzRWwOJcr844VWNXuo4NFnvL57arj1IpqjQy
39YexaHeoUTskdHAJmeEYO0XY4Lyoq7pYBFI5PqAmYDDmLNUHKP3cPpkM1Wez+xW
4crM9oCkKuDpBvfdb0WpzS0RBC1NzMq4OUFKnfSGP8FBdcJ6MMeHi9g+swlMm6xm
NITwYprPKXTPDeQzOr9RxCZECP3b7gJJfmyOTRZZhIFpVAvzxPSTLm7LRA+Idd/K
pvYwhj8a/I8zaSyp0cJxhvFgtVrVC5ZsIR8N72cmXPglK5z0dnSP3JsYh9UhfnWX
w6icNv4n7xMvSgPEeIOEFxQrsiSddvCIo1UmYOQG0NpT7VtoXBgIKZurvf3qRcbo
9M2jP5gQCKtkwSjQIH1HnGBrha5Cl5xYDSs1J3KSR0cR1FS3MoCygptEA9hhPP4h
dpjqioaIJx4nDlFVk7lY9eXHxDsIKdlaJ+XPpAWCXtipKdwfg+8vYa1chqeqAJUT
mp6pasHR1I/jH/vhmsTKI5kgtXoG/mgawK5MpwiYGWg9P4I6vSeNKRH27J6cXVYF
UyzQMU+n6sjr3VdqjFntINbtr+hoNw1AvqQLYzc2SJCU9UY1xPk+L7FiLhbCXYeq
CjErcOOXegbCZCIxm7Ax0k4q+sbwkXG+4dfOILlbrvQqCzoJPnvbg09cZvkx570r
/7WEjmS7Uhzjl/piswAyxsOC+4jiXikdIuhmqIxj9BzSE3e/3YcvhLGZOv4sM0NK
iGFLu04968uHHO9Xu0lJ0egdwhdjoW/r42go4MLhwQaRNP200cRPBZKDnA6AQY5D
qnQUwZ1siU+/q7BoZGELTzwSQ5q02QcINd3wRlm2lxCGKwdXIJaLT/A51wVc0WRA
HfBXQUrnXVptts7Ol8KT5kqTW2A1rRIpuQCNHnO4DPiAHf1VVz4LFTOh8qayhBy4
eSAC4UYJXBztDpLfnZES1Qx2bhXRTyU/Ya/3y5xDLZnIkikGt1cU3SQZwWkbLgjc
RxYBhkFLUcDQSwfqyaatvbHXYsqM3d9fCxe+sGYQzONYl1GCxmoXNNairInrwhN+
roukXc8xJWS8Z+5VseFq2p8dukKVHCy2Dc3gPB+rlvnuNPy8edlHZya0M/7R4ZXO
RhzpuzirjOwNZhgH3BtS48ocY78Vz60r1fphAfaTg7Yrrst61/7iRosFqdrCKOCC
WZFWBOEdYQeVn2VY2HZLuQRvmFiVxVs3bLivrrUjAHR1Xk5f6EtMS5HHs51ZfGNm
KP2x5K9URb1ANAzdM2zcovFR0n6qXqNTab1Q77FGcn9grO+KyEH/n0M6RRJZYdPI
bNg3R/kXHSnUSbJAMAbxT8YPpo6x7Z9jH9H0h9SgaVstQlOgUW/84miZqnvAUS1t
r7jUOXZ4cdnZcOCaD11TxvUFPShwCTyd+oiM9hsEkclStv74XZdfslPN0YJIT+ZI
1ul4GDk8G5Aj8GDzBM+CnrLq5cuKuoBSoDZTRVUb6spVffbcXSWyGqwa6n07vXgF
XVBxvxY3AzQb1uOxrClChxNXHiKgrDryA04fhjILQo6tQxDMjQSC+FK//TgCnHbz
xBdMqdDkFmfu9NzIdM6h0GrsaRvZSemCgZ/hAF1lSDqcIL+JR7Q7WRGFjfYsTVme
UFdUHW5dAiQi0TyO09I7Uug63fMf9Aj4nz/Eey1mqsZpyNEwl0RjFj+buS1EkvK6
EHzYy2ck9IYE+NfD6CydrHR4gnqul3CpGPRff37Dwdx0cIl/JGFFEVTHIhJeqbE0
zW0r5a0cp46i+iW6DXtzpDPT3s8dT1dT7cvPxN0HlhERYLsz2saANO3KZmFHzgzK
AdKVVaSDwfT2edpHFwdIOIMqrLhQGpWoTkF/Bk4rdg0j3eteldhL2BHxs+KfHsIK
5WvuWZO0cxEGYETu1LtVNdXu5cmHs1rdG5ZD3bWN6Jq8ieziO72s6xnjKmnM1EhE
FAMSOo1t1lT42UruLFp2Krk7lKodIcgi48Q8VLLYSdQWBoAJ2hsUijPRcx3TUl11
XLycE7CtzFZsiOBkOSCDYh+87MARNoQBRKQdIIorfD05K0e1qKUNsDiPdeqSr3s7
5ltXt64C3i3VgclLDMr4Q0VhELbTO9bZcLTLnxctK2GGVc3yixyE67ITSXW+P67j
a8kEp7mKINaAbK1iTWIXe0mKN3AOmx4Sg0REiO9OLpjttgodJTk8s82kHbqOUQ2n
cm4l/E3HRG0DVJhawdC8+PlmrQrCCEqU/tmlQm10QYL3JATbVAXuV7kEHpmmlHDE
3bMM7f1IjJFNkzdI4pwd7UbDzfHsznM1p0mdl9JiCbsjBIOVPmxiqrmSLx1h0zxt
vuQeAHYy2SfkAFaEmvc9sv4MGpZxJMgN0c0FsC6gCzML/EfkJrQNdWupBcZxeixD
rIVqA8/1pYH0mIb01g343TQNjK5CnRBqx7RVY9y6TcKGRWA0Ice8/iCPHeBkRFDj
7NceZkF2BBHZB+D8/rttsv7taITmvT3Yo28jxEuvV3/6SvsTyDePz296737mHHig
+PmR5Jf9FPAHilPJnCss4QqQeb150rA3B+VekSbavf03KEEdGqXQ8wBEPEqxs2F6
oHJeq5yIt3W9Yr4YcCPzAVA4DICnolAfhIMX2kasnbeEXYuvOewlh+dFAbpD2yYT
UKque0986aeLVyUicBPqhw6V2kyXgbnitPT/5CyYP1HwpB0KwHjLpNvxUNdo317+
4V+D1e7DFBiCpoVws4IvP3pJl9lv/xsiHsf4qPMJbSED9EBuAxbokMQuCjdruO1/
Q3f+SfKQR+G6PkyrztCMZLCYEvBm0zOV67ssdHzDJNo72ifhC8Lrwk6rfOVbNocw
0KgezEkg1+adXBdBpsG3zDY3dvTS2TfpAB9B0kBbcdOOzzlwcrlYsrRoXWWmn0PW
DXpcTIBvZdP33D91EgmZ/nTiMyTjosfjSa7FErNZjpTiCB0yS9jUWcv4+IeFEwNG
lgOldwe0WMW0qckiH6xhBNGrPBFiukqNiiAEc22uVNYBGlOskMsZgF+nIvtLjckQ
NvpGzzu7Zr4KbvdLQ9U7K1hZlVjAFhSfLYvytMNpVs1C3Tjxa+7VANm9U4idlrwy
7K9DS0/w4QsXUnL0ZJvuf5dRprNe4Z/crJ6OV+Pm8HK5b94uJVzKQYzvXjGclC2v
i8EJCakWaVtjfRqx8VYeA9Y7MJTktf/cRqQUyLgU7z6usRapGqxuOzF5j2PgA94+
eSklvHKzWPgJvDt69gxqudzvNN5HDMNCaBlsehrFtbwOlAZg1a7YubWYOKT+Qpap
N0v3wDBbo4xvsyDQXXunG4QW251H7dOT/1C9TqcpuRM+8p1GKnUsFytQNFqyBKA4
lZBrzwaXsBoda2ZdT9y5r6Y5E66bxfIVmFCjrbwKG8WlbABYFEPNmhDV5wohTf0J
kGC2do/mAP2WocyVv+dU+5s/FtW+3hHIDRTASTULp0EU6lAA66uvwzF+G1Ym4vyO
SzjlSgg0cjkAErWRqBu1AwNcAdTvg+S+ctYwYzmD/hQGqJSs4OW02c9nkGicMD0W
PBqne160GwBgCNOt6LwQdsf0Ftlkp5kGO7WXLmDtEwoEmLo9eC5lscmR6Cfym/En
WKLuqQ8Vj7t0hMMhmrWy33Bo+16HTK12n0Y5YQWfcsth77E5VCzjcsb42PSghSnK
WFVZaSPnNDEBjnpv7queEXyJjtHpb4g4gRg339lvDAXr6SR+mKxpQk2BsLX3yt/z
IHp8Ur2kshP35CiPNDGLVHyGhmsGnb6vgw5iSWOrblvGLR2iHmrHfEIhlB08HXTA
9ayCPvHXCQ99hnNcX7aHQ4N7y6Er2m/5U+P9zEEx3N4VLJ+1gOFasFML8fEvOms8
Y5lH57ALFuQHRGCPBz1C862rHPeSHotfP/ILopstOM4mRfGR4NX/gB3D7G64Zq41
y5CohD0arO0O+rIFPXRbP3FhvKYGBJjgfU1Ni1dbBsxvVCplARqFifQzmcaavmM6
tMa7fNF8ZyB18Ef6h1bSE/DaDyBbzqPedfEguh7Z46jv24ZzDdWZgcdFoeZTSDkG
Slxd0zViiyLzjDaTf/Sc/FHrahdz3iZI0b1/ilWhQ2oCOrVf5sOknNtiJNfXiUvn
NjYMKvHEY7hzJRiwITh0+ZEGlHEGzAKaArNgiwl5jdQfmBLzSV1F5TQGHObvI6Zv
U6kn6dZmup0Iw/8CrLcyt4l0csfBzalHuFcnwnUjcPpo7q4KFBJTiGWgeXAU0UyL
GgyYEBmYa5hSTyRj3KneIsjtlGzF+nWPe4AlRY3aVjM4PEc60AcjUtI4NQT8f4Zp
f9ugbyVhAwAxKwWOcvrdRCUqCWX6PtZrBtGpVcYhtSNMVNP2nfynwYX23BVW4lUb
c72omAildre08k5KLONva6v7QSlaKlwE5EOdCR7DUUFlEVdYJPkV9VX5Gq1sda1H
TcXWRqsga1FX5l+TLQ3IxJz04M+K4jQdBsnEk8zGykhc0fMUC3lc2CAkkw7hLNS5
ZIyYdR44weRQNZ+ooS/Ftwb+NP/9JrseuCrERLg6dQs8ZIqG4sFRlNU7+ILtuUIG
P1v7o8pDrgaYLvQoUK3aoFd9oScSlzFyVi4j1aVbiOHRE6QqywBmaQ/83pfSjEMh
sNa8brYoW5kKDQqDCFOXKetHa+ffN37lx+xm6pQw9NJZFrpu9bqkZKmTujpXQucN
plbtWAefbBCrHkOMFLRTplIz9DcKNymUhfd4Uh7ME2EVuuIMtWSCiAg5LQu6r0/Y
iPiWvZ+I0J1PKQxdcuZZLll1EKWY98FqyeGHNL8SvbTO/uvFKwmuoMpjL7q4CUln
ukCimD5OTftx75OxG5/bpA2dG66sgmu2LiuruusRwEeP53gQIOnFt090cJiUynFk
L3wohMkhwc7Urf/ShlCtFYmQ6VSM2uhNfraCnQ9qWv2b64MgALeXezaZSrM5CTSi
X1EhbJ37JOXh5hzXn4iZjopfNM7x3YaKe/7JQIqcjCJM07QSas9c+DTYNGMzb39v
uBNyhoUE3FX71HEmaiR7RSKcVvHG6zzFahBjT0GASC00nNz9QcdktOjfXx/zVmMX
rotJarz9o2yYGwkbU9LmxOfDhf6JKJoi8wnmr95ZPxEEPk9tWIeH8fab4B3mxRZP
Qa0hXNSq6PXT8tYIBbsd+tguy4X9RadWi/kWluS3zhC7Q2U3Qava5+6sr5h4ZMZC
yA2ztMhVqZVWEw1js1wEg5uiuljZgi4J7Bl89cmFknlZxLa98yMPYQxMbWOyGEB/
PHIU/xHeUmSOYHKl++hqvTI1lij8xPWxXfwnhkFJa7d3POwi0v3J/egNtRcq57fp
V3dH5Cesf8/yVAfci08q2Sj3ESUraAEvYHE7nG8L+XUy4ErkzQoUIU1Z9dLgCLZh
moLf2dV/L+0wP5wvChoeHyFLg7tFn73j6FHjnSly/xD16v5zJwIpfmLd1RZQF2AP
2M0F5oIa2RcfUS/F4qPvwWBNFa1V1uF2KvkJyiRmoaIja2CpsnQ51w2/DpJ2pAkE
oU4jr4j+dGz+DpCZ6xhuuNdfcouwJnze352lC/bBMK2/mLzeNYuJ8XVRJ0uzt+G3
yvGW/L9VQL+wxbAkkfUDl1ROSETTwmSvQFoReUU2u83ec8xovdTDhWlctcnAy+4G
WvwVGm41d9ofYx+cQ+1x21eUiaAImEVEFpTXIvqjK4tej+QRAQjIuUXuiq1OBCDO
8qv0MCqPCYnocCnetM+/+3ctrr0cs9cyoBimYgyiWoZlg6ffDW7oL9aTwbajgML2
U28/Zmx6728RT2IjzDCJoc7Mu6P+uOo+31FByrGqA1L5LUKncO9VrYoVjnURO8iq
B7kbQzuc4Tpuj1/dmJTRDLSsueQZHPBS+qnuv8o/odb+bSAigdanfLQwg/FMjVo3
Wqqoe3xQSzs51kmN2aw8wQyIlhowtDtKoUmjzplYHtHBr/XNCjwKVShR4Q5dtL7F
BhUu8e5bo2cQhVDkP3tPYAYJCRvWiBLWmQ4ymWjkpl02hixDScXhdzaIUIyGFxDN
T1t/QPS9qvYQxJs++m+vHY0uiUmcL8rH1Hr3qVjYSFMYHKsJDN7l+XcgzR/pN7LK
8uQ44wLHOdhMa18M5BGJC1UMunTEgrdpjGKluoGVm/oP2LoLq9onN3dVJYV8s6un
xyZNUJYzk1SYCBu/c6ORC/9F/Jxyt7V2MFWKMxQcMijoz/lsUaoy1vUUEKKnJyFZ
u1fxKJVjPfiPex0dtJMIp9o75HGCoITQozGd/cQK1WNWOrH0oJFpzLA9F3Jbk597
Wy1cbgO2irlRgoOnwEDZKe5TVozKPOr1alUubujRxwJvtzuEecDiuo/EGxG3iAgR
PF0hKIl+80N0E435mKzF8/4zfiiNA67jxeM7rRYi5WdgvF6sjCpMjSF+iFGd0uq0
n3cYE/mGirWCjU3qDfqFY7jgSC1gt17kU6QBztur5zSDeYnLmHEMuxeRLEKOk4UT
T82+kDYUoH/3tYpWoZQ98h0LHO6tZWQzxzkui0bRozdqPlQfAP0K+dlJYU3TP1MN
SgNbkyNeQMukgk5Nv9KL8MCwlj/S+TpG9E5XDP/UUJhbE028ur+kSmO1bgpAcDo6
YwJqvIFu3bIdOEHsKBJgR7vdFl0obz1NJQn5Fn3LnI3D440gPwNK1l8f38VzdWRp
ff5OhTuNsafTLMGhc+CKRWmJXJsHtNzHc9LIuhTw5YU9MuyCGm/QQzNm3SKxJ7du
pw1PwiaJzFeTyC6Shs2wY6sNpaPZDRAibUvplDMOU0Crc96XwPySmthfhmx7WsYk
Je6ySlRggqq8YxZpRhJN5i/cIrKqJNFiFG5/OopHDWZo2ls8jDaq1ft8c/nlaKQe
cRQqurkl63xq92u+BM5k5xqMLjja6wMxLOAqMYPU0O2inSkvOvWpkXtQVAEOMC8r
Vzxn5OAvex/X2hsKIrlO0FoNd72ZogD8YxxU51MSlkF708VLVNGQq0jT8eH4YbFU
wy5C0AlRwUmEuQwO+RSY72R0ri8lq475YOcCsC7KNllpvzD0VF/VeuKZsJLQNvbQ
64aXDEUlXoXcmBWxL+ZMHVSS959U9YlkQB6+aqFEwAF+k9KEKssr5cSqRZrPQ8nR
4uCeENT1IQxmHaZVXnRra0nIS37tUidBJOQLORQq8KTiaH8mjkm6KkMC9XCbORUv
jDhyU5I8DwQ+Sm0JzXF2uSPg1GmNFAfdGw+W46u7I3IcCci2PTsqFoQ8a4fH7zZh
lLvtLgB0noaeLozQTl8UXhM/YhZK4IB31W7Ues2nh5hv8JqREbYpO0UV5NYiOCMi
2u1CR9w5hJKd2OAWz5bJBL+TxRKZnB0KnKHkgYssLktMKEvQFbZcJi+ybz9SYT5A
nnKOVhZeg0sy5Gpejtwarj1aep3556AEgbFQn/1TdrsNIb0UX99f9A5eOq6oYtVQ
xua21+n6ZYPxdnip/m2fLlXKjZTaR/b7NSwZgy+a2hyyG2wB/zOGIMx6ike1AEHu
osakK727CxaNwjuh1dC9eX5n4fxIiUiGI7rb5K36ccC5v8iN06LeFBE+A+Byo+8e
s3y8Ks7+ImS6DX3DEHPM1BJz/RyKhAsp6xRjQm65zlwH75thkBs8ePEx9WjHFEof
iCIJwAjTCJhBMMPISc0G04i/Z/QZQ5TbgbcEwyM+KsBC+uBkLm0Yzu3oF4bpkubR
cnn9/Kfr+O/RQviFDQc33u/oo4Ol/iwKbeIw7NrGDsCVVhwqv5+TbF6OzbjWAxbP
MbcA6GNeM1kp0nccGKT9Fvf7Gufa1gqx5wp53IFU5+fbXLgENPIwsIzcsP499xQd
f8s3dhh2xBvHTNMLJCMwEvhguH8CDzx57eTuA3GO293Jls0yYxlgrqSDagRKaIJk
X1Hmyk5V6RYAiU0wT7hxjA5vZrFBsDNkn5Gi3cq86Q2Sj3Isaula5PZbqWzsT7am
B57rPzqv4p3QxU4kceocgS2eykZEUgdxYWJs4OuTcSeHkPQ8nXNeDu3Kr4Ni72SO
aL/H1nvy9cTJltIbORl05BnGsSnokXRRb/UuT+gU0xTOGO9dv94GnCm23f7H4oZ3
5OwPVMftn+ytaCiEfyVODmnG9xq3PsawC2z5Kh8fpxVtfSpuinmafTnv9kc09TBk
4h0FbX3SlkvKog4AEl+fi8iSpVeS5jKOqg+GGX3dzUG7KCOWzBIYEE4vdhFjRdER
wH75SM+yh5O5C7pmrZk5XTBzEg5ejBd70S6JqO4QN74jf/r5S7e1QGJ5Ufw4tjx+
r4jz0RNo6EVB2KMuQg3+NO7uDogvGx/ENW16YuWR9h63Scclj06z05kDQqxRqlv6
E049wMKlDjwyIVRxCtAVWTS9qKME+Yby/3bc/ERG1tCJUQgxSNKoUGVdvyojl4KH
dDT8ixG1EYl3w2BOgIAkKhlsRI8juQEcxfen11O4AUDvCcTT+nfAgldtrZGk7XNo
kpInhY7kt2/uITP5mTTCd1TtBuQ6Awy7/LNvZ4+FWLZIwO5vywkjl/W70KXzUw1S
AefcUmaT2uc7LnwZ/tPbDdXbUwjTa31BHBDzXvais/gGUjV/pH6XSrWkKgyc1nFT
Zp993lkySDDtqnUT3DNjvi/WnMP2o6n+j2zfWmmroeYjX75rdtWz0vcEbjBXd4c9
DwxNm/9vBkcoPTCYCxByfXk9KQAt4vmoyiOeJpVzdELQVDH4wBEFJ2t6vxwPq/MJ
jJlYzQN1ko+rbX2GECX4A6ulhVD2/FdA5gjpZTNxlabVtHw09R8JwFb83Sxj0A8G
/ICpohxZ/FyFPogiuuzhs61sssB4GXVLni5f8t/yOgqTOjtcxyI/fNvIJBsJpHzG
z4vS8viKl/MHbgXHNIANroLJIMSDg8oagEL+shLwuVcTaYIc5RKP6uejRCqwpoZl
amefaTRUSEfMQbjBS1v7KhZh9ZUi1/3TSWXC4U/DnKpM5l64S/3dhI0M6Fwt8923
q2Wm7r5YIDHAi88R3uQVENuCP9w37xcb9zCq2eOAgIWDcIJGZcXlfxgwPMfgsIyn
Yh2021zIj6vHnJOngQxGOPxo7hirJO7qzSDowhg91wXupbFvcANcxjiQ9qjHRs5z
QkH9sW9uEMGPyymut9ylkcfN5pLbQhRx8XN2PXBRLoKIbTpDUrXonb9SS0ClXp4C
1hrQWWLEL1VJHl/cSHcfcoeJ27gKLA7BJdivwMNUG5xOqaALz+YXrLKUgPfBh+7E
sNpew3+MKYwQxknekBZ1jFrURppYTihlHtAilVwOlm6CJHXvmF/RCYLkHzM83wq0
ghOS0Is2q/x9zDRz5aR9b/yX04quvNYaylHDZhTaOvjowyrhwQwzZusibb674/3F
08dDxqQpiFqDZORMcS8lOxu9C88KoB1XbQcd602AhSRObqM8jQJHEyybb4sIB+Vy
5N8aAKBSbMMz1nZuEa/1/7hOuRdzb2MG9stPdyZ6nvDXTbIRxLey3pTAHRlJJV5g
+8icTCkB+9ciq0XHu7CPzDRh1NZdFKaEPM51n/ioHwyJHfJd1fUykB3h8sM/lXAa
8DwrGHjJdL49f3+xsi8h2r5MxIa0oz3JLJY+oU3HwqKLWA4RXA6noswRCtSMZ/nU
ZpVdVijPO8Pw/pHbVfEfv62vc20g9xRMnBDbm0VDWhWhdlsFAMc1L4dv/a8YGlbh
WlljDnYRiKlaNTfEm6MUOyIFf6xlZpiTCsLGMLPxwU9gPSRM28rUPF7iF1juDJ93
tjqtvmyt5Vrw91D0ECZkbGcShUQ11YzcGy7CK41yTl4KrnJGrnb7BWFQgS7+Xm3l
rrUJ5qPuh5YHr1IHdVO7Dg0+L1klDMQ3S+JKxHlo5SBgAXIUw6+ydlNjKjPTBbQf
dHg+qV8iW/4BnBTI7VNVmt3XKnfLihSyuytrubAI5jdgk72j5Ahb5iSv5ITOtAON
lEt7cdVVJRcDrPCJtNWz85oq0qZmnBsHNprOvezCWa5gTiyhyZzYgX8zPrk1/lRQ
yMk+OXTU++uZBJssxCzNdlzQSSeOXQXziBkBFeWOX8Yd9yP8Dafu+JcB0tYYJIF0
td+xieLXEuMYETa4z7Qa5j38bJWhOb1eaIocz33Hcuc7CrtNeqctUNpd79ISZpAe
/Q8qs04jKk4gX1SI/jN5Nmlcpk83NgJs54O4v1xycDvAXiTJxqgC6vxaTWuMzHlC
jQLPybcQEJ7VbGkBC2rhjSPuSvVVYKQZJtzBlGTHd5FjPGseXlarH+51/SD1OC8d
nznFgdn+71TzJZs27nqKwP48J6jIdjgD59mdFkFGxdMF6pEt6g0dd/NvDNWEc/HG
ZDDSx6/Gu49/FsLG+lTw0KrzQ53VK74zCMR+9TJdsYrcqw9TQ3GM0RDoim5HCTBM
1+r1N2ipjUkFX8uwNc8NgDRvtEvmgc6x0F+ZgljPKUEgG/D4cU6reZbDvKR9vAyh
EuvDkXbykNkgWZP3fiqKcnOGjyf+KTsyE+IqX2X+Q5v72NtpPufC07lzO77LBl9e
bP5YrUCF/uNSEibM1ADEV6P6lGDLHWuwgIib19uTW/bs/UTJdD+bN6kf5w18LLA9
EzGqIoVh2nal6w/MEz2p3TjtfKOi+3hcQsvGu4WrQg98SeMS+KAuJD0GNRseGS0/
lTTIlJet+NOplweAebSBFlPYBI+yMMH6HOvzlcfcEi3QhQm+F+UxADSEibhz/O4i
iXL7hksrfKhTNvHWnllyjFogigSsGVdhwqMfWZ6PAlBzcbmnFQ8CZcFFauZLS2op
72gj380jX2gE4K6goiyRBy5vy6l8K8mwTpJ4deYtdjglOm/dQlFqwYJ/6ynDgV4F
In2zPr9RdpWyVQNTXH0cOnsARX3kJae4VK2/gF9AJ3YC6jsYo2b6uiijhkJvQVTQ
F+GhxjqZ92i7bC3KaC9xnRC4J+XJ7XVERY5ugcr5hMfOOY6n6AWEIhkyFzvI6ftU
NZCLZhbSHSTm5Sq7NjvPRnur6EbSgs22i5PIn90zhBgOZ/+3tcAMY/rT3OSisah9
LjQh5xpQE2UYwZ2iYOcGvZ+wgdY3gS6z1McOy3gm6IJCvt46URgPe0nkyISj6VKM
eUxuwcDoFjo9U6WOxg/SjxB6Xs8KwyaMGoMJ9OSLAdlR1WanI55ZsgOV+LXcnJio
UNA94az1bs/UOx22nRrdHQvbQOzirhRoBWrF83Q0IDfwvUSyGjrkZMFbfsHbfmTg
SlJLGWdK0oZ6o4TbtrKFzczu2+lt8xNDsdT+N0BUIFmuSUx/AfP/+jqFph436pzL
zRqj5Pf/q0BRQKkqt9le9M+tV5pliDK6pnfjCKMMsxehCW+A5OScVoQrDLSydYZz
42c2L2057m2hR55RjXoXxz2hR39Zvkz59JcD0gyARlIzQ5EMUyQOE2EhNX89a40M
Ct70e1+jFeUO5FcQQ69d6KT7HdBRfmKszh8XRnmW7+xM/k1ZfpJkeOYzIYJXtbJC
rj/cFEMXw86mfp83iVKXEPq3/8bu/WuAt/1Hxn5jCUAKONGSY/D2OKuu3C5eyxs7
H52M1myfNtugZuenkJE8I7Rxyooha4YOZBOzOm5LbE5U204xECRSJP76yX6s3tVe
iE0GU1Lv5p29qTGxZtMNXlKXWJmXMhMqMXE8RnbStUKKy0raLUWAPW2Pll10Rojv
/otiG9xUHtQlY5q2X6TwPff0hwyM2bM1xvj+lGXyz0iIigXZuP1fP4DWbrljg6oH
/TtbSNGFyryRVfrWz4CSbbtCUeVQ/B7wSOnnTLDBXPJhfVLX7SsJvUw1Vf0wT07A
iZOlX390fI4ULMrSz2y/+UKlcBgY9LhQnlMhJL9xsjZgt9qqnWztkx8xATQoQdMh
b/vXE+m8d/ji/LGRcUX7aUzuOi7jbxJOTHdujlXvnYct43sUFKNZC8iTjbz8qmk3
oryRUidyvPywBPhfhtXnSST8qfCZaw8cVPiorcX1A49j/nCUBiZ4iHtfLDamfnPF
uzMvF8W8HIP+9aqsgIgFPla+Cu49gb2S9n4CJrkGMpXD5g3Ahn1hx98UDZat1v0Y
RsLufBiT0mTrYMr2hXTTuxcRUY81+Mpi+5ZMZcYyxT9J/KUd2Q9wyaQAD28n2+oQ
MwSZ0SPv2hD46EGpwY2uAdzq1p+p76zcD2fdOW2WHJdAo1vmSLltuIRR4TF7SBEH
hor6scu3syAGY5uxhW7x7ydhm05jSWTJ7v721f6jgcQ5icgGSCnLGTAN1IYiAxqy
yMxFZ5hRuUeqKwfJ5PpzMgGBXZNBB0OiqR8VyJoTlXVac6PcwSe4LVUVGjyigwJF
nJcUGLmmUmHEQ2lV1dNdcZ6j9+7w9YTZKa4xzF02DgNAkIDMg5hzxoC3KHenFn7u
QcY0mzajOR303m28/A61azf1trOKq0B8XgqLxpc5Tz2MhVm1LLCHCoeAdB9Xckoa
VGreF8gJeQAuqe6drSsEmmkXoAlWH+fUqq0tYBjqDi9g+BDQZcYmCtWQ8MWZhVxN
X/1exHuivSdAVZfgVftQ3jCN9FaBBkV7L7AJaUfVz6syVPmX1YU2ypCmUnEIiOj5
rImbmynU3wHr/ChAC43zbVWoEuj5bFHWeL6twPED5WLb1r/prBEwwfGgP8q2B6r9
WMU9/tpPuatsfLew/5w140tLGlLrDZQJ8wanDzeKhkh95ODX8j7vxdwmnNDflSDq
sH8g9FGfh+nQSgW5f7PfFkAAMvcFkonxCSWJVqEwrbTuWcEAuzgqR+XW6WlItMek
uBD+OVv4GtgQKUxAvDjPqC/acIIBABOUdlP0SHUwL1RLMSI/xUPh+5Oir24xvq8w
F3tm4VEqHQslhrGFHnqRVZxR62mqbqe1gKQxx+22PA0+Pzen5DUgpfeYtrncWlZN
tZQYOSz67RMxdH0lOr7g3EwmpBR1Slv5x1SsuKwntWONC8yH00IPR9+sccXhTZzX
1DT9WgtG47gPpCgy30RFtfj8LH/4Z0jSWNR3SSlA/o+cJbQhzVbCxud/RvUpzTQN
P3xB78/xzH6AQRaFSeEkZcAMhxQ3yH7sEk01xq9nQlCdbibYija/ncFQjB6cZCRB
ah67vYqH42DCueh6gCKttqCM79EfJVAZe3fUB2wpeZh2edwarYQDQ2pH8nCEfbM0
PxfaYXTv8N9Rree653OR1wMWmeTpHPQg2qTnYcKu/5AiN0DiuRwGd3Yz8x6Wd27D
E+Rs2YRs9LUpff7zfGm1mBogjIbQdBWHhfYlXH7ubv8TBWCXlP+7rdC/Dy1Y0x35
eUgLhc6qrc+bxrKfpudim+TmhJxno/Ynki3K3ST0J0uDmBXR4hhH9bNmezzovzba
RlRCuWb4ugMz2lG4gtAYbJkgNGWGx05DhaqpNgQqRcyLc9OPhjBuvpa4Fm6OmAJ9
bD7p6PhIWJyzd4fSDs3RWgEWWmrPTNKZiliXAuyqq5eLugzqWzSk1bJI7ArxSsRe
D1YxvvH2K0VGEX3aKs2NKCraU/OOtPWQ2RSV8uvSPs1MgcEaVZUkTrZkAK7EDjcs
Op8dNVaPXzknwDMpi1+Y02YjzPvEwt2bgcMUiXsvWtz2+2teYwklcAs8Am0rWI5z
KRt9ee5VJkIuHX9P/rsoxY5esvnEb+KquUXCCh2CiUBLoU/6456Zk59rY9ZTe7eJ
XRCQxI9OKry08DMFfcyGrkC+Ep9tJy45KCqhwfdRHJVdGd2+Wf/7BpeTEnYGJ2Md
wK/1eWXsu4YaVRk9E1v9X+D6HCAsbSddD2DZwyYjQdaSNYu2stYb5slWkRgYWlBR
HtpMd0MF1FEKyTvZoLcBC33gC417Hg5mHwPcb0+WkV/+o3Yfj+cV0H4i/zcZ1imU
JmQpRT0KEx2dPOwcRXOwQSWKYHsH1mnJ7q+uux5PEgy8DykNdxOevF3awnQlB46y
w+j4/m80TmcvophviSRsVmJNojRHndO5PRfZRPEdE6Np+BlpzSi31lNxE9jrk5+8
22HcXHvgXsJQRavAhvyG+hnyAJbOkM3lm4YqPYlUViMoRW99dsHxNV4kfGQ0UWq1
KpPd0I1WLZHetJt4k3iJ/FtLk2cohpwhTxlDA3n82es7gaB2xmokMxDZbn3yacv+
aIRErppFVGttX8QkFbb+lekozIkWUazeuxlBxWaH+ltjG1odPGmVhjZ4Ex+mhxiD
40Tfk93fx6YpbgemU1h+zoPhMgTILBNHwFKYz7BXuLNo7Saqxl1jNC5+fcwjvs2f
rmRbWhID7MjxFSk+8O+n0zQ786+JqCchlhL2k0n9I5NqTM+YYcqh15JjANJGXj7V
QELCjUpFkRUJnHD89BkC3XxVkavIj92DiJyVP6sd3RU+Vz831dvKdPA3zlfYxX3s
VLANHwKKHqtpoCTrY+VLlbuLqLe2yXRF755OeicbPw+oIfstQVUzZ5qx5Evlomyp
H0y7RNxM+H58d0yV+h+tAamsmFfeB5jmeKOnSG8qjeI1MMvRb+4It4YDJxXzPduo
6/dQ1YuP5Cx8on9xsBvnZfN9G6TwGcUrLRQO74IESPbW7HelIcQ1X+22GnvtwuQg
YEA9FdoR+TycKLudl51YqZfuIgA68ddWYmUJsJqONJ80Jn1aFVYuql02Hyo/rwAn
0TClZsnrjgNMG3F/1IArdGrVG6LZZ6F08VeFmDohj+7ClxggJfXrFOI20qxCYhhq
imoUhIDxYQDg4xMNBsbTqztBQ94inYPS7S0MzC+561VQzRXDhivfLifdEkTGFjdy
HG4QvTHIZZ7BsvsQdPbHwLx5O5GOED+RQaIUOKu0nb6eIes+ZGxvphywMxYmgGhX
rrb+06hFZbYWRDwAiZPhAf5MUsrHIqeybCiEZnm9o21SjVfM+iSzSHRESjX7rWUV
81zgIDtRSxk5RgMlMvWbFAeT5RiYtYu8RQTH+HXnMgcFWwHly/AkId5mDFhGiBeA
7h1X20BuOnmR2TTxrwjkhSxt8LgH70C/36kyaOsph1WMpxR/EdxKIT+HmUQnErtQ
3GHLLCKmnZskCmXqcou5TnSH6AT6Lo4nU+GaDtsI0aTBYFTyRDmpeEWdNW26LNT7
U+1La8Uz4xt0hVufF6dgLuWIW7lpsZ7BFmrhzPkbs+6KK0li5C/VRB39VE43cxDo
21NKXRt+Nsog7lhMe/H2j3GsUFX1YqAHu1JHXYlJjpRgibenWXcbyVTHiZ/K5k2j
QLrBSxKl7Z5KrWkb+/knydBoI/ePkLxzLiuck4NQg0gn1qHVzmKC7zRYvjLO2R4V
GZ2uXBWrzHGVt+qZkYhv01jbyLeeDivMbW55r3/HhiwclX6CIw43LEIQBlH39pll
WhfEZgSO0I0chl0oeufCSf4mpvtrWhxyJZDKEXYnGgDhcMFaC1wbxDxS9AZZbBYu
UDxK5oCQlluTyqs+h8kWz8oDVsU56egwkU5iJBeisCN5rfUokcG0QN+Qxs5Rc9Sh
JvcOpzdIJnMDzk5enXtHLQbO8zR79EPnjG2+Vy9+Z198uJ8dvHxoowMI/AUHGb8z
1iBmV1zCsMCQQcdMDCHm9rwuO5cPqgjsboaw940Jm8uOuTutvbLukNEy47WpDqLh
E/fTBprEJDr9KjMUIqIkVQplBdVH/gLb50KDO0e/on+XPDY49ySiPKKhwi8P+G5W
xru1VzCKWcAgOb8iiD9WH5swyV266tWX8hVvHm04xIvuIam2hA3vFPl7rYbRAU3l
pH7o2Yoa8J6Qcv6gvuOI2FjxN0S0UJ285TFGYc6TZNjQe5jQI/TOm3PNpMtfJ6Aq
O6Mfw3SWpaS7z9+QuNornxi3dWf6SMi+qQcLQK/1PH2L3KdzO5vZl68/GDUHoAUR
h35aMqw12by8mL8odwheN7IMJDdOIfJ8hS2oB/GaZS2NEjMKzGvnhec7EKQRA65z
mfGi+ZuEr7INwT0Yd6WiuFcWr62g30+0imUGxpJ5TZx9/p3eP02O6pundVY9Bu/H
9tJICqW1nsRF4chLZqyNE5/FagOdeBGdrP7Lnz9dr6yXRTHq0W6fonrkhaFnwE+6
q/EjsWHwC/UQf2t8POkyamwfxYkbTjldqRD9YGE/tvB9jKL/O1MKuyWguWm1k91D
DwI3i7itRp7lV3/PbNECggO7UtN9ylHSQek1g4czUu18GOPnHQKJf0qGcj1OlZtb
wbfs7KjjHrAT4SkNB5Nh7W945TjeqfQcTO+ccfBpqgtAAUYHdWmXl8CBYUgQiY29
NAOzGKJxXGT5V7M4JaTbsFfGMsyANDLuySJQupkkAAYcnJKBStGgcgfOL6k4n4O1
RJ4+ekAIdRoQ2DT85Hryv+6QescUSOFwqnpfoAhufx9h7JkNF9Biohsb8b0j3sJr
7ynSS4zq2Qg8GphlLVM3sF7tvf5MzuhECTUWgZaPCpbFCU/gPvxTInhlv/n8Tkcd
H1preRWdXMkVstZ0g3lzZ9R+/ZxzU3nw/A9fUNA6uvM2BFDkWKvFum/I5zYysTK+
sfoQu65PkQcBPRySVcMhmAcJk63mHcPwBzWTU4NRjHYecF/ThjFot7FQMK79RqT7
2qNSOyWGXEeyjaC22iSZEWpaqb4PzjYakZAdODzcWlHGWFUTqAYjqxY/GDnjjk7J
UD0ZR8NEgevHztJgo7rZL9Zejzf3H3D/sWwXPryVe07Ne5j9qi9+7g/2rx5eMpV6
hkugMMl2w7pWCoq9s+uGAvhrEVO4H5pQen8pUSMZnWnaRfRjTAz4iogAXHiAJ7FJ
D/GtU2s/inAWrN+O6q4wxD24nZa8Vx8zlCkXj4IQXWhHHObxti6mjCZB0fKmWVN5
cZiIX5gfBiiEfQMH5K9tzs56uEXuaPwxddvLihVg06Ext71HDF9h4Cusq20GZVbL
Nas4Mb9S+YNLT5qMMH7SsXWNV9IWH3h+3ArU9YnEFoAVTS1+dceOf4Ie09J5cWPj
NsE+sVeKwVF2nZ8N8IjPuUhZdYXOKHEAh4pwO5t/K8D1ID8Va11rmgRfjLYAAnIH
9/kV5ET5uAhXW+RyJvE94HuqpXDFfzcDALqtGhepOLVMlIGfTyY6mYVqAfCZd/Kn
8A2wTyoEPv0KZnH4Il5D+j3ZM7oCH1uBN81E9b/GNWB7vRC0MCq9APNiWr2GMm7S
JM1yLJm8oF6duyzPoaTQZbBUvE2rl86eDlUCR2QsrqFDEd+JVuLC0vm7vNGxMBOS
fMz7fHCs3bsqIDG+cDDaGK2RM6kWsyshBjzzrYAQzIAPMnE+X0a3KkmEj1sdJrwE
KBeGUSmQQE0SNRVNPb547fsytXyl3nMKjnF5wCJLs9UWx27huxe8v1hDL/nZg47H
+YrUIykrLJICM8RULRphYNKrhd5IjoaZzpHsaEN3pbikVUWT17Br2AglWkqSAZAz
kjeYXMbVXkBcQXc/HIT3Tb7SWSzfM1rOl46VOupLoura4I1k/2c7tCvA2tfTd7Yu
SpWlmfZIBYvLBoRmIttoxUq8YhqhPIKok89D/JgRwSPk8C98a6F+CfZb7U9cTml/
OWKC7zjqAPoZe9rtdjq+8+3cAdvTy8auO/l3W4E6OMPIvuRyssSRfI1NxUAP85hY
5E4Se7+QdIfQhlGt2L6cFnYW8s18u7a2Q/YLaPonXZ2kZec9H0i1AIpRDeKBHspL
X4LII/QNaldZGH7TG37MKS01kE2hiDtsVIMCLuY/nESGcTdyuaFnJinpO/ctIG68
CI6c3bFs5/ZSEZTYgOp7FoSvGQIwJ4JihNRQXcvcoffiVTn17rm0Ou3frHUdD66H
sgbZzWy3Bkv1zodDKsXTNAM7OBEvlKREzzTM09kJZdQ9397qwYbePDHB+jx1oObZ
GE5+wAPPSXVTgq3jbErt5L+HKtnRfmqywSnCqJbMf1sdxajxbWJDIkbsMnH1IBtE
GcjnXWlO3L/kXVDJWd4RGLpOfJEmo9OwAMq5h9Jmo51KeSRWZYDfkQKQ6wmc+LCt
o8FexKeKbzaJpGA/NOZStvV3hSMJCW4Gm0gntqg7QOCz06JcQZEaDewIZRB8Fl0L
G9IDvyIGY7I7tbp2mDjAmcbm3n/aprknYmCwSTgVgAktfWbZBU8Ouevj5M0dQcO2
FozOzC8iLMW6amJ6eY98/7k7EJTYJ9qLdlwQ+iNt8mdf8heg6b4rDt5CLsC4l53v
GjnUq1p6B8uabXStKaOUCYJCL13pU3vUXCMOJvVYmSiS68oWEn4XjzVsSYdGNAdl
et2mKDm8gOjBA7M1VAQgRuEX2a7/RRaXBB4t9l9SsgwqNSFyk58WKpbsFQ585F8u
narfYYF7Zvjcde9f0+1LxBtYvaIodUYQmch546t+FJG1TTSdSqv9SBg+Hd4bU0dm
7W+ign2BE2mF2saSJr17BfAz2Q+fGaaOT4bEtliXVC/vQMiq5mjfRH1hRuqqK+0v
SCpsvaktWFuJ9h6sJanyBBD7u1Wo4ymlETWemcSHnwRxcq5cWbQPY0Iyoieu/WjM
a/7Un+Mw2Pk3CG5U8kk1tDd2Ypo2jRFWQXQkD3sBB7FXDBWk6t4Fv1A2kwfaS5KM
pFXQy7TYLVlZc1JWUYWo82JkjWKa20eGiHwjwDE5wzvNEyt91NBMIgj8rOrbNbqg
DtAnGw31frlGU8mIfc8m8umEFzHlehSUbcRAsdkmKvLsfYph4rv0BT3r0VUZamWp
MUJK15tC78GfqLzrdvU+2tkIjVHqQkEaEaJqBfVkHFaQm/h0u1SAljW0oUXqW/E6
Q8QhfAqn0qR7XSQo/o4Mu31rb0FHmX/OwX4iNuyxpvWZtvSFE23XcCuqrMl6hkDv
202TVF2V6tEZw2U9MNrflORFZvt0qHS/tt/8VgnVDiVo02jJ1FieaISjUuQ9yZx/
jRNq9tyAy81Holg5NDDpLfq1elU/TZ6YxLoXcg5u5PjbEcAWE77XGSJGJqZrWNYY
024GdxmvUtL3rhzD8iA596+petOVrfvJlzHrg5gi9nTGfq3+c5hbDJXByfzTyX1U
9l3ZABDkbQ//oHDtThwWWRaeIPULlli8QcCYTYb/ctotCsf0pt6GXGUTY5YG3Nkx
Zir8ZHry2radyu0qG9FOalPY4D2F+ynjycXBbvaZiuQzeUrm2cEC3yQTGXOXXrN+
JwCprthTCgIH99+0AgwBvN3Vkcv+Oo32u+nrk8gZ4RD0YP8gvcG3FnOeaBTKDg0o
q2p8v+b1IZL2PDoJMn+qIJ8ASDqfjXDNiiTpMjBscwtaaZFjdkY8LCS2Tht4sFZf
c6bW/wdKMThiR1sYPOFF+6g/quiSQYnm9IzZJYys9uG2APFZpyL14HD2g62GLBWr
8LL0Ne7giqsye1jFmGrUeBtuQiyXPO2ABzzFw2/yJtZ5U8yzDvrzc/lDyzhHm3HB
N6nZpuPHpWwT5VM3XiZjmmZRbUMkdxMl4gR0gsAm9x3T0uwYBaG0vECKa9ePs76w
syw7UiFk0Z7t9FMXy4h0VAYdsoBOJso6EVWz7N3nMCNh8U3wCW8yixne6UQhvFyM
tzXCFr6RB5YKgq2o7tfNW2xCefR9YmlY0q1Znb7vE4gmiVgrqSWmt9scgQTrovNE
pcgzkZxzqQB8knI0OpTZUHbzO1Us7hB3DuQwZ4Q+xF7FuUKR48INtblHD+ZyiVDf
LqhYktif/X8xD4J1Sb+6OAuKWcsyPk69pHcGl9Tit214Mr2AZgu7E+VrshAmsapf
pInS1yKIa9RELEVoUjo6Z0yDbIay3YlP90MgsoLvQzdg5bmxLdr7dBUJVFPy6uOY
f865c1/kSwQvJW3sa28VtZ+rFhDGD7fN8le9mdMmdMO/AV8aXGNqXflUcToOPwMD
QtvqgucGJUGXedL4v5EPEDXi0T1Q8Vig7QEPdQqnfCZy9O7FlUqv1lF2L2fa5Dgd
Wv3iQ19KOZhkXRPvkJB7CD5rspYVb9v6V8Yzt4HTXMzpUhHrRvKbwzK6993NSR4l
p976SF8ABidj4Le/P7eEhJIy/W7y/xKsJ5VbEhJD/WtBOAs9k+uVOR6KFV+ObhWb
rrBTgTLe9jRKzyQDOVATJteUFcSN91cynjRSkfO8ATUysQa97Ol/gZgvGb2Pwo4I
J4twkZMhB9AlJfujyNVxzok0qpJ5DU+T39Ob617kfnmhaaeieGf4QNdtCNV0EeQI
rtEI/l3WFjZqePZpf1/tweGDBMao2ceemaCWQ6HF0AMHy86ZpOPtdTLfQlaNXnT8
SVVIfiWVgSMk7QKbaUtVs8NV+/9n8dtKHAgdJj+XrOKKsf3Bb6NKVrKk9CLbbexm
JdZYqEjQsS1dcqx9M9AgsM54NpdeXIyyn4qlRSmt4fUZHGZB/87PQKkStMbHWuqt
InEhfkV04tAjpD1gf4sD5Q4XAdNymd3oT90b4Cx8cdTdOKKjzd3R9OqhDP3JS55v
G8ycRtQ96sOVYmR9c349nsBz83woUePASyq7kP4+nkPgTtPLUKB+Xuc28QiFhuxb
k8iVxoglAuykZx7B5xu52C4uwyNskeAMFZstS+0sH6n0UrgjkFCDZU/176hfloWR
4avlNfN6dyeCN8DeffkMJC+qaKmgra60nO5L7dACGGlCBtNuVO31Ueh3dU3oJLWk
DtOmDuSWvHpa0muQ+QmsKEJeAaTZGASHHJ4x9lqDe9P79scMPkEoCY+eeMHHbal/
vG7qwRiMgaBBpm6QW/jpDjq5DPY5t4ax+SNgfpiklrJpgpAml4ZnfLWSBUhxRf3C
aI4Pri3uydmvzeRN6RupWQjhtccfAhpQfKSeMI9M409BC9/KlDJBmCwqJFfaWZ1A
oSLPyj15ZD3Xq7oaogpez1PZkDLx4FQJdcdnnF5gOH3YHoQEcwKcy8FXuXtihrmC
l3ok82HVR+FURxcCCYHoJpWUaxa1D27gCMAZAZKEUQu3xgnvF8q7e5nObYGNm1Xz
uOdLSvy6tkw/dtv5lP17cvAH+eB7VYd58GmgM1PuTAXbFuWk91anu+7Am+guQuWN
aMVPVonfx6VklpSwXBNlfcEpkBs1j6FoYoegPGS38EsDmN3yzZ7AnPS7f50qiDg3
SPzNfSkjbE5aoheunUl9ezVjmwOPoPSLusb0BYCTFf6yjztGRIf+idK68LwRbBh9
3uXAraGsZBncHl7oiXe0DyqKoinRkSdGvWp5VO320pnHB2e1nGo9cch+3fe1YbVf
a7/KandmK9s/J3F/w9JjnLh/ovNqsKDXLVxatZC5avV0F1eenleWxLq8EKqummk+
uZm8fcHa1f8XWmC5hMsjYhDgQsndDRc0WxxQpPm4GAsmZzwN/BhkS1SEYB+4mVHX
5sUQgSGoHydGsd50TXNlo0ITPe/cNLCmyfMcxENEZ67VPPa1a6JOkbm6TsWYDs6M
jCxnWF78ROxJ9bMdZKMssIpfdEJMQpGJh8iVo9D6GEsSySA7AtYg5TQS+Z4sS/F1
OIJyPe58J4MJ/FYWuk+5spQu9Xn6IyDx2f6ma2PaES1492saITBpLZKcOVHN/uAd
ew1rq6IulROTg6+sF09kKtouRi/L8g2R0O3WCdiaFuzu6euCcO0xldO6papPkGMZ
Tg+EbrKlfwipoRscNHZkQlVMG650T1KhrQSPODt45SY7zAzOUv+hOLrwwPtYsJ/u
hv8xYRrhfqxzITlQZfMW3MZZwAj1g5/h9qnJlQ+66vgu1M0xO3i8D8FQ6rm5vNPr
MjZeK8HTliCwjpb2l2LN9djVfWzeHxwn21YDMGcflBMunGG5o8ud6a6RjKyAmaRS
FnzlZkvgPqFAsadCzSQVh2Rn6MCCxeiGwTUQATwPYAQ8pX6AwI/bX+VkEB9CxGLL
NhiyoEM83za2R2py/7YzgxJvgSd8yTcunnV0GHloqnbz/CLwtziO9SXY+V77al3c
X7j1R35YXyqYedv4ubvmLGy0P1c+PKyaFo8kYsgb4kfKCCLbagNus261FnUub/6w
uOV8ln4EZ2dziIAF9mXd3k8USdmrxGAX2xeMG4A2UBi0lzlA/FqCn7id+tCqslap
gHNuR2gM5lEFzV2+JWUwlAGxY931MUwA5Y77EZbEHXjlEPYEEq0XSTWKp5NVb0bx
/D8mxwc9SBT91nVeGkD/MuaxMPwzXWhNa1LLj5M9YqtGgwtJEHvDPaH08a0G8muR
8yyiX/ojahm1IuPMxqKsaKjiy8nydVT4k9ECkSNh3IzLKhbx+fazHj1zvclmRDY0
piFmNgenhHbTnq/snvSEmdVFwxXgbO45/JmslcIUhSJaM6N+/8ArEviuEX5hCmYj
ZRZ847ZRDeUN+xun87VKlavSa+f20J2lAn6J4fb5TnLRFcomZJoe5GcUo9cZWkIq
SyMI6s3Yw6TZhArJPNd9UIByYGy3LOEAn64WR4Z4q5dY/AnhGOjzO3XSGlxISlGt
NGNzr3S6MlolZvfN1tP0P8bIJ8V24Ue0fO0EsQy8/Qr34nS782+4QS0ANyEkd3Hg
O+D08js2ggJuuiK8dN/p0nIFQssBi7r7Se8kU1AHmghIx+DkgkmAbGtlhFLaqvfS
w92C47IifJxwkiXoXNJL3qDYCHBewNfufTnXGhP799hIklHXCXVRCdtAzNBYW0w3
nnbQbiJvg57EYrg5eAlJRNZ9Mlhqn4LGjDPksd2tU9wMt/6E24LTvmHPONXTg5N2
mIJ6ZEsVm1u4608kSSd29NXUmQchvddGlLWuSwns7vAgsffqI0/B2l0YbPDwIOWL
hxpcO29MZP0lnzmKcgnu1p7a55v164yytWXamrxbhLjcNrMOanDAskwq1bzSRFVD
Ga+8ausA72CT0k/9aAhRnoKf4LJINIqcOzSNOllzNT+i3IH0Kj730DEyB+E5ta1m
tAeg4usqjDUNpSumBFlJ4drBikmywhIDTSN3Jt4pgYj9b52NZLj4+fyKMDuMBCRT
b36aQoHyV826cV4vavCWjRvNSshp3Rf4YG4K59ws2csjjCevhtEEne1HplqEzJ7+
hrQCqZDxIX24CPGSrUoNq5e9gPRWRbto6VVvfpyXbbroSNR4TVvshBwbC5xVYb9f
XJQ2oS9ptm9SOWPLBV3NSGrh0RTc2BvS6vJZdt3J1ZRBpYbmWRh0z99/6zCR/XzZ
GK7XSp+dnHOBPIgTnpsKaPqwwZ3dWjuY0XecvoWo84azTyuzuom6/p6v1JZVGph/
Vw/MhdxKpsSgYmHfgC3lDS4WO8fukfj7E8z+CQxeIEEdhx2gRXlY2PWL4mSlnK5r
P4VkFLvNuTYoyxUwMnpTt+0RUHvVw01pBGzeyEZVeSeBKZFIIRG7Mn74CpyBOZIg
7fpQpXeePhHkZsemIoXI8B25i0SH1xDhKDOYVmEDWIMdOLsj/3RwLJI31InmmX8P
JD1jijlucJxYi+RkbJWEnl5N6qcDHx2r/qmQLsWY2yw2rAw/CkupajCneUVWAXQk
P0WhC+OEmObqJ5yEEfxpw2Z/76OyIYDolp0+YLC56FuqQgo9jfEPodePNNhNsLIP
IUkSIltmD55ZvwHKeR1o18psNApDzxjBK9em3zPGWISQdfH1V21sJsx4SPi/mT/+
45Bk+DmA/BB7d5QOSdTq4vf8DnIwZH2JIALBBulG9/Fg98bIgeHOMd9S6IS+gMs1
c5Qhj/2tifl3HTTMSx08FKZBO96ohGPKZleah1emu43AU+f5A50yKLy7L1IWgXtC
et4mjDxIC2EA/IMVYDPjlZJPnpiQd3BXc3yUem5PsXfLBoc4WnPYM+/2RjBWKmBK
7sX1x/Bc2+tRs1kcUi/H25BAzHoLdtSi7oOgqNvPnts31S7OwKjzJODIkJIF0esh
qmPJL/EubrXpTJebAupA1lYqyjVcLKuefaxqoAx85BoO4YcpsEGhM+S7GWPDr2qr
9drcWnq/sjfv5pBwqYh1psALwgn1Pzz7Olicyj2rHrFhHiqE1IUg+Wz0MyDZ6Ef/
fVnvBdugwDD4ucOVfl22xbAVZx9qC1FuW7fmWUGoCYZuW9zxCrDLwtE84UYvcdoO
vuizJMAuDVFL4OgmNh1deyzNXNXyXOpqUGactGzZOJywFbtFUJHRohtAWpVfvmuH
OuYabFYy0u2W9zAbVKsmsjS7e1oH9X65B0eB0F1lKPpmt7LIlSSHhwiZCutEUVWt
+xcdOSqaF2qZqpfzfQ3WbuqhQBzigV9pr8+hpCxzzPGbJIFiUrCrLqgdpdrk9kZ0
egWpio67vvNeXvUalol7N7ggPogk8fgRUNX2M9Xl1n1U5cb0x4tSweSA3umFmwxh
esmEjF3n1mLY2DJtCN157X50UyXpGvzc4z+XlYEDHs3wC3wg17Vic6aUPjgm4rvp
EecotNaRt/SG1dyqY76+xzy6oh/SEQbZUzA2/LQcFnRsjnO60CJOkzH/CiqYJT/Z
SHTB0Z7MYUX0gwSZFuRUhb6CkSBrMa8c8oh5SfZZqZAEd54K6RWb/SttZvYerCc8
wONrJTynol3kfiyvLnE+qLqwlN+jRBGctVGQhvT6BdBvAUG5x3jBP9pSv+9Jf1nH
Ws1jYtdP3lIKukMCg1RvZqtvG4nFHwpFHGhXx7wheFunpstZ4potbc5TZhP0GgB+
pTpfmb3an3HqXbu2m5nwLh4ccOT3lPtlplj9fIyGfPUPlYfgf+dqBAlDYqQxKAaz
wjIjk/xlsKOyv4R8jIotAyh63bN87h0C9bgz6E60M9sQWx6NbwaJTAWYcb2X4dR7
a1feKrD6mFLFK+vN7L0opCmHaB3wmnecDkClnS0Fd6vjF5fuujlraFjZNvu+ckyV
JkvwDS01FogTBeLIxYOwEw9DL2Fl57LuZc01/M4HcuErlY57kZ97az7AquFYKhWm
JhuU37KCIziD47qSe/ctd+btaSXQbA5WQwwIudzWgtV4ARnPU/JUZg/MQj3mdrSJ
/I+ebmP/VBGz4i5VCqXn9uONxvxMeRWqkU4N+/H1lmteN48tnjvrT5v9tXK5i0pT
xltVWOsQ8WyobsQIprbmsz3nqWCJ64ryZoCLS/gkHkYI9a3fpPIS3g/O6umifeh/
KDhuKgwDhGYtSbiMxBtMO5yJmGpuSzN/Oa/iM0UhFE3b2q1HiMtNUeq3X0LmI9Hc
uC9Drfrhuwz5YmI/6k7qAVJtzLqNzMVIXKA+E0x5qifBK8G99n6CNIPdI3KIsgpB
m4A7EqEkpa1QGIjbeVnHifmW+rLI6Kp5YbhtrpLh3cA2HL8/PzOZlw9isisgr1XJ
ZON0R/pK6yM3gBjWBThdLtg3X2fBsAV1ru1gmwbUnRA+Fg8uwpRo7J2/On7nntrD
0nBvxz+gVEdrKNFk7AN3gMeHMOX0EdSg3MHsrk03mJqB4WY/F1SIFlUamkK3d6Wh
aUkD+ncDZ7fh63tZhPBQQTs0Ui7+9pJliH4WxUGxiRjrd5Cgym1y3FMufeZ5CXRQ
NmauBGhuiuty0iRHeGY+OqPZUJaod2H/4L3ccLhLBopT24O5OYHO1BaVNx8noMCe
C3N9Stzthux/SEncJxrLih0fZEzXy4vu43RQ+dx11OL7w+YM9uOZUG8cvSHw1/K1
BiAPdJJfWG/fUmsXL1WC0dAFxRzWxMmI7Skws5hblElikJQUuL2N7EfY7gG153Q0
KE/tnofSQxSZAsZroi0PLdza6u++q/6aruvyexkrsfIeQB+ZOr82K0Q57CFCQ9Y8
MKJGzwQ64BCGu+npawdetaSADxOiTT83TN/hGVJZnPUL7q6mQLHjkTjRe+2QThAq
EitpEawzpgfvDP7ftAFcQr/wyGFEfgu6KPzpQmRb8OnSb9uzLFVWMUR8ZtqilfT7
KZ7MNP9eBZ3Npnc+g7/tYg2U9Z2eQFfSHIoBdc+b2ChRQi/+x1rWp7ag/Mk4n3kC
AEzbcqmn9nQSS857iRQUMjrrX7gS5tW8e2zxYRgrJ8zF+BZ5JUVO5QhETTDL81X6
ilCO9YJfWH/mxyL/a9VBvKgP91tfFFsD9MaJeIw2OhSdb1XQB/QvmrKgpZ+AV9cc
pGKd+xrVS2iA/9X1X9k1kqdTUmTATQ6X7njXrDh92Sbwii9jhOv/KN/yFX8a5fOE
uJfxMYPT5FqWZL8v8TQ652uf9EVykhw+/eUyQyR5mCUv6SNEOpPvk3A7Qf3MKe3Z
exHsXEZqLGfDh8CPFf4FHdJzjX2gLlXArl7jzXejTCxpd3OyT6+agKqOsdhA7u9x
AtPRCcS4/IBQSU9Xo4m0Khfw40nZZPqvqK3NIFkN0TAGzDuwDJeOK8LrLDI97Le8
qgW6Mn/H22PZgL6B+EIIzXiOhfWecZNzTNkuh3psd/1Am1aglUUynzM3P06NxIIp
XDXpBzSiDxZlSvT8u6JG87+FWEj36kqjul/82ZIh/0WMyjFUgKpUg0g6CazDMyaL
0IqY2R9JV3R0zoibXZuIRwQpnPHKWzQlfGEMVKze3mJsXH4RJPRtFu8RpFzyHMHr
ReESLrRYiX82k91vqW65372UlX+17sqWSD22mj3DjHfsLXZX9d4/ZLYkh/qYmR4R
uaTLfyYJbseUylIzGGY2IllzLQcQH8nkkpRCx8jAL0C9RMzCenG/rZVOmNSga+P4
QAO7bAUkoWyUBl3y0jKQ1gPgqArfYEvDuymekJrJL+QuW9oBVfFiHYD7ixIvE6l+
F9cSb6/9VA4U1NwOItqCh8QXphUqw/g99tdAfMeZB0K0oaLXAfauc8r3eLgE23rQ
8arjl79C0yoSAjPtlIFENrfATJgSUqa/K390z5SccIC4N+gYD8x6QrEOVP5JEKDg
ZYkorRvj1VP6lLYKIj9/AY3BF9gZQwORLxthjpEMZdG/Fypg2PN0Cx9g94PIzTeT
IwXdY0UZ07fksmQ84uX5P7jerixZreL8h6G82byJlTHKBUDgLNJHbegajJ21KLoD
vjQLys7xMwj9TEG9Xz9yvGrOlwr9fAt85KeY9NtU1r8lYRzm5tNxPK8VT7VfqLAy
nZsJIgbuWwXwyzUkdkxsvI2Ae/LsxkiLU2vly8uw9w+Z6HWTxkVJyO6Kh2g7gsWq
P2MAoP7TzBqM/IXP+v4YLnc/wEN4pLYLQPBUA9FBILK2mjJ+/dzdn6OV7EYmJUFe
THeFYCIhY/6ZIILe/Wi7Ia5Ti8hneoeuWDDRbGJPWyufcORs2v+AXWn94Xf8VS+a
I7JA82SiJLg0cCl4C57buSWOC39e3zwd6AbusFi7S8AQB+1Tq5SKqbub1Qg+jtl2
i2A6iCknPb35ReL6L5Er1Fi/TmFRNbamSfC9vlqRBLMaKRRAjgMk3j07sNQxT2dY
8kgHD1sbTwEFTlMEKGwC0y9uPnyt0cw55KPs2EVhTEl9vHsyWp+H/lVd7Z80NAhh
Ll9Dll0tm4cQYNhrWflNNBkoweFexYHwumIFZ0jf/Sw2tt8s63V3WyyebzDfBCj2
KExRNnkuVYYZQ26naEVPBtjUXry2L2HErVGOWK2t4ZzEZC5GXGhcdHgUMpMV1q4s
GXHjGpVVRj4upBX9v9Tqk+xXoWY2o9w56951cQS1WFjNF2U8YuxxM5xOtRQg398K
eWqsVJocoY0lHbBKjigW6SjbxMCPVXML9MosfiCA/wRZh34Xj43nvS3j9U3qrOVe
ssuQI/uRt4GzFq0MT4PYlBwVdY/CBPRJq1TFTGO/JvovEr61FSGEwId+3xAa+d6Z
WDqx0zYBwEGWR/qzHWzIhb/daJ2uVd5n9ROwnlNUS2K4TpWwGkr5dKWrtSTGAa7p
ClSKiY5wkkfB7DNTtP8n6WOFXIz5PSOkmSjAY21ZYP5qUwVfue3Kz23PGpILSOyZ
rXE27R39CTIZXOcBFoBqKUFPpPVEOBRPQJNnxNxhizQwDRx+7meIgmFHG9/qmhuA
PkTAXqvOZ4/r45MIdzTGinANIHkkNyDeg0uZNs8Ii1LV03clL/Gvy/tuxweyUGRQ
vRu8hpbyjHtPiFIlo00R9mu3aDq4Un5D8KhjZUp3liuDZOygElV1AsQU1lZadxZs
12rg7gUdrNY5lT8VJuXuHSSa0ywfat50i8S90uO6quCgoJgESMfZT4cx8yWLz1mR
7rKa+UKip47ChJMIDons4f4ovB022nZVYA51l6CbM9zgrjW4UVIxDhe+DkW/eLNX
Lgp3c2Fh4Pycptblhdr0CkcLs4sPzOZeb+Ccucz7kngRux3PTbVZjazKQsa9n0Lv
sPyikppE9YVCcBS53zNnVrnQOpN1wJtDtD0MPp1VYwR1UTJJW9WliGqjqbeZ+NK8
K20Uwk5U02WhlVBaY4aAKVsvQpbXA+6oYKTGty/cCc02nQc7k/Zn6iMOFB4ITVj+
+Ofux/Or3Zsa0ZjLgcAnkg7FJChZMRlEvek6KN3k4rGQQeHsJlGP9A5RT/MET4X8
G+PEnbZYiex10K4ZL1VsOUi1J9icT9SHgGVzs3/CHpsAkBe3R3Tx8hGtfWeT7Dxb
0Kbtad2E8ginZkHT/rg/nD/kvZuVlegxY+mhjWC1hLX7Sr7pcVXvEbSBX+gu4ePz
t+APtoAAiJnLNlsrJxiLdQ60myb9MS8CJXcYQF1eCdUxwBiWc4SoQ87vvszTM8a1
wtYfs6UeUnfjl4N5QdvkW3zxwJsXGFqTaGM0wuFz9XIB+fDkqCRC+OavQ20doUOy
lyl+vuxNRr0QRQHljn77iv8Wq07DanOuTAr4X/io+F9009VYNWH30in+JnT5eWQo
pcK9UqdbSIrqPXLuLdbzNMc/PzW0JJ4lL9t/V29ysMDKfGU/aAsCKaEsl0eT89a1
eQKw44a3ayqN/vbq5ohZJTahmTPPOs3M7W6xd2EG2XZTaYblj47JpmINL67l2Vhe
BI30v/cGVGd1v0H+4eY7dnbAL2c8MT0RY2erfXF0FrjfVoFDsFDJgniB1S8NJdrs
E4BvtGYg9zd9YGb8o3maRk0s0WsT/FEAM+qf1pLyYr6sQJCNxN5LDG2BbVjg7LNs
9ieGyeSD9cld/QDe1jFMdvE8YuGdH2pVTzUxifdiTTubZUTCM3TUF1+ZcNSBldDy
GhZjOZt7Q7JhGynZr45YsnHgg5NaX8XWKKWlWc9m2APVQCz2n7DBYeilsl497WdF
9j7gSUb1o5iGmHhdIE8gJVn3w0YZbOR+4oQujPgKZnzcpYguxoBJF+klYk2foVFh
WHHV/j8KzGTBeV8aFfnInsdOmfw7IaCZ6DbVw3TCvaa9v8Xvwyi8wHdWmVGns82x
IjI1aSOk/iNOaqaKD1QNphCfTg3uCd83wPbLuOruXtWZxU9IkMuHZE51pkKLo01H
enUX2K8qg7H/TfzvoD+YS47hdy7upGfdmCDlQm7syy0lworLSMPBmZAucMOQdWtI
LwbS/HDRswLzgl5TXRybaDy9l8pfDJfz3AfvCqhrtzlt7AOy0gNm3smqhrqvA3LW
SXwYK/KvVwUb4KsKnYvAMY6NHjMWf+aH0Byxws8XXJY7TKinCapuDyPhPa7KgkRF
noOhpkEpe6IdDggyer7sxPRmTmscDbAWySuZArVjjvC19TTGCX4Ne78e9vwgGxx7
oe3II0AC9P9ABW0jSa7HmG1NNWQIk7xa4VJrcUqjuBhNH1IergggNeQykdu6TXcD
+HyW9G3UELNtungK6opdWW1+Ck1DTUdC+7QmMrXxG+ZiybQvcYXxNNqf4c9zMCxB
L0XpMUK3iC6DMFl7nrT/rQZDGvfA0RAsOKeowSTp419PHywpoA7Z4VpZxO2eHp4R
1EqpL3kFyngsig3DJCOK5w1IN4RTMkRg9VWL6Tl2rSxOIi1kp6/Vxfcr6y+OZehR
UoAmy9O511QeavrhSMb6/t+AjlcJ229SM4MCZnZCtLWozQeHUlnVw1Rlv2StnETA
iyOcTTmvHa8AjfhVN/DncJ1GlcRLjJtmcgsGbDViMxPyI9w1tfI4Jj9ElcGeWW/z
wuy/uLc0xXgOXdVUngBg3a7UikzFwbD1IH05uzT57a3/4RF46uzHVaf7Wx3iRhoX
oRm/G8XiviOKUypaWuZLzXDhoVYA+WciWOSt2V/5fd/cy2hT8nyle0lDUGP2ZG10
WhHneIp+AgyR8SLH5NnrEQ0y6esbQ8cRsSG+CWx6uPzCRuRfaUCCMMoeD/qzeBJH
anmCHvEsG4AdUChvkMf4DMei+PRVej/dqpRVwoGvk2PFDiFFq7N05f2Xcak3/I5S
fvvKXeRtS8yTP6WuDydOWWuUF9U7L7wF4xijAwLBuxWa/jyoO0gh3y9aJ2xjHo7i
u4GQJ3/V+N9zhtX2vF+dTCf42bN4Uv+uG4jp49eWE7XBSF5zmN6vPLn33RGzAIaj
YDyhw5qCb8JyPzeYGpXFDBnvDnD1SiMpfGOTw6NQblscnWJZzFvc50l4diQCQIeF
yPK+j6CCNb1dPEQIsn10IoqGT9YoQLfmEfDAWP0GNRc0OFTPkCakcWF+JEtB11qU
yZoA5FNhxBCmIlWIBnLWl2VgNv94hug9UEprh5cSqVp7/3KbLvE4Mj0P0ttQW56r
FQmpq3QqPRxzSbQcYGAbukHvwMpwHhj97FItoIGTsKPLxRH3emw0BbvVGnr/7l6k
YmojfSBPOJ5N++x1fQDAq9vhcxFhwooMxRXt/up1S4Y5C/4u38yQiAzhcd1nzLQy
Qxo2gGGykK0Tb4L1m5cnxctJHfPSGjo0pdqwxJTESOe8YqTAFWLm521TXcq3L58v
TdPsOlCvh0m3+anIgpLWIKLXP4IRC+wI1vWrQtPKt1ZElvIRBH7os+TVpelXOAqK
KXbsNvkn1ZOrR/+lEPRdzH43rgfHop38dmNE8g7UaXEtWUyh/O/4b+PDgmgS+A3m
jA7fjKK2xrZN6/xJXtAS3a8R11rfwhblZHtazZIjA+54RBOOEDql9T0e/4A1Jnt5
S0qGwbeTOwiRtuNjLeMSwIsd4zbv3Za1SkFGW9oW1vo8Bb05sFIXgQtNvYBh6KkB
kenenHCKBsj3MKzIhszpgEJ9mE/dLS7nGeJdRWBBRWC1zKZO6wq/nOnqmVsXjnTy
BMePXlnlrmaC3ZwvYsJi3T2fghFthcED6VNm+1qU2qztra53mIqY1XzfMssdDks7
tMsd43sd69hcfnQwzywdhQOow0gj1r42C1R6yqIT/SHxRStJTrO4Rn/enjrNgAkL
lioyQg78NjCnGVMH2jMxHQuhcdHoVxgTfJ104b5vwARB7P3y/m2ZhC3jbpK8jtUn
ax/7ZeMMDmC8+LrNRv7OptY66K6d2DM1Agvf/W2bI14Xe6bpz4cRE2RERTRdaovL
wEoctTBdCX/YiITJb7Aj6JKFZpa/4CTtWfF0KkHHbblf+wv+IOz6g1X9/OBq0Qd1
J/m2XX/DidbOY03IIAiAriOvmbAXbvZBKCs8J82czd8GoYhATmip6hbRhISDnpcU
QKP3K7sN9AEh5DOSzXa6pag3xtdH3jrFol3jXK/aaCH3HzpjiyV6XO/O+CLT69GU
lbUmpeQaZDsoaNzkvU3GNv/HAID4uP3OXPD0g0wFDNPGlhBNQxGX4pptJUO6j05S
Tf8Bwi8vNzHLOu4OvDl1e+fPTOsiwUrqLL9X0CH7Uh53HlggqsGLr3cH33eU1VEw
8Qn9Fl8kkIR5zAcpxOf5NPtXmzoM5GNQOXSZQLhCUz6PWdAi6B1J9g8eZkL3KfP6
X04mesACs6224bYk/UhLdtcpV1K1b9VywD0jSGzGSikQFvb1VFj/EPu9tqTYZgRS
mGU95QCljsAMeP/mx/Wg6FW/8t3sT/u48Wtb+RJ4jBibGqATAKTk8uZ6i0RGVpvS
sVd0kz3aEvCUrMEI9bKvlMwLxUTL/bRv+WLkMocmxOvcdHoWGzHEGRWu7JRGLETH
aNvyBL1Stmncm9kexl4jU5/v9oUpf6dU0LoRFJVrTNV1dPla1JLmO3qrwzAGK76A
3JO/4xeUmphjGDrrjHXmFsV7BFR/l45N+IlwJi1tFpcoYhgmNdpttbfu3fMFKe7C
tZj08KhPkz9rAe8flk7nLQozNtsRwBkuIr72xU7GAdfxmTYBOmf27iPnpT3xfm9E
NA02oDhU23I3jcGUHlBFn08KUipYe7AbMF+juZLeCfXECP66t6F5I5L8OE1RZWSv
Pf9XM8OCBJ3tTmH3t6i6jy8eq2oERhH5xmv/q0jj1BUhvWeAkiwKzEbMVa12eje2
B7zdDvcztYE/0d6/FkoIt0yJ0IzlJQ2MaiAjlFhpWq2Z5ENGpAyCanBlGVtwwa0d
uLdOzY7LBuyDIHa5aARQxPm0NDU0/DacxxMmb+7VEweXsscNeNfTQFYHcG6mVxkn
2gvt6pe2Iux54fEiSxuTjJv/kjrmAS+wyxQZ9CdpRyng0Az7eiFhWXW4pCmO95Op
3JAFsqqrbxcN1+IWGWA9eu4jGwofJkU0iLi0Qju4RXgUcM7iqCIN5OtzRvRhZAr3
MFEcxXJtZvbLnUcgSCwpP6wLIi+bTT0HHbc17Gn6/pUyuGiqUJPAOW3KUEE4Y0Zw
SsL46xvSrVvvKwFo2kJZ7z4V+LhTrOQaMnlDZDgqQlhNIxixmN34jixsj/m6LJKD
z9XsFMrC5HlxmV8Thpe0HrMhwiO2gY0HsW/IUqgYMmHxSQehbvggsvPH7Rzasl96
8TVu4zbMtts9xceJwM5v/0T1MtjCFCnpw3Ut2TZWpqakeXw9VcSZJrh0ivD07yXc
ngYyGu5/FhNy0LWPnzdoQRqTRCPkPQIvWwuhsQe1eqkKG1LCUSAzv86XJ4v6y2aX
vVqLe0pEWi170eCqF1TSuZ1JCq/MWIc4Bk9AwUFX2ZI1P744PrfxOsI4as9L8STj
/RetAVn8CiOFNVoJis2jJ0CXOMzZckcFhU78rmBJFBVoQF7aPcpRWcctHJkLn4Zs
12p/mToErXymtcxbStn+ryTpD4LG3gPuE36gokX6GZ+bwHqqskhHmmcfgmOVpiJy
ntnzz4LuNZRVQ/qNcUuUtjX9N9vXIwkzbI4iyCARYra6xWbzhy7xdJwjnwX8QBUZ
AWGyUpxm+J+HdJacGdOhRZ3kC4wCetbCJosEFvjRnpNpYwDdF/k7BxZpqVkZe9Ep
UXwIb9GnY7elUFOJfkNC640xU+KjANP2ti9SQ5wKVcflCDilSnJJy2kOD+bDlq7E
GD0PfEaJxlr//oDEAvmwOAp/HSrx4jjBJkqGT41/pxo0Y9wfptUrAb7DVqts68qi
Mm0weiLqRfB7guG3qiwb28aI+uDYDl/E4E+XLI2eVHM/edDxwUL39JgmpE7YZnHX
XhhhBYGtKDLwe76KOc/Y5sSMmhEqXAYgOvNtsTDHkoJKgo6frDosAHpXKBs9LE68
qxQI94CDaAc+wP6tfORb6IhFqAqqFkgH1E8uQmvkrog6y9fKgm6jKVklh/lLGyyl
OFGnUJvvlfUzKClR6im0ogWCh/jiwYcBoLby+G0OY/yU76wC590AqHHqHYvVazRk
WsYsE5cQ3abPhVZw+sIEn9Kl+B5YjZpPtm1K31MnUW8x3VHDEdOI4rmDPgdU1fdB
5B1CCFUoVCUw7rjq4bECuaoJlhNqdro4iDPKg/l+bYU9/i21GOiDGJxd/9Ir6elc
/WUizqRNNMn61TW5N4eG3BOS8LSpMyTnJY4ocrUT+2VksKV7TizoIIhomF1iadkm
WqghulfeyvLnCbtd6jtEQ33Rv6p17SyOZJbvHOD+BZVVh09D6/dVAMGZHgBarBl5
bjS7IJrySI2ic88vNfP/OQe0XhbtwfJmoQHuMEJloDU+GrG9XlY+TFlEvPuRGQXo
rUrWTKZnLTiXGoRXcDoSQrp0vfOKjSgcCgc+tWLi2YTscn1ls0nDdNTazcX+Y1io
hz3IxUDn1WEIReQlfYCWVT1p6/TGJ9jDLzvdDsyuiZPVCnqR9fqyravh29tpbhY4
lbO7emnaDh2DhsH7ldgCR2gcWzAFN5jjTGynbe6LrxKtotclQI8irjUKewswpwXc
/fR6FkmbNh8hDFnSpOPKizO5oBFb7zFBjNFx/XRARuM33pZcn44LXIVzTb2yBDXz
EBS88ztu+p9RbqG9JJLLwjpWB48vz9Sb1n4Tp9947pMaN1eL6mzmcW9C6kuiZngh
gnGn9YEIl2+LR1ZS9s0Iw2jd9Ufkd+35bc6fRn3xfht/llyYU34vR5n6HYo+45nV
P0wlSK0tjg3mSWM2I6y4sk1Kf9UKQ72PnSLBM8z/F0BXfoxyoXYEJR0X+VI93bnD
YyW4z/uE0BX1HIADU5w1UOlEBCqA6I4bCJs/zoOINbkykWS1Abxr9u2cP1T1pUGb
WDuuf+8EDXcz0+1CkxUhH2l+Io9/xSl14NIz/R4vDhvzS64RWrtNpuUhVhFhtTB+
FP46hQmw4ukqu5OVg2XBmypVZUjwT4PjGMHZSpJxXvEF1FNZ9MqlPvr66t8GEI+P
Kv++6c4saYPQZXYx+WIIxAkclXmi8iUiTpF/9QnHqhIGXdXS3nCj2JdUWr3PEwPq
Ugs+6p3hajBy/kOANxW0NwfuscxPZEY+kNpHeEA+5QpNRpY4HDw4qrcfEKDT7e7B
GutiYhj++e/WylGGk6OvMGYGnpo7Oc3wHEx1osczCruGvqJQ583mm6K6zc3dUX4X
2rwk9nT4AGEVlBCivKfwEuVB4nQb9gx6i9qHP4WK08S2gKCkDrbbeDBX2/cr8BQp
EghHNU+qV76B7VyRJpRJVFh/smH7nNNJ0Ocd4vZd8BpU+ZzGaZwPCkc52cOjStQ5
0y3766Oq5Fy+mTxztHddM21uJqRwJn2M3xyyVTcClumLv43x4cIrhjK636jyv0iY
6+Q38QchCxyvB+4cqIbqjxr5Z5G6uXseg++Eq0ZKCOjkceKXbRj6YUjQ0TYM8oZ/
NHgHxSI2lvRwllwBBshXsXXni1NqRow5o9XXf5YHX75fv/tzC1Wa77jkalZgwduY
G61lByE3fFPPyivdZyyRgN/Ui8kYpPiTt7xbC3cyKqYoKBEfWCuecVWV0BhEKMIO
UFYxXYMV5lriWM5K9DQ4BdCbTPXx3eLShhV9Egxvwu0xPbfXHNHn/Uf4ZnrK+GW+
/5ozpH/DSqS9TDKIJGn8NtRvU082x538rmGqA9OoxnYE8hNmeRYsYefd/lseCae1
6/6O612WtIYHgjiyHl7IdgNak6xgIgCVnwOuDk5RM73CXn+aT1GeEWkoX5zYfJZ2
kaCPoympteOxk4wpEUAjJkb+189mYTIkPS6bpQJUBuVOMI3Fb1pPGkRWXjtLymly
E3Zzd8xZUIMKSAi9/XVO8HWoth5JZa7OGrpQTaIvvYyQA1cpkQ0gnrytOo3WGtck
UBhcbvPhoBgWzxNWhnhAGkPnetXzaonjv4slpSqETjHddVSv6eN4G+YjvtXGulwE
RGcIU6A8kLHw0zgP9nkRPKVT21ZtA/izNC0q0iJ0qj5yCVGrQT6Zs+frmT9yVXxI
b8DJjMyHDi8u27LTpftr7SNyoifzfX2j9STUfyOawCgJBTTs8OtDg7U+nhW2xzeU
fpK4HHMhRwJCSKcCEAn5hXrrL8mTV8O6MDfypvPk+htgBaSXAAMKbYs+F7CQNPWc
X4d7sSr9Bx/wBX1ps4n2aQq9J1FDWfFoWn6DDcymc/GuAIrXpj3Jzz+YW5lizbx/
PWivS4qeB7cmKWOEMeV//4A1/hnx25QFBykDoUH47BRamV0hsomnayV4w7L1UpzT
qkpaMVvtmUdgDyBkyR9tQBO1sce5ss/pOLaECXIP+bhk9VKo2N26+xf+xXgTkub+
E7R0t10MUESaJzPrlC+nP43EurNxy0U1OSsRGRjlNns1DdLd66n11MdfBMpEETDz
lf/cbm1wUzoJChnI1epe8qigJjoznt+kNuRQQsaugTirJk26pw+g6QNRzNYhJ7G+
QQwphA0IVQlcHJ0Selqmc/v4H8UhDcKTlXWI1+6dOP+lVR7rkyPxfeT6Izroma4U
anjGYzvZyKoZ2zMCWjraSZPBsgICHyttM+E39FHGatWh4+XFjbLMnGDhm+sIf3Cu
bMeTO8+ciNUvnBRDKNvEwVWkY101HI6Mbpjbqq53Q1qiHnsPUGfqbwlSeFVawzhF
hBHZkvwnDLGf1cuRmwjbN3OmuOUGZ/q4I2zfMbO2rJhvIu5tZYWk8nDQvfYI5u0K
tPWze/4BbS1P7vfft3O6dfdg4yGQO8D7vzK8nAxVkUMAsWTpB2qPGfbHV92F8+Ql
osoeopEaUptPOerPGQ04gzkQyPPtwP02qDpM+DS+D6fpIeSi8BPImt7xWPbI/Nm0
WzuKPru29oaJ+N19/DnsTRDyDWe5sLNn3OQd+u/LDm6K2lHv/rYixtwOrOuI5h6V
EAcHUQZyFNa3cFghmhyjDboD+QRlVg5xqwisQ9TGfdIxlOabrur8r1ZW4sU95M/Z
y4+MKYYZeek3NmShK5eXj17bluWoxYKGV6iDwJ6uJJBpgWdewhyd+RnmiqVIX5qB
hhMKEX58V1+v/kX6qPP5ZscKplDLQqlsKdpWs9cmDx1SlKECnQ7vl2v2O8tRZQfR
T1afgdL8k4Vi0dRDVDmYo18jaPaKms47EMnCNE6COEmt4kPEraH7iwW1JH+9jraY
0ZHQwpTOjY7teYyb5CnJdujbX/Ooi0b1u2afRqDWnNqMdg1PMLDi+b6U+QLsZ1LD
FPP7EUSPfBTO9d3tTIkzYyawKZdMU8VF/WwFx6jAEuz1vGcxHroFfDGh0klyTTGe
zM/GVrsBCuAX4U0U7VKjxxU7845rMrtAm3+iXtrOH8wNJlxtgZmTqknAt37GTFJ/
Qn/ZyqE2xfUUjSMaeN6fbvWAOwBBZdFsCwshJC031lq1eL/JPY/Dhs/3FWIWwj9q
tP2hZD2SkuoBDPEDkHafpj1SVVApCZWa5rU0wfOIOHg1m6wvd2RN9hKPZ4kp837B
O5++TKfywYK1FDBoai1D4g7OpfnsboR4QunlDffe3OI9lR0mYqgKAc9Pid40WwNm
32kq+KHtI6W+r153KqgKdzN58SzW7gM6I0kgs/tNfbed1VjxFqmjd2+Cyar/DoqY
/PfJqkKjcBo+IDMg4zYuveInglKP7nPmf8RchT2RDZxLsR4oqBW/QxvefqtFSRvT
VCQAZhWSN0f5rHASXBlzc8GG62U/82CPgyc9J2P495HvETRCsGOZbQsb78ccWdN8
oBifn9xNxHfPf/AqKbezbKmiB6C0aON63HELLybkimV8HL2Orqkwx74x2zi9R2UJ
VJRH9PeCTfoKUINFw9wGzr9Gq11BuTsPnGbnuIxc4y2ehimCQ//EuHaKbcDUNCCI
3emr14QzMDD/BZMh9jt9dH5qVvcF1sk924yXeuV9lLOus4ILHL2bFUbifyF9xSeK
Chjhka9ve7n+E6Jong4gym4c3C36syirGYXJWC7vZ9VpNdCkC4uNRDZvuFCzvG5R
7aIz2aftDFAeDm82OUF/6vPJyuSVNljhAVi3Tjsapb7YSAI0wonWtLhvmdCuHJrN
8NR+uNPS3yjkDEZVQxtSdc00bpM5Ai6rBIW4DZ/1LTjfSGiO9eZ0wzMCNyp17uVO
y3xIpd5HrqzydO9gRUdZvkFxfJ6eVSNXuFiN7UJehgMJLyJmMfKmpLrTy2vQNS0H
msWhbBrlozgEKS9MEC9vuVUBOiKxJncTVUCiLd/AQFuAYcc/TBaWeP/WCT0KGKFR
wy9DZXn+6Kd//mM7TEiRMqgDZA4F98HhUcoD0c6suLh0T3PGtobf47MbUzX7dm6B
46VoXqgEvInNVwx1qCa1addjOfQWQN0KtWP5o8mNxo14CremiBODJlWYyRRkaY4l
vc0/+Ob5dZX79Kc+21LAUaUYMkanSiE+fOQr+9F6X9hpaj8mAtoyuzdRZP89qAVe
W0LVtPdr0IEJ1pbNUwDPVNUiO1h2xrctpu2mgNzfpN3YFlyarGJ/a/1ERTpDVTsH
Z7HwiPXkjMK9SB35BG18Zxn2lAj7UQZ1R4yLbgZtXU9PROoly/qL77KhhnnQCpsa
m2B8CVmHrzFkDa1I1ROLKslQrmRLETXfA+gKUkifnMzQOHmJwudF9XxyasELDC72
5ZQW1gTQYR9uwbDerXIKwHRUx7e4pMOhgYvNPVmDSNIwcZT6nWNpKUHAKbzViWhn
aOOC9k33zvOYT4VkTOYpInnwLQNQEGg4uEZ8iEmzlLCb5iHCwa5hfdo9rOMVZIEQ
CvjxXZRXMhnFMJ3bCJFeG9nzt5OisEgnCo9RQl3Bzh7D9AMGOd4MUKziqrPngyLO
TY838MY0lAfCTQfVbZpy+rxSLt63wCAu/3GUBzfZr1d6ItJqgx5PpKiP+PKjjxRj
HLlHeAG9ADIt/8AbtaWoN9sat7ke4SXSU6nrzyi0sJrmWjA2e9gFlsWz2qzMpX0d
dz981K6ZbzSmAijjeTom2yB9yCPxGFtSOjwC3PTUrO/tVCWaWaC9USdoBSdKjyQw
lRLpdMlYbZ+AnMfwnNsSJOYy3GPI5satFaH2614V0CAu7Z+Z8YJSGKUJy51BbBC8
vzyPvq9iKCM8KWqOnuLkrhANox68pTv9w1MUA8xf0kKSBtBWsVJzpoyABS5MIdW9
+zvPv5Sc0AIVFz7ZWwlZG85Ukzvw9hnR/382SbvRwT72c/D/p5NcQoRtLTmkbpZ1
74Mh469gpvCfAdZXj9qU4j68hf57tv9P9ZrDk2Fi9jOAgs4MQwi9kcEzG+RtWdGV
/IaWxZG1vp+F4/Ldkn9NlfxRisWoTjmrvvvNHXFnHeVfIfOfZ4Pd75EfUIJtOz0m
JsaO5PhNKhDIDDvSQYNy1/Ed9CfEagj8s/pGXAM+o107Zq78sP7ov0ZmMnIgW4U/
Ca9qvs2e4jXdWY2px5R8ZMjKkdnkqvs54Hi2BYBweO3Hx1irMZOqu+7pkFCYZg0/
NbdLFquAPAYo+xXMQ+T2NDh446at/I93hiMF6iYTNWWxToO6YOyE2MV7fMSbn9oU
Gj5N64QsoHLD8YDVcesvg5zCsxIsYwChnT/iDpDYqCth5QNsAHN35nB9slzZYxfO
zYrPe3nlHY8Vw8vJA8QqDvaPqPQUdr1iLfQ9xPm3ILs41H1JTo+2M8wfieJlPQMH
9fv4iLBfZdMuPZVSQ+FZZ/as1BjOsTY8dhwucKl0osZS+wdPoNzLk32cyvDl5Kno
6Oha+03sjYBEDA9zZ9Ilq7buG6oYUq9sF1BI9vglFdF/5FJq1a7L7+8GpcQJcSsA
hqgzEz9xUEAzczbv7lah5SNcry4qHXkmYq6GxvJFyxOalnq+6LU0wgsSFRJu0SAU
SZHtFtT5U0cHbXQDmyrfsp8vYkeKzmSWHsTi5gqgZQflAWA7D1kDPbD16zoEMTZh
1w0/dAEw31Dz0lg8HVXXCWj5XNpaSB9h7Y8mnP5ShlPoZjH5UHg1Oqou/ipbKOSX
ANhN176FkzH4loY7RXIqc5bJSnIPrGfnSnSLEOKnnXrhN63SBu1ux9RMJ8EtGO3r
kgftbC1PV8QubN1XpctyfSkx2ubDh/cl5fK8w1IEadEdnMgagJjROczQ5nOpycgY
BVsaZBHyyLXI3Yg0eBo/7qsP9TTs3sxVZnMrcjNVrNOQiRVSVrRvWcKif4G4yVrx
GTHfFvlQ9kF2lfGu3iGBkDPkX0hYyPy/C5+ZDDyh9U9Z7WkUtZso7Cq2oYaet6KD
tXcch7c/On5QyvHpMES0myzW6pMUDhUJ94swcKmrfRJ6X4WlviorJ5xyRECz4bbZ
JKSc/bXtHGeBbwHkYaJXgr2iHe9xD7KaSV1WgMmxoiH90R7xxgavgj6wSzE2ZNKF
GyI5YIQQh309elCqFj2uewgN+pkt0sX7tbvD5HHarDWLDo1CR1i0eAvBrUGP+7Ya
Fq/XgFawePCx9jOL0FQtQ+lOipjsffkVm9bzLLtwj71IbEs4lY5HmOOYOjRw6E/k
VLCuWu3CvUWdvGyXNf6Y3S/Jwgoy0rmZrzz700OBx710xLXKiFV96+LYpRQ1hFVM
TCOLIKAtTzF5UK+mCk0gj2Ezl5NzNpKzRg6k4sOvdHjb/dxv2Itmw+JMXW00wZXW
C9Yn6oWHBJhiYYOaXYrtp/IbaXUPUZjOD389TPbxdAozemvmdUIu0YMruCoNBpba
lNvSnhB6X9ChFy8KAGAH/DhEuP6KqkxZTqeq19UGp/E/3hSbTSm2q6ZX/kZ0AlQZ
muPphWK+yC8hUZ2dvQ+Xga6XHCCXVSJrtS86xsJA+SxJee15DicZS1JasY+5jrTW
2n2tC7ZSCGFV8jWEWbwcd4YGYKmbD34ckCuBEl/C0A5opqPhUXyOFrV4nk9aChNt
7ZMMVO0uzplr5WZ3MGWFIN43NuwkkbP6CAy0sQj1bOEpqn5ak3jfpssosSdFeDOP
oiDjZE5MsOrSad3Vh9hircJgKkVLWL0gDznOCgWrPueCB9ketAQLyN3qFAToJvDc
wS5TbLZmqcH6mwIxfF6xr3f7+IDfxVcr09iL4vhwtR9cli9jgOY736U+KXLdUZli
3F63A6eERxxfnbEdtbZ1g968mPT4IvEcg7P1YjRQoZ16wo0sIrorkIfujw7MMBp+
vNlKDGDSTEgOu2CqHbXHX21SAHc7c6kxqIUb1g+agCJnyMjiQ3mOOb3CwZ+euFjG
3v9nLm6fnXMMsCCIJi56Fpx0ApK9QnzKL2Hon61nGhenvhZVntJzpErvIotx/ngh
Owq62OMNViIbySdjseBMzEi5yc7z3kBn0UFjXS1/Cx5xdEUZZ1V4v3JknXJrA3vk
tMlPzg3Zs6ufNhaftpVK8GMtE18V1j7Tm8Cn/gNm3DKUl/aUtQPXk4DPnn44tas9
U+lSSq2+M8VNoOnzf74NvY5wJto6QHOu+dYE1/Ri61vTA3FF2NuW3DrcIdW0z6yV
JXxFQn7bdCzNbMPK/gzDHSw18q6sedsoqw4CTc1EiF9KCZNc4KeffMggUpYrkc9W
fKxCpKLGCDgv4Phsrx/TuAYOHwEjC/ISsWT0s7GFcSw1iieT44FkJf5cMK9dVRQI
kczL5HHJRDs9pOXhJS0OFAt4l+ghQ0Rk1TEJB6ogpaOIcEsjWS5FWFHH+mol5yeY
jXV4//StKVikmzajURhLWvF4jzk43qnvqxvDwr6sxqOw0khpjRTuyiheZlGG0bbK
3WBD80cX+KXKLHHmTlZI86OpuG9jC9NdfVj9Bk06caHzua2AyCc34hL6q2R8jrAl
/Ic/IvDrGusSliZUp1i73+7gTYiygf5KpUfj9uePRN+EMLYxY/23yw4GBl3xl2Gu
kJEq6wRG6PIm3cOiDWVfje8Dop5z5vXPJaeyvXvOrfx0z0nZk+kU1lBuiMTgt7DG
zuMqluk3v5pEYNDzimp2aYG4G/Fs54KgPKHf72+avqbSUnOPESHuby/GhXljA/Ia
SYl8TVKCMqZkyn1Meb+9oAs86mJyBPB3jJtIP1ddTwR8rxWUXF4le9+y+aLxCBQp
h6KxEImhlHK8MXT+qO9c5yMSZY8lbHWlanwMUZ4hJTU1XI3SPGekTle6ZsZgHK/h
GC2KxiFLZVT7E5gOgrTL/Wv2eMLmsG1C2w3l8hrRXXo9EsRAkhffmV82lg37Bdt9
qju0CH06YLXFxEggg+w2dLqzeof9K4wJzj7TQrCRfyMJ1WMaMcQRKZyKT9IQ6Ia7
dJ1EXqfsc/AZ+6IPfaaOdiyp+iV5JkpiFsuPIlZmCd/O7hG/5Xcs3UN7lSnE72Zi
wk/67ImGe9sxTHf7OXTKxq9FuK4nsII9nfdXngkqVC6cj2G8OB9XPnBsNADvXftX
pXVMxbos4zdmMi6DqVMJ376nDhRFxGt1FbQ8GbKf3lMP06gnoZlZttQM/0lDCk8v
9yNG1oZjqQJp/IupRRaWXz1ZGkfnJV7jkRR3HDOr1fOYZfFpI/ZcYcR3LQWMDy32
saZmYLV/tbky5iJPejHSEOb2ALNREzHsx3+f16X3JFUACufR9rlDu8jGT1/ZzXbO
IyJuJVf5JWDucFC2R/Yp6EmUT2LjMgzgcSKeajZRX5ysLZOfA70r97SnoFtMvMTb
zjVcBFAXMMAJ2PKVK928XgdE/WGoZHp7Gim9NCsaUU07GQloi9N2thWT+vZBBzMz
UEQGTmKTkybEtZ0WWXjfh1/tGnP+w1+m1w9+cPQGp0lTfekd3WYQ+kL0Bmxzo8TK
8WpMhsNaY41lbEuiq5E9LlcNHA+Atdgc3CzbkCFzpeiCBPUYLcE2lzUevqjOrVMK
bHJ2XQDR81oMOr9DTmVzBPh/EHc0dSnRd1gVy0QAIQgOBWZcH3aYyrlqlwVulYz/
VNwF6BbCVg9eqgOMxF8bnN+vIp7nV5S+B+imZ4HiPiMkl+3YwTg+URe5XWsKSIaA
dn2mlF2W5pWuvkxdbMmTqA8jvhtgk6nHC5XJ/dVFLTbzRWTXD9Ty/3h5eZgR3M4b
qCG416titUGc3LWv88xHrIedUDGerV5BTiIlQnXzLfIII2J7KDT+3fpZtNZiQy2t
IgEJZ7qU/y1WJHqCZ04eeIkBYuTU77QET2GGClZ+/b3nE2jikjcRtXMaZNSomTSx
CcoOCPiypCzNWlBzzgeKZMrjoqmdOw2mg1zG2WewhMg+dioOXGXDT6SCP11BkI8+
1BcZuYO9y3iIsNjjKuzuuLU/R5/MwT1iXDEnrX4KWLSWI6+XfMl0DANR2vvaYMmW
JN8HdgOvUhj8e2xFwVhd654wsiHprP2n0Jfzk0RAMIP9rk0TLBtWa5+ORGOsAqJU
AeO4yxtns21CO0dyHdGZrNjT5Fd667QJ35duxrsEFAmDhaKa0CI98QfmjXAjsdPJ
SzyWWpY5HgL/ql+1iEtPhsQSrDTOOW9y1aJr6whRh0BSOLuKoF3/pWOGtKBJN1+8
M5De9DM9qeJd/92e4Vm6YWuBGSE4ifAp/wUv9z7mqtoXawgxGZ/7esPApmFf56WQ
S5DU5We4VQabdnBDwMy6iRgwpicBnjzAGwgrvhIRtASdpezllwWptz3keGQ1U9CQ
QAVtSOR0V23mOY/sANd/7F8UriyejTLpVEwaEdYhMnh5OmvAizTCGoR0wpFUej1q
NgguX+ozwuiSPdoE/LCU6XbWL3eWDqjP43iqGqMTV8MEU+Y9kek37lwqfEF839O8
8UqtUTwWV1o5rjBODjY9nYbpoGKY5yO+JNkLOHyZVXtXQfaNTmhV6Qd3xUj3X8HZ
EOMwZf6vyPyhw1s3+/AWpvX8Jw/rGSPuzWvMKhjVc9AUwamxqWt6RVp/xUdMRIuB
BuBiWH6tb7jqMuOReqaX94Nyx4UeupIUmuJ1c3geUeuBtnIeqwEPA2WBmQcGZklG
yfqpMWQJ4b/vK+qjUq1ChOEdSH93C5fI2yrSM9hcR//X1/1xawG7g6PHOKtlzR+v
0iagc0/u31ilNwFjXpK55soNUeSmfP3YaEzhD5LmgNgXQ2ha9exdhKr+XRFBBCRc
J8tSu+Z3qCgdbSf11kasfXICLVO6YCo7dnJNnFB/khebqlmaacJcpH2sVmfp/ISK
lm3V7U9P8vSEeZ7JoUeF+4I6AHKr0QvvotV5zG4nhPBgycTnNnPnajv9AbI/X4ar
kq43JLooPv2TVkWBVG+taXllRKF6dYUFxNCUilXc65igzOv+LsI65Dw6ToMwIQfG
grWfV6negXCkH/sNjZB2ImcO2iw0Ha0Aaw1JsTB6EqWYVZubzZw8/dPICU2HUmOx
sXdxa62aDCO5xiCHGUluSsXU66afn2Ua1KXVY62d3QlVbD2HAbDrFI0QDJhikgfS
GBY5G3/IJnjpHDz1xpt0f9dujmoR44HWLWb2+mOuXXCZo0M/w08owDvN4LjxPo6B
V2wTBhqOI0OTjBrY5NGGb0ZcQtVyv0c4jDrONZaR1Ius1X+eMu8/3dR+LOy8OLZx
IPKwNtO8MYqL5ulry+mh6QCnYUH+Jm4FubcdEV/L61Kx+zLtXB5xjpDpdX1CXavt
fikhZTDBl8VdPs3NhTrKFQCxDpjQUu3bbrQAZxfBiGGPu6ErFMb/fRF6XjoldHv+
cUAZM4/yeV19l6wv4LkAapoWNPc8IyDkdICWhDIQoUJuP3q25h+J/zFtVKGGDL2+
MiSxqTBEVq9YgpHMRNtCQ7y0fM+0hystKD5UtV1HujmNXdo/iluS2IFZfq6gZmwP
EEG42nq0UXqdaHX1K1VfZ6uZrLka3cHLeji8Y9J4uIlUTHhoC7e3j5LvjyvO1OKx
btVTwM8ZT8ZHEZJLp8rYKXB3hxB10kK6ibaSN2I86zMXaYpM5qHYkxEqvVF/NR1D
aGGz1H+xSLeadIM+3RFaxPnPeFK0cGCXukvth3jPe8Qwio3teVU7sCYfpQaR9CIq
lNqLXeCnO35bDjX3atTbQPcgYUHU7qf8yuD4asULkvCzv9W4XGgQ5wcXfKFWkfwP
7tfOblF5AwFdc+9LFFt6aEstuRX1SKuOAqxNC48/AensbH9oqLnTVcxObfqUc4NI
6bZwhldMWkmDcpcFTN0NVrOMJQ+e49Areh6pbfbtjHhrO8fDt1KOJ+VmDYiEFurZ
uuU4eL8b0tDdhX8UscnGJycCkXtmsrCiZLYx8jGVouxygaAJSpk+5HcBzv2ZlQrP
J6YGAw782WhJ7vxSNXK8zbPTxvSFMwrSCct76BeuMQubDhqh3WSwTlVFZC8X6QmC
hdB9QkKQ0FOsOHdaptZ2EzLHk5VQrNeXziSgTygfaIUY7AOSCJCSm5mTzoiGqbON
JCJ2r3H+jBvdpvYu7ElISBAmsb2g8SWpAQYa2Lr6AHA75hlHPUdC3dGJ1RGeEV3Z
CddqN/1RWVaBTKS+ymlfYf/RI+l2F3YjVyZENQ901nLiAtb5v4660xmr2Z6WD9o8
vYQ8gyeRcyyzxpUFBqoSMAXu3xDDuaYlIUI/sWeU92UhXWOwMcEdzs5hHrkDCAEZ
jFn32EPdEzbqrLtWBf7HGodegRX098oCd7p9NJAfhiz3A5GirLbPbj7trDmW2xqa
B8Je9XSjMR+qPyRB36IbpyQDl4VdvTfV4nE+IFffvixdVkPMli0SwfztH78+eOyC
c61apTtcwRiZhwFHFXG1lBt1AAua0lWXXivbD6KDzyKi4NXhRpeEMmxYwy8piB31
U35R19vUUygMyjuU0MWX+LXc81hmmqwNyyp3MuPM9YhER+qwStQ+EY1zgjBrwszQ
C1vOCDXuHsEMca4DUx1d38Wse87qbF58lc/Lds+y97o5TmMlQLuFrBNndFKcyUtW
xm5vVe1Nx0XTzF51wr/WsCW2CEmdZ0LEXvxckmzDtEW8A6FlqLJF2spjKElbDR0J
L1heRZlheBUEnvuKfZH76mfj3mJZxnoBFYiy6oRE4Fim0C0zLu7mPMi58dUAttlF
dhqTmynlKlQiATxUt9vmmZm51dqgk1bkKfJTQyoM+IOCjjzIap9nc+icMUEU+Bkt
ZBI+7EFsSdRUoZ6Poey4nFb/CDFZY5on1GC5M5egMhhMNMXZSeD8JLrMKwq5q/lp
4MQJmqsiz5Qo5iapW2lBtCQLyznC/kMmSzujI1LhjqpXJ7qloOf9ib3oUdSKU5O0
/3ZDh6WBhK0Y8yVm3yjcAhLMdZdJojEO8QrY5mLWz8xGFVlalRtHg8WHDikbEjYi
8xJ7nDqEWolrmNmBcl3iloyJ+uSnNC+W5y885Zmf4P3MUqv0hZ9nYD8sn7b7Ogul
BANefDTuCsk3zRHQq23iZlQ+NcuvsBti1wQcZg7cLvusf+reNsdCL46YGNo7fDXb
KgpHQrOLw9i+Q/E4ZzSRaJH4sSBP0s3aoPVK5KNF4HRdhsh7WZgK4hTHt9gQ5fLs
utwErZCySa+zqy1nuCPpxQWbZI96WptICXsTC3b0R/o6oZ3gEi60LCpOHGi3WNDN
YfQ636qkOsnjqHgCtxIIu/HnLWauvld+LPyYlAT64izq2WV0/Bk4K2M6Xd9mZvmq
JHSjLZK3eN/oNCUUf5106VFc1TK5Yt+Ay7Yms9SIHXxaZrtTzcpVNAm6/2dCuIsq
5U/JV0iRYewGh9hu2IVIEzlJrQWgV4ZXuo6UNtmjmRWqGFTYUs6bvwKMjU3dsmKX
ysXK9ciuuFHZ6TEOt12yX9qGT49H407ZNDc3XJk9fDEMwQx0lpxPjptyYkafouaO
tD4FEfiKqyuo3KqGzxM6dYHA9cUZkVibnPkTrId3u2JYy9Nf+5GwOUnjbQqXvzzW
TCauDMqsqGpkM9Pu33hSBYS/hxJM2DnkkRj2NuEDUsZAPhF9Ux7VYAsfKc59pIzv
wk2VzcTFKuBz9k2Ve9w6LoynstA/TyPRGmte4oXMG93JH90dRiS7jt1iNF/Qk4xX
WwxzuAERcghfgWbrhjSqmUE8qFG8063m+uILmTgg3Ylxo92WYtzzDIIxTzW6lZLU
i+DcJRCbVBGtciR8uum8+7Rd9SV1tk2IHXcpdfk+iYWiryDSAmVLLtHZKc2ryGh3
lN3JOGtU+ZNBsSQhE1Q2jELbIvFj0X4qXRAVBvaKf3U80vhdg/VIt6fy1iyRLPw0
rUfmk715tvHRqXcePJLnXTxl7BZSwc47LrCw+5WNUm0ezEWF44C2Ei54pVyJQ4cR
2KsTRxB/NdjdRv/hoYdLKMDflkobDmntR1nGVu4gfVh7kRt0WNqZLd44F6Uy3U8T
ZAxaLU48c6/R6YlptMlkJLQyMaOxDQfxsxk08aGX+V0Tqa81XPaRfdH6TF5bhm6z
c5u54pQgDLzp0XlsnoOQTCGyN/ixQryT6rhCJrmmlv5j9tJ6AxSnaVtzaOY/9R8w
fyYVllPRoEguhYmgsA1D4QAACylBMNbfXpGVHFj9zBqVH4gmDCopQp0gzX+ARK6K
Kb/EDQ5Rk65utQqFdNfdZgkFAvKxgEdkRhB9R0+dtwJej7crfgbkfPATYvN2RG/k
EpyKpGGmy+rm5Rxbg9h7jvi466zQX6yB8agcz2oIj2lLtI/ygugdPka5MNtyK44p
gyLVO6U8iFYQOQGd5a28TmaZv4c9XMJRSjy5/Skvw0mM7LlpXIlAkfD0k/fymTRZ
fNJoouHAPyCxAoSs3W8rp3+gdNVjjdAQYL5ohUemghPevDhYmjitZStWlub8dYYJ
DhMM9WEEzmOfG13LeTT7DJIQD5hAXxLkODP3VRubTUi+bHau6uQkk0V4DSyCXpwn
jLgRpHK9h2nM49Dj9csuNYmWrfKoWB/AWDmJq2/kY8Xe8rX73U3JdX6i33zR4/9Z
TB+dJDrZxl36W8LRRI/uSbp7NrpqLLMl2kkJgukhJMMEzwtk+sroSwtYmgfhTbwo
1gX87VohejyRY8a5b28IYCquE4cbdi0YpR/4aoG7eDzldpzjjYzOj0BTQ0U6AX6C
jKPN8nsA/7FDsbM2sn+A1xz3BkT/926HWs8tEGCwxJ9TKRTlg4+xsR4VNz4jRkbn
buIiSB7VskapzCAIbudY0Uh4OpzT0FAbE8znw1BA5mrOEOUpoQwaAL59fauuNWu1
IXUjAV5EAmpoKJovxp1WNgHhQM7eOoos5inescI5pUWf/p5ahrSLS5bIK9BA6VvY
j2y5ZiJhQNaqrvm6UKH36u9nyE0Vz0ffE8NAF+qlIYV0YiJUE+V+QfdNJ+vgzlr8
/salr3R0m0gOcdtDA6BM5uwNr1gSmQ+6kQfWiQvHUSPsb0XC3cyy6gtQlfQrSSzh
K/moEv3pUDoBZxFJjOAV7VI9MwhGCG4rCLxb/eas/QypnNhGTMPn6gaWnafCKuDE
nWD+A4nq4UKw6aRGev2w6pMiiwMFcR4zDQNKD6d/mVJlsYZFM88HfNPjszQrj1Sh
Z3gMePMiE0dIaMA0fLIjrFcQeVl85OYqabwfGVWXey93CDTpnxkJDAx14U306h94
YBnmMP+KqvMSpJZk9Qv5nlPc2BCTDPpKJR9c7DzVMqQgQALgzEz2v9k+eZVY2Zan
L3KpGUCAP7l6SO9OJ7DTMKQFPD+9hDh2h0LN31uZebWbWeifoCpxCGaL7Ofnrfa6
lMTEzL6mwwetIxJ2yQqJWKiXdqWluQW1aKy52pT0LFtaHg8xhFgs+GLZrHwT6LxL
LkWBLNIapEgXlsCX8MBjmpwYX1b9UtTCGyD6rCkWzGdhQNaL4twUFqmvV9vCoH7O
6hiSVyYxORroDbLIH2fTJjFvoF0zU6eJnvSEBii//TafoB+OHDvIaBgN7KeVjM1c
EgioKHeFt0p0Q6WsCs/HzfeABal8KMAZUHjWfqMfySul8NYia2h36KsvUBZf3GlK
RaiDH4cmkyvjbeCWnI0k05yJhzEusw+Il3L/yqXwH5PUloWYKbBxvJ7o9c+EjpnV
vYpafxQwiBhD1tCA53UuZ/Cy9dw5vYjZL1yXnt/uvJMCq8+jGr+xs0XvqJC/PlZE
nHWC4vPA7qLcJSudpf+ktQ0MFjQ16if/lO6O0V1Unk2CayxH3kR/U98Um9xywcPP
ubQ5aDWONzreAE7chfjiXnq4iQ7CK8hSDkdHFgOq8z5DnJ8Yph/ej9i1IJnkxDZ8
/0vGY/3/80ghv4gPHb64ccnLwZomYF5RDhgb1PgQfTChuhdfWqH+32OTkX/yCHlA
O74OZkQs7EBpZJyKAY6MiH3QojfwNsocZvaml+iCh/ZXLuElV3+YGAxV8IHCLVuV
8u+ke2uV/Lk7TPGAkHd/rab5qIpNLo80N2e3Wm3lgYwNZaJI29IGSBS03eo5BvXx
W0akmpQVaA/XsAdqO0bLV+milpoeghoKSS9hTrDGHHSGO2qanjYf7irj9sH8q4ny
S0yw0lPnsO5Pm6HjFJ25MWn//u68VFBHt6rawGLIkcqwxy0yWtDCULxj7Nn6/nzE
fzT4PcK28HWgG7YDNpKJBujxw344M902jjaR3ZUgo8tg0Eb6lAPuiKpg4MbglESa
hKBCUIRuJZuKM37/jH004obRmRjPYKlLEoVkjxMOurPwsA8ZC18JlddxMZLCzLT8
L6PFwYQHw85jXZwl74EHYr2i3hMaqZcwFrb3fusgi9Afn43X/yiG2ErQJRA+IFcs
s/hN0zGqVOW2ZZ4+Eg/KUwRV8LAvYLKOnGIgZ3FMgrAt752ZANW2WyaGcUGpEI2b
IRiB+aMOpdxdRYe5+T4qykv2HyOAV8sHBZHGfXUm9qflMx7bmGYZcunzqsh9dF9a
b6WaQ36/8gjL1Ge2iGQhFxvW6kVsGS7JVCDyPzA2aHBfWn9ksCBTnOd2/qx3h94f
oWiX6/Loai7rzRAqEPquYVuO+vSMK/K/6whyPDUYX88bgB/Ukb3ONEEtmgg9aeE2
YwVFC5c5i1l+9MsU8yzuBnyWROXour4QBXR9odw3kMxFDPfZ3nPxE61lYOTbmp3h
/C4weaXsrWTj1umQJv8prNFovsN/hovTHiObPN0Nsak2nZHVptAMU6TO/gR2vVnd
9+9XbmBa7pVw4VQGMkeY6Xo54csluoKXTK58PjKgLjkKnfzMvFP1Dmve/3nq1BbT
TFwBX7P2vJofc8Ql+hom9dHx5D+1DKNzyF1v4broCpXH7PLvemezTxIJHMpzh3oL
jZyFPYmdHKM75yie0R4+Y5uwERiML0ZjrSclgQllvukypII32mllVarOKi8KTAfr
yNcDCkACkK+31tiZSEzaeDBQGLmra5kgYNEgrWTQxEVkBtzUCyTH8ntpaldInVAx
kzZDpr1UjQyneGb+5aP38m+pGt2EJllBNZuScIHXJdCD4IA8/zgY4RXInyy6jEbD
S6MUvaDMokUujm6nEg8qDbaiJ715w5Khunw9KcYXDSk3sWaLxe/Te8RcqoMQQzGt
xUK73vc35nhTsRiw+gQUVp60byxBdni7aCUaMH3RspBt42ewB6UBm9YNk2WUdCoJ
vFpstZYrrzf9tGJVMX+lDePLj0gu4kfMwSgbrZ2QcFCXsvOfSsHjbVZI7MeF/A8V
vZlWL3yOyEo5aKMF1u4yF8eGVLRJ4mT7M4/Z/ormpW+Re0WHE+8se9R0xSmNtg0G
PyYXUHbt+3HIqqAV0vYlfMa1aKb5wDFNCKZeltfx/RJ973k+7C5wddDGOoGETcuN
HxpnarphZSmFqORxbFNdVROcYzyEoB3BosuLgmQIjVe/QPpTOd6Qf6fm6KGSo45I
NnBfVJRbfkHLEhAji2aq331FGabyj1GovhLPLWltM31Py3TcEZID0UR5+f6+WQ8e
QeFHvaQzIz5O70SaSh+o0kDbxfP7zEHnd/k18GsQGc6O939uGAvCJ33C/jZrzVDm
OObq2buJo8WuWZSwuk3gFdLhZMIQ6e3zJmiot0f+WR34iEznkTfx1e+BmMADpHez
Kim6FFCOJ/o2GH+tgTsoNuaFdXcfHl3XHvkyve9wFgpRfeX7GISHp5C533OC+hdo
LJAkWU8Kfc0ahb26ZHKq8Do5pNDsh2BoMXZ7uZ4rRfDwiIgxvKKow6IJZfRPzBVn
C5u/f8QTufeX+294+ncI8Js108ZV874WxOELobnUdEEHFZUOUa/4Th84evvm3dI+
FGuSTPcVHkk6Q+lzxHzhkZi8sP4YKiC+earUHsT/5lwuMDDE2VAtpixHrtmyOgso
FpDZLK4F4WxWytnwXv45uPRrcjci7ceT9BgkZKgH0ijBtDYMYpOoQRer7xw5/OWe
Sl/TNcAg835HZITtoeh7hgwvq6i46R8iupXEWTQvnqO04eHv5p4cZOS5hAXJm7Ui
rrog4sD5TDzk6eMJU1bA71Jg86kaq5oQlXIBosnGqGBrkn5Z5EWRxG5rKaorWwIx
z2jmc6JZ7ckiJ8xQBqcaLdiTwneUJeU1ztBiV/Zk25xZS9oF2CkTnBTj7+dnT5yc
wSHpFb5Ctd3EVEoMMRPnipSfpM5pyB4xUeO3KJNQAQUgmRE4Gq/t3DYpyjmdemkd
JAABq3BuXM2EwgW4L07yO5YEPFZYGuqPUAaEzDYF9GYgpBlkNG5mLTCzKKfERDo2
zfMUdGD7azx4gwdxL4oJbz05x+9GKcIN55OxdyCFZToVUWODHCzpB7Gd6Br2lISf
KmndrPSs69Dsp8tq0PYclWz1ZLtxNjEshAYwvX9LPRZoEyjK1sDiK7qCVL/perbO
n2Iqsoo7hHc1n98busTD5cRsjS/Uzcbevqm51h4LKvQpcUlvzMjZiqcPFTe1mpsT
JlwM9C3fzVBztRNGsjtpKiOrkQJfoKJnotOu67s1PqOPhz5Va7QuDoAeKopeuRS2
+W979qzhQPrMJJ9DVc/vVmebQYKoTmNtBQGlWA5RLRohyb52n3HUFogvc8UcAUNT
6bGKqgtyGylRfmj7+FqPbNu59wcPMwun2d4MiM6Bdp30+Pkh+ZAAaLat9JKocVBO
VPkWd0+uwOatIQ6aw8SAqP8Ql86EXtCvpr010hZAwyRFiNmbAv4K5Sj2iaNfAc9x
Gkx2euc0eLIuyWmEZqClU5HcPAGKl9NPN4SwSaqZEBkWhq03v9ISic4MW5KecpFe
kD2pRXy9EktXxrYErubVizb8lD1Hb7iYBIuOhJEIRaPZnSBxgNh0aIaOqcPkPf2X
ZBQtscFDenYiAqGANNTEJt10kUFSNExKynu83WqYEWz8SOHWoH5k4isAa5599wcV
wwTMz/onmrFUpeMayADK6T/WSNdjKpI72yLYgPHAfA+yT11ga4MDP5KqjskmKsIj
2UstUzHtlYJf+odJYl7OO2FaVtE+lnfLO4givs4jh35vDHLVmZXOwobVXPo3kvw1
Q7JH30LEbeM4Nq6TAe/yoSXBRWm6odS7gJuyz+h9wkqXuZHJmOmxbshAzpH8Zuka
7pEQ/llZNZ3Q35eCLNGI05xHotP1n03KVmku9gsDOPjDeZCxGnbbo6J+jGtQdlm+
geKD0lCv1M2t4dXhK2eKmOnXdL3dwXmW8ShxFpFcjYGiFcpYIs0ZNnZi4lVvlkLo
nbTIUQyR2ZbiFVqKoa6YcxTyGKfr3ND/s+UyLEqlBlLHeLgJS7FTaluLQkey5WtL
aMfMuGw1iuDgAgpsSGOOqRFrM1anwgUkQWBNl6Ra6zd36Tkp6jG9U8OGdyTL8CAu
tHzqwCRuJWL7/4K/CQc2VGMC1BC1saxqshmiBpUufQAXR0sYfHlYqP+KFKFnaeHX
l9FFZ7QslVPeBeZ0P65psdKAJt0mJpZSSIcuPTmHKyAjRvFd2F4wgqFf681+xBwJ
zt9V3N/g+Gq2HG2Gs6MA835YQPFg0eGte/mIzIw5M78vL8RLp6hLXkobh2y6QaSc
wmdX5W04GduxhW8Sha90LY+Z2tzkGbBeVeWhzYCW51JsOvB8UE+0kj3GmHjL+a8U
4WaH5zNpMN+7GFQWJrelioD1RTDLTwLc28ZKTMTUrvCkAsCVF0K2npTKu6IXtvau
/11adc2YW6SVIhs/28nB9pBJOEBmMWzxICYqjPsxqbPyzahAM78gTVHJYj8xgmQe
xKhyQowywTi4OjA1MQMgoObmST7Pj6Lv50Fwwg6cndAPVm1OwuQ1VIwuXn4UbCuO
4d47B3iz27YvfgZYwpXleBdiGdtqB2vc/8/IY46cVfOGT+Ge6Y4cDVNfo7Q494ze
aGYbD4/MDhZ5uo98Ptb9OP8Vc9vH2KeivnAFwP15bgoTJD3K2v3Cl1YRAcil1+hA
Y503uAxdTfMR+LZiO/GO9S7xo37mQo0ZHR1iFUi26KnpBoK7IQfuqJRWtiwPPq4p
hAlCGe0dDEtej1DOxGDa70yMkRAY2bWyiO58wJgcuFcOOtI1bEMELaZyCnCpPNX4
szZ4xloRW/DrKswx9a9VQMBIvqXuK8z61JL4rpUvzFe6RF00MZ9MkNpBs8F2zQ3/
r7bc48/tJo5quZUgaHSt7I+HD9kaSX1tZvvhBWlUjVb+/mkN77Od2u4TSomAEAFk
4ByX1CU5Gy5OeGdo+x8NUdgBy1s/OwTeUqfpxNlOCt6CC0rgxJpqLsJVhMNawnSN
+HWLsoeXoJoffcVvWdTSniq2JqT5qfol00WpoyTXMjC01PUlB21rFnMk+DksEpdA
9qxLqy+JqXg0GAR+0bs/Ze2zHb938yOhk7Ogb49gfKpWhWp4+336WNzkLR9v5jNF
rwKyAYppaM0VU4ttuF5hKHI9G4aJjxOjoBx27K3uE78fpmTHtgh6o5i88cMF6J9Y
55VVZUy/bju7rA4ScpdZWUMYzec/C+G/gCNPP+ju6nNq7KYTWZbE+suQgTOx8qz0
lN480gc1BSiGL1TtdkHv4URk72ZnCICZgj1n/vdn0MWDqbqocw15Q3w9cVzzAo8y
dNJhlTP38Qfm9/gmeQgZexdQWT50U7cdP0jBIRFCro1CFKcplTApxYCKy5mhSzJD
NP3cObWMwQcW32qw4ZW9koJaPXw/8nfc8nQr26GbaIEAD2q4hhfIDmubWf5CJ+Vt
rZvhW1bUZo9PYeHqqyhe69WMplIAPp+oxFQj/d/Uoo99kh4od448TVsu2+xeibII
P+mqWxDsowMw3F39NOHL3WX9MMAVMVV/ePhXTxq+nQ+ijjYdqnhvNlK61G0/WWAc
CDLnQ3dJWkI2u4xjyQ4dD1K0N88AFnftGUiY7IPMdZkf7On2zUTtB7O5YW5zoxJE
9Cy6+AHzgiorNokTr1rB05ibRQHqYVn74G4nmUs/Qvxeden/9Z063+baLPpPx4sr
3saD+Mji+bN5NnJbAlieTjLXh79QSXZsUjOLGWCSICwcDyfVFRVNu3oURkC8QRLl
G8mxK6BBddTdEs998FX5JeTGl9V0D4tsR8+uQWRyuh+g0l65RuIpnkz2jrWTFVFf
LQpgQZ+zrO5GHkUyMfH20HOQjC5xst6xI0oVAcAnPz2iRFcB7QWq3xAksPXGx5ee
uNNgSogsZn7DNYXbI4BsZT6f8mT5+hqnzDQHYZatpQdnFuWXQQMYrB8YHtZGs17k
Anov9lmLyviDLwPbD72itQggqQ5Y4d4ZX20/cK5CiNsMAm8jj3SZ9P+FxqHsmKaD
PrvhdSfVmHmOMImi5Gz7948ssh02XoppfWdOKjcfYRdvGOFAYK/dv/Q+/KoqiwjE
jvyU28DzT/pFdRZTGQDqh5ozkJpIXSMOeFnz75Ruxnyemi+enT5wNGhcQZTDuP5/
g1StMp/ejVV7zB8zn9JpD182IUqokuy5Uw7+9/pHAnkGM1oOmYWSROKEYAgKSFOF
ux8Oe4KeHLSszH0bizCC9nLE2AEaMya3m1A6XMhLv4sZ47tkrHzwQfwLvDe2Wg9W
oBPOScl4O9CFNXTfjQCZq+JIRLbiOtjGjbYFL7M6IRerc0O6FapEOqRvQgUKtP/3
enHheztjrYl/Ox2DYIkpGAcVJTEe+c4u7q+sOA3b2Vuigie2ycuyO+auk6q0njLz
qQZojn29sjRhcbGslbiPlmXxaNEsNLcY3KKSsHiqo4CT10gW4XRdFC0Gqg53xwB/
yQJ0U7sOEr0lu4P6nQGfBZg6jXVBj5WMBuw/qJE2d86RpXFUbS5wwy5m2aMCS9JG
n8AcZoZPo3kTRYCJ43UJkosXG83L8lrbrd+kcp8GpCpkGD/zdq924xleWWCumO+0
D/eVjfkQBnun25xqWhvLNZEzmWLUFlow4WYaFY0L6epu1HOPwe5v+mHu8x37Sq2n
gcRvTbRd3VwpopkKseF0SjOkrVMNwCDdy/wwwuPAtpwuGY/9j3cX0wrBMDk5YbUM
kY6uey7dDADUkFfjGg0mfuCVSUCh+LHaKiKM5WdfBeRCWtESGNQlr6/tkTZF+jTk
q+1VsE+j8u8wvz6cBMD+krPlPp97Vg014FtdbWBNG8WlknoapQiiHsGHbayo9G8u
gyCfzWkfLO99liH6sk431ls3fTIGGlD1QrwTneMl7T4b7+yc+RM3fCt6tHUzkPgQ
ajJum2ZMYv6Eiji7zwbZlS6Z/gF5TIrUwhMzltXdR+O5GiD4sEOVUyuk5r0CoeGB
L4rmMbmsOR3J6BDilccLQHt+V66PNtF2a78wVHjG/eWHpm50ELn7FlpR/DqDal/6
ftXnSmXHVvhecMljZpeCURR2yw+v0PUA5iXJRTBKie0DnLPmgJemoiFYmQFQjIaJ
UML/cvGSuu3r1bGwiQtuFUnYpzskDBxFzWdxicYxSfl0mkE1g8VNYGng3cFblXI/
WMMF/iGMQqodQa10Rs2FZ/hl9JchuZ1ZK7C2T4/Es7iForpXiaZWWN4VrhbI1myW
NbuOZo7jLXafPz/QumKoOJREP4DnUj2WbMOr7UYaxkYBTJmmpc/cPW8V1+XJfEWv
B9WeZ7+2CEskuL24oJmuqK6xV/oYt3BnzTEvZttvcQMy7ubizVzfGjt4KiXU+zGu
Sraf4XB9n3S7tZMNTQ0tVtW322hZfFHT8e8yVX+AOIRhezeRQGJp1t87N2BV9Gpx
6P9/k1ks+y5+DIsCAq4n0LIEqDlpJcqzsIPMMmUpqfsLaWqO5RTWpsMpy4GPRchC
xUAfSU3r/evNdkLBQcWhmb4at+u/Elx9TbeM9Kz+t3wXaHDD5a6zBVuCQmj9D+yI
vIfgqDuxN/iag4x0qZgVg8GwH7k4LAhoFhulKzMr93AHNFBquhgRf+xl8JvY3BLi
Xm3ySIJonPhqXHypDlwFG+HQJMdUSWp9jTFVSx/QcrWTeSoVdaljlXiS80phH980
WR0JQu2QumtEiWGRilowmdM1N65k8HsvdVSx117EikLVcEzWN4F4rYJKayjbaeq3
05noi0fqkyxoybWjHKygj683PAiZrleqCHzBkSJRhC4GvZb60JtPuUfGNcl+a9zJ
obppEjHrpkUIj/2wCAuJvCpGC6R7P/G0k7n4RrGNwXyXnV/Tr6gOvf7NOIrxoBJD
P+ZRDmHBTFPvY6F/0AZCBd+JYal69fTFidtiQ1DCTGKPyAyPu//BR4jOo2G8sCgY
J1ptbp/ozOMWli4MHa3Ub5X4gWFv3l2P/jlYuwvGGvad66stjjKHfIJ/L6+D6lLp
9Dt4hDGgQT9/MmImk+O1IECulOhl9+VHrRKqFkX5bcuADsYQAHRBuah8G1L+y3UZ
h6oZAUN6f6HmEdbT1EoxTyWkPrrXjnnbndzsssCm7HxlJy3Z8O2rU6TubcgfS9iw
9/QKnKYVhtQoYhHy9WT+tlFN47CWrjbf4xFy+T9mghd4M6o7XV2sIfLvYqxVHxvJ
FSj+HOUkwU6SqTyRiZWskj0s3YLWKykdhGGfmbqADTGJ+n0g7LjxvigSA/sCYIxE
5gN9SFAGVqJ9l6OgKpB5GP7o+f4yl4D3RGVycn9sGbSwIPrmrUvavsplSpeHX2Lw
RmxvZRr2BcnJIDRe56rFPaulrcfcMvwU/dZ6F2ztW/J2TlGyInDbxfBrmWH95IKe
f52odchdVFNCzH1Ayki6wrg7spXiKFwhVPa6pbTUDCmGo7Jp2NDATzCyWRylhZxd
4lav25Atet47rDHUUXaHm/3YZKoUEFBzv+UNrhTAbO5Ozjkm/86o2c7i/oYfNub9
H/M5meHInuQTuwYPW3y6yIOT6GxdWLAOZl28xXfr0eND4JR6qSDo7HKdQ8I6MoS6
kAjkIxbFYuaYHi4JXKmbHFTDSKp21I/oZwRv/DHDofDAZ3bBWQcPqJZbfPnY/oyA
8WS2PanuzJxuTJ3D/Krdo7PNoCEo3oPFS1Hjc4gxg664Y4HacyOc52LhJ8NPJ/ng
zY7ahZvrdZYfObBxA90WBp3hAxUbI96/VZ10as2OMAF+wgYQH0eoF+Ys12fiPr9Y
34fahNzAXQq+i3UacHK+ZLmPlmErbhXWUBiI1Y/cOu7c1R1LSLVm/j1XeHfG4ozz
hxN8zFFAGxz2CJ77K4Cq/XVC9mLwrX1wwp06Mxu3YCVXrwDn2wx3wdr5MOlSqsZC
ffZLv+JDRe61+++1559ke9Hkx1M6UighLI+2CqNYBxtKCrvK1qg1u64i1PMuvq2r
IiFlt5WnixMrdaOERi9BsMIUkbgleyHrK//q1QAp5PmZpPYjhqH4N1WwrDRbj4WB
sqCqWNOoYeqaVWXZOmInKEjRxyQto70IS4VpsC5k9Km3y4M2RBqiLeaJwsqNXlPv
TPsgBYjuBSuvI1LVrhj/wbxX0leUZ7rqw1vFrDdoxMYO9Xxyrt5PMverOgmiogzb
B7LBGQHyZTb9CdGT6EJ8YvE3nqjWR/v3VQ9KAQowGygHpfjTIpPObtM0yAV5mJZG
oGHWt6mKBFT0cn0yUl3A9Ys9DgcfIpfpXzP36+jL2OXZVyBFOl5onJSZQDrXZKnb
cGJZOIdNpgt1CwJoYwoNrvDm4L4jdOA7zWI4yK9LZwM/Q8qUMCL2Ar9utcE4l1yW
NYJFDsgUGO4Pp8odJzDuhdIuwEQKf3x5hcCA+jACRmP++xzn9brezjqgeDSsF6Je
q+NjNTL0X1TamZ9Vy/l3SQTKJS0CdDBpilOPey7EIQgVcTuLO6eKi0CnocJa1eGZ
DnEhU/sDJT5L1bektQtC7AZIlFjGFS7JA1zx24tU7umRgWtI0BlHcvR9Km5S4nKY
ux/DQfTwrFk8UAqTUiUdgaTONzb1JIQhihWLXPj1pjKkRL2RF0tmyRpYxtfdoeNB
6lHsKy6bXfjuHIZ1ypUN1rUhQkhSXbeqBPYL0PB+bZONZ9nImO6UzxDzL+wU1V1V
G8dbLt1xkZWUSda2mCs/wpTs4oEIS17E9ojBG+lLtFk9Q2PouC44YPHeWS/hN7yh
BBrD2Ns7mKnx6KbtKWmwUIPpkjtzsFms95ieBgAV6Xoo3CQLXNgWAStt197BBNNq
QKZd3W+RRiOWZid0yz9FUnE4kxh/894v0g0atADAhXieNMb7ptSLtQVjJ1O9MFQe
fqNKdUEr+VofFp1EQVlu0P5149/6BeqTEUSXUnBiRrdQwKf6v9wlH369eZdn6xAw
dvaggjOtgNgIAbLUqqed2SRzC3dzPutWFMUqnHELnX+wTk6FnZfpKLc7aSTmxy3r
heWCrL2Od3v25pEj/uEwomJMMuxTTsDKe8N7uKatq5/zD5BHj7gqJGdawlWZHEX4
6KI/7SGykSGt7J3wPaLhADeFknoW7T+2jgDNPCbtVh6CDNoAy1tCinw/KBfLx/Of
HJIGulJfvm6hoxATD3T2MHbFY/N7jI2PMB8YpxVgtTp2oRfszSNqm33B1twA08OY
xhpxreoc3ii8lIJDSJE7dXooU3en09MbkFf2OC6zB2kixPEaY3pWq0Gc4GxXwisc
/snLd432HEDstATaM7MM5LbiGXdcTG8C8S+xmDNoCpO4Gc5rUYre7h5PyZVBSsVB
KOvDbWNhhHoDRwk7dVPZN4X4GGfYPfYzKKzNtTi/NjUIJnzEHm1QC9nWBgyJtiz9
f3Qgs+hEcPxgA7OjQvJxvq4wnOw2n1vJyKltqsWgn0Jx7MZFtNW2ycAbXFh0ev+V
X++BzI6ra8QPyLHfWv66Dz9gB8yFul7h1V8ux3sPp1L9cx5t8shaLFtar5cnIquX
jVrIyvpd2ZMeNCeYGMANzUmIVF3al+bLakZ3kn+bvyB/qXi+L5faJD6u+cAB5D+h
6vDx1cL21ANEcHLIqLhW0uGOtQv3uUf8r0tglz51sMi0FcynvUdy2bLhksg0O+dl
epuyllyxe8ssmpBw+AyjsObK0i62kduLlAlHN/OYLIV1WBIxijpo5K88nbmUnXuX
MDcBD67KDe9+p5drihIqwOzX8/ncreD0I4Q5727bSpIbuJVGWVDGbtqhhTD511Ui
3C+tS3w9OVmXhPn9VAm9DQov2UfSvvDJky5CmVJjK4ZqTdvjnpNOg3742l3pWlUT
HH0oY+eZgnO4HaAqvgfX0GSSJ5YAJtKA1O++ysu5qjCBf2/HBHKeMVtqNfms3Mrh
M31vW6K4QPECtFaPYdeslbVV/H5my0MqQS5O9JesAQS/JSBXjNzdz39zx4Hi9geu
s3IexyqQtOAOO3K6aqQTg5YERoE6JMDQXUD85bVXNxc98D6db9FCZzszwtMWY2tY
INl7fxvk/ZRN2+613+NQ4Jue6lQj9tRdG58tUYmjqVgN/yjUEYhdCyvc8gxViMB8
hxstFYzmTdtNfc3gxB7bHQl2fZS38A9epYAT0VSGy/XN+RLuqOuK0M3/OZv2HXr1
LfcWr3j9WwBHJl6jBRyEXsGrLlZVkiIR3VAbv8MYXScRj50JQnu1dW3SXKc624Cg
a6Xgw3ObBn7vTZBpswIP19o/WNYUrHhP/d4j/9lqWMHq4h2Z6xlPC8i2thgLCYjB
LLxRIC2T9WMZNva5ZeEzqattB2Pk8F/CDeE6+AJTZTl1ytmTCeFBZxC1Coa3SWtW
joB5FbefnS1PDsDo0BDEF4HbWp70OMyGYv2l5pCttHcBiCVkhg0amIBO6phCM0DW
nv850qnWSqZVt9QmG0AODjCyWoJOXcBMZLYntIpZBF1W5jbRMlQxqLqfFSMaX99Q
IBng4htm7wA54SVfR+mt/eIyQceaMJCeDpzLIxM6A4ZQqUf86nrae/THYPLr1SZe
8209EaCNThg6Fo/UDCZYqESsikw9Em7KURKwF+c12VauBRTeOcFysk6vYHty/Taw
wKb/AddIOy6iEz/FpaJrVP8snnM2eRWz+CyrpBstYmmEWBOhzAzbbJ9CcBcE6S4d
4PuOrmqeGSBU5lWOAmFOjh1/xFC+7+LlDv6Ca3Lis+/rlAUPkpWZMyNqeBVyMauz
OCfUJhoJECEGthkU9SD1lL3Ajpy5UnldqGS62BmRCVYL5kHzUXtalAZ4ioyptrE8
2poW9c843PWBUJuWn/JWzHIYTp0hEbQqyM02eRqsGzbj1B07eTwR8c/jI6a2n2ok
sF66+ut4Tp0i3aGwQyaVUJXYQHvzxcJf3BefvjPeqRKbmGGBsE5SAx4qv/jEk8Gy
HEQJLHj6gy35/RAOoaI2ZSezB3DZ6PTNd5Q+gq7KiCX3tpfZrGKaDhfSc7pSO3NL
WrNH/wsEtcaJlmxh9EPt6QAH+oTBWjv0+IjtgSdqTzKpEod0OjTiiV13Qwf0D44/
fFYfpMxAMg5qzSUV+ZBaZIoZJoiKlwdOCJOC8pAG8cHjlpUQEZz54zm3VZnbhEAj
9ilwBYmVNiuQKoQSNTJwUVoq0m3YznwfC3s3/hgubnQ6lFA/sqWfEIVM+w2aryw9
HwYIf6tN7PYNvviGy1KHk57lPUw9JF2rKZrNM2MEwwjqEiTa8Uc2Zq6FVPAv5UII
FTnyjYNpQWDHirciU3v1e9yR0NSzmWaGmoPu5N29u/vsZWxw/xiFZCNbdcVJxY6E
HAtLK9uc0129Vr/MdY5FCmh4WacHmvn9kELszkhyhkQZ0apBOuWVSXCACScXfsBX
05MQ3SJ8944QFz4NJIPgmnxK9NFnAAKI110PA9EBOX3p6xfz2BKdcIYgMEzhxXEW
kpei5rh/+sRonHBzx+sGIEYedvibgeciD+7a3KFaDEG4RKLHiN+XhR22ohmTPVrC
5dwUpDtsj3+M6S6NW7dtj4G+JIzd4N/cVQrjDODAkv+jlvaVWvXJR5wa1RV03qPC
71PVToDxS66LAnR1Qzj3JibLdRSf5Cy2bQHXd3f0q7Af1TPhoG3F1rMi04iLxZxP
P2U3zxjRK0lus84B3w2qQK4n/EozkH9yQuPDwQQSdFhsv/r++u1Wg7bBqLg7zHoU
j0+fmYRFgFKhKtHGdE+eVAM+qdiP1eCrQQPPbelqpRHwuA13+BsuqmS4NUpfyGsC
HXTV0HEDbSAglJmVlXmbETT4HnytGEWEJgaT/9zQ8VKjZEzLgelS+X4QVfOzbvL+
zeFqDCk78tar6noAQ7mXRmCMmtq/mOTlUnToQPBJKjaCHB5MJ+YkB08Dvm2GbjuQ
SVzR5FOI2vDBYp5fahG3dtIGXxF+nKYTdKkkGzTQtI/+bF8FeZlrldWAiPYcBDUU
4V7RODBHa/pZFbQct0/o2mNXRJlwgf6q6PBl6Q2NpD5SqS4eYhTnLQ2/OzMIX9E5
KcNYIl7hy9B2vEexVmNr0KVgzD0dc377upynMfLvDIFWRToWi6RnIrKJ9k4RKMyX
Jv9SOMsLXkborC607/dLX3c8zdFQVgKvetrEge0TJr9THkAODzH3gOCHIpnBQ4/h
/CSFdFQtKD2hgUmjwdWEmApapLInuj6tGiHelkeyfTrPCKWpHfI/4BrihS/6rPO6
orPKI4hSOrdAWm5zgzY1R/DR4YvlM490bPnID1ckGe/GZWlx0U/y7W6Hu7e8ymPZ
gNNcLHKAY0d72e1bfcFbdu5ywbyfkDweQ0+/Yc4p1MZ7W0ISVZiga6ysALxHVXaM
btb5Yq4LRTsf3PsUEENaFOq8Ax9/4CY4L8rVrO/8Fp++JOxHnTga0QU/I2ca0TPh
oAZ723saIir5YohAaCBYXWaaZvKBCbBjHWSPAMxOhzaNQdh5f1eCiJ6/V/9B2HYg
fcM61CTO8gHKC8Lsaz4sQlrfS6gqfeZRP0rSFjrQKxLQbGhBCE0Z9CMPcwi1hS1n
myGe4Leary/My1fo4M9KMOe0vX1UOH6O6bbVqmgPuxY6WSkuSk/5mjh0HzdY1qPU
4OvsADDJUHI20X7viDRr5wvX/xWZWhGdt123JEifc8OJtnnmC1murjyXfGt2LI3n
rwDv399XQhatHM7bXzTJeszReUMCzlx5mS8htI59rTk9faDsO4BUtkFFL7VABLJj
7wVccrRKNj6mnmg/+vCylXj7Qfdbz9ER8rvGviwqDp284Tkjc7+iEFjZ8D0T0jBE
ZJ0BLKo8GmRX5uFEquSw3IdJNh2CbAwu9YIdD2wrqfrgcnO8EfcG4Haq/Cxv80mY
gdGG1Ie/llsZwuoGj4qzejOfRFb1AXdhnjzyBrgOAAY/nUgoN4LgHTDJ2iQMdNfs
ZyQMfCofXns5ai2UByFN/LJyJGvfLPPcNXCqYasXYjWesxOoAkRiDHET9VT2FF45
GzxhNAceRQzFtm0asBEf4ej1KuFpHbtUKAI9EVZ5L/s6mPAgwC2DIfhHBSpEWcD5
YhpzVaqoautCTjJ/h0jeyBPqonne8XWkRpXX5P3ql13T4aebIkuCyjOnoWn4fhXc
R9TZyhMxOEni9cHAcOFu8lLzoAGys+dqJ14ODdMjKuHdlFuPMOydKqqtApgXLC66
oWsltc6u0nq2m85OUbVgEC7GkEzDK1O4bXSXFVKEEx94xzV0U/6hMUJ2N/GRmHI7
QwthO8sDSE4fMabUgq23US90u11GPPmM3pwcJpbw7yKK3W7Rp1xPoTRUBDDGJfxI
lmwEE7T9r5Mk51N77XSuwDHOuF5w80AnKuRd/gFouVMnJ9nIfnPKG0Y8kMO5G3Ai
xQGVmWyTXft2DReoq4/l8zZzSLO1if7ydVJ7eo8Ps//V+D+jp00rxd0cUUagCl+w
L0sTiL0Eg7FhAU/LpvJEC/KZehH9tF9uOYhjHgkBXTD/zz8YOZUad8/6C2LKigGH
HBlFeVsxK+Gw0LZQG87ssLOex2tEtr3QpbQ5M12kpegCSuKRVfDECtrFJudrJidF
TKSsHRMyFp9qsX5BJs3kl9IjhEgswOAu1XuLSqG8mRqzDvgL3tQwJr+u5lI/6J+i
RdrzKZZGYjJdMfH+9VSFxLtyTHbi/O1D2aM8lZZWB8Pk9Fqoqs70hYG6n5uYZYmH
0RhVV8t1GvY/r/Fpm1XQDXsjl2DhARozsylJdJ/ugk/UGhaBZABy58lU7YNz0u3+
q3JkVJU7vm1wZXzAp547kMmOk+rPhHw5+9Bq//ak33tX033xz29/pptjBMqsGUgX
KvRIio0NYaUi5ZE1FyePkJtUOnnNlx5QgFoAn1fSl0TALXAQDJIxvHTcReuto3if
Q+V2KkIzYBoORLw6yH+kKjCfCHPL5k358qxVuQ0lOS7DSccYyLHohc6a8bar++7U
G+xB+Thkiu7bTZYEc59R3ZAbjykmZn3ZN8rWc3DWUFiUA5uG+hBwqOEdK/y7gIcN
BDNfiOm+LhCKdy6kumgCiPztv/YkR5R9hy9HWyo4HlRElOyO+051LYIqki0IpltU
LpN1YJRiswoV4a/3GjnMnAdvVRugDq0sZgmsqOa5H7632IOTEIS5+dlu77P2SBKu
LS3jj7A4X8/7KPDRK1VeCPsEGorVeFRrncgsy5sEduF0zOAgBibZcHht9eodFd5C
VLViC74uum2VrRwCYEiZ+BklCEZY6n/SOMu1YyaHEj5RKKo0wS7avV7TCuIfB/4C
7WHG44LcmLNvUOlx0a36TLcObUs5DLX8xp6yYuCbxxxSlkxNIEW+gdv8WHjtfdYo
NyFz495UFhCKN5KxMdjkrcza1BIBcvicQRtxAJaC8c3r2wZ/Z74Nv69I/Cy1zWCq
Sz7IeHQHOmg4b/585Y6KXYrU4HnLQ0/MlFJGT2F1+BrSv8F41wdk5wx/xoAK55iH
MuSYDHpM8arZD7I7c+3lMSq2PUGRG+wABeGPB+fjme1mxmp9J8wqq+eHEKrtZZ7j
J4c/6YQNQwjmDIW2Okpc7AMV7JjkKld/gxMkYG7oVdino+1gLOIhL0QKc7bi3d2p
ouYi+o37kE1mLbwQIQ4vLSmf38GrppvQUdDgBkbZVpHsN2UxXMtIkMTKJy9OCyKe
/7KJS3GX/iz9Oxu3cM1pJGx6Ghol+2TN2RVXtj1eWtebxBwI7hv29GGic8/ogW2B
nlIlgckCc/gbJNi6d2A8JYVr1hqqLGKLEji4/tp2OkVqLUTLWy4DSLREgLcJm7iP
/Q46FdvrrssL4Aegh5PayD3zCDvGBJJodycaL4ZYaRSWxCSa+dCAYO7gCzMd6PJ2
Hz+FrF0uVKk381TW07QLIhb8fvVOf3Sv1+0L+ZR0q1XeBJ0D8A6TtWgPUvtvsDEF
eY3cXaDNUdRAJ4TNNJXN3+SusA1DJ6Hwc18FdZ3ejRhlr8w49Q/nXN88VtLln25X
2/7rU5n+nNCzbt8lwvWIfEIurepfU/Mt27tLTWrHECJX35bflBLvVtLR6cvtPJTP
kq1+ySAjMNaU8cRSPhCArTRWRZKbK4qmxcuSsLE97FZq1q9EabWCF1U8W4dkUc4P
LO+LsT4NpNdHICZc4VR8X6VkEtr05SBht6MLDn5N1mSwAA5FeuZjHAjFts8k0MIZ
mbB+MXn2VfPtvJM5NX8PPWYNLixqLYNjGMCMCzp+hSY+VvuxvYbndgJlvDtx6czi
K99Hmn1eiztg9zdaOEL/LuV1Q9/wp8gKClSLAevexqgvTf1sg+6uQQLLf009G+cP
kpKBg6kfFQhqbrSwDIB8YhuhpqZsYj6cK4pUchGwcanj+mg0JfpdOMZQoV1zQr7z
dPH6+4uzjIdZX9eRKlOyx49RVRJ6F1FI3NnSIszQ4WpUsWXO4/sNNiHSetu0vkrZ
ub3IvQiy0ZpkGOFfxI3YqDJY/CAiZAnVG22WIGNHUN8TpLV3B6M7NeIDgS7f1lu/
sSEEnu3TENo92KyloP2tr1tLCwI+vpRGZPXsetlawH6IKpkDZ1fAD+/b1v/6getc
sDIkb7JKj7vopBN0/z6A3rcjO5bfpRKpjMrV3PjgJjI1OA14lV3PbCicz0S0L+0/
ZzVAhkw3AAgGcjrLcD2e/Qyzogfd6lUzgJzUpK+x2YIBdKt/nYII3EjDGV+vGzvY
gs0oCPgT7GV4L5D2UrVx7beP2wgeElBvDjdtl6PygWBi3FyOzg09ttgwC5jWekOA
9hk/1XRpxc82EDRV1IJcRPvMh/TRG2sAk8GSFmgzou5IIq/MPzd71QZmQKB2ZXX+
96j656fFrYmOTbjUytlgQ26tnguecYymp8EkfRVhDiNXee1RQn0YG0E97T1TlL5g
VlVBy0CjTItpTqA6pz/MzWkhQO9d8u+TqeOH7i/fuC4GJauz48QO5XD1RBEnZnBF
V+T3Yy+Jc7zqzGX3cMrlbx5UQuz9SCKwvqxqn6aKB9BKN0Psj9kGQj9YW1jDMkOr
XYeyJphBLTRecpumhz1wPGPju+i4/kOfbcI0tgvd16l1ETVcSbaLSghUUNg8DsLF
nnzvApO0u4MjVRACFa2DdOFGTaSIM09J2XHr4kLYfmhm81mn8pGzSDB2/RqeYQRH
QKqOaZDgZjfiJHJsyPkvpNb+Ml2O6Bluu3PHCrafdvaaJ71LWztm2bYM+rWtYdZb
mV9BKZNSstz0lzlJgrmR7BU7tvo8TVEUx6MW3/zr8DtAQPo5+c2hyUlFIsQK9xfg
7pdNzO91wmg4UqNqJOE8O573uFicDLAfH0eu81nwOOPhnxnjzlUnBiB1oqBnwEMa
xmhjanD/khVr7p52Rf/oZjQzKgvauGivayM14RmDvutZ9vsWyLgpKpkoWWFTg9tM
nxTFcfJYNlIhQxGytyTfiRxQBIImt2VgILkBG9CR4sQ4VX04+RUKVQ779egQ7IHZ
+rWHGt2MV8GLLPvdaFhVX8rf2c8u5mkat9QNeK3Ri2CwIDQd9E64dn544rTXChLs
h7SHi/el4RFS9g76elQjc79PIit1rA2DwLeDPdPJp1VWsMIQIB0QwjtkydUC3E/s
eas9e2VsdWTqov+6dQOsL5pqLZhjW9PgO6Jx4MuqHKAic4Q9CAQNAeOGDbA3znOj
b33D8sdvyUO9+RA0z27sL4Ar6h5qcBUCg3bzZDn3/aAxrazdDc8s92b+/cpZ5CqE
WO4Gz0DUMAlAF0k5qqn2W6n3bkpqpQ77jYVlOwqDPwa1/C6NEAm9eypJONKRDxG9
Sssw00uut8RDd93GPN6JVVYTabIw+5umOzZL7pPIl4k4g4sbxUCikf/FBPt3R5Qz
ssifAe3Oe0VupaiJrXrGgpnY+Rxif+y1me4M/nxAMEzq3AoZ8pnyHUTDo8jokIQr
YFF2asO21DjiGl1tQzydzxWTCnwFZN+StjQHtZUKw6U1GjbSzpLAr3E5/Pkhq7SK
scMdrp7bDPo6i7DJE5Lg0ZB5UKtttfYqYRVd6xILJIx+j5cuLy4R/D3fmlBsVLqs
9i4R7Oi6bXyAhdiv/A4+QRFctmj7cJAi2EylaHDnRY7ZmDDTuzrTFpk3VaESfh7J
u2n6ryNmYa1b0UN32UWdbokeTfjQC0YpzPxXr/W84NWhYHOo/YRne0VJVGWNou0G
8bDCXG0xSKGB/PwTK/2yVZCtquOxu6VhJfEn4wMgSg+5nzCj1WGaU8Bg0PYFx9GB
7Q0yTq7VMdI5Vs0kJVYdqG7K30Ro9hFFyNJADllXXUKf6gRVgpHcD/wMYRVBrHzn
Q9JPVq48uIKMd1LK+4SVvNvhyCKjl8biAk7IMmTMNnicw/KDLYiOUQPmwIlFh1rI
EJRHiou4NKooWp8HiUNqQ4x/TUGtWz1J/nWC8PCX+9H2DNXcyck43JdGJ6WN8gTi
HgtN8Vm6F93NTun/eavEn/8TtJb8yHEqpk2vTRrxzItvmA7dandXMavHKLlbhtLd
Wt/Z+3o6RNHgO0F9E1/rGZlNz/FNBl5kAs51yggORPB2bn9y7cV/Taw4aawZi/y1
LJfgAJ53+ET70P032wsErv//ytmzyYKS4NbHa/48C8Gjhg7TB03Iv9cWhLe8pPzh
cHnXpb/2E+xkdcfLQe8RBiGKU4Rq1aehyo1HHMCJi9RBQIaI24dy3Aa1G9q7vc4Y
whl90B6/iJ8O6AiYwdaezpVbR1mXwidJA1cgJMa3wsDhEJOQiP+ZfbqlTXzvckja
OWvHVrloziC9JTbrqWGTF4RbQDewmNzb+/Gjjxtm8xwFerMoZnuYTU5T5gQgI6l9
eP7GeRq6G3iANtq2ld55aGb3dDDb8VpnxLfjFGa5pOlOVnVczHCYqzeZmmQ7Lw2c
YctO2jP8MkeDrwjFhVuvgUmFLK1I3Eygz+pXziAE0USKgk2xp5M4wxp6qHgUi2tO
rfhE0tfW3hajOXsipWlsy8NCMgpNkemyx1iQLyq5ADKYfzNqW+K00Iac4ZLKzzBs
OD6+yULks1C5JAL0YH99Oy2jWRyN47OIGAold/SAPrY998S4AKLJ4qYpB7PevB1H
qQYKuMKmuMqUav/K5/FygaVrwKZYygg0CXQ8zmiU2hvB7lpSux+fKY9VUXIprS/2
ljiQPo/dOewI1U8/lHs02iOCI2Q27hKvdslKbmPQgG24jKTCNQLJ3z/Ui1INm7Iv
dj9eSsxwKVwBpo1dENoY9XQo53GrsjXNmCXL/XgmMPgu1mjdy3pLPUHTenS6QIxH
EyYBsTmzSrlhJwE21fkmGos4FW9ESONLsBR90ZzcvCmr3oOu0CW91jCVmpjVdohW
PjEdvCVJrnUkVQgzhKZ2kBNhz/ASP7y9YiGLEk9y/BEGso6Qanqb7NlxU9UY+LTb
skp1+LPzMm6+gKBfcF/55JQJ5tDsqCBUPuYlDc86kh7g3PGmcz+OuoQK9NetT5pJ
RDtFsQStm2v4ekChr4QIz6uqACvZyQrGTBwUBOf3fr7tZcc/fmU+8BFqTwXQv+fh
a5NPpQQWBQx5NihXyvBIvzXShJBPzuNsC4NG4ZSpW7WXbjau7vB9+AediWaYvB+P
dfgPz5w4cnVWF0geQlr5rJR7RMda14grrnGANf0jv2g+TwSL931OEUGG2+NVpXW0
BlLOLuCd2AMDjbA1KIJue6fd1V6s8/e75hf7t8GmEgJKQkUnqmQVvOL2+HgTL2Mb
KeNUV2qxT6jLSe9G+hekjcxzoD7OuAIFf5xosWdl0fGWTXrIj4pabi5QRTRNBcni
aKj4efV9eokVgMan40Ya086g2F9vk454AAR0i+Mz1WAVYDPx54DSB/J/2KYuknMv
80A2Cxgy9DeLdZ3gMpP+2bmcfOQd5h4fZnQPN7CRRxHW5ovKcx/K/EdTZ+TDhBqZ
6aaND8DU8Uro5T4GFGHP/LEZ2dpS6lz0Us0kPqGioFyX2T79vULpf5yeJ/y+9cEN
aK8N6V3KhOc5y3V1Hb6DyDUxv/MkhNSci4Qcn1AORYfs8VpX88M3YMU/nErVmMFA
w+mGOmPYRdDzgIxzYy2fSHsuafE7ygaa5xTGqcLFjq+BnuNbOaSKSwkmtSRJrtda
hB/7VUQqmjNzMdnpR+o2e8ZFIwPs1LDgpuwzIBkRBQLPMH7kSHL27khr2eX80J8Z
VFVEXeHr+vchob+J3N6gcplqCuxqPb6V0u/Y4CWsMOmLdq6dw0E3vyskPhvsBjLL
QSc66E5b7oQpaDtrTlj+3pgaYpef4NfXTvaLIjbxNYU9aJe8A0wUhI5JeSpxLkMf
1GvsGdYF4GATxyODXShKiUNqQiuaxkrMNj0DCRfpeo4AbyLsFv2mUAzrtS8S95GT
dsK8/J4GNa92NMC5/aD/2cjV5/wEM9cSnP2oxbeRNWbxWSq2XgvXyU0uHabxFIR8
X+tuFVAcmuyNZFqFEpJ6fgH47cvaMaRjGv8vkZrPXk4BA8NA0gFP5oNlsoHz2Jnu
LsozHYVGaTmQwGcBiKkn12kO3yXUu0pR/PN7NM+c6VRR3y3Z79acjF5NL/jG0PCn
NnZVc7eUXAt1G3k9j2HDlgIy0oonzzhT2zOkm2syil1GhAzZLmeRtV5gB7vsUD0d
mM5CgzYb4Evn0oFG9wC/4zG4MoM8qjbLEItt7VkoQEamIU9BBQmXQ5+FxPBaKuu3
3daLOLCwsH+YYZoPhS3fneTP/Br/7UJ5zF1SRyQ9uUFxPdEY4jLyiaUREFYdLctU
1bUn8z1iWDdsvvzTBg2lt6yXda3koOVrjC5pr9bE8+RpFoJf6EVEyxlxUP6G4/c0
XY4BwuIEjWpgVUi01wwbfAw+XDu8sn1sgja+GRQPDvSBz8BuVphhsiybx7hXE+7E
ZuFaqLmkS92pTroD7o3RjreSqcIiFV6pAcux4sOF1OTSBnhPvSh293UFPnZmDw4M
/t1VlnfcDPLiafFjGPf/7XwngTBr9uHXKG7G4fEsASSpD2wkYGylP2dW/KC4EAqI
3k8vTvcl3gdEQ1CDbx/q+8BB8gs4IeWH2Yg/IDxba4e1UEkvNSj/gTvFAhdhHUSS
yxEFcUyZfpD4CH7CKefO5dx+uD7Zn5LNin3BaWat8v7Fc5OAgxpE5tukB8GMWv0B
hlCDOg+l7a14q8hqV0mTKiR43FIEEZBpRuXAEeOiLOnsdJOFCSIJqPu2njp1uUOG
Il4Pn6OiIxw/VEDolLtIkLMkGrAxvePuWjLu5aJCKuf9hC0jvqpsft5vPe/YwAaQ
Mqqin/+SCozBJ0JJb5IoQokGpwuIQvXVhlV8pUL4Z5gUiVWeANk1NW6hh+5jQyfU
OjbqZnolWgVtKB1s6ImaFWoK4LBp0D6dOJQhVLV9ZE9+PLdAZQ4lqkZECv3hEUxq
cN2Td9K9+l22ag1DWgbReVr/4eTRCeADUMB1nLrLRAUKd22KR7GpeIryH+yNNkmj
G7sqV2IeQr8xmud4i4fUbVKMfczulNWHRcd3fVmMbunLKBM9NubbDVDf+Ooi4lLC
CntYa+loX56frM0mTAXBjfi1SCjdVE8nsGzPgIn8d52fcjy1UQvPSSVQQ+MbL73K
fyyy1tPjEFIn1Zk508AR1D9NQOsVUwS9PzWXEaVgJY+S4jhuKQJ8FD5ZEpkDEIan
evjCeWW+qsXF7fuK7yUoifHvJFkJemyrxj1RQAmUY5gYIkw+Y0cAubf/HLmSdri0
lmYCJHI80SW/T/QzGrr5Dn274v8CGDBF16taMNfW797u6O32fGJNO3d1TVqMfCF5
BYnhdMyKiDe2HXF7HYh3PO8UnJrYrcCQa8CERQg5OeZZJSF8LrZR4Yi7ZyjPFk5M
hyEfdWxGiKt7S9zsERhVRlOhCoAE//mJR4Fog9lva/iBmualfMrx0hOXqdR+ENoX
RxvZ0GXD8O8WVRkJBuLzVKNsqoFlU5ViC+R3Nc/UIiMjVie0QaZaZJLWDtO3mrSq
YQGIzqlpCCDl+Q1p036fBoPTZ6QHmAavpWCcDLfQnuey4nbqm8EYUPctidHymdSg
p3Ll9Rv5BO1SwkJiq/OzdBvWGJ1XPAk0wgQXxA3kGPa1M9gScnmKpvPSnsjdEy9v
nHyS11QtW7I9am/Nmss7HpxjbAWGPJFyWAMMOsWvtLeBKkL/FuyIpUgGunNSb8tO
3m51l/2L9H7ozZ6RDlTCW3UtTjUOg4+bPG5HsRdEbZXYbQ23VGcptZ0BXPcqByqq
gPCQ2EjyMukezx8uUnTKbh2YnGabutjV17BXVwQoM7ipGdjElFH7s3TTUlq0YyGq
zZQUKKdzMwS6xhBN6DeRkDqZ/iQ36OFIr3r335FBsASCf8a7OgSMAH5qMnr2jnYh
1pMAWPt/jA8JO/mINqZlXReCzKIqwim2AzJ402T+bdqtL2IplqafX/H5oWt6S2el
+1kaE3f1XV3ctsHTVpUBIRExtq95zAvVHl3xqFleZjEyyoT72lDXwD1H12wT07E5
vMFK1CQrYfJA/1QUjsRcRZ9Nz4xAp+OWxdGBdjX/d1Hx2o2KTCP9gAWIA4+2N4nY
+fhjIXIK94/F+7VkD5oHBqANo436g+c+TkNP7v7+P18Y3USHSLGdBtBP02lGe1TU
sFmiCCrkQNm2RxOCQRnlGNH25IEsPzWCZx2zdBtzbj44WHF5O8+mBiBwAMBU0Ug3
4fLgzKehsgeiR3lSaSsYdQnb22fxcQ4ysF2vgl5nCzd6IrFBj5CT9GZWwcqBdlYP
ZcJt8zea+qYKXtjbyiPtaEqG71YPSSufW1JwVCnc3XvJB92sGSewoSRKayy7dw3p
vH95ZShRhNAp3/i9GuWFqDLdomXoRJL3vOA8jhnT9SOayWr0xeHO/+fTq67rf5fe
Y3cgvdY1mw/VnmWbcq/rdG99Z7P3kWtRVVyAw2esWh4I0SCCNStO77KiqXZ7mxBN
OM7v7cAMbPxP1Qv162y7E61+tCQa0QER7IjpkrKZc2xi3KAA1lXhNDPH49TModXy
fRY72dFky95C4h4qlh0CJEHuZb5J/kIWzuTP4z7Pg+rlkFMhSEnqUl9s6Stw9VnL
3lW2XA3xASofTJpfMu8mXmFs76c/+2Jytk6+lu61k5wZZk9cvyyRiAiLwzCF5pVn
bXvMWwXquleWz1sfdqEXJufF5u+cAFGEAK38HaYASFYDvm6ym+GrXTGKzSnsZ0YE
66NUofaemMzzGd3Od0HbFHox4qfuJ2+48WwQ2mmgt4npzfuzOAUQJIdPw7kzWbID
JWNKE0aaYg6rau+1lALhhXFctoF2RgDQ7yLFAE/nCDnr4o5xNGKwbdMXOX9cxwJG
oYIWQiGRrkNyLG4ypjFaEehYBY2HRf8lMmYpE8h5EmbaV2ijo0O8fTjwANuINtD9
9Pk+XlrHUKhcqlf5TfWwtWtNxdZwGDNvmMdBvtBZOBOvjMPYE/QMs+oX2EVkGqcX
D7VCixojAGoI/WDdrHw04b/j5efv1y6V5SFMtoyMvzx17cr+LLlv/3QHhpTPwUXH
PsCG7SEhEJ416yA7AyBK9hc2aLzM7MNq1HpFBQleTj26dW+zG2QrmsvogfLsp5kp
JFnzpgDJbtKHSxDNsVis3C15VFIXFx0ufcHRcJEFJ/7nn7pi0Nq2gzZpTOfVKkpd
79ud59lSze7rR0dx8cAiOt3NAORBdNZ2pjVkF82IvC3fOj6qMFDr0XzFST1qd/SC
3DC0d3pF8X7NIt/hnom5976a5BQby4dTUmBac9iatqoq2e2JtefUPt7FNnuDyrxU
lthrDnecjeksfy9pyg5LGE4mlvyF55tCSmCB96u7TPUSc8MQKcS0QA4D9LpIP+YL
6rpms1IXRxeJrXjadm+u47aPc5wdABsaxEPDqE2ZCuYOllgiiyv9xoKOxe2zinO0
Vw1fXXxFsNg/m+ulZ8ZloqrszfPCxoqiUG4V++Z86bLZSDzbSbmn4ZPy/jxiMesP
pdtHlY2D+fIwczzpm9a6G3FoQ1/bP3b7g9Ml24qPkx9COFBdBgXk6XCLy7C2SwyJ
PBBkvfbstzrSl+wIwrOPUJNb5L3Fy/21eT2YIRpd8eg4yM4LAj+uYKQXzMvIj+nu
JTjOIA9cffpKT08uZPrDSR49LyN7+ZYo1D8qBjlY1S2yugTwV6WySO5uamI44WO+
mBpgbzNOhnuKG71Uko2/qmcHkiwYQSdLNcqsPW6KH4QZlk3MGKyRAmPiAj6f1buM
B8U0yz3NMnsNaWY/ayMSi/eRzYWSqKaJeYDwP/nes0VP0P1oHD1mpRqQnNaHR4Pm
4+Nhliw33i6szEdifAxPPTCxE9rIaqfnPHm+oXvhaIsoTxiNJwtchFmJTC0HZdEG
vacwzW3gu+d6mdUiwmxwQV5deFtj+6HWMGCKNtYkE9Vq/HeCvfwtxMo3O+zof3fa
Ct5A2WyTwPyfWgFIBjsa1GhfzNQFkBnQYUF82YMgqYlOYsW4N4FC8EaXKtPTLIo5
V6Ik32aT1haiMnyu/InWAFtOCNz3+P41owvzme1SuHIMwiaRy6AENupqT1fADu1B
Mtc8TxoWWErxwlBwm5o+XjxeMjuamiA4n4LcMj3ROzEQ78aNx7fjWAS8i9mxK7TT
iCGDS2U53rYkRl+1zaAtUHSEieSMCnYiRKz+WUIppUL0spS4ZFtu+80kXLuApEKS
9XjIAT6q4HL9Y0FL/MCDu8CeIIe5+94bv/i/fHeBmpPnYnzGgO2jnrdqyYPUE/8h
CvXfgniDC5uULsGhryaV7JCIoZCSixkcTrJ0yzR4QJ8EIQYF/IDY+2fFGSBUFvD1
6h/BR3s8kbScvlxCEKJhTBQo2vaJWkhWmayJnSm6U9CLd7B2K6szy0V5QlR3MzKO
wjg29W12x63B1FfwYu0kcGdPd7PRkLc8eOdPCeDuoVvkWucnr3bzuLOGY1vJXWvJ
SanEEj65jhGg6DXS9mIrj7/RupTbjK/oMpIR6kBpafh0V2LFIyPLGr1548BkkEhL
JfX/HwjV7RN4tdvHkxf9aLADFyDHjlRgvDIqWFOXwOWPwCLOuj/UrMrvYlmu2nDK
TS2fIzHDqAnbepHIdSvsf5Rf4mFa7HfndSKgSSJd7yJvCCTsCT+cfoOJrAEyZgin
gTr25McTB1X5iLlESTBGycycu2D3NXQxKceMctXXW1tJYv8zsKbcfCoL5gcOLkd7
MJ9o0+CX8YM/XgJ6Gg0ui21GaI0duVH0EL4MtN+TRCAkd1jkZLT6EuMCVfJPTCUm
NXtIUo/sZurUw4H1p2HfJfBa6RM63LCc+yzLB/PTDhKJSs82x37C5tqHuJ7Pa3d7
7UM26PpHIKQCpSXd5t23Th75aFl/yMAjDGDsL/EAWI0MNKn/NX7gNTngCqA30IaC
FuiEV2p0W/HMez1z4Gxo/ZoPjIloPSkJjqL0RKq0A1nh8Udj/bQRoLbctbu/mD/2
ofyFMKEuzjX8wzcHv8G2nRkP/jt3wn+MhgSBtwWD/5Cdby/lYkI0gQ+jI8MSZwGW
DyEKTQLA1CIwUkuCPXMkzdi1ZJ+1XtTpO1cvrUFztdGUnfZIiw8md3J5xn8zwQBQ
tKjAZOfDMLTCIoep0N1I4ZRZlXpq8d3ZO5H8DmGyCneElRWTbSQK0Vo+sVSQrtnB
l1mUuJaFudfg7VN8ha9bZJsoGXM92LE46tkbpjstytFUUtek7gnsxeFGgh4chasv
Hx0ZgwXhl94mOFyrDXfSQ6JTTxYWTQyPSieOcyP2yT0C+n2KKmDmiG1ceOuLH9di
ymu2V5vVyJOaV2gkMy9oMCbHYv+G0DiX6C+A47gyN2KVP1zSf1ynJyTkVN+gM0AM
U8uvDeAuwgDuxIdJ8opL+cMbSWZ+FppY4uMB7fnFoucbavutrD+rJ8f5Zq4lcXv3
lq+hmLeTudLPoXsSC5fHrFarLwFf5lq5WhdmJfpBgwYQMhR86tDqF+b5AGG1Quiv
onS3f+DFYSEWU+NHyQIHR5dt8sawJK+AJXby64rFYms2/mmy4z8/wAcfp/ZC6uKj
qx7QCV//2HiHbhOgllHGF8XaT3q/HvvJvjugaZhutM5rWR9qVS2r+qhkhfqc3TYo
csyCfyka2/EUC/3NklL+X6wcy4Jwrj6+rmneBPF6r/rPLHTwMlBLywTWYGkexQvP
/KvvOhv07BItaSaukkOzb76ZhcquX9XeoDA6k6tYhRJmfXc9JIzO5Zr5HwA1v3Zn
Lj9h8VHIrZaHoBVdzNykYFdIjro5PJ4zZH8jWm9k4gpEmO7s3vz89tyNR8E3G+9Y
LcZofQVYl4JU6lQPpMO2loUE0Z1DwK/mleCFwY5In9LnClfu1sqK8gJmRZIh7fmF
0WU2VLs8Tl6R8z0EdiDiXHf2C7KXJx0JxTsacbQT/8CD0A9qFyGeE+BWai50nlXc
9gdrPinEhyD3PndJRB/vCfRhs9uUCTEfJKwfuVKyVl8mVcDYkh0KXFY379EW/qs6
RgynxbY8yaIHkJigPrQt0/c4T5RZ1DT4hCy7qNv8MErmjOiG1PirrZ7wbZVJFBup
bqGMCN3U/4ZcO/g3X4151Y/LQdXbOBm6elDz2KjkJxifIEIkbPB89uShB5Qmnbu9
1lGMv3peamFGuKQWLlSEhuHaA5adV5zk6554Rg9Aq2XFPd1FfwkW++jMlMq6hkUN
SgheTwoSsF/Fi7XDaySd4L95YQjnw4Yk+Uj9wcx1kfpO715LQQ255V+rDFTt/8aJ
d2xdFNxoBYAA3U8b7POF5PuX/ZKHypWX0LbUdn+f8iNvY2DUU0ortFnAJZxx5BAD
ctbtnbzrzYCmpBzlhaRm8S03jyrzJAwEX/vQjptu09p3jXVWPRQzlBvec3C+mq5V
9pNLYz6fFT3cI7cNwFeAp4khWx62PPrt9R6SJqwPfqcMEBtMgyLiVorV0sruSNra
mDJh8MoVBw9KoQYLcPktFL7EnAB471GHxaXmkREKTtzL/Gkd18mj9QdzQQeRHmVU
70bJz3/pky0CQtr/eFepslvAwSq9WwmDL59his9kzTA8Flz4/zdUohP38EFNbxv0
BRn6MKiVbMpX/8oE16jso087skLSo7sst+S2ryhlXoAF9pR6RuWMkwOEeA13xlrP
2hu02bRQ3jOcVqPyl/BplkFiUkz7alKvK/k0x+NtRJQx8qahEGz0IWqYNMNBSsjj
I71WGRXNPn5ZNEgoZrvE61ak9tVskC+yN9bzRUFySqrr/P6cGj5s+f2l0c+dROQW
fktyavDfRZs2mrdhIFnlLqlrfyPJzU66pBYGsNuzPA+L/NaGU/SZfY7IiCw6CNWm
8r3QjRhXO/2TVLo6UOl3E9RZSJ6+BtpUfGqo9JdVAHtaMd91zbRwvsOpgPAr/rle
xLyjfLDx/VoPavSKjYFbSGyazVFL1EmAxwd5C6gNT0SG4s/+KU1zhKO9NiZ7dHhL
gS0ch9i79TFl9HxDLHAP8GUqUCuJ5xBS2GzoM/0SDdYnxEQsQUs1G5KGGHANhcG4
5mLsNOvFgIrAmOvSzyLjb+DDQ4QaXa4itE0bf1SjEjnFna1hXkf4TcLKzo/+wj53
TtBf9jo68dSycWwQCVZZpDeaYA6P+akF7pQGb9AddtWjcatYEpwJgX+d4sxDdcLM
OJsKjzP/XuloRY5JXwKx66MfDW/v1n5lsdLPO1tACJgZzNtjZJrWZVOccyqjO+7I
Xyirm28TnSSEVvEkCkne7O7VykIvs33W93fxaQhYg5QmURGkicF9OBkJw+s5f3D3
uN0M67ALFDiY7emoWW+JxpOfXexyc8Ls/AtrEUaYJve4Yn7cbxzviOuiJOMWVn1R
VmU7lNHw1VHzB4QilciWmyJzQVgmHDaosDlHBcVwpDvGZp19qwJuCYNtK+T0RNzr
oJc4FkIRc14rn68QNKZAXSganmPmS5fO5HRFMv5d6xlHkfQdB78jrwxQ4/LDikGA
qBzVSoABurQSdx55lW4HrIsTMuTkwDsPgPanv2HORq1DXnVPfoiOx1Db8VtjHKrb
WMrfFgtFywXKprwNjNmkQy/gCNndHgTgALpFv/S3AMtON41nO9ljjy0bhTsz4SGC
hqAXnACTewJiqOsUeoC1re1aVJ72/B268jpo0D1h0j5hgJRHcWlRLAlAncBrmrhd
omqj/hSSi5ASnTdBgpJoirvM1e8NZIe7SdJTIyB+2Nkd/lPpRBRxXsB6+c4qLAOH
zuLYEoG6zbF1czIhOm9vH5yx/ScJot3VUrIqPqw6dN8ne5+x7jPkVCdqIsZzQxAA
CT+9R1zpZlbdOrtRuUYFc6IIidzukXzkuW+oR7PpS2WNso3uNNnTpZi1La60HcS4
q4z2qvevVneC6dZUIk4SidwVv7Ksh6RRsQM6lPKlqyocq9lvSoQj5r3ATJppGER/
d/Tqhv9xhaTCX3KZNQ2uT6opa6ksrTr+1dkjznq2ubnN5j9OOdf9C/v5B0ouv3PR
VZcIIYO8x0wW/T/Kfus8a6mFXUnHL2Dse1cnvnytjl7ecmZnmKjL4tTNGKqGzCkq
koUJWh7jfZcJecoCnsSw+/cxE3Kfm13BTYGG9DNp/WGby4fP765HWHeaC7n1tGGe
ZB1jE46LyzVUOFUC1uWsXmcwuLyU3zurkQku8Wks2Hn5CpTnU0yb+4BfXh8GuRvs
Z1Tnbp+8ii807NCc+6VaYEJYlLqWe8ktClciomhDWi8BQRDtaBoNjq9Y1nUfkosO
3+xIZZDAIzMvwX2wH6ljIasbSB+IY//DuCwi/JB/EfxyCIE002/cAFuut3Az01w0
jdRCwdchVWLy/zyHO5ige3MH1UrmMRkB4ymRyQa8HdRdhfkPqODaW/up/kcjGoCU
AMVLKdBO8LksmwsWXT2hw2EbzmQx6zdpHypoGd+ecclGem64qnVM1uDqB7CEDrJC
W65vMwOD2SEhup1ALAu39/f1ZV2FCJJbG+OwQAhaLk2xk2Jo0zHGCRJqiwsWW7jS
eu7Dj2JwLSBuae6L0yfH6N/jRr3xny2e/iLTul4tqRwrj6YSgttUgv+v3v7iZDQj
qKX3JXbgTGFSQitPL3G9DN4PCy/3ZooH7R1TA/kF5bkSnbG8ZdYsOPB15G1iqo2o
Xi051d2SHL9G8nVcwYe++6f91PTymkgNOM1qa2bE2NylJ+mjOOowYhzgJtkHPY57
kxQuO5+Q9HiytOtVvK2Xmpzo4ynOaKyGMVVPw0x7p/S0S1vhh03qy5Qf+X/5+9ha
brBx32+9Rlr4QDhc3y8A0YM/FF1h9sFV5LABF8bx20O3TFt/pIYYE7LignrXL0yq
+0/RA5cvdkIMnvPxcavMGY5z5K5MJW8hQI0bpH5a5+AkSOKGXxQRWhCY7mp561Cm
j3GxAN9WYy9+LTOrO27W4351reNVOm4bDZx0R2zI/tJ4hJwNvuUN2OrBQzwnCai8
CiuuvWUdzIDggsp4TBLsepM4cTLtmoPA4qpNhCD8URZUXUzQ+79ph85xCVvjMrqI
KmneAl6tGXSAHxL7A+VgzRd8D9RFdCcHnrDZdsRBMY5Q1K4860e8eK9ne+2Nxlv9
Zd7Pi1DG8bCPSQCp3XXq6F4UqKlmG56nWz/i9DvwkAEraIkmlgxNO0D2aApea9rL
aDBaFDn7y29Itmmkg1ON1uxLUW6dqAyxNWVBsYZ+W3ATXDnmfM1gnWFgzZpusQaU
Lsym0ccL6y2zNE1HRDzZynPdyT/LU0e3CxMM/kM8iobNxiLsio2FjkRJArqHM61B
7D70f4rZQVHq22ZJz3A3wzPjDZ227F2NAQZjXrZhU2/stut2qBvd0ZrOCQqMAE+c
gDB37EK3w19K3X7mV40nMkvqSKM46K1CUvZTLzvMuSi/3tL0xdz8aBo9wTY4jwaq
v4cAWSBYR6b75GK+9Etc/UbF930zklQ/O6IM13GKIKQN3JiAH3omL3Ucei5c4V93
pc/j9/N1feuQY3R2E0cM9CKG9KZV3k1Y5H6W+4L2BA42kcU252IT6+mtk0rMQ2NY
bofVj+KOA5QxTVAxrN9fxh+L48mdbe8YkYDgfqCTwt1JJ/MFI7UsQnOl0x4RFaTd
gNHKkCCYYefG2N2hD+ICjMQ7xggGyZC49Bto0B6LtTJhwEuP79Z39TlXnRKrVvIJ
InWC/2udS85dg7q/Rz/cGM1OrVT56GdUsrG0iIKjELGa2oAvw9M0qvY6K9BmAz20
dWon0+zwAeGhUg6MLpqzTAc6vFMN0sBlDKQlibByg75P3vBJPfA18rF9c2o9b0Gj
i0QCWI7PIMHwFjCaZ/vvIJsXnh8Nt+TEtIBtoxcqpAnclotLznelXlx/xURCXRT9
DYbI7J3EyNeEFD61oyAKdvfWO7SAYe4i+TdAGPna/qElo/YPN0TKIFR6D/1ofS3f
zcnqIX10JOJxAZgRTFLp/TYk9v/ij0ccVMkN1oEJ1jzGsERKTBd3nZvZzFVJ6mlG
zwmwGVkJGD/Cujf1CiWbJo0Lu7L9OUGCOt5Vx1X0qMKSRQ5jiL44vGugZRk3OP2O
OUdnfJ/RAPSoc2CfMSVhCJJf6oV/XuA1sip9ZcyyfNbMYEDqU6K6XWyUSTpT4Tij
vX7YHoxVcfEwvE4UlSvKyNRWcWPHkgWQc/T9J2uiqQEJ3hkmmOi0bMqivm06+ShF
SdZtY/t/KyYkSnoW21JruUt0weLZvI2ptChjVr6fmOlkqADP9kJO37vp/rqxGV1W
JTqhaY97BluSZWeLTB9+ll5yTBhRn2i1nOv3bChzGGnMwmmpw41TfWPhOkujWLVZ
dp8WMQbrUT6/kZRUtwHY4nVxTDOL87UdiJnLPB/ArYZJBlmRL7pIKY/1RxLSL1le
wyi0HtqhB9e1VOjVVVMAVC9z0VqaFG1KYAEddWCrRhmRTzjm0caRRF+GxHCYFNGK
8sFhu0u5Np/qS+Fcz2dRJYgR/pLbn31MY52oqfXdJKJCnv4Hi9rsXriE4WxDZvDC
YbNzdqIi5UpTDcNYwP3CzopzcU3EpdphbuIUnx1zZS4LzKSjin9u+rgjPIv+jgDt
mLbUoqUjm1J7DsUlE3hSBLs+6NBYG3Ons01zn1js0wvIQuPkx0GYdBCV/W1mkYqM
yO4UtbYQMzteLWSueDJSi2fhAcOmgWgd6yNa9G01W8DL8AQ8nmaYa5VelYwgBUks
aQiQlfzscs0u8TdFmAjBTaiQHJFwFIHBGt95b3i8P09gvyP/iX/qj2f+dfuRtqPX
hAcYhrn5F+wboqP65jReslOAWkegPuzViycDuF5YN3bjCDGBcIiEKD652lf+pG9c
MPNxNzoiDFccMvVtVnciwzU0sAGHakhPsq9IJBNy+/ZhB0dKvz5h5QvPGnrknRVM
ighB4yfobDa1ZIyAkmJ3fjkX6tbyzcaD6NE+2EvuBBUF9Y6HIGnDJCQ+4nJH1K18
P3aaOYbP/2BHsKrHs8IFIsEpayQDj32WmxlqgNL8bmaNjRam1BgK6mNETlfuPlZf
kua/HTMxKWmqRsyM8HOLImtzu/EbsVb13my5B2XmCVtlZ8NISniGso2IgMGUqx3Q
85UdBFPDQDx55f+AhL6iGXgaLPFHmBX5K4B8b+d3FGGm+zHQRZ9JT4qFbj8z9VSS
RIeFKNKv6YJ5eQBR2KHRkmiP03NQkD7W22ZZxQzdEINjbRX/SOc2Ilfjg//KfkcE
XNwRTWY+tFKjWgwaadZVyvCVTqBCvWRuG8+zYPlxcdVdFLjZteQgqlktOcT0/7rX
INTmzhy6wSIASCKBo+bRtcPAcEn7cc3G8tG4OElbMj5U6yPBg02CxVGAp7npYAGv
QtTlwY07cvwMJFAVEasf0F58aozsdE6OEaHV7Rg9/zqBV/7vZRBKc1otrcNlIL7K
DZGnSjYVX849tSo51T0vBVlyNy8ib1U8vZNl7VDWXwfG0WOAQpq6RPziQYGv8WNU
n9ApN1iqPCWgLPM4zr1EpXPvMZMeEcK9rVHXhZRYgApvG7zFk4x7D9mX0a5YM5LI
fk5eOYAqNJ7XIbHEEE0ffyTpdohhzjhQoIiG9s17YxBQR0vOrxP8dFW1y3I3+VpZ
OS5w/h3y67BNg3Am24BaSZAZooruBmY9ic1p4MUIi9Fo5rN9+YDqnwtFFA4Z09LC
1boQYRZqXN+b+f4mMgjUatwM8TSbEuxRv0hEvkt6/nWOcwks07BB6uATgaWHzcIh
nn66rO+79BMiGeLwDOb2RMpvkn+MOITFQ4Q6wglUoRhgw+fDJJ20N8O1/2OUQctg
NtihjcAgsjbSUZcHA5EoY71uypcvygIbUiblPrbYtJTFn1P72WlkfeTrT651mXRj
f4TdzAiWP7n5oPxvvk/OMUGLN1RlhxXF6jBKUHO88xbUDnk9zRYMAtU0g389zC8i
Vhc5vaF8pXVWMLp7P6TIAcmuYhCNP57m4CS1br2YC4aNXkxvtDDCPZ9aJ2leQPBH
KJPwgJZl9MnDjZ87Wtc19Qi5lGqPx3fbMIinQe0BqIUP/hnFIGA62dPuzDTwAZl6
OMr6UsVhbVxjEiWBPRHc1wVCMJz4Gh18m2s++pl1fvHE8DNiRbRS7RtmxJmR/vn+
uR6/rjA954CA/AZzfC3WC9XXgiNyZX+CIB3iSJmulg5C1ryrxWBw6hlMo9+545pJ
JVB0+3WDXxeA6CqTJcVJpG6/X8qfM3b7K78hBeawdmeg3IF57C76F9zpGClhXpR4
JQfbMd6IVNN4/emAOeg4s+b2F7srbl5Gc/+Wi7oYLpai8b7BohAlR+LMBTfz7skq
wms1msKSujprtcOrN3kTLvSFTF2sOrvi8xdcBUZ2pZVRNCD2wsatW7CN8YWHR9TF
3PhLIJ52RyGKxh7qYgqDcx5LiK/SiaQbTbVdaoX1dYXFcSrFXJPaKTg/E5iQPybu
OxGYfm5+tIPcXek0gF2uKKqyjvDmru5ESu+uuKdS6IM8XNgP6oc1/XADaXYeEYKC
WjKWiVDIc5csjeBwJnTwFuQLPEZ4RZyGVNXQuPJJjp684W9oLLboIEMBHVG+a9he
Ft0Bw8eR3Ka4An30QYxl2YcS0ELUSlS+kH1qv6LtlZejkF2W6szic4MKjG9TuetD
RMAG1KZiktoTgSAyxGHH+fFffLDPC/vVdMS3gb6htCSqQc2gcZO6xpmGmR/RGfjj
Paq+1Qy73BForuEYfyNLDI6Cuj3KZ5Ey/KeyHHp6RSd7/wrzFLvmcx9CgD8GB0H/
l0K48tyGi/ekjc61hvVnPZykbqmkIDGOOtU5iqGtq1rE5GnM8BvUMw/aUOI1juyj
FWopLT+DPw/1Y+YbVKIQKxQt2hRCNDaRsEcxeTiPQt8Vb0UXrzkXOwUdLCmeBerb
s1eZqhjmesvGym+xtDWKlPAXT2ROFiNVuo+wbUnc62Z2afp2KxxIloV3JoMFgaC9
IcO3yREYi8e3F77gvSOXnX68DvGC6h4Gm9nR2SqFQrcdAKdI47HWdJaGbD8uNOdG
I1yswtApGi4DZEGKgL/t+kxTZwWREXVL93y9uQQz8pJx6phIhRFMlNOcNfbuKJf1
lYksyYZVHFivg/0AAUBlzgA5awFdNIIdrTxW0bWfSTiLDJX5BFpgAuErELzraybI
bmQ6UTZ1zcE/XlHq6OrhKPl87RLc5yhGoTGANyVjvPsxHer0n5fFx387UBm1VIMZ
1M0zv/fnq89mL35cqJ4xneIp/JUiPHG9cJRkviN1fa07nIbYl3PlEe3DvHful7/1
vcR7Wo4hcXYLMFA+jBghsTAT8DOq/Doaf19QdEFJm6C34NcOt9pluOIvonBsn++E
7TqTe/xp+Ah/irbvGj8OjKyWpNGdIMkpMIk8gRHPWNd41Tpw0tyxAFOqS6EUOeXQ
i8zQ6heEdvTlNGeXp/OzB/ayD3JJakQcrK884AcCUedbsu2sKmqvyt+1AT6URBZL
gtz6rSMXbl6HfAEJxOSpeXQXnkOeB5pDvSxl4dBwHEe1Qqt6V98Fxx5Ml40Zkmd6
D0NcQwRd/eM8MG+Gd3fwct1p8CAKvMjgHSejqfoCLtPs3TCFrCUoyGmtUtG/ZQdz
Q7VQLZEknTutsg6koSjdY08vcUZtOGjE07shBK3NXZRny6yKuJ581z3wdqN6ZzBm
bCDDPurPN2HExj7UYLJeqHUAgP/jP8JumutQDAjJPt8bkjfaXcgpPBBu5lg0xbEb
/0c/QlNYK9ls2iH/FMz+VEcmgp5Blv+ZZGzq4Ymte58DqS9nvrMWr4LJivYGwwY7
Vl+y8vq6Zz+aoCQxgHzafi29domcm9yqE8u7S50rtZvbsVvh+2zYFCGtXQJGf3qt
hNH2HZWl9A95oGuiJQ9QPbBz0zSQ+zKpn8zlvK+CdVGUSsY/yejv+P64Mxk6YCXn
mBtFgpSgOTu2jvNCS3VnNN518DTLdaPCbuBEZgn8cKvcfTwKcG/ljR+RycaQb5SB
vK6gzu8XJB+uyrb64amutPvmCxu40XWWXtlfgDmzFTejt4xRW+ZjbmZAgMuxs4Cm
RKul1gsKereXgQzhCvH8lSgMAVfFqFjaBwQ8a30lt0TIu8dGvexIyXeXX2lc/TGp
q0q45MgAzeVXi77Ez8WWbeIDzgkginY+tfuMVKKvMLtOr8CMNLliqMQABAqR+/Qo
F//5278oF1pz8BdPtEOZcNm/XHPqC+dgwgCzK3z3EHXyBtpWFRWyZl9Ri61rG6po
Ip3j7I7PmZmnKzJ7t5fp421VHL8EVHyPCs00aGxE9BmpWy11pv1E3qaoT5pCzHR2
9fbTtv9vY7x9daVQOyv4J8j3U7aviWFr4+0QuM/hGPK7HhX5OyrOApNUrDBQ2MPg
8rLa/SDLnqAc/rpW03IQi1E/uwwp0VbUygNHrVqPntzthxF2aftBiG+wZfSy3MfD
f4xVa8689lO9Ebw+EaH5BZp35ZfeunZLCFa985VRI1uZd0NLxc69l3t0YcnoCetO
bd/L8QB2W41831MYai49BgskuqEqAiY6rV8SDd++JnVpQq1l9CzvrKV/IA/BqbAs
fMoKM8SdoiHkuLnc2m+YkwEeBoUisT+DZ7xl8hIzpNl2HVQ3lW7GASzrOXffMn1K
IMyI6STgqcgmImIGo+rE0xczJ2GiZ9saUerBbv1SAomHEl3h504zOJztQJM1i/Jm
5ESz7X4gOlsl1A5ogfSChFPELZwZs+VF3VB/XlIeQucH+akC+Lcc6r6IR3uGBlZ0
E/MfcLrkq8aCE1I/J1IXxROAkNlUOAfCeUE7E4J+n1gIgAJSCxQrqzvy+wiTV4O1
rIxdrcTdKbIaEkPwcCqLYrdiy+17bkaktpjyOpKjnqcWabGWRW+pUUS6KJMQname
83Q9pIzSWmjDENCkVr+OQkDtmj92z7uGiA4Qau6EgCZNrTQacG8QXl2kQEFK6tuH
Bn76JYuCUjZKrdAcDgmGagY3ty91uKDindhmicSQyZjXPOO9S1x4/eRk/jL4E05F
vGtaztZivTHKr6Mr2KPLw2kX+5gGqRyFGqSedMJ1qYkD8X6kn4nI4gEmv1lVHpcF
mslnmX2vLQnlaKlg9s2Ch0C+VAvrW9bD+dO5mp1aJPM9wqX5twHSGSOQvTuAKxNU
+cuSYhfB4ZFKSiRrGk1DD6Xghtf3OdX3kJBAuDv3xwGqxeHZOlO7KPhAU/Ot3PBj
OlZ2W7N8ZpINBSRqFbhRkV8KmZQcoG1LtX+AzgVqjjK/4Y20VJSPyz8x64pMAG4R
FFn3S0G1PKWNX/LQHgqePLNBEua2VjK/swu9Nv0sPUIW9/mqTbj9hvuPUazR0Qrr
eoZnm2fLi0znEFgB4sMaO5QvDavMHINZHn5Hq/Nw+dhl8M4xnNR8rM5Y89xSO77+
6MrNblL1y+TKZwSo2Dj+8Y16Qs+t87TwuveJDYJ+jOsjzTzvQ4Q2DYfh0zRZg6kI
NfatOPNRW70MAPLvCNiMrqyyQGR2ExnCXumjj+yv9CAVhZADb1y6GLml2SAI5OCd
N64AfiVzZYNRyf0VVu9nPtj8yYTCu4suacScqSRlpWVBoCU/UZqL+rR5vuERlvTb
yR+Vwaz6Xi6G026W6ys+IPx+OCxR4B+U90FVRWjhUE4ZglAagUtAUMluZ7tsMWAF
acgVAPuYmKSB4g9yKsS3m3jJ+YbQVtIycCR/vb+7mZ8D81Pkj28QBvb1EGmKDM0W
Lhlx88qh2HR6bviHw2bFygZHCq28qVGwijiepQ6bf2Z/veZHjn/Xnl/Pdx0U9uMT
ZYugCTVriM7QwEnurvoYfI2rnC6FkHJj8HLez1DQOYoGyka4Z5ckI1OlaPsf3exI
e+OigZO7Y/iGwu4edJYsSj7n34xoGwAaitiPoaPVLxOlnJYUuYgS59+6vPsQgsee
yUjGt0DkaJONAsEPms8WKHNAzTf/1IoYyPcUiO1XnefLCi+4B7lGIhl7BCa4VaLb
fBlUiwmUcZW4uj9Kpm7m5QQ90sy3aLX+Q5h95PfUNSfiyKBM4CD8Ab/pjr4gP7js
mVPh5x+oinu9QrbvWfsdLT8vfyqiwOt1LN3u1zOqIzch/ihApzcqbLOVBxqxp0hV
GeUsNwDqclzktsU62WH5aEDJkqqqFGdO4aDqan7mKoi5v0cAJ5na17XLB4Xvq1F+
Z3YW3nY5cVmig10R+/PV6cSK0NmT/FTuFs7WEmwjiohDK24gutauNv8v4OcmQF7K
/GiOioItCtXTkEdJY6krVPR8uYLYi+rjnMGePKXR2AxiXZoUgLupVhpazmjtsYSd
mwigXpppC3tv87LET0uTQE1dqYQJE3rgH80zYHBj4EPDgFNSzyACAjrb1s89SyH7
05eHo5R8ff7Yq3HT8hUz/usJVAjVoGeG90VZx17pOpORn2XYK3HAfrgKFm/ovnJS
R6AHS4Wvg0gxhdu1jvcVz9+4g7N+zwa0Lf4gENMvQrjrmqsjJW5Kq8knJ6mxyran
uDgxDwTnrd3QyJvS27yb2qQ5XO0RrawTb2MCpesror3A2MzENv36cDMevAc0j+l6
6szRWDrTz4F0xuqWULu7v1UMI1Lntr2F/Vd+FV738vFLPoigONAAeH1EpefwryZG
2DlDHzlJryigCcwgyQ5wmadnkMoG5z8S/Mza/9rWvi3knm9+juqftMh6doQgSVvL
3jAEwtK6QW3nrWCO2nJZFSnTLjRjQSYm0coa1i6nHXhlLK4nosJ9QwYByo5lOlQc
OMU+QxItq6t3Np+3arF0UAOsZbuF0P+NNVWX/WrsSEa9uJXL5H+V+g9zkr8jB2Ed
sHCAwGbRTi00ikOnIHQSZdNUGEBfsejHxiLyUaxh1jShQU3KvEBqoEa9XAYxWHG1
9voVqQpOwLqIzvWi5T7FdqrlyKcBy0HvcbAxwNMHX0k5S7LLLDIcHXsWDmK0sICB
ABZKvA/ore34htZJd6JZ01HwBlP5mJbTaKb7sAoFFRlKKyiqt2eGnwz66jMF1sYK
0IGnyIn1nNWJ1SWl78cRaWA8d/Jg+XH4WUREPWmgIccQqAUIpTv8UOezqdhrYgJv
WC/P+jD5KXu15M/CHeAIDYRSav3Qt9EYyM4bI8HIReILayS10GtdJ8nUOGBJ+qFw
/bPysj/m/3mDCVLG1kcNjMAf5X9jZqy6d9ErxYZydmKmQe7ZZM+odBX26pIH9ECs
I68fwqKr/AFp5ovN35WgTQwWuI0DgBi2CbHjhC5gFua5J2AZqNtU9gSi/vQNTJio
GE1dfKmGWV2Mp39GsV5tvPeG2RnV8ty/LawRLj6lk9YJr3GCPB8oD3v2k37uvj0K
bta9hlCRhZzWpSVQi9GOkPvvxdbnqiG8vY8QM3HpdUxV/pZApgLP+VuPsQZoIQZz
gfsq20SG+eluZ/hHv3gZoy9Z7kk8d8eA1lIuTnxBc5HwNLSFAz6op2jTHi+QuRW+
D7CIgIoklUHN5ze9E1/juBfFU4PXXbo+hMm8U4G58xI+elX2rAQLyiSnzqm2QHYm
lvG1/felDZ9wY6c9o5wXOUnxZnjJy1v7j7i+tt8/BSHBhWj+HRnUva4K/ZkVOSHx
PoC+DGNF5YN56d3Fvc8oKiDab0HsJniZjBKixdlti1M62SGoYphCOg/jAGr69c4d
GE+LuvYoGJzL0UgQ6UftTjLHbSspLDZqXTl+qzuPPr8GPaEbLCf4+u2ZHnd8hs49
wmpvMGbSfp8WjsgmJom60Con6HwuOP2PL02msdQknkfy6MBQXGNaQBYe4XdN/FtD
pC94qCf5VSAJiRom5SLKFLtaw4qv/0t4aRl+q15r7J9kAdmL6Q6OhRxbo4jEXkxk
qVmM130trmWcjn9hZogMKQdSupWqwJJ0fSmilXz0ZFquLzhfdKkq5Wy3NikUmzuV
dzaZHgGGlqzDmqgkG4boCmJYDbsPGlAmeKSaWgtqa+aoMywFAnD9A+snhJw3FaDP
IwurnHp/A2GHoV+06reIsuwnjIBuqJwyNpfQ1Lzh5ONYqMXlO8LXEPToXAl6PcuF
EchNg8E+JP/omwA+zePInJKaI4xOX9yrs/5QHOJHyQ5QVgo7asbA7UB21nWolooc
lFM3I/1edhXnAVg5S+hnGPUHhEWWLi9gMalfVO6pPKzvDOSSvDfu7Gw2OmADPe5v
gWVT8xu/6HXHd9OkZqb+5AAzP+Bd+muoPM5HLIz88CDHfuiXu1A+3dcoCymvs+GP
nu2m2CGAovVt38RpTHaRbtnLEszytBES6z1XQJT0/ARTCZMUP6hlK4zUqvrkgTo8
KRBH2h17R+5avxq8Ag+mGNGmrMaHDQpxSUun9GFn/Kotc29xejUITclsG6LUC+gn
CxplHnvTJVbEizdSj774cgEZ8FWmqhYZCtVR2Lti62Isx+y5nx2uOjg2bHLquWCY
ZzhPW+FajgCNonZ3M0RIRcAmsxBGvC0byDL8a8UhGl4Un93wWE8A8zLUuNzfDMcl
R0PIlmZ4GApyihDUQSmEktNLZ19oUFmdk7YUrXmpvF98RTiClybf9VC4iLGbsKys
+Po54hBd8IbXrX5DoBr3poUUaRtKKs2O4AwCWONq6mkY3sVQbHOBrMmjl4XFrrNr
+yExftVa2S/Ze5mjQy1upWhpi++xdeJzOBTe3EiMj+7XIP2SsfEc2c8aF7XmC616
UvnaoWzdCxrbx38RBOsQVFCz21JLZj0uwT9p8CIOmTKuVWF00UMQHsMZ3aA6WdAy
A6QG4TxmKQpYVGGX3d+IVUVCgFVU1Jc7CYYrExxfSi/P04QD9lYSGOssL0n72gBd
6GWvmjrUpp3BR4DsCgK5+U41l92FDyhuUMRZZf3pAbMjTeo98HwmWPD8uqTIthKC
HB+Me+ZdIEcTFGTXKDvwFg34Z93WB7EtlOSCZGo7g1J1DmK/QWMOoDU3BO5hbq1i
PKwYB1HDhcJFGCGSV72lkLYD5LDxeNerNeersuoYcPnb/vn2RwWHAa3ss+cJTc5y
j6Y3PuCoCfPc2Ewb5bsbaNjJYuI/eCyCHRorstPxmim09ZrPe2B8EaIslE+ohBxR
1MC51O985rkBcKTSm6ku2p9UmI1dqeIXudP2CrChZOXLsOzxWxJjd1X9mkDsjdXK
258THuaR5v9snzcwSmmhsTRVrLn7KOtMD4ICfFMBkNDCvByv2SOVrR3OQAgeKTP0
cfol5hP9w5T8EJbbjr6f/u2AObqp9P//u6DmkZdgWVhki49LLc/wz6dzQ5ZD0cc9
uK+Z5bVjGUUViLPc/4nIY+xjzSVD+cIfzbhF0zSklKuhv9NsHCG63Q+l7OyyvzIH
L8perVIZ/RI97KthcvZrR1vb3I1LtpySm3PO0D47PbcwDOAyjnlYGGgsx7TCsXxk
Yoji29XWb2jXAr7M3v8plc/QsH+fMAjHqeoj5Svhp3mxqkYv2HqGaDN2PotJbEg0
Y+q7wEGFNCM+4/eYnFNE4o5UbZs16+SE4SIYPO9UN7YuVUyasm/1cFnDikls/iQj
pznK9vcfoj8BbdfIqcV2hDMojBP3FnbOa+dDBMCRqc2uNEMW7KnG3o+3nPklPork
ezwCuFAL/nHB5fuFMQUOQXKbiWl5FQN7acjEwUHtNoF+cUI0/o1z/JapZFHVEwuG
gPwroeTuSoAyTZZfHx6YxkCWWYV8+K2yClsok+VOM49lNO4mchxkRUU/+U0E+Nth
B5E26OXWEAsg9azHrAhzjBIT8L5kCCKIug+w6yPch4jpuEwVZ9SRAiAIj6qHJPhJ
BclUFMD/kQWfDUDPxDXJtSClHw6QyP+Nq4UT0l9+HNraIkOIMiyKlXfz/g+ujR+W
j1M0WJJoQywXzGSZ5i3spmNAgD3X6JGh+gMFr1LyqqVcj+3dl3AxsptBnRnt8EcG
hmhI32kz0I8lKwuIJPP9CuH4Hw810rvegOOAARgU/2PQJOId4yPUD98EfsWF3JId
fsnvC7ZSZ1hMAmzzOTrZgp1Z7ezwwOZM8+XZMLzfQklboqxMvBUf6sqB8NrIaCaa
sRPhN/n1bZ+UiohXZunzAWig/sZ6hgW4v1mID9mKW2z5GRC5ADHSUKB1fXCMwpe0
Q5ImjiBfb58UDaTZuEZ1q3WfGhOd+6jOwFhdPGERKgvwMSn9RtVAQqMNk0baPfrN
lU7dh5apNqH7UoRueltID4lhsh5TFaqCaCD4E+gS2AKSFck+kR+0p0MzRaNa3tXN
hY1tPIoXcBDT5qaakDwvbC9jEIM/Zkdd2sDuk1RmApgsR0NgnDAhfZEDkfGuVa++
Zv7QUr9eQ7cA1aKGYdO+NU0uzJslFnDnvWR6rNtcG4rjVZLuGMiVSo7mOPaBQ6JA
jyvGQsTlex1BQU/bMow/n3Dg2rY8vrzv9cbYxaPmfcppXe6teYciCk8wg34TehCm
LBlo7fj+JiRy9LGM2X+OLf/7MBtOEmuePALKregjpAfPB50wv+3ay3GHx327Uf9V
AeqDGBgMGFJucVT0foKTT9RW40RwwIwGIfA2GRaL209JyP2/NLubqrsR2bx1bjCW
xbpasrsTReYfRVTcgawRxhocuCSiAapbdXKf/wmRhbaCtm7YqC+XPBp+j5J4ft+s
f9OYxz2za0y0WNICOAVleoQkU1km43NYH+qVpnw9UzvwTM5cU5qPPhkI8hDW7X+u
+1mMiOi+/l6v2oqkxMwAbfZbcJIyYSW7JXTZHMUJvoLCwE8wLw45bnnuD9/lOhjJ
9T+7iDPFBiM0mxe/9jcmqZgEuJgfI3gHOY8n9TPHLVwU8x6Kye6H2nswimQKoP8+
u9FuPWZNrKPYU6du7y0cg3IkBzKFzgou3LPN4GJl3CMcOMqaQTatnlUnuc+e3/3Q
DZXiYOBP9Ku5Bvg2dlFeA5iienL4u/FyPlp4XztbgCQaeAd9nAJHcvShM2goJ4QZ
jMxQHZsgWnFBd8Ilo5WksSsPqEgLIiQtP16REFKO0kmZaMJhv+uKiY4OKAmAo9Yt
dZM7JkyeF8pOsYn4h2WuEJjgJ2nJGbKi2wk4m6+itC4QSopF5raywgQOgSCi7/b3
PoMJTlOqO3hZYLLEWaoAwx20mBrpRMcdUUo8SAmjqcne0DZFPhthNfQ9hOjtWeV+
wcT2HFijmh3h6PDOVeKDlt1s9Ymmaj6qX9uMmnUVMC28kyBkJHAA0jpSQlvOFJkf
FkNSKu/FG+MsYyqS2yb9gz+b7wY5lif9AN9qvtoaEn5BkiATPz6a0b2F90e5GQ7t
CTGutOmGuPce9t8/duzJ2HcIQFTAZT3js/rQMRezixUFahXhJx43UjMclOFoETxa
MlQYzYJfrKLmk2dWbHedNvO+nbRLCVRSH3az5ldXgJNWSss8x4nVXXCfI8PNENWl
NPSpxofaUA6mbXua1pPQlK+lyruPodN81DRDnZKasz1uX2zBJpuqn42p7e4bD83R
fUEqj9/ZvSa1umwk3UsUYu6AOB5FqOgTLtDvudcpIxiug2vxG2/ihjr5vwVe3Mf2
pvGQGEzsmljsW5320rbKbaURlIR4ZyvQQTk9xAZr6w74ncvgG+GUQIpGG03wWegR
EC++YOrXMojdMMpcqnjKPaZccOREoOdoUOnU2jxMcV9E/IQYvAedOfakXPmmcr7T
hmJHKxC2d7OzhWmQaU34UqYt+mQynTw0LSaowuv3KPUySoq/tXqmlVoiN22Kk91k
OHUMbHfCLFQ5M+1hEV6VrS//IVROXwKRe0jm9TfDb3dsjS7fNwZhWmhAD26Ze9BK
PIzRt/oczi7ad4sPw3dMJJ2N1kudeaYVzdYNlEcK10Rn60GLk16Btzuu3WnT1PhH
sRxrr/FgwYYoIV5Xv7GJdEG9IWqdAEaS2XcJKre0E/IMiytoZ52nh8bHOAxPRGSP
0YS8UbRstc25hg1kKXPx1AuN9Gh27lbj4jy7X2/vz4d+X5SY2vNQtq3P4GPUB3rz
WKCvEGQz3k3EJs8MQPEsKRk21QbwxCh0phLkauuD1GpBP8w2vEpiFKgpSkbZG6KL
KwW94618tx+fASRS39B+xUMjs70StEuknKCrUa17+n23fBS5wOLwGoLnRCmmvoc1
cmU8/2ZF/N/A5az/uooJikWoAknjhwTLsrLCqyLrqM5HUjCub4tNHkK6C4ICBsLS
OWv36FfEyfRBL8ci4ngJP9/NYOUk2IN3sm5TIEzR57QMUZoljJc1LYaP2LTORHHk
LG5JDm5soZQt4eUw/CUOlCnkG9O/Pt2n4976ztwORvQ84cRvifikyKupkfhVK0Jl
1vBpUYn0xihGpVSeA0a/24anmdhZppQW2dG4FYZ2bEhQ0KQhMyE2dbXVUAUkwRSO
0LsN6Yd8lh9kjECICnsEC/X8+OpYmFBL6zDL5P61zpp4OgV/+0X0yCsiBh0Kf50T
gXNswlzxRaP6hvlYn9HMXOzA4mIBce/QLfrDEHzFWxGHfCkIVSm2FCz7V8LS5Ys5
OCLFZCYuZ9jGezckTyrYHhCsCDRAxefa0CCjnCvhdbJPoaXEFLtQonrNngmoZ4FU
ewzCYffFrocaob2hXJqoAaDx5pYG5dS1yuVVIrZIqbr3RXzHPudATFvFUQj07ddr
J+CBoUe7Appqo7TtCbWYdx2Eu0NvRZPGlruw4P+ZeAg1hTqW4Rw8vdM4whEbhYUg
vfGhh76ecfg5a6qud+LaJbYs/UbM19ZjX7l1EEgS4lIof4hgq3a6UkL0S6aBhxVa
Wg6oKHv7Jv3wfKuxxX00OuduAEeDgnFjAgKgKWSriE/D0JypJ6wRYJcjOFRiVg9T
QY7pWxrsT25FHItAS5Tf0MfYlzjn0nEyVwtx4F50KDtx10T88Cz5FY2YmDR6MWiE
XXNqvFMjyKN9OBa3qf4Uct2cnlgptYbaAl/gTiCDlRau3nVXg5yhaoK93fJC6GrR
4ctf/NfpZu99EazbgWqTUC+6c++DlUB7C5Cf/PPLSlRFygRN1XQBRb7KrloqmCnb
+raRSdQxxZRXlhzpTM/mVZs4pWoxA7INPjUYoyS7vOpkTzkki+hDiuOVUmw9Ejz3
f9VnbKxI6+M/vdSn0F5DWDL66XuiXhFlWZlwTI64GawYLQqkXgCJ78IhH/QT/XxN
fzIrnQoTG1hYHBf7nnU6vUd2YuEywTXs3qD3haJ7n/R8skTYl/7nHpE3YqLT9qYZ
Ss9qD/pclNbZqnqUAvVMfgSEW9cCOPJRODt6+Z7sIToZOrZQfUTqim37paAef1io
dEUG75W00xOWaBuP/6jaedaOo+Lzx1vAj+fTAqG1ubGKiYQvOCP3lL1+YZOmVnXR
7HGfTjLNvvZ9IpCKXp1pZXLdmdJhvzzoBPN4rmH3D+uENAiVMFe1iAJxCWf4MmNw
fEMqbWzxVe1k7OQfRHBhOdsHMLdwb9XXJJxijXO0lnKZB8c2TwFXJsbS+VNrGkVR
tY6KpKH1+TVm1gnrSC/eG5ss+ZJX+B/f7WtHoHoxkwJQ9EgFEIfSemaE77nQzULB
kshuGN0bmIhXTnzJ5gtLU0qHuqR6UJ8pj4TyrWlOmeHcQk06OKBtNlzKqgCQNWMN
xd9QpMIg43kKeatZGqibZtGpY9w4R4vede6m4kuipWBI0PSJQb3IMG4fiyquFGla
SmxTE4vfXBPc9Pb81ojbOoOQMeCAQhlLWkjjgmt1xkMUCg05U7QNhST23MHeqdP1
AYiFSTi7wI2EDWeVRtyk/2itPcjHTvSWTXr+Q300jCFAQYyPOblZdZ1I6cafDUaP
xIF9kHiNIPJDghSt0UYP7w/v0LDmSXPg5k3wchTCfNJ0zJfGGr6Z1mFO81KXrk41
UTFYqhMeJ/b46cqxqMPW3/b9NCCZRlm/rOSEnRLDg0AH+Aa7sW4He6Yf7mssrqXj
9yPmucbQJYxdbBX9MG4Jv1lkYer7YgZVZSA5WZNdml9WSAwK3Mi+XTMEiX5+CIW9
Hkv3TUKAyEzk5UWj4NNX3APF7WWzUs6cOVU2VY4FUCI5lMDJh26+FSqDPErOCqLC
GQNLRtiL89GmQbxzSFYggpXts5KWc77qqsVWaMVATSETtXGBo0O5u362eTiCB0P0
CtAtLQRdoKPXBFONQxjv+c4L0jWat5UkHnmYbZKzBMcvkCpauyJu16h0nsCgPfGX
VDCaH6AVpsuDJmDCMVGOKGd2gF88bs3DICTuZWsW2TSVbjlW74I3xet7I1cFFR/S
ko32yt/kZ7iFD5YBBV6Ec/sVk5DFJNPMcLqoo6plHtewo1h7+065lk8WxjBL3hdW
tQOlLFueu0wvUFD1Dr7DJ2SdfhBoHTowwmQU3kMm42Hd3CaPaJ6vp03LTGKFb95R
E1RX88D8GAMUxqVAKCn+uVbdj9bZbs8uZs+Q+yYqWXWF4arTm1N2giHRGGGwRo1/
vC+06MAlgOIMO4RIEUhgXiCpVfZHtAXpn/F5abwdvJdOdC6L89kP4lSYskJ7yYbc
XHHJ+m+WjzFwXqi3gm3zYs0ejmvVZEyyw4tIOMFbLJMTrVQ5WFMEAV9FHUFbPlNz
ie2h4mKbTG8kiXKEH4Hjx559XPPVSeK9QJPFBjyRRrWSGBYLeaNYbnGo06L+c8AB
48E0DXfiAP35E1lTvwlZ/RBPzt44wOw6SeGd/dbRhO6q+fADMu0ZaVe0VD+jm0YP
RDKIZZJyJDS0rQBKzaRifWdN9xNgyIYZeUNDxgO2L6fWwluJWtjO6tfTQAQqD7d6
/DFLy00JwAB8ydeSJgxnVzOzIibPZlKZkCN7eiRcQuHH9TKd4uikkCHtN9aW6AEx
dXQK1yVNV1Z0WEt+oNg3hgsb3plJ/dNvoW32a3yzvdCsZmgRKaSNJDJ5Vfuxm5Ab
9DutUhG32KqEiWVB6jVnBA8tu1CdLdsfxcr2J19jKogSIr5WMuA1dsQl+vAP6R+B
k5XxQxusI6oT3USE0h4r4j0/sAeC3AQ9ireVSDh5crpVZhCWe1nb5pfpDzfmdG9Z
QZorYtDd9JZeJwQjPzni1lXOPXcPaVpuVM85hByayxB4ECLTiSUufJcAIILpkqzy
8hkt2i4BsSGEZWmn6hWNXJYnD64uSxnGYaVVeKO9tmIoffQp57OYmu9M0W91vKO6
dLVMAAJLD/HCZ+vG2n+78yRzDLXsDNVmy00cWSTu2P1wbQH2unIHwR9Q1d5D5swv
b7vs8G0oO2hR1Q6F4/QQHakVnCTwSnmUoJA0kSR3dmXmBPMp2QDT2h6CwcP4VDsJ
zNn3lwWemMjlsnM7ONLW5WEPEG3hezr/f67WUCs2N+DUKq+Qb88qMdJfSvGm2gBo
KkK/WQE3T81mJNt4LqIBaorp2LW3TTllo/ZW4Sg/mn1qSm67H8RY28b51c+8asgf
aA9XwaL02FnLrOCjxKBtIx/f0UBaeEGlGeUgkZefAPcu7aA46fHBF69JiCTXiKRm
FQ58pxucOK+rUJpe5Vhz1+XQZwVeob3ZuG814tguVfPN9T0Fu7diFoUTzAMdZ4FU
z1LgqwD0ELeELxo+L80BF+MzQpLy51WdKyg45p66aHIvivtBOuDdN8T/E2YHFtof
wbUKOCpyHIghjX7UV4ytxLEK0pnUdZASdTzSMDxydjsJSfBrf2FxFV5kCOKDyUeC
dyjS6o0RRhayAUBscazBYrsIG6d9Tmzh6Cv26qZt615hGUl+acgIwBb0HBV0a2yM
Lf5eS9J2JH1LOssCEOvPvstcJJkvNi/KqhyByTRoP6ob6y0U5B5cqShJvCN5O6kf
H4TaNydixxnsYaK/+AE34j/OdTHRpt+ImSxc3C3t4uq4/fhPjMo+Vp9+e6Yh8mah
6Ihd2LXlf3cY6LG1TmTtx79CXNEu6/qsrQ+SBr9/J57+Kazk4CS5G7ZsCocOsZbv
/35Unazciv660zp1ut8GCeGx5DAqMAZnQZpH5Zj2JxASDQ6ETLaeXzbpnID/V0D+
VO08HyEdq39meuVSJgmHfOzbmXyKM+72SdrolWT4uiTzRrzJClL0bJv7YUdgeNVD
FPYB3iJCB+QSHtQiUqCnF5Rnk+jwOJTE3swbjeV/xBnBFwOnAA3fomtnuJEiQVP4
333ZylIQb2qI4oDoogWC1+Ii3bbS+prlLaHJK3akBTXM0NZ9z12AABfesh7V0r9U
F/VkEaery7My58YNXrO5ey4KyRWVE5OOLtOl+GETYvvUMS5TTwxoe/mcV5YNh6EP
RTMzcqYKYtHPlr1j3BNx9gZerp2QB/tkpijJKCIebA/M1rX+hJ0es8P9+pgsegZt
0kQIDBgfpR4md2GstGiCOA9gOyf1G0FBQU+ZAl89O263atpueYuG6mFKEN6n3UVr
RbLMET6QoRCchfPPjaRxAZNLAMUmvPBGVA1dNGPWO1AXRwohFO59J1wfyGh2Y2vw
DXakXp/+3Pvgd4wAME3ZQoL+34HRtkue8npyHm5qGQKini624BWxA4crFVoCIOHX
py6WVPPisu89rSKmWdSC8iDz5WvehzGglT6yG8Zo3mtAzW7qfT+IKb+B3P+0lsmh
icsCT8sHWjSCDtnhQbL80gWc6zTXTFxNfvUgmWVjZhqwlu/6bUEr37e3npplIXtQ
3WnISU3y+cF3nPkXaXyrYtS8lrMK2oRJeb9Y1o8JMhjLKt4Yiz6K5vy/mnxzf0R6
2ffND1i+Lr96xfVKVahC4SXvXMbnKSQJVsxtcB9F1yghJEgoZ8ktbQM/620iMMcz
bri1DWJ1N7HJGJbmHGq3ib6NUk2uyCk6w/8Msv11y3FY9nhKVY4wOLrXoI3nMPv+
INkTKX7spCoCl2nL/ENLfSYno3uJoLOGyM1cyW36T2FCGyEfarLZKnBBxT7Tx/8d
+dLl8STv+VjJs7+p1ZBRxeWSNRhJSB4B50Cp8mq17aheMJI0TC1IeE7nv28ezlln
T89i2Q1tEEnaNDJXzvREL0j1fjRkj8WoBCuPn4F3f8lY4ZE1XUAVtCNwHUkg1Gfb
v4Bf5gCkGDkptQjKEEV+wRqzN+Xe4EGIuQHBD+P3bX6OYjnyVZKq5WE/ncOLJY/f
LmXKjJzgdwn1Uppc/dMbkQ3CClP4219H2lEAGbdtRhZNAKTuh6SoWDp/HCDI55X0
FHP53PauV9WwHUFZsdNq3TMeWJPxJPELh/eKKBeGwmo+Gca/n3TRM3mSTC37v2Bq
qE4hFBkSt15DTBVL9oawovJghqCv8JzrBmontp90D4I8REwx5OOkRS8+N8QrmD+4
ehj9mn1ELsd/Y8d33/H0gndsuVriPp5r5pOVH3r2/RpK4s0v5KjwYWo7G4LwyWCN
AVpkCkf6MW/bSyqtxr61N4uhkFFgWZKhUmFo23nCAequydvPLbsidX5FRFFBlv2W
mL30wfq7dZDKvTCuINDTIpFaJpMYtsggyo+g0bqi60kFq7RwdspEZKGwXhtT59lW
R9ufEpIfujmQm58UnOWpZfAAzvfG5CbZhRjfItsh4+PX8Yjla2eZd5AZxeKkvxGW
6MQpcIfo0Za0rG/M73Nx37eIr2YeAoaOZc2IpU51a+gcOqCQ60exq5MXGfL7zCl+
i8MQQMNFtv8HiIrWUgMlH+ZD/GRV8COsD/PjKs4F5ks40PlmRcxu3hnBuFOq7FRi
YeVl2lH73Q5iGoPydt46DTc/gBxPtphrBegjg8ENS742/A31EUfGknDG0WAAXm1M
g5aL1vtLnbdPNCNPv+6v9zmV7cGAfqpjiIqhSj5pntqV1Ga0u94xHGEjAk9mi52g
/R4uHEhIBb0Jam+brtzjJuSk45wsYGliVJIC9vmcGpiD7YXIEFTn3fMjPMf3toy+
9M2K/4Ts2WXgIxfqA947cc51vFj+/EEUfxjUg1tjg1nBWyYS/nN0iljXbtp5M/tC
dn2GhmDKepAmQ+TOF6V53u5g/qqAnMMK4rBc8up48M2ArjDMDCGaEc/zECBV8N0G
60Zj21RTJqTcxKjYcqxR6xDqvMhetNzBo107e+4dOK1nMh0IWPQGNQQ36hyiviqX
6khSQjD5ivw1CACEL5DLv7iMaNMlCUa883lPPM4Tw8JPdSiBkn+6W6ub4eXMopOB
q6mvTSbfX727xvnrULeAuRXcgMItukyiyyUeaPHwRa2oJBI9AlTqzWLJ94Ll731B
Q4BourFq2lH/Oat7cHowkB5ZeA0mqKBO1s3I95PvAI0dAGl50lf3SUAN4x40Oir/
CpgaFJF+Xy0ua+NIfC6Mffr2E9rKxVkHl4RmnPnXgSpJ6CpDI+Hos6Faeesl3ZY0
cmHV4UATgYbOppejheMVHDOACnfpmQKix9BUhMvmfn4g9SBfRnJc69Wl1gbdQHJF
wNmIESkdRQ3rWZTYCdtdGAfY/I0xtTO5BxlJIRiapNFcbghEVGUT27EeWEqJtvNE
uyWlAkPCxSs70t9b1vpDoXpf62yGif8C0Fm/9LKjd+oZpZVM1RKSW0whLLfpLSqX
0RDHIUdgcle9PUUaohn7m/tAR8ovXQn0HlKn/moneJGfXohWuAm/iuRJQlX/AN8h
4ZuzcZgkbGWinAfXUdd58eCHKoafB17WVvIEWZP7NsY+RlT2HS84JJlJ/JLTZesU
4xRC/oo8ckJHyx6WlubOpO8Y93v25gQGuees0AyR33XEF9AQ0Q/lbL8tpMiK2hYq
CBs9y+h63Y+rU17X4tDo2/PtR+238BOyofAbmDRbyKQWZ51YzqpXex6kqZtAmSkK
XoZeyPCHQNJVBnIY4ijGHWDS1D5jeYzknYWQMRRWPEH9qZOWwJWuwbRqRih58rZK
DVzysTkSwmVIIjNlKiZ8bwnuqttybXc+uVWt/ebsEg6x2pJ8jdRFe+SxVZMS8hNj
N81sH4KtKMUkhY2Ul955eDcckar/S+4BgKf2Y2zJDVlq2YCcL89yCXihEkTIJo+J
py/Xu+4tw5ohhk+RH/pO1tBvUzSB6V7QXMuIIIWk+/tatCZoGV0Ylljr6roValV1
oL4K00ngYngmzp5OpLsRkSZTR0cm5Pp3f7DLPOSdOeKK9VHo0pAxwcs8/akHffs9
89gt66vw8gQ71Z8a5kF3/+JQaI1LWKZWHBHrgzQRNCLtIOGbGByiPe0aKhcR63AM
QnqYqdileIwxTwxVQHdJmhz4eHVbLsVQxdMXV1tbXAiXQ6l6liLnXn4y4ZF44tvE
AWb6JeyIOZXsrO9F7gwFrIA1Qj0c+esIcCWX/r7ISOFXX8O1I1Pvej+mJddVzddf
++5NBnhr/HHHjCOqxQb2yC5h/s6gbniAwMD+uORNHTm7rW41qyp8AE95MJ1bfoNn
C1jS3EbMueSwdfhFdWs7pUX0k+gWQeC6kIPiKIyu2SPy5z0WlbmJig4f+DJP8BI5
EvujplS/RDj64gt9JhVbVbfxcAIfS6lDkR+UGayyOJuTzeYVTdnTUFcKB8XLtYPa
js8NqUCHwHwJ/cTSKXtl5oZ8MZZ2rlT/G7iYXrX2B0q+jfZszEWvNg+VePtuFt44
YFLHI5xiZafX8FupwfSFaY3Q7RxArU/XtHvstmf4vJ04opG5xT5PMab71WJn8fHI
SBT2mJJEW+4l+qMtSJ4e2hm/N1axTbNF5s1EpaRwOObpNF8ccW7yEMvxdTKvS9zo
ebIw0TT5YEBkH6jqvV80dWchBBs1EtcLc05myWN2UxulmESZk2quFbpm+S5XJkAM
9YFuMv1gTjz5Mkk3fQEn97EKKXvfR2hnigoGzUe+HctaGtpoJzVApusrWeI45ef/
zCvzqgiDVKWInHVEwqROeUd1n4aCytORgzpkeR2EhrTVDZmDuVnjSIOkPP6sikvI
OL1Cs24Z84T88tgV0VISVAvrfJho9NbZNOu/nygB9LvSIjYHbPDRG8e23UXAT2GF
VLMdenEoup6t7luwt6Vlg2wnXC7N+t5wbIznidYzxOujqMzxCcn5TiIzkER1r0Oa
fetayMPrgFsecrARKgGSJ1z/8NUExHPf1ZrGCSw1dIWpf/0KRNWyldDXNsaMPqsx
6CkeA/L9JTtRyiDiKjmucGuWaPPWI+APhoZ7XONc2disWTt2nCkmV3yENC5a8iq/
9kCgkt53rzgTHA7ULGXkCsXackZdGMiMsnmri6PhAwx76+HNO0E23nTVQQva6Pdk
nxrZUoDXHA4pus3A2X6cbPZpMwTyDipX0NwR15PlL9jHGKmJzx7cO0M17gyi4ORJ
0ugxjADqKYr02xenUZJgDxhn8jDhLUgfGQuj04zcEHCVSLqYNgOSNwifvyszqYHa
fqqRhJet/k1V6AEekePHDxdruwt9G1ozC2PeV/noaGfL6g08GEfq9qYKabAxGTc9
Mrycu79cDg+oXJV771nt4QoBpX/XJhjhNORGtozOtlT+FRXLwG7ePcWGuKmh6cc4
67t365zRUWf4ilKMEZ6DnpRcJmbQ2h7hXQDE8rqR4YvIJZJEI0n1bdmY6iehJ840
DshbMP3lTAbv11kVtDL7GhinY4TCcdI52i0qMGmYdis2p/Lh8gSnXiK52ITMjgQn
098Sdu3hOe+q35ZfncwmmC64fbEdTK2koaL3M3fRrcEMZfG1lwRldHzXqfiRt+6A
BUyTHh5Y29TmxkW1Vt1z3gcxOSM7SwEo6Yi1RAhYrJhBMHAbhJmrp92WQw72Osu9
mbh1ZZsdvKteebzTf9/BAHCLN0ZoS09Klqqhsnu4vv6w9YM4za1wO6wFxq+bGNOd
4+ooMbCBUEEE41Ut9vVFI5Yyz0oFrOcuLt9GYQXq/rA3mV6lCTpM/VvnInSVYBP7
msw0Hjlj/SxW49D4uRAV0hqNMdDUML/+tYDM5k3ZM9ZWKOpzQgr4vtt9b4AmonC1
TAjdUgXMel+Wg7092aTEwKu/Pi1bYZqBMIhmhs/B21sybI1+KjfLsCFpxp0/bguW
b97Z18IguX+CTKZ5y/kiJrCShqkanJKeWhP6U7DzbRJ5mPb9MhiUwkMQbCZAdmpo
FwRQ6APl/42DMJd3+0TbQV2gPRWq8bez0JCCeDLkBvYuKZtSnETsxPWORlDbL8j/
ucIxoqRnBtBoBaHIKY0uCnH/UQC6mLPxO9ZIlh2Awn2DEYVPwQy6Tty2BOs4HxNN
qdgcMPgM5JvjJL/uy7heSpYxfxQrGMaxHiOE4CiCla/5OuUt1ttszZQvTqwgkJqB
ZX/Ta7Bukk8eCjXyi8jOA+GHLgxN4xu4sgBPRvLMMxOTy3GCzqAM8dCN/iJ519Tw
V2KR3MNAG4KreL+aNtspRX82xfhKMqBOw8zh1RGPd30l1IQr69Tvr9x2w5BueK/6
XHztRB9PPPcX5MfQpflr3QwhAgB447aXPe8gCusc8YRq6c2N+qJHvzJ8L2gW0N9X
gMqG2h0Y8wftI6Ih8jBDAndIaEk+RnL60UPbsLhykVAeMDj48SyMsXldv8cNTvdf
uu0zAWL6YRlYGUK2AtIP0F1NmBll9NQVp6r+1Z27+uGs9o99NMwaPXlGV1t/QvKe
6ZVwfXtA9nx0mxs69TrRd0ivfXKUL1HsZy55EKjPhNnS+kRsI9uoWC3pLW8bdJxC
9wEfhbPwvOXa3KK6RCQg8fovnNa1Yb1K/Dio7uiFj9q4PXgDXliqJgdH0uWtTvag
qzwLpnK9hKhB2koqusHng0v0A3/Uy1uj9DisHF7LU3OEMabZ1B8fFeSA+khlM3co
Lg+KVhpbNtjpEZ/c79Uw7IdeCTI4Pkxi+GqRhYYHQ3hdlnHAcHkKKLpgPnfKSmoX
+4Xg+PRsJXOkEkYejfX59Bh9yRj/P03lh4b6RgnsJB98j1aHJFQbRlDiLAJ0fvqY
1QTc2bGwVnJfGtZO0TlIFgtnWzkGfUhZUqift8xsYzM6EX2k+gDOnPug7iTYEqYc
ACJEK609Fk0esuEAqhJ3vzd6CDuTgFafXB1dhlOYftJSOL0Y0mAFbc8Y3LKn0w5q
bWszZZTcLLS3CQ79AU+UkyKAG2+SMsvZo5pZqiMHH5Z3nZqatdkXx3peZ6cxH00m
lxKyoh2txN3HOCVeUtsHdRd8CrA9QWuC6YKLpw/UxjvTlQHwzZTwGdZGEPmZigVW
LYJSSN55bQ5pIm131Tf1fjBtfYYjQIbeWglwf1JHF0Z0wpcF8GR+6qec1dmA8jAW
82s4SYMEOd+fyMPU9JjGaGQc1keu3abY+LNxUikG3ec10guFstL2Ez8zJWd47hWB
GKjaHZD6SuHw+YTFDJHLPRSdmT1ELoRtlAIwl3XaKH4P5tdUY8NJvfMNfKD6TYI7
eUVY67dYFN1uwErIGKZQ6q+W732rUVKyro3/CEmyPKrZjfRbowo8udYy6xLRhHUZ
aNO+0iZ5y96zrOfxJwyv+5p0XwgSrob61p6FZx9/y8RARqR1A7jpJFk8Gl49qXiY
LKQxW0pMYFyXGc4URPHOxF7GuD/cgAdxVgzebgpkVTL5HXcDLSk2mSNkwaip43aJ
6fghW9wxD756PmLA3sGMPu+gsjZ7hLeMcpwXMWKhX5SJ+4rxUiy+AzltBbahcWdL
D84K5OVVsW0Lamr7OC3p5Qc0s8TGwFuRMFBVIhVgUH5ZA6DFpPBTW83mXLsHjlWT
7VzfJVblbGPlOHnGMQ5imogxu+oTfX1PDNonXELGOE48OIAlxG/537NZieqfIWhw
zZjvZ4HYPPxBP6eu6gfsRklqDhYQrpzquZbcuNzvtH0Aq4OpvVFqGv2A1ejlTp45
dNBIDZEGFmZzdka7LB0FXFbQ+Rlh/9dBIe5hhFJIuZYMkiNzoK3ECQbuKqD8I3hL
6TMnkVW45QXIyAn8n42ld6qz28fmrMJZbN3WfyDKPCQd3hsKyLlixY7dPOrDUvbi
LBeWR/iHdaka/KGoAnKfmmFvCbK3uTK9GLNxBWOU99kDdGC7TZQsqk4U547FSq+2
ieHydWBmgqECAuTP0HunrmLH07qIYzGvH0aLdUgQt+InJjlZ6yloesVOIZWDRr37
EOgsT7CIcdC8QV0qLK5cF+TPz51BUWDd9qZnRu5WrvEcVog9RhGAZrpPqMbiCpTT
1kIIPFOPhWaPq3FrUdOI2IJY5nxEUsYEP9RERrAubrObRSLCzLN6bv2PoKnvAQSO
g0d7OQe+KZr+ownbVpt5EnbVqLJS/v9wPVtYvP8oT03tyjOc3pUNleM1VJ6qZo5Q
/KikldFa10MiTX6+v7EJ5CmLGv4TF2ZoSQG1YAbtz9T050B7AzoDmZqguXlvs+dZ
pT76a79hbBHcqaMBQvqKDTogYSSPgEBy2RS2KoirpU4VwAAZjAlY3nFgPkPoBC0y
sSBIYWem90iOsv/rUzqR5lhgeWaAxOQp6MBuep3q98MPQuOKOoqcxFhjUOMzI4Db
44JY9JroKhO8T0iS4Tlx8PotCyCfVvJ3f58GM9Ad3uS1C8p1yPbKaDpShnw/4FBr
WqQ/k2rIhpMdVct/o4XoSuG1nVhbCvoth2ZLl2OFSk7VYvKYVD6rU50Mjdlg01dQ
Q60RIHMUpViIXBuBG1cTN8b26tbZUePuPGa7NIl0Tje9YYDysvOcXzIZ/jaP6Bms
RkOOAlqiu7s6lS+orh/yIpcAf8s3pmJ4kuBxMDkB1bzZ0uLrzGcZ+LAeFNF8Z6aY
TRxlGnNMVOgZlIDHUBAjcKxfQUEJzj5Gbzuvg3RDQ3K5bt8PJEKbCOH6DYfJTIG0
fixAQCs2Gy7MVPYJTIy6nN9UiNpj7v3HfkgnbiR25hAe0B80+Ot+a21pb0GtYSMo
XW4B0CvtVnq++KyL9Mq6/W6P7yVRujdo8oJutwTR7YJr/j//Mogw0GdMbYh3RlIS
LWQlFOTkrytZNWe7inTKleNcSPugcn0YKlj0QSAfOQPxtwkWQs91iFp45ygvIgBO
Yo1XskqWwyKGI+xIR5lekPFQO0eOgp64pt6YZoKVM44sIuohLZ6XWCToKOl2zOsp
Mu6gWyWXI0mKCFF61NHPdGFvdC5yK+DYQ5VH4ewNPa7qnrN9mcztz1gIMLCNKDz1
f+DaimbMrguhC/IquMOmI2beXmw35OuXbEpxj+4ZGF8E6jlPG0hw5JnG7QTldcsM
wNs7wL+cnVzkrYtbEWm1j6wz3kJdAAMO2fhyXIyD35b5QfzZmAnudWrzOOYG8H74
t9gImi/AOnd6UD28jvm6CuEB+lLvcXV5tO5QVHw8VJzIlbRqOgElIMSgSTycDmZn
BJcSOhntX+urPan7jnQHmgXVhNYm28DqnLI3OrBEJGiQTmepFtIZ6Ig0mKa+OxYK
/3cYe9A7AyxLKR6tyvCEssQ/G/VW9+uRRpWpA3FXTNQNuBYHVAiC7wmJfVz5YqCP
uT5Ci7BrPl0hShVfkgBfAmZ5GGm49WoAB5Y37+3xQViHqk3Nx0kzUe0Fjy39DuNA
sEyvkFLrdw+1oHHYYybN8sMsf4L7s5p5qUbU0Ew+qqG3LhD3WQ+vwg9UfQqSiSE/
RtPgrhR8r7upyu9WffYZDuRGs6Vg8kUxg5q5qWms0OWTcpbAtpmVN+qV9MUBm0og
HSdxRUMB7sIKMhiJ4eVEhCY+meXRQYeDi0xXvCHdghgrW3A6FO8eSNfEOniYWkO1
W4yQLLXtsL4STnxPDw4duNI/KlIJL9jByIy+Zlw7TMtkwrrie1c0ZGnW1E35Kbrg
+3rJaA+YirMfBdiK1WdnNmtC9eKUaS7ArZxGFLXN2e2VTPq0RipIfy2mNGx+urH8
cSlrHcoq+XgQB1udV3ApUExeAw0IN0VpmT1wNuR6ROFihUhEbZ7BTElmjxtQKZDz
g4VJOMNgExWxYEM0q2hbfhDCZFN7f1fgMu/TPDmlVAAD/WJx0FBqW4EVBR9CuWHt
pRcAnwtIso4vtqWbryjUQwafjxE7Q3j3qwmyEHgzYXRu8xfF+ZY9e1ycnmBtd3FI
p2QLl2AJjvL/xo4OW59B7Obsu+Ga1qkrf1egRbJbIxhyMD7xmpoM0gPSG5M0J5K+
Xk7YRUrQq2UH21qdyHfLnjA9GghkDAmH/nLEd7EfCPOiZeyULq4990iXx6r7f56z
KmAq9areFVPlKPbncpv8jGxPRuUlg9/++6WB4qvtG2cfAhXKQ1xCTADvw4PpubS7
FQkJqStYnGG9VhSR70nAgGDFs1Bm0c8oZCLPO+PeG2O1N11421BI9wrOZ2j7x5xp
c4RtpvFPqble3sdDXQiiUc6BhJIN7jFHc2Y8BjdXZmjcOS28TCrhqxhyh1NJwSpv
T6rAx4M8QyFC98PNbxySbd4OuwrnPTiSQFF5qVfuFdsE42KI8rnB6TNbY0MzKi1I
BRfxTcbb6KYmQzcnCn7SLFybT5cZ2wqyyt6UsI1i45i0wBzfOoTJg710Urg7m9dc
VfcwwZpa//yjnKoxtEWik4IzSfkDtIJK5U6CMJhQidFlqDQXCnTGp7rBLwntTzXC
HezMt9zBTWlx/N4piG2I8vIE74zuel4bH63w5qGvkrt3nvs2YFP4HR24Md5uuiYC
Vsu9YQFO49hCb7GEOC8OHvp1cpWj1OJ36YVAd2+Eke8vX6HuWO97qvhtp4T2KMXg
WMDpQXjMeqHRq1m5JuzI9KRafEzy/3BlL+vc2kdpNoR9p7Ck3XLRQVqH27gdjWsM
OxNPGKybQC4aYkZ0PDbJbru4zd6P5DZJHygC6Wbas69IXuLQLlSCmxbmLGDYZ1WM
R3KiY0cRubIp1UJxANhk9jh7OSwus3jo/+ECptmQFf5pmIrZuB9qSJqbxUKZqCyw
Z+DgZCrQwQnMbZw1G+zhCdFI+kgCX3j9XqI6uunBlud4WZyPrJ/CwtU2nQk7PDxp
voQ8aufW/63NePPuJziYNlGqLPhdO/qqe/fu2JdYWKDCj32J8nZ6FqbIZMUTHjot
uZEvOyG53kcRSQr7vC14r1IPOJigQDhT/VfgVG7ALVxp16iwkJjSu9Tbr1mAVqpz
rRVCuBa4yRb5u/4Y0BDe15h43aQukTfYW/UTFVN6CuvEql3s90MC2fyibxtfLKad
BXxPLJ5W9htH43772YfWetetFN4gGtlp30LwOyRkvEjIjHkYJe8NA41AmjLYhXYL
OtW2rGZMuP3hqFJxVNIRGepP3t0+64j3pUexsq/GXHCQSx1BpNhLdW/YFkx7/SLg
7LHdZsjw+ikHhUwVzP/spPBlnfprHVY5SnFJUEfscXX6Eu8w0Bg0f7kEkVyD6o/h
M6qNkFDe/QysAAZGIuXD0u4j1Rh6H2lorlVkU41erJNubkZrqDr+bHsYnfI00NeD
51RQGMaX3MCu43FtiAbKPBFqIJQ8LaOV2hwYFWiufoN2/b7X2NBGkat+Luq+MS6s
dQN0uvGizSrKa23rqtyvOH7iE7T+102HBXw7vJ0f7RuuIf/wL/FvagiDtWMwbp6+
Refw0nqO7VopWaZuopQmHPpT/8tT98Y/8NxlK4AEHir+FxE6Poh4xdMZvjZ468K9
CtXmDGqR/pxLMamF5BJqIg91WQmLgfUkHRCopcxWcpuxVA6dlHCLLL3NT0VtBaIW
/5Na3Wtq/iBYNlBxDQ6euLrUWCwkRWyGPz10g6ubocDoVkOQoFbs1swbHG96/zOd
EVxYIPg8EmMnTa5SQtQO8US/xAOb1SdqzUZ9mwGt+SGlOoHa1DpbstIGom1Zc+Z9
+WrUKcGrh+Bprv2fqelT9LF3g2mRdJ6+Nnt0g5vBjO72TtSnv3HWQhFTgsX144nS
SPV/4bmDskV34o3cW0bgsN9lzQmDDytZKvhZbRBXWjp8i5NrdbJyvGEplgQSnCt7
LOIjp/YoKPvhiJ1uAFFF5OZbmwDS29LY1NMXJrCJmhOWZrt0fRQi9rbPmu1Jt/jO
SuTQggxcSzfDhc7Fh4yL9WaMAKu89tcKvyaJ2uj3YfRy3lvDlwt4TxW/T0tBC26x
OJ9nd3TYlPq/SKYz1EImpmnAf/HlsMOlTCCVS4zPavVwG57nNf/5tCPV86TphEQX
RVGxzusWCQ2KSb2dDA9F7AB3HnmWGAylS787wjVX201l//oF2qyHAbI34oXx4A3S
lvc7vMmigdHMUbBG5hri38lexqpLDWfZKqFYhcaCbpyQm1HpV+Uo0qyInTJqmBlb
OqC8rfekWY78SJpFvm5o+26WsaQWB9rdN+KxRF/ulpN9RAA2sakgq/eZvyCf3x6G
+xgODR6grUDkEQMH6RDDrR/5ktrPaVii9rPB1DmKFzO0SRs776wJInWbI5Yy/J9p
mHdEEzWVUSyZIhJpH0PspIAqNrod5FMj2egWDhqxOnFZ64UMIEiO5vB1915L3zvP
VfODLhhmo949gV3tjdXafkeIDSXo6grR45HU8SbYcMuVhmn6jnCMAfl3WB4KwnkH
hWQIk9KW30aQfDIaROj5DlhSGijIOhFxr86c0nA5LNA9dS9UEYwdMh7K4Yo+qkRc
q2JBmz+sSkrQ64e/pRCa31aG3X4Ve2h2PAe3WoQUoLPA8JtpK5WwXQOACgRzHUok
RNmQS2O4EKLbPRpjP5vMtwC3m62d47qV8XA0AeZVUAXCty495dRouVGV7MGtfwh1
uWQzCPrYE2I/pnPH57qB/fd7jJxg0bfJqnAYy770m0bFVs4/6LpV1DYKR5loB45R
xcSyhWvpXK+Mujx9McVBmmsehydcUvvMRcV3xIVa4Rr7g5Ea5bDUOAgnMsfqT8Xn
1Mk5XVQXxIV2H87GB1KEdCDvtA1hBm2k4gn08YncmGsmr3DQTMeV5oQcFvs0VTaD
AohkEr6d+jfmj1c30/myPabn05ihcnaeHM0VbyDy92eG5llVz4IpFjLxUBCfseRV
kot4mcbitw518Cv9DA+U1bJxFZP/RBCQ/NNyoAbasfrTQjgnjGt6cmKIhdhW7wZS
g5gnI+5QkLsK9LtuU7cYUn6CMrZannWu5mlUAN/IGTlZZ9IKszwR4qrwkQtAdSwK
zhNN9zH9j9KSyzdi0TQgTj6cXrpWxw8GUtrdILzkDdt5IGMTfz0WTsRu09W2QVIV
BqEu4CIAGDj17ZUEOVw9qrENDJ60KAO8PioE8LhtysD090Ki7ghRL+qtS9w8c5Fy
gHy/O1WKL2CX/2qjHm0eIPM6WwsXX1kprh+760koxCL+3dxmyoHSLhG43zI4ZkAn
CM7bqatayj+/pF0gD8F1hv17keage/PQu6pZuYLq8Jdki8QMeataQ57JbRDIQSLp
r60c898Cu7ZPN/p+tlw7g+Qbqor7bCdlEaVkLSnLhYzVB7lKr74XON76zUQF1hxu
Evk8pYsqnlBsOC+uYbmEvuUaga7Q2s04OgJjo9RKgRvdbFO/lAPj7l3PGJdC8vNa
XpuKJ99FnfixDt8jZmS4q4cxlfkewQHHqLgNAntZqhmSk2QBhtqw9eAwrwmZTSE1
9mSKPmcxJF2rA2c9l3UqBwZ6+zqWjpeoNJpHrJnE6RD8lQSeWsZFsK07WU3DySrj
n8S5Aw5X+RMHOwBTkD12HYL0ClUjXaUO7xuVb0I5iWuhEQ0M5+D1vw3rJ+byW34F
Q2PDlYzYswoQmhfbQOHZvMP2RMgg+0+Q8rHxnkSyjJoYxidcRscgZJapgK+PZn6k
YE4wedlaZtLq7ZpFjmKdlvdG/hOTHu8iN1q8mn8AN9YeQ0QUSFZTSCLM7ZAszgXm
fIE/qx+AUlDQL+zpKjJAKD4nNBpKctFshQYxMXksjFvYeRP1jc7Zq7Ggp3lfXhOZ
mbeWazF3NE0DHMSmgSA47wWD5En4sK/Z8v50nPjHQYIdOvNz/vupitkbYOj8X4yE
srXpHJNhgDhF2ESlxY4IV+R4AAhEYs6wzO0TFR4bvJ3O/XxlndUZrVNHob3ehUiE
2DfV7vJjzJGwBMGY6aNHY1qKzGBXIODsLw4oZtJDyXGIUib7sTkjv3r3KCmkwW+B
7hWA8L14LVbRQW/elxMXuCPLLKbbGxbyi2XS1WnTjuC/ymHoR1Jvgd+kj5a6cV9O
h8UZm3H9aRLs7w13rsPgY+h+SvCNR/iiJL1uvu1PaR4xDoRQ0BZdDyZZjhYl58lM
2lPKSt43vodIiKhldOoLK16iYyu9+By11RbK6aKA9vVF8LKSPBbTUVpGD7CysZrp
B+7to6HLWinnyeGwIT1cwOhHN6klD4MXjwxH1lZ6iYte7m7J+b9l47lonXuJl6Ci
4G0GrqLKgzpljYnAZhgfYZi6jWAQSK/jVH8TCANK7GLLw4OfV92vAJDzsfcyOlVF
SexuxhKr7RqngREFNQ+X8q9vdZqFjsXQIP5a0wCv48KyWLlvEum8LUGJByOL/I/1
A0zvc3bwOv3kgrr8ypoi3fWaFMBr7RMXCKikjCY8zr8e+IOW1MBRBNIJbGiuZ8XX
GEKByZjHOttSo5wep7atlj36J1SUiULamkhyACYZMqUndacbaXLDmggUWg3FTWvF
j7MOblRfBOA5LmeM04fS1LTm+7DyU+xyHJOWj9AWujHcKPN1N8r/LPSM4dg9d2bW
B7RhxaSFF/D0a13ndhDqHuPDA1v5m+7Kw1Lm6cBuQzXUY+hyPE1GOWhBVh8iHzEt
hCoNlyFbtQa1ILoUMD1W90PAHZmzgKK2HO2T4j108dTD46SxCs02SkghByPFxbId
Kx7IFWnfT8ctyBp8cfGi78MVhBc2CJY1No5oZs5D5TooGWv1YkuOxCTlBZcTvXoN
TyHtq2TH56SRvWXkitsYZwj24VhMUUvf5kUqwTBzooB/AncgHozGwxMezY6VABHR
Iu2uhANgkg1/PQ9Ob9jDO6a69zi5+LgidP6pIjruHNfKZJB7lUQdZqvZAr0WXqFa
hdmewrcTOkdsCgA2ARw8xTdH/+RCHXnW8I90IY/SvDd0irQ8Kk+ZvotkCOgc9+kt
w3mBEANd9wUEMora23s4lODwyoFMnp5JXR1k4nzQrrbpXoYc9IVlj+f69ctsE4jv
stxHw9GjHzJNWJzUsjxPgk+2Sla4kLTH62egNpEcG8XR5MDt0INnTOrkXRkoxdB6
ar+M+Uw/wQ1JYTTUWdngrezbB+QiszqKXof8htBIltKcLrhLF9+ptV17c9jXeI1V
LZs7eE+hMAbmfWIyfaZkGb7EQx7wwxtdaZIReN4WN/7E1oPH1dEH6/yiOUuX0499
GqxAAxjBwGtu39LYY6cmd+Ndo+OO3UhMkKcmRqvhlxy6JLBZx9+pLjBjdLFzo3Yl
88wnjR5xnsAOLcuY6WdF13+LcWA1HftVoVYj+VKI3ibEdE+oqV0oeRTJn4h1P7AC
pXNgTJyqOio3wzbxl4qiF4nmP70agqHxxnnDVtGlk4pE1W7bJ40JvUxpfJ4n9wYb
4Zczp5A2xC5+17vjopW4mkQj1Oq7uGpTQ7b5onM9hZd1BmDyslqtZJ20UA7XRSSX
dqeewA0dV3fKDlZDltU+9yIy2oOXdfCBLMXRP8PeDc/nnymcvtxgUriakzRngt6o
HJq/XM2s7OCCR+mpWFPzjH9coitY8dnCIkExvGpQHlTACQX6BbuLk0VW+bdGJKsB
kVC7bUdGtTntzA9nnLtH0WESu3mkgYVxEojTIWuK56hN9DNKuOUqVBfhr9rIkYuf
9CkijwFtgFmydmYobwmzVpzVz7s5vqHPmCsV2hVPdIQcb4gXb5Mq/cSa9BgWZzGs
CbgKojxq5YMmwCyXTtHLgt3WWHLPap2iDFHkx3ZnEx/I17wVWmk2KrG7O85kIimb
PG/SKu/NLvGHqvTSMfC3z2H5LWXihDnFzlGbj5QU1LnrK9U+bGR40V8Tv6zAAwj2
Lr3G0vX1m/puU2IAQ82z4WUwZQk2CSkYsFgRDBv8CF3720PLIweFQqjxBmTECZMA
7BdOah0VI09fR2XBlFIkA2U4E+dCvZdTCr0RzHXhFTotNNnvd7XAu29Zuj+EMeu+
R3lB0S1FQCK375RcWHgm1vPBUAdEpsIpleTn+SNqCnhLf0hBEVym6mov9HxKh5tt
ilCh1QQVnEX/nN9bJOPOTGy5yU54UFYQmPzjSR48XNcktNq7puv+wiad159PlBlf
f0cRJHr5CecS6XEMiZSiH7N2gpnYEHLjaH/qEKJnu/RGt+EqIMSKr3j9T4lsp5XW
8oABm4tPSUKl2VMJV4ieduTMXnq10NEBcjF0KeYdPNgODLE+lToIk+QoFmIaI+1I
BoNVUxvqP1P1PWZy6HJG4AcDAS7NJaPL5EqdgmqJu+nInlSXcQMUpMknxtcf92Eu
C/YCKu31vXth77zy3G2JZztzgQb/1W6WFB3vD+TvQYPNo5zoi00GKbcOlKdY8xPK
psmAPVoev2MOQ8SxHMDVuTnAw6zpoN56sPZ+NbU892sLYwutdtz8B+Id6ieZoEHN
GJQSA7lTH7pHCnEYqQrOKV2M6Lx9xbl1iDynh9KLbULaY6vdnQL0Dfwv73DCUKC1
m66THFyh65BZnOYm547cl1MIQZtYtg6rd1U0HmpqSDdILWcE3JiIbMID4A+X84nN
9weDkKNqUX00/USRaMjVBrMTV+fa6Ej7LemfyFThRmEQ5P4q+yXEVezsYUvjj+Fq
f49pv112sO6rlMEmaSNxdSdBWWNRJzsy4W48S6CKR9xzkzbc2EPN2yNnKyVYadLp
/czwmQ31HRopUO//+TmCLacP/i5tOYXxD7zusa2b/dhqPHDeg0L3RneRqHjPxemm
3SOpwTxe5mdlW2XuLPJ8fv/uMVpx1Hj6AibdaCFuxThV+9NmQlCvBFCsHMplT8u+
NlKLhI+pcni/7fWw6EJR07prwB7GvxvRYn1XgqMOC44DilJYNb98RNAiu7t5C+H3
CiEe2RdsUcES5A2EjNePeRHWHFWMotM6zQXHOBHmonsczqVS2iekcnlG7P4hu92B
8HnskLKCIHn/nTF+8ohuKbthuPtF3TLIZMJSdiYba/q5U2dbOJqAU9XwgJ/m4ZQy
AMIQNe4XxRPiGO/XBX01zHUN0wGLqEIt3mSzMJQxVkz/q/d/JA+kmzy4Y3tJGf4B
UoElhmYtGy0NKG+Mslp0bZdcuZqI6bSMAUKC+J1SHCfcWKNAIe8C2NhDoFY/91Xp
ap03xLNmS5SfUK+i579MH4cgryvDNSn1+k0yxncsbskh+1D58aQrHRmg/MIN8v/y
VOeUQ0fwRarva6fQe8+Z75uUm0r4VNVJ0eCEOvO8Mz1bdnlm8MfX7uXF8jRK5l4f
ubuTLtpYf92D/lGAmvg1kbHn4l9YzcqRpz0Plwg9whrMkJkc8NBB3V15vghyoeKC
LjR06b7k8Wj3YnJwWDVEcmb4U1WvBNQII4IaJS53x/0v3y3WBS+4EMmZ2Ifo4EqJ
BhFObhlFnbONBGdoqbWtafNrEgvtkDlhvA852jMDEdVp//B83zVwbBXxqIWXgKlM
2iKydrFMQCbGxtL5QGqGbqJSNmWrcVriGAnEJzaWhqTeiFT36XOmyRCuyOwn2muO
6cZnj2a5s5Qt35RDLEgHgTo445XtRg73TTfXcRSOAzIolsoWFU1eGn8Js8Q72Tls
Yt3R3bwk5TcgjlFcjQmUvh0jqYNYwSRJaG/MSDugODWPMtlBB+W05QO11esonwDU
ZhW3ldYNs7pmCdG4MyIaaA30tyP201ULNLS4lNR/BVU0H2imv4i9ocrzW5zqU+KF
6b0RXdJb99NJC2tGFc0jFcd2BFluJZWzbmSgMZsj4hH2PRabpW2mho3lccaYr3Ts
iwXXwlG0KWX3ZiepIMO8Xm/gdfLAFaR8jQ6QRSw+dVzYGMTO2ROTvWyyB3vi5w58
Kp3k1R79qb3Lx854KHCGfurRjFJyXtIcldK3jI3acjNcMnapyXVDdy8IWjVXPsnQ
7WxaVr7SasrPiBPeSc0rWhYMgwIWSSw1OoYh2Jg7zTMBcya2cdMAII5kPg0c8qxA
+cni1zVwUDfbl1+P/Cd005536wA07NSqyNyRb/cSA9P6m+rWkvco98+Mcx9tHjhb
JFC/Y/axc0uOwvqFMJIY7+IkKxANkJgscazrnjvn19UhpyzLe5GSat+Rzgj0W6kR
B7uxB7J+q2df0Bj72dvRWgTx3PaTmpQHzL7IJ5hoth7bK/foxtQauylSA5Qmgu1M
bVXs71OmcOZ0nz/ePThcPh6qhFDW7ZHgvY+BVbJpI8dbeyh146/ze3JyIPUScrjC
XjrYLjXN/SmuQ4pTkexS3nS4wW0ap2KvMo2BIpkA8E0Fh6SlFXzlzGw38pxtQyHI
0Dyq2la7echNYwUWwHw86rrHvt0sEiiaCIAhX3awBwgb9flyH4fDK/QNQYtAaGx+
GBrMZfZ2iF5flM29wWZE19/nPZlxFVt3o1VzwgeCzL0HwOg9T9TfF1U8GluijS8V
5DPbx0LVhjVfGMxEmGSIt+FWspSvSz04eu61p8iGmxMbdQUy6n0IJvLBXBJlNJF5
KDB6Wau+kWGQfRqFEce2RS88d5cKVmhJQbBwXNRyp44TS512jw8qfitJ6oISP/kZ
dzZc7jQqXPuhmwJu/FP2N7XmcYIzGXYmsr0iGA4unLBReC3J4Y6cy4WPg/GkuQu0
ZASxk/Paw7gxe8+VLcTBDlCA9TwaQJ+TDSmZ3IVNvyIO3G/dWf7hzX/wlwNxZZf8
CuH81xWuPy4opPgJFJwI07cdHroYnkHqlwJTZXOwDmS+HAYU/2N2j+L7VAch6ruL
vdqzUVn/WcSn2/G17vH9/PoLN8HVG+ZFbxJK/dU6xKIDpgWym6I+7RkRzcamBLEh
EFWUoX/gbjk/AIfJw1boFbul0MmqZwxnmdD3iGnY28kwfwhwVPzXfu7no9uXWGwN
IMah9JlLutm1Uq0z1V5Cq6d3OcF68OEtVCtxpCpbMVtV7g1/Ws2wvLw5cWVN5Djo
OyQ7HkhdpMUmPJEJP9yi11oEq6Wg/K6d0kZ7HI2XN9ZJm6PVPzz/cszL9ORVTq8R
MgpqYBRLKPkoUxAzlRV2c19ttBfpM0bajrRKXGs+Ag3o0vspnfeLx5zNykZuARC9
ygo+BcpD1SsTcUy1J5kFCjEuqSbB5EzL28Y9ziytLS6DzOdWQXvKADZAiUpIm3EB
HcuGdkc7HG0l4X6LZOhOp7ZEFCVA1BnWMCzV06GOMq4r0USFfTi+Ru2aQZMkP1b/
OC2NM2JCbq5IP+ohcrfKKACC8g+Solkjh8+dY/0MA/8/N4KKXElx3lyXTbMQmCAY
55/I49hGyRX1W00n/ncHV6c0hzVYDu85li/RiiNJo+oTkTrq6EZavilGQNSbhGoc
Y9a11w+VriQkUN1LBwqmM6xMuzyTwfzZeIdh82SKFV+GmFrUl18qL1Q4dBOfeR0x
LO6E4D6QW1f3WHoCNRvpd7b1qmi7KPLHvLXjP8dG/NKAvF2hQBMB/mDqlkS3gku7
XeDdhu9/umTqc9DDFu5XqjEUp9PLN9iOG2x4ax+cYLy8e8qWVP1N2ArHDV3U6c65
TqVIZVSM5j9eHDsVSCypcuC2HpQNm+JMqtBqJrZ0SUjKM41488RvTp6YZjWeiqRT
EXT1wKHCokIX9y/jvExh80ePicwaj178c7y4nxcZJctI8iR30fbU9COSkmJABotj
zqkSfV5O9o/jsOqO3YlSEqeCuAX90Xgr+pNcJf0/FFF1hYcVt3OTMd8nl63nApJb
IS/8ealSOZBwvfDAGHQ7n+KQ0FwAEfmgkBgv6Xe3IrnuYfPwsVx45f5J6h1ePCi0
y9s0se/u3eY4DZTrJedDyjpfZLi8ht/es7+lWR6axwK/vWTLcRH4Abqq64x1JQOk
1Y200u1th4jJGsNB/wiH9SkM8SikQNpECTkD1+FPeXPqnc6Yv33rgPfB4n8m1anG
pZjwJItjmSTWne98r5me/4Eqe+TOy9hNihIuiWk0bJXuHAethaUkOP6z2TN0XDu2
CUviQ3F1OEjGcHNCZxMFerKGFyG6/2rua+tAo2jVYJbVR3fqRm3AsOViws3vcTMo
xwQc3za7W4uJiQeugqRlzKD38Qu49gsZILYYgHpCZM390aL48SbVW+F/AlRIxCOP
GxFbb5pUtR0DBmRif/XN7mVplSpTFgzqDtwYlcVCHMk29wZXHoUXZxCrZMb0Kuso
FXqj1b2e+F7A84+9nDeFVLyAQ0okLYpol4uM5NvghrRzfJdF90zmLqWAtig8FpZR
V6B967O37kRKz0dSOvw/E6qtSbH0/bIeS2LGJqdNfpm+60d88r2B1W3DBokdO6FE
/oP19mHQcNOiAn+fq0Exfyq1qe/ODHC+esxSpoJiG2QH6h+5DiW9O/LSi/jg84Ie
j4XSOkgF+o2jzaGZszF7C1FfXJIXhe9fuRMxPJKg0QSoDYJa2IdA2YGI84wyTrFA
ZsFyBCWen3M8bpIO63Weos248FoIhHSnzNqXq/R4hIWv+oVwuEL32k3TkOQt9Tj1
1kaq7wvdVC5ZaCbPx0FrQ1FrWibfPP2D9DK579vk4CXQEjaO/UzlvgeKT+/G2QQj
FXGDLutwij4RYV1J5kmtyeJUR8gzard6Uez4tqN8Q1UNju7lhCrNg83TMcM9ZtER
pnMbqxrBNVD6VdyNQJB/D+7KOCCeqa+ZklhXwV9AshHT6ZqhXkFjvnUBHtDbodR2
6QCglkR6AEhOABph8FBpDW5PBYMZl6vNCXVzVov+MLPPO/ODrSCOk4a45UDcdumY
CR9Li27OR/jfP7HPMdJ/xqY/Au2O5F/qnU8AmI2jWzhm/f7wf93UWn4Yo/8rPizJ
GjC/MhUctzqHXoeV3nn4I8oAmZsOIuRl3ffCnla2ia0LEPOfrsHarszjD/4T9Nre
Huw85AUXl5H1YR7U2UlWtrJsl4pJRioG0FONf0TnPQp/oEBhMQj4cHZ5qpUI0FvX
VYWCukqZ72BKAJTQkjB6sl1MCt+q+AzPTsApub1r/dIfzBKAy4D0ettq8ErYjU57
yW37XpqIS5U+nruYBTTAeZfh95gRWmK2XMomBiqGOmZCJog5ZuphTKT95iyYSYXd
7ipH0DyBecFibK8xqHwY5HPV/iFOefHe/bg4MDFHct1jkvxl99vTZk4XlmzM+JJA
Mck6/pcknRAgZnS5mFI9knnpoXSZI9cLACBqaGpgy4GT9TrlmIJQnQ9mkzyrwTYb
pWcUKmfnnky0BzpkukBrwttwW9AADwyva8IM9nQ1lP1QNXcEGmVuxq2aflN/dyHo
j2f4b0ux1OhguYmqJaaeZJ8laAbOpVW13741qfS/cy5rWtHn3T6TKOneCMIIQ2oK
WySz/wVkkPKLND3miyA+8x30LeauvoT1mpvmpdEwvDRsJZk0pgM8tQT2NK2iJ2k+
a5rtTiqrkMNy9ytzWsdk+2ffTf4xnjXitttvFIyV1BilAlT2OOlgV0kmtdB5bQJb
bf6l/tnTeFRAGSdZH6YKmZYPkR1wU7r3mAsNQ4Xshc6lVVc6GPooQ+ADxtP+nBTi
h7wLysSQyUAxpFCC2nsTq6l+EsP9+D2fVlz9SSXHmUATjwROHChDcer0xySWdFG4
7hkQPc8y9NPOavd4HWC0hPIquYC8IKNRJT0d1o0JlShOtxodGY+tf2UdtEZxPcxx
0ZelFS72JNADAxflmySSL3I7kxFzqG0d3iaYghwue+WsaO41zv5v3RXPMwzc+nk/
Z4HZc0noj2+99ipnFK6g9jQvavY638xmT7Ntgl1wbJHScBWwLT49+qCTPU8CM9Hd
fKqLn5nHIZ39etRfSA01bUF0wZTl3myz5+8WS3jX9Y4f3lt5pHzP07bHK7BksVqR
IKOCESEd18rgvGxEy4xUWimxA50NYTsqMQ0MYeb12kW637VptoZzoG7QXYcxGSjr
QcR8vC+YlCe+e1LiWfG61Fsjv33eX/wR+T1E6qeJtBuUSTyDay24Nzxsp6iLd/AW
hX2HqEnm57XhVo4F0VQ+QVuFsEwtHyZVBmooZMhkS8gzWrjqNt5xCaBUyyk25ViA
nLG6Uk8NJmsxkwu3b7s7m8j2B2V2iqg/aMmB8hbm3CVVFnsj5RRhXIu2DK55ikcR
OQO2WUysNAhjEkAwnVysuml9XxhyXT6MaSAoeKCvkQnoekg4rx4bhIkSVKTnSVYa
Gwu+aiB1lqq6I7B5gK+AopfcwglMEuXOmfJ2Pab409UdIL4dLeuLGk0D8/xHK4pr
VxuUbUInl7EqckywdZuYNHjUL8hIaneZPmWf7O+3M7LR3DjsAJ2mrWTG0DTOsgoR
37R5T+hf0xVqnHzpizeDeylcrgW8wC4sWGOR1VURO+/cbxE/Bhxs5HnsWjuQAfD9
LMutzV6vw38RHswe18MSk/6QH3KVCLfJXhCBrylNWgdbfzbt6CPn+R4zI7DT9hP8
RU6V98Ab5SW5fySyPgfU3bu95Ae6C/gqfv5767/9b2NtcJsS5GSgdkApZv1FwpYK
i1JuuEpaZGpniK21aeBd/f01eNzzOfTfJef4G9OZdTb5vOMugweCDBvOKmESRsW0
C4lrtjil8z6T5HNiut0A9kEonzanv7oEvkY8ZIaGOfvrsbZkZwI9LIv/go+EG2mU
QdYegNnJlAntSzIEwQ0rwLIl7ptaUDLlg/r+9QXrnJ+ssPpsO+Ypq8wO0w89FuSe
d1cBIQHTLOSA4MubgejO3SrBQWl+Zs63GXqu2An+r6V2CBbJaa+lOVkC1q5KrRBd
0G94HEu4XtbDExlzQWOk5sQsAaETgQ9MGq0fNYYaOz43Z4uVwYA+V648BKEh7Q25
//maEifUe63DwHXpRmEe/xJ+OUrJj9hPVI74ARzj+7TPZ8RQEMvGDP1QKlVpqAyw
FJT/mqZmeMqBj3GzkyXlRuliOTTVtGXk5gPdspYTflUjup9CVXzLehcTUiJ/hRcL
epOTI48JNeSavlyF1ld4IY8AEh3IBVCnk/kphNqxilLFkSp+UQ0eoaZRWE38gmyy
Ka+lZkqYiZDi/Xiqiu7AgPy+AstuBCKVjlrWEOg+9Dc2nJuWmsOZUsBfBPtvYgZT
K96eRobLXcRWNcti7GHhDRpZiMQGXaZMPlzECTY7KQTzH2QgPeV2WDMoRgmUYkh2
k+uOmNEPhGyHhhgWHAUPEzYhfigKBAEuVa1JT51dKh4KHTr/zfQhmQZYmk2wjQm4
c9mbe+hUcBAO2ayqsZy8C5mY+yNXvbSxMlQDW+cvtVOkF48OrTWJ/5obdqPRUe/I
pO9Y0dIcT/rIpnsdQkqt8+EtDWx/B3zN508rQYDM820VyeSf+02kFqVsQVjp43d8
qZNAJ85tdarQvdHm/flnWO8YIrDm6edZaryLws3NPUUjqFlAmvyYO3+ITsxzB/oJ
idM86MLq0QHJv3XvtvBJ+GG2tKT7EcPJAJHrNTAtAG/3KjRNXDwh5CkLhdH8iJjF
swCXEYEII+baVnv4eJrT9ffLojaPt2W8UDMNpt19G5XHZJgD5gaasnFbUsWEG0Cw
S8OVZsES2ZCKznPp9nhfHoni9HWE64O8oMa7ID/qVn+kc4hQAgVMq6yB2jZbSAYs
iH1uDWIQ3FKwfb5wc7YeR8voc7WC/m4VAu2u3Hj/X6+2VQk12i6QevEH21+kixE3
yOmULJk5S00R+Ub8iWXdjPBcNlpT6ouLD17cQMwypBZMRbLWVHhyRYmod83r3r8j
YNbej6DbL4v69hWqK/tppA7x/MPokfkTCakN1W+gRlPDH7rE0wU+cmWbyAier4dP
RVRhCFhx69x97LXAlF9BtX6NPHNklfR7p7q4FCqNizPKFko1N1NvOjZD6ueqdQFr
wVrDfNYdEOxvdRgDgxukYx22A5/xErTVU/ziX6WqJyoYhVvLRmfQBCMPlaVE8YZV
0MR9NC89opygeK63L93j/IM/vnWLauncswgzvOPdjrY457q9OaZtFSmLLTDRYm3z
ssE4H9+gPYprl533iz2cNtLCZWYRh/RYRGyHpdanFdQL7ME1vWvTLI5L4G1xwrmB
QZ4FtMGi2ojlgWXYF4Yk0WF1IWkWwKzoh3n99+T1taha0XRzPXOvJrjtZaIgNjVu
TWcjQcFRynTEfM7XZ5dyck7PGMgSlEnPU6Rk9pFRLP+n4Us2esnBSp8ch1Difn0V
0nLI4MkFUA+A6/PCZADuPFh5YoLsBatHM6pWSZucaZCndsDojKMCWhZUdastC+WN
IXqrXVSb84SnbhBTnCaNr7baJ6BMSs4JSIeI36HCmjjT6o4ilOBiHdARD1OuIiEg
sb/NVC5hBzof1Cafh9n/HYNcuW+FpC5ANw4RvPMS+6FLgBDn90SDWr4HpNp2ImiM
7t8+ovtIfiTUB42SmNaoILLsFqq0ztzAziWpmrHadiW5ct6VWWY4LhTWb7L+2o2f
GJ/oEFc6FC/LgTLCgypQ9AA6CCZ+p4dGAatQr+0BYLmVvjhy/CTTxhvrPP2teiVD
uMRUzd60k50hZ2XT7tWsbrDXpF+lqpmaLJCtnepd031DcVYPQ69xWa9Bb9djnfkO
Cz3UJaqnptLNWRH20kuVmQhhlN0aJRN8IGteIqywLBYj96Wkh/TPY7+y7wFPBhnh
4HobIg4CmYqdXNG7A6hHjqsaxcvwMlpo6E0tMMrVC/sWwUps+JTjg4qwrw9hWOJn
lXoSRSZWFBNyThe4pyQV55kSl9rSdBvZpnplDFa/R0MAJZPfFC01uVHr1sQD+McD
eEzXOT27w0XdjUmmjKNEzatttdMLIS+v6jhtdcRqXiiFGDI1tySWgdLC3NueJ2Sb
CnI/IYodcj9XbggA91f/BSGXSV/trRNWALO1g4oCPvqNJXg8WB299KvUJinj+lC8
hjHMfk5hAbfUOUjy1s+pOp1h7P9/i06Cl578ILMUWhPD1ZPlMpzizMbLPKGGLuXi
+J2y5f60wwCywnmSwhaA2FgH02qwDRChAqhnVpGWXz4i+0HVGkBMaHKdUpRZ8Uf5
+tsOvKevtIQFG8zJdCG3lJWdUQUJwyZ9BSmjtJzZG3NzE8LSRe7KG4PJRi8Nt24B
/FcW9R9tb9e7sdpjBD1SNCI4N6DOGxXZpVWErNdjBNLlP+V63w3xJqMZ/38UaIxM
So8wZejkPTh524gi6xnOkvNbX6hHAGG26Ro16Vv4mUJHuhKkUsUIXPeHXVxf0HWD
4oOvNAMEkmf85Pw1XkxBdm14gmk9rGwel3Bn/VLIUz3V6NqwvBrQEgbUbJx+joSK
Ker/E1CBATKWUsHgQF1k8DkYRg8/WDMtj82BCAGDtUU4zRI/kKFVPvV6tMS+R9se
bvzb0JuRiW3+ZALZ9GH4fE291BQUsOW6zZf/TcNT5pqBKeriyE49Os8blsmpvwET
EWNBUYcoL9ZH694ww56bj3fvANVyo5SetJ2XjhMdtHzcYxd7qRBMIMU5eJpmVrd3
JMMPTuCodWtFxjpL+Uf5302dLdzJnF5AmUatHJPFnfUkDN9k9ZFd9yhESSUXcrMq
pUGJbQTEKxRVA3VRfxwhp5rpDea0E/o8mTvbojhIpF2odns6qC8XETU5jabYpgQ1
mlOJV+Blm+DHOmxR1imaU0ApUpE0bfNXk0FTKMpbQPvaf7Po/cbBj4xxyD86iiIF
c6pBoi7oWftvd5O9t0mzPMYRlv1CeM65ckbVgrcgYTmvS4gpr7Oie6tGf6H0s6Pl
L4uI/3beVa5o3GtQ1wZo9KKiogd1axjkLkHXiSUNgVEBK6rsCfAy49QrE1J86y3s
ukzIw+z7LBy5T0iAoZStsKwJFF031V9Qx1zQtOpR/NUyFQchsdEbiUS7CmTMh0JF
1EFljIVg6CkG7lW9Pqx0Ksge0GyDhSQHvl9t0XvEHxV5MN3LZO4/0q7OnyZ0SQay
H9RyUbDAEh7xjKuf/NWNsI2n6DXA3VynXyRaR4OfzF2dGdNfK6GRO+DtHd5jIRt+
MpUecI0GXogTubAr+9/KxQBUMjLuRaQNwdOrXSmpz6Du7gdBoyJ+nj0K5hvvcCwu
oiCp3FPK5W60fRhTR8tPP92jpcgKKr6baAGao4yjPU8/B7xgaJhhyQ15OxB5tEaX
ZlE3YXWCM7cRj+GRCAcZ6if2xT6zI01xuDnSNzx5cu9ULLwwVpRZJcgKiRJ5xEcC
Sm86GacPW02xpngImbqWp/ENQ3/qiRUza3Hb08PegGf4DRdbdLDNnDerOvtqHUoL
Goay4u1hbTHQ9ZThoyhTdM4jf5LAnijCRuHzabmMMY3JFBXmP2new4ZsMMzDUlyi
8MoXOgsmksexOcKhu4XWHWcPwf0Hi+jfKleLT063StzPTgIvCu4XSgK0dXsEG364
bu/twh5GYatBsl8v0ILCvzmxq7UbX8Xc1h3XVpapearYC+9kzU7meVudQZ2Ei+oQ
Xn0I08BBQr/h3Z4h3i4DGS1Je9d5EQklwYVdrVpAL79XG2xXaXDD0GgeQv79QKoC
CWvBn331z38ONCRldhHKi/rM5+OMljBH4iIBa5UNLUK5yjh4gGiMPFN/3R5h5REp
DkCWldDOVr30l4l5F3daH8wIybGiJ8+wiAdQpW66KyuKVr9JNpqPqih1A04g2gPL
6I1dSWnWtg9iQMFVGx+ktauhQTw0VUf5MGczZ5CmceCr4EIqvhCucFoExJUHtI7q
XZpE3kOHT25kGj2HVoHCSNRxFr5X9rpIGGLWnA6Ek6lhnnMi8YIh6pEZlIqIMsKi
cFNssacFSdSbpQAZJ5dxhIvaEjZNCU9pxPuL/oa66WP+p36sYbxbXJsC1PoVZYdC
y+/nxISYrxvd5KQtARX6JyFUm51MApPMwzADtIb5+06gk7lesNXqgZzOfHC9uhCT
NkDq3BiagIJoLu2dbYOM0A2k7mDbNNcYe+DEVjZrHImcPsDG68gd/bTDurrg9Udv
llMXJjmL74cL/6r5R7NoY25spkiaiXutYXGPb6dwok3Ab3gasmToq1PiK61uJwRT
cYRDJKPCcfQgo86wi+Dr7z4qP+kg4+aCmLET4PVZFS9frrhHLdvWtE1m635tNN8p
fqIDdo8Y/Jx7f77B30EixxO0W42OuY3Un2LM3NWh/lUzy5Cu5G+TSlHDrQcnfDTq
nz/rCRXKbPQJl5onDElKFhox0xIjOzmDEmL5BGfK8EYuGsgM7N0is1ZllQ6ZIbhf
48d8GQs6bR6TMSPwAQ3WOH48WncsqlaZ2TlQZKHTue4dUFcn79JvD2V5+ioIsily
/jKHJu1mqn6ydAZyrCuJD1sq90VfUcZd4cIy0BRORlXa2dh/lPLqd0yTetOvkAsC
qM/5GXstSWnFL5i5xhckCWOIw0tr+dI41C7l+xEkEfk+tRpBZ1geaeUqmwD5hbEl
xrVXglypmiNA8Z1zAMuHqPTvbjmkmP6lAlzhlBC4XLfSBbwvi7+P1FVX/kVw8voP
zpA6iPyX/EY/NPL7zANNQe09ucxf+U/QPwuJZU7XKlxWiPR4RGGHye7hm2w5qIHH
ysXLKkrMGJK8lcDF8ufiHPKQZPBm9mm/KCrv7/DkhQc2sA3zX79l0JTvxFuQ8WW4
bfw/pQqlaIIdPsE3GNVXR0QA2GPZabi7j3YVzZ0IjdeLEYIGFcg3uwiGJ6zpqOQR
i8Pzcdc5JJWumYKxPzGB5blGGEu33Gt+uAXL/vx9sqIYePV/vNMjX+43RbX16PlX
mUiZDw+uBuLgCvOyCmklW8QlbXJRgb+5NW7Kz4+xEc6sJHvF6rChcXyUisYZGixM
AnHgzhgIPNObOYjU1tDzMn8aSt5GMaH1LLkgN/Lkkx+YFzBiTjPd25yB3n9891P0
L/oDJWC2oYQXnxOWuPSKOkqvU1D8MwmHB8GyYqmRO3ULOZXHVsIsPBXz3nEWIhhn
1C3DdH5sZkbhK+SDlzxYIC/EAD/7dedw7R6jW9N2lLkb2Al8V123VDvM8YaH5U7x
sB9Qtxp+RZwKloXU+jrSY9NR9eCcVPOKD2taoMfCbVvdgxNlTs/GliDaGEjYM04n
2NlQBNc1VduxLEAU9z1ptFzxTdOtZ72CIYyMc5Vhq8+w0JO2qpvVp48dXLadI+sK
vZFZtEBYmJBnsGJ80M3jtV8IiidCCxgL3zGwnWhtKlKcEcxHABItxnL7iJfvZ5Xx
dL+QhciaOlwbGzABEn0Y9h8jnsq1O3tTLa0wpudtOsDA7OnojBwJp7N2icuqKzm/
jK8qPzQY1y/E01eV7gb9Je1IK058CYNch35n/nXlqicHTfpwOCrCWSk/EhjwI3dV
zxN3AV6g3x/+LFb26pb9dc5A98o+BaHpuSaive+OnjnFsz/iNF6BJv5tRAx205Bz
w0bx+f0I/+fCz+jXLW8UPOO8+faeUBDS8RyCxa8tIDPnFlp9A82/yFSPGG/63lIl
fdB7EWcblv/pQ10uyTWt5HmrUoiyhdPAKNSaFzc9Supgkn3vh6y9zDQlV4tYVxUA
pvyqraPgTbPmfmv/8exmwDdP10dr18C5T2hvbDQcYejg5w3saZ8VEpZd9h7+sbtF
ypvXmDDoVm4pBgMQNrijKl6jUo8tB/TsDJfUKYMu9xvqcDRevKsMi3upoya1maVg
0+3iojw2KT/zEe7w27eotYqtk7K1UJ5l+nzI3c1levXyq8hukTxleTj90pxE205u
H7tYRRqmn1e9m537yD+jdZFZLDvta9o9RhaIrUlSno9mmpf3qApXgfDNLSm/5GMk
RMju06wnMAMETRhCzNq0TDckaZhPeG8Ey32NApN3n1rWdKfVyTTpjox7uTQYaZM9
UUFL8o+YNADMZHPDbDSLI3RxeeefEA1OSHPB98D7FxXPmDeAYNQWAGhfiHJeZTIX
YdXepxdy5mseUyBhxWnct1VBBOwE+5LzHL22pPML+pDWLPB5JiTlggyqXJ7dtBhs
hCZyoJ4AfYmqaFzfXCzqRbPWo0W/7cLC3dgtUgmv5XWElYuAu5jrgxhBY7XAff+A
YXmBv2uqt7OjRJEVe+DPkJEl0EXTzxsNf/A2Tt6cIdB2b9ejDhv+wmdpOF41BHVH
rP1/fANcAaNfsHWUQ8hSecDDv+I7L32E8HOuyDfVfX7QHzkIxGiqq/mvqKO9Dgm3
YD/DwpExAgGx6/7+mVG7e9m0h4Gd4iOFo/HLLYNNwZ+Jvnr++Bi8N40VTlCEyPsW
dsPE5J8byDk+Xn5jySRiDwmS6Ef6hMbnLoaHFnXYDDDVvUqpiFIAsUIkxi2XxJpn
8cnlsaZBQ5ken+handTjpWgfy2Qn4oGR+Ks+h/b7fAzFQkXpd9c7NP/ZGJz4woXS
XuJfAJIWBubeseVAD1AvC89aGnQIOX2+mOeBm9oxPrJx8qaMXHUYya0wTosV6cTo
obzmp9fWaPyN+vdeMWLCFo+LHHyWHVQkfPr6Hce3rdgXAed/s+kEmxTuN30Kzhzx
Y/IAgbZreNiW/87SFx+sXWleB5WM1WC+LKITgV5AgANVdU7VktQ9wC5JO+SeFssl
GF4oboOrWdpS9NMdjgUj+8fjzKEE4OWQV88DUTwccGI2+uNMjc3Hdq+GGmMKVzTG
I43Om19u2cPb0Kwdt3Rq1diuKbNUZWMqbHQ1Pn6avW3i/BC8W7HD+o5+e/wc8bm9
avYmajAsZpYYdZ3fX+tLiDkBCIqXO9ao/HtBw4PiYKoEoMmCoVLpIO/Ey8ZdOips
y2p/UeTaTwGHNH3hjiGRuR06aYWT0U2sT8UEPCa2LOzMc4/eYOgkw4vhDTNx+CH5
qPsvLaaj8p0uemKvdr5EK2dpwE5+scGm8HLbpYjavLc8GBVzgdlwUt8yWy6733AX
EbzmWniXrP4cIrq301JxqbXk6XVZHlHeuKmY4RPHXKjHm/ArmUCWBVMzhzVwmlhs
PF30Q85L8bNjanAkJsursGBfThpLX3d0co0OZT4iZORT7M9TEfITw6t1bblkUOp/
lxErtIpdq6Q5o9ssOaVIqcvzJErDgyQiMrArpmaTIlMuhOqwJ8agTKs5uY/r/sae
ryXe0/DzDN0mIk2TzKmnoUIkQZtBYgFEyWt9SfrVfRQ19dHlJSzzFTuAj5rdXOb+
HtNR+WfIz/nyTbJBnRV23V6JuWOGYVi9tfd64+Wk7CbUmBLYYaNNSBfD1OO1gH+x
gO7ENvvLSBBqPy1qI8VdLLBjY3/lOuGvxePIZ6USJ+dxW5AWKqPxNz0gq9/gJZOn
OEAH2dnJzhaSAfdbQqU4e0zOxg3hKZGcV1DQDbQF7H2gR5s9DXwpRsG0fdpGBopa
QIPPlJ3yeqDhdHqMhOVxSLAL3ueQpkfoatQYC0r9DL0LMXzFvZOscBlHgQm3+6As
1la9BJjf9smwUzPYp/b7Om9fE5S04I2rozRzQOoxhIhZNHL5ohNiyTc7xyDEdtdu
ym5S+2UgjQDnP97YADhg8rj5B9kLLN4O+oUQGhU0ZtXCAEVwxof2xg0LWQLY1O3M
EKbWHh5kM+Os7u+WcCvaQh+Jlo3hpwFzoDIXybneoXfhVGggNIh4jXtP8iW+00tX
8FBWvDQwh+dWrEI9PytywokU/es5UyZNEk1BgHkip79pb9q8sYNGsdWVGWLcO2o/
/QIXDND4kt/dcBpI/qbQGdyGshM6TcyCOAXd0vJPnkJL9v0Ud0Z6h3ZPaubDxXsn
5VviNpoCujS5cL3pUGSUslfQHfIcya/CZPojafyZ+ULz13heFEjThpMmtWZ80Srz
Tao3C97/qELO/uMEiOG+UOFj9NKIbJBkmrzsuxJn7H9Czc4L8fKyQpfZNGlE+BTc
N2fEJioh3xE9TsUAfC+HE6YLFwSg9ueqT/fIoYK+mXm+y9qw3vW856+cpc4Otzde
sRek4yzxppS2SNtVLLYdGpcsS4h0zrjbsLaCS1NveSWAgzgpx13ZWm+ZnZE33key
30ASp6KLbzL0Z7u+FnOPq0kJuh6mMgzai2BN9zE25Kq8TY1/arFoQb9xwFvvJKdk
hdiprSZZdvwSIbogl6xCGJJAysbAv+3mWBXSucfCFtzPRxP5p3e6hecTGUDBFcEl
ZeD7QRQQjO2joM+c74kOSbzCLEir3+Cix8AtCM4Sh9BDTE+aSddWVv7/rIB98Byf
2vtemMAzAjjIysHs3+5EWJW7TU6J9qLCvc2rHVHm+Sv5zLq4Cssx75p+OOD5/pzP
/1q4ntsXOFeBBWpNXdi5oq8QebRLsOKTMcl0W70amUx9WJdmvxG9PEeGd5awquIo
EgTSQPtftmUudQsEFAdT1LY3NIbFn7ALj/Z0L64gtboEbwZaYa54bEXdzBKgH3wZ
IWZ8rljRqNfyX7XvYTS7qku+5SbJVunawoabQQ4CfVsszO4Qb/4DupCo8TC4whLT
zdOqX+D+ShmQzqpPIji15zGq/t3Pd7te17hXGJZ56Oz0/cJ1G5geBMRAzl26hhCI
9HpVsFzB1zPQtwqwnu/TiJQm3e69isHFbI09lE2mRLtGy96PqD/iSNx5GkHYl52l
AW7s6FZ5dEOKIK4qhIQHuLELTsgI0Ih86BWOOKrwPdL8W/kQmMZRY588TGSpOP5t
0mHMMZ4jaCmV0NMb7yB9+245LKmFXS93sb6IC8YkoXyWzkVZte/Zd77acfbCSRRO
4zT3nHRIfg/n0WW8Mktg0YvjwNiXQ0l8MN3C3eMZH9eQxD+ZsWXcP7zk/OwuKfrq
h3xrOUesNE40kwheEz3lB7VizTP7iBMkseJzJUNVHowZ0Qlu0HoQc3p3qkPI5usG
yUUr5PgQ+kxRog66pPIGbF9bfXJT6C3lbRo/7vPs8OSZYl1WnB5WqqGgSl5nGqAP
GCXJlUgi74eRbt7FrLKq68SXpu1UiAtL8I7Qw/qfZ4KtyjHZuozsZqV5+QEdGyDc
czm4qeqAX9kWwDS8aJYMAdAOv0w2o5CLy36Pg+7U6aZ2N9G4mEOXmj4miv4gFTAF
uXjoHRDooyfRl5vBFOqI9uW1+nQzqJp9s/CIVob7OMBeVvTZCLS1dVMajnX19+6S
/wpA4ENW8hOLJLA54sTRhNs9TWUWYhIU4hZB1vPxsQdjDbp+ordrqrSDzEjkPMMG
HcNGsVL3rNbGcqYjl07bEeq/OVGd8VtcIKg6P5J4mKwO7BIcWoAZvNFfLH1qezGG
nDAl1o8jekprIfbQ2F2LeGkXPU8KklLgICU/i3i/u2CVRqOnlH7GFsoKUstBc/YT
YJ4Xj2xp4Rqb87JftbM5tPrKbzooMkbVKA7YS0FU7zLzBG++6LN6tNkP/BOZBav5
kzQfo+/UFJvfx0YFiXt2wK3u/LKcEGjStcgN3FXl0/5tcIt87jNOr0Et+yCxnoLt
HBCHLezCx4MoeNuWtS6U+M9Wt6UzcFUBmRzEDuRQA8zXZychOkln/Yo50jAJPntN
kuT/uPCrOni+oy0KIEXy597HEoq7PvwF+VbBJOXwiMujvm5FagQqqtT0h3l6P58G
+z/sKwMkpECUr5oBTAWD3kd7XnXqo0RP2I0ZPXkJpj8rujl08lQtMYXeH2xBqA5E
1zS82tdNhdgvl0ucaW1LQ35lYzMBgulQlLUolrOsv9B/emk7bZbVoIczSxXwZgqv
/bAudpvZZYr8miua4CIHIP8dP35CsUSLVySUHxF+O0JsvPYphHLMwkRAyb8Zmsmc
hfWAza5FKADzIVmI0GYj+GhIrVNPYGOqpCAYrMR57V/uTXRzJx4wrLN708e1OIB5
sKJzEqedtCpHLlmpfIIvOIamCih7L/YdL4M5dWpO7XHkeXvDH2mr7PrZeaUWJ9Ai
6KxyGG8IK+KcYxZByQ78/ita0HOKdxR3egeoxXHmrWiNupCZ1irEDew6fhiKGoWT
YTe7NimGnZAOlGtlZX3q2y3lN7tRFRj1Vc14B6cxT2seHqpJ8BsANiVF9MKikFqs
rL+bdbyl1wwICUuXYO8W0T7x8Il9ZeUnkMU/JqKqZZaYmNgjujnnXb/ktYzNQvCs
ptc8U5GENcAEQpHjdGS4/U2AuJxGpKyH/hFeqdJ1BoPRBc9czzFRQghvqJUpOy2V
c3F/bBs8wOuclxki+mHo/+o1GOYyPbqoH9NQGT1L/+ocCli52PavtiLlKcvLdNy8
R/nGpz2hdj8lzvuzXFeuvZaLQisxWXY04wTJr7UD78J5esaSqdHnvH4Rc5cjsyrl
IwmVU6WTU6nirRqBo2d9fKlIAX/qGJTuKRGOg0MDOVPyKUIL0r9Ao+2k0fMR84ny
ksAax69m5HjIGAkhNlw7yFtTLMgurn+12flYyc/OzKT1HEnLXMXodRuw8/qlRQun
PcT0nrKrCk5Zoh51P6T+xEyCHNrzBL5LMlycCvdOkxkfvEC9+yOt59jMkAePTpG3
nans0DESukIJ5Vsbamx9cWzL2ezw9f8nkzZvVWt3OIMNndPKe1hZvUv8r1zc6NnJ
X1H8vhsjDoHk/T8E9sTSevzEblVzVo00uO+/hqBroOtoewOorSJ90vxD63Bl1lFR
TNt1WPcwvJZkFSrXQnEN3ic9h3vhXmLj1SY4uAiemFalU5PDi66x5oCckr67hXjG
7unvKhA7CQ1h6hXaacV6iqUmV3lGVFvHc38dh+1ua0bYvd2sKJNoTIfoffIS7IdG
j13b4J8/WZ3UhmmWdCG7+urtGi9Vb8wD0uYxcjHyTvCrO2t3oboaLb8EFw7DoCNz
OVJE3ENNmwY+qNHY45O87QmRcxusl0QSnLWfs4eXyEU/XMkLz7WHrms3VhJNXots
e2im8IS6lP2r7zRKXtaMpQ2iSO8m6oFGXIwv5bGTaOzCmtDxUisJHLamPoySi46p
7923j2GSIQ1rNJyFkS30quxRM8/kUS3ddEecUz49v/r3qQ2kgrAl7vJJqr8XOgoy
zX5bI4D79RZL7+b+2og8v7mLDA2V5/y9jYp8hlmD/HWMjl1yd708tv14blDt6nmj
yBx6nkbWpRSPjWACm0eYTxhv2cmEAj6lfxMeI4Khm010n/DqlkjqA1vhZmurkgpt
a2scJ7/cT4gimY2ZTT1DJdhWxmh9+am2Pc54dflIWBgBupkhy1z+TFKc+pJ0lqcS
PUp9iW09c7/ILnC/3Zm12pt9O38x4WHw4VbIDsGIPytG76FILYbsbYSKHBQ6ufMK
aTXrMoJtAXUuFDQ80GRd/SVvz2Kh+8EcpJpTrKTLZ64xoKanF3WCLqy5P1lo0MK7
A4KnhDIwF0uZCLDTL3p/H+Y6jbHxlURX85+rxeaRMGXfg7dp1NXXs9lkNYMv64ur
PDj1sQ5H4pKQVmS1WTtoiltW+Kf4L0ojBjO9A8y7ulrqY3oV006Jm2YcU1HX8mk9
eM/K2gM5Hi9M1CPknHSyzeNHO9GIivZxb2pYBBz2Z+Ycc07Mp/CKv4QMK5fAYzUm
HxPvPhmbleewAOLjfMyPWo6uHXw6QeOjq65jdJj+aZd+RGlPdZ4E6eqZmXH1lJP5
c7Ll1CrUSliO46OBnwC2kCQ6TILcwUBSR/vjv6ZpABCHmfYLBFKg8ozhnRii8QeM
CJPag6k37Mmrz5thuiqwKgtnZTROdfWSWzeSM3Z15HoW+V9FBti+Q8qZtEmOjJ4z
CJMG3hcHEmMz5meEz4Kx5Qld8pn3z8oesHXAX9JOnXeY2btL0kFSWdswtcOf1yjy
qRGiACXblhUOBAJYQgBXktr+48nIBBFjaxVInwz1ZIgECblPHLyEqOkJWp/zpVs4
JF/XT+vWIbHmdPoZ3vKEeLCMoXD1Gp4DoEH10+TYC/N/gzWd+3gDm8prghSuZdKO
feeLtVGwYa/Ev0kpE9xiIy7iYK/n62TUfrFP7ZbRos2UQj4fGLJtkszMygOPzBdG
wiJuhMfqyBaHxQQcjOOvP9hJKkIGhBVKKlZVjnCa4r+x7AQG2Ln+2Hko9opYYRB3
Cz6vx9qWgiNGmuWm2y/S031LfD9Y+Y01E4/qcIBXL0abcTOCLgty5gsapUC4crVY
JsMU1vc35SeCjqO+sdPENQMj1/F54DV9ZJyAf4SasYz/ABCKhKXEW0gW29RUFcuJ
ve6UXDfbn66b+LSip9zCuil0a9XRKpCKe+KbOR6enbf4lA3BF2kjIW+Q4J4yzNWg
T8GvLcWytqTizTFP4WcNaV11I5AmlWrj8DwES/u4U3vMaI8vqZTiQhGXsO+clIki
puIZM7WSMghA6ZtCKgcwMRz19Z9/bkyqPbGj7VJeoHMXJEJbF1wvmZxuCrfGYMxi
tLlw1fftFeH4QuEwM2Jn/Hw9mPg0+S6TU0BeeD9aDkn/PpOhVU14xUHTx1Kx/Vth
jlBKhHKdjjxdeT3SykvhzxnCCHaCyVObnMLJojNDfDPTcog6bzaShexbRB/7MmY5
xiW9NJCNU53Ul9ja4sMUjr6cjCYOPx5fZtB87G3Nz8JRMLN6QGGvudBWt7+mFMB4
8OhJYb43AOa356wJjvw99jrIVofJ//tx1xAx0mIKhSOdOkSPKLtBJ6L8TGJ7d9cK
WHKiuozFXijJXJHbya2/R4lSZN4FY4WboMbq2Y1RY4qTiJWwMwuOFP3LSmiXNN30
bHOz0onWC7KLZ2u3yV+wEZ4Q+lylO44B0cShWhrLw26W65OVKuvPTPcmEbvhMYH0
bCQY/Y0ODV4Frb9gfTH1I9Zt9mJ43u8zw9ORd7m+YPvHo/uosEx+7Vhm51P9S0Qx
EgD+4cZjeQt7/0t2kAoYExVjlpplMwQbOGanWIxvWW2AoV/KuCZpZXKxt44mPH0g
Hhp6miFQYw5nvxClF0gWaVLPdzL8Db5dqhEhYHL+oavmwj6bTgS8hLrqyX7M0wtN
5hm8C6PnX/AD6d6jwzJwQcHo9p/Q5+nnfzFOmjc43PGtwhtOEgSP8vghKPE5rFUi
CIe12eddOSymbx7if9Uq72WpXb3DfOuq8Pj/UjEaNb3RTIs2r/ecYnd8PmA8UnNh
r7Za5vizz8jUe4SBR2Prb+wb1fSXVaSlPy7DfAMIneb58b7y4Se730vR5NFWxS2b
s84ZzihnP36ku4t+t4xRvumM/wobZAMm0tQVu6gvUR5uYNPTTMt1RB0HFg/BxeiL
56NHzn9zd07j7BZ0OfK6Pa/AwUv4fK+1IizHTQblBIaIY6ZbsF7Mt3usqc3b5qiK
vJpq8nLA6uU/crkxG/DaITRvF3uMFm/BVoOMpf5VOp+uwVez7it2dazMyGpLzem1
LqKzTODWp0s9xz17ax5f8bTzr3TKiH9Rt8Nip9aSENPoIYhqhMC0BtjuDMlx8ypg
45dSsv82Gth6tlaOjIrqMwhZyckQSTieoYZry0vjiNEj1Dl2zS6Y6rE13UM47Iyr
yTiBpPjidOega89egmTNvbdxj94vYsW6skh8Y1jCxujM6unGB/AcR9BEq0QGIk+z
Ikr2sv4e+kqivrqFn9pI3ttTgyDfrHQI65gWdjfLO9S/kyaSCa2rTgLHVd06TtL1
syB2pzKeUyfcRI8EA7D/Uhn6R/Hg/iuWUxeUsmEGXn5Xj5JKR7JWGjiH3g9YM2nY
6NBD5pvIeQkQ3GgF6/4mn9BG/Yfr9QZoEDRKMN1ebESbOx1/pSynaM/qcHxca1Fi
Nt84GzaUdln127EZAqA3dDfBvswJmmcR3dxhQYiyp8acTsN482RhuD6b69TrpJyH
tM+Ys8bUo1FfSpc2XjrczsTAqMTq/Zq5Q7oCqnQlnBMLKeXAVux8xvN0pGj7/dMc
9EVzUJGpU5SF8K0K9IwI7ARZ7mTulEMw6TtEgPZIYHJgzu4KPOhuW9UHnApu2Gdj
R6iYc5onwL4VO7xaSNKoWOWIynf3Tz3ZmicviRX1kZw=
`protect END_PROTECTED
