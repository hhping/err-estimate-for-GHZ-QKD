`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/dxaUVlf3egqYJgKJ1IQiimeGfWnopVUkaxNOK8WHqnuCJlwrdNWPIviZ4W0Z5Y
QhnpvUAWbU+TcP7/TAnx1Q23VURoI+4Tvo9/qfl8yjcdZWJlqvCb/oe6rrQ+m4Ye
vaXsFHh6pufyi9WBJBFbTkebS3Cs/otB+3Kl6eYhHj5HhyRcB3OzfdUtkB6BTI/v
HtK6gqu8u4R68ksA1Yp0HX1Xuu2eS/pC27OLX1OX2rewqd5baaag4HuDPALyB4qt
6XVVx7wAZcne/4CstOvIJbjIq8q8yEBBN0I7fttuhkoK6fDxoCMk65TofRUejRa8
L20YsZ3FFU0VSok56rlcME4wNbfqJwpxYsD0gdsVwBykRr7li9zRqeQdPWAj1CX7
SJDH+PMhWQwAXNe4WmEGYcxxglpqcHXM5Ojk9x3iTlhqE5oEeoNgkD35q5fgu876
F/ksAFwAxAIcmPK0KThoOenydaMjst6HLWWwn55+2ZcsZye+d4HUCYa79Hbjhb98
uhhhKkJvMkYnZY18aCFFe9GfC9lsuv+Z1dCLXXu4JfD3SXP1DpGzCt5PFPTacRCf
36Sv7s0aTnkp9kyj+1i+rY5lWu/tJFyV6PYIYQmJI7O2Tf7RVvwkEjZvwM9Bmok0
RsnYFEv7aOZhWuKIHbeaomQKN0mD1XGvM4Muc2tUECJWCz62w+MzZ5u9edyQ5yru
pBKspfDpgjwmkK0Fv47UrkN/y6VaTowv55ghbokNudZ4B9X5FgVPh/c5P5KiZiNo
FDl8ToAsh+4tJrKdKfEXQw6M65waliEFTAKdyc4+haBdTYVjv3uSZdQAZ24n+Owi
a9GfrPW41JcpBaBEPTSL//Bs33+U8kIMu/Nf9pI4dlnDn/GSAlusb1HWEFKaUaeF
RoBV48YU4h9Vjn+FEU+uKAxGTXFHrnRlEZoFp3N5D0o6iEYnuYygGFUBsA9ImI4j
u0MmMK/SMuaQBJrp+T53aHSFHSvLGXm3pkhqXdRs0LYKjEketPOfDkB6g0H2oSIq
W3VUHFRoZANqNJZdu8C0zyHPWoEqa49E2tX6J/y0ND100NPW8M49AfpJ0Jv9Qr+b
gEmXtRf/eEx6nqHIjHR2tDuM1e+yEatv9fB/EGTLrrVosWdnWU0XooNETwbiogNO
t/b/ZwNX6PdxDZTRWb3h1FYDnzBoZhpFOfO6yPOIKui0tJ5u4i7+Oo7XgDVtuP8b
t7tmauxyo24yDZbP36MSdF+ZHsGxAJNA+Lxj57h1zWvo487rUjQiUwY+Meu2Nraf
/cQbmu4b01asozgWJ/YDnevRlYXkDlpSlnTmSF2aQsQvQhzDIUFoqSLsVKgDT8Eh
uMSD5E93QcCGZcTF6ARIGYp3zR0q1doxieud1O7KhPlEFZ7lzxpcoiIQHre/nC/K
uD7crAk7kk66RelAOPD2EiFCCZa7fURDbfdJ6/zuthasxFW80aB5wGSFHatPijBn
clTM/VvbGW6WP5UpZ8yvd7lG5dSxCcfuLzoubzFyX6zu7TCXKrij3ryWZBF5EMOI
sWyymlHQsze7jWNzbklJwnrvFU/CxgZD0A+qaL47trldnhezON/aCP+2KToSo4IG
0qYWp3Qc1IWmmcTkFPIZQZlSPKhCJ4PFPrQZqsZlhoD8ku2QfsveNVQdejrbCBPV
GhwPgHXPmqrn8xv8ap5rgz2mROkSo3jzPrAwMrjFoBXDbiVKN/OaoZA4VdI/7Vzd
cZmZM4cPaKqcnWzGcHrL2BQyz1pvd1f01npa7wbQ5JcbtmXoLq0KQI99yqy6rhOo
LodkXoIzGysAOBf4FpKzatwEGxixXdHRWxnU3Ppm+1J8NZ07BEepGPioceOB5h0C
LSS0OfrwxVNcmWAQFGj1Sgjfpudvl3V4hT2huSFQtw5r6I2tPmozM+S5oAKexsVx
Dc82WgE7UBg4hX/18OD+mMkUhHA1L10+Kq0YxZ24pCkVon2yNT/RcpOBstZDjQf/
e+jmP6fxfA1wG9kkMuHrxTInf5uNJRKQe1xSgy28LGUs4LH4j2XRTxnwNaBN2Rdz
F56Ugb29ZWJxsiVyNgz65IKNiL5PChiQRV8fmQRIx0m1avQM4aZe9tvz+t/TwvIr
0tFGB+l1YInrioIWE3shoHmJoX7Oqngpbo99C/Cua7BkuJbCEgDsDYEOrdRUZwIW
AhR4OZL7PrLBltjEpVSUKT6mB7OsBSa7ofUZH/Qxube870WLfMr6jMy13j3wHyvr
KqKevmQCf+Jrx29F4f6KNVNgErVPH54CINOw6LvsRYPHF1HRwv50MtXumK7+arle
+zaGlROFCgQ9tXTMgev40dyNGV3NCo9x5O06wwLPz+k9X8b2KRTL1QwLnaNyYtq2
JmIOi0Egjwbk7H8tsbCSOoPLN8L8TLqj8Tl7abKCRW+xBGSobaic2Na+OCiaRC43
dfjENSJI7e/lBzz6dnlKI18Vs06WpmqWGlSRFXLXpzUeYVTxYtOn4MoIGDRFXNr7
jotUm5wVSmEOALGg8NV0fB1xJedmLIE0I87lSG6FRwWKLz4htiTxCfBZQajpSyDI
srBGnGB2w4xAf3qmZWf8BFOZfV3c8xwZ0AuLF+ZBboiXsNB106mWltQ368dDycP4
frAfnBNQVxye8AFp8P0kNLMxU6l7DLH+AMxBFrDEMqV4ZFX4PTD8RLJguS2A1xHo
DYpNr2SpsResSEZWcbzNCmC/Ep5nLskCX2peQdsTdzNDgf8Vu8KxQ3sxWMpjO9w0
5oAnYGABDflHQ1eSi38VIXy+5qga1Hq/Id1mhudHlTqNEz9w4GguNO0ZG8faSE9j
aAeFe6LLlFo4PuKbojJHdGCG1kEo8QjPyoS+XJVU9aX/UQlf2+34++/+rwvGybff
4HRjFJWJqmd5UE9y/T2QVQrQRpl92in+yIPN2FrMJnP3qLH68QS+7Ji9AHNTmOVd
sAEdRXKwKJN2tMJ2+sdbgmy0+1NNfXmhvbPwqDMgbXdVkATAYNnOMHMTP5QHyml0
nx1vDQ9clxYyVrmAUgNFbgCJxq13ZIVqtm7gVfwmcfRytfM8wDYCineLPiaVkbM7
RrnF48aM835N58rPwdh1ruaJNsC6GncDLRJ3bZg3faJX/qoS0lnxqbbyFw4LBe5D
5/2ypL0j0F+FTpj5Fm5LUt43R2IONPYq4qcjtm5N22ikZBMDdgYn5LlvbAWFI7jj
mwCsHvZ0ncRC7HIyaGW2PPCWIiVJeoatrRLPRLe5VWepcJ0CEgSXfyoZlUM8Hx5N
wgv4YpXc82WrOJuQOsDDYGlJFperk07zqNP/WIuns0okp7YQPq9CAQrC81aJH/L5
/GRr4asmN/ipA23VdoERA6Jm82AkW6ngei9xcIc9Ez2nvG0tbb7Jj3PkxqZoS9pr
gAJDTKAuZeSZ+NF7trDjODRwWI1mKk8xjyOJIeegeBzmawk02jl71PWvedjptUNu
acmphfGMWhreHUEm30SQQA+yn8QDpuUELLvs7CDzd9+/IgvBZG9ngV/wD6dSL915
KDWzowrQKhCLJp4iwR455ojuZBIqLvaPeswOamgcdW8NU6HuPIvNoitbIll+WvH8
0Qr5aclHYvt3ZWiUe3yfVAOq6QRoHW/9eJIW+V7uPFAoW8pPcJ4Q0vmXM1foc60V
mR9n3/H6y9CCoz9otjIWFUGjtwjh2d4Hc19ASj0cUGn/jmWEXD/H+cVPoAQE0HDZ
Evbo+J7tRPiWWJV+G9Y1U851zPNJrq7eWMYfuvwSGN223ZK+cfsgr/+C4IO8KDMH
Jv3NK1j9V7bSW8dOGBLUPonyvYflpragR9Ce/GNQLCg6WzSUlJcPzyZM22dy82JS
knU+s3g+MKg5cCJur19sELWQzcrtpnn6wUCM8QXyplz5l+zjZs4QmIllBxU0GQiv
+zOBmU31rdmt9/twUf/bJrU5fUyRJGpREvg6HMJ5DFLi4EzkgTlkofpLXRiybmsM
p2ahByUkCQqt9Gx8wGYFFGykvRpxU+LDD/VyAnMzIDEAd2i8t33Xq/ALYV3UxuuD
F7LD+Fm4GfELu1s1ijReMKxU01IOINEAjxmjAN47CTCUFvH/nV/crNoIhAluEEz+
Ku6jziYJDfeOCi+kLUxjramBEdCsJ5Q540VsbDihcgBNZ8Ztd82S/y6oUvXXLDur
2CkuAjWBvZbZr0/BLbN3TMP5uObMPY1SteOtBgdd8PzdLmRKFGjs2Q8ugr5ZwTeW
BLEzK4KBClYpvxZ7jdAF6mRCKqQz8bPPNAOMEr22H8jKuRKlmB8otNV4Rfrya5Op
jevmjnXvuQYhxsbE6x2O7KFujZkOMF73EBwdrKRWYg1WE5bAp6yTaLrkic1hY7+S
GFEsn++492n+tHYeUtx17h+DLI9+ofvwRCN+t0VK+I4s6Xou5ryjXXr+JH8+0Vp2
C3dl6K5ubtyneh14NYQdf1XiWwLoVsS06d6ULee/hkJ08ISL9K/Qt8jenKGl15di
YHIOcaPIkLV8bN+BMI51RSF61+ppdRD9BD8KnV7/Sr6LZIqyzqh1AoKKfEFYU3B3
+fhO8JNafJrC8+GPsgT0O5m3vRhS46MVceveQKTKwlTahv4MRIhAtPfnxVoR+n/7
0rcESTJKYw8BsDAF/UQa7l+Z8A7uL73w5pqAejmIvByWFAGiUi/BTrmfcpi/2TB+
LLMdkxp0Iuzmb6K8cQntUfZvjAfBcAvrV07OdDPw2VlPXObSlTmGkDWoV3qo3RfC
Ud8BEiTNCVMo1JHBf7115wqlIrerCqwa8+144hDXpTbm1/Qu1Vf0BuEAGxkWMa9y
TlDUig5vXGKysHpD1hl99llh09ss3v3XrvSXbDEdcmWMNUp/V7ZEwURwECQe18ua
b9PQS09Y1eZM5iQ6phXy2Ktl2myB9/FNVMGTFarTZOPVmD4StUyX/RVA2rZpaR+y
mMjxqBwywj30leqT6UQ146f/glTo/wQCiMBDN/rEN448wfVYmZ09iy9/siizU8GF
2BmkyAmhiUVTqYc94GsrmYp6dVPIcdO4PbwXWYTf9A1EsaVHo14bV8Mk2QN0U7qD
+ITo4fZQmeYNsZXCuNAYfR/1IuToAqlXk7QD8xEIT4aipgcG1xcTeMlKpf9f8jhr
haoAuiIcjSKZ5uC99QJPVRsj2aVWBGhYQd/DJz2ggciZ6vk7PD2xcjW8LMtsClRB
B/WVDNepTtN4uv+nENK0SrfLHgHdxhFDqDtK4Oj+0tAz+QC0+2TrGHEeiSu3onFU
eeKJDFHprYzxyFqHaohQ64aLg/1bPcdjANjW5ADA2fyzzn8Ydx9GwNTiTWy4ULpH
vgokZmQb4ESOoZ+XcMCy/RB5kiJq3/P1U+Ptu18ufCzzAjf3KezpG/8cGRZMUnjS
g7f+nWy/bob1iTJdRXu56c3C8JvHUv3nmgNEaa4fmdNLFvWFD0IWo16R89Ep7E17
gjPPJR3HOXdMLxvu/wTo+FB/g1OQcTEcUEj4BinPTEVtjJRyaTx9TyzFlpK1/ixX
2yS50YbiMW+JspVlcqpl7fStqyl8qHKVFSU+zxGbSKfbkDJPLb0VucCAtPcuPoou
aChmb7srt2Xj27D7vrxfLC7FJtYyi5xFOegshQgLTOKA0e3s1LfDRKcq9EdeaIDf
VcM+er3S81KLanpIn2heo+mNnKwh3CvjqgI8SUoyzoGsMdreZlB2wVrDL74K30uS
AQnV+a5GHaOHCu3h48xbmziV6sIzjCjE38ooS134BxgljLuI9jZHdcek2L03Y7Q2
JOeg5RJd8yR14O20HKxgqeGkg0cThJ9DzCArqMJgBPjmUdjXoniYDzOhmHx6NzMZ
PnlP7g1AtaFjcOuyuNGI3S8jarI7n/byY+WJGj20ZVJyMe3BLRJowdlPGeq9r/BJ
opoPT7zxVkseYcpwliC8i8fAsKiZB8p66GSZgtdiegBXOE9KdAJ0jMfjrmWKsjWb
nB13ox7uloQNjzKRAtRfH4vJB9hy/+DES+G60Rwf4xY9E+tXzcjEEuGSgBzDTvN8
PgPwdWC0y8qI/LuA9sO4i1ycuM6WMlSITDvQwk021cxJ2G3cJdH7a0++7KneD1TY
ZeH0kFvdzljb1yMxdIA9lcO1+DEzjUCXL7jbhTcIULilkRorRViFLLrR8NNHaiLB
w6a7JiNDBDiLe+jO0O4eriuHu0MiTHSl9O10iBc1luyZ8+5srah4rtyLhcHYxn/i
uax+Ha1tEwYB1lDx8/5M+gT+OcoeB1/pHkbRIb3DoqXKvnZ7ol/FGXvmQLjJ7a11
qEpG4BfJ8i/GPOYfXJ13aw6Kow1UMGzYDMQClDZDgGIglbnu/k82ZK93inLfZ8XJ
qBMThLKyVXp7Nb5Ht9DrZH7Dc+9GqDgaAc92DNDK3Inlr4B/tFE6v0KKyxJgkV/F
wBv5pAImmy94FX+tQCxD21EQCHflRvAsFs/oRcHjCEVSfyq6B4RNjUdDeARt7oV4
ekuY9IpH9NqRTIZ/jwlX/+p27r4WaeMOkNeblXNrE5RUsei5sm8o/QiGdCPO/bG4
fP/qIon9addl8Br6JUxsbZSLEcGeGDAmSUZA08bfsU535TZfnl1URTjPjiG0u4EL
EnSGYmhHJnBt70cL30JN3BMwPwOGvYMgWcsCoxD1kQlR9eCyuA//zopbCiRmnhHG
WTQazu5A/Obgog5NBWtT0dUDWCx5DNU9dImKOZXZ+2UI3q+ymla6sHTWVNAHppDy
5xIlW3qpn69VXJztlZj7ntyusu6kGWwfQWwcNmBJUMcJ83zKxTw26/xSaMHZYv13
wt+RPDUO0+Pbiu1OPylGUX0DUfHTVP/Ro9rszZGWNzXj9UFjNI3iHcQFMmat1/iQ
p0YAUKpKtQXbTaHOJ0K2EAuPLqg4YT87vM+u29j5ScU/CtcmdhmeKIs72cEO3tq6
8bFamn+DqSs+THA5z55dSOmZp6+tD0TQ0o1PZ6WM7yguUW/uDucOVje7RTkJHZOl
SsKw2u8htiIQxprg8D3j8NxIsz59J6rdZAufNwX+Ju1irXnX5EnddDhMYj2l7efw
pFxEcvju85Rrox8MLDU435Nzo8rl7ATPbl5fZNee4pOPuToyurlbK3IyP+bHfvn1
rBq2UMMfPAANW5Q4O/hXdI3BeA4bOxU1UAOfdTBOX1feuXpuZJkN03wxpCdhj1Du
EJ9zdOzcuHww0e504SHDyAt08x/KAS9BlSdAP33dblmKywq6QVy0v11YOjpIbqQs
bS8ZvRV8EOsgqX42jQnh/1oHgvo4WS32/49lDBBnQIONtCn4/dMd8/qtPkDgJZin
UtWYTgivr6xw0K+jW5j05+AYcxvEntf98CDK/U0clOU1XKpracCvOUKOkjel7XPN
33j726x57nbM5uV17iU2LWCZVbo7U37IWzTX3Y8soYix5mQ798ao5stzcouff26E
OktoIBWZOxWAl+w1Ix+JM23kmbo5Fty+QU/fASJVCEtR5ti+rOI/lUZdhJhLpjeW
KqEOzusE7YqIuTRCZC0XWawnnviBUnci/l3qsmAhBaQE8Y70snBKhnu1JwadfxOK
KMGDcyYSznNtZgHRhK26/rcFoRUL/axJzgV7PTHqUGs+ad//QK/nfqIjCFx0wYUI
wJ19vCoB1tsL3hylEtbXmQnDisdNdPRyLL8XDwnFQ5KLZcykk7x5jgV89TkAt46h
wa3G2uKus31WaZU9CAaz37vu3LuMNAyofr5LDRA1OUMIoBEcz2gAoCpBAjHc8IwY
HyOjdhJyglVfzDds09F21IhdrGWCLMgpGF+2Dekto4FT18EooSVDnCo7BtjuJmg4
2cQt3VDUPV5MW5LlURLpvGIM/qEYErzuaZYATklWfYfeBl4CwosjSVXrpOYut40U
5U61sw7gpba+4jtjd2lLUMC4RygOGnjK02gZrfRVz1fCtv5j3a6hFml28kEtTcYE
wrYHa78+xopHiyfaNgpxHdS9ZF9umCRrpBz0F1MQX1xoO/2QIX6CyClfckOHjqe2
d+IrI/EV7w14a5XkG665yIpTdnBG/3bg5iAzUWwaoRFl9jIbvov/agieZmt1XjFB
0o5FWOCXxRTU2QO54xzGwT1ofVNsdxEYfcgfgSL0L5yEOhOsRv5pghnU6+6Cv2Tr
OEJL0/VxsQH1jDxG6fEE+fy79PRSFjHqSBqvulPJtV5jr0fVQU2mDN0X9Re6+KHS
hvyLJzS9YQ0VrhIv6oKKV04glgWcggHJ83lRrjefL7pu5xXKThA/qMQ7e/VrdIoe
6xqDdU8zJi5JcBA7G6mzyJOGqW93y+Nd/oVcLBGZfoQ0wZC5GuFBs2PQjKNvOc5T
Lde/rBjGTkmbrgSVKywb+vDtoEE4ESTjOvsx7YymvNtkXcAfClk6b/Mw9KErj/Mp
Ia5tatdPA74KPYm1U/KPNlarZzTXDS1cSnx6hfiEdgC1G4qRakxd61Lj9Sb38lj/
eESj/tanPiFzFB9Dki7ggerRmjeqmBrW+d/RtOvSb0NX28QfdifN1iqp94YwAuAb
Lua3Sothmj9Z8rUmr/dYLitMQ4cdS0JvqeXfl07aQ+aaQJGhblzKxaMy2/27oqNx
QDhYq3W6lo5WLKjVAsKeL3OK+jQeSM8HIF6ZCcm2KdvYvJ0AgZVAl2CS5oO9F3mV
/tSlGjqft2E8EQDcSE3TCXSC4XzDMOT4dxnnKX5Zdc0PvvgmS4PS1xiCZO+DSsxw
+tSYIMGd92iu47iqwwyPS7XHLvywODMJ3rud2wsbGttnuO4Yw396lgsBvINgiJT9
uePF2keJ1yh7+i2cpVlIkbFtR7ZiAJvWI734wquWhPUaQU4iHpmSoLn5qJjmXFke
kKk4vhzz71gV3XX7rtqY4iA07y048WX3tkgvnj3Kx/EOtIBGRUbKOTmHs8wuu8lJ
oJvYv7GmEkPRO4ZhzfbytGWXAIPhS5pfyz7I1elko5AZdCgOkvmfKmVmBs2YxSnb
ZrOLjtohKGFAo39UB38SHl3hJdAajaB7cuDgUereKc68Vs2X6+aPGak5wsWdLKMt
5+W8ZOv/a4aPgkteZSn72Bi5Bzo/XkR2+/Jc1QP9cW1Lwvai+zvglvorfr9whZmR
LCbZap4YxeTkIJMZK42G64v4JYsgq69RVfdqmERRVJOZNB3GprNVJXpd7EzJRFvX
MavY2/MM8hIfxULlYqIIZDWFsM9GrypFbOy0KQP7a/ACAh3+cenXTuXq8bqW8nUF
RK4If5tT6JjpkYX8AEKld00V8f/e0bNBp6suK2wVQD6YOVVAI2dJF/0UcaBP1jKn
LYIPSsUzDJeTY+cabuGI3qJC3ji0jraS/JRVmx+Cyu9f7ZjRgdnOFLFajsaQQM7f
bc/FLgkz4laKljY6R01fppRQOYygNsvWlfLY+a4DO8gRzPQ62MEuwBofFpB5jF+w
hsGlWHGBQGI687unxksIsz6R97fPkm0dUa5LENKcUKbaYySdXtXQeXHWX1foFuVQ
9x1FvEB4JU/1YM95LYlRBsv2r7zsidtUt7BOJ4i6H1UXGLcMwHam7xxoIZO16+UJ
LYtYYrEmy0xdtXQ8boLQCIaQdaDpu4sQ9qYlG2fDHIBcmVaSF9HOH1Er+g/ytRNA
4f3Fgw2G1B/Dl18LguuS+YzyRPZZBit22fRRrlapKRiuDT8MgGQaTO4f043SBtpA
N46EB3/cIWbRjm4egYes8t+CKexfxoCjdrcQjX7OtNegwbGxwU1tlyARrfz3a6ZG
0ArzWuA5sb2lwiPFdL5cr9WrVr3JA4K2TqoEqlkk7hq9iH0Js4u9ofAF4eovYSTN
dZacufoa57FdnO+oVgWnbkCSmAuHyAYte+ebxTYJuhKqxZ1CRb+C5V7XcyieAkJ4
Xj9gfD8/gr+heqFDv7pU3iGdgOBPRsBkh5AnI62hvgZxCKD9qLnCXG9bnp51zS3Q
NoexaXjXiTt5onHlcOgPr7ZJmvJNB586PYeTXjNXLmlhnkp9Hty/X91m+PmmZUBt
pS54iPrV7pf4tU3u98fXT6g7TyDN9Wy+i7TVM19QeLq49lvJ1KlpemcNaTZn5UT/
lp3zjjVr98HJW/cbdtwis6JUYbxctWF4aXJurHUKTCvzHH4af+wGhsULg6SrXfLU
3UwAwn6byWCkKK55Z70DfEs4jHCbngDk83a3GOgJPq3oNgfLCD+68gEm5EiBxzh2
+F11xJ3QpmWc8m5aRzEMJazPyxrwQY67BdiD8Z2+/VwxmOyv2xZiDNvYmHssR5Q7
D5Fo3yAAuxz4vKpCwqkcCG17RCkEjhRCoWbvZSgLYTm35ch2X14SRar7c1UoGGgG
1Q0wM+NgDfMv4TLzfZTIme8FAjf8FRl1B+fmtw5y3KsDl6/p7c5+3G1vHpKFJOWj
jw2fXPfg0ZVJiizCui+l78CW4XyKcc8Hf4bRlN0LWbeS/aHCCGIXVZNYVKiXOpm2
z0ynEkL6e0xBO2LyDkYxa/ZxQm9vT682P5UoXYg9tP2OS4eVvIW+3TQ9xbOMLMtc
Wz+st8WWu7CpMziecdgVS1OzISHlhOZLDE8FaiNxLg986h7pG4czXMt99tQkY3Fp
YIqzn+RePHdHpnNTel4sm7X2HJh1XLQwKar1EKA6yu4Ych7XCSMx/y/+FpLKiAT1
pdH+gqGThudChj7GK6Gc3AQQyy+j+gQu1oG9Nz5hNXPLlUDTbS6IF8V40GYfszhj
rIVuKk6tDUXhHjCNb5avH/Vn4tWybhHWgdd+0uD7h4yqc+jTLE8pVU7EEpcW1Kod
/tHlP6cva6rd8/lbspv4Js/dOlIrs2J3Ce54qdp7CiAt2mlNd6IAR4CIdEuyOgm1
zCIE4zPpX4+sn9xwvx30p4iWuZmXw0NGzkQn0v6jA9TIiwZDhnMgfLUvbD479aSd
Bh21njzmYqB2rSGHCdMt9brSVf1kNVKNrobp2p3Z+6KVl404ggv8C2r0JXZ7yP9R
OSIQmxFPs1wJTFBoWA9VLypB502elqNbHLZ/sJD3vWtNjptW0Ma6hLun1cmCCo02
TrBjHXEiOa01g0rP/visMiY5v8pVzkSFGXWsHrbmhUkrbhN8fgX/QlODICm8G131
3F8CxZJsNNzZCYDtIFLANqTaxhzccsMgTBrjdliOtijjVIwzBGmiKFkEAeM+ZtgE
X+BKS4tzIpjHVi/EjM/w1qre94ME1uHYvYT52LmH89GxAWz8hU6zRtZkGsg0Z5W0
e13YC/25Yum7AfBPHI1/2IOzLf9VxKfMDzqyy6W0Oiq3UkUfYf/yVuCwXZjMae4P
9GU6qSD+TigxmPLHCHLKQ1+eo6VTvSYDlsDSOT03gBYRTHEuk6zT9h4laNRUPOxn
ojR+43G1Far9jjCHVcwl5tG0i+Itv5y0dVjAqxns5ncqg09koobhjzNvYWIImWW3
a+g6L9JcqzwGZTKdxwQfAQa9/K4QrI2K5GqPf7mfNS7UFalADuTKg6d+SyRvcBJx
jKFrJTOp5eF4wgzpvsSWdHUliqDWsJVrBndpGCgne/ZSFDQlfyP72GaSC6+v6CAH
p6inpZWEDN/WSHLYmvl7WiDJPgP9xR3dwxkUPVIW3RzuuEp3qDIa7oFI81R3s+ou
GTq4mCTXv1+KM0yHuY9SHsrJ1Fdpk3H+Ll6WvK5jv/aomuVMSDNucQFHjTUpmB0g
pkXKVluasKMr19WItV77OtD12BFWulP1IISpWxKABkmtyTM3g8WN+TLersD9u2GE
Vjmg9mSZKrdWnjbOybgspteeknYxzbY4asOsmyTSGBhl3YoO2HkuFnw5RvfSvKQp
dqBBVqIXWHUoPiB/T/GPEzgZs+79SZYV9EdqFx5znuRF0RlICyqU2gyB4/QiXfu9
IrxjPAsdTUAcWVd3B/x4bz22wPYSBw1Er6kgKSt6hXK/+NI4wABAjAyEvC0E9eTv
yA1GlcGresdXNMh53u+0gmGDf1Cz/rr2EGrTESAo6C7l7mvx9Qqs8bRed16gRGlD
CqH2NVx3SjD95q5FrCkDHBohAif3xsAGEsVRID/afTtE1e0G6XE84F502Ugj92+7
vdcze+3/E5iUCiVcRHlWZHRt+R4TGaNV+wCFJzsN0OAm2VZF4rB0xexWRkGCoFUI
aHah++4gxq/YE4Uxr8iH3UJhwcKWbyDus6EVMkg6lUoOhuGZcW250waHtGMFN49f
2Rx5/ni+gJJqJILtqColiUQt+SHcRwv2P1b9/wE4Ua73KG0v6WN+X6U+heABFbAX
aRArV7pGXWyPjJzEW4oKd0rwf9isvG17GFHsRh46bZFP+fE/FP5fhZxZArm6iiho
81NfTsDFCiFRomQjU9Lim5VZUjJbPczGC52yL3uwzYc/N1ryzrkgNdKnpE93FHRG
wgKTwlTGNaZHex4FleHc2Wfs8VwYRAFUbFDgS5qjCeoqn84UCjYiCPj96ToihnKf
dZ3H6/LS/vyewEdCWiSSraz3lqjQmnO/z8BFfIz3NH9rlAZEUQOZYkdQiQM7q7IH
JOF5hMjPyQ0Lagppc7GpdweEXBkRwMRST98SwurQwBkwk6kgLu3oREAWFwMvYPIo
DXEYgwLwRN8cige2fM2kOF/SOpdtR2rSxBAcvLBlQJ6vhC5Fk8vrHo03GkV0bvCs
UGLZY3dvkO4Lim28Qxr51GDgI0eCE0uZ6gS9Ke1cSopYuqMADfFrsdJ+r9RRFQis
8elMET7unKx4319dxvG1fbjisbBuk05Rhj192WtFhrU8Bui1+qH6PHu9hcgXAV35
ACP0CuamQ1TPaFf4Oeth6XS3n1R1RBKxYpXb/E8APHc/Q+UhmXLDs+sxxXAZ4McF
PGU5bfzMG+9mCcvSyBKmaFhE/I/qoCwxOVuxMAJHOkMC3cGxR+7V+GnGn7hVjlmL
o+rMZvK3idDYDRkf1NIrllUHAI87KsplK6qbVf5LNu3SEXsoZ4eR3uHsoCpQym2g
I90FsLG5wdiBnYbWOckhbpyuBZw+phvwIjUehjQSfJkgbpR0L52PyLHQDE6TQIcj
bWlVciG/Ui5Fft86ufbtuFXewjwIaqFGZAeMhcSZCl0E2Ndcc4e/wi9DDJowcUXz
CRV/ztDoeYrboIcvP4W41RJRZQx7CqTrOhOl/tbnsrml55VVjWNzuzomhCuuZZr9
UUudKgp2ZlTLSYhjMfMOBVqupGicZhwbJ0mlRb+dgIOREbKfWR1S/CYi7ZXD06An
WBQFxqiDaEXGYifK8Kid/qCqJyRQr3In0DQ0Qv3neiLR7kYg3PJqP3OBbkHOFJpm
A740ldiYYZTx6Enj5An/yebsyWZIvv+1X3k2AabYBuxQSydAQM8j8f1g/oA7iuXH
s/LaLoCPOLUdqWM3EzNSuSN+5Qi35MvIboO4769dOfuwUwI0LtON13L6cJpf+C9J
r+F0n1rt+YnFVy5OnDLIskk7mR514vVjrhpT+psjzXuRtvVbo96dZsGzKe1lStfa
6OCiZrwMtVN28pe4KXx42+wtnhz+LsCrLz3JL5o+zbHG8jx78+0a04eJFl8tZCyU
eqL9M7rAUxaogq56uCHAoWvR0kjY+/xDYlZ/9+FfAPlNXUhJUuUC74UrzgGb8Vva
hxZx1M9IMadsEVp+WrZqUVsrLIu0zZy6Joy3kiPzq/qd4v+hJOwta3T03wO6jc3a
HUKW1plyuGc9tqD6WQIYA1d+9XzwdlU5iLcDVTUVBGGbZz4Ib54NP9srmf7Kfx46
uNIkGgb1p3eZmet/lAztPPENl8JanLylbooAgqRDB6S77r0gT3WnnbS/bSBTROXK
GE7g2YtB33eZyRp/UJdgzPCkDFnlEu99sKNdn/BmDImfSOv9O5hjjXEui+jCX4Xf
uO+25BMrRJVylcZ3FJqFWEfWYN6LPPW6oy93eo33+uURX6z48d5Y7C1pxjpN0IMa
4/Cs71tv3XQjprQFsbP3s3RlDfX684HCDa95LC2tnZlJnTczeFJOTPRO9DxxlPmK
E6claxyqENoc13xwZRP+jXG8YI6jnTvN0ZY3NKQeG6yPn+C0ryKUVFfDVcXAEWfG
V4kYQyyR4khSaBfIECJoYOLGc/4T698Ws90EO1YUGcHduXpTdn0T5nXLg709beaZ
klX19KjE4yGd75SZfvyxmf/DO32ZLC0uxKOnjzap5EEZd8yKr5skpK0bVItwqltM
dib8lezY5aaG9hT+12zYPuUWWyIrFxZ0otD4tn5THluoAHRSfcXoSnbY57cWs2pw
6v0EwcVyRo2U/MT4IEKcSlb1JfYQu/byjN/Ak4mC5J/35a3gCC/oMMDCqI9oYC7c
wxNPqUaeulMZV/8LUjykiQwiWhDrk8FRkXnyT6xF4pfuCSOBg4dsXcFcAlpqXpMB
iyRNcTL7rHmSbUcthXv1uVF4TPFwM3sZ4FyOc7H64NEuDbHZrlH1Y0gV0xM87r1N
kCEPraJlhbUv0LXX71EwZHvdj29qnlKF4qMsaHmmUgpKapTgiR5nq52tD5d0YxfE
qnXqGOjF65J//XmgKMuCocubl03yQRZ3cwBnP6pRsmiG9xF3EgiXRhwzTetcApDn
dRb6aJLCzJFNJVkx81vwgLlOxz5Ye4u6qpTtXDnPB3SFkLYLslRWuJBnlgclT6k9
TaggLg7ItiCUbjr9DlIg07TpczJ7DKSbKan4AvdVFFPqsauEHeO5P6+Zg6gvHZDb
JCrzrjf9DYLHHJr6MY2ghotA3ubGTL3i+0T3KkjT20NDS1YbQxb2vq54LAfH8iHm
4IzpCKlWEjsMYh7CWqqPzqRFkvvhj+QCki2XVDRbCQghN6lHUTn4KT6avGSFLOc4
nhWsWB5UjonPgrj7bbY9LdmqyoxQ4dKfG+ZIo7hE6U1Ul9Sp3xyfcWIvgIwfERgP
bEwuf+N2Cntd3DaSOp9FsdLR+ODMhBcekb1SRYHszGvvr/hdb7M5dPC8WzOIY4jQ
RlRyQNbSBcCLhY1VjfOtTG4KIMfyY4AySnNPzRshtrtB9NaN7YIN1RJOnP5VBxuy
gq2Qdi8sm5Ffx00z12UtrAJId//DWrGIE+j8FbXVM+vqo+o43c2kSU6wu40eSEYB
5dab9NIQSb4D9sikUYU7cuFow2OHzhs0OC0+CZa0GLGFX/pBj1Ej8QroxjMBMGmm
mJQ+u0LubmqCWBkhvGqZ/7l7qdhOpxPUg8L2n2ewrpXSpmKu0HQGIf/srOherxSM
TQAaH4biHqT5dyO0pHZZaX8+MgPHCiS03p6SQtl1E7y58p+rkR2la70wTWHn9xnZ
EPXEezxCKXKhdMZ7MBUHpGfmIOPz2kklIqW3PKftBWoia9j81nduTD+R0ByB0CTA
EgXTsjI2Yj7WGGbv+iFm4fc/Uy2RQCqeY+OiMJvbfX+z2F9VypONIgcOamTlSs9N
ppp/MNK+fjrm4glY1QjD2rIi0u70VclgXm7S4x7NNHuiNfABpY3jAweZpPZKmYye
sjDF8Qi9CiUCORaFJYM5qOQSQL0doPQ3AaxZX+CgmFvcuHkdEuYrY7gyxVV4nYsf
mtJD8xkRutbsnX3BzdNn9G3kjLsswL8W1XZtl5OUe0MpTDH4z/sK5Wz/p0ym205B
sWeW50Wu44dkc6q/PQpcmqrA7GH/eB/+fdQaWwGgalgLoVTIRAIeMh4nhfUFY6z+
c2J3afgBexReLpC6MJ0FKvSGKIJPFw9+VfhWsW5ckZRRhkWrAujCegpTwxP0qC8x
mnlMOOxnUhRWyHeO4JdkKP0/bleTZWC1iW0TrQ5BACppAllXmMMGdr4if3m2Pey4
quNTs4F4q1U1bRwFU0iWDjE+sWPOWYqi+tNu1y15t9irDAaRZsFrJFoCt1lkgkAz
GCpzQNzQ4wdc5QW/D3CnAV1BxVYKgmhHIJ2bDrihPAFNEK6XPwsjoEzew8myMcaB
QatJIKV5e0gSxQKU8Q6SZWWwLrBU6ggbh4j+13WT9GqzHgWeBnv9K3O9B1+jocUv
5iXRcr0giwTiHHETKE2p+pd1p/D8OAzVqpvDT2I7xAXG8PSS4/JeMfQhwveNWaHC
y0xwQjNA6b9NysTQq3zLB/dTZaoajJyNs0nbXTBOds8Ryl3OclXc3Zd2128OhUtq
5Eyn9+Gf9KdCcTSDvDZU0zDvImPUJx+AnzqAFehWGpHEVY0jcVn0dz1gerypOvfp
ru953YeEjAB367ikaEv82FDJubqfryhPn7Ao5cCuNfyMzpnoVUaGKu6Q5m/qbYwl
v5ftoAwESWjVczxf5u2Lr4miodMBAYUge2S1e8b/eB+RYdc2IXl8jJLrKgBDx0x+
uJijs9zdKCb77OpcBQ4Tc6wB3V/frsrbo/yC3z//GiP1LMNlicyW0YWSJG6nvkSn
qGPQ3P+IWjwwf1zSdjrNd6XVJJtuJICnJKpkEVqura810C/NtmeU21b7liyQ0Ro6
dfUZQw+KE1YE+4WWWlaeX4Db5NYIQaWqxczoMbzFec3jhw021QmEa5bH6hwxAOD8
EX5NbhvMLJl3EpmjlaCMEzInzYva0CyC5qqDhXAubXGHxu7p8sYIebgQ4JK73q3R
erD6D5c2fB1gV6RmuSAnHQY99B2ceXjYjjSFv2eb6lbjS3t328e+gvVOptMm5YNM
TIfMqV/wEDTR16cuM+3oYX1Awdna+/xRGOca8laXHC+hqMwb+6mbQtGrsyocYBsV
5aknj/ZYjQL69sG3IzkhSrXU8eE4pAv+q+lhHv/yIIUn7gwHBQ3krRwmHx8f//yW
Y4loZP/k5yVsU1zz3jdANOURja7wIIBRTqzuturoQ11A7YvlZIIyYYiX24tACUr+
j08rKgGHGJ7iIuwPmc1ZgKRRgs4IrpfnI2sWVtYoLFuxDheAKhQ90vCjhB3Lxvyl
aQKMECBsP9VD88PvNh0WgybdGnUVt/ltu7V1iyxR/7EYV2FiUvW7NXaH5K07/I3u
p4d5XsgVs3nliEvLdJzk3vXKvUZ1EzsujVP2M9dmXVsHzY0vVkKtXSYS4Ot1V94H
qNeqtvlehjR5HHHekyfUiAWQkv/ZY+5bNth4ggeGPU0ERRMQ3ceLYQeBoH6mPNOS
qGTtEjYgH90jbt0c+Aqj2M3mGJ4TsisLRE7ReC6fJSuHVBg9ZNnFJEx4QO7jik6q
68rNFXmYxAGXGIFW/Wqmc55iWpv0VkYESHxeEVn7t7gIQqMNnAhQKQpf3BJctbtO
tdc+ftm1+NXr1YnGmOe+Ymw7mYBtVr6PdOToNG8U28F9oh6+inyTf9twXFM3eFqv
+D8T2zwEKZq0NRhn7KJ1zV75HjHX32ZFmU0p7sXpxAsElgZXqqRZRs3IeP5BToR3
/P0WbiYPcgkt9OrwwhLcm3kTYKy/F57GJORVHYDC8lAloOqgoDgWNeHKodSCQpd+
dRL7iUPPHlGpolnjNWRQ0qkEEvvXnHjxSJ+5V8TBDrp2mbL2zF7rv4D9rl7ERO7Q
TUqUvQOepk4XrJ/bGZkfpHsojrQjm195l7uPqYnxxjCi5/A7uEdiwdr+zFRc2og7
M2IDxZJOZoxdNOe3NzbDIKKuLp5ixA2L73n4VjbAhVMI3mYHU3cQ1mqOy2Bljlk/
7ZxxE5uOgyulnibl4A2MgeFENqg28/gGODpxK0v00gWqZgziGxus6fd7hYBI+qdz
X/J5dsyocf0zeaikPHbd2gCwN1D42TvrYzQpEwF5i8e4KeQFRIgMKvXI2RnqhIBJ
0drQokNhUnDfBI75cUXWEZ7iqu0KU7s5Dzlktk3h5yW37i0fvmBuLi6QjiopSKEZ
gOLBZC4aqqTUF8a9gHQhM7zbwAVppbOpQ2tISmOeRXz0OZLBiFWfy1FqBKkFHY4i
Imqme2on5XP8wnwpd/2cGw+yji5HPkjjUz8PjtRw9542QSzHhJUoa/r381MPTEOY
qRUeLS0f67erK2TMlQPF4UpAjBJV1b6x6iZAlQJGITX2bXTFjlim8KeoZGhKnQBi
KPt68RB8Z8edW56jEotorDFAb09iOawng/K0rD9lBqFL7DadnUCMXRtY9tq28SDG
ZbmrP3mR3VOG9pS82b0vMK41Vx+lgsxk8hlg9I9KNCg=
`protect END_PROTECTED
