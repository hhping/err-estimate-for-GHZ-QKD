`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/nSqF61n86EBtqumUTt5Gk1oOBAzdVrJvEkgHMQnHZLOxtV+9SKC5XwPyUK6wNz
ignavbhvL34VRPlxFk+utbmWc/0IGhGCaHNKB1jW2iJyGhtVB/YKMdn8fthAiJYV
Pfa+gnUI2FFcMqN8LwUNZNV9FE4880PVU7j2H7pptWIDtSnYKNTHxAZPVgTdHcWb
spnb5iBzjPe64m7ZjbrjuwcSTbxnlGb7NaOo00FEcSNdm+PHexXetwAKhctzno3h
FGD10LmfEigBCc/hLwSxS7pX8gfj6CGRAz3lGaKt7VIfC24sWUleS+BTkFgzmepr
bYaEOnzf2TCTQij1PBJ4AYe/V7Qp59V4FTAo1IGS5zJLVzcD80IoLiAa9fTJTqcG
0AlIUdquIypukbi3IN+sJ0CMd1ZyRQEiAUxSDq72JslrmR1Pp4BppH5kiMm3YUl/
NgaYEExtrTyJLgVX3l0Zp+rzcEjaVCT0nNLaavSxxeDnFH0NBgwglhXKCmyPvCxG
jBca+BAyslXBG84f7VF4b4GdJj9IWUEQ062yX9mvQlGNnw3CsYjqd+rPGsk499zF
9taVQQMWhhsO9LG5dHh+xmIzRlQsWrui/hZ4s5AL2iBPLGT5hOqz+NjcBHRwInDS
xJR1a0JKghYu7ShfDHsQhYKM/WjuV5xD3qSNxxcWpmEcKVGUpIgVQq4qJ/tgsfzh
yPRHPadJT+FH10fU6zzKIgtdpT6mlTw8fEu2WcpJchZN882/hmZlb6p09hvo8uIG
/jeiEY2WS73fYuFFl9BuXqHc+P//f6S9r78T1+ikg8qlyvKzuRcqTyaYVZbccBUO
/S8DqORZPbQgAmJY3r/AdSre1clOg/68WfOITlRNKXH+9rRHu8oYtJNEPijn9FEj
7IdBUPLVUvz0eZzguwtCCzcby7rfS2xrt0gfWVS17nabOFwF+UK7ZUdTWFwSZDMG
zipJfoo/jldcqZhETyerhBKLTslEDnvqyswgot+0P+s9eQHdP4vV2RtwRBO6fcUH
2EzsDdXmQNN3y37zL2wYC8y6IMEVb4nkLlMLVBqSNd6kNnnFW1QGvM5EkpzM6/c+
/bdC0nmvr0Tlt93s0H+EEwJvVI2lnC2/B11IdWDJKRBie4FMTEGuyPWE9DRIQtfv
iPiR9xoVovi/nefZ9sfBYqZEGM1aVgmikwHBbgHj7N05BwB8CBBCrZbpGI4ElxV0
4xcyqzUeDfDtg/S2x7oL62D+yEYYtlhv4k1Uy8ZqxMWhkitkTxZrEwDZ1avetUsp
t9fwVHHpAbh7RePBOTP8oXQqs1jz6GOw61uSnq52y6eVcjjicdF2g6CT9aeu7VO6
4Ulk0IjXPtCCkmwk34zXw9Ws1Sf/tkY4zwxKYk+mP76By6wSycxzylLGV9TlecTL
W+r0wdMhqvq6XUY9z+yM5V8LAtvZklzRlzPW6AvfjyetQPjudegBSN53SKWgzd11
4KKPbfj1fp6n0aoYx4liWTGf80cGEGugifUfjKuuzL+l45jZmh5EDAib85LeogKp
hHu+W8d6q821jSv3LZOJSPZsbbVxbt6TNI/bvakTm4NHqfRs1JQMycrtyI+7+MYr
X6NY7+TzApETsbMV1jkzWngnxSEV6U7su6ssCM4VeBC+i3E0poZvp5BhjRdWAhIH
Tvw0hsRzsRTP+B59kF2W/nLiMvEO/MlVmicQ0mteMI/wgKkeUTncj7sWQQdVVmbf
2J+0YtAFfQnlTF9PGrMzSOzXSvcoY/x/65O5KXkFJj5ooWL+U87w6xjqIjo7C6bu
DhKErR42xEiiMCaXi8FrD6aslr1c/vUSFbHs2CpjrYsrtQTdnbMy6Pz4DeThS1B7
GIbBK4ozkdCe5yOnUya2wSk4yA3KACImmhGvdQyxu9r5MyhfyPGiEj9uzIF5C7ww
mk7HqUyeG0LOnRhBHTwTk59G5IkDbfM8I5aTDew8ESRBD/IlDcoSSj4XYZm6U0Ey
3zl+ESJfYeiv8hZyj1vL4A8Vt6bpAOFw3fKJ0S/pQa6VJ1TiYEVR6jsnoMRznUB0
MwPyBWPWH7+1ExEsJ/PcWmy2yKO5q9Wfx0XsttGYZ4rBkX1QLfYozaMd2PZvIL+E
gxVKwgStMyVK2YEdJ3sEZknDQ6RHDZiBy7NIWSemEwJuksAH/kBdjToufSQjA56S
+ZCoBvP+8ecrGvdwkNbnCNgnUbMQnHn1J6YmeSAHQuY+RKekXjHoR6CVfneBZNYe
2GW5Keo0PAaupRZn6NvQih5KaVOg3YmKLOOyix+pe3qq4y0RGO7trflVpZHubPrr
m8SmnlCs7J5EkieFQ3iIdMel1I7nUARK7P89lZ0HfEFdw5KgM+KuidXK5JtthQ0C
b1o+6KGp8Qwc3V6M8P2UMJeOsTFVkLpWaYZdT5c62Kel8JPcFjKnwN5xKJH+pWZ1
Jo6rdxsDOU27auOyCSaS1A0Mqt5wq6UgWv8Q8icFX49huatBv3Vs3ELsX7cEwg7A
1MgeCOj+n8PL32D0KpY/1T57JTf+3xCAGGsk2oRT5Yt/ZznZVhnvhZFrlJrHEMwu
vRlkdmUeU6yV7n7k72G5Z+yAfKjpUnD/Qm2C5nMmu7KihAJgCBuj86LrSneJA+sA
w7pBAL+K6l75G5lq12EPA9jCF4mn+lXNuaE4nZKnXNT3okeBNoSLnzJfMIJ/V7WF
oRIW2pVDKeI+eTksNNfkjZfsLSSKp9eZ68hr7k5szUUICNnUUVhAxh0QVwr4f307
++W1FzGMa7LihFNzLck1Qw==
`protect END_PROTECTED
