`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qv2oGf11VdI3SE8gHjlA/UPfc21qyqe0aM29OwvVyEsrwfIBOSZmdQ1L1oeq6LWw
qPnLuer4Nja2BgP1jVWm3ngJGw0lNpYlbf6LZk2oLLwyx50BEhMv+j+wCVF7F4Qv
fT8A2jgOU6sqCRaH8Sm4Y61DiRir7rI7vw6KPJ9Ee5qLeAPZNJW6RvSuvgJETrHH
4TF/S8aoFuHqArH9okPSDo8r7IJZ+l4DAD4sL34+V1sVyzh5mGaxWTl8sfBd14K3
MN6H0Fpc2/HVgBnkUlV7cEKpqHNlR+PVAJ7IyCOaBEaoHLyt9Ct6VHFJuM29dkUJ
qZcax5cFQkZ5vLo+sQpbMqZKCrz7IlqzvUzizJ8fi6yv0//huuEPgEdaRY2zlhey
ByiIsC6MHgzGtvHOzOtalGlSRu8pjqn9dBXwMgFsILCZDzt/ClvgQziPjrnUINWE
r/ClduZoIgdukygJSaUCORhJOzgMFXpwJPXadw4vW9qkPSeovx7umdpCy4/eVLx6
`protect END_PROTECTED
