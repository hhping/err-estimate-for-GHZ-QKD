`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RP9/U0kT94m5785Z5wDkBWGJ1g4XtF+CzODzIy5YAjOZN/RDdFIQrwabWnmjCzTv
/EmRSUpHZvSBLE3RtHqaCRDl6h59WOf8/KSoOriPzmAzVW5rAIL2l9/KfjfsXkMu
/tJKqXp51mrUkiQTB77JIOv7ifJBiUbwfXFzGQP1SrNWwcWZqFCWlTi5rKoNPX99
kQb/ASbi3paJqyAkHIegR+vybf3kLe9bTmKT0/7zJ3hrZl+TYGMlJZytby9pBn8M
QYmfm2pi3rQpk4XMxj9646PnH+u/MISrg4vNSrNIeSnt8hOnWLer5WK9ZG43Hg7B
Yb32LwXGFnMcbf+ueQgefW1qCwlAGt+7G9jaAKKY/9y9TKRAY4kJqVojsTr762S2
NLeeDspTtc2YYhVraNn1BS0R4GxdV+OiiphI/l2RT0M+mpqSq2Rh1+F62rQODUsP
wDZjzpdlV3CDiWIahF4+H/H+4DzNEkx8WVQYEspr8bZ5kQPf52N1MxTagTR+WtGA
SX55PSoYifbq+WdoPw/zNQih/Q4YhwnDwjYSbEBPQjya4DqKJve1YJuudkuTHKHt
vx7oaCUi+hCkPCFN2vNGgLRZxzp18Ros2gFwWSjKGjweveRsASQP169CwI+V19U/
8KntTx/rtVUGP1p95Du6ZqIxGLfxm9EgQ8bY+UwAsnDwfpc3v0EhsU0OE/AqXxHh
3Y5fEnLWEmxlQM9CkrSZvPVg6x6nRdQkRe0PrAwzTzOCU8kIbKxAPLZBE0K8r5ly
kqumtDhCxXFhHPnownmlxf3xL62NA/w+fktaj2pVUu9qhmua1UxSZoCfz3UMDBJ1
sztjxpFWMoRbQmJ88ld1dRNkN0RBfdbAguTHZOVp6rV54qGbo6F4xRSI2xirVjNi
WVnsVAfnBD9Ckam1Mf8pfYbzD6xpz1V0glgEOn7RGsyu8e6/v/0+coL8fQ4MQfpd
xv2Qw75P3LPu0vYwDaH1xBfMjzwT0YR3ypOIDbbh8cW4WorP3Vvj6coqVirPgJg5
VTNCIMrRAuR60YM1mn2nJc1Sbw5IH/SaWWQVmPBNf2P7mlei75Kj/LWkJkyduDR3
58SbyOcSuvt6wZ961KRvur0pToJ8hSBsmdp9NifjH9q1Wr3BIapJFsAN1Zs43FPy
W9Gqh6C1oFVmK74IAuy8fsCcj/kFvn9yoqq/I5UwhyQKuBm/ozGCVT9fCBi1jV7s
G74T6KPIaMnJe/FOCY/PSYw5mdDfghPO8eZ3YuKZ3HfL+qakOzRRxHx/7GJIA9f/
0x+u2GDPaaZYYMMiCfQCXffQOceVi4uccP90IyIgfM3l83Kn5E7HJNLinVgkl0uV
dpZtXq7ozH1pviXfjO8ji8pGVRwD1EAZtbvQfZG8XoUshE6tU97HNwKACFyszjxA
4qnNqlD7z0zt2BOmijU7hX3VLAzdCD41KSerVMug11bxo7rWmQRmPYLn+uQjbu86
`protect END_PROTECTED
