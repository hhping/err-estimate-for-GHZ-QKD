`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jC8vvlCrl1LX0McMaE2tWv8g47FNLd4mO7+NMhgXeK4CByDr/9OPGC50J4yViD8w
bRANJr5jZdGbG9FtldIts4+V209zVkopey4HY3zG+FGBLmSC8EzsJI1w5IRdb6gw
Xwkcmcpo7+hTYBIMGNWhat2gmbLIFQHWIxOeJ80lW/TBhIt1SpvBKFrtwldHyevT
pUVE4b0R6W51posga+odBsoCy2+IQT+vapPTwPmiiuYecRoyLBrnm8EoOYOsM+WB
e0kfnsWbzZA4/BzX5uFUvLz1J/5QRDpSQUWZkg7lqWZbY9uGQHErrQKjIEboSBCJ
t1lhN/uoUNs0uvoBNiXtKa3jfOkFyHk1hwDuPoFLcQBB2PWu00XSRMS/euDbybRc
vP8bjbss8vI4KejyC1IWu8wp0J0ndm+ASPjHtK+/x8oOdRhKlAiH5HMFlK65dSqI
FdrKIrnlloBVq2tYy+1aW1UabRoXMskulkQbos8JVYbXFi8H80zLcYjY1mHGZyJg
lLUdFYMvwNP1mbsFmaVRz+bA/RPLDagmn1cDAZ1ylrlxRYtok94l66yVcew9NmmB
YGoGDd26+wHcMyIPKjMZPlTMlh8oc2MOYQV6bUQN0RrntwVrCIBgLRMpztqhuvEK
1/ZeO+sKkt5z+UHGiYoG2vUoydoV3a1gIAWDaBOw4OQ=
`protect END_PROTECTED
