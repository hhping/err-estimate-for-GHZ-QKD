`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyvWNOJ4l7/2VHTrum80R5MU8NbxpHbZqCwIdngS7AvC2OKN7fUSxvfx8bFuy3/j
M2sUrNpTY9ylApW9EIE+mrwXsHTKbv8D9QXplMYf6lozKFFT4xfYBXwcanGGHAR0
0U3255/btRCRM6eNJxxUZpiOQJvUpWGBqGCbJv7UaX+Fu4NHyLZMGQZEvQOQLau9
owh7tGlQikSJS6/Vfxj7ugBqAm4tkgfMywlC8G8jQTvaxK2pCSwiyuGJHNJgMHPg
H6GGb7d4OOQhXHHvIHqvCDHeFWA9TKy1eZVYwKexp5ReKNN7BqUGAtU4rnHEluzu
tG0HnN7Ao9wMYXat5IsbeA2hqPjTqHV4jfm8chL6yS/PnjXSvro42+WhwcrWudvQ
uEPqcbcV/dnuv+U6fNaY8bOHpJNa36nD6KmOB8YiYs1HUAf2xXVD50jgAFrc33ig
x55MxGikhHfF/GwUZdcBYtUJgTRrLOfOsDZp4lgVSzTfa3LnYi/3MtxiU5q33Kf5
MJilLZ79LYd+F/iMzu44IRX3sMbW8hvLde0IrCJ69RQtmXRvNpFVcWhiGVyYMTsD
fHZmYEDv+vqzy8CD8RldkUgrJj8VrBgPV0zeA70y2jevMjXn8Tqyioxvko52OOa/
MsP21DAOvCmO0vYgAQgJbRYNE6YpuvtUkjJPz2pNz06Ji5CXgvraKjf7DkFHIvIZ
cnmNXOjAwJgpnzU+fNwbAspu+ihDcA7MmQ5mUpcw2nD3UsJjS8Y0RCUfab8YgQj/
wfAxToCKY4//OwQNs5pPz4CP+ZudaOMK6di7UjXOjTEFkwgzn+z7zclBlfFFlSi8
/tzfsXeJSc1SzrTUTHTGuWxkcWMPgIISqqVngZBlCn/HsBVNJesycfR0qiiXGMqj
ACbBg46c9kbHGVGMBvKbN0utXRRko7L4boJ3qsiuH6etr2ld1G653CTARldQQKf+
w0u2C+9NwJXYvAtozLGPZshePDoCJC+t64g11BfdqljWwq6rK9Wo7sEJOxZBtVjT
y5Foa/jC6z3a3HbqoiijYdWWqOtE9UW/jNxcILW8Vl8Fc6/JS7ZLz7i1SfVl6ctv
cX5wi0gpdCrEnNR12vhnF1q6OasAnphpEweeJJXPEy/IOxCJsLNvaq0fewStNx+r
QkvAel0uLbpT0O2NqwZXFJ+SCqWU8iYc5Nj8VhRKsRsLg+RShsON0GBzi9seQyV/
+E+RqrDqQN7ZpSaLlzCuyl5P1a/qW1hQ4pZ20Q1mxSL6FrYDqFDrp3WzT3wnyNHB
HuRCsqUP7tbdT6jlbQUEBKVZGWq0dndvBRETXFi9bjYRC6RnSkpscUR7wi+CSHwH
SOKfmmfwGGmncuk95sr39ELQMNgTE4r64JI+lyUNFTSitfBIxo1BdWC2FMSvrvmN
BvdQIn6CuhIuwzlDZulNU91u0sGxFazukutznnDmY2BLWisK6P6lp/aLcVGdK165
86AknXRwvmxTImf2m/qj00Zg9XKk2v8M5l6soy+hPO1sicNZHV5qAtelMS3NIJGs
6p5RIInJYLR5davKRkA0csT49o/Ohzl5OdhQNdXSvojAhbKBaFQIESwa51nzIYq0
GQw0PDgbLc39C5VK++xUv9gH9QTIRwnT2dQM9WnoYMs7VoOkAPGHFADjaJQF1a+r
TnZzu/P3GzhkENbstdXc21DD/HP2wO8vHaq2whSE8+EMExBVNz6S5ccBsVoayXHn
xjG7ajIfR4lx1M21ho1ZKYXtQc02i7VRPwJydZIiA2NyJFDRJPF0BlgchM7Us0he
elrzHM3QVuzlV9BKyFIRw0JexAwm3abB2onLTJnJH2+SYmK/RkBrkVio+Gr4U5i4
Zw0xDiGMuy6rEKycoxVaJDeM/uR/uIHGy7IvPVp3tG3qflGXav28MeNf0KmytWb8
BVmyUSLP4RI9nzP8DbjCuHs1RSip0lWhMb2PwvuzUY85PYiU8zUSqUAB0PvxHTPi
r694dbnQOU7gAnay7kUcbu1UJuaO2UUlF7VgoJhuqNkfwwOugn7I4eBYkt+L9tZL
5FZbOp7HUzU0WXnzPGEmuT2lVxeHR4Ob/xx8fRyaId2v0usqwogFHgpMN3WoeKmS
WDE3bRB0cCYFuPPn1D5zMA==
`protect END_PROTECTED
