`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYY5q4tA5JG3S8fQ0c/HMfm4SdpgYOeU8BMe0Bvd7kR146gGHneGYhr3qJspRhZe
x7DE1S1382G3j3kXwx019yJmlTe3HraElJoPrQbI2yvGMd4aycWoMlS8y6sd81qM
STInmR+abnH4oFkyDsMJewW3lxytoOaPlCBzNRXuDK/rPkAvXtrIqJagNZkXdMVy
/wClMkSJers25+WNqQLBy5WFqV1FhUJHG3QbZF1Are4UF/WVna6pWG7dD+rNm0vh
sbZw8At9AzdBJieAhVLLzWSGJqVOFHHwWOrxQRlMde28LO2NNQU2hod4TBFzJh02
JXNm9aNOmzq8EBCxtZjL/RETl39K6Hx+fA8kPu0IxGDSia5cr9q9Vuhghw59i6pN
D5oMAW8Z75WBIJvq4X3eWdz5uTfIep9+Rlap95wB7kwcduW40h6p2Ik1zDoEUqFz
emX1uw3B1oaZgiqfdRMVN9+6J/HwXCdd72gCBUEycaYezJDek7/VRwfVgVA1Ctr1
F0dsAUU6dbL2Y2gDzgsl8whbwEbON6fky26E4PhVGf7epyRKqcok0d4P/kKX6HSp
ONoWMhPV2O0vctkmUBp893ZM+iyraiT8AAlrGMjIZWdMO0mmYoE3LDPXADhZpUKV
5c9FAmjLv9EGyJZfpZ9LwqUhLX3b+hDvt0Whbvvxox3R53dEmpez2moUbo4wpfdE
kTBpE27ywo9VHYtplwpQApH9x14nCJE0OLqPEpETbUs8U/scLZX7HHJChc3jrEO/
CXSaon2ZAKhuhe8WuS4ARNAP6IvHoDIqaALz9547REv2RKLlfZqGAvTjbh1+DGkK
Uy5paQNquHHseEntU/n++TFC8FclF5sZSC4keUvVfIp1dO0qr+4eI1H+q8flUkG+
q3wZtwSuD+AFlD7czzt/qZ/kv+qSZyBsTg1DocTK/2dxS41v1hjGV2ExuilcDwJH
Am7XURWMDKiEpLUyp3rTWDg8n415KDaBwf4XbhwnopvhZQDUYqMOo6I75cSmKATx
oPmxOvWyUSSVCvUBby9L0idJ5GrNtdk100uDOqnwSmM2IPLl6unSXLjpbtQSR7sd
BRXYSWPoRE1kv0pw8AjyLrZcOGxJ1UPiqEIh7b71teRZseADwtW1Q9OIBlx9ZFjh
HNxbCB7cISkxNj7NE5dlWtSn4KAVpjlpx6O2xlMqzEpXzg/jzh8Dj3fJiaVrJPzx
kSrbp5pBYw5JVmB8q8k0cvbFDBK4z2+05eGR464pMqK2bQctZID7oGtzDtS8CHsp
oVZItJW5JIJkXEmh+seyGp7uci0w1dkNGIq3BSquoYKI5CmHYndR6SODClIDckdM
CnTJoAkOyXEf52oiWGHq3viikp6nDtwRhKX+xsq7v9v7926KVybhaMai7UBNyA0y
AAZwA93KMvJA3xdLtQIG6Xf/wrYLSLd7pGfNxSN8RR+DwpK3BQyNt3nAUZrSG+b4
4THMML8tZUJE3qDcS6+9SglUOMKuj8xCZRwyqqGOQ418Pb8gWispXjPYg4rTBRth
LIyOdGl5JWhExSK8NI6DI8ssgaA94ACjWjULyvERUB8o9Ux1llR5aD4h4luF5x7t
U5B5rEJdqwl9XuwzfZ96TJPxvrWzwxy3aHNYD7jLMtlu+58QZNsNWzMLqaMdJ6FP
LMGPCX1bo++Fk4LtYj5Z58lvG/3Of01HknqvgiAi3YzkM7v83QwIScWl95A4+YMy
PSM7krygOvmShep+2TM4CllFRylflZHe/qYWWWvnFo2mNGdKX1fz4qdqtex8Se6C
aWp45ZkVXq23yJZwY2Cxn9XCw9eNXPSO/3jJ8lLi/f+vz5sUH0yNVdDY0D9A9sWo
f3xqqFWaaogpaR5nlJRK1HoRu+NjYGXELL/druHhpp54qUZll6Galr2vNwSCRgq+
pl5ZyMmw2nCJUk09XtfS5qWSnrjEHGJZGs6PkiVCVbiztmF1y04Qqh0c1UVV98u8
3lIofF7MBK3O+RMjoznCeSJYKAZRuJPtoMpIr26eZPJYW+G6VRPloJ3DkHonQzIP
6iMIaaL0eI1fYt7c9ICOENhSi9xROyRAyo5aC3aycgPbWqFxMc1yUk0VQ2bkP160
SGCKFRReGx09eKgdal0TgWLciaZKoVRlQ5SWJeW6RqBoOJOVwEOe47TnW/9RDNqG
ZcgNejilGBDlwGTnDSI3ZTAXsIoYoUl4LxhgYDDcFFlDbRWL+gdksruKufntF4mZ
T/KY4vYDPBWioKPMnXz2kIOCFo9lh5tddlK9tFJTDKo4v72Bmt/f47/yYnqYo06V
a8Wzy5B+Z1LuXVC16gYzr6XV6gZXpLdIbhe+Fq7zvtuAovB2IXEQ3p1+fDtJEkPU
uuA2zKVgJKEIY+wnMwTKeE3FEdaHdIK531RyvwZiSvw/DnI4hq6y8qD+J5Pybt9X
wdXYxbJAH5LSDVgY/ZaIDz+KEqr/5GBPXcoJyQjZ+Rc=
`protect END_PROTECTED
