`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
260LZMm1wqzZVGfZharZ7MAsZxumok1rfgpvCAPZy1nYoE+W51v3N8ESUaw1FLi4
yeotfagk8EdYRlsBfvA94LaHS7PFlJSMZ+SkP5HuKEvKXiXJibrw16JduUBU737e
Q0F9IlESeSxxirsvrjhJTjaoYe/xX1RNphVB5emHIzz4tRfyjjCsQJD6eTSV2gJl
Him+JxtHV1tH4HsapeqUZRQqt9lFnMDDEX1TGNBVvRYGNorS43mxX2DywvDluKvy
DvKj5HtSO3iv2zvfOLhCYp/RXspEnd1aE5xxfot8LvgMVfmLMRIn/U7EWh/lrFAB
AnhVicH+OPQTSnOxbWCtL49q+w56zC+Pfe3OmDh3nlurmEIEIE1JjAcAsba/1A1U
xKu05iMdgTvTo8qY+YY4GebHDuUNEwH/I2jdwIchiuoYyxqviaJqqY0aMo52dW3R
xw2Rv9KwuAny4I+vckeIRhTfv8e852/UVLNopJL0NALhJZVzlFJ8QyKJl+YJ9WNa
pv7WXAAAjcyx38GOAyMiOTt3TgNdgB9nweUgtyL5FadCn1qd6on/UO+uUhIGdPRK
iwCgyPAUIF0p74Cqe2/Ee4cX+Xp28D6vt85I9Q+jwmBkELmLIulHs+5U6RG5S3JP
s8G90wLYFn0QyMHVHUv2mkYPLIOLwFiLpTIxW0AqvX279+svCPHieGZqH7xGFgpD
+O0GYIRQYy7eVylfVQduXZ0VHpY2Q5yy6J8tR79KsO/nsH8AYu9bA/MDt2NCeDsQ
IGPIJW8HNpUhZc65GLiVNygVns3Aru6e1++axHN15XLS7PPJvcPp6o10i0MYKGsA
nqC0zTHsjO/eL7QJZVfSYPgKZI1JQRqOnUEKius7/w7OmeICOx9COGo4pHsJRLOe
5HZWFPIhD7eRYIiJzSGOUoiD7JgccpA3pHsTonGnHUozpiGNkC4qnNXSGaSM1EnT
vjhtEXtXxfO7FAuLPVZVQbiEWtzsFmHYZjgmSqsQwKA=
`protect END_PROTECTED
