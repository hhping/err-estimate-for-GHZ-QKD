`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRRXE0ssn5rG3geDmldhR11msCLB3uY6X+h+LK52SfykFVt1S+6TTmzou7G+b6iP
4rvIooJ9PH25xW1kLGUUcchbWC0+wyIneFKMhru/O7bEa7QjBr2P4uvwZ8tLuy5g
USRJw4ZA5Y8DBEPN3McePx3X7lgSHgkFn2JC4WIOz3bGp966YSoaRPdWnLU6X8vj
809S3yH8GyGoEAy+8VEXfFO3N7Ilm65YXgvyu8rg3JEEfc/uuZdPCU37hamBmFkM
tkEbWXurzMSDGt4CvDnzczwF9VR5TFJ/TuAtwxz0UIFJBAojEfznBv12BXObxhFT
1P6A9ILd2uhy6CjJqxsbWd02NaL/t+1NxCmK5JuNzYfQbi6jz+pN18kwkVJp1PIx
zVmq2dlz+B6KhI5uVVYhH2u7XFFUcHEEtzniUIGEYkGEZSSRUxBY+zK+67Xod3tB
OaRhBY/mCY17I3e6SUd+0hAF/x3x/dvIFNW4jb7MqOt3cBxbfDs4b8wrQeEIaD//
VYKRPaR8XytZijICO3PIcrhQbaRQrupmeDTX08cQEUVmC2GPEcQ/QXVW67BCKb/L
pu1N3BYpK98p/7B0V555W/u4G6204eDUlEw5kVp49V0gyX8u/mqOHGoC3eARcf/d
QHxtXMGBIFN8zN8SDjad6Aas0fQnfNWMtb/XzZdJb+2B7FETWkTbJTVa1026pWGr
fUwsVWJRECVEgvTIloioHJqXBZ47mJDAOw5mTNqMFc6Y4kAhRnqBBl/jlYkRnf5b
BPLZ67BAHX1tXrqgJf4l+dQ3kEZVwRbSY6Pc4puSBDBBxuJ/7loP26e7hH10J3Af
tGNT67uCl0prvEGfACcLbnEIfPJHFGpvwArrStaizW8cidbFzgvg6x8ivdqKTVfL
lDaNmao55gm1dOZ8DDB0Dx6Oka3jX5bCTkic64mc1M69VbzekMJc5FOnyqKvfJ+/
cyXeRcDc22A8r82Ri5r141qX3jiaUMtWJBu4Yx34/96dpA92pDJ8uYCB0fLxw9++
+B3L7JpKTQt408t/RDvnycK4/HQLfdTNpk3kw3b/BLvXc9Nti0CU3Fx+bjVPgkZ0
5MW59gCPbQNt3fPz+httaE4wiPmddcNIFY549wr8AW2sy/shzfB3Dw0dO45BHyVe
oXiDNlGoY2dBIKNGKRkvWpW8W+RCJhS+MhH2/8Gb2s3bg+WVh+5kq9ver2Y2nRfw
I0BtEDH3honSq3/xWbS38c7r8lCCmxWI7W+g5dQcEtjmzkK2biK2/AYilkLBM5gL
dFTL6jZWt8jgcnbFPJC/c+xu/+cdeAXL8+cAoDJq0Rs68qb4gvRsvDTcS9eRJ/oL
hd69EKt56Wh7VSOLGoaBrRiyGQNKzXVJzfUk/a/cO+JWUXhxG94YptxZSBI3bmRs
j6KhTGSE8/1LqfRTYrfcC4lP/AxZZV2DGmLwJiW4L6PrkBYvbRm73z2SOp53MQeU
B/NmDUH0jR8uySbhFyO/N3LItt6kSLFVmoRhDkV8jqjD/mPu/uCSO65z4H/Doy9i
C7J5OgV06//vKzMwfAt/CqJSOyha4vB23ml6cT20SrUCTwIqGhhZjq32N+rD1GBf
Py33bP7cyDb4joGnXGBKSlnmtcCw+YwaXzV0sXaY/BhtjBtJU19byh3pddh3zP2W
zbQlOr2oLfUhIwgZLbAMzeHFDVNLb3EDxTNuUNyIGpqLj4tV3Y5vWU1v7SN7WVxG
It30s91PJcew2QRWLL9aiIQiMpa5GSYl8lBqG1hCQwUkoBxHijX4Ke3xWXtMvoVW
JfBo1OPfHx4hlivDSezPL7SaAL2h8L/B/rUDWzpARrgs2Rmu6x4dH2TYDHqzIaKP
rl36e7NfEK/zKYTQn8ajE8KAV5LaB+Y5ykzX6id+MYpopbpRqXY3CdUJreyGHuzB
ZdzXv9VYPif+oZXmYmfm7AHODdsinYU0ImYcr6BVzwL7ybSEVMZrdBFtpfOqkLe5
LrKaRDF2Db5Uab4WEgPg6c1gMDtIisgZ3iBUZWDnBTKJr6U7tbOyigR7ORGoo296
NZ390+jlOm8M2tn6RYSEVLhQWSmsyjVKYL5ZsEJ5srQoJULl4sfD1jPflPsXBnSR
1ae2lTK4yKfinaFqh86D5rOmcewygjmQYCzPZvozSXpylumjM9+Vj/Uq0MVHhlCd
QBSlPd0RYg5wPwamTlUL8rHY6YNtH39j8P690KD2a0ku3NgSFmM+2QKdnaRkPn+z
zXt/qs0XLOpfnr46gf0KKL/RtD9HI3zGTdwR061Tts5o1sOuG9TDEQ1CUw478xyE
AY7Rk5tN6HjDZOeTOq5wOc0eq/VAwBAqAhXJNprsAIUo0kTRPxoGaUl/FDtcFEHH
vnYCdJ16gsWRcSLmtf/Oc/VYGTt2aIELxAHaO1XYlcN+Quz7zxXAgEbu7WjgRho7
Bjov8t1pglMXlIMJsKY2VLA5gE3kZSCwA4TsVeuvMdIwMfJruDGomjjK5a4RaDYp
+h1mwhavjv36aQ4u9zSZ0uMkWmCLx6Az8ZNr5e3oOmgTQRloAQCLenet/OqmiRt/
+sTkJDjEfVgd25pgjzH/Uy/DyzGWvwmK6sajTFSrw1BL96dYIdnEKNFPgjff75Td
4pFoL6nOHixcEgP63FVWl/AOATVjGOX/wa7Huw+yIBxAMgPn58f/UXImSnITxokr
NMglHS4Qu1XeL6TVWlxkH+BNeBNQ/SqbpGtCBw5Ry50BBMUYnn4/QFf/f0fKyhqQ
vTdEAMXwIYayRIbsuV+Z/W2190pU8uMA48Q6LApv5KiuxCyR0Pqa9BfszSn8p6DN
fe8ZJxIckiXmO3oWoBtC6vyeNWWyNaqkl60JmbtlIIayH9fVOkCYoXAcmtZlcWu9
ViIZ1vvdwBMw0MDfttjj8SqrL6VGyfZsMLwM7DzHR4+3B8dlH8vQsZlCC4xAP+mV
kuhP7Hb3wF9tfc0N9Z3VdR6vPE4Y+wrI0jSd4iBoGM+gW6pjN0FVPYoUMTkRIsuk
Znw5CrF+XlgnAUZy6yp5lQ1pWKdfGnLER0XGRoZpYdoni/EQaOSLzZiJvrkI7eCO
t2HDKVThj7Q87pdIVWr5A5xgaEe+1gPWugUuKER8OjGeBYhCgm0Vufjtot+iTjp1
jUt1dtuAS0Y/odck016u7c4C3RcrPDfbiRXH74/Vq8IHEu0JEx9BfQKXEnmlvzaB
0ih7BRwi4cpi9iM4ahED/jCwsg7M/0sBrgRihteTWbFY/1pi5Bhyr/SI1t69Xneq
CwYO3SA4rd33PactvLGzGaKAgqfDVy8bWy5ucqQsfOacKAQ4SgothmGadZwma+rg
T+j9Nw4nrO0PR1cSIfAqoiZmom01qgChEeMPn/0pbDCuSpNRferSMzrpXmljo7Ta
QB+HXBdvcRgtxWQxSNu/XKaE7bW0sA7Npw19Ee+sbKgW8kCX/DgSG8c6fNZFsDUE
H/3dTm526gIVUA5tVP5MG944FG5OcJk7fR6HoWD2aCRZ5GHtJUZlkGcW/0vNTyre
nz/tu3vrffo+b7AdJmw2EzE1U2mphhC0A3tyhwvJmVBOn/Gbsz3nOQUTF/QcBVqd
v4zw3KAqO+DThxU+kZ45ThCWKQG4bczDFYuLlOwWidk7/bx1gyrqTSAr88EKzWGQ
G3KXbFH67L+aa8pPww6kziKnt6EUuAUWGykf4m0gtAElb4jAip6tDM8NgC24O5Xl
zVCuB5NEuK3wTilyxTpkmoxUoHyPeuoMH/fzyFI+HY1LRf8fMqVoZHjTDMzKPM99
e3tzKj0Nrjh6QHi7gAHrDPlyIeFp4cLcHYAQw8oWMiPBc5Pv4sCRGkyhPCTK2z3K
czAit8vw+D7u4wNebV83Bcm8nqQ0I1LRQXms/M6bSV4roNq3kdfitqMDo2zFodJN
l5WW3/zLQgt0hxodOM0zpklbP6sFCGtqvbhBBPWDs2L4i75FUoU5b4D4o3ukBXlU
KHbl9EZGXy99ZIuaznQYmavUb4xYWe2p3+BGA/0A4HZNyTZ2cLbOnk9XNqyiMA5V
5+1RFpQJJ6h+r/QuAeP4YKziweNZ5htcTNAAgUC39Y1Jxr1AObcI0uD715RwLwVW
qphb0tTaQdgkV7GW1XzPpbcs2rg3EheIhDau5FsOKZVY4R6PgBi+qY3mbSHEMcKP
EMzbX7K0BxOw5YLG0JkcUz+HZR3Wq8t6tOOPwqi65ol2NIp2CUthQT/zlQ6WDCP7
/BfmUBLeWaZe+ZkAd2LS5hPzy9xAq6gujquTm5QquzQbrsUH5qyJmCn2TjT4dW8g
P1acy8HlZ7b9WMopcKfNPQGcQDoWwF9gQZdYveexh1YeYBIGj7Iuufl21ZA4YxVe
eTfcK8F1Xv+dQ9utN7FoQC8p8ktv2O9uzHSvwU8e7g+Z7iyV0mHI7z7qe4YPoFe5
xgggu9FqpoP9wq21nKuS1H/UYjyM/gbJpTdNXkxTKil/aHkzDkD20KLQ2K+I3ImT
jvkhT+4IAnTyj9kmymRz+VR33K+AOJKKhbPuqwPWTPHkUWLIZSkuCAEz6wLDeGj9
6p/KcSb0beiVBkepQN9n31bffxtXutoIrLW55DkjstMf2Njaic4kSmR+jf+xXonu
pkEvnQgSsplatqWw6WZZNiZyQR+9o6riMD6ELlF9OGlz+2a9kmWLkkr07sSfAMeu
UW1RJss2gEetabUrKYzQfV8XSaP2+tGWebxeYf857TBHGexbmMPTkLsyYWOvRUjN
mKWF6g2nKzVTgSAN+aeyZZSYFtOmhKGt0lYNp6ExEx9GV54afoXWnDFXfzKNs8wz
l5h4caAosn4GEr4hyKy2wbGlcKCHfAZFkpZnLwdn4Gq1MOgnqcBIq5j7+Fz0AnCX
w1lwGV8MUdNoPOALacd21w8gQQHtU6jBN+9CQHaRB/24r3NZaD8JetdTgqLd2bRp
IfBAM8etdTIjpeH/GQSls7/g6v6INLDkdsjIXWuXH7Gx7ery8S2gSLwzO8ufy5q2
32MDzMMWBbqqxLvVz8W5VSj19ABT3jAHh2ZzY8wCywN2gvSoiouBIn4ksh99yT8y
ytj21XDUpHRiGXzr8vJ3svH/hacoMpCEOJgIfChb87DQpI7fkeyYaw2APYSb0B+T
1FDOzsMWHExsxN+dhyFXsOH1UqB6hZsOLMOZu3vJYc+tborT7jS/2a8sveppVypC
fJXT3618WpVOLjDFOxW54F/U4/GIyFg8XxvkbT5rIWM1tx9b/Zfex0pwI9dnd+4g
efJp4VWPj3FEmVrkwDrm94GtgvF8nQ9WjBGX7j5uuPVYeHGs30xPIyMV08We3WnJ
RBcR7stWP36puIrArdAqiqmu0mPVMydIokd+Kx6J/L/+vw00SwTo9KkhWmqd2/ja
QDLMKIPjdzPoWImwPob8VDtC/XFixFnZCuT7ilJaLZjapiVX5ICh2amD4tF59jz6
lhySkVszJcmrBunewbeIl5gioIZQmGVh5pC/vX4Q2bXpTptVFr2odRBBktPz4l5j
pJnlk8UvcjwgEgxgg0+bDKFGfndip6HVLedelAo33NTBAH6bbMxaq4FZZa4/Rh4i
41zBD07hAduHxollxpouaPiLiZ2RENaVJNTxDypCwxf4cA30JdNPeGmtW/iCS0pG
lZ+b0iszBG272RynGeCkMIwYKU7WNL8ICS6TAurcsMy5FCIlkE/zte688UKK9DMD
VNXiGAsCaiAQy23mWIB50/rpPJbAjnnr37FHJvolZa4KIdNBSsEr2m9gkRNzN6Ik
X81SDPMN2j0tnZCK9D3fUpIkTWHQ5Q7fUvcM9zOd7n5Jj/kFHFYKX75vVi1phcmj
Zd55m4229MJ/AeE7JnTmiH2yCFuJ6WDQe3MqRPeleZD67XDpYMgejF/tF3lZr+aU
xbEO9uyPU9LA7vcAM1IJS7IcDqQZevMBqTQVtXp3vcfUnoFnAm8edX8YGujW4NEa
8Za6S/lOncn/dAbadl3gvsvvtEQUe5wpfMJd3HMo6dDnFzaR+bOZvHaQSeQ9UzRa
goNa+9tP54udkTbZXLlNPPiZSVsklCEleV5SnLbZjEwgI3s+9oT2fBrY9ZBv4FGM
hftW0oEath3KEiw8XuqU1Bp+f32d2bNiPYd7R+sPYfhf+fQpc+TrW4iu6u/UDAQt
N8gKzp7ZQY0VsUtSaqdlXcZtl1ceEcYvEUmZ5BN2kp7sASlTYEQ3hg2C2Ig9ec4n
uwtpLbQZDKVF16DS98BA+u20Woq/03d0egt3M9AMJPmRZxJhFXpIlhaeinvsld3t
1DMUtBxkLORlU4eoK6fnBWF9Y2m4wjAf+GvHwUQubzegc1chtcWGHQU8ssIisxYA
WwmTBftsJXCJP0Zt/cDlQsx6cPvuRd7tJEEYB21zYMzHPhUyjyIHjvuAUVh1qsbQ
/IYxjxhXGSqV2oRDcXp7KBU5VUUJHi/BpQFmxkByvXyW6Xrm1s6O0cqySFms19Bf
zo8f7v9DfoYdFDVZxqDruTqbO31rz76pRAeNPIoJFPfUVuXK6K3AOL73SxCh3IkD
nRLhJS9ENyy8T9rJJIcR1y9FJiRwtEGGJN4szIK81DzBJlTLKviEFZDYDcZW9uPp
OO7ubpLY9dDL3Q0fwR2mTe5K3ausrbybPqjRPvCdBE0oWvP1TX8E1JLK7R+A30r0
7M85vdoEjQjjMf8PIwqAzi2QDTkMrB9r9WBOLOh1wcwLunNNnZl2Qe2Ei6HCbJyU
a166MhKBOliXAIgF3WBt5xhwM0V0Niz92naYh0RxeYroxtbVHiQ+StjPQ1HRG+vN
loXTLvmJ4zpnQ8R8K8Rc3rlEC3FQHPpYPmnzML1uHost9Dnp9akr9ADjl+qNEJHr
T6chicoQmIU5AHCkd+vLwQayixkGx/02GMLBLFjdyXmIO4HToAj4tZv5qaYhIkjj
OkIVyHOjQHAe1BgzhK4cQFVok3lvIjcgjHxXkVuptUkCWcDuVj39EVh4EUX6QXCD
sGjN6R6o9OuIq/46EVdE67aDrD6KMT1ZTi4AepZfjtNdRt0pqUScIneybkaQ+px6
a7nqFIYhkxMJOUf5JaYre9o+WpEmU6Qjzd2y9tMfI6eOlKje3kBgBH+lDz7CPQwA
3Kk3405ZATwWF0TDc4mvtv8VqcZP/ZlyeewhG9VohOHwXww32mHcH0glXzIrHWio
mnlPJndtuYqZ6lN6gW1aCLW/GmYkWWVOU/b1i3i7yUUY0uN8BzvmEMyx3mT7AIVw
khVjAR1718anP9lquElMwhonTUmGU0WovotcsaXc3/Jkqp+GA6cFiFu52V7BoEt8
tc4SaGgSlyUxJsLP3XUnuSjd7EmDfk0f/ilrWd7DSEFSq/jyhavRU7zr36KIKe0k
ycMJ7nU3sfYsXWhCUURrBCDYA+o+v7RJBN+HztRMRqOP7HVLSGddJH+lhchRtLrP
UnOMUQQ9/w7foRhZbrHtJgIoRw4NtxQOxDm/n1h/G9qJE+UBYtgta3wsYz6UkKrD
vQOXCS6lDEaVcW8KEx6vdY2AJHjhZQR+GbNaSHmZ341XajoBEvyuW/O/VAV/o7mU
TiXHk2vZxx6NEMxGWj2ZU0BqYRHl2WhlkmJ+WXzzWDGDfArns4sULErzTLuw72Jd
BWjS21aOWfdCq7kdcHmadVrSEia5Zq7XT6ExYY8wEpOaazt7jxXsSb2TEez1FovS
0mkYXgC99+SCUD6UXBIJDrTUL94xBsn39h/lMcuiIY98buQggkkJsEwJKU2256Dv
ktAP74FQtbYi/y2gtK8xo3YfttyFO9ZtTRvbDagXIsHB8hTkLathTuvQDK5/85De
UPrLkdQ9MhbI8Wjs2jqdPugyCEmmhh9JZhGZTWhfs+78V1/cwCpARaYzMVxieBxi
fS0r5kgaITRbAdYlrWrWvglQf7/IhbwexLGZpkbj/vGGLVLznglBoAYrers2I1kq
NzM+eP1Hh5I50wUK7Z0F6Btd9pIzKMl462gvFux/xQ4a0dosztfZe2s3vqvmchLe
UteSGfgNjUKL93b40pvZb0x1d2YtezoZhYYTlnE/Maujd8hKlrpgBEJVwdyjb12I
ywpUYOJjb8ZZ5+ei0zOg/l57sLwDTvxuW7z41l82t3gYI0k6CLLP7/0W70bNn1QQ
Xjy8qNPP5usSJKLtLmEhMedxzxkcbwYm3X+EZ71sgXDRc1X/loIfh2bqjTYqIYqb
VKyjvN/DJsOUBJkZNE1/OU3TsKMP6xuIwTIsb8Q0ftoxcVinu97pzvTGxDu1M4f9
kB9DRyEDqJm8TjzYZ7hQnixQf1h/bUskSwMExgHYlbuOED7WPQojDOxRyJhUBYom
PgwlUnGLQenHr/64SQ7HC5k9NOTxUB9Y9yTQki0OHqCFKMPECnMYHIYs1zsEZEvS
AuP3VhCXlSKdSA8ikXuiEBWkzhmKwPZBaCT1P/yFceGTQ0MeIvOfKOAzKjN2sa1o
dbZO37klrg1r4mqweUdJny2Gd66x3bFo1fLu0U0/C7Fh/j47LjIr88yCsoo8dCmM
BxieKlOCl/0E+UQKuCQyWIHUtxrA+pEZzF3LWkGBl81hMdMnwDTjkrioYaBka9DM
rnpjrYPpQGMrwu8oQYS7mFNLNKxs0dxpTOWu45pQ+BfTdgVAH7key1kvxysWIDtN
3zRuFYRhHO4fROt4SxuOtZMb5tGX1hTfK3vyf2uAFaK0Vn346Rv0lbLBz1tqnrS+
mTRbNAm9H10qN2zMg7DNivFfJ1X5JX4ZR0LxzunAwOhyCGfNWCMiyDIEVXupw2OE
2NUx0IkivIIVmouLCi4dUgXQalWmUJfdRdf6CuM4LoR2ID5R+vYk12gnidjqB4xo
ErqIqoqgly7FMsp+WXx+1U/+EMHfDut4ihWCjhCLXown9ITTkQdhZoRujxdIW40B
fQ/NMAMyXmBR/ZBb558gVZrFXIy5ZhipVY/WL3rm+BSw0+T/kGKEXdEb1/K+xABe
OUZIe+FgfwKeS79OyEpCH8JI+GDZopOYSXr3/XJ5S4wdIex76eB36838SKBUKKfg
KPjXEc0QyWb4UUM8MXM4Zl5QH5F0r1tj/xHd24KeQCsTYD4j9YQ+CFrMEIEP0Llt
2X+arFYQxRYUQUa8CEhwhJqDgrZ6GdI50nzQzEkHLaXF6Uv4iMB0ONaeV0QZd383
92mUDrXwJDgSclADjy5uwWKpBEN4nPxy009eyN+Ny7mJUpn//dV1o5L/Auo4isxG
1R+cW/YapeaUsj9D1MheWyk0VrO4FTTwl0yLVoOCYOywqg4hVxDbwq+Kckjzw9u7
LRlpL+CxVBl1EVo1XxGlAqgJhv2oBNACnRFwQsDWEYCmwXc++kWNeqpKXnGyZ+uZ
OpuPbJrJC2VMkoJ/SCjq17ieOthKooPx2mIBzAOkvbk9plVyy3T0+Kx8OsrKhRNA
dGKgSrPvREYUinmIoiqdZxD/QzZYcABoo9c9syTPSNg0IvFq+NFwnGi6QRwX4X8T
ZSIaZmWThLY63PlASURotP6FEde7P3QygEZ0/7lRN0rlTAec/lQNE3EeRNmHxeFZ
NYUUPMsUPUsSpj3+X+dM6GXLm8DJDZYczl3ZrLiJ7bW2WlyUNPFixmBNfeoRbc4d
wifPiZ48RTsDPM8r8/+M/YHHo68cfpkqKRWDtIjXSU4Xlkr9UeX7qtNaBgPDXsMd
M08FpA/YSp0TTLpLNDurVINavtzRSJHr6D8HT+IzTYB4yO/s2GPGN2r1gBluF7Y8
0Ah3WqJBolnITW2ryfluNWVWphQOjomdHgiYl/FuWB2TvpwdjBY4yPuPfrlIq8gi
yh1lXj4r5jn4UPIxAJCabCVaAN68g/fS9P/DkeyfipLyxE1MD1bpqxZ55+vEb+kf
hV2lSATjK5I20E2GdRDzYch2h6mPUsiYuBqMnmpXeeA98Cswew72vePLNJq4NbZN
+5YS9sFoC9Co4OkGvZ9zTF6slY+ZyodNMraZ9UmilHiG1Cx7VNK50vv/3xS5EeEz
JnmLzNttWt1k3bpPQzgiAeGm3wqy7+t1btfYxFI4amJeTLHPXo5ijDN6xVx1Rd5z
AAGEPhV66V7tMkNau5RcDXzgk83qblWqq8Bp0RiH47T3tfy51xOr8I0gIlKX3Roq
FUJYi3MMJmPs57rxMLQm48xWOP4VNRtu6jR3KXQVXU5hrbBidi1U+aEVBkU8b2+5
xu13FNmw32WJy+oJO5GB0qxpYeTeWjUZZExFHeZ3ea47VUjK11Nr8x6lMU6vc+HE
a3G2zEHUYM1PSm1afCIZCNlAVgFCeRlV46URnHb8xOTaLM2Ih4Lg6tceIPHy44WD
nkhciMuro0M0VrZyuFLFciHcE2R7TbEAttCkKxGUu3xfwK6UAbxiBrakYZ7FJ0H4
oqarkapeJ72Mh7jlgFqbqjpsOaV+pin2oVUhMjbJVyHZjE6qEvHAqsMaXJ788uv+
qOecZ3iraR5qP6V5X2561mCDR40BcwGJohrsP//NNXUQDPyvdkeYb+4IpsOeKgDh
hUEntxpFYPW0OUBPKO06V0nwm6oa6Hpku1KHN5fLsFks/R4qLdB0nZVIeZRlLZ4H
T02W/ZmJuZJkAqqV1701GE6EvJViQz1GZcLpMighTcjtd+AnrxZHtVEeaQWWxl3t
nToC8/jySCHS9vx9vHhf5qMFmf9pohbyvR1FL3YYBZPkI9hFjiYgosI6mu9A8nCy
zzv4KzvCIjDo23DNTfKJf0QJrJLCW+0MTXzXt0t93UlzDbyDj8s8XwSFc9rKvt34
WCcJ3Wcg3avCXlKyZ0LAfZ3d5/RbMxd8mXO0j/qJwB8ZBxetZRfa8x4+TUmWkIVc
DlNR7yz2LL8YH00RiltpLFLGvS6F22R+PuWqwuVtuXjT7eeM0fla7SQeWYTBhHhi
/l7bpPjcUIZ9FJGUu7JCvlBJB88wzzKGFXU8WvjaQGOV/tV7cOODGJM4GPfhxQi0
Hvw45MYaGa3KejAVnf7KxJhQnOLJEEo9IEYKwOebY0LZMOL8yj5LM4eN290aMoex
B5urIplP7ziaBQJx1/YjbfnQRy4zdZAa4zVTWFvcQ+YMyP4rvXFGxQXVvjIO/gAm
lhMjTBHdvlI8bviTi+Muz5gvqg3qUNlqIPSLzqhUVQxf6EIjJWboaf0f+bJj+SN/
OhuAfM+As1mdauM3rzt0t2B+eyKjCywLw/Q8QGza0QDEsDXop7EgBgX+PSX09glH
FkdTLTz26xGIieAlpJ3Yfp5XiQNKq8X8Mlga8cgJDz2sUQlGchMu/f4+5heJlzm5
8IHzxfYwmBKFPXWqlvI2arEO43ECoojex1hqEilv7VLLouxjJTf6jOzog+l+jKvM
t9fKa1IIj69RGqZlIx2dtIYgpUxDCiDLpfS8sQz9XlHCWnCndC/ERzRgYGYL4j3W
2MEb/B1nxkMDffigX72JuZIocdYuNgW30DF5RaBQej7PwbJfY2dqhihG9LtqcH/S
0bjxIT1uEusJluwVhgNMwHioVJg/h9qYf+0j4sJo2r5dOC+A4mIX2Mp4Fd/ADfvC
w6eJD5ZfMD5NRagKm/ytzWmrEXRAgCDxbC6SdGhD6GbIybQZIuUneLnbVmtu3Bke
8fSXVzyrZEMFxvNYCq3OEKf8IrsLhxmpPeYEbzQ4rJpu4uJvzH+lnxihe8+o6Jcu
BZYUaK2rfQYclbJZ8AOXgfkGEIorsfSmyARCp4JxTUx3vnedMVKW7+8SmqwK3bpo
OhNVigSvEQ4dfkUAIFvwAE8rwdimOQmrn5PsG4hcd/ozcfGMgSX7I7WeZi2ZB/Br
2SvbMxO51EitBcbAQMJ0u1JCVKS+8mGDKOndeC36LZIsbyXCsW/La4FLIiCzvyMZ
2/D/0yR5OcdsV5FEzJ9kKPQORs/LiLdi0dYHooz4LdZ8dl8EIGVx4+3iNtWgREwI
Gg8h1GCPQTl7HlJyDL31BwbvP/k8ozdNB9OMjCMVZL1tcEs624ZaC/9hRgQG8Py3
6nzBX+n7KVf814dZ4gZ0GA5G7gB5YXW9UXI6y49NkpgYHCB6lJEubnzoGgN5zmCm
QfkyiDzv1EUcSQyzw29/xqErf/1omX4N1d6GIfAh1CYlSoTn1bTXAa8nbUbz11TT
u/kMqNqXtQPiE0GnsXwDqPxpNXF4BMHp7ivB6FlMInk6pmwRjYAUhnFouiNkCaxi
GRmnpivDriPyqkMtq3OnHzY+tqiwDr02ZXJLe+IDFv9TIlZlC8hEocNrJPl2A5Oe
+HAv6iB17ZGgos8tzRliKehfvHq6gtEaK1G5bGiZBRCURZqmx9sVfSQyTASbqLB8
7rw7u+3vCOCR/qxbqd/wwLlYLadSoR64jG6DRkoFdawXgRHjD2Kf16fcb25c1v9W
FLHTbsco7tDgKDVyNgHPiileWGKzqyeeLeIrYfKDy7ccebx09gGMOUuqHnyCeJ6I
4cD++cexzv+iuyv9DW6baeYh9VzWUrmcJEmEaRXD4vD/rldWoXEbiW0Cff/DGiYX
SIjR6+zWgkBvUBoBvUTMGReEF+asPzhR9qAg4TxlZwVCCDEwxqjBQNZ7l1Ko9Wpu
efIAamm56xLmh45PsmPpPpuYluJQN8Vigr1kd5xprx5UT4Lr8a5FVL/mPeS+kyp0
mPh6HbzGgihyyPy5TwTvD8xTg/FIgbXUzaPyk9uHuufV8Enaq81S6PQwGAErR5SS
PaggCbjVVdMAvNjpWONK/TiiA6D/gez9ybH8bgsuD9EgIHD7v7JfTMMsXZRWJhOx
A+KrSJWUFLml4Mzf11JE8vVWu5rk/wR/lUOpUFGNrinM4gmFjbqiLwr3hc56x/bZ
/ZaeQYkb29DtWl0EQofXG+3xpYhmtWfEJ1KZFX6Hf1ZCwNguEg0c/YDAtwxnANUu
RXXuouZBmtkpM9ta1k4mrVeFMXxaKINv/NRNidy1y+Zd6aBbXygxBGPXs921SdUq
nvkvp8rcJlxGIH9ntSvYI+FV7nNuoVtGQASvBa5vMglNJ5kvT3oA5EvIklT3ZRnS
7lODtuxcRm1UOxboRJEDcrr6P3JsBBNQFrqzjod2qGQue0YzCVuRxVdZTmt+bL+v
Y1+SXCFqXzeDY02I9332PeIlzyzGmrkROTqOto/bpqjcECsym/L0gOR/u7qs0Cfd
5HlAVx4efuueLwA7Banhj72eyWLA9JcKZmROTYS2SbcE6sDZGcwwtSAvgftGzrv1
eK79WLMOjbtYWjB8oVKS/9KTL+EED0BUswA4Kq/qm8lf6vVWAqVI7eltfg9K0Z5L
b/CZGnBatgrSeoNWcpqpS0uaBy5FektAC9F0CCzEzkooxnBnQ33LYSmoY+w80Naa
znJk8qptCDC0Ob9tj5wbPaf4LUl7ysMuVz6JD1yaKn+K58OcI8W4uYqlpqjnHVYx
jf5AELtDGPxIfjn5pmflo8vI5s3lQpizoiUVIFkagC0zJwdhnsrZ6yna18jaO241
/iCrwGuiigIOEvZtRZA0L8V8lrtTdLUIE9txn3A5v8FkcYrftgQQ+J0pjz4UHS1m
JGOKj92rYwxpWJKG/Ah58/zCCUJkZHLjRVWYZ3YNee/c3lANd99BntQ6ydg7/5gj
ugbhdACuGQJtR9iGPAKrZT24fLrqtoxp/VgJxGsLxCwxLtjgXt7LP6eY+xgcp5JT
9Y694xRZSUXgHlsIxjWK4jBbxFIpJaxXHApFl+7W9l5pBV9wLeTevk5kdy7BfYBX
mwI3D9+UdrNHhjar2oJnXGf/CkOTarb3cJsJFuGYfm7jPK+09NWmAb7ZQDJ5eUTp
u3SE1LI69zWaZQA1tLeeSI2jm8IuQ2UlNu31qCvxspU5MRrBoR6BMMeXz+Oa6Xv6
RWfdSn0V9kePbXRFjoEj4wppw+5yExesZ16XpJhho5cn3NrrEbr3zQJuifTXp2LK
N4aUozHdsgWcpockbQ/PHnPf6ay7rUoY/G6v++x3OZme+Zz3c9JRVZwj0W9J7gT5
cVUOWGl7KffAjjsVxQ9uNsEQJBRRioKGrPKJ5zPCN2p1NRKWWqrxLsnRCSHQQJs+
rp4gdGh+Ti4bUkcDOuWienMXOlsMLvktUDyHQ7oRQuqSS/vb7xFMfqy3bq8OSE2C
FNslKdEuZXFpWKh2zU5aute0bSHIiHMX5SJ0JjoKNvvEXVAvxIjBNrjd2q40oHn+
NZTd7sxyJgwBjbZbZVtCvzE6hz5ZIiBu6c5RjTOfQB/KARX0RXSI+JNopi+wShDQ
eZIFr/yp4wsGNY+YC6WGZfzuyfGCIdIJcwQ6XEGuQ9s1LbFWF2dAv4uDpCytWdv1
0PAeyiE3ATa66Y4TOhq2cgEFnGBHSYGLOrn0ObqEojHvAa90ScWQV3n4j53jRcH6
lHp7i2JNRXpkFNxp4nm6ULbruGHJwFuET4eqaXHQzrR6dtIIKaWB7VcM2j4nyUpJ
xLxF1SYS8K3o9CE4Kn7NXpHIPsOegROV4+mjlOnoYFM89Y8xt4gxX7hEdskdn2br
aFlpZ9QCrAw6462jiEZKHXL0qddhmZOb8N42f836UD3TUj3kpV0P/SeGYmNeAbzt
wXJKK51znXHqgS2JV2v0pcU8lx9rPTxzZscvwjQj2STON/xJVcnqhyr7K5BJ8iny
B28zDV+QyrPCIXjIJ5n0KqRvmDGT4jzZKJaETaHFO73uW1LO9AbknxBmnehpgScU
Llom5ntMPG0X6WuY5nFXK3wB1/UDijZwYTn6xz4mgnJvTKfztxdXmCawR1zoGKm6
mfgHkXCmVQ9QdZjnEk7GMPP1zvsTfOzdvu3/VfrF/mwUQAD/IOsQvvD9z57iCcJk
/FCO0T8DBrPKKURRoEk2bH6Q8ks8cx4z1ICOspdD5t8wzFtzFN3x4+ZFmNRmCSNG
ENNNDki6OX+MuI1CdZZkmcyjcT63lzknVlnsY3H87Dz+RkeC9yDfXutUqCklc+HL
vL9hpkn0CGQ23TsMOK5tfWzHx9QODbVsS7aveCW7UwNnsEI5dysr/oz/zypeROEy
ZoJVSZ5cyR1iasNQlAPtGTG+CYtB1HsoqA6dR9DlZ7zZHRVcOUxGauPZlYRj0XXW
GFW8/u/4W1QTWbYl7F3AQCLynbCAmNcU/0mKyJ57FTQiwv1eyFkaUaolCBtgCMlj
8hy4rNlCcbAOtE1RmPvOT8IveTt42gPMla9GjTgxUktitvG9AT0joQpYDdWGfDUp
PAR/KtFeFrx6bdVSNt42yqyuTifHNkdwPkaTBvJHh05QFgY05QOyOwCCqcqwT4rD
uFQ8LZpH/Mk75ePxnelF3HQ6qQyJkNObBuDnh22JaGGr2Z0cQmmLNJg4UrRlTev3
gmTqlFGD8J+3vcLwV/xpv6wSGteQYhLX+UgensaHJtWZ+fPn3vDjxoF4LvqCBzLW
2fl4QtkFdZa5lirURTJUoW13lBA7kUwHsRouD3Qoykf6OgtbKUwhs3d4+An3mW/c
VA3O+G0GBZhIC+xfGMUPdmIc/49c0wJyk61cJBvfXjiMkiztC+fgn3rMCb4PkYbM
2Wq1AjR8DPIpDKmyI8sHp0frx7wwwinD9tTb8khqe0kGzzv5nupgUN+cKLgmrNnN
2+RxU1eKVHu24kIqc1KKoX9HpjSAVBhyoVTHjZlDOHvAZbd0SshnJ0M3hbhwYNZi
NweF/4sQXl2ZVhcvi1MirDFszgODVjkx7WF17arr0GuSyx97QNZCnkq68OPJmNik
qJ/Beqwk9Xrgegn5myECFwU6i53WyYrFsWfNSpIqYRXKTWm8Rpkjl2PMS5y5gvIv
u+XuXdKQJSO+S0IYrOiJVinAAxbXF3uJi1Yqm3k43fQCMmVZdNYK0j55NkDpoQoK
DHJZ8zeGFnRXqV36p6E89YFqaMLpRuvccDsqfHKGe8lbZ97dbAnq0So+BEBgAtVu
Qe0V3MttyKMhph6oxixrQALmskylb5XvuVjqIXxAC4q2SQMeuWyowmM6Euc2/rXa
VEyo4GgUsLzoRhG6SuBNSptM2KlZl65N4msB/qPcjfiOT23MuQNlrT9s1QCH2Waq
DSm9SO8LhW6jhzqHMIOotD7U/br7fcEq77tO+d9yw0MXmL4uDtyGYwevVc3Xa9NY
fFg3AqecWQZ+/EjGrMMa8FMK5ecq3xVk0v3Le4M1BJSovP5/BWTGWCcT432bQY9O
siTSWgbsZVUFgpVzcL1hKpxS45kK1HZ/bmkB99OnJduj7tWIJebDU3ncN21B6nA8
CR6s2UFoXLq+aS5FjAfKrYxfTfPcy5nTbFmFkn5jESmeApVDgj7FlMvTjSaB1UhO
8XYWTOHyqHqkik1NdvR2hKwQ7ETHZjQUdfav8WdVjx4p0EE38R2H128NNxibSvFF
cLhJz1HVsH9MdfuRPaaOj17B9P1zHllQN645zx5yNc/Q7MDaxVU4z5LqmesfwhfQ
5RUfg0B/8DDfEX548itmeB3wElFv249a6Vk3u6bVZxiTLeI2cLdmDz7cOjHmZGs5
91eNchJq8EjKkfejPyPdejcpnWNnQ6/FvXwoqLeuH3xCNXJj5Z5l71WkQ/ZuLMo7
hmjipiOtnaHaWGmwHEUGTlEzaGWhbkCo18Z6ZceBDw2vBALF2oxPJP+v50YgX1ml
5mzsLGRJeS6EX7wD+LwP9r6rt0BNYIgwLI2JmbDQSWnWtZ5E5031Jatdyc3O2MUL
ythbuYF5yO2wnem604yRn00b9X1a5XcpL7JHqGZtRAXRXB2E0r9EcjjNcwP1UzrX
DWNJbkl/Io2q1tTm4q6eFYeDT7hNBq4mueDAsFQ6lEFa398gLJYUlVEQij8TVJmF
+y6qYEe9ltI3UdMUNt9Ad1WBm3D4BS9rm9qI16rGh5MBvMFDy6//KauuRND+ugUf
gfDFazOy+PlLcxzess73SMY9WFybOABdp3Rfg+X6yghephtA689YecSVgA8eI+fz
0/GSnSGIjrUTpqBTMDzg8J9SFBskHI7KLkyqM/ZaxBD5J2A2NVEqImX2XhXzCt+t
jEAYlc0J/e89I/ofxo4/zvJxPmzWY9r5Q+paqEJxtwu1sJqr89YRUFPMuu2YSWVL
992oS3z3Y9sZ3+tKEhg74+kIUcECIhIAgd+0w/ItGijS7xNO+fXu4Y5BG9+mLQEk
ne5rYthhsP715ZYRUATrvncsi/XsOtGEt74ZfofoNupHGRoGHz5xqB/KyYxNEa/n
3+aXatkz2mCdM9VeCcUiYR8WZDyzq7Aqq32xaD4UPX+pRta4mV6srsC7ZZRBcs0H
LKv83Ly5qncBv9oCeIJSw5ER3iVCrhJs4QN1PE44CHncmPH/VnlxeY36Y1qAJQky
2s5i4JSa0yivdaP1f7ef3racK0+0t+PUrBxPrOdGJXDpOAXcjlh6We7/oRHDa8Mq
Gx/6MI0JWLVLXpFGuEOzYxk9TvOMQENsxAttOu0MqSPk8s0pGLXphqjD5wlrNlXf
+DzyQ+F1eV9ooV1KKAWqQbPfrIKTra+YaTjQ0kZoWQUavMR4pEsIZzbUgYu07pQZ
kTd5DEdZdP6kMEMuer9/i+mlJ3K+G4PhBY26XFbnuoaMkyNT4+BEfw9fWZHGqKG7
lZRsDmJouhDdRIEyCVpN14BidT4fSmG725tFtere8a+ovP1sb+V7zH9JrFS2xxCn
MY8OYbHLe59EKOkNOMQHUi8uk9sbO1IiAcOCOEcfPcLf2G2v5yHVi9HuXkcz4oyZ
HVk5ijW7+ZmwKRHGBtfLCjZEZF5eb9IwnCTxn1Vuhg41bPjPx788aUB6n9LUhjZp
ESJp3nOPXEWu92Obhgm0h53cPRmPo3uqHVIUtPrlKw6pf4PCc6o6k6OLM46Hnc1O
LVWSDOleY7JSXA2yIWiyB6DFvovJlbxtYIY1eKSCLt5CwP3TKk+CnYIZDDUApJqa
JxA+dHO6qFm/sM49bFruu/jX6gm+BKDPFmZOp0EEf4wyEQJ1PlwOShGnIvgl3wYU
jyMY5D/WPZug5qR+Iv5W19TizudKU5lrgMxnWpTsQUae5Dv2Yw7+mxaKS/1GtyMh
ySwNwU/SjLHrLcFn/yLxE5CpQPzeEXmEH0VN07g+pkV1k2zGghaA3R4rmZZSdOGA
i4pV5BljN2knwojqE0hjT+icjfZF8fvzwvMgMDC053dTZ/rkyB1qzTnxmtEZwHdx
TmTmzNlN2WxRCMOQqOg3GDgdbGmYRblhrX8Gh4ruSJnPCBUG0frlbikf64wK6Y9X
rfbYbeXVlcxq3R9f7Wj9HHOLujYt2wtfBwK6p7x0IJEToW/eMGHTXBT+3lRDJswC
EfKiR0m2pg45NrjvERrKvSQDEdDWVXv596WJdv8WWouS/1cEQtW52PxCQtu/0BdC
Mtf78dR8OK6XryelJSP1se4YKw5OKo/AqDk8luwWUSZWMnXUp6HoysxAv9qm38KF
U0i6Hoahwl2cPQaDtyj5oqqVyEC+adFGszawpFR3SMuJNPK190xgDk+TC6eTBm/M
7GC6LSHHKjr9R9prPXAQ3/T70lReOAZ7AIRuBdSMALf0RhP2GQZpBRaWVLdfbnnF
2Sm0n7gswV6IF2YhdkVX3ZXD/ZZck47yxfO8ZsakdP6dR2gWoDQGICKD8X/kXwtn
ARydi/ta70K2VuuStOzTg0EkP078BvDZKLGzW4YwOOjOGbsbr9fAhNAT59Xf4l4E
l/z5hr2GFfV9pxfRcEMskusCTNluUS+UfeGA9bADkuU2DiNyj4tblatR/O4IP3+D
8ORE8pfrLaTc7LD32033jdieMCQ+HglHKRqt0bJaBJVMtJQzPENV8Py5Yi09EDuU
JmVDk7K1VkDhyjuBGfbnX5o5/et8MccTo0Vy74XXt3glRHeRR7MRtqMNRFb2/yeu
sqtyo9rtjM1b497rjpWD14O2Pv1MKkxeSrW2Axl1SQKTXeC/xdszC6gWhJoU6BEi
ff+iAHfKyl5YCgIc19gl9Lwnw6KRtqzesxKb7whdihAa/XD3WfnulYUfCW19j26m
rr5TT++aTiD+blrBC/g8moLiaEB+gykX1eGQ28IevVtqY5fLXTl8dii16oEXIc4v
ucJIwj2RbhF+1sQh3BaYxARDhiGp2agLfai7KC1hgBtYHt6P1KNFbmKXJhjgvyQr
bxcEUJlD7hTAbOfU3MvLZKLkv3SV8Nj8nGvTiywgXD07UXnw/T1QGP9xzzqZ0XC7
mJOUBP23/hUnpL5MSBis/ZnWWWmHN4WcAQdHYAsOh19c9F7+7rFw4Ah0G+mbtUh/
UZ2xE/5qGA4dGzx1upPm1D712sMIANFl2zyvlI/O5KUPNHXdGWns/e+GMFixtXTP
qw4pzWZItf4f/+hHOiHfYS+AXh+fbE2IlOVbB35bMQ4Ir1/z6bCe+qD+JDRuFHJB
PkSS2Utde08qSdAOILFwY+WT+H8BsEnHvYuBoEIP7M/vzu8CvCHNSYBAMWNodw+v
4Eesu/dMTRSuId2A3JV+OjWl/xOir4zVJi4udAQ/g7G4EVh/qs+2oneG7rzYsPfL
hqItySGpe+ny4mlC62X8tzwfJA+QF2qBP0JIgLqeurtnZKTtDHOk73XDwp3zFJ+u
4OgoVUc4YUWvNVu8ZB05eUccSyWOFmzdsMvJAaUF86eY1HdQjdY5TpiZngOh5QTy
dp3Mwjd7piqwF0fNQSRimXVPvO/y7NZbxjK5pydU5AfS+OuoYJPZESF1QDfXM9vR
baF+qVpa6d991qrGhSBuca81xjfvEPVv4l2TsT3TfXZXQXzDNRMbSf27fmQERgLu
LPqtDXmbW3fymLzx8o2IWyfWXbapapaBDK16Xk31Htdx55RSr0x0YuiV8TSKADf1
ntfVJunqq26hmuoLarL//RqWVZAxGFFs1NzvfW/IWW/fqCsxabPF8LiihOJ5TZz3
ubIPwmKbQLJgTKha64rDt2I+HeopqC6tuyJFuw6TO/0AEkPUKfUnrmTaU9Qyy8Ye
IZuzOSwZCPuTtxbkc4OBjEO8U0WTveZ23eBVodO654V/2NXeyZd7/ASc4D4yEUdA
CeT5J3w3N2j78If3d1gQIWwiGuqhO/4xCAv0xTdH/h2uEnAr3iWR8q3zXRDM8BCA
ns3y5/Xa63uudiuvep+t+lXdLeYGOvxyOGr3b8ouIFLcIR3DbGIqYn7WQQy9bbSf
+aSTgCtcJU630+CQFvZHmBUdZhmklfNmbZdKO2NK50XOfG8xMSraUmt4hwmhs5Gf
7NZDKND4/6nU5V4b8nTN0bosrwETsGf0EiJmfzhe3C21AfVuf5iLJdThZp9kldUy
wTp1ucTsxR2xo8e2d5jgVGQV1Fdo/Ippsyu8tEcgzUsN/yupT1bCeYqARFGVpZnz
BAOjAvvRQfA3U200WRNS+O+axUKpYD3UWEo3sSxptpnhQdKrmxmZwA0ZFfAWEGQb
2RpUobb7QPgOwE0qfvv4RWbzcEm5gLs49tqlimxlf90R4bv4vGmHQvdqGPTbvktk
aPnlseTGpPBUwdPTOUcZ/C5KhCP+3TmpGD/dBXpl1KQGZtby7eQ1wm4X1sQTfnu5
4KssQ0kvhLIWuCR3OMlpD7kiN+VaJWOB4XpoVm02bfgMPk9P3rGUbIDpCLLuxIJy
imXHOiVM3hZGngUJ7XK7pD9K6eDND03DRn1phmioHQrJBmzx9b/2sLO6HIOWHuJJ
TpROrdq6zdCybKP81nn3+eYCOkdaVZXuLqJNdVD6zZNSQECk7YNNGOVouo8Qk73f
yjQ+rIqBMkBv6NgTU3Ozz/vAWVMqe9y0LW7lQt8DgTZpojAA0tdMoFAEOi0Po2/l
2kY4SIaTILrRebN8uXOlV3QdYowhqDmXfUVj9cM02b0s3F1kMwpx+FrPFc0ckYL0
0b6GjFOLvSp3neBW1GrG0q3KaxYgQ1Z6pYOHdQKILgajrS3FG8PqAUnqUii9tLQx
C+XD94PJ7DiRDJhoWejVKbrLJMJWsoCMCU9sb/OyAIx/IKch6U7A7qEMTOawWzLy
FG023L9VkUGkoOAcyq2P3dJIrpjxz89LlWc/3bkXaz2I8oFmZKLK90+0nN5rMMqd
oDWwoOHo55SUi+BlF5XStPwaA/8phMt92E/e2FjfuQHLAXorV77M8r2bvqTMJuds
ruhLhY2sNFZrqJPi1GTNT3I4jD2QKbw4zNYV536iwUnLD4QJDRJ2oaGimxaLZkJd
TzS4+SsvVbKtMOvHxpG6Atf14Xuv4kmIXjI3KPlkl83GXbKesp1Am88tqP4oFaLl
4dy1o+MTVYYvQntKlzUc2olKO/NJP6+DOObpNSBmh658m0LGo3h8qpCjPVQ/fKNS
sD+lcrq1SW+h6ee/e29WqqWIuj5RxB0aUjoU4L7Q31Drj4S5n6pau70pmj9wKkM8
1DpaEjBCoLKGlery8HUpA32FbY3Gqg8Bx6p/xLu0tmhri35LLzn4M/YnAJIc61Ux
0AvCCxOEvK2JFw6/McQakn+ZR2i5lnT9Wl461/Bo+gCw60LEC9Q5A9WbgSBFhZBD
Vewj7mQm7xSqBe7/Vx1MIWWExYK7Xu72w7+x1mTfSjtAhtm+HXd85mFrIegtBwak
eeOgP4EBsGzKWhqH/5eKbRpWWrOEKw/AZ/d1fYQkCaEU7a1exmLLzYUcxBRB5lBj
HM1vl/oLUW5ESKuiFDoj8dKqeEiyexeBosWodiWlLP65MDQY0CSSBeMCL/3zT1LR
H7wtbHJ0FqUZmUZh2VByvy3JdEtM2bP3MsYpPACr458LRI+EDxMagWnLfUOqntwC
M9ie/8yfdH2DsrxbhNiMEFx74apQ/yzRtgAsxYiiN4GZKeRt3VQ7Uz59lsM0GyZL
dAdvCgf8zf48HD7Avl7gnwGz9wJBLBZrEtC1v3ls7OiYGQ4WU774fVlhflrATuNN
xe0pdbkBKMejWDSe1pysbjv6Y9xEy6mgYx89Ju75h4Ls65qmGVePzYbhywox1FXs
RwogwFl3zpShuBo+9AFdMY/ZOSr5/Ys34uwrxZUQc035c43qtke3su8kNUmMrNUc
1eWgR2KmZhC4mb3UyhM4cDWoumVFDcC3Pf39s6YIFNCov4XyPiX/TcpfdkYXdWHL
bTRp0PzDN7+uplgVsFEQG6GjK1aDUdmEOsXBWoaywSqsVNZr0c5KiDXRRbFFMWpx
We2cbPVuCtpZIYl0JwIMV8+LFVREWV19fwlNSpIkIuEy5THYJzXqFTGU7PXFNJDD
QvfTYWq2w8OxFv46trZqN0TRXW8w8AC1Gm0OYlfyCK3aPq4E+jsCFvvbbIqiB+uU
tM9Y+mj9nig8PCudbua2qBfCyPMSRQo7xndKdu4Tvaryhc/T7vJdrwqCHObjA/oR
j/7DDYxFusqGY2mbsbSWyvv0pmtumdCnrbFsF1Q/snD2CUC/854cKYP4b+8XAqww
WQS1eOR3U+AqCDjBVkQ9V7aicUp76E7hnZM++G6Umhrdb00m/XNHJQ05jhCSgbTh
RT0JP2sWbOAkpDvOQoefoZ0iKcI6EvujJtsCVzwp+XPJWDQiNwsOJAB9UuG9ov4I
xUlUH+kvigjBB9m/YxNqx6CA/Sft0GXrcEmpG+VXlbiTHUH2lNS2Ppp7/NtUSFJH
eRVjFtYRrjCveLo8O37OwrwxQZljNAVtok9G56Trg+aJGHBymYBJ7lH11W09jHty
AnRRDJ58oRmISX5CloV/X+yGnEIPHnMlsDZitom9Z6W89JNFH7Xyy/lBxJoYKntv
hWkfxk3Ux3ePmJ5kQCpDGyMxpSmTAAjwevV9i7KEFh2MlchaQTQfX5TZE1mPFIf1
sWKUvNK2jBFnxuT6JBQ/AKhmDOGIjNdbpXTNK6AHfOLB4OM+9t77hAB9B+ZIDr2H
/HpSRKpTUcsniRaswyFbcsJnPT9uD4MqrMaRB+tKIq5R8vLnJL7lqhku5Y84YYhe
mbJBk2Y4U7a76wP/fn/CxIZKmaP8p6R/UQPnmSXUZFl/91LRiCtxfC/kksU6wNp5
9fZ6MQV+WiNEDq6JMw3B4LnRzZ4HhEvD2HPNYZEnBG6yLsoqtvUz93QnzYfsKRMQ
1H77eL7gpLnYdPAq8dn8528fNm2dsH/6ACfXbUcMBS3PaCIaaqdi4dx0Eow2pYMU
aEmgGcCq2eqZ5GtQNQgWm2SCkrS+32obJKUvTDW5F8ix1k+PO02sBgANbTRb40ly
/hR4vVVwCRADl3xAE+UHm1+Rl1cUINxCKotmp91PLVf4jftUU4UO3/8jm865hXBQ
Rc2s2rnpyUqsu99JrzLxiCCO496+HkOJRn16rOvwKjqlK2B17Kt2VbxKbIajB3Hj
YrMtIgaWO0+Z7/lYtSYosCsnNWsh7NAK24bpBYKSATb4F5hd/KffI0hER8Cwz4vR
R+1IpkGd+v95L79F5htAvg07jXFxcFAqwTtt64NZQKPdqk7R/og4IiyA83WLRwTh
YXfPGnqN3hTYHFfg7teVUiglqQBt1zYAFO6tFGihAdgpJjrBRNJSqZGFnvRf2+jF
rp6djtp9+9yF5rQmaYrjaWR7r2M7m8UU1f4Ga+HNj6Q/idsg9imNolbUIvcb6Dt1
QPMOjmDrzBEG8tQpJjNwU8Sk65WB8GngaPTlz8//Jg/PKZIlMKnxwcw32FvYIT7M
gV8pyJEfOz/4XXbhtmyrrFlXhyqw71AW5ts+7FaIEII0aMmH2oqH/Vbg+hMNSEfL
lqoD1kd4SzNykMkCiw9d0k6K1uV0DviJHgZlHeFqWtk04NEeHnzJCtIhZDcHRdj1
3NBa6FiRwzA3bt33hxnGTQ4CQDNC8W5bp28JGehuu/CwKxvoAOPbL0Qh8gFhqqs/
fV9hY1CdypKvFiAQnBjQgu/GbKO2VbYemhpovC727X68GXc+DrZ9Stpp8/ITNiws
aoJ9uhCSWqRYOEvvan5tENEPeDe07UX+Bc5Ov/Q/9WpNPrvDlwOLQyEFRr0hRqJb
9EuraI1hHb0FrUObb42E8TL+GNjJiyraCPBFbX8GdHfRtG344g82Ee84vXB96i+z
FQb3po2Ox6Q9hEmTNg10SaW23LYI4/za5wbrnteRQu/BhofdVtTBzZP6KSgc4Fmb
2mK7wWq2+3YOLrJzOh9sKmpbouwGsdkj3bIoe6GcWkedDdMe5z+qEeieKjKJBHrf
khk3jxpML+DMy/d2GfnFtGgsggq1QqRpVdaxgW96bzbVX++0ongs4ez6YO6PjL71
x78sA/BqFn//lM82VaBvWGVgjQ/a25cNEchXmhxDXwCbkoKY7XM4XH5rSap2ITcU
Intr54FFaXwWVdv+Sz3C6NQpFm0KLbU0JXo4HDIZg6S+hvnC0uEw0nIsP5un5vxU
GPSl4R/hHcxRrKfAMm/gQSBc//lvBaYa7G4gnEDZJFmlLMTpZZQUfLaQoH3oDEil
nL0pqri1XokdmMg/a+7bO8jpUs6CXqKAnkjO71Ici1Bkf4TuQn2GemUEoMr6ED7f
RbuL+2pDNXKwXwAsNE+20eKxyZHBgXOo7x4StrRLFkOYCqbWl7wuN2g6SVTLLMca
46rIx8eytjdF1AXMoz+ZnnX9xp1/P59y9koHsOI8QbEZz3DkyPTCfsML+VM0F1F1
qMHdNJJLytaYb2sDXhG6qIo+NC4H4Lf2eYat1ZwExKkkt42tjAvQ1BrVl3Wnntf6
OIRJ82xCAEq+tLp7Xhkn27wuQdCo/XD/62wEcu5MxuCcGseoPOTQWMLodFZYsvdR
hM/3KmcqR7/2eXugvW0E8zpAx4iOzAhCIvLi3J2SdzYjSPdWCXMun9xYdk/VffkT
W/9JhsgAUsWfPHeeJCPd45lHJevhpfjKLLox3Qbah30De+sgbfwCfTCtRtYSSe1b
03F2qO9L7LXOWPDfjay3ddFcyZtbs/kBnFZobqJQONM+urYY3LzkJkYIhQ3Q+kzx
pDIYwb+7hXWrBcx5QmcR8ESR53o2GdBKC1XbjEthaOxulwvOiS8SPWDzzTWhgPhu
6xiF3fSub1GiBj/X55iN/ctdrngBKliO8dcfzNq//OWEhF9uzXbAOudr4Q/eWm0y
yEAF1UPdq4z6ss2dj5K82znFTeEPYL7VpmL5Z8nI4DD3oGYcLvYmjt7Wh0dJAZaE
eNEW6EtugxbVuZPGQnQTx4MNz96juilWgTkEbCIzY4qhR1IArtmok2wLdDJpIRjy
RMT/hEfJ79nq4xVDrXUpazM3yZoFaDQOkzA5P1QjFLVFU87LLjuXRXzB0KIRMGVO
OO2ukeilPqJxl7AGI83mttYfd9p9M7EnoXxw0SqHB74IdUSNSw3gKqWjeCw16MVz
vFiLYHeZuMnXS0ZiYFlaSHEzUYWw549LMcnMWAiCNKTDm7mz7TA4BFt0gQvZJbQQ
NEp90AUG8PWFtV1WQwNf3fjx/8yeFdKsoAcb5qNNPGuEzEQTgkb4uVUI8sIif3eT
z/PPJNCxGgD8NTT/mkVcmlYhATh5EShZcsSM2nJixJ1bu+w8xllpjCJQLligbBzH
iugFUL83mc/i0wLfQhgWLsFOnvceLSGB+2w7kOnLDOJOKOKEZoo7eTid7x5hcl1A
6zlwVaeHYThUfyItUeQ1T6887CRyH8Y5vpa/MofjEnCI2u/2YrBKd2ZMPk/xnsBK
/khUozpt4NYMwzlaQcOQ4LEPse/1+2hl55MIvwwE2CLCl6WEoEEfALJhOsiVBRb3
QlIGUWou2mtOx2OqTj2yGHMvqMMFWyBnzn1aOLxgDiv9WSqrySGq4fUR9PbVrDjW
9cwUhZK78S+gaWC3xRMmRCL/lG0LAhTHoLhJklAtCWZqAi04KoS4p7woIuR0ynUi
JjxoMCbVjjkvg//UxAu2IPZMxgarB8RxRDuxgDAdFr1rfeE0renf8z/CxMKAQfGM
rW05ZVxVN3pifNMnknk3YBcXRHOVP0u4A1/OYYf774B+/Vas+wch7cfm4252p4Z3
0Ca327yjU6xntbQM1URnjAzWrAbUl1hkDpmKpMWxTpVNFWItYu8bSRHxOlx0X85T
FBuUk0L9BcLWYt4pY/VEanh639CxDM3vblErh+jrpELwI3+hJ5LaPxoRzEB1i1BW
MGeUlSPqXcHe7WH5GA+2TC6GvcBivjOzQPnh31TGwImQ748+EtozSjkRG+etDpmC
luJpwlOVxjpPFyqgwtPPzgLjxHnUDVX2ARNnFXtBXrD1SbdZ74Ndq2dQYz5PctEz
NFmFS+34AcjFjhEMUWsupVVKMUt7WRGcjlx3hPoI1lwYA0IzLmEfpRG1iUBbdjui
LQFMRKegO2MXsASa8gqOJ6EeEF5gDcDhsgXpMOWQCHdz6ls9wj7FLzkUfLQQLofx
n/McOx7LuEmEXNtGopHvpLKqgF2MZ48132egS0ztEaywVwuLVI9kl/snhXAiaeHV
gmpFW+N7LGoHSdhec6yq51Mn04m26S3LwdOMfVbcHu3gkS1ST/7uZ4kg/SQiNQ+R
bnUbgAU+7aXfgLtlQT9xOPjjzaHbPgz1M4FunqA2bUy4xxZ4vBGBCXTHF9xFdVTx
wIuBGnqUM4F6ZTPp8oEJ4rGakdsROuZap6hwXycLSfXVn7gDe2cHRS4Khcojynyc
feC5tbL7tsjKNyoTJuKbNN108At7XVp5SxcNCMr6Ej8j0FoRdNj31ZU5O4k+Ixng
rWrS5GQBpoZsgNbliXS2r31/YKVeALP+6gQiVpSW/ZOYQpM5hSzZaojIZFycm3+2
uQNwNYrQlaZqrmT0Oqw9Q8kJOFpQH6Ddps/5trNr+BQBcJlYNA0k8Ca3RCOF8BuA
hb9ND1BUkeQdtzG5EjmwLze3vqOlLEilJ+xqf4Npgvu1Oc+jd3feR/QPYkqqhkpQ
KyyD/sr56vbJUUu2QqR294n5rvyIhEgwS2w1NikAYW07W/yY7uf1wMERj5gEX8gk
55tq94MvISa6rkEbxsqW0U6r0PFY+3A/uoX+fvGJKG6wOmdilUq1OkWYO5R2c/fF
C+uOhHDXPfs50s75VUi0DJsjwWrvxFN7cSkU7pBQOgHPE/jGA+JlFFOEXsZBBgmB
/krGwA54Ry9SqNIq/SPUxpV+2eQ9YRQwIh1e/u2cZYVvz7DUfEaYM2jv3GDV1SX0
dEetQ08d2ht3gS0+63CQ/pofKVcRrGf0bZ8qi+LGKQc9SED1ZVm16affVrmveasr
ceq7UzBEQPL1evJsjlHzr/gVl1Rqad7MMMmFOBpNj7PqLVKZ3O6yq2ZXkKsDxahl
0YvvwG8ns5Y4IHK17k/T+w90+/8S/sJh2cnvaRZ3WMUtIxHgw+I0sSUXGh/9/zky
eFM6hBWMLlUCtAMbcFKDEgHqfkcW/AVvYMNyRnrJBfKq6TZx0ZtiIhvMgAd3tQ/n
+jQUW7ZQ4qsp1yKf2rgARVXerOa4fhFMbzfWprU82UDWrinF+W07/OZN87gOK/aM
xwVu6qyNTKxYzvH2NQjHYAsQhnrIwhbgyWSNISqX2rqRnZ05bX2cmq4/qz/r9TXk
kXOsJ+1Yt34a1TeeNno6Ni/+o4CTwGI51SAfzAoREonsnN1HvhPOfpzOAmn9A5qA
0c515tWRONSfR8sQmc9LvMQkrDky5ftxARRaCFF9juqcUf9w3mva6tbvF27aIhqT
JtGT8n9O5k8yLVwIqAl8V84qbc8AEiLj3AI7JqMpoKwCOr0o7Dhb9jiB6LgMejpD
qFdflOSgb0BSwWrMr8RuqLA8836ezDDoE7o0FkbGZaLlK9RRAeYMFUiJeESkGG5N
s1W2B1lP6E7O1J3U6ZuY2sOwbfahXEOdE6DNA81YNwiCWTs2cO2uxh0hVoQIqcHw
P5Q/m7YpGWnbZwAzfjVbQ2M5rAW2USoELckHmWD9qVLGNMsYcuLCuQeSEMUBB/eY
tuXqGUlX80eKfhvoJcQjHMG6AvHPjZxwZAqO3SH9B0oUZHNlGgGwgylFPVmhl/F7
MhWSEQnJ+yzDhQMcqDCRvaPKeqUcj61LVT5+jcHUGiL9RsDjQKbnLPf2/pSe8M7P
Bbk/2B7GEMEHVZa6BEuHjAtVE58rTgD827cPoOs8SiSmwo9nKCoULLsHD+IZHOcz
+BAGetf0B7VPrFSLp3/o/rfC7QZa4wtM0A0DsIAXNyLpIIE8HIJt0mUf9berff0+
PWvBJOFjBVeM8y4lvejsEl3r4RfKZEocNkyBs2NNwmTX5946ZqPp6rfa0exNtOqY
ikKyQS1JvkihrpQUHXEy5hl8AH0zN2HizBfWe1t5WqSz4ZixanHJeFanZCvIlZJQ
yurSpTUfbPKCYwTx+FT2NMWoat0gk1tZtdAi6pR8qWJPdP3750k4SfPL5wFIp7NZ
tBPpkAzgnrJslnB5sVWlxgZ33pW1cCeqX300GJkpA6Hty/n/7sKYHf87f3uQgEc1
53Ypzw8Oidd5uGzeeWkFr/W/cs/jre1dasYHHUM9drUCfxSCeNmUf9BzzuTJUCJ+
WR948D9QZy/xoxQ4VMDqAX9dcbm0c6hU4eBPC4VdPI8Iln69TvJIveuF5qjPXJ+3
LN/m82fJcCXiva7Vzw+tx1OOuRm4DPBo5KWDjaBkr7jCfG+4dIUbLkcs2fXShgZe
Iq88YBqMv2/HV/U/V12f+cXqbt0M9qgg1UW9ebP5axfMaXRNpcFbYyWH8AtduJKe
HRIQRqRtLpsj2S/YDR8ANCed/DdsfS27Yp24amjXvJw9ef4g/qMgX3te37+DyHGB
oFMzRoYng88Gjcmun3TnKqV4fZqE311pB8e3JYBjL9zRlUtBVNqHWtGSRkeFCPKd
Cy4ef35NypJITuA2u4Dd8hLa0aUzEgZsP4MDEcp+O7HuCfxP6gdLP0LbeHSt5h5x
ijBYdLJOsTwe/6mSo2fP5WT7xzx+SD7hQ/OCG4UH4cyxUnOmi/E0SCdF512cd3WS
AT5uYti0pARFP1fClUOP3gtTtDtDI+wvNK6id86oHV1RY2QDaVJihxBrfyk25RIC
5+U21C7thh7i/ZbaJroXW8XKfuOt0Wm33jrc5+uuJpFPCuxBc1bPzO4n+WXXgK7O
EfCzZ+5w3LKa/DMcLtTPu/4zRgFYd0fnWdfmHU4Acio3HKT0Lx6HaFTQx+t6O/FS
/W96QktT9B0qiZS4JxUfJZeFgB3QaMUBy1LztWiIFWcBEkJknPAP0IxQpqIYSRvB
wqXY2pM5RUK3I06DcD8/VnOlAHTcv60K+8X2jcJw9OmSn07ciobJo1ekYRselky3
MXViWeB2R2csHe7t3Vc2NChDxljcZhChFi6AxBLifbYdETHxW+aBxDjg0XkOmsMX
WeOJezrKmz25hHjpnuLXgCw1MUfOosd29d0sxZIGRPaBmsg6VU0NG4a21H43v6+K
Fe6zdV5Ya/1FjuMIfdfuCZB0E5We5uwSqL6HAKkXK8oNN2DNMWPJZAEuuCGBbBew
A7uwPUNc12k78a9ePl8DvRqHk9zdot9BGX8pE8J9a7hPZqICt7qXXRP2VU66ti5u
y+RHrOO/dw56L/wZmyOZ8DAfjaoirERk0U3kAk70P8RqMy2yW18ojTPSy+DchIvU
dQLT1P7QC1Dv9LC6DwV//QipV47YGNJ9+NQyVe3naCwq/8bx4ljZt1C6fqYtd+MF
IntK/DzO2qr+HPDsUTX/8MPlVfST6667X7Snh0UY4wEOmKSZVh79OHyfCh6Q2Z1J
j7Fy7lwEp9E0vGQFgT62IlcUHw85EggRCeqH/fDEXXO5fnKREdp4kQ1X6dAFbhsp
rvU+ygczVQJ//iKq/KNdgTX+pw5dLiQ04HJU7b/QcTZ7EhQVWeZEX1h8lhGKe8Bs
qTTfkursSRpEjrQWVSxMBrsUzaVKsnn/fNhksAoJMcYL5YiVylnWiWGrrHLqDRf1
qGkPLNmm+eYzELdolyax2jFYEsBa6p+/DJDMcVn87tE0R7ZiwxnBUIThPm7TfyTN
tLevtElavOZcfXQAsOj46AkH/hmS76/fGF+QttRjHKqH9hsXHBoo0ym3BSXBUX01
jKhnkzjK4jcueQuETdbGWMLv4ABKPsyDTFDlrJunUk82MYZq1V5XuvJdWVOMkrPI
G5+xG9CQ2+EIWiAmtqCl4FhX6hq3zMPUfDbAgTqku+UYMxeqQ4PZQz9VDxGImjbK
venQia1qAQPocHJVYWW5fZv2cmptUg/uufaXKZ7obNY3jUycv62OaiogKSvYiGcc
5MftE8HtuQ6wCdfg6D5fUGqzpZg3U+PgXG5ES+bJOAR72rGcFtBgqDEpaEBOffLD
iwizGHuo4Uz7zbbQOh51VWYl1k3rb6cfJVRJ08svUUc5XBAl/eJ3dVxsjPy9LS62
QI2qk6rBn04hQAqUgdIVn7JHCY+uuNPUJSCfUCiUnz0i76CmT49Boky+bO2Nfmu0
pu3dFGPuYY8CeZ7FYkllZg11PsfKaWD/pRTXRWzIl9C8erynAtPHWBOc0cF4W+sk
j4xyt8cDQjZ6/dYiXMmJBIOa8Xn5oZnhBHgwjUi6nBbgBx9ZO3ZjaFQJAJMvHkrJ
9aPWiA26Qe4PormMmuAnx39eWLVx6kXjLZRiKt16qF9i7D1CCutqsA+O4GkLTLZR
Szi2SDFEt0fT7XLq2XJCRWBezlwCbwOZQ4/plkDZxb/0ACLRKBzJwwxD1IZZd6wl
whr8dPA84e8K5c7q8S6rj/l6uyhZaLQeYlECBGC08C5pcseV9HDu0+ookzthcUss
E2APoJG+/4qeEkE4RPsbSvixnT7VSA63q7tSUgXi2hu+1bRKZO9wmwk6OUoxqQo8
U3u9L4UP9xCOq2bX5emD73pQFwb6xabuqc049SJvtV4JhrAsmrdh/G6lDz7GUSLQ
NW9usin9HS5DKu/SGsYc4oz1d0o27q+zsRjMZBt7odnCUVngvOfruViwoPE6l/5O
aKhnwuyh/dQO14yX/RINM/WgBHqMDThiJ32cOly6bRBqvGwU/7mrbKKK87MjtTja
WMJ53PseY6iYlsa9IjICDYEm6niAlrVv1/kjQOSdHqoOjIySoWVducwRHkTowNmv
UxQOJQsCb007Fg6+5iAXSltglE0c/GklX5jvMh9e+owaBAJQZLvyZeP2VfGzL/Ej
e+NDcLlVjZA7VHyPcK4qB/jLmw2B4lspYesdOmzOEJ7gFZN5/mwF1A8cKtF3wFIK
F8FDYRYOZHg6q2+0SvyttUmYYkaA6R1KQt3mR+fZYXjiZHbL4Ir327G4zbu52qL2
dqahODgVVQfqSjqWSzbGPEhO+L3yPGuEk87VXHPJBkiz90lobe9XFzho09MhUeBc
EpRg6OjoAmhWSgzMcwPm4kVfgUS+4CPeU1jVA8LsCBDOTvovcR4PTsSbvpJZjXD9
K7X57t+QqVHs8/8/64/NUreLVnXKUGauP2kSi8SPQEB1Mui1zEr+jfMKjM5DLfFO
5ZAz4efg5PFKSlOovLZKOT53BVNx5ljTzjQa1O0TjA8J3PN0SPePHVjlQSEv6m1H
t9G3L403UFkUsITMY0v89FertuoMuzfrYQEWm1AaleJr3H0DPpkpfUWTx7geO9QJ
j8b8qJ+sguLjxCV9PUfyvEolH2b45Vf1OrGJ3Asj9aTE6EftkVK+YhJ6sk7sN028
TOt1/adistdk8Omb6nf5LwsWZd4WBCzPiRVzaK/0ZtfoGTpK3DkI9gLHcreBQnYH
bcRAAoisOJEnDPgfRZylUUeJqKhYvbfZkROqch43cUykX5nBu8kjy27dZ20UWYFz
Cax2oMrI4J10ZqD7nlXcxBnhvrvsrtQha6+LIRJKBVJGV9BjKgnI6cx8tHx5Nfsc
I3zBgQHx90qjYq9O95PpVmSooz9pke+ynxFpEa+5Ci76AcErS4r6P2J+fur7quXz
bs8tRpdWlBdg8/3Q60j+Hz3olztptTKF6T6hhuP3oh4OyXHA6L+sJEHRmOXA9EO0
YRdwmqDzsOb5TQUFzKoADa2kDu0FyXYJrtuTuAZ3D+gw5NlsSqGK7kR/NLLz4op5
cjOyeTw4Kh+0TNjFR2fIuocQeoi+XkBWzplpplM+VOnmSHjtMzC1GJdgMD85l1op
mdI46DLVOg/aj0OLLQv61FxTtuQc1oT5+g/jWMkv1EsdlM0N3AJ1qafyiXpC0xPv
hkl643CpAi+xr16FB68ftxKescJBOScAYZTyaPAlMyWLuE7NZRgMhwPB8mzWd88h
Xwzw5Y0mh1VK1NTmyAvW8ErOXzkT/AiQoZngvnCsHQa0k1xtEvEQtd9oVopukZB7
HRjyxuaijvLRlVjaQVOr+U0vhfFC8ih9Lq3+NDTzpaR2HTiwMvIfnj/fdPV5OqEz
uOli+n6vS0ATP/XqIZuX2zYvBL5oXsEBViAnXc4ImXPfrbGjPY7KKV1cGCJUiQBx
605dDj9n2t/vetnYSih+y8yL4FOhq6gh4YXb0eihFhS0hWTFFGen1UL0wT9kS+YE
j1BC/4x0iFOWxbKGZWczYhhqnpHVW2E06iWWbMvptapVcm3Qg0nFh43iOzhDkfHa
9WHWeFjzaUfV2vH/2iDX2ysZiJI3jwg2xOQYZ9gsfDEZlJF/5lHktT+V0IOkLANn
gUGXW6+/PxTlUlLgzI3SOiNDn9jjQnpSyaZoMhoouQ630VWwtNkQWspJrNZ/KqX3
Cin2FUcYZnGuuN+CXbqVYSR/S/JxM/YuKMHRAOiUtCvNLJXBpG74uvqUlDU+2CWK
pUrKJy2nyPCc60GPJJ6B+zf8hFH/Rs8QVsuXHSw26lDmALqSwgAlV2e2JqQ+bssK
FhWNnJT/YUN7TF/OOI4q9zu2hbTjEfwURDpL1BYxrVl2lEkk44WZ9iW+IkhHL/np
1OhJJr3ODyBLkugdAyY7W49DX4sfqb4yB4zblvE/Fp1bHKW1uRsO98jaL58ctugj
Eq0WHGhXqcKGl4CFwQR9ymdqbxYm5Qwb9O0W1xNJiducFGTN0dbeNIBg/ndctqW3
lBf0BA6/uOpHMHqABICSyDQWAHWHphTO+S+ElBXgjw9Ubppp8tWMo68oLNYFBKob
kP3R/loZmFSGWIC6uNjiuQTuw6LaycWCMlN2Mrq4iV4LDZMe2NckkBkVrV5Dbk+z
qQr8nZc9vELo8hYv0hih3v/Umr/DFAW4w70vHtO07lLvt0AcBth/TJsI2+3eG5Rj
P4AjralJGGNRjYaFhL+RgHD3wWlJJ2VLamWw2PPZREGaEpBROUcS6nhMkihHzzoO
d46p9tIGt3zwovre/SiAM4//cLQnhfVVGbcKEqCj4FYWru6c3vguFw+0aoEZ5m2G
US+N5UZt8SNCsAa46nJj+Oz6qEVZGVZHQp6baIhwbEjj7f6XCZfXzCBSnC64K3+L
mq+YmFrrJJT1lmtm4GquTb0t+FDXw2OIXQ0sDoR0Plp6GSZPVxz0uEHLcFdcxzlu
cDN657u8I11f9Qtdne3eCZPOpPwi0oOgU6vARUv6wiKYNzSX0BpvLnEt8rarelKA
2LzA5NiVdJNvgCALgv93ncYL4ImcoKexwZTs9Y9iCpzmMjiC2CETvAQcF3ENiqLf
THXBQeZbiZeTGrTbRlVnQVdNKiWEFyn4qJ0kV46r7EEjV4SyAyAUZ4IL/WMZx+bx
l1AleGDvZwKipE1FP73bP2yg8agXcBjWfj+XapsxFn1bp1EO4SUrGO8ldH94vQRZ
Rp67PosuuvFi81FV7rPqaLtATCunUdU2ID5WB1YXpIsm033w4d2/fKilCZSK9+kj
Rxm2T2oAnAav/RtN/XiYVLgK+ePlGwnqLPDEUs+reBzNYB5RVUi1W3SBpgP4BiEs
YG1q4pd4mRMW176DMbi1+I2aG4AyM5qyuoUuvs4a3XX682WNrvjdrXuqbSsFdFh5
IMtbxw7LswHMEUcMrLlA383AYt2Vnr6DN77/Fk73pW7xcSZAIhvHv6UX//5A5ra8
LVvbKIKi89raAMwnolweF069ZJQT+5SvuiHpevKTZyK3EdYN9b0tvaYplVtlbqR0
m3woJo2rgimffr9j15JwXznNU3VjxmE0fB3PBBvpfR1ZUidTRuRUNYQaIHruP2do
EEo8p2WHPaquEs/DcS0kyZSr0EC2PSdNrA6l7dGM/6ZvOVUF+CehbR+Kr4ToVXK0
N4nrDpXaF11upWkbPbuOimotzTI4ojy+qFqG0Zom7stlQT1FseGgj8732ZTeAqms
w3u68/2gPTL5Sz2erlMRNVkOdq2+xrFjgl5yUNAqlL6Yvf+byma+bsSXnSf1CjJ8
Kz9GGeHQxj3a2DuNQI6gJ+wiLwtyPDyLzmioyGaU+KaVxY79snzmD2HDGvjbEP3P
sMmVnzXmgc3i2F/q0DtmuYgZhOpI6jQOjNnzG+7mUAJB25Q/e63Xx90RhGZRcTW/
7EsTk36gaq0jpGhr9AJ+lQGm9dwLYcLDloPjGW1sToaAzh5TH71HI1tP3peOwIiy
1E8PJzmWQlhXqazluahzH0HJmH09t4B/f00QjD04wNmTqMyjZlHAg6NpE2i/XgHh
IAGHrQWydzdLB6FhEzKK3LK/79rPkQxIanIVeqwH8sMfX6vNwzzar0broYoKSJp7
D9O5nlx0uUcxSm2ies7iM1GZtSLv8dGRQc81LPEl62htjZsGDJzldy6bFLRdkD8d
VSiCOSul5EWKpHB1xpFBFe4WAvZyyESL2zCMMQH5BRlas5UrV0qgSrcqAEi9r2u8
qYq7CFB6voZHHZpO0+2UyIji9NBoQNsWpykm7NL10gplowubH4hyyhzOhkI3wc6q
G9XLn5saIDfyGOCrJii54f1Gm7c5SZ96C3ldGcuoosTsNQBwdiBfksmv4IuHsYor
XEwFkhorG5Gz6mMSK3noU1xE+aDJkDISgbE3oZBNWUrsiGREFLaV3faT14M7ZGcr
Rjq1XJmOxObLf20CQwpLqVysRIPuPN26lEvz2v2ZKomI/6ZUY3uxOqzQ9m+Z96ED
A0GS0cdviaRCFdVOVPiJDjNoZYeHY79juTy+6mnZfQ76qgrXFRV30Zf717Rvh60f
0lgkAkaJZ9gI34bFLaDsMuimzj6hf3XIVgjl4cxD04D446qmIU6HyP3xA4uah4/W
L0IGF4RqCL9C5AzzKuaZ533wSP+OeYqMIOPeC5C5e6j6WKYBsVwvRYjvjfQhJ+yz
alBO6fGspuPxGku7DNvrWJO8kFfC6IQzZspY3voereh4dY33zTeidCRxeLsxsAje
4vPKCvAEfK2vFP+piF5Y8ZVYeHpxQEYNdvd3ZJA3gRz5PeUmuP9UEW3Wrcjkdi2p
UAOlRGMCsVKIOGwTJ8v+FVLFJ+YqRU/RXh27dGd1EdZV42u/ehsWymyhhq7fxyHK
7oS5qybqv0gMTBgThBw8MjYmSHXkGCV9t7igEyTpdLNYHnfeB87FSBrxi2mRVyb+
W9FgDo7wXjPv/cVpiwcz+2oY7eTVTY5IQnEnt9FgbxlMjrSJkNkYd5ZVQq8Rx+1u
z0bSZ9GrmkVC6rZ1k937gWh3jucxJYt7xlnX5kYZbmF/RnxrL7ZV7EHC82Puh5+6
DC4/Ke6JRMddsYhal0XdmP3geBky/z/ZjYLUO5/3/LprFBwviPAr9rtBC8UOeBzw
oe4z3WpygESEfvWEDnoYnq4gTyWrlOqzGk3Rvi+0WnvaNoFY+ss6aBT7uBrJmWnc
824hit6XaxJ3+9GiDBIHUE3kddsmUqLO714JH72r+l5LdBnHWc4Oa9/FqDIo61II
9rEPnU5iWmTHVkMYwH88w7mZ6YQ3FvpvJlRHn7TUcElqtIoMoGRlZS/4S11yP/tH
C3tNa9ogQAsHSXflxstnNfb4Gx4vnxojfYb6swaQPr3JuQG8rZX7wmnsspsvQKb/
wTZbNG8U6TQBnf1qHM7YR0c01V0JYGRgfkHGJE8eaC10P2Bq1m7ekUrBDyjWswZy
QZMpiqKJttM92rMcbxMudpQnhzQlsVdSYH+4fIG9IuFcC9TI679LIjpOtN4GMNJU
w1LS1yo96xtzxfCyiFO2WmgBF0R6tcEjEAmR7R/oQWRxvEqYx1YJCcZJ08mT6YIF
YuJlwvsqo395qhsWaQV2kdJlEbcQmmo8hktmj1w3xBnTiLm+0smrDkVjO533Q7AG
qrDQDImB2GRsMACbXVGBUzLXNNYnss3EVQ1wv12cHnRJPfr28P8rtcKFUk8+me7O
CS6sh1cixtyPRz2SNw++XECB9lxr77fGwuRY0K7PM++5EMImlGJjTQCOcX1oQpOO
WfGcVC7qzC+Z0JSC7fQ9H8AvUgqeKSNhwpptqh4OFxF3loMvzeijTFL1FvH7ieao
ArVYarL+womoT3G9kSSbh5uSmN8gp9CmZ2ZpJMYx12kLhCiNkO7MEaca2orjoxbx
cpnVicj20VzFPQj4/7BdgMGK6A4iZRxevvHcoSNs++XbBDylUWiljO+sLUeNOj6x
7/Qa6x1mEuMDkl5MaF8+QAiWszCYUpAGljX+ScT7285DzcaWzKLCWo/jCMIdI3ZJ
fFO33Ow+6nBb8RAYTHEuO2IYLnnkUGAbNLiUKAvKcIzWv2ihH28njfMgElZKeF0D
AhbyOf7MFYkMnJm83wARnUHlGjvrlJFm+/QUNJL+mlrTeYq4bijuT2g4gzWpYFqA
Hwm3x0cllb3hteD9ydz9BQqGM76iyKJaqzj9zOLQodejTTzsPfcOnacmAn7KUi88
VOwVow3JmD/tENbNOJGYhpA80caVa1D1kqpeB2cqeyPKRB4JyC3SdEYXSDsgZcfE
Exn5w85ur4i/E2bMwaEsiLTgFlKHJEwvfHQsxqqiNHBBTIsbwq3/Lqh6k6wEg/Gf
Iyp+81pfznLf6xYBu3QIc4XNFXw4NipgLg849Mft822l0abtRDy83s6Bm7LooyLL
u4CDcLosplnlgp5u5aXS3HVOODY/hnezVJsEkEkX4YME5p35ndy3f5RfiKHF6kpq
Na7vz7ODjmEf7sY9TgiXEvC23XAr5HwD3Ymunk7V76RQXAHx3yPR4M6fizC/tmZw
DhNwM8DGdTihMYMrohs11oqZEEM5hjqq8ht6yXSXJ+V1XK4bLXfukBvvmebCsDQo
h8KmzY4QFK49pmw2J4Wp65/lqCWc2AepKky+hZU4hwI+VsqFZan8Abk7f1puh/pl
naWoCn/uTlSiIShFe5Qdn95+fMPWqtyP0oUu9KJcDPs5WjttNA2bQsLBu1n54R9W
uXmPz8NnhNRRi+nOWzg3lbbT5NEGsMnQrqq5TZzuuCTrxvUAedG3Z7IRW8rC72fo
vUk3ecsV0SiBjboPeGpOpvnq755b/k7SpW+Aza5JFT6rafa2AxtzAGwQhZzsfHg9
TnkZcxnYj++sBvaTZS2KGrx2tz9CanWLFvmDDX+Q7xAFCFRUd6ZxdpfY3WKphOq/
bLT+PZ+iflRso8XrcCCj/NlYEPCb/E1L48fnJJv82JONvqFW7eersjr5K3Hc5AL5
rnDrXr9vtH+zN3iBXCheU7eS216tOiyIN6UtgLEWgt1q8S26yUJxBkveWCHSvexf
WPrZwGRQPP10KUIU8DCi6tUGNnZnEbl3ugquh6d3mgmCLDCFzVxKFiZYTNu6/ntB
GXJxmwnMN3WgUUWK2tU+zRrgjZzzVm/EXClSHRVmzKb4B6E/zEKyUBR1hR4XK6I3
fhGgg03TNeSbVVXHNZgZKGSLhVoD9nB+XFjbhUvpeNH/qHOAlGvpfxy2yEl338UT
XKAMJtFC268lZYr1r5f70uJN86kL56pmtnYHjKVgVisTWDWNuBMp3XLzl4FsukEb
M1ox/e6lErXpqMGeCUKOaFTC4DQEoN9Up8skVa9NtrdfFnY/qIaWkyK4f7O/EV0m
aPQ/xURTIEPBjmnVkRQUr0kI8FycOVDE/mltA4P1lpH7qmM47/Qj7PS84wJZzzqB
VLPDm01a38AXXMlVp39ITStpPVsQTGWlUcs2uWt5V6Sie5alZgRYZEnxNT+k5jR9
4jpr5OheHeh3+JqcOq2YIeFYLjkbpbBQ32dBbZTrp6IaCrA7n90x6nwAMEsErSxh
dKPI8ysLwPwB3QFk+XnodBtQ9DABLTStWdJgR8o7zEvVweT90l0gM7+n64q0LFLA
MEp1GwjofhAA0Oc6szcs6fbN4NnSZ7kqcLfW5+RVLJVvZQ/055B/7GkmG2lDMB7A
CAxh0nvWntQRAQyd49UfxOqOR+t0DP8cbiqSBhO4sGJQjoWtHs73h4C1mtOPQhyS
r24oGKlJKKu75WZFl22z1QB+wGLQLFAWIrCO7jt+dWz+Fx57qhIxTrYw5uvLCDY1
lqdHVUXDymG+988h2u3PfLDWMM/sbXjAzK+Xb3FfEkuJBvWQ963wJfazVU7jLkSN
NFRhzWdM2MagO8K+OhHNVjhv5rrefV4YXsH0Q0ydChD4V68OV/neH6N3QjIKyP+7
JiDMD/AluyWNgUmvORX6ZdLgoJ6psq7yYJsstQye4fqIW/XPDrA3lMpAfWJiZS8/
N+L2kH4gC8BUh44o8XTJQcr/7Mpue2OoUeD3OryOEsDPzG8zsziCczj/w4HiGKaz
L96I6bFyZJQX7XMBpj9IQVrZH+XoZ1lxzLa1q0uuvK+wK4cwYJP+Ht1dt03CkTK5
2Jdk3Wf/Vcc1bO5LD39uM+b+imc75QUuuADXrH21aYyQHMrrpWK44AlmhMUlQZH7
I0J+TNIgyQgLw2NeQfzvltmizIAHThcaKOcQI/1HQKYqmOc8nFkJEWp29wsYqncI
tfVxypp9137If7tdQTyinl/QWNJgxdN17j0cXIiTg2TeIgrKaxRB/rzkenn5rLB5
hSl+xNnOd8uFtGTzRChnp8aPL7zqkV40M35iZ8ncxNb0UXRQHjPT5rDOUXwAtMX/
PUobLb6EjRRD9wB156RaSSX8Wv4mUBmN3475G/NTPIpQARzsyHgxA5+kANlymKDr
6K6PlqWVUiJMjaxTJTMcg4+q0c+58JcWgZxze6E/Kmm0210dJ2mprggnkGdPuv5Z
H43MJD77ZeESysDXWbbvqFzY9IJk6JdieCpFoAbsrNJPzRwwdyX/SHcUdl9TChYQ
yq1bPj/RHt0i8VArz66iJfnLTyHGiINa00K8YzWY8qyiDzKTEaB1XBHm8E6pN1Qo
UgXJpL7SrXDQ7p1+R+mudbuNrjHQIdYe6TcI2K1ohgqnO5UdjlvKH8Mp06TUCy0n
gGiVi9FTLiiLZV7cRvpedOVgM1vpbuqyBtlOwPEL+GBHqULcqXpMaUA3uvYgD02C
/bjmu0wIZyCiakJ0BoCocXiMFyhyV8Kahb79QUKOCM5RrBAgkKt9nGhVtu1KiZQw
sUZ9C3ZfTvOCD6Xpk36Obn3IJF1KTvd07gGsOTSJNeMmCq+cVyfxXnsdmghjhYLS
7eRRul/VC99MKVDRcVkn6fzoaoRf239RgX2jpGQT45g5wPJpOU9KQUcMfZrkBKY2
a5R5dT9WY/vq0KE724nAeqU0I6jGQhnZaGiwcBM+tky+e2UxCJOg7o4X2/Sn1G1x
jsrc2123Yqr6O0XWgbz7o/9GbbaKZjtwC1+lAzeTicrCzPXX/X28RADaXDr1f1DC
zR6+w00mG8/TTIRSwqXW6SQsj2msbYDJ7hB3sj0v8loSG1sj7HGrP0LJ5xg32iZ+
xc9riIkQ49g3LC99xj1/Y6S84ZUvGh3TuAEZyrAIpfOe3CCWfTtesjjVWrbWqSIt
1OekGPLoPv29eMeV71MwT1koyUJ3390dkcuzOvZzGB1Y33UewviVttI33X1j1UfR
Ijio8YPBinobd6Fi3tmQkCSoAQ0K1SizUF4tsBCKdum9yiczIRJ63vY25T7PXpo1
xnpgI3ch9Vq6v2hB2P3Lc0IkAWKDDQF8y8UcQrPt45vCazUxoD0337fvF1DhpQxe
Y6HK948s4nkvh8peLtbV3jvIQ+D+E0FajNBUAfugCHm6bBBC3ECc9MznalHb7cn0
Ku2NTw8mqBkI2599Ta55sPJscXDyAtXoRmxuE3Dm2mTLOnUuMxMwE8IVWkk8g2iD
VzV4dhHVPHj7Mzwg6Sm0OfQ/ip44O7DpWgJwZGTCtQx3bHRHSJuSB7NfKYC/8Xao
HoAYN3YYFa1SMcftmJ0SOns31endy4BsKMOmQ0tKL+Gv6WDSk3P1dTJiExrlyRei
D4LJQPZK+RRVI9CZ3tz7/0sMVOlv3UjwDCeCI3SYoK8E8VGPHU6N++QPatdNmk3n
noyLhy8M57tTKTdZFCz8fySV+as7vBT6aRyD3TxsXpCMLOTL2j7PX7931GPqpry6
IkDSCq9vfLhmaVn296kFoLWNSKLQcuxjLbVYL2YeoM1q80CZqDRScSqPNwB5mISi
pI+QHISts6nbwY9A7Vt/FNCZExUVmmr9rqfQr3E3NakDbn3KSAX7BOZ4tXhYFS1b
A/3lPc+L6lIcK5Q4SO3Lyep8+QPl+4uLGVU6XTkRjDTSZg/bb2l4T6oYaJEvG/Sx
Yh0HkfB1QH3M+YtvsPdlYstwpzOA3Kpz6sCKOOUQxzSAy8m7w8NZf6y4BZNqKoql
a/Ndq27bDThzPuZl1Lsx5qgi8inN+QBkKBFLXamIJgzd3vxXyvx+cqArTimsa2xo
y1KgOH6KE3Qrbqm18ds4KhX7m+yv+dGPlqAHOmuCspkNGYTIIGZ2jDEHkTb4nvuO
eA1qLHCNDPjbERtmbqAs80vA+yZJkOSppCdpwQ6Xt1jxxT+pIYJRSbOj6lSMx5lG
Xm9KkyO+PUJD5qwF4zxhuYj0X8sq4yq66KBtCC3NircC7VGwcn12wkdvl1ZKQjA3
D/eQDR12jW2ji/Q2zZwuJ+FF8mb4n9kvaNXbsSPLRfKNWXi5igxPMVdPltTa2+gc
KH5H7UvziRuBwrE4fvFsBGBC2ef4FXd63K5F7jQdAnG6JdKHVFx5jQIk9mKQ1X1W
6VJQi3sEvUFll+qwbt57AAyDvWJwL9P91wtfBLJDFtpW0PC4zHEo8FhQsn9lr/iG
6XwQrdMRCDknjmhnp7ZRZNWWOjA7e3I9nJiXgqpU1A/6dbWy2CEU7qEF4uP0wyoM
KvPmB4HlNYgExKOR57s21fLe/PZap3fvRjV/jmFnSo/yjJth0rSMSWplBVCjwhQt
8q9JE4P/kblzu6E+G8Jre48vxcAiM9qEPY/CIJZFEsbJw4xhxFARoc0Am9nIq0XF
6mbnuNt3jZkoers2Wj6vjcLIHAL21cXV2D+FAuRwnCmN5wjDNWGW+6YqPIkfeBPx
tihzu391ltfRBWA8a2ysYPnsj4QgTHVaIWWMMt+v3N/UVuMF8UVUMLnfO7piMw8j
KYuLeshUE7yJKy1Xcfu6eb/jOvy3EsWICtYk3mRmzJyukcfft1WIPLSuaPpS7who
ZwULWOpQPxqu7yQUOrFExepJkdy9FtXwkrH/wl1vvck0QkOq8vJhkfz4j8fejR1B
Ch7yVZ28eYBjjTFoPLAb5mwl+54Y3KDwS1VaiNTBG7JKFji6xsRvWGIAFkuvaoD/
1AgbMPVz3Xa0jXiuI+VJZAvFsDPgjCbP6Vyko/rq7rCAo1YyiO3e1/BCpKvgI/dI
FV8BLV5XtxB0EgCNE/toYK9M2ryiGSqZkbIVyNV2X8o+sYef9QZ5vd4cidhZpceI
2HJLWbWcZxjiTTlVFAgPJ1R0vtXIamFZ+jd6ZksRGLiFbwV6Ieng06db9Ga3aQ03
sv2yXJhYeLLXbaHX54pLbWVwJYLg7Xjw1V5JI3bnzZrHEI1KjsS+U8IHU/3t5m94
JV2ymN6xyZmfm87soB2zmTd3j1lFSMOCH59lezeivLXf7XUnwQp7HNDkgwDz8Uo3
2WESejZJl6yFYOlLLW1dhEU5OOU09jhzj3/1UNEDTbWT+8gU4heBEIDIDZcYkBFz
IpIPperViw+3uoqsMlU5lSY9ifaCLMNAUzfiJ86PP02gvAfvx5Z8/XDRl9ZOCACA
UnvPCas6KuZhZNLV3q/wmhp7MprCvtUmwEJ88jp6dHpTqBDMx5NG4nxS2kNe+kjD
exTXHiIailj6YgrzzWvOBCYIBrCjYY7pAB90vjuixhWWPUZyWXNcr+gYPCRNHRn6
fWPzHx/bFHBiBn5UCGhoKI+DYMlL/4yUdW2pGo2HY6Zsfnl86Q0aOW4/PLW6E478
Ft/oGM1Su8JgoeSSqau5UQrkI6cADwpTovV9VAzIUO4FR60EfWhM2Z/4ZeWPzIe+
U9HAgeWg2P4bruniqv3Nn894M7CNkgMMznucGqyL2PoNgE4Glbu257HrrmV/6vZd
LHTzvVlYKbmZRUE1d5H01kHZMsEwGH3GK9v30qpR63gFP5HIR/o/dLavJh4TUnum
8hcFCvpxRUkLUy//k8YUR/M6ABPtyee24zhEH9Nl57T8fLo5TbjYUWLSQ5gw0oUj
YmDXoeedX6Bs/VBSVQRfUvkIcQKRi8JLyOl4mmyChK0bxEFDTLvgl78v1dECEItR
w1Po19IIr6B88tC+Dh9GpqbN1pbe+iSF4EF0yHnaozjrp8V/YTAr8AJokDCvnnu2
z4Aruu3NWgmaj7oedajBh2Wzh9D1xooPO1GIs1h4wv/Mz0Shlgw5n49U8t56lFVg
avw5Yx+B0cVwrwYwdiIJLMKhRK5z+tywSSmZJ1DOoUK93Ndycwnsk09QSMOCimof
gzILHrjZTyJ6x1HOMenpx2T9XdyJrCVG5VrKLffzOa8NdUw9+xdqaBDR0f2UmAIf
YegiFswGP5bZjw4qg3tUmaOf6F5hddvguwRNZyAFpMVEpVhbV5nnlx8Eppag3fHt
nEtogczhwugtgJcNb8AH3HDlSiAIpbtVAr7othy8+TqLaFRfaxhcUjO7scOBP4pW
O5kS2Cnrr7Et6nVqYaUurhJMnuhimVoqFeWFa79AxCpwNrkCmqH2X4IeZkUGJd/l
yh+sN25f1sepi40JxjCY7gKF/+4lfZJEM2/9SRbN9+gI6DzDhaWQF/+XIZIYzn6/
erD487RJ+EqMkmQI9XEo9v4rcn6RKnjUbUu+yUzELGeZ2xxoCriBqPWPRAwECSUq
gCekVTZj3XT5VVgIqZjERIYK3zw7inFuwr6qwhZwYnB9mHlr3M+c52+oARrr8ZrQ
DBrz2Mv+D0o3R8eGY4tOnqLLGeGjt0WOoQbJaHGQZne1OQT54TP+fcm798Q852HU
pRAmYWQrkpeMjeDyK4QqRNgjeGrERr8RA5hTo5w5GGWlBKxpGv51o2okX0VWHs04
lFRBPLpCxOGgvOcFeMnJwO7jvyu6iJCXZ80Miehev+LLZA6jZYnXQGbfculMKidi
VniYrmu3+Wqp6Bgfz5lmSKdD9qadO/xCrfgZ72ZgqXF9knFdJ9s/LPoMw6A74CTY
gErJ+az11zh9WFeI0anOx7+BHN0czHvoVeliuBJV2B/SG7rC0HzEWT5qKX9RxMW4
dQnoXNGs2MLRLk9qy9uXByWd+8IF4GzXHX/lrTmpkAh/YUSEMna6+t7fmWEdhDlF
GW5qk7pdlnJJyHVvSm9j3qvWdJn+EuN5d7r5gVpJ8jjaFWSBM7PsrOCrfRQ1ah+S
ADNXOQ+g6zd44ysMLVvA5StCc3gXUFaS1JEk5gToLU+LpFiWVsZ/ayZS/87NmJt8
Qrti3+AwG41LsS9CGq38v7ajE3cujRG/9N8d9REIuXyjuenpkkmw3+C67huDJqex
9KY5XHcTp7SCl4266IS13qqIN3hlDdLMgJ4mvvVvX4iYSjpb2jDb58x0pTLgz0C1
W1lJj7fqru76y+yDV3o3mpZ5c+CHVxra5mFEgc0b+zjOAzmZGFlV5ZkDrnCgkEm1
TXvjffDvmHpbDwhMuQqXIjKNEULVYhiDb3QswVS0KQPzMAZmVrPmfyjuJrPylyvR
aNAWiJyBuhpl3Ii2M5BL/VCanQYwcAubz1V6i5UYcAjDvd+fnuUgTVMqOoXQzODK
Zbj+ci9qPrZlwI7KgztOiG6BXNW0PC4JAc5UbJnB8WUAz8ZKmE8qKSqXXVoWcAJj
e+LkXvpaEa2JrtwEb82ob1P3geNaNpoQX7uuwLlH+qLVK/HXCZehbTLIM0a1S/90
L6l5IT6ZIgthj4nj3olFHQinuaL2xrZ5eQN4bFmqQLcc0wZSFbFNgkTgjq5wSovc
YjDnsaoFcbFt2SpWg4jO/1/QIyPW8bB3p31UG6slGu1t5CPPpRQj22TVCS6q/d9a
4mfRf8ewg8+Sjz2j3m/HMRydvng9jnnkGWjA9h5bqpyG4TfFCxgP+FyWjE3Yu7J4
OL5jAkID8/VXJSnT847HldnipY51Z/mSbZdzr4hTVpY6DYe6HNQEqjN4rBuspfJk
QsmvD9+fBRiIxGOH3bueTl3hIxuMb4ArdLGucw5kOUNbSx78YetRag8nxnzNfBCg
VbCjqFTijcQFmiNZV+HzjdBFi69SI7K0bS1pwf/Tk/ToWW1CGxADP/UvPOA9+1vT
231kYN0FZaf3sJLJ/Yq+gthjPEXezzrRSPfznZCFrHx7nsTx8PLTy7macFmC63Qy
4euyQKFKpsZG0qwar0pLb1NoBsc6IzoaIEf4J4rBWoodZMy6bBHtHd6mrR97A185
a/MRwwFcb0flGMZTtepc5U9hwWwAT5dosEwzt1AMFBETBkrcVlLAXjJ3CbrNCfNU
7BRYs0AjHTXzCg3WfHnmvsJyzfpz4/ggf69sbf4qydaiXPKC2M/QJosMqtRMkxlQ
L/ZugH2jh4RR9yzoXPHPUGnFf1mEra5cCbTlffp/BKiDGr5ifqwBneupBD3XGmcY
ZTGe3m3DC04GrVR0daV9cyOGE8salZ6rCzD7SN2pAyPM0T49WF3y0NXS03ISDMMC
wghw7l/2x5kjpZiq3owMvIv0AZahSyY4/jkrB7Wr9wYbhZbSTixf/9qLek7VV673
WawAXMOxjI+pEbmQW1uDVHGcgEhsC0BjYzfhjg7nb5HA87gVayEC1BQuCLdktl6R
IhztjUdDk7F8xCjrGTmH0YJRYA/HPK23P271GV3haOa56aYXemAdLu4zttlabX9G
Pv8NYT/3r847dlAq/gNwg372YaMRjteqWhrIxCMwBP1PmtTwyQ/5RJu2jobeKB4/
rlt2F/Znoh5PtB0IfIYYa6Fe2UO40XmOsz4PS5+LPMH/x0gqboMX6wQgB0M+Crmr
7WE1RrtO4FCzElNREQDgu+AsfY13xlw049Ag2ow0lH8ringC/Jt7bNyLbI6XkE7Y
cYK1c4FodSu5lLZoLxdPqPvGRuBytBLO7JG5Mw8jBmIuY1QaRGehZIWQyRQf3hmE
Z3GQTpKeAYh/BnQATDoxz5/DYRFEs8T/JEe0SNcBP5/rykHwAtDzMiWIiIN/ke2U
nw9l6kwRMf0srjWYCHVmvloJNF3DwaOGLrO+eIwRXUYixA6nPBQ7/tt6HrUYw7Su
2SodylN1lXh4gjrYzUX8ZIMIYrDd5NhaFabzCZoHLBvyKOQKwlLsc0vDcofLQJEw
94hJfgkqZCa00jNNZNB9y+lY2Yqdg+PdC6i8x7/vmoH26lPW3ntaZEpMjZp9kmwn
oWb7Bt1o0jvKjuILLWVKRSoeMmzSzrWLEBVuiOgfbQdRU/N032Y1CKQOY4hwwrrv
L/VhxpIZN5TjjslF+K2B3CeaDFLmZl8Tl85ct4ts2X97FGJkX/Xs4R63gUimuYDn
zcIL81RzFtt4/UrzHec9O28db2Gpw7boUuHSXwrOafs25aM4fA5nRd8cTSfVHOWE
wTu7WfRQuEADkxO9o8srERtkq0jD9KxPHqY51cj28dcQRDYzVjqbnIlxa+3StVyJ
Wfm95jbCnMJGYqWwlgyF1o4OckYPWrEP3phFxWi5Ch6GLqwDA4vQj3Mnz8CCfAbf
6I+2JKpv6UuMxmkXH63GLx0v+oqkayfxb78g/CQi57B7EpdpS0FnIKGkaPn93LyR
KDm4LwMUhyHDkZ4ehwR9J2Jv1Pe9QiJBcsWqBShOXPbHiJmhDrN3YebY2r70VZc3
A/7nrFU62itOLgbCJYgfu/QrB0ZrVOqcAY9xLD1S37Ye5nkFEVGTNWz0fUtf+Ct/
HTKBDRHhx2t3xp7QHDJX7c1ilILZLv5YdimJeELOlc2A4JloIfuOfpqHYsOZN+oX
upSwgwao7nuhnk961m/FPrvlaY4kQg6Sjor0r4Fdsof4aGmOedzALfk9ln2xeeLb
4Ak3L/vxCKem5JAp7hQU1PEIrIvEQu9BqSpA4Xfwp5KEkmaNVnBlW1KogZjjMuyQ
1IuEVoSfhrJmH9zPa0PF5ot9Y/hVJMpHYc5JegQ2WdfsRJ/MCGY04xCVvBYZR79H
g/oH2UOF0RHW+hCoAiKV3k++AYyFBW5zwVf0Spa4NbpHOxmFBiwdOIUd7HI7YQic
FyB9Cr2rjo/a35bByFVfunNI0VeL6EfaJKVLi0Dsa2bM2X10zzpRudeFphpa25lr
cMsVR6ezHZQSOyyNS9viHhpsRgNJ8DkCj/S98k7MQvSJBY8ugrYV9PyaUosJKcbN
a8z4TTy50RIKbwpFY9cQoFqlbiVaQryAdrQfxrBBghzgPCIOXOfReviuTti4AAvg
m7BlXNTRSm49i1WOhPyTllWzSL1icI4Ko2H64LekofJ7edoDcOJrB5rMYOd+8Zer
a6a6WAo9UeftKaeRORw7j7PcmY1S8rWZ/XJyD/0t9INQHABv0Rfvnafc0hNbyLaj
F6sVWEWoPj/g3O1pDqHpmjX8cILwKZnJvzfut8iMZFS7wiOxVX4sVP+6OsKa5fFB
jsgf6hHGSDSj3zvnqfBYr4+tFwrUVIYecHRIPn4fXTl/KAtKhohoAjAmsmjvqDqD
lfstGH8v+/Ifeu+gEFmkjQ1hvrrUxy0p9FB8+A3BLJRAMaS3zsU7VQGIRfTrufSR
U+lXzbls/hhSe1opoVGRhbE41XCl+WhbpGy49CypRCMbkdeLW+Z1wr97hKFTYAmW
El2WLCmutJVF46aUKmREJ9qCD+VEgfW9H/Eeu0TOTW6RMmKszdvfMLP3Xe8wZvW5
bFDZUQ59TQar2wAM8HQSwbaTMS+v1QsEnpur0zBgEAJJ98ZQwVlTsx/wSKhrgTjP
grckmyhv8P00ofZANLjWEpryyzmHhRBgLx09RIOQsw3t7rd/OIIdTHgbEHUuiua2
CXUiy8LK0Xg7Ne3RPkZkUhYZZFfW6ammjYMOqSqzCN8eGCXqfR1gOvbza6WVc7eC
oCJ5tPyNUk0P21DlH9KiH+6maSmKkX3shNesEn6o574mT4ytZmCHl4wmEoGlTa3E
uYoKev4UAsNvRuSNMNI7hG/RaG0FB+9/PI1Sn7Uq/Yda8fDcN96RFr0PQ+VfV1lQ
zC4zpkwrECyNttkgdih0dXfkqMYfMSQ12PuiyFq3r15KaprWbKtKHiYvdoKkMqfL
OSHgmwBOGw5jaGdhhh3PszvjceBBA4Xo3uRv2iErK0lRAApfQhOvJKZ8LFpJOwYc
vglBN5DlPri4se7Lbl98+wznxco7f2czqR+AmuFgmUrJ25kmYsAvCWF1zfOxOtxf
DD1ajAA2utT+8MYHPMQ0LzJ7BYjUN4XtbsKynvDXt6U+jHOlVK1+EwAUWA9rIpsU
bUWuT/rpvYWMcpuCMpNd7hK/dB4h5x5yNxbYPHbtEF9ii28yxxfroHQYEJLFsZye
J6JEceKXYSgJm8FUWEbDee6kr75bKO+Y3N+m8s7WZmfDmmokZymdBU2OKDjGBSL7
TlCiJT6jdaipTFT17WOjuxgA5T3SeRo7HT8gi2d3fMAxao69rFPCI3Ign18BV9jY
NQCk7qxe55JYZEwi8TYUaD+xUvMiRYzVFi3gS+36R1PnUw/rQGmceGpk/iDY5XqU
eeOZdMiDS4wD0IojQXYZsp/2mjm8XP50Pxs1PGmLbZx4R2aYG2Rx3UQ3RN0UW5HN
MFynEDnUtQc6omIhrA0JGWctYzXnKiBCyjJI4HKo+padIIYBarGCJ4oNjdwSb6Ud
O/xMLF0cjjAcbGXGL7rZIKlexKhr3P6ZjTEgI7MBbrsdFAwMU3t6JfkbLFnDJFoY
GkPBbB8zdu0mRLJpXSduGQEd8KDn1FWzx8tMkX02flf+Hm7FmL7Vb8ARZSMA9DIp
w5wIbwOczdsd3lovhUCQQMsNvFp2aXQt8eaXb1KMbLjr5S9H/E4la/JedSG+gKe+
Jj9DhcGxaRum4Zdtr2k8ovinPHWz0VNePoIjJfFACaU85+cZfmGIJY0Vvs2wIQ2f
f3O/qBkE3vQNnVHO7fufxNfP539BiGpu7J5t6ADurKrxBFJmo2RB29IQGTHlclOo
REZOC99mKtmwKhr/0D8WzvSZx7Kg3Sxy5G0OjaasVj/qoCXkPegfxCy6J8aQmSTA
hqZdyu1fEyBoOMreKEDHlXTxysMNSP+1j33SzyVZZGoXK5Xv4ohsXg60/UMxwa8V
mXamok8sQTIoq968NUlkc5PzzVMtRFl3Fk4uQWVZlPGhExU+SfVAfDAGQZLQbyXF
qktRRgoTdLAg1jkERmk7UdlxQxsQSLPr4fwYtaKMDW+bUuAuo67myt2TR8O6cjDk
hJ4Kyg5LrfcCBLVSj85rBni9BxYWpjihHRqlP9vI8jwEflOysTOjeXC2ahBo35qm
VgyteaeTcEdjp5M0OfPsFSwY0S2kYS4TBy4nJxUrLQsA81Ek67eQPZFePGzr5l7R
XZV8VXjxyZNInr5kY1+0BhIva0UsxJiVj156qGZtztA7TQDJ52WRDsH4+au+Wt7J
mEGrIGCO1xr10jfmaUDHA01qKTK7C/eNT/DrulMO6TuRpasgYQqcLAG55w3siG17
NfqGxsh4GSPmoKpPUOvhbauX5sZ+Fb81tfLoMoo264FSy4bee4RUjWowqKO44ALD
L3X1IFN/MOz+61fBJyK+Lvm4x8S04ljqvyLzpTFQ9feGiOiTnhMIJvlnrb3wbBi4
uZwU8aZDy/1rC8Uj+k3oEwoZ7o0ERDXZ+oe1tf0VCc/zZBSUpEnw8WbgKTIsYmRx
63FUcyGSvg0XmYgGOFr0qSUXyGgK/4HtX5fujS9lxkG3L0ySCMVky1dXsI4/KqjU
Co+2QSvwRpt4Ssz/FaJtA6e01NO/bj7Tz+kI/pRDfgSo2cnz87/vYKafxAzM82Fd
uBqlvLeIhrw3b0NDbNztw6kKOKtAHETK0VNwooGi+crSoSkbzR7sxn0rFNo9TYoS
xMXqD49ALQMbbyUaU3e88Um/VY46fqkosn5xgRMNoKyXEKNlciR5srAbSfQSaNih
591yY0NgMfxaVWELj3qFsIwwXAVDYqPQpnsLarcmiqsc2DWRtE1eDW4tHJu7+x/m
hYDgswAHPgvRPqnt9wPtI2d49LD8+5eBD5rLrTkR0jAAGMGq0VjSUiH9L79ApMhl
AR2lZt1hrtaHXAwq9dA3N318vFeNmZ5x1VPnY5x988kYIs7NlhiMScgnA/4oANPy
CXKN3ovMjCRpwOSyzpw0V83AtZUJ/jalrN3Ko9cPcaOTKoRpLLx064XBtXfNVJby
SBfx5I0ogKT4zK0zkEEAmuFkj7plKLf/MBLCRtoRVLk+0VFsxQlNdp+lo8ILxtu8
JJ2TPJHMA5q1zymwdSFYzzEkW/n0pB10URXxYL8RSnkLq8ycCfO6mBrniDIA7DjJ
/mUBK8uhxJRd4jZN0ah+k+MnSByz6akjgofHwZgNbk6B6cF5FIzJHtD9XVdQNhiQ
4rwLkOnGetddInU+6Mclsv3eQJkCqC1vBsMQRGPJ7M5IxZXCMc3/8zjTywyHRw2T
HPTc6N+vAscwzB1I13zPDWTjDtlLqrTTarOoHvKda+i9FeuMUHg970RyaHT89YIG
PnbrAoQV5BHZIQkqwlzd0JuOrTQsYkfm8Dm162LKhOhYFwqOkwjx9KVrHbXk4aNG
OGmTw2oyhG5BKld4DxIHAfd9CSGZCv/NYkqtMP2kx0ifBR/BIhGn+uha5DdOGanl
UqqxfqphFVicHI6wO9Rnx87VNNMvqe5AuVlv9+RbmQzEGxedNZ2AYcwI3oJXwhKe
PO6HbwSl/CHH5dojY8muEYwnaahpfwGCi30NqW6GGmcCZ6CoXnyI6nTqBNErRID7
jpLVQX+6NhxtIZNpp7n6ZGJCfTF10Ez0S8+onnDrB0Fr9yxJVEMGGHiSiZ2xtasY
+Kpp9o/IMBJDkRp61W74rNa/ZZmToAkfsqm9/GSdhMbJQsqIgkjvbasO1WTRYP8a
iZk9Uzgbeh3cy4+vWAveL8DrgE4Cl2NRrCMl8ycO0MCP2TDu0FS43E0q51YkDtL8
0nUDbFW/6TCmMiMzY0ilW+xJD8Ouw/LcMzOe07smrPbTEdH02VZWO0Dz6UlaCvmU
PBqBj4JGNLvyoAPQTNwbq5vtut6wHHkQ+gCWTo8RxFG3ID3akWczx/bB2/jsZY2j
0DW/wrkKOfg3BhuI5GdDh5tQ55nGVn8qpHk62aIZfAmTKMl/TzoNHXAXETgXq/U+
XiynWUGlLWU11prvePdfQItckTW92PRTLZP4HGcy0IOgsmV0ETQ+VUlfUhOemFo7
liL6IKYlG7Nc1I2LBdnJOX6jORLl7ava0rdBDa7/sEC/PqkqR9cy2a2G2r0vze6l
GsYF43ud2UH7uYOJoiBkMJ5mYUTkAb5jRUm9y/2X999xIj0eJH5x7xE9x8MNI3qH
vZ6l5ZIArxQYNEzPXTFOo7MMAnp4ABNq8KZiZdubkTkyUD51JJRR3EyRuLXBfAAx
IMQiArA5n89lozv/ToLB+gYm/Wm9uYDSicZ0U+FM9huslghXZDdA5HcgyAQQ+BIf
rfTMfPC8+jsj5TK1CLgAET+NP+KVNl6uuZtk4MrUZFt/11714cTxKjYd6v9vukEC
PwG5tJRKLk5q2i4xjSzROkUVNjWQ8arcDpmy3QFI5T7owefeQPT7KQg39PWLd0os
t0mRR21UeJE6zPoStgCAsJAcVOoc/RAQ0WbbdYTXHbdnrdw0SRyl8VV6GKqt00sr
7XDiafhFfOHo9+OG6xtbnXFr7sS34sLMjMnlacMaJ1tbC9lo2Ggngk6fwsFZpaj1
7SeTqjqeM4SppNWeay+UMiK6tKWL8hbYNsSE4iMmxsGgCI76ihPsSaaNwzu/NS1u
RypGdf+u202RAvADL6EItuwFZ7fGmgA+Lq8K+kZzmGClW/0H/KV0PzEX9ujAHSt9
a4AKiOcxMum7QkAdmHWBpdN5DH9JJqDZQp92FEHih3PNOy8aTwuTyYUrhAfNQRWo
RYsjv+95hWfsWS/PEr85QPfDltnWqAIC+8m79zU75cYuDM/CQE6YtnIstkKkXzgG
KSIcujcc/4i38Eb9L28++mhXk0OaWJCrPRu9wgTw/DgISmfp+c5djD6dkr2A23ed
sxtgsQdTxMEgq79KNBxjrwkdUz9NZ3Rv1ValhcpQXFLkfmGwulq0JMAMKZvLbHHO
OJrlGsBqbwOn3FO5VQbuUjHb7RdvcAbqal4tpyBD0IO9+OWH4TefAHcdnmsKjGYA
jj/k1z1uOa492tyLVAGGXNBVnXcQObYvVVDrkl4tcaZwIa3cABBuH9KnK4yVJYDw
0NtKiXEGlR8JCyB7b2dizS2gNMW/mKQjKgOV7DvaSsbuazzpuosGnapOutNqKty1
Vb/Jzgi6RV15D6Ap5qXYzruJJKmkvbQCrqG3uiQLzJq+9Pqs+E43ATTnkVJPJinX
jxAlXtwh4RtLKBq6oKcO/+JiVgrDnMvlfR/4ptQe77o7EQ6DX+90i7WWo4JTsABC
Eqvmj2AXfGTmZuZ3xqheUX3YpxPAsfMfw/c3IHxrGYSh4ATYHZHgikNKcmHprTG0
zowMhBPeXwM2U3OZJInCo2ddvJD2tYRxb1gzw2Xz0zVRLAgffyekWFce8Ox7WWRp
DHb8Ga20B4mtiH+ZHAM8uGDYDtZkaMpqdaF/npaDUl9WYFEx0fjCJDrf1ekX17lt
10Xitb/yep/bf5nKOXv/3TYp09J2OROsreySWNIPisF+U3AI4TL30YymAuWyniCj
WpKweVH7fLMewT4TB31ROo1Mr5yU5auvUrlA8XhKzkuv/XaNa6J6V8cBpGRvUhqH
3vtKkk5l0piFJWRUwgdjsKvJEYGC2V8hJrA53KflX47FwBjlW6u8M6jfmTZuLGdU
D/Bx8HUlnS4omm8LRhHLeZmMMdwxoeOxYuzJI/0FXZyPMjRnVDfrRbgFpJs5zO3+
Qc6NYRn3oeJEv/sy4v7uHdY2MeR3UwAu7fpABZRXe9UvBlv1d0vcfVsnAX03EVgr
OfORmJT16LY4tknIumscdNlxICyEr0fzWTFDgRtROMFAMjNhcRakRtz8JE21w9Nl
s8oo8smyBxqtnXmUmgrnsMnARH3bQCABTd2jZon1HAIx7DYGpZPK7lOIWKqDAfyh
QYg/qxQvw2Pz1d6xUKPhzSO/LUNsG0jTtZRNvAM9/Wz9nxTchsCy1yLmWTVeOSbM
/CyM4Auiw7DDpY9Z5ddbs1sxd5erE7NnEQf5hbFbSPNnkgeaZ+r8tXBv0ZZ8B2CN
7UkUTzYKvHMhoTcon6/bp9ROMs0/LPLVOoFZUa05E46nn/xf+W5yrGtN/qo4aOLd
ugbOhttEZklXi+uugZ4futKwY9QPUBOKBttEdE8rLvF7Ge/cb38jkDkfZqy1HesW
o6+8w7Kv+JIVDiGtBdDRcUjqhfLWxe/vn6lnf5vPHBqMdueZyVAWmcnOG08shDdB
rs9dpUN1oFc8naa/xkNbT4rUqjTDExqmKnLjsAjZnZB/uR6eVLkGrJZIMtcqCHs4
DTsEcQuuIgIDTP4BUV9H1wTtO6nz1asW+rUljhzjOzuouGsNCQ5jggX+R8OIlMZo
qbWm5AVPpw7HP3tsz5w73fXNoOlCg4hwUU0VD6yXSMSCNuLZnu7/QBY/iIeyNXIJ
Moa4zcq6QXj1BLZk7oO9DzHHzIudubNcm0pW87coa1gvhV2x8D5Q6L2dlCPlQnCv
RQUd8v7F+I4IlIyMJt52SKn1vzqpMbhK0ZIcm+UeuZ+lvuNsYhhuD3aXNrKcYmlC
GLod5FqpECjAX7hT8QyD/Cy9GHHyQF/+yloTMvwIhE5U1NurxLomAnjtqwN4jpJO
QtKnC4fe8ZvNXiUztLQO5p9/bJVa2JYQi5O+oONOLWUFD+Ndd3ckX5Wy03OiWCtY
5f8KNsHx9PAi7a3Hl3Ofy2VxIpSPk14y7ffdgcT8F0iLk1ASA5ZMqRqrQ+8yxBgH
k/H9xm6vPe5EqFgX5r8JsjMl8G9gvIGx7Sw7DRt5tBE0kJRc98PEt8y71q4hQw5x
n5xYafy3dVJHPeqVB4yC+Fxc+p5CwP1jgaBviTlYjiVGZvNbMwMCHB83GAS+cTdq
cIfjqJTSasa+gFd4VKHPSBdbv0y7AQA/EyuQxi0laOG8NB+IGfOXM0aJKfeDADNF
17QqSZxrQYqbr4oR9ttbV96oKsOCiG1Q3nUEJMtka5obuD3wdQ9pMihVF5zxsCOB
n5M40gUf1FqIsETX6pcRlivs/g1DXcovESSR+AH55nXrfZhWudyvrZsE0mrMqp1d
A+0O4ycQKHDlwggwvWI3iyNVxovx1MGX7TTamEw4OWo7hyRG01sNDMcVrqIGoZcG
6sqDwOI7zDRYVJeEtKiEhs6ftNZEh5AhWOs88J0gZe7riQK71mVlguulJ9mBk1ZK
QERSHsbqAYEqQb84jOTjx8TGBe+GjY5nr7oUwDH2HgYeaXyRkOJ0Wr68feZLGSqU
H7QffZPVnok21xOS6YtFb1FG1/viD1S4uuxrcYJaMIhJVwlgqnJjcAGj/h1OEKXj
HuZdOG7VowcJKfYQps2V1BSU30xY5XScY9hZ17LsgHIsHzk73m0bizlVCdhNTCFw
6IENVZXokCSscJdiLS14aD5oiisidQ2KjSmktUzHZ1FirdciwccXLirLSfoJVmKY
ylPV5r75UBteUnjbGp7UN44Oby0cqZWCHyI4yG73VNcld9bfZRAB1NO1gX7l/1kf
s0HYe/0E3B9g3cnV3LJeJ4Kb5BndYQi+HZtFnaw5JgFimHvL3KJ0TDGs6ktO932d
LeKa5t1CzVsUhhO/s8H7q4dEXnayeXe8FO8OA2YZ3DGDhjz/usd8Kasw960hrwof
uC8UJF4YCVeFZ7mzRJlRkESbuNUW0uhjC/OmHcZraLALfoBhcGlSACAIe0fNmJ5o
vIWFyZ5T524XdjsVIeE2J1gzcaNGamJMR9w02py0F5DqUJjrjuN1G751HqaL0Ktk
2CVRKINOyUxQfVUTTD/em+6qe4w+4y/nFvYYpOZ8DjKMlA+etnlPX5yzkzMBUSfW
96XjbTWxA6UVy8nZq7ffqIM7qooP+Z3QZ3ICmJT40/VTUzjCgtU63SJmG4lfKemV
MV+doCYVlE1R8oZtCGyXfohXW8Xoa6bFBQh6UZFvjHVTbckqUtFSrHdkvzpIHs7m
yp0urrBWia+JzhLGVJotDO7dI5ZNrpsvh/5EXJEWiWJQsZNHrs92ah7rgFFu/SRY
iqojW/gCSOJrOYw04nE0VQfahhv+4hv3UyIw/481YAr+ut2n3iWK/MGof6tpSqjp
9yWcP959OcwjI3/G3wzBDJMD9j9kM/wdjzdytAhyBVtUkw6UWLBJNsvYqV+1xDuw
1AoQuY/Jb6/z94+CeeXpzblLk922XJMNeeAcLK+Y/CGGe/6cUCQQwZTfiR59Yere
44HS1uIn4PCxmS8WpcEfytupviVwEdEpVemel5SFtQnNxXGL1z90/eZOlU6wYjKA
xDpDx3y1Tc9iXzdEbg7mq3HN3vOzqKUi+L7Mq0P3GfGYqr8SqccFMJSgvwKouTYp
Kx60VAkqZNTSe4hgkSjhKMkxtoxAvXnQwj+XrneAJ00Ny7mZWSsuG7cuCRDmlKEC
+9J2zDn2RdzYvIEtkkl4WwJ4epiGu+SOvXnUv+eV2t9qN2+r3XF5v/sx8U7ysjvL
02s3OlK8RBS+DMLOscLFlDAQiwljd1XUjnAkBXxrfqArAx6xqmkQUEeoh2VTvUUI
j0Svg4z4qHONAZVumfQC+aE0lCEL7375ermGTFcYJy9Tp3o1iReyZ8Mqct9jJjt7
iWdVquMAGeh0gwr8MdgdsGUcSLeXTI2HQf51yIVQbqhKkUmJ1FhDLz/OMin2G7MP
k+NqaspJnPZ9tKwV6KDn18QCKSxA5GgCZe2FG4sz17ek87wsZ8/F4dNmgEmLCTRc
HbCk8w9/5qSsBFplR1TszPdl2Np9/d2wRhhDh3GiyfqiTbUBRhe+AzMZXOzuDSVQ
Fzz5CjDzCuPiZR5XnfJUmdKniOyvXJMZXAwcBYvNX197S0dKeY/bqCRXX0od2qIv
7yFP2RwiyoOxulHNEfl0PkGW99yk4J4Bylr+Tfub91VDAOF5F66I5A8Ob400F4a1
hvpfZeAMDWEDfAO5pgebuibFdwsm4Jia2lal/IXN6NJ0Ne9GvqS6hAj8K0v4h8pP
+vZEr4Xdz2YOd+rWfy7EMyPZMVGiqp3IMohLHjEVoRat2RS2FPcutA7zUTdDtQFI
nUCflE6IGlD6b1avhTg2xmtUCxORrthm6UoF9X0EedLPRUA9Nj9NxoeLP4eh+obL
FtJCa/jLSTIWPonHn8ikj/MeVNW1uwNLjRqd6Vd17+aKPXJZm52Vz3v2VRDUPbPZ
9kC2sJ7ctQbj9hpSESWh60yLv4zJ+n+B81KqrJzDnlVjMNidgEJYMGXN6VNCbgkb
mcfpJzy6x70TDl544nLvZer6YdQ8InioV0vGsudpfyUYd89UEhhj5KNXlZ28PVj9
RkQPL1qt8dZNJlhysCD3eBChCe3iwl+H1zyzlGClc9AyZ439WwVUrPUn4KzzoUYl
zEtEeXH/jnyd720RNYzL++jIRSwBsxyG7HNWoz3LgZE2lXMI88/tsJtegI2PXJDh
TZAd/efgEzoZYhjew8OBHNxyZBb4SI/2MoGD2FJLivr3ZOi5cju0PAaE5qWM2Wja
00IiGKs5Rax2G4fpDu1SOJ3SB8c8yggtMNmog6YDHcdU1qwXWy34hXlhwFmODRWZ
QMLH6UQIRPzbZcGXMy2UEvh5+v31rk9NiYLPRP6I5LOn/HFraBVaGYcfrCKhAgNT
MrAt3UmMsUMPM8o5CcgyXHwRa2dLd0/ox9Gh5DNUSyr6M2hwtm0iGSWx7zWsEiDj
wM9NGQ2hZlUyWjLk/FgXf8/NggABELJn7q1EhFJr6wXhI1zxEFQnAeO/gXeIX9ws
EGpxMrSNCYj57X/zaipZgrb5CpUKiHqLUfzCZYxOz6ovmo5XAw5xI5Ny/nfGBSAo
hk96EYzF7RNvO2/Y59pEc7rhnEpZp4HD1LwvLBQqy11qEjL1x7JYsSxMrYRiDVMN
r28H+73yuv1VYMIu/kuEwWx32CplFNeBu8zty7d6jIIVuPJuh0k+XT/BrJG8xlJ4
lJqHJs3oZugVSRqDvnueseKOZfxUZhNjXVTts3PRpjed4MUqcJbGZPgr4nEhTMM6
nRntHOQr2R2Ng8G0Tef9QYFGYzBDC+erEIpR7HaAFsVqKA+57cmpwaG5xk8Fo7B3
5KIfdyMSerF0a9DCm1B+/cg2Z0/S9OFW8JjPlCDhAQu6MLPbZrUA7IN7ZTa8RR7I
jqzqkE6kyzdSZKCwTcmEO15dyeroxTOb8dJkvOpR4X8yQHXEHEPxrU7yXaE53YgO
u5RWh9RfFSToZfcs6PLTVWuJ1Q/XE1F6UgEpXgDwEX6mFWXv0c5lEQh3d7J9b/54
XboMV7dykpwERE7dQIW6z9RuKNC6d3vsigNlQquO87Rjwg6SYN7U1EzE/RRg+kXR
m/nsk1NLxCb6vRiM/3nOy+rx+MaTZU+d/4VtOpeEcA2XYi3o0hct5WCzf9HOOtkw
nuk2Yy+0MUWcVESzwJ9/SeARRv7CMBymTT0qogwot4aIVVO7WK4ZTPBfZZDV3HwK
E3sk+LwO9IXdutZ23/bXCCWqY9vmPk8CNa7vh87N/YYRfNlMowYVY3dzh+RR2wOX
ke2FHYLuv0CdQXxhu1MAs5s4jBzRwPoNF3jaoy/OsfMH/1myGev5WWMZMC/jXL3h
FZw9iP3jYHZlmxGfmcW5tVS2/2TYXbrGR69O8dLsdiO1kpWGrskzAEOSGaZGNRAl
zRg18CXZbXbs6tK2322cU3DymLcy/GjS62a4jzVF5c7jhjsTkx+uGtgixUNQ3Zr8
tOKm1G/rctzB8WaOIwiKp1TJXDuWO73Zh4ToW80WeXGmJRwxs8KKVy2mJueCk0f1
y46oASaPDO+hax93sV+DHDn3GrJPpATcoCeakWoyekVTK0GPq5WtWc5iIzprXKk7
X2nwvmSWOOWwbZrfwb5lfWPz0dCZr+7JC2HYzYuE6npAQJYMUoAMfLoNV/N7fP9m
4YVWPTXJtiVByZDF1csGivrSx7rHDG+t1Kxf1jMAbxOUplW30Ja0LAGl7hw4BIbg
769EQ/84Sp8EwLZ8frs51fLVwHt4k3aIces5I22a41/0+l74JxX9MwRJTJPv5jX5
Ujelet2XFe4CqhVMlpXXNxOQDnJasSBSEm0u3+jkNS5bswFq3V5oXcVD0m3igA3b
uLFJgvpcN8z5QLntGWKos3ECSVaKV6jev50TclDjSmRZU8wvBzBQXFh7xTPTOxR4
iRH6vAF+05yFN7IsatAIACjoOU3Xq4N5PRxWn7eYmG1DrJKkxl2daN/fqARe0wwQ
oi4C46KCmqKXSEvCj2WSzoAHLvKo+PqpEh8pGNjy2nG8vZPwMXz5/5AtXksAl3MR
/7iqOMvIgEC6Xpfz6FmwgBoqW5aMLGC7nUXjmEuh+D00otbqqxNS2mX06b85XVua
o7ZkmoXotEFAbzB8yDaVSGfXj3PP7ieji9ky0tY4VeIGVzAuhSijVjORci7nveG5
tajt9Grj/aCY979Gaulo5nXzmu1LIlJs/fb6wIpZ59iKaBEpI1hVhckAkO9jsXch
ieJjAi+5jpV6WLCVcxQ9dEmX4idFiXek2eOxsm0X30Ca7UtkQjZqTd7EY/CuMAZx
MQWX6eEctSEQB+n9CjNZYyVSynBzlM9pjQlQ8ZrzydptTo5DipSFVV8fZCukloL4
rHP00HgbSS2FbNITuOXy1av/7M7YTyWamm29UFDLV4STCLrrKjNl/3Lwx50D9tAQ
+YFfULahloWDH4CogPNs5riDphkiJwS/N4Ex4OXSzVJeVLHb6ld6Lt0DDJf1xsOC
6z/YNGyv534boNTynPaOuZpv+Qj/Oz2BPc4RrlnIAlVT6MadwtmH71R8eBECKEPM
oSQRPtCCcBuGGptAgT1KF0ady5HsAKflIy50rkgUJfW/d/8Ln8VevT4PycjnXbzN
N0y1jNs2T0zvhsOrnhNubhFnmPzDx6i0V+6g/G2JXAbI1PP9UQZ/PRca4Wl1UfdL
06BJMJkyArzFlda2sR+Aqpueq8MuQx3zG2M5/aw3OO84VEGTjk89eU4BxIKVL0c6
oKww3Wyum0AmcN8Hju2cPW4lNHiaRwR65Ltov+PUgjZrUmgk+u61Xs2ep9SWZZTL
72iCDMwy4oNMTP41S+89KEPDWONsXQ0SblOAS1CElMEZbTSRkMG+QnH/vN9JJn34
lh0lIDwDRGb9GMm3h/SFIxMVAlNe998bcTVhgy6P52YcKd6T6R1NfmjdB5dNyXlj
sSN8U2BWJ47XEBp5rkJ0yDqzDLKj8VoVpvB4+x2GKfeBPg+k2btZkal3T6FQaRyV
jV4tr3h8HTFdlDEBmAvvKPLNyJ4jvD0q5PWI8p3xBAx2W1ZHUNFomIoelDKt1DIP
llsfUjLt0ZlqX5RxxAfT8ckW2oppLG0H29Tmjdc7OBfBg9n6mNU8x/kiOuow1NJb
aUm0z3Yd6kYRPTL0FDMFrfowoKGZE29Ula/06V6uSJmMSFMsyGcJUlSqsB9vvOsU
aPPUUkEMTQftMC02N1Stk0uTwUpxjhNJvQ8Ao1hlSMUFau2wl8F/lClYweqUm/fM
j8wKKUKQ/egAo1yvNva40dkNUIjWG58TDsPuPeMeorGrVv//RCexvGrNd02TnW35
C1RPqqh+2iwHYJpcgvhdK3i5mSLgFarQH1T7JWjSm1Igjb7Ol9oNIXU9Rsk1tewR
DkTxQRTlSYZME+7+XL3fpW35zGGUbqLWpgqOJzhAUAQ6Zd7zBD7i+BoNsc6N/ys5
eMVo6GSvTPdyaHpqcTMJvNhEVzXatIy86M9JfhY2Uj/c4F71p8Ewkly9XwQabiqf
cpc0B7nVrjjvGKBosrvg1Un5P/lfhZOjp6Kull1zEJtgG+lyZNZFyDlU/BcDnVhC
VdhsrKxypHp/VyoO0g+SoSksOXvP3OtvF8u3+r6BkrTaMwiiFfWVijQ+L0dGT8qj
RniuWad41/oiF8EkrJZ0iKGpUOdVXe4/dy46d9qLKkBNthft/6HFZDg47pK3a5jd
JXOPSC+f/OlQh+zJKXING0ucqKsyS5Ba4zA1pb0Sx4a8bI2XIdJnOG/65IATWfM7
21SOmjpJp98VaHBrWqvsZ9WgWCLM6Xb1g8jMW3/WKR4c8KM71g3WQtRfg+agNhtT
GugjYGjl6KCBjpH08s/4msS2IDRdNNbqMEASx/F7nFIyV3uGlaRK9lF4IqvEC1zD
+4B6CGP8Ey+/C7UuC5PlXaJ01WBeUwsZW/1+vsg4UCRgzhjVILwp7ag0BeplRZ06
zYpPupb7JIrHgoptrTEfg/zVwwBMZsZMz1JK4qHqkPcw9Kp65PamhrD6O7BypL+n
PfPShYV6hiDTKqxZD5bMFkL/bQrNDcJmo05VjnnEBNyc5ssURQULF+yeuVjzcHeI
+GeORZR6Fil1O7b42+Ehl9QS8Tbqr6rEAH0kADa390q7Zypm3J+sn1rmxeYviAJR
w/RG2pa/IBtMi/HaC1M8DOxfiwhbeSzTXcAmQZ8iRMZUlUZQdi1PJrsCdu6e8RQi
kC1CavF1cOfkPeGKEL+OP7PY5N1D29VIl9x+Z9B61GDn35mY18baa/J52sccAqR3
YrKOPUtxWFq7WvCUWPR601ZtF92fVXyKKu6Kas81WRWcWXrCrq2fIItjbfoIbuRo
6C5w9oTlQOXVpF6BggzYRxq6ugEyeqOEY+P1WWyDHzAXTZuAuQCUPTpTwtPSNj1e
tfF0gKNTHgFgKBRX3UbKmQNr18IYTLDTXcJmMXN+vE7vhiuehoURUcGCDN8x8Nma
tSVzZo4no853yasZZH/WOuoZVFNkGBh1aipXQV31s70NYaFHiAfhVPdK2iUXznRm
S5Trm1cLIl2V36IFKqSPtYlLnEIp6ZZ0/ImHZ04tPdab2TI982cZ2evNYMPAldcr
v/ivGSit0Rgcpkb5mHwkgVvoHcma/lCgrB74AfKP0BtcjlnHuOIzmFTsyfNBSsSh
dWEnsGsbYVut+3XJ9YQ/okxzehmoOykDJ6OlTVAQfJ4uop/rQjz5CJo+ERKCxQOl
jILfgReHZvYuSGvkANVdLssww+ic2bniofBHsXVutXx0q3qnZKqkN+IK3rnNp9nW
16CLhz/5Qk4RTmJB1QzXVyNmz/4GElE03L1+aoUjBM+5ndbenS0NEsxAe8SaG0yj
auERiLSU/4xONyiJ1TitfeOVs81TwaEv2fH8FgDzqQrBW9T3aeCexkPSdx3k6WHj
+wTd6Kx0Rm/XhxjlSgsyFPxsdt6uPL6geZHXpJ33gs1zgV1LMQiZk0lbzBrbfkxs
EqPQUHgphBRc1LDrxeBkYMk6SLJNfuYPRrCqmyB0vebL/GuETgV4GKBT9EK/wo19
bdlI6pvWU260846r+VaH8Msnd/w62XE7JqdT6OiqoOMvwsAso4wh5G+vgH6nZqnz
Vs3aDccDu53GJY+G3CTpZ0TRUxz4lkUPmOmaVuYz8Gk2fG3NkVCyQAnhwLis/VSL
o0G+81FtW5IubdlzONiAPXEFM0W6OF9dwb8D4SX64qS3kRfU/1pvjROHrBykeHok
eojs0+1eNmjLwBwgbp7uZB0nO+bHQc0/jJAuWh99DWKgckk3VAm3GfXWUtPIEnBj
XH5LMp672aicdm/xvv32y0ntKrHdrw+sU7WGCwUriAC/Vu2qUVkN/vT4CkO8OOnF
Wq1xUAGiWMssHYltwxREPQ4UQdbCSAu/7ZXYah5JdeDQ0SjudWocNj3AurSF9II7
OXKcJvSFv2EFR/cVyYxoyQ7wpsNCZxe41Te/ZLLFyyQ6t+gEAKGHcW/uNuWK+Nfk
L1xyQS2ltTgfka4THnVtE/CcXZYIaTAMqZxTa49tb6V/JZhWQUWvJsTf6HSyo0BS
EpuNfekwU6fkLvV0nY9Z3Rs4T9DDgfizO1FzVpP9X31MiRrjfwlNkNAE09ZsqpAM
uNOP7Z1eHEzWMRpvJn1C3CS9Ru5+V6kHObDtMm1w0+32Ng/iP389aPffv+ILnUeo
e6xiZ9JMVa0fX/5gVAuHVvqPQg4tgqHPC3UhPgowTV6XlcFZaUaSFI7VMd5a5ihq
yLaDBdyzntrjGesIz3CowIEBP3w3TvoSKusvwPVLyBxQ7Yr7wM8BRS2pVf7oJVio
m9mQj9IEW7FDAdBW29iw6gDbelnIQAKE9lL2lzWpfPjSj59H1LqOZ0FR4Wm6FwUw
ZV53+8z6SnK/imZylHvYpGOwfS+kCuEFEE6MoQUamg0YxqeJM+oMib+0QswWTzCc
y3OxNxmtzbYSIqC9N+QYSJ2uNsLdvtu2vCnb5ifFuqVl4YWD1n1WgRDZ8bGLG9dE
EvGjbgqI2un+4aAFJMuhqdyjNimHZBfDpK/lcTfvYPk4hG8MdXD+G9B5X6ro6jmG
6D5FTuupZNQtOYGz78mxxAGXggVrV5ND5CK+NwcM5v4MHNQ5u/6lg9kRxvt0T2HJ
12VpN0vPftylz3BtC+Se/q65TO2SXsoHeaVoeVMieUeOHrpn6EvDvbsake8I8Euo
UWTRyw4ah52O5nXhxgqRyL003fbHxoFPBC7xk8T1Bm3Tmg2VYXIjOJY1oR8pSJjO
sb+Syn2NIrNs7yjYXmTSxN+HtgliK63RXIZ+k/3gXAF6hv62i16B5kvfgCUNctHw
RuTJGMGI4Q/cC9EzAMNBvDJNiikTmp60H0CXhV9kL1fdpLO3BBkdLeHifBkS18BJ
e/Ta8D6PNorviiLQRb5lpv5XmAETGegdkKTRXS2kVXrojgCQfzzskIar1qN7/Vqj
7dtj5H0Vg8IFpfkfBkX7oEl1orJUu1yQ3M1utIhtyhNnoekLC6XRK/1H16tH4CAk
RRFnuLcbP4ZYAzrL8oipChWMf8NquoIaS7ZlDkDtPMNNaW7YgEr4e2bXCa8lQmAm
dqkzbTZObGsB/NL+/09mTz9YtdST3eNerFwtpmMxMi5TzxoCwHopDqNcCnZbvCuh
F4Hm4jc+rcvG4zzkdgEFVoOVhrqAuPASuT/4F+1EzKYa4IUpuIYbHrO5TVCcf5+Y
LSSeX+veNEOVZrhKN7WIuhAp8Fa5blR9HQLs2vFS9d8lY/cXK6eqDaNRu6ysC61r
QmovVFHxlBwKo91B2zMS8g9d2ZX9G0QGb3WE6SP2naEpnB7qxnKut6jYOaMlbFPz
7YVE+UEeWvJZxMqKVLoxZtyJgRoyVCGreQdALhF0gNrGg5GuQSRb4YH3pjwW9EVv
U1YjXoyS7Zurv7aKoi8wf2wK+MCcYUxSUpCPepGHYP+gO20XP8KZrFIZFImvtkxW
O6wfuqm6TAyfh7jFFxIhXqzhwg8A9dZhkNEH1l5IUxudTcAhIgACa5G/puprA8xe
1zDiaM2BGgd1GEg77R3BxyqDeArb/aUnFaxKqVY1OQDYXWXpHDUnmkrmLBquJ7iU
/itlxt3nvKa8HLFnc6zIo6qpFSQSLSbyUzyrHaSKhn+k4Vz/R9f8kgDj4TO66Jgf
Q50rl3oBq5a2URncLFJduy5r6Z1A3y+qK3cb3sctfjWShkhXlPONDfc+LTq6fUHy
SSp9BKViFgGme6BOZtTF4zGpBWWkgZVnF7Mt0m5Qeq18fCMrzepX/IoHH/cJkR1l
3sc02aoH4PsHJYl+1J/heDfkMAIWEhCWInKnTXt4NpGIikMS+zr0XuJe3elbxPkx
aCMlWccaZ1NDBWZxr3vq+vJxJXDi5BfOuXs+AopSoAUYr2jY4/uBJske2GP/jlFl
ldzHGH/kTosrjnVzuBh2Tdedg7ihgmI5qRVTKatG+CH/lOMhU9unu6s944Qysoxq
/vzpZd8g1ySs79oauqRL7LVoHoO/c1dzoFkKHhVSjtIPnKwdos/hIwz1+Txstmfp
tuuChWH+/gjINTEP8rJw7r0pwUOrOSsCeHpV5ojqIH5sdQwvJoPFgFFgZF3CEoEL
AJXnurjXNMERddusPb8HqCd5+h4PzNGQimxq0zmxYtJY4QzQTqXilQPwje5l+Cwr
vdh5MuCtQYtg4XYW4B/6RbHoskZIhqMOvyCixAEMf+oUL1iRiFixrIEjOgu5+3Oj
gUV5nblFuQR6jo1HzG5ZYIkNSaDoKM4wEw5a3qpNxKgniooyFCJ8/kNpQxOCezBQ
woE3/r1xDBrBKyJCumbjHaHJjqY5nYbMnq53jYEgdn2qDCi7ybHAw/AHsEhmDO33
nnmIUOVXlJtM8E5UES7e7TrOxxHww6S/eJdtxgYU/8ccnZS0PZ43yAElv9T3UCkp
p7Ag+v0LshE2/vDr6UnFtlk8xpJ+D/PxUCfVKTu5q9yDgRclyglzn8BwsYj+sBJX
6L99LhNgbDf1nLX8EJxz6hKvab6hvb9UvbeNQuutDR7Pme4NiMtTFg9SoeQ7qtn+
5ffpO5ZLFvDtH2UNYhhcm3JpE3igudz+ojAfWi26nJcHJGHq/8G/FTJwvRUNGSxf
IKPQfnXbqczqtEVt6Qz8GoiJnDtnymvolEAYRegw7WGu5pyk4gzBku0JBrxGb36T
hVb44s3ffTsAdTuMDl2eddEjMy8II0ShKmQ7OHtUEnBQVLk7a1NJjZop8vmq0UK/
Vx+Vnlz1tfU+RB5lEQ7aB/+Y+FuSH08EJ+buHXwbm5UOcUgQuG+rw3Gzxv4VzO2K
wtkv2xDHQs6KJm7FIoojJV5LSFS3WrAVe0WH/6D374WErP6syeJ/29RPCLFoGbg2
Lj0DWEAclqbXHAzBVIsmcIorshq5QT78pUyotRcUau8szNdiZS3K3TEKdGNvwAd1
KWLnEDaxBxpI5VQz1XPh+5K3rRRsJiHvVjB4p4eLSpGDCGKf1C6Hh6QeNNOtORnU
fhd2iH3HU1Vxl+DjkjTQIs3Zv1A+Px9+krXl7ZLSRDeQbjQHrTIspTz3UOfpeZxO
+UH5eG1SYpTGcoDYVqVT2V51txqQaKstycGvgrZ/foG3w6cOWSm2aXl3FeyKtw65
+7Zp1lUb1gcqexjHb5hgEijpq59SjxyHIFk3h2jrM0H0z5uqlcQm73ohOhibD/Uk
BQ9l8GikjvJ2a1czSRHlquDIsNtO1jRjSwnGI3fe0ym8yvl453WImF2gPTT3m0nE
MmeHHSWhwHHX2OyCfIINrXaGq2GxN23S6MF2S3Qt+SuaAUslfsQkmzu03eX/7kdm
tidHhwqZ/q47zdIsCXcKgptZC6LBMDws81+Bw3MACNhYOOKyJublXWhFO/nSjWlJ
zkjjZlwIuGOKj5jPof01w0LYJGC3NPFKRpxLU+UImtaK9JVjsXeGIA15mQn1AVPi
+6naZedlIZnk7gA2Cg9MyKywnqDoELb9RgzI6mpmUqZlMGZbyBqo7znFuDlFlb7Z
KDo6MEMpnWTwxZPqLyompdSbVq4IcZg5AQzU4ZowaIxXtr/8X1Fnaf+Ii2/w4iqB
NKPgG57EFBGyAca5PkFb5IbCK9y6j0vQI/sc0x5T/96qpPLZ9ldUc+HfUXHWNZs1
sIGGmAEDN+UUGXeacQ7OFYV0du+pAePwU2UmEnVA/vapo1fbbLm/CxfTiVk5RTzk
dlpKM/6S2CQuwBwP6m+cQlNKLryr9G4vqawd/csPPKKZY3fUA1GbIIggjG9JRPwU
0dqSGWd0lceb3DC4vm0fxxNHDaHcjtdw7HU8MXZaETT1qobBttIie29MbM0mFCAV
+SOaTb3tjkcFiBmRfXtIatwTANFZ+xC7+wQPHSlVsQWEavjaFS0YG/lLtPcgqHov
0sGK84s82gC1+02Abv76Fit9Icr0Lpvnu8ZGT3Dn6cazZHPVXfZbDFZBpXKwKrgG
S5/HzVRPWnSEGj7Oor/VlH4slecerDSAosEudbcC68ioLLV7HwFPHLj2FfDwgIvC
tmEjQHOHNLWIyBlSOrkqXDPoN9y1gVEn3Vz6cJBatjL7mkGmsNx5zp1tP4mtrAYK
PQWCYzivhiFQx7TdvBT892CkDZbkyPJTBJlpSfbyRAf968MstpA/dFI2m1QRnJFW
sDuWZMaFoIfyAIIW0uIfXj8inRibUYUND5DuAFzCawNwgfZybpZNI7mZ2aINK1t3
qTsLElwUtv/Bq3O3o7kWA9iPJrMW4+7E3+trwEAjxv4/sQPNssiR7AwEQVtMkz0T
SOL9HruipFYECVINRPr1ek5trnwVXZBZm3IFCfotYxO5xBjw3dRLTtwaexPADW7E
uy7M9yKqDuEvvoMJDzoCxHwkiOZ4denOGtArN6R5Vi/f6sGhaQCW+JgohUrr0Cqz
bQ41n740XabyA+p4rcIWYJLsu96pBd9yfYaZAhPMQwcMezVoEq/mTiEnQ1vVi55S
9pNAUVTLS6Gubg0JgnuIG+7vAYHB1mSK7rCngsG6tUiGzWZ4NmhABOVQqQ0NUit1
/2G3wa1tKQR1HbDywH1K8eGC+xnRPpP9VjWulRqDkRYai7okEaSfQ7P0V5fYPkcx
msAVGm4QsKWXZFPZI/7IuO/laA/TlL1flhGpjh4EhYWm+FzWuS8zCk+vkLESIBnQ
Y776OFL893sKIQ0nZPZsShOrL1s0zPoLM5pgmYpG8ujvQorAtMy8GFFsMabe+GzC
eYhP9UsfDdCRhcif1Z/fiFWYHx6MZB2SPmgsQfc6wZeWsbMk3bH0CVjbKLrOuWJS
fdg+LdJuBvQ/tfAwCKtkzxKhBHCung/nm/PpfRdLgqOEy/oI7seH7p2xv1QHcJse
QA1owXb5L2aHz+SfVsXyifr7FoOwIBHvYEWAjDJ55VZfUSkxeY6UILv0fPin0t2d
i6q3v/606R1WO6fDMpVkaAYENhapHLhLeRLnIKLqXXgnGtWxaN2ucz8vdKN2IyjS
pZvXGSNw5pZl+KVMBbeAizST++fHkjhCYxtgnnUD1+9UTcOHwYpCF0/d4h///Uap
WbgMA9TVWCt9YjehGXB+EKPz8x7xBcRR05x2JuIZKZCAjTN/PnRWBS1OG0xK4qrh
PYmrqHGBpTBwer+PvBD6l2lx5hAuqoX14ssf9UBGNBdgz21fWzz3HR0xyhp+qyzD
4DXek8gMJKh2pikTD1SA6e44ZSS4eHWq2xkPKfujoL1xz7PrEHO4dYDD/fliZ8D3
lTYZVGsJV2RpsL3A+hq4U2X7vp4nM4XNhmMCTNb+BHjKlvR/geQ+9VI4avFOlbjc
oV7d2H3lME93+XOG1SC9RspCtbBswSh4FO9LfOoms3WCxNFTOHziovLnU0gugWbn
RuDJ+eE01SxeRO0K1mdYKmvFukJWR+Sg/ieTusXbH3k7zyJe3NZtfDzGCwZx3mrR
DHew6pW0q6c8gu5jMzOVpiSEU2E0Y3F41+/RgwgDUa/ntgiWEbtjva3bXPGAWz1K
E1iedn3xcNgIQ01nVIglEd8KWbDeF3OIvVLDdWyg+SMLspBcorTApTmScET33Rji
3FjDVNbW7SYegImTiEhGEiDmvUD238dhqMwOt/mhfwyOunNMjq3HrPFm0HuI0MHb
l61TWBQ1R0rOajm4lDX9qiCqtj56Z5FKWuP3uIeI6+GiGoHIyh4L5MP+sFN/1UKA
t7nvGseT5GnrrAu8pHorJiqUNQa+weUbG/XEs9DJQ86C7Wc1ZLCVzx3SYIGhC4LC
Vc1B6TlhCyLPmNCaPHzFLdZpJdovraVdy+psOGaDGk7IMorREVTfA+i9DdTADUtO
eHs+XA/PPtymke37FFVHqbA3hrn6EovEueSpWvf/EUIKJmnCk16UpfBT2psnFzUY
scBQP8czuRlfrdPgQfwWCsZnKbK5r2/QvnzXKn2zTb3AFKE/ozXyNlCXWz7Yre0E
vPpQ6Mt+A4xTkaLu2VmPj7a5ZtVcCPN8hNhrb7vq3E8lLzfig4O/ujbYfIUrFxPp
B7WgxKO1j+vhsChUJ3Y8lhfVhAhsJDjdutUO8EMFW7NkfsYghIe2MxyLmUnrF9Xv
QI70lx8DevsgyK4aYTJD7tj70OfEfH6J3l28e54Nfu+cruyIm9s+ErV3heXpMgZE
oPzYJfVHkKob4DokObh6Ud61Yz2M5DuCJpl+DR+4d0UkiW0vKXnLBwO4tdNZdup/
I7zqYyVeJ2k1V/KZZwpCMJJTbQdbxxuSBW2PHZas0j0vzhYspNsMtChJJV0hLSlM
3scWsHY1jRV/AL4U/kmNBYly1QQAtBuYX4kc7FP3s1vf+hY0LFmgV+2qqnmlUvdK
SAhZ9muCoK/sBZuxP+3nq8P8NGphRwcV9kibW+SMexDGflBFY968ELn6aO7srPsf
TjTFIit8EBEU7im02fF3mUO2LqLgsQnuOScM3b+sM/hLI6g71G3xTcxGJILyUT59
BNbQX2oxJrfGxS/tj+Gg1ndoan9WtwEl1pfTYQUWj/vM2K9QfNv96vH4Q/zri1CI
bX/7b/D1tPb1jnRUZGIG6lDmz1kWKVeRaF76bQ3eolhER+6DVidkmxfAaq/oSON5
6lkBjhjNLicCvnkUtYaF/welAZEGcF8RDVg5RpuEs5DrtY59Y+pmgHfqpPv0uxBR
XSzwMCwS0Ns5S2QwFdYnFsSKuzZTuLHBGzwXeeAzDNLx/B+b63xVENK/0mfH+BGm
BDkUeOvJ0HdjGS1YbNjnyzy9He6uwLEY4pe9e8TGulB4BRCk21w/AQfqCBFWXd8l
AR3/VhOgfX/Escy21W3t/SrdEjC07IyQMmA/2xjzgQ51i/G/j7K4Is+SFKJt0XWU
Txm2zNpkWTub2cDFrnspNBiDqA3uPs0MT8vzZpHMsVMnqnC4swEtPzWhIWD49W9m
mbu/IGdRYKwp5p0sbb63ZAc27EmguFberbucrMJTxU0bvg7c2a/YPQge+9skD5fk
pzPA08m5oM6CPSSPK4kRHtLeAFvhYkaIYTmxLA0/5uqNa03JOzv9PpFtts3048bQ
/V0cbXkYkmQzn3WlT6/88SAi4w4Eq3lLGqR50FU453Kpjg50vAy5puv9DGKsCm3w
GsuGpUomBKJJPYNPUG9L84wNuPuFEnxlS1dKJcLZ1EBxrn9j+IVdW7qfwHWha5Qz
BtJrcgH6rXLzSBcJLreKdyBWWLvR3/AujUptNI+2IcvjsXMuRKJ+sec4a3lRUW4X
LxG+mkraRg0vVrE6RVVwUIHtagiQByD5kMYADoQE5TpBVPsGVY6+3n2QX0+FuFpq
Hhxm9lMgpIHDVyTLm3Zzm3CnghFDxazNGvtR5ZpaSXXzjOEigjajYpYd2AvyITC8
rFNlbWrMIL1GLYIZbVNET2+uEGtJVmwqMNXQCP+Ye/JZAGepIR1CAF5GabZjWN0j
rIeNAJu3xFQbkErrPrPMvLGV0ha61+hGoRd3r8I887Y5vz/we52KgcKatBF7bU2N
ZSpUwTM7CTvkuJm07HhqpOcNWb6AYOnSudh0+5jG1Udlgr0k0+homt6KnMZOc35V
RgzBX7+zhlL64/7FrsJRkZjbAfK70xhZHeoIGd1SeEGg6yMGkKMn7RbkNaeFBFZl
2GBUWn5xJEfmLdx3tHtbM6Kmk5oka88xLaOiTD38859ZSkHfLU/ZjgFj0BHKT2X2
yNTgjVLxknjCv6ivcr1kUCpuhqXZbYSk2tzUmjx2foXwLYFTXBnGHX69JKw03Iu1
xlLc01tSl5mp1aNXjQcjW1Ky9rUb0JMqzlI7kiaF4BE2ujvK+0ccQCmF15ImxBfr
Beu/m/9WlFbBg5rXQyJ+WBMYJW5kE0mEsjKTf5G8x+4ZQqeEBGGn7/r4y6jJErhk
/8pUkAgVUFcxKVDnmcWDNDIKQ9wnuOCfm1utD5WW25LoiyyEcNIaWsKRnmzaWTUm
HnBRRX0m30wjJlP/dHVtYXNF7DVnLh9dFr+U2LE/S6pJl5skPbEj00jyExO4ThnD
ZHAc9d6n2RgpF0tuomLMdXVvdMdE6QotAl/HiPhBzHjCCwW/m+PFgjlSb1DWTvnL
T07HwDm3SjbrzcC+pt8BtUBBX4aVc49ZgHwA0NEbUO5wQ1JazbOQld9u1Wd+oS6i
oz3S07dVWS3RcIy4pvif+f2rfyvn4gnF2EfAECTOFGPmQXKK3c3SyK4nFPOIAZ0C
h+n8iSc9lW/4s68PFvCavDrNUjFQA2Yy/rpOS+0JQxK3HZf50YDJOYchgWUC2wQ+
1vb6sjB9AE+qVDzaOIliXfMGgJHlO3fLOaf7cDN1Ofm3/uq3+vSQPx9KPxA6OUx8
vKO/K9Bs92BoFD5nq+K8sHv1dySNAiu917GhaaEt345sbQ0dm6AQ9qvWH3oGG95K
Ebog/KRZx4BA+34EGaC+14EWJyhkrQD6zBPJLDNf/gOeG6/iWHGmw7l/3/aXXirJ
Fatmj+nI03dyT4jstG1ZISwwvVcEyirGCTGurln3NK/GdDoB+IKUWvGnxwR6tCCx
ZF7RJKvLmU6YJiTxiHFBDcSr+72dSXkZ5FL9oP0YItbU17WcVS+GKIE8AgUCOJQj
VbHktXupPWUaL5woV/R8NA0CZycjnHfoEf1PKPHePg9p++yl8emcUmQ/dNu79UPW
rigzWwxT89X4KVeF+9C25J3zWQc8IphfPwH/K2Z5lF0F5QfLMGa66JVR05DtLS+d
P/1fGdF/RHcf0FlanuHhUdbVOJFhlAJjqbZBNBlc/flmNf7mErkbyKslywjK1EdM
s8SmPKA/WvsIW8EdRlc3OJ47F4Z7mgL0I3nQbX3Oy+4+zDg7GjLkmiHUgzu/BDq7
UCj/uRGhNFL55MRrOIHrQ3y5uQOgHJ9GVFW/LD075nHaOGg3tfi5eF5zaUYQ+9tG
MFPVx3ko/hxAAwpO7cjsing29Ymm9kU3VlVckY8cGaSO+qvcJwQLzFeY0mwRUblS
m+dPuP5NjUkw4jilWOiwf1kFCK+PmY+5jmvo+5iCsui6m1sVeuQYTrFTymd1uJUy
72e/Iwut+pQfVlQvaX9Cx4Su2xI0cj/COXf89W3vtqKI0LXIPjJyHLdatkcBHgvn
Qxd0ZTDPuB+jdhSAn9A13bwl+WmK6rp41POvqMftESrQu8Y559e0iAfC+5MfTSRq
32g9lqEdn/I+Mg8XbQ5f6PIQ/u+rpas78Qb1+T1WAbBC69qCpwFbKo8cPsxp20PM
NPRSTMKeXgC82rInwRgaQgljrBiT3Wuvnilu6o/zwrUqFR0RVgRVhKW5RLC/XoT+
OqqdGBBRxcSyNyalTujNp7wA13Mzpbc/zcfMeYwClyiPAwtQZF8ihTCEhKY6xdQS
3ibSAfeFYThRISoQW6RZCVKLFtdPPC3VrG23N/HkFC8g3jBgreglELiwLQOiKOOg
8rMJntJjZNcmIQkrDEl//38OUrPAS/Km547TWasKkT2N70Ar+RTHWd49b1VjWTPo
T1ymYFVqaN5ITDuZrYFVN2IGuAowRHsAmovE/xzDRG5Dh2loXu6BZWnt/bHwv4tZ
9CJX9yyOH9NKMY6VZLBWv4aMgbM+oSNwtzfIptpDTYFJQrPiLAfZS0eQVcjp0jt0
vrBQvpPYc+LIE3cLwJspY4wWjD9+NdT/g3osfKtl41uU5/inMF2A/awTc1arFqHm
5y9FjJQ2p3rTP+aT3IpVC/vdn8flwEoHjZmV4lGO7TwVRtVz768QnbCDNWcUIJE+
fMg9FPrhIAF5SbIgd1WHIH/8d/E2dxHPeo/wQHVSNFwGgyA3/hkLt7I2yYKjBQXI
znJFREZYSSPDZbaw+xKQJt/9SDke9jARzNLSyGPjQUQLncF9kUts0LU7rGFYw3oJ
eCTmsWuHw2B6ldwssdsFYnw2LnwGtyB4tcNn84oGbtXbGBuKOy+tRSH7k4rd5H4y
E1+ZHoVM10yRHWUG5FwqlxSGtUC05XuR7ZS+J3AKFtt+gZuDdNx43x9OXJ6HCgPF
yIi/YgK++RfbL0ZuFGY+RIZvuFWMx05Pf4/ss1z6s8bynVlEZZWBTgO5BiSVPRVL
GLF+2QOa1XffUG5wK6mGnakfHL+TX41luuX0yJYRkiSc6LKqlBKWJF/yIBu/ukxT
Q1nwjUPKt1IBvmxZEvkhQwbII5ipp4lUv9QYmDdfp+H5d0iQPppWHttvVrsQ6NHP
yGVfcKHqM49APgCPpJGb9L0WOtxo9LI6uVMKNVnE0iKUX5pljnwodi62FLVMmKFl
YOJHXy+0+SKkJQRRpjo5NyzQEX7MAlSehp0R6FjYzWav1Z54Sd1gwkal3+MONv3M
oP5qhUa2g5yk3wZCFaLbAOVtU5Cym8HcEFAFoO+bfv//saE+7EZtWA/t3WplXsaC
ttFDSyllAPHKLjyiXOIw65T50nVq7gzfmT3LN9BgfXuQwibCnxw5lbhT9165rhdC
+bQBAwMA5fg3fY2zS7uT+UE5ywnxmuSFzSb43z95OxvxhWXXIIRI6lF7slBdbwXr
HJcgDQCWPtJox/6Xs3OpL1Yb0nLgWFyrXmUEvEWod+D9cK9izBJD4dsCtIsriNcn
TqM5vVdoNsk9Fx1/bBHVt8WACqAyBqAYQd4JjsdnX1E0MknqdZem0ZdWig34goxF
7t0yQz7VUxm9ciAluXMtL/+gbvOWiyanxIgBNfIE0YI0lo/PQyam1cGBq/JRJecs
C4hYxgUdXz2USlHirmXYPktL86OmWdmCSkP7bSStukcqf6zj2NnvJ5xiK6IRSMBw
e9RlaJcXK+7klfdHkfCQRfxDXZ/Il8HZNktYP/m04Eb29QG3jB0EBmXhRjHSqUw4
1y2MAmVw1/vMtq7wq6VKV7+KK2eAy53uwfuV/Bxe9+hf+fDMdJL5wG/GMkcbKtnn
gntKWFBxD9EDBRTyZIxbAgNFVDv+Vd6b4jqCqv4rNvH1Z9pBBeFEr4ZUftKt1d1E
mPPgO15rrNR3JEC0MZVThKm+GwwsHTDI2ShknhWX/HuF/4WrFuK1m+JaUIp/uz1B
cOX/908QLHRCeVoJf7/hCQq5pfzs1mnaByUQaSiPwnR41bwbzK2osIVGz9oUenin
X9EavKM59RqdA8KdmcZTxt2IUiHuKimM0UovPwKrbuugY9qlqwrrEXTlxuQ8bVuK
aQzIgXe55O+Td7ATAQmcFkzvJg8qztVpONsTznK+YvWslsMuJREKF2KTQLko9/yw
5vDJoF8h+7p+339wA/98heZRH9mArGmqyQnac36Upr+Ro2jYYwNWjhnK4u65kPmQ
lL+/tJDr2NBu6/MPrafFKz1xx7oeaSi1O+0yjTmlWb9aOoaPiOuIhuds/RrKMrBO
7RrPHbQ8/XPgpnMMkZxDZVjmcbZnEAZW4K+0kAk4JNwNGvZ4scEb643x7BO6h/gR
Xl41+Z51VAS2FOXx0Z32yEF5lR4K9qY+/h0yeSd9MxM9DmaRGHehnWx87UflDmOb
hjo6xTiwqamXEK2Q/XBK409/toD9tQgr4+7yqxFlBGqlckk1bUBUuiQYL6L500VG
flaZRJtlWFMHFOwIWDJwNsvz7IaInH3yMiqfVmFweMp+JMq/xzWjvUY4pybd3Vr1
ppzl9gHj06PkoYKkzS+jp237006fNuY1jfdxZmOvCBKbBCLG0MeIYnUtCLcMe4fT
Y5tTbKCK7qgisIsVr1NMuEhvwfjCXiSkilCEMVuUCEUneMhxfSQUET/uHcRMxgL8
UdfYaDOKHvVvbXOuudRFRrhgKlKnBJndFbvGGyA02ThsT7N9iV/iYGz+y59+v951
SbgS/iatmy0rf0hPEtHM/mnM5zXjnpmGjQEdJkCK0W8NHomyozAWC57lwtnf9pbd
BXnEHgu5hP2HMejK3OftrVGUFfmEAuWGOMLM45DheG1LyAkKbyRsXpXQHLn13RCf
i0seNDOXaE+S9I5TvjqrvqHfK4XFWlrP9cLN4HCgY7ftSEnfnu1zJHwLAjUnrTU1
oMdAAwQYbHJjUQMdI3AyrotyIQAxL7YfEuLcUieiG8tXM1pRWJA/qGqreXeHLY/f
v+v+mvrzCrEXyVTNOxqyol+iHxI+D05GeF2iIYsOU1w9mnVvXF0XdjCK/gf5+UrQ
lZxgooadvR9qRgp6IstLhpXJmhmpuTH099je8s/wxrd0xRHNdWQ60tfvOihCDoJD
7qdOkoTveH2nRKghko5yAJq/J4WQQ6BbpzbK3pJYV1oa1sNXUa3fcgCmYg9kOu/q
gr9I+pIxtG6ZIGaSV/t8mFwT2F5C1uyy+r6ve+1oxCeqOXwgUvtb8CR2JnoVhF9F
kYqXn5SySwsAdcAeKpuwoYP0DtCHcGckJhamhJljbEpQhNluaa9ADn8nZlTtQbE6
PG2BY/NSCuouXDvT58zZCVCX7uoDu4nUHyLWgqw2i7Hn2JSpdr1BADvabMIEpc8U
3tBeyg4J8GSSNj7bW6ZRTUkBMLkkdLmDhu+vmyYDFK5WsxPqpNGHMjbJF/kN8w1a
DRir/6H7kmt0FLVxPdfb9KI7axYTwek5RWAXg466TdSTSJdKJs9cpz5x0zOBn8FW
UEXsGRaSsE9jo6qQFhXldJAmN53tcOZz+HBFovZvhnjLjDqbBXY+cy8Z2fpX4AL5
2YExtqv6Kh5dBBBAiLzWWjgXSwPMTWneprOva46JF3dpTEqcgRO6N3W6jnRhR7tr
/g6rib+hu63CKxlHUZFT/1zJ/3HUq8eMEKE+oLgBNUmJY51IHDx0svARc6Yy7N5V
DypdZI7SNjXYCiw84oJJr2GLaaHdYc74I8WTluWq6R2RKhkO97d5F0+V1PVmzfco
0TJQcDcsUvgGoomdvNg/Q5hWYRcl8ZQnShEznb0D2QhFlmraj2UCCPH28Oi907m1
7iap5QcmqDEiAmFkQiC/GsQ7nkcpc60Xda/EZ5t079NOVqbWr7TwUJrR/Wea4BVK
l+NlYT8pKonzre8WOMYFRCrO931IWpUmlFaWGGU4wRTbKeZu5FLOB9MKaJqg7OEf
qQyEhC4FO2js6L+gwrXjMkb6liMTzIAWvuZ6RrdljBoKhqMVNiHoUk/eUP1HIrIE
QnZAC4fJQs35DUwQJvFlshDQOK9pCs4YI4SEs1+jqfk8Auc26DoGn9Ss1rCudlvJ
ypsjL/4TBZJiDJaLoY9sIFoLjQ+TQNPNC9rbAxbcKy74nbPK40u64l+Fga7Fqfc/
4jxV3Peq7yTtdASBZLCkNXIF9+U4tFfnC5Tigu8Eoz8LU0hlv8pQ++6iYyQsF6eS
Yas08Hd5LR4p8lRo9PKv6hLkCmjhW0n20w8NafmWWndsUDcIJoUUgUhskDvP9VKz
tdLaEGN/SPvWFVp8JnXYEyl1nd6F4anPpU366weGePYoyfwVLKNBohai7wOfbxVs
KtQ4ADvG9I+WKCtcLKd6Z0vpDYU9Y+OQdf+XMXsus2iROsIBR437y4UyGgdo5YGp
pWHIy3OY08dNLg5XgLYTLC/ayvRrk2FM18lJIlkwQ7Ts4H1vU5MDdcSF+ZQKbwCy
mf7q8JPfGoqnMPFbl+zYtvjCWpSkVYBD4fhS6BEvy+LYr66lGzYK+wbXn1Lk/7sO
DNrqikQ2YbTwlSHYxEkrfYKZ6oywKPx30Nk/BockrrxEwgCVZ/ulB+FtJxCjr4pW
OubSvLeH/APP04iIk8LvDpIdzjzeGPz9+viq2gdQyRuNvd6jhxZMmJiY70yw58Bl
vFHIAppQ3DEYV8IKw7AbRedvuqaLXWVG4RR0CPuX9s8s8FQVJ7/ax1aJbc4mSmGT
39wUaMWtzGESTPohVBp/jdNq95BQ2eoUglMxKeGPCtcMQiQYxRISePmKy/uhwXIy
6N8saZNmy8sjYW+/mG4cN5jyJ7ATMK/aJdTBcJWJy2vd641eM5Q/U9FHKtw74zNb
6vxHtXp1582aE/BZm6wkQaPhKNANmczH7Padq8yuWMvPmyTkfbAavfYSGN3rppm8
WPFhjnmx0APtSJbYqqmvO7VJ+DEMQR/2hoyEFy/U53Lg2PtwPO3pzjZJISfQV+5R
N2sBh8+Du4kSH3hIDSU6Pkk9u+b9Jm0Q9wt0bDc0AuUWbC1h7Q8WFxXJHGMf4hcY
YKls0cW5mpZKqxk5/iZo5cSR7cCCTA4oPlpCVOVVlK3zDwtgTGuyKrYCSp1BjceZ
ACEbyExXZveFXoEeMObH3n20ZpvM5g5nFDNu1aMUP7CA9HvGa+0PcyO5bVWQJq6F
pbzyy+V0jSAy+CgV6arrRW7gMWv8Twka00ftZnNn5or7GjoN8UysvhcccG0zq2sI
hPBejBN9+2PmQ0HGBWn87y1MWebC13f8RKmYQZihwFsb72voKkgW5mwYgYm+nCyt
4wYdF/9NuhdjmASCMK10sR+fynH7b430I0tb4jyIx5zNNT24lOHLcs+c/5kVkv4B
e089zHyVE0sjhFhcCCEgfaN2REgnH9aKggowvBuLC9bPk34qdahMsaz7jKedcRTJ
OeCH7yMF0Z1jd1lk5yJ+92n8D1+ELvGa4yu2ashnyUtBmN2xj7bUu5alobe9mBIO
ZvWqv6QJ6AHntGO7T3i77uB5IEjG5dkVyzNqQOn8jlJhWNe5dHpLshn/C5dlQAFM
2ry0LaoHEHSnwn/ARIeojMB5w0W+87TZbjJKJim/izbHCxMOBR9mD7TrBjL+Qja/
SAE1PB5vLJUiZFfUydoPK6UUhJJT8ExglyCuZRwUKOkI57I1Xs6KkYedUJi8aD69
9potTIemd085xbB3ZRL8rnAX0DHAVQ3ovdw+MuRlL/khxuhz0Yw7jjA/mR9ljtfj
TsyM0AtdHjk0tNOdnnxhTtgDMyvb2AEzVgWSXNEsNhxf3kfloecXA5VD8QCvHoun
QrsBaLNRq/6XlpU9JblpP98hRX1Qa8Crk639lc1OGrzKHOAjfOzuLBME5O1i9Aa1
JquJJS5ogiXgA1ibRvDNvsx1fPblhK1Z6A2Rz1Pt20H2/TzxDGhqcBGDu1RHo4Sh
c2hoC0wLI0t+bUPG/vNB67QwfoqFErqv45cI6wWijgrtFt+Io/tzB5HOdgsubnCV
OKPUP5zLb06u6t97NjSlUVx/hhNteS+6aQU4dXnsTgKvD+YeFVe1P+v/NoN482jw
k40S5YmswrJRH2qgQPAAIBB6Q8PebgkSosC/5Ep3jqj9eZyI+RpR4s14WRzTn2V7
eOgLiwiy4XgsJOcwRoLctRBJdi8wQfVYiOpSb6GbCo52gfVdJACm1ldRCyoCmYpG
J0Rhvr2sbnDnemrNVxElZFDrKCZ+/bUiMYpX/xf/IJtwDz3/5Y9cBt8nZOnvGwgH
TC1oR893JIHahBgK3SP5M2FYrznoVbmLY1FENzW9sVaddAh2IofIpmNhumzp4B/Y
kJ8ADblvvIlU3lMlb8lbRXmBZWP2ArEt9wW6neMdhHxDcU62gEQjBpnOntOFvRm2
tpaxujVhP8TTzs6YL+my81Q6G7kTsznZcF8Ev91u5Tuc7RLbCw/FKW5GvJzhsvkY
gnWhOgUEPFxOCXno/Tbym11Zp1FPrZ/zJkUmtjITzX6q/1gnjl1HdbW8CSL+JRJy
2+k9v7B+F4fT7z55WNAWTYosiAmSIVvffRD2LVuRjoxxWBH1+pfYpoYeopEmHeLr
/bfCFXkiJkiLVLBS0FMLWqIdn2DroOePUYSa1Xs//tmr2Pf4sgr8CaK00KtCGqca
Y3htv9HaF9OC5uG1gp1Z73x2lrAs54gAyxe/xhRRzporjefPXB8t2RicgzuAbzZX
OR6PRVYucVyMELP8jEutQuB76vihkkvUcLdzwIymoZU0q6COwePUK6jKOXSFauJF
qyogLLMGVzdIzPzmGFQguk1XrDD0+Mc38BfDVSUx5OTW4CEpc4mZRJcMYoGxU237
AjO64iCj1MyCBnFyOHZzRuBVnZQFdKJirv6wXuB7TGiqq6sIpNYYXNd7sAqx31rK
kg+w3fgYBN60XSiskyZmSsTavvSKFEJV6PpPasf6uQhPwBy37aFDB5woGVUw1bVr
7z/RicA4+P3gh7U4oMcnFpTbmpU7HAXBdqcNH8+mmzlSrWsdM5pt5YLAFPuJy/VE
Vv0s6lrilm/fw+N0u7iqc9KtO0M2aKZI3c/MitodrF0r/jU0Nl6tnG249ogZQuAj
/X0fZSSWOKZfGsdZwgO59pPubEcTtfZXoGZO1bYufhcBoT4baGE9Slp+GelNa+IW
mNiaVQ/DvH3QTbzLYOrRnPaNvQ6M4oS2W2Npf2kZD4sfqDqrQHO7WfjL9xcaEXIz
ycr9+uV0BRiabmMAexu8j7vDg3pVwF8U7AM3PQfMW4f1WE9kCDrJC7YRfaXyj+iG
M2Tz+7qs0INHV9R5jrxVVjjbAWo/c5cQVigmb44dmrOx4i0Jnl4Xp/YXDlQF6ymu
rkXKMh1lWrvswHleHmeBPdMuBnSABDq7SOk18rpX7eO3pEHvCudsFqT4TxX0KPCZ
ujf/oUWHcRRSbIiElH9H84XkySZlFarmPI/hG0uCgphbrHUeWQ/sCCICeiVMsE75
NtkJqrGE5XxFs16uQBKGu75wbaj+Stlyz1wF/6Pi4R2lf5OyG7j8B/nsL6CAxjFX
miMxftlwaSdXr3TKUsBRpuMyk01RoY/G1T4EeiXxjFEeBfZilRRh/U9upMECRLsB
nf88+M/Q5Kb9QElb4Lg1zQuxpq7jDzVfz0bi8ubTSfCilVGNG6MW/ZiS6AyYkRgs
rSw5eGQqZDkFusMuG6NO0JgSwKfI6z5jZhWK5N1TN3qXabI0ORrLDTnrfoN+d9UH
J2U2hQqBthNmogEuQCh3PhQsS0hBUirA6jD/mSGtFX2uv0rEbMppGZc4atQ3jWXi
l/KO8ZocKELBD8OYP4cDmFVmWrz4SoC8HqEk/RtsJTcDaJDrP0CsLs+Y1fAK6F3o
xnR1LVlgfl0ZfobzWg2wdJ8hukWkQ7U8X7XpnjNHlbpLA8kM1Egy3dsqL7hkDV5/
DWBdsb7I6kUvmknIyGmipPgQtF2ARVOCjc0bsQLtB+XCeb4sVjVztNElsrhFazRq
Lv5Vdk8ycUbahlWrd9+hTP7sK2ok/UpZiImV1eutU9TlIwPwIPk6N4dxIGs4UhbS
4r7SU4AExm9HUIoMGQeFWsQj5a6K1GZW/8b6ZJJBbHIlVgecebdJDO41RBOkuihD
M2adfCTMUDLh+tGxAm9sB19+Tln9n6vHW+Dzhn3qE3DB9lnaQAzvgpaEt2iwJAtR
LkeoyOGHPi7UQGd9voxbU1JcloGgwZUEhkfWP8SsGmDyV88GQBBzZfRbAOCSsZK1
zpvz9+Yy9GAwc1b/alFUz3SdTBtqK1gkr92VWrHxB5SpNDFZ7WK4c6vCpEuzvOe7
Y7J8JjdvWVGvqGD3aHx4hH0cJJgyctcFL6dXBwFu0IYbzyFQn248IMPdzQf/9fGq
4TlXDhbZoRxnfA6T9iwsRyOXHNUYRy3y8aKw/NvcpI6V0K0gy4CJmoezPKbuqUL2
Wc8vaKV8SUL3zp8c0U9UQHmaRzYwwCYUlhRvKnHMeHruCxN/H1CWisYjZG2jn0cB
EnZBm1GPPBG+DYsPemisV1IZJZmW+NTXzGzCSnvnhm9wLep8K/7MfVXH/p79RB7Z
Mf3im0Ip6Nhj+FJ/GWxCPnSQiG/PdlBZBtJOOBSu7mM/tfq0/u7MgHg7EKwGyZCZ
kKnv5+BLT2lgfQD+rP4GMZCXN1U2e4T1VZ1xEe16wwsR7EBgx90eGFPHZr26/Wm8
075nrOd3myHTTvPbgTdVjzMx1PkMKCoYUtLX/9bv/BUir/1J+UbssJ6EScl+u7Lv
/DxVUhHKIq096fyPaafv7xlyBntb/QvPeec9bnIoefJqjtkAbJYG5/s+7z2c/MsG
G1eLjPv8CGkZPCH3HcnRGkBNEx9QN3CgC5Tit18tTIDTxop+yeldQevjBz6HBEwn
rfP1uw1U2quaQ1qmVnggzlg2HkCliGZHcU1TgOGTHPVs917ePFRN/oHIDRcOthh/
a7iEO7iOxFEBU6owaTl5ACJK4hAtjy0OpoGcNUKQ1W63LN3TZmBQl7dOdi7sKxQc
u/EYehArC6hahRG0rl6yg4Gc4FLfql1nTnFZVTassoDKT+53cUplDdzUnG78dHbB
ZjTHykdBHGDAd3Id99uyCPXJ05aYCvnjstCEU6Nvq4057tQhqqp+g5IF7mSR5706
cao7hszSf+Xuzr9uuXpVj8zShzL/PYr87FEoXk0ccLRa+pc9st2t+98Ku1TCSXwM
LYMlWFK/Zjxb6vZdW1TQURVHe/CVGnlVAhopyLrE3EMr+jWR84VEAEpIhXN2J5Ko
XVMMkLnavE3xIrGfvMUPZtEvYM2jgxYK5X5Tw2QfOk8CwB/WkscnoeIWH/CyzJU+
BTBjDI1Kzy8oTQqA5cTRlLvo2Zocy8KBXTt5nGg+MbxGMngyTc65yn5qnkSk7pG4
2UC2coZLLQvOH8eBKJzzkIQotQ9AD4L4PAymiFi9cIlD9pfYeT20zwTYlCwxGcIH
oJdCd2XrLC5BPlBbBxReAglkmvOzSh7xsriH3MErNFGiZkKbFSmI/c0J4MyeYZUQ
QtuvD1uEfaCrJ0DR+j73oNn2dJIs5twtvckdNzfNfJEJJ9Duwm64GnlMqkD3whvS
YbOgEDOzXJepQEHWs9dIIXskMNWN6xWOesrFft9qR2NOaun+Wgsls2h2Z/LrwgUC
WwR97lhPbJHHkY93+Wv+aPG1Z7Bu/khZ3XcMzABWqPc6hC1bmLRI3iyNNxOnFKUO
IJO66mphi5OaD2zyVTwz2K1IM6Ymf/XBgi4mKtyaycN6jAeDDVEmySdx8LiHfMPe
sQYNO99LPvytEJQuTE0fYWSyIH9hIBMeb/RHQpRet5VLjwc62/+W70+s6qwg2DEX
Tx9UfF0L0o5g/6hOdxpAtfpAAJz71kM1YbMAmm8N8MNfRfBQ+s2LdkaYnw6A9n9E
ONMdhkEFqhUn0ND47ozLHdRi6qUwaLb28FsaOeQ/i/xRHDa/IjzCPN0yC/RApSwM
aPrEMLPbIVGubXxGN+kpX1ebIJ2mExD3BIrpPr0pfidJSa9P0TJeAxBRTIvLf9q0
US4kj9ItHLYlwMrhe1HAFd9uTS0hHBSKqYvdruxqFBn03FzkVIkoVenS30FhTJ3r
x92LiKaN5jAs6y7bS7slvSPYIEjqjNis1EyOs/SHFv1HDsRy5uslToE8r0+f+yWi
r1LCooBr2Rh31NnZWFKkPc0x+Okp3oi8G1aIDgiNwh6S96yuhHxkPXlVGmrxOUJv
Nd+2XzeDMGh3fOkjNRYWAoTPX+MJBnQsg4RS0/RXv/s1ISnvVxOwQpjSgjZKdUbG
CKAVUV3oiSvLC//Gs0zc6bzYwFllD129XEJP50dHWzxiuTPF4UJJMWaq1iA72gtm
FLbK5suwRorjRwMZdoGWTc6oH0nlWlPUg4rx+Vda/zUHK9fKD2N400tVs6HpduAF
IeydVMzHnhUx0IFVTASpU05/Bst3kY6AWOtyA7IcePIcbuVlLunkd2R9upPYlqW9
ccaPElSaFOyQglRYpDAq/luQKjNjVvSlbLiMVXFM5+PUQG8CLg+c1pqBbR1aG2fg
4dmXE3ysJM6XP3oMJQfkzQKcBgSjvWDWkDH4DyTlHlFjb2InjRInX7Xe0cOrpx4W
24GXUI1MilETMMtJZVLjB35DjnayQLZkivOvkEQ4xUf81i8WU9ViQfla9e1RBYq5
6HvRPmU3QRjY2j/5ElCGRkONWX+FajhwzGBg6bNSr4kh8oU3p7u3FtT6zla3hvyJ
ZniUVgDe2V7fpcpct8IFXgBNnrqpA2oUf2SWjPzcPWwoCvEGg3orKFLEDr/lNWXe
lxZKRDbUAt3G1EQZ3GHJHB106mY8OyaDYVKEamj1JW8wrF9Tms6nRoX5l7ARL0ry
I+zHdfLzE1zF2dRSFKZZd2jzfYcMnI520namYyxZZPVMCRFPByvqqIPzi0/8OD2I
1osghEGMvLbOBMRR2yspWwHfrV2+01w8GuPXr5Qx5ivUG5FQhgn3BL0GIwt1lCSZ
HS/bQxhKHfJyIp0hFYiaUUGl6Rkarp2gCyHiVmaytfT/yRYpsx0A2BeKllR5/6+K
5KXJCH5vVkfp4KBjIqRLyt/TjCsoz0lED0KJX4B8e9ElMoAHq1ECPvzgiK1XuGRA
lpKqnopQkmJeXYvlKhp8Ol/uluh/pjvSXUENaZdzUEWMw9KItPyfyzEmN9sJp7gl
PJx1FzlJwHNBAVWa4EOJFkp2BWDAmFd3RkOsnJz9pW+CA058LClp35l7xotrSj9l
RUGc4Vt6AI9XRTwg95FuU6qxTn/34pNV1HAFM2UjozOhLCMUcSMLqE9HLuysqPK8
Dg/SoUl46RR52bV1il8sUa2Fy/UCAupyhG5LK6F9RfpoCULOoEN8+5YowpJhk0Hz
7fEZuCJXD9Yw+71q9cefLcnxOptgzAnq0pYjjyKP/SRVI6iAdHoxOyd1e2fup8Zv
BIS4YzrjzWgtvZjAGyzq2hKIjZWjb8HADNOIUI9DgIBSWLz8W95NmpT6GOQBmeI/
HDClbJYDLIMBH9HB19zXk223ezckIR8S9hD4u3K1qNMO8qifRJZmetu24Qhr4Wtd
E2WOJTfjnIp/7Jz8Jhu+5aRdu/kv2JyUh4JCGGhxw2RMK8fClQggqS2xsibzu+4Z
djcTna95huawHHx8oL/D3GZ7FzYqY7G6NwxrRU32UvkcPzqoPfGub2c6Ohs2d5OC
jOBqi6Yy3FcIYjVm4hN0xqMZUaG0JblFpQNvODQogwWmA3MuAO9sREi3jwjKf63i
3OFpvh34K8GczSW94kl4E/Rmzip7CmoLE15aI4Y7pmey0SYncXoHjIP7usmo+tUv
EzLg5ip89Nfl85RZ/xo24W/zIJd8agDJ/GIi5UB2zFrldt2Zf/encvikCc0J/C6e
aeRhh435K3Bk9kWrml+0RPNGTZHAN1b0r0Z/Jo12/NrrNpry1KifCYlSWxBoyOGI
x8W6oVbmbjOJj505HWgQoW6i4wqTD8ydWepc9+Vs9Mg1Fmf3IvpNkZIwUgHKy6Wb
1vvDp63qYNlv8Ezaei77v26IqPBsbOyA+GaHsQbFuCDiRai1eZEpfMG4NIzs+nuI
JHGQ06it9TjFXGRBwoQLyEHKGyxqjOJtbERk7McI6X6iNUdZGK4niehGg6zb/sqF
pU37dmazYUVQoYp/UFcQDR/KCiZFMZaavuX7fVwlPCtPagR/c2wkk+ONXNLTXOYP
B7LNxh/y/uzhZlBYy/x2DSRVvEacL+9D6xflHN72g5vUCWlU+oprOpOWknaXlU5E
/r+sPGR7Zq6RStB0gfbBw1hIDIDSlpuORW93j0raLMExnRz1JHVzE+OWdMU+Dzp5
fjn5ytyrOeTH2lrTv6Vky9hTIWNasVg/WaLDDaurIZjeyRy0sbtXgP96X20N8ybQ
2vsTXdFYzigecM/j8a8rUoe2dlCq38sG3JIHOM/cGa4QryKHOEwVdWA8uCPldlWr
Wu0sRu7u9fM+LVDf145Pm753GsIgVhT54ZDNUlfs0Tu+9BnFVdY2NxKs9IxqLFtH
/P1dCZd6jz/2TYK6qEwBcHBES4qm+g4Na40zw+qF9iSOG0vn3CDOmxpPtWLwPf21
Lj6hcwTqQO4EWTchs0kMwf4lFGUOGqcRvYGLPiWxFaOExuyhCaZJWHSYcIOW6G7c
jsUmjt5el1BH1sdIa5q6bNduBNByjtZJcWH/L4nvmxACBxZgh+/x3IXe5ZwOXsF3
3k0BVZ3asdMUw5+7S8NlWZUMiybH4ontWp+xfrIIBYC7bFf9vBGCrbpTSglYlolA
u4Gh8XWbOUlqBQkEjb1I4wPBfOGwfaDIc/vhxraARhL34j8Dnq2RLGWGHuj/ZWE1
m5q2LsjCua3IK7ziy7/gLGhH1ewrujRTAhs3KFJo9fj2m+/BPFygeja540vV6bLZ
UZIOGT4qMGWkzCgfePy+qcbzSdVXTTBJ34ngmIzD4cCuvhgGhM/4o+7xnA06/OS1
bdY7EtmXafGRp+4C6RNCtCKUFiVvUYSCgsrfQ9DYRg6yBTwhkF46ZmMYUN6eyFB/
sIsJB1oMIOIhT84PR7qY+GCqrTXNo8o3iCf06WboquSefEEwYoKHTXhzktlIFj3M
4cSSB9lEDftL1M5pzX310uEmh+yvAwcwLg72rqCJRQ6IJhA6YvN2zyIx1mH3cV3H
H5uy7d2Qa/M5ydhNm5V4Z09GcTSmRoxoHFoBExAh/+wj5KN8ATT3t24onco0HGnc
8gc77a5OKPvXvMVBMUP+ZvzN8gC1pe9n22jIPkJT9eBM5HjPq0vE25uTJ9hwkOdd
9tAJn4t+cn6AD574V98srU7f0Pj7Td8LKwBtEaUoSyI0B9bYIZKpZn1aDS9OLW+e
QDMRbIDu9uMQnq80bIF54/U3rcD0PL6fRewlNOKudlxVTIyNj0XRVLMrFuX/llGJ
mIm5TZ8S19wmwrJv94aStZuRosky0hHMQXg2vE8yRT6XQmmeCJwjw0R+SdlNyN1/
h2v5TGdXZgw7ky/zo8Q/PdNIl6g6ltwVZoRo66BYA+faO5bEYV+MgeJA2QanXivg
vZ2hwtGJP1Fm2dgGruzs0frxTlQmuj202UqLKCMrcV5/JJRakb1WU4N8hwbV15II
jyrtTWsLLaOl8jREC0AsbFjp1fu+ktidv4TMjM29vvUkJE9kgUzyNUHxUM5Jpbdg
T8GO6ruXWADpOTa8/QKCefcnvqrgVtgJY+rbqyniRgLWACgdZVYduRbRkTSCLHiN
X6wXthMKzIEKTaQ4AggQU9jt2lTJ+KoH97OKXPo+9+2rl8xK2aq3hc5Bip3ieqgE
Msywcecat78h4f72yMQJImFLbP5WSzIzLqk3EFBCNYHph8HgJ3f7Nf+3j9KUzCiH
tuO0h1f2+5QJfQcbeaukNm/rjVprJ6nEg9Y8g70VOmtHimCYTiD0whkN/UYB7KCn
EfyjcfvfiYW6dKMX3YPWCP8d7r2e/wmMoalRYBtKZd7kaRYFO9CJjcqCt4O9313f
M/dGCs9wUXjPy4SKSkIrdjBIHoevD631C12zkyuqF7WZSYCZEY0XznZodazWRUYI
k3hL3sJfgvbRKWD21el9kvor/7hBdDy3+tFuSuStTqrx9qRGFWZauXvZlPAn3Kyt
N1NKOyVkF8rsRPPASjHLSUqkESaQdwhmEcIjwJb7DCNauLTCfsAJl2vN/EoVZmUW
kabMWfXO5k4DQnNa8SY0sRWOVqTF/ZOFpx2Wt9e4J1CeFuuEk4SFkaAqKZ3pjX08
eNLslyjLIABnoQ7vLWCvVHMoXksbPf0OLKLMpPt2UBNjyHlcopEr+M+K8OsNKX46
IHT6VowQwFtmYRxq+IDtTdz7wNBsV4nPorNXuWYlFsVwgK98GW/U29yMgKF+gcwY
2TxRqVt0GASPpLNHEzMqjmvC/eq7Et97ejHhuWq9hbVk3PZ+cx3iwO/3TNiKQAUH
x8fOe2mvOEAjRt/HlHeHldKn4R8vdsllP1D/cBmv4ENlNCLODwsiMf5jF8RE+5n6
Wjh7aAcvAJzmER/RfU0QmN3k70QizLl8Y+N6CV1q5FB+QZ4q36vBpK1XZgj0iUCE
zL7tLMxGYBfAygDaUBFj+dEwtw5tui/KOELSpxsnqIjVFD9gblCTmJVhT6ajMF+p
2cYjXI7tpwnSYvzzo5FXbjKInf1HV+sMmyOaBb3W6ppMacCMlrO4kG8WCsEXq3y9
2v0AXxWhzps5v4g71oApdT3C85obp+aRrv77cxZEP7McBuSCWtARruYdatO1rfm+
VbnyRCFoDz3UyJxyCVT7KqGTjCoQEvokH8mV45ehfePRyQpGUlweEtyz1Boe00Gb
yCNILTPGqpsk3g0NyaL1YPun1YVR7R42DmAprp8ZcPgcuH4NJndzK1hFC82BmJO+
OeJZJSku1Gz7Ku1bVv0U/+fMe84oi6sL8RPUsRgZjR5zVJLVoMukY3CS3ZSOeB5r
bp9iV9rg6RN6usllA0Z25jcKR+XdkxZHXF7vnKKvnlJID6Y6Pr6l5GHM/0P7Ce1Y
rEEm69wsLi1maRGxaFTnN8x5HEKH5dF3NIQWGPj3a0HiN7z7ldbQ304fEQL9rngl
tXds/Fa+xwjtkytDpH6ZAfV0gj9iD+GmRlf4Aeu+LQvdHTVaaeebQmH4fMUPRG3L
BL3lbAdUVqPRc5euIqgNmJXd0V0ahpjzbn0awxNYvbW4F0nKwoCueSgmQrqS3Po1
dWJ2cDz3GXXg7x6kPtgR4zxaa48CQvqVimC/LSxPXwALnfKO2PZucZA8oPzCstsT
Mjt9X6BSXxi3lzXSQ+KfV+BFISaFSRrnFb+vB6JLFevKHWRlIb+GmGICTSPvGuZ1
WRyAcMr9iIDgF2z7171MqBVCkcVkSa7u+E2iDnz3LNHqdXsq5X9ekfYu1e9u+clp
4hxsR6vy9Dlxx3JonUqTDXUb53XGb7/rWuXzspgCAXeTvsYJYJIN2maAzoZLzrvE
NVpK1d7Fd//0J8TdS+mvVuzP1LazlKfL5v1WDYvqbsNoqUHHBGdk24ZI8k6xnUoP
MnpkXmACCK8YkzdXklE5VHH7RbhezDv1DIKd4Rs0ZX/vzN9f+FMHVxja92WvHjNp
mupg2i1cRGGeCtxaLI/cdCaQdug90LYvl8ONB+/D4byhLajBQLgWmC+m83xGqwvK
0mmV0FOJqCFBg0B7vIqkcEbVPqFrzQGssN351JcwE6gSpq77GAqq3nY0GZHevMAQ
m5HWjoGsKVakRqirSt960OPB8jXu0oDkp/B6Fwrt3mO/ksbUsPkDxlYiadQ8jAYc
r4MMEuL81NjyPGmPevU3tReHATsfFgqL+wLG1Jw7KSITfE90vHjlTmLxVAWBVEHP
fHQW6ly615OtHCJVSIp4BZXib5LsY+I00izMdUwwSFidCZNb0valuv1F6wWaJMkn
f/Vuqj0zOl6gfUl+s2fv6NZg8oJVU4f+XJJzIIWVAeyMsNZZ+A4gQU+BmiDXSzE7
fOILQxdCYwOXhGeGSWE0y/5+Do2ZivildOQryTAMc6BkMJFrFWY9JWo5EF5gbeZy
BHo2RmZw+WYCYA47MgsdMDUdhkTci5z/GA7gXJTAV6fjLlqNZcfQOq2ZMeMTr5a8
vPDjpKvau2n4p0lHaKto/zFLZBCR5yR6bMDUMfmWJJFOdsmamin22qVf9wde7i4M
BARhE5akI+4S1o135KkPhIRoypOroJ+cSWHrdhnR600gSoe641i/We2CH8qaaVgM
GM3N7aKCVd3/13zLs6WvOs44rM4AhKteZlix12K44DFk/Kc5UuVQLGaqslt7fP97
e/ZlVY7Q+vlXm8Rf45szFZjr30OoJ22AWqq+wr/JJLza2P/bBncaC17XF9uy7Boz
0wsEWrvlJ++3K/+aydVBUkh9I/sGaA4JQ9VYdLu8i7zki2i70IhWVFh236BL2L2h
DrTA5uTn+mF1jKNtdmgsd8gzGf5YrYEOKlIVoWJDRYC43fgtiAae0L+k3kb8J3he
cE0fNamrAtCqfcknx93Dz5jQDlayq15uPztxcwmgvyIuhVZBYrMuSQ5KgplnwEme
2uPUVLCiQXsYPic/LeM+0BFvtxwLGY7g2xyedOmpQP8hmBOA1Nl71+miErf04uIP
YJI6bp6FBVVGFUCCNimyAdPwmOE9nlVpE78rVv+0wZkwSmkrX7os/VNPCoUKAm3B
W7qvFWFnO0P0XWQdhjSA8EciVsVO6pA9mngii4BlNVQ96+Xu+TKT+YCoHHGC05+p
3v/hg/DIvSuCa6686VX7lBozqvA32cetXZGFsj8ns9g02UgpSWW1HEHjvBqIlW/p
okK1x4kcdK40mowiRjzXgeDpFRo+xUZjSvMXg/AJff25Bk2r5ia9XT3asXwC8O7z
zsbNRrGNxm/Nqhbp73HP9C43VM+uzRl1oFYIh4Y0xzRRoFyUxbIxsWeIVAadkDzF
y+UHkqgTzwCEk4/KoMF966q+6sqdQrPEE1o3smVo35qY73u2BT09MOmaTtsrAWmX
5PLok4+5A9FO4Ab5fALfrz7m4Exjve5ApLZyiAUUvLcE2WPS6lq167uaxcCl6cUF
Ki9cqiFdbORRr9e1kPpg9GqNNVMjw5Y2GpioFQiEiw/qClwvWA4NcA/H5uZ9NVrw
lsS00hFwJcRmpG9v9XSkapDr0OHEsss752GVuycofK1EzBEE2+6liaKkNms1Rl5W
Evg/V5pi0HQpSln9oIRhRARy5ciBK0TT2eyZr4QaHA6FdI76DE91ebZFBfuDhX8y
fL9rUcqEcKC2rC4VIrBtiKOcjQLFc4SmYcOkNeyjPLbz4afFq6XDcXmfzDbe+lKW
j+iSP0NT3kMJZiAddVrrr4IT5LusVYGtZnru1lEF0Ibxg3ol06iVG9nxGhGn94g3
cMZTpHrwIFlmXX5QVuzChYTzeMKScbRshoGRtGxN6L6NFErRW85hMlY1H+I/GgQC
GPUrehx+8yOwNEIrkAeS5GCZgniA8D3Dxs/rdQSaex/ovU5aAuus5J0wbhjO/WPn
c61oF4UlB9MSZJKaz4KjXgySdTZWpRtpmHaCnqdxw7jnbcjDAyAa92rJMkbrli/T
dL5QUynBCIhOvPtlyciEaeR9n7uVf00iWrSKzELLrwqT5Ig86V4ZAMZi5Hv1eEBG
MeBPi02eQWwuCsvKOUvNGwfbO+h25bPzQEN/Q00YbXXD5jWOGgyg0N9kkThdXr81
D9vLiz/Yc4v1aRRLYajXc86+3EEOA0TxCksiwQ3E7O4SVzf0xrrKhcT9nafPluHC
2ujNf+QxsVCX/A27Ikp5/wSksQuoJSunpmf0JRdgV0fWHsIXTwB3tlqlMQAWOYUf
CHsD8KAQwBRwEPfj0FX3UQTH6tYAvE43dXomVlEYWHflOO+YASRQ/sCIsixr8c4h
mf+vEmfEpQ9JvHme3QM48vqMRr9zGx9TkpLcnJDBGdsK0pCLMJhHICfl8D7b5mCf
whgqrlO12KFYUxG0i1p731QyjMdb9w0fqAtjy70dgEmJDSpQpwILFjN+vl1Ztfve
AZgAp8AssrIyreGI47qCSOVPgJqEYShn5UztrKr55THMSGTUXSCzIpk4EGAp9IPL
w3JMoA8dkcK0pTggeBprA0AZ/1qdvxQ+OeVIbsCYTjzaDIwVIYvHKRp3PF1Is2Iq
3kyFQPhWhFyzuv/q0npFtcKg2OMuk7OhnvD3VOlMs2fQisCI6iluhn5K0OM+9lUd
uZVDYSONFzxxyHIqQuaKqGhsckkfctwi6Mf6Ow7Oia1MYwxZX0TAKTjGb3InuXyS
YbyTtZrgBo4cUPksnUHBhnjocWiNVGLl7LAJMGZC+9RVcMU6aqkhzHlOr6kQteAg
hSNvLV0kzo/xzOrDSS9RacQW21dLgOmozSRjSqGz8xlCEngXJNX2GyK9Upit3DE3
5iEmZ28lek9P41x3PgJBnwGedXytUNogodVM4m+1WTEKvsDEs7e/csj1P02lUsXz
BVVVfiMHFHq2SS/oOhdpdmV7RbY90d8AQo+2Aj2ov2Tc7D1tiSQdaET5ngiuA7Sn
0p0T6w0vu0eYOVPV4kdFCLty8uutWCg2I2ODTyrBIENWiiZKREAyv0MDzJ1qvrlx
ChjA/fEvMUlyAWyVP+XRd9UteyHYlFv+j9sdwaf9DZjLHe6gm6ZFs218O61uoryW
ck4Xfn0EikQ/V7U5PnwmcGjLSRIukxi49H+Bhe67S6x0bNx4rS8CMy3RJ/IAwYXL
czp4kiQAVfSkfWxQRMYJ4oBmxvyds+y89DpEjuNujBHK5SHEZqlqFKYsRoJOA7OT
OA7oDfAs2iNs3GLUhLbrcYoJQ9KgHo/yT8VULwR/WDqKB6kASNvts1bHihucmgOO
Pv3l+U55KKlrktJFa1DbZuvrGG26sTVoj4G1qie66G90NZJolJcjLFq5qiAsGugl
Vnc9GUw2SQAlNADCCmaUkTvVZjGQ/dNLMm21rHCV3LTqJW8z6u7yuKkCtaAjZ0Mh
E+oNwEYQNZhjADjlK6WPwxAGpT79VL0Otj859Ppnf6MSYMmEzF4gmGM/OqWw7FDm
6dsyvcmKxQTp08/uzqmYbxM1jvI3BmRbOWBNtnWO7MrTh/ZyC3q1SjeamgwKbAUZ
VKphwhC+1K3alJPkin3/BRNMIzPHl81+7qCBBpwxrcahPYQXlfPoj77KBPY1ey/9
LHMM75Sprlw35Gw1mFEExkArRXI/xohRC+s5upbaabVxA3MpyCCkcsrWFFAwmNqV
JrPwDkSWPHW9LeanAwC5ymXTU3/xNxz5Xk4AogUa8NKPEt8ZwVQjUSwY0Q2RcRze
CIzZrBsx3o4QRxpEJLXX3cGSm9dq+d/E2RFe7Taed0eRYNsj0yjpbxeSy63xsNPg
ATpVuTsE1SXy2F5rkSO/BpBy2DMTv+7YV1CFl/9yTLY3ccjJ6lgbgAAyhzUHkgHT
yiuZtHvMZ1I0uRdhfMMW1Q71hpLtTFhLhucUQI48EVKWBJL/1+dlSLzqSjMdANAD
eyELefaCV67CPnfUY45t/Nt7EiBnNUxu3y7oIMdOfIOChqpMxk2guw2Zoh0GBvHW
JrIWa7NPl1ZT0nvIeewwlfWJCEdOaqExt5KwPfGa1bFAxc1Ua7hyxQ3PbQZlDEXA
Tnc7sa2r4nTFZhWkZoCkhKqqBzDAdbIHJ0F7g4lICe5Lf5cSANzQ9HCVwKgnDXln
7CjXaWUmTMX9rHoKOOZH1M8lQBn7zdAghf8mDnV9lIKZI2gD88zzEbndFHAXynjN
TehBb6FE/2a+aqMQZgyS78bgEm6e+tEf4p1B136EUxp2B+ZjfGOgt+koHPXKhEDn
74VMzD1/nOTa80MxYDJpU1bHpfmUNzkqfl6IZZ/sZ8ymiE/siIHciAK+pBC8RiNH
wa+7v1Q8dUKlxjST51q65//eKcDNsNf/NkqNqxx43igWNPS1oxp49pYWH2tDXIWI
23P0jEMV4sBzajh9hu723r9bmD9zJrAr3WiOmi1vZ5er1XpiOHBEwX65T4WSCMwX
77rqdGuQo6pDOczzHC/pnAAbqD5pn4xROy+y8mUR0rFQ/4nedtIFbFgEazljX2y4
RhtWBPMQKBWBhT1Xc+oZKXnarrR0qe5bUZWEVJJ9GZca8G+otcP73yVC5m0evc59
4eEtl0fhA2wF9Vv/Wp/U6I0CTimoco4F829p2qzIyDMvA2hluO7c26++HHcWT949
JhiSHlGRvdurjJ4CX8E54xbVZyBqCxFXnlGJVIZYE6mtZ9jutLG1xl4DhKd6sRtx
wgmfu/r+/a0b40t0C710ia7ZCPzzg/Zo4gJyUWcVcvfGEYIs9Fgv1KoAyIlop3qv
1h+XBSU+oC1nwVRu4UYDlJqQZ3Qm22hqKnryKYxWhO5HQcDCCxIQeSSYSyp4WSST
1pz4hC5t57fwU39ufqDpxcvFJvz1STi0IHn5tmyPUjbdcIt0JWFEtHlsR2KS+W21
T01FVRRd2P00opv88LvjsCfn5vZS92S4ptaGz7Nu8HOafnzumCgAl/2Gm7msq57G
qY45UOFS46o8TrwOa/b+WsoY/Li1mnqcF9lMzgn6N9R8k2Qe2YkS8kH0dnbBfRap
MmsFGJN9xp4k6p3zk1EEZOlToW3CbcuXFqeRGFrXm2afJK/9nZ6B9i0ZehR67yD6
Ml6UvisiSRQlkhaXo9WL1y7vWGg7pSNzIZLDFCWTTictj6yIs+q4L5ZnBv/FA96d
W3CQPQwLXf1n6J+/vxq2jAKXdvBKKlbwco4Uxep3pGUN/8iqQ6ji7C7E4V0OkTC4
PvNkFKqjNmTgESI5BKuGag7bNHBglkigCYpfN0dKY1J76WV/bS9Vn6/bV4JO9Dqq
z07eB9kJBKuGHre+smix7t/jFMIcpAHhcUGnRNkzsZchwWzq6xNTD8m3Sk7e802t
rAhcJQ8q7sxqt4qDjlNHSu0NMox6Y16eTCij+odTtBQ9hE9sqDeIh0FDJf1uf2jl
OBoPkQqJkI6CXPw0zDHKiYr1irLSj7yJhM+RtkcGls1U4ryTLZJC7WiHAtevfDZz
r8sPgakOnmbfP384IDHuzf2j59xm1WOM6tUSZWLNcbHfj7vDUKdlFJnVgYoyg6qr
kvSeE1cJJ7E5VpoRWmaSeYySFp+z/WV+JXzhP4bnzfr8GjPgcgmcnxX/qpLB3E9R
8byjwCw3b6x4LN7h6Q5Rly1BARBlprRUkwKIqqPwCelsTJOz8Q8v3bNzk86hnQ1W
6omnWlvMVwfh/1g+l9Ry3KSL3PRdmeKl1ggZlCrqK4pKQjTDX2w2Fq+dDahQrBrL
Bv9bziZW7ZprgKz0SyYvT0o96aKJV47frq60wF2em3JGOu65Gf6hPXOXL0zyQr8I
FyYHpM62Ym4xD9mZWOjHhWBolWbQpxTcbS339hozUPmICvQ8F+JSOL+a9+BAL9d8
ezjQ6EgLlkToMswVGJsJeHkSMa6UA4gXs6w4vc4H3meqwYKJRNrvEaFZarTi+iXT
JC7dTjYBMAsrh67MlUoOFWgFPn6W/aMql7hAcw9lv9sZVQw5HSbIFxdQyfbPChkL
aiH2lGqkrAzsC+sxfiEQEVg1kTJk85KHh8deoJJPkSrGxA2vCVUlS+V4HSIQoI9J
6pbZIBGLr29k0iuD55KEoxOWtrecqve8N5SfN5RDD0/T1oNQC15+/PcEnDk51gXP
LP1Q+a1kXPuXNo5zucGYMiw1HJWs3nQqv5rUeoH/biYvszF5HPmPEFOHWdKaB9w6
taF97MG2sZhL8lHC4nYyw7wHgTz7kLG7bzRVG+LK7KngAc8P0RwJEnp/ZMJ7Sv97
Bc1k2r3M7qU/F7gSOEBs5w9uoReyUenXmoFndhjpBtxw00i5OeyukYH0Ysq8piop
0xjThN4b5w8WVHZDD1AnOVo7c+mONHJywOHBSvufyn1v/QORyfs2xy2gIpkoDE21
sMgFY7JEA46NLBG+hHZe41EEbu1Z+x4s8qGcNghPcVGL2QK6J01fkrl5W0y7GTC4
Ud38FVfrdvmhYnyv4Fugj60B2nKCRM/XI3U1mRxB5zB2uFHruZnlp0b7NiwM8cEq
Rlus6PqrCDEoZG9Y1akQt4FFomZrJO98HGIA22YMKo1HgjhHwfpucYKA0XcmQVNH
qc13CHxzxIkAg5v6AQtdVpXBquG/cQCb/vYJY+mYatiqVNU8oehjPXyGVmC2cx6c
zo3OR5qkbKsNavRDEhTpSQZ2/zYLAyPLanFt1zzoEs56YjLD5aNforsg6i6QfSdk
W387ueH/tdWGVAyYU4WQfA3oUUAkJLOf27Jd1TBg3vjfpTyjuxxyjiuwVLTtDuDK
UkfMJTDPudowhcZSMrmVTcCvz7Fq9JETVbuaPsZpsh5kHRBhs7UEIu4pDakWFwMb
EcCUXlkpgAv51EHNlrjJ1QKRmscLb37zZaFl5PFpmGgOhkbFTlBoCxam8Owt9n59
40+PWFgT1qdINQ1bKO5A8R6fBbGhoKEfDKoGlc6hNyawab6UPHJ2niCguxihFozC
mpIpqCYMXFjU6Ll1XtQsbxATcdj3f1BEoDMiDIvFn7Fi1SiLhhkvBg/Xop9AHJ6B
Y1JdCC5uVTXnObvFeXLWKp9TX7NQhhJHvJcoq/y+QY80ran9kLoIFfqiDvl9fNZV
c06bBGILXqGsM7u+43D9rttWa+HMvglzXdb9DUDntA7Ce415HPW9H7TBEy6uk/oR
iVb04s1PaJmQUCfzZJNRC9IDwLw+NHI4Cal47GBbIoB+QsuYSgPZ7wPPt8J6/271
hjwkUmBoovCszgCLzDyqSVFrZevLC/rZJy0K4oE3vMyduN1dANtJbZnKjxI0Wsu/
dcdV5jI4tksQnZce3EkRlW5TPxc5lIMX3ZcKcqoIobgtOsUXHNABMQ6lnZQUO1HD
q9j1UffAX7IPgIo1+XSzsHkqbEo4vZm3+WNbdl/FkphCt7GvEhRbLSTaC77sAHGG
qftkj42E52Bd+tcnoi/msFPWvS7IpbFwlxWtJe5SWx+ZOQ0si/oSvysCZGfOmFZ9
2BA4Sl6PK+5Ckj8j5a3Ueelft0SUT5JbQigeoRupNvPXeHXlq0bPlMFL8CZscIT9
BoQxCrtkxkEsk6XRmmByfAmEucxMjBT3tOacTfl1y2gNYk5UAkg+4hvpZusjQkBH
SvVpxz11Clqt48NlsolKlXpIYfw8+IFxTkoHo7kHT0287T2N841e09MEGx06yxI+
qMmt433wc25iW1ERrjJ7CjylPk5gxN9Vl26e3YnX8FUxvQpZmCcSHyscN0iPkE+S
FxOH8tBO+3F9Q5MbzBcTX+XhfoAjIDYkIcqDuon7WfhU3G0G1YPyc0a1JKF8PlTv
aeuHnM2E8aIVOWASCBRpcez1CZqHptxcRC/UTd2qPAQsVlUjKJHVxPMqKy1xLrjW
iY3DyiXUyIiHHESH4Qxdb7l4i/iOzwKRPJkJF/WO9JVXPx0TFWb2+ZBAA2DJcS3P
DSjWevF+xr9BzuXhT5Gz7wYaOxlThP4ozP2TEJjlKgt2u862x9Z5rUfQ9U8Q3r9K
2FyCWkv6ZkLGnxG/efhzVjcHH67M3ZPJHcdBDF9beTxY0wthi/pIfOn0hdOrQ59P
uOJi3vzPgtHqtENlC1NEJp8QI5CydY3YVatPXyyVwBPha62yVOD0Spsbywb1zSIa
`protect END_PROTECTED
