`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+wM981/75wvt04sFyLovNvGHi4oHA4miKnOYSnNwL3PDHhMhTHXeZpivj6C7ZQu
1wyz/C1iLRY3jq67LUFYPx3MsOzOVJcimhEV8QkSRB4wxwW3CbegBqutdmME7kQc
RtgRFIPqTMrllFQgN3ClyIqvKjavRE7CxUFZOQ1RyAVosdFYzCAjgxfoSHtRF3yW
5hkyaLbSErsCroxqReaoKL0fEoiE33LbcDL/VG/Ykm/0YU/rpF31/ZCwrXqQfcWj
eIZYpiq0kAkyFD5yUzxiJd21JCP2jI4VJooDjsrVPgH0wa1zddRacTnZ7rEtY8Mq
VnFjgymUySPLp/sw1eMj41WVJUNYO1YmaqiAR6AWLNQnvVXKCFn5Rf0/T/BNYTr9
FtfiIe0oJ/936J+5DuFuR/hEqzUdKqJkQOdbGPF5NzI0hrgK1P8dj2qlh+V444RU
UogzaRnQk72qike3mpyI4JVfdcGcYbaEFbHlORR8QC/DYGa+Dmw+LR2AkZKMEAmn
3P9dwaKx0ia68BbBKxkeGh5EQdhFwQKmooComwIjInzzJQtgyv89PkHXTDw6V1tq
KTmpuPtMIJ4Fih55cbvnk5u5YTbyDyZpqupLieM6kGBMY27WSwjP+wynYZmmgxyp
QgHZs4cevSsIuZGLhr5ZAqnZoC+Q0xIIezXkXbaphJlcX4ffQgsmWpDQsivvJrzo
UBrzg++25TySWHMxaXY+6U2YWQ2T+L4BI7hAVMAM46w+41y89gSI7EIsPHOG6pwl
a0xArANPzq8tTZqiHfYpWUBbR07Csp6lZvm8tNiTq9Mk2xcRfs/EP359f+KAnaML
LqBLyL2KK0cq69apcei6Bqc0w4h2iBq6yRMQseYmwAJQ4io+WZG8GyWC4xiwMXvE
aWeFpk5WKfxBXHI/OpS4jk1MbQf7x7OtDqRtY2DJidv5B5Fxf4M5Yg/t2ZT4YiT9
3mJKmy+jpo3/wDB4FsxPX3CxjkRUfjelgZw6JoGhgu9DGt1i2+lUBdMi8wsYL02R
S2jDvRyjqUwUxlZWOjx9H3qleGlLGegdpKO/mFtpB+NsJmKvettnztYhn29OkkEw
a19PJIwe7/gnpSgbacCOGUHPkGbAEzktfrQoqyNih5f9Lz05fxeM2Dg2hhpBtnQr
38jj6GoRs4YWdAO7T6PajfpAwr+hs8dkyS/s9vN8bnvkECVWI5eqlrgjmKRD29rD
QFONeGUx9dXahLIWeVGQrNTW9L9xVmoRj64+VCwTaMCvEFjjnFXIDxGdNWWbiDbd
7oDfMa2Q03MwrjVoOVLkBRrEACtIB0CuUql3/ra4mmK1QZK7Ln+aAbknKX6nEdlM
ao3Tg43/63GbIE9T5cvjtJMEUv/wN8Rz6qex3WAcGVFF70HlAHGSFCTMDX9v8zEk
uUD9ujpnHcHdF+MpplIdHaF0v60894AoIUCFxse5TPtKuoP9TE2XOUd0YVa1xcZu
NMbLrH5aK34RRFzG9dGYrD0aywuu52fYj213DZGmi9wT8/HX/CKu5gzIfaiHtszl
5R9eGY2QX1cbWlzmAQA8WnpNVKoUq/KQf7c6xd772TuGssH5m7rz2129iHr+yjfm
mw4BCSIrbQgmDNAmHKvlvEPDTgDKnTnCFEPH53V+poaEabvOTCYUS61MltRmVkqV
JJmb+wtlXFcYWfxiqTeVha8FTZ99pzecQAQd3I0UgV/4BgYk3PKT6mteo92pxTyz
`protect END_PROTECTED
