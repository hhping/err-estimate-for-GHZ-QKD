`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAYxf1skzR2ihF3IpnLve/GCOw5Bt4bb3iK+vDhZFyCZ/RLZFkVPMj2My82b5L0s
4ksbdnfQ9/fvy48yrn7yGg0QqUIymMyNuaP6vRz/L4TJXP3mwLivQ27Aokx/B3C5
FtGcF26WiuqFLXYbh1fMSPlwtiGeheahDNk+tMLRXAt7ZnkC/DkJOdS0gP/8iOWw
xqccNC57t5DSudeLIniPelbsDsGPmAViCqAZsMiQjYT1XhWYbT2yCQyPf981SSSY
1SHMXJt0oCy3tR08zb+DOfrRc9Pc/WGJWj+lMYocrPhDYjoZVzxwrhSwSbkfEdtr
NfCpGvghOvSQQ8tGy0RMgGRGrl7SPI69MQk6A6ZmoZ1ZGUhv0TfS5wIk+/CqQ1b0
frolRs0gc9pYoHH0sLeRi+Dqx2bnQT3Ga4n5OVPYfNXKC5/xovz5d7P5O+9mKQmi
MVuXS2/o6NTy0+I7I9HaSvFbGEtjXytSr3ghItAz1t5WbEfAfDZa8aoSxBjAuPfD
rDMfyZOfMUciMIc4uCZnrJuawNEw/TXQ9KL3Gyhx0m4XisiSWgWWH+NDCamAotdj
OTIJDPBysFWtapnriV43mxNGEdLXgIhqkNTuqxrZCAf6hjNriz6n/9gJBJCDc7px
hXovblbsEpgLw9qElnugJ28yIADkDV7mMjiU9nxsj+Z+m7Y0e1AeYAAyUNdIV2oI
XAQ/q/BXnhEMO2fC26CzvLyLgQHSrta2KFACczPWfvXqftdtpYO63yhzoJzblOWc
W7lPXpNZ0AtcsUgj13g1/oMSV0z1KB3v+eRXK1VM2Hli1uPRaNLpYnJeF0PvAj9B
9imOafHrl0ZBW+1sq01/z8f/boS+N2j2h7OdQunvEIDr0nYc6rgJD6HI1Hbjx7dj
pUT0XVq7uzRVnfTfRqE2Dm7I1wrQ5f2TJjA8kVsPJE2QXvSJCvFlFSn0rdIMyTjJ
YLAwxSPJjDPv1c7yMAj1HRn7mQUMxZ/290HfPcrs13UNtF/bgE3JPT9brgXQP/yf
ok3211+dJEWcrVVxvGAdMSaj0fuLz8jhGVXTlI5IfAK5Wi3ufq6B6T9G+bMmGkHj
mwQKvyCcbqv61fp1vdO0NvlhlanV9v9n+V+zoR8APR8te9R5fTzhAd62BldU90la
Uw/EBsWnc6KYV+ur4ZPncCAebSDa8SCIDcyySuT8Dh7Z6qcOPeo9tYkOnayveOex
lKVF5WkroK60hvLXkM/oPk3N3pO43ZzTJ+SQluFszqnZo5Hchhibr9OtHKoQebJg
qmbap2XrNHI9YNEuF5lM8ydFCSNim5vHk4W/qMm0d04z8xT+iWFurWBOXqFednU9
EwJ0ubPb1G24l7Sy/hA9wEIm3U5TmqkORyqJS3dv1I0Ic39elvQSd41vopEntxjy
maah66X/K0hMi4zh6+Ny91iR5H5+DM0BOXPbYYg+NSri0su+MgIkNERvRlThOcK8
vgxc9NcIX/84m5dHWXC9aETXh3gV1b6YoTKqCKX0r84MGCX5uk0wOsQ+HfZZT5xD
HL/KTq41F5SwdZVqR8rAsRjcBB+Uywc6OOmseIY2Im/DFEV3kTgocAmzjYmASUv5
5QAECkvTQ5ty6G+YeWPFsXtO6w+MqkwBI2fuY1hs7xPZlUjve9gPQz7Oet29izCM
hGajGQp9vg5qTS/9P0yQBw==
`protect END_PROTECTED
