`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hjubawgg5EIUHbw1uKxtr76QM80ZpE75TULI3R3VzFVS6//SD3/2cc+a3GmMjiwP
PVg3mx5GWTIY06/kUP5rSNWJx+AwTVdxRAbjfQcwfImCLwZV6T0sjrfSDnQRR7Si
tF6LzzFCESZilyBGcf3V7jNSmHO99v8pUJ3PmpmsQRkKGPlJonmR8ZOJ9/P4SiMp
GTBg/T9YKZTQFThBByKwhtcxp12Kb7MKq+uHdUAbvBVKtQDs7mxVUoiv6us/mAj8
8xPPGqjC8OkKHA6zSv7tBV9Vg81NNnZSi1I8psh14o7ifHDn9IsXo/uOLQ9Zg7c5
6AgMS/az4r+5wcLvaDbdNgi9bcGUCEG3kru4gwX2TSAzSPgcqKDyM+Rpie6c6e8s
sikdQo8DbCeE6ktIx71wERe0X3m2Q9d1mn+X3YhQ52PAGhsnPCO7yxhF3KIduMFe
Bu8u5MjT+SNglNPYQ4BwKFzFrv0iPUFW5fb7jWxjZb38DM6d7lNc1ZPPoZ9wyPmC
0bzwanr5VPmqzWd+w+FLy+hlQQmNcZs98qrr8O7wGWI=
`protect END_PROTECTED
