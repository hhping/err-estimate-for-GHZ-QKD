`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXT9WefecjX7hTdN7IdeT0Etd6b1lSNABDu5cfcwHXjXSZEEm8wl/CKFAbgH9Hne
yVt9go/sA2z7GtIHhnDf6yKK0TMrAjjyQVFYwBRRK0RtiC5Qn9XIUFYbRbdOoJo+
tBiCJOk1ej9/UK9vNGWyZaADT3OpTOyJ/VyNQ7EFu+0ni+EO23D0ffbDlxuItX9Z
ZeyY7LLDzV5OHf+GYo7kXeK/EghUXQzi+Q7SzUvBI6C0+u/9P6awZtlHdmJZx5Ke
/P5QGN0bOL2YmBzUghtPQpJeUOMCwwNAf7s756PHdoWCd7Rl2V2H+Ks4LHXIa6Yc
o4J9kimaugfGkOEYREOy9IFcG+ATmfMSVRZAhS7syN9TTBX+X2G5fMkyDbO/24Bd
iR2T2DFiMJE995fJV9QmTM1h94Jzv2ke5mp4Y8V0GLZG10R6DFjHFzMpB+8bQG3Q
W+WqSq6N+gxlGRJh44q+x6etZcwAfzSq1uwvGIdFUqWbH92Pas7uPfzzpjbk9qUq
/5DH0pYmhrObEF3NeJ85iiCV5aCPmn6uDigLlNqwIcbzzseI2xVJvUL8PjaA6Dwj
bDnO1T2fk0rIsa2LqVPxefayGoaF8Gr5JYklvzuJs5ICnmtHwNPIAojd8I9kFKPg
3QvpdlTPpgdHhQJXD7Xa8XfdVRbKuXkOX77fdRL1+T7JQI8Qz2MaWzlZmqLj8VPq
+8CZo79OcAFq92d8Esmqnsa3mYfM68DDMdFbBjdepX3VQfy+3bydSyB3AFgwUxU2
Bfd6HGQA8WNJ55i75ULboAZd2GMGEK4q1YE6brkfOyy+jU4ucuGJrI79U6UaA6i2
sWl9/ve0k5EsnFlcxftO+VWKNTHhC7N2nrd0NhTd19I1tqYv34MIJV/J9KhejL2L
G831EXI7W/Zk2n2QBvS9I07H12pwWFNL5ydXRBZquHtt7Yd8FAsJjhRJsLoRyBn5
Xe7AcqQ7opZowbj9o8whgse0vt0KFVp02h9Rx0Q+AAL1ABScJwbduHu2If3txlJ/
lfGHepdKmTtmLBSXkMfltOULrNhrX/9VW3Xnr4WkEaSGDr/IaVAxqRe3tgoFkg2M
RtpMbVlqPpMXXMoBkrCK675jtNk09vY4v7g3+wE46SRuDFGS1xmALsJkIExJtpW6
tgG3cJsYc67sXOz0Cb8ZOIZ/F0tja7SPB0jQAs90bNiVUb7BYG2gfaWoHWLV3tAR
ZY0+IrM16xLIYF7xmD8EiaWfT+x/8bowK24I4icXVNtW+gSwJhntjrTGdr836kNC
QnIK/Jcfc4fOGGC7CKDwrfs8x3/8il46bbwkrQxNrwSmwNFjujYFSjw1LSR431cA
zc/O+m+CNW2hyk+U6vL2UnG1wpS8IfWp6+nn59h8PaQlm81GdGPc+crFfsDD9lkI
Iz3QRgHnZNculC0yCf5J00cIvAfyn4MuffrQSU1ErSoEbuUXUNIPI8NIm2SauSP5
QN2u2XpFMC+hDcIoC/qrfkVGiF+wdIZ2Zvg8mXhT8YAYeh5aVgBkPd5RyAokEiAl
t6PMbt/NsgXUg+jBCnUBsbMvovJM+v7NUB4QM7Io8nIpjJoiKeVKyB3D/p+QCZ98
8/vkLfHLQsXN4X1NoG0aS9Eg1b/tSBMzjVxn2bReV8qCsRZFSdMt/y8rt558ry5p
m1pkfpDD2Nl3d9WYCivLSOL0KxjWUQy3T0LzLXt93MQtUzGB0Xg+LqRtMTht93O2
HWyIRyYEC9ckWZ0Nro43IqzHgUZDn1b1TEFzdnlD4IGVq/7UO+FCVMEq8/csiIk6
SLBrs1t4BeanHsQmGX5ngbyBRNVpYLswif4EWQVIyTGEka7eHYUYLjd8rIDrYIDs
nPhVObIIIA+8feDE781PpnAWLAgNiQv8Q5nKMKHvk/kMf669ZGPzY6s52nuKAkYA
DjLlz3YfVWyr/jA9j0EJZ/MDaRoGKnY8w6GW3ljcsyYoMA/VG1fksxAUK1GaUhFf
v5Z6BjEQVjvPD5kP4A8zwtHEEjpE/zhtVLRRj5QfLDST7D1qrwUle51If4FddybQ
AT2fFyWLqt02M2n4wDlv0vP3oYUOFARyAwyNJSA9da7VIg1YW+9OplvFyegwN/04
YpXE61fq2VcbStst8FpNS9q1LvXXuiwCDu2RotrPMbUYe2HRewfVVtPp7fDnTN1L
LQAuP5pRBGs1gJVtA1alvrjkdktlQ5HKkGvHaZ0NHD02ydR/kme1QExmAK+XswIH
PjkufK3nbgwnYiccmgJVdl1KnI7PgrG8mv/XqKzY+sNqXP/xcITnoTPIaoSBGUoB
5sTAT7vXPGWv9jVBKgvx/Ck3r45TrHWKHQsbW2RbjNz8UCQPcjMffgT5wbiEoCN8
3QkpyiOmiEVe8FSdKbuIPDj4s3qFPkBA5FCt+FZtjQnyeq8JN05y2SyjtDOHzE7L
gFaX/fsgkAjJc9H3l/eXuSY/MsAFixnEDtLEQ3to1x++G3NlpWdshZkq66BLjA1H
EBeXcvMmrMx1FKN65ev6ccID6lWCcmc+PFWXWtMeeKlhGxGmDsYgZgO4jH83+Y+s
kx0wzrfzq3GZF6Id0NbxmkfdKFdnyCYXIZe5QpHI8d3cOjITATNJqxe9DUDt2b9E
OntOIXNN82tNHrgIV4z82WR1j2LdR41k53j5ZJBTKgQFIEvP9LY5F+Kxjjr/b7RZ
6ov/R8liRE0Z5g68/H1G+G/Kn39d+pp+qY7YOywoEfs1dM9jqy2yHFypBCusMYVS
ZEfYwSSlO1yiwmFgmgCkvG7aDpf91S42+1X+zFHHhU7YfKuOzYcTnZSuNtUa18Rd
l2p3srpLj0/2Lxj71MWb7X5kwRNo42QasgAdyUVjz83dlWQiX2PEqi5DDl3E/x5r
sYvok7zG0/zyF16juGESI/gFlBW0Rw94am02cLETc6tOsB3F1W10PBJqWwYBwW3r
ztacAlkDdhzXpAUrny7c18w+vxEpC/s5zBRRt8oLQpQE7fi/ttlEM/4uwOZApvJH
aa4jSCJ+8+i9b+cxjH6p0RHuCa84ojB4YQYeGbNQt31O6fXGGiAkxJD5DsofApNk
VMTCMS1VJkP5NhzvFZEl7wENSTx9Qqjs42tOsTYzWSTkKa8W6AsxTQEF4qgvGe3s
Hh89VogGIIq7Z3VjYtEbWgPlQkoTYJbrZ648bPPv9HBHBHA44Ga0fXI8LijLbR5c
sNk6DuUaW+4k90Vfr8ZpNp5bGwymc8ByRgvKa4CK1oBTEAhOhBVqMSdUt1hprL5w
xkwBGco9Q4N8Ajk4DqhnvREzf1el0HmpBfBgLLcyVxo=
`protect END_PROTECTED
