`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KT14eW9S88fh5Hsn2MvsgTmwBKUscYwt2DgWmKi57i+936zq8mYFc6BV4O3prAJ7
/7VSsuuGciHDKtkb+TfAZsA12F7afkQu352g9k9MIsnTFcbDAVeqjoeadOp4APtt
zJu7UdrvG+aEj5/fxswBdeJlr8825W7R7hjqACtey1SyJbzvq61RlUVzIMC2cPce
klj3ws3/5OtESo2BAC1ta8WIQl7fyU31dlXmmyS5aOjC9VyYjQG3pQD8YTHrUlQR
qCI9+528hPoWC0eEWwYXIHUJCUDzVQpI1/rx6RrGbxGfvHKgZZKSjoSeVW5try0R
Um5efGAGmTT1M7bT362hpMQ9iDk66KLfJw1BHdQQfw/2pWz+LMcvn1mOf7wynyC0
PSmPNSr4KBwhyE4ZGKsW5Cxdyyfr53z9nO5hhoirVWOBQcpe7RGFh7v1CWjS+vOh
0+d8JFQd+1BC3yr6uMBOafTpJwHUqSgCOHdHDUIbBuCLVqYYL11s/91SinYCRdRw
3Aribl0kzylG/a/A6y9p+g==
`protect END_PROTECTED
