`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iK9PgdozP2qQRMFEwY64fetZu/HMSKNGn6RWBkt7c0hzjg1jTo2Og8LfCh8sQ1e4
yapmXwYWxNtyhp+Y6J/FK/hEFjZLmBWL1IR8Bmgo5iKo/SftR/pUuzBtiBEpGUil
t1CQcziOMPEVIgM77mlRh6dHFEQRbm9cYG7XBMcviqfA6HU+nTNWpaoWGG/MM9LE
fFeFWK49vBgj21PL1PpNoBGgoFifVpF59cvLxIvTTADbC02wsoMFaPlZtSEblSuY
0TNbcGXVqmGQrQZO/JIko//agOLikm9U1K7r7xwqchDo9YRIEldEJtb/V7MEeauf
MP4Uhy9piRmNIAhlOQ4CyRsDgirViULGvDG4bQdEpMDEmo4kRJxRHqPBANeweJBG
4PIqIPm5T02OA/Z59YdJ26/XT31nualTAjdHfKvpZWHKMx8r0a7DpDTvJnpbvoae
JCcqR1WdU/KlziBrDDO/d39Tj+4RDAsUMlBF3X0a0d0UhYbEMXvHqadRM+BG4W4C
qzMYtgO5HN/hXXNToDFkwP5Y8Hnax8oHeSwVStASOnTOi8cVufLEgZ53RmgEepjp
D6aIIGFVzcjmlJF8en+gjWE874R/0OZvKAmVGVvdhN5tyniK/ZEB8q4OaSqK0BUG
Euw/xrQclg7zwIecjyNo4o7COIaOHtiL4ow5SJqIqGQ=
`protect END_PROTECTED
