`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWSgfYNSTjYgrcK4huv08kiknrD+gZLYa+klYd3V+6x/mLTfUaJhf0UnwIpzNRex
uU40T0cFx3JPgMuUo/hlQVextoYADL1u9ZIoy7Kq1ZQawcW7HGAFmfMiMj6boN7a
wUQxvTAf/zG8rn+I5BJ6gEvZ8V531mEfYJnCIQlqdkldliZor5/u5wp+j1i4Wf48
HXLsIEqlqTTtrCu28n7HBzUJAr4sTYxtLdrP9J0B+ScT1jiCnRW8zqjojU5ezZXU
IgCGsMnRJ9YDUWArcXw5x3rnaf0XCv7LKAlw46waFkHQywTyZtRLve9VkPS5xUXx
eSjqIa1UpRlfR5NOZY7bZoZ7Jo0567nUsJ+AU/POxO7JSWqjvHAaVuQRBUdLlVeJ
FQAkkSgDuz9MQdOf+jCwdgsnPw6uLwQRKLZgdTP3xtNYesuiHAw/720IDNAwYm2T
k0y0SJgTd8xqjiV2a3mENYZNLK9Sm98AVRRxh8Rrol5sV1Brit08Slfk5XhNW8zh
ukXL/KG04kuCrwhAT3SuC4nwNUcQfdqkYM41wnvE7EVk8Li+rUPS0iI8oOp416w3
+K9cCdDnwnls4QJ+6DOg3GJxT0Qheeb0WZNt51bHQgOvbePSFPzbjRCd0MYShWr8
phIjtC6KVGsY7anF67AC3K36twQvMydlqY0V+RjNUx8JsQHCiiAvXBseDW9ytdCG
8D1GBofAJutLl2+K5xNYik33IfArZPV7vDDDQAAMtpcdYUXzOzjIu0CMHsV0nmqX
Ylv0o8Fu5Af4QZvDiFoqvqSvVkzNsizcJdPm/L4zTcDeBFTNFEcIW9yEGIOMhmU6
kNbe+YUTg/z4fEU8KJRazD66wT/LQp5HxXCGqGEa6LzZV5Oic94Ym7j2FxTXwsH/
o30ll4O59N0pRRllprFX4tvCD7Dw+JahR+Gx6H7QlZ5/nSuree5ITuACcOdfL2NG
bDWs6LfH+hLeN28aXMV6cOWtcCLg8ZeiM2NzLymtXqwyxqHBWTGuxrey0UflBmCY
E5TuKGkHmrRCYejYKpN3COmrrVTepHDcqIb66QN2DZdxlngZlK9EevGcXbKQNpIe
dKNEAXVKVX9MRyH1z5ZLH9RBAN+9CNWrbNSf7lKqbuaJy6sFHWKGD2Zwl32i+NRg
61UIT61vfDKSOj5KB4I8IFaV/+22rt4Hs5ZZgMb1nwsH/tZbMpQX66kzrtY08vRZ
4eiAccXZqjUK84xUKWyQwVjm9nIk/1ID7wIqloVnosg4+zmA23Jgup4WWCBGZA5j
tUSwD002NxoYCp0PIav8un2cXzQFFWv3ktSqabV6uYrgYQOOblXA+Si0lGs190Nc
7sN3FScyF06sx6vfHNdjpvLgJRwJuDUKjsyF4FY51nZgjbzk2RzazgRNE5W7F7Cq
LclzNJnUTXOnb0c4uz7YhAZy4AzCGeVpFGI7TaHJWQEv8GUf35dMAgVwYQ0i1oOO
lthn7tVaJFqzcwEi46KjU4x2Q39i3vO9dH/LLynkeATg6zwZFu1zwi2YXQgVT54Q
cFLmrXVueqn9PHifnkWhK6aBFm4xFg/y2vQYgmhuzfIl0i2bglWzEBEL/D/paUZ8
72IvoPMobLjh+8azWIn3RfQNUW4VzUMvUcSkUtG97H4ilJJL5rfzGGxT4yL/8GtK
qtOVVZGHhhSUKbdZderlKPVRc+tjkyw7zcz3eUU4Yzvn270mZGgZ0LRzhXjxpIgF
kXTDB5Q06pcLsM4iKEyKkqJQs7Q00DQW7cyNHWO80cfahtM6i7EDuYbGEQU39AvR
Rf/Fkig0z8gvJq1Lds8JV0gcfD5+GvcuT1BEiv79QeQvkvJq28/Fs4CgZ2BBSfok
z4DfoVghgoFNmkSz7NS061xVYhlv1qeaBbLPRcXAA3wQCotejVzLyqv7oC3yLxPr
U7rfP0YQnymEdHQYWqd596vHpJtvbH0Dby6y1+RYIR4BbtpMhkKTToq2bF9Vo9a1
wrJMfMzr4L6VzZyEJmHBEqrFF8v5Jawzw6sF+JcEjfVfrH3euNvzZAUwgeIDulgE
7T/EvGxM9YDVKpb0vfWXrK1FpExZ7QVoluNU+AhpM4jzYtusV/UmNSuQTVdAFa/u
EhoTS93XvmarhgX8i+kK0Ja0F6sEQb6J27A/rF68wzR5BLCSqHTCfAMmmRkCodKf
pBPfxw+5fPqTLEFPKkW0gtxorwuNrpz2dXbw/gT3FVG3QoJNN0bqHJtkN4cIWGka
3ijGiJcOWuzWTSuukOdpE51CBxYH9eSj58AyleD+YjCUI5NtzM8POqvcPw9muTWR
9SFrtyRnxMaIl5G6sF+ud0Cuf69qD8NUDDREQE7Vwvc=
`protect END_PROTECTED
