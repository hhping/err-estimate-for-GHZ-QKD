`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUUMQ0uqdfX1kA4EQdqr9bE23ECNxv+jydHB1whFsZ0W+llSE3W+TL8f/pLNsafh
hSkWq1BS86dlDzUV5NE5xCoRHEhGm9HkBBPskE3kjjdL3oBO1wJwiB1TuwVBuISe
TA7O/+nhp4M2EdF0wIfeBHEz8GTBcRDPsksfbSjvx2P/wTIb6zdrth6C0ynd2KOM
LN5YdY1d1wreSbJV9H2FAeBQ17EzEyq2V1X3+qQFRH9NaHNk+HIDxNMJkDKsYZnM
M/POOQXdkQzaOGFnjOcGAtB8dFAtK70v0AJ/x5SV5Kl5qKsZRDwKvDBtH9F0dWNj
Fuo0gSIDUQrqxh5YBFbMBYvlBXUg8KavNAI6pUVhmoRDA4LfEJoi/Gm4E/hl46nm
ytkfn9sei/4KMC+kVB462yqv8qmhYraAs0MHz2X63DOqT7PB1wXnbvLOn8OmBBot
l72/ybnAn6CJ9cRtSZyMYLNpalcbUf5AygIKzpZHz0WBsb7kbF8Lq+oD37a1SyZU
zVk/5T6z9ks5HSlUbk7/t9ovOBML4sQKjFCZ4XBco08sV3Tt1SsqTZFT9gePWnfD
E6s0PP2RLEDAwx5+FXAR1pPqvvbba8Ghkun+ReVt2prFdtCKASFHf4CWUqxz2n7H
q5UaWSv8qPg0Xf5pmrshTx38ymL4IyzAbBskbGZvGbn+B8tiCnb6U86Z8PaHcvRH
4RFx8vY3AHO1ugs3RckdFhl5/G3AK9psv9LX5YqNHabb59oZhCcawRekJodOpWFq
y81CzDIh2s3AL53e6wL2ce/lrMqUD/s4rp4k2DCcz/iDaggBT03tt2RrsmBtOGdG
BER5nRZulg7yMbhZSmpVbZmJCDbdj01BQxQxqMSVbfRwAfuq9nxJ1CMTR7avNv9M
E0KuP1lTq1XDg+5aCF0l48iOO48pwURTegjdj3XgtpjRDAQQOrgichb0WqavIiD5
SY9bAt8YkAVEny3ItrilvxSmj5Ql2iGXlYAZ7x4SNvubwgavjKuO5Mk603VnJxdI
Afukrgx9nQyc56hfTCosDlqV4lPISCHqXtp/XRVpNCqj9RPlwFJDMsQ5vuE7XQHr
qBUj4CAdkykMyZRQ1URJWpiTdzkc0aQi8hJjU0d0ln+Xq77tS146Cxltz7Ak5sje
WZ9UQXg8J2AX9dJKkL4nkUwNm9EmLMFjZIwaETFM2XaEocnf5MHZQf64+4QdLciP
nsq2JODVhL2ATuaK+9S+0HkuGxcdiDghSjMjfuPStkNzbfFKkFWE3UsHKMaZFHQd
`protect END_PROTECTED
