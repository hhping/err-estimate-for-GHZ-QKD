`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btrM9K4KRDmLCl/aL+BzmU1/ZaCwutqUyH4TC0k1dkkE8vbGYYBJqKWTmYIqBsDM
TpNaQJS4GBIfGpdcGTX5Et0bg3NjQwAUAqbkNJUmkzyDtgvvbrKbkMQEk3joH+N0
Rv9KPWvQfhsco+FWMPUNg/lNyfbn12GBi623kyUD0AC55Wzoxjx86OlC4Bl+ONWg
MQbgtkv9lpJZa3PKMYon3ITwY1gfv9dXmKkjubAgt/+oqsUVydd4GiAL8BWBSYay
hI41JRKDEhxsl0vEYMN95hMzkGFeKV0qU0RFGb8n/pb2A4LQR8kuyTJWbGBS6KWb
5oXGlpyx7qV9wxtJilcleIyYzozGFhmsnOC1/uHnU4boKg/o8cy1Ns284mA29gYf
3fLQzFOpo109L7VBnrD/BIg5hYA18NLlC/IzPBmncVW1PygnRSqO0eQeWgH7ncw6
bEClczEt5KX89kIKiNA1ZDpLCmus+1ZNyFi5ueAPUQmdeYZG7RaZ9Xe6XUY4WaTp
theX7TarUDMSfK3XvqNJv35sRk/u4xIk80NjsqbPyXHxPmMqxuuOugTX7a+3zgco
PdZ8qG2MVbEUFLV4SXCqxRIhyxBiMnckA6LrYDcY/C7IWdnQE3Rvd/SMDt9DakDk
7tiNPBFKhjIuszeO+GTvG2lFlZZjc8mXX0tVUaovRMTf8p3tPjoy3dB18wbC2ypd
3YRc7PHHdMTP2CP/c40JE51qTSUb+vWeTc4P2QiAYYArTLIU72+GBgUWccPAaBZn
ZTphjs1oR9CclMwaoJylO55VejvV+d7h64VG8L+rZZme6rhSk1YQw4AdvV+/MZug
2TWGjqDdgVRz1qLFIR7aqgIuQpp61sJd3kHkL1WqeDn96Qfdj1xlAu2kutK6NbeU
JqriGyO6m9u2JnEYSNoCbMrdTPRw+FWqrDbtDals2wHtQBeBhJg51oWBdfSf6feA
YfLMVC7jLuE1xo1LxErKl0z5PTaJ6722Qm4mexEbfhf500mVRjK0gvWPmAiEpfY4
`protect END_PROTECTED
