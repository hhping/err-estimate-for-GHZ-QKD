`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lqHDpeaRmkyO6HFBGKi+qLn4usyi9YM4Qr2SPVxKFWCmKL89B4SkoR5ylJFzOrr2
ZEEu85jz2HwjKrkD6Ja+aI9yOYhG1ip+Q3d/RVCl2UCiEE8YnMyBFi0HIXwYhc2f
MKpmEY7jwWWwHagb7pzHekSYeJ/Wn/kxEiv9GShQxX8MgzVf1hOlNe4xRjDMGZKO
pvPi9Bt5pwKCE+EXGM8j3U+eeWo3OE6Nehyek6odeAG5EQ/qRUWDQV7nqwXXAqAp
oqZ1llGDRThTS1EI6xgQk19OSJKOGSUly8quLQ2Zs5lbike0JQzY7t03CSBzRowW
Wp/oziP/Yg1GULLyEIV8nX9mL+rqoayVAYg8EowLRKiKjXiEAsmEF5ErjmVOy6gs
yMFgsURsl3c0W5SKBzYeQ+/YxHcAEs31wz2aALFSt5gGG3Wr+W2eZibAyTu/swNt
sDC3BpkBINlEkgS5Cfk3ODrnOYq0sIGUy/3WCCcT7llRllD+mF5NewVW7bduXmCT
7VCvnjg0jsxJu0SI3kC0XNlKCw6HJHXOWqsprMO47WJbeQwQaD8Gscl2UHWwtlpc
3npnk3K5Py9JAeMCWCTEMTAvV0EfDYf6WYfGeF13qTGgpahfw/EO+wnyn97RsnhI
6ZjTh661XSOkKyq2PYg6OZqz85EyNChx5oZQjTyM0i5CoW+lwqov80OtoiKEKbko
Dha3qIukyZ9V0tk3rCUa+mF8HnMwR/0oTaMWF+Si9Oz2UuDv4rBAunkINgHua653
QD8ytud81RGhrQwiG8MU5Q==
`protect END_PROTECTED
