`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0r78YUYO0+7ACdSVgOGZbr+F5LGnjMlwomd1ISj7lbU4vK9wcR9eNPLqoten3e/
2+LRSw4MNF0Y54n+hYl20kdZlPZU8sR3GdKWekMsfD2b0gtSTriYDeOMaQDwVEoW
s546t+MmnA1lKSV5kjztbDRTbDVK7v4QItzXU04omn6+lop/zZOwZVilAMPQttd4
mcTHMcxH6uPcR57ZXEUhvwCQ9Eb2NtOa+PPi8HqgUybiOkOX0FkYGSIH548gQD14
2MTsQp+6dLhq8k6azyyKOA6eKvLKzYRjd6Lwlao18ELhs1w+hnKNgcECKzo5cHrj
XVA+yyBlPkjDdPqAk4hYJc+CtgkwAV2oft1hhSwhrrl+ptx8RtftYX5nNW/Z+i0N
0nDgB3Q1I0x6yhndu0ZiJsXFFK5Di6vuM75eR48YDbjTgKeQHGAy/KOdMvoOM9BR
`protect END_PROTECTED
