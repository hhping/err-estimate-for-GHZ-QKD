`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFmBqyoCIFx4B6700O8FLwsNXIdUStMtNLnyF1QQRXQP1Uii61iXYO+R24XE7mCd
5azq7ZpboTAoB0/U023rZQdDmVVuHnhuhAJv2e9yIo61glXLc468ssEPuACYiI3C
++I9S86yVspRsyvSwXU1dnr8zXfut9GGICgs6BrqATiRrpapfOm1JMl9bI1v7bY/
CNEKVZa7qe3/7hZCcRU3PgiT+O1xqHH8NfFpHnwpmtWxe7twIcjjCvIMVPCaCZY4
hlsGngZoT5XPO6ObW3OlfVwmoiSgcDzheYs5sDuqrBjwWeJQvC2BuLFdMi/zYJ4P
VORiaMcyF3q2tkOo9mC0ZQxfDXTaexLaSBZnafrme/hwhlRX6SGsLOIwZMk4Eje6
i+vml5Xm2985Z14ZNqXBG0JT0Zofuj0Dc8XDN1nLGUxIL99x4EyW2L0MZVfidPCJ
K+mbHBe+eQjg2cEfIslWseNg9ZK7hJ/c3QysYVuhFb3l93v5HTNt6lEHa3rXA/r2
skTDdy41rfAOrpRG26LP4NyzsHflRDL1Bgqo3NAo9bklSC1fpOmJU/mQ3AHmrix/
ZlzIgdc/6Kh3Xx4iAV7VRnYOdJzaWyMnBl7rda9xr/wDJzFzTE1bk9FY0Pj2BTYy
W8G4LVQT1VdTPL8yFS17TvAm0PrfhmXhMHtcEARAIViP9aUT2pgxpD0SC3nY+XjA
faJRDCuno0lh8hNImgmsApICkQ1F3P7RgSlkhKvht2yJErdCQnVCQW17q/yM7F5Q
giNV/5wPFP/4cz06iq5WK6vbJAU1zgQPYZN31lb+CkOoBwEkwmnjnXQfdGIPKB5g
CbjhKi3ec6fuLjXROYWu189EtO52WwhRcGmocoEx7JgGMLKobtgRW0QC4k+V6j64
0jIJZqwrmxQxjNG0oZzyz+0iho9mjrwi1CuB43Uq6XIo5FmKOVR4bbd8nR4UooRe
Dmg4v97HwJaeebPDppOF7uFyZkhcNK+NGxFTXAWYld2tx8T26+BrxY+eSPvbG6Z9
dG/N/5gignjfkHgieHyfeUXCVZW4AjsAb/SJg82pe3kkMXpRjqdXijcAZEMOvFZg
ENLcdPft09xV7YZQ6Hk2kNNFZjnczrqlbk1B7OYjSAPujjOt8JkJkH6n9gvUy7MU
HRejGDNkPVjwzirpuDloBGPk+NBrwMpIZCt5OU6hCI4=
`protect END_PROTECTED
