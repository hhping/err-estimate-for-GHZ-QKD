`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cC09rtrdM+vJW75bWrmiEIDUcjiiee38ckjlcwn2G1FiASkDiY3GyA0cX5D5rRle
aTqIzRLo1q1IIPrdw475tVaVrOBLKnpQUcP4+8cR9412Z/iOgzj7oM74RYgeQmAV
URC1nlqW5LUbonxYkZQWhHiM7FgseSu+9WetoS2ScN6mQ6J+sOQZI2NdZ8Xhje4f
PD9KsVejMOk5QepLLocQ8XVQMwL6x25E5toLrW8929BgekJxMelCuEIfxdr5cYyo
ImITuDvbBPTGmp5PJH9YLVFSbtNilk1o/gANOFQ2RBULcxMba3fOgIgnqI+xvRde
BrOE5fA0246jcP26Uuztou7jgggFJGo7nwnnqy3J/7bAXIM9lCIdEVy1LhhU21wk
DNH6/IwHNUZatt2Xv2RyYA+jAivqKqNaeFixAexXjpkW/FPScSubJjZZFSuTrS89
J+iGkwCk9GjT9hbbQaLZm+6Uwb6euLF3xsMY5E2VnX3ZehxcGBUv29oeAAID8Vrh
/YP/ACM4jm8cnevTXNgEnnlgeKemsk4dS+P9WgEC9xu8Biz/Pc6mA7RfBagmSSOi
FbZFI3CzkiE4I4+JqPZXX/9hWm/e2nMapqhPG1MCHV2AFmOrVbmokFBRgq+MbdYP
1WWuon1lxJc/FCiGwTBsXPIDjtcXyXAB3upCzJs6RfJESa0iwcEYveMzUue2E9XR
42G+87qskQ0mfCuN/KdmT/al4nkI8bgctUBjHxVR76OcLq3QdtwvVYTDiQiBJ3pn
fTcCACnArX2mgP58EpCPMz/vF+ykMZhdCNWPpknsw3AU5SDGT16xSBcR32MPz3P8
jYGGBi5EaYSo8+ZaZyyXJlSYQjRLyM2bWw2KbSqLHKpqAIHZgSd020GKwkmTMU3L
USR9felW8jRARuItNhbCxH77dylysnzlPUL5YIkWeE/tjkQNpLnhMQ5ONjyYFJ/V
/4ChpiW3ERtTZDPJHXRzcu6dlUnFgHL3qulNoMonupQzhbJw/BG/dj6q9Yo/Sw1G
lDfDs8hB/fL897/XQsFSS2ZuRWTNSHmaDKJMCtUg7LdVH96ejIV6uqgaQ8Iemnfc
jJKvpHblohBjTnylptqLoWoAxMjfLdmwRqK0TvkgpIfLbNJP5FbLriPPVZv7wWMZ
KxpjolTkT21VB/QXxK3Bs8/s8Ea3ip+qXH6K6Ixlv1gtzDQ3AAE23htcGzCl8OX8
LVKMK84zBjirU3yyw8BkqymOULRDY8MFtnNabHRsXZaPLEsexmfKR5e4q8UTA4PO
q4ieyH+FVMSw51Cloeaz6Lh0O4AUcZ15U3Kir5pfI2RFI16OxSsNb9zDnAXzYryN
tvvRQYEX34QrA2cnARpcdEBiXj84ry9pI8S7pYAyYlbJiK+LLtangmXlBTYxH24k
CmXt7T4brBj5LtQGZDLEwdJWBUdsya8FTbsQGfv0YUHYkisp4Ex0RDTazi4ZskCk
x/pQzpzFlNCIBdBFof9dwjateHdwN8WFxg3wmrzbl1JSu5EearpQaR32BlvGRHvi
Nga0ZcmtdGOhQ7qzXx2HVr6yFLg/gIkcwtrZxl/QVv5TCdswbW+qSudLJ9zzbwdc
4xAzQf/N204SgZEq7XGISsLwZkfBXfd/So2H3S0UI7gf1WrjsI/x0bBG0u5C3zB1
nLe4ODC0P4lAfMOfqgMIZAsNePJK2ArBpqkX/7J0ovhhbr1Egf/poVUi6HHEJZg/
qzqvBpVQyI5ZkCdBsbtNY27nn7KO948fGCGKEqrmeB+W5SXB99yzph5khD9/GacV
q8zVhoxVnFNI+pNxYsgM2TzWWyW4Le6/jpdOAD/c1KXEeZwv0hybLqpV7fW17erF
9wMzDPAyX4YdJTzAt9PVZDcStf0UafPsxqd/U0a67l9yutHexNzUqq3SsiInYt+/
X/asx4xJ/98EMJzAPt1/GC0YZp+Lfir2FIhRCWC0suf+t0NXuXpSkONpYC2nNhsh
jOEfLS+3aC9zxSdCqtlN9HrkT5jNMXBhFlesC4eJKA+yZaLtPP9E/+nLVEUsz68w
S9XtI2sBPrZKptmqSGrnHGNi11lYQEPtIpITm6Ksh6CaRI9oY/zdv3HSRP+JNZoX
HBsdYqUXd70aI1yeJIPvqNQPkIFN4c6K+Y84sGL07DO4hb++lYTVweoKARSMgP8u
`protect END_PROTECTED
