`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IS48SnikLu9cnkIZVA+nj1achqifjFY2z2c+YkMZM9VnyaX2Y/i9FpbdVZmeOa0Y
u/yO34U3ux4FF+p0u7f7DJkZ7hwba0bPLWvAOBaNAubttAiifB0HXJm7tmqvE7kx
8ge2SvXQhAXzA5ui8NLrm609vnPtwN5wiWJjvOLk6+0Oi+CENSsAx0IqqyiIVY/8
AYK4POUXjd5ysQrUU9puw7SaVAFj0YYDdMn/jYu1iUsoQL+3aiKQRchMbwZPvMdi
3cpJXf3iVZF8dU7sjLGt37EkWUTDHcH7wZZUFPjbGGCn9QHwto+HXCpaHHwCgPuR
6+YHOIvS5s0JGqnzQyjuCctM5FyMl29UhGoAY9cd1AO6GTMbrt48wWVv198UxUJT
Rw4BEpMej7t/9x5TJ5H2i+ycguu6UvFYoSx+xvRl6BnaJitpuJv7NrNE9P5ObArI
uHif3D8jm+F5GvXXsZYAPJOxZtZd4yT1N/aGDEaSGuGo8vWAC2qIw5hX6EJDxFA8
w1GbGdKjTTxX6WyjkEOAPxb0p2FVJCge59NvOC8+YVh9A5+YeG0nFVDdE4712pF4
jiN3LOOf3Xj4L6TWjkf3Mzb7Vy5W7BThzNgnAIx2cpQrXzP9C3OHPLxKbtME3kHA
URFANry5tLEEAzLAuNwgzm4ciylrXlbfZlzJzQgAg/tBMFRQK5LCAPquzRWg185y
LTc5NDydS43E7DIouhje5UwBFmpNwowjxdgpGb/m7T7ydPrU8x+FC2dvGzmj/rrn
iKEDdftm+ks9gD50smJRdvWfTn5MOXk6ZjemPWoLaDCPxz0o+tmn0mVog8eVqsm6
OrOyNaT1d6lVsBG7Pq4TsxSslC2IdTmCBMs1NfxMtXS8Czh+/FX+Blml6GKwSRpM
ESUi8bnt6cd1elOEqr/heQ==
`protect END_PROTECTED
