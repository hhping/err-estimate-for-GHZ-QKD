`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGr4tKfcCr37r7q1FseN+UrrcfIO/04mQUnNiMHWR4w2BA0za98WA1xDxOzfiHwO
ucjDb5iHizy/qJjHFBX7BE54T/BAyCWP+MfOt8eOVBffjdLOAGqITkKT+omt4EZf
24YOAQbmMtMBhpHv6rfPEhvNyke2H5ddEiHeWupvzblUYECSsUzdr8itJfCUKlJk
DlnijBkHd8vjtA1dI4DSc9PgivhjVYDb9JVLKFoJpbq1x+tcsZlnv8YtjCvs/FaK
MbjfrjTNW8/QMjo7vpogx3OP6Ah3aGA+iFUKL8mpaPdV76rSB5vAPsnMZ2v4YE5s
jPBKw+9iBAXO3CJgfgpcOuPvybd+HagnSazteZAuC3Ve9qyb4QNMy08aZWu/Uia2
Wm8vYDPIYThClisAvAf/iGTvcq+wwzkpUqyW2+BM5rAaMmrh211HLhi15eSv73Na
auSGXNusXP4R2+/pWfvEOOYQlGMAaOCsF0YkJQjJvns4vCZkA++Wkz191glGz6hs
R8xJZ9iXLXR7BPY3lhvnjPWs4fUHRllgdRACU8jbKKDrq1xahiSsjhw0KwI01Noj
u0h64I7wJvCJRLV997RvJ/vFKHHMLX0tqyS8hP8jUG/Fb2Np4zRjC5y0IZCHuDyz
EXh0nxkqOFdKHqhv0LQUGJ8aiEA2R0aI4ehySHLbxJS6D/YOpB7Nh5JZHe9ERy6t
kJg23BV3RlQpY9O62SsXeKwMjzRPnlQneNkuXzQb18FefDBmaxBdayACPR3ORPbv
ZhuTainzAuldeCenN8rw/af0InZz08k2R2W3T2Tr/Yl312jVw6k1jTvIJibbgjZV
Y4Ic5qBGo/lBrY6tgPwNKoVWSk7vXisEjT0DT/yneb0BhuVl1LP0TltDIZC5uphs
fXLlsUyAtmZ7nU2Nee86tWjDQrb2EHgC0dMWKSelYJlvtFqkutjKylTGV05d/xJ1
nxQiTCXIjLEteAKu77/W6vmm/uZ5RimORKdMamPPdX05KoBab/aFDk7zaruMbRhN
zhdN3EUgpAYpCEfV5QtxWh/+axumk0SmdWfbiw7Gwne8JXKG2xuwualwwV32cYJi
R/gWxRc2RzFF2P5Z+M2IvqxHIHUjmxCGhhL98bKdbObkAvQoGfBEzOEm6dzkeU4f
WXP27XpzXxW8JXNIZe9tqyZmU+erj8kZyhdJE45oDIu5K3E27/VYbuJRsAtA7b8N
VmVzLapiXl991IQ//4SzhCbNApKYbMts484OOrEob3mVtEks+0uOfd/aOuVwiyYZ
hF1hYRuQIt3EDufkx6QpudjCyZRu5hTCyeHZ7jz7xNliCwZx9rExVLvpgjyOg+qQ
3P8c6GfTPCjPDNtf/q1C08mm54XFaKsq34ZAFtpfcQ4ElTV0oQdMQOYdV6YPLi+l
74x+MRyItqWoujsZBujAi0Rxidqautu2zmbfVI5cBphni5EpTQ7qd5rLqxFQA0zs
YFdxLAdyazL3nldKeLETyZxuhPqgWAMI3AbbpEzsHQqP0d/lw2+Bgxckmf8fA61D
cDXORynMuMB4RC8lg30PgBB74DE6kxFjQMQr+7nDHslIMBuj2H1mj7Pc5nW4WhkC
XNejjL4rfCJGnWYIMEBRIpzbzHMN3oYTS+nPimxzXTys1Sz8OypIiW/FbLDTPKla
S2mfWla4q4MY/pFpGDN4konORK9FG9kTYIx7rX3ealkxmrZLPFoQzqgRgCOyEWO+
XX3yGIOe93kCOcqL7rpb5hMhMDwT4VckZBLv/ShLERzaAlFa2nQ8lxkSpnEldCd6
avTvbXmVtIOdL3JdRoJAdpjZcKGOd4b/rN1pmFMMff80hXmuXN9I95A27moaQjwe
GkmTUMY5wzS5wINgna+9hAcROoseXvsM5UO/E5rk/dQFT+ZVh4DVDmU4rmkkv1Im
mFmUU9RtLlgZomtOAxpXPANidIeY3l3ShGYJuVMaF/i8T9eKkVIL0foYkF3yiTC9
RfpRZQFxmTQ18KMYfaBXVa1KOMntR7KO8kNF9Jqih1ZlLDhvw7+TFwluyH1NdxVV
LEjN/c73AT2Po0/lS4rrD+ef67ECHntEDBHKErb0sGtFlVtXSu/F6MKEg9SHSWIZ
mZ1jBQx7Y32NiAEqFH3QdT0doFPHuLX+XrTj0hNTi5phCo6AKsHw0PPUHTXH73Tw
JFSbv+0sUuY33TVxEXQZBGleyHDo7TNks+Eki4E/ZxfGEqSofZyqpYb7cCNC+CW5
T5W12qAFD50g5suPmLxQWI+DMyPM4sLBWTKSvjW5oL8Tvn4z93I2Y3U6Or6HJ4+C
TImpeE6XQ9dpKo+fUkxFi2TIdjBYSz7+x7RhhVhW40y6MyxjeW8DgGtU6KqBxUB9
`protect END_PROTECTED
