`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDJF8OkMvQMxiJi1LQnY9oG8rBJ3TLUdQp32NN9TB1h/gNePDP+ozM8OdSPfidvy
+sM8jw6BNLcFXvj1XKKzZEAi4tZXYNQ9Tw1k+y0smbfgcUE1LH9L4mlMA4cLRKm3
8e4k3vVj0D1PsjBbBvUWRhawYVDEsihPC1ZNv5dYQ7Z1uR0n3JxC3OX+nMxggM8g
FiPdmlVzHVyhZB9OSp81nsLtdz4tyZUVzDCtWBG1FA5KIMuqWgDxdxxy5u15VUxK
fa7oi7o7eoce7MeT77XibKDflJT9zEuw/NgNopFjtUsTGEi0XquVVCm3uKCa1Y2i
EiJ8vMdK7HLPokPDIOWqdzclFNPUxKH1yK7gFdyvzY9W6pjS6ze0dhueYiiHYyct
5X2eGBSHCpOsokWHqLhsNmt48zW0PjH4O2phLQSMI+LBvXoxX8BsvBoxYn3q5bhL
LZcIiKbGpFI0Atzf4cS7AnVQX1WIDQCfldLnNc0g27CYDJ5yp9qhukzhCDL9P4Ke
txDz+o2r+qXqD7bCEMz49N0/IszhacMFzQ0tXUi1Jh4HmOOAvugCfYgv5J2cKxRS
4aJC+LL6p+qv59fkd2i+e0dmwZ4tGlpEOACmRuX+RKeYMpYvsd/9NWRQPtGctyl6
uECeHLz/JM/Hkc4GFk7dbuVns/jb3PqZp7tb+AIwRWAOb+wg1NcOuppaIGd7HBxq
kLJ6BLnpFH2/BbDba/PAwbTop5Q0S2qVpLYGcVVARBnPH23ffQwXRHxu4CDnBfrm
NBfoQ3C+Uybsy5YI2nhebMs0MotpPUpskOrIqLOLS5zKasetVLJxDa+AXfSxamU8
fy9KvHWq+7zweAO9kVIQpFoqtWJqa0j6P7h+/kvOnA9iMnx9CqvaE/8T/7SEwVvn
269ceP1jgEql1DuVthwR+BzABMvkv0NZsOm0DyFSDtCimwOHxfaqVtDffztoAsJe
9H5vcn23hTqzNNfwilze0HHzQIukU5Iw1vP/rykIBYYV6LtjY6z3jBo5SBd+jE0u
5zmbOzNAA+D5mYRXO54utqN7/5h4zEAkWWzLNKeD5PCppXJYuT3vgebHhgOP0fvC
zaiikNusgBKXXSYpCbge/MijJTo7AODmV8JWlpd8l4z4zE56cnubmRxLtySCInX5
AwsE2DPWuK/aKJyUaXhkFUqXBkZpsyvdj/4Iug9X3oFblTSeKlQJ2S4vwnl0XOaO
PqSpzeZVc+WMmLHxoXbcwZhkZd2ekPALjvejwaeLgu9ZOh74IctMl5T2k9jUDp96
tsGPNWKFX2xYBVauWvN0fBWSUYMmnqdNC4rvvnVDNs2Crl+x46vPcw2Nmy01ko/H
omYpVODN88ixKI92B8YtJLsR6WOEOdfU1AQsLIABbNmJdASCDynnLgJ1XWzeuuL4
jPhjyqwDa671h+3ibBVTCe+zcNI126FSK2YhugqsAygPFnHxYscyL8JJ4ehfHNbF
YrVj9XE8Mifmi77MJeOU8ANU+NiihK4mexmR8V8EAqr7BVJaNRo1g/VjQbdZwgLU
0fXh2/MOWgiYfAm2gutdeJ2GRIlLYUf9loruzsPCOTl14dsEm9/SmFlXhQorUpx/
bu9iGOXKcXZxFoi3qILZF7y9RXpktAISuoQ9kx9Bv4Oxn7fWejHHy1uepATvHPLT
e6U5/TN9bqARjMqIELmvCGuO94ieP6yS40BItAAg5aAJoWGU35t1aMEu1dFUvHFM
7wxvOBabVaae5Kn+OkWG2ipKkmxx8vnKg9tJsWSiQuonI7oHTIUtQXSwMOE0PKYn
tlflvFf7R3ptN5BZVqPCWaLaykyZobxbb5yfL6upW5ubMq5azQ44zn81BfoKM2Gr
+VpFQ5Pk2nW9qmRS53V+JF4nF60noAk0aWapikDiJDW8ycxmDg0UURoQZe8VxapS
IUtzZ/GS7zw5JlnukjacnbfXVLmBDmeh8y95tSNggzxrrTBYWXHwjjxEa9X9nNTR
JV2b8p9fo4+OAF7jm/OlCiT7krH1GgRnc4AbgFPBdetHeMXMpckDQQEfUk1RWFSi
tE/7fxqma9uR8xtIUcdFdGk6d4JUy5cWssx87C+LosK6y5srZvqx7Qc662gdbzdf
m7mktzAHiRcLkYQqCo0X9OYeZFrF+9yALIch1vucxX/lbbVyBL1OqfMtSbHbQMGt
ZoKbOp4BLFOP/bcychEzNwYq1jxigqvWADVR9pisOPpI+Oyc2GXMEFEONVAcoOa1
LSrdFTYKwIBDwB835St3+hRIcYafiLWWJM/uxVZccRNRJRVnJhyPAyFvOuSwedll
3+IB+jrkmEruq/MLf/2Q5+15872njmWr6QTIzXnpiFAO0FbdAmg7csvwYuBpxw98
uK0Mvm81NhDaRl/SFGhoDl/huA30DfNkj1VViybHZ34YWCDYBRJDWeNPPTHcIo+7
IUPG1JTsRRC5WGyLP9CD8EA/mzuyYsAg+BofEqY2S0620jrYmW6uO8ATNcFNDD2V
Pc70lNv5r/eEEqfG7AhTxX7gjPNWWvT5DvEhm2FOW0IdlkbaECn13j84XppeU2SC
VVxww98eRVitmopyhsh3l91uXtdq4Q/z4gsq6KKLbRJPwEjMlJKZLKh+01uHEtlB
bph25BglzTar65KekOZBu8oUHBVEMSjEFLldRZtjhFryh5D6okEfj0cD0g64spHw
yQ3/FpUhefVY3llF1WNokDQDjhq8aKNdm1DgfVqkmmeaUZYywNPYX8mzmhSCX3Pr
3CbI40SJkpYMdgIyZJ6E9StrobWZotRxTNcU4NvPIQ/hXVNUSaoda3kjKAVJNIYy
iDVdSVdQUzyJvoaCcw9ijfY42C64iKI1CH596zViD4ike/SaOObzDe7Ax18OVaQr
Uemc/eojLs/vI7mqUr/Pk9PQamx3Oy36W8UbuZcYpnzD35yx1M+3g7u6fLcLUfyB
2eJIpbayYfzMpdTRiJX93Ou7iL+cJXlFZnoKMigQQrD36dzsVNJ41U0z3FAk9jAb
jevPnb1TDEivAga+NxLfspAQJN1ddu0lxMNVERP48Vz3tZJD8FUN2Jkzdizv8Slc
wtz9anVBSIE3WMiIa9qK2wMnntC4B5YIsvHbAwEXvdVouEn/zaZyEi2qXQGL6MnN
CKgE64xRMXd0kAHfmuWcnO2Zkrpq5QqjNcg+7kExLdKd2e1SRX8R0a4m5R7OZBjE
Af19vUMbQLQgl9VTydsBVaMlcAWSoE37V/KSThZQZjDgtnswNBw2mOxfxh+PUDl5
VHTGY/zLIb2lRNo7P1gCw6/CnIsmdgBW8/EHjq5dDKRsUe7UzNJ6vnux+rMvgpv1
2031ME6ALft2tt9Gj3EWUG8shxu/XmGQLb5a3oSO7E5hS1Xa/0XuQ2buc8k5NM2j
J9gfQgBbQTq6brpiwoAs6Uj5DJ3Wh+3H3+PoSgT6TLnbPUa9LtDNkmFNv8GKhwNm
SC5r1IHpevC25YfiBjvjnDpWNuRF5VbL/1gMrtYY4KJaR/8jLHpuG7p0yw34FBDL
7sAMFaAfNecv7pgR40t/Tq3xkO9h667yp4+5j5qDe8kolAX5RwZT2Xk/CtZ3S4hE
0DFJLJTiG7IJ8RFk9y0IfY0voblEgZrgNZcPQVnTOEaylPUiX2XffhUPmrtsP76r
vgD0s9+4blGHjxy3oyZuyGjf2NPL1GIqRygL2woOPgdewFe6LIz2El00DZKOd87F
fRv8WAfb3o2/S4z3otJ1J4SFMFd2xMIgvDGh+bnPyAEg/NSKxew1MxP9eyf6oDxx
Epap27K11Man7h35qdCuphczWVtuf4NInr285N/BOhSjKDjb6hbWqjy2MRWlf/um
erd0kIzpaOLbBgIM0FGrmWB3trXa2LeX8ANMjAe0rAd+3UxHTYx5muApI4J8kpP9
2gXEqGbd2XUelPOz6gAlg7BCs4UQOwp0eHfeUQ5Pxdh6gHSNxJ4ncOzclQKI6vXy
s9nJyRBu4kMxaKxHu0hFif+4jAfyWakyAiDd/PfDd8SGsNgp74DLdXS/T6iAaUSL
OaRf1sq/JbBDCoo7BgchIUO7SRBcjDgfuEaamC8TiuTE7vW7CjZW+tIVtzl5y+La
uBwMpj6+CFTqiDM0B7jjase+cEDPO3vX1j/PEPf4CQFVUiq9Q/9GwlIKeQOQ+CXb
FBUtVefWeG1+72NanE0Ke/Vq2y2VLpvm48pPpcc2BCnwlE9zOeSRs7kM2bggmHcJ
PbgEPGuHhi7uE57hpdPBvxkTc2VBc14yLwGV7vkrJoseQ+D4KXDRVphyHGuve450
udx2Xr7byO18RykRxTfcXeH0oqfSOmXREKbf8+5J5Z7xL9jywsPGaPDd311nOmWW
98C91s93LKSGeRX2AxgX8wRHL7+gRzeEryjK2LWOTRbUzblOElw/cY6e6t1eYKDU
Gf6HwP8nZOK9us22+A4zcwUo3O3MQSTfhBaJxNSQe9UXqLeOd4o4SwhbR4a7poGJ
pSgzC/huYOVAbvDSnKTe1Qz99OVbyNfNpZDcgncjrnEZVdhsetMtUc9E5mPqZ229
E4em5JSKNFakaB3BQB+Jp2fE3/jjLoCFm6ja4xC+wr9/GINkZctLNSYg0GUcBqnd
pzyP/Ey0I5gWpIEDIiwZ1bB8VumhYVNOgc9MjMiC8eNs+TDWIDgL3WSC5ammNJaH
SqTW/LKznaSmr2RDcK6vtEe6BI2/sOIsaeuNgtZprwy6QzJbALpeR5L7rPeO0Roj
OyTKedBm5qBJaRCeD+khfX9bZm+wXBD/JIWb1KrcudUQCz3scpGeYtAdUeJwP1aC
Jt9LtuYw/RJenVb1+BrposbDZ7y6hzXQpQiVjgqWuB1hGFcZdlnastSGhbUrqbSr
nSkhyPtdTamjv0ofvrAdOpWzOazFLiNgKcU22A6ru7s8nZc2CNu7OcC23esyxBMM
TnZVuE896tRzearxo4ssUxz40BsNpkhlMtwf/MdphC4HCC0nldiX3tVnP7EX8cBQ
msGl5FDo4GWIoAi3U0Z4eV27eIvGjsjIoJRnzyFtZ2nxOO51evo605y8vjLgPKr3
a78FmDHjNVa6M5SzC4ekRJEkLF6nDJAMcRFevkpKjZpxJ8IajTPQDKkXv/EKlVw7
LSvhjWNMI7ZF4h04WRr9xjAOIuadoTmg6taVvvMdNqiIg50B+srJBICQG/cSMVdr
dijh3uvQKPd4EppdI+6AkBN8ft7p+s4YrChIWDyrRqLOdKjl5P36+X6lOQnwYdfW
03vQPpYygemsKhZABq0pzz7gQ3npdRgrM6HUGJs921p4frUN4t7BIIMDhqNHKLyy
NlnZ/mOtSGOhv1Nn6S0ma1xsdzJ7E3C851MxQAxlWuij1APMwHv8ExxQfGhhZqTU
0FCx8SlhTbDhrEElZUU/fYiKLTzzRpNy+f9J7UBWPFu9b/wuFH+hiBPAuQ/gIF84
Ej38PAnrWYurFtrVJHjg1lYQFcsG3/pbjOZhTQSPnBv/TFfSwBujtaaqTuzUj8Bp
SmshoM2pnT5KpzoQqtq9YVQsLOxo6cc9G/KRrG25eGQk9KErWeS9T+YRCDW6x0m2
/Ym3+8Z8MwphURW9BOaeNBD3aHgpVMSOtjfQ9Qs7Sqk69Jb2ZZE4BYGmw/Ma7Wnz
5xY3xmux7Lw781TFGC23xmk1wO7pgpLzrRp+EhopTcQadZ8kcBiVFf1T3ju8ZOc2
G4WThi5pDOFnQLGNvaEji/Pnv5Ey8gRFVupqN+rjIhMDVy4AkmxOGPQiHFJ93U42
56RbPGRyaae14JqUCpIBXDDCtgF1J6ZJzf5toWV65IKigkysjc7E7w0ebI6RhSPZ
4iCCSGG5gfkzwh3uDldBrVngOY+gGSXob7NctQMMLvzC6cKzQinhVPvkiZa4q2xO
Od6Zky+rCeKodhelF+sQfA==
`protect END_PROTECTED
