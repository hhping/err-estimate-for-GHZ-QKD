`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eOXYdON5ckF8AHiPVAoUOy7pyuClhQrqqx4FsST0C73T8bIbxYNRSkOTzKV6Ic2
Vy9koDak6vXUhv6xJEj/klbsKVeWeThWA14lBB1z9yMIRvnlRfV+li3RBBjz/Jtt
JSXVrYvHAG5wuaT5cV+Y5R9A3SwjSkTUKaVXuCeH8HkUbjvt2NfK6F4NRuty0ZSc
9c1T1MPvoWbtz+LsXVrHm8V96dTKkJ/HpbSbKW8JvcGSN5MlNdJClptNxSJPphBG
k0Se450kDe27fRFPLLDb5Jym568+08mrAPewDIrFmUuaxyAdaC1SQ+pmjfLrqAQS
S/gVu2fKupq9eYhF5aUEeKGu7DL+wRdwlDoBdgQOccWBuQDCjuhhxPwjZlvmy+5s
MJzgpN9cMLfU5/ttG9JWl4ay6rZruE350kaXDNpuZUHi9VV7HxfHJ4k1ZeKXQcGd
ZvbllKPAy9N/MeBU60rSJKJoGSr9jAJdh0MhhOeQZk9tGIa6+IEzBFXU/tmSjRrU
unOjQCziVMlaEb5SaKuBHHwwSwwZfzMAB6ByDXMJYfNiUKyCqP6UdthJ8dUz+nhe
gIWU8IQOGMQsqGca9K9Lef6Onie693HbcAAPxIVBpZjQcHNeWZ5nbYpoAiHOXgg9
YjaaFPyQbsIJBHB2klKaIbszvYUoaNWhaWOuBk+vTMwc4hJxMToSYnIVzmM5Er8u
LuOCm4ftt7lqRYkeoVh9OF6jzW7Tj3yjl0juNeglncevTIaVt8gx1QkrRE1J3rtr
/oZaFRL898d10V6PzyZKYCaBAq9figKsHSC9bMkrm5rLO9b2GVZG3a7m6f6GOWeV
MTcDZfn94N0uTQg15XhdKIV9nkNbQZ/1b6DXe1H8UAmoZa3BW40pjOBdP+2BBVUB
lehHbZh2oC/bF2s3pcL3ofo81SGrpQL/uSW/rMyxXWwtso7PALJAz7FOtCZOkM5R
wppyP5RmeZY1nvj+LMZg+w==
`protect END_PROTECTED
