`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PAzZgLLHRMW9LDXVWTf9RJSNHGlGjrJRKUl9HZsvZydI7oawN2eq38nqGtbkSZ+
AMHpp2mgWuqZMv1q0L0VWrJOYTEsChWpB1wdvyobZbzvKDwMayqPZWCT6Q+fXNTf
V9txW/Eps9+wSmN1LzAYMZZIcjK+VHJ0nA1qYcj6Hs8NXxTQNgxOZTeeye/Pv+Lg
FSJJkSS2hCWYMn+UGWLtrp8AuGoDwKXtfW2SSJ6UCuJ01revcg1h+8XoWDo67UfA
IUDE8jChw4GyzR9HKkkoRhCNMEA6YmO2YXvtvqRZrCoPoWp8B252sJlB27QzpvAG
3OF+jylotLUBcmy9LxCalHJDZ6Nl3YiFthXlGHIs0l6IykZiDoSpdnFA2DeBrj9W
yuecQchUvVG9r8C/ufCRNTEYujPfDnfmRvr4wNuzL3cW6CwjEGWmRdiV5JDBf0Yf
`protect END_PROTECTED
