`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOQ2bqvZ6LhDpEfXWTdMt7g3km0Jct3qABQRc/Lj/nStxW6ZyXYy5rOvQNt3Kd37
A2uYLz4eUby4zzYpQO9U5OgGgvMHPTKPfG0FECJdnPvEckPDEKEMzeG3h67TEa1G
4QfFuV//O4nlYRjy5OST0yR44c+DhfElk+sQ3XUPaN7K8WLjHsOLx3dGUXecMyoy
RkRqLpaG9UEwRLlHx0F2J2yNWCVGxNII/EIYoA59h3dlP1XKnKxDDf4K0vsxOimW
4iq3dF03zWSQuXZkHBtsZpNV5HaNlI3iW1/OdxaveVRllqS72Dbbis0IN9XsqDXk
dwz1r+Q94o+hr4keaueBAbVgmA34/U3bKbZEcyutIswK9mF3sB+qSOdSVg7M3Ae5
MenKtmO68VUSu2FBddFX60lPmaESNYK4J6wHIc4RP/WLxbiTwC/l3hX6asRUfN6i
rRDrafM4FdlvrTwNmXzKIjANTHUsUTeAI1whrFJVMqd2DYi0H7U+57h34fp+/JH4
U7mLKeoao9SbteZbLjMbGO9PZ46FIIzuQ2LUI4IixRQii4wIGOVrQVBd5BaOxu/h
gevkdzr2SJKbCW1MxoJtmEVonr7O31Y57kgEv4JH9t0cwZD3A3ISUP1FY87oI3lt
w2v1yYR9Gfu4WJKu97rCFOED+f3G2F8u8nXFAglMPmhtTGL7OfpJVHmGsMw1ZNmM
5u3TjHjP0v8sYjYMy2kgKUw/odsknbk1J6VNupLVX051HxGPl3U6Sro+VivtwDgv
XjJGvc3UK/2YIh+y1vYhZqp/KrYOme4qLcG4fGprjFNuI4mJKBZ43gBdF2MFdO8y
vUwkeb2RMe/vCjBl11omLvJ36pXNC1yGwwS05CPztPgG/lIMnywudD/k15tGxwKH
9QGuEte++M7e7lBLy1rbiqP8XagFHjUZ2iVD2sey+T0St6IuvqKYnXZSk32mNci4
ssqK4nOdHCAh2zygYqwbmAtWiyRSchO6e7TnIip6R2+DheTDH6EYAbdBmJ77DxBy
mmdXFOCYEC7CkdniL9SrEs7zXQS5vuHMF9QHiVnjs9A7Cw9O/V1T65f53odjxgSZ
Lft1iPsFNg3ebE30I2aGZ7r0cw3MSHUqlxVJmh50t8FcUn3nf9+qkZSuSMVmf7hF
1U2OGvoq5gf83WdoxOk2Xiy1pXV/81leDyLT6T/Ql5eAonvXY5TVC8BjEcKlcNJA
xfe0s8MB0CncFz0NulTylR6dd8MNIz6Ji8+g5LGkZAriRxJ0SbjrjYt1MuT0VItc
g2rx9Om4ymBcEouWPLOscdiYpxEmHnvf7S1R8fE53aeY2B3MwUOplbamvJ2boZ9o
EGGWytbNIb6ctOv0kuOLTKzb8H1EnS1u4dSEXJIjNvpcanVoAPgSwVIi1ZP+PmwN
Q4WdDE5nDyXFkQc56T9C7R+Res9yT+8++X9z6d4rJPlvT4nQ+wNV8hmUZ3uz5R5o
UfuAm/bUOQpjoB6v+AamtY15Ql3pS7ZFTQYgolG4a/zXV3n5OMELcxf8lIO72UUo
t/QQ1m8fz1CGxlgLm8rbOXLNEqtvumhmB5FItEBhSP+tYEKmQZkXCK3k4ZpT1MS9
YAOUmk/wqleqZ5zDSg4cIqQ+wG42El9lJ+FAghFAMCZ7ZtrZj5FTGsdqoJ5k70IC
XZFri7u2eMfJCcSBEYNG71TXOfqXJEgAsBxIh8jxrigGo8ZNyaeXt3R+R+veYiYt
x1DkS+lvpim5sccR5D45w35aBAuO02lr3yOnC262BxNW8dakFqWD6RWZKN+erFwX
nMf9Unv6jPWCuduRIU6xjsEuqaK5Nt7ez2lVly+aC0WZZKqy5HLzXgeslpYLSNAm
dH2QYEJXXYo14qyyk79DGbl+vwBFLBNs/msaeGUWPQ5k11tlUJtiu3I2V0yUHQ0Q
7yzDFqU5UJt6hNWGW2IeQklAjPCVhfCoXqC8l1cXO5wYFpocGTR9lcWVsdAdHEOW
fT1j5mSwjKE1OhxpnjbeIu5LO7vsmzRS/QZjRP9xZgvqMx6vDNBgO0uKhAZmupKu
HHSACUvPfzYpIIgUSjiz7aq9ZJ1zIYGLoqX1v0Xvf3QYsuOSsSY59aLmrbB57m5Z
GeIM9Lu4bh4EbVd+Wr+YxLNAoMsXgCa9Nt7//zhEhhL6X3Gsk0FZKjE4hO21IjLK
l4MWruATFzKWaxhDqd1BTji2gylpyr6bai+d24iPUPeoBT8TcP0xsHL532eojdaf
xqIOCbBrTqZPiXTdYXlYPg/Tio+Hy+VlY1GolSJliBOI9QEujjQKe51QOLXYJ0z4
M+mdkb/BMgSNIL+leYv0Rt3CU3Yz64wIkkJPyt+4H5WTo0fnS0GZdWe2sdqrYgve
f49QuyLFBerORKETxrPzL0KCmBAMII1D9Ukggiz0UmdOCd8x/WYpY/chBHu/HV38
3Qglr5KGLo7pPdFeRDw9oFkbywtf/3RfK0uUL2sLqC7QWVgwrYHZ2tp9PsCPkWfZ
wI3kXmTp6/xSGnP/llvLrmn2642COkupxQoJd91U+HstgN5N7swUlJ0S68P05XXd
SxGoO1PAYbeFm6Oip1nybJR4qTKtdSFIQKG9m6bDJpPmPLjr+qCADKmuDwhttDPq
rZwh6RyRBelGs4x7hntyOpR/w+/j2KSZAIv48kPYaWT+sd2CaMuDiwPajiVZkUxF
6p4jtrrRKxNr0MfCKfPSrqRqum2F2adcjZKrSr/n2cmcOiAxFvbnlTKQ54n9rXLT
5mV40TIEibApMgD4I6/rjpqLsXMwepT4qfwW/hmocH0=
`protect END_PROTECTED
