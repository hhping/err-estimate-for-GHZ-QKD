`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
seGAoxfdl30cxyHuSbjgRYSAp84TGD2MumE3Qz1c5VIELOLfeQppCmE+VeBjjFg/
YyU9J4u29OHeeMI4dIlSifQNEOFUuuBh7ijbBuyfyEODRJM5br94u0RJTKTcAf7B
ap9Ph4EY2E4fL0ghWCMcLXGTvSu1q+XWu9a0VkOJislOd7Fi6iY0sSoWrwNDWqkQ
TOk08U36biJaQNuzMDABNYs115fsfwlCai5UqA3r/mB98iTSVJX8ITmuLXNCILLo
+WjmDKK0H5iQDi/2ZEthi/+/ATWZ+7UwvILcOGAq4JTybmqnQ7ryBzQwExbczRkY
drqeVgl3PHW72m+f1Tam9LvVbYpsCME6mNV5F2MGAC01UDdkXjPY2fWX+rqTKnJq
92QBC3mWkg3V2lEPIbpO9YvDiCXffzIgATcahuVuqX/nmD/J1PLiGpv4LLnVBaCW
HSHG/XGRzE2K6tLBzKSWTJjbFShE3P8HIF6DgGzIRG87W6xEp2jQaFhIUVB25m8j
eZcQpFGQmUoCTHpJm/vSv7KYy+dLEwPMNbtQRko3o/1FH2mhHh/iUhkAYCz7HCwo
`protect END_PROTECTED
