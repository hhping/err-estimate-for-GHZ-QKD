`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhNsyB2+QLe6ZTrOWeD0pVfzbuaiE0kmvE3GJPG4AAKuotXnZv/gdQDXuPeFqBNi
jqnMLAtxYok1D2nRCJe33YuSwzpJsVSwRqMFO7YzFnY9rMoWuLy1bp7w9NAT+Enw
+8FT8Fcv2W+BnOBZ3zgGR4KNN9h5Kak1XXuk+g4BoRSgNetnk5TNiLylzPVe+1C0
I4Lo1uU6I/cSLs/6NZPRoEfuImm9Fo31w59g1fVtH95d1Gme3PKMz/Hq5U8+U4rB
XbjOFx1oga1GDOF9NHhSvVTBWFMdD68uzOoi3/xRKqS4rHXXdSfawICYzVEO380C
fL/gECYJfiUKERLRRvjjDYuZsFgB6SpgAPToQRF5H524ed5ygBwIHB4Jg4t9cs27
ryFn1oB9M0NP947jt/6nYjdTj/2f8SvpUK+5C89YlSzub4CiDz5ujG0rXECvSvjJ
1dcAnj0V7zqZ77gJaxrEr6jdnhhFn3SJm1rm8VzbqyyplblaChz/mK2CrK/KMrwi
f8RJLCN/4lt7nTO8ulhfA2bfbzm7n6qdER+a5owAgFXCY573F3tlYmyuuqGgQhOm
IPkVR/xIqEUGKJfi2FEDqsimUMzM0SKDwtkiICbgEbh6KdzvXucjclgbh7fOm62L
JHBKsKZzFD9lOmaaXul2YXO9DNkCql8P7AuzZv15vL93uYYX3UsgeTcbvC6LPI1p
OC9XyiSl1lyshhYgy82nU7iyzKXgjWi9wUDZrjy5XP6utDMzJm/PqBibLS8aFk9K
svD+71QX1Fo3RVjcCw5jH7cL+JH51i+gzDmt86rz+R7YT/iHP1oElD/qr5aBjTGr
w1MvoSc2jd+XOf4p0wKzN0aXAIzaD+jG/DbZwAlbIDGFsN+/rlRjXXj5uQkArhLR
OLdQiWyhSLdtkPIt75b9QaS7KOIjC1jZB5JS7Mdp4ynCWTTrYtJ0H2qBcUzJl5DO
L7nEvzyYIQasrbbzHmT32lro6bJZpsfgXy527w1i+VSLc4SMkKvJdKZyy4ziCfGV
I9NXc8bsIOpTSM7NDxRv/PHjwnlkExie8FY6Jff/Bewi99KwV2i//ZVAV6n5qGcd
7FhAmpGLJUae6BUfdAofJ1n83gP+bkEKts7b0kz/8/UOUearZ7JUI/coXPbxWmbp
KJ1m/IYxdVcQSy24uAdl6pr/zlTHawkZReQLqCABRKyWV5k4yNQ3xryiA2JVDdPW
4nUHF9dRJivHTbDxtKL3sg7KdIpu1wKE8BiuanccU7AlJp+W6cgeUVf+ZsAytUoi
S9Ikai43NFtJJyexXmQTf1ujb5Z2xNMfYx2NiInLBGFhe24owwTCGSjzxdn52N0e
OdXI3en3cC3CCyiDhq2NhwTMErLpbrTdpMb08XeQTZODZlU8s6Buo73RJTBHhIXZ
1KAsRx69st7mMu5+M7Fs6FzD8eCH9HEQacyN8zxYIfZ8B7Og3IsR59A7qurqjlSk
ykA1imD9V7tXn354DKTN/SghquVzTXqN5avhQBvrOvq+TMjM/ybPuk1jY41NjU/K
eeKPhJej+iF1xgmvdSC9lO0Xnnj1iNeROXn18tFhoXOtUsE8YLpHxciLUsdXkQCj
r6P2Aua6MlV7f5eZJ7Jqs09VTRmYm8ELOjgA2aJyG0qELu/1oyX+UOGnBOs1fH3+
RoQvCjTTEhleolOYHFb6T1jrMqhoCq07MAZVdzAmIP9xytbz99/Pc9pyV20kXxNN
xLUXLIQ5XZ920ox752vmo8JbWJf9ZcQUYOXH2JMkGV8QHy8Jb1Q1So6RNJMsy6LT
gEFMMJ8s/EdpNVp+QB9x275h0ZFKV4N+jioGkKhgbFn8K27B+FwuQFiNhszaJsg0
6pWHaMIlnsuDtSLZDB1qcoKn/cz6D13mMGds6WmSMuiovNXGrgd6+oaiv34iAVWf
TLDzJ7zpVgrfW8CG+kgIWKGKrKC4iXHy7dHpOn1ps3g=
`protect END_PROTECTED
