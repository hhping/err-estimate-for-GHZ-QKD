`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iN3fTe+FiLRwEzDDGxmbGxudHT+D9Tkw26eGuQNC+DcBqiG/cU/G9W6Ap35BNm6p
6ndVssm3iqsPJQu/jtv45f97vijbqO6V6bE+P5v7cvDfkjr1V23NP9uhqTOyJqHx
Ky6GjOpC3YU0jdrMHQv8aT2e2xFdLZcDhSFoIFMEUWDxkjsLGOSYbzbuv40Guz+4
10gJi+DaN06Sg0zu+e5ujS4PrxcYA2bll4rKYTWhaRi5RSY/J5c7F5JJJyTMeoYP
Jfn+NMDEXEsVMsP0yTORpMxgIFvEISuUHSgObocH/WeXys919MoCTeA0An6KOVqQ
kMT5ZrYapbS019v9Ym52wY89iuNAMHMV4UF5zeAmDt/AgwTRkS7+2t41nfTNuk6O
Qfna6QKbbKF8OR/4ZycaSKEXULFvBPCJliTc+RdyAphcWmZIiQh6IQvmC2F5AaqD
vpS1Z/wPh/nWYzg8VaJkdtTfJD2Fy/ppMsIXyuOSAv65dS3pOSwE2WW6Mk+C6TpM
0ZzjI+IIBKgk8pV8mjDGpW5Nvbd+//9sIcdMKygiNzy0q2GKWGVN5NJkvMuQRQGk
PwaHRfKzS1Vo6Zp6bDJGUwwhN2rFti84bBLg3gJS1uY0kH44UJqCIrZ/HKGWqn1M
RZ8oum2mzcQV3Ulk11kKmGHV2mfeymwvfU2kaVJHhvrw5wF5LTg5vSbfl0sfRuub
MsPlE70oJvwowQi72MNasg3XORVvfAS7/QMFN7L89ZFvjNSfPtl0TrOkJFzuMHPI
ONIdZzME0PK6zDO9CJ2fpYjvnX70p1MY097gFES+n1Pncd2fUTtXOLUoW8/DqHNt
jZmXCPssIFX5LqQapj21sfgOCyWc1bhyzb4xz0cHs5aiibbciLhDhOb5MVm+GYUC
LZYsc72jAgJ0Dl+LSwMF9P6IwyEUnT4zhPSNlEmdxDcWFuvIboBYO3y31qOlMlu3
1ZksXxwMwEQdIocBuYzhpaPApaan7schmWKNmA1Q2CN6bsDXwF4mgvl4KH0FKVuh
qDCWxijmPyyw3zlixWxjQvTe1osjXScaufHKmPBE0PKjmnvdOokIZbj2WhS9RfR7
mI0F5Q5AJ3+BHj5wKawROTcmInZIK6vl4cHdbXeLb0WI7w1UhYNldxh6vaMy5fSd
FCz/nAsJPvW8Z018W6fsa+1VTlfWOkxHhzQ8/Lv+qQqbY9oBtEPD9BVVU+1C4Dof
Xd8J01QM8+Po62bXEtfV4nQoHB9y3R5bTjAEGQjJj6nC9/hdy2LCXn1dIkitqMzf
HeOhTN/tIFmr760k83zyvNZECoOPJ2jXTKt28cWXFVo=
`protect END_PROTECTED
