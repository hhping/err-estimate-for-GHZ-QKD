`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ENIhD21VzlVoMMJl2eNN9oYbrDsTlxU2XAlpo8yJSgcvX0BnrwU8QV5KVTDYwjAj
X6f78wGUI2i7Ymd7JJBp77Jd4jEVUEvq1t/TR2Q5GB/A068qyUI7gaexelVxKBti
6oYsbwl4FuwjFdnmxYIvi/t25j2XX7agboUzPKvQHCJJdgcoFKdWQQrRf6mIwGeF
BwoN128nxxV1K4We7hPtIlkB15gocZL1S8mGlORJywd4PI9cuZX/b3Ho8MCZ5VN3
MdpNLcWN6i5RenUND3T/IohtIm0nQBj8cXUfZ3tXX9aZyiX2x6g1yaoEYnl0S7PZ
M9USFD1MCc0ceus3CUm6GmrZ3s7sWXcqYa3kqUBDjMIDvBIX0x8rMazLoqws1nOE
QMDbdsK/eDk1wuhi+TDn61cL1wTAwzwmnE7+G8x1f3k7WLByON60Ikq+yNcknS+n
aCGNqEgGC8FY2s1NeW36KU6qulomDApN020biFYlDfpeGKDG12/tslbQCWRRcx3s
vPdSPFI/tCQc7g6q3CiQ75hfG7yZ3mxuxpdEf4CVZ1i/XPFE27us2TOd+ODuWj34
lsMM1cL0c7ArQ+D6LlCUr8XGtGduYV/JmKtm/1Zc/6Grg7WSRS55dsiqJGv2Obr3
6A/TnyBe0cr7SxMQ7n+RpqIaUTbv61t5l88dxggzl7mlia2C1tSA/3cF9tlVLKDU
BOPJy8bMBQ0gFimB/0g5rwIDp23QZv8h8jGEuh7/tpLm2cPtJOK/qwDl81ebaC5U
ZiIsxdUPe81caZy5zolrmlg1evaxvCBQrz5FLdhws7rxtYGur0Jvitr0u9NQzNav
Cgey3DdWgZnMSiE56qvuRuALLc/vUIlQ7YpGqM0xt1eMx9nT60AelK3FnkV3UcsI
MZOhi2vNL4pvMIRQ83nyQR5HWPWfKvLp9FgsVe71t3Y8eIkWfhLtClQ+b6pcUDSm
7H9sccjZEMI11/XGTvY0wlTbNbBaR7XgIvWZh3YU/Q+tS2oe3+PBI5oHUcVGYz8u
zmFYpU678QnYt+FKUYxgV7F1uIuzYHwADH5QwGuT0SV8EofsMN+Rs2SUQhZ2cYFJ
oT8c01GmQgUd6dMlbjpZksRihaH4fPOeNegFBnRlXxwUQU3eMn0rREfmOnfX4HB+
pAnre1ixaBN0GhZHWLfcmNM95F0yTlfOeDF2raKPof0=
`protect END_PROTECTED
