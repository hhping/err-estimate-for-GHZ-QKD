`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDOfWh6HkIIYp0tf0dBDOj5ktB8JVGn3NCbqoYF04KvQk4Oq23+7OfO7Hc5sfkEg
ICZWm2U8gd072JWA9xeJ5rdbKDHcJgLiA5Yh8VtCloBVakwVK7rv7y51zz13xb3S
Ivmk0/wgLp4tRAIsuJbXueemN+gecCZFbdWNtELq3UJiBLj75NdN2pUyIgaS88E7
3jdM3ufNROUChscpEeFcuOqJWZTaR40VUn8eKeFdZbs=
`protect END_PROTECTED
