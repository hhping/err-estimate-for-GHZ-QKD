`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYGxbNvENpQm61xvqhnuEPeVvwdZnXhPXTd1czDGZKC5/ERzhpGZmwOgHB5g78Pb
X8JPlge6d16iOYLCzKYD30AZbeRi59lOANRqU9wFDiYKlgyUBU0CDjAwUg3pS321
9iirSNeDh7SvT3ePIrqbfcQ55uURhYuvTMLmfO/iVdwKLF/963f893uL20lIV7Yq
FbE8zZMwssfKmHfyrfAae5cVxC7UEgwPT1tkYk6HIQ0qwLe3iGh0G+ilzTazb6Yk
HqO9aPX6ewzc8igmax4gUvfV8R/Z26WUnDIPGWuFrNZEql3Nmfk/ahIYwk17xF/n
zTg6j9xed5c34hfPoub5C3n+AJs5RYnZBc9NGflQYKWosBrFuIVXBDJMbt7hHUGA
6lnNMvu0/RACxz+z0othuDi5nEpuQxqJTZKQTzLv2+rMqXQFBw0xRGkVTOiOPicv
RbwXk1wx8kkrzlDJ08/Zfaa67NqzHlIqFHN7mam1C8vc1aN3ZNYjmNz5rjekoZrk
9ZK8lY0nEPVtLjRYinQLvbxbgWYdlm5+oIyHiUuoa6xNjxOxOEp3RkoWqcBy9O1u
axeY4AkvopJfw1uiieRtuyC+ygDajBQdg3NIZE6xWwfESwTYO/iaBAW4QC61YBsl
Kgq1rrjeklpn4ocv0ivx+A==
`protect END_PROTECTED
