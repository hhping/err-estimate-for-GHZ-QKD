`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWLJIV2khtzRz233svcdHOXg0+WlSavIA99Abez7kETgEgvITtn9W2rGrErTLRV7
B8k89QW6PFLy/10XDTTUA/X+JKc2GnomQVyPzyRzdorDww8xqSikYimEMR2JgjD4
tmarrg3SoUHNyO4evB4qHjnZ1rew/EVE3rwcPCGYkcpUBRU6v9BgyFegybIxHt2M
76HWV8Py8YnFxRY14v0IrxS3SVctuoraSvqd1hnsLerVT+J5FxQrsQhDKZD+ZCuK
tuK5hOoflIWi78C8AU1Qt8T2OmETuUzwLGMOIrIcZcsDQ3pBaseqhrHE7zjHDruJ
uvSWbeN8E6GmHy2gwvHJuXPZozm7Ej5PsHSWhlgTQWfIvTMOi/rTs1BZpBsbR/kN
PFYnytWVsokgCqkKtOapE0EnVZ4TP0G0G1wliwPQYHOtVNkPSYiVVa783LEBpBKR
HGSGB2RQpizlpIj6PcHij96RhdULpGiTrzdTMcuIlhk9tsauFCG/7/phxAA2ChiJ
MzALmYmZtQ4VgRrbYt8r1yzYZ64L4u7EGws0llDk7OZHKygsmydJImqTtXaygwcc
N0Hgrt0O/TcUFifz4899r5+gt/EN3H8baUVR2Yo8QaWbSWD4ZUx/Ve2GAm/vKcSH
jZ150O7bey4gAn9VZXqItZyZ0RVDOYS+1rk1doB8wUfYL8myOcB81cJ6U0H/UizA
/ojSV75zckNSW7OBvmFiN4i6Tp+fCTspVAUlc+zVjP3/G2V6adBm1eAiDupxqqRP
GKM4cnpe6mq5olMm1UDvEfWQkcIHrK26YbDYQRXhuaV0SQyR74FOY28T2kgtpMz1
28S/0Ahf2iURM5r59tQYWz2cdJ1lohS3+4oRz6EX5RyNcaytQria6aOo4DtJ86c2
4CM6z3yAqopM8ESqzP8qQeof/3ankEUuDJuIA3tsE4pF5widjZoNG3IDYdiFnCAR
nr6Z6dfvWIsXhEa44pXic8Y/PLmTl8ou1dRTgtbXOEuCGzbw+ioEcTbLDQqLxe6d
X+2Y5BUMXJQPognZ+e7XuCnlBiQuyd29phoOxdTtAUUtwth6AI9yNNzU/WrV36YJ
OE80HEHCg0IBSnqchKI6luw4C4RhzETqqHCPjOn0+izt42tXeqy6+XbaUpNqLzR0
DzZKHRwcQdVV8e/no2NiDVljyRem03OdFvOZ+ZFsXEgEH9WbXNYhJPm1QBT2WF6w
pjwICad+rrgH7YWOrbpGZEFf1c95p/aOGNHNiI72jqW+R6ZRvA9lCtrpkia/FPO3
rUPQROh8Xho6DDhcSX6TPsDlK2gPYqX23MOgRxwYFvqbE7Tnm6Ilm7VqxA/pW7UY
1B7M3RrL2skNJa3AMWLsqSPDd+WJ+xah7FKpB1ci7xfjtKwcFNzpi1UolJcWEo0z
rXsOV6dCcFSfzh2EMVMMCsmCNKTpD+8HfPJP1SZpkIAHTJYUdMVbE8WiV5nMoWls
8/x28WU4N7c2VrrATbMCDg7ceu22xOzTRXe2ZixWwshp/hPL8/JUEZywaI7Nx+/O
/v+hJFpysSil0B8mIAsmZTbYyTWrVn12mSLHTURVb5u8f2XV1WBGysCxRPhY9ySF
sSbTEZE/mwklJjQpNGh1WfSjhDaPFy5jZEa2AkkSQ+P7PlbX8hDBpmJGAzDQCz97
F9zEjGEthIQFqxDGWRBlZhmJ1ejVNdUPP21z5kzILXI=
`protect END_PROTECTED
