`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mZeWS3dTAGth/ETtv2jY1ulKENLFARJClK+iBtIcbXo19ugdzwZHKZRFU34LPeb
A2GAHxNx6ahMiLTX67CgnQ/YTkkrenbunYBtrtRTNap4EJI3Sb//5MDcisRAEAKd
Uup7az5OiffdJIoyEtwIkdTITRh+/LL4fXfNofQ4o09NOrA/xEnVF1wZJCkBGgY5
Hj/XjVeRLdAusLkBqHvm5aOYZfB7arQWilA2Q01V4R/fUk1XaIxc+Vz9tE3Eyuuv
rCRWGibYryBWKRnW6evB+S/bFeHjbgwaMWJ14ifyRaAXyHfefWU39/tSg/lkeevu
DFyG25Jze92UqGpRlt6Kpu6jYX4JmD2D+R08leSTsy+WBgrfFVv24kLhccaU6BdF
U5JDZiaAmc2dafLi+ZVARG42SH2aaO13mXvLcZ8G8w2sxt0vupeQakpXldbQia06
WgcZiAp9KKKQZdwGEHCcFLQe+gjSvTUg/+cvY24doNfLUbdXEuYC3XSZpCe06cry
3JBxccx3Y8hZprrZ6fphq8F6hKTdqE5BHa1bP9JlL4rgg3joFmCrAtF1s69iSJPf
o9ZEwkHgNgYHu5cuU3ptI7TuMwhwdR3YzDAkXCgJ9ODipVYaCVVhf/Wd1j7QHVda
CButIKCaKuE+QSe0hxu9ic+PbmgE1B0g1hI5NakkqRefTBp96qPirwvtNjypC5JZ
0c3qappUtgnu6fePpgX3GnRY/tNKuYGcmnQi6OdBOv0UJOuTsVlRIVBevAz5oHrf
uKnz3cJh9OgY7RVdATFeXg+Vm4tozCnm1DDf7VvLto2FYrhOum/v6tfr0sSiUKs2
OJwGnC/+XPDlVT+tGbuvU2brt34DPWAQcKxNqI+9sLb8PCH6j0Ybd7/97kC3nRdi
9uwxdJLzYdRsp1R8yin8pQkzTNN3qSvXfKtLjG4GRLKka6BzukNQogdbQuyw4pMu
tYgM6umNti4gLnbN5br/AwkIH1nwhjNYVqMm8bKr1eLfVEZT+Tbo2rWUI0C9av/p
bWinQcX715nXyYi6imuh+PZLlXJwxcKJGDJ2FiO+a3oBA3cDTPwQWy+1gWOxnE+T
F/ZkkLid7BjAEEWGcTraGQDcvrHohMokQC44+x4IvhFhp95hSHlflyoKg6RzRqUe
xzYlBGou6mCAE/nHJZuZubHVS9IN4oUb9DR/9IopOK4P5EOn+iSdVqHHPcIWXo/i
RmfRIAgmSd9YzvkS13ogb//cX+70BDltBg1b+zCOlGh+iispQOkgyqGnLEbRGPZp
+SMb0vWrKL0qVJqeukFqhw==
`protect END_PROTECTED
