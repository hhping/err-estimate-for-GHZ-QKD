`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gBy5EIBJw8RC9soKL0nP359qbPKraoG95B/41lEysV+45TRVPEyWvkbrpLjwSiP9
XjuCMAq7yUasoaJmljHPUGf628UcvnTjIQ5p7gD16tubDXeCzJmA/G1LFqhCTMWp
TWivFyK8KkOhu6GNgsWXGvLxYWiwUYjy4PCyyTnzHMNfV9JSKwg1rpfARCKEwNZj
MIqXwHDBd78mhlgVZquPxWbFJO+PWNNdOEBto7lr1IdYW0zBBdJOQfrA0DIc2tB+
ySFQjA9ZYKk2Naeuxxm42v2cK93xyYu2URtEDlDFD5yTRlZzfPtKyBhOcLxEmq1R
XuBKfv1T1wnGlHK7gHSjGpOoyiWAQVXLuqPBbC0BzfQuXC7hyhBY+BNUUkHVynDZ
pS9jJGbOGtlbiLLld5KkYORweTVqiSCdGNkmCrALhh9TvlNTOva3CVm5cPG6/kXZ
zaSvNjhnk3Qr9VGaf6JV+UbBQ9YScs4R3k++IIlBdcL+v3bzGvNABvRd3YRSHUR8
vBqWPK/mVx/6ysHiVkDu87e1fl+xhYg3G7FD6Rvlykb5kEx/9zXdQgxbQezEbHyx
INxnjQf8qytPwdu/iBT1dDVerqTm5b9i/FZUrqDCKELtQmksh55KcsiIX/ZarwRR
y2ReQa2jyLfm1vJtubUzjS8WvVaUCVeydz+G2jqEmMuv/YhToCaBsNLDzFPk3HFN
3cZC3mJx5Bg4i4uGve0WtPwpgJnVM9nhbpDMrCUTsessOaw/KCyPTLDVzOA16oY/
`protect END_PROTECTED
