`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4404A/37lb26/bb2YrI0MI/ZUolLZ1Xuco8FkJngD5pHiixltzIj1yWRO37rfYcl
B3/29sdeqFVisuw1hycMIrjBmc3gPlDVUcIpvbiY7HoxNfbLra1jIoXzyPmsq80v
K8a5yOk9VOymhFu9PrWjYMhLCTgkOnUESgrf8y5DTfX6xeyFhaFNaOT/k0cV66u3
kxLrnEn/KsFJgssPV5BiPeKKAQDDk+y9tZT4KZSvhX+cIztN3qd9NYIF5v6SDPaz
XWAGWYnb9IT4YCH39cTQMNgX0HoyyGCMpHHPeF4Io+fWoL+2DTDwRujnHupnftIL
/flqk8TfXMZ8FXXS5i7xvqz/dxRfLxOyMKEJ2DooWQkFQmAF28JZU5TUxnSmWsw6
sXOOpamUuxoxeVU+T5S11aeJay45ZY3sQnEn4HJD0CCwPZaswH6u06ze2M/AzkEH
CbJ3JII2s3RnVRoSWdMLlSn3exTWrI3a5ylKCf2MIf1hClmngTklAq/LPuclfZIl
OsIzdU2mrDuvqiw1lA6npea3mfZSLv8os9+RWPZC3SMR//GAal7wCnSWYziQSVm/
d3gxO08xC59YvAc38dWarr6HwRDKlMG1l3jASYRIfoeXkSwjAgNUuxpuIpfU+f7F
0vX2vidjx6N5l/wOs8Q9mPrrrMXwZix4wVwNGbJ4/GjNV/7viQaauBCjP+slcq/F
9sOQR/pUQgkzdgKdr42Vre/EIW5zsuq70/CsgXaYBuovxs0qeXqYJjlyRo9eBXE7
lE5szskm5TQkaym9n/nT/HFCN1QZoNQ6Hcm6MHwyeLm+kx5IlXwFIU5MRPfxZYop
DZcoPYvRDXmYSCozXlRZEpega7LX/Pi2eIL+OkU9EmFNmYmbkEA0ur8c3E98mGLz
5UKj7yVwstQgEtM52t73/G4VklczFKyOfoTMmIYLRauqNQVXw4hMSQNOpeWkv8je
8yW5EqrUvVk3iyO1X+CMOXHTqxRVp/02Ux7nbXbqm13GvUoczf8F+VteJgRgDHEl
6bRUVi+VwPyrLxOnZ1DNUAwoWmAncxrgCsVcw5XRf5lf3z9LqqfdZZhpgXAlkKLs
yEn+/KZzdNq1Hf8RKdaVg99qqU8kCo+vm5c75YUAFJ7HjlmHzWhGBk+M2kkcm8Np
vTBvx3bLUsVzcqj/l3wpUyLAjTdC2zKFqWOJZz0cCeeHqZF3/vM71L6wMqhZrW6n
ZbeE+oGTP2U7yhXuXmbVtb0kjhdtCl40Ipisyl9Cp6WJbEuDIYZ4V3ooVkktRtUE
dWe0LXQNq+fkW9wifbNERgzHdgbzVxcbN6C+7Sj93i8DAzR1KxngSn+ck+4W1Mj2
/xZx0twdSPqAXqsoHzXxSjF84wMHK8yUmH1tAdwPNltsDhui/j0GZ1xMktYrPxPP
oe8pOdVSV3b5DY404+ZRp4BgpLQYKR0gtRZXv/4ph1SIWjyFVX2/drufsynOJKlN
62d0lER+8DC6A6AgL2+R2E+ZbmipbEFBJPcy9x3T5lC+/J1kwfHjeaTtgbXHGQZ9
mT0gFCkRx6HQXL9Ij0Y8q67iyLQr7m8H8OKaLjfDvToqDtaHqTwLpLX1rx8y5n4F
xri4nRgqkKA8/1wE0mWj4iii6vutOjDllXEEq6CCM71xVcWxkIJlm0P3WiUEEFdW
49V7Igp13BqvDYoK6Bzsc3y+/xcREmV7uvLZ2m3Z44CLLDszBn1oz4jbJ3CR/6Kt
7YFyEIqJws5CXFSd1efYIWMmq5zEaldtpDVpZacq979uy4HvAsKsLIPwIRCx5/3m
AY/diltJWYrJaEScsEh7OlH4wk1C2/UIHchG9siu/8udh8aCV6w28Oa/w00qvL7r
CkCkH2ADIz6dx9LMCDeuBhbgHktX7POhEnjTOO3fEFYL62Ncd5+WgGZkFd/ZQp+G
lJwdOsnujocmRwpiGua8Bu/lcObshzPQVrcdgzna1gLaiGsGagIvPNvQuoeQEsqg
b0pojX16ZuAqgcBqJ+NJgL1oS9GDHw1/F/VMxV/LbIRc/EiqyVqLqdr/RcDh5pJo
+AptNoBtcx/+713dy/2bLyK5OexbeUuGPiJ12jQU10nqL4WslhJC5vwwr8CM7U+P
U6ryjV4Gfvz9ozb7tLob8gFnQ/E639LoqXS/2HPQLEL6eIz7WCIAw0FpouIi1fRH
jULalTAbSnzKBpcEdNIZWf2K7T5gZZRQQ8GtdZ00VhnwiO2ZJFqLrshpg4pIzJPV
H/B2GBw347dEgkUJ/b0mVWb33maTDYWIuw+WbX5iz72KBjO64XtzBYElCytP4Z1z
x2Uv5OHr8InTHGTVb+Ugf1V8ztFw8oAvu+wcJpSUG9oucwKyV33T6s0Atzxhfv6O
IX2H9bvRkt/0W1gCGhdKxTahZGqvqe2Y8DhIUlfSGPSB+tA7pHdBr9Br2YyiwzIb
VZqDBj24heIvE6U5rYkXJsarowPuKpJWW9MEiuxKRSANy4T1Vsqjy8oCsJt+5pLa
yRejiK3r2kd/wGL10IVBf3bS7WHZ7ugt2QGkxNxKQWsOsfx++V2w09uaicSGM2Cx
eDxsurNCnKbNxi4+LJJEsOPolKnfWHc0nhhjiC875jk3oejF6tYGx5iSdtrR0X/3
9fhuk/mFCUKyEhNc9G2fcDLHUX524eiHHFHPoQIR3JqslUOy/hBulS65f8nyJbIh
FR/BPTqjJW9FjTpGkgPvrDAf24BQMKyj6OJUsre+QgPJzAwRmJoHRsBRFifflnJD
X8NQRufdbtWYCPJ0HJavfEF/8GFCym65qJ4NHNvKru01LJ4eTulRKN//ZJ7Qu0ob
VDsA0Vnwjal8EwmRPyZ12oRSJr8W6re5+JMnR3GJrOicRGvz8Z49SWyjgNujXwGP
MLffJcmC+UFfXCBl3e8oPUIlhrLn5DWBgDQ9+cy3WlvyIlVR/1Cb9fcngX8WWhW2
j/KAykb+XkbUHOjLDeKJO9gn9Lb5ZWdSUf+rksRaLUMGGMlWDRKti+stCbuU0r0d
4G1mR39JJGT3Bj2uZ4ee6Yrv2IPUTwziIds7AGtIPLPGyltygXMkp2IvSHXf/KOm
/vqZZ/LT92VBVh7g3XXwqINU1qAFAiU13PvreNkJrD3PMgEie4uPjobvLVmSxekf
bN5jUfnK5c/u39Ilh3NyyhFwrHJfgmNn7FSXDM8Xpzyr1NP/xpIXjj1oEScn69BV
uJf2Dtr6LdT9p4MigPtOznYsTrPmeL0eI1Ar9+ujzjtn5BlU3Cs2+aKeJFYhi4d8
qg0dBpmXBV2mhyWJLM/5HfVYi4mQSA/tDDA+2KzDxKhaEv8NTdOrICDHrEv0qH9m
gP7pIrWWQWTQ9OOVRfkEoLfdkU6V/Tx5LenncNizp7TDbJQDMd5AnlaN6r9u0pi6
8Upw+1TyWRBdUlmoRl5+j5r5ByYX+RTJVXgEHVd867o2+vSGKzpt0UFp4HU5D99z
p9XtE5qA9gzdxSGXemD9Ncyy1vXfH57jmMPP9RdSNYCyDIkWWzosB+UW48izElih
Jomybd2dYQDQ0Vuc1jzz6SUBo7PYzBahili/YTlJ6/KfyafKtBUFgzNdxzf2UKd+
M4J1EqxTzzWsndrs1Dld0oKHemo+f6Ne0/W7X98ihHK8t5CbJ1VbTCMDB+arlAY4
8/f+6kFbl7uQNW32nw1Y4pAv+pMR/OpUsfOzpv8k9kbrC+/O0FDZhndGZjRL7bsV
Rc9ksOmmAlZkpvvOuM7VDMyjD5rpDYR5UfoATh2+B4W2xvidyQ8/QaIQ7QhFfIGJ
uX0Ha7U8jMZ6Yz9et8B/JtVkAjj1RLkUFTas02lF9nMklUW3qWGkHuqcn/ey0XRz
UnusLQjkMaXdQ998Wxfe9QoKTsQSgZ+FPKaUQ3DVH4E7hIRdEDxERKALxLq8guYS
/43AXRC1U59GihRSGol/YFf9HLAdV2tZ1AoVkXah5uigZ4XRRIP03jSJzpBpy/Wj
j9ksm5RLvNF9FaPydbTMyTTK6b14KslXDO7TjCKbYDMp61VZqu6iV+LcwgryxKXg
frjx5MiLwLM5ixOQK3R3GrvaSuWN70xveBHWrWfUZrQ2EfI+0x0mg516bKJX4QJL
KPo8icECZSxtdNvgcS10/yPgq/zkfZmnKA3l5mc//q717+m+wJQC3YRrJ57FpXVz
caV/0tzdsaBujnAtuKt+rFrNH7zg2gr7GRreribP1jwPlqHg2xxopZ545nvr5R19
3au8dFMHV3zPypDEoGYNyokU3fKKhfrL2V3exucuyIV8AgQwhJxgSf8bucOIC1Im
nu0jy9r3/sbY8sGxfGpiT0twKaO1mezkzkOfFyLcTgfZ8LXE8LPnlMe+dLGs55b6
o7e1kf9ZZ5FhTT7OeW28FlVAJTcLpjjMZ6O57R8VEkjM1lLOXcYvk52B/RZvkERx
ZPmDko9GCWjb0gWU6o60S91Qm7PFJDrijas6qmnlTEcg4wvRJvIarD4BZnPIeDww
yGikm5BEGL8e0GzbgfCqmoBA933FnHu44wwbgRbgIkmck6S3d4qsvwKV+F7KFf1q
PFEyduy7aMlDVOvw4aF42bgPIsOOceF4nNbTOA6czBcTYW2LF3+lvU3ul/5bJFL1
YO2t6s5VUGGFFH1nBKG25/2PndIvl4CIJMg0XKHTEJ4ebZ+ZP+lm+wjITljzBMNt
RvP+NjE7KjJT3WhY+xQ+WyJ+Xun51ibja66MlEVXajCj3GE1jNWKEsRoV+0HJ+gV
j9nyxzcTRdVXQz4hiG17/kYiBF+4FvqpPMAF7W99KNoKIPpvHLORpi43rwmZNIaQ
i9LR9aQW0woyf6csyVf+1O1UdUHyStZZjRjNxWVTMsgI4x0aE5VoIIHrfso3pk6b
mIW/UWxboyWkjbPpgAztWkRLpFoZRpM/Y9ltKHUKgXSEQHT0bpfDMk/4oZyelTnW
uBUymDmpA3MtYs8mmoM+bQ1ywDqiF2yzgwm1K2QlN2pwdKaWq5k5TA9KEXWqYXF6
p9Uu4akywWBrLu/6M45U6CJ1tQKorSXLTaRf1W+Jr8gIuxQb7Y8lxNYf35QY2wIt
mEUTFAP1mYvKhjK7htYSWQebbqd84G7iFD4LrGCXcENy88leco+1yyfJZV3M6q1h
m+Hyxm1YJ6vBuuYgGtJnN5nJmHFt7vk2Go4H8D4kZpfXWXHJq3GXjxcBEDisxTxz
GHBTwUZXx+QOaqn47FdqEEs2iWAcl4uuSpJV1iy1ipeoKCKSnWfNCVRyqHyLyTBB
9bx8m1hMtRbYMKUp09sg9knMZod5b2/KAat3U7euO32oysGJl80N/8Bz/tZr09G7
wv1pndIZW6edRqP1bctb07sdtQdTGtI9ZY/OrUqGa6WHojysk12f3Ai3vvlrjeNF
UCehI0IV2uLaFIPOv8I+xSwvGDHcZAvH5uS1yoLCFUkvrUYMMQaDUr4VTFTGucBq
guB+wRUSgkO1n94dFqb/N+cs0TZDs5EfJjh2Kvrog0oWi9JKRGkjdlicL/P6S3fl
cUY6snqR2Mk3qrXg2H8/gT1lSaBm4OJ/zmcEhUh24fg7Fc1BECdTcolV+Pcv2ELE
1qlvL11326aKKCI4z36thef3tWTLNhn1/uXvrIjPCHgMTriWdNa7bOLJwLLlU15Y
Hvd/zEMddl5/8aajXvtxA6oUZJrOSNBvSZHZQs8marI8iKbXKRJhKyOhwaJkCKrL
jybd3KyzPhw/yPV5l8Ym0R5+sHyaDil+lO0ULwwC9EwEYAmWDmRMBolEM9TtOemm
Rtya5/kD8r6J0W4fznQJaldqa14oil5DGLqWxU0kQjcJ/IfcPnAvaA9a7rVljJyW
mVLB+STDgi8PoMgTasAMEuudielVSarHVkLPwv2EgaBWR8cIIPTGDIIwWoWIRNtv
Vcfi/FmV8lAjmQIpNWKvi+vy3607w0v4y83lvYCIgbMdXKt6SOwPUlXme5oQfx63
eImMCLPA8R5zgdQe3cdapDrdiWzRYSMr1niBl559Lc3UFxVGtFZzuNr6kq5WMHqq
2Xtydu15ML9vdC7tOatgXXSKLwPkuU7HIc+ePuUUSTd8yCBwzv2eUTdQfosJjg0l
ZGBHfmaL58KulpviWYMn+AflL21VDENOtMH05r1Z8EZRVsrUHhaEXI4QkOpc1ZzO
RrRy+plrNzaB6MYwym3ZNU6ET8EaSD2u1iiImB69e6NiJtr9jVHnwjhR84OLWSn7
yomUps39mzm1t+GF/2A8NMZRq43lN00fpIYfdrx3In+vefYQLKv4xjh2PweALKWl
UxqAVWHKDghWDTiqx4b4po3oQknUTiLSl4zuujQa2eSON3vPaZ8jWIP1sFGy6qvn
rXIoDhoaBEmboDrMlkpJ7TmSysYJ5JraYVhAmYOj2KnHUoRvbGAgLautkN2e/kh8
kfoyowPbwAtfA2zvwg7xJ95q0dhsYZGolZH4UY1gZYH8tPv5E/T1Ak6SyTnMK/vb
fQrwn82axTBzm4Rk+xvCtVOCUutVLXFhRmpq5pm4/d/XqwD6yAo01OsVJuGXRBof
yhRpSlfQy+VRk70LXiXiQCUmL+HdaCBLi6MiMQhSGPel8YBc3nFlH6N3B8k/mq9s
LYdv8aO1EgiqoF/tyYVhclnVHUWAttAuej4jCSbbYYemEwA+KQIZFHwBrkS3fdU4
ybfTt0Ib+0QywYEF6kke8X7NGjg6MULsyZOhPRnCcjb1jyJVMzCUB30FAL4QlhJY
eoUZ22KqizDvbyFtIrJlOvn41Chmu4pqDPbMrtTLkOmd5G30FMf+C2I4pIUNFRZj
dIN4JYBreOv99qu9K48UKeWzNeid/T5gOhSOhEAjFPbaRVO6OSyyp7dBtJFh6wPO
zoa5uibdjbgjHCSlaLrveqC1cg1Orbn7DLi9egQVAziLSTRMVYdb4aQSys71bzwB
PCBsUCJ7STG+eMjM9AjqH4Qwh3b9iuiVQHeUr2EgX24n7HccyivXovgr0lsZ0vKr
CvoaZYefKamfgn3oR3u8mtJfoqA9m8v5aBWyvdaG2tdDP3UjwHRsBNX/maF7cw/B
d+81iRszn4dMiHli5bZNlFi460puqbLtAgn2kY4a8+COOzA29wJtwb55j8dRiE2q
HeBMoaBppi1o3PFY4anoz9Y35RNPrnwBQZzh2klzxoSZ6LiGcBYcdh66pYxNs7x/
JtHM7+XBvXN26lFyAWOfL5YurIjQpSttgY1AFbCEcEzxfrxcZD1Yd2zyXVWyqYRV
Bleu4UaM7nS0GgJfSmK6l/6WQd74iQY3yoZu8NA27+lbkEb/SvIRWm7IGtCOvfTd
sjgpD7wrdniV5M0vU4iCO406mcfsw9tMf0KbCLfiZAZcHxUEmYUVkICTEM1hB3gd
6MQ/jrMWJzhun+Wi2Tbqi1z0cpwrDpa/kRPDloKkwzhd7gH0ejVvrH1sHsvR7dD5
PZCXY0pIlnFKve7dvjN7TP7lm1GM+JKwjWk6NtLusk89yVJklLi4X/4h23LQ9dhG
wKN/0IitvfGI+dvtS8etHNmOU7z/lEJ5atKMa2ax+D5uIYrH5cMtFyxpmJ2Ladpn
iDajQES0VLa65v3DViNAGfcdqjv4vPFgxfcgCS+hhZ6N7doQwoCflMxSFFASOa3D
BLcTHpKWMh2CwfghSsVQzaSyQjkKMwm/2hd6onVSmQsijzHW06PWId3y3He1ggH8
Qo/40FD8cbIq1fSCZ/7tib6da6j+zXLn6x8B6B1VRxHOA8jTuku2h6VnNqXMSYb5
qYXIbU0ZvIVSENpU3VD4SUapSIHeciCxa9r9k25pHB+gAh4NsQpSaqFZ4WeoP01m
esXe4ilyWcA4QJN7uIx62P6fRP8dc/NqSz+sZq4Sma+XqPKIJBTJf8me1wsT3L+V
4BjyCe+I/gTokMhX1h19JqDGcnzZQghZ3tw5dfqiwCDJusFUDwub7MoMrRAbMmi5
ZJNjo82Yk2wcw1SdUjJCzs0oJPOeypwT3hExMdatSfBE1kKBaFzcT/jJmRCge5JN
Tyx4QJ7u5D9tMZdRWwSvklAh7E0x4vJIv4fWAMkPKjTWP8gXoLDXeycKVCcQ2EwZ
Bc3axLISEZXKqt/gRC19MoVVapRPJyYk0gPYcx8YQstWjyuvMnQgkueDGMmLrGCG
auZX6tCg6lCP9zrIZ7b3osIrmPz8lSChmakDP6eJyJti0FPSjy9KthCB3zokC7B+
5RAOQSKHOaBLMwHWzVEUPP3Ycxz107j00TfllmpnpKY/QnOnjp2fRAND5dZV1zuf
NfnkgSVCbXOOUTz6oTR0fow8GTOOk8rl/R7ffu6EPP7yuiueWGQxmkoT7DSy0ohd
ot3HTvczMUKeqlKqbmnrH/DaCBDK9+zupZ7A6H/HOORfhOyuG0T+Lk22PorqaW6+
qA6B1mXqDvlMg9WyfdDUy6gaFeoQmxvlUabhnEC1BQO9pVpBcP0qYhtB+yW6/Nka
cw/No0MS8tZGXNE16bLSOVQ5MrXo8xLvoJ/eNq+jhVjMNMkOgVQvk5+3f06WsSZx
XAuwVXw6tWHVlXI8tpATrWPbxoZHU/poTHP29kbCia/aanxr7HZgpNNBGhJHdaq4
My1qbsVZV1EpRD9tFHNKNg4Rzk5ZMtxLu28OpN3smHCVbvWwgd5rJ2abcI2WrDlE
qDdGFzuW4Z/GuoQmwf/KvTcGzuRSLLdIzCF6ttA9VwA/QyazIrYSHcamTOnbwPED
gIMQqT+GGK1XUWypTjcdoPPzq0vrqfiIn85o8opjt4LrMnSYwAgXILurrCuoiNVY
9YJ42fXIy8rF7MIX37akeCfhSJBxobxeA+Wt1ujiVNkxQiHJIiS9tYdUgCbRPh/D
7tX1ZPVeXWRqbQFnrt7EGhHzOuP7llWKUIT6IfJgHMvA9empzw7W+3/Homx9OFjo
NG5SaCYqUVkmrY2+FqpjRmoRjUserdxrkKscW4lV+PSqz8b9Xjte36wCI3fSa/lA
WhPD+LmEf+B+2+ohSqjPB0fDX723Vh+dXxYGWpnYGIiSwpGeX2GUwTI9UTdT9eJi
RYhn8kzgoucRP1eDfvcPepKSdP7+T8GGgCQPlX3iwpqHV17n7PiJbB++r5BiNMMt
p4dEpmYFP+FACUv8j4RrRFTYUnH+e7RrrcbC3HV4jgTdKWC9nOyBkjmecHZ8sE4n
wUmMmT1PTamvshpcCv/72XzWY7qnhp67AXt7lBuLILxLap8jE246YFDHsvonKf2O
sLYLnNo9/YHAz2JBG46ln3FLXtUwKvRMtPwArIOzg0BU4ATFta+/gcFsQ6h7AWXx
Sckhg4q9VPPKVhurDE4IicqWRFOhXpxdbKnLJfzBD9JodmfHdK+Y4AMoN0gk934q
i6v0Biex2lo5InYEYbYZbRwqej370wfc69YmGFBM51CL919pxrilMuqgbwdM+t7U
O6VUCvxXB7lEGIP91ZEAidsIAc8bLiVYJ8YKGsFaArp2jylJqaUR/zZk6Tt1FkXi
QdktRC3tSfsobvrMKKFQUGvE9j8o+uulEgZsc10VU1u9iafjozW2kI3KammH3vK+
XDdt2amDdmzwXFHqSqFSqAWSnDuBZgHvymTVVhV9cOrr9yC3HwQtDisBGnerwFQN
UKgsEPVETdBibr/zAWnKbhUtnsR7zpgzpW//doBXVrGErkvkjeb5JeZ76QDSJtMr
rEjhtJoIw3AMVI5PVBtDevd7QN/VvLrU1iPyhF4L5Nx7RnUwPF85OgMoUVTpJ0Pu
rxUez0jyB5E1jQoUI0M9LfYjawppmPOFzkbSwFQJ1ubqHEqH21JprW8REo+iqUC7
emv7kFF7jDtD4ak3MiaagvTOqNsApPf9y8GISS6GTwCbGVI4uYv0Gs/4yNNg2y2L
M/BynNkLnfX4EZhLc/KgeG/UEGBa/nH7eETjUpTqfFPHpkf+ZGtQCkjOwa6DHLZ9
uMshfntXjSQ9rq0R22y4IW6cl/XRkKCQZgdFC0zCqj+f3S7H2MtFR5E+PlP8sThf
EIrJwSxMs934Hqjy2VBQUP+Pb1Ojf6PIzknAcK8jRcAM5fcOEivOT8j7Kl6kHa98
dlv21UJNSpF/8MwNp8iMeDeogQcI/DZ8RAuPnBu/GCGbupq0oduRCNzY+J4XRSno
J17gikXGgPuHc8JeIzKcB6/ZbvSXx6YqeVhWGjabKrf2DTgRNPy64HeRn2bYZEFw
+fqpmYjSfw6bfY5VyVy4hhkMJ/SlwTb1LvI8QqqXMogVi8kOYLaQEB2EsonMPRT9
fMRIqoQBHOZhL7GLw4V9+P2JcjDN3IwRAgWqcBryAskL4Wd2tmzpNPLQemXGjDmO
2YH/mi4ybJZlAILfLg5xZEk24GyfjnwIBnjLc6WZ0aTc7H9xh2OXUDIzS/hnRbkZ
vkOk2Dv/lqgYedoTOMA3pUy+9FpTYhSd35lTBh2PK0mwh1PnryxuEFDpbJ80LdoH
fm7mg9TW428tyoyUm5u7wYfv13e6olsHurzSl2XxysP1G/R4hq6a8h5NA01MNaU+
s2RkRlBXf5DQXBm3QGm7BExCYc0F4eLWw1K5MCgac375+495YAfbJLrPTz8yCJED
xDEQnVViFUDV5uLgemVBl+4u9BFrlMC118TpLdRmcPCKEdMRhpZGccCIhx6bSoK6
Ygybu52er4JOAYL7Shnt1bfTNcQem9hxbohsYjnRFTwutDB8guhSU6JHZqjz/kqD
zc9YuKdMrYfVa9IJ9OYR+jGGjIgaVOpysytmoJ/K7nT8GfuDpPFKjTd5Jhp6KhFa
Xju/UWMk7IrL3zsck1mFtuDW7Yfy9loY0+UWMEzYqzQ+ZlviSv1WjTjQhKU9tYlO
Y0EudXghcTxhoKjiVXDhAaLdigu9NdRHwTRVGnjBzTtrbShntfIis1qf9JudXqOl
sRBN1mmci0PN2K64Vj9SYQjq7/e0p94cZN0uk/l9q4v9bjOqYI3CuUIFsZmytz3m
Z0zeAx4lsdIN0lTA4RcoJ8g+AVyFK3eRwYdptWzfIXjNDwwiS0bHXbNgpVWgMKLr
BlFxANs+x5DdJX7QW8JsIchoNKG2OKeykFMuA6qVfwejsdQG+vLCStOKxhTs6TZS
G6S1rOZhFlTD8WSqKAf54tUkJctdK4shyYRKTHgLirHpwLKubxwVxptOgjA3e0cJ
0qHft0EwuH5GHujL1RiNYrEp6N/kjC2OBY4gNB4Wm48ns6TStv264/H2b5EgmRKn
ymxfgWyulHSHFZlSaH4rjtvD0T2I/Hi+q5Yqcj69bdj1JOhgquBSvMsh+WTFuLrS
Yxy5lu7dKnjIIZ2+7pJR6VoWmPbgPfjY3dQjrkOIxn+TJBJeXqYZK7VcRAtKYOeH
zJzX8jF4r3hBKT/5RVHvNhz+WOiXsooH3lvY9Tvyx+ULi5MgUJK5k4tcOxQd5bMM
dXTxSgjL4GUEyRU2wFYRGKLadQ8cbCv/vmJsO1pF6YR6S3CIbptKU/zN4u0DgEYy
3g606vcpwqqt+ihKCF91SO6P5s9sApnUfuOuhe/oSEYyqEx76tx/jQnWQZfaRSdY
M9cV8JZtRPXIy7nKvUXl6MCb5sUjksbBSWQHUPxedjhthmSd6YPKLMPQB8fCq5SD
4KoJN/2UG1SyQya43F7OAkEG3KbqXNjhMRDlXwL1LKLhzRR6plli3nF/7CZfeolH
IZNCa/qpuoNHW+8t4/GetZ+dlE4iBx5I1P3LBn0BhSv3fFtstEV+silfXfVpqPg+
s01qkuoYVfXxJNfmZEZzTGzht+FgZu5g7r7qgF2g3XuEBt5PQjxcXTUFcn/yE17n
6MQWAN+N4Vxif5aOiPh1jfBuvloBxu0mNdK9ZdJ/af4uZ29NIT7XqaoaEx5CJXAn
oUhIAIvJQdPV92OSjF1QKRiCU62aHGyj+qJ51jU1tWkJPivv1QwpDiX5d04ZnXpE
kAn3dPvdC21tSXh3epLUFPooPjUykVBn1LxyKpzfvZQEtq+Vy83Qf2ePw4kkbA9z
TFpANoogF1DmbhvMUi6qj4vUnzI85Yg6Q5L2t65RddsET+N+lvIt+cF8xErmkUbL
kcCBpJbXhIS10ORwGcBK2Z9iOnKOrKke9IxiSUf6r10x90oZbI68t6Jqf5NVe7H6
IcLyKRm3BCkl0k5K6CRU2efj6i2XSEU8qS6Pd8Uxk3WM6EGa9d0aZDdXV0wNa2Yp
xUBjWlYVQBBFFwRnDmFwQjn1Dh8+ti1hY9RrDViRo9mJ9mHtQs9KW+ow4tsl3dNo
U+hx9M5tL7kBBnE9J7x07CoA9bYGB0JxStIhKiBP1sFONCkTBIDeUFleaFlyvW/p
rDbEE1xQyAGyh1kpCKUsVnoJyW8RwMmCaorD3MxPs2T9/SMOYZzv7ZV2Nufw0FNj
WYKUTT8+LhOe8y3+abWPBo8BK4tyEmwsXAxD1ZU61n6qva0V9o3Ze0RAZscZClor
inNFAj1t+pttqZxs5xF6dAuH4j2RJ0LqglwBGS+Yue3WeHaVOs2XhWbfBRiwzW1J
BUUSyISj3zPqCqwLWEC6faxdumocfjuEwEKLi5mAdOv2IMn2T2DqlJThmwJ4tigO
ovcz08Fk7MMZSigUUHObXLx0L3D23qj4sHNlTnmrL3aurhA/KZlYD1d60IL2YCgi
pElv3Owe4bAZ/hHBK+c6/gQcY40qHHEt9kiEHojFKa3d8KQG+AHrKs3IgpPzCgNZ
qsjThanlHURsFp7ohSaE+6gqzPDPK5kwEWmFVF3oeALrVf71ugoGkno8JPohMXTo
DXKsma5SzIoDIAd/wdIYNMqtp/GSTJf40qFy9/ARQ7qx4LcgdXzEBfO2fyIwqTwD
IWFyy/iPEAIOGPDduCWgYF4xM5efuuGeDwNjLVseE8hO6E6a4bk3TR578ThRvNcv
gMAUc6QsQC+8RQd6RuqYPBVFb2i8wG4c9ozUSJ3DGPZfRvX0WtcNRczCVKHUZSce
Dl41sDUSm1ahcCRe27AAPesW8h6Db1O/n6Glao7SvHChMmHmIIzLWBddKknth8dT
Hp1q8SOzyi73EbYdj1kTYogePXqPZ4rdahztlqGG/a36cRktZW6i6rOchZ2RcIkA
Xx/cFU6gfjjy0EczEL2rX8up9HBvr6+456DFjqIt7KGGVR7TnVVRxm1nuYJ/KwRI
APH+LUCU8Mq/Hh3BAFcnUL6CDUDoB9kOAYUS+PR57yk3oYOPfAAwiv9Lrb/L7Utd
aJOPx7F3JnpkKFJFdz9k+o4MaPfXY/US+SQXv2GWMR/11c2cRW6ogCmIYBjc/V5L
uOIojhiUVabydy8zJWzyn8B393/nftEoccEj8znU6/npHThJb8GS8nGk2ZiNTAUY
pV6EiLV5K7AfLIra0mzkPnTkskoeTuhb74aXMPrP9HUuSwwjXEq68SXZKob4z12s
w3idGTpHWutmo2jwTIUuaNMhI05ImTe0KHmVyVduwrW2Nyhb9Xn0edPbAjIy+5UZ
iHUazfAk5Y7T+h4NpPd2Vpx/4L9e+M5mYCoA3oV5SgrNTynGhqxWwZ2FLbqbeKIx
IHb9TmzHuFnLCzK6CoCawXpNv1ng2ejCo7vqUViw46WJLA+0l43JLXm3lU3Y1aOB
xm3ocRyXyfzPU889CNwyzXjM3MhoHf4X/ivmZUtHsqO9D9q+17f6Ex2I5HEItxCb
QAeZI7tZhPa+LVvYdMXVBbciNzqSiC+Qj+y/7K6EWmFzY1NXSVxU2JIJFdUCHm0u
QO+SADF1ykCUWEvxQJwggNgbsv/xOXZgNzJPUiatSM3T5Z6fsgJ5wDSXm+CoHB6R
fjikECmqHm/eIQK+VOJ3f2WpLcF3U7QtWP2vbtsffvP64P6g5vDD70d0/++2Y4Au
C8LsbEGzJPtfn94G9jEP4DGO2NWDp6W4xSl5sdlh6OLsck8GSjevJjB8ljBhyRzr
pTxNJCPhRpdRBRxAD1eGVHQjpf3uVcuCsRtkvy3eDNcvPvd4F6iD5BCj+GQSbPEJ
2rS+XPIGm7BSl6ZPfHR8hrUXKZkGAki4QClJXAcRVIKSDlPCyGBDXgJWoYgVcZZU
p7VOjhfTGiyc0TTO7UFb38LoFl2yoFBgJy1yvv00XoJS3lqx51+/QfGb9edfQlBl
pgzFSu8fT+DlhKE0KJ4bT12MA/ym5rIVRxNHDLj4mqA7hnwbbNCe5DPTRxg+JsR5
xQSt41paGl38KPVgAJ+dwpKi6QlEEHjWmIeVuIi2d6TBQnyjlCIrqY7C80UXi8l9
30poj6rKxI6EbH8PleQNptqsR1n/KHSifBtjx+RwMqJImfS++mzfGGAUxgLOG9E8
iZRf0e7Q6Ge1xgQc2JgQtOJyPxfObfKGlrrba3T/TUo2rGB3Q1zsnWvsFGipVC1x
iVCra5vcjzyl76xE6xfeiaAWlZvVKuZ5em0er3TZBm3LneuLrn9PwFslOWiUEupA
5gpmGV7VbBXc+Obz8DJkKCX8yJ+uFYNSRUQyQHNsmd0Tn9T68YKoUXP++fvUt7zG
omLo/ZKZ59eAku66ryZBWC1fp9oCfmGtGxTfR8x6ebj4v7gLbnOJwjVDchu8rXbj
0DqomE76dkMD9vgFNV+qYQyz68s3a2NC/4nz0nwwtg30gluVhIZd6ZGMU4zvL+mV
iYYhCpip7Xzp8Ki79X9+8HrbjC5c7zYd581SIbPk4ZyUI/Rw7ExLwn71F2dE5FTf
A3SCoSN8JcMFdXH1GsKmwf4LhyYsQ1pSQotd4/QI40r0Q+LfqJXsFr/Fo9B4/ac9
xWTgS9cvWWgdsylT7jz3C/8R/jKWA1W9DevdvPhRqQ247yO4J0Pw9XN8TdnZkBkw
e169QNmvN2gZObzWMSP07Q5Mx1LqRob74mvqxfuiifMZxMoTMRfs2xyyd7JkDGKY
zwcV33tfNyVlwbUjCA7IoYSDZDKgqc0PCKhqxG7BRYp7MBuEriEIbCmBLBGTJowT
nwOf4deGTNJOxqtVXtuimfdJv2PaG9uMoDdPBSVOIjgk9S5J77df9ccyyhASr+lH
6/CJTlskV4Bi8sr2lZI6K4MUgys38ZBbqE7I3NlBPo8uWM2Bm59x+CLOHR2FBLmz
KG0elYm3OkE+PMu7j8FxGzYMmzbOA1WCP3O+jDxW1EgqNurOrG4gUufCT+l8YEn0
ZYaqZiFsrz26k/KNGl1fX2gmyEL4jHspTsag+3UeFxpevcME+ASP5/hQ+uCa3QrW
7wfrn9OrYCea9wDbukzQPChZz7SHcFxk+sSKIj+LskmijOHQlfdUrLX4+Srq5X2e
udg2DvXV0IjUPix7Qo/WvyHXvFazaYV0LbaW5ZRzUsyC0/zfGEHdFJMrIwiy/tdD
by9rULR+9ClMb3NhmR+nyecy1dPEHyosMVfRY70HDgITgj9GxCgFi6llEc1u5p7R
tS7yc4mlBobNrDk3cvhWNsE67TyXMpvj+nMfBCIK+Xys9UeVF476EMxzbHNfgb11
FEq/Pcmo1x3wgd+j/S8qeOq6d4cXmT0DDxVc0cTUiZAbrKdNWHBLwoxsbGFGApUg
y325+O+X/n8XIT7/JgDsKMxLPPjeuWGOK6S79jAKAQ4NLGQzsZO8nRoFRYbhaEn4
+J9ayqkBhvM2jaeoKNNqs5kVuKtPK+H3CtNM7fMVhRB8jYGZb8JhZKeA/2v2ru+F
gltPRwybCwCBOME0uCpnKZoJdmR30d4UOoAQTKr1yBWiP+RZ2+wsZrCRorhaewnj
wShp2AcRXQEdxOl5qo/5anFgUF+weKxPUU7iWdqJCt2RkYzy0vPDpa8CjHTVOrWx
d0c8DgjhgNEXSN7xh3CXIU/OGAlAKJwO5z989HlH7wC5SNmhPNw002DksD0p93mJ
i6+OIvy7sW1pS9vrspFyzijGLXddzOJJoiAfpCnzOLFBT39Vez/BNvCqNAe5aE1q
OJYgLTMgyMfoNCrN0+uQckSkZu2gAoniNgfHvyuDNCj/XQdyO7fz1jV19pYr2P0s
bJFE55Wks4jSZ164yV0AqNw23wODzONUxUJ8jDE1zvkdKBqPTVNWTWwLaNMsp84w
ezCZ8hqdv6/1TSKe9tLHPyl0XldWRBsC07SwTMD/S0w30QERH2BiU89BcxzMEFoB
RSHxDsok5o1Fs8titOAIBTucpQeNUQAh7kif0jEhN8y1oJMGhftJPwlHX156tIu/
k/afCZrz6YYsZG1moshhRnjDbfFjHGsGoO9pAg9yC+fqjFBGKGrGrO7sxWms1gXa
/tENXHXHAsL+Jy2SxQxOm8yMPTLz4T71oJyWrhutEwYhuoitA+TgZf4hajlFKHC8
fyI1swYuSev/Znh6FK3tvs5gdQMlOHZgEsoocQcD5t/khwHdVXX9Zs7oo1DA99lJ
MdDhH3LydDKYrhWuZ982AQ/FJ4JgwNj/oZs+HCXLfYLTpSd6sHu3l2Z45XiU0zCk
gOQgaleTigpaBznTbor8lF1HxcX20Y94dnpsG6hEyVvYyiG5TqLpD7YVF0htJotd
o2iDNr91MSzctPzJ0suWmOR7uQ8jXb1sP9iUvm2I2D6lyHQm6oOLhLSiYXljVUEV
zvpMzzhOxDO0WAFAJWAf4FGPhq0gSQOuGLIdyU+GaeqlZyH3P8tTr9QKF2kndI1q
AjrAwhaCQGnWZ7Z4scWHwhhFpsG9MGCJnoi0FZNRWu0X+DDWT7XaKIlPX5/7El94
Ut8iZFj/lZyYNK6dlgvI54+rydu+LtvDt1qXNzXYgsZf9RPhSazkmxNxc3c00sNf
/uMMRjUQE4ujPZlriwu+wka19VgkDZ2CpHSHUm29YPMYWQIqyjLhnhWrtUGsiVtp
Sq116WfJMks0qW/dYHd7GsVFVlsC1iWu4ZyLbjNislO3RdyMTXI3vCQu/4juEIYQ
Z+4fFQy8wx6AgQbKhOM7LXmwvG0mA1pvNqU+GkJQ8gvZb+GDkJP863uOz8HZEZ7L
5A9wD4M4WiiEzIgkuWHk+UYi6KDlYqscyWMfAJSZYSAzs09hNJJ9W2Fep4X4HCb6
2sbCCsEz+NcBX6dE9cwakeH0c/vSAnE08tBasYSFXFpjuPcU14pPwJIgrXo/dmO3
fUMmgmndFd1LpfMlhN8itagI8C93P9kN5vEE5otyOT40zDcIB4VZCcbxhsTTGscz
JmPtPHoI8h+MmNopEDXBPntCm1cW+nsf0OcvfkokHmyFWkJMGn/ecp7VxVJ1Op1j
upJyj21RbIKrcMSgPg+nS5hXZpVW94GoOEHXHJXZ+s0ZiK0w9VkLh6/w6rIrvpz4
jgmF76CjSMWKs3E4VxNhoBADqFZMVDt7LJeLV3MGgaYtjHpHzRgRBDKgcCZBWPFi
yiRifwM2HIv97MhI3dXuXVO5v+tP62bxJYK2bZGl2ZMs2WzMlwowSbRvEleDsFzG
e5Cyp08/qvmsHDxZxVAzS1rE0WGGR3Bl6h1VWmtfT4F9ylVo60DZG/QYMpDvMMjV
yZe3gt19sQGycpXZh7wr90YKg6UfReUNJ0HLGMnSFV3SpnZ5BcaZUYqT/2wmrUNl
E5zN9M943e0lo4ID/T64os0icu7O8WCWJK9NRzLpiHllqdzrxKV8nh3pb0eU8tgo
91PQsXHodzDrGAzoJpldPBK8bZLgqDTbIkimZfe5/AOncftgTBFzSWzsbufjkRKN
62vLZPABK1ITVdozT83L0H9mAdmYC2ZAo1ajNYc5pNLIzoFXO7ps433BQ3wWkMSV
BLapF1MPJ4zglZS8XjQ6+l4QzC70u0tB/GsGxFhPpThhN6J09bnWTYGiPKWk7nBQ
J33QSqEIhTKR4piHhkLcST5GQxjGFksjuZw24alTfRKUpIqRfeOGdzkOVY425y3o
baQT9gCUExJA1Lp8JhJfodgxI8nGZcqA60+jYnAtGu9OPhSQijebstpTA24qgcYT
GUZCLMwWHkbfMkpxP7QTVoam9paool7DO1rSbfdVOLYVwwUFoWAQ/8i2jslZxI86
Z/51l3zvOS+wb79CZxqt8PzuFoZyk+TdOdEBWaEq5PlPpQde8hmayW5NSblqFvKV
dZp/QENCAhkFPf8ajyTjXNtPxnOaFPuHEiFWUUQLpy6r08l4gRyTN7KBtsgEGhT/
28XkkNv2C8FrFDZ5cRWwpbGT9Hb/JZm/znZfwGO0n/nWlKvMuVo7+2cT831qFeAR
XNnqBuNausZ0YzZp73HPnJ8RwKBAtK3a8UelsJf906bMGjsitEiY6dy0lms1LqSM
Svk/bvzLpXIFlD4/7ruBxAixY5A3L0/U+JbnXGH7LjRHQyyyIWwObddh8aBSIV7C
xE7W1csdg2F8uIwLy+RtwxxLGTFrm0vEexzfS2Tj33Xa+TD13oempAf4SMaX38xU
/bxVCDuAxSbW5C9dFAm2+Zwn1eKnDCTj2rw/GRO3hqyBgQbKYIyeHdppzbvtYALG
sJpWxNnaCBa+2ihMHDhg/WJPrHt1Rqbt5nB1mnEuAMUma46LRzJ85C/OfMyFFHBf
5QaSUaQjRuE4AxI69GAP84c8qSqK41Ro0axwV8qez1YUInLhX4g3xJvnxYglMtCW
b1WF5tJjru6HYEWD/qi7E6s8T8lW4BLRN/2gXwcoF3sMPATT8AiHamHbVMwZc1HS
WCmMMBjWB/jjVLtmw1QH3ZkrAg6V3IkFBYFNx55+ceHVnVtY4SA2zc4YLcsd5DHZ
KrWm2+qTn0IqMABtZ4JrpEQXM+c2ZXeQ/EseEwNJxUVt7Q4fuVvVMY22nAmMwdW5
uS388pFa/46yWyvqx830Uh9Md/4r6hXFiM6B+vZqhvlNOEHuDPk2AMWaHZa36KQ4
B0/9952eEISBJtriXhLq+YUm+ayzLRd6D77FdB2tlUZbEbru3MADbUILvHmILtus
UQ+rXcfeIVPFLEA8uarNinyb8xCFYG7jKygBotIaunHTkCvLKBkIKhi7V6Tda7FT
ZpOd3G958WjhpKM+63qGNJSwpZathLxMOGER8pUyiHY7D7Rv9QJMjsgfn0HG2VW5
MxLvrZe28lrqaXm/iq2/lx+UyG+1Z5wr8tIy+eNHsq6Trb+WGhoqxgFVlbBzxVU3
jvJczBhdRq70+xGxhbjGaaU8ASQwZZb5YslQqB0fU7tp2n4zLSFdtxtKNqhbKO1M
IheikDv9kqeaRxZzLCPDwnyzn2KpZDslN3swIdcf3orogn9gCLNbsMikXKoKem/C
woVmCSLOOd/HXQ9QwvXBtXHK+FGYUAkwuYP4YD3yI4Ju2gQMXVwp1n3BTZQjj25y
q97pMZNz6dtHktd5b3TlUeOq2DoQY1yNRF39hVWwx+ihoDGC4qhBEwhp5TTO24BI
uhT9i/WJwwQviPNH2CLa8HD10hUN5z3G0fXO+VGqFmp7xAwPxumeiuN/RMKHe7rU
v79S9rEZhsAelwoCu4SihdwdeFqk3ktwHt+W30qU8ezWk+BX3ruZFZ5iXKcu8xxf
AvcdTFO/krKbuyTtLdWEas9YFktQ0RCboFL6SkV0Olj9eFJPeN7fdi997/WC/eBE
O3XqW6mxS9MHYTWs2IiPc/4Khzxh/71A5Re2SB2Ac4g+YOOTy95VUD2odH44agtv
6FIlbGjUXEgjwm1J3FFRi4N4su6fq4ldNzXi9U2keMlATRyVsMTqkXPXX6BSoR0e
WT02DD8QbgPg5RPilP+/ylWhlLrjYEvQlxJUAiw4mJlz69n9DqSbG38jhSHp5ISN
/UcnmFWv3SMxXBCEy35WJuMofnSMon0Xxknztn7wUiFB36tRnnNEOucDaBrjkApm
6kkzc7TCyIyr1SYVvXVCeRXAAHKOmxu2MBZW/7P340LRp2pZj8SvJBN4gxsRLRR9
d7KBaRnIz0Z0uBpB/uUxlrHjHMDCYZjmYWhYAWD5oDJ64OnQAoC9K3xdFwyL89X8
b1zw6HW3/P3LquCJZU+3i9QN62rgKRtiLxym57iT7KXhM0dyNBOe4XkrlIcNemhk
7IW8mafbn8l7wCZmEnlea89kFdZqhL35FacCbZ+WVgzWgnhj6j3PuVlyWuVWkAMR
1FqLaMueazCFf66ATlzsdAKZkJGon9oB+ilJ9IGdB9S9T2YoumxnBTSaIYuzgVS+
3wpm4FPIt0iyjip9T7Hc/mkGdeDJp3tpT4BQLXb7R03u0R0Ca1iFMeRqNRLSJJJQ
eeVjl0onkdrkPGEc5gQz+HdRYTwSuAPzFHnytgFqc+ORvItyDnwq3IPwcR+NyHAC
iK41ZieBi1BH1qjRdP+lzdlpAx9TG9h4fwTqAppcD1TdV44usOCchGrfw8HBKCkV
nyymRi5ezASLzrFox+tEmYJW2cLWNxyHPyqAGQYErg8UDoB4/5eRVnuxFKD6v2p3
Cds86gdKGLH4q3netXd9bSTA13vZu/nUpXcxQCb+9uySHCT8g5aOiINRoha24G7c
jMm84hTJfh7qo+d7MN+ZssxbI8cwX9+ap4ZpQ8FCkRXV3jPR69j9QxJ6xRvwT9Ik
UfJNReuqZUZ8BhEjsWRbqeOzcJJFUkUqjDamrc6YsWZ/zgW6BFen+/28T2jwBAxn
dvJV2DsDBtVslVgZUkSvqy4vqt/6pzdYe25PBVfiBfl3/J/eZywK58V+V7sqLmcs
2+vCTL6fVNDC0NyWQKVIGVZeYDSD9feL+c6yVactVAEOBK7Om0IR4xqLOWTJ2CgH
NECcVPrUVMKVVCVeSaBsq0ofSq1R1V5jftCnGzpU0+JJiuwzSkEBfGiQtr7ZvWu1
E6lHWlh82gV8vM6wLqqddzpFqXvb+MBisEsNAOaPMfzZc+Ecm/ssWbZBfWuzqNXJ
Asw2VqrlQpNeLz3yHUpDMKs8GiwG5CYjfd8quioe3Z4fRYwLVi3ToiNM24ZPoitB
PQVaooIMThXVK/92sr9OIFRl2Kwbf/KIOlvIqozmCOlP9slJagnP1iDPPbDGesA/
03M8xfZ/kEdS5xb2BEzN8lvhFAmLTECg0wf4Ca/EpO/OPKpa1AkSh9mEKhOuZvpe
0TMpSQ2XzyGz481YouZEeNI+rCLBtj+pfm/Blto80g95IEcQ3Du7OCSpt+YVY9V3
oDSN6vc3Mlsa6hgxcaQkTxNB/jpSyBd1xEbbwCzeXPg+pE8C+fiJMkopgSeJHPON
J6/JMDAMNatKO2NyJtP+v+fj9yTqK9OQnuotWtyiWxp9F6D6XamgUPrO+j1CC4AR
MML+xH1UYau+EN9x9QaNGgw0UFBotPiFIT06YBDnujNFaswiX+1D3+ExVBbjCQd5
qBb4JdHZhf0Jr52ncm7UrQIk6f55m5ZtXv1PmKbiaPdiEiwKYnJ5HLpYKjoos/wz
Xcb09tf/bd3NmyGKW1t7lBkKKAOgPnNkL9ATLxBr7kBmq3jxHj7NkMPUvj6ByU2h
S9J8f6PIXKT8liSwCLUfiypwFYGFaTm0Bcd07XG6TXWNUa1Cp40cPS9gyEZJtKtU
VQVWxNAsYzbXqNNVDmYglwr1cAPcrROUaY5GofOgrCgDAlfkXwctxZcOcwHPIZqy
cPqtU76OShuBCtf/cq3RWZtrsHr25Rmlqt8Dn4LFNmC6y/6tziwMdfJDkAjtO1RW
YRQ8vjOx3tg4HCVvh8QChHguXU20WlGbSUZ/groLr7T1TGNV2kiC3FE5vygMSr7M
WrggylNq303iNGaDzdhTQj+EQhTD/une79kjWgaiVK1ZPpKNdDMZaj7cxOoS1FXD
JNBRzQQFOcqSt8Z8yK+tLMIT15Noz8iVV7Lg7JMpNLjY+v3nl+1DF32Fhtfc8dn2
eYKpKAK/mE7BadXt91SA0cPHIn7Zi5VmUEmpQEdG7Mt6g2XPENetKl7h8V18rwfX
lniQHwCtlpbZj2xPm42HNUvh5cfeatlkQVLKofVbPL2NIjroBb2aTJfxva5uQK+9
JsZPBGqdQIhxYZDWEpARHfSURpT99s2oqFns/UXvBfaGp1YAuRbtj8+rcDJMIB0g
PsYGoCv7gNRaJ7mbtoWfPK4ODBcD9NjBuf1JyJFtIy1pbhsCKRItpu8Pfm22bGrG
FjG3WHwD+Bfc5efltmBErtBvBHdm962uFguF4QEhGCGo7LNy3xTxiqgA8SlaHXE6
Nf/oefnwOZ01MC6NBtjzkUi8cU5O5FGZq7SnhJdHkL+9KixPpGHi3xdls5Izs7y3
O6rHZzJEN05tilc0dYqQlxRRVbXnk7eVuMk1+GQFaoWBe4FBvEy8l31n8DlBRBxo
DztMbjKuDsMrXb5Wl8wE/MIm15qEgPwUCezbjYMEEa1VznLXx8QtTYFQ1/kYD55l
SPr+DcX/Xf48WpUirVhm2+0MQhmdsZT1ShsgTfez7tIc9PXdFaHP1lNM4i8+8SOg
T9nsI2ngjsyIHjhylO4lDrcBo8MjvTFlnre2ANzGMxbE/TgjatQob+SjgciYmkut
fFVrjwxGfITCfTLTT5TPJE6xq1hYJe3dEeVyf41p0Tt18nl1XC8PnRKXGRL9Znxn
zoMnSDNXGCeiSrEkJtIEZ8xrYdTjiDoKmnHHQMGibq/OsoF0DEKGahXlreGLqgFr
DsrZT5TMsUWQs6paSpznBzF5Av5DnbAKVYqPlQSUBVMj1oAJRfdKCllRqxbH8Vzc
NyfJ6j5V2iNwnzyasMfeqKDmhLbPPNk86Sodr/6ChfM1iEDr44TiMgQZD32f2QeX
hJKoysu7ZakKu9I7wkTdKVwY5uWoIKlrd3cXWRqjlujjs2VDu7YJ//T0TEi+Ag9G
FIxMZbkdzSmrXaUPgh+VK2kAtzOE4JS3yL9w/50QWrat1MPO2GUVLXEZCaMikld3
wAyHH4gJrxPo+v+isq1rT2/c5pmXh+tvAoPYVedKcZxRFiMGyhIBLkQwo4gFShht
W6iDyTd1EXw90W3r17ASaq0yWheweYicWGYEP6382/3t0tp0kGv+rA82LpkwcA6q
LzSJYYQY/Dpa+WBNTZqT7Lf9poycNanShcBmw2hAsSX6R8MlQdxt+v3kIuGbmrJd
RTjaHwS8NzzBrnirVqeqTjKrbhpn8nQl0JAoifF/imiWDsC0AoOJNMTDL1g39mkG
q74pGgjDMBFVEg8Vz3XJEvYGA/0e+s38WSYAcBvjXJwvmV/UTPw2B1UkZ321GulO
ZFs3Vw4CJpoSZxNkTVVLtsBvhv/mx5YTVtuZU24JDK3YbfGnZZL+A4ebk6SplA3H
46QBHDP+2wNxtCOH2cwHSKTVWYpSfdm3qxsnb7wJC4miaGENZkMsSNmbukMAwJrs
00ns5ABw3DjxjAYh+rYuHXwpJ2nAJ/IuQOKyvBrlATm4Ct3vcXrISFRuTIeI7Vvc
Nbf4qpfS1aqFgeifeP8T/orx+qcnHippmKHANIZ99N3ze7zDCrPGYTWoIINy3YlU
B+4rKwhGZjfAoV4P9ZV1OI4o+ndxq+74o8WvHi2H5P2dlZS8ClJWAg9l3LnrSCSM
VfS3euyu5Zi307Xxd60TIy2sPzryDTLtKUWrAmxUMCu183ZxAvXPL3geGJjV4ZpP
MQivOSjjd0reSXUuphbExnGGB3xB2R3J7a53aQXL1AFcWDxOEZcvyH83gEGz0DAP
3h8cpaL8djfHVM62/deqq4RA3pcxneUKEKjCrgdYniQGK92zPBfuREFWSkY+s/ti
A4CSHRWXkQUSN1DwflpphNiBSW399TVisZzdqc4x9W3EkI19E/YBbBTnwlcSLzxj
GzLz0NpnmYYVxB89j4r0XeZHeyBFnWgtll0Z08FBEIyQLIfhSqDvcj3L108wxFJN
76+Q2fuuVhfHqzDpKPxZmfuONBvLpf8i0VK/7QsJ5UZooY1ECrtgUp5k+NEzkFa/
/3+8lcUYJx7Nbur2vrcIYja3pGJI6aCp6RqITIKhdurMT/YTNH2eT22ummdR1xAW
FIx0p04MED/jfSc/aoqswmoheP69FsnialC/jRq+UEZrXfRmdn9hjdw2C42hFHNM
/EoOWgShfZBLVCHJ41ubWyEwkfOO6AyFzfL1boP9vDsaeP4Znh9MgcckOCFLtc+v
t6+nHr2QOFl9U5lLTpLBVbQW5+kYJymHN923EIezwEVBrHQoiHBjs1mAou0tWLo4
3oy+UhcFKU2+xY8Xk02/oirIcuyhcj+oYTBR10vnQOYn+ziujV5/CML8K5zol5Ui
23qp534e7E+XB6/T1a4JUQmr5nj/3zW/886Wwg1xYziaV7eXKAFBc5f6Lps/iVMk
+SDTSBEHhPeu0D61HMRj8zlOQcCaVNiSTmLBlMOtpnCzqQ15eLuI9rYXS6E12tx8
dbcyqdM3ShpR6AmKtVbLQImiNgcepsgroTywo4M3t1QHiT+zKlJvfowHhlPPkjLu
t+CXTam7pCVgZHQ/NUcUZtctbB1UtMZvyElW3rgkZIdPee/fplUwHprW6VzEdKAb
JK1GSbX5ODBcyq0nyogmocm0iBCyVwOx1NTgMCbfZ2kderDjEQn2Bhtj6v5HwJ/J
MBN2XKQM814j9pTjj0cdLSKkeC1rA/SjqYTTk1P086+KinrYBvR6b3mm4u3DbKfl
Q2VKVJmmkVZ4vqc1feqroasIoYjNZfeXQozyQ060JSlZI9hL3BD2TdQ85914ialh
Di33DLirFQKn9xC10E9sZ4hTmYvJIQ0iwCOAuMrgz2cWGSJ2vPwapkIVzh7XP6Xa
KyVUAYaomg7/YyiwSfg0507mlbRtSd8zmZRP2D3VaulteE5jSDtWAP9jl94mmRKR
lcPj/d762djXIA1xkquvg6WhKRZKua4fKW+sEgSe+FDV1SVjyGugVIyQacqwsjmy
t1KKmuq6LHJF2MrfoZUJkiXVc09dJWE7cnjxvvb0MDoYzQDYO7l6tyChbUnPdAeS
F9X4MI3xrBCkDSOG062mHDVr2vhjR223Zc+0PlP7FSgIH6rIMGyiJ8jq/ErgZXJk
QY7pHdO+kpTyyeepIRR3P7uma2wLmDgvxERvsTlLQ/BcpvJCu48uZYoxUHy9ZG7Z
0ZsZ48V7bPfaH/29T9EcWDqHMJSzP3nmY20vYwOIT46T6VDJeX1ZzuPk9asXHXyK
rF834UE4/AnFyXSowvWtE+XZdHYU5PcbSx9ZSGBknMY0mg6MLg6jKScEHTgMy6Fs
6yV3oOjRErfGYjHQ4BHuco0xUHHxh3ZfFy3GhdiDRjoViT4o+cQMXx2L/jskk0Ut
JH9FfV7+jWr0Zvc4HRUz4UFxNxdvzK9FfX2o7wktreEtemvSQtDkwvwvfPl/aKrL
k+4UwNtNvBomui5fYaXUbyY/FeSFqBxBqnuTNgB9lPALZGKZVkh1C5WXrKk1gnh+
nCyosc53tQWKPScPQU41dSItxRcTW1zFjL7RnoG8Sf14wrKkRFULkoRfksHHxHms
g7OHlTwk6IL57xRyEv12+yPK2CPAh2fTwv3vVe1vQ8+dc79tGw0vYqSxsx/pNhyM
tMkOVFweV8WYikGc8aJxB7o83U19P9hqo/KUBwm8o83RSLVUp1TyxPQoJMu1lBuI
BVOfdr6bfD93qQSo6ph/uecsD27XJIlTTG7qIPiNgWOjA7nYZn55Co/oxJK8ci/H
J6qgbrbk1HRFsS5SCeCsWuoOa0/DeM8uKFbMrYwLNeoUDelhtJYExOv4jAOrzqK5
QSRYL41RoisWodlLReovFg6edRkQTizm+XmwQSw3ZV3DGQ2xm32jQ7sNTTgBAaqq
dK5GkGjnj4V6Y1MZOvUptBalBvLEi9DBKgLaWdie89J8ORrtCrS38GqDEcCXsNzr
igHJBV1gSHL4WDqCUEsIRdh0YDUr7o2BBor50eEvfeLYIebm9JoDy9Gb8GIKm15w
/Y4pa9YaF95RD3dVP5QGLcgRV6eWTVkZ2m5pqpvkr31SCuAivXws8UCVPEFN7tK0
azGvGR0LAxbKPOqp0FBztiD/VfC2KIrWAXw2o3qTeO0H8+68scErd0nFDM2qNV6v
LWsqiiu3Ix8FBnb6Fglv530qqE0ki767dtYBL6C4NEzfgdOeuRoKbJdDylCRhb5A
5z43cpkBs72iWjNBWRwv4zqNPj3yZLK8Cehz/oYPwhNUqu130kqqUObUe5I8aCqk
XTQtNyFazKXMSdyQgPBCXQMbvD4Qx+K3Nz0E62O3oU/GMyCLyxwEZz2diEigPVLe
ExvSexnBfCT3Ycy8/acITvQbkDGIXH3zOgHh3XACZE4js5mHmOm+mW/Gr+jYTeSv
6Zz3pRW0MtRmMVJaLqMEILNih3JOPMGSwwgHVaJsnK9UNset7zZSf9EWOwnH3pbM
GH4T3lcsj0H/mIqRCreE+ChqdBc67bzOdTYVMDqIs6y9fZuTTaIinQLRGPUOM8kY
A9OyZXEu/ycfUdERT7sB0Z4radv16B58ND0HVTRB4WnSsebkhNCFocCVA6ZS0jGy
pHW49KrzNbxDNNau5ABNC4uTCBT5kph6g4Aymb5s0HgB48dANVuWYuONFYlBxLn1
/a1tLcZbAfEaUQevX83Ym5xZwyrH7onODfDGUvo4ix8wb0sSD/iPmsqn0akNX/Vz
J0OJvxApkkF4OlwsT4H1FF7/EXVxu91Yviz2PMhI9amFgBazLOgolyxA2o8tT4zF
bJHpK+ezqAYpWpkUlUMud9N8KUfOv2Zwz42pv/YPOiAGvECnK3xRFcO/Ic5EcF9X
KP4QeAJ7Q4IijsDT3tuXAo2r+qt9dEtMBOuO6eMMBKqeZZTOWPgR6TaB16JJSPB6
/6ZMoLkb7DvElTgfXyW67tdFVQksVzduAgLW7jN+uRFqT1EcxGMNRkjBgMl6QiyU
mk1vkBbQMqUMR3ALkcmEuMhrP+MglXjxbzDwMAQg2XDGugxUbtWDblzz8gx3XWEU
bvutbkSj7TMQVMVYugSo7+bjoZvJ86bC1jh46nMcxPL1Tb7AQEWgDFs7lI712HPr
aEe93AOqjvHL3c6m+F+GSce19EkvdjF7GujhIH4wXKaPXDJ+8oyrPcS+Xy2ZNwNo
Pwnd2ibd0UMbQtfDZvd0T34FJLSxzkjSCL39+7kqF6tkWcjJMEpD9ClV0+uR10RM
k296SwVYHv5da4L/ON2n9iGpwhORg9uEnTiHFj5koFG1h1AgHVCN+I9td0T057zh
l96lUpkNR/6+nkIJxTdNMT9SnqEg3pthKD69tQyemC60etbYsBX7NH/sHKguVAAK
iTVYidcp2tJXgjXKmBxYzmjJN7Nbzz89R8E0AjQnLJYD9ct8FiSe8iqMGP4mO4IR
i5/uW7bCOoF0dWMT5Cp3h+5xFYnf2jNko7oJYYMwESvQs0Y4N4TsfNZSFAaCGAvv
cWZf7bHjbrIitymIw1Ftm3TY9FBj1AF99afYKdnKpXmkAdHWIlRJRogxk0ihH1eO
AmGxLdV/jyc7UOZZRTnPYFhQj1pG8UnRwD0gTvRQcZRd/VGp0Uh2yvEiwlTA7ZE+
Ee8eMp1hCQsDTrGYYBxcRN4WmGXnVMbIhX7bhSxcMIpFc9PVsJfIvS73FgNTGaHJ
w51JmmE+1JcyRGZGz+80eiQ69kjQ1BThbXapPRsL+FMGiGMgdDEch8VIogBsz3Tp
Xqk3mR67IjcDnkYhdZ8vpObDvGUfTFEmoLURMYijeF7YsVOtM1j85jEoAREXq8df
4Z1jYQE7I8+qMEZuM7fwN5D/2RIu7vLx79WwqZ+n32BlJfYPXYKRsU+Iby75rjKm
xejwS9UyWU+BHqh4qCVX4HXQ+2xgspQXS5k92UPtduMNT16Due+2Vb+Rkh2DgzGC
btg1qDoYKgb+D0xq3Y97fb7nKokWq0JZzU0kgz2Cdlb/dCPiSUoxHXPqfQV99TSA
8calh92ZZ+JXevyahXJKzDwGlTWr0szUgMgrg/K3v0LE+B6oZ6rFQPR2ocp+Yv+k
ooL8nhWcDlyKloTQTz5jTqePAKgHVkYNXf7sq2bKGPbYWk1uZj4krj95KGG4tORg
cNV2IymDIhK2gfDRz7RA/D8jR2AVfYGm8efq2P35WPZXqJSw9xYy6beGqG6c3tfP
rQrxPjuPVMrbENZpN7glVaEoQbZcT8Q17ecDYjsWpbOuo+TJ47qt30HzRKdbAaZu
S7bMB3K6u3lSbScd2HjSVm7O9PUdGAqEGKnTNLqrG9wVhV16T6quR2imL020O6HI
KEjvATL2GHZqs69BbEHjA4cOaLMHyjep/T2c1gbGL7ilmY1vKQP8d0frT2G0RV9w
sSpr2U0zECqtyfHzENP7c1XmhX5kw0xSZZTbIhaD6T5ACX/ucC8O0uPAAiPyiU0Z
wjaCYKvvMmh/VGEthjvdaiiyCsOaDalMAbxhZE3vYv2mNp6SUMZ5jcA29IILZbVa
fdmGkMZ1sssAn7F734gnXAUFGLySAW8BesUJbguYoASqDGucSpfOFD4ReZR4btQ1
J2ogFy48chFmtFeCwq/VeQhkVKc+yc9ap4+4N7d2V6eSuc5JBLEB6v52bJTwQV1X
yAAX7atW/cJ9+kvU0s+ZQ75/vIXhuqD2ZKsOo2FhgiwLjvThYb5LqBZo3Z3uZuly
WwJ9hFjHrdYkBVX7crxQTBOXlNMcQMqfLe/rKdsIuM7AbQMn4VyekGvpCuWgYrIR
p6EsHoafgPK3B8TNUn5rFBnK0KkTVfmxDYOXFex6vt4N84CujeUL4tp/ank4aHmx
Cvc8rctp9NIwbrI0gyH1zsDdEIiqdXPBocuYObhUOl1qk/mo8cR9AyFKbl+x1IMV
WkEe2d7d04ELn3rIE6Z2BSn18PtIDkEd2c2x13KC1/9GrjmjLyAQ4xRh7OLKB5Vl
AZCNYsnr0yx68BcEpWNczeJUjBBuLF161m1fWvn4nHYsbOLsCsrfVIcf/Pj+f4ze
ybuN94Q+Mk+1ZF0fph/E8iHpeUVNGdf8jtmJIuo3wfK6am8ZfeWXDcHQ7J9eAAFd
cJlVUmFdYXkUd+UHAndduMyX/9CBVHR/8c9aJsOnNbWUXFaMWFqs+hkG7W6EZ3d3
D+Ke3voqSZz+u6HqIy6kKlQaHylvgWIz1njGs4diUXDhUO/fZiJFCgq90IizsfL9
1WEHSkxaL1ra+gANoDyDgobpETVJlv0mOj9NxfVGIFgFYuK/7UN7MeIzVcTyWrMO
cmWx0aG7wfV7mCCFCzP1Y7Fy/iTSB60lc+0kx7AVAfPxscocWYFDvTVj+Mvhp+/H
2gXHdF4jNAwxOELUz7VHGxYADJFp8nETIbTLIVMu0GbwNN6HkSR+PTQ9Dg/A7arh
uBqFssiv3Izf/AgHof9fdFfvHmZqnFkxqj5CcioiCCReEhifIUR5cPqj+xiSMvwd
7fOc+EeMtBs5wUjEPM+myzTmQ5hDmtH8xoDon6Gq7WRhh7MWiS7RMGb5duEKhovV
maMFv+57AjORJwbI9oOObFw+2gcDq3dR6i0XKLFC4Y6pztfrhSd2tryPSV2WAR2s
ELYkvejNxKtDaBG2wemWo/vaqG3XrUgjfSLgwQ7QNkjJZXreRVR/wi73T4fjSjZe
SEP/81yu0OBJyYCy8aGQVJrHD8W5zeooJ82dvQWxruzmMfvfSJlmdFL/R02o5iUU
3ZmFBXvrDktaNn7JtZ+t28iJyzIpyOp8ikELR9boJi7kc95w5nCq+SFadhoZJdrN
MpEq6zx4qDRxrwF5G9FWFUjP+Lr9zVjApRlMG5Ya8RhxDtmDwEUX2VFP46Kdt+MS
B9+uW1uUhyOkljnuzZwGGVM+pjs7oorJVagEkyETnrr+BHms3RwU01AS5E2WX4JJ
kQejkK6B6hl9X86TuVYlLTiy6Hnkkw0qmjLy2PsgHufroQQIEsiAcXc5Ns1oCIWr
HrQDzdbx2SNGReFCWxrWTjU6+sz5IBsx3bowLFbGZCGy5H677baFmMV3A0pKrcCD
P+mz91vjwvEpCjDCSdjnD+BOj9p/4IuqoYPq9pfHhRnwzIAZfZ6NNs/wS52ww0qz
w7wSNB1GPeeMLFNag4McL0iD5ECpfZ5LkBAqeDuNkFXgdMPmrlyqPjFgnOT7nKz+
g6APY6hx0ZW3EBHuwbzbFkkDpcsmiWR+29H0O2zz/lStZ49tYtJZS76Ne4QLmfHJ
D5ipytkcs23CPri0QT4Y3DbwsT/0CCqgtkB7/nt6nn9xGJXCSOGPoElyHgSFX7K2
/wOffrpe+Z1j3e2aYVmHkF4vzGSlQdFRdReZhSJYgkckXGDuyNdZn1QJkNKj6HMj
MDyx1AqWDBFrmimYMLUodcmURpaaGZPsJe/wB+fkdddUkZUoTFb72fXjPV/2jTtT
aU5k1CuiCBjTnBWrnu9yzWvejyH8cAU6o8B4QLfIuu408oBwnTMmNGdTxuBGHXp4
TsXsJ6Al17vPPxsxI7Cm4YEGO9+1NT9VO6XDPfs8dZHh7IG6EMmP3U3yYiW8ygT+
Jwfx9ZRxgTWt6w3vAa1e8yOcnc2wsE48uzJTGX2OC1vieZGvBoR+RIAPBttfYHiO
pYSc+0I4eif3zYaREwAH6JvUZElXwruFhHVoudios9MdMOPI5n1AU6/JRWre7VTz
jJLtwuQjoTgwG+Jh5xTZr8XXDBgnCKI/MnT7+8lFOugDo5Hsho/xRI77rVj2B3Dq
CjrUl9X7C6Y0eKfNiXRymacWfbDR57ia0RVeOo/Rl+G02ckoQkMTh81bKuO+3wcR
iDpOUtXswMsSNyGFjyO+0ewWDRdXXAvcypa+A2uDKMZrASzbF9tRKorFxE4BlNdg
sO+arJf56hrUhYO1Ch3BqNEahKK1UknL9PJF5e70lm9m0d4EMD9DQi/x/cReX3iG
38mAMi9UTu5u7xGUyyfGvq6BtZTBXbD4aqtqxRmnd6q7FEKI6dFk/9SWMug79DVv
wqPPdIGEU5unLB9HXItz7gH9xbkKupqlMYZHs6MWY2AZhJagw0+TI/8kfa1Osl3H
pt+K/NK5jJ4eKSCCF6wABhAfvjc5TTTxU56wdIeXXqqJVabWqR2FF29kyw5+4PtH
VwPqBPOF0Qz19fsuM50kn2URFNjBgOr8SVPhen4KqjolOggu8nOtZfqwzMlDFo6I
RF/wqLWxe+Qn2Vsp1BHSzgvs2rqAa0s1gNdGbFKbMJx0m3QCwbfJb+AP0OkBlA+j
ch38lWBL2e3JJEKLsH1qlqADdFXQasomwsV+xO/PaXFhoVz4su8zYuCnQhruFnTB
VOxFKLwZho0JWBev6MfOvdZ0p5/A9+6FAU0qjutawN+LXDk9Ne9ekpEb7x54l75W
mdnh3/QQmCgc1QJEdSYUDRtZa2/+L7ZyYGu/fWkpex0DX+1dkN0SWNcwL4T8IXYj
slWjnmWMeNTkxmaKnt4/Dr7Lvg+UZZoegPV0YMAI+SNhZMle/mWW8eOYAIiyCGPd
FZk+k+2JfJ7oFVMsbjoEZynfBC4Wq38roZRd32smzZXTuah5/VPkZpGVRjwcGwK9
RqxDqlGHdz8NypWFzZZ92be0sWSVJDqYG3X5abtDd8SpTOjXa/7IrbBCNVRQZqEM
IluWNi43acA3qTapV6ZXA+qHwRhJAqvydTmalVqR0bhVzbTQaks6wscelMlApR3Y
BgL1+9eDmy7DxDFB8YqtBVbgDdspc8rv96UuQoWCcLuxAVmnZ3UQiRumR4z2IjKV
ZO0h1FxImeA7NtZQA/KIGtDUvR3mhpPzQ4HpcZifT72CavRHjXbfe6L4C9IwwBAi
ukmsghxon2gVrs1ggtFesWlBo6lEI22WBZSLaQGBy/JAH+ziijIs5p6tZUx2i/6D
9N984gbHXBZRUYJnOLIx6dwl2m4mYsRhqng0/MtPhq2M0s02owyD0LLWzOZZcvWu
HerO78jnBvYXRJivzZJGwI3qYPzCySeem341M7+lS1t+KCKbf3aRDRx7Y9v9keuM
wCwLHci8TzAPpj7zWoc/zS83p6HjmFT0PrZfsSqMynktLplE3J/E9Z9up93pex2O
SKG1Q0q2ylgKqlGUvpGH61qMd3OPgxVy1h8azZuD+j736CilgbpSIHV9B9edC+qc
Af+/+66toSJUk518NZ33GrvXS1jbwtFPt8WwNhiQWTSOYPh07NBlNvQuZP2K22ae
XLrj+mm2goBQN2Ka0kdBnfzDsMGLgSX9/F2xbevXHP/5nUzq7v+doiLp/O6yAnxY
q6Iscvv2RfwvR6A6CHlDHaxdJxzzbs4lupTvVHS9qS1RwEQSo7QIIEy+wgcwwSSR
JrxveLNNkTWiHpBGG6WXPOlMXOdI3gZZHrR6jiYJzZtXn1Uw1MWY+BN4FjVtewmh
lIHzbGIRdTVDJ078OzEdGprTrr6bLiBKekqcil2aBx1BOCExVHLbwrnJ0MSeJFEB
nCqnryYoWW4G7DKB0vI4kE2Ks0nAGIdei21VxxeOn3JVC4uJ2H2KYojJuqN45ERI
Bi+iIMyIkTfzr4L5GMqEAchh5xpR8s09r4LEgQ9O77XL0pM0DPeOSI7GjaZNqVMb
+Wt0kHi6/m0nowmt2lp4AkzTOOMRts4g/IOZJIBeA9WeYlRk417mNq/FutFYglKf
ud/KoHE4V+woNQqdOrhunTQ9Zj4epMnQVDL58ZU/nUYTeE4g7BpWThcXxRy1a8n0
e9r9N+9CVk4VJYASDYBZJQMKRqMn+ftQoOOMEpGdSZTiPqMtLJSOJrFCfuRaFm+2
6SxIBCQNo8Ccot3qbkkTD3mc9ZigPW6PtJwNKQZWTZ3FydHeyo5fjJ1MJHBNCgVy
vXGj00CwOKG22DoKUUVlgNSCAthjmc7coVG6vuwVpvadI3tm3H57/ONedNfhOeD3
atl3f2Nzo8s5QLH1rWZHTiwR/smNEyxfB662ioeCodOLvJcFmsMW6wckGY5I9Kb2
2bbAj6Sx0SZWnLUjJ7W7uZvCIPLO55raY9PuUIR9lffCO43ZxBhqwZNRGpz1YR1W
p9Xi2xbR6KUeSL/De04tyNHNxbhdpd02G71ZOGMrsw0Y6vXGiCdjhabBG5HSQOAh
7w06InxbaELyA84cDMxP0w9sQPryQdDIgzk9EHurN7oSFjRIXeYjf2jRUbe+AGre
1g4zz6f5+lD7cvLmqzqU6qLwXS4GCxrDVQegaNfT/We2FweXkvccQXVwk9ASUP91
3wVs82edVMA1MSUzjxmbiMZx76r6Sdl9a6jPsVrXQtae9RedZtDgaVCD+Ud3+PtJ
bo+OdiUGWU6UMdqGpc4UqKy1ur+E5Fo40TBSOnkR/BTjfX3e0VfWJEELEHI58r4b
34s6GN7p+4VqYAtv3gEnZgcw6qzYIKVibGpUs7Ik3s6qGG6ai1NV26QCzbe7g81P
FNmYcCgiJzEWXBI3I2SbyiRLXZKkCYwpUf+k8CsbF+DHgLNLsNIwPcKCzLEpQWFQ
NwvtEY2oP1jd4XujOOE9mbtWeLXIVtenIoZfDJ7+uZAzstoe6LyiGDTvdsk+b8i+
5VjVg7ChXv4zX5FLSvsaVSSiov67IILiJPsV0OoLefl9IAMuWXI8A5LyIJUCaKNv
XALJ3iUENf3VQtVYVgBqhFShg/M6NhH3AJefQBvLrULdhQCYXM/IGFKZTh10xasg
GlQnB1EMgBo5fWSQrtOVu1mBU/0wLvQzF1pS6ifqLttGmvuRTteXECFmz3j+u3bm
0fTjTKn6Jjc2Ibil/8vAn2wcv1PlzokwZRxsgC2xJ611E54LTGQv9BPtHgMITLCO
sHEFI7KWy1TM0XF3oKoVsmV31YMtVfyJVrXdshGH2w0b4asUgGW6hwK/l1V3fXXX
6ECwOdO2FNBiObst0YQ3+pz7pTWdMfbW69JspW0x6Hj96/60T2LuoVlUAl81ny36
NjwUAEL0WafVrs3McWzCl+dejdkzxkoosbLfGyYbt3sIvZxC3OSFsvCUWeWjKXNX
7LPSqaQT61b1ZcIt9W6KJTDeKzSPfmg2ZBeUmeyOAri3eDVxH7wqCnQeKPE8Q2gf
44zgAONJTrFeMbGF4XZI2fvfKOLXnVdGAO4IIY1a25Q3AWS+1GF2tfPghNc4Zes1
9pcZ+nUW6nE1Pl25Z0Y3m4/XAcU/HzuEWVObOYYD8FaZ/+bZfX31P4/OcY00DGqb
JxGDY7T6FJvZcm6Gcq4URxLrirJ5ml8tgMgn2thsE/hf+ExyzFkvu+zeeFtn1Bnr
fRPtPMpqa9Tfo6qe1sFMJvKvrJdxEHOR39sEC3m3uvsyT56JCVhOPUF42BIc8rDA
woTtTqWDbbgMuzEGwoApIyr/IJv+2GNu9qU1CWCHbwGgLkiU6FM3U29FAQqT8nJ3
3vy71nVMOQ1NN9ibqkOY6H7pVuiB3mDMm4oFCUA5WNftn/43qpfNpmNaGeupiXP4
v3XkcC/QTF9opDcH9F+WW7bnZhjLiLaeTWSgvUlurFUJoVx3CEBuAUF2rLk+BemE
13StEfZQMgKobdeusWAsuon99keabrGs1h+Y65SfvKcQHtLLlxwV/mwxLiQ6/mN+
5/7qM+C4cdPy0/7dIokQ6ZzMQWeFQbbuSYRQY1Sh9Gj3LgJLWdE5NkNUh2/nT2xJ
0KO8ab5hB6NKbBcKx6pjgnhCsp2pl7AwkeFGamwdyWyO2WPuK9KVg7qhYpJbz6g1
AsqtpOwtUK77/nxf/ZDSLhKeB0JKVoQS83oYSCEl9itqMLi74PH8APv2ntHb0HN5
c8fSxcW7mRMx5tcGDOQ4k3tncrS2jX933OhEiLswTzD0Kz0qMaJNzA0FT9ntfiRv
D4rKqtmloIqQf04Zngf/o6W7G1ekbY0KcPLPiS/2LGK1oSYl9EFOKg10kQ6zt2tm
X97YBvdGBJNAlvpmKp6pHBtz+UEM2wd3X+fSaLnGkbHzZqAH/8CitNg2Clo2L/Y8
XDFhZUC7WfOi3rRnHQOUGBtosmmbAgDPjdIUu318TLdbZSeRpVtZ3fd3oSRfiQm3
Bjtb6p2VoeWJagkpsMFkHIZefgmeTDgA2A7VQDVWI1/ot2EtW82r+jac/uOBetNn
90V2Io/SlmuvXje9+1h9hoJoGzOdEobeCpwvXnsUTbyaXd1aAt7ia6ShRqif2FhN
h1zomPuCSGVtEIPplXPNhb9Oam7yIhT//ZbxyjVJtCuACgnZGq4RCp+ZU3hHM3x3
mlZwZ9zn3Bw9tea61XhDX0IVhNw+HBguUaykcxWSSeKxls6VJ6pPY28mQx30psfy
JBcyDvhwaevT5v45ENHaSB+CIM3jC85zpv/r079vH7dS5P/C5QcznQv5cPNJAmT8
kjNWq2e27iF0Q8MwXUpp36kFWKnXeJDWaSXXK+Vv0lnoAxcbjSrMbpd5q2dqj7b6
oSA3uwL5j+8JUD+NvE38mMB0zhiS1fObk4keF59JQ4f6iKjmsB6pjCLCNZIc3JRq
F3dnqDeebVfw6Mmyro9GRVI0JJirr80McNx8CNZnyUN2buDeWfx5yhIdEc5TdCi+
D/uNOb4qK6luNLJY0RR9aYZ6tGOQuGD6oHIG1MAl6TMr8lcyWwflHBZwwROqW2l6
+d8dWFVH/eSBI1wRBV+IIRFYWsz2MTRNnQ70iQ2+Ap3T1Xdw/TnGhn6DpGiQbMWK
aMCfITwbv85iH4THZtIyZxB7/NAFbm/Pjn2If2eWwIh/+JwUTTlEMiV8JqwSzEKm
nFGQwbGx31GvE7SvEuiFEMt7rE+Fo0P07fDEy4HmZcuC+2AfYWUjhXbKv/huvpsA
C0vO5jxVr3JkjEPxtCPZSIBP4jjWw4uHsiarQeQF2+ebBwYRbDclm0c6kofa1V1r
o2uaZ1xRsEX4zxq2mbz7+APKrvopwI7K2y1KubqBGKBnI6wzJz5fPhP5RH34NAVj
A7LmGIC8i3kstQFyUoJ98P2so3Gtfnl0sC0213od7weAq28fe6+RutVpZh5gZLVP
tF3lT6pDQ0vpkhL/3/TFjwjXbX1jU+wH/xasspEnx9lZU7OJZwW47pEKwNvrmS9D
pZYXaxhU62zKqVwxVKUwkldnvZCsp4tI1Dqg85GgHkwJEi+dcGwlq0miqId5fLIs
/HvHcsYWhlDDaJUBGbtOWpA8yaIDIN7Nj34c8bafakrnNLiZRnTctKUxei++H37j
6gNMkkAD5hKqIkAEprmHyb05ak0msCFUqchjEvFOE7Gy1arDvBSjNPHVw1HV/e+x
ZrxdIkBzC1Zp8Kb0pXRw6AXqVE9byqMFKuZenIbri8ibBejT3RoJVldHjiz7DneJ
qzziAqPoTLMbjz+Q8RPSLdr1zfmQ12vhEgoYNG0ZoAZgzOANkPhNKp1q9gbM8yh0
TY1UhHKHqSKp0ONCDegsPEOrb1i+Ku1B3POMoM51wJcdRarCvhV3hbNJqCKkuR9a
08jP5FMJ8WLuwG8DXJtCS2/NHsx4pOZ2Kw3ZteoAvyZxBwf2VoFZTkiolyynCPZC
f06A9VQJsgemVYSH00DnaVS5MkUwQORTu2vG1LNhHuOlTEmf8XWupkVEjDO/W6ZT
lYdX7jxaFF4A3RNMtNrbk/1EbVFpofmYzVXPdAtEYrbapl8Cr71PqcY3qH8Jf8vx
uiHkZ0xtb5uRTLrTyWctrTCRdgV27QHH2WlZrUvjmhUWR97Zq+O0Cfm9odo98WFx
JKaA4d0AjfokU12pvB7gtijN5Qhn0oS/43jCXFY8b0ONz/Pt/Nn0alj5dDhJGuZ0
jHXC7rMGYBrc/YU7gqjMxH8CqCMWYjhA76bIuSYMAEwjBT4hyqteoZ7S6HNapc4M
Tkyyj4MNMOX3ZfvdkBtXG1H+5btWLNIskARPzKzovtFNJj4TaT4VoQ5+O7l/l1Wb
Ey0RtY1SpeVadCdqq0RcBgI5CUtxLpNslkUKPLuXYOn9AFkClTlMsjjQDI+pvgtg
GvDmCkchh4bEaCHMJlEeFBmnY7sFEI2VrerLv8t7TnMjTytM9++n104uBmIHwM5P
uVPdVYt92JfCnzGCTe3ygPTUiOzp5x7G4cQetbTpA6p6NBfbVUQMsZoSit4bYGwt
8WGeiRfYGNoem3f5uaSDnMzoAl70zNNWCV5K9M2lAcNIrlbYKQAHnTdTUQWkWBOF
80m553puZFY15SKFjwKg9jSUpAXhfwlfeGKR8IWseRVBmVY8O67O8vj1PGMZEhnk
rqVi3phSSoOz9KEpVV9bQdFpSbcrv9QtgxtNHYp5wM/6qo7bvbHZANB1CE8hUM2R
N0KU2blS/2TI5NyTD5AMYSPq6iXy8UWeHHMG0sFvkZDi1QruGi9T5VytJBuCTD8h
qOPCQ3OXN9pKoOYTMi+F7WvkWGpx//Tt1zQWeCWN4zf5i0XmVUXTxLCGbvjzJpRi
H5HUoabgEevMoGh9DKwzlc6pJSPuJlXQevptOuVStZ+UZuMGkQnnfXjVQjpdu8i4
/o9CjytahHShj4TxolEjXWBR1O23dWTBZ6/PEPeDpV6HFmW3EvZ1eTMbeTAeatz1
YJlVj8E4S9Sgn+Q6xa7mTBC7uunrw71o124abFhso4sLqIq0b7uuwLcwNQr1VTpy
JUEKv6OGqHYj7YNH6kGQR/c9FRJnLylsn8xB0N0N2MNapR3S2OFixaREAOHq78v1
+hCgEdjC0F/n4gcM7oWJbhNbCYM3zlJpCG0BVjjMH6TreW5fYbKiG5qVOegynPSj
KV99Rwxd9tQWwtDq+Se59IxzHlf50Ma+Y1fM769ZtzOlZvlBIiYkCbE8VxTY/36s
7cgcdQUJkorr/eMzOskOFbWC7aliHsqXmxPKyS/7GBIR4B1sZknunY4vMnVwVNBY
Raz4OUjeYOh06tx/Bzy0E7TtEZAHsR9R9GjiYcHwyQ4dGfbktfeskU1/pY0hQOaR
LCOl+cYpPxBI/D2WRUWIYFpO9p1lMCgd5g5PwU/Rf31DhTEotubV1Yf0EhqaXcEV
8MClMOW2FCuaiAdKu/10TfdEB752G734/IyCVa65A+riFnDvrWaE+zCSyQLDSiq+
vIhlIMdzHGj5XdJY1iSEQA3didJ9IBiJRidt5U2ORURtzdB18g6XqXZX87B6rq11
cFOkn7z8UlPV8RVSfdzNpqUqwX8ElpIIGTL+ql7qSPhvHjLAhXRBhQa3zpKoEYlI
qkqI1HxTYvxZBLUfVJE+BbHuC61YwyIE8I9oTaDSMa+2+UCUlVcq8qGHDNP+Gl05
kPvpvCOOkXu+PSsSwtFZix+fkEwOw5R6TOKBxD1fd4ssSGAE9r2IX/MCgBZY4qzi
fOyNOBq7JAXOIOh/+oI+okRkujQqzkyaVBe7Glwdk/CZ9l04aPAOrsV/lqr5y2PD
0B1jDydMBwhZEJ268a+DaESSNzlu70L0W/Idfcs0Fj05LsKyPFUpLF+nJoBQQfK+
p1QTXJk2lQTy2QStUdn6a2V1XyFgD8pv/CbxrWkcCNIxu841usQNA6pw2Y6bLG66
08bwpXf6x54h2UaIaU3V0kuYViOImvdQ0qRYUDIOdYmTZ44M3X3r3TU8tubQC1Q5
BsJl2ijeQbzbU1YXItE8Z+A1IZi3+iWQg4b5NFASMuc2eX6Be5VpaiWOX+TnXbd6
F9o42Pe92GXGFdGa0gyOmet48MRyFGxXdrNtyOT/nHTLyukzgVcxCKxhOzf+JTTC
RzeqSLHcnDjcWLQOfpsschAdSIGN1e+cbzlx2hgHsfF2qlzy486EOyKjnhtFtEIi
i3FMwf450Ubgui0qRRcJq2sLKJilZ1hUjpK5PNRDR7OhaU1ffIGP1QBWLKeKX/1f
nmY8kDppPneKBu1ZTk1TDNMM2UjZlILHR2+mglBK3r9IiLFVN972KXSN5XP/maIm
F0bgoH1C1wH898d6ZW2w1EXVAjDVgt/7UUviLz05dk+nlZEqbqfJhRPNddYcKqLL
dZpFeRx6zIqAxi0t5BW77BnUrhvlG89YhPCB0MpsVqXrmfjGfKQMXjy1IjHdG60u
O3iYAKxLjqCh2A3LwEXkzCvb6Bu7/ZY5z7KK7hzXHGyC3NUXspNZ9o8FKhzewqlA
ri6y7/ukrE7Mms2MnWNw2kBB3dSNw2+KI/dDt8am9HwkKrkNfBqEY6sYiiUdBtGh
mLe49etfMibHhpoF1ZavrrcFf4Io4eBEyebGiPSe/NhkRcofQlbyvXFpnSxnrO5y
VDj9KDZb9ixTEfyBXEkQvKpYwPsukzejBlCC1XGIbl2vbmv7vxWI4473SVQ+tten
eEZEjlYnb/bdS3KG9PXt+67cbAMKQDe5edblOI005DjyXyeH06xMKUwwXEXMWT8N
QY6xm6jOOPoJhY++dQmInMY6G6pOmS2spWLDdIPs7zz6aG+ECo5OZNbvfnyq6n/j
7rai1V3oALs1fNOxVHJzF4gM4+A3Biqwn2zXmNAws5A12E8R44r+2YXOcLEz+w9p
BX671T3VKGE3NSAU4P64sIo429vMEh2Nca7RYhH/lUv4imfuGCu1gxexS5wIGZMi
U6ONfjq2FhdHjWw2PmTGgd0f7AjS2pYJ/TwBiPY7rQE7w1abEM8LmX6JFbGf3VzM
ixZNM9BzRgcUhn8Vs05UlRZtOocUcFp0cU/wbUhd3kanHFQ2NWefsxvWiSrQXxxu
Y8rfvaRF8i602KnOW3he9bLLpiMkrnv9Ib73hxYdqHpZQ8kMzWFwipQc6pKYfWnN
2fEaZDAr0JxQP+7LU4rzUfBDEipSZcSGW5OrBJxe5ND0GUOUWW1p1dD4GGd16uUA
jTuIsFer415qHtXRkXMeJenHJbUghLCksvJ1/PNvxsSEnICLE2UZgC7w6kcVpnii
PDElDIzHsptV0cNd2G8KUe0HaUqYu4I1b2HeXPSTLml8xjk0L1aDEXXLrpsw/5BZ
LPQcGPZZV+kyeeZIqzlksU6aACu42L/ZPVrMNF4lZMjBBifY2niItp94YDLA4Ksn
3tWWM2rxgBlG7lVBhVcE5HaEcuCtGcLY7wRhMIiotJRQ62SlSqWDfPRAUgxmETMf
lKy8kngUwRacBnA7UO6UDjdnrYGU8DzBSKazIHLcGacjhi6LfBZmc3dvtcJzbXtr
wTW5+0QELWBOf93k72ZAfOUIBZMlfrGNP8SvAI5cK0pfAKxZhRsMlJ6mr0lhZABY
KoNPo84G4deoSg1DIkUzSb7PK8gT0cz5NgY6r+23CFPK+WPZVcu/FVnEuc7AGpPo
H3dmz5r6oQEwr6tK+eE1eQf0lgWK5Jvkro0+vpTHO2gjVynKcU3ctSdOGyZsdzYH
ddupJru4qjIgo5i4fProslMED/LAL4iVjAaQ0BiNcf944DCP7+9EHHhSkKvW9Zyl
vdo1OCDA/nprmTx54/n2OadJ2qsAVq7ECGROsg4DGegLoIgrGRFdoYODiImk8ebG
DQX0CWYn0IiP7kw9rOhNtdFUb25EjYW/OmO+o9lOzRjd++F06wEn/XK6bpPRkj1Y
3CjN7rz4KT9s31WUwmop5aBGZGmYfWXWXBy0rdN5qu5fgxbf1/fD1nBXsLC4/jyi
JTmnSjmCviDON4IeRr9PUNyS1wP22OtYaRj09X1lfhfVPX9rDuX6HskpVlUKXnJd
p0VIFYddBTRFwoKsD15/Ikf+6CEDd6QgqpyTuq19ty+Vd7z764my8iPI41Iyxdn9
PdoUJFd9Gw0eOLiLHYygs2ZJJ3MhjBS8jfR2dLJO9zPyXFb2AzOdrf/ZuKtWXYLh
S3qJSeQi+aSJ6CQa2gPlBKculORyci/ZKUiAROdUVMMKiaGpLqehBIyMty8JDwfV
nMd2P+ZXDZztB1CikZTcEu0kx/x+et6FJI3Q00ZBlMZG+UUtZEzJd/XZLYYy3mrJ
Fb9tFAPRYo3LUg3yfInA01JVhsUpRRq4ov6G7x11k0ZOcqJ2jMZTNYPdamSZmeAJ
dpJfAjU8hP7cb+VAHTy7vddt59ziR3rvC0WeYPubJKFUlMU6xcJTVcZhBqHCEpK4
og7RNBWDem/2EkwFrRv3h6e4LFd/1s44udoA77/Njeimyl/dmld/3PTf5nXhVfbP
2xpDuc2a3pJbsiLdMkB3V8rqYAhAXAYZ5QUAbuq6wLr0RwrZdI6kY31XBFTKsPVb
1R+FvFtxIjXcN8xquiaHIp96RGWKL+oDFEv1lRrdBAdqYiC9NzTNtoQ2DUu9FodK
LsdWiyZZ//Zx5UyYX6DUsPXEZcdPCfzyHn3SiZv9h+YozcNSMT+PAUzqhyFoMmGO
8ZVpjLdtlwqyYzXqHYklA7tV/CAsqCqm0sfEoKNqAtigRKSrnf4TePBMG96NxZk8
Bw+Nc1D3Q5pDuDnMwvtPbL3MlyQRyKOHOS9lQ8HMxAMKlIeU2/20c25nguLbEdNK
+J8pyiFSo6tB1IbaGTdVepybLNYXXd2fGtPpud6Pf/i3z5ygDWCjDGTcIjMGJl6c
r97gWy4H9x1FKzaN5uuanAjD2wpdB/DvOj0GTptffKkb8JIOzooTAgfIOb//UPEG
xCHgCuuBUkjG4bRyYCs7SZCZgNhBXjlT67apiAXRI43fwerZqc0JimrKauJ09+/T
oryMzEXB+K32osvLvNJ+HmSQbB1ypf9SThuyVkdqnSvz7yFVEOJvfEC/hmvcP4dO
9qK2lk/Hks5GvKFCZNnFJHVdH+fkBhKOh5fsGMpZegLs3ZS564X83+Qf+UADoFaA
XhFrpylAt7ZV7QwM9SBjWeoOU+1SXNeNzgOs2zN+ExOjwSDArzpGwddjU/NGzJ23
shslfa7v64Q5I0TTMRVOE4V3Cz69UeRWrjJhn1xiaZjHKefYfBpRltOjYr+S5t/n
8mwr9Mns4DLCm0RXncpHg59W80BTTGG05TsRpAP0cHYrj4tiS7kTghlZRTS8tcLt
3jBX8F2Vv6ma7pKtMCjRpcVknyKzl+trCI6ybpbfofOnNtwRGX0mD/Fbel7p/mb7
aGGHr/cnI2AeEyQZ2s6AW7Vh+Ihbr9sOE7v1lL/K60WnIsx73jQ61XQZ6+umuloK
NcJC8cBn67WYvYIEUSRCnC1QQYNfDMrkuFgXVu1m7TWEmqTKPm3w0OOsJpYIeapq
gpmEiN7Np5uiXHz4XRFkpLd+XnXQfQQOeX2Jw0hn5J3u6RXJBGrZil32v0HL4iXV
t/eLkPQ7d7ADV6E2AaVkp8IKA0gvo8VQ6zStsa64Q8XTSZddDdum4PB5VZpkA+Ik
UNk3t+OdxsVJNp+4j5uIkh9BQiOed7a4NDEBOBjKCgkXVLMLmqyeyVKK2Kp1EK2c
mZGaJGJzVlYT+jJ5RKKY4DoDgkqZ2fOlCIW8W1N4hLxVzHF/aLyDVOhMtpw5GwxM
xAl5uROX2gsM/Mcsgu2rVQc9ljJJAIM6QlnLJsiFoV4NV+v+qXsNc3SqBRBbN2rz
V3HYGUOG3KlgDO6Q+MC4zWgeFfgZ/V8DxZkii7ofgNe7eihVn5Ny9XdSOeSesfp6
+n37QmGGQ0MNvNNhT0OcWNwUmL+h++qDdGZAkvMAq/5l95I/YdPrhy7ILllcGkVE
x17u4tv5kcaLrr2pJPMb1BBEkBO5cfN9sD0OseLYfrj9dugtk0swm+ssmXjGrPFV
tOYz2cDw8V5iFRYGkg/lrm/TqVUPg3VFY6Pjzc5qOA82SlSNZaafCHE/PYCLb/DX
ATXNIuA+V8cvTvJSj6gKjU+pf+5RUzYUICQJoBZPfcwTXte5z+40oPQPo/x5TgWL
62PFMn409XZ1ONbdQv0udAu6AVaSsVulGmCJY87SO1ghObKRgrD30sDmQCjO3V0K
9n+xcht7WJ6AU8SaBEjsiZkU0ZX0BqyJocUMk+vnlcLkeZnquIG0GkURsgxlorQD
U9hXKNFZOQeB7Vlcgy3siuZyPS+58X55Z9ytFBFSrPucZwDgWfU9/olCywicQ8y1
sBqOP1mkDFUv7bx6KhcJZLiDjd6UjZ2cKewzSRVUsz7AQ5AiLH0/Dmu1eU2DVCa0
lhGESRMOk7bJSaD4SSIJn3pi/ZAldKa/AuD2yq5AuHai7KFo2imspn/5hc0QfR5e
x8Xr8E8JzMq0Ql8m3YEkXSxoEPKiZbf6jsrRMnKSPfA2AkDVThDwqNs4Z9GGZJSm
Wikt2kVob42XUCDhepQbSXb0TOb1EFxAptFNOFKPsmwnQWtqWmRkp+WYduO4NJXr
uUL/pRCnRSxFjCtY6lOq2b8NEz6QbAzAPyGNOW/phw1a0R3pWR2QYy9LHiwJyZ9J
kLIomKwbpVdh9XPTSL7o8o7sUCUxkL799wR2iENoUKqu2CiWK0QuiyWgzlijjDuO
CltR4HQQplna7UpKmEMZyu6ufPkwyyIvEcAI7Ix8VLYDPzlA6wpdA9wAY1v0mqU8
Hoga+QdJa1zPsNbGy9EI201yxu/c0xi6bPP/+MM1wuBTCc9pRb06ECF3qqSeYPEO
8lBtwChU5lwvHwmybQWwU5GTjxXuM1z8kM7UQ/nRGMw282FW28RgnvagVi0BQjTo
uNj9D126hUuFXYSx5L/i5beYG+6Jh+RwDd6To4dLPg4cJXDuxPb0hZC6x17JIb8H
DpJ+6g1pyo+26o4XC00lZzT56XZlLgoUhQ0JlPzXIEO3QoSWiArfzBm4TNp459HQ
EK9hUohstt1jIiC60ErAUaiwZZAFAghVxI2JzQ4ZF5+wrBa3BEwkKqs92Rpf1cKW
GDmWPGx3SPhDIrqNE1ahWS7vSFNe9WoGTK56ox1jOn5wFCQWUtpLWjjAxV8WGiiF
sZ2/vRYX4QyHgxZnnqtrN971M0LHkofWlZABmDcGm7kT3FHMWBp63mQONlwv00ka
UrRK+UlHaJjhDPtya/kfbmNs45sM8YHvYf6bHJFBZ2VdtV75d+NmjL9TEUAnD7b/
NP+xRmIaz/vf0tn7oo1tOsWGGXKTrK7v4KGVQEmOGxpDicBWxNl9Qbohm0/51TKB
GTtp4tsujGmnog8vsbsiB8G8y6YvFFEJbpY/VbrvDdB/abOP1txyqHbTPdp2dqVD
oGTAjon0Y2A4a/gr8NMvuJqE4pyFxcx/turKEIr7wqauftLEQXfn+ULyD16mUJgo
DMzPo47/+W3nSYZqDpGVHo1VwAcg/czfvKf8R8VD6JYOdkuV1H7g4xp8gqOD4bhB
uuNmeVJRz/9DjGLdFfff4eA8LJ5PKFWsDCohsxvS4I50HEWUu9VFeP6mLb3rV66s
9CH1040n/CxsKcKuuBZa/TVnz8GzkrqP3B6l69j8t2+4gh0YF6MCL+R4IE7WAfe+
/8p3fKZE6TbdyWCQVRy5kTwny4sZlAj4gWBHQN2ZgVYzmZT6cu9016G7tyTcndfi
eq1dkA8P10wlZuO6dSSiO2Qk8mUA12Et83Nd9yXQLip0Cbes1jlj6ib/CUnwbuSo
VjVdG0NolIfltu0fI30DXSWjRbw/v3/gQnVfLpU0X0JtDp8kBsbzJiroyRtm/zKf
5ytluw+buuxrBvjxZ1dxI5cvx01QZkeNDlHtsLycY/h6nS0PF4w0LduDIhU92o+N
q3THzF/7K5hrvV+KUe1wB5xb3pOa/IgZjPWaYH+ZWxFvVnz2exR/YCYIRQ0aOIng
mzxAcr3JLMqMNyUkatTDzQyaJ+1q8WeATOjDdrUSjZLCBO0wEJDTjBzh3GLabZGI
UkrOsrnuG1kXAQsl/wdAxlH7wro719QH05kyyh0WtqIutECx7qaN2INI6TjfUJFX
1vq9Zv404p8g5CPlV0mm9/9D6pEyzzvFV7KtkXdweMhIh3QN0rYXW8AqhDIq9KSV
OitLORH9Y+X9ixBLJ0UYkP3HFWX6NxeAoIXfg/GYe8RmQ/bMxzMSa4O31HmhoNvC
eSmS7KJkUYonw+h9KJENnr1Elh/N6h5B0O5sCMHTjP0ZUMEQVvvyCPBnufNMFcsz
YP+XyLyFHDt6bG0CrlpakK5rwvQK5FiOmAEfWQeXknko1xS2amQS4E2GYqLyVhAW
Hi+LxWJJJ3I8E23NaBgrfu234Ufum5mEEJiaw/8gb24jjThPHWAUyAurl4XBuShl
cEuQIQHf9YvKx2Up7exHSHT1pDw7vQn5QGRe2fLmomSN6FXRCMtG/zlQVi7r7dr6
Lz/QdMY/l5xPvODWNZbQTsfIHgHYtvClEslZ58t8x1uQxrcLMCXBUKU541raOO4b
rxeyfIz9gOD+JMTNxhq2YDCK6RMCPKF/U22AkH3yWQn08ntrWaZQJRvdV9u4g5Tf
f6GE3TZ5hcdTjU77ie5624BttmpPzKHa2BAhRHBBWRbFPs+Ly5piklWBnTHtDXUs
lakjV99+VoiwvTBGkwPVW+32jVMK2Y/J/zyaQcDohZZt4CSwq8tYZUFjbmLUk517
QyqGdWStF70TvdT8q9k+0acCmE47pLSsIxL67E3DgW7PX63BvnzpNPs4v2PxX14D
PKS0GNCOq792VRX5lrDyf0J9JI59AaxI0FtuN1pR3PxHGLplDAjTA/0l4OwpmyJw
1AzmE4OVXQyxhJma9/w6dAhJosDd0qXKdgHgyvoetO0M0T1xJxKtK5viar5ErnOk
oFwrsO8yBGKBKVNFcPoT+vSa2daVfmEXDZr57u/42dbrU/KcHrkBu22E1gUURnhw
9jpqbCmEqF9vubL+MPwjDoZmpUBs7UzOjMuaC6ALdVO0mmOoxPVA3Rc/FSAGqub8
yoeN6YfVSTvx+XBlyhR+vBbMx4WZCDN4bqwSVCCa/p5K6AgI161oL+d4RDoORnPs
iVcD89PpnnwbR+CV9KKhhG6LBu0cdB22ESjRadjQJC4IWVGRr5yns0mEPeuTT5oX
d8dxuQ26YFKcWEl03ssGdNNCeloZ1mGrlXWmG0gRC11gGuExX7LEwjfcuOu+0oSU
SkkhE+luSiLCvIKcSYY6cR5ieQGM84HQottChvfAMbSmUhKmP9mrYtQjPrszOsX7
CkszvRLge8zfu7+ZTvwCQ676mwJkcBtxao5zmGx/KK8h6oM1QjNh4oW3KV+mx6Za
W/KI8++RudS050qnI8EPpaFpxaBeTluA4DOHju9MQpZ53LJAtzCJoqxEs+JPGBqa
R6T4h/dfnzAYkRe79pzOJXkTi26WGQYtavmpdh2HV7nUkBR1Vl9Nc0TZARUZohEg
BnV58JHsZplaQbkAO49lPB9IJbdgZiq4GJUMD1Nva1oMCt83OBQB+LoAOBFxzTrM
GBV/diwRS0rpsdjlqozwbhQgSG2vexQnj2oSZDYAWSD2H1O2EchnFBFbjRiUAXiY
EQxZJZpdb34SUZ69ZShVPV7Fs1dsRpR85FLJFTprHHhj8sbcDSYHLrD1Sb600Slm
O0rolpFzbOjJDjKwONnjcJ9dwnUPhERU5A+AHLv4tFPZriROz0rpN/8pZsHY7zXD
ic/RIsjh2YBG+3O+OzE+cjBW0uMr4C7V4g6zhMq7PBu0efq64Ikr/Ai2X4x2zqrK
dTz48EDkDOxtmrBestOPMTJ/MA3qRwywERLOebDTStkTe2sxhcxouS3GGAdkjO/L
jvBeUSp5CDnk6nFPk8OcvCkjhG4Srcii03K3noDcPU8rNV8vOBvrLn0AYERXPCV9
4cKr+VpBseTGF4s/QlFqmO73rC0GSKAYooSzGIiP2DMGldHj6S2rAW3h9HnitUXn
6PqR/Yp+4x6Q9pGh/5/VuLcx7iH5IvmJCgmlrvlfqbILLoGsLJasuzCo7S3PgOoB
EVd0qg9NApDZBu9r34J7d2EEj6q4U2sCwF+VzXpsaur1vS7Y4RYErgLTogq1oXXQ
IMjgwolxHQY09g1d2Ihx4MbVJcNhJ+Ia+NW7EkGhTiFVNqGAuE98mn+jDs6xuziq
a9WxlFHoy9uatISMDGoFYg/qJ6cLvHP1ss0HY082VFfiuc2uoeUDRX1iz7NC5VB8
YO8s32/RlIuP1DRpjcueOBfWYfvAX9o8cn/IPah6sEGV0GmSJLj5w/kYyNFySMc9
+tiecoPqhOtm0pRR66ir9Iw9AX6tKAGOOUf7fVrUP+EQBdC0CTzewW+YOMK8C59K
7A32MM8SWl4cgM1gUU0SUIu+zRUH4nk/gX7GOrN8fZNS6deedk/H+6plaNpvICRZ
cfX3xhFme+kvpk0l3HAsfcCbI9LkoIYvNu8WhWXGcpjwLM7vkcugI2qaMCGU74jK
nJr7dbOYM/dT9gKs3hNbKqZ6T2qitR5ganX7HMQQwVu22kg6Yeq70oBOnbdzB2in
SW76UKbBTb+eRWgrTWnMHoiK2IP5T8X9NV4+LqQdqpuO4rFrvNF/Sede7cXqDH3a
zAdAWCiRrfyV7HUHMV2dP/jI454XL8qod56Mu3teBu4sRSiQo/NavjBG2n3vAJIk
FZpJeYIzM3EQYdL9D0JWTXec0ywb5WJCu/si0X/Yelo1xurIRvht/qNw55Y4MJIA
wzhFtevfpQupwWgScEenSoLP1wBptVCnILrJNAq7N79okdAAmE8Dr8hXWsZlgpp4
G9S2RT+V0nCY1nE4Yp0nmv4Cl7ilQvdrpuZCn7AcQnbCHBVWte0iBDlgqBibn4nO
kpGC91HAyDJWs9w7pOvJfzKjIPUy00S3X77nDH1aFB/njRcc3UnuhVYTRcexmHG2
NY5LLTyL1/Drm4b3G6P+VdHQg1mTD8PFlqNAzaGxT0RZBRbywML+CGo7LrGsEUwr
qbkMUJYZHwMIqv9ClvPxO1vHZo5iQltFcd7a6mWI5prnPjZmDcHGyFRfHBsltod8
B5X75r/WHMMEFiiA1gpFuG29wwp300BOFMdPXIgLi/NiR1KIAkac2fCywLTphJRY
fZjQ56PuuDjzf3dfdEM+u5V1WEQ+gmEMISa90KMNoSUt9wljIcUNNF4G0srMSxfh
jvNDp5rX5Rh1siXKbz01w18hgf+3kaFYBNrQfZbuPLRQWUq2yFCVdpZj5PUGpnkO
B4Afmt91vDvzIn3wRDYAA3/LeRbDUUu9llT6IWCCc+tnEWRfZLtGNc3G99/oGhE4
ZQUmw34XhA1Vvm1e8A5y5kikXkEXr4qtOAgW/OBBkWtAU9NIEZOzgYY3F+BSE4wu
49pMJkW9Vo0x91pEswGqfS/Z/iYDjChBwJ/ktQevji0Mf97rZDS2n47LeHK4mOHI
hyrg26WZ40JEHLIEdojVQExW4hmcf1gCmi5c1cMaCre59Ffix70g2cBbOXaoZq/e
J7m083zIGoFSPkwQ6mUgStUz2SogUbynU8YeE2UAWSLnHpBmpHR9gzPFQpnbgQeZ
mmCCqvopWIPkwHSctdnd5GNoq2Z7zOCOrLCjow2AnE8/1Uoo2ox/+TcgXJzlsI/K
U98wHmVDGrVb+7bD8JXMD6xZOaf++mYW0MubHGsso4kOyzDA5z1ac+XDTLjCfZ5W
c46bjURhiuUd9o+OKKLzoqfDghGrR1b5dGiwmebxbAXSLTObbo7W3kN1QAPell4L
wbByo4RQsze/JnwCsTYxIJllScISdO+9gVrmFziCBfrOq1K4acofJboS5a3Y2vzx
6LHqutp7PBuZms4oD5NENjGPgtzOAYZV8Jx/b/+ayYYOxEBzPAR5vED6nL9rrPOa
nMo7qhtb7gn6BqsqBMrevqxwSF7jH9sVpmAOdFa6yKR/uFx+RhDSxvtO8ZOOuGOh
8jSKzyzyY7dnIkenKCMZYl8tULCDxmo/GFytX1j+434ZeiTwRh0D4LTND/edxS0q
tlVjMvjYwxwYCO608CRjP3IhQPXYPm9YoiRofcZvgP7S14CFdffdrcmy0Ej2vHqo
Hw19IXCXC/04osMZoUzHVcoNWMpntNjDe8oQc76UnaHY7e55lP4rYIIpeJ7E28rl
vpgWTmkogf+rYLnPaiPiFWoYWDuEg4pfIj/976CkHX+klMxykEmxnfPYxatijwnN
/jvZ0t1D/yEJnloNHGd79TsuZ66UHGk4RmGPSPWUpmXfh19vKju09j+HdUtOcSBl
ZGVQM/dht3+IRq8XDWg4leky72Hu/RNKhz/hoZ0lt3JklDIHaBDxlvH310aLPzrY
mk5HMMaywwKHkBORJBxMo9LC3HDjh50q5De8LmC94ab+gIAZyYc8z3FO5PP+J0eZ
V0MYUrTYk2OaRyroxAdWO3edOMtJAnfYQ/EhZ+chDLHLCX36TIABuMZTaJ7H0uQP
bjqcuM/CjgHRQalVfcSQmog6+ymTUKlmt2ed5W6VmFtmSTW9LDtZqSeacf3k6U+/
3/TnIw4/loXKRrSlyl1G5HjtojxqCOo9a+XQrSG0ZEM7l1LhDFCTnhVVVbenLq+a
0PWLPRcV15vUQlw5dTi8IPbHc2zuxchEB5NqiolIUJHiTdrUJsj6QDsDjlf1WmZa
l/6DBIpiA+832I2dfc/AxwKY6oRvcrjwlU3NZhdkUM0gVdTxwbX9u4v+OJ4MXqLX
tFQQEA89goXLx7ZqTRhey59HKZ/RDcxto2xQzMac1sXvP1FChWvrt4vNhRc/IM5E
N292zBV8bM1yLG4b8T1dmlkijjy2+z3cgY3ono/NV3eeM+9+G1cSophwp4Bneyqv
d30JXq/AWVZF+olAHSsdXuK+PDzOhx+hIBA8+P9uyUlvNBtr82eqb33NdOqXvqWL
gLm7MglCNWdA8rckjh7DdXLnPpZqHaJEtXVV8lf8h2gVXBijzV3YWyVdfNIZJ08S
rG+zyuqAO+TncUu5wYTLwDKYEYiu/dT7oo8m94I/DDrkNaPdHLhPYNiLvCa04OWH
F/pjqOAahJd2pcE1XMZxfi41C5/WF53sHT7IrEBJQ2Ciw5SVqbSYNKupa4VgkeNZ
Pl/2t9eA6TgWpN/thVg3+I2qmdQxh27JYO9pIms/t01h1BHBEBspgNidncVwBgw2
sPhOqffK55E3zbq3N+JVvQdp+aaLshBi/oKygfJSnGFVtsuqR4F9ogE332xyvFiY
a4C4sUI1pN1YzcLzHizc7zWaOlE4lT+jaJjg2NHiu7RBfgzOwTpJ6FFVLtsLLCDL
G8adqawNyD4u28NGWOFwOZEjHu+HMhL4vm6n70aIniXmwbBA7DaDrANKySLnSsk0
Yhl6n9PGk3jMpzK8xma0KHaxYxvT9w+CXMpT+oBasRdecl3tFn8H9KDO6LVVp9FY
iPsrROUdSeE3epErHcdSgUR8jsd8fIQ5sYKgWEhczgB4SZRivxabDjvdSLIPeAK9
JvJ+kv/qvr/5csASvLm94cOn34DWDSqPkymHobsAZyTtgE6POrOovvpNSkuyyLvW
LXXKbRMjjswR6mJrAHZ7Ha3URl8g/dseSnEkB0spBNEs9YGjUgOQT+YC91Gj2W8K
0b6fe3hhtJHPZvgnVSF04y88zjirt+SS5p4Y+blFYjPgMnslLGpig72VBjqJDh9q
BU74WklVPpEDIPS/kuB6J2BigB/8RnUlyUTQEqTSpDIhzD+dlRRO+2/jWmllcZoL
DB3QP9wo7obgUxnRcuV0g2Ln8zMpJ0qmT5OVZz9VZSb2SVegcdNGLN3FSIOifoN+
Ps97kq1Bg3VZ+S1VnWBE6sLaqa/7nydpdRly9mCpNCwNL998LY0lwFPhhII0DmVK
AouU72qH32Fs/BdRgCG3B0MH6FgGahHYDyx77I/oNYgn1xBfPyXAkcMKpT7nTvZU
K85wd6JCfUevLnBGOzMWonafTRVrYkwJk6rKCCrHj+LfXwa0cWn67wmrkYD5ZaS0
KQ2I+QRj3CHyBa5mFNjau+ZUAUxRzfREA0Fj90N4kn75k+DlRl6YKUP35+B0e4RF
qSJMmkrF10JVUYdSB75VsF5tQKNqwOTSUbgAg+XnpNvJ8BrLhEcFWuuJPkd426bM
pIwe2qWkT1zDUgHsjAxiHD89WI70YcCA8JjXkY7DKT4/tpinR5qOs6rvKp3d6gXD
EE9Axyv+5w7XQQwnblnTJqic6xVzoAiJanLACo/BoAyzvM1tg2yIQs9OsN95HcEe
vzI5vi/QCvNmyO3Gr9H2YvGA/79VyEkj5PSQL35tcDuTDEpwmLEPa/7nnRlwqlsG
7zwoIowMd5x0NkhyKoCoAu3VzyfcRwVwU73K31ugckXJIDw9bRp2aSIZ21u9L13k
cQo6fJUHiiqSjAOyyJgPEMh11VlF9vcIOAIIKwR7/X6Iz6OGUcwN6jAEYc//WalE
jvB02/ciH3pVGysLKztNDUATOMbBwGsQypAEPO0peg/PAZ/kKcdZroXzNwpKzEDq
SPiCLBi/0unc2lAXzMLK2Am+HpcRsGq8szICxSKa56Tv+cX9xip6M8CsmfgOQLJN
gL8IhOm3LpWDmwIm8j59PgBd0xxLQAWaqbN9BDMraePRM8AgHUsOCpCKbU2y6lxE
2rtsSC4aue84RQXr+rZwj1xm0OBpRrdrNBGNiKilLMC5XijlYFqQqPTLpOQYktPf
S0+2Na0OxEn+PIbyhk3rN+yjIrKh/owSj2aqoZqEUIvmAdyLWFWF1Lg8EBauPAL3
JugBYFPaNx0BDXqvGPDleA/Mc+5zY1BCbN8ErviIqHeKjxmOAF2g32kPuLq4Mho6
K88TekwqLPHegl+20JSAefNPbjaGvZTQnPDsyawhCnAVsvKYVmK2RNmaY+5hgaLJ
VDdhM6x7E+SY8PbLZhjDfZsX50FCpxR93BX2jYVck1OcPrWEtZreP1G53ULSRpRj
SW02vg/IWoHDZ4VY4tU3iqJrWks1tuRBOGCKsZakld3mTX0lU0lGzhyn2deD5JF1
SnVtL3ZXBUAapI+IE/ax8ayc1nAX99sqS6pUjOAT8FOBzI1eYi5KrelsmOgzTeiI
ctnHSc56bwPRj16YY3g1pgS3JoqberrGrhWcrXGK8k/eK2+jmmPs2F8xc/0HHIFC
LglFA+Gzfsjc9itbNJiyLTmc1/sAmibKjei7WjfvTCDT1GYh0TgmDstfUWhW8wo7
OZsYiNILGxoyN28gDIWs123Tj0TMGMCVBGgcmqhu8J9gwCRb7SVv5s6fUx7vwJOB
dZYT4hRH7NTYkBKaHogv8LA+ab4zFx8udiokzxraN+7z2C8kbnC2JJT9Jhy5C/dh
Yh6Ee3qfbi3tY9loy0A2WrorarofcQlQ8g2lIGgKDpsUz+DFLw3ySR3aD7vfYCfA
7JBYrnaA0V4yD8kNsdh9kyFj3UYxZfQQ0FLR5Tsp5WAll1e/ycW4MVKOIMs1sfk5
ldRg/gBJEl4aVCa+eVBcTSYXWSpo8tsBiXaWr1KaKSEkBww1xVFuuAUaqMOs1Xrg
7Jr41yB0wt6u+S68ZfvegFk3Bb4sSdAqIkU8IT1GM+TLN76Ot7SE934gNgP6wzqQ
avcnwx9hfqDJ8lHtc7NZvYFiuh0ZhQ6p7b4Q5zMejyFl8+6UpiDjMPOuUkVK9rer
+csk6uttzb+tpcnGd6YxE8VwWM/TvJkCzpYjnX2sKSPjp50fB1sGk4h+VSoB14ei
NhpPx7x2sUbm6zoF5NrLovhmVz/5H+Evj5fqVj7D+B1o5pfIl6s67rp2WeQcKvnC
07veBCUMQvBduH8auYEeZfhXQRvPA8FyiuvgBVkMMXjKUp/gv8TXqJNgEWRQY+R1
biao40ln1SJkPq/CR+ZMiL8s9MScT74rzWiMpglxEN3UYP/2IqO54mZuMbPg10gO
RDEG0MpSLrAs6PSZ5ia1hDhvjeOMqk5ZtEzrYSvH1mfDZNjGS16FEGOHnTYiwC4j
6YKyrDxRSLMTYs7pe71uZx8a1fZ9U5YNHIl0ki+2oAvtK7tScUUD0iE3d6L107Qv
dNR1cD3myuVgmsn1xLm7bEFODFdOWRc2UfDboEWv7qsXHDKpcfI0vidkEfzghi7g
4fVi8RC9Py6Ckl67sdI7sL5PYrF4LaklZdauCWSsHXtkb/pbs1/kidxwM+iNoAYe
wPZdeUARih8RxV6vvU1t6pLX8XShOsWj5eg6XojKQie0b50qKJS5RPhe9uneX/nH
VwzmSCYzLkzeDSoYItYPKUaerrJ2BL1/A8AmWnSXaJITqDMn7KpOjiU7anRFsPKo
IUwYjOXqbh+ui7RDW5WXsa6akaW6GrWKo9J4IThn++88EcsNTIyhSSkmm2ye5WTT
PDNzaxkVXU1/ESt4qUHtjUruVOujL9Dikl/oNkZ6y9xVuOKWbYIyB2BCeb8zSnya
sD1zoaMfDRqYC6bGly0y/HyKrZ9pZYUMaJfVerzcO+cpqYLlbfDGS0ox30Q0kd8M
O1sgB7HnlxIHkJZwHGBLVDAe6LgryY4DSlm64u/hH/QFKZ8nm04iXhT5fVLNPY+X
qgcBa7ZdCjE4Nrn8hqqUGOZ/EDFYS6KtjnnVP08FUOLtRPpSMM3J+IoJjOP0qOuq
mBvFBNgJwKLikT+DmS4vsYSRxPfp3EEI7c+VWLTmfd9HwlDLK8q4jp9iWWR883H2
kredsqnN8yXCGCyg1/ksp2x+Uiax1TUF3SM0IsbIRBFDTVSLFbMzrCojxHTvmX7f
laG/C2/Z/+dfXf7lTLdfOR4bIpV5PaymiI1DcMANtF+sJdXnaXgjLlMjIS06EURJ
iKi9EnA5spuLR6AIn3/zKUJZvRBDg14cguVuL+pyY+9Vp8+bzpul0kNAEZli5ODj
d09OKM5SGIlPfCugkE0JO5HbUO5GblMKr83g0PS1Uq/A0EOB0x5pzyzrd8SFgkAr
j86fhLxBhX4r4c4xuXvbcMRd286R8La5Idd1LTMy73mv3GqO0Vtpa7k9i2N52QOr
QXhb0cPyr4iuQPVomH4yyfyZmNjestYJYTUoZYKGD9H+amWxTUiQ6H5q+Z/EdyIK
S1QNygQ761B93eW8wa0O/5wT16auid+0NLQiGbIGziiv/dKNY6+IWTwFey8k9J6u
P0rodJ4GeOPSgQNVF3n3g9sblkCZU7lz1xqTjIYxw5oxnaFJC0SokKkdNZrqGMjP
NcHHS5J6UHt+J/EigTTwpIGvouL0m36MMLJeYqskF0ooy/skyMxqDy8SGDLl01Bd
h6wITluJOZwyBZGgN1VbzOBqaIlfSQGyDMIm+bs8YYVjJzRblAz/GbHVkRH2Z/YB
3MWkJ3wE1nwDuPMHHUM143WG6COrETBdaDDdoWgU8+gjZ+mWJvFzLBZhq5Qquva0
QOQhTay0cXQtApcRU+5DWvnhHFHu5kSazX+QxwqV1uTl+JO4b2S2zNNZShRImglv
sIZmq9BJbzlWW9v2Tb8iv3vWXoKll5YgQVKkGw4YYf/xMeucmCr62dZT8ThFeYky
8MrfwA4lwu+716fWC5S/ZuHW4s3pQSt0LbAp8o0Mk5RUUr00bBpmqnOUkC/A2kRq
Tc36CXRam1nENnDr8TSlP9N3WIficHsfj14LwrZc96UwdcxoxHpzW1Z6QJ6xjYpr
eV+If/Ermt6kDdJbASyxQTURhraU3r7OSiXKuMwxpG3UNDxF1djl4+jzFQywGscq
1ZrYQAM+JK9TW0L2wTn/Ok3tXQ+/+rX/Ixb/aQEHZio5aKmR/Izow/Mcz1gCWEPD
UzRewV9Dp3qNJ+jQXwBaDS7vvlpeDat7NWQ8ZceI/O8Ser3+pq4A4gjIPZTCTjtr
dkjtf+oFvUyewUo13LkwNtWM601nt1/f4H3CWGbIthYPPwrfgntsTmixBaTRCKHv
CUzbre74vJ0uu+hU14NPlLySrcMkPm4Aj0CEP6odWgZanA3DCcqeKYS/3tSLuWBL
At+d2+zElQ8NZ0VA0ZEeI/yax3Li31bU8ASQD3t+859EMUwKl3h9k28XC8kEqayK
n3yZEUnLq1XG3GPkmAPiRVy2bd1QhWB9d70Bn/vkpj2Mv6o5KzhApq2szLiLzuVJ
KIyTBoZEQFAVWgl30en55EWRqe7/8wXgl5KOpVan1U4qC73F4GdC3jCD5WqCMIG7
KXF7rxs+VfDusXM0NJ3EY6C0mZiF2+d39nWJ5CfcmiYId8F74k1bV5Ie+aD1HNxy
z9/fy8Xz1IHh5aLa/AyzXj+YMZdACGZZO9tMn2tHiHHiozWIrkceaytC9CLlvz15
txc+sVcx7vhKH2meUF4v1fl/TJwsWNHcvbKOD+gcNBnmJ3BwoRn9IV0TjUTFgSz6
YHe2tw+NZcwJvSbAwJRt53cq9K6biAD0grScfMISm9oSCbLnNPDcTJ6YeFwJx4qL
rub6waBaG6btQbbEXeIZmEqUNRkI7jznCkyRmDmHqBay0mpbPkWLKpj8MIT6wqzv
Ql3p+8Y1YaEBaHH+xPFdGhgxuZdyMzEoDdJlGw8ddAvg6tvKJvMNRY6qiCeaFhNf
nMNBRt5tF8jzzE+yFalWYRgJJbKPmvibYPM97faHah/kRUtHAvY08rmxv9jO1Aj7
qXwSaWfXsvKsoDekMgvk/XhVpMEJIUMxg4DPCLBg5G/7wiBOI03vu1KDTu7I1BTe
8u2TeiPWVZOdu3ALRJHTL3Vo8PL3G6MWQJOkKO4HxKR9XWvt/nBKj671KiNWz/17
eoiCAjH6yWNIQIU/jTQXhD7zGaINgcceWMvjUH6jsbMKK3NiQCl9zQ3tHpbqzign
Q2nS6UoFK22+tuvSoCitgKX0TQzrcTJb48CAkcAk2GkiEJ1D4Xk4zVAx38yxYwDY
eoZkk0gTG0Zh55NCGqo0iYF5qiy2lXw4BvIjpxNyYbunVYKDBbHpw4zI2I9T6Znf
vH4wAdgldW6yFljQX5lCBt8nYqk/HVWpZG1rd5Je9h6kbFAtdlEWhmPJ2WP7/3Dk
/4Sf56+1uGITqR8ij+GEom4/DdyVqT8ngTAwOwUQ0oug71nb99iVrUtY9Qkb90T4
ZTtgTKZrP+msMxjfT99MZ78Q3uq4uZGUmZjpvDsnUG3NFCjuNOltBMPPGC1J48UW
iP5bFahH5gzA9TUdXbOmzLMqBI1uQZU3HHiwPsCheC5AkgKt5gPPdbIaQdpzPLnL
T3TBdc3MnevRY43F3OnhLruIeacY14NFgA3m6rWo+pZ9mt943UH/IpH7l8k1gGvb
WYp4pyXrSmu8JRDYy7oor4huBd6ftnFMboKqbnfs397MBkVfVArZI0hVdlI/ZknA
ZnDSGd+Q3+Pw2NVpU3WHqmNrVhTMw800CrJmztDUOPyKYGYRyO9k+Q1OSJ8Wl+fq
nSTacUOsF9DVyhcLYK9DdonB7jmY2D1CuKZb0C6e7c7m6NL28HnPkfZe/Eb65mZq
2VizXf8bSjAh84K02chDVJC8ZzOL/hrjpu9tjZoBMRd5ZvVliCvxwiMRXPiJa68v
Ky5ORrd8oYM2ghEgwr5e7ql47JRsumkWOOgT809KAwryMuS8ohg4fTeUvKTEAe4W
uZTogC/RPE2FSPErILUg1k02gW/p0IMzNvNOgBWDrTbiPnf1Y02UIOl0JsHsA3FS
EuQgAxM1grcuhl1YlOIsSJuLGsF5XoJyVqMDsMlLU4pVNFtU3C3slDvPXuUin7KM
BgcNKHq3iOsTDSjnuWMg5zmbR8DzYVv6q7gBvgs5TGd4B/j5PoHKdm76eng0q2Bq
99KCtcL5WzYzDVUGGCr6q1dD5v7To5pLmK70lhMOR7vU8DWw/03wFTAKnksfzVm8
fHf0h18EDW3LqVBM709afHcUhmtdp8aMm4Omj5EhmPBsD19NyJ/3Itv/6xF5p+8h
S57LYjhMcE9YD0e86gTVw+AhVGLbQFMDZk2wgGoDJF6WvNkBX7MPoMbmBMOsWbKf
x+h/9ai5K5jS8yav+kyhjZdZGH9snLd7rKl7ocHuXyzt1OY8CjiVLBKTY4r1n72N
vJJFFL/uEWm3wknNYptSkeQVSr8SZIA1BqH5HCcVM6whcbwZvdKYuxlUxL4+jJrG
ZQp2zbacL2p3aeQh66kt2NuuxYFk1sqx31TsIf149cO2MK/LJdnDj85XFXbzohjf
6vY4oCW/zu9ve6//855AhEAtVv1xDkLUSj5MTHG5fiaxkJQp6om7oMzBOIdoczSq
+9kH5cKupGdETjXZWTqVQLxc3sieShnzkSZ/pmjaM1B8d6SyiTdztIAcJRDs2YmU
MXWkB5gFRY/fZF1b3QON1muuS8b9Rz5eEyVTd7jVcDjqgqXYMtnCZa/bLZPzkm0r
LsNvlVRCks7q0wYJgTuCld49c2xPM0odJWTW/Dcz4QxJJtj176tQvkevLsv8bfUV
xie3EBUwWQsxLbU9F7kdKRbwArZjQdopEO379vRH2czqLnrxPtDS1Vv1FP+cKyQz
WFREUBKwVoqmMG/LQJ30tFCsY0/6wg1r7l/Eyya7l/nN69fwttobvRCm2cYsNNAa
a6eHcKQCPF655d0ukTq+XX+7A+K6FbqXujCyHy6sCIT5ZnkJkRwys/AFMcTJfdaH
bri2m8tB+8RHI2KnUGKhNReeQ9fYyJtrmC+hoFufvkKHeo2Lf+dG2ISkMsuWD7IS
D4RSGTwgX3cNUBKoId6zxg7FlS3ZMahXvZnYHd7w1Ej6mZkO9T/mRO4agyXQAatx
y5qHhBiCtVcqBz98cy28OXzV7GxCL3QeiQtpoQHZ9kO+RLFjov+axuc+vAcH0H1L
aKQKlpU6OfMMkoXl55GMQHibpvUiblYJZYaGqEW8Eh+T4HgPgkaLkL1iGWbbZwce
l1BWhRacifqyTKUyT1hiWHBG3uKXW/T9ANEv/GJGZQqK30OWOnvSfXEqD4EdO1JS
8V0GkDXegCWoqPg3RjMyUtuLHd2Q4rZaKqUgt1tRppXraz1aWsr0ZEZud8ZkL/3n
8G1kd5+bJFekz+i1EbAS+u/anO9XKq5x3m6ESdYJZGgTOi69ldGhT2AcIzUJUsyr
Igp80jhegpcnzCU/Kh1XayafktvVnTYgev8Hr5TwsIhuIY1KLJboMdDn3hGx3A59
UUQ/5IP50ttbiwtYa1R4wUr7XQewKLUdirypZSBaD33h7fGUnLo+dQ67oD4suyvG
jIeygRixl2mg6KZa2zNkeJtOcMUfoMuUTRnjgiDEqWGLO6hFlcxNrA+XRXXCRAqx
jzlnK0a0uhv71lSpwH0uA5BRShp9woEbUkKLTqiWXgM5g/nOBbjBG1CqF/FJQvZB
9Bw29A5qoabPswgMgfxA++l8um3848vYHf3FDtKzjCSnwL80EJx29MbxyzmPvB88
ZUSx1ANc4D9+lZxcCThHOKajuc7s2LUzC15B5CbjCw877TVc42d02v7X/5eGmxyw
YkNqL2l7/QVuOFsUd2BlcHp5/VhMzjsCSCIT5Os8vkGGOju4GzHQnRLNvdBfFFNo
vW3W/dL2NrEOCKshGAgt0BdYelkIox7HHeBwRl15KzSdB9ObjF3rkzrKPbqArw/y
AFjb3EfMpukQSUS53sWjIvH3yeIS38ExK09rMn8xql4SvL69lj+SVTFwDxo2/m/F
kQ2G35U0CtqIlmTNDDUkxzRwip6tajeuMIxMaLqiCecNLwmF7Lp1ufiGXXmjo/Yj
em8kwiGGNURURqilfIhsEvDzGqUwVtpU/7Ge72pV0XOaCHNdSr0CkhzQ6aSc2l4s
Kt6trLe2ncVJLZuSq9dx8oMF2vnDtZOrj9+IfzVFqSg+2uCbLplyIf5+hhnv6LH5
EOytPeX9YVx+TOr7Ykb8QzOyOHg7dcJdObGM1Jo16Ub/3wtJ4yx1PgOUOWQJddW7
haMSy3VkKNA31w2g22flgpjo1vHq294ugKMhL00fxpKGaQP+6ND1ixPUOlpt3Tzs
c/u/ygPTE/hwpI8DVsWBacwjmTN8XrMgHK2fn9ku+S2MGluX0rDw24V5SQD1Z3fj
wIycPplhJTIRCeWRfxuMFjy2nTYMErVyL2qF19tgh5upfjx33+8vBZLgNsenfZg8
f9ZJ/a+TNBccu8016CTlRG9t5Qx4oA66+JcCC0juidC9zT1QdFKPJsBi42/KIfjG
GAaDTY+ALVxyA32QaeX5Dt3Vbn8Z1V25TYNWH6mGtIEfUkTlYNUyMDgw0ltLa8Cm
BRvf9aLTx9u3tAYb542aeegMkB9Q2D2Rc5Sz22bF5BJjv57JrZQqiAYNQkueSbi5
CyLzw4AqGrdBwgIWEILjXVk0wMAYVtDIpVyvLM9810rJUUN8ybwP2j9QAKmhshsg
OkYsR+uzDDXFKD4z2FiJMzrbiMbaSRbZ0XEEHD2A2NRmtdpZ1CTvdEsC0tQB/Ke4
xfV12IadkvujQ5divQjMEQ19Ki2hxSNyY2XwL1l9fZXTTX7CfSJxXeWJ8E3+q8qs
4dVv6Du8B0OVq2Oo3rZ7fXPGvgSrYA5jBbWuvbcljZfwvW01ZpxYTCFAR7u6hYcN
8nGyQszEJOa2XJF5OnX+C5BPM9OsswV5Lu/k5TIDpVHxsPEHOI/uAZfx3GAPxNdy
Hr20uPrMkMAfxRVik8j/f/uyzNUMPamo8b9ceOOJRIwyAhsxe7c87bSX85IUKn9m
Gu9PJfNdncR23TUMxzowKur6EA6Al9BPavsaUAzTJ1e9X5zCJYaTsrkzOMuJ+iQf
d7USMreMEC5UXR0vvfV7sa/BfRDJrmjjEX/EnoLPfcjHVxDP8qdsOnzQfN3+EABx
+yJvzADml3UjGR0y0fPgaZGAzwxUdUmJoL1cFKbZjh/gMeW7+cJSG2Td/MArknjZ
fDwXTCiG5DflVdQr4iHPbVBQnPy/pEsLwDq7SSTRg681I7Aj6Xuh2is8JaqQWU+H
6kOc3TNytZWYPs9d6fQSJW5Gq5qc6150buewnaouuPTgShH/v11or3ix1zu2D6Np
R0QXzcF7vH9PnWQVdVMUFGVQvvvXxhBwoIEddQX3mGlVoiuc/WP7yPNo6cW4ORlb
Q0kTvA/5unKp8H2EIEB346+Glkod6MTHEfkHj+hfk4XVypnbtDoENIxCq+3WNaG4
+gLGXnnCP7AeWAoGDyl2utXXXIIzDdgt6sbMdAN4/tztRxOSuYor3vlrB0vLtgBv
t+rV/GmyE//DApnPMbavu+C//02jMIXYnYTfXIUuvGSNYIZavEw3qI2nRsJnzNLt
GVVFmXcykd063NMl832lf04ijgMiaf6+2/LkJVGsMPjeFZKZbEfBsnIje9Wp2vYz
Ceg9OZyFvzZ03dcqp1+c/6rHCeolegBYwIFvOQcp70qhu/KHmbjN1QlQv6yMd8pn
6qnIgL9WyIS4gfQ67rZl4o8uC/52BoTSnAZ6pxCpJ/juyeimUEDECQsuF56VHjwG
6QOzmijfN3ll9L5zCrWAPiGtrxjuhorsiu2lsAiK8t0c3XxnG2Oe3Dirm8hI6q2Y
vUxfW+IoxAJ4eJLJBiotk7hgLbo5oNXdxoXofMV6M8x+lxOqiu2ohRCsDjBsYVRO
/sxywhPvc7ag3FNX2+PVlD+VZntnUxU2IrtKsY1Yn46qKMRLcFvUhQQb8wYnO1Zb
a4BSz87ELTT8+bgQd7VJLPagTslSF156XcaIO8hdWAnGVjmM4r+JDDp1OD9LuKOt
N/L4+Ie+sxTV/bHY0kpOfauSsSnKE4D4N/NiRZWzuuHPcCp8xTa4CgQzVo4LLxRr
3IIbBz0T+BqOhKsvC/tx18kPljnR+atIU9Y2cBENyRTa4yJg+zvvSUEE2j/rtAgD
ZUfCEXtLhwgEFN/OkGfOLe0lWWNQIUMFtBOPI365AApwHaMaRZ2c54gFrgRLDcCm
zH3uF+SG8GuAPEUNRwpj2hRNWS7LqNYsIWV7RHA7W6C2PeMsyCWYTVHiiCg7FVfc
dSkRNje5s0igdCb9tsn39y3DEdbnA+XDPsfL60dnn6jBu6+Hvu8P5b5a0wXLzcJb
H0zEr1kHPo2tU6jumXroor2bzwll/tauHXjn+kTho2a2bmIz/MRpgObCE2fCmG29
vs69d0Ey7iNRNPn/JBW7FE2lrZ2XkDBmdKaaGP4SptzqNuCIAw2Iq3Jty43HM+Zk
V+7kY13Hydt7fH29G9Lk0jeZfen3iIp+OnSQ4jEHdlxiDghYsCPRQWckhEncVJhX
ypV/btqsV7tgmSPPFnXyChfssCvdJt4+a9U4/pi2+rUi7BEuWmkYc0sdTdJoSjEQ
nanDsYlIpUczHNjfJtEd0uwUOPYESTBV1z9VH1shORyY8d592XpazSmeg2cX4XAK
203bwuaofSgFBCcWwsE63X24hSBCbSqj+M95OwjLGUXOsxBrdOlQY2LXfAKA0I0l
e5ir5MqnOxmG2voSkVDulj71DvTUr95F6qMgkWKzQdukSogGGsA88cwxhEpnEky4
/Jk/txKhdALzv1BE24HkyYrqQmOVHXJ1hxyAdq/bFLv/jlqtWpjDzIf1f1PNxQ3V
6UVPsQ+k19qvmj68VGiB7tTEp2O3jOjLjxuRFqLAFafNPe8hi3DRY6cZMrb7MNjH
UETX3KCrnYO1IAl/CjPib9o53fo2YYlr+2uc5ZQofTAwYRmB6ZvYLfd96W3DrgKX
MhsjGTSyNou9Qc6v8cXDWrMVK97HtiVkZuzTvP+w8T7dQmwFsrCyiP3XjB7pWCiR
HQkWGmH+jIE5dPsc8sTJCKzwZfdzaDdUjEY1D+RvqkcKkn6LbmHNtc4QXGT/81GT
dqC6bd0ovhlqesHfqlb+xc1orwTaeDVPBIO0yGiqdrJiX+GMYWCHN+RfL/1irV9q
7roxPTkP+4QP+UAi0rlVKo556+I2MsnxP+d+btb35/ox3Xq/wc1jiXMmmY8qRJMI
97+DIAaW1RuhGThfjIl6Cq7a6TvTfF67q5Ky+vBZl4DL+goW5Z8oI4oy0U5VZWgm
D1wYkpknQ+NflHedRH5ktbEO9pNRFEejIliA2vZv4x6Qf5itJTQAQ0itcerm3uXL
uAutc9+4yeOxSUa6VSQ8Z84kh/rZeDw/KMlhTg+yqJRtYndUFwnbh9pvNljI2a95
etDXN1OChof/9yCKTrHiapMyIgj8RUpzQLvpSujfKukxZGfXqhYv4VQgGLp305EU
zKZf/VXMiMx/+WPzm4b6GjBWIaMmuMVvFYf7vqZr3K3Irfu2MBD461bjP10937mL
4hPtDFNYQ0jZsh3gqY1DLO1QKsozKvuWa0LAuWeHtKzzHG8zaUxBjL7pj+TGN4aK
kGs4VBjDDqzTSD4mGXYSwPCoDLXiJHpvatEDpBj2FQX4Dt41iFOQTQwmCJmSY0H4
A5Vq96yB7qncdYPILc/1eG8bFdB+zdtnO6zI2123Z9gmJlwwSIpwa4PqdvkkIY9h
eOPhLfCpHkFxhhEzFu2lf273jm8gadjMgLxCSIKVa8200DroQ7oWCqFEPhxOKfBI
gczafe5Suv6DoHaHZJKAw9ZltG4t3TaoNm8DDpAuolFc4NGqkT2ygJ42Xe9f+J+W
c7krABaE1/oGo2BdVhHXptmEbRP5W5Ir9KoSjtVMKBXddzuenxYI0iIelS+2itUe
Phh3QYuMQQCQ/YXN6SOxvjsxpG9DZeM3BghUlpl1EmP/ZHiej4iE+sDZZVw1zsQh
fdaBsvRT7RI9pz6dVya1LF7pPPjwPHdDpKTe9vlG0SvJIWvldhg8qgHqrLiVLkSj
3Vn5Ik3stTRRGp3WC6YrzofGyFcW3uy2ozk2A/MVfPqTFanmagmP/DGe9+3fEwPN
dOdslNX4ZrC2Vpc84iBqOIh7Rymivsyhi1lfFhHgQPYzqepyDYL+JOqIIRj9fh++
RjDH2PGEja/WzTB5vWXBEYHbjom8eXrCg+HE16EBPlH9NTBRW/tmEq5CBa6YjGga
B0F572HG1ldafg9eKimZvgWf3nMLOyIunKE404uer94cMBYKjEpcbqaXDlWFMn0/
H9aU2CYa6/wQwHZNQOphLc4UCMbe8hZSGbWbLOpVtlxJ75moBAgVrbiBay/b5AwD
GECasPXjQ5QIDKoELy65YD5C0QB4gmR++whX2uEfYnFRQ+42Xsm+KsYuZEzD55ph
XHk6w8y/VzexmOdM3duDKqvkMSZlYz/eTXj0gtqAIvbi5wFLz586ntRzZH8eUBX6
3P2mYjKl2mfofrgXoeDmfDqqAjXausu0gy/WxkQOzVxCYT3YvMrUOakag4CsOot8
lvCXuyQP+rx2c9gs2QannPpSGrYYBQxkrg55O3a0xBBlFkR1KUKoAjyO7yfTbN1H
Vv6si1Vo11DR33WOXz8XqFXQFN+ebju/DezFKbbB4DfbEP+d0ENbAAaG6aX8pEon
LfH59FWJb3r/LDsDorejhUDc/c9aand2hcTuKsGJ/lZcY0gB+y9lEc3g8JQkBJ4o
kMxMcqaMNUXfKJPk6A70vC+5Aq5o2Dli13MHuwUF9ZmYOBprc0W/U6/xLNeMrqmL
IDiHx1ENMCZj/M0Z/YUaptcYzFdPny8y/Kc5D1Y1RVq2PSfYW7ajQisyyfXC1DrU
ycpq8WSWeSfTNOCWZSEjEdazmdVtPDyOvIFXkT+WMphPfnIXZE/ShjTqerw/aLKM
KbaUwAVy8lEA7C6Tnh41bvgGQJWspkymqYeRDrVfsfaLo1sCb7Kxzq3NRdJkq7H3
cFfWnbalWMbcDRIl5s62rf1oA91FCjGaGKgMgjbdp7kBGojp7KlJ5u3ls3MXOqvo
4SWcb3vAXiYurOw1ohhhiPndMqrF1OezXzX/hdxwbg2FTfNyf2Ogbwo8ttw3Yi9N
ycpoHpbq4d5Ynmi6baRFh4XuOZmM1+jKW3nTvZRY9ESYqVF1YctCi2cjqYyMoE6O
KXnwGlc3UcIYyUkClP/6kWUumzUwIFrqrOumjmhBcnI=
`protect END_PROTECTED
