`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6DLx6E8r3gE7KVUZ0Y5WXykAZR8QKCfRwVbWjQmSTpZ5Kz8DKQ5HHkCYGJwfX04
viXd/FDOe160vEWeBCE0ki1sbXl42lRTugH3GfCzTeUzCgNL5q/DmyEGqwVmx3s4
N/agNY7J+xCb54ze/HmDwJASlbJ00Vnstq8TwiN1s9z4Zh+uhZY2ox+niFDU0CPE
bzFnK1SQPdMI5NGpBuZVx6k5wxMJ1/wr+elykqVAVfOlKPR4YYmBWv7OQYUgc1pR
KHTh1X5khFD5qMGzb/KtFuv7VAeVtEogn+qs4KrQIOvgg81cgvfVcyRF+mtxRFVE
09WKhtJqw1n3o9X0fLLmJk3Ez2UDIFrst+jXKgVmZDzB0uWl0TDafdAGSARqn9/W
yQoe5kYG9/b7uv1oLxCqe6eNgayDp62++vnhJgztToAAzRWmB670um/kXBjnhhLh
Wb/wkOU4+lG9ZxUETyBLekG95uBWjXYclZuIO5ugUlh1quOuDW3vqiWrVSmv1yiW
MxxGtOsP/SHHXP25YSHCJjaJ+hRknqKBbWJU+3K+HbiB9KQ3fBHFJmaBkaqKs6K1
vk05rZCX7NqAmM0TGwOdzg4BHaWkf/GHlhFd6VqlSMCfn3vCXjr+062U8bVDgKCz
1e6cGJi8OqOtH8f8OewVDrYKM4fOeCsdQuL4KQahGleNzHUVJpNOx+wMqc9dOKar
uDbuSQOg+e3h8kh+OOrlutnhKj/nfHpVgG/fDElmqug=
`protect END_PROTECTED
