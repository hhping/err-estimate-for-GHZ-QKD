`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqltHcV1ZlnQzm+Eiw++ht6CgILjH38JAF+SUyCJfUWfXDauVbHJ9O4crf21WxKR
yKI4ie8n9p88BrQRYgTw+g6RoqAOSQrWoeXF5VzzIxnGO7LORDuCICOQJ2eHsJco
c94xzPCfP1O9y/y1SdYG6cAPhsrUE2mmvpSDA9zeUbWCT1PXKpSt/K9Nr+E64/F0
5rpCKd1lma67w7edBFKaGOfRY8Gj7uGtEzZ+LxILaIJwf/TGZ0US4nT9dv0nd/4w
TkexdFzizMjd19QQVIZv1J2HDdDFTRxLhyURGpalbpsybTp0BqnJbC8WilpSSW4F
qSEvohzEo+RRhbjo84WWMaLgdBY0M4TZwGYcH5hjkuJKuj0/CuP5TfWDYvUgm4jw
yRNQdr8S5C/bunzvtpZCZXPNrg1R9luLiFthQ1Cpl4clL2AcoGObo0CXpvFkcjz/
oPVwk0t6j81KXKXUKPgA//DRdvg647egQg3JZgggbiqNRKYDC59IJMV2exl92/at
75rE/UXMdR+ZCi5xL5R1WPmuqQZdBhkmVszp6QxwBBw1lF6h3ikbK8I9r4EFfi4/
Bp2G1JgPXGAoY6dUpvxvTSO0RKSn5f8Qr4ypLkiTiIjLBgitiLlkCEZdog/48gIq
BYRRV9oDZqR/a4d0qwgM3oN8GcMSVV+HU79n5QS/f1sOMn3pc7UXLzpIo7Z6zd/a
XvsULZYzJ/yEJDRK3sLk8XI29jrJhCX46NDsKYKG+QBakSdzlwBKhglIoXmtpRTG
uYLlTF9/ZSTi8RueLwN7Yjxuk/UJy9Xwy0XEsBdyG5M/GwsJ/MVcLxcdmXz3J8d5
nnpIsHmFN6+HBvNmZFIrrDIpOTktBJ2G2aEgxJc2RjkAioK4yO/v50JNMpjegidN
`protect END_PROTECTED
