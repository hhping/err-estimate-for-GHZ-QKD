`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfIbNkHnzof00h2ZekL73FrLxmBCOMMj0iVJiXfP6YXvc2QZLpX2Btp13o96BwnR
eDtS3vX1EjVzRHP2OmlxSFl0d1zSvSEaGNJXC1AOKqkrLoAY1TtJ9fVs/b6eM5gs
5ZJ7wBncU5HY6LE8+O21X1uHbDMJgP/qc4oEPz/dtvNe4/z9+260VhCYd88EqCrI
Ze81n26MqhhYn/hvYrFydNrvjhjBXzMGauGok0H3E5GBeIDe0MppVpRorN1EYOKN
tQ+iSs022miui2w6Brz5danrZ3vZ572yTeaIahheUpTbQ47T4XpF8cYQBSR4BFqU
Hr+/tmHJPazIMjt5s7KZ+vSGbLy9oPiTcNkNIhJf8rj19WW0Qohak4ceGIid/dO+
RF+6G6hKZadlUJTp3yGaqR/lmFCPFv1HkZ7xAns++/ofCfi6VJOJYm5vSIZIrvt+
+bqg2MxFBzbkq9pDKFOuN/s8p2YyVsE/RJzHWRA+ikWiJUQ3NGZFmGiXFBMoSIux
v6ixdKFaAbilxlEYglOEekWMh9dPbcBBhVxOYrUpfVjbq0THWOX9P4pVFRrThR+s
pTU+73yyLj9sT+Polo0W5ZVoo4CHaR2PZqJL0QQExIwYL1ZOB1SpHZVl13L11Q5V
jHpi0osz6EyhK3ajB7/VCeLIe+6ThWp/lsrCzFhdi2XJYn8HamCa/YM2VFXufRfg
QsDrfBVIUYScHp7/nDvpC4uQqtDVhgI8IdARfg7nmVLf4Mi/zHmu0LFOtkcHyoiC
0BtZClV3cMz8Y4D2altOGaOlEOcLH51xopY2U8ITIDe7IpKg74kx4V3aGtDB5LVE
RjNMDrPgWYdLCYXXvw4WoTq+pVlnw2Y52Mk9axFu5ckbGjYZ2g1PGKazQlOWQ34y
to1+G47MIHy2ZF6bCAdKmtOXUwSnILKxNLpj/X0wxubXNJWQ4qzfrwXeULPIB9ef
apwHhnOVgYAKr96rn8PY02fiajSP7BDvyxoBSWGCmgE0VqHKKKXwzlWPVoHG8rtH
`protect END_PROTECTED
