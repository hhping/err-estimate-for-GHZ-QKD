`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4NNNLvqMuo0S7ZIQkRiCx/C2v78eNVP52+zhUByXSdR6koQzhHys1qoKDqgW8rZ
aPz9kpDpztmQavnR/Jm41YNY5xyMg39bHZIqclr+L2UNbqnMEUkQTWPhoitVTdBf
v2Er6ZGlU8yK2H/MBdCczPxEYo8cBQT+LybOOu8CqZpSqKHjF9DYfB7stYgzqcHz
77iR2V6CcohWj/6Xvj6tppihnPN8qlmhh6/UUi7CccpWxbA2Ll4+rDX27EUoJcMj
ok3QGkgGXf3WJLGReCvazBFAKGq46iFs+b7Xe28KcDNAD/hvzNWdNEfhHlMuf3hz
N0pFfmcWavLSv7Rsy914PPSa7YRmMAhFjCHJw/eNz1K5kjfUxHxiIFcZpbbCE5At
pzFpXsewhRwWeEvfMdmC9w/mLGFuPQ/0d/R7lofWUNHAiOxzrWrTMVVsOKBxmf+2
GVpdXQrtBz7AgUeC3gD2P0BLGIelegEtYVQZzktIfWujEXSL5kZKzRZZH4+MyxsC
nfqEMWhE/97UfB55NGOqVrIlUMd7g/nNLYwIrgPsXIOm/KPS83Du83QhowoorUJP
fLJ4jIZtRj+yMurdiLLf+ICQ3Qbs6a0byTO8/+Zu0OtGj8P6dlZcCvK4uCmvmw1s
h5F0lFQVFJfXg0z8KMKD8Quea37bKAvncxo/d12jM9PD5BTqGHbXPpTKNZ66HEzS
M2Xhqrswa0HQhYXq86P/UGaDrv/tw5Tt7tVgNpZi7sxNZPhlUtGJf41W4ciqTBdr
WXkQMJj2QlTOHP/d+hv34aW1/81WdLnKcIKUyS0+gti7kZkGzjLhOA+ktTDenaTv
OWhWZkHigAQQ1szWnTfP7rU+PGt982PBqzQLOcqTAngS7spDDkl6r2uEZvoQ1GS1
qFy8akk8Cxd8SHLKQAXNMbnWXsZMxvgt2Wfh1Ty7cEEi+LYZ1M5S638ICecDLWF8
q+uXnCDpPtH29dnthd69zConmwMXTDHW0qJ/rkp8mpd7yd1cWji75Tj6umzE04Q8
YITFxbVhAUD9+yNIoQ3T9eQbjTaJG9LANv9YPss/3IibrpomkPh/9wg1nU3LAZL0
7ljMDA/uwaeemShuo25PPM/WC8njA9hDzp/cTO4ynRWOJuRfWMpzNtIi5bgTAvqh
2kRE1A+g87/qnYHnuR2wWbBol3T+lYI7xaOdO+m00EQXmbNuWa3eg+N5JtrXlRRz
n4oSG8GATpTAnrIrH2sjVi7QtUlqsT+nAJJ0VbCtvMzgmz1q9+QJSjTF68qtmKn+
Et9b/4oJq3SM5Hxytac9gnMujLCLG0UYG08uy8Yh64y+S8HCmBUXFRt+JfBU2eh9
wrUBoW5edGdEp5rOqrYQVTC9yEOGlZCxCE1/ue0aBTKcHJoQNMWln8Yz1h5DUgoF
qPg+viJlhgpMvnqceWFZ/184/81C1Zg9Ob1I0lKTC6ms0Uhl+ceC88SAJfag4RDp
Y5nCzv0cDxdCKlgiEDam4Wc4/agOCKDPLKQ40CMRLoRfc9Wa/xZWkjkrpvFCVfVP
AqNMeKG2jYPeXy8vcLPSgLhhhS8wjEsIjwHwsBZF2PAbmQQRUfir5Jdid0me0VyS
sUCPopRL6v9TNaUi7A5JjPLORZjgTCpoPnikYSUK5Mt6TO+H/UuUvfkWsYQYBOvj
kagNyPLm0wMO68kZtZDepfXVlSsrvvuWGc/qfQB8P9H5Jd91RNaosSxwjWLSeB1q
NnKBnMS37yphS3SomHxtyw==
`protect END_PROTECTED
