`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gLXs/tHTWMifz3ehJ4v5iVB+BPQdT3JLe/WlYNnsl9hRNS14avaOxn3mdEZeLUZ
ovKk2+Ca3LoLSMGgQVVjYPVK2ZKEoJ/FcgYTFJJpPoB66qiBL2stU6wQSDnSqcgL
aRPUsaQtptzPJ5ZVE/PMSimtu5Nh2RVYwMaYtodAvLBm69KCmoQvNWmTEJQD7wQm
P+zYsIGeSz7W3u9w0RgbwmFBJDZVm6S9vBfaWWjdfSYgqmYRQovKBp0AByDuLrRS
oCFptME3pTiw9mwzCiytQ7RtJ3eTbzvhmwpK7sKW54kcAPdj+AEvjiL3QBhGcw8w
FNsJhnpk444mOVyvXiSXOxRsAkGE01s/ICvJlpjVcopXc5BZ4EcMB0denEMBCGY7
xGyacqwTM5/kp962Ynbyw01/AHC04dPn1k+1wKOD1lHX1jRv8cNIfaRRxCiWdWyR
7zoJOVUmdKqnrS8ZY/nrnqlRCJdCbhgIYDxvvxOEAmuukd7+L4uZc5DVjVIduw/5
RysY7/pf+7mK/2pYA+l7NrsyGrHi3JxeY/U5zdtdT18gku65UxQqtmzg/jQ7GNxu
tQHGRNe25iYZNfpQdszlcw==
`protect END_PROTECTED
