`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VgOV9bePELr53nvtMXEE0e6gkvUcSJEqkkh71i2NWtbVLo+TdWRfH5GDNhMGnwie
hPmeqYDkRth0enx9iA5aOlk1VQta4yvYQbvd9GmWS7V0+8d9SN0Z8/wEmkJVD6Yd
ENVQB2tLCyVGoDGeL66ZEd8TmiicgI6NQ/uVm+W/RocPcYAYvkIJN1jm0fUCSPtH
2pyi1IZh10z/WO9EZSK2jxP6ItCHe6ACccWWkd4W3OvgFWHcl95ywUwt6FBzzSLL
dnV4QHi9VWRAjr3CbJyl2Nh/nn9TPRRpaYTsbzXUyuTO1VWINJJSHF3LfEh6QMfO
WeaKbUqy3cPDm8hsJiOdQTUzbdmQP+nGi8ejdZtK8gJPZxf4CRK2sKg6nOsol60Q
vAiUldkc+o9AnLMzs9QmhnPvdVGJA1dCIeheFpkK1Rq5kC0GdqdmZ92bmVGUCW0J
WXkVCiYShn9EdC3G76tEuV81AMhKF5w34puAYxmwNXvlnnag8gxVcVN6me+TrgKz
`protect END_PROTECTED
