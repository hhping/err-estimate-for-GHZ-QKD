`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5f6dMnxL4rE/4boR+aLNs8jo8EeUklF2NRsk4txs8U81yEO+u50BaGH/lBnfejMV
YzN8qsnSTMH/Fi6ef9aXpUrXtxTbMjZ35L1Nj4kwuFf3V9bgTvm0mUqN3HFYpe9f
nQfrpSxX5hxZvsShcenkbwwb8ipQxGVW16eV2djtiWAst56vhrb0MYkwAB4Dqoa0
PbAj6o7SEnwPUzMHb8emaI5lUfYTYvhieS/0+BMZEC1wa2hsc7wmhElyUMV4jfyn
TwA68O7dLQD7laIUMnBExMSf9Hss6tqz8aLPO7DMwhT3jcF6ET+lrrOuQLzOPPmH
ycSppbycpa2w9IqhNOFoWiDqA5zDKRDYu4dPnc/HwvIH73+CFfSgHybg1OF5EqQ1
MF54GdoEe8Q4SzVxINyGxJ0AiHnDCJG5JFDxM0PFqrNFt9Hjty3TE4hA8Ecax0W9
C11Q5kX8/510umXd2UtXnjaBd/IKwTXDXwYdJKJRNOvAXEwnW/XGsiRh8tnBgH3S
`protect END_PROTECTED
