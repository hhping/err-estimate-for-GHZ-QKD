`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dj6y5lKBgGS1uPmqQAGKePiFDD+9wwwsW1Yah1BH8JQhVCfHdHy8eyt8XV9B3dg/
7BJ8hehMK91B3F95NdeUyMW4VmewJq2+wcKYnBkdTQbBmuLnlXBT4uYSRYpfhx2F
nZQI66MpqCPTVS8iEoSSFmk3BE4RsObw2r07LuerVpWA72ut8EQLxtQlFuDUwC04
LXVz4h1iEinde2miBK6+n+lhw9KWYeeV3UdTC2jNfigMCuQcNG4Ocj6Cuchv0lfP
5kvQmdp1iXzYAKmvBwBcvzKX9Fn+tjvNpHKXQULsoT+Xzb+noYOBSAki1IR4Hfe7
DDZfnKPNV/mPTOgfQ9w7NIpwcQDH73JHtvojJRV1WXZbMfvnvXr1RADl7JX8Bqrr
zePrhxQsYlYoxxRFJMJFMgiHkS8Hb9I4fS+NqWxIf8Kxn8kjQU0XTd67P4OqBku7
i8zSMWD4Dzk9CBsEagyKQkRn9gKS8j4Pm04APSPcmmsBgEDD7X2uizCcLjOoqJIC
mkHRCyrSsvY13cwUrbFvv1gzluGwi93wNsu+4nRO+BAo4vrM8UMhfYizktVdjIwd
dkCtJn7u0BXMX4EFb34ACQPMMiJFeM8ieTeMJGWeoZA=
`protect END_PROTECTED
