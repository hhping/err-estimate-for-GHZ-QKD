`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6J5k8VRziK+fF0rgU/0cEZyQ2C1W+zFJBAHVLxbGSz96Pell2mhp0lCVnWqMHTg
hXLRENDu4XyDeBbqzlpCxl7Ds8UKVp7HkiqQJ3H4Ct9FfU/XvvQ4sU3kqiBQY3d3
0AvY6qKLmmh02ZdQajhbemL+2xQcs8gcxOuAnBuPpogcLXEm3VNXG0vNfubBnn+W
B5MZHntJk/w9vtz6lufTVV4WU24EIcbM4vkl+UxQaOoad6YUds5unbAkDoSPHztW
/1yrNdsDKg6ntXHNL/PptuKJVzVJiHg8DamuiM+8Z5Np8cUV7NkQooTcMlrsL1wB
toRJJB6yD2n6CswqrOGXKmlHSutkrvp6KqW1duwc2Whhelw4iAaSH5KBqdxr9uXN
UaksWyLdrH6/k/EWNKnTZTpeMtB8MGL6h45GILAu5d2ORQ1yu1r07q3POkc40DwZ
rZuK+uApMnR2VG4vjyK17PMgFP6GGBhxeNhGP3uGQJ3GW5/oRVHSlimh8Epmqa4f
RnFAwGmntkYsxkJrEewbMOENF0GcD2yTaL/AQ09cLt7LnLZyUprJyK6xlFxZ1jLM
kojINVh3orn3waztcM1g9c4muuTBp7T6BAmCbzR6C8RKf9VxuHRvvgVxVskDib2U
VXAP0fMs2zPihcbbponr0WN+5HkfzPa1caoxNtD6++WE7wcYHHywCI0k+fNUFxos
BnprnlnTNY2Fpkw6twaWNDq1UIvt43LY/RB1Xa5Qpk0cXY64HCL44msTRYIVDe3k
1acVT/0+/uF9tY8IN1U/g7iko+/3N3ykfa2kmIgOrjvWLEE23RED34jPakTkc41s
3ZZIAC8ZB2hy1TB8MNPhd3bVnZ27FV1F+OsdS6zp63zRIpGC5KYh4XvQ4mhwvPUO
kOPQtksRSJWLz1OJiyW8XzD38WiCnJDeXT+KjWzSo3rDxpuMFUGiYzRnBDRfMfmk
X0TTDgTi058dl9pE92C7I9rLyGaKtLmdFyifBBQa1Ix7FhBAXOvEaMfX7Sa4OKv8
WrD0TkUHtMDyLINoBsuD6RVAiQVBnGznAIeNF64gZceBzHt/f5kWko6qeLdgR8Fu
qG+iFpQzZ0UIOJGWzVw66l/4aR+SBts0Sj0XZaXlVy1/Hn+JeGL3omYX0CYPxoJh
`protect END_PROTECTED
