`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjVLdCI5U3I2oB6aEZ5MXicmGQxNtdSdB9ZckFeFCvsvGwLnkgdYZVBDD4sypmVS
jEC78sWlionl3y8hsnBYnv/PMKgpe07kWYNrrqKy7zK8OxVCSWL/kHfib00odMwP
Z4Ut5+XR475pcbq2dz/5BE6rYEyZvGmNY+/6hWwKnwbifaHWRzhhtEDOK238AqOF
L7K1Cl9atSIRMIFZkkiLTi9JSnh3SYjI2OSyx3uBram4vhU1urSD3ByUh02M1Oc0
`protect END_PROTECTED
