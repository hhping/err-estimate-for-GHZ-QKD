`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMTfec17fptlSbTmjxT1vk06DKDzAuObTx4+DiGkTEuZHguGABpfX4KQGXZ0r1FX
GjEaN1u7dVZQy25tFxZ2DuT5n+mFbA2XACLC/ok3Dy0PLPoFW3iUNpsnacNXPClU
VuRUpb/otleZ9nEMoYbjdBwPI/JQAYTmB19jZFEIBbdpkJ9YtpdRfoAztmSeI/6h
kP/Gw7YXYwVxI8meujr+bersA1rZ+l6JmRssyWuTP1E0tvSG1It3vJjSlNWUal98
Wvimuxz7loWoQ0e2JfaFNUI+bOjUQVACs5hIERj6QtjlqmQWyM67rhTErC0oPQap
kpqpWE/Gii2B7DGk/26cK6rAgxAuhfD0ck6JUX7vuqK9oz3uTbI7ZY9Z5fySF+g5
+iqVPUHbhNUr4o2MPxA+BBCU230XQUU0NMLGKZ12bhFgYd5icbzcReaYQc60cbXf
cO5vIqZxaWVopzBp6X8ApmSZdLBtDxaWVfGLxjgGnZdwysuH103E8rBv/aLtb9zG
V4zxJ2KMBY4rgi0Rwr3KR+UEUFQmuYxgep6ap3ktY27Vrm7hRlgIT7m6mnYIaUmF
foDSJAfCMCHTr8ZL3otEEdco/OcLJsTG4Rr2tI8K5My4788yKk0nFXhvbYJw1Em/
jajPJw2ZDRxljf0YmdB2AQm2A7OAGDgdj7+plMFFjzUzOvq+DUpxrF/p8J4ttTqz
L7GQPB3QPkrqZ5giWbsfBQHRdc+90yeQ923kFsjfvYX7mfGNNysVs4ss19KCRfqh
QdSPXkzQ692uKHVOf+4VKzUn7hLwCip+qnVzxT/uj4ER1wcJf6gYUHw78kVdyzTB
MNhGLMD18vhVbG2wOUnUoWmheE7moczgdURAZZ5fCi7o7OKxyzFuysuirg/AaJZT
mfwofGUSrgu9F5ldLhUMp87Q/oT6YOzjEEPtQUamuRfCVNbOJBvZOJKWRTHoOtya
KtGZ5MaJ/7R0O5T3ZlHTwFBwCkbgcV03YVVOiOAJz0Tl+tkB39NXzZSY16diidXD
CO79k2SMiQWEDZBthxC7d7zmLkgCh4JFhrkBVu69T1KGr9W0HGCFJp5FLMitGUjw
xdbIkqDgaDYF8tBttLtgyvekuEODDC64dMpUmTQ4yXyr3y1asTfth35puGj44dRk
XXEnsQ6AzJEDgfihap95gHEFlmd3P7xke7Al5EzLVh3tZ5ngkUyZQvuHtPZi9FF9
5cqRpdfgHTYwdZW78FKcMgcCNYGXRIJO9dlVxRmpgQ3HsxOVu2foFFVYXc/cpUgz
OstH3MBn2C0PLeLR/bMPo204znorYc+k4NM3WyELtSaNGb4AhvKNYAntpJFwUwnL
TrgD24Gm3WWrQYSotyOKACfu4SBjIeI6zA5K9I0ayTD4nfl2x/U4/Df6v3Hmhk+i
HtYXZtNKOfN/PmcP4ILbikI4PkzC3SEYeWWb+XQTskPVMK3aawME3f3420+1ElQT
0+Gki7AtMaNOkVx3MaserSftsn4J+q+6sjgDwx7f0N0GSjFfv7J6L5FfzZNbv7DJ
dLZuWsKU+Ua8q3KiQnOiuKVB5cbPKpEamUqee0mM2GC1HiGQ4RimA+B8Rt2Y55uD
RR4Ng195Qu4LfSf6l3Igawe9wMLEzXg6z0TQrAkHWrVIkbf4Lfbaa/Mh4Z8MoHTv
bN4k4r9YhcgwBkv7qugvWS93DhDVWv3GiceuE1mtpL06hqsZ8PN3VR4Q9+A3Lbky
NLyAUBGCXO6Wb1tJFm4TAlVGO/nwIojM4j804eQU3n5hsdBngwlnEgndhvaQV/GO
rQGUQBiY+lWqo3Us5BDfy0b2LVCqiGH6+RT37kEhvPlKpJsUS6SqMVm7Uf1puMZd
GC0aK4ZAOjmhR5IOj7UDOaJGmDy4ZBGyXF2TmMJm1/kTszPq58grVicqpHB4HtYq
WG628mYBeXhe12+2DXP65zsKRVDO/dD2qD4VdzaNiXVCDnags3y0VSn7fd4SvnlS
bc2LgP5lf8hxx9H4jAY2ozMX5XS83tjB7MohERCbyitY6PMFZ3Q0Tl9sz7dRDj83
0TpCuZjwOcDJNU9mpeXpstjLL8hA9+A+6qc7NvQfeNiB7C+B1t4+Om2DjQ0U/c3z
UZxWtiAm1sekJ2uqF/n/ZdKIN1D7AApy2nnxJsSLCj3p8y1tE9WKPTYVlmun0lnW
WuEjtbqmbdtykzIWlHFxDg9Dd5p66JAKuy1nn7NcrJbWVOomvOEqOzaGDNYYezqd
njsyOrjUtXlQBtWVb0Prnh4bHrgUxDsn899fxzOyW3bb5++WHDqXjr8tJ9dTOp7x
YNgcWkex/ULfYKVhR5sNeolizEjAmwWYod6dwzAQifk1YA/QmUZ0P9SIgMIzCkXY
EcJ0dz3Rdsd4LcmtBFJyBF0Goacl3cmmzj42VfVbe5hmPZYk1cR8bt5QjJkgZAXl
3pw050y+60DlhdLuVRVoEuIWc8Lw7IV/u1z+QknLbGW+L5TGIFrYvzhzXSRTwXcT
6aVeWvsJ98OKh+QihUW/PYm8n5cAnS4c3KvS2RucGS5iucJIv8cFo0WBGlE/Ko9t
fTdMMHD24oAwHObNrRWg6MOZuy8SCZM7L4My9tGwafz+7XgfNtp7igtacHXEASRY
7vSVovdkHn36fnda75qJgR03ayA+9DPToPSoPPu/+1M7fiilf3lnuNjwNnYkrJ9h
MeHxZNWslQzsU1UXBHesEKNZfSOEq2pQto+lUFHF4/aq6TS7ZgV30OSOfiCZhf74
L4OQ8vSai6sfTyayGCpXhHLsp92BzTuopE3nUcDs4gySJbCQhBc9/QMGcWVL0soN
lfdOjXpAUkvqeLViBEvCctH4U/RPyj082dAAUOuUYnW8WrNONXxBHcXTthiqmErw
LNoDJlIorVxgcDUgz6xSp5xWoJOTvUQGVfHxc+zqizHLLz8swCP5PZbwxYgTm7+f
EycmYaZOWXU96r3Boj8WZBUEupwFl5eIlkJBPh+BxPHCV6ts/TEsqfnh67zTgYpb
W4pPxGFQ2CUl1whxWYaEU3Gbu7dYAtovCmXESJqHm9Eqr8pmsg7UuHfEJkU3CKOO
MEgLQ5zpO4kHYwRR3OreUYeG5NNEk89+noy2tt8RVROSc7c8SjBZ52X2VODM88QT
rkCjz0VimG57cgLmZhS3BIx/g83ersjxhPfV1zfb0dv3FL1ijuuKFYroLRHKfi1N
6DyhYsDIQx4C2rhXLAfOKUQVbzcID8TYNQ0KdNLTwPhjZF3sWf+leS/7VgCQ3k/9
CjvxT5No/T3unkabVGuSdRM9RMmDvwdG1Ys5+Fcp7hWuEm8owAAjile3fv5TIBei
TRzzVbdr/akgOFZ3VnISubNthDPxXieRjW6HfnDuuHgGub6GcO6naK0zAsi4ZrdF
qBzjeScS23KP5WqEg1UK0upIQbYdVWUkEzOq8dT+mloj5CdJZac2Xyj4SurgSheD
BohZEjqQm/mFCrLrVw4dO9RUn91eyRCULQ9XCvBqGHRFTeCFr1J3pPSydCV7Wu5w
rO8G5ZNoO/XHt3Yt8Spw82YBpVDzamT6l+T8x5iEb8fJoVAGbNHByUmLkagZ3x1b
czEyq7xdM3IVWKNYi13AYhzIPPbl9x/n2s1Ut/J7ECzn5Bsnya2prRtSEehWW1aP
dV/zYMleRdwT7gF0Ko9+9lPKSE0p4WEIzw1X6DNCSOkPP5XEK5F+Iyyen6usRIDZ
gJv1qim64mGF5wyUAHN8IC/T9rdNfT0qhK+10O0tGie17oX2zKebO2H5WliId3rB
23hPWjj2KPmjfSxfA4dY+wwZClS4CizSnywaPqSEQDSdXEywdAbLbfjBnv/sOIJi
NSw0/O+gLm3adsZLrAlHZrM9aNj3dMTjq0kZ8aaxgBxT6ny7AoPC43QgkZbYtrA1
DB0X3jxDJs+NXAsWW2zANQXQfb3602/XegyZxr3nl53Id2rNNUO2gYZhdgKHyaC5
jk8lEeb9nvs3ZFP1FGqG3tnuNJz+gWr7400TKIk0MsRM3AlTKlIgcWo4Hr1uOnIn
BX/IxzMslT4zV7RAOEJYxQKPgYcyAFpnEsuQHegb7sqL2VLUZMI57zdNSrGd6KId
1EaCp3Bhx+QvW0/DPVALgGgURxR/ioSC180MX/juhckFKczokI2CFpKndkwyoxt4
KjiVeMfT5iOasCKTfn5/AiyQS5Cy1ed2xGg0hB8UuPfdd0U/yQ87lUnl4RBmylHA
soHMMY/2vdubC9wA8HR1qY7wm+zjPquT0YD3cdfyp1Vob9ValBTBDMh60/uzIUxE
LERip/IyFz9UXwu8Shbg/3/ULTUvnYxXWVVLDAzZRmh0wmORxE+Iu7ZBgS+LcFYv
HsaHidAttBDQWNtp+jRBlomSzAkJCWOwaQayZ9or/YFDIVFciajDwIR1717hv0hF
hTJLpd041F0As+pqWFPabz5ttaRdGHhuCCoKcaszLp+Q8nr2IKRnwoyZPWqtJwOC
b6RLgV5AtzKrxX2wHFHyEmEh+EsECm8aV2QAZE+Kf+fH7nLbTfvpX7ChisEB02JC
W2iLeFgW44P1JXNYO/og6cFtv29iCGa55WAVG1cnvgXbwFV5aivRbyCl6oAJp4yU
ECDJmXzeeNoYZymkS7L8GE3q1vmzdLgivMRCkrJdAG7aEmtbWqpPLCdpLhoqioUT
RwtPk/WNDUMOKT6IpW4udPmu420K7KXc3XDQZejH2V7b5rByCEEK1G4aX2SKi1hB
amEa5doPZnDWmIchqgvT4pN7b96J+GZneVSqh7Ml/dri6mw9e9WpvkakAehkHwe9
3oc2MAsetzi5gy/mZJu9mrASA/TzC3/efkQVetRLjqfbNaSM5tClHRkTj7gpcYu7
quU3zDojAKspSy30PsvdUPwrQplzAtPHD33pF0iiubX7OKVblYR67EKObTlmPHQt
GGCEIfj0yw2XZtuVTNxvnye3wXLST8NbCQHhSInxJrzZa2eXrZIQ188curw80RuY
ZXsc6/xTIMC9RVCJzu5UIX0fKG+TcP6noArBp8PGTU/j+al3d85Xw/swRw6xgVC7
CMzQ/2uYXsMXUEmFxlFy7GuGKv92OGjLY1qC15draAIBsnQDXA+yy1nAFc7IPC1d
4/QkwWctiGE1iftlXWIOBH32ZFXbwqs44OH3oersQRdoivE5VrFHqikrJzaRabzc
aFfa7EwVCJqEHib4qIk1WO+aJ8ysq8s9N0sy+GJb+cUooW4TvIi2M1wun4fqU6TU
Lrpxo3VvHdmtKrHGA/1ypnPAW8UxOyal80lZanFd03cYqmRkA+uMxFb0V2xjua3N
/v+ISe+e0mvlXg4Sk1VT/c+AZeM+A9Zkegl7eYaoX6Ly1DfKlmDACxdsywog3aSk
jxtJCCXeATL+lqr1OI90ZV1eGvS3icnU2cg7zfDx3NhBbKIqNa9jxPLdKptjgGfu
f9lz8/tTfsPad+AWTk4uSwSKOw/XcQ6YQcef+VKnjIHii6rH3Mxv+fkQnnzQVJIe
lUgQ7RyM/eEHCetHVg6Gr8G9n2WNirXh43iGYZ5aQ6dIuhdcf5P1Isr3T828XpIO
QznHfwi8r6qZmlQz1Xfq7x5HTLW1p1dT5MaTJRMofhyqMcGhUNy7DHvqlIzUGBw/
xf+M4MwGFF1k4DKEEABld2TPkvA6iYyGSqvvAOJquTlpQMMHkCM3d9vRu8Mk/Q25
YuN13jCwwSH5LzW547h26aEje5biOzx3FkkHNbPOBdyXqI8HUz0CptuXCBTK5w6h
X1qRZWGUwcuD9SSoFUuRdcIWq7sKHGpU4Vx1IFoxBlBGp2R1tVV4uDQ3X/CNejW2
fJtkON1JEIXn90PpMQCzZPXl54w4WMnZyEnwEScaZR/ki26/gWOqB3PYQn62IC1V
wjz5pU16vlAxrx8LG/WH1ggCFv+6ROj0A2WosPMTGFJ6nH4Zzwb0E4K2J7KZuL2X
hBOCS2SRYBg+QSKp45d/GpLbAyK6bY17oInllglcVB6Zee6xpu0BPtTgC+cIShvv
VzHJ3wCg0kSTx/xgGGUV9oXk4kyJJbdv9HiUctCAAfeAd8grk2BBhoEFKngJcwrt
BpSQOlbmFil1DpTVUg9j/hedV/BANXwy8B6+j0Nw+YC5NqyzgDwXBZTJ1X5W1o1s
LgNxVoqKqcpQMPmhBvDtfrdycu+rjeHbuGD/zVKzKhm/D77BRUGEbuLFkfjSaqmp
SNrzLNkiHYhUyEfl6G8SIXw4QNudXeF3hpUd4WXfSHusd0qGZnSkZG9xs37ZnGnw
hR9sHw/993RiGOCdfPykYD3x3AcI/jR8YTJOTWBSedoLkNxIB2VhuOU3G9/p/+HW
2xiP+RnAzeIOmAYrfK5p+XFGfkQc3vW3g8DebtC5YjgptH4wUX1ph8+D9Xqapm31
cHsNhyVAObyvMEpiBcHn51XxyBpyVnt4n9auHo200QMUTizxLnOHf8Zdh50Q8h/Q
SVXRJczMxr4JnENgAW6NuzqUKwO784Y1EE5hWBx/dfnLuTXzyAl5O1Xzi0Acegxq
odvZ1KuUOUVqchZjBv/2O1tZ9ej18eSl9anOiey8jmFeOyZ9J5/2x58H1sV0mLMS
ykKXaR5SvmPaJ0EEE9atD6K8ADjyrfQz04wWGj3A7jZVQmpSCrgSFOMHsBDbcBSQ
G6BwO/nKnAPvVaPgJsOemfBMUkbbrx81ghPC7yl7t0s3+kwLtBBiRK4rAjpFn9rn
z+7pfRtTJcCeP2HZR2Ue0jdUtopBO1iHZnVL8J3UnSyY6rm/wQUD1+6LrfU9QHf5
BZPFKbddh3KBoHGTHmCKWkHMYHxASxYn0gsSGCoGqwUXkbqyYRuGEjloRKl9C+Sx
I1HUqI9Rt09WrXmkeSlyfmhPHmNOFVutfKjEg+EE9nOiJAhw9TpRC/hkgcldHaWP
T7TgkICvAX2MmEncbJLSxkL9lZP78wcdZJC1UpOeKRLvZeLpKbyfH47gUYTr8WZE
Wt+Z0/rYsAEw8EB0PwDAN3telFgjWL5RBhgJGlS6qCyyfbndWnh40rn91KM65U3C
H5aswIEp8aGicIH9OtwEstUpttK/FPAve//oYZlOrbJErBHioQ10ttcYvmVjl3Zt
8kaaxGCT3s/0yB1/JO3KU8hYWeA21kk35Z/ASbsRiqn1FHxoqOegxZKliuug6q0s
NJ65asCFXVjc8R0sf3rxP8+ZNQSLSa641sJuChjYlULBXFVJykhfWS/r4B8L/++m
W8rE7JL70JW9xBK7wuyvjp8LEp9wuMs/FIoCDlj3BKfl8NGiAnce/45SlSIi9yD7
NhoektOWm64o9biFNPFBD3R+8BbU+mF9KYImxiQW3Y/14oElSXNgmmil8vFYHgXJ
QMRDPdrfv7NLLNIAwTTX3ZNqJAg0PJTknIJydIvGd9SsCqCBTLNye70+VGzWituP
hJw7/qg0i0hb4yAcWLBqz3C9T5oqlFR31eC1169mLa5YTg2nivjeSSoqZYJZeCeY
vqLPh6nHY8dW8nte7RHU+OgdXGIb9J7p9SIkSukPR8ScRknhJbhW92QYYDkQE9KY
/YfwUQXcFUQEBrrU5psDtJDtToFDqujmXD32UIYGBsXJpW4w9MphGVewknTetYYM
uD3UudsZ/2596WBrANMJk1lJYFeDoJPfFRCEGb/m2z+9nIE1KdBrwynO94AVo8XL
doGPxnuvqqF4j7XaWkcQ+3zJwj0YPvMGyRi+zEjeiwwMWXyu2cAp3OTIeA4SVK3p
Tev/nfkRU9gB46mfoH9W5P5rLs1YpR795nKKis3QZGq+Z3DE9aAmfgneg+il2za0
ptxG6+HOvAcQQpx/tfJMmLa6byinNfu3zlm3sR/fQfWXrutDJTMMgFCBveZ2GZjI
dcdR63wEy7VKu0wK0QDFoG3tk045LhLmFXjwvu+uXljdZR5GtZNRIHUDjmN4G3JN
dVqXbxghjLaMtldrGkDFdf7InKX5ajnlzaFBiBqSvWR87za5DCEQIMR2/OE21K3j
TzGh6khQxj+5FMyuo3xf/nSVcj5i7c5lOEgzqKFB7O9RLcfkJYXuEt4wDYWAsyIm
L6+yTEwjHGQqYNAlbG/CzpgkUqVBhZ0SRV2loh9el6r9s2lNM8zgw+IBIM+Qnzze
ijCpLT8SQ4AQC1KPitLXWHKLCihvn+1LYhaqEPRdbFetOiTcVYajJt6C8ehd/NOF
zNeryVa0oHQs4BWX5PTHfU03VRIHbJ7zJv0b2aBviDnrPwAoVgpjYBBksjmvmgJE
1++Xxm7FOyrKCElhOjf107tTNlQ4dcVjTciEPJCkBex7lnkOksOEgu8jbgMBWJ1H
J3erjZYCCQotwI89JaL91jzvcydaGCCwk1gonb7GDtP+merTRpXG7Z+DjeUutEvu
3gEcBTY201X1k+RreZ7gMnRuO6nFhni4KQTU1V3uAmx1eBdftXrTpar7Qt/4YYXh
hzuVan2kOVEmaKl66SgcoDVsQxUgNEbB1OWk1DMJ6qLyg4wW2L217v/GESDDhBFX
oSRWPieWy+m5PHOMLtHNRSdqt9dvUZ60DdKVf9KOqsl/JTYOLxQRwOPDeBwnbnBW
N7h2J42JgeR9rSoNzzifUZVdzJMf7Zi0i0Zj7TfO137eciWX9DYos/KchvKHbBcb
3m5HRlZFpfecEON+IMqWspSsSWq+9LKF/kQS8omFqgzcFVspVdOXfZGnCfCiTQGm
f4HmPVcKMblVFI5DypYPD+DZdTcozBWDNKmfbyA89pAYbhioZuKVueNEnzkYhVN/
O3V28jfWIbNn/JOV+8iFb52fgYsCA3KNdLX5DUsRoXadhwMhFBfItjl0qJHd1Guu
`protect END_PROTECTED
