`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FnLwKRvQFsP3QaOvR8HqOehpiD2nzzsjh9e9BNaKbZgbkL1WsSHheLwGK8faKcGh
lYdT4UP6CMdWpM6v3rc/gOkitMDjPAAzZqoZ82gXH0CptVWh1ODB4SJhwIU57WgC
rdOgSzoq3rx8sW6XKtJyebP7wFKALnQ7aZi6uTn+gsS98pODvFdkAkB/xOs6wSsu
5qCz3ZhX88STCXvkqvUocvYciL1myaDknsDZFn8v8z+vijRPqh92+y9mbSHEv4oF
CI2292Z/zRbFbFuxTYWEFZ53aE6q+l+zKpqIoqos/MvQ/ZBoXDv9F4WmnUrn8NEP
LQClAZhbgQxzCDj699fnhnQ/9v5UBFJmYoR0wBXDqyMr9cUsDZ3VsOMa0RWLCszA
WsC4sW3PvrnxRy8u7QoAmmV27q5GAjRF3g1EHi67gRpnVpbCsIXTse8aIEfDK2cQ
4DZB204jywXVZebFs4dm+f+7HMo+0IfAziIJT5YPqejbo9XnutgoZXZuzgvuLk1Y
WC4FIXC4148y2QptXZ0qlFeRHakO9JJHSt4CgTwn8lJea7r9r8pWlv/vnZH2tnBI
rVK3gYh/fVHw6LBQClEvX9qeOUQT3Zc8bxN027zHsKcglbHuRSdn1vh0JC+WYC3H
Ry9b7e8HlDFnoHBRfOx7lg==
`protect END_PROTECTED
