`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q57dJG7kmBqXshs8Em8Xvi7MiRbpYgM+TepWwyFrr6glBd/uES2G0cKlodZrJ/Ki
Grh0iF7DJqVFgfUff+FjI3oei7o+PnzZpAKVrIjWeXTAadYiIrBC13ffsAHDu+po
egeBLgoKyyJDI9C1stN38QkSHJ+4ks5BYqlIn04zr+3zZh7kM+D4ogwfvYEoeBsX
wixrMTUGmhyAbn8SH1SxTcyhWPAqiyD7uy2wt7wJxBGXg4g1VZiMJ9AaWPipbR7d
1hcac1OaRuqZjii8Rd3Vce5jEpmukluvSmctYsX747tESWhk59I2FLDlJ8ZWjJl7
n/3juB4M0q1a4Iuzr0PZ1aES4mKiJa1sHh04UVSqoSwERm+fg7el1T1O/hSA9Ds6
MTNls4KZuvH/WOYgsETFsGw0p54PnkpV0P6HLevg+t7mfds1A39H6wb8ouP2/f4N
RsHO0pGNih6d7KJTVPj4M/e7ObVqjmcR4FFMF2B1qChGvHE0UbQDYcutUuRMyHo0
E7qEm10tvSXJk7yggeH6stKdejRdMSKxQ8vP8UeveZTe+qJnMonIo+x3B3sYWZlB
ojrCsnS6ttlzcLTa3tugrT8AdKIQqLIeVum9IXhTysLUHYtJ3XTvNQHju19h0IVw
bvItwEBfxRLRDb7kXODqiC2nDrkmsX2gHs8+lKW2uwUNhxN9DR/txL0ZTqo3YdYy
acYnDuUranhYF7rPzCuqwcUArt1O/iua/zfX/FSFyrqkwSdnyv/uL0YaXyOoVCiY
QGF6RpK3IwcI51nY+VIXkqstExBhIi++KzUCZ8hBVHRXyG1XoZsgJZYIq2jX5Djh
L1IOiaEW5j7/tDDCIEsRZemwEXyG2agUsp7gz1eqAE8lotJogkVSpMzNej7JvvNx
Tor68mZu9bPs3vLMUSUb5/WX67EX4W6QhhKERzfS3WWdjH8SwSOyQ7/Jsg50eAvD
75sFfbGTWO6h9ayjPfdjCUX4IzXPqDR8F497QG+wnxomiBt9FYft3tFY25SL6kFe
TOBaOGGsjaw5PkbVehwpafZvnJrnALZGqPqcQziV2hXycL52YvDhciXMjAK2GvVH
yPoqNVFpaSa2wqvod8qFAK6H5dJOU41llAMpVENOuJIlxxMFltU14TZpjlQeJcy2
mgUY57uLc6Gy0HDXAo/KxBGwhkq0x70ZTwD/g55uHjceWLGVkFLwD6crLeUnpcyM
n4pd42Pj/VxOHF6vRtBycEZuV+d0vxtO/YsAaw8x0FnPiJJFc00fOhJfYT930E7s
+Xjm38qiAEUxjsuicOqAsnncnkQyL4g7eSlsW5FTpUwNbMfFJSawBc7CV0bd/jVA
QwOCoK20f21ocfD0FJNrjYk8GbNq8xqqN1MzDZT0j8ncoOhhru2W7BSKh7z+9iHa
kTpU1ntFbnjnuY3w3GNnwCbPCYTNazP3IlsC7EWPBVrqBRHcltm5ouQgufxc2RLj
gOxx9fxEoAbMBYIDjJkbCy7au3noCB+WqFNyIXSf+4o=
`protect END_PROTECTED
