`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D1ZATDomkA7eNIG2Y9xxABeUFmOIIvlXtmN5GE96oBKaCcrsw5noIfXOopEWuBgS
TD4vBaP2z5hEIAAfXYPzFYz5Mz624joD54i1u7sfjmM8i3rXD5+wdNpJKM6Dbd+e
PzqIma1jLlmJxZbUe+050p9Gqde+6A7NWn70LagJXJLlGQkPbWz5GzRJ92ifgoeC
k6XWvcBieMLx179cF2Nif68P75s0f58+CXmPdJa7Slzsk71oWYt2YeqyU5Z6c1Fx
gdDpsXlUS3tZ5s7cRkZx3anQpsaq6//RMUKWcVWbc9oDM6elLDuXY2VpPUGmLnix
9w//wH/4cbos++zaySIyLDEJ9NEl99mRM6cjo3kBRqi2uhutkibfsS9hfqmpld9y
Vxz2oVOh4vq9+labHq1SJzmUM1Ri5I0cGV85nB4+cr9HCY/m7Gxp4zmvmifHaiHU
pOGPT+hkLgnsTRieBIoM9K/lW0SWwYUk8PwcX5TLKimP6pzSFyWknpshsMeRvx3Y
PbJL0hUyj0ySb/H36waJj9Xji+22fcLa+WhaWRO6O9vxZ3OJ5vPB3NqSfnUJtH7P
d2K6Dz/RhiNaLzxMwdngSAzQdQpmqhx9gYSpq6tyQ1pyqkmS2utpjV50yoQAyl82
fHmjotHIhSV5WTpxdCQDTmT3PZbMRVaMsro7iBUNrfo=
`protect END_PROTECTED
