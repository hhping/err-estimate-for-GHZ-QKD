`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmWyf37CEe3Fk7GEhamxYbaoNuGXlgMPiLR4s4Z+wqQCaUm4Y8yGRFuzxFxly+NA
eODkciDvA30DePlRPxsi+r6en26dPkPg0KJzviDv17ZB6PjDsdoT9l3hk0tOfcKR
kFEZgPbpDKjLqvOAc7syJpOPDN7oHOWi5xdTq0puhCKVpu5P29OT3KmIKJcpFhvM
lSkssMO5046jwT3fpM1HkFD66fG137mlLj9+LHhw4CVYB1L+iJtqxS/N/MnmqVXk
YKAIVO1Kj8GVlqoZgFgH7VGdYykWt4KUbR4M3ZG2gMOa7MHK1KGU+fdVlQgeaM4v
lyAHH/uTjIMaSz1n7eDYhFhdVxw0H1L/nASnSGgggO2tRPAmzJVT4lbj1ysdA+i6
zHdUlxZhiyCQxWR0Q5CnDvYWLamAV8Ifzj19boGf/uQVT9FfqEf0vrsH/C8vsMWG
+/0Oo2nO3orv8cZ83FktlKO8RM2I9Yk2PCAG1egglLmO/DF6ZW9TwKsIq+8W6Idg
QAuPswKwQallrHNSE5fymH7tBfiy6XDuKLF6I58gk7fTdg6JdtE/miZHpqVgB4JM
g88SpIF+gv0wYku5XVRbf/lMioRPk3VKLFZJFaYQV5iLAAfOIuNEH6V34phU33DM
KlhUHFlmOql6Lu0/bn+E+DpaeNI4cKTRVXJzj7KZylFx2++rUJ6ODMiY//GpnhBz
COWr6aqbs3eqoKxrJEWJM7KfIC8jFFGi3Lt5JaY7BoX0VZQL88xPF7Y12xNs0dyd
GLCAvUqNHAW+3ehzLkykuWL0LM5p7ONbL6QAVt9omnIQcYWoTtTMO45eLxxW/qxq
eAKWJpgPbGeEasUhuqNYntXxoKt/eNQkUR4NvuxdYQKYpGAttY3hKlV6KMxuMAQa
sT9Im919iLEKG8KGle4oc86XarSBMnit3PN50ih6lWJbcxeiOfuxjzTmw8Z7d29Q
M4VQWA5fMCQpwGUR8GAP8NdqhXs5/j5F7312vvesV3q7PK7pF6Ey0y3ejN/lG1RS
g/ODL0TsnrBU/MP+6WlR+Lmr/pHmaIz1fe59rgUhdsqsJ5sTTxRvQVOAdZU/HFHD
MyBwFZ0XQjlSqU5mZj2W3F4xI7D8HeQUPdcR10pgqGXRZv9jZQljnaEiuSixz/9p
hSzdaFiazlt9e6soj3huvIfG5gClWQstJTjnNfuiM7ZF9b7WG6w3vqKxLK7lJrUC
fRlmqoQghmNu3ERwK3TkOjLrhMmsQa9TUt8aLWfp9L5DTppU35gl0IwY3U93j95L
cIw1ql9Hh1jP580/jSL0H0AIIZulanJ3vN31TN88P4JLLehGfQGn064qLAPRIppQ
LAGjkGmg0cwME9wdk2S9mMNEnbudE0mh912x6cK2a7GaY2Kz8Gxj9GAEfq0bdiRC
QmGOm3zhJoJTCAGzF4PZRSCyjq4ik585bDLLo/XcdsUv6VI9yOWSo7WBAbLISi3Q
z3UACruhbmiR3sv3bkhVbQN4cRWGNIruNVH13d9BNmN7k4IQ57dQIeQcpxY4+Brg
FLAkYlz7/Wjc8EYjY7+HwtjO+F2aJBIbX5VKFtEMmMwVb6btFC0vj/gMbxhV0OpL
Kik3YpwNYYReU+3K5A0MesFcKzaRQcqUWfi3YypzMcJoUpJSW30Xc+XoAeR1px8q
nALxtazg9xYhfUE8JaJ1w53Qq5bzqwURLQJAmNodklp8R2EJNvGR6cuc9YtrAZ49
A8ccymixUUdM1oiOpfvz9SDmGFwHVPfvSDB3JHukDoh5gMgY6XDTehk0WgfTiGWM
sBqeWngZYFF7ycf5gk0a71bH3F+HlQZTdfoWhaVtL+/dBhPq7GU20FvaW0nWmVhG
nyrUdD31wmK51fAm5I8UdMZFjhPU1caGdZYHFGq883k4pW8wnKYnegZMTnCpV7fI
Cksg49cbnvZWocRfk+lbHA==
`protect END_PROTECTED
