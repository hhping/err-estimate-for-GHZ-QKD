`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNPN0k+B1jFTxBeyJD6zWXDzOxpEO5dWgblN0/n7i1Hsw0Z2ZdQunTiQNdzQozAC
A+iOlnhNTel8Ly9xALHQqfMfHSEYRduZKsnbs973NQs08fGT3au8UEne1g07G+Vq
90qdRmDNBLBInAEosdguNMpzh6qhcnqe4yYnMiMLyi3AIcS2I7yFVhhbf3mo4LzP
Ijdzy/euWdxzlCxh4J5n6ZlnSIUAL69MnzvGWZdNxGYoTRPl+B6JkW2MfHqijj3b
1TupydL20n0QSNlGyjtI3BHm4bDuVFFmV0553alcSxfsw+Tghp9yrD5+AOe+6xt4
+qzZitqbChiRlMoCeUdowqyBtpqILqi+H6niCxoCOa9TTheR+pM+b9CwrqVJQwRn
ZBbHPh/4NJeiwVBjQgZDfQV+U7zS/6mW0J4oibvMThjLQIslnhxJtUKMy31/ahot
re1mM7K+OhRmoLUGr5FK5QGa0dC6SFaxrFhJWckS8aN5Qr3zg6bAmN/MgmdtBLU7
cknSkdkHAYEcG6gSZ3nE1/kkz/PAj4QgQJWPzDeXJ0lB5kOsF9Sw9/KP7hZW4qiS
Z1E9Vc5PmA1XFBkNjYZWWP6+p3satQcUAVLeSTgjiRCgiLrHhdvYKxE3JaWPLAYu
OkH9DBKibeQVKMKNiSui5sXSUFnRwytgMyMuzETkl9L9aBi6XrD6aqEDY7k6heOA
B5Xa2H6SPhDj19gpWuz+jJe/JxSkwi8eNNoyB3eKSbTEyNXEfsnmEujyE923goAQ
cm9phnMcjqPdQT8laD/SYrKRZb59q3TeBvlBrwguRx8aPl4VzZBi400kEahbUesE
rFL/U158lFKf2bCiCTa2cAALRunFFffhH9vTxKgE8VDwSmpk7C4+2ApUQqm88CCz
tHjsHKm144xwp7oGGCi89C6q8IYRtI/FuWJu3ujbYPmBoGmFvsFt1pd+SXVkEZ/9
GJyBGiYx+rAWNi6oWzRq2Mg0QrDKCGYTbu65LbO2j5QEPigd9cmFg7+PuTcRmFUQ
XjBFyF6z29jLZMA9+I4s+dyy15GauKc18l465AqRFdQ1Ycw+yKB9K2yoMML365Du
Si8WCFyemkzPa4MN+bZbANUqRK7syLlzJ3/Mh5wGN9xm1DHT1f26ggLatE58IY+7
j/nebsErAYoChUNJI64vSM7EOjJEZyjRNs/T5ZtB7f5fCHQXUrkq2vNp+cSX+Aem
GQ8GXXyr3xEE5H8jQSdH9hxU82RZRq90kkb0Sk6PpR+lcYXu2tblNCV9hOzMNSG4
nak+US0E1V7aKTbwDFZOr3dVaQPLFJw7KHkyF3+60jTb5E1YqatfZV+dwJkiTfen
VRgEVDp0ck00QfjVR5Mst0bX8BmViz5kkqi7WyQYqh0BudwZS2aMZEHdYLrEPM83
lVLEkHFpO/psN4Vn83ONL9A6NogPi0mofv+Otmi4+gk6njbtseQ1jOoRedMJDNgN
fhClP1fH9CF6Ndz4XwWXI5tHfiHOvhdw5NzFdXrmGexsrqkMjQ/i/ioVK6BYNaHm
s+anRkF5t0U9A7C5KGekycevT7ZUI9AErKmvBYzRY4e5Su0u3wKrC1oIDvGrS8/V
dyY6mhRfVFZbX56deKszrbQTbitu5a6EE6aA5evEYt/FBeNFWnmXxe9W9hO5jmei
AD468WlJqKeToSm5d5V5dnjl3DADbTub8/PlDrfvI6duVRktBG4szRDbv/7jN2X+
nz99KNIy+hTvUJgSEqMHzpWO/PlrhoVVNgI/0MNdw2jjHuIJMMLuKfjFXUYlCeeQ
eUzjUk5iHdK+9EqQHsCdfayyDInWckpOX4PPAkmp2fu77RztoHC86qgfRCSk5NTZ
RKVJYX3Ge+AFueuXujQRz7H7qMiH3TtLGLGAl4sawh9oWf3H16Ej+N2ZVBc3Oq5I
h5v57Pcvc2oR8AUHXkgKA08mYc70r9gpE+Jq9zc+k+cxvuQ4/s3WCdROINjrD5G7
AE2F+SltqVaT9SQGaCWSnqU694wH8o+n+ZlSOgf/I9SXeUxNujLsfdVaYt30HJ+D
8X6oJMCsUYI6xBmRXk7Q1UAy9HIH8dZS8NO4OhBwYRNqRyLE0laxR0fnzddghBjf
7UwPzoQJ5PlQe0t3oC1OyVCGN12PXRBqQUvUq43kvcszo5I5+/rxnww4MQeHpak0
eaHDMWqs7cDfORSY9ZvslYu8Kij3BcCQCL2QQD6ej3/8Em0k+WETKKFFTeGjeTV+
i+Fgj9hZKcL/jMhVqpjlnl2pSc49LCHQHo8xNiKov+JgFLb1Bzi58YEz5PznzD+R
DMInS/YEZYXCVo0UiOt8wpXEMJk/a6f5+zGsWey2vxxybQSRfwouwi65Z3+lzBx8
3AHrvZafEvFiCkm+AAY9peAXUorHIHyz403tyunKwwqRVPWv5xV0XtyBGihGqzMx
u52aM/BF16a8ut8dyUMYBN+c3QeccBCKc0V1PBrI0+8MmQLhrLXHmsXip8FNZgL3
KuURBelJRqqPw6TidjzWASET0ubjkOc6AdypEsIA6FAsAg+EhV+L+7WmPM26iNAg
QBRR1lHSH4jBYfXxUxwFq7HFb8ecmpMgao0KhGd0vyfV4/H60EO2McboAt1r8M0x
w8ig4ti4i1zTWM5ZjfQeN/MxAxTkrtDSKRH5sklbbK2u7SlZ7w+zgkozJCFcrnSc
zBP+2EIMkTdO2n2wmjKklK4UzdQ7wkYs6xu/gh7zC5fkca0yE0y5QSAZ1ouSSUbt
Bl9R6BMSPy6Sl8Na/U6/vGGMHM7mMCcaXbL+dExuNb0pHRhHhRu2IxOWt5Y8JsKA
wyWiNhLam3aHYP6oftRtgT4OYRKF3oYN/siMzErQqeGpLLevDeHnAljGXdr7gyB1
hCiFvalmPx4TKmpzo6rSNt+IWKllGjPx6LyNw906pDYEb8OqxOjK9PBL9NVzYwbw
9QjrRydQoiV4CkZl3y3Iv/yQaDMztwHMx/llSp96W8tfUH3Z3ssa245l8a+h06ev
9ILcsKprWIxTxiIelWlJNy7lOw4wbUvyO70IAftErbPvDeEvPdKRkXTKcubi2i7b
oRCHN4NZrI9ISOzEmXp3haUjRMxGo079fsZALT6qf91dEHV2nC9u9PzalO2cS2qz
N0DxwTw0yViqgQUTT7KMo1uo5+GvC7FtxZ8uBuDsZX+Ic3Wvf9ba96X6euJDEBXF
lVJROHY1DXq5dlg0uQQJcjDok5TN2NudKvWX0iOy20gSn0QG9TY/Y5SbnBc2BCaP
w0GtFOkYbUqyeUysklBxRAHjHlamlxkQpzCjx4pEYtFXnr/PR3MTwmiYyfSh3eFu
wv6/vMc97w13jLxKXyo2awaMKYD0yR829t8gTCb25gQwLZVy/BySXTk1bsbK25I2
k/8F5ZmhNDV+gfHLGrIZMaBUEMz/Abawda0mIAXgBymImF4DJqE/aoGXkiT2OAbU
EwzPq/Iw9J+KU1deYvFQ7j7N9mgLsqoBTybAm5XLVAprPnHAswftMIc7lvz96N+y
ViHdZ1eSFYARqtcy5/MNQLHCq9L7j+EnmWmUD6sgUaXAGbiSMoMJJVFLUcVr+my8
DnQcGf79vG3VO9cMNHHPxW6cfgBCNitgI3zgqAma4zne2m0WaDOzLr8aWnzd6gk3
D62LEGhZ0DkTJhxQS0JGxgkPWCrih0uO0MmAAV6AIC6AKkmBD3RuWNtNkc7rnve6
JMQWncUMqDCw1dv+PMVwbiYDah+w4+J5Yr1NAWisl9I1AZ7kATguuod0MXmYP4wk
+rX/nHX+3wE6JChtHqe1ZAuvIz35rSt/ctkdHD6Bfi7KvMgGguVApGq10HumyRk0
MW704DNqLN7oC/7yQLQRQ9VbQZ+Pb0xsz9rGArQUeLk2bDy9FbsV6+Bdkly38lm2
tyDw663SaQtOol8wt9gr6qb1IM57Hn41dbYOtcNlRIWEKuvDCl8cNF9bBNxKiYaK
xiCSu+xJEUUEzPFeGR4njcSgRRh7BAVoiGR8+H447SzFUz1aiXFueaLhDNyJXZsq
8PICDm+ve4OisPdvWGmh/rTXScDp+3+w7R+6ngwYKQKXzesPEEIyiTcJU957hWJz
8oHDdjAQQNBBcCliD8Kjt2TuyRA0zI1BvXick7QnpYoHgGOZ3uUsIbNOkAk+SUij
rhJUfe4Bs9y8CcrcFb/gtak71q/xe6AtaCYNcotQMHcmiGdVNUmt37y45E0MU2+g
+5Gk1f+bxwNIRR7X8F6x2eF4V5BQ/lRK+afUHELdT5vYoyzf5gFnFDEPSMil8jIz
ETJ+G2/WBbWN0kGOOCzGLx0lATZB47RxXcMMrk3667T3qIlpXBTzGN8RkL/99IuT
rZRQj4EJJ2k96RUaMCOlhLKPneQwVanKuumS4XoqWR3TMNfJMohjP1FOZiQNxSut
y1TjkFA3ZJ9LLanm56LdQA6Hu6gHb/MpaNsB5z+KZzQXlToCFUWSFKshwf287yb2
GCOKMBxiTNMgPy52G1lCNaemX+JhXjgOPQgWVbDPH0cwDFrDySv5n6dvcBGU5TSy
I6GCyyVWjfXin76Wv4h69Em7AyddxCuEhCF/Ko04ehUc+VmWiR4O1MpXtHpSdZMK
Szor/kBPf6DlKV5jyqvsIONfNavPTlthTrXwr8xL7K7r/Nzv/ZOhSI6ivbqR6D6z
WNKVIHjjlupbSpL+Zf9HW7ECRePtiR6C1yjyVvg+UpBbOEl3lJt4Jjvw+KUFUwri
ykr1GqlUDYasLoy2LtoEELQwHwxW/4tHZY5ZrlcvXtWdZql5WREA9MOfkzv3NR+M
l3j4xw2+Z5AktdrpUN7SEbZ6NVF9vDjEw7Ue05lcm56xsvv56EY/C/cOaXSO8oQe
ylFa4tOkfp3vzjgYy0zztSBPrCJjjz3b/FrwuM4OET8IT3fibXcWn9lGQlVjiWxZ
Cn1+uiHc+uE0zkXaTOnk4oJtrpi9CKHPnaMv9H9Ktgb7KUD/aVE4IqVkDQhbLyIw
m3jVqb/T4qEZyjmlZ2900yeQOMzxgDKY+CRlJxuwWt2YoGodvDOrOypAQYGWD6lM
QjaIpOO2NbLBd7ftRsT8K4G3BmNbMDVDKJ+EXfZlZ4Dh/sEm0+XQ733GDTRzZNb1
0gHUq+Qt+fHHeOA5iapxz7k/uw/WcqAedxKq8QaGPx2MGlkNpLc7p5GgQj4H9oSv
OtTvY+VPQoqMUMlY+11VmBwTt5mY5HehVl96KiqTQ2pXkUHYVnp5PjtOBWUt0GG8
um5qRgSqJF/3d5kKH7FShmSWOpxnkXfW+OUW05Sf0Kf85szC8Ui88LdW9IFyTe5N
j6KjfufLXtBvskt3dpmp16Ai+gjE16/lP4JG+4EQbWH29dkCDAkk3/PnRIABdveV
D06YgtLlQ7sR5cZYktyF97h19tVO0MuvVPD3cxRHsxVVyIxti2CBcmq6cCjmg0gC
fTKCyAlEYkBd4ZSPlV5PCvBOdLbCXcI0pnTMuuKl5E6DQH2vHnHUBNORp1/nBFMZ
Kmt5gQBZWORa0+g8DQTfmVRH/aGVlNaVF/6K2l/mEpcy072A+YEtX2+mJ0O4smIO
gLEt4C2KBFf92FLo4ZC3fNpVdWiVzJjXmwilPD7f+gukops0TjzaM9hO1zie3TKH
f/WK3ll72992lNRzAwAEDiXg/z5HyK+UBlJ2nA8rmjyww9ciYicdt8FE1hxOevfE
zU4DOFymowxqDYf9A3UgsoVnzQv6djxNVjMm4z/ZKiwBa2xEddCtPXuUBQ2++ugv
6Sl5TCEPp/R5APdQwEMD26oTWZRFBZTx+atgTv/YGkSHbiHfzcBfSos71dJj2fUn
Ts0Gwq6ZGD3PPoNmMQbI60zy2coSsurMBJDTeFOKeGzZTzBybYLXTcWsqzmn8L1S
xbAVfcsSRpJOVnzIkBCRVzm+RwJwrqHediFR3HUIBrnRb1toF5NJDB/3K8ZtWhVR
EjRZbqysmDCbVvDl57qDQCSaEmx8TOUQvQLqo4zdlcVRVguouYuwm3MW/qmVFIM7
KxIDA9ZkF/WbE+rXg0WBRZD7lPG+8LQW7c9IvaYDyQE7ES2MGJQa5Cv3kmOKbfm6
N8mUI4EqzRfYQynl2jx50UKEpKWiVsobtu4SUXl9bC1mIADvjlhYEX56/k56sEgJ
QalL9z9qHmFnY2TS8Y700YZajiFxcXyg+CjM8ydAm77PfqWwTkObGNh4LQ5OgriP
2EKUHhle23+cedJfnASZyNpVShHlXvkBpL/VsQg9kHBxZ+ZXjT468cXFrdYRV7DC
MxMAoZjPWLqqVJPK4DY1N1VjR63jQNOrBu+0F2FR3joqGCwFMPGa7DnyfJIRNDZw
1gS9TLJL30gBtvnkUq/orTGYevy8fwzUUu1elLj5rVZRFc2wO/0GCZwWgkCOty4w
MA07fIN2y1ENmIVtT7dTkRALkJdI/BV8ZVmhdnW+mIkhRVDNinQmXFv9khdxCc+x
um003k/TjVtWJ3s01UPieL/Spc1gtvJHFFDBOA4cFcfCUaLN2LQz/scUhjZeMBuE
ntwoi4ZU3FmxsI+MuXu8OKddWLnpb3yYs+Q6kSthqqWX/75U0IiqgGagsiXF5v+Z
NrfK4yACm0cpkM3uyjAipGvDbsGKQEEjWk47RsKBTliu9CHwBaFxA4CPXXXW8YCf
936gBDv/d9fr1Z79AYpPnpaWTw2HXkHXTMW4jbOWhGdUYnGklEClMQjheeaT9/8z
fLKiDvfdIQesWfW3JbDxw/25Bb57bqng3xg24ZyEeJ4PvmQLSMTu2Us19WtC1i0q
seXrxBLfocUiwC+Z9wSpUZ2OgiAn1NvgwLSRjSQybzXZzGm3LTQCK+swR1DXjU6t
fIkeCz1+2Ke8DnF8Og/RCfADygU8bdfBznKkfVKNVwyZXl645VapujKzq9Bn2YQn
6lLzzMDQtUc/uQjongTdZGLgR7rufk/09uNNUeWHW0BCGzkW5+EAlN9D1/ol7G/j
J9/KbljdBOj5CHaFhQy5bekHDXOQE4HwY/1BDOiNYF2qFlkReoUD5I7pp99RDR4T
g1xmFbuA/5YZUGb8QuOlHoy61wz1LCpIaXBB+GsLCtvlLGIHYFT6EwROpBZvnag8
cavFUOcMOkl/Di89y8q/gKjzaaT6BpCNcFxXneoJO+T2DJH+84MYBU4gjNjoyrDX
LOu3sD6VhwyPAg6ZYnOIGwDNtKNHvvTALh6zHFO/XGYZiovJQBUHYO3I3kjCFujY
vXbFLLV5xSBafP3nUN2ftNP3Txw/OIRdvcWf+ioJ0IHoRYc8H2QLLI96IiYPjt5U
0zwXa41xqMBJ4L2X5sb13mdICXXr0hk6inzNcoIQO46U/8oQwiRFo2JrfgRVu+N0
I9EctRKU6wzyEtQR+aZK7mpaj2TdaiHz2WkzONJpb5wPGP7TGKwMl5i5oHttmJfK
BSNfRh7wM4i6UAMOrr/v9xBNSx5Zfjl9QfhsO9Jp/nby7jSV+PvgoYP3o6HjcfXi
TFqPipMPWQuPZjDdzd4FHqHGTr3Q/spHZAmj4DdldzKQSkyYB5nG2GQk9QuVc4Kn
7cIaqxvHq6ekajuLALCiG4T7y169HizNj0tofxExtOPZbIgz0KqKd7WxdSHBn3DJ
SgwWxGddEepeLfI3vk+gceEG5Ndgu6PgPMAdCdclfmX0QsIs+GQ46V2aT+sQgJfj
UVi1EG3II7qmTruLtIcEcJ/8MEWRpNTc901W+cBh03qgOVTcxA7846TlCsaXvvH6
5VJc8zJ2Ztf2RR/Cs3T45C07Y2OlWzn22nfTOPwF1cJVT52P+R3vomXxpUfbzI3B
9jqtOrFlGS+CD+GQBQ986LDJ0QsDtbU5G6MW+gBGyqagBr6JmQU4H03uiCD+rhIq
JmTFmmvPRbmWk2LUk6ptkralMf38j7KEnJ3HNtfBBJfaixlmHySa3brjpswUEdei
CckrRK4ChhAqISqmSaOxfFDrurOKIOVK2+BfZx4O0A+a9YHlLHXH2wD9p5maR9GH
GzK8zwq2VEbGiZ2LipYV1uBrjh75ulcqD7IrfLSv/TQn7mpziu5iIMIJW/WFTQnA
VG+4N389aMdxYr/l5+A3vIGvnEQQ5eNUTNrgGmLEPhQhKwWRnoHNzg1hedr8LjPT
HIW8XwrjcbInDo1JmdoC39d3z2Ozg6FtEvL6fRctZ/jpzj5+gpsiBbNIRBrD1C9s
53UKMDqCbDbgpKsO60CKSANdXON0nCx72smtzkA4RaPXoghShv6uwfovYNcwoJ+K
rs8vVqYIQpLGfFtbFGLGDE5Bmh8Uh6/KMvhvXYwmDximxZyLlpeGn7rVnjAYrrtG
aJPpopa11q6t/TvezNnM3w9k084FaZLxw1hMXVlFFE5sX25MvrQmYgC/SdBvuPh+
QwrH/5gqFE1FLcrllytgh8xKqj6wXRP6dDvMaYb9oFU1juleX97vfyDCyy9w+4Yu
OqF1NMgnYC1Dwjo79F/zpmYYDr1/C3sBRb6A3Jwp+sTQje78FRJHzUGNXQbUzDSj
NdpebDCYA7xBaBzctbqlI4dufRe0IzatPjhEGMyxSiV+ZQdFgGZA9nFiWTxDzQda
T+8t2USntvscTDOr1TKd1EqGdjHq0H280nEZTKcHMVU2eVtGES8A4LMstd2QxGAp
rkqGbcJAid8cmI3vULjUFihOtIYT4RTVzY+/+hZ57bp8WftytPUPAUiaCfn9flKc
7oBLlMs9o3P7fxqgVHZa07vVnE2no28PYqcnKghl5avJ/m7Qa7O49FMUITFdMXGM
v7Tc22gaz78yqdH17gdnT6f6Dqo1qXT7afMahC0ptU1+uesymy91qh8p9RGVGQca
NDmb+19HK1lVJt/fPYI5ZvY1hhOFI/FTjGyuVzFJkNMNH44+O77x+ihnm0SrTDZk
2O6R233cQm5Zo2wbOBSN6cedCrzIyPJr2/8V+bmdr1GY1u0n0UUcHgBi0WP5q/Ys
qg3jdPQEeLZCKIED5noosvZyKPTtNb9vhGjD262Z3UHmM92/gcip9UmXrhh+1anG
3FY8uAa86ScNf3A/f3IkVMj/5RMM+badwDUJxPQtJMXlnKFo56pS/GjEC84ozEW5
1aLznBRx4fB1q1CLBLfZB0Eafz/35U4f4cSbGwUvaayLhSNw/375e2KmCb4LDHF+
LYpWh9+/vdrz8/S/zXzgqG5B0T4r6OIqJ0M7saf07ddoWtbbe1hf977Z+UK6MUn8
R4hDY3GGTHD88Lil1IfTMV3CPXMWd762NIjFUqbxToUD+Tl/ni/B6O1d8pTDvavU
HTLEXHr7v4YTdyggxCxeLRg/qIvQEEyWM6lujoaPa5rJ2GBT874eubIr+Ev5x0s7
aXxUmU/0NJaVTEp+qmaRQQkBVbPieFQF5Ep3uYe9654a4ONF8e3I4dFcZnWaBFv6
q4yu/6azmfQF1NQAF7bLk7Iz5amXxXbl/ByGDyNQZxi0qXlZLqkI3EBkUTNvsjuY
NyGcGRG7k8XHo8Uv6DYj3H4BraIW2dTVR6bxReD6uZIIU+W6r3F7YFrT8o0P8nq6
CO2aF/EwG0L8qLRd73N+jodCeHo1d9mpufJvCZA0kIQ7Wr9+FJbOCLOuz00Ivajl
F1+pXlxY/+cV3rDhNykJtrwMCU5Lg8aTbAPUtYUoLPGmwsIztcszrjOFsY8qOGuK
PF7x9L6WoVCOaPTQuXCkoLVxFQC20/ecK0NUhYmJRyyJ9b/9tu+f7fArODe6e1RJ
IMLWnTU8ykB0XZPhhzxlqb6xLN9HZwyIFzAuIzi+W4cAnrHQPvBnnRq2b/cZT7Mg
bMtM+x5zFLrb8PTLibLOc6br5z1vooZBapu4533B7bW8cUc+dJSz4E8IfjRyyPIH
TEsRRU2Mn+jgg/mUs/L/5QYJ4fXno6/zVd4QG3FV1OZyQoJ/XCeyr6F6W7yEEzu2
IUqOKwDetpBxlTNBSEr5fJiLB+9e6WBiFlatL8BHnIvxaxCN/CpAywrMSO328P17
CrQxBm0FqxaZUBEsr2DVfFn4zIacPT5ndqk2XoikttqfyU1Y1N6qC6IaHyyibvCz
SWil4ZseCkTdaPdO/05bYXpxO6zhlwsVjk1xuQ2wCaKiZT5j/VGfirjDD0S1Uk9V
VOEtbryZKAc0Ch6dVv4/beXjvIyM+n5AQLjqx7Jm1gM/1D/xLtk4SjfjBlUf27nV
Gu9g5w+bxP17CqGbluO3JrZOFb4tAZynetGVKUs8Iz5D4YURCv3CcHR41yP4dCK8
NAiooIkRfiGKH+ef2+mL+GxX/8erTfH2E0AfGi/2hdJcTs7upvKAVs7fLdp/AbqC
HOlr/1pYUgrDvbOhYuTK9A4zG4tCeUHVdUrtgLK5GBS3i0z2IUszOGIj82JfeuqW
lgQbBqckoLI41rMnHFozvv4lNRPXUvFDqYjf6VwCwzv+oyrYx373pMqXrUZswQ9Z
iUhsKOD/gtU4FtjZhgSsdvwxnbLwstwL6Ffxjd/SqlewSjY0wuUVwPpSX2JLWVy9
SwPQOvYmFvEAmNpbERcqE+Cb8Cqq/z6WuocD4YRblziBH5j0Yr5uK1Ffl/8O+YSV
kOXuUf7RmaGahtcoZng/0o5s31sK838wWiu21a0MnkoHKZePvlkPdfmSwoBmfKbu
TlhHQHLmetwyQ/T7Mu4stB82MZV5wTavCotXfQa9Pe3i9zuWfHGixz3PKlzvCtOC
GF3KYSdd7uj+x0B5lERCAuztgXKCxlYMbUf/0viRDwntvMtVzUe+NsPtuJaAyzOz
U9mn29e02Dnz+z8LKf8+ZzMHxojoe98qxlj+bx3ondDmx3SeBKY0O502gfl+l3Nw
m7M888kvJjuu7sH8sv1UZTSlUWhdFuv3TKpxveElODo/ceuPB+2nBAR04zoAVpOl
SP9Mk6ceGrBReL0PcAMQzjZR1603d6xiYZql7U0UzGg=
`protect END_PROTECTED
