`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmXrZRJ3W+40ZTOD2GSfwLFjIzWEepX5X+HmKwDwQfV8urmaXXsXdxEKxku3KBHo
6qqN+SD1nEfVXXKEeoWOAkhamCu8lVcB5od25lmA5XsM4be9WzLULnb0pB/7xn1C
12pCsVLyojFcQgvgW3xBZvIKQlhy2OiV0AX+T4/OXLKkNNT7IjcPokyc52HI8gmX
IX9yhhg7mYxjiN3BwWtUGQpnSlmXrchcQNxQO9nNnGnwr5FpMpmAMveMMImHy/gz
IcmqsfQ7iKuVDsnhOaeUReXXei8Q7urEGsg9enIkcuf0ELl3YhgUKgjGROWHywHY
RYfKcrTqFx8xQv5uV3lBNom6Uhvfhw5cjmJZ1LfBXhhPG7iOlyFNsOF1ByOVPxyW
/zpHDk0Lw22NVpTDMOaZ8+620cmaKNY/RWSYNlSRxSx97kzdcGYnjAbX/LvsNGO7
wfZNXRoJRuKgMdZSy0UJBCY7bRHHe7EGmaV8x7OCacVwGj2Sg0foq25rsbgYiz6k
vhoVANL60Sj5IsejlwuJenb+amaf6hQaANoH4h9sXoRkMGYwiUf+uXt5bDp3dM8x
UhsDGfBD2uqAhwVPAIkHLmLgjkBl5t3yVL+hWms6YuqP7chwoa+HJlf7yx9j1xls
PMF+wDRJipez5PJTcDOdnmGCspR3ZrvONKeHXUc1qCVKWQo6MyDODceqtIODKA9s
M/T4LPRXJmG8EgjsdBa8iG1buX8vKkQtUYZlAT+LTpSkuPL9/NDwrIfsuORvhxcc
8wacqfepD/6nhL2/alApVL4kLP9o6CEq9DJhJbHYc4/LGQYgFqk2QOEedFIu/8FN
hPzsyusQR51C5CHvqcWuEwaVL7KD6xzztWk9PzEIK/SvSP21+6TW86IQ06V1cio3
1ryrrZzHxU8D9Jv2GtMTJeKtBOrA296KFiSTcaIhvXFJhoWDvzGWQHqkqahEVVDK
wCI/uLumU7c9fOT52JRqB1vcQwlgh1/k0lt7vmk31j88efksAKMt9mtA5hrPw/wS
yQnYUKU8dpc/nnZpXyxmGxkct9Q0ZaxzqjRpFqYb9x9Ag3rbrhHNYprF4ZKdLNEU
YXfjadqkn8uvXuLDa3pKfTZGXdx/pDa0XXE17wHPevQsCOFwHZ72l0USGcu94DWi
MnNO0l1wdb6gyG8K0vXe6kq1jpTu5ZHxVoWoaOU0wCuFL+jrSpsEbVWJe0LbEaz1
AROBptNr8G9+4Mxpj+4/xWZdH6RmHM9IwCVviuxpjg5vHuE2jtxAhVEn8qLDYE2V
zOOBCmxESRGqmgGc3pN0lyCZvfF7biYo7ob9ux73STzFpPaMYiXXJPKHAfTl6kF4
Y/zdeWH4NLBj5lL0z0WfUz4jbdAX2W47QbKKQolFl6QZjTy8GPuNZzTechMTkilu
Iz2hceY5VJBjEjdCwN6GjldfI/kywetNm852C2EmZJA=
`protect END_PROTECTED
