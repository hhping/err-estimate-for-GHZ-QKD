`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OrdiaMgvaLsZEkHazvExui3KS2z2HzOe8to7GfWD9RZTdngiYLTScuZ7OIOSOap
MhajNWZIphQliGVjq6AhoQaRl55lOsql6aVmwAzPi5/w+UeJ9kQFxG7kDJjMZNFQ
jzsBoT2CAKQL79SIkZGcGBjsngIB/4tbH7awvNB8x7Wi+vK5iimwH6w9qftruitx
CFvtoBXapom8zvpKFtZ/9o6oZ4fUxGrHfNlGozbxWUJUMTDKnMtXbgon0EI1JlkH
MQ5JIG8NWlGA8z/KyWcbO+7UJP/XAMYNNIbTrGp4rnhxm/+Jbo1UjNVgXqbJZJBj
xoZIvZYFIcAHIZoO/IBv0xB+EUJzvArqb93+68aEpxTstGFkk47Zu+N/PUxO9Avi
L4VW9x/U6fuTqvk+qqgSzNpww/sur7ErwDHkrAPkAjqwJFn5+iGNnaeW/b39zf9O
2XbUjMIl2ZkSbU7TG4CFSSvBaF3bAzaRftdkba4bMUN3+zIz5k6O9GVzu4RRSL3N
wVZDx6qUUxjM+tZo0dd0tEU5NNMXsGa3TDj7odPO860N8ZbPpH5XNRjzTbFR3L+l
`protect END_PROTECTED
