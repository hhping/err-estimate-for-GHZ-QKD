`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvKEURtjyistLXggtnlT7aETFrjoO/3rvh20Hh1k6FYYd+5RzzCgC+6bOHTvLAV/
7jeD0xlyYGgQ9UiU9msgcAh9VwO7Z1c/O7efZP0ud5qMpSauI85oaYLvLslunRuu
xzquPmvkbW6R3tNPKNUk0CVJ8LzZSHRuL20bEbsy3DWekQzCV7BWL/vqbpypbZiK
4QaFJ12tqPA/evXzon9xeY2vGg93wJsPMURZBvupzQDGo9MMB1B5/mQm/McvPi93
zGlkEOfB/vpJgZEeLtAsV0u8Fmgzi2WrZ2tcs7rlqYbStAFzapgl82GcO9pENx1E
50KbqxKjNpi6ZyBCGZhdlNxocjTCdwIHnw3BJnfQSBLw/zt/aOi5b1tP0K3pU2Jt
2CDpAg+pFgPy51FHxTECaww5zKU7DJ/+SjX2ITguWUq5mpUH98y1/RvjmEVu6IC3
yQ8UZPMTxyJGxDn8RNvq+6W42xFjA7dVNCY47xkeIS9DrCML8LyVnqFi03R0Mj40
Qs5wG+WOdnUNRZBukKjTQgGTkvK8Y+u2paqvdHEXG7MpQVQnuEE8PRBtXcPcevsT
KRgy1keMk87MK12sydeLSpcsitJtUzYqyozk0bFGtR7b04K8zY96WgN9MWbEWQDC
R06fzGyMVUkbpeeQ0/Qz5VV/KtGbdrmrMhxhFrrbn5gnDnPpnuY+gTCXgqU01ULs
Kkq1ihbsiAvSZvLSNqaWczhRUh5JTWFyanp5azN2HkXjvZP7eI3AN8CHQ6ITKhsG
8a2+v88bpTrjRp4sXody9GU9+FplFVlRVWUZd+kbckTqgXU1AfHPvWCg8dowTD5m
wqUO4eyyEOUbrG7CA2Bd8ZxRe9WHjuoK6pUMxwHHo90GXz71Qs/4Hm0RVtpqR4th
91L0jb6AY5ojHBYaKWjtofm2+SZ80HvXY/d7Xo6MPYM1TUz4Be6tEJmicbMQChdG
HxkMPr50oOMDPTomY76t/bZanWoYGfLJrTCj7hOCJ8k3mk0TYmBXc8OOeEoqXNn7
RIqKSGSClCpZTnTFqWQnuboQ9e0mjfDg9Tuu3rY2IXntMxe0VtFLw5XINjML/qdz
p8s9xz+JPHipOmara/5N+Cd00Di9p8pWjbhgli0R3YpBJz7sTSz8k506niQPD5om
zN/Isn5tphfN2kAUFvOhDJdeTsHrfc/8xMjtG/nLhCuApbaXfS4Zmyr/tSs+QKtE
IvwZqLVcAxxWZgt20SfCRWR4CdeF0d6taluR/gq3nS15OQd2ByuB4ZBfQori+PIz
fdzqZaP9DxOEEv+qHg0t4MCaBn29btW49DMmj2nHammA6+yUam9xO3eJvcmde6Rh
JuYds95xgCS88PN2Ib+fTmK+9QxyshdR2SS9gmSznwuIXclv8ULTsqEtDPOgE28F
Y/u4rd30MRqhX21HAwwQ2lUD4s7YIn/j1qNdS+x99FYR1znmKwqtK+nrJF3g1x19
VwrhidBD5JesOE9/qyrCrA==
`protect END_PROTECTED
