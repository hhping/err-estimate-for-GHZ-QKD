`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bI+iUKtjri6ixPgRDg/dnRsogpv4DxAaJRnWObIc5xnF74y1sbzsqKPIrma2OQaL
pS1YNesXZwDHqItiUpxjTxYPZo70PystM0dGWo+5dpv4F9xsDCkl1REumoADlQZS
UzOzQJPxcqspX36yDDmFrrGBPVwq54f5MmQ8fvLqjM0TFJshFeL/rLnxtfih2gOI
Nc6KmB4r2+Yqt2E6MweFk44lfH9V5i3HdU0rQe3pjbPGheM3XgBwd3XpW6RmT5eu
JBDLoHeMJC8QAV3AybSkg+fZqN9AiaFyqNz8IgmYPTiEsvrOsN+fpSifKwEQ5Lji
JomiMBPPafiZ3vLeURYFC2uepWyi90k1fIHrXzsG2Lw=
`protect END_PROTECTED
