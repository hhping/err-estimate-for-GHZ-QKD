`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgLj10BlLFfPJP2mKHGkdPDzzHg0kv8ceE9kJEfJMD0VO+JP+wyOrtoTozn9pvsa
hjLf3z4bmuTMU7p5T7ifbhJU8hWPB4yDszcdvGUfACYzyIrvoRe+wwyd1VqOJV3u
NoDiAJjfbDV3GwhCFSI0HgvHOFZkptNx+mKJL7M27LoKSYzLmwO3pWrHR38KTD0z
J3n2Pl2Z1k7b+kMONFzHfaJGYS6i0y7LZU+szcuiguDA5H4tdo1HlmqMAL3Rcskw
kSTNT5z5c+ipzMVKsgkNE+XVgq8s597RQ2bWNuR5F8Uz1HllsTBw6VoYzHUS3X33
fyS+j7rcj22LVbUhVKoKnrJEWufB1yZoTbBS5H9bA3jM4/mmOVHzxrXLIUYxFLI7
wLX1b3Rp3FxfGpejW1s9QM2iGAgLCM4K3C0tZ2BADRYSJwybE5LAf5P8W4WKFwE3
prFZyUM0RbVkRfiHVGuIDwggXFtYEBi7I0t1g/wO5q/ZdmeFLe+ma3yJD1F9sSYu
aOpzNOMAPmn29g2m/TGJGcvU3Ns1kJLymygIrTnkJBtUNEs7W/MNJMNlxdgr7Uy2
bl8/w5fKIUotd53J5m2HhW0yn4qp7LRtwkY3ydrDnGP4XFWxg9VlPj/KHgab5rp7
WWg+rFjcTRLW3j7cBeKY89heGZ9w/GbS9M9Uls1z4jC/GN+xsJ9bKHWyAAxD4wgs
FnBq9O54XyMba+oIRe+8g96SIuhW/+HVs0oa3cLfAuAXjX6rdhXA4IY+kzaL/IRT
/iERIE3UWH9mwjD7/W/wI1EjpA6XkNO69+UGHloLRO+wkYaGEPdrJNnoe85A3/n2
5rKzZJQkqzJuawUk8iLIyvyjQQY/B0UFsYRgPZV3J48rj7qkUODMVICRynF2g/th
T3OwUdn2YojSmAYg2NmoZoaWDllcrdRmYMZaIw82lu77HVXaD/x7bhjWGC9ivn1f
VdK5z82meEdBlTEyGjv92s9jPXxTb0ykf43hdTkj9dU2r9tmxWhi6Ed5sjnUml4a
8ivHcMHccD+jGYMa1q71rZBFV9SWxMHvUwH5HoIGhoeqW/BTjAqZB3n0cxmn6hQk
JN2/5PvIuJuP9x06Qx1kNXf1lDJ08s1kv+w4voAxI4i6royA/GVIm/t8hPXrBp7c
BjkvUoJ+inKjH4P5t9FC9Tk0JyMkjy6R5BnX0JYXLx0WZecXWkAScj+kz4T+DKAT
vob272wVMF4aXkkNGEdbAQefhm88ZzipAMsTx6lfvJI=
`protect END_PROTECTED
