`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYTNcbin2hYg+ZkV9COL58jbHlawRMlao6v2kQcj3eolsa4W4eoEuTCzINuu93SD
p7UOATO1j6yk1FxBFYPGWV26LF8U1P1Y6IjGPT4ZvqRSvv+96CGTrpc+vGQI5P0L
7R5I/kgjQbfVSplCbPr4S2mgXCHUvXUFLHL933CnAvAkzkfpKQ0ErKm9sLRo+ZIy
BBbdEyOMLv/fLfwf/go2O+kQnqMR7gD2GegQ0nj2k931VAT/uHNGa/bJ/tJeZZZy
zjUAcz+I0R6lvN5W0AVLZ+LG/jD94BDMJJdcoLlMQ//YoHO8sDAUOcBLruNxzaNc
uhlS2ElcKM6R74hZdcbwUaoLPYUIRBLbMJ0/OlaLdKFxcjIWwFXXkZ/oYliANy5f
c9vw0LFmcIc2ogGoiSIu7eKWLjpRuwDEa9OMitiTW/QGavLTd5r3Yj9WX7P8Q8Eb
qMHBUsX25NE+3n/rOjLT5HrDvpq1W81c5DNzmX62+aS7JV+IC6YQofIw+oWvMeg1
bfNiSfAGPU6unqAv4m0vqIN8tAeuUgEKwf59Bnujz8vvnh2ysJl7L+3il+cZAuTp
+/+rl4oKGYgxyBRTU9Vk7T/Rdyu4UDTo9gZqi6iedzQ380P/eBopqLl1mLKmVRXV
fhAHIsd+bPirmq6+NDr90x2qH0wgReLcspfFCt7j/bfx4Mz1Ct+xTNo5Y5ChEbma
sE6wYOfuiKCplO04ZolNAVzlQjBMBGfhSC9zNf3/S/i6Z+giW95z1PksarNuW3bF
DeGmlV65DsTXuPJKwSIXku//QZP6WxmeuPoc7oJMwXgj8Mwb0dHUxe2FkJS+oeYk
5zFmivVAci0rC/F1H6NXpXBW4d46C8BQECYOcd6BDalm5KadOJhUefGEph83rzVA
g2HfzFuNXx+YnUhneSBkJlj7X3AJzJDhqVLJCNcXUwAa6RTPAFLChpcCuMAEYIWT
rGUOoPcCZY1HouIOMMmSANiETCqXutywwv8fo8Jr+yWtaLMcaEvk3wcklcnLGF8S
6RjyUo6XzFdg8syU3ykFSNChW+d+YjOrCDjUy2Jll1qVG5OZ67C8AsAwkcqqVRPG
TRqqUBRFLwvNaWNjv/A1TgdwQ6wjqS7Z/PjySIjP10DjmYiySw/0bm6TjdEJ9ho0
1t8feT8HzAmHKIx4V6BRVfpPUk+G2CWUH/6rSI6dFW+kHc9TtiyeJORW8QFziCdY
KkYlDpxBQbv5FY+h13WT89Lxqb33aupiRsKSHkiDIhk0d3+NclAorWMTm9+Zcdi7
uYsyRBSSm37ZeXSUjQoW/9aY9fqNoO8fGX/EZ5QhsupjzfKRSBvMCB9NwGKZOyD/
TQae/ZS8qVIoYELhWvWewM+Y1M2xXnGueuPYuKWM1NBxhlb13TWMP/2+9Cj+UT6T
W9ZfA5Hie3zRyqPRqYWMWJMxEhaQg7CWN3vz/EXSV3sdnh7RLW2IF5wyLhTUDIWj
q0sPGfRXcGPxs+phiHq1HZybYVlNzitBMOaZwEh9a3qm+c+eASeXFg9Q3TeJt5bR
tq3XgCPgS8c212D71jS92SnbBjRJHOg8x5INL8luJXz+hJX0q4wMne/DhUUZ29Q0
z2F4MHN4uxzC0FNNgjDDWec7iMidBSAv9mvTxEkyImg2uFQn/WD6vlfkTqasIq2q
y9oN8rHPHhXfvEnqfP+2yEe2qI4Ub4I1jQeQjxkXSv8UKxG/RtPuuOYHVw0POHz3
A7o84sDaBQIeGt1eE7esvmErl7N/J4RrEb7dJOXXX4ZVsmd8S/kW490PqRg0HOm1
9K+ZBHOEyWiMEskoUiSi8aJVJB1Mo9fyUkdxe0ObWfL2X8jGf/QeVIxDcyVjZdd9
ZW4gVCl4DhVqry5BpGXn5QHbD5OWIrRh2wSweOfz9M4y4Z7wADlLWY10Sk4E6l6H
mzsOuCR+3tGQBX20gIxuF8XyFMtu80qjs9/xbfpTonZh2y6HfMGiZWyQAM+ulYW8
AiLfXGkWGLb7RjSxGB7yEBlpCD3hZscCruAWJUuXsa3fK77U2g6RYj3UF2AxdY1I
lDUXx41me1nSAJakD/VlxxBIEWRZXsvahatxWqWuUyOcXp+Vz3SxxXV3qIzOUd2w
SIz0bkzBtjRcRGwwfJ7hcfNlfQGKiFPjgUOTZYJgB3KHiWCiby+dg1cA4iXAVo6s
rBRTlX07fJTfZucwa237YAw3gJlIB1ZjenCmsWKm3G2OV8SDtQuNTczpPypx9bTH
vvbzrdR4fyvjmDIlluCddbTTPXZVziS4BuU/uww4hGD3VCzoUYL9TElJGfDe+sc/
A7aDoenXq14dyxc9bmOSGnzSWzN/sRMGsIRGR0ZTFenbfw9u6+2jBTFym0wK1GU1
cNePfA9Zz2FPh81ptQVVMYr5GnmBM1CP0b/Byc7cH8H8zEPetl2eRWwOS7LCvwXs
fr86Q/xCr/h558xc4h3x0h32PDd0G7OrxXL5Bu0aXDffHJd9qI87H7uCyQxYYFB7
UwCrh4iOYukZ/fu+OSMcQxr6iRhaL0Re9CCONXP0iGqCzj+7v75ACvmlcEVPV0ef
iXmX97SUz8F1p9+F1ECvNzoKFBjhPC5mm8DHBGHXx/vDp4X75EJqYs5xutXfsWam
Nruc8x9iIyEIFIdtg51E9q2okd5X/cYaJcg/ebhYUKRDazHJFH26Vpih9sXaBY36
igJ+MKmo5FFyKPbIqtdndXkq+h5Y9FO8NOAZReKS8AUN3b3r1P+JTBmJJ/g0TgqH
MhplHpaagbookS32FbUKyaKluUr4sRU2OwWu9ALWdUhH814FS6AD1ee8R/jt61zj
uIIRnqNNbXAOXxk/k4xqOxf9NePA3Zz83AOguM+OHVuVuXwSZIdl30DpteKvG3XH
TEQfRGTjjo1p2jkct4qQzEipEMqzCJpVfQHMhayyzOllocaeKGXWqndyi8uSgSjf
/0EbNkrvKTAfYxGRTXLcO0X9fDi1By1x79r6/Et1oFMV6dvoTgfNLw4hWRwjHOfE
8OuCGSZv/V+offiHLs+/78szM+6LkNuhZBHmeNovvwAYsM460WDsTtLCRmnUfG2K
h1xqLhQLhDsqvgV3AQjaNzBAmUegjoJFWoM3mE2TwPHBxgbW8F6ZF16DLE6e6ZCW
9jhliBOxWVFVw+xHaafoRFGa9HFkcHw9OS0FYSdrL2TD4BmedJGbrhtx9NuRDzfO
Ur+5D+PvC+hfaEapP5Aa6kp7JfjwozUrSyRz12aQO1dAt3GeS7ejO1Bs4x6nDAf8
rwW6wjfP3CnlBRaXn1oyhKWKA37gL3x1XmAL19UvBbl/YiafVuuxHFJLYwVp9Bya
SZLUvoDXCCNkFlqplTKtozoVKZ3JPxAoOvvXICHwOUJ+GkSRNZdzV1jD6dXh3F55
UCVjaF6G1Pbtg47TeM/4iSRM6EZ8BQ0Sv9Mr0wfnfwXEW5A1lJmJTOxtMZfPA8H+
Nn/+v2JGWNf0NKh7kVUpgs4wvIRta+zvc9UTSuB1/qav45LlGVOxHZYIu/N849oD
3Myz7cDXDvj/ITxWQBWnasyKpV97MXpaobmWJW55eG0ZyUsVhfMi7eYZEdme2+3c
4D2Uh4SxkPGsawROcQTwNN2SY/e40R+2PKNHoKudieNX98FURyZlwXBREHVYEN/a
1btUI8zL9k/Lbaddhyp/AzexS1NpZfZ0lBPS6mY6Wj6SuCd8tMgAMFPDANfv6PsE
0BkpoKeuPB2Y7kNaRcV+tta67yRj8eyMas4ceEgFrxhcoYRoXWLeEie9zOYcS0ll
wiyjzH6elgJ6IuznLcZhLF0OfPXc/2bkH/4K0VhketKkjXHEiE7X6TCL7L+d9jap
BsX2XAoM+RAuBOULv8JiZX/iss2Ep6KmKZ5JTOdmd3o502/5d7cDrek1ic/e+gZa
YkMq2rr5MQtea10lQ0kzy7ZaCRKBKxOLFOQVjlXB0yyIPLYe7a5vnWTv5y2tRXSR
D6jn+dc/0OlzIQsAwg03EmpBq41DuQmNshA/kTg8sfq7Az60C8naDjrK4NRrecJ/
kpnpWj3cFiRHKJwaPjggW6/NrCWnwxmUGknHB6eO2oLCZxXo8Sf5H2oWgbXndCoW
cqUIlqpWl0mEuXzQMyEi3Ov1YzDyVf5o+16xS5QESsYOlU+6zpX97OezCgYlHV+H
v4rXRWHAcoJfh7nT1joAfmqVUL8L0wyTiJNFjs9xm/e8bvCdDjeoM7mjFHEOmHRZ
LiYXdoC+rzI9/UlXTDOv2NCahHDWSL+tXE7HiL3/T1XT08vJlFANVOCEH+8LDN4R
UiBasL69Chd1T1bzJW6Q3fVhRS/aeTGfpRIgqQoBVqWiMMV7dq6UIEh3ARcMpt3x
OJkHoj3UvDNmdlTN3BWynr6r+cp+KiiJM/ouYScE9OzIFPBPenMt4ZZeIjdOA1ph
KIdyBOuloSDtH9rZ8/Fq1cP+0xPAizO3ajseRiEkbbuKND4AqpyX3T0Tuyg9RbzZ
EWT/zR1h6YJ57+p1CFEyjucTQyB7b1HimuzNgw1wsR/uyJ2AVAgnJYPVEC91lA0e
NGgAqc1Is+iZsxzC0xve6vVFSZoYV5IHaHbP280cEiGkRwRBwlxtClwCMRas4lRg
vj8Q6r/32AkUxKXPYbSuYy2G4kEchWNzC0VPyL5SKISeoJ54TqGTrzAbrHNvC2AC
ludkGBCoivSor+JWpS8pUDPE0ZpxIC6Nnk1saEi3WdbJt28K9av7ehOjf++1GapS
VBOvBrOKd05xh1qhzt3tTC3jEp0xzMRokCmEZYEOif7ssKSGvqRN8ebpwUb0j2Ue
/goWxS1gmvUdR7KAGLoSRJQV5+Ip0JDWkC4nLAoEizaRdFXNJS+jrFe7NElndhrV
fjVs6ox3Cd+SzN7GgzP8yeVYbbA+68NwmRZuBcfauAM6HLHq09mo60OSTlUUTIpv
/nIGYdSVa1kyhIOl6B9x9TlIC1bSJDTWwo1QEf4w+EG9FB+9RaNKChiPVH3HuiMD
83DJtQbRlIUHqcYaM1Eowb5RQ6imoZFRKKSCxqW91uikDyqfo0fpkUBY2U+QUL+W
iqzN9XODTr6CTnerXdSSnzBgAl6tm8z2K8p+7BbJRsmvvJxtH12VqvqmWtEIDUKY
4CYuDkuatnfbA0L0yKHdn6Sptu7Po7xD8Bv+KqQtyW3yvp4+G3AEqb0d+Zuu8cT2
+0cHhyaKRJ+k4o3875D0a5At81HPD+pOt6Af4UHGAK76A3yRVIVDONph5LYgkSTH
mTGYB6wEMHOOV4G1e2naCVVRUVr+mrdNbR/A1uipurXMDRqoTwgnU92w+c8DVPOP
07kezTqMpS/b4bmTkAsQvlYhldrWzo5ZRRPtpv1fsINX2DcgxbimOwB5dblspdq5
1oLl0B8SXJBhYRlzOnCCD0dgyc6Wm5dnkfYk5URn7Gk7GE95Z9mRlRjut2ZDYKGA
f/ZqrHV/Q01paFcF81k849tzFFmxnfdDMYXoD3j4UhC24+BZM/djbZ1I69Ps7Xja
XJNC+brmS2J34smFYsdU72TAhECDYPIaOBp2+WHdN1GQrVF1rpWe6FQrdBN3CEBC
uGhL7SOa7vdcKaaGClAOsjS6n6VNmwbKh7YgN3+jLO87zS8QapPTzTEke1s5Q2tv
yAv303/+Jh1euzabaj+fxRGS8KeVR5RmJlVuj6Q/4TtReKnnQ/4i3QEiY37faboP
dQ0REmRaKGVx5nS8sgrDrTEpL4xvEmAaKjqOgWMFgyx9oizMv8Z5/cB2ONzyAwyS
+BeA4/sTYUsXkamJBrQMny3ui1bUD49zR4dxk6QvPXcGuDx2wud16Hbng/J1wevQ
w7OizXXcCx6v4x9X1x6SbnkrS/puCTg9VefTMA05Sr61IeXWpsUmcIWttZmGmNZ+
LKFNYZnHTSn8N6hgOopj29Y6kSPKfw/9U6M+8UbEpht9a/N4mYjyFWaE3l6UWVRl
ZQ6WEGfvJhrCqDG105SyNm1RylIzK8o8/zRnG/BOERSjnavsqjJn+aFhpx2abPM2
uirUuk0PovVvCEYZ1BnHincxmb5O3SogGSsVopxGsx7/HljaN3covLtdvcdFJOpV
/zfhcErLRGJAkGZm616FyiX/OD2qmGmZcKwCkZ3ds+uw5hyIzQz/dT2yKgsefgsG
PQ0Wm3wH7/mjnNpRDRG6FGfhXiWd7iIqLtl+pNY9gVPrSjC+fuEPT6qyZ6+UCQEu
Jx32i+LRHxAlj0hR96q+N3C+AgMfSZhJqyW4+aZOcKwkZFV4D/vjlKorPiDfw4AO
tj0QsLT7y8YrGyd0704k+2a12JEOgRwG2TXuApkIsHasWoN18a6LxfWkyUYo/HFT
Zg1YrKYfHMysZnoZEcaHD4uPX8fzhKfLEZ1ljb+2WfL+BSuWwYuBpHRaXQ0qa/nv
qCHQfmOL03ZcArNMUo3oJ6DJ4ZPDCzAu6Jnck8Ae99HJhrMbj8pwDN4d+m8Rc7JZ
oK6UQPU9c0l5Kr5Ugj0IiGozebmoaGBNAzO3sJJPxEpvvweIrSkp7vMyK6CcUGW8
C6+On0d6/7a0xOcQP9UZEd9PafpRfusNHnKBPw9lLkEIfQfOOHBEUZstcXmANE2U
bhrFfwazZBfByovg1w88hRNhDvVj3Fb+DvZeabOaazE4x1gADulTayJJj15yRTAp
mVRXA80eE4N+sLvAFp+vXyVUIf7XVHQu676uVdXM62eyPcEUcOylkvr0aHNY2cJO
vFEUlD28Phvs/Q1KLFMC92+nAc1W3COKC0/73sExaCpNdAHj1yieeNL7wXYYmu5E
p8t9cZi97ImRcdIzTFNzD1mpc2PY02KWxy0aeIMbcARSeYdptoDMlHEAtPZkpoFK
DktNsv4wT5NOJMRr1sM1+4dD7CzM9dMLNzkV/U1INZc68sEV/4hLTYY28mECJi67
L24PtIDIRX7b6HSqQwZ5UnB0ANOMjf7fda44o6gh6HNzis69SmNWSJNaMXj2wi5h
/vGic+UWePHRkUQeCTmm7r0TaX66XreL4VetBun9kmfHxF4aya7OMVVTv97AeKen
UliB0f55uLHW9JOV8i+9+IXm14RtRapGeswIWqIXWAXu6VwOUYdAS7Ecu9rWWBMh
zAf+aXpy/AFqnMPkyKaBCIUE1ISz0FCh8o3ZeCBLVPZKNiUaYUNQ8Qyj+UNNcgCq
JBERXR3VE2txmi3imJIeD6j4gZo31dcJpII3bSoopY6c18zE9hRZu9tzGoW+TDcq
CR4d8UAnJhARkoPOV1aX0ulK6iAOgqxm3xAZIOcdG8z24txmUF3elxQKcACESAKU
jpxuWsm1w8ssOfhxBn+Fo8VyJ+7i2K/weyRWGKzPt/yGZMdK+1mxuCxGBLZGImpS
NWuRBlXQVpeMMHBDF++N/w+cK0Q1EG+nJeAwoWy7Y2GGrOFcSyf10hi3SnZKvdIC
Y3PS9FhuUVLGh0pz/QR3Y26fdo0mOeMcnzHQ+LmJsNo4Sk1Ao8a45WUpNPhluAu+
BZxUOGs4uqlT6Gh0NNqDYS5sIYkNg8GSNR73aFRyeYdNNDnEH/dWwnBsaQXBWSwb
01GSaHwGmlbktA6vIyO0pXVcHeBIBvTC1DYM4hKRhbGwDO4DwglVZnXduZwxz7Kr
aC5hitEvGp2mKVU4NiSXyGBNmi1sJUQVxEAbRP9B0NkTJ2RTDzfvYesRKNH/6Lm4
EhbgeirdOTr8zOEE92EctXz9t0R4/wsEBWVSoHqbpUZ0GFvmo5TSShwDOB/smbrm
xUArFapORD9LPQ/R9Vjx/yPRe6u4/ziponXPJlsQ0O66i1qEHqrPzObPSAZZvudY
jzqWYh47yjEwsIne5gBum35Q3i/byRicwDQliYFuovqkkrdhCz6T6NdfgG2MV6Zv
SGUCkzIT2UN6sxV71ojELYTQlLPMDIEtl/2cJuiMZD0RwFkP1/oyJkHU0z1l8BOW
k7AzQROsfqFLmPPhNKNnxB5hcWYxNCzvwX1paJ+X4t0w2hfQjUQ7B8Kh8AZ4DKqm
OU8HS3vty5LzzbD31hCFJwuBSH0EL9ZjaJZwoCcQFQkJU4Sw0PgHT/e9LSIE0qyC
XqatvtbEbFXtnq39TW8oTo47NLMteoBLOE3KAgNX16yLreztJuwHz8wTduvpN2KK
Un/YfT332hrTR6nAVH4PQiImCIfqGcPRARpRUrjMHPk/gI5kdrSDTrcvEb7anr9Z
+wo9kdovxQ1FCgxxPAezSusPfz6/4lnZHsYAIksfnRXxADWAyj0fjuFeE+c1hD47
lz5jvbhm9LylX79x16RwTTiYmM2sKRN7rYxW6cohuFzzWtz+WwfK479HAde4xqeE
2jhYTsqS2SSsYbGbuFa1xjkXOsxmZycI+V0MrpnwS78tr7WD9PKLl9Ydc1qBBhmQ
vaR4OQ0JYU5SUO/RaWifLF8ZHeI/8iwU03Vt42EGHNhNEO3hkK3BM9Y80ggG4M9v
TRypnKfIYytW8KA8lGlO7uT/CTmRue5R269yE5LVrl5oN8VzCtUG/yMt8XyivGXO
iDp+xHquaQSiUaHcdrAVEqLd5kui7e7KsseotELH/yKYgEguBQC2mXjD2xkkw50G
yAHqxFgYy4klbV+NHPM6Rs83VefqcFMybEmCl8GZa3y40hHBu2fP8zpgzzCwTAUm
s2PcBMliAKEnbRtWFnQyU/mCtsCzNTHGEArWzyKY5p/9hmmwxoRj9j3I622r2c+u
hBc8sx16NLmivkV/ecDkkDVjIjhxt6DAIGh9OP46Q4tp6pSkyYT+9uc4gaxBkrtH
wtzvw8oLw7oLrHAiHBpY16iJiT8cDJItf+xIsMU6HJJ9PD4Rd35W0m9qYWZ9JaSo
E0nyiyJnVuKHsPTR0nKHL/Aod3AmbHDsXRp7mLuVnuGcy9cvHqSl98XLGcUjyubn
jl+/ecsuW9OLxNHMUa5NJkEMohR43eZf8enmVqvDt/o0E9auZCQchVmahVEAw7bA
vYZwFcu2VNVpPAKX0+CUiJuPdDxmHTau08utVFtrrPktj/hqTp+XLwS0B7ZUIeTy
V5SjguDWc8euJJ06Ncj2xRIiZT4StuwIylYUntcuYkewhl/Izu4ecoomt/ppNb13
C9gM4ACORi28AvrIrmEkrji5MYHeySpDcW9mJtKuRwPV/tE1vEBnd+VmjlbsGA5x
IuMlqdik8RWLck4r8A1rWUPyWTOb6RjEn/lmjcApn3fpdAAVY3R538zdwBCv3KJ/
WneS8IVEytena44mEWrmuwVA2jL50ZQHXPb87P8kJgAWd3d5AS13UE2ANX3PrXwl
BQZAvvAJV+qEppSYRkejSS5IAdVELQr6aRUu2/xMMS5KaAbfp9RZ8GMIMp/1nOfu
nH5Ay4ZK0Q9L7saLUMVF42cSAVcPx5sXLMl/xynGGmWM5AOlSJseFeWXj+f4d4HM
YLCQYIsegSQLeWIhDF2o/8yCqvkaii5vYlZ+gVueLyFrDbmIqpaBiIB4MZUlnSK1
u5YJKpNvLmgdEKF43X3fPxLAiDZ4WTT2KVJZ/zgIfk/qySdBXmR0r/Ntm9vwcdto
zSp2xdg6sibD+S4+qZzac9dMW5FEPusdDKaqbeFrnm/UaWVLyIdKazveCg2+rVT2
tEPWBQZE0e2pP4OK96uHfZSlm3tk+GX17YYe4Yy7KQkSsp6czZ0qLSCaaYWp0v8u
ePpGC+HoCS3gdbVZl5dma0itjJRXdK+sxcV3amcE8ExBcs0orpplPFdPBFvfylwL
U+HvcffUz1MkgeQHV845w0uNQ/I1xV/6o+lSv4pLlmtTCmwKTAAKz0pU5s/bhIED
FqXdbBRlamBATRHcAEGP0K7glrmosMA7WM11zygCDg9fQhW3dMa8X6bKkheWyMug
j5JFPGmKjG2sVY3YwwZkoVKe+cllMGeFhC1mpnNLVybV6hUQ2dsVrJEZ5TExkFjl
dC3vWGdamjLgf1a3AdFVozLGRu2FCXFby90HPqiNyvUeH7k8DeDsmP0dzyGUk72k
Q2MsXI+mWnvaM1ltlG00ERN2acQRti/GV/Aqftd6Gy6dnpigrRKUaGk0pizSOyw1
eB/8D6nfwyI86RtGyHi0KFkJzhlbXRTXeIzz+4UiQHzm38u9h74VCUSOmdohqy7U
dItKjoeWyvb+9in6Y33wh8jGmDv3qvQsQALX1owrXrZfNB2Uqfj6jcD9NO5cg2m9
hHc/qMB8pp/oHGR38foPnECbsAVxAWMWqheEWuHRuZ/HHLUf4lKxJrzA0DaU07hX
6Rlx89QVjw0dYYHSIPwDqsdQmlPXnVXG8iXEB60zogX4ajvfIWlmqu7FpsF20cXb
21YA8xuigtZqev4RJmLp4Yb3WSgjlmeP1p0h7KPY8eTtoeqxy/ECrGp9WhviOYa7
p47tbXu5YZ+nHIPGhUzbj3msaxvK6JAtHTTHS9c9yAVTsSYNulwP278S1jYJ+7tU
mxFFvpRc9xslYxJsMW0N8oZ0Dv+am2KevQpqWqUvgNma5V8wu9P+XcLyVy0Dii52
m2w84nb9P5iIUVWUx3wF5MkurXgk32L7Oqs9JSeOGXyCDfZVR2B8L6ilRS9BW7Hg
OQmeWPpE1ewUr73y7LchFFoGcQSx4RMmz+fIYO9EFMia+I+inlo5JQYorFv8EJMK
QQSaS2HW2znrrFAv7ZsndLqi1+pHKMNqgOUh3AmCJ9gdggSA+vWSSiZR740hvbjI
GoCYyixWucg7WbCNrTqk8/HFQpVBiDhV1EXWH1pzz+ZO7mAx9Cfhh3UaUgi4hKmU
/8w5PnA6YU44TgOj2ZUDB9jmXGRRW/TNcoJM3HT8lNU/W2/hPX3veMNYlwYYVhlo
2Wo7j2coNj0ktDhQ/cAdGLk11eu6coEzjfknpR7cbZjFpfY1u2oUdvgSPfBqeHES
CVL97cacuQBxil3QAoYtIAgfz9dLSLU8RyJpo7zegqXLl0c+tYylukNIiAEu4yaS
XXUCLex1hIGBEvvyEp4KgVzdv3a8a3jJ6VyjMGeHSsLXNg+qp0lRrhfN778giG8U
24FNaTRbHEN9x5bnLC5cXcGewlwBqZuRCfxdKbVypxvus2cvxnnzC7KNtV42vr7d
zYTruS7hIMeDUwCRaxff8Eu70Rvmin2NM6v04gXO1xPHIqnrYJ1330GR2jNiVOPX
j5YGO6oMidMaP2CHXUCiIHgSl/KYNb2PNHReckEn4QhIGbZed1+YAjYkbvh57DFU
mwDUZRYFs5wOgGvnf1w3/Heoljc72fHZulrAdkH5utSNNLjNGUk9aRuKNbcu7tNJ
OgieODT5lawxl6LjSoxQ3tU60jYRJ11Yupr4iKZY4QOWAO0Y5my5I1OcxGYQ5TI0
U/nD43ULY/rgu24eiZpePgKKa9kHELajoHvS+sXKarZ4AsjN3yfXFZAdGirUDSFI
VDSmPmOFx0cf4zXZIW/3s9VtAf9/FZdv59gtf3J+SQD/0ChxwXN14znh8D3CDjHY
B7R1j+9t4N2oZVBOLJMjWg0z3rUtRHiuMxnhG26UmpRTw1NcXE12rXdz4TNxEsbg
HDDwaNAK8AwhlP2/79hUEW3tkiAOSao0qNFbfUUZBo/KMtBrCB9yDZzyb22lfic2
nlfW+OC6H6Pjo/zoNfqLPOaEwNQYbggZWCZ3ZBlcgt9VFxTEgMaqViBUAlQhsKh6
7SGHkw8Y2MQMuXO06b6b5oIe7SMtDCgmEwAQSMN0QiQucY2oWoHmjUOnseTaf8/8
DP945a8FImpScdqP8Hm9EEwBt4SlF92fk+r/5dYqcTljfiKd3ZOxeZhWwTqWcjPm
qOkwiGbPD6cXMZsV/rXn3UPGDu3NoSh/cdmc8NGvTauv8r+tGpM+sN9eWpe61t1S
4TN7uIg6JxbElEd6SFHqSDLVUOJxcnCepA8f8ArGnGiPLlWDzlZACFgImNkm3uM4
EOfN1tgRHdS3s4gBnWWsw35ePyDjVJsHMP2Pln7oRm1KChQ0C1AVfxg/eIOf3RyH
AsHL+neZ6N93wCdr7LZStMIB+xFodzg6uj/g4qAGGUf4aGbzx9YtiSkhu4DbY9+L
cgk0NTEhjr6628G2Y3rr1TpyZJH58WDlXtiNtOkF0KG8NGKAgABvg/qwvtuxcd+S
Q15Y5h0Jy1ZQVilNeUm/dGfX1N9eBXSuODBCKBXEIgOQmHa7zlf//+uEmj8Wp15R
vvES3HRsiQkTTHX5LRNlHGe8R+g6+sezmWKzWKus92p+IHC09skolLp7Y7jThctk
bNHJXHJ5PhF8ale+Lk9sbfQk2D4uF+OmQ7CmNKQvtdU/Z55waadg6iWrl6QjSSJ8
49y080GL5u5zrmu4d/m4kRHqWw10KwmuXLdqYmdX2H4Jk0+TQe/I9A8yz0Fj2Sn/
N2wu2qpulmUACYuvhLhL3o1FmjpenrlKDTOZMLO3tEjB+0G4hxzMuravuxTXbn6V
tBMUeeJ1GMIHLPHv4lTpjAyb5b2fNNWjVF1TDRcnfNz4iGQyNsmjQZrSp+PbEI59
RfNjwMwqDfA2BmsN58Us3cKcApFAmzc8vrgvs8l2JdKVaQ+fznvQxk+nM2viJzHP
qzKan03uvuS3mdNjmnvm/4SzL8dTsM0+qHIQhKQrH/raLM+FDXX1ZUYJAvyEAmw0
gWF4Tr1+2rOHe27j8tDG4gQHc2RfMpF/y10K16ho7t75roSCRPy3vTA/d26z6uXi
agK7z8IBrh8QpVIRGnfVqZPLB/WPhSamOi6W2NFSjzZzC+AAPDi4vhdvuM7rhhhA
MYQoMFd1NUCBRMZ8m8M551s+9lZoYV7YtwkNnarQiR8hcNnv+zrVGBoiBoq/LzYB
IU4Y86AM3507Ku52e642ZwpXBtJlmOcZa0jGo7o/GOQ9CuFHF30Px7SUJFuC8sFI
qGfK8CrGBNmHSzA64yafg6wgbEGHtoBL3E7zi/u9ZP83auE5wZfQGSRCA/IRYect
HHkTcLS2chGwbJ/nw9aTrFUHE8G5S5g7DUaLMIydui50AIykvNCf9F9hK7l9VkOK
pg1G6svwBjafAN9vtcWjwfJzeWr13dwml3AGZxaniBTUDgHwIuLWU59kivTfw2Fx
9lZwLr2KcTle8cy68aMCEygJiLLnAafEiWXrdcRvR3ah4NLw/sryLAL70C0SsczS
HWkGLh9QHCB7ij+oxXH+9vhOvK0hZphCyH4XxheUfYOua1VbOefmvsf4Xupn0PL3
emtN75cAXNsYDkn52QXVE6xYBCs73pGc5Vnu9hprbdYDc20fYpQFKJPGlz/HDDAO
yciyfEw88h4NoBFjxRcD6n59Jq8xrQpJiIIXXYrRdUKbknsm9gVXnBKI77fyNgGe
WKnsAtyDYEeBaR00VIrNiF6qEC0CVO05EyHZsDjr4YMHVfVlrgEkPO/fkYSfUt97
gcJ2eeSVPf2MsNefN4Nf2ega+GHPoCmr3F9NiwoNi3SY+gLRgLszhMxbqpUCAEwi
JLZtNYXzJ1NeSFckJktyIqrf0J49CXC7tIWEUAkTQDuQIVJ7hjRrZtapEmaedIEC
VcxGSPMNu4lR4Iaz+3OFV3ISo6Y4UIHPUptGj1BoJfrKtZpmctuFxQqeJvEKWfKX
rTD3IVlPAoNFkazmlxXvmk8Mv3JOubluL3pfKaycqXFFP6UG4y9vVaiitQZ7VBF3
FcR6PYlEmXo2fHzWyQuqd5UrPBSfBFu6j8zSdxqn5L7LolGcsf8p6/55NwoTQ0ev
esKa8feVShqs6RM8j/Oq0vnU33bM/Vpakc+bJnr4N2XoJzml0tymqu8eseC0JkDy
/SUEU6BxgWh/3i1JkjX4F2ZbPW6Tgf8X8nXTnEA1ddUbd/4pzGvbqH0tIdX4utRb
iQ0F06etxm/eNsnMoDjGSx2Y4PQ06XnwM64/e+jmCxXJiVdK87CgYpUf9kXeSOYR
CKhPS9PJKzkmKz3n04Jwq2/V9diAK5vMMlll1BDz7WhFbKOuwlvjx6akx9++mChJ
LNdUavDneY5HRNT5D4zVEqpCSXdsM1trpcNW/TV6o7VIwseKqlHm03T+6MM6Y04K
IMws4Hj8ZGNSOtIEYYHbfNSNToYVtz8uOZhV/DvnKfSpc49T63AjadGW2MdKD/0h
OWgM07r5NJXqbbOsLETfaJo15DJCfG+we3SK+zyeuBG/xQ+Z3lIVbHHPNbdi/Ask
J2EPq81PSUJs4P7tPrGRvKkMaU7vp1NuWwPz4CDZCMoVQOF15ZntVsr/9nkGd21g
zsWejF6Cy6VYNhyOruWR2+MnYCorxXI8BH83D0t2GCNw0mkqHdSpCkOzAXVZENVM
kcmMXXWeXFhm1qMrLxYReiLR/PTZy601w+wYwSibnakSdyalJnHu4UnZEntaWxfK
o8jbETfQySP1mcTXO7PIJmmuCvCKwDwZTdMEX0J5KMcUJflZhQ3p+JNGbWFlxtfM
9IYdLVPSObbdKJIM1rtClEQTmI68DEp2MX4ht9vKhiETcxglUrftElLB/kdOWipZ
8OmA5uYt8h2YQ9jCxwEx+Mt1EBgfvg28GsNjYRtP9vhAQqGMmylIvM45UrQzKpxm
16ZKKT8KOZ1T7KjBZyYTPvXNsNM/eibj+JUFTyzg+eh14wtFyoMG0L0WeI29S6lk
hvLYlI28N2aK4wImJ7Y01mmwKSN3mFc0ZToPHBfgTw58ZVYT/0LgDSZK6rszj8zq
2LXhe7Tko6VjJkYyYAXl15J2dREqubXonrZTNJBoDOQ28SFCebBGSlZM2DYVLGvR
HLH+vdB+RRD7hRutTd43wXtXviQpTBXJext4+Y2INV5ABUbYCgWUgHSW5NM8oOki
fKYk5D+gm78l1s9wmMK4s+ZgTue2T2of3pzewDi8mWF2D1sK4uuX+TNnVV8ZwVzl
XBxhg20nvcPUqqfGA7T0D544NYLwiCw6o0I6B/m0hF3pSM0eyl8JTz6Xlh1MtZQ2
GZ970a8LQTg+hZSZcVcpxWZV37kACZeU4C+GEmcRRdJgOfryX0juFsmsjzXGGvCd
MhQ4MozeXALfT3+fQjq8hLsCTVHJnTl09pJagmqOHq2VTL+d5VB1P0s8p6O0alKI
s8kivzVVuY6cvGbbqhpzoJvuNeWfvB3q4XW8m3sLOBhgwp29myjUvx06MkitiWsI
dN/vWn1uB9Jbw+dCGA7+E7+MWFM17Wp3dzBaCcft4JwAimHC4STkpBGPvNaiDWV/
ZWcNErgSTwZu4gNeT4eBYSuqsHEnBo5PFzdKdvDicgmgxCFRSHOfJZpdb/uvYHI6
AN/7Z8BsxBemmAPsjFFPjj3AyIVohzc4SE8XpMRgeMdzkuyOnM+7iJWW9X7DB2bH
CSSCjeE5ljmQ59KBd5ZpAGG63p+9SObwuTnD7JY1U3Yz4ikbpXJztYi0xMp127RF
9jT21FpBxB+NUEBDqmJAHAgsNy7CtwI8Sb9pgbZTNSfFZ2Mj0YHiQFzcC0RvO+F9
OU8Y1Cuvq6VoXz+4/+JkCXkD3mv/k2hLCM/VgyyA52qqC6gYa+MWcjVTBVgY3xwU
9BmdsoTXgRSJx84JeVf93UmuP6Jte6onAVdXGA4fwujs4QDfVJYpzl3RvSYpL79y
+jr6kP4p4KaM2L9iFlU0QpQ0SoLH1Bkd8EN3IiqMSnt9L5Yrw52bwrKJMvbsvDMI
aUj2EGBJ7hDBWw9YgevGpRP0NBFmBsQ62lYbYiIxC6doDPre92p8eZY6gNC3rD+x
sqwNaV5kwmz4avSBlHOeUHXExXovny1zxJjC/Kqz1bcnPYNk7ofdhI6ZbIsQgkWj
7p89JRyn5CCZCdKSfBrzIDTA0hnQku3UYpCU7NRphHqSRTF7+6E8KFiY0pvaufzo
mQiH3ESHVUGzNRPD8DvtZpVcbp0GqEfOOn0A5ydXiNProccVdqB003nKDCnXwRSA
HH5bxiTigbzZAi6wZgC4DdiozjyRLBKJreOLHN7bzk0U8N9CXienjRJUcETQdPsP
Divv3eQgUUgnFWF7yLIOo1eeB9GceygcKKSCFGkKxzHDfMK82FWL22WQVF+4pTMn
PL8uaK0bbwMIwv7Nti9/0Q==
`protect END_PROTECTED
