`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XbT333qz/PPbktgJvUlmVF3Ea2cmwLZ8PsWszk0zk3gJSgdxiPQw7P0SHgkJ4HDt
zbqJZWANY0M712rw0qqLSSs1dqTFz7VqR3Bvfz52SG/eyM4wYVxDhkZpB0B8Y++x
r6DVYJiCT5bNwPi0O8RONDlVHR18luSqojF6GMLEhuOPIWK7qYLhu588+OLcngXG
0kGKuUGXdjFOKac17zGT6HLP9cssmyMJy/APC+P9tpUHwdlFUQBSfoqYKg9EvwHo
7qfZzvI38TJYdNUDBKlUDvkfsjZ8yiaUAK+fur67Li0mCA4Czj5dyJoStmewAZIX
Credy2XG1hqiuhi7XNclQw9ch9L2ZZ4tvPCvqnCYe4fqlf5NmvCa1msrrgSSg/W6
7EpfoSPZ9gdBltSh5+oIRSeYvfbzzueqdPtUh9V0QNOhcgcd/XSaOanCklmGP3y0
79tnCB3badf3tugPN+vx0REgjJI6ewlk63O843IvluyXdno98mKxAAIp/ZmED8vO
JkJ8CT2+FmuToI4dQ/INKQQqml6DhiywnIBfWrTCeFmMUa/H8TujkVmsiSGFPyWM
RYhtTDO8zzOmcPYbIKn699E5kp/v2wtFjzGSA5VfvN5aF45089Fzmb7Hp8TcxTfy
pEhlZ8SGJWzS9xaPJ6AExfmR+13ehp4c7RCOCd5KWL6Y8Amp+K6fk5MDZj8M5uPT
lB/GaT65nP0uOEalr9sJ8D8o/cerwSBhzAKjvJx/xEfWBAO9Xu4w3tWAz2MEzx2K
VpdBr499qyI++DrWb4oTWhZ04ZWLJQBP1FaGTAwy9TXYhxfrdmwL28bI4Psamhfs
z/jXl/1+oX+G6E273MgZuchaRCATacOlvE6gbkBCUX4lnHXc1r7zoZT6jdynkyOv
Z2rgIsy5Erf5k9UJ5j7t7cCcXqTLNvITBbgqpGhamFyrXZ0sljjc+zGJ4BZaWntw
aN6R9nfQI/qvXHVmgxZ73Fj2yVTVUmZopzDw3D5YOGcTSUE/ndi78uf6ToU5FcKO
p892ks78wGqWQo5paSHDN/6Py71Osa1ll50AM1e78c8sRp/BJqb9ej2+CpGOyIoX
vNrJ/Anl3ldKcGxj55/7N1jd3L69AlBLO3rOplEnpztz2i+8WetJWie/zECkZKUg
bReTPutBa5JfUct99xa6mAXNRpLw+/Kn9bWFVRBbdCOAdg1np+vg2+WeP8qNFr1R
x09aCyQg67FD4GFRPtjK3NjacJ/w807TFtef9yRZZr46eKs7Miq6dsIIoiCXUP/M
uT2rl7FWwvKP1ySaU+vFe4BAjGbjgLgVFv/hW4CbCg4ZnUCvwBhB5pBJpkgUYZRG
wzYhsa3kIdqDorYKeXTLDmoLaHByFLFswxTw6azt5Yo0m5i7JjuwtHMdLHg+kUD+
Vwzvx9j7a3q404lia++ryFVE0fZn0QPv0EAnz4N9JDl/deXzUzgmTB3udWWq+5GY
ehp1JAKhOoXTkhS61SdKCCrF9XWa8ize94QQYVeVU70Ji9M1IRMdRoDXi+SZdQeJ
p7MB4R5cyc3NQtzr+ePLdSAUU4XCjF6RN7mzpAVFJjYFr7I3YQJCP9MsRwohqQDf
QWMnMKdwA1uAgBhK/gUxMDVy2tM+VuVSCsCJdLLFABwZ/63jCnK537vfv2HEGTFx
aSncii2QiWuHgZOwsh94PczmrRUBew+fwYa6498MevjRLR2nTJ1EhDhnklQCePme
W7Gtj/BoTnveDwDhRDZWkB059Mb85ZE7OflhKaoM+6Dr1ASwqnd9xOOtjf7sRG3B
GlIhTdeptZnNdYq1RUIwv+5IXpJCmoyAAmalyMrMi46+xKC3R/ZsDv6jvonwuHsI
N3u578iUinjdRf66MxKB4vzCGvC+ZKQoHKS/RXzwTkySQpUxBhri6/iAUiTt/Pgd
FOVGFcj8A41IHluyOxvElA==
`protect END_PROTECTED
