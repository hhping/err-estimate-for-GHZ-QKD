`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EmOxMp0gnzfJ1vEUW4aN/37tDkv39FGPsMoh9QGG2Y3ky1gkpyO5R1zRUOwb2TCB
mrV8Ar/cPOmcMPE29kEUFTbXUiHJOR7OANvuGwlER0uzC4nHMlYprgVnDhKLmj2k
WjUEFlB7REnFkCAItEMH/g0fPbJM1Nr7iyh83F8il2rcLv3fzWkpLPz10HAKGYA2
iN8KVNnucku/QhrhRnsNpr4FnzikFYBbySPRovAridMDy4g64FMgGoy8QpEurwae
pTis+KFBaOoYsO4iXLLIbsyl3EbEBMi1Zehpf+ipcOEq0+e3UPKQ71H0WRk6AyF7
nEzIgjvlV7GRRhb3kRBjZbFkNlbYlyu5wL0RaVqt5GXoglyDFhLKaBxp1DJ9mxnc
QQVVGGxB5Pyg1RtI2E/aEJgkKAVKok6IixpZVdUDSZK0igcUaAOWP4YI6lQiqelh
VB1vsR9dgrvO2RIocaahSiYwyA4c0t0322vdOpLAguLbbli8a7jHdRnPkdNSIOLc
cHl0v45qpnYN0UO1UymB+23dX7A3xnBkQiN1gKBj0RzesYdILVkJD6V+xnXYJDYS
wAYg/3PE8SLsHDQLc+KLqNF2hVSU6CU+bvkpQGT0UFXrBT06SnpG6p3W0iLGaqsJ
rCVdik6nRnpjaRqaumF1weBD92qzl6B3FQNGnngCngOc2Y/Jgr/ilmbOpZY7QT+S
WTAFa4oErKzfwvzOn9YiYMyxjIN1IJldSdH0G/lF+o9SbQ4PeGvQCXCCCPXjgq+1
68LEH4p/cfkkmGl/R1NO1g==
`protect END_PROTECTED
