`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AZCDfmY6gjgYv894g/pwsocGpRX5IuBhIi77Mx2wDdkvSl3YGbmS5oeiYgQ/sm5m
Y+hPI0C2hkE+04ypULV9evXW2pPDXDjlfV2/1+jazI1Ss2cPuBMQKWdqHt9m6agA
pk0nr46CA1Rb/YMngVnJ4bLqUaqgGoub8D9FvzK3UyM2uB4/BYdbj+HYba20A1RE
pxIlmR6wCf4VoQqEupTkcgorND5E7WYgBtr6cjpKfxCAuWgHCIGcm/0r+cKvFeoy
xN4CZxmqJQieFD6joEj+/GFIdVtLNgq5/SkFJjBjIKyXuMGwyPCMJtRHwLTMY9r4
sjwQ9CKmj/Wfnmieqdy0fRBEjRlT255za1X9kB0uGsnWuk1mHsee/gIgM9VS4sHP
NueVZt7kfWixul7RTw1kqoXu6H9H9pOJfXdKy6VswQliyVcRHrTeSWEw4ZyReQX3
9lOFx9wlT65+DkNLetPFXNCS4io5FR+jgah7VF6bQl4wGRMhvJATCkORhgLdQMpA
dDPd8dcavo0DOP3SUnNKARfc8+zD5GN7q5dzP38Sq2QGWh65pCTTP2fzGfkDpQzr
ILfsHg3IBRqZTGqRrCq6lVFyBveHz+ghvyWp0Q+41QmUsa3WQfHwh8gGg/Kb5uuh
WgGqXj1txFgGdHRrOXieecLHgwOGaJhb/x+GHcBUl87kosxEWC9QoSvt5ccic/GC
h2RfMlZpnlYsKiFlVBLeypJkHfSMp5BU+Pp8Ia5Eq8R7Qwon11WJSCx5+F0isicn
KOOfrGkmGBUUFjWA8mQem9XVItzxGGKmElJlaH7RVArfB+SM9R9g8eMerpBXzILy
NVHVKNwTBM/x8WdDH+IDFP0BrI5y9bAoNm0nBVICHpqrF0NNWR3aLkmVGi+dMZy1
ZZdbFOSkOfF8EuKSvkei4FsaFozcN78u/QziXbveiDt33WNUPatvq9wb5K1fdIA5
CfnaZ/yJmcve/6dOoK2rNBUwoR841+2srVaaBivqByfH2KsDUDFjbI89zLjYfKqq
ODKYzP+KCdhTypNC9J8W9cN5cGmWQ59qlVp9uguiFX0eyfvYWBls2TowTxyh+PHk
iHjabsc3VD5/PQgYSG4y/4oe6C+aX5VULTWu4ue7HrEgapCacj4v5Z+fJON5THEG
zcLeotuWbebTA40aX6V5Dujzgy3CXB30jdTWrMwNiUO4WUb8vnBfMxxB2Mluw/rZ
HFws/8j65wDXI+Th7ID5/evtQeB2RA3QJa7bdHvI3VsKxQpRoaI7LC7e0/cMKbMJ
iFHCFkErDWs8kF8zBSFfPd06nnxVYZ5dbmssxEtXhzIuaDLfjeyr7adpjoX1ByWc
/YU41BfQMa7J/Hru9eTHpj/oLR4naos5bYXuSkZZCZ8h5gh/A64TYkGgDeQWpp69
rIuytIEf1aHmYykv1NnvnzUAAsYjkQp3CzMGLUBQfdJFsH7ZTt+90joUC2XJmMbA
R4/nORDzWsg7YsiKqs3+XFx3CvDwXyIHbcR9e2Wphpo4BkaNbqyviO4zd5TRHThA
f5RuxF/dZuDc+y6EgQurgsqxwzC5L4yoRIassBbwPLAz8cVqEop/N51OFKcx7dLk
IqtCcyXeuUfbxulDBjMs+Te6SZrnb3kK38WOUaLlewGsc79h3jMBJ+LIqJXJNMPi
VNa3HiGgB0j1Y4fBfBZv4tYy5CNhyL3Vt8l8Kh1ftHibbwxlBUoUHDII5JRi2LO2
jmTLaVL1I4f0JDlANUuQBdBkM+cIcBnK/AgFnn2sOGh6m89EFvD6WpJzxc2eiAb4
i2Ls9kqRSB1WUQy+iQDBO1Vlr6KI9KKM8JFmz2SZ+pLPrCyElbm1nExfQmJ/doKF
Rt1OVST+g0fJ48c0vSExqtDGnL0oqtp/L8UL2O4DfkFsTc5sISLwQW2CvzA/EzLH
8tdmbmIgx+huDiRqIu6FklqR3v1RQ8+1GkhFSHYo53rT2bJd30obewxcqkjT6brm
aLj3x2j4rHgBlqA36pBOFV+kSDGBx/gx4jYeDNC6J+OWzc3+Fdvmlsd206jRGDG9
VTYKdCaVksFtErB5ueh8cHvKtvXV+qCkgaTLWMHyAIX7qC2M3jre7vdA3ALX2Z0p
l67X+T5ZzwbKaoCEAw/YUNQvpvdnb2/DGy+0F+9M0ilid3kXsSFT5DQmWZXivjQT
G3yD5DH+WubnB43sN9S82mx6x35hJGJuqeuEwqcb7I8G4GGH8ZIJE1t7FtSokYfp
7YClNZLWFTy+eGur4G9cXE2r3dM8io8eap+09YZ5JYzgJn2kQH/qi8dOW5HUp0W1
HNPj+LWiuVyTMjBcMuDw597+OHTHMUFoZDXjS6nvgUlMZzmU0YnIWWeahENtavDV
rsK/T047xcxuxZepP5B4kZ3n6alOmNaCJH1sJ0HzqI+JdLxz4mZLHi/GijRPKJGV
1YXGu3QtMc9is8/kqHui11Ucx3JSFl+A+GWCVZp4+Bgs+xEHeFUT2dWqTsDX0yxR
Zz+1ThIl52pRY6KQZA6xr/DfjnOX5k9sdj5uUyGb5MyQy5Csz0Pu7fhh4N4g5Q3w
A4tWnDdtCKmJNNnUPccHJIENXP9BoNxuYyWW+bXYTHzzSifkoZ8gnTfO4zXh1C8j
`protect END_PROTECTED
