`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lk6piskdUglfccgadaSwb7G162l2v0K2A/0SgGrF0LG+NfpKXCnN2+skyNScCiyO
zAaJ+S30GhHUplmfy9KEQipHfOwGO6sXDcBouVryYHfHL3tt77Ds3XDgnRUM2dbz
LO1JAzqSemmWS44yOX4Fhgd/EZTaSdBbSdgVCtQaCwfQgLRsqTrfjg83c40sAFPj
SfNdHEdGbWae66vVqZqASa64W1Oz1DJgjRG6VKWEwX2pkIcU1IHysz5Kir5u9QKL
ZsKpmUKsNCyoxgqEst6VOR5BiYPy5I+hn54eUVEi2oPV37O0woypFZF3nRlaEq6F
V03b5qUh30xPM2iWuGbezOXSsU82EI5aWL6vXGGVc32U5e55wrtBV1DpJlRQO6N/
uqbngUBpCxpyHyQGd9dF+zbalkYFIdqydtMnLDTeOWOGrfRy6tXQ4U5DANvT5PBd
U5IusPIjLGK6ukwQ9oDiKwPZGZ+1KExpsTjWDlda8nq5H6+58C16LTjHpFf/S4Bc
Xx3hNwSuf5UEtiylXGUVOQAAae7WLMjx43JNr5UACpU0UU0BqFF5E4y1V+vBG2Un
AjDK4WIx/zsuSqe1TC+MzFHsyx3eZM66z4DFJd+tR6ANj24o/OuHJVQ73Yu85aRd
S6/CQBJ1OL3qGpwFiORytYOS1nto6rn9p+GL3p94AZNeTm2IeG8X5bUAR1LJLwsY
Ff0Klwb1CEkr6uzDPXuzq8JvwhnNeGujHI5O/cgxUNs=
`protect END_PROTECTED
