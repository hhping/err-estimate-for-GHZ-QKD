`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INJuh4tLwHkcRCtYCn+d5TNCnMSYZp5n6U5Slxjrw6XwPgWo1RFW0QLECLfpOkml
AYg/Dh9R3+IvL5GT9Aj6i1OgWt6MHgvie4kjnjzWXTcSGHd0FtzK/rCwYIfQTz01
X1fMzsFxJ8djJbOkOrld38J52LtucHdjXTjRqJgeq4vDDhps8y/pGXxU9mAdhRe0
vHzTXMsBsxvlrTmoDZKyx0nLlnSn0Ow2pLGz7ccWyTRy2OTYKcwLEqz2P1mPHD5v
Mfw5+EsKWJ1Ze02qCV2RFnuPDTA/70o90BQ/7g8PLD/VktEKii7gm6ys1k3gnhQu
gDnfg5z2/NC2q+Uw09tVz5nMM82nrEETvpTywKAQLnaj/9jji8YQwHaHkqXHg1xL
EnKP7ppEZmmBGWpuxI8o1ruyWhIVw6q2PXJ2Xv9A46idm6vOIRS22GkLTndrLrFK
gPjDGiuddcS07XoLlrMfXfQre8hrO1056stq56yZp28sbbKBEtGgHdQeBN4LJTwq
z3A7jhUhupMDeSlihttd1QgX73K47JHGabf8BAZswmjeo0BzOv0VHxvKBw9fmwL/
E7Cp3FLHjIFrstXMV7w+C4OwbNSmiEmzSwahViUayiMgXNCEA178rDuFNFmnZVp+
oFmEyVjSn4OuzvzxSdViSSjCDKbG78KKBPvfncOAsfpvP5dxcMqizRpXpc6Ea+sr
zCd8EvBBG9ML61jRPjbF5D7eQT5GZuVA6Jl4AQia8XVwtqMngxvX1QaM/aZ+jK3p
gTp/zauWgajTBFlYZOxCn8CXD/40xYz7w9HbD3QW0Bo4Af9gO4vprawo12XIp3l4
J1MYSy0lZHWwirkB8zBSbxauBWNBtS09fDocuhy7E9l2i97QV117OGKd4y/UmGm/
FGCxt0VY7ABkmpEKZ/MerGHAgqWO33UYTn5kWdyZwHZMkJx5cnNf3VrhfHYhprFi
IksNvV36X0ldlK0k88TcE6h9sztGL2Uq7BHpkhgeFerEltVRNIyVCRma5gK44RGT
sIL7BjqeoAtGrGgtj8x3semsD1AgQhRsPcYA3KUL5ZoErujU45PxYyqNHBOYe/UP
zyMTyeHHQMU5a0ENUTrdspDEV7QIObmb6o5sQpE6EptlCQleM3puLBxt450CeNhj
EJsY1L5dhLKevol7mYkT5YwB6cXTsCRoI6fqPrp2cahjXTpoy9zOT0JUr0lD86eu
zVWjea0+4qwWdhNRZHUIswFh+FklDRxaCc3rOE3Z0P1EqRpAtwXu27N4otL9KWhM
+pDSyMichi4Brm3LtAIfWtNEs32tI6+DWBIoQGwJLQqGfK0RD3UJskugPibTUXn7
k3o8Ab3VybY5RJfXFc9DqBrd+IrWlfQBWWAHIgJNS9vpG+96q/sIHgSqE9LtwiPM
DDD2O0vxgrEsxdaqdmHCzKaf6Pl+yk6F7W5q9ggcFcAef7d/alH8LnKblRQN9aPD
04/YhLz00875TaF7Hs2igsq8znk54hKXSoYFlbx7uN3YiaYGRLNvvfbWcCZHoN+B
58VL0YcRoj8p9MT8iUZcQEz+zrTsf3rUNU4tXD9G1mBfyVOnKHThpJhTqsL3DJJG
ymAvqaH73+smpUE7Up0gZ5wANHnFog2L8JdkW8Gpca1VoY5a63yirngDR2hlM1vq
FJ1ugw3Yc2cI8JILopvTpGXneUdUBAFVa0aXTIvoPl21g5a3lytVFn8FsSkNyvhD
fMK10c2Fw8pqEe8VD+Bxu44yZWyYoQW494ovZom45ys7RCwKt8kO/fI1bTM89J0u
otnQWbKXdfWcg7cIhgCf4opOOS0jeDIaAgdEqsv6oxnzXWRtlCJqTSH92VYhrLEZ
Wnvlr4CNYi9UGHnrVjBBmhN+8K8izK4Zc5HpX9LWLjvl0tDVHcpiihQc/SSmHh+z
4wCgSV5Orp3aIV7MoIzBI3/mofFCMbHNrYa6bK2V59C8HOjZeLLn7jJ+LWwlPtji
h7kUAXsTvjRsquLXjHAIMS6jm6r3BIFDYJ0lbE6aldhztcO3guOS0y2B1B3kQOPt
OHJrK5EXqHwfBj0I9VhCmGQ0PzQWN2YbY3qMK9inzj5bzTh8an1T1D7uHD/vWgvO
lMkQbYpdgyt7eD3Lv8s7AENBJPsSbwK05h7NNSJPSzJw/Ax2AdFtc7dx1oiXvVpy
EhlHIN5Bq1YhkC49MRVxPL5V2olwcWZ9fsulpmhxdj4YmIqMeTVPs724q1xtxvnX
4DVoObNrYJSjF2M5SylrgI8LuEU0cTzIpsChPAupETgEOtOktmcEorP0GkKhrMju
TGeVZey10gh0Wo917nc5ByQroWTjQ12njeU9yJMQNjLnsLW2w8wdZVi8Szflr2Tk
9kVCRrFysij/TM8PSo0anCVFpFVaPJC1rK1KqE/UU85YqKzO1Z+PUsbt28oWE8r1
NNPJHR3lsRRaBC044oeCB3MiPGvYC+sgDFTu2X7B4D57DlvVgKFbCd09Y4KTgg8D
g88h2YRdHwaMtYbO5rggfqe+WGPa2ygGDQn/2HhueqTOulqce3gbxvmrAxIqJlNr
G2TGv/w+SwmGjDzrPuDNtVoRyUq1XGAGCY+PFXSKlZ4X0d2JfKkS2CdEgmraMjvm
w71p6ivdp1yi3cyOdP4RinccHJE5lHT3eZ7zur7ZfGckGvdMXYKTYCX8KKHEkjk0
kVJr7FKVgHwsbLLOx+7+YmTUno0b7kqXTGWgkpcx1382zIqVSBS1AjZmDCSn2BOu
wfKSCdeID2nG+SMtdSAGlY9C21jpXORHTBCAQr2LmbOF/ITU/Gl3OOhyBDk0+d1S
ajlGPGXxIfr/RGb95B6IN5c+8+LOYV8AK0iclh7v3Di9QMFrA+wXYA2UKbv/s6QV
+sWLbmWXzhHEhTIaR2lNNQHuC7thj/YG3G/HkAyaEnM3VGXs4fSzr/tKAZQdrswz
zuFQXYteHBOaJ0wgrwua9aP5ugdLmnaVAwM7wAw6Y0wtCnQDm7Ccrs0J8nvht0n6
sJbAjRR7KoJpdnfhnDdP3S2CrBz+F4aHujbkjE5q8xOPoE7qyhy5gKabAFAAi9B/
ic9yvWSySqeChLsWbUUb7OQJN8eqAk1q2M6w9S91j+IdhO2TN8gNOMctPAfcO60E
H8fwVfWTJjgE8ueZ1NSgaJx/Sn9bqiAjw0Y5jzcJI0qtYAZRCFZ2R3KbAY8F9jjr
pVtXewWLK6zt+RGMcqmjdY4WAfh6cPnUkfzb0RQMTFlXoeikueX7ZbLn4K27plxB
nQfrJTg2Hb/m2nZdFBwjf7LdBuUm81cAheuo0U3P8yZveppJA4GJftzDslwwh/wE
xn1+7dLJSrrki9MgDH2rF7cLUDn7f5YJsiCu0JDdyGSYcpB23Qkjd2Iknit3H80L
nU8aWa3Pl4UyOYDm74B2hFxs5gAoDEXKd9MO6eE2W3QP3IwyuP3C1EgHJ7uOo/1D
yTyE2LXn25A0HXrN6EuGoZ2PT9kVF91bNMJv8Jb+XOQjk0duR1g+G+2X1ZtV/V2I
DPamLTtnM2F5189Pm4NfTcHrT+kqXvMp40a3smMBIVVQIaxZeIylVTHVKLemGFt5
x1uYkBdklpC66UpJbsDZwg0hXshioW8BXWMfK3KX9nlDH3N7A9+gFErX6i7KDSvX
gRk2UtJZKLcQMtJLbqEASyXRaW5jV83uYx99FNWLGh0JlrTeMi7jEb6dZqnF6HMb
DqxyIBwOGa6eY8hK0Ipvm9pMe0kKEs10m7bCj2USVqFPwVdEfHhUqy8dRfwMbhig
UfNMXT3fwa9u+gvzseX1zlgGkiDZ61F1sKunGs0f185bgpEEVx1WyTDwgic+3QIl
A4PnmPSYiCMrbBZWWaIkblwk8zz4b7vP6yR/s+hhICWQnx5pe00ZsOBTYj6ruM/I
dO2D8kR8f0xQwcnEeI6OxQ7ZlprgveSul8vvDC29aeAtM6Z8ed7b91zqcG7rFAP0
kK2RHyWDGTCA/XUwWgTJNpr8kS8t3vbI70lJIpuaGztSbaDOhCqv1HB0zgOsNg8G
G1kmSPI5Ql0skPB8D8NmqVJRs2cxZJWNhEZ9W9jiNN6WCqlkj4y35goxuJwjvpwX
P5os+iCXRAEn2JtYhHy1pshKAP7v+wzRK40q1MuWca/5IfBmiOfpgp984pCPEUNW
rmmnoprm5QJFyRbZKOszj+yXhe0HVp+yhFGdYG5l4jEW7R+uamovtJY4YNgbvDff
5IYLPIQYGMEiSCnRNQDFhxgiZiISnT7qOR5IWZil5lFqhorWwgFCJ+OGL41kZlFN
tg0Jh1t9Rm9JBy95f62zppFWO2QcRasDmdlrAC2FkKl91I+0U1ADCSR/+Af4Hi1i
XbCtvn2d+DxxBJvlpAzlquj2s3y8Jmd3zjlzrys4LT/93XfinaZfl/DggnLNKo0H
KIQYPh3A3DWtVvMs9Bpc4RzbXufnyjxcnUNc1Dm58WbbM7IsXTlEHIFI+NFbchRh
`protect END_PROTECTED
