`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wHiMKELMO7NowcIhcI6DiYczdUKZxaV6XINJsffKycG7iEwCwN6dHzhkjGlgwql3
5w7H2haumsgEvWrhd8bt4qcDUa77qDvcMUgFyhCuJq95T3podDe7fLDFV6SkmmfM
UM1HyrWJdVmoMjfM0JNutIHGj5ZWtwNjCVwOt7jPJCkyFLXOtiE3njkCBaYRnUL/
gI1Ae1JespkZ2iehVmY8NE0qngFaz84OHbVAUlqszHsNVSEP+w1epZuaKpq2FLdG
wzHZDpk4FOZK1u73iiUKV+nYCNu8SVSwIYkrnZ7RVZYiGA6ngmnkie7+OB/RkMIm
ehUEzhus3YTo41Ky+H+T/4QZwe3lme9cP0h4uFRmHCKgPEzul/fllh+CXWFTq1wE
xGL5k23nVWKXrYkwwllpBGyGwcAGX0k/JBVm0inCjcQOkimZ4g5/Ryujm5kqzwVc
dS10mUnx2V7vn1CCMrvA8QKzUI+BvJgBr5w+6A+qe1yo+nquwNtBT1sQ/1iMpsKG
`protect END_PROTECTED
