`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lGKwm2G1EBIovFEyVWp+oP3hbQxnAJPdnlf5Cm0fMw87c/Lo0S9aSbqMsxhEsG9
t2W+AqcJbHcFpgLxIFItd+2LyLI8PjpXn2PbSaa3j5/WE91r70Oovx80CUcvO+MQ
5kmfbp59yQHIKLiDjZBDFStusEKCbH8UsxS7v1v1rlIMI+IHhX6Kwk4EFDjE6APc
pawtfbJvqVKzS2tTiFS+z746iLWcIbgn/YWkeYIQNWCNzRDfEetyApN4SdTUwHCi
SBwPQal9NwkazFmVEXjA66xin9w4NUTfnfpTNOk2VILS4ZGnibqPku9aB3uHTA/8
hd2bPogdPY8ZXWgTRLstbP74Q8nUXtOxTGaI5xUci1SJSAoctfsSwc5Yy6LzyfXR
Q9AYC/r05+/f0+rNnp4dp0tsxidrvsWB1ppEe+8ihp29EoT6GrSi7u9oi6DnxKts
sKt0bAAclHKn94Vfr3Z/kT/pYZ0fkJgGcMeRripDPActFzPiFafTG8H4UG+EV8GM
bxUg/KABZL/Vfvzj0qeXBxWTCYv2G0XzlVf1Ol0HnKyA2TDOdKIF6ZXUDeLm7bCY
LJPDDA95IU1afwtX93liaM+mqntaR0DCu6L/MfsLMuvfu89eAHRsiuScQKO+XEfV
8L79hlUixHZsgEohA91PKPLOZf9Bik7lw2WDwiQ223En+cklJzvmXEySgZarErFV
1JxDKsHNYHz/htbopGZ6/gA5AXxV6A4TwqmMh8R+qEHNBJcLT1jroKvHgxtfacfV
IEa4hyT/QAxPazU5pH6gBfypEDk7NFDVLNGfmk75Ufrub9rqfVpD0adhKjmd8xQW
QDVFOacgg4mqLa5aaP75RvolpbYOOrRX1eL13wEuvqhSagwzqpajD7iCqNug1zU3
DxWJRnCWKNVoouTnwLjMb1e6X0cUp/dlR9cSgr5XwMppmwGfFFR1zKqMihMo22IU
PLQEGLssqI9StYFiHTNFZGnMlflxN8nsCwAvkFZUvKTI1PPjEpqePzfZ5CdxanJ3
TwxqTTI8QlTz4kuFluHW/2xhE7pyPgRud5QaMvMR4qjSEYwb4o0IkyohFyeZfkZA
35DFxqz/PwgErUZatElylkYyCDCQMUFLqLKYe8w7q8aULJNskJRa/kQ8zDPvtKrP
LM5E3slocugzr7gHhu40RV4kcnYwD15oRcH2u+vZ9TJd2qfiJi/XXtkhoqy7/uS4
BxTFyo7qT6CLyaZ9A8u7pBTOeSPEJVQFnM0ZQhbMrRZA+w1NlpkURtQp2XaZfSXM
remYiQRNIQ90ELGGXwsf9tMODGQ1xvLyiN7yTDuVQTBGmzl7B/+4mybvyaovzSrR
dMs0a5SdaLeMuEmqY3EMZGxct46iA2ZxGIFEl0spfgKqPz2QNFpTXb1EavnVPegF
p1zXFmJhnfL2iDVBTSPzaEka7f/gDOYjmIs/fo4xnvHLXU01Ui5tPqOgAA6lYvfz
cS/k5adXK7vaudf0Fn2Ww71LPOs025D95BXVF3poYOPt3chbVD457TrN+Z7eALsl
tBqy+rXt30MZNRguxU5GibpTiTyTC0xcHFp9Vcs/s6sZ52bBffcmWC5KZE7qrGws
zRH2Bn2QhHPWJ1LrrS2lpHTSzwmWJlfazkdb9M+kCsmSHWZGQA/PyYIoWTP5mfMt
kBWqVFaZRaHzO+WgbDFNUwzjlZfdjS3My7xZ9pgRb3QG9MxKS2jxRtwzgTbUQTch
`protect END_PROTECTED
