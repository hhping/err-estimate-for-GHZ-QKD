`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSFMLQV67795rQV3e0NDTRue0lkZ0yNqEvUn5ErM9ixPW+v8LBx8QDgBJTldJXJf
K3e9jpKDHJ4vARONnNhFh79N5JO9lK87cNEAnJU5/0CLLuqRp6HYpxPoYxm7mIcK
tdgOqbX+TZWkNgLE+zEnLwgoajIij7YkNGIKMGKUv+PXTmy9I+ykpzjVgylHk85Y
v2s7UVwh9KXZtBxw2vZLY4Em0hT5rcf5qy/ofDQ/Wy8rhfiaSrk58VwQXhgU2/un
kK9n1/MCxWTGL39p+nO9Wc0lFAl3LnIskLAWP8u0X0gMw7jRZTvh0JIyJMi39oDE
JcpJReGHCnYXZFzoW/XS83VrtrNZvwBFZgUUSI0sXwmV2vetOeG6EaeFLBnmfO19
RqBf2bt8XSPQZghkEg3Z12K2MFbudjUoGHn2clQB41wqXH+TUfr2YJfKbuz/ZP0T
RqngSyBwz8cWpSLkBt6fd6KMKnF6dEIxUWEcULwZSOzzJrLI9n70uuGGvriltIZN
oEaCqvxuxCSm5fKO9S4dW3kfya57L20vVlxWQmjdrWm7YqnCLTPMMCHXyKhfWyc6
UFxSe/0dkNuabPaXuduuS4r5E+eBuJ40izb9QNvFz8y6ykW6t25j5t8lk2XgJ3AF
1/BvNxoH5YNhSLQ12ys14zR3H+2hxqUPsXvjJUdzF+UsnW7h1/FwQUsHWPkCd7qZ
QKPS6+kS0XjnoJmn1hplK8ci3z/wXLEpPwj7y9vK4pwK0OL6fviauDmG+OnHEUfu
spf8tDtOl3aXSAwG6vzs703qqCQlq0U9P+WZF55xJQv9zOznHlrabXhrIuPsyT1o
eco6hLK3ubNU8k7ylJchhAEDir89Vt1blvZoz5OxMpApPF7yCHFj3JbVNpe63oHg
4WHbG1u8mL9/yNITU4v+ziYUbJuZYymkYKn3wezIr7C79T19YVkQyxxjF7HwQBgz
HPNKxlzI3sJGsU5hEWl93k3roSEKCNSwENzgAXzGHS/Syrnvqsay6jHcaAvr8Jrn
653TgNEQ1rWYXrQlgUzUGM6QKvh/6Y0EzhjcrQMceDc=
`protect END_PROTECTED
