`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B5TciHeDmEqClvPBl3LhwLz7Fev2tpnZVcgQYxVlOrQHwgnzxBQOQilKEY/oRGl/
+JDfiMVlwas2hwW1fl/Xk7R14vlAscbtHjV5MZTCOUAzxLly6EkqoiNlpptJi1Lt
i3eZTXnZyvFn6ppM8fwHyBpBAW4Ga43IjP+q0B3r6/vTkV00ZFJCWquJxJMuhHxL
Cwv1VgIyPFyIn/p0gHteA0fbdrD6piezaqGpX9SaJf5gV/mmIrL+xiV4TtAQ747j
s3YWzKAVf+bu1T7RKAfO7TL4WJsuMTl10qIkbIm2JIJbbQR8H+Iu1HexwB5SsyAa
zJS3G3p7y6knEK02lEtCgVZ9f5CCX3agpPqGRgJPKo27DWkjENc8UMVJ9G6LwOtY
ygiELKVIG+yROaJ9PI5S6FeeHLWamNdoMiBNs8XGVLheReV/p4WqnW6+0K5FwX5F
n5eU/sy/YDhnbwgCgyL8FO4YJdFLTv/F0o/3DBViF5jHzk0IzoPBz8hkEHAY419S
IZjsZy/NlLhNRj8h/6nNqIbsJ0Cw0giNFFiPIr4zFCnZxDSJn5bn1Q5VTUDXQMsG
CcXLfPUH21uXYgpQukzwcAfvRB1jtgW31yXvh5BgFI2Q1t0As0UgBM3JnoSFj/kP
Zaoq5ki/NnMD+GW9EOGfuxTdHN8ZHBMeCl2ZeeOD6j3zt8vESgFd6kxsZ6RSjzwd
+18aMZSoHodiXawMzcsRMP5vYo60TsEVTBCoOrvCgjteX8y56Mn2OFbB5WpBaiK3
W3lKuhFCDCXVm/8u0CC+nS5Z0xi7rOe+yzmoKMD4nan1hco0kgEUt0al0doqjtJl
gYjReWkA15pWFrFyooggQ2UmDi363BGzk+wJa69Asuhm+o7RWz0fmbT8+PA2id8L
mMBOH5mDj92ExOcrxSVrarUeAq/bfiCSE2lisQ69zTXtBzzQxo564TYHfrWKUN3X
fuXW0EBcXDPLBzPqdfdwQbpKDfIsmizBEl4VcQHuI8vws/xcB4FLdfhiV/gt4yuO
fqAGlzFl5DriI4yMXOodRC02+F/NhKU7Ozm7ZdalhO6kEgi5jVuAeEfiJ356a9G9
yvevINbHqN82Q7J2YAEAWMbvFiPF7Pcp7cl1OkgQOwQTU5IiNLATbuxBij+YtQoh
mK2ENxIwLwe5V1xtRxcslQOC1ZpmlGBEesm0RASBKbqN6ApVlwHfH6RqnMM3L21V
fI5QYHEhVAHdz1yQOUQzUZJHxdKIGZkQUgleIDJwxzUttnv/J83YW3BAdbWUA6Bw
exjiK6zLPWLOCyuwAg5+0aIKgvzyI/bPD606wQW3KT7EHkxHbbMJ+fau6qZOLijY
e4TJfvaNshZFoR5fFLBn3wFZvuuWz3h98EEeH73wlieEwL/XG5+IsfYsaclz7mpt
avjePfODUN98W6GJRrqQ0IkAk53G5Q7zH+WjvrgB4sJwZXt/Tdl9gq4orEzItAQl
uJ42M0bKj8cnlqRs5GuZdfHJVVDXVOgGRr6kNhmyaPxUQUz5OVxjKqY35Iqp8fdU
k9c+3zkRUAdUfKQpTVeq+0pppYZg6YFaQ1+4QupevpJwxDhcAI27gjMLUiuIZfjS
xOv74B57QM1CfQUYc7+GbW3bmB3qdMh7mzzrvM8trXXE5dW5K+afSEeNlfXcpyul
dmk7h9c8g9cet19TqDFFR1yyjcif6GJXw1srESAo+ErMlo1FZ7Ea843Ot8NSnBTw
+tz3oXTYOBowed7kzk/VHQa7WJCgSjSH5HsUE5z9b93Xg6HNHssLLyzKQqKlrHaI
Fm7L4iNv8bWuOstd5txbhqPDrUGBlqQbdN5aRUiAcOJjKga6aq6ZtxByuOnPTVKt
QcrhmQ0dII1+/P/lnjfwlNqu67ZSiEo1cb303kgH2x2lcSKxv5pkZ23wMOQgvD5T
wHIknbHPOhRARjhwWPiT68xmM12muM6afauIjMw28Js5xQxHgO6nfCUwIXwWDZFG
`protect END_PROTECTED
