`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnb7iu7yO3JkiW0dmtFV52dcps0jyi5IeGqNwptqAzHp7Sb2Mi2BnMug6gUsGLHR
+kcpjD+W4bIASwJu1kDP8L8zbC8mMwxJcivZIp49wSdWCJHCyXhpklHML1tXvEsy
d/UeB2n5crFFDq4cvRXTJMBiK3+CZ/xSGz0fYL5xilgu0lYd2KMNi3k6+NXPvL8j
dHi7G63kq7m9KetWhy228MSk74CZX7vNONgQyMCCUydVG28KMSSWn/bZBPxnjzhE
S+8Bs/L00ZUZPllwFxvl72rBhAeKWR7fR7ZrLlfc+UBRwa2A5fClHEdQrfE6Dtvi
o22W+zwczZSQAlH+vMK54dmKI4oPSqa2K8yX0GXjrKRTqh7FLo/QAmxQCtczjwlo
RC1nrOvKFasiig7Ot94DE98qToOSRjkmBtVki8m3vIe0dUkzoeXeW/nsNo9CXtM7
N+tQzypOzo5foN1R6tPltQfcaf/6vM04OvIxFs1urALIF5+HwvdC9beghIQaL2K7
ZgscoOFXTFJc4RmiTc+LnFSnd++BCzYAp0X8fKryhan9tzJfBRNEi8ACsHbXYMzd
21ed9kn2lC2Eb5ZDrRG3VQK+H6qMS62EHFrwrZwRAaIbX5pufQO7BC6oG8slnSKk
RLbGBv3PbaIKDM5O20Kc5g==
`protect END_PROTECTED
