`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzQB9zcbsmx46OpIWdgrzJ65UIaDVd3dJ4RoZfVHZ49MSmIOBtweYaI6IKx+w5t7
kTLP+ndxIsn5XcS/qsS+ydFoXaC11kkEvlnes3ZXSYWmOVrN5kyOep5yWDf+RFlg
4ZLqOXVYKrSZb68RBEfwwLR2q/5zYhGxVRNVPKAB56RQ9rCWmzqGh0InqAjJhAaI
0UMbVibzFd0/jMNcBxJY4wITCPN0ydpbQ7nJxYqK2fB1jlEGBTkZEMN9s/VVvLiS
GFP/5X5dsGiXF/ZIzf3/UpKvaWTyC3BLKDR34CmdVpcLdUV+NHKZY33e0T3HN0T8
yc2AtV64UkTMQw0QTtt+AiPJ8voo+LzKtZ4fDDlWx77deN0s07MUUnh91FbI6T96
RsLy2QoTrhU2ggJiosuZ4YDi5q+Xyv2HfqAabXN2QJdDqQsDGcWtTcENffgjfRvh
Gmk6kGfpZOLKYwxXaobrWO3LtSfhMx+xhYLgGdr607B3LIEAJr+9WePn9DiIZ7uZ
pj+PcZkl8izfZ8NGljoiWE0CITV8FESqVmh74ql6aPDMg+5Nk54jcyE2j7w3sifk
J5TH8QcpGpL7CnwxELyUIdRtpS0SCc443dXniQnMKoTj4pZBWbe5zEX03fP3heE9
0JvbnrquAzYxMsD27z4TszCoPVbAkJcZYNDtY51fq9xUvReYZlYe1N4L2Uex5piZ
IUql3R43MR/to0YTIWMAyfYTCcyCC902j9wN0uXglTtprh6OlTdttDV+KWKVmWt6
FcfJqSN+KDB5+7mtnUVmB6GTAxU12VstY9jqYI4P12gnt2wNqixsRPtG6flj9L5K
Wtvu93Ynr30OCmyYbhjCOGafgVajlYT/V1CECsFLWlUNkdPCG3Uqj26y2CSCgzZ7
GqW7JD/LpZu+P+kkosuyRGEIzr601a+nJK/FsFd++aniutIA4sLcCi3wBoX7C2ZR
mgGRXQulp+f16mLdEaAvgRthA2VCuuyKjgnYmQ9f4jQ+jnlQeNaC+kk4pSBaEsxJ
F7zeruu0Qd4OTe5KK8bUJU3/Ivg71mFiOujBpJaADybu/lefxb6z7BSKhxDHkQWp
3p9iedMwPwwNTXO2t2fJyFza81Ih2OPSU4ji0FBL/0UfF3uGOI30gfcEf4GbNtRy
S4UPc70rDwe8xTU9CFC7u9rRVbBoVMsMLTeFbhrTn7czdBNk038O2PM+at9J3OXS
nU9PtYdC2fO1Cx3svFRp28WFaE3Kgk4Co/nauXTRyhwLKr2ahvKnIyyVUgVK6JDa
QjbnqtIYXBL9ybnZ9oW9vHTCfx5tFKgvT6Zv6k7eN+GrGFo/K3k1xU4+dfGvmRaq
ztYhO0+cSdUmA0rD0BTTezKCJUqvDQfrEvf0YfL1dkycFBcW3pBCkpifeVflJJoj
vd/qXZJ4NwLm4SLSxQOKJ8v9yRifXIfoGKD1/G/rm1TA7dmq69+VRjYSQqK68+nZ
+zgpn2BcMzzstPhZgIr+48n4qNSaddvY0Mt5iFpa5t0lIjvwlPebDV9YYM1vPRz8
b6WijvXznGbeBEIExTUfsoTVmYPomLOX7zCi2jDqdWNHMNk7MtmSr+KA1/U6Mu43
bZtf+AqUxR5YfvETgBlnfrKvSwKw06REuwX1oQFAdeE4+WOO3qjETlWmql2jdsqC
4aFqS2zm5YI5mBwatc6nIJVvG+tqqTHWfwnKKZR+jM+kcOwrFYc4p+B3Tj4XqKGj
J6QgWMIMEN5UM2OiM7/Rug/1tSIn37UC5dtCOTXEsCdMwveQ3289fuyplJ4rLhwc
vGdtP94cdJEyeZfxawmM1ALTszvw/nEDpeaivf0NASpFaW7+MU3Qhy0Vt5+Vxq3B
PJWGKQ3gIHyme/R+zDAAAW56uAizkfXEyAXRfOBxcNsa4ExJ3ZPH0JAo/XWMEjiH
Qw5tZBlFwVGaua4ZnpWM9pLZqdnzs+X+UjzL0KygtdK9N+0AnvLWjii1ndaz8/MJ
t5/hMrFa7Zm7VTGCByaqeZubIWBBt1PtEvz+h8OID1YyNbEgxJRkuZ9SCpzor0CA
`protect END_PROTECTED
