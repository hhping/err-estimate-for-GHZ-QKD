`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kB2+JJ7DTgF1s9yAktDq9zRGJTJe6jDhjlMp8+y2FDjDUhkoNfGmO1SWYHdB1+xN
UG28JtMYWNAMWTfaa4t3H94BDeSjHTuidyyaxo8gDpihMaLncX3PDzTDrvDG6a7n
Cp7ieUKMAnIjadZ7DfgfOAwIAPbNaUTHVqTf6jtKPi+KG4/jHa7kZFCBx1GyAHm8
ETbDPY6oFINqsTWqsSN0CobvdK6H+0sNiVk8rhcQewPjCh4Xx3pmkiC1CczcJHic
UfmVyuAf6wIsVDPfzo3Dg/g8vs96FvZfH/jCaKlSo7z66LDEyLUh0S4UpGFmORaz
Zv8VXH/FdsN2zRFEAElcDfi10sPDhiotZ8CoM3tlisqRqcvrgMLi9swMn8zCxVwR
KObW6iFUrjrX29IaoOE63E5MMsEP50ePgpYeiorPwKCZ1BsjpBpKF3D5WVronEOP
2ZLXGuGMaxntBqAAD83HBjRyp1K9qAlCDKkoO1NlQdQY1gST3AoFgf2x9MbuPPwW
rb3MRN/E4FzGX4rprUDWKqCL9qnU4jDux69XUaWmiGeYKp/6VTOTk/KCL89xKzAN
Q/rwZB1Hcypghu6l9SGJJ9JlUOEuTHIVvLzJbIlG+lve6rHYk0V614xBo0OnlwO0
zX1ZxvrwXKhYfw42872tzVN0/7gvXOLFhjl9xJv/IlTNywssAlHD4z/HqYx6KGhN
ST3N4NdX0diWM6JUISj8SxJQFPC52IlaeUJ4La8y52FuZMNROWCx/1MpJH4gDZIb
zMp1Lo96ww0j+PeiqL532ckRME2gx2L0VukH5FwAdZHeavv0kQT7BxAw5/Qmye35
mLHIni0w877ZNsyRazAyTBTfyy3bBLQJubVqSiDjD3pTkXJBdEAEN/mctnZNx5/u
kAOLUlHWOgqbg8E2ANzt5jfs199a2dsvRxh751HF8sbqZqX/ktF08W+z3Ao8+rKp
nHNOQoU9HHqeolkkaRMGJefO6IxndNPmHG3rf8/Yji2roeDdYw2znVny5i5EqYo/
zM+NBKxyCqgTB7t0vOepI1fxgFLWNUJMjSBAAH7jbz8o6UMx3p0hhntLGG0hPGSA
gp1eFvD9YNjrR2U91x+jZFeVJ5FByEXdm5sS5P6DF/SlmMUN7C0Kf22P67CjMTi3
CqKDI0ipcC99GMbR9xCM8KPucq+koStptNLYWE0juk2JhRu7bG28mOHtF+sqotfX
QxbuAWarfZTTWh+k1p02DN2aEJw+7txA8xmsEzXhPFtVUg5eeCnNuZi8I1YGG9MX
JEhkZXSDFil1fAghNuZqde1jxh/DCgYVUukaUj5kWGXl3zq4A0S7QyFH6ww6hu3I
JzitG3EZD7zCIYa48ZXK/A+4+Vnvxr/vpEEyws2OJXu12H1DI37cwLp7Qx+iKvl5
idRvd9NFiaBllL8ckhpZycvKUZNy87LtzmtArZbgCDi2A0cDxbZ2VyKtvqpM0kbA
3cHhuqEN8vusEpY3W6aXA4yPzv5bbGho+6fAKX58wUIMG9HqtV+q3LmK/oWOI/f5
ddwGdcKqGRWnkVvLjWHObsWdl43n1AxOgA3E46wPE8mpGfpwXGUCWxXKi8ITZuzs
F+HV0XrY3dVIjDB2IgpoX4Sy2YYOBV1JzXeYjFV6XgleNj3l/aZouvc1tZJg1XBB
EomZgqOrwUs4VJ29oyTfqOQtQDwdxmpnG3GysKXVu7IJ8q1KNIfhYWp6HsMYLwuj
Y+TdrAXLKyaP8zsgEE74h3ccBbmzvs/OOGIMK1Q1HxJPLUQWzCWtsDqaNjVFk+Pq
A87glhgYEl/uxxt+GAii10Fpnj/Wf00EDZmQR2vkbIUfLj3bISSAcbFsbO5/4Y/b
TPnnREoUMY2Gv8F/Ojs+EN6mBe6R3BE77ImrTNpT8H07YHyQHL7gQE1P1uqlZHkZ
PI7aRITyi4KMSAF0JfBvfjXVYZsgmU3LfyjeaA+cDsVSod/6hJaL/PF5gspG/g2j
0fXEhmw5FNhZ+p5I1Nx1ZiucEvk4+RUeWSSPYZJ4bAf/GxHa+/qGirp7MSkvEovf
6wu4Xwvty6MjrL50ex+TWGJkWX+qYZyLK2ly2kLaKNY8Ce2qDtlvhNbovRL3UdKY
Cjf0LgCeMy1alN/wYW71awOfunxvPN+mEBOB1TyRMWzII/FYI2J++OCId0jF2UtU
oEfgshomdV+8zg3LlPpVdw5I5yekMKwsN06MGC0IGMAM1Ko/jePqWT+ouBC65HK5
8exMgA7g1z3yWRlCkbxTSa1H+622py0Qi8B+tyaFUYevF7KDwdL8UHlGDmvWJn2U
DTFQ8Z0fpg0eJTCIkJPuRno13kGVD8eJVov/t9fmQq8498bTc8R++FKgzsEKwrbT
3jEkENWBjwwqc/IqUqF6GAEakoYc5obq/JLFu2F/356Mqp8m3KjCzMWLht88UfTd
MLxg9FjAV3qUjVf7oT4dQeVMu1uRrgMQc6w/njxIdWvj14wcR1tPrn8d8wWV+b6R
3cqLL4otEKtE68KRUSomcSShhOv5jGb8+ij0WSCSMadbgZ7K+HLIitaL7XFKGSyY
IYIHvPS5jU816K9gflzT8jvHKSDTmd2eyZvFB7w+9H5jVdjZuBUtlIjBWW1xEyqT
2AphmsGrg4DSZp4PBSuoKeQJBUWYY83E5VBx2ivPbP39aSmMcpIIDTutei9t0QM5
E1GNNS/DKFEQM8wcf02ot1dFm1tgOlQ93P0xF801u4DTqi/YBmH6sau6xZEVdDDA
jYUWkQvTwg+l/VMePm0nb7zGsTq/Sti76xJ4mjSJovqyldIBKhE636cZNRQYx4bn
hl5bwXFHl5T4OXxPK607v/HeXeDslPoJlsxbdNTcgIWgRidVfINUb8c+Fx0fj1Om
Kl9asg7Gn5Z3iTvp+QGUWXiWCXAFepmd4gsCViD59/rHRahaK9bAI94Gzlf3kEzb
`protect END_PROTECTED
