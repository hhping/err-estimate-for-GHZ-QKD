`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/IzzZzNqSLXKkUuwiq3lIwmmeYmOzmGU+9uqip+tpgGtDzNmXlNVgzaZOll06Lx
xlmOkERgN+gv+8Iu/eUIK9k+7nHsIFg7R8yvc2iTrMyOJ/x0Vj0xwVohk70f35Eq
vWvPPeAf3+DAeS9Cl0q82RWZLoqzCe70xPh4e/J18yCdM0KQfUXVltzTOL28TnZ5
UEUrhcj9tmaSYPH58ENwwTwLclvjlVL0ANAPdZoql5La9875mwiqiRtF7YZk6APz
bS8cgkyY6gyE3j8Hb1usXiVxxlCdyVdKsUMqK4sDTkIz5K/vN5TLXCD7bn7K689G
GHTAqdDUr1FzqZExQSyRNEGPDCweVvPLxRtjMbIh90BIWMlwPXJt+kmjCavYICgp
rN8mKvCpUOoRHptFtNKwy6ZM8YEnZwMBs8CoP2X2i8X3lEI2iP5dEpdpkir5xELb
9ktm6tJYPGVBwW/shoMdvw==
`protect END_PROTECTED
