`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUE4lKFQDx+7LPiRuHDHC1gsGah7DfQlhFWMII+XF0YnLqnE/i9h9caUNl/NCoKL
m4/7VdaF/C14QzUC3s/sBjh0+QwlR0PlH65lTeS8wQSkeQEl7cYMLJJKvfjoZZ4N
BtBx4jOTkmh1D/yn0ISXr957bQvYesoA34LMJJoMWJBezYh8iO48yN4nqfsPd3Rn
C1V5F80cT+UOFz+RcEL//f4qysw4F2QhXof2cIHP29FYx6fSVf3wBVT6gEh6LujC
4GMcvJXomPwzpxuda7VYFOQi86X1CqmTtOPGeh9ELKLKULWOstOWXdoLJRSRBUQ4
apwQog7+jCKMCLA88cW6RK5QZJ7SlHveNw7BtElRx0tiv//mSi4bl77FnkMTKz73
XnjjCgbEInn8kipd4F1ATfLNE4ZKcY/9ZvHMc7bsmcRHCD2XbaxXimqhVt2jTRgS
cEqEknaQP7YSvEY8y6CoiRMLMExVAwcBaPlxEmUOROvwE9fYs4nyojYw3IlPfx3+
A3qg1P6inbIUucQW6t0NpZBN5DUC2IgxuDODvYP9LYjXGj8crUuP5WOMsyofPihg
uIc7HoRUv8Y47diq1QChmVKFFsGDg/F+ytcnkNXSY4QeonflTk5uVm92jHH1Vblo
h7WMrFYiYVSPo9op26PTG3QJuiIQE49OJ+FzQmHzKnN60PhhyN5dhAKwlozzjMdK
JongNYy2NWk2voMGQAC2ECLA4El0odJ9vSTQag6i/TWQJrwOXn0JoTvIdbIQEb7v
gF3VkuQeoVL43i6fZSaw4zclCfydmfaTlmhNtqvi+sq+wPXb+PVKJD+kj2YwCqiI
`protect END_PROTECTED
