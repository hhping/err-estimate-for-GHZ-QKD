`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2fOWWcdS7UVHz3kTmw6yYWAeGqvQbWJP6RghpzzedJCTXMc/xLqsVk8fmlpJ/UP
5PWFHL7ixGdu2WTsHrX/X3vP6UvVgGOc8gMba6TJO5ZwLX1l6fagKEok7rDtzVVg
hos2cIB6rKF69isl6IxD/Hy8qamPfrOT7wakJmGYGXjzC5C0LsdyMakZifSs7sKW
rzQRnMpDG7XWmDL5TPGuzbXe4uhKpXCTgqGCl0QSWFGbx1vVaHm9ArblnklhGoh2
esc9bp/dNw1bQGb4bZAJIHx5+8Q/DxXIOO9pO3aGJEGi4UYZBuFsthCVRA07iecD
9h5q1GAxbuTBfNAk0gkKWpjqhB6O1w0eP2vsf26yi2iLBbFUBcdH8Slcf9lvtcOi
mixPm20dStJ0itAocDWzjG6BtIZnFfMYfx79UFegD9Y/coCrZ5UzvvRZoGDyzzHP
mNBQxLDrvjmrpVSIsF+myec7zy2iVbb1Jb5C6g+MvHnOyQpqngMDuUR9osNbJj5M
yA0I21uQ/meOUJUsHipx9e5U4ryOkP6yThQnJWdXaz77sI6U/uJFuoM3c54t68/r
rouBf81U7kWqdh9/qM4g+Qu8pqRDD/LiCiir7kXsgQs=
`protect END_PROTECTED
