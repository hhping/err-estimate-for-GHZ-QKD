`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zY8f1rav9SVrgylnTjEO08PmvZ3VceLJln+idjy9Zzbt/GZzUeKRY43NEacytf2X
iaL2XCP9JQQfu47Uuc8G1aCyAOocH3zUZmrP0a8jKIqrbtUjTLtIk2TurxZcG04X
HGif/cU7g7UyMCH+izT6iq/Dcg04eH6iPjUdcPklZw2POggE5y/rtbGuIW3vuUl1
f/fOPooPlE1OTJfRQb858iDv1YYkOmKDgxEjFfLpCm/VEUDIGAud9DAaAG+l/39O
pWVqmP6sJPAJ8EFEyI/Ju9SFo5xXq2/wRKgc+mgnC8PI/fIB8xgK7nK2XeIoc5UA
Mfw1xYEM6h7anZi76cIcP4ddYdtkIPDAVz6HRW7/gzoFcdDV0alBjUKW+JQ7UTY0
96Ut6Z8AzsOl8sdCaABM277trLIHxgERLfb3z+Q4gLimUBlio4YgzDJ/QovZ8lIg
XdaGiOztw0glpQvIsEBnQTbtBgEoS7yEHN7ildDQyyYACygr+6fXTE8JEzskyDfw
+yy/M/Tcn5B2gfKkDxAoQ3F2NWYOe5cBHIX7tcSiPSs7Z5jz4q55KPOTdHO+kMpj
sLmonrBs+5jC7hDTHEQ5WtpYZmAHA7EqwCEdn9TdQn2yIVwUyy3FpsIVvIv0qGdd
4vZpC+Ya+egO54zn59n0G49+pIuQ54rtCYqbojrv+DbkKQzn11kEh00270gTWdnr
Pne/1NY3eNpyDCWLAYTMuQ+J06Va92ErLfKwIx94Q4w3sMt0BcZ9rDcAdCdQHJrm
TzPMJ+F02I5tjI1zrIUoP3uqwtwnd6E+82+VIKf3q9lOsqZp6Q17neQzz7YjYuhE
58uXhdWarFPU+a+mt5DmmUKBNI46yx9j+RQfBK5b0ymcsdg9XNkBsFV2hmvj6EFE
v172fRqcOlEe5zrVKR8vyE4dpbZY9RcqiS2pxmPbM1OUjwmQjtrEzPNWWhojZz64
RjFaQ5sWi8X+Awf/gnNdufE3cxNgU62fTtcm/kCc02YajWCuNrCoZcl1eI59hLZK
uQc7cC2KX+Z5Wy0INGmffT7j/TC6NytujewiIsmh6JraFjWdSB6qrobp3kIDXgv+
Vz65/of3g3Fo6lvnPgE5Tw==
`protect END_PROTECTED
