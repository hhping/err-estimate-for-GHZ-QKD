`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqH+V/p54bZQjR1ZRlpPV7HvswKPwMAxOScwKpZxDstIWyD27sf7Vxw4tfzwH8oq
ZHQrzgKdwfL8O9orVVjbTnn3MCw04IL1hZF+9cjNMmO+DXX5p7uIalGXdL/VoZkI
DM1T0OkNGyAlxaNEjY9UUOrWAOSMpwnpyd0CdeQiEh6L2AqOXGZ5qY0quMgujiLF
VN/fhRWQr2JjrNsyJ6rB0WKObgw6hPO8zZxNJvB+hQImvFGH+S7QpApZ4K6hNa2m
YN0s7Rl7qRc13II3q9Yzyw30rKlBzkJFrfFWnJKIHPwnyfepZ4gvASYSFN77IrfY
ODDqX9s8UaHrLS5smmXgJKq4eA48ET54DTayb7vfll1LoqDmAkXTq3Xu/NG/WVxM
BdiwWAohqqd+HI7lkgkXaLx2IJjXhLZ48yLHLkPJlppYGjj/P2C+pSaikDYNHmgW
a77wSF1mlOnxWt6uvCrhxLKD4OrzqZWZVnlNXSDa6kEmme5WVbRSF67EAohgTw1C
rU0Uy/oUQE+ccIEA7/tet6A9bImLGB88yzxwiId6yyDWDVuKFa3FdO26arejzs9F
mt/nmd3nbP2PTGfz7zb1cgTTKGGS0w7jOluDQUPBaSyzDI74zvWOtH0FAnCjt6oY
ZdKjoJ9OkEbzL0q/es3eymQ8t1Ra+WkG3pco1+SYhVWMfWdOKeUk6xZVfpejt72/
xliw8FRl6yNDJFbPw5LxdWlpHpmW6pgIA5bgYgiIayUMtKr2F11n/1b6sWYN5QPB
7JxEP1RgwFCU3vciqbcnEgy5afcvWKEBczFsnoJDCxER9mociAfMNpPTGZBRIFY+
c6keiGJBWlvj9BftWtck8yymh4yvfajaxIMomrpw6JRYEP8pQg0BRiivjTm5DKPP
6m1bO2ch4ZV9NWJ5T3ijReLwQIirJjftS0YyS0w6nJ42dNxvCs70SQMdQ+Y5o4iB
Hc+nCfcoWuBpdZZAjG4fMNKgHcZF5T6G6nUGTO+Aj525GQNN4up1tlAj8Xw2Ncmo
MC8wQiMtPWZDPzCTi0PrM71gSELtkhsWRXYzc+mcK6wPu4uK7zfzGxgjwPftnf40
xk9KFPuBDVNuOs+xSmbzR3ZL3reKjHlRZq9+CfH/La/xZpBHJNiDG7omLDOAcG2F
yTKMs5frPqii352kqIU5850oJoGqM87LwlReQX9Qz29Ty8xIatOn/Sdg0z+vRpPr
WwTxmq6T2/GYk4RxEdF/NNC7DmdJiWfP8DpUuV37e9V8mrLOTt7vDeMW/Ouxt8CT
ZqCWGmOh9+HqM0P2ziPLhTJ8egXaBy4CmLgtua3ZV0bEbb+EWnrkaKyOcjcR962n
y9obNXju6P2WZhsnAjNkUnlhC2Qy7SpD5YdI8nUMoCIyC502vDMwwNLaUEIiq5H2
kGw5rDLHsKS3FXuOP0jI1kv1iyffeeR2LfKkitkhTaepEr4S8mT2BZxZPTUMKIUK
Zmd/xaWCDVfDRF5XGReMSQ==
`protect END_PROTECTED
