`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3TjkNdPCFBnTq52qgZk1l5ntvM+DZ5MCOhye/reY+ncqQjOfM0FJCrtCAPFDOMX
IlVL/bzwphV/4rClzaGEWTUMt5Sli6bCea2sZlO1WXFUN/aG9yCwergPlYp9c43u
90uAESKq7sWLYSND4V5htTRyMvyCfggxVsrtm6Fc2/BeoiDzJCYfXaMy2qv38b9i
BKGV6VPlS57ntOcyapaCq5/jJYCD1LTAKlXijCO32z9TfGKHg57tVNjRUKwuaVbb
zLY67YGXv4tk2gzrqG//nI8rGLnv6E8CmSWBKbySnO0Jg3mQh+Lts8HHLjZhel2L
MAgMKo3zU1FQtHn3Ztp59/5JcIYJlpSiFmKsV29bVzSO2mcR8qBz2w5ZbGxClT+y
4pz/JIaNuhzPons+fOYivkNEW51F70wxfHjOgEnOyFvpafBb/7rhg1g6HNKBipHo
oXR84Kvzt9JD7mvtBbW9lJ666rtP38H1Rn0RXDok0Au4h8l3TKCi8cEkkJ1LZHmW
YE36uWrW9GKpdGhUrGaE6RfakyNO5PTKsFXOmRzIYaUybHPnl6eu++QIr7QJcnru
+c4kT8lACMyWcpVslB1QBt6qlUjNth8vek2bv47y+qdpnwOcKqACH9ZXxjHjBHiI
WFp/3gLaGOyE0oKgqqRVW2fM+KyZDbsggcloqbCeEaSQrzdrf7FkeDdGFvm4NVLY
tmzMvPgA2kge5RVqDSeyA8dVxMgOYGJYsL5hFYMW1ouRg1VYDFu0mm2CUtY9n4zY
hwP2GdpA4iP7ccifJEaZMmcvcGFOn7oz4wgDPbNn+Q/656kg2WOoWa/7roi7EP61
Bze4vmNYS4fZjgwSfe3JJIP0ugB7wbpP/lIl9DeYkKmXaNnjP2Et/aMJnQne+LkB
WfQsCbec1/LAwH+xe7BSNtSzn/NE+jtKdd5rPLXb46EVJq1pjqk02XrFK82vc3FG
OK1wz6zUXm7lt2I+8apO5I5BVvSm6ezvsGNjoug3dTZ1cUm6d89B3X2wws0uf2s/
zJVMrdmfxZ6KivSNSaPSEi4pk/Yz4cHcpAkUwKkANRKmpF15iRzzTYLW7x4PAxKt
4RCapxgFXCKzN8T4UO8UCRlYU1Of0POv6CFDqNYdG+opqF1vfkK0M88FTFPaYdU0
YeyVK80TPlw47O+2WaYbVY5NP3enJHnM865QyOWKNVWNvlGthAMEqtcq7MIWWw55
HvUALLIConfitAB89FQP0wXXCzIyWsRXGqMbkhWqk/gNQHuGYbTIsYsHmhrWOcC4
125+W5NC+Fnx1MXnORw8HgbhziF66d1gGvZbEAiWeKuyKvDC1pllK3PcYgpq0/FE
Ubei6xvRJPA3rcVkPS7sZnljH1ifCO/ZC3hfM4zMGfRMfzMcANaY5/BqqJCKSJV+
L4eQixB+WS0bgySbfofNfF3Lw5ZlrtQyVIbp1BQebKQl8SCBfdJT2dMK56UKvrQG
lJFuUJMm5E23tWFxgfLGyFraOJHaerRfiGof3WTcbQCteR0cxwJ6k6njtSGH0IZ0
qwdCYrvVRnrUgaYPSFMIrFzDxwF1OM61rzT9CjxNtloG/0L2YLsRAt6APjVNzyrI
sUSdTG1j48WILyKxUdy8gnvfEAaDeKQ7vZgB8sAO1z+exYVPEKe+rvpp7ocMwxSk
BIlFx7eYDrRJC1Pwzw+BqXYZeQwpWdJaGT78wfIhkBeapjTlBemj+mYjpB4qi7yI
rnKlfuBZma3dRYy71ILngAZnFw1L9wUgnG9MTf0+k3dRu/ECHWxFZXI85Hq5i2tZ
Ar9MSgGSoeuExWqob2y+DrBGlyk0WunGxidVvZZsD8R7JiQcqldH8161WZ/Y7Owb
NiQ6XZ4XV5mjM8hFsVzuG7ouCoU7hEuT/+yUvhYiH2acR2wAKYwsxzAxfusfqe8r
RvVji/xEvlQsW0WvW5J/yj+0DRrSeE4vu2zg+m05dT3N+fsOuhhQkLgc50xcwklv
nBPwI64JQDmSJrcz+4ykqbt9TdbtH9N2yMl+2SEN1CVx7d3ZwATfUA5rrqNo3m46
KO6phWiuUa7QClXSGex5Ggc9hXijXA0Ww0YgYW8hZ1SWjaURuUOyAI4LwheTF/4U
VJCKFiNFUTdjWaLNIm52xKtIQCZJedGhXsDWmn3bmt3CFpDDPtMMOOZdrQnaEqk4
xCRhaLRq34OFngxiYGJGoFtZFyyKrlpsBq5aJWjYouBu5b+sXnhZiq6c4P51hU63
lPMkEuG6zGC9DtGQ4DqRL+q0mv0S3wzoK7HabVKV0S6HRAD94fdVGyR4mGK6TJ93
CeXLh/gHAgtNLF2Yx35El5HbAe6cfwv9rzm+7sPwmS7loD6MkbirrX3vYoUytGIr
Iiw54pHjMQdmLVFyCzpCmFUit8dDW0475YCVpomFYKxTXwCU68/BJWYndYYy7AaL
mH1jf6gObOxmyoFfsT/kAkNRKsied5Clct2Jz1VxqgZBFdd6pdcG1YSlFnr+v+5r
n5wHlg3UuhpTQ4+xZj39PwHY1e4Bv+KGcoLW5G9H0uXDBBigJEi+UZQIVKybNBP6
usygB9uTrlBYCTUqA6m2gsZG5I5OY0AnayBsoMXL1hxnXArrq0WXZ//I+jotfHkt
5H49oXbFpmiADZdbCJYJgNdUOvaxr00c1fJD/yHS8as=
`protect END_PROTECTED
