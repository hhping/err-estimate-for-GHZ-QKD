`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6cEYk8gJWslpN929OLED7z/KYn1y3OaJA08W0ODdczXiWQuFnQRUz2nH+SwI5u04
skS2WNisTywFnjy8MBrrwzLCQxZJFu6X80NG4qxyjdNZyonOslegm5pmcdkXKGIY
ZnNasHEHa+/Oo7vt74XhNcCRxqO0h1pveK4xP0arp6J7Dif97ctLWuzik1ovU+1p
xk8dBEBVzKu4VfbARo/Cx0wJx2Rgpmzm+PFBvcKl6Q9lbMmEer+HOCatviD93UJ6
G/OVkSHIQP+u8IiJ8vEaRkAZHxFbIdEBWAM8Utn0/LYIXJl2mgMKKVGr7NFV4CN8
acYNAmYthBXs3By+dkrKxHP5KeLe64IfMOlZcc9fVohtp6aYZYzsb8K7uBcIkjql
+32/gmZ2HiSP3pVgjp8FHISRg4TjG5FhkzqrMd5+MJJL//T6L+IOofJJNT4Ucqsv
YDt1RZPYPDBmQAGJZYwD62vz/zF/AfcFf+3QGadVY2G6LN4ywXaNhS86dc8RrUXj
ZDlcvvUZFucOcau42tRW4YFJv4mAyY2okiCJDsjrFtdXPKU+aNvtZgW28xUaiMqE
313CWy0w99PUmvuUNCvCn0NaqYFuL6b91F0AfTUs3wPo4hR4JkR6/a9q7wE+6xdo
S3whDtIosbw2EW9Ag5RG3r+GqKs/zUauaX0J+IJqX2LYRJhoUdIBApBV5paMNXly
oeuuRSjeVLHq93R2HGE3XmAhBKrYrVg/AOFhRkPWxRHt0W0ot/k9AdbBJdFOvmCB
hBdmiQp3lEdrJby/m8JgmlsUhPz82PAopzlJNp8AIHGR+6dxNls4Y/gYz23Wy0IQ
7m+CRevopzc/pNO9wRdkCfUDPcXyvhZLNrWKJ6Xmem0mVDuK2oFZoq2wxv77Iino
en62BtQSJ8gUMxLTT1niBPwVH7iou5pxdg/gfqjdE23VXNTMZpQKdqbiSCemrzyb
ARpo9kWGbDvBb9qbfiwOKHtLsr5HZIxLtjehqwXRIF73GA3IcZqTF90leWsaFVz6
4q3AH4DNAoF0QqX74SB2pBb5+mje8O+Y+Gih5LHIeopf8ZNGVRegZMF2u+D8tQHf
eqZIkCCkSk24N8EkBlwicrd0cpJO9JRcTCUyY8aZOHJU5e7ANT1oyd+oE+GaGTDj
VdWrGJHw5Mkflyc5ysDHFuE2GRMc3sV+mM2L9C0wMD8=
`protect END_PROTECTED
