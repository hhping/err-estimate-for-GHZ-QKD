`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9u3H7ESdD/2yHq8zCDXhy7z/J6tMZYU2Ph7/ExCXATBDEulTUt2v5G2XJc5IG8g4
OOKUQ7WiLFGHJth+0Sl0sIq+NLC2M0AHrgNIeQbr87irkCBLd6zHm6xja5qOfIvm
JWGZFxzlNktX+zxK4c3r5CBJS0CjiyWvHKesq2dyKFH66D2WD26aRjv0yHYUyClF
rfdudl9HskzzeilTe0MQEDIOTXowVHIYOyLzWOgDu5fkvOwutWcaGY/2nshibWXr
QJG56PlWGf+k8hkhIGguz1/zGD+D+SK58aCJri1FTfNxwJ8jeKifXtq+YG6PYhXS
JT47Qha9vDnEKEa0dBtq8WjNQnUJLkXYnA+9oURbw/21qHrjSuGdoO4+B8zLzfW9
/qn0K8gazAnUQ0CjYgMEtH2WgPsfxl7sqqKUzbaiccvSHlRJnrcMIO9/xqiuHZ6e
jGbl6j4WU4NOZNvcZ/qZVe5yW+f8p9zWyvJSaD9Oc6FS+vnQ0FISwAeMkFRpwLLE
9p4NRVlz3BSAUWdlUMNOzkICnGLKREcQbalOELyyx9Jp8SIq5yw2E0VBMGMSQU3X
lTmue6EqdaCtYBKAgydvvZeabBuTYgVkKCC9NxaXGwc8pJows9gaSWCpRdey7NBA
qzNUU373nW/EkymYHzfEL+h/eAYcuUUD9Vk2lku03v/SrEzHx5XH4wMbS543Euol
xUfaGIRiIl5zUlsYa2IgIriPO7YfKfUO9yLAE6BPQja9eEG44l3QvXkPomAxtvO4
tCT5lOBuKxu404zBLb6M6kYROzwdGOKev7/Nyu0X5v/cR3P8rIE0wAxmsgkZPv9a
r3aZqPZ3AOqa8QIFG31zo4/o0HeWRsAYDJXV1lWrEDRbpaa+onX0znIzYoe7O8Ez
MY5/bfvhBTpLPpivisMMtj5uIU6QEJcfkz5MljTdkth/DVIY7C7bWj+WDvkzZfSI
T5LvgqNep/ChB20xS5E4vL5DYTQetFh8NtOBSnh3oHPH871r7aaXGTGr72r0TZaT
+ZoqZTAg9MIIarFwduwe5/btQZFMiU9zEho8SCqkfnlj4MFqCK2IKHMLkh1GL5bY
XXJzODf2Vvwv6Yoq68l4g2Onu/iJ+ZehdxWDCe+VTjco/EksvI80tOOS2PXWm26X
8qOzd9qkMGv9zxkvjKUvsMQean6nocS7iaSP+3npdqRBQbaZNOAtrchThYWevunz
vG5seL6AsFywNrI4PvNb9pg73AK5f5JV07aq2ojYbTekOqje7jJXPjSC/EOEn1qu
UODnIOBJzoB0/YDyaRGf8vbEA3wLENv0K21nv1wIudUcNs5lLxrC3rpAMYzp63RQ
RGBnu+J9YrP0gvMeCzua8L1P42ymb7x4xeiz67OkCTPOtPFnwoYNskJuEZuRYe6b
HFMqMDBzMgwUeY2/D9Zmit6f90OiJzohl3CrVx9fJ40TiogNwWorw/caiBLq4XnE
LYGww1AfZ8JxIihLPapwGFLPHRhqyQVtPATyrvokzUeavusxspRswBMqPUXhbAqW
NxHJlV/IG8DqlKapx87h8HA5QAvXdK6JSUG/JK9K0mA4iOPihKV0XNeTfQKBNWQN
oIRuYI3UxsCVfUcVkfrKtV8ydtStApik93tzy5olrtm8r8NmVxMWkCkdoO5M0jlr
3QXAVgt86OD8cu7C4ZeQrWJ17fpoOG09smtbVrAtT2plCPI55Ho2TGaEHEINJZAC
DWjrKNOGKfgk5HdqQXcOU8FCxbZElUHumZXxK9Br/EAnJVsmvH+CISNk96z7yRZu
m3uwOjYXGDq8SVmWxYpl7w==
`protect END_PROTECTED
