`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5Zwg8zGTuCpGqjNj5zUXWIzjZG3n+6lI4D2DsWOQFW0LeoPDT9ll8P/DG8pUEc5
kuvnq5m7Wi9VmiNw9+vdFUtuz3P0j7MOXx+gj6DqmxGQ94bNGbrq6aIi1sN+7d9o
cgjQI1iz2KyUFjnaX3BdERQZRZM45XOgHpENVHx1INNbPKF10DgA5Xz6BgkNM/nl
wjerGP06ooIa+uaU+j8llwvtK3/AkaGc1QTXUcMRHp1DLNP5QNdEydWfAstd+gBq
QWyJGpHE0yZw9Ni7PL5J4wREZhdoR7HGug8d+jjmYohr9k5Udmc/+UGoYw4Xjcuw
fDuZNUK6ag52w7ST/8qyJXaFSQmLO/M0nEmjK6Azv0LMDYwZbX3+ZNp2DU6uSPxC
xMG/DCvJ8cRiESHlsq6c4A==
`protect END_PROTECTED
