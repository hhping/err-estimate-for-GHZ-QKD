`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2uNhOCJZaiTME+GxJjnxwH3lMy68wCgzNeckd+GRyE01kO1guEnS51I2mINfWZ7
90ZkzbX4eNoP3Bl/JAtvUDYt+z96u4MvQNb+1C6mgHNnsCuGP1MxrbEKHfladP7I
uatxAzKHjYBRdomJQd0Qn6GR7Pm050iNC3x5tfzqes2lfXDchObsVdubC+EDbxot
1rXiZtdwVcHoxZhi/8pztcJ++RAHvPYZrHtEeYb9dixZ7Sxcz0kAgjjutUfAlLUz
ZCouQ3sEE63YAnUCUBDePuUAUsd9AA0CzkJQNW6k/cQEXuX5n32gDyi+2zYLW4vk
+5TQsb/THGLLwuCqfNLf/M69nMPoH2sGzoRkl+oRrKvc1IZUVRFqrH7878VgiNll
6oqy+K3/RvArF55YDIcntYmv6g67yOYQb8YKoEhQ6kg=
`protect END_PROTECTED
