`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9daKShqVPkOgrE7k85Qj4NLyDucqCVrGGgu0QHw1toUtrPA6EIBn2TSSKsqZeK/
KltAAUSmqlAXXfvkCJU1iFXMyw84wjk9az765X2QQgSG1JZdOWb9kXiJvFVExCQM
rhPsBnLJd4iO47bw16gMzUCrcZMn8PD+OE2wSLjGrJMLRbsBtidBrqG3uYvy8jwd
4ns2Jolodmc+6mPc2KKBrjFam7Sr6X4lZ8OfWLtBgxTu5RgJnl/36icn1U5dejfd
DeUs+a12JrKW3C7k/mK+zi60vQ+xhh0TzscSIq/LjPjb5M8bAc0qt4w72QI8l7n3
Z1qpK6vHETpVqbqnnlkeuRKKNXeEh+WQWlXR3y1+YeqxgYvvwpYRdh1bz6zMZl0V
eA2PU4wB/g52JW860AH9BLY3lXt8GBQ+lepUrcpVW0FGLbYLM6ArWJNHc2DlpfY9
4HrgeFwrVw8SDU3gp8vQ6gvgvWr/b8OMKvoroaxfWU7D0XvCISStI31sJgH2N6Ie
lHe9SYx5OI8AmO2Qtqyd1mdPPjjYpg8ZcUFvsaVmahDXELmj21aWobRmKvyTU5Xw
aSiobWEs9pkcu1/TWymfdo32B42qJ+zXHEjc/yFALAJALN0k5X08lYiqZM4cCZD7
hmyfj4BCrgyfTW3aqs7r14AtkrnO70PQCGa2ZckEISbdNjFUieUxeofWAjDa+vzS
aYcZiQavOOuBX/Vurj3tD1Y0GG48CmtbZw3Bcz6Fb/LG1Dr8Cu4/NpvLka3VZ/qi
6zizdcK9P1+GSbtVSCx7FRNHfvG8IKFui0ZUZEIygC1Zb7Bl0NQKAqXU+Nxznqre
lP6QiEHZYLDvaa6DtPDTuH8fQ4jcS6n4vqbkoL4A3mZly8vuIkkyjv/RxMdhHndJ
ExiAdHm/PK6Ot6li3RRjkMLmNSseZAXlg2W0jIAluB34P+1Ncxo/ptR6CJDxfWYO
wrSOTUfrnhRRJ8ZKO7PTC6PNo/AxzBusEzP5qQkaz3Uybvg/Lljp9EXv/FAecPwk
Rm5a7kqe2VWI+rH2Ckju8nI0ExlcQN7qbfXv44JNcDZwNUQgg5OHOGIHuo4Zns3G
REYIj6V29lM80dO1ayhU4ndCvj7mxLTD8C+6DjMtLas4uyI6YJTg/fPYdghYe1AX
7ZwFxnk6hGyEs8+NaBajh550VzDDMpPPZXQ97rtw5uD1zm/RgvogGURcJ5l3+//c
w2lJTpP2EL60lxGN1+QroiA2CnygnIFQvbMpEUcXTQGawkgsyWOfDBreXNc0lJEG
0P4zfDWFNCYa6MkKKEhOHmOoSTQ4xBKm2f6PUBdBpNpkhEMiT0JOodn3zVldw5SS
3wGJXXSgb7CgO9T237rbunC8KZ0eYlJMSJCvSMWQDiQBgismEzQuqGGzlwHHKO33
eUF8ttZPRNk9iVOexYdQzaKtC/snSqL9HJW+5nyA7zTK67LlElEHf2lPl8cJr+xk
mBmqXU4EsbepLhjPWoEgVKJrG9lLMPEXFB8eJZSm85Zd4vi/mVaJvEudqOTqybrO
lhD6PdYUzhvLlwuov+IB1pjzU0MF0JUPxwVgbn6I5ZXt+PfdU9xsLj+TTSOPO8eR
mTbsLklboSrUtuN/F/8XF5s0txuffRLuI9l8i5fUHjUzcKmrRh+J1FqeKafSfD0+
N3bSnumrzcpB4V0rnrmYzJdgPkpQJi+FzlzAbQcuSzXjfmJb/VEcQi5qoJwtuaXZ
9z40N+deAItL4kORYT4xaIfYyg9yN193irskV9ql118ZVZBA0G1/CFu96qbAG8YP
ECUUql8jq7KtnaSh8iCPCBs1GB60IAp2YLh2AW6LsgCHYlgmCAUJ4RrCEXXEAJe4
HD89POsQZs8fAMmXe4evyeFVR+SUbBGlEHF252KjPzgJrI0A+FW56chZGS+Ynx3a
2JKrjkb2xPj1fVXOaZs2b16xd5l5JMCDyIosmkZUlP+QO2sJQKeW1j/z8maQDl7v
E6AyXxFhdcOaSEcxqgYUiuHegFsP4Nf1714s6v+CgPHGPtFb/rDBHfxKaRJu4mDP
ix6GcrfMcrDA0xzZziO2V4m738a0sfuK5TPOG3UGKG47v/5ztffTIj/EsaSIPeEG
+xuJEVh1SEVNqz5eUShta/+ph63+oTop+hZvHoVV3ctEJIUmzn/KfGC2fYKfHHBj
6IiWR46+I94OBxnJTDiaObnmwfgs7csO7jDjbNoJsUBvzftUZWXrI/G7DUH7dcxT
BWHUDWC1078DYGvo6T9ISa1lox/3JJza8UPnmf3HciPrT2kq4ftQCc/lmG5lVhbt
4gsRlOHWqQYx0w3iso6FFMW2L7oheK8mmZ9HTCNIOSSNbFae8l8Y6PSXWbIHwJUU
d80HUTXBAFp7Ewdb9gI2+VSJ9I+590U2ZWn98PzB/Me3B+xKYbEDMgf6h42i3AMc
/y0NW1qkQjKOMb67ZM8WdLtAoDax2zlJm2r69xzMAQ1jzdmdSjvI4NPrHWmCJzdC
M4AjFmCJ53aznurLU0zHVQ==
`protect END_PROTECTED
