`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHvBuLTq/ONMtYF41s8CBc/viQh0J58H/Ep7jFN4lVUT3Yp0qIs1DQ0ncsvdMLe+
AOnDJGYzdO1TTD/HEYt8h6c8vKwrLZH/lbtM1MekavVYHysEFTKbx0n+FVJONfg9
nkYiOkY0LyF0MVm5BA9tJK5ms/fgSLlletXUOP80/8TQD4VN9CaAHv85VivAkyE4
6kVJk+yMrrmUPvOMn6ouSbbdx+1tOCasekdqgZHWc+Ogi7F80b+NEwSqNFY+O3J3
8ZvtCEL0rYwJpJnuSOPJObRTCmelLuN3n1T7jqhbStECTO5Kpvzlq3EB8Z57fKnE
J6dATgANqzxlH12A0PqVUhlXwDUrmkHh1S8b4+WcohX7B9ZfbnAusFg3jl63HT0K
7MSr7b8fHloYADrILjo3eaffDiFKyfnpYZYArt5iDRuSFZXX2a31VpdGbJT5lk8A
Z/eA0b66qMH74cR/nvwpteGJiXsuO7NF31OIrMEoV6v71apqejnbm6INj7mMCL02
ZmLgNtC16D2cKDisFoHf0hM6wAmcGFu2A7gzRIyyhPrQv57lFUhVTxdLtZHcTD9c
Qo9XNsgUMvDydWPpoLb7wWaBjnW5ESrgt9bR8iPyVxmFZ4xzVR28+fPwBfjBUudQ
vg1/ROHNEBOQ6knwv8NQ5xLG2yOslBPFOGzkLSlGw4tfMdb3rl1cvlyAB3CNrWLv
nOFMbPz7y591ebPxZYeN5W27yGM5785Lnt0P8FdVcyRbLSF9uRHAKAhaRm5sZzmv
4ZsnwoMsQz/hejJJ99MBpexfSN6DejsdIkU6E/7M/gHnnyOffzrZACYh95PQrSJO
KN0/4M+0tYWLLXl2oZuKY49c3tjW1IDqW0SOUDfwXz+etaxBqw9SYIzrlQ58Jtc6
kowJv9JE8b/Krb56ai1r91rRu0TDXUjuFGYXJRCHBYiT189RjWXFX9dJnZlH+21V
Oktno/AvPzB39IOvH1A04mRteq0jyughporRk5FnAKZlyQ+DcellmsyDjN3IE7QY
PdY85mF53KjNYZkBYpMzAiEHNSACZ+h/bxiNSJZIZsz66tmYi9iqgq7YVTHYiHA0
5W+SimxjuzuuNZkAKlXfFWAYM6Yj+yc3RDozaQAx2rP71oqWFBK4Q0QwMBB5up2h
wI+LW0LJVEi4chSbZDqIASMJ/6gKm5tHmIHQvsSWRnnosxRK2ILOaSuZ5vBIrrLK
aFIq92jP5MWXVfWfx3wGvksKa6DCneJxEv9GRziOtsHQqU8ig906UExe0WOqg1BU
EqTmKJUOiyymO7REiBiiL2S6FgFw7GQHBpVBkd3JllOkQeV1CTxDywU92Ok+163j
0QSvbcPv7IhRg3A+Gle4oa3f8jRLziM1YR+EJTzChie+V4kK2r5Ax3WSbFCSDJ6A
OLY0BWHLWhPcRWjx5ttcVxeYjieZht0r6UjfWKTruPp+IrTAhm7hGN0bDpFfTS/1
jPXXJuc+H/724JVJNBpHSRyldCRqkjFTv1uEQ9dSo6b/jQ710Hu2CbDUkeXEAZ/k
kdmYjYtV5EVClS6eoAoA1SDrJ2aC6KUgWTD3F/IYZJorIJJlE4d/p5zOQf3HAgLF
NiODmakAFaXOyXPyB7qPMaINpepGm5+ezCXBBCHjFY5zdRu/SaseHiJsmlsadC8P
0twYKqi+eRszOxndr98eVJhIFdVJ3CBBHMZTz8Xzx3lMKo7cGRooxUnxvnsaaCfp
lXvC4QY+y1Mzp3W3XC0sOgOFJQs3Lr6GtKoEU6bY0Z/nT/OZndnddT1Nva618sAx
3y1lNxXKi4U5y+bfK32S2ZhZ9o+uOdHpXCDNMRIy+wsTxXdifHgWWlM4Z584hIMn
tbfXitWEjVbphCee2W9e5dFrjMgzrpAA4wpidl2+sJ2n7CXX9TzyLIOLSwT9DBAX
vPrXSi8ua1R1l8w4KS7uKZfdx/M+e75Za0+2DnNCKuZgFpW1hkRlQzUW3NuHZ5o2
0Rth7z6rmvZM8PjMLJr5QoUbn0EZA7ZojhKIxTyMk/6iGYy8PQP6HFLg8e5DQGZH
6BBGZdu3XqIbV4rBtKpiI4OrfSkIUu6Rj0QqR9oDiMvhouZwOcrO1pkfKRKkO+hU
H8iOa5isW6hJSYrLfmIgQa3zXUIql2o02I2d0e8/+K2HJ2ZgJNp7cR0BX/tIqSD0
b7pkOZbBjffBij4ZvYvKRKw83eQD1Y14Q1kYL9V5A4J3OSj9A4qv/78UAo32viMg
JtMzWUzXlnOm7M/Aclz2r4zTAKIWRCCSM+PQoHwxPn7fN01n2O3SsM9ozXhlEN19
7wrH1ZoKz6K1JoGTYbASQoj00d8SAMQxEF7J+GlRzHf+SbWmhRkNCSY5uIhuke4q
GcQdRRaivzuVc/7fZOE7AfjWjgupkizyFCfT4S1sCgPyrGdB9QIfG1sAWWamXwyb
vrgk3qIJ6DTuQsgZRmrFmExT1SimFgU7Zvd1xYFfctTOCIZlt2i+55lAsEtCjQ/Z
nyjjkN/2dvJsyGJKouA8/U7K8W+0eUj6rqQmEc74phcdEzLmBepqvS8vrSe40UW8
phI9N/j/AvTvXmiG83UAKX83UGPgh0Rg3aJMUR5faqkn4luzbdzFAoDHCRwYj3JS
CGKLPLKyerpKgY92eftowDtO3mmn8vdmO2G15OKEfdiL3/2U4wOrNVpArw8SpcwQ
zjoK6nP+Qy5HDdKo0Z+Ku9mFtB8ClZMWL2P/szV7VkTQ/0jSYl+4+dGAwqEHGZk+
Rw+ZFCG2sUAKUTwFEk5sXVwf0jhy5cS0a8FhFHzbs2HqN5h2Z8WuDum2RufoSjxD
mmjJbUXErFdeQAto8HYGU/zgVQaq1tw9tEVlgIOLjOWk/s0V+eSUA+scdVInfIIx
SyuiqldJVikCQtMW+CXMVKzkgGAlm+IGljHgdr840Iei66JtMQE28pjqBDT+TWrn
gpbAbwjSxcvGO/+6a8UQzGRt7fkdRSUEd7cDciQb8aezkPYBGjoZiJ5ilYInle+C
aZtPFPPYDKr0VRzVPaBiMO+6YXqN/gmvJFPD4fXzxIDAo6wYnRxgGF3yN2cPb4sX
4Hlg6jGrdhcWfSpfKaW/AikWxxmlqMXNtUxR9p4bsIHQLgIoKu8h/vgE/OEPet4I
CeFLSqiv83L/rHU2GRHj+6Ub+LXR07v6Rv21Z1Kgw299nW92U3uu4adddST4lL6X
5OjQgiHxyj8vjfxmSDrqmom9mVgIBnmUsVEp6XSYGgzvG0sMZC9+d3u9Rv2twnBF
R6jsXex1gDGeu9C+NVzCv42zxnbRrt07VnrKOQfBBrPxQms9AGG9EFj+JbtSlRJF
d2KopBFuH+RZSI6j6iAcAW7h0G/bk/V6KRu8sy2IdMP8ZU5dxEVcj03UJQd3Y+Q+
YW2Q66QRxGWYL/sC/vF3/2r20tS7yjDEmD6fBaDSS7b3H2xCZmvmQXoyOxh1NyNm
WN0kdWnGxpFmDViGcNzBx5W7B4Uuw0vTXf6k5LDCvq81PoLHy5tMM5MgmAiPtfBI
GFcyWeRAxSPAGp55KjKdICQFl3CyhUV23VGbyYhNBuJQrF9mHHEf9E1P0N/E5Fmp
lNr1NNhfEyDJNZRX2pq/C3v4eE1E1f/SusVfE6Xxtil7TekQQH4H5//ZOdWIOD+M
iiFaa0zTDOfura7sNssL74Uq7Zfu/PIkXyy222XJd4AsrVcgtFAzHoWwlPMHZfew
T4EFn1T7xvktvEr0MDWtP+NgQm84D3YBdQHbhp/kwVoRz5zpvhTtpFLrANEWW/Jr
kpq6yRsNF4FNuuydd02tljtKoGEZ8kZ70APsaOb/N0xaUM7dbA34lNSbDVHY0Oii
fWXEswxNHbrWcIT+3sKyYKHprwS2SoOVb+rBPqOdMBiHIBEZszXqgrKufqFW3PEP
zoQOUJXki0Nz+be3W7i/Jw==
`protect END_PROTECTED
