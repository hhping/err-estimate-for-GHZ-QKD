`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXQmi7KkG8g1SFnmGTUvSRj0ei0XpJ+uXEbv7hM9jAX9FgESir4XPwJjPoK5SLBD
5WQgZrlRuNLa5o0hVD1GaCcu76FjX0VgVxO522HGw2le5FeRDRwl2bpMYtvYnYX5
Mds//34IMDbxODoFI9lDpZxMwl3EHg1NyL3wlNM9uvZPs8Mg6dPBlHyqAoRhYr4o
O63UgCOdbuTkrk0YfpeJurgAGWbrCVr3GuYoDfK32NleU9W2UPDfcQL+919EkKbn
ScQuW6ILR4I86GKvjG2rOyd7aYNtyDSH/Ox9dMzeU/3+mmsAueQ5fCICuMr+dCyM
XxfyfboK6fAHhRIlUZBOR665daTWmsoK3gqNVr8DuzgdV0yGWbJlZJ5iYCOyB6rb
3KPJ4g41c0yHlcKBlmoc6S7JXDM7vuEOWBwMMue89UHGaPe4wRr3iqiQxsTneOyM
cm5YfrslydfA8gJMxHILYcZ5VWdoBi3GgdvkCGInadk8nlKNYnG1Nu/JGY2Yp4tQ
th0pG4AcQALG4B/vLbn65ZYjTuyTerhWiayK9B2jqc3IGyy7yg8O88xqQrMDB8wK
DZTz8MY0HSBFLsL5ZMM8etA7HumEnmIHAC1yU1NEY0iC9UFTU5pzggTYlHkkPQDO
aEbrnGZouvdVeDCpwVa3h5rEUoyGEDT4+t1LQztsoNChZmbsPzyGnBg7cFNuq6pC
jIubJ98RVcT1WTPl5uW5n10QGV3Xa4UxMHO9lsYjquCPlQF4YsinTMmVZNKj6M5q
/JKbnKXfw9ucffLIj4ezd2oX5Z5dZYpF1RMnaIC2Hys5R61ad2QODJ2duMX23l9I
nalFb50/xGDnAzuuU7D+AZI8RXlrj4ZQ6xwyIRLBaVO1MWhWtOGZHtCkWE/gGuRV
5c0z0QSoTrfIyj/pH0hmTf+hhViG5wPIp0lyUN3mx28t6X966j5SAZqDiUKjI3r3
4sOQkE7XbD+xUefKEuOlwyVv4Xf1bqdE2W7/WSWdw4oyRk8ctEBt+ZiWG63KUgn2
uZ/fGD4GVVGpGtC2aS4tisOrvLoUM+pdr7HmOfpWjq3YlIUjGxfzbW2K0tOzjFT4
cXl9tTVyzJmn58dAsHQa5DnMpUX+ut38kHwwa7XeQHjaE4eYVsZTRrM7nfuO0Qbh
MWiRHLDYhjF/hYTuuXcnlzpLkkY4RhZ3kaDRt8ZDwzgeli/J/FDSC2kYOjSICEFo
1rAKcOYuOsJU/SZF0hSxDRg7m3Q7gOcBWUNljm7tA3I+ZvGIJPz5VVmpfx0ips6O
5b00gym9nx79PEuIPxtQKi7clXjRJvFwDjuNstwOVeqbafqeqxCPMoYDShx2FFst
6xatX2ezwHRLkAZ0mS04gVK1QNny7mNdwAB0llFbI2DRb1ypn0cgt8TX++cH/4CH
LkrtGLKj+L77PetVm1FwRuvpFcwNUeWekK32hR5/Opzd5P//s5f2/sGbHDNk4baj
dRgL1N05S4F2l4AnLz0iQQozbCkhdYXUBbYTfD94Gr1qeDm6YdwiwTyorGz5nRgy
x0Jhd2Ls2CAzlBMN8pH0L8qiQXgHvxyHZsTuOPuF/lCAXocdtL3/6NLLw34aHn7l
jqw9WrZZdXZVcTsa/fbR6MfAqL6okib1R65KeftPU5dAYI151adbhbjXLYiaBfIy
NtYSiAa5Bc7TT9E7Vsn47pml6Z2iFfvOlUgih0XvCYkVFBDqGjtPu/OpHwSLRH7K
NJeDNE+lK8rI+e9RAJB4JgrnXJPOfBeitpJUMnxoZrb2/WVz8fAgJH959/rSYOO8
73oghrUfc1vHLuiuX3LJtTJl/r5OKHMy+oVbcwKuapneEpTBgky9pu4GKmYOQmiK
ux0qHxIUTjha2Br5uBQZg7RrAxqe8BkvXgk6J/44EJFHyCsdNReW3vph58fHm7JK
INPWDXH+dpDgcYpg8luxwY1mnzkXZlkbZ0lFKn0ZCQnjPruaKtsPgG+Qhv9bNa20
n3qZTo2XeLglk5jWFmwBlvWVXxvS1AeHceY2vEPYXLVLw3OJaLzczjg/kj0izz/f
yWy5SG46ecUkFJgCz38hOkN0zRvG3oI1PUaewRY7c9jTfsPSh7gqKhF3dl3bWbtt
fLwUITTHSDOzQG7pxYT8d6afeDIwNTwfi3f3P4otH+jxojJxgJCedacuwKEjn9Bf
0KBk0VPPHqFP8E6cK7gYvFYxITa8N7ikbfrI0udnPuZAdXPp35cf8y4fbhW/4X7M
21ETjnhhxh8CivprwkujLaYBmZVLB7o+3e2MAx/VPsFxMyAsRhhhw40GYqw1Q3BE
/MNybjxLQbO8WP7ygggMYIfDVbrHc7W5tN1L1yU/Da9S2p3ehkPg5HOOMh0BJHW7
oYL96m6pybhnDQ9MwIEBiMHM2PlEN3FmYg5509uUBPkvOOazvnNLK4HFgrVX9qY4
Zwhb5Irkrv2JEWA8aejY2w9NxHiJ7feJGKT2ErDLyudPLghlAcYHd+wghM83i0CZ
U4R1gK77EkPnvNlaQ9X+3tnnLFpvWqiK8CMJlxBD/MZPZJdZpQKHfrSP6Be2QyOH
FHcvhBjGV/rYxeYh5XnOrNvtUq6X0dW2hBi1wOta0FwBzl1od9yPVFS14Rqi2E5k
+Rr7856vc9FwPTlOXW+Rahlw1vuqGT2taGkKcaaK21jRs2+FG77sHyiExg7PkWlI
GIN3zlwhCRD37yeA4VPRm+Hv64cBIgrFuMfuVWDlv3um726g/67USrYT1I4yc05E
iBmy9PAjAoG4Stp2buMKuQc+zuf9Z7txncBFniu/NWKMwBnjIfizhoCrXN0CMaxC
NU9B8b94eRQnvIS6g/sNdvMoPlVguxpuTQ2yhclmNTsHrNcQ8+e6KMzTxBo2rNzb
JP6n5JQrqNURRHo/iaI5WQ/UeQpTFufZN3tY+AfdxekAUGUM7koJtR3NrmHamxEF
x+wbySmm6yuWrf69H26Lrc4DINDqdMcIxlYIXEU6nx8MdLot5wrjGAYULmJDnKSz
42vr3dfpIWNQ0Bo/uX6FoOCnijOpP74m/yMysY6QPWGWDjvvVHRbgzTksnNzDcZ7
2/g34VlTA0mIa2YsulXiHyVukSW9g8gPEcVWecKNNuX2ri/ISO4mDqbsi3ONG84y
5GZSRENWUPplWRvbMJB+vx1rIJwfbLt4BBx4n6SL+wdNULC4eUem+e8/ZyXIUbAP
fEGmAq1FunSQOcqP8mGAr/OoXxuBTo/XBaeH1lR5gVPSOawB703yvhBaRuEeIIqp
rbig2VAFqo3lvzl+bXJj24AcjnPQN+wVtcRlYH8g6gejmWGmnYIb9+m7HpP7cPQI
TBgRTzKzUkTBqzUYRg8VmFdss0U5hrIfU+NgoZzYE9DclHBmRaZKgeqIgn8LjY4Q
eyy2SryMZ251gonVqLFWQY4MW9CnO+3EtXSpP/VIXNFU7HdKXOMis1/jcVoXZ+69
kfJAiQYiTJ1WhInzVk0mCGXekb0vthAqW2RzrvDeFtl5r8nHfnxZUgMAgR6MjTOV
WVLoykqVgby6bI3RpzMJtx4/e141Z8CHhAo2zXzf4LjNV1RrzlmlnT3w7oMGxXK0
VTohEPvndwui4wsNp+QIc/uO21NzuMzs2/Vsey2KXX/b1fy7HKjOgJDxpfUyB2Mv
ZzeZBlPJZ8p4bllahON8IiLA93K679C1FimBNGzrrKEn/FoHAYbmrjlkeBifPQVM
GzRScgVSZNu7kAsNbzqwvABatAbGWa+jaVjDZghoFOO6q4j14RCWFT2bZeugR+dK
5HiBhnefmaLE+UPOUvtB0uI4v0UqbsRKNWrHmr/SRM2aqkARkz2fjGdwm3gbeQMM
Q/l19eRYDcoYAEaw7jDJhcK/UZ8YN90xans3LaE2+J75GgJugmPFiMdM7uvsHHxq
qNGiewUNdBzFDSdYWhgd70NtLsWd1XA3HQEh8shupItmDt6DfIU7DxnH41CnQ/SH
BvjLx2YuEqisL6lab1Af5PD5Q00k5QN+7gqsRviBodSX/fS0gYjyL341KjSKLdGc
GeXXdnXo+I6lxK68zWpxzD5PdtBKRtL9eHGKfJaE9wi+P1NM3gD9uHnbMaJ4YPyD
ueg0anm3wvPztuMsQ/4YcRSauAfRXC6MpSY1zI8mY6RGdALK7aDVK3nLWX61jD28
RRCVnjOASciCM0WGt8BN5W6V143wMNEzNrzKSvXHGGwAi0fhLQtsY2Di/C+vC8my
vYWoXH5eDJna2DsP8SKBIw3p8LXNY2OAHR9Z3zUZNfcyZSsBiKZ24/LVQqRodRaj
iosQgDkl6HnBzFyFgwlUA/TeUohEp1GxmE+At1KIycwLmkwLJbxKSxGOo2omhXZN
0C/mbQQxVeg1OWXyxzMqupUEd9E0rb7jlsGP7aamb65PPkP8bzO5gllC+1JUxApl
KeDqFqGLxvSCLDtyUKUwkumdgTkU9uRln1p3ouKNJZR2PnXGZ8zsLeBAGTPIveSA
DmRWrLHO0Odv08Fd+yoykTxMtRr+bqOreiGl9kRpKXMDGIKPBrKhAqBnGL7udKNr
z+YXOGUTloL/yvWk5wciaX2TWbR0TjG/w1UmhOh1t1adLqlNmA9EVHhfhrANRv7u
0BREnLTixK5XylWkoomGZr9IOq2xf0ht51mefbPe3wtSj4pXiTHKf13N1ONb8OPN
Njt/5Dw/4Fdp5vzSspyQ0XuEzcijQ+Ze6ly15Xi4VTe/0kL0af4QobJsAbTDydzo
YYHGaGxseLQU5LZeJDWXSao59sePzBdZUVmu6yNwN9diibiiDxt/n64J/kQwr95F
ySHltw3zIg7gM7KcqJiaLgaIW40WLCrpAx80QM95G2zlGUXFbVyAxjewgqX3Do+1
VpoN6hKLfDwLjKzhBNStJXc4ahS1Em+y3RzsKyeYciSqPAgMyJPfT4QSSpL2AXty
L714+18pacBP9M5bvwGXSJ2g2NbmiUxBmCZR0SRK5nQ7/SPJWHlHHa+/0BjS3L3Y
J7WVEBxF1G4Smc0VXzjaLrsQdspqQYbiaTX5NN35cRhPTC6pSzvFFSrvhQzrxXl0
lxvw3nfwkm1I5bs2CwIEZBXPn5dnE2ypkIMeoKHPUMhJrd47HsyqVPSr1KOkB5H9
AnNwIurdMidc8TwtpcfT8j/RbOn53eTEjUx3LOAGlGPWiEKAIvGcfzGhjcgB/B3c
hDLVPW4YSkGiRcDBLdMWa6Z2BsaVqV1i6edGJtdxOq57AfOBR2yvdcYtEEwOPpC2
ytg6CwPJPGPvaoSQmqgWEP1dRtJmXUeQZxB/izgzcH+H9e39SWsL2s7M1N26MkfH
FGuUaom9NTd1vTkxCQHENWCQDhKOP1ccKD/OdI5UVuW2V2wCpq+RqdgE19ZRrE7A
8Jicp6UhbVRDMYUkKpACF7uQ5STGUxL45NZ6d2PuXuH9G59FkOnm8PdDvibcRo6i
WMYuPMvIrulVScQoinS/mi3z6rzLQ9Mo/vTNQBJwQjT01ThnrbZZaxWtOiG1vBF8
FAFMLkqAQwoWp0Aunzx81nBpuD1Ygzv0LzJWvU+OD5qEUc+r7PP1p0oUt06rhlGK
udUH+Vn+ULJE2+PNqzrU0FtP4dbyNhfL9W/6/quXnQed801fJyKNiCYq1gUFe3VL
bOQ99NDvbIrqQWo5ZNitYg==
`protect END_PROTECTED
