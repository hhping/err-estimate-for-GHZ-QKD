`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfNF/MUsS4qIKD+7OV7JLWscFAHLAqZEA79i6zIyNeWJEdkG2ESDOzFP4MfPtdrC
nmEXg7kroPUHdMTwEWwSGy5ao59tFYyEvqmfHlvxT9o8qEDvpN0rSmwtW8kJT1kv
zDsdQTNVXUdEwgCzzjm+RT8zfWqijKEH+fgZ9yUyomRUec0D1IMWLz1DF7HfHuEL
ArOBfDNKQaDx3LLdlZpFwwPoosM2joElCN7KT+7BmiBjxuoeTxUFIPhBiAZL7Y+j
V26Zrd+mbj93L9WzHYWp6B0SYXD8YexoVKVSJiBOvEZb6mbQwoAEhe8wUgRgxnXj
L1Tuj1nwo5QRmcG2T14744rGdDfwoZNysg7DPZ7ytjIxYpgPsPI6a8BNs5Gyu7T5
FwXM7SH21Sju4ElChe2jxRB6dkU7Me1RFOF1vfT6aw4Irle5HyfeYQCGjy7vDgS+
7g7jNMAg7LfKO4l7WML6rn/ajmYtA7NLCdDpbCZUfxD8SpigJ2vDKgey7zC2i222
x4qjlZfc4md780EymlI6Wl5QRR3+1cKziiKXpmlTzkbBAfSuLadmam3WRmczRJPr
oy8GjsKcpfMscBVffd4CyHBaikQoTnYHVxCa1/st4Kcceqh4BJq2Pgn1e+YDkWTH
`protect END_PROTECTED
