`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Etdr1hRl6jysdK5HuA2LOXq8NEjKmE4n/FHppRto2GYaKLeTItPRaIQEN0Qvmiex
YO6jh7EbAQf59yW25OD/oEAXX0w/2PhNL0FFX1TOxmKPOqRkyab8B6MLMzwioV+w
L3yVBU76A4Va5GVjGfOjiXa58w3n7Vd8YXwt3C/N1AWhD/22SkhP6lZGsde7FU/H
/evCjW7D3fUJzTOSlEEcSEfy/h3JiVYqs5wjfwXlWn6mfe6bWyi/UQxCTHxFJggZ
`protect END_PROTECTED
