`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGLwYyRxoJgISEZ0fJHT0lc0CyOpqc8W89jv0h/hmzJhclczBwdt+/dgimidXiDs
/HBHirWXlF4TRbSOsnsqv055vog+5a5/GsKb8oEsyr/ZeLiklS1r6G5qIOokBtJP
8/b7DrlF/ZSF5UqsPik+VE6oezFRjObfDf/axY4N9KqXwJbObuVH/gAJzo1GsMA3
YB1ZgTZhnE+ZdaPqdmZCLYE1UIkGueJbIgYbWLJcHwe8F3CZaMnmLPJqxflxG0XC
8xlPG9tN0davnH4zsbITaFXF7pMBg2ps7LvZldk0jAaGlvjEYgPSheeQEgIsiTYx
lB5EelJccWQ1zd5h7mPjj01fTvzWGa8vgWHgU45IDIUL4TC7sR9xLYyw2GVd2cxj
NRdmszh2/mqrUFtDPaL5UdzaR2Y3nsZXHAi0K0oCi19zVD+58U9+zRk1kDoGYuzL
Ec6XUywaqMLwnNUQUnff2sSjuse7XwjvA7NQ8NaEoeBBcnUUhlYfQInAvmaOg296
AA8+mA4Ztav+jQpNzzn57aS17wwQ77TNMsKqmXP2hnBrQtLkteZ0quWEQblyyI1R
xGzEtkXyBV3D+epMUM2V0zjczPN3L//C6wqr45Em1G9AUqabDtlf6K4wMSLICVJO
yM3eVu3TD76oFUywGNppYdurY81UrctyRgH0ba+CguInhJf/a2QQvpR4bwlsGUS4
QQLoa+R9k+yOCn7+Rvv/6/bUqoDcfI0WJ4isnCxscVYQz69Gf592LUhbpPBWTNAt
GtO+f2JarWPCjbm0CkLqTqXj3xrTnu+MorKfkAODIlqNv0w69AasOIAU37FxghSC
9XmwtUIf9nBPGZuwPhG528Jmt9+5WMCmm77AEMJ/d6VwifhBiUkHPeKwZi1Bcl77
bV2hXI38THWQkNjZ7g6DXc+V8JOu3bVV/otTenznipPreVReOPSBaBowruQZMpb5
0Y0N0f3Kc6Bz4hFibZ1w87E3MkE5ssj3TNNPnLlyBSGTRSNbBC6Mh9S7wzg3KENK
nAyEfIguRF1V/d+xHdEECJ7kv0niVCXYxqVC0cmmujfdxgZDMIDF79FPnhtAsGX3
yO5EYSWhzqd4ALc5J0niIFCcqqBkZNrnIMctat66zKZR4f2dP5bmX8+OWYmP6X7L
ngDDytX5yKlvwdgJSmXY9y9kMHBbHujMcqUz2NjpEDjTARBDnurEnp+U3nMEOzFY
WA2+uh9uqszUKAfSzDc6BUGQw1h9Qu7Qoex5zYNDwSi6+D7UlhHzn8yuYBPNjPQS
PJ8NS3H+Ov4o1g+M7yhTa9MhkhWmzimWs34eq36vsgIMYYuQp6jhHC5U5zlacU4V
O1Qo+k0TnV7chdAWiMBtWD2C5aInTzdaFHFB2LgQTjtWQRQORQwy2Q+Y92Bhdqcs
0DVCpOUt2dgffY2cIHMSmD1blzP+gZ3UWZslG1sPSKYKfBRwST0xW3X55DNHR7kg
b4tAfoZmLv6NBR6ZL0qogb8w+oH1VKsW8Lk9U/ypUZHr9Ve98s7apKrnGFr9zJmU
siFX2WDHjjcxMDNUQb/yynAVFc+aBsamCfbldRspf4q8ebI2UcLi/DblETl811GC
qR/qkafhTnlMqzhuvEkKwDbM8JDHh5/4sm3JuCxOhN4gc6QwplRgd2mvKDYLD6Uj
BkbHAZ/UKJDIdGqQFjm5RQBioosBRgRun0aNvPDBmvPnHpucCrFF6YXtYvvtFTET
7jSTthLAaCM0ITM5mOIl3DSMwOo8hECgVy/tg/4kAH8fzYg4uJsVnIGC9k8fQojh
CtlCtbBTfEkB+k09xrOhlY4vz+aImFc0NoD9HLimSiBSGx8W2TK0WAtOydC10Q5M
VXeLbGF/N3XU8oYYvTrj5IbqYn6X7KGIKKBIA+77rU1RwA9+CLDgY0dF2YbMyDhq
bKdNXs/wi+1yGD0hiRvwgbFiWh/TsO0RfjyxjuQVoLT3bZWEik3f+rqwwaA19kqu
O9yk6rhNqWTMCDVX+j8z32uPlyszpU+HBapbQ1nsKup1G7iyN5cMHtNDTPtqApEb
e7PdQ69nCESS0ZXh1KPk4iHCx1ScakBEZmG2SKy98EksxpJG/ElwwR0h82gXAnaw
3ylPxDMoGidPY+M/HdCJcecyB+g7RnnC+dTChvfeeTynQfIHPv47Kfeb5oHAmSXW
nq4nDzxmgaqV5izpTGDTicaNnZ3vlyki7wRGnWH9b0kTM2sH7tczMEwDycUC8Ui8
onmUDHq1mLzUzmka8X1m9R0jhgnM+tXhiSynOMdCt8UaGicFf9S1VDWmNvZzYW0f
uEbp1SNOfGm4MQo50cAXUWiORcQXL8n3fAOpGIQE+bnk+FWoRJPBDkj2ET5EOb/v
JSDzWEKJmflAQ8iTbpxrv+xC2/foJBPYcOHFkmYoP0zZvBjiL29mEXjvsznHW5QJ
lo7fBdIAFD1HT/G/zg6z878DpaDFfpTWDUpveZxCF/h32mPm+M/MjU5aE0THNMn9
vL6GXPHI5y0JeMs6y+Ov6a6bYAMMt9Q1Ez/PWGfzLbfVPAPt5P+fxXWp9TrdZYIc
tL5e3u1M56Jw6iF+JZHyItbyitMimtqYiR7JtH7zDBRzZCokcbJh5Ci9jQUbvI0R
bN0dsnxxNLUHBoEU3BHKQ8Ssc3qSY0mDVjk6FR++mL1Ur/sN8mAhxtXT4MC3JxK1
mEmq1bTggk1eP3HbFnuQPx4ZQqnHE74KfEmFX8HIEBNZcWjzLLr6jiFV2eLKiikL
+iHpWcmdjghZ0YHE0FuSG9lQYmibGIUkv96HSIR+7lVNmOEbbghBagCwfKpJA/mA
aMUCawJG/pdEgbG1ff+Zg/l6iF2otcLUEAKafpbDgvhAWg910uj2BMexPcAY3UMh
NQw/HPyK7i+k/uqC+BRm+33/WDTXp/2ppL+9Xwv9pChIfMUBEjjvO6TVye8ZOheO
lFOLT98sLPudrJX/wO0YOOb63TjG4qJ3cpKfZ0r4qVI=
`protect END_PROTECTED
