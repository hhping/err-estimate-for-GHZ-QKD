`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2ZBoMTdQOP3zB0fF4fhb+vlgNqYZRmvBFTL8xs9FJaKfL9mfbqLaO043zzKKBDX
xNLSoKoWAuzfLS7C0hMfxHeryQJpo364KjS5btRACl+hUKCMEwxmvAPEFSf/O59E
qS5ND4xrd2bv+4TPFWZl1ybdrLBvLxLAIsKS69f6v9MUqD1Z5kjO279gV9g2OImY
aNacdWwXkXaTU92Rc35kfceBHm6Pq1VJOgcc61y6YET3BcQdS1d+EJpMGQVXjZTe
CJfvs/Yia9zzZfnJnMognNaX9lGLUgk9gZpYloqCBpbM1NrvXRE1p4HEQDSX2iQI
N2HJuEy3ykey2HrzxIBtUc8OHRq0XN6Kxxiyh0i/wOtkpU68zcSa/9gWNuDnAfmv
KelPYNajenigFADktAWPPZ0neefdRHejb+miX7N8WknYbmUWw2ucNBstp+dnYjg3
bQ6Dpi/gq/gqd/DLyY3KBkP0Wd2tyk+OiePrUR3h9q6bkKggaN61sGLXrUcFGQKW
Qy9uJji/o4HmPMyRx8USFiDZhsorz3iYGhNf1tpO4NQ8gLPasg9EQ9nRZbWm85nY
i9CbLmjmr/CFc8fSITbXKJDtv5TIun2mTIjeHQzRkA9RKCjcrOKF4sZAOx3WORIu
NDnr54aq+eiPTBYQeGIMemj7QPR4dzfHAKIIZy2KqxycNN/6IJe1ULlP2TVUzmQm
e87OUcT/j+EEwEpZkPukkKWdtEqSd20EWhujb3FaMH1hOZN9x2oo3TNmzeaRuNLk
j7Jt1KeWxq/qiDWG2wSp1jkKSvCDSuP7G8XyCAZrvyeJlLgsETf2OVLcCFncuyC3
/KaTGVl4GcxaSO4TCwWt1vd4GHqeoILp8I8WktSJfo+LSHQtc6KIo+8iDzi0w8BH
LIIo7yTCr/h+FfiG/lnzahH1+oUzKuxbHjLT27n+YhxCP74uuqer4cw2RUqajvLO
et0KMBrbWU8V+MItg8/DrnRflIjZ/3iUxQxIOl+sk8HcCBL5IzxY29T70BsGRD3s
ZdL/Nv31x36kbML5czaVzLcFztJfH85mxxt39KDwyVQrouzLQUd4pFrIckWdRpxh
Dax7BbKTZwhJa3iA6e4P9hhfV9GH3Wmh2dCPRH25UNyhed+qli2hwTXUpct9cXab
Yn99y2SYcN564O4WvZZxun6tX1gFfEBZGrSJURGC3PDJ/p4IFylTjm0MYgamG3KV
8VhbD7gTVfA/npL/A2JH8W5Rv8kCyc8Lwu/hmGWd3MdOz58dK5C3OzskksWGtL2b
8jBkEbEScmDCETarBFmvPl61IbyXTwJz/SDsiOcTtw5T5n0U9wC2AZkgb/Ccbttw
8NAiaAML6nt75K/KToYboCEZU1DbCTO+en01OPHYNQyti9y1z3D7wqHNhtGDC/B/
It6AWHa2lOSHyQg3oNTG/oJsa29pfudw7QagsWBlqkbGyqSxFgdAfEdkQf2UN6Tq
Bewlf09nPl2ljCJ0p7vlheFIY2v1G/0nCZ1JMSkPqgVYYe/Tk1Z+MxqDFVKL5jor
MAsBh5ID5Js7z0j2d9kN5nK57BblIwlCyR7SA3xKaxMHUYRY1UTQ81u2wT5vZ8VS
Fnb/YFzNmLKYrp9G4a870LoQJNI7m5ovYC2LCqdVBAZMRyhWpt4WT4z1kYvBhwZq
I/CwyzpDTk3c6MscLRIo7P5g9o/Pxjsn6RKaWwuOuKTTHbXO47kunzDfqjQU54sn
LgzGmvCtj5zm1fceVRT8iAObkCWpFVAfFbouVjoJ5NMmPja8Jff+w4NTfREt10ML
NveURRrxjd2LOASHSMhvdEASzqXNMeYfwsavSnT/oXX0A8jK6VHGr05ubRqO7S8L
oaSap87On0Xt51jrz/nVrwlCYUK1Nghn60htSjXUgPE0Q3URnc/gWmls++nrszQy
BReFppVgbmq/pBu7ZJWvdvPRZSaYRtX4/obJam/PY2AWX5DYfBtp5W2UcwxPUusW
qDqxiZQjNXxxFAzg9LvFxmguS//j0bI+GBQ6uG5LpFv/KIG6urhjLw9ZjouSkRT4
ZZS2QI1vP/t2Y3LMDGHuVzJiiLfB2aEpBJFsDKr/sP7lfGmxX5m+1/fI3JSZd5Di
YfCTygKFd0SVorg9Qtuw2HZJLnMp4SBa1xSgGOD1A/Whf55PQC2BwXVdn82CG55A
qhqFPd2TFRLz5SDFeb0ddmUitFlYuVk9RRBl53o/inSD6w1RJEU4XtDdDp2NR3TB
9jYCkTTjFLWIAb0jX+LdL3HOdqD1MXCVm39YzASVfsQB0MEJLj7/49oZvn1Dr/eN
R7OXaIhyqCFSU0zbFP0yh4GhExNNTkhOLDcyphjWmS1Rg0UYaaWdSicNzXgLoxFh
iXFZjxa+31VziuV3+UlYVCsRR6onULiFIfJcJPZXz3tQyIMvNo3/4SLLAC5LuAyb
qFYLUym7PLWjCYyWf9DIePJICM8luz0PFGpik6K3+4ze+k/ya+Tl5IiSNzw7BtwS
sKJTDD2bNTVK9SCGKMe4zR9qnp+3VAd9Xh/BYnjlgxkyCYyV0fGntbMCB0FRyC+k
AfWGs4low5iS7EckFpuU5m7kbtfCB3G4ODAYcKwJh2VnegyYSRiUQ1EFKU9QijJw
p0gNwqRicRjBGvgbHYJ2ntCGYiOuVd4K95wrcRhqFsbPm4X7nYOYVVzvvlAyP7qA
V8XnpSr0c6FljJTZOSCKKaIYjU8yn/VFepgM3DJXUKd1GrB/asuoDhFsnvNdvGvz
8kUKy+abuLWMGIJ2vO1YvrLhSB/kmGE+LXrhZkYeTwoft+hd2Sy5Juqa59cApURb
6+QyRiPgi+GLB8rnhS4Mdd/oEI0R/rxTGrozsVRx6IZHA07TaMMlFYaW+/hNWJFI
41fq3a3NXiTZNNfQcv+EtOr9sJoea18ss3Yq8DEb3CGSb5W0OAcbW/7ds9g5Ps6Q
vG1tn8fy1eDkp30eoViAux0FzPPvRv1nq6GtK0MrK9vCKK2f2qsvHgWEijfr2o9d
RkZe8IxsG1MQJ6NU0PQifBOrUTNKwGeUvAMBZ2ecufAcaasw9VnQdQw5FtYS2XvU
CpLeN2eV+YFqjVev5L9GgPikKD+QfhedYsia3lM3s9hEdW3t7TcRIgroeHsgclx3
LwLlvenYAmDg5GA0bA1tFX/tPl24YMK0lGcKC+teYekR44zeGUcuSUFdiOT0NhwG
arnR62FriXwhMBbFVIS22TzijMZQxG4nLFqXCPmz6wqwwZ5qCvugL6fysrHQIaCu
NEa9AwMBLyZAIwtk339BoY0fcmbaVfzPU5Yve5xx7LM=
`protect END_PROTECTED
