`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQmhJyHr3Zb0fHnr6qJUbToysSBIR0wEl4IR/GHSNxGSzmEpqJ5TsCgxPfYhRqvH
HO5h4Eu6eIF/XcHPbQ0yaaJ4CGCvHPJX2ljJ8zK7K6NJsc6h89YGNiSId3/wGMx3
VAeCOnfi5L7N3nn09t+KmQJ4lPPem3BVr9Fc1JBfBLV2Ui89Gr6813rJwYXpEmHn
w1C6BzJcYrV68G5+RPo06B4tm5BtT+/Ub1XX/MLbmsSYmb4UL70oC0zh7xeQsQUJ
XOTeTS1WRiwq6SFr1YZkoIub4ZawuIUwl90PfzQZfuira4+bHz7L4vnEWHMiAwN7
lLfZ02sMYyKQgK2KksULs6zLZGiTxTtp1dTwP0DZfRKBJPopT8MGzeFZ+HhMbul4
nZKVjnyAtmPbLLCsvi0Cqq8ZSHUMSQQaV3nfhAfwRUKn6Vs2ujYSWHbSLWA/kcVL
WondiBJ80o/sxsBV92g/y98ceqLLaYQAuukYN8lh9/De/PZWUMQz/a5jaizHuXc/
bPPsSmG2faPHk83WSHnWJrqSBDSXei64UkFsJqnYuMmG7zByfXV/Ah4TVqYe09Ag
iAFsp8LPXcq6XmoVC0z1aCUXGbBo/Bxs8QpA51gWm85F6dLWG2dla69kPbAFkfBs
T2EHhFPYfrnfrclKX3pCdbIL7wzI82flam2k7UDcg1GO7m6pJMpTJqw8BAA5PsVA
xPB5Zb+OaVx7kySGaZ0g7ktdYg4TK0BvSHUq4efp5BPR0IfdOXkBxVPXolGKrx7P
tn3LWlhKXJVEcMmZvsmZkFG/GMPAcbntSC3722o3bQ0EEnqNlWgPneVVDRXX1egb
DdFd6iSG6CsVGMTFGHYn0zZPOXrLnWQVjUxyzIwk/0OlS6C4Tt/xLfLNHIXsljED
2Iryt9/Tef2B2TO/er4sY++X+p20baw05epae2TRXd63DcfI3KIKcOt4G2c3GbHX
rRdle4d92caWkQGvz+WO/yvRgpidkvmDi5QVr0hljWeD7cw6rYhUObYZakL5AGif
FG3K08XFfC7H+0eSrH0Qtq3/wvbV0TuI0HJxddaJf57FaJU/AqfdC8UC3QhKK45V
RfGxG7oULsDnZTDwu96rwi+F6a29nW8hTEl9y1dZC3jzEsrUp8tbduiOrsKxNHrk
4BRUsSmX/DfasdKOg9SHMihZ55TnPUosXgELcIp4KKs=
`protect END_PROTECTED
