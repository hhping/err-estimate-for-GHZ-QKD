`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qk4nr0AUew3YQRtTleu1f0YtJiiFZYhujbI/GQpeWsMgDmcupmpciFh9We/oIvth
vhgXx60zJ7c/7ENNdknSsUHuq4M3t9SQlZfm0OrikijfJgiBpLhUFMJyQMMwAH69
J9XgCZem5GZcKTukvIKQalL5Wpz+YtZjykM95ksmQOahKx/E1TOjMuXXKO7KAqD1
S3mmqDkRw8DRJoIFgOjFpWII2n2H0AldEeJr8mk3E2j2itDvqxNMKV3rVO11M5jj
2GcJjfFywQzw+ZNnDl8wYaH7DsE4paHJyQ6I206zerx2r03EYWvOvp8KHKVi1v8L
QcmhLlXqFjbSvH/G7xhHDywiRyDJiAa5X2YVr8NXmm4=
`protect END_PROTECTED
