`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vesGlKrBf2ZaV0954LqM+xcEGhw3OOm+PtqG+O7TihLRyZIZ4ldrVTV+Hk4GrAwk
czLpCgYkgNXbgfLysZkmhT0lqPM7mheEftztDTpAbBpHAv8ahCHKOj077o5QIXDd
xyhU36gHpR0CWIzauQZOcaIUg/MRHhta2s4OQRVlWGgxFCgkFzS3kwt8pik6RxpN
pFEGbUsD6EvGWa2iMqc8SumIbuyLZBrHXpLiGzrwIt/sC12c6zyTK9TxiFW6sOao
8JxJ1pFrQnTp08rDo3UyDBWqojQ+Qhq3oTCg06CuuiBWCM3ANJQogYpB7QOfeKWx
R3Mz6GfpmG0fYM8CbLaI12lC9QyaI685iIKh2TqZ9yNvqTSFgAsBnKtJVk3eE8iI
jW20KCe05J/ppvPMXInpTkgIbkZwdmIDQEIaFpbXDT3fSvuUEouIVGyjUdaEXxE4
m8dzBv+aoOueGgSx/xT087jOK4SFLuIQ4057DIIyx31Uymvq+j1larnXsaK+o5z5
+0H1Mv4jhuRGeTBhz5DmYxPve1fYsfqeOtdV3YToCvnw5Ekez2knL50ZN2xoUSbs
bsIpQx2TF6bDODPSREQOK8x/OsweIdj8313m1tN7zPVCePGk2NYKtUDoqBdtnC3L
LTSB856ch9a/bpBr5qYdIkOdi1JKM/6IzhR1RQ5TnBTu2cZGK++7JvC2JczQ7URc
d59eQji/296wtrZgwctEum/YnzNK014qOc5UZLzkk//kivpWOBJS3daMSqFoWHyk
rVeM/tJRLVi6FYC7spq/2bup5eq34hhYZcCC6GR/lYsyDm1PXSGsuupRdS4Gpblu
iTcI2pXltoppDZDSutEfrwT0HmOlMgUY6OLGfz+pOnCE8gFfzn2V+IgNi2zWKMjV
AgfZjxW9juCcK/UByvlFsJNlESCnDOl2CG5TEo+uGVc8X06H0e0Wo9JA0hby1ZE8
aFxUyfWyW2S+wjDUSkXazNwQxc1pWGjKANLeq5F0mVBrAnIHLiXfRDf4sM2s0e8x
cDdj4UIMUgoc9LPzl1CONYbdgUt20TiosQ2vneV4pgmlgD1Iew2AdbABnC/FLVVL
kM+RJ24UyEf6CHmYzUyb9fHEp/BzECzo9lY5Wcf0UKjgcrV0vfGyT6Q8AQHeMXg8
9A5092ErqwbCaYgpnn7clF/a7yA/AOjiRHeuY24CiJbSlxVq1ZWpsgZC7cUfT7jE
Wjj5zriKimKQMOUA7E6Nxr8+ff4krC26PAdcSdLDxT9xKzcvLvbCj01FVG1Rx1jR
8e6WM8coH95omRSv38a8gQZe7Vlyuiuv5/CUqhEKYMeoGidw457V929CGzLuGUor
WCKeMzxNmusNO4I3hq0USFbqqP1inKgNFIYeyJH1kImAVC7dyAimAodHa5sZalau
tzuBID/VJg+voGz7r1e00c1tOmd36l8Jnx6v1H/Iv7+h+KbR1TBtVwQ67OFo7BSD
OJesHaUq6nP+ovFQdi3/s/VMAgbDOOXLv5PQIW1/MFPAjRPpot72RsvfeThtsaSw
Ua7NrbEfluKjKtxRMEWA73BwbQny2iMV+xYHN4jvsQ2l7GsDrhMZYT195FQCjZMv
Nt8Sm02WgJ8TpYtciT0wMbNol1sn4bFyIVQ5IoreMNa7EPSUE6KeRQDyreSYZVh/
qvaDbLN52q1zd6EcvXBDxJK01H1zmOfTwoPb8SToiyIDAHGDHyYPaO0/CYjon8+B
HuB8YB6p1e3hf5YYErJbI0Hdjd17oUpea37SmkMrfzYtZq6ANArqDmDmz01K+idb
qvl3huJJZNLr8zchwfM9Ghy083zez1pyyWmu5UdwNtxERhzkheCjB5mOoU+RRgLZ
QK6Hg6alqmDbQzWVFEdjubu5Cjybd/DMeF+5A3AmsAGZd0O11wGjr5IkWHWPzZV3
nP87azfAhSIHiykA4tqKeSEwdrbhibvWdz9V6iGlT7l3TuN2QV+qy8Y0x6uyA8Ra
6oAeVwBZ7eZr3i9VGyJKIz9Dbq5tnfiWXEWymbyZbh2x5br/VS1hKRq3nev2uBy6
i4vqv1vy27Yxa6tNIhdwJeLcy8umLzFROfFVB6/a0H4l4cBP5h6xqYgi6gqahvzT
piFyntQjkKtoRFziCV0PhPhHTQgyP6wGYVpbVtlbnrjq4GqXLIEYLjZ1HHeKsLmr
Rmlu5Ix8IiEMfLWIs3mLznAAWpxD5B4XdxcclofDx5DTzvhiwHuUb0+W7Lh0Ts2M
3U8uJ7C6TyolT1lkjqIT2OGmvWlZHcsRhwQDZsXq3RgC5c3coUq0fHqlEMuVsWbq
DYEZFlNv6JWcSrZYI+ae8NEXfNg/DHQIBn2JD5CTJqCEM8/re8MoDVtNYPaWEA8P
eNzzbSlVscvDt1kgSTZ9urPt8sJdnww9rxGTOJvHA5hjHkNqra4Vd2CuFN36Bqb+
e3AWDbuvUC7aKuEJCkdDl+tKLEzcv0i+tWp9Q3Om0z9/LAVN0VrJCfq8WrX+cC5P
Jy3fGp621uDOYiTQ42Xi+sYVQs5gGxOzKHDy2+mx9qj8h1W4z7kCgV42EED+xiwZ
F1mcBu04lAdDeHwgreFVXh1S/NsJISdkRaWwpGJLtPXVehoa3TIDjQsTac2TbyxQ
mpbl7j70RjzhnQgvzWeQu/eVPzhr857naPSFSmDBexOlJXPKFPWsHhJrjr2nv/5D
7jEEl7Vhvtph/qvLmI9rbi/BK087WCvdn64tuzY87hTYvqjIzPF2h9kdmlc26n5V
h1fYlNiip3jJ6mllWwuNLXlL0n62vu1oFvQ/9bIzT/qr4KSJDnFlP33aXs6VYvYk
jbx0q3eHLu8A97fjmMq5gpzef2zKjzo9A2OPIJcAKsgXRSPRl0++PZpbXZe9EmBC
NTGYDIlegRT2hqTqEoYjkhI+OkphBbHIYkOCWwV9kbovqBimzjBJiBMzmlXkfhK8
Ku+ZRA5whn44NcoIybZk0zV/HJBAJFDrOJ6wnuubyOCzoBZ+nZhzjbs7I05N5XkE
hf6IdSTnRNdP2zQvi/Hnt9rSLOpO54iNLy47nIJgrd+je6EUfQ4VziouuljcDhzi
dircuvKQWqFUMGoh3WiwKuKShm3oyrRMveat9/FfR9qY2HsTLqkijDOXuBo0CaVm
DEJOvkADndtc8j7A6JOmMdAmaB9A2VR6nduNTP+SWzuvZ9qHn+RbJddwAjHVvqi1
rIqbUlwXinx/bTGaF4PwUpIGF46uB6PwpXk4SeVLSwapo3RpUZlI98niOVmBlPlb
zeyn5UM/bBGe/qNlXh2oKErsl3a+P1O4mcRE2rsGHZaD069jXKDdxZaaYPDVwQnL
0b9oUujjD4lymnHD4Q/Bp0II1AtWUQTqgmhRbAFNQRdC7kDWptNlChPrz4yAj4hl
guu9WvxU7frAD9YyNDARIye0u66ThqQ2g5lOGiP6FxyNyVHbLlduCBSlGUP9qgUF
3pSSRVaul/OCFxTItibgaqppxsXeBO/CxXhAokYABU0kVrNNUs9dXPCTj1FJb7U2
5HjBx6yqdkjqhj/hWWMaTWfRGMoXb8HN3q37zbFhPjdoF7fSZOmhiFIP24e5NBlC
4pG//04/sp+DBAw5+fL0bBrEhBkjhGxm4fhsEELkDu8LS5njnYG4/WnvfcLNBSJ+
Jlb3ubYU0TazQLJ32fX+FeSmX2u+ccuds/k15A2rxoJhS3yejJNI026xbDx9/aPV
Eqo12PU8oxFtqBP1zQ205EpDCaYl1+s/fJpiD8tUMKQ1QjA6fEO3COXD3ng6ODWN
7ljCADPSJaOcwVuyHYjo+QOTsSIN+ERDd8uHBM79kPQqNaI8emcYfFatsDzvQ3RO
qL/O445/mLN7N3fdHyq+JzYtv6C3c6gkbCYceWciH2XCnOYM3NszGFbdV47C20el
xHJJ6a+wbXa2Io4fpkSfUnegKKneZ0BgqUu4btKlrpiPhd1wXGR/P+nPt6t+hs/Y
ktZFTIRxqUV+/rgpy+BKBwWkNEltBnsfmns4rkRT6YwCiU6NZPeHBA8jQzcssZKn
DT9R4mEeifETHpwMT7zy0yuVi66yNq42W69bq3Hz/gqRxAfmS2RUC61xD7G3duXl
Wq9x3NwIJ94HPt/Vyho+hx99rj58D5GGAgDrW2N4ebsNk+ISBNV5JAJwyWpIDnRx
x38HEtHl2ZVdBiWu3L1z6jk+AAJB61lk8p9YHEwZBOFUEU0aRdDlbilmIc/MDA0G
RYovfLvlTEKkAbid1LdYHbwhVaX27srU+VWh5sDqv84wGLuLB1unR5fB/vYVV8Cj
ASONtcMaiTWtPmgYgiecyvO761rTHgja5SzMLp0z9RGOZDYgn19EJBSoh+sykrBe
tnnTjRnLD8xLcE/HUv2VrHv6jI9mS5mCJolLMaBJI5F9jOsaAv98fF487XUzLz7Y
QJ9XICwYp31Kb7H/DKLxqlsyXdMStr48zRi2gkHLL2pqggxUdvfH3x7RdSThUSQM
AoisidhZX3yXuPKMk6oTcopo8JepwFzLUtMRN90gOfwsBV/TYuKwV41JuVqmmSay
HhEXsfSXBJwmxEWE7ZhrUfc3yW0mCiD2AK3bnj52I0K8XCt2TzIoSFXsgM4q6bIU
N9dCdNms8a5YvZvfSUJCmaFjlIbkW14VDsj+iq6B4xQnz1+eqeCEAZCYY5mtMRRD
H3qJDfgdiLXFzAMnttl/uuN6aAZh5YfR5m6sBDABX5mMWHIyIRLIrx52qCWpYKjQ
h+UR44bqBtRFo1NQP0Oe4mXclN+KVlgVZZHcugCb8JKGpUV7t4Rn27N25SIe6ToS
PC8sSL4A7zDtvyPn/S0vGK7oQWSqMhYIM4/fmXP9ZJdb6OyjWoGRiUJ2mpvEqPZE
R9pEpoMHzj6DAqq2FpIZisUqphIkiO6OYaXn/sqa8+P/T+sx9nCP3Hxo1rjuWHlg
ypLHKOM+2BHsw+QU8JHrmilysjZ+hGggidvYEsmh+NPGnQOg1M765RKAKoEuhL1y
GrCUTiVkQY7T/w5QhSNJQBvTda5NORva+I4xz+QLIOlTZzloQ+2rZjUmgtwtNsIh
Z0D48AaHxP7FnHYaQA1G0Lf0DkIWGjvm3+gR91cTCMdZGgS7V8tX8GrKkceRYtag
B5xEV+IvU/9dM634y3b6RbmCC7M6UJ8lCjTe8OqysAESbCQDshnzPdn5JiY1RcV3
KDA7BCrjeGmeqag9mpLE40vjsBtKpEwJ29Od7GHxRL8uR+GDRTsDbJ0y/bPliWrR
KPugONWulKf8i/OFg6C1evL7/gC/DgO9w+bDaQxsucEpWCNpjfZoM3aAoqo9tvZP
XMyHag3GAwAbffBNPJ/LAP7XWQpVLt8pd25ecxdvKDbOeCywZVCuMlY5EFKDip7+
XnilNT60pL7iiuhGxW7+mwIgQNtVgiCIgBqdd2xcrLs8OYl38RMAx5Aa4/OcCz+X
YFxybtjJkbBuC7oqOtG/+SEXiz/tfhhYrj3WP+mWpmv9eGhcsUSFoM1Iv9G/z5VP
RRnRM/+AiOPQUdK0U36desCxApzE7qj3o6jg2nN0iN/YDZjPpJ2IhsW4h32WDxbA
GEmXmkRkHCLoTvAL7/3TjdyC7rF7VxGpmXXgxkvbecJgC42WwLJWldxEpBN7j9G1
bezHwj7oeCE++hBvGNuMkyEmPGXSNCRuAsHlN2IRCAZJdevJcMloAaYDoYYobH/t
GOScmFGPt01SmrIkuWNuA0ICp7yD/aecPui1ccfi/qeTIYLp8DFzoijJ7DA8cUXB
kdfsFAl/O2GEmbPGPynR6Koo3G8BCu8NkE1vL8su1PI5hcroiInB91NnTx3czhNI
Ozl74mSd7e5D9An3ZuAin/PrnXaPr0YG86qDN7CoArTMGUshlRfouxn2RfvkntLs
2beqNEL0ICTWNYgZVJ72ybRpM0wOpVRf1FbxJyQB0EtNdgdLGgKQ4GeRTybtJ9U0
2HOgKtwAnW/uzErT1i4vMGU8r0qcPF4GbABXxOK2ZnTWCQw3vusCsUbvD4JdmZGT
iTGbMLse6oP3gGNQvg0xzTmf9J/yrHAm/wPdQw+Bg3YwmPY5R8PPWrn0E7hm+Nqf
y3bUg21xgKnouh+C7mmkq9NsSshNC2CBuuVCYzzYrI2zfLUN4FG2vNSfbv/NCG3B
BzQl0PmcNp0L0pL4YPUgqCEFWrdZfXrfSbO3IqpjHIqM8gyvxYTDNkOI1UGulXeY
mMwNwQk2+fp0VzUNe0EYwqnN4J8sXpjzHmQ59a8WbBXpdYSUC8ZeWDeV6rnYNMqO
s2CqKh+7+oCKCQMPH6tI/YFtW/85ZdO0I2nIDlE+ynxtcuyBohh2tfX3GAA+jNpA
wuOawCSbad4YcHwMWhn7qq+tCkWVSaqNH/YTgfz8ggZKclSqOHMjBiIbgNJcO8UO
SHYulXfuNir95QyXa0iLdfkqCDXOmCXc9gkunJ7XvRgfEq8RiFTvnl1Ff3HrUWId
YkurWn35YwqFsQ5X3GtJheyDisobEMAtDR3mlaHTiKO/BlDJmlO6yZ02pVh1TKW0
fQTBpaW4U6LFxqI2thVvgDoeI1DCNpKbTG3Stf1kykEjnMIs4Rf8FAScLdxBfVnK
ogilghXPWGs2c1aDC5WXpVRckhUMqHdv7gz1ToHo3s6eTrGtmX5qJ0qtLWUFNTTS
mAQRrmshVU9pSrQFu2JBz+lNdcJ09Xk95gvbW1uflpiVMUNOMSaTkIkFOvv5vFtv
N+EV+lNcoq/yMuJzqJvRBBuc7FJcoXy61C7RQypT50BUCI6kVMtvFjyrPuqVhfoH
GlcrNTMJ10Pq5NczbPOcG+RDE9IilWjNdjwiMcKZNNL4Txv6etKNmf+Dsl/YyXYJ
hIH+1rt18iU3S28HoS2ZlHJ8J8urEsLYvqVHo3UlyDvibLw+VdyyaMfGjAN4t4o9
1pQCjXj0AEJTv4ZbSUVz1m2RxUmdLPYYeDrIOUDyNkSsi9to/n7mP+rMTu4IHL+f
pfmztXQD8GHw328UqqBM512YwL9RrPN+xiiu+swQ0xOgT4kr/KE9Xjb4TS8KmO8f
b9zlXn3j3BvZuv+q3+4KGTZLpZHiAYIheF8et2ApJTw5CbIyDao6Qz2YaWW4zgMA
PtYPq4TRdYL0V2jKdCFjiDpVruZIclaz3yNqSqlLZJHMnlG8gOn8zGlP1MQNJtTN
D2We3QUlPTuYK5T1+Vfu9Xq3WHbu1LVY31BuFOgKTDv4BbowqAXynHadm7Jb0Iei
Mzw17fo22BeZp5vbWwgdGScLfoV+KgIKUL4knUDb3v2QeBVA6JTVf2P6V7ZQNBTC
qtFK2k49h9ndS+cOud8MKZP0QRUbySOmYVi/wwAB9GYCr8hPdrMYJn4U3eMccMn5
eT16a+D1+14siCvvgTc33cirdidfqDCnY+Rv2vzXz8FnIkbOZsudDJOvEFD4p4lr
2RSj8BBun154LfUQGhyav+QuAZHOUIUENoUuapgjwGCd70rKISbDCOkkfGBwZSa0
vC9NA7nWDR65lEZdB+CDYolpWpXbevw5aupF+qZZDeg3XX6OsYaivsihqQ2f++gb
XRQRQJla5tN7ZCHEg8dPmr5dGIHNRm4W3Yl1VINQzxjDpG9V5LIkfNS/i6za5qBN
5AeD5/bs514u2yww6LU0PHpzZegXV/wGYF8IHGdPzb21dOusMLTZmXhRDbgT8V0S
CE9NAZWmtHudGwjBsYPNfErir0PuZuGWEB/XwZxwEldOuGf3Xd0U1ihSc7kh/wWb
YEGTKswoXWKLq8xL7srOpUFYPoGG4tdm70tZEJJHs05DGYOKRBt9WHwKkz2FWH7t
z1cxuuT0OgLzuou/8xZ5lQCIfzKirpHjOfBZpcWzu0HfNmzTxEG0rf/koimp0M7I
brBlCoMbB5Ny+W0DFUzXZ1QhYNrS+aFFckJXrKxSdQk+kjQZSDRfmcumr7IQZNsy
/WGKGq1xXCkPQFmvdbaMVvcgRmP9IU/jimW2Tczi6Xb2V2KuFjwwR2l+L5DX3z6N
WwBE8K9j0GUtwJIg/T6c/rZQWwZSIv64kRnupYu+r6IllS/It/fCU8ZzV5NPRu1Q
+VfT5WexJKEElYTmUT1Og73SCmJdKw8VRKDw7CILjsJYN0QPqvInJqtwCCrPQBrL
sSwbYSaLdbGjV1NQ9wZndwGQzDASYBj0Lu5uJGmMJUDIPo4siA4HwNXJ5ZJcNUi7
XmtISjzbBMvRxML+SsYRoE2+lm8jaXTZIKB+triUWkGV5mIoS0xlCfwLPyiG77Mz
NUxLH6x/OscnNaMRLPENw/DDbTl5EiSG6vQVtm0q5JG/G49jGCRtaqT90FVto13w
gMNyHR3K/wQJb/k3PO9yA+ErdQ6y2yGix9W8ETS1/P5IrxoeMkBJznqHORf8J6KE
X5q+6Dm4RuJ/J1KGK5o3mNVKX9nPTHVO5HvQoqKQU1DZvq/0WE9uYmcytRSqGKra
LfTu7Uw4gw4/cJ/qd8nj2ymUHcB7PAl1akctJXk894kopYtM0URl14J59+JY7eRd
hplU9HlRacxRJkYS7DTlM29hhLSTFrnzAWvmagf21gtx9pppc9TIbJ70DY0cjo56
DUcsJwgIXsIR8xwFxQV1yt1XAmr2Qx7VjmS1D40wcH71J0JrUTogo7Psh3dkpxsQ
yWM6cbTBr+g7SpZQCsORPTaZ4P0U18NDxIO7B/KZ8HFNp53YbVlUfqJVw0vK2gTC
jw+lk3/upi5VdqjbjUYacvggpFX2mk6tLRrGX/qi/D66BTpzfp4U/qAOsxcxRC2L
y/mG2TZl5Ll1A2sQoyaDxPMUYLLhgsgcz+4LqYfWYnN0bxv62LGRPKVFe+iRwR/5
/AOhTc27FBZ2pc+pIcagh47B2jTrC72UjWQ0CPdc0aopDtOXk0rsfyE39Y/bgNTi
6UKsmSOy/RJVMNDSKDHVNy5MtTK73J852jWKumatuIFfa1fpLTJphxxUqP8bp/Iq
3mYS7sQqclAq55ZQBoitniwZk27E2V2rRz7l3rsmoM+TPbQkOqxluUD0msO/Unsq
vXja4hfb3IMRh8W51CSazKym4hsU6lAWNDRkAWMc/SkfJEZs9Zj1jxQk0n9ptWd9
3YONHebNd4VZ1wIULJeFdRk9gqEr2eukyUcyqHEdtc43zW+zBFO849xaS6Snizat
h2zoxto9RlFLq3lN2DyBwgRPoNBJJrVpqg9Zc9C2HxHh5QMPpbXQ+kvGi034QYWW
v9fAxHCoFoOgrqWe/ppMCUSl45kIkPzVApMUih+6ENUVT1zkibyI/yJ96CZggsUu
JoLj3DYZxtaDS7PID23gQsrFzXZ6OD3xANK9x0uQxFl8SNEpHJb/7YnZhaPSoLvs
8dEClQSVG5EjdrChyr69cW0ym9fE6EXaiAVrSKl2p6nsUURtrhLbtR4OtbS6GE0q
pslakLstVp4GVnD4pFM1HY0pphKaMWTbyETDgNaqJeq4ebHFbjMy4kYqr1NR7UvJ
RJwRgoxTP0qniiFgE8TkSiOiUvQzui6XUSOPBsehJ9iqz4Kwyq1zQqXoBTiw2H15
cFNHQQ8CuIZmbPNMJH1yxwwuqBSQbmXM/LeA/d9Cf28LRTuyiGQhf3VC2D5bzluR
sZ7WwOPcB1uE5VAv3hTsEbeaDZx9Nv9btsCb5JbdB48ccS3bnz7h9CMQGdLkAZVB
izlpyOQT0mC7bg2tdmcdlhwXlX1R44Uec5HmGILPTWzRsLxXlF4GA4aHRA2bGGS5
ZUuOsadlmWwmDqSNDnEFzGqB7ABVRDAJbQgYXZnRGuaRMxkmyUC7jvz55eCGfvW6
4qeuQ0b2BXSh3Dp2a17g+A+f+MCQPxclNKQXX5TOGeNKsvS3tX4Y0Xnf08uK4kAt
5wlKqKtqXy8mBbziSl/nSwvxaec84YJ4iNSUHcZV/0Cn2XpFLqMhgrSRZyFoBhkY
wIPrmnVJK3HOYsldVQXpcVZEq/RbTsW9fEgbGt721VPw7EFw8NNXgH4Mn3A5iJ8c
6mlmzuIx8Pk8p7doOCIB0YPLWP212t9LpO8YYdv0Ce8U9/0IyQAbkni/4gEnPd8F
4UQw0IWUWtw5pK0MuKInoSgCrzMu/SqHksyo1Tz9vHuHVdxsbuTtMxrME2VLt5Ha
gCwXG/fOIOiD5rxVQKq3lrMkrr4xFbHKURhh4XdhQl4gd0lCyNhlx+tWGnRITg49
gA29Wgt7huGKtMg8HeEifhBzvmif2tMOTRDXiJjpVc26T+ZvfGjgfopSroQBphwK
gGeQY9P7Lc7E1oh5vU/mR9tpocNm7NNrRmcxOsC10aHsSmlcrfs85goNi5Lvmx/H
ncgDdrM0bqlTjQSL9FAfykguhemJfdAXU6D0K5Fx1WkRyU9GlVqeCFeYWxMby2Yn
eQBSPwTnQIhK3yccmmyg2m/JyJgocS8XLbzEyKx1zI+2yMgohK6VcfCZ+kwUyTUe
+2p/dQq0vNEBZekPVrpUyH6XlKGFfKMlCyg3jGV27M0cqHSlzarkVQ1Ttjwp972o
cFvacWamEgLtNmPb+2VgaBapBJt3JNTs+lgkLpu/s3JHyQi50ozYWj9UCWZhyhW/
CpCtdecVbsjXZdwZOplr0gEm+yMbsTPxOF1DgkanqBrZAUB37NHmWFExkvdtAUWG
X+kj3sxIMIpk9KSZWyetntXW0ISmtkUZ7jtongzzEvvsemrakFwW+pRGHJOLn52h
YDI53pPkvt5R4+5u11L6AC0kUBuKXLv/9b2ZE5r0a2kQOreWDDrin1KCfEVwmikK
T1jYfAgl+9hHDyldzOvn+WCp/O0xf/seX0dqKQdkTvayBPI6laSrBWvlOt5WAYFn
yFc8+uu1aw2B1RDG0KtwC+TidA1oPZwbsIZS7IFErAWSoDJ3r95FINn3EsqT/90o
e+wDGV6r9QP8qolsJXHUQHRFxSfDFUvYm2zY+PvZZtVbn6tSiUei32/qU/YUD/he
gRtTmiDO6uZUO/5NnMFpAIIyfQQhx6CGqSSurG5s4776lf+1EbkRDC38J3EApOIc
ECUAYu3MunJUSaRBjm2ZYXyjtcCdhkObdpuwz2pK0vypSNtNWeZInWO3ODwp0fKs
vpOEszmPodZhfTllMRMp3A3KUpUSNjFGSlRXJB5LFn5m8O3WOMOyz7CGHyiUgirN
bzT5+aY7WVp3mG6DZPp1emAfJIDKR78SZ20lSKNMkjyblP5POEFPPQMpy2PCId+j
n2yIUBkQYX010kryL16qjk7RbIGOwGI4j8lUmaaTk9ndYev1fJHiFVZVZFlgk0qp
W4/9xD7jxj/alJp/5lg4NbxhxEbd/n71jBfumEBxxvUfqhugeCeCAsBKXnCH5jrD
C2i9kYCY++5/cEYOF/dMMWuwLBJ6mwVcrb8TnIhEb904jOT/UXOEBVhjtyApe5qu
dJG+orbEXUy26fmUayH28SJZHmcx1SjKDZJnyw79IqEmsCK0/+aO5CKnwdNfHu/U
1+Ey8NH4UtcH47K4tETdndrK0yBiJa4iAo2u9RSivOcCDa9rmn3jtgYl7SWo5DBp
/GB9kJ5hQ21ZBaMrWjv9OvjzeXHQBPkZzzaJN+gkzySxtAanZoW3npPVtaYXT8o/
`protect END_PROTECTED
