`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WU9U+isUhqhbHyeHCmpKRuVA3+eIoKqcHkNarYLn+bEVnwhRlEaWDGFbFq3Tu+ok
HyxoS8KvjUdw0WdR4Dy0hY+5wp5QVycOnVPHT5NNNnn60nrXp5S7ZSm/zlu2dhBS
vBbVOHusXBZtlIECr4Yxdb/IkgB9h9Z1bfpctsDP1o1rBUoGGsqZsph1ehvqBnyg
qwPMeDFuXPRb8IJ2fKR0h5+IROhiPPPj+46OfmN+pBMeQySZRfmVEdpp32YHYI59
cn7MDmzNYsTvbjjPFFpbyjp6QmXC2IR5Lpu/zzRl/eRF85JqduhaGTi0T0mXBx0P
RZF0Xen88WYet1AQXM9jjTdIO5dnsuUkxLm5VSRtNhxp09mxqTm2B8TxiLIYUkHn
z4Ey72+dGZX8ObL7MJHC0Son9x3B2vCMZcUy5mtY85h8KH2Nipw2Iv768lC61io4
k6pWIE5J+j1wTZabBr8Uj+Dm/kG/luMbDK8m8fM9ua6oAaHVL8n6JAA6lW3+ocze
s+/1g7yGvkbKQrjYL585DaErmHeFh3IrFP4E5lwCVpy7Ip53AEheBR4txypk56ww
J7ShBfPyoDmZsKtE7YexPv2HXGfufpqafKgjVLQf2iXEZKRgxf4406pTvk1LIFfF
qskfDHWGZZWkXJ0Lk+IfWzRZq0/L8w5VR/EGuHBpAVFyYI1Rdjsf99IZcf/OGOQA
8KBUigH6V7jvukmy2wM4UaJBcpybm1vwYwgVHqB7yNCXSHQVyZeLdRlvngELRoyb
pwcsIohVI3h8Ol3XLqfgVGli1Zyyksymo3QOGkom7xygyTB2Hv79nxJVrZdd6UQR
xcdCEvC8V75Ecqf14OTCCL87NoRdlSmlvAVtuHYjKVGB+mIcTW13wNg9dhcereBx
c7CFHANfGkR0JDxUN8ozSDFtANSyDTUA/fMWUzVueVwCJ/KQKoVMwfZUx0i42sAf
zZUmUIqjQTdsJNO4q5mBF8U3pEs+Q2+GR+qZXv4952kbPosUETnwOU/7Phu1BRZk
zZt7Jr+miSwa/9aeFgl6yY5iNJ4Hvtn8KhMa6E6zFNw6R+mPAAID1Y8n6Mh3zo48
pTix3ICvyCl0LozbkWy8mhw373SUemkQf8YgV4v9AuBmiWdV5zj70j04HR6IZ3hZ
ZiLDOMmZGJzrZB3BD9AMDV0ulE9ZWUK61pXJveQMLV++g+U3DVie6t7oVR8KuBQ4
dJ/emEy1e9rhlKLpFllM0TdRqMbdTMMO2o511XCTyCUv2rw43dxzJ//msJvlXlqC
s1TFJeRADnijHivALfuIrBrXhmv9QCeJpcOg6Ah3UgiYxttu0U7rouDF6XbHxzl8
/xZE7wDf07jCUckAxYcyB8BU6Hq/VPL8sCDn9hLYPnUtmNBS+tB4Iz0yJUr7verA
IhpIApxH7W09Iw8SDrRLeSsZC7IWmZ9ibkVrzryBlwBx5AvTp0inghEjqj4o6XWo
KJekEAfHx0S/O2e50unDrM0p8Pr1+E16oLJMGg+Ed9hOBb60XOvHj38wWwsA5WOJ
Ea01pNmapiEoo8avM+RcomqeTO2TyyEJhuyhoyrwxC4abvK2aG8LGZcn61v6Txjo
lT6Yc53N3zq+Gh9DqXdvzzTCgEarZcqCNUM/F1/el/8TGD/DkQQEJkfAH0fe1bS8
6429tiPr9Lsy/N5Bcq43x8nUbsqT1TgGzNFbgHuCmqJfhHLRs58AF7xjlsfn8Qte
pfqtKYqrW7pc3pfcZZiqeBXHpKO51tUP/cEEZ0zjMw8wdCmt/CPDtkf71pl940er
IgANPm8sg39JJxx5WgdcfzutRn+sH+RdNeZNJr4C7NcRei72oKj7cKHzFebTd+ep
3B3+cXYRk6sMtaOmPBMIOVBz9vecGg8PK1/AUdZpktC3DkvnpoIeKineNymhY5op
pvQQV9wyWigYI/fVV5ZeyjZOBgmCc7sIRCpAlvSwrH/xCcJtKO6KLTiwuCB64uUk
cQLYVJNCJrEEtiNt/JTKCuTMrmTebq8UI4Ipj/+nfVMy94JdM4VyuC8t2Gl6ZHCK
rAfofpYjn5VKTY4VZ6GmQgcdofpN56ku8xQgiD+GlVJw7i6sBTRaVvvRzAYwpSWJ
NwKDm+vPB8O15a5mBPcCyYW3i9obRDVxlC0jevtXeujK4EJ2OLNGOrI8lEonb2Bj
O20DrOhS9o1QgGC3WWnJLjnGp6En2EhpJPDAjrmTSnSMrwbjiTqDed3InQv8Dtgu
EGZGRZhwQYgXgejaEING5HkRPEHRRjXi3055Fje7V0ZcrsjevmuafXnJSczAVDsM
tR5lhSGgEvNzxvjjfmn6bPJ6blYuhZyXtLzs6UmGw4XWUtcIvfc4QNuT8l/SxlEu
2Vy7fSLFs8sGp2swWbWZD/EJkL+W/kV9t6vFSv0tktGM5p+mhG036BiIcfq9SLOk
3BsJBrrntmfXmV3A1MJU+PphRLEg17QjQwlIOrUaBwCqsEQh3uNUAr53IPNPnID6
b1Zoui51WtHUIwI3exVkng1NUs0mfVsonHlBPgxwnWd5x1bj/z4/5NlkRDTpSeWJ
Onv7H5aA+Eny8zbLq+yZMrPHZTM8so7Nlmre6S8vzFKm5+RDEKYpo5dZUvaTklnn
3JpDkjFJa166Ht5qS3Aj1xeaj5K31wQAtH0BtT22NPe077Xr6IQnT55Ya+LTwWQM
zSBs8M74XN9jfPBsOF+Ja2OjINqXer7xKGkNZgCugxvjvWmEkBt2Q79w7iSfN6ky
gjfpyapJ5RySI1iyc2Frii4vwh2Z9igCxtGERFoAaBSD9Gv4f4F8mIeKZ2Tst1BU
16xG7IYliB9kHfAkBXGsk3pg+aImKuihq7H57j7nTO3Tj5EPv2bVRJMbFwFeyDr3
+rEVQpSeXv9Ox2M8wI34s5YAJF2TqZSBT5GnzBgQY6+F7JuTSKNjJRKVkpgadko2
ngoL5jbxCJ6NyGmTNZ7lF19o9T2AlJsPHJM3WgYI/mDdiOnpp7M0DtUVYWFtylbh
5Cb8QoMkNoqOzJ77RKoXyKgw7xSAJrP2BV/dTw4lSpuE6FFGqOTDwxxc7GziOu0p
xEQWhapMLKvo6oc/iJvzRA==
`protect END_PROTECTED
