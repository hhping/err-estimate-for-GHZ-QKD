`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQKywfIbfQEByXHqHjSDlGliF/AIOMLPZ1rJ/C2yilHnL1uW3uCFTYee2LNh/tDU
cWcZ5j4rN+zzNF4nWQT2oyiEjUdStXe2C7vqF1UjoiZKnrKKzXwVQIyG9galhXwx
vSFFVQqK7cQyE2FA7MIxO++rUurge7w3ikjUt1cam9gVF8GO6KanTzpHgfPfZ5X3
D5bWPBMKhm4ErArKrvppsNLmujIRJqznQiWTU/UKeZuftAH2PaikCT/XaChQZRzP
LolgyrS1fOOl8SQHdTBLVKDZawzddo9XBx4o6+9G0G7PlAOxResEjlQ73vX9dT5o
E1VL6sZ9lkWXbtbZoIPy3xR/3JJqi0kuhUMm7072qj+w3AlPqguydKvKgVibn60L
V9kdD9YmAqqI67CrYJOFBnu83qdYsoj/oaSFaS3446PDZ9/BHQTfyRqLsg/6fieM
/PxOe1jg3sgHF+Sk0CewE8TYgVihVgtHmPDQyi/kI9Xl4yMUJ4kF2sx4ifusqey8
LkblnPj1fp5raIFVtjJRRiC4yKZpiSgEfMd8CyC180yvlzB8ggZQ6tD6/zX7QZgE
zFHIYG5k4q5ks18uDLubG1xJynTJmmluHIVtxTxnlOg=
`protect END_PROTECTED
