`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEIYWApjGKBGJVgDL3XTOKeeG845QRsgFig1w9x63KBXF8qFt4ZRzpoOSDSjgjNp
6bY8jz8x1v5KCjfRXmGcIo/+UKPjp0F/WwH0+Zarfl2SdAZiN1rudYWVAN7LFZE9
O9YTvH9se39tTcmt7lQrSTHG8dN13/w5uRqg6Pg3jIlkjm8ZWQW6aOWjrFGLS2ES
pu6ahpkBn5XbD3A+9Ob/oDltFElvDmgr2CqOxzz174BA8ocUgsi/K39HRd6sGDzI
Y55UoHxW56mKKtgAMbfWq+vZfrzz6hZwcM8ZcpK1U4u0TBiLdwEsqbIsiWSXIpVb
XNqtLZjm4j4kS27HJ0Ao/fw6QHHs8bzsQYCD7e0SgaEZKUqrNNoi83Rl7eFZeAd8
3dFPwCIo2HLQuENFtdUwJdgLk/MLqLvJqp0bYG8sfVtXKPGzalT00LdGNWOyZvH0
qkIs3py8+r2X9wdWh010Tpf9iuqcwCHEtFPRM2y0ZTEYRr776TP52lVdL4t6oWgF
HJSx5s+5iKQ8gV1b+24TaFlSAWAEDBopYDfBW1jFWR52FKxUPntCLoMb4rwlpCoo
dwlrHmw+YKfZkn9xzIKAlck/+ht2Mqj7pdeBCmJ1HiZrti6UFGxXEcW6AY0xLFZ7
Jhm2IXh56sdwYeAEg26TynjagoHaXwXB6QJysicBDTdrn/UIRY9CZ9xe5heLgFKu
1Hl7yk8p8065/qwg7I7GVJd9KtKU6CZamVEI9VbWqktapaWsVBCkKGjq4LvW83tP
pSZKFk47B/DnjCSqQo93BP9RGfJK3BLb8AUB7m98EXkejNVBa26JPO3765LS2x3V
tji576s6cVwNp5DpYmsyp2nSCdnbnegHHor9tCrjw39OK1OhL0gmytqFk3qwSPFA
FSuQ7lBheyHQHQcukGyNLjFxUIn2/2n1TLpnNOEOZpU+ALUTpQPUPVy6gG555oMT
cJApo8QbncZKrQHOwQa/wcs9Ry/vdlyn2BpLCVZwi3UgFqGk9JtZiGP6gIPf5UFy
1T3EOruY8xenMuyDJf8JSgax0ZmUl/E2C22o8zIysCBevfEkID7GLllROjZCUTW2
Iehg+4VhrBHTOruhlEX4HD3LZp9dhdwdt/CBuM+vLmfKoxVir4yg4LwbUDMFbwfz
cm4Wsfk6hVczyXPPDq1/LXPyGXC9xt/qIHSGpCZV8LcyGe0X3IVpmB+w/2J8zZxq
ol15RAnXMadb8lI74LFRjagTi1GSEHlLtJhdLStvkPZxuCHDT23sfUkAKGSaf+mE
yBLiYJDm0Bbb0dgmi8dQ8jpy2MP/ya/cwHgwetiPPoUIxMPISgA52u5+zKjMmEIu
OMfMxjevTn85MXCVuNC9kapxEVuyAC9WjwlSxL+V/xHdMshM8Misucjlxi8W9VXk
IPbzpCx1Kk99KndBgRrD8EHG09ljBe6Ij8XrYUL233C6+SvpVZQOP9bCGjPmAzWj
93Rfb4kmI/Q9XIdhPjlXhWrqlu4a0UR6I1bbBzj10+oVi08t/8znvw938FNy+jXO
NlRG5NAC/350pPZ+/WGZLbvnImX0TAyXZ0nRFbjh3iH2i0kdI77oc5Ndyz2wiP8k
XHP/BBy9QHDhhvQUEDt7vFXUNSDEPLNRm0ojqyQgpX8t7KYDsfPJx4C5UKkKGCZx
c5WlN78ySmREVMiQ3gRiBYCmmU77esjy3P2+axrENvPW2RRA8qlTIHCErmKsXL3N
7xw5pmmnWOgRGRF42iAHcKgPDMXgD8cLrG47Y2K4zWl/8ojEmCn35jneK978TQsb
OIEv7Ss7kqHxHACxnEjbrMGyhm+oSQykD1ywUmqu3OwkF0wkbqV3HTgS10WrukPP
ZMlxOYu+AHQtPqrLWHaXXfub7PCestcn8Xf6ebIT6dQETF8bRr0oMWdbuEthbvr/
BQIm7PQR1RyS9pbrwHc0YGEQxAguymlmWAryhI1Q1JHzRqEcX69Oa63Dr0XmAbVX
hg3VjtvNmsPpRjFPKTMpdZrzCRm3jScV5ZNR4RRfqtKoOGygNR6w7Dh0wmhLDIHr
SxvFq26+tj/834GmtJ4CN0EyTdDfyQB59H2vnqoPBCeT5+5K+xDDj+wZ3Yq8NZCp
PMm+yy4K7hWAHVYoXV5jbQRVsgK1qzjDZFxn+yvz6yDIKz7DGcDMMbdVcGCSoucF
FdnaZXl3nkNm5V2Jt7kFyHW4tRKAExQwHYsF5iySfRkejJOJwy8SYiY401k5raeR
pvmeK2GNM1n3IDAKslvDsFJZM43cGEAustROkK9cEXgHwY5LEBw0b5MYGaL12gGu
jYxz0VIVItUx3UUO1snYLa5T8tYRqMfcn0xaszu+ktDQUOHpkiGAli2q3XzvmDLO
ujZgBb+PdZr4aZp0o4BxcZxZt2y0hRLfGsUNl7HtSbyTEslj70VtNklnC9YE8Vc6
g7qS1Dmb3s/0oOYkSAy0IiLus8z23cQEJoL/wQqZ+aWryl77RnzW3iVPncpfvnJf
U8aejY+KJ1JAvOVqmE5qrFf+PWa0o8QWVIfibnRPf1Y6f20hNjgyRuMFc+rITPIN
N+oh3FANHOFjyfDlZpivFVAAKybS25goDR0zHe2bvcmR/yn6TCpU3NfTU63QoRB5
ntLwewrV3kdwsjpG2+fFZZrJcuzxf/gCtyrLwTdWXciz4oqDohF/JLwY2L2Q4FBv
KluHtTWNx1qWw3DqTNs1CFCW5iKBqbJoTBpNnS4OYj5DCIS+zlMEVKU5v5m3sjLN
oi0UJaG9LNLHPmWPQbXyDNZRI8wcnOkek+7ltU/PuyLqjw2axazY/rXnYAZQhkHN
dtIWl9gabpAWu1MZ7KU/ZzaKtqtxaB/1RySVAh8Cr3KToClp/FjempXxO4XdRNSg
VFDszSz1Lz4d7vmEws/Xmwff58mYvLoaLrf1K1pEn/TH01wQoXyIYCHYy4B0fxOO
YQ3j8UUlacwVSpowEZ/WdI0eWc2GloXH/0I2sNYQ0Jc=
`protect END_PROTECTED
