`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Seoe7/h47s8OChf4tCmdfVnt/wK0dTMpfXPKu/MgrGPXvEt7NqIdFTsnOl8xN3vb
To5QbTFvck5G88Al6/aZ4ruZHivGZy3YaFsiU1ATmjEdmSVhrKExi1xtfrloPgN2
sfORuiYxBmrpZrRsyj8OZTyw29QETfOOVt+00VuKI9EPoin9DaA+Qpw+2QdDzNN0
Cnvp70r33ftZfzvSq+ZBp8IM3DDuruSnIKNdM8/A8yAiAsha1mvYKN7mWiGgZ/oK
roAJac4NVpwIEHxW1hUIZpN71snByYz3bZ4p1sVaBsWypdLV0J3Axb7JtVSd6tuC
80ZpwpyGmrQSDJuzJ/on8j6QqUiyYjWDKfm5i/TF0Hr71k0ZYBAhIWCToCxZi0Fr
zHqFklCstZL1tz3LpZU5zlg36gzhIz1mh+g87c7RQM29xlxv1S+xTRLD3WfaruzL
fyfmqwsvaY7uhDU3TXxHl6MJJgRNLq75BGEFHQNSQKngL0i4nyl5D0ZINInNjZe+
4FQcubIVPHEb6YolcDnOHtasPxuvTfMciBicTPDDcdrDMhNpkqoIDraDMSbXcImu
q3GZ/AOE3wNq+C+SBZQ+DikNROyXD0GAoOWsMfxrWeX0SCah2omAOBHqKUiftnXn
5nyJbHs/VsOKYd2I4DwOztsXCHWEL63AXHlVRv6k9B1Q6umUx6iDC2gx9waQ1EqA
z7GiFdqQQENHw6TZwjlVPKZYAj/i5jedRJiA5BskD8X4zMatvF5+ZtoExRJSRL56
1ODsO5nHjQtjF4JECFszqVonZv4ruax60AOn3DgiiZjq3ktMTTG5A67czPv6ApiF
XR1OHyCDZF0vZGbpW/n8QVZ3iP3uyiieyFLMgoQCGTfyzQobFTR0GTlcZHHFsE8p
UfdzezPxuEvyAV1+0x0vLe4eQUXKc22spduKJCs2KPhPH6Yebavc9Py0r/IkRxAP
IyJ6pqJVc72QRHly39np+5UJAUR9T/sLxf+xWPJ1cDUPwpblFBgbxA2CUMYCaPL7
CzefHPhuJpnh3+cHXfoQgu3k9Pi+b21oCffGY38oNpp2SiWEzB7urf3wnWK/fKV2
SvcKoNar5PCb/U/znP/vzBmyRNMj4hYice5qE3PuSDSgSvrcctY0rFHUidF1ddiq
2D5TyT80UsyXKB4eL84lA4jjzfmgkUwhmvWTRkgJMAcWDXoVOGKBb7b4x6MfF18i
t6PyWSDpDgoRhm0LOS1xvM1Oyb8lcHpO5rFABrajciYbdvrkWlAnJHBu0gC76pCj
kD0sBr//U2tlqIUSHmdkX/y1ex7EiCcPp5AFzeNGmQ6vWRZEISKGiX2Rj51LTVmn
8sXPmgAvvGqBRhFK4ovh6nMI/S7WC4RIFnfujhpp09N7BSKazbIYPV64s93587g+
CA2VA5/5ZC9oZpwY+I7j4km8GGCsmWENiJlysGjBN6YrqMR4O6Zf0j40euLaWp/r
ycMCVewjYTCCmEVVE8DS2wtWQhJVUkdLaz69r9yeE2Mxke4K44h41UFIXsZVTYvQ
TieW15SKm+lZ43RDUEofUSg9dbsz1ExIVFdt/nNZ7kGVLTVY0RjVUZftOgQr7EhW
87ET8hujnuEx2zgQeztrpPEA8yIYfV08RGz5DS0egxraHE65Fdn410RSn5ekrxG/
XChK/GxqOebXwa7RlTITKndn0/rok8iw9W3pjpNnGgi9SyMWhipZtpLzgHRCvjOE
5OR68puCRm3XRWR4cwDOK/LMJ7z0ZCl3nNnEkmBN4kA=
`protect END_PROTECTED
