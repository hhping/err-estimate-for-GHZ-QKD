`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZKa3da8X/Ts+8WGXO4mwBM8m9YTzDCORz0wahPCotfchxEsdQlMruSr005eFlAR
3/xo+iecdn5lqILLfy/ZVqlJziOcESEOWT64c1522P6NB7dtMb8/OsyIU9vA7RjT
joy4XxD+BDVhCK7bJQZXVVfwUsh8L5lyUxFEwXa6m35NwOXho9vdJZTiIhQNxPRe
xlCro6vvvqrfcIEnGIk/o8FTlDQg1U8lpcJFnPa19XLGxASjmGAEGrEe47tbrw9n
n6v3fly4VfrRW4RQkamyx1fiwzHeZzj5YB18Z64kdjkYulxzkSiHqc7bojYrj6Lh
Ukswxf+Vpe4B9feQB6Aj04K+QJgwUUzFKCyYbjMGU63iKZPcfSx9xn3+QBgBajGC
4uQVrEqWEhVESOhs8mOkxcvA7QKH7QtcTA3ko9u0Ls4LFQ1mSr9eMLRPCETBVD9k
sVJbPDePuwo8/sqU2+P0v+25lGccXH20/g0q2QztqX/c8on5hb0BjQiP3ILIMcJw
m+a1R8NRghJnB2uGhXSK6OHNjbf0RkpoHreZBxuubdRcqLsqID655BrpzM/25Tno
6csgkVYtl6q0AHb/tSDi4vhk5O0os0ol978CQ+2xP/87yRQx9J4GUeQYQo6gTy8M
3rg9P+zfr2nPMiWSekwMW7B7KUZdbJKQRnB5V/OXFmD3xgWFIjek7zKB9aucrLOU
RH5e0NSws1ktXJRIG/EK0xoHRl21l2SXaZfByfgTEyJtsMphMMWHfTC8ORSYUSCl
nCZRO+JH8SQlr26mjatzUP5rBqgOtvhg+v1nQS12daiK+/SQeOT16Vk+/msSDKfU
rw0ydW3QRyJb5jMMRsW2ZYQNWs32myzQX18d9FDYpeOrN9ku3dTH5cm5wQ0uWQYE
uFRZg4pSmeBqEOqKxeGmCessncB+2e1NYkpxA48uF2A/VIohizDpOZIws7ZImMDw
agT/3pN82uoj4Ko79qi7Nn1MSpk/qY93uOGmQLLsekV5thqKgdBR7w/r998TEvxF
xkbql49u+vGK40+mPeXHR1otDvnq7fq1zruKBGzhr8qOjcEHzOQrQ9GsQXdAWFge
nzUraOWSTkhK+JiCdBV7HXOdU8cJK4SOsN+VL1oyzmPRNIv6m3ZJRrBtMaTtldZH
YNbev9c31jcoDodQKX/MELQALaS98dYGi+rmrFfA/GllScK1Zd8hkOtJ0ijHIiax
/VS/d+XN0cGUDvvSCo/l3ND0aDQQFXVFbashu+9T2vkP0r6R6P00fZK+9Jwennln
IRiqqq/5ZXvJ+CwsPKr6wg6kqwOn6KMxWjPyCqOIOp1LZhz8Xg+5wb1P0BCTS7ES
cR30/AFPnC35cApTCriNWWAL+jvl9V7Rc8vwR121AGwneMBLlNnmwh3/9rVYZkTy
G9odxu0WEKTvBB1ZNNzmEfnDR+eevpm8k0sZ6soSijTNJ1zX0Ms+97kMAx2t1uZg
4z4n1Tb1vApiFyNS786KP8WsfcCj0TH0+3C1kaVsIRSYlDnjUB1XGblMB+2WSPPW
H2vy80cySU3hEydB9eji5N90pGnjoVI/7fPJTqy66EYfog9I3nEP4+DQDA29MMwD
g9dNmLYwiXwPSlqdpLL9XAXxFx7WWSQHw2dHqPWztnfAGwAd/cQYNZRjksl0qv6N
MqVNIFGXtG/D+qmoDL1DccZfvibLxVzLYL/crinQf8eJ5ke03r5wL/AebHhdi9xE
Haz0vFJ+8wEyAsKDyX+C+IWMbp6wXIrWFfD0wjWaRkQQTW2fsDEPPdbbUAeJhSkq
DImLqwW2t8xDTyxou5mynLZ8ezuEs6SnRqeZKTAjh9UjreK4WzDl15xKgnfD5gD8
3zePkUlVC1COM6c8bjf/nkD5LMcmav8Z4z45Oc/hshRbfAWbvRWnWW4mVLa9bxfV
HApswf5Q/02nMqFRnaK7yENCgAUA0GaI2iijlHufjxAjVX04pyz6XPs78PZ5eLTJ
2pzRNSkgIaa4f4Fqxpx8as1QThf3AvZaNwHelIIupSuVkvnchrwTjn1zAm7dVyYR
YnxC05CZqnB5ii9ASVHxf6HUPx9CrbK6/NqOAF42pmkoviagM0qBbyMTmJsPNvZq
gWTZ6aRm8Et9X4uQaT2gwHI1+sdk2zPSECAsYonThu2Mi+j54jCBd1zeyVZtye29
GKCX3FNX1CAQuB4pwjey3wI40KfKmQNT9knmno5xzAWM5cGt/tdIiFEL+hgB3xpP
OValExjxAuLbjjDFPXoTFw==
`protect END_PROTECTED
