`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiZLlDvhZ6WuEIYYiortRyyYs+GT0mEhzYNGljuBa9I7p+rCRcx7XMDlEVXEpGD1
WNuWv1aOQA75Ok/LV2gubMx1t8nkXYbo10Q2XEgMHCED0K46a8zZWZNOwn/pce8X
RBDfRrbitP4dRyNoP8ypoeykA6Ulg6BjkmtpKoXVSnguU8aad1X3oe96GbzRHuYo
pFo2wHtNt6r+rbzMHVQSMIZ7dV+qEiJMXOZ4yJKHzMujj3vy25SHDJh9vxYkJvWE
+cO/50pHLNjUv8QOnebTFQzFt3hrlH18iZf8wI66YyUavtC4JpKIHHzj2PrU8IDK
dnyksIBUeKbQbL6W7yOgoLFG0uWX0RQzANOjau9taTYAF6eDzM5Z88Gb9VrtBMWP
+zBa03duLdtaobS/WzfeYwmBsyDfcocTCO/3Xy5+vvL4BZO9nONnc6sfflchWa16
oYySjbdJ4BFvI5nXrF6Bzosb36RV9HomJUIIQO6qqDU/jaP8oQt8FoGqJtYa+4fi
ZFHOUdRE5GwvHc3vOxi0gO/7zLIqzEKYunQAQk9ycLU=
`protect END_PROTECTED
