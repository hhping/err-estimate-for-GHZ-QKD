`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fo/yxEFo0Qa/8vQZiLwJ2FlTe4MNu15fcWvVjy7YDbvSSDelhtXU4AerHyX0SyDn
1b+qjpzgrTotryHr3erv7QTlFJZwAlVZy6VK8Viy8nnuy36In1PkSQ0kaSUoaLfj
FW2ldLiNPd68reibTOypWmdUtzETgsiOo4ZWQ/tay8nw8rosXhv/ryb4WVmT7qpy
qt0X/x7Cl8/6Q25srMqM7LKiVTXwZeKqbYmEgwTGZ+oPrVlEkpraSor/gpLmFXgO
K5KEFiSvpu4nyKvnt2F5M/3FW1Wr9RJX+n02IBZu7hdPGX3Ibkm0TExDsFSpYNWM
vAPIhlO+uEo2TFxzBxkxRRRB7fcMjPwbNP/s9VTjNZ/4Bnx7I/kPqoduvAq+2AcZ
BpkbewDTBxbJ6P38JTXpgRh2KNMFX5OpSzXATX2Z9cR22j3QWRQPrmq6j5bIv/RL
t2OA7vMxVsyirHAplxvGogi0R2vCgU589Y587UtaPq2iLvRGvppCTl7LtSgA6KLD
t4DGGplz0T07JKKuiXsiqr/goI+LnAgdgSv+axrUF8ipTSuRcMDQIu/vuMNGQol+
S7cGMPR5T0sUXoD1uYdURPv7cHcIiNQifJL92ayB2cgobyKT34DnwX53yLUI0aru
VBaimvxrs0hqGCmD49N/wxbIpaaJgPF2sJkM1drXO8tDZ5JPq5tnWOMmnJCleBCi
oYN5Xe7ijChuogHxYDMyLreeFtL2VKg8KBngPlRF3vCRBsmqjslIefarZUpVwBt9
1P8OEmrOd1XiGDmynesbOg==
`protect END_PROTECTED
