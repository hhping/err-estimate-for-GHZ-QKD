library verilog;
use verilog.vl_types.all;
entity twentynm_iopll is
    generic(
        reference_clock_frequency: string  := "";
        vco_frequency   : string  := "";
        output_clock_frequency_0: string  := "";
        output_clock_frequency_1: string  := "";
        output_clock_frequency_2: string  := "";
        output_clock_frequency_3: string  := "";
        output_clock_frequency_4: string  := "";
        output_clock_frequency_5: string  := "";
        output_clock_frequency_6: string  := "";
        output_clock_frequency_7: string  := "";
        output_clock_frequency_8: string  := "";
        duty_cycle_0    : integer := 50;
        duty_cycle_1    : integer := 50;
        duty_cycle_2    : integer := 50;
        duty_cycle_3    : integer := 50;
        duty_cycle_4    : integer := 50;
        duty_cycle_5    : integer := 50;
        duty_cycle_6    : integer := 50;
        duty_cycle_7    : integer := 50;
        duty_cycle_8    : integer := 50;
        phase_shift_0   : string  := "0 ps";
        phase_shift_1   : string  := "0 ps";
        phase_shift_2   : string  := "0 ps";
        phase_shift_3   : string  := "0 ps";
        phase_shift_4   : string  := "0 ps";
        phase_shift_5   : string  := "0 ps";
        phase_shift_6   : string  := "0 ps";
        phase_shift_7   : string  := "0 ps";
        phase_shift_8   : string  := "0 ps";
        compensation_mode: string  := "normal";
        bw_sel          : string  := "auto";
        silicon_rev     : string  := "reve";
        speed_grade     : string  := "2";
        use_default_base_address: string  := "true";
        user_base_address: integer := 0;
        is_cascaded_pll : string  := "false";
        pll_atb         : string  := "atb_selectdisable";
        pll_auto_clk_sw_en: string  := "false";
        pll_bwctrl      : string  := "pll_bw_res_setting4";
        pll_c0_extclk_dllout_en: string  := "false";
        pll_c0_out_en   : string  := "false";
        pll_c1_extclk_dllout_en: string  := "false";
        pll_c1_out_en   : string  := "false";
        pll_c2_extclk_dllout_en: string  := "false";
        pll_c2_out_en   : string  := "false";
        pll_c3_extclk_dllout_en: string  := "false";
        pll_c3_out_en   : string  := "false";
        pll_c4_out_en   : string  := "false";
        pll_c5_out_en   : string  := "false";
        pll_c6_out_en   : string  := "false";
        pll_c7_out_en   : string  := "false";
        pll_c8_out_en   : string  := "false";
        pll_c_counter_0_bypass_en: string  := "false";
        pll_c_counter_0_coarse_dly: string  := "0 ps";
        pll_c_counter_0_even_duty_en: string  := "false";
        pll_c_counter_0_fine_dly: string  := "0 ps";
        pll_c_counter_0_high: integer := 256;
        pll_c_counter_0_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_0_low: integer := 256;
        pll_c_counter_0_ph_mux_prst: integer := 0;
        pll_c_counter_0_prst: integer := 1;
        pll_c_counter_1_bypass_en: string  := "false";
        pll_c_counter_1_coarse_dly: string  := "0 ps";
        pll_c_counter_1_even_duty_en: string  := "false";
        pll_c_counter_1_fine_dly: string  := "0 ps";
        pll_c_counter_1_high: integer := 256;
        pll_c_counter_1_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_1_low: integer := 256;
        pll_c_counter_1_ph_mux_prst: integer := 0;
        pll_c_counter_1_prst: integer := 1;
        pll_c_counter_2_bypass_en: string  := "false";
        pll_c_counter_2_coarse_dly: string  := "0 ps";
        pll_c_counter_2_even_duty_en: string  := "false";
        pll_c_counter_2_fine_dly: string  := "0 ps";
        pll_c_counter_2_high: integer := 256;
        pll_c_counter_2_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_2_low: integer := 256;
        pll_c_counter_2_ph_mux_prst: integer := 0;
        pll_c_counter_2_prst: integer := 1;
        pll_c_counter_3_bypass_en: string  := "false";
        pll_c_counter_3_coarse_dly: string  := "0 ps";
        pll_c_counter_3_even_duty_en: string  := "false";
        pll_c_counter_3_fine_dly: string  := "0 ps";
        pll_c_counter_3_high: integer := 256;
        pll_c_counter_3_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_3_low: integer := 256;
        pll_c_counter_3_ph_mux_prst: integer := 0;
        pll_c_counter_3_prst: integer := 1;
        pll_c_counter_4_bypass_en: string  := "false";
        pll_c_counter_4_coarse_dly: string  := "0 ps";
        pll_c_counter_4_even_duty_en: string  := "false";
        pll_c_counter_4_fine_dly: string  := "0 ps";
        pll_c_counter_4_high: integer := 256;
        pll_c_counter_4_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_4_low: integer := 256;
        pll_c_counter_4_ph_mux_prst: integer := 0;
        pll_c_counter_4_prst: integer := 1;
        pll_c_counter_5_bypass_en: string  := "false";
        pll_c_counter_5_coarse_dly: string  := "0 ps";
        pll_c_counter_5_even_duty_en: string  := "false";
        pll_c_counter_5_fine_dly: string  := "0 ps";
        pll_c_counter_5_high: integer := 256;
        pll_c_counter_5_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_5_low: integer := 256;
        pll_c_counter_5_ph_mux_prst: integer := 0;
        pll_c_counter_5_prst: integer := 1;
        pll_c_counter_6_bypass_en: string  := "false";
        pll_c_counter_6_coarse_dly: string  := "0 ps";
        pll_c_counter_6_even_duty_en: string  := "false";
        pll_c_counter_6_fine_dly: string  := "0 ps";
        pll_c_counter_6_high: integer := 256;
        pll_c_counter_6_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_6_low: integer := 256;
        pll_c_counter_6_ph_mux_prst: integer := 0;
        pll_c_counter_6_prst: integer := 1;
        pll_c_counter_7_bypass_en: string  := "false";
        pll_c_counter_7_coarse_dly: string  := "0 ps";
        pll_c_counter_7_even_duty_en: string  := "false";
        pll_c_counter_7_fine_dly: string  := "0 ps";
        pll_c_counter_7_high: integer := 256;
        pll_c_counter_7_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_7_low: integer := 256;
        pll_c_counter_7_ph_mux_prst: integer := 0;
        pll_c_counter_7_prst: integer := 1;
        pll_c_counter_8_bypass_en: string  := "false";
        pll_c_counter_8_coarse_dly: string  := "0 ps";
        pll_c_counter_8_even_duty_en: string  := "false";
        pll_c_counter_8_fine_dly: string  := "0 ps";
        pll_c_counter_8_high: integer := 256;
        pll_c_counter_8_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_c_counter_8_low: integer := 256;
        pll_c_counter_8_ph_mux_prst: integer := 0;
        pll_c_counter_8_prst: integer := 1;
        pll_clk_loss_edge: string  := "pll_clk_loss_both_edges";
        pll_clk_loss_sw_en: string  := "false";
        pll_clk_sw_dly  : string  := "0 ps";
        pll_clkin_0_src : string  := "pll_clkin_0_src_refclkin";
        pll_clkin_1_src : string  := "pll_clkin_1_src_refclkin";
        pll_cmp_buf_dly : string  := "0 ps";
        pll_coarse_dly_0: string  := "0 ps";
        pll_coarse_dly_1: string  := "0 ps";
        pll_coarse_dly_2: string  := "0 ps";
        pll_coarse_dly_3: string  := "0 ps";
        pll_cp_compensation: string  := "true";
        pll_cp_current_setting: string  := "pll_cp_setting0";
        pll_ctrl_override_setting: string  := "false";
        pll_dft_plniotri_override: string  := "false";
        pll_dft_ppmclk  : string  := "c_cnt_out";
        pll_dll_src     : string  := "pll_dll_src_vss";
        pll_dly_0_enable: string  := "false";
        pll_dly_1_enable: string  := "false";
        pll_dly_2_enable: string  := "false";
        pll_dly_3_enable: string  := "false";
        pll_enable      : string  := "false";
        pll_extclk_0_cnt_src: string  := "pll_extclk_cnt_src_vss";
        pll_extclk_0_enable: string  := "false";
        pll_extclk_0_invert: string  := "false";
        pll_extclk_1_cnt_src: string  := "pll_extclk_cnt_src_vss";
        pll_extclk_1_enable: string  := "false";
        pll_extclk_1_invert: string  := "false";
        pll_fbclk_mux_1 : string  := "pll_fbclk_mux_1_glb";
        pll_fbclk_mux_2 : string  := "pll_fbclk_mux_2_fb_1";
        pll_fine_dly_0  : string  := "0 ps";
        pll_fine_dly_1  : string  := "0 ps";
        pll_fine_dly_2  : string  := "0 ps";
        pll_fine_dly_3  : string  := "0 ps";
        pll_lock_fltr_cfg: integer := 25;
        pll_lock_fltr_test: string  := "pll_lock_fltr_nrm";
        pll_m_counter_bypass_en: string  := "true";
        pll_m_counter_coarse_dly: string  := "0 ps";
        pll_m_counter_even_duty_en: string  := "false";
        pll_m_counter_fine_dly: string  := "0 ps";
        pll_m_counter_high: integer := 256;
        pll_m_counter_in_src: string  := "c_m_cnt_in_src_test_clk";
        pll_m_counter_low: integer := 256;
        pll_m_counter_ph_mux_prst: integer := 0;
        pll_m_counter_prst: integer := 1;
        pll_manu_clk_sw_en: string  := "false";
        pll_n_counter_bypass_en: string  := "true";
        pll_n_counter_coarse_dly: string  := "0 ps";
        pll_n_counter_fine_dly: string  := "0 ps";
        pll_n_counter_high: integer := 256;
        pll_n_counter_low: integer := 256;
        pll_n_counter_odd_div_duty_en: string  := "false";
        pll_nreset_invert: string  := "false";
        pll_phyfb_mux   : string  := "m_cnt_phmux_out";
        pll_powerdown_mode: string  := "true";
        pll_ref_buf_dly : string  := "0 ps";
        pll_ripplecap_ctrl: string  := "pll_ripplecap_setting0";
        pll_self_reset  : string  := "false";
        pll_sw_refclk_src: string  := "pll_sw_refclk_src_clk_0";
        pll_tclk_mux_en : string  := "false";
        pll_tclk_sel    : string  := "pll_tclk_m_src";
        pll_test_enable : string  := "false";
        pll_testdn_enable: string  := "false";
        pll_testup_enable: string  := "false";
        pll_unlock_fltr_cfg: integer := 2;
        pll_dft_vco_ph0_en: string  := "false";
        pll_dft_vco_ph1_en: string  := "false";
        pll_dft_vco_ph2_en: string  := "false";
        pll_dft_vco_ph3_en: string  := "false";
        pll_dft_vco_ph4_en: string  := "false";
        pll_dft_vco_ph5_en: string  := "false";
        pll_dft_vco_ph6_en: string  := "false";
        pll_dft_vco_ph7_en: string  := "false";
        pll_vccr_pd_en  : string  := "false";
        pll_vco_ph0_en  : string  := "false";
        pll_vco_ph1_en  : string  := "false";
        pll_vco_ph2_en  : string  := "false";
        pll_vco_ph3_en  : string  := "false";
        pll_vco_ph4_en  : string  := "false";
        pll_vco_ph5_en  : string  := "false";
        pll_vco_ph6_en  : string  := "false";
        pll_vco_ph7_en  : string  := "false";
        pll_dprio_base_addr: integer := 0;
        pll_dprio_broadcast_en: string  := "true";
        pll_dprio_cvp_inter_sel: string  := "true";
        pll_dprio_force_inter_sel: string  := "true";
        pll_dprio_power_iso_en: string  := "true";
        pll_vreg_0p9v1_vreg_cal_en: string  := "false";
        pll_vreg_0p9v0_vreg_cal_en: string  := "false";
        pll_vreg_0p9v1_vccdreg_cal: string  := "vccdreg_nominal";
        pll_vreg_0p9v0_vccdreg_cal: string  := "vccdreg_nominal";
        clock_name_0    : string  := "";
        clock_name_1    : string  := "";
        clock_name_2    : string  := "";
        clock_name_3    : string  := "";
        clock_name_4    : string  := "";
        clock_name_5    : string  := "";
        clock_name_6    : string  := "";
        clock_name_7    : string  := "";
        clock_name_8    : string  := "";
        clock_name_global_0: string  := "false";
        clock_name_global_1: string  := "false";
        clock_name_global_2: string  := "false";
        clock_name_global_3: string  := "false";
        clock_name_global_4: string  := "false";
        clock_name_global_5: string  := "false";
        clock_name_global_6: string  := "false";
        clock_name_global_7: string  := "false";
        clock_name_global_8: string  := "false"
    );
    port(
        clken           : in     vl_logic_vector(1 downto 0);
        cnt_sel         : in     vl_logic_vector(3 downto 0);
        core_refclk     : in     vl_logic;
        csr_clk         : in     vl_logic;
        csr_en          : in     vl_logic;
        csr_in          : in     vl_logic;
        dprio_address   : in     vl_logic_vector(8 downto 0);
        dprio_clk       : in     vl_logic;
        dprio_rst_n     : in     vl_logic;
        dps_rst_n       : in     vl_logic;
        extswitch       : in     vl_logic;
        fbclk_in        : in     vl_logic;
        fblvds_in       : in     vl_logic;
        mdio_dis        : in     vl_logic;
        num_phase_shifts: in     vl_logic_vector(2 downto 0);
        pfden           : in     vl_logic;
        phase_en        : in     vl_logic;
        pipeline_global_en_n: in     vl_logic;
        pll_cascade_in  : in     vl_logic;
        pma_csr_test_dis: in     vl_logic;
        read            : in     vl_logic;
        refclk          : in     vl_logic_vector(3 downto 0);
        rst_n           : in     vl_logic;
        scan_mode_n     : in     vl_logic;
        scan_shift_n    : in     vl_logic;
        up_dn           : in     vl_logic;
        user_mode       : in     vl_logic;
        write           : in     vl_logic;
        writedata       : in     vl_logic_vector(7 downto 0);
        zdb_in          : in     vl_logic;
        block_select    : out    vl_logic;
        clk0_bad        : out    vl_logic;
        clk1_bad        : out    vl_logic;
        clksel          : out    vl_logic;
        csr_out         : out    vl_logic;
        dll_output      : out    vl_logic;
        extclk_dft      : out    vl_logic_vector(1 downto 0);
        extclk_output   : out    vl_logic_vector(1 downto 0);
        fbclk_out       : out    vl_logic;
        fblvds_out      : out    vl_logic;
        lf_reset        : out    vl_logic;
        loaden          : out    vl_logic_vector(1 downto 0);
        lock            : out    vl_logic;
        lvds_clk        : out    vl_logic_vector(1 downto 0);
        outclk          : out    vl_logic_vector(8 downto 0);
        phase_done      : out    vl_logic;
        pll_pd          : out    vl_logic;
        pll_cascade_out : out    vl_logic;
        readdata        : out    vl_logic_vector(7 downto 0);
        vcop_en         : out    vl_logic;
        vcoph           : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of reference_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of vco_frequency : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_0 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_1 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_2 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_3 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_4 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_5 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_6 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_7 : constant is 1;
    attribute mti_svvh_generic_type of output_clock_frequency_8 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_0 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_1 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_2 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_3 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_4 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_5 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_6 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_7 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_8 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_0 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_1 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_2 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_3 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_4 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_5 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_6 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_7 : constant is 1;
    attribute mti_svvh_generic_type of phase_shift_8 : constant is 1;
    attribute mti_svvh_generic_type of compensation_mode : constant is 1;
    attribute mti_svvh_generic_type of bw_sel : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of speed_grade : constant is 1;
    attribute mti_svvh_generic_type of use_default_base_address : constant is 1;
    attribute mti_svvh_generic_type of user_base_address : constant is 1;
    attribute mti_svvh_generic_type of is_cascaded_pll : constant is 1;
    attribute mti_svvh_generic_type of pll_atb : constant is 1;
    attribute mti_svvh_generic_type of pll_auto_clk_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_bwctrl : constant is 1;
    attribute mti_svvh_generic_type of pll_c0_extclk_dllout_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c0_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c1_extclk_dllout_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c1_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c2_extclk_dllout_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c2_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c3_extclk_dllout_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c3_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c4_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c5_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c6_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c7_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c8_out_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_0_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_1_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_2_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_3_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_4_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_5_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_6_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_7_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_high : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_low : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_c_counter_8_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_loss_edge : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_loss_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_clk_sw_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_0_src : constant is 1;
    attribute mti_svvh_generic_type of pll_clkin_1_src : constant is 1;
    attribute mti_svvh_generic_type of pll_cmp_buf_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_coarse_dly_0 : constant is 1;
    attribute mti_svvh_generic_type of pll_coarse_dly_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_coarse_dly_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_coarse_dly_3 : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_compensation : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_current_setting : constant is 1;
    attribute mti_svvh_generic_type of pll_ctrl_override_setting : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_plniotri_override : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_ppmclk : constant is 1;
    attribute mti_svvh_generic_type of pll_dll_src : constant is 1;
    attribute mti_svvh_generic_type of pll_dly_0_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_dly_1_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_dly_2_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_dly_3_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_0_cnt_src : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_0_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_0_invert : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_1_cnt_src : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_1_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_extclk_1_invert : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_fine_dly_0 : constant is 1;
    attribute mti_svvh_generic_type of pll_fine_dly_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_fine_dly_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_fine_dly_3 : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_test : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_even_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_high : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_low : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_m_counter_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_manu_clk_sw_en : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_high : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_low : constant is 1;
    attribute mti_svvh_generic_type of pll_n_counter_odd_div_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_nreset_invert : constant is 1;
    attribute mti_svvh_generic_type of pll_phyfb_mux : constant is 1;
    attribute mti_svvh_generic_type of pll_powerdown_mode : constant is 1;
    attribute mti_svvh_generic_type of pll_ref_buf_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_ripplecap_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pll_self_reset : constant is 1;
    attribute mti_svvh_generic_type of pll_sw_refclk_src : constant is 1;
    attribute mti_svvh_generic_type of pll_tclk_mux_en : constant is 1;
    attribute mti_svvh_generic_type of pll_tclk_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_test_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_testdn_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_testup_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_unlock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph0_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph1_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph2_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph3_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph4_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph5_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph6_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dft_vco_ph7_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vccr_pd_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph0_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph1_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph2_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph3_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph4_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph5_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph6_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph7_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_base_addr : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_broadcast_en : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_cvp_inter_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_force_inter_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_dprio_power_iso_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vreg_0p9v1_vreg_cal_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vreg_0p9v0_vreg_cal_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vreg_0p9v1_vccdreg_cal : constant is 1;
    attribute mti_svvh_generic_type of pll_vreg_0p9v0_vccdreg_cal : constant is 1;
    attribute mti_svvh_generic_type of clock_name_0 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_1 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_2 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_3 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_4 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_5 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_6 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_7 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_8 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_0 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_1 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_2 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_3 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_4 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_5 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_6 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_7 : constant is 1;
    attribute mti_svvh_generic_type of clock_name_global_8 : constant is 1;
end twentynm_iopll;
