`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yr4aILUAGCTE11hbkGcU6QBVsftcXTUzsWW30bgg/rC+NM8r1T3zC8YVSa5J7WL
Bwrz1JZrZ5sXWmqMpOIWdHdWFLQxZnMlGX+TaGhen9i9A+F+J7geLgRukRepaXo+
pqB4uVxQFvUjLMHIn4OmZPY1I8UF4DKO+k7ksLOUWnl/XY1C8l9SjHP5rk1IJPhZ
zVTtTggB5aOO4isGGRTw3gboxfsL4/GRsHoQeqnW7SyB1ez2Pvg79a6MEB5d/hyw
nk4szCMTsP2ejqCE0FibQDbrBf00LpnCNGeM3zxfsYzJu9Jfdx+BvgZk+W7AgzPd
bsZQaw+u/JOBfBBF3XuUKvBr//4ojzvs4L4AEL5vvGKYj6uxPzgGIkH5teMEFreY
Pjw+Jks4c2aiZeGe+yzy5kUd21XuSD1tPA4SploARjPoEMPzWhw56E63bX+uv0PM
ooUKk1o/02t3K8WCQfnhpPQ7Hr/6mvENB6NjMhGIK0aJ95CyoYC5I0PL8GyXzSWM
V4shNgTD4lws6OUTYPuDhgjd9BA9AGwkEQDcZqzxUSqwFa91z6q2qO4FAEh6aYOR
102VLwFqMSZlqAPnuzC4gqZ6ovSxyEiQmAkuFhHQ/F86lp7EwUTrHUrKgUq5lEon
6dx4H63TwSHx5WUg6MSkXwSKm1HX5jF4vM635ePpmUzl88lLC5TQ3n4ZKZTQBBO6
zi2yhAUoU4xxSW/ECy8iQYqNbL9cS9Qs/8sNGuq8GIWO2DH8pywVlL54r/gUAu5m
cLYmAisJxseYYz47IY15niWEOwGrQujkoS0lgzF7H/683ybWb+cTFGewUurDNLwz
pzpsjOHGE53YiAkl9RKVPVz+1KP2nXxcSjlryoJSbVD3BLfj+REpNVGsT5i7Ux8A
dmhz3ot2uVLcZuoySIn8pFnCBFmc/KQ3MrGlymTMHiVOHy4ew9WzYeT8TtMOti0R
LGMp7DfQTu05+yn2gds01D94V0vM3rJ/Xco2auT7xVX7G+jEP+6TdVkw3b/XzN9F
cQ0qA3eL0+fLKfoJZLpSsGWScUbvgEQuD1yGF7Zu+TClCJHBRsFlz20Cvwg25MHw
ry3xDgaN+u5s+VTTlY0jUKkOkWLk6jRMu30FRTZ3t8yezFCFJVQyQyExgc53CVT6
1hg01NZHc2ixDrHYBYib5QTrGJrxQtAevWSvZ02JXeeZBSDiQDNuSPtviGZYzimw
5lQeJJxmSoPyIMiIjh/bCWKbWOMgiuZD9UQr1VjHF2f6QRkOXoiiUm7l+xOu93Nx
J9XQ68i7Pa78zBkOKhRAGZ9aBfdKB9ARm2zyICYT+7IRF/IzlsL3gENJU5K1rNKb
GTny72VFUxr2rii7SzUQoHAgHxjU5SXQsGB2/V0EgRZ71tORTqlW7m+aI/q/3W7l
7HzhMdARsQ4A5paaa137JXk5j0omoV+DpaavBCXrZF32s7lmgHkfXJAjXThrgz77
C35B6rTe0JmhVUV41dRmKz8gB0AkXkA8AojkqUedvCA5VoAIs33ipGp0/dueDgy0
xnk9vXQFpjNiJj63jq1ykPtD0U8vmUj3CrjNbtCNg64nlrbdiR3DJu2FitP8gDR2
FOMAOoPDmUHmG2WHhZTo2zR78ufR14xNIsXaa9Q0+vKXslg6OLc1DbZIpM/XWlNx
bwA4eQaUcXTyjpzHoh0KhSqJlRPbftBh2hpcbLRWmcuxPYYQQlgKhSMDjHck9Gia
21xUqkqUFL3aVV1hJt3J8huQT8CVpct9Xy280/mUX+DhF52XZ7C9TwLNeN4EWzw5
1xPuu5U57z2S+FdLRPnloA9ruETx/L3jBRJRSdyT9QUgjBwsOlJcayHvPMf8E+ej
vJAUgD1uS/3HcSkZZ3t6WM3Qnx1mXDarH6/ptALVEX2A3A5YU70A6/vlvby4cwYV
9oAdlEzthTbLzmeBqvlYPAlpiT3594ZiAqMGJJLgALQ+bEI0Tlhx88059QuBX8pG
aUeyRi8ZaRPJSaYdmHAcr6SbVT+g2r/XTCRIRJO0oTMUPCd4fvoImMQSJ/VwUhoN
3vnLIgOp66xPU+5xBDuS2++L1Pp0R6Uj+imtQhL+TaQ0cUWX/MnuoN2Ae4/nRCbC
iMWMFnvrE+sXrMKzGC0WMf2CYSoyVkdSdA4DW4sT/APZRsmOxcyGlXG5vicUebCJ
FZ/wWKIeR74xm9sPpz9Ane41J2QIRJVGjmop5pqp23Df3txYsr2lvhI2Xoso309L
0Zrom+s0AOiw4ckmOA/LxLP+PSEfa9jogV5gdIB0LmeetRb60dtb1/vnliWYy5eq
UNzuxGdvy81oA5zDQIDNrxepf7LBXjmG8zArxyBNmFQ57XsVHn70RU8o7/BWFvjp
vi8kOv12l5EX117FB+efDZoiyO3Rg6hqJgCGHYqIH/URGEt+78rgOUDRXqtGzhwH
hIyl80m+Vl5qt+pXF7hZ/PnpS2ktRMEMmrHEhowyPJhF5dLv0v34TSngnN/ppSy2
vk7yKlSLR/Yel/Qw4imjD27RATRfg2LwysoCRMYLahoUyOiQwPi27AhdYcqbUZbE
ucNXN7E/QUMKxCBMdll12btkXvcwnlElwUPaEpAIOPo381cMh5boRMsvfCvo24Vd
YhCI9PLPLURUP00RbcAJ4Qc+4afLxtWt4IUKDOdgnBNYbSi7kZFm5utqwBwYO55V
ThFfLg/2VuVstrWe7dW14zIjFzVD2UXjEd21zn+E18AAKM+rnOzhY5ZNYt8D3FFO
zeL/NPHdZgq8InMJu0NX0RHTQgV6+zQ9Mwil5A+i0SUi63zubiN54dDSV/mbo6Mu
R6Oxbzba0myVeOLOEBwfB/rAobunOOoKfMGrSH0snd2211dJ09rG9ZVnRinB9jYM
VUdXDO6q+DOFicNAR50cLYi8e9HOqKQcUqQuSXfoQQDu3goBxgOkrqe3exjbrZmh
sN+Y+CignPEkf2ywCPoaLsWhSsNLgntcyvs34vBWv8ZBB0ANREk+RPa+pkj6APjd
ktCtMcI4VfjHrpn0yEYqjEBf6o2IQqgmq+Qq16n/XnrI7ptOSeXLzN5VmRapIMmY
bzfYJm0W/Lktrf3UBkVcOYwdl6kyOtNlbsb02S7n5VxEZU/VlM4PPugkEA+8O/e9
lUTuAb2AgYmMoDoytOKCnPLHxCBbc8x4HJEM6QMPqpMVSgFJPucQwQ8VAxupMjWh
FVbHIy4WotV/g5uSUb+1H9bB2TIRIEQkZXEqVoxtMJZr0ySkU5ox22LzCK9cZ7c3
C5Lx9F5CrUsFzRU2VVImqVg/tsjYhBjHvVuyW/0Cpbcy+xaGqSy60XduoxyM5p2M
859m5ThuXcSgeGRv4arMlBrLJ78PzPNZ4t8WtruZcVAN3igz6cwxZdbTr+a3XMgv
5uHlSe8XsBdjN/59gaufpDUbD1AW2zz4+yArBSnBPiKBLLLtMoy3IiiZgrR3w2gB
7yTS3O/ap7rEPZ+6fLZ2Cu8eM5aIgXjA7j9p7vKjbHW5jqzvREFDelLMJUFzOmpI
yfmMJrf9sBkzSygLgiCembDh29/2bQrQCmUADE95TavGllFbghlXq2g+NCxKqOA2
`protect END_PROTECTED
