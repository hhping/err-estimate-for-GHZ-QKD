`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqK/0QWSa/fi0S+128oESwqfhEIwa9R4SnC+JerPr8BMNC8JeWhKTGGelcL7ICLw
qTIPXY1zL1m7578EIETcTN40x28Gr9KTxaMYPmB+mDx0TkJB8SdpMZDYLpjtWtmG
rgjpcJAozq4drC/ZszHVf7MB3Vxl7x6H4LXj/dp7My0j1KR4ik/X8vB2sBLwcnJ6
8RniPI0MSY6PUnUM/i9u4hwU5tLbWf76nCSPqonZNPYWGnyHMUZcK4vpAxJQVdBj
zrHM4OVe3wChSAZ/fu/+cB6bFyl7pGwPbtD4YdggHq5LpisHrkQTaN0SyiSmIBSE
YTrkP3aYspwEDCK3LI7E6ovrxZb88+ArDWV8WJi8ZPQoczvCKF/COGeMwE4dNDzd
Iciut7/MiQpIvOVOih7KAABhJbSa5fxZ98gv1AsopxrnzvOOuRV8JcfPdoz2JcnD
EaKtCpuMB9bHjE5mbd1FPbJUJ2hqO5OZuP1BjDBLYuKNEXGKvUtG0u3hQw5W8jTg
u+BdAAdZliVQOSLCJDQ32H6qz+XbWvf3yAYCf5+KkByORLpG5c/wPXU2YvoyyWlN
CLYREW/30yhJVCQ4MGEMwgJpAeLqhUZ9LogmrCev+iYcsi7gmJdJ4NbyYEhqmsmZ
Tc15vDgnAhq2UAOCKFIA7Cg0pRfV7eTT67yBZvrBGc9PA05+ccyZP7wYIx+yjved
8ZLYYV/fKGSbT57tisksz+y5H5DrX6PK3J0SujHgTzUODUAhQEpS9b7L5cu6JS9k
2JPS7JIDBw20JMuYOZLN56vm7uuwPerXsucUK+lItO2fwyPt87sB6fjI1rN+kuv6
ciOT9KS1/MUfdBIhmGNaj4Qf7zVu9cAcmDCdhZ5B/xDZ22v0vWtL/87aVvJCQaHm
UqJDLYQbdzl+60GGFvSV9w3/LqK0p528++MdJHHHYdbjXvYBir4M/H8iI4oWjWXZ
kmPUTBW0CrKSdwJ7w1fMiCK8fmavXpuJpUG1olTE8oc99zHkkVKQsfzjqKvJbtRv
aVZEFHXYtk4fN6iIpSTA1qNPWMFP2lomn9Eau5pGd4wV9NsBZ9JXO0ke7D7ESJr0
KTIMp8IIKrz2+U8zBY60xpHqE4ZP5lL4d1L5adSZHcUiw0JlxCfMzt9DAG37tu1Z
bx22Uyobr9ylEjIAuVmLIu4Yvlc7n+L+3hy2VHdcjezjGPo2lLYfENBb8W7UNAWX
pfyaYdolal6LH86E3yVRv/hRLX4uJH4dJxwfz7+ikJHLKFIKYmgt4Vmmjk3oeUex
Fp3IbvjHN7QVwo6BfHUOxBbrlK2h2/fxTeEspXTZONChNGZsF6BXTQABD6pemxSK
KeXNZ2lFpZIY7cSK9SLJrNc2flcJlZ+VSdUH/FC1MoYfZ0eftH+9Qn+jY2lSF2s7
u9doByjM1OoE0EE3R2i1X/zQri6tzazI9Tphtnogfx9TzBPygcVFyCRWHO9dQ0WR
tQ1kJkqurSCwjEMgzDAaT+NSI0fbrNt9RAv+XmiXo50oMNztNoUMF2X7xdRMSSmK
aai1lLO2Hk8Uh36q1dAeyNL17mgufd6jnBDIH/Bvre7ardknIVr1P5V6lU7uDK/Q
tWRiUg99pRjFcZ4q6ePgRCULmygzNsm+qbYOwJnJGpjKR9cGb/BsQ+a6QDGdyaFh
elB+OvZO1aHnjevPi3PY49JFWPJZ+KaioiQ8lS9M5cnKK7IHNBTjTwKFhc8QPsz3
DJuHRYb4O99Mx3wlaraJZXK7ZIUBbDe2fMRIlKag8qYhpzSJeoaVj/6paOPX0uXm
uFX98j87GKfpIw+o8mRlfbDCfvvhlLYw9tuGpZIWIeO5fIrVMC+wlYx/LjxRQ0/m
2efBMWX4NiYDTvIGrkLR9LSQD4/fv8trIwgdv+1H+qlu7lce4d/GJiMR1RbBtmtx
bVMXKBn5Xwmo32fAvL50OWjRrFx4HYrjYuZfxocuZ1zg2rril+AKr3peWSnqLOLQ
t29khFCgRAlY9HFRWaJnwzxZMm3BJOvwNJ0RN6a79JepIb0Yp72na9QcbOFyiauh
xfNxn32PaB3YpPi+gzvulZsCFz7CmCyCSbFJGk+rQAovIDnWdiyVeqg0YXHtgy6m
9H1On0a/RJ7DQBtTlSXexLNmh2ZeAUdrPT//VLsOoKTibaKnZvfDmieQ0WpJMDcD
6ilrHg4G4Iabk7yCVj8QVXyPBwZZek+npYTt6znVF0jFSu3tmVUgIrnCnHGc2pYz
wWP0mMNI3svZf9klV5jhGgG2BTJY6hqsqZ+AUtgCnDZSrRM1RMTp1b7YFgJnuEFt
IfgVibQtodq8fF3EhCtmYjaxvW91JxtscMuONsxNPsAPol9Fn9q+6IoKBuWKghq3
u2YcfVDKk7ry373lncUN7pO+tN7R0ll/g6xvNfV3hbJt8xqk5t5+WPgAlJsuNm7D
CAlJEcnU7x44lkkR98NJRoQ2aa15MCcNnuai7bkHnxkB+xorUBdZCM1XLKeFsG8A
WrZURtEBHrR/RCW4UXqR8hp8VgXEPp8ysUgWjcmhrFDBm0Rp9aPp/HCW2W3X3hFL
nVRupINHYqSJ0/zgqeyCtf+D+Sxdf8X+HiUB+BYaNBkl+r53Zq5F3sMaUtYJ+Xtj
pN+LdfuM0aVfZth1/BZGjaMr/daLOxXh/UBPWjhoo1WCVTgHUYv4lHMbrv1fggW6
IvqOgisEVGhT300VzWxMmFb1/dtxxJGcFhXe1SG11O2uaNISxZM7L6gxcpaWL951
dv6IUS+y7wideD7nEsYsFmZkrFClSKfHhrH7MSN3ScTGkWN+N9/DBNu5of2wAo7T
agHsCNGVtqlR9er2VJSjG/wqd5e/U9fr8qDgZ7IYtAdeADThFXORwAV3/jcjV2nd
iMQKCeBRUz4UD28u0+cAvQFSR3lJtXuo8ezUSqqjZ92WCi7E/5HI8E91nPgXQrKy
8Qu15lR00PH3ohi6sOHGDJHwFPeTCvP3IsGPugQuO3fS1psoRrHA2/WkfChWuUKa
4ZaMtcniY8aniVFu0PKc6WEOJeXBfxcHwBshGyLTR5LrcNp7fg+yyx51LcEhyMEi
5W5KvUT4fV6ZvuYClzFtyTLHR8cvcAt2+I+61Jm/qtz/os7xL6CjCkOM90xhhsB8
yQPy4NmirsJzmU1Qrsgks8ibxrO1kKmlZgbWCOyGlvOOWLi6hRjdGF354dVDD/mB
RipTy+zqCBVFfUziHKFQGCajTeHqK9q6gjF8MipWFlvQY0yviawkSaTQVyVPcumB
Jf6mMHOmaVs0zGnscZVwTMuoYlVsOI0qLu+C5NXYOcmLsncuVxw55K6FTnqGM1eF
MzpzY6c4m75WB4tgAXaHwDQsoGTzOiMR7zPH28SPORg+qjD5QpDCRQHItRJsmovW
fh/gC9EGGlobTPxxRi6fmjI0c4lph9XTA7nJ5gE1GHOob7E33xxsyP02mv2ejq3W
IstX3ZDGRcbMNdmo9fI2wFCHr3liHRNypcAGVwotnpUzAAvAlWenEPSEYvgXqFdU
kW5NTxO8qAp+T++pYEP3Y5eG/pCvWG00hix6aW6zyLCuXDNeT9Wf6u/xZgJglT/6
Zr/RjSNUgTGmyORLS/p/wanHw6vmKzmIefDxhTR55SDFUbXCyR6nXRz2MU5LCuMy
4aCSz9Inc9/BLQ/JHuMxUC2j92vg/7EgGI1pHBAx08KgcP8UfdT3YjaIzRqprDrv
ncxP13JvpfcqZ7jqU8416BVZ9m1rSQ7mAsxXlYeFyu+gDPYrvbijiLYhrVkHTFhN
KUU8TGHAxaM/bd3NjJLFSkppgUsqrVXSJyZaT4kBbPOoyv1MZ2SNwL8hZYKlDTMx
c3Lo1rcYYHZMhXt4yu0jabd1VPna7SCS/9VPEaVKWzrHJ8qdgeT3AXDGu2nXySEo
rxc7iUyOCN7Z9PLBrO/bFI+bR/7E3hyKkhEKytwbSmLnmfhbx8MxLxulytZL2uZR
vtBXsH1O+3IAZYt7pZEeecvMLzCNWLIvb37I3Qeo+9fL3zY3M0SshmgQvuAeDVS2
5OgsEAARjigrneYfje96kh7X7WeDC2b/Jhisl/MrUeOd1Z93l20EQK91Fph3d4Sd
KIreXjeyn4y5TlrSfmgkh5L01sinaYfcRiJIXpz5U3iSYndJuCSFFtaDBX0u2zgY
AjnDFOrttQDubwPlAqCiXvIEfG7di6lPNXImnzdk0BplaLzGCv+YumIKT//L9N4z
3mwNlnPgz5pZnZeks8y3ZVbH1EJdr3Vr4bKcnu2iaLYPeW8DCoENIpMtsyCOylX4
GR/x6tHQ6b9bK8r4+c9xJo/uXryu7rI67nV56cShU3UQYf76v/YlR07VhjutT5R0
3JzGnSwAqpjosILYn1sRdS1E3qexEylTKgJGQXsqQviWgsqIaKhQEnQpzMCkET5V
W6YPP0fLpgjyW7GXe8IlUTvhlA5I9zrxCShEG6tWcxW5km0QnqFX4hoXl7KttuGE
JX0UaJEYtQh/5zWalDToaucjY4jWns3lvz92CVOlNEYZBTOFY5Ph5WNDcIZyAkcE
BdsYvGmzAbsFb6ThA5eKH+AQgB2zPUtuBsmj5wCb1RMrOc8+iZqUFqgEquKp0TRz
//NJO56eNxFmxt7XVHYJNAeAT9UW4Wz+6cTH2UEgibs5wISmdXyye2tz7NrWv8AU
kFxRvxb6V4iYzDWOAFAz6lkyE0aY10t9QphpijhfNcIJ7UDW8Z6WqO8iGDDP743t
5uWWh6bX2BYEFatFYStq969Ql1qH9Ox+bVMdG6SbhqXi/rwbTMfcV90iPQfEzHUV
VdnEXbJOLbVQYIEgc1x/I1fW8ASXtYwjNvA74YBR7CxpMrg9Mbpe63mGp0JsaDik
zZdME6+KXgBCbdm/cvUs3heLZoGDKBCprwol/lMqhUZ+C0AlRxDfloaz4cDz7ZBk
zjSxOYuz0CuIy2+BhlZGpYRPSMCDad6bgpoz1xP+UL+DYGQblXZCqho+GrNpU1nK
mUrqE3LvXV3Lg3ZpY+3f1juweAOvDOdhh8gpuDu77/dpfgHSXHkdrZsCXsh38ZjP
gjTDLuMbj0ewsNk0uPI4hjYbvJoAJH9F+0/lVLXMy+0QnXhW1PzjYT7wM27VJPEf
21IZdB73A6bHtfvOQd/MRC+rlCkUwOWLDEng2zXxCVDzA9fqKPaHs01ml5PLdOkt
vukOsFDUBu8Pi+382eCyuI+fiR5qvPD51zGaquV2HLMzBv/40qCcoVuz0NjaoO9h
V+/H/QpS2KlDdwNbCjWhXk/BxTG4BzH8NnD6g91TM+vkwr/9Dg9nodtq3cL0NOCr
LH5l9zzWt4us/IvYEIkG6KU06pPFleshZ7EXTdZY9RASigvIpsDOTE9rZ/Fjd08C
taG/tlSuyydYzv4OIdxr5HgjpCYKkhxYC+RghzIcnsFhbWsnbfwnvoWM5sPqjIpe
9X2F+5AA0oqLAYqFAyiTckVdGjIrf6u5q3hOaBOehC29kO+xi2LkVR7hWZoELQhm
c7xvGA+8MyaPyg6PPLnZH1URIN/NbrleyolOAbUgxRFH0J/HYTgDjgVaS/5qVlO7
IV+3Wpu2h1oI1n3RXWYAd6Avocxks+0ve0IriGqBkxJuZ2V5Zs1X67boRicNcHL/
zkb9izCFKUjL37kYPtq0m0WTUEtrY2KIAZ8O3SBX5oPIB+3+yUTClUlARAez0K2s
BbbnMLszRZE+NLM84CzYcZigen6Sdz3N5hgeBqbv8jaM7QyUFmVu1+6CLArE05i4
8nSCzaGtQ38BzjZFy0ihlyPDW68Z9/ls2qYEC5z9+YRcmriMGSgQVXdpAEvQAz8m
fhIXdjphLIxEyabwSRXGlEqAwg/6UmjCMx9UVKiwl2BZ9ba9VEBC61AlCyc3fYzp
Nh08XyGKzbhz9XX/kUWJj7pNPf5KSX98JiwHwlSJY9o5oPfnllgDWjc1EzL6ERvr
JTt3iRWFLLwhqy9wuOg5NQjqQfu/q5kLMyoKTYwjfZn6q3Nqeo0cWrkRyPbveS5X
AZH75/wdHHVnKA9yct2M6DSBB2CICCTz807PGXQIjShpx/PjwXYfbgmGk5wPRVqe
fbNHIYyw0xPduDZq5BPkg5b5W8czwqcxSoBd2fINNWD+wNhzoWm9517klnEwyaQ6
tMzDCE58io/JEeHrvCGEun+BhxW0G5Eo7RXgzH/MeN5XHjEu4F9xrLS0Ja7IgA9p
jN+zPCxeuLAgvJLmdnI7OhBDQrL3OOkj1d/l8rIOOBM8qNhP0YsFLcEpah6hBkjG
IzSU3lMOvjTkj8KW+gAEekMwhxiWd/upX+ThqaPqx0dTbpmbei/5nkvkTXK8WSjq
IG1NYW8e/jF/DMN9YPMUOtONIxNzys+MDf3X0p1Y5EautDRWCbxVlygPkeGi22Vj
KBO6C0oPJdxQ9+/kO5nnEQE8Epzpkot/o8ur0KvhHcT6+UA7FYHKcnkfnq8KfmQS
WumDSZQ9kbn63nLuMhrsNFzLic8Wy0V+siMPDPuGdpcv6BJ7Cp0QWIbdKLgpAJp8
i8y3NekBCCRCIqkD/jZ7JByNGKVVivwBh4QhU/bRSgvnNRWwqrfmkCLBLmIYhwPi
JtWRBZQS7jUJtOcaFNajr+3bLtJwp+XcPtGERQAu3cctfYdOOc46Rc/7WQvQze9G
NZPR/1ckVy07vlvJkJoDdYgiFvQoDijR6iX4pG3nDA6QH1Bk5t2Q4nT9fkHhZXsT
SlkkkQfFaW0x/qjw9fiLYbVAJ+WppJeydzciw31ntOX/lHqnQ/wI1/q5TuLTuN06
KVZ3Nmr7vfJEd1BH9yby0AuTRoSuz2NBS8kojk091cO0yQp/0NRFpcNPyMK6IQTm
xhCrUS+K0uxU4E3aTYdc0dTVPSDqseqPW+/Uw4sMNfrdzK1lLqgjWeOiij2B3PhF
9RrFdTQceXRtvqzcDlR7SeODSewCXv/I6DeBaV1QxfXobhsVJNj0sNTk+DLQ8ZfX
d+/NvClI/ArZR3qSZI0UGyd/2YYwLSsK/ql5a/NNk6yl0TLyTd/KzKk91cQmHNAK
+QkLr+trmGxWOMB38Ga6fiPUvprAdWvwjfgKLdxhGtDpG1bZYbvH8YaIGRPRAuCS
FpzHqvTvbGSksCyimcfL/qa06Hxo7NYT7j8eyfgbw1oUq/kvJs347UIImwtTdr5K
DRPNIpw4jz6BkrN8bKly+sddtgsNOnQKWRdsxoujoHTzZEU6F5+fCGdZnJdcUWT6
wdIz0J/bcg9VOPtpRFk3oNXVndIJaL1xTNWDuw2sQzXI49fIsyb/D2sgRPRaYHIZ
Jp4Qp5aaLfZfZwNLiXAnEo8XxRkryo1tJeBt2NgUdN5HYThilSla0DAzH2Ypr30K
lfJL6zrJEitf8Nr3qZZTxrxGpj64Xu0T+4B9bY45u9FCYt6zLsRa6zWvCCLcRSd0
G3mXTRm3DqGZkeZ4d6qp/ezZq87CP62W9CTSpuBFOOkmyQjw6kj9ZP0cbL1nu15u
Ifm8Z2xv/dyqcEivhgfZHnepWB1wF3pblVcfs77u7RE56BG+qKnrUOKwTy5uReEh
FtvmRBaF//aaMQnxKHiow+H29Bz0Yj9kRb4ftXpW+JVr1XE4IRcxML6XMd15NEO1
1gptcmXhN58i5imptUnZ5AcgT81ZAR1qxP3Jj9D5WehsQ7GWTJFwhvevy4v53vB4
ANodxFBzIjI/13IcmhdErXftVutsqmvkUuaRxDjuwZr6Pq5iOZdacZjDQWWJhdHh
4kDDub8uts4gtILv8TcpobQN3k1J9Ux7IzY7a1pwISiUF/Nu024hXvibN7AZyEG/
16iMGFHpjSn+rd9wGxu4pdgsehjoaLDFHj2mOamxtQK8fSfbrDzIP7mIH/djrb2S
fiHM4LhROK/V1GIrJAH4SZkYabHgExu3wPcSrqV3S+OZGRMGKDOYu9sM24Ffm0IH
s4Tz/WK7GhCNzDvpsuSCp5HObaYrLiGdeow2vwyJ2BY7D/vPUXTxOY9y+3OwoDyX
SQGQ/wQb9wg+KNtWv/TlQbRPvPCngTyIB/gtRRR5LieKJyURinvADqmqo4Mnlogb
t27u2aUv/wYgsrhuSUMknKjUORgXBvuZUfV8UMI8gGszZjzOPQUX7jV4e9PuNL9x
MjlkVz3ZiOB+3ZonC/HSy0+r4rLbf3MzI8viPs4Jc5w8UP2kpd5Bth9/jR+bo5yZ
TSleqAHj1+5xvNxwM2WbTcUeqqgp1417rFaOPDRnFeCnglfIggbzqvFuYLoMbmgn
9bEHZ+C7wwLRjWtec9sIvyGpMwyIC5rFlo/W+WZP1AK0wexQAH3uNTAyIqzcbTSg
9CAxydDBeuBYV+IfY7sNuKJVlE2lpRzyd3MOHfSmojFCNH/jsuf3Zg3yXCQBo9ul
q1eRtpu7hunc7PIt4z5j0XCSrb2ujz5eZrbmje0X7tbA1LSEEXTbjiZX4IZGM03y
Se+2OqtiNhfgscxRofM1zl/DsPkgK32dteOyr6ScJKV3kRunmJW/SsZ8V5tjVtRR
rEqmp4JeDgh4QaRCAmXvbd4OzfQi6MpKKt7mB//HU9s9kYRy+Wsi65Oq/ZttTkJ2
i0ZcTeTe8H3Qoqr7SdRQAPnYAEbT7fhjIprD14AM73Y+SYSi+QD66MMyAZi8kg0e
CTMCFwngrl5n9Vn5h1Y/Czz6kCWRf0KMsAwZCYtjWKMD0gQaWFE5i5VeGO+eMzhL
Sy5vYvlVi0ilB3uJjdODaA1fZi3IjtO1NSbq2xG/1Sw6mDahOC8aJF3H/qaODKdr
o6urG5UnOpcBK9CXUrXXtqEVrFACGhj68Mf3DAOsKMsQo1sMakCKTALrpfUWLIyw
OvvbyRIJCum00DLpnajyjOciin2xczqk/biSHaFFJqDgaziA6O+HDKoWlST4+0SM
/WcszRBx07OB+jZWXjkbowKAcphFguPx99VrMPBVrNAe/1uW8+HV+hImeQIIR/VG
0b1vvtxqMewRkLUzbGMMPEJ3gW9OS8I9cQoFq2RG5yoxeGVGCV/Slx1Gt+mGWW7d
5zNqRcr0mSnYD3FYQi2qu4wf938wfYXhH66n2AcNhWobqgj0CM2Gbhtmecvk+d2s
rkrx+p0h38ewIPyUlXWEvYNhMA1Cs/8y54baMJ9/r5hqQa0n6mLJIlOOM0Xw+ALn
HLlzPE19jEp0l08k03c2cT1z7SDi2QjvJVTdyoZFbTOGPhUqXgLKgF8KJOJ7N4Lt
FOCgh7AAV1rFzmGXa92Q7ouN2UqxW1JN4xw9sn5m6gYSPP8p7ZHqYVR3QmK3+kmm
kYzTb0f6Ldq1cmIokQVHuvkhQPjTnAyX/AYqjau4c+OjOfuXy2MkmQz4PtMJFOxP
WtxgTSzt40ye2p5COufFEYPiKKJ8y2BvntLJTZV9hHtxglREN/e+Nd87beCqXqUO
z7RH12JbbEIJFjYYU2EBXLmz8SfGkoJaSrGetAjFH7yWZvH5gprRfhXEgdK9+6/r
6Qvm796Ne1ArAvRhqRSfl30X21zIDz032VR7DRESjKCrMtANNfWYwTbY+Mhwh8hj
drdCw2kuWucm3s55R460vim7m2cOn6NEV8YhOeh4jSPZNU/bacf7GakESBfhdjF0
GyVho3oc4RdNVOOpXDrYlO2WBNVKEXWHyRJuE768VLq6ldk/XTS0Xiw0+fyxoZdH
usVGhpn6Tc5EyBlKSy7jyrhkrJ9A7iZfSWxREpHfJsd6iYipgwmeNd2EFlf8IYM4
fi2Y5iX0yoFTbV6xIuqFj52QIqETjDbDPax5xEC7aYHovpSdthLNEam6ovFzDGGl
Yrv+wLV/J6Z59GAm5pufPO0OUoVk2RqpQgD8Ku9/aY1fAXTFyVzH432EYKAjagb4
TSYvndOwge5RQT//WLCf/tChJno0vWab4n79GrdHwCnDxX1aSIKNGiCaCcypqsjG
8T/WujlmyuwW3DuFIWTlMvHsKPTdEJLhvATVXhcHIe5LL6VVi2ntaou0rxS6+Cg3
ynaDRAn1Vq9V3J1kX1iIiP6JKImXxghl4VXv2dLVLxuAkxU340U8Olo2YYZnFsMI
QkkZx8RKNDtcntrNtRox4ktm0Yu1atLyxEokXeKweNDGsPdRrTHscy54tMZ7XgGd
u1uQNsYtk98FJkmVg8MqvLszwCcY1VMiZ3GF/ArAIw23OMNwWv3C+rojTLE8clbk
NsezLv39n/HC1UQMfYGBGIYsJ+I+YyUdtNe5JZocj2NUv+x+vhgUqsyEG1zgQBmD
OoZsS/68pm3L4K+So1maUwG5EgPmTw1tZ+GTurkJRjDtf/NnDHTU3dEPGaSLIXrR
eB8eenaj0YkWI9GPEOqNdIf56SDzSYEOu/1e94XN+DQF3pZ3eDfAylATK+TCaDMP
FdAdgQ4jgdRkvcrw4Rteu/xnpMz0Qw4O0P7a33bU8gMb+fbjqdpyIB4nxnS6zdcW
JbxjbgzZ8yiTEWzmKysnptrsmEn9V6uB525Og0GU75DL9PuU6iaTLzHmfdaL4Ska
OxDM8EsHZFA7oFc/kbWmcGRmfPIYkc3zUCKPIRk+AlnsqJ3fGUcBms3u5pY6w5+5
v1ex1xc4KkFvXumg+ts3ntun4TveGmGYxBJ2zRfi6Aa2htRsHwGvLIaS8ZCCdrMo
jtJv7Kb+joHUZTZXbOB62vLm5m3GdQcO0WfriQT74yTpqHr46KGysy+rF8TfztR2
NqqV+R0X7bA0fsjlS1+lQ9KZo7lf5wEijuBHomRYm5QzcSmzk2Evb9mOckYQRWz8
xs6JmibNmG1Ej7oJ/b2iLcqwRwn7FyznhxotB0zhm7fnkRs+22/YWM73zENaIw/R
yfWlCu/cWBuHbkU7Xp7nOBhrolNhWMR5+sqqNjaOQLG7pwyFtGHAZG2z68jWA2t3
Acd6XYGjQo/FH+gODOUsOh+/v6dFAgN807IMAQQuzP2b/A2qnUIU/lRq74MMy9OH
DXK5CRskUB4/Iy1hLodhvrE0QdHPgoKIzUtS5bn3RDiC9I7OXYb5X0iQqztPJWsa
xk1m9bQWs6hYbSIEItLuf7/hJetKyN37TuDd383nzHreZVAueAaiAeg9QprbsxYt
kRheZuuky50vwHoBeh6N/6d5bw4EwSsailchJtoAMcj53tYG/YZlvwLBjOOmqgeN
LNYuYtK7ikoZ5zxhy3KY4Hc9wdErrlqMcJLbAVP6GqFpMZ5lrSSAWmrRvJ0L/Oj7
tg61jv6CSq+KW4byWqa8yxP8b3aZttOcImbq6p0vxJk4di3NIPtut2BELVGIBpSl
Lg3e5rAi0hnNU789Qe26UEHBUoJcKlilKtbfFPtwSHkARd+qAUxgqBxC0lz6eXDX
+ZO0ZYOJ/lPQ3JRRXUA+pzcNfzg5imEkgGf+IMQGBFNoHx3lxQZiM7qoSnVz23yd
Vg/OWtCfQkLrI7o4zgA9ccDAeY7Tr03YNLpAKeS0GK+n81exJ+HVTU0C2cPHYxTD
/0vzax2b+ja6u3CVXD2CZdNC5pMe6nhmzddPeD7eKwA4XVodAV5mpfXNEJwtAj5M
6tGD2yIBu7roUUnKtJL3xQNJfZzJp3nqcnSsDXpfvFJUYeDIL85WOXgC1TaDqC4W
G6keujzCwWqkN/4HbQxZAi4RxyS8gWix2D/MZgRUXbcRzKFrhotwWcl7wgt3fxQh
dFZ+YjKpev49r9IwmJcshVtUvmmk0bsTHXZD1emF5bWvA7wlU63vXJza4z5M6WbU
YXJAhHcNUknkj6XjeNHgIPBuXMxAPWoOmGjl3sZ1RqxEwL7ux+Xtq0PryZ+iZo9j
jaVvM3Vk7lzaAxxjimZlx2sxlYygdzPJ+RerNGu289FSGcVzWZFOTO9qxLzyL0jR
qkb/UkkoLDAp3r5DHVRLcceal38uWHyrM3U8djYyZKslNy0SJyGLKItZ+Dma1XZV
CyHpMjEwDQwk+45Jf3ZNuz8jhU3xif/vLdejQG6hFTlKGzFgJb4Ihm9+gbWUc30/
TJN2wCDfwU/41qfiY3H7L8HkRzX3OVaFH9SFJV+AA+0uvxGwu+ySQ/DoqtZgiznJ
NBkIY77/NWGz8KoPUN1p14P6zupWqtOROK5nbOQxUFdZ2WnNW00OHf1Qy2ePqwM2
Bbrere7ms/GXzw/C1e7JhLC8aIsUbjCaKhYoq2aoNkEs5CTA6vu63plPVIkL3rOm
NabUlFOk6ygAltuKBvO85ff0S8kVvwo5rmWcZYSbzpPpuimMTYBKZL3OqlGTHLgN
kDoSbUmlipWbizozdIBZcdrV/DpOmlTd6zoGDq96krxzZ/8oNp59ENTl/i5tREFW
DFbSeH3L1nJONSIPb6Nwx355zfjOHv6vAtbjGHpvMOrv3J1AKm6kPDvUenweawOL
r6erP9h0cuVNDOTD/XYvoz5IeTM62pUiutNBRUbEuEeXCAxFeHN8WQcEpOMav50M
LvlSJ2lvm2RJw9IRP8hLrzXeMLj6q/0s8nQ08TM52PT6djnE4SXeF8aMzpG5Dx7/
1TbQdD3Fo+GRtrud6pKJ/F2OlXn7h8m0Q8pNKH9hrX3LGJx5Hpuul2X5SSNSs3vl
F16Cd+f9znXS3YQmQGzKWBWKox7S0h4CP7gPlLYskD4hGfAf/0Y+q1GYTtBmI3nR
zWoHkWV1zuS/eaLx511t2/Q96f5Io/UChRpO7xFwJp6qa25JGr2L7B5JwxoQHmoK
KS9e3p/99I4xc1IE0oFX2rNiMlvaG5SasoMaK5iv8OvfVmc+SRMw+esHCVokVl0y
fCyMxvbIeOZA1/dK3l6/78BoShVMz/IQovG6iR7A1lBjF9oSTl3focZVTYcZuTSE
kMSr9tT/VWpwUnDwOFv5DOywo4E33Xjz1E4akz4i/DLz8mPcY3VOLG0qicV1nbe3
S1zjyg/bR1JamuXgrJAboHVrGlI2msxN2mus7fKaYK/LPokFcwYeuuphweEcPskI
G1AJ4YFQ3eIWXlJ0/zQuRB0Ox3JnN79s+FIqljwCvg5Eu7m9uHxxhlxbcTyXE/v4
xSO14ybAV59l7IRrLLWBNCAtGT4y4XAVnhT42P5Np9TbEIofwptwcUoueHjBM8xm
Pb4uL2+2rA/xMB/eBzPD2yVHPgZwKfNE/Jo8NAvQmGGbljUJ5Sef7BYSEuqDwOD+
/g2HisIYJ5QL/rmKnjo6oCF5IlLx04cEYN6zLodlscgBcsDa/10txzPxX0le57ql
PlruOVB5jCzs8rUU0OQRxmDHcYwX6IKlox8reLZhm4+WDmBWowx3q/VBKFsCTeHq
0Wu3ZcJ5FiGTIY/WW3326isjw2nTVpTiJm8Li266b7D1kjZ3FkjE5c5L4FoJQ7KX
BH7LYoM8Av9WzbiP7oVEzcgtNvGBPjhKUHYjWCGYfDJpVnOLc8tW2XvTzPDHCa18
asW7Yp+0F4gAYr8kzR8Ahr+noKU6t/IBzSuVaKqyb/7eIkLR/k6UpXx1kEepxq0g
+nKpO34lBHKdw3GGOiW9a1NYoFCUw/tbxIjDX0biI+SOfN2fbYPVE4GLhpDG0u7I
laV7+gL15GHGk0fCjNysvgyJAa4XAUSmyBzCswV2EoBavGA3+OVXZ8IJb8xC4kh5
zWJYMiAa0VT2XdEbSII0IL5ML/W8saV5/jMYIWaaCA3RImhXagwq2NUHqjnBTe6V
aBjcww5hKxnRJZFYSJuUe06ZKi/s/+5NomBpIdgbqzRtMZvkxl5jB3IcAJHHbUst
ymhd/i5Utm56mNSy6f58zifkjZjncXbz3QoVHD5WgaT1RtfqXxuTWlohLLh7Iyqy
NT1gu4IqGZyi/CuhD6FVeTC/4xQaH3WnPKLkBEEFadAjgJC2IbK+CuOwPYRyx/zE
QYT4J3hVPhIJVl/kFCHU9SGKGRzFhX6p2ph1xeXAbv3+0j8boTqktfYclxvqDtKt
L4QWw5RFtz7+xqbl2CHG/v/3nnvt2TpsaxZeZ58sRaKHUqxNN5dq94ww4GlC/1Oy
JNuTmdW4brRAFGyiVcTHkKf8tmMyL2WbVsU61Lq6J5IXEWEgAioJDxbSvyxjKoKd
x+K2Q/8W/QRE0EJomjxWRRNdkjaW+9MEKxZ6MEY31jOREecrPe9kLlSGBqyGz5QR
HQ2lr+ersah8yxVX6vZ09nvRzdpXcpvdj93rVXhaMZceoW+Kx3++36aAMIhw0oNs
JII97v5HJxPhb4Jo5GGl2L4AFVxkJfFhmWXMnAsJqhV8hI82X+Bzw007uw93Esgo
hKTCoe0y2cawdbHqrG9A4Y8Sk8Ae21uY3YZqezBEgjFVJ3RJLkB7Zs+Xee5frY+q
IrfdHA3Ji5hFdUvQu9oPWDkLLEISoNy6wkxEH22W9fllyXfm2Tp3SOIZHwX8xaxm
0Yy2EcIqWvkT3ATYj/T8VViWC7/NuCJUolsbB21G2jdjbJCJBRjGaWsg7G1PglWl
E99t925AqrRyRriwjGTvG7O8jGq8Rf8kVA4G4nGphaQhlRN/tCKLQVE5/Av3k1fk
uk/EpMDv9P1SJIPNsEtj8PykIAS4HbhPxu8Yj5Q+OftEexukmyfOdEzlEpdTOYDs
0hAZBDoplndrGJCWxXw7/0VQlfq2z3FhBaTaqLOKpsBH9oix1pzFA/O9NJ5u7Rk6
PYW0KV3WFl3EPzPnBgDi9Q9GZXNKb5bw0K+M748KXC6vtgnJEcTkERFXS6J6sksZ
qZJ1k7WOtpK5Xj0noqa42IqFnAXeNO+1VEEShF4fnXj2JQUlxSWU8Mk0iyt/odFI
kL8YRgN9iEn3SegRPOzyMkD3qicohaZo5VKpW3mswaON6jUiJ0DEzC836YR3Lhzq
XtHDBlQ/6PdVY2RXXXzeCbln9GJ/4sJ40Jhi0cJPdD3CAxWZLqc5LKXHoWnDhbeK
Ju3DymIYnU1YjXYLPN5bB0AvNujZdpp1myycBBP3bZSg32Sy8/1wdmgpAuaaFnBS
Vv4+BuGl1gqGj1FBx1DUHOzSyJKptTo9jXodBdvzW2vmOUexEKStTvGqUwCvZVgR
fGxx8Yw+RoH1UMhUgw0O1RHL+uGqPh7JaLypAiuufgT6UZBdhBGxnKo9/wjPjmWp
fRhwYzgoGseCDpfRqDVV4Wux+w0h6g8cDnnfgWqh74eMR89O4QKGZZ1cndoay11q
ZPoT8sTROBo1YB2lmL7o8aAaNQPsXRfLAPzhVAHv1czPlzANc07hqI//PvGQWIIs
nnrjymCEP0vI/O32r/YClat9qlpDbIKLwOdJwf6vltKZTo10nAqr6Bx55XmBMxsy
U5tkpCQGzsSatIrj8QduM2aRPh5q/zg8+Y9Hin54iJSkAABqEj8r8za8SYHcWDX8
3E8c1d9oERIHmLwFOp9SvJbo4DqZ97KD/dkoJPWdjbGjzqxd9XKuXNOrs2YjY3r6
thZwmZXHsJ6/XvsA1BSXJTiiYvK8XDr9Ljukrt3ZvZWSRh7nRMgl6N0+UE9imjI4
kv+5yubkhPcKCPzEF075HKW92iFFl5+760NRBJx0Mr777TA3mZY5642uimu9u3gM
I5kQ+keYSMhfSpoyGER4M54+YeyPIUBUkXEg4FTstBucfXaYEHUePiCqNdyS2RhR
uTA9t/0jeXhfXFJXB/NfEPC0LkS8TqVh54tlf5H9GEt4pQZ9t8qr4rXBi7wGr5En
B2ZLditazS1iJK99FAKtmtCHs95ICkHnhySZ63WqKpFU/1YFbqE+x3K6azFO5z61
Kw7ZfHOB5C9f6gJYelFMUIXXTP77cbUvuKy6wd15/1vndXBqN+ncfRar6dM+ARoM
Ityia48xhVEyWvGfU4gqyWSqENpjm6eEI5J01/jIQSls21LteeEMmOGtDFBhUg0Z
rskVwm4HLdErTcAXjGkfliTtwpS5PDwOoljWrejsaQbph9+4wC24NFl98nxyxc25
pc7iJN9lysq8qyy0RZ13Ayxws0my4eSiTwbHPuEQ5ooYMktOT3QjywUFxegF+KBY
dVk7qOEB19uxlQkn9G2Q5hcmeycYdVISGxZP60f+FUUz/6iSMlvVWSBtRle+WdQy
xZaOqQYBmZo4vH1je8C+vEQF4JtX5TjepmWGlgQXclwtEZy0Lct5gYT+MmMvslaP
weUuR6UrqHI3jzrA62VZmGk7R7zaBjeCv9aXt60l19HBtfCSOFv8/vzbaK9aFp1p
jQ1D1GZwkBCLqXCyEe/ay2aBO4uLeyMKsxXEdLC4CnbZL/1yGZY+1uCeqtGgL3o7
jilyJ6v2dXxWEjLtpe8qM997yzCKqOmCtewUYj4FJO6ao5QkeiJOumIbqYWq8/4a
RDfE1697AcnJY7syeEvXOpTz7CfB6esh9XZTT/DYngNIZ9tI3vQTM4uGdZkr9vN5
jeMWUTqoWOCMJaqkBreUW8ozBvHJBUbkyv9AtDPeXzLXxUZdxGl8FY2b7yN08R54
tjQeTBlhA0pGrNJ2XEoIUH+27Yw6Bkm99aREPGe3Zx2IbyhLqqBv7Hq4TPGeZ0jY
MfwdASC/SuGMw2bbscLMWr8v+dH9TMNnRTie7IfJbXn1Z9GKvc1rbtbxI1whFCS8
3BjMi7+naVLRcxWn7Gn7sAysM3CshxjWmHVYdpxs/mg=
`protect END_PROTECTED
