`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgDYPdCHI/7qeEBj0l3Db2zIxjGmEC8GvCXiDDwBShzE+OE6ch0y2AS5DzuMvc8q
NbR8v12p38taCUNrly5Hz8lsKjrlN0NcEBFcCZxr+DZn9IvYEQG6sTViRdiarxTt
7U6UdXLbD8Kdb06nb4ogzWgSo2mHSH5Gximi6GCNWXiIigAUsahCIHkjSafsDv9J
j6FRvtoYQ7e/vURzm4ucZLrH8SgKi7/JEZGZabGfL94D60f7ZhMHqEySm4Umt4oo
lmU2fU2PqF6y7BDIVzwAE9U0Tute4yxIIuplAFTywps/6ejqBHKWgIAn5KjVPy6t
COZmI1CUvcsQxsa5hzP2KXaiQ+Jv0w24fBWaJB7ombeiXHGaysZOh+kia8lkryq0
ScFxZnFOPOpYDio4oBCCRVQXMVZdnfTwV1LZZnCjTKTql9EszCtdn65EjuylirsJ
CTsaKfWk4coDR8hTUWRczjLMMnjn1LPQxMfcZtSOs+6QyEy9yo3r6UUQ5Ppsdsw5
M4cUtoHKOS9dQerg+NO0Fdf1an+33iOOXK4e/ki5QODBEPVOX1UVpN9SZ4W2gQVJ
5KuIqfzj+zBiARM5z/JH+37CNijszeGFpZ3SgMkE4Q0uMhf+UT1MQWy7aj6bYAmD
chC/QjubfOeqplNNAoeg2YIWrMmHxjlrGTmErvctSEbIa5ths4YHQ76ygFSv5EcX
DbCL7yteAM4NJm0/nb9Xb/oBqVapNR51I53ndE4BLh7hCZhGhHMw4ONNVOuRfNrm
u/sWWpwyJZwYoyq1Ms9X8wWcmsxXmzDNjDTX7LvigPbkBtvtTVt76FpQvHBZhHDt
BNjgSop93dUPUXgj/TmQ2nNGPA8CXhNJLwEJSVua0MJXsVIarpYAxOmtttA+iHe4
N6TBfwj7moVOkSla65CR0GhdTGW47vn3VfyXso/isKPmgzNOsyBEZ3vILM+z8cKF
P0ErPcgWdCVBSFXODyBtSFD3VNjX8ROzay0emuwnCf/BA1Ey2u94aZFgSRIpv4RP
MDZdZX5N0QjUtdOQ3JaoQunRbJqihuosEvHtSVCIpl1xIAG94AMATGpHVdCaCctX
`protect END_PROTECTED
