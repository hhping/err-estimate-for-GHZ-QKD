`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TcJEUAefnl4tT704TqxHR/gPIsSM2q9rAIQo7eit+tOTqCLxUWWSxqBzdtgsA0EK
///37TiCHR6ptXTxUVbYbokc+Sa45bZhd3TSf30F8kUmYGcmV8FGplSSoWni0EZ1
fRTebtl9A2ZK4ncnFwSykrHDAs15y2oHAN2/nckIUvpvOdy55NEX6IDMRHb3Cza6
xHVRotITp2ItGPYmASf40tK3tDkG+xfAHXehLdKNuunN0f6UklJBAWo6I4nr3e6t
+eOdjd4JWwyyFrpHogt6OKme2yjaE3HymUd9pElr6S44oMLd7W+34EqH/1RhZciN
lpKu6jjY+OgKLzpw3/E6YLIGYDk/aQWBtEjOZE4LRiHXwS00uVBP3++c7en4TWuE
dSo5P8TG1bf79ij016+/8lc1U7O7JTpB4/GgG99NxcRejsJX/OSMIkSjacrkshGP
b0tBfNBvD9yFWsbe5FBF2pBQUHrviffJdi74l+e8d4xLWv+/0RV01kSlP6v9toge
mD9/2kBt9va5qyXYrRSUgHatewXlWoaJ8wHQ11LJ6ediwyPA6GmqeDCseLh7TSdb
cJR153ipDhTr9ddzleYkpx56ouUlQTN3iKwkA4Ipz9IiUXYFT5F/I/JvJfyS9/Av
fQqFidUOd0Hfq3Av/15Y/Cu9Yby8vomVGN8TghlDMAc=
`protect END_PROTECTED
