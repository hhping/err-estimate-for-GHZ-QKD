`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZbGVAS7yj6rs1QKhEp2+tBgrWDHONQMjhwNBjNV3lx8wCoKqXL8k2ELquYjGtB6
1eyB2Idk3MD0oc0rShnAE4bytEv/z+gdi4TyGMeoDzxgYSiNVJ3j+xyMgzdg6sTD
e46ycwAVyKLTqISyFyfG3EayAtx1FQ2/6yrthJtQnuIwSzVJTBQiokm3FGEr2cKv
+B/i3p8XZ9w4TnYLMrxzFnyCOc7l7M70OzEgYzGk3PsR72RDII+u+HeQ6B97ESD9
6zKxPuDr3fdCLanNiE9dJC2qv8FZMGEP1RCKcvOLEj3cSjvekTKRcfKoE144kLN8
pK3UnuaB1m0D/nLL3vUcjizmzt8Ga1X71XAothkG1nuJHmkGLMBmOPIcSjyG2z6w
Z3x0t0DWQStvc65oREVHqw==
`protect END_PROTECTED
