`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knavFBeOO+QkwsdU3kW0nmZXxXcz6QzjUGVq0Tfq/+sFinSxCOsMLJe4/x8E1sUA
WP241abGSSxgje9EZktlnaxX/rCbSAmjkWHC6YIzHjO0DONETWNiP0ublJ+ZG4Cp
4oRGjIgkwJzvfadENYgi1XtwqiV4KmhNqyTC3mcZLm04BDtNA7K7X5WdqPvO7KBu
+EmnejhbtRlnSq3QNJJgf7Hjiz2OLJr9tKgUjYWYKlefKNGDnt/YfWQkiP1f+P63
oNM2qJPXukHTZQaTBf8l/MQggCUGSPjzwqqGUimkl2YuaWt4Ly/XS1NkDTTqg4d9
pOyT2g4N3DH0zpftbruowRBq4JUiQJOzZJ5fFcFmLpG7HmFa12yL7/zOMHqUK1Lr
kSOs3laPwkqOvg9Jk/gkakoN3i0OSVgjnRVth9l37bArZ+Afeef5d3TswbZhZQSJ
X+tVOJriUr8qGFNd69nvtZjqe+RcUqpQGiC8DlOMplzCjLQG6Hcp64YyNUOVpNXX
MhmVjR+1d1u/ls0vOqjCVKCwRBR64INyIelZVq8wfVSsSTDU/BXFvgAe+7fEqd5/
HXhKbQO/nlCZfKqHo6bsDWmF7L+rZyybuFvlYl3teqYmGYysLfSALwWagC0ZAb9R
0dOv/86DNSYWAD/BLZEAGnUD8x13tAHOv2nhQKiJ/F1rK5W/0i87qSxAkkSEg5/1
menpm8lW7LIjFJqx/qBDVmO5JhqgjTb2hK5WwWbF50EkR2zwEflxF40NLG4OTtxA
p2gKQFydTlZgQ/epT22WHyXTZXjkRgguJz6rpBWgMF0zJORJV4OT+6Pkd/gd+pw6
wX9Aw9wbf/tpQPuAjwMiR036Vdqv6y+aTb4kHLtykDq4z8aekqZuDNg3studCHua
k3N12CROgAGYZA2HLFmgl3z0xSOrKn+dBbFdre2jxEYuGLBlgTAIQJ7BdClw/kga
NmmtcT+kukIQ1fdjypJGidyF5Qi/imyMbgHS6QRMiUwEm5DCWtnkjEhFB4c9mDMX
26zRhoQs64yw9DgtE4/jFBL1lE9tf0xwVW8tYfr4GmrclW8c9kHa1vIxR7724Tfx
kVUFHvla9xlgd/+pOkokyrXjoawnkc32ifVnXlgAcwIANDbrCbieWqycD3wkvqwz
`protect END_PROTECTED
