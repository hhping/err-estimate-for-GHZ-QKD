`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6Rhj74zh4Ly4Z4NPiK38BWjwHiXELca6cNX+gXWHO7SRbLL3FacDQ56flpY3uxg
DAh0s0QWOtHFjHn3CPE6s5nkajfxDzqO9n6llk7mhOWkmpCpEnxZa+oGFvVaexIM
StgInNcjt//I8Ojkhr32+RxF/v/2pur0CqLoPB2rCumR+DQxh/MJJy5Ta/5Y8TgU
VlgMKM3wyNQ1kIj6+w2uoxeI4yl+bEAf/d7n3XW/mU7sBH8PyAN7CQudiymMOywm
rJ1/PN2hFlCHaxqurCHxGEd+4w3MF8iySPNtvOf6HuX3rTMTGM210LMP8cRj7IzM
ouY5JRRjkOW8LK5l/U67hY2U9FlMKadyY8dPpNYy7bt4u2hQfOvEHk5Jd/H1ymCU
Lk/ybKEklsXwMgubpSWnmfPNSKyQO67sgEUT0z7V4YdnyXxTu4a32cEs827vu8ui
2dBAVM7kLPLiRpoGSNdIQcggCall6L8q8CoG+ieW54lSjki23kdq/zkXUgtNvbuX
2eU7klqGj5UCejlllbmOP20RnP/dRXem0fjrVvf6pldeKTCa5dLYHEb1Mxpyonwn
DpYMQ/sBB1EE9HVKk5I4GvRmZqK00RAVp0xscNxgMj2/gU7YudCbJggUEqWuSqPp
P9HkJjxGiZutq94BjHx52Mm2SfbX7y5V9yYk0sUIAKBVBg3CGPI23JyLPA1QBuEs
tMaJAW0Ec3v359z/y6DRXw==
`protect END_PROTECTED
