`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DrBn5ptBZ2/gKfz5NIywQMnNCJrCxPI1p6hZKniBcLeP0h3YS/mKCdJyG2NZBSP
ZTz2qvDpcCvLfQ6Jz6BM0zn0K/U6GCZmf39zE9wVDc9okG9+WfK0PQOgw/qt7IYM
51ruboYW7X0YRokghMDptfT1oSGgpQ1Al5TPQx3IPA+/c4xrMqX013M2EuEW2Tf0
gG9R+V7uU3mtjNsYSHFA5qPcQkw78k+hjJX3cyqfIQaiO6vtPSceeWPgDSOlHuH4
VGYMaGISRO8sLBRus7x3lA5lXSfBRKd0CcV+dVDI81QEMB0SQqgdb83leNTWp70k
ucAVZ18fIT9A4HqJpZGI9Tney+uoKhPRO40TNSumEx2VM/h7XiGqvu2tcorZ172S
MOY+wy1NinrHtAPTT86+xnKWEnQwbWZDVcVQzvachvSEqQm+0od1ByiLzMiF//dX
89YD12IkzVSIvRJQbhTRgyZP+xk2CkHjkgi07CIOSdc2o0/Sma1m/N0fSgIyezg3
hlOM08csvECEDqvosLKCgx4SMVgLE6kBuvhEAgRjOtyxmPcEo1eRtZGmIwNjb24t
QHVQ+mgQHYchE439pDMVk9QhWUbEG/0xfL9XZHvrgPVHZnhdAf9rPJztQe+wUCjz
`protect END_PROTECTED
