`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTOYCe+cKlCK5VXpZ1sYqmd9CotAFFfem+QNarQkbQM0vNCACl6iFHEKUGbbuMVq
TyL8gwqrMCv1SQaXvdNDyceFROA5VqelMjdS9L/l285h+pkMvp2ivYnS2HTyJ4NR
ynt/B0KOCX59UezMQB+NdH3XC9eizMxdzfCyvREPyBDTNWfmFTMGq+Hv0PICxT6+
vILQLsrmODhxCJCqZAt9uC3QTVYqLBk9PPhVNYls0Agpk6cqIWWNrgIsrEZB819a
tglqI62DPOMOuO0R4PwIpz5POtuObJJpHfKpGH8T0vXhXi6HYCSKnlbyii0jaIEo
w5bxlaclayqf1wwqo0XQrgS68xKloiC5j1DW9a/uQsXJbMulhkRjYTuXXt9Vckuo
wWkHJidPaVmlYT+e9VIEvwNFQghfspLmTaQXNcXATpzjQiRhq/Jo43t6DaqNazmE
A0CCjVlyO2LkQ601+E+wdBnJftUnRShpgoaSND2TnyAZgKbK9ndl3+4PCk4s56uk
`protect END_PROTECTED
