`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thPo5xxUi1qOdb3Th11wm7jgwken5r6HFfjABWHYRS9sTpRgLEOftViKRdu77x3F
vwvTZulpMSczbn8Bd6ususwGWKSkN2NuWGjLWfkbOt69NCklX5upm9unIYqP6U0c
kjhDyCSMg28ckEVrZ8iGs7Mlqpdk3hDKVjehYRPzOhdM+iSwqQ4s29y4o7B6ryV+
rnXy2VNKslg4PULGvZpskQf8q+R8yZmlqPi4VVZ3CQITG/rPgqMyTBMp1XOddl7/
gGaqlwxf43wesUBBD5jpQC+GKVuJT/uWZt5daHspsLdEWp7XM8hbfyE7cbPWu2B0
0U0tvVRRxbtj4kAC1dHXmnVoVyuDkeqeeBqKfyYTwJ8LgBeyZJEXtY4D5IDpVoCD
NbSITG3Ixg+BjbxR7BnMxG++91rK/xhEiu1kRpFCNDCeeIB+qCSdgUSx3b6xPR1q
XnoI13BWBMi5rsqIOb1mATUxKqMmfy5r7/JemypXK5aYUL02ZpC5AiI1OuQjWzzG
qzywZmWd4T2XIVFkfD/6aDO1Y54wh+LFwFV1N+7mhwArD9066p9IhiPz9Fo9A27k
mDZlqUkPh02Zl2sDsb5DKtJNwkk+TgvRn1eQjA6Y0N5nQUluxrFXJKsIJWHBm1gZ
jjfqvGi9DrRSpt757H4n66L2PlGkVf8bUFHX+KZBH03PLnABG85sfvgwc9g/+P1f
lDJs+3PxhUE4MJxkLbs1hU+VW5GTvw+nVzbcyBBK/cUjEcdumniY26mNEwOzQqcT
/DESd0pbEazODQFGtW9k1ceaatELrjk1RYe7RZ5/UTtUplp1wdX2KnsrUFESV0wq
+Ts7yuBufzICEvYQRFqcZPnNYDkuiUHut8Wkrl5IAyqL34eRzYGoWVPGH3sERhLl
q6B3ZE9J+Aw9XPgJEOXFD5EGTXKUf60qdtUPLQFhUWGsomqeTTEuIX7b7vNfzV7o
i2gi4Ja8y7Ky19UXYaIrZclY72DCzcGtECnGMMddQPogMIhvWpLjHkJUOCblh67F
1Ps5J/bw2uXtUgGJa0Fe0iu9xuPtMGUAKxFJoBOUfyCyoAcfVAbyvAQ/Iz1JvgTp
X67Ex1Rt3OMsWKJ+WFChbu8CUj5EFVaj+2h3B6Kv6CKTRriSbBrjuY36L4SHQpNN
Iq9Bq6wwRU+/K1RjOaaKe5BeFHRytGT5CP8Fl2gNs4g7v5tUtMziestb+5Bd+T0U
T/T1pdUxNdYQqTL3W7ybo3peinLDztq9iLjDWUo8NouIoi7mbGTjc9JF5moFsxgW
1FH0BmB9BdV1NSAUx3+qkB6yhFj7t5M1O3XQCntZ7rmhS0t4H0WfPc2d3qI9/kg4
la27PV6F4Xxfa0cD5u/S8jqwB7TTVs8nxc+nDsP5a06P/NGa+paQoR3feLv7UU2r
8ZBwiyxvn4O9O3bC7ypPpbu8ywDR/0+rG6guhwFzOUZZr150jyKXc2vz4eZ2flYF
on4174NwTBvTkFEvDdS5JtGBL+KhNYFB+xl77+A5+9X4SmwxWCYil9Eg0LEv31jN
MQ7n0+MAbWpAA8tw/2RkYSr3N2GvljzXZLmmllfaPUcCueGGz5rrtieX+lThWqsL
otpJQ7Nm+kB9k8H34tqruiCEQWnBhHtRnNNGrXUcyo1qI/NylS4zvRFyw46SnPeX
welTHs7alBTTCjrHV8sNlRvLGRR9LPpnpOxjaVuYY4LweCExEuaTrHT7NXU/l1dN
LdpD4Adp2jZbOdSGpFGZ5QsC59fq11eGEO5EIxyBAmbarIgz+0Dg+a/sjQBEBSIj
2qZVVUF0kyQZoeZi1W8MFHeBN6ewUntdpxoGYcTkPdnGHc1ZoUvjeOmcpvZuzek2
0EdMxn3qcym7d3cqJN4lA7orRbkt9N1mb2ey/WanoXPDWvtdoWa97eiXrFEJCpPi
R+F/tWSq7T+cmC2utHa0xzqQIKZ0ZITi9Tf4tLz8h4yY336KGmf+N01/df8tVt8F
j5QUj1ds42oK9BAgQdnaSOn0swwFZDNK2Itow5Prj+6/N1Kh8LrSaP7uvbujjBUW
gdyjHJOBa+52xn3HEYfB+f7IDhsXoRX9wbvEZxxzA44+fyqoeKn2f7de2VVEpVps
yWSDLPVEedj8pL/f0XxnAjKV4ExD1kscX78wYjoRXMOKN2Wf6UZui+G6x9NwI1QO
VFk5qAxIqENKzbCx7pmr4w==
`protect END_PROTECTED
