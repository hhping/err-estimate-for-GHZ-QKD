`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvYbqHCmclwQ2FgE7eM+oVImL8QcGnlM12XNDCxqsjs5lQY6WiZ3qSEiw1L0GEdp
tqyIccU48O7Mq5nrgH8Wz8P0S2MA3SLRBLZOJ6o1B15kFs+6ezRKeRdLH23MLpNr
0ArIVljCq9hpNIwNXFvEebGY8Wqt1HqK9Mg3nJ+p4VbAzBZPUfzxa8fq8e7LRYvY
kaBqTU4MlPediZNwC4V0Yuz+Ch6d69MOU/3Jsejo26rgX02w0bNnrSAC3HcnWE0O
yzlk9MYW8S/4ZYQIgjOoHdyGyJlms4KGPfzmadEFYUH6FPkNWuPk8uX9C2SVI/OY
j9oQhne0Eiz3ABvfWWmbyRio6S35898KQ4WjdI+S2aInOO2MVxruVeMquF43bBQ+
jua8RWfodyQjBw2NMHhvqWKGIThEw3vb+uWeS1o8mO+vWOCbHIOqQYftJ3WB4cIE
QsnejmGktMs3LqjcDYUYyWHqbxWM+QlQzMe+seKN8Ya3tOP41C14YbZ33fYfrROi
ZrXTXZuRytd8dN/S0sJCHjnuO4YnV6LrAdjRGuBUqhHj4tLPf+th34K89g4FKiLe
EXId/9Zn8Ie0fAxXnpKNKnzOtt1zR3m16fcprtuvMqc=
`protect END_PROTECTED
