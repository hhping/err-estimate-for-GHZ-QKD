`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y9ViSCtJGQ/9EoFZnmoyL+X7CA7r4c9kRfZnDq4fpQyAjI/IJatO9gsonkygLsGR
teiSn9CstPQarYmlpzef9bFXE9f5Dr9XzOLMQnbx6SGxRg36g2quMj4rwCPASuu/
tJ6PcZ4nduAugVcLGEtLqc+/AZY4s9mIgs+LBSyrYk5jv3anTUGgLUf/5qfjdBV0
8x3lkdSSvxRHSXC2SNpHPGC4kkSH0qJSYlYTIxLZLWnxE1Wkt6oldBRnIMWMVoXn
VgvqH0yDcrzX34GLe0lzIzoNLMTWbdRCKtv6pDkpZjy8uxTcdhEMM/Ary9tiS0OY
+IO2pXmmHqYzqBuODqUww6Kydmsf3s3YHrTHxksy+0Pqe5rR+thA6+rma37I+hQS
X4vE+ujA+O48kp7OkptnBp5rvFHmPtH3l6exgPycupghsA/fBqzPrPgcS8CipLDS
wNbSw/szNWGxLR8F8Ri2EWck/ls+bere/fMPqb0pyCq+OP2ESnNi3Ku8FyIkPfWf
yEQtZpe8rmWEgckA70QeLmGz1Mxz3GjCMLrER306CUhwsbF1NM0loefV+QzfrpO1
7c75gjimNYV0M19JvqpSeLajUwWw27AtkUwmR5rrrpDlWJ+chOHvHJctwbK2+mLI
idHMJ0MOY+CHCbE/gZ0oDIiyDwLuT6nmAC3UzdpEXGECQk9RoW3WdtI0egFZR9to
jhs0Pdgn7k5EDHwptrF+ITXv6HXpduZSxkyGCmfqDoUY1kdTlgvMRZEk9exj9bz3
lXuWuO4gmvy2P0KwGN5/dzlciHzMlOnZ64LbHEDT04BQZh+v2ViwLJZ0H8y1775a
u2wZV4Jim6ggriB5G7Evc1SZQqM4PtyC7pqDkXqp6zsjwkfDPJPGeXHxe4QyEjAo
z9HpRfTBa6gmGRXF4Rv1RKnAnCb+F+Cw3IE+Gt0K0bwzXDB7QPaMCsG+JHDIz5zX
OLuotOpsbp0fW4CgFF0tUCtqjvcvoV+7NS4/Ar5jUFweIgvQjpF68uGlaVhw/wXe
7foBDO7RRhwQwTotVInqyL0d1FGdx0XajcSOBoIzW+3zGLkWQ0PfVXHoVCQCAv9m
YKd15VXHIWiPatf8+tPwuQ/HTClnzBpQb1y9sbuOim4n9Y349XgmzvCA7jo4NFIR
GqeDu8A8uGXzEzIpetFvTZ8DaR6L+ZMYmaiaeCzwNh90D0WJP4ds1qKZ8yAbf6dO
GCmuUWcpyH3tfDcH1PuQgQQgIITQflkzMPVMv1s170Q=
`protect END_PROTECTED
