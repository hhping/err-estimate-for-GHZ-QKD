`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QXDeD9wuNNxaNkhaWyNUsP0M1HQDfPQKu1ARQDMjQkpC6ib3i1edY4iibuo7Q2fL
7sjC/Les8vOqK+8217K5+6p36Z2XVh3fL1f/NiTaY6lGvzw9MzQzYiOd09JmO8tw
2YBHKjgN0h3lY7w/UnLbzaNRH+uwakjlecFSvwviYLZYobuULbkIOso0XaBDv1To
8X4ObnPBCCTrU+dT2t5AgQQd3BRYlu+MDQA9RemffuZ9MY2UjC3CJnFyP168EyTd
wL7NcIgaElTo21wC/R0UDFNwRHbWOaAiElOjoZT6zNAYF5JtlzkdAm9yZFbmLovd
RZKBnZVb5MJOHWK+Y185ehWQENYKB2yr15f+rQesC+8upX3kldwqEacbbR9CAG7A
5Ls/N1XoD40/qXetzTMdIF1x0+9S7zN7Y/+xg7sb0uQX41TTYhFzwNO6k9qUzOPu
PE+yGsm+TshSnPC8/720bUbh7IS9DEQcGjBWvrfM99T6o/37BRFlQoqHqmRdp4W8
FG5D09hgnMG1A/I4YIn2nFCzuxqmVnecjWB8+0gBrAGBRb7SC1bQA2L0q+PM4fwM
`protect END_PROTECTED
