`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WIv/Yw3GQeofzQq+uRxDatYsuDfKeVOwnbO+NnJ5mOljmBsZmkLWcb7NgjtQDxhM
kO27wpTWnxdejdpu71Nh7XTGBfbG4O9uPAm6VGBRJxyhfiHilxT4Gm6vsfg6xcA2
535LzBzsQgLLXDJnXGi92yUwkrlMhCGFZM3dNXl/XO1UvzHOJvbxiD6ruCWRVhyC
WrVCCkrpAJaZm7dL13vz38i3BzyGQub7nN6i+kuPql4rBXesHei+/lj0BFmGn1Vu
RomvCuQTrqdRRyZLBsKwMWgNyxoEphGHGOB3h6zNJ5/2BLuZaxyqjtBsyKW7Qu1t
VPm+1LbN8K16IiSKrymD5m9SI+EmDoiomecsJr+1B0g/F+2/I02tWE3rCT//yksa
PMeL242Ce5rOwox2CyQ7b2jtCE0tB9vMInuXmZDAx1snq7JtvvW+AQnX+lK9LgUQ
bPBMEETkcwNujQlworDDJCESDZV0Z4D4FrAjaBTv/cApDtm6s21sGr0BVtnHgO6Y
nHY6YmGh6sL7tRRSdQA5HYNIAsa5Gw6Bp+YNrmJK32r6yn7bHlTfDPj5B0h0p/Ft
6pr4XORN1QTaW6qdZ8+sloJZBt31Nae2buDRBFs9wRWZDzY7FuS3AxlkzRidTPEX
XbcWMM8tdaJ2EGAS3ZK6+8iYTgc6/NXES1G+8rxY3Q3MeRUUECg2Q3IAVdLrmUkC
wTVooDfWiYxmqsVe4w1n94vjAnVhMGft1pIA6+7V15vw0Vj8sEyeBYrXHfKS1bTF
xk+ylkv+DyPQfXr88Ius7v6U5TggEiuZTikeTM62z+JRL5zRkEnGSJZqUlYGF5Ux
Xg4cmn6jpksiMozftfwiM5N9Q8zVeTnMpA+TfTXZYz1UZriImykifeakCEVRp5Su
puswlo0Qv1pwSMz7NuM1lTu7/py9m5qxF4WY/FehS/Ut9Wxv0abKrnUNGLRJ5PYL
z1MNCB4z5Tj4D9bbVybK0hzgHaFVvAuNcZkGuTx+wYaDkUlkttu7FkXj+XDuMxvA
v+Y4skAOuBm9UlMewtZvHnviHR1tBDHTySZEc3JwKiU=
`protect END_PROTECTED
