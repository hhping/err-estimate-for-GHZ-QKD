`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eb5+6rd6sWKMylDcnz1C4uyaHnPous5XIOsvpl5NtasAgQCc9DyzUq92dKYHjHdY
HMpyH5mnIcp0o3VHJnVjsaZHfHm+DGNVUr10L3nAn/p3nfTUGU9U1qpFidLHz3Q4
ou/o57Yi3Ve32Ru0wtmLbb+ILRAnBVLtMjUmxubB2NERDDJhuQoLCFz58XhIA0BP
vQEH74j7og6F2JXLT7s6FwvZncADwWNZ8lYxhXyr//VyltWTArMIzDhu6RMNm+rN
OhJVzr7eZkH3KEoZWV3APBLdkZY1LWwCmuLRRQdLD1VlqShNBUTdtEzsTsA91euq
qMMFLZ/kYPKPFbJ+AdA4SiaBCyfpXBd6qIf3WeBWu9G8GpVkUH90XwufXHrcG+WU
bTI7aOZPOjwKcL+vBpPGzvHYbrAouZpbuR/3V3mLOmrkLwkpJ9PRrbyBXDBJz/fM
fz/hXF0jU1yZFLkb7+88PwEu+bOWErCZ3WUSGUYgn6ZUbZzeG/LD4tfIBpjUw9Ni
mbdmNiys76g0vO05GgcHGysBw4xFtpDG5AAGVl1j1F8NaVf9NPB6cbO0EWOUwtxM
d4StZhgada0jldtRVA0Y9tUn9NOypK4dXHETf2B2JQxQwLtrxrrSQZY7tcfJDILX
M19OUyiTcQ2qiPmfmeJaad4S994hRWXMESd3uG5yrgjEvTQX/1RibF94uMuDREUE
`protect END_PROTECTED
