`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OejJk/2qTIhs3zG1aC8djfwOcagEXBL5oR90W9D2h/TI2Uxm1k/0AIRRfnw1PA7q
vxe97J2dgNUqyxkNH/dRqyrAULVHHcfmM3Sh4JZQ3fPX1DlI4Whk9gdYEQ9nF/nB
PZDVkIP4k/FzcLpH1YEWrirYmjgkNm7nK1u37xzeWck7sLcp/MLNBct1Z4F3zKLy
sgBajR/2wrKTSSXYayYXAq1trSwDf1lV+m4xgEitWlT+1qwmZYIk1igtpINJzwbf
m1zODITeZniVUiQ/CNYmTVfPvhzT2BhwvFC3gRQJ7nSypnFNEWpQk8cSOUPWd07l
+RK0Bt6lF/osxdfTJbx9qR3kI4JiHLm3JTGJpNlOXGU+XlTIoN/I/45/l9gpfGqy
ff81WzAAOe75NzjPbJeTU7+3T1KedPv6irPWzj4lg1Q=
`protect END_PROTECTED
