`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqjIfzIKSzeaLMi4pCAEOBFbB6of5HxdeVcb3MGQKuuDoK70QHP8lfWVV6e8QWcR
X5+Up5NkfINRFNAizjTFTa8GtFQI7v+9xd7gKiV07Q7ERkBj9vVv6VQt2bquiNf+
y42kamE5kHNveNLFdo0ZVrpR02UaCIvS4FzvY7hsQ7a6BViIayjrGvxvoUbWnBRN
aSc9zq4LAxlVr4Mq6VJVZZjK4Y6KkbYSWZ9PHDGOz6R1+68mEG3gUSjPDys84dqA
OmDjXZYVGQIfI6c9SP5VXtBCYMbKHHnYZWpfOhIMme32nkFxTlxH8OfnOiwqdbnd
oOU2rZHRgWJeWe5BkjmwimvS/3URNmJ6ibYKMqkUhFtEHk8mfPOyjSt8/6BLHdFz
PtH/XvBfMGblyJ6rm9HpA4LpUmPy2mRJwWocuVXqJusmC71GcsOGP+jgfsQ4M0SU
saYWLmzl9xiM9Ad2x6RTTsHKdYidNYj2LJUqrAnVqBBr380KD0Vil35jCvxZS2yt
KKM73Mr63BZdig1DRgyyjFGp7dq3Yc10ghEgJHnd0sUtPLMHtgiuh96wEsuP/AHo
nOiI3VOMZc+w0cIJr5t8iIh6NufEutQ7oe9kec4hKQy++pBLh3TaurMpuEOTo8KX
24TVbsM8Xri6fNXwk6Z5R4ZsD/Hvw54jZ47pD5DVBH9qkOnd9gg+0HO6Wz3xMXJC
0QJWSnDmPjCx0Elf5Rf9EHvVUATAv/I1hySoZtFJWlJcytCiN4rISyuejnuhh6Rv
11zT4b5+qjNFHkJPJ+BpUKuallmg7EWpvA2jUgI+gd9NH8fH/HR0cSvyI+E3FvDR
XpKraiDjAXbDnZuymlFYC7KSYAboZhcvT/Y/8py92QqbVU71rVPiQWKfwd6HhoLj
2OkNxidtgs8YDmgK4kmD6uLkTeJL2IMqjD6gviFYETq+NIP3zeojk5GUPnvTlTHm
HBsee1oVxTP9nL02/IXtQK6QjRMctydEWkKsjiv+8DdgQMnZRhI02CcNm1vU+Dbe
AueVzvD0zKNgZY+X3NuiRQLtkc30HGcAntprXL1GP0F34Zw6ovCZkHAl+ejEhYTT
Dbv7WvRo+TEBjnpVV/nnJzR1xDoBAqRXjyZ2VeUYxhjCx3TpTCohY4aDH5jTLTW2
zukKuetR2ApUp+3EOJ7101EaKbggVdZ2wcut6i8dUt7QdHA2kuIZ5151ONORvZ+1
UK8gLxNbxDHyuXrFFG0fxJOCsIb9syYcBbVQICbDmVyq1iyi4IdoJ4QuuIxGOagg
SQ261t0qean8IB0tjnNISgZuSzIo1JfAGfuhV5LehBXQwDePUwBwnQ3N5oEJHCAi
0AYblAwOW3fxVfOr0Nogu3dJQUaav/G2KE1YbR5Or91bCwOuyoXdKbdvYxBDFuGr
zZXSc9ozTd7hMcfN8mJ4xJhmjmKO7U5R0PKd2WkoH8ikMXGhLaQMurQA3Va4yxJS
2kTv0IbXZbwEFSmgf56MU3SPLTxLJDgFz5eyy8D71A5hlj7PxgaWc5c/QEDM9Ufa
SXtIm21wuJ+dOQaCbzZcHDYrjDmCTxR6y4m3IEmflFcDWmaoa+BvvG5VdsVkIgIc
Wbvd0JdsYErxlB5pQrthnzWNDrizMIy2Pc3criE7ke93onrkpxrnxFoLifnG60cF
57IWYHYtfi3oG9FZHkEDYPHghll0/rQcx2lBuCTbMDJyCMKLp6O6apvGzvcA/E7S
mQOZmj85shrnsfyewrVLEoCtRd4swHk7cNUY4PAmEN0HHjZNVcSGGx/9Ig9Sxouu
8fEwUxqzMj+3pTPd49chcyOn2ZRWI7Mx4/dnl1HbpwyDZVIS9XeyO4yQuANqVBnJ
xuZ8HTrmDfIaqzYfkT9hCtQPCx2rircvKg+cBqGNL0oo1L9vBTbpEyZMKoeXdeqK
wgQ01ZrBgAF6IfSaDucInbPJxC6It7p8L4thqD+rzpkL0x36lQcIX+WjZ3KgERvi
Pi/rrG1qFHiHOMZylKzlSbBYEiAKygTxy9mFcyBK6lJuL/WfHqoy4SIf70Lzq9qp
a8nDa/GJV3DOkmE71c1CT/iDXPRCSQfVH3FXrq/0GIQ+a2LPGEGz3HPHDZGQ/cds
+Ep8GyL8ZKLx/aw9hiPB0HkqURcMobgGOZz3hDS7EQykjlRnkkFMjzgUkiv9/uEt
SU9z5OWTyybco+LLhJSQj92Z0+Td2fDwRsoxwEnlJaaOoeq/IkCYYLY/hoeBZlgy
MY7bqU/Vd8szPPH0uvRmynVEQwEJk3ASyKRMs9Fn3QdsAF5l+H7/l4F62BwEE6gZ
r+irzckLVbn1Qk3ZNT4RIwa9Y/RNxbf5TeoZBFXLZhGVhvytdchS3jrl+XZz3Lup
j9YsuCQqNSlnjT1mMDAc40IGSake3fnMkOVmXPXjQoGhTyHoQqT+luR6wC2SRvTr
W23FYJKFydike6v0HmYEnzr8n00kfv5cylpunaiHw2A0qyDGqJA51GoYvCUA3kcU
CflzcCwk1qeJeRlnyHD8rFSEHaLjb/MDNhH2w/dC6r0uxEUmZOZx973j4xoxcKWf
Z1zuxlmW/t/Z4PAFmgIkjtJO8Bu8a/bIBv3XoT9pY8tGlHh82fjzxuiXalqEbzfI
/qd+DNbJ8RoKvIjKufjdDAhlCKS1RyPZd3zzAqHe4jCPORv/KZaaGt4ECNgIiaqx
9Jw5hApbNpRFbMpGp87zZCdA0BX6euk/FzeI+LQaz8dz3MiFJw/7VUkBXPRkGb6b
QKzPm7PvbU/tCOtPUBuY5fMJNHH4nAQjukMcHPUo9ofQCaRYi+VRuVkOjeyqHFd+
ED84EctnoiUw3LqZ4GW+y/+xu2zt9DMqU7qIIiH7qsbKO92DuEUEam2ptgU8aqCn
DVDvh7goMl6yJoEfrYmG/s3aTMVQsYlH1ugecfDZELiAGuVCzz+E7QkbOfmO9Cd4
aFa7FYiwoayGasASp4TdoKdB/g1kVTgRApVBy0zQgLG8wEPjv2mvdGrCEdZhgP6u
Z5ScF3KVYwAzAGzSwGXVV4+A9IsAbMNqaNoJ05Y32d9tfldra8MW6Eo+tPbMHpPN
MdjT9smNSAWtz1eLAZduJIIqyoyv1yj53WICk6D6n6eoYwzJmXrnADYXoLgB/Rgp
tRvE1Arpny4NEul6/V+CqS4unnzkE7u7WHweyiV7uuG0LTZBFozH9Xl20Ll3QVNR
ekBRJdqSS/E6j02XHgPJBWbtI3vpzy5MiHUAw4QwyRnAUGGkBX2hk0q+/QLiFNyQ
JD783USHwUxjbIVl7BVDgQsjFWzsmiaorcZCHHMbNyxhpF4Iku+w1PeUzFcSTocH
`protect END_PROTECTED
