`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yb33n3W37VNWl4XW/UF/4JtMZehp02lxIgSsTOo0zBYGz83TbOE6qkQBGU+z54n
eWaIvMk09in8Okd89hmILj1cfSz25mwCe3RDMiIkmN1jrg7OoKNPnuUoKyH+E8c5
/oHTvXTpOyvqBx22b942cpZpTIlKm58TYEaZT+2BgydOTzUw09e+rttpumzBBSyp
UcgKusdRLvP7Appz8LJbZRMkHmnhZJAB3kaKzNaftjgvB2GTatmZ+Wn3O+9bS71Z
qdVM/YHF4rm2CoDSZzbONbvLdwaJ38glt8SQF0Mxq1D7KVGzS1ybCc7igKQAJd9n
EhiwvRO5Vt2htVS12TpLqwW2RU5IolnmezkIlwBFeM/Re9/h5ciunGmsAxBsoma/
gvo1TbE8IjHARuvE/6as/Ez/ZUit00CwpAyN/OF0QjB+49Qt6KiuwH2LgXIGPXv4
5Be5GgaIljhnuk78LVN16/iIHTZ6iRCD9OfIZS0FCjpjBxRL4h99RLa8Zm6m7Iu9
SWIYs3lTaMIYou06xayFe/fmvXPVrq3tWGw3wKbx7h7pG2ri+FE62WRx9HbCcV+m
K+HmkW6h0/Aeq2l6jD6DMSfU6zr3Iglp4eeUx7BrJaxFRb7FDS5/jL3AJJNycRGa
QvBjkVUGckqf1ICR4Cm6fxDECs1VrZcXcpwh+iB5PGQA+ebSLBVlZG5r1F5Q3VgI
s1zP5x8/vey5mKvWZFVdIYpJG9mopI7vSZn/sT1mg0qY8EC8mV3dtArqnKNzwm6R
IsMKkGUq4i+oYHRenZnvYEHqHIHgY6E9s0X3YbEfpyh+S6pECSZI8pJv8eCukHus
MnuDYLreKlPVM0X5vJHClItFdOg4ZM0vrqSf2VhRYB1oQN3qT8DcUXw0klXwAvKs
U2itmULIe2srjxnhKMRxbkNzQC5yUmJCa1hj/+Qa6H/B+V6bxUH5mvHLlQytDH9l
ltlf/fOAGGDiRgV+itkJgIjq3WrOIOC5qD+2Pc5M7PmKsBsn5sqI7s4vmz9MIYtE
c6ausdvKdxiTmj0DtO3eWp/wJmeSgGs39n0AuIsM/e3c868ow1NhhPeueNYjs3OS
6E40Jxx+BGe2nyZV+R4P73RqXUEkRcigE6J93lid3QuCblXPDE0hEmLViQdZu/nc
NQm4wP5zfVdRNnIxRn74mIhQLgnLj9Enftjn2c3bqPMrf5RWgDGDpZ8UQh7Hh2C2
rxI0GA4VpG3IbDN3mEdHmRRlDd5Xw5K87l71LggiOF+Q71IaTMk4v/71VKHMhOyW
mSA8nI+xR0Njdey9o9WI6ve8EuHoYB+qAeU9GzXL0Xh0VCV8nyV8uRMuydU/0jUl
hARgBbzief5n6PcOkiNlzxmI4m/L3THFUcaPAGLcXcyFUQy2OpyUy/+lC2gA/X7N
FrukBq3AUiSdaXVFpzyE1sLMyRHQnGQ7XnBJ7DVnEjWhu3Tgo7S7tWqhqwKAuChF
9dy0ya5cu0PBjCbvi46ij5/SHnMBW6I75FDYSoHY8GufyGl62vVLLoSvvv2I00AU
a989kwniTFA4hfSeTbSYjVXf3gBzmcUwGbh+zap14VJfzhxi5BkmrQu2jBj8wmNC
kcbGiBstiCzefoQ6LDo4N0Rzf138tKOSR/P62C5Z4IGqfM+p7NK/RykDYQ0vGzqA
vVfzBTu6WcSyaMnWANT9Bg==
`protect END_PROTECTED
