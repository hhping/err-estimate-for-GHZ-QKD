`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1hPJs2YNJ1wSdVCrBdCajtVg66FuSV2jv8D9Da0NRBzGujHq3LM+yi/uBciC1JK
i+mx5tuDPJpJ2UlL3TJWB0UYFllx9YVysOHlg0b8vwnuHGAx4QGA5uInxSywh0OK
11G3vOr0bqyIH+aKsdS7Q2TEmxPHdoPREhYtRY6MIMK/CU7WwyVA958c+UDJ4wVr
Os1Oa3Se5lf7WfozuPVEHt7HtjkMKcr9r2npT3Ky0MMIr4gjhCLNWMu+Ddp75IpT
EZ6cUZy1oVrbb3bIYNoSEtnb0C5V/RJ99U/WMZh1hqzyVaaq2ZOSZNFT0m2M4pWg
EYdOur26kWRjUToIfIdYWte1MbYF0hDF6rs339a/VFetpab7rh4XNfTX9RAF3c3H
KtFndXDc3x27SeySR+tOHx74vx2PPn2FRl5WUtdL4j8Ljpr6yXY+8MlL0JqigYQu
8PSymeAaGRkZ5HDfXPZzgnqKsrn2EdHLy56iiFlLTS6lfakmVGKU9X2jOjST46GT
7OnavLvqUWpS6zmnZeyVNoMvRZVWIfeIBneQ497ScXiIPQ5C9llTrPmuuix8BNcZ
xSumpK1RWUiI+BbLnNJnwhx5rktKBI1XsImC5+hy5+znO03lH2XgjcjqtTYqXRdx
X5f5+lRbgRUMbGCQdTIKKRMl7PFMVV2mzeKf7I2ZpezlpF9v9Y34NducrbbgJs6f
JOIYlDfyyTNBqds9f8+qIG9Ssg4g+Qx61N+GwLUM7hZ5Sqmqv1/TRz9iVkVV5VPq
OTFJS/pwgLRlvsnyouDFsQTXo5G7z/CCDhNE9T5HXp8D0zNQtpbMMOzibLtYPY5I
Yb3hnyPsbbiBfXwO+TwHKZvmD85cVKiT2vuFk0JguHacaXmOTTeqpsZMwoGx9Qtu
9bIkD95ALXLU25N38Len0xZFWUsvlSHpDZmBYACjGTOIzHl5sjM5UtEISfCRG7AP
EAEwVp6lU6S2JtZOBHwhRmgOTPj9981syjlXB5vmGXG3vFkOhVG4t4SrrPorAD4/
DvmkGGxcKJd5ruhipDKXEkGHAWUQtpShQcyeoIC/tSKn74rDElqQ3r/ANmPTew5h
Mn06mDaM/5x6ScnQliq3idttW9bIIS1mweMGhfbwzWzOwLm9YQ+SMNNRdiiR/uFe
nvhd3zgjn5Iuov7r9EzYJIDQs/TeLT3qWZpPGgtK2AIBJHm1XzDf4HhNSCR1uG/C
eSY/u0pfcdxQLs906RZdzEBL0gpfGV8tYG9imcHSnEwhkYEUN0MaO8vlEGzScKLT
UDWdsiujPC0NpQgDxxxYjCsS5MNuTmhBnB69z/39u5rSj3nB+U3FrInNzkhKdldJ
7WBQ2wnmHlQKMCEoAIVtazMCHBu12HtDe5YpyNkqzdFyrhI6p25dxUpQxoj+/Unq
bvXGEb7icC0YLVt5J+rGrEkPf4eg8xq1XtfbotFNh34DtFS7/rZ/2QZP5s+qdIls
QAeXdFNNtn9GqD5GK1TYrSvUaNBJypf2hfrNT05aZu8k/ZCCK3n9BO6crdS/f9ne
AFsWKVGQXcq2jdWi0O6kTwIu4bMAoYXBc/xJGP4hAjSt6W+MfTdP2h08XdLfDRfS
nxpJgeFhrtQI5qjCjhkstFXlxGNYByyx1XVfl3JvygnQB7Mprnm+KY2GGVYJmaon
zWZfGRoktneMYHt01UPOKfCdIQXd7H/yHWTGa2DAFsu3wJ9mE5FlpHJcpa2Clt7G
fUyDS+loczkC8ot4ISMcr1BBAgbAVl0jjHB1N0weVGyN/GPxNOnRvCTCVz2MdbiO
bgN6uWlsLgj9y0vJqN5pBIrORnyT+pM41ywk0NZfB/4FoCCfaYt9kSvgNm7X10k4
XqrYblaj+kEfvhSyQk1JadJuLtKwseqJJtmQBPy3Ii1l3O7cksRQ1p0r+hEEvk7l
fGC1B7W3YPyAnCXnrskeBCTed3KM1SJVKVuS8NbVlTlJetYp4TLJqigWU6wLC8Dh
ngbzpmd8+fv+JobCqQMsGg92su54Prie4wpeiMCF8kpKmGhzDgqJkSszmTE/N7Hs
iEIoO30kvwInjB3yKZpHVUL5HujtOeR8CiR5B0eFFDDPXLuw/I7QQDNa9SGDrBLl
oMmU6GJuQhJPmyi/geODhFt7Zszs0bzLh6CrOnkIL+e428x4/eTpGsKhZ6fW3lqD
HxA4UxIqEgMPBG/QW6Wlx96WCGjVr4IZXlSEw0SZZcv1f7zUwwF99RYuaNZyDjG7
DyVEQabNc9TEvFfHkPQjNDJ+QpPQv/ES7Mt0NX947uZlKptVu4faVtrC1tuhx6o9
hOA7hCJRDhz+dgBWxHoh2lY/0q18R/A/7D8ULP3mfg2hYh0zaldOYxfhOcQ4ff5U
F4KNhaOuz7qVIGJdiTNnwLfaRsNDQkubcMtLRuQMO9EaygUCxfl0lJ/YA3S/C2L6
Rl8GMC7IArCpBLSG1a4/hb5v9k00DXJwPQgVJQCAAdjgrBPenwGeqd6s9Qt4yuOB
s4ZlUulaw2oSk1UYlMOAFTotjgtl3ItyfJh0FiVQmrvZDaxhI781m+FswfNvvNDm
C+9NTACAdMN3eLkccAOd4kA+gN32IA83xMIEXVgWyn+Y2Gv9K+yORnG8KehvrTqf
rsxgISR/FVMpMpdFjFDs5oRk4MTgbZT/uOaIb/jK1chCwdJysc+C98uFmePgYUVp
1ewGA5C8VNGUwEGhQZ7gSj/CDheWox4zboipgKY17xvQnuR0uYhn1IWtTg7AUwBy
V3O/v635E2071GK4lmNAvXfKun4CnEFrGktQQ9NbY5Q2KjYcVG6jC0uiw4tuOyC/
diTa3HGQndJ1dy8+axCLSsgUgD3a1WhiZdpOWe2HpNGf1LSx5HMJd4INWtTL3VK2
4k3LVjqNnpvnzzcanMvtxHNqkuxYd0KNXUucMNqY3nk=
`protect END_PROTECTED
