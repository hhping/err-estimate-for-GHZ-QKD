`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDsjT8jUhjdQsEAEkzaGDYSENAgiXgmZ3/2GQAf3/EZ1uEC93oPoCTYVLwNOtnpj
KYV0g32Pr3tkr2dr61nt4P44SjrLiP54isWipdz4RKGP3zG/Sn8M2sY/VidTSXIH
FLhX5ipUAxE2IBCJ11jor6L6X2pV41n+N7uaTM6gH6e0P3H5Gg3q0q1T77D+8Bwj
yW142QEtpDAuxPpO438+fsBEqX6pya1oTGLy3QdbY3HIs+e2bRTorML368g0h/WO
TSosQ/s0e82Roqqzw28PvUyF/kAq8YibPrZtfwUMZ9Xlrc0pjUln0gVc22Wn73uk
dU9ZnYdB+5JtdXiKkqkwrQLsFTvYyMMZxQ2NCjLVc+v6/PM+oEF1oYuypR8ReDnC
AARNP2v2N8As7NXvC3g56ms9weysSsRzfTSi1srVX1jmFEpXv3U0SJm6h9aSkG5a
`protect END_PROTECTED
