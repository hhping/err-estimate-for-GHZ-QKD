`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B6C/H2OONSGjQAvSY16ckiW+iAvTKyg0APIKwkzp2mYwtNXfSuZyK69qGsM/8YUP
/tsHNsOrg6C/MGA/Naxu9KPvdT4IRiIISqa3LJjWCxOHhvY+mU0ADQZf94KiYp6A
8t9yeFpSaC4Od0Q50SQEViOqnlGe46+zmNvgppEJiRxFXjascCxZ2tbajfwcqOG2
TAdSGYtpDDLmJ5eHrJpOkm/EgfmhkNKFiynUYuPNw8G8foi82E0Ka9TLNs61Idga
CXxkSCFjtbiRhBE3wz35BHNujnc3TVOTURhw9COD2MrFJ7Nes8Ko9D/+8s6i+yJM
BD0yrXkYQxqOmoUiHIEkU2DpPwoLqLRGGZ4IBhJ0+P+xeZ+EEGdcwXHMSMLrm+Bf
/E0a7Zr6iFUB3I9yrBWwCMpyKObcuV4UnPEHwzbD6BSPHN91ceRyfAjlnCF+ijwl
AFfcVW5c5HK8RptQXrNCA/Mp0QEGIIsr9EYlvjP3dQqWGJEqq7xj1jNzioXhgmQg
+2nMBqwuc9AoBliFc5CI9QpcQL3AwwErckbaZ9vsNxOBIdVnb+m2wY5IO/vh7tzc
sk7evYzM2OLYTpBadOPZ/Tx6klpvWG17V0UAHMKKcsuMPZKyDcQUbTNtRJybWDlD
wcA4Oq2iFYjAFgtreqPHrw/UE1v4CdB9zjZ1fkpakNFLC8unP2wn2z3s5NWJw0o+
oqknI4w39xXFepzVgHWQ5XzLNmjcN+AsJnTDSJ9MXqjUO44jXFLsN8htsiV8t1uk
j4JplirXAA0g02NRkgkb29Rft3+3QD1/DgtwTOqIjZv9PU8eCZ5J/ZPXxSu5jcgw
RYEP/trjzQRmEYX0c3/At+aj011+Z0MRxK99pM4h+eJCixdp2exGrrp3OINl8Xso
TT6R0+YdIPkHq+O+GzGp1Dh0mScrsorTeJI2YmdBL01kOlJ+CY+h1dvz11lNHshq
wy8ptcaV/w8WzjbS79m5Tpp+AWm3zcSHFL61Kr/NrnVCiHkrmVA7APxvWBg6DuB7
ODLm29IEdy1fd/WBgXR33iZL+4dRoL+hkUlrz5mABSsQC84OuOgOdpztpPtf4IgM
wcYcFBFZPsIPKDLv3uAG/+AupXmSvszuebz+ZwEXl3ZM+woEbZ5JvQCusIOci4vK
4v1/T8BqnMiPWMsdMBPGI58HOAas2j8vzLHSycLbuEUojowkCvG8jlpEBbXDxg84
YTHDAWAu3hGebQRCex8HhmVGzIItHkkfxAcm09wAWxYPBSIFRMK3IoJPhsAyMoo9
Dm20uCMLo22afS9SeiwSBdGfsXM25yOGYSm+Kur/RS97UXz4l98iK6fzs2TD3GqN
e9rZGU90PUyy7Nm7L8enQ86o02Cs5cHvGeAu67GeIpXgC3oQeJBLSNbZKP+eSbpi
T+F3U8Vw0AN5SqVPqnJ0OSXadLWFgClEIxxaBkzsCeW6VQ50npb+8NjAsBwaZ2na
fPaXZiqGCEbJFvI8s3Ca9dQWd4HDNnjFdqdU1I+a9wJ8w/MBvSqRKmkq+MPJYhbo
cdfnKOKZUCrSVMILtqXVm1tAWj9jw/CxNaH2iATiCmWZHguAcTIBgWzN3B5p09L+
uoxBI921Opuz7O8Lbl+1X0sfAqsXBYwn5XIb/owL01SZJxmeqsapYBIpFfuMNeWW
DwIYcrUDgC4QwBrx/sq8zN5oip8kKhSjYvUx8t7Pd0syvKuKEbjwMnaO4yFwl1F4
1rzcGoIGnHUgOiH4/B1NNUzuYsl60hjgfNxMepYBK7LDK0cWzd9DemwBgFdsykvn
WkQiBO0RZPK0KFyXlXRXe08aR/qPe6wCtuzQ9qPYXSAvXBo9Z6WIhQOzwrSyhGsT
sUl7eqF89dV1O3pT084rgTfL7G7Xb/6VIH8EBcGLrarQ+SXl8f2IrqAfoHYM956L
ThbuZu2QiKbuxlKu9NdWKC7rsoqR8fyyh78pWKosl2v5W/2JJLRTOd8Q+7bHnVUx
KMj1qym98gXgi4e9IsyXDKRgfEpa2VstLHiZXlN7clmQt9qtUqJ8dKZyDL7Sj5Lu
LF9Dvq+kwYk/C+fccZbLzVRErfq005C2277T3vuZLuvo7klaEgacyAFcB/yetldP
lJi0JkhsMSjvDk6j64Txq+4EeTxUPmCY1prj0nc6cqJ5kBht1U3qygYCLesbijXG
+XT8bPwbJNCFybEOL4QASuTlIjn8RtCElw4Uw42dsK8TnUdJgihyikgPMtVQgca0
A/tKWEMSr4zebUJC5HPMNDmMWXr6UNDsMSt3bQ/FzPyGfoaNVWxKbSjT4+mpY1U+
hxQfdVWeJmDQE+pgTIwAm1gj1iduo/PQpYw/8nXZDaYPvFrVrk3x/dAfDsXVZYu8
8ohv9VaOcL6sE6CV5DRXE6Hpne7In6q2wIEEcKkvkYCp2QelLTd2P3cL+EmyhoyU
YsUn3C85DPOoHWoUHwwdJ58/LTtqiT1pFRGy9euB7a5Srcd53X3ww5PM3cReQpjt
zK6ZFvaK9dBpaiXkbXaEhSchvx2ozsZVlQZs9/WHg3uYGYVA7a+PALfWPW6CXWWB
DolRCesifKSnI6qjOM78b7MJ9+MbmDtWSvgLgeQ6xmiiAqmt2/hPs2s5dGbPRfTS
dIhbgEmN6cbjOsiuKsN5m+EhSovrl5mvekFIRBccC51iL7xeaUVpvoPHbLtUCo6D
/PlLjg9GucPICBTRkanV4Abgm2cGQknIEmiikykD/MQpw8OTrr3Q00HJ1bnaUIh0
jOsYICxCcaNiIvR7xVQHUdrbyMfdpdoIT8CPIz4HU+by6Xvinl63omWyN2el01/M
P6BF+6JOXu87b7Zui5RfAXiVS++2zSn0yNwkgm8FFk8NoMXQqh8RtkXgdso5CiOC
aNvywG6v1eM5rNwAwoTHMgSz1wlxybTkYuds/UeRn4CtQwD4ILFMFu3JdjPdIRes
bm+oPVACn4ib1JPkunHbc076P7nGOXHjRw8NTuIrbjWKPOemdh5gdzl1em+Y0zUD
DC4A7KCr0CFTuOEzlFhcGt7htp/BtVix2UIYfTp9EOcWNtWRWcwUIxtf/tbIpvCN
L9fh5bLPt4Vo9CErHrCBLkBcMgwt3rDRWWZsFsRqqAEPYT3VYj5TheeTHMZUOjbb
FCC39aWprELJgYDMIoL5N38n36eFRP5ropcrmR4GeqbVPufI+8fLshdUllLojw23
fBVfCEjHho63mmQQEX/4JjFSlbmSKMQ1LcKI/8QikjtE5NHY+yCD+39bDLAiomrC
xvXntgx7m+0fEWkMLRWgyw62neCILK9We5HKDXjFEnTvNYstrWry38BdrxnrQNE0
JSy11E8XhNl1AnHTjbxeSnQvOmVHXpmxleoRUiRw6FfiYFOtSFqo8K7oyu35osJ1
CrzVncC+mHsgwYS2DqB5qdacoDESINBcBAWSV8sYbAq4m+M5Ugsoasp+FXuq7uq+
jk7kk0gORITjes7w8u8PCtNSSCVqj0rq1m7C3IkfXRohRekaqrP+lBI4XkSvNW4w
r40G3BsOF5+D+txazshqFQPuj0xUqtoCPl4LJflbfAOqcJ3zPtOtifUqBuonkjhj
HSqFM2IgIpMwexXWs7uiM90xVC+y2ivSb0xvpHy641xioElIEIwyWMEvJxnD+0uu
PL9UTpcphHpS353m8+DHFtdDnq6GjtYmLmgW+vevSH91pbxRBxyCXz74zbOrJu8s
+UQQMKv6hlHAL05bZDyqcREqGsMbC8wNOQtD9g0d2IBuxIDh+L5VVRi9/bghu5uJ
5MFohjG2NbgSO9rx+p3ywKHtgdZx4ZERKswmpvKhOKqOTelBPa5CJS6UGCAZqZgS
T8w7cTo++lYhJwaFi+YuBPIPcJaWg31PDkBLBJwRguzrlD7x24aAPSuZeLKFaztm
QK8AqwJMIrRmYWsvE14JRb1vLPZ3ffY7EU84/4bTaUrHnSOXiGcGBhhfoehgovQa
8agDCySanWEI8DSsKQjx+O59bL2VYrWc74zdEulrCZrNKe9YNMKVFeuohpfCqj8A
c2mhU5WaYVp1lcpjaxjBxBsqE83XXSLlMAJ8tFXkq8vw9jkb0C41UbtXhZiwIw8l
Qdinq1UOcSD8WVcBJX0/nKpsxqW+z7obM7qxMAAuZzclqWwwO2xxllA+58VINKAx
xf6OHKvqJdg94WdRffCglv5c+9QJTv7syaG7vXaGouqwZkbAsgeuf019TNRcG4Or
a9r6bne3D2N5dzPy4iQE71zsKQWUnQcc8xsTxaqRyDEb+cankUDSHR2DjEQqJv2A
Dl2Z2xVFI2vnllNSeQFsP2gCPs6CKbnOWONRXg9/2kJt8W9TpjV/bVJ4uHC54EIk
4cEwRUJk61mLADsGFy7a8LzwNEuh46t/fyDT/VZC3AGoge1TqYHAoOUCm+ry+qls
p4C95rkO7PGhTJRa7PsdhOS3Mp3Um1xraTz3OUUK2YEKkGd2PqjixUnYB+Cf2D9Z
/hRBFSmCQrB89ULBD+LVw3bxLR/bltoCxkujPi12A44d5GVbelIu+0KssjGgXWc3
BEeDatrRspU+CdJe1pl2cyf8gYbPYB4eK5PtFsjhzfgJlYVf0lH2r1XMYuuQ/lqs
enm3EeiJJocFUTeBkRtYLxf1LBJj6oGLRsjRcXDrSbmy04LJ7n1auc81l7sLtrgO
Z7/sGWTe00dUTroU25mk27RLKkprRHHeHoKhjxQViFfZUsEExuypqKzQuWSlhNYk
/yUFbX9He1x7i44nACuD7VS+DnmmN3FApEJ8SkmDAZba+b2BDl4FFuqbkanHQqap
BFCUI4BzYu2Ex6FKt4RjsjlxvleQjD4Q34wnGh5+5j4DzA+l6P5g3fGJSs1VqKMB
4ob+xfKERykpcnkoJCHL68EtMJ0VnaqD3HK/ssYEc5vl5K3ZZT/zbrZWVBJ3KOLl
n2aYTxD4KuUvXGPMDLLdwFo70yecpXBBRzszY2DeTbRRORRNdjsGtAiktlSc7R93
CIeyb5qXbKOizrmS9jrG63DuNm6AxXdEBvDT+EsvE9N0vErpqUETwqCwymC1E/2C
Pa2Bxe/P3Ras8k7b02le/mKfso4HrHSEY0pXhOsSUEAqdXMjvDZ9ePRW1HRKbz8D
kzcr7DsossBf6dIvbNLaJn8qdx4t/YaUVoJJrWq7o1sTigwQ4DJrVZM1ZyCEh10S
bLsRd/AKCG2XQLO+yykDULnxIvNlRETxBvSw0bV37G7FWzXD395Uf85B37Zdx1u7
+/WEU4F5A4RbhD4j5Ui+D5KBEd12zhuaSoDe7VJfV0TbdrW6iJLKZmi5I84CNuTN
pXYYQpPFLB0bg/htUTY/eBpseLnmFIDhLSXiJQDz3QpRcgtjLV5bq9DxdNNWZhwP
5u2zEsyVcOPeWgdy42822sdQuLrdS4mRtC+gXx0+87lMcxC3Tg1EAZpXDvN3gyRQ
WBQrAjy8vlBQeUg437MvFnTcDfDgLBOnCJdmdlaYNGArR/qeMF9ct0QwxWm2811a
AvoNhPyVdkZkKAem7HyH4SoELJy57yytVzgwHkVLCYCwjWN8T3Cd6tRtFPXXwvbO
FaxiyYtle/DHoCZ4Y4oVQ291VafGAw32/e4Q/vU6xlMyX1ceniBpv8oWqZjWrT1c
gunNZaN2sFwkxPWGQDBegCddoe+V1BvR/XqqtBpIrMMb260lILNJly4HWdJPYaBd
fa0YWyq/+gJtaVJIijxjEvEshrFOh46f2OzH6iUbv7pn2JT+1NtemEjZpkhb6Wq9
oYm2rwzwZHVgsVEGGAXd6t4IRKhOzmBdUHicPbP6WzvXOnukXByUEhHE2yc/rmy8
IaT+Riaxh3aomtOaz/dcW8/07TTFo7YxSDfYu84pVttIPpB+dRFM/Kuip2nUkNgg
U2D6FUthvIFC9l9p1fMFHqTIFJcV+wDwRj9K0vDFYIs=
`protect END_PROTECTED
