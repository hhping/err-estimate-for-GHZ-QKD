`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvNiaWkcZZQP4tBEhMIvT0Hjy1aB9nek9WCxWToR/CcERBq4Xsic+fWAOQNinNb6
pgeQ1jAhgAmtdEyttAyYGwlFz/Ecpj3B79YX6amVNxXwt6oYOoePoxCb/T+RekE6
RG38B0UZ7IkJGvi61P0BH/IW/BVopnE8HEEuOuCK7wvRVEtgIkQMhyvBgVj3XPOV
U8WgpToNOqlb+UkiIe9CEHLJBsspSkjwFxUbhvged2s+ag2Q/6x7Ai3dvFMpIG0t
k2K/FwDyqEU2h9yo3M+KpvtQr9brQqhElXdNYC/Mm5SiCuCTzWImr3kKE7pif6pz
J09BpdgoliGxA9lqW+Y8KwXXIF7zjvNvQv7W6HpXA0OqYaDEZsjykSrbuG+cxSBf
aw1v6MJ9v4B0aF5036YCr2aqwIGoFsTMYZ645PqmJOsG2m79MyFn8lnQEB0+ZftL
op10ANfgyoAd0tHXFMbJciORIDT0XCcKy3jMTgMYfoQeX/GDBiW/3hfDfHOjWtKq
TbA/d55HZOLRihk9MEmg2QBRx+eE6RNd3YMbrvVsEOHeiMYXplUmhAEYozGb9ynN
Wr8Z2gKtKBtFh+3enCGxg4TabL6hL9xL8UkqQHCUAe1mnkouFA0izYc1krsQH/5l
TZpRWa0KRQHkSH3MOpq2ng==
`protect END_PROTECTED
