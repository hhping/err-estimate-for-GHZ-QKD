`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IsXTon7jvZesn0VERn3BfB4rEPn+l4d1jLb/xWPRbBKoQDw5SROUy9t64DoExc/c
vbuOBYc7Tq7xd55ehjFMW0ZHT88yWycdfjFeapT88YyXlgqvSABOG1eKew+SC8cx
zTlF6YwwWKodZqGYAuv8s7jQCJTxHGChwQOMa3SXGgbA086VWZJ1Uc9SVpHV0c0Q
mweOqqx5MR1ldP6t23kQb9MpGtG06Ew4zgXf1SYvFLV2gXxXtpuonhhm+qYoDwsV
yJG+ylD+o199P0DyIqhuEpqX8NtGI4kKgwXYbht+uVEFBVlFAvlXobh3dLlGjklu
utS7n39irbHzgh/LyosQdMVip4iTs7QpzxXSTSEIOcpkRYQm7Ztar7K9YhG3XWVR
MFdg+EWV8EpmVmlPz1UcESrdhGKhx00LO9BHADs5jevxrAKAK0uh0mDssmRZF/E5
TfjubJjFMIa+fExVGBkdpbN1anlt6g6hzBUk5HTVNjLAs8rLxqwOBnLRuGtvDLwf
We5QZ7X54XKOL5Kz+MEM8KD+2yCTTu3lQbZAhjCwL+IDTk4IkHKIumXvLt2BJJ2H
Zd3ihbiXHRc1RpLOedI1sW68AJO3E1JylKb/9IsiCo6Ba519T5Kbh+r9E84wz8O1
nPPT+/KXf3u7MgLPtB4yEuuYAh+YbKehwe6FMIKK/CUn4uNwEvRFCyJgwLd9GBJN
I5Sh2T2eOoKMqpbXLjy5FfugYgARZJNcAiUF2IAdmDIe1zuTDn4fRorvy5FelYM8
XBcu/sWPAkvMbXbaHUcf0EiP5zzVMxyKcPZrhGOGxSL1GEB3RjKdtBQCwQ5x2Afr
x09Kf9vjVsi/HyZ+L3IdmQ==
`protect END_PROTECTED
