`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
biGSFSjHBupHMlPuIVavKY/oJ5HLwR9lMAleniWH43di3s0zY7LzmrXTZ2cVqrIs
nD7MufNgoihR4VzaIJrKf8pMZSFad7vsWQ3hfIIcYaaVBtWce+lH15oI8KdRC9A0
pJCrogVkHL8OzSkrXzD5wZnrnqRgB/GWlzrepxonyEcxQrXmc+5PlgoYD82BIkWK
EDM/82LHHxfZ7FzWMLWtqXQj5C5qjGAuAoLj7IY8vDPibyr9bIiSkMIXLcYriOWr
JUaii+2ECVTHhp4Y4babQabdC5GtE8r7gAIwGHp5hXgqWHqzl1F6VDRsjX0NVmd/
JJKnnMo1p/SLHjNV5sld0vcYToKjQ4nobB1ewWPOUowTukziekzAH2gIP5kXR76t
23eN783e8UgwVcSyW4LrKMKL2LIoIR3i3JBYwUcxmQ0mQK1SAN+GHu3zB/BRxD6N
ks0U2MtKo0KDrypz52Q+Hgrbcex3Ul/U4t7iRnep9qjOONvlsNFzLnU5d56aqfem
Qx71QZiYNQR3XmOVyrjZQtmSjjuJdctq10rz40PDpSE=
`protect END_PROTECTED
