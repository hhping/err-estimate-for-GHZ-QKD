`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hMuDCsnxA9tCOdF+UJ6OtRAmxYVF/lWG0ACAwmRt9a+HLWsfdDzaC/Ay/N4YHWi
hxEoUyzONYnRaeptqlnUISORSAEbQTTMFjqthC3UuBysr10Ql3EtUcOfrJn+JXOi
9lJ71m93Y0LJ7JlEtJN4pVZkB9nysgoJkPMVEPo4wZxtkueXgY3pVBZaYmJm2Xrj
8f7b3bEgNoSlBaTS03sqWVn7tWcwzHTGYGfcxIhFo1YNg1Z8BaiFsrmej4Ko9tn4
HNWp5FFs0qrGzVR+S5Z6pvWEbcfGKv2qAHizbR7w1AAMjAdmYN4010/G0bGmLs8W
6vcVlfr9vYWPik9vz+aN2bs6we4nHGIWvi22kbdT8p2iO/SjUyN+9Oi0k8dylXqw
TdMV8ESJ4ld/oH68e/aSiXpMKu9ciG/iaFpqNKX7q7HsJVc48UdpsiqpD7d/5WQL
2polEU4hF43SUU539yftqRHmpEcxWRpJa6HDe/vaJdIgxXnD7a5jTyuijI+ffUnd
wXXYLFYnw7IPbAgD2XScYbWfNdUjV4NAMZPeGfroZ1oIz3f5h5+VUKcI+LYoxCSY
8lpK18tea+UhRRFgGduxRLdvAYzQetUd0FbPxHciRcDq9q0WrIMN5ZtCbW9wwVRs
pNfxNn/B+YfKjxuQCLIHfxmjqWPoY7iXzY2OSfJuXynwWj9+jf5UDDjF5yBxDpYz
`protect END_PROTECTED
