`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLA5AeGCu4FuvaViS+9yvhEzPPIQHGPucKx5BcwjrcS/PJEhp78YH3v++aJdHs1w
M8vDYO87MM3/5lF7kx9KR9lZCLbSTY4dd2cQ5XKL0vpYWEcKJnkpSJ7YWW8f1nDZ
a8KaQqvLD/S2IEtSTSujuh0qCRN5c0b1vzXtByDTXU+kNRh9QqmxvhuJg3Wox1K/
tIAXhfozZvddGste/qYOFRRB4mfnxyf6T4a5a1mcmi6S/v1xIepWhU+th9RZyjeO
IPmAjm4MQeBAr047MkfPkcg5LXh/zKlwfL+jgr6beAaAa7hjUWrx4kKpjeAHG86X
6WHqM5fBc/YyLAnxYlv+00frK7oj411mpafHU88CMvIB8Pi5K3RjkhJMwRZvsprU
T1/xsBO4mO/f0hPX5dHtDVSm6IJOA9X0tVXqFQjmKKiTYtH78EPW9BMHqCROpFr/
kCXjzzQmrj96ySFBWJ07LXHYkOTHXb538AqEzEot1+gbn3ks7C3zwC2YMAxQRk0V
7drZIQ1b0B9v2c3cainFsPc54XdyJUM0SOHDr13HAHQvineZAZ9PWrQnzcUNLlbS
0K/IYhUm4lmyJDZcpVAC4nzLfyZVDgO5eZhT0/YC8KKbPInPqfw1vfDKMUDwIbv/
7RK9XlzhTJXNMdZQFHqn7e7X9Mb87yCFvvITqVJs+RYBDsXGDf6532fYhxRhmd2i
YXRSdVUzEp47NiZje+vwkdZLiXbiwSVH8Us7CV4XNA6j2XUDG/YynCGXMztP30+F
1pv+BLNnBQx4wTLFLAZGn5VFYYD36ABHAGSHTdzf3tl8+4/jodAKgl2OhEu5Xy8u
gTr02KgUXW+yyKsrVQbaP0EUNfq/sIFmhg7y+eHxab7Inn7FIx/W/38NjSev0t3W
Rgko0o4HuzAHbIcGDonzUiGrknGUi6eSfsAQa90CTns3T0GYAK/pC1KlzCfCGCMk
1Jjcbhg/AHCvjjh5Nm9KLsvEWXOpD3j4vSTm5owgd25iSFoltlgnfR/jUoNoMpgG
qT8xWSEv/F2sMAW3kGMB9HS6hmKGG0Gxb1dN8/Kvo6H16QscDiC2HybKrdc2j2DX
irpytPgQCCsjDxe5Pl8iety0cEA3xkvgyqQKfixIV8ByCM24U4qs5jvhG9wRdqLs
89FR+ZOEI5+FkHceDiIgxtgnKC5I4uHJ7Vjk6+YZerQrvw0WXNse9onI4+kL1PNE
+RlvLVXkWAwBfWKMZMvYkhD47IvOozUXuMO2ARWOavqcYPXdw9PU+azrXqviqbgf
GRmWNLKG/I8FqRftzmF+LqzdF528T8LS5gAzR6UIoc//SCQnEDfa2eCzM+qAH+mg
sMQn1SJ/GYmFBLXHFS7Zyl6UcaGIoGz3kRRA3tLoSjpGfWqDnbl8S3aNkdZGV2UJ
p0NVWnwqYiq40OsYcaJhhGMsASDy1n9e6EFernHj0qBoZ0cW8QMYUXqQHlQXASgZ
X18/d47PjsUgmlBQg0lEYdNcFLZPvyO1sEaHCQwrsyuseReWjGDsR3Oa9+eXXMUm
krMjYZsNQ/y3uyFQDapILopq+ais1EKURrGKXQ7fYyFRHVtdsiy/Fsf6eNOn+3/u
WebMQFcnSZT6WyJweq4Qazp5BrXxmoyc5OeNTfzL81IBvz1qMxR/+4qCxDJ/PDp5
IGk/DgU+kVK8eN+QYz2LnCfvXJvb2ex3h2DgQ3pwIwBsRnApPjlymvyU/g35thON
Gsq+xUPtFWJV+7oSxCHNVcgC4QGSWd8DVkff5XDyJQTJWTOYuaZ61araZV1SSiQ5
kn49VRmmEsWxMf1SMDi3zh1CPeQwHIjJMdCe+dYtUhtgNBQT0yPpnMjIrWrVuUXH
CHl2gcPg2JawH+wetGufMzjpepeUpf3x/YIu+WiD2asyY7O+1IfmBc1ilmZgi7pH
57DPGS9dbSbm5kk/oRCXerzqdg9OYuTTD5SawhB2zhhsd6DKVYWDPJDM45O1FPAJ
gVHG3zf/31P78B99AUfDc2rwVfF5MErhkZxNX2NBfqk=
`protect END_PROTECTED
