`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5BBcvUEsw/HVwqFLCqVhb5E+ms0N+WZ3HfdZV4vyrw0+B2jpucXCfbLaoridRWDy
DrxZA8Fmsd9xEm+YaoQRmw05X4OXTnkhEJLWOo3Km5SbwW2USrGqhW+wjKmoq0FT
tYJhHSI1d91BjtEpbGHDtNHqkulp+g5sS/teZJpz+TZqvjvG1TOjKVqYGknwrZG9
UvzEXBJeM45Hf9Um/ngxKgYFQDp4a54W0kWHw6VWvjDQS9xfgDpmyY4gz/94IP3A
yGQbbb91Sd+VWX/mQwRYhRMIza923HGVcPE7qivEU/Ka16sRpZCx/iLW5/Uggpi5
9m0NED4g/O9zsHXZng55gs4KYSfwhVkVcRQ8XK3XibgyN6lbYBimGAX1sU/RUScQ
RWrd/6AKPIH2NpT94+ALRT7K7k0qZQniTwuyUTnbpdiLn75TnUQMkxV4oaxcMO54
58Am+7uVIARqJoIvk+Zubq1PZ1suQYoi6bOXHST1tMfXoGw/di/dF/a74jMQpEn6
62toFKOSc5ZGKdg/ZEN+6inKFcUrg7t3nD5r3kSYUlfW98Lf3O6r2Ymjn8wtfEPH
DU7xC28norpUICCwi748O/uCcUpJLbgMVCDMVkML3eHP2zMSGLDMLhV3DzBjNX8i
IYeGc4qLpVzmtabTuDbx/FO6KnCYLlITFXSQi41EZXTEWNnSfaPaSCqLvnJfruME
5uIsAofgdfilY/4kKClFkOvJqCEoffVngN3WBt6Jx4p0Jb20vL2U9gxH9RDxMbY+
+Uzq1CXiupry8e522pUW+q+v8lKra/6ylV0ns3wApBHSDOYm1q38+6Y93IGbL3Oq
SkoyoM23tYez/78HohYJxLyx4lQzJbaYY6ubwrRs5xBjxuZYng9mM+luhjBXrtQe
/Ca3pEa18raGiZfaqqa2Adb7uWTo0OpGfXoGy2CwYwfAwDPcmvmYq+9VfR+mRXRv
si+pTqXcPbUmEP5gHOv5dluVvdR9QrUVJUBPZtdIq1Uu7f4A+7G/K0MmQ2I2rY+9
+jGZQFVswXx71KKWjoNmwxmiMvwW2BOjb+2LYekVtSFULhe/NRCuqAWKFzRAn6/U
ppBxBfXzDmLwKFGuhlbC/nDxA/m0m/ku7XjgIYc+nnQGX3I04GBsHJuXOYk1haUP
u4lzrKoXDUiVfzPOKpOGcPeZl+bFlYaoevvsVawrJ14=
`protect END_PROTECTED
