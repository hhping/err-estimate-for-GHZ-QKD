`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTq/2KoUpTmaXVv1UjM8e9unZxer/9ePD10U4DVMdFmqgEeHk9FjYx2pZ09a9krg
yz+MYlxS3T6iGwlibaOJZy2664+p5S0IOY2pNphW5VYbcyS1s9Y1o0BAz581OrJw
5jNx1Gu/HUjQHDHxUcqLSkaJThm9oholZ7WQaBo+HDVhYoUoaV16RE4sgd1x92T2
5qfJsP3VJMBxzYXzTF3AfJ1hk0nkvHsTFmoZ+Yd0oM9gPTKrTjyUV4KRyPIKXyCR
58cg3qhEyRE/78ebZgEYh7WykMbIyRSiTLXbj966AkX1xr5HlOOWbLGHuXqDctcm
oclsxJ0iJaImSsQUGxck4WsNOcEvWZAWcW5qqkiMtWccHN71N8lsOOugEKpJ89O/
385WuJkDAfKUq215Wyf2ZOT95zvD1GlDdJ/fRgSv9jceUAkUhTGnFqM9CBZRc/dF
PuU8mVTPd6RrMaouqSbCPt2Crq90dP46Jzx510eODpvfgpCh2+OOEvDu4Jkus1ZO
uJJIYD/+Hp1v1VEILgo1sCKqKHaOVWyZsNeOxdE4HYpDrkSUQmrX11y2uhaCxM+T
1sjXZIqLMB/PewKNswJunxAiKTRhro4YgOJ3b0kRi51DCma5RCsHgzSfIz4xTwBR
dV0fRuXox6DV7uQXdOV6PU97Rz/xwVdOTAj/m2uNQT6PmNV34VmxXRR6AEReOkKF
/1v3k+nR6ZXuFHTDnnun0QEe4sLAeOVmgn/PLeJsi5Cx2dBr6qIKrOKP1Xbah/r8
P3+rXEqw3BpPk7u1l3k88XQrWE1cD98DCbqvqayFzLWb+1tnMifQsjmqRaAjSREw
IabF7sRB8q1YTTwSvEjB+7bDxlUXaWZi9cY+Lykh0re9L5J9/IN4hxaGqU7Icw8g
MVEVW9FbinVqgkBfH8QdXjHL1Fp8s6AGKaeUNNAik3wLfjv9minq4l/bbJjadUpm
ucE+khCzuDnIpkDK018ISrWu+hmzVrBAQun/f4bG3Mdkzy2/llYad/jZqoUFswfm
MSBPM/BVV2xkwY8P+6efU6CVtw4196czZMXC0T4rDvE=
`protect END_PROTECTED
