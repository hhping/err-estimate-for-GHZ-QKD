`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmMo7UjvNuCVcawpcqVNwBp3gFD2G/R+/yY08w0YNUqYbgWRUHuzNLb36Ykegc8+
GPiIEI4NUsgx1uTCpmx0xM9iluX3AYF23thw/wfVZVhlesexGfsOxiX6kTVJnBJg
/DPP1mJd/s0/tNTK9ldbwQpGyzLYpiCk8vyr742vELvBeORB7Qa4WQsT0x8uR+UG
i93e96XYyQ8XmehlJfvPfo+pNfrjBVDuOln/o+6ve3ErPE16wMryvFgzwi04zW3p
cd06bWI/V5WufQc5+nx9RGpkWZhjaqDoatQjLo4vsmRj4JkTETp+fzXtzs9sPOg/
p7m4b/gdgN3E2PUA2GKWTuAIK1Cr1iqJL+msfCGSLjxFWoz7xFGMK8OgTUmkcT/N
1oJKUsP0hhDzYq503MLmLJDGqZq8zyMArGz8mYtyKtULius436Yo2OXkJ2GTMVeo
cDnyC7oScd1N6yTqrIoQ0MlhSdC6S0WwYWnHxGtHBNMcXw7KFGRl3wJwc/Hb6ITJ
4Dq4Xh2QW5c7tkMoMMEkmYM7NCZWggMgnNqkOI5Tqlw=
`protect END_PROTECTED
