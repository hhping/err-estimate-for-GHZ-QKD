`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0w2igpk3Y6yvbr2SNMKWfY0m7nnADYXR1V1Ms4/Il07vQYjbkiZ4PqPVNZJvLje
dkSgyAB3AsihX2bJ0yZ3lMTD9ZAa3r+HFW93PGaFscQ0qqKHqCG1o4uMg9jFrvAH
ErHHXgwMw3+5IWQp2IQpcCPi7/nEvjppW96zeRq8OAof/mQV3y1GyVYAjeBrLwIk
OyafvlOsXhefAlvm9qgo3a8UZolOe85Q1xqWNJWHfdLZydp1Tc3WWRiIboNLvFqb
9Tv+GDKKrGy368ypa7cJb5Nhf2HpNPxt8K0KEialmxfv7+edW14P0J1cTGIf5t/o
XEw01Civ2S/l1jZ2uZoGjNMPOpPy7LDH9eST4rL40TJSEe7p6BZBbpSPvV60/HzI
Xh1INrD/UDIe4VcaRq9z30wV9xoPDBiyM9yFF+GrgmbOoXIxIyXaoPP1UxyMBohL
nhJZ9WpYERBTHDTfAcmgoC1joyI0ju9MZ+cjYmtmjaZH+LIzIuIemeM34YTczZIy
nBrXbMS/ZvLD1sKcRPujaIVGTQNd45Vr9BHDSHYou7G+a2KqDh6yyj7GOO1eC3/h
hnRyVLaHmB8pyrX92i3q1/tOgBeXYrhOZgzjr1bJyofl/TWjn1Ux2O+Vm+dmpNW8
1xlq6uy45DVRBSaL7iXRgQwD5gVQeRfY3NhHvi3v2nDXKgEmSv4l0aAaYzmhDHkY
0pcN9K5bI71QTM/WMWsqARsvw6DHbZoQibRhpO/+7yO0XAD3Vbj/sfefwJFIFqTE
UnjTIRII46Diw9DHsF9ORSH+tdNvBnekfp3QxvaRB5LSCotKOAHCQyC1MuCdm7cg
wTtAR0eFAU/3D/q8eSXtDHSe+aYEadqsMSJXldOl5S75w6XU/zh30rWH/ivKOo9C
n+iIDwtGgznu2oPZdDTGjplfDZOCsPqla8je96xo6L7VrMfpdZ3vu/gzdbO1wNcd
jjeC7Vp06kTwgriruCHFWLoXSq8Us1nye9SPrA3LUhSMXG7slYsRiMXWw8Cz1Fgj
DFReYN40MGeSqwKg4fRYROIbKSOkf2Vmf3FPBY2uGJlmgsHL3/LX8ueRUsPW8Emu
fLZRygv3iwSV9rCnqF1WH8sov2gmSs6PX0tvB27R4bjdWPHH3wLtda0AXTu/aAm1
HYUFtc9IaGs449SGIvAPScr3MdlgPnzwgHtb4PhY0sFxvX+wyknJsOcOhSiDfhRR
Oe9l6bOJLx+4ylGedCqOwj89oJbzv/1+LpHIDECZeEE3gSLJTmurdfoGkQEWWPZm
nGXrLt9n8NNDQd7JVkSopCFT0dWae6Ny5b7/oHF+j8Sew3FERIEYc+T3KfzzcqTV
mKFbw1m4nrTuKKIf4BxzPWlLaYHGLLvzxa72iCc8PoHkAym7hBxwOfyol+FZBKeJ
RvprMFNSG1WzxTY4hdGE960ysgJRBbK8JFug1pwLz9n6inyPbPn4diofuc7WnyE5
LJ68LuUTklee1Qqc1sspdw==
`protect END_PROTECTED
