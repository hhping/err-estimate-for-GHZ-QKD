`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsJs+QbrSAg2JVeqIdJIeJI80vVPFKbyurwTTnm3+7DZYQv8vri42yws7gFmzxOa
1Xr4YibYahlscARINuikzrY/kgJEFNnyuLn9GU093MByMsSx0v4LN9aM/vqpklNL
h38t+1j0OkiFaBQVBWl69aWE8tx3fuTk9vMN1qpqE/LEx00AxyJgy7aZAB8yp9eQ
iD4VDkpZ3BgHQh5fVUcfl6tMfnPKmKbhi7DkeQDOf59XNuujbs/P1liQPQrehHLy
+awxXPmIgRaT2g/Yf4H5u/E/0pixKxNLPJ6P00j8V+VOlq9z1ZnnzAI9I5+BdzgI
lA6JTYPJjL4+Nq5CH+fQrxmK+rObjnEfwvrXnnMaidpz1zcXPvOirK92ct3Ksj4V
zJUdAOBWr/0hK21bOOBKc1TdF/NOkK0gjEUBvX4X8Qh3molvuGJzO9LYMQymd2OB
8461at7CGP0/7h9PZ7kh/kDBr9I7dUGwg8RXGE25IDO8ZYBtI/fNkNHwBcrPlBX9
Fg7dsGYfMcHAoh1wwbP2dqlOcwbLiSSLINKsdZgn3opCc54dAP+NB6GsMA95wE7f
qqkRlIIk3XsAHx90PYXJf9lbgLY5mT5+fQyeqyUP92fh5cNi6C0jsFCjU9eLYKWm
IYv21cS/aj0Rw8A9XIh1BNURwg5oMsmEbvs9jP+G1uKH3i223KTyxO8wbUNqLQyt
hpX5AWZOiQgF97isCrTMN0NuiLM8jglOV4d5HSOg9y5af6/i7DtJk9UCvDq3ERFA
zYq6b4idZDs7Qn1xKPMCqnupJ0/uiip1LeW1+kGyEUcj9VvD+8S5X6XFAx9Svgsx
86+EPVT6ithcXq08dTCdvKyQ1uMtU97JWYCOHAUqkys12Burbq4jifRxAy/8j1Qr
yR+eSnWBtLr92vrlaypwVOR0Lw/mFgvwcMABjCpDxcFDFFJT6/gMHIOa7ibGLpwa
eV4oI5Ey4xEPNaIUWKXnCmz1PkYcS7SZDZYZ238+2X8zD5xYHGvsGUjpIE2jyuVv
Z9dXte0zCqPVaGC5if6Ub7aZbjFUyosZl8ddRtz36F9Yct/tfA4LgOrn59L3T+sH
J5AcmGthZZxXm5cj/ui/T3L9Gkm2WfCVmaJCgwB2aWIKFiZHf3Zb88lBOYKyhLNl
ats+lssllm78tqhA66W8lSjlXk3sA7l0XsFB3xbN3dfkemgjAlhllaWWxQarHEjX
aJzKRGw/NI5LLQhpUB9VZqGNIrtqqAoDAR9Qxcc5UWeFoobb0wBjlzhNohGleZQo
6cAL25VmapHpVRfYDjQVCukG3RggYdeoYnLuNAQhW8Nr64YMCO+313ZF5kfdwXXK
sbEscIPBArotEtSSDSaeH2GedPBAHgWpTVwxwb+xGmbPtbQgOy295eZBzb7GJWiZ
Hy1mUg5zspNvv0bleC7If3LeltXxNTDfJJoy6xMPSveOmcgqrOJoGC+pkmqPXKJZ
Vr+VfLs765McHh+ODEy+uvpr5A+Oi6pPb1ueVtveMRcyoM5Gj22+ZQTiaxTQ6u09
TkiqekTivum27s9ZJIr1PyavndamQWCc2L+16Nly1b3FKgBlhI4ENgxbA/+vvfD9
oW3vX/RVTehS1+6PyF/vpkxpqP8qnUEMdyaaFmQdTTrD+i7G1McLDnvTxIBzA/ti
KYfzuWXvV0pNysQTcD8rhrCzP9QNUjIUo20y39n+zqvj9OkLN40/yFVgTUrWdvln
1qv3HMAbQNXTcE6ONZBuODqOWmxASBNQiKi0jIyFyrSpyCob81pmrhAZpU1RcOZQ
VkgFyQo0CgiSBXMFvSC7+Fd0zXxUR0smKwfn+7koEALl/UIysWLUfZIUzOfS9nox
mzsf0N0PGXJrKi3OO6LXl5DvoqTRr7TWlOvWnsj+BEk3G2AGZwQPXI992ZHLH3gK
hxlzwXQiHw4NAbg90i2jxMealCm0wS+1lu1yGQiUvLE0h0xza3OLGXgMEW+/Alff
gngb2sgCcqWnmv4Np6YqmhzNAdvZxf350+UnI7haUOt6HpVeYK5i/4SliNJWQRvt
MpOBu8WeN9UYv3ytpHNAcjXoYt4VbwzRTM+CLkhPYqMb0rTF7BK+G2qvCR1WDA4U
lSkw8fgUNG6h3Bo/++y8PFtl+WNbIpJ2zmobnW+Vt9Nt5x+3VY2JLHYGSkxtonCw
LqaK/L9YfUlN5ZYJbCFQCL+Jm/67gV3IL/DMjzhiOt0e9YjEddeC+9CEXe22BhNN
DO2Fmnf7DTv+VwhF2Fj/8nHRwdz5oXMoUe3xYYWXnG3gHDrQ7gxLjgPPc2heYBtZ
krvfQqV7ycnI+YsgmzASDDeHILHN1KGrDgOgUS+7m6/sEOAyVux38KTSeEQF2ym8
Yz98qhr0O1B7gmL2PEAJ4y3UwvNG96bJLvejyBCWiQtXJ1L5uHe9uDW1BYXEoK1O
fnN55V1nwOpHRZ0p5l7zHfPL4L6XFJ7bmeXWpiBka1JZAG740hedHgXdyM3iPp1p
p+J6SojfDOOOPBp4bryO8lcSgGCd1jISOH93VpAehKRCepzRlz2QvOojCnEPQntB
KKcPJUgI6tAWBVi/B/PwMnLMQp80KmsWRhcGSK5xF1haRNQRqmwvHxUttBIqCgAv
VUWE3obSGJn1v9A9CP11MUmqc8EPk/QctWnJ55RZk6nIoZrKNdt6gyRnxZj2rbmX
oJHNUa4ykqe6rez8eYzd3tCBI8uxqbEqqNqOT9Ui+SvRndJiKV29bqYualhm7+g9
Ah/Pl9MISLYNiWBx5M9JgJls0blmVfry3aNuArn/UY4dg0wY6RwP+kk0E+ioT028
7VU7tRF3oYCWTlMYqFx9cIfJVubKbaDmpQsIhN44ggWksaRBh5yZ9Gxl2T0rkQyA
s9BEil0iSmHJArBFLNvfPpYBSxKhiQG5GMTeZJl8RzX/1sgJGHnG3NyefVCNTdDn
kjee+kqHdLQDbyNnfmLdfkQORAR8SPYfaxT/Q6VYjq4dnGYATcaFJO1qF3RTkqt6
0VMhdbNNjQYA3bKuLgccAU4sZG7eh05hLRrTS7+uSZpg5T2+8hKRKQFvLQ+Zl5w8
IPECLIit6rrAARTJBTYK4rnCGs+J24lm7fWfBS2hM/n7PWNZiV17T66V4v7Mtxxg
stYsnZEdFcGMbXPO15nWKsR1K5mDnm8LHdCt0EFmMa3w1xXwVIg3ace+pD4PC54p
kkI6HpG0lVLBa7G0Fr2g/Ntcxxl7mpCijxC1dGymxiTRe+sXq5St0FRBm3jNdCsO
Rp7k7DVGCFU+GAE5rAGN3Ceyqv9a0R2msIky0tPlT8J5vUisnjXuu8xWjLTPp9Ct
e3FxDEp6yENXORa0e8ei5O9pKPTDb+I+TaqI4IGhaGHoSDp/VjiglvqdNVkXXx8y
AJurGsCCedk/7QPs9AGAzFS1QH63MWAthiGUweTVAPrPHnUMq+T6AW5Zzx68d63q
wNDJ+4p8Ay6unN3TYujw+N18sMOW04JKzVhLgwl2z+XrAPyt7EuzUUcftnv+CCW8
KbW1mDv4Fr0neJ5sCALI4VC8XifHIdsQptpfvs1f9jV9i06Kt4LHhAkdPBI7g9H3
Xpv6z5dW1sj5Owo5DtxEjhKtGVUX0QDJlO/2x8fdWx3Y9qNT0T/oH/jkf0i2OL08
acEgxt6scew1ifGc9yTS/cJkhOnHQ2x4/M5LSqjGRh3OY17xDU8OwlaQaFVEQ+Xb
tfB9aeDBoIwLIY2ST4ZYG+mYcY6N3hqUUxWCNePWogEVuWM4nx0zXPNC425J3Sfo
f+D33z98RRsoNbzZAofOPB+Ua2AmdWkHHZqKT5mB2NqsPJBufkiDtiJP6eUG6LLr
MKaXLl6+1A1wRtx+sUyKLYi+SyyeOTRH0h9mejWJt+atqTeeEDShFp9bqEo6oMF1
15wxKDIye2Ni6oQfUjTCsAkBdUDs+7S9cAbTRq7E7WpzD5TZC08V1RCfOXjPSxnx
kCcsJxrSnyQ9AhjILgScHbjBPGomLH7Nu1zEiRoV+NXDVbnmh9nZvb6+CUs3BXZo
uLfIXdZI9cfPjNOp+ub3iYkZCUPW5iwwVM2gelZygysohuZwSC7R7bWMSQ/poDwl
uE4gtZ4MQKw9RHTBzlxM2EeYQm+/lMO76hEJUDqtq35G/yP1iydt8It/KKOCTGIf
F76ylkcL0noPjKNpCjZFbP4pP0pjvxwwXjmvvRPT7U4slkLwoy001n/7lw4bNJVk
m96FMsHvvQ+GRfVMNZcoKNNX0oxcrkHlTxx6l7RYg5uXoHBQFAkkot4F911ytlkw
LU5OtCoqKdk4317W3WNz3MJb35NFdXAZe2ulNrcwfUGISLgXaQyJX57KlqKahkqG
fN4Any4C6aHab8kXqAGbnMYm0hyARt2kXi30LKKs+IzPGEfP7fVQdRSrChqF2+x7
yK8rqMgckls7wxLdmLZ12+uuqabp4noba90TK6L6GuevaFHmmf79N+27mLfx6cKQ
EJo2HY2deuOPJbJgB5hZbbq8DXq134Q29ybRCZibXEKS0Utl7ihPCocKAG+ZvVno
0eD/ulZFzBnsU57ux80wDn7b9T0tEtzpxxnzHUyqaryGt+CAP6CLaFJyoJ4FUGix
v+LP8395CRHJ1AMdBHAOsPYIR0xpiNiXPAUMd/uxnjNfnNxvxK86/C4FbptRNkab
TQE/MCpvIDjvEWHLEMhX1JN1s2GopcKwpJtsRrlyjGWm3s5xXif7LdvyQb+AOyZX
W4N36fhW5B5RW9bFKH1VqhxFnJTKdeb+udr/NaC8kHretUKctNHbCosF/TF0TbhH
4nmrCpZ/aEfzwhXM1Ln2Ugwt+B+i3hG9tiNEjMkgcjW7A3fYe6GwYBtTCywedIjn
Ha3Ir4MnDaq6pBg9cmAPgUKhuqCDKyk/iH++UVJIxuSqujW+XlG9NlukNDBLHTrZ
q0mqOmJFTegfBxN4nz3jdAoxvfsyeqyLlkyhEmnmKoqri3hVYZZT1ixDMYEWhwKm
Qhjg1tfuK/OsMoogr0vce/cisoa7nXhlkdHRfnw07EasAezS76Au88LYBWSaptHd
mi86haSiNYJpM+gkHZijdxbCBcv/OAaIygCB7imKfNeixTIRVR3+1JHiZ18fv42Y
50CxawQEgrCFNDORO4Qyi9VHYMCV3Dzq1YQORPLVs+vwmWNwc9xEH0H1g0jP+vQM
BRKmZZrM+J4rfvKm6ep3TmqRZFkfH+Oi0jMA0pc+0F6yr8f/IZOAILFXkEUo+WuS
GsJ10fobMOQ2NCq8UHR9hA/T6ZE8c0e2Gh1DKt5GedalX6ICJ7lv4qYcuXrZZCCI
m98uNPEKibn1Mw8reDry0yK39TV4HhsgyHYhfm6S98zYo4FnpsOmIAVl1B1mxn5L
I3xMAZAR9Ei1UUnDUomQmXjZotbwJJTUvHp7MPtS22vr9sjRT7td5+sS+79Anpow
aAVad/MFta9UsWYIlO9DeJU1JnuCBsB9CLvI02DqJXnfU/l39hRZwrOftRBb+FX2
gd6ocnujdnReq4rlUrPIBei4QNFn70MSJeOIlW1M3GA4vkqHDrUaTSazdP/qbIz9
lvqL+csTJ/cXQSo0XqVTpiIS8+4mzaaWLtrBNc14lWZAv+iBb4BMeCV/xrIKnzEq
36WaS3DhUGHAKqccGJPR5sSSFeF6Gj8XXYctst74Gdc8AixUSvrq/In7UhSQGJ5x
G6fmG99emr3BQ0jXtpQJtUl6AEqn3NCmiDI2/AeeSLd9lY3xGj6lJI3r4uw+RLSS
9vTC5KQ5KjmvhxR/TyixOesvehT+tGbwYoi1FJZBjBdXYfSWbpY2NfXizNcNOuPP
lZK9KBfpK52AdVWdpncXEjIBoyM55O38GnKSQ/cD8Cd+Y1LseDOpMeCdaIfGpi+4
4Jnw0ZsnUwWbcBNJRdX1Nu95LVloTC0Ri9qfjW4562eDQT73CVQPPMdJzGpA2RUb
+EelSdft0IVFYaREABjVHDbv29t7ZoTWhISknq3oDNqnmf8JvkvJWkUeZ4Jl23ez
cRNRMrtMUnAY0W1jOb1ep2zgKQd4cRtozDqIALcWQCoNWsDW7ftOkgdgXeQeoBGT
KHNXuxBsBI2n+RicUz8gtfz9I3Nsr0AmtPLA9SoJ+cVCpqDib3ud//LuBwtGrw88
GzKVe7+Z2bytJKWdd51u+4Jdn2zbxBSAhEeS52qlbKy4SWClYsQulYy/ZxHDcFOv
6+s2YONKDwFGvqlou+q6lp7eN7n4qf58iD+cslde0ehVS+eaKa0eXGgGpOVhYAQt
2GUKyjIcMQK9O7M5AjuFF2NCMUhSwqmyfGxI0WJPvhq2VpDUpo9+YTq3/ug7WAAn
xoQHMokC3uiSNZIxmhCq7AwZhj1i3q6PmMMoAcMdcDBRTr5+t5nTLeiIUv5Q7F7n
J9cMfu+2ZUpz+g0RZaiDt1Oyy0s7S9kZ5noUtCwlfajbJlkse1J+w0JJqYos2N3h
3deQUBzvwpqoO024tgfoyJwNgk4QCm7vhgeBWMvQQMV0EDu2MPJ65Njgcc/a4gSq
3Krr1LntVafMRcJA1dAUKNkDhsw+0Ne41YSy3R/Gn+/F2zZy/6/00nM9x2p8sHag
AF7ra4uTMOKa/Ere4aQdVuVGSjoQfKQHDo8bgRRnNY7M5qDh/MP3MIRZ0Oi4NuYE
AjQwdZLf1/RPemcuKg9OkhWsKkHtsuQY+5lE0MfsIdResoc4BlRu0Irr/0b6CYlV
PYJQ+9souFYkOkFiFunOHVN5YabPqHSP0Pg7rV4UxOGKEJRQ9NumKDIJVx5ZDEGJ
+u6GWDhK4j2gmfVQBHNIvHc5fmoeTtIyPkZ3oNbaRPfO3mOTVzaV7Q+f72QYBr09
7E4Moqtye4lbS/H54DvMK2zMTWtdEnGB7y5X+mMSzstyiFn1TVQcAt6HiPkptf8Q
WmCwdWnN30DP21FWCuInCn35rfCV7zCv1y3PxifbeIlY0ANUP1WuETQrI1gBYnNy
J5V0DiFWAIssdywhRTnYfLOEEQDJpJTA0ovhXOnQbUgU2kdCUP4QUrqFRn/gRpdy
XeSzcGqjbemP2tvns8CoqPrTBTr4g6pocakuV+6Q0HIaCN6fKuzSQgdiXw1Z8+8J
m8sBxx+0Z5NBicKxszdV1jWB2UcfTmOFfm4g5Xi6ufwd9HvcH7zGjGc1cr4186KT
dwKunizIu13PtgD6XO1mfx8Tnf0aMdTyJBfvJTFrtLcywF9fMTdCqTYeztV0Zlkj
NZPaGDRztcj/q9hbdtuHe68/aqFWW4Zbib87V26LLFeSRmHB9Vt/GkBX3K1Zd3rN
Q7W2r4koz9cHu2AA2lHBpquqU2aO7p6xl3WYarG6xuLxi/lTcN+w4uUBJ4hAB+rG
O9Ngetj0t/koTExTc/UCNz1uwEJptjlLsYoUYOVxNYKJMX2+5oj7OqaGdbAnygzR
YY6aZTtMd22ZuLoXWlHYvdAaqThp2XoF6r3Wyo44wYJiGPlrm55o0E+TkUNYIN/e
eoKNH6ZI+a/pZsCwD/UQYMZeJW7iWZB8Gg+pSEwHS+kMhKG/AjFkx6/j+K6WVfK5
T6cbO3T3U+MUEz8XKmL8GM73g0RuvF3K2hXoLGwiGD8qzm0DWiUoiT9zhY4sbOVE
K3gwjbiBcwROVPAMllcPcB8Z1+kdI37TfXYyhApJYykT5SuUQ9N8JV8vaLYyOmyJ
L47bIX2FHb4FTE6blfAxN23yDo3Bec2tau2wqiH+6BnAQAUy+q/s5TNUExtCK0y6
J+g4Gt3no9PSStEc+zrkSDh65olcMgLlaDQn8kFtQnqfodXqQXNDXMDflNQz6ymC
w40oAknagX5k/F0YBYUU4L2aee/4rbrmFOtWjBcBBUxA4J4ai3M3+6UBhws/haDZ
ixboI7En0pqjywFx6Lqj1Bo/eV5vfmYXkpw3tok2e6rhB1qmtT+Id1unetO0XeEV
Yg1H415Vm9k2V6fJ9Mv5/xOozUBnqv0bq4/OPLZZTj3nXyQ97NJNmVL1DZN0uoXB
8JSGRWkuP4QC1pAzPrHmylZnQ4O2ONm4Oxx3EL/j46XA4hua9wvd4iqICW7K6tlg
LH0XXrw0uz/rCOCxmvdtP5c/0HYaCPoL8uMrUSdOoFYAHVvQWJyD++2RzAUMPn40
DxcMrFJruoMXgUt1jX2d94Xo/j6KM6CQcj3vWaDAHhoI6ZrGPJOLBfDRJhvDH5x/
OGW/4UnbAzQsNjDznXXpllnADXdgSCJui6kfV6g9M70J3aZc6I5woNOJvNDMAPos
Flhy8mdwfTdGN7V8eBRDRDeT/jPtNMU0TWBUSpgiY9xoFBqwL4JrwncQjtRkYjcg
/JmUu60quxUyR8AXfKnILaoWUmKr1OxpNspt5OThlss8Lq1vDl1/neSwhbhZ6JNv
yWUTk4avI+Ps8nmpjHb/hq6rTfgxgBEd/MO3OIKyjIPFfORbKGGoH7vkzClAwxFp
T0lfj5f53o9tEbgfIc5OY8RdvRmvY1s65hyiPipHYuzSk63H3ZruDVmp7/LSsnvT
+4j5+eZ1gGDv0763FOFS6gZPI1W3ws23zwMIiaZTRNiIGoOPaULcdun1Qxf4up9S
LShcPDOXfwX7KR/yeS4wftGVQi4ftBxEJTWsIqycxUutwIuEkKKWiA4CY0iYWaNw
pIaphxfZgjYe+3Av97i3YaHgDZRz0y7Y0AYUK9DYnKI1PdYp1Gu4ytAUjozrCx6J
gV2mPJW8I3LOkztUd1QRoTVl9zPpcYQbprW5ArXs0IK/QHYmEBWjRsZVOjbAz446
bmUZFkIV9hWqrKFpDuiJAIPosVbYckixAxt98b696Q85Xf9MCC/HedjgsDbgNtC6
Z2s0coZnsNgONaBoJlK9Laq1Mvs0Y1jSfyl0gKZBrjvh65jDB47s6nXg+8+IVqiB
YxCpPLyUrJIzCimhxGHpQGd7EYq03EkjLpPcOx4McKayoEqwvbYx22Saf5F4fvCh
8P1uwkit8hhViMWtGQXAB8wrXFyN7iDFSlKnL1ONrdWdzJyw7Rz0/Dywcsp9fwtk
fPy4eAY3N/1MGw41VS/jfBMeGNZenIqMuW35ltOkqldljb2fkfYb6/aY96OvtAFr
I8kQoRkvRGSlMxZ0ayucszaNy0BHRuyFIQWTTY/4iSohh+j7DLSpY3zNaQ5s0Cma
u4WXu4XSKwzKmT0R6Ls6fBF3vc6Gahhi3bmG93CdxpZr5MuaCwrXjNLxBqP4zcb5
R5n9HFe99yHQjzwwufiRAEN27FZIdj6zSLxgSThZ0tjwnZdPDSZQt/j+x8Q3tORw
zcyj5G0r+du92ZGkGHJKCxzSusm0LcOLKASg3xgCBFJAk6mGEYEuo+bJKt2iN+YW
Kuf/+N4Hdm7wgcSffxN8dlTPYfuFrf7iQabS2VybwOWqF1RBZQsLjx/fZZIsd0CP
E0bJywVPgPdCe6vcqchjKRix0mDHICHsUSut8cBYSk8EVCEakaBGUa4RQMJm9EX6
OYTaPgwDhd2GBdEN4VGOTijvXEZsWNWICcAtuvUNWuwcr1CehtNcmB+PpA3lqten
RlL4z10xM3IvCa9fnLz2Pn9ov35kvKdU64VYe7L7Zea0l2ENgegYzAC1Gb/5BAVN
OcG7ZfC+zt0YTKh8yoVFH7YnstOyEYyejqnhC0EO2Bpm1iC8dEkRj+ngeWkhOwQl
vhFJneQNG+UtVPGm0BPzQGdBJtd6LR4P54mBUn5dUhX0ZEyEon1QgubVVItMRUWJ
EDwb+XgUuIbZCLihybDVApz0j9nsVG69ogmDT663rALnIvpbQnhtDOa86i+XJGEh
Cg2RYsSgqyfQIyqOV9K11ltydpv3hmutidDUwmpdwngU600r+UGuTGLfUbuo4J0A
bV+AQiwwCxY4vO9gub8fVSszFomlHrnyl3H7U7IocIxEOv/zW3Dw4JavlvE0U0/b
/0tbP8M2sLaaMi3ZAqvh/X+TRl6EcV++GWsyPamv+L0EslJqmqhkBGeqxmsSLPLi
oMwL8hjmIq9CPWvxuQIYWLCNpfUPWhrhxi7V03WqtPFRk+3y8Ixa+6wt7R9+J+wL
+yezCASqcn/0VBWRFho/XoC4JDjrFKnvzrxw16uSLTTnnmfMXmF4axcszwKI4O0S
2KdhQgGbUVxrLWzR+Grvi9Ph2Wzk9iZMtQrhV0Hrlw9tXeKi5mPULS8uXpezK6nT
pyGg1jrbOetdvgHRllLu2ohqG4Ojs5M1PygzpYv8eeYGIvfbUhJLKAIEY9ArEx0S
A1bnK7GOCSzy7hfaICejHEaDOUUCCSrJo5HNvAhLiE4DF6xpgbi+LJFl4XIm00ma
z/NMWcP1wzVkSzTjEsUybp5qmREB2Lla9zgc23J6NuMWUdOixiksO5zFTDSzvfOk
qlg9uGikGaOUCq836i3u8Busb/7OE35bIChs5ZmVY7S/RvWklcxIM8sgmGk/RxlI
7Z92RTzosIxn3RcrgQU2AMkcuGFVnwNeoAAZMYv4c35bjkEeD460qb3ORC9hQgJ9
GJKbSLvHD49iisfqLiywx44NyrKy1CNZUF6YysuA64HYwS3MmehypcM3v2M6EnPU
p+AB9qLrZuEut9hxPF/4/3EfO+o4l4964echgB2X/ishSBedkuRPjW6HKog7ikek
SQA+N1Ur5uehTbORctlk+NTkoJ7oiK3zvif9JQjgORq1x9WaU/EEPtxnUzV4+nsb
22+2tHeJHzG87MOJlf3A5SrsyIhhqbnfyh0iLk6gpoN9cP6Ix3OPwUi5hd05G3Od
tiLOYP7Oep1i2kUkJ572AsS4I1eby9oMCjXP7DyWh6mDee92UApEDTLMHImkRdXf
wn0Ub8CT25q4JL/6GMugT0Lk6LL7ZO6/86Zp0W7X2xEZjqhIV8b3y5eXZwMu6q1Y
niKMHlHGw0xvlnyWFFpzW+4eKpIYZrqkKWrkHDTnTczV9J6eu+U8CTY7xOJ9qbYX
TVO5gviUaEsiwnwq5xIJOmlLnZWddnteZtzWAAOXJWWaqcNl87PPU2T6uXMa8amX
xXN8isyHmJ9i/0gVA3qWX8u3gJ/9+utDr1ZpUrp2ZM1zM5KOXVL65frjOaP+S8uJ
ciQVzZ1MnYxfKcho4pCDtUMGM4S2l5CrNDcwpHHU9T+zQ7akPH+id5X0/1jO0J7Y
X35wj5iLFh3JRJqLCPVZPokC7U2gXa2tWGaOGErEeeoieh0VmO6VsC8JYp3JIFCo
/IqryeSgGDIgcSRUIK+Fyku5RhkS9LiP1d2S9NxVDjNVlcosur/qHzZuJYIiNLVq
IyFB/uyk4y4M0QFa9NgUXB0QHT2W8ZAvSs/EpNeAuplfwEEfy2lT6G9Umcscp4KF
zaiLQrPaZccuAlQy0koGbI8NzYdkv6kl7mqqDTo0AzwGTuxjjzzqInHNUpQ6FW/D
C4ofUijwHLPj4hzRQR3RpmOGbblnhIEe9on9Psq3irWIWp87X47dTCF3wWHK/1i4
oNMEFt5wXGJxPtjVFcEBARTR9irPKgPHhoixJFtChNfvotzyaby3S+FkcmkCTR9n
jI5mVdE8Cpftqi7JvW1HQEDhO7A1zB9mB4zPyt5ruRZ5gF0nF8yMpDsWD0hr4l3H
oOffk4Lktm1wVkCUkSaaDDdQWe6dkOxY3KtlPgzJrCVNlNaf/YicXWjFXet8d1e1
EapF9g6JN1pcCLMkvdCcy0GFezIME1XBcWvL38ogBp7xO6bOa29Zb5UL6IQX4Ii5
B6T0iM/T3JVwt22yWZKGH3Du9RDbe2ofxe1lBtRPuLaiHroW6NXoOIVDcN+A2LJD
PRV+AeAV2K37mhfkOKm88FPe3/XMN4sVPzO7l09KOP0qe84KJDarZ0+4qah5cfUE
FioNJWEgp7gnFdYU4qtemg4lPSIlJw4GXArB1AY7adQGu19KdEaPCLxevUBxeviA
XkzAVVtbp7gpjfZAKA/JIqtdVV2pHs6ArFG1dSIocC59EijADPauuxg9QG1CkEUx
M984Rv0L8z/UlGXbP5nAPEd3yZf/0kk1Z4tPT4LGQnOxdqXqtoIlascjMuiG5rfC
qaCHsAquCNo8/UoMjGPh4aacX5tZBgBQWnumls9JVUene0/W1zSh+TCycLvWhPDV
WdImbprMdUyUqnfF9NS2rTIqUaAqZM2IiTFyJ1z0DTt3O0ag1AT1QFLdculXmVR1
QOpn4Q7gT1Kcsr491KuNOOM3UnsDFlsmv+6GFrCnSRayQRos3NqZm9lcWpeuuuSm
i8Rs03wKrLmddxL3Obpo85JTn4yg0DBk4KlUDqHqws2xoYqqp7cFccXyv38JLRta
IVUamHnhDG2OQyuKudjbGbY9Ii1mVD/2yO34eJ/yl7O+3jK8bUC33UEUMH4nDUWq
CVxpN2lHBTwoomnRI0/ATpnOC4WETVb3Uj8nggJcgm5HQVGvX3BnQgQv1bUrL9aX
daYVzXw45abIHrYeDTOOvQGL62QCaFyaLDd20lqKgh2AGypOXwCr/37xcRg9uRpg
TraumDt8v+2QNL3uSlPTAG5EztGmEhYytWzOzV5GPjDDa9goIt9ZLZT5aDuOmA6L
014edWpcqD2o4E5Rv4Q33w71Ygy/14TmBy2DIXyVg3ElRaPk+f0I0eOcrMhsReME
H1iDL8J4nxAIufDIwdiHQJP3upkK73gW0k9qwpMqMArgG5FhwSwryANg+za53Okl
4jM+ou1x1fOtZR1bd82LPqY6Npkm0VSuUvh6L6UrixUYDfi1l/XAPVg/lVMFEHLD
FfrXwQGzMhlLmWQdapF3BNJ1bUdHnqDRcBG2QxoTWCaOmWTJsVHnEgD+nLamzWjJ
QoqtGz6UJyKzsh/Lj6n0ccFf8LFM4+verc8FYgyF+2j46FkSDc6NwLifK4/IeDsV
c6IcYa50RFr2O98EYgx87PVeKpDBqlNjN+5Ae7nKAcaBGT947FI7qMN8NZkvBgxq
iSr/xSz4yGPh95DZDclFytynChkwhnfebvCo5Jph27by6GexYEWOJyDoseniB2oz
zzqgmMXQGh4GIFqVi6ikXHIxagm4zQ8/Q3+PCgQoyq+LAHu0L8QHcsaQgd1hSfHK
EFE5LQvczYTfE7ToRr2oAmCMYomhrK57gXM8T81ocaXMaOgdvHTX8UrtcSxVB96o
7rhOIQsTL16TtwlPHEV28n7l0Syfn2gRe/WNKgEKTmLwVmgC80JTKiqxcg1UlCns
h7x+DX6fzJbSQoHfUKoEAP+XBCM5GJ1mlXMcy8+rrYmHUDG5VxFioHmOJbEPT/b0
l0pjFuIZNHGwuUV21SRPVpLncEaCoekX0xO+8ImjyoRuLiC7AbQsZJq5PXA3Qcuu
SPBCXEu+DMo4DIAIOgWBFmA7irxZSiuvD6Yt5Hj+o7qMCi9VoWo5dv37/TSKWgKz
sUMN6S1YHTkouT69qO9HlOemhdsf+ArmB3MAEfi+SsQ1+MtWzpJQT+DhZYjNT5fO
YD336zXosW+2rhaRbXYdVYeCQ02PfgfSFVfgV1/lZuq6filPUoFpCdmCls8Nwsdm
bZvV/u2/bmfznUYyw5YwLHYpdHvzWs1d9fOZacVBKEc7+ndBHTdzEt1USBv7+ltU
GL2qBm0qFLBmplKGHsRwxlXWNQ9lyqZ+Efp347qX9KQvPIx8eAAS4Fd9p+C6yf8l
Z5CZP32n01t6C6Y/2LBTuduK6Xfxma7P+MboXdsl/NKsR+7zl1+TgMPuyO+98QSt
G5jjeUCcLPlLp5bTuDB0GRw6OmrCCl3CbxnGZ7ep4nKU8g9O/+cKqtiPFuQJEefx
uc6V07ks8uEM3u60osIjJKObqbwLdkqVlENGLVEAlfcDUeeUutg9RS2CCzdlda9Q
5BZ+Vq03TI0ayJhiwAn4oC3Ox7eSpMkx7J7STWpM23sCWIm4/9RU9wqyDRInf+3f
VYbApuIBzB1H27HkiD6BErqGtwUaV5r07vYHrYYi0lFGkRSI5Nk20VzYNLeyc7mz
VRlgUu3ZZ9e9ABW/slOg48b/c3GN7RMiCMfWJSa8tZdW6wnM/g/JMR7gqVuHbfzZ
UCeeQHu4LWJ17adEJaK7zjMu/LtNVUjjRL5MrtftB/tj/3OUDorlak99B23cnp2J
vI0Hejv6yF1tbFzYN6HzWk+peBOr+BJN7kaFaVddb1/zHnse5xbJhRIgrQhVOu/E
ukJHkQYR5rdwSX4K5MGsooYw6gDWjcEPuJU0q+zpHHEXbWawS8vuj0Xj0SZPkmU0
fLq8y0LnZj9Xfmn6MT5c6/ZC66w8XtZhzFfigGCjVIord16WgQT0S4m4h7vLNEpG
1ElopLt44mMxW21+ZPRhJ1kKPXsiQtNVb3XQYfb7tCi8cdVSMldpTEl+M3hVcFTp
ATKIl2liqFMmfK5XfW4jmX/rO1agrUWWajIV4QzT9Nkcgrmj2rhKh/SeJxMS+w6R
CEru30a7JH9wxy16X0GHKpvWHCZbm8PmQD/0yRxHggPqGJYCmkwMu5jK47CqCStc
HidsVHxvrIuVLXSkWHOhZvkR7kM2ZDyh20gE4hTu93bSnTDB+qCIilTBiVtE54na
16i6+VHQTgeKQhjetZfBQO9U8y15Kj7YRzq27ICYTAR6e37reG5Q9d8vaqMrrNcU
LHuEWGn3ngxqrcPSKVHC30mv0X/nk9x56PPHYiwthTc50jY4iSHYrufQl11h//mG
GR4zPt1UZWNtrI9SlCVpRTZCn/g72gdLoL0iw8mhJ8YLDgeeXaObsv0XG1ktQcwd
7Dl5IsnaAYnridDi7aVQdtQUf70E4SpE6XjZ1JcJViWIwipTpP61ZdJSqIVzn6L3
bLJ7CYaWpfv8n2JeOtu5Ybfi4uQ0Y2TujJIJXtEgDw5CI/F57I8Q3y4UepXQsjGQ
wAwcC6yB8iofjp0CKKwO7vS4Zibc+F+6wzjhCHqRAmEcjcWHPKOewhIcEy9bdMGU
BfPJMahgBm5ThH8DLzf1LHcPjDuvjzI5aFze3U1ie5ZA5pw98XeWW3ErPuqayg/m
Yo3UPf4EP42TP3Err0UhqSM9W00IxDh/TxURxrBxOS0A0fO2s+K4+cm0h60Wf1QZ
ogPY2GddvArksGpvNbkCCuXTtZXiSAK+mAa8NmgTgyegaXQLwsGXAI/tMqghTjxS
oN0arHtY0XjFA3bDrNN9IVOgX1O+3gYX8qPkVydjP/2ZXiEc/8JDqXAKrpuaoJx9
XNNConleak1VsoOXOaTY+vsaCvcgYqqoexML6Prwb9pIXqxFGxQuN2tDeob2Ica5
qtJDsMfn/0xj7YpbGIcz3IevUy1htpbL7WL/nsxGaFZpg0YA07KZ8u7DGnPxJ3VJ
VNIjgGcU0JCTX51S+Hot4d2jYfsGNo574ekUEYRHQlINcfPvb0OZpPk9xEPfODsb
fBf3UYswHkH2ahmNKpaWI+5XljJSh6dOVBIe/7OgJmEKjvGXgiqUmO6NulPHhRUu
KQGUyaLpYthqwhP0owk6e80cNjjs3nOGh5rncEYUvjx6kKQNdOIBa211U5PnyXLt
WKCzE8BoODW/zXAwgvWlXJk9/x+3jEllZhlF3FEEa5Dt0FZ68+pgpc5kOqh7u9jK
PSThpNE5VPLdsFNc5K5yoiqLYLIONhziFvvsWe0Vk86nzvVuZ1DCtywPO6n/skfG
KUbddRVPFaNSAaBEQBXszBa4InDi9jAmN7LRWKijKhkY0hQDzOjE7JR+h3cOyeJh
gPJ+K67uWgIbF5a1FMv923cf2+9oCtygpuvhfUb91IRsdbZfTGmgIa0TKwFVp83t
FyqiUf5BfUIf+WWZLb840Vpsy9NC36qCwxpeeJXHblMN3fs7ahZDcEZ50YpKFtrG
cVx0mEz8dTw5hbO0SodUgJL4syXC8wHJnBbAwz/b8QQT5GjtHyhG9j7zpeU12G+y
voBuHQtnlyxzSgBV9wDmNguvhO8JgCHBmHIgSooWa5pF3HDUwZCZQ1FNx2VSbv3N
9/HE5NaXcMFVInNwJL5FpVjjxpGLgrYvhJ9XDPLtsU8NbC6B5rilAYZBaj+MMaep
y6AcDopRHaRlAlMcTdZiFQ7WPmQFECdtWQ8EBCiEHnfgSP7JEPQXqPZmoVI2xoGI
U1FXBE49nN7qj3ZIpf5eD54MxmWk+b7C8LuLmdLslnuN8LqGA+rNViKem3cn1lDG
V6cTOOn0Y+GDV2Oy/9XHiCO+xT74cRU6ePVGWEmNiZKsQX95xwr8wqVpSEO3GGot
MAnqaDmLjCLItIxujcI0kVTfBzMdHj+QdHB1Gz0rxnJPxJfYx9RzooTck4eaTogB
+ea613OL47+nFWhgPhbBbn5MSsIh9iHVpCthELF/z5cUwIAiBKpM0ZvWRMTu65Qx
97rumLR6zBUeSUHb3wX5iDkFA+fZ+EIxtMXfFA6TgFfqSd//ZhBdJg4XaHwKIzZF
s0+P+4BcALyL/RaeJdJZ/K4GyitjlohrYLgxLbtLluv+tWHCcNmTUprffqoQiXr4
DVrz/B7U5WuILkHapF0pRs2ETjBWK0gCDhQZKYtWnYKDTrfEiGY7iVVZTW4PX+sD
nbDzFr9zrpXcKoYqYmC6IJ5lVLYfHqpI3Mq8ZPxiby3K8j92rcAynMLoK3596uuf
U+A/9NXvshn0wIW40zIIEaVUJVs/pyItAMKSZheGHsrj0TETXYsRQuLl1EOaCdAV
prT64aO3dE0QYUjwkc+9Yo8V1BUWk6BVd5L3ICC0vJtfHzrMMOM2FTdFUmxFL42u
nr37D+iqZMtfAwI3jVMvio+LOcGSJAXd3PZLek8paIWqojpgkQyXyuuOTQslCfx0
KVBEwUMalBQZIkNxH2E7Db0oGaNQgWwwzKRlLp1NB0BIR+Mavhr3W5coQ5ZQRWne
OM+Af2Xmtq/zy3ciq03w7fhK0ykUHwzlyFggvT7Z0akN5JghlmmaXVjzhfseiZ+7
AHQTjnGn+hSetiiAQD9HUZ9izXhwe1GhZ+A2g6hEQ+WzkaDo0KjTOjWBnf6arM1f
CFMVa7DRWUD67jmsLy4e2JMwTNQlaqWPOc+ZsJ10UswWBcyi0IyhvoeUlYrPlKo3
i9zMOO4Dlqngs8ZflIWIH0+nbAgPrJ7QAOPN2W6VulVtETfG0Ls25nlK2iCaSKM5
QJI1sbkRnGi83npH9wcsPz2DqCxBKZ0VZMtt2qCr769tm3opASH6bs5u6MiRuR31
cUokPMN+OteD/NfEbY4rAkovIT/WJt1B7NdfVsx/L9MlHKVOTOcMQhS7OGLYTNi7
rL/FOUcSH4eRrVEHDANn+9XHDiDdlhajfWZROkoKF0Z1sZhmtbuf862JP2yIdfnZ
jF+kkbSDkTsj1lgbrWVCNh1b05i7NpsP2OBgpz+qF4JjLA2kGq0FyhPbZwfnw8EV
9vhtNE8U9JhGlffzkxnyzjCwEEDiirUk76tiF90esxpHh8vLRKHBK8UsRfnetJ14
lJ5t0EcCqJgQC/5VMhmROcAaV1o2MXZOJO+qzjFxuhbr/ryAGHB70vGVUIaZ9vk+
6ACsF1/05JlIRCve4pASCYMZqr/mkpcHiYG3PJZkcCeVZ4ecNC0zTH/f/96QmRWV
5LViwqFEGEHeWGI58/ZUeY39x9XYmfO7RNHfZm9+XxWI5olqEyRPJj8athBN0Qwz
OHlLMJWlEa3LQPy0NrIYgqeKODdMo8/lqedf9fxr5EY9FDARwMMXQlxfBXHZnQww
XvuTizun0HQZpL8gcqM7CJXpXRt/cX1Rt6ZDWCwMn5dbBkg87Oedd8COplNPQPIS
oYHXiYyzsehf6C8dYlHLMuLg6+j9MLA/QWi2Nu8ONVEJrwNp7+AaSzwBX8HC9W1E
9F2gi9SALArcMLHErrzFth18asrLbALUG4H4HOWP/UusZZ8eSI0PnoD/T8YMm+3i
foi5Yf4b6swFhVtJkgy43A1RZh+PrOUS7KBFHBB2w8OHepodKC6TKZvdgoAVBCrH
UfxVz8tM8+q5q2M+oXkfeEuwI/1/GX+etTuDuPzqF07ET88KqFd2KLNBwo35HNmS
TUQQOeUr+Gyww64WweAI46nB067VMX8RRgNXUPLM2goHumaVK1KRXpIITcBOr9vm
22lUrBbWLyhXCQxGOAVhabn4Hks76Ib27y+e7Of7LYaVLzNz+UPKXlLXPwex81YZ
SNnMyr7ylpC4BU1NBb4f0+e+czrOZGpbmCuppS8kLMcUsSzV5uvJANMkz26mnETq
Zilip6mM/FXh59fONXMBheTvevUajncjI6phw1+9+J1n5eGAcCyOlriAWJlGatK/
Bjy1AWflUGaa04J+Ja1m9JXW7/RNQCJCRSL/RmCbFtEyfdHdqpfy9km+VFCx5ulX
bY45D1P6FCDKYLAx/ElIP6NIEe/CKfGtuEZ7xYOfox+KzQ+EAt5NJVzlBQr9WJe8
cWlC2nChv+M1Qo++r76006ElhTeUqhD6RUN/FIWK5aFO2dU88Z07tfyB4O/r41Ae
fWhHS0r6xuZYZWI4Q5V2YsEtgZYXukcPi7gNq4PfR5l6XVAXS7fBVICqqFIvQp39
zWATVPcS+ODOhiKGRtQhlQgjkvVWxgtSVZm9kmb31Gi1vWYvvXcVDxYAeSNz14kY
3GgPgD0ESC96trRmo2xLiZSGX7k52V/TlK6v7muVVWAmu5LMzG4k0Z7rrmUgjczx
q+v+C+Ec3Jvadhrw+B+tCRbrw1XXuEuRG7OOl5s4O+Gkg2lLNBicjDHm7uijuIHx
8A4pqumOyajXm25MHarv1XP93qq8RrTT6y4Aa7XzxiPvbgYdbP/mRV6yKLUd7p6P
mAh+xcK6UReS8jHdqhonWrHsYssYYcium84q7uhMdsncNR83NBokL4kztO6+iQhR
gpUpu15N1Pcrvco4IXybjqeU99iAv/KOc2kgQ3nETtq36CQd0CGUZEhX0yMfDwD3
7iJ14TqGa50Nt7JwOh3EUzM2hUN81FAmg4ffyLMVmU57iW6evJtj2efBlxhzjfKj
Di6QWdc62fUnU7687b6UgUYJW+Q0TNmdhkj+VAze47WGKC36Qc1u9iWYCitYEBtF
+NWPMABALdIGDSUleG2hIQHjVKGryKneM4P035yjP2kaXbTmvFFwlflhqUyutd6l
UgVcgdmjHYOHgTZ3s9ZG24c5i2o1F2AbV/YU5mWclGypl6oz/OXHcTyjuc5fm4dH
lxEnae/AUeTEuyftZ+UxvzYcy8yp2Y9vsACZTpuNv8rEn4nyPAwT1EzemkW3G0xi
Bi6SZeIS0uUWZsZBJVf234avhozrSDm2yQgA0uPje19/UVTlJ9ykxQ4gGcN3fIU0
sUAi1kAcA2Z7LU8H8gsSgM8THUme3gtmwSiAfQEsjg/hH0oeykX2MEKUBtOcUj/E
mFpnuDLhzegCKQLtkZlmqyaIC1kQDu+jjs2ekAdWFuQV6+vjwn2mCaVXXFEVwv/8
L9OcKCIjHesW+b2Iga7URMG9Lp/S8lQpvLZ01Zn1wNIfCv/RhfUMqC1SEA01+0MX
nnFLPPhEH8ngn0PoBpva/c+Jl7HvUTG1c8R6/spEp2vhtoMbPilchS3iWUKeRt9U
o4EVaKc/xigEwXwwB5SJ9k6xUqxIzpqj2kkMgpMHIhEgPl/RDUevfh2FligsVi8H
hEEOS+2uYXeNruA1dArAVu6W7Ly5BwTmJsBL7tlEhJcclgDfUL2yqyrA1UP4Ci8z
ynFUBtF4DNPJoUskgZmVM9fud4jrN9lT/WZK/sG5MdIRIHj+FYf6XRIxLw1ct/1P
VniicbPSoUOB2T/cX9+bDJQrEy255okqLkpU8cNMJQRNd7baUahLoqxQATHX9HoH
QcfXv5SqYi5E96V/J8Ab9b4qJImcVMODR/VXul2y60xDBNdPdNQYb5ul0A+OpgcH
iqugwekuElk6iIhutK4I5V0I8elYbrB46/D7tzOklKqdLCvskqqSgC1LH7S2JEHd
1OizkarvrGm4FA0KreI+vln+4SCZQ4nVlqJW5d7SfoJnxbydXybb5A5b5h34Q/R6
zofNGjYZ9BEE3qHiFg+uPTgSOr6wcaoiOv7f7s/rMjyujiJvigpusAXIJaMNDgpL
qstVkrytA3gbuySyE8RKtq3JbQU72e579Xqp5uYQTPKrJLwRYG9CZ+IoDH4OVlN/
9KPZv8g+JQ6Ew62bPQPFy3rXtZk0RgKXMIdQmwItLS904MIj0zhcaRSX3S8oQ4yS
eJRxt85NxsDDfBvl4O2Lu50CT0Y6Hla+CEoWjwOa5PA4/L9bgViIour5nsQvzED+
HLJ4U3ifuMLNqpHMeZpA7S3z2wO7650oyHVAJzC/1dfRckbHFbva9M4mEKjQQbO/
ijTe98CXFwyF7L4t2KOzLegvqm+8GXG2TGYreaX2nw48xbsXNsXNryrRhPGFTMmQ
eZMbiVOUKNiaDtyoywFaNr/dZ9AWIdttI+88JNXcnQAmrMd7xFTQpCnwB/sj50jd
9DZq9ZkXgrseZslLI0UUknlG7FHctRpkAxJgEpN2x35mAjJ5YrSH7JjgdTE22suA
WO6kNTIQFO8d0+qhp92REx/xBPy5RMlUFvteLDFJiDw2z+l84cpy0WGAkQvSq5cj
42IuwUVp7QYen/VLNGDTuZA7jC/DnX7Y9/77OmnezmR2PBM34J2pDUTsYFob2BlU
pi+lpxTbP76/rLO/sz2F4ljnmCyrI3Sh37e6X7rJgzKz5m4f6m8AiiA6+TD7b8Oq
CThAI2sbva2d2QofsZ4Waj4GBrs0q2E58oh2hfTKsIgOKni5fsTblKISvU3py26N
KEEB5WUsJho/4C/4d7Yo/U1rctvwanKFff8hNaOZiRfGerdycR/yyB5lGvMv6Eo7
iLjMrCUJZGB8MSX+FN1JFArVUmFuOJGg2nQlf4tWRPKODs1F6AVUREg7jdV5oU4S
uzWsVSyf5MaVjji9tRV3+jYhqRt5VTFHiDCnq1myJaEoNj1EuQSYZru1HJ7GnNqA
rs0pVj4a3VhAaKnQoe7EIoFyFXy9fvz/S3GsYbqGzEXuyb2sjsudFj50CauhUiNK
6NJXrGfcFBztvIDb4QBMwr4gMQN5Xaslw65gP/Wr89ZYrZ0pk76T3ukqfdwWAN8E
6RTe0tUsoFsk7sb0z40V/knhXWr5bilBIbnJmVbx1I92BtClV86Sf5aUHbfqCUe3
KDKu2eGyDMHTaJRmwDQ+gwH7vl06tCYyrYRdZ8HajLsLz04SdO4+qtQlH3YPyoy9
G6dQUyieOuzzOPPJjlPYnoQQhXUyFnv8uzQ9BoHv2qmXFQI6E0gblljY3i7UPher
z9GRSpaQYmGYQTGg1wLZ15TFQyIOYypZzV3CfpVtx2JxOySOwbEZz7NTTehEwxWr
xJrxzrra8yXxPLRsZbbgbsP9Y/rAYW90TsSEV7AGVCLVV/81h1b7b4ym47pKWOAv
tzDi3DOLkb4N6qpIkcW3g/GGAqrNbYX9izc7a/mnNb3gEi238koyUJgIIWSbDANI
BuE/RX2W1QZ1X8N4cRzoWpbz5OCRjaEhGbQTNHjSUu2loRK00h11N43NQH+1OPwi
jO1MRathANDhaxsJJ1gqKLYTlyGtzwVSeRSyqnVjK4TGhTm8alh/9ATyZTnj/32S
ry4fSFdj6oNShXox+uBGAV4DET4XHmj//TX0+mzgApBZgQuhD0UmHbhA9zNbfBqx
TZu+VZiSaSI4kbIpSFiOJDYhbu8QoprnQsmO1k3B2yBZzMTmdLK2wB5Z8klIABWu
MGwrhQQyfJ9HTgHHgbZaZyF68Rzb9j+06clTxtgz8K0B17Wlt6Ks0n4Pd5h39zjN
k5sbptscyFNc526eZHSXvGJRpZ48lC91UH+FQGN4fVGKIvLnXi3KPY6AwCkozo9L
H0FlO1dMWEqLtCZHR9tasd133bBPW2xHXMtjDQPlTo4z5+QbplU13fRs+x0BT+or
/Doe3ItbzQRr+18cRVymTw53QMocLsPDq+v/ZCS9+A6zGCUcKrxnZipOTl1WRCOZ
H1ubtjW2QjN9YsW6T/M99LhmUHq+3rtFyC2qSKOZDOnmrVG7SHWiKkp3JpFtMnIF
TEOJMquZHoKOgVtvFi+0xNW6RPmPQUfD9CvaRoTlCyknkCWiyoYkGUR/huoAFL9g
iVybPA+C6Z7fowb9ZqSzJic2k3jj5As3uHR4I7O2/YyyRpx0tIOhEgKB5IQNEMgg
/bwj5QNEfUbrlS/nPCFbNkrGKPLavAjRaE2C7UJOM4SZ6PfxPjW2poctZ/R6mInB
6kSKLJukA7NDgiDS6cYtn3V1cCFNgDJeHTuagRk2PVmicnWlq/4ybLwfCzNgZJ7m
jKcBYYFFOu5iNv7Ok9UvmmBkvSC5FlE8q2TESz+YaETXjXpm3kAer5Y4L7MPsQc9
IDxWwLOQfitjiEBUJHDMnw05R3FkueacyKU5w0pJSOEcJ3VDW8h5l/tjKopCi/YD
oXVeTCgexUZkK2D/fLsMI3EfpzHzUoosPg7gHTh6r3CnpMNZEGwa4ils+wW9tvjc
m1+ebnKmL5ENP1Nra/TSOHZJEtxNt9mMhWN4/ov7thG3E50WCAQ0J1VXlekADzf9
f7CWYAiEBQJ71H06tbaKpYbF9f/pRpmgCerT//tk8GF1Z2NEqwktzKe+A6AImDbd
Jz/AyEtqh6IxOpaGMxrQRiR5gcBJqGr1qN9idH5TVKZEg6O+W315AXQXRm089cwV
+ZTvOnlg1akUxgjeHOwY/72Q7dJNz7+yghb2evklMFfE3rvcDbnaFpeF5AgTvSYj
NJ2ZFStOM7etnireb2jH5of+TYMLpe+Ck4EXl7Y/yvy2oWoyjGfEhBUL21nwb5F1
FDqJpg7Z/hFpS0oVlUtE7IZCsM78oLk5o3LVPNZJTsEdRmaOeW8lClloTMLmm8pY
umq4fMWPZwzxtV8P33zXqAMTNvCey2iWZrrN5nXmYRlwrz1B+fJsa4tF1DOlHD1O
umsScWn0SFqt7e7IKmxuDbOqCSnXqPEiDmxlUlM4P61pvaDkKRf9ptHHWeXxxi7K
KPIpCnUH6ywlyI6hzK9IWlCZ1kv+QuYOrQKhSHamjUJNg5m1UZMwgbn4r8xc2qxQ
Z5zSOS7VWRC/iAWQTB6yiCIW+qn1uRdHs8ztSEdLAlaNiU0UvrV+X+GWt2jDpY2x
C73RlHV58kMIeokIIQsDbgf/owC6TQyV9wnyB4s1SGQuAFA13JUn3w9Swnb7t5Jt
XGt9vCjiGXBLnh7Vva+6u+gR18vx+FuW3ZJEDIjhvybKpfKn4e04I3KKtAkWQ3Ef
R3+/lTc/TS7dt9nhzWWb8W1au0SPeyBQm+C4Btsc10+vnuPSrlwyWRyPWZ/7ySCS
5CoFpk1ysV5vCpYgMdepLDTXFcGi2wqdnRffBcgz6lF2S9ibgU+DxLVVcBFVvU5i
4TT2Ybc6ROiU5RLy9x/fIm+PZ9s1Yd+c/cqT+oZjCEw9yWxtlUqk45PKsNOzvuti
Kf7HM2LBKYHKxGBaeuQG4KHhdkq/SFuZoJUf8tM1BwG8KgPASFLC7Tlsvt2YegYb
A1hGg7wpomQy1AXmeiWalnYpTstogrtf7lJU/sF44U45iXcgSOE8+3yNrV0zElwM
rLyeI9AlTlwkM5Fm7lxHbqbt3V5K6c98JHd/6A60fBBbTmlXkQxh0/V0En3fGrep
R910wq2u45iBbAE4WeGN21bPajRuL822nF0K4YoyPZVJvppItwYHf8gNoDhqUHlE
uAlTP2HBL7wRTS7zkqLPPsciwPFfkEUAQT9c5hIWhdEmeDgHj8b77bYW+d9J2ykN
/3TOVZsaT3wUc13xHhtwLUM+VrYv/hMVFYt71ATPC/XgqOUs45JD9FnbxMNFM0yT
p1gRK2l21OEbV7hOyy0Y/dtT+Ed7/71tuXmFe949U4amxfcoIm8opRI+e2q7E50u
d7B9I69CmryCE0OTC4OmM2kjZVDefqkkyvDW7njv/4V0HRTw6SlduAcB/fo/fEls
zpXNISAA6v02CUt2fY/kUuWikEft5lG4bSjGVvPvdRPDz1BXzbqBtxi9sWm80raU
DzCWonkBM5JPaCO6mBtsK9b8I08SIqVb81m/2faNUUDEC0rNCeJnjpxjVmxfwHsH
+gzWd3e+HCIEFbIkht59fgI1hJXy7qf0QlaCwHC+Yh6321vJ6sro+t6AcuKFpIhi
1ys1b6X9S5G0rb0yDb30ow3k8ACeJbHanSDFV/bsh9EXi4qLu9xNPox9EW0/7me0
lrU+yGkzll3OlPYrnoZrU8+vKAbIrPOzt//kuE3FD8w1AKu41toNL89F1F/AezfC
OPQoC2ca8wZtGXw9UGK+7lwLnQtUpUgQMsjGtrmwWMw2ZqR3RqHXXtI9N1MVa1lc
RTAD+ZduPbaRe6zpGQuLxw1ONgefHEspibEugXFYXDHQ7Dk7tirdvwZCNmWS071t
eYjbNuXvqCDWY6wxycb9qol3/Nr1pnnoY2I/iuma8jitllrDQhcVQJtw91mahIjJ
uyPPR5MGO8SaGU9sKO9YuhsVX8S+wj1VTi6b4gpjfjZQWN/v99sA6V8asyypGlt+
Je2NW+7S+nBR+TkUOpLZr67VFeE0yKi1Sl0zV8I9cXLjoHzenQ15Tko5Xt07uH4L
6BVZ7+Yx5hkGABG+lEE8sHHimzxMntqQqbXiVamhuqze55JH2apFPjeS30BngODw
VqS9I+vASmni7x3pUQvJPMJMN5EMD04o7a/oFx1IBaEF2nFtznz8yVsfpIJcQTUi
0lG39SjuZKkfuyzTUwhwM2KVcI16F+9/yZV42Nwa64AZCbn6twk76UiFSmFp4SZw
RG4rjm1FF6PARvGVCDnMCFmP1WtfUOPIeflJ9NYrK36ywoeqnN0ZOXHbpvpw2dCf
ZpXCpsW78IltL67tf/5bk9SQ6f91aS2HwJN1zq0pOC12Oq+NyYoermwn5cL4bAKc
cf2WxXbk/Gr9o7orxVZYQ5Vqm8cT6TicpacwQnoBJT7okYOMABSz694DIeQbsdDK
37dmhhlXxmjiogSWW0HSJpGqsllbSfCXC5zoynKZFSNHHGYLTmEj7xC+QdVHGNtk
suh+i3KkjUilKgwZD26AXHY4fNxwkFQGmDEHg+vUsjrH4Qa/IJX08i7ijCFob6XO
6I1yH79MFSrAjqPzzfKP2usmMDiIkOmtzXnIRZ+i1WLtSylYOWI+FSfMkzMGvYe3
QCtt7AGBa25ABYNlnaztjrKvjGSPYVfpC5YIxberJpn5q3MBa/ravPCOi4+z5Q3U
FJ8bO8VdPZzz8o+z1aYEMZ3zs81vnt/jsIpFU2qFoezBw/8GNbOoa0PbAVSEjxlN
FGgaTY8u6CudxnjFvkCOSpiCuMnadVErxsbCxWJeehXgjudpmDtefDnteW+lf/P9
qid10p4GEuF/6ywoJg7Pu4vROKotLUEBAN963SFEQzvOspAkXtvhgwo7u8EMfPNr
xvguufIe3Jrm0fPocida2rrYG7q3fzcX4Q/1CEjDnwMFCdxnHURG8HI1a1KXA130
5jmNFU4Da48CEQCeqSlJb6cLQpRSk2CdIP1bBywETuegjsAIRtsjgfgCBL9uA3Qw
GyVVxcdYHfbtZyFozTa+dbMqfTEWpeFBop8sfG6XFcPotM2dJCGpEdPTus5LOQwE
DCpiiuq4H/WMbRZR+qOMVB9v9tE2Slz2eLXGSoGHh65x3uxhrf2mZTtWy9N5DzUo
/SENF/NzM3j578BePxcv69eeIdK0OFZbt9ZU2o9whrkuP1FHKtAow4SyyimmUVsL
I7gMKIooxlBF2Oi/dUA1dLO8EUi+mBxBrgtA5dBQ3vDMlf17BVEJRJwroZoiOcI4
LXCbuvxiiPmQk6j8PEa0EvLYTMFi39wzs+wlZwPuAsuk4TGTIBEl7W+s6VieTj10
ASsftdDsECNg4zK9RmueOUjoMnEst6sbxD2Tq/PGNTDJ35d7EqLltqXtrfQJ4X+N
cWPkdyPp/kyCakXcTWKr3+CCQsi5RuHk+qOzosBZn6HxwS33sQnNT5wFYC+d3i1J
WIKtF80PNFs4JX3EJEc+1En6rwmkSaF3wXoNQWh/Tsuq4yZcbcJI1BkkIztMliEu
yTBFBXa5r2hTUfbsfqF38b6xVp5SENPid4hYhe2Bn3VcgdB5ZLxeVPgBeTvwvWAm
jqubLKCI+WRAeN5affEw12I9dVQbNaDv3ER+Xd5BaBvXa0ZIcJrw78JNSVEnPAfu
iH+Gpm44LPYjp/Iq8qOlugI8kKZAl6WZIXfGqRWRVPnDldbr3NLw76hzrusZL1QP
8Kz2NrgARsty4Rqp70qoOrJxJh9OcRXFnMg2ob2kaTUEBzzN/ugMeZbPSV8V3BHa
Vo+PafQWfYF7jsVOl9xGSrdnqSCrEWXcBKkoSyiUK+mYra/GKZJvICIuVQJSPHdi
bMWD8LkOcXyaHYvHdEP7I9uMGqPdMKGanFNu5Na4ZNE1uWAE9FivP1Ratch3Uqte
vmz7ObM3MFs0Ig+XnXQxNDF7gMGFhBH2F9N74CdseB28+Uo+CJLxulhGzNS2cOh6
TOm2PZObvkFlULwI9jlAjE7/V8O0afOQO5ykt57yLNZpzYRcAbpFwHHaw6lMeGWN
uQWKPqcbHM00QhNDyhUrTSoy0zrvmowuy516QYeihvdCipP9l3d+S95kFDor+1p4
mYAfz4eR/4GZySrIWtCLz8zNhme0M13TP2dJdu3B9Znd7C+ysDW/oTlL1e+9fZZg
8VdnJWAJjxWT/oRgKIim4qR8MZiiygMldkS7x5VOLaLOlDh2E53rhEfuENiv/MOG
+CJiJuIFH0YFkuf03QdCwZL55x5PhoPcaHpifY/RNfwZiJmkIpJE1yK5JLEB8vVV
kGUuigC/YlV+TjZI3i/uMrGEakeqzZNkhm4vwQM/HdlJCQFpWqBvvAZvyzcO1Ihw
XN6Hccm1QGQhG9AtBW2NT/h4J8aKI8z2q3FkVrZIvFiEm30YGfbV0F6irEQgImal
JeVU1l2zf6gW2dRveMy+eABz+cUlgQcg0Do39FgY1G26+8THWm1CYWacTFMeypuU
xV3+UPaqYdvmwYNXFL6Xig0QRB8FCWqvh9nP2K4daTa6DIUB0ab+FN/EkHkPALkB
OK4nCzSgope4fD2L5dpRbiDtKDB8yLTPEqo82AW21CnWiNvKKtD2y5NQbSVlFaQF
llL06HdHBQdg5uChT9Nh7OEd7vHmq/ukGWPF/R1KqEOQXMkUSY6nWK2qdJHJhLn2
sgJeTibcQ7M+qbhf4YHyAgBLdEjRdk42Ge/mKmrcXNlGGFgv8qI5RhlHIpJzoyhk
DyJTcUlUiF/+x28nDycUgKHhBCXKeg9IV+2mIWrqHcg+3t+yAf7tUPlUJCm0nHoU
8wXAsysLyx69ywesIHyTkDfXU1awmEd76l8Apm/45XGK3w6jC+lU/D1h9h0MsJ19
cSD6pK1I9gK8q3oWbeNcgV+S9eIpLJRqT0CeDLNfkGp33Xm/eTkGr/DNaQC7JNCy
Z/oH4yEz2L2RnXwica7vGIYbKO3d5bbnv82CCPaoQScKsmnpW+rfnMO/3G0UFsVP
pIouaLTBkl4LtzEOvBJDkAPqis1md1k+HhvUPtvtIMqWOEHS0CwicD/BPPlvZNDc
kmLCr+FE8ej3m1XC+2riWzr8AnWPqYpsGq+WhatQ+htc9nG1Ds3Qf2tCOHlmtQr5
6V0xrQUati/gOC8368OBcAxGWVAVLyuQDutki8Vs/AxQ73ztThdDOgvOF/OlSggQ
NzC6cobpAvNWoVK7XyO2oB7WiBJh9j06khqEdbO8GR+laS/g+n5uoAN0lBy/DDCH
E3Md1+KQJO+96I2voOwo/09RhuuAzKvg39fXNqHy19A0IbqbOTQiYtfVJxIurdja
///gmaosDBrlStdBY7X5TxJiM3WgecNYRwwLpTbMhL9FlIxKkFZcAIimMRU03rsb
pmNALKgNtwRbFR77nX2tf/mRzkKNxJQ30FK7t3z6p0UZFN5MvJn+zOpbboEqI6Br
oJtYgg+26QxGSZRjJyW/UTPyq0j6QvK5qbXZh+3M9MLJIsvHFK9Fx2b51sKfogmW
L9CcWB3lUJYysS3yU3+gVUJ6lIUKRtV9MdIZpnAvktJdxCuQETRt9V1ezNS4elDt
LfeLFVJUqCW3aOZrhyoVBSt1Mvx9AY9qQANCcfOCzWjArarLyuUwjZGsMWTDxMOM
Km8QYY9Z/Po4EqMGE5MX5h1YI5x+bzEFkrFkgUUmr3Opcz4yP6Ma5LLdSkv4jkMY
SR5gfoc/u2gB+jSFRzwRlHmbMs0V+hIp+b4X8hps0/T0ix9Z8b+R4x69kCAoSVnY
RKpGc2ZQ4qYq4GHrbXYgu2kJzwqJW14+mmJJWPhc+XRrJBrEIRF3d+mWR/mBXuuZ
bRR9cGYRboO4XSZOEc0Phn5crYLt1H6grmoD+lP8Xb59Yi+xQ7VTLJWh1LwqHbUi
ELiYmBf3wCfH8bb9mhu4lJIbM9xLh5v3AIGNxJhfYdudEiWDquewcUpQp6kdwMiZ
izvCmlKq9Cguk4pSRTjsVBZOq8oN5DCmjfayTFx7vG22LY2gMLLDYDxj6fEmxdlY
CUdbxE/sZd1xqxg2ZIgftx+SU3WNiGIRW+h6Q8l28s/GSPLD8TdSeEt5YNZePbSo
qlVkb0qoqeZX7hV0qMWp47J4EmRONaN5snX9d0TjKVlY0O9DYUO1GvouPthpb96W
UxQON9S6pPXfCDXXQkHliTgMRl29ByzOESOUEujBtVEBycEvkORgtKep4lUsnm7c
S659z8W/SCFZ1P5Vu8R+e0CoQHaC69/GC6zmqiYFrS5Fy2J1rqVpFsPlCi0tmMVT
6p3T7xthQldg9yuiEYmv1STvtzFj7KKtcZTZrU44zOhbsWfNWJpFqiQfjzq3lo09
xFUxBmbxuquxoWfQ1q80a1NCGBsXHv3plIo8nGbkxA1R3JEXt1XJoNczMy6aJGcu
SGAYhl4TE5wUYuB7Sxo8LPYyjKE2CKEEo90LS343pxxlQv24vj5XvwqWF3Snvs/n
G4iuBqUjbz/5lZsNh5sqW7MX6DBGrtG/TJP+p/qr3vOWcCykatj0cxEHhf9THgEh
ljbYnjZTN5x8jRga38nDSmv25GxvyKr8P98V1WW53/IVqu04i25Nu6TWW6ngVTis
cOo+CJpTAcGg7qb1hv5l7P0Iz6X2rIJzMLKDz8RMaMj9G639Bdz/InxCMaU0rQrX
e6QllCEqanVpS9iZ2UpxIrqKOxT6oq/4/ru+dFhUrcwVAk84YsbHrqrbJEZd4d0+
nVcSBk6mzjjCuJwk5afcxR9iAxBx7Fg16yOd38308mIH4EkQcOYosEpdhTV6tLq+
nMird/Bb76XSGcH88RAbMjmTApCRF/qFNu+FO8QDmHRuo5nUWhYMt5YC2DmfE3xn
lhS6XH0oplp+5oH+LHpFoMDPBGXY4G0b+E7P1XtTDXDcyXVoYvHHpTp7Mnib0tc9
MaaAMv3T9vJ5I7stoGHjGOfCp60/Yu3LOCWSm97BlaVxH/WAqfzJIUpkmcBrGvUB
As7yIMvI6wyWNPPR2JdJIzvVpScIN1UMgx97d5YXuC4gF3mtgVSHAAlM+iyihXrd
/jPxg2CGfL2USnslsRz1IJIbcibnL6L4iaOWX78g4WLL2XLQ8L1ra+g89b9zzJdt
BEt5agZSnL9RPOqZa/rDhv2Fit4M10dycSlAcwUZ89PUqI0IDmKdgpltL7dWm+KB
VsrrLzZWenZqG4+EcKBx4zpWs1+NbYp4zOzek+2htkjec0LTXHkAKO/wPs/pe+p0
gfCe9SCWPN1gAbeus2dHja7nSXzjhF3azWLbtFAk88NfjdLJuWSATh3SqdmiwXVK
Yj6gd6924+dkMyr35xpCnvN8qliWc5O4M5xuAV7bnWEDkhZyFhsVpXJk98lDD44P
V9D15bpjAzE2Cg7HTTJJM6daKn/Ii9KKBlqI4+VYcrPs9ubq7Tzt+J3MTz8Jmtwm
HV1ti72z3pSnMGp0wezPjy4yO1MQhzCz0uFc2UOSvvylTjCE5UkFE9AmrUzxEFN4
0+SU7z/rBTdLCFWjGUZeT67TiDtjDjmJty+7xVUY+BJoNq5PjbVoqcffcGbxNAzH
tsgrO7sz4s2py7fw5bGM9r8IH6Qh9F2hmjJPz8/qj8UsxhNhZOdK14AG0M2trEwS
1T9FyWlm18uMQTkaUQac4Xiw34jBlDz6tFmzmFx4qq17QuK6dIePOJYkNVYJoZP6
33M0BUeWgzQ8bsdC46q5L/6yO6pnFaDlrSALXz9up5E3hx1d0ZsC7t54Hx8+agMp
goKK3E2v8FRINauHsM5i1UK2N0Dw8Sj+fGNRLRGFUT195tyQbWfAY5AN5wSer22D
fsZd1uphnYcdx1A75n18Iu4dkSe2s/eSd1WBF0+aSBjdTutxxvc9HcLKh2chee31
qQKVb0aP3M+60vu5egKXDVnsOii0ORMWPTBor0yeQTN7nZIMJZdcQ551Z9cFx5ed
PA6ACO0PeL0oaTEG2kvh0X25vcmgguS/LFcSanhk7QlS/uDRwMeW7p7r90pGO+U7
9ATFH5XLKck/my7TeI7kY80sWP8nvvLSf6wuYXFMZKrvbo/SodwAvW/cBEOqZMth
K//wwwfIJP1q1P7lxAdaJ7Adm2MfMIxEaGE/L9PJBkSO3mdyguc6eOUtxsasJ19A
We+rH6qkv+c9iILOXQ0qTx8Qvs88iAAOuJsry7NcrU90idzyQRCPOBE8p8hxlNbI
R16DBwntr8NtXqG5Uwpj5TpoFqmvIhThe052oh6hu2nCns9JMJX43oHmdvHyrSWC
Tte4ycmlAQL0O14U5X786iUS+9PWYyit6VzpqoQEHW7FQ0ZsKj+8EuQObEY+3+AF
UeQNeghn2AVPFpAmq9Sv0mkVnSzRtrKHSAfVzP8efmeAfsflVdHEzlR6WDbceZsM
5kfBBI3RD0uadsggY3N+ac9o0Cd+1M9xVKeN9H/2waZ6UB2QxQVLEEo3Ktz9IMPg
REmoi7AM4joOMpL7LMR3G2ZchHim5HXRF7wYw2aeUNMKQ9O7mdS+W+24RC9ayFJD
1jWyDG63l/9DQOOzh844vC6Z5pJRig/rWM1PQI1zdpuTABYIiVAhkIecJgo6kuOe
rfJF3KDVUN0AnPIVaXN9vPBtfyRpXezPdIkMhWfxccHHr3wGZ99s3BHipo77Dq46
cNTipwHYaVly1oDMNTk9Cny2iS/+8KVAIARf4RTnJxePFxKayHaSw62TOtaQjTJT
dtvg37Yj6HyroKcFXF5Cy9jH/WdNLjHcNmhiixzR9oZenNyQ059p4u9aAF0/27nb
jyzxWULdZviwifzZyXEWoROBupftBUoqPUgUWuVKTuOfcaI24AZ8CoWJy2f1Dht5
HgPOTgaOAMIF0diqoDL+/ne4P6lvFAuMbuX4Yh1GyUtg1sNvtMYMCRw++UFzpWAo
p7ReDoVp1FavYDMqmLk6Q1EXSIa8KRN4A+AdglS4mEtOvdgEUAHvY9csXh3aCH/X
HaPVMY8QAV+8aO0N6bzhv4/+U9dQVf1kcwyarp5BFIAPUC0j2bXpqDwQZegy7xgt
W9KSuMPKSZZyq1xRfVM+C7URpHpCfOjdrWDYE/gWon5SCck5sjjLtJuHwJ3KmPuO
5YTHTi5nfwyW8LxjdBYM2tGDheXc4nDIvcD7JQS0rn4Y6I65M2De/UHQ0sdh6Q2j
IgMa/va9zpVc2US1h6o7a2GiEC0l5cZkevzV0ag2lXnH+cwqJOuX7Pmv/Y1J7yMI
CpxUZinc7TpzKX/ELP18NCGlUZ/YJflyutcH+r4+CIV9k26jGJzDs4HcS5WDNFZc
zBO5dA/sN285xtsiBaQbh1tOl1xoDR2BKx+041m40MP8dV47ZHTOzr87TIot7Ez0
eRyioD1XcXQiSV3sgPN/RAQxdbv0KhHO+i+WX/itWDvihjL8bbm1m++pjUNzUS0M
llIakybNw11fOq9fDqYkpfXipMH6Yj+CPKL0rAhDIvHprID/5aCz/MWhqJfMhDut
CxExSUQINZ/Hj7JS4/ha3448jd85kc6Fc0QPUShGKdmDRt+TW4qhn5+yTyAANxoY
+WOdjEhdL0ntf3o7oeNceLqgK5vD90yqhbuBajgGyA0kFYnikp2Y39rbIwZ3ysrs
574ijAETCCB96EE45zR/5YIZZhTzo24bYVEfRymSFK+7WGQsTa14lU67mekO2rnr
VhRt2W6hOyLO3SdAr1cdTwHAOdWOzo6HTdyzFhJx+F3XOgQRaGUFsD3Pdm0W5cj+
PS92EwbMTOrW0JLewrSkos2Oz0FokHu2uFs6H3qP05/3Be2u9oBM0lsoqan4Wbgs
C3I70sodIZilCDwoBj8ur5aVVHdVxVmBeDfhJEmz4jJlC6Izeym/6a+LM++IRKFt
E++HrslZVOg3ifuXXLZBIsGY1dluaKgg02QO87DVqPmQ++3O0xmFLYxTy5C/HsC3
knu+9BBH6X+6XPrVHbxhW/OxBODawGETQFJk/tVo+ejWc74jBYyfT0thdexmzduy
rWYQXPhB114E3pnH9d1ilCrTG6GbRYGAij9FcKnw/KcJ+v0v6x8sfCSetyMa8VM7
oaQroqZtx0MWAjjztvgQNVxGtC7pe23UuovmVUDYZoP88/MwWGowGSHp8cKUlnHL
d/um0UQhaFxMWfj8WhpfchC9n3alnI8wqxLiGN4ZH5T8jsinfLhKaDOI54HX/KXQ
Pj1yXdLLbdXOQqy0/WEMojRVosjn+gX3DS0wL9Q7J+yFLtlCS+yXp4GdxVdsmjX0
lgNCJimETvoFE02DP09Vx71i96d1msxFT9zj8u2KXhMjB6ylhTm3J+0ngNRdBtAJ
mrrm1HfAWT2PPcor0ne052VdfnzlrmCqPf+yj0BV2JYIjn/LX+zdzuOzPpx7mHtE
hE6WC/Em58MqxzKxcaMQGxB934EgZy/44FGmG8paPsWk15d96jeKw7n5NClJLvF/
SvV3tY39tIfwtNnYjTikfqvBXJ+r9ahfkiPdvC4cL5friB0O6JKIQmkp/sWgzW5D
VPlRShPEmL4egNgPbDH5/SPDI0qHg1zE8Vo/5kwmVHY660pAL8K3AwCM/s7zMdQe
9n5PvyvSccIIw/B7yCFxG4S7m0UeDylJIc6gUAuOVzFeDJvdONIVDDixdb0AiefW
JU5AJjXAWfefet66q4+N6ze5tUpwj5Xh83h+shuM64hCbuVndRGhTunOaoaQx19J
Dfw4CkSShqvqtUUVGe66IpL2HU8eqU4mNwdMB17vM2h8Z/garZeOoxhS+iLrEfeu
/o1Q/blajvQNURV/WTvvS+aQliuh6empuM5c6sUzzPS1IWmSp8M3dkdDQVoLvQgN
0hqEnYt+apsMghdWP7+gUXQqpGI7Bb41dpRXZEYCfkHyzXkcEs91jG4d/uJMKnPq
IHjP405nfyle3k6Cmar0X/gAG4f6DgGOEXQGYRG5w4KXBKI6YSZ39uVEE1vKJGB4
i/x/5Rg6jxUwbl/rh3bB702uD3r74APcu9xCdYdsm4Xu1Xq8wjBK8pJx3trmvmXn
XtFcfagCvdeYfGRcr3n9OdIq+EK/xZlGTxLz2oCgH3Hiw0f2cicOX/yCnbGn3+xZ
Qb/KQ31rn+0Wq0Ol0Cdj5OKVC3Li8yFmKT8f+9DhWul9lFCrSx6S4N9QsVFSmUVZ
h6omf4BzJXGg4ZtqnsqiFSgGjbIJgDIts9G/XzG9wJ++Vq0k00H9H2FESt9SFo3k
3DRf2w7/xAlQQ4qZXtzuihyrwTW/ip//37Vqsxpj5nr4WJmKRMMdAw2byBtZD6Sx
dzVfpbFX+JPkfDH8KtPsdZL6BA9aMhf1KIDTrSnJjPHs1GTo+wHBQKjx3RLZQ0/a
xkqpDTc791hQc1HeiRJkLrfoozXel3pJpkoMctZKL+Ll5OxvsCdc/RgrW1ZzYjCo
Lyqx4eLFg90hp8c5lWJawbf6KDoZn0wsJMULW8ULmtRLzyes9casXOO8YmLP1aRS
MijeHcI7Zvz1liFrOU+lYbU6W11RbzS7R+jnqElerpC7KBK53PS+xQ2+sJAX0m64
U+02FMrQ2oKR/MPGqJNSNHhYe9nsaw/j6rlNrW1OBcjQAKQkERc9I/dD7yXOaWqR
MIzULWfxIHfb/LDYZKNM1ELavpl08OgFY2qMm7BwD5ke2TRAZ8Sl20jc+cviLulW
+u4OCE9QJjGkn4pdSupWn3pxOfpjm1gaxQknY9F8aqfDyxNF2K1xvmJWpwBpZ+Ab
CS/J8o+sDG+PJJSpPT6Dsgq1tsuB+7Zhn+iiSGhc0nB3/+yujV4/40Pbn9SoE6Yv
FXT0ge+GkHQPjhQB82NAtRsgcnjWCC8RoYJkz6WUnPnxIX5ApZYiho+dTxUEaI1l
KZOydEvrcd0SqXYTK6mGSqKDjlOlouYZLbLp0cCeIkHzpLYCo67xgCvRQFcZJLrl
nOtx3dTKNL3UM3VWIxL2mr6sEdcaS2ACwYyzBOzl16XF8K4Aow0xWceN85GXqbBT
ZCgBOh86T+Oh68bW3akgaFhJXBvz+czc2f3UmzHaD0Ch49yAS9+T6w52uLQ0bxxv
Z0LiaasiKvVE8TpS2WJyPw0YKGvTNBqVxRdYG+9/Ku04o7pXxC/IlEtGost45369
uo484u9HWl7Pdt0UQWmzfDAOChzoyiYKsWJEaM+LcD/C1b3VFHEpUW0mTuSIi4G+
90Z6BhLvA1evTntmqPXohek7yB82YwIVQpk2L16ePiGeO04emZ/dJ4QEzYBOj4ik
eFP7A+AcwGAU5fU+VQ2L8Jh3kE8uAy/FGec8KY/JIMxhqjRBvRGaOYvAvdC+lW7j
TMeaXJuIJd4bK+jfZXeQ12wLG3BrQEMdtFtebGFPwEH1oLGpce3JYhFEJEos4hTS
gFxaqTJ+G1o+aAGTiqcAut0ogy+RRuuQSkKN4O8lS5p9v8IFm4X56ztFUO1qW9Ak
SemsaKymLanOOAYdmaXaeNQZlYHhKXNOfyIkYYDwFL/AO8mFtGxFFg/ThF9KGqXI
5SRlT7f0WkQgT6zUYluu6sA0JULEsb7A8/6qlVipCyI75UZDMJvROybZesRXiikD
HjEsnHXCboclmDTa2qH6vGqqoHdaItZDu34E7401vVMyqPLT6CQKZv5yo3RhkJvu
HlxO/qpSJukLKincRr2a2JWV/dj9Z6uS+X2XiqYSdD0ryBDZZY3Yvu5jHmmlqeKL
MlYILenJsnqC/leYREoi6zB+T9P5LQgy/qExADjE0xFVO8BOd232yt05nYf3pVWA
KHtVEyuyMidZ8TR/vN9BbT0CFqLonNS1ITpuvhDiYrdgs4uqtCbMj9cFQ6tQVrvw
+jQ1h/C9x+0ovP7Ua0n8LjQM+o8VpiWFhmhjKWfwdsAD5UwHfWLZJErwBEWqOhsg
oHMYSijrgFCul5DukoSCvqA/B2GQyQhoxwSTVaOiUvCPNQIRN01XS0T3KshkcNvM
7O/1AErW7LfZIbtRumqD/dUnETBVRD2GlI8YKbKdlZidcGnX0co+UTMkKwzEekto
XtZ7tMz0pIqmzrpGxgJl9n5wssw0FL0TCIomG7PxHAPaGC4DtwNmdRgoxwWTKJIS
R8U7Edo+Tsj1ft/3UxXK/EDGAqtmXGMtfeVCKTv2bCCDF3YxdQB8JdcSrmxXDPA/
ehlcYSR+yg951nWzSsq8AUhMZBXz+ldhZ20fEjes53F3GYZuwJULLSLNfFNToj84
ZjMieioG7Oa+FnbBFTkV8N3tIlv8Lbn3qAMWZAWAnxMc52boLvUFg0MtUJWY3UI5
nWPDVKx2kUaL1s5G3KgsqVTnDVZsYya/s8FJKrYSzkGP8Wa54tILdj9VBYJ/Cd++
HCsOBFS02IHe00Rxw1yyr8AYblBaX+fBYqF9RuYlJUv+ns4ALb/ufkRXQKldAvuH
HMjC9GvH15+nGLbV3P6BDs8fCtCPkFWz/pJE6JiKYn9r6zheDqaYtzcc6Fi9pXG2
yB9NLPBVRRIj4wBl0RyKxniYW4EFf+rE6jv5X0P3bW/97W9P9trFCHqUZUGvCNCe
TUkRs4T+sPaqWtk1C0trx+xEKNtl2baP63V+EtptUWBxpsoAHJgFVqEKQE/vezGq
xF9WOyE9AvqayUgMqaJPKcz93pRHo4v7ExQJooeQTNQ/fcnhZydE7k4+DwFZjk9G
iMF8PbXEWjsBC54K/dVW2G+JwzgJoRKe88UEyX9TbsnLb+wMDwLCJ5SbqQkOdMQr
FKxZWjUoGk0twIZy2GHaEDU90wNIbM8fVawd74YCBqP2w2K2/G2VZ7eY413vh9Eg
8314f3rZfNdApY0QbqbtzH+VnxLs4YAXaCEOcGNh1pAXUUnNtBzfV5yiYKldlHZI
FkGIEMQKkGN8EDmkd8ngEr+OhsGoF4FclyBLVM4vvYcpxbD4XfQ5zmaz7fvxPX9z
qTNykRSUPZ0vwwbgzhOLvKO/pFrXOBhHA1zdGGXxf1ugb6IhVwTYu5Y95kkh83fr
HTZwk7ceuwtiBZZLng2pK2eFiRstgYSYCtxogvDqkLOOLTTWqCAELLu1Vyhh89Q6
e/KtIKX60EF3GjE49HX/out1xrcxzvKjg3YlP3yr55zyMRV7d1z/UgmsGBeS0S6+
voNggC/10q1889Tat430TkvxkUGCUffb4Bxl1hM9pkEYwFMu0ZOgJVT5ZNyZZbbQ
nwubvJ10x+0itodecpk7Cjgwi6NKPfxCgjBXEowEz0jQ/0bHikz69LZuXsv6BiKg
2KKkNBWgmcjtwfKOAXiGr3FpKhtIC3CyOnfMGnaqr+HuJYa6Awd6xJxENTrSizCO
JNCjrPQDtRthni8nMSGkZWae3Xaxn2UJ1ZOnHuhzGRrRC0ReyXUIZvfvcUCmErc5
0Uf748UR21e6i0bUXsEz6fyhn878SjswUIQnvrEkdz38WaYAi2XkChvdGZvy5DGk
4FYSu+cImLK19Ngn1qYZ8L1ld4nzcQUcUIg36w4NZlPktFTtbzfdUeARBSYUMhLO
TJq/x/c+RZg9SeX8LEbnVtDEnv3ImJ8CxDT4BAPDMSuc8WbNZZFdD6cyKtm1W0+V
/mO7fp6vf2vPi+Er550r+JFMGI8OrX3f4AMYAghC1TT8hI65KzsQwRt4djxo1Q4d
KrtzXjcF9xapCeI2YUAqk//+0U5WEAmmnECs9uMqy0zecGPoak8Ci3RnDn4Ykgpb
tDiOC0hXCb1AWxN+ODJWAmhIVeE1MN9fVzsGN/exc5pLjm1K5yU+HX7vcUdK5djA
rTVqHi7Tr7Bs3AwtBZWqBeGp55XAgDjCoDbzlfj0MNViBEzcHTKUi5q+twMkiCBm
GdvJwpniQHP4mjDwikhlQhXNFcg95v7iN3pxNceyt6cTe4P4l9qHfQ/vGYuK3feM
QylW77p4D2MggizPpilR6K5rbMvyTvV9lT4GV+bGiUGf4AuMk/jhb1kekgMyxPTx
VFDoYsQfTq3nNYMAxX2V82aiso7aKS1nrMpYkIG35lbQ9Pde45YgikrjB+x8xMMD
VD3YcTCsA5HuJwdTWQEGCqh9dqpfpoFB4eGE9zBhin60gNv0HzlmEHmqErfpa2Kd
2z2+pziYuXaAHJgW1Bgf4tWNt68amMBZzqo2d6xlJ62wPFPxTJVJsCGNnJrW+0zw
xxzx9669Z7oWTYs4nuahsWJGREh9wW0t44nhEiSszXAGtxYcICCrpCxcr99VhpwB
oLKqYAcOU2JDU1G3lqTjS+mNqT84iHBZWP1+Y+eOyh97QJtwsr4KDhltzkrkOQ4Z
PSZ42cdW/i6pP+WwUtSQKgbhSOTmd69ed7QNs56GbII9OAtoxhXr6t4T8qcgcoNn
E1ecSrlsDm3bB5gtNQyccLNRdERpeIXVo2G7oAii4qkE+rgJQvbhTL9NAlcQJ49H
UjnNkYdEwe05wpvj7YbJBtAKw94YaCTwb6yrF7P1MP4OR0GK1DL7yIus3aKg+zju
nnzg6LJcqaVVsST2A7B0SfzD+UFgA1lc5Dgr7W4j74GNE6uQMlOBEDkn8xTFDC06
5i99mnRsMiDWhDTSR0D/DGaGN6ynjKTgto91mn9Ta9Ks+deK6CZfExVAPA1aE7TI
PahO3P+GwUkc9023OOeclO1OjII3d9WHJ26QNimJ6Oav/uOTNA9krMftMa+6hPRr
RcSkxCEp6gcZgjBJkuFQ+y1q4rkis5neYjDwrMLIjZm4S9UN1h9+9ojVZ+ewD2+g
+fX0FYHSLz4eCn67nGxiuByWr2UjW4fu88rTkfAQUetgIuKWtZx+9Ov66qidluuC
d/wRyeKPnbhfKfC7txjyDvAFceEI0Iwse/8blhvilKLnB5eHQxw7usxLBzS22WLC
hJ2eXBBAc239P0gtmiNqiWcVuTXc3CkPo12mvqHK26PdwKyFIb2mhYiW40XEDdUk
FHxHnnyO177xK00g2/awsViw1TtsJPiA6uwTiJHPKsCBTDsvH3TrY0rPe+VNhBZX
ksxfYRjpopjnrbl6sy2y4VJ1qou8fn4fyGHvstFRWuBXvfgao8kW+btw2d1QLtEV
W+XzXPgwmG2puwqtGKAAEFMqvZvcULaqzaIKl+XLQXNHwwGzaUMRwGtQCXqnRF5V
pQ1XmZ7+iVsDur6QLmRcg2O3bmrNHKS+5MWWpH8rXf9TPlhoU99VurfebGnFjWdK
ia6ppTEnMsbYZJuQ0ZXpdKVTrV7W0TY14LqsPoqgFJlEfo5IDXzV2OJFBORMmQD6
piCqck/bN4Ldka3gYjZe8aE7L+YSOySLOLqefa5KdqIgPgADlFlGJucxKkzNqc12
NqhbXLA/oCXDygSAoVi/MUVJpVv16tERktt44GF5ajVhdc/xe/N8kulShdY8yvZp
Puy/HsGAyZ0ocTXpmEhZNhC3JG2iQ8nuE8P8Hot/f0s1EeezNu+bkDNZUhsnA8AJ
ruYXC0xoCN6DmeFE9sxKQBEK0y4L5FSPKl5dY0dFH+mLsH2A+Md+pDCprBVJj3pL
PXsJzD+9xkLW/4VM6/afkZSPEQ7Kmi/goOKXvvCVP/Di4SyD/YsF/yDelW9rV5Fq
meIomi8VtulBFsB5V7ubNTt2abrLJr4H8zU6cGfC2gfgFKbLUhGxCZIR6rs0Plu4
lEaGIUby4FTF8aECQgX3w2egvl+h2VUAKhxasC6Agxm+3MAeHiS9J+XEGkoYkNnx
/5FRrN7s8jtG5xVMwskei9oe6lgCr+tEplxkF5+R5VrSm1zwioFnI2tV+cvXfRxd
elzZYCl9WRdAlYMMJfTdBjrbwXnJJTd2sDyVoF0Nou3nk0V+3C8a71V8pu6w4ugU
DNxiqt6LecqrrdEiDYZCaTdxfqhwQXEP/zo/NdKI0/xriLG1Tt9XRqDKVFy7Jinf
jkKLw963nacmqwf5fCP/CqM1fck04n6Ja1ztxYGna2Pk4kH9UhXhlHawSBIltSg0
za3GnK2Z1gPf+IB6a3wZdT4nO8+i72pr6+UViVZAA3nKAcXojikOYXS8e9Ia+jL/
fFMNi3C5oO4mWa5whotonu9Z6Fc+lxWc5BW6vQ5a7kLYnKQx4ku/NuuQ6ontvOrl
JCPcqYTW/gfmIoZe1pKwBcfZVounRWv1L942kE8ip+Tshfmx60KC0PLDUXGyvuBa
MVNj/VilLdeI6/nUqbbAkyo8T0BrcUalLnJdQ7pdilU76djE1aC1cOzdr+zviNvf
U7Q/PeGhum8clYJ8wvVY+33R2z9b3YUlPzw85i+pqYLEugXZp67dbEXnUnGs/kiX
8o/uiZUn36JdGRzXgcLshlNuLkesxd41A5x6gg/xYt+y9dYlnqLhLTwDmQFyXEJY
jyLCfwbO4mqcEevQP0PmHApK1iyXHd30pNo5zJt1hSTt5a+fW6hT/95d8YxlMXi/
CMqAO6KlJDMeM3KW9sRaAwag1VkR8cUJH1f73THw0xFeB+RMWnlpO4kDcIsseaqt
VpW42KqXUu8q0WtHofcuu+xAOWUAFuWX8Klw/+tHbqe3URISQbNRPKoIK2RusagR
JwCOzlKkOXlVKW7J5qRAV3o11RM4bB+itwHsJcLNobqfGRcruBhPN8LM/KJ58eN8
kpLL/YqVlHY3BiZgzUfB9RmC2htmatrsyV8iBGc1BMA/7svADHA3HCF6hnrlF/ir
83gURChA3uBcLHFLuOe8Rz0xmJ6dw4jzi2lHNku9C/k7ZA8fxykx1ozKRFMX2F4R
UHZQYBFS0O7lPXyeH5xMWTXgZW7ngic5SI9b8+jzkf4GX10E6zBkYOMDAQx6KnMn
Dc5IvkJe5YIOKgacn7I+07stCW2tnR90QlQHuZ1J2sZK2LHgdhlsZqWcrv8V6lpI
FqtgpayppbFqfDn3VCwSFg01G+pfgGHLEnaCQ7XEuIXduMxcVEgpz0z1JSxulGxs
pMEfP9IvbIEQxycLtnzqMF/FsOaIYymNvbiDqUAaiVMmA+L/st7zA7USIeNrKbGz
7hBadfMyhGG2i/K7Dj5+r4PXdiLbiPJ7BpHNl+ursyApw/MswkMmSli1nnolXuiK
Enn9BDdiygfs3A4vGkS6y1yj/LBBrC7qoKrOQPwZtc4nNvlGo0jHkfacYrqaeiq0
UHislFgB4qHvuzia7lsQvvlZFajtB/7hweCAoz655cE//E6B64GAv8kOvvC2Zypm
ENnWLVwr/RUgz5CC/oC0qhgDLa3fcACT4y46a91lqZGRqXTCHZAgjR/VOOgNo2TB
44fb3HbWNdxCBbqcR1Ki6QIdxNzACnWZqymfMrXglhsf6WH9xjRmcJoGDl4/+8VW
fMQEiCKwKuXlP6OJEQWYbQ7G4vi+TydFc11Q46/LYGAoGJc14NyKpg62NvWRdqcB
9rmWCZEo85RinkxvIh+BLVgd2YGB0tiSR9w8IpTosdq5OBBmaBtM8S9UQWAbbJhD
hOi4XwRvrP98y56J2Ql6EsVHofMYKGBY8MFG2Tgo4X/d/FjUij+/usIGOHQS6SS9
9h/03XELSfF+fbcGRDqEQ/iE4vJPfF2rFTAh/A/6ohNrNoqeaZE31mZZytlx99L4
jcVeEVMVY2m3P+vygnNy0EpkDUT68Jl9N4FHbBJiL/15s1XEm0od0GL9CCDsjKcm
QPH6e+vRRaTd+4ewAQBOs474T8AHKMU1Ljv1V2FxvwTEXxPF93LWtoQoRKIURcfP
iURqikw/L+yWaX/e3WcwL6tO4x2qdvGhw28ZOJL3XaWHrXQqZPtj1Ls3a2xuSGyu
bvCQNaCALEG/ylFtPA2jnUshnavBPjn+g+gXxwL5z8bva6qryarqRTKNXWxgC/nv
SSS1TStzymx+07tgE5ydryS6OQUEjsG94dCQH+hoLTYafGUm82aT1zSjUs4oabJ5
SEIE/mEu+EOkiCl013YzS1Lo9ftpWjIVYoc2bdBQisGdhfWRcC99SfYQWfJQs41c
9odQR6rizbYW2uIgrfe2JtOUs31y+zX0QCD+56YG0N3ASvfipPKO0otn3qXHMa1c
0w5hl/3aNSP1Z3qqXgbs4hRN8ZQOIRgsEtA5xp8Wbbov5Vh1qMagqt/4jP/2gGK5
Cr3W6byr6X/L6Vg1do6DIASvBDhOoAg0qM9LCt3EbXRuUP0/UTH/gFBdmX/+W+6o
mc/+/vd4mZR47h8vSKQNv1fUon0lQIbVKkubLE+WQdoJFzMN8MGC46Gl6GNZnb72
lAQH/XxMm67fS8Cb0CCjxZr+8PHRnk2wEousNrOcLeGZ8zTFq/DwB7AlbpUrKpHp
rnLDTd23SPmKXP3Nz/fq7plToS90segkzttoTLN575+EQi9XbUBhZfKFipBMNiAq
1uZcyH/Ekg/qZn0iHf4kMAlymTRsJGTzrDchiPWDfF4Rmc42HP+mXJ30v677+YKu
lE6FYruSxFQ95o+t5rb8qu+Q5qt3wVNEnRaaG27uokzgLMwoqhHj98wKAvOIi1a2
/pJWRiwr2cEBsDDsG9Ys7K73VEBqyvCXQUOlMzxOCyd8DWLW2HTmMJRn3avHUWy6
u6eVq6JYfsKbIKitprXHaD12MuBhEtssQcLvLZ53tK5rDb/TTXvMcRkmxZlyajtf
zY9FZVApdq0R/bdVOSpSS8PwF41rTdQYn2O6PgvTflx9x0PDowKcavl67KiqiH+W
hFR8xI2RRQXt/wxUsgEeTq2t+DRsn9+MjBokkZpEK0Wqnf7U4WHtpbciMFB+J8/l
z4I+dp/6ymFycvvRArKbQgM30B3lTpM5GauhyLha0nZmmM9Zt0oam8SOdKXB1U3K
qT6oBm0g6mXW5W4mrngRezz1hkKGVARaKS0KcwJDCujuUNoGm4VWlBzx69PrmNtk
G5J/wLjdD/zNlEX+amuZ/dsGoAYmvdS4uZdU9k80xwyFGa7O908K01vgybhRoBoR
9lHa3Rtr7AzD5941S8l3QlgNulYsgj2AuoGXgZzOXhkGcH6M2clWYqRiMtm5AOcJ
zwhwhxRv4o9SFHwgoHREXw7MqdCRM4ATMLNcFRI1UA2y7RUMLcqrDhbndMlC1uyc
sMZIxxz4Pw1F+oN1Ig3Sb8q/qg2geJCJxhv4GMS1UL+jri28f8ajJw4SygfftX6O
DHzrE5dHeOB2HokP4JQ0SR4BdXvysgWu8/G9ROSWQCsHdLqZkkbvdctkiZlXFJTC
L4pOU+SnyR+qckyZg2YYXaOpQtI7vbwd2TOD90WeuspJXEmS28X9ecoj3hrjV1YC
AQXOsSIOWvGxf3ZSdknpUDyU2YPgscFTlOKSM4PuB3+z+cRjQgszfkLyYSeU8+nl
pUmEig/NiZvfgP53x7TDwiJPk1ml7WZK4OgckUwsPRvnImuqRi3kSsunqeyRPYny
c5fThN/EK9hlxYELgWUR7+YhTRXYC698unzs06tAa1jPFg0dA0zQdza+OX3gTo2Z
hvGxUJZJmj3Y0PDsmpPu4V/O9dJbaYIqNl/A6UX0/1PmrAJLWsoRiUJ/GX7RH4OF
k/Wh53Me+uDTy3sLTEfci7A8ytyBko3bJFSWbUrfB4Qxp4Jmur7N2FIacdjiDVmR
mNd3x+710vgwpMhDJVlTJNjdZgppRr3nEX6/ZCkB6qj4oZTvPUc3NlFJvLZ15+Yo
WBTclPay0kqOhx2Z8chqIgBm5KIh9qMAU2wdRPoIwJ0e5bTF6gCbU7hvLwxLIYOm
UqBXdWl4755HDJow/9uMsRUVIsVQHLohduLpCM9RG0lDuZK8sKgmYFFUij062KWK
8vFQNA4kNnD+8H5myxmSshEmQoLRA7ZQGX05syYUPtf3pQOujY7c2sbRzA0s1t6w
jl6ew3RR/6A9cZ5uagsoYYn22uunThWu+R2hkTzCgLhJCGMjq/U3mGXyyGVgu7ft
h5BB1b6n7jazv4JHscOEDpomSb2whoB4Z3owQRWYnoFy0Lww3E6phKsso4QRDZXe
gQgFERH/Xqi5LRHuVRo6XHyNIEqVC6Lg1MOMKoIbIEMudHRm8wLPsbFajuyDa5xP
sByjPO2vFLfEvkl+oJNluVufCB8+7scK+8wlWnJzaY2O4VRnR+rjYjXnDMQqRQPU
awKv2Ft98uumzkRu7K07mJzOFc2FCbDkDRZW1KZILiDMSDjXGZOk1tXdCemW2F/h
yFwVGzfYos/CoDk3tJ/eVvWu6Pk23dNydRZ4Bxdagdy8LR9fbokIa4IA8qGfeYZH
06a0YFSUlp+y1aU9wSRJ23QyGoX1kRMr0Zdwa3ASC3o1SKO0dEenYO10sOuxnJo/
62fdogHrRhxV2IvGHizZgZ3nRg3+P9MLGSE+fK5wCSjRZOjDKqpbfPpCWcOAREmU
lutGjXGvYaXWP8SRD69RtZjFJttmSiwZ5VeY6L+qXeKQ8wZX6gJ4MFn/yGCiCD0j
adkaYEp1TAGHf7QP3yagIPOQySsw3jTD+H8mrY0RBDTXMcvo76Uz7jFyn3LOserj
w48nN4HNxBLLfsBeSJ853nwuwCvUdZ/VOHbWU6ic2amC+/UbC1tpX1jcE0IHa/bl
i1HAD4OkjTk+yKsCYqT5fBtPG44ar2HHW6QPh/VJU5OUQ6IuHd1TXiv14qh2KX6l
AEFxv7G+yfYa0WFIhdxfj8QiMYOTc8aM/fcoZjJbXmg//MmumtIB91eu27YfEMMr
BKMLWRXoB+2r1AY+sSa2bg==
`protect END_PROTECTED
