`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KMm/P3cTvTGI+OLa7C2REDaEQC4HQ3T4SZcE+iKDLIo61O2z8X/y4XMDaybJtuH
2uE3xusjY7ulwvoELQl4eQR8AcyYT/ojKFsFp3Du1IUhVSSppEZID7puNO+ndS/H
k5mi74Teq/w8yH9AWqi6dNQA50SPWI9cUQBAYhrOujCSbq0fN7+xCmai5OmU1puf
kk7H1mdlLfBoJ2E0QWfBLN4arpmssMZ42UetzHnK7IFhiBt3Wej2JOztID/ayXrs
pUlLeOOfVsmrDD4Ixsu24l051CM6rOijhk/8ucuwlKzZaLvptJKcKDA9RxFZFv1g
dKdEbMz3Pe7p47KLQM0TxeZKIVMGL+3lqnFaSkUCkaw11wX5vu1k4+FojqAlHHdK
ZIGqqyfajzeGdbenyj1L3pZj9pkfdVPH7xCGvXQpmU96lvccW+VdCjWu/hx7m76m
bz3Kcay3oYC763/xcwVd/w==
`protect END_PROTECTED
