`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrDYnMqEPC+WH5N4mZ6Cew8XgQi60zhv9ogE45juedEtOqITP3/a2Eita+8MGuxs
KwH3cgewtsRBO1+KqTAbrNucPsit+HqqPslmt5jAcD4zQ+0c+zg6LNgVZC0Qr69K
MKQVQCked2gGCVReJl9mILDIj1NIXNuVlvfWl1v7jbC+W1+b83yz+jvRGp2xCAis
SXh0B/mn57eaEj73z9rXFwRXJlh+PWd//SdQlp4N6+NoyzMmqTwC64YRucwM44uH
ZFBrfU1kfVM4eLJ6wOVbuDucgWvPJG2I+ie9T6tGiQxcfNCunchxTjOaa9RXO8uo
Sw23OUn7wxrLmReB7RFkW6JIzOInhXdAO4nwfQgqz34tOIJMYXm7Mp5oBS8ZyI49
Yno/obh8LB1lskoqieuDRM6kY2fNKPh1gJUUdrUSCPLTU+ZwR0fD2O5Ixy1JSNWO
AbNvRh4XfLVLOKjrO2z0Y7G/gsor6gaJk7esOZDA40NvjGxpIrFI5cWBn1a5LybD
L5xHdo96/aLxmB2Kd468sBp59ipu+Bfp5yQhLd/oixAr6MzJHha6OoBPJu6Bvy3+
ZlF6RihjqIIaFbdEBVtkVw2gBDRhVYYcgjNiLQM7qiPmvRdTQ6ZbZRSy0ltLq3RV
PE5Ayf3KW5PKxSHIYC1IdhKuBzH/jOcCiuHtUCTIORU6mK/BpnGmPK/+dFghd5Wn
syQQvoMBWQYthp2cha+9lv+nql3af4aFXzAgvKOMjgkaep123/oyBcLlKM3XmkzU
LYB4UZXWL9U+NxV5DIZi7XpdIfcP05QTfcqUA6ql4dAbOhuyf4CFDoZC7z+2i1WO
`protect END_PROTECTED
