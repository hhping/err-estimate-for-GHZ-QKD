`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X53MlwC7YShEovBDLEU+K50CycyXLqg0lNfJb7pqY0d4wSvHsTfvvmBXX3t8XPXv
4ev/5BD+zEF02qKyBMtDDpz51sVZOKmC7u6LIuyRyQlMHMfcVrYpip/XlfYTlJbv
3TXyMQ831Il1mMGxInTfGKutHfQ7KxVe5fpksEnaH/4kXA1ByX5xLeZGsvpf86yF
C9OAMGxfdSdM9+G3rAi7mhHVi8wGH7F9bEjlFQret/5oHX8yxHwg/F2Rub8WiSD+
AjOQBOzigRbjLY7zCDz+JPWPA6wqOfnKnQErghidUgw5madNmaO+5E3oy8VtSv5y
5jOKtRx7UYV9NZlAk14D1h7pzzl28kO/bItk+Qf0laUr/j7x58vvLqo+9Zbn8KID
zgvU3FoZEOTapic2vFtD5TVCeITJkGhDkHbSw9vNJVL6qHmxQg/2YyZyjeTEIKzm
sT9hoRFLJDx81733YUBTSQLUZRi+JBSnGqe4vrhVdhdI7fdmt7jOIPiBAhuhGgl6
947HEPP1BrfXQtHM027Cc8bCLNTCfi+GfxOvHbjYn3cWLcyx7cp4XvaQr9afAF7i
KyQRdKTV2J9bGGlgAs+6906mwyfU2WkvyMUK5zjwphUGA7p2ex2H4rekevPRfcBB
1CbIRPw4Dz7SQUMSmUwOrQFnNki2WAx7wxcISYn3I+Pne6TrXVdNopT1QRvzG9NW
JhYCCZtrCraeopCfRm0A245P6hUz5M+kLh9H5LC+0xsVPJmkV0hA6HkN73Nb/VVt
iV3kG7BDWMXm2WgqciYz2FQvolcn6w/srxdFN7UedV2kf75HZWcoD3tBi9FOQ0t6
Urtp1Oy2JwnxR5YE4JARc++LLbsaLj1gFj2r78PjBqe9FxWRtFxvH4vjePoAoHUc
gd4o2mngbUq8L93EEpNwVVtlxAiLC2A66EdIpl1uEO51nch0abknK2FuTfELVCNM
hXMjWXkIQvett/YfLoJeb6OTFoUU8jBMCGlu59Qz55mvlocWBnEAOEflBTOormdE
YoJ3MXtVPR7/kx4bsC2qQG5a7E0OK/yiAgYR0Ug+7sPPrtq8RjhQBP0Tm2/JZbPQ
LFwT1goXcGB+va4PC+XlqhM0kXTF3ssf5xEYdFgKNVKUf+3iORSlxyHmQ51JSCT/
EkOm5Eh/2yJoXQgUYR7Wd4VOthIHcizK43fMxrER6CBYkeLsMSh4DtkyzOdQPLqe
aUcfWJSJ+m2SpGty0JwKjqk8I4PUvWFkP/eF2wiuGZUrZzuqWp74YoT8mrfngrLT
ftF2iEeRINjTUZJ6WEVcDaPyLQHwJE9kPzDw9ja/E2LjKaH4l+/qwN/Kp1B02bJ8
ewPD6KXvBYiIhDZqj+yPoExFDESo0i9QX4BILjP+AJxSd7HnGDN5xXiZbsXYNS5s
ZvGSwL1qRsZhSnryK8Eoi6kIk5Rwq1p7mBl4zPtg51QZim+qx/4Yjb+CgsqB6CJv
8kXPJgaD6Xh5V7qMPaXhDVwAgB1a47sb60lKHGtwrWo42tXlfLFa/QBWvUVkjmWr
fV8IM5v8zr4Bt8fPFApj6PNoXV/nLgzx+UYsYhNS5Jw=
`protect END_PROTECTED
