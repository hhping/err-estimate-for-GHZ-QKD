`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Brt0C2goAL8pEZ439VdkVNWbRIJhZfajd3zi9igP3MCu6wRJGEuhsi8XbCEubVn7
oYCsSwX560LoU0wfhq083OLytqniJC5MgWuNDj8a8lBZ+zEUk7Jqmo26b+wKt2Wx
00j5Wl1FQCk6IxI6C5bdXqZAmH5mYfm+xehOgwl1YRSrbZgnlk58cIoiFg8jBVWj
5l3ZxClElt8GSg6BDLQYI8nAlz+CHo8f+XrTX8kqxjBlX1t7T9UdNbVXHwmCSteV
h0rpxJLGhkVrXQGUxEt42qbrHxNu1mN62EqkhuywnLHjgZvpTh24D+upSP/vAWcz
uiKUIvnbMofl9oP+tyS0QychtR5Qe7POrQnvODPelftv8kS8oNQsqDhUcPOs/Wkr
BzK0YSYIyEEWg3tGCPx3whj8CD2dnRV45q/EXH2sLvXza0Bv3FpsQnyvNGTHwHzh
oPmyL1XQzewvPRrfByW4E5RAKnTTELbdgBffJHFdJwTAoEMVi2Zf7Abhij/6nVqK
RVYvsdg9CfMpSc1oPKNGgOBWmxP0JyosBkPfEmOWl67Jgh6t0euWgtnua9P+dO1c
MsNi+/DIe2+0u4aUad7VIiX7c4hoaiRcB+J9MHil6boRVFWXNNQodnrI6HMSpEo0
`protect END_PROTECTED
