`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+aB+EA/r00oEC7kksvtX/DvIMlvqrWSwGpO6OsDipqAYO0Ee9/X1pPOuMqNTEtb
nwvoXQaW9LFjNpksQLTx9k0RRC+HqjnhE0YfuK2tL14Ll+Z7W16mCnEXZXaj9Fsr
gjsMgC3Xu2/GDEYjkjRvOHOv2yymQVGyz9iCjDmoMzZFPXvvbBOdeB5jcD2UW/XW
uI2M1Z8ELm7Gw1F2cLgbmM9VRc/EpyYLF4j1qb+gAbpjYaHvG+t4NpSBL4EUUCaj
tG4xdH8Ckqz4O23mC/LlRN7aUDMWk1bjOKNNiC+jnllAOwP0z1ydFG/NjRw4eJQe
HIWomQvlPgl8xTkruzV98EvZyXVl8jIRaJu4Ij5CHufgcCSYCI0v7IloEYa39tO8
`protect END_PROTECTED
