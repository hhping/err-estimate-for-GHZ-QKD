`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQcYmaVld0Gbn289l/hDWZAim4vewPj1SyuQfesAbLAHXbwvW9NzWPr8xl9S4J8a
mQfzrnynla1qtK5a+gQ91+/AEVpRFxDBsmQr+pmLmZGpaSXlwnm+B5z4/5SM1cfV
vew65Q7821o7E8BRS1I1LEKNI/goXgKermmFDjUDhuPyazRiqkJ6DcSOUDV3M6Fj
n1uVUgFAB56d6p532AF2drM5PlbhaYjPrsXLDn3ph6m4eb5NW0R37M6P7GzFLoJL
sgxepKUzs6pJtgjE1amxYOWRuA8hiXqBXUKZgaRehmLEH9F7oCFM65pERgxHa1/X
2VAe1fJ7gEsQ3cCxCYiadbpOGJ5hlVIF+5H9Jc+W+gbuo/8O/Nar1rbnh59X2Oj9
y5FXbvzABOpmQPKT7n/v8ktQ7apKPA8JvYXvh0+Z99r+pCL0DgwDtlOVg8nLFGyO
K+hrtTrJfWXygSFdoB2v+aj4zzhnLtX4qr7x/KZKS1Z2NkH4eAyelr5kWts0fj+7
gI8Nm0gni4KoTqqRwH2LxVarS3A7aJQaXuI3i2tqrTMDc2zQUQgTl/FMkODuCu3g
HxNVUAnWyAJwqk7TlxsgmJ0F7hI/HUBQxIQyqb2hQI8a6FdZ13z1a9maNxQnc93f
GBiXt2iBwTI4Etx9X6SrxHK8lpYXtJW3K7KUQcyEPNjKcwTa0v8kM1YxDEkupPeb
`protect END_PROTECTED
