`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mPTYMW+FS0OxI4V9Av8vqy3Nkler/N3O/IZxdwrF5tEOKju2LCu0k/dA0fv8gjn
qjw72zjjcoetF2MJecLCFKhkb44mknpwr3GcEKAcMAoRHAwzOP+GLiB7dRSNvVyP
OlyqgfToV0zQiOKzHDxrzMCUEvMAXUN4omCzdZE3d41NeAk2CidyXbroYrbpLxpf
Sy8xjHbGRsRu8ptz7AQe8Dyc1QHQxsYJIzKIfN8dMSSctyy83FvMyGFAwGOU6Jw0
3+ovUSxbJg1bP51dPLfCRoPF6z+g22WShrm54JEnWpaHW7Sbbf0LXCgTQcOVSgDK
KhrA6mHOVAu/iWqvX7y1Ux9rYsd+tb3uBw2us1DAf7w1FkzHSVBSVWEWmDyKhTtZ
34bR1ZqfcTe7HatzYYZt0muNEsPln4tQ56xK8LlnaYv3a97effLEVeAQnMRoBUyS
`protect END_PROTECTED
