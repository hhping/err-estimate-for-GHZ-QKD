`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQ630+wFEzyPRvRBgtR+rXsqo11QbHqe0/QT3toCHdy2Aew5QBZt/f5uB5wmjUpY
PeU+xh0Eu5xf+9aYOF8PrJIQZbitCz/krDHFp+kh+QC25ZpCK3YN6f5gAtDbK6eZ
ostXYxbexxI3a6Z2EPKNyLT6rTyVNPCxYluXeMdGQlWYoUYp498XU14Y2q2X3UZy
EQ+WOF/ilfqEjkFYLtdRvh2F+ZbWFgZpC8BvXubyF5MDzG4NSwAXpmJhq2jwgSJz
KBFAbi2+J5W07hnQosGGL0KFxXwUniT+Tv8B7G5n3cHdKFUw+wndcfFSv2M5Q0EL
o8TqQwbEAEc4PzUiqMmQAzbUpZYwzYiVXfAG8r+doi8RNITzNnKTFO0IXIeosIgI
C1rMMYyLceWphxnGlrFL4g71jMPXKvDb24AVZ7zITLs6eZ8e8o0T4ukarnyZ7OyU
KNUrlFMw4pORBeKHCRiZdVlYcr63wVzQtx9LCi19G5tyXhDYS21XkUMQ2fc89p2r
LCwkWHAGd8LUL6QKHb49qoRzjfaA0MwvbZv/9CcWhbKsJIi6oaWBSF4xNp1+eSA0
5o7wvsnFJu3E+75OEUf64nqJyayAgzzt0hbN80PW8/bYjVGmhzk2F1LPHinyVO+1
Sj8PSNBBO7yVYqLTwvK5EKHg3/Tkrp+ZYi6coX6+xK6gKnuzsrSGENh3xqfnM/9o
URurj3lvaZ0SaQUIcGr5hYFQQSj93ln/QQKhx/xkajIYSMYyL6apbyMRldmL8/uC
GJLJxEAqVcj8nHtsIPPP6lUEanBk0kwJ9ZndA1pmoI/Jfr9gyh+OuQ6Wgjfyv+GF
dp51sFAr3U3W0+ar7adVSSa5jP4s/Lr7TULam79l8xFzve1sLjJHN+6pPJOhwuyg
c5vOZkGNdrgfJ0lFCKWOBJ33RVaCdezEXDSWxlI5W5hqJuxRIiy3y+OO2t8evnj4
ObSGhRMdQfeGaOB/Zk9taQMKvUQomY7E71iPo8r0nJMJBNNokLhLg9XDMc2T+q2R
ZGWunvVilK3DkJ75cVwN6g9mN6X3VTmVQbbplAc6mxwTJQpdENXTPRaCfCVBNDmV
664566o8LRM/E8kgk+DidcO7zhVPBvGQ5Ujo13P8SP/nmADC8t4y1ubArfrba1Rb
qEPFY+e0XvpONnpZ/8V6y9AmdBb4/R5CRauXddpt+tboHtNhnYzvTqP1psiaOjig
56qb7toxKsbZDLg9TSvwJFs9z9XuSXvV89g5mjC3b9sXLppXwlRT5ZRYIg5ppw/T
wQY2t3A8onKS7EgwgTfkMFPHxE+KaOZdLxriRrkFvpQF1aOzCll9VzO1YUnhA/fp
3NNaK2sQ5+xoCLtv0X+OO+EJ4iElgV0bIxEfQ91zXBHIb9bXGDl5b+Q7YBU3dFaN
IKof9cLq83J0NoyDIC0VdQaQEVkizYdNh20On5UQwhgUpUgEvdimJ4VbnNUlBqa2
DgISx8jU3V5/7g5aa+1FAr7KaAFRz1BropLNleUElXM4zR9urtTu/d/oSbX33eEA
46F9bPEhMj+A+uiXUcK0EOdImxA+VsCO4EmK5PSGi4gTyeWA+t5Y48+7C0SxBmyZ
G29IfCWoPnEiIeltrVEgvlsiHPJQVPN9u8VpyqZ/PQGwhvvdnK4VhGB9a8FE6XCX
JccXMYgRGUhO4uq/1Jn7XquqmTZpewZGitxCa53QvkG+0q4TGKrKLi1MbMGDNHOJ
zbV5yqHAXXwmL6PIUIsGo/LzAgviTmo4oQ2wA6Hv4HGjkKW4ZjK9mR0Z1N6o0W8P
opyrzdKm5quA6Xt34our7DUHQoRnTbSngSxglY2TSvQ6RNVOQXicTQfcDmamI0Aa
4i/EjknS6xXxYDBOhO1yrvbNg39f+decm9m9bF3B3q8LTlFi1IKEECQtu7GcDMUm
0ELnUmGOKnv+3CgDpX36ZqteAu7hLQtLS6hH6uZm9w1WHuEujycc4qYnMzQl1rZF
LdvPq21fj02JUNdu2zlrqyAblOa2ln8XCAjrOp7bNTb8KJ4YnR0V1cIEnm5TFGlf
in6tDnVIZRw1cZlqqRNHShxuXH81xm7jlK83BkrEtUgO2qjoPX/haqofTOagZYIz
FzUO6phKjKE2Ua/LWFSxdyQp1BNlFGFoNLPVl5IX7rAputH3GPg/6Sk/KFR0SaLx
`protect END_PROTECTED
