`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uu+gtsdVw0RLJZxE3isKivP/PjP2VU9bu/aAa0Q+DqbbAT3N/kpzZzGbTPmvi+F
LIqUPfrEeJtr09p8XgmVCHvmDYSMh7PUe7Vo5b8mM1ol0QAFsc9qeFmh164MNfns
kct5W+Mt7qSFHJ4IayveptMT8ej0VMw3m0XG7odmF4yNqtHdbRF1qbZxHCiIqC2w
y0vEJ1RxNjckWBsQR6zQhu4JihdFib0zQts5Q88ItM+nSCrBHhghQNzKttFbHX+o
EYSMfscZON30ZnbfR9m3heRx/33zo7TIaOj8s8o6U64yp5ju8q779fBxaDIPLHT7
C2WdBAWB2M/N77rWbjepIzIIpHxuiIAvIse3t/J2NseFOBFEJRU+V6pUxH0lMftj
esYmgtLJ2vz12qDvRqqP7wvbHNNP8a4NDdMhdgurvmHoadGC9WOobfIRSYYdmUqY
6nItgPPrBpoLdqoHEeP6Htkg9OBqInWp03ItqXwanUDMpBAtUdRPr60UmbwqqBVt
F/7drfQ5byK4O6kQHJPq8pnz7qeiYGOEW70jvacKUQO7K47xPPsD2mXa60bzD0G/
2q6nkWdEwt41LKWFyV0VfbEDQPv6lt9W2lenzqbIj16AJ3H+pqtRAx6p9OYRQMTx
2OUiXeleHOM3gorOHtwYLKi8hd3L5xeO9DQTS58ATxy9XF3j2UogxQTJ9+fD5fn5
FnTa75MR/VO6gzx4kV9x6IRBUTTPWWnHxxNvpsqZMZ7WEWtyihD1Lqiiovp7wkWw
ZdI8zsa/DXgADM5ROoa/IfAQvguLU+2HvS2UajtLm3PyCFdGp1ECf9DMsCGEbQ6u
HFBbua7EAsayWMd3sz49s+4V5jyC36Uv1uGYQ8GtheLYKf7HEi1zeOjH34opF0h1
NDy13EzgfSv6upGfssXwGuQF0dWgnlGUZ/klia6VPPPQNrCIKgTXb0TJrpkKt78s
dib/eu/CdFWvoS7N7ubCWyTQIReqwYhJVIdxol8+a/tIEX4WfxxXE0RxCZIUIWCR
mvItMoad9WhOBSPaeA5nv64ZYv/5WXpwO+LrbKUqNL3W+8AIE+MUuFIuXTOdhquw
lpJhrgQ6/WqsrPHUNLHpfaiJcX0wSRD7D4UsT9gMCUJsOZc+UWFtGBOx1LaTlV46
UHH2kKvxOBhL9/onuiVAXxabzxUVV/mw3Kmp72d5WqFjBEEaIzMkes1MkfVz/2c8
6doKzeDeXT+kUPdiAbToHTPjVhCdwOqpvRcRzqcsWE8b90Rcy1K+QpEKWIIdxxJe
j4GSpk8OhRex1oBBacax3XmfRguoLA9EelUz73IpgRxM0p2A/cRmOV8TeQjd7kLL
+rf3Ge2WDR5hSGazKQ+fPOHtyQHg9HJYwf0eh0EyTF5Yw59jA9zNPMOUrAwq9mb4
NSO4gLBwJjahT5iv6Gt5xVgPyntWfwHa6ISySaDYRuBHQ2/aw9g/pnXNVjchzOcV
mKktvCzoYvnZv3EKckRrsI0PXJ9SGAH+pqbY/aMQRjcRRcEnwKds/+dGUTlT93R6
wdUYIDxR1fgqLTtwBxCPzJRrODJN5hGVsFD+/0yBE3WewHFOrrdYKZLuzChNoLC4
COKv/mNbKZfK4k0w87FFAxVWpbOiaRmJzjqW9EJuGkcIYa0lKEYUjlYEVZkbv4Rz
0tDuBjXGOAu8UBPieDmwba+9f9TZrn4MtWF/hKBlmE1m2RSgZEVXxSkgd4EWhuse
ChcKFeFRrQ/GdGzCyfdYVs4Fn1ZkC0N2b7mg0JQIEB2IhucbwkZHh9ISj+78x+7p
44so4q1TKUDZRdn7CGeM+HQQ1LIjW2h/XyjPRKTy+Nc3LvqhgMR3x+UUQJOZoK06
VLGEPC4z8dwCIePEGXS5qH5/jv8QIZaigJSl1Bpxqhs=
`protect END_PROTECTED
