`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ISVg/5lbs4cVeZdxvSBBbfjzVaLfF7MvLNKlCWnySEgFCWBNNzOZSX8x4lc/sdC
bMPguR1yBP/uFIDs/5c5nfw5XmFpWMhp4uPAJGrjQp0LJJSejiZYPwPXcZ9OD9sV
xfZjM6OOMRI25ezwAm74eMD7Bhu7PFM/TqDK3r4grMtYxyb8xqSPlqfuNEqMydRd
4f3QDHhODQ1t0UF0fyqcdmapN7KI0W4aaaSfBbzS5/V/IFBvSunbDlruH2bVD0If
RxqRatbrLDFh6yscYMxsAM/Xo61MdP+lWa/NePPFCgWiyf8aipqg6WGgiSx7zN/z
YLnOU5ibiq6f7QxFUdsLYFMqUCVU12EHtAQP/J1HqCp0q73iXhT/SBYhHTS+Uwxk
SGYBDOAuHmw+06h/sbUODllbpV7VHjqOCeI5VVIlC2Vd/VC/B9IEhqVnm7bGAvG2
jXALhwnC0BfBt1vZ2XDcA7T6jO0aJMSXaYnOAlq8FSozcQlMD8KHvsQIkX5XSdSb
I8lefXuwRztC2Nhy+yFTbXiGkF5AcRWIH9eBizVCUI2pD/Jz623qt+D8y6X5zDAf
yScL6GLweBt6E/qCVT3wW0DzVV7flsa+UlISB2SB7lPIT3k+l5FZds8DnKXrjw+f
`protect END_PROTECTED
