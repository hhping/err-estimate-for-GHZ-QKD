`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3S/go2x+PIFOs3vKACAFt1S8fMUqY5YqWxnVzGirXqvTWB0BoKGtJnHc/Jgkrl5u
qeK4Fd34cCvieQq6jjJynz0qoBjsrcRrupHZdvAguhsnfUi4ymon+qeipEBTecH/
KuAvciOmOxFH7oDr+eeBnMlpt0N+P1nGqX0F8cih87UoucxQIAltBcNYt9GaYwFm
aQ7xhB16PDFtPa8KgPadM8gHJQeJ1Pe+GnBT20+uJ1LBqgMxpjxVUav4vD4xDTeQ
GGG5YW5O/AuvW/8Tlep4VsHDi0tQ9CcWvsb23kmrSbJ5qeOPoz6aXuZ0WZyYaqfJ
FK1xxXyzJbUNK6iI0Q7thMfKrgMxBW83rke2XtiYW3tOrgi/TBSDspAkQYg19J8T
DLeCB7h0jfSaezNkJHN2viuLoRvN4K30vmTeCGYd+/1PKUs4wjuUs6QY6qI6VveH
O+uiHFeCHgBmhihnP3UfRQ1mc0z8ja4/BzTvQ+mmFnlhxLCZqxEjS8LNB5MjBmmb
adX3XIEZtJS5OVlP5t57jAOn2egzzMX3FyyTw/rtyOw2OVdIZADPBuvDhlmW0MiR
oKNfukEr6SyiOuNhWkWGRaN4GSZe/33bgcheKespKV0wabAJ+/j0yn94XPTDIxKb
WdCDjbKauFHM8IN5wFk6AZxjvvguVoqSvZO25W8KwBlr7ZkT4T+ol6VBs+5gRXCw
ePEvvWl6QtB86GJqSv2iB15eKoVo8dbDoEQMKsv+Y2QLJo2wxDM5c51/9f/eSRnt
JrldhEEax8SLmJZRgWAz2NWk1r5FMDuRIFo+qthLiaFYo/QykRt4vMv7zdDUfdQi
hg6bOY+sr+mOyzcTZl1r1lvSchRVLzRnuUu2VxLa5HufMpHOI6BTrkhEMcZzP+JN
MsIlWbEEbQJEB423hEnLWhu9CR35CD1au5J+DxREDtr855rfnBs6guxeb9viS3cg
fge6Z6zssOqgLjFFr7pXTIu8wvRA+kPGHG1uqIa+0tr1hJLiDP7Cy3BF5jqe6knV
i0ctW3D4kolMdcAdL841cfpmXA22+fEgiFISz5ztC3PUpScDV8x0PLVcPGxGUBT/
`protect END_PROTECTED
