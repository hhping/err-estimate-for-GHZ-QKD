`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
smEG0xXCU2uir2rwLAeveh3cxfmLJTAn6jTrO2HwDhkd3zWXO6QhyA0ZcoIG5QB7
EclqQLpc/SvTvQ8H6YMHEtmmgnvqO/RUURM8UzzsCYuBI4zjGvrRqPxc9v4U7Fx5
UdxP0gtnjq4vEArzv9Ns3FuKcDTg/ZMj/t1Atq8zFAYa9eHXShwPqJ9tEQanvySs
lDPY8NnLckJVJ0GURK7i8aXvz5dkk3e2u0eMKTuEr5+JETwe+TZVF+4TkkvvWssR
aIDfc8umbqoCmdIz0ji4Fnv9zQZXt9ypQ/aKfHSdj3CoDsBDtbbqZq1fhSOGyrLk
d02E8W6L65L3LZq8/odPOe0XPnVYwgMLJqnn7Emt+zZSGGh43+ovxFH+QB4aK8+q
AkGEJ72SWgj55oCj+C0wtLIJw0UVlu4NW/+jITuWnQJDaww1t5048c1nYLk4V4Tj
ITAkNnhqxxaTDDT3RryI/pEGyOtmGLrXSyfx+MEEujao61MXXZ2jGcFsQ1E3Z4gT
a8FfSjZLfJjx3MGXMAg6O2pLbHJv5aYz0KUk9X3n0rqTopUymVqYiHDudGX9qxpq
nzJ+GF+ovaN7tOibarDzAaijjOO9kI5VVO68F1NHUKL/OVmQFtgOS7w8uc5rq4kV
C08U3BQHNi4KDwe2I8tEUGnbNyC3/KSGw46OyNjRfrMScHzqBbTmJzpyn9vWAe4z
br9fJrO16JsNkmFqvz74s5KInSiXVwJb7kYoWv4henGf0E2mgGoHY78JKSTxx5Oj
6GLCdrmk5wl4BbWY+MOIie0A43fN+6pK4u3aoKIUx5VZbSi8/fffnSddSKE1d4Y1
zaBwINGlP5Wxt07PkZGrAA==
`protect END_PROTECTED
