`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3mJ3hINbWVhb4KW+ea2Ln9pInbV/3o1a8iabb0eyzxOecQyLXSJkSVAxKjF4c3f
TVbcbCKwDj7x6orBhw0V+kN8iSPs2wKXEHgV22oJWoKCYAz20GEwzoGfLS7z6j91
la55ddE2FryWDn1hS0K/HX/+f4dz+c7XRjH1+jRQ1B84yytTU3OGzFQ4CmfxrosZ
lF97uoH2wpFZgozXjzygn8BN8KSbg0mw0MQjJvf4WVgmixb/PCs3rpxR3KYdkIDJ
cv+xnZ+Sa8tMbQjgrWnczo0WHcK2v1uWG9snRoc7yO6A8Ai7WsD3mKe5HiDdHRLK
R0hentG7MsmZ+EY559TUL+Ky2o7f6vgAfuEoMgcYMtm3y/5ZydesWEsk2mJTzFVo
9bok8kxRjXUkTdsgW6+B4JAibPwKUIGyLRh+emScBYYbBwzxZM7u/xw/wzx/Rs0e
lfjHjo++V4ThthcdR29Trp0o7dIhbob5NKbQuCszXj52pdECNtuDM9iaiQEBgXnT
db58aSDUONlTCVBFLONTsN2yTOvMKqYBWq43HLyPdlcQDo13Z7ltRMBuPcPamBUq
Afn0qUoixgISQyR3bxMN/cNJbpbAB+DsCPY4EhzEVQscJfRoJgp8g0eYs0W5ESXV
F8vhBvGxP985dkKD3g5k4hUNRFSF7ZIaVxDjpRqxpRqf8OgBCagI1XWvwJEBr7Bi
qjxLe9amvmLt4lDO3hAQXJUX1dsHfvydEOhfbu/1DHHYUVuA5eczF/tLWdOm6MD+
ZvfW8TXEO9gQKW3RBQGx/yRutfXgY0+etibtIvIsL5rNJsUOUesYO/oUnniw15um
a+MA5B/UPetvtwRjnASrmmU23Wls8/xtzYx7fG3z6tPkq2HTYQCOI8nGMKeEUe6M
OvCNNqOY5XPX8xNz3lMPbGdjakZJUTwSSBHq/9yBu/KXJRSmR2EJUM052iueWuus
itRVO101QiEvTN7HOL4B4h5uy880aSVxK89NsORsH1OwubbygWAYp8BztXN+hwoC
d5nwt3X1UF3GRVerr0xNwYarh6CAzviQJQPn54av2prQ460pl+oVlyxfZp/pwVlt
dYXyHUAx8tB95xkIjfmsyTGrgB1/z8DCfalrzAVkLKjDKGjEASx6zhRyHn5eNH82
Zl6pLXORLaJ/JA2LPdBZpOIGmGZvIG1cJi9TQHBBRTuDnjVSzr1ubLaHFDgfsRw2
S8uuBiw6XJI/BvTE89tBRS5TZ8CakuR+tkzQgWa/9IyTkto6DDmUv62lTLSkSn8B
vgtGymVoriDVdFrbfrBwxdn/z+V4HFkz9HTvQREBH49rYYMybedZypGKs4NkEJ/f
1qc0F6uBoRmnRYoeph/EQvjng7X1xKmhgIsnLts7DXHdpQG9sInpI/rT4eC1QTHs
kBiezo59Bk6OrWkfas0XIA5WxT9wcxTAQae3SG7C2V+gEho+g/z4wJgJYsHo4uJY
48PQs9f1XiGaOH5AnUUgCup+8xsfUOYu+k94tk05HZUEVC1+KPOC4pAXAcAnEm8H
YfqPShenb08Sp83rlwxKciUtbLFSWFrGV7tj1mPgWeu1vGpt+1tMWkZlpC8PAorJ
cz2Nf8XM7F4YVCm47f0r19RZuR5Ax3TlKxs09S/ODl+MmrO7mUXO1cUOClU6K8iu
CcJi/BO2+dEidlbAuUUQ9DCKH7fr2dQ/4I57ykCODxLuLoP7CZnkQ00TLo76Xsy6
6rkaFQayumynYSUFl+/T8MnvXBWNwEjzmYnQfxDijYmgQPd8d9DOe8oBvaL6RHwS
WPxR7YbYXww3yjhKnz929XjSXVgUkVHg7LNHyvI+I325vjlsk1R4A0A26sqJW4wp
uCiH2QH8rtK1OoC7z42CSiNoxwbmadRu/T8F0PeNnjPNIEWQW5xjBf3tcLFkafW5
E6OuoPpeh53hSEgmOwwnh+GrZiNTJnTHLa31Yyvq323GRGUe6fx9wLb1lrAHSsBG
TS7mDl2qqyemyFF+hwI+72JYD38g6jY/QXmZRtOpTHJWGeoDGtM5s8c+EHXreJOd
ULm1/cuj9Z3CAxgz52+kOQJtH8vzXcuGysnBHtYEds8gW9HpMGCy3KFV0XF9yE2c
2auTp9LLQvEjJiF12F3N63hgAhUEY08eAsLRnzs/a1uiAFQPOlFSB1e+9pDuq8Yo
S255WJmT7l4CKOO7+hU5pLwqB5Zx4iEbdtzjayommJe95IUM6Nt94u5qjrGYOwx+
+OZlQcjEr1c9Pm7nLHesRDrSKTEH+LemcCUzRqitMxIXBn4ocMWWPVcY35pDgDdp
6+lTbp4euF/gkyVvfNB0s4VjMzRoeyXuXelbED+jW6UGvK9Q2DcEmkvLu4rWAEab
sAH/4PHECO6tvi6WMTPck24a7VeHIPUc5msa1coYB8nPmAFDQ4p9FIiChuCFAdVf
6VwhtRaL3Qvw4VbjlRwG9mW/wlS0wBOOZn7ZeL5bc8nU12YG0hh6I+qfpx3bstW0
I35rl6UIui1T1SkBYI32MAsSom8dL5B0CbDJ6HRWcDtTsuNeaIoasNNIJDlq35lB
rU1UJo+Pm3B15TkmzC12B8/PSgGzYSxaaGSs+Q75SXnFvSsifCmu/HkINto3SJ/q
PTFM6VH3irRheNO6yhNtBuj2f6u2mXJLiADdidV0FPyi1FSAEeke4jP7qdHO7zLK
PZFdftNFV0YB2XtdMliFYN4rTxlYl8mmZ2EC03PBPJp8SgzrRsykC9FexmkTTnr+
4Dm4YDzsDd9Gc0ZYSgY/96kbeN6BNL7YyZo838aRVAhTqJZq+QgFD+9zdSzd6WEj
mEX4IoEaexDW5qdMbw9GKeT9GS5zWBHqyAaLIRvTNk6KpiGfOVf9Mn/AA0hr0pCA
vIF8ujYLZL7emdzuT1d8QS1Pvb9Azp4917iM8l7mSj2JltBFk7x+F4Zhn6hzc2Ai
a1IWSNDhX6A952xbKak9/GxMcJHuhNQekvVfZUhAHBwdQ4obBuLkWlaa5PHrd9sY
1Riv28Ha0w3aQIFPzy6x18jxGlEwmEziOoCFvqyoNnu3ammMAkTBGeoiHZAqSSFy
BS/Eu9DNrY73lKx3Rn24b7TQcOe/BG3wrYFKTLmPHk/NT2Dls4/uueR1A0cigavm
voT2L9PVPHiMZdVyjw/ho8PkoL+IV1mqDgVghejDQb+odmj3j02zmO4/2I2GAa5s
a6nKvOpo7qhFyULDFyfTLF8K0q9/9P1D8DxIO0DOieaaBgMHHukzU3ed0v9HSvar
EQBnEqtrTBUaEQXpQRouYRQ0+7D6y++0MRkGPw69hdGEYuovntyZqYxklch89H4c
K7hS4mRqg3rKheAmvBIgy9rNOlR7SLyzo+ouU74YACkjaY2bnD1pvGyGsXUuRr4i
IPG4Sdq1lDKHdiHYF04GMzX13gqaP6pj0WRpdc+UKd8RLNhKRg5QWTXNl1N/ml5Z
i7ZXKM9WWlu+lCU+yEGMeI28nDe8Nh/oMnGY7TG5oyXdUeTA9KxmmcDnxgf/sxUL
uMnrEVv2DSLidWayDgBRJYviZknecTDpXbx8dUCwLaA5wTwrqWpCZiV6OrqRXGs0
JuDL28qcjs+bFQ7yk7aAr/se0AGpxuwAoivgehdW58tJ/fomzwg8pIpENYPeoa/Y
YJ/QP7kKG0xId93IHqZWV+mGz/tmap97qUu6RUbc7Ye2grobhZgeJkrQlwTTAWB7
4+IDE3YbNR+qn/CE/wkkCMXsvkta1Ky7xcAn20oRLVBBGIkrIDFY39DjEap/U5MC
N4jCyoUNTb39hiJ29J4sWbFXr4mcAaKtmhaOLoKLwjyNnAoFF/a+e72FbRN43ADe
i/GlE2TFEViT26dlNzvttqpF3mwPWao7yB/KO//iyjUQ0P5A2hVNCy8is5FG42Qj
vBhcbtbV8btlCpTPFslbnX1BbkZsp8cc2q8QQg+ovOSwJotyxbGd5a5xDONRa2Zs
hHqhj5ENcl2eKSSfNakS1FLSXgoMuyL4+ds+p1zT5UIm1bfMnBXIxYAuZklynJos
jddks+hnMGh7Kvzga0HEtNsdJ0QUBcGJ/EC9XbaRYOzzKEbtcL5qwX24YtuPnlA5
nhXI6lNNTf/XYO8g9yX2Z90mgEJLVkqFeGmegRM1hhscwf4niH0o5DHXixfHjsPk
sB4zDPgChcCl0PunDOCZJCo/fnROBzUrdlIOiLhOjE5S9EEHRFNxhvsDXXjAcaKV
Byh8oi/LrbYPLwu+OKLZCodAkauWgNQZ6jckCf0A1RfeacLVcx/A6uK9sIefKpTU
uDHvvM/RKn4tXv1MKnJ7R6Bp17/RJdxfkQpe37oy3yY4THgJ4f/rDz1LLdOhEtT1
l5MQcKTgw761nd3+aMBsGRM7i4XOwgxG6914WqUzhN+dRwGxiwHAZIBbpP2Qtvvq
uCo1Nw6VhOyp38xKuHcgfozeHy/++b5FqBIJBS7fHAyOzWw74GhuAQv6nDM2liBy
qTXoFsNEOmFiTCknwUkPd8nFSIjfdvWDsSu6RNSh4MGrRsTHUH9UPaHaRD6qFr24
lv/HCNw3/gZsKoViLwlDeKirVWoGtLWV7jkgyz3ibbKT72tFQ6M4V1Qj3N+u+uxN
8juXy5QH2CwZnz2EJ9qdoYAW2y/DDET3HQqgiSfzAQUDH0m95JuUVDRwan8M/AYX
tMfCEpr7niRRMgCA0EALQBIY1SPmFX71MtU3Usva9JBRTRDmR3oHj9n68XRJSZzB
56x3NiWyeNvMYYsTdzIAWgOJhHDI35s3VsK2xO3rQsqPobYdu78ESJlo5GoNaulh
+eKgxILfqiSFCMJe1VPf+yez4jHZGN8EguWHGDoW/vKvp28QsLlk3ExUl+70J8my
pYHnyYgrjQ6Zjhh/Wru7PRp5+ew1eNCW1QyS15ySFEvOJTTSwx0pU88LqGBC4Gx7
NN0uudNIF1U35IHJFdSkMtIRX/mhHji4MfJYBC5F1BuylPHQ1/4JruLAdlKE0RBI
BF8EtP1cHoAzophI4DKTPkyYoGLTWXLjWFgcqUTAHOD9tuDcNIG+IoKn+nRc5F6A
BaEGQdAWulBZcJh7zw/UiDkMeuuZFbvLVjyjjschiqASSlVC2Krmo8KuxngMuilS
EW1WXYngni4NB0jwiUyLUlLban8BbAil45yGdcESWzxztoPgldcxoiw4SBlU99Fr
M871ry8rJrtfl5yxSflYZ30mOrX1SJskeJW0Dj2JBFBFaz91AdfNa2zLvTiMjpKS
LNgauVfLw4fZ2k115K/lPnm0Lh6AeVESoBavcRHk/+k0Ia+H8kvyeqySSHxil8Lr
6zDuf1nVWkZQ6EYRe3yA8j3PbnAFFoLhqMTk27xe4VnLoJnDViLm+RWuizs6xFJ2
YLQnH5bYwvHQJwVMBxEmmE2FVaMeVFBb4ddh+tftfPP5lDfqlBheuT+f6R5Kg0Fc
LySr7u+weOGzXGeWlB9vhZ4rVltcPzKXZcpBntPFFmjqZWqfG1CGP6DJG7ozfwXr
k7LDgxwuc866G7JLXGyaFexxvFzwfOqm4oZt0S+r+6+dVrUzbFTaNhQC0UdyEI/p
YR5dRyEt5oWkbi0RSCR+W9Nypqb7LOuRE5sqVuCkIyr9PaNy4ZKMolGYRccTwpbd
nbPXvAf0O8FktkKkBbFQMssL09dwZ008xfx97XyeKLhl7AEOSkB2gtBnG7nIHBZY
M7mUFXXmhZMTrcKv308l2EvZkfGuivQILM/BfVX5w0Jo7ljPwCsujOvE73PhWQ//
8SKlBxjc+smk/Pis3cLSd1uMMaRCt9gQvCH8niJfDQWRNh2QdiSOVRmYXmD1pzdn
TxWDK00BsgZH+W7NqLTgXxEjGU4sclbt8RR8oY8WSgJkpdSqwKTNhGQY8zU/LWqC
I6Bog1WumKhQzkth0JrLJLU8OZ5VhW7MxZzxxAqYjH60l1u9yl1fMt4AIf3sNbC1
wWrDVl2wzGojXEiQzGbfQw==
`protect END_PROTECTED
