`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QL2KLPtD+bYSa/zwBJiP7YNeMMjYjX7Nt0/EDXAJ0eNz/JzH+L0kkhppz6fl6gWf
oZhwx37C5zqDgAiiPZSH9MVkVf/kAjPiOu14ypiQN4hqDRk/a+ntKZTzbLuORdOr
zFYIpIN+KKJGEJ9joemlhNs/Ag7tMVb/59UgTWLvVryHNjwNQoCZbjVMQ3k1Gbea
0T+A0Q2F0YivtJcytrRpPl/aWzQZ9h4n4Ua6fmpbfst7sV+KfF7GJek+gVOSNFZa
wxl/D2dngAnN2ASE6Er8Oy4a16gqooAbDdA4ylh6WtI+j1xwIR+NfnwLceqkGvDa
jgZgxLgT1LUf9C583s9avLfrZk+G99xEEGbez5YiAlZbEzdfOMp5yh8XmGsE07Wt
tZDwfUvS+wp/MvyWY2hO27+OWl3nC9rg/snycDESqsjmenz0UXviASjk4bc83iXM
IRzxdfTrpAzCH0syLbCNfZ2ibcA4sDNAHdfR3BZ5pRmuIMmfSk2nEhHzL8e0yZhm
nWYZXeB4xaSP/gtMfV9WEv+1UMhvfLGXlDXKRKGS0h0rh4MjnGXJQ4h8ZusS8+ro
kZJrYZQnIEb3p1cfCq4EyKSiJv8WMMenB3RZdyuJCD8=
`protect END_PROTECTED
