`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKRiYkqH4XWGvBWNDHTX04H/WrOiT2IuF0ZBU3YiVq4W+GPZheDTbBgWXnPuCysK
RiWDopvBZRx6cO4CTXWXHk/7GKW/Wqhso7rUoQXZCKRYKhtLpsRWw8dtR1q5TQt3
z/1ehBcbAvcEjPIseC1kMVqRZ+oS4p4/VUJn0gaW0anOqSofIXGyqz+1wtue3MRA
cpMIzgT0GUjCZWE1FdEYDXpV5IADHP9xlHP4Mz+uKdaM6NbUpCZ8SiMBxwD7Vp9A
I78kWoGFX5oTx8y0nPvqtPqq1r9IfKT0ls8lcB+JYMIhoR2X0BIIkYS+B27Qk6zH
5bPS702EKu+GV5leiCN9Uw4fINHbQIeRgIXy8aXqoyJhTfOhlu8qZNwCgdaG9bi1
S1tp2aWmXFxzsewD1lU/5AAc91OT0Z2o9RUEeiLjA4uyoL+JSL7sgh5vlDuhOpWe
EiCYr2GT15BHMLEUo/z0R6GkpSIRPV7C7SOcQkTGvBzG3pNNvP4N7DvcIJn4UhVn
MJ3p+VcwPGiQJqggG77GfZQixHOxpx/ZyXCoNczuU/bnzpt3lY6K1qo/fzj1G7ZJ
0yAGts0eYw7JuoExX5lvjVr2F7GTMtA9MsC2oDb0XzxyvI6aTo4CIUAoFaxuzqje
SkZtBAm+lBP6VZkuZcjGeY28bn+I4oJMi0fcojX+jDNZmPoJuEEIA6VlCxYZe/bH
2a/svLtsCEhLHbRKbE3iiahFHq/d+k2Lb4WFMTnnpQE4Bq/1IHXkM0FO9RZm8fsB
1uLjojcu7jOPH1975T0yKAz9s9cKmexhdCT4TdHTUAJCw741i2AVKTZrnCYlENYe
pdVBeb9RZ/AEbZD3Q7iDEF1pxCaagrDXgQ4boOSM7OfmYpcYFbGupzZpObrVu2lA
lcdIa3zkHBLYDjCLG6vZKecX2SpMkWdkZPmjdjCqzjimtraWPWihiu4+AfKYSBs+
23Nl46XrBp6I0fR+tdioh7x2y65pI9BXHbWewPIi5cnfRg9EgFnNzuS1g+58pVrF
nntI8X5ny6VD2L7Pq2oTaP0Y2uGCE5XXpWw5TNplQoKhe7vQGYM5R0PNfS7K+vAT
mufDU2wGWf2u0opm1tTI8kVVykomdezwsO9i5MMJNlyXXZcqYWIRtuEa4CMfAAJL
eSu2No/DgoYuVY7LShOCN7HH6Gl6LjH3ts0uNK7hl7rUZx+d/qJIeEJAqZuNet/o
GiJku3bX5zHH6tj89WVrgFXq7lq7WH558hGznpdYCptdR9Yhzk+fX0o8qFpYLEhx
6S8pBQhJj5ySGW3oJ0rRLCWia5NUWQmQYyqr3juhjtrmza2oa3CQRm/qFzahL9uO
Vs55C+9ZUfnu+SXNXzJsB2gKe4XrZca9TAxjEPrqWROPmQ+6aGnaqYkwL/+R99Rh
EYWDfKMFdzF8r0Q9J/OPahh8ph+fzTehqid0kaeoS90nwaGP8gmUvu1R+xmq2Yia
z6Byxga6yGFfbm7kbq7yy3GWIH448lJ/ldDctPfXQ0V4p4sG+Soles1eCL7HW48L
43n2Q/pyP6Wq9eTaq0I6nHqNtUVCphCimB7QSHQFgT6UdF1A/9QQn5Wcl5WVDUyM
fTxhWFC6hJpGSe9gn2YCJqdG2PwqFsu+CcBGt024OqWLf97Z8Jjy13KAXf97vQsc
zCUdgHsIhyfydI2jm1E7cPU+wy7vCnp4a/TQC/rZxSi7d2wn8102aZIlwEdUhg1O
NKa2GnCiQYH+h3PHOE/KTgz+TRC8zGwB/VENeEUqiU+hAaRosZB+QzoCUcgDZ3+/
qtLEIEHRSqFVhB3Jefbn2Ntj19Sqzr38uNQI4ny5tugoRNPbBGoYQQd5C9PvJ4TL
sxpHI3YKrAC5jXqyGQ9lxg+ojJnM0XXFPf4YW0RYpxhsLB+q2n9IAKMaR483uDWT
s67l+ZoPzZjoLU+BR9uBLFbfI0KtWS9z+amDMWa7oUkmtus/y9nkFQePHDIkKvfj
yYhR4YmnjfzkkDDWdJV6WdaoGAhyBK+L+skJDpa0NnQVPIoIPqRQvi0ktNiH2stj
q2Xgsprt0is5nJByJF3/AIWL4mIKHLLzOESksVAOwnZfBXp7KSyQS14lBP0j0JNJ
Otr79EZ3zdn3EZN9P1z06UVW3aTgecFbs/CR50F3TGYifORTRecQTiCoGPzF9hv5
ay8N/ICLzaNgCLE4T+uh5Hd6Oha2JxueYNk4jZISJkQC89lpdlUr5lkgW5ZtJiQ0
aLIwjh1mRMd5qFBCH8P6xdawuD698+g/5SpAMRiISm4GtWHCBu79Txe8XGfe2i1k
ofC+GB4AEcyQO65cmYfoCqmYTw6bq5O3uswBS+HkKwaTevOxaov+Cw9Y6aG1vgfP
qTDik4TmQ/AZRh0Yucuumpv7OkDs1vkCvtdmq55O0UU1wNBPIXS0KCu8mpHB1Elh
QvD41OeNBStLO6M+nJRZkI5G15HMawTiKzCj0JHJUE+PKW5ourE1SzmidUOubNr4
wDAqlj5ys9HVQLx8nhN+DDHV53ndRhEq0HFdbIqbC3v/ujOG7FjjNS0NW2+DyUnA
OBdSztDuICfYhzC2YyNs7BqJlPCza16u6+Jn9YxBIlePExBAW4sjelblt5kLynQ7
vW8hh+6wEAgICdeELoPOHHOhcjcEva9FNyI4QDMRXp08AaRnrEqLiCt6NueKqK+V
kGGGtZs4S8GBFeIamkrB4vHtEnnfgO8Ims2VYtAkGHupRDL1giKWCPMJTbPoqsDm
G9g5Anxh5Wu/F6qLpV1xGoMXWbQgPob0KO+n2elSDXPACCr3dI9KIGNYZKn/Lp+6
x4rPsB2scGyZ17ICWD5hB0TqR4+LpTmbk3qeaS3tbftw/9ERTev6VbhzngM5mS7p
KBPD6hpyClBpR+dKJdTxd8BKGDPaLZYmXpGuEkbZhkCbiwmgZaPk0wEoBWd8H2YT
9u911TnBaNfxXpVVbIT5mouiqlBeWNhYofXMPmRoxNOOkkhdqgHB648a6i3XdmkT
PAh7uBHL6athrFH5FO4vqBcKueWaBoKBHRA8LdDbOj5DLAu2Q1PkjDrEZhu38fnB
3FT5XCAHUi95PyLIUjeS9eXyebolOs5ODW9UGx9kTKyFxCdYy8CVxs5Q62x2rZs5
qpDl45ul6rFCR1cN7vzHpTmo3ivudsWlw7u6YncD20BcOz8JRwad1mIBR5UEgaKA
FwUa8W5/+9hjrcvdxHJMCY2UWcYR30euxjtA7bVfnZRQLObq1lT5cY9v6dYL7qTf
uTUhRVLRYqhlDD4mwi7UBe9/i0x9WR9KbUsY+wTV1u5vmiwtoCLT0Xw+LIhWzBdN
PSi0M7/eyOLC9ZhJktlbTa45vuri09D3O8+XgMOXWaHtdSvbb8S/QvRrIKy+5NaP
6zi5aRtk6cU6J5r1Rt3Gv8UW3hvpiIt9AF2gEwv2jxked77LOXbsZOrGhw8s5GW1
cpPhNOkPdDCztZBkX+ygs8ePa38K6PHHrnHyTfGRXCOvUEitWJhLhZBr4T+XZu5x
ZB02q8j0v1/XgiNR9VU4Uw6DQtZ5+RcBUrr6pBySCOdQu1u9qCmDUiFjfdEciWk/
j0GBD20qsDdxjnBFdd9wDQFFLjXJeVHvZ7gghuIKNw31RuDZpHv9g7UNMwInXXUz
B9mGgv7EiiLtpw7CIXS7SemCKWI5ixcFWS1T59Lqbr8AFnLkAx8RghP+mH0HxbFg
q6nbGrriCT/J1Tly4qUQZC3DqXJlUbS/eOOUzsu1JpwylnTi9/Dcx6zkp4YPvXp5
Kr6XYzBs5qMTpiyMIrbQmxMF0ZtTg/7YIuDdEH3iioF5uyyAqxraCZNQDKjdYoRW
k9Ie6gVlevKc2lYnTFvLK/C8kHpYJcMnzeWavCJU/OhJB2KCOfccL/Ohd8uFhqvy
4UN4jor+8PqH9RMg5cLF6cqllCcfQQrsNpdPDENLapzEK6z3lULFdqriKdBfm7D7
XzkLVh+Cw8b8dBuBAYGXykI91iInSr8wl3fvmscwSfemhmLJcfs7vHkhIdGdbhNO
TDNARw40hUthHyXA9/L/KII4cfDkqxYQL0iVBy0wz5XhOgSpdwpKmsDVqn40Js7u
Grla3HC8AhTbeNzCzcUIB8CE2Cy1G1QG/Fv7tLeeijrzDF/9FN90UiEje/Gh+LrO
O/wBSRn8mV8ha7UYPXWQepRkf2hGcFSlJVWWA2GGZLam2RmkJxI94uqKMuP5E/gv
StbJQUknk6TelvXHfaIwzpUeQuPpoWsu0VWcbYfzqNDiHPuwnbWfsO1+gaRf8fNQ
DyyuPUWOgjGbkStyS+CMh00pYq2BtDw9yp57VA7HsO0O+xpXYjk7/uMFfI2yXU9k
8x183cW+3jXpcjmoXwgdFdGAIAtGFmvW6dLtLlDmrfQs63AQ3yfj50TR1IEcs9pp
`protect END_PROTECTED
