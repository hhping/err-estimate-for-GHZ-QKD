`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qu3C9Z8l5Qm1RVjsWF1cltb8mkNBujERyG/eCc8qjl4wE9SwyfROu0PrPCM8rTHT
hgxe1sEVcTjF2STbcwpAOneHBK7jsV3Q0y3553nGKezjjOesL1TkGAxoIJFwjCY8
tXLaCDbFkeH3Qhgpoh60VV0WnYg6ewo8c/AsNS1njj5N30rn4XUr+6ooePqI0poh
m844cnBPcRestjw+9TvKztgroDyqe+c7OcVqo1Bz0Vm4solQ8Arl3OjuW8YVMaD+
cx2XzAQDiqOqZ9tfBPrj+I8jKjFPF0r0kGIxoTb/5fbKTVfpwhPeDe84+bauF/UY
EU4rnnnNUqFBx7Gmib1dt8pO1OqxafGYMs532yFSvVbwFhi27jAKXzsDDh64ejD4
gdLHz5vlpKVkes+kF2hUpOdVe+ILxHqHnXsOBO4PS59gKkh9GJ61Ol0kbTE/FMzC
CeQ7nTIiAHSeZVAapVXWBJP5dGBFVNdungMu9hIPZvj6eamUFNkJC4lRFDVsv1t/
2gXdqzxGoccTjJamFmY0EZSj93zUFrqAj7z7FLEkU3ZFlJ8qWRCxZHhZHWPQmxu0
lBhUS/le0sZB3Oy75wWAp8HY7jrjZ28R95IKRgQSsAXxs/KLwUdPuiHRxf5w9Rxo
O5qXHIJbsOIjGciB/59q/+SDqlyuSZMMJtJ5EN+4/TvU88aZH/bQXZttm8ysYOZ2
EKWmtUMYlrsMSpGJEWU04JRS91eV236pFiXCwFqtkHZG5DKPAxYD8dT2+OVec9bL
nZeGkQALyNnK7t1ijuYsG6+BaVESc1212p4XB+nvpOxz5UNoK+IRLsrWo8WPaSwV
vFJ5WZmMEsW53oXE5g/X7BqIgJHGgZuy7v7tBl3vCuwXLfG12Ml0e8BXeSbXRK94
VhebUCDr0m770I23f+P0Sosre76yNjKtjyRgzS6/FuxQw3jBjREvJdCPs1bOUmbO
Hqx38yuAYqEY+oz8HGuu7g==
`protect END_PROTECTED
