`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmZmpDUKVtWpf4dQ+Eq4UY/M5QHP2PZOs49u40Rp2Cc6MVJVP9NnmgP41fn+tZ9n
ORu5HNEwRExBIiSbbPHNUdvls65BmNUlkM23H5/68t0su/srQcz/a2kfZg8lR4bG
ZEgVZMN+Eec8DquQM9zk3Gs62RRGaksvby/65CO7CGOOOdTUlgmoYXa7ptf3B4CR
vW+pplRf/lUTXTpcD8/wF3iji9/jcik/71NTg9iJREXpI6Ef2F/ps1T/LaCYPUgD
`protect END_PROTECTED
