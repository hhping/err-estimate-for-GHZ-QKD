`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NRJVMj3PH6D1mkXL1kLUMyKzn5wWGQVlzfR/MBw4w+zR00RojDAx1fYIKECs1lk
A7hCiS+VStGQO7bU7blBV0RZxk/6RD5e+AwrRVKm18MO5iCgfThXyEKq4t5VNOQm
juQafYlmwsNgHyiSiT3CFxk6bDq2p5dtTG2jklRqltwla3exH/RM67nMeuhmveG6
`protect END_PROTECTED
