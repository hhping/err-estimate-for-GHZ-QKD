`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+xuKPjsPdPwfqMjXu5KwG9pZcqbecEObRiNW4/H64bGzf8kE6w7L1ergZuCXTMx
WkG89AYg0YufSpA+nyrHdJpn3pkOPS9rnG0vx+72aHJ4MKaRboCLaOZRVBWQFOCr
Mu3tnU3miW14iTXa0AAKB63cQEB/IF0Vbw/tDBI63FGOLTPGpzg56NTNpKyfsML4
6Wdp/Fp//7jXSswp202J1xr9hDXkHeCr2WnEFRa0VxIJ+ZYH/y/KWzT9HkYa3WXY
GYRx4Ligm0vGCbisZBJ7lh65e4Dk91IquBe9Z1TZwlllHRn2EHvSdFe0FQfBKbja
IOTAoSU6xGTFbVxxr1Nl4Zew4SaJ0fwIT31SC2Yy7mAlVjaSkGnSd6yx4qrDXcHz
ZZ5dw4tBvMRz0saGyJO9stljngSj1+AWSOswp2aoDmWi1oFjdjj/wA4GJ5neejkx
MFjNKCl3B21OkmsSQSsYHz25ikP3qnNz0zD9EwIM0habP525GOadLAbg+mPQBfeV
mvULSfJfixpJPPI80jpK/F1IvWaiPvPvJZ5w5NuCKhGPINpGf7ApoISjzJ8MxhSd
gpQ3bSXn4owSEUcTKflBPq0NdnwTU/vWE8kHA+nPt/oRoM1x8cFMrmQFEqEdZ47a
zS6AknwAZkbIeSkkNufjsDYh9yLKOc2A0KoqEurRn095fflTDFBzmt3jYMBfuP1z
TvcpqpY3grddjUBMdZ4dgHKjt2vk0FsnaDsuqfNnAebm7oii+aMFnbYO4taJ4Qae
67Qqk7hSpFVKXH7H1NPNiJ23taNsdrKpv+g97OgnSD+279tra3z8U2W14x5fh7Ko
BhaH6BPzGketg/jVtOLJ/VrXD3KJ/86cJNSsvvgRoqmqlrX2P0Tb9AftJK9NkFJn
P4GKQWx0aQLeuVRdt+7r+1sUyJZ+zw3SlWt/mqBFXn+reB7yXLh++7zCF5Zzc6LP
/LLFIQpwOICcdrjdwFciBh++9oJsTs8KG1UVDOZM2nZxqgTXtMv4cFMcGt1NK3tS
VNW5oo+HmAryf/5f+LfiZQ==
`protect END_PROTECTED
