`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F5gDFAL/k4qMiC/Bjfqa56VT4YKLFXkXF2J1ja3KIa5+z6l7pTpdvK2zggGxv8Sb
kNUkkmxpnZ+PLcW33btSjv2J+TGf3+kbOdIBwowKGGbZJc4OVrroqotJgTCnoWvC
K/xcBG/ZN+SIyOlgy6Q0rxUjCu2Hp065wwvQOmis8xHCzrsfMufsu4kO0ei7A2jH
Z+E4AhnwOeKlGdQlKVHZ9YWDlh5eDNGtwiPqPrJbyZ5v7KliALv5rkOKup6t9pVe
ltpzg9lU6mLKPNpSu/r+GaLkdF4gnfTuzY/reKIGlG6wO/zfLmcPPyXTTI9ge+Ht
O5pd/MWArBpQtNEW6xZ9NgG8GKxGMOoFT13BDOsF1GZeQI3F0ojURwyP19EXNPmq
TCjHlGj+kSiWy67kQErJgyQV59gZP76v/koW1Q4Foha+VjCHzdqXKfQg6Cm+V4kw
IfTUOSzay/qFN/CFzLlJ534e+fef7OyWtQdoj4JdG3injSLKKjJyTlF2Z1mz0b6N
cl7xmWjlP4CX+OGkSrcTDd1U2L7zOW3tFLszCS413jQZ5nOw5a/gJPQspTrtjm+Z
`protect END_PROTECTED
