`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YdzVPeqeBwrvcFPG1HOD5kt4JFV0bbpvNTfFwP3CaC4XDamgMGTIWMxxAdS5Od+S
SHpm69Qm1u8XSacCPstyReJ414zjGxY3deSpSAplf9Bav2E7meGP4ixfLV7KIpFn
fH6J6zpwOLQBD172pZQ9dAZzisbjHkeahaZ3LyR7gGVjZnet1E+XqdTI9X2SrAVe
hwI0wxcubL53WBdHD3WIqjClNvIqrMhuG11HGbTIzxe9nDfUpoRKRK8sAkpO4Iec
Si4i1GOZy0yFUTKVyWVN8ON4kIt/4+DNmKQLZ24hG7ZDIy3AMug62Qt8F+50JwHA
zKn6SVlxasKMzpEjJ/SLCRF0WVFA6DBbijjkZJ5mTHHyrwgyQCf5Db0gyKFxnAec
OX152ivZKR471tVjFlTirw==
`protect END_PROTECTED
