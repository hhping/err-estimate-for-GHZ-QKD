`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/35bdJWRFCia4/pf6hMfPOdsmbQvwX2M3TSgdjEwyzwSud4RYIB9oOsqmQIIUG6g
BvezRg8t5hUJQALIFnNokiVr7SHxZelD/4lPAXID8hBgdkQhhA6fLGXx86SBms4N
tBBvp9E/3tr2oBPsLZUXKhCeOCBpFXjsURamAqJUSZ66YRDFYu7ftfEofD9oa6Er
kU8cHyydwri0f4+nkEYEt1YrNpcTKwuKLxuHC6a0hfDckweaSdzyyN1nwsizFI4O
ZTt7UuV62af+07ehvSgZIhViKjfM7uNVJ6X3nCb9ujEaU2j6GRihCL5PyM3d29cf
7nhiMsSaw9p6UOrR/Mgav+y+vaRUx0hrKoWL2Lp/vq69agCoQA5BcIL/ZcqidEEx
+sCJV4zfAXQEWuHjoZk/Tjo8EF3vLXTTgtJJgvB4QIUND1yley6G8WBIvDJkL9FB
rwGge9Xgc7QWKsKsOyTfnNk8+YooUi7Y0BdkMj1KocjRRLKKfDSzJT4o4ukVkCcn
3G+2DG6UzaCZrHdJbfBV0mOew3bdkNVkVI0vrGiJjv71Rx6F4wOCF1Kou6U70kXD
Iifq+mXZn51g43nSY6qToiw+zWpwFyGNnPhWSwnQYkQoB09xKyzx39r9njH9hWLZ
rYNK2fWIFmBxCVpJmUEmAGMoHl8+Q+y1uymts3cb0MT+VdQTU+OBtd9d5lpIaIAr
E7H5EbNXc91qJvjcxMdSqfJOS9sdEHcBD6CpnEOf1tc59I+/tgSwOWwObzenbRxD
nPn7fqmd0QFj2oeQOlt4S9h+YCqBW3I/RZ1sU4PV0NVOxERrVBmi6ZzRX79O7yEe
yI9fTyuLVAE6tS85k19nHGfbA5H3Ez/6g+Gnxe+PZlWFBD0oChVpEMqaUBl7kVq7
yj7p8WJEZie81IW3+uc0eYCtpH7RL9VrGm+vEC+HxcrNZa6yabbSlfZsR6UAZ1pL
4lfESpb+Y/F3d4kFEw/cCBeU/iqZcMNVUomck0pL1g9pybgG/vka9r0ufBponi+z
R3ArYc4HcpPINTEET63FwrvSYzbiDFDLWpo0aH2mYuB8EatBvX8v1SfcdCw8eOeQ
xnDRLVQv9/LTnT2GSDZ0/UVrwuYLCp4kJKbofS54hJ6JQTCodm3GohnHqW/Ij27C
Mix9EfKrol7acXKGv8sLoY2loytwUvRZxfJ4qxrMObVWSf3XouyytMG1whzF2w5u
84meI7Ftl6DGFa3zHGnrAQXE4+Hr5g/SOuyoSo+LpCD+7fg+iWVvLt+cz/uW933m
V4rgRyq7xetrrbRcUGgylMNDjxUiZBPuH76h1DBWoQHTHYKH4te+umrOWjNBhS/I
Api+sNob5WuocX0EWlyNYZWzdS6aecGtdL3hcvWeB1h0uYO1pCF282ym5bHv9GvK
96sMm7WZsqYXmUcdU8rWHBEk+4q/qX5ip+DV8tWO859SJ/9LjG4/VP5alPup6UsS
dGYNdqqyWHqbA8Nmv3YJNq9DL2YkDcJm6EukmWJIM/Q0rd/z754zrxAyjOmJHJGn
wGF5+N8zgSh3UDPv6aZ9o4YUPM4xpBmhEhqfaYDXhuKk+PwoGteZWSj8DOKbzY0b
l8o/ji8y2LrGVaUv1OhHM5WKck2gHYatB5XsJPQ0zgr70/t8I/VlYAM04ly7/cKD
jId2vncuobHUWLtdU4Y4xrfF+7LeOcfNDjfUjx2/KLMQYfhi41aJiYo5LmAJdCHu
2ipr+Nm+3slEi12UQZWhAzeHoerNx9dVZ+K/VpgAjg08/y28S6JHdpyqfzlqrAKn
kKAzc0WEbKKci9CzUNrO+t9CsMdfJV9IPY6G+7yQro25mCIYcDqPenXlvR4zURzr
ksgy0LSIo65ZFPDTiq/sZ/ei6VF7+zzU6RH1FxyYXVFN494638nnIUDAQyAEp57x
PwVFhJfLKsRGeZga/e+JXnhgod7eFDZn6tPtKHtKoJWmMF65JetsihZY339JXA2h
`protect END_PROTECTED
