`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+9Ii5sesA8HMwalG7cScZy7jcs35Npr/xdPq/0PugMBFIPXpFRawPw80LwX9qNiz
ZYpdSpfmqd6SO82XKqWVRRmoO4BXSI6CsdWMcjXZYNN9g86dY5GZWjQIdTLbNjCa
EJvCiXJzzxbJrZ1Gsuu3h2Lvm4+5c0xXQwZQHJN3fu/zgxv9MQVXNHorI1Chj5mn
Meutwzb/eq8e0cPYFAdiYNBwa7pA6xTmBxGTOI/MP84G79wTp2IzBmq6Ogy4M1Qy
obacW05am/g9DGwZ8KT0vuEn33aNcJp8Ox29ihds5upzHXCZOKQpKmeqyVVLVp9B
9zsa08D6IOMm/G1RozIutRZ8vLPWLBs7+4v0tTr/mxqih/y75zh5xxOVf/uLrOo9
BwGC+VURuYdlwk4ginXt+g==
`protect END_PROTECTED
