`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VNkbSo36JT6NbyPYFGmdG8PtYcMmD3sZePibfbFVuaW4joar0VkyAgy68Fib834Z
B9z6Z0hX9pfGSp+kKjOK0cSF7NBdF5qMMOzRylZoJMwh9xvfIW6S2agnyvl3W7g/
F0fYCrCxTSqVITtPrvUxVk3ubG+EIh2biG071wndN8ueslIHzOVeoVhWGTl+RMjf
EkwyjCykWPIFky9oaxxrIief5xjSbmK4Ef0eRQ5G9PwHrRHyP3dJzHW6Wig+u+y1
b4knouaRNvNi9/pqvuBNHOdq50fzr/mEn9vPlCm3xArkRGWOjHhDVatiJQ0iQ4a7
f/Sh7Lw3tlX7+LVkb5SQOt68LBhaWRNGbM095i5yrJ/9x5Lcpi4WaicPcoemHVGb
hHvqbXovkYlv0ID5fzu7QjD/IrRLBqQgACrw7+AjnuhgEv6O+/FyZz9HeNoQm3fm
NQSrMyJ2/3wETB1RbUiAPGa8xJ75r5Z8OfvwKiHIzcG9BUzWayxBbm8UZGGPhe2k
kC3mJvaV++MJjVlEVcniQLTHyAN3cjtFchniVNzR+PjB3Q7L0fwZvnRyTEc7Mine
EjoVKAN+olZwBk4owZM49S/nyTxYUSUi8lu1Yc7sNlILGJFeetYQtkzJEuf/737i
pT/7BJ8MyOaSYoYcY64YxBYgP0cxy4PY/h9nGpvc9vF6m4gMCs62Fe2xG0YJ8MHY
t1XX6wpkjWF9ZWAPzftIGUs+pY7hj57yRs2gO5c/EfJExxBX1t0Yy0HVasWVEn4n
HnhwTjLzyk5Lv5v1DHdt0zGu2l/E7laBmNU47BgVxBG3LE6TDaTMCxBQctRYRl9b
LjFSWXu5CAN8CieAzTyAVVobDWaPCz5Dl/ShE55U7CkX4pJF5gQBukRHFtWTccqN
OUScjHqweMwCBg+gh11tb5ZJ1LgtVrQ4oEMIZh37NIZXIjMhqNPaCI10FpW/GlO+
kGVT2dDVhue7M+uetZJ4S5yLYI+FmHPhyx4t4x71GK0=
`protect END_PROTECTED
