`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rq27vzXBbQE4GsjGWEv3nrpHmclp0Q59t7Yg5+vfnPr5JT4ITmO/FsDAPrA8pZ7q
xsPRGmuIpj2Ujh/g+6lAiDAR5sPlPuePtbO7WalIYrUlbTBKLdUWU+CIjLFbVpaX
wXC6BneH779EiU3njuh8iYXvdfvXDZsfaq+UQ26O8ueIPRaW68cyaUynAS3adLn+
rcT4ZAmwd4AfwqWHcoxM0jk+BFd7JPIUUS3azLMoQ9r9/zrH5Z1Z9lnqRorp++gn
kjWWXjSwSLvgiodmWnQS/wM9yBDuUlqcEn6Gsxq6ERB+DOioeD9WZko1A8aWX6PX
gSdX6gnPb0P+9JgRrAEB0sHokbkV7P1pFPuOX23DM2f2cfmGo1Y2NQnf05KoRE3N
oYhMTYgb+0haeSE5VdtVX+Nf9/twFJ3pwyQwQZGMVJwBoln/TJRX7bzn1VR756Vh
2J6t0aO/OylVIFOQwOdsC2Utn9m5GYKTRgSsOMm8VrEZmZOXMoO1+NoRZBajBBy5
jhNJOrjfc4ypVUN3EBykEO1hhDZuRqnXWHImVaKbcZKmR3wejEV4Q4nGKjYwfcaN
OK0ZqFisPmzC5a/V89UuZop7Ds09z63zeBC8wr5LsaI=
`protect END_PROTECTED
