`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rr959xneveC+sNSoAZGBjyubSGt6ZVTJCrK8JBQ1qQf128vRs+WcrJNDKBUgokKX
A6nPsIHjYIP9Anew/lL+S75KkmcFuRT1XnEBLothjc0qteVlIl0NQpHwJzRTt4UJ
niIcwyhofypS6tm1L0scgRH9GgRkdCMGAV5HuYkLoG44A2y59aX1rEhiJ3KFTiCM
OxHlGsf9n6Fowv+SfB/oUfYOG0f5TXO7WfWGxQC6vAaXCevP15ZLdSy7nJJoS2+o
rWfok8p3RUMyKxKwvWAw/YZpIVlzkAJ+we+wP8WUIDnfuYL5+usq6KPJGmBsSfQp
ZcfYrFhKpdfJfrchaw1BW6nU9xso+f2MVycsIMD1ChLWPj2yTXgeuGBlxSU2s380
VsbbtacscVMI6+4kDR0HrOag124oAEVeJt5ktsBDKtNtWBXUpS8+P43QK4eUPBCD
LTW2NWYvICWo9TmwaFL563FcrHcBvSA97M24b+EemyX36n83uSlvTWvpKabI57hu
G1E1YfHJEC4vNPp6zdyVLsYBTbeYELk6qzOmJzkl7+7j6sDK7sLtXw4A3aIadn14
Fi0NsGMWewB4c+M6KUfbS1IJ350BD9cn5kNoieVYqHBKqAQtQhfdJlsmMyc2Ge/+
HlNjpxfrrve9sRJqOk1KxxLPSynQg9G+7p4GSrrbTdQ/TBakMNTKDynSNGlq4Z6v
2h1sooQbldGmXzyTrwKJK6gYwP9ZxrzRC0nPOenmZQ5E2LD8eRIy2Hf/ZsUf7Mki
4YexaG+kE9YdwfiWADEOLFfG6/P0BazqhQWJaTo+xXzpdzIpIdSJ74ofLHaWrYKC
EMuzuPxR3QzArbLFL8qsuc2ZZKI7cS4LvSfotq0xV9yIyHFF+EWR8MwvXduaFMNN
yhFR2pKjW3YFzTjcU2v26Qw3gChqGPhWnY+uygWfKsA=
`protect END_PROTECTED
