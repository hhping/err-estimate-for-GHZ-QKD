library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_tx_buf is
    generic(
        enable_debug_info: string  := "true";
        calibration_en  : string  := "false";
        calibration_resistor_value: string  := "res_setting0";
        cdr_cp_calibration_en: string  := "cdr_cp_cal_disable";
        chgpmp_current_dn_trim: string  := "cp_current_trimming_dn_setting0";
        chgpmp_current_up_trim: string  := "cp_current_trimming_up_setting0";
        chgpmp_dn_trim_double: string  := "normal_dn_trim_current";
        chgpmp_up_trim_double: string  := "normal_up_trim_current";
        compensation_driver_en: string  := "disable";
        compensation_en : string  := "enable";
        cpen_ctrl       : string  := "cp_l0";
        datarate        : string  := "0 bps";
        dcd_clk_div_ctrl: string  := "dcd_ck_div128";
        dcd_detection_en: string  := "enable";
        dft_sel         : string  := "dft_disabled";
        duty_cycle_correction_bandwidth: string  := "dcc_bw_12";
        duty_cycle_correction_bandwidth_dn: string  := "dcd_bw_dn_0";
        duty_cycle_correction_mode_ctrl: string  := "dcc_disable";
        duty_cycle_correction_reference1: string  := "dcc_ref1_3";
        duty_cycle_correction_reference2: string  := "dcc_ref2_3";
        duty_cycle_correction_reset_n: string  := "reset_n";
        duty_cycle_cp_comp_en: string  := "cp_comp_off";
        duty_cycle_detector_cp_cal: string  := "dcd_cp_cal_disable";
        duty_cycle_detector_sa_cal: string  := "dcd_sa_cal_disable";
        duty_cycle_input_polarity: string  := "dcc_input_pos";
        duty_cycle_setting: string  := "dcc_t32";
        duty_cycle_setting_aux: string  := "dcc2_t32";
        enable_idle_tx_channel_support: string  := "false";
        initial_settings: string  := "false";
        jtag_drv_sel    : string  := "drv1";
        jtag_lp         : string  := "lp_off";
        link            : string  := "sr";
        link_tx         : string  := "sr";
        low_power_en    : string  := "disable";
        lst             : string  := "atb_disabled";
        mcgb_location_for_pcie: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        optimal         : string  := "true";
        pm_speed_grade  : string  := "e2";
        power_mode      : string  := "low_power";
        power_rail_eht  : integer := 0;
        power_rail_et   : integer := 0;
        pre_emp_sign_1st_post_tap: string  := "fir_post_1t_neg";
        pre_emp_sign_2nd_post_tap: string  := "fir_post_2t_neg";
        pre_emp_sign_pre_tap_1t: string  := "fir_pre_1t_neg";
        pre_emp_sign_pre_tap_2t: string  := "fir_pre_2t_neg";
        pre_emp_switching_ctrl_1st_post_tap: vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        pre_emp_switching_ctrl_2nd_post_tap: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        pre_emp_switching_ctrl_pre_tap_1t: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        pre_emp_switching_ctrl_pre_tap_2t: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        prot_mode       : string  := "basic_tx";
        res_cal_local   : string  := "non_local";
        rx_det          : string  := "mode_0";
        rx_det_output_sel: string  := "rx_det_pcie_out";
        rx_det_pdb      : string  := "rx_det_off";
        sense_amp_offset_cal_curr_n: string  := "sa_os_cal_in_0";
        sense_amp_offset_cal_curr_p: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        ser_powerdown   : string  := "power_down_ser";
        silicon_rev     : string  := "20nm5es";
        slew_rate_ctrl  : string  := "slew_r7";
        sup_mode        : string  := "user_mode";
        swing_level     : string  := "lv";
        term_code       : string  := "rterm_code7";
        term_n_tune     : string  := "rterm_n0";
        term_p_tune     : string  := "rterm_p0";
        term_sel        : string  := "r_r1";
        tri_driver      : string  := "tri_driver_disable";
        tx_powerdown    : string  := "normal_tx_on";
        uc_dcd_cal      : string  := "uc_dcd_cal_off";
        uc_dcd_cal_status: string  := "uc_dcd_cal_notdone";
        uc_gen3         : string  := "gen3_off";
        uc_gen4         : string  := "gen4_off";
        uc_skew_cal     : string  := "uc_skew_cal_off";
        uc_skew_cal_status: string  := "uc_skew_cal_notdone";
        uc_txvod_cal    : string  := "uc_tx_vod_cal_off";
        uc_txvod_cal_cont: string  := "uc_tx_vod_cal_cont_off";
        uc_txvod_cal_status: string  := "uc_tx_vod_cal_notdone";
        uc_vcc_setting  : string  := "vcc_setting0";
        user_fir_coeff_ctrl_sel: string  := "ram_ctl";
        vod_output_swing_ctrl: vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        vreg_output     : string  := "vccdreg_nominal";
        xtx_path_analog_mode: string  := "user_custom";
        xtx_path_bonding_mode: string  := "x1_non_bonded";
        xtx_path_calibration_en: string  := "false";
        xtx_path_clock_divider_ratio: vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        xtx_path_datarate: string  := "0 bps";
        xtx_path_datawidth: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        xtx_path_gt_enabled: string  := "disable";
        xtx_path_initial_settings: string  := "false";
        xtx_path_optimal: string  := "true";
        xtx_path_pma_tx_divclk_hz: integer := 0;
        xtx_path_prot_mode: string  := "basic_tx";
        xtx_path_sup_mode: string  := "user_mode";
        xtx_path_swing_level: string  := "lv";
        xtx_path_tx_pll_clk_hz: string  := "0 hz"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        bsmode          : in     vl_logic;
        bsoeb           : in     vl_logic;
        bstxn_in        : in     vl_logic;
        bstxp_in        : in     vl_logic;
        clk0_tx         : in     vl_logic;
        clk180_tx       : in     vl_logic;
        clk_dcd         : in     vl_logic;
        clksn           : in     vl_logic;
        clksp           : in     vl_logic;
        cr_rdynamic_sw  : in     vl_logic;
        i_coeff         : in     vl_logic_vector(17 downto 0);
        oe              : in     vl_logic;
        oeb             : in     vl_logic;
        oo              : in     vl_logic;
        oob             : in     vl_logic;
        pcie_sw_master  : in     vl_logic;
        rx_det_clk      : in     vl_logic;
        rx_n_bidir_in   : in     vl_logic;
        rx_p_bidir_in   : in     vl_logic;
        s_lpbk_b        : in     vl_logic;
        tx50            : in     vl_logic_vector(8 downto 0);
        tx_det_rx       : in     vl_logic;
        tx_elec_idle    : in     vl_logic;
        tx_qpi_pulldn   : in     vl_logic;
        tx_qpi_pullup   : in     vl_logic;
        tx_rlpbk        : in     vl_logic;
        vrlpbkn         : in     vl_logic;
        vrlpbkn_1t      : in     vl_logic;
        vrlpbkp         : in     vl_logic;
        vrlpbkp_1t      : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        atbsel          : out    vl_logic_vector(2 downto 0);
        ckn             : out    vl_logic;
        ckp             : out    vl_logic;
        dcd_out1        : out    vl_logic;
        dcd_out2        : out    vl_logic;
        dcd_out_ready   : out    vl_logic;
        detect_on       : out    vl_logic_vector(1 downto 0);
        lbvon           : out    vl_logic;
        lbvop           : out    vl_logic;
        rx_detect_valid : out    vl_logic;
        rx_found        : out    vl_logic;
        rx_found_pcie_spl_test: out    vl_logic;
        sel_vreg        : out    vl_logic;
        spl_clk_test    : out    vl_logic;
        tx_dftout       : out    vl_logic_vector(7 downto 0);
        vlptxn          : out    vl_logic;
        vlptxp          : out    vl_logic;
        von             : out    vl_logic;
        vop             : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of calibration_en : constant is 1;
    attribute mti_svvh_generic_type of calibration_resistor_value : constant is 1;
    attribute mti_svvh_generic_type of cdr_cp_calibration_en : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_dn_trim : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_current_up_trim : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_dn_trim_double : constant is 1;
    attribute mti_svvh_generic_type of chgpmp_up_trim_double : constant is 1;
    attribute mti_svvh_generic_type of compensation_driver_en : constant is 1;
    attribute mti_svvh_generic_type of compensation_en : constant is 1;
    attribute mti_svvh_generic_type of cpen_ctrl : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of dcd_clk_div_ctrl : constant is 1;
    attribute mti_svvh_generic_type of dcd_detection_en : constant is 1;
    attribute mti_svvh_generic_type of dft_sel : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_correction_bandwidth : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_correction_bandwidth_dn : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_correction_mode_ctrl : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_correction_reference1 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_correction_reference2 : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_correction_reset_n : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_cp_comp_en : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_detector_cp_cal : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_detector_sa_cal : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_input_polarity : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_setting : constant is 1;
    attribute mti_svvh_generic_type of duty_cycle_setting_aux : constant is 1;
    attribute mti_svvh_generic_type of enable_idle_tx_channel_support : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of jtag_drv_sel : constant is 1;
    attribute mti_svvh_generic_type of jtag_lp : constant is 1;
    attribute mti_svvh_generic_type of link : constant is 1;
    attribute mti_svvh_generic_type of link_tx : constant is 1;
    attribute mti_svvh_generic_type of low_power_en : constant is 1;
    attribute mti_svvh_generic_type of lst : constant is 1;
    attribute mti_svvh_generic_type of mcgb_location_for_pcie : constant is 1;
    attribute mti_svvh_generic_type of optimal : constant is 1;
    attribute mti_svvh_generic_type of pm_speed_grade : constant is 1;
    attribute mti_svvh_generic_type of power_mode : constant is 1;
    attribute mti_svvh_generic_type of power_rail_eht : constant is 1;
    attribute mti_svvh_generic_type of power_rail_et : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_sign_1st_post_tap : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_sign_2nd_post_tap : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_sign_pre_tap_1t : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_sign_pre_tap_2t : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_switching_ctrl_1st_post_tap : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_switching_ctrl_2nd_post_tap : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_switching_ctrl_pre_tap_1t : constant is 1;
    attribute mti_svvh_generic_type of pre_emp_switching_ctrl_pre_tap_2t : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of res_cal_local : constant is 1;
    attribute mti_svvh_generic_type of rx_det : constant is 1;
    attribute mti_svvh_generic_type of rx_det_output_sel : constant is 1;
    attribute mti_svvh_generic_type of rx_det_pdb : constant is 1;
    attribute mti_svvh_generic_type of sense_amp_offset_cal_curr_n : constant is 1;
    attribute mti_svvh_generic_type of sense_amp_offset_cal_curr_p : constant is 1;
    attribute mti_svvh_generic_type of ser_powerdown : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of slew_rate_ctrl : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of swing_level : constant is 1;
    attribute mti_svvh_generic_type of term_code : constant is 1;
    attribute mti_svvh_generic_type of term_n_tune : constant is 1;
    attribute mti_svvh_generic_type of term_p_tune : constant is 1;
    attribute mti_svvh_generic_type of term_sel : constant is 1;
    attribute mti_svvh_generic_type of tri_driver : constant is 1;
    attribute mti_svvh_generic_type of tx_powerdown : constant is 1;
    attribute mti_svvh_generic_type of uc_dcd_cal : constant is 1;
    attribute mti_svvh_generic_type of uc_dcd_cal_status : constant is 1;
    attribute mti_svvh_generic_type of uc_gen3 : constant is 1;
    attribute mti_svvh_generic_type of uc_gen4 : constant is 1;
    attribute mti_svvh_generic_type of uc_skew_cal : constant is 1;
    attribute mti_svvh_generic_type of uc_skew_cal_status : constant is 1;
    attribute mti_svvh_generic_type of uc_txvod_cal : constant is 1;
    attribute mti_svvh_generic_type of uc_txvod_cal_cont : constant is 1;
    attribute mti_svvh_generic_type of uc_txvod_cal_status : constant is 1;
    attribute mti_svvh_generic_type of uc_vcc_setting : constant is 1;
    attribute mti_svvh_generic_type of user_fir_coeff_ctrl_sel : constant is 1;
    attribute mti_svvh_generic_type of vod_output_swing_ctrl : constant is 1;
    attribute mti_svvh_generic_type of vreg_output : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_analog_mode : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_bonding_mode : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_calibration_en : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_clock_divider_ratio : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_datarate : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_datawidth : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_gt_enabled : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_initial_settings : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_optimal : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_pma_tx_divclk_hz : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_prot_mode : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_sup_mode : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_swing_level : constant is 1;
    attribute mti_svvh_generic_type of xtx_path_tx_pll_clk_hz : constant is 1;
end twentynm_hssi_pma_tx_buf;
