`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJoosRNQdvSAoZl3w+Qmbha6iO2sJKoRIhxt2AEUOSt+gKg8AkFteIgO+PMZW89e
P02/f5CWJL85cl9a8mRV6g1JOaEU2O2vyKlK+TuOiPK6BP4y47KT7s1V3DxEUgUh
HKFChZc9j5wNdfXXq4CricSALyJ+hBB6se7lH60j16f+4+DaMHRKVZ8mQA5DHbsZ
9IRFXnMBkAJL8Mm3b2Cgirc186MESL08Wmqs12zSphy3DsHF8qbDz66gZ1H9E9u1
s5bnn1WE+AWPnjeGewcVfVq6jrPPKJgSJFLLraJ4B+yneapt4sG31TsCxFb/CE81
LzFSD//1qUpwU5VbI+489TJh6Jgo82wMh0y5NGDwUxP2Eo9Yfv5dW07FO7PN8erX
pRy9CqrhorXktOWvMKDtfyIDmd+ZXMT7bHAnSWzqQRCp9TMBG1mCXRCXwkhbIX3l
f9M2Ttgi7fnF/WxleyjkieEPGCyK9lgxjJsdnVogx6NpF/EVreZXWFoZ8iHiS7tc
XVrKEAB53QKirWsZmV5lB4bnRgG3yuuxnZqdMmiiOUUxB1TShDwS2NDZfd+PTQUA
mUyxC5wmUuNqIguxzarK7bP7JDFKKm/0qlhFfKzEib7Sw9LVEcVPUU5mVyJk56Lg
Utx2AtFRk3+EMA3nGXQdf1goBQdOBuEfu9+CZqu3T4Ewt+g8LEvqaXPn3KauvX0o
mj8MfvUZ0G8xIfuEHC8HNdy4TmwYYL4XdqWPMYW6FQm7o7tZBX2kRv7CbToLVp7C
Numl80WmeMQwohdRzzxZpC9YMiS9GPzc7OaNaenb29PahHXczXl9rZ5jkfJeqKwq
heiGsynKjEP5/QejEc9CYq5zF5ZhIo7s4yrcYUvGhj1juXB7b1a2ut2yN0ZFBqXO
MBWvxAgnCIJwCBGYppRZDApUrAxgottWX1PdWIAikOs0pYvnv8fE+R7dWvLISy8m
+2k3O+4B6X5zl8ZYhcIFPhb3MMntDYtq45KUGJ3x9x57XDaE5zQqUCTyYRz9vsjc
XObrea/MxMkByCo0E0dIXXlaKZOdTQ+hzHT5YFGe1mVVDYfSt2m4pp0XY/9px+6j
L9vWG0Zr+AbeM0P54RAOnStZZG6/Q3s1x6uq/9iO04rqP0sxyCiz7fnu7j+clwgd
yHxp2MA47A8f7rVgd1rhGIRI1MSDjyWLb7PGFuj1Geg7csXwpvjNtwLzsE2ijdYb
OrnitLG5T836Kgi/wHW9UpFp6zextvtac/twTFUpy4PIbxBeSBQJvAg2BVSDQBDs
yNPlOlcYZ4n/R5uX9Z0l+5qKuvoQPurGE7TzdeGStd6WnoO+OnS7vhXK9OuwVE04
umOiLdRzj728C2x5Z0V0TY6iozEgcFqQkrfZh4y9ilIeYMfv0Q7SHU3+J8JGjkjK
RSy+TyDx77GB0Uq/BhpDppEnt9E4SlLFRyG3jvIGl4dEDlyrfb8ZOvf+pS+DZjqQ
uDrvgzkUlfoG0NL1VWZBUSJZzDQnRvNeTqxHGkgpbvpmpCDjZ5hJdN18/A1+NNkN
Yme9Pm2jnFYz06Rq16ZhVG8AglO7peYftXjjwqAHHWsA5EhlX42b63hr7EcaeuHX
j9VqaalDSpq1Ub8HfYe2V51mlY6rC7kHadVd+pkx7zOKNACq7cO6Hj/iz8F5xlOz
PPP6xV6AvRz2PB607hJ5o4BrO80QeR+dG9rL1NL9kU9bv+T8EfkdXHTfsAeybDzX
Of+n6mOtdpj6C5uvbRH/kqrwJrxPfZA6LM97Go+tZ0PXmAda8ksi1lcV2JA4xMdK
ollQGnjBjoEoLDa27IrPfeiWxJ68nM5345xAnPhhT0ZWuixIdM+CRpvvQb7VDDAB
/fCJbefQ4tN2DDd2UuthHcGxFNdnYkGYkeQ+vekuh+FDN7WTdKKFWbl2NGMVZU29
uYlzKcBjYn4aOXeLMwEgGq9rkC9YBhYFcSZl6O9ZxcIPsVLXpGMK+gfxiawhvgAl
xbJZRvrS20dWAGx7Iw3t1wg1XsZTjf+X+bNBkbjfDDcKnW9dYgcsYYHPAlwIYruH
FB0BdL2VzhFB7fa5xeNCmhuDJk1zuaq8xDBnn2PYmo5ZBfBl6AK7rZu7rtjDLkI5
CuhXHX+Ht/nLE8B8HsdA/i7eFT3z+6RPeiaLbL6MEWLRbvPuH9aswiZyueLCpBBj
f+4JImSM/eZVUoE6Yl44bz7HhSzhD+odnMp492aFPPphReZG+xZNBF4jFpO5uUH4
9/R2v4pKu1Sc2ivwHLL7N54DnTN5CT17e0yLA/+pn/cyuFGSYrTozpp+sKZHp6YJ
5mmG1j8Oub1ENQ7us/dOucXF1wVST2HmQekXZOD6+TkDUHHm8+dvUC925L8zrK8x
ZRFnfmY06B2bI/UYSx7m1UgTTh68umr7xRnvaArvyyJpiCtYyULzm3ygObGjrdCm
f+5lMIM5HCVDsl04AcGkmQ6d0II80vF9KfJ98mceWqWRLpNAYsZ+49/Kqtv+N8iW
2HRuxNdp6LWzA2jeFm9ZfCHihS1snqqC+oTKPoLU8Gtozm4MEPmJUVQTbIvkY+UC
f1md9LDTcxorkuiuSG8ro9gZxBbK6MiOvtU85P+fhRPvWZbIoaAn8gJvZb7m47eb
wSVgFgk/26VuMeQW+1aO4nPbwJ2j28FVEw00ztw+IP6w8E/j9hrinelkVDzjQsfx
/EGiDkWaDh3n/S95Sh4eG1DapV1frISuAVHbYjInMC8vep/WFdXpLFiBM3BY7olj
0cYCxyKgXL+JjaJIFEtBpNhAP5UVO9+VLEPA/bQ9zzhfgGsQ+/sv7rKYFWvPPVW0
JCVaeo3KMmlYNT3W9kcOl8VM619TUsTj9NPgJii+zoqHCL9kTNLdr+A57dWKG5lz
VBObhn5x6kGEJiuv5gF5ZHBFrj2mdSmy65PPZ8v6qumEaJZs31Ozx+rcVQdyIb+K
zbTmdP9NsZZTS8zqGvxy4GFO3N54sd4QLUAX3Z+XWK8cdHr101PekCRo6lT8pLRZ
gSqbP+PbEYpMb1x1+R4+j++8vvGarbwi/lO5UC7l30FEplLuAj9y/LrIoibAsIi1
U6tXkFQ/vOhht3VbnGEo3O4H2OdDglBeoSu2dSxeWIJ6RDs3nFc3XdWExeXBNF9a
HDgVcGg/cFrxIfX8vye37WyDpqI/w5gn/BtsPbYGTK1QQiIc1DlRR2/VbTfFqqD8
lsSkdY8Yzubw+X0NbWnmBkW9Uz72G1QjHDH1mcGcOFuB5mDFyrl9L3HuYXZaZ50X
sVKbaov5JpHpPsOpDFC4Gl4W0l0pUxl6Z+ticrFZKi0qud12FaiDrM4guJYLiEhF
YWzvHde2Eryq1nPSUVRr4z0qIZxtkK+u6CiZ7Z5djy1S23OnksLGsMmOHrW9CHHi
iH2DUBUTz6bIjM/qN9a6tGsEcL1KZ5Xc9qsmo9sgu0GYzRuvnacEd5bttnIy0BfF
D+1oVRGPwsgC10K52VPBzagQ25m7JF7WoyQ61hFFMVZa1w8XA854P/ztYwNKRibi
oGnyweIqJd1HT2u5M5+NT0VXEZg0HB0AHDI0wpJ99xf9F6JEFNZ4PqQkSV7qHT97
evf3SkuDLaLVPu5GzmO7l+xlewzi4MF8o8PgFdKPqSoSB3CY3R0RzaaCQjjUtJi0
YgzmgRynTeHqzNgADeUG2fsQWgxYhhu6OdhNFng5tV4lhUxjgRomNuucTkK380eb
TX7XH1QygHsr0diUC4DWQtAI/A3nJOkoyJL+g7s9YNxNaEXtQ88JRBRa+LcufjTp
i1NuUxMlRifMYtmlbpF9Wn6laqoGtXVb4WfynmyYu3MiNa3vh2pYC6AvM24XxZNo
hxp56Lr0opoqUKOfDprZMRqPtvj5JqLdWttUI0pmTsPtOnYaA8yxVUqCmse7WYhB
wv3H9uByYMEPNbjOF7rUJc8QlxHLdre8CW+kl7NzOdSBnCuRuq6uaWsHh2yOtAh1
fnyO1gRfiqgayB8Pc02yaVv0rFdC242P/IWuzA22uxyypdn1OCwCxgMhZmK8aZf8
auKloDnjH4ebUQ6aNCCGNR/7i8Xylth4nn7z2zg9eiLLki6LCPlYsPZhRh10iUyN
F9+pvkpQU//SqRDuurqXV7zmSorha3lM2ewh6+fI41xdkN2A8AmBvsK5Ygj9A7zZ
oSLcv+bfllm7AXFRoHLUGZXTyjB0NVURa62YokLvLMipJALXjK8S7iK42qXmi6Lt
E0ekVr/h1NP/SoybYILGKULFKujPwO3Yi7MmkFppdsIc/d5DUM3btsfSRSOnyBdL
TtPURP0/zxt0qmxVct6lBXmGOyKOAHCRunRzgCLTxcoUgmLxS1xLsNT+XrAac+pG
eC0oCnusLCnYUDnzpaIxuW6J7NvbzeeXUYz2Dv+z2QON2A85mmTiM3YFWWdmLtic
JaXY10BYKCOFuRhvMK5Cw10JH3bmyUPmzJDfiZfbQBPSxxWZJW6hA/ulvmxeOWR6
pXlpiFk7jTsCHf0cjRujd69WKu1vt1E7YE2S6fTU+fDtGukR/AJFdmGBdTN6T4Gw
MXEJpTozXoAZcJyypXF7OMXysScApyBhojIHPF7FOcH31hoV1UUPDa+e5/NgFzMq
0DIIcNm9ndoM/WwrWW4j6W8RScQGkHEb1iDIX6du6IvbCdDtB3QWTvpWqpHjHO7Y
HMlEuKqUDdofxZ+LhtyEE47vXKLUnz4cSWlklpdC95/KoGEqVNJNQJornFQYs1qh
FxQ1T+ZGURJ5fgqxCTFUrhkGs8KmeZ+l3YeTHUhUJb/baivtf2NUiColE+H9Rnz5
U4DuMOMTyihcCngbVaDArCFPP+/wXseEIay2i6X0PwcYVag+HTFEHGJjG7oyEHYh
uuFd0QGieDLmWm+A37NiBd949HReiRVWQNKCFlFPRPIsCbWWzlGH6S/U97uvzl29
8i1O8n2/lBbv3rwIySHS4KuXXc9xvpKvY+7GFildZuuzuyGkSMac60jW9jAP+okM
OBXuZguWxoWWgxa6EtJGjUTqrG51IXVviczV7LYdsHc2Ofg4oh5GRjqtMTzWh6F0
HYdCqR6/v+BsqbIaf+y+yIrrU9X6WXyjY/MpR6nhYd4laPY8d14aVumtvK9BoAT4
x1tTn/ruZd3vvN07Pszo9tuHwoDZpJNagz4EmOhGw/sxgFvmVfcUUqfBFrPkDYu1
+jUOFXREtNYqkM2T+LJRmOIek0IocpdK9MHz/Q24SFIU0fniEr3FTsPdxq3/HOxv
Ag1Uq3wHhnyaytNc925hb6sHeIqX9AVg2AwlSFqEvA7jxei848mXZB/+5nS4QuHX
isTEjDLySJVp9qBOjElIj9GMtrKdOJSj1meqGERYnxBDbJArTqIQR9m4LrJEG4w9
TtnyXWjS53DYqxdhgu9shZ8ui+5V+hFMQguEcbainhgS4Zbn+60ftvlilYxWNVBZ
0CveYXdasH77L3wlkuaj1KoNOsImOiqUirY7BOg5qhuhQc5LuvIotdP1Rt3uqYS8
HWojs4beUGHZdpdJfez/cm2zbJysNe+N/UVfv8OXRMbIFXqs5K6jh3ZVBjFsCBJf
YLP524ctH7/dtD1xeDq7ADkjqlxRIcVZUEgmsfoO0vtbuInteLtnJwOMQsFOnKkt
L03DQRta3UOQHT8okn1isEGT0uRvfpi8Av7DPoYuG0DEO1k4wkbw25j4b0NuR034
W5jDd8Zo6Ub/JYYJMcNNiLbW9UNlJuYQaPuAqBn3MOK08zjWGsMMZmX892Q3jOmv
5cV0mJppC24LSVjCxz8C30LuRyjZ41XL1dBHRYF/rpE5ouXgRkc1BLqgAUImD0XX
t9d00E6YUYVPbwQlPY3enDWptMHHHeRA8k8x64oYWjUZy6vFdXI+4WscsFkmC38q
pQTD9cLgO/XLkFEhYauwZAP+EzQAJpA5VEuEeky8aFr9HSvWZ2iLjQvhYDySDA3K
JdTC6RIXIESj6qXsCbObCm/KbWYq0hfMHWrCW+wRSGVcrRG/DQUc9bctDoMjSDI1
3YP9LrcWh/yAVnL3vuCFepJFSN2wqRUJRCNUS5ikgaT+3c9McgDhLIb3o1ZKxbB9
SYOerzbgwtXCV5Ivx5IT8ww8QhQrvj1Twf/lTebhoke8XhzGX8MLry4CObUZX+Fq
88/lD6lo9Kgyd0HSDLK/bA5GdhYqapVqf0p0tlPQiTvrd8ZyaI4zUTZkVnsHsRMW
8YpGTpTXV/f5J+vP+E/eXHcqoGwRw82nrcJ214530EA7iQCHtH1jtkPervxAzhrE
+T/taaDA5cyRIYNRl/uf2iOx9Yglakue1pzGkyK4rYUeGaNoBbqmPlaS2vLQ28Q5
dad4QpyTQW5c+54KdzH2rvBZqHEU/gnE/ZM9/dgS1rK5IHXhhmBfoalxvmNfZO2i
s0RYkHhKig+NMmw0NiAbCJ1aHD5sT1GfBwAm1eSrkcgd74AkKkVZtqw1dwRpJcxI
txhVUtBcVuu8aHRzifUIy4OUSKHr6AN/1OigxMUiIV8vfzSK0nI8u0HNYyja+zdj
P8S5c26L+nTRKgbmD28vIjOtMp4IiSiKQ6zoeGp6T8c7mjOvjOApk8seQKZ7sacf
P04TK6k0USle5XEZlmUGGC+d9ccEr3u6fMDxXaseBe7v6NsMh9eCAsVy/bk1zgCj
Q4NAM3wkp0SfgFXgcXoOIQST+zfP7vq0QQXc1uV6LwM4Dlxohf5WrFWGKB+s/8SL
rRgN44ZCYDpZMgLIosrkno9qJ8I/ImLfuH2hzZrsruvpx7RtNxQiexsSRnPcOeZB
/87Qz+mBIGsxtKLoGNlRe9ZIdnxDaIzB4SOPWbEVGACKlVTWJUbnhM6xB+ApesHK
vfZykNzsLbttvpiXH6mmOTs7RFE4/E2pd2LEAebvoPiFN5/DRyLR2SIFzyUPhDuf
jt+MWFTK90oxLMoDgJj+KgywZUIXh/Iq7sBEQYelY1xLUnn07bhizuHPfK2nwEVd
W/NRISe33CXf9ZX+t++h+JVdNtpQMhQ5dxGLHYYwVWZ4zUyixjv+TWPCJo6f0yH/
ztBWP0E1lUn7dHmxBTP4QZTTyHEPJS39BKjEX/9+8oglxU4CpajvFe5PtGkToWZJ
j62D8w2DcGulWwWCaXFaPK6Q22DFJECbw87vzdtMYPlwvjuW96Yshs+nK+wQYuDn
1ixsQwsm6fJblueB27briGQRQ10HzITzjTmDbQFEBZYcosekHhgtg21g6Vm+bhpZ
AaGzR3YuBezF4cz7gwmtGwqFnHCf0+rXzyYACT37stP8qvU0Ns6W4qG39eenMHpW
M5WGBAYDhwiNeIS8RRt8v4/++khvQ6HtnCcu4SMFQ2mm4hB0R8hxKQERHZIJo/QW
bNQ4BFsSKdZWNeYHfiGB6Jp/BfqKlnPfFHmgmXxtaBsUEbGBYG5tz5c3HHcsAe50
Mf4p1HadXJuNfe7oMV5GuEupF7vAwYmbce0d42khqxDjkNuCtz1blfD8sfQRp3G3
axXNWz6v70ln8ezMuObHKRHgeEPK5/sy/otC3VWuC3qRGcNcS8WO+LiQvHfBrinw
6cbKuyKlP8zeXzNie1EM62TyvhKMYTiJHQsgg6TnHjpYjXm/KY5xwzlmgUDdQeb6
cYoHtfICcbgT4XjWXaiwtjSATmyW7kvwv88+EGeaWLW7AqKMRlWSpr5rJDpbmseM
pb2Ed2ITKHkmNWyaEN0xJDaLXv6f8tyclh6Gv2jzqTcW4Sd7prShz3NwDmKqRGDQ
kJva3xD285zNdVN7Fh1nuRXBxJM033uIHY6yVpWRU9Ev0rcEZ5rovamTZ2KV8LjM
DKsjgxtgMxkyDxjhgTYKFqlMVuCbW6C88rGXPD0O5YQVZq2UDxkPyKWLRiawgzQq
/00sJ5ItcNfq5yJoX2BqQDIff+gp4h+QhdC+Bk4K/s8+ZPRzvDBveFamrWHuFN+Q
UFAN6Sa2Moj79H9jpnvPXSwL70Utna7UWf4j80Kzfxs2HE9D3LZetE7bJLqUHfhj
dAUywZk6Fb1/Ro9JktR+vZmCws6IRMpJRV690vaD3TRVkPPYDNd1jbiRebeR/Ap7
CR9OxSDtU84XaL7y8+O2gPLWSQXf8ckDuwN0Wg+F+N62/Z2w2jwcEx7Cj97TaiOW
/lXQqOOho0kxHsfb7xswzX6+W90ImfdLa4jqP4KWJMSLPQti7tRiPpaNmXHrS+ne
5I3Pumw1gLXBEO2BrQRlDIS5SqYXhoEy6Q29Fw8f/CApC1OQ9sjivXPgmK67ixlx
d8KVfzCuvSy5Bb3ymMPKIiIXBIxS51O+8kly1MegM7efVQ03q5KUiPT8mIGKb3xd
hsl3xMxQ8enQ8MM/obfrHnks62Dgo8m/VgixHaJrG4rUuL7ixgWmCIvJZkXO/zUg
jENmB7sLI5lmcY8zvpoPRaK3hjNicyzTP5cfvceCtvsIfpK5tvA0sosQTdCuUjRm
gzSg5RspP70YJukvtCPLHUCr08S+mZw6T3V+J60W6Q+g+vmkSl3o60PuQG3L9WJ9
IDgxzcQNMr8en+/XWw4PZH5JMUUPgVirq76DndmeVtE7Eze6OVezi5THEVqE66ie
vTd7SV6vqIE0C0hU9Sy1CarWYs5ZslnJeCoGc5VXlj/XstwBJLp6nctleEYcckub
LobkrZ1j7bCUEQNuZAIMq0GFd38zqYgO4qJbBJin9KEOO/TPVeXutCjRWMqp4sF2
EgjLceTJdDWISy5yCX3NQAD3V+CZTzzHeMNtB5g6wOapShruMW0AUhxedHtAZWko
whihHdnq4Pdnp7cfgPwzQ5eLHvXwsN4qdYCI307XKDWmVp7RH9PG+TOLsi/PhLOg
5o6O0IFYAvsal9i0uk9jg+s99QfR/w1j5C26gFLBjXNrJsDowjipg0t9Swk48rPJ
dD8OXfW1Y0iAqW7u+DMfUWJE2svIPKNQyzfWJHVGxmwobDf11QBZq+H83htceVIc
APllYASiTB18YvyBlWrMMQGdRcrfbp0ctNsW1/7LrNtW7ks0zFLQAiRH+2vlVlV2
OM3Q9rMmby546NV3Y6bWXjgn2+Q9Q4lpR49uMJe/eigPUF/NEyJIQVVrMfJ2+xWp
M1iEJ7Nr6dEkRsB7/J3PUnd5DXV/KUIGVcY1VUVGmt1IFLYQhOLhY2sJ7Ln0zQAP
u/0WPfq39ZD/HwrEkYgdssVGgKQZfyX1PmNhMMbsx/gqpcg8M71BBzwO1ErLwKR2
F2DREI7/kr5lg06lZKYf1aZw1KB+KCAzGPxU5Pe1CVEGPil5D/ukMQXJ28s/tZSw
CEpoacG+JAk1KeATlbtpqhnMe8ln78tBx8IdM0rqCa4nULX2DDY4TC0svUw5bi32
5NNiOyalWgpyJ9W/g1fWY1ghz1r6Pz2NnstsGnd4Q04UD3Iaky3sNT5Zp0jlLbdm
HEpNklhVnSGCvLLyveoX/MvRdfGntrqVbOU50+MYFezsHDr3n6cbw60AihJHUZb/
UG4Yam1pr81oAXHbyhZygwevzBbV/8eUMjCaVjGgcY01UDiRNJ1l18VDI4xF3hP4
CGL97Cb0rcNC2ISqQ/kGiuCu1j3jkjwPfAm5qrox6yqkZzPgUqvOgjJn34/SANsr
fGKB55/VIW7hSuEWw6MTVTrQ34CfmKLRL6juhcmThNasG/UBBynZSBoHE42zmxyd
lu66LkeroTrH1p5jq6Rk11wdKOv3a/xIR804zbAbP1hx8YtNYGJTRsGRw88hxLYk
kcrfN+vwKdrU97A9B1v8/uOdK82erZgADL3TlGwauHD9wTkSFPLmWYJqpFRkp9Td
4taZXuNYT2u7wrEMTLdJkXyD9ZGUWqiq46VK2S2QavN2AlM64lqPuAvuRNAVV6zK
GHRVKy9lPyNAupsRL2RBLamiDSYkoFp5wGr+CTRRjQoMkA7hatItFMAJYb+sGZDZ
tUv6A2uRZz5SnXbigcFVn9wdFTwtMWBmIdk5eCZJksaPxGN5IYxWL0aGW+hglqPc
lVpJDtkThF0VbI8oiziyvmOTQwe6MkEgCy6QRNu4iM4vRYRb2gw9+oQx5QCSjPXe
zfaV25CqAAh+GqZAmZgPCGo2S3zOSEwVIaGxo4jwQNayPMeDQuVb13SvBlvmgVca
gFruLGcXAA3SHErms75fDdcmNBT3JzWyZozcz7buzOLeCZcRx1jfwyeb5GryKVwd
xTFDZPqxRfmBCmUJnZcnC2g532p9GtxegeM+HrYYzSCHGHN8ShXS/GS5n1O+AKc+
nEU+6UI46FgnrZibchUH7X7xkWrGDD5xhpjFLLWJQeI2VV5j7mhMNLCJn1lQv6q6
eGHCikHeKmkghugMf98gw5XYUYsMozUtMMj7I+J/jVewR+AJ+uiagvm7O6zcGWJJ
U0ZKCR8ho8AxMvPPRpTvpWYJRUfu9cUwjC3VPXF2QuHUIZYwqqTtppEgDGRKXSi4
dw4oNVOqjZOlc3csF8ONQ0htEP6W1DkM5i7OOFRJQW+HFqBvZpzBbN12jJxv0iZe
0zQq55sFYq1udRj+BcUrJUei1dunBBbHutuu1mgxZvqby2S2jGy20Ckl5NXRCwiO
WgeDksxWFRuy/Uuy8iuvb+ww1RbWeJHsQjJy99kJlHdtK9+O5FMy5k7R6hu9UP3E
GdtD/1qe6fkO6P8V5lWxPTNhGvI8FPiWUrTIz7fRK4T17hDKFQC9azw0Hg9AHoBH
NLn8pvGJw29lum7y++2MmjUu5ydRVa9pWSPW2O/w828wO6dISM0Dj0q1h2x0YwgE
8XHXCIyrD6AS9tZUpJ8BewjdzI4664c1LtonXuNmKazWXXF3PEbpacEJ1e9wZf2S
s83znyTs0aQqO+OQacZljLjpz9jPG/b7qQnQaPxuw5cFRLfYj3j6Os9cGAVac93H
OhaPkOQjCC0Opt9etkyi1FqmE7pR3Rg9l0eFR36PwXtYpAemPipu8mTqo7hzxw8H
xqh70XNfscoRQ7qUoWTBh8746ZYModeUz0UVWCqIAykzh1K9WXiy38VRxxpwB7HZ
ib2CaENQCZpDMyvmu+BTKZaeQhlsqRkyhOK14dSHRQwqsFXIKA7fhKDM+XSl75OL
krUQoswBHHxtSmSBrsDV3O1b+CO9jpLuWGNfamOZskVC4GNVRcTR+BaCw+F1zYiP
4TFBGQjYU70m0QmEs4G5GBXQJfw6idNgmLQKKoB8Ds0d637W4zdGGO81YMNpQB4W
ZVoAajGlLgsnrwFWnSCeLDFGg6EiCp/uSgL24MrfSMTx1VK1cszSXwjmDEjerS+k
QfJ9rNrkIM/G+NjMjwzUPJ11EkG2dYtsH/roV/mR/Ffku1f1W3OG28jOdpAYtS/N
StHT3fCIWOkkNb5U6j2Qr8e6GkXuFDqtdLLhOf3HX6gf3Y9bFZEF1AqCL2kYGDLs
3XtzcfZr9fT3Zp0otchrWTfv7fmnJUYHfSMk167vUVTyN3aLtodDrpp4QmHgE0AX
us9fQVcs9JW1sna0EY5zKHHlpDMyt3wcchNJ3X7XQRNd+ToIa47rjQNWBOWHSEQR
dephMi0IpMk5CGeieh4g4BdtDwM0mCS3ZkiCc7RQIEN/kFUksFtMtPwbMqEpdP+S
o108jXbhIRWwVWqBYV2LKYkxTne5NjEI5uYLIbpj9njEZXsjK5fjQvMcziWF98Xe
CDlfCi2Y++iAt8rzYDFRtg+XgsEvkg6ybN9oF7KUhA63Jltlpdgkq0OMNMwIwCbV
OLKWdTI2puE5cLsffqlQqzmIA87kSOcwjBEnVq765jmXyJ8WE7hHTk/vs3l5I4mM
dYPz+YOJzVA6OAlktSy3P4ZOozxcU3pr/oKEG3XEHPpC4C0XKEP7yA3L2adKKRkF
/BrnUNYsj0sx3JNNGpzX0nDH/xnS8wzMUUqL6NQmg+69/9mYCVYY8j20zK+7rT3k
5Mxiq3sj7P4z1Yze7bWItDUzqnwDX9KI0lYjdHvf++iOiVInos5BNR21NmYRnUa0
IinmHGp5MKhXPDf3BKUqo57j+BkJzJS68TIuaEdaKEdpo8naKS7qMT5ulRF/ceRW
GNncs/eI6Zt+Y0f3jK1twmT2+x/rFvRsSTRIM32ZgGg+rNZEndjGlhFDuRiJ7shu
FNB67WejbmNR6ja4ycvxP+lb7o6Tsgtu/g4L+Uu7Y5Mytj0wQs/IvMTRfFq0wDe3
8wfb8TWQTnaSk7kNz/1eet3Y4OBHkbBKKAxopZ2YThDl58sQJSs1N/iDWQ7Z1bg+
fhj3uWo8sOEAWOyVGYvpFMh2aowAOmr9uyen7BAhWLnzSvo57fjL1OxYWspUgYgC
C7w9gxyA/GhRjas7ZUbXYxwYJWeVQhrnIrBXQG3OXON3nw0s9fukxeMYUbHQ3/Qd
hYtOXnSDLiBAB+MN9i7bS4GAMufMa5rPzvug+0qVyjnFIT88A2RZL1ls9ZSC09jm
a7BJhv0MOQzLR2aZsVJbPyo9tVIffjD0tVj/lUWKSwrh3cQLr8KV+pkcMWryBMf8
hh55highWcDGkwqCBvbbCac+ppmrjbWeGCOHCAaQBLyiy2IjeE5Ro8PoEUxmyrO6
KeWlVkG3woGD4zZKDw/J41AAIKdRoNKQQHFSUB7XDqBxEAv2KYEg02d+X/vGhrJ3
/CJ04h511XbbDYWiqbI7OMY4VzqwOKcZL54taLLS3Hp0Db4QfPVanDALaX28ARtY
htIyOoyAA4y3kLqhhjcU1syX12MQKWtXAtVelAgYX1y/OFooMOOCDKkSnky8axZm
PAJIakKrhgcOA4C2z1FBWIRWi+hFOVKLHHiXKUZVtiR43gfL2xC/2xxfY4vVVhGd
Che659NDPRWGUDIDoal9+6mTVehrg87Ku+vjlnSneIJViRl2Bu7S2sjMz37P7BbU
cY3EYApqeZwxxFgzgVcfFkFpCoX6I3nr+Pb4udWlEUbO2FRTW6DRtLxnsl8WwRgG
myydUC9Ufvc1tnO7fY5c4peGVQx1A9NVsfIczBAXBZyPc1MWOPdNXsLYkQMNWCaA
UfKlSViUyaxCovvvyndz7EwKrgBLfTCthmpqvfC2hxQ5OmAe6g2gWxbLMYRXOvVV
N/NQimFfOBKpD7XAaNCincrU/lR4VvhZQz82s8n00fffAQX5fr1kMF6hr8N6GC0A
4W8ri3cxuGtkO49Hu+Gmmr47lOiV/2DzOMW25d9RtH9kEGAkjxi0nm0JS0XASXYh
cz0qUMVoV2qJxCWr+9yjqNOWRDVKmU+MV2zJG5A187quiOjac4E+Q9DDMhRbAu70
aQeDMlwJp+S/8mMSnGFTVx4Cxk/JiWJuKS1b3TZQKm1luUqAFSAIkukYgIB5wnrX
zZzIroZPKWAnXlp9bxS+Q/H+w4fwz7C3NRYAN0IsMj3ajeGSSLDndT6hPL58aJHx
iDExURzCBE0XHWzFFJyU0tQ1x3IdvverUUiwyJewAWv7pXUQjzqqObJlb7J2aJJM
haEqY2/a5k/b4+wKkn5aze8KnOi4/uOKPc67HNPoD/LXW68/LEV7SOc6n54Yy0ui
5oXu99UPodUHgMHJxel7fqDJDwi9M9+XKCD8apalKY/F/M5yPwqtHo9/5AxE1LQZ
BI4CuTiDgct4M2Ad7A7u62l2IAYA95vrLA7MQL6xD3sroevAOCfscPYtJt24Zi67
cVTqpaUHtHhndX/h3XIIJzbi7MhEPoxcvKuHiv4kLdzuFgBL0GCFxXCzcaP+Vtn1
+eOZ5p7mppiT0kCJrST3fm1swmz7d35MJB7yS1zqSdY+MVlVf78rAJo8Hx1eZgxi
eg6PGrXwe+hwuM3gHI1+tPSTnX/lNnvWLB++NXOpNKRWEhS0mPdwZPE6L/JaUgSI
1eVpa6pg20CCE6vAtYPwiDk9C3O2g/Ydr40pKqMSWrTM4aPS2M4/cIz829VACtmm
igIc7ZHVIBSAsbW92q11+v/JMmznEVKo5Ch10Por4lEFry+mS33KSwWyqkGp9NPs
ZUJ9jeaYTZMKNHLC6JCTXm35fCppXsDDShjIUuhts9NF2+/U13QJN4pYtX1aSz9t
QFnTR6/Ev4EebZMVqfnkb9t27kSAXW/777BVw2jFIrGmf6z8jkQqBQ6l4bffbX1/
wl4DkRfQ5YmHOjluqv8JGfO8QUctS3HEHGjqFTyETKZR4VYYl51E3FjGWjGiimsd
/iVB2jlHWZPpAnIfAF4Ret4yWppBLAau3/twpKeWGw9TneD7HKOyll2q1MmFVpi2
+cde1jYuU7YDKRPl8KSpSFYdSMtvhi1p6iO2740Y4S5Zkfqbn1EXOZi1hXbDyeno
1wPhhrGDbE8wqo+aBCpLFnmI9f1OVPMNoJ3auBBUUqAUIT029/S3oQXabM718uBN
9V4Bc/jNfurqx3StDUlj6d+YqQWO9vZQETpeQWqB73naEtin5XJG2mmHq4syuKT9
nMD9F1zqbTh05RCnhd2LIWoQASMQCniUIFyNP0m/kH1h+jl6ZxAmI35cpJMOPpeO
ELCUVGcZzrLjQ5YGYU4a9KMmuclk7DRu1xAF4fahMB1xL5QQc5ILEMoWdu0zjrpq
Hg6WXfdAruwk1rekwypFpNenr/Hw8D6h6AdNqgRCSXG7tSXNHym7iCbh0mSxsjvt
sJUqk9P24UzWhexZ/xILpnBsAD+o+onjyXu/D7yvAYjFS+XlCOXBU6FJ6kH8IRQX
6w89WO4KHaOcS1q+OdTEL3tSol5EcP4TpoZXNpO/h/HRwY+E5v/l0IUKA1ClgUBl
1cm5G0yp098IfeAPtTN4urrTCTEkLc6ohYZImLID25MuenLeSRCJfrZ6qXzKDQth
kNDeEVgJczmMftAdgHDMbO5EdMhAGrX027Zs7WtEibxaQn4nX6MnWa1yIohvCM0h
eHM+cQomELcd2TIvobg1fDDSauib3PTd4f3v895OJD/URo/lewXqZmH6Aqb4t9qg
f5EL67Qhbzv59aF+hau4T+498vl4nX349tMzJN98c74YMZmCRnFKTO2cdKc6rrnE
RRm3IvBTujgIjk5E8mWHw1bsnx1HQ1Gs1ApERF/CqaOcCCrpI3KhyRfgF9udeuj/
tF0n0PlhttiAHh4j0+j4/ZwkAjcyQBC1vsEmOMOGcmT4De7bvsyXWTVt0JEsgufP
1bZE0Ctkm5MEUyBRr0x98vQA/Tk/NdeEBhWH8uUSWeQDZLnId8TipLAc3hcOpGvU
C8mDVYtiIhqqYC6HUi2d32C8oL7fRseFjEM2UyTXnjT5LTGZnX8DFLB+OGch4GYT
oO+sUPmAh24W9doaD9aY4M5ciMiUrHL1k8vBn76jYwgo8sg8kH+MUYiB0qHorHwf
xkP7/Ayb4UdL4Kw7lzTTJ65QC4n7TV2jcYJxbDq7gFBMLEYCzdJaTAg98WzakEjo
xLUI0H5hb2TWCWYJJZOjO/D7ppn+NFTnN4/FXTwT0XbUTc/NGaAi7NEj6qgAQ3Hy
kdMGsjW6OAuy/gxpb6LIH7I0AAXneUhu0Ji1XG9wgBdAXcr4awMSvNEbs88wC1BM
scm8FB2VFk8oDytgtwx4MXLORDXSMAcfOokKD9KWa0D5dSTw6RN55aBXvnRJcKdg
9aLE8cbB6fNTYXEzA8Fn7OjYEWuJXtH5qRvG7IjcWkYFHW1xi1dWOuvlEpgrec4P
Y74yOCpB+sB3+Z55qaWaObCx5bO5d4ObKnO6oRzcyr29D1BLUbRB9b1buXQMbRd5
aiIXNGiW2BHUcv+tAz1iiO+jvv0xE7AJMqFyirpuoSxVVdhqmSUMJtvfb0Hly53U
Aw/KyJpYBy7ddqISxZsKI9q585jBeXaK+Gkjb+TSeKiIQ/tF5mwkCEmM6MXQnMfi
B8cidTMcKvBfKwsal6Mt0uMCaD9HGd+Cyv2hrZVD4fp8QLZBDO3UYwzmHjCyJH0s
/LIq61a4SOEUXyXyoPvfavM/6Z01TAHrh+bIIB/rSSLzHwNAIBvKb6ZL8vNURJ7e
TB+HisyHXmrueMWjvrIsYZjIdMwctG9oWDdaRtu2KvDa0ZiZu0ToBnq5bax0ctNx
cEb8BT3y0sUnHCrIFAjIURz0dyev5OcfgInDZ/VNbowQdQamZ7thuKsit5zgCtQV
xv2UZTDetYf+9hteL5QU+0W0SRsRghoNygdLdUbk7wa0m7q1P4YiNQ/7AEVrOCBS
jbuLiSqlUSgNHTfWbja471CbVegcqEQXkmVSpQe4OpnYNZNgz4qWJYMhfQv/peWC
g2+c6rcyrtsTAmv7OSod5zn19xLpn01cRB3XNT0gVkQXw/K8VV7/yg5xS+rPi8he
b4EV4rQHtqqcO36zxAOT2q8Xf/VsNSsawbXE3w5fspqYz4SNUDeXcUsvPSXGS1cl
V77ECnrP7dGQSLCYIWAc13ZS4MRt3zJlIYY5Y/jNGM/K6qMQT05vnLPAhNTjq9SS
tb/1DqWIIf+7kGWBs/BIgUEdrUzvGXN1DAkxklcyzFS21iw22cj+GqLhHLPOE3q0
qTcliJ4GpXJmJJImpOWNDO/qRBwK1hPziSTrg08HurhqSAH5SwdX/A4XUheoUAqw
USVJncnlLvtAXkgjHv4EJ5S+gaBEVWE0QNNy2q1nw4/Cp7VArS7/OEC7rHa3UBx5
nQYizZ0TkWvCB2U+ii7O+k7ekPDMiJ/0maCcO7qal3IG05cetABz0FuV2dqJNDx4
Q9tryYiceSPLMJ2C+ujIpiIrLqx3bYWjACdhSDKOiz/oH+DZmKdb/gLT9l2iE7vv
qZ3A6fFGOBxUcRooWVk5xLVFqouCRh0oik4HjleeXTO8I6yI30Q1t8NvoitQuaBq
sOgMCRHJdTS8LKyM/Hxzv1OBYINHATDFKG5TyQXBxddtqiX6Xtsc3TTDjQxwahNU
2OwEXm1M7w3hTESYcsvVb9fDwETFnhDutg9TtEuFhDIIkB6el3osB+w+tF76y/0A
6iMrft+SE33kKvn5CL9X+s3El9rEZb8DVftZCG4SM6hcAA+3R9j5oAhm+ilHuXya
YMnc0Xr/D+8ecz9LMfDxG9c/MSXeaKduYqV0lGzT2aaAJkfYWTrK7AI8Mzg86v6a
c37eJisj1CNAex0FHuQkv6Z4Tewam9gTOOVFj2TSxU13X3d0kX/w+e6oKNfp3MWg
QBj8QQNgamhjy8xi/F0KqKA/bgcaKOtFnVBXxOvT+rD9bBLwyCWXosbOTSlJ15MN
H0ZQoV1O1l8uP0FqYtg8gLoTRDucGEWw0nGElXQPgpHPVdNMGTgn0ePNLk7l85Vp
2Udo7r7L21u1vSMnUa9+s8w+wulFhc818rOw37TCA06Mv97TkPFK3OJNGdvqixDL
gCp+VUp0sVu7N+ONCOencgHI51vd0rXX20+MC1MrcvGl1k+Bo9mMZwIsWqL/T+nG
un7B1Pqb+hrZHmc6qZYyriY4q4BVthcrMbf/Uhw9gbkKdEeNonFonWrrIOz+hfSF
5juf4Ew9yFPoCii5MIhgoOHh76FRUBOq3oM5vMPSWJkp0F8CZ0ZOn9225JXl3+yM
pfcYPdMBpzA71uRZHzZirHuyXb8+mwG7hzXVgFdXAbp986vPk997j5hf8Fw4Yocs
0WJQN+UFOPhskqqM2yWeEV2MCXX3jxOHsYbTcel1nDYZ6VwSMaCwJWRaR15fvDto
ssKeeXH8R7S6wEE02Mvk+TTFr3tpWdHPayeGWHbh1e0SfJ0I/St4zdTt/SoazB6P
KEujv0xTOfqE0hv9NtIu4njz2jeu9WjLLYnsyg8zJXhzAbRcs7Hw2sv+GDfpzBCz
LtRTAT2yPGkM21GVOKwlNkMI92vlWHUdiUyvQkqkVVMNAGoFtuNC+E2bStqrW5cP
9lkYGfbsmdovWEQGlukWhp1vl+IArK3mxKNMmdzi2Z3gpFDhjf9XWbspqaCbNjOk
aZAYHfQ8e9UJBQvadn6s2I7MKMJorulgqfcU1MtkPTpptBeXvDFo/14QDN8R9M+8
THiq+w2KSteAOOgBQKhvgdHwGxiWmhluBSABdg1cuKnWW1n6j4TuZ1zLeUWm0+8Q
FmR8trOPeqUPvVty0DsEAcZOUCzYGrqJJyWJVEj1OCivy7tV6oYT77eEB1ExbePH
y63XMotUeWmNXOjkED7sxCqhxIXJSm5aXJCGQeIBt3biyN9+CePuf4aWttbHyLGI
nK1a6Rfat6xNPfgaNbbdP03xSSPUNHylpgYzcQLMZQNeaBFr6ixcWx8kdETRxAiu
NUX8AR2dl6CBK8oDDr0WwcvGvnaX97JfbJyNSi05DYVjSFsIhjqFBuLFU/7VbISL
TP0GXz97SZhR2bma8KQ/ar92Ni3C0CNHnNWtZGfBMPpaeE4ywxi5IVDGY8sEhEJ2
QnAYrSFVhefIeCqPj/xyXOG4y1NUxs+Qe6eyu8o/v8c+Up5zOUU1oqjOKwp4qM/l
TonPH0xrQWbw5epZHjEEzEDnAb+2Zu+ilBTlbvfwMOCFKVccWVd4kMeLn0VuKCR+
KkoTFa9Rhcb6YZg0oIQhx+diZkj4cTR1dBMEU+M5Kpb2zn7KWyOtbi16VC1x7JVE
+3Vz/42Knao2glIJQOQqp0DphSpc9wpO1peWPyq3BtFk3wyCEpH0E3TwduA67HK+
TXhHgAO4fAblSxTVlBu6oLP8srMy3v5va4hdvFLdjxkyfMm11yhpAgXjYoxlEcnO
GV/d2B+aqUHnOMd+DPgIXCAIUgigNmW9JdRHtrXmxciadj5bHrgWxSbIYF27VU/q
vfCtSEQvCBzC6paP/l6fSN8tUDPYiwEBYnaenHCasYJkUE2fuUGPCho7nvyXm5pS
ym1Lee/jIj4Zrmm1rChDyRg5IxlLNmiO0laVibRVeGrxtq1s7g2tgIldc3yZ8bX6
6kyW4rOr3dy3o57SjDcTS06V0wRApRNd0joGKs54SfI3L+0Izw6HckLz/LWnyXVZ
eVV3dPpRjv7SanvzozBTrejPefwEUQ0p5CwKwCrUoJPAHhRK8MEH8u22DqE5pxk6
bvsbKZWTOpSUeZoCSOhaKq65HNNDXP7Z/P5JifWEdW8QyGr3KmNPoCV8lBqR9TCE
z9zmBw+tyD8NJuzCIFGHtbJmFqe+YhtOX0Nwcc4KSUGhopksSVhQlECKPHd/2ZG7
dML9VGs4nldMe+E2n8g01k29voGYrIqWtNmiM9FAONDEf7PpODQoqLn1lvdUFpw2
/xXYOCwDFc/hvrxh8DCfhdbdIS9kQhcSNyJSN9YZ5YQ9WMedlr2gbxIs6FWijHJN
Pc9JIYpOPTqzxNcXiWEzSus7YN082TylDZupXYFGNd6+YDmXFe0sZP8cAbcMqqjK
GFMFgHnSffS7fHvOTybTeUK8+2TRU44xjKJeSBWT7qA2Eh7dGU6a+UoT9iBuaJhH
ZW39039Fbsw7W+TqcXUJmBTaynWidJDS/I4Hg83RLXjwue9O80Vx9tb9RWNLaXXw
MT2c6hZ43Lj3fn0GR2qoXQT1U3aOC7ieNumlO9Zs9FcJ/YA3dMp7iepyMLdoxacn
c33b//g+eGZKOJ7IWWXDez3DuviDCvvjoejsRu9e5My+gaQOeb0Q3q1MamlqBTOt
q7JCP+zBfKE8hCW0pss1sweJJ62kQMCL7ds7rMrsHqMFi0CC6sDTgI/iSmbE5CZG
mA5JwBv77I/38OpjQ/z6vvsZ/yi64gNETaA1Ao+GATPpcvAZpNC9bPyiQbweWFlA
fqyKjPFvIj+L9IqfNrSHaXiHQZWJO3qS/6SM4C/kPfe6+hH05VWDAvtVhE6Cn6iR
ZVORjCaba97hR/480SSasLCBzBRI2aYJiZ/1YVqmfvysr+mqpoPjGCHQSIJCb7PH
jct3Yp+eUqVQJnSddn/OCTaHklstw67abSZp0qZQdGtyacZkL5ZniZNJpCHe8voh
r9JtwTPQq1PSHtGIUTPjOTl+wzc37aWtab+mWKcPd81s/lOYBihQk1ZFI3s915vT
uF1QCVtSSCTKCvNkIdqO3VRyIzC2MBLCvdaq2ibIESzCDV3N5xWLRJSIo06WDhx6
bpSWcxC8JJiHGtX5D0DX0Tn419WxIRsVjjRGruiPJPEDmwJjSA2RiPIegJZuz5wU
qC+W9GWaFfOCGpJDoqdB7sRupEA/hW+kGtmvymS6vJBV7aV92ow7YLluX1H9fym6
KdLdU78LXG4Eyx7xg7maIylmWQyjTY667eH3w8d+hI9ptB6htvAOr9cGcfjiPQas
xLbjn0ieZOyzKwWGVafSkMIfo0N6qRA3VbbXcZ3XRQALWNIUG/8KtvJzNNHuvDAE
GpLtwEpKiEm9Ec0GQzh3PEe28UT2UzkyyRqusS+fibw6t9hH2ZGMIFSjg8xVu2TW
SG1MKjM2mhQb4e6STS7Url2QsdY5pejO4zSdVJKArjzguc5MW1MO/Sm5qkDpMwtJ
+/SDzGY9LCXZf/7DDEkzcfQl+z6PxACzOoYdM5Eg6l8l37TiPPzRP02nKr5zgZ2y
0VG1L9qBOGCTgyivpkXp9mMvdPsViISxf6QjQv/4bsw4XU1ooL349vwcmymFrqxp
t9ynuAfpsYVaTCtnN42tqV03IM/U5ZjU6SSWtmi+mtZ0hPcW5+ssHdYwO0Ss5qW/
6N9ROjH2AjcoBZ9rB4yrorC7rUszch/KT78uJX67eLPgSAfxq9xjYFv9MU4QQJTw
JRFOLPaIOHfSASob1a15tXVFva+GgmQpkGC3X5/i0QxYSQlGiQh4NJsaqITtesKN
a6dtld9iuiCSMV6NiNVdzwTxzCQNAwVSczNuZOeYpwvBAjn6aPYtDafVBKCRqOkl
o4DQA4q8LANNHiEVGBZcZ1jhqFxu6TFkZIaIXpsyt2gg66xxfU0tb27Yq70asrpt
tbdAxAbSP88yr4ReY3VKs6WQqgr74aJnFqmqHKPcNuePXss9ptjmlOgQUhJ5hPg9
sC56fVZsc18urQV6vF66zg/FJoCpxNSyUeHSL4rHuZIna0QE3oO6d3zsdE9m4YXO
x8cjx027ZpTQmOElkrIPLxh+ToKwQlE2t/UkEIqb+1hFPBRCLQ851ZqXS6l1eN8w
O7tIHUajHQkUrPaN3sy4Vo9fHqCvx5HA3UNMaCERSZp0jLkWD3zJr6M58Srg4Wfg
ssu/YtPIHhNX1YBxL4fisBKoo0vQVwu7HKhZaTul/Iikq5qJp9/Et65gu/05GH0v
uGD+OLa0AnSsQc67IJMWYM+l1AI327hvDBIuwD92SakXewCy5cpdI3XdV8NMP8t7
NF6lvtOkgoTc8P1SiAIYDRf0xH9MANnI99tWkcADcN1pTN/2E+DSqjc3YrqW37Kl
UHoCuP/UEIPRtTIZ55tZjsadDFRm6lhPZm2eGcprhYENH+BbJRHM9NadWb1h/VqX
Md8cbBkIIBuWCHziyfyM1pDPaiF4mq9BZhJZBwIC1gwSWIw/XeRiZI05zq77P0L2
e0+a1K3R6hBaqCjRSiG04gg7/QhmGcCxR2f2O56SOtKNy5CH5lzxUKswwzK2VDWu
hQE9G8bhPlu4B+n/3f3A1/bCcZcaAQFqgGq+SVvKd6LogMehdW2mJC6q95eA8jMu
U+WYG7b+dt+HuQmPSlu4ZBwKVg19ZQ2Q7d2jtvLyDP8KUyO/CIFHFLTf1ImZc2Ee
N+3ijUPnePq7ak2gSUVbdH+BSf6usT4WouUyclFaDC8Ur9OoaZ3i3csAMFOV6Th2
6FtgDXGi8QAlTEZYoxQa6t0J7RKt6qIC3x6iyqfz6ool3hYgBGA3+KCJkloOxDQw
MIu2SW75K/gxKxACwF3JJLXHvfv2iEKoiC2NUAPxTPe7LDWDiUEbxLWLC/b8Otnt
/MSqgomna29n5IBxWmEXeLQzSaJlCUzhJKM2t31t59RzwHN8x3HrMKqAzCoex6fA
bPfTzTXGWU/q6Fgu204T6d9B457fRhNLbfKhIYvyC49glNvt1zHmu40SXrEO4UfX
SCbkvZZsZp+VvcqptW1uDgAGcp8cb8e1hW+zqkDarLBQYIz8r5tsWzJSLglFAK8X
vppR6lg4ToIBLedBfZPxheD5hBbC0Sof0BoB1MtCsdvk4rYMynS0KttEbz22vrNv
1LeCuHemFYE+GNDoFzMGbeP16OEdSdq1LS8n12u9b8OBkQypYUp64sB1+RRpvk0P
i/4SSXDGa5yrt9yMEK2vZXI9wHcIOqLf8988fBxoDvAftNiHgsV2AnvzkR+pV/r0
ToCthhKu7epQpMlVakzVe5+zMvL99zJY2l5HLDwT1y5a9QznFD9xhC5KVAEXtxz0
CsPy9eNeXK3VPHEyNR981l2Idx+GygMTFY4Smg4z7ldC4JImpckMi29FuW6utHeH
gFksAeCJtk0IDWspdfEie951PVGihVGS63SoriWOe0BTsJ3n3JaNmDMi+HBLcva0
KqrMn4vcDigLai9Mdm29uqvFOhVbOC9cosHWppLz2Sy2GdqzkC7ANuAbzv6m1jTT
kxIieNl7mFYI1bvbtrGXX7OO9JYFb45CKk6rmrH83BTg55xM3dACgvM5DBuzjpCC
cwTvGAjiPPTfsFVIZ/sgvdLwXBvPNp7nmPvjoFQqIIkrL+Eb4hZfzG3Lu3wJY6o9
kAcNhykhlR2etWUtSVkDqnRZ83h9fFZJ9Z1oXHePSrGLssmJbA1lTtAg3Ny0tLC0
X+mo6D5lRwhtPiDDET89FRVSSooFeDGuApx+vF/SxfrNlgzdAz4eY88PRw6JHUhC
Nh/XQJ/EM1NYQy6tn5E5vqiXqg8D7wXe/daOaAjOcnEO1b0dTwNErThKMUNSspPR
ntcg6JIgiH23xCR8a3nH3l/u9mXRTKUz8CGm+LA4FDaY5O5j2QUYgEqr44Lhj+VV
PG6ZfnhcIROPHsL0PTzgvUwm8EAyZV8hfn+PT2a7FMb0E/K2bQ/veEeA3qck+qnC
tXUcW4b0+H9zm+7IX/T0r/L0m/j5hVQ8SGpbZfX/KwQBmVNzEILKcuoEqPmi580/
DkSH8nmcbWxr7FeMZhfjAzIAdwJZJc4oTYZtjmp2gJI9UrRkrLAbLfn29a9sb5gi
KSoxzVcrkSEWgdhT7I8rU7CH0PdU8pZnHsrI0AlnID05VG0jHLLD3fgZbxNv1jUI
DZci4y23K1Qza5qqnxlNCcQDk7Mv40pu5j9S0COpcxz3UGal3C4WAbU5PPfdKCnF
6agzVQYKGmRBz7HO55c1OlkCiHWrOKWiCrQTeH6LWarfiyKNsjZGhpiCCGCFyC4j
s+/XxiK5ZcpVr3fOIPAyVadyzf/u3SpAPAJNR8Fe0EGVna5F1F8UxAMxRg0l3HMO
atSBYoNSJmlYFUPJYbcUws7LZ4cwz11TWvcfw99N5gd8xBex2j/d/z7Kj3wE0tW2
K3pKxbLX4mER8QpDuZDssWnXZrtgn1vZQLDuq4DMutPX7teeDTG2yZ3jsecHbTjg
OGnhPUXAjCI3d0izlViZZ2uu0tAQa01Y8dLQujmacW6FVVsFiQqv+otqXzMhSDWQ
64mG7HqJPN5ERU/jMHMQjEpBGNpEb3HB2VfKDG1M8xD4pWeoyTaF7xKKdkjuOahv
8dXYzkZHO1jnCeU1mqM9znyW+hTLTQqlaiuoK8RGfSUspCYlC8Jk8xO617PMWXVu
IXxLKR8ivS1u1zcsqrzIZTG25o6APfP8OIV7Dp84dwF3YUJqP29kg3Q3rUBmA+Z8
5bXXMn6Dhw55B3JSZJ3uRXYYdI8PEwMFIu7qlBBstH+zg0oQWvPgFe1AIv0tPRff
DDXmoNgDAD/k4GEGzZnsyEayeMgM5jbO4UbNDj6bhToyAqkPAOW4BE/71bK5Z348
tDPSqSJQLBnxwA6Zuw6wtEOQPrboM9ve/GfmF3TvVz7ImHp6L+mnSv2Mx+OJx0qK
YvWmN3O9mbnqe/8CaArAL67U1Yl9dPEmOoxZgXXSS1KQ+x6NxjfHhC2dVRu62FOY
aCNzAJFWtSnKo8MFVKBcfGuvCGUW6wrzuy8sIAZw129hQ6CMQhDRy+F+XeVwcZLL
GZJbwHIWulHbr4M9WBbHQY+ESGIgh/ge3j3htB0+L4+YH149yXgukmO0MX/JQLLs
UsO+5czdATWu6Kh2H8afvFaRg5mtgMBH4+Zda9hukGdbpNK+ciuilNH2W/jXh7Wu
pKXK0u3IgNM92VLNkJKT/XNmc06iqyO06OnVqiDPpuK6y6sXsp8KJkMOWjD7fCC3
oRevs/VDIrra7EC+Yfg7MBiYFXnNwv5CSk19ffTUAoCs1BvaSILKQqhlZt50EsCF
pB6hiRQ+Xu1Awq0sTbYEn4R3hXHQXMUDIMAUYcHsBOFT4iwvFpdCB3a5hJPhDPLL
dtyiv5fJYw7HJdKYQ62ceds9W7R4Q2X6o7/N6j4sx659ZgRbzgH/Y3PldBqIJgIy
MES0D4eDcX857r4iYRBovi6lBSNMAFtStbZCFF2LTA6pqoCwpB6lYr3o5ac5GquK
3yIFW8GVNsJ2R0Hme7ub1xTBDQH+rzVBCSaYjQtqFRTHOwn69OB+hJ5lBLFQzM49
pn2tJy2bANa6LxPQyAH0Loh3Tpe5UH7/B2JK7S+LONr3BSmiE8nVCuPEEZNDGW9M
mABWAqyQ1dOwL8enhMhSg7lrbQRPEwN4Ra/koBtBU2Iwl+IUIWQ0QlUD2DlYujIi
uIs29/0wA+zgqNlzZeoEMayShmQBaQkHS7D5PHCRrsTCxZ71Z48u3/GMxjhMjoN2
WJvX7GmlvAAWJuKMENWz8NUH4OZ61JvDqueYijesoCbwpm8BCqDCkLlUTGrmLDkD
3luTyVEDOFgmFyjLwXMlFED3zII8T6D7pOGuvcTtOUfaeu2VUpSOw2TxEJgmJPmY
vFqgJolU/bL5fmr+mKL2BRD9h43qGLA3yv+Mx/1FMOznL7n1Wb6Wega12/nJfVnV
YJUc5SDYrDBBFJY09lqrtvhB1XWYLk1Ujg1T9OyHPCfKp4bb99JGkeYWF/eTDZgw
CdO6IvV6IC0iiJl0E/2UGkgfFmGJfTHaMNMX8BIhTi7Tbrs2tyniiHuqdlp2i5EX
t1SQV2+y+kB0Wbo499Ytjv/Ht69wv20vsMOGWx+xoiyLzQ4C7VP3MtNEi4UiDEZr
OWieiGvmVpemschXZuGKqvmIdEQJJdf/AIPwG3QKppEwGR6JiTmT7mp9E7X5YZLd
qIf8zOEJTqBRdISdwXfmhFGG742zWfAvYaW8EQ7LKQOhnCBAsUR189LiiFxh2LLW
x5faslNWD4bVq+SPZlp1C/K2BNFk63g/09S857DHayEOItGWPX+oP9GZWehDmaXd
GYju6IT9cNQIUn3pilmMBQHYHyu7hvPMA0rBGUkGltr46eLMDiiFx6bFjaT9nW+n
5CaeNTq80gzIMGraAyjA6kFsRkpNlX7pcwAB1Ee+Uas6vY6aNhphgSev5OD7F/Ek
UMDq0JaYcLjPbzicy5PT1Zsb1zSe8rKGOWM+4ASjj3dQtYq9ubA3kza0m6u6xL6X
eIYvxTAbnomT1A8uYwvoxOCh8rjT5AMaIZSaxePoDKPmQ4Qzm2j7fr3n/9A39HYR
1UuQ+ukME9NhbrsxkproJzZfdcL2SLr2r0XgayCmpiWA2bhMHBYVe8s+S9toUYvu
ElE2deN4k90a/xR+pPdKaUsfDUIfn3q3opLFiojwJhe1Ev1x87Yp9cp41ZR6gc2q
KLToBswGTP9AaMzI3U+CRCcglczalTfIb4AvEa7l+CqTEEXklJo1h4YhauhBTfBW
1TQ1nzywk4kqzbzlM4xzKCcBhTcrvW2kbXPhWDUHwQcovIdlQBUyzeaaySUVhZsU
PUZq0CwtZ9mRI0cRRPdnsdhlZXC5komdmIGfvosxbF9tWAMPBPd824FYSVt/jhKs
v8mmivBJf0qhD6nWMgqU5Kt4IL28IU9+JoMjy/UIOsMOV1i3xHpr/uMcSzFJoPKF
EyC7/861gzGYCEVt3Npo+5yJXVreuvdCQ4wN49JNogh1/dLiu3M64M2Tu2hVwbIN
0KdXxazgumdHw7EDfDGvmxgjpK/kQ/304lkY4F6MAh4He1T+HfZU08tkNC9Kk9W4
xmde3n7hG7giEt1q0ALjZGjoom/p2WKwxxjN1sBSYGK5TIrJL7RyLMpxDxs+jhjO
Ljab5cC/t2vOYKLvuo7EYAsRALeuHp7HSfoXCmdhQLm4YdQZv4efGjLaFuCiN+dW
2XpJGQLURgJL/eh5X1tmdLuQCmUD6FsD/5WLr+mVfzReX3izRGcFVfC+2SbUnebW
mDZ+qxSU9AmQ8SCZnRoVbnb2MUu7iS+BCGlG/IcPMeNkROY2Uxe7gC6f5db6Te7o
kEy2AEeK4IfSrLl5PxB9F8nrMYQMhEw6j8e3ZY74cv3F2+ArB/QzstHnFIlm4gMC
8wk/8qCPqhBjtFDuOUEYqmbhsC63eoajL/dWx6s6iN7wobKkv0LaB4qjOSyemCtv
7cN5I0YQZv869yuvD+F2mi9No3mrWfeB3kInCTaXhE2wz0H6X+yE6hRYjfkWIWQa
i+GWNpLLehZesP8ITY5/SU6eRYEHLZzum/IntDXjCTJ9ZvXZjNfUzZ2EBpL/RFkp
7I8gYEx9Kz56xnNaaU2tMjl+Qpu9cmg3TaBJZ7Ofiel0AAWtsk6lI4F9zq6+juE6
6sMYWllh+NWyW7wVh82imf7iZDUiB5MWhoYvna+SCO1mYc95P28ppKMNl9TxoGwt
DXl53+Mjw+D8qGeiaIQoRVI56WnFzKwJtiUUQ5VDKXl/lCFpfMamcvPCbgtWdKra
LiEETayMcJ5IaoSKwMRs9YCNoUQO7ZDU/7SOusgC7BZORGi4kSlJ9VnMZX4g+VmX
nzBc77gI5ATKmgD5/NCl1/hFgQVo1r5orpXv7i7b0YTvbCXJJrqIp9NF2SfHAae4
NdUuwPeZLt+LThQ6TzqwfHF8Iy2dY2Z7vmU08GkifsKKLtxyAvZfEDHnO//GgLRO
hDVsQcZeY2xfO0hi0sKAyY9j2PFWCik+JnYILfnMQohoT8YUcYEdKep2d2PrrQBI
MZjV+kNWIIbUOWGhw6DGypSEebZqHiHhcqivNpRdrRGtiVTc9nsNsd6/1UUomZew
9Npo+4+i3ZE7Cxm1dVCReKRzHn6oXw3fAUvP0QNO8HoOeEyKGI8Dupa2yvhv95UQ
PBkmfwKNTbzTf0tIbn1ZG5VH27obbBHG9oYySEf+dT7bYVoY6vQPOcfNW8wncdkY
ZlFjFf0tgbwstPXQEdzE/Bjw2ir2zepxobD+WMfyFlcagasmSMprC/zDYazvE//p
YCszW0lcRdD/rXy8TWwBdrANVKVlIj/DfPiaLhpwkFWV6xCVNd0O0dsvVhJbxjUV
Bj1ZZgBgLWZ0huCmquaukcycFnSMo9I7vLzIPASd+ZpweC1txlwG4e6YgXw10T25
/FU/eGL+7z/DmPMWfBE4aBqpPIuCPfJkUPgneOLl4koXychN9PuK01A1jDDj5bIq
PuL9qAnZr+8YYWrhuzZ6L9dkmzOV8tUjVh9RnQbgfVPaLq+LZFBeVUCn2pY+LV1t
9CSSQTwQMNFAdYxNGBxMd39gtfUCV7rNM3O/GjkAiPVTQcrevXupg5sM1MwmKyyN
ehB6nx2h1F9D5CsJXucHG9Ag4TKt9i9tyfJ9Ph7B9Y1lYWgnRaWQiVgJ4pNhAZK7
T1aRSgHRTrWT2EteZ2zoZB27+VooeQ1wilvwWq8gfP+i1c/2bWZ+hG5Fai+ui18e
1ujUU9A8kBYaH1ambakQEQnVbD5ubbs6Hcw8w266R+9zxZ/AaJefO7f1Oxxiepqq
x6J9cy0NB9f0lKBTV5wa9hR5DCquiEENYlrFSL4bap30LWzS5fzEL6y3cV0vVokS
n7VjDNF67HKZFB0NkhdfsWMwBaZFdPxMiQO18rAumXxvZ3PgoKK5modk+T+y7flf
TiTynnmQuSMZpDmTPfWI014y/6eLwlwEAl30HeWeZEtj12PkFLWeGJteK7/wYAn4
b/1NXv0b/swLL5lPFzJllc8vTNSbAHdy4NuXsAz7kmY57cqFZGsrvpZ2IwTpynV3
h/XOSTi5AI9/1viv+jDZd2R2P/LfvPNLSJlEkWNQE+IX3ZpTzymcRF4dkyvmpk/J
rByqIChlVfMNKoNws/mycPq+TK70N68bhpBoUpppCAFLeKTGu0sF7byGWm9N4lRU
FNca/6cMpX87QjwqqRpn1b047/z/aZnaw9LnyhK/2PpBj6tPWMpIG5eTtRR8m+Q0
kWnTqOl584YZ+oUrBi2YXk7Kv5f8jzw/hEIyiAexJ3ZeeyXH9uxJjfgIw6B+bW63
vLGWaxyhNRw2rfnkud8SrDB9OCPxLicwBfCNvN0V79Gsqsp5KPzTinIi1zyoyAzw
DOGC1dTY5Srd9VynLJH/lrpLYsuQAtVElpC6lk8Y9SYXgIa63cuvrcKogh58cmdv
QvnkTGgBPD0f6ys6HDCGb246ClT1HRB7jgVhL3cRccKUKyoRg8uVJo6CZqQ3f8q0
I8i5MUt2YnxLB4CIWaMjS4dY1WuYlQW/J5pR/BMZa2WDdIcT4gwMV16yhGXLz+ul
Mu4YAXXMw8eOH+RkqBJGRr3/KTNxsfZWQBF03Sd/EPRGYfPK/i+3CiCcuvXKG+9V
8wkTblxRnzNvvya0zpx8CxwLBmZ0w4wwWyZj4Xa59rjBj2Jxa0NluYM5R6gevJz7
1E9HA0Ed2yIzeRfNLRp0l41iQoui3I7lFPvPUy7vQedhJXR/Du3XbqrSzvs4lS8r
7ggNGCfr5jfqrTz1gr9h9uvypQzJsXVFkBeetkxeey3WwJ9RlyvInTemRMjabPVX
d4njCKl92tiaxdDfSIjzlzKx9acNxzsz2XOLhlTusm7YEnoYwnc+kQc9QuyTVnqq
fAa+M65iAzHb0ypuwl52pmCzz8HlfkGFfQ98PPRBjDThCiyr72OhpH1hnBpNz85l
JhMWEWCgA4tNPb5FG/hR8/9Wl92XR5FT+4OKXeq4s/KDsP9dTscMN8Jww96VQnpJ
O0vw60ioO8UCubgvAx7XQu/aEUxZ0C4qUZLzsHVC1c2f9lIYjDxPL2pyFqif4S7c
Bz2tGHMi269lq8rUK0wWqZZuTrO/6nm8GysrohFwdTmhhiPZyD8UTA0x+kILbOva
WVXyuV+0O1+jwOE+1pwzi6qv2cYgOuagQAmgH2StPkid6wG9ag1MwPYSp0pP5cP9
QrX7RpBLmQ+XCylFcg3fx7OyoF005xDQX6bxo1TseoCZYh/hYUVX/A5W/Z0iJxaV
RM4AG6G5vErqVaYIjFurjYXZd/UFi76LtlRwBp04McU6GWPQYUH+t9AbVsVfHM61
jpdor6HRPcS0/HKNycc5SCTA5JefOhsdVGmMbACO/L3mIN/qk95YI3Lbui/qFo8z
2O0JV9M8fhgFUryBrbvpQi0WOCGSTNMjQbFL7MwerQDJt7TWmZDSaFo6TC37NQI4
Phri0ikzqhWrXa/QNIoeMW+tZvyhIpn5EKgWRNhe879quXB+hALL5VRTjCUMY82/
3csw7AsGs4bVvgol1CbSzxGiiRLlU5blJKGDdUDVChFFafGIS3nAF40bTguCENNV
uW+jnd3pvUJFHIfiEwLprEAD5J+gCIMwTSmzaiMTVILvfKGJ7f8JAQSDKLjt+LkT
9J004p0cgRtHHtQNzHU+VqvwIyhFUs2QNVADCGNsKrING1351w6ZrweoxX3eToB6
GdxCE4wfpQwr00P6lUyjs/ogw3wpU8khgyEFmFBIruzdJhBW7wp+FClDXuC6xiVQ
KKc56HYNV1lQeQ+gaQuvykfEHyKcnuyM3pPRSwHAsBD5RBzZa02wHec9vcbOzVnh
zrHJmy2427x3LM2UToWZh7ogRUea3zFYIF0rtyomZQQkgmB55Dn2cXIUKC0uF7Cc
FkgDDNfRXaUnv5NL4ZuvtNgxBaKk6MI3glfXY2XCC//FoGtnTVGNL3SDO8yoPdkX
IYr8Jh6UyESwnVas+UsKmt+dJJYl1xptaVNDQLdYcYzqhVnRvP2lEuwOVzMz1WCf
kU/oIaNQupxiByEetHzrY9uMXeacj5TUYZBhZFrK4c0xuzpMHzHu4jtlRM4GfIgR
tEpuHFKSN+HYJWppc6PnP2kUUXH3Y/qBX9XPb8ylktDJkx+g3+tQqnpH9J27eaMj
PaIZjywR+SVPqKuQar5FPmL9SS0RMMgDLRLr5LuFuc4gF7AtaDAlLp++ElsIhiHr
3ZjJ1U5VSqUKu0WGMJuL/ztEpjFomboqXfajNYdAEiTMEcsniU/lm17E9EfTU7ZB
JL/gFJBCxwEjr5jG8VHwK0AAz8lZ4rvh+pL+UJHzmvUkAavYGbTvVZaInSCD7zYf
dfOKqjLGiB0UfIFnafetObM/NLHF6wD06jYo27EZF8jp1J5ts8SQchg5viQ5GsEi
OQyAXyVso8nb+4Fd+KrsZtHt1WRUefUCGo2b0dgahy3pSO3zABsWq3FrDzwCbm8w
J1JvBjuR0/lK34S/B/COCE0ChDGz2rd1xrn6B09KwdcSsUhXphX4bk0iM0cehy+P
SS1Z9Q9yH90XmBe7pKT/I6Lm18qzh81vlyKvncHc7ncr2t5hKL6KKvnlsoglVTQe
d08/IeSNxpoKmmj5tb58fIKWTJqGq0ItRqbo6nF0H+/gFdw1iIMw+gd+EHORmOyt
Xj1EThlVYk/+ufhVG9UH9V5FKo37v1z+xP6t9e8o+HHmzpxcHWAtZE1Qrin35h0s
lm6OsCbnkmKn18o4g43VD2QU4qgYkIHUB/kwpzODhT0Zct+QP73u8/qRH+bKtI6J
/wTqQOwEfnlX/OkKRq7A5nMovdBJJ9jVTibdb4jqD3DKmaoN4Tc2MUiygYvQscq0
GEMncC72MUlBDOQUXBIpCKEMlmBD5M2MWjfJaKcX3+z8NqQhMrT0R/Y2a0v7Pjnc
c5VzZXNkGBb6YZ+zEz/zz5HRuqeUMtJQD5JJZpo+1JpG+24wqS+BFC9Ou9xEWyvk
Jeejex3iGSB5yvwlY+cgxjRr8X1mTj3s0lGSCiglxKHrmPtRqu8FNnUrcKFrW7O3
2dcaIrzPZavEUM+sGuG1D4SJfYn7mJP5++SYJnyZc2s+KVLneF9/GjIr/LqUCbEg
9tWYOj31IVItHHtg4EdKZd1nsf/e/ukxG52YhhNX2ZViPPjkslw9A77WWUI1k7b5
NrpfuxjWu1zq6UP5BK6jqcYIwSz8d6BUWV8ilZFsqMjjtc5XmwpThG/ta5cRXw3e
BAX3dZZn2pQXeLX4kx71VM7XXPS/FCjXNVGwzKN8/PstL3IedyzeUrNKO0Nwc15g
yRWaNokXAgpgtuYgdSRSoCvq0yqazVIAU6A8es2cXJaOyjWPL32Zpg06BeboG6TN
ebtmX/9p7tHHF2lJMBuuSSlXjbRccTCEYMqgvUsXJzL35S/K2cPO+fvpjvAyoCo5
uUzSOu+ikA3rvimQUZeXnwENmqZjzAfPIYNk0M/b3ZENkwwRc/LV2aQmH8+SibDe
Q3tLzwpzCsHGsm5w5k8Q87cbCKtpeustZ6oK9L3bZbtJ4qhN2F7kuVhBqjhXn5Q3
xTlAgYS+LbBSKIe7VegWR6V45LumaxAQ1jVE48a+WNHS4vEngdvgNhHynuCyi1uM
MSnGdhPhkK18Ou/u6aGxooX+ZYS0b0jcpoLh23HVn1EVyiQ4c8tWSWP5DFcHOPl9
iY6Q+9xv/cutYcE12wRMpMq56QCuv+kTwAbuPYskznvNlo2DNNLK21Q77Keunpp0
lNURD+1apoipuk67nVk1Ew3Vtz0JMRzX3oYuL39z33oTuEoOkZV3FGiVh3rT9pjl
GxJiUJKAZKyqhgnYoshDoFfhs7iUrEggXF6tOs/uOI2D0+8Bg2WhXlqTngAhUKgL
pTJ26u0nZ/sHV2IC3MP1y9JwihhEmcPxhbjQT/ssl2N1Kyyehc2aRUAp0J04jthy
MO+ms2m7Wg9roh2AHdhXyPfVb4m0bZPcrmO9ua8IFW2QklP95t7V1GbuimRtWeMJ
F64azmXd+aSj3LT0zoBLfyK5UnIkykSsG5fUnPV0YbvyhA64Q/0wIxbNMKvJ95Yg
aY5l6Jvz+4/mqVeG5Wc/UkpKs3YsxsctYZzpY9gcv8+gsn5xEihTYO6+F6z/i6uR
CA0NgSduKe1JGgBxyFj7jX0a73XIz0oYM/SH1iOfPkTuhYyzgXNYs0SOlrM4NGlq
VRdLS6r4E8ONG4hzicWIpCTPLJUdmbJaDikNxYLbmoR4smYBqmvWNzRG05pqcrkN
dGtSX6/d3ccKS2Ns8SJKcX1HvTEdOuRxapPJn9b8OXyuwA9wqTi5qRxEhXZrs4sq
jyBIJsqi91stkp4+udJ7bB4YGGc/eLudkwHpapPUpPepg50pHfVTPf9ctt0GjBsq
c58kgpiJjp82x+/hCQQvykNBHYmChVIjHzwRuHkmIuIGtbFc1GQpLNofOJoynNYH
/hFBVqXLm73OzTL4LhRu8MoS8C9R6Cps2gN+LjcfuzZnsLPGbtVLqSdr9/v/y2s1
p/ivu4kn59oVJey/ZofcBFGGAk7o+A0O28K5odYE9W+/RnLwXGEdWQy52MhlPL0K
Q9D7bZ/BTEQdYA9gBMFWfBl0hIS5viKstxF05iuNvv+3PNVu5muc2Y0/A+qbsLPn
oKbACff6g1vdbLCkU/m7F8NeYjLvx0T+Yu214Y59tJs4G1iCHzHrkPdN8XRAMG+0
foayfO/Zl0WJ+W3uTQFipZ52kjuOUsql3IopkDmjgTx700NCm8XWp9XHlJWxi4Z2
FW1N0KmyfzD8paTCfIHlm6hcRps9AEkeItFs4y8popTPHKNreQcsEQ4QeAmRkk/T
r3Nn9kJqp2lkIZ9Br/6lq2MkYUuW2oEQISIltMBhcYZIxilCN108XMjVUjOS32OX
jFDtS/v8YmzdrBHBzR/LsZ6DTwDcF8GlMQV2X8TDZ3vBIkXkBQFaXhhYtc+PrCjo
3SWLFYxl1HEZH0UTDTf9D05UVfCvWdhT1Qc7iP5LaZwQbq/rkSQBStyhP3tevJnQ
KPRv3ovkKBHtsfgGfMkkrptBvPFgfaxwtxnqselaMKjqGF600hFQWo2JP/dFMq+P
AefQ7JSA7Up2CJYtNfQ7j0zvrKFnNpNK4rw3BkXAclLJYLloz8bp6/RStaooJ8xu
jdzn9veLj0a5DBEcxsSpMlyCElciK2nMwu/Jg5LuuFqj39061mFa3exqWzBT+Zs+
h+B6Bb7fCsDihFQEJ6VWdIKh0B/2lk3C3DHkL4B7q8HUt0h75m+vFSE5GrhqDUW+
DVCpbkE2y0wBfzuY9cBEfKhJqQE8QyTvwnH8MDSQWQF6m57JngX+cCWvsrvtDo+N
d11tozOhjxYeq0hjeEuso+gUdC4CFS/JHRaiZNoXgRsjzAb6FNfeBDLE/AC7gySA
VT8cat9yM2UQFMXgfrLRIltTDOgFD23d9uwgFC1F1/O/7XTxa/5t/JQ9+d3he7wx
3iHSyuQ137nYuuruTDxSRhPzX4XbYiupIBZbWrMq7Jse0pFPyOjGhwlca+QRphsY
zddIwCxBMrlAz05bnGubr1x/1sUzTo3pIeQ5PWTdpLC07LKQe37bHMO87x29J4ky
Uxl8qRytf2ebnzc0cT95ykAlo/EUxdgNZvhg5Xr9suvXD8ALS+9BziEHZ1G+fFX1
FI4lJBzJz/Fi1zkEbH1p7yNfalHt2p86wKa7psVM0QTL/zHmiG5QeiTQFaVsGrly
VggWt3vfh/RKSPoI/dVa1Xzm+X053QQ1NzNqHWI+xqKsBm7quAlYdT2j+tKKIjue
vT7YjRfhRZBfzpnmjjIEWKaH6z9GtFkVKqUIl04GRvEPm2m6BZRrd+h9R3szRYQL
EXbu80PtFUjRCw8AcIkX8rtLcMXhS8Ra0ed/RzXmbPpG/sn7jCYFVpnXzrIm6n2n
udZjQ1yml/UK3jvWhswLlWBQ+Hmic6Qe0TiVO+X6w1VE188CJG0fGS4tIDxWJhnh
Fy2shwgpOAnyIY8EHHkiOEjQdSG7IQ9R8J4LB74HlkUo7PsDpQsY93aXjw1n8JHM
mm09ABGCZxbhnfG9TVyuEPwXigug/5VuUN1ARTMc7hf3HYOFXxUolYgDvyH+HHgn
e6UY6MbtUa7R2Is035JmGYX+EgnSUjL4Aa1uFfHT1pGxz36VV0TDDX40WyKhoC+Z
2d/uZualachmx//65aeJtkbn76z3jVGnwgjsg2ZOIx9HNzWoM7cFLiTYRUCw+qaV
tIk0sn8RYqjMPBtPDxM0GYEDjdv4ipNq9lglmkSSPuJJ4w368fpKkWbH99ACCZrz
2gcFTPaP6F0N3XOVa/yHPp80GJAPBNJFqaAuIRzS3E0WBIqyAw/tG2jAA8G6AByP
vDk5HDA3DpgyY51FBOhhw2iOE0fwn2kF/Th/pAUUSL+mm6rWxWGeHV3H0bW4hudA
/85ILPyMXkU0ylNDTqO50Csw1dBr02y+HAzty1ESjPL9XHZvzyewQJPPc1C7aNLG
kgC/xpDDuQDEpfHzY8IAfZBOpBbFdOnjEg52ErTUpesFifDJqFJFhupH3AsLh8xl
H7yfYJWPehtSywa/iETaRADyVX/CCKAEX2YGJbxX+0JJQ6t4cg61nOJ26b4Bb3sD
6WJpXpDAipOYFbT3MuiGhybxoDNO7W35P5C8VKVqI4rTKa84UCqUmGEXI0h4REhE
xggwOWiHWUDJpK+6OEA8YdKjdMAyiyqstKE8lVeWja0HIWmbXYrrzzZUGHJsRQsC
uRPszfR0YmckzWALBwbtcxOmv7/Wl+u0LFz5YyFCJ4T7iJ8PvncCKV6NUx7ERp3d
9gk0cgieacTyzf498y62cpVID21mQKjg5vKn/ackxxXpwTS34SwxJ9YCFKb19PsE
deeyuL9pCOnxkudXXWBrdPxaJ2y6HMlshLNnP6IQF/NTKO1erVQ4Yc5184dhCxdu
zgmjJBw1UUi1ANPCua0BD99aTb6HPgy4BJ+Y1RpoHdX3ENh/xIGqbboz8Y6uesjk
w6jwQyA4muQZG2UE6YE4geFbxf1NHPoNFb3mKs6YXq9WlMtWpXcuT4aQsvJsTxwk
g6ai/33eqDrg1af0b/KR1+f2Efi7rOSDwGPvENjIiPUMrE1e3kg8t9OVwQxE9SxE
UNPAFMHgcAjHLX7/AwscFSmBXrqwXgFBjz1hr5tt5yCUMHrCokuPulITw97Erj4W
gj80PT+zahM6YUIBGiEA09lg/elmeMQGQcF/KCSwDKPHLEc9m4G+8073Xfh8FClt
iDXZNqDPc34eHyFPp16q5jFdgX7/o+QDtVAEny30LbXa3pXtfeimU+wK1JghPxTO
ItATWA52q9lCjSqxegTSL/Ksf2oE7bLuxWlN3xwOtny5S7LywYjHzWaLvZ6FUrxS
O/F6N6kYvHozQuPel9U0csucgo2TDMtpbVHtaDEIBtvf4kGZBS0N1K0KHEPr3nmj
kO8nV4JsQ5D3adwdK4pv5OPIlGcpOvvb60sObVR7BNLOFDiMvf6WBMIkHxg3jZQD
EYPLIn/nqZ1L3s09eWzvcVPF2HFgtmrl1/qI1PelzxJO87XhJjyfDjfyI0Qe/hRP
N6uI4HxTSoFi24dswfXaxabq1opZmiWoN7udjHkor3hwx9SH0AesuCxIsdABsVKC
uohp0sh0EIo/aTMgRyTVpy3Ge1oiZpfOTlno4foGzQ6aQ/VIE1CKMz564A1PUuXQ
uGSWHg6ZS9luEtjT7Viog4L7NumkKprDafIYNUW2Zxqx7QwpraqNfIx/r9KPC6Ok
pysa3VZoUnCVkIy2OsDiGRE8g8uozu/CVaShtSvxOB6M7zCtLKBIYGE9bNId12To
aftbpPuLe+knF6kwDS4gHkqsiQEKj1FG8iEDkqqdHkjiA38Kyqx3Ui3E8m2NWii6
m9lWTqvYy8v0wOINsjIuptLoAOFjIo+/RJkVHG/stG2pIlj/exe4lIJaZoQ6G98o
oCt+V3TIZdjzDYZPZ8o4VWwipJz/HWyIvhDogewtbxZg9D/ajkXkcMfJ5KWHvv9E
Bv1nwGowC44UJQmAj6vcFnies0Mpg78clJTacDjDKWWXMxd17zcORMKf5yjkiEwr
FfhMBlsLUbUIHgZUzXkx/oAdD+S254i6q4oVie16pB1fiyWNjBF5a7WmxzWJPype
+Yp0a53ffgCSeZBrZACqdxjno7M7V58p+2Sg+L6P2pq2Xbyr1xNJTg6X3TX94n3G
8BXt4DWo44jW5PhYP6lvQHvcsfhySDLBmCjsq71IJuZhyD04u5zhQP4d2Auu1W3A
1WJ/wwkLTr+DiepMa414+nZTtpRV8XU8qVtK9T8mukpDjFtYyMCDTh4GJgpYaoQV
93GDd/VWt6fSu/bYDOZX3ghH1cvKlsudzj8Cmrx1RJviDrATlZNZBy1GFpkyU+FF
vQn8JU9bnI48IEWdbCmCaz4jwby4X7Hx2KntsuptVCGw/qyEUim0Txmyi/lSyZyh
9KpyT6aRa+wyevMEwj8VCbRkqu45sKofR6R4ONcoY03Ew0VRiJttj2+fX86dfaZB
+31bfMtfYqh00suVP9mCBC1+vY0k1L5EdCmwAo5MkH20e958vxK67ebu8u8HVFRF
7lPLlmG8HaRvTGPOYrDWcwH3DHXY7RpHEF0NEWaSenxk+FLLob+VbH0Up72piuMe
YeH4rQtdqyg7z8E+3gsOEVDO12x4wZAfwr+/zV8g5auGjpvZuCSlF1jZ8ba/RA9/
Fxt0ubE9bhMcVs1WPxhIe/OboqdiW6DUtVWWlRzRysqF8EZbkgPq+rKTMaNr50BI
+W7LbK62PJ6lEjgLhrEJMFH++lp/18Fh7hRfkHbQ9b3+koF8o3wmid9Z6EvgLTN5
mj8/zdHOYKaeUTTrIvRpVwxjQmo58AtiVXxeC42Vyeqvt5Isq+GPugGjTnaisgzX
chCEAUgHw5CFzkUX3wdm2nyaHwwCcjQvVJFNp5SjJA2B3w2tjGmp4Kjn3QfRJscY
uxl5r0Yrsh3fhqp9Ex4pP7taa8EKvnwpggcSoEFHz0x+nTkIp7zqF18ub/FlUpIE
7jguiNeH7sYiNC4UjgSMIAVb0q5Qov2YmIwTRI0AXYKxxvvSboYpV2KZzWihAjpT
GB+7+mC0w17zWNPxJUCClEGPeqeLUe0wlmFVK5/RAwgr2KVHjQywnMxJLF+GEc6D
kb9Ck55aE9AB6ZWM7gDN4IZQqJkPev3entNsnfxKVzdoEL71tEBRx7ZcKTr5pB6y
ohX6s9y39fJOwmOCJVE3W+g6DGTV+l8+FNiX5cNXTtApjrh3CP0uYcdHrdphHR/7
/5hVkhW6SPQ4Hu+cle1EGXjgHp4L5PlXEbJpunqQxVDVCZR/cxWnOyCUmv1RdP3/
9s/i4ZT7yPx5pNY1XDX0UDQ+EBW0R2aRpNfjlohAmdCr2ZXjMxQcbvg6BPmVq0fX
2f3fS0ZjWvk6/NBqpoQJsKobALUr7rI99g6Juvmm8OKFZRXqXkBMQrKmGwBlAgsl
Y+RFwfB/sQnxjXhCYJ/THUlI3p4EfTwbhAHyxxHaNIBFDCjc0T/y+GXVgKmXeZZz
X2VLAakrgyiiHH2Gr5dIerw6OTuchb3j/WGDNPKIvbamh7aGADqsq6nM9Bxf5r4J
k+b5Vw6uIzK4XyND+nf3yRPKVbUqRevPbS5HXQFLre59hPnQjNvDQLEjK6k7yOZT
IBIH5BFM4E/Lea42upFo6XgbgsOysVLyQcWwDz+VWgZ5QDoh29QMnCNWujkxTAlG
AP01abm0FFU88Zwh7NpDW1fS72SwucSyLE/X9Qihclf1GFyV7HhZrCOYhbYV002d
WL7if7doOfb+y7nqv9Wq7SsyNsw98w5An52SLDFR6iJ4DLj2jIfxaWAxVnLJiJgE
AiiuRcMYFtij+I4seRdGAYf9FNSQ1sa9DLAIDkN2DE8Bbb0hC7zds08Xmu0i2/k4
HO3Fc3oZ60l/1TSb1jfWUjHqVbY8nKau6juh6Utjq8coL89walc/hW/FgdMYR86r
6thPOUb8KTfAevuImWPwFPPS0fI8pKEp2E6eNF0uxaeHCjOfmVUP6UTSrgmJeaDu
+FpOrjDt841oWuDUtmzas2NL+GWQLM6jQ70qeKPg9vxIgup66Ve9vPsAuREKFnGM
cXpGHdYgs2Xbr06hQhoqBoylCzpR4rOqFvQTkdJml0TtEU9AU6dCFL+2qrMr4gh3
rMwi6C6hxeIFG1vAm6ANIt0elpc/Ln/d5svDf4RPfQkQf1TDxXkttdzd6prriRWC
RjcXtjns+1AdhPGzftr3eoT2Z4oOO+Iq1Cj0w6cnUcljNw4fmHr0/kfE5AIVMm22
+1JWU5nLsOrjY4L/NysDprAm0NuDRoigvbz6BpGdsc+mlYY2aS1nGA1kie0/1vBy
Ae9/mYqc22ShwEviz40dqpWOVRmvBu9M2VPImdD/W6Nk0LIwLOJniLcTk/G3c5/s
dyzf+YYGSwooK8zWNy6sSKuWsnCTs/yZL1MknFCbO6J1zSufsZTVxylMKRMkEorr
wyqLneZtTCeHA8tTCOCeEw1fM/7yw8uw9pcKXvtWPAbOuEY93f8IjBHpdru7lfQw
mHqtf/wHYBTnshH1ptspy/J2hUycqGiT+bgnjuPhcw7nbv+baxqhiB5Bp8KQGLtl
DLFPsDeEfnG5m/5FY0eksI0CQiIfG5RSY08O/TLM0EpkKR4vGCpdnu/NL3eK4Fft
ka6U11rzt2maC6zYP8lhra/enhlY02U/JvSI4n6iQEzZL5dTJxx5N96wteydqOGQ
IWIijctTMczGTEj9Poaq83PENAq+GQGmkRd+UJAtKz6c6q0HZ6PbIfT4uXkK4xTh
sj1i+2oO9z890nRbw/I7QTLAl0G28XYqJ3WaFkMG2Xl/4PWv8ymyK2GaEQI7nXJw
hWzFLiq4WmvGT/XJ5ULA9ttaJTRoz6+pOHEf65hUL5/WH3LPbqYpu4iKNgc8xI13
xD4zYXix8hh8/OiRmO0o0Ha0I5UFFsx0frMG6UrMB4orOJGDseb3ILjkWDt08iNP
7YvBsV1JwRaXkDBp364iEkoL0BsZraSvFTWaif0bOCIksvdWjRTeqzRrK68t09y1
D5N5Ja3U0mCy1mTxZWVXHFOm5ozwZKSKdk332blBDp4K/Jfa9lqxJsOfVGbf4U/w
J4nKswnjXXcvQ498cXfaP1gLxILDiYfGgxIv70hs6RBbLNuBjySJFNxuqrwkdgIL
jJoP10e57Wgnms8FXcclrmpWx3SsgoUuj5GhjP0RpCVWIIqt9UYLSYPJ+tanxu8v
t3tRUUuHFa7mJRIQOjYnS4ryIAAd03tO//Wn/rthLYKpivoL5holOa8IVjDJE8fj
efVGjf7sAdCoWboMaCw9b3OgDUVHaj+1YpZUedRJFijvNwIKfx0kCKP/8imJj7k6
KzMyPY+XJcJ9thflPlxvKrQ17RMDxwKHiIw82CVRoVgIRc4RM6YyBD7/HYwVePbh
GKap6Umkn0uSHQKKSxA6xTjexc29HNYs/8P8oTewS3jdCYeYSfqlGTFxii6KT77L
3pjsKwp0Qy4Nfz5WenA/t2OsXJsRdjAHqwVMUEALQO9zl0bkMqPQDHQUxyZaCf+h
r/JLV4H24Re3dzTBQ6KYtZGElhugaBZ0T+NAMlC7mc3y96FrPqV6lB2OuI8dm4Lq
LYz+Rwi2Gf8WpD2OPFisuAEPP55uCXagHMIkbNVjgmxzlHBt6r5MxYJuFexFq7KA
yeS/kQD9A7TktY90WDJCG6GvfUS8pXWaylIvXvEdhWcoHqJ4fDH98cbGChO8jfb9
Nb3guZVMfMN7x6vpCm9s/tDoSYk/c+sfMQahEGyRc45g2uMC4Una1p5AFMIv337B
Rv4GaPhGrrw99vyFVbYYIchEkHCqwNEop7ySbB5nSDQchi/3vbaWdB/0MSrTAisD
j7hLALEvJPWqGV+KCHDZ/BCnxymVFohE0Sndi20dr5K4XhrzvcKCDCabeh66K7GY
mAb6ns0lADpOIEAtKdDSq1oPEUANzzTunUO+khNEL/rWy6kwjw6/mv7QaTUuZWaU
YokwDTLPcq77vE0ecjLuRyy+neVYj2ot9QmBzKWTBcoxEVA9WL7qCYjq76QwHUlX
nRbktb3VUvRZA8xxbxpP8PUM71+Hk8uXijbO6btNth2AY3wkZntnioCQXEPkIYX3
fom5ZPCu8LjKcBpsfK77j5g7/esC4XNZ0r/jYJyJN27nizMiDj1bS1eFyc+caasf
lDEjXBzmsNfh2Rpmk+35SXq/l/chMZqetTwpSCYSuH0qBBM62UGx6S5TKDE0jOj3
xbid4DkvOLViPscqBJ2twFOsiGmIuSoSOj5EC9UHaAmcqu8HUWJcJWtf6t1jShT0
KKWIdg1ylNjW7yEtZ3mvniPlakFbQGz/CL7x9SxahUBL9ljTP91E62hllpYtvftT
j8NDZGjiAWg5LHLumG4HnMD/ZquxChNLr9oEPmRiTxmas+gyxy7oAg+5zJudKwsO
rrD4awnxkFf3gZEt1S9/JA44fWSGKcxZPRl0kyjK3uiuQUWdIBaUa8jDgyVqXDvX
odVxydtDETb6cVlkKvNzFUZfNe6VrcHKZe4s2PTBYAh8A02ZuI1GbS6lc366ZL/s
bn927ppTZDqcEHU1SLmbID6obHHGuTs7kH4wENxDCYpkKm95i33KoujiRKCLBwHt
Xj/i6SHmlpVPm7jD5MibQVqBu9VZxzSRm5/NvZN3S83WzpNWmAdOPR3vmmkQzon2
CGbGIRcTDTcHae8phc487w86zTIlOe6MlEbI9WtCrfleI2udt7hs8+e73v2dNjV5
MJzfGsgDlqtznGOEraxTjhU1oDYCSCjMpBzu/QgB5VApVZQzKf6i3HAhK5WfaKfQ
2QWOoBHzkdIQf3XRWgGH4UyCXxSZL5csFC5Ru4u023zqJZrUB791oS8BTAUTFqSM
neVBiChVDO/m1BU9yAinfAQxsWvYIke0N5mb79WuYFSXhd+HWD+OYtQ3aQ/hPW8b
j267K+PHKQOKZXIqwH57ne98csJmtv9ZlKniMQS/vgQ8/G+zoIDIMxJYLvhSZorO
dhL8HKk7TrtAjT3UcnOnswTqMeXb9ZvAVCT/sBRtvHlo1UPaqh+Z/zUExMnI/pxh
H9PDd1kLrNtb94ADC2FTin3lBuixdqEllmV24tmkEQnhY2tzwlHbsh8xm3pP/7AK
L0v1UBpbJd7JX6nDzCMG+Yo2gkC2L73RGwF7UlGh1gDRCyQbOM7+ozuMb0WC6Arx
WWd1LhmVIOB/IQiJ26W5GRIcL70YMf6+ItlLo3C5/OqQTWA0SPZ7zMCr+oDHWqrE
g0Ewz4KtWv2SXsu3wgTSKlXkaXVQ8BTaUyneZw3cYEd5QvIZKtOIzk78RbYTwObt
3xSNAGeddu7PdQrI6xar2Wn45jsj2C7QjevmKa8Md9nnktWE2JkpLDzYiJhdRCkd
iRWdmaDF+9kCJhsj3F63Vvp0ulCjx7rN34Tqhm8dNrLmxjCgerHlU+FmldMsz3a/
QGN7icAU/RU1uQU1rVWb6M750bK92awaB+U/oFKbU5CugVhvLvcJg/+boRRDz07j
sfqNFWIFh6hXUy4ATc1JaMUpCE1GTCL12LwgaUqcs1Q0e3b74Qtde+6cICvVsLle
4G9RMj239vcJglb/LxG+l/6vlone4VuuUiVtQwsajsdyOui1kFUYnzEM+2ywhmwQ
XFVDucwYeHCwHNu7rTnNtVlmYdVIMt+d1lP4Z/n5vb3XiP1NQua0+Lz4raiwin66
8Gqje3+/psyn8ATaT7djlz1yI5xrNsOjLS19JL29tR5SD8Ql/QlBqErq1F8CSb8X
CLci0zcdnm0y1B096Ad7+pjyb+54jERY/FWl4Uu42GBxTvDbruQgLqgJz3wb4yZU
urwJkKUK1ARHZSdrJCkBOBnSGozw+2EzOywq5ol55LqLNt9rZW8hOfS98q0TJg86
8hHtT2tpvIOdtulu2b4/HA4Gz3Yyk6lgNjdDmu6GWzJDaVBV7BYxNWlz9AKwt+Dh
66oqQ+qcmIg4Fe80zU5yvroo3GXpoNpIkQ/BC/JNYBFSRjWm3snJyVhxksk/nIQh
t1jIJUleQaknwARL3v4zZyNamDGhafB9J+6ReH7ai0nh9LQ6eiMOC0rsTuyOf8t7
bcu1xDggXVJyZ3FruxokJQmp/kf9I2ITeCiwGK/Q9XFa3mGT+y8akiGOcDoEPZNY
vT88vpT+bmfDm78bsAPedBotSYWcF2gQ5TOO3ryucCfd2TvUiwew7bbOCMw8AYYq
+p7UtY16TWmS0fChQXL1CBNAOGRWESuYBZbqXDvaPTFBii260IQeC8P50fZQd5TU
0EuignRhWbMyIImQ5Exdd39ey6qBxDl0wjzCOPdmO2Wdyl+vG7VNB484Zk2K4aN7
Xupacl+vuTVYjBPK9h8ce4STdU0Rp/cWdklDNx9D0M9nG2MKwJVIP9NMPV143P6u
H1Nd0bMOAlkArH3LjcjsZIl56zTpnP8dLPTguMJ/nfu2cC4p1ZDjkWZSckc0v3B1
Zg7rWyd+a9+YQPqoflUVA6zUVWPU4EOpXDAkK0Mt52TD3e7lUyQKyTAb7oViWc4J
bOT21BRRE4P4gHu5f8nuqo9Wxme/zybvxgF8Mit0ymSNKBgnQckZT13WCuC7sbak
UHVCcjqqdlcdkoRboBEV9w8xnvz9Xx0ux/rkaLgFgW5TLJoIG8VUl2hE2pQG3puG
1tpp6N3fFzB14D5pzTe7KS56+099fHPdvaYFwAL8puO4A2qaHXrWIHl8yioeYXfr
RgXT8pj2Wjh//FIa/S3d/5bclTdXEG/gla886UrbgvSmdw0e7N8Eo241EWKMQqOM
srcpOZ3qJ5UmJ6FE20hZxKNiwrrR4v/z0e1+0i6hMxUQEYiQoPbBCKdxSWPjv67+
McxNG72Hi6FCSVYbFbJ/QW2/IiC4i/E1W1veV07ciaLW9I5y6GxZ1oCykW6vgtKA
jQk1A71WK6WzzAOMSS/hXzzK3y8XfdD4TgLuM2nMw5o7vn2aBzgZSOTUey2bT8l9
e5r13CAXYloKyIpTd6kzAhGP1NrRp3p8eLw803OB1xKqmZT4mr5arrUTFiIp141r
tXLI6/bPpcK/SDJflmtwGHF1PHtkMpFXeSjgoxjV4G4iyyHOKyIx5DO2I1Dfe/q/
FlwFNDzd7amAljR4nK4bboLHLjct5/A9jMwzjWbZvOwNhXQixjA8k2bfHLi3z5vE
WuTIzZ6oJq7mBBzsZCDc5bD4gWQIqww6gQ5IGKmXhpPtxCwop1+oG+q/2uvfHw/f
VWnBe6ebhXDf4SiSfAbJkF7c8OpK7629y98DR/gersJ5sCiNfJFKoiVJWIufpnQV
eAxIqY4KSGTanaGkzfnQyrgUbymBOcq959FrXm8gz01dbzx6bnUvo1Tndd3t2YMY
U31LTUCfLBqb31pvXGoo6vFgMiBiTHJo9JkaYYZFDfeNg9LIRUUox20ziuQf85MU
Psq6iDU6QjptKork1irPJhMblNKQV/uxPapa6it8CXBrr7Qmb/miDGEykYM+XsuS
0dcDjc3VF3vC92EzpWapyGl+JjKbxWEOOSSfdSc796id93d036lgxNyFQusmaIbd
o7ZZu/MXSKMNhLPRYUg1RMhKGeuFC0N+ZEJ1jgICbV2xO3Pvv+/m9gBK76L5DDHF
aslCLIEfK8ZewVRH1kkKcAQSN34HJQzQek8ZjFleBi6bBHPDuEhFNIXOW1yj/KnF
1/hqDVVp3/Qz0TVwO5lvF/PvYVdofEXMNhUbSAogoHAQBu0pPwlHi672MCwJmyM2
ImrHHGIxXZ3ONoN7XzPZ37gEhh+Jv/XzNphyuv2FJpDJNyZ+8xAz7lrjdinlgJEV
f/RPhxlwZpbm+wRjV2DLzpi+Iy6qlpwm35gCrkH0akn+tFKi3MpznSYEsfoU/OpO
qwbkAeNUU6YmJoBFPWgLu8qo/1vZBD/XUpD6/fOTO3rzgtqKDs7G/MzHsCE+vide
iRLkSMNM8XEsFg5EW+eqjZNQDPINjfu41b5O6utvlhJZIXJEh/YVan5b7X0qOMRO
FM4wV3fWiHUDcRJWNTSzCyl14rijZ5S5BydfrS/6J4diWd+SNWBUqBxAsAp5jCwa
Ma2ToQH356xg0Lz8ozuRyM2SrHx8mqsO+o17bo82Uuo/9MluxtCWiMTf5UCIiwrv
5FabALkNBhmOh8YFduknYpx+fZyEtdMi445S9VQEj6RyoW0i41Lazl1u2Kn7gxZ5
8uuMJE4kaOOhTlkUn8DUpqBOfo0/UqJ83pFEcJFQwEvsQqylmyD8LnYfbxOVelUQ
3z8Zw6Dzif2ScONuJEG2A4YqhdZ7AWrYwid70QBoN89QGIS46nNeTVB1f1KGnbkK
vnDoLmBmDJNGABr1c4eRiM1QDJdLgMYRaZBC7PdmWBepBpT0K62dk3Yb4yP+COhh
aK6vBIqWDbhXIg96XvoiyK6XzmFuvVSYOagPrhcVdChYrjEd5hZlKVOv3XyTohmJ
7QYUEMYgK1n2iW6ouDuFVbvNrGy14c1F38tgnnwjtmprkjRoHPRCi/zJkWU6r5q0
zOBQUlMbIjFj57xttgZ6eB50ot2V8MXQYn+T3xDAcDoEAQQ5GgEV9JNdRka/+Bdh
cag6s6SkISRoX2edpSQLJJYP7Wce28KBFqIHqRnYJrYjtF5clk/JsHa/QLEzmm4U
J/FB1OKnfZPg3Mqe7QPPZ1SrtmHQQMH/FEHjeykDeSH8+fVvN83qMpjQ98aDFVRD
FdIgrnhwhjnEon18yj+MU+KYnwJSrLKgbzVh7Sk/Al57IH/x3C2fCzA2KmVZOLQc
ImreZx9gHGKEnwP3T14eqKS7oarEoKXxFhqKQ7gn/9wGoGZMgMei2YW4E9BOJOUe
DgjC3I+pkO6aNRjyBG6igpbyi/WkW1IVEGMtfUMC8bEeUV6JgnRh5dKSsmNzX1Fz
uzRDg7PU16UfFCWTuo4EY6+3ZRpUXt3nTFiaJMtujwIj2qrMhPu9rucWr1dCvbwl
mal7+FM4Q6b4Ie94yw4t1Fh0BHYXveue41gQMADZrpwlUY+6qgO9hSvOBNJc22VI
S7dWEQy5gHZ2LRMHb93yEO0nDi4n096DTZABZizeyR0lH8Zft5UMecN+j3yrgGeg
KXa6GGKyXgyxEMcPqChEpDTUnNiYrrYhaXRMVpwJD/w1BFYPbpJsywgvikzQ3xSb
ax+zUnGBMJm1W7dFYQTsqkfh9sSIJPwwKH2dbqJmQMC8u7z1WNC7bVrRiMFEJ6AL
tmSRKKkOYvewh2oOUsHBxRmk+DBv+q+0f4uVbgZV/Sld7GMdclYa6HEm9B5lwTXZ
gZ7iHBtZ9YIym1ofHjTxYGmTd7XLtzTxS+uVnnVv52267DLDYw18yPOWd+j7RmDM
fhryE6NbU6A1T1sPbtfTmotKizwranSH9953kTSryQgOao1EhZfHtxwRp/wphcy4
ixEy2W1hL+/u+VRtUgDlkPW8u/PVFW6N7pvBf9P5cPNXAl+vgsPedCM9NMjQvAPW
PwzzEKE4MhgNBMKTkz0HP0ovNfS77yP4YWnZrKmCvVQHHUP+T+IUymF5xwPLV5Md
FHG9RAeV2/cnOmvdQ4MJEh9UUQWTzL9hgcjLoi4t0jM8FYX2TSkadt5EVsOZDghy
dg0lFWd2gUQgCJnmaVAbQQUlkWkiAmIzGSTUEJnnyvARBpd2M9UDTxY0xVxCH06U
D3E3DxE6WqVKAVZwUX6VndpGVbnlKXuY06jGRVQuVrCNT3bPk6qyRPwA2uM67tk7
6w8IFdOx/KhWOCrGIT6BJwiTWItrMc1xPFrmFioz2B+0lfAMoPc0WOzTkNGCcEJF
BPC9T51HqsZw0Xgtz2+ZxbNQJOIAzQ7boM2Q2IzFmt0cUohwN9eTuyrQ785TA9TT
wLyvrd7jMxET/xtBKmwAWXxbIxc+YPVSSwJ1dFnxczPnEBHygmal2zPYqd4PJTD/
OVXet8ZLGJStaDQgqwX9xXHB0hkZdo86zOc707UCNwA/c4FBe9AhqiCWcbTKSll/
BgGo2PVAvWRipVnDoIqgnEuSxKlH2got0Ob6ynUM8CSwiHBdkEKu6mYvX6gk/oVG
59xQbqUpt3fU7sxC7S/g2Y8fIERPzFNvcdwgK13okDA6I2NnUfPQvJndItec7lKe
1zcmH+5QZHoQTc+pLkwElQhsPGe5eoahmgatFKHWxdwQY25xEBW/JiPbZS6CD2Ny
VsTNOhcVB5iithAi3DH1do46qu3JWDrLDkz2SqGlrdDVV7hWxTQ5fkU9qZiYRU89
QfcWtCAGsobhikeVge0PZDfKfLYQI7mN97WCYPio0IRmnoXRASxAls4o7u+A2/7L
QYqU3iTeZtbF5nG2vzcmH/1bUPvc+yO08/MxwpY/C5Bf/HIIZVJByutB5Fol4PS5
vYK2GxolDniPHgvycrNXjsYNplPWdWMOfpFuZJfFCna2ykSRjE/BLS8AaK07oYbv
PZxs2fJD4vi4Z2E8nnxHGh4lZ2v4pZCojSR5BkrlQnGjiWgZZVxCJwaFxrgDrTXK
FmVcizeaSVWPrCm6cjnna08Mk7o0znOIZvF7ZRj6DchDwyd+n2eBy9TFRVHjzGvq
pp9J9LR/TX4947n8kY1+E7HhOPrq3KlnfTzD1oHcg07IeVeWRid6lXGXUhdy3aQB
VJFpJUfGpaGccDtatqbAa97zgenskFpoEJUXfCR5yoftEdKeXOGdNtJZb+16QnQf
vg1sjFimApAZG93S/rPkcdXXot7GnzRPJt4c1cuwvdGKfaq6TZvkr6+VJ+0mAAB6
FJ/6F6TZs0GRc4xOGTP2XGuTLiI21oHTZPLOaTJ43VwGtrDEfKWZs3bOCCAyGo7D
Kyf/KUSqTyfJc4XgohBSfMwG+S9a6K705CEd0/At98KheYZMKz+7RhZz41rnGKyC
BBlwmT2cxnPQzl1MIkT4kyQNpv8cYvbrHRp2kjpyJrXfgcBNqSRVEkJtJW5u+wtu
s3FO+tBCpPfgsVCpVG0kKM19H1SLgNtLnKbiZz/z+vLXlN/sk7zD7Jb48gtBrn9L
37cvqSr8mpklBuZmG6xbvJVilObIA7V9M8Iv4OJVRrX134S2c2/K/3QkBpLbBTrG
6LwflPUp6jl+BbG6yc92gXB+LAsTKc9gMbqeqtrYiehXvxnnqREEi4xtymFeJtAR
4Jy/NKpMZ++cbSOv93ZfmKDlR/F7qfA/Ueu/s0wbiPXeRe883zZSuYih2GaABj14
BAe69RRzg13b+xtQihrPP2FfhuKU3TIC75IyGQhUg4j4gvOrc94wGv/+44HQwunt
Qw68dmmhvnnPgwSrmyiG0lsJoiuzcQ7qgDHjt0RMXVAyLzcRcIuuLoWEseKbWzds
X1pZCy6C/1bOYRGPOelG6XvEvbWnoxLrwIIkjIrRs6pF+PRAKZdkbO9D/H95O/+k
vzNIubSsATRp+KNgCbDyRGPiebtTb7ZHpefZqrimECzoRLKVDNTYqBsC1mWs+aD6
TXSMVeMEx2Hiy89ZpQ1jhvQrjC8fqNWEiBl7PZj7Qd04CRcJT9AH7SwTc4EkO9R/
PPzdxF2qTABZGNDUbojLGcZvCDLnHkiELmIHvT6bNn9K3+dadPKRufwLPFIHHj42
cQQug+d3jBCySuFnwrkKXtkHgaa3EnN/sSMO6Deou3ZXl4bpO433wCmdic8GTkkP
s44T+Sjsjpwk1sTKnxNlZoC6Zz2QFNne0AnRisRxOsYraYpmkJ5KmhJuWnNwpvQF
DFeX6Z3lX9VQQs35eAyuWQciuh2ROSpPmZg6L6TOB2zMl0MFKLcrbmUBhaMHjceV
C8VXIEQwf0bxnvicbL86QFS6ZbEsTz4vJWiMUOaixX44uvJ+cCbnYoi88WIP36+P
efJevarzHOZyu4F4sV60s3n915ejXEkgXHhEMj7WEucbufySZncGHn3+zLnlJ45y
NilvygAqPYv9lMr7ytFQhKlBJEoSEuZIdWK9q13sbmNuIZ2aWOy+RyEiHx+TdnvO
l+u/FvEc6i4+R+lHitb1oFJYSaBSLJnLxJEEL6qEuLeWTFjNGptruochJYIuABYV
47bkscmSGxL8v/pQqR9K41xtCuwGvngj70Fs0yAcjCqrM5iSm4MX6h6+sDnOgaS5
q2+tkF12vhBfGgqS3iNcXgjqp6WzPBz905PKPzO1hl5qeYc84upmfqbobgNcb39S
6nMkwbN4qe96GO5BdBinCJmbjs7KbEEcX0CIQFXfzIVPVoMvUtxDi9WZ+AZ2LCp+
pIZv6TwZqZkH6Z3rUfBTAwzo5rqiPgQgk/bOvrnDRl+w2qAEFuetwH/uPqZwzlTp
yX5+djY0Ui4PZHMUVPVXPwPKMIFfwlyObGXjSHtEt6zuw69rR3JnHpl0Pt3vtlm+
OzKIEC/7i8svEKL7umzV/PfbYyQUcgZOUkdJB4yeTRV8y36J8cIrSd8s+DzJjXbN
Ic/VDrmIKVB6p7CdMQ7sgjq53wjio27IXZbrfW6sd5DYctOYWRvm5OjU6TrBN/vR
jY/5bG+xhT/bwXB70TIlKZ363VcLsc4o98GVY0y1lwuoW4KJ5uwOhUYZqNT28xd1
8/2cGLgry/SWl8BrAqSug4os4fkCfi80sHBCtyY/TRXKdoedaSujzV95mR85IomH
HjqikA55GIbbiPcFVbwY3+480hh2HT55LpyxfTCWaIlSJFWcu5RiDHgMVaLYQWrs
WK1zRBgVPPQwRKl9/dqTS8FBqwpZM9NdXfRiwb6/L/992I4gQ0PFpSOIfaaPqrhu
9oY7hLCSMbiV1EQwYHLb4ydnPDeIAIY/Ps0bVnXv5pgrtbynSJFHVcIPHy2564rZ
y11DcvUlqOAA+wIzIFlRgiQTb6XmkSfQCOJUmIYepsPKxNEZQY1Tglk/scXY4fpy
nYWADX8ClWv1JS3X/HozZO6gLkgj8jbDLTyJcKDUSeKbW0KFQodGZivRe/SkOkKW
lEBmDBKTBBrmyxdZGTHiKB2o+uQs9XzgyBN1yb8yPhvj5NWnbIcFCmb77sDwB2T7
EsTW15pVzKb5010VmUXdA8c+42WN8iePtJ/V5q7Q65G0Lh2GHXSEAhe+6ElADb23
ojI27YeCXOjN4a9QFm/8ZJUsYf/zLf4lWobWRezLnPInmoGThPZbONHT+2pyEQCz
Sa8xlJxOPPe3YkGKe3dZ5edNDSec1IoieHu/KxYnAY5FooiHVTGrNk9zXcPhayby
mdhytWHsLgUu8Hj/kjkymoZDtHfJQU1smeFEDMlnQEidRYiDnde1Z6LHA/xARnSZ
q+s/9973kd6E3Vfj9/9vGxEZI3LLg+4xlFbnVDrR7NPlkulTxNm+ymnnX2j4TcUw
FlNhh/e/1yv1b3/LOzUvWBe+Bldifgvwu6w/uL6m25z+XkeE+NvgDEqkK/X3wAxI
FcOscIV1HptNspWnZGi5aayXTotBTrnabkE28eFWTNqfqIE0H8qZ5HO1ZoU0NHm4
JDvOUZf4kqWMNOO5IgZKTB+ne/wMgvJEUPB473g6t3D7JHK2BNdIrHql0Se5Ra5P
+cFqRKESv8q1MMBQW6nzdKTEqSFvn5ZGqOBwSnhMMGoLi+OhPjq6oZeQkdNp2jev
RtbdUUmSFnflrw5o7kygv/57zBvjUubV/nOj1G7CswJqA2QjkYsiXtEbMLdbUy+8
/dTnFoOnMa4GaWhf6gw4j/a2E+xQal+fujHINO8wPAekaU61smOYVZrpjBAmUWVX
gKC9gFQP6LkNLSzWtoPY2M1PQlESEwMRR00Ls1UsISnv9TBYj/AVebgkw877ww+C
zWxHCgVIubqnCVhlfkipeKqA92hEdU9l0a5D8PzK7FtoLTlLfFs2DWAnR0DvdYtr
E4AxsFmAOHEWmoAmgiClhjLUtEiWeMAOuALJbhEG47ILkRy4+aaJ8ckHANyMVx7r
XhbHxusDvMd4/hDGlR/UKqvGKpx2dsrN0FvKPRXnpI9KQI2aywDFNchSpJCznxIW
Ol7GjXBM4ltnLyZH2YLXbHgTavkb5KCUtL+SuRREKpSxKg335z/kOHVXy3LOlXgk
3Hlh5Y+iIbQN34dIJ5D9siTwCMxOMRgcr5kriSAY7Od8pr5sqdr+2zYGO+dDNK1N
ad4N+aUVwbL17uDQeKVYPJCrdvLX4p73xeNsCcGFlD4tDpe0+j21sMTdX/CaaMSm
MvrkJLMeagXJEQ1Yn4G4SLfJvcCmmI+sDQMn7bxI8yIF1SeB5kRTfnIjZj9B/eyl
arQUWLAqfZ8LBeai5To2kPNRj7UkWnFbCsTMupswiq4L883ZoPQaUhWVKOihMa+B
EzKL6/5Bf5RjJz9bi1L8TKfU98pVZ+W8Cr1E2zLnOyL5zFhUf9rp6rpoB1i46eUO
Vkbtz+rF3ii2a4KxeQChKbkdJpa647WZxz4DEFQMg2JE3FmPXzpC2yhiQR2N8Fhv
uU7M+A7HcBj19p6fG6E2wNi5Ql1rGNAh1dNFSDEycwSR0u1mlLsPmSwKPgCzXUCs
gw0Dg0243iFm2butDpcGaWT+V8unj4NmsQ/g07LouhxJESutxm6+sjF2gA7XRi6A
ywLshxjQ5fiLWyci8cLVg4Zj2hjEuqPyplp0CWwhDSFvqnIAd+EnzI4tnVg5WWGW
x88adS8roAuYKLvHf41HjOmtVO2WXu6uoP1b/CXJa2ehNFK6a2gxxB0N/AsAhVH9
TKd2GL6oMmPlE8GRN83eku6cz+q0O4V8XmE+MbbG41ZU7Qc32FWqQenT7M12tclj
XIE4cPTMWWXtHIz/0+KYiKYw+kqE1YhDpk0D4WE7b7KJc4ZjVc+hhJ3d01qC1qI9
cT9zUiAcXFefHEQ5t8hiGXhI44AvZa7HJX/w+M76MWvKj0KTMOCa5q8zIfUvCdy+
BA9bUEusjLS+1jqqfJL3j/fjoekzH2UAJDndGfWgbX+AVhoBVFTv+syYx1Ye1siV
aFc0dPiU8xMptXFtsVNN6yEJml63vONHL+ybqUvbvKWBmDEL1rZj/RwoonoyAKxU
eJeaifof33BWNFnlSk95KowWx7CDNjPATCPUBEBNAxutiGhocomosFMhLze729yr
uE6GPRytJn+Ak612QtG60ofpIAztMW65e/6mZvBx6qHjh1Hr4MmCo8aGXocf0/Cq
3VTNCn4zBPneJiw4jTQTrCcZVm16gRSQ6mrowUnFcyMZiQ0wppi56//czCTolTOD
0fnVpLavCr2vG8jrzlgk4lotfSN9eOSNKQv/X2/s9d+HRNWPLm7pREYAx7k20Wma
VfPdV9VrLymz+ETCxLcImsjOqMqE285WwkGotNz+V9bIEa555g+MoLBplXA0Ourh
BKxttgc3K4Ltz5ND+zbTpV5tQojd/DKEE/y+dqCzspUjzM8vkCcV3ClFg40siJ/H
MnxiJbYTs60cOoLajaJf8uNwWy9xfMwsUPfKKpXLXq1JHD/h2Mx0CVFxbIpqgphR
yVfO4M7MSXxdTcnIJYa4eF98X57BnZ8SKOc7RzG7/OeQtfe6gyUcz/gaQ09+CvMB
Aj5X7Yl3MPWK+uba0rxbYSBxKowKGtZ/aJ4esInR9U5eC51kuNMsHFnBUTkRL0iV
3+Gw2077kSm4avoJmDd3okOQWg80YyFDLgZNwkvcHCbdT8B1FWI+A3PXkMcvrrZD
sHNizBCU+vULZDwkjjwYUf033Sgr8+nfLvhQfa15Z5ONbB5i/W/c02Vb/4s2pHIi
L/FgHgo73KagQot4PhLVPSInsqKgmH9QkdH9DWSq/wuU3ZZ4mT86s4k04E+XvoDQ
+ygISCggxRCjyxa6Jy+EYbBsYuWhHvDgKD8EnRfd1XGTOLVYPENbFpiu5YGKkjGV
3uiFOVPtdPRwFx7TJq6nMguZ6PxN0bGuQKvIR/f8N8tuypZ6a63WHJONA3TPvRg6
Itxaha2UgoG/6cZyPVp4xf0knSh592yRBnb1K7KclLDo5wb8Exd3nHis251ftZIu
3yQ7aUb8Jr9XfMFYo6KWNdWzw4T0Oo25iC9VqV498HyaOi2f8gFCLZ1KB0l5K1Zy
Ltqt9Ks8+5kjqwOCtGFb8ToVLgSSHjiYemWlG5t6aopJ4S53zJq/QgWaX8vi8sYU
TRIA36n1y6X/bj1ulwXg9bZtRdrTeTcFVY8BvHcSbu7upe6MRBWaQDkBbnQOQf98
B9BKU9ZIq5ijUJeMDqHx1UCmAKnwhBHbmSW9eb1GLXAaD/FL9zOTiusstLjH9EUe
eR5VYWQ8nj+Zkf2GqYtSql25G3P3yDBaG4q5sD3xZxfPl+YgvpErLIEvYiyPmT58
y0+nJMIG/La23ie6Ff9WwpV7acP1/yXfwr/PAGuQsXvRWHod/LLJ2vmXVXUAn516
Irv8pSdyIz9cQOloT48EobuEl+GJhp7dbFy8TaE2WhkQHzyv2pLFkBOS+5FimPxa
MEEcocv6AOBOaoxdTh0q8EPIqUEro4EDLWTaxwGR1rd3iPyvx3XnrV2zpgKaJ3wH
zSLCHXhKURxYbPqoA/2zrmtWGUmcMLjFGF7Fls/M6Drm2p5co+76R2k+Gr/1STy7
vO3nYMjtL421d+usyTtmcxqI69En9SP3ZZV7ct/5Fcj9ALN7mbvk/M69Sn64QAJK
PQ8ypMyyXVNDfFTGhXR8ZxTrdWJIXpEAo7h/9FxVR5pKPXhpxQlPj4DyOwb45BKO
HDdOz+cRVHJCMmYK9v2RETvhlXOkxOrpXl5kpEfPqZScRa1Go8dEAnCh2fWYOxY4
rBZEXxp5LRcdzhwKVOoWcf8hMdIsApuybbNfEy7QCnBt7N9oZK+CFH2oLtMbEKK6
egU3xjdNdwtkFPfCaZtWn5B//Mg+GDsYiGnaR07CYn3hFm0KStHvGLkb5Ra4YUL7
Ld9mZU8yykAY+dMvQeUyd3m8IaD/vRf1855YrZq3PRAU/OOjgT4ep6IKzOVm1DWe
7NMdWdaOXUeTZHHkeU/vlw/xG3lxczITGezL8CiFkbpLuqhlYbI21Kw79tDJm0x8
KCoqDXQkYdwHQVlReSJfz8hrOOmW4jOuZDflCBOgjUr88p9nZ5NaiKphycWFnB+9
+ggPGtrUsBWY9Ium0A/wfkxia5K9QXG5Wirs1Bn9iCYEN+WXGIR4k8+LqbBWUKcF
78ZH0qEKybMd90n7f0P3fFVi4ZCaWm2WGKYwmvbtdbk3OQTnhIKJXP6Xr5LB7cj/
H86HOPmHkf0DaZsTMqI0hbSm8j1ZyTHPW0LfBov/aC3qEeMbHgYLXHcydcHooR46
15t7MLu4mOobUfAfj0R07Fejkyfxet6K+g+cfptjTxn5L/FhjlTWB2F8wvB0oSdN
6QkpQ0+AHA07syOUXk5m4N0NWZbDrErmNGs2QVS9efidnBjWuZ2AaRHu+UDe9hs/
mT018MI4QFU6kdJhI6GTTqPGUXjTg7oyGHYDnyVu9ae9pnBtGRq0jqQL9Vzb+HNr
jkNts2dhZFbhU6IMXCo2vSmwPckGhK6LsBfxgYWfa8mGDjv6EkJceLgJO+jzHXee
hPPkWpQyJtFFR3R/Xv38hvnAlmKGpLFqmbUgvsxkSn9jSZ4OKU/mVEnnUyfj5508
llr76IimE88CaHPbLuOigNzVVo26jUQdcjcqm+NP7Go3mflGnsT9jrZx7vAfCycg
0ZoZa+IV3XwetTF4QIxl8hPyIKMo9IfrE9YN13l9BLAdGVXUDC7iHs7sufUA9YXg
4/4/VTWAyIJ4wqRy6qrJ/s0QXqz93DpmjZSvc+lAGng8naa7YOaeQAKyAGkLDAAv
AnEmqauk/00036gdjPGvnl+nxfiNu1Ti0t6q6Mk2KSsKXnsO3VPhluBLxpOtYQgq
rLL0UIcB9feeZvwBjdaluI6lk6mNozUgr7i4aWeB90b8QlEsdMGw7beuCHdgAI9S
bgS5bqjFdi6QLH2RPxD4GfmrjOu6zFfQKzKJqmvM4x958GZHbJM4bMajcAbS5Scc
+HtB7xLvWYDhPrYYveWTfuXDddKJQvvDLGaSSIk+0z2hdiXzodd5/qM6AuBy+jFQ
PTECX7h5xgM83D9t7r3ojuiZJnZOEShh3+FWR3qqfEizMtJshtxXI/zahGI0dO/G
ufy5vz10MaNNoeu94jFxgcamdx0KW6Mf7pWDr5ursqPalgxJz6pAUO/+bgZrTXe/
Vnd1AwmvXAcePaD4RkeTKjyXZw2ttSFGfaOMH3LR//UJ5im2RJLYUHRkqgxkYiKf
4XUXBQREHDqPsyMqAob36TNLstVqiuln3fziJW41HyCZtEAWKQj1fUWgNTaGTWua
Y6kzRAMK9mIxWS70aGMv5zh60Adp55MaM168TuVOAEji2wx3xPBfIm2DLVXUm9qr
t/hIxJ2wcK0lfosWQ0HJfTy6SV1MoM9QEVV1wCqjgcKDpkVAZFJf+2cOhIC+t6CS
voTOg5l3DMlp6qLRr52nM03kIvG5iHqoOmLY557NTv8OJHpARdvm3wYbsnuSh36/
LXqHuMtnqcuJTLHRaV83rvk03KMkQqYiQYVjwPWUm43GTCK7EBLtvttoLpPK7XbR
3kojEgb9VPjzq/nLdiDbFiGL3EjKjFq3PI7II+/JZMP84rzIM+jVH8jLgSM3gEdu
3ZFHtXiuPqFSvhpI386qH0UbhShomAq3yJwgcFaacTsFUOPF6ZDckX1Jir/gYGdm
cdORrKEnABUVLskO22Q6b0WzO+9NGV8A2++XOCyPCc6fZVyHRg+jOEiq+KoCQla2
FwbHAY86Upala51JQZfjeDYh//Xb1dpMCUA2GlMkQpkWo4+9HuTN/qbbUQudNq6h
V0pFVFLEwraqQ6VnoAv+bGVU/mAuSDhHI3EGNIfClkgK+nzOTrWL1mPbe04K9s/7
woVegbywIUdoMrYg3UMeg/z/HxlgBGXAJ/y76B4prkvi4QU7CkRe/jGNpT3LdVnl
JKa+aVAQqs+OcOMyd6YmwQrrZLFzUyNpQZLlUqNBBRe/Op6/ZEpIeH3L74HoyyLe
ozzvmE3mgix3xhJ0l8bhtmdNJI5bY+4E0VOcUcOhj6zbCLt0rBaWo27P0FCbkCdq
NFZijl/CPrNf/WZTe7C6y3PH6MLV7GKqHXH5er74C5usVDpTv3slIDlToCu8gEdX
1TwbaC1UKfQ6sOmLOdEk4jFPgIJmR7EwOTnkq5OIXxsFwbTssmusiUU16WTMvgkL
b2mYHEo33EfwI2lxSnpgdVqsz9+7LkO2FAzu2zt0Cnp6kklG421stcRfSm569Gcb
Alaq/exqrcVkwxNX4aYc2RxhOqVfRMgbaV6IKzs/4KEL1zEg2YabWPmXwlxwdHDt
Dsg4yDgs8cz8VNqxUkB8ATaFbAyPfe3WHm5sjuqfnqZE23HRagRiFONjD4PKmtRF
/U2XrrR3JEuI3x7K/82RQz9QitlTi6s+Xn/jqT+V5jaRiz6SSZwhjliAPmCygOsP
4SVjcDEPjnJRofJzDnGdRxPbGqD0/X09zpcP4LQAfn/uneVidxqw7cnF0MlwNSBB
m8Apsi7FtyfGHmixSiOymT+OHd1QFUquErtRJqZg41eXFgbnHO9NjPnRcgyxhbkw
g6BfiwVKLd+3RpUtIHXkjC+HuPWznBE7UG7pv7T+X7/5MGlRz7bIKZgWsy0qLFBq
a6WfJMBLx5D+CPdCrRwo1feZD0UJ7TEDsUkZ2BjnqBdShI7JF4M6kZg0pJ3J1QIF
S1Zf8ioxBUeUF7ljytMXlt3msmWLjuIH/G7YWy4ULAmSMEs5dGaImaIuf8HmJSAe
aFawab7ohosSGv4Xj8uiCnBiWV6wtq4YY+A+mNBBiybu1Va66KbEKn0eH3BV7C+B
9X8y5USje5dKVOtT2jstydsXz4lgyRFrw9LbKP6aral5BCOAxEV6QR36UkwmkX7O
lfEy3reEZaZleUAvkr/KvgEUM8p+IsVrXgsKrEkqhivQck4UkYX78XselGFnUwfb
43xzIgnNYOE4euoUoWH5qTsWQMxnllsqv70hzDFfBVOMyKlKDGf44TyvgunoSSLG
l/2l21iTvc9M+JYEp3Z98m5rX+ktIsxpVI3uWX8/i0sEgxAhmzB6ZNEX7Ukl14m+
0IXatE6O2LsJA9sqGMadwJSk6IBQzV8xiV7tr+KvkKFM1e8WopM/inKQYFlDSRmU
i0TmzArwM56M5fvmLrliMZLoK5ZKfaXyW0fN/IZF6Xop9yW7AoTB6JZ+WHdiIAao
a2Ae/CI7Gei2UfyzPnNOGfwVTqV46EfbSpXAkrzuLFxhrk1NK54vQxFObIS6nNFE
tzhIZiiykb6u9D3jU+xFxwlqb1ApdkpL8UTWC6i9ByrUAd6ySbU0ym5RnNrbsufw
PIuhHJzKvFupu2pIA2A3msqv0Wn0JTTDlPlYhJ+5vhqd3A3+Ho8RjcMQAKAbQvgu
4hXQE6dQyBu+nFJ3FHGOmf4WxqP3FzYczSkbyWSKAxT0QSzypbU1YuO0GDS1ZTei
f+9K7jaNoH4THmYjxf4xmQOAp3WGmK/ZbYcwxdNeBwTkme9lkLfgqse8euD5A/+p
IP+BB7rP55mDuKi1xmlfwQW9xvtbXnUUo7cTrtRFoyo+hTwlntXfS8HRuJUaN0L7
OIYc10p1pzUc3/5b84wMqqATCXy8RupmgO/hf1sR63WCgxI7lQdZcFwtnVDtyYO4
TBBDDR0AhO49Nyb48k3Y+V1w0/hrkL5j1RZvioBws4lEje074SXUVDqcHPb2EjV6
AzGA16cPW9C4KTvDtnxy9GrrHMscGEfdr0qxniwldesGSIbVSdtztq/ZWKtMSivo
cXT3ApRUoe8ifbJgoIzXwJ1JQzWJR8DB3M70dxR/pIJB3SdOY0UGYbRv6MdaF97C
MU5h3MitE6CDkh0OKf5CECu+UvP0z2ao7sV0ityoL93/gYZM/4OqeyoluOJwlwu4
3OoCDHNqTNuM6Ks/XEAd26mg4vBJW/CSsIUxwC/HZO2gBjXFViow/Wcr1fxykqa7
NBRwINxq1smnCxKMDO/cUMgfDQbbl9nziyxaNphe3+VHquk9bS4waUls2BNB0Qpj
FjeNTJ1PteuW0t/2dt3XVQRI64Ab6JnQGfoIkgE6mQZMi0QM8o2S1S2/IONbiO+U
bVej06nLszVZWAhHwuPyaFSAWg+4Pgz21wsl3cFDyEbujhlkw+CGgbyqFXLi5ORm
kdtpxoxyRsccDEL4bqHBDHP76ZiIahRmqMwWa/DpusFwiQMdaZtfENjn3K0AhKO2
fdjSNdodKIPFp3xr3G7K9I/HRhHBGBIHA/hXjr2d08UcKGgsqflNCf3iarLF9zP1
2uvpXSeEi/CDvmbq8Kpp981srlIp3zQdHXGYJhPBXfPXT7RIdtcUvCGm2vy9CMux
2LBK84/+74ORwIcZEsk/onqbCBSJv9ToWXu4QsZzQfBLHQGyZLFVxvPuI8evjktI
p++4i8Xr9w7fVtw1wsN6Goxyv8qVi/A6pmN/vLdYFl7g1QwL6g/8RR+yGG4xKBsz
oggC0A0Fq+HbnNc/2lYbJlkinRClrRTLOaG7jNFUYeyu6c8Tire6i/g5L3hmWT63
jXlF1RrHc42EAh25LWy90+StF3Egz3pzWgJqfbYm/vnhas62KJSY48/7pS7uwqsF
03fFvoAJBGvI+boIyge4Z5RqoqivLvHcGL7YAxRPUAEvR/ALwlNx751QZzOSGypp
hlHU3YmXk2uqXLqcXxCP7gd64aRY6qJqrOwaFXciVLfHfgaSF0OoYiEt9wBWQxrS
Sw/yrCAgxIR/1ci04duHkTbxYHWWVv2ovLRt1t5w75cFJnGQ9GoHllM29L7gTY1C
0PzKuVSaWurY5pIl2Cj4Yk5RG6TFetUdGq/QrlvEdqjzFfuVvoUi5dA50Ph1+UHn
LaD8c0oD0CH6OZg5hLP199MsEfOwzAOf6e7pB62fShBiPIjaL9y+ZjK++b38jEQR
V+hpVR88x4Jdbf9gYEchxuqC7O/YnKu/J31Wg8CIBEh4pdyT5Nkt7dNjU/MxQO4T
wYbqgjN4BqgagAjINiY118071OSYEFaLURyiDR6892FAjHstCd3Ny7ekpXLuqjKb
Q9TcRv4fxiuDtbgVIQIncXbHVcpbADt+fLu3CyQ0tFZ7iyKLRcf9oUrdNWYwSLFe
saFbLimNiCIf08bczq4oROzeKvYafxMljzl9ngS5E8Bcj0ETEgTsZ2rvnIsC5olH
3uwfiBTIy4oguzO9USg4ncdy8QBAHpS1v27pjJgu1QJaMBPagfqYiHjPS9j1++uI
Oz8jlKRs7UANeFAcpMgrd2ZYHnnELAOIRRLq4hDti22hKRWCgs2xhlIczpUflvaC
V9bEon8fbuWAKqoYsvjnAd/ZvO3YplZBZi4Rzo+73OaDE7jRQImAXEGOn7neKQEp
LUErEpG0WeGUyjc9ZOOIWXawf+oExnWDM6jvQ4BRm3+1/NefcFen44CJ5VtzxPQm
fTlpsJEvpETbCrE9NQd0vEZhhPat+symDbgeieMB78AbZ7yredNlWkLAayLdXsjw
1fRkQh5iWUXq70xYb3cW/5tXwb1zJhkSPyF5si4rc+aAz5DE1HrxMn+Hz5KR8Ktc
qqpjdkH5ayG6/BLJQDrM7K7AVkNFlbJAuh/bPp1qL7s2hlwDzQhq/Rh3xftnnZtP
QdrNqLUOQyyEmYBkl3cvwa2dDwsw2XLVvSloso1Eaix1lnrb8moDrG2ScyczTIcw
7ufu+0xhr4Vr3+qNWqwJsZElOpBazgK/sEn3VhOmD3OT+6vlZzamH8wZcyftfrd/
MMp68lNlyhcIphkKd8a6he1ynFnc8HwIwxrO74m2tHLQVGkVWfWZefL3JimhD9ew
ghlTKHJbVJ4nF5Q/W2msuyvLYVkihuDDRXDJC63Y7yKQvib0lsYBBucJekCEyOjt
twmZcA7LLdpB+z7PBTaMJ2Bzb6AXyoaZqpyOSsLjpMeGGw1ZXq4ft5XxEQ8KUNtR
5GQzl/G7/88cw4ZPNBNqM36svvSQTd0o339kP5rEMPIoQQk//Shc4OYrwokpyIAB
Ely/g+ySDVUUhwkty0cv3mjhplImx+4Jswv4HesqzqY4jF11qwayoCqZhKagKxis
8W0T7YqWysZfZmL78BiEU/4qnVuiKHsXbXjRPTgEF00kgjr6roL/oGjXsGJ5IXNJ
26vPKZryxlMvPFh1zYTiYVhwyZ5VWdCXkUJjjpP+toKh/b0dxYRd+26L17Kb0qew
Q1UcQYF3fZurZCDb/xDjIKwkd7VF9Jy4qDXfD2QGp9ehZOkrj86SCxldo3Y809A4
/fptTvK/N+Kh4nn8au4zhqzjfr0lu6JLEgvxC0y3CGUhvTnOi/kKiomUs/vvnWP1
RiE/DaSVUPRAb1C/W6Uo7FFxFXZIYPfSAiFg7m9ZVvZ31AqukUeusFID6+VvE9Z5
N+q8DsPUhM7ar+6OzCMHwGt0RH/zjTu1YvCwG645ZtOGviK5b96vufOWDhGHLjED
uSZMtu95SCbyMkHF5HUmX7EufPyoo9LKFExRM0Jgpsa/LrjE0x/uuZH26zkRWu7+
j1qhvJ7Rg3kf18oPWkMmZpDwcvYbRnfwVinevRIdJiYD+QhQq/1GMFdWGo+bFR7O
0N464u0JnYf/+tPk9BnBT8Yp0oUNffj6FhogYSTFp4gXCpqq1jzTrP5FwNuNkrvI
m1VSZKMLupY7FV3BYgnpNZOelH6hLJWtwQFMvh/VX6ZuB8264e9I5JxENfwia9tu
7S3JKzBfnCD/c7PXQ5zKgmkaC9SaAKjrCByIUCu85eTfRFbUw+OUfuCFoJz90HfO
AIXcbDaxl5a72WAZPssDLFCZ8K6nuG8WujF+BeN5y5wqLWTb0wU9rr3e7ovTT9kQ
el4vN1psO4N4TNbF0JHlBYwSm2QNhy7TTWhV5vJF0WYykEa8PFwtkwn5JPotk71C
2CtXU9+G6znum0RSVFFBQ5zQAW2WTnHZ53TI74Tu5toQBNi9WTzHrI8DszGFbgwt
03Up9d2bIdsxe2KSSPH70fFzuCpbmI5jZovYtho1OskFfDWfqoVokWZhmcVZl93U
GX4OiFR11Vzq/atO96hiZqTvu+0z9bJ3VDg0smyTSFGDKJQvd+0jvdyFzi9wPaOj
OXBPnhCWZK8UXVRv5ONH/2txe9f3vW+gxiKKoXQAMn9vWCu2dBiw8Fyp9m3B69tm
aXTDG03/0NU68DIfntmxyrgPETYY/q8/pLSNaWftdHQtkOgMW5YG6QDwZdPHdCTN
WixzPZmcs20Q8PZSkAOxqWWpa6TuqRBjMigSy20rX7RSf1z+pLqfVlecO9QJwzCU
xcjI80uLBJIjPKemCT+vKLjlbPKxfjKL0sEDTN15qNhp9JSyKH/0A1y/wGRHVORR
o2JK+hKVutIha+imLlXym0ZlSb40CkvpLb/tsYqZM3CSlUgCEQ+7nOPm/erNMFnG
6b6sg2Srk6jdkR6jRsDEiiidoHaDnna9pLwdXOg6ExeqFum4YA0STU66sBE0rdad
pbDGtpaC15bYQqYON+X+f+QOQHaQmPcFHYBNpZdaddCRsLY1YCkeJQcd+009IZXi
57rXpht3/NxH5mC4HFhdRaV13PLyIwSf6G7eV98Qu0JACFeuLwHS7vUGKK1WstsD
xG7U6ImjjK61q6CTALcQ9jGM+m0+bsGjfo87n0AgG7akl2kG8NhBr00fDKx9Crdf
SXeHsKV6svKsXqAXlKtD/rs+vMENXCoeOEKPAEFru3/ErGoY/IwfOPxWXETWSpEN
o5nh0Dz8R09cJ8o9OOZAdqknwm9qoOOc5U7Hwz+lMz+JzM6kvkFKDI9e5GdsmoSx
CB+SuUy5kMmgLHCxLn2L9bILbxxYTGcc3GbpoJqDR5BIGYX+89c3r+WcDQzILc0z
IipQPfqv4DJF95UCZG/C0duyaiRDzY9v9DbiNE0uw6mx0a19uArdZM6MCd40OX7A
nn5nEIj5AchtqwivnRnrPQfaKTaQxK4OWw65JDQsBD3r4yAGC0b6bjgHmDiqVYSw
M80V2RtNfPIcATVywq3eWv9QmVPLxc8NfSidcXK4H1uR39Hk2T8SDJ3G8ncEIxmu
USkR2suCD5BrGGv65eJEVMkNPV7ynuG5MPDDXq308aTPkYurUm90iJ3wWSzOoWJm
XT7aHCiOYlsXV6U/y3PajC8qU3M4VSAfxCImtHTp3x58u4oxzK+pvlMblcEkWwyh
a06dZnR0AFfgNcmTdf3YywlrWMUlLThLRWSu9V1mAxckUjA1aLLwovg4aUZpd34L
3meK43DQeIrxD5IqesXWFKVLEA1dHUWSvBAv1zNaAL7nkJoD6sfOCfGK7KNsgaUS
qRZW5PPQV1/y/69MMPYLw9bHFKJ8FN4TQvJHZlkP68AD3NqRJp/QLN2qfwSyBmVU
1h6vGvgQy627UGACQ5B3GQHe2hXsonISNHuDfKcIu7xxpk2uu9AHbybLTD8Txgko
gWoRfNRmMlk6RPFsQE+Jz/OX1rUh/YXajHpn+ULTSYvZbefAvhVUxA+IpzgA6lCk
OiaB45MG4VI/vh8Au/Ki1PSypGPQskvVbwJs1VoArKJ4p3LXIHFg25PRJedN9zOA
DIl6s6KOtWJVlb84IHiYleQhNhHnwifss16zH3TXyjPSnMQAo2/wJ5qR6WFwc/rT
U0Xn4hhSRZh8yFGai/32yachyZiChIP1yY/eMPcAsJua/59dT4+PxWiRmBMk7Tvv
5AV0kBxo/WUgAQioCJHYD5oKOdggRuuSJOtNzVC81jcs/dUOKdFlxhLt/QX451xi
nSFSI5Flz2v08aZO8cel9bOljGECfki942eopBe+VJU65LxytI7QkgXIsbC1+dFv
lRD2qwn/zsWAf845ASBtjlFno2OU4dfq1kP4LkYY4IOCUa64CjRwnIaPf2tn2sJY
HvecUsyy4blQncpHAIFOFSB5Y7+f7s2/0i2hL5rWI1RoO+BJwMHRa84n6oEZuZAV
GSWUgFMXfO/aMetMC+us263EtSI/tSRyi7UGao8FtLu+Zs5PzJCwuBTNJDTjrmcL
P3WrGzByK+MHONYu4yLxQIxbpvW3vx11ej2t77wkXA+T2sGKWeP54Z5GKLlrUuWU
Isn1NyxVnuvxW7AKbPuABISP1ypaqqZeheexv75eYSWvocrGsdvAKgmXkD5lO/Se
6rM4G1K9LWnFwLS3mgImmiNcSLzaLBx+9DarcJY7KTOIbVOhqNC6BPOyX+156SL0
3UkwYKdtk7omhxcdPea8mszKhfZnsNBs9B+jrz/MGT3GfgoJTAy/xHX9zb7jPXs+
8hXd2/t2XNS/j7lBCB4+NKIRxkEKKArUTuT+y0R2lCZeLveOdz+SwbRYo0iL2KYk
oXwltAbZjRjwfspNNt3kSF0x4uPkpe9jVmUKOeNXXRO/k3WdUemK8sQEWqqwGfa5
hKAQd3RAmL65sbUFtCv9iu7dly/zCTuYJCADrMrI8pwcrwOhcW0gc+iZRcgWAQUY
Rwnyhhl7oh+4/4yPsNXrjnXVMIddbGUTXIUu+PUS21phjtoUpi3xgW/CyYrAjgPe
tNEftBAv3XV9UDtDYBP/07ChbTxg6g1+ilk2eG1S1arbREP325yCX0n9g/COFdzq
mBmM4qWFWlQNgqU1//UIwVWYOoi+/+ZF6x9sAszIce34VaMWH5CP6W0Qg05MUjP3
nMDkIx/duY+Iz1J8qWHzgXc2QmR0F/yIOfFlts08Pu5mxKeofNANi4sGRddutJcB
WbaKH1OB1NqjMJ1jIk7OIpe2P1yhbVaag7xj2pqNnruTNbF2Exqnwm46bSu/Z50M
dh2gRtgyeHJM6hX8PMUbbsU6Y1nXf3wUV+ej20wWJJ0yElD3SgIlYCaVLShyRBNy
bP1lbFz8acPs5SqSBqmIOJZOQnma0Q2qPUx1eiR4269SDQpDxi+TyTaqc4ufm3zy
RPGqtMWa+JzByubvJKdl/M0mckUz4kJHt012E4t+w5n9dpuH8TJA8ZN2tdGZcF+1
xJfCptNwbq2w7NMhWnpQERrqmzAd9vyE3QzYCsZTdpC8w4PRgkGgf0zzTcaFlhrX
Yx6NDib9IfR25bKrUDFz8W4l22nLZgV7fGGPkaycG+lsijmR7/4J2sPLRp1t0Ve8
TMS5LHyk2YwRJxocBIqnNCzk/ZA8IXOjxf3euG54gBaYbEcYbeMXOQD9sBn/f8S8
FQ8B2zR4cTq6cUJUlN98CerVWcdS62YTzDzMaVkGj1+08xDWQtmfkTJqDK90bJtz
fsfCkApdDwln6Aaq+dy3RdqSRgcKOPcr1Ep3u9ydh7UsApukAdhQRl5WYuWgUQnP
66DwXLEgeyL42FO1c2zqTp6jdhYZsjS1tQu7C31pSWQ6FQkVioHMSyTP5FSflsGl
DTKlgprwZ4jRDtM12Ypq60iji6at6ri1j0KlRcojNcy52i1aqODj8pz9FbLi3u9X
AIMz715IYz7Og3ceQH++OXDFMMUmiPa4IUxq56cOeaHVIiPBZp0SWwKiJuwsiuYL
890B9UdxMLg47whS6R6AMEELnDJ2yMpGrmkxP48hrksazDPCa1ri42sIJejw94xu
KaxL3dJr0aATZ5VOhihXz8Q0fcYzPOTNovPkBugFCTufUfPAgOFswVpgEBz/NnbR
AKhcDY1n0be7kzpgjoYH7uIHfuYuo1g+1+Sx8JkdKKkLGw+THLbKWMtPOz+RqQV/
v/xCBwQYleCJxNFiV1/yJsTRmI/STYDWW+Kf2Ix8fRZuAvZQEF/wNYnEOxLbQB26
be3gvODUidOmh0z0zApBRFrWqUMCmtAkORAqTzQ9FG+NSed062JCIuOEoEoy0bZg
ZRSw1d495L/4e96m8YuQf6yMt0MezxyaCestrHvvFlls80VkiMHmVfwxZNiVceDh
TQGihiltK9cZh0Rb2U5qFvXJTRCNFu2arO1NJLVR9mQ5m1FBXcOtJEjmJ08ANLe7
CUvBNxOFdlau7szZlMtLy7/xqYrcUbFk7oWDYyd0WanhkJKSZmgifcCdhWk61C+P
Jd63Mi7+i8SAPuAjVhKNqLyI1VTEqRBr3GicrkCoBGQpB6L/jR03yT0ZI5UEZnc6
DuCKoNkGwElGY5r+sC/RDmFAWIt+sVD8JLFws+MTlL3844BQQLXyemKDfWYAL9AY
LHAHdODloxcGdzanvlnJ6YpKOc3WvlXy1ULmE6DAo1sFP7/vS7KYhAQBR2KDpvFe
vPLVXIDzKZmuUCwzmgvymAUfJEBwJ9e7xkKQnTJQrIItPEklKiLD3I7DXhOrNrzx
+8vuKenPk7vn130iEyw2cjo0HLy8sPdxTIAHwKkvUeoUQGenfW0If+lb3CldP8AF
0TziRvAjxuoUFbXP492ljJtCBXic+90arnwjMsZVF2oyohu2gIsfRmPPYrwcjv9k
bPs9yIZazOxxSLYdi4cKsllXY1njT0wCej4HZC7zBQ9GE+hc1R4gVf4kZoudOS/n
QDWZlMh1sKZ0H6fqByqNr6vFfpfHP2/oDbsem51Nwma4FvgXWz7oOPcL3iN8FvvO
jPbmPTf3kDQfYLnqAnUzkRFaZOyb0E9nASuOJElLHwyVcGNusWzbQIlGQpmRnL1Q
ig+1nbgpg39eFrGsKpKYC7BroHOLRY8cphzRoReff0LyWlwfHN1SC6EYLu3Q3V3T
Vaci/KCDpo14Y7485wVqnf5FNCpboZ4CVYe0SNtFXdyatuMMak7nhhCh1EXF276l
O3NZnOXKz1GAaOpsCdrgRvdPiNhnUSgZTSP9dH2FdMraV6A1YmOFRSnLsAeiQOh5
vIECi1DcuKTd2uo/Jx6lSQXsqphlr2gFlHP/ZImwU4si7Y9EMyE88B5ear4iAX9L
HS/izr5JxHg3aucdhJ5Bf4GAey2ZAsjhr8oI1ip24fUt5X2HFBJCVt8Ror1rNbtb
th4n8cwsojnBlHZAK/OJa+1JaN8jkBu1l4ckpqtdQB253ScBXkeDdZM8HLkEV+bB
5nEFBzVbIz9wj7focTJz1AnBsMioJusaF60l+zmINmbg7Set7dsZ+p7K2MWmUvDj
53mqk5ZxMx06vH0d6OQHMZPGjWALcTtgwIS3jU4y/B+VqYft9MmsimEj3oyR8X3z
MM4mc+CK5i0UGA4E+7spV15Pk9/GFZ52k+KEfmRbsRMnvyzBOgnF9oTM74SUsTrK
CB2DY7LonyYCy58YJRfcNz2GZgywIY+2AAdsVGEgCgFOT5LP+G5c4A6SCVOmp0hw
CMYt0ytl49t/bycSFOgcMFpNNPszBcA+d55KsmaCl5z8E0XEr60ot3pmIrpYX9Ay
tt4dFPMA+Y7cN+K8/9nUz4tIM8Dun/rR8XUlNZgbpYCE4c53ca3it7iWCiyVL25o
ZRmHQmiHWsIDTkCVng7MnHGb7SsdWc55SPYqNrhglMD5pIVxXfmKDpx4uqc9ijt0
rISPBJNsqxDwlw9yQEYKjKZr3KUx5qf5qlpi0tpTONJ/C19hlYMPOL0Vmf8pE6aw
ZG/hdK+xI/GrA4X1t3YzeTlwDH8nf3O3v/y1khln5/9fNkeILh9V/oABUAg5+Af0
g4VaLS/6iut+Md5SJOLGK2g/4qw5JKF/MEV4y/Hy/jWA+wo4CNI9jUexJGNxBCI6
s0gewFWZiPO7oJABR0ZcLsHtrxFsqPIah8kcStHRKAxPOXHfOxhtO5wabOHPk+yq
h8UROmW4Pu5aBl3bv6ZFjp13Ts6jSRlGa+FgTlNHBn8UG5TVkeuAfOjh/uI5nWkp
CG6o8K/dh7zVF9un6CYQyfTsy4xYPie0FIqs8Gife2zb8SmbzRZ/9iIalN3y0DgB
4VJvt1GjGRzV5zPdKoTjLuk3AOU5dHeTu7tw+RuCOsXEekHb41DDVCfoG7fRB71r
ffpelLeZNGwZHI1AZIgRJ+qx3frRoNji4c48XdvTdz+CR07PlorsFoiTHPG9MkNx
IU1gzoG+OzLjt7HVutDYz0WJol3244qPjTFSOsuX8ptyu/flDEbt6SXVhCPqYLRs
F+Ib+kwZsK7ruVoeOPgdoKdLzFkutSBnwMHLNLamthcpJ/ehrdZzFM5hboL38yXb
+wR0dgM1w898UKNOa6Lnan/g801rJSln2A49HwsiZlEYZ15bzE1UJ57bkAfAZuJ1
r+fnZLJ3gdUSBOXbhRvPRBoNmXswOUtXoHL9wJxGpA/iqJFWWOlPmJPG6OHWCOUu
umpDT5gHSX31UFIGGUdr97DZnxrb+5Z6+oMwgvBtJusjUbljH0uISOLmps0dvoQA
cblUCjepM/zrEGPC6r0sB52xtuJGd6TkBh6dVJxZB4ESVZo5i9nP476nmIiL/nEL
kX/qsLCSLyXNs8IG0mF5KGVIwI6hBWRnm0GgTPizThaCuqmU7q3EFUFpRB4mNkkN
pPSNHVp5pFBg47Kz3KlaR2N4Hg56pl6/zybpURLjw6wcwqniTReuVmRPXf0SG3EP
6cL5T8ejZ+C+OUI5+kIlTDkQ2i/43aZuntyjnVQMYPURGN9XUkfS6GzL0IWRXVyu
qUU22wfBUBFOTuJ0bcAxDmgp1TJOGebD0dNIsepmfvE9q7JE0EwqY5mBRYrI256+
nLI4n0qqq1GyBxY9uzTzj5DMOBfWVbfufpwvqCvQ1yBY1EXv9134ICu6okmsCWko
jShPkjFQcUJtiQAXoHqHxqych0FwK7FKztQItP7BnZiDODJ4j0CSyf9dtAhBnIun
iThUKW7GIqtmcDepOy36gBGoat60GMl5c4mekvHEXIOte7ghEOSMcgi9zQueWfCm
1iPqFFm64PDtqe7B4Vw7RCj08QYJhjcsGhaApCkIyx8o7PYpZtlOQPaHpyP7luku
hHnjNZyJMihCppfkVcj14EctauyaxYdi6DIY0HpSBlv+GmeLSu6fT84OBzo1IzIS
evK5IBEFNfvSWZMlROj0TBpc3lyfqPXU6vNhA9lS4t4SfogfH/qM+ikwR41AEI+c
KpX1ool8klrWSoTue1oczcl6d/VkC+f5p0fIV9Iwn+wB/qe8hdfZC6zdAAqNj0ZL
vegmZedVTE5wUGvYHflODpXGIu5qwDsKEG+ZQG/jwo0+SxGejdUdGrvRuZYe/2zV
kRWahf++5ME341GMeV6jjfwqrY20GI9WLN/cIWwP3Qh3d/k0OAwMC4EVbauyYaEx
t5fkmlwzvYkFkAhpD4Hefr6MsLV+IjKeeaBQy1q1ye6FdYb4kKsPlKWqqiO7eCTw
k1NtEscTuMXkBebQN+oe/fY9fHt0TBeF8h5PRCT2F7b0f1ZJfsF/sb1ZUpjNslyD
bp9zpWJZq+ex6aOdqTt8SMTF5aM0sbeuAhCRITwOX8qdKaFjgBn8ySJncDmSnnyZ
2yHmhWUCprLicViyxi2QPnqkDWRrgUKGCseu9NS44Rcae09qayq14+dCEzK4hvNF
Misqvk+LqvL5LtT0sEymn6SywWRco0+NFIAPO1pqJ09jLWtY9/sILi3MRTXaAS3b
ZIBiA8xlhyC3RrFZyf9c8DmNXA7aRCFJNcApEGii5BO6K7OWrR6oKC5cAU7Lqt5V
iCXOW7Y2ntFQAj/q9lc+fmF/MfDVBw0fR7iDX6/WoPJ6rU6RFA7VEwNuxrTdCTCK
SAfcKUOOkgLtA5tvY8cUZnjnhRJpr81BSsjuAVe8dplXqn4IRa4LxSsdspNwva4Z
tClTzjMp3HwkDfxVOlvgS/tJ+6k/Qje/G0QINv5/wdjeKwvaRe1ofYKcsT6slGSn
+I622LF1nqEmp92jaGyBpKe1Lasbnx7C4RiDLGEo0g6iuYop9iVCLHLmu5Vc+AVc
bXRrhS+JKFP8gjur1loalZf/ENcpX14s5WvyirLpiWilupeLRc5G/7NDTWwJF3nw
Av2kUPeUQVMfp+rgLwrq7ynKirFCGfbiQKjQLZsrr2xk1O4gK+C7dUvwziM0kyTP
pOh2pWM7WTg37LpGGAd1Pfzwybb8tx+R/N+jVNkwbL8mAmvnqkhqRynhRNn2e+T/
pYAV3SMABov68qRpXuA1oe/xFKqjHTWhLiYVyKEYJMu73M+04aWDuMCjX1ugE2v7
yEgxa3zNPEGiLl0fbZ1o+ZG27ibNOlE27gi4BMsSqMI+E3u8Idc2kv6g3ENnuefO
j1fH4W4IemmJrVF7ejrWxhMaNrjuVN9g/D2CveQVHkJyp3w1st9HkmVKkfpsp/tT
BvRzjtwDkbTj6WfFtDCkqfDexCjWsNno6Zt2st2FiNRLWjP5gylvsJ2t04EKntO8
jWQaJFw+6NfrXCVymU7Y9bffwID7A3Wv+5shxO3mWifEe0b2vZ3ZFS8iqLAV/Hqj
HaH1PKWzE4EP2Hnc3EXWQy89MtBUq0cBwiBjd+1FE8/PwufAu6B48bCDvExMh02K
1SlydHmHWB3gumeEaTRtk3fwA3pjKzxXgSq8Qb8hXb/jW82ZptE3zjwmVdPKj6GH
EJ+wrhNWpXoqD0sG8F4ox0MjfgeCYe8TGUByNk/lQ1KiGQkiaocS95L1yuzDUc3F
MNQzz98EpeQW2XDqiCq9lY5lLBRtDufnYy0eeGfs4ZK4YEu1WufgObqxMuBZbrnO
hwNB+k52tkWkNWH9BB3xPNE0KiSWd9w1l17T2UZ7j78YGrJ2u64h5b0pM4MF25V6
AfeQStMGHeBGsQiLwWHF77/ObAPls+5qr9UV+31tE7RPxK+Kp/yjmHN8/LnN0odh
hC7iGJQnTUTsAnQ3rN1viVuFy2d8SYN6sNrmXUjC84VicuogllE559jbdR9EGmDz
JOft+obYCLdmpnY35m4G8e8qkc5LZBLvhv531udnYNvZzE3UALhH52I2zLjX+J/6
SWAvXZPl74cBcJDSFOwnEKC7GjmbJqEuSbjTtsIRQYMGDQJ5zQhed9Wo3J9gE3H0
0X7ZUJVpeETMNQKisXx4c7QNU/8+fDMCnWiHsLq07Ma4w6tUbim3hA8V0zVNdjKr
2Aw+hF6XzbPw4Yg/fLb56s8X8p4RbFkDl9a0WvWlDhOmHo5VcM3Rlr4J5lvIMbcC
/E8j7Ck3A0AcCOUenW2Rx6eGJWBUhb+oSCr3dX37C6gi6QB6QhtfzcQOFH5xMWXK
K7dZV6pygXyYaad9RGQByQH9juX5NNMGB1RjWzm2UxcPAH33oDewrL0Rv7yeZZh+
YOJiF6tpGj76vCzl232LfB99uRxOO6W/c3GFyKgs/aSCfdratzzi0mhXjY7yuhT+
sMXBpAJEds0QHMwT6EbC9aEBw0zUnqczXzCitKS4v2VACxSbS3zEjtMzEmdk78Of
Hs1MZZSZUVAH6fgJjvC0e5+lh0fr/NJskRgUO6fMx9+Ks5A/Lh736Dy1ZVWFHhfb
DvTHcm28F8ChBrAsHC1LTZ+ukVUqi6GQb74hhF41pgF6rcAI1xzvz13n5J/zTWAn
gtXZUsly9ELV/zlpDBl96BEZEgKP1yujLTaeQEmZBMV/ou+LkqU2nB12q6fdQzCF
7o3MdWNbAo1rFZ24G48+rau3SbuNXEHehVkIZDvOhgREu40eKnuM2wNh61Zi8L11
hfj7U9mQLHLBXg6OyDvP0giAhUfWNsFpCV8r8fRw7+GQ/9bB6XPumrY8KTphlUAx
N2hXu/3cfAeGb5ONstKnU7mHa1xAuGAhG1QQeVsnYTlwjXAkiUWqbYGW2sFy/3nz
Qh9GDVDNZ2fWoGOMZs9RUUQQ9WBVLJH+kw+MfKGo0HdY9qRY1sQG76rjKwNS3hsv
05vd5VFaogz+gz6Mloytx7F3/2Byq32m0QDkTzyZ+TFnzhcOhyg1ruA/uExHjNt6
wB7onQ6ssssIfPkHNNrvtToOCbYRcjFD8Ob2p7dBpb8Bc+FDoHyuHtNs115jfNQz
kbN5qaf49Gs4ufEppdjiS93qiLwvm++H4HVA0a4Q+WGaYw32ZvsN3zpDCizDk8M7
QDNWuTG1GXYaCJa/Xbs7rARcfLDqMNPFqCUQmC6SA935y74q/55yHOTIfJAuCIyK
lJnL8W/pOPBhROWd9qBYQHSYqdyJrkh5ZjOnDpcMlYeOrUY6oOqx7R65+y9jVNA2
uxPWEQXzuolA9uhqqZNIomXsLLKkVfkVOZy5gWcLBJr5eKxPT37Nci3zSEhcwWIT
FBBedhKuiMNUmWptUyQ0Kr0I+or2uGrQ/Vd75bwP+j+GDP1jYGD0IFHo0CMDsKtm
2kizSWTYOLtqU1x5bLflWS6x4p5YUs+tqaZmPiIcJpoaaz5O4s6h1e1iAXVFqVaN
KTnD76eEqKfB2ogflSsRbQzEvo9gaclfVLvsPMRCbTwr9rh7C3aOA4ah0C0W06dP
v2w3sFuyFbwmWSp4Tn9Pu6ATLCr2UEiakWIYBhTYR61u7+g1bufVTTaEEeSTRvMP
yWy5cR70Q5AS5NZnG/SKdYeVOMMZFYu1pw0lyQru/LJnVpRrRriVZM+aUcz9VjLZ
AJ6PPZCwcqrdbiZBXreiX1HAvQWHrHILeT6LZ2/LGs2ryEsk7oDCKo5yt0TpQ9FM
dqSUOvG1YFLRT5ZzBaZiGjdpc/js7Ywniojzx9b1si+twnDIh6vbjlohDzZG8CxC
rznzyzRLngdwduxjxBSgoQfx+iZ8iSoYPW+9WBu6bs6Xrx8LqOa6LpdgxfiqCmFB
gaoGEm/eH4E29fTSxRMc08sE5DSjlgOh/CU+XfIC4xpoEiAStNMO+9Phy9RQqYwR
y3ktUGjMuX0TwQMBauW8h6R8JPB3rssufvcUb0Ocn9izKdsVtT0jlyPAscVi1T8/
gTAGmUWe4CsEw+/iVp67OjkJ4sq9l8uJVVKi5kIaNGdFo9z+yUxhNTwQB7oiS9ZW
CgCwog5fSEoLnMHEGgJ6P5iN3KD6ypsv627PLQkDHpWfPfOdrNvb9HEiJ18ERkGO
3gBeVsV3q2jSeSI+1s8IPN1uzELyAG9ylkfvKWYV7ct+24TvT5HlYayhCAa+H9xp
sotRgRjFtd5WsmQyfXcD+MwbKsD5mmNqz2Y147/1yCPBZJhCDdsSXcFnwsFV29o9
FUwrxAU4GWfjcpuSbFJuGT7eYU2VHSMnkIfQ9Llgy+AaaLBhisjK8rYAjjasak2q
qJefQzVDcBqGn/+DnivEKsA/AWubKmQUxP6PjG2UA0hSvM9X9DKbOwXFPF1ItLb1
VCWuDUf7ZYB9QluuXLL5ZwH+zxOZQ+iaq06DH3yHxXZL6fjaVU4FKtVz4d3bp2iV
zfLM0MZzsLxWbC+pDuq69CIzZsuMFr/3mPoZ2IaDTN3m0sCeEA7gyua28DRXt17R
88MO8oj3y7p5vyggplDQrXlFDzalqp1WwokTZjXdiVo/oqQl1+rsqinUyzzw/dZe
pX3mTTrjc21d3PIERawi608MvYLRL2Sbx4QyhTAUX0D6ghB1xNfKQmL0Z9iGSpL/
ojylV9t4rs8KWp4c5kpwRNHHZxcHRZ2Z7aF7rpKjHpmjhgAlfftEn7S5wzX/lAOS
yCnu9rIpxRKxIQpAifNReQmnwMOmDsBcf0LfdtXihZGD8EbWXKykq7HX3tp5jCtr
e967rpf7FnaBZKFAfDIbwaEfPzywYgBZrXwRwqiAn7GWtiV7lsfizpAB7MR5J0ob
j9bEbmAyrrIr7j4+Yw+9nTuzXA47mgSwqUhdfZeVmh9/lyIjXqTomJSZ6Ts18F5B
FNUAMq+cyEOWln1GJujSh7YghdEUyQb+4YNleDkqsPkVoDCHHsQik6LZtfCJ81FQ
O6tcojCtZfP7oYocrzXswSmLj63LFQbYfDEykXVBC3puRbBsJa9hxpUHcENjOjh6
kk7gO6zJ73GzG3xSlofsy8bG68p0OlmZWDU9opiwdWUl5IPOu0RT8i21TJpv6hH4
PSQiT3SADrX/saEpqx/Ld/RYv0WbARy0VFnZtjbfNd1vYT+nu4tDYl825G68wn+Q
F9+Xm0xsFt2Gdcdj6yQQyo8un1p3N4PqU0DIVhqlBgdGMAhl+5kIrSn+nd/cef+h
YENVvBKX8P+4cHd8tZKvE4wDD8ZnVvU2oo1qMjCEEJcDtj4/vkH2nrSLWytS7FB0
dzwvLh3EKqdyyBFT+8rFLqsqw2I7tgsNNe3XrKUDEHbMW04qRtRtEaEWsIhRK+9n
iBeHnaqDxBW4hwadNjzzjUYliAxhZizZUylgdhtYFU5Nntkb5dYeBrIfSlnmbr17
UQyRjwb8DSQYHDJ2d5H/msoJE7vQ8u6RiP4TUCAeDFmnfAYPZF/NaY/fYfIUjapP
tXzGsLRpfwMLtO7RUs083eoL3hHHZEtI7CUTT3YxCdGWniAZSUZ0QtiGWzMou5rl
plSWs9IF3l+/M306MLggdiRrq0euBfZcGoGE3ELTdKetMGmSN+eTTR/xkoRH5QEu
eZzHl/ww1RlukxebLJy9Nvs4cimTCkhVcmPADjMU/M9tEq+YyAV6ZhqwX1JsEm7D
bTyaWdL8VWrhlVuQP0M0E0UZCqCTgV87jVZc11Hyl2Vtr1MoPY+c+N1aEyPhEarI
f+tE6GWDB0s+n1VNY1H90mY+REkpgM/UMxxmUHRWZJ5isARGVG9XjaLY1CLIwbik
DjVfUW4rw/NqCFooidYjWFjRn5SokSWUrl6bpaPRK9bOW+LG7Cz0wKYHoUlrT7k+
1KzrKSYpzXzoxp9G8X9EO7FxQx0t9qYCWi7M2I3swP/hZFAZvpz4jmc80ObKOE3o
R2QkeBQepmxGISX+DX7QDXyr2RQbHgwhlrbyg9dlfjdd8eJemA5/nUXew06rOKxe
m3eE/DYppG92HBiyM+YkEF3E2Phx4MfQcq7c1vQyUZD0rfutniNJiErCQcr2lRaZ
DDUU8AfcihJFqKCDCrE/9Y8uYqpeDoNEYWw++2OxoUZzT4YFe50Vv2hW2/d3L20l
56J1uG1Cm3cAcTqLIgKZwAxcytrb66DxA6SotapHqQyVGgHB8Q2+6TBhm9HrRG4T
CgFJaGNcadFiNe3+Dh5dAVsFVD27eY0kUP/FKp/euL4iT6mGPc8Op3jyReQ75fg2
Am3aCJDtswnGah52gY8B0lafDc/DYVa8fZ8EgIZqL46441jXrrBukzf870nVZpRI
QSCDl0UcANIj+Nmx4QEzqIX7GUH1qmE5/d8KjZeoWy4g76NQO1qgSJFFVqBt0HFZ
Zrjs62Hpj/A0DsIl17RpY7SeJ09ACMoqsM7pjnJtbfHOqHPcmifnXCFyBma6akWA
dcER5POTTPaO7i1VHcG3OO+yzPq3g1MMHVHgsHJAhIUPJCI+Nv9UmT2+yHDWstHA
8rAm1u3R640XS26pJGU9NneQViK/ND7Vx7JenAqy8BwL6LgmuCi++Ww5N4+gqRlq
wilTcS8DEf9wTxCrrpHeG5mIlRmGrH7y4ynvmT5n+/1Zv8zzKc0wPwkr8a00Vs7v
eadgVlZ74Oq5aO867E5mAVaLGmRwY9I2tt/IwTXu5AhSztWtebL1aK4afcY11lN5
Ty5bSn1bIgoACTl4kRj/Gr8ifEg7kAreUQHNJhuseG1KHs8hqZOOFhoc27ss6aEn
fj65fqa0fEyzaJpVYXPEHASbkyTEDJgUdP/L9fbG5yMVBGPem5WWd1WmOncnkpfi
hOMI6TCb57n83YRw9pfQs+rc2dO176RZSnEDsbMttyneM8kw8ZiV+pjLXmRw0Ei1
21rtzoM5q6HBS7LvkMrEOPZUPvojyvJO8aDNMfa8FltSD76MsVC6/ZMBzlriMrPR
0gosWOyuMhc4HjcDwcWZfBoCTwv8Qv9eBBEZskSYEqUHkg0uqt0UergW6tvrGKj+
vE4rvJu+zC+9qeWQYBfMFNJNuXkKv8eafSbFibppm8iSyjJwCrhFKRMbThczx9PI
iO7QHoFeeFtVJ8JKpuv7hF31JswYXtm9DDGjRx9An2fWX19yDyoQ8g2MLaZHdBA0
i4WbMEpeq1sY06gyEAwU4bsFBUVKe4EdSP47UqKEWMFOYNrdqr3PmRyJmZOUjdl4
v8YOJWczSe583AN629Wg52hKluse5E6Maw+eBGU6a0ARzZOm/svldS2ndhCgamd/
vQzSMm9tvRtQjHrY1YQ5tjv5fufPorMVwrLbiMNicXmJEUGX49vD5NqPxJA2+T6c
xOaRTXTUPx4wILUFr+YGiRbFfCpQAbhLQdkLvF484NNK9SAhH9xUL6oSOa2Prp/O
/WXX6GKppM8Tzpoq+Rw3eWqBjA1w57gIsQ1IjNQTjeFqvHM2g92y/QaLO/E2xlEP
ojhRdHiMcYBh5FHDR137U9kqSDdRkm4FButd/dyNzf2oo5/KPfvnw9PbCG8E3Ock
X/6vh9TkGeuGoNol1l3dhNKP7j8cOUxg5Br92+DiZ0YCrsE21+8p5gZjrg19hpEn
QwwEzAdghUHNOFwNa43yKAK8pZZbcClPtxhCoXQ+y8znhohxgJA1+1OljqKsXYtQ
ojT+7PDK19GXxCajEasQLxYkqB1XGPaeAWK/jwMdbUjssnEOEwirBAeowpK6qFdI
07tq3rKCQZaHQ17KoU8E7BsXN8FP9DZC5/COlULJqQeb9/R8nUSiWJyatbT7V0Rs
uP3xd5BulxE/1aIDnzkQlB8HJrd/ZjPkr4RdGHeE/ZM2FjyXte33NvoK0qbf1mJp
u/SLSLQfD8I4XXJsF+UM8nWdV/x4/SZewXVVMqulyAa9trZs0L6xETLk3nE1cak4
GA+2FNPep2/R+cp/FWzrFbT9RZ+oceluHhytUk+DHbfOcQv+5dREqI0QXBd33hFl
KAFPKRWHxsQ8ad3Mntz2u1SxVc8KujFYzOv/hHQ9v0B0KOcqPpczQ0KQDGSYPSIV
3xHbxdO9BfKCJGGt67BrzzzTorVtKn0zKE+HQ9LUaLEQuyCcn0UVaSYPtzLa4uOw
k3MS3/WwBKkNPYOpUzf2PUvImepHBC5AUnWrWT2uoK34F96iBwlwcqyZKki0rGQi
sZHDie2j0ZFxDNvfYFYEJAcaiUGtOMBeDjuRgAh7dQJxoUv31zYAkOFABATAUWA2
aO1/355XFDshdY5jHuxfzpkwcB6B5eq3WibEdYnvOtvbu/ZE7aXwoJKg6B3GLHhK
/wzWVsjosHhj6mIJivI+lkUhd0FLOXGzPeOuU4qxRiYlsY4kdsbNnCKvNUYiTOrd
EwoK73SQUV2oq9PMFuHbuXb4jM4g98YbqPrkfA1B/45VzrbQhl+UAqsH2J9FRo99
aPqCG8BmxoJmhkqypPh7sYzfTPB9fsvj/xSgzNn+fEgam4SX8YYQ0kHx9K5tv0ry
t1Ds/8k75BzAh6CapjeOYDXLoXxzszCDUPLc+q4t+RbQKb9qKGZMUsb2cYuJRXKY
VjdsFDvbI8emZdsqeNxpNrwFxLnm58pDzlSCx1fAtVw1AYISw/RBYbo1zOoRoLI2
k+lpHgBvNKWuSiwt6m7sc4H4qvnbiTyxP25ZSh6m5RPIf+F1FzNcNKb75FH5lk2x
/CeQ+nzNMt/3BSMKoddLJHG/eO6dgJqYsKuhA9bZjuW4NRNbkS1AWhx3MbL4aAYY
HpUKWI0x1cEQ0ucUiI/kJ2+ubXoYBJ4kCGCn31AJHBUOJAd8yDoHizEveLuUyx6j
F9txlYfUOWxIshQ883195s/DYjVGIdnKNyxvEiIdeZz5VYzjsSHYRS4kkeV/seiX
liVRqgLk1cW92mXt2wAZrY1aY23u2kWiLW0hCw9SgDEnBIDPgEk9G0OgmZXW0cZ3
M1T5u6DJ+C1Z3tDpf36TG9/xh6bWw6ePryjHI3NHlt7UcA3VumK0mwFrq2YEC3la
OUuEQZmcjcuA2BBBoq1a+zOmuzAHF50l9J3pbAkuJSuQIZCFx13dYK9m5IrKe94J
ub+tTGxnPxNLORRKsJx8xy+p0DEdSVnX6ytg00aEIfw/0SQfTIaKJPFTfTBJb5L8
zirAR1PSKS/B0aqG1PaIaw38lmpYCqNor4kHpnBgdmp+xGK6Vh9vSl2n2C0KA3Bq
UL5Pmu4fPwtWGw9HUdbNHM4sZ0Vk/3SppRlHGyCr6CRnUqe530aoUDYZ1VUrbepO
+6iyRolHrDM8E7INbYE3+8IwjoYhw2wiA0WbNTENHDJ7VUFGQDDmWOq94BUo9YoG
fXBy7cBIqQiag99iBKxLkF9zqJ2lUGlT4c7NeQ+xjnsjVkJ9+mIaJ24nCDqDTeTy
vhLZ6HboRFsQxcJT5kGh3krMzGFbMncoJCXsaKKYlbVFnQ5bKsuBXd/2ZLLMpvEJ
hE50DE15EyV1clXODrtQI3V2N3z/DwW9tE+P+pnaSwmoFt7mu0yfhHqAhxYoXR5v
crmrpi5ees+njJ/Pwh0ymdFvnoPu2ugi+CTuMWpHUFWplLF3+tVtp+nD3kt4gxDZ
VCH3w8ekxe42QyXYm03fXyhV3+Ufq/338bjjyZZ6YGyvpUQiU8rv+XAg1DoYGtJm
tXYiVz4ZIFBKpaHBjCG6wsRJDSAx3R7frAW/kpctcSwq4Au/SHAUUqQEyF1YkrSo
x51LqvJaMJ3sedf0Q2B65IBiXDxnRzKz2SlYpmqdOy9DMOsCEE1kiFItXmi4FVA6
SEALZhk76JJmSzydXXy3eAQEKQvz0yj6FLrMN2rxB88ef7jJ5KBJrwB1lSJVQxIc
xetEid1Wh3kcJ1BsoTELgDQHYMMC5FjyQH05c9OG7dSeQPlS4cRFTHz8V7N9Fd6h
hl3I3EYfZ2575+4rCXHl+1l0qMDfDTWgjdobHISxRzIhv9lcOiky8n7X1X8PhfU5
rz+Cr3isAhkYtxr4ddTA30PQquOaBEFvTECoCbpHD+Izgrw4M9KwdemjyMpgBWyp
PAQrEl4makFLc7zD3rpvCI6vb7QtdKcFpSqbwKs3bg35VfFcWeRXm5lgEaDfLXHR
syGyG7l6whSHHvVuh/7TOXVQbnl6Zk8xgHT8vLF5yAVvWHS4tqF1xKC73TgweIac
dvTh0Um/tYtavDZzfeqAOb6L0jAreA3FFIBCfXMjCVUygCTfKxgXozJjzQ2QTt2q
KV5ZYB+BJdqHtbHN5vJaEmASnr6Br8gyeEO+CJrVKBg6uHwU4Yet9Swjyk4oO63O
3SqDsP8/FPkTxPJEXh0ypBnELFlw9E5EiDmCoBFhn8uX+wJVKX1VsOKvsmDkY1Bj
N5Pqm56EFKZhR2WmXVIG1Llv/PlrghKgiJx6q2x5ckDunCMq2UTusMGJelooekw7
ZZilvfAZgJKXydA2Tv+FYz5Ta1W7qddg2OfZ78yob6f57bpKymrtBvG4jfUIghHP
EPSpTV0EAxoq9Z/Regm07rTH828E6EIaC1N+bCBo+L4QtdGA0H8Q00We1OrPmtUf
Lf0vEYXSxE9NnkMpo+nZZIBZbvTFSLGjMFy31Wdg3Iq0TkGO4rPy7UJ5Py3zh6yD
T9Fcim0Yn3hyl3IaRmA8aq/Nu2xJbaEKDZSJy0mbl/qaOkrv19uGfYX2DljYkU7g
U2ZPSCoj0Ts2tqA76QBKy9tWT8v5ZJd2ezGil9JW+IEmKQDHHbRkkLZfUA7/Ju/E
gMijKueJny5uEADV2/x6HzM6R2pSltcDsSuVX1OsrfbhJt33u1sEqFZU7T0WNeZv
tjnWtUcVRdZJQWbJTaj68SFNgZXlR3z5BCvTY3WlgRdHo0wRvsRX0ic2RcIuL8Ge
lzUFaU7eyJAav0Lz/AsUxrvHe2HIRFJyIAVd2J6g+gA840vySyblnrKQr06erZaN
RCJv9PoQP0Lcx56Lgr9Tp5Y4O4DyfuLVGlZW2FanWFvCj/xsEGpiPBJv2YRXOdW8
wNj2ApfheYW95FLjPShNx6t0hKTUlI5EMNJDEwcjvqwQXp/sCAXEKn9wLnVAX1V9
apcKa81BUA53DXwmsSiqS/2AlBhoxxTN4Dgfl+sLm2jvySCMKLOs3zBYgFaJlGz8
q+RMgp4L1qvGJKXQopPTznX4wdBmg8kvjqIhz69DL0lll153XFGMNeYgVKvuOjqk
QSubKB3q2ddCcL2kNMTE3F/or4F/vZYVGD/sJarGfBJK0UBm/wmLnckeWyhuVJ6P
xuTnSTTWCSoJnu/mM6EAvMQ5RDs9/wWUjEhP3yUr79TExfk+oJBN94pIbUJpVRKX
g1aqAVDb3MErFlxoltGW8aDoflzEtxEVBT2GOsDd4D/ENh8WAZ4dSFIeyYg1PyQM
WCuQMPJhtvILCYnuLP9tRezLdkB8YLSq/TMMr72TXsj3hVRCz8UULJKeJpXCPHuP
cYMrl+RCkQ4LuInmSq2FVe4boP2Vhb54pEblrAa00/o5/43r7T1KaSQyn057rm5l
QKK3x9ow7KqmmBw/srQI20DGNeTGsyk8i6jQmHCBHheF6a/hPuvWZgnQM0QGI9gF
08RNYCujaBm1IzmF/frAtaVlESv2YGw9rzhDGdF/99LteLIA9yq6kKIWgbK0cUca
p/6LFWddoA6xdmUWLEq/JAnYjSCLvOVrHeQIkJ3r4N2hsDCiBSY2mPnt6lX4Q05v
1jmCnH5WuWfITFx2qpvY/nbFjZoga/NZwZgXtXcQuZAWyrbpdVsoANYGFi66NTvL
IJTeIPdsIsAmaBFcb3ZjDwSoHkHKI+QJn9u/rOTzCaoj0I+x7cHFMSX9/RfkZ/NP
PKxSgKCEOAWilHFd+eGWiQs8Q4Ic9iImFRrnhgGDl2rKixX5J/h4LRd+T3rEB6B9
Z2W3Xjzc/eIL0XdMqtgv5UqBuBPjn2+F2CPOCdL23JS6Hby0RaNIjzfqeyuTahoO
UHTtZ+gVvY+PInyo2IlqE6Omq4hRj+Lrnj+OuMjl7+3KdqpQM7t9V11mOO6PK9Cm
thyZvzavbuLoG6hSRsd2p43oA7j73Ku66z7KPfXbBIX9fAdP2POx2miuT2rUufkt
DiSuKuxWAcfFH46atKvd3zThe/poGSxrqzbHwJi4AIBjqZlnWRz0RAHO/PP7VDCF
Ypo5aIONTWl2etfgPpgK0S2Yx5ukCrGw8/V5w2J3lvOnfumIwSofs4Q/nXcNoGhG
aGweSIpHy9LN7slNScYVA4QVfeMn3F06k+al5Q62zdq36NeH4axvuRYuUaG3pVn1
Lm0zC5pu1hhgIQzyp5Vv8Ir+ob5WYoO1WYuh9UKMTr6hMIRNva1xbh0I9Rno6dh6
5NpgAVIwshJ9jrnrEkaHDwi1Bg7FwvmgMN4f5fGjFeA2nED5BcINP3bCH1CqjM86
Xh57nrW2WDkJ7ghHbbFRXYBUe2IHxjASD5YCaaocvOAyfjXNxhjn/bn0t+2GZyl/
wHjvOh7XKxKASvGSK4XxthSGxyMtbbotH7QCeFXo8Tegk/FroM4/oSQ6DBKBxQcT
C1vL2oLHhE6ncqlJbz6S6kkEt+9lQP68qARXy8QLjHCv7NlQB60vTIYXxrqG0jst
xbSG31xhYAeem9MwHEBsoum6SwZMibMMnWaQ70zuzXnQU0k3wsEsCAvr4OCJleYZ
yL2P3Sstl6+bVYmI9mXAVDkjjvznQhffferG0gdZvHGpFkj15rzUKj83HfjP3SJA
zjyy59OM+Go2hAuvcH7fKDuNzz6AyH4363t3P4kABUR9ciN/qGrd41VjjcPoLBNG
vg0u/9LmY1eotvdPgjNWGFF5DDpcEhvvPmyr8F8ZG8GA+MtBjojucaKBwaVALTdq
zP8lCIDp1Dld3QPxcCc8TQ90qvzqoKbvB9A8fEcaBkvySR/mZ7tEnymG4z8aACAQ
oMAEKZpaz7wTZBoDt7Z3sz58/lHytSzu08vypvEXrPlTNBF5WLKonLGDPY1zX/TH
1RQfWcebW3eGdkfwBZGioIQ5XABpkwKQOcUpsdMRW0QEW+BXRZyXBzuNmo2yCdLK
d8l/+RbWyETwAfmC6NyXEVTL/gHkrFvnQGxRprhIbdSbD29DK91gSLKf4BdvXJtZ
hz4VGExumacBBSkUUpbq0mJo3IFnIQQ1iZObJhgQZvT1h+s7vDkIQPV5l5kBmeUT
gq04ipqSu1fpRyvzTN5Etl97m46EdOi3SRH2RdqgL8IVO1a9U/adPTUBonvCcrOs
D1+iefKWQI+uQipJrOJiccn8G/nEQC/JPUJ/8sb5kw82wYNzPr4Pi7NNwxHD/K2i
jl126HGUXz2qzLaDmFeAYdrueSlw9V4zfVndp3wmmLUtA5lf9vTQ/WZryX2k6A0F
OYDo0iEwwhkwhKDFS4Sf56oO8WeLZTUn6lAP7sA6Wkdi9ARRQbH66DA3N5rEILYS
klRrjIBRj1UWb9cIvgO6vvK+3N4ezkMwgAcaT5pciZFYMM7VKc4phXN03mK21yRD
1YEkzEoAqBsapsR4Gb9IlLQtxc+c5j82BJbdahVUTDmjkQmhU+1hy3UkuUuVe5v6
x/enyiIS++5oPSpGb01IDEnQ4qAAMNLRlVTqB02s0+v8fmHicNAu9AvXCWDdsEPI
kR/TgIZxXiULSmJZ1MuL3/ZiEqcjvZQdDXOvsLMyqdAwwo5XwVvhk7ZTPbv2nv3R
e1BGX9t1Kzfh12WtEK1RumV8yLtouvB2EXLmVXIIMX49dfRhs5d06NiW6fE6pTgA
vzjJ3miPMyLuBqwP3qgVohory1jRwuij8rwtVFVH5lg00C9HGCwnqn32dbFHAit2
qRtRwYrnVPp2kNzAfsNLwv1F7fcchrUG8rqzPo4iB+uuaV1pfpMtkB9Wumc6Sr6Z
1j6yRziU/6kOSLvdPlrd5pHgKrryksv5qtPq1kJtm9IzkLKnVCvP8qaunX0Wws2P
QBZb2tRp18p25l92Fm2BdwcoId2uTGwb43QOQfe/h4VksU1slPcWfLgSEkF8Ew4t
UGZuXeo3wSQgFEgi0nbHt9yWoYKPb7Ce0EcNzHlIMZIV/W6mbnB+O6YH982Za7fa
LbtcM0wRxlQY9iOFMOt7YYViOMolmsp6s9B4mZ0N2gDM7UOOQ8OF9a23xMFp9wAX
Derv7jG+49llGsGAeNxtqBfzgL0dj/3zEsg6H5u3W2/ACqCSNk8ngIq8MAjqKovj
IBD4jI031bVZvuFCw5pmbT0ujo3bvfrGXGH+0tKh/nNDzoVgM86wEB2psUkhoiDh
yizB07SlzVvsSnsFg3hYgBWYQO2/78RH41XMF3QG23PyeWt9OwULk/d5+3kYN++a
cJth4q2dG08pg77ob4jCNIDJpRvXCjDUnZp5rKh/9sZfgwIxxdZQ43/0YVD35zSz
uDNLjkUCzkQSbKfWnYO+mQRsEu1U52On1xUUxGhkDM6dlYRWfMZyrEwWVLnBmNbQ
iL+W4o+KGnx/CJafaK9Hp+GdSNvsFWvYUj8fdHehZpzOqLlwoZMY4sD2pDmqxwBq
k0aWBHxjADWis34ZSPUJ0hQu8YC2FoBKDpK51nxQ8JSy49KZ2EPgiAXxnkAxVX/N
Ee/NsyxkRKFaB3bpjZOyk3f4Leg10oE/0FxTN9TYNS+a1CyrzsczEXCFzYFsn3Vu
0mn7eJ3c99oYTPJViwjhcWRwXAXZUWUjDu8zgKWyCKblDkQNtINGPY9rPudCP1WZ
ls0xL95IgZFH4dyYorMxD3HUVt7WcIrzT0xUQEGwAGNHkQdFIHTVRCbTNp68u2Iy
ollIhHch25DvYU0oEyos1CW2AoFydzXznT6HFENRfhORXfepGjw3apGIqzUctKIp
zWcdio0H8bKTneCe+MT6xFK/EnvoyTUFfd39qOG1zMsb0gaOpKCgJLvq8Q0cIGJt
lp3ZdrrdKdv8nvIZBDaXn17opBgdWdxoXJOXnnsDxLIBIueolJtS7t6bQ1dzQ8El
qggh33DIJ0nXNYjp1bThKnjy0dk8QeVMab6tRYMQqw1FIatq7MpPwXKr6aHkwedU
rWiRwgWnAtabi9FQPtDtFmrhpxz8m4haZq+HHCtYqIBRPesMpzTs2Bjwe3WNa3Up
0blqb5zCWcj11XDxl6Ci0ZQqiH6WljnaqqUeE5mbSpmC5zRuvZ85HHTCYR3JT76s
7qFrsfQiHQmlITHWYHbXTsrvvCgZr9FzEBeQvnvHaMabkgpEBLDB2zIAvSugWxNk
im5ClQnyc43FqjMRD7+AfaZyC0Jpqf4zT41qacCkm+6fSS7b8Oc08yk/ioo18LKB
+1t3I41O03j7y1fszPCQ9r88PNx3iMA69LjN6nDs29hwxtMQwlZdTa8fHjHxM2Fk
lJB2Sd7XPBDUjhmDDV/GR+7u7NnH/eNR8ZZ9NqrkqAH6u0Oc5B80mZnwT/veXT1d
zr8eOCBNURFz4Xgatd/yJZj1eKH6urfoRmPorIpuSvyQt/NpUwjcrITAH8MFK9cz
WEQsA20rZMea2PSXAdpfn+x8tvaciaag8SpiD0lsbjwDeQebCTIUZ6mGK+wFxBOc
5pDX05XvEgrBLeaRbFm1qQXiic/YWHowrMuTWtQMpThEpssyCbyVI9rPzvob+Vi/
HXW5SJx70ckuppuVIJk/w0v7aqXGAEy7dX1hsg6abX13fTSdoIxxvOhIMY5fHL32
Ojn5+6WUZldPiGzxDA7rtMrhWqzUK53EbMo1czCGX68BgoSbucQOUR6nordN+N2J
Dhs9GuH3k2r0ACjZFktLh65n5b1Dg/0M0Z73PENJa85qTltfYgbFCn/3Ow0ajjJL
45X7VBzmS0lgSXm3WdnM7yXWa/Qx4obJ5cPmYfIHE8jyUtClQUiwwwQh4NAOeRpJ
zIWxM3xOaOCVnEBw+Sey4Exu5QkvosAyFKBT5DWSBPKTSzr+YIw4mPFcDnOs0HlT
AtiT6t7xo2kuoCRt5bwB6dQFF8WvVgC5tLi9TNLiLTcHRYLqCX8gRV+CAI393Lum
FWpvX3Ohq/zt9U2teqCH97p7vGWjV4m7ZqgNsnLEtAMyKgbIK/px8ZGK97aJOR78
kNL7KrPlfKbtSzHMt/Gv65FEJjX1V2dMBeJewpqsyIhkRs66IZJyjlg/FBQ3EPb0
AUpxsRNB5rcr/NrdtYwwcNS/harsQuAC1dIjQPL8LCx8ZPgZLbpdxSGUpqXSwRGe
5TuDl1LhRMoiCxxxaBrTytLdAF3jxze0HTEU7jIvxXqAcHV+YWCwkPQ7Frs0dVla
RAlYgfVv7Sv1kcD50PEst4dAFCOxIrGAC/RoiArN++haHCl1uKujsVyf0JzULeTT
71yDWCjnfvPcXOryu5Xefj03aTkVCaJp1SNUVLNpGrY7nq1BfZEqpCIDtI16Z0hH
sjrpifXKRcm9jhF4fXOuaamymd+LyDmZjdVse4Gj+FwMBKNs8sSBEtBYgx2zvDyF
EIN5N8WTIEVO9pcLgpqyX57cuMQvvZsG5iANVQZMlbZTJwmqHiNmQkCFrhOXuQM3
+xMzQdvazL3YvRT7XjWn90GvoBQh/coNj+NlVM+yatttG10xJjkN7zqakcEbw2Dl
RfDfDt8T/D92bHbeOktaZ5gmH5rV/Rhw6kJ9l4JzycgXj2F8aUk2uwXX7WpDEiO5
BWo7MtPz8UcNUndC1fmePFb4lQWMPGGPlZKWu0GXJ0eyubA4IDFvfZVDumamtiCy
3JecvSZeLB+iGUe1w46hXeB6Ql/HaNZmozb6NO6rYOE6dLm63mfY3o5exckegFJq
mhHC2Hhd5LGQKMk/VUymDzPyuZ202VXrLd0kFcMjQnDCABYKTQWq8xywh2K1Gm7i
6GtXA9NlHzwwquFx+U19RA2rHakYpEjzz4oNoEQnxRXjBXPCXzA2YD4yf3cCDd0V
us7gcVfQ0/koV596SqtHUYQyZHQqTQ+F3NnXKXMKM4C5RsbBS8JltxdtE/nobd0A
k61hAabwOCrrpqkeQUP2Xglt+Hevj+DL15LFD29isKe0RQDCuA3uCUOiuTCg6gaa
vjaqojk7Ly4Pkq+5rnrBLPuSaibZ26w+1QN5bgzfaHvA17D0PZfiVi2jLqh6fvo+
3sYmVVcCN5mq/VgQa7damJcFvhOjOndQx+7nPg8nYtKkr1qGTG51be/CC9fYaZEs
4ZZTWDERbQGBB7ANuAtNDI6ekpXgDnyKozZqasyRETCz4ynv0xzvTeDWv5S/V4Lk
V5AgZgnFn72xgexws7BWWrUSqvwTy6f+qqw29YSuHrobQWUHJb6AuXKZj4E/wNSS
JmompQ3XXm4gibUQ/SUswsJyBT8fBC1B+CMhtiNbpCS2LsPuCMgRAAg1nYZIvo+Y
fAoglw0BqRtWWwK72kMwzEZmNLCoM+s29R4mY+dOQ38P9xZA0XDArlQPw0MxkXKT
h6vctQB6uhyJE7BlFAN0RnPF9na9FDoUFqDAGhNI/mwyX/0hQ7ChQ0QYZF5ofKFh
lHl9d9/G4bIQVREdaSfXd1qgqRCN5M6/w9uRbw/pGKItoyoTTUqz0KQGkDMasLcx
z2F5NfoIkSEQCmCfEJ6xvfly8l/b1trqE+LZ+QG+fTt55KZWacLYZ+qT6Qq9BUVZ
b+FfxkZUM58SfknOEsOclC4zNQtuwL+6EOZ5t9jmLo0x8m/yl1B4UA+4aUfBSchY
JzdT3nGHGLzBPN7U4mGAgl6NsbIsnYllaWFT/kTkCVUrEvx1Ph3N/MvR+gvp53PH
NIBPrRAlk8KTfn8XLZLmL8TotFgjfYorF/Jgr9EoUDfKoa4CKDjtcDCojODxKDuZ
aMMFXEmpbO2bzzQ9AsSBFpCF+Ml9UEfnnbdjakFS4jheKqOZYce12WAKQw6sXvPI
A4gZpOBBIsr6DlClXAcpjc/EhRMrS35VyIiRusx8tzwbnVbdWXqDRkMcDEeMfNnm
cIQLcdNGVTKUawUpALZsXAs0rGHhOvo5wHjb4j6kvBguP/gu+PzXsxKjp5QF2sY9
ge6ujpvDHgdGUJ3FRDS0gaFwBKPpLpd+UFeyh06C76mLNByTnWIK7Du5YUh3Bqda
geu1OdjboRptkWQeYm6bg74AkrRAAfN7zPYJj45lxnVjYpj6ILzSssOuBetmeA26
xx6zHVymW74NcD6JeXx1ubi4+w90HcU/9vdBzpqJfoNe44wVH5/AYeQ6hwkGimDX
FesQC7xjab9/WnSHbePUXQF/c/Rxc8fAdp63FlTjEIVfVyeGKFY9E1ofX+Z3ucsj
NysSTDlPyA9cEyipyoQw3dorS4V7etoy1QbZ2YF4Gb4VlOO1MeppgR2huT36YfdX
eURXVMfGfjxs4ChT3Ehwa2s9Kk/lNKpSrz3SwrFQr7d3WKVu4Td6klMiIJdq1bz1
e/uKEAw43WrSVvchDq4a4JU/cvHZmbO3FWgFQrSsyAf+q6RR7lIFm7cKx+XBI7Lj
LxOTNyeDnaX1WtXFX4CUu4Fx3qFDByoVtbyNj05F6K2UiREv2qzls097PD0WhULl
dOBn+clx76zVNnTKzzKNkVSQELV153BipZSzB++PGHzoFd6LpwYOLuOQJjSTrKN3
1ImGeLT2eoYqfNvUtVyoyK0b0v83dnKV/rctoFyPZCcJm939+axstV2KYKRwlpQM
1n+aJKK2lQ7gG54tHO2sflhIu1VRYqSP1cYnx3D72ea2rXAWeGFOKvtX+xgQUcTd
Cm55M7IZ+kkWxLQuMHfYYpRDIbvDuW9b2guEOea3Y3noYoave2/wdAsj6um3gZZQ
lRX/w9xqJ69FCwE1uKbQg+64scGX3w5cnRRGfuM9lrZbHYnGRC/AUhhy7XprSiMj
xo9M5XmbDj0XhosxNOpmHaJDoO+Y4hvTgpIcxIjoKPzNvfuKu8lkAvmBOIVzZouh
Ui+naP6ZcXQhZj6VxDdWcXcNWW0F+EMN8OeiOZo3JfyzZZtqknPl4pcP+VBnozVx
ecSab4dhLLh4yWaejgHTZRunF6ETwgqo3poXEgGr4jIYfa5SywXlTZG6QQU5Xtvl
EnAIBKZ/OoLvs1rfCRiC0CkV+Vl0km8lawd7KL/BEdD7MGHvXi0M2RTdY1QqrDnP
NiVFewqoheN/IO2WQve97V8R4zdRxq6pYqNdqrvxMowBPLD1+imehmy/8PfT8uEH
hMDYeO1Zsbl8OEB3IZMNLonpjTmh5ZPAIErrNm2HIJ4JjAt8Y7R2r1Z3Hs1F+RGn
Z003Auc0DILm0uKi6aC0lDOW1yGTTnmGZ9JtpUmB5gL+nuUOBzgt6JskL/kzjsmO
hejOhQeXSa1hHA/1aNx/bjL0s7SOt6obE8iKCQUC2dwaO7QynUKfbmsHaokK0AmD
d+xiHEOgyBE27acivjmiN3mmGFDjtrPpKLS0KcqdU8UFmOZ88gDhF8FiOktJ2b+6
ri7dKlH5hkIJYHUqftDGi1jEfBT4/MYaEW2lbGlM5RJZoDSJArUAwOKxFG6xyOAt
Yx4Gcq6khUFfGRnBwYvofcQW229bsoCDE7TkfyfRpxPZEWI+i5dLjrePG9C/bNyS
J5+mCcVcDa1/ShcI8osuBPVo71xFbg1o4CYZrSccHKQ1luRtqRkk2WS4eKWzZZpQ
D1LUX+L+s7tVllHL9vUPZnX3noJtwdelmv5jRf5Wej4nbXyK5tnM5GxQWMLrpDt8
Upx9Klc4tLiSmbXn7vkyzHM1tm+/lUbLdWWhXdewiRA3FWGFxN2cELvSZJRoe73u
TtFtnxSuYbnMlKzSPT7cnTGHwkZl8yMmlyuQDrLJeVJw6oZfkCC7Ro4Ao9yGPHHS
H5oqfb6AXiH/lcHsJYmSjFnQhosnGuSW3NBRO5JgN5IQC/E+8Poy6cKwR9UzgUtG
fByI0Pq4NSrJc0r6o3AaoR7GQowFPJrIxQoRkDJb1lLZyapHl96BSFwxfjBpQC5O
zpOz3G1h/osAC5jDrfoxA5O32/0UTrZNu/BOY74wDEud1W7mMVLyLZz3oJxYH2FZ
76Wqnc3w07seg+dK5DA5t0wPVfLf7GwSgd1Z/YXwnn/clx/RbmdAJNTsDOPawmoB
SQJkoYl4UpzQsIpg8ssg/QVCiJgxfgnDf7KXfoigKGJ4e1MEtAFqsM3abYo/tlk1
FoZ8i1y+JHrNqVvHzDkSQgpVyFWb6Ov+LiMcaTichem4oYJbF4gPll2o3+4mf3Rf
mDijT4Fgnm2nACFnJ/Z1VSou1l8M5HyBg5IkTt2KRsHG/UdKG79NvuwwPRfpL2FJ
4UhE6+BvwZMfIH5kh0b3ly6EvAnGPmlaH6DrTlKPIacODb7UmueQz4k7OxaoOuOn
lBAO+2uungZmo9gLnHiSs6U8enQK4Mv8IWo4pXhbEIev1qs3DK/5DT8nozuTcirW
YpGp0t/onfcfdS31Suo5tf/Y8KH2bOsmYT+96WcbPCcvdZvLSIgRpjkuYDyhSANl
PoEnlJjPYH6ibcxbEQRmsLJcPLC9iAH0S41U8NnfjUuyLriPE4GVGc95CrjE3xTI
pO9/zy9LcEpCfXbhdsT45QjPWSc4zSd42HN2xJHGJU7C+ZGkXGImBXSYrBG5WxJK
LpuA7l1bvN4cdaSSmTFDeEgRu1rNnBai1N32jZy7potxf/XJ2uYZzfnqiRFbT9pv
FOevFKseadpw5sVWNOBDf/FHfFp75nn1k9OPNuSq+H8PRMM5/rHopD2tvEc0cDU6
V3ttlGEwyP7iUS76TbL2Ya9KlB1C8ESNk0RHF1CU4IyD90UWEI7V48k7BK5N8mDy
/gwXzrwxiEgVqUr5cdOpSlLCwZ0UE2XFQWqP0jYNDwg/V4KyclyhGW0SdFTZ9kUh
T6phuNtJPrPvyK88YsCst7q5Em+WeHt3etI6WsZ0i001t4FbfpMWClMoCJJ3DeZg
fKAiYHJuYDUUnpPpkIOqjPnq1KO8ZTw4MlZqQtmXvMS/g1dryhNzo7HxkLBZubV9
eUIPCgYfg9AUz7eq4qowIwOkpDqOff7zwe8QuRFVD5qPvH4p6jWdd1n2QeUGBW41
0BFy6jGJHsyMdqMiqEc8kd4esQxzPxUwY73SntKvJBMWTMo+mZrLKUG6lr6R9Tjb
HyecXFvXWmO9H7Ei2Z9zVnVFi1ZJ7yext5CcsB3vKSOaXAJkRfuDtURHY42fOtob
JSYTtiw0HuZ6MTHz+yVEdwCPe9ySHJ5Ca45zJeS8PTHgzH8FcDuVbPq1BFjVrPwW
TYtIbBT/WYInwjmGl4r3kekm2+/CR6DQfd7TO6p7TVW2lgeFA5RFx0RLrXEJtNS/
oiEw7dWm/OVt6VhzaFcIhPFjETVpTjlY1cCfSEgESvxoBrgvvSxX0MRB7GmTwJL+
WkvlFwvUUsVBPs5mLNH1iNUP7BYcV2i9M0brdEonBHelp9rrY50xBAwH3uQnVjZL
+fc+V5pBa/ese7Udh/TjJWhnWDkTD8K4Ki4xS1dUeN8ZoES/y28K9UgZZEMlhHSA
/oURnfYI/scAwEduDlXLFbqSq7BHH6D/iJ8aLCnQ/Ml7a6UqPeZUQD+8lCp/WgvE
7tnFkiZfP56YoTGfeaPw6VB/Xf+Q60jT3BOb9XfT7nRtg23ePJ/sb5g4W3GhzHKJ
Gqj6S5RSalIo3cDWpXGQlkwOae5M1IgIm3T8/Gj+qv3VQ3fnKo8E7ElO16qeGg9D
PhZx4wSOjTaTdLLvtSGJdoSm/kp40IkG3HyrDdLPbcut+E/ejaxJIq2WvFMKjkJ7
QbRY4WbEuLezcCjEempADeVjWj7+qyhdIkQbQR/IlTj6KxY4AlxulkFsx7jmZyX5
GEQvpUkCCscNPfVScbQZy3Zm5EV+gUtChjG4Sx3DTdWXOypE3r9+jMz/lPXX28kc
BN2EDSo7PRVmZfQkocOWcnUxi+hJfNu8/LECNxfPoazjJ7fBY4y1Y6du910mla60
noFKzflwwDJIQRyeY7Al8H1r80fdpb8fMD++M+h4eYmZK6lzgywkvRODkFlMeNpE
hdR4LbiotLsZ2BSxdB7Eef8QkjajXlogdHFfk2DUlPIIi8z3lak7hqf7StdTtZUJ
YA0CpIEu4ddDDdcBLkjM4AQ+MkFZw5V9r/C+oS7ZFre98UN1FwjzSgt9dhMoOUDV
36HjA/Z9sePAZMssyNef/LtvwToATtQ6fsCXnMBBBIqJj+ddkiJZbfDnnPSLAnE3
uO3E1UeOe/mU1h1hJPbjUMacEesjaGmCM7w8eeUZNeJYUyXr9ayP0X4Jpdvm7dyP
34c0SCZyEuhUuUwTv/jTR6zmyERks5Fo5innr85QNHdnqV0aOo8gJ4fDDeC6W716
u91rw19fcevsnYynpyhu1YKAQdBSdruCrfBCKhGburD27Y/LDlKYBuOEEgYiwUvN
wFHbfGsBXUsXLtdjjZ7NtA3SX2BX8v8jprmC8DJMnqkcxxCcmtlzgH7TFv6Uh14N
kSNb/9B7l7EPg2Y+KRkvzoRvDzEa1Q5ydrFFgqjkWqae/VhFcxaQjY0h/0YDujk4
6Le5EL3EOKvfzokjZF7VgaI+dahVrOvcgGF5UmQn6VsRG9CXvbL/WwOUZvEFP/Mt
MFTpiuC1sWD8PKCfvoIMp1OdYhmg0QdR6fc9cIqtUKS/LGVBBD1ldpmZxYDKn7iy
X7aG5lt24OYxxtLfabinsi56eRoeBP73GX92xPQ8xSm3Men3hVvoiPXQmXjuwuDD
jzYSXpN+y+HEz7ReuklLlt6DCXXj27T+AkIv6tD18RQVWiNu1PqC1BPBwA6bD+zF
mMFswTzhOHVHH7pHMU9Rh3virhvc1hWmmPQ8rkmQ9Le2KGBl+dSulm7B1d+MznNh
j6st7pH5Mhaz0C3FCgRaJw+PEzUxvVGL7tCwhf4B4fEH5umISqFVzEoMbYGcnD+S
ceWOJqGt7swRmSv8cFOeVUj2HScVyhCueMRVe836cDQO1xgFwwPJvLyaOd5uArQ9
Vy6/R8lEeibvL13xnTbnq3HpdGtKPUJnRbh/rruyNQ9AOHHHZiMO3FcqypuWGjtQ
ZNifZStewfB8Rx8XnKignBB7ocUPkybZWakSc4ZyscqKt70fkCjtlWABOQQHdUTw
3Xi2peZLRCgEGFCkyf2bwfr1wLs2Yfu6XT3w3mozwNIX0ldNeSKfej0o+PxshL28
mayUbKHHlUx477lnZ/9gJGSFQHYfPMbsHLmlj6vNnp0FoSqXbQg6XK3w0Aj78kgD
UcLAKWq05UwVCDyuTtsoxStuJB/ZSBiDpftTezSE2eUAHM0/0CGL523wRy8JS6lR
WPOg/tXm63iWiwc7KwVx68fNrA8Kotu5blB6MEUaIbJ/QNKYBzv1rqrGaMkRxfYG
Z7iJJBiyuIYY/F1yFLqmA2RaTmM0z5rux+UxvOutnIa52q7f+rSHKTp8JyXolsAG
CvoJiZ9+rjgEd6fbtjj8ifRcvGTenKUtKBCifDb/o1cvWqaVbaUBeFn8peLvp7lq
kKufAaZE3nu1o6v/BkmLhQAewfJPirs6tli6t25rHcpyBQcP+mrvqeqShQ0DwfcU
ym4pnYxS+vemCYKWAc7H5I0Qz5FbcJlc1cayj0QHAn2dVzIZ/RGoLDj67oK1oQqX
HOYFpxSaxu99nLNSgQ6XHLJzjF/X0ecYa+5s2R+RPBtwK23EI1CO65iCSxoRr4jO
8mI9KC8x2vz4dgHzfJpXb3QSRyuGhv2iA5vFeAEWjvmjW21WfeqDrSD6EA4Pa1EK
zxevM1bQCUQoybuuwk8HqwVCwLFD6wMX5CymXFRcK8Zufb2Zj5Dy3/njp4dCr8sL
LYiG72qE7dvLcNPR1FzfPbaugB2XT2zhgiMqqU8CoB9TxInWQPFtu5lzk79Fm1+l
8z4mGC6xrRY9iPHOv60VzDn6WlDZfWVOocv+HsSHYFjcNtBHdvvs+CsHjrfc0eft
fxBSuGKl/nyTXsaVp2q8kdQBP8yKofTw2T44ujfGsbDtbLmq4o0M3WVnODj6yyhn
V2GNWk4GZGhv4XoKEYxHMNVDmdzF2BDbcCAac+k4T7ztDE8Tyt6qvsuALNZn16ey
DnDssIwZUTLlAdTrWEloorFRY7DRAjjTVTNgxX8V1AT15ULY7mjF2DLCQUQFCsor
XfYN+jmkJ3SArtSPdRu3HwR5Js2JU0Eku98tl4qnHGhOWngqQ4uQhaTcchXr7iyp
xKpXt/QgRFLqmKZ5uWomRie4QIDe9O+Fg4XDWYOwJ/7FssYXGSXcSuX+ESo5ao4H
75CWQxugvpITu5TC/pzfAb3KvfIP+fce2T9MPecY9BMA35tOI8+yUSj7hnPWiSkx
XjRmi4SMbf5CXXGWN4uVKSWsc8h9lVCFI/O9SXbTZc+xUBqjBcE6HiGf9NHQW1ok
0zyjHfk+g+K+1bwHlnMa9QTUsr0a1q6PSgHweINAM27ZQ9Wcw3MzUK8PCNayLlqk
jg1vxsSbcaciazpCWyw9f+YEXNGj+I8u4Ao15HxrkB3NEt5lLtMSVfWUp0Arep2z
zFfOmFVRYVATOzYwNzXQDW4E3Qc+Sy3xE6+hy1EiAA/Vq9zcdaP+ZBrQ45Db/MZE
dbUudW7/3NAMAHSrLcPtzC7YfpzEDrNB4R6GZ6z4JAd/tevfuBQ4Z6QKT3h/IfZ6
++0B8tG3ZA6W/8FfRT676FEB35WvJD/7QlVlp76qdl5HFFgZCjz9N3O8CGj1HRFF
OX/iE6qsZbyLPaHhcSrASmqHL5++F67WtMRtExL4XVBkclOz+QHakW/BPIAjjmaB
je3tcozHGvdXnyluBQmCkKlZgDZBHAgcVtka7A7U0YWYIlXPVFPRDmoAf4xe13vm
z0jl4o20JsiUw2wDg/k91OE0CZVEt/50h/yCF9jHUyWG9s2/YRpfBGmYxp5KMHiZ
Kc9zQQUPA/FEsuvRXrKiZVPuJlB4SXu06SvZVeYjdd3Dt+uCdTzZUND0QZfadaMc
gcRQqkAPlFE5qrQTOtQLjpYmJMQSXc/tfj7wMl62yMmQCouUwOFg5UT6EHVobyMl
B3mRn2uztkbSWLC1r1KCnlYC6qI7IjchYpOkW7jlAF+YWB6xIapw3VWbsRGu94NE
zIES59OhYLrzDDqIJat9IXo+HZGq2rUvbWSu6Ro30eIF7wLk7ik9JMl74OFd5ccT
vGqzSYRlZvi2+3qKCuZ/qs2AWHLF2mg+VhmsMHhm+TxEeXMdod782RaxDmf8tLJL
HPvphip+LjkrsOLYuJz2S2ULqXvC3Xp5xPsZu4NYg2GpfBpj8p3ynpcwzS0MqUi9
vjMbaDioeK64W4EcYa4GprKv2u8LPM3doy0IBDh7BLPXIbg1IxXj19U8/RJwaoKs
ufNLvm8ltvv0ASsughjIr+HkS4wLCb7pzJ3H5/dwfEiD86gtVDnHrCD3vyx0jzNc
9cjhT1WYjhaKNqrIc3T5QkV1gMtREfNn15ZCAKKCd0DmG4l1t1PqhZmRBSGSEHfj
pfWEcM0Vn01gLLEHlaUGX+hyKIdi3tr3AfxVddb5k9yTrq1pdErDmoo3xauuEYpp
8tfr1yZbrniB/FBxpXbwblhm9U7TXHaav/jl+wUR0O+RuLwlQOFMxtNfR4JKQ7rx
Dmq+M2b+Gu9o88U+VKPu2mIUdu9NvOwvcT72UQo6LdTQDVnUhbe+XREk0msCGQU5
I28q219AtETTcDIEYLnfPm3+TscdaUshptzEAT9ujgCmjCx98u+WU8K1jhOiYNee
0WbKNjE/8u+kDFx+hQ58Ivkw6IdO24mbB5hDIHH0SK/CqvRGOY+73n18txeu5Hab
ed2M9ZI4D5Nk0OeMCnBhI5rA3LBGRgZPTcGnPa9XQqAeuUpTqYePGdFuLP5gq6/T
HO1SoakCkG4/PahM+XAbAUfGlN28CacBp3yCq0zXeakwVsKZOqLON6RA1MpH3kwZ
QVLUUHPSjPs3GAe/kUIhraz6zYfp0CslrteLAEAPSuwQYwIQYbEplpAqo4fNQK3r
R/LgLw4K1pQznOeJ9DQ9fanUcldJ0Xby8jfSrWqpsQgw7GTCRA5dcOmR2Z6L9KMp
GYeJKJdx5+JGlsaRG5t9eXIiontUmtk1NxjNXWFgzGXqGbuAHXlGRyAAIPKK+Ah3
wIVbTTmDZAaVNKmIWUuW5r5Na+6zMY6bbCG382FhUcZx5Km7J3WZgbN5VZZdbWM1
m5ifC2l80opPttBQyRbTFd+b7VjsaytsvSVDg/hkCFy41eVeKCxA8xigeDO3ixd9
Jvx7CXkEWKDC+VDVa0CUBfrVNldwONMIOfAfqritOI9Dw/v7Qq4/YygGP7lt8JFQ
2g9QsIBMayfGHX6QNNndzmdaRZbGXOJbVczg61Y7ABvwXqE6wsNsKsAyZjiOxr16
9KRLE03fRF7KLo4jxL3UPdsleLHBeo7XPGZ3VPV1s/e6MjSyFv4rGwu27RRqXUzs
8T2og2y7trXE4FQ+w3DtCKcgV0ISFCbEzpcJqX23Ub7E/bUn/PlxB9veuilTmnGX
4pKQLc72wDBDeSmuhZNdx96VQ0i0pmTC/LIaaaUjBR50UZyvYQLtY24cH/ezK/zD
mAwySC+R8hxpSEZkuKvTOzwEHBM2tD/vgn07IppVOTi2VekoOpgKV5/iJNsJEZjV
Zy4yrXtyrkiUxEc/lRj1dJfUqJ3Bu1V6j4Mfm04rk0O5Szk3UIlKJM98f6xwsWiP
vPspryKUuUzD2HaE7oHcBA+OubswJSI5wPF03MtP+4m40Q1r8wgUEvUiOiqnIXdP
o+uni9QZenn4OQnyTvEPgbDfWEyYExQNFiJ5AlUEIG8lOClj+er9OrxH77axjknq
JpEcKZZITTy9ZbuzIsnQ6asC+sRrWNsxfWu72sVyhFEMRj+ZOq6fz/2zD/HpbhzQ
pzm+xC39yZJpqFIaTaBlZvzio4pRMdC7xqvcg9Y+Xt8pOzCTUeEXPZeFw4KhCbRl
ctj/lih4MhFBKesbzWqyWuRS77Gn0hMqYl3mjwUnrjkmxKmrJ6PnZinOD21x6cvZ
zZ3J3OeEr2I5Js/6DlPZwf4t4rIpCqcEQJULBBhD7wK4VRsV7k8iKgS8A9JaT6N8
V3eB5y6JRTOCnEkWMbVS6WNEet54rTgGs/MUurOXUlaG4BTj0/UM7jeKGlds8wIO
DOuc/6NJwM2dhtChTxi1ZOlCs8byEyTRyN6lcd4Ws/b9CrHTi4AMJauIuLKA4ZcH
KFPxMBDe5W4o+R1xJB1XnXwdBxnzSvpY0NGfsZimkGoFtvJjzJMypmdmrGl0/Jr7
/rlCnRuPcsOIwxHUIFrGFXj4acf/rPg38iXUrdPxKjAra7RQZIzFUO1/iTpKPrZO
+eKKxZb5YTzR24NETbiL1PM+b59GbMlD0LMQk4ro6pa6fsoV9BU0Ogq4eVJj7ZZK
CKR21M6cb1GlIBKJCClKzmTsaI0NQ4nP/Pn6pl0RUa6zLVUZstvgnjwWqDItT5pZ
/q5Z3f17ZuesnLVq5Xr2Ay2Q0DOZLCMlsYhDIf6ejKnCTErxr2n2EfwgikDFvTM8
at8uYxIdYy30QHWtIUxtQwCX1vIxNpifxmJJaWfBNv5skN60X90aJ6L1JTHCChiH
9lokjkt8Jp1wqwsT2WHPN8nlm5MR5DnFc3XbUMqxFHSY/6kuX7aIOgLAvDjYd48C
W3Dl8G66I1h+ph9CaMKYx+fuk+k2Lsbv1ly5RvpBWG8OsCnkxj6rhe4LOHaknIsS
dIPpQgJc33i5+NiXnTVxK6jgp6JEv6KV9Vdh1Z3AQRVP9OohVz8UP9bdyePkbbLW
zfx71pzN2PtDiyNiwuW74GfF0/HFQKmHBwnWoKLKqfqt/JOZCR/pC+dyObWxX1bs
HuboI22yggtoXGg4ThtHGG/T0MZ4eCYo6ObUkrzn0fyabHVqonG+ElYA2n2ktifZ
sZGLW3h9IwaRpRmAI/BCDlZFx/P0Ur7lwtWlqDUWwly32ogXAJ4fc+GmxypeX3UG
BZFTdfjP20kYZkLTJ1ku1PJSfuE7a1V/80AG+ODkIxUi7k3XwelLl+BbqaYQAszg
wv8bxffebTlQilZmuDHx9LsM1832FOHTzi4nGokjwsQh7OPDNkl4CYGBE9rDey42
d+qaHhn2BfGMs++nYxQHwoJKEdkZg/9YxOncmjhY1aDSPhtNc9IZGnnYKPmUCcUq
gGIfkaoG0aZh6gRvNEX8ByCNqNDj/JPjM7AihWdZVwVbr/WqfPhTf3rDFAfOjpru
hJ/PfjS74Ud5VN43hxe8Es/vJYTvHcvotQhOfQ50tW1Gla6jTbAgsvoZYdqsoD8D
OnfOBDBoPuCiyLmkpV5uNusLHS+YywN0sERk0jxjarfzf/ncP0c/xzk5SetG7Gsv
cZbqbaDKSm9nq2urVqMHkpAgUVDXkKTgtmP1Oz0A538Rwvha+kCdHQYAur4YU6Rb
h54eYn7gEBgIfrTo4e0EsKqVv4tiOBOVuFp3j75QHjGRyqAWak1XgdqJayEoHMix
AQxx2tZjcBzXFq/1ut0VzZCOI1IZTkLHq/P2F9wUHPwTtrIRrFFRoo4+p26XwVt0
I+/ai0GvRa5pTVQMAJYXk8euWKBMFEMCR0ZEnoGmw0JorE1o2HRDCQ0tg+VXicUn
KJZA120M5fho1rg5ovT3pUH6t9yQZHioZ8HC4ktMx9L2WpQs93effPcM1DkuKCPg
98MzCJCgW/TMRQWGSPeBgOX8Wk5Wuc/PzsXr2l3zLm7mHeVW7nEVKXc1Jv4VGT80
9AD1L11bWkInN0FqKyuR2Ip3585xB+Ss7NxYLjZ0LIWiGPSQFoH+oh0SIJQPFnIb
7R4gpZE312jj96EN6jJq4L1DpDKDclicAe4CsqXgEOAJpxauBq2J9wWW+qe+FXef
ilfdr54vZybaC68GFbILFEUkpwHSwz8/c+a2si+pyz/Zu+ulkvtvEVPxrwuvlQNA
zej+n+EWo5WwN2FNTaa0M7YZLzI7r8/Q6GVRH7/uoq3uVXhisT+//l3i37sU/CNx
J0wvTjFtRbb9APSvXPDwSC/FPIGvcZbWY3PONK+a6RCz+691okpxm7Q8gaqFLCeM
ON6jXhtkV0xf9A8xJsgEk23gMeDyKS3T5Ye4nE8J1Z4api2FbxTOSbOfqDsafWOR
17rcwb8fD52RX0b1fCcF/Ln9+hZLomhcW6rVp/mDduhazS0LoLMmgb8f52EDBYd5
sFJKCDdFBr8LCVM2rAFYZqsr4nxOTpPBfc5FEl0P3jYEvUEMvoq4dbIcbzS+LMOW
YWfxy+TOrOxsa0Bun0VGcd2WoZwpntUh0rP8R4tbyXQ7i0GmeUSqFP3PvGMAsfbG
qgZpTnu6T2FPHcwzej0ISOVl3vIlsFdlS73Y2pw90bvnCOPziQa2RsfPfFR+blxt
ySvPFQW2pt9zHqlM49lOfUAkwJ5teaSH91ZKPrw3LmbrBNI+qW8ykF+DLvWO03e3
BcQZkeJGlRabxIH63p74Al9Cjs4OtPS3/74O0L4timsC2oBv4L+zCtBtOfiOa34C
K5VvXiRHesf2s5NKYBzhQQ3xMExHVXKpF0rF5FFrKsKsU9wasYxWdc807e1FAPHr
vm5rjIBcDwdhWvHG0JnyIuGbV3Efavjl++xz4fFwDIYxU+zKuQJF6th9dpReCDoo
6tI4MCBtL5wJtMgvfLsk/Iu1ILUn3TLY7avoC2Mq16aKQYi/G3tbWGW0AFEYKnU0
bJmYsHs0DCTphSOH+To24LnfmTIbDh9mU3qe4xkuHu+CEjM5v5GrZoT1cBfOIJME
0DEijKoJOvidX4NeGxO2X2S4rR4qJLQi4IUca8P72Z7uklVhCqwgOFYc2Z04S5dk
qbGqj6fuS6m0zkqzYF+rkmUiBGqiGuF0SykHM7INLhXRL7eRMGb6nMVnZw0PK7m1
7yvh6Z8lsk4KeSs+MvrYjYffAL91v6DRBW7bWWA/o/IjGGAb/2wIOCp9KrKJbbwU
K3fzPpTrgjDpBo/rxXmoux0GpLOxtbx/aVSNV3gq436gU3ToifTLdeO/YrJBD8qm
QRv8ybOsszQ5K2uL9zB/k8cWxnje1IOGfFbGlClx0ql0f4NVuxWpapxc+2gO0grV
Ia2LXuVq1iB9RjcHNgUmUZAbo7sek/GfXa1sMNSPIEFRWSaLYah/+wvR10/R5G0m
p9C4RXr5wgnlaP89/EUWowaY8Pnvgk2FUU3TMFJZCrNd7ezTMSJn3WKVbLYOJcmU
RixE70qH3zYzTVXvOdTzgLiVIDp1xOJqEfPV3NLCRYvNtHDPz2nmOZ0veACw1Ang
BsfJEzafL0FvMqqKtTpFPS7g4hpXfnKILdfCr6IbnBIvj+Z7wIFLy9FwNocOKvgS
Fe+sxA6T36UyiEGQu309WpAqQnCesWEG7z+zp7Io3VK0KWt/W2oe5AWZREFjOSIP
xIV5Ja4e2Anz7LUPTnovyBgfwiUzOKS7qX+qw6rlsiYkHUbj5xUCdP5DQxgc5R0c
hzYs8Eo8JaXVHTX3GYc2fOcY17DUENv8QbtlfLhvrwZta/i480MXLUqHllBfHRhh
WVKJEXntaepxxAEkQjQnZE65sceBdeHY7t+mhZO/B8FzuQfmh7rZAxS0pBLZNvvp
o6eu/02YiEA5KcKoOGJ8qGCy0DuhFcq+I3kZdh6Pw7BvVuPmd3esZ7H3bczhtn1U
kHQyI+TjcFdx84n2fmzBcNtRrY4lGCQBtURWC4Cyjz/s03sCvIR89eC+Mw+imutw
RPDkTbOVC5JFqOE3wh6kSS04AwDNWH/byqQ79YNEAU3SxOJtnSTEhqDxFpFxWd2Y
qeBDz1/PCmsIuFvCCiOft/OnYDxRwR5jBITTXoobQ3eZyi6nKvmviBkVwPQdrbdO
4UnpePJ89Jnv84r92qQx3DiccN2tVYWOx1Lrp9HH+/YWVU21d1bqcSPfAuNuAZG1
dbO6wGFFHXVgCumh54Tg9bj/tIrwlyiU5gF/pB6Kbk0QeheJ20LtuM4Sfy5Xf5Ix
odSQIsVhGTCgAs+hb3fWthCVjemWFXINUl81PpJC2oFhUbxKp4ZpzW6kujqacbS7
f3vdUH3wdN5y+Lx89GbXEk/yZuVfvqXUQOllamzevr8epJbJ+KvDK+81fqz7e2Ng
OJ9DTwRsAIIu5ElhNStxZ7edfsLSQDYnyJBnfebLFRXxcA7l66MMzEcVmYTi6til
0UmCvTQoM1TKwLAe0R2UbtTjFOyTVMBR61NV1EGJV0EXaATia8ECpX9hXsk4BNow
cFaW0YQlvOwdbb/IrXcBGpFp4wNQLZw27POMufJ00nBcRE2vPKKxSKz3ziKPaNdm
M79DkPitpN89Xi4eoIpS18/kAA1ys/b/7AZjhRo95RZqMCnRjhT9vjWf+++v3QSl
x4K+nxWPCmsfDDu8Bi67ZHru4P6wsJ2XAh7gPMOWrbWB2RZO1jzNFpgHG1RDazD+
c886d2eVSqEqnddSfxlVC3+wgEp5mK3QkJ/YJktmwTaauG+vnTvxkMy5viflKKUI
6mmbeF/x9ZQQcm/MBxbz5q01H/YozViB6CcI8nceq07mpbAebqk6noWPk9GMdgWU
TI7IE4KVvM44oE8jLiSmHB6yHhPsYZ290MhRRvdagdDUkaVDWgHt0MKLqSNjdkw1
GXk8iJkrctnkJ6fxX3fGprSf8b0uGD3G19zEqTj/ftfJjTiaIGpvXg8SJkvkXtNS
TqVEDo4LYeyRhN7WsCbtzJekIb+QPQLF6C0Ev38jhOzkq6c/puw7qh39+GPWosVF
r7A4rDfn6Pmr4o3UmbeahF3Li362mH0vCaOIqGxJnNQ9Ss5NN6ZLTC4RUGIkbIRD
GPY0TD4BGGvcJbeghOjziKIHc5WGmKj+soAR8PVKkDxRVqsba80VWNsxVA4gINkN
P5Pk6k4JWEkISd7W+W/9YYVtHKb8agMXS9H9Qv71l8VnFgQU8CI/fH8ID/vlmeuu
kTmbr0zEUAN1H3ryN82nkrc1kXJEItHBW/IMwUrHAF/7BRgX08XsLKgi2WYSzjN9
tBsxGmZSbkj6Si9lkwI3e3Z1TJvUBJ1bf84TYuROZcGk4J1tVhxpb7JYb0vjfW5p
tXVXr9lhQhJOXe12c1mYDDB5pvdWReV+9FvMp+eKHvxws3BaypW6I8Xa68EUVpc8
l24oBCqCQdWZm9bN/PW/7eKN0XbaYWeGeD2iwTOXSQVD0U7Hmy1iaOPRfIysEm4J
uranXxP7rQpyP1DouYEGMPbOHiRRObcnaNYBBV2t2H/UQKy4LmNG/rDLRn9bOYsX
AJ7UchXEREapEelU/efDAwFSBCkc5PUnq6/jV11lLLwG1w/G2CEgo9P1e7j8XXpn
H/DADo/ONFBdPj6aRn7FM9aKR0curE6os786W2OFziobh/hPIUg+dmh2ISvOKf9/
STNEsFZVDUrgqq1M52Qwx+jN7PMm+J9R38X3IXa2HPjtkbpRMRiEb8PKnvvmSkiB
2qOCgzreXYmBBD0c8yNdUW5IiydalY10Xdhh+2/cjC3TE4esAh75gSZuYCD99i7g
XVQnw+bpoEk08X6aZPkQxstFxcxECapEcY+i3s9+CGrsQzfqPZUavScuOaUQFSxU
usEUMu5XqtAfBYUltUx0wZ77gMR2Jj13tqZoR21btJNz/YpYq11sq+Z3UDqLHUHH
qZUvM6xiPz3dJ6Ip7P+Gb+eVjudv0OJTSAGmRjSgN8wWmVsaI90gkYVQ1Bp2Cv8e
00matQZaTr2L/r4lIkljoOVyiN82PsNNBm9PC0/N4PtGnodw4f3CB5TnK2G5UwGp
VbPKJDh0pwMQapCcD6joYdBVifih7tnn53LB6VB7rId4CQ1/mVY377PVFTYqiueQ
FcnHiUZY8Njcz9toT1UerhpdkQQeHS5nP/AYMAkAu3q/D+smky6WBJFKWVF7PSvM
R+vH8gFSEYRnomEt/c1sPHf0Jibu0DyPYA8HkyFw/S0+psToElxZ3SjrDir+Hoop
dW75FY9ECLBVPutZuQ/e9Hsuok7m4HDpPqc3WeHideRrHIDeFXAoAOZU+BJ+yuE6
utiPMZLNKfx6zG4KoqPnfChBV+HvBVhgwh4cMhWj2PBXVOo+a5PY/2urhMjFejZJ
m2S/sx42GA+7fPa4v4BBNzfQW7OhEqbDac8HlHgonSpdVGu30TO0Zm/CiaVqE9jc
0a2dIwBC0GhVthE7obs8Dms4jgwNHlbXekIMkhtb8yp79I1OmA47SxRqJEDeoFpS
LJCaXlj0sVoO4wz+bE7IFJGqaBCtwn7SJfWrPAjpy6ZCT7o9v3lkM9A11l2A+bF9
ggK+umgHUKkd4OryLtzgh+cFzinGSBzAHMAMXHGL0JGhV4cuJu/kHUnv1pgIxi1V
CIZBPstsKjXkxwTBwDZJx8QrhHKOARgmPB63HNL3T0qWuizKpWuKXRQyNdTWq7Dw
XnPNgue4gfwg4L34jHn0MQX2lkSWEnJ4i5ltqcOb8ZyP4QpAwI1mT4v8o04M4hyL
kLa7lCcXjB371ZA7de9FAgbH6C28NoPNeE1PTFzi4RejyUjMFU/jOcD1TKSU08B1
1uPo1/Tf8nq0sUwlOYJYHadOFB5lhNvVpwIUEr04p/ILbPY1GYrXld63kHstNbCU
ZS+me5DfstzioiXCKsh6p6g8G+PTMO3e6oGnG4dCSHREXtk6l1A5OoQ7iwteFqDn
VBG5lANM/fFfUIG1Uhw2fzEDGfiMZaoNFAIzge2zgnJUZNUK6x1emzct6VSzLZlJ
gHzp/QXGoL708q5PgBJxQMvXUwTnBPDp1l7z0hNA1wC7WOC2pizM4hh0R+vMN/SH
3dS3NB6XAYZZ9IhoV2Jn6Ov2MmfMyqX0IX/mJnRm0IpHp73H//8GqmQgno3TlTD9
7iaYz7xyeBjOzQRy8+lIjxeFDVuCNwtu9hrzULdC6a330/0JZv/Ty4moeZSC4mW6
PkmHcb1UobBhfDra+LENzBXM863iCTQsu58xVUb3e+FJh4JPhvRkeAVqeh6nCsMH
IDg3W73aeaf+OfKpOS/UKS+jrhiXMBSc4BEBR+AWIU3bzKZ1m2gv615gsvC/Y5wM
QelUfKl0+sVVEOn9LdVX/P0o5G5Ls5XKZcW2rZqM5SmqYGeue92OFVJ+r0q6q1/q
MLJ8Kn9BdpJEDEwqP5MA0Aw2s+3QqoQvXqpMDLUfTWwN+A2Qd9pgPEmyxRTT8to+
cGNFEE4UbHJwZ4I9SY+J9q2hned007Ul5XGqml9XohbiVwZvKBZROpX954XWOItF
5tkUn2563zICptXvB5eYV6dmwYIZZ7OPzQOU62QOWOshMvp98cPXLSpljcpQiW/R
z9rHl6t+AJM35/MfDn5WP7foUUDAfRv8P1m2JvfZ+De2E3WSxqV6TNncJFzhMBVU
qOdkav954iXgFTfIRMbqneiMZpdsLM8bSJHXL5lLlFzDaLRG1wSB85yT00b6jT3N
U1gkkhh46dCzrcxljnRgN+INVy2FU9F3GDXofS6eSSZcml0clMDZkMgcq9sKt4W1
2ZAOP3RIG2J9bo4doFRmqlmJvQ+RPI0t9Wx2lGY8x29yuJ1MJcI0vyn5hYqLs/uV
rdTM3O/cU4auWI0/+LmnKdU+1NDAgILq9wP1Ak63lludie+0swWSOSS4qKp4c1st
sUl35BZaNWqQzT5tygXklRpLfI9tteSdM7wkf1iM4cBrw8NSY9Bgh4GgLnpofZDc
xmcQM3AUK7EEruZHg0IAf//y4q+07Q0IJG2Hb9+itgD2f6RtOVAi7GWRs3oHKiGa
AD+tfy56trK5qv5xHECscC1AXYzDXnI7ZlmUGsEA4b+a8p4p5EYOOd/mURvd8gMn
sT0ikL7Zf9HUHgXnFaLYiJEYVVNPBJiP/+LAKuGWrKjrlV+2uzQWXDq0ojL3Tzpg
rCkA6OMo0gaBRvuM/cLilI3LSOcVLHm8ryg7rlDC2ujUy4fJwg/PG4QU8tNRiA6b
+a7Gm+nUK4cry4WgLQM/PkBX7M1cMv+PXIYkkzkz1b9xOo+JXSvSDimeFyZ8JcR0
z5v32/0YRUeha81M8Zz9+XOCyyC8ydT/TYzSZ+jrEcdNj2Mu2PWwMWerCkDWhbn3
wgIyZKlZb1ELniRRGYqcEMl7neeaABjFGU88W3jYZ9MGKwehjnnjLq9nBQMj3bPD
6WfxkG7LW7A1HlRqWEHSG3YFFilRhykCGuHGLxhXhFWlcsHicq+YOizbxNx3KDnl
YH0H1Cbnb08XOHOfkXyhf/2NsTwzyopHNbNcXS2U05AlYF9AQSfXWAU0UjIMj2yD
LE5BjZA4Vl830wQglFSIRKc6tC0wpWSAJOl5CrlFLht1+NFEzD2+fFNuWsaHn6+U
el/2X9nuKp77nI2rODaX9kiznAw69q2X58klYvIbJwN2slVSXrytt9JZbS1l0QkJ
NlumpvWuqquoyedqzzWcod7YxVfkMK82r3U69Muv2+yJzUk480FkJ0ZeEgsnUXbF
NzSuLp/q2iQofA8Fj3p5PAyz+pGzHTcQ7XHEeVQ/k2KxodSpUfnBJJec84IyDYnb
nKxC0E7EQo1wU/i/XEzshRsGAVOaivZG8Z1ke1SQl1s+JeLTHjXxpZzdnmkw4Odl
3oUlUqKWFjFhKgyCRY0y4q53wYW3IZWNokSN7QCODGscowztYxMzftOiRmF2IXNI
BRCzkymqqmkvFrI/+AfR8aBwZqxspF1Kw6lYetyrugxMihnq6WqTZiWqb9+3YfAH
2JgAPczyQ8jaSyYei5DTTVi4LNXFwBmfusff6Vz7KoKZt1Ynr9TpFL76+cfNW+kJ
fp9Q1YVwi6uxDDsJm/0SxSGL6u4fl+sKIHkS5xTtPkI5d+55MfoRKJLATnyYaUcG
94ceTa8/jPnQLVbci52yA5k9HXwq7BwjR7lMyVmdF96bM2+lyXqBLdNmUfqWsckK
WA6dPLVFj/eyv9icGx82r0WGVW0qu/AqIIAlVJt7FiF+CUDGN6Hyq8CuKKBuJo8s
L2GB/2sROECw33roDgkVh/p98eCZ2rJwp5cntJgnfKdYpRK8ZHwTXWs3535lw7JU
NUMZYpQrFHSGeAZ0Ryvgodxl7dwIeV/wrvp9b9WSRTgwzw8xYNmrvNk0PhSS1zkw
ubofnyUwKrt8MBUs9qzfytOjqxAms1yeJ01leG9xzsUEHvN/TgcrLl4cfsW71Cgv
k3b5sd/AZkNT7qCOV1xP8o7mzJwC7qCWwWP4aow6j37Jj6YRwEhjO7O+bMeXtuVb
k3+OUG7M+SHXERhfXW6w7hZnUoZWDmDf0o+TvVcMaTWFuYcDpiwPTayjwhPXMlmu
Gic/GlucAawvWDJQFX+KkhCyVedkvCXE5FUl9OqziAmfSstndk87P3BE8+FAtOXw
sjmI8Lab5ZEmE9sbvpdThtAF2ojM/ugqlAyPQ8rQfSBsu536wiCmrN8owwdBl/tw
kAfdBzNH4+GJ7av1dYfySiR0zGaCJYD3jolARjbh1x8csct4nQ1ZgIGLRX+Iip+i
lywk+evV58m3AYRLw67PrV+/P2q7HntvQ7rivU10FQGiFmO9p2rw3SoiCo/kGhTx
Gt1DADWsFUTpYzGQ1Lf6Ti7vPIfgvJ8ffA+aRYD+pfKhk4qbtU3CBRyRHtQEnywG
yzj5NEKXf73opgAhteG1vsowuyKAF7zZVSWRYpP+uRg4iS4HDJK8GUkymhBZ+49z
o3n+kNrNnxB4KpGWpREQ5UPZA6xhUAGqB4t2AFwlUEUPOKnOExBaNnTBLwqxWaJT
oGo66rCyJdHF6+6+/8QWbKkKZcIewlRmrMxW0FUiw3QpQhsn0pTUysNAfHwa5ji4
29GDhJV2EX1v1HE8grZutBB2LssLNtwdKODSnEX1oFqix8fjhaV1wks/Fkzsihb1
t+Ysi86zchaZVrFOIbF5IsjfAOtb1Wa4qQsTBfvmx6hDCSkfV3fwSuPyIiaX89m0
G3RU9+BjEn/IdfSgiesUYi8vNtZsOdNm3SdvQOkFQAenAIluNbI2FJFV9FZ5+jzN
xS9nGtfXs5IDdtev0o2MpIKRT06E9TnavJE++aOgvjHGz6GmFO499380qnH6seke
4HYovShG2x45sEIID9s7Kj3m8vIIzaDxMeznr5wc8IMJaGEZ8C1SawwifVTmg1DH
8O8/keEUlZSichXctn8l79C1nLSE3c8utoRnSHDuNgc3K5NHjjMcOqDmKrQejOgh
SGZYot5szxk00SkL/ifzqo/UjACJKQE1Pso3jC0LNOYOwRQr1rr+lY3QDjHjwVGG
eoA8sM5YOA5ADPlav5GGmX5iLVEZDCH981x+CgmVb+gm1Hv8VEzenhOfO6d1me9C
w1LPJOVCprXqppQYbVC0m4HdBxKipg0zOE+5z5PxTf698895WXb5PGFEYZgPgTMK
k64zicNKgmxpkxC+OiypU5lxdVESNnJr4VMSZ2nyDfZfd9Pxo94NutTzKjWNgRu9
7SDSSEZtzcceZCuZ3D+N+YLY30BGEcvGZ8j0cccUIcxH15kwIFtFxs9RK1nZIAv4
jn/8Iy0Db3XPwOcDzSpSdOPuCzLx+EB7sB6DTH1oT9/rcJirSUowoFb+6Inh2ggz
S1H8kLxaKQk7HxuSHbxkjII4nJ2HIojYMDrCxncX2VcfY0KVKiZvIAOsU4G/Mp4T
tvKjXh40GYRlWauYY0/wpb1XChJ+UDdO/YJb3q4+P1YpjwSK9DycZ7p7yb+zULLg
sOGcCUwsyFeoAd7aDxQt8RAyVB39NPM3/71zaSYKV5/KBUYiCZGz7PlhB0xIKUOc
lRTfmnJ1x+NVoEob6CGXqFFjbN1TdYPmQnSctpWy3ly+MBXUUw5ziDEXdsr8AFw2
zlgz6kYScsGGc+xchBLWxJH4V0dJDFnXLzahuWylEpMl4QCmD7r5mUwRRoqQOdQr
BP0PlUPfncWKIYO3GIY6kbFbjM6w264qjrdGImtgBMOUyVBSzVMQLIRs+1AdlU2+
eQxTdhzZ97MOIMTEA/za30/+wF/pB+HyKfDYc1cB5x/ikhqF7Niaawqn5kXOh05Z
w3F2xM9UaTjbgG+jOBf/LTzcf9j8O6kUQKZHIJR8+DJRXbK9Z0/ViJajj3+aUDYP
nZwEiqDisuVP+9396nCRXC9Y4zqWk6OUaRZniObKgf5vuOgHVRkqFdrrf6HsA/H1
NPOaIci4ohbuVmAfp91Kutf4r6fjdjZnbbe7dIN9tVQIMa9dqfpKgj5yAnIIF2n3
rngZx0tmk8f2P1Qm+fLycnrlegIyUlxX5MaKcPvrIBbyqNuyX3jEeAb5//ygWvki
GSB5iFOBOf6LPJLHBx0c/Qjf21gbk/7sT2QQrO0Nqe7uSgeCXd26vtQUkqzWAcxQ
/ZkLhm85h2dRHU814Vq3nf+HL5UEzqAvQNktnf1drZecpm0DYmWpZvdAzmSPMg5y
QzvwJ3LCdOiWWhqioPQNEYmP/RIAse9Scd6Mpr6WwFWBJT2O/a2a0kLV+VWCtkSI
ThLaGxXZ21xj5ooTGzspZYHE4nmgzeYd5yLxNyyamTqRydb1H0hN47FXqcRStnXs
+Ahi1lCHgKRE+MtmGQ0ri787l/EK8itDjUoIAH2GCbR3ytyL6IoISqWFd/+ub3Dj
d/DxEuNbT7dtWxeKLH02pTVOkV30nqhJOJ6wqYj/BCZRlR2qic9bgmhgTlAwkTFT
LU3kyKY3Tk286nKoJ+wGJRpiXCua1qRx06t6zUhigKSpD4bSkjgfsQzI4qDO0xpP
cgBGxcMns1AmhrYtC9qDbePzHS4/Q7cQkG1tAoAW3JmDDMBnwZnmaluHfNWmviuz
gmrAq06+GMN/yUpKA8FyynutgD/YGfN6htB6iD57HOSpW4bbwmJoN/obqm0uQb9V
3f6XlxjKxSIncuySK0ECpgzHE3yCCFXSOixZPN2o1/i7F4Z8Gk535PDNdFx+lHyz
TFWDJZCqvQFJC0UaOar7TKc7DgRNzOicXyvHZxGNFC8rVDkV/CBamEPa2+wFDmnx
Yo0bc591fE3PbGHvDzfHpTbn+Lh4HBlvOzGGj+7wB8Q9/nzcc2D7/9QqFC+gvCBz
6Oznv7LeKdNXrKN0NGaat7ZEMlWcgKpRdlqNbxlE33H+F3FdIYsXdeAqHDnZFYdp
/6d4luxLQJE/l/PHOK4BI60ssltJ6FWHe7fDr8MyomiRYanaNL6k4CFlrp7aciCC
SYZCaDV13PdspnrlPm4DdPeBV7Go10jbXCtakI5aTAm9JouXsNuw5u8yoAtBIyEH
eYyu85JntGg/BLfHmd7aHmill0OZU6zrj6WLOAbQEqnudnz18khAYbZ/L7d7hwZY
JB5dWEnCDDxNp39r8rwnD5ZOsLX1pYine03r8GUCq8IxBGgVI+Pk9QagLCQ6xsTa
JwcxZwsg8NfxIVzvwb+mjF9/DMWPyFvGZE2C2hAeXlTmwJJoDp1HAAPzO8oX7fdY
VL71dACdANtNbjK+oK1ivgxXRy+UZ8eI2yZzaIaAuV+nuK3XGSFYmMv8Q0vgBTwS
KIn3q1vRKaXCnH70RsiM11aBsX6oNJjqyh3vVyBvuC4Hz05OCysr3VvtuqalHx9O
it77n2DcN2YrsOg4DVa9EJP0jRKPy7dPWgm8ZfXz8LDk6D77+o12zbmGatyyV51w
sOppYUNPGdHxljltQSb+ob0eBLQfBLe0cr4qgTHClXC8mecM6GqmEd4NVbv91Bik
3s9Y6F0OGNWq7wZiPhzBugewm+ZDZD8QILXfen67G9vuFGepRbpbaEhrX5/6dxnG
op8khau8pSzg/iZ3YZRPjzIIFDba0ccNLZZTkB4ljNI/Y0jUCr4sX5xENu2X7UTi
HSusckYGkWqWqMa4DbeML0xKJkO7E+kMwnRsy/J80DLEIkGZqqPcGpFLvbEjAvTi
JCsHfBOFKuZoJTBeJbTdiQDNrtR+2Rg5ChgbcGUEOO00xLC1XskIoIiS0Xd00X3S
uwc9bhiUvsB9iVpboDXSuXD5DevZWZ0F0F97Vao1tDuwkw1hN8gAaE0Z9K4ieuLo
5Ap1QcQ9sN81Elw8HPq9Rf09BQ8+NN2u/v84BEuHuwzvS0hWhdyAIp9BG7u8x2nC
bhN0IPW4sgGtA/dXrcDyHrH5gkaSiMVXzHrs/yAJmaNs/bBLGCDRwI7upHZ2Tveb
D2vX75IV59HF9JLn7J4tiUe4E74+wNp0+y5vuma8gzqi7ZBw5FRZGb71JE+ptHuP
PoJnwHSj2jhdU1giIXYbI+A72T+1hTlBO39igiNn2yaqCq9vecKzN0fuE58PACQg
HRb8n0pvpkGG6YdX8bibhMzPC9qxc4wCz+YrmOW7b3lKUdvuEdx9DhVwmb84YSI8
DW0U+k+Ns2W3QYKiZJSClnhWURvQRHBylH3qtJsuoLJLc1+s6fJhY3z9kovHXCYa
JouUJt94ufd7TvDoMk5vTjzfHnad5lX03WLg56el6iEtX7THHenrGCZVjtvxTWTD
7e5BObGADXez+FoK8T7ZQAQQlOoVLELg6qcTT2bEshc2Ix8OJ/+a/YAC0VGX7szC
jGhpelqZ3XyWEOEf3aRcuzc3CQLSU5QSJqWQQ5pXBoiFeuUVYiiN0vZzQ3Nry0Uj
ic3oEFlpRMuPYloVNvMhk1yysMDFhCBlruzX3h63Zy7xo0ijJtZ9uEsjzifpPVEi
mmtUr9hn5DZg5dbOAouHcu5p0gO9NTDx/w333G9MY86DFkTynmOiNPzAqYiat3mD
Z5MIlw4CTeG8En6/ZG2NY/QWWYZoRfyNnIv8gJttGOnIn2Fw1TrY/seTpOy6aVua
DkrK14XyODaY0Mm1CJPr69CnU3ZEt21uuWZFMXSeGdiOxGPH3LAQp12Yf9J4crkr
48TD3l8zhY5Eq3X//uPcl80Sz1fpfgRlE8J/FJGg3Ke6Jmv6kCrjMR9ss3EFH0Wf
A5ClhTqQYi0WmaOVSKbWEIprGJFpgo3eFjilOkxTHT1JjlpusyhFe9Vy/a9KdCD5
YlFXmbkqCGHnwPzqc/4JJSr//l0aXdma8nHEYo+yxv6rAaOi9fULdQMbPzUL9f8A
nUzw+k2w5hrC9SNwFZWHFOy9aNqumf0zOwj1u3w61ObIIGh/caQ5p06qaVEdN9gp
R+Y0gYwgv6zNinKgr2LLW6NUcE1nvQg52KbFtAn2TdZ85MWCNCwGJZSJr37oCPLF
RpDQsoV6s0Ta+IMDsUhzh98xPA7pqbMXfZ+AWeQgG94LtpGiO3oJwa82ygtyP1XQ
fUrtf6kyLbKzlcEWXMIPfi+OzWHQuuXbQzTpZW9uiJKKs93Y98PSjSNdklZhkcEn
Yjb8t7x8b2/ISHsomqYHN/hC9LEafyNELxWkvV2vSlp1VrI4e3o04IegqVNaT4K3
eZ09pG4dypNt5Zi0jwYUHBGX0c+gVcP1K/fJRMs28y7s2Sku+L7QxynTIKcWkV0A
LXbJlyO4aKSZprHya2P9Pevnbz3Bixnn5vJ7tOkFMGP1PFZMcrFwwgyG5VFQlicF
W66wfFpxgDWlswLCQWjDqa1ECZNV6YQ/Z9/+wSD9AkqPf5+0sS6nY6NlEByuaWfp
CvRCMu0/XyN/8ErttUwpSrGn8UUUFIBxiecPGWIHvz35CjiLedM26FnbUMrIWjFu
WDy55jQUlF4eznzbEV9aYQRRjKlGTjPQuLLEPjn7zZKYRbDfpomXxy7RgbaCJCxO
2cskaZOBzzP9zWG9BTNmgZ/Q53Nf/GrWVibcxombyN2zlP0RkUKkmIpSdzHTNfaV
DsPZK9QSPGjX+omVNgBk+ca3s15IIM+2ryNWrQokUEJnxTSWKLmW8vONSHYYCRVx
cD8XIFKMEnp8oTR/GbgmYP5SzXlUGrfBdewGYSRMLlq/PomFpXHwjFqBMkEt6ZaS
oQyLzB/y++2d3oPZrwiPEgwK3V/dXajX0n+lR0w0StPFuwFj/eL5WmXNFG+g/O7I
AStuw+z5jEoo9HLRERc9aObLzAqca0QwMorObOXSoLcokrQCI5alQRWNMqXqPh9n
dIkku/89n/ZaUFvKPaTJMxgWqC/0gynhSGGEoDWPh0v/bUT3oGCn1NguVb60eAAM
xWlo7gEQ9j+3I58J/5iFa/+k8I/YQbNnsb3LW8jedwKEJCvVPUXnAiCNUT7WOtBS
tA01+YriZ25Z14xNF9Rzx4JZ4CPAZVvNXXndSCZB6pR0WRue7qiqgqmPA5ZS3tw5
38UG3FRBBaRrSpLAFeeZRDj51ou3LZ0MV5bzmWX0tDPNJmyg+0hpAG4aZ47j0tYK
bcfnz+e4wittOk3V8DcMcNdtdRV06vSvsFHxp0ven4kyNqhK0jnJOXpq0we8Lmcf
H70BAuiSSrxLKTBeJH6y5PeUfKDRFg9FK0BTe7Yi/A64oKj2R8GBfPniEcCVfEAv
StBCYSRf/gHmHfxM8WvjznzR8epM6MIIguiN82sF1CTiqLbcafVOXeBZ86dZVxj/
dEfdE83gZqcl+6Obw896Akf2/jh1qOiGc8W2rXjhVJMiDxXR+R1e0AM1yh/Vq68g
PSbf2wsj7VqZYU46zb8q28VlaJ/jiZjzTgpPfq2A58qoIRq0mUlmOGu0CV52XsfT
UV2b62A2jF8EiaFprbl2XfmLXInZ+/ico9T/zg+AREPP7yQDMkdBpmJ0T0CdHW5e
3SDwTWT/Rjl7Fylwnglx2Avar0uW2Ed48m8TlwZPj1ms9OQkvc77cwM6VbLksaht
oUP9Xkm3LXX1fb3wYowqySdHLsQV2RLPNL5A22vVWSipu+5qSPdQjtQIsPxXiQfi
xyjGJsHOLmHCeKCPnYy1ZtDp7j6F58TzGSxqBfeQec603gCCLi4z2iH+tX84y7ub
85CL0HFs3TOyGukvx/Mb9TxBqnG6k6uTpr/um1F7Z+8zxlDVeNwdD92+uV7+91Qy
6XGDhfiHyyHZEds/uVDTaaILDWbhY1snWvPUAzl+SMSRc2y9PnJbvO3ny8Z9A94h
w1Boy95Kj4LnGQwj4UEnEj/BOMcI+sLiK8OErUNWX6YVBOxH3RoYze7sj9E4fkYX
GOhY5kwItznSqiU6l4VU0dWM+PHRlWKnD8KpMHRDZ1cuLcPmxvIM+GUzhsvClh0b
RaH6NSgKF+e8hvrdmFfZwpfJMUw2hK/hqwrvxXSEqnqqrmho6xQglTuoIYddjvoB
23ng/l1nhIGfpV5+dCoi0rEt6bgVYggOT6TDUr1ofvNAx82LspRqOn8RedqRi7m8
T+gScG6IRBn/tjpZbImJ/WbTABzWLk0jObjyxFTw75ZeexOdx1jVaHZOOPK3FATd
D2YOiDAr5mcRqBXkJt5L21WUuxuYijDpq/ZU3sbEHCqWpID/Y6OLM8GA4AT0v+MB
riK3P8ikI6d1fTugE7XWvIWq5RtxDhXyX98bNrR0vYXAzT4Da8I7Evbz+AFWjaR4
58j5YEqp32A/XIvjeu+r570TtgXm3Hie1f0TjbP8VtMnFQ1GAc2nUktzM1wheBY1
OdJ+oZLudlsO1ZkZ3h7GmBM2pyeFQOX7PvWdKm0fM0+MrHh6RuFnlZXiY8TsbyQ4
oCjLlBtFnWDH6XMUnaor+70Do2w0/zwLLTwQSI9g4KQ1iJzKm00XFXoqjfVuRksy
pQnTxcksYza1FqjDopXSU9S1DvWF5hta+mUpD82jno2hypuBuHPXM5aLn5ArSex8
bOM787OCQQG7xOCwHOcbqasizezI4A0LyzWPgWQl/zNdx/sUWhMHGWUe1okhZWww
cpO+WpfFO2bj559iAT1RqbRQkKJrcDGMFF2/o0gBQYskA3ijEY1GshwM52APZFrK
1mqVl13xTsQ71UfC8ZTrGYc7SL0Q4/Mr0/vhjc64fVGvEfMS2jGW5JV6hqCUrbgs
q+DKRpjkLiN+5kfbknX1lElWz25sEX6z9Rqq7sCEgb38AQCc+MZOlT5NmENIV5LL
eV3mwChiFf8wx/5p83MIeLhWwBdB8HbpCMEThxyT3R57obFI7ndvDhC7UGkelkce
jZOS4nodZi9vBg5DNYmIvYcE2P7nf5QtMSoCR1mitH/zx8/j93Vo/63hLdFe4G4O
oH9j6fDVSfM7oFslKXC6GWyrR9csfJAJBDo68N4viGAOvXE0WFyzLD2nxflWENjf
EmFPSC1CtRlVD3OnTJCx2zFXMbHhzN7XnZJcuwlai3Fn4z3kY84WauYW8+1CWScP
gF0YKg5o/Db8oiNKberVAIw+5LgBNVJyTzGTaw5557zbWKTA6vdskjHySZzNJLUr
+zqj/Am/DOfz3xBExaO/mjwf1m2o5EqaLWj93SJ99U16gL3bFqfC9XTV5wyvKYGG
FcYdDgnFjLkk727yohXCDOC9smJk4Dr81NLgx8qCTwpsbp8x5WynWsXII2e34Hp+
L/idp5BSyjL974PKh3PmAn98O72A/x/Z+sHj2buWoYKJPEqIyP2/fwQFzrQBi5T3
y00J3g0wcAhi0Jn0Nmh+NQkWrOaVY/MFJ++2Wr+w8WHN1oxOlCGv6Bi6Qbph1si+
f4WNUHgSLQl2iqSuT0RUAZNxBZq7mrm3KoXVxl8n6NA/FNH4gr3/alareKsnFocP
zb70QoQmFttLJqgFKjAcWD+meomY22WuATr6lcRV6i45191yYtYPcphme6VoAAfm
AlqZbDfJNV1it7QAMtYY2otQA24vZQY+WbtKF4JM5ZTzsxC9Boozq7HU8HHdKa79
V+P+PxBmna+vS9sqNdve9ONHsNP6drIA8xIjwlIOL/wKDcb1s1qBeH8uKrshuYZL
PgtQWIk2XSUbB6fdXcSuLpfXIaazC3vOaknfOSlgwdAd+DjGmB49vHEiKbtpua+S
JJ6bAWXazsRuK4Y/pYDiR0PIG0eINLj+AIPG6TDTyvQhWtTkDGbDCE5rM+Bgp6MZ
EJdA0hdRKCiXxHcbiq7lJvF9LLruqLB6B8Os7sB83KcSg+xFMtobJGyW7DhPDIYB
acrMkaG7jD4cSOo8JdqyYvhzY2WY9bOWw8+xfXvjDd5YnJNKHMVnF7goxP/85BTW
mwfHlYz6fhmpE7BkDGFG2giHLH53OhAzH++/SI5YvXGJlSqxwdWeJdYVvadfVfIi
oqs4tb5rzq6OShWZdPOxA6oDMYE6ky8Lb3/14huXY2F0LqvnIdsrEZ17qq8j6JWH
v8/hG6hPvyN4qTqwp0YhOwMcKNF1mSjas3gbQeLFbVw7jjXLsI4tB1FkY9RfBT5H
Ea58qnpXvI2b4bZCcn0Zv1CRBJAfuBDqLHGqC92ALqtA8Anioxu0kA8VAxtGQY3F
bFlY6COpXAtbHo4M10booCM6y2gLjhrfyrlCv5JQYbfaj26jfuBUuQTOIE49ilkD
z7ZX7SNretE7849HWOV6gcK8NirZ+4hNr4PAAS8AV2w+6zkyciwtJZiyd/rR64gZ
eBmEpZGZgbuTH80zTtsFVsMCJPdGJbZK2njB4j64o9wwRxfIyGyazL8C5vX5s1UX
aVHkwx5FtpM0vLrIbO7oli3dsGEZ2ykgFmGIGqdepFmTi96syql5GJy1QvYnbg7n
/fZEWkfhToHXLUoSiGJ5JBegeYKoKsBUkl0Qh7kiPIGTRul6IqNBEnfVIx4CMjf5
8zh7ZsSEirdOOBLo8ZaOuhwd1atgn8oatLKyQB9AfAcHudc0oxbh3PQRLvGYaPBy
IHs+WFvd7EG4JZk7mijkOymmgZPzXAmIHHUn3czih+DghP+bFE5mTl+KvXIXtiS/
oJsNJXJrQv63BhUPIAJFjXGCPrn/L2RVqcdjGlvSfqr3d/o1OZ8S0217n4WDN0I6
ZcbAggRYPMcjGWB15dX4aJJA+g9scxXZJK+yXYra7UEhk9AEaXZ07Yd6xGYX0ZBL
JiNST1GJ0638miG4m/yy4ctxJC96phbqDaKwhUQjuFTs92Cmphesc45P86rqcL2z
BrRGB/oC++n4YB8eiL8VKdY4kRP1gE9c2czx/RHUn3Ardf5U+OQ6RaYLeSd1x1q1
Ljpm05GkFgzrIigqbm5QH0cT96jaR2Y+5zluhtVht99mkhPfTEYmKGJ4o+1Tswvf
MLdqKJWw02Gj7TMRW+ZeilXeHlPmaHximm586pPRxeuon+RpMbajPGJjdIxX77OK
1EV+TDRC8bsaKbk/MEDxeEZu6n8tHYPxKW+WlcvM9GGUp9aHGYk8TBdnzfPJD5LN
DEhG7q4M8ia9iQrJVmWiZQrF7lyFkZQqwxbTpga58PIRY0roohkC/y5FBWZuDovW
tz1SZL3Si8oWtzoRBby64dlPlvkSzlxJAbXrNH0wGG/nCck0QDe8faMjCu2QiIEs
HHLZierNkvv4En8I7U9fCxZo32kKN8o98PcibnihPAU2A9FMphI+so2WwvJGA2Y9
mKqAR+IRCkk0tgKDJKrsICAGB/omr5YHM8IjX1yEUWc1K0QaRkExFodqDv4VVCWO
CY3AtgBSivHo4LBpikLhgqpfnLJzz7WPImqZNcVTe3Gnn8CIxmiwRxbIfr09dr3o
Jlhuezp+pdIM8iN8wBvXOe4yn3zSCEBFZnFMEU/60zfcCT4VnV5qCLsA612mHK+j
f8goKM7UTqCpo266EES7mMhca8Xm+lJ5fHpN6Z5yBoHthwclZ1V3QFUOjbtAKQS2
cGEfrObD5FMknbWfP6FcZypoDMQ7M3/rJRN1kkaAqF2Ss6K6eiC1Ao8llg0KJo7p
0QW0dl/oAjzr7+6V1nGKz2r4n5Cm9WKGIURU/EWE0ZxMY0HltvM5e1hBQ/zt+VNn
M0PWdHqRibnDeDDzlybAoOXedAvkgOw2tIhfXuts+PA8wXB+0JdCaLOtbUmVKlfU
a/e7rkFfryTGdacSZILv7mlEhVk1K0UDznj5EeKSrQt2cz2OkH7iNURsxKWYf53k
VyzvjleshaY9WinVSvuAuEVL6khQvxm9otipGAb/KZ4Vyptluq3uNBgJ1CaDGLOx
PhscfMA7kCNpKXqLkuP/BhfPxVPqyXUNv4E/qfYrGyy6kZ4lpP/uDZuGTNArVOL5
jKDjymllKfH+hU3kNtnHHwmwQd+Eges6Et4JksBN/VrYUah4d77TYXlHdxfZkDWo
cST9RIJUrA9AQ5XgYLJYuTtIsCVfQqs9GLUke5VNFwAzQvQnWmSHMxaeYxRQuhDl
X71CZliviBVOb/IeTGbikT0Rrsn+axA4LGZz6HLsqx+jVV3Q6NM69u51Maq/6z4r
mU5ltXPCWwuvB3k14vC2fG2hbxEEcGeFhmXxENQoRiIM6vxIDteiRjFVJkRcY9ie
0q20yYt3y0dW+bhQ7HqXR22hu32214PhyYdNDbCYuCH3hZHEsLxLHLIZS7RO9mGo
YKk+zKxndoNjYjU9aWZ8N4dUosfkKWesdrSnM8x/U5r3tXzZBYx4NCO/MerWfUXy
BIzVjjwjXvkAHCKIW07fe4/YDjQpKRJZ/qX0MWxNgtPR1QDy22JJFzHET5aA+z1n
V/tP+KeGXFJIeEWBr7HNWIg5LEXhNcVMGd7aBS15Gz0Hv1PNUqsMLfY39hGXT/Tr
PGWck/SRHhOX8qOzzgJna9lNYPKqJOBrAYMTzkJ4NmkOmMfDlVMob0oX0YfXnk9j
oHtFlxCzfxAEOdaclMDMqQZgVuGmmN4Ew7fjD5EThEG2MOEvaevQ7bDVWFLQnlQH
KZYKhiD0IqNFJqgIU3me+/67x/6qnKF+iMsWhWYXRDgEk5U0e2BbS0jSUNIeWGqh
j/uq37L7ajkGLay8Qtfe16AWa9ZPyw5HkfNMHI7mWSctdxCnftj/7tezcpG7KJXU
bKner1jfLalhvfoTPGh7s7s+Egy4oDF1C6y6+7BN0d0ybVSlvX8lhXkgYOluI7c7
1AJgzy3rkwoyAfAPVCe5qOfiPtA+HRp/dn0vWhu/W8Z+lVVHjA+uqR4tMfdcDK2e
rNHNQwjsSBT0GaWvSx1Isp+Zj7ghnmWzO8B98qapnzHhuotdCPRlRTXe0a3XEGNi
1eZnhxG9lVdV9QLj03Pk8b7hZwVeUOkkWqkwEfTBg778waKpF8wWiJ6QURDqCEoP
aG9wsbRp7g+Nn0hADJxRT2wWouFklRLJRYMfJFFTelbRIuUaQYOyhOpSYeCRWuzD
edPa/M7yUASmFGwPON1EPgMIyC3DaGECQHHgVYYqeFB3/B23dqJS6tssmNSefyvI
4IAL5L8MMGdzjSzYK3bz27A1KVaHr9yb27OAgn3XyEsSeNdmvoMYlG0TABXVNSRx
CRcaq4SRtQRoxsRE/d8+4t0g/I8k5vAEwLc2dQiSbOCWSlFxtZAAM0YAmTNOQBNX
kqPvQraBgUO+ab5RS+Rjkw2pSOss1neGxFoQqveX8KnRtmrKnwOhFbQwcXAilE4r
C6mLbnmG2oxpMpgAxQtOBdpaPbyowclGLSPZ6QoaCdofbS+gbTjXlpiT4qhTFaRx
Tqp5lmiH0H5OWVY8FAb/YjOYcs0o8q8aLHJmPKBPNNCqd8bM2oRbrcbP7lKtXO/z
4nH9mk5SPwU+j8gke7I9irXg6AYbvZKNDNpj3yPAX1B6Utt5TF+OwM+WYZz5mFnv
7Vm5hjWP+Ks4VXDhQAnim99a4drbgzENI84RL5fLZySrbzoIp3ahu7RGCx57ay92
7Nr2kcZ6nx7Qy1RP/W/nC/UzakWdHSFMp26VWB04TfqmxBqyG4pshQ6OLcmkCNdS
C17t3TxmvfGwnnbppHcM7CrNOUpf3eDLvysPQTA8jSd4In4ThMr7g1rCX2hf+y5L
l+o2/X6448TV+gz8/tGMLCU4CWclPmU7tLnStOCOGjsr2tkw0/IRHRkCIiRCU3sI
ODIWK/CqpVpio0S/ovezo4tbBWGmpUO2X8Kz+Ld8mKmL+es4mbkb+ZB0faaCH/Zt
q9wDkwgzeTnuwCKFBaBYOTV+jzsejqB7mbq+i6JSM7aG+tsOb82a6UZq/J4TWOH6
kVRH8kzrI2AKulXs+JUx7AAhdE80DfhhLcVkyV5PaVlmkvkIqYLNlS3CNkfYAOrH
rc0OMACzDJXxl3JKNnfl3tP9UdP5Rju8htCO3RuKJhrW9WicQ0t181G4EIhxX5SI
OqReS09+idjho9hxLBhDWQRyhYweqvX4FHnFfvgZy6F2fpkx8SlRMvReRLt7bDzB
ytHwy+O0OAThQKwU7Tjc+jHwCJVIwax065IiqR42Q/6ePZadKOWhaFxLZCdyFewX
AexCtdTRgKGU2LOaDuwYOUF0sACOieSnv2gBhe+/UtyjgmV4u7XY5wLva1UFhcqA
I12g4/bYy3uvYHBgOULnzeerU/2gOOzxXp4LJu9XnEEFw2nEvqQd/QQOrEcGq1UV
DSLkvy/tALo/RgF1xyfc/KPKFVQrLSkMOvRy+J4+eE/W4YCb2AC1Y2gvSEZB7efi
QUIhsp6CPLj9k3LimlhEsuvESOXHDs07N4GZKwQ1YL6wYKeDITm5uhgL1Xh8749Z
Buiqg76vQxQyJTtlgi6Q/r4Ch0+3eeSkbmJa5juwLsvS1A3+fLINX0LGgXIA7qEX
xriMjIGywGxDuw1BQ87HmIwEtQv9yNoCzV8ohkPqU1qianmHnLA52F6W+kITFIGg
HhtDG2wVQqgkoZGVVsGAvfyPlMqdD/M8uY8ngT3syyvsiBeEI0mTZSnspc72aWWu
D6A+0gujVHv7uCnKnMXh3q/HRPUkRAevmOWFdsfbMclih7g/2hxjaPgOdIsHOAgX
adnQRrnrPlewGvQ7cqkUDC1dcCKWfJbJS9WRwO8aZfN+1QV983Bz5SihW0H+uwqr
H7xKfUz9+wKaIJAdXyb4g/fulr3SRJxkCamRBUHgUU48UNtKjZk72fFBYvLcEt13
L6rbO1E5nC8uXyWkrP8bx3BXzbtDryBjgibi6VqLrQ5ZnRdn4TG4LJFlaRHKZU+j
btWpRx8jYjxvo/oB3qjXimT9RoBM62hut6BLWN9W6wFoX4uJk/+irNH4ZI8MbUu+
1D67tIon0WyOLb2mjwjQymXy8SLiXPLHpVVhIKQhkEcJT5fl9K96qwSSaIpFe+kC
eY6bUqpveSGMPAAr8bXWAIikRdRR0DYvjhU1d4rPsSCHuB2OlQpNZSSZWVZxQ1R7
GYsgJnTcSXlN/phm1bU7aPTBdUAjArPerxp+rGwPpufEqCEjpK0ef1v1Mb5ntqHf
3uczZ1GT3D1M5CcusypvLi6LgV4+E/8icFAVmj+o0hguZ12y80mT6y3iHK1dCpQW
M2cLBkgGan6gEI5XTk+sWRehmmXH5dsESgwX1bMO16SCIH+1214JKVFhKLvy6yXF
Ln0X4TuP+BTz0Zo1l5ciRUVnVLursIGrASFBmT4fnhfZXGw+4FXvjlY4N9/dVvMh
YW5rYAl1ZLDCfs7kEDf5QxiqMBgiX0VdwAT4G7cxsmoMc9DvC4+IysFGbmIZczN8
afuhx84YTwR5bLbC1cE7wio+ubhJSp1hTXOPqOdGGnz9Pd35waYeL+wRqVnmd4uC
7gJ05dpKi7KXBQFEBBjPwMQglRg6ZPbepeniQWoYG6gpns98FU0oxEpkr/4KuTEn
K80uJric7qkpV4OGBtQ7PeRJ30c5YfhH2PpSEWDt68N+Bu93g8k7/Nnu47ccXrvF
2LH65oSYhkzT+GLervVUdaOXVeFdB7amXg8V0FuwpHfCRvNasPeZaPi4/XPb94VR
oktrk79CbbGLKOw5qK67I9Q6BiRgWH8PM+F8mm1j0Aidq86q8ebv8Q7e6JXtRJcP
aq4oTfx59/XzhhbR4I6uP7YVk0jMkCvegAFvvGkNigYjrgF4PlB1NzwgrK6XzJdl
6fGmRxIgEqoQG+l5oRBqdXrOPuopOHIXrwMGKtAu1SzS8JMl+w+/cKbRYBu+eUXf
2FUzXe9RnzdwgFoHTenJQ2FppfI5LUdAE/QCx73CDh8FioMciOY4TrSO5V2UIG3N
6nT+/X1zmJiBq4L9ujiMbz8FNCXvvHs7PWwl6VMHwdTCIKbvEHZtmZPLJVUKTVzB
0E7TQT4QSYVaqqGK5JcHq5CoNB1UZMDoVjnReTuEH8C/Dbjo8rpBGpLgQdL6l2rS
YZAhV71wZACxzGkCzRmyGHxh7G6i+jpf2C+uv+T4eK/fyQvSroJ8tdkzCn6h1Cqh
Oq3Qfne4Lyz1KqtGCNSDJhQAq/0mK8hpkN+QsEDMNMdL6mJSeDZ4G33n0NgJmj4/
QNUmmPGeZuDugYXncWUzA4V2C2/76SjMNm78Okpx4lDs9dYP9G5O9Nv4uRZySsZl
XsuFY+nSk1Hj3TzJH6k7iGGZdGeqiAqKtdY1kJuM90APIOOlU0tM3ZQcv+Mc1lOt
xwx6Y3bpin9ol8gq1TuqmBIOB+nTPdi1j9MqAZe8sXrqFPTCdtVDOQB3y7Dip49e
Cnkq1cIOYUtM1tJI/TG5U5qE6Jcf5LB5hXGnTgJPhjxclpJRfuTvMKLpVrdXOHdg
ReHsp8q8sFZqpDFtpD5DN/gU3UQ8h6jX73YgwWmo7EgBWqbC7DApmNUXSOvkL23x
4Qw1jGEy91b4MRmCNwWQ07cG/QpXJna8ZhFdd8kaXWu1uh4j6Sflc55HYIKhp84P
q2sxpR6Pgc+FwArYN/qGWfktj9F785E1YtnSSIVchg42i7hHTwxKaeeocJMN9DTq
Sdr2BvOiMWV7e62wx1LsXMzt6lYr5ehUl0yD36r9mlWIoDU3rDh1iBhJA0hEW1H7
BDkW4DuHa81zIYnR61wHJfjkBWSA2nmVlJceTkjVRC0Aq/fEjbEtUo38S8LnmN/H
3glYbk4YbEloJs9biY3z7k4XiTWmV/HFNWAIilTBAi4GV9AQhqTYX3c3xGPJMUGS
p+h6XMdpub6yR8VrCJ5MJd+LIs4mi/5MLfKP2wxNfyU6mYgYLPxTAAAl7Tf8gQ0h
cTwWe+9rjxF7ErSwNScUIvFwgbEAk4GDHicMTbOY74DXfdPkjcvJUgGMSVCEe2TS
eLTRdqvwxwEtxLW8vLgfzF5xf8QnVq1uTaHw/deU8oVvQLiZkxsgi0NS5FhsZkhc
33tu3VvZWQOfS81Ct0TSUA1qRGqvGsTOF6IBb54d2+aAb4VA+N4yTKTDnQqsIZ4+
FyhCdpQ4mLg7hepmUjnUxDSwi09+21/F9pGlSnKsY0o8G1Xj/iVPntHaRbbQZInn
eArPc1APKFW+alu0IT1HXlYa+6CHUMUAR412wKJalf7xSIru41ij2AnbfC3hh0pR
o+EF31th4bNN8HQKaEZUnR7oyZfg8dUNVtUYGssjjw8vVKD7P8ixXmzldG4DjJrs
Iyl6WQzIOq6pCX5s1K2RDD0eT0/DTJaSm7onjUzXxQJSjVip2ZwTJ7ytqnYqQ5t7
hxuJKBVJHT3NrsWqO1ZS0xZhEm/K7u61V0hWbPb1yAILZpyJ1EZ/wpgtkM7vkjMN
Jcp0KjqGXt+uA6K0YSYDoiZp/t0ukBUpe9yK1wrJWbN9d6+mAlqZD1v2JVNvDMZq
5NQOaQYr726DPZlMX0pVXl+g3Ff/Wtmz5ZmQzCMJXzp8wABJVE+kkXsFFXIAom7T
fa1Yq/hA/pR6C3uLmgjP3nHgTXua6KztduKsjiU7UNPsphF7vI7vEArZSJI/cfZJ
KDDtxdoW3jURMhMnuW3g934Rg+UWkxlSaO/cYdZnDdT3mk/zcphuP+fcnJP4IH6n
VtEHty1YRcVGWHg4SzlIn8oiwOXJEeRT6Quf0itCGgpkyJN4+Yp1JL8MkdB6mgCz
zUxcwUQcUkw00fyP3280OjMbSeOpWtYEKYNvJO6prthqHz+yqHUk2TLYmDewkf8G
w0ZNGIYL88ho3vPQzQfoPZqQ1rOaozZhvE3wOyYdZ2AJGE5oGnIsYLy+2hpti7EB
UsITvOVKko362pJvXHsOlKcjIabi66KFYpEY9y41++VEscA1d7F2lJslo7yy3RwQ
CHeT7qqnuXVw4U1SPqJVd1h/Yt+RbYlnI3delM4uJLZdXhXFnUAuH1YyZo9n/tp0
CV2vHCY0zBORqpxCDLtL0VuJ7uxxBmti8hDepne949e2z1uevpSvr8HdjfxKdgih
O9YpI2MNQGrWdNpFwCRC/1+LV9IOmkzzmDs7uuViSO+APfK3prdqQj5RC56/8rL0
ipSzYQP/YgLmE9Y2baw8CzsYDm80uUlPbjf62sYykSSW2GnXyRLOvbscAqVi/ey0
fJhV06mx1Q5DwaffwCUeM1CNZamD5Onbn1ILeBv4qgGi45QV+NQaGZXFHw23lrCF
AsBQFXZObwNMzO4OIL/9GNYg2qg3EfAB4XcTELCnJaGGxEn6/+okfL2JUh1gZWe9
GwGS/hnhogRT/MchqugzFn4+VglT0+p1PCPCUU+8OF1+IqgWO+4h4GA7KpZOLaxO
DmhXlIri1itcb+SGPJzi/K6fRWL9yMbu5DYCodXmCuO661doOa45DhboKwnxwKG2
i4agg2jzLLqwLIEJJwpq84tsS/JuzH1ARYwCmIHPjKbB5GpX1fcDYx65mdhewZsy
sUS3iv0IEusu2BCVWmiIoFQdTQFQ8mTj/8rUc9/iLao+dKlGK3Jt05SFPSgSXqeu
t2cEAicWrGJ5s9L552cVaSvMfBIwwmvFmDyeNNH+hsiMgva476Aqkk/AtlEZsa6H
d0ljp8uTyif9kxzNxI+E4zARxVcWRV4JgBgj6vqLC9GwHGh8SgATMm2BTO3o8dkC
8TwbjRA2aSdGBaxJe4dNJg3V5i+4eDT/FC05Y0ez/Hl/ceh7Lg6fu6LrRQJi3K0d
DqqVwmt/2UlIBwCtQVhnfxxvpxvFP3rPRBkiFq+RB15Wm/oA7tp2le5924riB3xh
UHTDFqJHQwCXBTL/x5vf0fl6uzIUXEUl3y2KS+KD4yAjgcUYzpIED2PRKWKHnNYE
/hwy66YiDHP70dxYm+w4FOetUit9Ga5jrxbCNynRFx1ehk4XJTSbnGk7AnmJapFb
4EZaT7YBfwDkelUFFH103HbnvmSSI/zodkQmz5fWOC35uzvLh+E74qQpbOlu4vsN
skXqRhGPCsjA+9IxU9Mi16oi6rkxUfjeu0RWdBvMVbNFCuK6ZsR57B1SacbVp7hg
dcPwzyYZWk2K+xs3mg2HQdnVNtfxZUQ2Fji3C42DIvlLHt6qJr1+y2qhkWrFF1ug
tCcTZi6arMCSaA06u0vibum7VKoJJT6JC9WKHeW2qeGQufMW2UAp+v13Xmcs1nfM
afhddVjgkqubMxUJ39oMO/8CKXUMVivpKb/XLzRCrfkrKAq+gsl12W8/0UTztE/N
8LcZ0pMNAvAd9IlmT0SGSkCQQ+qK6LJk4qcNglvx7+/STpOvck52gGAv5jTlgp2V
kY6eOsTcHHqFsbeg9wRMJbEoSZOZjm7iiUVGw/z70bY/84Ha0mNOYacc7dof6Dxi
gruHetr8A2LB/WZZoadOz/tG7A1VemXVzpaVZ/zSSXoTgZEkSNXQfLceBT2AikMA
s0cZz2EBnMtLWJES818UVvvBoNoTI/c0BJOOdqpzPB83Sw+bjAPhOxAHQyBk7tYJ
PSu9eU/I1Kkp329fR0I1D6uZrnMXcWAE+7frgc39evIP82HC+C8BnELtmQ36P+7k
hH6iSDgQhZE2uIF68xpYZAroFO2rWeF9R7I/kw1TeozRIXrJ96urUr2qhEwH5WfQ
aZsZJHOGP+BVg/wocagZIwjBh9D/PlqysE0WzKZs+OMcVs2C61WUW6Hxf3+tm2hN
gYwxo+xfevRAtYIhGUhqjm4EpMM0dwldws72xgT9ohRmbH8YxRqPn9PM5IPMfE7m
WW/9NmNXPB+eVUxLAopJ+jO6Af/UbFOxGrd80aFu4/r7fCn49/opbJgXKjIAsRTa
TbZPS7YEju350tt5HEYZj0J2F1uFJBiMQ+4YAAASHhgTxSCPcaVyYXy6erILtIdu
GEGBbFS4Y6QwsSBtu3H6hkfHhgxCOLcWnnZZE5JXk5MCSEMHAKP3uUJYKEPczb33
FoI2KwslP0Oa/7R6hqrK3wDDTwIa3zy3MVK+VvH7Ex7uzfDUYtvMFDLO0bM7UPwg
aePfZyUt/XoD3Yqol5tEdZQJMSBf2YnL8XVRkyhBXjHvm4L7iMMiH5Ngzk2xpTjA
H3jSRIprw8wbUzvfI2IB5uOD+JBiMhAA47gwwnKJAoW1kAFOIXm2uSvBkb1qjl4O
R0nDQEliKZp2H4yR+GdP6s7mfmX7mPML5sRc7mHv8Sf+ke2RndXrMSdIah7FZHSN
nem9HGkrdHXNaMG9DDu6/OHYq6D8AlrRMJdsQGodeE07Av3ZZnf0ACfFyt7HbA5C
EN+uN6bxA0imCQetKJBQwL6ToOG68QzYsYEnVzFxb/Y7TfAe0iO1H7BSG6d/WqKU
/Op2PWhiwzbTp7DJ8JxhhDdoA0fRUAGCTmOQtvFtGsj9n8JuPBMBh6gk5HqIjseq
RKzFE/1iluhw2zWzNAE7NQI555BrG593qPr0QqaMZZaewiMPW2Vnffb7GOpfQ2BS
0N48CuHLgUdtKYyg4fhSFirJWCQ0FJRYlGLnqv32GuBGEuTwEDlf4OHlaPTxyij1
ZlYh68J71hO0GyyT6NmJpevFA3Y4KqvOe2mqxGT/sIDM5J8iRrVewlREB+0Rmp7Y
X4H2oPG1xrimbD5V/fcT7ymX/4UBdJ2cvMWRkApN/E8fgYvl53zSkiqW1GQ4EEgM
k2JOAcyDCIEfUcIFcBtdG5cRxZ16VlHYhvwBkF7nPalWq10mP5Osk8eWKuNGGkv5
49rLoTSjk9Y2umFRLDZBunDysOQLxWS07Fv+cWZBtFSRuMUf2StkbH6nXSGrUz+/
6Z2oIv/hD1A9fqfLKziVaUeYJzW3RKgpVQ/5mB7VdbRYmiWt3ftS9Q1+A+Lbfwq6
BJqoBSCmsKbsV2vFAH4ZZQg/nqX+qtSdpVxL0ZRLQs0VCIIHEaV52kUl9y2iXl1V
JvmYcy0RgHU1ldxLh0sOrzxeyvF7/BAo7jojW4VzqkMStWYfzHjKFPb/LfeYzOR3
EVz1b1rhRhN+KGb6fI1Wjgqo08dQVUj7YKTKq0x7OYAb7sIUwEIvb242TKfq17l8
LE37dX6b6e7MPtqkurGUoAM8thynYHt+OYk3oOw39uU+DIwsFPai8qOOjJtGOuIK
PyeZSGRwFfdqdj0MNeekZi7lpgUyg2tBC/lY7LKgtJgYCYBBaA/Ngp9YoewcqChz
CHqK7Cd9SM9VV4agkFvVuXYUv7fdAQsl9GOt4EwGW6nbs35aWFvVckrwA53W98Nf
oWoqsxz8aG8pZs5boO4bBAsTPskN6gSG6UXqmCdfIgBggQwC3U0r83eocaZym5xZ
zRCXEUCaEH7PdNCqBwBlXcDlTfJqb9EpzARUqL5XKWBJBj/ywvN2J2XY5tocTwzM
te46Ke8OWGFAxAZBRQbm4Sxx5A/aZH0T9ZjXQsyXx9N+wQWQZsQS0n1+2oN3+cGF
0TQei1dsI3BHZfd/pHJza0g8KVYRu76teR4yehhVthDQ+jlbvQJKwh8G4C81/HIv
rhnRsOC3U2tJhWV81PhlrOC0PCD+yfBRln+iH53UPooHPbBklwbzmrQzFZa7lr7d
GSTEntF2vMYBDWAHGwqXq5qvRiQS4MYSpZ8f5VghfP/VycUt+oJ2SqDyqgTEkbg+
J6YZVhWSaUm+nNdE7RiPdrCMPOTGIaUSMXmHAqWZg2RlXdS9VmQ/90LU2w6BSUBg
V2NXuSiw4NIdyGX4M4S2LwVahArj1rNfM7YNGbIti4cOqo4iXz32fuGVm5aKATEL
zt34bzgL7/EE43oWpvIgzXdN18ntyetj1L11c8u1S6lVeJ+Po/TpXa8mneihRem7
UiskvDIZoSwv3Vc9u5F/rOFuNu88mr4qLqlwkgBP8tLn/tXKCIeAsxlkljTu927g
nQCVd3g+8p/lGB9yhVr06jIVrR3hP8H3bN3kpZvXlUx5LAQ0gxgGJhZFBTKebwE8
oGUafSDeGZRvyGPaK8ZmaNdE/+pEnDlDtCzGk3re+ZSwRsJ6YBMzKRKr82rC0fyj
8DUDJuykaoC1AhaLeXnqTKdY5fghBsXo2OOTCfHO38T6NrtN/KJQXjOuZYKBLLSg
GWMOCSiyLuKmInkE144tX0VCkzpMMk7n8GhPWGz5kU9yG+6afDZabph0wlRI4YcJ
K4KP+t0fM7k8zhO3SuM0PdvNI3Zc/kECIzr1PsKi9lCxB+RFkNQPBNlvp7VkM94l
qT+eh3qjmVXYeGs993ZzxdAkOkJAUNrBHrKCz+Re6ZUKzVUztKJjWNvYFREm2daI
EjnzFBDcdGO2fU6uW4MdCPuqyIwYQf+7bmb3BgjxWplRgrJ+yjT305dWPaia14VR
H0WOClubLrgeEKWyvB9qs1JhHEl01btE1gkjl8O/XY/kvuaTDo0ZzjMCmEDj3UK9
W0YkEw4KjT9aGHboArxy8g9A6p2kD7YPM6XeZc140NvuO8Ig4tf1EfEQiq8Sxq8k
g5wsCqgoNPPxVs8ApVYp/ddtJkMlSMbvFlaXdTj19GNg39HFliayMF3YNdLIcHkf
bIHOdOlahT7S+kM8VopX7eLbw/xVyupWN++YPypUhN4gLrDZ+fHWuXexyTE+EcCI
3RH9jO0G11y3nODD5bxx+20MlvQTowpVfBBzIWPT0luu/E+9PKKpDjSZI2IvbtPL
wJrziFfSOxNZFZOF2TqiQUVbpNG5yb7OkJYuIz3nR84e4wj2WivDkxXCP6dkLjzj
Qc7ZY5NaQJfQHi274Mm/TY/SxjqMgvqhQ+YdWhF606uibyen/+CzYSgmLQzdoVUX
+UBI+bJSjXnFTRfk5PRf6JPKbrAl8DAv3BCY+NWi+xKcvkuD+e4qEQM0AOv6/szM
2u/fI80BX/jgTdL1U7Uir1syz8MVqkNWud26X1z29V9Xku8pJeuCyMxx2udeAGq1
YIPK+dKhyHVWIevsy077i8CGFUUyKJHSYFMclZ9/xEn0FEt/VjKlAlsddTlwoztP
xuvBKr8UrAdmFmbLU7+eki2/FjGk0zKSsIemT4bnl1DHwo+9lt9EPyzTiSPBNtmH
GWMzaZ06kjznb9i59NT/pKJ+oBV84zXvyOBPPdXfU24E+3akG+TU2KHoV+VXav5G
99gnneLolb2QxVdXSUn7QjL/PpYnUVLfYOkzi1gevthGfKdhs2RhFT3czlJoq9o+
pajiKdXGZQqvYExEMqvPhr3fiT614veXr0XE5qz3AKwkjij7HTsrsl0J4rtN5BC7
NgSRKHtS8iuxambwGh8QL3ii+1Nc+cXPrf1npXi4BuMYl3hSuPpQWaKSVGY5+ux0
WnJ/X9IuUXpK7VdO1qzNizaSoaPMZ4hpx2qJoCuVwb4UWkeUaHCcstBdL83Ttusc
7IN+M4D30ipmIE4rh1yJp+6B5CKtOpVn5jDKQM4/UOTp5IDkaN+7HA/vYUymkigw
KFyP3MuRJjkltdEyVmXVXGyOholyZAci18XIjjO2+32YkIlnQCavi60KzYbyVvdp
N77DoiTf/OgpLZEb1G7DxLh4T/F51DXFR+UaAH+o/ceIA90fzuIZz3D4wVXowIAf
BkbKPAyCl7phXjrcW4rN/PuMaKjRLV2tbJyKmduBx8HimE21bD2ti7NohpBxQYiw
r9ROOI+t/PUrM+OX0+/958C1nrTxyLySxsRQDGreASxXjD9NKA468cZ1TuzsvsPD
UMZ2jzKEsRXXOme0Fl2y0072zJlQs0lHb37mzYi9CiMmOd3JmTF7k6DEcNqOfbt/
Ia6TdkS5s27qqcKESX3SEMKW8F4mptZSKCKI/Kr3oI3IbzqMsSpEtgUuS6ePmJl4
VpKsbrYXytEdtTVhSSxyLaZR5iwXCrDAHc9jcc3xg520PVxEHPO7WUbEkcf/6vdk
YCGFeFzU8kAsIxW1NcXN96UgfOgY7CwdbnZC8RCdmV3BpbQ/FoQwDaNlmlqwQGFH
AYLQ6YWZuCVMh9Ag0EwNgGcLV2wT/ON0Kz2K+CojWNLQL9jQODfZt6V5tG1xRQE3
fCOd5J0SLmYjtdGtISLQJ6LikddO01nIK6vpiSXmrLz9dzISdcVl/0kvqeyL27Y+
Sg/2CGq2xhFp71hR1s6X0cOyXJgx7ck5HvOBgdtOohiqN8VQoEgg5Rh6BLja86GK
QnYhwSjXaHRAqaufK/S/CmNsC5T1XLjdjedkNFxSdXwX9JU6lDr5xH7+KAoVcSEO
CmnUYlUJdaMDfFsNghIuuvV3xJFnFFRPCxg9m/cY4Js/MSnQfAA7Lz2dMFgr9x1u
oE0YmoZ7TmRhRRSQ1OuiAeLDkqkXtuaNwbQzQkxLb5T9VkdPjKwXVyyUXcscL2fj
WzJNzmGME94XJ+juNviE3DR17QeDHMFyTq0ZFIhC+eg/lVq2Cz0zwg078G9XM+4n
egnfa1OZ7Bz04KqIpY0jWtuAdTJ3x9t/6LHfa5rYtxWccElabmGCXO7CDGTqSEr+
fiX/Gw7UsmOcRLw6PJBibYEmn6HG/3Sp/zOkb3+Sisd+j7C1iRbzN4RQYkutNgZE
rxA3a9oVqcy6aBfIvRN+2ZcFmVBH/QdXFb6fbOmQpQsmMwLRaNoaYiClpRQcxfsA
qYs27FKArX6oBU8ryeklSfB6C3c09aBrUjseaBXKYx8NlNEhvn3twm1iS6zf2mVe
uLLF8g64CAJI1MCQAatbSdHLU7GPzAve0iqf6gPIWGyChckY6fT/ptl+dVnboPDu
S9MvpWTVFYErGXo+5/jZ5wpLf1LfKN1wdDGkXnK+jEi/l5VsQg5sPZwCu3xBcMG1
LB/VKBYdrqVaZPMagQzGpKL/eIATpb4EZCDmA+Q1iORxweo1sy8S4zMtEOTH2Om7
Pj0qv7TvLMbs+9BsK8mnIAEbb1+B+ZN2WBrQ6szTh8+c5a83jGOvLYDl2SiXOv3F
Q/88lqbSGQzsf8QVLwWceu+dv074uZThvY44MPeofm2/lHPlf30carkCSr2fZw5o
Nj3Izgym1fYh38C70y1JYcTVFu6QaS22TC1qrfw5yNJt5huWBPrqAmV2VuRVOgoc
lP5QBPgsrq9ty/Bk2jxsjZKsx4QviVXP5JinIguKYNKdPGPK8eKJjSPTlsXtoVc7
8UAxqlIkajr+ogPjdbVlRXFPu1cSXUczzbtR+hu6xKSTathwB45FdUbQQBoWAGNJ
r772CdJskuCF5zCxfe+A9SXIn5d8//fffZ5J3HQfI6W36PfGytV6agaWte9pX0aN
ZwSZAHnyi6TP02d+tc0wE3MFW9GbsMqgHIi+febExtfZmWyMYsLrWQt8hXRBAzIA
k0SjgPKaqSXwzD3jYC7xjjNmEl79C1jJt/AghKY0MUd68hGCaqGy1CSA1epIiG3S
G2yXQyExUQvGKS6GYUxJYXbDVtVCSI6x5syX03Eijy0p4qEHluzkQhhFzsNV+CZd
fMnHtpe/apVm4ISr5c+QI/BTXgnoPoKnL4dNrjX4CaOeVaivJvccbNM7CMwoMDKT
60opmr6PeRiS0kmkbQ/2Fymw9II+8xgrtgZs4diB5A+jooidUH7GFK8VUSNOLZlS
58dl+TwjG8RnxZjub1vpCGWuRqh1D4GvWhLVdEM+VWVpUW2JOzFeOF+y4aAxqOk5
oB1C/GWD6UyYSkx4oAvwA/iXzaGp0azWB9Yyqg/Q4PORm861h/jGvNpt8rk4wZB2
yxzNGLdTC7a3WIQ+MdlTCLsveys41tO0lT9DVlLse3Z6oJgKdryGIKOZ2L8OEb8/
sk8QwYDTz6xlzDi/VDUWqoEnld7/fFb3dwRcJmUbZlPe8jR7A27qshYSXEl56hoQ
UJyTk4mq4/mRJKdFmHWoXr2Vf6fGQC+1QYsbgmGsUQcL9+VotTr1JYjp7PA6X13Z
ONeaYfEcr6CGdN6MXOqANbeS6x3ZQxcUHc6B5xD+Cn4iiTjpEjcdxtJZ8MNdyl5R
7x0ZPC97wpIdkbEykYgt1RoNtrt7YBgqVI4/KEHna1HV0V2ZAIScMlRWLJpUaS/N
T7qbAoBc7sgmZolu9V6Wabtr0KflpboJfrJl6cL37aCGddI2YHZ7sAVMRWdNZ9ll
YEq/3/hlGXHOMpqDkqiVi8qpFmI9B29vaxD8X7JdKT1KJ4+7yF6i25/kg5fUrYT6
w4mERn5iMEtEv6blPdC1KpEPMhbGlMIq1jJnJnCUQ3tVZouRVMfPTs/ksEsK3SGf
YYP4U9UwP2wgOlHnmYiD7ib3kjaDNBpi0jHBoqWy3aeSZUyiBgD0MXOqs0SdJpK4
WdYSlCGLmxmSyLmf3zu5eO+lbWpeBc8yTZMyM10w3jQw2vwFoAT3iUHeup1lqqQv
rcXn7hwPFN9qQCRAt/cV320WCHuuIbbNfd+BMLmf7GjrnS4HpcYAZxHeRBz+dW2e
ZywPCX8wA8O9xIFghJKDY7D2XXEBdJUSkj2lCBXYUYZrdJWbzObd/x1ZHmS6B6D/
VumI6HQUugR2/K0SiiEbMf8qGvrzIb4icEz703OwC+FUjUMP3nMzFd5dro8nURk2
GcCv8YC/pVzGuKZ/GbokM6z+XLKaxuUXE4LZJl9ZggBGPqFQELr6z00AXSAC09TQ
vK6kMqjUfdMtTnASxuNDbDo2ug45h8+CPiOj8ki8nhtXtDw/gZuwZ+4IUHefoeSB
geZj3VJyh2KqJFKXFJC4CkhwDkekIuVJU1bhQeKWIIvm/uZKSDrsDnneWLx2b7s4
M3GNrc7/56TITCiXHscG15AC8HideKmU6Xq2huZTAIOClnanoGBWnANd7EVRI2Rv
rTEpsBXLMM07hWumqx6AE6rIUdttOWSQa3ykyjphIIFEwlxqIPpMYVm89UNKG2jz
3AoHAi9doPtgcHbB8mETHgWNuFBznO6RzQ+gRdFnaElRotoxU/ldWtlJUtaD1lWO
OhOOZh5TDFI6YW/Z7M4WffqAVW9jv51SgIvxmzVNSjgIgqHPNxTK3o+Gb5aWzAPc
a/BO8N5wY8LmOAz4SgnI15zB1L7pZFyxWNpS2xzJHliOufRN7Ac1qqnF0vKEfdzu
DgObMIPbLmOu6jGCxOl8nKCt6IN4R3SI1NLLOjHa+fq6J8lZHBu7cOp7P4ZMs4ag
QaoVy471W+GFrxuebcVRwpZINbE/4nrg3rqkYI7fElY1nM6wHdYuXhdGWcXt5RPX
Z4eJlgPXI3PGev7m7X/8mJFJcnC8hmnda/S5ariA0Io5YCWu9J8jYHiPfJLEPDC9
vzZ3uxM5LXoB6FGCvUmCvpQLd34SM8mUgngKH7YGXKnVEkE7cnnXC2TZ7bAynVLD
Khml9Kj01R/CKc9xK+i+9wqIBl/2j7IzKDE2BJdohQggaZST8FtV2PVWUF1V8rKr
RD2Cy/7+ppJVfQvp8wXMhHVoBDoYpM8hKgSixx/4ItQEcle1yj9s2j7XWxOcGnPP
pAu2XyCl4QCTbGlTBbbB6eXPXPTxXUIzws1pd9OuFFcFbrd6IVPiy6LwH7dt0s02
Dd5Vj+MRRk2vyOOXWrByTQk3LSRCL2cCMVj1xi0AgWKjSHjijpQsI14z82Jt8Drn
zgybqT4M70ZtRMjWoQYDnwtsnxgA8K2gzpIJsw/pHVD34qscqtp/YOob7R8m47f4
Jmorhl07TXVuykx5VGREF6imlxoPMYNlF/OyFO/PnaUbZR1FAVb2mLpJM330iEPi
pawot7qTxpovX+PIENHFBWYd9r6Oh86LWkq/U3fMwmq8cxPpSGwaLzQajmNG6qpn
lky3U93Rh5df+Dj2zShvkvLbQXwGwMOqlsbnuUWQSn7jglvJ8iznZX457iUGyOWn
ZMV3cdAhS4wqr3CAKZkk2Yxz/wk658lNAmBX+AoRNqkLl41aCyldIbBbNMnTqEpx
8s18g4+cxcYcmxrpHkgY7JQnb2yN9PY9TWwLZabsWiPBz7DDM/PD6ObQekrGV3+W
+qWJnIJEe1zK8kbvt47eEEOOgepFPrR3UYaaUk+a7tatK6S0FObbyfsd5LWdGbz5
xJGzbfvhZm2V3fTgS/wtF73X41IrG6eT7qpC24o3eS6daTmaf8h0fSHl/uodfrV4
Uj6N57Z6g+DsqKezsaaHIqV2/evkDONeIDy0VdLdGPx31aIVS0b7JNSAmYUSUyd9
Fn6zpKIsjDVhP4D5/KH6qYhmBFcUGnSM9dpG/9cE9zPiGf0v3dnAX1lQBRZmuxWd
BUFr9FvNyXn4+D1NUBvhOY5YaAehYFUZiLX0xevETKuAlvrtzem+pYXroe4aCl/M
sdCwjAcZe91Glz2Twfyagd9GwxSxxQNZ4QKZr7XKeqEB2+DLhQUDA996O473ySKx
Pqa3FjlTHmp+/WMtiKTK58+3lNTIsuInOvejk+z0DUMrc3iKHRLkSRXRIqCofg4J
M6tVZlQjfhvC9zYnkvhuN0z/yj9SSpxGssB7dKm8h+eHvdvWxYCxExcWmHeM/3nu
CbR0i9G3n4+X858HSN68SRkgqrPiDdNquy6MXqbCFmtrdhVcfeVKzqYEyOLkjkVl
biE34U/jsP/Eo/thRWMBT5UNwBKHlNm5g+hoPEpTRO40wvelHIwshp3b98L7zf/0
A7uFzYumqP+DZ1nSBqJ0KFbP+U4e/iORiaSUxBftCnXOckeFFYR9f9WZSTnLkIIZ
yRHRnxBJqh3lLy4HByM+62J8pffJpNheuY+7UZKYIqRoXxBJbeC9M2mGqR5oyf3c
DlufkF8tpzbX+8RjnPdsW7GgSnI3gVgGc4wI6DEuhxHobDq5cVV6wBHxzx492HdJ
WpHOASeV98QU61wpe7+AJ999Bimo3pCa8N80g7bVSO6UjK3VRheSNK5y/myMuHpx
32Ab6YL6vvfmc1QMfu0RW+v6Alb5atYl22Hft14tNvhAruldxIWkdmigjUFp+UmD
S40M1TZzUOlQz1rOjBrTsySn0S5Jph8S8h1s4swWXKlR1D885eyqyNTA/3VEiu3b
2kBe9y9t1g19qmY3JwZq4n5zMQwd+g1XLH5ge/cLU5aIAvIrktKJhcH47VXAKckH
o9cU2T1giKgL12TeN5AzUNYRjilbfxKlUnIM7UY1QX0pgG+VXk1Zs2AuJnKNlTa7
zeWbmla8jJ5HIzjelaWoQ18XbTJykuSov2EEVlTTITZhaih2bJfmhfJmQL/AlfHx
zRBTLPP/i1mLB6uxc44eoOzOJyw3wwWr6QLkAS7z9HfvSqUrw/kB10aVhZY2+JHf
Wvltcr1wtH4352Coz3c20fGGLr4Jl4uTeapIIFSNvVbZ5XunZG5AZAy40aLsTe/E
TKIYjKXHNoFAv/PKQEFIzR6W4X0Z/5KSXKPKHV2egbWeePTkWsLZ5mLCd+6V8yag
i2l64X444CFHUVmCYrlg358pv/lCkCk6uQnTcNAHalJtRZw2xA3cZVc4OZ5DVoQX
BMxFzF1hmrtQOhaKVE7MOChrqZkZJeCxoo2h0YdE/8NwGrbso+KE3iDgBmFDLGwY
KlLlvYj2jpiv5K1bZlojDuK6Ufm8hnGFTjrrvUyOyOnixKvwZLvoCQvnSbSheU0i
IeKD+n3U52SC9d3og17sjktrrQUg3J/BzMMHmuNIw8KpNApKQtB5Ydk0R3+FXZ6y
qZgbBmKlFBTvAWNDf8OYlzagaKZ92UsBhnfFHPlXoPLjG8uvMCS8fy3QA/WbqPaA
oJ1BZJ5fZC9x71MsJwCtRvI1vB/ob+MyRHXZrO8Zv6ujPxSjQy0ZgYefmbauv4PE
WsD8RsykMQRDhAW/wiDrKKOIRY/4eRt82uiMW7hUNziQM9ZSPIgzHj6O+WPOhZun
U93iB6FR8VRcvoLTwtRQWDbPyZE4wIoEXzCirjgE6HuIdqrjcVjIlbfntH/lJ2IZ
jO3n9bn5gDGdBU7F1UzxMtlTVX8g1vVNfP1M3yLOpfLJFYR1gR95GXJag352s1vD
oVpxNstCne820gociN9wUVdTOoBvNiRjvbJvymhA1qiHjwHOaMkkqS+3QkFrsGJK
5QevF9Svn89vaK0rX0x+McX9QyKsg+LQRCxbxilHZJ+8hAPfoOJUU5aGmjjF2Xpi
XhWTwjEuGsYF2RV9NIEB7ocM6WFUYRZ2s8Ou4bSjltR9R+9WJ+LS8njJNpk1UgbX
n24/maaVYeSXMwCayAaFMLUViDdQMUfcSs19wfQ64VBkrlWPagRydKlawo5rxzFU
r+1TWtA2OoVJZQ08HW459llyzGBfKDQe4r8lNJdVnFtVBTrykl+TEz4rYYjMAjGK
lsTQLVvmGVhL5ZZmL+H8oD0/wDzMzqFNEr6t1ymS9RJaraCUhkL2FiUil5R8RFur
PVL4oIBt/lp5NBE7nDZLxDbtVPBI9uituB4GyYoAbVtOVkq0U4WOr+Cz+DgYLddY
IY0gKvm05JoIir2XABurnIYgfBulZsbwCB4wgs4Zu+GzwOKfL9vGYxwjHF7buzhF
4XwqXyrZhjSXqSBUT7QF/G7ZTuFWwfEsaMlrduP5Mvx2ZbauHp+zL0XwPRz4i8hw
q5Sl2xxcecbZ0BgDTYo3P3prOBlNiq5AD/vRnOWmkKDVuwGIenNkZJ75189vgEPj
aahtCZorl/aOsEKwIBLyeGRvUwjvoKhLKVsXdVe4TpDCpr8xnBQape6tiiz3EK4D
bJhpsERmjr3y96Dny8LiaacvBf9/wLovgsJE+SIj20Csp0ibbj2RyKOMx2RUKoXV
bBpcDym/3+DiJQlRYoNcvID1heTSPhQov3J2KBllk3q78JhqYK8fkPwpNOONYQz6
xreyvRxnFJrhdcKiDtTsjfVvHkcsMhiVwGM/Xq06D1YvZu+hqOHCixP4bnFex+EJ
QN0s8VJCsXT+CJsmtr17uU74zpYVQCALlXUNPUcWcoaejeuGS3O3s3zLpJKgQFz2
IyuPgAZaaY84K+z1JVtl+dJmbMGmQnbBfh/FPg7+dqksJn40PPREq3bXSAR2nFP8
BtLVZkM8Ruu5Pezet+/NpCz+eE5enNGPEV+LR82fFioMjdWEm2bTEEtyjW9FiJUi
DVJkBAMuE60GuCpADbVGbyUnVdY+DZ18lnhjGzF5H9KxH1LYzdXz+u/u2HZRm1kE
/GPNE0PYlER+irJTN3WGFcRFn84X5S9OVc4ErfdOenrMERXn2APaAx0v2Ws0eHnn
gt/DRQ48RtwIUwmlgWPzcXNgYWZ1pRNDsHoKf29FBJa0UAWHHZotRTbZhXdh4nB/
Q6tU7MElk2VQ6OtX1t/glbksOF9OgZP2UQck08PxNCTM+CmnDZNWZwtQ0DMWh9uk
Vowa3RweW0KBHK7m2LgGV7B5UfpoyqWta85D89fwCPvBsNwWpc/8RDvVmrCltHIY
HQQ/YOaHEOzaar8rBppcIVsC9hFGhnMDbeTRxKh9ROqnjChMuCL5y9+g7uREttu2
MV3A3U/Y11GzKv+63mPqM8xhVsZgBotGnj6/gXbLQ5Xtdpa53lUkclbtTxFw1CM2
610aQVyqOnRH7njm1fwLDmk8heZ8tayyP/T1/f6CzjrwOwu9ewdx/mUsxBHlYWFF
L6S3wWsgAqWaSoaOUVGwTESEMgHaoKOy1/60vYkR5tSXkf2X6gadqsPowh1OJQc3
a3R8YK+rwlcrMHkWZ855OfSd60IGVBQ5q0wiPhjrkTTwJANLneKXQMXelpPy9upy
ezXOouUbUAFGeOBnLSn5wCiGxyJwMqDAJDHqA7HCsZosgcDV9dmc+3CWWmamjOUo
2fJEKVuAoLvfT6Zesw8lgL7VPbt1XNe7V/3QfkGauM+PS8Lx9/yCDOzIDGQiZU3R
XOQES6L3N6kJSDul6O8GqhnuFJ9X8Z6nk1eijjY0SHlw90L/HAKUx9hGDN8egbzP
OZ/7P4vsxHgpHLfCCw9/hEMa9QAHuxcK4er2QMEZNC/ynld24Fwl26+cC8teSgYP
ugSA/TSUwjR3J9Q896Ey9nHo5cVk+r/oGWGSHMBbxLbZ7SXDLswRVFchkJQPxuM6
zDKkLKaGJKwHGk00tinzt3CgK8OXXWBw5epX8kXNJxNAEM861xDiKgwKPJ+TCet1
Na15UUbbJjN3kliv+FtZDkNQlZZKmYb54lOVugshCKtLc24APnxm3leAXVjQgJrS
x/loGBO2/pDbMh7WjvvuPq+H6vE+mO227dFmpozqy61IFh7FfYAjfSkW0K6pT5lD
C31i2+eBcAjFrlex/GnMmrS9DnGAk6Pf+oWoPkqggZoPmpfmpfL/m1o7BNOag5R4
lN+79PxJesk1taE14N2kdXeWC3H2tcbnADbN5EN0c1m8EK/eTrcOY/BTHCK5Qvzk
BsO1ZYnYzoLk+IlwzXdFxjZ64ChaHDgnjXcDDgOFmqRDjTJnAxIsHVDSHmJ/3/SG
GCs3sDMdj2BfrPWZunTd1HeKdC80crHU3shPSPxjUetCg81IqJNnP8n/G866h1DG
KoAdgGf0jRqWr/1r90zxC/E0Q39dVDo+ljwOEHkgflFvt/KprAWy3V7NOkKnK2UY
5NOfNI2ZhN0LsZT09NfkJb7XcQ8uUdgX88mDRf8mxsNei/NaFCQAiUsSyQ7W1Ppo
SwdOc81/LQxkzgb2FvSsu9sPhgDvf/CBs51/pvNFneQ/QsMvj4jybSbgtMH+cWeJ
1pOeUnlARMMQeuwhRvuIDrdICGsK0HcUky8hbv6bMG64CpeyzV9ccXzDs2nxDB1u
UCoWFHJBUipSkwn1GZ5geiLSyIiuWmCHDl4/fSbVdybWXjuzfF1LKWRm89luDvcb
ClYq89jg/BCCfg1GS/Sdde2OXIyZOLX9AZYWQvOEpgC87IQCXlgSaQJhNsA4WEzk
qtQPVRi1Zjyw5HhQk7m5/9/Dljhd8Qo1+fpRoAfZQzsw3u8bW/s5FxL/OW+NCsPK
ujqUcf/rq2M9Fk7aBmr9naJpcwu/6RD/QldQ4dY6RtFM0q9uF0IQoL+rP3qIYC0c
3UURm0y6MNlnWiFhFVz1zu4v2NbwjMnG23OUfzp5uFI/jf+rQXrL+1v+5g1RG+qB
eASYM1C9lHD2DEhfYRXdTuqAvKYIePl+XB7Q7ZlIFMiu5RjB/w2Ata3h+f3Eno+q
JtKNlHCKI/n4N8qZvGZXXBNA5rhqdH12OPk47eG+/JtIPx6y4fI9XGvmatnKXGcn
wp95xVgUx5AOH8oF48wrSkgn0/EO6OBktV+pE+yQvzqjV4IKs/lwemGV4KoP6l8w
H4hvtfuQFijPCgnS52j5yW91fd28LGf+GjAcZ5cUPIvPAydLgRHs3WSYOXwy1Ovv
qnGr630e1eAEM0RjqckBbZ1GppYhNfz6Z7dU5UrS8xmtR6UniKRDzPFf+uDHh2Bu
Z44N1s60XLIFdfYjD2Y+mfephwf8AvYlDyYL4Yd3JwOS5uQo3aPADS+PgUO8HZJQ
2SlD9R6KIZqbxdGLtGlRqrBdGJ7JpQ3LP8jHtNVekIL7hmHu7uV4h8hpX+al8FqX
mWhxSOQFVbF75tUvoZ7h5I9uS9FUhDq/hWsNILGkjoi3DWlyJGmANaHxL9A7o6rq
QbbYjsTvybpE2c35g6h/mxbkPN2D/1XpEEybc3t0UNuX97a7oZBb9KgNElI1vpTk
q138MheiJG/TX4gXYSqGqK7MI6LJDNMWehYm5W5Y9PQr8j4c00DfHgElpnz+939G
NbjaP+KtX0E/FWtMR0nhKy+R7/gYA9d19VOvKphZ0fT6NIO/ZJeNGPYveMbn6B3U
AXK1hyFk5zwDH5anNZrHZ2NN6FKhKov9Hto0wfREMX3+qHtZiEpTJMUCt2ysXnuZ
DNdA78epkOidRIbifyyLGHP4GGT1l8KOGL05eDxsCsC0jIMLtYZKGmDXGsaVaNJK
b2Ts7ttxo7+Y/OKUWTV8byWJjxzDuHLl1D3JL0/Aztb7+n89SPtQMhyjkpuKijhK
q3PdZcYlR2a9CRZUoA1Kv29asgHjfyFg3otxIfDTVmU+9N8nx53oPHf9T3q49F68
zfOagSDtcn4z4vz0H9FQH9GcTl+Q+f6xzxXcF2rMzKXZ5ZhH4E9n9C7PSeOHo4fV
66OO+Fdrli+JTlYmqvc2nJrR9/vu1Kg/gQgAn0TcxMOk94ni9P0TjhbUiHdgWBQd
r8RGfW3KmouEZY0AVTtskf7n3Li4ue2jeALrjPU4yXPJAdJTt0WsmCdCqhGSe7sv
wLcle51jn5O365d1akUUokx02vm3L1fwlnXcLMxA3AuYBmCxsb6Egc+Sam10zPEF
jrBvLzyAgtMSeCTFEF0GxKPWP4LNOJiOIkVwzn0aydV8kXFOREOWF0hBZOBq0y8N
tFj9q18ICJGVlNxnC8XGoObvUlqjY37VokjOzDRqQ+cCuCZQl+PLTL0M/oPNqZth
2P5yCz/2n4wudQ22HwRW7tspDB6TAYEXdVb9uWUavbTTuMq064ChHfN5d2PDK1NG
fdKW2YmuY/MuxOw/1+P7Sc7VqFKh/zmJDh7Alo1AnKOEwrkVnXstOCCe2jjn2lrW
gTsu8apUM+rjuOLwC/e/zgABSbaiULdZATGE2rrYDSPgybeuMPf1iD44xIq9dCT8
ESIOQxkFSelpQ80psRwhnXb5OX6JHl8a7g3Wyfi1ojweWDQYpXnD7P0z+i8wK9Az
KO8ERx8JlxX6GJpv4qCJ5DczhI8vVm+W+XnfRH8ptWkNR8CqtnD6f97Bw3qJAu34
uLYmmw2ydZYNlgz0MvOqTlcLwpSFqFEKx+OBejOmDRlZkMxBFHdWxvWbGfBADXaH
4L1egVZ47UwpXxg8H7SZZgnBoIbyk97ZefLiu9AEBLZTamDPP5X1qVz4ceghAVHz
7DN7lKxBkvEkJyVCGh24OtvF1qV7rZtBOdHpE3pI2YX4+aMPUTSxGYLVi1LxYeu6
bHAFYepM6ey5BRha1iWdat5VCFEUvgSdiPktxt1IpK/ldAJyXeHdV3qvsw02cvgd
EbGzPV6qWWTOUlRCrH1jSpLIPRxB9aI7IId0NCa01suaU0HLe+W4iyheBYup4kO6
xDV5bnJviBQtEbBILqS+6Nknbzpoew/pYd7kRiyd175IH5iGi2P83qVJ4a2IsCYg
qXa3Z1fSx8nT9xfjw5tnqH0u+XQOO28uJ5t57IcbPpCNW1jy49U6nX57LyriF+zT
3Pc4gfWov1nsxI+g7jfldmIaq5mJjr7M0xXxW0b4SMtazWbXbFUYa75k4KznjRSY
+8OQC2siNxq75bFk5NODfOb/ZhUtpGcpmk9ktHcU1nURH7jB+0ZuNE/HRcGvgdzO
TRg8YZd7SSSN/7dOCyPtSSC3pRCjvmPuG8l37AI8Mm2bWDvb4sb047uknJ9RItHx
SC466r6k33ApRBfBqB6yFRVj2mBQ/I92XYTpqaBgxsvjB7aQRbDHIrrhOM70aigg
Djq9Co/5/D+zN4PtqZeY8Ms60eyhXzeZDZ9HMlcb11buw9thotC7OYlKgsvIgJDe
qltN4qcx6RHqXrLlOM02AWnzbFxuw/VqzySTPKkK8EHEfvWJNKmaXp6FSKi4JevY
4H/XAtIsZxXJ404XGYNQqEHlRwRbS/O1N1DLAvhJOZ/eBhy6Q8SHuUwsVyAJMUb3
DIzbcCautPczr9Fay+LXPCVWqumUuWtRIM5R4bDqe0Bcj1swCnaZ81pliN4aGceM
zFajATGlUCHgX2Y0G3CtLea+BhxLe6fCwXAT29z6EiESZNIL4dJ3V+omWsQB0hDC
wy7Twep65wuztUi32Fzu+d2IjNEK3McAMcRmk3JtepLm95TLsDCXtBxx5XKmbyjT
UaiA4fwerHgl8l1NzoecEhJHpKqPszBVRkLvQVB8jmX6efdwK9MVfe7dhcQiyTy9
kfRB+PAXZUsLkKy1GO4yM+tqna+FrvadlFLxr4Hj5l7s4wqpNDBKPA7CbERDlG6C
p3r2TfpEr1blMv19mpP6hoY1nUpu4ueg2jytzfaWt5IfBk5HssFBmp3RCTLzOyH7
/gN89kMByOFeDAXVry2jQxYoAhwJwuhwwSeHbv9XdN1l1y2LTJ5m354+VDTkCrGj
zu05cocp+XIMDrUH135RZf9r0BLbynDjYDzhkEd8/BrzidWaKRipm02t+5f5TOuW
d0erMLttkNS8exqeEtE8vL32ZYGqVJ4dcG4M7DNIa+1SzKub+5tb/5ysb1jUwyhK
sYeQVCzQf9LbXA6AtaC0FPE4LQawGzApRTQx/aBpRz4Cc2d5HUczmd18Gn/JRr5h
uHzfHMseA9sAKE6EkR1nl8ZDDnrJfoVijcW6zLaYY6jKUEDblM3I4oah98D3XDxl
rXSH/iVGhZGsBNorhR0yAgcigxUyvTVQitpWoe/0cObIV7JGk/tOBJc1gIMOFsWy
GX5R+ZY7G91iYoJgrS49NBbmtRgHo41rtfCH/VGc0vTI6xUfG/eBKrUBYuYpgWe7
pZpv+OdfhCXqMVVYBZHQI8gpc4ymAeupKdePERbF/mItIPUmj3Jnxt1VeDIHsND1
jzvkNE+48d5B4FksipBqxXByu670OxZ5k3aVzbKvHh7Gd10nKb7WMEMsZq6BLylj
+azXTRDki9vu00Ae4lRk13VwD/AuD++wVXkCwmKlhrDr+tRvyBGSWDYfYtrww4e0
mm+6pwnQFyupzNW4Ipq2ke5Vuak790Vz1OsN8gtjFkzlIwvcge7eYJmwYHtvKQvk
BG+lOf8VNUdzu79sMBWtQmcAgSOFc8QoZX7pDcZCJHSGZdEuwM2qR/Q/lLLi9+Zz
dGvKJCjKrjBGVJg8Os5NwwXaXLeyIVkoCzNCcq7f3xp8BE7uDszHZ/fCHcboleFU
l6bjnbSV9yx3JSYsrOZE9k8vOXl6Z8tACjOpNv0/NewW1NvFm75XEjgpYbYJ1D5F
afZiuE94xDtVbdQJ/K2pnV7aUBdX+OX9EhAeAZis5+1Spd5SmFJ4hEVCyiC1Lc5s
R83bscL7QVUW8X6V5Xw4mPln0SNObFnxmqqxz097f6DIHJib8MMXtoxrBhfi8ohI
mVWnDrGgcgXb0KnLtTBo8wpYXscC3XbE7cb7HO5z4BfeQZtDU1fq5fk1DW7Wyt1U
QjL5U7bBAmLB2ryDlIJExZbY//h5Rfhqf/Fp8W8GrotQcmllxhGJRATvEoqnPHWo
ghWN72kFv6yd03vxPO7JHbYk4KCgpH1OOr8vm1t9+OKRGOIueNaU/jA+xbkl4TRq
TPxmOByCCh90OcDkYFOjhXenCBmcFC7bw1jy7uFrJBgB5gDuvvF8J9cxI+Wm+wjB
FgWSHtUw9IbcrNIfsPhYEW7M6SeZUNPKnp2mCF5nxlaygNJJ4IkWoE3rbn8k3GbV
zZPGENkA8/3I1GWNlPAY165JisQfAsdHX6nwTP6LBsnK/4/DBocgO+OS2Zrr4IEB
s59LlFGYfCS/Vb4TACHGmd6afwV1+gshgcrLwFlNfowSfdCU7R8nt7PLSq8E05lp
s/QdrcMTdp/5pKj72mpBJ/1DBgso8r1XDf+ZYn3Hw2ZA3kWAeNAYEkR0xwW1fKCe
AjPLBaCLUaPv4C7to4MLaIw6N7QWIGRJdDzAH5Jw8q1uqsY+VdNnQrna+ACZD+3S
68Vj3T08MLW6PR4nrFjcBkP/NNNvAW5gLjrKt+YhJWNw0HQC7nqpjHX4iYZqa6eK
48SrcXEhtjnYdMS/hCGrJRzmP5RQASQ07TEoGyTaBmTqfS2pz+HgUKSsRSv+rh5H
1Ka6VslrC0ryUgthWrYiwnP027np5sBnc0RWQ+P9L8jho/I2YcIRVlbvTAUYCmb7
aJw/7btEodbOFpw4LndU18sReUEfDDrg/1ijDUFaeUwMqhpeLTARq7qq3O/04c01
UsPsoMOVa7DPr5xXBxHb2ttkVe07PUzmioKHtmkUdXY5At2ABb/VvCjUO38xwIaM
9EHNoXu0JZd/am4diUoct6kUS9NDvyARovfBLDxh9/doQZviruZ05eRNrnjSH/DC
h5Ahnvut91fc0gtl+IJyeIxq7c7XaasZP1T5zwpOWkRf3VoZ7bqhq9eosN0LzwPE
rtMxeR7Q73+D4O+IsMSAK1piLomEhwIbXvlrQ/+bt4T+pGfCXoiAJnFovh20CIFu
6eB8VQY2qIUl/7XVmFc50wXCFO259gf7CsHfGVG2mHBqHwh/8PPIsGlff1pabWYv
Db3oqsoVDeBPznkrnuOalMoqberERfLhp0A6PWzybXGzdjYR4WhUZon9k2Zb1ttA
nopravHB5StlGmzg8Hf2gWIKVKAMH/yPb2nMpFT4c/e0MiUH2B+C8XFrD/M1O8vo
DVKVhPmIrJXrTPzvB+wARxbM7BdHcXwC7xqNtGUYwK9DaHgQz6HV7Iw+EvnVLfyK
1773Qb4mIn3HwkobzbsmJLW8nb/kTUY/ESesHfvLx5er3Rpzu7Xwx4qx2D+7CFkr
TAr0N7WKhaAjMPDjmpuD/jX68qz1UVlj7A0HO5fKg38aPJ8arxvu3950z/3CJzQt
tPwyHIpPqIAzoIfc/4MLk6grZbZYpNzsUAmewbb4W2j8Ef2FfktxR3ghvIgHlE3K
/GqMkp/eqiEhmbXc8JvnWL+hpxdy7uOu48bsTc2SijvnHUmaBHCU/HzwbdLOrQqp
tjFGp0VYBoVYimQtm46V0JaD3gOQCsnCPMauJ56KR3yf8f6RID1/v1xWij1tfnbF
YRH6GaJcXdyrFtJQnPhm3IrPUlzdi3o6B29ButZrl1hfeFFQNgHGPif0ji0fAqaT
upDYtaGCCez0lGsDJH0KpAyoS7WuXtYTuEdCe0Gh52U91uVNhN/WcrV6WdQhe/pY
P1jo1jMzRrP1KOSstAH6IT9oX9E12qZwLI2hFy0fcEusrq0EKt23Gku0eUeATAka
6nEujl8OGkkbmeS8F7XNrN3yaG6emmQhdP8OJj+5nKzmCRTC1ehI0MKw09faW99m
wmms7dPiWs22cnmdwjy2cEGb0varvE2Cw8Yymy0XU/eS+j0EQo7AWN0/0oltgyXM
NEU19dzMJYYleLKSf42wEDUuC0Q+1dRwawmbxGEeD8/vp30SFh0ku6q6qZ8IWjfD
q8Urd4vrWkKKpB8EqYnyQIMs1T9iRf6Xnq5UEHpH89qcO8dU1hDD+i1OyAsQ3OxU
ghjTxM2jfsOYwGttn5cDHf+MCdlWY7/sNjeMByXj6NLskIkqrwsPuNdbgG09YePr
ajDgvi8nH/4u3iaRD7tcWKzHCtxL5zb3+KaAtruuJradLW9UVvCAnVpV1LOaMfiB
IbCjeoFOIFOCqZ9eJO3JzM17OxjMQGMKJcCm71OmTRxiN8jkMNPsepUjbPxHMWYQ
/tzPmHdE1AAaY4UgVSxqNkVP+UbLGeq0nrJMpGui5vgntmncv5ZFRFYTAzIDWtvT
nNV1Ve0DjgZSZLjO/aAqCbEQM09OpbhVB18vLY0EnLhRRt+XKj+AjiHCmPIekyM2
pbPFA4+9Wxsv69QyQUtOCBe3OdiQr/ESPFTVvfaXJHCmJcx8Asfbs7IS1RLjBq50
hDzFY2QqQZ35Hv/T/oydYFptbwdoWxf4rTvednBf/IQhjGBbhe0FYybin9L4iKcm
hGcMX4yzYJIgVwqLaD2juzST4wzR08NI1USL5rmqO4GuiBVgnFDqTK/SL9jZHtgi
YqPJNJ7TN1w5G2sJNbX3OoOd7sCy7GPeRxWtcHA0vfaYuGtVfaD8L2mL/U2ZwrVj
eAoDVrp0Qn4Y5L+WWMZMEuAkewXLPC81VYN7qUPsKaIgtwKvgmj0WixgrZDGxLrF
QNaVQ/c7FSqiDtAXDkignXXMVn6t1DM5N1amUp9R3YFD63OjWYhtBaQDcxZDxqN5
EqFtHpGaEqvdeqASixae9mH3ciok5slfweuvfT0VGU/9J21/L4VQqpJCPrjzc59T
332v4J3cdBLQEwn1cY6jrhNoWB/mprrgMl2KXsWB8Ub6D9uZ9LxR2i8DYz/Tat5v
yc7mxYbXJRIJYBM0fqqsXH+TJRXQx0uKhh6VrigbEwcWL//LehC8+gVNuXT3AcPM
L0qJWRwolu3dxCS0AR07P5Hoa42jDmDMDe4myb9dKNRksggBh7Uve4saN0IZmJdv
R1ScXhyGgyMX/GHGmD2mlXh7QvuKBJn8rzzWSOD9LulaJqqMDgDRsaTI+PWe0Imr
IEtQ71O0gDWjKoOVI/jpD9gMV8HY1frPgJqBm4pT0THmcRXPu4tmeBPxvKO+LQOK
7dUF6Vq6h9/7sZC/bPWUbmqra0omeDJrJytU1TqCXNO9b6Qe1U0DGKIcLWv0Foo1
SAWN5br/cgS232q7PEYK2qZ1ozBW+ZAkl58GTQfd+oJwx8aGmk848nNUWTfew8fh
JsBTjk4Xk7WObnhAYTee+Uuj0lqiBkqTF9hVIVNAg1p75kF1yClTEUK3iNRR26H9
ihnzg9hRSlSAlnh4nPGQtwtV9//j1tE9l61ufr87XvaTMlX3dIkGyxQUeVCkCRoS
mUZkvzxNU0f0qkF4VzroLPO3pmA+s+iWtQ+EDEPpThZLu5TcktkvzSqwoaRc6jBz
C2YSUzkNgN36N5F6o10F/936MX2RxXLIXZWXtwAuCctF/P/OIk1iVmuBPpBRnG1C
dksRaK3lKbOJ9W2N9QClO88plCgFUKtLiguZRBb2oshN3xxkIaR8FooNPYBgG9i0
IxL4wa0jI4yLkij4e3JHl/XujpRzBE6nF+VYJ4H1wNyYimuHhZtjZELTtFez1iaz
jfPRauDn/z+v4uj8b8oMYzja1yNaeT5teq4efpei7fUwrkNFie/o4IqYGEljRfY4
JE6pVaPkTkiTPNJ8dasmnAllIhY/5uCvzMkAfqqmEls5PmejxaJ6d70Bn0hsaOw9
bE0k6hohQdp3GiuZU4Uln0XAP8p/Vbq/p1DxEBdeBVlpEIHwi1TqSoRIYP8zSGDl
RitI0FoOnsCITsvUMehGMJSxjWbqrPjpkgZUVh9idP3pCmnFWONgLHqsWlOauxOZ
W55QcVk0TWqQ8QXTUpaRHBq52msun4L7GjLrb1JVKt9TsBm2h3QRs2hutKAl/wTi
9ft2BXOStTh5A0CvSEipy/Wnot41wwPInIiw99zAf1ex7JVGgi242vEf2VToT9nH
rc4pyjK9gwiypmR8QyOsT1AjvE5qY5cTyYVOxH4Z4TL28VcKT+MLfWMV6PlGHf77
RcDW1wlLP74JNyCd8TuKIDP9O+D7u7NyOJPjJGjfRC0a3zVmydmTm0gfghDxoFvl
x7qKKXaYgT1PEK8TVFgVpHsbBFCjTgKOvzo/uJpyxJ6nWaa73DJaY+eL6ujJ8eO+
RItVvhz8KAKTWVBwHP8lofO6X0UNxtahBNp4XzKaa+/u/mvJO5F2DUz8qWnG/csS
oSDeXOp8IpmOUiIFtnyRiDhSb2qfohR0bMHiUqEdJH832Am4YnejQCNWRs98qKft
Y+yfVxKx9BNvo4TIk9/ZxxGElViq9G7Ay4wZddLywK5tsAZG+K8gnUYxW8puUig7
jVgpjvjSuB3e18lZWA8lBpt9SKWV2b8ACraMPDSiFcrgoZu/dJj593XH4VGVJMDa
RBmKPv/f0LIORWB8FVsPzI62rwcWzEamh2wkfvGdoyK+4Zlx5CwoqtI1ya+VLYbp
EnkCMZ37X8ckw6DyRBm2zEqCMnhoKMvgxubniimm/Y8CvXrmjh5PGm2XlSJXfaVD
2aQWn26eL/JbTNjxsLR7Ykbw1rfRnFVKWYiiRuyG/GaawxCAwTXVr+ZQAScyezOD
y1slYz1UBrJOY3+03ipP0rTvFzhHRojo11aS4GzN0a+uqhvpdqxMvsCaex1fru2+
+nqZLj1S3dGx07dQ1dhZ6Jakc4w7icKi9TPX2FuLPJXJTghlj0Ui+a5nWPn5nzUc
S2q70Th7SvZcRllI6APaWBc4+5c3xvBEl9Mcd8Zccfpe0mXmz7XMKghnf4sCLoPd
v2vNzCmuaP3kr96VRIY2qK03jkAmVdD2ZTT0+9ETpltG4zl0//RoGetY9/GeVo+z
ljsJSIISWYoYilQ3EPlFra5D2h3HZHstVG7H6X+YcTtwf80q14BJGLH4wwit5H2x
w4Kz4yHtLpcxOOWsxHdjz1u2WaFRnot//sP5bRzX1Eavp0KQ1LsLF4U1PN/llL+M
Eg/DYrRcxGhL6aePvClJYLqBEmQCHiMsP06wVHcVhK3mafquV6q8QZ7yIs+4n2pa
sBOw3t9q+nowvNR0OoaoZMT8+Vcz/dZmwuJzxAC6uKjSgUHRFJLE7Dmvxgbjcffu
rx2mmHmVgMotkywvOFVc9wGelVBhr7gYrQGz1ZHE2uw7jr1snta4iAB77BcX9ZfG
wyYw3FKskOlKRc1vB7LJupWvv5FQutJ/RIIgQ9gybuWTDBs5ZM6EQcT5fgR8s34Y
3ECg19Zjjs1lqQ5rcAKfdHi4RZYMiEt3FJaSTYRDj95UP9gNovcal2NQMDiRrl00
uhyLVyIB+ibKpBwFz/vSYvD+hKsaisCeITEhxB5/A96EVCeGwVbRhGhz0OiA4bF/
LN9F6nPQnskYOKdpu0enAfKMJTVzwGQXXtlKhvr0eOqPmAEPMt6jjYoQ0ZwoC5OL
+hYRN9H6jwt0if15kITekwEW/NkTPqTtjFu2CYC9+MuEntZuhfygabgIqTQO1qOh
6n3pCelfoHXDmzpMvsv90VfniwFW1kpTJzoTgWPupWXILla/JPad54n0111McsVj
zCTkFuOc0I8dXKGCn7HuY+oGch06fLz4rcQqYCjfPi19is63U3+NAoCNP1R/AGHp
nkMZqubvci/VI5x82sRlA+QMArz6wIoNc2REhi+ThTJZInzKiSzeWHGtZyoUM4wZ
mYWY96zQWjcaHQ+oRuydCOcXEYMXC6BcTEr+uMylhrhI0FLbjjIlOPV95cIAEM6l
UuqOxHLaPu90csWXowcYMt5gUwUb0Sdy0WZNt6hPnE1j7QQIcATnRAseBSz1BP6Z
RxbAmhBbY6MEXhsEL3h0oChAhtmxQEFABKP82ae4Xi4784Tq6QaU8qLI+5V6Xa3Z
2W1hjf/boRWQnPl25hVHqq6MEGKj2O2n0MjfG4f6T57hMjwaDWAewMe3rMF7r+jm
ilfq1PL4x3xKjNBFiO1ll7WCikvq7l0L4ku0G5Yw7zdz5M8iPyzzcW4G4GKAna2k
vPiAYkPEgYMX+0FcClaIsc1WeL5fnJ9QJ2hbPpoycnBv7QcTPG/wxyiZGvC3vslh
cz5S3r37B7/9XJl4m2VLl2Yum3Jd8h0FOZ9+hKmlH3X5fQkDUNFwGTGrDaEnqBaW
SEInHx8guwfH2f7U+vL8YwrGVvVnIm9F83A0bwyNwEeRu7QSE3cvf50qCyTEANxf
UdSOXSzfwn3Ig0GINPksUDYVfjqM8pxyP9KsRsARtM602cqhq2AM8o6jp70F/zEw
Rt5hSOGiWVD4Gy+D1G2x0BEoLepvwkJ0hniHdxwagspNme3G8zAMh11xNQOkd8H0
LOsemVENhrHvCR/wi1GgdBLhml6vVxT383vSyhplRICE/T/lan40vetDxOMvujSo
JphIatpzr+Nr1STEK3TrSLv/JkGxAd+OQy/zSSOIqo8oG7ohRTvlC3OYrGJhJJeP
C2TUjGTkxpQcSJEP4RqygVBryxAsNN2mtSal+hJCPSVa76/kTRxNCfs5atfME203
K/O3y2qFak7+XKUQp+lD078e/lhdHngHYhuR5i45sPXCio1Tej4Zmy+z4C9xRcj/
4BeoKiRjbIIf4KPfpmwQU+jGtOR/6JXDL6e144Sx7LwQer5x9ZowW+6BZGqSq6xx
tG8gSdQtH+IKZDVgC5otWf1SYuzz9ZrkZ5wwub/SmVjdgop2qG2ZrphnQtVUyeql
qamed5IrAWDQoN7ZHpCfFNTL6cwy+YVRgsRwoEMKqVR9K7LLhY2CF4GW19KU3dqy
j44cmEaGByCXepq9UGWQIZwA6ruNYIr9wVLC2zKJZBWLRcacbDxX+G9KUtxvtYa0
tRHdDuDW3XhodTvstBmzKI+9OszGfiiCvns5JT01iG6xA6NV95v0bJ+FX8pYmohy
XPJPAyTTkId2KfG/BX/6JTZLChvzfCdefZxWKxsF9zm67SsPgZqVPj7kA4ROz52C
JzWuTFL0HlEyFexuVBOZW7AyuW6PSs9FobvhLaAYTiQiuLnMjCOWO8YYIsi8d7kp
DXA5GXMuco3Vql1DoPogXu6pECUlGrMTnrOOdeIKjFnZE344K109b0ME2anph2SV
Bk6X4ykTFoRvPyvJ6NMzU/m+3KfLGh1Bx5fff8rn8pusiP6OOMma4mCtTzdfhhgh
MZY3Bv2yrr+pPwabNNeQdJMHhzQ+Ijv7dMVzrMplCX0NLTt+lXu9HKMHtUJ7Zkgh
ji1/Gy7QKANvV4X83G62wAiddxtSg585qXcunQUVehg1fEMB2S0zW7Mw4J7moTGG
M1JR1b21IlDz3tVQQFrDMM+FCLf8WLnbycQzvaEQihJJqdENmHemjhPlGJtUwDMi
QGGOuPxolGH8gl37iq2l/XyHwCO+BhHC1Z5QnUZ2SLpLnDE4mMS+fiHoLGc+Bw2h
3S73lzrnEMFWoLNiafc9T5HC5+lVAQNSh0PafV9XiVqQ3HuTZZSeUcO0POBf2pGY
mbIH3OpDWnok7O1q2plfmLslyLh0o9LqanlwNZ9pRm2K6p9ubArE9Av6MbDS/Qt1
xTFeLGxDc2pqVxsa4MmTzbTCjQcK5OBqEKv+Sof/v38fJo3ZnAybVS/ULOZgAsPJ
5i2NaKJg0PTX5ftfhkL5yuhziXxJ4LU/qv1UjaTsxDnfae8pG9VV6v6+ph8SJEwm
utlSpaACeTQzOwJa5NFhDBZMfl753UPiWJNbwVo88h4u0PtjeHFkIGpqT0Koas2C
qgRcXCAxpffbWO6iFkRerpX21OBPPo/xXFfutrB2BmAsfrCjTnv8bESOCWkQ8/X6
B+xyERbc5KVMXr6bn/QPxMiJ2ZT+6VCzwdGz+nZbJsEyJ9U6JSb3CoXJXnGYRt4S
5TwvmPeWsm2Q8KrX+fp9PUas8FJg9h/7KZR1CmrHoY+HybvTjrKLN2mgOUvl5ETA
VHKXLAlbk8pDJ+oDccqOZGS0ijoKh2NAL1/ltSmpg7/xMRy7cvR7So5fIBLKtYGv
A7aOFdWYUnutIQKP5txL5ZrtGyY8mjMhsa9dYAQB6imPksVxxP7Dj80lAEeLjIbQ
yMXoXgtBRp2QURKEdBF6oOuLjFqNXGh/LS3ENeT2b2I1BqFJ9da3jVQtcHeQyOU4
yrfBUUeGxyKrL1AKpPueM7+X3r+h5sP2CsQTY+c/Qs9UgOjMpd30XkEbonqeKv08
1ZJUzPlsSWs64huayFm1LpQm1QLIo4nWMNJYWJvPVV5cRvUJNvuuAz2TBbrZujUN
0q59gcRaLtiBVJ0Ao/MBmaG7z0ckw8X7piic1lg2Qm1N6cCTGntHLIslkiklsBep
4zrs6TZYwiN/L+nfRYMKwp7/RvoXof8ipGEzbva8HwzPON9gNbha0Y8285GAZfTL
3qTDOIcmPTEYsLWfAqIPRsPprrzquulagohFNtPKgIjbGb0J3weCSq5yh/pPfXPN
Ko6PMfrft9rqA7SvpNv32tL9hEUAFh2dCek9z7kk5hWm9TTVmF2/H5TEgwsB+Gue
Gcist4UiNuwi1MyXtpPHBLG6zhyyVV2XbLgev2ibfnbevmPwRCM3Ekv/Lp25k+bJ
IZIZD6cJPM/Nsem+wAWZNTm0iVV2NgoPmrx6sITB3rRPnSvnqEoDCOAI35Gph9QJ
vLDC2l67hUKPczLkvYntigFaRquxuw4Y02qxHHuklVaBTDFSbAIqPFGXP8NCFLBY
L/nsUP5cQxgOzvN2WVRe63S22bVJZ0dFDPohvf68ag5vMgbmtT0xV5UjuooB8Pvp
nQHNj1kQ77JFQn1A8vuKJrtTLhjnMecaNXuGdhlBJEGxVD7OY1w1nRW4W3J31B+F
m8HoebRlvUGLjPW2jNVuLp/cUUOnP7jDV+PqryqdKtZ9nkUH8H1DqKh8Ev2zWAWb
E2qCqKWfxqvifctuS1TIyhDBx+fhCmITD+Mew2mDjZJG489qSXFusz3SR5p2/TaW
w9Ui09ul/EcG/eov0EGy+xamIDUusgPxhgoQgK8+tzvYmIf7nkhXzDUhW4Lnemzx
nOYuG4Sc8ES4c5Z6r7EpV+i2Wat2tuJZZ3Dyk0ds1CGFllqXjrmoLrGU1XK/cfrx
2q7dpfEXLLSu6GKKKCAD782pcZ6O7H/YQ0c8t8AFBGZZqArdnHHlQLIAY96UiLTN
STEpqVX0BFodyX6p4XvMTaUyej98kVbkl7VAgvxuLGum8XttEguoDepRgQ+gm9HQ
/WISIISqwMOf/9EuQKtUXsEOxJDZF64MCcsL/slgo2qbIBWWaRdunIPepdG6RSnh
77tyKNyChqmppVbbc1kyQ5oqDC5LTwjy/RlJEw6C2vIrmxRO5jNSxd1DvaE4a4Jx
U1FcxsOHQhUId/kW+V6NeJ+NE/LDF1Q7G9nxiBpNsHuiLfrM6m1izl1J8VD8yb34
lYyWVaTjSO83sPMpV2s5gd36Ss6iblHr9lIAY/nWk6rkL8twYFUUeFx1T1t/EzVG
Ts/2WbpF6+plg6gkx1RXm0Ys8QvtJSQ4Hr7a87irdO8eWvulmCbdPXruqtHyCEsT
bgTRNVVx35gqIO5ixLtuX+28syafGeOInw0+64Ud9CQNcV1w9COtYumrauVCax3G
+mTTqFw5xVyF4iXo4afD0g734tI/iXxW2jD5IbkniShI9iKTim74jjmOmOkNIY66
RxwRySowYeH3s0FjVovoQHtNuRvqWs2i8p1hPeHQkQ5839//Aa62Dzs93y5Udjx2
hudCr0xR52283Xj33pgvhDnGpUdhx3ufFv3+ze9pS0AzoDzOBDA9KAd+jSRrU+u0
Tbf9GRH3A6aqoLghhsP4ZI1Wn9OgGHPB+jId6bRViobuQ4dVbOvNi9D4jXDaSlGE
Dq4CIquIe4DifGJY/nBkyDACbMdCPG+WS8EdMPoWCOLLYisjC0/BUdADOrNRLvv+
sLCoYOKcjeCWoDlaofNj6pn7YKVe0WeZjzhlLvxOlMUQrOgWLcbQLOIIzTAPpvEF
4wy7/ycBzW69n3+b0VUMaqJ6yL7HI1ZqxrADOifr8KfK7Udxkw6GbAlcNvBp1Jrv
yGAfdPnUdh/VrFDZnU8r6cUzHJIfGabmD/1caeoRX2Gu5SXaEPvVN9tOkYBBJVxk
WGRKY3yL4bqThyp79B39eAr8s5SaiVddRz/Mcg1Jf7NMhi+51i2Q8X1LUb/HNzLc
iICGz/yFlo5/ZSBnDn1pn1oiZrYHWzI0twqDkR+tUflA3C85lbLXOFwhdxE+80rz
BxotHc0a+pv03WybuYHVu3Wp786EO2wcui1izlyzOM8/V6IFcY31lq4A918E6K+X
1qJ+avt4EPoAb29vOTSTY0gF+9THLLQRXHzwPoxZsDqDcOW/p9Svt0tbbX5LYShH
noI5EIxRmEbcGHsTExZc6ZGHG9l2/YwGp+wrvO+36+p94tN69OtNneWsfDTiFCEw
PxIsG3bn3/QLcuDMjEiaeM7/R60ujBEmA7gsEZ2eEL2UGSCN6WvCTqQpG/oLqAG6
nCX5PtnasYQigp/OpdaWX3KUXQo1vhJfk00i/V15ECp4wgQwuO1ifX4CkBM80Qnr
LSt9x4GfeLaOsaXLMKUBaf6oWVhySR9NLNy6AdqDH/f0443Bt+uZPNI00nUkwZmk
LLnerHS6KBxzZLrOFrsxhxTHcDvrz/zAwtjSzCOsGe9LPdORym5I3KGRtDHp4ngR
hpBVEX19CHvH+Kxg6Np2wr8cg2wpFcHePtlOQ+SVZgdtoVb0jottJUnzPzHTxZ3r
o+rho/rFv5p/UyBrO6RlpD79oO1AjQPVpz0U18yWnMOnrv6R1fVsfQ7R+xxAy7PO
bIwN/5z4L+CdfG+2zuu99NRUbnj/A49LxQtk1U7ACv7UGQOsz7ul/TrBU0Z55Yoa
Xpm2FsvZ9n5NRcck0RE1xqrWB2VuH3KFmDnKbwFz59CiJ65WE0mxTFY8d5zCrWlI
xpqigh0PIAItb1IRZ7EMNGRZqfy33g9o76+jq6neS8ptMEmkpOFL/D5TgHcESLdA
0K6KrvFSs0W2jKLXh/8bXISObIYbzxfI0cDh3v23VgtyAWubo4sCBUBd5FU5KqC/
qcutNaGD0fa9JItL7qRbqpKRzTRuQ/pGLY2OO2ASMmNAqOJghlvIYa8twjxoLXDi
KOUuFiIxg7ZR98uVzfSXMfMPjJs9iJdumwYUqDCY/xg3mXrLt5BSMvVb4zRSxKDq
XpqhPrcGEcGaeIoiWlYmvc6Wex2M+nzp/sW6llqAfgAC9AAW6UIJjd/v+m6NKkkW
OqkMF9f36/rEWLq0BMps4ewK0Au7qcoDgp5MshTXXm8UQB8LN333thLzi+XqBH6x
Rg0hwDSoAGsSs+oQGG0EubaKRXoCA4MRn6sFJgCWzorri14THU0LL8VrhxmetqAI
FjbLYBsWxw8mx+oBee/avj1dfrt7ceLaccXVE/tzZ8l8KymAbZvwr3xv8rNfAPml
obgnfXvleO8My7LG4uek0LRdccSxLefsdM4IVi5WZymRfld2+FJrI4PwLJHySZAZ
4udd42Mfdr9TdiJ7UJvrKxd5Pzid4hxQ8/fSETJ2MXUILhAwZsjxkuULMYQ/3Fzh
qkho/Kjt8+3brdtyvFGbLOWDKejpzfF6r13hl8miBJAj0c7lMvxYkYrLV0SKX1d0
WbbORVSZ0wriIUA/luFv9lOlLvQ4PfOl9ttg1hRrEucnL7zZ9qEUuIvDqb1fHu/e
/pL+q4Ld1TDKWQA65EDW1Tv5M07xDRMUyktsvj3djs+BjeRmKVupyHUTKdBlaAW3
5eyjPOYCDqCmKpBEV8qDmvFgVGVNfuEX54pd2Yk2cFUJYSAlv474cICEp+NXAJNS
fDd8tNit41kJhxB70SJNSsjIulMGT8aOEEM4hj1QUzAySRkYW3hCSmdKRNml2ww/
sli26qfHHsJr+BLHTV3krF8vfQ+jNZY488tRdA7WyfanXQCzX12CFIduPCy/1kym
8aoP++rB4LFvitwMeZAs4FmSBHHQ+OtJOiT2r57CQdD5UJUCpqXQIWgvdWA7syy3
QvQgIsGrLxF7+AR4H8Qx6Q1LC2yu4h2yLWrSoZXT3nqVBfcxmue6LyKx/cLeKBx0
a5+z9+NfiVnWvmaqJLBzEkDA4UCzn6LJSuArqmZH+l9oSTMOTwzPkHsl0iczaK0p
6zE4vgzDoXXdFi6iiHBVP4lQ+i8mVohZa0MG5rcLz2FH20xhPyJxoLeCadRLn+Op
IDUQ+82rSOhLk8Wa7R1tMgt4qhzBk74BiP7vVZzsQEcs5G90uzKch8wFSAYrGYvm
SkupE34cWLariSFaL473uL1O4Ikw1/fxC+lXRNSTIc1UZ49qdjuH3YRqLdeR7hdB
V6z8rg3wxJ3V/oPjth0LfCplt+hZjLfBiL4pFHQRsXt32FjetRTVdTr5oaKyxFQ+
sQ6Uqj8UOr6ZB0dEYT7qaAR0eCERVOweeZQ6aaa1S4oasQQjycW50acLCiejqEDW
ri3xCSrMwxTtuadYbQHkae5Y1Wwk39xNrAWDuV50xs8IzbiafWCfDC/Lq2uNr/hW
lmxmyVxaLiEEKYdHFa9J1ob4j471hooLbuGYXMO6gL9Oenm3+eC7LZ1/yXxgZn4U
r1KuPJWorAmNIonW/coWtKve1YWYkXx7ZmRw1w7RovjkblLVBJUsmEyMbmzpcDbp
eOb9mmC2hw2whCg4b5d+UMc2Z8XgZruchsc0kskS5PYcjCRZ64q0krW8JjJG1KEI
Nj7ODEaP3CakkMvG2FuMTdi/P0OmYOVkbksyxqbHabByGo5Aa5nLyJzJ5B/+wjlG
KK5QzACjkRyhQPyIq8HaOQk06Q+zWr1teb76kIMigOJDfTx9dt6haxRWAAQ22gH7
gGQd26sRluxSSa9TP/O3cZhveIDODz4Wm8jSGEVBqkJzA5l/2+cOk7vtwR2UWs0j
QzRsL/SdQNI+g87NSYQfhwSOBLunhzAFQCy19SShII2sUF9lyS9Nsv9gW/N0Ar/T
C2kacbHMbfxcJPIjNqOqm1uSqnBvCyo3E5/aFCIMI5+hI+SULKb5+JRFvKMfAlEY
a5NfDkVFcyd8qu3KW2ae3k9dGSe7f+2shSG15GnHlVuYc/U8fZXMJ68E/tXeB5/P
eEK+s4Ft3VxshRHUuHl7wfqhX8HJb0OlBe+HrxZWBHevBFx6chNavBzb3J5cm5pe
z7i8fJ7gNfxH+TiOXa2AAacUcY8PIzuABuvRfNXc0m8vl69aCXjZvUxqu0Ff+utw
f6QVA+EZZAkO6VC0OekrguHRLHO2Bnxpv0Nypu158Q+0AKchuImYJMG7qnRbAMpf
2PAs9Mr/ckpqYAiy5dOXjufsrVrOCxcCPpDmLFtsHRSYC38CNWXUc+v7GBJGSVPk
n0aPxSZjJChOTHCwtgSMin7WuqIgRZKes/NfbIUiqPwL30hdZk5sCarz9z0JMlI+
PxHJN+BJgmuANvRwsy9soA+nUn4fMldMUectGxX66HU9W804jsW7boRBuriEqvlP
0zMQkl41FBbCqHRmZMJ8OM/AcT5Yps4QJ5QRW4PiJN/+hHCLN9S9Ouepb3Z+BkqP
Mh/dMfn/3GJCk2kyESgU33e6vie1HMokWlbO8htiN1ubk8ZTZBFtTboY5ALsvlfN
SpQ6YE0AnLcPzc1kO86FyrZUUZVAb4xaMmNioSayda2nr2Fh9PgnQHlorBPsk2r0
Ae1tBBEqgisarWXF9Ooyk6r5PxnymcTlkCdCRcGyKRuUpyHYq0bbWF/pFtHyegnP
Yd92mqJXLNJ2rPWyQVFLHBOml9Qr6vtPmigEyh6UtoJ2xj0G9WwCfDBwF1o8c4yN
QkEwKzEQXPaKHu6idYTDvMU3UHZFmPJ11CIqU7h1OpChoGc39I8h1w+rpLZjtz62
QqhgA6oo919QdkHGgRUghJ+iMpvwmCZYcsde+Pgry4m2iGwbc70LnbWfPkq3ON9b
sCIzSVLeFmBcnzSCdr3ShiHVu75V34+YS0poPR9MjkaXWiAxmAwFQZhn0WfyL9Jj
KboBlyt1du4NpVDI9lFCSViqDubbAyjs/hmsSrR7R/3q77xLSu89FIoxQZ/WgS9b
QlDs2cJAw8XteCO/u6omMdhQ2lDrA8uneD47jA3KMR5OiOVaDwF+PBNvO89GlKxs
UwHrXFvX/sUsbdmFtxubySndWQhTN6z9eFQafrh8QNYllibevyh4EFWjPCxmQKyZ
o3rp+08Dq1thmIdmMySRGq3ycc2svKQtTo+HIE2Wl1LOksJd/E5HLG7GxNbk2eP5
NlpVigl0l4Zcn//wZtjIZ7ir1Pvo1LswOvqDujb9abndI/MhaCH4orcFl8o4ko8K
BH7FZbGmw1KTpzwJthtfab2E1UnRp94V66jUxERgoOCY9ZpoPArmzMKvx2uU2+UI
76L13g6jh21CG8FDwvT5qPEBUBJ/AJviH/UbCDj63Qk1Vlcbg5mCd1BBFswvll35
3yS7/SH9dA4vQab/JxNg/kYH/Rv5pDlklg2la3dhPSXXoaD9mBT/Cfu6SOdRKOpn
LDfw2yl8qliBJJ2t+Dq9H+guxZ3j8wp7zkfoTdAMlTo9bUITj9/03AYIzhODyNiJ
82mEGaiG4JNFCiyxNlWC//5aRjyoly/kz2V18XwuZ+Kv+1k9bITRM6gpeyuF/+/b
QyXX9v3N6JzRZw8Tbb2WKHVyF4gIVQm4FdYU1baJrUhbn7Dh05DIus+ltK31bu7l
LktpRD7uwDCTSV8S/EE3meDB+S9hV45Wa/eICx9Z/tFQa8KgB6tnIcLMxOqCEgXs
3eGuHuwkQ9jknkcdoU/8aUQShV7rwPLnldZ6Bp00/MpgXJ8n5PZO3CX7uC52k/5q
YSSJvr/bOzQYMy3pzvoklXFG05nwR4u1z+5y9WqPvnihL8/RObh/+b/aARPs0Zrs
nHeCNTGNynkyuX9nFPdH7XnnvkTw6Rg6f87ArFtHGLti5FvhEKBQI2TfUDRSjOeO
1MZnClrDDEX3N2hLlgjx29tybGwN6eBVObl9LkZRxdHtQGTmEd5ncXTiSAkHbQNS
cUXZi+Exc4fWQ7SqI0Ac5H2tvv3P0s4FEwIH/7c4tllZmmwqy7vcdVCRdFqFdymM
cbdAB5tYWI9gfAwnbKbU1pLDoP7Ryt6lcWB4k1lvv8KGj82Op1XwK2dON4/XqPWT
daVnfzfqGLLNQDyaDIyl/P8Ls/Otliww+IRxLkmqza+M751R7wkaTyLDqa9F1dBw
PtEGvQkDi2UYucTq9S5WOwKdvoxP1Orw1e/S2IsxcfiaYxx36FUs8tf4mr1wr2IC
fbuJpTjiQ/RbJjJ47cq9+adHYTmDlgkRSfVG+uFA5fz6AxhZVxSKgV0mgd4DtD60
ZTc36G+prPt64+E+yfbVYTBGjHCy6QWm44g97eIsuU6TFPN0NL3bvhiJoHw4l0xj
ZJtetn461OZpVolyrw5TLAJpvfuB8pobw77EZt5p2QBHijIA6CbAT7JNsXItaW8h
qTndTuE8enp1j/4MNXO82ANzO5fXRwuBLeC4MtqJlO6tCQb6qMNvytRZ9Lnfndny
KBs9cJMKf077CStX0SSqLwnuf12n1GN0e97tjXcSh6xKt3bzjQ6EylyGF0L3dhG1
ObPkwnuUcni/A2Aw1WJ/zHRQhmpFBI9bGhpmUlNgn1LHkcHZLFvtmUXd3tpx66kz
Wq1TzNU3Cfn80EbogFtC80UaAFbFp9GfYEuvtV4KBQCuFuJrWiY0gKCEh+lbyywz
Sg16/XNyoqthThVtwG+vHGy+mjfIsXOkhdwWtnz4/jZJA/rpxVcSV1L2CfKHlIrl
7mkSrkvl9cLCKXuko91x9IVpGAlOfBaPJNssxWtnfP2AK3lOwSyNAopwrDU6DE4p
OZIkbDz+0yNUcau7QX7lK9csCYksHb9buLl5UeDmziFB7n//lAZioEQRcYl/OXXZ
z7/XbTKIzzZrruy75WPAPPvHXZPc3y8XZGofiOkHsSqdVQl7B4Aanlo1Tt2XlqmS
moBX3225sZxCLvfsx7I72pCK73b6HvGENMipEdBR19DLHWfs52+bfAJ6rKHCDBzi
HZpmdau/3lGApIBASQdu8YQz7D+luQH89kkxun6cY/4a9WUKPjol6MERm0cgQwxl
1lpsg7uUAIek/7I2kFYwun3p/p2DPJrbnBCp5xY6HE+eqs2quIroEyH1i5TKN7nk
HtLDDEfvNWDQDoB+etm9pPqLdqM0/9/PxXieDCAmmA2nZirRwaLTO2Ob3t/ZGJHE
LPVFlVclXxXmDVsovr+lsAOoo+4kh83ektgFjnnhF7yTyDH56N1k9/gh1LW/Ys8X
vtQ2saDVHUeUe1MPBJUBQcmSEovrMHyUB59BgJ542aiFVwyRWD/TjfEnv26OnmsW
vni4uxALWPufVHL1LOonzApamck3gVrWRJt6EjL9WuVja19cF21uoriQxwHHpn23
BHr8H4UzHGHsMC9UIosA2amQh29fUPs3TfTSFrnTJKjU4SmVNdvo/79k9Q+qxrJr
0FqOkbvOxn2CaB3DPAAd8VFb4Go4xEFc2Yp6dhifdpdoeYZLFyQbzFXAHced0lto
7yrKKeqK1L+W9zfHTgyqfUv0SqoTlDOThtmdR60czWjHOJOpbBL+MvjRKYtVCPoz
B14CVtwp0D+AKeODjUA0fS1F3ewIeeg3ri0eYXloybsVH08CfewXouy15ghI3ltI
jPy/dzBI2MF3NK4FuLbr1nTiPIbG0A16nluEN30cwcZOY2wuWKQcZpXP6Zn6lAl0
H4FGhuHWbXxzy3E87FJq1cQQQyFahJgtetyNBC8KWsz+4GcaTu9PFQTLVc22pJ0J
KO2NizMpDgw1PGhujYjCBr3Dx097ZnRiisyP+AZPfXaobHxyOTQ9JT6CnUi3OP5V
lpC/2e4o296+UFpucjp7qjSwA0TVmfJFWS1u0NdBZuYRK7rFGjqOY5OxRqRe7YWD
53MaRHiMX4N5lRLm15X/ySkaC2PDQlB/rdlRo7YSb8kSG07mtYy7qucDl9ESGcaL
evJCuZEnWiFKdadqmxEfSsBdSlLDCpUllbClt8yPLjf7Z5WH0s9YMo5NaqnQSE8b
CLABdQGwCmpib863hHoSVGhnnrGKDbLDjH1kYOX6pDlrz/3uwOURkMY2MLcxPRDG
9BYGLejLgwaCPVJfYFIt8tyUxQ6XOonN+I1uEDioqpRfk5HVmmOK5pMoWLc/6Wux
dVkmI5IGVHzy1kDkyBLub468Gxl+iMkdj3Eq8/YRx4W3AtmrBv8Ia911xuAjxulq
ZuorQodBEs2DNMmo5QLQJwfznaC5X/HHNMdppBTN3s6DhIJgOkmYg8t1ATpdi8wW
+zt0nlsq554HalyHC970Qqzh1ySEdckq9d85G2qTdeO5NmvQ5CwpCj3aeurA8ewD
fNkuUZaOn58qGDxsl0h/UXCDoPbVTw0qR0ZvKt4mK9TFYtnGjAVWHDfU7OrxP4o3
OIh/lJBHEpEHU9crqgAeN/Jhr4V5auU6r5BSyu5R0HGqTvDHtoCKFPf1I/s6oHL3
BXyJFdZ8lKrywTHH28xSZzvLB4y5cP1qnh0DbOHxEf6oeHs/OzfYMCFo/jI00rWg
teepKvZBZeqbp4vntbHe02g1FpSE4vZOPy0OPybo0+M+XdHw5LqwmFHqN0sc/if7
nJLTdwHw1rUuISZA3zIWBULyQXx+Tebsr3aiTe4uyc8grrS7xvK0FZrtJuGrD9Jv
cuGaQi/tGvcV98EFbX9my7iUoCUlp16TW59Uv9os1P/JlFYUONMaL1T/JyMYnqoS
ngoWXloXYWCEUWxv3e9ztmGBO+Ms2Z2ClqrB/6vSqwi/f1qAQHejkqIGFsbnvumT
UWD+7Nbe+Ax7qSAb4M1pa+K+yK3IR41N8fRtmRY64kkhQSXdjeDYDFLvnnnW+mY3
LmnKhjdsDQVwympwTqvdUSVKPHZWdcyGbk8D28W3LUGHkt68Ms9HXdEEiGAJHI8i
KVMid5/BMTtjjilHUkjWJswV+n4TmQwX4Rtb5C4DJpY7z237TeuG+C+y0M9L+zs7
1kD/Cm1rSo3l34dRkTo4x8DYEHQvy9NnHk/9JIlbMgwUkOOcTCnMGDd8WQsEseQa
jiBTIFaxf2KoDjK/Pkz8ZosXITBbIRkduASOftP+3/VSAAPx9qZZ6ES7W39INuXY
M9hY7uNsrZYyhhX5h09pDAVK2UjiDPYP7RK15pMURLrNZKAU2siwwYpQH8cvG/gw
13ZOJCB7riZnJI21HmZWll4WrJS18xQxnnQlJ5q9tCwUDRwrz18+1WJ8pOHBzP7N
ABKwG0KiNxfJdjaYE4vBFgOSN7sBYuf0LKxUi472PmwnUOhqtjg/IssjJXIlTQIk
GIo7G6wuN4Ze3JvKN7eG7A+paWfQqXd9jZ+At6tUK84uHBzV1J7VCCycP/1ZCIRb
/Nn1QI9YSsd0PWGFRjn4e/LBN/MzO4/hcMwX6U0dpwCajOtkgH39WMXx9tE66eI5
KMYrCkMWp9hwvgQRAV8uxkhGEI7STSH+55kDy2Hb2dv5mIiw4LNgozDnI4Pu+4gt
scj+iSVGZMvlKtCTyWc/CX9EH4LZy52VLGS3A7yzCmeDPOnAxwHB0j33hfLoIP9n
eoOq5FYEZ5YSKMW/z2weTlINk2m8X+m0FR8KdnI3Cy7pFqkEojiPyFYtdg2y10kR
Vt4QvV3i6zxOkhaFWpZQyWH27PrOu+5Qq/34qkNW3Z3nbMs7u5cczouyrHToLx5x
jIdqLY++CcGzRhhzb/hwiOJPNFg0ul/a9hSLF5en6wS5T6pElr0Ii4hXUA+edldB
h2D6AvDNCrGOhJ4DCFA2702iEI7cvBvRR9EQBCxJ3PgIFBQgjBj0iCm7YgB/XKTO
c7ZylVPSqEM6xyqyeLrBIL2OA0mVD4a0YiAXsz1SHcz0DIy2v94HzM/uYPqePxJu
HHKc6GVCGnPA+1ZB33ry+9MzwfeCuehFPQNjqPJUJ2rBp9s4DAoSfJOGLA0yMe80
qcgB9Zqx3v8/aBPhSOYzIgtohSyHIvdsStGbA+PFOGQgQNDR1crN5jRBtdDK5xSI
f5sh6GFlReW/k2UnuJrJiWMXx2avdit+KPTyStnM8M/RAXcwBngtgu4TkSvvbDfF
+qvSl4N7/+V52xnW/jPtaXhlp8P5gjMIMnYzIX5BejdC2AOtTQDy/szBYJ84X2gj
HaAy2czKHZGtScszO+1cEm9Z4P8FkoQhTbXCxSY29KMZmC6wlzt6QWhQwAryQk0z
v1GKvbM6lrq8A2HDBSewl1mD4u9fD6Io9kAQqPCKT/DIoS/4AjIa/2V8RnfH/eaX
QmYKnctU5VmPs1tl8LYMo6q0yvbdlJ/4C5jp/frwtEEBom5YZly7fSQ/CuM5tgG2
w10f20ji2BgitMqFs0OoxmQlW5yUQNGAV8uwfiLIHkQf+zsJ72Q6MTF00DohOItj
JqfvaI63+WX+BlwVFyyRmWslFWPpRZbVeUU7zmxWzSGxnvhuwLPyKqcKDCBfpXJ5
L1LJ2K3L7t7xQ4JIXF9fzF8yg7W5OxTY2v72VPdUZFECWYH0r7jVQ1sgg01MSNHj
TxA7V2AheDlv6GrCNi9uY0dQKQ18HwauLXC2mxx9gRFjmbfbcZbnYRw7DsNOIfB8
bHKFkhFoXaN748m0Nq0a4oYjtnyWfPTPLIf+DctbhgOO86MAvIQmWqNybs4JSr32
f9stQxX5GCdYZdgw4OIuxwL75JT1jDK1+wcEJmUG1toxi//Y6Jk7gCGYBxUal5cQ
L9Zz6mQ4r6uBw9dANnRBKgKPXHdUUqP3n9LfEBubU61c/ueO9ZoI86jPYAw1hc89
6cMYNUI7L4vBWC2t2oMzbJ3uezkalKM9+XrwTE2UdTvW0Xdq8pJCS63B2c2ew7XC
lTANtK4EtXM6cRS72xAUtq7D8QdNqtmh3BMnNaHHFJhVmwBhd4kbGbvYCUdgjtyA
cDTd0uECmp2ORojMU/+oaNbAif41TY6OkVBUkGQE3tPY3h2svPVVG9mw1rsmtxXc
9tpbkMtloyOtz83Qaf5QwCooBKRaz4QEzXag4vY8OESM/R9okSI7nEXAuh8eTVYX
bzHs41h+TGpYIOzFKTPImETU4GkbwjS3pF+U8F4oVbpUnpe7sYo9VpmULkZ92dDh
tK4TC1fT0g5h34JoQYLFvgI0p6YIrcy1NJMW6N2pwkZyzCDdtg+uzcpgInabaEq0
oBc70f8zU3o6aXqFXxkaPd30Gp2f4bTyk12LNokn0QQmGCweVnV1/8mnwkqgirR4
x+bsXiWX6s/ONecjAXOrhjMJopIDT5s6ipLQEqk4LROhxDK7jRC1ZrmTrC/wtDK/
7fafYXO1GW/RqenkC7/BAa3YRkLK5CHW8GFlvHcUoQE0tP2merxrVPvuhyLmhr+M
GTTHEXYMFIQSWSokTPNCYKHvrlnrtoFF7OkdtJN1ONJlVotdskxRt1NFpWwZ8PGP
HJskY3uIe+rtpFJdiFPBqf/sQ7KwHFeKxFBGUeNkY7Dy9+3uGfclGmqi0Gt/eDDD
LKWfWXeDxEqxvyh5GoUzLzbnE1EmKcrO0WO+6jQJVaSFUw14siSLen9AA+EUxfsN
uy0SL2tFisyn04mhJu54drJ71CYuXL1wjse+xs1/UgQ5nwJA/7UF+HoyrW/Oq/SG
Q3b4N//B447J/4jXNDoWU67GblvzqG625pD/pv5OPfJqAJzqyvWLcZKchElRht6C
iIFyMyyPahfF9PGJbXgK+/feKRdfQMeBXODTf0m4o7sqmcagxUXlBe13qtMtDXkp
zGchcbc4iSxnq5ahf+yY8m9i36+H7/51X6Uz4bkFPPf0wk3OdnHWaODOC/JQoOJe
e24dxXEENTBA+ZBHEoaW31XpwYvuYxUz86OeNT7g4G7OTkj4xhb8Vf/rKyVMiVf2
yi2LW6EasJwmk74y9ZHXfgb9mxIRepNcJFJKTkY1HO77uoYDDufUIm/Ooyi0p1cF
sPGCC+i7eLu6e9f1uu7q0rQSHNNuzWKVYcGv5cu7UZ/M6H8SFz5EZjEe1WdYi9rT
g1qeEp+94WRnIX4+kjJqjmHh+26stbScYJFgZaZeJO6svNCs/RDaM7hbM6UUpGRE
IDlB2BYgylo0x9wcl2/tDnj5lxfc3W7gAJ3cc2yx6T+AdmyEKOBezzYJ1dDBIb7F
QsXJWxUh5veEmgZfKrYFjCq7peT5bqhySht32xQ80lQOJDTB3Q6mWLw8kV9MWOpU
C2tA8Ct33qC9+Dv7FLXsuBAKcd+OuuNNhJRckR8m73spgEbtjCve0p77U4++olJe
Ev6+r0sc8INELjLhJVu737XYM0UVXBdsPC2KBwS8t+rG/Jidfyryhx1LgldhINqD
amRD92KEyHh/8mPBPBDZObSzKC+A+3ctV35p2Qm44qL65imdn6/c77tE7F6HXyfA
gTLHepDGfcKAieOvCNrxZtkqNf5J+5mwJp2T9Eb+QsXQCYNykbvlcr4JXReq7MSh
xqF0nytiOX3OPL/B6YSGhn8bj4k9yCHHrHpNIN8Wzkz8a3F+ktg2oJFOqOWM2HKt
T5LY2ejjceqNFEfQV3YoVGApotPmN9KLAygp9qj1q6PUtq1D+1TljwDA06p+meG9
8m771sgjJHON2JS5S3mQw/o88zqxwXWfcVY8iFEwoV5cqqv93ZEcYrkYvRZ0xATg
8f67duCGKec3EYS42IeX45dGHPBuaKVAgsDdDm2hsWhkj6dPbwsuCBWDDUAbdoL0
eR6AtUVMjxZE025kF9BBjrCbGXierUi+cVnLvV4Gq9LHpSlzcMpTHm1JlHfLbkGc
eunioNX/o7ZUdV6VTuckoDPJMXXzU/ELGdFK2UoWn9a/yl9rb4lQLEudaSAj6dy/
yA8OWjcC9dWs0pDaxHvKNfgJzPrXV+2ci7j/cJaK/f3+cJoBDtHZ0UOIuscPP5Iz
YMeL8nFv3/lFsxmUSPbYJMU4pXRkeSr8ev5azDBIB7E0b76vj/ZkWzdAQ5hz2xNy
hX0bNRjlto09Kp7YVXraezpzCF4zZQxGopb3b5bXjsC9hRv1MDbYe3hsPNcr/D34
9MbA496j+RHYu3UH09UwZJuTuodV0P8hnkKw20KHVstSx3tMyD6bvlAqQtbxX7Ya
x6CnT29pA6+3mWZejygQSBPHY98fGkgCCxub+pwDKLHqN9VVI8bKclIPuRvw6ywx
CsJOaYyC/MYOuqPa7l9XTAgW31rCJHdzkEr/O3YNFUR5ZYovCZuqRgP1u7WqJHRV
rN1h9cfqJi2BDuIV67Cd0diRhKr3jSqRMyJK00c2rUUda7HwmvY9yqcelhx/EpnM
MR0DS3dQvx5yn3iZY7lebI+hnTDfdqbdX5q3+wVhcuTwVUBYg48ctBjt4tF92yPx
zz6ZrgXvyalK8d0VSvbqpKZ7RwY/oUKuapP8fh0OkvLMvk7Wxf/FBZ2mxUwwbg72
NCsyUtEIdRZ9/vfhSRZuebJZHg3gRuKcWLSyMRfqSTmyIM79XCOiF6iQvF5HY8kX
mUPkiJW407kjIjiqDyrdjO440db1xAOw9NJyRrCD1KEO18dLrHAZgTVwhXubQoby
FPD1+MohkVdp74lXx6lItHurMNMtSxaakZzzrL5pcz+TZOabu/6emBKc6au4yhe1
JHYiGdSq6RWQqNdyXn68u/ycAEKMAlu+4wkCrsErhD/MCFLW4eIYz131DnyY/olx
3GVmn0Tjrp3Uit82GflG255x2SZstFKlkyT7T0Dbw5X7Ewq3nldCs448VZxoZQSn
CWaFJpBnfnqU185RRNMYfh3zOWSp8G9h3lGy/jYr+XKHCO9VNCqjsRH1fT5vu8Cr
OH9p36UuqM5KWGt4pm9dPhPKnrVrFUsQ85dB6eA/Kg1u5/QrYjUuvbLT8kUmFfMC
1C2RiFFDhCbHkr/Qq+iiS0c/o9twN4qejExV49NjtBf7mTusJJZLWztv5XG6m/36
o0IjPH8fYEI4FueVSxyn5rP9fXyw78kyUzsesny0AlFfOL9abqlLr9CtIkDnCI6w
p3OkGKdULxGaLtOAPKa540ID3KHOA5Ww/VxeD5WwteoQDNCXOGGz2hXg7Ntjq19G
rv60JHc6R3dzr1jlXInHqeAmNdvrq2BvdHMNZ4SRdRh9Ioy6SgcrSMkbUS6yqZJE
/JP7EqUUZJSbw7qgQZsdsnMs8S9sojrRpuGHi1rG7DHOQlGl9w8T9N8N6ctGZnC/
fVUGiMFXrG3GwvVg3eh1LQB1sjuech5Mwl1/MNBT6MOqFl2GBCklhdaADGiY2mQl
bDj8HpFtRr+1TO+70Rb6NHM/LfZBfVj6mYiZv6ZPPKKRCKqU6L4mIJB643aLNC7z
vpmnLm83atKh+Bjga3ZTzdWuPUyD3XqdW2aLETkK7pQuTglGxMeBT62Dpu0M/kdN
Ojmx9iJ0Mvd/ylFpmSRuhVeQcI2tsWypH5/74n104Vu1Lbl/PtTUQtvBznlQEB4d
E05bWohSpVuzna2+03NKVJlCMoOV3EzYi20j0BYRWf0yvKgs3+XZDZK2mhxA/phT
R+wlKfg7b8k1117vmeHgFDaNez1GIYuLyuEXDbkbYfD3s+oPVrR7YkN4ILYtC87d
ShQft6QRyJ8vwnAQUHEBl7ZyLu2Lm0yO41G1pQYd5niR0wavZxckgbsdAQ9Bku78
2ayIpJXyfb8v1JVAOfTI6xCMvDJrlA2/xEdOF3DqTFs9e4eJidZILWZbJel4wZd5
2GzrOSSKua1jLetuVndbjXteAp25Vp4eUI3BQuELfD6h2Xe/AIpWaL7UDnmGFsfp
y0HJucpvxNHj0xm1IssffmzfpkLX3veFMReNTN2IxeSqi0umAqik25z4xylBvtqP
l7ZU7pTEFsLlRn33m5kxg64uvPR0g2wmCS2yufABgfHVmhwTF4G3FGFuCBH9HeQF
iFW+8lHIooQY3lEx2E1+vEUKmdtQLXCHAY8yybjaoPVT7ov+tSjLsPulfA7+TGMc
gg5YBbK0Vczo72o/P0Nu+hO7wgO8xhQOqmmrWNGkmZeXW7iV6irAvMqzjZ2U3Jnj
mIUawLqw6gD38ss4dQqpn48UwyWi6KM9Rbz2KOnBx9CfkAxZL63el6ECUYZnfVk4
DWiPyQ8RxD1+qM/O7px/g7LiU3JbhQcLcwbuc8aSqiCgVy+kiw8Tkk0CQsLx/jNA
P3pum/nfFa2m3ZTjUDrmNqWsAD+DQ5A1TRmqsd4S0lf+Vit29+CukaojfFUU+5ym
z0Tb3x5v5fdybQvv3VjvcWZ+W8wC2m+JM+jenpbSmF9kBcuzdN0Mi+ufRlf5Zqrw
Ei6kszgLyEG2gV3Ey1nIo9b1iJZ5w+LjWOoVR9KZLacVnD3r5Omb9OU6CDlr2L+r
UKC2XsDljY54bgjvRScYv/k+GXD7oGSpFJv5gwWSFyJQxvUFUkmQc7LhV4xpnvor
PNvjZJVBrW0Fh+XWStX9r+2QLuNzn8e8yBopURPUOoHWgnXybFM6EaKFrMKX7bW7
jTp/EWnWBy4HlkHBk0GkGg6EYyVFYctx6XEWfYBNGYI7y7F1fTAhFNVc3pW//Jt0
zTi2h4rhOKbB5Sw2I0CIV7iuf/E1hkaIEWZOmUe6Vme7K2aAv0CZnD/FmLiL5VXI
EbwspiuS1OsqgH7eG0HM+PbAo1zgDlh7ngvhHN0+i3mHeMXuP58Ewwb8UeRRzsiX
zMNH0p2Wvn9FF7tJhf6PHarICyY+lbNw5KGa8mkbDxNIi+yPSZydQN1G4jX8oQXQ
znTRcFEUsGVez72VepMMcrHko+vCuroKMeNWYwhUzPRO3ldUpdQEyAB+adkTP6Xq
xH2PhB4qd+a7n4OzaAyjPy0LPJaf9TFCnV3IXZlx/t9dzoA8n+9TsTqATkYOsrNv
4cWhHl/oFr1J78+yH+nSv97TAMtTKpEndHqNMU4omvMX3Pra+XietmqC5JhuTXVo
AxLyS1FqgO44ZHLSau9u0+1s350uDEivZ5vDPayKYh7GUhuZaWgQwu70nDuDnkLa
gFVemrAhapEU2SUyJ2NfZCsemNgHjAJfmxe/nddSABHt1GO+E7jXqv07Q7cSAntU
wRPyMq4RE7oHSpMtB/0Ua/7c9AgTYH/TcHKjDrP0O8NUqq5QMNEetNd6Do5+3qdd
hOLyweOpt5zBVnA2FDrsqJ6XRjMHAD5gO3seLMThC6yiB8WZ8eilTjB4FEu8Anew
FHm0fOXgEXuWnGRvbZFM1BANZ9xVcF+jGXZb+9dXCgE1Ta8kXiEzFH9bnTGRGQuv
vZz783BtL5688/454sLYLoqOsDzrCkZKjcCJ1xcLojW9h95IdhTlqtmR+prOkg5r
Mdnps9Dw/ZmrWrw4jHNhewTWj9xyto+g/GfcMoIBSRe7nXQ19OpqWtTPleldKwkq
4jPw7uvLdXjjbYIFMtngj1d4UVSM+vHJx/o6hjkPcSb9i+dMeH6+TNhNqE4pkfR9
kQKEwxwG6Mi9MH5WsWJ2GO351/b1CDDTneK0JQTBvdwnfwP49yJu3zPyM5wB7gi6
ti247cTmT010AFV61OMubRQ0TIdUFfpdG0EY/yOY8kjEl83agp1Hfs44OLQPxBeX
t10g3taTmaSZeuMGxAmO19uzv5nvAa5DTDJ8Yyjt/a7tuU8Nynqr1pUbnq1AuBlh
pTv90J2ZhGNRh4v/okJf4A9bqIHqUoM3B37ZbW4eHU4blHDj3BUnn0riFWokX1RD
s1s6BPFHBu3fbtBFGfgZZWngqC8FLQSIyKQOb7tI8GP6S8Ona68d4HVrdvzipcIT
6OocDSA0dPDc6iiJGIDcV+aotnhy4QOrXgClpB8gHL7M8rJPgEC89gaEmLTABAuI
DvMI/wdKNbfuwN1oGYz2cVew5q0N7eshdzHEAtUQAKxsR+D6B5odr2vjrbRnkggW
/kSx9Aw7RkaAUi+N91Gu01VklPOsTeR1AzHnenvdtPTsm2u9fc0ex/CCpkpQ8tWK
Lq81R43MqA2Tdr5fCUL5F3YU1j1Yhop74QgprqruAzq1U5biXHW26r0YMGklMeGO
+f5zJiOSiXPeOxwxBCvrUKcNHISiTGI0g8cfcYxruU5hA+ktqaR9pOhtq5+HqLzV
qcXDhUY7YTXYR6tJ2LLAsM0TRyb/C1Xu9qh9yf7Trs6Y7I26ouPH/q4zZ/LtHBqY
yY+VkKm8fWcwGLeixALH5z/qWXc2u3yxyUsy7m1lDfNpsPDRomiIs0vK851Itxpo
C8dMLyUx3HsdtYVgw5z375QlGZyRbUIX24HO7rMyvvcejY7dSR0boY72lB+gMckT
IUsd3S7jg8MnyC9SNNqXp3rojjG42C0IIn/p+GabReqA7zT3Ew8mHae7BFXGWgOJ
gRTCItP8tjebk1a/KkKmLPcSyQ2KZH51Cc368KWxNKNayXCvMeTddcURLjSXSsah
L5sBvKmg9BltqW+VxW3I6dX5N3irUSpAtfvannfm611caoA9FkYLRbtfwBJYVOIU
jsk34qV6FtuPnGG753SU8iapEOta7i7lXRg/rgYbyEhWrdsGdnCbIDmTDAlGv2tj
ml1NxsvnP419cD7bywIX9kHD1Gql2/nAeASDzMoEcKP2ZZSGSNU+XbvwT/l13ddJ
RuVDRCYYIJUOASGuUfzklM13I4wjkRngGRRSGyM3MtW6yOP/QBxom2OQHwsG4jPD
N70wEhtwBUQyyq9WYfo9vk3iZbfdHZbs2O+L6kEe8KSermN/WAwzGbIFpsc6YGKJ
ijnrpJroaEBkh+KimAw+mZrTzR6rm2DCK1N6Tl7nKN65ncmZGI72nMDo07vzTPAG
CvAHLyWPw2k5G3T+eB4qLwC0wRNE47+LW/MrUBQOIJ6ffX3xuu+qbFHAsDHeikQb
J5nSie1zu7lByrMvlaBWEfom9QKZB9CwSANiNULSQ7qXP5DmO+xyMbfXSrx4P20N
j55mLqoGjmpKLza4tkvDXz7WHYf5ct8XiXCu/hXC/nj9p2eS/hhfaR8fmU/O7Yp6
LQkF3cZy+s+nL4LzV9y/HI+qOKQ6+3twFHTvQfWBW9uXSHUGrnhtpKqo6tQiAp38
KTif0wUSBwPSNskqrt2N85rdtclGqJwW63micMY6Fboo0H2oJPlsOHh1J4T1pQud
IHE+rjEsQzqgVRVJhmZ3Z4ABQkD8FyVZNE81uuD/h/oAxV49ZFDmO/+wxgpW8cFh
wve5H6zo5rtCm31Hoh7Onoal+afYb84TrFpj1PthZVzygrf3P5w3GJ6aOFeOn471
iIIal+lXb+BpA1I8rmuvnlLV6aADThuBZOXMxKFEE9oFry6Jpm2yfX5vqTPdYCxv
u0tIRX16L/GAy1qOf9oUiKN4gzSkJEdkzeTKUvkIxc+JNjVeGyzOOwXVo332ZizJ
iM2m2ijuxFIYoquJUVHzVtMV8IAKDIcax0enj/tson3Dvw/gtB1ZE4ixL564LVFA
CQJy7Dj8DfzAxqEDCvYzpLCh1YMCXvFhJiiHdbLusVu4c4+TOeYS5vasxtKSSaiU
2bserE9hs2EVD19grw8UA7pd88l0MjWIZSEL29NO7nolx9HS+xO0lZWTPEiF17f9
oV3EQqWU3noYVDduEAnhUt9M4SRQyoRT9JSrySNW1OGLDgyZ0jIYVQ/eaDZSuyax
FXVgB+fa+S+N6oQLxPh4ecfx2bl6dcIQ5FYQf0qIra+tCVbVMmUTE9hcB5Igm6t4
KkgXWBLp8GH2Xq/qFtWdo8XU6XPiPSE4SwvRjBuxo3Zmj1woVnZXxOdZ4mF6Q0UU
Er/dGMjjfSbXy7Q97HMyB8j9kOUChjA7vV/Kjl/oytXpSVkSv27H7g1SiraM7HLr
dH9g+OWWDFAJf2ipU0yMhXnKX/9NtgcA4gWfH7ib/59Cuh7lGQlf0GNLy+omLho6
AqLg9YVUKUUsO+xbwJRLsR0rNKSki40Z9aEMFdYIwDpT/tB/cbanLZBQ2vs5TYks
9Zx8vmTSOtC/fwTj6uddF4P935wQxCQpqGpzEJi9Ekf/LcFV2wtM5/fTYiPz8d6Q
bh1kr+3FYLz7A41yMM3FvvfjBG6FJxkOWtxck0iuSGz/XEzhtYHvnb8kvycBTWaJ
uzvRZFgnfocfBEK4Ax99jrsgDv1W4OINgfelDufDT/RWWs+MstBntQRj2y/bv8gU
cYHtHjzOO90ZDNk7aX9zypK0aURJ9jjGvZwYAOwu7MVofqihY+pto/W/C18epnUY
j4Hlu5NTV/Yl+aFQmraoIbIGLU5N8ns9gVeCplRiNzrxnkBiX9vjMh68A7iQZZY+
Rvw2TL0DZhOfJwvBCwMcHXoQz2gb4RB5NjkTfdpIMDZvDYtdEc8ffGvLv/svruLj
UWt33+ofrolJcJJ5uPrIzX2HAFRxOw1WMdvKv6yHccxN+ubFgOtTOKy/MhQv4LpX
qfank945C9vARpDQ4iAz+mJK0ngNQZjQULDgsSQ0fZu1PbJUUXWKH10cg9wD5en0
2/bnUo81QYjdeDUlpqtIZDIUlLiFZg1mFnZi+djwwHS55UUva+cYpye5B4UMxR3K
3LSZPvkluvlC9ZEZ7y5YZkt1GYyoSqv9gqBDIFhMSOwwlZ3IqOLd+tzlpDWEQcz3
SfWmLyVu1+02q7sBq7Zo4aALWA4Hp+c/j9MSfsGNMkmHF1MI2YjcaRLwPlh309WM
SnZIe9JLnACNZZLeBKdOBlVEHGEyuxMUazf+WLXvGQH+uFNZJ6UyCoLxVvtUMcc6
xDMSxdoGz9Cj0Qb4xhHEuFEgzM7HVwhdW4OO52ByDHP1zesKgUCa34p4+kox5nw9
kWO4xwkb3nmKqXNEEjn6x8l1L7qj0L3Uc46w8NvUWgEsIj1d42oELIgFaCjUNWoH
sQFiZjPsbV9hiuNZ5ulcr1Be8mSeczDqaUmSK3k88mhF/x0feDhF9/mf60pfQcSa
0wPi/yf21y59AYTEx/2Bh8KpJ9a/tNYFdJd9/VmQVOvxbU2t3s5FC57Wpj8670Sl
USM23SLIxoV9Z3PyXl4DrREZ3Uvbdq7wNbhzY1jED7wALcMS8QViqUu4je/TOiQs
Q2DOg8AGLZNiWiXjoNvTx+1vaP75dbe09+W2zHpgFV+nXOfyOLfufJwQdurYj0mq
likwxwf1n5ihDF+S51cLUsIfYMbEOa4DJKheylDVKzfdTOvC9fbNMPU9D9w++3Su
kOq1zyqrKPf/fy3vl2BDZsu9HBEVdLooT4q+b8pMKOUzRFJxktApMOat17g6kEob
/ys/Mj3Dqy+HwELWVo7nViIH7vky2UxeYna1HgwkKe42g9h6NEZeYbllrs12YclA
oojbvTEsehBgXpW1R01UiojA37o8zBOVWmT2wVNISH3UKdYQ8b6DY2lCBndRF9Rd
w9k503jfPBlwFGo3J/gEdmctVzsvIQAWfXrg536SL7EbiXwLf2/uSbXTcM7X2AGJ
QxjpR+3GxlaHU7G5kTV/9tVFTuDdeJwuDsAWyE/1/EBadeZc3CYrD/UH1jUqzk7v
6gkiuAiphfHonbG+xgl0iVP2qlUy5SG36evie/z7ncYM9iJJfxyIMsKP3ijtmMud
sBNBFdvRZTzm2HtLGb1eQcHG6qJ7Y+j2i9eIsOPegnKGBUDzJqys6vBn5/1FDuvY
epGYezTH73pIuUlQ6Y0CaXLbldYolQ98SHPEIRZbXIAfvN9CRiOOArCCV8mbn285
ZzqmIqCNdmPCXLtcOlhQk97EDjNq+AH9KQ1MwKVODmH5Me+hYAX6q3+f7Z7kVArI
d2IEnDfMSV4AwH2rOTyuXZp8yFRYQy57qTe3CC1lSnXbFBXsKipRwJKYpehslBtI
QGC3+uObnFG635/+H7p68C/pQZ/TnELz5RCXERApRsSAh5dxjT5WOq4C8LHx8f/g
WazXkBMavHxhxO/QrF3QWu/0ySEj5u06gKv8/9v3LeWY3ramFY3sXFlaRoycosZO
kzoUOcLXvnwRlaLB980bL/jOuBc/TKRH+IatOq2L36oPOe61Z/dUk2nJocl9e8UU
II/mRFaDUWlWi2fUx8Yjhw/FwYCaA+OzoqKuTYLixeqcGtkMlTysYktTuYwXjg5r
6BWJAyfodftiHL4HkgbFhfkeNfNYfMMN6inRFSgyV8oY9aVZ/L6IfnDx5/65VPZ+
GXYyVzTsK9A5X93uV0N3H7SQZqTR7k3SBoEKZg/OOc1puJGV9l2ElJCWoM3Lp2h9
8JO7uGXGjUIsEF+hSSi79QXlxoK5DwKw+QFAjaZI1s4hBEfkFP6yh3M3i67e1jLv
p234zs4zh28cfP/vcjWTO07dVAElVnWWD5j6TLtwybE8+3RdUPDLkcNC64XjphNB
HqJfm6BHOuPaj/ZYgBLXE8NjPJze3rlJ9gStyeG/8530M+BgeUcKUjtnzQpSDbUP
t6C79K6kZ0uHs8dzuIXyaeLnhm5XHUd0cXG8vYAmujVc7kxjVLPVS81Nhh1Du7C1
CotJiJgNHiSyXxq7SWf7TQC48J54nUhy9eBMc0DhD98OhtqLS4rWctEu9bpcntJh
myrIHWB9FkWWRFj9iVupkxaW/xvn5O88omWT3izUkfF6fopqMAHtkT3lPbNfDssW
lBlC7JAvvVpRZkkUxqWrw0/STHb+Bgu+LOADJts9zqVLZQkfNAYxLA5EqLD8QzNo
2t1LG2ytCE94xUIG20GUNv+lKvO6tYN88QAg/L04GO1o2sga2rE58rSqd6pBUqAS
m+WO45rFi0Dc+rSTb/iXxzntt2eSWHSrMUPjU3gdKuWWule2wL3SMup/ya/7YfRu
aT488oDWL6OWxL7SSvYVhgDpNc5vKfZRvvbtslp+O/h1khVQbvaNXZrBGTNd+p7Y
cPpwDWL0QvlPUDO0FMiPXxOFLubRRvlOV5mtow5rNmSbAvreygps45k+BmxB/D7+
bHyAE4h+5Ds+44EzXZvVmRYJp77hC/Z0l9ur7X7ea8KHEIo//7taQLTIF90BeAYU
rzt14POtr1BNlCV5LqM5wkjF5NvG+gkDophLjGfrifOH/1LUN1E7vFoB/2e68S1K
QfGnGnKYhtYg9O3piQECG4T9vDoS9zvwHL6i1eOft93v7ZXmPXmWjOeKz6fUa0m+
OMZLNTvG9EQiBPvdtnB5Z5pwIjuPQDmSw3WHmsmXKds7yVoMnx0wW8CzXtmu2wwW
Gr5QIAoBKiGcdcTgF4tb7R+d5fwPCPHUEwjAp+8J5pUT+x05vDStiLbxKyrYuDpC
+rLoKD+k0JTJnkBfe634RuKzlG+im7sDhrQIj3Zc7o6D3eBBHOehTze8XaPAejHm
7REbf5vOf/DWuk1ldiK1zuFJpri/sIQe77K//RFZ+aWD656vl0YAzDkgjFqLrxx2
tdd/bb03wKMaD7EJSHtpOTp01ZgJUJMCGBFkJgyYeazo0WcnNqUDysHaH2bh2dnW
/SJPwmTWsZeWe3uZJGnoF4+m3cq9cDVcvMAzRkgcSbFxUhJSa6uBU7AWXoGOpy30
rGyA4uWCmQ67+1rfaNQveGcd6o0uuEQL22ow7KCbPinKXiDqs+KrxtiajkhQ9iMu
RGSHJyqohOOMacc2k415CxaPdQYU3UucBoz9LQX3FqlF7Q6zsCS/pO8zbQkG9rwC
55esfGvHzzXtIz3b/c1cu51krrKkHvPdi3qB0z9q15w/g7vExA53r6voZt3X3gnI
Dk/Pcs5OJXhlCONwQ63UJA+eQxjEAaIZno0mVYQPsLKdLOyGhRRXD7suxwRWMR7a
imuWgbdb05C3gL3I7JGfcXRIwUv5heAyu5AsyPEvzYeomKVmdBHuOuSIwBeA96Hb
7FORH2fjS3jcqu2SDjMBYRu/S5iFUT1kDDOCSH/p4adtZhH9BKpb2bL3COYl2Xfs
ARvViCwDdHoIdGWHiEHtpU0cEmxpgDL7A+AG6fPu6OhXZ8PDRQXfEdxqaWPKzztb
vM7dPOjatETRzuXZ3No7VJZGmlOcrBUCb2RWelCmSWnEJf20V5/NDHtllq3NfkGD
rauNxwp0eHT/XSHVH098wsKl66yfkZ+v6Azt+LSsBGgiK3ZdT0+IY43WerT81tKa
Z2U0ClAjNW4Kv0MRvY+B/fLy7J0+1TUR9CZ/g4EUt90KgEakwJ513t3YtKtuEsy0
ZBvDQ/otPVUVV1mngBXdQI7eKivXo1xSI35LVSkm/EHLj6v2PDPPnD+cJp+davGR
g63W8La5bXiK2WD8nUUjod7HqZHlRiMldqXx0v9iVivRh/UXz+5/5fGj5Gucmvs6
C4CSyZFXa+lmKr6rIUX2fZ+0QStoxCRomR3ADWcpwcKC6KIlJvlAKWpX9kZYygXV
GIBFXNkwHok9y4G3toOyqslol9Zhr5l6RXycy32oKOxBA9GOE+nNIeWJw7WBLNtz
Mn2XS1Lq6SSDGIgRMAB4/eV2bKXVByndiYJVcBdAL6arOgFwNYtrQG4wPwqpseWr
hnzETY32/FLCmKhk/jrLlILzC/nNJxxDmNO/GkR90v/kmwOFrJlPhoJcKc4N3DZN
t2lfW/tUDF8FpYOqodJQ7ZwOV4lLwAyLJLryj8YYCk3QpLxL/HQHb8CxY/V7AXil
/QXrQqbajyOtddjkhsZGOK42VwKe9fSOEpmuWVcwUGxvfufm9E/76bMPRQ9dF7XI
iPzIx+YOtpi2Ne5UR4On7CSV3RnoTibrOkPpOUIWz0Yz7uTIMi5bGtfmaS++Vw6x
g/W3dc+OgH15nh3AK+p0WZWc/yfD5WCDRDFmmVpYsMdTD9j5d3RHCeeUwIHHUwF6
rmjcG0Uec3o0106l4jDXEcjg05IeGdnNXTB0KbZQVxGm9xch0WacX85OdvQ9IIY9
tA0sZ6WNPhXs4aMxUSjDz+QTdcbRjGtWIQdUr2z4hJZux0xWMsgW+xDkjU5gs9+W
QkUrHy78FbSmCrkumd+dOTfwSju8lGdyxPCqrd/yh6mcpsGhr8P7ehgKwq/mId/S
mmAtJ+eZyJz3aKxGgJJqk39hnbCgxyO+5vntGn1jcBuMmn2Mi/jxmSTVhdJIJQzE
GzbJSBQN6mgzs41jUZ1m/j8Of+95HA0O/Zueq2za0Q/OOiM4ODESe1cF2cjqx2nG
pUx57F+YSo33R4k1aBmy3V+UXRGEqmGiQgL54Gvh58g2m9jDH8MjG30dXiqDFMKc
/eaGX/Xp4ZPB07ldo8Qmx0rZ//rF7dmnkQH2lqt5GxG3dp3gZilSgPe8B4bOZVJ9
yql9BUg2zEJ8izB+qIWhj08IBXjIjfngsMXZDRyOzgVCzsdb71dY3M16lP1w+SJy
+BNhFqmxN9kks7cUSAZy1EY+OnTDt4YliCkY6mqui+IAst0n0Yv5m4YFuhfmdbGe
0D3rqrxs4MQEvd3tu819iyin4U+QaD1DZuJFmCSDBdZn3Do1N/hOEkTnxfPDDHEM
xunztViR+tWbbzchfNewfeGgduiphI/ARkFf9ANCmiLm/KiE7t7e+7CHRG3Ui/dQ
7zhNJUNcnLf4IH2bnOp+Nt+R82H1YADalmSU5tW/BBiT3R/HUvkHeZuI0wDjmRqE
J9TsqHHwiUrNphu/LZ4PxtIhwo0nL6zHg/8ZqZSNT/SfU+xAmLq9GVz29V1SWDxT
7hW/xY6Ogs0reMWKv2zy97utxWKOqb1UXt8bx6mhlNe4chkuUw36UAJh+jlNp6tp
t2VXAb7ZIReziQTQkvWmJ6C0RoWlCWds9o8UYUVkb1S2e+RBZRR232B/aveb2Xg+
5TfkIAYwYefBwQ/TNoeNb8bdtQatmsMo56jk3yc1ayjK/NX1TAQcQTxNGMhMa4RA
YRGXp4PiMj9WPLUEmlxdTlphZOZuwEllSHrnmW5wwvuTEvaA34EmyriiJRNvkkT1
4GQDZC4d7wXz9klzW8UDyA7KB58c5R6yIifRpY/wyXPqiQGzDxNvg8jugYLzGrTx
fsQl/lpUTdg3sj9P2tecMyt3bANr2rNCqVLFn+qUueKxE8QPu+kcWiI/HHfcD5lq
U/FcFlTCXg7RTJRw1SGyBRYQRXhd+2+5lqjlzdFHvBfalHtYPdP5GGUPH9aYJxC9
RNytQv0gKdV5BqfK/58RGjS4ggEFJ9CH+eouy7QpoA0GGyLOc79NuCx7uI0V0eIC
ypBUfUP2lpJJ+OPJn2UIrO0dtXjtRZcR9sdjywBK914TuzrYeAkykmCPfcsK8crn
AXllFv+YMkS2m9swRDJYb3M2hpc44rQ1chc08OqraW7cIpMn5zLnjoqAdMbz5Pec
luO5Ub1N+VyxtkgnRorStbUqY9voi45e23pkadHV6QDklzwgAjHVYUZypyBQFS0l
oFepTafKU+nfayBwwvuvfd4KJoP3qC94DLybMmyPH2iwZPz217XQecIn8L32xYwe
BmExnodoNMz2Vqwvp8FiRPNyAi/pONLJD88rkS931r20d9fzDpq14fuscF/BsTce
byG3D3Mykq32a3b9u5A4H/RIdfWfhDADsGJKyXa9dF1U7h69PjmiJloa1S6qyNBY
oVYMBROd5Ikz/3X02GKGWxRO+ifhnnaVogGmEeTUw352ZjSSCvbSRzpzQ2TBMn48
50ZyepsjXp3dXudEKUtSqSa9W1kdn9pKbRijMtR0rsM3TDOGFEsaexdlmxYSRQXC
zobqEzdbzT+ECPbKozLXwyoXGYVj/SUUr7lIfIJ+g3XwTaPzdV/JuktQ0Q7Z+Ovj
+qiEhbEdUaNk8XNx0m97Xs70tGjbIFqrysa0G3/QyBH3Xwz4hyQoSjsEa6nF90Fr
W+JNlW8vflp5Tw6rH7jYAHzLc6CRO1ZaUjFNjosqOMUwhtH86SJtCNJmyGgWmT/U
iiE7HzT8m+S9SESqZSn1/H3AC2l1KP8JSAyR/iaVEABW7BbI+j9SkAZIxDMCmc5f
AMmPeBW0BSr0lubnghBm60sFn0JEGNXvDLGLBO+uM8bjorlV7oYYsgL6GEZN/+e8
e85PGh+U9RWswUwEA0s1ZNYv7BZGlSRs1mFB9PNfidDS3Ga0mr0MIx8JSi0oz5L7
zsX9AcaTDrEsGni50dgjZDL35nbUb7VUdlAqlnQDTg/yjm9kHf8HdDbpmp8Xc5Pm
wc2vC5s23IAUAfiaG+gfxFMgXpUGIyaD86H7xzvWd9hOGKa+8//HYlJNAxhhM9Ab
I/mD1o+eOe4LWXAu/eqDRFaZAtUFgO6s1Je4PnD2b5WCpXkTjnFfJsC4TYU0F8nJ
O7AdcaAstaeE3u2EQjDS+9r+TvgH6+5z8gpFrweJSTmaPRXiAWrSiK1xsaipm+ZU
IVq/MyC8R9cnH0jcxXfZ3irAg7li5obqaP2ZP8KqQcedjJEnc3h9Yk8Rp7E9Ik6Z
yV8Gs/+gtIzcRXkwnlDTZ8SrqmMDg8BkSEE9DxcsYH2LglgQ9vjhlRVe1MCcUJjG
cd2fKcAKMIVTqYKugyajtadFHAYsD+5bv/4LolAn77wHdS7eJbv+msaCcsqp6d1p
aJH+FKONzDY5Q8vLtN8pSdjRWykqv0NZTCxOuBOm0CxyVb3AUUnkRVPyy6d98HRU
xe2NFRClnB+5XRkA7Dq0sIb9BTBaRP03tiTvbH2Ah2sSipHEIXrRzWI0wer4yKbW
SmIwcnOIPMTTPGasaFXSXcEY3ucEKaMWmvPNWzNg+3xiTQoTOOTEthRzXb+OqLcz
7bsZOp2cJZwtbX21fPlz2KvKIQMrAM71YyB1OsqgyC+Q4yLZj4brXNSOjtGjAucn
nySavT1Vzx6OeTZ3897f8K4i63Ni01t7iTrYVZslBDhXZecC7P29tCzhW2RPB3xZ
CT6MnTnLB+uVBSKgnZyR53Uexz9/TEfgSt+xT/32qaH59Mg7HHaPk3QXQEP1K97Y
1kiYle7IexWMsJ8ZplS6SIGZQw274UXhJcXFbK/T1JJvtvQGMQLhfpg7013zG+DB
+cy8BEpYzcet1ff+LieV+CgoTzvazLW3b25453/thp6lawJ24BzwrpIlvTjsFZEr
hKJ/IGX7DKCpuEKUY1lAivfzUM3d5KY+34XuUriY5Lj+1EJ6TrDFSiiXP3kdElYp
b9kDVpjP8wQ1SHASAv1C4y9s+oChfsv96el//98prPRnDmHms7sZXOSbhaCNscTb
Eo+26IX8WNzfkS03xzGb6VF5V0AbO5Onz5+08GRAMEkLYlRuwQgBqroMyw6QrqrY
sGubYBzbol9VA307oe5bIbFgS5bcwcLqWYVwETSvmg/yzdguq75iUiny7oyPGkUZ
SM7gjKdRx0itcUN2ao255MPNoe4RF5sGFuSuSS/KbJ3KKqZnfHF3KTd2xuDpQwcZ
AqWfLmFPTPTuC6eCmBV2HIYtybck8e5m2apEnZQZPu78HSonmJrkIC/PzYf7rozO
F2vjbVgo7Wn/2f372aBUVjJubjibU5bhSjYxcCFb9GGYw8u0+XKvCRIy75OV6QVI
F1PtAD0No0jpC64MPF6TFHOME/ZXEZoj4qL7VJcvEWTpxywtXnISpvlN8RPxAGXe
dr4mKJeidqY3m8lO8nme7MhrpnzWm8UPseVaTfMCkdwjTmsEK+eoBSk9EqhYDuVP
YNCeEJvdyzXZUECttzV54FY+U+IlmBmyOVA4IIlwQrIJskGEM+Z6MozusG+cjEbb
xj0sSMzp31ehbyorYFIhz0JF8QcpEwDyvWPjRLJj1caE40oInppmu6yNypxxaO6G
4BTvHxOIeW1wmM9IW4+AwQF/Oyu7v/CaPJcsPP15jJFCJtdW4VOyWRxDpSkivv7E
1BgffNFynrK4TBDsGPc4AcQcu4wEn+j3AHNMxBos6A0d16WH4ZxmHNYLspCAZ/Ym
WvTjEDDIshDgh1HuDCy1uXZNszoYxyut1RwOkrupX4BblpKIzVio+aPVjQWkzYvF
UYmPOuLUSWeGF8yNg92yAAYIaMlnICG4MzKmKSv41MbDPBlprmkHskV52ps1HZIh
BE3eXXZ41vo+yFED7B7d6tQGXNgEISDvqG/J+oxYLqoHa4fjw7yJzSGcAy4nsfi6
R101D7DISZfH1tDmo13EaSocRUr0UYZKa74fsrjDuBEGk1KfRToQgqRLtsIW2hb5
rKAVg9rbvIijgDu2WqHVIo1hDTH0hwqqP+iQNTYbm5sDqXp6KpQrcqPss4VWzdbJ
JFyXlu844SempWwKsMvxjh71fBS4bF8nq6XFPoY1j+4rVJs0OVrODSM29cup/4cf
Yj+ajH2QMW3KeTc3n5nE9YqdTeDwYVwmuVcnnOtaipM0sntoGETcIL6AUvZBK9vN
b6RzVahipJdkzjy9sRsYpL09FM0m7gLCzB8OeF4/OGl52HY6GQFZ0jlUExQsmuGO
Ys3AtFXNvrqZ4MzHr4ZrPL0Jt4pvjKJusSX6iAxIhATeIneje3NDfj3Ba+4Cw4lI
jakey2hDiOCmvtWLkqW3q6jK+OTLMEuycmkle9E22ghpsUfg7KvXu2al50h9pma5
IHAkEjJix0/o2pqKy+mQYDFj0z5FniBoQRPyI0yIvOLPWglsXSUUXck8wubXyQYA
GSnZnG6MJzf7bpgVkCc+NCzFEOgZBUcBr5UL24/RcbE9vhVlZqNKVhCa1psv003b
ukV6isW/KTHeL76hjYXAcqIH1uBxNgwaP7rL1T0ZG7J8XL4EN/CXpup1Opq4M2T4
xs9IOk6pl7YvaCWG4oMNeDmXsqpW+wAm4Dm7pqG8Emuz/tOHJcrFedpNr5l540bB
mnh6bxVAIC5vB8CyHigThUc2npg/2G/ay+iC5sg/GqqBQW+03Q6LFggyOoxdcEQM
jCb4U6tauL2CeOI8NbaFFdBZs5olskVmdWnlUdQ32CkF95w6DPQNuyf74JPkYvaS
RCCe8N2MSNpKZEBBXHAVm8TyfnZjwD7dL3j+tUpBCpDEYiRfKAW9zy9NXN2eePX/
b5ABqZK9JY+lgDX3VfmISjCCbVUBbeHh6MGhCT6MBBV5a38UAS5mLKl6xCjz/oOK
6R7f0bC+Ss6br35DPNiCOV/65f/QOslSVqGGGIjfqDc1y+VRUS/3F//7S6TrITei
vUYQAQNJ7Dg25xhiBh/0kPurnYY3zxVfkfZiVM+9a3478tj7dTPXpiE4krbr6ape
bGxbHGzSZOxoUIUJ/XUyVQ8pCSRTEixrGbkEX/TpwwL/cvUV9l4a9OQrlGID4I7o
SjSb/2SCPUbgnhnH37pTZWEmoZ0lkBvBc1kqN5XcsB6jc0KinWol/gCOQpwa1IwP
Aqu0eo5sDSqE1wit0KlOhqHUtsi1Sc1mDbrCswlBnKMZ+xey5BgySNc4ab9j0twd
BT6JGEHoqmrqdSkcM6kjRdYHCebGoP40c3UapuCzAhILtSTQMEWuIqeIGO0qNHTB
sEL+l40BBjzskWzFWPo9Q6FX6jFoqERW2bBaD92Zn66gdIdM70b+SUX404wUaRI4
Ehwm8C/DocacA3YbzQDIfJ892uPsSWWHwWDcblbNi6HGEk5d0haqALT8FZBCvl4C
lkro+zcYCCY86ekgBXoaakEC1x8Z9F84ytb9LvworfHPSCR2nIT6t04PP0hwa19l
yyxmAbMTpMtar0GbqM3Od9c336F5u4fx6coYzTsg8kIw679svMt0cx50HLkCpmkt
LZRiYUhVezQ/VPF511NFXN7QiwMmwoO8dJgJtNaDVryv0H6dx3v2FZ5KdO56YKAU
9NHbGYkId0+74L3xM1LuAWD4XHe5wLPJpCFGz9KZHPlg+rRdPZHGrmD9Uof3Scqy
5VRx7AQWBZpxqFL9vRyfciFAlHqAhvLgSWyLfPXwLrZgDCGDvhmvkC7Qem4m5Y+o
FTeIGsivo0apbu3vP0Kg6WL81MPaJwepJAGHFrCdqqV7CRfQIgcqrlJw1C0rIi0L
WEBJv+/ulGDpo6iPQHFig8KLHgCRHv+9OwEX3TwIm659N7RXk5uOPc0/dkBGLz9K
J1f/NXdVbmCxA4GqCaoBZi02X71m+AILMuvJKz/yttQZkNDB9deZVDMSaNAByldj
pPR8iXzBp26OxvOTHvCfwPzOK0X3DyAqd2lcUjr4UZnEu4/zAR+jOfiubIJnpnDj
2ZEw3FGN58fxe9O+E5xCs6PSncs8Lak+eLl7OFpq4VZH3/niEYMffYYAv7juMNBu
B5rAB0fd3Z4Q8cRez9mE8EqHhGOXinwI6TJ35l3BD2/yA96U1YqDRRJA/78yis9f
2Y526oixDPQTbkVI64B7LlblAn4Lrn/vptIICPvH4ilztSwoYevml2Qryw9XFIRB
C//I0eG1HVVMIlhHhCanrQ39Z5JqfSTayybzj+tAoNpUxC0SBOYihYXBNQPgTMAo
B1dF8ES0Vg4BynF8sP1ySMRK4qfOBqI8iE1QtMZhOuQeBfoMOzvvfc5GUr4QEd6C
8W6K1EFB5h9vEshpqUmWjANOHsNPJ/SfsEKSD+gxOfdeq38jGDzeAJKHxrFwzhb/
XfG+B2B2l2tXS0p4EF7/KuAO31h/jfKDTz+u6V8HKifmh4l0dmH4WZQ1OgT24sIl
UZC3lNx4HSp0J6Iw+LtqfFHb1mMQUAj+BWrF9xowT6v2Bf26jrXUmCHwRAzgqFTk
IoLsERo/GUU+mQKeziMls3K52AVit7rD9/ThnlYS36gZYlt8qrzb/zqLkc1aBJ/R
ydtf70AFtniAZIL56JTAsHvsnlZxHk0zLyND9v0E3vqxQupi3BvV+/9HTuezLyxn
wAzp8T+CjBnu56Kj8eyKc0pgZqNp37T5ya1nKF6z3sh67D+0fm4jE5wYyk8KC3Ig
fRyHkhyHtE+2ySxTiWMDhF6q9n7UBbDbdm4litetX1WrxXz4m8Coqh1uS8Q96iEp
XqgbaCoBJj0o9gAM5bF8ind9mCVPnWi2Ls8B6PAgUOgw6MIL4FiY2gQqnDQA24fH
CshILM7eTZgJmU9KJsVXh1KS2IAYT+ufRlt4BZ2Ew+DWq/uUSpIVsEWDUp4oFmYN
iEsaXMnF5b8wsB6oiUsxplqjOzzg7B/L+fXPuXdFdjOBzYPk8QAmEfWTrIyBXzCQ
O7w5A5JEiT8NZK9+YWYugdQieAdDkGAZGxgIlfYcDV6OLccdzK6YQUM3fxNPa2Fb
YxzKBzHM+tsM/BNOZnVm+4/zn60lJuZCj+hDXmnwHwFAVwzpzRhZffhv46KV27Xc
oxjoKXE3/Bynug310206H7VM/QWqrYG8hMuB0yaksO+aTEu8ThsMQpJ84WW++YGV
eWrexhNB7GW8W3dC+elXNhNRErgE0CUgs5sXymDwyxKnmRRPvtFe/lVQzBj17H0i
ZemAJn5odqoVscSrxUSYZr8Wr5p+YuVlGBgzYU/DvdTimV5qnNT4JSaFClbCjRRw
CDkrdg+42Qh+IrZ4v8VV3Z3ObDLnhS5GrQrD3aAHBEXNHY/nvgQG9jKONeIVak35
sAM3hYn0pseCibU27uSirSesubsnTcEm5O7W0QfI6vzyzlB1rR8ieC7Q0BvFBd51
nvS3HlfFz735ao+pGXCgLx2+dA5e8V2Eypgt/l3uht7kT4Pi7EFbZJCXA5ZBvYpo
KXqDz67oy8R2cWsJSo2/Wiy0FyBlOjbKMrzNH4BdQYotZbkMJLFCbaZLzXyo3/nr
nPXkbsgPkGW3hZB251Y6Q9EMYGUNF+B0r94C9ANzXXCJ6rPGgVSQ38f+/b0tSsei
lY7g9WWDme+QS06DuiDPYIGTnbPMl/l/7FqjHraUuS944epCay6nYpekVWP8XWoI
9kVtZGneLC2cZilVmP82WZbnxAmSvQIjcaqgz+c6kJuj1eRBpkOMAHxlDRyJCGBY
NNySXvMybvtU0Ahk2lqvxM7saWKewTGMrvxMYrKEPeyGL4JqDVp7oAQCw6FHuAR+
Vvhorq805f57CdGxuACNocNN2ZDKvjRnO7+JadvUcsAgFVcl+LMAhXI7WGP33YHC
heIaVyE9WZhIWbeaFfjd8oIp3N3+MMj2HO9sZ84ejqWSLCKikdhm8FoVr+LftRWn
fL3uEqvehVkRLHeOwTDFYDnY8cYAr/6YEdNKBIVTZktntL3qEmv0CNykI575P0pK
mOuxaJcVPJAPHU4+goxn88qBO6gOlnxB6rTZGgs6+hAS7qpTSR4yuFxaiF3i1aXd
FxOKfNiW+ioeA3zQxBG5wU0rb9NOE/Y0oAzOciE5MnBEWxfiEltmA5tnrwp0r/+K
IGiqZxJNUiNEvOO4+YR95BCKVpP+bB7/Dsl/rYcEP83CiWDX+PILIp8WSP7ZSXZ4
Yyu4okqjpQN09RNZzTjxhoepUXOqFAPEqoAOkm3AectHS138tr5ByjoLTTrDNt5v
MyBlSxhGZhSQPkfyy/XZWJH1RVfNUhTWCIeTG+qMJ5AZxK+pazkMkhc37KMHKIRQ
FjtCRoSe4nNiOZXVXr2pEaSoRJ1BoAne4LocMDwfhmpm4YZgHa4UCLfjAHfC5hoK
0Q9QLU5vCK9/wXd9pdUDPh8K+SMBdcC8z5icdxb8MgbjpjmpRf5gpMbwNtJXwnXT
aNJIUzgy0mCWlRq0aTpdDvjp5QyNOAb9PPnOu1RkTw1TGJ4BWWNswQjUWcpxThvK
VTLfADXz9Xm2qt6luj5ONvTj+Lla2lKgCNj7VNz6Ox8UWH9lX0ElkGOF4BeTioNU
/SJB2CpiHoCMdFqqvXZ2IDUBfS0SpwC9Sngk9GRSJQnVT6vTDURf8R4vykhHxkmR
eQ6SgX9ufj9YWQttLgjRZXn1lgBzWf+W77hWxRzqvyJ1ikWqCuUZ/Mjb3L7YD2dR
ZTbT568+EpIPJiHLhU/H4SlvOuN4QOovX+sDR4fPD9bMRn+8Hp9u3gu88djEeyvT
1hyBKpC7eysKOTtzMxeyD+atpDvjZNpoMEXTRR5bu341PEoEGuQ730C0EYLJhRqT
na4tMSdc6ZFTuGJxL8JVukAGW0LS30xDqXFITR+7bEtJUr7u3Fy/rC+jTZJCUhNo
umcIKocM3Uoiy/Y7LknNke6OeJVPz1Vgqjq804V4vn4vX9KnYdv5f/7x1Aksgwpz
UU/haNiikTeS3Fns3GilyUtGEQY3oXTHntZ1+vLYRNHr9fl8TpRBpswiudNT27gK
CjkimbXilpJVX8s7FScoAkBSbJPcfQpA77yWBrUaasGqzBL3tI5t2CI+rxEu7Gyy
fo6urY0Bc8YI+IrRTPM6QAe7+SdE2kyyGvtOgfJsnPbqAqHwsJGa030I+9xPh8xB
yIhiEFp/vdOeLBX66gH2C9NKEfVboddaZqLPDeIMb7kbqDtuR/CsggHWj6sT764M
mBu/y5QNWgUm3KgR4hmNuXv6UxXbbl5ZMVpzrqLobKm6MEE2q8xhiQwONvWAUo2H
XTBAWR0w60dzqgH4exIAZr0d4AS4QmSFr9HI+xJth3idghAZnufVcbgB/USspFTJ
lgsq3IzPDMvcG63rQJF4coX1pc04wrELQqOklcCdzRjy+p6rZSOYLnE+bjPU9Drr
zMn1fSkfiHFIkER7sF89xRxvGOk06YhAOgnmu0eJnAwUCuqzPN4tl1DeuX+Az4Um
3O4UzvsmU8duGepGa4g4pTH4KVfIOJfGHf+Z0iRgM3f6n4kowL+OOBDhoyA0xSOv
lO+6MM1c2SxMEcxXPtBbq/PAsCcsuXBWoNz6nCc4FNOb7sQ1XeNv3XsTbzgD5WD0
5IuZRt8HJGKN4b2XVCO2GrsxU3QA7e77LidHB5O+iBOmmNjOYlMktbMD3gHZyDOX
x9ZU/hLTgQd0G7qlSAoAIprPYoixkcAev81ETMCO5GeZIvZQdSXmHWPrnblfoDnm
ex8LlgYeJFZWjf7fjk0nDCvTdh0sBz05AmXIcDMXjF6zghbVpuuU0u8HCFCSZbce
OjB4rRJDaHTEU3OpSt83d9qGr+4SaJEpSDBYLgue9Shlm7lSCc78PjNqrJ5Bc4vO
7HKRX9COgaeXWj5P4rBh5/zFZEmZKCwWOUay+Vt7mcB3+5DKky5CXMjT6ZS4Qiw6
R0qhE0ylTv2FTbk3W/OCh0JTnqJfu5/Ipw8gjEq0hZAjvAT3ujXvBo6rqD1nMouB
Yjs6VOhBZOu042ZlpSU5Q72oP9C3O6HsYtl8iHjlt+HzfiNBnzUwnmB23w4rBv35
Ayv/ijhITQu1smMcgy+RKE9vMZ2W68dIgGxzU0HeX4WztzvLp+ovUhFgXwt1uDPy
At1HtINSGp/aS5Dv1CdkOV21zaXmq7bmck4VnXC06n3rYvB/d/uewdTqskVX+wl5
irL8+86FNVJicZmpWi3ScL3Z5Isito/FYT/nqH5HetUUA3Yih7rg19o21nHsCebI
2ytAzltih+8x6sWovwyC2MjLW8PKXvWoZBg/8Vo7MzYk+LfdIr+EbR6z8gEnqK9X
/qNzrsTiC0atEKv6mHo9hZyRGk+YJB8hYtZcR35/eBtEig8xVdpgIxTD1EJa8l74
08I5J4flVJdPI+QMQc9xxZa1QPTCBvVwAUjThmWeL0l0mSNGHNa73KDIFBuKoAkm
0pSOKAWQgLSUXWXSfo2o3aJPIEkxETmUezyyAwcUT/53rhjnQZvdzI5fvHd/N2qb
5dxJLgxS1rdRSP9jJvbG5l8ik9IrLAmwgMO4BZ+R8HCXPcubKp1JOBz4KDMffe24
i1eLkvbM0x2OsYpCrcrHJt5TF5RNpLtKBcgIsDMXb3CTerr8ao40daCTvHNQGVaU
exdMj2oDc8KJtZVFaJLaHAwpO1EwMwc90MgO3ru5IbQJNZiM3S5nRmxi/jRXbtjm
EnylxAX0eDkS75uFWXVJ5yLTtm7Brm9qCEhtt+T3d0PY099d8guAitDuP8y2VOUC
pOOuU5qcbCLupnYdFWu42K9bpE/fhjCMCIxwl7yL8kaH+g0rN6gcfpRJpxO/Ud4T
exdu8neECBWkwG0wnsSfKfkxS9DyB+K6GYg8lUysKhJq8TuwYZzeYG3Ms4QHi/ch
BblSMKfTHqmnWYL3s0L3cfcqw8nHmbTcQJ2ltCtzi5kBeehmwKl3Ru5ITn2qJWgh
sjmt5tZzF0C3hZrIWHmqJLVdooHfN3IZhfNAvmBnFySww+xEUzmPMnBKaPet7rcl
2QxYoc1AR7NU0PfTHsvk3KVrzUwJjgQsf4TUGlWbKNRle+IHc0hCAQn7Oh4oMf3g
29+gMlxFKkAzqKGhSoaOGCXVUr2u1ieVBauWtor9mkj95VAVMwhSjy7lSklTrP5U
45IZq0MjJdipfuskxxwir0q4VU69+PjPVoJWkaxbnqnnR1YHhZpoy/grAGLbPGie
7Gk/zYecVtJ/Dhy1J9vOlp2xe0iHuPxrqh6djDSQphvCtbMYCi492e1n9ytZkehC
X/OW4mofFMAa0aA0i5L/KgX7ro9DN+2AnZ3ZFg15vnOVT5xBNOCLocNjGN7MufIf
2ZU74+ObhFdl9G08YGqHYpqxbZKw37FIaCjsHuzCLJTvymEIAR9O59DGoUoTiwii
mvaC3fe0DA+IGRw4KUCWIITu5S/uwro75RmNjQ776a9pKMuNBu2VVcfiNyWLHBGe
NPdZNoAXX5EEYGo+2SeUXaeMRLRSSSVZSc5HioW7eKCSHeCd+8z002RRAMunIU8K
zgcIZYGF8BRNRbdzUMd7VCZ/MqklISd+OwrZJRv+nsN3KrYuWfd7AnCo59h7D4iR
5fUo+JGUgTlDbgWdSt9ekCA6DYvjWwA3QU4vJ0LUjBEvU7GY+lC8Q9YdZAcE4JzW
hs7joiPlI4YYmp3F+9mg+H+SaLsYkL32jWaXABTCl6nZg7Qmmritd5aSR0Gcd+Ks
icllCuGeAiUSl90ExET2Y5ZQC4wZ+9UiaA1RQIIx8Wp+dTwa2/Fp4r8BlKOZzj7v
rHpxnSk6IK0D4L6rvHF0j+DN+btQ/ba+a4GrLCu9GEyS9L/q1e/ttfHwUl2Bqges
mkplETRiQW0KdnEDcqjmWVdcqtwPEfsh/BfSXEOXm59HtGIIA4jYSso7NaINjHHg
bQ7SllTqfDUZIKPExWNGE5yuSpSR7ZA1GW3JN03R+UF/VJiZZrTBFLodfwa174PJ
95vIQMq+8mJBJtrvcLCaa7Y0xZ4M5csZVWjXo6oeNYJKbK2CshnLL6loASit/ALA
FG4YfrlJoPSBEO95s76jLvJPATWlJTSS1vGN8dRhTpS9y+XFc8M8hnHntgxH0b0h
rA39SxCvl0PbVd+txSCeE120I3iI69JQZvAA+feT0wMlG4naIoBMvCR902ZgLKmq
Xj+CDT7fq3jvQ+aK1DVu0LZDLQA01rcNY9eVjGK9vfiDwOp9ac+iNFtADcWehXQo
FgG/TpY0ah6UmxDcnKlIAwQQvB1svd7Jl5xs2oHaEfFX+jMhrML8aKSp7H4SUrHR
0HQooTifk5n1eQHk4IopXe+KWal0AAKrcnooc+0zTkDKCcb7KugJYSTMAl87O1/a
6Pei/MWifswLyKmsPmQJ/iikxraYm3H2GaZSx0PFqJgG/vxzJksVPk/Ms7gdMVEg
KqBSICgvAinJrMC3BKm7v7r9e57sCWS2A7owY260Gcv0t8H0XHirWguc0VAGdk1S
K15uulWjM8Za41zjMSDr+C6UZ7ZspgB7beawXXKR9OJ69CripxfO+JyWy7+Cbh3/
flCL7zVgyP6ZkavNfoDbKkqCNiqEMuPDy/eYYO/7vFVU7T120n4Ja2L/qgcFyvN2
FTM4tb3N6olWuuP/Dse6owuG0kHi+wAwa+yZSmweHwuRPKbL7ym1iJORsZoWp3GP
cGajX/zL8Xya25CjCYUoaUYS3t6zN2Wq55wvy/MqgsGfbwgQnAwyyg16jt9HrvH4
cxfxyz+YEciAHXAqnT5yRz17q9L8lesrnIevV7/KgliCO+loMKHTrrNZqkppsplV
GWGxSBz1afxWBoaihso2czZg6oqmyLmZ0C4U+jPkaPet6fJofo9/VFUuBqH25jTL
JJkTAubkrznkL/4Mqp6IhjmYiFbZOQyqKoHMdNWFNvKrV3eHfNE/Cm1pPN5xavTX
LwwEl8KtgA502so0ljR2jwQc9HZ/TOooP0WEjeWRzDMH1iCq+av21rTg3YcnBPbB
0RKLdOTDADMCJWOuzJgGCVNc83Ct+x/xI2kQmpTBcnU9qSZFT2KEt1IkYC8+2bDD
pXn4x699gILaSAX1bJKYzTaUBiODPDJEc1ZzsJfjVSTxWjA9HOUSqUB77HG6SoKA
oIVRWmE3xFhn8biQYqkowFPMQWh33rh/6PQ16rgZzyELDlsBSkdolE1NMiHnENyt
DY7EfJI0DhWRaSupQe64VOH+1gYP3Z5K4BzG7JJlapaNd2x0XmC/twvLyEdBa7Zb
bQNmaCKcsJuyO4Nls3T8q6ZEDE5FmzvZPeU5TtKzv9CXG+xb/Q0C/m2i708EvJnr
QHJE9hXo3q/GagRCbf8G4kNf+djeFKf++/uFtdPARTsuuPXG//1lI/dhhZt3cXV0
1ge68VugPVPeRHbwQ5dELjA6z8Q6RNfswQhK1AebqxmaVYfckV7aOOFwQA+jYsBj
OlA6RLIpNbRlqqhzjYI9XVXf8QsT8Ts608rFTYHXMdsqjxijzSIWWFcxP1muqCwz
tvKxIkIb3TOcVZbL6w0ZWsB5oFrRmaIKiMdIW/QDbfwMDtjvmqMB24jIJjFSvJjs
ODOHT1ZwbGfYOPYVJDI/vo64bw6Q1Z9HNkKlUx849+8KL0hkGQGdf4q7CRbczMKg
E/Mjsf8Nyam6RWUQTYFBlb4bEKcz+90IMC/8LNYQoaOcxFiRfoBJGgzpyrbSVanW
oxDMK2sT900d669snTox8g7U8jZK0fsYr6V4XHPp0ID6n8QNva1f8kzYn2Bm6wKX
k8R3NGJOuedDIRYtc+VK6QwvI90NatgalbaJ7zNXaH+dsSVlWYzDly3DtTpWoL4o
U1Rr5M51f4EED8u27ensFIxroiYZ95qTPxSgovWhT1nBevS9ZuowOUm7IUzadQjy
2x4LburPvJr5D7psv1QAGAi7dJh3ZrpTec8Jle+uH82LI3b8HMAlvqnNIaIPR6GX
8+JYAAwI0s6Bl5oLd1vg4mU2bFGyRYmieD7l/CVHGs5vd2vT9y7X/MGEQmwnQPCa
X9XET/gSDHqlCecvo03wXNZx1ZQfsKyfrBr0/h0zkv1CJZZHBlURkEFPMKHW4NYN
l4gnOw3quUYChaLRL9drn8BdpXxGI03vgIVe1viwwfAvWvkBZpzXLUzFBru3idXZ
O4e91eGqMGircKFnwAf4MFdSqPOUc/WoY03TjlWgR3KG+weqijXoU2evuX9HV+XZ
s590Z4uwzXfuxoBTsG2bwWirvbxJmojFlHoKwTwiyMf+M3BssFkU+aTQBtlKWotP
1OTcn1i4Mt4aKfLAUvaNFMjOe/msswv7EdRGxI+aSJxD/CKthWCHmee3a1zrfYhf
k9txi7hyWRavbTNtK5KK8crOY/qik37kJD0iwoFiT0QMuAvNwQ8jK83JsnpQhSkV
DojbZnnAIGMz8jExrE4dKxZeHnX35xtsrW4fPsT1xObSX62nx+sqzzeXQqRJcQ3X
rioX6DmV9sGQriul4A1VSIFMornJJniTmV8IcxJIwy/Kf823eb5BXdnCYJrxuKHC
bZKMfqNuKlFjzRGpAo9HOG41MOLcm3JFLRJFitAYVRtAqvhoQ2eBXXWEzgnuUzwG
7iOPg4DqdPvBbsdz0NlcdW0ldDF/Mrkia7K8XTWocw8TxxbDknTjBS+vGdFWoZOn
AnQ5raD474o9rL+wJFeZfamtANanhn4mHVi13bjd/1eQbN7eB6rcz1WRk91twpJk
7ac1aMUsmHz36jvfnH20lRTTU3bYETV88PC6agHuq+c5Zkcgm6pQs1c5Sjs1LAei
vkcG7K9ktItXata92nPh39HG1T5aWAPXcgpILbxcuRrpzSjDowqf4iHnahi4yhJe
tg3NTzmFDaU1ETAxlaBW7kH6iKfQGbwccCVfB/ZBcES6RSDjE309zUuZUWG6Uj1S
elG48Fk5oRq7AfPonmFQ6qtpoiRqDYCUqXpXjh8HFgIqk0dm9xvnZvfAh4y292/9
XddNoeYZc1H1gc9xi57bY0WSz0QVehpeSV8BhBmhAxvQDpnl6N1eGnyeoqGBfjgm
Uh1N28GiD/E0kHMO1u+godu5mLP307lmr7jTZw1h9EMqOOU3zXl0DONNKln9Q8BJ
zC+hm68r7liIFSofN/7pqAujtQD94jUQKXq1Apnzj20gpyf1Ul8vDKuKd88NjDCr
IbjhL89g9esSWOTua+XGkt/+aShOalYVs92Z5/6Dg/nOfcdCBTWFxy4JSC7nAWNl
rQyud1f25jVXMTbmu0NGklaGWSun2FeVHALVOB3fPqu+3v6aFoxenaQuFe1DV6r0
X5v5Ytt3w4WHdd/2D6VvSoCEMZ1fdYuxcnMcKJyGOrT4LOVA/uAx4A2pqLm9EZkZ
4PdCM6w5Hd6Z9/DYX9pkEIVvMNsCDcvWmu3EHOS0EdBNMV//USY8vNYqY3FAzewg
6P3B5CGiyDeC6aAvYu4487qwuRd3GoozbihavZVuIPIdB1QKxm90YznX7CDeaH+n
5gCWvcJKC784MjUoXQuCWXbUWwWoiKStGP7FxKRb7nkJOehfrdrCQQF1lKSQ9A6z
FHutgL3ut84nuxVXe+Q//zjXGJ/UVM2oaRZenNtQT/d5ZhjX1Y/OZIfs/qTKcnCp
xjmrhGrxE3kqtEEJDqp6JGX+ZJrSB8sQUpopxgBKLhkRsQaeNo2QfEdrKUPrN7Fj
4keQTj+z6ef/mp0eQLHEpO8VTsHEJ05KkNPleo/5JSgAFJdn9XpUo2OqSjg5pVI3
8OavS2xDnqtEUIwGR/KIC/YwR3YankFvxgSGGvkijYfW26r38FnMUxje6N1NOkca
Cefzo8mvEvKYyepsTVZAe9QBuQIwrnz4sAN1Ky+F2aq+8SRGhGsNZnqCMImlObpf
B/5lpAr2xX0Tf5eTqmabvY1CVviuoRruKvbGYBx1ozwcweexehljgugUfzCQw2c2
H7YDfcZ1ACrNBvcxpxQES39NG4vB4zU3RTxo1Zq+00IddHwoqtMmea5no8AEWzXk
e38LDpehN1cRejYEfUrgncqVsierb9Vu3MY3ZodH7+1Z9Blaf1O6aEyhgCiwvZfm
OKBxpo3azmlkPkVWqQMrTmItZx590xbzunfTVHt3qE2+94O7docR63wu/TM10b5b
g1PS91slLLESs8MZBBzcP4xy0FD0ccR0Pm1ZDhd2OXABzmxYnUIK++gF9aRx9KUv
CSJjcvK4pOViuvWR9z4CL9rDPAdDM4N3wvwywE7ZM4ke0+pHRASVGOm93Oz5MwB1
ME0FgPSLo74KUGxLH33tQrtTLIsP6fmr7ukaKmRdArf562isNvJoRoHFTvGqsXut
VwNyXVz7nLMsHLAwTyEB6jELUN7nqU33IQkeA/vi7Tx+7Vo540V7j36AYHhpW4YH
6uuR1CLOH2oW7uwHm2z0N9ArkO3uHKIidTMtDES1/XCWinTbcvsd/TosQPPIEild
IMWI60sMYAtJsX0NNG1izdi6r91+oBiX4UtYsDpabt1UcekGaEyJGW1nRnlklzFC
OkMN4gMMucKW9p+BTjSR3W6fWOBEuW3rDwf1DP4pFtalln6KLOa8plSCnR+d0/ce
cIhYJ940W03jkIg6YJeJug1td5XJM1loSa086lLugZ1p5Pd+jHzTv7Z9hU9gafn+
W9zgm6uNgbCK/Q0GEs4gBYzzM4diX0yX0bMusWyeTB0DI1mDJsOnQd5ttqq5vhco
n5boR8dgGPbwmVThzpn1qQr3Mx9haBjAORcARO7AFhsbgC3cqAte3S7h15lLNgmz
i1KoNM3yGFTrj9gz1E2vTQSfSnSAAFc95XSIMd3pSL4Q017fKuvNSHNBnjv+MOdh
Fh3qdVamzsJs5ASfJLm0Yj7g+vz1o7qSTsIYUlKBS/LIdoBotNHvPSsgZJt7pnlX
t39j1NPwCjoaCsqpxO/paTzqzKK61oBGLAiqQ1xOgcg4jNZcW29mBTT1mM4J1dJx
3mcauiZ0+c2okrjlN+FgbqkWBe8q+UHRu7ZQt2jPtCFQoOStc9nRUm3sqqwmsjLj
1WC6bYrLibf6L2aL/0naosztsIdsKJCEG9ua6m9mPdAidOCrFBIwk5FYuxTaonyR
ZSLvJ+ORdipTOkIJCLFCxES31PEYm8EAwyVoX/1W6Dd1ZCWDfv2aNy1s2FP+sfNg
kF0Igm8/nHfHD5MUgkuLsBd5zgwelFOP7jR31QN1D/ZICb0E/71aYMikoV3XXzt7
6ON6DD8euDDUCwXXykKDa/jPIdcBKt0l0HEopeaHz+1/6WbM/r+GlO6enQECuK66
f4r79nY4d5gog9Lw8A/vkca0N+uhmD8Xup5cCvl2cltMYarJg53ts8f+Y7N+if9x
S5LKCjWDdHNsZkAbyqFGRoKsxNXvJIOi0wt1YfoDzKBiWoVg55nKm/i2OWY4jnb2
Sf59+n0GBjyM4zzdSH18erULAFh6lnrpcM0rUooBZt2RrSl8tbirFX9m7qejw7aU
RDwlFB79tVE6AfUoBjMTHt1PQP+L4l++vzoP+PEi3KFnUwQInNoRK5MmqUcPqDNU
u2EuRLWW0BsFJIRS9i+TeyP5KqJwnSh9y58pxJNs14cWNsAJXpU20hXdojPwmciV
zis6BCXV+bRsFLrXAQ2aVhkutZhHH/n764FGBdFVsssPI5z+HvIKrYSxmkm8y+GG
K+R1n/n8LwDyYP8SW/fkzWptM53lGrLSp00MnHOZNwPdNI3CegbTu77ZOE8UMCM3
kcclEhhlv7qQOCu5BlQuUqHGJYVrGCURcCRsrkVIZQAgXEKx0KaXtwNrOFOnKQNu
6HF63+ngCtGWZrcRVMVtnXYrQ1DqDPNIKi/eDTuJpZeEdKLSVE+5oOItEzd07PlE
DKwRbDo43L/+bd+uwObmJ/6j1JpV0nGBnDj1rgn4VTnPsj3HNxPVuiG6rgI9St3D
l7hZSOU8yXos69c4WJuYUKYiVNeC8489XSVuoIve/7iV6yOJWoeH61bLOuSTVFIX
zx1eDpUezNLiuJKaMBeQp7AlSuFXzFk5VfOcIVMwBg/uZJoj0cIE8TTZhpPqy2la
OMuXW5m8OPx8L/dOnaMbMFSNwxyEetm2KYs+vK/KIBfxN84YuQcmt74Z5Vaq44w2
g4+lzTVZBmp7dIjPVJMIwXez0/C2A91drmUn9Kewm59+urm2h2L+f4j/qaaU/86r
Abd6BkeRc9tDwQvBd3zJbQr/wzuWjMDiqzOiTEI6THT/ymiINo5HIFAMNqQK3zbo
qPDB58jSzYKDLKJSF0NQB9EdnPt85YC3oFPeQ3w0uJqsgCG3aw0tQVeplLkQ8GHe
iiMunAdX2KntAq6Un3kI0SRxqO9zBMZi1DbnWUw3GvkM48I4mTNC+NHNOoYKo70C
G/GzZl2+XjN3/Qv81DD2jTYmBHP0cd55J+g7Wy1DTz1qoeLwlfjdfMWxwLfWj7I6
q1kaKL+GEGwFZiGxZLLUBM0dbxDkmC/Sd4zT2u3Puq0kVFrBffqqktKG2Mr6bM2D
3JRE8CvtxelpXe//+8DuVkWnKzM/GiQ9x7JRfViozs+juxP2uvvgy4YEck7Yg/RU
99U5kis2TIOvmehCjSpJCQYeTdMK6P/QmkHajPYGsxMSxjKL+7HSvg7/0kR2fHgc
j3oIkNEye4BOTIHLoepAl4yiAU87J7dvFAR3QYlwoSz89vhP5idTui/+AQNbz6Om
7K4DWuy+MKUlPdpA3OYQfoff9oATmV/TwiHxUJ9vH2Svv3FpDPjdat+gaMxHZFvW
gh78gSGUriXTrLHi0E+wYfnQ3nCWbD7SLIkAIYgmafWCGtbkB33gvUQfLjnc/m2m
fN4y7E/M5tVBfJOU7rMEloPspdZJnhCZA3Vv78USEtg0lZzfjO9aBiCKb3iB7e5X
WRxrEDA4HDbRlso8zp5exgTDlj7n0RCUr1NvsJ1QSnkuZQ8uUfO6ydIIh1JGrS5y
Ot8mXF2Xnmr0zIMXrC6HfwC+ZiGAugy2J4taKg8E31Yce3XiXA5Et/IgR2Rtcfp8
1aoqOLR2fsZwtXrlGZKUdpkntt7OF7nxJXmh2CG6juOUdSdHeIu6aSRLJCCLRdHU
Zxcg7KeEvUYr9DrOIJtvjKjQ/VYiuiOWZo8BAKzVViu7tDD1HCd0XgW1cWgHLP7a
Ma3SPYQiKIJ0TebASwg3Qiz6usfkacilfZCz/vq8zRTMWUP7qVXRKq5zEJl5/d85
4CB4Mfgr0KLIe1cvstebjCCZZah4RYplLnBcygdNbELCw33vFQPCLb5Ku6PL5yFR
d8nwS3YSGjKTZI3E6sBcnrE5h9gsWYkPjfniEDN3rO2Jhb6FBquq+5h7xFJgdvW0
2UcL7Ze8Ob5nG3W9B+MnM2CpUqNt05ZmjoJf7QMyQ3XhkPCYiJn3pidfCS/9vOAQ
16+ClsDfzQkADaJoJC0kb0zUmk6QX+onSVvLALoTzS1hy3CEhj3kqf0Fuj2VY+Q1
/3oW1iiYx94LzkHVf54GHOE71+NCzBXoGX/gNCTbHP+yN3YTR668++DPXkxjLrZu
4cWS8Qe1KKRC9eIPnPltYUnh34c8pTh366Bh/jSUUBP8CeAmSdr1zW4tCTuZYQNS
EOoVgd9Qx9g218i0fdDSCfQmxNzbVxH8T+nw7o1q857baAVXPaXMd+4IP3nD43vK
Jy+xkKOk8Gse71V59JLsPw4Iwxt5wHT4+uh0b1OMqbeHVvnJizfagTztPR2rLKek
sgwXTVNfm9mWthk7X0cbFR8O1gSU7LYutqvvDYnyaLJ8AhpFWHh4rX31Q88mFijP
TsuYwnq190awOK8QSU7P9cIUb/94hJr36qNP826ZLjs7S0njULK9+cVr+Cuv5KVq
ud6gaPkUpg/f48SHSn9COoAetESdKuHnrOtUPIgB54KrDZZoOrYck4sgLajwbne4
DBnXMmhkNgfUUEWotEt80r3ZXvHXfywj/6I3EQtVZqCNlVf27taOeV1dSnPivNoZ
RbjpQbew5HKfWP7EbG0ACyPWISP6CQnle6QKh4ZibFqkxDb/d5kP4pf14sKHjEUX
HmO2spT7DsOXh/REjDkoSA99tzpQZeUgr8tDkfkna+ncn8NFUlH7SfNnloSl4oeg
F15FUJgknkXUD2NowWUdRfkcPNB1wSLP6mEhdBtlznZAJJD6TbL+9jZGeiMSYNEK
LplttH4AkGg4yahL+4Alf7A3MRPOSJcb13HnMUGtBiWp6jpv9i2Bck68xj5LVtBg
ULVxfIxJZtV7Dw5lcI8t59MkflrJL31kBSKIYoUoRaAHmMeGG4JpVKZYmPyA01o4
5rqRT0Tn5xf7gQTDstAbtIX5K7GpNuXmFVfLeOaSwV4RW2imc165gSFQKFnXPGZx
q48LdL2kc+DPIXZRCQ+77NfREeduASQ1UGMZd6E6M5PK4JBb4xEAfc6N4jEGpNql
Zu3IBjMHPYtJz0Qio7BzDrG+Sv6A0kYdOeyj6A3qG38i73Dwj7MEhf7QSZrs3s8g
cY7O1VKuOCwGja6Q2QidCt3biBbs57ezXok/EITX4UhII3841YpQ40Iv01pCtNJl
dB6RToFzTy9o2pYhhrJiiAxuOPOB/sd7gqkHBgYiSqP0SxMX4V8cqPhUwr3/djui
IiJl2a+fXMxJ5fRu7j5ZriGSUkycRR2aW10/w7GsZ8Gk61Bci7XjUnxIt1yIC7aN
Yv63AYBb4xD6e69nNqpO3muZ0phbsOeXCG9jxkSlvQ1pVCPAwN3W/QSIdaNL11jJ
fJhWePx2h7ut+eKnpn+p5+XFO8yN79DxFzehi2zLQXE2t3bwomPPrtqQQwSDjVnK
2oAEJ8JZL8FTntYi+V+FrKgAQ0DFeqoWc5rFYxAPFcBJzQQgLvKmDnNgeJqYBeKj
7gbD7IBtYh+iFEeQN7ovx2WgrVuHaCifUk2UzZNfxNpDsVT23KL7uiXqouGLipo8
uVPwaOJL5PhQmbNc98AgRqnYusQ6ZzCeHoOUOKtQKp/PLLxny8lI+U+YHcRmqG6V
m53AhldBawWtwtOY5hSNH/IXDW1gTjozUrU51vxWaRQmaIJ96SvuhXlgXwJ1uOh2
Hp/Z+c8o2zM1uK4PEcHVmi9BnRy3PyELOGDrVUwDI2hTDZ1/ilqwPH3ilRPwF/SB
g6h1XkgpHnbbROct+pRcFeZyglBRwVUVreZTbTVY8pv0RnnpIUjH3cmrka3wZRa2
oOm656vMa+b6usUcpoZ64enRXMKmRqOMHtS5GS4RE1hgwR+/ImXt1kSUaCES4YJn
OvgSRDGUVGvkekGjYZcmGv6Fgesu7sdFbYYmfSzEnxmVDZnuXG9ePkMJ+iFpPO6a
UvP2FR4ACXEtJd1ZzMcQvjN2CaJvxFvr5Yf/HFulTlQ8SW7mBBNt4ZJxcvOAaovh
5SvOrbIsaM8snhDm9u+dHMYwbvPd9ZopYlJNSYazjfwOzdLI82mMXxHAhidjs88G
8GiCDfhm+uA0nk7i12XgNRqegFwZh9fTRkg48i+88ALJdjU1mCGKEZ0OUPcZBsnz
zkRoBOGzDur1UNh22fQTc4MNFadsO9XKCX78fqrA2O8AUAL/b7SnecFLlV8RhfFA
RiS8KdVoZBGuGvK/R4pkKv1hTrnIqy2zxx4ZeQFjX/PB3aFwDo6FG2Uac3oryh1r
tsFStWiI8uePMuhv30+EE2l3GWxwv2Ti2MfmOIezHsfSEB2q9qhEkAAnvg+IFcQO
chr33jED0nUprEAr8KRRWMvW93kK+9wXbAsA3C9800eZsZbDAHXycouL+RxzM5Cn
zDf1/9IknGoU9jLoE+/10TO5dBwKtqJQv/eMFs5WDeRceNjdmQbpI+ffl8/JWBGS
toSxHU8rORKULDP9Aov8xGXNoDsXbOGBJQ9+zgUYYL3Sn62g6U10p3215zPYwtnA
OMQ5SNPa9PD5Kudw2x6GLAWkxrXV2rPUiU+isvXjeMqjKZgBIgFXdUZOEBYRiU/o
aqMD1ixhsNOc+hmXW96w6YoqBczWj5mBNR58cYR0oq5pYVjGmlC72C/Y6HW0gIpX
LFDNUZubOgLUhIg0PbypBxwlefXCC2Y2xP8bMbHz0t3b1S5o8yqw8R172NfxAzgT
ioeiKrl2P7f5X+sLBXfsmF0aAlAKLEPiKxkOqhyl81DINC/lcxZx1kPK0xeDtG1H
nLt04vgJjgEypNyGI2vB40tiaHijpWzvsB0e74DEq5vOH4bLMYg/WDdpIHI7ig92
mkPr+byGr/E0uAn8gFvY2gbnJke1mCt6EDW6CVb22eD6pLAq1Lzunb1fg8WsH+1M
HhcMuG9vY2mOdeOs2A0iktDWWOj3JMGPMuz3hL9hX+VUUgKfbBmaJCKnXRfka/Bq
0M1z4OdpIc8FvOc5wqEYyuFrBeD7v6/nuf4Oakx+J5zWD03dDso4NUUcSGCVix/i
wjD2oJO9oRJa4rfWvwGOaAQ9agniygc/oAOhQuiFMl9IPWcitMwe5VmoC0kWhQLN
BTfJZnrDXS2Ewp62PLNxQB2qvg3afTVgBsZI/iUl4CLdzyQY4JFoBBih6OYbHhLd
iA4NRrtbGxb2zzkHMQqWA2LdVLLEqaEifUDyj6O3G6U8UKjBme5+0mYLIxGFsTte
7jeLeJ+U9wS4Mgwi/GPbdzxIh+gM0PFXx+p67075hnUye3apH2370izSBZx+2lWO
fvtBLvKw/1NMZxdYOLLlK2chZvh0OoA3X9k4gKRo+8xoQdl8pMsMglBoC1nFkNBt
WErmGug45+SVVdcM/JtmTdvAVHolKDsQREfVcSYm9KZsLGp3LjBaTq6Lj5+NSUyM
Ob77mjvtMmxLxtrCFPIJIzTFRCo0aIFLgjC4hwkHSseZxIp/UnH1JUarK4Jn6VVA
opKfjxHhLnLlvckzeeJB2X06EIdrG5KTlUe7ccPc8HqCzT+FJI6ozUbEMmVkzkk1
dy+NqAEDvz4zFplk8Dp8uvzre377JhRPGlitsfRcgZscOaeQGJkOO/M7aOPS2tWw
DyKXN8x4atu66QHAWnxAbHrMzPYZjpN423JhQ9cWPf8/yPnEJ8LZeXQ1giO6oIXM
Hagz9pmabTN2P7FYUERidAyWTJpxhOa72rZeKJq5gAen79W8UNABD6CYhS3Bbw2G
VWrrq3E2+3BW5+k421Ua+P85ug7HnU5mrTzn2vimxtJjoz1kpjU86UB5P6NXXC3j
vSUknQLBn5Ty6NbdrbZTAZJk9JkYf9sigl4ShFn9GeIOKcgK4KkkQvrjQsBik8du
PV+BTPEaiSNuVVBX2kQMCmuXxtGRCnUcGJni8Jg27DxZbWmvC3dj8jVjocc09Tg4
9NIunRHmMWOhIRYnRJi8nP/8OjDG8ShMjyDg7qj4hUfxV98cg2GRjsm/GehnIJjN
YTLcfuQPTC3I5mVgCBY/FnMXKc/8fPO1o5Pvdy+iotvd8BEJhimbDLoaEQWS9LgI
EX4LY0AgChQhT3uTeD3QL2Wh+pywdsraPzdeQpUdXCkXco98sAHPgUdbTIbUgT/T
jQXrzmtsrOSSsumlvxt6xZ3AlZv1wnQmA7ywtGV/IDL2mU/mG2fg1ddnQq7uiMl5
BJbPeB/Aghldv3UDH2UnudwqKB9k09ow0KY/iVsdrZhh31NKdTcxYWxAoiS+ThXf
Mxd6WWB49f/av9av86Qv5e1OngzkOREg0UIGXrju8HdiFn8SVDdby2JiN5Q1ZHbl
jpDA2imzErS0ea+PR5IyDH7tiERtVajLmDNGVSkWFcvj/EV21BUbUd1inQP9Ce7e
A92k474KQrZtPXf+o1I/QOLOcwg7Qyi9BmNIr9/y8p2SzmEsVss0Leses8Cy5lbz
L1VXmiMT8+ll5dCHaIdae7hiLc44XlPkOReEMkEFJUazyc9A1KOhrAp/W/xhfr3z
FMCNPXZdIoyGOMbOu993pbEQfszwvApRiHCf2VPumHOeaSneC3N6clr7yXN60F3R
7fCkVfJ2vvO5yRb2x/eg/cxRHDZGTmvoBLBXr+6Y1HI6Ni0VzW6PKdqTUHPrEtiO
HL0Zrty3nqC37Ak3xt60j5DTJ6obX8NVBL4b0MiiS3YvAeLnwK6bacnCiSXorS/N
T2hRnzsHt8TQYK4lqLpEWknDyTXZkyoF5TIPKwiqVq0uhQVydsFAnuce/YtLXIsM
WaQ26velztv+rtq21IOXPrT956ycm+3aHDIuAQM/CSt3nm66a0xHP8Dc8wGih3ML
8F4xtTwSO3f5q1cer4zKr0/A3lC74x8iDumGq2WMbt5XdBlBgg9xM0IvnLqnFb3n
IKdsgzUGr+utOeygixZqpnxQUz0Robz83oy42pejwT2omu1hzXRWLFVg0vKPXINY
pVLvxNejiMI/yvkD1xBkvneU4Djmiy26w6mFG9gerU5xcJ4BLLXo69zHGI3he47h
VYQ6YhszjC1TQVjcuJc37BYrQxXez9yKVCHOuNF7PhtCI0SrBJ5hQsNDuU2iNaXh
rRQMxC6LzMXF/GsFLjrIClXOHJAPRlopDzNsfBFNv9q7bItp5TST+LX2sq48D/r6
XPD3CmSjOv1iXg+8BUwNc97i4/M26xzgEtNw5RNZv1ubNNqBIdPBwJQ6LD+/te0Y
Zo2d6wStVVdqpvD59ulbl1vxol9JZGIWGGGajRTGlk/JTb7Nmy16Z0or2hGIpsn2
yHDc6GzQTkkDR0di9uAmrcRPz1j8/OyK7LK3KcupnaYh3qMM1VnXSJ/+0JHpCgQf
P9TcCx9sCND4iyJkuCZn4hYr3ENcjgTN17xHOUnKFLXQef01R6Jiz5co6hQXPGXL
tSCLe6d4o+GaAfKzgQYKDnabZ/6UotaJHS/XT6/MX9QRFFQ0btvg1nYxRUlCRdcO
/7WqpyA0lNsM95Pv27xhREac5r0lmrLarRcD/3FA69ou5G6u1p3nvV+FSuzpb27I
Pn3qpYBUi8R6dpiEqGy9gtmO+BWNqPtUlpG58OfBvrnAaeeZt+FoT3Bpe+Gc23g+
n1TRoUclX0AN9EA5L935SxGEnM7YwR/tZzjfSJMsNLOxe/IZwAu7RAcnMiUDoAC+
DV/SAktA1EnhOdwpip0VDldaTj0ZNhNAdLGvwsayoguxPazi6Cw1QmeeK3u5vxZ5
JI4EKLjLPpONItKyG3bi5vLk9SEMVDMDGjyeJzdbYS3CWPeHUZ3gOqMksMpHUjCN
Yqab+jBeflX14iD6w0UA25EeteiJAQBH3Zc//Z1Xr5wMN0gPf1QGhoctKaIyS5Fg
/qEQoSQoaClxg2+FGOe+QXXx2Np+NE4xDBY1szfm/8IZapgX8fWW6QYFaNa+LCr9
lJsjbXF020Jy6ivU49VMA10ybKI0TtVfa3R3ZujNptDU1ylWu+b9n4XdDJ0SUqq6
gVWiHpljguXc4Ouv6dM5KB/n8FNzfDixyuMIZFsFr351M7jHLdL5qRY2xE9+QbDS
WJTgyreREfmy+/cShlPscb2RZIpEOJ6xE6i4dHkx3oiBsOigFaL3wF63fvtUUZ/X
Jrcb/t628ehalqRMRxSEnTpCBdTEaumJ08umKNwtZE9s2oIW/zFfHe5F8dYGpfFY
smCUuB3HA1eMKlm4hhifKXb5cxJO5jVdXOVJNTLIUyElehyOaVKsFDQFUf1q6hiS
4CIecW65QUnUmzs1dUVE6srrQCNXOQoMVLuWKFpX4XOT+tCDQ1n+KrM9CJs7PHgq
1oFrXTVnuxdIOpn25M3nGZD9lWwjONPUYiWzg+Td9s/CqHbMwim2yAaoLKIlv2UR
b1Io2ksMloXHjmcAGbZ+FJ8+BYIJIhzv9VysuE50A120bORd9H6wVkrh27/k3wfy
mifeJPKm2mToPgs5Rt0ZAsOGJ4VsY7kGrxVV+j1rLDKxR8k6v5Wnym56fD8gg/MN
niQYrXvfOH+C5qdzArT5lNBYH4aTvq5ZyDjCuECsfAkLItIK8ykMOXpAFgMYYgn7
I3Jrrpxyh4fLCB+v6cvf/6/9G6rb2szKXy4rfC8EbnZq4buvS7hnVtmZ74J9q/Pr
NyAI3WIH7drhE5M4JuxmOKxWijZ3YdoXMuMfZcMTzK1+/e7BGl10CL/ksGuC82vW
yLYpA5GakpDkoVsEDoKu2bb3cvYkQB2BSBkonow1RUQLUNE2mifkRcQcaYf877u1
ARbrTh7dgomwT+ZQyzEWU+R6hLTh6y39WFhiyTZF/d1inZinOwcZskBgY9s94i+u
f/o1rsg1xqdT/RUej41PrmnXF2h1sQjaoXZ+MOUKl8w8DZUldICyP/RuXUFtJD77
0Wjj1IGl1gJfM/36KBuPjQjvzQxSF/uIBr/8dIkNyEbegwU+qiiUcc1zWzS0Rb/c
PmBC2nvk6LNxSn6KPgQxVFMmZxn9x0OgOmHjbh7wznl1BGEH7mzbPWNEV9o169vb
B7E76NVLWtkOHowWC4bCF7Q+/jv4bRbql/1f99LEs3SEvLX11WJIQ8oIeYpYfApc
C7g1xDBOVgOidsfMp/8j8ZSB4acO1Obigwkd+QwUXuzGy//dRLtPNpcZq1zAGawT
6033g3+rM85hyZzSY9yiPSY3XbOYrOCbWDjDimY1HoV/SS1Woe7mAi1GQx2cQLox
FHeqmVsjoPEfzbunyXCC2Mt6UrIhvfeLPP7fLUw3OY4jW7wD74TrJbcUDQq5IPc2
uc7kvsmn26EbjeJVaUR1ifuCl8NyuEi2Mk42qV09CrFBWOdut88lwZ68dPlMr9Uo
sFgs2eEeAt1799FH/rEhDJ2L/37TGtAZp7ioCVy3u6t0An/ripMs720Liwgbmy8J
I05MaEVqLxANVwxCp6XviAfYxFtBMH7l1FM1CbLbI9QEzo+Dma18aV1laGDmwzlD
0588v4m9zlef/ffLJ0VmT6d2N3j/eFXlUO8kBpksPo10/ovz66OfRmQe8oqIqcKi
DQ6pKhQxNvGCDfVdbJbhZl0rTTLIPp1kJyfeavADxFT+OvHh8K9hydISK6bbyLpZ
zVaEk2M4bAqwEDwURATHbH5Sla4lOCNLPHgBtQoDvS1z89yoqyQUEKGAb3k1AbyA
XhtS4scDtwZNxTXivYooc49JAevhiLq2zhc7G65bdmfn1Z8n1Caij/wlV2p1UW1Z
YjLwI5kK5WFrexj6EW5vN8BCKne0ImBq3M7iUP/p4Tz+AQvT6Z4Jxsx8GuafKWPN
UW/xDLwQ7mUtmjMsbNpxKPN7wQ+TEB2LqU4X2zvYzF/ACwKen+hK6Izg4Rn/H3kn
8NDPyDLloH/hH/3X8geEAoQTv7LsY/1oRaVJuUt6uPs0Zhvq9WU5CXHQRK6n/VaY
qCJhh8spnOqTWNWWP2LzIY7NLo/r8sEQRvb+s2h88NtuS8oDR7UHi6n916Rp3o4T
oNTKkqJCgCZdp9Jm917vpqOLZZaG7dAy46g84IlE3kJsOV9a3QSiYATsEJVPALwT
xylcaVGnuxa7NZyRyeGrkLEtxSwquWfq17I2ZG27npqUlgQvlypxKz924P/jMlPQ
mzHMxmMadz9/N4Ds/zmYV7CBNV9S7qk6bTZSRcFmMxnRPCBIdOFDeXvtGa1E/Sjj
3e8tU30m7h/xAc1A1S0Zt0V5bj7bDVSDdATY9jzIf6YTLl8YQOaaz2Sx2uCSl0NM
nXvMgNhYsjIAyogkIKYm30FlUu/k1whgCENyC+IyPsLFhfDX0SsvBzUR070QlJMo
edw+t/kNQPZ4Xa/3OfF66CX7zjZE7ax/Bm+bGmAlX5sMmeQJQsWVyFNDsOzggGfB
Y8Tt89Xi6LsUBaVCmfV3jInj5z3iqt/Z9OMZdBbQUX1PEMm/vQXTuft/FfVrErMw
3+eypB71zzf2LVspdVPBBL0+KMgL6pQ6uoQkfMjdtGQ0tTJniLJEfmI5Rkd/jwj1
lsV+UK0TniUD9ERJstYRoFATHIgbAF6vX/CgY0FRRGR+5IDXswcg+S/X9WG5712G
t12maNptFIbMdL4xwz8taseyPq+O557xR7jGyWNtWEzZKiORK2VdGU3q33nEHnFS
5hNw21qMOZRq5BuH8kcM4l+8JqcDIvYgoeVDgZyKHQr1LVmBF50w3lNS8Sd2qqAr
ktoT7xwQpkQHgVUU2U7zYo1pJH4eHgz65c1yNi1KbntGsuwCT+mQQRCJNx+3d6Sp
BGppIQNT2liTgGyhFAUGSz56cwXhB6AHEbC4Cp9mODhjxsTJjv+NG4i0ZSb3B21G
jddzgACc1fN8/F3Z2uKl4wnsModhUYD3bCLCzUiqRgsnwwItbJC9jzRwciVqVxRS
bhUI2n7DFkACjzjmSJc81oFPsfgqJR4CcGl6lFoE08LmNnXms/LTcL5pq34Ra+Pq
FKbuMEOsmbnZvv2zb+SM2Kcv74OpnFvrDkhn9VI522n3zkkSJcknAs411S/DzVN1
ZvWqju7HuTRWUa4evy0ARDRcqe5WxnC9I0w3LlW/GS0NB0EjP5SJz6s4WWTCMu14
JP+sokIUWbAXdORksCVVOQD6y8Md7y6fop13awnuUv3qG1A5ut3gY+1MCIOdyW/X
Sox7nLclZHhADzIAlb8nOf7AO+PFeAFy14vEU1PJarUHFhduu0aGWP228pcX85Uf
JNQsDYHO7HN99CIY9oEYTnoNLJY8SKvhb/8FdPYvGMSDfld8DTx+482ODxbkUOs0
C8fwYBq8xKsTxCEk5hlETlGqxQz46G46DM0Q2vCTuqpryJK0CkWu6GEnWlVhtY/X
KvSO8ZLJvUDB2QCMiPKirUsUoh3YCHO08W7hJkpzlMjOGfwd9pp/Z1Xa/zaOOa5F
LckEBRFmiSBVARkg/RN42DjjSyhM/uAczh7iHeFT7HKMN0ZvGzfoKFueUQNfgl0W
0iFblGNflq0pvuOE3bsghzNZDkcpGZL0dHugrwkYabny6QWpuqkM2IKPzR1T31eU
uYudq5w7V9Bue6dnTIYo6/4zn8pfJYPCBQ5/GOKFjpLuIpyEQl7DLqrF8VJapkav
Yqn1GfKTBhkojrVjYaIObSUVrfQO5Hh1YJkAOxeyRsz2uATIUyEW4LGgHJQX8pdK
yUgSpbHBbjqXKfGPdhzI6pPyQ1T1tzCoIBr3HVGgvrLv203VHdEzBTtreJj83nQK
8I4JBbeiyi6rH9CvmOMaaCa2R1YsH33lwy6DZcrNWKb0jKlKo4gpVlBA6JPC68hX
s+3BaqF7OQRMwdoJV5m/ehMCbVWBu0f4nJCZUMoDnEpe+C4GfjLtnac2bl+hdu2+
EpBxY0mm+ZCsY1UsfViwoUatI46F9JFjumXMdIp98hMy7jBT4AuFNy2ZbLqc+qK5
Y33LZqyXyHO+lv5VLbHKK7lMLvOIbviwcnvL8wr3wrWFRhO/bMluKxUYlteqI2wO
LEZTaXj2xshXuitX0aWRoUEDV2qoKj197sd9aDUxGQ+p7cCC7cBYWkGWwbUq8OjJ
yWryOughsZ8nU+f05WydLL4ty4ZUW1p76lBxoHb+OsBlrd5BB590t5GgfAmpstGa
SoAD6q1QkS59eVQ5NWiZnrFRpaf1nsKMN2niVGoOaRd9p+2TXOQYFZrSHT2ZnZiw
LG+b8b0EgXU7YIg9AA30wZt0tyD3SplDw11yBZyExxlwmJ2KfYi8lb1/qKoS1v6e
nrc0qgcuj9FL1DByiry6ORNjV0Dvom51jLfcAQyVfOTV9R9o9yFcBxQOW/5LUj79
5qqgBARuOZ5/drcbd4ClFmaLKctp1rjUoOfFdW+7Ieu98Fru23B1Q9pUaseS65mf
fDTDe8uYxqDPatuhbHbJGy98RY3oM2bKOx9Ypb35BCuI3HxLffUceAvwrmYQhLYn
YQGw6mOHHEypZKhq08TbtJwyIIQn3zFpCPpJmxEZDznXlQd57v6/MZ5BavjjuekP
xx8Mqf1eFjTCwDwxgPFxKjE6SdLE+jVqeUXxI+7qdAKK2M8DI/M1t/ZuMFtwWNz9
zowxS4eNgHLtdnzIW3kol15sbdm/4CxelFQoyp6D5o4wgHIZUGuRWXEkA0ylDVkU
+My1U92DLbnu8RY2ojyuddwwOPN9gdXPQ/8peVSuNn2+QPJZT51HBAjMnxanR+91
+hiKTAcTS3vfNaDZ/70zhx35ZreBvHDjORZmOlHbimV1O8Wp7B2raaQ+pYtNABjK
vyv8HqyHrAgIBvUT5BTccKavT2rfznKV1gjbimNzcW/mmLQ9HnCylCf+8A+fnlMI
2ZLt0X/x8AQPmZSHUhJihOQj8LdWCp+DJ9igguCHVja038IRdzREg7FYiuu2tORA
6aHBFcX5BkPYoaeZu9UNJwHCJ8K4QmnrpVmaPL+EeTrHfI/GMM77allQ0+w9N18p
3Kp6TwiLYXRejsCVbPOv3HYZPC26ndx5ois0NXoP2YSF1o7jQeymAVg8udfjK4Yj
vnIuIwzaSMH0OPdkICRaDGegM4cJHNi7seT125O5HE5r3EoDVC/kuEOrGVb7ivM7
XOSvEaUm7c8B5gU6hJtcU9schn6MMtgLMNKx6cdaNWG614CXQQvdoq7D/0NR+3aV
GJWYoMB+qG2nnbPLPGLc+6JLVrO9EA4KkE+3WWUX+gaKyr/Nn/Tavc6mkQu2QGil
YlYksTHwzVt0XMiT9JVH6NM0k9U5KD9PHm5GOB6+5ItCZXCcFLUon+LXAKRHuX7z
WykZnOt+P0nbFr2WI0t33DpGkqWpabCgPrHgUyNXB1HrWJv2KQ+IXX5a83zTln/d
5UBJjhi+RqOj1UmNtBOfIWpuAE7dPMnu+oPLholkxucaK72GTmxW7nNLIiH/ohp+
e/OUZPSIi83ikJB8LwfZv4LlCwJ81CYPZe7RFdvPDx1V+295oskH4K704tiUt01C
/NUGmOnscrI1C6X2E+FomI1vlzjCDhIws/w/kLjYU1AHYcQ8Ji7WJ0SHTLQK1m2f
vg/1P3JPrTt3UsYFTczou+ZCvDRvyS24l9aCxyruRTu1MXrtVUoFPB643K4a6bBx
7m+lQWg+sFkC8SQ1QGDOsBarCiWBPJN9pe7+/pe4HwLy4WIXi/MOK8uz0awNG9WD
TVRNlselILoqnTHmZeZEOREGI61vSksHyGydoWw4qHKt9UBRKQl4yp0vusgy6/5l
xomgHDfk43sd1O5ZtrV/czNHM0y5LAxDM9YEcmJzHdulHKYdxJvWboi96mxnHU9+
viMIY9ydLu7H88wdhwuHI5HDebhAf3tE3SK+dgpLFyMTpL5ebI3f5b+fws8YxuoK
HQ+yoVueIOuiKQEk7fBy9/mmEz9Jr5RtMLSTiBKGk4d7KDEQ0zAsCm1RuY3fajWa
JW00Vj8g3O0TjiiMUrddlRX6g1Nx8/Wj7iwn+YdXYVkNEA1Bcgr6wkoCbpDoTwN1
kJP0KijluDHv8hbIlWbzdLXSMqOQFuHzuBQLjNFZywM1ntJwBIR2SGBunpZaWUa5
LU6yitF5jdVwNBlP5thfo8V5CDgcdemX5BoDKg2yMmbN9qV0A9piB8kG+9BxdD6P
qr/gI+i1IXREaRlmdsFtTtZIuiYzUmaqNAQnsRzc0pwjhVesj0qTq9aP/M0rdHV2
R/CBsy15ZxbcgbYcjfvGZWTNYIQ0Ziuw5ArahT4nL7Oi0Q2WB0P2DctiArh6dtvP
GI2fiISlbw/KuaK2f7JTmVMdVHcXY63hOp7tv8dscK7AvFgwIKdDOHXVJyppkw2K
fYRMzfXBKReiuuR+aw5UP1+EIjHGiN7q3yu4LofU59aSvYg3YL39slsQVc+WSgUK
FGJWAIxBUTAGLRfAzSpmxIG6VgOcJCyGJvjW3ahIIZ1WXQ8Fks/5ZLSdQ4oV0kLe
2J+2br2SUNLOHn5SZ+HJjY9n2iIRkykc0/SSwCOfxq4cmyvTTd32BExY45h8hL3Z
Z4LdYIbdzEYLn2ocMWYqQD8n9sUTnj8zDzoyGWhvJq8uZMoQ6arAASJ6MiQM92DZ
rjhtoOJgzCOVoZZC6DsnkSQ/8M/lhivwCiDX5pvP4/5o+aHgX9irnkn0dddC8qm9
TVLureNcKNtdGDYtTAORzyhQ+Y3oEJdK9Ms2DUGZUqKGUtfWL8LreyQyhz2d8a/v
gFEyGEP4g0CGADDELwQgOYMK2+QPBjIJWpKCLASW2M2Ounao/xC4U7CaejvQX29j
gZVv0vvEOT2GfrFNEgk4CwHs9SM1OS/7ZdVKoc4BkOi9ICMiUnpbw8s+b0fGJKNr
Hwr10qq0MMEOSLE5JPb+HTuEa7xycVjjJwE7L0djmst+jykNesGamMUIjBmjJoFi
86ycwqWjrCns+Wa0CIXjtIKJKmGFQX4xt8IkLwJvawhxuGoyEjzkXZZ227YjsluJ
zdYLMoU8Hq+N9aS1tsn/XWb3ZnLpyA/x8tvonzEjpUCiBjca4KitGgwnCn84lVMT
omFdQU1CTIEc0b1mtaGF0valKR/hgjBVEUbYuLrBs6ei0TWNqQQNWgH4V8h9VTUP
UpoIY8XHNzEhPj34blCBjkt6TKoe42gm7lOl5JB8eBnUdmx8eTCwFRaWIhRb4rAP
QdQYX2vgljHG3UwnH0jVV9EWEy4/vmXXJlD1vGuIZH76TEHNBtaLeN11XehQHCqZ
+E0hS+VD8qMPvFJM+pNaaKGJOdh5z4jCueWqtun1aJFS8M3L0cYnPHal7PVTtQ+R
ZqU5QmqSwiVDVkOcZOse9C+RP3A5sh0FPzKsUPxbU4OXIYR07b3my2XKH6xyBmNj
LoirIVMIURS18UTe0hnPgq1K9isD0/gL1zvRIknDwXpxJ9yxUQpuX3YF81TDy1Fn
5PBKGHytAzqZwQ/gjigvOv837L9wBoubN8dUl4DVKV7REUpXiF3Q3Mb3HiEsq0Fw
tTh+ynt1wcXm+/NJ2Mz1kJ01Tq9eZJpXpC5Cw5zSmj3Qu5al5VcxkG5largVr6JG
emH/IWjZsp8nj2nedJFi3eA7B2+TQExLjwGJfsU+qrEpaDRjgVFjhCq9JjakdfHQ
AD4kfNicj1HsjkRwgiQXFbjlCfgcCY8Nr8E0sJxE17XIRV/BUiB5m8Fhq0jYcHP1
75NjZ1Om3BQO9IEtv+jv4L91wPOvq0+wGRtNXJyfPA8RnBLDP54I0uzWvWwiG1hI
mvvPd3Ga8h2R8S4Jw92/W5p7h2mHePN58KCtA+icZVzvaHeazlK+0D5JKiAcESy4
CH1I3bG2eIt/MvRjC9tHBqPK3mV/FvSZbW586W2ztBn2qZBLFSD+DazQh9/AZylE
fDz8Y6OodssyViLGHG9GryVIF4biCZuQ+YeUoj7xK5m0Ta15ao8gGGXfpjU9VZ+v
AMzWwlcBJyOxtBCGSrCGGuIlIWQTBy68rFJlqY1or/09A2k5uglhSq3WObzTeB3S
lB+R8KURtb78xyhe0z6U3QDWpO2kjjCGcbJqNyKIlRiHLMUD9c/OobyqI0PeyJOC
iMgYsrKHYxpS3RS47Z0rt1ctFTHLjvFP1T3wuGBMLboo9BkS6KkJNTzOhTBeSQqF
jDMoSPAFLX+ZTnw6xfr2NEXe8Ca3RqdQym0N2xZkMLarEvTmGoIIoUsx/8rJ7NmD
1FUaqEhe1Vg/Z3psrtGoDw8UyBUUsSv+wSMEdS0xoHdqtyLx4KQQScGbeSjWJ5Kz
lXtUhfR17BcfBNOlh4kDRHpYsi6D1Q7s6q0l4Ugj+ttjDkfvYFeIbjTEG6cOuEom
KeXOCdnkq/7kB73AQ+FZeRt7tN38+VByczbN+TexdWd3bsGa1Ak+Q5pB1ZMo5SC5
pIz4xJg+3I7mvFCTS55EoC+KNyz3Lkgs3lVQIzPTuvMAvd+YhU+mg6888p9T4x9h
dAxh69o/cp0rgZCjmvTyGf2fyNp3g6uVEdHLoF6n3tCarU7XHpAyOGba3v4xA8pn
LOOcw2hpdwLATNjQURzTC0IuLmiEBH/yb0qglNtbLT3fyvM3rP28lh3wFu9dCvFP
tHK/KRD5wHjQoc2WgALhWiBuQrD2KJ28lnLWjS116+aHYuKfPLPKTMkP/S1B2W9A
ym6j1pDJIO+X2hCeAMhl57XLLPuV8pEW29waD7tQ9IWO5ICEHgE96BVzAAIyTAVj
ySFnN4uyvWtalD4Ecqr5ZtYsYm946ztauMUIh6XM0Q6j2EL7rxPO63X8RxcJnh3L
wrvNOha1Nv/DPICQn9bTtbsloGpN6Oi1h70yXY3MQev1PC/z5l8wrwHfUfr5TBhi
xGX644a9EaxG2OpJyrL03jSV5V6KDqvVuKPl3cRSnuIQw5m5LOMk0XVvRVZE1bA7
TSobL4F79+VutvdZg4PIUzJm5+akMHrJiZdYJoK5mYmsb2/+V7JEUDb1Um4EoZMJ
L4ouyBmGkJmd1HaWl/ANZCWci63bAPyjjBvOW1qo5G1XhsIw9VfMuPfzoSVvf8mv
ow80GW95FXwJoNANYCxdvkw3KPkv666Xqjh/O+Dk5K7tNn1y0RivOD8IIeydTaom
IIWCJX3cIAY3gPRFNr1adnaO4GQ6zz7GC8fIuqt+tjHV8i1oRWgWCSR+oCyaitiC
vmBswHWXy2ftK8kSr/mQ+6aKT0Hk8Hv3mwU0wicHFpMbfFWK0iS25MrPKHx4gYrM
AC5zDsBV2dpbZlGx0cy9tjW1NEEa5ILkbBkUGsk/TYXSxZcPqVgrgyHWNcjxbO9e
QL6zz7+v6OMrNCGCDcU4bYQ0P+SrAShdCtUQynkgi5363r1U/sEBMjG7ok1qLz+b
uYqr8ZMbzqoRswYi+Fse9U9tT51/MgD5Omj0XB36N1YAeK9n/YgxkBgd9AlttzF5
VaOzMC7uxiWPjy7n2bAFq2b63mFV1ZcE9UakzDvIFBH+zgPxvzypQYFgg+K++1fQ
zUA90t3UM18m1IVpX8RDdWAem1j40vMGiIFm0EoVEefb3owCjA0YBgng0/ymcwu5
qdn/XBOGwcF1YdvnAHOohwgwJkroNlTDWCMpg8SSgo8VtrqdoYiUdC4DLxzHv61P
BOjR6duI+LW/a9w6KVGww9Mb0sJuLK4vXRhE4T+mt799kciMhcje3GTNOiE9lBA1
zBnwfUBisYdzj3XVsIMFs7EeDvRbsFAkDuMcAlkthpM64x/QEOvMUIM+pocnAn0Z
kafKTg5rUEWd95pog9VeE9Oeh8LK197QLZmFZ5mjOeJeBswVmQuYcVNRH5EpmEnv
8n0SPhv4CubbMNgQkndqY4hH777DsedZmmKGlvAdAxfCotpJLxr6QgMtFQHnPLNF
J9TNYqGOewTvF32jlrmevmSxWvXHiKsloKvXU2r6sO29fmv3DDbE+3bPjVW+zuTO
sGCPU3qPzL+5Q0cN2r50Rj3ntVnirt8sVLs96kin03C9d7IbUHUCNn7LfTdD2uvp
RbbSQTtrUri8bk+YvguOrcFOOyN7M208AYFPcKO3LHYOYy9+o8BspQucRQVrfAET
gxuEhHhZQCTgBoDZT3dfxMim/qcBFxSSNzbMu3R1VikGTmSAqE/PGA9QQu+go4qg
NDfKJpt226LgsJ2mf0NgB7J/w4cA5/a46Rx+SJLA2ICtMcYUt4/agLkUcI3qYX7S
4yp42JXPSB7bW2X0tXLoHrcDJn71df/liQYoTsSLsydih3eChoXoATfxSGrImR6i
AZBfnNRUpOr4rMAoC7ASHPH5eTK2qkXNDnIV877EaYvfr/3BfPu1rZ4JCrS8q+Nm
R3CVYS38dbb7xUHL99ffoz0nz3H/y7QRkAbxYW18OB3jbnh8mU+dRimLVvAokxVQ
tIj0uYb4YBt6vAnJjhcKS5n0uKUeLbRS4ejOWKQqV0QRTX/3lvD+LRr1mHwnCql6
jA/WtMCYB4WfoQe9I7TDxRqpxlLfCa22Bd3M7/HLUAmgUcSfu+O/GA7y/PE9CkJJ
bmXR1lpUCaGk0UGNfHHH7oS7joGLGqh7CB8kP1JTP7rp8PsY6dA0YiVYcaq4E3dE
8SbLXB1UVB24Wx+TGV/SuImzoDI+Z+6OjuDzH+FW/eOCHNLJP7vnx8VoNCZAxYyI
32cOe5Hy2VsuK3TkDXbhLhg5Dchk6t1qkBNmS8j6UuLApCEqVoz3XDyKad0seeGv
gDKvTCWxe7kdBZccbw2hTNvmo+73Q3Wu3ANtJTpdInkrRFpRPlxsqgAypxjWgzuM
B5BfTvqDm4D+dktUtFVNJVr9j1oB2JIIGWNDGXPu0lZHRMI5/C28cxfehVs29Hsj
BaCK3FNB0/pjc5fkXS/t+Q2URQaArHVhXUKxDGF5A2j6/X5CjuPthkMe5orzKRFs
2zwX+7eRqemUW6zCkWAgZrpiv1OnMmlmCWgOWYOkMgyH9INgXZTsxGKFhucly3k7
1XZMbo53lHbk717iCHJL3+QO/lmsQeKuoxzMvMm/FJzJOvvIb9s7scoww4JPUrxg
utdxlUquQN8FW0RZRRS0+E+91Kh8YkcI59IexHuAZmPG7hOu2PRr3aDQMM4JsAIa
GFFlnhOBh22z+AfIGnfyLLm6rwaZZqw8rN0cR35N0WqoPCAGniVHGdJ5IO+qpjBp
p7l6GUbNPZm07uWwlxEh8iI3k00u0vuekGQ2al69UqajrzfQXEZ+LL6M8jYKi8Mr
PBZVZBXQDwQ+YX8t8YFZD3Ond8ax8/vpzRynfi0MufPkguGEnBA2nslMvdSWoiWM
TXQJHIItnuXXfX6+10o0TYLxTpztmP3jxbtWWluD5ZDT1J5E1jSou11xvwE8N/xG
Ev3xDD2ap3HnN6CcrOMenOyLad50ow0gkpMYdLz9yCK2HVGzUjOTUZKkYFLFHYSj
dt+Dw2qu1VNbJdJRYRiC/o+MmSIL5I8G+iAjW+/8SaiU5RciJu7F4ieKlPqUgBh2
SYGSwfwHlkGxWWBzf+l2etEIwcC0Cabg9sDYplO80n7aINibjBQzNyUKV10FsEkK
nADcD1MB7mCVwVGtsihnPjT2m4iIaLOox4KO1H1aXgFMco+g39oRkFN6Q/7tcuk2
kIup0tjOkHITU3QNNepwoWbYv8zW3yXuPw7MEB1gDonm39sH1SwTE5kjY6qlArae
brCO05+rksKsHP6mioP8ruX1qa1WOKMUIh1CWFwMbL8q+4SkOrRiBCLoCYRHiyV2
7rlqqnSqqnK6QXU5PLROu+V81bVCZKgu8lV0P8pu801wXvlSsTzh6kwYurKCrNOJ
u0D47eMLIQ43RZWsDnOCOT6V5VP2J2JKYJAf8sOlmx+9u9dhLWdR0SDpun+9cwaV
OhZaCQKg3XqwVf5/+8/hIrXKcK+SFKAfVxq898MQ5/V8pINqDrBDvRmFaJj/Ixwe
LXA0j+Z5cfhsPRKf5yVIFK0GaV1e8lVl+62qQrZy4M/tlygs4FXCIgVEEu4JuTk7
724p+J4fHvCDVVGUOHgFyy3KCwaJCQdm+nwteRwUDrSc6wPH5YR9kKEW3MWEr1Qk
JkpQ1Ra82mdIS1+KK7h2lNhJmQuCI7zkjHi7qqJcXnOqHfVhUBzpr/hDWrfj0xRv
7z18AZnqwiKh/XoOmkLDNLm5ZkCZFDVPWcrv29GbfgpOFYr3ihEsChVVg0sEuVjJ
rO38vk3rINnt2Vg2pD0anzkRO3BVH7DdxRFO8Jky/kJIWiLcEIcQvfmNV4cH5Ahm
hwNOsUQPC6dJnbHz7eE7VdHes+DWyp0uBe3TR2vmTUWRnLZJbVO1DGX7MBEdBtOv
oSTP5I4JU/uaBw3P95qVYdpoE3fGkRagDIvFtSribQqLaHIG0aK1RpgDqgDLnzOA
OQdfugB+pwfg/qYY34kUZZx3NhUfJwxUJ4+h1XR59kEvlS+sLCT7/JGUu8Asqtfi
bdQw+98XC4CR4K/pIK38wkx7cBibEgACDXFnzJgxAKwY+jmujb6McwIgIxUrcq0T
0tUsCZGH9WmVgAzs6Imiv/GEum5e0n/65EBefHHn8ZsvhMEpUX3LoJf3pLD+kcId
rG99DEdgGB65itR1MrfwmGsCFbuNbdeRloDp1SlkjSl78V8PWufx0B38pQdst+b/
2ArXyYCG3GJAC50Q/7BKk7r7651fZyNBdfJrgcN+HScR4gYzc+5kpSIFJ2Qu/lGy
UBjNV9qsuReg5ydWLKeucB7gLrWP/aJXuG5dmiuX878KFa6JnFEG/k+stTWUC/CX
saf9OXxY6sh5Yi3eKawSId3z7Rg6Y9LZED+yJgAza6m3Rn6mNRkGt5lW244CQeAs
WN82LngYum83jXPk1lYoOvVJs5mYaiAHW2V0BmAb60fxzvNPx0kblajT847xgimY
qcybvFmRLzjaBpiBhQe7OemSwHEW9SLI7KTy/jxJquKlQYZgRtTZcKByzSMohYb9
DiSxqBLW6w+6sjuYAdK93nPj1vjtZmo36KK1UwtYO6bIP90H3SEpBmeWrKkG+qon
wrAb7r2d9irUyItwep9EZWVYW+HN9vPTgEBOJZABJGwoZSW9bjeZg+D1tKl5ZwE8
Q5xOE0pueHQKjcoa59xbc8DEJKo15w7pgf8K6PODFar5AZ/1Gr0A/4mBpPFJtlR0
jZtBENzRAdVMKOpMwtpIUHI4klp+llf9WUdXtudL3XqDM26g5q3bP3PEFGjsvQOI
cOZxq8HihBKUPwYVH6WgvsLZ5AHwYvsTp/V8ynenkKBeVpgwv6NKaXJ3nM3X69l1
Ld4kV7ZJHU1xZrP8vwTLwckVfi8Q0+TxU25opi3/mDTHPikLk+27Uk/7rYaWu8fj
1sNdLBBanf3k1Muo/5qaKcdxrfjxy+VZJFjTTNMd0oO/afWt7BtMVF5VlS1TZwGf
ZoqdSdrulAVB7J7XIh5MaT+tkzWT3ORKcxgh2MqCjXoRlNHLhyRapTAr8e64wii8
O4N8VsJ50UylUcI13XC9xCqsrrvt4GjDzaz/CfHTy18qD4xnYNuPmd4w4M1mveGj
e1vB0PWr2vJ5bKoTolJzWxnhYFiVxqEeEfEC3xwQmRhoIdXoOoIYbVp6njfCJ7bB
WeNqpun0OoV3PFlZ14J7gfn1XX6RSNilsJu5e/Oi69IiqLEIBk8kLsSArlPNvVMK
Ag5n6wJ/JXaDJ/N1XWOpMccQMolq968qtdeQ6xih/OukNTBdGkrst0kCOVmJTuB3
bxSASn5ThI1oGNhpHMpuLmk2sSf5zI+pNvz6FQGjsJDco+pUM72bpr7OOyn1kv0d
gGJohxkIAtpyE9jdeEo0CIZ94d75QklF7NRZeG4ipwtye6bjuhn2b7rzASxmczjq
+w6KlF9O7QCYY8T0GCyoHznHkl3+TtlNPD3P+2MeT3MFUw4GVakaH5c8DllnZeg1
xqOKcOm8bsC6UTJ5FEmlD4fWdgRjoiznbYB9u7fYTgEHsNuMamu5G8UksmL/t6LJ
Uy+zdnaXoKGP+WFVnMsWby7EjBeYzLR6doja6h2y0T7jKVvVuWX1Nu56bDvzW30C
kdYSYGhiX0fVyjSk3LNbHU30vJ1t5qfFAHdTKw/LYyx8SxEAdsNrbMBZTA+UPtxv
SkctO6SFkvkuok926FLqZYROoavY7LpDPqcGnfiaPTc+r6pdlpJPmTfypqHJDqDO
5pdxyTiWb20tB8EFzk/G7Z1c/g6JSPF+QzxMwws2ZMDEU6Ia/ZvEtGX59J5ddOze
j00kOdArXwhnHHbOuRHkYvj2ZEMIXMqQdHsvT7bgrX5dInRQwJd0bIz8hpqFcOg/
9/HHNwPc20zhwMXni/176VU1iAtfVl7iDMVNRojPR+o4XS9IBWqbC/JwoTqTj4f8
aPzhVuDDSA6U1vTy+zthJwklsbBt/JUEY7snz5kRBN/r6VtJHWKVc2NLmBMCsbLC
ab6T4eOaCnndWR2IE4bA/bEpzF4Mc7wacjjT/viAZIMkGgqs9zzItpnCYYXbpZDF
8qim5UmM4hacsqJNm3aSOHklSgOZfUzSCMldb0gaPYedKbKYERJlH6MdAOFupkNr
c1H/haPm4wnja38Gd2E5ViMWYGBVB8QkJfbw0Z7fRGA4fbn3Aub24N+N/ccoSFO2
HlG7K+aoJkZVEyNn6AAHCLa/AKiXn6o844lhfECOI+cYnccuewU9y4BYdmecrUrm
59ZSYOVrHraeZnj4O9rvi5CSiY9PmBof0GWabLJlPRX3Y4OqTILsRAgxk5P1WHRd
9klIXfH8AzRZSPdJIIEw+o8GoRjkdx6txXOP1adnakIltGnLq0KVGpkVwIDLiAd9
8PUPYzbB0fenlGPte3dOplnpmlfOZ66tzsCg8RN2U9Dj1bw6lGdjBWmopV4m2nfn
hQHTwPbJD0OBgKj1ao06l0ejiiQukZkf6Z86hOJsWPD8BqDvKS8MfvoHSPi0z1+T
Ww1SYtVpm5YX/JVsa+AbUeuHACsR+/yuS6ZMXg3ds5VvCodRduIiQQOhB+LN2o9Z
SHyN0zm7AMEDvvjwcdVuX73vjwaWBv056hiQQj3oiSmZld9eYShDJ0nmfDo0l4vM
RZHbwweaagTglVTwGL25SzZz+n5M6UiDSu12Gr6v7QPUEvOMB1KC6nWa3QkdUAvl
9VjMF/aiOvciZ6W2IYgJqTpPRjCTTcgQg6z639Jx1qKbslBYFw8BOT3sTIeyTYDl
2OLyRpEExzeEoUNFvGsYpgREIZKQkIr/ZUgFPV10Vb0lJlRfD24L7E/hb14iL9rJ
REwJQC7vlY26c27zvQYjv+tWYMuSeWXNKrUlU4NIKDPDk0c+wErpR0jEbBHB2YOh
oTDC/89SOeW0BigK2ReG/nDyOk2lv8+mtlAHz8V8hxjiNEYbT7wey0GQExPZ6u6a
tKk7sg4lxvfvFaFKIO2vsRckADXnRBCgBGqNLMzxD0+4U/DGe7LSQH/B9pyjmO8V
4x8XOdLQcv9JeNNgH8rA7yKuvCY/NetGdsXRlPCgPePLrWKj9ugs25HemBRiaSk4
s5LOUG4/w+SFNEwav8k4n1kF5yeSSSGfw05kRwibL6nEy7cKCPIMb8og047TUWIj
F/WHbONS3zjG/f5Nj0XpQbmmal1fZu8253i/lwbenjcDVJSlNEvZQA+cCzQ5i2Am
/043tz9MUL3X3cgqHXbgWhPUe4L1wCRz9VOGetasbFBTqr+H12oKvpN1z0oPN1iG
j43cdFVSoCbtc5TY18tVWpWSNYQM3G6c0LeHNR6y/JbZRO3UBAcNjtub5FAS4lpA
8pUPKFA/Z0BR7clKJxfct3KHgi8ufNuZAqArku5RdZQ+FRIvgjL2YzNg7xXFi0U2
asGE3vsx5AygrDrTKTURsF9N1bhgTUP956iE8n96pABXaes8s4zY/ung8R3Ht2a/
446HAoiW77jVxAVN0dRI9vRW9tjie1cBiG4aSQv620CxUnIbjEB6GBscNzhACgDF
a6Chm7dWmmyTszEM4/YO8E41JCZWgsP8t3nBnhwyC2hvTgCmNGS/vHeANqNkaj+7
SWRf4OELNclLs8X+bA8cGiH4mPa0a1w7+APZl8+YwDWm4qCTpYjTJ0N9Pg8w0Sh2
FbJLvONY8DFx5xVViiwG0Q93aEoRfs66mD+wQdBDww8yXpDHoAHJxOIPz1/hT2co
Z4GsDToYOyiysLw0NhMY9AMmViAJg2E1GpZ4mi3ozMZh+Ow6INfEzU09ukevc7CL
9xplIpOiPLZAwSwiehuK4f3r4XDeQnbKeBGjlktfdrN3mKKYqkxfGj+874vB5Laf
6/jhrjb6lIP6ekkmZP69lytWAoR+WIftWL01c3a02ue2svbLHX54EMO/vcvtx3Pn
x3Oa8lxILV+1+SDJbuEcZCUFAHTW72tatp4JxySW/SYdZKrIl8Kx4wt0FqTa3tYV
8sIkHRnmBqYlGBoJeB/Xlm8v1Qr7ZxDR+4XK+pV9z+97+2p/cEss7fnkELUgPcwv
Y+6Gh6RPR7Dw+67K+08sSgJjgrtALVIDHhsx/JTq/iTTopI9r5oGk1VDd7Sxy4JO
uKqqhCTd7NBvgaA3cdGmtT0P6SoFfUu6A5ff0FFJjUimeyLPLfbWu0A6SAUIYGDI
lEA4s8OvIEwlnYYnbvDnHfdQhRze40J+iaeEC6e3LilZlTm76hNBR7CHMcwullAL
/yiAs5ZhF64Iq82A6A3ke1EBrdbZQ0FnAGbQMpunCByHB6stRyufjrBziQMEre5R
MpuJqNj8khROZJYxtswMaZRv8KNw6H8jOwn9i1+TzQnGNyTeiWxLq/qW5pAgeWhu
KiK63E1tVNJzLdsnPqZVNmnNLHK1WPcaelyMA6gOVnI6YKYBhyHvjvsklRrMI937
sk/JdohXARF6JTIm/nn/xMEZXmgU94HeO8TDlVmOLFFPyLbsuFm8/p8HZWOgU2o0
Fcu5qf1hi62MVxGQZypTigVx/TpR/3hkko5GFqNzOl1mrMSqZz1HlMKKXPRtJOqh
kr77DOuy/8iU5NUE+ack80FnqcwcEyVJVbISc3bGH2ZxgUS7Z5lxMjsC58H9Icsg
xfpR+I2xgWuGVOIuildFZPmU6PBVRrUJTMNX7QxNRdl77EreKZE4EIkzqJ2tzxEH
M0C8gwRRmsKPQdqaT3LrZoA4uzsiQ8neh6Mum2O5MyoRZxJ1DJBwp6yPpaRTXcRh
NRBXLpHY30iOinF6ASzrBGEIkGSUJ6cqBFKwftgoA646VGc8tx0LuVgMcqIqT5rh
lDEV4+uIX5iP+D/m99iJ6hRiOGg8yM0DprSM0SQb1KdJBaCXVk8ztSHk1AUxSMul
FokzA5ckLXoPt4itgBjKKXX+pno1lzI8d84+F7wqy/6Qo23ISyj5tkkLi7lR8Fkq
uVu4HKiop6noe5fmKqXIhbTV9pvZkfpFD9uU3+rUmq8s7UtCKh1/JPRMfBKWQhA5
erlYqXUICfogRvHZTpDzv7Vy8VJUgkSJW07gXuZZXCgGCKMJHNKtjun3uqlMF//T
mR6Ox0OO0+NXetoXQIlO4mE8w52YSAw9kQDQouvuEk2uPKJ1zArTDjm9MEvBrLCQ
Y4xbl6VeO8K/hiojVm+f+l5fIqn8YhzVud2zLwIeb5A7OXsB+qsp0uerVzbsI5EG
SMzVljw1X2fBeHbqsIjRszSGvEnBtAL9SlxJpeW8YLqOvXwXf7mMs2mBfZt0YBGk
Befqx94QFdz4ApZ4pPBh/CzJPFyzd1b4PvCzKB8vENGUGxWzN4lIBq796BIBoybF
aeGW14EPuJ/cjTVyv5FE2SeJkZZv9hUomVCaxRYBMlFCbuog0+2aFxEYvRNbjXXw
F62tqAbEIF2e8RjehuHfT/HPrUo1O/wQprqB54D4H6e9u3A9KzM04IPlE9kyWqSe
NL/YVYDW74f0V0ZFcjs/uNbJQocS0xD2aesQ/VIGO/MKHf5Rl7nDno8hImOXb6Gj
reAEgS390PFOxNmPZVXsO9vG5rAincKZoG6bbcxH7t1WliXKCibC8oW+PKlCcuNr
idXWtbXIhGk0S30lb/HQbpeBoRgX93l+t8kwIth3Qeud2KKmFhYeEc6WnxvEOtkx
lcVsN/6X+xZQWm8/WSn3Uob47f+tkNdLw5h00R+6Yq6tr9SZxo/sB3EJO2Ot5Rhb
HNcOVP/xy8Nsid18IJNzB2P9k/7++HGdqo+jYaAoNQpO+UpOneaJUvyZirCEa3l+
aZ6IUKxhaAfPRDShqs5R4yLGV2bWPs64pCT5XG/ISE3TujazpgxbzAJ2QTLJkOM1
ccc+2NmLkNuSlClENCF8zOVzD9WT0LIOEuKOcAr5NM46SNOnRan5fUP96Jl7caH3
Nxr0b2Yepd6sqEx3Xa4xDavqUl3XQkY0cS35wb98yKQpua2xRgUHGQULjaJFhuDt
acx+NowhhyGqWtASyfuo12THpBKhV7XQnTYGcr6ELvTmDGdQEkssK9Bq9G7P3NcJ
ZqmDHPa3qh7C0bGwsolhV3JJbulYksJgHJFIYw7NoQ1FAf/btbNKa7+KDrBVamlG
4W57xC9V/rF27TSy5ue6HdxKYDHtjeOUunTQ7LhSBCDeXhi4677Pf72y3fU/DMqi
bOZVL0sF1g2hUGSuspzcfNfS4HSHiX4jqMLpBHbd3IWYPq9IUpzns8oAIr/3+ohM
OVSKixTJsMGSpsODKbKKuy0WtavSJ90yMPqWQcUzG2mVpFntIaPxVf9UQjwYvp0S
Df7u2bnQ/lpJLTMvFBc3BzsS3hCTtgB4SVWdVAJ+BrNapt5MarELnRkzxESEEtxs
+j3qXvIIo4RB6yLhHG5BlPHkS01ATjXePgJ04VUEAIGqY74/bGaBiOB4HmGIJ+69
PGOcKuq2D81vZVUPTbyoxrNY1gE1RvBa+QwpUJV6brWLHALUUmtB2lZXGIzetK2H
UP9lR6n+wmWK/sTBEGe+b4izOxBuP3WjXy08+tDD8bmd9c1w0/jWb/oGFTb95YNX
/PAcwLL/ubRgPwCY+x8EeQOC1aHVWWOl8jTQOqABgVwV0+Yb6/12O2TeP60r94Oh
n7h0xvbSICsKL90gdaY4cvQfDoikFI/cuWpbQuz10WFzfeYN18PC2uoyEzlTTq1Y
Yup4VyDWe8VIsgld/LZqReLbvLFP3AKODOjxqv9qcvfdXY0cTN2GPS9mSWLlQSm6
2zJRvNsh+VC1Iu3iZampVmdyV5RZY53f95xpr+lXRhbe4jq3TTVsTIG0oGFJxHhJ
HhhuzQMbcnw78P8Z1vnkcfGotoLmv0/1LTZfFEbsWHh5/qnPQC76j5KHBO4pmXTL
PHrJPBKIgabqEpUsjLZlW7omt+LmD94LhZ4tPLe9buNEhZMNFKSYjPHAQUvtn1fv
FU3NDPgRR4PQjHE4taqG5YEJBdSk2plWD12zsUbHa/g2agZX+Y4Bo9HHTQ9GAdyo
LVTQPJ7SW0Zib4ZJ+NgQDnjFiDZagqtDrYwZp5q6cBy0hvVgUlVqw4ff1AEZy+7V
A/rG4PZKGMZoUFjb2+FH+klGspJQVCffS+cYMmc0Ioa+ClPqZY7oNsq7wlQl4gWI
q9jjOsKX5IwEaa1u39FuOy+MxAE+7JrpnQaJKMocg7nb9wgKtM48F0k/l3/x8CZ1
aY9vLHkTmoN1e7ygaM9fvqE5pfdcF+WSM9rPqKT6Osag/08/m9EOYAmVOaYtdQrH
6B7DRHQs8dlMvFZKVByZZAuLp7fM8S4r4O0sKteTRvTCsFAxRVvsWSY5/696XbDR
3w41r4esNzpt/unwHAX9GH33AAkkg+ybEvlAsRD5/B/gytNIuLYUR1Jc6obkW813
PkIDldXk1QtUqRdiNPdqJleOP3c33ZaDAkGJvfg3vGvXFd8UKFNGszBlpo2fN0uB
tCY7VymvPnIziUSyCMN/wfgXSWbH4rS4jk2AFUDvlrd1YfAOViTy+EF+b/EEbS34
Dh+nkWfBTikiIYAm302IGF6DNepe7ykK0EmL67lwuS4WdYbLVCpkAGQYDd2ov53o
ESUPlLk68PWx4d5RgaYoMAfLDWTOFaTakH01LxJjGtiIvwAn1RCn38k09ZsOTb6b
1Sa3M4TpuS/soVP9bbhbIhiQuxc+TITucci2baQyo37tnuTGeP72VDr4+ehS+AXl
PCSlzHPVjSVR5KMg2D1zA/pcfUzg0x3ocGLyrC0D25rSLcrEEj1i51NOs847LLZu
zdfHnTskqmggiBt3bR2sMgmsF/YexZxs2cVhF4AUECvP8xrtZbXAzyxLsO1iC80X
SyMwh09ubu8EkOhjC/An9we2yZSahwgcU9J4Gx7AvF1580EXyiNvgm5tRH6g+cAO
nWdoZP1qmVjKIiVww9sji94vKtGqxB2B2MAci++bBOkD/nXtjyy3cXDmXdR+wbbc
7BUwPT3RrNwxQm6nGn1xhKsm4pC6WXq84xPvsAG/g6kDJj4SG1q1MmrXsuqTGmzj
Tmw8mL/mjDousZ0mXNoJT8IGMwj2t0CFUcvx8wxo8a59sh1k1jQanj3FpP7k0q2h
V8MUxjzNhdOO1ID4PK+MQuQfvkwPgSmldqfu05J+9tEL0FUGnrQRRSh783dLrVAA
8PN85KHNYdT4DM8bdGEUd/Cg0L+yRtM2ZK3qZhuNF7EUrxqpovLTy+y47Mhw5BzZ
b1kMgW1V4FZVp8WpyRlOAjlFYrLwHJHhPAPvXJiEa5X5IbCDhjsircu65nnNENea
SHTSIHUjuNTyRp1Eu/vrgudUDGjfql60V70SwFvM1aUW6v2ibCR8MVpkyPC0Q13O
AJHFYU0TqWvoD0SjpyeHQBrzlJdGzCHgd0gCdZixwdHMJFAxOsGNb7sucdmAOC/P
iJaZI1qVMLMVQW8vxi8Miw2cjxsUl9UUTh14RbOSfRIL8SG0r87PGe9iN/9ErpXd
wWobccJTcTrhlLhVQ68vrXiLea6Jj69Voo2zX4nGR/djXzpWOsqcMTBwSlqwzsg+
mIIC+5MMYDABol7L1hzp6QJIi4VhLm03KVPJwYrydBM0ai8EDRAQ9gcsNJ5C/OIb
T1iWnwd2DBjksRzSEXtv9ITpng7pyAHsThJdIofSFhCVnjWo00+/mAOWpGrRTmz9
CxUwfnJouJOF/Utk92MQA5MewBVx0uirhVHObGSoUn9flO1GATih+uWtFzGjlWxZ
Bhf0Msd6caZChWglyebQE1EAQnQblCJfks8YH10+JhR5miTUIBbLwfosiYeXfJfF
LwD+2QEdN6YKxbAPjpKrbB+pXDlJtOZ4HxKWW1WDZ72UOqkE9u6e5nvFi4eceq3B
dJYoU95oakwMOjQS0JIfaEpdj7duMhP9aF5kTjkMcmuQ891k1uui+YqvqNOZ1EBK
4SowYHp1GhHW3HMpVyrwqhKd0tNJiFp96QZsVcqGCHPOJsT1EZREpl2s/M0UtBtC
NQfxWRMbomTO4idFPfGnZ8FWdxUUb2VbC2Ija+oE323cVBVu+Vj0/VeBghRxrch3
bSKGYBkv+aaXQJ/YvQPQx2bxrSx8pwx24MyxPpUyEqucIw4C6ggHKOprbDMDChDm
XZ6s+r6prqM0Z35554JBQwA/acLDgXF9003rICNozep1SHI2lLkGkKj0ihqBpzS6
etQ2wvlkono0lkk+yMH2JDdmKMW/H7NRNXRGJHoY07QJSdJQuy4oHjiclbQdiIJ4
9BiYE4KsKWMT5uS59GCe5KP/OXmmEFfogLwl/XRQZGbxlYv67UgixHusQ7kFukki
o8FIyzJ0VEvpu5dda/wcRJLnx44jlumc1j+VXiKMwp/NKZ49ACRU6tJT+nK7jT7x
VhUdE4mklFSrodCwORiEDtmByjs6NLU/WGAXN876Q1kxBgTyyN0mUVpyzh+NVsuJ
1WDQbQCfdDYmQXxIFky0oukxjmAGSra04AH9eAsj++EiUmQwsJgsGks+oVr7ApMu
eDGRx/DxQTNMb2OnvJ+x9hLatMCd9BoEd5XrKjIZuW9W4m5uCgLaVUYtGjVnPtKO
LoANt3/BVSMoueioTm6iFSgZNckqFxpjWfMyu6Dzasps9xzQBLc+ys2HK1lCYauS
L8N76D1PY6lu8tq0O1BshYRXGI1oF04KBoZaxjb3N/8Uatx0s0IqzPCDr6lP4W8K
9jMlYQ2SKjTBGI22vRdDpJt9q301swIOfBkg5GukXckdLkuGygPwgHsMyI47ZMwR
W8SsUiPvORkypEqUaTwgB7SS3mIsIMLEpi9HSVccVu02P40ANRJQOuL+i1SZQYA4
fG8C6u2x09sBTbp+ti4Qn+xXo+rKpHdv9/mZcvlH3i0pvdX8XztDfnqBZTgzKdIp
YoJZWxcYL5fAPWOCUWVhKPXZPUeHWraXdLm7PKfrdYvjBkYCaiowj8aPCLCHyVho
ZRAgu75HzuD+Ycmic2pnQCqtjNiACjzjx6QEjjasPBm9UnMsofqoqWOdds9vn6kF
Fxgn1CWXSwG00E0l1uKMeRXu+VyKPPls/1u6GaeQrY8sKfm5zgHuf1urnXBmA5yl
v3ASsjmWKgjkChC6FjQEAzrAc8kzZAX5mjsaUV/3gKEWfn8kWv5gmsmUJiey1Ica
bMwPUxF3vuaMvbEv3BMIHYFqUhkTkfeTpTI6HbMdkQpE3TOGWwl/3XA4IYQNtSY8
8CejhIAGuFxLoKveXYe26EXYJz2+WIgs6wC90p+8NGCeaenXrSjzDMB3QC+6YkQP
hdaX4CMSxfj6RDvNrFA2GCbgxTgSqvepPQZGM/P7d3XJT3lbvVimWwSbO+j+Wy6I
Ff9irAfLQrgz51NuxqxgQu+frfQslsQbV20CdwfeOZ5rlw651yBPaVqSgu9EeZ2l
Ic8eO0PzGfbEZr7qWFxuAXK0S4F/NvMrdk1X+SUh3EchKT3FZD7RCEQpxp56OB5E
oqW1/m0kQbqevddrw/7TzVDTKoXLMxE3oUl6hwRqXic5CY1i8ex/6Z0VJ5DKvdJI
AY7TWuJD7cm/A9CFadlcMbsGVIhygP+WjuyNjVo2wRbZbfKLiD0/eFx88PH5O2Q4
sdhb++lwYRbXwwHBpCusZ4R0cxJ6WjObHftt1BR9/0ozQbClwuJyBJTcVmHM8m8K
GmUbNfuq9FFnN7EEVJl7pRK0x0xLiac22cE1Xb3BZqVPxD68k9FTL8q1vIBjlo/r
om38x5gvLpq4u7+ZJz8GiSG8wSnN5vv2Fv3Ra8hzh/PlTGQ1mmPXbhuUoN/4pTxo
cnHauL8YmqSNCjjGpz4zkQCfSRqHzJ7qd5GLOUkzdKCkzuqWvDnanHNp7xM5/qYE
VrNSNj58cStq7nj03FHI4PtTzY9BMf2DRw1mPAxxPLnTaIWyONgUVZySaNd7u4gI
uXz6Psq8gZReWprrgl+jeC3YwlYSMy3AfKOuEv+dCXKdd1WA9H9WalGMhxe28xap
+H/9LJV2Uyu5ULij7jUtxAfi5+JsvedB1bMyup+amvZdD1++Rn1cmgJ84ECWjaZS
/aq9JpPU2YEGrFmbLk2GEkELpZcbqK7TXAb5BFNnN7vJQMZ7+OFGNw7zh/h0UfuF
/sj+MNpCSoU7SOeP1bC3hAwkMYsT4coW1imgYNihVEAlUaxCh3lGtGWObio+OSI/
uynC9yo653Nbzr4pa+lID3PMqW2BZFjRA7SleztsnvWAoCb6y5JccxQSJp6B0nmK
8zKZbvd7vWxmvsq+CTG2jIAHZtn9REhN6bwASCCrysvJb1+fdyVlTnEHKdFKE/6E
FN4oz+zST8fLEGsPgZgUAShRyxU2qwkNPiOuBOCHg8T6XhtJdHCV3RRUfGK6+658
Tme2lMe/BFdXLp+hYmTehGVua587I+31gIkRh8tR7iHc5Nfk7Ut+9zRpwT0jp18G
L8sil8YqTmnrjhTK4usj371qzdMVZMlYK6kKCYdrh4JCPfC8I89e9FglJsH4ejl5
pfRgMuRb3NiJCmIQFcZTuyJ5Gs123CElU08npJvE7uA11JPnnxVopNISn8r0wHNx
AAfWOT2ItWHQojJM98SKP5vSnGot9ICTJ05A/WOALu5XZORZppoYPDZ0+su4kY4H
/+15uniEqPDSojmpreK8KIth3v0F8NM7TqzMBnZgtwGsxnNJ7w2XxsjQ9Z6Cie4l
8XQs/eVDMRyii+IkCEWiXzZGSp7aLJiPBhR+q5gPzVvom5qqWqzPNo5fcf6wxovE
zRl+kyFMywl+TWcLDgURJdAu8TIBKTL04QOSnzj+YKAs5pTLKZeN2sk3If8IfKxy
qjwoCjr+Jm26cquiEmF8fmMDYkqZUvGsTcCMbXIh0xzSqZr2lHV4WLX0zK7nz7km
17DIQCP5FjkhmjZKF/XE5AS2ybXhqG7+cSYBj/7rZwGQqrymZsxmarNmG14ncgYG
c/WlU6yO7qbY8422vDa2YAcACmf4iCvdZyiKLLUe5/N62PZcMKUZMHMPDKwkNQcH
saQbnTsTca9eIvNMdiN16ZxZJQrFoq46h9T/L0Mi571b9fq6Cp/ha31HrtDZ+goR
G8NKK8wTDVupb/P7iva/HeirUc20vYo0iO2YTCr/qEHmyjSU5ZY1/EExco+JYTco
z3E3T+JdaPO/i78nZt5hfrMbppUcN3q5PZ3jkZF4fQwC4svxUtq8H2ruCQPSNR2G
tKfiOts5jNxosq3airUzHesmCZUkg+1Xrgemxz/2S85rfyPQzZ9zaY3tQ+v9d3fc
ad/5c3EWfj/1U18wb1XYAkGt9UZT0COmH3bIq+pFAFjc7bHca/bxYd+oU7lpOw4T
OZVSiOwjswaN1rCiXaYkw8YDLHBdckdrUFK2UzlxrENzXkqblFIxxmotpXWViYEV
aI9M0GCyKTMRzyEBau4Q1QonkcdyLxjy61Lem/npliMxYt8q8jg4LHZ5xiVpvGPO
PjzUby/EKvSnmvq2J/NbI1bXqwTHjt6otNXXlpNopNq3iAL7FNlxbWsYPYaOpNaj
fDd5s7J1wXAVewhkq4B9f274zHoaor1PeT+3KEsuVc84axr+iGNwKGAKs3y2YbB+
ASFnLX3Hy30meuIjoG4/Vx214K5sxrilwnTWyY7S4lBbLaIAzf5BrgPBUMV5zPsa
qnAvo+ETF0WTVyOKKzzva+SIj7Mfi/j8dSgH32rrCmtE65xguFbqo7aYqHix5eQ9
sH+E0m5s7p+9j80xYEDGcyoTbfmjDrUV4R8YEL60+BPvPZY/ASID7ZMXACExuOiF
jlsymi962b+yU3qlkIV3Hc6wsC6nggtyByRzklyMOEqf6yV99CVfacR9fUb2lxCn
0c8BLvSAOs8qpwLtX2xj1BhSekNgNIMFSaIQasjPDraBtFiljBf6hMEYKeSV8h2m
1Cn4OIEd1YRFQNZRv28Y/MnIFuGGnsXMA+NQj2fSh178jWTVv5Xk4A7P+TVEXJoG
HZI2QtL8+ZAFo1lbHc8fawt5sNbgWVNrLxYQ6Fw0yykWfhDgUKnh+Py/aZgo33Jq
0zHjYvrrJi1EJbA0zeQe1bzs7GbrmXcYaWG6Xjqu/uGz1VD2Vn+9mYLohRYwWZ72
xrnXttx/6NnXZq1yjepZeqvbKqSeMDjovwUjWnGGxPUJoOAIW3uAdcWv4sH0Ba6n
NB/6+LXqgLMApoeb1HtM54oT7AtllQwlw9du5MaBk/7GE7QAvMf8e6qGa0FRDY4r
WrBlDMZOal+q7P5Pib/2ClddnEVd7x11wfW3u4j6MY8o7G31sm1TMahexYvg3zWU
yOvObMxXltvErDex6SmsQuCctRP6uq+2BluSJdNVWTfIdzHRN9xEXpej+IbTA6yq
T840A84d14vdZmdiqf244WPaKvvIa9DfOtG9gdYS91OB2G7nXygqhh1QgT3Wjd7Q
IRB4uL9Nr1Q5phSfIbAcKIvWZdi5R7kOU/QNN+VVTHl63my8nWjaAsMs2u1sgsFV
s75uECleeG16iRKuWS16+PGg+uojhZgZONGe3nCPLROjc3ignDpuh0aMNRsCY2NM
FER9zxsOBih7M6odmf/MsmXqy51TTQohuViv3T1N3OX2bpn7x9btYcHwm72NdwJT
vH2JxC44DdkTMVNZXK02z8h5kg6Fv67Z9RQxdeYpuJxMEJklLA4muhBp/Vrzycdk
yA+LgRyezoh8RwX4eg+WNbfrYK1GBUK96DHAbz2EN7XCnZUlsqQTFDiK0YT3lRwj
0rRVT7C4DKMfwyU8/73b2rQHw1mCXU3WM+chWvbtqI5mLfvi6FDZB6WgJMIif3w2
wP7Qnwcvkj03aNuzaWLRbQb0DpSWJCTo8Lb3eluOA0SPsGkn+7oCm1AaVTP7W3jU
ELmQ7EobxPMM/mo5Q52TUyMrAaHNyTHtVGh6N40cT0JZps8fCF1jGyNhiuRW1r7O
H5P5b+qzpEGfuq2ABYFoxd2C/bdfcW/hv69WP5LIk83r2nLSMbs4ugPze2Ra9cL4
27SPC8T50EuVdjCPk4VKJAePNon3owKdf2CxgBxEJ3lbF0UOTVpivqAz4Cn101Qh
ogMK6SpZ5pfJXcZw8FHmVsalb7KzcPJ7EBc9gAT5tE3SbEz2kqBU+weUV/rPbd2w
q45opZdgOR66YaBo8AJ7VjDYI32a4IoeBwpO2713fXJBnPS9O80LDtvLbklzyVyz
isZtOmud/6rymJTxIrlEBHTDwanL7QcxYHAv5lpckx1oSUpvABZT+1Bg/c1psGKW
PrnjRn2kPOMb0X+FGrA7MkE4hAjM7ipe1KwTgY8cYG3Uio/YXgTWomG1F2Y2pFgk
NulgpvREkADVeeZhsXz0aanzS+u6u3pus8qUay3XR+2xOAOeu9Ga6QgRVwHjdAWt
uTn93YKdtej+0MQWJxFFmznRnnMtrQe++aT+XvopfjUd3bsrhCC+X6sRKSKfUqVU
Fz0Z7/yiuiz0EWClHGmggxtg398ijEgY+m+g2oVn4eY/3A6VRZQmfzn7AXMxFRuV
2NksJM4Yy04Bn6zwG9Pa3o9mzB+ekGkBjiGODzX2fLv7NXtWnr2BbtL5ddDEwoWL
u6dzXJFSt1FDF70WHfxAUU7LbSiJ9DGazuu/A2tEHIsLO/MysJZRuPaXVZyYdJAC
etEKwHPeSmR74cWzxBEhRa179xFba8s1aJXRKK1StkZUTFrZvXo22AoN+9MlYym+
+ESA6DQ6cNRKpyZLPL7aMX/455ihLVUAZfYT/opMLHvLBrvwTc6mpf0yC6rhPka/
iXyP4rqEZb0yH5KEOqDTd6DuLCKuHlrPzsrCjwJAyJ9vcxcZzbgCOrnmjURj2qMz
VXzw2MjKHkEgNZrqbYHqQRCioSDq4haCT9pg1N7AX1OIH4vlK3upHU4cOsiTwwSL
E3khBtfNxbLTa9fyHX8S3+LNtgAk/e66Um0Pcanz5BUSTr7vy1tarBimIsUuFMbE
bNj5EGnVFm0Ghh1zSmx33mxuInxWIWXxOKL7LuJjZ8oncNLxXylkdq74vi8+yPez
X3rK8TNe8EL5yxzs37gIqwZ2rpXGfAlxieEY0BmTpZhYtQYEXd6bYwQcxkwfZlI0
QN+2FnIIe+lyTDM+GGJRqIFr9f3ytYVJNCF//mmh3emj5U6b9oE/0HCNqCJ6xDiE
wiNavHaNRHHwiuWKZGVOhfTLxvWrgu8AXS7hXrjJnfGhktuu/mpxVo/2qMGw55lk
YRWt+1iMTxpPBtmoigUmHE0gLWmj2mmO80OvNVfj9WdscIGMjcVgbhurL71q4xZV
l6YVhsOUCNFp5S6Ef5n18mFnj9dqZDwi6m9rv80Fv8q5daxER7UdVarR89XULrPJ
4dwWOYdQEKpJg/mPoyrrrzogQjoOp9Qby4lrVhl4Fs66ItZxnWf610kK4hgscOUt
d9QWTE04DIMIyHhpljh9XW1ndwYnWzdOqzuTCETbvPAJ06eHyQWGo9LvX+4cF0ry
KNvrd+rOAZaxXQbMtOun+4r4rOfEfuOLyt6V+aPBCzCgxTm5CgzWWed0n52cwnfJ
Y+sdFE7xLQMXAK2g6niSWNhYiRGfMRrsnB03XB0I/MHrJXJm8Tf9avBpzors9A9o
km5tGrXpWWGQiCBwlpmvkbUn9ZeDvFtWTKMPJUNA8AdDiS4X0jMPaMGyXFYvaFPw
EaZMALk7TM9qMyfU6O5GK+hH/rhaQ1J46AcP+3Weah6YnDtVtu6ah53oXTIc3R5r
4YbKhA+Z2ScfLIHmo0ESISssnYwMze0QUPxIXz9RhQwEQ0BfnE1DV30o3amsyajW
QxqgHuN64SVRWZz5eei2Gucy8W0ANQcblecAb5rhDZfVAAAYtpVIZumgWLrjayPq
m26ezKqcNIxjCCybdaDRZHXN+db4n3ZXuibjyvAgrX5O1Aiuwjc1YONkqXF+e4+1
iVPeQiZ5PKA5a7vmFOsZqrP1DYLjsvjYTeT4/SKjVZvgGAPGLQBqCWKd9RWDIerv
m9TXgt27y6MvVeMKbbiZdgs3W+vsl7s7WC8nk1VFyiqzdbaS4OaWXiIUQpQ9Mrpu
fchomuYQ6T6tmC5FcQV7mzu/04m8ZQPbiJ8NXZHpwXMr5WlDJfDQ+52sZNeUsXHC
6VdhJ5/sUud+UoAcF+W34E63I3a/clN7CHSKRdAIwRoQkGv8d8BkHn/r4dzr3sAP
ilFxnmZhZ2C2AVldN0G5ZOtVWtUxP1vDrexi6kGJeZtHXY3Y+g44b1PaD1HfVITT
jveQS6OweXccUWkEqjdhFkyyld1vLODIoTDrKkEJoQV/u2rp6ddhpFUx/472mu/Z
LfhiWz6zJF2TAkfPb/WoQngtpEO4kXtESTTc6axdRYXrfRTH8+2yQmT7p0YJqlhW
ybpir3a/9wcUDnP5bocG1D4X5IoCKMr9/HQ4O18QPT42aEmUBto22lDYemCZ7sqR
eR3urFuJQJKHBwLAKjv/VO6/0brOwWqJQmeAFWxH5rp63yvxXPAfN2G01Nlu7DZh
RoE7oLs6XIclxlYP3AL31j/IFA2TTjXw0ZZiGjgClaJbmNCEQkHktyKwepJ4C56f
FoRIrbj9HoytbUXRRI4Gm0ZDXjo7425JZ+AmXet5gCohuW8imvdO3yZ8jknEdELg
PX7xohP3yygVGlRzrE+n0eGz54B1yIyfkdWCjWW0JT4ukBTxEebwYeUl6C2lM1wC
RQsRZowRdSQlANf7tDsqdouvxQuieFN3o25WGBbqxJTFkDs6fzBFNUg2nci1mPm9
V4FIomKhXCPdZSyNdaIudzLNOF3SgqTyvly6UsRuMiU2DgdyE5RvtxrJ90iTxxA3
gduiktVo7foezWgaSXpAwgNSFfhPLmokIzngM/8U5MprioJ5TEAT4DQKDI8Z+iRY
Mq1NscWH8psXPt0uQ8vHiP44iTOrd22HPUwDZgFekA8WsxHFXEXQ29+/oGWf5NTF
HbOirMR7Jw9Go24gsEOHUbbUV2jrtzI5fZ14VWHW6HYzfUjq1TX7+Nh0JyI7/qe7
/7H9b11vQMBMOSxPuAQ+/FOna8Da81n7f93HQsfBVpqcns03RygV4XPnUXmEx3Nn
0lF+9Mw08GKE5x1efYoFjsaItAL6KVYDDvrL+mOfJ0qxqgSQpOV4AQwQo6k1jWBv
F1K7C6Rlz4ADjdtxSXm3vZg7gWwD84sJMEUHiSdPRad1US1rP2sF/iOvvUcb52B3
BswJZG2uo93Rk9sHxOTSHUjiR8G4XvdIPcDZyMqwbTBuACPU0sph3lTvbbzHNNWQ
rzO+FBPRyV0nT27zJIpPDy9PuhQ/sK7TzmaGovqf6Rj7JFBiFW5L4B+d3YbVuaUd
aqWfzNSKiUBzPCZiCHELkSeh0c6wPY7A91xJjpFYYjUxV3fQ81qq5SzHmhUliHET
cHsw00mfUR0Mkxxu9T65Mx71u39lHttrm7MQWEyhhlEgjEai3aoNEv01bJvYS6io
8xE+UJV7IxPRsq3uqvhhS7uVQgMPPQPTeEPacfFirf3uo+S4LOOJbnzzyceCOBkY
UCE2cSRW6/GGf2IJUITEdHnkNoXnI25MdVxP/smE0BPtksDd2l2XvYb4pYE8FJmO
EZqUDGiWyNLEBr+e4eUhqrCq/wcoC2ucrjfl8xdRc2dSgIW2ezIxYh+67dXj59hs
3uQo1zansptV4F1vRl+5N9cIiu/DfI9ATqcWkkyymA0MeZo0XmbHMs52T8rXpmOZ
HR8kLY2CYb5n+XheXW8Z1D5YUWYzzVY8r62MjWsYNu3fk1Y5BHaKRXbMAdruOg5H
d8Hk9XBnksCWykJvQkIuUydluAjIu+QmiasGOws58oBWDCDBsc/idTlLbiSr1HKZ
aqYf7d4s47rbARAfEVWUGZrFm8/blZqvW1Sh0N+HXszY1dXurkQMJIXtPXfAEXf2
8Ia9qdiYRBQ2VC6uHPA3ScnFoi5xpiADJNqSU0TsqfGZi7JIsvcaOZkW8urEYU3u
dClVb3LxsUKajqFoxUKK6QxairCrBe3rKqyhowL60t3aGjfXsBcPjKY2TzQiV2It
0waJIysej3Q6jKzaUV3JDVrOALsDfbF6o/botnF7jAb3aMuQr/LPEMvGICYs498w
MDnQOKOxoPBCCip186+szK1i/6nHgc1mG2ubrcQGQrFDeyvS50Wz0+ZH6ZkW3kXo
6SaijO1EGxp+YcvHaAgogXGevcAaphMaI42aEMlCd2wrPSl/h/MsVmT3v0ZUKxmK
PMPeA0NAse7f/dBGXKNg3d3CDN9tW3cJrZ7OoohV3+ndCh+cWI0XYoSoydKeCL/g
gDt1visP6Kih0D+fBtzrOHI+YR1rzrKVi/C0kwQrLAL0NSx1a2a4Rn3ScG25Sd7L
OXTpfLvX20AHRr++uSOBzQ8hBeWKDD4LRwpUeMdhoRPBdqbVKcP/qUx3L8eaGjtp
eVL0KfxDKoYl1XSlNewy7qrfoD9gVyOLRJmKAXzgqQQz9/gG4xjqsYi7J57t4gBB
NHEA7X0GtA++Q5+imfOzCddUN5CKrqRIaeceGb+/ECiUTyausHgwcyxDTHocZAOS
3OFnVQeDz0Gr8/t/UgZC1YyR0jZs8vT4HuNYeTw0JHXRgluULGQXouffDSYWPUfD
6X6kcXQ7srFuqwInPKcAHLy3BluveYKhfKMc84/h9Nz3r5yd24XP+SN8amk5JQlm
rGDxJhXSxW1y/XgxUjY1EMo6uRmu9R5USeHNM6bkFLqVmdltzAeQl4qkisilV2Qi
yCevgPwk4ud1gjU7LXX+5i10IH2HHzzm1QwcgZsQ6slaovRJ+/VYx/T+iuakyQz7
Ckowqivh2jk8UFSMzKib2hHgUp9mhVfFy9FCYKTmPrWYmx2jC92V3Uk89Vb5AcE+
33Z0tDYc10nmHsY6t4iAa4gg9/RNeJfl3JbSIxln1t8rsltY6xfjFxmg+FU3yD8z
NG8SA3HG05MdmrummAA1QL5dGxMRuOqQpexN6UwcS1bnGI+fNrTpPfYmfV0tekc9
HN+CFG/txpCYOu7sG5AKSgz9rRG0BfZlJqcvlhoSAECudtCgHiPd8p6/09wO+PP+
XkSnu2oddbK5i0Q2aOKRPDdaUtb1O7PGpDQShZlR7dCb89N3f53tcTobp7LdlAl/
p6I/FqU7uxodo+XGuFOTdomZxuKPiazICa9/Z00crim4BmC69mYOtYh5Pas2DXqO
t7SG8mxREfdI842f6dsl4oqQk38XOw6wfFdKXFK7hzdf1fwuAX5vFL6BWsRt5/P3
jJrMGDj7rrMc+nmoBG18M8ngyadYwgm/kjm0PnN4HlTXqaFWDSGoKWR1/f4Juxaf
Wg9hFnkEHsF3W7GsupbiqrHK1FnMGV/MAO0u+BudJgbGKuJ4seVGchpHmAjmzAh6
9nYvx4bJohzIpyqWL+aqwAxtvjlk5BC6SIPWBWGxNIwuny+7xfyYO01yYt/ToB1U
xSZO4qQiupjcTiOFsUBk5ZtR/kdDnalzOAqd1LEZ2iGVBhISKC1nh0NGb4WwGiXw
UkEFyKZZ+uK4Vm2Uxx8Qji2wUvB1WRsWYXaGADONAzVBnr8drIjOPiXWpJjJYKA+
NW3ksbWDGTFcEmsi3592an0is6glWWbicdK6Ejj26NPt+y5Lf9iufEkY1SFrUwg8
HZavPFeUtmFiTUeNmviz0TtbaQkNrtDltnCpmf3H1PBhpvfmmZR6tyY+Rz8WMqFk
hzVA0pjyTdtVKQj2qQ3/bp47KPhLSVfFOPlGZs10FhJbpH2vYYQWwCqGiL6cKXbP
ppdhm8MGTExitXi9KCVWYZUmo6TDLCLC4p0aUACFDkFBGUAX8UCcvykSBTO7GBbC
pDdP80pzq0xqKMYke0hYMpCoe2e672uz8cJxLcMCO/zmVSYNA1/wJTPXMOP7gEmm
xcN3dbp+gMAJBI2oMwCNEtD+z+hH5M3DVRkR19I3/k07E6EZTiygaVL2bqPZHWte
hxqXy3T7UbhAhHSXPnCaVEw41aN6kwhUAWtWqnk9Z41b4PAJI7x37NWROug2OwIs
I4MvAYmqeEiPQahZDly+VfaZglt5QMlPr0ltOsywevwjnA9pUTtg+ScN6gMxHOB0
AtggkLmndsabaQnBOQPWKGitsRrozRBaqX18s1lLwwdRbuiFYAQYWoSQMBDZlJOm
0s6UdoSsYBgw5jpF5aFHSLV9oZxwU1emrGcYSMrgyE7CXtqtsoepKpHiRrug/WKo
qfrsfywst1+t29AamkQWkPRVbkK13qm+OSJmf5I4HBnr+MVlxftxd6UC8FZg3oca
vPZ/i/f1wCAwNFTkYN5eJ0rZOrLsMngc4WHyt6r8K3KdRUrEZFt+y3CO7Etm+MpU
3DCAKZQ/RY+uxEyVYHeHWhQjEKX/Kytq8s1CxH9Wx4l9WiqvaAamp7PniFtdmiar
JeitQnTk7sAAoQmApHT9n2rO/OwPj6Bzn8cQQvRg4ZVhbLVyQHKNSkKspWPfeecS
RvZs0izko+rAJhAyLzQrcEO1Hl2a/wb/QLtYf1eCAy7Ek3N+N43l5W3OHSS3WIcW
Ryed8yZMkmw3sv/omr1cP00fEBHA0HwcTzaZEelsjlHXBNBjS+qoHWlYBUNXWdpX
lp8c32kH902wNI81HPXwgshUw1pxQNVr9XvmKAr8w2qZ6wb5FTeEjDjpj7D9/H8v
YggAAUCf6onOxbpjUuiic9stkah1s17tv+pQbyXMgAU1z66i+yzyPccAoVm7LgV6
iFTSakgNrikQIKkzNDUU2pKD655Lck2KOI2nF7BNVYg/fTGUi2lQvAw0pNG1S8CH
jNQJs9AkLF8aNCe1vhQp5MXnFRxedu46+WXQHHbkqyaEL0JMWqqvVD7HsKmMKz+4
OdoXLrWkEhmI3sUajaWUFxgCysZ+pjYpWaKjnpb6dycL0qykIfIHhP6hmUSmK3uP
RsoVW+BILod2ZaL5Xj6hhR9xrCygeZiK1yFUUqlDHQT810xkm2CwZOusubxwPSJJ
r4z1BPdzCs4+CiAQ378h8sTBcMerExai/ovYfzR+R+qIqLWRHbc6gGgNAXjcbwHI
lN0q5AvCQQWvkdfkgDTQaMfpsVaD9ETarCLR+0O+0rknN9vIye1Kg3F69U0nK6Gr
YIiCvV9xTzhGaSx5UggrG8TUZkD6z3VRnB7dnoAW+FwFWCSiaaGxopo53LFFQdAg
IQbwUUrKr/vJj1HnMgqFDJRr+nOogEqwnJnXWQXXeX+IynK13mJFn3MPSfqbd/RJ
r7PrOENLb54900H2RNErNr9xmHVufn/WhT2aHLubVb52y92oSHqWXZF4AMscjaU5
wWvwcmAuKZM4Gt+lZThDwzsOr0SC5BHkBsxQlkYFdQEpyTbuGL5mpCjA9ny39A/A
KgFz9P636iUwtEUt7rHdobaeu0bvpSRTAp58RoKvQMK1IPhSi/+kSzUMjSLI8KoJ
vzdClESDtTh2hQ/ti/6g1rG7CLIahuIdddgbJg3nq7AQ4Ei+7XYd7OAaInnrYFuh
ybbIYFgy7Le4AUhOzJWz7ctpZL8SkYq4e5UuTveMEYn2yXbPwajqZc+OA50YNbP7
VArIt8ZP6VLFlPzfU6MLXpokKlT/TiDg7XFmU+AGn5geVSYpRuFBE++Q0KyFvOv1
bovs/Gd1KsGXey1CLb/RyhK3PpTv3X5No3M2gNTeh+S9r3Z747KgizKAypLnFSZO
CuwMRRQgT8smXd6A7+ecst9YaP/fYBc2B0kH2RCd+e08bNyWiD1lMzuB2IVGIVnE
Tlr/DrLXo+0iDhhiOF813X3Z8baskNQfkHcoWCZM0WcKBe7k9QaTBuMGh1tI9cYg
sr1YksbcGlWMHqT2rRNPl/o1LsCCm9X1ZSYoBP3XV/kjrmYWj49Khaxoy/Kb/bOU
bghCQT+PHQG50GJ8w8tKz76JR3B/G4U4dxTsxRCmJx6iCpi+OHl/UrlIm7caA9Se
KJsb9r3sqgtI1nfmrPkXvqt2vIa5IJcjgCM1+7/CAGYby5BJBM2cDrywNoczBCig
c0kkwGCL8WtZNGoWZw4TyGO9qeaAFixIcWBKPzrZbrSHb/Q606rdH8oFm79LLIqv
mwtr0hhqiLXSfXVUgjOceRtkQuGsU0XSpDAcuQGi3XrFJqUevbXui2l5taXgWvEV
kkTZlcDIG/lSfUxZi9iM5WyMZNL4nxQ4lpPUM8cw9bRNkHMqTfuVWbp3Fl3bRZHa
vhlyt+E3kCeIZnuKeh7BqNG4GaO9Hw+PHKxHoAbQl1RgTFo5XM8UnVLPGo6UoNkt
EvOOJWg5Ry9rf8hvH7Lz64McygHNvP/K3farVJG6bZDMRkTNC2/KZdPqvitpCyqA
pMeru6uxpPCoXMhZi/gO1Py/sp6q6LK2maOSyrdNVI3XCVDA+GnnY2ZcN/ncdf7N
TaPhGXMkdQsOxHKv7lsR4J+j8lypN1lbxPjjnjYf5zVNdL4tlq1hnTQ3I/TEkR++
xY3bqd5W66NHv1Jpw47BKVaAc+dvw8o5djKQd/jQz86X+wO7lsWWkqVgAcipQote
lsPunglHAl/OpwI5oPXWhCiJBDQQVzbQhlsZO3yEJlSbDOAzxnJ449n9KCwttLWF
pO7t5M5kH3Hvr0G/ofG+wvLl32PwQleAgDLYU7vTFlCRCpZKi23991jgSMiA1I+q
lR132/YdiZSt1iVWhlthpL44Rftky/SISSnN1yg29JxW3r1Xs3pnLklZHy5zlLVa
aPKIyNQnEsvO5dZ6aDhiChNbz3O1bVW0cXp3YBRMGw7gl0rRGrNGXd8BYN2e+Ya3
vZOQ4paRBHcWNC2RkkCYD0MuSDoCkbAff/eKOhRzHNPZEtkTm1c6rqjrhoRk+N9z
skG72syx0u+a+bDsN6nUhNVT5zRskuMXI/+XTVXKTnQJGWRwse0e48W+CBGavEuY
WW37VMdTu+7YwgcWspLm3Xi6rB/9hQIkqCgEstZGUYLjPmHakDvdpkxbHrtqub8f
lVrmfmQhtWW3Q4QIgv2UM8ozN/f0cROlQCYg+03/LPUdkWQMcpILys8clPor8Rcx
Bwiwd9Tb/tgZY/IhDoxITvdFQBOB61HsYi9Y4OIKfVTvFzSZgpPDo07dtgRuL2nc
mZq6Eh5BHr2QsjFx7KwrKP2vve2tGkPjDu4RBDM0KCAy46+/XGGd7SZuUnrGSZHb
85qa754iGeATMQkzdwN539XEtCvYONngDExr1ehYpheHH/c/9cKiZ6tVey4WRrWU
ahbs4xMG+00iWs+4Xy755fqsFgtUE4dwGif/s06/CBCoR0XPQGqyphzM9Ja1klfP
sdMLmaKpiryi9jQsxLx6uvemcW9mWAtyA/OMGUkPPiCtKhptZfOFS5mGxwTQrE77
gI457YewW4nqvEqdpHZv4Jgz13G4gTFcxkLXx1mw3Ot9x/astqg/7rV0zsjIia9n
T2B4B83kOdGVCUXtDHRYh2Kt4W7DHhmV57iwUGNR+fmuEXDoNWHlYZeYmNcVztcV
nJjoxG0wiLOcIFY8/y4B/QbAG47+SLRmdmddiVv1WxnOflllv9OlDrQZ4XdyBLY8
Yoi3LmkgKz2L0MvxsHxg37zPvYs8xWsvwHhiEP1vEGnzsv7mwt+LtB9l2CljkANE
aGVbcCCzwGFzccdpSEO+qbB1uJnyrj2jdWV/4eKoRjMuC+leFZQ06tMDXPXjQoyE
GFtU2VY0GJ//cjvOxuPZLoFWa6s9GNkLsEDMQsJ79xIYeCMgmhacmee/w/WL0Xnw
gPw8a2hqjWaAMY1k9lP6myxXav9oPehDVqEILsHmn4F6Q+IIe7YP9hY3Sx6ICffz
3eB/E0HJ5R+YMFeOH/QExo/qlVvcrz/2iAEv1dkX5b9iY7t+Jx/EBGGImJcVtwCr
OrKvsJlQcyAN49syI0l5s4DdNWWC5d+V9PwJ9Ey4PZwBAPYxIC6a2fQ0ytjTuYPB
FM9RQNWT4kmGl9XMp05RJmaUPmRjR2j9ShIns3phgC74sdCv7+WM/YzuGifX23Xj
QgbYrogKEJLoQSTehiSBn4GuDAhSJWan3wU29/TEhOMS4AYPWTb2uyCkU+9vuhJr
VTY1hrpYwCdM4vshsKbXmbw5vANfDIFBU1GFDKj4VJ/Fmjm/Lp1I8u0s48eNb8p3
xFXAnI0g9xxabf7t76FASZ0mHYElcIVCK1Q1yuPPyRK35d3V+/e8BzkP6eFYGdqC
mOmEdwG7d5jWXnCzNhuTv/szFYUXPE1NsaJUV+2Fy3z9OGJHB59UTai042guOKnn
/FeGUFRY1j597Y2DVin/l7DcVBfqRmH+LxAlN8XAml1ExSLdPi7zieqa9GEqbGev
ssbJ9+4dpn6KoDmxvqmZHQu0dASTpINnzQ/LYO/JsNa0gaG2P/F6U+mFWo8sxckP
8o7jLnXBbDN7MpQnHWU0GJH5xa+9rzvVcavSjmO0VxyoKFITs35meeoLnEaosjQW
AhOaDs1sOgqW4UJcirLL7wNbaxcXAtRKm1EM+QYDrW5PcikovNm43LbC6rT+CGlb
zmtFr8oHd1iuYD/P9GYeh4Tv8xD2XlaMtijyz6k4LeMRAg80M5oKMA5KbCkAAtSA
z5JS4idDPJ1M8L8k81VDuhQzRm+94Na83L6/7iZw1o1+PkJyppODYO1OyzckY/cJ
BcbgbTtI6q5Z2Vwovn9bOlJd1YcbD0DPSoH/F5LpTkAVp5Q46/OUZBMRQAVzcfML
6dWM3wXdanE512ysWOi1MZoSytsCd2tTEPFvUVIQUc8Ey/QzEEAemQeJEWTJh0OR
xcuFlUrVrP7nPHq+aHKRU7rn5t/QBfKqGBsLLRcgt4lu7o/fikWXqRgUdxOFVnPz
R/1Bw7prnzzDwvCZkmHqciR+e/ETykD3gOfdrL9qadfNcQuTyxhda8jj9ezQsu5M
OBQzkKEGR+3N0cZeCEL6cVikNk6VJDFaHbjHp13nfnDZLdIoMiyiCVDP5Pxqo/vs
w64l7O5y9xyeyHBEqqp17CnEfWVrZJsTyIkheRacBOixY6RUGc+2V9hnXhSdS83a
Drldvm1m5HhP90MNlyGHYC8aN08TxY2b6f6CFmRYHIVgdzFy/485Mo+m5p2WJ7Op
glTno0H47GksU4Ew6jKaQTifGPkFSZchKTXRwBYmGb88U8lYT6Qgz9T0bq0AAcNb
qRSaKSDBq3k/Lw+Jx43KRUbXLrj5hUeKcLTa2/7j18T3HNRs5kQU5dTC19MuA+Y9
6BTnXLpk36jQrCPEQLQY9jBnb2sj9qDGm09++2H8xrgvzdBNCnA2ck4TZHRBNEHr
HqEgSVArViwxPPhdebL0z0PD9atVJrjGLZq9nyv5j5KklChMzKYHA7FOazOpKPqz
yJb2+GbPsEflD0gWVzJrBsX2AhxaXVEiTa4QURfAB8FRnX8eq9d3sUDWgsUDeH4d
6PCMxPn5z09ufizzm+qIth3EGs/IVwHdIzW2yAVQWLE8h3tI8+uLCDETT14k4Cqk
PBIsMw4xvthCq72WZluEVAurnyF5KPG0qXBZdHPjAMhh9lmKeFdeFpPHtQFDLs+k
qggBlSJ+tQwkQYQELgBzb7++WPm/H0q5goIIZvsHgUQZsRoYPhHVZz5Xr5qG+GDg
KrxaNtK0BWG1wlZ3ZsQQhrJxtwMNvbuA1QS7IwwyAaNmEAFnIOjO39g8Nv7HSpLH
sdNIWUfQMF4ewJ/Nm22AUlSgPA1rgLWBRJyLAzTskrlZ0P5Ry1nlhBPrGwAxEuG2
2rYfxtPsLrCvP+p78nVEjy/8j1cNvf4WVRGZUcTvCL1fjMbqePxhIb3KdC5tDlXO
nF24F6uydLoYsLDZba1FtagiORi22N8bKeyPL8/aYVUUjIan2L8RtA2+DOIE1J+z
2aR2adeSJ+lWImqGHbRhekhbwqPfBpluaxrIwJMD2o/FvAhH9bMV/zW2drXmWkX7
tjENr94lJX9ykhvUQeLgIHItJaNyOKHacLEbwMEjiVBrrIX2WvfetpuqY9Ax3YW7
JIEn12wJUVcCRY+5fksyjqUnYJBQHVzD1BJmphzePBGMZUn36594+Hs2NpCyYckK
f654l3Xbmp7dDaJnVNW3EAHuMelEcJIN8B1luzDOz0XIWiaTablebxSFYHCCOqdi
zArdlZEEmeakI6mWYlktKV36qt6SCq/Vp063+vE9qoTARhpMpRhUkHLPzwxLF5D5
VAG0obj7OPzRHbM7kPB+1H1gd1oUqFaSSOCs71ILBwwL6hrx09etzwyOmi4YHTQ6
lW+ukuy42HQGiTnQjBqQFjOHkKUP10ML3j/l3lHZXMUxxRvZWViivvKlJK6LRt4C
TfOKI/Nnxt1BKxMLAt+05mEHGGcGKiEWM83r2B9sLYRzdura4NjRB4Xkz/UFcZbw
7WQle/84bjY9NJw+1gF8QhHTQcoa+FaPVG0wz1IyTxvHrwJBvB1bTBt/SNjB4MCd
kW+vH/sQr/Qd8zWsqWv4C7PSHaJZzEoRYL63fCCwhzZ/RLiAaOhhIqaEry8ozGpl
dNvb1eKqHZ8/FfZTol2RzKdOjgKhInMtqrIW69vJ0ug3H61gUWHWpucs3pyooLJK
ZpqqdfMhLpClSh9I4aMat9GOHXb0mv/aMB3TPupCKIpXCdHLcQF2fj3/t/a/6+4v
geHqJCvx6eZ8NZ/MMFuYQ9hDQBkKpcRcUFjRT6bjNMQNziT8q57KgEfcnVjri5vu
/jckFCAAyjrY5iS5GmDx+8OkGKUU2qSHfod2pQfFQlB6yNGnHhLVb22lK2ncOLs3
9+JRye7qtQrGuQenHs93XDTmYJX4NyUz0h6r98EcyifeOioAgklNgb2i1BGa2/N7
/p6mEjLBCbpijWio8MD1KuVDIbrYFt9wR/YRgBoNVJrPwyJ3K6z+sQYJoN0/rOTr
7Bof4g2x0rZHrb8IMr++RTQcEzxPUQnaq93HAKldpAldl5BArwsP6PO8a/fI7qiO
GhY4ho1fC5KxlUqQEkpYHimTbJ/xibmJrmStCS9hp6QXvaUoiC1/hlsv5RkTMsBc
kWAIWgWebu737odRJ1PP3bACeH8OHvUivfo1uaCdDLVIW9Jb1Xvi41q7xyoV+DSe
BV5KN/Z0DBOSS3KrNvi0ZlbNvjPfdlxRTt/B4dmUKsUNlAoNap8SD5PZTvDr3UoE
R9tayxgW0Ug3T4YuPHjefKPr/A4YC20CjcdH8+v0lfMT6RjPH7uA/nUGJSPAwIj1
C/9gnVWSPB9185SG8LX/EHTtPYirwIk6M06iohkwEzz1d/N4edfQa+5X8/VTd4vW
KuD8Niu9aOasAO9JHYWn+VJim9hNZYpQMTjza3eedy0WNq0VDoL/9hVvWP6oP5D9
kC6IORpb0xYfo/3oJ34s5JSQiz8GKPmhFopq6xwJT3/EUR2TXqBU0iTKQZJ7fSb6
0ZXV3R2P0aFh/9zzYhyglKsSPHDFeXcgR0FHf/M2Vc36WrQvvjCjnxVHAbQbkMWD
q0J58ZK+3dHOZliQZdcuTZhDCVMFdK7WN+x1T/vRa3qRiKkBmjwvB5mkowWwtw48
6wnryrgEmtWd5wcB9K3Odcj6tNH4MYXYjFsRkTPPtCofxj1y9Ta0mrUNwKl1Lp03
sIIMebreVa72rD2FWRaXkcMF5EuLnY/Sdx5T5dXh9Cu0jlP8HCv8uxHGanJza9rY
sw1GYoa05k2QN5mfu6gUzg4q50ZfcNh0xDPz7a5zcQDp3Vyy4N5dXwzgIUAy5l1w
a6UL85NFqFvxKMBUnk2PTGctN+61VcUJeRv0AHY9w6Iuq/DyH8TyGR67piKTXOKf
9kL9aFpwr9S6VpLfmyNVwCOhAVyboqUDG6Iv2osyQvR/sAEfOF6tg2ucU7ryYY99
GFUzeQ3Bw+qvXgKcPsGuJtDyLTCexl85QYMMSmoBerdvYNRj8cfhrJWsVm+04gbL
bdtS2MqnXS3ynVgoI/n64tErHzHmbUIZlOF6LwF56wZmhZFXGRLAgN6UbX3Ojr9r
Oo2xpOEuyIxITIgTveJ4rNlkBgdOwRKM4HVtjl6tfEfUQ3nhERwA7WnO9NW0Aupb
9xLXuzaelKxHaNHa/Oy49uce0L4tCUN2JNkxf/vTl2/AsmUQxpWpnODlLO53XRot
w9CrYxBqMK6jfZV05C65+VDkwXojAZG7ijI8eGQUZFXKEoW451Uh5Q8GJ8JPBer0
BmOZ+0BqQFPTxne8/ZL8Uph96IJYlPOyquY3uf2LaQBdJs8lg87dIPw1ae8W98/2
CN15UvBDVJfakAl1wGKKB4b4K9+oyb7qqxklKu7eor/muJhwkJq4m7z5dfKyAn6H
ITXQVBcVna9zpPXjaDUz0tGDK9Q+EyoUXd4acCNluLrGDCPD8XXiRTVFySxMFOhu
wjrRxViVAsV58X3tcKHeQLZmB2OOPe0pw/OxF0oN8dKi2eSunZnEWS7olqoMQ7DN
98RAGl6bBoMpiYHVybwIbioNQ0J1aooDQeRqMxV00y0feVbCjnUzfcf1Zm7Ufkf9
LqeX4vfT845VSaM+4XKS+8db8t2jHGrwEt+QdWYEuDBOrWrmALVm1ovgHEGHy+Pr
lcDsF2YVejt/hrhnyAHqOJ03ar53Z82kYEHJEgcwMfk/nr/i+5qUljrENXIO2wn1
Lx1oxUSNL1g7ICcslNKvoRDQU+ve7cfOVhmjeLSOFmoSx9M68M69ocuqOLgoqVFe
aQzOkhXB9h8+we3hvSZeQqlvP6G+FPMjgH7hVnVOL+cQiqurybYYbn+9kMhx+14I
nC8zDeY3ZA+7QU+XSn4nOVbjegNpbGzVqrvtTNuZBI6DMouSue5fZj4o1ap/hFTY
o4IgGATnjESAKThP1APXjCVNpIjfFDiCxewrOVV8/1ykGEKTPWSO+fFjqeSDbq0R
gS/KKNZ1yImMaWU5etIML3Fd7AViGIlq8l7/fDyn4CNa4c4ufcoqK7I9mp5ToHey
gFgrFbItG/nCtXGycfPi3M0/URmcrkM9DxHZSPI3RN+2YAyr9Ho7yzRBGjVXRaPd
D2IA3BWXvNZMowhTajrxV0iXN9IWlCzkDU/fKK6MaAh05UlkC6FNrm6U6+LIz06u
GbiydduLitFFxmJ+9cln04bBnSjzrPUQWNpSk8dYBr5sAVYcBhHJr8jF1FL++Snu
+tRY+XLhtQ25Wpo1U0SeImaiBikSa4sai3TWx7gZ2z97qE+xy/s4pY1LXzqfnZ4z
EajX96fzfZKc5LK8Njn1KHk+hVKPTvpTEn1Nhl9Yhsv3JYzXyrJsYMpDWqZIVzPf
hvsVzK+TxP5ib5Xj/0B36TDeVQ4owPmGBnaTUB7lGDhdbjVQ4/jNoWI8quH52/TD
3EmoCjHOcb2ZGsqSpJzyseQ8EuX8OThYniSdfYuVmH+q2WzGUULDX6j0lQpLVfvh
ABK72TsAU9LcRFE0PQ+qp5wvbiCY6htvJ6DFmb7sYARxr8mLK6XXoOIKsJq1LVFl
6pXkELXaecMB+gbn12MPW8Beu5806RX6G9XeTDkeEKXhUwvGN0btJEKOTeH156Ap
dr/Q1gmPbz/yi13UWVGms9AbH35W1E8ObLRuX7Do3IxMogscGxS2s/zt99GkaQ56
bR9DjaMSol9xnDJ/wJJeixvImZy92AK85DD20/7lPxJSwu9Rh5bsYS1MACGcAX2z
Ds8slgY1PIZyHx5PWSvdJxPInvkYzO0JzdE2vFQnjssQi3f7T3/M6soGMeyuv+F5
EbdgI2pwJg5kVYMN5nLVIiv2Kg6nfXIfzr3amUvNhzdvvdRGKpbpIbUWWNTHBINm
ODFPtJ7OugzRUqzPvgOfju+Pr4auFx62DWv79BFE6OrptyRZ5NFuTk5hYVpgGuVa
J4z94OOL1U5BxxrfUYuJuWRy+8054Km9Ck1WlrlsJZddtB1PHrcMt5/NStIneCuT
u9x4en0CbOrq+A8w3s2o48BQDndeHEqCnJy9dQt6WqxGzbNxRMwBoptcN6YHDBJA
KJSujjrzBIK2MixJwRefqVh5Gg3w078PrqAi7ln39x7z7gffuIGAkWBQmWaHAzXA
GkSvlICCWO6gLbieiQXs2z64wDC1znjcBM+8dA/V5NJeFaqfyIjQrCmCqAymQWLF
GOkbAQpCl70xmcPzdqnZ4YuG6R5DYHWG+setTuEAvyqrrp+E0Z2ltZdjJEgZvBNI
lrTre6hOYGKeoNm4bbgtZef+pXoHVyLgNr+ncXUWJG3lUjxGKohSMSIphrLzPjuj
T6TkaJxOAlYG8Y+ss3NVTJcFwE4ilHQyQ04FhqXdjHnxUPvQ9SiehUlIaixaMTvv
UvH+BXqTOkbQ2IyKuPtHxQWpYHjyEJ02X62gMgO7mDXETAqfadPkL5WnukHzs6Af
gRJZ4xJXcpRf2Ag4dtT/ZQIdEUTEmtB9BrckHXRToV0M1AuN86v8Z5+v73KajgvQ
geCu8TKJ48mD4sF3G+NBHKJxjVSSm6flRsOTiatebp7VO7qCuYv3pZu0YqPOJEa3
6sANvV9fwMOFg9WGYlj9ZhfnNaz4rA9/u5EUr4O6NrFok/+5PUp+XCBCiCrEHCSv
dUx2mUrJJat4KDl4ifFw7iBx041zgY0vXLkruZgc8ctK5g505GPvodBl3nLGACtQ
vKkzIO5TM8jiF1WAb7V1aIux5AsiIcUVmJRdUEMoS7EIz6CcnOypJ67jjwCaeS0m
9iPZeIlWjO2UNIzLN3lnkhq34qd9QDZFkiYW+uLhRbAQCMOOlgqvHm9EkH+7poqP
IO12s6dGqD3aa4S3qkEEE6xWXDCxhLOx4RNZd0gk5x00yYxZdLNYMxOrE59VqU5b
blPSQd8+1UjQ2I2Sc8zoUe3qQH2IG2FOETxAN15rca2Fhf/jxAJINm//p03bvRuK
DtNfX73m1ZC1dxPwu2NhTMyNZluBhAxAQ2qqU6Ck1Pp5C4vJnDGlLQfyCS08Aj5V
SJo69190N6vInVeZNe09SNLyG6TQzxXmzxDXJcI2BvRAoTv+CbHIC005jDLVep3K
JLdqFJ9osAPuwjyv527QqqjzCJ3KuASWVMHoilSGArxErXI3UqhEbgdDxfP9VA4J
ji5E10YUhS/qNBt1I59U5PQtza854WoSnCbc8g7s9g+Xq4rsUfHU15cVE/52Xl/n
TIaO/j9xLlOL6N4caxje4lUUWhB8A+KQaRRkXl6yXUA098urdH9JDhu246XkgxAj
nNrRf3cKtKVv1tfxHE2HQ3eRn1NGjBhG1JeCMV113dSebgftqxrUzcxe+fxcJ+an
g41lgjQFXP46Wm8gsNR14l+1FS9JOYqVgQfLXn9aOxWaMRdMV33D5ZW31JH99dGH
IJ9sybzMt2j6vFp2rRNL4XqIzyWokIHb6Uu/fhjKuGY0jp0hXSxzMQ03UxMs2Brs
f/3kVFthdppXgJYD5STEv+tzwcfIvcWVirWpP34S69/zDaQI/ti5w2tBu5A+9z2U
MCytifTtp3dfExe5Q1bkyCThoKI/WN6LRBj0soy+MNRpNaR+rxGlidaElwfW1NXv
Mb+/yuXkmKdOUXs8x9XXXFMkZKLdJChlck0+GZ2ELnFVhpv6II/mZojys+21ASyD
oXT+rQFPRV7RbJXI2ih7fGPZMOt6/nohjyKHuKgyV0mMV4qnq+uL2cGIhn11GA5M
ExblYbq4qkW2A2D0s1jYrUyA4+S5XgU7mAY7LrkklLQwAZJ942axHO3YO8QhIMPj
/AfirABBImKQwtbAjvxBzwsUQYUuBAM8xTROHQRaI7dHBh+Rppk807MfQGstfH/8
VyhpVHXrXX8UojjetMtpDxl/0z92n4ZcLXhXvxszhtxBVqx0rbKl9dHwyHkrCeFD
v8JChOOH036vDAz9bqalElaW0pXPN3x8e5A8uy23V3V2cfpiFmsTLGyPnL9jEnQc
RTuiO8DJXmZCZtygS+IWo31cP+Oikrgw9HR0UpLOJM9Iy3EGiSS6X7ukp2gLUMqd
4eTLv//aI4V1DHZk527xcKcoBjdCGO8gVXopoRYgc3bboHPdWU1pGCgnpazW4/2l
+o3cDFnAQi7i8GVSdQaxWOKMTen/Jj4GYMVgwoUrznSWhAudw+GWo4Jcym3Hugz7
Z+Aiei+1sOGJK1FHgBRIfouzTUQFObzj4KuyzOSv2sIytE24GbJq4kkoAFui3SfD
l7pA+bY53PAjyeo+8gHV0Bzah3KsckZ2wLSaknOART5m+lLVXsW+8psI0rWGzAgt
QZs5BaDkO4fvxqbzAqlZoAUqO3Z0A1ePR8qt0UV7oAYP+OKPvD9TcMZ/O9NQEQgg
Ati/2jumfoc/ejgo3sgNR9sAzV5C3K309d3tTf/p5oKsqi99EMdCwkUoAYtmau72
rljFeAQPXpb7dY0zMPloW/3XrGgjZFtOkIcdSXNV8T1KNolzzFn/1mqfl3Sia2tW
XR+QU0AGzL+0S02sz/hlKz1n6kiye1Mqd6xsxIppZtIZ1mSW+Bql6zlBedPwPKc8
wO9bdFqLccSpWCAQfhHiROq1kCwdZMTyIdya8r7fRt8BCiUOl6nKVu1EnXM14GRZ
fNvTy1IcCom9FiYj1ZWkmiTxJXe2SCpOnuPW1I7YxImoiq/LexoOGnSSPfbgXhJF
8oRIhm+ahehEue6ZgBw8G4JE3D1ee4Cbxw6owmK7PNX1X48AGwy0ca+oZXHTYUEK
/1syPejghkOyLVcDHyfVIGSQz5tBMUwoTjVMMw4pnulL0dDLlPWU1MdxW6DTs8MG
ttNA/RhuuaGaq2035RVtt2cNtHO9uwrxvZC5QQcbUWwHUVbpnYPlukINk6aYUhBB
2WHqJbW9j8wnyZvqJFfNa4iX9BkBEF41wPKfSjbA9YjBfEk2DxpXHZr3Uiy1dNa5
zbPnWD9GdC4nNRWW74Id5VocGlKnFghhyUipvO3/2hWUSE9rNWGurIsMmHYtkph9
Dbw9N83ig38eMbJC4Nk6fyI0KnSmLb+JUVbnBB+J2v1PsDh4dboSxPCXuDxwPIOI
dpcl8+k22cjGYmmUTfySWdKvM4adtcG7Ph1ohoWZKmdt38Lk2aYJwVpgk7PWd6K1
QJR3QRvug7wty/m6ureSouAc+AxuR33HIW4q8Q2JusnRIMIWrBgldGfDppmQqhtH
UcqmFE/ChsfPbBt7CqbCEjrGL1b+QRSDzsyCXHx8pv2hcC94SZ+BMiXSj5++1eTr
tO5Jhr/16rgNXku73RgmwlqYJxR30/G3/yKGs8j0wHNGcNKbt5Cf1piMPZX0bJ8L
ILRfOz9w7SChOMG9nY+fx8IGGMnL8yQETZ/JEDx/wyI0/WfPeNbvTt2B2tJy5qMw
CAmpY+ZmeXzcPZuSGnxsjGjGwsoaw7StsxwPBIWLsoEgwibsZeNz+KmArfuhGOn9
3LA8mQ9NOWxOUbh+zy3v0fRmc11LI08JF5BqU6I/oHxz5/Q7IIaI2Nbg9DfPBYXP
tApSfbJSFIkbAcDi5iLAlhFjRAnwWXN5MuhFPFIaZjGymwWRbo6M4PXi70HKAz28
0ZounIgSq9acj9YlCpII/wY5R2fHgPtrGxdmUfLjQ0FYBsDXotAKrcydEhlVeYZO
DoMZmJyt7xNuWp7aLJc1CgjvzcGv2rVM30Mq8Evn5caqC3HuQnq8ajkwN9726ai4
YY3na/ASfZlozZs6XyJRhUtQrWlCTsmzT1Vc4KaZ2AlGkoQqkAvmGixuL9oe+q8R
4fd0IV4ytEBDiDCPhUChF5GSoGlVN88XA5qm7CsvivkvHsS0hfi2CzpRwki++xAz
yTMtdYkTfPheCT6FYD4fN0MCfAK1YeLEPE5139FREOVBxsTnPoVNTydJD6yiWcQq
5FrujuYjAtR633H9fWgb9PORwtF4SZ+cyRyAsP+ctlOYD3w0VOOMhfxcbOZz3Gx9
KiOdHHMQaBL5Kygixe0LHvQFW6xw5q9JJeuw08qnut2Te454R3Q1Z/Y2/JeLERyY
0kYZO0qqb8dBxEwZkKlv5+pfYyEFy6nCjsXZ0OBRxHHKKPhOmG7zCb3UkTnful06
fE1gqJymPHJjo4WfdXhH1NaGkmkJELNZsc/JM0LP9LJCIjMPSnQcitSe2LNwuUVt
nmuYiNsbHya6C9vsCP7DAdQ8oxKUazA3lMxwbxDJSvR9uBR2eUVvYI4yS4TIgUNN
Yiw3U8nBjGcNUTVaSOiNE8SF70UP6Rm+obwY+ypBt0db3HutVMWKL/RciH0whozu
gVFO8JvVyQRSsGoFftjPFwqhZLWod2/AOvnDZFxBgO1oTtZQC6NYpf5kvxPGYdvk
/ciDx/pVK30CnXSJ9rPFOb0AHH/Vh0Yu/dGw6abKIw76brmhhkRJlyWWmwI7QFwS
8UD5OVrw3gXTYo5WLQDCM4b3hZ297+QfM17kDiajbBJEiC7PnzeQjfHNL8XxEVZk
Ljc3/mT9sMSrcbifenOX0XwHv/MKZjEPWKCEn8ZyK17DpVZvRs3aBbtoZySjQmgc
qlv4sBiKAOv6tTs7FcBYp3m/kCjaLpFV2aK1Gn6xx+Rcb4YiWXml3ZfVBUnol8Vb
WedKFV7NxiPqsqC9JRzj2lftaQfgn2qoIM220XPRg6aUUZtvezYeNuRyOffLm9YQ
QJmpnlSaAAvKKTNpBiU1fSpwSJ7ZryWGf5zeGblPkuPHjktvcDXmnnAMVsLgkK3K
777eZzBTGlGQnVNBpJ4JbCcWoS3Q5lswyL4RNTmp3d6dvsFYZ+LLVKFKepAAVNSs
riF6ERrdVuTMfVf9FxUf/vCT02HGuyC+b/95JrzDwS7x8T8I/0pCaiegCIdHK5SQ
CRIaDj0VP7qpVXBtZ5mqCI7cDCNtTS9MraWCQObOAuf4wHbyZfvTOh0MvLfmclmw
9JLXdT3MljvB6JS9jwe1JqtPeePYkIYYDNYpDmK+ItK9FzW6QELUX2yHQXLj6+ZF
N+VvRrYmHtbqLJbzAS3XoNH+9WS8PLIKp9s7QIbTt530J51PhK5y6YuQZG1D4zWI
MmxRIaJESIzc8WWGb9x4jqH4P9xE81m0ZBEbrwRtEeI2tgTjt221aUn64QtaxweH
NQYd5/UnOTl5eKr4VjCn2SYbWBg5qHDveoaMYaObKkcor1+KQBw7f5O6IgHxfCJe
nLQc8DlDTdnS7zzW8TBHjFxiMk01YXlFxkLdoJ4qGnFasSaKl8OvFc5e9O47WmAO
2I/DawNbTpAxX5lQjxbCnAHNP+R4+4H8iPdgkedLVy2TqaGwxnHGL6luNVCcrilN
dQG9qLEacyLhldV7quNUnpYePhCdyVA//HAMfXrPVQFZ/AwnScV+hjynGTRikgMB
hjMkQTyOG4fowdtiKy5jVPYSJkQTNwi5vUO2/V4uxRxizp55lGmWynPUAATXZtvi
YxuS9TLC5QqAhVuyZXBOlgaFljDAATBoRhQ9QHLpEx514EEvYGLbV12ffcM5KGmI
iM5k4/nRof+GhXWmafAqwBnfbf96jMIBfLlXkcYB2kbt32wrRd8+MBg3W1YZSrtr
sWJoj9Ehck1ut3j4a0OeCnM467VmrcogXLYnRBJY6IaGlRyobYS33gixOc9inhti
FwAQ/61KmNJY5vwuoHTCFqsteeHvAS3xv9htI8HPxqHhqNKVtOdyZgLwiBbrDMTX
9334F20wpwEDkM/JVH7Wp/e5YMdkao+iPm6GAMkacXOKkttWf4KIvWBmeFuydRP7
QQ/e91sRHrKShSgn/iiLhcv6YvM58lxjMjbMsqXw/TJ00sLEESk5E2W/0I8Wx0KR
aVjxfD5ATEQSYSFtE8CZATLrKF2x6boFZT3V43QwU2rZjLAvQs8vgNgO7QeSxAIy
QQ3R/RRhOw7FHhcg3mRfFhTyGMatXB9rzMsfn+0DQYie6FgtDtEwXVF8WXrKlWx7
PX4vPlQPeIWm8vZkUrPWutlDZ9y4ulaMvXvXNYhuu/+C2w6ROOAmS1UI84t7qgIH
ES6yNuYx1T836VAtrVzk2jk2A8+fwrtsiEBke+G1XUz7GlzD3+VFyRAOVDnGIQPj
cH1x3phz0Toz+iMg+CtZxA1AcVX87PYF0GDhIb0l+QrXZ+tmySpR2HTmTMFEF9YG
95tiIk/YCKsso02vu+U68ulCAvRBXG4WeEhy55yakgehRq0dFdMxUblELDXwzlhr
QLU+xURhBEFtMcy4DVSkWCLRXRRns6EqDONU1tvTxOQrPqd/g5FiLrdR0pTz5r9i
qyFHMlvcDpywOQ5fQaIdUX/qu7LOnVDyPxc9STprILdFF5JIm+LMDwZ87QkKrNaF
DvBXaqW/Nd5RermBf9lZWwzn9/srEO2Brlu3mEFIRhmbxpsxE7v/HkkIh82ozUSI
ewhQYo6aMrn0RBYgpOxvWkUq/kMMPwIShbem89UBsXuBF7Gvk0/IrfWP1Lp3ZN+t
iI9p7zxHrQmymmtbHQjTKjI4NVf0OgklrDDhN1o81QKSEznfEf98R/lIWlfNPQiO
+ZrBLH1xBhONRs4LSzLkyU5mY/1eWxEwNQR9POM1RsTl1NT7LMp50N516BboqTdW
dGTUkDDSEK1cwOGd0NUBexK+qFr9dbphcde9j4cl4b8uiFkmEXo51vVcPZIdMXzV
yS/YEol1bwyuV9kD3rf0MHZSSgwQ0klU0Jg4R61AX4fZ+n0czUfuL0S3voDjc5ya
u8hrg6R8dM4VZ/HYheTlu3NLt2A+33S9U7WmX/JLI04PpoDjOhUKLUWJkZzRpoNa
keCaR07TnYH1AMZv+BqmfDWaTCLTYLoLlXgclM8A1mg+/d4Xr+BWkqOfU90xxl7S
wdp1+PFvW49l4cHgucPe0obeT0qN8iyDT7RTZkxvbsPtHpHr3WCkU6Fku2jhHzIM
u+ZXFLkLEOCrC8dbiaEKzEl2IodnwYimYgMTlPk5j2aKuFaDcZsufu8dA8WIejhQ
WTvewkUTySP/N07QBpK05bSG1qVsmCWMbOBwhxfmOfm7HutHHXZrjt6INMAcrdXk
CWTeXIxHLcsW9ROx27B5wnAzkyFrylr4TI8PrXuw0AeCw1d1z0KMIzqdoIU7zWXl
7dS71OqLqIVnlrItg2kjsz5VQ6YyuPduE8LTVQmoCYimufYNWWR2DcIsCHl/ujJ9
brdzmcpZlVz0+MyjnDH+xg6sRNu/JrF1pVQCRF8ZBUnP6mdApOFUdVMM3Jwur7Vl
Am9wBfzQzQyciG5Gvp8zMi72J5jYNtneka9FVAc8rSZj0/X1RUWnkvlzniv5lkt2
vj8EBfjc2B1suYMYTAFTGrwdwRoBdMtAduvBrNKUbNuDhz9UZS0a3dlteiOOBueH
QM3r8QAQxOGfyRQmfshhgj1JuZcG+aE6E6fLU2llf0aAQ7ZMDTm9Wnrk4uwtmoAW
m415pk2yQMNJYUc7HpGCw9gB03kNoTyMuPB5oeLBMcap5po6wdSuBbRRZi6jcgfh
7UxnOTtOBcJ1/wT5KtBcIbcCGKisbMa1ktqDtD6OOCW3+seLOaSaypeBaCp36DhD
5nKi1aMfi+n0CUlzOJ/PQF3/N8s9XzWPPiMUYi9fZ3U7WpiLEVmBXCacs18RPYiW
1QksBAHksEm7OrGJdQu5Xb14RbTkBCypj6ZfocW9iYmCVHP690SFXU2YOjpL+t56
1RBrq3aNa5xul70eYBjZCJfetdtKnKjbWFXStUuhg1XJpY1IYky38AYEwKMnyXbQ
tgnoEfH/GUlzLitdBCuWmq0FwvVc/xSMao1QDc+TYlBpdy8ly66dD6cX0ey3YJh7
8UcANHC8e6Vduw/GZj/2xaeyEpo2UJX/QsYtlGRtonLLlZ8J6VDzb+Dq2mICeXRs
HZnW9vZf2l1TKcdUOAoDuw5tjwUGTCK2Dzi6b6Y7tm1iT0PrBcayzOfvV1lDMxMf
+VbnObCISBCqUJ4hoarxKH8X4+xxhd402dDmR6ou3L4PDaqrQd+RVGFvP6pbivWw
xkuVR7t1i/MuhKQ0rstRs2ojA327idnXdwoAknD286tMH5uKsW6TGLzZpx9M07i6
ygHua97X1Wsaoe40YQW6QNLo+HjLtXJaDvHXBB3JsR4hwjfswd+6ZU7bcqe7EDqK
xw/2E/e0cqrPCsINCABN7L2h6O6v87tEpeQvduA/cXisjbcJuVIIfSQmeVEG2kOX
qjnwSk9TooD8szW/PkU7gdTRZfYx35cdZaohQRNFDiY5AsZTslz1AlavW2D7UALX
ffYqQCXJ13mg00sx/pLN52Ao03s/roaW5T+VQjwG1Pu1vBxtHXDC8sYOEU47IMeW
vta/WH82jhatgjzZNrF8fuva115jPbUyVtGub7gImjrT2owD8thDEl5mc+UCwGix
YBVtqfB2Bx9NDqH3WipIW8rTMpwFBHntC3uVDH0P3N+m3n4+gvLj6VzSyUBFscO2
RHD2f+iwKa2S5jbwypUWgiVnKnk55gxfhv2J6t8ZMa8gO8ojzPGL6uC79LEd5g1a
3h6kUDvBmxmBktelp7FWQFZ0EOEwxn+kVBRRu9IFohnW3hveQjOp/jKdE6wUHu73
Qxr5WdDaCNDYQ2BjHVimtehAvFu+K3VCFiU5Jez2r3IJQNPv27yy6n/5sp8lSsZ1
s2sdPOcFn4iWO8VAJXmOcU5NBwWyOxY1jQKdC4MU3IsFbHxS6T8czbjPGWrdxEGn
yVcU8k5V0yjheGSHG5DGLuQMP+vy7s1a+iPhSY3hbeyBMcD6PAHZzUGtKwOp4qcM
ggZNaRdUgi1kcOefN4M/+5/X8GzCHZ2+8O1Bw8u2/5lezXlOQEe2kjQiBPbeGY1x
3npPmvdy0GEpVKfdRUAG3T7J4oj5kxPW1qAC7JyJTMpzdip45s1Dax53Ef96DaWF
JYqGBRawB9loQVLD2o2QLDj1mC+F4aUxWqOeprF1G04xDKT+cz2Ntt0Oqwlq4X02
zDz1ZjijSuWRHHjqKUGIzqd2oekNZZUr1Yy3/oCn8botLVONQGY7PICE4N1jhGOG
ZE5ux3ZaZuExOuon4IZ0AFhUOUciHlBbWB7kKkrjIkMSbQ+nEa6KrYXW+/BMFfKb
Gmt85EkCxHTDuZuXdlJCKA84IkdkEAsePlXDgHesl1zPRQjqnHTxAijroezJmE3h
5aJXaG7CN5NrOC9EGR/HAKWE4x2tYG0XABkMYMJwwhjrkfYbqypCAq8TKL+HpXXX
PvDmteFaBF2Ksq49UN3J8m+Hfx7v26A85EKj4lJH6sugUSAa72JbVdeZong0teu8
MwWPd3lmNAvEHVIBU5nj6vDN0rbWIgvAYT+YEZMI4OGedGy7Q++rmwNmaUj3d6cS
JeBEECjQty6ablZVa+/K512R68acwEFon0u8WdB8Ztm+AO8REXuSVb6TGyaNj4W3
afVIXFVTOTRTYdQUGLk25qX/CyTW2I+UY+5JWajVpC3GbuGE9yM/AbJOjYYN4RP3
KNIOMLYfz7+X70ID3cdJ1zgyVhpxhloDpuuQixEOTyAOkLvJKSeSX/93SSuL71KK
O4qk6sW7difZo3Yj6ItypDXpZTJ+EQt2rneLoLfaX9IlAsPus/xJhjdYVM8MapaG
Ar8qsZ5Qz4crmZ6jRenTSNfAveeiksWOdO0idr0F+B+fE03vZfDcrMvmk4YNAPC2
5o4nT4uaXkdwHXIsRhtV1W61+uUV4rA6PBLw2VSQsfD2mz0w3KJRzIApN0XwkL1U
hoHN2o+p0DUoz4a5joD+OFAuEk8AdwQuztFFrBdRAO0yhnWjl11KlSAK/o3MKx5h
pgXr2WZOHPJgyCcKvfnN5DmQVwX9BbTyVYIq8gy8h/oNTXQJ56BDmeVn2QH+p96I
cidpsBLfjTSZhPoOirwIa6cUV/lbbYgXEeRs3G9CsRxn2yO4jwv/sgeet7hKs+l2
g7Mq8i3eW0XwpTpokbx5GYzssp2Q8DHHnJ76DXBhN76jH3MefGSaII+PwIbavwtS
lBhn+d/wgywrA+asJc0VCI7sYKglfp7/WjyC7GBdOi5lqpw0ig0o/D2D4QLXCYTL
3HO3Bvx//sDL3Ay0RCtJ4TMtD9ty5aE4oTHN12rbVDV73ymq8Q7TzQsFCAzC2Evf
dekNe48d03VkunaoUNrnhfIuetuyzB9Q6/2X8tTjSkDeQM92k8p5/XXhu24rHBtj
wEguAaHyCXpypxpCCUbggGkK8Ml8C9LeInpRB8Ax9/w1Y/Se5eKQ8V6NgYEafsng
hENKcZgr122rb4b70utjmVDS5DjZjxvPliBZyeITG9pAjziwV9M3xaTsYDO+E8gz
Eyd5L76S2JZHhRCdN0iPx/PhyplHH6tk+uA9nehyeeEli4EHqO8sbzrg+f5QY0dy
i4lIbZw6BRq8O/SfS77mWFdEjFv0Cr3fZZDBYySpzBn9SwiWPKio0+y3ixqwgOR/
/NLJYsQB/yTOoHIbU9LA5OVd9WGPSvPXmwkovbsSkq2mZZhovR1aIB9zNxbE7lKH
YVbl9M3EIlpBwuQ+Mks4c3wyEW027DUAiQtyFkkPDiwItY3c8fJDyg1CyFu7RhQe
qJVyDa80zE5UqsvdFs1EW6RJqv8Ov2EqNMWKp0fp0vwUsl0JhT2A94+QhUbeZZqD
73/7lXjJb9P1hn5nnLZG/wBMRrBEACFaUWoLEVzAfpV7Cpnlak/BF/eExQlxYGQY
R8hUktzTR5ivd/7eYd2WCoc5Oi3G1roWMMcwLEVYtM0YlZ2dywk0KpjaVYE6wz4X
UJmGO5YL8BLkrZBhUXAZQb4E62b0AxqqfTxSYR0r46KIzFfzIsKDWqsEcXxpC+LG
mbe6n6430VqnO1nzJlL825lTOI4LnEFrNEvOl4uxfpHosYgxE0VG4EOqNj5R6fRR
M1P1fG10I05KbdmzjT6UzlgS2gQ+gxmCIB78VBVTrBi+L0QSvtP2it/7j6bliRWA
4jUBxfSLsOGVTld7kbUpNv1nyzbJNMYnyhfctRXQZXkE9GytFDZzpJfQzq/7HcYj
ks09zK2RzHU3AAswRlbNm3+iRx0eFj2t1bDF7pLa6kchWjLgjgCv9q31CREsFzxA
2FoiFzkZoS4AzvEvx7Q9O5f1Nrx2Rgd6AHdGkQwCnzP8HrLXeD5YOvq3e1jwUA34
ZXgJOA47lKTwaBEmQ3iVYMTHFC7PdWiPcDvAepzc8k5SdkOsWWt4OO4pZQzgF3vF
fupB18gU7LOUBS5noOZ6h1imEs+NT57niDnLz2laUhuvqsrM1nCeOtfSb26A0utO
rlRrkv9D18qdk92+Vh5n3PwgXrA6+Y0ZycpIMzS212D65PD9+txVNJMGsXN6kNZ8
mzIwg96U8Qaahb8HQQcENCI6EMeOF8FbYnPI9bF1r2f/rXtriUZXFp/VK6MtL5iF
Em6KNFw3tUOJmz60Diz/O94Gh7UsH11g+h8pWqJCWpPuvGu45/xkQydT/NgftvdI
mN8VjeAwSYbPSISpmUEkj1qq3ar75H7uP8i3shZi3NI8jsPoVHAEpAzffkio4D2A
cPQ0SQpXifoxDYWVoYJhJfghX4WTc+Qc3lX2Ok6xytVYis8qctGxp0iH3/s1zjpu
tyVg/w2EGKoPFsgd93MgOnpXH+vVSkv3dh1BMt3VRGL62rVLId3b3+GiXcFFBooa
v5/usXSXy9UU8o6DhWxuo4ZrT+jy5Y04GwHVVfYRHe8okxFgvULl6+4S0fdANA71
jryQLLGsB18F6LaOpx79u/jwd8ckeF89ouJybWimo/8o8PZw7QRZZZw8GV5KaMUX
afYeOC0psM3J2U2pSilvcFfGxhwxo8ftqEFRVHpA+yPHZRN3Ucn5CuctxxTwpwzH
125Wrg8W6WnN7xsB/BsSLWcQc7h8N5thX8Tbe3fGyYs62vrKpZh2iuAwb/zOQ7yr
qVFsjWtXKfEwaFL4huQ03UXlc+LCUKrBSPPfBbeuVFICx7XVyyqHOyQZqBNcx8cj
ckNlU/XMktCyvT8IaHyPNgdlHIH3jzHabYq+wYGahyg9EN5Gsk40ZgoYHxUvnrND
mE3A448v0Gur+KzXliA+o47yAbo594XuX01moYeWuvoYffILsaa8HV02/GJ/vAtJ
9PT8FDpPyBSXr3FsN2Oi1Iy9AJhTCf3Py7F4qFz69pMDPFu6oZx6g9iAy0ejfnff
rAOQfxuDcP8g0O+6kIbrOBWhEOP27MqcHO5WSfFotAhDEA3FcQ3tlX5HcnDfrHvm
pQXnb9zK9Lcf+pq1MBaHlzjZ+G1wzNY+3X5v5kNL6zxZceXHhgmyPKG+lEn8YojO
pzRMBciP+VUOqbvsOqtrE/aLSo5RrOJxqPVr3CuUsmL65LAjkz5fOBIEJhJW3lhy
sOBujs/+yt8AuChaOJBFPprxF/e8GuLv7TpZbL1ue4oUPEx4WDYaYHazfkvcTOhQ
+bUybUQJ+yBAAZD2OXsC+I/Sy3SVnPXghcXOP1yV2aYk/GlFZRClTi6Xzi/3XFYj
AyXu0x8JU1DwGVi73ioeSIaZW5vn2NTU4kf9qCwx62p5wXFzieEcnNn1Y2Nb5fNu
5RD8pnR29txy1CnTODa7fl8r3gScwQ+47x6YEK4e2/UtxIFakfqbKhs8rbn6a2q7
x2Ptd2mX9rqq3z8mQF8VAqrJNzwAv6JgWw6/yiVNdPjDkGq1YJlNasspr0BYnEuE
fkePtcLCin4+ua/AMR/zyM4vUcJu5UkVDaHe6FzKZuWFIaLtdGD65SSHVeT1htp7
1JC73Y52BoJDbooKqjqSYOwKV8XVT7+gvKwbI1RkJeO96BPeUg+kyYUBjgLfRZWn
f3ZEeuhHobo6n6N0udHzKVEQcxXAzCWwyIGL4xBprUIeidio0yHBvz29eIUi3oTS
BuAd1AS6iHo71wtclBLNKP9fHgiD14mdDf9WVAQC47Cp1do9wVaS7a4zuW00f56p
OTs9lZFFEKD6i+bBWGxLVBXmDjpWlnbTKrXECBR6YsMHcVxsTq8MRZGlpWkDlOJP
6cM/YpWcrYbv9WC82Qh6Cvs/hNU4lMbgxbJ+2cvSUHq/k1/SLtZTsVXZE5tZzqMx
jz2Os/8IuKEyyKreGQsqKRUT7JwOfBDhNCbBwHbf97Hwuxfaz7hyfEaTXFW+//A/
UHNfNgHcCCnqNPjc6QkZAQQcZ78ZvDgHCa6dfqI68GsbWW92o66X0LVmh4FlnnNF
EC2DnlvBLnQQDtGDlwH+Qw8msc7fo3RFIPC9QK3ZiAn1cs0kqV++AN8I/8ekJfM7
kjffZA70Ct9CRnhk4ckQlO4pqX+/S0BGtAv35HG67/oUygrQKdeZj4HVqim7Xb5z
1p00zjd/vbx+ZDSO3hPwUwRahflEh0d/Gbq2Sh97i/JJTh8evlHYlWyAxuL5+WRl
tBdcWweEG0xd4Zl/stfVjxoMJq5aZ0S2hAf7pAkjP9bvjt9F93JTlXI5tEdMTLB9
e6iUeoZ3cvo/wStzQJDPL+JH0ZmNj3qn35EjIGDV3FBgBh1PCMqMRAhjQ8hi7u5h
+Qpa58vHFqEjERl+efOqm0kDLPlXlX9fOOavDx1zspkEgVqjc/f3uAqjfPAeBvCg
S5GrdKiXiS1rFSxcl6MLY63IfzpU1oVqn97GkqtcYDBRs2t+tAzEDk4rK+qGHhHb
uPuR4b2hVKLEN0OKDp7bSMxPx7hG5dJgdxrQIiQxARXPzS+MTIdtEjeiAx0Yi14D
oaZ3abCtT3TQELZoObS9Fgnf1E6rUmKw+u/9HGu7faWGMoffe+lkKGUgPO+YjjON
APlpo6cD1PkpXvDgKoCwvi+xQYAifTUZ35mS0gnL4X2Tdod/o18Ev+kFj+5Bs4yP
1zgwv+UIkh/jRr+uvOTDH5YmiA6BeVd7xL5962fw57NMkhwkmc/7rOepLP3G5n0b
iFnPf8o/6nbnNIWu84YeZHPuCX+1U5n45hm7m/DVF/o4fAloZZsieh5mPGfS4+g/
HcDk5T9LZQZfcevUfqqgmuxkyqv3K4wheGSCpVqoEdZzdqAg+58Zi/k8Pxwf5G7g
KXDkYZ4hs9ZhOp/vKcQ+449zJykcN643gmvFgMgwKI0l0mPBkdHrkDJz9QgFa6tM
yMiAEWxwoGyG3jfl/NRuJDHk5wtgH1b+s8pogNmUZ8NgKzMsIrDp+5D1o4fdcP5d
KBepXc1Je4o18d5CLV4A9A0m6dZXJVjIat/uga8GeV3Mk1aX4A8TM4LwhNKM3x1J
FxL8Yq8YTA1DHg52EF/QA4gOouv5BFB0PK8F/fmy9R5aPU/iA/wL0UH4w3bgG6m4
Wy4y5Z0dj3b9Myrshp/GbrOe06Sb0mFFADZLGtBxPVPWeRQlB1AbkNvAvnCHzMG+
5bHRlE+7tALZMke2ZXl0fFeIj+4Tqj/Ji/E/tq08XmH4YaulSrgM9Mxj8jFIL8qd
Dl9dxOhPozfUws+IfNRJGQGXJInvzQVq8xYGsPWLpqYJxZS+ihC374z3MYwusnfV
godq5JeU6QYman7v5H7BzxQCwSbrRz8XSnsELPtlNEmkcjeWFxTkuMUHzxLvhWQz
xDyHQuABw8KtTkuQW23EpcJnCjDwmfB15WX6dU+XroQKk+F4D/wzxq6xHrkQnYmu
U92TbMm8gt7g0zfANzvsU2gutDTPFg9J2lX3Nt/j1329iAtkfTOfOj80ZGC4SRhI
dGzdcXn0CR1yq2HoWkHEjdNDdWSGK5lyc4Cy2fR+5YCKFtaGhznlwssMms5/MMuv
ukBFRpPqcVa47DcE6fCtdmsnEsAnuuKvJ7NhNqO9ESm2sa8J3Y0SC2WTpTDD6yH/
YfFfO1Q449IP9eyIC0k8XOQCbrP4EvTopOrHKWzlBwkRuNl0UBRGUO2Cgp0ECR+v
yRUeR8YJnUM2z6jpssYzVkHmn8pHELLTz3jg+/V/prrzaCt9fbTjU32diHz69DUz
A7NZh9I+CInWkDxY9aeemrvsGy5B/zPUxZRSp5nuwan3cqFqajyThiN8M/5UKCA+
giSLIgjhxzQ40BxdFb81S07huZ2awTMOval/Baj3eu1XsV4WJjDBhfFTz5jmsNJ5
qj6qL8F7ZDqy3y36aYuRmUoXCZwM20WohO7s44Ls96wu7kiZidVzxkufr8r6T1zJ
8CNlFNOf8wJeeSnbnFy5vXLtBcbNCigBfkY4TuvtlFyRFdiJ2IT0wMfPczpg2czj
fzv/Lok51zYLA3+mGr0bRRx72b2GJP7BvbpFLa2BD+HlsGh3/j5KYnAmD0LgdeDS
Vwz2mu+VQyuy/CMlG9JepSbzcMCHsGO00qLevGpIaBDgHrw/HTLjc2n8G6FDb428
dzPHvXUDKhBrKISeRdHpzBB5r8Z1kzJkN2RlUJJhfoD0W6Uj34+sAVIfQUM5YFg1
09URNH7uiR6hagJ847+2Hpl03BJUbf7KgUVn/tGxcNatXfU6tEIBSucQ8mwC4v89
9tQPVr7wmAYdUtsMwl4RsMjg4U+bzsXqR3Hx/ICdTUpMu62xffUeTk7NOdQ58AQn
CQJKNtrTh0bg+w+UN20TwbDb9e+89p76gX7OfpDmm1dPZxoJO5V6tYmCHF+/QheD
F92p0fLFHNzzrnIstavi91qSaaE+B9eLFw2BZHd5IcF2ueqXa8lI1AMb2UtP9XzQ
BVk/Kb2hmHmVaRxME86zm44IwZIubF21gJqSKvFS+sM4fHjhXssbUQy3SDs/f2N0
cE4DJi9qMG89e84yqMlsm45zoEwz2JoP1CgYs+H7XTMpFAgPQYSRFY1gMad4WTGP
vY6D60ToBXfky3oIo+nxHDLUqPFPgHxL3vr0zn/nlrt+Gc7YF/gry3KzbD2l579h
/i6a6tqUFlnI95L858fba+dOrYc0xiAQFXOKqmafftfjym0sDd/YmS0ASJeo0Zzw
M/Y8odFcbd1JbeJl2cyUeJaPyvvxayISEOLRI3thIOum9Yvf4VC+OS5EctJ5wLd/
hLjx1ycfrHh68RFQ4dZQ+dt4Q+jlIvostwS3Dv82o4uENfbAPpWkvkjsz1m3Pl8M
SE3qiR1Y4wk/OMEJfdXCNGQXzGLWrLqiRA6MWqmd4Y2LirYuA6YeL+hhQbiQGgAM
jFGmbtPpuXPZwu1bHphyLffO6VkUC1cnGGHD/HFefZqELZqJ1jY5nG69gSo1Hr3L
w8wh3kmm4GToNj9qpeT9lBpXgYn0MZ+vVKPrAbgM4dN/lc59OcAzfkcNbPlGmFSz
FMZrXYbUih0pLUCeQYOHeaTTCmAn4geBmQl/jfU5703ZGzHyV+UWbJ1B0IgfRvsO
AW91DQ8Rp7t5vQ456at6SvtQf5Sl/qPeIoKyJGKKv56Df5R/NmwfscQH0cqFKeQf
qWvjTvr9tlw0cxdHg6jB1YroC2Qt9SkiTfwtKBbOM/095OsIRvhowOgF7ZqDdheF
k6nB5gM7vR77J0ezJ+HEHZBadySmrR3IfSHkm5RxVsSTPN9VSWazMQl7XfjnPeAL
roqKuBjsZtZirus9iDQcb6I6NtVSeKLEOjHuBMgNQEeav1WCLewsSbJVoTkbq+55
MmqS1mRCiSv7UAVCT3H05JaQ6YciODLql/t2GNRRpEPvUjMZhOi1DA5Toz03jdA3
DvAeKQ3gue2PGOhMTqoNOTTYSIr2EAOdnfXvfVJtL6lEe8Xem2RCwAUYPb93trDC
RYFof4cEUsuHDSHzjqqRxXBnvB2F3kX/P81nYqBNJq7LhliHVLlTxBLa0iXF0lSr
aaktFatJ4X2/Sfml328Ng9e9mgK69nj1mTv92Jg1zBoOf1GffiXsujXRRAYYgt3z
Dh95TR31/U64lzM/9XvBx42wGIvFWn1ejDtDYP8Jck7r6hw0pnNCSLXJEWeRiYv8
iB6vh71iHmwhazTUxopxahQnnXsDiqpOdvjlLYB0fdcBTTpTkFCL8dzEZvaTQLND
pag/Pxry/czQdQpcJCf8EzmGNcCYOb4m88t6lAYBPxCdHesNk75bH22leqs7JIXF
waxgdALpcCfqWlyoID5FJHulAqsHQJEVhY4HKyEhjFEIuu7cwN4iol2a0cepDO2r
zzRKG14yoN2nOFtLHkUg3cYoa9Yv3e6SMnNuxYCdkO7oVOtddnGLevYP6/uVzBPn
WcmxmqeCIpbjR2va1o7Mr0eKdjWPq00BEN3cTfpkB5Iiy1MkEFjP15ZaoGnomvut
ZMuPn7ndUgt6YscD40SURF6Ah6nZNt++gKLaK2cUMRUJoWdDMehmvBhqnoUCG2uT
uhx3eQws1lP1M/Cw872IYfCxq8Nfj9+5FkjWvZDZjnjEKY7HhXhP2RoQ6DorzHaH
M/ncpHrzt71wfoVmLXsnbZsBSB02VNFQCQdHnVQlMBzQ++PTp8as3dhjB6D0cSc2
wEJyEY9HQsB0FYrBqBzcPQ4oHoBCKPjF0c2b+BziQg5h1FummrjQr+Vgp0Fxx51R
sdBQjgyixI9ONRGDSoA9fcAyf8O08sneRel5ayO/6nbFXaYce9rkM57/lGjIcaEO
OEUbswfcTVUJghbCSOi7JLgkU5oErzutL2508DhOfETm+isYzFBBI44fyZjTujF1
zOCwq59gKBi4SGGOsgimMtZB78GtXHSQFz8u5VdNAfA4Elpf8/Uu+Ih4/RtIDeMI
uyEmkY0TzeNnEUScInwPuFM+0EUbAwki04zHrMvni/62p9+Q9NxxnpWR8kf0rkn1
yAmfqxioN0mPaOuKdvs9jsZNSZqEYWadK06dKGSyBwwnf0zoZqSLyGYiaig7iNT8
PLh3K4KpT66SVEGkCBKh92Iga0E6wVWhKFP43M6oBj4p5hhguZbJVYf5E4O8JbOi
5jbBoKpFF5kpKgAQyWFN89768VO/fin1EXA7QoU/SfhFy8/mTu2WiUJqp+bH5UQI
Zyo7snwla8KSk94e/k4DrgPHKquwasMkcajJkcz8yqY3+cpH2QwxkT8vAc0DlR73
e6db/MDicS2sluq1hi4jvI3RvFWduqrWIgKvo5UJ8xcYGu+ce3HEghd5wC4UiC3P
EKonmP0F4mHgOHx0XG11EDXZGFxJdfaeVmFELGYgBOY0QJLYtk8KEC6/VAk/2NcC
v1XnBZb8WBmStEGucy4Wo9HQpWqGD/i6tukWm3bSkccPNr8yNH2p5dQJhmlw0kXM
eW6OnL5EgLF2vZD/ycXihd1JqZxxN/HFxcz91Zi+Ra0FRwviRC+H0mHw388h4QN/
1d7PdX6zxz0wYUVrVZeK0BA0HBWxMLTzLlTsxq+4V8+8xX4KrOqp2tUt+uIeezcN
oG/oa7WSvQ/2uIMMKHm9/ojblJgAfiB1lwyxCe82AomnHFIxJukKXv6uUo4PmXn9
2f/fKBBm+0iDE0thes4Pt21NTzP93K3kytdqTRgpkpiJwalNQCpQBI2e+7p0gM0J
rGx6svELiAAP1nHXWYund99o+XA4UJsngqIuBt1Amf8y1JJDZ2qXAiQS8ZFUq4Ew
uWE9cf9lKzoeKGNLtCF1Of9Dr1a/eN1nBmHpz4TMXIO7yTw/KxShr0EaIOyKh2Ob
Hwdbi3GY78nMusXrgj6zcfmXXF9e2UsWJOpPMmNxv8KJGx13XWk0Sl/FPecFPwUZ
RBsG9L9Yl8zdoZlJCUq++o7xJ4yATc9DCIF4NWZH+UtcKBd3fzHlyYGINPyRMYgN
IDgLkdv2yF9oyfpg+0cC0tjJyKwgdfO3zxMe9Ycph3VfEJIanaBoNcaaD2qzXk6Z
4qkBeU4CdDL/50uYqZ5aaeNjTO+ckd7aJmKlGH8aJd20MOJUnKgEDzTwTUyWapWT
71+7ECIQlxJ7xGFxMNBhbRup45x+S7B5pPiZWqEwWVgJH6uN0R4QQlUJTHcE3/Ks
9uLFFOJU1sfcfpEUvGGtTpwk85FOTVCRPJsl9yXLGe7q93xQq2E2r2YtTP1XIglV
uNmultEo+TJ6PJCsePK32Ph6shVXSmEb9/NmaFX+/hH4Dsh+TCGIkGMdw/pF6fZj
Ws8AFk0jA/yBZGFivNBqUPhpcwEkIl79hgefhmS+MNK+ZvHQKlV3HKGFci7p5+ZZ
Q1cHAx0Ut18ZoFw7vghvDqmDeVKwKBHeRJD/bEVmif9/oIM/HXuaW1d40eQKV9sI
QvkZSopU8jKnlujwDYoTJUxToQQMu2TjwAqV7kp6/DEElQGsUdNZ+WyGHtQxo8JL
cKu2YaR7iptB9T2RRwt/R7zi1Eyjob9IBFtdZwiEZ2cl3Q2KESdyqLA32p89aqTg
mPvRRJPVVSRjpG3BfvU57SD9A9AMx2bad/99Oan/nkrA86KKH6rqRIp6kTtbwYOn
XjkPKuqbwanX2oLm6d5lIgi9zrSRaE7snlvW4BZrCLkQiSKtOrtW63Lj/+IU3WF6
W0KQSJaB8R/bbxqPzeFprgCjsDtpb+CEOgypuM3clcNGGAb+fkPN0P9CLU50BE8O
AKtqOkZT2e+E8FUpAE2llTTVDDOAOjt9pQiSIjNHXZWqUXM+DiFGTxzACuKlc7Ji
C/6OJwtySNUELQZ54Dt1764jFVcZjlh4Tjas+F1oXZX/BeygbOqiDCrgXeuhiTQC
AFiZGf5zVHMTzi/acXpbbNtIC2JQJ3z+I2bgJ8wuZIIX4bMNmT/8uPLRzch/MnCq
SFLag55lJTNR7ilwwXWGL1u8gtCUz0XkC9gfczOemgB0uap9ZwbCWAir0CBHsret
/f56knjrvF7pt2xgTR5UENC8KHNkQN4nUZRidMKRQFIO5Gb8TP0D+g4pBjxKSNFJ
CNRU2KOpju5wBSQ4aeYk22czCeqNdcshh0HbdSltaHWLqww5Sns6R28dPQu2ZUl4
H+h36baoFkUHhNluy4lOdqV9uEAQj6z1YL/cGjHBXSVQwnVcgNei/nxTkIrX1VUR
kSWK2MdXM15a/ZT+fwc9/09grwx+ePPdeuh2IHrXU1kVxZc2aw+TYLweytlxGHqR
V3zlKoXofLv8V8a47NPCBC48xv08yga/Kzo4jUmeuaiODDasXTc9nMKQ+eXVAs5f
hsjH4cl9JjQCCc8kvV3AyJQt9sk/M59KxcLfp5lve65obukDM7bhPvsTjBoFIufT
5W2EhZz+dXMlTW+/IxRO/UYhfJeWuAkpQjnUnPgerR6oGI4X4kvbaWYSiZi07nNm
d1Hpl5yzPomv8XGuXM/EJ77aTdgsojtQxwAAgNnfGFziHyhZnuMFhqmiAwVbo2yk
1+KYQDvYMe4uqg3LWoxHzI1heuookASJWW2v58tYkItRNfZca82aDlgzWQXi34z9
G31cG1+usWQJnEaCQPBMxH0nP/DPR4uzKTj9yaeV9bCULOAC6Ou3dhnVieeulkPD
TWv3Fb16fADabttdqZtO2mHPn7MR01dPYMEAE/Ya6Ouot063hsRoI1iMs4/N0UiM
XHq450pxiKygb6MUgL1EyzIX3lQW5APXnBIyjohGXZ6ywFL+2ww/4fGCvY/28qaU
LsBivJKL75xx+fCv4R/P0eV41n7sJfY1shhqzdoafiw/HLrpyhRa2N2pGqz0k/sS
7qS9+lHoqkVAesgenhC6TiMqHQkOloJ66i5Yp+RX6cf1hAV6TZmQUtN7aQgIb3lV
xGEmDlMnHJi48lc37ULAzbzagnUW72NRrexfWnNPUSkH/H3Iib2/RQ6vhvYPl6el
QGGS/mk+nFv6hyNo8dyRaHBZMwEKhrDe71g05fkpd0fVnk7Nf/11hP1bCLe0wTn7
Tb383vGtlxgs2cUK+67394eS6N5W2SirHQSF7IN1F4omTBbBv3/PJsHbVOE3qCl2
Sf4Z6h3uZvvMLgLhw44j8Y/o7UQV3fzIR6QKBxqXQIVw18jJnYIUneveGqfbWDzl
R2U7rfzjz/sn+Z3SHk7q88D30pgIiMx8NUeFF+cO3qF4I0Mh+o/bGbjfTRmIqPGx
DZ0sdpVT5dMqndUUMd9E08i+PkxHl+BirnNXbJyv9zTw6xbA8Dx1MDWWHtJBE/C8
Vo3j17jrPX8OzQtBSUhwhGcK2q0kylMmu97MJhYDt4HRtY7Q74LbyrakMbU1Dx8g
hIQhucCzAkkCbttFM/zoTe0ES+vxpM3MIqBUxgpUKouCrYLVWtqIZChava/1A3U6
c7dPoGPOWwUu+knQ2JvhHfW7vcaj1Ve7PidXKYLphdvZWVxpoLSvnR1mNOo9O1Si
uUxnSKtZGbF6xSKlrGcnCDK5sPezRluMDBN9QvXXcVh2Z9bl2IVavfkYd4wDuJN1
7A2+aqtL9k4GxOQzAGkEON/TlrjbqOpJX/XZMBAZuENKejY+fN1xqVhZhtix1lVC
3Jf1RyJTla3APzIlx5oemjQbl/Ky/jfH4Yik6L8h7LsXaLfGMPePDabpV0i7j97M
SwchBEguQBjLwjb2hEvV8tEQZ1trLirPhrS8FYDyh6bHM6554ZWtXtbzoZupfjp2
DUsBH5ws11qmuYhlJMVgXtisP/6rZZQoJITwV4+pbrluySZ/40h+U7yHZc4sL7nk
Sj26YfPKJ2JusA64wiIVWR6L52Ce72EDgC+VAqpNyg7dO2P+reFBkPtUoFDorpHZ
yOOlVnIoM4Dv5Aph37AKXu9uAdi7BFpwmDshuno40rQnaUPOhaaNEKhJl4yyj+RP
8XCmkcf7EuuLlNu9+IQkB0WsB53F7up07/YcMnkQmHHj/0/gN9wuCZtv/AtQ87jK
pcqpgWGNeibtihwW5aEf+05smxt98qZyTwebC0yhFVn140MoXy263ALNrHAuVi3Z
sgAqFWuuPY4X7gEyVd9+5ObRDE4he20HUkjNiyTQt4KoOHYhGBnaUJBL83+g5+p9
6WaueE9+sHkDqUK1sm7WsHi7ljVmxoo5ZiyPf58lMPiuxwSObbpBhsIiU6Vuqs9q
YHZVKdJxwdCBl8BTpjdCYUkgxZkF/QX1gNQB+M9V5TVq8CWm14rQFeXv5L18xaku
VdgWKlmcn9KOXC8ZwHtcYQN4T1Ave8T2asWjaXxlSCDXf5KKv6vO9Ph5byAd7AM5
CYGzA0MUDyFqAqC9gODdm9NsBJtlXmaZIIS5zKY6Tm6NM3vt7ABTSnh56nxFij9D
oLOmntc44gyi8ldg1lvktMMtZPPoZJoL/Z5hFi1VtmyO/U6APrPkOpLWgH0pv8y8
cRCWH1j89sPJmP+JmB76uWhahYTlCH5bBRTAyv0YWyc/PgeN8qFuBdpppwSTm2Ow
+q1SG2bboqnraxTw9fBAfF8r/r8bcHl3IIOz58ue5oNKO0DvA+Vu+Lnvc5towH5I
FPS5KAvWPrDJ+XxCbQYsXHB/SnsKU8Zlydi7FoePCaH6Y9vW05o5789lnzfjYoq7
/iWF/AU556/b9h1NxaLgDDhX2kzA6pU16XeX1b6ilbwwwOfFgvugw9quQGDQuEPI
oXkw4AYfp9ahwoWN0c1LIU5f+F35Shwg/rxLYRGoalkS2KDP7p47SHj3KcWxMwmw
v9an/KL3R0NRXqWXtOwGbSO2Zteq3BDYugLZL7QUFvxVppGLYXkDCf8R+OlH58uZ
fHt/97IRDLd2C0GRtV+1JEDSS2g2I8UhDRE3MdexHrhFU6MUzgyNfwDpIYDnNME+
IqcHhqBQiL/4veM/tw8s31FJPPC27bM5bYh46vNaqmwdAYjmAbKApH1hx+UNcCPv
Ch04//u0YgMfqUJPnA7wlfxGi/VJlyIVGUa/9IdQnyReDfSDEb4jjGgWyXA4ML7x
iKKCnCIQ4EBwe0njfU1ke8onsiGkDoMBkpob7T0tP6rCOPkTYfr4zwxvtMZueXDA
dezsQ03FnJkCmc+XIWDHzcnUNMB0Dabdiba+N4afgsv7g2FoZvQRQoDDA8tSMkU0
exZqk1KizoRyGtDw6m0oLmR5CAt377EQlNPPBtYR5CSCaprmxjwsEYcXpjbXQf6f
gTGmY6jz9v1SxN6IjhWZZnAV9UnQkx2B20o0cFGmr0q57x8qp/bcBmJj/+FP8W8I
5OqE6RDMke8eNd24fImpHeoU6XL3O79x+vsTnJglgft69HJcuXJdO4aDqgTKwMx6
sLgeV+z4DyHOx75JYIg8kdoocpX88aqQ07rny9RDV88ocr+oaWgB27jfwrIIJQ/m
8Bbqxt0bTc+t0/CXz17s8Sd8iXRAI6TSMhmUwUIRCuuMxpe+sWdSU6i3gsOcGnM6
Ogr4ZqDhthC6RrWufMahZ6DM6Uo9qpMlRW+lBJrRbO666YTD2LYCNVQO8RF3mrVM
/6v4oJXGq9GrOjvpnYq39VcsSTxhxc6rCiSxry/1iwG3Ah6bYUbLyF/4jMlvmyBA
QnQiTMHlKbtgY1Z7tawL3iuCpvTHBmlycSOLu2a7AetrZ9ecg2R4d1dWijT9ZXF8
7YsTrVMpeokvpls7e9Yg+Zp+kgo/RRPs4PZkgbpFb4kf0sjU82tm2BmI4sx26E/W
/XqXojx6jRCEBEuz4tnmUBtEibg7dAXD59adDDczahZcdSaJ9tpivQ2cSp1jADoW
z/trItut91wEnIejFLr1hJqXl2iteVsfaSU97/Kj4yc+oS9LqODHYQT0fAohjOqS
0V12hGSjYzw8u5Qgmckq6MD3DcI0nCwOQfZNF198X24nJfeC9kiOLB3qjNNncMoa
g/mRe3JKKctYCxst9X6b445OKNyrufAiIpSFXxt3MpzJb6HzzYdPY4ixn6EOxwqk
OJT9TdkU3AitsgEX16wFbo1Wg+oPRpvXB+BIqsr8mKb2XEKABxhkfDJ331pYQPYN
FtK/oDv/gau1yXlq9LDFYukA8fEItfEqmT1MOeVngMYSG2tG/yvOFVa1xGytP7lR
zlf5aKSB4lJpm3+HHFNQXGYiaBd2CFbUlZ1U5wHY/aQe0oH0bJ95NFEODJpVx0n0
upJcLQrpRRVa25rOAKv9eQZVBWcktZLOeBqLvnwSfijZnK5fYaQ4QhE2aiQVBgYX
N2UEgI70wOGv8eQwL9jBG00B8mcGd15mGAE6fOn26xFbHhbeFxI2phEIRCzc952o
fF24SKpn0OJ8zcKilgSHjoW0GB0DRsv9+Rgahjh7BdrZhco0CMjbyu8AueXZDXE1
C8Yv5DUWIbx5/AeWCkyXnefI3sAi8SIQvn3IDskOYzp/BhM0OSrLmofya4gus8pI
r0TTEmPqYZ32NF3F8UBEoa+SoZfqzFuEPnCc+Qx0636exhjGs0rBrJhF6GwCenLx
QcQOIwW+tTFqbChWwbTVHt179g7eP+B0//yZcqWXLagAEx0g7Wrln/HG/jNHSwzo
Zq5YltWSKTAElqIZCxZRNMmEXqHs46LW7Gcg0bYdV/iseMibOY6AQWn9DGbSjDeZ
Hcy9EWX2vb4MCg7fmycRhGVA7QuYfC0SydhSlrhREa4OljciedAcvFojs2Y/FA1s
m1JW9wbPcIdNunNbjZTnk2BDtcwHSvgxB5Ak+AvILk5E3E7wVKhvLrn8GXa4hWqf
rwYqebpRf0IEa0Hy50knRW2JISJNYtBa3zTR9/AOmjJK1ziA/MSzmOxjD+x6dAW+
2KIrB1xh/KxkDI6vJFI26NLGY/GDSoK376ycLjMHUgwhoX6ZPLYW4M2yTQcBOZqm
jBy1yvyPFT1Mqko3bsOg486zaWsI3wPeJ3/KtXfpP0eVOa4DL4wV7SMihj0JO1pG
2DbGpaqu5InvIRrNnX1k0VnMRSmDIfGbQCm9SrUe14R+3LpdPfQ8kx7J5TQ+u1Wv
EuSwDwuN/wgWqZ0U7g19d8m9YAqWP7sIkJ1CN6iQYj0rctLKVgfYZXeqo0//CEx0
/lpK8VN2WKL4hYYvokh5bFBkBDF9jxylkpLBSvPQQMutLkHDkhLcO+1hC292ogMJ
gHdCUq0y9nPH2PQg/tF8fo4TSxASlNxFITSx5LOe8MQHFT+2uhR/qD3c1swT+jMi
H2iLsTTSFB3zgpIIIwED5ouw2Qc9GWfUuaX/98jnSyyFb51eTj3pHiszxpKuLy81
h4raspyExn+ENT3x1DuY+cy6h/kWG/pAZwSlMqTWbFKUn1y8hZ3OB277IFonVj1k
O6Ip5fJoWVpPutjRwCeyz4Rgzrtz9TgFp/XjKwmG74DRhaYum9KgnMmeJmaqZ6dG
JEbQBHaeogu4XZrKHdJ+ou5+xc3wqGoQ7EibyHwiuiic7aciTSDu59jDt3UQjcWs
GQLfgGgA21WNqABkcn0vnlW6bxq/s5MD7kkXsvlE7SCVSLi0ScGczhQNUoceyGG8
khb+O5dS4YPqFQivxjeYo/YCvi/q03sko5QTLbrZUZ/UESZJBB+i1haCCPhRJ3Vv
jjpuRp3M0km31YNXnutpyC1uHdIJYhIs+CGGCKNaICRj4C3G81NU1coj4hAWYqCs
+psEdJcuS2w3r3DePoL5Ffrq9JBWtSt0OJ0LOaJLuVs5aeoiPXi4CLK5Wk9Li16B
ZPRDNUmVJe2o6vDLtK792na//Z4oMRG/hbZz0D8FCOF9ATbWdHpFCvfAdiPsVDmW
CjeKbdDWO1J03WwWY6P1L91zeb9OAHSyZkqrG+ZVlYiGWFU6RVO/WRkqV/QmApNd
wZAcd8UFskR4MavLso68Jdv+dVsxgO1Ail0Av5CBRQn1oF07Ns18mOhe9qpwcZ3x
APZphFMp8JOe1syTc7HFW18ecMFti/8ZqyaVXPej+f7dWtTQvJVTc5+FejqBsYIi
Uthr1KCnuMDUfwKFEwdWhVktiTlSuCS78d9SU+ttT2r1Ep/KYlPDiGf96Wth6U8O
pvdj7u73XkTV7A+D4JiMyohEKvIEohsIokMhLALwoQSEE6vEoKdSUJWMyVgsWVje
ssTyfxMDh4n4YOOEMsFEGuYvJLRqwkxdr2Xe8aABoQgl/BvaA3G63qbTGEYcr/te
SqZTh9oUUn0DiRtmmRliGIG5hkCOWHjbOXJN9X8Zk7L/t5z0VzwLlwlLQZYZ4S0u
DgG/CksKUly0yhUigXP+QF6zt0zdEem3QF/3VerENDVCy2P0x7MaN1IIE94fnueP
NCRyKzsMugHswsk5M0gXNXDazObXoYEs1KxhujNLv6Q02Ih9ymPpoCPsEhTbHaIb
OHwXZxgXng6fcXRBfWScDLDh7kBaD2ti++Jag+I/uLixIAU3cT41WO5fgzX3R8OU
GAIXDsxaouxjOT+xSsplXgD7OLlHk/tV6e/mJD8cVtGkjbYjjjkzG5MH1JeORpy9
U1t8RpUFP/6j8JaGdeuhmKqLaV9qf5WGfBNDAZs/dbLL28yZ74QWdgaRCp58eZJH
C/NoXgy6zX+Tb1Miuw1gZv8ZFYVuz2pb4zbkYQuL0wauShXERS29crZyC/G2JLLh
9GAIPHDHwf8DzXiMW5DuEFs+6G58Nb0gS3+mWkrZcVYnKwsOfnpfhV4CdJTT+Vfc
xTwzCwX+Ctr9nKatCnacJyi6L30dfjFp9yNF7dWWe71/a35+xygSYDlziLxPbTe9
bPn6z0Wcu9i+Gw4kHMVABKaeL7tKbhXNDGUqePUItvWPi85qFtMEvLLjaUmPEjr7
XG3ZybGgh9SXVkY+BOD+3wN0LGLg3rMKkBEoEMmHTFu6CxmXAjM3Ymi9CjbNzkI8
GK4Gvqw6GwBiZFuU7jQFvY0KE01gD1nKwGhvh+uznxxVybgfVRaKeWORsH4uVZCG
U1EEZAQENwpxfe5Iiln8K+VR+eu/c6pP5wHm/W7qnP59AhlcJaEh07O+kmTopWcE
PRsAdbVwD62y+hLJYCHUDJGyKQnWuK66bhp48BuAkDQkWLLlTjdp/S8cd6vgS2z5
90FycAMtRMDkSfjTaNz6jcZDdf5u43WeuwXFFfpRjkoHQVRyYtLKEDuLN0qtbKOe
OJtNNNcDmiDShI8Yc/aYzoR2Po8RjAsiJtlpmj2mMpBYxAmQ04eGoKT4zTJ5VtVL
mP5oPBL7mSTmF1R9hIloBqOB+3DZCicAKrbgrM4tW6+pWHVaetd5bjy5SGBxYpMg
/1+L/nE+qNpdrevh301IFZFfBG0U3YqDyiy6YFfLbkw2HdQwAIEUbK/zRMkt1yOS
RevA5J8uFSBQ40lUpIS7viI4TMUE6hu6dCaBEPnjyNVoB3HlktLwK7bIACNc2Pv7
0eg3vS1x0PMNuaY+hen2mHjJFyfamraQRQsTPKOT1tvNSRpauHEZNXVyEyU9yyCy
Gki/GfvzGhKYRf/gtIW0g1Ae5sqAxNG1vYW2NiK9WbmG+l499JNCw8fer5rRxIbj
HDJfARQlIefmGEw0Vr3XWHVlXhKYXzZa0RfVJunDNLkcSMNkgFTumA4vDzKWdJd5
KbaJoz3mNH9F3pEEMUWF+Q2P7OWLZX7P2f2BZ5Unj8HwrzWb3Z/TfFOeLQYzG+EQ
eaHkSPOGDd8epXDrLbpjTXF+NPZsoBvazG/qekuDnPFx5vH+B5MFzh2hrnUHi3iG
+PN8M8hfAOkseK38jntg/IvLXeT+6sejXG4CUWr7AvN7ZNH/HvxoJ2QqPvV7SHyv
4SCRIVig+g+OW/awhRerokcvgnMP59103eoNPIQrtOS3L0JDdn90c/20i2w8D8nU
8WEPF1wHcGU6FxGpQS+cDr9pr/mrRbUUjJT87N4X6OSdfzn4Ang/yhrvIKjT2LGM
/H4Fio3LNlG4dLVK2P37zTEOVLaCwv2Zwc4N3l3k0maajcpR6lHLKrFwyNjwskqi
NACWbP6RHPrVRF+7NaelhNGLVKp+2nfKdpfI6ai8PmTLe66fUnQVJ0JDlUUkm4HH
dG4IjUJ+8azCOHcJFf6y0FzMIkq5dddVHA4wUvH9A2FhchlRs3NePWC8CJjUV79B
jIgutsDsQqE4m7abNb0bBaoXf9wWPvp1bR16mzdd63bZ+IfiSGS0vctHeUgb+SPU
pLZsJMMmGN2iMuK434enclOBNFfAv5122fW4Y/wH7f4yZGEWbqHR3PTlCirQs4Iw
uPDX4ZrTrqVMa9RZRylgM8UaPFdpvD2xnj2VGz0E8HqgHRlvZrjIvS6WEApRju5i
Nf+/rwT7qMEiA1KKM71SpvDySA7J5Y1tMAqp8LvbVtKu51dR2i5cAlp6GF8yMFPz
0rw36NQKgd/qAH0NKvRuGE4AeYeHluljxfzy9r4xnX7Ls9m/FnD1uxOf03h2jUBn
6LRqGE2BW5+HFiQtiat3PYFKwddtObTsePGCLrsAbWeqx1ORxRnDzK5NsHNQTHs6
ltgLjTr1vapXeUFkLJE6DXwGQo/fCPdxFA79yFTexD502ksoOfzIRoflcy4rznFU
foS0f9zODka3/5BC1f218li3bLWhUup4xD1oN7dy9xD/hlx44l0oK7pVtejc+GeB
glSnp4ti9xpYRCHyEZ6QwPcDD7pq2pw890jh9GmrYnF/VyN/7t1d/eS+mBXsOm0O
QzbVaYl3qBm8kIz0v7JgVHgViKSqym3xg7+4/96hpaMclGQSQn7kbjPFxzUP9Te4
Prd+F3ijYMKrJi1703Qo0WrKz4fKOUcfPPyXHV/QMT3X0KDCcZwRgbdbwBHlD3Ks
6nRz5sqoYDkgIGz4mUBl2zb8qfwvmVoOgyVvXitCeJKXQyD5I3QYpjxIQNky7pHI
9JB6JnsKMNac9VrMITBWLoeEX2YLZ2xyOfoudZE+LpyI8JeBkHgknPVimuert2qn
KkWsWpwTE50Gy2J2EK8Tj1hurnAWNYuxIsZazSHJX/Msgu1tcPDRgjHi1SWAo6z9
FUwFW5b07cgYpM+PU1a1mvbyFbOYDByPZnZl0CvPLjOdcxcm59asM9TPxrtNwapK
tgft5/i2Oo6dNtyyW0sow5WQU+908oPI+uzAYg7BDBnmlzdYmKtJwAuHEwCfegZq
iLEbmJo9G9sy58cBWAxRZsNocfU52rrcRE+5oHt+Yl9KZCGJ8ph+OfioL1C4dWu/
IKsA2qY0ZhJcubMPJFvaL8s59Wga0re3mEKKGIFS/C6o0TAAR5Ty+sG5E46xbjjH
7cQaQ5XNSqa3N4sRh/zVoQ/MnPXNUwRhIJrPZMf3yyBHmnM4keJWVjEWK9+I7JAK
OM8Y9bgkQSm3wzc7rBDv3HiwhlHkRe6SA0/D8jTLyTA8l7NpEEPbWO7/8ncrK/G/
Z5GrnfITwR151sIW9mXWu1uGcxW6DD5yq5S6km+r3Rn6/Ehp929b0aCji5DvFYNv
hhvsZ8ChYee4Qk0y83ObLQJzygyuThmx3R2inctvrGAw046FQxTVIdDwuygJ+WBE
zMmXv9MzQ25Nz1+kq9rXF2pFxNWA7sUPOoDdrkuEXnNkbYbyzq5tE1mGiBn5lXeF
qxQxlRf/XJvz7Oldyl2he7WORyWDwt5aF1sP0LypuvfmvCa+SFOraQN5ikrxslXM
dglZYrR/iZGI6rNfq+7d/VmqqNHmXJp15yYcPwMZjmGv+VEH4QwbsJYMfFiTXiHh
7P+NoTt3ewptbAV/NLc7wpEP4WTkdtn1CnTvDrw3H23j/+aMpv2oEQTvBil7wh2K
c+3+w5jSmfX2pqWj2Tqrnr7gB/lP3iN8aqUuf4YYWTNDZZWPv7TQ+fY1knA0y0Sw
fFG/sznWl91sGG6t8eRu5K1xpkz+wYwQhBENumK36k7H5x162t0MWt70DRBV2fTj
GFEk9DN06xr8cw8caujmL6d3k2rySLo05H5H91VOvYwYkJj60Bh/7i2MvYHIgAU7
2BN0FuVDAHNIfjIk+Caak2t9w8mFZijer8LbtTCvbvfwhg1uGrt8LjHL/ZcxdhRn
rb9jVh7xgEqdBuaTtmGnO/iwwb7qXbYNwy9vxvrlewGdD0/FCsUS2FBjIp8A30TL
l9LDkg4xzqjKa9gh/9aAX7RQfpvX3kDArCCF1X55UK09MHv6adJmUmp136Y5bPrC
if+phFqMaT24c1l68DRpJz14eQRGe2PgFiurQ3ti9wEK5/LREhmlj8TJEYsdysHi
j5NQwfxxjiyo3AwLf3Nd89YvvNkoToHI2rFYBVhLb4MNSfGpmWKeh3PSV3aXMJ+R
NiLC6YsGWFv8NvskgsoZ5suwBQahVvF/0LWDp7G3ipIYz93pLlquItwwmgyzWuyG
wh9lpArk7J8pes0ZOMtlwQZP6Bey1TNmLYeNUP2gFWe4WAFdU7UsUtgPF0fRLfh8
BGEbNZN42PRsG6NDjc2SQDk6diHPKnw4cSgWTVH0drb39mmOf27euUMvILtNwJdx
KyxixmgMQTRA3im4MQ34oFVyONJ4g9fVSW0NotHFni0vL9N/0eZikpBJhV76QDDW
DbC/gCj0kRhAg1P0zHNMD6UopEQa7o0KpyHRdM+71kZ+/nGpXErFAO6eE6Ing1Vz
Fmk+Ze9Fn8jSKXW0hC1ZHnLsGvKpIILcEVUR8368+y+DnbNrQEqLDw5yL9JXfzif
6EXbbtEKlMivLAAC80p18dSa6u56nvnbW9zeGjtff15X73DihtzqWkERnmXt6p36
t07vZSmtqzwokPIPsnxga1lY99vSf8+Ox80z4xvT3uMAH5/ej9/Qff3ba9ZRDFd7
WEYb6JmXL6SHkd+aYh0mTlY5vd4lKzLWCPsss/iz/tgK9Fhg3bR2tuhEfmGcpeV+
84wBfxsQ05xCKVFFv/kPBZjwcksRJg3wd5Q30qNxrKCxGLfbbAtRKnAJECo0uPgy
k08hgJnAkz2YVLIidEO9/BBd0cFXc7Cb+CJZY+FSi/iDivzL5d7olzxG0+rm3PF9
WbKnjE+l/fJyYp9zQjXVpLToC4rCbQCyeXcPVCZ04zIbHZWyqURMk/za7PdbmCpz
C/Uf5hRcYqoLMb5VHhwCv2PnD9N0lD9o1W+6rgc/DcJy3iUTysVwZgjyrDlp2cT8
ci0N6+AiScTMwquS75r3ncPJakvXkdq4j6aN/4FlA3BJwckk1lGmg3Skxdbk8sDG
Q4evHbhMeadY0QlX7IXQQWbHzmJShI5tqniN0jLSqtpnmz8FK2dyG2pk05vwzv3U
8T5QqVO0HyVozODEBq40acXgpbwROltZdfffZ1S67jnf6AwatMYwt2YFj1ejdmiS
XekHkv3H3kKtJxmgebXYpIkNk3vqo+zqEUqofB2lndnLXx3Ewryo7DX1aXzXdOyH
2fXeEKsai//5+cSUL9BL8HqbtPRbNzmkgydVk62LOAHIt+bBfvXW9wp6qpIi7o0K
FIh4h5bW0Ki5zsy50wORk+Lq9p17uew79qKH1USIgZKwCVGKPCXDdtwn7r8mtWKx
JynodPCvMMnrkWO7lZc8yyd9JiMhlFlzjEGgjpqdJzuPFKMahGVyJhR02V/FW3qO
TcTC5W/ad5u0UvNcfsloxkik63elU8lZaawwqvXg8/62+D6f/f6b8D6C2NxTLoKO
N5zDe0dOcqceJghJoiXtD+NaQHSdJc4umpuVhaNk1H6B4jclPycPC6a+KCH6pY0j
HfduuB1ZuMqZRpXz98nz0o7jfVHIxCt96wynhg0xJ9mV/8uSOHrwUCaxWmGBatY8
l8iZwonktX4csSN+wsIHkF3/OdScYyZgml/0ji+MvkCISEjGr8sOri+jEmJdHOS3
DSlIXlODaXOUxyEqU5e+Pg8fwl+09hiqk/iwskPcBaV8/LLoWFgfRciD1SY/TXfP
Ozvj9+QC1E3MxjfiiGkBzsc022GbqC+363qwuhikqStjTFGNf5KrYLWkbciJuXcP
yzttvPieSS2vu6vIMbRHv0QcS5woqheXshv7Ja3YGoymrfWqSzl/WDnOoVkicK6/
g8gDSlL1Mhoij2CE4zTsJFZ6hDmOM84X+RKNc01rlWfLl584GJ3aK9RhTmFAhQ4E
Cc/QPWPZu620kcj20POBVI2yrAA+YGqb9cEe48hlaT47A4gTjyaP35o4pmzAHlBR
eISeNoZjMRPSe1G3SQVTArs3stU0aVDDzjE2jvs0pkn3G/tErc2Kc8RCXkqBofMQ
OYwlDw4ISKgt1YGueSaZwD+Q9pDLWGE4bwkCWGb3Nyh23gmcIt86qzur43O2wLfY
hnfOKgGU61tvMWd3FvSszoqGUnjI+OkxGyKJ9PqUUpwd0i6AATjjLWw/Q2bj3eQ0
H8gTmjEikOcyzkx5vCNblZaMatmRzIlAuunXbT9959F5L87RqF+S4oSkzfijMIEr
rAb+a+m7CnFt0mKV9iIYvQSi9YhNYhE3Ko8yp3rbWloNwzmT+K9XEpSYf+KODHGG
0gnJd4BhfD78os64vKcbWNHCgub/38EWZ2JHJ1VAkzLc0pSCrhZ16wUU5D+/vaDf
+lKw3uFyl2YWLghj3++iFMpeOnMB21v7K+tpLwLKuhg4RDwrg3hpyNjwT7hdtVZg
bYAr/h8QVH0210LGVcOaZIl7yFXUUXoR/JfCtFIcOqjWh4vV5OhLTv4z6u9cA15k
QIbQtdCVxYHrmTumQv/u7y+iQy9+Qyix3FBLh1SD5Lslf6eRS2/okj7qFWEb0erh
V6AzcOq3jZRU5+M6IRsAQ8HNwFdMitaA6Bb2jLChA0GRNm7bBD85m263wZ0UQqrr
WrY5fcAnbcul80SHJXex5pYpFZ/7wilqd80uxyENoXoRXo5tSo/Is34/Krh8Jjiv
fe+SbV/URnEBDld34DJKlTKImWmz5mcyiisYR3Sal+jZbGEz1DSsVT48Mxf0i5Et
8BGsmjg3ThS7oWRu6tuqZ7oduiLw+mBmUFtx82YPBvc4lORpPlveWFn7LcH8xo94
aUYrTVMARFuSHPwVPI5C7r5RkOmb5imh+gUMuEk2OsOoqw2hH0tYeb3rwCIEfk6/
AJf3dvhXLJqwkNhYqK+w4/8gILIH9ntbymMqMcCtFs3ZNoiitmyob0IqhGELuXt1
075vUE+qYBGbmkWYhuxW1PE3Y5210WLfQ5RAlW4e9r2Ko4PDn8i44AN4TsIJMuhE
piANIzMKc6hAk1h3CXFLkfsE7ewI8+ODjoqqVztJm5XxRKfG57K61Qe/g8RCqxbE
YE7L15W9d2w6GvjS56kh62KZ1rP+bRUQZ0R2Jq/5etaaezfVcqiF+N0Qo/wyxSJd
XqG6UnHwvwXgmDF8map5Fa4udBASdSXbQbp87BQJI4uHBNtXAETKB0V/R+8Hqk34
vWaVbxJoYvJrfYxH+luERfu+XfBOVjb6udMGd2HJqTKIDT49bPUosDM1/H7CpM2M
E4xAfyuq7hbe3YVN4MNUcUYWPZaKh5k78KxWvjqTO3sNeikKZmoll+Kztht57syn
URnrFSZ48C7YSd0/tUySfO2KCUISX6CqKVNdUoMZ7DbVdGeGsuji102gKFzkK9je
1he8YJJDAHlacmTbvhQKtAo1NUY+DuEkNq7jU3LwB96Vo6QuDdH91TmxjTzZqpLy
UncBuvvQ9e/9Dy6KN6kzLHhGskChu1zCTEa/R0KV0kyQEilY973+wOGrY2hSwygV
o9Z44bGIi0jltYk3g9L82EildwnVuW4UhQertrqH4RSPUbqhBUYKrRT0Oe85r3uD
gj0CMNbzLdcMsQUUYOaO6JRAevLxJqagbT4R82j/YakO+PM7D0ZwX9BU7HVmIoga
LK8jV2hceXvyGmCUlBzspL5lo7mc8cs5GHRo8bMQ+DxoP1yptB6ttGcVX7xakYMa
MmN9YcnlAt5lPstmYdREaPRyhmK1DgKuFRkcO5CdGv0RUpxWWXXa3Ow1704O9lFE
ejBrYdAitMoa0/Czk23vAPBuZ5oyHp1fjBbAb+GS4k+Ii8Z+0LUcYhuV1Ib+UmMR
8Dp/bfV3mrRseUdJJ3xtEb0A+sIIgxgGheWJggsAINt+UrcJBKgJRMcr1h53X0d1
pbmAI90wpoKC3dW5/tpv/+uNY4Y9aIu71LiJ5sH/mQv0pgqugm13vJxSpvkwROii
7B6gZn3Etl8h8e3YXTNIRhSEsn9n9J09082LHDdMWSimtxac4ievOi1MFQ+D38eV
nFOujUV9qZG/5UnWPxrkRGfAwWh5uMAYXA4I6NHAUn+6NdWPwsHF3ljL8+YwbxBG
yykgGM2ZT6pkm+BPM4vsO0WjUXj0LBhhDlTwbDxMP9XePG3tx8yJ5GmaVDfwZmNu
D85gaeAvq1E/j0yobi0DURk0ZuA0Facusn1YYWXe9GWk/mv6vLw+88mj6TZYo8Wk
UNRMLy/Yn+5+HJx5yZGqDsx+Paaah4knhLR13zQTdMqhCiuBIeZ3Ahi3S9Ez53RI
SaRbLzHIqCGWJEzKzywgEic0JlF7DUjimsVJbna5WHcgYoJdID6OjpEH3jQoAkk4
63MceHJetigNHraiKZ24Cq76lsZCqhKmpg4yOG5nKq3H6sT7h0IrmX1T/hHXHfE0
Prx9nbMpDSI7rSuHk5BxIfEv466dRddhajlSYzGz3UiNzJKr17VuJdRTTcMy09Lo
W3AZCnM85KUPha0xBfq+oBuJbKHt1DX/OM9COglH28pAcQvlJggFy1zqChtAPCXz
QxjbiY1gOBA+/xeuw6DUqmjCN362JE1wklTzQgoQF1QdUN3R25JqaVG4uvOeb8Tu
H3byUlbtmtI4dQsbi3iN7/K9U6a2UNlrRzZ1IzrspNxHmgQKiVyysT6W6tSguO0d
ydwL8+7+3kfe3lb8R+4SUtaWsmTrd/7e9BQbJr7HtZAH4alBVZHZNC2hSfTNUhzl
/lVE8lmdyMa2EzuBlC9QN6aMDDCur3hwFOvI5GNBgU8VlT4Y+nUaLBnu9MDo98BW
hTtMhDe1zmsCXnabYdS6mJuMGUeLj3qChkwPcLGVurqlLHlD5k6nUu141ct49d73
+MpHJoqxQDkBfkFQo0SNc4dDVDFkVfXlZoAdjlAq/mTb6Fmo8w0bahrqLHxlzNT1
/0kPq7rkZj6avmQ3u7GXVkutC1c5c/lox/q+JkIfQWvlkIWmUyj093ojQsdS22XL
Q3nYnD941+nm9GBRvk7mhqBS5gJ9I18teJF5lukkfeVkDQxk/ijXASlKddOIjk8V
UZ66hX7Gx1cqmQvINsECYPg613rS7FTl2e9ygWh/lebr3BAfw8STeSNjzRrKyV74
r/HG9vqJsvAiObIgZyvQ+27GqYR3cbRN/poNcEp3TFkQk1RgkIz5/bLWE5zslUFy
L6pdrm0njjrCpeCRwg1hGw6zZh9PmuLXPBT8j6p8ZQNdMvEI4tf21uTCC2Hpm46Z
+gtWYzodw1gaSw36vFDbf/mJYEPa9sBsTTFT2YIMeMnZNZMGA6trP45q+xKZ1w+Q
p4uAkAJzIJOO4GEGV33JuS1LcwZloi7TjzcAhu9ELYUDHxN18bVyzVtS4EBon84K
mbECii8qV+DD7dXBg4qYxrN6D79WxWfCYYFkEqv5IxNlkjHqA2WeQIzeoFanEAYr
4RNCSBl837UZPBwvprv0tNMCv52dlfI+Ho2Q7xeQPYWd5M3VUzznd47tYmXk9XGE
5SDB3fSUi6ck2QoPN6NwPX4IpsPZ9IMSIpM2TxOjdtg5S4B/NYU2SioJ9U0EbnPg
qHZbE8Pel4aTHd5/1YQA78YvLM4Os2ecdqKgfDSe+4eEX5vZ56SGryvRoGTQBGYq
mvfgCtrR28ed6DKDC4yFQKS7xpr1z6+FYkmkOuVx/RNC+TrHGFRHbVyECAlaw40K
86r0J1MTYRVR/IDyJFph77euX1y+1w5PVXwRhybfGra9OSYVI+NXS2UKNmf+eFRX
sgvi6Ut+g1YbfgcsSygl70ANHBrxielxbbYXEoST6f1k2oWvNUPHLwTKID0Ibw/N
HApMlQiWO9eFlFKFC5Wj9Vly3NZYYMqaEfI+SxCvGtIfEQnXYOhGRsgetv3dFnKb
osAtIwAdsPEqbQiMZTiobrhdDvyh5cEOAU/vsBwpCSEKi8VKG0izuTlOiBe25dr1
TZG3Wrbaf9K2lXsyzebBhqswtDDuOy9flNAeykBSgF+atKho5v7CItXuxGtDH7pF
4kbl+E7SS3DCmG/qd7ac7jpLg8s6i0trMUOlQscRzNz/b33iYqUKtdsUlfcoi9s1
OjUOdlKd5fVm+ntkVo4HXoPyw4LCUSAM944Vys+6ftVjTFPjiMZH0IwynJYkBMvZ
YAYjKb/pS+IPAza129+YZ4w9gxijMXgrsh6KZi9SbKk0n7nBG0l9QjrpXEGZ4Y59
K2hBXDvkxU13M4N2CnkKeTjoowycGSHGjPjPbTadvGCMijeOVPIR1gOawcwR/p9O
dq6DVVEYdPhFl0qW6/MgNQ2S2ryP3WK2UFfdX9ItPPi49K0MsB3f6SGC8/w+1cUg
Wul8ZM6Q4GVYkUMl9lijjcj7tJByVk3mSvf/JwffLSk6Eic4UzAlsZU/G9OLsG7Y
fKMkbFmvPSryLlEywGFpGtQvcxBmZcChpUnfgbElAf+YvKrECAC2rwM0/kopZmqY
QfBE0zSqo3tMyOSp53m6hqDszz8yCVRBYmwqbD9DbRO+WgnjoARQzZJU60yfUdJO
1RDPLDrup2Uy8Qaf8JiFFHkTZaYq9m0n4qiPNfSU3m+cKiBhdaG41J1dpbFL5Tco
eqZ/mwDvcLwD5a96/bRZS1K0/x9moIwIWPfYNt/2bgGog/DNpSsVSktTDxUwE5Uj
XlXvRg0a995lcCOx5HCo+VOmz4JRliT3QfuLheZ0GRyFzypdW6Wlfn3f77VHui1Y
L1gVfe7usgoZA42vr2/REi4WHfX0ue1KdWVcp1awgTOvRm4lZw86YXh8ssdMXggc
ycq9jm4cT5sAJ8dMLyyMsIDZc8iwRU+mT2RZJEgzE4uL/rVeg9gs5hDAD127WLWu
blOTW3lRSUnQWTjYoyKo3El7gszYopQ10usIKlNrwZmvrUNDtsZ8dNUfZvFVJEWP
FntzhmfR8hckEQ0WWBpwQRPzzon/hqxvJQTLD5Ez7waMtdxD2pk7PZC44/bqwV5S
oXLWyy0zmWbmbu4rpoP9Qdhf76jDe6EXwIGQRq6aHc5cY8+x+MkTG+5o/19TxgEV
DBYoaVoas7dtkBNUwcJ+BrQtZJRrI63IuTcghtHBt9i2NaPay7jNOMj28/Z9s6nS
Rq0faI4oaiOhq7wHmuPD/C4mJmUsQodo4GGuhuMlNdwdXhA2bJKiV+Za2E/lZ8jM
g76/83PsmbQTHL18eHWa9wS2ic99ShqxTT8tx9CVMm638OqmL4vAPNaECM4Y8ljx
Gmjvqs/ZXsGQ0xE7YtWqYlHnBN4UekcZdIG6OsWNYrymQlOcPVdIW2Eb13iSX7AM
G3ZhvN+wjIvMU549fsY02arOLwRDW9BqRCjtVUXErrtzZfRkdtXZheX5Lm/+lDMm
NECymjkKbhzwur93QBg+YL6ladvPEiZuOTWLNUWTdg6WjRt5yxLdik+tCNQYGtiK
U2RuQ2CZPTDetWNUoR6dVOE4qkskti6YoChiX3xJQ7eeKXXsH56/WB/isH8+MtwW
OGRmTt22elaaXGi1Pg3ilzLArQ6QC5RoUMKvEPvZQNY6JgsOndWTZzZsjdSiBfUm
9g67WJCr/zCS5f1Kun7lm/lMz0isJeNl6eB5A7wNMHDFmoqUdX/MTH9Ljk262KSK
rhLthcL/ZQfuGpxdN0mSPzK17TF87wExd8ehl7PbCT1p1/f3VuAY60j4AurcIqZ0
DryV2iceAoHDzyG5HHDTC+COgcNT1jLTSjNQ4CQ2TRFbVqrJVZkgrX3lv4Hvv48q
f6nkXztDUhaBiTq1MxMr7XNja9Sq6JMypYwfh2THKfxhaHRcO4xm6xbC04UeaEg9
9bkA3IbJ4FxXwElGMtGuSn+StetQKGWT0V4EsaqQhTFRGe0tvKV81D5IZA841ykU
dG6InArFwIieiLrkXcL3Bnx/xL8ClF98A0VmrCu5rLru2EU7TGWTsd9y64Uzb0g0
2sA2aRT8n8aXIKJqEKUk4vN7Wwl7RWHO9b2GO4KXcBe2U0cwt1mak2Y+nV+0fO6S
dbqWmAnHAp00N6f8rgCSCqanUTmYGTrPhoqM4l1NqxSQMzuXxdciEWtNaXaM4gfm
tdj/mhIc8jnsmi6+gqX3QmPgjWXWAiGS3FMS8d0tK5fLa3Yh4ng/hI2987DfmQQh
UaTmTjPr6XCNAhPRfEtFORbZfrfch3bV1RRGjxiPUNuDwL8M8mdG3d8qdqFQsyTA
IDef1VBgywRsXwUi/vFuumaLZAjuPBO9hOtST24t1Ff8HLLwv7wymeosXYLaOl7c
urt/jQsPY4j6ZDWqYhr3GggE1gz87BsaS290lkD0tqAOkZKJud5TVsk537Zwasrn
V1hGBJCvSdJTOZqTOG6WxMkGp4zfZiwLitmjL/ZOmiL1vayrAM/oAL8mY/OEycu4
JISqwSSAFDfnK342Xxq8YHRgYplJ9rsHxs5BEnBwgAq0L2wDfCig1hTlAiS/s3MZ
MqjbiS0Vlahxw5q1Rca7Q+7A+l4Du0yCG4ee5ZY3HFeTZUie5yRE58+QaHqlbW6o
m++Na44xt3+tprcAP2XgpL6ZyyLI+LApsTFwxi2GxB/4fWoFg5FXG1n1oswbsc6C
pKlWSGhPNiwENxdZ+k6rT+4zce9ofT2G4v9/Tnbqx+U89DLzsRdKOdcSyJhb37Rq
WIx9r3RfsSTyVaNqHUKC3YGY757Vj5Ub475tbIMzmPYbDMOmXW6nbevzOLHzoU84
TQzhcaWf4XqdagJkiVO83OwCo7/N4jO33PAVqoaQ7sWbN603s35YXmYkKZSKdL4b
jgVbJl7oMpYQGheh0ZjRZvK2og8fQvv+rgyUJM/AJov/KpZIU4n94acbBSHw0lm3
jARj5uWOFHldNDln1bHmfwMUMdBZknusgEzt1s+/arAqoJC2YYwRBziRoNpyBTKs
gLGAfbW+n5E7OZ7QAGkAF3um24wyzEad+LBqbAGSJzx0A/n5RV7Verrp+Q2bqYT0
nOLkMJaqHIagKfuVwCAKQ7YOaaJH3r5OTItE2dhYbe1sM8auCZcszpieefOeaBYE
UgcR1jGjXz5iDSyONVBEqnvI2uTqEwlpeMQi0PqCLWCi2wChofjp/9YL5bJT6RYI
H/h1wQlWuwengNjBMEspFUFt2SR0lgBrqRwtd14LKVUoBKCwM67nlD0nWaI4OoRp
+DI++srcb/7YhD6wVlwOntz+t23EoQ4S/dcUB+33HcgP665e+HSnd0MPdHjQH2Ji
+poVQTAkVxGjQzEvOv17hgOqzz2YdFM1vWQXvt/75R52U60XBjIkDJIKP2tmxf7I
CeVq5Dacyk9utces9Xcffl8BgiYNxgm/EoT0K9ZxazPBGwg6H214/yZztWyXQqWv
0ymu+zX48bwkO0ONhaEzfsskPkMkqJGTnfM3vQI0TQKcvue0Gsy4D9XclaCCN4kR
NzVbsuMvoI8VO17/qZ7D7dFB5+4ydHTHeMp1L4YSS8pqBTzLBkz5mJ83xShvv7SW
Iq/8UCiMyGsgsD+HOcAEK82Zfr1Gr0RwwZWvC5lZc5PCMdoMP8wO7Ou7qc7eo1A6
Obp7UlvVKnmrFxNvmyLgyyCtEUtRueawdbxTKsKm812X1v9G0aqH1GOX1v8fJshp
9+178gSi+rlMcwC4SYQ5FKAHuXG4ctOatvj910LQtkOBehbX4qqLIH19LqAYEzH8
ocYzWWzGsHTYRdR8lDrns5bX1D9BEwJM/h347jH0+CDzzQPpoub5gQ2vbiqmMjU4
1JBBvaFptc0xDD8HykhvbTvv3xo10Yw3S4/AgnDBcHQeQ0vtIPVw7IqcDnRcylP0
fWxFDl/tnQI2uUxHvFkZTGFuy5pgl8V9L9fqOBrTvIwmVvct2CGEbLMcRPTZAVwR
oBOk+LOe2UHxG0RVuJO6IuaPsI1KuP/CtOrCU+4npzoVAutgxfJm8CZDCYF02u3t
SDEMewaUr8bgRuCg+DqgMxNNMHok2sRsXhsAzp6pNMUXx0uF8j3PaNSYpJYLQ+iQ
7eSthyGEd8QifEHy6QKBxOhJMl5OtKjBl86K6K+vjMrtzDiEdC8m+ZVhsFBtegeP
MehwkbjXGqAL1jTQmI4nqT1df63Obv6RSv4+5iQq6jfLXA0V15UpYL/5wjrPRRoh
HbshqCSPoTDZhxwH9VdnJVF5fKrArokdBUIo57eJeGKtIW3XmpeYfcmdD73LUxMp
exDg/QfIzDHGf/hXoovWq3k6+oNmh4Q6VRzzIdqm8p41GdSWD7R8CTLsSIUP5Kr+
ozv1+Aey1Z7vhKoBwwOvHahAddi6N/qUc2TuZW5LB/nzEYNWbP9rv8HHWZ17DJm7
2xnqOj1v+hySFrJqlAxPkwwSLR7Q1S6TyTBxM/Q2qhhcSG1oOpjl/TiF2l7Dg6jQ
fkuOroyPVRN1lDiuJXDxjcf1A8E/Cl92rZBChh9gJz/NgU1zr0JD7Xr6MmTi774p
oJf2dOhC9Z0Wc5g3B1UMLlosSyZWwN4deX6ITvQapVNFTs0GCDliClUuoAbA628Y
1sX8YiEidKNMPyP7UU/h0+ICzWQt2a1j5E2MCADB2h6q32rjftRjMmYJYTs8qbuo
VCV5Xvl8TN+1wOHU7EqL9Q92HjMARrMufYTfNcYtcZcmMvwaw1VUEX+FLKBnWTQ2
ajGDsruzDagY/rK5ZkefvbsfiER4Se7aaLT/l1i9JbxluUx0GFoORV+bDhSZsA5r
eSQKzQnlP3+Z0hML/gCbi2JHNQQ7mNSawMNzQbnaF0Xr0Nqbn6D4lYLvptTlDe4p
qfDb+2HLSY8xJ6QufmHFuLyDaRR0gQT44IjAEeIbt7oMB7Q4mzIbxKRAOQSOh7KU
+AyCpubth/Knp6aA2oAelKi7Y9B2U1kc7HmN3NOTdt0jdjnajPWNEB56DbW/CtQY
A9YoDctrceySz5jPi3TxSey+6cVJ3YcO0L6ANPKcYc08ZmqHe1R18Dy8kMmo3HoO
H4e02vuBk4BvL6pyDjWXtZnnc0041YJYw6Oi/3ObeHITnxnCG/LTZB7t/Fn6m7qB
wCZ4Vl+r2A4TjIx2RC5RMY28UA7A5wXyOg4x9gWBHDoMCXLY3EdvduIj+YvSL5qe
NuY3iXiP3FwD15GZzHZWOI3wqfDQCXCnNpFJBSK50G1wZfdgIweMr+wR94u7DLsY
GyayEqcU+vFNHyY9V4BFiqr6XJ6cqxDXL4lXapZyteyb6phHeiW3526Jjt5uqMXr
o48gPf9UpCzJz0p/hT5s7t/41U4vpQRxhxOfmw4FTpaPe+xVU5o5ytb+k1bBU0pE
a0VDDpvp+yCVZtoWczpu9/UnwHjhyknCCyuN9M04VzI9/ky8HjnadNFndmDCiR3u
T+JHMIJxHS3JxUpsnlo5C3QCEJEh3lTD7/0rDwmJC7RT1JgnW8zbsGJbj2/WcqbD
CHwjvQkOerDku+TbFukoAZgBxtGVzKAQt8/f9ONpXjkf7svG60rtLBugXD0I4PGx
kNcKr3OB67OLyDoy4VIom4QJrrZXs1zKjBALqeAaX69f9DvDV03qhzHsrJ5mVyH7
XPxGsz3JF0zImKMnnJU7YSwtvCDbtdfAUx/C34/I5F0akKQNtTTAxm1iGwyg8dzd
Qxv7EHK+FL/Nk+JMcL+AWE2udwZubpgY/n4F7o1eF3a1a60Hzs1vv+za4tbIEL/d
SHiDXkjHxQuRMVw9D+EAecfURk+O8/uGXAC5s/nTF6fI3DdV768c2U5rzbYW/jFq
HmslYwFgit63kFTyY3z3GuKqxuS41Bc7wfs+jNHy8Jva9xOUZcUcOIz34je1Sq0H
eKKMddXvKbdAOxE058m/N9BTAdyey8+nJrX2741PzmrYf1FZpQ1Y+nARRnaaDxzM
LwtI0f3R3oanwrITVr7bE2xOpFRzaKaK6CfQizGM3J/jxdlz8BMW3BZ1HyetteAV
HnxXPKEGLyJvI2f9AZkSKPKUNNLm4S53CG+hLWRwQe/ae5amvdpiV2q4KlbeBhbq
p0xgQXHTK3SwV7NVTRDjYVX12YFvNb+xidHOoAaF0HMJeZIFi80WJxDMbHrxQq0c
vLRMPZhg6WFqjmHRzrD7AcqBUR54Y9pDEAhhyC8j4XZUaY08eM9ec8n0byn1oTWn
hA0ox8LjbUUNubw40xDIjO7q6epBzeckxuuoFnydrJegOwQGUZ9QD39ddYGJF1TY
hza0yW/I7yT/DTY9M/Nwd0JERPdle4gBeuVZJyk9MeHA06uTnsokdmfZ4XdHHBdR
6/2JV1tDjcxqYlITHGvTCcjJ5xpPtDg3dtIcFj8FyT8AFx/oC4i2m/q1EQbsfPfG
XT1z3Zgdtj33t1JMnina5xx0M7uV/+1WGCWqDLbojHn6sTqxUxOLZUhsR1OHPPqT
HI1a7UurOwtBfin9P+NwfIhmxC0e/ZJ+T5ousJxvw3TWtF0/aNwYAuDtj5/rJzBd
p9EnuZOQmIHe8qCMncJwsF+4xQpYWNAK8LZMTmDt4AcSeSpxBK7oGNyHnF92WQsV
zhjqpb+OloDyBJY6rgDJWrSJ0o/37Rf2FxkjgDNLiJ7rmttxKMEpzrYBRPb8z1UC
dcNqwlmX3pif+7rv0Po77MzvibNq7QPUNHBGVpuqxdEMID3ut90N4C5UkVY8kg7i
ZuE2E442L5Xvt8Sxlx6IKV9ZEL4B+A5y32vF9EZ9L45Audgz2JvVP+98/492vGWK
VVQscuecvXtx3mdEc594HzqYwvq8pXSsp7GcLp6T6f/DDGBM5vUqZ89h7AnfN82O
iaosHN+VoJwn9zr6+CFkTCw0Wbac+RjkUcVxN+MfK87PM9vbkeWtzirsS7q5LoPb
+yBvlcAkfssjZdWBu/RsQBrdNDk737TQIMbtye1T3TW/Y5BO+iYhJ9kMTmMlEutD
gVsZWnHLI1vRFrDJ6dk/gO161hraiX7PmItYcTtQOpse0Uy6dX5eUC3aIDq0QkMM
H5vj7SFjfpwe7PNdt274kiLlXeJkKr2bGNGZcQSy7tCIPcyGSpuT5Ka0pzXccJJR
dyUclLmxHLnvFKYAzeGHfBfG1kqqcvAT7jrMWg+ksH6SwgH4J8JVsIDrDEEXsHZB
zlVFhPDRD4exHLpsgcn3u6mkTUCePML3RPDeRIB+JX7gFJv4OoOKVwE/ivEjML2A
l7HJ46/WaGigH0Lpy16rtULNehgMRDZDPsh6QQREt9e60ZqoIjO8bluHgDI16Ji0
b6QHBE39stlzZSwgmDs61ny2rlSmOCn6m9Uz8rkwyHL3r251TuPNZB3JUhpu2mAV
jQWfO7ENae7JJ23a3+0SW5G8AwXEfjllUUHXbRnmCgWZ1Q7AcHPgdAJWnsRcPK7m
oaTVG+97haTS4hudjY/p2UNt5Nd23U4SevTqOiXoAYZT0XZhBHvgBz9t+sVHObUX
Afw/A+/Fp0UJ1llowSvbPVQ8JZvN9LryZbAJKcPzc7FVEnsfkTUVPtg9pt8WHDuC
X+j058ydD58M/xUHh/BMNV4hPGjOE82GY1J2czRHNHNapTUk6Q5iGgLTDE4XEh/D
T24uPU9m4rsahmD0vIpu98D42k476l20+zR/IMREMeFkJP41as/biH4/GwOyBBV9
kNHdeUJPN44avGRJT5i5Bl/dPot3zUd8cEI341xSOKzo95LYECMp21Yq2XG8xv1w
lOFdbtuTU1sQ4Zilhdx7jJNN0vMcuQo1nsNNpYcCfQigC355s9s+8Vt+sNE2i831
BJeKQmzWbLTnYEqTMU6doRJHuWpWP5gQEas6SzdWqoeOxtYAk2bp3fQl/xImOcga
abkcMaxoIhT+tGm4WZqOkohYS7hXKDz9vJ9orcGcgJ07mwEJ/rC9uL1Tiy00mQVb
5cJDs7QzfmwIvYGuMp1gEZ6mQd9ywmCXd7onr67mSzzh0Y4+P5ShwgLvuNKREoJ4
Drronhugd91dlC9fAVrFDMPtJaXx0Kbh/2JAe2e2DbffCe7E+K24Ro5h7jLThlkj
Eim78fDcec7Dsf3txtu/oaw/Ng+7qySSGskdlvoljbTXYTVywZOeSf+vam3dFDgi
9SNxDjuls8BpvwwySoBHH3rnxphY2oiVhv8/i/QiXyO0s7T5u9T78NoOeciit9Ul
IHIP6vjyPOYZt9SN6DHPR22Tai0VZ85ewY893SWJkoAauirnwwiNy7iq4T+uvCep
dAQiXwoRWhYWoZFYrDgaWyh0/6hZgVT0bRKcGLZQns4BESvKKeEqmAifBJxCBLMP
ey7DFIDkoeU65GrY5AUXnU7AgQNyFeglOGVOx29xw0bWC79kxOXkIrBa0cp4d8HP
6jJYpSQ0IYhCZ4D+6nK6SmOSKbu1qJBIaEfhJLknWQkfjo77V3PQwUivoBeDkGxO
ua7dEzEftVfX7nD/4cwQSXEhUMa3AXw10J72ljPP8BL4PcTCwvx4pY7WvBhtiNDA
7Kn0JvAhlhHxSqV55OnLduAUfVCDXcj1YVRe5EaKTQcDd/KuWxeSckF7r2DBn70V
EjcKcaBqb2dpQKOaCXA7GwHsLtr22jfxun4EIS+gx4jyoDTUR2Haapao4jZV6lTG
Uga1ruMTet6CYnvERGg+LJCn6eo+DkZ31G9N4ylW0JB4hyyf/A99F/sqKFK+0tIu
0w2d0mEKAK6oNZgONiCBanSCmx0uzq4pnk3soW8jV78pe1XKIi8jPH8eR8ovn4xG
ajhVqJ377tKXTpnq9uQyK3A/v4lzbwWfQs7xZ9cPE/RvBt8A3wCbNW1zOejMg4Bg
mZWnOe8fw4DZEKe+9bWdJ3wHd3fP9thFe+IfgJETNBH43xZGGMe9lyk4HY6E+rz2
5pXtSdNfq+74yjTbk7eje49DOh8B2A0znlaRBZ7epgN1ALh2lHIO9BQ9rhAjzZ/x
PYxYxAi0xCrzbJCKLnF5HQ0OkG6nVy5aDMPTKVUIT8Az3/5xUaC1OyruR6MeZyIg
18EVq/mu9KMAH4GifSFkq3lND5M9LC75mn5u1zECOv4uoFc9iGVgfERAFam1mrDU
ztHaDPpVAhAnPiSd42QWAhaZ7q3S4/2HSl/MuyHdJDMdLq0BxJEyT21k2E9fw8ud
yQeOGr01dxgOE2NSX4S+7lnhO5dgPRy7EbQQZhATeEYM1Qp2bM+V3fHyLn1xN6Aq
4v9YEwvoP3PCx+2khitn3O52HmF7chzOK3RUfYTZfJ0NJSNU/gab3U+cAIuMBmbH
xsHNQjZwkv7DQes+slp6sV/lIUz70b9GuT7f3PxlSTgwWve54gs5QPqUNMIwdXP+
XY3xhpLzwFDkxgYbab5JnE8Dy9KI09qvAOEDRTQsfc2KT6N/cjifuItP1vJzK0f+
pIqVMBGM+3IbMT6zQQdfxFQVgGchgE0txu0EC/12pK4kOcfzPraZKFzFybA+kZlR
GTE3C2zpP6Bik2/frCoqmMutFAomAJCm8lrpCK/tBBbhuWh/adm4m9GZSOqIvMmZ
hMB3sCGmOkbWc5cWAowqnR1rFQxilvOrYzLQK4A1rN98/GDgxMEvVxtwjNS408nn
/vc+F03AzOFRYXh9ZjwXaK9Fh/uBQFall4bzQf/a4O1AfZwF4VlS5ShJSKKE8xz1
PKIr2dAGgpeNLx/Jo0K6OJw5TK4d+0kEKL7uaQR1O4HEKXkhjO0yBjAcbhFjnsOn
XCnChPLEN1x3x1wHeYvYrtrCiUQsubWpwpvBSj8+5foxjl0+xMKcSzUi3UPyaKHI
TI3G5cQ6BS7RU2YFMZ01rbGjBNNNez9JQeUYO2PZDGE9ufMg7AeTmQ18H8JaFvVP
oW1cgcn2FShHgnl9kq9KA8MbWhvct1cPUIXx1ov+P4mDsh5lpaBzNmsAYuu+Lh4+
k6C4yp9P4IzQ5o3y6ZYgyJEmOH/4VenUII2eAZSdt8qopxsUZ1Hr83JtzpMGN20f
KRyaoz+hoMJRxJ64WGrOmc7QE4yHhmoyLUyMfqXeiqmfFdhF3E3fS0e8dh3qW7G5
DZMDZ1meXOUmK8z4JuDBcnEu6WYG5ER29EtgkFoKshWGlB2lCx0w5jVH1+0FhOkY
M94rJe2QORNCgUZVhOqALdqUX43gwammsPnWYEfIJVgsX+aVNRny62JuLTusFpGL
2EWzf6AfB8asSCf6J/i6EusVXw4FDqCp7RPsNrUcag9OG+53DyDRlyTuJQ+a+iUt
wVGQDvqr1r6amUjdFgSRtzq5aNUTqHCq+R0JyVM7S2CvhEvQXkn00uW+vn9A9HvH
dHKxRiza1Xh7MJY7IyDB5PbMhy5MVgTBCRgay4u+bDiuZDyd9v5rbwof+lE60JKj
/izftdvbzNw+oVl4MW416lgzDBvkcU2lc1yuUlz2TuEzF8FrfOhJ+xR/YltJ7gVB
uxFGUvIuTAXVDfm0l7pYt17b/eflK9v1klIzAKE/Me7AsqWT5ZzJaglWModt+TtI
hPTQlr7R11jmpMt+yhWrEBKhEgqNW9r6OHAznle/n/ge9f9scxqyqEz55BTjxlCl
GyuWBf/wCT+eRfzfon+qPnO56hawcC6FveioRT52FnRIOJEcO8fFonsWEPYGGzNp
RjFff4hyEtFkoJ7mlGDltAN9WkbZXUen4CUeeIYxcy0ZSM2MxKehmoGCCGF7uEzC
eiRoq1Zs+rEg/9VZrv1CsR6NEncwVkoO/04NUR3P3iO749mVlqdAsV+ZNmKzUxm8
/DadPcHSUAqjCx0Swq0dLiYHC06wWhhebWiNJIDYvVxAdz0fQ9iFEcP7EvVVqEjM
fG98wKcHzrlWRWOEOsdWkHrg4sVzrMh9v3TcRVL31h95MYivgLLWsSMCo2iMvEfZ
HwtIKUfCFaDE4BEcmItdUcewf5mBAAjfDDdx60jRs2fqz3fEOYcpGZ5R5wwX0zaB
exVVUCHUa58y5XfdEFMl3t998e5GIMv0GpCxY95VntMB76oFljgQQhIim0nDSzNi
ANxbjSWUojChFq/Ny61wCyMx7JBf4i7mmaBf+n+mgsnL2E3X4JoCQzbOOHnCksxW
sDaQDhsYCnjZ1J8306MFuXVaVX+OhldTgEGPoTRnFpDmlcmQu6jUitNM2FvdBJhn
pWvoOyx+wLdJ8eCG5l/TNaDARN5pYXiEcBwpezqK+ZoTyP4Yuas9/HLcbZOgQQrw
TJN5r4T1UDAhGqpi7noDoirRQU6vGvjUjTYDx53h2r0676iSxSaRvwAY/G3mrt9z
YTXYxQn3wHwlntoX7kbZcJgdEpFuCOe8qNqgv+UU4O/qYV8zd65J6YAH+gDZFsbB
n9OQ4ROqrp39e6spOKFFnM7bOAdqXbJkDUHNexK6S7QfqVrEsfOKiQL7WPUzfDak
65d/FaBBHT4RBIzYE8VhVETz0rWjmDneqcEOuHFT81n5jET3sBDqyNi36v7GMsTi
LHsyhNvl4gtecfyeVtuCWBxEgF3ReB2jThMER0QXurbf6OZxOR/mo4n9IDhtjCeY
HswVJITr+t10ELgHS2fHtOO+4GJjxH+O9Lg7PA4WSWhYShverY1yllqEgjD6FpkQ
0rk/TxInPyrFO0V1hAOBE+wgims0uEX2UrPWzK6ygQ7bVsZ5Ve+8loMNI1X5G7cx
KuqJKmrTvLum6h1kOSWlNhKmnpQOMjsGU0SgXZzMu/5Tst6bhoMLr68+M7C89Zcu
MvVo8/30O/6ke4XXtxSyYJHCp2zfDWsZQJq3f11Z9EG4TiSxmt/4cC2hCWDXOg88
zphTAKrS4VyGbf8ncm8dBpn/UWMDDX6AxhnOVA3T0+HzM9iW5wmxpoIFT/TfTUqN
Z2zGorReJDK+vBkgoYdJVBJONfT2zimOux652sNvUtNqdj6hx328l0x8T66iD0ci
uk5uz6irVfZ5uCNSDRk1rbyBOWGym0osgjadcgy3hTMB21oOdjLJMQAGNqE7WIYy
txJo6lvOSd0DQ3wGZsj9iRTr5HUaNPdwGlOLUY9/3mM74UXEACPIeCnhBsS1AezK
p7TSVcUlRqiQiH1I127iC3S0e+A4VrT/PkpsVaLx/VLHsFpOB1Ef9Zx3d3rjfnM6
gmLNy4qwYFQGazTtg2oY0D+wSFjWZpDi922O5W9l/vdkApwlLKCaS1ayjaHviz9Y
av1v7FhskkEgG+a0f51Cxg09MRu0X6I2TC2K5tnStzaDtO0hy+CIlNKsV+69JJoK
q3E+zOgmm4qmqRfVxhVlvkzad7gm9c05LAb52b6Pv+PClc+soBxVOe//PbGNdt7z
Zdme5SreeoaG1JpP3gJcpJol3jViHtf1LcFotefcUfKje7qZ5yPRUAtz6yKC2kTm
I2wIjSNqWcfXOMa8UtRe74HaYz6xQTPBxU0JvE/XUTL4RcKykvKARDSUJ6YVvKpF
UJAjHNnzHcqdJolyeNhqJtodfagsd1qyTCjueZsLMwzbeWynWzPYVFO80LqeeWf+
JoCVatNqfaaNR2y8ai3RAhAqMe2ws7XQjIxsXYW+rLI9JSgVZJVjNJrgG8fW/MXO
pzVhiG1n8s4ubmwBZTcA13FSGu+Fl+GYth8Bv/ShevFoYW/15GrDj8QbyRMcyeAI
wlVC2TR5fIUSTbMiPhPDr4YLri8ZLYAsM5e6Z0P8xSNBEKpSizQrkaf55Co3YX4K
f58eYevJnd0tTLQrLX0wrUZ5GfeQYlqZGjkGA+A/ooNFVXMBG1YQS7lce7fzxRTU
VNyjTGkCdo4LyQbEK+EdAy3rXrfIyBQ1WT/1LlnIc9d3zik59XL74xRRzsHaqbr0
xBxicB4Oiz40sosOJNizIY4tUxxariHWxRzyUSYj5jmqVs6madsI/H+TcYX8l8AP
67KXWfu5Mx98lg5nvUWPeMCrvqJUgg5bltXmjK3RyyztAIbn4eyU1Fm+9j/sMUa4
SNbWXGqgCSHT49k3rg+1edQTBgJXMvfEjd4g9xaKfuq/J6T9nw36JiFVneQ1ivdR
Ssa6XAABbMnQbOLVlVmpKi5yU19br6XOAaUXbzID8h6+B6OQx4qioJMy69GvZXWL
xidY0Ce6McwwMQO2LeCkzO2BZdqSJQcqyyOJTBvSPUcr/RpTCYMERT+t4U9Ri2hx
jg1Ny/C6YOXBQSeMILVi84OjY9XsmZ+pTq/q34gJqU06h8ByUufj8zb6IAdZEWHL
A/879HaQ/VWvFRdVy6S4kQ0mFSRvboWDW3xIR6/3/qcHnQQLpMHxwIWTMHXaP/4K
OmGUCqY9QmkWFCkb0mvpjsFYn6Q46OV3L7vw8j9gB3C3eHVZkp9vLe61ug8G8aKr
+7ShT/y38009hA7+2mWZBkZmg2eTx5Z3PzbBue3bZErdQlcbEIfsv5tsNhIC5Iy1
GP9Qj5xsLHLJ6F7LTd6U9IDg2Etg3h2U4P432nN90rKxVdfgA14V7VkTvD4HIQBE
XbChuvLa7CAvYlpdiCn1aAGksMo2NuaK/RqqbaMKF4B4fI3xAPUn0imLxobJHr1d
A7zT9p4ZJSp1g36GgCD7pJ4W2szU3QcgLEEh1KqvbwPtQuCS42fkwiSSx9MCUl/H
eS28rI7svKERI0eOqFaZl+7t/QQKkK9cId5nSLzQs1lJMFk2L45GaZ7OR4UcOGE/
xWHcG4jm7RCf17TLLjVXt+FQr4k/dxN2sPJL2uCEKmrFf5f8QvLviOe1dgxCgsB3
DkTM1pJe9qycbv4SoyP3laTlFwM1qWyzTdY/qjmFHtEBpcJ6idnPaADSd/BJJ0LB
yeDm8TS/9HpHhK3+kIu384TJ5hleW/GCK3Bk4sE8R+tGYWkAi5SWkyqaQYTz5jme
qQ19WKdF4mQR+DpORrLTcH2cGb1JZKbaEhoanN8auflr/lSGuEmIAyjT4mBNUbYo
ad7qB70ZO53ru99GU/MgxxRn1i6doRaz02pBNN/9HgUYHZz+M4hXCFt9PxggS68L
4MPxdeoHBvz3Ovz8ByV41wnRa5yee3Ut8sok7JuBXJYTkbEwAyt6YmQgVCzyi+x9
H7Ki/AfhUnkyDwrQWVPWpWsjg2wKdIjEeKC2HvdPfFIzeQlGA6M987tTaMN7PzRA
cGXKKTH02sj384iHQYRhR63IJVYkiPcpLq0B2rrqoFtxvrR9M961yao8pxnNYLwA
EMo+Bz0KLahwEO+taJR/tdWkIG0moJyn5aV/itqR6MrYBzn9STgDLwvo6CIWHGwz
8BblIb7CvuxOc03ie8LVVI1yYny1opaZLA+1NTkrkmqsLyWXVdb2EVw6ZqvBBZrC
fVzMX/SrZE2Gb++w6Fj1PGS/ZoKyb96UmTIOZLQNLdRJImw5+gd3Vga45P6tmyD7
5EFxQWEIlkmGUrb8EQP/XvGqIx6Qask18kPylXrQrtcANiZizjfVdjpTgJqHR2o+
iRoF6v+aR1Oo3oAx815giRhkX+jyp5fw4KNcZDgr/lPKJWQ6YTm0oOfOP1sYHGwD
2RvYZpK5pRmLoTYrQbT/MiF/MYNh0UJS/n6+M7UEMXBSJFNw2eNohEnwen7pmNBM
Qd0p2v5wxAelJB6KtMFIBGVCO3eyfGqniGS1lkPUp6Bt/rrEUdj1qBJtkn7jgDmM
ulSGmCI4kEzfPp+yjavf9rEnKIHRlg3DxsjapIQkkTmYu69PeoOL0bjdvYD9448u
LGM9DiDPgsKLWUxPP6o+ddEnFdy86W958H27myL8F49Fp0mMwA0cbFaVdYrPG7r5
3PuUXgP9FJgTTAy04gcULapy2YtZGYYL9GTXMj5329FdWmcDGRz9ibe6S+psDbXR
r6kVsExCPkpBG5sa4WZ106FvTpcqkzmvA/908yVQR1b6qpxOhoL5SSfSzQcPG1+N
bCw28uRhbRafPBs9WWZgVpadcj0+08RT5lUvjoQC7+fCP+664xsRs4EoSNF1HUkH
tD+CIyBkGmFwqHni5EZS/YlC61HH5hZ3IPMEiCzXzo2hpI4qkdXU4FvL3dUWo7zC
plb6zgJCGaGmhrZArcBiNbCpRl9ycLJZXTPWZv3sE+Ip1mFF16hgCR+gJhviRFad
HMmfclTWKM/R3Es+aeE+bfDmfj1ufik9Mt6oexUHcbKG8dQB0L76xWSQDjcVezSr
JnfGmzucmdDRDxiUkfJDRAArWtVWJmz6VibJYmwRRalofvj/fC0+1VrETeYFfLuw
t1xyy/r/ZtsVPIzVN/9Euu2nX/I1p9IgyD+1L7eWSoxROdcHQkZoPpALm/o5bYnq
g/OQf9YhYdEykRbYijxB6BMjduENrPOOWG9euuvwRK117cHG6FidddRSwSJyefIH
lTFdSVI09EZkUnUw6/bqQa31maC76Sb4A2R/gkvcPS0RxzKwCOAIIhOBJTALnp5B
uwkEspnrkrrXHDb5oYSRMdLak5HwliaRcMflJ/3cnxetDBTUZUVSKNPf53oP40zf
pFtqRmZMTXvr0no0247TVkY4em4fGb0aOTjMSg0RPCIZ/Fe9hu7xEl3eNC/HvNGX
Pej44mjGOkRwL65cOcgoB9dT3b8iMzt9iaQ0uv5xoyojCreOwJ4ki58d8iFHHVaj
h4ygVIKcbFR7DfMk/UnR4qImfEqSE16aueGdwj+jGfDAHW7YFcTiOLuJRhRoVBbS
ar7Kqd52uSXG9HZwoausVn4woXJIJwfNmCNCWYKb74wdYYaQHHiKBKybu9Lb0ycx
yWgd22Cooy1YAWx5F2QMZRdeFB/EE1E57ldxFkJ4mTTrG14KCSZlzBDTnEwTINHk
YhoEfQIKpjPxVnIZ5bCmlRTc5kAWQpjhDmDVg6fRyaJjpS226/0JXhTCCK9X47Oy
Gwv6IkuLGKaFX0AQKZ7nOLJkDs+6dhwokjcMib214IRL5W6T6JJ2eC8XasvZQTuI
nsba8q2jsCuifV2hszgJN5LFCMuQojG+IAL+LN0+nNb0FeRNhS5tVUpnwiqqY3O6
mSZ6VR9MTn69gFng22n86JrkTryjyDNQB9GrMbo2cx1jkv9IhCekplVRbrscxV+c
LCy0LFDvbsONXpoBYIOW6OG32bvUpwcX3b5XcEt1drSPl1jcxSoE7Zqng4JcjX7s
DcArQiRUuodex+P9nI5Hg3uyYKPxPm8UsOE+vdmvj+yca2x38/dkHDzvum8ejpi9
MCR7MFwYJftINhxWmTAy8d/f/9cUIlu9+p+hraUdjVmMRMx3tGPxCKB0YwHwDL3k
yG6zHvGQHXahjrB4LJe6TFF2ex0uOQoHkrqN8sR6UQDDdXEy9PMFdAobX0o9VZMr
BQemirCP/mcTfE8uvAbhjtqDaqvkBhbvHZg80yuXtZhCDs68OUaLjdPgHbXIT7Hu
JkwiWmLGBLKSo/WciaFKaoa00SMHPJMbJZQYjxKvYNOaKcaMPh7bCpxifOW2WzjL
PoiQO941tr/Ssv0ZH8SQ+PoU+IAJuR6h9w65EUhxjn4LN3d/pCr52W5bI1tQYcU3
iVdEkNHqRRVLoMlFMolO8IkqkbhIwnTspOHKESvsuwjtb16ZrgoZzX24UAVVMDi2
MEO6ciPdAnHoe6eQz0hFENmaCRSuSc4tSteBRVw2b+3ga/+qD+T53wWGJSk0Wwbc
FqWZvCaw+OpPGjMrloj8N8L3HEF7oW98DPZa3knGlCbyEYAn+a74Xg6MHxWFvHGW
5rhtvBpRcUDZTrV74vAxgBoWnlwade0R5na9OJC9mXEjNTsH4IPetbJ7gkrMHp/m
CGEvChni0ujcohgyR+ksp4Slr1HhVhkZGB8xphV5q1QJGSQgvkHadQSPL3yHnYhu
tl021zDdPSB2Ga1WVjZLLbWURMklTt7rLK9RpaCML1lCZkesOdbEsF60NChRau9o
FBbsfv7A8fPfuH24P9nPPR+UothrMMlZ+eytK3hG5vLKbTRm+Zmna4sc4HB3PxVk
948NBKxflTRKQ6VF3kfcGc764ziXzngJE+RaYUN+9pJxRsyX8xTK4K3OuLSwto8d
c7dOE78druh/exGYnZRyYUL5IpJIlhAoLybhOZr13qY9XlyNCnh6QgH/L6zBxmP8
nwrQAeR/HQn8aFsG/SSuScmXnkUxOGJCElQKTZN6DiWf/Bdv1wtPrDIwwqY6gV+e
Ex/ujUTUIfxtZSCQXCI3fwamJOgXX0p6Wknyb64TTuuTwRDpOpsI1ZZesgRyH1Is
wL7rNKGpNwImKCn2fnhDA2uX3FF+Z8sTunggSijW0DMeUtnopVLqZVFcbRKfM9dE
pEQusEBdwkCDHZnqBwiDm+mG+Ea3OxAGQPwrXtYJuKIZMQ3XIeXbEkyknieit6t+
dqGCNHomDVyVO930f9SnRk/rkwiakrNcByWk134LdAmbADR2f8W9YGSRjL9yMQKO
Ijjju9wbEcEkp0GCwW06kyGFAi425l+fzfFXgsnEz/KnMHeEjcv6Ae0vcQDKgMfd
om5aSVvYccevh3gx+LGVGK5UiRn7inuT0nzQTsgog32XxIBSMBHfsPIxaRRLDgEP
GaAh1VgAARnhOEeM4VefAU6hY4d/Ic1Wokfw4hPdCb5535astfC7tpFc8U78psIw
R4+jYh6SEEAmJ9go45FHTePY5qP8y52wO31PSVM6ljj8ky05O5JmxWq1JYTigdE3
qSaACjRFeuQJA50Bcgo+Vh3pI1l6dAAi4HZvR0f7EWtXp7tSsp1ttXlFFyk8/u1m
dozc8z3NQj7kVJVhRBZiUX2xuCAPjbPNu6S25bBIiazXqaJose78yUokThUCd9xN
WGuwMpPbeIZxyjWk5y+sdLdnjihb3dukkvNDEgWqKwkBjimUICQIft8sT39WUHM8
wG/puo5rcMcihizzgjVvpS21/y6/vcHAi2wyuQU6H/weAiPE8lKAOMuq4PtsNkfC
AWXKVl61CRBO9xgB2/DKsM/2sEABidIq+8S6hoFPdokpH6Q3JVv9doLpvOuvEi3O
3/14GkSj1mb7VykT224wIQLilhNpWi7TVoph3tSNWLfPTqHOU0HQHJE5Fl1g2DH7
miT6qszN95tMpeFsrTNkUcxiNyz0VbD4KZaLR21flsYw7xccYHZ/zEX75xHceV2f
NZu98q0Z6nCkQzzaG3XTaPnbZ5zfitNhqQgJMdokAxHatP1DBwxA7hfunZD8QGvM
js3WT9yzYK0XAcwhVkOtGQGIHVvlyzP7fIzraIth71Upv8MYyMYqAeMFnaRS5qdT
cR6PWMJZnYGHdXoUjgslLfZ08pI9h/OpjXFrv9PQIZon/0vhcedVS55i8Zoi7xwY
NbAeFZl9wFoFlWXi+oKT4TvSGXWa775egi0xp+OprHcmyL6bY1g90pCZm0FHsDUx
sJFja3hyYHrGE7D916ALQlTlbZznNuOmrgLLCCWaxD8D25vuNfamN9brmtx6cuhK
v4EinCT1S9JXW/nzlvGFJFSRH5gxUZL1XlYzN0+sXN9IARwyFBnE0dOpaOt0coyM
Kx+3CJwW+0XI1QEF4K1pLWHCIP+TanNcwSsZrQUMgMJKX8wKw6IBYbHDGVCTqBgA
YA87XTLUhKGfYcONBfIJawf+KDfRZmDzxma0xbGy1o+8NntWnLWxZKrqlbL9aIVa
oP7g5yVqFk50+XvCTyC10g7wKVqmBD9wjX/d1KvTWyZss/XpaAWF+dnG/CWS1Nqk
9MRSPbSOnXGvFWPvwxne7mvHYQOm80bv89gdtRnx+4nXakf0c/yCwCeDMcIW0web
OID91CvzSiIokHRVIf4OTsjcFDSoF5MnTW8AG7XRGNOdG6XktYytHYBRyeGIw/mb
ypUIOOoclr21PoD+6gYzDJp0Uv/gBDSM4OZlGa7Q/H40021XhF6Yfi3xSAAQZ5hu
9GDBCTKNQ8LbP6j6lvaueWEziTwWcXEDqzewjTV42zokI0lVtChvqpF/ccIb1pBN
O+wTCq65B2Iu9h7rV7fnOZ6Y74Ul1wl/rR4jw2/KZAg2Jr+cU8ybd4BSp61nHOUQ
6nIums4pxmfrsyfwyTzC8GU50sNMl0IOozwfjYEpTpdU7ZiLVu1vurEWmLZ8t0cZ
ECN8wJrFnStgqXz/9Feq4AmQOX4/aC3iRcN1ggRr8aphU2wAan2IW+smgOv7leYb
baK9qtfYm7uOHao/czKI8wRDu2ULdh5nTfq264iEicXkQI1fEmLpEZa/67VTIyP0
kwXnI6l6YqfAxJJTEWSxJKxRVp2/ViwE1EvmV/2Tt9Ha9dqfcNBXZeS4o699Pao8
kLqVMJGvvDi9U+Km32pvoRRklWE1mqQ/wDIFxVfg8urQpQxt+/FUNctY0IAIyPK+
V8dDGzOr4Br8ctKy6IbGmBTTRL1CNFLKEusnQyfUv2p5oZBy5d/ryQwJhKIgtshZ
0/MhjOx8LUF/Y6ixcYlZEG0aj6TLlA1pzgbFGZgmkqZ44v1+5FwfNuBhYFfBYcjO
n6jXQmoI1jA5QTSSEJT/GXMUlYAWVYB4zk7lQIhtia/+sQ7XEvFeKsVwH6CoYNsL
WKZSwwqRE9Hsk96IUZPmw0fAAPsZE3a31TDBugy3mEGiRpMnwpJwFR6BRhNnIIR2
72TCPxF7vpa4A+lOjgo2+j6UNAeI5c4qU8FX6doyubZT0GKiBWE7OBs54HgGdNmT
TCyxLfZrpeIUNZhXYAvqMoR5bdUQeXv34qiYMDa/6NWA8+Qr6tkPuQnNeTAFrJqC
Ahnorgrqn5AqDqRdB4OYLFF/S4tDbsUMDwGNhRwyD0TwKx+RhphL0HDjBa6ja249
Aw58gtNSSjaincxETqXjobFu7cxeAOY95Lj8dcdCGUeLpQIJUgOhChyrXkA+o0zF
qj4xN8847qwVBxtX45fzKf+H8ZB6h90XonGG163+rE21nyaPxlq2wVBvuaHC+clt
D3G2LHVUaLzGnh80cjJhtFsQ8kLPJKZW8V6/qaG0K5Fqon2qUlllxZMNWe3UqovF
7O5X452+dKpDU3CLzZxCDQyricTEUOPmgkn/aiCvl6eJTEUDOdmhUQTffSWld5Tz
oo3U+G+C6s3Ayckx5Qg+QOjG/pKQ+M8msoYLmeClD5WWOCF5CQ1Z+/GtNz9Mc+7y
QadYKOeTGv/q4Zgq1YlaEiWb464pGPJF2+X9XDlrCWrpjvs+HyI4Vp79BSmW7Bp3
YuTtmYZ9OHR5WQvWFrAquRDSWXzloMPO+ep9J3tuesdcKys8fO8oRYRJfJXl822d
O6GGoKAVGt/vsmhvbEIbPJX6qvNuni5Hj2t8cmUvn4ajHCGy5x68kHrPegt1Fatp
L+1BgWHGlLFVTAx1lDDGBjL1aU1OetpToaG3t9BUe73Y31ftdDoJI5woW/UpwDKg
0WQqK0vPr957WjDxAi0FgIiSkvlE0C+jTtsMN6OidxBq+UadRj/owHn11PISBqak
Th6ZTO/hWJ6qSDSAHiiHvo9aSqIIGw0IRP1SGCNkDrKU1MwbxOUFsemsrNnBNs7n
VphMiqoPTFnNdb38kiiCo5UHg9X0c9mu0ShyGlLDwx8PvdNwka7PFRGxXKhA0H4W
cTWBFk/Mz4WPI0W+L/VVYI49AX6ofkOUlabPeSiW7yYFC0XtilN+JRLWMKcyPVvn
cq+n33QpTXkDcAyuImE8AcV/v2BAyAFaPs2nRW+9JeXdV3WJA35vKlQXJyxGZb1P
1XMOhOZlau34NKLIyrWGkrSYu3bZLhI2ahs0pKmVkn2MZm7UW3ZlYnB70GSqsNkT
iXXli/anwhXP39UyuWbyJT6J3/OOu9ZHofSf+gaEgTw7u3mTh3eQ+SYLE0THuhgn
e+RUmnJW0dLcZZ9sOorFiW3otjtI4pyk1P2CkSqfQwQ9Ic4Ca4YyEt7ke9KSXEBK
zZ8xJj8r/TCgfOWkoJNM3C7/GNKXvC4XJKxs/mKu0GO8YFWWM9TVFiahbiIngbcU
ZUkdvXKR2XUS+WKjWpp00GMIgHPMy1xKo2n1ZZ6KcseQAT41u8rt4iiO+eaogu6M
IpXgQyZ0LFRRsDylXaaK7dAj9WMueyZHrtWJKdOLVL2lT1lOK54JiJ7vnanCborT
3HPiEQyfGIN1Kt0InvFPzAXJS+njoca3AeOYCaflaq3jCTDerfrvXS1yqJTqrju0
E1THaMovlqPwZ157h+dNio7lPpoEUPLR0v2SlWjEMfNF3x0tL+znNuEEflno0AEZ
4xTpObDD7OFSe5/2+uvg654IssTvkcEI6A0byfFnZgj0n0Xm6EIpGVtthKo0TnHf
+QpvZBePdTEC5PeYQIhxE4oEqCT6uDh4QrgHh7WOnM+hol/+5vpR9lcGUOjYTIxb
ISBOBDQOvs1oizoBBTp2FIMECtX2ViIzA7jEYonYMroHJu9CYhfoymRWeuQyM5Sz
ZfTdX/kc1pvvjU9oJHOm3XbqvYyf+HQcEqmTxKqDAMCmQr0DKPvAJdiRtXar1Al/
F/lAoyw9YN7XoCnEkN/8Hnn2Obz68TkUa70RE4rZ6o0Y7YI8vnbjDzeN0n3tcG/H
9KwFl/bKovS8f/39itaLJnq0h2X2UtaBNlpbSL1j7dSQGUfK19AYkq51UR0LY739
xEEjMB2b7N+E7lxfYh2JFR1AQuSoHOXn5DUoGxZKoNLenjjUcsytvM+g970WGIU6
dZKgcLan35ED7xOQPK1XNp+jIO9A/19G6Q0dGP98JnbWFANfLZTmxvvQZepEVTNF
EIMzwkW9gR8Hk/rBag0TbcuJp+5BDqzp/ipGQV7BWPGsTo0sdyrjvpavOqJmSZsS
ZFCVgelRMt3K68AmJT7NHyVjt66F6Gcugi0F1Z9tPQoZLDHeK6Rwl/9WsXGPzHbF
nTf9tIUqAdqDSHjUw0FYwVU9wFBYlEZePPsMx9gT8uDZyLmMIQc382epT7bk5GxT
n83wbZ4AZ9AsfCrp6jIvkmGqtsfY6qOW+IQFI2VYnOVmHpbUcJNc78NmM8K6YGVD
u9hEKmr1NmQXwlYilojFTvKKqZiT//w7zyKtf68cbxtr1Skv8uBTXAXwE7Bb+pg6
gv9HH+6I5sWDZTen6AkltyJrEDr6adqkMqKDUQlaNyOsO+GnLKzyHdzG0i8TOe+i
pqzwctj23QPve132MbuAOpdGgXjoDz4tYCVk8mLGcH1GE1DEYFhNnNycvc3b0dd3
5NPABpyVwT8re4XYs5HEAfGfCjcjsGT5UtjaI/gKnise7R/hFzC1nQHpZ7OHZsTf
57QzyVVhHSBNk2KTV2jlYxDyRWUyhPAo5YNgqEas7sxMULBcobtL1ZsnUIMBVksR
GlBe9ZJxJM1ocb5k1iwHl7c0C1NuEBPQum1VL5qXcPAZHXYXPmpfu4pDgeJXBHkt
YoU1nEFhf1dbclAb0uz0wn5BblxN3kgBnpLXU/NRE+6oWKw75Bira9OHE75oqMlp
JKcAymU9zk6Cxr7jR++5X7xofbd1px4kt6bhIL9LDVgGvOVuLbnVPtuNGHWK38K1
cUqGvjBVx01Se7CjaID/W/AFaPbucFohpGtAvk4KkdoLukebYfZhM0N2SD3FBpew
Pqvx7boKwoarutA6+JKV1bhlwhSq7ZbDIsCccOUEIDXhTvHP7FkMMoNy/6ssERJl
cmmc7Y69LoUshmuwzVCQYIedLUitorH6KdQtcDLjcktkwZMYpwLHyRnHY88JmpMH
uPwxJTJ/3uqlmp1rvZBuplPi6jTBuzTOcEQg/QcOA05A1FuDOSRlH325hI7q/MVX
8w9NOaQyMunJ2iCf8AagdsmvpnDdZFlv/KbcWLNfryGCEHZLbIuNNy+JBz/z2mIj
bSx9wOUhp1EAxQilbMA/2JcvtdRwFe0/1A1vAqC2iBQtughT2iCFe+JsSR7EmV8N
YtapUatzryw40NxTYrYtN3C/wXYDQ7z4elQVF/4KIfi2Ugd7RAvWsFvAnNiqmaCI
oaihmVoBL9Dnd+NaE1tZvcLASyARdmoWaOZWGcSWL2/NWLGf7ZnAQLOWuD80L2DM
pFjSZ+ZHU7jmKvfJEWMbro5Fkul8plxQAnv1kwQTX1eI23jIk4TeSLgNkzTQLJm3
XSMgVZRWNVKuZ5IGV34GBZZppM5rwpQcSV+Wc9HRLsDcoUepxLjZBsdqiVbo/19N
xCt1x4AhLSLBTSUorMmjiq5OfQDYm+JfOG+VEDqJ00pSmrIbxwp3iMFvtcqvSARh
28qzm5zqydGhNKw55xH6raR6/nREZujABmoNOzIZoR9ceBwrOz6KOWJak/eegYhr
0E6d7yk6jf/0pmJdUxjg43yCHjinsaBAch6fYGf0RS9Z7EIA3nevG+Nrw9BDPs4q
qsxMOoWlXjWVg/WxogkoQtIukanE3ezG/b7Hh8U/G+3A+4Yw4uaGDcnHmUbuZJ+N
GDQyTAZLMYUbMYDqtmrordcFMkFCb3pBTaDJK9jzjscocrujrtgikVmWan9huEWG
ySBhMwmpyLS/U4P+38j1OK68oYGmavtNyhw9UG6U9uLT/3Te4dxvG0b9PfnfApAQ
OdgqRcb1Gnkm/ZxTl31pPqrLg02KO2RtJHrmrWR9sAMqDE7ilVmnuIRaV5GBE21O
ECYxWgD6MvEigy+2fPOomZVI4vv4CCsnTsdXOljGAY7Fu6Ps7wN7LCQpuQrq3Ihg
REY21KADR9lmjMHFWjgDWgq09M7LbK+ymKxz8gETkRHCOZ/ndtkhfBmmVwJ0/Wp5
tjM5HWzonghzSW3hkabb9Y9uDfSpLXbF0Sfct0W7OkI4KEgpJtoX8xcdhvq0SUvA
DVxnSvk1u56WVx9GGsyPFnAx3JwoyjbwqjSqGZr2JtzOHog61gdDftYXTfIzjuvq
BRPJIPA/bECkrQmnnPmh+DgBxebYiFO+58CgdrlOJD5Vl3p2kl7QNvD/FhpSYmoD
jYUnAij6uPWqrJjIsL0spNKGYzRwHP2VzVqRhOLUYzVKCxPR0D6y3faWQx74oThk
66hQ/Q3KDs4H1ShZTxa5pPSsRaoVNY31/fkRV+idfts3pgrS3qeCniSKi4kI3Zfn
XN9f+aSmyYQdlehEdsaCBextYUP+dDtaHUu5hM4kd4lzYH66x5/e9bI9rH4zkFEh
uo1vbm5et2ibU4qHO7uZSG2SihPdwLvLJKpgJGxI3B0Oou/TOFBspuNeK8bdIbPw
I0EVyrpeNaZFce2WuJ/UGOrdVX2k9/8MWyR3Hepw8p7grQ0iwsqsDms3i7/3nEMD
/cviJFRg/o9UkRWlPIEiwiOXcpIUBJjugGc26zabpJ9WBHcmgYPb8i2XYdijCvMU
q8B5hGl7nY5gUKVCawn56/Kr6i78T9W4oAEShshfNsjHDb+neSgs/+uiHzA9wtIh
q7/nJSffErwF1/Pz5FRWfAcXRJt6YMjS4fx+cU490UaW7C87oO4LU8vZnyLol38C
X3K4wIHe/X2i6YOLk67SfQjje4RJwQOKEgfxMr4UbocgYfN3XpEomMfW6oL3ZZkO
X8DZoqflFVZBceFirXAF6I6TdtDV06H7jjXeNO0/pOg4QZeAuv+J88ijMq8Q2sfc
I5JEOXeeIKmPWDCEizBVMnYWmajPMrtmkkETuRmYM+rQAO6DNJxaaYSFhJMZuIJ9
yMJpYwHxo4RXX7x1kwJJGh8qbNhuDGXjsv5YRFXUv9cIo0apZWN5yh8P//oqCeY3
Z32C2pvgPI08iumsanW+VktuwH3USedZSRzQ5CA7g3NbcyM3LH+yc3TcOX8Edlpx
PNPlKzEl4Bh7vDmrIOi6gXzzUh2P0VH5p8vCTmJe4M+BoCN+9axxfM5Gt4RgYHQr
RSUZZuUduCPAbL+QY+8p39TkHgim2nE0ZF7JdLbUdm8nKAyeKz7fZxQphAr/BVtT
xbZHf71MMH3z5PTLR67zUwnLWnyY7srSVvN+LUBr/jIh2E1qrYcwLmdyVr7o49Wq
k+g3QxBeudi/fSsJK60WzXtSv9u3gvNu5i3EZ74WcSwFvSAzeCjX+QQoiLFCvyqn
Asaq30KagHLMCkg55lCX71pmDKygEMV+gFOEXDN5KyZZ3JaPYmGlveCo/BVGuN/M
ixGRyw/zef3mALojUVMMJ7uLP85nCsa0wS0KSB2V43ArlPsjkBMsc1ivFFU3DAEB
MLOvMf8Qt+5i3Seok2BJZqzKv5VrBmN3rHqNSRNpC6wZ3yK6997dSAMt0I3kKI47
bHRsBUJePWXMkTF9bkNCkBfpsNxq6i0pHGOnHldLeHOtbK717dcD9M+aGVwo2f9J
GD8rybRo9FfEu2m03G4cEkkOagh/nMqgf2QcNx33tyZ+5FF7myS4bbeVCIun4Lbr
XdSQDpXEhpUzMIJI0Dlq8slxvfbS+nsHPQXHfPgmAUw2goyqRxfI1+a8szwNUf2v
W/JKdLPbgTT9UOY4qbr7CKIea+D+fRhHjkms10z/3FsPpHkNiWmyfQCH9BOyaMLd
cqKqak+w/hGKgCGSFiecgdKLlx3cWskn66xOY/2+8Zb19EAK3QvT4zDWsh3TtLbx
z3oR2n68Hp+SxRAkHn6x9KKkBh3jkWiurlOA7lhh6SyxnrEvUecYM1UqfMmtX9ZF
BNvV3pqVy8Cvrv/QZlUkNqM5kISAn1xL1IvR96iwxVzs6rKnkacze+5biWndtlkv
Dl8rRSyscBGDcIf51QVp2pJMuGhJkF4d11peD8PqkLn69yZyb61F1SIFymfctHMY
oVtyEAybe5LhW9GTDZLxfbUXxmENja8hnhJOFrHqCJM2zrt+u3JAn+6aKFCB4VH+
xdksmwXXew8GRgvSxPupPM5IXKayl4nFqqrDWNMxg3270KxY+G3IWtbmIyOax+8P
ZpL5O0K3ficrSGI/QzoOP4ao1jtnztmmHx+R+qInmp9vmXE2wpbpv/qf9e8gCGpY
HMjlP6XYUjcuUi3rHNLzBoEJ3HyF9BCqOcDtmPAk2VVO4ovhBLXd4H/crRfa0/nN
LccDN/hV2uHyHXW/+hx8xgDLz5rlpVtFE8nPBcbW7GtKoHfgJdZ0VwNtTWiO/4Lf
tYxAvJkDZMsmFQ4LlUzUeoImlFd+z7/2dPcb0dESkd96q3WHF2NR8yapY1wTqVgF
5Bonaqwty3PAgj9FLgBWX3dbw7HF/7rOdDLqPlut9PdD7At7lscgbpAEbDLQ+Awt
rt+CrhiIpMfnyclgOSrwF4wy0BQloOUhkocqjFtXZgFb8S63pMaWY2VN9lR9s8oP
ifzuwCO+7y2uALjmGxW6KCylxampz/KTl2Ri/Mw9rFXGn6gJc9PzBGclWWtRZ0H5
2rNVlVVT3snSCGgeSodKlsWsrMXI2QBzjC7IeYs+6QBtIiruN+P1ooaoy8el5EFR
sTD/Jqe6iiTU1Cww6Z2nL4evZdBROfQu2coTp+gwKebCj5BkvkslapgWOpG29ADE
IMF9Jy3EQZXmgeQLNSoxOYYQEVcUq7j+c7c1HE/jagtbK2GPXgN9JnKuHixGHNr8
Ps3PXvlZ7UBHOrkqgYhJsUPk+ABJyjNHiiIvlMYrxim6yAEGJ5bnGLDN1J+Lh4rM
lFuhviICS4ZYTzFCKO96EjRLD/YdSgk8M5ujfMDU/tZQnnDP9YIAiWTXXcfRjOPZ
aWvWepv5DyIXJskxRMohFmB/5cjDVIb565e4DovUER41lyCkyLKE8N0K+fZDwN4Q
AhHGRoj0o7ZxvFuxatCSBNYCZDN8NPuqYLBstvnbONbWgiF7Df+GBsrMb5Ujwgbk
dG4ucNr3dKFEzpE+MZC6bMtKA1dL6ueulG6uFaBPBJS74E7QqImvNO1Y1H3Yu3Ke
KkF+801ii5IxhWTFTJgG/82tCUPVgE1IlY+x6N/g5Uaq6pZ732xgZkciUwn5hMUp
x9qzv5kF8HZJuJkaiUzlC/fJ7S4msG00+wFttGQPutayl/t7aA/BSSAf45ixU6zg
0FSssydIpjj1jVtC6KrrgBHVMGwS1VeFEbN1RX/LWfyGWuIvd/30UpoMAwiv8d3N
gl+Lx1/Z+0KifLKrF4J5r/0bOsG3hGRCjOmPUHem1Rhkpxx5JUb+PPGj0pUe5CuP
8S0uRg6Cf1ErCyOp67TxQi1yZE3zt2JmR0BzdEDfmIauf/1y2iowHMm2ciUtP8fi
HvBJW3NMe2BxuY0TTp50FyuX608/WrIpoIcuRXNeiRV5Tmctay9uubCzBGrGuY4Q
JXVCL2dwzV7REJgiEatvegHCCaefC3AOuy21G0MHL17bKGX+VcNjUGYwYvgkix/Y
0zZli2yomrco7LMreop2tMHCM34f9sqO8Tu10HK6+fuV5IBtMaFYZ/C3wgMQiVee
/908jDp+wLAuDswYMmaxPzpYvTSNsaDHmOVVQHevV+1hCW46jy9yqdz2e/LUr8uz
AFXcMLhscCXjKLJzN3BKZSklG6YTHlj7bIc2KGe/JoXSoyU0NJ87lWYGYhju7LIh
h5XZ45MOSODQZrsKHM29jOOacC/Q8yVfosYepUUlMDnOJJJu+mFM9EoPdVe6r9vV
ZM3NE7MT+7PBkXfCDLUmHclPUKzzkE/8yNeQ/Lm3U4C5O6bveuQAVAAnWGLxqOoA
8dtEC2wzu64zfM/C7lfd0QqnVX9ZsYi3yvtkw4FIulAdNzni9aUHoLrQKA/4XYuR
GChT4eHnV70XolH+wpRQvvJWn3d3dnZxLTOSJWRtmq/OmLaHFFvwCX6z5jDL9q65
tj2TyI2Zx0n6C8koeXr0R2PAHOfQuvUFtYCl2yIo+/WcI/wEaVcVWbIdoG4hMgLE
srHUaU695kO1jGE1F78DfCp+CkJ7XnuJySf+/TFAX+JNbrQTj1pn8aEjpInKhXNF
BfdAUvfyW0FnIHuxJ5b10KWParfI9FM4J5DlKhkP2B11+u1ILAhkBjkYDc60tTs4
tdU92KeDeSoCwx0u9AZ0cIzlacgXg5LP+xMXUQb8uiNOM2eaYXmizfJ8E8xcJAY5
NnywSCfl0bV8JS/4Ksva72zcwoekvKCfPolNNIIKcFCWYLicuNopMFj8n0+1Mjuf
svOhgEagii1BJdkzfNixRxOoujtnkOxgxim7p6+AAwkllBJwOlE/i0atEEp7IINa
IQFc88h20BlXlAZ1PKd85r3F/BZQK1cW3u1LbJHKWKn1DQvXNtwqeQhqkpZxB+h7
kiovd+ziA98bYkiILpmc/RpfIbqU6ZkW4+GwkirrQjZVVKJePJ1lUfv5aKbrR+tE
fV52JzFL7sAc58UnJSRYJuH5P2zcvg7bvoteAh/CmnRDSp6FTQ3IHXvsnsAQ0pI/
1e8hAh7ajnQWaM40dQOw+cchrKZ6TCLlKMk9KB7TY486rXqfoN+d0sVqnqkuywSD
Q9WbOFtk215PtG8n0edL3MOw3RWKhBYlEn7nSw02rDPeaHrMI2SHvL6Pw5bPRd6i
WDPVF19sB3iDUGmWS4vVZ1jTlbQZayCo1Jr9ZI68hVIinsjbFCNGU1+xSyj3XMt0
c0wJeXXksBYJXN08q9N4imTrw2dVUd53+nbJgK9IjvMgT9F6m/nRCb9WMob3CDqk
OGsmXaSt+mC4xzlTjabDz4p4gW3jdhxuLwS9otJRczutRTYemjpeC/a586HG+kKa
/y9MGonpvBwp2ZZ0V+7Sux6qQ2nu9RkCoSDPMhDIKrIjVRdATiFG01ypABpIj2uH
iV5GflneZMSxIsNS9okzuDBlHhLVHyi9iuWDvdUmA61lNlqV7opV0IBYvJ2USo7t
6qr40XZU1C0wAixEMno3x5iJOgOJmCs+gxTGRktkHZDnyNwPFsXE3Qr8RRXxj/M4
3pXp5Bgt5SIBMuGkEfPGRDoitkw3taWjb0mrm0SuCBGgeFxj5xCeFk6l2V1zTHA2
vMJX278cil7hkeEOu6WEE77C4b1odfPFCIqDB1R8wXGjge1ZbsyuraJcbTMvVjTN
s6Tkl/KVwjM0Q90ti15oAq4STgQ1xRyn9MIOsXRIBZAamNrKjGhqb99MuS40YGh8
DaGOvg8eLIsN9P5biZC/VZfP3OWJi2y2u951HanXYtQHnQoq/YrE4rXhOf6onsIu
1UVZ6acY+Sy+2i1Xc3ytjVHX5hIEyd49/xdiYBJI5cXj5ud1ei4lhD1BDehZVHFd
oIKSVd2LrwwnCo1ojN+HXvLCNEoRXjEK5bnus09gRdkLCnxzYqR7gIHJJwpkAuPh
36CUTcqbD7PtMM2rWTwNHEJfbOEaaknNpttrgtt+lhjALtYzAX3iRyBGQOtOQRNq
djik5nFKX/fsFe6BTpv72S61a/5cQzKfDAwxSjSEkO8gHv2222qO7fV3/fSpSf3L
WlFJasaaRabv0FkQq9katDzcFVWoNEP5MMqZAAmYCkjva41/N2YEubYWMvlCyDPv
/gQ6c5NxMQp7xzzUmHv5JQolrtvMZ0aQudVoC4JBqJ27GEOqJSI54NHV1gDvcIym
cvo+GU/T4+wWCa4Cd8duu6Ids9I3HmYM/kT5Jjf5BlgMVrZDyKQyovN+oLYS1XoG
To1Be0iG74ILUUev25kahs+PWKywXQ9K4wd8dNd5o6vbFkyaGs4WjujXoBpch67H
C4Wgn+I1Z6fmTY82bRa3aYE3Rgb2HV9YRxjlcaqVzkb4fbLH1FyVcR3/6Lyu3s0Z
fH5auW14qBIbanRVHtXDHYijRFxV+iE8AKNK8DlrT1PUqXJaqbCLe6utWb9d1Uws
dEgTFb/8m0/O+rjXXaV6WXGdrjvMUWW+RRm7tX2jr/ILe36VfY4+ZzstEpBHL+RX
mUJ0jK2cVOc6494gx2kFwtiYistKltqn4SfCzy/SlnhHLvULKwO0li2xismotRkH
aKMR20YSCDgSV8sIkNrP+mFGzQ8CvIYttsIBPljL8yYRHp/RR+1WP9j3EyTCwAAY
6V0lWbKaE52hUdSNby/9VqTr0RAVcapesKmcNJZJuklFWZKOyrBa5EPd7egPpjrm
jHntPXTKs0qr85btWWQxfiLI9oVVJ/OVeAAe6GkAiK9KBUcuQNZQEclR7vSJad0+
SMf8fsUbczbTip/GmZWU8seBJNg1N0Ui44W/4iwtfNfaoFPHkEOzP6/CaHfxYGpl
WTyG7Kap5D5PnZHsskcY813KL1wodjMfxCWLkPeDswHjiAHCsIm9XRasyoflTv/e
7CInP90pl+JGceXGGN+Tmp3kP2kBiUXFhQckDQzSwLnJS9PYsU1XqA3jt9DB7Apl
TmMLA6+P5xz5dR0AWrFFd6SnsxmxZnZrw9jNy455psGHW/dma2n7vOquVulNY72N
rEko0cJkFPken9KjQcsStLVDRZwqYWJuaGwxnqCShTj3inYERbQX0IU72Fj6/9Aq
sOoWAyCZAWKfpfsoLUcfG0J646lg8fgLATfwACr1bJqhUSIrx0V96ZSbxtWSS/r2
4mC+/LVikgUl7EzPFjrAQB+u5Sfiq7hY8QiPUdnCgvjFSi98rcWBgQUe4bn+6E+X
vJTEDONhVEtFHQdO62vIozaFojoCOWt9ZbcGNP4A73QHrzSHjK0qlbjrRK1qTT58
bvEPPpx17rNUgOT1vYzMUNHfuTSxf4xZIypRiLQ+gTpV9r+kokIKiALe/C/pPUXJ
B0V22GRwIRzUF+PxbYcHzoMj5DDXI9awGxUvR5ShJix0egnDLIS8IWGhtiWvGDEX
H2j7S+YUh6q0lErOIzgA+B7ebTYf0RZ7OIJT6I56BhmEGP9X3GwyUMXmvXV0eNyp
xDbHb/NuHFaYy5qCZi1zdglJ3SOlLh7yzurp2fTjO9rNwaCKiyDARbwEW6riwwPW
rDssrcJVE87bas3S4P14XieMhxxdqoezeGGfHYT6WfkS1DWRwJlcuAYr/GgPbs8v
vPGago5JJm4cXgHUKLXOz5WF1gePu5pbLHijpvUjsyiSLbcf4BBlvzKIVO1A4D7e
73jKTkp057QRtr6gYkyT+8Cpw4IBHnc6401PqScDA2qToGFPmfadDXHLCv8PKpUx
LVARyUIUr8zvFxctG6cP/+Z+Gvze9eXETfgJxe6o1hoiYOyHZo++4kycl8ZPhQZ6
8vJSv4XureSTnb2aL5wNLJOXW5bhmLfhj1b0a9fP+wDCIdMgG7e9WsjKmaLm+rki
D3go8GFv4WRGdjcZ6icsGq7DUwZjGaij+8zzBLwJgb+o8pkh12k2ATLbn1gyDiEu
ez+B1EsnFshnzQmuDSFz4c+mjGwgqfht/Ydds62+06yOY4AR8rF192ZOJVBQuEYM
LzjfNFdbnByTxEIf5SYvH0WcU58hzA9BjN3POWHw6ThqMSiH8MRzYYfuhP9BGP/s
uYrBYvFhdUAdcLyLYu+Awx8XfNdw9YhKldr/RE0B4dl1orS9Cd1yd+X6IAim8WDn
4MoQdqVUL0SNKmNiTQRCj6ZE+hNWfhe8bptKnXRVCqiSkUa7RBSCvPbsty/xKolB
iOns+Ms1SyLO7n7he4kXB//61I2KbR3oZNE0g8iyTrAXAeO2n5jePCvCA5V7bsOj
r2KTrARAhimyjYK+UPpEyKXyLqw/fS737MOuHzaSntQAlAuoPqc0YFCVbmyI4orZ
TnjURemyUBPiQsd2hmeGD0Qg2ms5Zfsqk1nQfACXe0Xhbi7+swf2yffn406RMVyl
HS5FiEYi16QOC5L8Yotjt0tIoAMdbhvNe//RGmd8jlAZ+HX2vAerU9BLhs/9AuRT
4RWGwZoXnTK0Ei5X35Akw5MFnDAL4Sm1RMcjDZRv7GozUkndbWsQVJ1A1Anm7eZZ
J6IqWhilfZbFz4rUKif61PZImfKETsM5vw8fetVsj02i1s/qkZ+lengmfXmtpm6k
QRNuLKL69H6tISmbJj+Ujit58rKe75DgL1K7Mel+vtm1i81IZzwPmD/pWMk2rTXF
PhPvn+gw4loJHU2oSJm8WyJu2a3jHL2EiCfq9MOBviUKTvXhvk4IWTSyeNIIXn3c
02eslDWNeeJAqs1ZojI7/nefcu/dRtRv+3WeKmTsxMmnzUa3EKIxyxQi6Nq6pCbr
fG5PBGlNRV0BvYXo+99jTxQKOHndbkwrb0MesMoG3pnlvFc29JTy1G8gFE+i8CEB
KRZyf/aeQwG4z1rHnev0u4Ys2v/KepaQzdggOXhWVr486ifDa55rSfs8TjT7rBs/
2HX/UuYt16F5KNoONkGF1YrdMrckENsjONPLPkTB4DlQJ3NHFINqgl8RNkMstymp
8xGkHgzeBONOek8HXHK8kkD7uFU10ArP2eHFf1uaIr6icKr4OGJ6QPq1/ZOfzfqU
EDSnVnc/SV+nsLb4fqIejS43nd61abB/Utmhr4FWUiF1MnFtqn5F19nfjIN9pUGx
m5JfjhaFEd8Q78wtl/jwj8lhBaZIzhjV1PpeZIXY+dDow3kfbFNYzaT0m+haJA7D
rSmUbDcHbbJY3v0kXKanvehISxB1oeV+PlnIdYbdvxYwvkThn6p1QUp9DoFWYTC/
cS92bSMmV8zv2sUcvDkOqUYYL4OWYRAqAUFsc44ODyx5Q/RqPDmzW2hI29LiUGkb
ADpHtNyIjHjiKpkhegxiEoPiRDuEheylpnQDLI2mIEcXWZLaQAZh5MiNOwGE75We
p+22oUh+CvAf+6fHRDnDdw/dV4CGN5sYGNhtZ2EZp2Bt0vxCZuFz3rHMOY48gY5x
lUWVJcRltOxmoe5Pe6KhoAx0FQ4mkB1OImRfXWtIAWy4ycrDX+qluiT2EXL1Qpe/
hs+Il8N/y5ykMu/KZJoA2RMicIwZpBLalvGwef4a8cn3cVqrFOCmadeE0QnIp7fl
4aCrhPYit2hl6dJiOfTabGNFF8M6h2FSsk2fyz120758hJdTm/LR3xWulkxKcslB
F5yEp5tmsKbr081gKhRGi1K7T8JiK2DhGcifWbxNstZ3ORJNQdDTrGro+a12HHp+
7wLmF4biYGXho3NvRnRXXygZCdBFWDINNLfO2WPQ+aPoj1SLEDnY2otMTI06p38V
j7JRj6YVxgTPn6/Jp7BuwfZxcMLTfAF0ZlE8/TJikU2YrAJIxN37jeSjjeU2wvrq
tND4/pO+Zjk1GZIXoudH3+lejR9IPpkOHWL9vZcVUrkjIUVMUQk4IQWEQtCqa4vY
wiSH3mPLyjeuUHoYRdAL7d2at5kfBSgAOGgspGBHUhvAbMNg64V+IrKvF2P2MQdG
OW3htxMkJ2zBZ8Ux+LR6ZIUIRBpuCMCaQli4Vfr0ZUeMsigbEsqaRuRxoHtuB6lc
sb0Ke7QrWCQkOF/wxP5p3NkLrl+Kma+DhalMvh2+fp3IJHTFdVJb47Xm2EDf3iwE
C+2WuhNs20FaNnK07ufPeyAef4t3A+0i67mDtJcRxhrXTftU55C2GM2XKhrdX/V+
YLLuqph3/dcp+2IWChN3cze3wuhzlKFpcix8pOJB9915aER7vyFVgsihxNjFo948
IlAIFc98T8OSgSh1x4elNxmuEgsVbc70l+0UAJTza3CQnd9DLhD73z76PI4Im4t5
NxnH04b6GZpmXSR4+HSWye1g30gulxiv2ywSs8tvrAEXewNqpgTMF4qhNA5QJB6H
m/8DEmVm7V1aPxN9nHXs9+I2S/LG0cBL2xDEZgosj17pqUHQ0Shtnjm4FVKtobpY
KU8hdwUdyln2Z9erQDidXDpO7gw/KFsne2c1nACiOahJ1J76aoOOc3tUIJp6Ymb2
/9/ckWGle6bqkQivaWHTPsoX6ZNVJgfMkQjfvPLeqCCu1cctbG2o7TMGmQkTqp5H
8c8dFpIJXYLF3iK3/+xtBY759VOrbYi5CJBxMhMWftkwmcBrV0IP70mHezX70b0O
AOdmDdGOa0lHWayY7gQYxK2nJec6VrloAeukWmxuMnP+nEinaRJgX5TAv7i95kgg
lAE9taREZrG3aWLYsn4T6XcA8fEpNWPC+F2+YgaAKYF9F9nm0k/WUjVCUf2hoG7Y
NBrfPa3aE0RKU8ymYAG7FvuoioG3Rx0sS+lmD0SZ3Y5mZeR0JWOxAjfMNYfvr1Ty
h8tvmQ1vHwtxZhkP6FKhy5oCfKIurBxS/aIGAlW3Cav1b6OJVn1S69R8LOPiJqLt
3uUlsm1XQuadRYXZS9RE4FJM2ABvKq+3ew7b2ynJ5QxkgVNamI/wj5wV3LYHJDT5
cmNEwDuYQqKUmDLcv0zxtbwi6UzfOq9GWcKsw0KtIUvM+g5KkzRcArorpdu7G2Nr
3EPMqm2SdhXTLMsC6OtRQS0Bw3hdFdFt/DC/xOxEYmsL0CavT5/Lriu8T7SyZnGM
bqAZQtwaTGTnAFaJoX/mMP2ywf5Tug9vpkYAjJBIfehIqB9HnfWiKhPCR18W27GS
3erdEx9yZFm6HfC8x64D6nb/wqDle2mCyLwh+pu1JA9DECvvD2+lQYh2N7u5Xnur
Pba86BrOhKujrPGrz+brwwnhvY+hQiVy6MiZDrwTbqcaMMRYA6x5bAr2S/boUapH
H0FqB1Sylhp4WgZuDqOOg/7+7JtJmZJsJOKQxvvF//xKbos4frb4nEjW5PLfSHwc
sQiNtZpw6/cYIKm542e2/cgJom87PzGnFX4PYkqL4LPpAp99IQ7Iv3sk+lle7BoE
k8BGa1RI+Mg7IkmXSCAqGe8m4aCc5mHHpIqR/fU9sjw5zC3KaoM3otPrMrEUSdVi
TWohvVXjMSdm/8518/rE1cAgOcdokAx+EeeP5Hg7teo4gPzjUZ4HYCWzg1Ov1g05
TBTw+QHGXNWBm6bD4Y0pRIsnxdc863Uwj4pFRMDTfdAP6CvfoVy1Um/GKDYigVXo
5M35TvBNfDYz2EhOAYJJDPta3qknOkhT+FUS3Rkal6R9YXHpalNmjonlATEgeC1F
onRF71Hjfx/KsElfmkAu5gPh+IIkOSpL9q9xtHpEPHIvEkdsKtA7BnATAAlTFSkv
17q2rQ7k2tOuXTAekDfvjPlvZUd31inyo8NlL3LnYSSHcyaCctQVVjxjse4nfnlB
IbO0j+8L03kaR4CTeyrRsOOBKA4KJzXtfxTr8n80cm2wGJNGDE3XaVkEptUX/TeY
1IOgNkQtZseueZHMpArDUXMla+vtCQFZMfU6xebAkLle+Wgx/jKuwA+4vPx2l82l
4qklgk1PXVtT95HDrllE8xdRv57BnYUKJIw9XEt8Z9gL25W0oCZR23vA8RgeqZJo
DRrV0YfOFuCmYU3DYSz8gUTlknFrx70IDf1gBtDQUA9JTw3R8gKVr8gnfBjDUtG2
eKqnxZj9sHPlGW3shWp3+kzW54hgyboN1xtZA/0B7eKZhsd8vsA7EFUCKOhbfHXq
nKYKMMx2/zrPWXKQ4lbCSTcdnF8our2i8xOmF0vC1XEuhZ3H4nTIRm1WAiI95T+k
E1y0593hmvt4Nh4zOf0sZyIWvFeDQnOiBrmEvnMhO3Lrtq7ZBXh0uZeZzj5msZ1R
V5jlGmDYW/nMJqDUhliS624EpDm+xlExUGEaHzi1IUI3OD9aOHp46LqJFcHf5ZuA
46VzAE8vZEscc6wz8gOxLyTjvNyvrDl3rspHE8esuRKAFWVTLon6rgC97jEx9wk4
MpqnV122lIZZjfawMX8ivKuMacXprNFawfnXxfXbBrueca7vHlCZUCfWtE0qcP3Z
Cb8qOfVRetkikoSFX+r76BLAOnF169uUIrstmscmS4wuoJfX5jdnPvxZayS2hWbk
Pk2UJ+j/dwBmJBAb2FA1BD/F/0whdr/V+T7KDTDPQg8+cJ+M2+76nhHW9GP6w3Z+
f13sF04Ba7FZHjMCIAr+B1TRzHcTxTvXh4KUh/7zdyvLYqCfQwSypG7Wpmaotobo
+36Sulgr7n+QPQcUDleTxoztszs+ODn4HKf+S7LTYPaioJb1xZR0PVnWfiwvKg70
0n6DzGyvnslxTZZWAZu0r6cIvhyafvkF4NLfUdOjY2JLQ5S8WX+FvIw5TjrIRFUC
OlMG8cn3wf7rba11kCZfl0gW3D0MnKU0weqWnEQwVGUYUHSDZGAC2J522fHkJ71d
x/e6tP/xZa4QId6+ZdJg0nNYHgNDY6g9CgwGybtf259wVHZLwDQxlBE5Z0tw+yF2
f7ILd68TKXyZ8IM/nsZbvPZZDWq9iEtIVmtMm5LzgPQty/QYZIqdAV4PIVCJXRJf
DReuBpnsuO3o/UUh1rqfuo7sLRNTbbArIoLMPZyuvYbTrSfetkYk+7j1ZJXekJJH
saXaWuOptuvSisljcyks+IyPjhCGO5WgGZpKdo6N98J+s/v7n3aJXX5cNjDKP5W/
8cPa0o1+aXnZZNsmAFufylGBxzWxlRueX5PiX2CAnqBOGK+Y5QWcMRgBYTVNq53R
+VWSkGVQCYBOY93vpA1yDu2qF23TdUMDUcziR3JlhTlvdBJKdZVNxiRrKifIOY9Y
2Fdw/28G0rgHmpJyVr8e/Ta6CdgngeKQpqXoPATsfZZsLmuimnBMOZVQSzoEipnH
/nrWhybxvsh1rKbLqohMRy3rsOteSR8JO9dQuI4by8AazGAS5isEfTdkMKMKYRax
Yiaf6cAnwUeDsyP4ecKFFDIgn/8a3USsOnJYECwLizs0IP2Jg3xhCvCpB9YuZD/l
adcfatojHRSSnO/6uHz8mOmYP2nbgKcKFkANHLKMbsM5V+xJ/qp86WLCH5M4syr7
BT4DekmmuXqllWULtgzXR4aCzf5zp41hujVWe3fQKckxZArWElECt4xinX7F4h27
aml4giowrGLKD3imzi72gRRpgtuYyR9F4djtDjt8D4f5Pw2WW35fThlhCV1VyLgc
KP/6EIaCwgu4hlnq8KyIuP1wzf+eosV8K15P3HlfV2nkeQPszakEyE9ReGiMl17Q
t/fF2XB6hEmd8/IvsurxfA0rXUXndQiVY/qo53xxCzRSLjBF9duWMEMKoiVwmMf4
8m+iZ0MjmFm137kkNn2m2hs+CFbc2SEtJd9aJFPOd/JveT4ZwCrN/4eptUCdgWDV
8kPIfZKjUJjgqxICmqAD+D74/QomRVfAMT1aAKT/QzspXoVWvgS5ZBBBvPbeRO+P
/r9s9iOJ8HtNhP8jtvn+khOadOXIC7MxktxSgduOVrvxdSYTFsfEWpEtTcR1aunO
4k3Sswat1MVDSbnddX1eFuFVmDkydAK0/hTuEEA+BBKo4ENvxfc4dsFa5N3wiXQ1
WPeEIdA+kBMEpEdh6z4hCdpatY2nZkRxVFd2iqYeH47GOBQhNjHYogk1r67HK1Ik
OqT674QJBPulyVmxIdHGsbcQ27rx9MH+MvTc9KHGGiGJ80Jg0n5e5Vpy4snoHzeg
Ip5muk1vqaQQDwKgg87NxXxp2sJXAkzoRJWu+p/Ht/0L/DnzpW1kqZoflUXBqhgJ
dRMJQAKP3MUynKK1QbcMyhZ2amPEMlEo1Y0sUk3KW3ZeRXrxeaYxCxNfHRmdB2dq
KM+uDE9zULFeEi9xMXfDdSxKPNqJ1oQLI21IGDbyJAWDZbv2hTGIDsHULBMLIYnY
B8EI29Sz7qJXt9AiDmOU2IkzI2ZX2Bznq+iZphjODTwbucWxZed6faA8/OJwgDxM
1uUNx0FVbRah33S+caMY/1V5IiZTJ3Do8hFKA4zy3dGKaZEWDY1YRv4qMaewrdjb
zmeFE16+7sIFxRq6WO55b8p9cuUGQiOe4nj8nvePMSYXEhx1A9yacSNfQUeBmm/h
kN1/5tCnTxMlIzsEdTb1ERVbMjt55RU1rdwaHRWyE6QIR5yEwqSrSznBkZnKLS8e
JsBCXk5MAAZ5o/l8icF/E4ixTvZNBlFuITejZoKJf3pl2OxjrX7E2MDhA5plky3+
nJVvOZnMLh/uuc6vmJ2BRcncj84hF1OHwzK/Y66fQUPvriCcXBi/iCymzKl6LKbr
SsKDqL+VROvMPmkLTvMbaxCHzIMWSiejjrK7O781HDHlYawAHBkPK5I+3CEbe/W3
lK7xFtVQm47s1dsyoJaUcewlfpAJ0Cgi1byYsaeKRsieNrHEWZUP63ifnml06gVs
txU149xk6yyjeGewM0slVgzO7T2XlW45Vqz8JfrMUsEfGRxr6L0tyYt5bKtcTQu4
oDBs4gU85vgydz33YjqjsDJuL7mzMu3GHDVKKUmACORhIPKWyxv7t7SrrlG4vS3F
btRR43PWLH+zWyJ8pfkcFJg2JFDc2PuclhGukyOGpnPk7BAUj67icBoUkFdBuKTq
K/pqeuhcxdyVzz1wSJhnMmvXbdODibw2hatLQ9RNT0NbvcQ53ZnIp6Tz4nisJUJl
r0LvCFpin9e/3MWROScBM+5H4v9R5MpLH37DlQWVCNQRkWKy3vOlJo5EYWE/HFOf
Y0ol6N/OYhUcAbLInvdyAytMoRbWyzDvNEdT8RcYSgGhSHzS9HwcAQqebw0elEfY
yFAkWwX3940S0XMLMhTVI6BS1lelSJu/kjZ6YxfXgdJeRDNGONjbMVfIOMCgEzVB
zSYAwEdxnEtZ4Io2SJC0aH63h2dl1rki/idJy58qhKG6f0MCaFpCcnwxTu3MVLiL
qjRg0nYl6gWIHh568HIqAklfY/cDJdhLSk9gMJ9OkA8EJRPlsjLQflllXEfIV1xW
BW6YtcezgZrJ4jsZvNjR7X3Q2IXi0UlHU0eNXrKw+073WzO3srnKNToUbieDrtcb
YRt8e9COZ/MmnqRhOPMw57PWNGEvhrAhyhKbIk5KgBSEQJ7ku1xap1wrYP/jN0vf
yJ0ljAEywjYJgHifwQ8qr/wFMilQhX47KnYdAFD1ErXuDKR+DTMFMGL1MXLf9Wfa
UMcnejXcTrtOdSRjMigVItNQ6G5QjUfTcsKMZeYuasG3ABIb6SshKptP7jS+rQlL
I4s4QNEEt6el50EbYXBY0jCog5uX5NcPKk9lo70HQFj+SNr4WvEZV+UbGYf6d/f+
HL+YkHCqftkdNTlux91YlUIKdu56KvroG6oJ5YuXhV3y74OSFferzITqk3iKaLBD
DmoAJDg49Gh1cQbek+4y5w7ebb/Na1y+y8/LCS3fUdmo5jmPWOphh+7rCuL4MzYE
BOHcq2H9PVHqo09K0PuNKY+U1xoWsOiugnDitZNaxEQv9rpo9cjOcChbPgtEPraE
n7NweFc2lwfdIZbRUOlhiVYraXyZYUIGOI5rbjSEjn0xjBzp8irCyvYzuVjj+vwZ
l3xWqvfT1LSDCF+Q9PO3DDq72gB4Z2BBZ98UPYFDafO/+hlJQ7JjMfagxaIfHJKm
NVN3niczfCIAHSMVe/YuniYle0JW+kfAhTiwwF4oNCP9eiUXEHZRfOUT/T0Lzn0f
cFMcLelCP1rtolAzolIGzygToMMMyyU0qVru76CPgtw5aQHGdPMlyFAITlmfdcY5
+lN1UCsnPfpzFnM09kji77ndZWSATl+crsEY4eGkeWePYt/0KCIjxXl9+2vG14sB
9OswVFeyK6JviZ2BKLqJF7yQJXFppowcZugaUu/1kawrpV1foD+nrNiYCKjTJ2aR
BoH23C85GCgyaNq4MDwW96Oy5ys2AfuMy7Fp3RW0Xupoy8TEXdJIuL0ZQuBZgM/t
2JFY9YsdrO3EwyXN5ITORVLDSfRK9I3QKZaOfVGUuHKn7OskJawDXCi6PVM3ZJNT
F9+k4Mus/D0QvUAYoMDzFgx9BUKH2nkM1CJJ0zdZdCYDTc1P1jcdg6btX9T5ZSkO
l1AhYENI48cRUlyk2g3Ur1APqkG+TbYEAIqukC+mRbRy1bYOlUekqDMOiDmXg8id
x3ECQVBmh1Eo6GakZBRbTd0EdjGECJcCo71XHwkuNUjODkgwYceSwQq+prrqKEl6
YSqjzxjBSBxUlka16Bw/BPLriG1E55akk62eBWREDivqMiVb3VlHgIiqXfP0gUga
TqumlEnqzJjpiYZZ/QzNIMY0Fm2aTpnzSoduKwk6NMBrcGCqTBkm8kkws9bU60lS
/zNBjJR4dew7+JrFYvwljJ9yp8j3mZ+427arkP2CNblqECxvuDzFkV/IJfSuBjfw
V64iEr2qYH/6bP/IT+PCgu4SVbhCiQOX5Q7Id1jzrkzeSjB4+DXQ3fckp927QK+z
OGPydNR93lf+lTw/9Lc70lUXojaCxq7UKA7Mm02zactCDBacVGMgK0z2bdzgNM5d
F1mTYQTGKlwGw8BE9echbm8AabUPev6keTbXn8HrMKCr3CDF+Tn4N9OS1AY2oedg
TmSMqad+An3Qduwpp8907GHsYv4DZr6sC4o1Qb01bn28aW/a+qjPTPT1z5QC/1wX
oAv4nclhX05dGgf/R6CZzSJJS88vOHdUcDfodrjVoclOT8HJjQrP2xrsg3omUI5w
npXbuEMPn7IzoDotdQ8I4SieZwaHzf1OfT9BBWrOJ/fYBir+pEAGKxojuwpXEHlR
cr2dgSlVs3+nXyOhfE5KzQR5ZqxuNRwiCnM7NOWXzhZg+Y5z4dLzTaPsyHu7C8yS
wKMFLW/+jcVPqaflkclDV0zkkrucv3PCO/ut+eopWocapvvUg0Ms5c/yBUPQvTL4
esjFDZctbBWHnd4J++xEO4xFzI72CIlUS/9ZZqXwUoiPDrAK5UtCkIPpAgPyG9Eu
QgLFoxwn3LF8mz1DVpNIzgFYJ/0oYXRaDXV+tshMAyGgB69E7jIn8FmdDerukSY3
+1CPqEY/iHS276A0BLlUaxolYAU1i2lvG2vfi2wbmm4WMaHErTUObSZiNk1fUm/W
rFFvSseN2IDexj9azIaYxfpqVbVgr6QO0xEeaRO5ZpqbVoHWz0lx9Zia1Uv+et/0
Dt67zlC9iVmHGjSH8Q1lXSnF/D+L9w8GBUeeNczd9bwZc8IbYWAXqHu23ODGTuwa
YMF4DSxNeV+ryk2wQOxud8ZyVtaS7Sev+a1gVdTiuRnYjU/T0Kj1qBbaZGZ3CG97
aLRWPNEbb3zYbY+BgksJErfKzNFCjpszT81M+XVOvT0KokfryYZfCGurkIPcoW6C
OpqwrqOv78dXEFXYqdHRDQIZJCncCOGMDfgZDxQS0Jr+Ud9lNFCbCBMHaTz2DyZu
usZZkee5WnDDPOaAWd+/0TevnXHd6ES/Rg/kwe+Zf5gy98Uw0Kc7djM1VghWsP0a
6z8qlecyy559H96t8efQFZg7FN0WOZ6JsTt2enj8wTwYRL6l8ipH9L2zLoRDEEiF
9M5o93juyJ7j0OFUAjI5W1chlaYViUkguw8I0fGIUWWRwSG2GlDQPmaJrdM+fmBa
2Ps8chw9SLIBRh6RgbgnRIPm+wfbZ2rVXBGi9QUCuy4VvJJ+5RIW9+/AMkAvp2Ax
nSes3wKnYepX1BknBNznjvMb1c7aUcoXrnWLtmyLbd9iwLYc3ThjgetKY3QFx4S2
+dWcCV58rjzNcgk9OkHYfiXxvX9sBTDEns3e2CmrLGJU52z5QsGXsx1G8J+sPzAZ
X76rpzxyTGGzFcjTlACnTVYX9DxpM1F0+BnSPzh69kgU9gXF+vR799JeAYqothsW
WZX+L9Hjc2RXNxS26OE5G9c+FrIGFlfLD7lJbXPXVsq+5zwbPrAvBGa0SRwFbgND
PM7ZoJR6YFM8W0U9TK17HyFcHaWr9oEbJl+OPax6HwZCTRi0DPcGk19jdjsTxWux
IvTyXj9vmoDJRBlCYlhqgks0xPpfjXHJKnhElm7A1TuOC4nwcx2YOzI0yS/LAhJn
sQQeHu8Zd2hhPN54YAAdh1LZ5GhyjH5Y1wKo/R+5GMPVb9ExlQsnKDezlb1iHBpf
kliczG6A9CHxrRzxsigDKIjlHi+9dPhNDR4Ar+KkcFp6ugbnSvjcX8EhII23F0Vo
G3K+ureRWCk5GIwmNKcuhOs8mJdeKKq2yPERoM5jeuTyTmTkIbfn1tCw4IZWMD9w
rUM1h0q3+TAWxttRMwFiXfwPM9j2drlolGtFkaC9UPEyWpQahZIrdZ0QVXTPoDxA
f3+1P1GvOy1ri1eidf5fPhApGX/0pAOju7S308KNnKGM6qEQJB76eGl40uNHMVOf
HuLGCeqEx2LIHlQ77o6XfVI7aQn8mWbLTFigjId4otfPJDYLS5YENVd1JxCXWxTM
OZMODVfvWqHCbVXRBHQ2kuv6Yi8BoJ2j7SFNvGfDg2iZ0h0ZfcR0nqmU6ba6kn56
oRaIeZktIcq6rcgk4S6hVZHKkNKFgxXsF/EmYUWJnkD5TYuydImbTortFVVQqWCu
m3vmofUu1heaLMWO/6c/2r4SAMpRNSyICT382laYYBo4ZLOtCNRbhGEIpMQjd4aE
m4SoNPRoYE8UNDTIDMY8byJBlb9FDptJaBErEVPuH7cqCvcuYt3vatUZspK9r+5O
QSHTaffmFEfSkD7XcTT1GJxy8zAZ/O7xHkFTJQFHRzOzB31lUI+/q2PLtalVNZtI
xxVI+AfStbpa+l61Peh8W+qByNPgNsfRgfZrkpgcenLVxbOKQAoS6rJGLmHWR9e5
CTLP7wCA0q8GjG0uAKYth+K3vCswQQUUTB3fICh8V8D1NtUyh2zBCTXd0+8Dnq82
BSRhAC0Y1p1MhewF+RDdt2AeZCmzPT8C1XowwyfHLdXUdYUzuDdX0C4lXf98ZHjs
4D9QCinNoS0pghy67hJDb5p4U5amA7r3wmz1OMS0Qj4ouzQxFftEElqaMGOIcG68
wwkc30+6Bzig69w/jrpMr6g+2brt3fLdspBng6OsoZyADGSlmkiOjBfNCDFFEjWx
ppxA1XLYxQn9WmFQjtwSSB9tedpVzOq2Tfm2VL/NlIyFKvfJJkr3m+rDH3PsMN7y
DbEg7S50wH5Oc7812JHaGydBmKC3RgLrH5il2u8Q+v+lew8pYZsg1pZtnbBhmvKc
A16ZaHvXldtKCYYCz37Fy+K4NiUnyRY8AQhxer6XNSOcdMqQUO1xjn0QjIhZUVmA
KvADJtcQUTAAbw+gDhL4N4uvgSj4AlwIIevq36wKjrWoPbt3AKAO+eHBVaGoHBiF
TUZ/1AllEztlntFC6FXnXeEImMLCEWd7BKb6IQN5bWd+KaznTD0QOiwsC5Vuk1HB
gL5y3yBK8wG0rl6GHNpH1BVtJJdwcDuqpgK9mhUw1dbmFOg9U1Dp2bE8WmBTLd+X
xeLD/BUJ0L7gMStfrUAePlSKGN74DV8WzMf8ZsvgkjJdnlYaMkEFGWzDsoL3HiBM
Ab59g8IXx+4PzUPSS+SEXG9hosbMYRNaxB4ADEyE9ykRfW5i4At5R3CGB7Zj1nXi
YzwSKKnJHtVf5sakwL+bSnc2cLOKOYt5SabrjH6F1DY+piVPD+2hjgZ0NJETExEr
2JhPCVTaGdOMjL5VP1JoUQUSnWGcov375XUie0Lhvv46FI8HqtKdGoyTjib94PT9
5e3CYpJT5giRnsrXziy5W8KK3BmNjr4YzOt25kkB0UtrenNWCyxbGzePp2Hwhp5N
ChLUhEh2I4lyb6hEtTpaIODij9Yns921sdyovkkH9OdjgKq91yoAOB0yM5MtlRGB
2SXKnarxsIllpNEIuZWc6QM5zY/qLJucttfYh1gtgmf8E9e4FlGrkis28vhafOVG
Bp779R5WBcaLUUcRT4JTs/lpPPvmHQaYXOeBTDkj7pEx7SlGDDyIZhzqawihjoel
P5K/RTAwvJouA9OwGKKGmQwAQfjnICJltsYdElBOHR81ugyTy5wUqy7Z/jeh5iMJ
7A+WpIgca2E6IpNYMPm29l/PwIZDOxQK/Nb4606qpFRtf4xZJcLBiHOw4tsWNfhB
4+ESi0zfE1T112e/cU5+vQe/7YuwPjNAmL1pSZl0RAuRXVf+SZHQFFbkn4DkjdUA
tYG/d4OORz9KTI45JlVTmEifRoyv/rY6zAmLNM5yUAuhQsYVMx8yjNVgtBfLbTzU
ncHKMB+alnPo4Rg6YLpwUu1Pf+t3YXsqoWYLqOIvwBXBrAUF1JR1b0ijm5GfWLR2
AVY08OEexf4y3yW3jmurUMzBsE3OUvUroAeneOj2d/iA8jYamnxNwU3GzMvIsMVr
TsIRvqdNP2UPX1FnPvA01KzMCVj/rLNfnlzB8i6/rYjs1r0MoJqf75Pl4eKrsW+r
dnV83dDQrH8yt+7jE2lJnKpKRh+u4XTVtek4h/dvsOCOdQiuMHr5n0myHNkfCB4P
R80cW/HKqg8KsT5e4Go3vQKicWAnhnTv+nRi7JhKYOXEUOAGLApBmFnsSA8EXx12
DOEbTAl3DSmVDigZdiEWf2faE8naiF7bZOXKPPP6JGZv5WfiyS08s933u/o9yo2N
2Jn/cOo3oW/VYN5iMZ3bTo/Yz8sSf/yqZoSGR3/H2nfIuqPUmq+zxjRHMi6wFLfj
S6ngpGp35GgVh7+ukVPnHyzs6k6QAY+w6CnmwPLdC42vVLbBjiMcsZj6B5WJZLmU
BSB0g0Q0kN5cBgwI8uTzk7gEVAwfS3i7JSOEbxB83nTTMkXSXxh/yG/RnK6m/J+b
u5I1uAp9XHav6+FzEo0bUt4O8jxi/3irrzWq29F5v6h7qiyS9lKHfPsatyulO6rH
w13VA+TRQTb/H8DmyHUpAyY2WkVWt+kACKydVbHGcWYHPhDlFJeWWs/pYPb0e/7g
lRVyV+yCpFzz/8oU43Ou41K0gH01HmJcV2XeXb2nx8mgfRF06CtLBoK1TdOSkzma
oQA0JGLb7orZg/ihOWxEvCz32N8+zmSCjIxlHOJmhNyrH3luDSO5+jnCtbsZ8Hxy
5t9w+Csg2ygMXyWXM0eaNRc8VHhm55Z3YGN0yZwppFRiotriZqx1l3rRBYQAyJRB
VmFJBKUov5UbQF1r/rZWZWaRpK2MHooqEFyX+TbARYD8lEVTcAbdKHQwdVxOckpV
/0/kDQ1mnczrbUUk7WhhRTv/tWZcgwAEein/qvUoWXyUt1FRpxb7f9qM/Bg5QbYx
W91kLrWG/lr9BQgZBprec1rdLyqKcXis7pjEsA1aADAeR0pbykUihvAaPAA/NNrj
wusfAkvz+bZ53Lqn/n50Pb2xW8HA9C0BkjgFr/JaWfHZwx9rbn4sa4G32muX8kVh
MgvhBStb/Qm/ipmMW/P0fFRJwNT4SQAilps9oAFTTv1m61ZE7auThBdIu3e+6yZK
Xar+GDq9vYL2TL8pZRO+QLNijdIhOUopZWJruH5qHPtRyRY5Z8Yo0jWSo6TRFgSd
cE2ZdqiMgSZf5c9G442s3bqQjRwOMLzlMqaBhF2vlSpTHEGZT61GZWWymizU21lj
hulnVZqzXAOJW67bFOi5fBghUMrdacL0cKoBcfMkdO1WLnfXOLakl1bW6SaO0jy2
a3/m4z0zmFqDWE8tWlIbsvuOVN8gXmoWxNNt5dYZe6DfxMEKN7dFm8NcA9ivgi8Y
+8P62//0jR/+QwYk4ZKzDimGpvLZDuERh9VwFLgG9nSixYBzuwOOs6kz1ALMFFMS
PXsvgkDfI9utAX08GaHhFvvIUb6alh2KFs3N18boeb0cbnDmw1V3LW3d2UklM31M
beLwF+J3njtf0zf5CLgNorVVP72cBOSGBHomIrGYvb8mL1BYhhrCKJmMMPx5W8Pw
2Haw77B5SDj0x5TJ8KdDKv+EuzuBxQNKSPKfz08blcf0z245lKX8KVoFV7UUKkIp
VuKpMThhMMik16PRwBptm1F7hrd8PyCqmiF9jnD7iedhpqzBVmMyECcw5V7CWz0K
habUZeU8e+6D8StzBKrkSbdsZ4MsRHVULA15q0BOIXsYiQGrgPQBrCRyfRS3WQyB
BYG97Duc560dQwEp7o1LFoF9P8Y1tqB0qBDNjS0Dj0cnBgx3x71Xp52WAJRG80cU
XH8mEPf/eQaT4o1x9ifVR3WUsorq9VlDTCJbAolpIKADUDoYkwPkax2hWfSdc+FH
e9gMmrg6uvj2VPe5XVJFLrQslNdRVVpZydY3N+VvWaFb/73JohL2t49OWP5pzE/N
fFN5QjgPe36cn2jdATaX0XzByzziVg4bextTGA+qjOWUq05vJ9ZJfSts+opkRXbj
EbQ9e6YdM9JqCpDrJD6XP9hjUNqv7Tp6E9y93u6R008NDtaCVxtl8Xn0NZg+E70m
5tj2LKhJG7H3im/sJQ+TE16HElURJNF+vfbppXwCQ6OjjwG+M++xrbUsRvdNZOYB
CEY2rTTyrPMPiiE6KnKshAB/bDTqiZ7RI/YT39KRejhkopWY7BjOhtWBpUVyswbI
bsrv8+AlnbV8rpVLfMgd8FuYjETkE30Yow4zB49girQgQaaTkQg80BnFMR8hE88z
DuKeACElfMjeYtfmhU26AFp+XitJk5wlKxwzYMNT5+ghLyaZjkSYl5myGezlAWYD
uvBXyXtmpqedn8smYwULyIMUQ469ym4VJi9ngHo/Nedu9Oqj4074gogmRe5xjjst
7xKdwW/Ikdd0Q5rG73mT3qkbUHAdtj4DFVYDs0AE7rJeqHmyywfgGWz7Bkkk1NUP
6qKa7WW9etvWQSG7OgfoLWTe/FzauS6Nfl5gNV6akwbagwnX5pThbc0m7KlkOaJu
DDxqBOavLlgELVO4lfsf0hrJ/erbPF52w1cxuHZsc3j4ms0bXM1prwPq5iCqW30A
+FHGqpQ6hEYJJEvZh1IhEFKACOZRtKAHueAMHn28wFX/tGedSECUdoo+Mty1W0MS
nqzdk+VPygg8CVlpB3dAG9Phpfr49NonA+Fzqbn4hPZ6L+b2Ygh5SXWo9fJRGwqL
3mSqLdS/TqqDBJ7WasYb1SKOSbGNdenpG9WwFDOJwb1yDBrLcw8Ivqg5QVSqwFWO
McSisFGp/yGO0DWdnayu7vMBh35Kh3O9QKQpAitacgBb8X3b6zkaac/ZrHk6aRxc
vRRY2uz2XkHmh+IshQzyh5KeGUVviv9gHJ1yHG2VtseWenqUs650D4VTJ8kVidV/
pl6pxsjKIRvkQDOVPUYROXrQ+szwqdPHe6kWhrWGmzt3r8hSvivZkQsY1DVvHwX7
KnL0vZZHMxsusL/+8hjeTTO3USj8J/aAwsxn5Z6YUPTmKAuties+pKhMfpMBP+Kn
EXaKoNEmjpuvdER73tJK5jT7vwKEev+regC9SSxL4iRugTyjE8coNmZdrMK6imuE
8FE7EqDedgu68dYXwitjCK1N0kLhym9vBO1gxXTSLGl+2dKyplJngX5m0vOZs1sv
MU0kZbEIo5yj3c5+PgNe2w7wnvba3Xtbv9SCUu5F0q/gtypgML+az3DqH1K4ixDs
GFkhsGMGjlKg06aIrcOU+UIpLGtVxC8X7sZdQLOESH4mxly6Z9SPJDyyVhuzGdJe
NdCgMvQoInxD2DL2BtnAzGM0k3ElW5V/4ZPHoyn13xqD/Sd9wnGrqcEbI5mMkNEL
yEYFXhO9JLcB/bEHOC4dLR4CKXI9fx51T/xi6vBUK2u7JOFQsvSILEvEkjHmsrp7
r6EN7ODDL+88A5tQLJya5vsc6xuYMItb+UWKJ03YW9KHfB2IyUO2LiNzcSwo6E1j
evdYTqMLyGKcxHU025ol9Z9ZJLUKy+1MTyQtSydLxnIwusFnqOqaWPShgrkumNfm
J1XzzGRTdst7Sb1HL6jtRlo2GEFzQp6UVo53gh/gxWk13UO7wR9iRYX7V/8PuNGm
I9RU0zpsbH3Af8DiLyOrWZ+SQDYfeWOlsuIuEByOIXKwLNLsq48mKZeb0qeDNWbc
pmDFafEmf5yVMIECxslwx32cAuj/w6V1PXG9ryd+PnXJEqXU8/W6//5QluRg4BVg
8Gh5lDspdntIAjLrUPdUg4iCq5H+8xjvQUZKJJpZeDQ5z0SbXiTS3azhRgOa/0w2
wO/VihL1y0ErgFpSr4HuXaSq+oUURPvE2b+n2hPyA7y+/lDXNGEvqcHnneXfQh8d
dXybfyIGIFC5DBvUSNOK+1/BpQq04JRtVKLPtLonE4JK8KrOQ+GbIRiZl9wCTwsL
9dCjnc2tZH0UWnsQrR59kSsEXF0jb2e+yLVlAuaTmjbSwUKEL7GPXdNi+YQHSOTh
5Oz8JFrLH/93n2KqQ28vB3qaMuZu1uBtgGWn/QU1pUuZo9ppe7b4byY2YDsmdJIu
N/tJXcx2iL8NOVpBhgl8r6KE08ZNQJbmkVaq9yz27z6HcL38Y8pPP506fZc2EZOI
zQzMkkk04kNU1v8tC8PEUbjj1tdsTog7NAYRy6S02+N9MND+fdlcIsJxD1XFe8UR
cTXf8ZFn4ygB4+c+oDldZSiqCrzYkC6Z3es3ahSj6GjYIs6mkY7Wr1t8MJu4s7Sk
x30+hYgtOll8eYQ3Aju+gWvTHo9g96weE+bcHMmjpeMunOh/LY/OIgXoQFZI86//
zfZamF5N3Ihg8Z7DLnKNdGB9i2y9nktYpgPzpaqY0wNmr9cPMRWEZ4T7pgqKMfQQ
Ptt1vem0xXN97V2VIApIhkFat06sM6hOkUsPSgzZKWfKENVNmkpLVNPTuWZDqnyJ
260LexceFAkvJ/7UvF9MezcbtQUPQO42xWGjlnY6qvssOtXsNCWRMbraufVcM+w5
/Yn98D0Em2QDj25k4Xwxn1wGfKLWL33E0BO0pN3LOupdJa0BjhnKVVOA7dWty4xU
6K9xxCYEDf4b5wywN5hCVehLE/7MaoIXACIfsjrn/S2CD0xJaFsah+nkQ/f1uTdx
tGA2dTiNqLI6ENQmmV9ExYQPMEO5iFjCHTnUQvzdeEr/bAnQ6pM0ClpBrNHdcy7O
VlZoMfucp+T9zT/L1LYYnLpcontDLZ/AR+YHXXG1L98gq3rpcY29WHqomN1aPYwu
9vDZH211QmBTzEiIIzBU6Xe2u25BpRINyTP+EhkU8Z83bQOnIPg8k9FRPxmi6Ror
bdiCRa0KDn95xjg1+bKRLWuy3m8rwv2yGUlC2TzUjmcrdd9Zdh8Xt/B+CSt55IB4
0AkXnGQCUCT+g3puUPCmpb2FjFrtCcLLQqgr7gC5ewjFV4NtW+/QwR8qL3zB3W7V
geY5CHVdbe2knhMdD7qIcZTc1snwxoZ5W5LQzNHxBsyqyNblWb0PedcRyTQsAdAU
FOpyg2Zry5gg8OnZyhsQ0yTbMe85YVVGlsbRJZ6Z9BN3cWoXDS1gYPc+KMSz8l33
GHBwW4fXktBfr3C4oC1dGgeFPVivO02Jblmr6FKtY86QfGAgD1GmY/KTMHjV5Rgm
TxQYFYIfqyaEVZAlPuIKYSQXE263kbaAUP9sIG6gRJbN2icrnW9BuR6//hGgx6Hc
h4tgImIsizmG7S5LbexdHBcdrlmQZuHq+wG+PtnSrsinZ5Nz/UBxdLia1dp2eP+v
x7LVFCck5irLfQb8Wzc5/M7sxmPG7Ma7tI4gzHPk3efFQck0oMeRxDQRTHib38SE
7NnH/6oJloDAsEY4uFMX6JxFL52WxHBHpFhzkuV19dgMEcsfECAYtZIVbEkXj+FJ
DkhhyiYo6fjOlHvV9B4Egi8fNjxzRTmd96pzsYoqZ8YcbJKOQWVA+/YEUz3QwlVa
sfAh6ceWPRPQfam3up00nVcWcrenWumUmxSTFEEqeuCk92kNume+9+sf4idHSC0H
S0BYMJkThH7JE/Db2qBDogg5lfTdfXYxCeqkGZAp1T3AyvUa48JVtAJiXCB7x+Tr
j0lkKd+X4DZP6AVIcYlM/zZUk4xiSu5WgTMnD1gdWkAMtEv3fq+BgnbO1sxWlCRy
6Op44pyGF2Yuq43dpb40BwpTB1w/EhzCtYKEEfnoqgBWdSxDMzgkCRzW0TbtJ5oj
MR90TtVT2HRS3Q/+lkb99GBOSKyQyPCkrP7EO7eopyZC/dKWEP0pK6T3rWchu4XC
/iHJ/UFJd0K72K1SB15h84BiuTfyrzLV+TWTUO8Z1r/wf4qhnJYeio4QNYiJTFtT
1txBEyIX5rFheMOOeAx75bDkm6w3z/TuwQ6BEz04Sd4piWlbXkDwdjYUoHFrOFh7
bJnj38YZgdgMAfRJAbcdieGIJO/gl1FhQapG2gcQB6aJzClpk1LPDdLnnCrleN7l
ZFFvyYBAi+5FgO0URmz2VfA7Wjtyd1zJ+AVUjnYb4Yc5IwZ9J9LXNqMk7SfR/JVx
UE20jvh0vo02hhHQqQkHLTNN28gM/RvFCedQrOGgJfGhCBRz4o+zWHhLNISeTigU
bTEvtdsLy6e3FKn5NG/Xq+36WifyMLdzplkBQX4/IsYPJWlzeEp22yYnq/BfhwHw
2LMGNvD84YB9+SdWd4QjgQ+9mkHE3uTq0jt8isyrEHU0MmlUIpXh+omwWtNUPWRp
FLxh5vC8XgBaUqO459nMmAPImTmTxkHnxZBagREEw/PveEcHmzwpAWSSThYpABF9
zSbkntITep7sNXsuyU/tI8wQsV/W5+Ei6uHBxkhBNb9tCHPQu3F1raM0KMzOXFef
b9qiM2eVo9qkffn88Au4CIm0XKoYWICnaE2GXOVmdayHzF7Q6RsMxBfRYBqSyCZF
Js2Q3k1y3Go3AgNk9h96i6i+pDNpcqCth920rvMklh/mYHQ4PmXgDWmvYEGAmnOm
AXWJpqDKX1pKDUC9+093I5b0rssNkbfuh0jd84jRZ6jRxsTkgaXk4+Tr6y2o1CFv
55OU8UNy4Um0HKYmGEv0AyZYuxEfZSzS7pi9QZfot93mt4BIaEj7xiLcL/rAmK0b
/x5Jyfb6wcDSC4thCA55k5u/BO5sNURvWt0MFOqehoN6QIVL0cP3zZo3LNmOAB2A
mgjNOfvBfc2LdXe/c2yYLdt8qv2RW7pGEjlwSHw9RfGgqQxJMnmXwdF+VXVkREgj
yYt3OQjA6aXWk3J9f14CavEftcQvRepft6cqvSrufriU1VmXjyw4MxU8Hiu2s9fy
LYjoURCE+fRG1PjVXryRCUnlzg2HbguY2aPdfnTT3gqCA1f+KGq+VQeNCJQdg4TG
p8q4DRp90dh4aeqWp7RTrPtYfxgQld2S51nws0n6kb8TvsEzfXjQQkVGYNDb0tkg
W2ToCVZhUCuRrf6sCx+iSJqd1rDq1mMtu+szz+ueYHAeJfgkvMKhehgzKAtxvYA3
8d/5j0JPkHHI6IE9GbH0Fz9IXQz4m6g8w1seZC/metu8+HsY8rBHbZqeDGZWgMo2
E217PsV0VnjYq3Oh851XrLKcCjlyiyVMCzI4vllWK5Axodabk3QNvxoqOxVZGz5w
3BelWLftkWXcE4GVR7PlbY9wNgh6a5PFJq+x6d+0Z5wvLw+HwQOU8Xg8mtyBWEaK
B7mmImYuiInYonPI1ix35K0ka8j0M36CIO7U8bcZ5h+wZwLC830FXsK4b++zJEAR
PVNqzvImuaAt8ggTAmJy3hu+BpVzl067XmWHK8v5cZTgM2VTo1yzRFWhJ8/HYzug
3lBc30c2h/p9xIjt8lS2q36Z8qVU+1VkcmarjL7LIXxGFkqvZw+qhBYl5o1WiRhG
egZ9UCDJxqlYgNI38W07+cmDD+/r+RDSEeCEJG2tGXdxWtPIiAWZBKgF/pA3V4ew
t5VpB/UzycaZQSzrMLjPCdxmpmwSIp2TXC/3wH79Kr0d98rhCck/8GEiMUK9qYUI
fKUdpvwMnM8BZAUe/ckdaE1w5AfXWdpa2cB/VyEAehlxr9btr/yeQ+SGkeyfvGA5
L3rnOHCQUkQJ38yeEWwc2JmaXzofSLxHcPjXiggB0GroKevS8NYBd3olwUDggZK4
cO/p5yMQxJwrHBa5a1aQXIWmKxx3eyHHOHLwKrC5YHI4ZYjgcD8cvPOKbluyFgPv
ei27TzcmkRs9cSM25Hcla8FHhBIgJGZWMBbhhJ81RbqH/s3oWjNvwIsVchj/h/iT
x4Ht13+mRCdWk9SB3XPsSLT/KFXPdVkvx6YdctpdPgoyYBKD1mU5YI9m385MJnnX
71UgCMcJlXFJk7cXE4JUAtIEmYUsrGTT+wFpxyx47ubSYxF2586qIHu36m2Pt+0N
Y0vv5pmvJoIaQFy9pXM0a+hivwjxjCmfaW4oS15TQAI3rcHMCKGVKoWAOT8ZparA
iMcAcR0n6C/9VfT2scsVknOYsSpuv3ULVAwtgjwhT2lJAZf2SHYGgBfL5YvXTav/
A5p7H49hhEmUcSAt4z3ud24HEhB0v8VOiLtCK2qcWPfcFfkgmzrDTWJTdmB+MxMd
tg8QAXdC91jTq+cbw38JTIcQz/iGqTlPLN5WLle82mhG+FVDqvZ5SyA9sH2CDA5V
4nhKRPSpLOM6fBDGI54MNFkuBCITnA2JEnk6wEtpyGN8Ygm/Vsb+0e/Jkf3AVztq
lBuDmNgp+nWpXTn62f0z9+Bxo+LKr1DuKgPix0vd7wnqud6y2Mysvp9E/MmEx7FW
gtdYO2d95wmSJKVDTfoziELoOcQqI3rEZ5owbrAeYT08k297QrmPjvpVbjaS+20x
ED74fPizX5gKN9Z2l2+u7lfCIbvhHE7Aj+C4RP2ubEdGFlVeFqhsviAYQ9ZW89Og
DtbydkoCFHrztracLZljOBl/CGo6hpb8Fxc+Oed8rLEHb09Wwz4BZ4rSO5UIdXve
qlYbghyOEZ3RM2QabKk5ix2b2iH1J4j2x658cIYCnoWaoSe/hqAXCsa6eiKxEN8c
FOWtyCktWLxbr8wORsvA1hf2djlH3CVceLy3Qt/YF6BLwwAtdNaZHyxYe5HYyOb9
J1gSfR/2iS/ErOQVc9yB9x0imtXRmOoUY2TdbPHXUuhsDLul8f9OGnTi6LnqSna8
E8ZfUoOd8zwRb85H57t9dKVd+4zgDFVdfglciW63Ml99SZbnW9o3a7TyLB6sJB9b
WIsBsDlfupAXf6VZ4G1Ug7j24TeWr7nkfzG/fueahaSGs5uW1QnLj2xI8b7BCCRG
dYwZGlMmZX4uk+JkFzy/egaV0F0oFiOJaINOaitqghUONRSpsJ5RWrnJTHCrcFEC
xsoggGwzMk42/8sEVx47EPhwcOkln45tnx8aCcsOY6XKlFusGEULObodNI1RHLx1
DTH3xMyMMl8DBQH17GIRP8XphV5ZnSZQzBoX8yzzxBJI266nbVoPZmY1Wlt+bWnC
PFowhp1QAbAcEJMAmbkgenDn0FXsqRjD6D4txq1muxYn2hiKfFNCg4jYfDK4vWFU
bikVc2HMIlL6kN0jS8fS+dAPgCAtTf6cY57CPr1EcsCMzxEpmqPN7JwNvTR+FXpb
sihU0mLFa8Idi1yg3SkO8eAQGBIWJAO8y0Ekh2nTKmQXTmOMnmwS6ij2GWwXmUus
zQWIGdAFDxo1ZzJuebVdnsNZDcVEO/vO7OPAcBDiDWpe0+7x2+SA+Ik5Rekdiovo
C7l7P8O7DMcw4ahg7vK1DxzIK//inglYwyHJbVkfptj+rCzBvW9/h4IdfrKnUEmF
tvdRBPAGzc9QiciHVOTEwf7LHlBufFLymkdzOTItgfCyvSZFtAEBgsnXNAFBlogQ
q4d0hz3tSlZeIpJfkCwq5W8nNuncE6RzPUnWmGJqbkJbgS1PSAFioYsTaihLIQhV
adfFflFHru5V2y4Ti0Yz7ct4Cj0PrMGsBIEltfTl5vTVd5uP6lfU/+7RkzvcOeew
bSME3kWbUeKdaI9DQBRo0PFWyCQB0HKKAzzeyqaA3WxnTzFVCIK2RvbuLasshMjh
nV4Nw7Y32tkubn8aSbgVis6J/KiZ+mZdpWDU6vTFZB4VvSPxCkN1x0zGt33vVKch
u4yOs1KWl4C4DTxsY4Jdjrv1LWa6o2RRO3j8gjVk1rzXLt7RyW1ewKRg/taT9jjk
F9vPqs+hrAkVE3Mww7lMdDpg8revkQO/+OXuuflCC/SCFc6xmADyHqLqNNYINMwI
CgDbumut3k6LT4YgoCjeu7A7gE6+W/u1Ki3+37IGNZKHKh9rYeW2qwmxDElvLVGH
GfphSGZ2Nhet6p6K14VpDq8yY9/aqP59ngdr2qGRAeVt1EV3GgknSygI5vSauIOw
bGGHNTe9q6BHgDFFObvvkEwLBjBIvsPI1YWZYmU8LUS7nTsoZsOpCA11cOb9W6gA
zTRUokyhW9kDLboAId77vU5tYWz72OVYB+EApgY4yBABbN6jccIEmHVxl2FGxlio
vZwXGvpjE8ORbuSRvBh6/BGrEZ4f46PGvGC43N2ys8pBDg/SZVvULS6bm7gEQeNB
yhzWFQUU4ZvQ/rEYAATdAc6dNNIaCLc4iLy7KdJE/wQfO5lRZc95XkUJDCFtij7o
k+DR0oTuKEu9go/zebAs/PytLNUOLeVu0/1rzT3EiFEKoFeHH89sGjyv3Hv8r2cG
MR4bDVj2AV5ndmpCihEhETpTX52dtgQyNqzBrhaw7Z40m7+WQ9OPt5L79WNDDEMZ
c+Zde2TVCdqnbIcmeepYPO/3k59MNfBqluLi0DBBDaqo4Jt+ieekYR8hoG9fDiw4
YfnqFqOutAqe+BDhlycKu+vbLOqMh95MyCHK8hD4vstVKZ7kphN83uNZvCdkCVr2
ujzFUELw/uG/1wIN3WB6ye0hwiizNmHAgXeJvslM+ix+s5XFHyJCPRgoXSWGqIZc
6Q3GlRj7tOIO3I1ThvmTxCNoye7geTAeP9+xUiTcgXDOvN00win8z2DAmoYh5FmD
nV0zduBGNr3DMTTupQr4VwVih3fJHn61XjMwUtZYv+oPvyNSCF3AO5XlouqIc/xw
vICDjFAQIQoLA7s6XT+Gs/opDgGMwF3Irm6KhvY7sydMu4gP4NOVdyNDwD4DtFZr
6VGbTlFioSxpZYNJ4cy6mDgGUZ5aEG5tMDkkEFDhxVe98rHKbcZVuJMLxI1PN6AW
Cj+I7cKUQfiqM5Pjq4HovFz0LJMvahxRHN6ulJiCdSLnX4xOwpkHMdkNOGnBqEOd
Ihgkb8M6M82tSPiGwXgpZPnj75cbycR0O5BqdlQHYeNVLDc9eVRmXZgHXbUi6vI0
Pg+A+lCE8yoKP2GpotAU5cVsigWiA/FWAh6AYx5xknQ5FuUfsz9YDvgiLOAuRtWT
6eGVAlZxqPzbaHyAl6/4qSfZxZuxjGLtZFjhldKpwvKLXLI7rLMxt/PJYFYpqVJh
jZqVVquNJL0lcm8oDeg1l3MH7r0c36mDSsAE5TBFIXWm5UrGRT+ilCM2HovgXoul
M1EwyotfrHQxeRBYc1WiYNU0TmzGStyNpqRrrhDSaAwIfrUZR+qZrWo3TBMg80Cw
LZYx8QO4Y0EaehXdMVUk82KEYxwwP0ApX/WLBDIoYG2T1I3TAx2Xii/ON7vPjkx7
5U8JjLwG/6NhTMacUqjfMV4WnHppHqaja8jgDmH2kQq2ef+LQH9yuEtDxHDlAcpB
mBztsH4Gzy02VOYyR+WMlw0JsF50ghyn+o3oiyQHP1u3lQBEpVOEGYuTOFiP8YYa
eCBrVqMpZf1lVp2jSPbFLrDW7Aq+Y54tlsgJ47YKdIWDbFGZhkHg5R5DGRq70Wgb
WWy5XvDpDtV/JBAYd5+ifVD9TXOlbUArmuUP6Z7L/OtjIQZwgKnp3+e5A99YTPkQ
waCzzukoovuaerAmLzwpUlL03OkAcoCxV8B/OCV7UzmkDDU6hmjRc5fXaeveI2ol
b35QNtsoYJMM0jn7Pwdntg+KVlRZHApgDV8NT91Dd93buSYEog+C9cIbvbCoYLac
nmrZAwER8lkStTh2ItkSvRCE0bMoqd2y0aqtWnTNwu6QsopZi4q+MMqnQK8hpJUB
tbcPgmQnjPaypqk4e9NmY1xzdps1cnh703E+qh31qzY3P9U8Hln4VL6QuHXNJRs+
EXopRO3AmFcdDbHZPIL1GvHfcDYJpRZMHkc7pg/ZKB3LtbODn8kh8SXtoWY/Y2Rq
fWR98iNNgC1huaXhAu1J/U6xcdueP7PwtW8RdnnQP6NvJACNHCPphywh+dtY3K9L
B9pJLI8v/E1lnuORZ9a3gYJ4NzV4t11eAoDWX0RPrG2emrHiRiowCjCn6SMPCLLl
bI1ttqwHg6leibgxeOcG8BkoZKG6C6gQ2UmE09fwFeKRSI9JPsFgvzYJpknggfQc
HFd79toZBSR3C6K3hjS5T+rUOkW+899hYSVBs9NTvknPhN7UY+A/DtuYK3+7xjl1
kj/uMil/V98lnfdj0GQ23bvPzsFWM+0EIk/43UaIOMqC0KaHkrersH8aCLE5PHL6
of2hmbH4Q0MHg9V+8JJuW2/0B136rA6HdryMFGq59JnoTd2JsIx4pWcm25/nhs1q
8m0HVbwPaARoWKHyuFg0Kcv0c9ny5z3x0PiKTLVMQRAw7OmALhOItUUbq+lpUbuL
ETQpnbNkUdOA4xvUAyBofMHvz5ZYP7btf5CtjqltXVe8cNlcSG4+AwIqpWuCDy6P
XP5VAV1JNSPFzUSOJGGodGjiej+zaLNDMgk9nVV+I7qzsExfsB8QXHUJKhNY6gaF
5/EXdAYSZGaAqRxwDzP8WPOrW7/nVnRhJafKyjrC+0ZLb46hJd/wPO+UPvOVlymr
ixIDsBbHwGWGHTtuNorZMBz0cYhSJNVWe5qfUssEtsUj2pHZBKy7YLZ+fBTd86HN
f0fMgt9IHkrtSqZThbHtbsqm2loWR0okrjB/fOiI+CqEVCdaZqjVwV6h7Ym4HqGf
P7HH5ZMFADA5PulqoqYumiKYIBiVeg+Pv4ZYS3aksl4jrtr/P54VRN0noGRFjz43
y+zpg8k3sS9yM5KH8ghDeQ2AMBCk4ACHvvkFqyQaiigpsvcBDDEDLXXTBtuMhbSD
QodGWIaFI/gbqE1zrLom6uKAAWFjL90tEF0Lar5cjALRwOFKaZg4aSWaVMQi2ARL
IsskY09ifd9UT6J+5WGlDbB2E0+TElhgI39mOVnh1igQOmai/uTWw2eSYcg7yS/m
RynCkNTojpURNEQ7mv6WabKQxm+wQpgem5Cj3ifz5N9oPutL6JaO0FnebHZmvz2B
rRMs97aj12XU+JMrcpi7S6ost3KXv/GGOFDCnJAeoLjHaSapgmXr35ofhH6FrVbB
JZnV98XSXYm0Q8cWbbA7lsP0sshp+jdTAT0FfCgwupYM3vC/H2kJcV0uILlRHO6b
qr+7hZNa9iaPyYFSEgVDunjnaYZYuY0FX59B4+jQgUX1Q8KfczgTxnfrNzpjfNBa
tJ5ChQjxP0nLuKikeHqVMhXCMv41t94y30O66I/qKGFTuIMI7du7ZV51tvjzlYYx
sD00os0cAv1YrGkcP4Dz/bXkB7OQP/fc32DSXzF3O6BHGGEI8lReVZ8Z9beO1j0f
KU2zwPXQ1FedyqDzxM8A8nXhaepwLI/H9ewl0E+a2zopTAXPWyxAhTDbxV1X2+qG
i0cyVPNv2itTH0xOEGSP1cVUB0+Xvjvlj8EDRg+yw3eq4njyXl4MVyC5NM/wAQUF
s5WIWfevu3kQZxZ7DEAv5q0+ouMC/ofXF+C3Ihc1gBa+JFbEyNMyyVI7E3GX/Bj4
HqJlJp/bIJ3iXn32zQ7bqIeTZVteKjnXlTH4/IcUa5tK6Hc3FLEJQTTmLib7xiSo
e72S6RzU/oMeOyfnMFqOBy9vJjz2YukdIbX14JUP86rXkWJJogwDnlXE4v5zhErP
mfFIv2pP6iSg1TA/eCCq+9ADFXrLvPh6t33MSht1knlVCegtIKma7Wr7dOHn/+SM
RodTUWsLNpoyA8bH2XnjMJSBO30PE9y72qk+SMF/vF0u9g+iUev2OP8uWYVbngPO
KA3FOgZeE0ip10auDWAlH0oay+8mcUlIqqUANN1s7gzwuSqEMX5O+8FJl5GSyzp/
lEpijDEQGfQ/Wf9T2/q35Y7xSY43w/JaJe8/TCuYJl9RCRiyQftY9Iy9dhdPrKyF
1eIF7+Zexfj4+4/vl+hu/KrEtg8hc3yTXJ5RaPrH1DYbElgZxeGdnP9+UegQvbWz
/Bo830whfvzGIIWRWitweeszXxx2TxcS+NuU1cM9JLTcFItGp+adcD6ZmuvSS0w8
Hr8YFbY9q4NA/PeNoRWlreI1jq5xMxaApw9Qd16iwqd5gxBLeh3vpFrlbCvgZNkx
4+6j448tfFKnXTjLZqgLBLLYT1a9ekflU+93kEl9yrJGcEjXoXEWI00FSWaR1wpd
Zizoh02an0hT98lyKLEfTM1GqKxLSazVRPTkkpw42fQJhWpQYiCV1ATkBRD3Wi45
yNUg7P2vZLZO1j4nXDrGEBx8lZTsCTHmys+A34jWuNlAF5BbkrmsmajwIUya4v9p
J12mVDQ/gHt2LSGRa2FjvQjgWIePac/QYRZoigSja5/HhIUbswVdtiGquSYK1H3d
XdHEMkDuKN6ngGyguEDZcR8KmakRAZCB/PuOAgvsw/aZYcDj06i3yatc6vdTyPjv
6hj14cp31jszGzUEA8gchcGwKQhv5O/rMGjb/51j744SFSS++kzK62vsOaaXeY5j
sH7hXIlJgkXDF14oc0mldHrSWh1tHRJNsH8eLwDksoYL5Z1et7SG8EKvY24XNI8r
p8pJLcHueFSwtuGLKVejflp7rOh5lR0evtVmEzMf5HZTXGTxcN60KkrwpOHjpZa3
lxODbRB0WmecCU0Tg1bD7iZAFjrBKZ+ziXjo317Ch+B0uSUhn3fW0LgOGsvDRnmw
hvehOJoWhC2LEcJYJF8VVFnxcQOC/Gme4MdVS9O3RJH0T1d3FBtjRVlNGJfff7is
11ItzGTHOvqjwJmxX7Okgrb46/I658tzTSqBRR3dHrmEIQ/EZdNSB06NC4thqGeG
b9YjE0IHQJBnEFpC/l9aJA/o/VneIRh8NPFYEUlGFNgp6d8zYavkUqohml/0aGQu
9swGQCq1qo/++tdwrKP79gEz9wD3Zae6ZU/0Qs8gRmJByNeyZR2nlasyYySzivEp
FMleuP0/7PeTw1dt1pS6M423xyqrqDO4wVAOUMJAaxStRSCOyueTefJckgSyKVcK
+noBhDs0e7LtP+fHwcbmr/umlOKd5aFm0wswfZrK0KegSWkY15fvLRaQ6miHxrMQ
Btw7P6OLE5+ABJHuIUYk3xVUiTqpeARVo08PcX47w5cavL6WwLwbUM04AIWmrbjR
pboJaLIJ6b8yeBRgnfoiH7VwrMH9WVIxNge00rSmMhd0budVOycBetODWJC3FpAs
lPvfEtEsIjiJBJ0gYzSQCZ3xa2uxZiwbygNIDfFAFPjiKU1VfTjtWBID04pkbG2g
29eL7FyjoLJdlhMlAjHzh8n/8jtk/LV86PpS2+a2U4aFHq1QjjMIOWTWwIm1LDa6
s4iJtZ/XdLDZjylyxVRDyx6vPUD286mbLtL7qe5CzF4oJkRBhluC7H6BcoahMWNR
Vwa7r68YPBLkMN22KT7ew3FTcSOgvyp5sBVkBEhzAfOLrgvrHkYAOFmKKlE7HzQA
MpaiaVaeHRHSOuwTeFpr30EnJx3kcATunWT1PpW5kPLhtmlNjiNr7JMS11TywFYf
XH27D7jTUh03xbiJoKYsqc4FkFykSkYSqH9hShAp73Lkl6CR9tf96KnraM7yao1M
4RRJcIXz1Qo6azTFvD3VsiDoy3+01/t+46iIDSapGCaMd1LEbqoO4pDePLcHoNmz
zO1qJvG6uRXAFd5ugAT92mCgOkN4JX6P0PIKUJO4tgyo80AWWlMUklrnC7bVfao0
0yh1LCr6+x9nMGdpW0AOpTnZb+GD0gpRT2+Dh8pTzpV9M7+yAAZocUj7VTTAOXyK
L5OIFU4Ooj173DRwUJclgR1D5Mk86aNgCOUqw8ODKc3KxyrCcnskcy0rebGj60wJ
+I6NcoB240J6leBd83YMqAlLFgdJMqaE97MkV46EsXbSKzMJc4SZuE8AZ0PB9Lqd
T+CaLK2WQLqEaBI4D1KpYBJLl8nlbFAAwcv69zFEeH6J5qlIOi1554Yl9Wrm/5dA
lBdx050RD7pOvW4ozoZ9ynskTeaJSQMkIWSiPlfm4mK3rXEJMWtO3Y2hegW96Dc4
1tTVNWr56sfePi9t3/j76SuoNmfsmfsWQ7XdCjIGhXslCLlKDW4kMVw+ceAUnEaf
IW9NOH+fK7jOmf7/CQ74mPc8hCC6LPc3mpOIEw0Brp+KHSyjFMKKy1MQ83Lc33VD
cCq6iy2E1W39uFGcqct/7HM+EZbjGRCLiQKanuc/7cgzy5ka2IwS+IxZTB+uUxdX
UCm+60Q9i4pkCPp6HkPfzasxTrUFrndK+VZ5jO5vCSpsKNXo5jOvF3q+68TrNqZw
VUAt+YgW8bzUG9k329Har3gOKo68yvV60+3I1zJoNZrrpUrWEPKucUR+T3LzOkIV
OolS/wISw7hCAnRt1k2ZIKK64VwEfbsCz4D99gDSF73kkcmRzZVkamILhM7EpcNY
ZodrS9TElU9Iuz3jaVFgNEXsjBht22i302jjvSceGcuImLj58j6CpostrY4h/xbv
Yu3+JN0RwZL8WvF3xa4varDoN0gydIdahrO2ujg6LusXzgNhLCPQccOnN8pBqDug
MpMNDOEHerDr/D+r5/QH8N9a77cvV7TJwIxI/ud3QFj4dYP4JarJM82PqqbWFkeG
q8uHDoOvCBCbKerHpeHbAprng4yCsedvT2qX46eHARuyYTZtXu91icQxqDfKB0Tk
tmoNYF843sGmaskBVN6B3o/F3QK5tWbr58kwOE/pPZRVlkaqNqjcx5RoQeTcQUxB
GGFNEeA6wH56Vmzq+rJBiwa632wIKrH06+DzVwceWiiQJD4OB8l4VxqNgLy/Y2Ms
Dru8s9lRl7VPpnvulxGVYsvRSM5LqNpInHRmm3yRflI8G54s48alOIkffsI7spzr
PDyAgMp4w9jQ/X6qTZXK/Ke5Ux8DAfUjDiJj0hIggJa0AuTtraP3TQ3kA/IT71JI
YECg+vNZ3rIlGwwhpAy9WdrWUC6DYiobUsgn3ORAfFBQKwh6kj/ZXDcPj5R3CDZU
tix9asXj1/5yKuOrIsQmUK+31/iumKwUXenoMopgFar5xHpXHQq01YoE+cLneICE
5hWA1hR2FSORqRFNYStYKZa104vbsO7q/y9ykV2j04V56izLUzoEDszLPVPl4MJI
wkI9e+pETnKnJMMDXkPIts4UhOUdEr5ctkTZ3GTJf+yTmAyTJFZyVKPU2m4ydEPH
pHjiz8xm0tJATEt8AWbtVMiByk23gA9H8L6t3JTv0T0mub2WLpIy6GUVPfi3J6zh
G7N+SvU9svjEN6kejKe1ucheqryHhtp9zi9XQPSlOHCDyZTrhdNI3PvymYI7q/i2
NPq4+p+pPgyFqsT/qfkLJx+pkXeSgj9M2Grb885Pa1GVX6hL6mFxQF21zUoscsD2
+U/+ZtzbKOnLbse0IGl9H4kp/CPjUFWNDHl7M9PbrwKFkVBwwUb4zvsDLk/Z8QiU
96DDfIPSUITSUYlaEcrUWzmUapdnY6452AMn5XUyac5oFmZZQQ93lz6bHQ4+WNmQ
YY6/MdIGnoeQmsVUKLgHIjykjasutxmRIIL1DsS47OnRtjGvbpbRXk7nEU0084U6
qkyDZpni3befh8IkgEggmF3XHKz85qpspOfTnVwcFXaC3T+g74NugjFco0rFJ2W6
rY756L/WSEhdHrmiDoK+i3M0E8Hv+cDjGIocjhPMkMLkdcir7fXx4dxZMnkE182w
rn/WXFSXRvJJlZnW199BP67TlRSxMp1TvOBga5M/w5/64y+Fj0SXWZSLQ1AaXY+E
yyyedJBbJHQDZZXdmvXp7zF5QBHQdmr3biLWPTX1vkI7fDzwyJzEZX+Qgc+VDx6p
BU5gx/nWUE0MMhK/xZYeo+NywX88v6z3cUYLORLIbX0nJQO5R5Bx17JtOaHFu4Pb
fslijUSuwhNUXnhFSGpABDeVN0UCzVtVWErAcOywKh0pS9WWx6FTE2JfEpuW62Fa
7+bpn8JZ3ubYDo3tEYJs5Iv9Pat41mGohk6l5GmepE+KG+xP8ya9rt+8O9H9p7uJ
LLXX93gr0fnbPE9FhV5biXvcXBjJRDTf4oxkkxJF79DL19bx92DkUY8fXK2TjGHI
dPrMILIDJT1OjWybtQQ8dYFzVpCrWh6N7sDXCCn3Xi8vCqOZ3FsnSztiB1y6KIOS
oJLbOqNn9kzed57/SytYl6PhXGfGXQbAWUKXK32GJyC/VZaGsLXi7IVxk9KV2crR
AweUnrRoBBqlcHWjTHdSdYU0Q0//pIj0J/R/9nGiMtIAVG3dSdFq9a8ZHWZgw9H2
vBUs96l4bk9zV7vvIOnj8tKVzl4eBDCXlMTDacImEwPhSMupWBpheliiEIfIlQxM
yueoIjIGcy5nvnZ4ZnvYb7A2p5LPziiRp7jJFzJmfXVa7aXFyci4Y9X/VT3NpuJ5
e4vWpVW4kAtYmCXisxrZzHdAsnRe/dagXOEWrdag7AHHwd7vIRxlrgplvlsLTC/6
JmWJ/pBlw/UdyalCcav6KWBqwn5QUyTaNMwMxFg92LKEfMb19wVTZxzGMPNQFPsA
A8bbJGzvQOdKfk1Oh8uvFs44ahGwsvkSLjg7oVEUHDmmdvCVonIvXMrj4s2H3OR9
RPiZV9DTenux+rbSEz+EdH/Un9PRiBSfhuL2lYP7WpkcDZcXYmPKM1b8xlARTXsH
tFPAABWbfmr0F6/8Xp94MBAAbwSwiSZ6W9z639QPDzPlBlhmwklC4uHWUTm/dqDP
ql4w/rCm4HX5ovkVo/bqW5W2ykUyIGMJXsiT8USSunDKYXxEafWW6/MMdYyff7mU
DFlA8kgSFZPJLjADSM+NEhJViU6ElI/jyqDmLmPQjlVKkOoNkKMVkkP+0Rz4gWl1
cnDiQLCbTBvXiBnhHw6Wuwyu9dz/3zWuH3RAxO2qpSyNC7AXQ9xPcUiNqiufgSVy
IpcPXeeygdMxfqgIJAvjr8FpKIhK4rhQ7w0wRQ+yTWl6a2z8Pmgc2NToFCpou81q
4gqB+z4AnTZ/CxEe9AyLwaL1fVeT4eM4QUvyM+XojbGuGrSINqbaHa88TKAoiSec
v34JIYrXOc6hLtgVVXtycTdVgEuZu6eTdw0747RMekUdjzzfwGw5QWG4PsDii3pg
WV1v6Q9tHHCIkg5IOj3+/A+7DaPEcrH3CJJEApMwhzeaYC3/gAtVaOdTt+ZBBp2v
A3GzC9d+GI6dJICVdZvqB01X03VjtLQpGbnICnJmp99Z2TqiFScqjLSNkDCjgyVr
j1ocqXqsvCVji2U3V06e1+RTkXitKw+6ehebr4WNBxMbtWyNdT7fnRrotynm29PQ
YfYZjuX3nSz8vAxIZY61V0FdB7f5LISRdF3j73uZ+xcBBY4pNjW4ag9BRcOhzetD
LXXa2iH4EiZd1CaS4Ysr/+e7X6ii40YGonejyxjZLD/Uyama4xaX3qwTo2vNUWCw
JrOLMeNxGvIfES3N0D/Fwq5EmHQqBrVLqLc7RVII/3OokAnk60gGfxWU/o4g3alF
cQTVPDPChQH9cqefr1FrVn8Nt0N9zOqvGB4j+AUQrJnUz3EkcgWc42iza2aou6EI
bSGQHOJf2ebn9p4ByIKOUS6JqWNhN9h0f5BRRlCuiQVomHCGM6EXXkHed7DIza/z
V8mpfgIxzQqzNuLknXzDkWovgCBNyI4I1qyavA0FVBeFkJi3AjVrJlzgP6D8jClh
kj5mYBjBKJGfgybGaGovO1Z2QCk3Ys58vewjQjuYU4YIT20orwz+dQZ6+E0Xb2gN
mrG8abPVZ3z1H1CW/bKymsGDgBrPOPqkMo23eQ60GFKXi1G8qRz5aILB7+g8UUaA
m2i8VMfF/3/cQMk0J06Nm45aNLVj6RenP4m9EfSuolHtohZKAGo8UtmvaJbGhav1
A7BFEIEV1RsB6MOOAZa2uu3XRw813Vr+e1jPplJ3PQxCel9Cd1eKQZQI/026AW5R
7y/1xw7DH9EqOqKHNm+nDnSIUMKiuOfpCXow1XdNGnsWx6a29yscRvZicDW8EZcV
9wit5xVu6r7WPrtxhkSObYKPFKrN6Q+CG+hYASjSMLtBn819DFXvs4yOSSNjLbES
yEmugcXfBTeUuDLpWM4BllB1FYE9ykJ17wIU9EGO3MP0GqcUVeM5AoU0xJJIJs9f
2rI8tDca244lQzmceOcilrii0JmLQsnSiXAN+woL7sFGqnm60HiL3D6o8o6cP/6P
S5LX1ENgdo/tkBo5HP0CXJWJjKJISuIzp9BYrXEioUbJlg3hcecuhwo9etPSgFRX
zuPk59TUS0B7WrVAVhSJuUVPjd7d7UiVywEIpc2HxpsHcyJazQ+7NdksqGGGSQ5C
XdhPyUuzy8tGQQFQd0qU+mDUWSdi3rr4lyqnXRKmQ3dDhJAg7yWm00lSBkrW2T7f
OscC+0fA3LuIUjv/eyO3liBESqOtnV59kftXDIwD6QDzs/tB5Z06hX6oWBvt9UCO
CNbFrZmz7CMfUERhpIgWcVN5LEBbSTTU+8l7rUNBF/bJZmMSTFHihvbcUq+cDwGG
v4XvWbCJ+L3VRhADcr6/WfRQQtPlOyr3eh8u64d8gDlgSeGg0GKlq1n6PXm60Atr
82uuC7upU5cLqoBP1kvDf1eSB83OzkUde3j2RH6R2qv5BSrFTS4I4rgtXXkZdA4m
rD6pEUY3bMsKV2KvjvoRND/FUo41F5HL3A4NawyvaQWoGyIskcvbFvuC3C4L6ME3
ojb5JWuvzE1xBMG0I4X1jC9cp3rlFylwECIwpUvi8jn8pN4OjhHTJ+bCGUEZRRdf
P4wwOcidGKZ+Hty2q2ypRd/0jdY1R/Dj57QJWomCptloGL70fJANncsRXpbPC2K0
atgtB7XpqTVd9iFVa41R8hC+by1MwN11QaYfhLWGIG+cRaNQHLzTGwz+Gcb13FlZ
v8MH4DYYMxu38nKUxM/cbOuj+k95dUfrJpVwMb90aTXk37WTdzRM9jLOSzHhpHHZ
mH1XrLqwRI+Eavqbn4bMnKIEfYo82AacbZzt+ul+E6v1suut/j0exjwHQ79KYyNe
wcNTeV9FejbbiLAmyAyfCa6TVJoHK1AGLH4MwsYz8qNaqAJdi+AcmGJZJ9AqjAnk
CakS2PHghaMZWW/m30uQ1Z76z8uTea8IgRQTbNY8/J8AEJeKf6OFAZcQAcwRWwDe
hD2j/1XYMm39qs76L6wYncaAcwfVz2RMnmZNPLfAaCuhwZycW9tDOPLUhz1P/Y1Z
13ximz7Vl9gIaQdoxcLeGn53WrDE7l9Iw5D/Q/yfntW9o5dU2E5+ggtU9kRmzYla
7QFZhsabNnP/mCAS+LBqisY8rrDKRuwJzeK4ZaF5WZpgz/etPx53+m5Ai6xXousT
b3h7/zSuEAGOcabq2ozr6bMM9GYY8sVvJIn589DjE1ueIzM76QiKj4/Ju6GcJ3si
5RZz8jpC2NLhu9lb5zzXft1EZtdArnXjoxgAdhxrUWGPjzxXlH9rtGeWnT8DdXT9
56MtS2dZU3gIEu8dfdMZa0HdZQvv0KcAGeizwB32Vu14fVXNKHrjePydM8HgQw8i
1MZ6w2qel7KruN5Jd8+F8b9bb/QyEsQWY/T9bBkUniQlolOErFWXgjMs7cTkfM0U
Gs6lea3h0wPkY8kE46LCkQ/08XCGzdsiGPQogi8CPoRy6paWoHH9sLlkowbPQPnz
XRzPWoIJmb5B4O9cIIItHijA7BXPn61LDggXTLYh5XBzDtmweV5Us4VQKtVn2XrG
p1UCgyeW4cppa1tvU+Jsz8LrByKYrDwi9kEFozZVi/yjYES0wczFL8lkNFAogrVk
WFmevgtq1kpGTfbL1r3J0S1P/XcftUeCv9Xg5QgEOb0GqRNuM6A9oohUz5nSYM1E
TKuioiIMQ5orkiWFRgjhOl+GnTfJj3sIZ7JPdQSewkrnWYMKGGv6He16tzuxrPB8
3SEBciqHpw7iLeUYm3D5iLlaQRrICT/2BKFGEJtyX+dBiat4sbDeid8OWERQPHy2
zU9j+Hdb6Zs3k28MCju6y05/2iBZoW3kYDyJ/bfA0RXMahz6JkOXmt/irzJaueGA
3KZQuO6JlCRbvq+KEeIAOYgZCLrlFRka3NswnQllTvyOOeu0qZ8Q6UWoPTwRhmj+
VNJxdiWuYND/9kPweGAsoREwLZN1qXF9ytNFHaYuvWj7MtHTAmlQSWhz02NbStH5
di1lBdOhaH1xZ+sAzqJyQfCkh4TX4w2uXBpk40Mm+Vm+3M8FRkYUji/MttgMbqKH
CuCd0uCIhvEsM+qlWZTY8HxLzsHQDhBQ8W2W+qj+PGDyk/Ss6tUVhep1AesZf3qw
5PXNGY0n8w026OXauuQfH8A+gUl8B1vL12tNNVGNODG9xTuGiRC6DnsBi9OTH6+J
MbEE1mtDOZsOiNdrFRx9vhqiBnkqf1togASL4lwhANOPJAnFi0XPiRGouek+OZsQ
ncZxo0GS9VTRqOYFxOLnX69ha7ekfxdtrcnrgqL3gEUmCHO7yeTKYXU0wJBzL/kq
aJ6v5rOQToP4sBUcZAQBxil9m2svm2z0Z4qisVhrHgI6A7VedQM4geoeTWaFsh94
8Qa8Ln0IjnDtr59o7noOjvjtwmM+45Ua8lCW8RDvXdI5K8MieyKJyM2Xb14qZlnf
/WLADR+os88sz20v/NttrD92RbVLfwEAKFdBTm+Wu5kq7N6Q++LAZdmkwbIfCOAu
nstlpKsApf5XARWydQ+Ph8SSXqgDTmP6AY1C+VgnY/u+pSVH/Ns6BeN/NAppH5gO
x0aFzEF13DDsNIxXskJwD9uKW76jJ8wwYOZeUqsTdFlgWhkpn0/dQ4ncV+MCBoJj
i25tnav8w/IZn7zq7EO9s+riWAJ1pE+nWzB6G2qM6h4FYdqR9d2jQV5JrxA5wYm1
xHpGYGM0xw7e3NWT6DjdYpM+rWUmjVMG3ATh/T2gjHHtGeHdGHh3/6w5om/eyVtU
dFghtBGxnaJ6TY/pUFRfGTy30bsXvBMBpaR4cUibVfldD/FMAO28x2RVCcjlu+Lz
mR1H7n4KmEIguiey3zR2MFsvJxdhEfOasdm69vG8vfqiLCjvgM+r/bWm2B6J42ti
CmtDiZJPxpv2AL8CrY1VtULDCal4k7BKSpu3XkTCHsfVBhuWZTJ8S+n4oI0Q1+qj
7eYrX7n4oLMA+1Yoxjy/WTL6rgV4XlqOztRO2BHp/MJo1UZoSMaEOpNiB7r4STl5
OYlre1CjW3RoKvlCw0ilHkAdpWkBZwun8fP3U7q9VjF9Iwet2hpUQezTaistPzuj
bwglOlZ4E2zPb67ZYkK34dAH2cTrYXLnY4H6rRHsIzWwNrqcyrzA59cQs2B3vh4o
Bsr/sOzal4aBb+IPZKIRkMIoN0cGrG7Ci33m0rQlPy9D4KS1JCjO/XXF8NiagY00
dHh6YtC6Q8qyWZWp5Mwk1COWTikWWLbSY9VFyF4wtv6Ld1JP/3b49AE2cTm93HUn
3X2gdiHbGSbjJdANHACRXG2zUxxIp6BnTInDmyqBqRmZZCtdzHBQwEqQu4mz2yac
/qv9ngJ93EGuhcx3z4iWhmO0GvJoxhZ0J3RlXnH5bfuoIIBM14xUdU3DgccUPxkW
sdoIPnnpjvxJOHkmp9iU8XQRtysd+1f8ZlNcXYVTgYReQmmY3A6vMDjnD02WzlyE
BpyMsnxWHyU0ANr4ySUhkn/y56ORWrrPIDyO8zVWVyPQll+/v8Gcvol/sF1iJaMa
D5zcnA4+bf7VyBlM9oBA59zrk9Qy/jsQDVjxVqujWQVT66NU9RryUDHuIjy27T7R
k2rSO1WcBcjOgiuJuXugvT1AmwKf0p74NUPxGsvgP6xOngWjkX2acaG6Qiuy+Zw6
Kpo6PJ8iS0tqA5k4b3KLCsl07BwyK97dsyVYzKuFgqTiMiyij6yYwAG6hKUknKEa
vjvo5k9dnUp1JKxalfpAjYrm6n9F22ynegFLZMJPNICN7RQ74kSjqYSI/yDcFnQX
LL1bW8NsBy04pxwusn85+3EJLi0ZHrT6pgD/Zxar18oWuekWyT05ICeMvkjRS7CU
4bqpcShsD9Fjp9Caz7W2sp/Eqln/tNT+CET9qrK6j3lcX2NVewGWusihDt2Np37f
C6CZXrNwdmxatn3VFhC2BC/YgaWSXxC6R3fS+rau/i/CN8R1eXj+gCXSQcMjmO5A
MvBEBsqtJsRmFm68ecz4ibRTT3IZGnnKUqE22ItPJBc1jGLQTokc4mlz7h1NrRPW
yrDguqQlLJwk8hiTxfgeyETEOLTvyxqQon2MlUFWBLreanSdUnRWbXY+9UZ5Dsa8
CnihrG5YThQqYCbhTQP8oRgFSu7ABpRXtHDonkUS1HJYdfDBfjf9Y/qTxoPz49A6
6F7Kp6HRxupLYTsFK8v2/HJz0dOBmZwzYKPBor+G0aDqKf7Tn+WU2pxs5b7RDeFt
+DLZQr9hy7mp21+ZEGeN+sa5/6VenNRWclJhCpIJ5NO/BM8SyEfc8i3u426DjDxI
pUXrdBJdNA8qOQJh0G/a5UYMs8WOjufjrVF9gcctHh8lmrbCsINcwlmzc9V+80s9
rIMDInws7RJZP+6jVloE83w4MmWkHEdQAFO14TnUU5GJ2t3WsqWugEHmVIV5sTsH
/iVR4mIX5Gc+bdBUTdTxELTn5cmVFkwaWq9czsNg4OE6l3jV4uH/+UondsS7SHaE
36LVGJW/GHXEcqoYqNAJxHgGTxmJdugstSKvq3kXoguQogTFQEj638OUyY69cnWO
vsGEJjcY3Z+gBwa3GI5q2KxjMSgNY08lBgjd0HVxjNJQCi4wkUJjPRV0pgPzOIox
Hm7jhkpLVIkTnqBDWP0Dx19EKyUSWsHOD+A1bJsYjTmUq35LKxnNl75M5T+94gZB
hHkBzMDooE82qCdSP/22GP0F+zbGbWyE3WRI2WizcWLcIBX579naHaTACEdxioQp
IoCj+rkA+jn1467VXiMDQoXzEZsxjWELSJhvq0wG+OW8zyamjJDfx75TsyIuTgA7
m6QhAksK1PmwkRLU80TSkFOuGRGlSR2XmrwQDr0j9ezXXlzD9efxMCk7pPI/fCZG
RSIpSjRDbkZZhsqdBI0jZrKTqrsYWfDh2kVrV2+J3xHkpCN3tGK+vBBXoNkPdJea
52uCh1ehLl61j12XWyDj9EuID8sQU6UrGW81nEYxihwze0rdb7iGhaEJCjeEJWj9
cAk4v3lSx3HPPO8kR2FvuL/yph611kelWTDFPoBsjsvT2nbkuJjbX+uDjzrshb0u
pkNzVYGx2ANxbC0X3h00eS5vhMY6S5iWPihtYXSPY8VwbaFV/tyVFwX+1gb8uN27
C0RMt/D3nitd8xDQW6XjXkY07RnbATx1tgkBvhlJb9p3YGqLj5Y4I9pcuAxez/7l
gpXhrZOiC6xgbwcWtqb3fnlF4kwCl502NsqM5pOcezMD9YeyWdiQEG+y8WqiuOvs
oI845EeFwl58pvNUgfbUU0kX59E/FORqjWOXmNuJ20XGsZDM5QYr8IV1aYRAzI26
cG0bT3aWELp/u97BMWbKciohXKUKH/0ZEL2aWjINulOHCZM3pSb2SII+43G8ZeNS
zOJO10y/wx0CJWmzwbP50/wThW6oRUak3vXg0FHlMzsWHD7CI9NbdXVjX7zt7XzB
2xn7dKyABS9z7wMh04gmVFB9TPF5k7/bHS0R32w9YHvmtOiFMihsCoKMO7qyjnB4
kh5kn5hWD/QWmLUvNjABqzBzpzGN/+ZIwei5KFP+YwBOwPVu24V4ftzfeDavCGeW
r9jNIvfcSBZts7xF++1daQRuIwyQtp4UIOzoTwcDbYU/Virol9L1N5y76Nm2l9Hw
lDe3vhkgODb57V1TurFMM6jJYIfWoGtlvyOO4I0BlXKPHhKqp91SkMDPDSkO8euq
cyOaiPBp2d58VjhoA0+o3vciPYRT4Z9GiIq3rR9EpWbLHxMkjxxw4F88MCi8h5xV
iF1snTbmdOP9wlidezDHStlMRg0ikjjVFMZIIJ1w0kwceAa2PvMRZmfRXB+7G7iW
+/jnZHqWWh17UxgdlNnaM0EFBgWijqWqT8/tnz8X2uAiM5LeQPNBdRSaYTOVwI3o
MLgn9uQa8gQx4MQMiZ7fnHj+IDXf/4Rmn7QBvMKgfmNnOH3IwJPpZF+a+w8Js7LM
/12Zoagv16VBWQGRhy3zrHdPx0hKSLBfALVQDhEV5ZVUxumIYWp7Mu7XlEg3Wc7R
KyuEK9w9wXyvIh1rP4ZZNSUREFKN0PSWVg5mMyOv9kvar3qQzNB83fpSdRDL9Gr6
JXX+4HYmGk/XggW4X7sgbkR01fDKEHyt5Ee3TcLOInXpBq9un4byTtfcNM25JRay
Lsd1lhW50YRHnMNpecqgVwQkMx0UwRW9wdVY8LMSr55cek2x7ysXrdIMJwuojxoH
jwhuMK61TySMuFLMhUKEecb3qkWTeoCFudfGvoJsvkRxccZfHFvW7ksnzH3OR7ot
7EpuwtiFk1p5v24H41Qu0W7SKyDkTEhyv8svwZFV2IAw5X/BxmngApAqKQNntFGN
DCWFQhi0CQdnCwndPTt/A8OmISuMrixgxAM+dtKsC+pS1WfcX9a1otiPKYdhJYEi
/J05tE1NSfHfatb26+8eCfY846pD2V6beR3jI8sMtgTBrZ0GCjSoDbxkzrCZR3U7
/klLDxJmn0AOofj5pYuMYCts+TFQgh710xeFV/jAr96VO6gKhMFimI/lUQaFtrhx
0KAmOlUss1F8iaq3JYFLllv2KX7Z7ktPbTg9J0hOfU6JDv/e8xQiAmIIF66qzBSq
hIJmYNd0zszZv/zxPRo+zqGz++LUmbkzFdjlCEUZe5X1Z5hW58FKpW3x9nQym8PQ
0HxTCYJTJKxVp+hnbuwptdrefbHS3D8gbezKWVbKr+Dzgx13zTodLlFpDoNM4VL/
/Pe5XOwkQUibNWQ22R2AGcw3Sp7bI5MXmAapCyoc8u+NFswcdI4KKYkQrPJqjxF+
7axMBv8V0nMp0m5EFG2qjhjS744yw9H/B2ZqNRi4Y7AcWo/izDrZKgYo3RqT30N4
J+Bb+dDCH3pJP8j8fro76y213IfSNVIFureQxTOWdAjxdGNiohSXYo/aJMHkauPG
nbORZ1T2JdF/TEa4toPWkwvSCaCgnvxXXLVrQgLAKjWZO0zuchXy1sQ0IPdxPkrQ
npehcb7BVfAo0Q2px736nz0+qdkVC7sBlbR0AfOaeXIIHkWivKaugS/MOMzxRiTQ
rv0UfqNBtKoMWNPE4jaMMqpCmMMqXQMBqI249zQjp1Iz853htmUzX+P2vBbKIzpa
3a7KNp2lmyB3HHq5BDhVnXdPaQuc9tLUe8kk5CLJZKMz8E4e7ZjVu0ZLyyFCJGoc
7lmyWfztw/CxD/gMb/KslVbEb96WEJdnFGGUcBJeZZwrK4vkqcxHJM9HQYGV+qv9
BUPVIwvZGYUeaCI20UI2JW+Z7bk7H4PdoAZplXIMLkg2ZvDbpRMkzXYpQWlDHB8T
4MTT0cXXTNV9Sh4TinQjWttxxIwBIHYLEs+pvgyqnHx/opOCQlez8Vupapcq6Sdt
pRJEp88Bs7cTHvAyIIShA35YEB+YM1850ahg3SFpnYms8oLFgH5D6M5OnDgvxoyB
k7mU0f2tcHr96U6L+VBC3OoQIYV/42On8p8KKelS6uhdkMxW5cevStl52uQt3Siu
KS7JehUC1cHw70PQaLCre4brnP32R5pG0pEf0kB8/ab7q1oxEpqKRoXKPRIvMEN+
wAY/wLX0saXb6a/rYNUE/76BddM5Eiiw9pDrY3E9a5Sdll7zZqrYNwglDwF9j8WY
54LVtOAOIcJyVJnYIk+8NoUb++LUInvRA/rnbO7gCpDo8ro0TqSe9aefiB5hZsO3
PwJYizxOW+W7/bUqGhL5MV5t036Sh0cy5cci2UoQUdvyXYpMcnD0J8Cj0vl+PxeF
hl/iKUnV3MEXUpUZEYHKzauE4e/tE/D2ZrbKo7ycvBtT7qX3ZvNrSLQNAbP9WFRA
dI9oPbmpHgn93lKHUrzGbdoBiZsvXQWlAdske/QYAALsLf2gVUi1HFQaskpvy31g
SPcQAMYxUHkhIJk3n12p8SDSBxuaysxkaBYTKKO7qtwuqps14adilT7IWdVL5wlB
tx1+1whp1ChrTboKcRfOp8VJFWa5rWq9hQNpeL92D0/aPKYgiO7+egeQ5NCVD6LU
VoEiN8ySpKDDh2psDJmS8Zwn/lQ7Dvr33A9dVzXSPHrdzluiIZb/uiUsvDw25EfX
xi4wVNXQhHqck9ndsdPj/gdrCb6JV57OuUVZw1Es7cewrNrbodSdCUabJW7Ydpi/
GXvFob0NLZXzquPwCVg+mOfAwh++rxz3ChxR1ltf63oTwSllAZhFdADBiHCitftd
55iDRhQ/0LiEWJDttmtEpHRmo4EBD4xvEw3Hb0LSPmdVZQ3BcmnvJstKtp7dIN1P
m3Co7K8SHpFun/hR5Z6mkuSeLRWUw+UnawIBhO/w5SvuVhbf4G3qdGqRZytiRvVf
JV+xtquI21cj3q5DYnn9DnoaPKceABwi+Eq3iTsbVAVkPooLk2ggzXEtZkm5Dlkj
x/w65t0RFHjDbTk3i+8o70MWsWw7/Kq3+5LbzSHsQF0h5Ma3cbBhd6PLyudBpRan
DXodO6uX7f7W+VV5qukCj0L2qSNwC05wf/sI/jBgedNTXUt96dzLYTf49EfMJmCc
8xC25zBlMXulnasEUcIR0buteSezuVKv661M7Ac3IpM2JYsNjqsZSUwfWxjnS2k9
j3g4H2OaNuTeuKplF/lsM3Zcy3S5mTaBP3fzX9HEDnHGv3NgnE03ONOzA57nYzCp
VxnCFUxjUZMk/cb+jjYByW3WyOc4EMcKIJ9Q94LUHROuE79/uDqGfUMFJQU7BLsx
XJGa116cY0ETeMI3MLq2XW4EbqDTIQYGEBGwI3hGZ26Wpw+SFnPX9EvCcti/ekDp
yDCqdKLtKTd7vaA4KMkVqhe5sFMZzbhQrn9GG3LIafYeRdEDaJ/c4Hh0Vo7CGpT8
GE5PjEE8JEFHY0T26z9ZOwoE+emWnVJF1hdHbaHwowD63xjTB8uOZUsGp6pUOZMs
sMoX5LiAxdmHSbREOFGH2Nv+jObdK7dWKtS9bJbNWD4IDMbcv/7k9PHvz1/9tEFn
pA7iTw2nQahu4HULanpp53pkXcisPFWBi+8cMJqGKBJ+kfoknSKv6C58CDPnPDmW
BWoW4M1mq3hbmfK0EYREoXyyhYiOPYmvzAEuDyslkgre3G0jaWMNwiEeCQxA1o13
qw6c69iEOmikW+7rqpb6R6A8AwxmY1LvMgBKjo9e9DHFh8EHawh8i183ylS+jAF1
TC4orD3ykUbl0tbZR2pB/1mDw0mMl35ArXBZ91Uk9hzBcMOHT0xA/g4jBNfnWKUJ
Z5H7dYtYC/7cfaB/itscl6z04GY4mRxy53vDPvDulJKP/wTWYABQPqRfeUhqN/iF
yrrhy8DOpldSCpGAzEzAf2cvJiQsl++why1vh23NBJcHoaD1hl24OcxEdxGbDCJn
qPHcrC/KbovPGncILB8yPqRrngnVa0iyrGzliwmeg4+6c8ZQ0Z/G/q06sM8OHjrt
/GWOwe+okUIE4K3wCx5vmWD98el10mOrVQvYIkuRpNYq1lJtwDp/PI/EinwNnwX5
DhoglH21EdfMRcWOkpo1N63zuuB8DCgvUJ2z+cPG89Udcy+26fNZllVRdZf8jknj
OCz3sDY+F+H82ElOjaUr23MdXeKZhnCsx97VwykEAXhcWge9RzwxxR/iZvFUzR3G
V3hPQdhEqA0bb1GcBPEQCcRMy43oBxNA3IKc/N5MgXBNRDlaNjrA/cN49UsvKzeA
YOIYR16ynoh5mS2DBFknbiuKPUe00Lh3dWrWQqT4S2vJ/YDgzJ0UHVpFm3CCJW0p
poo0TZjc8YmnRebcdJ5fYiZlalyYntWkWrAFu8WKckfZCYKRcoU3TuFbULNxvsAc
lWIAWUagBJsz3zqvO7p+MFfCA6YjxrbAXHAORWtXKnSPn5+p6dnGYUj6BDLO5O6c
LiKCj8rhlpy6S/bQMYkjX48dIsLu7g1f4aPqJ4HcqXlsMWjmbUbNCz0H98mfPgRr
oBYHJ8c0UKt6XvRvKfPdvyduM+TABa1cAnQE+bC9P5QxokVa/SXs6ro2Sb9rxGWy
oBlFg+Uu7KX9Gqgck7HXMq59ezHs10p8qA5ypnud3PJjMBzYLt7FbJP0F/hk/QXH
BmErgKADwL9FDdJAf1oXom+dSBHApyRQ3pS6ug8kUR+5uR773BwNcbYGxNpCE3DG
A8iVGmNNpMFonIUPH3zf4b21A+XFLlfxvD2Uft1ZEYlkSxHCV+eD0VdRfJvab3/l
tjnC5+6S2dMIpkJm+FLSnc7hrEQml4pYYiK5sf3imfiaj7RT6ZqJpsSlmUBdcBbM
WEKccWQI0swe9CkwSsNnEN3yildscsz6sT4VLpmhLD+ARMa1H3qQPLj5HZv7bdnI
5Vfy9YGI4yAlddHbUfAY+RQijLGNBjBg1mMmfJuBD080Rtxe8YBwrizfEyuEm+Pk
jAp2izI0iTIVRptFao8lsFv3w+YaI7CAy1+EshwrV5FDwnxEFTP7+59mKNIdR9N+
Yp9oJxXqzYOEzTBruk7G8eDwFvKjReleCquGNAXCDvvV9GbgejKzgcYGIDJrmWfM
xWGxEew2s/EVPBmjdQ/wCPezG+fTCT4vT8F70PpVeYTx6ff/DWSnvy9zdcG1PdzX
jsC4XTMmMUrMStd8fr6j9IEjr8QkpRNM4rifvbjPKfSo7cE3r09ItdXJ/dl7BzJS
4IgkAqQuVQcY43bZ1AxSK3Cit3SfYrbcroGrfsQ5t/VGCdSjtEM2XSBx8jDywNqW
MzDo7d9E3u+Lk8nbLfRgFKnbw6waJwx5rVMeY75a3KspxEu1Tc3EKQ9h4pzyH1aa
bnJDqeD2NG+1Y9wNvfA0Y9Ww5g2bDerlZX//21e88Jh3N7362kj+9A2osZ2MJXtI
xt4kq3FXltx4UWEBOdFY66B5fUDoUgl7jk4LXdT9HLDdY/Srwi6DVwjDObcfPwV9
v7RGaJuTWdYTq0rZczlbXORsYrJ+OHaW0gSlnjYtlWog9cjK+hjdD4ms8mlSnkPk
iFhPgAFpR6UzZ3gAPczXwg+RUCA/gacbkP2s9qAxvZdPw9hhybEZZkWdv8WTaN+4
+dnHCzf5ct/UFb3dgczeZUCQUoFutTGKJeva/7qYC/j+TbVDEtpItu8xvt5JFXk3
ZJy/9khYVuLS00bdoB/dgTqqLrOzwhKUWaI/V0qvHAjDn1nakNTxOVFj/WJgwBRb
DV+IAwI42zlzMllHXRo/cVXRmWmDRyzve3r3HqztItgecPsN6dz8zhaEgET4kivF
Nz1ZQYwUPmguNNJxv7rLixoQWJ4dAy6I2kuh7bQq4pp3/cOrU7ptszNtb1RUWVNt
qKY7VOc8F+n/WkQ5w6colGPfnRrP8AZrPjXkwrEecVzTxKhqVrIAAGPVJby7NMY6
Nx0h4uSs0dRmkEqr1/II/pUYcHOOEzfeN+hc/8raQCexvQaP/u+QA/L879ElAG/s
zdls6PXPQijk3a++c22AeUhKb7ltQMVrRyF4ApMWay8Qxvf5q0fg4CjaLAL6kx9+
BoUqSwXCtIzwr+YRqohlPzNbwM4h+GsUoaix8m56wek4gByWkVND3kaX7q4G0QgS
7PwcJt6EMdvWdunLckLOzKAdoEeC3TZsnJoemjgSJ2MTD8ZN97gQ7CmgzgSk3CzA
eDVcIJcfNVi7k8tHXZpV1sQCmbeJnrjPdH0sSrRXhMAYxOn4+PPF1cvEIQdFnXPL
g4xiS+Ua7h+dfrKdLtofBGotFbsFtU9CXGYs95voWeBt+jgs80CYPQw8t3wnKmOL
SMbaWZzTS9un4gQ67jg2i/sz+tfZSYKs5MHAS1Q5yXw2QnXBluGa/aa1DxDQztNw
jRqz5Bgj6RVT5nSDTjqtdszatc3JL+5R+tMdq0knoI3+HoKD7LznZkHsinBbCE8t
SQZ+OLVXi/XbdrmZtz5s5KxWAOXOJsma8Efg/mTCYycxcA6/1fsAyo2nAsQfrRya
QQhcX2BL4vrWqUmaw85mOZdymydax0MZQG1LV6aW5i4LEjt++xB3dZgDAE8/eBHA
Ddc7PQ1cxXj8tfIt+89cky2wKiLe8ehKZYa3nmDjotcb8TZ5NQ3n8y7VvcmJUEMh
ZOE6AVcwec3hGnNX8/v+IcrBoGv+i4z+FudQSpKs/UJTEabXXe8veoUkRBnLv4se
58DYWfjXnhoRQKnuXoJfi2bSwHzO9Rt41FFIW9TRklntZdjFmih+8O8VsqKliImb
K+bXUqgMYZq/QXY//PWMRGKy8pXqGtMkUsJ0fR9xPlZtGPx9IJVO7OS78Lcqdglk
WEOAkyAWJN33rDMGCga78GKPfkTRcQFaOjyD8diYoIVlInMICE7MVSCzOWyJ+Xay
QXhuXT50ZHQ1EBAxj9w2dcy3Ng8SGIUEFERW351zIav+OIMrdvSW0oApwmzVJjik
dakvUDLEcN+ABhVLcYncfj89pgOUVjf9VK0RUTmGDz0qr+PP0yn9w5jiP4CKLFzl
8hbVwq5ZGHaq4jLSsuXIOAYrZW3NNwQAHloXCNOHBDiCkX0n9xmpsHyU9/bjP7R4
gAFuUbZ1T18oLlnckyc9LDkyTrz7RdgPLRsdaNgIyqX41OVJ30J8SJW8Swr0u8Zj
w9iegh8ZW+7uaNZmcE2dxTXXnYc20Odyi1zyvNLKOiqiYAzz356Z0hO0BGQg/2Xp
ACD2Ar/W91z5WCX/GULAxbhFsIiYQykyCuHEuaC2dmiwKTOxukQs59eDzgBIpAz4
7pk7SNw2hiZuFlGlFjuoPBYkJTluB/w668XHfDJJ6FpMmxlxSjFDn1UgT3EKt2sy
0iiviZMqWcoOYqHzDT8H+K2BEukf5rTlnVal195UN2+QI8Y5TLuxp+fu9LlCrS5P
j2Tm0VfJIFxlCyNXBUiIx1Kpvu5EkgwurpmOsb91eLCTLh0vZ5wbvEFBQ5ouN45b
MJw8PspxKXqopS7Fw6/OBWT45BwTuHzcI1RUsdepkuhMMbsFz2Bp8YHdooD+Gh5m
N5EgeiAmu1+q8IofCWrGs9SQ/LgCZMIT+PI1Nt2cg+UrOIBzBZrg95kS5XnHV2ZI
vSZy9ktnQELe1irNqlmaeKEWbxN5aaT1E/NnEzsetvRosI4C6TGk/WUAaUqfA3o1
JJ4uTTGwvhQPA+p6tcWKLn1MiGfQRcv3P9KLebqz+7tlQerAJvR8Csh1YXtlVzOi
8FcWUxLnpmUevKpDfqLkvRX8uR0lzXsz98OVS3G8wCbdfpmC0Hj4dMtBw7hDrNeD
zOwdKzerO27yyMytnOX5uI5kpsSC8Qu0OSuAwBpFyk713ksbl6fJgi9a7Bi68BwO
D16VqhwCXWN5pR1Q8NVKOAA/t1utwc7QvImMnZ4IBrXVJ1XsT+/netmqVsLMEo9F
3YGgBfV9lx4sUWe9AVtBucDRVkYsj1FHQ/WCt31JajUgCGw+1u31PkuEgZ9Q2XW4
njY4b8V+vHvitxYb4akXjl31z9LyDUFJXgtl8vZJ7yBC2sNBT9wpxU3A9AnddCoZ
Kl8qG5UozDnsWJVZJZ1P2qLo2B2543Dx1FiOknp67gmpcODVGNJXHtNRxivravQJ
15VIGWqhGj2NR3MbWUm0z08EQh+Ljlf/kXkzB+eoW4MUd24F+VBaiOJSJCXH17/E
27+9tMwqdQ9LRWIRIYiveS0a9HqUPQtMPwyFhtGs7uNShrwy0S4xBo23OgWvE4xZ
bWn5CdJ2+BVun8Fi8zi37YzunrUARCl73n/uVw4hUanzmsatj7DWfg6xsr0HFndA
K8+6HI9+hMzTKdcTItaoiNXTeOyhhUQfnkkipYYya1Ufi2FxqGwDQngQTECcbPtR
uSjGEM3r08GVrZkqg5u7urQjaksNToDULDl23IP/jxdC1R0QF12rbn7r2jaNSzNR
MViKvtSOCNHfCtP7Sy/O8/bx3nzQGhGOQH3c7t0Fo7aWHdofZq+LXWEBkK1tie9L
khEiKNpVLgfZD1VTMojHIiIBN+dpZDpqxSpBCLKMoLvYfKZdwUiNlhtBf0gEehWC
JbHwv9T5DlT0yy3PnQAhOM/g2kz65GkR1Raz9Hu0C07aqdV1tQZKAXH12Yv+drz8
BbqvecxqwU68jJeewZLiNz6ScU6jEMB0t3wnw8pTORMOvANOoXdHIoQXxkBy6hIV
eibHNkL1Wv+Qzu85lewxrhT/94sBlg91VFQv2EjNhcTewX+uJgSiPOmG3Yrb9XSx
C34RnLF75CTkQdWZ4WuoV2ycYdKqftExZXDheas5VWoURtNUES90dVytWPajTlr3
/3Luwx5+yrMFTogczhdKqPArIRnvc9E5AnfGraToXGiJs3aOKsfNW7vR9UycP6zf
RMFuMLKzVNRQJ1bbxkILmmJz8zaH3tm4bp/cK6Rf1QJOvhRoSBV3KDiOJpZxdR+m
oB3Z7gHUbSlC2OBlFWcHL5TPSQpfTjHGbm4abJL99wO59oJYmL7Z4NhIRPDzt+hV
n0i11isoj3SUJ5jr6RdxlhDcjocHDO20PVP5buDXQVfMOLgb/U3dxb4GEn885Jlj
YlBPI2rzOiCza/F2WtAWBWqE87B15WDG4jp6yvk5s/xGH7j0EWGsYdi5Yn/GB+9M
1mRii5nzwR2SqxItrYnrtnC0ealU+HlxaDbVsLDHC1VH+dBAYIMlMfV4jAOX8tb0
jYS+4ihCs9SXjG9us6UjLq8T0GoGa7NXV6NyYjWVeYbA6bGCMyaagtDSSjY4U2Uy
6gylDB0FDgcHQWW8T7WSQLCD/8TB8trXrK52+1BklgyLyhiR1a23BiyZuskXco2j
7LZR9MJedU/tzImJLfs7Fx7kcYmSgmSS3PLie6wGWrSpfgfuAsf30z1tQf1G40n+
8cFP7cm1KcNphKUOl3LUvuMYPyrdVZhnY9r9N3FEWBrzkbegmvhfd9cEPLy8lfM+
LdEMWZZFpni8dwo4N2K05D6YyEnrIwcBsZyQWeQFHSd9z/MpiipbxTJwnZBJUHbz
3r6Hn/9ZbsFnJXpaj4Bu+ex3qWuES2f7d5HnS7vpXKDLCDtl0vangtQKijqoo/nh
RhOUKViwAt/2pbHXJNUFD9ymUP/jCXl6tcI18yxIFnRO2Xr34TVXEz52dNbKp4bY
E/BELkT4TtSkwctXQmODE5phZd1Qdub5tOU+b3P82roxB4K9FZ6zitTcit5jauht
/m9aLzcDn6MXd52rvqyWKoXv6QX2SzTqGx5u/a+1GdiYfdHilWCmGXUA4QEc8Z5w
o9enzBRFNxtIgzrXwsnMoG+YR8W1pk6ZKiYiz/chkTYjVuPOncjVUpxoPWxxSPH+
O4QfFwXVL4cI9w6lJsLNc1CmP5NnFQndrupWmpSCek744njw/LJCOCCeGwN+mYpR
SyJOzbYrJSIkO5b2Sd/yG49On9VXt3MmM3n2fwf9P8Q5G+6fXTELTh6sba/7eUlX
aNlHPnWFCkgOIsrdZLcK1yCLd3gmoSrWtjgzjvgcEe/vDBAlJqMQSEbNIGoiSJTB
3cj8gMm2noF8UvYvxcB7+bGulJ52Cuur5aH5Y3JGCY7mntzhnCtw3xKfKmSvV6OR
ncEQY/V7YZ/6Sj35NlxLIPzuV0xQgfMcQ/zzqAt5pPfLosYcLHthQf3ZQPTed0v2
7SVyac0qLYJUSGC3fdFwV0NpIdftwy12yrvVispK/GIjZTHYwQmlxYPPm1stYpeA
nR9Lua/0uJqO4Z4AcCxHcARROQYfKlNe9llz/uyPzCu4bU5eeWrROxkYCqrN7jVP
MHEbtYTCgw1WrmMxNl1E8kz8FFH9TRNruetmHVtmzyAy/SZpGke1J26qVyR5p6OL
+RGDoITPukQjXgl+qb2tu6vT60FjIkaZ2gWrgGQK6BmCLuhtE8xafD6HFOccshiQ
EKSxJyCpF6Y9wCn3o6oxegXnRX73HR0X3ikmQ9sUrWW1qIrMjx/8B26toauYATGm
3BPTuWmqTSxxGuUjpP2Vl0Up9snFqVVlb4MXYTV5a3lEivKWeGoebUONKWrwIzt3
HeBOwsQRVYJy1a/LFNmL26HTmhs6HCC79cIQvBvNBzhdyCMgpNxlM1dZRaADkM8o
xbjgDLxJz4/QS6TkpO4UdF+1HreH3M/3DltrBiXIU9lKgInfZcrwS4IlgSNgBr97
CzFvyrqeX0ZqzBnBenlnjqINs6JqMZTz9cvGDsPoxdWH+KYE+hzFfilUZdFo6JHG
5APZYRDkpNaDv4i6htU+5ZXsrPdtbJjSxXAGmDF5LytW9V1KLn91bNh70Gl39hRk
efba6QxDfRUMnVlVZiHm47adxibtvHTZxTc0Eoom8mtqlMCC1uBvtPvFNvLcg8oV
MNZGlnVxvV1ecaCS3O6ftokJC0InSECpicyEZn100b3TbB34rGqDi+Qd/Y2lyC6N
Umq9iwQM6v0oHanQB9S81UpC/n65TghW7Ff3zlrmWSD8i+MV3cggwk3D1mLJxNIq
N8tRoRs/wSBQ3sKqr59Ns8RqTTfuYY5z0Dss3gg7V2ujd3qC0Q/tHshdLuy1s2Ez
LJHtcU6i0D53GenWUB6xvh8YrzCle9z7No5QXpuFxzEWMnnJro4gC1szE4NMyIvw
qVCtyQiIP/YRQi/32idsjTDO4dSoVk4q2G1ZXAqZHNEBl9xYkaDNvkLidrfMwl3x
2onRtV9DjqHXZwKFB+ZzotLFuJflRSiDQLMpsh+vQmA4WZwAbqk8/KlKwdSenyjd
0y4osrmgNKGGyr57h+upEZgiNYKBBsruVRCY4dCo8R4MWZLzdF20q3yC8zyZqWQM
S4351ppdkajH9LskyVkLrWKMXueF3H5b9jP/mz7oRKNGleUzUb6EOyWJgZbdVtfP
LsKttVYG73+V8qtvZ4GUZ9u8cKQ/SgkkwhRYAH7vqgzSt5rwae5qb5FQrGu+UHkO
UGdY6c0YscPekmmg981Wl3/UR/+RzTd6eVeEgH1cnkZs9UoypHXvgwbdw7Qy5M4e
ILRFZlUEOJUAoHMm5ontsidwAlCVDoWtYkJMWWAWMQDDhlzdflNq0E2yAlafjHtk
doseEgMUMDCDuU/i8OJW4uCQUamLktrx9U0etTgGGPxa2tC6yIB1/ShGMF4RI3SF
hVtWLrGlhPXWiH5CiyVwFrKw2uqoAhEHL4c+QQ1u9QSjZOOB6dN0dh3OEhYCy43p
QTrO0FoXAph8AXLih67hMVV1ULkarr2Cc3XUtfUZSXmG2gtctHOr+9+ghhBBcD9h
dh3NlK+ffFHu9m7kLfi7YfzEOXz+zLvXXgIQXKa1xRJvm7TSn/irfALcw8SPmooi
sWSqAFH0Qsm+yypoAmPTLIHgnfo1mmVW8WZ9yCzUU9IVJh2kf7SBwzThBPykd6Gc
6s1N0wUjhTmFKBwHMM4h1vrPUqnbpo/cI6nMJElITvvNvErQ063JfNV9Fp2H+dQb
MCZ/s9pUQWViVow25b5P418HnrJDCpn024E8ES+R5geFRU/T3n4NsHCxABDgDEU1
NvFP1ZEqiWAq8KYQPux6+MdINeYli8weN85/Jjvbi+Ve583XhZVX4/yAyN1yhJ5B
2ktZSfAEOfmOO3XJzSRf8NZpcsxRG9ThU+kegCs7SIsiVhAejfgNMmlONwb+6sYb
hhK7uJc/Brw7Ma6IQdbaJ131ZEVZeytiB6imklrAj197Ng5peuFudHRGUbPDBmD3
0XmXCxz/cgAKIcZnK3DYQ9exo40PVjwi7urWYAEg4RxZHRbbycYLQg89nVgAJghm
MhAizrTsGLDkQua8xOdKRJu7t7gflM4V+om5z6eDsOPYwmS/NpVuCkQ04cz34sYq
Pumg0q+ZnZrJwZ3xU8tajBNIqkFZ2a2vkSnHHrD9b8E0zjYuF3NY2A14+AaEN9aG
wpv74Cdln6wFjw5fs69/W9CiftYpgtZg+1a8L2TawT2Y1CcRDzn3aaAkksuBJXIc
pF1BbLzCHhMSLZ1/wc9pjmLNVYyZl6HmUBKA1If6hql3Ca29oHAkVJib2uuy3RIv
hMja0za1/cebScRw3LqmmjcShLMTEM18AtRFD6C9YlBpHMTLiFNSC85p0VG2LYwC
kHxPOYD3FEq/l8qC4vmX4CIN9EysgTrKLj9p2ShnfxhaoqIraNFKZ5WGQa78lGiA
zqVLZZPUOW2Ph6GKvUS7BGOOc1vW8K/UJ0crbbp6C+Xwp/TLdbhNs1s4c9fGrIYb
gTcHbQ/5SlUNJoHlKyJQOc4UoC/T53FNWs+30yS91F+SFLd+QkZSKOfdE495jLVg
bjwT78fzhLkw5HR/o1vcT4kLAcV0b189+z8AeO7BuHxMz1/Sj2YTqNAe2vQveZN7
sl6RNfvV0+5BYmqlV3qV2gnDglpGpBFoaKIbG5JWjN/meYcwxgYJbE1YN5O4y/uO
bEpf8n69GSmMRKEMTrTU32x+qeAEzIxypUIqcNKwhW/fV+fmfNui7TD+mFOOtVkS
HFDkgdK6Aqhxl7itq+bxRG7nTLqlbEbxgfMyO5INZyUlGo3Hp6SmBwEePP2cgwty
bNC56qJc8xVU9cbiMVVA+L1efHtdUGnSHg7rQ18JFCDJz+mtiEGg0LNpdjvlB5gp
42dOigxGbKmKk6kHfBW4KempIQIJ5hbJsXP61qkOPkrYCAdgi80Vg5dxmLWiqYlz
Pu72r0xqe/J55Nt6x+kNMGCvKnW4mKv7IGkt5P+0jlFf77SgFbAF6q955xwyHqdY
YQfs3WyF0PYvkAvgef6u2sLE7UP5sYZwUW5YSKGQ79ZvBHVYiCxzDFkrIFe5XTGi
gPmCVrTyBa7aibxodR9wQlmj5Ld/gyhMnnBNcb/AkFDpMz/BQIDc5wwfS99WFUUn
L/YGFAUBVIBvaz1FBIEC22wJVgq7jCMj/SVMlrZhtHoYauOm+CGb083GbplV8nFt
OIHuYlTAXlovLVuHqV6YrvFXvg7j/ieyxKSzCIMA+XhCVuVhas3sZg51qgrgAZK7
P3ZQ1hB0abu47AneQF9jS8lQrK3kLj5goG6iM/E4JzX1HGlhX+zL6pUakmacaXgj
7hqyrNEB43zq7vyaP8OuIZ94YCsbOR0Mh26iRBOQy+MVwAy+x1h3KjeKNlrpuSSN
t0UM11f3hTF5b9SrEDonH3Zpxykrk3jq6pflFGhJBeFivk67CxCLDfbtVChXDdnE
UiHVnA1deLYPNyV/rbi1LnzPRqffnXtSMQrEYtmZkd72wS9InqyTymAeqWOZIurB
ziELSRsRsmrsCRkQWqvN1O7eiUJcrxu+6dX29L1sjNxXac7xUJEljxmHPNv+VRRA
wi4SXmiWs3QrjiKNl2Z4693Xl31dNLQUR6A9QSIy+FR/Ua9pk3O+FOpIaCbin63M
InaVxVPOa3aA0XghHw7afhyZaraTHrCyEbo9FMPXo2fU4+p1gucO5cFFq6XZCm+K
lU9f7eFuiqQeYnS+2CrJ2+VF+bHHRYZNlbGOQz5kz03Sj05ZTDNE4x0/2Zzy3M10
dr5panN1ww1pQPR7R98s5WQmG/f8PN3azQKp8u8wXI9VRmnEp6zNAKzxRajM2xH9
TxZ0vScR74sH3lZz91riPvcfjjFqw7eoRSXZhg5cohLPTZCEgvmrgg2Fu1dSNO4L
Qu269SBfuSbym/JIb3GzTmxH0jVtdQ492OvhYEcMuacTR6xJKLsABZPCPk0CHjlo
zFz2YY4lCR0HD9Jjsv1fH3TYXRCZbtno+hV8mN7+QyUrm5Tbz3VS7CofNq7zLJK8
4aw6H4DRt8/hd/o3MD5Ss4Ywa1cPGYASo0xXh7JyQw1PV4HWvXnp6+TeVkp4mtUw
WVM1s6qe8OF79gfYOCS50QpDrzxJPyMl0mvwakK0lIxQlFeJgot3gca1mre1DOhR
s6KcPrTSV7lkd6hbHibEqNviG1Hd4TrLMfFprYGaSNB3bO5wh7dXBv7BH44oVMtC
xe/NLBwI9EAzLMOhDofnobUFcRhbhL6JeXlmIVQnChNb026mrK/uukUgvgQtNEEG
ZxFPu9esrSS3KPyRNsIYSRlt2orFMHz4LUkujRryPTXXQA/KTy5TJVj/uO458RPK
ALhg+abkn9HTZWOcTo2nSBIOlN3Hfk5hKRz6znK+7jHl6H/ma6YqKW8N/bFjSDgy
U0RJpbjSmRaT2BmQ9U0G00j+vnLS2seWJKSTOXV3TTkRTr7sgpMg3ci80cFGgV9n
GnTqULg23/RENaVtlwo5CotjJUzwgrRWVgOr+Bn9FWBbDRaI/kti5FN7QvfcoHmi
T9rcD/troSmzzFrQ2rHxNpy/ZKKTA8LSqA0MRohFQi2Rutd1b/roqsV4+HMspIby
pHJ79tW9bb9IlUoD4APaphy5Ii0WvDMZxnmt+JYmqks/s5/1hjPwMoBGM5FYCd0V
jwCXYd+khABQ9T2wMyvKRpX4eZlidTdNXt7LuPo5hHxaW8snPpp2VBDVQQO340nW
sPZkOaf2EBY+h6FED2p/xuMkinZjW5RiFqNUB0o66AKfATMuzjR5Po0vMujyF37T
fwtRCIcDlE2ApbuAaFpAhj3xfM964HACw3eB1exmnFDtzBgor/oA0RNFibPWaeY1
NbFFdHqWkbDwuLytwM5r1YFMVWPIfjGfASgBOhgzQl+RyuSQ9GHeftw5XN10n8TZ
nn5y7Yj2tD3zwNMEe3dcOLf4bfTC1QXmwc/7PkOAbRmNpTGvmKCjrZ9fY1pc4F0q
Mxp1IyKfMntN8NDRaitpEO93Upl4GoITkWBDpUKGzN6NdwvNgzy9NOP4+F48eb6u
F5GmLLwVmBnDG36nPQeTf9goscXRYQDc4pKzsS0w6ba4uAx3jcKV90I5BHGPqRwO
4pOn79kFH53wD8jIhwUFmpKkQ+1FpFmlxyGs9NZOcoHe+8fGgzt3rf1WTRZFfEOw
Hgpj0FMu0n42Gp5ZJv4/HUL/22mzwY+v86Pit6lZ4d6kF0/byNgrBpB8Scl8eqzW
Kez6gDHeEWKUh9akwHy+S+A2QiIp1WIIGfaa9xqRnSqZ/vHHxZKb514OlkJ/cmHB
96XXu0TsfQIlyVGmbloohxH3QzUkparOUqBOIGFGzDpXlqXrAHOnHK7fnxq7mu1w
bv1bnJWJzvrVKr/zkLP8GukUo2oEp2Xd/jpuJGi1/MdUqRfoAPS9EOyJgoiAXSlu
hva0uMDdREOTWvMk7QXxSxFf1jr1rN+le8zUteTfnhDHN6uGoDuV6IpZgxqplIOL
THpLJeZjbgigrenwmzv11jyDxep8joQvSXCIQ4gPWzSFKeflDN2EQTiYgbPfoWNS
qv8JtNkiTfbm7zd4UTlYqg8naKNsVr/S3iKn4hiqmgMPTA+LkGseUAQ3ZzzqNo76
TVukZ1bMYlOovkCMCmKjIOHTwAKpQJGymjJnU6QmZv63hTSTZSU8m8Ym/uWumfkf
gYvQrED9pCf7kiyltFfN7kCXq8w4iFnKvoW9V806mWSmmQQYezYr6E3+c6wwFHx/
drLAdYhl2Q7omQ1L6LE+d+EA0LE5DeEvHgNbVr+osHrwyGTjluCO22UYCVaPJmCo
gfOqgEevBeu1y59JuCp+4nfrBcHMgYGMUZp8WZYF0LtX2R8G1x7uBkqoZY39QCc0
NC7v1JMRuzEib/qG4DxWqFkqQI4j89r0eRf3n9m3VtEHm2LTDN3HnuBE7YZR/xkq
aCqaBKLuzfjxd4IN2Aw/e8z0tQ4wWGbh69XqwdWxPorpqINH668g/KGdvOXpevPI
1gtf/YLfMNAKfgzNhbyzlHo+NCqXVIAqOOnQTqmxWI0yc/0OLEmb8246pZ8GUkqS
B9CxsdgZCzudng71Oxv6C1huow62oR9vJXeGp46yKgawbJyrm14ipC/ZDO9RPym5
OG39F8JzcuUMUfKBBEzFD+C6FcO+hj0bhUfTL9bpcyN9bGgpIngWIlrJ3eaViSuq
eM5H80pR8tMs1j7WWAzHypv9YURDa6sKZhLqJHdu5aPH4JF394sBcQkeBxTr4hcD
yxOqOd/qCXcEzqK8Vj13zWFPSaX4ghCmXPJSg3KsoOMx6ZIfq1rl+1t/U6dLxABv
23xGQLAeV146dHw1Z2CInwXRTwYHarh4uiv/Ve9hdqkhISWIZ0zPtM2+/m3A6NGq
SEfU6qGFJiBSH9lS0tWJ9k/7JCHKtk9heD/KaSY8eSwawjQl/QwTTKWPnHwVt7XM
W9yIIerIFW2StrOioDpmGfonpS09qOhSwENJX2fRbd1KwDTFO0cqj2G+En99b2X9
gwPLUIh+CNCkipQ9alFKv0LidFEU3kU3AEWdw4IVwU5aN8TxDEVvl+ESnpgpHznL
3jmFxeYNyIYhAr3PJppfTkxmd8kCTlUWzIBAqH0dE1TDYvfr/B+X1dwwU9mM+axQ
4N7lQqEzaQpCrijDse2Ldlaq6T0L/V9MAKUdzOfycyycib4QTQRkzomkwzJxJt98
8DTlemGqFAv031fAL3oCdbasUoimc4xfvzLOU74q8E5Txycxp+4jVxHMSzDBuh7f
+JRlWPf9vRjxw0ZEXDLJuTeL9PgsOaJrnoLm/c3DUJKBqVU65/bmby86tY62bnXw
mnDJ8dh4Pxb2JgSIuJDD9fpgKS7UCC6BE2J9hTGZLRD32rkymBfQM6QJv4eVfKfV
m7sChXx5qdWe6cUZxZHqd0PVX3ATh+ML5DYVCLdxHwgrkIfSZ/DjKwL5Mf3Xmqxs
lSQLveGffsmjaHFRaBUFowg6jw3KgYi8fIYwRS8PAL8YD7RJ/gndJBEiTUUv//OZ
0Gqfgt/bobhEf1EanabNvIgfBBl0Pz09LCkt50ZZq2UBomIuT57wCEFbOQn2Fqzv
OY2qYhakJhj5nirAd4sAzWLXWvj+GDLZj7OyLaRq7/5AMk0SNUT1r3yWBwv2Yqub
HYpjl4B38CyOJrz1muQr5npbn8xR4kJVRrfiZlcOLXiE9mv3odN3fgX8T1BH48tx
jJ+fqiMSJDKfqQ9P0Yj8vcZ9hxXIAau8yQsjQhsS1zuc46p22tdefBdIbOxcRISt
7wCCxQHCPDhBJfssOtDh0E+nQUYN+7hBXsfCje+8BPrMviXK5RaInfE7uz6PmBKV
jborBsvA0pbbqxp8D31/KLQDhdUSKiIUPTBzpcp+byM7eIzYztqqSatOws4QKUNU
HprYci02aPcyregjM8+J8QiyAWxWOfd/gR78rjFKvqs8QNhoPgc733dVXkmkDTKj
ZkukbIrdfa7yRxjFL+eIqAuRFgHx8bO64GwM8SERyYzON/vHTVK6ooaUwcWj9KgD
Q60X++QeMEMCk1PTjUw5AgUy2DFWbmRP3sCG2dBb6dQ32h7V3OxjVxLOf03wTnjU
G5d4wNdqk6bhMTl+bT6RNeGy+VHYYNdgqCT2Y94G/npTGZBTKNniQUERB0o02NTF
Ue0jeUarUXB3SuLMCjaumFiQ4luM//kxg39yqCRS/Klnv7P1PbRNHbEDo4hQXeGv
/CW7nrkmbLzU4pInZTiobhrRLFC5YUrKt1tnUeAvccgqU6uLPU+KkSpc48srIQAk
g251Z4IS25dC9Ir+jkDWk6IxpCHmLyujQ4+JHDNFhpOVEwFw9zeUZohfMUILJIiF
rATSH+iEtk72jxO/9q0GHmxjmSNb/DKqjMjPWRYvaraUk3x8s4Oux1SvKTWyYKBL
WMpxx3lPQZGzeo+p/NI/bbstjdYD4kNHgyqR6E6ElqfWCWDdFzCSCLm6tNEFNyzs
Jki/5UyHrRn0KvFLiOenHMJBMz3eJAnSaDeSGzKL23rmRuVZCya2cli6nsw9mi1W
up4CnEKAL8uUFTBZ5kLE8lSMeBhbf1jQNXe6vFGak/Z9LzXJOsLZ5DZyPLbVGLat
BAI0Au5b3Ydzpw6rX6YawMFC07BuaD3OZmztL8Qzq2son5louhA7hGae5/Wjdl6c
WEL4i3XgIIC/qGOdIPIZ/VEHBYrh9Ah4J38rHC9PBudz1njmgc0K/1aW16aMrMXA
gY2RToT9sO5peUuottAbGc0LITEByvBT7h8/gjUYh79XqIDrAjziGVOzkWJzBL3Q
ZvNXgX/hbzf4XT8riBhNGcovvVd0ntHF3I5RhMjATD6rmBzVqWecTOLMF3ssp0u3
9uIqJUt53Rpbjn3QjQknkgHpB9sjP7GEi61OIAvICLHTBKWlGvuGvVoqkRMYxdf8
cpi8oX8Mn9iqIBoRpFlYwruzFL6pV+g2NGAJlX37tNilfCtSp82juiQtQk3iJTtt
X1bojRZBqDw4AmaUbvnPglD8VZagfqO5YXp0niHMlvQZenqX++leV6pLzI0f3IHN
sNpIA0XNJ88+X1rgBeMuDpUjVi/MPQamG2t4l++xSwoZvfFpC2aI2ORneNXhVNE5
JKYcnrugjm6aNz6XmS3R28MDCmX+Q9CJUqct/ySbnzMfIrQQdbQWxaiXJGmiXP3I
YgPPHsi/0JYA42Sf0u7j50ZUYjO60jGtJG3UM5BdI3L19HBjAK9P+BVr9SoznGmN
4ZYCUppNREOll/mmBaOJoFnbkIhvFMuq5EPDiEeTD+qNXFmREJbz7gV8nXdA56Oj
RaNGCjzc9Ohp1yMIwsWyE9PKw9MKEuoifar9Pn2hbNardP/iPHXwAeu3M5lvDgWV
cO6I1sQIkb34TTemoONfQK3+/wNp8RNT5aTIP2Aa+XbkEbcz1xDGFUpZKrRGIVf1
TR/bHYOHH5CaN/JUE7vddRXuIvRr1RPQnL4fajHlbvPKFTve9hpmtTwqtT/9lUg4
QypF0XHjMcUGMyOErc8YJPgDSm5R/2PDA8d23X6fCveNH5KDLWTx+hM0MXhCfwwd
dp9ln48MbqvyYC7L/lOFe4KH/7yexz87hZ+uxdEuqVgVPovlo4kFYzSY5c7wfmv4
pfDDsTlv8TiqEOf1uYSREXr6YSD/XCZ65tnF88QXuyjbLjWoyY7+bmwn651xNrnm
GS/M8QfOPnMRdlzW0iZS1OF24p4949+Nl9fC8gutIBsAO47bcttVk+YmjHxTmNyc
0H7NvhjMYfYgN+ay4VKXZjcgKwpQODziMgrQPXeZwPmVbw38+AUyyFqXsh8Ktf3g
J0Mkl76wD/KQ+luhRM9hLUAiN5D+Fc07NFbaDW8YygAOId59cyOeq/ZOq4fVhfvz
tXayYoKRDOTsBv62chER8Oc8vb5Wtg7B/7YOA6EKfaiQSc3sv/pBN9ruDB5gcNEv
02kZ2baHzHodnbR5FjLwzSdgoeyjTcN5/NXV69bdzDMWKB/4QUsaKDsVqFVx3SOJ
xgNbbbI5lY+qowlzDbMRP255OxqKEvUXpBHI6AI/sAHRHR07LMxU15hJkKtAMtdw
9mgm/forA5PFj/IjvWlvnhQcaNUnnoPT/iAhTqd/UgOhjpC5gT4bb/8uUbgZIgVa
jZ7hRt9SLeRF4rzdHDdF7kuc1dLaQQXTl8ewNpwwI8hZ8Kwp6lKexfMq3vOOLHIE
mxxzUM9tpGUKo4vTYpaBWrj14/2CWko7GWGfTqx9pbb6wUsXao3fSDNuJWCMRl4f
CkENCNCG5xFJHY+dn64SYznPylYeo4cp0DVP2uZatak/Lkj/noGlpfK7xaS1RMjE
rouDzlhtEnRHwIXYd84GblUjNTGvFIKgIdNZ1iY6Q5eivi0D9y9tZktShBx5P/pW
/+2cc0GE1ex75OtnYsG5chcrLe5WHduApMwEQtyXlybun4nwhLIkzPW+Gb8BRIIn
gQSG7vty2DDMcxtUVHdR/NeJt9Axu3PgdLstMGtFflPMAuJgtX9ATzwWveipGHXU
6+XZbY+Or4MwQJeDEOnvuX/xy0PIqJm8Hicg8/+fxh6xn6UeNyRsMisFtVpsGl7B
xov5al11Di0nQI4tQtswMUTOBdqWD/lwZqtmcS+WvHG5tmYuMWWx0weCakLnXOvK
8y2fw5CmVR8AHU8VV0hZ+jV0vqynUmXKmK57yXuD4YaZ/cU/ELtSgQidNu3q69lb
2pXPNnnCuLZalzOP84Th32kjM5/neY5qN3FCYouGKkdbmVVsbjK0llczszZvtuLn
LAxC9aV4fnHg2bjhlpLwRj2xT/dq8B4rS7Z0WiST6LQgUhK5uYlf0tK05Y5yGRz5
zB23lEnwdamaDpDCDg5AzsTxG++pI/d81QeWqPAxR2uGo3rwNE8fgi6o2J5VcxeA
HLVOwNgnAa4/4aE/qf8pvoeDMqoaT2/C8QpkGMQiOx8hrZP9V3RGexsqrbEbU7qm
gwVCtO76HpU1OKhzmMuY8PpM1fntckSAwOaYJgUsrV+JTkgA063JyEaT6fGMMD/1
l6Zpy1eaDtWz85yKojHZEXMZegD9IFYsV+FesLHz9L0Ctye63FseuujSDAGk2eAy
sIERMq8RqHyUN/l0x9MOLZfSTHeHMPbZLOW/lAYd9NMNJpeOSSjwqNXbQf1yCEU7
0ougsU4bM/30xDgyGK+bdPYG72Q9Xxh4pIU/5qm4iBJUOU2Ev3jyGA/Wgzpwhtsv
14XXVbhdv/OH66gzh/iyJw6ssEOOR3ECVUZjN7iUP773IAWulDdMqSb0lp8TjcY3
xMUN4kRt6ki3Fpyms5LVR22vPkqpB8HItw6opKhFDohLmWIdcF8PmDZgcYEUl7dd
RNLtdamcqIdUYFGoAFgyXBdg60wsOFBVMJMsNnf8Z68qweY7JhG+NYiEhTI4lOiR
uWRg4WQy6ML1bIKdmC6IglJJtVTBnCQJui1iWDvSHusg8DIxkj3fFFfUihIXUWcJ
F4HoQ/UU7xijr7qskXd21QMkbVMmutLPgVz1aQ5ry2wa+gziRjts+zDN8uHr2n/D
hBSm5uX0DTb0N6lXrb30/OxEfBLStwjJjlsc8TFSMX9HgOFLObr3BQg9f9YRTt7x
WcU/pCf1G6Ewdi2he0a9705gMFMhOBynjdGXbQqCueqhSoL/lb7C3ij3mFkdaZpC
M8eoYZx55NTBggCVrIPLvk6g8Bvv4GVRkyIb9+n2Aus3fMuF7rzhLUOXOe07WkOc
q+Tn5iOb1V9MMMwRk1eglVeEb2OcGNHNYmNYMF3uFSIzK9P4NhNfXko9dnAN/YuV
Y6l08nF+ah76lS/+DMB0hw4CoFhT3XfENU4v5taKLbbYs6xY8QRlmagzJZnLP3uZ
xW58PU10CgVmy11DPZEd0GXs56h79EMbvBs1q3L+1kZviJf8Wp56CwtTyDRiG3gL
CzO8bbXSWt/HLs4krbrF9MhoKJJvFbms9Vfa6Q8OEqs0oxBITemBIycxrWB1BaUG
8BgolyBcZe2JD2tafVY+jDFce9Cooo887Aa1VB4jUYe/74ZZ//QskPuW3FzB6POH
1eHx8V8wkDVh9yoj3GMxwByFjYsevOHTOiZBjqxstTzSTsaSoAiOjru8V97HS/qQ
u7AypAGWhlz9p7uCav1+OtVBqxoaNn03Ax1kLPhQytVbZkgP0Sgrxi8ETdBA0yOL
TzMaumPd8EWxP2Iv4cX2qjq5WO450yxPQrQ5yrHGhoAv7QNNx4GR79zGYFJ5Zrbs
MTO/3KzCWtg8VgtmhT+sjiS7Zf9Nr9l5XcAxXzzI+xBTkNPklKGuB6rkiWn74Czk
NYwPHC/tKNgqfKRIAL51/iPPEVoKFMXdhGTbZKmWI+VGqcaSM3yjdhJNiPzAEp5O
by42OVMe5ryP3VGOxjp6UQPey/GvZGKBZqbVr7KtYRb/TQcPmGE+Yvcj6II1PLvL
xtr1XbrX0Ppmb+2zwvdJ7/hqEFfGgB9HsujtUtJ1dfcR5h6jn9hZs3nE1Vn7p7Yk
XtDWOlrZGSh2GbrHCCV7YnJ3NYpgLXXavEFmtK5dB9ANvw3xuT7qL0YU22G2X/FE
jP0JcxFRi6gtBSfiQa90eaG4OnBzCXQIjcVfqeEXd0b3pTaW4VNbTBUpAx5zP2q5
2z0Cw4f+ViDfhIlNbbSc6CzeRabR3oATKUf9E4jVuGHS1yyaz5rjjfq2mBZy/nR5
dEwJzGoGXtAzdPcIMG78BwOEmvhzmjAU8/xmhYADjX8+1/0DG/z+9swuDqXgyQzA
3crZTWwCo1w96cHq3cBhTTi3aL5o6Sv/CqvMp5EocJ3LhEFQ+apBuVGYZASC3bng
6ttlSRx9RWEITDN0+vWoFtk8ZvPeqsyFM2rMf8/dDbPvQg9/44Y6u62j9J90t8DQ
s8oA361tEM6JPwKD9eXUxCDa1gUoq2abqYizntSZZbf50YU+Lxsw0m2wzfHl2B9M
IwKkcv0dZS8mgaaMydEtWXofNSUOcAyvwNno9Xy7+EFPjiZ7pDsUEHhYopQxssN9
WFQmuUTH4rCaH4TWXdt9X8P1AaxQW1xsSm2Hbh9KVoNCSaAJ0gA1inLvXJK0JHC2
6NcM3WMTJucI477P/zL5ClEQrVmm01GgcmBraTQYyZPP8J6gwJH7QYnfiDUARDKK
7VbGL7VSDLrb36n8SGJvYWweudlwprga1mjdx243HxpoRxvhPNVICAmPSN44ffhZ
v2QKlr844tguf5EQNqx/Za4O1zwGJFfOS//64R9nanmjxP/EgrjNMMv5TF1d/R4Y
8YAahtbiBw1KKCwgazsnr9b6ceEKYCDg3DUTU1eeaCl7CBIL73D3flHqaZo6VtFS
CFWYJYQb7amdkzsARcr777LBEgWVtAJSnZIRHR1RoVadvpO195XRoQqLEEYaTRvj
0vUXestvuWn3Ea8e83Y0TnPSd8tmy3FGwyL7sRDXcq+WvHsVVb86U23grIWvwzZY
c0pHt7O3ycaB5IZIxYR5jLIamHesXYdUjdyAdNXf001KiD/Uv06tdULmNCGoE9Ml
6BKod/PTjZzjzBp5wo0ZjMEt+PPMdpOwHYLBxRyDXgQJnVbP6XD97F4ikfSH8kff
1/vRSG8eAWF7CkF9nuXDGk5nAZBZdcJSFVb0b/STD0yqxzzkZ5Lr9DnYzywoNug+
wmnFZcS+bQNnpqugeP2c+DxJL/9ZztF28Kn7wuYlXmQkYWrVSyYKyml9+jh6F5T+
nxPIzKejgOuhaneevW/0R9NS1wKPPVn3lbRAiGSlcsAEClN2x6VI3yG5vkjz649j
/MC/8awWR0rsGKdEsztmIDtZHvFtunxSW2UfFkRNL3SrEkN9SbH4mrEyoKmuH5R6
i4tkvD/elQ/mDrgfpQpml9Ftr19sr3R2QSMQB0K4OpC+2z5CYnlfxdl4hZvUDgNQ
EMroT/RgZ7t/QLeH6ScYJN4e06RtvR4NpREpHX2ejPbYm6V7BR3Uhy1o72oEv8Im
rexqX4zsDGyxbAvgFn9+N1NuHOasHRnhK6DTslytCBbbquNsWF5ilfQwoHu4DgOX
Oq7XZyutla2SJhGuP+iUUS/t+3CkXSMpDRwCJAGWBnZXA8s84E/7Vq0cykyIG+zu
LKT1ti4aIFLPATyPzjk3m0ykumGvl9BGEuVvXx0WtpLgfRGI+MxD1cceD8DvO0Wc
BtPek6e32CZD78GTPU6023E3l3bNXX1rHsPU4AmnCxbkrXH6IxOovJ/V0YacvzrM
Eh+JsTV7Cnnu7gWjHN/qDH10MRDb6DlR7vBlRgqyiBV2nmqgJq78vOXXesqzFVhC
inQxHWuW+7dJnmEH3ZQzGjBmE4+sdDl0hl/3iCsAiE3XwNF6VlADWY5cwdBK7TFm
bGFDybl9p/mDJbnIBZfB3THrle2kvxAdZ1ciNuDQQYMBOEFDgwCRlALmTSpjKc2i
RUWeGT14GQkD4pzaWpgWpeHw9FvUwx4idyz3zz8rPWfk0qqe92x/gWtFnHxy7a8X
CWISHCWb5jlt1R+q6G8ip75RM+oVvI4nFDNquz6beuBtrMwl4HVE4M1alt9p0HRq
i4A+Xt4sz+qQhJlQW2sJsbDuPrk4e9AwOFWhHzL37VZ8cXLP2tvfEuodhF0OzpOW
EUriYBzbtOwSpRGIvlyUY/XnSKoG9TAu9n01su7oj+ac5eQPrkirDleRfI7U/8Ic
CXUYLHFAiH7NI3KL2CYBRN+ihodZ5Gq093sGo35jS2EcQc+GzdWbkSyQY2nFIJD8
snH246Ax3BJuBqKwrBVK1ZrnW2b+YePZ2xHV6xagnkXr3ATCqXVaFq1/mBS65RrX
XXPlcf6zm+/bvCm05qDeUmrqPbX7uD7q7IPm0se7uiYck3m72G3nFlt4HjJZcML1
U6E+yuM3FcrwJo2q/gdcK8L1F1WG+9kKI6gCcDRTPvQrnTCPOPc+0v4VneJg+b7b
EzebUWlXJ6gjXtgqzfzG5tSsSfAneKC7LD7xzd2697den4Nw/1UsJwmLhirtXUgA
0J5aCJ6fvL1a77R8e5j1qgFK6BzSIwDCXiswRfwwWWoqpQVC0Cb9dH3in7D2ANmi
T7Iv6KDttn2FkMwy/JVla0G2qt170A3+1e19pTTyxPAn5wZ/O4KSlPy2JjDZXMzE
ZrWuLT02Bdoldc22pFMBh+fOgBTfwxCWuWeZAuVe6X/BtGkFyaMWIScVpfKXDTwb
Ujy8Wweh0pRHFF1BaiI0AZpELhuzc/r0TEzgNILJzg419kd63SVfTVX2s9zy2y/a
rlSW9tzz65HORoANZTW9etz+HWeiG665a0CKvnciu1oT8xAfxLwdpZan2bAaLgxc
3PFx94ptCviB0biKwuiGTc0zp8jq+zp1X736dzJiuWlUm+YdvR1DGxIMpk2v3SIz
2nXvKpkNSlCM3+JnnZQZmntlCVdAt0fvYvcG83y6etZZCRh+5e86q+Tk/aRSc+qB
ItCGRlI1LKCsBdRsuYHladdpFFSMLEDtwTo0EXQr6CrAKGPgrHIfVEejwCkiF1jl
M9dCs7x/yv9ZHzq6Zs5r73xpRvRwBAdcxg7aQKWAFLuElrjgVDabppDbO+FnJ7Pc
w80HphEnWY2fNI/vOct37byi5rqitA0w/V2TMLNEYpRIQXU58AyfpUIdqJZMl/jn
MYj05+7tvJtKZ/UX0vPQJ8ZdgHWknvHOAoMitqEaDhlVBpLDWwKxG7mEU/FpP7FF
7gvS39zDq6/S52Frwhc6CX5KLg8yAATiUKRZT67XMIg4yxe3C+dpWh9xvyHOpFSo
xqJJvd+fhJHg23YNatOd5e28Eei+ESBR20E1gwK2Ze568pQdHNB7jngvbgPyl3Qm
lh5ITqf4ikvPdC0B0kPf9RHXzhDpJeyPYHg9TrEYXWTzYzRRiHVAob/a3hBug540
/o6L+I9WZObXFinZzb/QPqgM+ycZjjiZwqwrxGH57g4KHpVuFVzJWoAVBcdnstXQ
cn4KwnB7wunnK8QGWDxz7hdNkToS6W7NC1hZz5SRkutPMcMO2ayBnVz9+fC7neIa
xVk26vwIltMj5S6/szxDo4cP6lxcJmXWbJuUH+IGe/8bVihNw1nxe31LhKStWftA
aGrBos39fgxoMw7C3uJVLPHv2814WgKKlX2lz+A6akdhkGPM5HTSAWl+1rmOGNFw
aTneT4H0uBK+NIKQalFwafhw6wACHJO2Qblfo13MoP54s5sz6eR9vSyjpmXgIDCD
qwLkSrqvGFOwFtETKgmu7Uw6Gi0LOYUKP9Sl6jgCZT8Wh4simFMB6u7QrIHR+X7P
1K/0LC0v7d7FJOuPjvhn4gyTLHbGv/KoFMf87K2kn5y/aJciszy2qUhzedAmNQo/
dWG4NzU7Og8pQSBf8yOURCjWd9oggUjVF4uHYyPKDnbFZHxs7rBOr3GGVeOAm2e2
zlra0OjkfxxXIsPcmuKMA9BQv3xHaSnUg3rB0Marfdi9Udqj/lEcb6rXw+w/GCD+
QQ9UEykrOZgOK0k3O7G2dWrw82a3gTcXwycJDQUsZYgoT3FO4L/6l/Re3aY6DKgA
9xaPTRD5I5ltIt72G8w8rKOHnSgrr8KRq707JrrIxBaZOfg77XXzgPYIUyaH1vEH
GZuaUxlJPBj/3zmqkFJlHqKAZB/Rc6MuRzGvIbGpKz2HGzh9CXkXvBZlxDgE6rDm
5dhuYb5AZDj1l5T+VTb1NG+Lh8Ms9AkAiBUA6g/gk9CbtqvbkOJDPuX3l+CpmyK5
qErpSKVC4/aOGO/PkYIL7zpPgpjW3ArCu/Fe/mZrYqbh6AR620OEDTSXEYlBvB0H
y8wENci0zBMq2mV6xcGyuarqLRbUJCas+GOaqjqnGqS9rYoSxxQMpP3Y/zcnWNfS
Bw6IfP9Tc+6hUaEQBcxjnYjSx9JmrZew546npXh8fXC62Pm+kH3GxI5ECYm6sfbP
9lUZSk3X1RsluhjtUZ4UtFdqQ6vd8+I5DUgffmVAObmd19QR4EW+EBPVFCXxOlly
YnB7OFPNXzYb3kXic2QK5YBFocS7PlZ8p8bnBSPj9P2ax8fj0LVA2QquOO6dRrGW
FMmvpNTAw5S8C6p/ASfy/jn6AqYmBtXdYgCzptZWJWRgETVfbEUPR9eztZsoB4ss
M8Kd3wYC9KS8cYOCW1G9g6XKeGEpzWigygMZGNKgjCJeT7Ozy0N4FL+399UNV/rA
P5o506xhz9vfdcSiEqnVBAPF3+89X6t7Wr7A7C830CC3A2toAHJIhoiwOql3A73A
9urvNChCBxBYnLgmwZgxlkP0J+sFcT/36foer9pAkALFLjXqHLvVvq0ETbEry+wu
0K5xu7ivvaY3CsPpic2dQiDYzWqkknxp9LYgr7mHYW/DKwUFH2qPQ6c5TjYrjX/w
N4AO/q+hZGjRMijfN7FCGuIN8+fZJT8zOQcx1oT5+SFhTv5Q07wX2aTyRlTZyhwo
QkUFo2TsugPlx7FEYuY1IYxAIFJxvRNDAAlZf326Xngp7Ya3kPrm0tyxvNvUXCAz
ANB/htSOnMfbq5f6KC5lp3YNDwTt8/BUNpJ676mPVd/hH9aYpHqw8lpbJZ/4W7Hv
7ZNxe+BP4LH6RiJ80Xa4Pt271wER31AlRClj5P3M4jucO36iOPmeh9nXNOLChVKR
Qe0a1CIDWZHOpDYQVR7kYLKBgOBlKUYFqs90f1n3CzRYiZ6dyRr+jmoW7lCVFhVT
cRx0BqHRZiuPrsMLoXQ7I94LHXI7YMfePy4MSVDfsCgSjoESjAXMzFDDTb2jhWvg
RK3i2AtAIIpp4Q4Gk553CKQyyOrLD5IO+/eoem6qq0Ns+H+YtkY8E8sD5R26ekKY
qsa0K4dFEgEwXPorG4TOU336o+lmKMM8PM12OKSN10aFKHO9xGOa+pt0OlEq+M+A
9X9WZKkCWIKqWg9r39KWih3ZTvaGW6KQsFXnG3tjeY28emmA5iyz2tFSEmtwGcqL
4FHXEPmXlsooBMe3MF0Rti2j+sqQn+6T6zDgMvR43QkCG4VUnz7zYOolDh5ocRDm
yyXMPZ5Bt8iy9MrDpbe2/fBgw2UMFT4udM2QcXeAqr0GJGIsH2+lB5CIbIcbGWBE
k7Hi4g2rCVFwAebJibNzfCBIRhi0FCZcUfb00N00nKoAopHNDyns4OK2l5PFQ8mE
oz7gK2Ghhefy6s1BZ/Zm6NH4XlSXCuSOWzF14AOKehr6Ff6ppCPTJTGGmPFDbBNL
Bh12HpkIeP6f+CWEjXYE/RGSXZ9dAFJCJtsyTTQiBBL215PrG/f/jJN3r1S6dvft
ySnoEdfgePa75ntbNt90CAvVYiZkDO0D0reZXiRpBWXDL15AN6Q//jC4JOj/3TSA
Y5Ih4MCT31+PbttttiqFBBvMUvXbB5eNSxSikrFQBFcpKniCGpWCNhikdWCHP3oC
rgAR5l1Flt+fSy8seDGDVSjNiByLjsdqwKptqFmKKpaBtFc4hQzqymokcRQ8vCO1
NfRu16xp0gka6Bpkd9wYMCimmsGdNqgsoU1iccndCsTtgh6rXJUaKgCP1wo5y2uJ
TU9JW69XnzSykC4xNzfYWx/afseK0Gti0Pt8rXtvkgsIfIurIwozgggGPWA7l+1w
usHnBsMunh8jK6EPEiDeRcH4E0B0zPllzgmx0oYE/nklyCTvLhGxkOGaiTI0jDDf
YNpGQaVPrNugIvFUvRpStX9DrCyH0TwDT4SKDMdzZQeHt29P7vystv5wL5mys+dz
YAMZdnV3J7fKjNGoU4U2w3VXetsoA5Kj5p8nFjb1N46O92nGbT9tbWPpDwr0ClSS
BA49DJnsQYQAqFYQdXuduWzLTf1x5Uj5IKBaq466Cx+3sNiImQnKeEMKrOUxlxC9
eeNAA3F5wnOu/K0+hpkjkrom7lL/H6EObKk/cVY2xjP7z5d2jnpkHxxwSQFCN7L9
AGwGffsr1cd3w87T1ib9acVR/e+XO2phN37ILfpsVx5s8Lz2GkpbaKXEmcVavpIP
hN4/N5UGRwNoa/WZ8C+MGdStWrSLx8NcnRlWl0bDielihZ7vPQmptCfmEtjYV+ON
L3RXMQGpRV01y0R1mUmRLM/jD0/skHHxIr0XcwmWcYJP8dYzgLtBX0LGVLz0CnMx
Ymzw7mbxucUgjC4qjIfS4UZlk9Wgbc64DqztYAvt7gdFDhbhCRHxo5CIPe0rEab9
Yiayev5nSWqW+i+pgtspRu408s7YaevBbVTdCemRpcO8oy/gso1k2ydAGNm+cFJ+
dHH7nisZzKuyiLxDPPzTyFgN0S69yJqb5gK3g7TIBKyByOniF5OlTKxPa1SpxPKP
hz8uVQZXGmXgE/be6+SUIffCAgMLnE4hm2Gjo6xuFLlvPD6230kDvXVp8UMUC6Tu
1IWQtBcedcJOj86F0/n64s898vmXmUrifMEC2Om2lUVeGteBrJ5xBhaPJe9VInZ+
qxultCUoiMJKeumc/7CTTmFYe8dIpTiHprskIoatzX0vcMW/l69UmBlrHyyRScrL
d+3szv1qikyt1jv7ZkpeIyTEHtEyI+KTfn/nh7RlVjQqdOU1uY0mwrvffDFgjXMz
oVjkNAbYBUjKmVHNApfZm6rTnAbJKir496+KMDZtnQcp4ffhfAYmNN6DyvMi3SK7
gOCE/GKO2Ls18ba1uIpakaVMRhrXBasyh6l1HieiTR8vWPFhl3pDfgZspV4ekTik
mL/VEW3LqDdXCOmA9myIeAdQIZCdS2MtSXm/QwcT1MRnSb5Ggn9TontKjJaVbPyw
ejBTaN1rZqHYAlCgpETSkgOdmA3VxJuRXfkdPGNd9mvmTKnSrXpZ6MTUDO16CwyC
JAG6gvv+Xv9cNKVa5dGGLHOaPMbQvsFV1V/uKFFMdMq180B9K6GKkUxlpQtsz08d
/A8aYhGCzxe9WpUi5Xhk/ZJ4pigQvU6YiKqSeASv2L5SY1e1E2YbYx8Qz/yK0CTc
Lvitc8lU8dioAHAqnLpk6YbSFtT8WOqH46Kcik2wsdljnIFCY1uqUUFahcFXV20x
N29kRYy2GIYrJXeiQ3t+LtO1MMtXE72auddSRFygw7FMu5xywu6aZboEgA2Lq6um
NgJBPmW9ZoPn3Lf7EgYHEy0rwjHfEmCh/O8mlPkDUoIy97bh+o1bFyZiUoxInZnk
3Utejyek+VzGW0PrpQsIiqxBWMuPGzEIBJasMUbzHpYFFrOPQct1Wl/P6SETXTNl
MAmz1cz/7t2mN90kBgo37zBtlVMOaeMUBQeFj3CMAYT+WCSP+5IeyCw/luMjAv2O
dcuY/4Kok3JX37GJCNLWRZWqjPwbXGMZs37DcDY5JWIcBFVET5kKxd3LKNpbHYTC
YYeRQI0hVlwOxXYN8bsiY9GxJRdc/63gF0AhhWKB9hemKLWp/22fTsgwGfM6vg6P
leVyjJkUKC//fDiis9tRWdMP3nTYBxNJlnbW5wIBkOB1HgvkIiLsA0ahMuZPQpz5
Y5tFdkyyW/1uq96K21g/tGpywe2oiCtq562mEMzh1fucFu/ZFYdFT3hPvBo55EGf
xQKqEzfBFBrbxBsPAB5B1+cNzBz9XwdiWppb1gtu9eTelWojOUAxxq1e99dA6ffZ
j/EhevERkChGdws1Qer8lRggMpMpuYF0vHWajH3z5cwYlosXN8sYwPWiIyjtdJgT
pf+gTZgYASi9cZVJnpmyRusBcF6G66lnLUnKhLpnHm9ZRMXsk9ERtC1TxsJyn15H
nBNYIZi5mEAfUVZxfRHySGm8I6imkHruZQrG4F0kDqqsSuPIPyZqPsTR9EVlfM03
Il1L+DMXisTcYP5VJ0r68ARKnf+Bjj9S1kY9lYPG3WOAs22EQuL5uhTRTQ2nU0Ke
aQQhLokdfLwbORsPaHxiGdtM4J0JrEWhF8oAB53UxbyFzHWxG9U9ZhPuHWEIQgLY
mnuF5HuiQ/r19ikrD0Xhl6n2wbWWIbjgUlyG/oS9tWdESQjhQTMxgNyIDc5ngD26
Os5ZYCXtN9LkjjchFwJVVaMdWga66ZGhoCs73b4CjNpUeXikZHCp5PmbbUZg/XWA
OCKD35ODlzFmUlcHu+euonBPj24NxZUOgkhXJZyweBf2Roji408uuj5HjGv+wlGy
ZgdI+k59t+qYYWvDQbuJnyez3DM52AQ5dDhFo8srHeeCHqnPFK5j5hfkS962mNjN
EP59JscGVYAaRMUqKEMP1I8J2dYCTQ+U37CIfNodaL93/8cIsnsA7HWKLqKrvLsQ
JGEYQunKZr5hYdxpF0ks+VWi8f0lp2/2pn7rbqQkMiNTOIqmGPkeI/5KBop95Elg
22wyP990p/0TPX97fmZjRwpcEDAkjb/dUJ+WLms3H+RoMtKecov698bD1xEdx52g
6ORetpy/Qkx6xI7O/fCQJOc3jMKKE13k6EsaSr2D1a9fBmHAklSzmdf9izP0jcZE
6I63OrtR6NmfFUhd6OOLSPdV5q4JxVgwv/Msl1Yz9XHC12j/UskkWc3q4juc1BrW
a8gdyq9Ct50QShdacIukeZNdhaM8OjMygTCifJlJFESKe8rDVVwk7iTp/UdQvzBx
XCHPPZjXQ/u7YFebrkdig2taGCJN14jwj2CtRFSAq6m4mydSEdl+Yy6Ax0EFA0UN
D1sNJdmBkSFgWKga+1l/oXyNnMG1uEwwSHIUIoYfzz2R4HAGr3mD7z1Dhc7Fi+zf
r2uzNG+5zRdIF2mRLmv6/mSZI/2Uclf1uvn7w9ws8bDJQOXjnTa/910z+oLXdvl1
H9RlCD7RdwQuliTkFy7n2F0Zt1DBFOr6vPn1mB17gUs+U2T0oKgigKJ52BWJBfi6
guQPBsreONXCPE4TJtcn1BpsmOWte5SfLo5y17GoDRvbdXADk+52t+pmjTL3gtQm
ZyeXPdU778SDJ7Crln39DJ2sJcKxC4C/qiCFIzZAtN+IWzE3fB2WQ8CTqG/pd/cH
WwRLHwny28LCaeyrc1nJ+6eOngjoe/a/Qr5D7oozjr8hcQN3n7qDknV7QDlTb2Jd
ZMaHjRAeOOf0c3PPPanT3o0NyXL0GnGr0la0z7qfGv2VirmrdqTBRcZy1iItNJG+
Pi0vTPZuaeFadHWmDtwuwl2MmTrW3OJIxPobFXlfKdsb26NebaxMNK7v67wyilZO
eoGd7kuawka5AZMUm51WY9adufKShr8lURfLHW5yCEqYUk6MsqiVDXs2U5FhhN5s
yKXXpFH/NJ2sj9OO0qcdpSiBb9GOCGMyL9tVNLOw2mDkO8azXNoTTCgiob/xAQoA
yEkOnogp1R8Q51RaeiPLfbwD1Vof9qj+3PPMKRD0+pUDc7nKCLSvwSKUgE55QiAP
wxJXcOPzk3IDy6uGmrOEbrc3BT9IBO8pRA/s3fGyel966aLv8Er7dxCDn8U+C6Mf
s4P5Hvf2WP075gF/QIUneYgDt/oNlfYhUcog1l7+PxcQm/k26cY/OygZwD2SuwJO
ApkAAIIRouO2VxdK/iJMaaJHCdf3nEq4k/ZnpjoC5FwjypyNt9IKI4WtyjpG3noP
bi7hYmn6nqdGRfevelRiBQdLXbb5rwbKxTWYNNBzWlLfhsUFpAL29bmxu8hJVo/t
Zg4VCRRQDHu+A3oklloJ2MzGAbEfcIMRqZYTsCzefxPeY3TI3f7358EGJHyccnbH
DrpZL/eqlAxoolhL/Y3L+TUoDiZ47pxIyoiqozT9SUh/Lzr9DxC5Cpp5d/PM4WEn
vEN/5FKvfSfGZ/0v+4OSzImQ5ece7txwqjkcqgITLOPqqwB+VRu8xKoUqc4JZE6E
Rs0A2SkqXgUPE8OTZA6DvpvNruv/+AaWq6+Sw/26TpXxCqRVV52hpUK3JtFiJD2J
dDsGCw2AqmN5Z4Rts8+5he5kAiGiIk7WUACr76XcROxIMcQ8YC6XQ7SFAjwNwklu
4b1RM+AzhQn8OQqDJ+PX3UExsDs6nKrZVypcn+cUUN6jurno4gzLeySbR2gKclO6
vclVOAoE1BW+mBEOwN/fI8A8yYLuu+1JVf9U2rhb/Xs7170AB6fMC46r9mCouDK/
9OQ2huEnPZjsOKCw5cTQ/Ex+IJcRiLuS7jnILwr0lpMQqU9lo6ihdsYr/sYqhUQA
odHdLoqcf7ZYJmkPB+y/5qaM/wZP5L2j7q0khNZIumXdamhS9faRZCufmoGCXGCs
scZr6yXc9rRyATyQupRzty04VaPdo2hn1IzSX211tAKcio+jmmEDN0X58PBmO7yA
UQV2CA8Db5LBzWipfxgLTX1roslKl6KKkE4b9+x7gtkuCtlt5d6Tw9GjZgYHS1aW
BJZGgZ6yQi5ztVP0eNrvdJbEMJaEPhcBkjmmX6hrY1McY///sJHxVWh5zBemP+bK
1KUyIkfFUy5WQIDFBjTdxHupjEv6JX7DskRjMdokhgSm0LuduO7fHLG/jhnvKiLJ
fqy4HAa19leV+ZLZ5o10REbLtVGgK1oRDQxJ5ihwKuHRNigDsNVurvBlBGlFs5zp
UxvyEq1O0CrzHfz4O/0jt/eZ9N+GS9PE/eEeNEWNe/MGdCvVOwcKddX3f4JLUEFh
T17bwIyKdNKTX0J8WRndqdKEaLsqwz9Q7G6/Ues/L3T6uI6oaE+ecpMmhtbSwl8F
rYogS206ZILryj7QIsWrV+Wf1P/Mlu/DBTshFnXQ7D+DxBxZXbMJFyaFhz+GL2Wh
j8jX+GMcDnXYMml2CFffcVPLrP8PkvD3b9wTEsZrJG0RuRvqoCdQz6UPg/IE8gaY
CnR+sKOa7Bm/Ej2O9VRvWE8dwbSQnhsGd/gwc6Bjk0VNqtJE/SymRUvqNK0FgzZ5
o/4Unh2K1RMEEF7DeaXY3dyPvJmWTRI3gjSFmRFMEpjVJ7rtdcUWQ3a3ujCvUoxj
Cq8DpDwH9EBK088rsAMYaVsbNNDlj94yXlJcEm5wvpIDiuH6m49f7Q5GsE5WZ0Sa
B4p8e02TqkC7yxnRH8H5Ag+nHohpdaW5cYTNKUQySltLKrZ+olslnq3YCF1LDXXM
T6lBC+YEw0da1qtMbucpaFDF3zKsMShUJLepLc/3o1xNweeud2Qyx5oVlQgdAbEH
/dGdI65Cdyflx0pjEzcJMaaXg+3chRZPzZz/otyE1pS6gTJ1i7XhI6Tt2s7pBBec
kLZ6yRniMcxXkj5SLb+JtgGhARMdgoHXY/6H/er2doreat2rCBvbGKC5WCX09AbZ
SIHl4wkjsqrFtBva38s7r1t2juqcFd9otWLBO02QKXWZiNjZiRoryHPOdC1ZbLl2
M4MwDijoaGGyBMObqHNTmD8P7laCwIOMfXAaCBjv7Lpzcypa5D4Rtqj3kZ2KIxTu
+qD/snZ3HPLp4MN9wQlm3T5yloeK5kh+qn7t00DrdD5vk5ZmOTD7G7ohi1ErGMW1
XTrl7NWDITAq1xV/MVeZG5rsfeXfLZtgybICqs4IBQNiLEubHvNE1rNT9kW+bM8G
xdakwPS8t7JkZ9Fe+QZji2I+rxtTSNlDC75dTmhnd+iV3euD7MiYectIbu94saTT
ohSI7TBI3/Lh3d0FCiKGwrWzNNXHumaLjyUx4rQJVsa5Pxbpw9U2c5kvYMLnDmpu
WP5USgNYtOfcu1q4XWKy+y0Nd0b3cF9yX2pAjaYUv1LOyFgV2/1KjHspC1VJ8twQ
86sTQ2f7e94CNmwqsmKh2Cdl+UW8zTsN9RL+us0nCTiOYG3i3lP8kGJi2MrmSU7T
/1HYixCBCfhJOKNH9DlrT1SKeJmTG35rmYtcRGwTcYuI0FT2u2X5hx9t1Z5hEHoc
0iwexM+lOUiwpDZLKWlkAGGy+E5Auv7JQoAsotBfvW0ltd9rGX0n/5a/WvOaIR3d
hUZ8XDa0677SrKrFoCQtYNp5TaQlBMeMZC3sPPxgFMQGfueyEYWRCbQVclx3Qa6y
cFeRw8K3ESA/e7NFregv51LwtkJRbTepWNacAAhXaoXxMqSlFtxzRIScy/pm3+rA
MSisSySpHz5SL598D5TSc+pBtnv+nycjUZHp9qeYS5j4m4glIWDuYl6e05vMc7OS
rRUSf0bly3C1eWXyZIddPPD7tMLpw19OAxuslI32tGYo26IptHG0wKLJ4C3AOfmN
lpLWlAfFs+zE3DS+rU1iThdERW7kVcz4aEPMNg35FhE9Dn1TITIn6pw/r0tvtYfZ
sgVFmqUjmXbsXeqo54itdqJ5bNi84GzXFI/kNFJ96s9jc86W5S31S5moqzhdbkvF
X62iuG6OuOUVVEn/w5cyIL3x6TambPCSwFdcsbYcgnBeC3qV3O0twb5H16FPv7QN
MS867D5buIJ7o1f3P5rhkiA2IUGvJ1SzgjBzlchS8IuIMH6oKSC9upzUTVgWRA4e
5D6ETs6hb7mkWfsrwXyjdxbxY7I+7oJu4reIhxZ1MRMZnBR9omHeRaLDtkWlZhUf
iZNLPQfL/Ebwo20k87EyXwowKwK48EO2pYgZyJszdJ9nedSfBUm9nr7pw8AOA1O2
r81jHSkfn3bLIm7YalcOU2Tui/iZFEmZIct9/X044o1/bTP9p1lf9cy0c3Z17czN
dkXCnKmaHHDAirhmiHSfw1ZMj6TBOntYy2oK2KpsLP1nJc7lhGZWZyrZP1YKY5y4
Amjr+fT+2hYUBYPRqah9hkBjXT7PZyKFZjOclznNb5gJ864Fuy1m0HtvYILShUma
3dH5yPtyfx8runD+wZ9ZF0iX+sRyQwKRiSzXQSHVnMYw6Yej4S69W/hkqSPLF4g4
Ex93BAcpIYEf4milHEGsd6UUpo/hPLwKj4glsGcoDcAakWJs6rq97YmU5BwsEj9V
5A94wnVYfvLITx97ZxCFZ+M2uUnLnC3dzycW0mh7MwG2AA49sk57P6xBGt3qollB
EShzO8bRnhNNLwDpR2gvrPEskX5+KVuAarg7OnraeS2GoaDJ6IbzxOSolw3qtn58
MeHx3dTJ9DHMkTZs2pjjdtbPMkMgODXJH3hHi6KnPvU/mLayfahO2AsgwUjO7edM
Afj7HB8CNlZKHhF8AGYalnkxC8v3njfkXfFOPllpONnDScYjy7VSm9O7vPR8bFmh
i9v6PGWyVQxsmsEBPEgJ15tqf/c4430CVzJr2KMMeZaNQSOhbSMuVpQ/doGGnV4o
u/j6+KBWP2SCs6fWxFjU09E6aSxHewRibOfTW6zYbQztAXFvI2OKVRyay/a36W5o
jDHOE5AhuNhb6UPlSnwdBAPI7mOIN9LUDX5GaYjY6Xf8+mh8oyAAthwllo5QtV2e
VfqyRxcog7/CyhB4XrPGWPRdY6hJDDCUEUSWw+DjN74pcN4HLcL+mfeAh5CFml5r
KvsCl5BJKKwsjG2KJDIEzkyv+LPDnLOwXV0ecA5c3NGkmvNTNaNAWkD9JLpIFSDC
w4OiZHsMzH3TQTo6OpoyqkA/A6iRN3LIz6RiNWDKzcMK/kb5YEZYQ/HGtXxfc3bO
IVLyoH+F+rpVv6NjyaqU2yg2C8ZBgParEI6pBj8w6w8szHBk2os0n16fdSWz0YCi
pKtHLUi5hBvrZfIPlGOvgz1bagJhEo8hoyNeGrLBbhgs+hzPdQpi52evzHSEAibc
NRGG0JgCeMyKLighcG6FdxTIsQ0kIseQBZhZzZK24QHAfEkKNeVasVk14nLANR+y
7bBAwDzcxE8kXnzYsqkJRXRb3SjrJWNFaQzxChF0oPe9fI9LZkFncItyJnuTE9Gh
LBpRkuOCe538lHWHiYGf+S2djz5ybe5piXYoFdSRf7EM/VX4ZADyC+A3ZGfLODgO
YkOCO4/PbXe8VFm9EaDqTMkv4CeX0VJWNkQuYjXBJbBlI/oZmVhQhY4npiOTIe/C
TkLdThbXaU1oKkGBeBwbW5HROUjfB9QH3DZmbZpEKXObK/1ebSYPFDk90xH1RLWl
Po2kJY4HEEef8QZ/g6x2vRQZmonUgcQBCpVSNfHzlcv03a+M8O61+0WxFb6KdqnG
VCn6v9PAgPOhQiTOYTw3jCkUINUnDyVgs+Z3aw0V32AuB2Pdm/RmkaGCA+R3a1lE
a13V+QX1gozztxV72FUyZH3A2tdnpJI0IZ0qw1CmcO675g8Ls31MBHkMgmzY1ZJ7
myrtLmeCRZZNMfoOpgvfPAMcQhiEzI3sMeZTspCipNQxbMYyIKAasEHnBKstkHA5
W7gQiBYD3kXlmfHTTT8oq+DeSVdN4nzVcVOmucLcFwfZ2J0sbf3zlvwGRw2BdGIh
Rhwx2So17tUjZAMBOaVXPSwkzHhslRJuq7dwXIGirH/QSqPy9O9ANq8gMWwQnUBW
Dty9UCGE8IyWXC+qzh+JyYsAB66gVr+omN3RPu7739DhdWppeeYMVcflPIiOaQC8
uq2XX+Nyff7kKz6zrDfYGoRcUP54R9nqvX+fS/bI6eeGg82qh3tB0OgJNCOov5ya
fp9DMGE0Lnn71sVcnQL0dpAgYDBqkFj5RuIsaYtzB3jKp+xMwzbOzOwlBrOqKTPt
dT/mAiUYM8HFx4CKK1TA3xM2nemLDmGyytyPRBYfTGR7JIYh9IsZKw33plBQ3zEK
r8j+DE2I064ojQklNKlscv2EPII3m+jjjKsMOVRpHzHApGv6UgqTaAATWO4ChieO
6vo6UslVwnzZ+9HbCRSI3NudRsjLeHptmj/ULBkC86W4wmSBe2OjHPNmY5UAbxMQ
RLfmPGzMc98kOtbNMRG0OzgHncqRgxcQpUYhoB+f0s3voMVVAXlHr76jc+kdWuQL
jqbQWm18UdL+sAY7GrgcsYtVltcOMHjB193Ntm/cUot5Ils1zNuzshlC+WZ8CvdO
BWBtzo2g3P9CUEi7qUFav/X7NxuqebFhMOjAR5lTOsej1L3br+v+cnMN111mgQJQ
gdvubF3n8nKGzkESRDHSWLcWE4p3HHNCaug2yvVCj9RGTE/yZSrZum7YY0svvXnS
k4Wmn+MXbHZYzqguerc5RhK30QdhCf3vRgrxc0w5snTc1YjeP0ZrTB0ui75xZlzZ
sVj+cUVpwbpTz5UrAP+98VM8rHgz848iAnwhc+Nu/Wvm+WjMZTDj80HMqkt8z136
GsC9v+3ouGb9i8cGD0Eb2MjHebEdlfkLZ1Q8yx/U4uDLkpqLdsKhVIoxqeNltHYF
oV5x5wAFlrmD+9vceAvsWg+NhOQdv4BsoB8cZOT1Wov1JUbH97dUcS7/aMCJwau5
UzkzDWAUU+p/PfoV8Z1mBb1jv1tRMf3zkD7nqGtBbg8TIgHagx4zbARRDGh16juy
qK9bqGHspHA4JNKMSUD3Wvxfyj+WLcZLMWwya0/mTQCwlTHCNiZpSb3RhsuwtfFX
lA9faKpY9tH9qyvt2a0nChPO4xiPw5MWcXHIyhH51LwcZZYOyagCv8XozaF7atLB
WGpAaYn4ekEiih338U5oMpkRfKyrb7MtY+MsWt68VIH/LodeResBmf5255MV8nsc
6G3HMD4EIGeT4+aLphcgOBV4lQ7cZ/eT+iaOeyQPlGkYiK1164FkO+RxmKXs9k21
wWovGSUdUqD3W34tUcUtj0SC+GhM6iTm4rGJwkYuMqVVWIOgIVUdEE2c5vpDSvnJ
Q4i2dUbl/Zg6xxmq8SWjbYO/Aki9HDEuy+0vIHrdeV+PGIMwlWaosCl3OoIB4Jrs
cl+hWz4NfpTFFGwHh2BesAZl+meTOrSQ6mgQkczk+EffOLYw6+AktusG69TGR9bX
Ad/4B4gTysIV9k0N2/UngzvUOXOaOp9yovSR/N9ODQHpfMfw6tBTrQaLBfW94VTm
Km7ol/OGtmgZQMBUi3GxOkv3d5BFObAelsSqyitmCt1Cn2+N50PX4s0IZc33L5zf
L/r2UKnMLMOCzrSigfWSvYSIxaH1oQ7dC06rpj84svyY8KxhcjUYkzTqtrZMj2Qc
EZbND+vwod9BnPZfIG8mxjeXtbEUOqxLFUzC3chMVfGvBncQemgPFkpj+fBxrkJ6
YQKofP1rNzecHGzzunyEJ4BvbnLZgJ0xdlyzwI/0CoAdF90ic8Wm9JsbxWtCEmAQ
1CEPrYaZjQbGhHwsWti/NI5dYe6ZN5dDnEzkwfERT2+7UvXwuQhAMkuC9fwkCvsZ
6tQ/plEDU7Oayx0k3vWP2hMOdCELJnTNmgSvV+rDCCYK6EH7Pwf6ctCUsWsH0XcQ
0wDHvy0Vf1d/vzLnOwsVs2bcefNBElKlvvft6P3yQkc70ARzRfV/7PzJ98jnaoMK
G33Bnqov9BB78rCPiq5jxuBuHo8x0vrz6uP4IbaWc0jQgnN4jdkh2v6j/JFHlszD
qCojXwiMewobIKjZLbjOtyDKjRDxmYUtQVRRKBISoxZxJ/2tJVUanGl6Uo/t7/bB
pe7TNUJMo1Cdl81SqlmFLddhYec+PgQ+uZ5af86pln1FqwFCCeKFxk4bA3NJrsnI
sbq+FuodrwQOUEqh87eiuuWUIpPo/YqHVyZ2BcFR0RKKtGFL7ubhLuGhNQelH+Dn
BZCUTTd5FDBad2i4PP9W793FTJtSmbMZ+JJArwfshJFSSxsv5pP8rye1hH7k5ezW
Mnkm5l4dDf5iB7OdA2KELBhjNHzb9qvLR29WoVPxfHzLlO1XEh81Gs6NqTVtm6We
IkyF2P3kkRNb9kz2Zyp/vvrvdGvFth5IgcFQ9KQ2y3gD91l/6tMW4qzffeg1AWRu
hIjwjzNkhnybAeJT9+fhGQRJ/YEaGpmu4K2fFSPGPNDVnBOhGfWoJD7kBKhlePaI
ByuZB2CDSggWSqkMpgv23eVxgGIVPOdSKcefe4920wx+0GczwkRh/c+FZ32ENQXE
edS5jQrHWms1XM7GqXz6KJEb+QPX3/H0BFqt2goLyeA3bDhg9C6x8J/G34+SrKwS
5pQ9FQaDLe6nMQ2YZR//nTwTLZfZ8Wcx3ARQJXk7NI3whn20txZqo8q8pS7bpvtt
Lb7Scb/a7Ne8xBoMstX0SaBoWSG7pL7eBPLYVuEc8ReEe3Sk6tFAM0DqtpHG6K1c
sNGZfclZYfBUexT8dch8v9d7qQBR+27c+c0n6WdkJVom84rn5+hp5HnKAlPdQVK/
DXpsUfYMaoElCRkLujhDHHBh9d8YBzgs5AXtRlUIJlCOX3ooEupYZk4q8bsNF1v6
n+DRuM9Sv78rvLHKSYus4aaRp/PG+e1z0FpUZkKNGdskF0fwjcuR2jlqNhdCl961
/DlXyyJwN1LsRlmhIFwgGQI/Kw+Cbe0jiInYVKIl9DaEinrvToPYH4zK60TqUgyC
ZB9bEPsD6FIYPksdc184nNC1/ooi07DxkaFJy+gpnNnSSW9Eq770K6VYXpAkrjSu
jFVc27Kfv8cYuoIUH7WrXID/ADP+WrQnfOgwLAzFvigH6eepnbSf1GBX8+ZXC5Ps
cNGDTvM6k25N0jFB7iHmh0wKi5kcCHzmRojQ3ndY7FwxOeNp5COkJ/2+llTP8JC9
zz106HmD+f9K5UNQa/G710jEi1RloZ0xhxN9plvpW4Edv2BFIQ6QpTOxXjXakVAA
BPGSrhfTYD3fFLBQE1WPmabuAQDnsWeknjwIctlTRHsm94toGAACYDO8kAG5wvBJ
Ikyn4HLDJa1qoIDwdcWYX1YsNHPZnhtMV457/VE+1+zmn6o83g2vpHJwWD6QTQWc
1d+gcQBVRz4rYUqtXGK4/0bAszk/aKRBILVIxe7zXXaInrTLT2FSUZ8MZf4xznz8
swZPD4vNuN5GdAMwG8auxvTtNi5VyvmJdK37vAecg8HgFFMx+/f+McGjQJC3cRWo
6TOkTHCCRPYToaHznHydJC6N8CsGRQ59owTQTeShZ5W13ofiHGg9yiQ9LHclfgHg
4SvzgGihpeUwFCnfKGd9o6xfGSAE2kAnlfvDuGCpKZcRj23YqaIYJ8t0J47dI12K
eFbVWbOSPLsnB9GQnnmeRJHvQFqpKP2FHDMu6WYBiHC3Ls+6JzMhfR7AandVUtrL
WmnaDfw91gRtpNaQXkuMphIqor2VwhHreTjb9dIWH+FtJ2joBNOEKMJUoeAwZ7JM
4/rTOQZ9GqUbUoOMTJKUet5kxyqzZp4ztO2s66YL2lOvC0aEWh30OQtwgt7btJo3
0OgPCIEbB/eodLhDJ6+S9vlB6isMQ1nh9ZewR/rr7uKv5dfvbM3vs2VMfDrz/v6V
aXTrQ46j6z4QMxecC6WOVJISPuYrkxsXnS1XLZsDQHdMmvmhS231us7xWjRsVEiC
wo9VmcA4aOrV8b4j+gyndcJU3KQXDWjKClmGKtVlSQwbg8K3fqPdcYsAolbrc1lx
uWXKP96apnO297nlG/LJRjR07MhcOOKeFE3kEBmYHAOhXDWHn318Ej4eAb+WRyfg
H4TXdNrLTVTLEqm5CcIIvCWQO8AuJNlddQIFGqnWunBAucl49xU7fdtYdnq7gGFA
MCnJkazkpOnKeqtssTVTHtnlUaotqAIl3hg/H75y8NmlfezPperyGF/vF2r2hE/M
jIV5I63hWNiKRNb6skiqhOuCqYuhIUDa2rrecCpfW9PfH6hyngnVzUFsxUOj2ogY
87yQC1sd2e9kaBI5+viaTzuzWD2G+elgpM1gf7ixGD9m0ckF40/qYAQVpdzdBr2f
bEqipqdGAttYAZJJBwmh3zWJVQHhNM3vftKdHdZuUTauORkSgWbjs9LQ/1U3/koE
dpEy8EFTHLJ53PdGAS5v7Y4luKMhLX+qmkNPX0TM49MI5XDT23K4vOs/FRBTin16
icJvJiVEtreQt9YWG1AWppsDmA5D0dAqB6Uo8POXXBovl+C+cSU6AAZN45CX5RdO
DqrrWdriOkbnUxmtcMfZ1Ghx26WDod+UdJSbAnv4Q4m5qp4mz0CsGWO778PShy7P
wZDBehxS2upnm+vTt1rhmB7f3AkmpmO0SxD0A2yijF37AVYkll73FVE7DJTU9VQz
s9l0fm9pyOFgd94Z2dyJ/zM3FAkcbG9Btr2HzyHUr38mtGgb7gGjI+RT0RbsXaqx
L+OxkdX6C3JCaTRjFzZ4jc8t2lvHF45kGLMYGpMJ3xYIBAcLVkXX0LBghzAmE02B
FSbCryHVAipfNLvusZNvDxb0Bp5zXYiovxttbeiKT2jFHsCD1qr6JVU4I1n/5kmq
yOBhYr/RcWoJDJN4YGFuRaoICl2QA3woZZeOGtPZh47ShL3yLYOrjVvX6besrx10
Rk265nd9Gc+dQKcQdVezj9fzTKBB9k79KiuTr1xwXKd82xmzKrl8hRNeW9eOP58c
64HwABhxOtoOj5ZoVlOL53EDNJRmkcde7Sl0Q+zrs8tLMvya07k7r6UNqTObQhjH
zshOhsc5etX0V+zTQSJNiwWc58wULC5mKPXhJyJxVODpDFf+0MCCrGszR1uh1hMC
Y5QQfGqPL/RDtTYFOGggQ8DOYIhnWAPBS7L2H22olfwJBshKKjQ7ekIqZ12fJkkR
EqJp+g3RdYKI33U/UcwGr7FNAiX/Ip9aO0CP6VxpzoWgsQ4TL3cOEpV6dR0Ly3Gx
YSMcbsSV1NNgPUd1zeSXvMuH4QWrOzQE8lWrcr5qbmBopaViM2eaEmJSHrXe+hSB
0Zb1SuCvWo788qo6kQ+9yeqgA8c/9H3d9xvfbYLjlszpQWddYxeklVqTjlcL5TCE
9mk3/A7+6MQfcKPhjZhPt3GujIQiOVBgGcsxB0PEVpBObXfu2tAhVmo0SZFawl5k
PFRFPFyUMwStcPPh9zq15pqCSa9uUKLt4vQyoa/FYJ56LfTqjy4uvOmX/REex8wL
Jk/N8SxQMGPuR5Vz0UuwQOA+TJczG5LB1JqvcM46fMW+BgXmvfvzmE6PyGfFjPJz
5mKWruqhhrx7M8Xoh9Xulpm2ZSeF8r2aRCXmL+xLAkf6/W2mprIIekFX0B53+WMk
R1xKU+xzjlFUKJ0XCyHzeaHC/nMI1s1MxVTMLptyDW0othpyVeRHGdb+7C79Ybsx
xcB7cfgbaE6yiCEfLFyxRIlGQUCPUi6Hij3OsqP/vCmW5XiQBeYYi5caket3VK+y
K0Wt5xR4kMD2y0RHNZUubqGj1U6zGhtV6L7ni6Gjja6plQC3Z9H9PvdPfD0jn9wi
PtyicCSjijO1k3jtgMdscNBU5i1v9X4oTz+/P50b7FrVRPxjyYfTG7ZWVKiV+vED
TrXn5MIveqIQjdZtSnTAYyn3ov/itJt+IT8GywoZLaqjFLwnn4x8hhIW3fu6BC+S
bMTKh/7O/87OiDBynQYdIpUjRZCje6NimN5jsM2ByqisTGvMDVEngoRgiI2aWfkb
2iZGDHYi7ECl6IVnMM7xbSX9fGBmRCstuDNZ5l7JvvDGw46mlNb5l/oEJhmw5h7p
fqn/x08FjHmK0Wu8cmSYDNyyZxDn+JBD9mdbFLuOGYmJXqqE9tlub8fuysZQy4HA
NTejcL2bK297ykt5DibN0CIX/h6g9ZeOxjlkGzPfoCdbdsW2+9wnvzDdVFgEj8W2
OmO3x+EojyQBfbH8L8TufRGoIDWnUWUQ+IhBOSHK+N+j2ubuoJMJrkILWE3DcpZ6
Hn4nIYERnWrIe4wtB0zlfSCsy4QYx6cNhR0tmw3qRqhy6hADNEn+zU3Dd4hN08b4
qHceI04GnD07fLSisWqkn5ya2xmVj4uc6jeATlgw3V5k8rQSFVPaNaZGKFCq2n4u
AeucDu4M7KFZ5LOxS02OXvrMJxBQbkVfLHPjzlBdHBB2UP5w0ifVxO5Vy5jU30HG
ZFWqMGXgXBdz1KjqATGUVQzmXJembst/EWYhcdFZqExe6J+cloMQiGXeCcRjqdEg
AJO8IkN0xRn/M9dBKkbU8sx4wY+KdXEciF0wkw96NDNEY4DDik4WI4E5wsmR9YWj
0iWMru8Zj9hPn0Id3J5yKbX2Ypkjr/6MEo7b0L8zuCa3W5f9Bd7XjK6qJHhEqu1E
h26HiNVHuevehWU/NSQ2maaD6nVj7diIqZNL7TmGgpItsbglPeFcfxWRyydz4WV0
DBsYus9It9GBYLrCfRA5dPLPfgYA9fFe3h8Ec/+nCOqhSf4Z+hOh1bSN0u16fMk7
R7CIVLFhvTTHG4IZHSUu3bBqQM40BTbie4qKVLyuYVkZpmLwkwBZ6U6aCFIK+uAl
wx22AjZSP7PYOlnuPgmGGopvJ6bC70aexmBG7A/YLAtI6N5W9/KgcuMcloULKpOb
t6PhCpebMt4LuoAMtmtBX6pk+S+ycNLOXCaZCuTt7JZmY2s92nK+YS2brDS8YzNj
6WPvR2cFuf0j3uKS78MI8qH+8SseukLi1e3VXMvQX6MjYQbud4bXsfBoZhKdfw7e
W3+BED8Ze16u1w1I0/OTCT9VhKpNEBFKFw29xQtGm8HDc1tuuOGW0RUPCyodLvXY
tVZTssxsCzxrTsNg0Ypo+D1xzJEsD6aeD4OS7gHOl03RBeCZa8XeORYQn5YBfM+j
Yy203hocMFOo3ziibA8059m0YrUUukOLI64kLMsuGE/6h4eCgW574gsI42arFXXF
MR+fASE3w5BG8rCdWs23S8jGqPvAuweWDoM63uOpn3QC1nR0FmrOwREEM35zgddG
rVhVtpIv6Vw85HBCT05Tcg6Ycxb2N6Ugw4Swdgiimuhh2ha9pEMtv9NU5WxDgUGk
DT8X4CXQnLPBwNn2aDXANqhRQd+ybYZIWNUZLY3F1g4lhiIMBZocN3A7Fkh2dxet
54K9wmGYPlSNANOvXmRgQH6Yo7gSQyfwTF4jur9Ksb2lG82IXgxKselSiJHQewV1
rNKM3NZMyCfGToudu/g7GalRvladZqc1f9L62OnSys/+97CWFP/vwAO964tqKp2C
dXc8SB0j2AKts5A1uA/BIWzU15xuTIcLucKmAiG/zNwylrsnjzKoTPVTsnSrx+4y
3zcnY9BFHaeYB6BQlOF9jEA+Nnq4CCN+wFCnfQkN19gRiYEpq+9Km7phHknQcujo
IysXTralut/P/61tkG6NizNMFCK/jryZeHEAkIV+voNks47ac0KJiR5vLlQyKg25
EgTGiCW8ZCHZP+spjFyHCLRgS/UOH92z8frZVUPYPAODPHcgdcnRteGLMNQYAW4I
sRh7SMtje4ijkXXzp8pMfJ1hAlk193/b4SdnVFUr8g9rzAc8cmNovS/mrKFTAGMw
J1qnOP19uljNFHhw9d02tuKWZJU78FgqdGczyCN8Lzy+pfOhxG9wGWVHmgZrHVOb
ECTK/bcX//3tQSAafnK+p+ISB3UfGeMmn17xQYGctnTV0IERLzZdENF/nJklM6AI
wNaSXBvIhH0wx0A0rlwUvwM52ZdJEjTBiQoqm+/69SB4R/fmsXICixZxUkcZeEon
vsVcaOgW/5m3NZn0iLUJ1470U+y/aDRDkg2hauhy9fxg6A4u5edHtetjubVGHUpv
u1/RF5PAYQ/TtCRkz1WrAB8Qp2P4+duFpn6gHCkc8vCAeYeCuOueTTGG0uFcTv7o
EPU6Le+xl6HmPeftt/alFDGmt3APE+MMuNDhksOZr+OX+rhthRVWi013wZnEHJIb
uH38cQq/BfTBtbiwxLfwy66r4a62fpXivbDir3/cjeZ6Y4adlyn5kCN5awVpqo7R
tTbtwCR7lUd1AgZgRiI+BGP4LCF8VzbRApx551gpV6oeh/nJ9LCEZ8aECnEaNET9
l8sbOFK/qaBVEoiqVKuSH/PyiWWlc+JUo2di3reEh3Pn8lAKHUF13y+lAAfrbiUk
OcdJ8vXyxdLcaGHeekLTkrQuPuOZgvdF3d/J9fYozP20royQSxo/D0X9B/CJpK/Z
ldMCDlE7En1VoUQo6QHxfPobpwzgRpVaIO70UzNO7BxEYSBUVtAJBJcPRyYCqWwK
409HkbKP2mnVqii2p46kao9CwQ448fAFgMGIC0gyTnYxwwO7Um3CZxbla1JNEc/V
/OLUcGFs1ryQBpmvVPJbM/mVfJiFiWj+Gu67D8a4/k/PncSizlJhBksZRuPQQazx
WtP6u6R9YSDXBdqxfzx7xF7NRAmDx1Xob2B3ea12LKRrtDZZaWxEfpaWr24faidJ
iCkuvvZuU80Avkp1QkCWTVEJW9iEaiTD8UCuzrUHFLB8N0oMnQjuXQEMGunAAtIv
s6qgqTfpKXbha6XgH3MTXMQSuejkIP79oayMRVcJ4ImGr2DvYmDP+USU+qXEUCPH
H7331tJKt+6IqaihgPO3nTwlDYfNkvLHhxHAkBbdbfhKu/sa+4R3tWR4bO8ew0O6
ROpgKxHsWf2HLy7FsZ8pw4jYDynxHajsZM+XHiRlKR7A8O+/uISZMfNVsPgcf96T
lZCdAx8RSWSuH3/x/nbAXAf0+sMS/A4AVKg+8DMoSaUrnQcB/PxfaBrzq2SYKdyK
lfJG01dFNf7YVDR2diemvHiT2S6sb8eRCHxBmm6sPggPwjmcG+mVzXpqdywtx5Hq
veVAWBaJq3/3yWc+9i3IIwVHI2yIWEpVgyudqiSjtjz3y3kft3Jgy82owaP+kNBT
fzRjs2GM9mSSHO5K63eVaTcEaYEgnkIRR9VbgMZFAVec8AvRDp0LD+Q0uXzrz8FF
33MGXUosFhPFtihsamMUzWWOotkAuAifLqaHEd6tSZmyl4L3pJICspoh6TUg3j3Q
mPNvdyWk/7khe8etWK/TNN2S/n1nM21t6peK1Inc3x4G80EtIT5pRabibLTN+phe
NXzGs1CV2jax8x7X43VHw/41nmMOQqed1y+9OqkYcB36E6ws93Q9aUTEsMn0IinH
tJzMI3cg8EpzQ9G1MeAebMxYIaIi7MHdQZmljmzazqUEODJw16MCYymdud56VQQL
vOAspHBZiELDHvzXkBvM36EJhKoO4D3COOVZqXhywX/ZWwYFBIVYutGa06FKy8oB
L9miNS4N9AnrJIz4s+ooRaobFQAl4zFfIud832RENZrnHlWxUGAGzI2cPkb9eBjv
PpQPZZWDvt7DE99Rr18hgWdh3fDYcnhy1p4cpanKTLpDgb0xUEEq/9RaFrzWM3v5
q7QE5bypCoN4hl1obwmdpPb1UzDLoY1oVp8kd7E0ogR0CdILbdvUnZwlvSXwfqRy
0Gt+ufA5cYY6Bor4WqYFtUG5k29iJy25BKI/igKG43TMfja+v/AorybVnC5IgA/d
3WNhDUw2+uoroUWiS11Ez3wu5PATlchkllYvtIC6NqCEvoG8TAgqO552TIeifWiv
+nBtQaV603PwhFYTfKnQCa2iqkFoDpJ8DXWzxYy6jtpdyVO4ZYrYSMRDL3OBJXlE
CZCrTtBM2i+zHHxyz1lfPk+O0b/t+bl2OAf7645uowkf73l4Cpu/mR6RyCYRf2RA
Uhnw8N8z39uJ2OrX0WhKyABTJDDe641jg4WclGMdjQfAFMkDJrsLLxXeKBOnYxsV
XzECkmU3lpbfyqYh5F0jRxBsbesDc3OD3WMiOlo/mJ1yorngalaG3ezvts6QxkgW
rqlMQX1XXa3+7T+WInVYlBJ+rPKouKC4PzYXO0GMicuxS24CkyHBPXfPFudz+CUb
KG9d7zEzcrXA/UAbii1xKxL0IJPTsCIiyqAgsMkRlua6afiZW93c79DKmJqL2otm
c1VYHqfSecSQix20GwaBsstoTUmV7eLUYB5UOihSXQiXgimHXCGCH53Sj6BhmQeD
dve4LN7PGlr/OWbUdUFr/Q+Jo0nXXGuafZTXRa22l5CW5RYCRLzDcwEOzwcUMAGp
RlZElSFVFqv7L8Vk/A1zcxgzrdPlTWv23cJt5W/2Bq8jSOxXSl0avJJlQiLVbw45
dW1psx8zKBfeEmJ//496Wp+RfdsspFU1Du06PwmJ+951OAN6wqU9WcOpsZH5/Ssq
Vtqk+nAQ0TLTwDLTNBF425o4X44KBQrwv8p2BqSLHpORb4XOxx1Qgo4a5wSCu9PQ
/vBUbsWx3SvvzJgSt0hhJU7jBmckF5vNGOLKeUn8qqHa6SDGqd1/LrnWWnO6Vp7r
WwqKW6CfoXnGEc9vtgwhQGPfePW2Cukm+/bPcdcJML7AcwhsMRnsRVVIPx+RG+5F
bOb5tUzIdTCzQgpS67ZGUZae8HtBeGvlaOI3V/Ho//6ENURJyZqijWL/aL1F5sR4
fihNmbfkSx25lA1vv4xpa+k7nUcV0B8wult2ZJgZ8yMUbkv4CdSuNDf7L7ItevJH
h5biXkGelONX0KrMXOIZg9mVr6s4RrVA+ohHRJOfuICbIovKytqkESbPlGAZcDnM
4Bn4+jacAtCbz4ax9Yaum83FQaJBQBDHDbTX1Twv84hTcc0meJTxQbF3zuQcnkH+
yMEN7xcXrwIGjUAQspOWkbcHgd22lK8ZVW+ZMJMZC60TC9MdjFbx/3jEEsuEZk4o
uJnl4U8x+FHAQ7AxHPV7M5319di39Mk0GCnpoojOnsqfSHJPGU+j7WgM6D82W/ur
/ALCxuLaNAjcPF39CTuj0alJnhxc4bRUpDYBBg3MRIKq9sdQKU1ZW9Pli4oT52Hu
fL28h3niP/hCfHvKmW4lKeWDJ15/qr+hS/oYgJqBs2PmVDE42E+nJPF7odNk4dH1
NZFBMdPquSRqp88x6KI3GYvLvpT2fVgajOwKwLObyrRqWHl0TxhfgBm624vNR8HX
n9BaCTqZ2GJ/pRp+llrnurv6kFLGJ2rZ0ykc1LaGNEoFGSFbSrfriIZKBZbYtSSU
scJrLjQCynUA7asbpJwV21oRnTlGkGhfS4FakjTFL+e4n4l/SsZ++6eAtd5YPGs5
tE9+a+kk01FdiaNVf9YcNP26OQ4wJH0rs2b92EFVUPJFgAVYKu9yyoyKSFNA6Eop
i5r7aL1p6MR/VqfhLSmfDbhMW6u/2qkZbLhAQKqPJDqMDYkAqvRbVi36YnE3VXkE
H77YFQYHyrYMm8ihn+6mQRTykKhjOK2L9/iR2Gb6H7RwrGtS3Sz7syRHxI35rXch
/ZxUrTtS6+pKeEXoJOTP+RkmT+gsdMYM88BYN2uY2YrQ4pPUJQ0Q5I9n78TgfwhE
jkxb+lMpEDrSAbrs7dMzwG/Ou3dl/Z1YuUI/gsi5WnCPtbrbiIuKAa0Axa7JJmw/
Gd6xfXLtPLg4A+sRhWa54DSdu/N9NasMnu2Cn+ccbFEJcUzceXvqCIMnD3IXm+sr
G2httnP2WdxvsxSO50zrqH4fgjv/sNyjLbw1BdhlUVNAhm9z4MTwHSjN0b072dzv
lXw8NLkYtwpUIhxjP86WpUtVV8/itP0JkfKXGJFoFYws3OktfCewcDK9sqeNMOPE
JwFYyB8WgQ/Tvaew6B//mnU+gF6vjZXTbL7wJ3WkbT5MEPRmCKhzpgyBCRPjPPkt
qcZ/AjKi2xjshPqGm+TNkd0H++mRJfVPw0MHm0dznHWMeAhETDPWtxtMwDt36OQx
svYT7LYUjoW5YQtKtciAaJuC5mZi/Dgdfc5SNlIufQBm3m16PhJHHCXZuVbe/346
4y9RddeEy8sHfbWdf2jHu58BOMxdsYcOsmSSyYUcW2XDDp2v7P2i3PZvFMQgpc8j
iu3pcyPeOOaYSPf1qxAhv/e8R7IdM68OQG7Q/YaEZy4oa9Wsq8h4gzgxv6NOonHj
j7uK3AAlje9fk4sh7us4GDCjQHWBio+cW1LcHMgb9QwUMwOru3R0Tb0JPywV7HuQ
KAEgQypirIEVb/8/cy/0MUEKtLIObwIctNNYZ/ov5GKqHpZnJ3EThmtvvSvdwqPY
w67WAWlQz3/VikhtpMLWsRlR/kozYBxC+FYFiQxoLV0En43S/2+Xf8xR9oBQVrxS
Q2Ema63K9v8LZvVu8jvLCFlXQjqy/7VORaBxVRo7BzPgRzqZiQvMjxbo7WcDeLbd
3WSG815/YK+fBqhhK9jeEhXuSrCEbmVP6GwHD8qdP/WLDjckyik/cZXkurH/cx2f
iI71JQiYTf9WIFbnXpfV+0EjPIGDm/gXtaGamPAWx/AOOmiqx/QI5WneEguEh7TX
tTGgqZ0OvRcDi3wqJbCRch1jMsvvo2jI5LXQyCt9ew32sRHv/s6yr6ozx8/KLH5h
tN1BaOw/gbnlwb5OzoE49mqkoujL5eAhguVSRrbQspv4Ml+F+YaI40/StP6t6jCO
OQNW+30tCDKjfpYacdWNicBs/t+sUxQZZqMjY1x0veFYjZfBjxxzYqpIgyvj9puY
f4CGEq7UMSos/r9TIDBuyndxTUctzzU5Vu3TVzzTODInv+iabGHwPumPDZlMNk/c
RTMyHiBgPHohvOoHhdbLJJKul+Mn8KxU3bQngfI8Tdr4wJb3UYGlh4BSfXnegt03
Gqnxz7zNKPVTSqzYhDf26Iv17ftu3Lf7/XmlGzijFFULJu8ftvR63noo3xCIggVD
HcQS4aSQsJJbymtQeKh7WZljWmhi9inleBRHqU1LVUK5JwmQsnypg2jr1IXrD47i
KHjCUPjjswIkt9buCcAmtEYw543LxgSQWM5JLtVnnqtsi9GpUxnDYm9q7FagaMjg
sCZzBrcQzZUaBX9sqvNt1UegqLX9Lqdvf5rDw82B4NOXS7OCfCwadRl94JLPFw0U
txGH/+HigWRwIKbalElPaDSLPcNUz56rzrX96LLQ9FvtV6XOz5aFm5YG8N/Oy/7b
lTd1i5Aa0vEEsUMmZjzEYiY4yasWqVYIvlDzhAlMt0G/FIYY3HeFsu1Si/4A+TwW
pkT3Hs0eYC20opIdiGM2aP7YwFyi1fpSs6xgQeHjwx5Qv6fWQb5FKFotIRa6rtny
Jqh4OHTOMMv9WRFk0F7gF/lDNm9nP84n4RUWxdnlP/acM9RSZ/l3OdsVJPclzA4Y
+pX4R2/rzeAKD0Fnco/dvKmMArvVcKcwzPSx86Rho+DydjF06qTFrgV8iydoIGo/
XCXdLsl0RyRLY6bjqJam94pl4wTpE7EkS1C6fOgQX/ppkC0/edtloe+dRFE0Ip5f
31UJZa++U8MZVE4lPNV8n3Gd38qNHU2PHaYw/zkXXnQbwpMwgBbnbi5lkFVZ4IIe
Sdj2yW7ajbFyPkmEuPxsZPhuPDnEZuOLeTILV4iJA03nRXv7WefTsFzWNchfjNka
BHwx729hKZBGIofwta+h9fb++t8EVdlDmf9X26xa4FwuxvGB67xI4OmOYnP3w/9t
MqN6S5pCKSWlmQnDfQW3hbHeI1nEVNIhqIQmbgtJmx/JTmxePAckgDBx+A8ihopJ
S7VOQSuunYY6CsNQnirWwN4Rwx7ZbpCMwnVqzNn1/ZEESoh7/RPRM0rpJTG8AlL2
c9kK6WgpFG6C1I1dhbWwil7wKYkXpqkdTrfBW9M0Aa2eSCtXpgPTkPQmIaMWJ8FY
5Kf2AeLUkFlMEYuT7/eK22Fln/ZXty5HlHwtU7A3hHJ806tYnHPz4RnerGZwlfMG
OFjrnflve4K2BIXAJVjOt8qzl5cjNnDW2AonfB7Q3e9y/jAQk7WQPQNtAmulwzc8
Csmg/mRPbY47DV69oMpUGjSwOs4eLczS0osc64V4k1HkAnAK0l2kxoUuzHrs+uw0
D+UprQGoxtJGCPdBMpVkOypKl1v8+liZuwIEx8r3ybtQzBnwaL5BzUweuvg6FJoz
V/gpg4z8xTPOfx3UuAZ+ZW4llM7ETP8N3oLRqTJbbsMX7/IA282ViZqea3oF1bvE
sAqxXub6/3AOp1tTL2lpAbsltilst662uRlMDU3bJoaO16w6gMsHGXkdEFJg9mHc
0KVg1ADfjSWlqPKhBmMOZXqTZzBNeZ/MqK+uZZc5YtMzSrvHww/afgeJPLwSw+HX
kDOLtP3pD6hDRN4259b/LDUxVs45ouI8H6e49zTzmFlnMYLOKhuZ0uz1hiAA4kE1
9g14ryALmmkHPheIMG/Y43RHJkPWodJfxdZukcGw2gHG3HLguLZbG2zsF6OL3BDl
a1CPlY3am+dqhm1WBk0hignl0XAzT5AxHQ2vzd8hfq8z/S1FhLnEPE+tyAkhtYF4
+jyLsiDVvpSuWWvylEMzC7aGdHJghTJzAk+YkZXS6wgMs7iphP4EsHoZefD8VRbI
EFWRrSWKDiYmWpogaCj6JOrcMFFwNScYxLvxZcMLCQ3Sc4h9bUZbf4LnosmAhhQ/
dVulT2VUIfMvCizTOTphixf69XWkI0dvNSVxRqfJUDhxmIkMtjdjfuEEAE61hd1Y
J7bi+zAXLDQuiWGzI5cdvHVIgYnfLEUPXBjrAIxTUBb+B+oabh2tmqci/t3ndNT8
TCabpYqwTWXTq2YgZH8+Ue4Wlr62pQJIVZdw2fkXwhi0k4anVA8F8NmfVTxnqLjW
tcKTXvDSv8Nm66QeUTbb5v93U1vWsnNWtPb7/ebS+N13Wjt9y/lNo+8/Quj5MYOb
uFKozvD/KW/JWy/tqjFpLCO15PpWdFv2vtAOzsZsqxaDLucI9tAGDODzsAUfZLvv
rxwA4BetxXRGzfb4i4GgVD271kOvG0DqljKym19qzZduv3wiJ4nzX+Zm6ELU7r8M
xVY7l4aCMvIJg4/dhx1gta778vNYvzLd6zfAeO/UHjbhpKZvNnzAc7eugf1l4oKp
eL1Jk4w80pDlqz6iy+4mdOR+yj1lcwsiOD1HtYOKPRLi2i2lyqk37p5KgS19W3H2
xTEpagka3kYUE3jPp9H/rNo5URouQX/4oD4Lq3GbWJJR4iibY8Hvc1jmwTdHeyce
6j4UKrpbef+igPZexXyfy3Zoml6jBPajyQFELUyBmwmMGY4RQhrsDJpMaeaZmf+l
CuI+DZv6xeMb/e6Fw4w4+KZzblpw5Bi1+NL8tyFlBC87kk8EeSSvoyMTaLmMziLL
SxCWH015pYe3BmD2RhYth1hEjYIkAByd+p5qRR740Osq77IvRDip7wITBuhEPpXr
GpymDFU3zi5GyPkhCLBz7vTMYi2lb/PgbPu1StktM3g0arca4E69BnspMWfTq0ZR
GpR0QdCbG2qduFf4MgzjMp+XZRU4RnDQYlnw3Xw3hIpK7OiL/DEhliZXEBwVRuIs
kWEajRRoYEK6d8DnJm3roJ4rT6xyIkwxW1sjDSVUHk6moWDCP/I6xwqzl8X+hfe+
jAE5Y/2R+HViRjUKdLufkafKAp0BGd/Y9GvTFodN41p0HYfsI4th5A2AJos22W7H
H4VLT/6mG/HW2Z69xu6OS3CVAe/ZZfXbZBQHtQzy5s2Jdk74FPeUErGifzFblolU
W652ULaSyxU2eHPKzohNt/KAMrQUQP6tTHkGpUgANy3lF8yXJqPU7LbX0/kff9+p
539ossCS5Hz8za44o/WMz6L7rbn1Gc5oUqtLIihMW7NqlRjNzACi4om+bulo7ChM
2aXpZS9yjJHahfgTuUVZEMnZoqwr0Cms6m3A5/OwOMhc+BSgjposT9TWq2ZJFqwi
EYr9At6R4/jeyHC9gnD9xlcnedKYlukoa5D5AC8nnAVSzqXrER+ab8y4Jyhd8tsx
gvnWtcuubibq2ZVehzW23sDbgx3gXGKP49mCskzUwherRvxx+EtsvbPb7jozcmrK
SlESG5zE0T7fAFx1P1VPz30WGQQTIr0pJuCCfLIx2lR/XM+EgRx2FcKEP+9T1G69
7UBuFxQXEerN5ikgqIAhh++K+wuTj2Nf+2qWEIBieQNBdFKaxODSSNk8eHaZrYVZ
LGMgnY/XSoSDlhz5gs6Wj+DHoatnfFCLeKiCCuPOB0Psas0W4dxUbuJ8MlelrNrr
5Dj1UZqlcRlejyUIrGe1gMwK2uKl66UKczPuI/vVfs1BwcAvEpPf2A+SmbZbebic
j/UmKrbDdGQ1P2MKELElR23ILbarGiAZElOgfbHog1a5+T+6ERQXtgOL78O+CiO6
bi4fl/VusGpxcB9kBXMEiWevCHWFZvOotf3+Evdpi6QrAlbqv5YfoXGVsV00X9AH
TM04UhIKfR7iRrqM7js6dKYtq06nwsTRNL2MVAIoEw+6lrvHGdgd6Wdx9soP8Huk
QQspmyIvJ6v8+xnmGZFjqf7NVB3bq3XwRPOQxeNQVq8bA/G6QkbJkGR71XDJK8lW
rp5B5jheiskhlUb6B9wV/dhJ6AUtOd238NUVfrFXgTy0TQgB4Db7zXsg+Fn3tNR6
1z6Su9WuE2SQhX/GcRWCmlyqLx8M8E0D1R6PhcDpAn5msipujD8oqWc5tfsZ2JyP
MGXhyM8zzxWkvJIujsWAt+41oKUkAN7NhMb4nNy+CY8zZ52HFHDmggf7F7OY6CVS
PC4vc1Xtb1b151bnNQxziwaWNNLzXaHJJT1NLZA3pZkAEwrCqR+G71oFuW1TZqyF
93M1RBF8gARUKhzrTeWRPvwSY90vbjIEG921SVHBGBpotikEv3LtuIpVANTuBtU7
xcSnDypYfYLtZ/4as+9ZdDmt+rmG0A8Cb4BUkUQTOeVQeX5ADTEF+jxUyGx+tv/t
RjDWsuY22T5MnqBEoSvm9flkzd/6yzjFSD7Wctd4RHb8NhrVRrxUJjs6vsGF+d6/
4PRNNIGt4UC7/dG1YdFFGWpyeFSaqrTEXSiskog6THHwm5G9aoXmjeKP5+HJejMz
6pT/mE3b+oahWLmGlbw8peCdgibRgDdYfnHo/UH1VjI42W5MR5dA9rXqO+Kz44nV
NY0pOZxPT+J6T1RfZfWdA40h3bH/cwr2ayJSmfwwyxf4VvjJV4I8TnmQmBzYstsX
aPJcb32Y/V4O4ywar0S/JKMVdKaOHOOzZ1Bpf9fzeZ1PL4XEkXUEGsINvCxmwJIe
yAYWPwc6L27uAaCWenZ/NaTGBx7WyZGPtpX5IpsXr1r2uIojrjtiOoUHznPV3wja
VHAuXhTagR8ahvQdJW9fuFOz5PyzDYUX/LSzEJ/JTN4tosNKEUNjyr6E9zn+JEYH
T4cPo6JsROxCN1qri9wdm4k3boIeDT+1yjgzCiACrj8+qo0/6IDXTggnCc1p2IEy
lM7tXuy77OLCfUQ6OXuPjOAyKxQH6fr8U7tsEMsgZemc5pa7Ec+fbpzv6zbcdc+r
0lSVQNO69cJfU7+u6SUuqouU6l2sDwV34d9m6Vauub3L76flbmBGXNA/6yvqyDtV
hPKc3J0SyOY2JNzHRELlfxrPWs7fnDpHRkFY54UpZDmDgzy7gg6f06IkFwpJKgWe
xk0o46kTpCDth/QhHP9WR0QqomxqAdzr/XzOoUZ+Ta1zyOMosIenQ8mtkfARtiin
nfH/r6zZ++FgXzbpn6B2NnbJm2EjVPeUOTwF4sXSWqbvEYco70aFOTwKiFH9aHfn
VHFH3+a6lKrf94kTQ5ws44BiaSdRkTuiMKDWvorqvL6B+x1/wabW0x0gloUJJ/03
1ol+ctVwqZddwAmrIn6szIUS+8NZnJVSfgjj0wfF4EGrThcvlJmw4tNX2oyILRvq
k2PuEfdxLVkR38YzNU0URNOT3ie3XtXZXa4zZErsK4+vG5myL2T3rx4Mwy6VQSO8
dvn2EfUey/e7m2vlahekiLd6dN07xTFI4QgyItx8tQjX5+2X81GGqvr25MeVD9BS
MzrOKhuYBYcjAJOIFRklLHDHNR5W0ogGwXv1urSdqMCKeND2bBv0iLSyMzbkIAHo
JMPhJzq5CRaAGljpjEro7kAdRBp7vwG/NeT9DVvXWufazZUqQDUud2mA0LOfz4PP
pA7KpUadeigm8nEUc1jiNj9P4PoFYEuqhAoQj2EGaN0GGGk4lZeZ5324JmNOckZ1
dZcoIL5XanY65eMkpizeWf0rs2czDs/crcXrN8jZ3r4JzDtWnSsUPikhc8JbFGDb
CLZC1GQ6uz5muwf3vJG/Nh+c4QiURwSbLcXVbu3Cqon+fejKO6DUlzF9Hjf1jgfV
DwsVGnU9ydgkBneoXoo2ShMk565plis4gezHpOnhpoX5qGpY62OWSpSgyEtEH7SE
mavI5/NGsYuYFPulkZsZkOsAIb+o8/jky7ePzntsCsjD9ILF4CjXrIlTH9IWd93B
ikWHX82VvRbzxKeTHmEStIhnLKgfDkqUuVUzapLsXvCBAPznf2ltEqkv/1SqaQ0p
Of7iedyAkJAI1ejK3Dme9M8J1s5WReo2lmkYoHa8Pcfulqo4daXexgvQ+JGgpMvz
P9TZC+CbHwka5AqBMracB+0henFWW2pwwhl23yJdncx1roy9SbuIe2pAx7NDQpQg
YwfG5RYETbuPyZ2md95KNFqftPCKVKH9yyA49oDKQRxdUBD5B2pxbUvBX0usFnIS
frcgwZZSC2FIu13S2FkhyRi/OVvradc3SgijrHXH/NiBiC1N5bNoxiSCUTN8+EUB
xeetn3U5CRLBi8SEPkquK3RDkkP4zz7c5lapJ7+OpLr+gilLo/b419GzWtLbEAYw
nHzZ9cNubY2MVD1jJf2ypD3GQReL3hC/NqyDtWtYly+gs72amQaW204yWCJilQXh
dO4pklY906vvBBZ+y+lfZ0EUc2c8g9RUimlnHI8WqcvNu1H9mO0XOuWEFk+VNXgq
ah0etrXJHBqwvKq3hoH17on7kmSSiMws5jfOsH3P8Sb2ObSDwKZE8lLsBwet3uoB
mE9Y/I032fbJSHC7JbmS7XKualfT+kc5VJWkGSPM6zDVzwXS3hu1YA0ZlSWlScUk
V4hvyeh/rtGDeeSxjO9pxpyxOOcDqyyfjjqJDvqhRahb8n6zL50TOGe56cM7c/3p
rdLJdt2gN/QWCisjQVI7onoSLqcIEAKwW2O7A7FvwtXoygsconRL7cm5fIUK/iH1
K+Td2q7IzFyWqZDNvJK5wvYDS6osi/3W43bbM+WN8eX3GK+GohUUhNhSOr/Xiy8L
ZlC6djkQVs6GGeJfWaMv853PSi6/Uy2eCYsvas7KgruUePq5R/irW6Yos26N9/uO
wZE8vV0UYoh1ySp/6xa4pHSKdD/Y5bubYSx78Msps+8R6DjHfgGJNsBm4qEB8DAm
ONWo+mIDjv8JE5Z1Ho9Dlog1N/PQkRNSjn/oRfGHsfWYLgDBbnGN2hfteKwl4Q5L
TUcuSkjMYXf68nN4QHsOaD0A4P8Lj+0BM99fDDfW2mjWqffzrmo6oeOZQ2qO8kYJ
BG4aIh7s4aezuwZdfI1KRnYnDoNxOAcXHggEPXcB5GKuQBkOdij4bF0PlxeDD0KP
rXnx2f7Evvi449EV5ZxpmPg1Yop9/1CD7un1oIFHBe+Qm86UnHuwZZ8BslIwNLva
p3gYWnPl3asBZYP/RMGyzJHy9fWEpp1FVXbZYUHAr4JF9oE8K4xWaUPe9cA1MoYp
u2m+Hc8uQcUBZnNGmkQTCXJHOB6VvTCXhKcXnQRjz/2g3ChBpyuqhupF8JvXeYRQ
GzO9OJrTN+vw/ocx5v3TKseosy4jmO4A16iVilU53ohBDhcUSUmn9c9mgrzQykko
afvg++YZUJ/v4Koh3KLtpOkgg9Jagex8MfTfLIXLxtI3L71jp6fhJzi1LCQq8EdS
lcmCSs00CvODNDtjOxXOHsgy/TEckDnDRRjySkTg/qMt1FMCrT5zu/hEk9/rPSfh
7Yk2kt8deoH+S+6YcP1SiyynSQnWEczpHhyCWCi5+lzf4JTj5hYdIQiGNPkqHgw+
r4PBeRPwyCfgPxHIz5KHIcXY4XqPpN1e2K+rTzGNq3qU0M5XlN09A8maGsxD7TQR
f9g5YTE4yppVUEPHWSIyVS4I3VDAJ7ZnzL+wu4uAcV9MHoTuSxHa3+Nb9+PLeSno
YWmlPhrpZik7KHqk5G487jyOehcUr3cbsE+JFl6INFQ3rZk8BWycr+Dg+ZMvjCAN
njNJR/qWQigpN2tIvpMMvlpoLvLNavw4XoH1ytph7yrH6E5gY82Zcp/DnX9VkqyM
4xvipb79fhv69AUwFdeKFz4kBp/Nmvr/qBeweis2o6oKxv/UJmKJK6RRlLJUD6rQ
IN7jkKt0xM7TeOIgiBPc9qVu5Savr90Lqr7iHHTGwRmMSVZ1Cf1WaIk8SYCOKBTS
YCeOjBmTdZMm8HiL4myc9Kn7fxhmUZ71/pu8cMAQ8jzkd/1LdcKMV06G4J5i37P5
/h8mjkjv6IbnKO3q28mndFSMdzseU7nXfQD9B+p4i9hhaxRzrMfrZXvZta4KeTMY
8xNReQYLa4jhuAHGUVtHRXJyJ/L2QfMKxCrzzYxISZcnqrHtn0YbC40F6JRDcVBt
FDbHd1xHoJE1xzVb5kUq3Yv9u+RfMe/UB+kw0rxNUji/Cm6gchE7kCxlMrKT+AEM
hBPUiWL/GcNoBx0+speva6ZPATRPx7d5O8XUagPjdNsST0fWaf/bdsvU7fxMorhQ
5yN621Q6BQyq+Sg/3dJrA9P/SahmfNoL+DS/hrGCPO4bcr0j5qs0rIPOIvztrFdH
hlgPUBDqUjhb85PxwRN1hl9Nek+mbmmgnI4OvQ9k88oVGN3e1wgYEoNU4jCnnUkn
+pPX/niZWsXhgjevnjlcGvXkhmAtHR0lyYg3uXZXR7DpGQetEhXJn5jB9tUGlFUH
lMm9xAokSPlX7YGaASmHzMv+oodLL2cnmxlNbD8YBh/1D2C+u1hN6qJ2zk3W1ZC1
Ju4C7TgB4F6egzKkWSnzBF5XD5JL89TeytiEo9iXTW0eThG3dzZrhlNDOBsafEXY
M04KLI52xPPEkRjEsXWeF4yBNc2vcqlqDPS/FFxziT+d3o5yGxPZptUYHE0HECSF
lUp7hJv+3RCuA6yMb3rOhZoQcFSM6uakYL5TjB4WK03FlPcyOuXzGwRgvhMVqkP7
5uXJhtyzqLplBfttKHCfCphGhrqvr9pUfjRUxWj1LZCHPsv/PKq/cT4UdGW+P1ZZ
qGt7VO/0OdOcpy0Vts2NTLghEBztUrSAbberLyHMdi1VpFRfVFikBYotTp6qrmxx
TatC3YrspzaPyAc/DHKvdJHMIVB3Ktc3B6Bn9DgB4mHLta13icczQU7Y7ob3Xkwa
m+nAQTF7UL/Z05nqpvXiZNsbAXE7/s6F22ou4NuiLcrk1Rva4ZWSsRVsQrBEqZVs
s3g7xKgH5KrRL9H55K4i75IeP8uSqD7TknRsFcJ3rs0lxANzzWFyGJPPg2O46iGU
85bX5p05FcK4nKIjqzzU7nRqReUJ2LXsTDJ0bFPJr+TIgiKZ2at+gEbhcHlwUCwG
264xZ+3zEgIhxlMELPBurAZIN19CwDhIHs+p9LCMgrsXSTBw30yMG0nVHrcplM+p
E9X1BPbqEP1EK31F/bjgH/JwPSdEHSDwFRaUKj6tEgxfsase2IAWyboT4kFU6GK+
7KedqxANX1vDnFS7n5AV2Kg7jZ0J+mn1cexgLNZwnaPKHJYQWgQmpj4oNafJaaKA
9CKGDNTDDgDzJYc2l9qBAGIEUSxdMq+YU0uk2sgQPrBmGScc17SdaLHs5cltCxj9
yM6JVYx5wZ+B3Ydce/cD6G5KNRF2QGhOv2+7U9iGR4bjKZGF73iU3Tt0Dt1U5I04
X2/8pPsxjsfYySQdknlnlMOlhZ6f1u9gBiQDS/febaMjiseyFWBD/gbTLhGr6q6F
kTozVWhOl4kl1LFQyf/4aRsAI0EP4KDdhC+spYZxjkNXpfs6Cio5cTRNy3BY+8S6
rEt2x08HW76GsByiaUCKZBsldd6ZmGc6+m9S8YyGPyy3BTiha/V5dzJM4ak6d8D4
vRFSSeFLTRzfjXPK/gsyplGM/pjMsslqBxFa2pDaJlbgPtl63f3jBBn9gaqw14wz
OSFI4kI4kOCznw7AyhoJodZwubiFIKySuTrKYCBd6ggZgwcNBqEO16LD7L9HIjaX
qOX9GmlnEEshVQeT5ESXGjfCn9SLwsES2BJpiLOqifmMjEB+6qIze5NTt9umFkgI
ImPpyUdsvWZaKVEJNL2ElUR7WHwcEfJMGIM+jTkQe1u4q+nTAv1L3y0vvplMZRBa
VO17ikOJIKRoE7HGALnrAJgMY/BKIb/q6wBGG74xU6ynxbtWcUbVptrR0ocsPCEI
bNcpMukxaeKh0EeOOLNuNsMuUSsDIbAqRbHi+K7bhV87F/Df+1TrSfSYdEtjUrnb
SsLH9IEbpz2qu+NpkRLpYjHjhnW83YPC9hUQ0cK9bpwO3dYbuJpdDC/sjyIxjk7n
lKoNEhDWSY/M9tRH5oJxAz8tB4eNN42gkeHQ1M/v3YQTOYAGGHnyuU3QFPloSvuw
8q23p9H7YUSapsL7i73T9uYySlTqmMZPGsdgXcbpKhrtL51NRRoZ4fKQ+2Rvwff5
vtucZoqr2wZWmfRBwAdeHJEfDYS0sdOR6qOm7auLa7I8bp5E8g3A9QA/aScK2oKl
5ebzUh2i2uLQJ39dAvVDgoznLAXP7222U1Yr4AkP57sQ3snXhRBxzYCwi/03soTf
0Yqum4cmmsAikMaLR1epOAG/4nmAYYnQs9MXrSFaQDuOHC/mnZ46iVwVw9ziGJQ3
7bpdyXRSa3xnxAWv6z4wp9awh/q4+yu6M1Z+vw2JINqt9NB/1siuGT5zVG2uzZLP
OTWB1mURPKrCIrd96sPKWbCPMcUhMLdruVKdYZ8sZhbs+U6z9VtjYnIH3Rphsq/e
pRyRE/onfFIJPGkIuU3qSlmljU2CO7y8BqBK8chBI98mReAxVXG0esAGj8HjbNvA
iNOGoEdLiu0UEV3yWb3EkdrDXhgch+GyixfOZFx5vW7Fcb1rmIC6s9rUhj5X9Isw
nGhcWTQBGI4Phz/ldc/83l/PAVuJ8yaHCVWbuR7Q5i9pDKPtoQ1zoB7Vr9uA/dLt
tMPa6ciuasWw7qZAEdQO0o1DIkCH4pYnfKpnn0CwpYeil47DIJsLrLk2Z2yedsS2
9uMxWhOJYYbbU4WPrIsqjEb3CvaGN3lghiWbNQKdXpMJV5nCINR37RkF9Zii7Pza
FDkzjR+PBm0gJTlgAc62ub6Nxn7NXIGS8uQMwoOSqg5teW/RCuNMD5jYOtoL6bFG
gKD9XQkVmPlPtxfFRW3PZDEpK/EUD0KDOVfcoNnJOx2tljtCqf2E/Ugsg1QnS+f6
q2g2C4ykTHypk+00+hk6PeXmm7DUy0XlOiGho2wtjEcrTnh48xjHw8UKvHtQtqNB
0L4zdkzcoxn82LBCE6HNXVmpEHdrlkecaa5rPMdpGK13ZB5RuUtqu5FBidopzBQv
V0ADUOVJfxX0B2albth2xkrEA032sHS2id100BQtqkZemnlD+3UCjur3wxtpKoHc
ajsKpn6FdkPUHuamiUkxQpdER7gf8YmolyBYy3BExxj/7Iimyc0G14nHm9rHxbtc
U6d4GVh/ZagWQNbgyr8ZRwovNyhkFVp28pgKWy9lCRRGK4vOy3bndbgFniUkPPHt
yiof4a6180mv1qF5EFyqG9AX1s5il64rQtWc88tHJoHwItF7n3I+bOuklBF569Nh
La0kt2+OTa/soH8n73s0zTp+X71sqHj1OYK2qbLc49YUE/NwAXJfqQbm+ciENmJ0
vXnrH/yi8Etoy8zISAVogPJB2b8A67X0ASwzvzdv92lrAuQcrnQ4lbj8Ov4HYH4R
21lKZmB5jlpkP4CYI5hMLIK2AkLCSXfhtfYo0ks0e8VY/cnK4NgNHoT+wLdog7I8
l2FlseW/v4TLldlfi01dBfYB1hC7YN0IFwudtdPvRfxFun08j+SrNyROvkTyzHM7
CsaSom+yhJdajsEGw5tAey7s92yB9M6A+Y+m8oZnG0EwGm8LcHtQ3Xbcug3IaxPp
Lyh4pAf3avP0JKvuEsJ8t7ZK12iDXPhdGSXscR+fPsixEwtmAhtoUU7V75prwloQ
poPpueDkIY5CYCYXG8u1FzGkXpyn8iEYihem7skKBT3HxS72smYez15NkNcs0+mx
ug5WtTxK9AZ1Bg+zrdIYA1HSZ8yQ7fO7rkhFXa7KOWRUGjPhrGnCDIvL2Z5cJGTR
i7qWmeainP1OLE11nZOC3d7nc4aQlWpF6jUTY9XTGb/cTtPotWb70TOKGIJ6/kfY
fUiNhAI/vjnek5CCQQ5EWe14s+S9UJ3b32/oxSFHdSyNldpDn4EaReoYla1zm7zU
DnRFyU/vGR8L4zF5FMSyxUP8y5l9fbvpFEoHIvbCstjJl/okwulBDIwYqCuNPSxx
Onngz6zTsVE9YPHrbQ573p8wFa4EogN2YZ3SnyiCRIvPd29opEh2c98Qff8CrLLc
SrfqQXmmh87LJU7HDBKsXB1sOgPGAWnRwip5klJCrRozbepuroevK1tlONdjShgo
Qw7IZbla1/WLudO/TpvN9AD3s47N3EEykQn5qFj6E4mnrjxfNTN5iIVOjL+sM5AJ
R9Kv6uRlLoT4oT8JuklSGmJf0bUV4KMWVgcMqUE4R8x3gj/joCw344g8NEQs6lG8
tl3LSYTpAhd/ca+/OkouyWQlbG59lPk/RvQ2bEalTRYpq4xrIa0yEXNCbTY2yssQ
CxRRxSnExaYNCFLjbOfC6kSdzdP7pTLaBArppxBQvhWdWBhZ288wVUFbbVY3qlOw
ucnoyrMyvp81QH5yZylkN+CfqLmkP9vMDkrmP1021fEHOx9Trzuv7Ue0cpd5DXkC
CLGX2wK5Q4+QT/Q7PydMiivxQ2G/Dl+sY4qbQl0LZ7oRdXrSlIUAAGqwwNEmomma
wLn7L9JFuH8kryUYFC5bGK+I1nwBplj96ZFEHpu1XnQfa28pRkrnDPAwQf5ZoYFn
1ph80tBVTOR5ohIqD12pvD3uyoMu7s3ZgqFalsn1KUGW63dTVtBoFJE07uncp0Ws
2tdRarmAkyt8DcH6viyYcwOxXCuu0gpKRH3GOyVfVJPqZL5XIg0Xu1BcmKNqv4sw
mDLqwwkKBgrbrfI4CbmR+YNqIImW2A1bzx96RlsrqocrWpjwheKpHMLdme3o9R1J
cG+zWPz3jvsWweKLjgwKE3jtLA/tLYk13I1uUYYmQF2hS/JyM/+oDdMKWpEIFCPx
QBTYp1+qTwSAoEStNoXOq/l2n2O25FX0FoELis+6uJpprAvYMN2V6p6MlWfUwJPB
qzDbWCwY2MOTmkCVdehZTA8MJMMf2dx4dqGYvr4RkHVUhA+bqKnzsqqoFkkN46Yy
Fl92314WSZmvc0YOoEGpn/Ux56Qa3NHK1iRG1b4RJEFOu/PzQqHguf0FFP9Qffgu
Fp+4nJalg0k24L+tqkzH7Y0F55AV8e7CHeTRXGCqGZFQ74B+5lu2B5xc0NNcA3xy
kmE2QzAe7c4AmIk1drha34HVzx0eh8dLUP78QrQcNVAJjANZnAatgGzyedwsEhN7
WZXLh/qW9Ys7jtD0jMutjTx3MzXJov51dumYnPUUKvJh4ZhHrql92Uld1rZes18+
u/NRymo0TBlHKAH/uh9lm6OLUZrDp/av31ipRIy5laHo7N2iSoev7U+adGPC0fvU
J0AznPWDY6hkX9NQKQ6ZhodQ8hVAkNWbX6vuDKuSQxCzSk24b+lJqXbc4Ec9b5lh
O91swqPeXuQKGjaHMgP7Ho2vRf4MIj82NJ2CrR3FsM+KRz0XehxgH3wE49dq1Sdr
4eFowhe7u0cQhnAu2ZArJI+Ie73JRi9wW87uyqpy62T9RcqOuZzyjSuXBLRRc7wZ
7DB+fZvFybRBoXM/Ibz3sSFaq6aBX/MyDkpL2Wu4Cf1o6Ao1qz4ptO57mAW0/CGg
1v1MJLkDk1L8OYgTuKY2bFgMMGmuzXHrHOtrv+J3I1Z8Iske4SSyyFJuPm8GGos5
cr8PBuDZjMsssK5pjE2ImJpBzF3XJDxHYgpLkZviPGlgf0bCeGgmP0/H8PY96zPf
zCRWZf5JQM9mBzDUkNRtqp1avMJvabREL/TrKmcnvFz8ghwCPrsqNETo280rKaCT
gSKHwKACUump+U10XXtrnZxeEnDrroqnTDDJZUmE2ImDy84dc0Ij9WZ/qxRaVI8h
4Tv7iMzSfA+gOhMD56fpDKDwexBeSur2DIyP/2RKHQYO6I4jHqC2GVXepF8c87I6
kdMJGT4OstS5HohLuZ8sUoDMGwaYMRh0qO5Y/hRmnFHbUV4EGKMDFqTcbIGug8Ll
s5YCwzY6U+52sVfGBvT/SH0XpWj9jWij9C/bkGKGcfNJMet+7gBvbC8fPGcBjLwR
EJ1xJNQ7YAEjY4SNfJxYTW7Rk+f1tHhSchQ1dek1HRkiNh6FYyddmWK2PYkkVBUo
e0shUgbHV8zP0QOYOqRofi2biGMD9Mkpru9PrrRNfJLXi9KhLSwyv/8B6PjcuXkg
bwpZi38G5YIDMNljp6RB6E8zRNrccsU4/KZ5wnfA3gQsJxKcosfrPEUQC7KArJAA
UaGTjNAYauJBREiWlvJnNoXPvEpn1BD9wlK1pW79z8TtYi7jMZuYi+9URGDqaBUl
houKONS1ufHUnw2+kFNmem2DlFpick45a0GfJXh0e3Zi/bFAVkE6XZ/G+Uwx6PSd
4n0lLULDI4hEXB+gxnRW6D9m/QC+UTJirJpSJQUU6S5cfXUHD9hx+TLkrHfn94tF
ngRvAe83FEuodj8q28lR4Xmlbpbzlf8E4GjTUbWfCuNlIHStkGGGs6bud+ftoA1e
RQdyIFk4O0Tl3LYMGoUjvGtKmV+nMu92Kusj025FBxibuNuE4R3+DsmAiM3vVDON
T/K0Ngm51jOygPtXLHF0aEZrCLFMq8adV4rKEIUbCaghIu9QlbmVeo6q97S9WweC
0jp6EYUsPpPGDjIu08A+8Ni0DXR6gnuCa8ZUXSRb8/Hw16JBbsyDUsaPCidbtx+H
Eli58Rj3fXbTHagfRNOhOez2bSBxEgcdeMwX5IBNdxAz+M+EKJDoYIcLP+ISVsgA
Xs+U2wuZAtvG3AMxeZiI4BvevUQLY87Hyi4TPzXb9PhqJoRdX7nEhs+9l/Sab9lO
qO5pDU0NPJxiaa9siHgHrgBjeB7Zzc8UE4XUpf+VllXXGSxtEsduGAZOFuSiyz0v
1+fiV6f/z0mSYTOFhKFTxB32931KUIe2HT0aYh9eg0Ax6UtwcfKtFfebJBVW25+X
yq2HRcFhkAqkin7lCDR7joegO3iGZ1UUHEgimIfPG2CTIHWJCMm+qKl1Tz24J4CN
6YDbKIzsGmWf4pedjbKMtz58fmmhWwnOK58B+MiSHdu0GMXAOxvNdGXyi0vpmJ0J
aeoeYG3jFUhKY9wtoOQCFCbLPBc1ErgFEinMNz/7zamYWjIvvKImnMo0fbsbhzWk
X7OqVV+PpArPpqiX01XfR0MQ20BpSSgcWnutQX44FHV2jUWxzSAQt2kO+Uic4r7u
VnS1pp1EcLiWCRKHFJxG90uje/kpVPHZHOVFdA0/LUoSRR3dyvF1CoYx72vEP52j
HX8pOXCDEdxMnAWtWKekh+HNrsxyHyQT+zaibvceeniqkirjAXcZh2h+uPf4xc2o
7Fgd8SGXd/QSCeVuI+tY7DGY0dM0R9GQkBZ4jYVdjJ5/f9ADRvS55jnH3SOI0Hcg
C6sb36QR/G7XOyx2+El1i5rfCtBW8s+9/yDDLmYP62L+fdU1x4Jq3U36d0uWH17B
Dlgc2Y4NCSsMuPTU3vWj9RoJlpmxwUOxigX7tIm41W6t6NPtnYfZSrOemXMTGOZa
rHu4dzZ/Dbd9PEIjzVEEkUIPzH/13H6+EM7LV6DF0zml99ocTQerV3qAlhjUF5Ev
p1YbvNz7urHFG3zbxYRLIcCzPempBxlNCSJuzR+oLfYKi+Cg63/osyYKSMHsDkyy
con3X18lCM+++6b6jMcTUb107Ywipi8PNWWGfcnBvvMLdnsddP75VnNe/BYhoyDD
e2DTjWHqFF9KQ3upK8jSJ51mstVoUaJ+rZsQG/wUDyy9EiPYFs1qXOdeQU3S7PcR
bY19kXWBQHOt/iEFX3a5kD5YieqtcplQLNWoDVUWyfbDB+5SFFv1yozJkBTuuWU4
6NpYl+ec/OZ9Q0EvaLd+zusEguE70FY+bNP1m5hG+aQm/kR+zZ6xV5tResG1To+r
tbcX2+h6S6JRMTHltdvtwfuPHKNatxD9gam8UO52chh04W9wILP3ycsIzm8LAH3M
77FbawHdISoz/qLB9JohfoGuCck8cXOIGDu39gWQFdJ8Wx7PXdxlmVFvGKvRe4FD
CqQdtzehIKwodmsSMsygAxwlh6ZzRzKy1d2hm8gYBi1HyVBZ3LVgzBJ7BqOi+4m4
7Z+RxZRGW6ebJ0O/lOtREJDoSlACkEoC+gyfaTfW2g/eLg9iSvP2mT3hCdHaTWQs
hWFneVgVn9qOGiceGPONOFXD0KwMngJEGjFaoP5y0HFZuDdbcPR2N9HmcxsZyviV
c0kFAi76c7Dy1JHiAZ5oBoNrVWUFXfpfS8koyJ8QqoWkEBL3t8gENG97mstpfmNg
TicxJup9bbtEtr4WMj+NJLDPEmWlok6L2+cv4KU+9Ljk70pMR+JwfF/kCSk+7kU7
JEUzuqNQpoNlODiEfKsb/MqSzMFXFsQPpgTdSf1FFtWsGQAL0GQ+tY/sln/TPCzd
XMIdnWgw7jK0Ai/kRc6zotzEyQ5ReghtdGITCYMiYWeJBc3UuBDSobxM6Ae8kXOK
V5pfZDc3ky06GJFqNI8+sfgFx8Yo1qeZPR3f3T6lma8t9nGZsBFmzQlCGY0h5J3g
uOFJsER4LHdnGpSSU2yR/DjEpIP6rWW5W/bNrMp5hyrZ2CnbGjYHK+sJ5acYCd0C
P/nJW4D9OJpontpOh7/GfPPY43hK2jCqb2kEVK3RUFTLqKdEZJxjOk3g9QAuCg4h
jOExwTwLDVb94QYFqJc8c8SRqRVrjm6MuPktq25kZAeGT8GZz5q3limbQZKUCdI0
H2j9OiU71XB1D94a8ztAFq2W7A23/iKlB9U7eMUi9PsHvo1wW0jV4bjfAKHkSWFw
dR57cvWZS2eKet78HM4UDSw0eApmCazXXIaCCzXD8LyttMrRPq7YJVglt24t99AO
Op8MjroO7mo/0f79nhFL6cmKg6rwveGPglsKzINahRaacg2qDPugTG/yuI1Vg4su
avtgRrwj/OSGqtxDfIS4xii5Fi5uiJa+DQ0Jb3s49eKnTm8MU8Un/CcYH6hd7L3P
qy+ejyygGQIIh0tLuYBng8J6PCaEnYgzhh5JwcChy4g14Yyfj064ofhDB9Lqo6KE
mOIosg9j1O/XFAAN2nsosvGpvUfgFmPo0JAAf1aTHmRZAZnDUhODjfI+nAjJBZgh
QoMDsK27TTSu6WJF6AkYHvdEXpYFvhSpWulQdIxHY1uKY1gboXwjn7j2s0Q02iXX
+8EXjhzqyNmLNkbh8e0XU1tKJCYtaYFiallmWI9AO/ScfcH/V2pZtEvkIeb/o7/w
6ISJ/sPINQLP97rygPApHqLMOOVSzF75JPwQG5CfIzcVXbwrmDxhYsatfBFrXaew
aeES6l7eBAUplzuuVCEoEUniemIbj5ebxklY7KJ4fRTBAUihIKc8DyOckn4n29gS
9HRhJbGI3zUVxZu39z9ijl2T/G7tY9YYC9Px0K3FPBG2c4konkA30bJeM8QEr9uY
hcwkZMNGkyJ+yVNwwY28Ce/L1s2MxiMu8OxUTRw3lsTe8Gy3Ipnf2n8fn42oA2yJ
4b/kpA35qcTbmYjlmeizK9/E0XP98PkhwPA4SXPSooZSGTUcv50TqSYVxUjUK3VU
eWFfQKefZQqJBGPoK8lCiyz5JTfFKujCoZGSROLK78kRRJfhpcuz6gV16HHUxkAS
3nxdeHh0fU3Q43iY98utcu9VmCoZosesLiCUoEBdASf0AxveXTQhB4s0/ZS7eMAV
p0QKnMuogMp636nIGLb2HT+lGJPS1RJJBQBzw75k5jlWPS74RKqgCtcboIi1O+hb
ut3AnWQYokK+yp/4laIGNdtQoyq41Dnta6HHjeGugrKOiNtYxAMsi2su1Bn1749N
jii8wiFZapHJYaT75JUva5SI5S1KGuJ/pxsGtJlkmla7iTPcBwskDlv1PA98yDxV
KFl2G3wU0W4updrMXIPg8Ai6MOZC4HILK+zde/xYFqphKoOOWK/OpN6rnwSzsJ8Y
4KU8kRdfoV+HCB0ATQW236n2JE/XH/z4r7a/d8Ke5T9GxYmeA1gvvBQ7ijw/glti
BOwz2VN/IBt2lak17KClPTuXRjt1Go177OJoYXcJE1b2mJmj68VLbQKQDh3Pjpwn
/hR3vRFALFG5S4U9A4/LaoJ8JI7CKKW0U3b96F4sMjZZryCJW7+kcH9AO3jVsW1U
f07fNfgMIkzsgYW9r4WeGqotzBo0nppvXiTnSxNf9W+aigHop5MOP73XisKsh96x
mrbjQ5gaClPCa/IWzEYheWNz5rbtrEnPK2yLTsKvTONhIf2NUUbo+2nL/8IVtAuF
dWjjt7yAqahv+KJ93YDMCVCWbmoATyTzhHvInCFVEZ4TSL+pC0eJUi50WyS7yw54
Ca6x1n95/ZF1sCd4/jHtkB+4SQBUeaRCXYN6sotR2HM6Buken8L/gVbw9nwSp1Xb
4kemeErqE84s4vgbOJiwwiH/U4vSNLzvIYkJrTddh/xIWx7nEvjxe1dKFgwqrXyW
ipGNtAxb3zw8z7+iHOR9RNowTLDjKqck8YzHN2/OfaQSvNhxqcd18i9ImasryKid
r+7hj1D5Vbqw+B9k0IVDJGiLOAkBUaIJZSXJUTQiIXZQi7wd74KvOZANG80gxPuC
tJNnl6fuUJvJ1lQXgiYJs4oIAtpl+c205ht9Qj96sJTEPAl1/NQOPdSNn6P4Fkcp
lGs1hJ6BZfqCIW5vJsVbGox34zGTtVFKmedmrUU3I3wc1DSa74NwnRW6Hq33q/cO
lC2wL00yflCDKn3Bp0plKBajyIFLoR19NqBx0ZmzBV3Somt0D8HhulesTTk4V6oL
0OXU6uXtK3ZVfNUWE9cHoJdpCW9wP/eQ7Hr4GSRSjnDZoe4UNl/90s0QiQ16dpnE
hQdbx/uN17h3VZozqSYoQVyRX1aR1DwM+r5nqYv1czhmAd1KeJx25AkdhUto86HD
2Tatoo0AywNU+unFDKSpplClTiiFjdzcwfVEFmAsPYvxg623ecVyTvtL/bX7Re8r
jsQKnvMmvrrpRzfFbRXXb6ssdykQzS7U2K8OZBvEtbT3mmr0EsV9TxxyZs8PiO8S
K4EGI9QSYI3R9YXSDowcTv6PfgU5VVR2dTpZdPNqef6bPBnj5kLS4ugxiot+IZem
uuyNUWXI1Rc4XzjtlmaF1PVZXUtMh4XCEg8DG9BDGUdgmRnXmCEfllF2olODOAgS
g6VzWDN6Lpov5x/eo0P7/UKUpKzPXHwaC+EsLKGlpMCOAkpWPHakFWpGtZeCQxtX
pwakvmNksTrnHdiQkXSHYbmo/JalYl3z+UjaAkcJ/rY3Z1G4OyJlcsSEFGhr82S/
M6ohCKMM09sr3JidBRm2V+iLRbI0flSywIjML7CVtdJHqCWKJgE4SeGBiHr7nQfG
5QnZVHw4T9qplevpjNz/LQ5AsII8kDwrq9LZjNq6hS1R7HOJjyIIp51PFlrM4ysG
A23cfTOjdt6OL+a662HTVJFmfko2MsDOm5x5rN4tF+FO0v06DOcVAh9R4tT04+lN
Au9wu38v2Y7g/PppeUyeNBaxbsUQTP0H5EKm1HVSFhxEKnwQXXa7ZFC3cojEp1xf
GtBflae894E5CNS4ouvQDvXB4PBMM0UbFcspppqHk6ZlrhUhOhqwMDExgP2JmA95
+OXgC/Awo2DSWorhWVqiIC/hDcnLjMqoR1EbQhOydq0/eFbcpcKFJ6h/TXR1HVNu
T9G915T72m6bLVclMLZDAh53lEJP1rWEuOBxpK0DrJJbPKsi8MwLlD20uFIHQUee
fs/g5mZ7TBCD0BlcImCgpQS8PNmxdqFQA9+5QsJqfDNjrQ1+8F6oywYzsv4cLFVW
lqpFyEPcaF6n5BJiSU98SxhnrC45ocVw1wM9FZ87N3kBhW39rCZiMoCmxpXXAgGm
wfhtyl4KhXKymNq91AL4Rqdfdhu5rRZKVLmyJXkH8Qd5TQ+XFnXfM56Hfm6RG8Ci
prmj5o+ETTJR+N2TjJFupWu8drDXMe61dVmi+AVTccZHCJmTFPViKtGaHBnrttaG
HTbe807eOBCyhyCX5Q3CefyPkiJXe4ww39SCEUSxGjhiemKAB4Hn0Q5JcOFxe7yo
PZur8GcenMpK38VVI2U24syalAS2XVowVTfn6YoOXDJWcK34zKENEKA3LgOjqEPP
/7ON5/60vuP3yxACnk2bdBHbFpge9al+trnTM9/27pCeXYj7UU5DM4q5q2Vh3wwS
bA0Zl8cxUaE2vots4k9uJdJPlZOvWf9uVjPpkjYnkL1H06x2WSCqkgWDfJkV4iOU
dbTWLQpnHwUW7kLu0N6i7s0Ix+YvxVcDM3BpnXRvY72qvNN8WegGjonjA541UYX6
DxbAYr/EbpFoDROnC1RmAdYuG4guBBa9Mbs1m5OW/ZbF8cORvmjllRqWX/mOFK0h
d/BJFPRJzEQ3MdXI6l7GXibnjs448uxqk6dh5RVnZymmG1/IX/bC9EsBU5+n48iI
H5ekeoqRVHQ5gn0XVEyzDCKuvWjCE+j0d3zXH1bZW7ylHCKrYaeZNNCYJD1IZfWu
z6qeWCddkEBH+PQJpdL6cfpBKQLJ5lx/H6Ey5Wz/KBKI9eyv7arnuT3dcpqMdG7x
IOpVEzjLiknIj9H20apVEtGawcQ/7o41RrQe0gSyNW1cunn3FJ8qEQdbLe1TBAH7
fEE14YGE2qOzfiByZaSVWQXhmwzJw3fSabsstr2U0LiUUpfKo7BZHfhSSPsmi3ez
ydTIatoaUppZtS2pEA+KxL9pzFZr4TyhhF9NdAJpbRh3qkyorrGUGwjFGV+tCbjy
tu1Nu+MUyDhfQjQ7QcPSN0sC/RduTRZirPE/HACIoS0C044afDlZmQcj3bWzVrCv
zDmjOqLUvM3od0EX2mLzMKyollk1PdObuxXRWKHfrOmo10EKAqNf20JqoPWiLZyF
RYzPMaPGfgRWEQZ5+Skhrhb8NnGb70ES1JXkdmC7GQGYIPrx+TL485fsODUtshWV
w/eyWDY006NK9Ks3VcMi1fpReOj0DFhgJIe8G08jpoNhQvW+DSxsi4LEonfkJYiP
OQ99/BvEhgztF87Jndp60URVUCAQC9GFH6XkPU//cIG8taXraJmlIUdVjf83rJPE
dh5MC+FUxAZ5ixkxM6+ABV6ym84PPNr9oAsLGzej60y0FkUIp2T/IFYqpl5cXROf
IwpAckfWfU131S0siQcoxk9aedr1Xh4WvP/aCJBC7RfVlqWPvOAdGGETpVUOk3WT
Lhd2Vc32mtAt8Nbv9WdqLKj45v9lYS+ZLpUQMb2yQHn4bl8ZuqC7OEjiWEskllkf
xbX5HLFbp5FgFnBASDqifoO+SaEH7De8wBAnjo6jkHFWmU/u/yVJN9mYZ9z2f+1R
ZQUcge9wtgMTcuhCCJslbU3s3Ghc+U7oj1SlV67pv2a0NubJLc+SGGb1XPSDpOpv
5mpogm7snpCcGwWPiH0zEhNJoIdBKNPMOI2DJ85sIY+kq22eDOhPAH6mmQmxiubK
SMTbvhtjm1Ars/zQG+uOHyryyAz5VS1K5iQ4mLVOiNuvnK8bgzlI69B70jqEZp1I
71Qa6aYjcmbo2FNra6JsqN6PhJBOj62st4Rd/qmlu6bqdjuUERo+gp0eWsPlrAFX
K0VUOipC4OtIGP/8S6CIw92WeFXrmPRwV0Qi5zxXx3th/W1qSjzEwoOtXP8e7Moo
EK4GIlx8OaAQtiTNyhJnjcH1RyHhAXW04pjPQfZpwgRaL3JR74w22AidV9MwzLEf
lRuezQ6w8A5SRUtpfj2WWe2+0+/gC5YJJbis0RsW0FqqXhwsgo/2u32ccSuYbVg+
1q98rOoAFPLWHHkCrB9g2ZlIpoUGukH/8WKXhhMwnPYXBmXQWov9esjxpBkcGDX4
ZOiU77jQAOGboijp8n8uKlJJ4/BfbEnhjtYWdSNv1yBGfRvQm5r/lp6Uiij7hkmB
8O8jdnzeDseurv/NS+S3/x5pdysoqYyNN/sTfC9RE0wQBPPSkToUNhlNyDyLEhWV
XE+K/xbBaGdaBChZYuoKdqfEB9e0hPidd/p4ZxR1qzGq/hmZlTjyGtpIc3ZilBbo
WcCPFYX2aSuIq0ezHOnZJORY/VcuOPfAygBAGQ1im4cTb4WQAl0myhFPfOLAnvmz
Zcgl/C6Iju7nculN7lweZzkEHTFLMBQFoxvgCM97yAmM14hUSblcKrXCutZkGbEY
CL68eZUSd7clpRk3i0lFSwFarfqVmhUD7S5n3yy6dy+PTJSBZytaCtzFKdRSY3Fg
GnxaYEgquEU3tsy/F8CF9DNGLc/XQ8Tn/ONuxd5HTxo28WyAa/mTvyGXkj8MNRow
95vo5kZXVsZ6lDJJ12TTLz7vUOUIrigQN6Q3k/o+s7C1oZjl+M2AxokA79Zr2YVg
j4KKz6nKYvgglaZFFspZ668SyZwz+sajZWPALoIYngrOmqqnW4AG6jAHrBOyjoQ7
N8wxu58ImYVPjeB0okQImsf1RLUXtXw4cLEITBwaOXCXR0mLrtQL9q+eU7E07fZB
g9QNI/XmepYvHL6E+BPpmNTxJzCshuXBku3sgG2ZULWHAvWF47OKxzgZOlrlxfdJ
zvmabEONc1yhNxrdM/ovZg15K+yQY4v8CyAgpNfjLrg3IXQaxCmBiPIuQ5nz8EhE
muPUDJqTwn2H4fRsiV3gLYWI3jTyZXK+xK3sZ5dSOhX8vwiON++kGVtmTGIxYzKZ
nkT3cPSotou2hmvH94rzr6zL1qVzof41uomEncjCUdQJ9A4xMLAg2NufahrLFlhE
V+XQl3vlg9E1oWtHa3Ygjqru1rEOP+9lTK25aF+CZS9WaL9/8A7/jRuAtSc7x8xx
R4gvkx4OyZLPnE6a2m4xT1a8nM1GTLAwlb/nDQcgY7jaK0hhU1A/t9R2yAxfJVtH
i2HXgSj4vJubaMvuJxjSe7AsYGCvjysecTxKvyMHlXk8XAjFSvXYaBR7N8beQEx9
z1XOMJO1i2CDfdq04prvfkMiZtz1riBdGwKOmHYYs3++HKwMKtsPhQdiEIQ7PKxG
A61fsKbf6Ucmqcq1zYj24uZdJt0K5aqsvLvaaUmBVaUSHfFWOtLAQViMYZF92OtC
VhXtkZDYAsLt1GQVTCuvfQcbCj8ov29sWlQ06R8ljx4tQM2EtgjIktRvyXKCdISg
mU+aFHCifxIHfKRe7S8R2Xr8I1iWVZk7u2oBZCFgKncbVBn9I1Gr7nFOqCxixMBB
I1qQZ3UKNETU2YGb/EUV1nDaqSunBgF/Vyjd+I8Wj8uj8BGJwtJ+MohNLMBnEb4Q
eTJ3pkPSQ9PvSU4SgnXU1HsooZUhwqFSx8ZxylBZx/MkmI9dok+TTaXAG8VlSEra
X6gHydaOYQVpiOeivL+m4PTzW4RB6qrwzficGETBMudkvdytE1LkFtctRawVrMnq
ufvglxqyv+i19vNBubMIu7NN6+EtV5IKeb3eZU2QrBeZs/inZbKqH9AfBjQZ3GSI
1sMFcjRDqKZc/VkLayg38J00VJC6VZeRiAU9HLMY1loslbzm2XR+m1arhPWvMHpe
H7deiCSRxnOYcbgFU7HUlTUjutNb/zoBAKuzg3fNz0YFvcAFI/kBMfUt2DeuiU2E
1ZYHhd4V0Gcwsy7ZhTZMjYki+ilR4t+7oz7EVfZqdFkoVVCrBqO6qVKmaEjRXFah
TYVWWKvxQ7xbHPm4g3Oyw4QGvFa/ORRdpBtp9AUTL/1SonuvOrLvCqX2siG0e/kX
7jAIduSc9U8XhEXJuoxpLO/fY/7wOg+PUPlQ50JJ8KITGniIYikQliY9HqjzdJ5q
l8mYf+hbrUob/Wi5UNK4IG9+0NC5TeoWfB9LZqJrLtdN+OeEoi7xMb+zM/M5iuLX
37XWehTQ5RvIbbENBz3mGka5qThlaeWvMgf/04wOVAI94G0ZLzkFhyEG36h1IeoI
+gfSZX/9n8uP8K+PC59woGWdIUN24oMadYkBaVxMFzELxfnLhGtaUO7XHtYwHI+6
XNQP/VwQ8jALcWWsJnsImL2WT1z+Ko66BxRTbIPTl4oDVAjvsas+qfLH/riYHBKo
JKmpWdtX/EWsv9eH+BZBZMOvkcS59rHM7wi1Xb+Yo7xcrFZ61jLlJqKf9C7H0a7w
15yZMi6gxJS7AiRipil/Lq0tV4ZdcoVaMyh0JVGw/5DlrFNFjvQmG7r/IQRTMNr3
fyVdvP0aMw4jpypBDybUN8VOMW8s1OvNKs6dc+oBp6aJCAf7nKEZSJ0cbYU4KHO/
+8byHZN0WMnckSdxRoW5NCclRboZM9LAO4GwjAA3IHlNFAM42RFp/o69aH+co/bR
Z4KBoiTLsJ/oqlA+FCUBXfCsZgyIX+hf+FJPBbg/uuw/hprw4gvoLJGRnhZBklOc
t/oXbsuzziBcBgzDOQlm+hr7K5VXZHB5AGgx8s4EyyAVps9D5YQ8t9xUis8YkjYe
MtVbgxdoOg/3P4jUHXdNEirg4QRg26F/+sbxDU/UuEqb1hoyXcWfYlhIyY0xzyrz
NFn+ryPnH0dik2oXCD1Wc59egCqhNvJdOZ5CbloVKvjzIIb30MszGHReFoEtcKsL
7KO+zGDdGQyNeTtCjcLRtIGG9xqKMuopP14nCqayyv6X/58u1EMiej22VwHPFe+l
SYaUVo00oBifvvxImJVAtZAFv/vdhiihTB1P0aCINhfQAJYZ801gCRHdqqX+YVqS
s6GOfGtk7IBGy+CkRPUoORcuFWazXDFhj8N3W096sg3ADeJp7/bGlaFyqkdniRxw
qJcEDt7T5NtTZt98lMFqjN9j9i4Jqp+QOlLuShPu8pfxbYMmo8onKBqOdTVCZyll
mxuxtxWjM1kptRpnmTVl/DeC2AvbZuwA684BS/g4Z42efgVFueErx1SwvN68Y6Lp
KPP/NPF7Tvey3BnineYvpk51FagrkWUuIAH/w73VbhiBG4iPXpfz47/WLsAL3UUy
51eS4juVi/ar/MKmgLWM3b8JEh7VCPakF07lbyS87zi0OaC/UySdAKPZ7cFFRB8r
ietMqQdEnA3rHp8lhC7g/cF0bEwf6ASh0a9kkyWzZSO1AHDUWjwDPwvGOoP4HptW
tozEyJKQDbhzYU/hTxVkLzsZeWU7IFGd0UwxLfzAmqs6Znt+YvloXFlxFv2FUFFY
8+lfFAsdKvV4UFz59/2zyONTTL8kZs28STo09D1qT5VyAHBq9fHMlWtSGPIg/BlU
wADUwB5qKJx3r0unxH/vfoJ8E0R5vc/yt9QvD6Ead8UipcWIZVuMPBUmNr8tUNfh
UE+CPpQlNG3s4ZeYSVFOtbWDlZOrPtU8WqMtlOgvWb4SmmQb6HZWjMw0yisNtNEu
BuDsnntH5DToLkXtd3yBde1XbWi9U/vI2emUft+tREbMyBAw8UQZuGMNflkz8io3
n/kQ0S1duDvlce4jJIa/LkGIQMX66ULFWi+4e+6YLA8E5Z5MPnFpbC6zgquQ3EXf
pC4U+/HKkAwLDPXZXjfnQLr0d6Vn0WauHgqV3LJ//e5+pYUN9VTmxL0p9tqZTlHM
4HO3ZiGMIiwYpNG0bamnCC9KgFlHRK9Px1CQuLohEYLbWFqU7b55WDmTYVzLetlc
xBGq5B3tmbWTFwpJu1puLgQ2f7zeoO9BxPsdmVwK+rjoDaNjfazKeGYXKLshq3C+
NILF2xivDUiEvjqFZp/gDLPOQyn8pOZ2aSZBsWIDWLf2plBDrpfHWjr6tDrFSr1Z
GZkr0PkltDMUFR9gWsf6qPmjP06aRZOHARMTY7TFqEhCQe6ONZk187aN2R0lJM7R
1JRhquaARqqu8MFGBGVYxRZrYOjjixtzQnrQzb4MDiDZVBs8QVNUY+Lm0QBCHxnt
YLBhQaQiVhs5KbpSjTSafEG4D6tORfG9TE5tH6hxJO0EZdi0OIT89Sg5YnHLjJAv
VAVm0ZDP6KrJxroOWv8nI1oMWTUSVrKrCOxTz8tRkBAZWSoUIDyE73Y+f9fKnK6g
DeEDRFR/FG1ySfQ8EbjNdRrjZDUzJG0x82peGLKi9SRb10GgjVNFyevsEqV9Ndsp
uwYcfNWHnNKJl2xTDbXRb56OQk3Q2yvvJq1ihnYFcNYAwVlUD16+FfdoYpGrD0mC
raChmN/9iHkkvRxkn/6GojX70vjq479G6vLtF4Ih5IkKvg1yEm9kTR8ATjdFvdaB
ApwJr3qcsR948yxdq07eCcwQOtYiE4RFhxlw8x7+7RVbBRam82Q+hJ7iD1ieQw2d
UChkiUr6hD2GLOcsEB24bV8ewwi+MsWiGLTnreqdFSdcss5AzuGUfc+EyvnoEMKa
ENctvH025J3kR2B6yCmwpa7wcyZc/oUqwkwFQ+EwWmVp3ASEKZw2bLoGNB3TOp+C
4Ga7Z71w4IF0kAm1FwZGeKXNRmtP+UK4ZwuSY/G0lCN1rAeZVpTLAiJrYzaMjc5k
AXul8xuPunNMB45U2RIYVzB2HafxZx1Auw+4G6CJOa3KuEVAdpk5LutGeuqBYMcr
XJA5L48z6fKB0A2FuLCxtf/LufxL/U41qnDfzD+Pi65OsupsZD8sxqMClLWcvjpM
h+Mw5NxCtiK2WJ2wKCStFyVywlYRseYO4kZ94NFR/g07kjdvPGYAG5HJn4aaBLAP
IFb44NKJtwFwTsRJcgSw46Nb4tOKFee+w1iLwccPB4llweH+x4kvj6YbaPeoYKki
wLPOuoZF28EDZ7W3+CTRhD7hBNueAfPOMv3yT5OuSMAoZG01O6rGql032VrDs3sQ
5efIxin4elnu4FnTAGe1amicUwjpfm/RaqdFsQ1CsrFQ7h3G9IDhFLfUk7TaFezC
V9hxCxbzGiRmwPgKWww/DvQRdW/h1dfcWJgdK8YobOmsk1Tlp5KDQ1m0j7ADW9vH
ZVDo5zyKzv6sWmnqk60htt2okABjtTiNDWFE64LFdXMM9MYj474rvW8+7cOCw0Xw
lPPxSQCGIns4n2vXcOw80KrdqgOA0UXyz1CbSPrpcvb/80wiHr1frgsjBRBQcXE2
Z3l+hRaFei5uRfcwKzB4Jn3T9KYI9Du/i7gxKTnKktqE7y4fcENN7GsOZWTt+4Xp
cdTTsFbkEDDgPKxkmCTOhTkRfhhOQ6hI24DToKLxSoSBNGmEu/dEkr/NaVRwEq0F
qbtpRBqRuKRTBdyo4jNRCt6SAqa7sWYLNym+MaYU9h6I4jHfQH/sfXT0Inx0kw2p
aiNOq+wmbL/l9F0wCsPj1/Px9M1diKU5dIUg3i5YCf/E7NXP1Arx+pLhis6cW8pa
RmOyuR6X7z6Q5zoF+vNDU8bzrPiKJt8DvWwcErjNCZ1X8RgCOFDBo5adLxNy8drW
NWbb3rtNLr+s03WcwkatGWabhsw248YiNBneV8Y+h5SW7YOiJNc69eEpSDXvI8Ro
GaayjnwK+ENedNK62Ex0e0d8FhLSsr0RA05Dzpy/E04bvxZF/Q1mMaXmUQ+VJ/5p
CU72LSN42LGG9v84kSgDqlH1h2M1IehE2xXp5H3llN/O0SVLMdp6q1lUBmbAXd3e
zPzvhh3DkumfTrl9PTNA/pGf5kUe1H/cpTV/9RAmRoJE/bOxuG3AbpyxRpb63g4u
zadL6pO8luuXv7YAj9H4Hh4D12fdOoeXcnfxvNpZbK97KQisPyD7BYg3G1lAElxs
HnXm4Mromx1k5EeCvP+MPPKedjHGqffNX30aIUWiJE1ZoR2YwgQkrwt43eZwHlgh
4SR4j+FBwhwnruFYiAM4n7AhlUDmTznnpQyfC4D/yPp4cFiEzeNl5ed3TAzQYNE2
FO//Sch2zv/Rl2j/gGBSuno31BCFfh3MG8IMsWrJsHk4I+glQ6cPGWI0kEILRyhk
hMQ/SwS1SPQy6EDnhFKOjgG+Okc1rad+dL5VPEJhmqznz2GAby8de4JXM4rcxJnu
wCiuK1xrfqSyqjpXB/IFmtED9a0bjyH6spXhtOahsQhCwnaPEgAlMG7tIPS3U/F9
i53Cm9CiuCKUihtUtnUSCvBXXKre1boLaeJ2hKlqiNsh2ma2FhchUmmSkNdwMseD
buc3uQiyAkqAGibKyTuf2JVE/CbRA2UoriMQiRFytHTb70tXVoDhrio8R9SYrVBF
II/K3sXh+zeS08ubhbwB2io09WP9t6xQgOkGdWGdxx6IQAGX9GSZ7N30nSNKanP5
vntNS29NHW9m1Oq/qJK9KKFzSXVlJ9EF526z3Q2qkf4miBRVShDvs2n9ViTTZO+7
y5/eCC/HFbJ5LRo1JVQgtp0PHKEJpQfufLzGBXZhnM8oRNTiMaWfojvWwch64zpp
Mvoav+Gxzo/LhYZ03TbcrpcBGto+4Sq3Dgdneg5Xj289VSMeMHwctzkTOovcBb0m
nVqQ1yuwN01yyPUVPUMLzOFObRtuWcmYY5oXdRCWNLDJ/Newb3vkJiE1TJmgDHf7
D+VPk3MV4Mr860z9HWgk/E/+TAhXeCiGkLfgbWkp+mslXWcF+kcWvPuyRQGRPKqZ
ykSsuugIVs64OzrkCyanrsQMWvf24B+DPnugNbn+1/1sqP8xMBl8WO5bvYZDSBga
VZXQ0LHMDONIT2bfTGuLHdVGEZ6mLJ4ZXLl/DVrJxjVi3svA6tIlrRpIqIOY5RdL
GZJPrdoRuGLahMY5BdRErnai8Ua3i0exA0VwGsJtpZlrEFEnWWNYhMHM5qO5tB7m
qXWtDaq2eTA6IfYD+KTRYfJ+in1pExEJRJ1y3jR8VXTo4LRWRRWEnbei64R/9GkN
cj4OSOphgErhywNHbU69vOsFshORveodY396PtGeP/wwRKuAmasWOdCh/JBya83/
i56SPiRdza15sy6x8zxcZTWyWLdt8t8+PuNZ9iyB+UfXeJiX0z52BRB57Fz6yaYf
kPD+1S/mmB5RNaCFXEKj+KTkpjgVhKqltulNoyGZJrFilkgVbMR+DkbHcF1Syi9B
+xe3iN3NZiPpEf/nXmXG1Ky3iYcxF/XjOfbu6l0VzNHrEJ0vrE60tcDdOVTiB4pc
ZyFIL4z/rGr0sn7H+ej/OejlHdvB5ozLDK3uX6Otm+b8oz1SYHvImUlNtnmcJ0zY
j8HARiH3QhaG/jYcMHLXSuURsYj6cwrDDegCcNdMKqmuZqcF8rQhk89mRdLP9/DF
fpzhZ5Z41iufnZVGg9SmCeYPqkx7UeggRB/qD/FafLcr9t+799S9EK6eI5lWtgvG
L8/2IZEB+HQGvoFJBE77d2LiQI4xZmgs4trO4j+Kp4tqMGOHO6Ypy4mRPhTA0Goz
KUrJ4mCcOGruNh9s5FV2Bcp3VVAg7tPP9yA5JQ3WL0U22YB02q/txABT0aHdx51x
gysUB++EqNiZDskDgCe0wXAAuTQP8vnZ5OkC5HSehgHHA2epULz50Umo2Gg6gqtm
YAgjnUsTo3+TipbwpFRqE2GuQZ17gvhzdnNUJ6Nq/GcqWD0UbhLN7AkgH/8H5cat
ZfDvcXrr1OnwDjflEO1DrxT4gXW7AK0v0WWzwh741uTZNNR16AzRoZidhks1vx03
swgVXwDWm/sVXZQGw6pv/h/5Gp4hiyfqjZfddpX/RVCLo17/p6jK8JtK269DvWrE
msSRZl60jD7PAEJD9av2QoLGL0WGlHQr2sJGpHkr+j5ZOCgZvOsmLzhB1Gi6XPKH
Hu+gL1uX/MhSriy7M01NIX6t4eTc58kWfZkhc32B2TCHUvB2Xq3xVnY2pUB7UxsF
rIrzQJ/A2prZu1KaGT+mDKiOXpwdXfG3zguiLtU+0KaeJLYKDgBxZ7YebatzPeWa
KgkNsX4WK9Z5uJ5zEwv8YNadTL9jUFHGJgNZ6Frnu8fey0oVxvMn0PHge5GofQa6
zgU/qA3X4vJofYIyX3Xi56ACZypeKWvvuquUE4yQwMky38ehsM0MtqgOeYl6E7qd
6WGzA8EZ/eAJm7flPBanNZ+kALPn+9O+PTLOchTVaxhQeaUrpNqHT+n+7OWRhMFE
keH7Z3+Roe+++XdHNtJGeLk1O6h9ohoByk8H6Poasn54Qs3A8B/JyigF7f2rFBAW
VgAQzlsELoTLhXQPMDFIZa+ZL7FBplzBKNcpM1eCI4ZjC8Moc4LVEHz8B4jkzOxr
FdlfPjpCQANSKZmBVsvpYb0x+nqHdmtnwIP51ADTYB3x3d3bHe6dlbyowmhbfonO
Xv/gkuZ9/4o3uf7vLCFRMQVWKActOwYvQdlhPjX0kZQmtIa2vWFW9QDi8AuZmNhu
nhAWl9RaKU7ZQWFZUdsTn5gHN2GXO47wTJwS60FsZMVCBXBcfWNtDd5muA9UrNhV
mfHtmfmMV5Z57cGh2rG9OXtPNIWWZzq/gvA64RXE4S0i4r1hWiVwzjnM4vcoA+h2
fq3EJFzg4NJuJ55rZEG9QidmdsDfPch5fSlAR3z5VcEFCYDITLmXuPm5AI+twhUg
AuNMkBQEaP1DOB/qOQ/W30R0nUdtf7R8E7t/5/+1EC7OVGmQ6jL2mWU6UCE7xbHO
BCP5Rv+gBgpo5RzmlTt5iGH2ftqPRIMKQrSfsJlKmQniOCbzwYvxAKOlD6miMzEj
o+hkQxImC9SLf5dtok+1HO0f+yGMgnmmlUby1U2VpfvZdr6QccAznBmXu2IPgcRL
PZPyP0wGI2yFZbxTh1Zux7hh0XaIE0t1LQ613DIdvofRORIwFf+HVONQ0HoF7bpZ
8V1L1PxOsKgGA9mYc42j7I9CpdwuKlSK9ETmvkA1iHMuHFuO0eHFEUByxlXC/k4Y
KUlmElh+gXoZY42up/5D5L4qyoh88xX/dKV/bHwFryfqQykAfCGxJ/UJKV3d6M6t
o5LqV0hCG8up+9Xja7lzT4KdqLexP+QcFq1XfKM6N3HLp6YqgaJXmatdHB44J0kq
XrEHy/MZJc0KL4Z4BxhHzbWBKcen4QyLto+7ibUFe3haT2G1NaHYdZKBGIQSKpF5
Mb/nvYN2QhG9msJDFhx3nangJdh3GOrJTeKmA9oC03Fc2GD+0gDcVSB71WvjMSWm
coUr0me7V16dhkHHgOXp2QbYICQtPWHzGHWAFSDjjaIygHcBg+R2t8LWXruExNg1
hFcNGL471PHELNE9XpBnOTkYTVyTcZttLpISZ0pbFQHK8K8spIatiDrwRHv0OPHm
tWIfZwB5ApzHclPQjpuB4G3hEQD3B/N4J5XRHaQQBxV4BLOX2DLwjHTpOeqnsyxR
mhKIN1hdJH81OtRu2ZpBYaPMLwmlLq0q6WAS2O/IZV8WNFr6exB45tUDb+wG4F15
fPpFNPr1g6eul3Dj82Q/hPZ/N297Yl+b/jkpNzCzykCvhca13BdY5iIyJsCTMq7q
LI6i9/r6YwUHJypplU2grAsv/p9RxIFRdIjbg49n2IklwBD/4BBbZbSzbzAgPdpz
QTJyLGSZqPts+LOxMxt5+azJGDQObAa7+Sg3gZB76AKRRzXURY5c1dd/wlqXl2Da
JprzDugAuI95I/AZqnlOHWRTvbn1Jsg41bJjTCdAK73gq8axsxF4zs5Jr3ME2eRz
O8Fkkt4oAKioGvfBJ+Nn+c94mzU9piCfsOgoEYp/y0rDn8Y/96KXH8Ocvji3dEr0
y27HLlpkH08+d2kHvGCl7SmzfAFXPB1hUYYVdspYqLjsLGSip9tOe2PTExDfTTO6
yUB/R/jlAE5Ya8gYhlY686CyKsJv3vZ8ZI62ySV1KB2oTWvFTjtzhuOQuxdK580+
YGApqj4Tl4xe2b3GMA4kTE01uJOs3fS3MTz4bnsZlTlZmsxerkxF2AEFYEj7mfsS
nNXmHNYaK1F1lXp45hl4yvlKUDamtPmBhohz8BFrir9WZEGH5+NLbwRJfD4sxO27
ZdESNG+6WJDccf3PPXtqgHJx1t/wdVXDXtTWF6nb0km5w/wap6kkIcMQ4yk4nRa5
DtHsU6VfCz6WCA4T9aDjQAn0YNV0T2ebW9Io3aAcOzDjdAtiTJdOO2KdF68NWI2y
Yn0WsSedpbcFUCdphaWf6KMvn2eCvBfhR76UTef2FY0HReHkNYWdsps261s94PMJ
c3Nl5F5KRPd6DUn9KYQDIV6Yoop+UiK3X8Y+yKChlGdMUpNqnb5qzBkT/YZnEu94
Cci5bw5uBw9KM6tf6rLGBrcF7bYfmh6e4bYfVhoc78kFS22LOiylTJhS3ckY5v6G
KMBF7V6hkqC5od2emmXj14hEeTdC+3G8Q/9s4+MbCP11giTZKVx98fIRsc1SB39Z
l4f79Ry5imQi2BtCXZmAFweGUJQnanzVVYW63TXvZ0ZoLjJP+ZoEQUVe9BBonHje
Dmhney41N+bJvA4nJKd7E2mpi14bHr+BoZM2ltFxovKpp8wxuju/6b7qfc4uZaSK
RI8re+B6L4TvfDXctiUMs4sVv/LFg3wHQdhRqySbS1oZtgQSDVWCi1MX3/foz9lN
/AzYBuo6p++CwxTaEkasen2VzrsBw7u1GsApkk64kFEbeB774TsLEIEI28RcLb2I
M7QHV2Jrm4Ulq/Ut4p3SfyDSev3N9GmmlTaGjdBIo63li+52OpbvauUWbPyTP5yU
0nHzYZVRgg86+zY9YGKarzgaamkJKo3uzPd8II6OZHXtkHn+5sZI610MQU6naR3b
GNR5k8yCYR37viHUjuitJTPCgFCEf5JdA1D4JwyZaVzWBTzCHkjz9VRxnM6lxkyT
uYcBOP3AhEYeGBxFH76brSqVS7RMAfSrGgfkFLAd7jS6AaaYjBVUIxPuGDO6glo2
VaGahI1aZqdH6LxFS8O0S1wPNEHi/AD0g2GIrDWj32NvqFMw+6KuqTWf6kJF3z0Z
yi7SLDPSwzGh0egtFAw/KUzKa84YaGiWXQd1942itEhWY6GbtWsC8k3vDw8AGmLm
NkSVgXxr/iViEkjhLv2RrPPAmwxK7tGm+nsLQCPzoboaZoVRtp+4y6GTmrLPGvpH
650jRxloM4+D25D0BRip0OaQmRvmoGVR3DIIvN0uZ2cPWmjQLzpBIc/G4l3f3ls3
hH6n++D9qK8DHR1E2sQLLhJECC4pW3SH3uJqg9KN7j1Lpnjwb4weaQ4EWWho+hGy
qGK9kwZlVVjMWMCnJpYfFrlbhGogbvfFW4bMIdznDQ1oNZXfEMcpgh4zO96KLvm3
jmAT8c8AR17Hb6fqrQ7/lSMC3VgDHZgB6qrB69iIaAfwunLmR1qXO4L5++Z9lY0U
v5IpA6vnJYr4nEPNgl3lAyaICXDSzCJsfa8Dm9+sHuUJHCqWL8semRIwEIuqhwdS
pbzjQgNLfyzPiQxdJUaul4cS2du1gnffwBuW1IsjhoYx3+ZppbyNvqo5AWG0xSRa
BcvA3CBZnOxQsDwoPQlvTLNEZn4gNQQ7tXJVAiWz079bOTzPSnr3tyFh0v7PoOqp
hqjYVR43aDAEpUaPMzZ0A6/HfEuYAPejdWXhO0DVCWAJOByhoA2mfkYY6CFC+tMf
FCRVWyzkiowhoNYlkw9JM1QsaKcGuNsd9ZA1GQFmGYZcirMvx7fFGC62xtr6180i
JvNJmSMe8MzuSw2v5V546JY5L6s2F9/HQZTG+JYwYpLNlNmHvCRumnBkl0B+4l8U
cU4qBCQexf8WZyGIEXiZQ1jFWsXIvoR0/Hu+UuSHgYu6MnQjevITSzXb4hHt2/vo
5rh4J9vAwbAricdHO3YVJOeNHx+JSKjC/QAg1N7m1PrDvfQCLZLfWIf85MZl08+5
wRkORgNTFzFoOpfrfjSDa+qIbqGyvtDYKgNUjdb8MmXO+N/JSxodfPvg+6RFuoNc
hACV+sRxhsYMzNp9CPywd5mIwuq2FymUWwvKjl+D+6KMBb/VPFXDpYuyb3/qdikn
q/tpjganzYmTXm+QCcv1RNrIu8cW+pmukWF67lrBW3KehrEC9epGFWwtt6Skx+4R
rG/tdKbxKt0vYZLOL6vScKZ7FoPCwPFou8f5Aw0ixnmiVQxPRSLCOLYxQURFpyqd
NHhf8kC6K3v0A2Er7aZg/O12xMD5g6qeQ4ORn3KA63xWaHAPZlUdnszGJ3g/+rRw
KAUXhFzgSB/QSGqo85GWjiNwX+W9WODW9QdTmTca4BujcxEW7m+dsvT00imiyNQC
py5BZuJLKh8oLmPuX2hx3NM5n1+hhCgy7u1s9de7EVO2zPbCRGAFd8i8uxZdf9N1
FEJM7XxTNtxPigbbEwzZFGQpDvE2sLznXZBQzMRpTQe64cCkSz2B1mUt3i80ZlmP
Zq2k7i/r509PbfP3f7IryRomQ550bDoKOaScRr8fqj2kVu6bX+xCuNnLEh09Cn1/
dqKAf2VAsQOcud1wa1q6k0T4JTAjERRmQX0D6/F6yyh/WDt7GpGSoOw5uRuzQQbA
AHNY2OcQRjAlP7ZRu9ERZQm/PMHnuhTpcOzZ+vrTVALlTTp2VDtD3OUG79Hkof6F
VNWsyF857tp12Efg5Ey36NosIqLudJp8Zj9cgMc/vB6xLbzbegsMMXqSICVhdSt6
3X1PRL0+wNioNN9d5aDEH1gR+9Dm3nodtPx5db3IfY6BB7G40XElo47ecRuO/NFS
FdBwdB9ioSDgwgMQldy8KEVMqII0RmFCMvU+PH1xEdGwnDR4wwZgU/tvsrrWmczl
/sZyy5Ve/otd/E5s2U22nGBURKuIE9PyEJx0TEUWsBjyvXRtOxFhYupmNOzs5l9Z
INXPe2pi+TNBhfYEICuZSwUxBxOxF+2lb79z53EKKbvRJLEAlpfSFZdXMZX5l/xK
wf/VLnDzimOvAswtvqFV2ftiENeWCA+YxncQ/PbkFnnCm+4QjBXaKljXkDblaUBk
Pz8gz/IS7tsgpjhN/UbfTSdrjvHc3XGQLRHciAG1kJmGdkOhw4M0mj1d760JHkvi
YDBhO71m7ipWMIKPkjyzlNKhO3nTD4LwMLpOgInVKIzCaESZUQ+NH1DXFzmMweL0
BYwuFq3BPyctCiNJrMaAXrekKb/NJsz7+ypSUHCfQWkVLUOL2uHQNOUm345z9rlW
coreLWjkEtqSh4zz0OTarHIoAEX8Va4Mz6q5EfgzGT5wUwMtn0UOwaGUWp7J/Qoq
+TG2XPIPgcoDpT+QI+RzFE2bb4NgO7MCYoLWaqC4VLuCtjNWigqJxW86e1CHM4S1
R/64F6C+7BzGuarkV2YgN7QFq4ZEL/tzhVTYuKWerbSFwAxGQFh6nVaCrh7RV2Rr
YDgh/0Vy99SaCUKHcqmWcFqUo1a2gyk6Ek7cmD/eJ3TzCDjThR3+KgZoH7qkLu8B
amY78+YxPAL+Deoq66v3moOYdzMVdukrKWuCGghq96+G4RtKY/f8eWooldM0SPDI
4CieG37PJPkwY2/7xht2XLTv4tBelMJqQQTCHA+srW2w9pDod8Kxg4VwJA0sTRIw
Zxndab74CVjRyqQ43ujHNPalOt3m/uUngjmSV9cM4J13CtT6V4OP3r65h1WxfDlz
PfljsWsgm9V0mJF0Qj6DU5FAAKoCTFgGkAuhcCWJFUWSzSHHE2kgT2wmsL0zDYw6
Du4hAUrLa4Zq3fXC5vkcl+RKA1+aUX5qn6QReeKk92LoWRVE/SOB/b9UQyoz5/Ce
R/mY3t96cwxiYkjlz9R2VKmARYOH6f+ara0lARq79iuI2r2Eiu06P6vZ7t8RIAgB
8Na4oxZ+IVK0OY0b2a3I7pXfcnryiSw81NAE++BJOYtVoZJvOxyG82ErCW5nB6N/
HGoqV448a2HBJSUSeNUHzt2EVN6amzncqqT0XAW0TAor/TFiBfKPfp9fZGALV30/
9UqhfQbaHQPUscNWq/4s4ULcWhGpGDyS75y34VcKrCsNcB1ql03AzSGy2l6d8C4Q
6mvw21WY4gKfW3AUGQZiMuC8SkEkfk5KXBf1I2BurJzi6o9GSTfuINRV8C1wGuCZ
zHeeiVW17QccD7ny/FYpAnpUsMDFkaz0tXDOWtKvH7iW7tIggAka/YmnMIRZl8tG
KWKXEUNcX4uohdHZhkUyi/f5ZvIlFT9iIEUhoeejfVa97a0P4ey9TMP2RKnE4MlS
LSpw2rAZFuG8YyeLWsYomiUEebshJgS6wviTFySY+5JiIM0gAdZq0ifYZX1RmeiU
LxZLVnG4V58Gukf9+xMQhRR/nGW1QPiFau/p2P86TPLgCqy9DYEYZGgd4KdUjacj
YW8LcnxD6aC+7n4EPCsZwzSUOGG9GTeWM8OM8KPf8Ut2qPfnHwXniw0QKKrC04yg
7ByvTZsLpahoI0Ru3E6lZC97SP9rRXytA0cQxeYcCbpz0jh/ZJp8RHSuvG8EZhhB
j5/QJK8VUlRnxz7RkRyd0EIAHYGxp/JIeOGxdeIdIAyJZ5DkRZ+Vb5iVcs5orZlm
2+zMymZPBAD5dS35hxoYuapvbMG9ds96/t5GIwAc21ohw8OijJr+f4T5HdmpFuh5
nNgwtjIJrH/AgfAceFK7x+oMW9BfRg7kthI/AlinHgdr473yWy9LLXFMuTyL7R9f
NU/KgrNmiq7epSQfC1lISnLekodu0q9nqXMz6i7neZHPFD4mWwyWxswukRjknk1s
ZrxDCNLQwuX6ghA4UK6YXIQ63IdWqqOLnp657oObjJ8F3c0NKQUZi6MUA9S8c7t/
c2yQKFiRy7HWqNlHNx5gPi8besnSZmiATqfMjEzhuan9lIsRCywAXKhkj9Su1foz
CPgVO6plCCpC9U6aDrmEgbVa0Dpz8Ox5oxJu2b9JK3hEZ0zHs17g/Sg5U5cOp/I3
aAOzByxf8tlXBAuiYOog3zrm8nzkzEiPqfNyXx06J+Oo1Wfd5/K9WK0TFWTADGkC
uiXKjhfrtm1AdhjvqYJGUnQntXhu5X7/bk5NUE7mwUzeoXUgwtqnsMIjW2aFBJ8l
UfzDHIB+0Rv0S4/eByMAjW0ZQG8sDidGjapaCruC4cnrU7UIPQCUBj3sKDuA//YK
es3fwJHjQX9tjOQQ6lSvBZfayoZi6S+BnbQaGEzI02VbdVoJLdV5ofM4UEffcksZ
R7gZysjS1fnWqIOujurVWKnSBGQD+3cJBvrINKYBflYbLMsNGFdbzgIhBftWgnW3
impCjfwr99QblmLWd+CTtTyKbEp//xNajAeC3+vL7AhoNdov/N+ZO/iaYg5ZtLW2
mEpF8bbg7XUlhxfM1THhOk/qiHdX81fl9/8kA/1C1Nfv1D8V9iVKmeoWlMPQ/Yge
AKnhXxFF1DMuM/VQsXc2jf1Aq64fe7pbnGx+FrNK2taMDf3MB6iHN2wUfyn6I8yo
lpyYzXwhtKDVwEELeqXdtYfjlQtPZv28TYSCBSzMgb9IS6uv0w0YCHB5/Ht740wf
B+/Eo76sLn8esDDsExVGahuvf/M3M4+IYmalay2XW6vimqQS1yqKWeF2Uy8cx+Et
o9uMO6egtfyFLIq8TGRawkk4z15+g/zNdyLywTUEpAYiELnw0FN4dZP1qRwQLl6d
zwp9POQ7TIo6AB4QcsYSOK5Z0wd9ZFdCoxPP68+yPa05aCv5+NdtYv8p1LxqLnLO
VXFcLOKFhabVQT19R0OR4mGoMgxsvEdUoAd7dbpkBENGgEbUoVHt4skzOebeumif
ToKGcqdCuLpLCIvxSNN5Ckz361DCXyz/Vxvr90WF5cWYOQXxZ7tmB2w0yW9KYRet
DR/d+ERwKB6loCAWaefF8FPAym0voglvHUTprWTJziC11gRYOZtCobhcsT2Yh7XQ
ZQurJ5KXgWwgjG1cu7s/ysOBwUxvsjpB4kSXFvJHnxB5PiykeHFnyOoDVqB/bcqe
a/9YIKkGNt+AnqMAnXuZdkXWgVNWLKW6lnQJCqFszowICxPFAN31moO5AD2OriT2
JDo8bG0j+q2/x13M7FGuNLPNm8F1XBFK1SDACnuNesOPJxoWQ1hAKChXCuVVhrn4
RmEoOnnULMFE61Nbm6rmwJG8aXA5CxHAivo6rz+5UIYwNkR+/UjuygUmBXL4Lgyo
7rzyRla4ez7XP/ozG5K/LNHRVGFTe7igtoI7lQb3YYyn3csAzTQbxHxoBwEl+KGG
mz1uY2rayFnjVihBeaHVC6G63KQ26/aXQfOl3qfejHtuekiEzvJmiIaIqKyyYWyy
+vMk/j+qw8LmzStBsqggKHrgwO4YjST2uEohOsznJtO7zG0MWG/lwvCaGItTljC1
9e/jIqYrBBt+R9YuD7jfR4GpWm2XymPU/x/90UbF+FWCbDTLsCkG3qIuHlMBtEfS
5dLmcTIQanvm+KD+wrvFIxIdys3epFopq8kg6ictDx/3BDxC5HvebekJy56JvnEp
sTdZgOq1p+jpwAMNTul9K6MODCDaWN1QxITE1qIPbBIrMyAwRsaNywkjhlz+YrwP
R0B+1RCvp+kBSFBTSHry+9kGM3MS47ccTc5YtRwN2VrKnro+kfTB3iygmDL2SaZh
DjTWCNDoChoskO1ssDiLZudzpJHonYH82r7XLesxQGqPyWteVCc8Ct3PhQoO4Mr1
WUuhJ0PLL3A/raxNUZODJQJIVLdcj2P3UH52srDjHjF86EgVVvZr0xgCuIohnKt7
ztUbUPhla5cDLsVZO7Jc4vWSmFoU3/0HFdMjByk6w1RqmbeBeQwQQIDQqYDgCbnD
0Q9UdP8Z81vUJ5pcReP6HtroCJfktMzEHlzJtgZjPDRq6KUxpEAaL/wWdhsgvuAz
CkJQVJWOlvZ7sbmf+k/bJRBhXyiHjByK+WBfRAEVj8VpdZfKagZCMOReVDjgowMH
aGFXouokSEQDUkdT+J9/GrWv931Z16ZJUHxnivhL0MLE8uy+kd5tRxLKYkYzio9w
URH2VJO6oNRi+ja/MNeG7bLkXVyT618dv/WvbVlOOuMcMbXOsz+NQkyC6m9HuBef
YiqTxaE3T8UKkROZItEoNx1jjyGSyxwZeeFPj3qul7rklHsoWjTJo2VWGMcBS0nZ
18jFAWqp9xWFqutNoQqbQCy8mock9rhTdo0sE9M1yEvSLlEPwoh3WumQ72+UQz/U
PTdys3fggvE0X/rV5FVIvCS0GJ02A3gWqkyT4jC50J6O/TMxANBmLnXAutkAAnvA
DBQFeCQsnHlmAVmvrVOL/61wGYM/f27BNchLmA9ofWcoWefeS8ygkF1T0J35OaHE
0wWWvNVHIfoP1lqWStcnHTCe+/zoyA7lEcg4G2cSTDkZ3t5hEG72qAkljjZLXpoA
RI3V17Q22iMgIaOiwQxmOTSMmBkUhMTWYYTzJ5Bs0KaKlZ12PXRAEnAxv8Y28fxI
7hxSlfYDv13XZxFPet9CgBPosypIvFLrMBY8bq3FuJJiMeHgxVsnhpYgrAWIOv2f
mblCX2SoflgA2y09r0hQiRNf4fjJXE+lWNC28B4W6aQgZMR8W+KZrk/RqeyAojGs
Tev3E+9D2sXLqtwjaIrSlT9dtuPBQzdxBluYsF6YJrfl/pubvA6oK/s7u/rKyWZg
KMUu8OQGoM7FhHE71oJIbmuEMvSDlrmWJ8ynago2MzqUNJYohx3uZM8LwZeU51Qp
/VtZ8rJB75XBL0jQAWuNUc1zxuod/D+oGGO2YrfGvmW+TFSIX48g73xVoqVyGiGP
L/12SpdePFGpb/NOhGlYlDwVz95gK6bvZ9G5aUFH40UHpzg5DhpfzUu/0v5ZZmsM
STRoNkGX4OKb/iAMJEv4mL8HELhyIqG0yXoZmhJmqexmxmI+1fEnJJ5RT1M81Di0
OcsHftQz+5LjjEd5tMufrnyl3bg3rE5mW7Xt0TW69LA9ig48mJ5p/rlLTE83/A7s
md9K/YdAQ174RPG89pFWtE+88lQYLfZ+UTkrQlMPLruL4kHSMDwdJou+u4yNinl9
0e3C8KAkUUdGt83rilIKg48a69BhOHjzUoLvQGXs9wFCbVyXbhd+SQWltdssUIMx
tZpiKLJIpDmEF2eQa7IB6tth8nhZSjDNa85iWtKRAA02orUz2rjO80fN8LmM5UDg
nDAZ6kZK3tuN5Vxa/KOg4ZCdy/L/Pm9hJ8N2WorI0tbDUVOzSYwT0Uuej69zCDch
ldXsUf89Fuzr42pea/Dz9hdCVk6ymD9+cWxAXyou2n0/5BxTNXsuT6muXbG8GeMG
Gx+4Zu3SYg/kAG6xJTbD8RWcbxJHIE83d3+TTpxFlHqIzFDrQXzH65oLzLmo3D5n
6vBg2OlZwrmtWMy7/MWleVtNbrs98jeyIgh/b7IBtza0gztf9isWR3R4kdiB7gEr
up7r0j7U25eB4HRHo4WRIv6GQaLAPRXlRVaBfgu94jZoyhCKQzTWv1rsHuo47CUb
8th4X/6toKx0pFAhVrJjCEl7GNSV8mJKjcRzbhKqYI/9Dj5feM1wECgMu8Em6lVy
ka3aY8nzGCxrmZWc2/hZE8MLgi2gg/1OFk+wv0w5xcKU/l9m1+6XOEnYw/apRG6D
4d7ASpT124Q/2eHmK3aAoYrngfN4FjL2veL3QH+2ZWliObcqMEyd07rRzm+rs2Q5
ADL5/3YdokXL2ejibbDcH5FPpQ6exYAwOdZuVUOdI7I5LpLfa1EM4L8rcdEbpNzI
ftN+JchoRUTSAJZhPvd3ITkmAV51OZ6TLmUX154gFplym1ilyv7Y4o+3ariEZP38
C+wtVzKh8ltcsP+iB0T2e+Kk1h5rH6UQ7mV/rkJXpkQlCUov6u8MgR/BEe+thhfc
VTTy27EvK715d2YewnjtoJlFJDWeJUxww6bBUTlEKq1Kcj+nBaaRCnAq71QTAo9x
jd71GzD/TaSoGDLg7b1+fiQ0gJvIcx7/D12+nG7Kwoo7ZFv0POcQUfRvKGqJwd25
edgqTaB4oixKvdRgU13YdjZmoH/oj+QFIKc7G9dvdMMgHHo/xset1OXo1pLrfBXD
AfaAM1hEhjpY2M+4VVAH3ynVFGnWQ8B0ps/z3s3YfLDEJez82TPaHvHu/qayU4iG
l1qQDIHNxK1RmR3/FcDFLmEgDpQK5JlB7STGpm04sRkM4WUA2PGI0xwH91FeQOT6
OCMaXOPd98gEwyYm7qBBVdKMYIgD7L5RwGpmz8tercDISoYBKdDx4BnMw4ODjgBs
W+BfyeRgsOcfMjhu9BFr2QL9t4VMLfBEns5JFycxzMOHnVXj31IRqgnSNQXOnpxl
CHZ8ou04ygf+4bwnDWj1amxl7PEw854vdoNRewJ2swG2lqnymYrqRqgOzQUOXmQl
Haq4mBQ4/qefsd1125MF+kGOjPydN6jMylMWh9wn1685uP9JLTSt2lbNH3BOElwg
mBEEwc9eBDTweG9r+8TKmwRG9BV68qH+3gweDwmmidQt9kdE6XR9DoALTFehW1Vy
sB8plERzpCTHreGa6krOiQvo/G6QXFhq/1JIEpV4Mv2TmXASwfJjYrGXJ2/3q4nP
1SznSXcdLPNA0pU71+AQcfIodXF+810lpVaPwgpTbkOYFFc9+XysWRbSPxAovG9P
nimHC4wHeZ/7WK0ZtbleSfbUAhHBd0p/e+kdzOhYpGtt5TN4IaNxhoKIK/5ICxGQ
23JwTEpzdyxNGj4TyZFQRYo9TYUndA74uJZ/gFi3Z32Xfc1ti821HHRQ9Gb78PZ4
VCmeNjwHXVX1/vL9ZsilExiVmK6suN0pfvLyUb1h+qLOXjLQFu2P3o9EBNKFMhpI
YKhI6uv5LFLQBp0wCVj5YybemYhZojGS7RknLk5hN9ZfI4TflDjNUlXY2Gf4sE3o
khuUyQhYBAYVmAENVwE+A3S8+wtwX56CLeG/32vNvLvmy+MIPl/7JlClyhD9jj7Y
B0UWwYtCEAdo4EdgSIci5MtbEKUyFaXABjz6qPl7t98FTCMOM2ybP4nqM8105plk
WrGh19YE5wxUzs3MlKwKIDowHM64xQ05StGSc/zniWe3+Fb/wTau3N6PsWOjGGYJ
VV9YDPNNk4Ol53m8prVTE3/bgxaIPfsk8WZjc0pUr9Z5q+He+9ahYd6Q7LZivpKT
Ww/MB6CDXnDro9lqhv95qVYZl/BUwlr4fXleWDNByoSEGSBSChgYuIhb6O2H7vih
Gx+GvVOzWQG2IHTf0dXsTcI251GVlNeg+YpOYqPioC/iQDRO7jP9/wxkONawFsqY
62twaE+owyoDZGMV+Di5ii3AlIWEtNxm28G8x2XOTYVSAlY1xw5eKFGuZYei231r
lHpZ+MV0t/CLbmHy/hw3RXat//ZUxZX5wgb9sOzrykHB354DB73zsN1nfLMLxf3Z
7vDeNC+04MAbc2FJCRcY46YtWUw47W24L0cK7bdsm9KjsllX1vss94ozq8sRb80L
Gl2IzxYK7IW5sY95YeTmDk8OpfKEy1J8CjvZTgxYpvwV14cKNZS5ZtV91iVrWU8g
iLOR0llCmiS0PuZwbMJeXDhmAlcgoozIYV4/HoDNbs6dhTYu1cLGfXt2VUeKFoq3
71zDkFX0cb5pKXTaErbGgzj+s1Y7R9iD+827Oy3n2OVYyacHQdsEkNr55TpKwaMQ
m86t33nTKvV8Pb6iNqfFoyAQMK0060Xwbsx1DnUu8DIs6IUmd/BTpOv6A2ZgAzX0
zaWtEOM8vszjuSB2VXVhx8k/mSK41knKD6sNzqLVxnk4gmJQtPHpgjZzkUbpFw3r
cSZbL9uS1ddso4hwzOxBJ273sr6bmYNMhZF9KtNPVQoi/3PK7MzVgwaLRblfEj2A
CQPo7KfeleJXOJgQrwiIPbHZ7T6EaWkgAusGE+37R8/ZFN0m04/fUQSLqsAeedvq
mEfcmHiaN6NqYdiycFBaoHmCJu1HMMBCBxjk+iLji/jZHgJx7KLDlZrelpQjm79W
3KIGAd4wdlVOMY50pZ0l2sOM8uEMWBF0rDeQttS9H416UbrDcFDL8zQKoJG9Va3i
gsNxkv2JkY82HSHu50yJ0t1qh+CaI1CXJlgTXnhQXQeysoS4hTxCvEA76mOG9ghq
Gz5V9grynSys3GXbJ+L6/KDijZesCpbxFzAzPYNZWjQZ2bZb5IhrdkAeGvDK7G88
6fk8InFqEyaBOZmvo/yTKSu4Fe2E81qksoAE5o7Gv5MKWfkOH/ITFQrzJ/GyGB6h
0iZCR6wup83xtk/v90vsXmLQdw9UkXAKeHQPM0Hu5ENM4Dm40pb7Acrs9/KQ6Mn8
0Q1iXIzM/JiOlKgUqmTtw/VqjDTSR2geSqTo/xweratei1cYic6efvMRyUPUv36X
s3LegihZGdRH5K/Q/2iHIXFt6iuIQ8rgNA6OA5gY7geni3l4op1coZkTm1BTqoWy
ZepVQJ3qC40bCQCUXwFi1HqHi5arWSz/eVVOg7dA9al96xO4iGYtPhuCw5NFdg1A
cHslMxR8lOs4n198zMJiI4AUiJbPv1/oswFj/XN62ojDg3mBJiJbxCuRQ8pubo63
6ww1XdX7Av6mznLVDxG8+OYAK6QttpA826vI59l2vQ/cTL6Ji2V/bC9hHI+qEpxw
Gpbwrcw1jcmJM3aY6WPd6pPp9ne+Js58p19P6a3Hz/Pm73Gt7FBUcW2BZ1hI4xSz
CV8MXuxDhS2mle6wpMQTijHV7Two76ctfybDaKW8j/Std/Qv0c+lc+Qi0Q13E7we
zKMRTrR1hcuReWXvmt6FDmrx3mmt5IKkjwlEgqL1lu9Smc6kmmPRQBOz22lyXWvn
epDKup/vsd3WxbsdsKfHebWkwonK2bkAXXxnYB2fU07lqe+nZjFlqXDpVe4LsPlP
0OZ5lU/X7F6blmUUi5mrUOYkE4stom0J+iXhr6bMXBWSH4RaRe241Y14kkm7A7JP
Mx8XwWZhnOL/u0lSamgFsyscdenwBdCzPeS6wyClGzZQsALTc8VPl1PbZQhIbdCY
mIioC7TUOHzp7G03+i+g4/Kg470DywJmt0iBxySnaAinK6HANT7m7jxN4Tb2lCq9
D+t8go9RbusZh+mydLpGClkNdMR0UxPyb+Xt1kWhBx/zJBNU046YnEV7D4SGpzI8
zPbfLFyJNKjAq4jKh6SY/JL/Q1len0QGDzvL08CXCf1eAyKMbCMFOc+potaRYFAr
gJbZdOI5C29Sb3d3DfOUwGz/adzdUibyObcSXg3OOrNMONXXkKbVJTqrFLLYBu9u
1MifpwEb6v7EFcQglPeoQQZD5pZU2u7u/kH6yPJsFlNS6Y8F2g1wb9TtmRrqDCUK
ueX6h4obLiHPBwxc33KPYetUGf+GySEywUfrDO28JLqHrjhn64uFmDWyk4i+eytB
E1Arij542kyAksP2xE+Qm5E+L3NKa0IrQk/dgcfaGXfEP5jn3RvN7CLtrHJbsb9N
uUv3s8f97nDOzjwBRtyQlZbv3ANQAKR0dq3egyDaCZMFnxJm7iwKnOH9E72aAJNU
XtC5k0nJ145CFxkf3Lt2C347RqLQ+Nh8HqP+uQlUmECTIZ1Dwz5W2sCDgdMgXjPA
jyTJPoXZQER28RAnDa+P+6IulGT4hCZgJJbA+GbGwFU0zkSAeRLWWC/jEX1O+hcK
CqLfEVbeiDM4TDjTpPuiw81wXXm1jyVlsWx0NOF4Z9d7mjh04jb0qLaIKaQC6uAF
5v/9wlgz0a/bT8tUjIsB/TfaivmpDRyQGGfIvOqDT2de+M20CQJeZYX3UjolscqO
3FOyNgd8fYjyMHNEwixKERHnBW7J6J2o4ESFvh67BW9t3b4AKl2b56b8DgeoCFXE
JYKqlAdARk1Qs49C+tV1uTGHtbjqvn0EzlezoYxfUxXo57+9RG1YCb9NJImZ1MwI
QY40nIPZxmyHVtIMzVISWE3dwdDvj1sAnvgEsHLemjxmsxdWsKefIFHajLUnG/3U
EQ+3T7NyPuhkZiS/8Se2oH58ccD9XuAsOXd2L9Q31Rzu8Ja/AXt5Yl3DdkRxdQNr
bHUwIP5NLH5KIXayWFvZVtAu4U5s5zD6V0DJeVDS5uMiIzbD2ccYeSedMZ3mxEcx
RvyyVDTpmK/G9WqDILhhOzEzipnvYT5whYpJ8Dp3xN7DFeworAaCwwupqNwMH1ta
B3pB47wpR1V++AcNTnoLOZRwXuluh92l1B90cfu+JfN63zhaIz9cXQqKWBxyaqhy
wGG+beIEGDE+5XiJ9HECBk+IfMj8pHZilpPTNJGyNtaM37Zt/vMMZrMl7LaYeYAh
NDcOyoLNt6iZN9crj8eRR5Le4jlt1Mh4K/ki4ZqFD2iWKx8AWIds+CiINFanGL2p
iZS1vXBD+hq0glfhL3I9Ta6szDUSGJQ71MN15MO39VI2hqvR7L405BuHchK/X5XW
F4Qx1H8eYIJmGq7YIcjDjV5+hqnBWo4yifwcgj9aXxRTo4E9hpNcIjICa52aeU6o
X1KdW9j1a5HIbQ094T2ecPOSsVKGaezP1oLi0vrK/1QcyEBbih/nLvnzbWpvGaQh
q0+ir4MCtsd98ogw+o42FmG80qSVMdGJkeC51l8GdILXeFVXLNnewH0MKuC9P6YL
sgDiQO34ffcqxT7AWKZ0O/2P5Zw6oRLaTWjcbYRDHyN6JTOP2FPYJsDpDePSeLd4
1JDrb2bEj+DQI32K/9JpVG0gvIJVPSCfn2gVZTkuUezoKkeP3sKN9GInQ8Qz4DYQ
GqQiE9DYYMWGZzlMLfOvLc7ui9Uv0IfMDtPxLVgsOS54Asa8bnuJw+bXjBnQ+FJr
2ZiLKwFUfooIMKWtQywZeOO5/b+e9pTvn5BBEzROpZRCv0P4G1uLGUB4WnQex5Gj
8ZOqASCrsbuw+YlOH/iNHYRgy8HqBcJ+dVuY2UzurzcKCvbYiLTCkv2QtCamPTbp
U7edZa9Cz9coHrPUDxaL8U6g2aioePfumJUEFVEHucit3gnzEkG9dhsKnuMp6krr
iCAqaq3ZdynUQSiD8QI6VJ2HrGSFvRZ4+oXTkhr3wLI1dIExs5g4jPCCjwhlBdpz
AQIfXs4Hiv31jWJ6CsHTNG+Jc0W8oTb2IVZP3IG9qqpowxzDl9wWpRlsUzBqK/Vb
xypGo3kzKg8CWglhFtqx8q504t4ee/Kf3iVQOhFtDMTvA1iwJaLazwSi9s/pxNJh
wNACUKnj0cYnT3LdQe/6C8pAR7t0Is3V3qm1dp/cN7+Rgz6lTUALZj7JT1vJt8Oz
vcaZSig8tZFyuFezAeT0TtE1Y5curMl9s5zQbhrehCueyU/0ClymTy4A64jziwWu
cpBL3dUBwO2N0H7Tfu8bgfOFTbviDuC+AL/HJ7aUdwU8lR+/RDLRBJ/9hB16zjZ/
NNW6WlQoxl6kqW0IwtpXrjqPt78oSA3ZfDwFmjnwo5zMQJ8BCxxioKPTmiKmoB20
ZUh+H4K9YG5+qYZUWlhOpEh9NfWH9i/byanZtnhTRGKn7j+HDee7S74cxFCL7dw1
OuOvTG3P0TtckWDBp7M4NE6XzJj1W7Z/LRRvCc9hg1J9AFpT/BdfnQmhT/OYqB1t
SfrVaycrZNd7SG+g2MIEUgmKX6XJRU9xvJEzQjk0Macp0o5A8U79ysju58hQmjE6
5QXgE1wZeRoud2S8O7boXfCf558cQ/qHu8nuBRWYke/5S2Pds+WsYJwfdqCrbAgM
rsQjTPg7FJjllqYeOPRhaHPPE9NY2KFg4jELbgbvFkWgktjeGdl8laTveQX6myt9
s45246ZatglDratFkC6fccQx+1E70jghYw/dTwmLSwZckuD1JLghG7kLiC5GbKya
DLGWseapQv9QlvSJWYTQtEjsPqC50ZoqXpgCHOECRG7uuq4EJjckSb7A2JsfJEgU
kuhFfPiIbxGlBSJIG0ftlCl8mdCBsHgvBAVwDDCxy0DA+EPvS2Tt3LfEkd7qptah
hm28cM3KL+TcQBObmMUR5Z6ijLI9s+CEql1gvcWWDHLR5IdUsE1Idmyu1HaUA/J+
t7O29IFSykeUS3EemVAv6YW4JyU31/eDtevXOb5jew4zSeWYKugRbTTEYziLiGXi
sExdwxbbJq+u3Kuxe3wYPMWCmSNYezbbkt3W7eq2hIvInM3b8p5Qc9Pehb5GyL9v
xSImCWpS2RTK7YSobRqfFOqKUPjiF6ggJpxEV8lue/xB8gyEkjggi8p3Dbo3M/wv
WoumdZuDbt5ivcHiQBy1qWkNMC5nHJlqPum+yyAP9MFptCXnHIKt6Oxh8ocZIsj0
XNdbW6CNYza8cp62I26lAkCm/oMK06tricwEygPfRK8da+ueJaoZlNC+uKiUMqyS
MY4W5oKklVnroszoDCP44hLwJQyjvMBuL/SHHCYHjg8EbMHgySlkxP8qpGRNLXHW
+KFk3LiHdAQAO39v5R+JPNoSKU8fgjFWDHY2mVxR6H+c0aW+wMjuatSp9pObgFLJ
P46fwYb4ik6h6LLmq0ubHLd/KKM0YWP71dtwgsKCbOi+9eq+TNtGIPnANKbLzrYV
ADawyjRKSOmxf1yrtLZ90dCFcBdmTgPS0Pus/EPNkeqM+sVycbvOUdRR0ZwlCjKP
GsTM3g0CLgcSIVtqcfgQEE5IDjTlB9pHQ/aQVcAUMkDJ6vifzCycQzbf7NquOI5C
7OddFGQfUCipmyFlM4mMj1rfiPOFWt/ioHDq95SKikIPPuhH5mIgvBz+1aL3e4Jt
J3Jf2N3dTRpkhVw6ZiKqJf32cXT2UfZ+5UdyjcZ8kRU1Jn+sx4IT6iLv9qKXFQNj
+OBk/NKFYtxicLIidueEoT2IX9oM8Yg8PI6ggbWOr02IU0SGCEzBpaQKp5ePSqdM
q49gq8XkCx3vmNb815S4dR6b+5RI26rzNC+o7sbjibhuRm8jdRnn6+LmdSH9YsNV
GxG8kzExJ9/tQfI+p6Bcqz2PFq9e/iOxcSAd4fDrrXp41I16HupSdLgeAPOGsE/8
iNJh97twKYkLbyherxmypmwKqycb8lMFxzNgPCi69krKNkU87BBTWKhGXD+ATq/R
R0iKuOM4lz1RVtZ/R4Ixl7sNmG9L8bKj+2pjCZbKpA/6S3CDX0/jyUyJfzsNeAhc
xYgSDX/gpXJQpz0xkfQTqPrQsDuCVU6fFGIxOioFZO0ORH6FKlHu44lXE6Xbgafz
gI4Rj3krtV5AsGexLkD0daUxsnWp/v7JeLEZzsdMWr2s7cF+5Wv2//QG0AGkh56G
jBLGEZ8MGTfc645NKMhgP+sH2rK+dIs0O89iOUV12MbzAowJND5cYKTTjgOBXEiI
yOVX+i03Jf03OEX6Tk0BJv/suEX/1QcJaUY4JyksLvoStNcV0VIuUedQsu5/rVhy
OCK55maoBpRphHFDMNasd3i8TS/IDSkNuIeINXj0p/6lU1b5ZmxcxgbJ1GAD7sLO
6NW6JGie9OlfwjvKzR+ULdhSqGtdg5S8KYTI2565fita9vq+dK48YVz96LchAuk4
mXOnRIw5G0YWgyCo087cGXs6nxf7OiZGIqfN841jKoC326jESCqcpQzLuA1SBs1J
BwcyWj0U2EEMuLLn9+NSNVhNaFMI48ehKK9xMBhcuev77C/DyhpslPxcEpaU/7Ek
lql/aac1SfF5GVxSbVexFEJw7iB+ouoSw5r/q/VceYtyNqqzZuxzdZl5d11yRQQd
yVKHbC1vG8SKRMjbzbziYpb5fa6dtz/9c1Z95y1RHB3dbWkoXLtH9xurz7VFLBKN
5JpOt3aYxpOot1sem3kdMl8t16CW9PfCCap0oB5vSFyshEDbTeCZvCvYyXmar6eG
kklmGuNhg8ZHu2IfMG47yD+s3jWaDURyQJpMBhd+Md65TJMH3CXbuhKqD7wNnuOx
X84NFyOGNCaMl1b2Bt5RklLuXbAbJaAqkOiYNPIWvG1re/GNUrXLCUgL+5nazT+a
jfi+61lO4SVAyracZ/t3ClGoRbhw+7HwKa7esbrDEezUzxWnqNcIzk2xmNa0Rci8
jnizK0KUH/ABOCnR2zShVe3Gm9TXXKPUUfI5MuH5BJCxVvWsC1Pd6CNA6w4iJN6d
aG6c63X0uIY48LqJT7TWlFM9kIxW/Eq4fRaGyPlyO1NvWONYkLk38+KOPXJBdwzR
XA6kAAw6JLy8lD44l6rYN0Kgb0H8D0MqJ4hO+mvLNmTdNIUSChw0YTyYBKG7FkQJ
1SLUhlueCiHy0Vd7I+blPJ/++rcUhSxFxbNORREq0NAor90GvQ7qLJ0IS0GIFr0A
jEEStJh5oTqCcmvzb+BIt2/QKdty63I53db/+nDPZuq6ulauBm1k4pMAXQnphWFH
nu0IlD3vghxC+OURZYqUwiifsbQ+OOemUJmP6Z6uDLXnt1nwaI0Kp6hRu4AI9fvu
dGj+qYJ7k6qQmW9SQD6DeHcCMbCpSyMFUK79D2mPBr8Re21dhh47EqZ2/WLLdFSj
tJkaiz7Pwss6AHNxNqTzLgzk4Io7nXi+WXiKplR3AEiV5oxi+vi7pmUqCiFXX3sL
lIPq+yHmaxDRJsyc2rz7jFVMxeUhgCwu6u4yWDVYsxmpqAmdMgoYxejXuUkgoZvI
YDKCy+fxZhwL/gUBEXotRB/M1qzlZ+JjTA+4uzRcwn5fHWFq5dNKrSWLBxk1E3Mb
W++FE1BxV40kqLgH0icZXwWKpiHACFharZiyTOQvQpF6oScmKLuWBCPPnI6VKKrK
tdk4L/Rd8fk5BQ8M62Lm4xV0eN21Q66Twuu8gCmrrxmNUy+kGSEY528g1VK/RfUe
YXSq46zCLZlZqeODfPSWosP9Kaa7/fTxfhTj/NmVYBDcd1SkWdu6zW7MNWvp1uMi
jv+rWQS9vrxgEqdWcLhWJ8nZk6O22GICdhKQMIT628g5wgh7YXyTsx9tzGAsBuyY
i/sc/lR8IE4nL4SXqVpixpld+59oAUZ4TsgLBasxOZr1kR4jQKX0cSpnIo1UvR8V
nrSKFjwd6zgAoQNHt17ycyQX3TyLwuAN/o/MoizUUUwJraxSZaOLD8OqlE0iv2na
7taWWl7O8DywW4KoGqL6S8CyLxV568OyuCPPcwL6XiCJiBUDpbCHYj5T8f2DKgd5
/KkjJId7RvM/3dHZhvEg+SrchEnF4T4SzMh5mikChOsz8L9WLt3SHbcgC0qSQ7sm
P5kqfSjJ/mtK2dZy9Zgv5CNhWCwOU/eS7pXLoi6qIICA77Jge2DpM+Uo+If3pLlu
TV+8DS7KGCbI+68KWsCxn9562AXjHu5E2H02wZujR4LpcOIQJwyuAQfKP8n88ThU
ST/KJqNH1zlSBCHHS4AHZxyihfvSjvfJ0HFB5XivwKm37ESfcnGR09W5DFMbovGq
9EG4/nuKPY97MgfbjKBIyQIK3mEVZA+MwmHNVdfLPD/PF6fnTPOnGD0N5TIm1K8D
FMMMnicAc2cxQ+NwGvsXKN0IibMI9x2dz71cBMKXn2DTyjsp7zuVNP2fNUzzU0DX
xHQVapmJaKUzND0G/Js9hgrbUFjb8gGesrDRLYEYvTHHiUEk+4Lw5xoqCoAgU4xa
rATnDHhnOs1VzWfOpeS+RBIUO6ejk2pKp/BrfXxKjPUQcTH00BmfSeoJutp2V2rE
uwXp5Q/FgXC+HZYN26ofYNWeGg1I/gB0DxkrBe2569Kg58vzcH0cx9//+XuPJMnV
PnpIkZvH6OixKq89rf7qLX+5RC4kz91qMwH5Y/dpBJ0L5powhAf5X5qXbwni7JyQ
BHxvUuhzbS8CyVA8uPykKcIc+jfu7lU8QkP08VCWE1Qnf8Lq9KdhKLY9X36e/xQq
Cy7sfsix5xzKwKzryfWtPGAu2ghI0EwR5tVUAR9kPw1eA/oDdYTl1GFS4IRJ+6jF
PnZJgfjabz0ZmMoOFE1cY4MC81F/VV5LngNbZSt49cNjQ76YSVMUbaQQtcj6TYe8
MGa9SzeLNLQm79hmaYlMYLkTAZeRsEw3Nzg+J7Tg/6t/bHgkAmJJHtOR+eauLgzV
rRbrnYI/RRETyH/zEgrbr81b+rYFjf+Mjqxr9daZBWLtvzN4sfdLg4SJEsNvBZ94
l2h9pmj2x2tMuVmefK1xTASD8LPy1Qy4jSmiUIxXinMzvNz/Otu/In35kSsGINnb
U55C0zcanMq/gLuX9hldpeW/dOKqTfr4doHOu7AZUdtW257kbFVqyxODusE9NMgQ
QM3w+QrfeaQqGNY1kYdGVE1g2z7vwOrLU4eYy3L86+0DJRV7ZXJbHd0q9Y//eJW2
B7oDgsGHMuETG4t8ALXnNqPtGOCPto6NYVUUbtpPBmHXDkIUWRjl1U9sbRE1y29L
3g1+LqyYVYWCy1ERY/CguBLD712spjH1s4XKehGOenFOlm3wIMqDqdrsSqolJlgc
P72pfIJFNvAytqCvQkTwFdwAnqw7tPeMZ3xZqLiuZuqCVkripqjZ2sevTuqiUjJ8
54AXRZIZcSeOpTkq4na6lcJoODcfzzuxrIC6mSSa+Bxodav75wum59Yq0B+rNBu2
yIh7gWtxZ9UlR2bskRPr2f0fyG07PjK/OpuJcdKCA3B7OrCMxf7YXhNKuOFiTAvA
+xyK1v4o34t5ZM3sxPglxacNk9VoUw7F6rFDsvQx5D1rymwVeRE8XJGgGEmPakln
mBUoTsj6nLY2l3b2GRtB6Dw5iEX8U67L48q919NCN/wfYdscsM7wbbevYn/7A3Bn
PMFWHVn2WLO3kaAG/jDj4BxoIDwwEMS2WReMlZaLEQA0OViSk6BUl+yVoI+uXVa8
oyXsWwDgA/+3Uo/dm/2xkyCQO1+oPbSsqxRUfyLJGXRrNEhr5kVInHAecZ+j1rzY
wYd1XwcLqRG5onwlZ0VVU19XR8Nu7+SynXLgssrxbUOeNo3WX2aScOMxl14SXRJ8
9gps8OqG8Qr5vTv5hq16NQBdGPxALQwJ5vkb0YMmhZiwW1rD7vLWUB/eO+ENu73Z
Mcbkwue4Lm0HbjHN6Fc2Us3EqmoFloU8WN36W+tgDhkiPFo0h5Rvfkh+CH2mzURa
eYJKB9yMKs4HSf4t67Q+9dEBhQXORk70UFtb+SnzXGHR9RtptHJS8NBlQ+qiLAac
Wj67bKL3oA9gQ2JhRHTGnsiN09EJ5yTQHMspEVCQfryseMtGJgfkPQGfwS5B0hPr
Yk3yhQ6ilSi++g/biTrQVHZw3USYHCddA0eZQ/v+V4GOyAlGyObx9yYnthP5nAbb
F2MKJDxZhqBQCmP+TQSHdW6aaWSAwyoN4mSzMECzXjgIVz0KzqW4gnYihv34fF3K
nfg78SE+ZwvoBFqUp2zT85KtFMTe4YCbmYZjQDfquNbR2xjxJ/tk0jO+p5jrQyRu
755q1GERBUoEBxjw1/HOe4Itc2pLSkFuPcnSDB5gEWVWZyt+GabjsrGCt13GFWRd
sQ8gxVw7yL8YFeo9YcTrKgwbjsgTfmNojCckqYYgZOSKAHd+rZt0bBvzZulJfeOr
uriGN812XdoSMGywD5J9if+cWJYKlcwf/iT0o7tW6a4j4/vQwiuoMn9fI/YHG9zC
yLO6U8STxK3BwLglzk5ethdevYddpwFlYm1kfK3ZCm2vBPwdIfSOIHC3pN5YLFiw
arIkDFRQdLaO1wedrLuw+Gg65XD+WNrwHD3HDwlajB8VNHPm878dXg+Hh+lNHXhg
ON8p3CYWajKVmNOpFUaU4sXXxXmLOlQaYmHOMWpn8htpm1fyGT9wnAVQOAfR3lYg
jiJwqu9dUb761MuIGtn50t6aTLgZNwFsU3PE6aeWOzEVVExaz45L+ZKmobc0vfeQ
bp+qA2+1EVI/oFaUK8vmWpPCyc+NNhrJnaBQkuskJJRHvjuhlGwOG4yIieGQvTql
eK+bhn866l6TKl1zj+hGzmcoX38ao64+StxP7uoL6BQYEnH2X6W5zilue0MadeNg
j4iyZQeJeZcZ5gZ9jtBPE1Q62iGlgiDQvC2o5IcvlQlxDcTRmp7op2tFCmhKdYMA
/998w7AambLrE3OZuTk+EvDq3hkdkcSvXb3pY+4w5U4fUrdDC/Dnth/w+6dvztUK
PA+zyvkIArqSM1mnorPd93iD78YhizVnM8DdQ7FpdQVOKsjXqFnEpvnYova96Rf/
rnMBSnxm+axzctqkS0VRg+RGV9Mcs2ZpLbtHtXssDvh8Pn1aKfWnvVzIl3YkmDjY
qeJ/wsam3vLyJw60hRUVUYAK5QqRdLnlGIUQ/dKQibLEB/yw1EeaIpJ4c6+mGDPX
7OyjF4+90ZNeXlzEhr9IfNFemqCiKf2r07O3Za9CP/2f5PcNK2AQ6Lm0XqgsVksm
PC80ZrZyPCuYkJRq+1QzX4E2KzDtz08hN/FEEFCrjxlkm2YSlz/H+QwRAfpIO2Ru
WVGYwcLacMJBK5VYl+HjiURYrkxdbOnevj7MvCsPgroqPzQHJHlMi8MKtQ/hekk/
XKrMSTJdrphexILfQMokC7hN9EuuYq5x4QS9rsEn8Vwbs6oj0Gj/FXcCvwxm062v
FeML4pfVBkUw5pRUaeaXpJskq5WPl7RGsu7Y/h7EPch+aAwfJxvGm80K80wRfQ6C
+lq9df+hGBLMnsRGUGzbk0dtyT9yWy9AC+UgsmA224Lb98tNDUnyLHbk0bh71KBc
7uJ4F0t2ylN6WcZ+lUM5AjrQ0fugvf7HzEYxmkSun7R0cHeHevP3Z3rPKZbeoMW2
hfyq3MdisvRxy2UcDwaH86MEt2MZzN0HcuoWVU8zgEyNirQBcknhFEQfpIisrXz6
mTJwy3+ox37sZJzB0DtpJkZ6xZvSYQCJsatlLV7+aowRIW8i/VmZ5XKSTHVdGWGS
RmX5Onj50oIeIiwClOxYdOC3ZhUi9Y5lcMdhwfKfiQ+wG/tLDBcB2yaQhi0L7lW2
HsIzaquyXlXXCQmdEQZEU5Aet/fpTcSNwljUtIbbCsA9vdbcBX9OBDStxSY8ZT1l
x/+LeN8+6Q/D/FdzxNDxzOVm4Ruc9HUJk31Q7hpS4E1msBOf/IIyUH1TsQ02cP3C
nvt+1bdBKT7CEGGtHfnr0FZwv6kPcAeF+2ydP6V2x2lORIyiFsUaosqYRZ4Plcq9
15pSMl1zdWK5ggpC3jIy6ZOKxyEYZOq9Zr+jaaqfTFgpop8JejrHJTan2o7Lv41f
yxEkvm7d8/JT3DkShfO0FLbthpp/vkb1AGX1VGH7YJUe9gVXnAVCNF3Q2x5vQ3tf
dgIghX25503KkRRWDbdn3Qbye9pcC2+09D7z3YM5gTBnW/J95JEKseVU3M2pCAmP
O5+3Tw5hMSWW7M21qT35pbsbwhsYrfKy5bN6CW5X3hiL8mSdfTOck8EeRxCc0W9h
6qZEPeqt0OyVZNjsd32onbpUx60wNA2GPzF0lx70Px5fLXAjsDTkxnv4PkMac19d
YzjycsnPSq7Ig1RiRjDtV9yC4MmQ/+mERMIRyRX8f2Wc0eQqvpWDOtrq0ZCpVpw8
sPhGX8E8bTFlpsEu2iT6qCePcV/Ljv+IBFWCsV77LqqwAnGNFfelfT2eXIaZbWmM
W24sF7Mji/BePdCahJOaZKMXUWiEdLdgSTekbNGbQnhnYsMZBBn9h7pCFfBPt3hZ
GRq3dfQauFJjUocghC3L90qI2TTirlYClle93C9CEoUBRadKn0Gf+TU/NmLYHpWj
5M5BCjSDccPmLqimi4y+Ep16fUkT469qmSgwqlXCmISlxtawUwzi3UokBSHQRHof
dvMFHNEenrQldM+5vf7bG+1G1urpr6Yj88TzjYD/fwbSQvItN9c3nYoBEjXttqCS
WUPpmDGdOdOrw1OKO6Yls8D/NYRNBGl7YxJlXZAsu7m2YEMDV1ferJXSeD2IcPf3
8W/nENlNFS7cIMFjudLNgPjnLVBdW/2ZcLxTssZ23Y3BHFMlePbxXNloNUTZa48T
S8d5m5uEEHPHvmiO+ZruCKxYZDDB35gC712XAy/O8xhWA431eBi5nW9kJ375x7ew
FTF2db8/MqYaNcCYaimnLI7PzWDxZPtfWG7VehIWRlPKx79r0R1nXduFqupDMnrl
egk0e9rJu53AmICT9KCq8MmgzXf5xKs/JKHVDkNmb5ICiFC4hMTB/tw9CyzAJVZF
8+KXCdzuRM96Qr02ipEo637OPtbV5moB6Rdj/AHZ+kqlHuxZz6rWEQew/RVZyeqw
4A1VnMwvf3x69I+oKxx2n0j1H7DK5HYrjFzMEuVtVvqZusaMOvjI9DSBhPWUzwbe
DpdIEDXt0vw5xd6xN6Ddh5KTwMgd2HI8uT+ErwsQRCQcVeukDhm7ndt/jIp20A+9
LgeaDe06jmn8202BmVJxPpPwZPDAKHGFpWQU9XVW2N3u3kvjO9pPyfRHlmv+UnWK
xQn1LwTzU0qs/xxqxlhkdWpvj90rVHnoQN8y+5hFWCmrp/eEz4ty8Kkd+gEPDA4W
N+PAOIhS2gRWmTxG/+WCj46OYlyKVHJYlHjC4V/iXQgYoIl98ThtLhCxrsP3K/F/
Z8fi+iuN349RaYIg0RgXqtZlfr0KpiOrYg+JG2MmXcAy8cOwnH7RsvBjTp1CQvdE
YmhcqbJvrnHN3oDLObtzf8ydXc6S5a3ki3ZFubHvE/PXXE84pZPhQjoVSiT1o2Z/
41tXmW26IdGV6IZiL6clYQwNXBvm23v19ds6j5fsw5VBQuAYbgxKCtCD8nE8OATV
xbBGVHpXh41hUDHaswACoIrxSb+ufPAYyxRB8b7aqtoRgV2P3GPFfQGSqMGoNzAm
Ih9B2e+NS1mvXefIxprTDGniEbGBklfSV1ySoXehx2/8nifm4llIpNxxuQ94ITiu
x4t6jaNnhz9gnEOgT+ldVue87TXHY49MjmSpqCEEdKA2L35c0Z8yhiQ1zdvoFha+
IIjadtq9eMErJ/FLghFpaduTvlZsDNKFfe2ssEyk/ZbCzdYXGub1kb0St+l2SR6e
DwwPfCa0aRfiJYoo6L8iKhMqVWOXwuKg7wDAqErRQSHoPDinugxgZultGVd/HBz5
m1zejrFurIqrl2voPFDiFpYwvpyMRB8g8pj5C0HWTbDWPkwe0jDC1P/ZVvWYfiut
q3wsQUjNylqdwPbPVvvGg2TtT4ShsFRMa51mn+KcjcKguqx5GGSeG0c7iQbGgGPm
ObPW/84xjTCG5Cbi1u6PEqBk+VFNyLYmPZDwUS7kdtTTPiQMK7moTpNxY8MDi1sb
pGwVylddv0zqOlis2prgkiA8lddsHVxzJno6UDeFaq59BQoniFu2qVr4FX6fxc6O
vWX9KGESzqxlMPgAhgYnMew/cNyl7Lma327PWjOg9NZ+eUJLQvFkZcNdrxVOhmok
a6pLlSACg4Nbgfi8kqXM0O8dyKrAB/gavKViGxKdEjJ+hEaen0ZCFGxaywuBEv+a
orRqMU6Oo+8Z1zfe1QpC6gw5rs6zB2IDTDKYECRanI/WIthSbLlMkRc7BCxM4/Sv
xqZolcF4nBE/jYCa9SF4RgYRRVo8K7Nxg/GtKdW5e/oTrpwb++OUah8BNqypk2ZF
XkfUUYwP1UvhDOPWou8u0WBcT++7fsVFP7KML5qlzdir14ThGLH/OQlBYaQIRUim
WpZj5SGbCYe1MIMHGdtH7XlnfdUd7dX8yEISD++aSy2zWpTCjcHkHo7P4nQm0xCT
miTYRJ1mVHPzliicQAtF3s9H/70mAybgeSaYcPWIJSV+EzHnEF9yovAtR26CjxGu
KFhqub491SlQzu0ume9X3yTk7J59FE1fXmNRhC7HahoMtl+P6wkuN/0kwopknDrB
KeFfs1lvscvIhKs1JdUTi3fabcFWyQu6he/Ns5ItDJKzfPeQwhPjv3AMsUOScfOy
kc5JY6LjMF4nZrB5TQqaWAOM16GThKXp+NH4lrPHJaP+yzwOx13Ts9LfwHHyMie9
AviYVRn0AgcxFuQr1dOFVJds+V3LNa59S4xlyWmloiLp7VHSUHwaf5uSqYlroaTk
SLDs1XcSNARhiuHFgTkRZsf8fJZi28j6b9wRsNoHrMgzfjUT/1pCSAP2RTD3jISU
grhCE6ZnYYLYmr848BM0ktTlZs7xUvWVD4DVCBFb+skrzzURg3kFUaAoz6y2vbDb
kpSxmdEI68hvbqclzaHnE7g6RXp7HI1eF9XI+TNy7CerVzVnlldRl1df1A0sf1Bo
bFXloyVtzOudcNBmUHoqVRI5medK2ELZMkIYBDpAj+iKO5zrlWxSwzcYPdgNdN9u
b4oWleViHIzQxK94vEstGRXHb6ghoFjn7vV8LD3UN8u0AmRdBDw/6Q58T7RsLFJi
b5XCEHEr8HVheX1JJBjen4XpTlU0KQVeRIdoinGsL1Ryo2SdhoD7YN44zF9wkpbI
v2fNpJCc3/37vSMpKjO1fsMwaXUX5BYhVsgCPO8a79kZkKt0uBgah9edqXHCe/H2
In+WtFkJuCI4xvol7g0SQYVVh16ELPltYiPNVmj9b0bnWh2zxfSYAgvZd8FeYaZ7
Ijtu8QS6pRuCJ07PHKIfMmaAQT2VaSNxdNusPQT3lxy8PSRG7Xh4bjTozVvWj5Qn
Nw8TIeXnjwwFGRVlv3aGdxScTN9sk7oy7xebBlRpKRS3nGcQcEi62ix+Q+gEK+la
AUYbYpuZseZy+RJBRNsSqp9b5sqj2NfxRBVEiVUX3b0csRNI/MOJIzch4+gNlEux
hxDiMv6qdOBLlw8g4bhr5At1gm11rqExzuzJqljvKz8y6wEwWZQkall73GI7JrqP
0zEovS0lIWbfU5UULVaxEX1LYX0OxP5KfZwqItZ3Ho2QFfX26+J/3rEBZYke5kd3
jS0rKLJMOOT7ve3mGJjJqqBuqWW3kKOyBwlFd4u+9jcz6tMV9frmzCFF06iQb8ka
l8comCrrnhbIDZtCmtZUS4jI27RrucCzqZI3rDBogvpvJWxjgK7qcjj2e8zMvxVH
aVFM70PSjVfNlIhH8fiL+Ragm1lwNMu3l5UqmhDY4pKlgw2BoKRfva01oefDiDCR
JIXJnRW3EGBqTpcPbA5nwBZ1UV4r4kflMMfI+iPhv/eulnnpI0/GGSYJxXdWwsLe
SR7/3qbuQBG7qxg+t4GYwVGims1DVGmTIUw52AC45kohUlemmEzgSiyv3d6ICI6a
yLRsNcHwh1tQfyuJS5bVc7IzF70MMSHi1J+ohO4JzA5p399pR6+B5Ju3dkdMgyWs
TEj+nZxx663NUjCiTGsDQwwm1VohHb9vjUx+qbqqfdB4je/sTSNFX9CizfTC9r4/
6RuHHrtQfeF/L+2ShY4gcP7dhSErQOL6NkTMvl1bDmfVvsd/qwxcX5rWKeUndJ6h
1aNfsiDafhlCaQeYPS/O4Lsq1kw71twZn5RLNr0n07AIyE83PwEOGOhReg5KTVwd
w14AkMnt+UXrzKtDyNLjV7C1z0kPZiVXWu5LkgeeitWuSRq0koMEfqhA5vBj9eat
4FVnobWryIN9gi9y+30VUk9GrPXOOJanygIDijyKOjs/Meq1WrI/7PoiZYRxbXqm
KRFaE9vuNbEikQLmH3NeI3UjFTQRYfkfw0eX7xcvKfVYIUfyZZ2pSIcRbsOm7Mqx
rXmL1zewfD/StFif8HEEsWRJwcYWLafg9IbjBsmZk8dx5Ni2xoiTJ1Yq7ndysa2f
Fi/rXk5UqabuYhSDrEZw/VumomUIlCnTRJyWbEhloszVdfUPBA6eEON6sAnvbsmL
oBgNaBYuR4UOCMLF6WCB51Z18THIEvJnJ0MG9M/A8d4LFku5rlVseAWEbSVPT5a3
HEKgihlJAalzjQ808wpsxnlGXJKF4p6bAn1MIYvF0D/FvX270T8u6sBCJD1QQ8iF
5THz+0k4R5VE33D0OUT5VBgzp5dokfKwLOKGFmv3IC0RvW79chjE6OvJUbTS/d98
sbLc/5dNvs21cPdsnw1VSVBSk5oPnqv3E13fgrl0aeIGboJuU7oeqOL+enG2V161
dvvoKpzFTcYT0AdhoH93L4WTMA3/MbYSLvt7/F/eMYws7rXK388fOdHOsS33jsJT
8I/Ft53icHxg+GbeJEJyGi4ULwKZWdmPdEjrLKbnQbNa3hXcOZ1xOjunbPbazTpv
+bV+vw4TYEUbUGLT8Frb6K5euZRXrQ168Dtr5rMcKvRiGdVRRvkWk/ScumYRZ5Cp
e/BaSV5j+CJmYEcb4pTfchcDViO+4Kj69AnvzWMO9vDsmU9VHUo5J3pKAxNC/oiC
HUe6nKG4kioQygQBm97oEKmgsZ2X9NwkXEGP+gujU5CH8/YY4KsQffh1CPXOlN7K
tuRrhXJx4JFZ+WQRMQGrSkaU31VRHDT2/8QVArsZmD6cw4yHbEs4pzhdHNNboVHt
MRnxh8V62Eoy7veU9m3bFPuImQ6TOESa+4OX3nuNbrL2uZ6CvyK7QNZQ2RtTBM24
5TOPw0qJBvL/aXlWsY0VAsUZC6AiVnC3xdr8J0GgRTxYJQ7Sa8U46RmTsemEPHyk
kkEVEngrX3Sa3Zml6Lbj2GhEyYibsbbjX1LnMhUWLJc9h5q+RVswh9N+F3emfQTh
Ga653BotAWrivXztLJyCfqt/kNqxgpHNk4lZSRehpwr+XeQ9hKQSVDo/bSy6LBC3
fj+F4BNgadzifZl+DhqOlK6c/IxT/KyhsJpRFQTGlX6yN2FHvwMVI7JpJMHd99Et
+/PONIbSICvi69/6556y3E8u1AKhD7uazJ+r4bWqLwnVdUyygx6xZAKIswvNDfYG
1LpziP/7VaN833SPzBvlaBvdikw7zpOl8tDS0iL46RlUUqyU4YaLjDMrxirj98aw
VNr5PYT03+sCjrtoQD77XvgW0zKx2fzjwuAn/ks6cfQBoWCI4z+SmJ/CJBRoEQug
NPP8L82frH7GuTsnsNp/dsytkU1RLvMnI00ruNxyEigMuaBFzeDd8a0AK/p9g2b3
IpAvzJRGEkI1q2FhSHa+xp2DNJk/n8aXYCgAPk5Vw037Re3/xlbAv1LXWd2l47Ea
NwgmwR5XYOL/1QPv0zZt8CeNY2AsCIjI0A51aq5LZx2ZkGhio2c+C0gyJ9SGfHF/
hgz8SM/r5w5fz24zUmo1HIEttFxiVsChc7mvTs3VvvjbsVqoEafSzt43L66/HRrW
VrIY9zH9uNsJAwPsbva48TwE9eKh22Voz7ApqFw54pUhuR/qeY3u2RZLu1CGC8lB
LhUoA845SKqIyIYGXzAtLpDy3OiOzWwVHcGd/uYvQc88jaD7tvKwzQYVKuCLoMqt
1MzXsGD6PR6tNGUi2vDuMTfHRey+GhAS7D26BoJQbKzZR8SfoyF4Ae6jUAnemfls
up1ZTXBaRYbZni6/CZ3z23c+JJirzrKdgU/Rw5HL+E5ZtW1fg7yhM+IJf+wBCpAn
8aspTeggwFAqi3L48wWjP5dVG136kGEypbZ5kBYY5zQ63qJbDmDGgTJgMXkQws/K
Jce+80La4aFZPTyn6L7g5qDYzM7RzJ25+POxjIcjT5QxsMuckZr1kLuwpklXGK1x
pESLOUgFKuNwD96vM2Th13GvC2mlxvnwygzqx9l2bcupoyPY9T9VJ2mRs4mg77hS
ucSterNDw/wJS02vc/DMeaLg+VSTAYodI47EPgdG2U58lizfYTqNopOUfxNofbP9
wdt3BZGTnissMD5wUHNL479y0gS9dfwJh2iG69bM8Ff+ViUwaXxEuK9ixqkTwfO4
6fX2ZtoRm7W94SSTe5hicJApiPnR8GSTuJ7l6XWCokqNdk7NvRvhQa0wilGPzpq/
rE9/CJpZixLrpsTUgshNKPcpIcqGw/aqhAGqJNHnECWE/i+RCM7XrYmL+nZZxbyA
ZxCxT/Xj/8HbooDRlIcdOacBOXJfroIwmno7WcOQDFdBwH0/c1AJ+yK1h4c2j6CL
esxV0Jv9mZzO3vhyLG/5U7gnB6prbnBOSp2JkxWjlbNRkPuaA7vg1Lt+fAnBdVr0
Hf0p9QKlYvMIAiNwgOSE37jp63eD9gHxWD7Mk8EciEWoq031/JD3nyKX9EpWUlft
Q56AdUh/y1WgrPAD24qmbGxx1TOe3ZrtkV0t2d4kFRYPYh9vm2k3VMdAgmLRp8TJ
t9cS2x9CJeI4y/K6Hsf5Rs0Fc2tGpn02C9MG/n2VImwwAE3GAMp11dN/aMFUiKal
XznIpQy6D0v2V4xtveYSbiqKvcpVZTgL2SzzOcfl0Ub7bbM3wCbbtbuIpK+Xzz+6
gntsQSBZkoTJ1wDFTzKtoGkSIjg6x/fmgSaZaSCPUCQsW7fB6s4LeBMoOKaj3TEF
uHmP3vgYaGTW5ityC4A/yFNveuf6DqaIAvH9zoypQj1qk246X0DWHsy67iu+nf8Q
fBe4HKHqmhHc5Q+WvjtWDvFfQkopc/4QWwilmxGDVlvX4bdMFyVlxm+lsTFpRkz6
TEmz9hMt69QdsT7IYFkFaAgLliQdfvrpi4ZqwXO5AZWN4GBeuwEhc3G1qL1v8Brd
f2Jik8QrrM1w1FV8Eady+2rj4qZPEvrUXlIbVyLByHk6FJdPV725mO3Tle8ZH/dV
f+05SluiLikqyj3If59DUfBF/da12nF4J1SJWUvITz1h5GrKN3d7/NEZGc1ia9QO
RdMQBxt6SN6Pj1DiZa5Cq9U9fcWBlCIFT8dzHOM3D9LvlRo+0Sl/7HvdamXWz1cm
qJRuShtyW//F2MxvIzCnpsAUMIMDT+gPty5/WY22U03nAe0eB6KcPZCWWSNIJ6Rk
IdhnTWUorWxu9Avqgmn4OXDVCtIeVGMbYzgnOwIYfx0XS93pbPIWeory9TmldT6U
/No8qiMlOkEe+xfHFVGINIMh4AAb7pBkO1uKorqjQrfPmc9QnYzpzk1nnRFCxXhl
BG1Nt35/Ymflo8/pnGSIr2+iGVx1RLZKTzTfuns/We+xB/FP118C67BEpbPV13ff
gXadpDB5Gj9WLzJq9KMQvJtaO+s0QisEYJ+mHPccYNOuDJtz8r/HGarjOR2YjzyH
FSpZBATOucsl1d6ZYeLtlN775dMUf8H30JnyEPOFeEdTcVB1nGmfn5l3zBMhVcRX
+4afkMURtXlQXpICOBBZpsyid7SwhFBDgkA/KTS1fllQ9JY1l/6qZ+aGwximN/qJ
H7yF5wzpje7R7nNFtpuiyF6K3oTSjf1PX30pUXljo+3lSNT0Cf9qJDygplqwTcL2
Gnxm6tttmFA15KRZ+RfjhkXd2T3qTDRo61r5lnmXz3WvpVGuaYLLfcTCvlE7fUn6
tdwSuYVPLZiRoTbGQyOlteeK6NE+aFHOZVq44m/CL4DBh2CFHoS7lfC4xYomWasD
krEkuMyLOv602sUALRzjqlFGWAz8z+NpDYybsXym96bDpGsxX8NOI9jvfzgQ1bop
+mmOCwQInGv+ce3F+AcaqKGFRdYodWn1NyTGLKAR9dkM/fmO6WS8Kx6P/PxAdCz1
nMznXpUue9PwgsOVXBLXaxv0+zvrVxQ7sivP7WM5YhEzCXiUsp0xQoK/5F6Gh1kU
f8VrLREtUMfvqwFKgXw5asS/7seMOdftUWZyzBfgdxRKOpY1Fvqzp5pDXYM8d3nW
NtKhP8LX95Sq9m1o8CY03LygzERvF0EzK9ptMq5KBqStv9C6TlDm33oTNJylX677
vV0wMMUx10WdzVfw7bjg6zk5K6ARz0xNXoueeOm70c/xAzA8+lOwaTw+ZxJEFCUi
ZWCRwfuodS29OP7roQEctAKPxh2m2D9r9ebFVhRXkD80DV66hB/foU71Uv2YKfRH
OQbfnOJx2XkrdvPdPoPfE271ajYx2sV0i/0ZvQveMTxPWQM12UvvGGGwoerZJLBU
E7Iwyp5Z4xSMPckkhkpMVVyG8z0QC00er81QyxQY6F2OJZKYgAb8hwNJvwOM7QnL
7FUJZeCYx2J3hYe3ClFr++wcMs/Na0vjJUOiDduYYooPgsKV8RZJnIfRcWUlumaM
b0g7E95UlbK1zNpSbRSNwPNKnhPrNBAlsvT2tWYOS+K0+aSl4nUTkJDwcisE6nH9
Ta5rZ9o1UV9wh5yQVK7OJi4y7FfBxCN8wUWdw1hsJHC8dIcLuoOZwqNGZud6tX21
eRUOADLtIu5j6v0VNkmrdeppEZs3O7mWvuw4A5PFXf/USEvKStSgzmLhLCivPB8F
vuTbn1xsCM8yf19YGncx4hiJmbu7A5iJKlsPsz7mpsfL9FC++c5m214mrqYyjuBz
RJiC9SsEudraQ0UJC3CUnf5ogvrW6CHAjD9A+6Csz2xAMPBTybLLHU1FiX0wh241
X7Sl03BKu83cyWx/hj0GnA==
`protect END_PROTECTED
