`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PH6yy2IvUg9n73MDS/cwS616pFIkgU/ZoArqaQpq5VEXiRU7Y6unU6DCVWrNtvqE
3fx2P45H9n2S1/BZjIKXEgYjK1Ld9pilpjsG2KrTaKkKJJZfh42+f+RVHP+JIby9
iRyQRs7lC0CDCBliHrzWWFJdnxhepd9PJixmLMWssCbAu32lvGOoL660lbVrqXBg
Cjuph1oKLYBbRoaAifuKCQM3CLhikzRtMfSwceHotSpc6+9Bxr7Be2x39veDTyYj
xgjwsVoFSAwPtFL5XKLlZifGKXuOCZNBmljr/la3/FHbCsKBkgsRx5a1MfI9PSOR
xWBolSxyiJYwE7G32xJgq9lOUX6+H4UE/Sy4eNwU2phc/18KMgdkMPBM0plaT7Ko
xPKW9Fdhy8mbEWPx93B43UqQMiNfHPJNaDl4SS8o7M8B39KoAtDi91ngJwYnHNcl
sYiZ/FuNB/yjlD+rFzerolJduqjmUbL57GRvyTKHp+XEbe+idTt7SjhEF/I/fcHT
eEaE8Vl0zwFUELa1322gRnNU3NqA1VCoAtG99anuHZxXt+Z86FPrAYzI3weC4urJ
2l6jIG8XhSALJeWWTGVAr4kdONG/+Iz1gA7UuWL5RsCnqGwBAU2y3dBYW+VpW0x5
JBzXI6OQW2af/ZazpP7yYQ==
`protect END_PROTECTED
