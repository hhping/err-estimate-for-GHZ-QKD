`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPoneLUxqI80pQ0yFowdegZ4Fzr9vfkiclosqdXrUv5MXd+IiITm13FSY4ACDuLo
Oa7Ui/yxh0hAWvy6O8v0BrL15QLU98x8rvceyV4sUV1ur+CDrKLCfpq7h+iQDKp4
3B3vBJnjUlLqqjhLWr6IsMtPQoc3fbSOClR+/krf+vvYaYxuVH6tyAJZrAIv9qST
QJhyf7ZAGkr/m4FIsu0K860jZ/5X6x/TuyECMXfTHzZ3pew2nuN2ODkMb+DtEkoG
LDiYqhEHiW8Gs8BN8h4aoUE2kIzRsCSZXdjhksIiC/23b1Tp2aBjuvS1GHMHkh3h
tQoUjKnKkjtFeHU3X8n9PoL84JA7p8yj/waujp3ljaRMI7WUCfJmT7NzRRlTE3to
wgjQjtFXhUyZIcJwiRZqD+YewE3k4HU8UKXGRxSoGwvc9fDvjJBpYG1pD5lY9VsB
`protect END_PROTECTED
