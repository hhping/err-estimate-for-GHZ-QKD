`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5XjT+MVg209gocsUZVUMJJSR3Pf7gmENeFAzfJhy17j3mBPbLQWgrZBjn54T0KW
T+YghMNE9hJDcU1BpndD3FBe3WAwi3vTXPIwzeaBHJGXaRSA8uilTZ1Kjz0k+HKL
Yp5f5ik2Kkw1SCqB6JWePXVT+ZJUx/5ennHGWZeP3wFAFkljQkqmWUEwaHe+BNqQ
MBtSTfoJdVj3pqPl/hwIKMyKzgkSe4Q71pM3u0ceIPhmbnTselpyDJL4JAKU0Fqq
V5agi1wOvxGHdLRi/+TkMC0IN7xnhrDPZYwzpu1im/wHuqIoaugR2URmo9aCFGWE
wZ8/S2NrrkjTRYKppJ1A0OYpXONBwjFIM/Iy1OyKRHBqP3mIl3eYoIk0rUI0bPxk
8no55ixFREXZbI8C9t5IxQlAX2q1Xg3FFijYBwqrfOxwu63sJMKvIEipbmbSHz2X
kaYjYFf98EdOlkl/wu/c/Q3QBU+jwmEeaR/cqeB04dEWrLeZKf42UvVOre8tFBSq
aatmhXYlnwva/lmoqQ8kR1ylKa6vDwIP1VnFZZRmpcY+uPQ6iH5tYqGpo+pZGaSk
f3wCDauCnw0OVRmIzYYZtUJGgDi0f96KIbQTw13hxLZ1WXomXugJtJEEBJAez7dN
Z8z8WmmkMVAmKn1SSlhc1CbXxWzwHLxOwzLfNlLF97iBIGrbtZQlysco10OpSzyk
O1s0H2QjUrNQPjJBGinz7who1GeekhbOX2OKHFs3TzIILfFSizSTkHAT0g7D8s5l
sYGlZeo37Jj1HDxobbhDbnOlqhYhAw3BcZHDnTy49L06EqwpfR+WFWnC2zwAsLka
gvCKIvo1/sGaaMw7txU+aqqTHK1iKIWbFS1f3zGqYteF2/jNHr/S25gqIT0CA9+Q
TPHzTXhG4z0Ci+sgBeaYmf2ThR0t/vNoh9zjxgqOVO6WcCk0PZDOtdPz5xrE+uic
uvOSV25zYBdPhlMPaK88Jdho00m5HgYqRQZPZufQG5lkBG7e+rXJsjhf/Om+4tNo
rPE6E1d6+BtJ+CbAWTk6+5xLXstfGgK+RkrEP9CRujyWdu1EcaOKvR/TNIQDi1tJ
LHfo+oox4gsm88ld7cdbWVHSrwIKMClX3zDDR/GARxzihQeZPWygy2uc83ZY5FI4
AKS06jW9CPgY5V6/dHeOxKW1wnLIjnDnVoR0AsUnt165j6zD9IIvz6m+wIx+u+lD
QfOZVTWPWOUJ2DHglO3Z/LmRgvqrbkxwH3MM3qnCbXacxn9ZDhOGu95xL3CcPHwP
OJFwbEj8PYxKmLWQFVHMVyduJMIBq3ck3Yn1qgODgo6O3qnmI4SVkW+lMndoh9RL
vgZYWHctUfhgheZfcjysZsbXLOU9dK9ro3bVHpsDhZKwNewQ0P53FCtbOWpU76KQ
XNTrQmZST9l0auGKR4J6fOa3QahwVINrUJR4DlXbYRh7wtHH4FL075s5WnAaP0ZA
Uf4kd49yx2uBqeVBUNzBpKunwIcvTyNMBCnLaZES4Z/L/uJ8CqeFcHWqKtbB8Wkn
MV2UtB/ivPGRgF7BfgZ/8cGECKN+jvZan2+VEPxLfex2dNqG6SsAeYdRfa5Z5w/d
+K0zahUTEszdOchmUmvaLAGU07dFTlC4Rl1ZAbqYhqXe9aO/JKWL0IF96v8G14Mf
oCVcM1S3ht4O9n0Zi7VXD+I32XAiCQQgQEgwAK4pErP0pDy75DJG0nrfLQztNePA
WsknQZh21j1RDM6px7OtfEpEmeV9c9Z5mln5fsNPGoPPweiRCfhn4RSypBPMkgWV
05rhC4bVtrL9Moz6ClRChMUzOiwUZ5Z5Njk7FltJI+Pm6VqLx7EpcB+ORPLl+gia
ieYrSkGIRfY2iv93enotqJRVj2sWvEPAcAWJeL24yN9ueyXwVTSHorEW2J/6gPdp
XpXp5EdcenoIh/vLyhjomHT1LIXwYvXuPQ1PrNhxrWV3WZiFnadyweYztUcMvg12
LEOEkfPN/8aIY4SDqwS9iBxekCPM4C1xXnxi9o76pMIoqImrU2XKhqXUCqEp6Hcs
42GIm12wnbhY4IOGouxB1i8PvOseugTIeZ/TSRypc+fFru2QYbG/UrIVA5U0nx9m
/l5Jve8+bLnwR8tikhd8JN4okhvWCvUJvCjbN2V4ph1P+TazP5lzCWiB91L3IoOM
p7hUuFC3k9Q5QJ0Z5KINqv8Eb9fwda7g5hJHmMQm7yxZGratYs01y39PzwrVsGNZ
quZY6NsJREG9kMnDT7qlpnmmveooOuirPyykn2SiNzN1ujbbHKWodNZXtvXZMVyT
`protect END_PROTECTED
