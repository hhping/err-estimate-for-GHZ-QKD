`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbYmSYzgOvGXus8Uar3pZQ960tJukd9SojdCOdbRX0F6gG9uTOkjI1y6LUrlwMrg
D7VtwAh7Bg3ZG5ByVRGA+P7pyH5zyfbns6Cv4AK94LyeN0U2CXEPY+PEhmnqIwIt
85VT7B+2NDJ513qyQckyviJSYoxRWuc/lNp7fJk+0T2nfNRVYM4JnR2IR75KK8Mn
haCTA7Q+/U7Qc7UPbAzOVELfW+XN0bf2HniwzA4yMGoeLqul7vrzxpIY3yc+Mv4d
JLKtrMfdVDEpDUyKKA4YbSQpxmlLhIgJ4NcJFLmB0c6y/YKsaiSvxQ+dN5CFlm3U
7EjDJIcz0A+JtuZJw1OXpnYGxQqXbkiPH/qj77MN262Ysi2wWyJPY2mtBMpWkcAV
UvnyKbQKqvFgeeBUxXypp578ECtTxY/cQg1jj6GmAHWrSVto/Okbl4JfR1hLijF9
RndIk9G6X1uEhUAQK0cDKfFovk1Ug8rm2d2UZllOKvQi58jaBJIPalgROOKxvwj3
6Bj5ShWDeaZkLp0mOrCDd3eIcAeXdfLbpIgWhMw/40ETtRegE8/w8Q2JxPT4ziTx
VktSXTo6JYUdTvuSJ1IjJchwY70fHn7GHF5dSPwWiRyMKcIutxpVP0VSiQEK9RaL
15Gtvf/NXRF9pM1n0Z/SBxNeqiob7NZXdQJofvFekW/yI5PTVdqeBVpGulWwe/4Y
X+t473+7Rs8ehKdiuKA6AOdfbJ/zA99J34dHYqm3qm8FBfQ4W2OABX7Dno1rLD6e
mgh865FUujf/YGjEjCG9N7Lf9W68QVEdAXcq8P+le4sie7SQ9/jqUreQrjXBqbeB
kVIYVVJHWwrmh1yImlRHQUM6IyXzOptJ1ZA276wWnybPgW3ifoEmZbwpQGO+D8id
RHlVpo/+94lJD6a/RvpmUqWYymXemzUjgTzpDnpLUQEymfRgOXXwyDupIPzXke+G
wmiv0u746pqAqXT9M2mZI3uw2z4g2fwlhrivCQz9pz0g4WenQYQw/ltrzIiSDLs4
QfyRqjNe/Sixi9fiXdjsIrZ4FuSkegxvR2IlyxWnKrhXuZOO499gQ3lmRqS/vR/c
RwcKRjZZIzXO4xut920vlIDEFatkzhz+l9o+XAsN1B3QRQPTiGUL1BC2V6Jb/lvV
RETpW6osHRQwxlTrlswe5S0DUbt8CD79ixpT+eUbyp8IhOPqj3hl93uqD6a9sDX6
Ixwu+uzBuuxsHa+J/8LU3FVWPI2PA2A+AxYGv15fYDpJqOaIuGZZoZSCEmZR4aeD
Db0GlkXlFPaaVD8vdCSLGz7T0eetQiSdIH3NFPQC/C4Dxwt+zfIwSW6ksrJqir2x
DMjThBozq9lCCGS2hAH2FtwFcMhApxlhMoUXzpwbH4Q48/lY+fXkk5zUfxVp0/ui
xcYB5kPsRInHLokCg3RDat2Rxbb1Y5ST4+wK4t+nIsYy7bDnPfysg6DwNTZzSiZw
ucX5yq0k7d/Kl70f2XVSojDPAiUK5gLaZe8Q2++IDeMF/XeW8ip/3WYmptg3x9Pg
LLxEnxm3ZsNWbJKjgNHukSDaG0xtF1TO1fUJsZFIHdk5su0IyDp2l/I7BsYljSvY
8diE8wkV5WCD0oFzO/fXmAcuePvOJ08NoTz/FBxvPTFDqlGTyIweOVzmaQP0KvaE
73oPZCabqg4wia/mvTivjBzuMDoPEMHgy+E9wrIeo67OLzhFNZ7t7WKc5LeR1PBq
yVASDEfMczIlpTwgo4OnqqJa8cxjUIRbnoB41xY/Q1oR0j/uD3aDX04CAtpiqRgt
IM+WLONKLI+fxhSL8Nnb5Ty2vzDWmLa6we5L52LdEkb4Pt5LiOKlrQ0iqZYUvsju
QSJK43uNM5PWrAVX+LGyLSvIIPQJdQidGJsC/fPvYE/9Wa+chnhxbOfjkJGUrMzM
sgTRAaU6DHprPWNvxukwO66DndpnMEm56C3YuUoHZlAXZ2eWMFFjE0/hI5k9zSb2
6WRkmsHUkB95FRSmzEi86LDSojyTNs0G5hzMatfbVZHhhzOZvT/CnEkej/325BVN
ZW4lWB4fF6kSKBsdRMOH/0urcFUKdwYGfuHITPvfNktfvpr9F6rL1r2vMXVU7zVg
Vph7Zd86lAASTz6WdLRl4EAaa876VsVA1x7899baqBzTfUIyE6di1Sna/Ym1aNN2
ALV3Jp3d2N+hiOOHk/9gmSMYI8sIA/CfVkLLOOm7zIFXG+xgB3+/VPvlk0djS4cJ
h33IHXT5Gx5i21x13TSxs35Umgut/O027FzAJhaZGWEjCIwkR8F+4qeJkzV8g041
g7OlNP3rTOPXbCglLKYV47M3uA8A92Llf0KwdeHO+hbNCKTJo8nzE0yx827/lUPL
qSJJLasCR8FyenCRAYYdtI92KHbKKYUwDorcPqPxu2OQG9hknvYId0CD5BoQGdZD
/Ln00S4qE3oD7rE5EWarjWRxvlPK8n5HqS5oYYZMFPt3xNygcwl8j9m4iub2i4yL
8XoEeoB9MHPixid/rZFY2+OFOUPNA2UiilcvyqhdWn0YnL+KIhKi92AvRgRtRh+X
bl446DoxngWzi8sjTY0v1p5ywitN4NLHqNHBNEZ/6Hr6OlJ8UfzsKahyFs+CKE78
55KedQD5PKZp3ItjrY8H5J1eaSx/kVEZXy6JAQbGQR+7CQTck1BvjoHvcnfXddLE
KEdHZ49swPGWVPd816qFe+RkoUOSJsYDSP6NjrHSUhvRSfH4Hv7LTQCPHtc5s/ar
IF5Vrl/sR4VAoRv9Zc5x51gMG0VfWYWxSJ6K8tM5yGEwE5SBITfMWJVovXE+EF5R
5q9cdTJGCVAwL7ydJ/RtTDy6MwJq87ITzNLzV6De7WajBH+8IJ95NoTdC9ZCcgjy
aJaabr4ZjCuRPnmFYJR4JRrqQZlUOEEvLXYDGB43JN6JpDRPzdEn9tu/RWLnOQhs
Hm5og1PsW+JxYWOc3wC6XRV1/02xLQY47qr2KRiQUhjnwZjnQtZHZmBTFHMVFe8Y
5ulJIyAHEBwMrQH/veJCfLTPXqxzfTTJmuSiIe1PX8gzxSvVgwC2p/Fv+9TcEfPe
fCuzvSpEyR2yg9rpIIj7sJRT5PR1Uukp0OrdfuW7g+m5FbSG5p4Q4X3mJycZmIBT
29HvlZM494XceqsW8CynVQYsDno+VoPnwBcgiBaNXYVE65L0Ii28AXlF9bccK0i+
rlZ0FYmEPjA9VjzhazPHJSosKgMYpwmKlwKf4TPOaOf4ADEazPWFJosY9ghnOUbG
bxJO04Cbdxl5UE0HHTO1Vfv0zSiPgF8HNHq5pCuNejanVjppjaqHYeaWFvl6xult
NEx8xx0qTz891s/OZTRHdOHJcpRd5tTG9wN39LIRTsD7rPfw9hKlCplbDJgw3ZgE
4mJ+TudnyV5v6W6Kkkj85/aSjrNGQn8xDa2TeUC0pwWTqI/WEeYKOi0w5J0KnqYf
+oKd8TTnfXGNu429oCqGpgOShhU6rqlDs6t95D5bOo6Mp+T72qCW8CW4y57xy41c
rN46K/nbAqOB7CpvCS0PkKCLd1JL7o5f6pSn0V98c2muYGmYZfIoq3TfHHNny2sX
iAXmdAFjNqp0IOcbKe/gZDeZWDBOqeg6oOVbtcSvJ24mjwcYCpx9PuKLKdgterRK
hka0znmH/3EdiJzUbxGmAg11eolPXO4y1EcvtLXt2CAcGyIEKsPqobOcTQQKIqUH
lXPXREGFyLvEVb9TgQMBOSpOAYSe45HA83Ftjs9yxEJwJCR32j+OhrcxgbiSwDT0
jgUhE1NEs4EBZdjXHdAlC0Q368rwTXK/k0WDB/tpIRCEBA0xuI31HGS6UuC9Ar/i
lS7Y+/yhhIzKXh1DCDTGQDacx7MBiLm8806/mus8p/8JKtcb//h2EkjKsJmBlQD8
r2EJSvukugIPPMvuNsMOjYEohIYMdmSCPndsYW6s+xqJ6V37e7VnClP2ZIaI+fRt
HFlM/PrqNpkqFcU2tiibsOCNSBkq3VOSptJViWXrPODfigdO+hzhd/oOGnRqZIo+
kM/g1WXCN7HZAc073TjZeSOElbKrIhY+X8FPIPIYCQAwVLI/lYy/5wb3fCTQpveI
RrLfMzaqg5nt3cMoCwfmN+CvhOLgzJpa26pKajGOguBJPc0modn3BFtEbQdeCw0O
dEZTvNtHJbQ7LZ6KO8IU2GlpfH1eA5gZrmvULPlYKl5zQKrD1sGTyvOKDj3d+Hfh
6MSHt9g/TAWyPftu4dZLuXxi22B4SoNkvzC9myvcrqkczOr8hynIFs/H2zis12Me
OYRGa74KbUJ3qsi3+Xgh0PHUP/Q4eAM5eaKxidm7vhRO5djY/JZ5BrnwC/CtRrFn
UCfGbno8nrpbmm624J/a9KY8HcwqTLoA61fCMOzFO6MCgd3bDIk2Gn0qvfOR5OyY
1rGtCiigwxd1Ud12+1Nc5/wIrvBZiKHHUnyYFwGyow+38mSzbotcfw32qHXKHP7u
WxjLHZicJ5U6gc5oBCAeH+7X3ltgJwJQfbipWZNVMzYKjIv7zhFiyYTcTdPQaTsv
81WXJ0PaSN2Q0W3GXza8mavU1/J8oTfQgDfLv9IeNmFxx46wAx14JuYXDq+q8rAi
iXcqC9p1vP3jTeF4VPZ9wpGyIq0BFKCoPUtJr2bzBAfPYdkwHKAsCNNM6Fg6EJ+/
VaS1wsiCJoPuZLOyKlIkQs/piPa/joBB5Ln5xC7NcyvSFRAbJhhG3kdAyExmoOx+
Q09sqR3CZL5lzEhgKi3oMwZ7JUOvRY0PPdF/mT97lPSuAWxteo6ynzWpyW9SXblo
0FX9XoEeQD1Kkbi9ndB9UGwc79qFfBVgtZGs7Tg1EMKPcES+sdOAHTP0GNJ2FtyQ
daPoSXo+cIoCVhwqVt+A9A==
`protect END_PROTECTED
