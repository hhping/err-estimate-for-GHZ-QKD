`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SWtXy+P+IB+YThRG0v5hYFH9HaJriyiJ+lqxhUDxn5FQTAk/pdQGDwp1Fwg+J3+z
qmh/z4xHjWK9MNh8m93DcGarLWvQQY08CqQzcGpt0RrDQa8WFKlmCT0rYfxzKWb2
1PtF5CfDo7vL+lyT39/Z9UD7We4G8h6B2HM7HsPwkuS+i/edlUn6ro8Zec/sx2bx
R4YS4hRwHtg8kPuMSgiRH056osv7Ay0z+CpTGptcs0np9w9VPbtPXHEkpai6IWj5
zZrYwI7QhLarRCAi8/G4Weq0KEhGHVqNBFj4KBc/VMuxjHZg80axZa1XaNVdNUsY
3xNbT+910GOR6xN/ftm+t3p26HXhhtw78ROMMcTOCxYQV60d6OFJRc3kP6z4dMU+
JNsfWvfmYuxZ9HczJUO5bz3zLFHKHpRlSGEzHiwsuqmxRtD1Qi0UCOEvkykdqTE+
fLNK97dDHKZoE2rSDffDpDJkeo1viHT864ZQIWh9M3Oj37rEmRpI2aN9wJsR8brw
B2wMtzimQtxkn5XNQDUuAc5OH6zFdwtM5pWxB/6AZp8yglo0nBvmSReEQoByxDCU
agHOpm4rdU0kxkMo/62pBYlxStcWeGAreEmyVd8K+5VRKKhePlLZ5HFhfIrgQPPv
T7PlWwKxTrGxND1NH7uYVRWL893j42aYBy2CH7gDQD1vRpr9r+RtaLBIpEJXoJ+K
NXyemwrplRB8y75YSmlOMr5AjXZzUM+18g9pt+sduWWfYKlcaxsokJjYb+7RInT0
HWKGMfLR2X5nw4hZNucK5RtNLtiYudZuEC59Z1Z+1xvFwtrvlKXS25H2ugut547O
DVbPtKuDoEYpy5iv/dCq4xWnqdeZ3qLY9+wY6YYkbZOihi9BR9JsP2nH8qGIF6Sm
IK32WwyvcFn4PKF+wKumIWkaTH1T1kprU5I+vd+Ti8fbiTi4Qk+7dKf/JLWEzleK
43M8Jwy9fdu10eqHoVjjWEobpZVWUsKRtYmq7E4QorJnLthALKPQ4anXJA/Mf9V6
YF6WHs8XvYZLEsCd0BH5DFLVMIOrmH6G9d6QgifvJr5w0nW7nHww+lDNyLp4BYRM
x1K9WcvYKNBYsX+AWd8YuEpxzNw6YdRLne3VCfYTDYttDW63Qs6ca0Wu1uY9ODXa
NuKYO0n36AIaUezHCyrnJQQt8UUKY+X6bFQG4yDbd55NezzSIdUh7zDJsYp1mBFz
A37SzwtShh2tfMDRaVHddIcByrEE8R+NjQ/IEUSnENPHkMxkEq2Bq1saQh45yQBF
`protect END_PROTECTED
