`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDL0bUr51YG+XrxlbhnFrg3TMm82lwYC6Vdjw1/9FsR2EGzGTmYWhzZaIbfdoWTV
aYT5Rpg3JraYeLPyBhpBK27TOdNEy7SuMQHMD7UgRYo7PTeRlgVIARg0/BktUvie
TOeK/90mN/xUDEVe3AEE2koVBMVOEKL6xbfP+owp2NhufJxbyBLHr18LsR8U/UM4
1rVgnV2ZpSpYL1BKC7fQ5lGM+AX/A55ZSl/5GORokmKHoI+DDSWrvK0+I8ksOPWM
KvWf5/zHdJNFMzmq6REaFsQBkQ1Hgx7v/Worl2LIQV1KzYGGgHCM4um0NmK8+orw
LEBaRoRO8T2SNVOYBoB9TuLTQi8sFAQOdoeMnjpg8BaJkZ9vw4egvrX8fBRUn4gf
/Oiq2lbI8j0fypku7m/sTY6onQHVd++3qfqzAFtyXXhi5eOiKe9oC+CXnV81zlI4
opTVlHXY1NXIc62PPiPJpNiuo9YKY7m7pEq3VB6km+sr5oOzxNSQDTpIl5aALqQD
+bGDTDf1nCcwNY46+aT9otGxXeLhXCl4GV9csWa8ukcKsAyqi6aGJAP9oBZAwKK7
uhriUA1Pfz9NmYhHvYp/ZPrmzztpViuShcJOYA9EIJ4lS9QpQ05CaNdg+TgGaG24
3VZML3lvQZTin1LAZcuz++S6ktOYoTEwwTAkREidYi3NgfNzG2IEmUeBYIWsfmid
7m3hYevl2pRAij/V2aj1QvwSzjoz88IUJg6Blo5wKOj/NI83+Edhis/1caecKWyM
WcNSAjpnNc7mi4LXlV3EP14usDBI5VtdJYl9IbMj0hgS2XSWUfrdcCp4KTE/k/Fu
oYPis5zoKbBlLdmMOOk3MSuhIenIfOm1+a1iH7lY1pniXJl0qakrNbQ5gyMrX93N
bRQIqXtrSUQqNtqkYSD79yk1fprHvONgJxDwHF573Fm/7rNAIvUC5eKOQipLIQAP
if/3UMijih43HDHbS/I8h6neyGg4s9EFP5IqC8DgWOlfYpLif4ogEnZA8agXBzo2
qvrAJzm1gl3NbuuDv9j3ID2/9Y/dqksKiXTsluwZdff+BpABW5jRFodgCWAElzUn
tBzlCnuRl37aKkFBETck5RqqwZwPxLjcUY3kaW37aY4t9BlzmSex9CanKB+Eu3XL
k5BJjK7iKDSZiCRCx7xPoHuMCGgQI70vLvpeZcrkDNTZGqr60Su9e5YxySlUp6nT
GsQRq3TMyVRb5ZxX0idHpc1AjiA3GlluTWaTcN/l43OMh+lSjsAwum8jm3GnlWqh
hKTytVUxtu+BVcdGrKVwMQeROzFFYJrh9SJTz1HzA7IYTcMDbw0hgGESr4j53vEc
JN3VFgEdkTNi80kbStMGzSbfLdZOXPWUeWNWyEmVexEnxhRMiDsxTb+ep7Yz/EsW
kuEKlUs1SB/kS11u7NkYLXQRMRl1JP9MGq+5gTpd6WA11BZi9oxT/nF5gjvd9Hy/
PLn3HanaRu+mUP+ITbffUyC+3x97EXzwvIfmkESm1Q1fVIvjdbeEqaox3c0MbvMk
ENUvLr92E+Mv67DfsQAPkYyGoORk2u8FB1bWAYzEt7P64rJzsNHJrjXd/tj01PQB
ymJ6t+2ZUq3/djFBgQa79e4YQLSMQ4h6oRBcxDoPwOa/3zTMZg7CBRfsD4BuagyR
hSZVvj98CHBTCZzz7/RMEXdYqgmCoQWyS7bHf7SULdQ2ELbrTvwS5BSjZ0Jhz0Ah
4COn89wjKS3UcYn73ASlAYrIjMjedMlsSmYQghfqKh1/OL5fAijBmAemZmPov+VK
quOklZG1QVDIviVempmnrz75tFesiQJU2w7r6HDlu9t3FQkoBDLact0Hl0aXzbds
swutKvrZb3Fct4vWuSNSN8JDYgV0FkVj+f72PAz+gMpOSQrOv+3NKlcCQw8ih/mq
6/73zduyqx+kJKXf6XLfNx5f3pKj0B/bKFfn0uQHv+gjevZ0ywpiYOXQqcikQbjA
xiGjlhpj9HlKQ3vQJyKtHxFkwRunm8/+GeXNnJnIsMVnaLBoykraNyHxo1s42bog
IvhUTuZ0zNrIlCQn1kZIz9f+2ZTV2Wwloedqp6K936kxkpIEIUXsEtKFU40/wF1C
x0as5O0XLdWPSftdnnTHYu68/iJYllWi7OBuY1Es9LbMAhk4ws77df6HzPGTsWDE
AH1NDpqaWn7T9q2rRvCc4gHIjyOxQfWARUEDC02X7Br4guV/7OXRGeNIqL7oYTyg
afeoHes/t9nNu0ZBKIkWNene9npkgPtuE+8RCs/4xhMU31AQs1U6KJEX44dCIu8R
xPTK0qCq7ivQ/UigrGWSK50T7HIASY9klf06cuI7N1oGYxgeiFutUc+Lo2Sb+VUO
Buc83Gxm4n89yVIObIpdx2hYH4xkj69txGqFmEZnJ8wXQqF7EouWVHYlZ8Mc5IMa
ldKPLh6lo2JdGwFLrzVl0EYR+aptiLsTYi4RAA/I6gcQSMZGDQEQhZtrte4psLs/
K6A6Z/sBeo3VKtck9O6OWHy+x/IzhjfoCiECt2edE4rOF3Z+ABO+glKHe0kH6ypn
RprX2AnxukvY21/HisIv6DzEY8zPdiaUkHKlko+6rnbiUm0ZBZNzPioZDdxiVEaP
67beAVZ2C9xRNjogEeAME3knjFZ0G+/rlLoQz0q6fLC1rt+BMsx+6ojn8HR2ol++
5E/SjvgvqLbD98JZxiEv4xOuyslm4XCb5ykVj4/23aqYbEOJ8rYN8TwpDCAMcEnD
SKWRsSDqhIoqn9sfdb+AINbiXcvdsX/9hjbRzH+auJVCS0cOug+qZY5F/Q6k0Ujz
l3FwL8wGQXMbpFnCu9ij+UyOOMPG7ZgsSquVJdpQPMjHXvK9AMip6SC+YVpTxGsa
rpNsWLjHGUHlvTA1m8AhiaWkWRMi0IavQfAq+3P4rVbUih7XHafbWKRdLTFnP0jJ
sdDG9MojydjkPUIY0ZotVqRUseswEf/xZbgUVRbFAMpXzWJUTQ4CzM3cZnAdc0BG
CJt8fEruMo1PvLWyQ88denrgtrXzPmKP4z8r44z8Hz4reb6laZt/vbTczxF7tgPb
RYP8kExXZNnuoCq6lxDu6dma8YA6R6wifeRZ7honz6W7iUEoO9jIn71bMqS07bvK
qR1Zv+P/cYD8lyZ9z5NebocfOuOYrPmIoti+FMH4VRg3TWJ6d/eUZPJSegRT2S6H
YE9HC4PQtKjLMB9RvidkJ91OeqGjsORGOVvhPUuLynYJjv/UWFMmpsdHu7D9Lj+i
L+adi7NHHM/2MqOCUldJz8Y4rCQ49vihi8Cda4933D/FcOrTa70WTvMIIHVW4o5a
CIniWgraYC0vI8Uwj75L05lGjths7LNDFYibTvV8X78PEftDyf1Y7MVGLSDoDG3T
eHc+seEzjWtYRWtGL1O8hDO4gnCksm+cy3Bh3q4q7PwAuN2qcBrvF1XeB/NfqIS3
8WUzV2Ml+WwJnofrcU/i6RUPBxMidWfM6/mgPlrJq6gXB0xW6uJdUhEx/R6l7U/9
5BWigvAxNCeo6D+hkp0plgJmu2ja5ZzXI0Zg7ukDQ+rh+nd2UXgqWS2AbH8/zHek
ygg8dBlqNxT2S5uTTjRg9e5XUC3XIlTIH4MLhRQQjv6xGlcxuyN6izz41covzi7P
JhJKhzZ36IZvGRSagu6YJuL3T6J5KnNOz+AabqcHpMojl4uCEI4qJDLZwOIpxbxq
r3ZqxQHxCpnE8Jg4oaALxfJuXuZa6A9OZSqoBdOa7iLOvFT3RCyQ2lBo0AjUsTZ9
YLzHJU+OnGoEI7fLL32HgShBoUVSlA6W93BwTYaBTmqQk8C0v3nUWBPwY4J5UTmo
SbDkDv5K5Gc2kJgNDbJHL0Kji05v4qkBwAUhyibBd7rU+UKjihVrjGTADx+2nXis
Ffl541KDFqOsxtBNRkhFAwtPNVc2Z6CQABermjT0qVLc97qFpYrYh6sNa1zbNLL1
wD0nlR+Rrz90EUsRSq7/qDjWa2oSFCdK2dZMs7AtVj+bAOYNczquoZGFwcoczoEm
ezkU/bW0hoa1WpEvK2ieovk+7SyEGFyPQCxVWj9C6DyqlmZS74UnHUjTZjYXqJd2
x004yZvpnKeodHuHgn7WCFIz/GOLY5Hj/uR5D8Mp4EBjuiP8qp49CzTlpaMru+BX
nEShjfd0Xico0B8u7WSY+FFh5HNeTZjq93ueOfiukPw7aRF2lhqhgAFUwejLpLiC
u+VWs48OECkS8cMMD4lYh/QMRwobumYpbUUnfCyvUgAlqVoRHnqVEoKiX5Pwcd5q
fzVTvJHRux39e5kljt2sDTYZ+2QHYX5vHWdk1YWQOMaP9jmx59d+2Y1vTADkgsyL
YqHH6dTrmCujIk3tdk76L469TFtw1+DCI+Qw1sxauWTaQqivt980B2V9GHwHh0Le
oZo8JcSUPWnwBKLzH48ySdgcJAJ+sY2J6Jz09N89+7mODKd2pmkDC/8c33FcanpJ
peaOzpA58ucR3ogpvIG8eGSPJ8epMiLVCIEXEOsbO+pLUvpcV0t3K8UPOePtMNmr
QfDRiMsDQQy719kNtLrJfSffvXqw3RX/vBDWheE7gtRsvJnQB6ib32n5BHHrk90K
taKvotXOfOvl0X/4MXsYiqDshndrgMquy7xilEcFrio5VDCOtGTWvO8yp/qRRV99
kfohvdR9/yNZcup0N9WmLDnlZQNP9wrnhvXFrNF8WzG9VFcnNxlbfmt0JhRYekE5
xlPHlDLKHOqq6jBBf+1L2ph7si/DUI1BqqpCPt7+FRrOk9mNceNRHJAhhmc3SJIh
G9dAJtb3CdgsSRrV9BFyU67Us2rcey5ywIeByQTMB5yuXo+FWd/TagTMjotIxh18
FBbvB9e3TekKdBpbddRJuVotW3wPRzidjIX0tR4yj7CQGWhx//lLF7V/kgG3fETB
Ou3hCzRmNmejCgz6sQS5XvxJkz1j5+XuzMwzrfV6OIMKOipKijZzzVyvl92o2rS7
Gn7aVYCs5wSCvSshY+Pu7t0XPMjVLjWDcSX+KUw26c/sR2H3uDhv+sZKm5u4PTKT
hkVS0zaZBbb22abMl42ovh84nRBAZmJWfd9oKvlqRhwxHnVN6Y1FQ1cu9WrbTY+p
QcoUJNUZfFqDFOLQ5gzgapHNrYIcyQaMKR1oRcuuIOyCnGPHQDGtzRSqCE/drSrb
BuG55s/dq1lygkrPe1bA9Q3/KlPUjKXrJerxvjag/QJ+cUtt6dRn8RqpGIWg0Ru/
BvwB0T+9UL5p+02qVcMKsZA5mD/dBOU6xX0x4daBvJVE3Cq1R08HOjAzugwhfMif
V1uxGXJ+FUL9gTbpowUFEGyWwiuT8h96iZwglOPyrFhlUb4ea/+P5WHKOGPXJlQ3
TyPXY57YtcBo0CTSIpfBMm44TL3CrsIF2VrDqFcNWZBoeLN/bKka4vokspHZihrJ
Yh8ZqN8y/+8fBJ0LWare7sH4IVGQbwaQQ5vEJfqwQReAl0vw5De0IsOxZPEQKutR
BH+T1Z3uJ5jjyKTB97S54ke/NzjhuBxB5RNRZt+D0REeaTYjv9BTtEz+wcz/KnB1
LtyqfKKp5d67dBko3G5eEykxJtGvhyUapQl5RjWw62w=
`protect END_PROTECTED
