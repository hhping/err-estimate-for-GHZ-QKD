`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9DLBYRFNNzLTtqv7SaglFSpLvtHRPb5r4eEhGEh70fBE2l2Rn1vOt8fd3ont4BbG
+h6L382fhEm75EnijubvqjznCf17gUuMyO0cxk5O6CO9l8yyYtFuDf7vaWIKvBTG
Bzp1z409QfiLdET4ehspQfDqe8XAPuArVZz48PVF5Od9pp1l6RP1C5HaMYq7eR8g
UHssOXHF9CSe2UjjzrYp2m3WUnArNue+dqJbWY+5K6uXHLHL3Cpl/yiLWVtpNK+u
egdtjU0vMFmg3a/wxliPluQtbVxl1mYJkGsvpgp8pv+mSd9RaxYVCDk6ppADfrY5
n9pHOhPH9WVXbLFuOtgAoZlKXC3HlD/h91PWOVhcSlYrkh085IoYl6PWTQ8FjT3f
9o/tboB0iHRGEmsu9naRh/vhZQ5UM2zDEYhHqQ+YmriTKdZv+0uu7UDM4MFyNngP
RUGahNtnJ0zbmIFOA3A1TEQc+RH8ufXwvrq5HUxY/oxcN5WhAWIU+TIcUg2xvYWh
xtMbfpVdFqfTwZDFk7vXlfqyHGDWjTxtfWYwWHeMu4T2Yfe52p/PCWeNmL9fyN4x
NldXJNgQY/Zgl8eDB3ggIQhpVwUpSlOXFIGfN0fqoCvnW5NJ6ftWSPx17gJ1+Kwe
MKBPmBylKbg0LsCCXM8r1FvgIWMjJSW/PL3/kiMBo3kMAEcBFO2/YkFR0yXtO+Hd
IkQuhl+CC4NFf8d9qOjV94gOppNh35/qiSS6PGmBEv3Mbl9HVcxeTe/GRUpJhyyG
UFVvjUvJTlbjW9GyIVAXWagS3Fm2QmaPiK5tUhJfMGnYXbewxbJvlFpa6ka35URh
oiFQTE2OlyAy2eTg/d6SHsyDfQ17tKCh/Jzox5lLQ1IVoByEU1Kn2WQuKSPJveKH
jMD+qV7L/QvIAkY4Ae2W6s9TBcfMQ2oeCDCRClOTEuN6exfL62Bo3sc2uaohUUSJ
69FGjV/DhExrRIL9WrVEhb5Ynd6DSDKVRTG6AgMiNS9q/mqMtj18tsjHVvm0ne9F
52N4HZX+XFq9ONfIqnxzuap8xS/+Vbi6sr0pffsJ2d0aaU9FfYe649zPECnQsWXR
+yGfJQKNC3SXvCms0Mnm47zEz9WnhMSjcweKsXCbbN+gWYJP9Frr623eZP59oGV9
aM7Wc6ANf/QBmoAC4OsEmE+IG30fawAVPgfWY7UnFl5gzrQNP0krmf9UvesBNMvh
IubMcH1uOHC/Clrgi3UbQ7DWiM9GrlV0ZcKwMxl+hffuOeOp/VOAtESldoZ23bSe
OHKKBVxrVoCA2mMHlgoTAguemBb21YLaQIhwMFudEWamhSqssLKNQfb9T9F6gkKd
VwyCz42uNirfqXMoMehFAJ/p5AIze5XH4oU+9LZaRj5R3iTZWMdosMVASpXjDz9c
5+6Y0R9q3h4fiDpucU9q7k8VkuamR8POv8bsjhEhntNpFXceAUGDUPj2ehEZYV2B
jSm58eu5CgfjRNScBViYLVLBaXRzMevbIPq4+m8X+OFn1wHm3Y9WKw3LxOrS1dZ/
SeF8bnu1zKamyIZVmvv4wUQTWker/v+WAYLzwVCgtWAfxZXIjRzFH4WTDWp3ZRCD
pjwjCGm92IzQ65uY7cVDf8XvYX4YSyvt/4wwnAnFHKNu+IRHYS/CoE5/0HLzKKVa
9eKsJMtBbbR2BRaun7r7XvvEnR0k7DhnSjEL+mHhIRxMCxFSms84tRaGjJhBQJ5L
CUpnAYtDVb8rqEQAzmGIOJz+XKV/Tu/a5NZoN9ZUIkSZg+fSKTJxj6Slmqeft8xB
4Xih/9J4cF3tIOtRPG+rcm4I23XpBGnl+Q1LnwJxSX0DFfpap9NpkS8ilksgewbY
UJnB1x9XceYdoMfC5Nq6cGOIZnKwfnMUigAu69rbkr5YqLrKS5+otG5luWqVgzR+
nNiqbpG5/1zpvYvrC8slAnsLKAakjrdDOknYxmkrtsREPikrVlx2OUFlk+8SnJw0
xhCBoL9L4vOeE6LZ5/luZ2i1gHOx4gtV7Rle3dPurDJuTzKeT6SbR0FO0k5zTYAP
2RWVdDutsD6FbZYE0+VLe3QNmmVz5AroUz3jOdqr3pEjmFZ55fUt+/qKT5DIerMf
RCzaiX8GoQAgrT9lseLSW1Jb+O0Qys8Vh2mKStMclO+ETQR7to8Fn6XLUVE9OrIL
8SVrTjQyZwhJuy6cIWqxpVW3487sXO6MPJSPOZGGI6nuENld6IXLsP8U12rNUxOK
dh6evUR3xkAV+212K7IRVprDQsZza/WEr1K0CRqXnj6OAngt58K/xBI2B3KUyw5g
`protect END_PROTECTED
