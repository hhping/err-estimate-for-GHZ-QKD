`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xz6vRAs/1qidlqRDlkJQRvB05Bjmp9o1YfzqwnWY2PHrfOyKYURfp68WoiJsTsBg
X6UAY5o67A45MD28mj6iQa0MqwqljKz5yv2KGgM2MDOVm2cSKgACDd31aw1BJcwA
yYo2cy7OG7bv1d73s5LkrgyBFcquSE6mUG6hGAu0XAH2IWyG9OfJsEP9Zd/iuE05
1rMK23HA/4YMo0cKbLB2plVWQX6A/5VRUuY0UtmgT+xzdRerGWRKTbG2Ejt2u5mJ
MHtlO8rumnVwzjvKZS/Yy5xQb5Emt11gpn34MTVR0KMKHKw9FdcQ3xIg75YG7a/y
KEnPi7XdBh8fNjL1PCVcWOwr5znNASrgHyItgaGoBSbxbPSHDdftZDFG60vXxvdS
FyrgZvuYpEz/rsHUWCTCD3LB8nLZ0BJ6OiBQaMvH8Sv0dELzZ8/5h1BpiG5BiqwS
0hsI1zsdTyZ/vgacg0sGPmjrjVI3zX0wfwgbxO6faBdXSzTCZNAARKTXQDHq5IIX
s3AGP+DRAooEpKDnkC24NuMsEcR0cbqgjoeRhlkRAtNVuCCQoetJJDVTIaFWcuME
jidgWtJeUJtu/HL8x4y+zWhWQKKY8p7/7VCotbZRZwWoNdUd2RQ0p3rkJ4gyZym8
WCyYtXQPIpUFO/Cpp+JvQulm2l0lCgNqpsJ076aBL2WKgl+3tDXdJoW+SDBeHk4M
ZLzYImbwZv/JOEz6v2fHL3LLIZaKSCcz2uD+E/q5R6o=
`protect END_PROTECTED
