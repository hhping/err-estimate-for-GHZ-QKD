`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klTbwm2nnICKdmdnxF0+RtKhJtuh0al+7rZiS9Ktnfa3h+MFB6bbJ/+kSPOwFZED
HmxvvhC6pjvUxHdP9t+N9K+3mGcecdS97+oa8+Pgp2dyjuLhwSryj2GwzwNrH2ON
prhnczwcHdyOqt+sbM0fY+pMt+Epnbpz917RTFbYOW/TXrktfPRZUyrtRZ1mC1yN
5mMSN23rSEy2ay4oBJpPTw78dhX8hOQdp7Cp3Xc/rg74MYK/yWnWHK661g53Ry7/
OUSBpACKkQaidHaFpx6b64bTyKMovD6qvV7J0mPtLf6o1XnXwYV2uOhCoEcbaGrY
Q/m9LAny8d7KB484TkAucbIXEHu3ofRwFhx1MUjXZsdloZcbiv0lzMkHdVwF0rT0
a3q/9+ZtA9OvOp4JxyAvUcSdl1pAaNKUF8wGUbYr8RxmEY1TB8CBNpM5nx9bltXh
QoGi7cKIMDsa/buvCsLMXPNpXW0WNsHcZwR7SbCBEc7u5Y37cRVp0st7EbpttyuQ
4UYQvVu8BZt3EWeSWDYPJLxING1gFsf0Zjvi106rReF8XjXSj5SsrFe5hCpbSg8e
dGsCD5gwbBUjaKLwuWnaaGMSmisCuAhhOQxZMOL9RilxbxayRtQbfF41y1rmWo/4
EpQqf2Hr7dJ6fnqxpEsgPy4i/lJOv9huiz//i0ECLzQ=
`protect END_PROTECTED
