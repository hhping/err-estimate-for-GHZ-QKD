`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjcLFLiuhasqGLXc3APhSMSuMeBFv8KKwnNdkJhjdNdb97iYySSCWQUa4Mn76FNx
ukv9RXCuc1D9FIvLOy6WauWlF+Yotr9+wa51FEc5Bm2+4ovTKTmH3J3hpUAPAoEj
rm3e0KGOei0F0roToESNBPq6qctxDrhLRf9VTSqCIwbq5yaCuVlS3cRNPPiMGZte
sCHtL7F0adjV1XjbyrZxDYEC8wn4T3UF3B7uLJ2+CW0C5HkQqNMmYhN0V/MDRXLg
WmKShw3jkdRXyn4vVsFkg9Y/u6p4eo9B7Sb5szgrr6PTGx3oBEZbQ9/YGFYsQZ0z
nOL55RAip26ktRXpnsMcKYUBnz7CtkrFaoNxPzwyM12q9R1SbFTmkhZXdDd3+TLs
OXtaLzrzX3C0TcPHwwD6QpiSdIu0if27Mi3sYf8Qx++aTAuGgNmb3HcuXgHDeWRr
d++Q/wKrS2lil99LS2qVngggmc9gn63LeHgToVh3KxQUwm+7vx+Z5bwYlkSPLGYB
6D4pEDwFLbxyz1UKi9b70Fk75H9oEXpRT26eGU4kU1sD5u4W+R46OFKS5LbTKN8r
/dwAWWMfdmwj5KdsPg8M9AJlxZecxgszcj1Ok1FgzfBIjmBSLGAEt02v3UB/KW5Z
KlezHoYcnaCChvIzJIIckF+fKquZpZbZ+AlGvogjq2fQ38hZldnSMHpu5qgA5sLf
PGHNEMt5LsKdxDa4p1/drmmbkpjz6thFxj+VZKlZFWWUFDYnwcrNzMZjz7J+viAr
+zddB/Y+4WxWU5TDFQlJAw==
`protect END_PROTECTED
