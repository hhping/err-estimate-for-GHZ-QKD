`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgL1H9zN8u7/pl8RzpKBO5j+y2nFi7VIiMcoNyoYE85Cn82gS06aA2BQaLiM/1tV
kAOLUTCRxh0nyVhHXYfM1I8pW0vK2aUNYXTHeJLH3e+G50fCQF2/LEmSR6WCmgNa
+Ma9f/Tt2W1P3e2TnQFqwQ/ukfnvYEm8bc9sV38AXnjIWXQM/mW5vUfWy/1w2oIc
3DU04CdRB/UoeQ4LuQ4oElikF7AwbcwY2hFEMlGUfcYH+LBlEBldx9ghm5Mw1Q1M
dykER8ccfJ1v6243Vl5uspmTtOBDs7mvMWsJ9QlR1wKxir8YXnbHboDbjgwlWCaE
GcN1PQ7+qSmMAJQpiVLF0D2RMZZkRp5k99b0cdHI4b+RLX2oH7zRQBmapMN/Gbpe
xV36PRKGguEnXC5uVETEJ5ryLqZ1Y1isCyeBE+5G7m5G1mRIBN/2ilwxWwWkQtrv
s1d0NY52X6RXg8e6g35UlX14/WtEiXHqbsmCvvX3NIwVCDpNHDp7iN+Mz1p5t1T4
LmJIS56Ihv2PcYEJuI2kM3zeBJrUXseMQC/i+2dJlOufk5DEoqpnmCsib9WIJB0l
LoQarTc4c7baFSnJkjuppDOpNPwpE/qhjyx9mgtr28Gp3NSSg9sUQHCedu8ii2jF
eSIZf2GJbdiiNYSmfHsJf17TdiGw4Uka9z+0JYQ99Lc/TxJazpPqd7JoiSD7bwPV
zYNE6fVjeaFLrsmU2i1WLRa9Bu++hXeLkRYkCZgZGQHfqT5VMkiAU3/nyq5aM8tU
UJ9mScvI/j9Jhs4DBACcqqWgdUfZI2rCuOCOhNcIDFMYdgODEFMb5ftRIQNJpf/L
npx+PAyl9pDb/+ainglX60vqsMIh36lWc9/N5j4lcjvagsDunMoqIsRitCLUyvdV
DzY4nwQ661QrYJVNnITiVtnsdo0fO1MmQqAwyWNiMCVliftngwAl0FOBzdI9735j
NvQaI+wzuYgwYmC0m37pM+fU9cCF/jzGRJaiX08kZySpyLbZwI8DrSTXm3OxmuwR
y+NR5C1HC6pYDsqpXiRW1VwZH5c+a1FTN0y0lhLCfYWwo3yqxb19APGFEDmqJf6S
1GGfXdtDRV3ufrmzVTx8Ys9zgFFCYpeqhnlxaBzSQcfwNf56VbDoNY/SgCsaFXN+
EknZ6QC/Wl8ar7BMbpIVMe1gzFyBK/nEIUSzte0NzMjmTv7+axtZ0aGMHzckE/Qq
dhn6x65V+CbZmuYUk/yR3TPIivY7WxGzfZ0EGErFUc8Zr0i6T3l42T1Orja0srAR
2gaxFRKlGX5oTOpmSTSqSqSivmIT/7K2Z2VIKDBkacThhzETe65Mwp+Mu7MVRsyA
PstPp9suT7vaBbi7RlGvBWTyMa9Bqc+oLhC5nkqJAa+DD9rSAUjbanhbXQWurHkW
o2AZTCiWqRC3zXPqS0LjD6F5EQ236G/zbeT+L3P7bQ0jC7P4vD9gDz1FPhAxdaLp
sZtVQT8oWMQC1Ao1H9Jy6rMydRBV1pnnqTogmE3odsxBwgi8O6ycuVbgUIkSus6K
cJv5rCYQLgylpq2SFjv/7Dbr6t5Nu0AIMiVrei5Fxy7CJGEi9p1br/v+e9nu3NF2
PtAto3hOIHt/GyT35ncd7FtvW+vaqwbOunHHA145vfsxwElg3TKO+UIEOQeLqCQH
AjV94YWtpfFE38yWD1pFz2NgPiOs6ZWvTMXoIvBsBK7flv2E7XHBZX5XjuZeBfDb
OzqysizzhbvM8t2eEm3G+aVxaNCFVo7gqcCHmHwby8dEkKamHAZLAhUw4B6jJ+YD
TtvDQwAAqnrw6iH6pvD42PnEWAqyNLUdps3J2NVeYZwFPGoPvnhka8JAbMNifKin
KY8KV9JWQBYVu/D9aTdgU8pJ5QAc1conOyhHxy10tgTTPclF28w1MzvpuG7XLTm8
q6QGWDiVUnSxqRNhGLBqYeYPv21TcGk2CBMwkJeEY0g=
`protect END_PROTECTED
