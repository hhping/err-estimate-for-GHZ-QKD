`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEfJfbN5az4nk5DMDfAFqLjdIBehsw+V1abF4ud9G16nJezyLL8vD2xIAToI6c7c
IW3yOCGbRWy0BoSIcsPYxh7MRdPKxX0L1n8GhzQprSkEkURjDlBwUjLyCEeQyJEN
r65WnK9JMQkDyqYqs8PDpjEJ0YDXiTHv4ldp5eBVgl/KCLPhBdjmPJOQ9t1DG08d
JQz2aKl0eAFEErXNrSitOuugjdQJoQMn+mkc0JgmSvpxpTi4g016/hIuzj4d2Eir
KGwdNbuPylwwLgR3+IX0Na8kFC74607geIOfWkardyXiq0etTde4IW+pkS8X+629
x4bWaj8pT0rL6sbe5Zde2uWGlAjTu9VnTCuUr/zJsuRa77CI65iaLEN/QSpYpHX5
BP3FWCHXfJeadRDgaebjT9raNdphT5RNGIoNbcgqwd+gi66kYFB/MmDIIsPBJ8jV
GhnAdbfLTcnaNA8mqKtxolAY5odRPsavWzMJQcjhjM24Obpei2Pgn0cQhCstlKGw
08gNn46O4wKykaToCRmYR1AdlggZr3I4/86LfsEYgoRhlRNQ7HuQc68xSYfxfDNj
`protect END_PROTECTED
