`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRt4FjbfN0EIhc9KCJ5Gmnkvnx9VYjdnv5kZyQnHr1zMFvQvVAHttngRscBiMTSu
9B/D/0FQIGE+FcN+HGym3pV7QthAC7VmdUB7rYlITLmO4Osy30SZ0vmUaGCHriUw
SEzh8bBZmbi/Y2NIigrcZsmOOmehla8CP4ZFfYN8sE/3wbz8lbblY8hWBauTrReF
irzzsEVFJn0XnaveI9rhUyKGhduwNJ7fs1+pt2Fv1iTB/DR8DpTZzMv3SUImBJte
MrJBdpwQp8szEBkB2bfMRsPR1eedvR2ecfA2RKiZ6fGyLWuF+nHCRPB8NEA6YdMl
wY9fDcA5O2g8EHRkHjKKKJ0I8ZGzF7uJuIdi1O3DfYNlidg7GOciygxn7qtGHFhV
Ya5IPkwvBEHvQjZnZvZwDHiJPaYFDCO23aVlkDB84qzssrBtNigBAK3Rok0uyBl+
x9m+GmQh+2GW3PJbdCqdiag+CMSntIjIe40oqAYH//DxpPVrtTcQI/b5+J8jTZBg
RTr55H7yju0zRc0CqQK71aDbfSWU4QV3T/7NaJ+KFZovP5lBqm9qMsxTF5L86Xzr
GuV2m4QKiEqEsiBx6EaDzaNmZOZFn4P5KHdNbmcK0HVO5/l/jEH616dtVOVa0eXE
2zX+NgYogvv0U7cEmtkzV+lPmmHJ4lsYmzYG4eIISfMb7VMcMAjqSYQHw6koPqp8
cLlc1/h4yS+X1UrEQyV2xQ==
`protect END_PROTECTED
