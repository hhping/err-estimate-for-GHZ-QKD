library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_common_pcs_pma_interface is
    generic(
        enable_debug_info: string  := "true";
        asn_clk_enable  : string  := "false";
        asn_enable      : string  := "dis_asn";
        block_sel       : string  := "eight_g_pcs";
        bypass_early_eios: string  := "false";
        bypass_pcie_switch: string  := "false";
        bypass_pma_ltr  : string  := "false";
        bypass_pma_sw_done: string  := "false";
        bypass_ppm_lock : string  := "false";
        bypass_send_syncp_fbkp: string  := "false";
        bypass_txdetectrx: string  := "false";
        cdr_control     : string  := "en_cdr_ctrl";
        cid_enable      : string  := "en_cid_mode";
        cp_cons_sel     : string  := "cp_cons_default";
        cp_dwn_mstr     : string  := "true";
        cp_up_mstr      : string  := "true";
        ctrl_plane_bonding: string  := "individual";
        data_mask_count : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        data_mask_count_multi: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        dft_observation_clock_selection: string  := "dft_clk_obsrv_tx0";
        early_eios_counter: vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        force_freqdet   : string  := "force_freqdet_dis";
        free_run_clk_enable: string  := "true";
        ignore_sigdet_g23: string  := "false";
        pc_en_counter   : vl_logic_vector(0 to 6) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        pc_rst_counter  : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        pcie_hip_mode   : string  := "hip_disable";
        ph_fifo_reg_mode: string  := "phfifo_reg_mode_dis";
        phfifo_flush_wait: vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        pipe_if_g3pcs   : string  := "pipe_if_8gpcs";
        pma_done_counter: vl_logic_vector(0 to 17) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        pma_if_dft_en   : string  := "dft_dis";
        pma_if_dft_val  : string  := "dft_0";
        ppm_cnt_rst     : string  := "ppm_cnt_rst_dis";
        ppm_deassert_early: string  := "deassert_early_dis";
        ppm_det_buckets : string  := "ppm_100_bucket";
        ppm_gen1_2_cnt  : string  := "cnt_32k";
        ppm_post_eidle_delay: string  := "cnt_200_cycles";
        ppmsel          : string  := "ppmsel_300";
        prot_mode       : string  := "disable_prot_mode";
        reconfig_settings: string  := "{}";
        rxvalid_mask    : string  := "rxvalid_mask_en";
        sigdet_wait_counter: vl_logic_vector(0 to 11) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        sigdet_wait_counter_multi: vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        silicon_rev     : string  := "20nm5es";
        sim_mode        : string  := "disable";
        spd_chg_rst_wait_cnt_en: string  := "true";
        sup_mode        : string  := "user_mode";
        testout_sel     : string  := "ppm_det_test";
        wait_clk_on_off_timer: vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        wait_pipe_synchronizing: vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi1, Hi1);
        wait_send_syncp_fbkp: vl_logic_vector(0 to 10) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0)
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        int_pmaif_8g_current_coeff: in     vl_logic_vector(17 downto 0);
        int_pmaif_8g_eios_det: in     vl_logic_vector(2 downto 0);
        int_pmaif_8g_pipe_tx_pma_rstn: in     vl_logic;
        int_pmaif_8g_rev_lpbk: in     vl_logic;
        int_pmaif_8g_tx_clk_out_gen3: in     vl_logic;
        int_pmaif_8g_txdetectrx: in     vl_logic;
        int_pmaif_g3_eios_det: in     vl_logic_vector(2 downto 0);
        int_pmaif_g3_pma_current_coeff: in     vl_logic_vector(17 downto 0);
        int_pmaif_g3_pma_current_rxpreset: in     vl_logic_vector(2 downto 0);
        int_pmaif_g3_pma_txdetectrx: in     vl_logic;
        int_pmaif_g3_rev_lpbk: in     vl_logic;
        int_pmaif_pldif_8g_tx_pld_rstn: in     vl_logic;
        int_pmaif_pldif_adapt_start: in     vl_logic;
        int_pmaif_pldif_atpg_los_en_n: in     vl_logic;
        int_pmaif_pldif_csr_test_dis: in     vl_logic;
        int_pmaif_pldif_early_eios: in     vl_logic;
        int_pmaif_pldif_interface_select: in     vl_logic_vector(1 downto 0);
        int_pmaif_pldif_ltd_b: in     vl_logic;
        int_pmaif_pldif_ltr: in     vl_logic;
        int_pmaif_pldif_nfrzdrv: in     vl_logic;
        int_pmaif_pldif_nrpi_freeze: in     vl_logic;
        int_pmaif_pldif_pcie_switch: in     vl_logic_vector(1 downto 0);
        int_pmaif_pldif_pma_reserved_out: in     vl_logic_vector(4 downto 0);
        int_pmaif_pldif_pma_scan_mode_n: in     vl_logic;
        int_pmaif_pldif_pma_scan_shift_n: in     vl_logic;
        int_pmaif_pldif_ppm_lock: in     vl_logic;
        int_pmaif_pldif_rate: in     vl_logic_vector(1 downto 0);
        int_pmaif_pldif_refclk_dig: in     vl_logic;
        int_pmaif_pldif_rs_lpbk_b: in     vl_logic;
        int_pmaif_pldif_rx_qpi_pullup: in     vl_logic;
        int_pmaif_pldif_rxpma_rstb: in     vl_logic;
        int_pmaif_pldif_tx_bitslip: in     vl_logic;
        int_pmaif_pldif_tx_bonding_rstb: in     vl_logic;
        int_pmaif_pldif_tx_pma_syncp_hip: in     vl_logic;
        int_pmaif_pldif_tx_qpi_pulldn: in     vl_logic;
        int_pmaif_pldif_tx_qpi_pullup: in     vl_logic;
        int_pmaif_pldif_txdetectrx: in     vl_logic;
        int_pmaif_scan_mode_n: in     vl_logic;
        int_rx_dft_obsrv_clk: in     vl_logic;
        int_tx_dft_obsrv_clk: in     vl_logic_vector(4 downto 0);
        iocsr_clk       : in     vl_logic;
        iocsr_config    : in     vl_logic_vector(5 downto 0);
        iocsr_rdy       : in     vl_logic;
        iocsr_rdy_dly   : in     vl_logic;
        pma_adapt_done  : in     vl_logic;
        pma_clklow      : in     vl_logic;
        pma_fref        : in     vl_logic;
        pma_hclk        : in     vl_logic;
        pma_pcie_sw_done: in     vl_logic_vector(1 downto 0);
        pma_pfdmode_lock: in     vl_logic;
        pma_reserved_in : in     vl_logic_vector(4 downto 0);
        pma_signal_det  : in     vl_logic;
        pma_testbus     : in     vl_logic_vector(7 downto 0);
        pmaif_bundling_in_down: in     vl_logic_vector(11 downto 0);
        pmaif_bundling_in_up: in     vl_logic_vector(11 downto 0);
        rx_pmaif_test_out: in     vl_logic_vector(19 downto 0);
        rx_prbs_ver_test: in     vl_logic_vector(19 downto 0);
        tx_prbs_gen_test: in     vl_logic_vector(19 downto 0);
        uhsif_test_out_1: in     vl_logic_vector(19 downto 0);
        uhsif_test_out_2: in     vl_logic_vector(19 downto 0);
        uhsif_test_out_3: in     vl_logic_vector(19 downto 0);
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        sta_pma_hclk_by2: out    vl_logic;
        int_pmaif_8g_asn_bundling_in: out    vl_logic_vector(8 downto 0);
        int_pmaif_8g_eios_detected: out    vl_logic;
        int_pmaif_8g_inferred_rxvalid: out    vl_logic;
        int_pmaif_8g_power_state_transition_done: out    vl_logic;
        int_pmaif_avmm_iocsr_clk: out    vl_logic;
        int_pmaif_avmm_iocsr_config: out    vl_logic_vector(5 downto 0);
        int_pmaif_avmm_iocsr_rdy: out    vl_logic;
        int_pmaif_avmm_iocsr_rdy_dly: out    vl_logic;
        int_pmaif_g3_data_sel: out    vl_logic;
        int_pmaif_g3_inferred_rxvalid: out    vl_logic;
        int_pmaif_g3_pcs_asn_bundling_in: out    vl_logic_vector(8 downto 0);
        int_pmaif_pldif_adapt_done: out    vl_logic;
        int_pmaif_pldif_dft_obsrv_clk: out    vl_logic;
        int_pmaif_pldif_mask_tx_pll: out    vl_logic;
        int_pmaif_pldif_pcie_sw_done: out    vl_logic_vector(1 downto 0);
        int_pmaif_pldif_pfdmode_lock: out    vl_logic;
        int_pmaif_pldif_pma_clklow: out    vl_logic;
        int_pmaif_pldif_pma_fref: out    vl_logic;
        int_pmaif_pldif_pma_hclk: out    vl_logic;
        int_pmaif_pldif_pma_reserved_in: out    vl_logic_vector(4 downto 0);
        int_pmaif_pldif_test_out: out    vl_logic_vector(19 downto 0);
        int_pmaif_pldif_testbus: out    vl_logic_vector(7 downto 0);
        pma_adapt_start : out    vl_logic;
        pma_atpg_los_en_n: out    vl_logic;
        pma_csr_test_dis: out    vl_logic;
        pma_current_coeff: out    vl_logic_vector(17 downto 0);
        pma_current_rxpreset: out    vl_logic_vector(2 downto 0);
        pma_early_eios  : out    vl_logic;
        pma_interface_select: out    vl_logic_vector(1 downto 0);
        pma_ltd_b       : out    vl_logic;
        pma_ltr         : out    vl_logic;
        pma_nfrzdrv     : out    vl_logic;
        pma_nrpi_freeze : out    vl_logic;
        pma_pcie_switch : out    vl_logic_vector(1 downto 0);
        pma_ppm_lock    : out    vl_logic;
        pma_reserved_out: out    vl_logic_vector(4 downto 0);
        pma_rs_lpbk_b   : out    vl_logic;
        pma_rx_qpi_pullup: out    vl_logic;
        pma_scan_mode_n : out    vl_logic;
        pma_scan_shift_n: out    vl_logic;
        pma_tx_bitslip  : out    vl_logic;
        pma_tx_bonding_rstb: out    vl_logic;
        pma_tx_pma_syncp: out    vl_logic;
        pma_tx_qpi_pulldn: out    vl_logic;
        pma_tx_qpi_pullup: out    vl_logic;
        pma_tx_txdetectrx: out    vl_logic;
        pmaif_bundling_out_down: out    vl_logic_vector(11 downto 0);
        pmaif_bundling_out_up: out    vl_logic_vector(11 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of asn_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of asn_enable : constant is 1;
    attribute mti_svvh_generic_type of block_sel : constant is 1;
    attribute mti_svvh_generic_type of bypass_early_eios : constant is 1;
    attribute mti_svvh_generic_type of bypass_pcie_switch : constant is 1;
    attribute mti_svvh_generic_type of bypass_pma_ltr : constant is 1;
    attribute mti_svvh_generic_type of bypass_pma_sw_done : constant is 1;
    attribute mti_svvh_generic_type of bypass_ppm_lock : constant is 1;
    attribute mti_svvh_generic_type of bypass_send_syncp_fbkp : constant is 1;
    attribute mti_svvh_generic_type of bypass_txdetectrx : constant is 1;
    attribute mti_svvh_generic_type of cdr_control : constant is 1;
    attribute mti_svvh_generic_type of cid_enable : constant is 1;
    attribute mti_svvh_generic_type of cp_cons_sel : constant is 1;
    attribute mti_svvh_generic_type of cp_dwn_mstr : constant is 1;
    attribute mti_svvh_generic_type of cp_up_mstr : constant is 1;
    attribute mti_svvh_generic_type of ctrl_plane_bonding : constant is 1;
    attribute mti_svvh_generic_type of data_mask_count : constant is 1;
    attribute mti_svvh_generic_type of data_mask_count_multi : constant is 1;
    attribute mti_svvh_generic_type of dft_observation_clock_selection : constant is 1;
    attribute mti_svvh_generic_type of early_eios_counter : constant is 1;
    attribute mti_svvh_generic_type of force_freqdet : constant is 1;
    attribute mti_svvh_generic_type of free_run_clk_enable : constant is 1;
    attribute mti_svvh_generic_type of ignore_sigdet_g23 : constant is 1;
    attribute mti_svvh_generic_type of pc_en_counter : constant is 1;
    attribute mti_svvh_generic_type of pc_rst_counter : constant is 1;
    attribute mti_svvh_generic_type of pcie_hip_mode : constant is 1;
    attribute mti_svvh_generic_type of ph_fifo_reg_mode : constant is 1;
    attribute mti_svvh_generic_type of phfifo_flush_wait : constant is 1;
    attribute mti_svvh_generic_type of pipe_if_g3pcs : constant is 1;
    attribute mti_svvh_generic_type of pma_done_counter : constant is 1;
    attribute mti_svvh_generic_type of pma_if_dft_en : constant is 1;
    attribute mti_svvh_generic_type of pma_if_dft_val : constant is 1;
    attribute mti_svvh_generic_type of ppm_cnt_rst : constant is 1;
    attribute mti_svvh_generic_type of ppm_deassert_early : constant is 1;
    attribute mti_svvh_generic_type of ppm_det_buckets : constant is 1;
    attribute mti_svvh_generic_type of ppm_gen1_2_cnt : constant is 1;
    attribute mti_svvh_generic_type of ppm_post_eidle_delay : constant is 1;
    attribute mti_svvh_generic_type of ppmsel : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of reconfig_settings : constant is 1;
    attribute mti_svvh_generic_type of rxvalid_mask : constant is 1;
    attribute mti_svvh_generic_type of sigdet_wait_counter : constant is 1;
    attribute mti_svvh_generic_type of sigdet_wait_counter_multi : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sim_mode : constant is 1;
    attribute mti_svvh_generic_type of spd_chg_rst_wait_cnt_en : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
    attribute mti_svvh_generic_type of testout_sel : constant is 1;
    attribute mti_svvh_generic_type of wait_clk_on_off_timer : constant is 1;
    attribute mti_svvh_generic_type of wait_pipe_synchronizing : constant is 1;
    attribute mti_svvh_generic_type of wait_send_syncp_fbkp : constant is 1;
end twentynm_hssi_common_pcs_pma_interface;
