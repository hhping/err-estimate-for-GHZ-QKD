`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/MuGG3o6NqUhn8+0Lxz4H5kqwTB8gLMb781B+FWYAQcW7YBeHWLBbnv9HVtvIxEu
JJbML1gktPpqd9/T05Ogvp59AuBjQqbX5ZLIRnqOllFsxnq1B/8GUE6OePZZfdvz
KV1Ae09xT3v3ZvCjFg+QwkYPXuvEBGgbGbccbqjq3YUPByYAATflH3BTyySRcfo+
ZaU7twCMiIIkc5jL8fgJYbAXLUDRGcVHaLEPFjriJqeRk1a0VFNIEJED9VSMbP2T
ERjZeu7Qxq74urd2Sh84nY5QfNmnLOnzZn9O2YjudewfYFxMs6U+JsAj/Oxm/8pu
GcJ7QOy2XzNSICbEtcTFKdtnNSyQWmu3jTVLAAy9NdjmSfdkk31i/usUAUhFTcAQ
6GGksaPEcaFOiqyjY97A7MQB4xC8iAvlobATg1SwnV2nW5ZGiCNjMBdq6uAx6Hf6
aNr8M6gZSHXGlSgwTgeN6ZHintWLa07E42RjknYuEr2az/NBFvPFLh+NSacBgDTl
qvFRj1UCQ3TS0hOFJ6Y7cp0sj9I4qaT2TfS+wpKJ7SHQuRbZ2eVq84R/1Juy7kqC
Dw9k6YDwAsST1fSL8P6o69eWSUIMjdPxW+bX1+tWgke/g/HfPT0+pYBL+IKdBnG7
L/itw0A3rBSx4KtqhbyoI0XB2SMENRudy8mwIIWz2pHjJqXD2GN+06C5V6YiGrnN
7LXz2SIUSJhm+9W65OHUKckPqlJOdXLl8niGfG875vGGK3xykumTw6ejO1VwQFym
A+sIjdS23Em0wDjFWONSZNtZkC+0PN7oELtpQRuI5CdC0f90oCKZwt9UmgjlFh6J
1uynLKU9tEAHaHKO8iKgwoc1VLyVj1bDvCdl/MlBcoBK7lVXIsAyejdWFiscNAkH
PtbCvhV0sauy2Iq/6a2DVJa0+yzmv2hFRTeqCoRPoqx6topNO4cDmCLsOug1yrBW
tJG2saDOKQ3gOT2KEsho/OHukzl6VmOUtL1VYCYDtv5yH8sBVN1oE5BZl9DNXTjU
hdBYJ8Jh2Q5VEUTECYqDIMA7IrH/dRXhsI7mqx5PWKyz1a3MYz+XVD5LBPanOzdS
nBfKs6BfFlHiz1hQtR3y4OPN3oy/NACeiqwAStpciia7P9L5CHEMa4C/ui8rl4Tj
GyfF7lRGvSju+J95E0k+PeRTyMe46v10czkEnnBq00Xqxf0MeITkSh+FTls0lg5n
jXAWZqHKE8of2Waf5/DYfcnwmKLPVRKsI9rVSyUV6rsfkMcVK/lb78/9vyb9gWKy
bKTSkKhvwPp+JKv94Ap+wTMzD5VQ/IC/ZzETHT+d+jdq4Pmyz69c1Toci8AnZN5q
p+2DjqSGWzsXmf4TOZnL8JjFBheAimHFOcaU/2yeHvtozpUDNVWuOyAptrA3Jd7s
cmfwdn8k9z5nNK1rFCShEGql2ODrdePRxQRewLtXVsbSs0tilVDdc9LiEr9h4Lzn
HylJ8X3JD25JLbzxQqbRxg==
`protect END_PROTECTED
