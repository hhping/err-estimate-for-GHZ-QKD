`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYpfvQ0ORBhOCIJQ/9JKN3tJg1iyb7BWb5UN5f3WvKA4/frZc/WL0kBlTvWBm52f
e4VsFW9k4J1heK6P3ukD+iBaKA8Cxpj3fi+UrZw6dcKSFxFkXNJjvEhtbADY+RgZ
K+QcvA8C/W1mLlb8Tfto73wwU+15ikg1iw86tOC9RFe18n5WUx5hHRcDWtPkk2ec
Oa/VKBegS5ZQ8ImfkD5swE4fT5YEfqqSXGhYLXXbxmjRa4fwX2F12BJsKrkfUHTx
nZFEQaTyg9e+tdDee4IE/UN3vIXqhOLcgqpEyIVXB9+kUQ6iIRJ5wc3KX9J7sbx2
ctvaRIo5LG4TUqrqy1ehUgrajy5DORJh8riHa2wt+SOE0FYTV2v8k7j+ACJG0+f1
1z0Mn7tikcUuTm8VYsvLfGVOsdfYH4oJ8ADNpjekGVLUVCK9Qv0wi+7rhseZ+gd+
CFXT5LAnuQEIgDZXxROxWrPKeZINcC65g1UlrotOYaIIfkQOu8Uq1wttE/3wPw6x
HDslY3NCBkQa+JY5LLpaxp67vbjsuisxWdOkNFuBpwbHFE9IEWwPwcGZDjGFsjww
rHBjLvW4I8YeiqF0nYmsxU60vJEUwmtA65Wt13DGhaMvyQbGIL9Oz5tfzOjQi5N7
enaoRxndT7Enn1qUP72LyMbEp3rY4Y1qjeLuGTmFl5E32oAZUEiVrT8FXRABAGJB
NQnE4F0nT/PMeqqYojLnbTwN05aLipYVZ3jw7zSGjUMgNRPYMylFAu44l/Kkqd7z
ZwFqYxvjgv6oRjNKlVDT9wHnb6B+e9Me9de/MeMS+Wo3oec8CVMIlkASWpI9s1Om
c9MDrPHXP2pFA6n5q7HA3Ny6W0VUJm/CXpMJ2KM3o+cwkM5/EmEmdahLFbUt3eoH
+dyEuIFpAAWtnFYOQFaPi91ms7CI8mEUrerU0XTNYZcZqJrFdXX59dUELSWrYpz9
zWDAArYf2IOXCQHf5cuzfAqbT/5D3WJ0/7X7EtWKCOj+Msw6qX8fBT39DaM8GGP9
NXJXkJvwhpmbx/6z3t7nAgtOazDpHWa6+DACkzLMsxW281VFrlYySt053u2MMBPZ
BfmVBcWwFaNIJwVQDjBPXIBlfAlMiA3RgnenzJIr/R8O6EcyWwKgD8/KZlMLUPhz
jCpdUPVoKDwz5rEEj6wDPKBsK14j3BosMZ5VqFH2JvoGXKwNlPFDawl8Fv7R3ilT
af7NVo3f32VHbtdBKbtkXdtJVbFvSXmWdnNnzCkUoEG8nsZNbWjtHeFo07/28sAk
Hv1gbXbUokpMqbqNtWLqb7lKiCBMU9Jvfa4nO9uFpdL0uxjoKpxd8kvohHh4j6zp
wh8u+RrhcYt+AK8DSx2Ne8mG5dyH8t76nudzzrvCA7M2mOVu+Y+3etAr9xwqz1qQ
qNqc1fx7sSdOm+ot8e2naS0IB+gUmMPLAYAchYMUOsjPWBrUSid+XyXlCq9A18WI
PPjFrBswaKMa5KYu3W4HuIkiuRv+xUUGk7fX4ysISgVG53+hxgyDkQYXIrzZSqpH
VxTR40a0SDqpHYGHTMPTrDNF6UzXkQY4oXWBqge2P5B4MQ4TJmdNDo+X69FxMBAu
nNmUEnI8xdWY1SxWdgTXs1DRJPqeQMIInpB4N48MppGdY5get6ZvKuoHY3phQ8Sq
s7zpeUbWhiGKH1/wtxUPUinmgdNAu0E9fjaCBWcnQLO6eneWVCbF5UlrL5HTo6je
nG8BSefXraG5QkztwpulPvG6tdlO9mcRrfAaQ3SpDEy6v333E0zUSt7tMsivzFJI
zM5jHAZ5PACdMxWXxyQ7HOZBQn1ycJixATR2y2rDIR8nJvTrN2MPgcOvHGAHshqj
jiokeoh5yrvx1wXRgdyRiOx+ZYcV/p31Vfh+uv9/z2EafFEDqpUpYFs2hinaF+rp
0xI0pMmD1iMUqyal9JieP/y6YaDzv5r1lGKEVdhsyMmlA/jSeBZ2cWicvfPwqYVA
Y5gEZMFd+nYsH/7JliXqo3CoEVog/ItFz3GzKyL3v8lh1yHQcvs5PWKb2OoBlDMl
4Ybo5JktoB7dBI08ULs+6aQqqt8N50IrOyV1O2YPUXr3WftldsvwdxOmpHoQiiAY
YdsNcY4alyxjXbY7EduqMTKjYBK3wjiRNWFTfTcuWIblIiIS4kOk34LFdJ+/azou
6ZjpjDVwmUG20uniLo2pp/0ICXutYbxXVC/1bT/nVH3TDMU8rwwujO6k32Yq/CcY
jNa9dRqmbkD7YJPhXXetbfZZGHkC/XnqfD4YovgSMbfgMxcmuqB0QO5giSupDynw
+X95xrosC5ylDZOnX18bCoBZ4BX4FmbJBsBn5QromZQWbFYmNsCSExTHsdHKwhK1
TEY4qGfZpbJbltSPKn478dSmTFMr/2MlS8IeDpGW0lXdIT44j/pjkQDHc9ZSyBnu
N/QFMKKRIxQ0ASnwrJ/t8UCzj0QvvHDdksia+n3ga5a3CaUIi4PTicJD8jKM/5lu
h0JeQnjIQuIi/PuMhJn+ghROAVMgaE8p73R0ZQWour3is7TSBp4rYDooRdnb9/lX
mfFmUYplbcRNHBcdc+4KJoDMcF4lEHFoKaW955DLbMzbBdYnkqDlUNPwh+LgX4EZ
z4c3MJFETC0IvctHoEUF95p7oo6oTdBar9FvUmiuIcqjhGz2q2j/5qTeOvkq18lP
4P7t0G9tQwT9mB1UWssSnd68AInQPUYdDcAqrA8cengcdGsdVz3eqEA3gcV91ScC
V03jBuhm2Xx0Y5vW2W30tchL+3nxkDdokvTiqVcjyLcaKQ5REn395c2ubRE0V1O0
sw2KVJabkMHrhM8YLS600KI12UKgzaZK91avIwkVMxWlldUgK70fRawRBql1qwWN
crpHRCIVNSRnyRfPXST9tZSQHM2z7uLvBhaaYt6AU4hXWKH3PjLOrjaxQqVvKfNV
/bze9md/tP+vsrxBjvsAOfA3Z7bUG2dlb1xTt14zlUh3znR28gtDZWPgQ89EIElQ
NI1UZS48YV02+6ppLOE2MWqaYHaQMUSQk8i06LqKv2uAQBYyxiOqrp+7Nx/U7l9y
ErtRHFktLocMoH+/6Zx7NIZmJCP9JSDozsIkJdc6fblVwqO4CXOG0gZ1cdrwY6xN
GJyqcQWu5vjeAxxvWC5eS9unTJ6TLELz8VNqSZ+Cb4aafq/uS4CNQsCMcnCsvmfy
a9kQ8BvlArT9ijI79SLkRAmd/GlITMiwQUoY5JcLOV3mj+izGi4Y1qPoEbQ8tqPu
GZPyfA0+/KVe4wM6R7YCfntZzfMBSRLb1smj0BK3vpqBLw8fV7VNBwIMoB1XL7r9
II7TXhFbTV7L9MlrnkNcOfTw9tFRuCpK5x+spjWi6ITw1AQQUWD82S0FBlwlrOFB
AkscpZ7BSFurMZ+3nt53y11VFYZ6o5bfBWzDidPqWjM+T65OW2jQvD7ttr6/u8Z2
bYkaBx8dGmbKaOZR7rd3e29MQ39D47f64FibYgiH9oiBpwsgfyhfQU8411AAACtR
n2VURd1XD9wUoIG6M2eqIgREFhUWQyrsWRBhXl+nixOTke5PTTgly+tVE7TU9xKC
QfuoUhATqzWsTJKownw3W8QLSbPf6D3SChk5snPB2CFPi+FTLmvlqA1RFr8R/Mm9
Aw6TM0vc1JIxuX65kIdK2ZUyl2yMUDF8RUmxn6C2E7FocDFQZ1kz7pXeXwQ1+kBa
Y+OYs3YrqGM56qRcHWkS3R9C21kHFKohZRTaiA6pcHOVIyza/Tulz9kNZO7NmzLK
xB4GlUcCu7oEq9kfbK899AZu9PAYJjBRgCIoVzMTleU9onCkIOL9yj/4hft+9fWe
/eL/qTNSXqmPnd8eYldIRG6tnn/v6dOxIWGLYrvQswlul2rOyo9JmGqYfFBpkAch
49QjINecGXnhlddA9A6+WDcCsJOPrnSApyX31RyNjhNtlYoM76WxOvRCbJYHArgS
kLVQZ8sisePak04CXsQEhzzNZSzbMj9r86AOPflFW5k98xOf4Ob4TEKA1MmOXb5T
5OG/+ltttEWlQswt2gaOMa7zi97Q3LksFcYPjnqEvQK2+zgLeCMmQR8xswGLAR7P
qzt/dMLWHfUif7l2R3f1Vejf6SJfVKNM3AUvvrQqUJ9Kpxej8+9pwensN3PSBzOT
2/q5zfJ77FxaN7VLJST9G6GFBmo7JXhBqLw5lXTGTNCFrIkNdreObjq3XZZfXD4l
8vYquDfpJfGwpsVsgvOG5rl1rYLuSn4HlAB2w15EA0Rng02W2rPS7XJdxaZLd97v
BGwrpDXm0kOSIy5YS/2qhDlwFySid7yrliPveT4h30H9NDSOvkWZ56SHm5BJx3+H
gaJQIdgZ/wAH01wGVgM9z2qjgMJ3KZwS/iRwNlXJ3J3vJ/jFWam2PvTVfyzx+4OE
/ZG0EDSQmfxH7A9+kusRh7nMX8aolzTyD9UCcw5NswYm+EMK6FMutKcyhJWAJbO6
sFf5SHCmXT2MaO7C4JUnO0ZlV9s9PIzMriNZKCmBDjhwO91+ghve/HuOE5V0vdtR
KQAZDdBSnAjrhNLem8amw322Zg4sRml3W3KHH9nQwPMiPQ+AVd/dRePp4WDJs84C
QFegBwupXM7lLs3uow0iIGnrtRWnC2/FyNGDYXKXqKplSbHjjL9zMwUi7Uqy6aUG
jOBg6rUTRMav35NGLvdjldhBPHzEGD/hishKVYtw/6ZU8GyVAmWMEhv6gFDO5YdD
TjlGbpTdJuOtakxNy8NrfpOyrtMwSducBZrAN22jIC5/Amrcf+1mGmAc0lxy9duF
NrquZOTBuwQTWOA8mB33Iws4c+MkervRIo/MJsKE6oZsEcjNKOK/+1zxnEERizFf
BBR8QPrZeQFGLFcWbihoA62pvNzfGD1FCM6einQmsU0UmjHj6o8bwJCqbPFCTQfT
cDH338U3mYCHhkqEGkecCDbnk2v5A7yQ4J/9zqLO//OzUFayN1+oe1HdPa43iKu4
DkvBdwRUh9ycRRGnEnAMg8UKxr0I47At+9OiLx36Ey+MDbzzAGHBGkSdvgx+nbcD
Nor7ZyXzqycERsmC5sgqZmEfIxi6B0awBumCqd3/sA1PC2syhh0ZVV6XSqjUPSj8
7FGe9RfGOXTxrFg8YCV5q0btqtGV5T+GqJXZLYcvnrIO8jjH6VA970Czm55mLkuQ
GESm6/RAFrO1SvuWAyn/9P+uesyAUD030VR+CSprEBHQ/OOoVYlQPUi/o0v8Djjc
+Jg9jBQLciIAd6dx2LVFhoiHh/PsBFy6/08DA5BpSnReQd5B851eyfQ13kbGj3Z3
P1W7xlk9TIFKQN8fOJd5aI5ArF6HKHqjv+XYewozc3EI2QOGuFO+7U6/KhOITbmY
qT+Vouxz0IYArqloKXLP4Ft1hhhXMrq29RlcI16UmPWyH9QSTRKkQNtOo5X2QGco
5zmAWOh9Jk8mQARrXFhYSMy//TqSGuIa4JZLOqxpbn56Vv7hjiv45pcTHMUR33zI
x8Y1HWVTB8jcSw2f9fOyanjDYo7OqUasYOUogNtNKAXhsoi2V2/WM4a8tCW/LOjF
ADZ4DX3Ftj1a+Y2RMFrlWlsQWahEm3f2jfjzJ2iLBH39kIuyMJgzeALLfXsUI3GN
h1oTPqWYRCg8UhqoPkO9iQhxvuIGv+HkCizHjGX2DgjjYqpn6kN3gfqiR0NJozkz
gHegomKMG7FjetcFMl7E5CugLZJB/9kdULkoEFq5mF99fZbWAg47S+pY5dbGvgzp
QYRZSWzRgRtcjgTeCG8z1H1drP/Fsc4VqTTTPvHzzVxLTvJ9CnmVx3/mRFxKaVms
jRtdFG8mSa9HKIuhmZfbgfegzDU9fXoj0m8HHMGpjIlJSBJ7TXX9JBvTtiFzou6C
K2fpbIfu0lSSejac98p7LHJv3x/zJOYUrMmFMPPOZ7EqQlvL7qpYFT5Z0F4+QsQZ
eXG+viGHQapVxsNwc/Uxb2b36zbYppy7xHSFmGZL06xWv7wxmmzophm6Nc/Atx8m
DsqrsrzuSV7y9SLNqtZ3zYKqhc9V0K+88i9VdFPIdrXd4wUZ8tNo40O2z2TfYqks
3k429QmVWVU+JkkA4ZzuLoXj0uLUmYap6Pe45M8d09LNk4HZfXij4shuNGv4PTlb
H6ZPY3ftqANI42ZZOZlhnqn+c/HWMxPDN0/wPVB4F7fBDRFn1e2d0C99LhABSMyq
PT0Ccng3kl946mFG71SEghULgzpFu1Ze2z5hPG/s4rGFrK0Er+E483RLQYj9XxSI
7YpGZwAVIIk4ftTKvZjGbJzINsEvtFjY+qs08CxOMpCopUR5PDPCsYUtUW90z5Df
yBLYypoVJvhGwpGh6pas//+Zpq4EZ/JN3wSSjvGY9wRIC+ZUsZ4a/YXySPuqu904
VAzlk2KBNC4p8DDbtJO7SC9wkJ2F9jAnwPLasr9YkTPOkMeWxnOrItrmDnX9agyv
DmtzjBrC83wejqySgga5oiZCoBUR0cZ7PjimqNCvaos5qx4ckAaofjZCj6o2P9yT
gJJy0Xex3qxLravPUfxW0g==
`protect END_PROTECTED
