`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCQBMWSx5sX9xVfey2qz6Tlcfyh8jTMwoN/0d8OHAmBqgr2AmrFLw8WjHVIhhFl9
NYcmOG0tgj/PYIotb1jKYFOECh7oqvsKJuT60zEfNYg9hHrOwLz2uIP5ppUZwShr
+nWp5la9bSoEmdkJA/GzP1aczjzpaLh4vgC4A5dSncLQHRPhjtFPTm7h8PAa1gGW
13EL9vuZjEQdxgN1qFAS8kUrekotyd1V9LJsRmCxGXOn0TF6wsgO2W1jtW/wkV2C
UwG6+EwBV+IcCU+NQIstqhA3ddrbzPaR4vlEcG9sUrDAQuQXAPsSAzqKg02yEG01
9j7Ks/7NKGJgMAIIzWAfpIJon6YJ4aA2HZbJkmp2Z9aZbkpuMZvI7MDDpU1tbPkR
7lCJy/0oYEDHyACx2PI77x19wEtIW+GrY/V47Tc+z6dtRGomImhdzzkeS78b+m/s
7WG+g+IBM2kcHKU4xdVAgFb57KvNe85ZBeBcVe2NYQryyTUnWwnYy8y/m1hdkQId
D6dEtikWW0mr3Z14729dC3PsCOEYXmIA8RxZ/VGZ2vn/W36C751rfOn0+jVOLNJv
aFHINPO9zIkR8Df8B01Vetlc1zWFTxUdNXPY996L/Ja/l139AYkn3EPRiEH1w4/F
LlzAxb/QZ4kETIK77kVVAw==
`protect END_PROTECTED
