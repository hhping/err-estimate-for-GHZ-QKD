`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYEjoP76bt/R5WdoiJdXggFrEj5vJmMgzRPqTBV/XaJsLV6SQY4Wzu+8FWKs4Z7B
1Vb+UoYmYUgpJfybfGUuAYBppvub1lsz136ankcjezaMdteOwhz3Fle2TMjaH1K3
l03cVCeO/eN6nqFiiaBBQ1cl0hLIjIYt/vBt/Gwq5+V/HDfqOQ+5t7BC0cydTqwS
t4iemyqJmTE2EPMoD6i+c9M5AOJ1nfNkdgS/VoujgHWPuY55mS2U8Kf/wCOBPWQC
WKAEmZwlrkNGNWbdGuD3p9Hy5BuOFgV7TN8O+uicN+YBtY7MJFdrDFfcUjuFtBWt
38pH7BP9K2Dg+un6kdDP5+fhIu0+mhTCRDOnYo5D7uMpbtNDDQYz7ji2p1ZISP0o
TOJ98jTABSa3c/5kZYMY8IH4Qp75meCJ8CPpOnuKcnS79yS+URaOfLWZZjYp5r3i
PFw1j2uT5CTFvdH+uH6wcaAstSHmLsAtz+jcAPmmVEAZzOt5ztxlwjMxu9bqHcQE
nwtJyfzSy8ELeVCqZkElNamQznSkXw5RtOd7jTdLCHARIXLmyAk4UU1ZZ5HS5nhv
WbhSDSBFjnUvFRte5pI9pIPODq8cKibklSy9/57jRefujJPLm3ZeR3Iv3jULeGjL
zEb0OtiVrwefOQO721S5CHozf5Ss2OOERaLAUEoPlVCaEWAWvLElbMx6ZZEb7bvC
+YPa85zIo1xRP4N3Lpul/7Oh8NMt3Au1uaI2XdgrwYdU51B6dqrqTjqwDshmOdJW
EnKXYa3MdUZlfEvaHkULJbNOBuMvqVJVm5H8B6gH7WVWS91lf73/onhN+e3KcEQO
Vw1eRm1CF4M1sus/dcNoEqHvJ67APhP7p5S+wSex9WwoXzEI8wPGbZkfeqnfyNDc
M971sRfZHFWN1ZMrrKuWngVI8NescCpPUSulht5y78Crq7EShW/2tE7xfMaMzAYC
zjN6zmy3YhOOApjyUuwekBUrTHnqY1u6zpgdWIVqFrH5XntXjWo7roe/NNPwnzds
0GPqEH0P+ovEgy5jZKh6uDm9ZkzXU9fOJ7hZvWspP3jo/LEoqtKA3SJ4ly5WtZJK
P2vkU134QkM86z6vAdZi0dWFiksmkznoL5ec9xYDRxOAPahKrgTGq2LVscZBIyAn
H2fLQTejhURpxjS51GtY388x8i2TYSu45cacg3HeFY3yNM3vLMozXnr0tbrVSDrU
rEZ915hcSEUTPE79jZp1zlLqN+9VAHFuhAnkWrkUo94WiT4nNwUscd/AFLxCfOiE
ZrW5H4SlO7t/yoPXpf5vwjrdRG8B7V0MnI/PXpf/n3K9QbhFKeBdLHQWTz2wHY3E
kjJm2J6By/CFoKltrU6uXonRXrCv7JFRH0WR7nbWe3LX7jJ29gj5AdA5HYvF0HFl
xRHRE16jKi+SBVwiG5IzazCG3IYvPlLlx8lLbe4xIcJHO040l9luw+ObZDRKczzX
cLSvsi86bAOuD0+ac2ezMp35VrW2tHR6AtNbO4fz5c3OsZbQ60aXhvUIPIw1mox0
w6SF3aRtuFTcgt/e3ymOb/i0/dl1oqbccmrMLDhinSWAJ3JdvF9TL8cHyt29j0qQ
c4GcR5qEIGbT2+ScDmqlrLaKWZ6HPpOjeCXyIQMQtq0cY16MfpSfNMQscXRrBo6J
FaCcu1B0b3t1ICjsCJyxky6pXPeGtNumly5bLyAvNnvfEc1llTkDuKE1o/Haj+7I
p8T14kMdroFxqsJe3MPPmE2696Q1j0yZOp/SfsKRq8Y=
`protect END_PROTECTED
