`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6p2l/756Gf6xgsfwT3XzUu5ELudagZSB9I4ucS9jre/p2Mt6zLaYOoWE3QVZu7Eb
42rmPGXFItIH5cBl/msqvLBTU4O64Hr6CFTna1BwXEBgywayqSt5aUq/8ELrYOeV
Cy5NwtdXoq7dRt1pPtsNMgNw+vcj/2mjzXyo1W8eM/CltHZKKVO1nkdZzgVEEynf
2jlJPadJyhx5y/M+tdr2tcjPr/wl4RByKgCvhKopB+virTzhY/ve0+AwUAeeRUFu
K7ipbyJ+VYULNME0Khy5J/5UHkKhelz5lr0X70mIIWAqDJUEO8N5ZwNR1RuYICDI
3KYbRt+GyyzLatyvyChJlGAohgLg7NQBAqXq9nWyDn+NBbyl9lPvs/q1q6Mk8/Ob
kN7biSz8FHu5/X8W0XR5KiC+OpwSR3beZGJzbZG/x7fhIvoopbUHc4rAgRPdvzgl
/EA9T9IUfVg8YJFnBrG9HNw2oKlTejQWezAxpzqErEbEAYFFg9Y9yCIsnPEQnHw3
nuTy+ksTwK4oFSuZKIPZppx8D+XvWjeJKoj87uQFtlXpjkDPjjCn9sqKYfKRF62V
CoTsoPHyAp7CDoHzYUZkw2kLvYSUMTWYYqZ1Q57YrPp3MplNFUmeETrM71OzWjWQ
PaEQOSwO2bh5lPCQmFSRinoXmTNJScQpN5mylAfzaYV7SlZdHF1c+oCdQw/4lfk+
MIoq5lMZhqj8aNisJP12Lf6DNOVLchzasNgPWQwj0GWegrST8I7TSRMoJKlfWvyJ
9jefVyl+NbbsfRI3Y7fjclU9R47eanvjdKL/hyRaaNw=
`protect END_PROTECTED
