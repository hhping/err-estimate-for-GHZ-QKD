`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
po2kPLPUCG6RE0d2suXRLjL+ukvCrPqLhgnIMFh1Q44Jji+KEjw8uho/t2zGJZcI
l7zgF9DTnsWio+x6hAcD3B9fWxm5eNUFElPUBSFqa4rRDaaMM87uzAk4LZaWlWDW
4IJliXiPavWK+0eayHk2Hra5qKf9rqwy9KNBcBo6aHW7DczGyWN2J5WjWeLMMhtC
gUJjK2Ch0flvE9diL26RFbAffIEU/RTaOjAfV6MUg+OhePx21Ux1RT+QJ0b+4b/t
FqkLwAOh/TfslqzAtBdOl/dP559zd0u2SdTrNmxnK7TK9oB5Fzy4jQ34QAxXs6UB
JVY0LSxb5hNBGMQZ9Rdy6joUYC7RbsL9dinz9Iqns7hkDlSO+Q057WLxfqbBMqTP
nDZHIdRtxF0Tbwnbkr5UwfjcJLqQ//ktp4f2nRzLX2iJjbHgwm13MzgMrggX86lF
PZfFB1BN0YDBcAvXtPKhXcAjU9eBS9Tu2Zs/L19iWKVFpUiPOXv8gKBgMps9LRZm
pKFhYEbBm4hjZdU1QtR7MCY0UfXvWL7CQt0h2VTxRQLlMWpBDNIYD3/1nWgRbNQt
zGw/wvFMoq0cCb8ouAMBn+ScGOckZHtk36BSc329sUTppYSvNmaBQ+egRO00sZkx
uly63Ll07XiRPl6upDjRxAeLnbJzBIh4JvJQpnVWsiL1svk5sMeHk/lqne8IjW5i
WCR/Td6W35Tv4nqSMN9JON2RFmxO8V7uKxZB1+K9XhjCuyAM0t4KeAh4Ds57g81u
9AsWH6q0r3qCyPDwPu+gx4pLoVsiVasKHqkIPj3udYfnXvldSPZwCwI4Ibbbl/ZQ
BAThRhc+6xTWZskvHq/aQXLUA6UnYw2Hkc/jrZRBgqjZawhmJPl+VxwNwcp2+Q+H
Se0iKwtjj2oIMLVyPuPHfjQTWo20pfXkdMK2dfYjOjrX2o6sGCPf40kU27SADQKs
cZhsRoq6jUKHp4GsRePRY64h5jmSoNs7fyta5n+ZXfal+dApZlwmTOKJUSpySChi
XN4vqgI35otg0fs43fKtveDE1o+5+Pg2adiKZWaDk7eQq1CpFmgjmKI58I4mF1rF
W8fICmZ1gfn4P62Bj8y+cYsYb+nEPesRVTLYHDD2aOorRQQjyoRgPILJDgCwl+Sk
AUoom+u8IDlyxrhvbHrAeWDP6SUN4yMDBJNNDYSvgyLI+eCp98CFGo+OitQK5D0o
rs//WNCLc17v0xJKa7JBoW3pWSCtEOAqFEKo5fBFoMvoS0BgDf1mpHWJ/oemS79m
2ruOwG6QqZjo1xEjJ6iD8bTFvGd23as+K7Pk6y1JPV3gZP12FCd0f+hdft72PvmJ
s777EFHQXM9Nx1zwrBkAj29d1qsP9Yw0U+YvKPBfSG2CWbi8SnYWsxZatZUa4CcS
WX3X4GDmEKYFG9l6cBMMyGFDZL4yQIK4G17KBIAGN+rrMFe7XbaTZ2iA1ltZDYbr
ouFBM5PCW33HvPifKf7EYOAWR88/FQFAbioFzVcrUKDjqrdrdsc5KKXMS85Z2xzl
/GoUb1cKoMbE0Wc5x5for739BA86qmpoVmYoReHjzT9s/+AbJnWOTjx8DSJw8Y4I
NE18k3o/TJqeYCZ3SeIPc+MwXCxIS0CBz4JJaRHzjcjmRjCtv1YNFr0i6x/dacmk
a4oVVnSq/UJgeYuhw2HyPxF//877hApduK1uRktkeZ9BtNup+Ke/cDID6LnpN0W7
OCQQZ7Iru/+BmAoDaMAtnL3VmzcfB73DXcXlR54yxTMEdAEz8GSru4g9B6XeO207
D2/jBifiTVMsLWrgIg8Py93xjS+vEsTlJRUhP/CjhNy3NML0TgzzAgyE+7Ng3YIy
BNLHkCGXf1pDRt3cV80kmxuRAg/dyfn7/yGpFiOjf5eoWdP5B/SLtojQ+PoVMDPk
GYVSVkC33Z3scEHl9NpWd3oBt7YxiT6fSXDl2SMcbQ3olzIqcpc1E7ONADuX9AD4
SayU49KS7VR/A66P/m9a3loXzXQswziovAvRqRhsX2yPwAo9rtNBhTWTaDMuY/1f
mVy4dLYL6zpsx/kS2ipx/1h0PJ5Pyxj91NwvxWoAVgLXX0J8UtXwEp7txZXYiTbq
/xyDATiMAkDkpCJddiveudqjPnXfTJ1clHhmwkm4YFMmHPHMmWMQNbB+4tCnZ/LW
RqTBbDcKIB6UiKU/P3VOSUiXCQz1fuwtALH8y8HZ8RvDiT8fwCy20kItNZ69z9nl
xiZdlqeDTPvYxBawF6jxxKtATiSpf7Hi1mzi+6jnGtZvuWvSepCfW1W/bFPnmliN
GeGCaJAV7PxticCLyO66NGwucfL6k5kr5GO8VRS4NVyTUqQ+zeeLpwC1JjSYi6yY
F4SIfBoIJ/2tV4rPZ2agjwIST2KshedCcan2NfeWZxVKSahRi3SpPK5ji6MlkVV9
PrfhYFNxBzwoe6ynpRfQ9CieKNhQ5C6aOQS5O6L6TSohjBHIOHX2eLrcHXxq7gG6
G/EXAFrmY1v8VMhCWssQnw==
`protect END_PROTECTED
