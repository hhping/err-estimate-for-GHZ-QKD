`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5UoKeNlNU48jknZl8Zv5ivtmzkT80Ic5XZqP7og2zmwz/siXQ3OC2A6NgkPgNcyz
0hha5yTo2e7npdlTJsbLzeuZ3xGce/otk7jaEJt00CEUjNmbddiTH3PK+LlU9iIl
PgdpnUUSAa7KqF2IvavvuT/rVTDrvtqk46EmlRXqmRtJKIwmXdHSCQJmAKxzJK4W
Vkqfd6QAKT/wdtHlnNBc3ZnuAiEdZz+0OafmcappYGl+qmLs62iE/CGTKi/+q6vq
v+1OSxcPNCWu63kd8g0IEG3N6R7tWdMth+1A0bFADl8j9lIv8uFhSF6avSCkjKOE
8hDX8DlmGasoPjONyGHX4jmBWz8/aDreWNKemRo8qjtUoICglSjHe2vNXWxdEfhS
tmE7m+i8bOop860xllBOQQ==
`protect END_PROTECTED
