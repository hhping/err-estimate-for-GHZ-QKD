`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30jjfSqampnfRCtj1puW+/2iysrvlvrcTDY576P02qn1tiSwwA85xbjy2gLQQmbt
gz+d3P5TKVguQmDAcv19z0vNPiVrbgAkgH7Dj1Bi9CCaoI+Z6zjVIcktWKK3yBkx
bMFChcDsHd/kQ9RWiNgeshCICaFot9eCpGZMny8Mhnl9PTbncJMKXm72HfwyHwaV
EbDPM4c66CLeyvKd+iRJvZWhGytT4mYjIKoQfrNIEiXLRn7ddcwaYTvvP0kSOTP6
ao/OShil4Gw+XVamI8Ro1BheLXRR9N/saKneXXQWGACj4/GmNvDH5OgwFphkkROF
OguIUdV6z3+Yrm4aalPp7dzIBQ01YSe4+6L6Fx5MkTh7HJ6wxOXOq0akTR/q5f8o
MUckadATClHnEo2g0Bp/SY+EF7ttGpUIID103ikrvvpEAkCoVqXMRj6+UOfWTKxD
rKbyWynYNrb8XA74ri6V8QHeVnsii8O2FB+RnZTQ7bMNWZdwfmSZM08V+lKAw58/
PJYRRlZ+EpweE+yGYj7xdrNn6V545W6Gzx59i5/rkaxwXcgoDc1vvGJPBZRarwCG
1XzjScZvm3z5I+eJ6kM2uw4U4sxv9thQR5dn0o37XoeA0TT/awaqZjOVAQ2kS3Ke
z7MwMNXIP6QvnyLl15UdeuaL6KPn7wZ5hgoGLeTlAk2cMuYCMLlDMoBaaFiXLxcZ
Jkwej44EEoenBjAvJOZhoEF/6tKSbShWppnZEsRFTw3sg5CWX+q0mwouT+6cqo2Z
yD3VXs1rw/XEKafIfDPNGJG/LdXUNZ7eDjok0VRze6/BpH8DOD/d62oVL+slD+dk
bx5f/iGz36nHiqqbxwrvMI3wuywbTcjtCZaIVbILk0ANBarif6NYBfjNA/4cNmPw
HQjP2sIMsTvVQBFNlMMV1KKvXhehsUSkyl/7iaenmNdhpPPx+vWjeaHwAMXnQrPz
Y/oczNxNsUU2ZvZRlzTgHd8Y720rwZ1d2WkACxMjFouSFNXZgC26uxFO+5rg50ki
hU3sIeoxYD+f/C65JRK5rRNJoy55SecpDn43w+a89iIfkOTg3aMDC40CIGBBnpqy
GFkuvV33adOSvkAwgWZk2ZBwpWAwm1Qtv7lhZX/IdkSwA64p3CPrc9dbeFHTO778
j7MWb6lOTTSp57dSjJmFKo4ENRblE/CsS/oatA0FaWIaB360spwNIiD9UeYzZIPo
Aj1gkqSCC6lbAZHLAVPO8wkwA3VuxC9VDknLFy2a/5DrucCBkRIpdX6Nr+De01Xx
qgvCnHHSLhwy7ThGgZYl8muvCDWkjwS4woVSIuttYq7bA/o3s7aV060fwHoiRimu
NQuz0x2r+ROlv5X00J2yg0TsmlO/XiUrJ8M98Dw2uoYjuD2vfARwTN65vLfiXOeI
Ae+34yD1LBsBhFbNjFiW+A5sYDtGAvwlvx2f2UPOZZcc0a/0ot1kdPq2z4Xm3Bws
lIrT4VHNaQhxNgMdjw2HOn6zNNRF6lknfEXIw4rn4ACCDRu3qirJA9juGQ3YPUcp
Ijt9KJ85WGNMmUkrAQ4CfzYTYP2lXBEyKHVOrzxpbk02e2sWNZmZLwhhCRscVWxd
+Msgr2eFFHdTon3g3f/icqKVybTakH5S9IwmS+FoflwcTxkz7UK8SIz9/6kA/Zg1
XYoyFNx2z/2Ly31SqKiiOk1UZmCnN0ws76QT+PCnZUTsISvafwI5il9EZlPO4Fhu
6RiNU4Rt+TlKXUrdF/wWAesCcyRVDbo5/aqO2s5WNp1HcQ+4/FwLy2nx/+CSHBxC
4tCkBn7JR8Y3w+wBd0NtQRst0NWRkkY8Vq82o4gmBk/KK+wV/dMc5yInmWr4G4A9
AKObwgXautm+M7ucYt3mGvGdBADx/PBHq5/KHRSG5q/8s6/ZDLKTvnfVOwbtBHHT
Kxi+p1HdyBfiX7rWKAW3pCUTZrkCbG8xc7XYtVOuiMTeaLXYvTaiF9tTtsVB0jXl
iORLzDJzOWsPagG/MCD01a8tGnjRRi9dmdoeCPCQN91yXFk3Dr4/VcMa90NgvFtj
GIRkSlWxvQ0w7EN1yQtwkMbxpr/AXofdUDxffGKbA97+hrCVZpPAvAHiE6whDTcu
dtqyyAv33W9FkVx40mfxAaU0J6WyTBCp49ihteMARy0+ADkfjGVXWjgC9YIf4mYI
nAAzsk68V1yl9kC5Kh25aLnOWzs26SdjFtHlN/Co9FmZbKuknxUJJhLHl13S5zNP
XDUXQqY4OHUb0vTaLEwPDXVeGDL2vZOQBGw2TGSL6M7xhbAREFfZMPSmWUSDs3cM
jxkhjUOrAqmU7nQZ+6Wc71aval2FqCPaieATsUz9gtIsGIGZvl0rkeZlqfusPl3o
7fwoqIa2JJfRsTxMoTthBzsJ/aKdp+8inYYE71XNLSO5WYTh16MFnhoE0reFf53E
yyB4prl1PesJ6DWvuBX3XKy3w4Wpi6dg9S9cymoNAmCTTvE8yAghIADxmLSk7fNU
p4dOTP97zXa1KtW7ZvCcoQt7eEiqMBCOcJf6aZ8hXYRsMSOwAq3aOWVLil7TYl2g
2Msjr+nTvbZiZdR3ny5bqVGFr/3/syweFKS5mBs+eFhJnvuZV8PPfm25bu4tQCat
gsHhVMnlIL0DR0ax2zuLjK12gba8j+lbKL/bsvK98E/oeDwJ5aHMMPNOfy4sBmTI
LhjYnLBWLHsYI3fKU9DxZh8NuUxgjKmOtwbO4BTYzJYBdW9eQYbHwBi+de4FTDc2
1KjdjNejHRj5/C3d9yXgdJS/2ju+FBBZnzWcEyBFjEkFRJpb3HxpBjYq33nGnc+R
TAT0/km1ddYa1Em1Tcks3Ae71EEePIzTwQRrmceV29Fh9eB/4YK20LRCHUNI4aVP
n5w81LjkZkqAQTnc5n43UaOSd60ObQ5gqnSxjHhwdol/6XqHN643MDiv7nCe/j8P
Y9gnZ2+iGUVXNUd1j5UFEZaZh8x9v9ymnVsH22FdTeXR9WiBYzIWIGx0LaZoYqIk
eYdrhPVa/Vkhz6yRR5r0y5w1k4rgiReGCGPYKHHMLAiW67kVFJ3DC3nKjaZmN/hY
G0XUezqodF5D3uLOsl/YVo3OW+MnkJZZBjSwF4ghJlzqi94oaToSHfzZJ1INW8O8
z8IDnh3qlfwp/huABdD6rqWY3xKUD1RSEQhQ+/Cd4AvCtyDu2NpXdcIYdUyHgJ/9
xwZiO+Nb/ro05O6sQK7zc5Jw2CkrggTZoIhVZVFK5yuOxWiYZ3MX8ytH6uosoijP
XThJrVj4gn5+dUplsF01Q4m2m2LjOms/PitvUezDEaj+LOz55cJi3u0kdrkIcH0r
L+78Mlv0jJsmTp5Rpjy5X9wJmSbHgPGl2+qXitEYscHj5Z6+3FvLgmE7yywF1cIx
W6ktkC1gafPSsLvY3xxj3qFmzDsi6IcTjTSerYJf8RUw6273sEtD1Br/BKZWVgrw
QxOlKmHr1eacWQ9R2Tuv+WuKAlns8Z2rtqDJGHFmbaEsIDPP0c94gYoYqUg5jhdj
hdXxmjNTGCi+R8iQg8aeXRaUHoRvmb4CZwjNoL16g80JHsMp0b9EwW/6hFrc/jc3
jHeOIxMWXskr9n3wWXhv+n1HOqqtTNyARm0ktqZaXrTRpP9xCitLXEbUxxMZZ0Sx
OFkPQsUAGKSFjmsKnsaxNfLA3TYhSu8Atd7h7jNHlbBI/RVyb8Zlu10kBHiIpZ3r
pTkZVdXnp3xvzWzaQLFAm6lJnA5fL46owupOh5/vqqSeAZjHesNLtanQREcxu7et
o2mmv58AsVUdAT85o4+k81Kcdn/kShbZ1l/Tzv0tZlsyFNdHoVZ0D6e/iri39xqd
nye+oSPGumYxkQqAQErm0m81iwNiMUxJ7VWnbsADSjHbTIySlbSa/MTiBJ5E0T/f
pfWAKETUgdP2PM2GE8JR06ePS8xNI++h9lsLG0fy+LSE6Ppv0A46+p6u/MwgHVd1
gWOdkha8aQT5NMl9iZEWbx4bn3tfTyf0mEptPioit4x4WQSD4r4cYLwLWyBBf+Sr
owU+FokKsoXQaxvZk8jz1XV6pAaKpr4A4mcQ+/OjH8Xcsek0Bo3JAhvL/TUotM0c
vVb+Nhb1eD3gOwS+/X/8Hqhc7MLec1qwBhTrnAJDrR96f+/0k8L0N5jMmIrr8XMb
THRefMqsI5yXE44s7F2C4bkQ4/YFeP8BIRtgxYHs+dpiiV7aYe09RDB9LFzcVT5o
lruBnxU3N54/8yJtCcZhK3TIrN1vqBlcdS1sDlDUXs2UcSnXqwfGjK/2OIffHCUg
9vJPmC04RK7OVPFPxeZ2I8831VfePnJVTYSa57+Kq29SIMEJpH1Pbv6lp+AhdHiQ
oRgvABVs4DqCh4kNHVkDd9+coJ8ga3K+PHwAM1AEMYHG4P1dgvv485kxkCT8+om5
oBB0MW5esJuTeZbkFLnm0/AXkV731iDuHM7HwQG7ut8TAd/qVbBikWxr6o9zE5gM
KvoM9IyvW84As0PQAPGMZvonLhwTdQO25QllGx8OsIPsoWPWug6XtreLoCuifDmS
NqVJjViSa0+6RVjGh/+wQ9Ozal9+E7lKzLGXBdBAVR4uzlGj04C1DChfbweSqQxV
iONGhJ2uIR6sgaLiSXyU4cEd+1GIeuJCYuypmrRrD9F9FzCTJz30kKExGN1M8YS8
sdT1wxDZX18A90uUenQAfhcsRRTs00Hk766TDmo4lK59a+mYlD7qwHGueMFwzOw4
SoJmjlgNnDqpRdcPFS/FuodbHJGdpV0scIY3M9nP6/alSuv8gKgWCKOjYvGSWb2s
SWr+ckFTwLXYzFaLiBiiC5ViKAv/3Qi8tj2apTOOsdGwT05TfXOF023xLw3ScfTm
hUq2mK+jdOHOxIbxvICx0Zw6AaeOe8pLJ/zMsJLtvXRdlgcOhNAOgt0bSs80IDtt
6k71EUkS9lI7zHa+o9roxfQ20Kowfw0sN0cJFIyYGTRrHHKsDVDK2iphHLusOMZ5
5J+dvkAJ+mO69ZJa8kSsOP1UYb93P0hr4NducbY/AXS2wC1Cw5l5VMctAX4p6kYJ
NKgVUYxYUxJskxKqhs+IB1lHLzrjB/j10Uyj1yxDcBpaIOrj3MrnN6FZ3EvHqYB6
3EYjJmB8smp3JfVnyfZ7FZ6uCp4XNkvorG4JU7d/1MBhI1yClBQ6AmiJlzcgl2j/
irNM8SeUh/koUBlJYG9sEzvo1mF+Nfz+TEWWxvgXyFfju6oEVnV8gT6UcZWaFpa2
JAp+xPO9x/Zx6Li6ibNokUz0A1IUj5gBLTwpfvuYYkiuaibd2WCuU9+NiZFHMLmX
ein5SVh0OZ4Z0r3QtEgwvvu5Kkh8OpUcdU9bJtQvCyfmAsMTdZdrVOrvHzqqqD9S
na9rTzow75PcQlmqEtMwz6mJDFmiJ+lPu+kiQIwuRhWEG0pRJImDiFilWqmvw2Hn
U5vogkv1AExLOVL2f+nLhJBy/lAjx+s2aWSf1UvDRI5rP2iNKd/5JBD3HahEtTCD
k+puGZavRktyyDN19zslWYBoiJUlWeWbH6CdIXTM1ZzmqXcnh/eY/BE80uSSWB+2
oCOoAhvePRkMeGpS8ObHiQ==
`protect END_PROTECTED
