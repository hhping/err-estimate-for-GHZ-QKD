`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uiE3XNWWU9sReWKATyfaEPKVN0a/6RTSrp0NsdSmdV/YLaxGa6eeyAeMkfDa6Nm3
KGs4m4mQwFavqhwvMeOIUU8xdphwINYEQlLhNMindNCb3IDwr90N0qpThqYYfaHH
ytAPNa5iFfDsIH1uxoJ2iQdDOprMK2+0ZHf06UpDwQO9Lg9PHQU8xichsqmr3EC0
8neG6CXjoblDMy9GbzvQ2naLmBIGnXGz8n7vG0N45FUmr2N3n2qNTs7tOEJkr8Y3
5hpMKnIPm7eb/Lmfk35qTkPgT14fvfe9bhqLWrT1gYkRxG8B6OmCwEr0xoq+83+Z
/bCjhlQ3SqRszFPDWeaClFoNThBuzNJ/l7nNFrGgN1v5m0iI+6WUYKII+yVkYMZt
gnF/ndjuzH2cS9rcJ8QEYD2rFh2jbfOpcZ0hIpJO6AZV9gvDq4ssT1jh6bbj2XV8
7ggSkTHUNDKm+WLHXG5g4e/RHgcRHGHPOXjFAxUbNkEodUQEFMl3jcXpZVfmnCeq
qvQZ9OUDYe3of4xo7+I0vApGWOLCwOzLreqpK+NEzGu6fKjEddjBsvNl4yZQ3VHh
SuM9niRk4+OpVbKh0Rn7JIpzVdBJlg+Y6vU2WlYd/YqWJHadnjP1ItR081XwlaOY
hqGOjDYy8YiAxrL4Der0JhPPptZDTlIs9KiOta1yH/BJW8ASOCVAFyJQZlM/Jk38
`protect END_PROTECTED
