`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z23wJF9CTDIg7YRqRGfxcLAD5ReNUaAJEkoAUa18EPQp8spSyc/RmoPJiPj+pN7N
yG/ZUO/5SqPbJEz+VIcrP7Oy6aN3SGPYw1yiUyNOt2adJIExE6vvMlDvp3Rs1q4B
oWATMKgiRvnvIrQ+XxDqbBYNv/SGVUHo2TWuBD1rX/XS+juJ0YjRwcTZ0w+4NKsg
N/rQayoRA0ckFSr31KmJMVB/es1zR5y6kz/b21LqJszFY24uIgzPVuR1KOA87c/k
E0m1Z8biBDaaaXzuY1Kp4m/n3pHQkI+bPNT/L1y5eg97Me7XVt+FL0BF5i/S1TlG
KJpEw9W6zeUVSyIAaT3QlRxqTStiMldTK+bdN4NcYGfZUdou1jA7IqqZa9ITj6lE
`protect END_PROTECTED
