`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0Gv0R4l0OkuTpLA/4/HOmUVXu0SUEYCa0xqLwRYTW48LBzqfDg1cy0D0F6wqSZ6
yL5F7awaKFGnm1GpWaULuZjG4rKVhvldEQMUGzYoChLPgOwFz2iR8xp1uEa1uSdk
UwF94frVc+P23TCTR7Y8es8HYbRLr/BxSh3HCpXZZPb0beIBYCUS7vUc4BuAYEIZ
uxcTz1MxfaTMgZ6/ysDkN2o8XP1hKS+FGGBKros6rGXesiT7sjgDZT/JUm+hwkvC
TErlcfuYM+ggj13+7yUsGTpO7kyZ+WwMIAdRY0MzjguT+NNagtcKEuQ+U/XNkjS4
bboPQFuNsDW5Z49O3+I2cf5l9YDOX8rZ5uFO9Wa07RRF8YJRnok3Y6dctOLfa2/r
ZY9WF7YZBCUvge9Qgs6IeuVcbEVBVf9ubCkwmFsN+S9lAjyfc/CtV9YDlQMAzgoR
6lWp0CCnroiDeG1vJH+u6PX+mzkvI8lkvgNOtlWnGcR8VJV0VBlsWc6fWshu3iT3
OvE+ZwosIT/m13VJ0B0IjKIFT3mgNUxKl5WlKfs0ZOm/B62G8iYTGKyQnHQDENyD
aUFikC2WNtOn6lBxk0UAVi18jMX3RD6G+6Ra/1ip/svo+zaTBa3g7UtH3v6XauUF
eePLquJ9USx1+bCTQ9RiEe2PFLpWnrWnTvDUP5Uesvl/6N0BqcPIkXDwWoHTPYwA
5qYCk45VuCVt2GY0Z8rqSXgA9BpHTu2Iwg9nQDI/ij6KicCq48USFueXs6mMxrVL
aqkLGRQhF/MAAQEnLuKkDV5CgV/67P9aW/RoNYt7K2lKhVTvgWMD2sQPgZLYa+Tu
ryN2LggEFXFdXKxUl8yN1jWdk/GlYT10W8H4BwmHyg8SXBK6eonlM6pS92rNbpMy
0yaoGM0qyGwnREDyBlefyvPfPf9SYnDtEYqQuBkhN1TpRvYzOYFgHe694TRBd/ma
tEs/x9PkMxONpfcYDO2Xa0VVsWITLzx4GvVbTcN94+3Yhj0Oktv3PJ/KfWeCm/9L
SZkJEeuOnswqHM6WM/T0mKf4KneGVvweAmDlD3772aTabblHlSNlZFcp9EbVqbGE
qNX6c6Esd/qgrKVq1kRat7eAkXY4IvyL3EQfMDuJm4vgYzQoKJ0y+IVMKOsUDzSw
9oyoR6Tc2EdMTvJdHErr7BO8327yNNddSyTGYkk+w1e2tIvfGxNclQ/KXxgk/Bes
4Ubpws9D0uSBgbr8Yz8oD4WzUgaI/qI8a7z5aX9d4iyhR5Ztphvgh/DRxA8H76JF
wiBRN4tesMA+++TZDYBb6qFEL3Tprl/NN3/j51YZLcZVE6kx/YltFBCNlKImDX+s
UHw3Y/hi0GCidIWurMeEWutbdOFtwKNoYEgfSCSFwtVuTlpqk7WfPcL8OPzzGMJo
GbvTspNFgSoPvf3Si1Nycrp010C6dC7YYP+FX9vbiJtLEGiB6GMGwURszSnX65Kt
VFbbhrth2GFkqlwme6adcP/nNgQtDQEHPRDwCtVnKEPACMXg7cPfrDfPzj39INod
eWHbocr2vQsGVHpv177gip7nD6snJHQXuzhZ/UfebdYjANNHXRMcwETBsfgKOlaK
bX1/gLzhEC4wCE+OPLOpOdqLIYmj1k2TbGvSEAozavQVgs6sDsc6lBn1OcEmdeRu
RMcJYoSTP/xcF3Ck/KfZjFa7NxoDugHR3wnqHbWZ8JA8vDAnxNxcOGqqnfUeTSMw
l8vH2HneOWshq2tHL7f7nWImuAurvL6pPdf5iQ6Skn/ZEb9vAAxHjKQufc0Av24x
jshfXdLZdq3XneWrQ2tcocB4yoT/STEF8KxnuUIk/hPtaHBvKeQLZNwCtDdgf7NO
VkjQYVOg+Q2Yo/Ko1BYCJ6ysrgF/MG1ZTjRiBgJE5N+ZN1t0/g5Z5kA+nG2xwKQ3
j2K+eW9IWp0l2dzEoq6E4elRy8qW7oa8WoOmHExFfR5Ze8zZz4PNLBZ4jKqsdhI/
eRjAXMmpry98KWWRibh7Gvq03qL5gLVBCKc2KUiEwgxVjTI+b5e0aTZ2jYgFzEGZ
9Mlsg2eFeMf76bjs5U65SAuVaozqbKXuBnC+6paWq5/PKQ03Y3uCydCRWG//Ijcu
xRl1dR4H8YztKLrY3Zi8AN8ECYqsbUVRN3UO5vy6NFMYUVhNWKcFgYziFAmTXBSO
Izr7AVU02kh8bEsQaSEObpQpC5gl56AO7q+h/U1SeFKm8wc0KhXs4ncQOOAPcj5+
M6BPe2RIBbVXlJu9arulevOEE6Zas8N69UM3maN190Spvs1+36QFNN191PUnjWgq
Ri3z5oXPCqjwePFYmuEZV1Y4HOgv68NpL6Boa9yVCTglTNfZLq6mve9Wy/BmcBwP
BvK2c5/5YBl3pnX5raTjLsSIq2k0EtPQZMVF/LI+nwEnFCi1P4A9GYHLrb0NA544
FgYExno6tV5q0+G/Ns5xrQSviFGGb1qN4g+0FtLVVyH1b7pI7fQkzTm3ZiFhHY4A
sVwMRMV1a04lZADbN12iwuqe4kZ+4AtYRP3v0AzUpNIcNTNJWOg6PgSg+KiCDjZ6
OCA7etjqz0EjJYfpag/sIJg5AHCwYUSBIRLHUyDJxo825alS//ePx/t7sQylMHGG
I3vm/x/9j2k9MQigTdT+iXw4pCJJByvxFlk/DuYsegY=
`protect END_PROTECTED
