`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BPX5LX8k/XZtzfYeyBaWt9qB1fTa3QOlBR55z7OmEFTx9HC6ymN3/jj78+wsETAt
whp19Dh7LvHDigIpb5SGVeTVD1ASQvs8/vQhw2+cxJykiDQ+jj4AyyA7de3EE38f
pKAyRV26kZUGypO7tbaxp7BY2+rHbI4FKGuBEiPGq3uJxCiWUwqoRM1dZc/pqd8x
1jg0W4Ji2/P61RFbSwGocbcCcHoQ3xBMr07fsqwcrMXn+29mWzeCj+TWKk2RlkVR
cPvIgCEYRLCGr4LjobdnrnZZGdGVPBEW7B90lIdh2qJTpnwer7h3+ndXzBwXbCnC
iEgi/Xut8Xl0HaX/8KtIcVMxyB1hbUTT9hJUe8cob1gwAoHoPqc7pLQoX/xwh5ft
ZY0rebQxzM9//daqhPYQsg7YRLfYSftsSr5ndjHdLWiYiieC1LDB5suqGMZw/M+3
7ANvThYG0nweoc4fJeIES6hUj2SFSMaG0hGzrzKt4yoU1FkNR67WljkMsRh2HrZA
WSMahs3nD820zjAWqLirUjA0CCxyQh5Txm3oezAdkNk53LjIo/WfBmGTux8STXD9
HlldUs11+rCyVK2x7Wx1lvvYMYlwXfnggnIjnsu0uPEfRZxro1wOfBhf8JXhjJii
JtPcVCaaRP15P2Bqp0oQUU2jN04IpC7jIQTXaoRQ/M6vIuUQUBb4xU+mXWjwikXz
b40k6F/8gQb9eUV1HToo0wYBGqIr6njiINyZ953eGO/T3zs8iheg1ZTqY3ZjGrEc
JPwXI+FCyMY7CSg/atqifNQ6Y3+3qBhX3DvQNBfPSU4/tbRhU3B/lmbAV4H+pnda
pAtKz805dy/X1Zc8om0Fdfr0i+wmEyOGLfuafj9aTdTTGHUXvdOubOZNdjSwhThu
BmZiHt9ie2+mEpGxinWvRSnLQHqvaw9goGlA9DRTwbJeiUyxxaD0So8Ws6V2pVTs
X9RJJxXo5gKhuChPNo7Mftdrws2mbJpZCFB1+JShbfumdkczAyp7kmcgG2COSoTG
b6cYDoI5cQuGUFlptWjqDXSQBjUYeV2kEN2FwGY0HC4g/4GWT+ogMcuVFPEFOAKV
EEzDRXhiz7aiA7Gnv07c3A==
`protect END_PROTECTED
