`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TEEOEQB05Rw86HlqRFkPLbVVtNdGTY+d6BLGIWJLpox/1i421Rreg1OXTOJ0bxRo
HSekOiZn5a4ed71jMzpAdY2pfk2UoFMTwiciwhjJTv1UsBRMHIgl9diullTzN4SR
X4ffcAjulhnJEutDe0CSyC+2rIq1jHyGFpI42C6IymLweSunXczqRU0qV+dudgI+
PL5DkTuLfZuN526OuJRVMgPp+CZKciNaJHFJ9D9voZ+ZEesUUbZsslIBfXquXszC
ZUNP5k9GFcldpc3+cPcX96R9Hv/yuvV8wkKg+5ohBvC2pVJ+vcWuIxGsOkl4E1F3
Iv7Z7Mr4Gu1kN0hlKCBMqx/W8prx4ahMndacCJjkbyQmnF1JKPeSuUJuA3kNjIhC
GLEJVqsEwj7JaX+YOiCfQQK2cxBSSda2l+WQpx7CDz1qV2JLRcJfj/K7WCIKAMPy
w5R7yeZ2Tuiq5bFJV8rMw2mlxPiz1tLTLBohbzdCe2DG5Y2/DT68rS5FnD90D7zs
PDns6Z9gKdgcoHxk9CMaAnxm1RJXEX9trn9h75pm6estxV4x4uJSm85txv4Uwxse
jdvIolbptFFtzLLhnI/lcVsbiagyh4h0VPxNClcfyrsGdzkooC7PsxXfGylgqVkY
/PWTuZBwplHFmHAR7+Qk1cd79YWf5fcde8pimcECIz77bcIYwnTWfXF3BjH1JfpL
`protect END_PROTECTED
