`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbCSa6gL5SXp/jj1xvUtIJn2Yic3xjYtxhPSvmtVdXOwHkN7m7NjmvfZepqFoTSA
FCIm8raUOSXoCkmbB2mKVmtupZKGc/xB9WmHKx90oLIFRiyoLuTIJZP6moNEfZ6B
j9mIoRWvXIQBBNhFr8CXvjHVxuJ29Y5/s01qnM2VS9meAeorn4NzDNNKAcYukAZz
dTYu5TLbU/mR3HcwuHneNcaQ8947lLs1RkKW9LYjPALLHFKe1C9Em522dLSkqZu+
YC8j4J/eP9IRzlZ9E8VWNgowS4um5AEAfnGblxJMx7WIJ5OR3jYLDMOTVLxvQ/Wo
H2IU2BF/XufxuBZW4yoqAnzEjK556DcRj1SL4sOGaNI3Ntkqx54gOTqG7oiGicrF
J3im/vxbCDWOfZAEEl3vMCwmtpqmCxoUduHsOB8p54gjEWXqQW+ZrKMoZR1ZEOC+
l1DH4KT1IrWWtk0bMbLHkhHyqK7yyg12hBRoOEl9B02g76yi9FAFOecwdMrASwjT
sdvQf2hkU9X9cvgJ08WdzU0G7F64VC3KYfmBNJVUCmX4yzl/Wp8XP3OV6YQzH0eG
RqwQ8AHEDCyfBqupY+qvMFN1zuAZhDMuV9YMMRlcUNF0PaP3wpwVIKEq3d0/RXGO
4REiodqG8A2CAcbuyESZZhEEK7FWpI9jO12zGuOfEH2y8CsQPg60it6aScgt7ATw
J7ZNsuQHa664wrqdV+/9HohRgA28gCnaqkQ1qZRTDTmG9FdyvhVqUZqcAq46rDL0
0nI5uCBnz3NA6w031FsZz/2mlOabgRCfG/LUYTwLZa8ZVS3zOQ5ROwwUfJgpmGhV
Ujtb0pK36/iHWAj2KAsvgzMyGzIvqN3sbtEogJYjI3inNasmSOms6C55mmrMvdHQ
yQGAqM0OnC+WLtwgMhWA18SiWt2FxpmgfhXnVdwCLXZsOlD9fPSY1k9K1C98x+s6
9uvDplG50je5n3A+UJC6ejK34iE4pPuThGXELUCfA+XQJKZAFt1X5YbEe4x+7dlY
d49Y+iS4aowaOmRCLBUKJS48VcLVCEbAI5J83vkXN6NaGRj/H2nMbZj1TOQa+lAv
XNyodqG4bGC3AeMWb+i+mP5S/UQXCkJyweOXqI25ZQDALEJ9d2mIj4d73UDkbzb/
0bFYmgU2kDt1W0PyVbO/XAcJJG9I4CZPAg3E8X6BbHEU2nUtGG2VR5Um9fTMbtT9
67ktncV0Er0xf7Qa3ryfxyF2/zihu1cBXjHUUhYyKqjNWLkPV4bRqopKJiW+PUuA
iuuzC7wJEH6r2Fhleq23PLxLiul8W0ZmwpwfW/gEeVdy77uZiGTUtitLqQqsZjTu
`protect END_PROTECTED
