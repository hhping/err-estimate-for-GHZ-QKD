`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6KROsChFx8SpsvPNpBBGR005CyXI7ZGqI1/2zjVqNuCVzlGtg56G6kzXgeB6wR+
AhNeEIazo7ZntaUGuhPkKJR6P/Vu1blOXpta4yGv0uDujHjmtvS0ZHP7uL5fYTu0
OjJOQ+tZ7giR8y+XH32QPeYiGmoDfeigRRKzc3MeU208XcN7C6EshVlFWI5MSJVv
dHu0qVwWLwBF59E/nSBPGERUCvw+c24scd9DgpnUBJMbZJAiEkCbwrehUCi6jKSG
UkR9RoEydkGPe+5WSuhhZx5o3b8VHuP+04ZQT9Y26yI+wJSP11uZJuLq+WS53jGL
yvVSw6BMrOo+3GY6KHp24sNSZ3YPA3M0bgL1cGMJFPK++xD19aAQidLgmZJsZess
J2Gw53DrSK3d330uifnzGTzt3cqeoRR/YKodalpb/FMJYy3ip4hD54FbBGWlDPMz
PoD35verMz+CFFSAubxJ5ct3iyNgdVgZqRlqjOfhZs+EnXpC0bOGUPDf8tjHeIbk
6GQZCS7TLHLHpv+63yOyaA==
`protect END_PROTECTED
