library verilog;
use verilog.vl_types.all;
entity twentynm_hssi_pma_adaptation is
    generic(
        enable_debug_info: string  := "true";
        adapt_dfe_control_sel: string  := "r_adapt_dfe_control_sel_0";
        adapt_dfe_sel   : string  := "r_adapt_dfe_sel_0";
        adapt_mode      : string  := "dfe_vga";
        adapt_vga_sel   : string  := "r_adapt_vga_sel_0";
        adapt_vref_sel  : string  := "r_adapt_vref_sel_0";
        adp_1s_ctle_bypass: string  := "radp_1s_ctle_bypass_0";
        adp_4s_ctle_bypass: string  := "radp_4s_ctle_bypass_0";
        adp_adapt_control_sel: string  := "radp_adapt_control_sel_0";
        adp_adapt_rstn  : string  := "radp_adapt_rstn_1";
        adp_adapt_start : string  := "radp_adapt_start_0";
        adp_bist_auxpath_en: string  := "radp_bist_auxpath_disable";
        adp_bist_count_rstn: string  := "radp_bist_count_rstn_0";
        adp_bist_datapath_en: string  := "radp_bist_datapath_disable";
        adp_bist_mode   : string  := "radp_bist_mode_0";
        adp_bist_odi_dfe_sel: string  := "radp_bist_odi_dfe_sel_0";
        adp_bist_spec_en: string  := "radp_bist_spec_en_0";
        adp_control_mux_bypass: string  := "radp_control_mux_bypass_0";
        adp_ctle_acgain_4s: string  := "radp_ctle_acgain_4s_0";
        adp_ctle_adapt_bw: string  := "radp_ctle_adapt_bw_3";
        adp_ctle_adapt_cycle_window: string  := "radp_ctle_adapt_cycle_window_6";
        adp_ctle_adapt_oneshot: string  := "radp_ctle_adapt_oneshot_1";
        adp_ctle_en     : string  := "radp_ctle_disable";
        adp_ctle_eqz_1s_sel: string  := "radp_ctle_eqz_1s_sel_0";
        adp_ctle_force_spec_sign: string  := "radp_ctle_force_spec_sign_0";
        adp_ctle_hold_en: string  := "radp_ctle_not_held";
        adp_ctle_load   : string  := "radp_ctle_load_0";
        adp_ctle_load_value: string  := "radp_ctle_load_value_0";
        adp_ctle_scale  : string  := "radp_ctle_scale_0";
        adp_ctle_scale_en: string  := "radp_ctle_scale_en_0";
        adp_ctle_spec_sign: string  := "radp_ctle_spec_sign_0";
        adp_ctle_sweep_direction: string  := "radp_ctle_sweep_direction_1";
        adp_ctle_threshold: string  := "radp_ctle_threshold_0";
        adp_ctle_threshold_en: string  := "radp_ctle_threshold_en_0";
        adp_ctle_vref_polarity: string  := "radp_ctle_vref_polarity_0";
        adp_ctle_window : string  := "radp_ctle_window_0";
        adp_dfe_bw      : string  := "radp_dfe_bw_3";
        adp_dfe_clkout_div_sel: string  := "radp_dfe_clkout_div_sel_0";
        adp_dfe_cycle   : string  := "radp_dfe_cycle_6";
        adp_dfe_fltap_bypass: string  := "radp_dfe_fltap_bypass_0";
        adp_dfe_fltap_en: string  := "radp_dfe_fltap_disable";
        adp_dfe_fltap_hold_en: string  := "radp_dfe_fltap_not_held";
        adp_dfe_fltap_load: string  := "radp_dfe_fltap_load_0";
        adp_dfe_fltap_position: string  := "radp_dfe_fltap_position_0";
        adp_dfe_force_spec_sign: string  := "radp_dfe_force_spec_sign_0";
        adp_dfe_fxtap1  : string  := "radp_dfe_fxtap1_0";
        adp_dfe_fxtap10 : string  := "radp_dfe_fxtap10_0";
        adp_dfe_fxtap10_sgn: string  := "radp_dfe_fxtap10_sgn_0";
        adp_dfe_fxtap11 : string  := "radp_dfe_fxtap11_0";
        adp_dfe_fxtap11_sgn: string  := "radp_dfe_fxtap11_sgn_0";
        adp_dfe_fxtap2  : string  := "radp_dfe_fxtap2_0";
        adp_dfe_fxtap2_sgn: string  := "radp_dfe_fxtap2_sgn_0";
        adp_dfe_fxtap3  : string  := "radp_dfe_fxtap3_0";
        adp_dfe_fxtap3_sgn: string  := "radp_dfe_fxtap3_sgn_0";
        adp_dfe_fxtap4  : string  := "radp_dfe_fxtap4_0";
        adp_dfe_fxtap4_sgn: string  := "radp_dfe_fxtap4_sgn_0";
        adp_dfe_fxtap5  : string  := "radp_dfe_fxtap5_0";
        adp_dfe_fxtap5_sgn: string  := "radp_dfe_fxtap5_sgn_0";
        adp_dfe_fxtap6  : string  := "radp_dfe_fxtap6_0";
        adp_dfe_fxtap6_sgn: string  := "radp_dfe_fxtap6_sgn_0";
        adp_dfe_fxtap7  : string  := "radp_dfe_fxtap7_0";
        adp_dfe_fxtap7_sgn: string  := "radp_dfe_fxtap7_sgn_0";
        adp_dfe_fxtap8  : string  := "radp_dfe_fxtap8_0";
        adp_dfe_fxtap8_sgn: string  := "radp_dfe_fxtap8_sgn_0";
        adp_dfe_fxtap9  : string  := "radp_dfe_fxtap9_0";
        adp_dfe_fxtap9_sgn: string  := "radp_dfe_fxtap9_sgn_0";
        adp_dfe_fxtap_bypass: string  := "radp_dfe_fxtap_bypass_0";
        adp_dfe_fxtap_en: string  := "radp_dfe_fxtap_disable";
        adp_dfe_fxtap_hold_en: string  := "radp_dfe_fxtap_not_held";
        adp_dfe_fxtap_load: string  := "radp_dfe_fxtap_load_0";
        adp_dfe_mode    : string  := "radp_dfe_mode_0";
        adp_dfe_spec_sign: string  := "radp_dfe_spec_sign_0";
        adp_dfe_vref_polarity: string  := "radp_dfe_vref_polarity_0";
        adp_force_freqlock: string  := "radp_force_freqlock_off";
        adp_frame_capture: string  := "radp_frame_capture_0";
        adp_frame_en    : string  := "radp_frame_en_0";
        adp_frame_odi_sel: string  := "radp_frame_odi_sel_0";
        adp_frame_out_sel: string  := "radp_frame_out_sel_0";
        adp_lfeq_fb_sel : string  := "radp_lfeq_fb_sel_0";
        adp_mode        : string  := "radp_mode_0";
        adp_odi_control_sel: string  := "radp_odi_control_sel_0";
        adp_onetime_dfe : string  := "radp_onetime_dfe_0";
        adp_spec_avg_window: string  := "radp_spec_avg_window_4";
        adp_spec_trans_filter: string  := "radp_spec_trans_filter_2";
        adp_status_sel  : string  := "radp_status_sel_0";
        adp_vga_bypass  : string  := "radp_vga_bypass_0";
        adp_vga_en      : string  := "radp_vga_disable";
        adp_vga_load    : string  := "radp_vga_load_0";
        adp_vga_polarity: string  := "radp_vga_polarity_0";
        adp_vga_sel     : string  := "radp_vga_sel_0";
        adp_vga_sweep_direction: string  := "radp_vga_sweep_direction_1";
        adp_vga_threshold: string  := "radp_vga_threshold_4";
        adp_vref_bw     : string  := "radp_vref_bw_1";
        adp_vref_bypass : string  := "radp_vref_bypass_0";
        adp_vref_cycle  : string  := "radp_vref_cycle_6";
        adp_vref_dfe_spec_en: string  := "radp_vref_dfe_spec_en_0";
        adp_vref_en     : string  := "radp_vref_disable";
        adp_vref_hold_en: string  := "radp_vref_not_held";
        adp_vref_load   : string  := "radp_vref_load_0";
        adp_vref_polarity: string  := "radp_vref_polarity_0";
        adp_vref_sel    : string  := "radp_vref_sel_21";
        adp_vref_vga_level: string  := "radp_vref_vga_level_13";
        datarate        : string  := "0 bps";
        initial_settings: string  := "true";
        odi_count_threshold: string  := "rodi_count_threshold_0";
        odi_dfe_spec_en : string  := "rodi_dfe_spec_en_0";
        odi_en          : string  := "rodi_en_0";
        odi_mode        : string  := "rodi_mode_0";
        odi_rstn        : string  := "rodi_rstn_0";
        odi_spec_sel    : string  := "rodi_spec_sel_0";
        odi_start       : string  := "rodi_start_0";
        odi_vref_sel    : string  := "rodi_vref_sel_0";
        optimal         : string  := "false";
        prot_mode       : string  := "basic_rx";
        rrx_pcie_eqz    : string  := "rrx_pcie_eqz_0";
        silicon_rev     : string  := "20nm5es";
        sup_mode        : string  := "user_mode"
    );
    port(
        avmmaddress     : in     vl_logic_vector(8 downto 0);
        avmmclk         : in     vl_logic;
        avmmread        : in     vl_logic;
        avmmrstn        : in     vl_logic;
        avmmwrite       : in     vl_logic;
        avmmwritedata   : in     vl_logic_vector(7 downto 0);
        adapt_reset     : in     vl_logic;
        adapt_start     : in     vl_logic;
        deser_clk       : in     vl_logic;
        deser_data      : in     vl_logic_vector(63 downto 0);
        deser_error     : in     vl_logic_vector(63 downto 0);
        deser_odi       : in     vl_logic_vector(63 downto 0);
        deser_odi_clk   : in     vl_logic;
        global_pipe_se  : in     vl_logic;
        i_rxpreset      : in     vl_logic_vector(2 downto 0);
        radp_ctle_hold_en: in     vl_logic;
        radp_ctle_patt_en: in     vl_logic;
        radp_ctle_preset_sel: in     vl_logic;
        radp_enable_max_lfeq_scale: in     vl_logic;
        radp_lfeq_hold_en: in     vl_logic;
        radp_vga_polarity: in     vl_logic;
        rx_pllfreqlock  : in     vl_logic;
        scan_clk        : in     vl_logic;
        scan_in         : in     vl_logic_vector(9 downto 0);
        test_mode       : in     vl_logic;
        test_se         : in     vl_logic;
        avmmreaddata    : out    vl_logic_vector(7 downto 0);
        blockselect     : out    vl_logic;
        ctle_acgain_4s  : out    vl_logic_vector(27 downto 0);
        ctle_eqz_1s_sel : out    vl_logic_vector(14 downto 0);
        ctle_lfeq_fb_sel: out    vl_logic_vector(6 downto 0);
        dfe_adapt_en    : out    vl_logic;
        dfe_adp_clk     : out    vl_logic;
        dfe_fltap1      : out    vl_logic_vector(5 downto 0);
        dfe_fltap1_sgn  : out    vl_logic;
        dfe_fltap2      : out    vl_logic_vector(5 downto 0);
        dfe_fltap2_sgn  : out    vl_logic;
        dfe_fltap3      : out    vl_logic_vector(5 downto 0);
        dfe_fltap3_sgn  : out    vl_logic;
        dfe_fltap4      : out    vl_logic_vector(5 downto 0);
        dfe_fltap4_sgn  : out    vl_logic;
        dfe_fltap_bypdeser: out    vl_logic;
        dfe_fltap_position: out    vl_logic_vector(5 downto 0);
        dfe_fxtap1      : out    vl_logic_vector(6 downto 0);
        dfe_fxtap2      : out    vl_logic_vector(6 downto 0);
        dfe_fxtap2_sgn  : out    vl_logic;
        dfe_fxtap3      : out    vl_logic_vector(6 downto 0);
        dfe_fxtap3_sgn  : out    vl_logic;
        dfe_fxtap4      : out    vl_logic_vector(5 downto 0);
        dfe_fxtap4_sgn  : out    vl_logic;
        dfe_fxtap5      : out    vl_logic_vector(5 downto 0);
        dfe_fxtap5_sgn  : out    vl_logic;
        dfe_fxtap6      : out    vl_logic_vector(4 downto 0);
        dfe_fxtap6_sgn  : out    vl_logic;
        dfe_fxtap7      : out    vl_logic_vector(4 downto 0);
        dfe_fxtap7_sgn  : out    vl_logic;
        dfe_spec_disable: out    vl_logic;
        dfe_spec_sign_sel: out    vl_logic;
        dfe_vref_sign_sel: out    vl_logic;
        odi_vref        : out    vl_logic_vector(4 downto 0);
        scan_out        : out    vl_logic_vector(9 downto 0);
        status_bus      : out    vl_logic_vector(7 downto 0);
        vga_sel         : out    vl_logic_vector(6 downto 0);
        vref_sel        : out    vl_logic_vector(4 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of enable_debug_info : constant is 1;
    attribute mti_svvh_generic_type of adapt_dfe_control_sel : constant is 1;
    attribute mti_svvh_generic_type of adapt_dfe_sel : constant is 1;
    attribute mti_svvh_generic_type of adapt_mode : constant is 1;
    attribute mti_svvh_generic_type of adapt_vga_sel : constant is 1;
    attribute mti_svvh_generic_type of adapt_vref_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_1s_ctle_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_4s_ctle_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_adapt_control_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_adapt_rstn : constant is 1;
    attribute mti_svvh_generic_type of adp_adapt_start : constant is 1;
    attribute mti_svvh_generic_type of adp_bist_auxpath_en : constant is 1;
    attribute mti_svvh_generic_type of adp_bist_count_rstn : constant is 1;
    attribute mti_svvh_generic_type of adp_bist_datapath_en : constant is 1;
    attribute mti_svvh_generic_type of adp_bist_mode : constant is 1;
    attribute mti_svvh_generic_type of adp_bist_odi_dfe_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_bist_spec_en : constant is 1;
    attribute mti_svvh_generic_type of adp_control_mux_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_acgain_4s : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_adapt_bw : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_adapt_cycle_window : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_adapt_oneshot : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_en : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_eqz_1s_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_force_spec_sign : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_hold_en : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_load : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_load_value : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_scale : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_scale_en : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_spec_sign : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_sweep_direction : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_threshold : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_threshold_en : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_vref_polarity : constant is 1;
    attribute mti_svvh_generic_type of adp_ctle_window : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_bw : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_clkout_div_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_cycle : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fltap_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fltap_en : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fltap_hold_en : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fltap_load : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fltap_position : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_force_spec_sign : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap1 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap10 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap10_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap11 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap11_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap2 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap2_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap3 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap3_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap4 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap4_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap5 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap5_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap6 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap6_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap7 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap7_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap8 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap8_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap9 : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap9_sgn : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap_en : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap_hold_en : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_fxtap_load : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_mode : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_spec_sign : constant is 1;
    attribute mti_svvh_generic_type of adp_dfe_vref_polarity : constant is 1;
    attribute mti_svvh_generic_type of adp_force_freqlock : constant is 1;
    attribute mti_svvh_generic_type of adp_frame_capture : constant is 1;
    attribute mti_svvh_generic_type of adp_frame_en : constant is 1;
    attribute mti_svvh_generic_type of adp_frame_odi_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_frame_out_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_lfeq_fb_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_mode : constant is 1;
    attribute mti_svvh_generic_type of adp_odi_control_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_onetime_dfe : constant is 1;
    attribute mti_svvh_generic_type of adp_spec_avg_window : constant is 1;
    attribute mti_svvh_generic_type of adp_spec_trans_filter : constant is 1;
    attribute mti_svvh_generic_type of adp_status_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_en : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_load : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_polarity : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_sweep_direction : constant is 1;
    attribute mti_svvh_generic_type of adp_vga_threshold : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_bw : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_bypass : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_cycle : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_dfe_spec_en : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_en : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_hold_en : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_load : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_polarity : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_sel : constant is 1;
    attribute mti_svvh_generic_type of adp_vref_vga_level : constant is 1;
    attribute mti_svvh_generic_type of datarate : constant is 1;
    attribute mti_svvh_generic_type of initial_settings : constant is 1;
    attribute mti_svvh_generic_type of odi_count_threshold : constant is 1;
    attribute mti_svvh_generic_type of odi_dfe_spec_en : constant is 1;
    attribute mti_svvh_generic_type of odi_en : constant is 1;
    attribute mti_svvh_generic_type of odi_mode : constant is 1;
    attribute mti_svvh_generic_type of odi_rstn : constant is 1;
    attribute mti_svvh_generic_type of odi_spec_sel : constant is 1;
    attribute mti_svvh_generic_type of odi_start : constant is 1;
    attribute mti_svvh_generic_type of odi_vref_sel : constant is 1;
    attribute mti_svvh_generic_type of optimal : constant is 1;
    attribute mti_svvh_generic_type of prot_mode : constant is 1;
    attribute mti_svvh_generic_type of rrx_pcie_eqz : constant is 1;
    attribute mti_svvh_generic_type of silicon_rev : constant is 1;
    attribute mti_svvh_generic_type of sup_mode : constant is 1;
end twentynm_hssi_pma_adaptation;
