`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Pd1pMO5jgLYZTTbPlAwNmIej6Xv34oUDtgTdyhoteS9jcitY40CT8EBFqI/FfbW
TVy2MlwDy0ptqeLOdUY/4eOVPjBG+OkMQ5pdaNmZ8zOabd3xf8mvUp1nHKm0Tb0S
zF/Nwt3rF5pptT9VAdqs9o4ng9cSZvSXQMG0jOBn2VsFI4G6ZyptXUCdlF44VJX6
9MLSu0ipSGAFFxiwkVlfbdTrt7MsZ+fZrF+8HAjl8i+qFBo01DCuiZPUflOs9YZ/
5S41TMc41PTWEe6hig4QO91m9VnPt5KLnGkE0yiGEcTSQU4PwSPcsVr0APcbPbxI
JjfgmqV9jh+NJW1MgAvNNhIzz1qOMfZUtgVquhq5Yc5cbXPlG0colN1vAKnw894g
tsODD5srWoohOISS6dfbzcbMTd0XtP2nbusugp4ZVeY=
`protect END_PROTECTED
