`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XhHql8hazgt14LnlaYoDiuiNC2HhQbXXZstvRiRGdzo+3Q7FsL/lzThSBnquYbNw
w8um0kO/N0NHX/oyOfx9nuqAQXDjE+XgLyB+g21LyGj47RQNEyd8meTcYPy+cU1h
DpHH2xYwMu28bgOu1has5s1iiV4LfzKRzBFEPAk4mus6yvPgl2/SwEPUKsQbPOSv
a6sVWW29zYzrHC0KLZ/Eh57540EqpqJ19r/civpFRXYhN1OruaMd2KZS8uYuVFo5
BFEZbxEMi7ohS1MpetlhCVqcRHmxqWjxeYQIqnKGw0Cwd/M5BUd2ydsBrQSTI4QD
/WQ5e2yDcUB26m7eEvnPvixiw3AHQnsOg+G3sxQCiIHu9nS8H4b99dbc7MVOqE2Y
KDiYnLb//74lS8ChB1ueuLFWsz7f3VNJ07JWm+0+9zpK6exLRuMOhjgQ1y0s6XSs
gIFRs6o4HioWAvD08bY5Hx8FsFPvphg+6yQul7xt55kPA76rxuy8qCqEOjgH+Hgf
IjWLh2ouIuHF8ljNoF4maGLVbb6F5FspoXp3thY4SCgqlxWKC0jgiq/sieWSOCeE
Ej0QCiF30TZ/Hjcknpb2bk8TT5dqC2zqnCSNtOkOUPJbV4VA9tv1J0zyOxPpvXOf
hcFtciKaENQCP5V8lfUGbmEKwKhcgdDZTsJ+BcHGZmll493VMMwh5vHi4imRRmDZ
bbwzsy8AAB2PY8ECWYGyoVOfS06glXgglJz7c6h3ARGGZpERhQXckd5vaZL+IS0j
36p1uJR2WBkSTDkE1XyvK6/RKY8JPpVkk6NXswDKQsOJavbwhir4i0D0BZUignmX
PrMSrQ+lEFOb2gOsfhVgoz3uDyON0GQZk+m0Cec5K6vCLy/a/X2U1WFuwQc5JSX6
nNpp/+3T0gLaSuE5sSuNCLH05g4J6fyAmCT2Nnhpac9XiduurVBsA1k2IKNqvDmL
+U7eBAkE9/7XA1F8LtEMSTZXNb2E5dxHFSJiho1aH+5OaQ6z1JCDpSokLQtPUP68
gNN+BAHy6Dw98L5+PrvkpjQcTBM2qUodRX9nJ313b08XIk7CRpbHOlQh9lKNELFi
mQRZ24oM0o+m/ByMVt/an4CWW5zGm/GHwNAbgaIK6acikeDELxD3VyGApa6K1frn
Z3c/+ezMa35OQV478QlhNsgxx/YOs5pWYaRN8pni/Y1WvD4t+8ZBrp5ygybrsKgw
aLYfnEyFNIaerl6WwrlM6oIH4dOMtEMjAVZ45gBhIGUlWZCwpBlMjWuPbvCGKplD
xKWn6Fg1THK0lED8Fu/fP38xuW0+oYDUfWAI5/SvJ0LEDodLIHbMRHXAkjxJ8tCG
1mmxuWnMapOvjOlu5b9VvPY9vkSwJ1T369Bxup7y9H3X+u4FkOP4kui/SYFZXQbD
LkA8HgVMFaTTBbIx84vuKFcqKbsMbHMr0vj8mYqwSgwLqnmxZPRLl43jIjjzpZsT
c8KMMGXLy5RC6iAHYJEaE7EC0JMqEbJnTCSUFfq08Tu3gW7NTE+o8qDHDaZotEHj
0ZXKCZN8g3Gb2xv+OB3JDqc1M2UCFPB0D7t/0lpmQExQfu/iUAip/vnD4BC7uvZk
vuutfdLsIB6pBfDf4OHIJiHg+o5ZQdZfNBo4rQvGx8LALIM2IViaAfJ3ERKOjNqF
4co9gQwZpdeTIVBguQI7z8Eo5y44b892Ee/D224kcZ6Ivr8QpK9u/xHFnZiQC8hr
MUNd8LuXMB0KJTdUFoAVX/nclcXomODdBINcPbiGQWoJWaP+EbJarzSar+mbTXq9
wi312SF6NFsfgNH6Ui6uChhI0Jd4qK29YlbBsD+W1nQ2hZKcdJIbLT+KgD67nGvs
bcMfBHtFBBj5wtvNhfsPFNqjbee76Gy/zyLqIWX2i9n45mK8tMvT6Ahg1MhSsA5+
TjOdHHjkzURIck4T+1x5ii7AaoO/mc4p+AuiDsJCC9Ys2nPitbbsl4XfpMznm8aA
kero/F6UidQr2XgbdBaH9Orshhs1ZB1I5D3bhmJK/aJtMJlgQRnVtbdMJGI04SJf
6qu7Qhta1OvKOTde2R2ffau2uvssquCOmekSxaYNFUd6Y+4AZKyTeOgLbpgTQMNJ
zmRfG65VlYTcBHtTXXdxoRnt2oulPMnt5/+OLEG8cU7sa4NlU47sn9d1ARmy54Kn
YGS4OWZNY3Wnm1ZBmmwQYwbcRB9/fMyDCVzkNik2y+0hJkJcxgxmpljvncBJ6u+Y
eWrRXkpHi0OqySTweN1Apit4XQT7ugFB32XLuYvBEvFWS9UdRCxbQBEQVmIuMgUl
inZL6je4us+qr0G9YkbizwKKcQ5IH3EdN4gF8m8FSMvXBlVVKXLQ6ucbZEa01MU6
`protect END_PROTECTED
