`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjqgBmgTUBCzPbc5lNrH4dUSTybH/OnEqvFhwwQwws2OMxHilFNpebTU9WOA8YSS
rVM6zM8FFclJ1qqAbkN4gFAOng4P8lkf7R13Mhl6Zm14F4JD14i2kw+RHK5smrvy
BTAdsC0VC7H07s1TE3+CS12SsTD0eWEp7Uu0JFX+50lDjgSgZSqLy3l81duNvb/o
1xS+rrBj13OHT192RuW/S2Fwa95AuSFBLvr82zNOO9VQR5LMI9ptiD5J732UfEfb
d1XQIV1gGT2b6WMWmBHHiJEu1lu7arU8joePu1cQIoRCyUjceQjfE9zgwl8auOgK
65roL79q7qXm6eK0OM7ecP+pFiI1imX1H+E8Pr/MCVXXcvDBrFt1UbhWSy+eVgW2
T5JJ3VX6bX0HiSXvY/x6F+ExZTe+1ppAOwGh99paa3eaL+91utWo1RpZUbNNRPFZ
vJ7WJsfSTSqUo3eg3CYB6A==
`protect END_PROTECTED
