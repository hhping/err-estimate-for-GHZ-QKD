`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JefcotIoTdURPe2/mSS0hl5ZCPKVYVm/XSxqQWSidjkww16xy+3SPe2m9BrbaaBD
AlCBKruGboEdD3mpyz18mOyfwy0eLHQkKCu0oGIAS1zjnlSNKn/B2FyUOOmHCvY3
MtH1FirXv3mCaYrOnAqHz7wdxPrtpRvH9N+mRm3lNgcIVe+ApltQWEOTWDzDIjmG
560tkcSSL5CgGn+evvvfSPtbSoVsFZvs64JHkmsu//aqqJHbZYeoSYl+Q1Qife1p
Qk2kDT1POaUrT4hfRZpAzqwmPjLf1mI5fnHXCJqnfHcPaArLCCuoSdd/IGaSI3VJ
83idbmezSPJ5iJSwmUj9EawS5Jvcr2Om3TLhfPJUUphwsSjyUNMvQCGNZsn8yh+s
WjC2M34Qz+uec76qcLUKv0Vo74GSAEvr980G/WLyNqUQ2fgIBHAs80E403a5eCFd
heVPdTmo3wJH5UDnM4xx0CjqaqoA3qa97SuYL0OV0P80F1IpGFQRBAOqaykbmz7o
05y70A7UkhZk4RVX/V+lzg7xeMY4SNOHtjb3keYSyhwq543jD7Hejo7olJfjz61o
y5XxPJ8vgtmD43QaqQ+LyNbz8QaNGBhXp0nVlPt6J6FXUoEAGWv8JR232MYpaeAZ
G1wyaRZqiqOIu28n7+NFT0XrL8SWEMXr0b11KgZRmQ0mGrzTIElZta0Awo4uNm0U
6ASHKkSPS5MmW10M5+dZFkwy9NeFlkTVfvU5wYdQgW0oYZqBw7/snAAUFFN9hJYx
FtWtO6bm4wBLeMvSp3GZUXD7+NgBYKXolC1kHLlEW6VUKPOvt/NO6u4xqmBSXtu4
MGUvNhfTpUeZTM6yhBSHE5Qu5xUTBhdL+ZCPiFJ0yo2jRe1z+8mQMiNMf8JPLctc
jXveFhxZeAsqlM1SgGG/5Va2QOvY8vBWF1sIV/ART52D0yr0Wrz6U+8qX32ILxJJ
T/KzWlcqyElYXNaBzBceqT9x4aJH0sn+57YxexaM2q4Ykha9QobczdSw37oFV+B4
6v5CTJ/GK3rtHgWryBCzl8OdQS/KCS+BmViEcSToj76FSbaMQ8gMc7JPJFSxS0i3
Hzw+u4g+Srys/WEKnxT/3j8gNkceOLtLWPmbW4pOfvjddscliv6iT/Ji6Dj2VHCZ
nuZCY+0hGVR9G9q0ARImt6Pt0UCIbod8PVuTYKq5/p7mtioXpou9ID8BbbfyUYKO
nLya0nGspjVXgsl4xpglXIoC+pCAWotrKEguZfipdox8vPp+dxQ8PGVfRITp5h9m
WugTyn4pfX6lsofw8GeB/tbc4r4keuAzPoZZUHTlcIda1TyDKmB1Rb0dzuBkFVCL
E4nYR+aqXAPnFa2UgY2dBxjvzq5tzK/QhQppIbqG1h+6oRtIBODjvKJtQXw73qaT
aZ8Ii2HC2GHB89QepDchr4glqX/DDUV97Nel3lNHmy8haEM3PefL3eUtWKcz/ATM
bPfqr8EbnCp3O/b2pK7ZaN/3WdGEqkfAFxC34iIWLI4rKb1DW9Mz8sKxfzC8eYq+
59ihhh7Ygu9hYgHQpat2xhfWu3lU9ZAbmFdZ3+7ML6zMIzduXZTSNXOK47eed93d
KSx5U0XTtEWNl/1DIBaq4/++dS0UxM+GVkwmKqa5r4cGgOOskikQkYtlDZv874uP
bhThQ5avsLpSjx8w+emjxQHWwh1V2AJpVMQRcj6eDesyEdXTuFs73RzdJnkExrt9
nUo9vQI5ZCFaAvDS12rxrm/EZr/w/1NJaSU1QT9NKYehgwv0Vhy+j8ObvKkoYzor
CB4UGM9bnqloqY9Jdl/5ElL0Ue/lUfcV88Zjqakra81tb4d2/Jnlc3ywpWmJbC2v
Ll4l1v3SW/sJT1r32+Wn6/2BGSwc26A6zVsxI38x9pIFLlsybPmqLdbGCbONpOHm
QiOyaZ/RifoOxnnsbbCBx4EEasBNb3Y1b6qC5VeIFPA6jydhYoMKmWKDXvlgpkQt
oF7ZsTmQJ0kl3K7LQA91pp3QhDdYzzTp8v3/yOyBItUP9mGjVt7JywUyB+vldTCh
R5H9Fu9PXfehZ+HmpHNR7pFDytdN4rL/OUGYOUsdVVTo0TKOUg1EwEg5qwopSQ45
AxZCquiY/o3aduESEEFu8N6xxxaOP4pTyqbKORwW0yYZoNhTXzkUKn0p3019TKJE
PRt0jbaiIAJb26kXK9L6B9SLBMB5HVoqkh7qd3dHqrjU/gmKZ8cAaDoJhoqzBr8v
zC0sxa4FEIKVD2enf+xPWJLB5Xxr2pT34Wq7hnTUZWGYwBD9Ob73N4FDzgd6Wu9j
eCwLpsXA7OHAbOodSSocgqgdbUAcQSgwxoIDa/n4l1fojC5nrmGjSlLdlKL/9F8O
uylSaZwwUbzIuYZd1Fiq6YhGC06LkKUpubA/O4uPe8402RP48KIMHLAVHdRZT9Z+
ORtQcfH272CNogLNLkJ287VO1ZBcCkwtv+2ZTA9CH5lsqSbhEX7fxKUQCICfWXrZ
R5cH0c05WOACNedGCKTWzK1rNxlUYKcFpfOl4EThmlR5Iaw7il8w9xhkJiwsJXVA
olauf3TdSmm/q533n0OkvnICYutxofDEPnVlxiEcxBerFsVAJEetUT+9lJ/YXeRB
i47EtdOpsgDuUfWrN3YHhj+g399VjKjEByVLurCoJglrc+B8Fkut4clwWiZBF4pb
qhIy0VN8VDgkWkBvPemMm/3NH0W8Rr4YWwiopdYKs6FUuGOKEb7bnJ/ifDIcTn/L
2dLSU4pbs7gngraw6lVYY2WU7Xw+6VpVLWfMhRTPQOpcOxdzXYcJoehnRZOSgrq4
L57Zjq4XixEppk6mkywlvqzT6haGLrvqskjGtroi9WMOtSown41YNR5Ic/SOONbq
/056fMyQisV2GOK1ZrIPP695sGLZuBnGM1wKPxTvIebS64y4qjf4ghf7X2HKWFAa
+RlbXsylTpWXIcJvMDe3QOGWCi6mDxoy7nIkuXOR+U6WHqaxUF1h32Ny5z2pDSX5
nN04e9HHQdBnGVVF7Tt4OymbPURw8Gg2aW99k8ViJ+23G9YNEsL3VfPqc5bFbwpX
2wiJ1HKDy+gh+bR1nnZKej8wbfD0h4hB6qJgtf4RXY3tNCDytFpEuFgMQXEMV/If
SzW+FlWR7i+DKFS/9gPndvyeqAZ82+gDXnOHCx/qKgxviLNqzSxkV/D/+W8T9sfC
XDFJ2wovZ7wr01eHKZy99pQb6z0qJsvbwzFvc3F0ILcK+3BBq1AqGSbraG9HoPYZ
PQn1mLXPXv+34PbVHdNLNFjl7DnsnAFN+5gU1UgQ0B2steIKEACwe1o952vwvHz9
h4fjPzGI6LN2C8USQqaCgrVCypUWndLI8XFZwFteDR0J4MIIGLp6LaxR0AWgQJHl
3OBE9y45ptQcja0fhLGZekF5z8j96vSbJBjP0NHOLYkQ2J2FqVAM/Ji+Bt+aI0EY
ldB/uA+clJut9p+ImtsoFPCKRL85ysHNtlQlOK2MxgWtchlX4swMWPTvrsQkvLYK
98a5PKPH8uo0Zl2St8zjzLikj0plVJP/tE++wbtKnEJ6pcn/7u3zk6z6YdUAMu4G
pQ2CcrYg01fNtgrI7y3qkVu36PNIlC0ZvpsLmnn7QRBDIQLV0s3joJ3Lq9XrOCMH
Cjk8RslGZkaMj3wJGh0Ggdf+LlYY/Y/pbJhpTukh79HQDqTUTkyZ9vwr3sPDrEUn
1kiq5GJl+TWyy3V1nvvLxoL5bwV63O3DT3u8RysSHRMeBZfHTXIrXCjX+RmUBiyx
eWcvbkDycUJ4gl0ik56RWkjBMWuGS3NQrLHTjrc/iF2S0dS3w79dtlYMXka9vCi+
TKBxUrvyu2hHcNyo3+2i6XzeynG1Sax1W71RX4b1I8M+L07LzeEJW/rhjKe/4gjw
EHMGX+iPgs2JrwvRjlQ+0EfeISHN+V9829phnm5a0TWn4R6pauP6gjFhU0PNCakk
ducHykapi6Fjn3ttl65T35m+7YXQgPn6Tmiwbw2xtlEOJOp/UCpxxsHDxUSfjwzp
yRdWRPD+1Du3OzfvrGFt5McP3Bjn1FuPPMQ7KZ8pN4gnuTRMsBANZCDng5ul22za
ZNUmrsFWFbZzfHUxjXCq4w==
`protect END_PROTECTED
