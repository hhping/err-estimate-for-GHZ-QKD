`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
428liZv4nse0LANfD7fCJIbpUjB3XFw/WytqmRWMjPnwpvAcIh+1JVZCUMBP+8Tj
2gop1n1+HfoWWpKbrdJdVbDgcLy/Piy4cPTZiIqqX5IY3GuF0gMWXQF0FwV1K6nT
eHLtmznazz138COSs0szaSKu9P67ATGxR8GqBNZMLBhVO0oH1n+c+ammqnLigjN5
4qp8WPwyk8k4UyjRoPvRDTjzz0lRhp/Z3DP0e7z6YHQhinhUaUpqG85+EY9HEYAO
0XiYQxwIroNH7rY7MiV2LT/wUY0Hkgl/UG/QdN6m+bDudIZE2r5F0IB2C02uheAP
hP3y9QGNX8OHkVr80FPWQouCWHZ84ll/o+LkFP7argsugTSiE7IJoQ5K+VdB3CF8
`protect END_PROTECTED
