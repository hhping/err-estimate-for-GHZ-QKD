`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rf2weYyRK5QGDXI/eDNewsHLgygDrnuB/lwduBRaeDQ7yjcQj6TlmmMtntu8as3W
ek7e6fWYO2347couRWRsFQ3QBRQpSWc6+23w7HXYU+tPW6o+gkUeNlPnvXR9zlQ0
rgNQewGNS0gggiMrlp7ZDWh1E7it+28JKXsvJaDyHcG7t8Z3X0cUPLXKXKfM2xcj
T2f9/qnwYFVMFrloa2wCP3hCnIBeA7tFpJEbANSBFCUsELsFDt5w1/vEdeTYTffK
KmSTYQ96w4ldCq7E+LesAQySrasIetqTs9nEtKbE6oBzIicKl4YSfbQfTkyt+Mg5
PTWWL+c7yJKuju+iXq2zjM8iurQYTzafAUweRD6VU9+E1MmrdaNzB6q/bG76AIum
omSPyTCsDWSIndxCekN2luyF4t3CIL97rHHU4qtvmd93gxGgpo44nVQWZZcoAnxQ
qZ+8O680WNhfXbFPvU+6pI+mMrAn5GMfRZwxxo9FbidfMayh+k3cmyJr9t6xXZyr
hxLZnmBDzrebQUJ+5bHqHw==
`protect END_PROTECTED
