`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QW16zbMsMv81DJCI4OCxFM3l5zuJw7npZMTOjtaPDJkT2bs6mNZHDGhEHYQT1WJD
yNJPm1tMfNhVBmx/ozY1B+A89THBHHus7K3wzRWH2BDcSMtMAQfQfZ7wqcWOthjR
om7G8TNE40sGDgiRPIt+jK3casCc6YlUROCHXApYz3fAEGXI71wapLTTLVxe2GdM
Mo1Mg15QNjBtDJauPDTGjoqSXe7nR0bjsMkqtJSsfkSmTJHH3DdwXZ+XapYkUNLy
dB47vs8pIQaCf33zXp9g8Cl9xBHKCERSO7/bSnd4zLePvDKVY9gJUf5esGLAX5sg
yZ6sT2gmwk+zWy4PguyuF/IEocylnSh25aR+YNfen/7m2K6CpKhJFo7b/o8qs4U/
XIgZ31xBHsgP087WLnU7bGHWs1FHDAUvpOuJVPoPXEOT6KJJPT6qvteequ0YBUrF
TL/aqnD8wPjeTdVsT4OwdMh3XX0esWBUFdsDkE/S+KfIp1o3Lp9gows0Or3A2jt2
+2TvAZPXIDiQZVPoVpk4RZUJ8p1GeJAwFIySEpHpTSYe1pyabH4N0xt7SvC/MvTt
8yPlAtYzhd/SOMuIZlm+WXE5F6UesWjaF9GblFZiZZsPcuTms6tHs2QlNBwaG5iE
4NTyJNPpCGetllzZwDaiDA2Sds88S6YeivHC/8AtweetC2XLADvlCZ86iRPW18DA
bOBV4xFtmtrlIN1sQV9yjW0doXZsdAx363cIgmn+PVI=
`protect END_PROTECTED
