`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TLzuxH5DtsBFNNZeTcrieCL4Xw1tT+dkxmDA79KP83DUIakQBdIDOKOi2qBshgd
HLiop8u0pKLnsTZRm7Mx1yRHBsXsKNwCKIgEXK3WiP0lsf6U8GDtpSZ+ZrnIFM0k
o2JPAthjreuCtwrjNhbK+zNIGjX4rXtMrd+NvXdj9eV+DKqrKyXl2khT3F9QILWS
Lp+8HLf1NcpXilbTqHQXLHWENMlCZY3jM+Nw3FgMVOcov0TDXWyXS/EOvGZvWMIv
as/HUU9KSBNLNFNjcFmgw8dXAuQ8rM0J8atQaCPWyOBC5A1olcUX7nLW1KsHc9UR
eApGPEAJJlYBVR1Z/vDgne+6/XlzrAwfPcTxEYjUFr8=
`protect END_PROTECTED
