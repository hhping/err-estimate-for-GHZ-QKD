`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tSJ/9r2ZYbEPvtOGP0VpqUSfm47N97DtzOt2ZI1SYYjlO1JSJ8PEG0jPP4ygzmul
8rEvB4IaiqbWvy/dE6kERtivq/v3LL3Ozc/Sf7MQV3hryvNZdoxSOvhkaxNxZiaZ
cjK3gLVtT+Zm/ui9v8vlSgS3nY27s3ntcOn49Sa9bkwCMwbvz+R8MuGptzXWmrNL
WPc0dSicvUec3F45ntBfa8dzS7DFnrbZh8jMwWlHaBabjofrJxN80u5h7uapWIRU
rBqNOAU1Fbsxxpd/I0qVmu9y9Br0DRXjo12ZNAr2rYdC+7xryl78AjmXq00jSiwe
S1wAry4eUSdCiUWDVhR439y9nVpz1ciJfS2Siby3zgrVdTY1wHnc/j1ukGGqslV6
BO/+ybY8BXIZ+xD8OYJWaJ5etgG2qWsjktnL9UayRCnKBqPZXLeyuTHK/InA7Zvh
zFu0RqMS6YlIoI9CR0cHRyMPriH9iruB6zaveLkykVr9Y08/0Domu3XWI4AAP4hf
9Qa+DkfrjAc1DmP4VtpP93SKAyn+PNNFsmYnK4FXceXcX+E4e4xodAUL8cX0H2H5
nC2HMzZtn2vhx4Zze/tBls3s4gjsUzsDwwKFtTGakK6M9j9KhnMLcBzAJpqG/lLY
vLsg4KdPIwnqfh5sMUDRdvrbSvrQrtLv6BGOaqlCDK2w6p/6nGxJjn0t7Dxe6/Qi
KL2KY1mMOsFfbSqeuEevlomEd3TRkrQ4s7ZG08axNejG4HZdajhDgklEZYX5ZiEO
+u3EugeB/PiaGX0r0Bv9ydECT+J348E0+QGuJqdAmu1xRtiWKKRQhKXb+qi8J7fD
wjABbR3VOMXoiepUl2/0oCpzD80Vx1t47sR2PSnvD7YWmAEIG3yIGV+2odMuyatk
rVQHKiChafeP10YH4OEuxbxv6Hs6kY2IU3N2G/9Hy6AaXSYINySA8N6gdjB2kG8R
SDhJ6knLMGb8u2d2kBCGMFDg5eKWy40DeHbplsf85mD3VsLKBGGmmHiSxLHypyPz
FXfAluQQYnbBkHoWZY+nNhoh26FxjfqkO4+DaPLQGAYaOJSI2AdEbZcP0xhMI1ke
dx2ge3SBriI3vOtRCXb2o4uQ8A8JMY3tYSv69Owd+uRPgs3MQTet/pliCXomuvWy
QfvbbOMA40w2MRe+SAPrLiliAj1tSL5msaQMBKaLYf8TZdxCN3lf1hKu1vpkSWWb
dm7had3cDaZc0ZeUEsyqqkxeVHx76SEHDb+YWEx/Z7V3E/eFOGWShIq3C65263IX
0ukeCX+ePGNyAR6goDvFNIB3rRV/ToAdg5LhpTFkH2qg37LL4IVx8rlWgTtScyJ7
88sw8nfKofopiUpciKOnqUlqQ0gDqZ2bCuc8AVLTWpRAIL5C85/kC5q77FBgyEcK
zmH33Xkcop4lwzXgzz13HG5X2wBTQfXUqIEvW9wndbIrb+Fjc2dYIUPeoTFAvEUF
iPtavOumpzHIzE2cBGQCl0TkNpEN6AedJdSrq2JsXY51dMh/fpqcLNzke9Zk6S4p
i8K+rZPxWkw3em63omYDpva4uZ9IOI+wJr2UdHdMp3LmPMmdSAqcqcn8uuP/00lC
GE980rh+FHGbQ96E9S4jqEHm7UBsglRJmbPzbp3iVr57PrdvDIboJE2XUljM5bCU
LLdI8G4lnI+UV9Naecb6OSMMOX4BsmkF9c9FTUTtPD9ADh2c0jzMysXvqjIaDzdF
Qh88KGAYtBMZFgEKgBf0436dz9NgB35dJURzCdANJM6Pp3Ansod0NHC75UuZvxKm
MbkfC9ENyh/Y3VFWHLRwZTrJmV1LeJRBNgEOi/DCVmO1hiCvE1FHTWYy5e5SljE6
Otde54e6QA94rKYkHWdy4KYGZnvfGuz85QMGQTr6YDDgmPD7ykn4rxYr08xkZjye
XCGrZvX5KLliBegMTcYFKnz749FBrD4NhiK+sWQhixYOM56gbbPDQfpVZKYHWyQ9
Q/kszzEnxRA7qI7QPORmPrjJSkg9yYXlWBoJN2Y7ACRm9YZAqXG3PXCUoCX+xULQ
vBMuuPiwFLKVW8eVLU02VKlHGH22VJMA15sqQaGieGKh7hZ+3zzK2+ir/BOT36hD
W8baTSZY5nW2AY4uFbT1bi9gCPJFt5aLsxeekEp41vHE2oSFL2zdRhqJq5Evvv/E
+Lk4CJIoJjd1XFRDeSEwWT84yvnXfg292ImuLuwjVOqenD6h4iQxog3vc0f3JFJX
gq/Khn9/wwiLjU81b5GhE/7yBG0Uvpmtru1GvbkuNTFirkCbyRqQ3M0BfLueSact
FzwBTrMI4P9gdEWYh75sj59SB1bZGf165TwfDAJlHk5wchtmHIFNEOisx3j9QJ3l
M6yifKpxJxw0RaDJtd/Esf2/Y4N1iwnyZ16IBo8j+X4TEYjdiciU9loeiB4ufzgH
zQuFLjb27Au3ACIgyad7hrbqHgEFCJfa7aX43WGbxmsy0w59efOzmsCBf4kQjlRl
QjOfgefsYlXoWpHAOE7facYIycYxrX0j9DM/Roi/W/S2OCVu2/JuyOJYWh/66lu1
hXqbhUsFZb2ajgduL4ZXtIJeei6ShoW4/0J4BMcWEprbi088vPsAK1sl03pyY4l9
T9+Se+/qxous25xA694zQgkr5d325bfGxzKY5B42ymN8ZikfiKw4WZxfV0aT47p6
QmkxHhhPaF9XSnSyB67D5w==
`protect END_PROTECTED
