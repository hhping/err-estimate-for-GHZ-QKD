`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zif4B/DaS319TQjLyD/V3KAIXlXujR4sGnu3fDTOqvTiOjaZIJlcYznGSxuiMezk
RiPOkwN3Uwtf2Le1rKbkOSD9iZ1XbXQ4peZda8CISea68aiRegxo3Te+4J6KQ4U8
u1eu2JB/cbo+1kBBaESqCQXUjBehzCczhB7XUCZsRDdBtQYiQorpimOUg8y36Wj7
3wwUrI+0+eUz68JROva/SGssXNHWdv0b+sVhz8Y7nMtlTlanPfjDV2H/pCSSKow2
8djXKMMz7IRqwjDHgfDKIjzmTfndcG9TU1wWp9060BF4w3x6hGHTnfv4xNXBWwZH
af/kvXYQ8JTeV5pjkNcJCNyKnVM8BJ5Tkl3lNUx9TWi5o/D2ODescYxsJlq2xxM+
cJTZXFkrFvvOhSgyaemFQ9otYdfl8OQ0c+gGwUdhqLGy4zDGDXQB0Yr+yjeyVb70
K/Gjlu0ithJXPP8ASfVFdjCnimO4PcY4PaxPP96gcUQ6yRpuz/2wqKNafH9XfrOd
eAW2wMR6vqs7mz7hjc538zof5Em0sgKML5OMWCu7O8cnsNYmpXIsSn73pS4vvvgs
YcPMS/VHUEtWlDvguQAS8V5kfngT5MbI6PmoFz442wZV2NQfPf9WrVPm9UjlldC/
dlbq74iuWydHqMGtupVj8GzscTFZtTXmck87Ml1eIalEh/alPpsUW6oi6ZcgEK15
j2q2mTTJ/xgXacI5hJeUfg==
`protect END_PROTECTED
