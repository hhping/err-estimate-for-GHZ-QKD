`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+d8kMljDMz5IiOorXKCmwngSw6mzRIg08obA7kDsaxI5sr9EGt4r99mBv8Vi3+p
CqMnrbgVcP6SaGIFQqrF6DtZt7+qZetawSKWTbnExHVCAUfiE/2QdH3T7hGMx7KB
yHmqy+StJ/3yb3D/2ozqeYpGqcwTt+9tLEN9e5lpRj8lgSMeFKB4r1tdwONHCe/W
Cwu+Bk1/518WyGxIAgXebrXIEv1ywNVspQpQrg10RNoCV5H819vVWywa3nkuCgR6
LK3PHisculGP3mQveLKriXnJjQKR4b/pSPkYjmFTy07O6f/xW6B5Y514fjNIv6MY
ZDmIZ5mDu6wSoPKcsoVa2jVvxv4vbf1PXCVV/c6UPMnztueHL4uhzW64lcHeLq0l
ekMH+P/Z7DR6LLxOoLIB4gdD6ql7FKtcg13qvQmwzCLjHus1KpzDQKV3ws4WqKQ2
/QnYElV5ffwjBu84It0u5BzU+bC24JQpPeskSytTN9f2pEilJbi9oJfxTEqntcos
u+GlpbYEZ8XbH/AWRoSBwDRP3cUc7srh7wYqs/qd9Gk7r4x8AHCY/tGp0sl8fID0
x0HbkrRP2jZ6aQ8fMSWJ+XVCSEPe0sGBum3x+WZjq0FYRAw8P0gWjtAxK5j6Pkjg
0YVPfYAueJMzK3++LjTvw9B4DwRsHJedDl1yGVI0cFBVjswJuPpor1SBtW5XfOVn
jtNccCJH0kFnyONFT8a8pSkHdfRcRmTkIxxLxlNYf8pBJ//DufTC8uWvtw17d4+a
F/HGOO6LAJtAOLyICl+L2dfOjiHB3SQ2jnOxlEF+hGNZA/wI+PjX07LqFM2IjIuH
Fh1xqCHZADdv1i0w9agNZ5Mn4I8SpUv9q8GUjDVTNjQT3ZTdWv0Qn2cIOIjkzm3q
KoXT8K4OE7J471J3a7bYDh4vjw+p3zDMG2U8tpWJph8hkzDLugCekGquIvQbA5P9
VPRaf26kKfROOj/+loG1x/VVZAlAfLtmDaJJGgTYjhzB16AVGiYBZ05oPv464aW/
ZZpbMPFwz48ICUpMpV2y7/pRzk4bMT9KjLbLQdMK02J8tbP4JHmLxYL7i2/4LRz6
2FqAK++X9bRWgz1g5TCwmo6wkK7FnrNvjMAkDcafN6v/6ZCF51vFnVlV/MIGFx0X
mPAse3/DY1dbZDv07xS7Q0BQKEWi2hP4DaxKOS4xCnnPpU0vtWG9SZvWQQGZqDk+
`protect END_PROTECTED
