`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2suwSCMbuUM+4p2DYnrY/ASPXLLWmobEKo2gmQ9KhQSrkbQ/44TVuHmJCERKOCu
52Wq6k9N6kqLWRJY3uo/PUAMNf/b1c70Yp+61AJvU0S+tKIzUC9R7pOs1ti/J32t
Xqr25LsjglYhIZahI7q/4yOKKsl6rPoxikC1BMYiGuGaLZKTNP39wiIWTMeIVclj
Tu0hy2OmebrgwIh0/x1vu9IXl/55T3O0HExFcoY6BEjcVX46ZBWtnx9ex3CValWE
pJ/2IZShId0SfohgEqcGE0Lu2MZMv3otNaBw7PdCw1gMzOEh/lbpliNdcYk7LqCz
h2EBcxzM//gHyfNNs/N6HdxcW+ptgSEjAzwuMNjbiTztq6mkAJ4IUrvOG3n8kTE+
pXX7rt/1LFvcn+DLkW+QJTZBCTKtPdbnnHJKwLkjQIq+TdmnoK5aRCpzu0vh9UTU
wUDbXoMQebN+ph9qAYWPmwz8PM85kfeodv6P+6ccpILZml+3D9jSAe9GlPECwNmV
4RkUJAL0rL0rOnKIA2LZYpnAmW1IeSbscfokpaxVmVU+vjdL/Q046yP5V7ts9siD
DTLMKhWwYCRyeAbMlenROMsZ4CyMjPPLVx0dnz++WPEQoWT3/BWDQUbuxDXOY/Pi
zS2TQqAX/T2pssrpmtQYCOzN1c4I/J+h8pK6SyGME0tS9hQI+JHgy3g63PHgEX8g
4EWq4K5VMheVT/eBqvZ9KpFV0wjQt+LwvCCQr9zDRk9kHjFmWYwIYztiZbstgrE6
s7VoBYhXbCJXlvnhNgzBnCXHvydR2dITgjW1T1NQz0ip/vo7ZppVaFLqXjd/zUgP
zw1D2ROVQzC1U/6e49GZ3ArA0vAI2GCVg+wKkGjbjvFE7LX/4372EZ0QKqgV7AWX
np9CjBOFUjOxhBhJZJj9VC4xfBnPzBwASp2C1X8mEMjxS6jMTOKGRK9Oum8I15ni
atfi/aGDwxIYGiV4ZQJ0v5Q3CiL4XQSEQCBewrCHjmAsIxHbLM4NDhju2GpIsMhc
BhSPPB2/7aH5/iajdelUd8aHnwPYcigBECRefyc0ScTEeQCS+EYTnCaElB63aQIr
IQ7lVDRT90TkFJT9FbQ2eJeinwFXlmNrVOLbUoFPwK0bXgJt85ShpaiI9lTqKAPL
QUgkOcxk705+MygK78gCONCFyLVgPA6QrJ3ttuLMbBxcZSEZhHhtdn7hexPKnf+u
QPq54lXSFqhwB28rBakFxpTgm69b20S+34lxQ3H9Qs/1a4eLy5r9Susv/LikQtCV
oNTIBeMTk2SqCF5/vii1ms+uSBplGd+wfZbHoJqH5fZ2Xp9oGclFpmfDfcGPXlJ1
`protect END_PROTECTED
