`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmIWsnI2u3V/AaoMnJ90SyAwhSbjIu2doe4UoM6Bn7RpmnCpQAdQfaHb1KHPhuU4
CMwFSghc9SYrysUFdhytKcgAzjpWsSB6mLd8zTtQ9pK8zT/VKWySeZRNbcMzDcf/
ieCvBin0GZzpDmidpSNnBLgn6pScQTkpJ0hjatc53JGm8mR7Xq2vCG5W25NmJbbe
o+FLmzTEmeWGtYkxiVJsAFYOnKTyevrc3/8To9HEN5De0YYjlob8SLro1iNB+Tdc
pVt6zDRezbQJkjlHwRimR8r8z1ey8SczW+JGqSEdPFYeD+oA1CnV1I9kT0jT5hxa
ZmPN3Lkgt7SAJwKLXWfmzpqAY9mbBbaanrB5w6cFxcdD+nXfIAHPJzUaW0K29P3m
bQKbL2Pfe6vE+2z4GmNut6ou75fCvnFui/Sk/8LmrAawTNtHMFU200SBBvAY4RHx
emuKszJLreMO5nBm57Oeaud/X9+kDIHRGYhOOJw4HpVCfScpgaBJS1z2sGxBxoa9
faI5OtUWA6bIGAkk4F7dyBlneutA21/dFP2Ke0QNQQoEkVB8WvnCJ8XXLlcXxSgl
ZVgh1ZdORR3MauIJtf+VR3gvqwqD9TkdLAP3ynZfPWxcqxYjhgYU9miHm4Hj7xyT
koRHLUnzcFh7d2VA9n6x9ikMSUzH1NJdTI20qFcn3jeg8eXDahPOgGZySbQkW8zw
rJkbaEA9khtpiX/itDcpBF+eniM7G+WbBVVjIb97FjlZd8P5++HhN7VhKxKSonkK
`protect END_PROTECTED
