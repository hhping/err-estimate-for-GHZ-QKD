`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ilq3sB/Lt/8H3V0g4E0t5DW5aWCY68Sw+FTP+kR+oNHQAI7CHbVldRT4KuOzmytP
Wga/OF7jzFc3ic3pcbxcmLfj/CNOHQEucxjkgSqt3ux6k2uKEL51ksyWnLcD91Jn
6jRGQHLnPqSEeUqxhu8W2A+IBnlUw5j1CQWnQnV0JuinT37I3R9bQsGAW1ajZyvl
QNo6eKltjeDGTh5TkAKAiSPY9SbbheGADP2s0wfC2LGw0LYY7yDfnrpct6BuqbLI
GrBDcUbyf32LBQgfnn/ltIh0o4WBuKenmS4vryFpOp6H4nVOUSaE0gPiW1cE6lMe
bB7NIfL3AZzoQvB6dvSFPTqKQmUKvANYFVAFY4K3WW6njLAcwFUAT9z1orSlOfDQ
LlrWHLf4z31lUXJ6rmH/4CkfClFgMQynf89YlLAoh9352u3kBGkcDw7C/ERN2SJZ
bZotrS/7cYMf4cKP2kbf+2cJ/tGoJu3qBpE6v7rJ2tzxA4SFu4+fISMGl13/fRmr
awcBpNKT3AxNT3Njaa5IpHvFn2QYWNVPP91hslDW5GvB84vii09unoymZ4v3JzLl
eCqJMqdI6oheMXmM6FRwPSExUPeYuWgPW8NbUri9WLQi9pmYdhLho5c32ryQ3fZ/
h6akhtP7mB5sCmEmUy7D/BEc5uRUbFP/q1Ub7wqcSlxzGESObMeWyUkgYkPXab4J
0hkKnkUI4cLbOOWq4RX8zZXJWPVPl0gFPeMGB1LdCU1nVIQOlwZgL0fm2nme9y0K
5tw7GiQf1K9/n0HC2s1a5wAI0lEGj6LOrmdLDx9NY56ZAGHeFlEe2gDOc9K8usdu
DPNRc5kE04fxAugAZlBTRlp8k7nXs3us33ZBuh5nJdT808+pnA2mIr9sdTT/OWst
gRnyROFH7PlWAGsCQ+t5KziDBhQAzQAhrvcdXy0Sm+uKA5bYOmnihkqu8A9ufc5X
TMuC1od6RN4vM2Yw/7oo/dbN37S4Yj2LOMucDwj2H9BUHr4jLsIVnPec0SbKEzep
YTdJLQfoHhhaAvePswcmeg==
`protect END_PROTECTED
