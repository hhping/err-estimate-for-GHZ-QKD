`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBAOmSu8y4JgMw4Pf6UU+VtD4hXf2lQZW88xgDjSKhq98TxfzChY2ojz/qQjnMFK
XFumWLmPm0An/IAs6TkATf1E5sZq+g7jYiJ/VFHiH9Qvc4/IR1nyh5jUaGoWbUIo
31woyAekqLUlU0GWvQBlwNqVuBg7mdmQHtJeark484l0SJJMb88aJcO6aAt/UCur
UcsHWMHBlPERZdVSYaOVs3NeI9u1RNt2lfsJYGYAHTUPrKU6ksBcgTOGTmKknDhs
xXxeLCqQvQ4+jKMjChy+rMJJgGuEpvAyhMr8ZskAahhMhKb6ZJwUz/t3y/ErInSo
HVnx4qhs9R+DpFY2kKf1ef0fPTaAKlNpNkzD8gdKidzNUFIYDCi4dGLu3lEzaYbL
NOY4u4pzdQ2ItYPsJGf14lHmNxLj7Niq01nQo9GRBMHW/0nB2BW1yWr+9v/IoKBv
kjXF83kTSZZvY4f8mnh4ou/jy3OVOXGiTDxFxfF97Kn+8jaHyzv3wvscIVG0idm3
k1uISfax5hLpNAD4Qb1pVdj7ur5IobhlqG9367pU2ehf+fEcp+OAlTjpL+FCStdt
UtAoPsfuIcI8WHNbpULd24iS6DBGqd2+oRjMlnUoaqGftn7rYRuWE6dFL1wflAja
DqCX2c/tMiX35xmC4KltxgJaLbgAgvBH965rd2R/cQf9hr2EFJXkOpgrck772bMS
GWVF2hHqSL/v3rgWdnAN3yUQpqBf1WKd07T2ynScUe3Lx+557gWWoZ8KvmEd5tls
bqp/QMuVW+fGyukmvU8DCb7pQacSnf63MCE2F/64CTaJvBCoQgye+Ruyzy4igybr
lQVW63KTm5GF7aREv0uPmydCiUbFv0Ffj1a6yIH5Htgbh9mNtYwF6CdxGvqlNUW+
aAQxqbzy4v7tJ/ba2182zzv7Le1XreVISaXzC6J/VUvu0qRD+CcCImRGeDk6Sr7M
32anc0y+apaepuKMwJ1s3KL+mZ3AbNVDktQqpOCLC7JU7kGEjdtMIUWe4k9IacdN
CAbxe17j6Q2pDmUybisjOBxEkWRpkEwqNKRSZXUcr6TvEYIyf7kUEkmBhf8ubv/v
fw1SObZpOae8AmSNo7G78f4R/mkNhsEHRDsyL7yyIxB/kYLajrmR2POzl+BOFDip
dtkc1gfxl9aLH8qrfn7RtvVpYUWOrbdHEK94uoVNGH5S3aXtci2ZymSoxljlosOl
C2XQBBtowUhaxLK70LIKilrLK886HpKRPZ/zeCproaMbSI0zLGPmyJDrhGUSHcff
+M672RB54alSq+jKs8xnjgKBZiOJ37Y2c3kywA+KSN8=
`protect END_PROTECTED
