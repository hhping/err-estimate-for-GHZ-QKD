`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qvRPXdccnUd9NxW+EX4KgMAVH3glZa10vTLR/iYwO7Td7N0SirVVGJP7Ag0kIzD
27aXQzYLJ8YrJpeeQA8rYnK+CHciV342ZgpenGIORamUIiPd6w0D7uoJrtqI0Iz6
O0YdzcUUfLqnzFOqN8YUBQJjdN1pZ90XB6nQmgvK7hQr0zaxdI1BSfxbmo+Si/PJ
8c8+Tdwt2pUc+Q6VzQ4LG4u8ndEUyLuxbWBneWfnsh1Qo36g1Y7BRApmI2/iTMsZ
MDDPzZeNKxDyNW1nniM7Xwr1oHWsWtF+Q1k6C2I895DO6SWMUctMXarFXJf4iVuN
eGa/RprFzNygSLZLVCdEN8lFeUxMjqrzyP9Wd2g+sNI9CZ03/sQmDAG6yuq4+g6E
kj5Jrj5BmsTkfxp0qNuftlhD9n2L47NC4i++Td2Q4GHpkE0FwqWXtIChtWvC4G/w
A7oL1wSolqe2yB/gj19ct9m5n3v0vnbc2lIFWi26rW8rgDrZCyBY7X9ypJswX3FH
sOQWxsvym0fwtT5KBvZtpeK/+dAIfZN2penURwXQGbrgzrYW3KXDsV4CsFXqn8q6
mickTIJqfUWZPPnSGv8ibyM9qe6FuQgmH0QdbZmf/wQ=
`protect END_PROTECTED
