`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6cyn8CQSokoUaGOMGW7OPwmEwd+ydwnXNylwQy23exCMx7sS+jpN9Mbl2H06OaV
ZKVdlIwyN0vsRRSU8aUMKlPKzYMAF83Vh1F+Fdu7jRXKcnn4U9MkooQRCtis0Rd7
xzTHD+37UHhhhvjbt57otFRYRwZ7Ly6+3Sot1o0A2yu97uskk96qlHiB758/7zkh
08jijBWA2VR5U3VzXjPo541MRBtQRnphSWfE7lGpCsSnAAOYUrpf1Bu/4DS/2GrC
1VjyQkguZ75YBR+zYbEcAT0m1wr6QwUNRmtn2Ex3gykku7/iFA4KyjdJknH3h7EN
bFfCcGMlXfpetw9QRAx1bXAaqqEeshy5gHnEkoGq24at1UOxxRLMXZrMb64aG2M7
Hiyx9Hki/nUnJBjZz0Wn4t/5nP5VPB+CgnwhXMfJWwBHD5kuk29lAP19Cc+C8aaA
2u83Ev6aRMVfO6rNHKRlQkBeAi67bzL+9nQI9ReaLPkubrDW1dvL4b0YuFB0rHlt
Y0ySzMB/bCuBitiQJQ+ajE9yncBBHaa0f2PnA/KrDkbyiU6stbgjMiGE/A/PVXQN
ghO0U9Zt2HE8a3MXTs9iieYesxIpTjuOQZWD2so8LcsHEP3uRktoMHwnVVyM7Rhr
P+ZM2rQwtx+Q/vtcAbkvBMX/PgHRVniMpec9NVr86Gco9CQi/arts01k49TAit40
nqTyi6PjhR2pWbpAfg5pNp+8UuaCqdRxPBB1wM1Wa9v/zRj1lzHjWRHJEBBYCpMY
Skv1T10yu6na/yEvuLsa5bT/I31lx/71cMLNgmIdom1pL/ESiAMkKBgHjoiFbSoa
zlCmBRrfDlsUg91AjE0u6IQvocQ4ul/UZaq65uo0QLqqQR0DWkvSR2YB3qk2QAQM
2oNt6wVpxWfLQuURRzdRMw==
`protect END_PROTECTED
