`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLCpU026jhBGgmls0NCPFZWqF8AYhvb6WQr0V17V1IgWlSgSjQyVYXV5Z2MtXZwn
RrEC02l0Hbhog9dJG0lyvPw2GpWuBiLgkiZH9ypA3i6Sc0WPrMiNh6s+IPvAgyTi
H+jLN3CC064/z0CUaD9eIbUlPcYK2QlBH0PHqVeu05Ao11WqB7NwBoOWYWM8nZNP
r+YIClVVhP5yJ6AOjWpuMJgd7hLKOz0umLuDq3sCX2NU3Yo7p3Z/PpBMb/grwrHD
OamuCRuBtr09P6WjrZPMiqqPt75zV3OeVZIATYaUVvo9rJV4bpbxldNXrpVh/Fse
5gIGgvI95pXNBO0l9ZwxOx6L/73S5RlVzRKeHMB47ki64sZrGi1AMtQrTizc23QR
xaNz/M5XlaLM2r61+N0BvziTEIl8VWGtIe/ZorTWYZHZ7aTUxQGppwvB4Y8AO26E
gCLES6RpTkQnE7QL6kf+5+Uflu5bvaJ969YhuQgpZnzsmmt+uearxlVjmxk560Y6
RFzmJi1OHkBfsaJdRaVDKevaj09OWNwXwr/Zf1a57TGaiUVEcMmhU7ivQffv8p4g
`protect END_PROTECTED
