`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PH8fYqwI0z6HQ2X0sxEaU0y/MRjB4xkrSbAmR2qmULRIKdysQVCvvEpSfhvQ/XvF
qV6YHg35SZn/kihHK8luYFZtath9tt2ajURBrpU5SnvEF4XmgBUZDe39LcilIhLR
WMTBxnBq/YjZ+IX95SWNm9QquZbexVm88/IARrMhpJiB5fUE5MhWOUNjAaziX8Jc
/70ByvuWuhlnWQxU798hvF1a5cKbMDtWsZY4vHBurMU0t/wdMu1CyT32xEGX8ZFE
84SScjhqjG58rNcybgspKdLbBn55ko+XqRQfTDb7/Mh8AtpoMGhzWflbXI+Sh3RT
LszWshi27/LBSGvrVHTorh8MWHBAO9x78Whfawd6I5UmlurkUDgBWbO5IGuSKkHG
tcr2vPShZDG8qCV2RAjjkkSe1akk7e/wzBJ01i33iDjht2noPsz1TjHa4iJzTdOe
jF+iEyW3fC9409PY0c1E6VJVbz0GMHE4UBJM0yUiFUVnvcClXP9bMj83WoRVlPPL
lGkp/m82BedbzNwXypmXY9M8psItiSasWofFxfv1gHQukYOO0joNuiPYgpP6+wws
vpcIVZ8fIR36Kvk6r320/vT6IESNV02NY/7x8N6q/jZCPS4xnKKTbS6d5ifGTJx8
WXminKiwxrajkcCQwG71JtDl+cb06otEYvQNIKmKVaXnqn9VhbjsH6KCDaOLcAZo
7aQkhq4oMs8sJPjiMIKZxxP1nnZALoxYv57dPXGOTbJgwcaD/DnKrTyeWof7aRug
eRzWcje1YZbWHFHx6ZnEdBxVNIju6gAb4+SldMw+rvCl2QUj1aq63u1aoJsgafZT
bQLqHQNgSsmzsjpoqJlQV7UjZSXsNLYqEMwJXc8IhAwEwUoLNk1miP93FsSS0JFE
y7QcSRa1yiVlk5jASBmOou9Ilm9HP4kKNvMgd9jXlI5T1GYsaD0v0vraAl5TVZrE
bL4Tr556wyYMi9qYKdbewlodi4ZZ3mYvzvSOhV2GAcEMzddGH2tL4Js+EPI9HOiW
FTHccBo9ePWIOhanqY7YG+iMdda0kzF2+RVJ7VocIi2mOD/TiZM9w188K6qUPgY2
nmvdz+CxbrtOtn/ociIQGwhj235jydEcGy8FDWKME02IQzChTNn/YDt46U06K0gc
1bz8mGjgaPdxyo22g94c5jVU07lCl9ei5wetFHiKZdjuSyUIiIGxwxwXghuxwz8d
8+HiFWeUNP4PAomZ8qZQridehX1tMd/M1xX90tG8Vf9aD8j0BuiCvp9H0CyhZ25U
y3OelPz/1hHT4OUNccra0GbMm1ylImH9yA33MLLgCVF5fQJXLhFryKWKvpNTJZQQ
fl8qUugEzccOla4BtLWSOBLhZGnMhlMjyjVxvbBgqHG4beclWWyy/oJ5glbCHsKy
zqOeZmkMLAXwlOt7MEXM2BMNySPKKbMlqtEcRTclD8rb0KMu72aH+JDs8wOk8TZk
x3HnNIDl6fXwJJrVu9DCfwf06eIOUjOP43u8Mo9wZoiWPbfDNYgIGn4ZZYHIbch6
dUf/MnAwE5OkB5Y7qs+f4QcDkNemrQxQGbAb7jSVu1VuFVTq4UNo881tXhfeb3EN
nerI7e0kCHeVDC1Vuc1jI8Pg0H6eIrFul9goVMhoVQF51djFS0hgGyzAWzRU6Tvp
spkaIztw4tMv6TI016DtNM7tvWxXgv82CS4q7OvYPSAqxlI3oNGlCeXjqPPmZLiB
ETc+Wc3EQBLE/Ybm3eW3XD1IZ9jDFEf0h9hxUtT9FGqZY9Xlaj6c0JBARmMyQ+V8
BjSwjXeqdyi3/E0DGJJV1gFrytNo0nFa9MTNGu00lv7HSjzYuAAp7xNX0mYuzAyK
Agezsjgf+x8zfoJ6TB3vn95QX5/267PtNwzzOWfOLDAt0k5/ZOVnajLYP6p6Vq9p
GtlQZHEL+TBTHtsCpeD4/o++0U434MipEgFbfjsfCpRRNb222d1cZULbwgUqiBP5
nYxRrZQY3+91IxaJ6FV4VmVYqkhWX/YQYtvErAlyJ6NOn3LeCZYAwMrvTX/DwkqC
EHRAqyXZJpAdtYYabVnAtqLqYYIxAdRFABHFfzOlVBI=
`protect END_PROTECTED
