`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQq1JP/XDOPGLj0p3d2f6UesJN9ayG9WW4U4u9vo2tarfPEMsXwu8tBnKXJIUjx0
BHaNQEiA/eFIzyuBG2v32b1giR5XHISAZRnyHa1Q4biHlylzwgJ87R5kjeq85vsa
EJbPmpP4EWcfqDaWrV+FzQxDmSPmaJ5pql+D/GPUl55okFwpLana5pRVNqhm1LY0
/BPAD1Qjd8T5PUnIg5XjwEi3HM/JToyt4iarV0yNxv1928UYYmpRc/0yaswhedbw
j1UtPaXmqetX4/gscWbeEqrkKg+WDlnqQ9n22K7/fhObinX90d++WWx6IP69HjXa
EjIWAX+5lgWAO7hL7uYsBtY0SWZlKujBm5tUZfGv5pq8CdN8R2Wc1Sn5g4bzO211
cT/cYmpL4AC7C/maYs4IiyCiBDQTcZaNLPnWpMidtlfLrMeB0a7lxRrPLNgcZ7rH
MPlygNy14YrkYfanV8l+fGRo4KlHN6aqtsQJ1afPt24+EqyKkvRIvi8mb0EMWQmu
bhjFiexBK+RTRM1TR/+2Va2k7LSXMYXax8r5iuA/SMKwGhfZnX4BtWWy7bDtPRlp
G5PKpSkaAWHRwJEmm2H5YKtN726HCkvvKtucAkZJvJH6DA5AoavVO+6jLMfg3dOs
wZChwcDtW2UldNpat9XK/vvubxuhDZwAP0tivGenRoe3XZlLIGlTpoGk25HJcVBi
j5BjXnVNffk3s5vFemMOkpSGB7ViIGRWRDPii9gnvxKG8opPouBF2CsOQp0KkifG
39e/k2Wjpqtp6JYDfweFbmWg3qOUd0kn1MZ54TDyID3CtJ+Awh0kC8vKvScl/r4s
pS+od/ZvACdFL8lp4CGjS1xaBXN7ptGb2ghAY8EcxZ0CogSv2YGvk+qKNwHWECqk
lySKikU2y15rmwuCJriGywuObWNgZk3avjKeNpQQVhLks14IKfLscWMvyMYsAf/A
W2bkqszV6SqrgjJrPFUQu4j61fsRkWw42XP5+mFbNWrJdeTZSqVudwFTVMe3tpC7
BedGllo8nqfupUifSh+F1yIpsrpi6CuhadAXF5eYj/ChWO9+bobqvitw2NNYLfJF
NIAJl0rY9irNAD6YaVAm4h+9da8DPZFswzRbvSQ3s2sBEvYf3lAg2Kis5m3DsyAS
+NM0OGSUFKD3lD4xHYSVMwLBTCvZYgGB2ekz3LPKZs7r8ReNpnE4J5Gg4toEfZIi
xs/wLQtf+DhjSy2wO6Nq8uOUuiJZ8wIKiQNbiI0npkPiukdjzFwJoFM/BNTVjjSL
PSPNFJi9K3XcY2APSdypQFkSuAiS2UY0w4TCiRMu3OScr6jlm45w8Ctj+fgNE0Ft
SIdm7JQWctS4qdFps+VDu+to+l2X7OzflBD+EoKryZpXmX4wkZGxpejpIn5dFsXo
b+PROMDI40DYqMIThLOfjDWsXGttLZz7Q9z4FezBVrqxV3lxS8nqpv0qB8SVI+r0
NX37tfflIml6MnQg8Gknbvx4TMyLyZjSkffLtgxxVORAKYtJxdlArPOBwR9FJJHp
p9YMkRF/+lqh2U3HvGXSJBfVMLt83KWCvIFTDnHI4y42cB6z2v3g0upfGAsQrsiV
Whi2qy58JuYaCzeoSIUYoq09P0IexIyYBY/lUtuK0mWE33SAnv3LibUGaip1ZrFW
a4yTsQLppwRmMAOMcI5z+wiFVXrYXlqsSv1hIW6x8XJH70nCjALwJITiLiEEObn+
bNiGZieWAgHAzqX4MhLrKOqjPL0El7dmb6KU2o/zsGJkzRLwGkN7Zxozm3gQ9/Q7
e52ahJNXXgtKc5B01sTEI5PyO94yK/TDGdrEB5LHUYk=
`protect END_PROTECTED
