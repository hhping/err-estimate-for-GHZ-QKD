`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3F54w2ocOqzOP01GzwNusIi+7HmTK/iIa3qk3rJfLBG3cwAEymlUpS4tcAX1U7Q
yP3NRXWfaivswr5XCTnX96NhkwoBc0ZN4i+RISux2GdrXTj5vv2XKOHjsGtTqRLl
S+kRHREJ6oNqeS5tLONnx8454jt7OUEff8pbgC5/1r7XVuQx6q9+ey3uav35y9MB
bXtfyNuRj08FBeDh87+dq8CQW2HWqBSEJ642vAViRM4+GjF2mkPtAjbVNOHanrjq
XeiMHE0fVUI/b5SHqSHuJ43jEbf25uQ4Ga8be1MPSo3BN0yvH97JWAHXZua1nxgB
DcmGfp3XSZjgpZL4NUjNnd0Z5cLMS/g7d1eAt8SEpkVeXEtPIVzMoQo7Fy6LkyG+
mIve8FWzPsBYdr0shuJnyqbV/PLZShMzVlJl7CLyj8Idl5eIBgW9hj4Yh1aC/JYd
1S3w6wfrfCmcivJBMN7KbyAQzpAfcZ/Qii5LE2co+rI=
`protect END_PROTECTED
