`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FfdNK09YUkZNmwJXLiezsxG8PpM8J5hvKLT2AwVNDrWWo4b4YlmSA0V5GIfoj+b
q9JD34F9aiXkcy1mQWIXybMOK/6469eGYxS8zxZ4lSa8pEiSzldMYp66NoqnPPte
6NbOfrOFyyqNOcoDFsRVWYiKoICAMoCNZLUdyW/sKnMyg36mPWfaRZOvkiW3dVPa
dbU69Yo6lss1meJNXdXnkRkEyoTg5XM/p+q7zLvnszj0upa6ZyF6ME293xS9TE/i
Kuq32ZS6yEAi0At+jNI7nSSvdGF/3B3CYOpz0RiYG8mjYtDfOooj8NTVYle8u9aR
HuudCKv3xTRNTqLQCI/hKhAalDJH8SFRhVS57L0QeSqlG2QPdgCH55SFKWRNWCXb
CYMMZtccl+aZihmhyy0bjOH5wpthyCqB7Lz42ogNNoU=
`protect END_PROTECTED
