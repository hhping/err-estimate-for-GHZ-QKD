`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfzVVA4fRN8F9dNLi8CAF57gLQZiphldGwfeNyKG2TZ91AC+F68QuALztvdZfsOA
P2pVZbt2pXPoXA+H52H1DWSyzb4TXBqibFhu2t940z3bHVp7pQnZ77N/k7q+MS1L
F3troE+iCCj5eWIzYf31roi/N0dEPtrpOkHAm45GVZ/urTEYg+UMQ3Bg3//c81k/
d2/APqGm1KeyFva4QEjmM3ak4HoXRK2YbR7/a2lLMo4NWPz2psdvzuVk7WFx5pJI
cDdZ6LrkpKgkN8V2e2MvQsSx7gmYgBDg7MksGaIErHBOWECcnuQdg/kYJX8XxEUQ
UaVnZXfJ0iALII0yZBT9TtyScQDlddOfnFeH+XmD6D6ghvmWR6A3tUiXtxUVLYoZ
h/XMmGp1fAEEw8Jva6W3/Cf/Wb2HPSR8NFSQXjDd1nuoz6KwE5tRa73zXPfMNNgn
i79TKmAilxnGS+RvXlRjtrqJSLwKETgxJyHMdY87I96FhEAcSPLS9SGLukrl04Tz
AR2T8rL2wns2BJAo+robQz6XHMBhaxgLz41OZKgZulfB1JQHCcwK9UCjvB483FRh
yh2EPtGHNsUqow2ux2XTrA7uelPHLeV+AgGdz4Ns9fm+5Fo1xpw8wHfeLS9ZOOdB
ifivujtMHNc/XT48oRpXj7ytsMozYC3JbOVuK30L1KWzDGIIA54jV0il4RFfgJDq
4C8W9By4wNefIGKecDquoSDAlDELiN8GmxU2WBa7nIPOlKqbk6M1WSUU11ZbVTDf
Nju0PutQe83W0K5yhrIYE024z7aSBwohkv6eiLKgkuy5IXHCoq55DHizvshdXf3C
TaVBWGe6lDwBj4w88SP4RC9boZw7hFEPBiLPcdYq2DDfsDsTzB1QwTNRLEr4htez
C7n9VsU81LZt3JXGROLloGani+sUq364YBQw3C9Fv3SI8ylMBK6OpV2vFRHv0e82
k24u8ZQjNCgn3C2RWWNvv8ZXx0a+M/GmliSNoRsBJ+Zk2c3zjPmf8eP0WUKZ0PZG
MEtN6oXs6vYvaRI1z09yD866Lr6iaBP+GrCAmg73XK7hSI8jVl/7NQMELy5oD6xE
gQRWvbj4E/xfEsS5oRceq7/CpcKHqLKqZSmRNSV6xjtFG0x8i7xbXdcIYOqmoQkT
MnaRon+gFb7Qw4Mb/2y25i+NabxQWuCXuBqpAn7k/YmDx4Xh93Fv2XASSjbogckx
3YwX6GSMdBD0UODHR+5CPAwFNMu3nYzANfXDFDjOgsqq9Fs6hl0XPiSfv0X6FegP
/0zdNg0VPi4pamYjxS/fK0iDFJME8GftG6aNqJYD0U4wOLGoqFONDyp1OfUt5Rv3
ABDZJIK+jZ6CVdcLibJylUDJKYkiArpNojsCW3pRarJb2RGxvJevyjbcjlxzw7yQ
kJtkrrT5m69OaA2Vx2IiatuzjoHQUuugcqIPDBjJvANSy0/q6mLuzmS5uLIGL0bI
RO+ocULY85T1La4Rxkgr3iTcBKooGbRJmCxZm3TKZnfv/BBbfaEGWlZJSjy7iRiz
/7ov7K5ZBDKfhsgE4oXzAIxtrhe9ZHcocV5dPij264GBndmCvDm/mWFSaiOxJkRP
M/zEbzgqSaAtlgb41ZnJjo4HIKvF/BKnfTGnH8SHatKrr0ZNQK9It5Boxc/iwvtl
4Wy+lqjvQnYrHVfHHSKxgrWFdYxbdWkiMl84y3myqOkL4aUQHP1p/aF8RWBFmkCr
AnRaUgXnieEkl/MNiKyRMbkPdDWu57qTMDX6WPNRYmQRW3gRJjcPoDy+UyEgZ633
XAN0I16G6lvp7oQJyNJOdrb8j7dZZC7FVK3oi7dZ/a4HoibPvMEP8k8WgIsWz2uf
M9WY9jJPLfyw59QxZzayfN2yxFIbxafFP/kmpIHi3qqBUSQ/D1eglNUi49PccIDh
AAwOJHzNw4E/Crrzb4FmstAmnDGvca11E7MrbHGOUza1Z/zPO1/oV7Bkgn5OODzW
FI88HvV7eLNkuPs6zV5QwWDvBXriU3zDQOQBdR8YaQ6fkChjXuAXwcAH1vVCzxBG
sLHH51cBLgTsn2W0lws7YqDJwusa5FoQVMJVv6fOPXKUh6NYKrcAw/Lom6o6Wbfp
aMZUd6fG+SmZfMjcN1sM+S5NsQ+EwEl2IPgHkPIrtoghX+O9bQYLUUIjK7GXw8tb
FBsggqM3wv0DteAc8v0qQwUh4E3RzMQ8lTrSuL1CQSndbeHFp2RiBDrD/zZr2EIU
CRSSjuBu20jFXwPJc7/0FPwOVlOUWzf+8KmF98iSg3qLwsNGP1kajwcCPoOO3lsf
WPY6mb/urMaCdVwYTuGjV9/X1zbqCRkYGoTOP5967F4n2SUl4LltltiqBbLkakl3
DaUOOkP7Tq4vYjarakhjmYbiIXQNxcLu9YYIshQNouUn5/s8iMQWBi0j8SYo7lk7
1R84hfAwbEiWcHPEE1BGTOF7esotAjTOc2nX75vhqBe9Gkv71Mofj7e5mW9p/mun
NfjYF8asKN4ZLkRGGr3CND+STHCJO0Xnh75nDSdvWpc8uV5K04XyEn9fTUSB/hAt
cohwmKf4aWdFOlJZjvfRxGoIrTqhYQ8wScokWpFM7/n4TMGVI6WLSVqP9kwX7+V3
9carroEh3zh2kaJRKkDMxX1i48z0kllfAszOhK9TSKejZbm3ScJ1bfWWAlpwuYU6
w0pW3mnn5zGWo3E6DLvznpb7ahPkwvhPvntxY50WDSFYi1MpKKLqKg8f0XeDkMsX
svVik+Cy4CmBl+g4lQz9MJutw4fvRyrbMk20SNDBHF7eAkUdPD5cL8ti6s+5HccP
1TVTOIqOoMrqux18x1usfll45OIJ+dKTGICSvBSqeKjgQItvUWkxK5TBltYKXNfc
5iGVXDhILbo3CY9NRBAvAVirKu8JNq/oKgS0WJoEOTPMFfvqB25/0KJ8ZVd+R+Wo
51Q40HIhkmfKKLJHB9g3BnpmMwooCfcf8M4uimOK+ucDdBrASr+xkf4fxFcviZrm
epvWvrN9gkCgLTrXlwz5Eq6+tYEp3/in9oRxJ067ZQuNZgqUfkGZMFlnVaPF+TZP
2D14SS+0L8T8Brf5JLzHcf6IqtnQUL1HnTV00wXk4HRY7IhaKMfSmd4Vk+C5J+j8
Hrk2Y4Wzu0/AJ6599qw/sufYSPKlxU1w7bA8OmgU0FMZ6pqND0ReFduu91yXeDd4
IqL1ubV8GZ2FxCyUKkGDnizl/mNI+Ej90Cat2Wr+I+jSr/GwT/uvYWVc4XzgfaQ0
JWw4T8fy9DCzB98H62QqzB5lQkK5d7nyST64h9vVPX14wrJZ/DaCkrHqi0tPisQN
ORUlxwX9flSVgn6s8vjS3UqvhzVZEUc3ksIF2Q8tBb9S1REhfCY3dGu+OIgRsz80
/fzLZB0wf+DQeMpZIOVBOcz5pHCusA2r97BWoH8tCdysSaKlUMy1g4NnMeiPZtHd
bLJqBkn/x6YDfZBPEHuZFEKagdWQva1F9FTLw4yug/vdHz3/YGIqbjHuuV0J3G2e
SSxQ8XMm9q4ODYEv6c1sBBXwcz+6/Fq3kBBSSBtC/T3QEbC7kiBEu+MFkYRp4ZuR
sINvSvv4fzxEdzU5yTE2DFm5+0Ni4gmbjjNclqPMSNIweOqKU5R+CfBUrX03tJzC
kJakIo4zjIxnPtEcC8d7EoXTjlDbR8W2TeYrdwSADCkRXwC+iqZuVmAxlGvkHSW5
VEAqmEwU9WUUs3OuQAXs06oFXwkC/8T5Fzq/fF5NLiD+bB8tDHdSeKWGPv09O/yb
6V7erOkmTPByvsRSIJrkE/LacKnApPY9wTybxrNVkhUlBJEBj+aJZKMqBYIFeuRb
wgpuUzdRu40RHGfZYF2ycghRiAi3Gw6BLcgJ97dhGawvineFJrjkhAmcUxHIZxNI
eZR2g5qIYxlgHm2V/Tnl2y5oS00peY51hNBmJisClu/UDL5SCJQBAyXTVy3a7vW1
dtvzN1dIY8PHtiBTnIWpX5RbP3O197nFhhWNWVS8+JqNG4I92A1bKLVVq3CTpXpz
GR5CJ1ZKkRsjZVKRdc91HPiTt7nvlhUdx/4IhANSlLbhsAeWuIAaKO81JWJp1ee4
nfprKjUVT4rP8hBLCN4tskJK4e6RU7gyc0vqYRGRo86dn2Jd3Fwsl+AY7V4GQvyX
IlDwiBf7P4vm24hzBhTAoo8pUhrF4G8p4zhe1+2It5dCbKADzGzsV41ljewv93bW
XtPedLeJ+vqKRVFcKHgThghWnWBEJAYh57mcp1EWDSnNmr9DKtSnj0219kEOzIDg
V6cbRD+WvOffalPNaME+yfDG6d+huneAKxiN3vY24lU2XczkSwv3V8S5954ZQFQO
VwdrsoVyKtcWtex83GAXHwnr2C6Sg3i9aahvgoK6llODV8XbpzvvkNKCGsY05pzQ
kk49+Xx1dKs7n06wWvyIuZqwPSo/KAFbNPjYkLhnZA/V2KKylQiPJRWCvSy1sK4+
BW3uzfoDilr/npgJqst2iY0kYQxoNJKsAivNnUSCwr2vzcgQK9LalwbR9nIw0bex
jnPeXetTwSayllESdzqbECnFncEo0MNzHY6pEqFgEHWpMNkqftcTgE5LGGBOwpsJ
Ytvz2jDcaPqtK+qQRz9Oiyigmo0mKlCQ4yYyG9+Qxbno9cAh9M242IKw96m5NQbR
JXkF+9rwndg01fec9TZif+FgR4RAWhmJZXMOsO2GO8nmeKRZuTUL0HIbzHInDN+X
346QSqwrHyX9ol5vH2DJXFYK/qEFUmSVXZlBL3Q/yRbaNrgN1OIAwunAbZBFCLKs
xFxIBYWdFh5RhLeYu92U/DgiINBTLTY0y9/GtrpTKkN6tZGaY3Yl/hoDAqwXJ0ne
PTWJDy/ljPlePOCmng8krsPrZ3kz7sKQUZytlqlzc1DBmuGpn9W2CdnxptvgyeZk
7fZkYQ58+3WI2iWGLqpIIHWkGya6vhNVaIvXL3+X+tG2ao7/yAY7L+etCv8E6g1V
WIzr3m2R5mplN5yzB0zIYnolyvk+CPAHe6Sf8rXWRz0E4iV3hHQFejVwYgqImcvb
Wpl1VfvLg7PGXBVC9hQXG4+I7Xy8s2CU29WI+sXiPl7aNdmo3m+Ywir5FE5n93D8
htDhWpPXgGJhbUxmDm78Q/oYthr/UGhPKVREMC6+PK0Sx/Yj3qhaBT8V0Vhk/o8I
fbMEDwpPW1YoGDTxoFDB1oNyCvme1hYznLPU4Y89BKYUqIJQ+QrPKoRBgff2f+Qe
mQzgmSyePXYyzCTOq42HKFLmPK4xIvmnZl9IfmmYigfz1gSnDPvKVhfUQS1cOh+t
YAiCOEh5sAKtiBz2vyu5c9gAqhClYEWIqFat59aw8mHSzLJW+6sffA/YQrDMuCye
VEYdUUDwDk6G+QBeYGejOb3LCFU3WQLOvrjGaGI1EBgbMxeSnwW1Csc7Pi00RZtg
nRZkmkS7w5MgBo3we222De50KymkNAQ2ZKYUKVUskZM4Psb1Z83UDW5fu8l8Egmm
FLULrXJ9p+CK4QUYjIM6DBampC1sxB7WoRsxyC9+2MA7l2WujHNvxGusJSrpJ9Jw
QS6IefsOUkZWUeY8yY3cSfhCoq8HvqeYobdCbTWKRZ2pzORpgNjbBMj5A9YTSMZA
/sBiCMG7bdJdGJMKhm2YL5oIByCh/No1YrQ9PBDCgMREV/1RZx9i2KYbOgYT9e75
0DhpghDQ0dOiD7eQv9S+SaceNClgEXBxrHdelP4u/0JJzFIpEKxhG/0h/BSymDzK
0jUhUj5mVBDCgopBJS27QZsrN00ZfF+57jgr+yNGSenxrJUBHMXo3hLtX1OXANbG
0b2b9AIW2PPVsHJV1b2IyKJKGdU1YeQT2yafYKb/jtwt2oohQ8TMlki38xi+WGKt
If7TReYwrZqXGjoBQ8cZBqy1R4oZwL9cj78BQydITCoBGtIsAmHKao3imVX/aXSS
ey1jT1fbKP0ycmFZ/UjEAeexW48maKRbgcYhjKhTEr8/3er0aDctBHuiM/DPDsAG
QP5BBI/15iKIxGIgt5XZclMYgdQcQq50SRmirw0BEbgSvksYY0q0ys/dsISSenaa
Dz5qx6lF22LzSPaJ8UrvExOxleqcYWBZtAbBdb8lf/+KQf6NKSyDD9DD82vjU/IK
qEZ8N5Y/ZnM6+oonHqHxAFIRbe0mhZHQlyqVY76zF1nRDIwwWNIxTGCc1g9SU6QS
raufzMxMxBkWg1bSIBvOGt/qoN9IDqyjk1XGtfMre8alHEpn4vMlaVfGKl52FzKq
J2Cm3lAI1pY1dENwnglSAMUxf7ZItet4JDdc0pkCXz49fTOAjjDctBPqXag27Z24
zqMe0wNP3gwmRxpvH6qSlAgcKHSQiS0+8AHAdFLbvUHOOqjidW8kmW6c2e1YMyJ6
hcFFNRq5HYSZAGbp+9BHFZ3BPBcw7pvIpU7pt3+kCLcwdu9Xr6Z1BNA4bwEf0NGx
Imyjm847lFw1l7x3+sxFE6Q+Pd5RBccULEi4nLS7/ABuE9VJh7PB2fs9oen6vWqB
5mwVpuU+nkQ+cSUzeaHlZ7av7ItHhzoArCk0cQ4QKDOrMt9egQlM7Ru038/L+snP
T7eZjc5J5qP77lzyC8rYMrx4oqyFlNA36Y7r13mHUumomNNlS9GV7fgClspJ4b6o
gfBmgdeD63D4ZnplFvHNwwzPQ61IomLbN2Pvd05ClV6n6YLy5dDxRInt9ZMz+pDe
NFV0Ao/0U/9IWxoUiH8lHwu2WU6ppWvB2ee8PBB1yte43cqnEScabJ03Rx0hCNEz
U6ziXpYC+5qF+zADBLEpPZi1Memu1T+TjuVnA9dY4CxDjK0PuasrdrE6zCJRhK1K
5t4rgAJ9dBNPkpSI9wFmKoD/zpLTIxllzP9j2PUpv+3O5m8EK7CahEX/oseMJsiJ
7RgpKIBKd71C4Oh1wuBsDjtnBAJ0K9wnFdY1KCYYU0jjjKkBH5rmJALoZVRdgdQG
k0tXR9Jt0BNW2jFyq280CePkg4VzXpaVF9rVMc1t8mqVg5OFAGiy4ZKtuSAE+Abh
QVC6xpCHMtuXq6KTA+k4y+a3aWUOnF4jdqu3oleW2VEbA1rZ1aKw/hTQ+DomBFqz
7xMvS94TCGoF+3vYWIjyDus9mPzeXmtnk+1qDkYYfulYJQJwcfBcehgDSBXOvZb4
/vlNxku2hIXgZcOLEoQSOAd9dQ+YHBcBoevo0SqgfTmCA0KNJLqvUd1jr8WiMj4T
zE1YIFJtp79Et65KVVnOKcT99daD3k1XufTUmOj1Pks6OizWbUpnifwS4iKn0rue
cGWdjL5i6hx5G4IKr7+r/vAFrnqCEOkaROWSoEVS7k6ziJz3T6M5SWOJFJf8N4cT
bwdgeVL2c6WroQqWhDtDPtrHzQ+yuCjRS4FgC+tRCfDuno3i3rTcJKGJBpvx+Nw6
sC9Io7kME0sMTmDKDIXNJn46eRFzUP9B31zR5uq8XtJJ3qgiJpayRwZB/xrq3FiI
Sq1G5pOBxm6TVLxVQ+oh2kC11ffnfPE9KaTp/JBscQ0ihW5UtptiNtUsqjQLDfPA
oEUZmOIL+KXNnVitt5PpYZm1n8A2Swzk2nieUjZiiX8RiCHoGV9qRl1S8OdnqVrn
dBU4Pa4N0sRhMb6S2HfglIIe8cjUSVICYhdtsFnt2c0Vh2rQATSuybU93I3CwySp
h3A6WQG6ECg3TYo06ydMgWgmS0ZabG9zxDjh9uy+Y3J83eAi43pJySVcczEGShsm
j034lVrmZNRWTGFvRO3TreXi/Mr4DQipgnxSn0dWCLG5JRn/L74TGSDLUka2lCgo
zBiXQxbAt98sqXLC8fju/UvRYX9ylmj8r0rWY3sj5GO+/QkiqJeQp0jHcxWKKowA
+B3fUydTc2vriFca65TjVPAUYlC2ngR4GnvMvjAXW0jo8QJh+GzMnLXJzSzJryP/
1CBL8950ym7m2hGYgxn0tDU3sfXd8H31oNI+ZKSWXuZ1Wz5Z/wn3hDIemvu99FGV
3sg1CFy8+eTBTkEi4bx11GVwLhvBgNpxVrUa9s/mShr0v/n6FRRD38ZkBVc60Pgt
KV0RUVDoGbUpeHCZT7GAVSnvdvG+XfaUEuY/+LvK5/VjI37rylkBFwmOhUZ5f0/h
KM1woKYXjo+79QSk18rDpK6Q78NcQpx2eIPngdpL/DjV1fxbVqClxn+mR3ZJrSnm
I+O3zn2ekCL7N0WqDWSVp+TAi+rkmh1xsbPaGlbNydpiO+rQIf+uLSC96/hvRr6Q
pOvH7xxlTAy71HG9VrEDKnE/dHXSNi1y7wmbWBIA8zsopRIXJjUXsQ+DcruAk1y8
BmUw2MMIigKk4S7Vxpm5pviysl6zGKl/VDgrpCrnjR37LITI0ZW3MpGUrDiutoaZ
7pcHo3+hYwg6ngI96jBWo2wFLkHfPWXXwuAmcEjzKrzYSl0ioa2hNAp/dnBLasod
kam1s2etRsHAeD0vNX6MziFobH3NGJKwLnmxkXv7GUz/MZM2MQrS3Ng8OfsqRfB5
fbBlZCFdOa4XnI4JWOne+ZdIYvN/tENf2A/BzeIFDbj23a7q/STKDdkL1ZrZe0SJ
ml3KjmzxBaS7jgeIv3zPpSwHHvMwh4xAyARxZWbi9wsPr0RU6Ryh8nmKaIOylfjr
aG23fx3BQTHRrHVcAJfjEKYC5hDl2K8XyOP1VHQoJrJBM32skBLUUMlOMjQKoLwa
2sIZ5DQEKwOBfaXgfMOjGxHAoHBIohejEm2bUoyQewJJOaAQbC9+sShhGylaEE14
qtpb4RYGFDkEJ7ORbG6hcqhxtAx/W3p97YGLVrfij4PgGLJ/uQlXd5Ej0/85O+KZ
d4fXJclMIn+jWOEptMtF5QAPhAeC+4iE+f0O3qK5jJ0E7BfwYp1X9JcmFZa8Pk3X
bSNhwKI3gpO8+ahUSg+KawGwB1URP5QqvQx4CPegXOIYWN0s+yj+K3rW2TUwRTdF
Bi7qgpKqgu7gfa57lG6oLuePm/4h7cdZxfoeAyGnNeJKnxCPEkCMv3qiiIST8Vxy
FwhrdX4TghbGqvw3bttC2hCZYJZCdL1M8TkisGllJKWIC+amPB3kr1yqsvzXRZTS
RmRwUK9OIXn9F7Of7Jf6pFcKzGRrzsyv1D4SjPFkWBPka/EA+cdEAogZvAGIguND
Pm+Ud+log1AhMw1yrZwUbJ6WWRPzQhTYaKpzMrvqgajWQfOC3pjtON04M1kQvap3
pFuYhCmR3SC4fXfPzyHt7GTwkEN8PfX1CJ2p2A4bOLMX3UFRDxDOa2/RjiDKgfYX
xnYzyUjvb0aevzagTw9eIIzYdCVp/io7c0HfajrPhi9ruw+QNjOGfJ/ikrLOHjWy
V8OKU5Y5suJ52TcHxqUt23LtGGhO9MoWmEa+7M+eANilUZpH0Mh654CPX6k0NQAw
RIvlmaINgRGg4ZYsJq0lgaZE4G0CuNKKeya3a8A30IdijU3sUQqXe8hxjvcTYW80
M3wbYjnPthNsGodSAGCTidpn4bhmKekzIcZIr/PB8a/Y2la5ssfwEsEoRq7RNK5H
/5Xa71u34GyS3M4UGkN4G+KuyvuLcDFy0Ln1bvRUCtBbNXiP8YdkvzfHszz5Uc6l
vqfRm63W8xhHwBLzAPTnyy5aDktcWjuBQZsLrxIiG/LcYWRvMCLoyLMoxtJ5jkW8
PhpRtmp6LsGsWJ4aT6yjV9+6WGq8B6jOiSjZCLuVSHyISsKsmUFb3YMxX9vGOfiI
Vl6gd0oUJIytUTnOiW24hX1rQW1OINBtVDXEio74CYVkazuvr7QcAU9XMfaSCijl
aqr5e7sLPRwvJ4Zvv6Acv5ePYxv+kOO1nm3H66UV2M+Q8iD2OuwD0OLkep9w93oi
nS7xbxGYuY/lkO4b2WSH6GWhMebq0Za8AaIe7k4vhxHoZC0sz8zpaX8ZaKoxOOVl
piN8rjfy5t0iv3wbMtWFEzjsMgSabGJfd7EBXSGbxiZ/QMBsC1eC+OgEShRu+702
aGEDWSiP6hKI35UlPxHP/EJpzhiYhjfCP+BGmUPNpphLnnY/k6rvArfwwRUVtVKi
zpzeUQ2wLByxrni2pNN2ApYpLMzPE31017U7yHTNueazsrNAqPBW6XXni0QzMm/4
B1NVThA7st9hZ7NpjOyOWjtDNDzqMw78cAyys3IMFnb6BSKc4eotfkXwEt/I5Vmo
zaQNS0qvGkU9M/ti6KDp5BgVi5SsqAgZFMT0CRawjj95RmxPwAvR1yzRfgUrhiHN
uyxGMq9pon1CPjWqXEjdPOKdWSQB3f9PN+7Qu4haUEckoIH8BfULraG+fS7HrhNu
ymXtAQMyG1WPbTTja2Bflu/MeoJe3/CyB2VzIV4o8BAl1i+v7KzqvFji+Jze+Pwf
2xTq9RPldXaMoL87tx3oKhcS/R+/thfVWLkg1l4KuTeQBWMeHyXUhUxIhUhv6jEk
P+KTSzAGex9NVKfyddzolasfRvur99xSI3lBw3kxHOeftwUno3MBWiGGnzgodn3y
3xVAC6VZ6y11r1GtFJnKBTcbkjuoOAZNseI4oXq+OSclU9bldIuB4+GgvUJhcHlk
YXTkzHXq33BZz6ChsLUIDloby4KiB9LDiyvEZzHGe2BI7w6LzpGZSbzor/zmC+FZ
ojCkxjPWdl1DoimWfVaR1fcGRNVOLVkuCMU6ot/QCuPSJ1guhNO7Kx5znpJbPGCX
E4IkRxEQfkVPsNqComW0TB+HgM2x1VEHJYTbYAKnqLQZghZyj7SAu5ijqnUoIPlt
AgIEQcYVAe0Ncnl9xxbUe4SqV1Atx90Y/mYOXAKxejTe4oziO/pThSIVp0a470rf
5Xb1KDx2KXzyCvRCA42qpYn76rlKbiPN/o4bMMo5lGF18c6mJEqbLytab4FRlUwt
qvu8IzXBYk/vw6S9HetBPdzxQpJmmCGZgxmx9G+02xAqkuSUWWdIBRIONhiMNYEa
IjmB/gH12q7D8SXsz8/M2eRb4ocXxyp2TLgrKkTbuiWwgP8W411r0tNod7mtbSr1
xduVlYgtV3ZBmdmff+GQHlr3MMnDX2yGEXVuYLaoHL1JsFP2TwLHyKAJ+RAVOxma
spu0Tv5Q1kA/kFvw1zvCIpTyzEH3kMDFwnoGhoQvqq48fv+4gTWKxFoPcMgl2bek
m845J6qft/kgqIu5N7A0PXfltOAw6ljtncHvNPMiEpNw3/L7whi6T+qeavqnbK8w
A1NqEKVWHCJeNU34dm4t9hEfEDToKAIuZuneLLRgMJsb5tAcu07Sg9+xyjPi1AKP
4ySH6+pJNqSzSj713HYy3sGpG9XDVxCZkvR5YYA8b5h4j6ki8iR7CHikRzxInqPs
T24NUJpUPSY/LVYx3/5OAd9/qN692QAqyCGuGqmMBLFzZYJbXe1YkTPOZQM8233J
NTpFUWqB9xIQGq/ANEETzeCgKSTFWgtKrn88x9ya5MAPP8ShjitTxN4aJugqeliZ
gz4xOWmZVfteb0SpbFDr7GW4ebH+menLZLj4f1/7rTT7XaEgGE6fTJtKLF+H812h
clRTzk5DOYSSorNlfjbftciVcZ0FAe882ETyZlpxjl25oZnj1pCWpKTiPeZFy+yU
iFMWSbUFgiitjCEmG20iie59D2aLBEGUU1XCAwtJqkW3iMGUBf0rMx0TLWBPpm8y
TpdyXtcSAxSD+gyz4+9MWTZD/m1QLWCrMGsdr2/iYKWNDFIayvmdcIV4KCLPXkvP
cKlp8bs1jmvhrTeUHkuL/INQsC3h9jcoqqyFpLb0Qao8kW1tyDSLHxDXsu7abGZz
d6A0v+qwCanF6AVGYKI8PlGey20XclzsTIRirYal4Ze5gbIdcvf+fvsG1Yhhi0fH
aFg/sHAyJYGr8UrFCiwgGivEj9GmxQm+3Kol5wpaEqQXtjTJsKRnk/7dtFbZazpr
unFeANzktiputiDgy3EQSQlHfVH1jzLqxcUjJzkK0ITERcMykgZU2bPzcDJriOBO
GOQ4Ako48Sel4uahqwPG31RxA7RJETLMhUDs7y5rhEW6AyTpQCILuQYR9idd4LFX
2fl54K3kjSYDY2vkSErQV7y5ynqp6er0UP5Ghh7ac5gaAINMcqt7+qOmlNv7GCO3
5nty0dfWwlPKtF8GQgctp4oJQflUuZUT02dz3CwhDmsLt1SYlmclBD8OJOzSbLUy
XxO2hKfLFabc1/yX2yNaoKGMjRxn8COLMFARZdIAkun6UNy9kmcc6ohLflc4sinh
ren4EtND6GPpf9HDCEY6sDkskvhi3+rP5soFuSArPRRZcj0/h4tP+C0f0tshtLZb
WJEnlaohEvtwoLOiYg8CE5/9uZuBt0Zs+7snKWJ+ytjPFK06pHUD9R7KtML30YAc
/sLSrIDny7Wq/7v8JRhl2A6xIBizUFLCqWRkeXrdgWVzc+/hf2vNFEqJObIJexJy
5v3RM7UOt9/uZSDz5FYywmjt1oR6mXSP6oze+kZC5Jp75wpcAH9rPR7TuLcKrtOF
j8hGsU9ciGDtu31GC/pBKXU+vz7kehRP84hlF5jqqRtzbZDpmDBVn1Nk5881kwuI
scf97e68GLd9HPNKJ3gKuzTqQsse3/LXDVed1elSdt6jaUZs7NABaWyvNj7faTsY
0J4x+zyr7kXQMZ00Ydilkml9lGn2L8hJp0U+sjwQJFM5BTyDKZM0ky8YC+88YYtL
CTt7IGQ8OZT5ew2B7Unajvz8tZqp+bDSjaO2tUif+2HuXnfBlGxNmeOfB1yG9175
5kHLo8N33AnknUSIoBL37V0ysysKsJPu78jJXE99kMtnR+zSWZMtPyxOMT5MBdbn
JAAtdPYW/XaLB1clPSi8jUYzNUeZZCOrUJcrNJrIvKSbsH8XFSIg3IwtfxYK4Eth
DVNoyIEl9lZZ0G2IoU6dEeCddrQHpZnTlVrZDsZW5HcMqB2F1ki9NOxh4WY4zO/X
VIrUzv9o3Dft5ZlJiaCZzw==
`protect END_PROTECTED
