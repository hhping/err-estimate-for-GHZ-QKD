`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDG0ifw+66Y32OATI8KHI7vX7fFFQA0Iiev3kHIyLEoGbMaHIv8uWN2iCuGN/tX9
cmP9Aelocvjr4w+G7HBZ3GfAKQODwOMnqj3nPvGyVmiBniTR0jL+KNrAganIF8sw
VPSkyCHwgYlIdb1AtDafxcLEKo92OI0gol+C9rFZhIYBe0Sz2mVAItcZGBGphmu8
sKYzSd831TUWeVM5AJxQbqlV7uMecDodsV4DXwjsE7MuVA67DthvTLPOEpSsu1PO
Ey9ueEMWamQbJ8pRv12hV5DGHqNFr3f8Whm+gXh62aAqUplaOak9q3cp32sp3oTR
Ppq5gHMSUZpEx0xfpqenREc2cMVzZZl9Mn++4mAgudwnij6r7dn7/epdMEvdGys/
GXWdFk0m5XjIm6xM9i28x11YBJYCiL4JM21Sa0ZoXNUlJpLE5iW3t89PD9MVxDwm
SyUnIAHHBUzTwFCTAZT9ww9xZxsJg640l2X580gFvkx0WEFYanOO+eIw1ooixMfl
H8n2EPyy5/Gu2imkn+pxlHsIfKkD32BwkY8eCbr0cyw=
`protect END_PROTECTED
