`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tuxLkBN0PAu9t3gODQ8kcW4CZypTUIdvNaVLOnr27y+jX3sc6S22jNw9voSXnyHZ
fgc+L7NqpdTsL2YLWj4Gem7Por7mBfBS4zSl+rC9sFebclXiexGCIhWODF0MfBTs
abU6CzbEDnnWgzxCM5uRDZcZdFZQ68lg8PHShRsubITgy9+ADhvKCPFxEBb5s3Qv
vuPaKif2rkIN2xOp/gLzGMywk5hZodZzRJ6tIpYn0zrd6Lh9j9LL1pJTF31r+q6g
1F1b67RNCIAW4RPI0bVK33EOKKYovbm8B+pwm+QG7GJFj0t14oN+P5Fqc5tMD6nt
C/0mUx3rwaVNjH7DtB+YKA9eadQ3MiuPu7MxqBOlttigsisJ5rhdbm73MilVs8E7
XQ6OygC+818bQ8KQg5IpxmgW/jUCJXTEcGMCO0rGzHRpUZnHoadKRtfh/yfiuCU7
n60dX4sSpjIod/dNWyRWkW4t6CKkPpjUgrOxJcJGsWgri1LaAPGwJ/ou5SVj3iXa
IG81p11C9GQ8+0Z1jbN7/q6rMUUiabPWkwRAH6yMLt8IVEYqR2+IEtXkqdcHUAxW
drQWZoZ6zqs17gmX7rTjkVWhijy+LZX6XdmVuAM+3I1vIVs4bQS+ZAHGT2Cv/DqG
cXhQgDADHvzMZuLk9yQj9igDEEttNqeOiHxlODxIA1dPWeE2hlINyhtA0TehQ5bs
Lj6MNUzKHGCKuF9u3RONEhOI/bselR+AR0/hihAg5sIUYcp/ahsA9CWjJwl3lY/Z
`protect END_PROTECTED
