`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VWRth5V2cei4lLy4+TDT2tKRhNaVLWiwSUeE9qw8Li4P7sTRXULcDJpmg4MgA3Vu
DvLepR4TKJ+7EqB/r7lAzpKk47KcIffFwmMEPZ/3ti1kRP5DLGbymz+o3xNafa9N
R8FT1nijUWx5Obvz4GyzXYAr29C7EMzBh43v5FouXt0UYPCTd5N8b+WaqCrAj7Vq
S/xQ6v4PTFSFYZ58Nox/C0kvVPd3dBrpVrXSMklMKiBkXCWnioVllXmwbSMPj1E0
nQ+QJUz6ZV1hGmhQRpsk1j25YvLO7+5A7n8t/SWgxnLjR0KtgQ0bIQqwkBvJBueP
cEpIMlh85PbYLgggpNzSfIQE6dDn4bIutpQQt1lfhjrrwF1tHg9dzK5twaEeyiyA
U6jzrG1sTHxSpmjIHcuMO10cGkaZ28JKTxHhBMUEj8Z068pq9uuYj4vjAoYr1auH
2rYUVHcusk6gQ3jTHJqJB6Fj8XOT+4gRi4F19rKTlERKZ0Rvo8p97l6WilCoJj/k
/nyoAC1B/hi3yk+lVMY6Bk7tkCpJ/vBRIMIHFRMQAX9Ly8HZ3WH6dGYuOU8OMbRq
S33sQeKWbjxX+81+bpDAUC2pKJfw/XWusIcQlboodZWHKTIoxoGRS9EG+LNjn7Jd
zFNpDpzvK0R3RUDxJ4NCxI3nXq4JsRP2/Ke4vVUm4c34da5jwySLwI4HNm4n4aDp
WkO8iUfgcMSHbe0qvWc+OatmzU/92+odfkSZUJmtEPwKgNWsOvegkKqjvRJGu5ZG
Kte9BqbHcyEq2Jb3MURfBpXwClvNgSN8dN/ai/h8Mdcf8F6PGmHEWlKanQnmrFpT
MPzWAh230xlhL1O4vviDZrBgxodjBK19ucYYZTXD6YRm7GAapSWVqbZWGS9x8m/a
hydOBAIm+2W5j7XAB0O4bcmqBWK0LJu/UbLJgUMAVL08Gsouao7gNqlmN5epf7Xy
X0EAbQ/sDKFii9oof7laI4UfSlyTbfhiseVTfVYneCZS0dsIa0/copyVe4ZfLiE+
gzZUyyRHp6IIi/BayihBmhiOLgdYm+GmdBR7I7CjUpp2YJLoFETGa2xsnCs42t+k
uezupMk+zAsInDE+mVZTvu9ER2irPdv+8JwmcXs5e+6yzbNnk/m/leMz6D10xUkf
jXVppnwDw/+ft6lcJreOYxGP0vlY/f1u/CYPo5UhdXXCEdKQBzLisIH1odVZotCn
5/6lPzb8U78AaVifEIBgM6J+HLMjAsLHRUNW2sL7AlekbuuHxpoZjcMWoSLXxL/J
BLIcsj+5jfpliLXFmDDOPZZ+JEmLpfphM4Jh2A3QCyeNYoo6NnIh4aRsG1F3MSD3
bdd6P2Gz8Cx4nyIoQm9WXWDFkzRfRXxYl+B+B4/AA/UrBZyAxkVLh7MMckP5/jJd
5V6JuOP84fdehaz8CZTMg5Ezjwf8YLK2h045cdYXulg/gx5dlS+r1PhBgiF201zl
zskwZnemEBwk64lBMW14u1H8q32Qi9610m6BIW8cusWBekTkfKevcI2tciBGOT6B
VRdx3wzP312gE5pvawjGVPfmwJQkdOKjAvgzUKREGHE=
`protect END_PROTECTED
