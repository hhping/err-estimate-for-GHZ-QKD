`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElyNRO4b0eVwZqxxe94/wCIfxVi4O7e84xCEYSO8i3c6k9kZjeF4xQR2rcU5cjfc
PiVy1wn5cpnMpeAg8Em0Wp+L1tIH8Vr7zNCmrS7pYuBwB7aJkyAaNhyP5BZd1mdE
WzWJk0p/zCmkgrQlBqceX8jfCEQjTbtO6ETAy/KiSW8YAzmRIzn7A3dSn7XveOww
ig1abRQnq0RaMO1EI5exWLdqVKjCUGmURGNyx6b/zxRhcHqa2UFpx9I1yjuSs4rR
/GlRTo/DtbqiTaWPoq6Zi1Q/xMdn+wbG/grSEyjLGt1eCR81EsXcwxccRNBRXwRe
q+knj1NxNB6S0GUW2I1IQUZO++ytTFauUVo4Ac+WldkRkwdwElOlZ6OBcd/hXEXp
OZag0As9+WP8+mgicwXOi6YSVW3sLK0HzaTp2P8zsCnhHavVGiSax3/4+WWtvD+T
kwcI5U/U83INNvXTGppSxgctyLbxSqzY/VzHzuW9V2PC0cngzRMjxtVW9WDUVERw
0J/Lr5wdudBH65n/dKKL3Me4ZHZAOB64uyPvwF9D3hsgnxP3P1yszSFAYuBlKy1Z
6N55AMSAuo+nGUZz30soJVm0LhGRYwKmT9JGT3l6Mi+XFb4DYzYgcnAFR9nTPxH0
bFhzaCKN6AWyU5qh03DPBd+eTU8YyHTDcL5VzlWKUaU2MIaA9qqbpuiCe2W/hXXe
VrN+/XIHB54CqpThJfJSyfmK9rW7o6hRkBpu1YkMIfwA9o4AtQgFtrDPudbFtxYZ
ZRibS0Upx3lMD0nGN4O0/+whrxMXhK6phTrHbnnCjD+Ga3JlhOnb8OuV2s0UZ0cd
uJM4jaI0Z88Xc7OEhbxmJS97Qo4kGO9v04RObIt+UpBBW0BtPKZqyb36waWfsetE
FsmhmLVzhcwZ24Xd8t7HlTLyVDBVK2EldUrg+yKsmyL9+6jImEKIDD9UoSEAjLCY
al9WQbofYc0zHbhLCAA3Dm7s5jBBbA1kvOk1xr8ldVtxNn++9f0RhYYuNqIs3bNm
17/z9kmB2bsqHcp397KPDzcpQQkSs/TjDgtcQnO9i5E=
`protect END_PROTECTED
