`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kselldIw1dAyBA7sMMZunATgMakTcAeVF85i45pkjtFxBinwp+RqhFLiV9FmOl3h
cyF6y8mRmeHxPJaEkUak8XgCX6fiqBYxIykN3jkx7PXnYMvxWR1PANgpyrFVI7hy
tZwgTKNuqyUc9LfXZ/2SwC5hALu8qpakney3JDT278OF9Lm2HG0clELV14dp6vZs
+/jKLkVFHFg1Ng8OYs7I0fhN0Jb83avs/rSpnkBMj8DXulU8nZmveHYmTq8RGPvC
yYGWPrDQSsedoYThg0TmK00y4ojs1Hw07drJ4oEfoEgAUOzJTZwemgEZ+199XfxU
5PFVYeCdE1qJjLeNgZv30Lb6UmJFDYbIP8LC4LU+4qZhrV25/TJONP3pzTzBChRF
c3U6/VYqxPxwe1BOsUcEg8YoZiQ61yHMWvXEGm4qmMFQydraDITHeykioP5UZ8iG
H3Tzn0pk9vTWan3eXYsM9AoyNphqAfScNSSYEP7FW9s5qr3HpfRqz+Qe7/d9HThD
+m9GyQoimiVVtjhL+8GEhjUxZvd+2RQGZVVD2hfAgAGslOIEJgEfbWq3mYK+ZGf9
QPvwb9aSCEvwSTm109GIGrhAIKSYdrkhZZX8MZhPv4052lRjB8kIWKtW3l1ExFfX
g0GcxPol4E4qazXviNd0tYW8NjeG+9o4d/r+bnOs4hgV3pASCoxEPqONtBp+TJ/5
38s54GrvuYJ+d8Vkzo89fE4e427XK5W5ltQu352vaZuUQwCnBVE9m5/rBz0ussVs
B7mKja7hzQ9rmm92V59t0pUNowmqYu7a+0HVERzDRsw/aXTtSiIX5EUE1A8s8d2x
FJCTvcCzqW5DWaCcxAM3wgHBRMStZyCaR7G3CfI/2KzAJwHUWdacDlOyBcYzzOaq
0u5Sudfr43EUWtM6/Sewxn8gvhTkBGp2N8SJQ7dg9AqT+nfv+rBecrh3vgFTzBva
uKXaB0iXVr7ITu1LAnL8Jc5/uC+8FV7bNMvoVsQ9WjcBnDDgErkyEE17k8UbDgWl
ApkJWjrRMGUBtTfg9TkUCu68hfZEiUo8imE7O+QlRQS+lKK1kshlj8vtHQv39+Me
hjAKlba6rShWx4F4UcaKHENP/TINQCEIHJmy/NNVhRy68Ul/JGjU4I9fhGnu40u+
UlowDsE+KFfEmjdzWrCCfsNv2lQIES3FKBxI4faZ6gLPaC1TNDCd0Dio4NA3ioB7
OLyBbUEScDGKGI9aXrvKsA/vzqJAR6a4Oei2VkG3tWWkvpaIBWfHnHEBv5A8yo5O
XVzyR1sFOhVhs7aFonQ8Udjx/6DkoGrXRuM0CprP2GwugGx3BOyG6ewkb/5pvlEa
LE/RV+qazMWiNCjDwMznkLRcLSneylgAIX/ABsCDUZPdgWj7dQ0K32D4KT/0mKVW
Hw6lnn/rI/H9REt3wTRSBZR2ABrRBJtELdbZcCvddJ9cLahNsvdv9mR+3T0v6Aeq
ZR1mrE4TAzmGQflXxxnP/Bss6kHOuLClVSeu7MLik6ruMaDp6EJt0DQaMStxa1fm
LxMDPB74ZL4UZNbLXcPq2RFu3dymDbV8hDBN2ukRueHZ2J3b3+3lbDejhlTyoZ1u
gRFq5Tqs9VoA3mkvZoz4gp2+kAgEjhNnFKHCV74J1ofLmA1amh665VYho5CGQOiY
6mhhXjzT3dU6cShJcdhtDNyOvsu/Isa2Cl6bx6X6/XvSVLnlvwfe5Gost0fL6eat
o3Wcf9DVcB9CM0mg72GQMzEYnMfF9ei0ZpkxbRCzDOSIQ6aKrgd6vqxZ8/OPQPGx
KT04Vsglys8YPgqXjg4koSWnl7vjpM0z3jTXt1cyGJg5OPF1xt0cK+LAzsPd+3Nb
dU+G7lvcln7FnSVQsganmCElr5zvhim0/tfXTPJ3MdcJskxP892bKVJS78hl2oT6
aD35I0NHL7nVRgiSi2h28LVNNeI/Edpz0iFk7WwwjQctBfu18h0VnVAXz3tGutoT
3RtlAx51WQwmPDcmdkzgZJm/ElXCA7WBwg9MVF/ig43xff+tJjgpddWxDt40nciX
UArsVrY3k7wVB7TKeofbhWmIKZWVNVtj3nItxSYitPYeujYwctmh6GX7o7Kf5WsI
mIPJ8wd+cN9DtGlarBWvWrKN+TW/OoAGtcURs0Sr3uc7xXLvvgKmF4z0doGui6Qv
L7IXGbyroOok8uCTy/n0/YbtTbTbTS2yfNx0h2AeZCX6LUj8vLNI5ia9/z5HMXmN
N2a/2qf3ISlWj1PwhRyyeEiI0gyMKypmPXm4x0/1lmDr3+7p+ggqyCGe2oZa2ge/
pKfDbJpzbasGhevK1H7k8HHg4QYVEgvskJcit8DD0CYa1A6eED9jltq3KzNK6zFA
496DGez7wmAGhTS7LZ2wylOmN/NJkOy5vj6s71OlSeX664QyZ5GKBkyQrz8bL/Sb
2kt7IJFA6elZH5Zi8o+Papq7zD1RXM1TEq2c5dJ4k7Fxeu2AKFnxu2agt4NDngLt
zHDqHhzVJyrohnKyA1xJBYBblzx92Bf/iVZsBjj2LNsMiKnyW/A+CXsK/rV9Klm2
/w3WdXsZBpgeo4LylRRaE2Hemf/ARr/0GRa6zEYFzVX02InwQwsRswy/Lq25TjQW
5ieVG9II0BHn8ZDtHwdKDErBZuYmpgxtGEaB5216zk41Oee93m5zraG3qVCwfmVB
L7gHZokgnFzu6YSuziB61PQT01JMXObgScs9bckClxRqQJwTlgq/84PAaqvsWf2Y
aCjFiyEB0A9k5Es4VrRJEDA5tWo818b6aKD+h+W13W6/ibzC9pm2CUdHfD4R1NIe
Z/FXqBF4BhUEeQl+tSdQvIH9F//3D3VZEYjuqnOXc9VRmwu9w398X2dc57a4JMtA
68/yDDhuX9pM5/TRwZs8+/rQa/FgbYRI+kxySHGOuzyXN2i016sF6RPLIB66EIIQ
XQgrrpLbGd/dYCpIIms+k5iD04eT48kBO0zHfm6iqGevhEslJeg8grqfvRlRhQVQ
QEI8rDi9NMSYFfzYNo3YzONF+NWyn74OTA10b0Mqjm8KftKHAUQ76arU5u4DnFcW
QEkBLrDqCmAR5WJx5bDW7PNPM2ZRUrFGat/P8tvBfvwxhSy+ae8cROdSD714KXFO
K6Y4N6R8mdpV1Xo/0rTx67/7Cmn/jMtYGYCTkaekNPzRVtoUVI8jIDieo2Sd3HxH
054aThrl9/GXfPJPt7dpFB3YCRt7kfqSHGQm3ij3sceFrMEQId3mcXLMqactLpMo
MCfBOPAMXyFVLIQtmOtIF6XHhbd/arFeJZ5EPvWGTnsuZZDffUfpnTUFObB6MLvv
A2VwVWw0LCL5dm8OfU44W6ZkaYmZ+8ec231ngvKaOle3UVNxTZ3jrkfcgVU4oz+V
8NAaEN5iWQ1YWYPL+x8SlN1OrjLhdu+E0RYvXKA1BC5CP8chYwtYSXZ+EjequEXL
tUi9hU+sPwcofTiRoisnIdc2kbfRA5ehsKgO+9OmMHYFLHmuSzBz0Nhg/lfKGv08
3jaGw83aVDSEhsldsd573wMtDnXzjibJSQWRgnxNSQyJ4WJeG1gpVetMgcCn4DFr
+10KJbI36g/3ZkJJMB2TeyMFIxHX2l5wC0oBGfW6lofdKKyXE+XRVlkxhJqWCE8/
a8PlV1A+mqNjtvtj8P3VH+cOAx9CJQQQGJuIt2zRRFJ4rnIK2LGC4QQj268omQ9R
ETtW0WUUeMMG4eS+QJTbOvkS8EfBhos7CwQVGz1y80Xz9jcC2PgTZ6BSvQBUJDEJ
zM844RXd0JURS9VWO1/qyVxpZ48QRhLzhiRu8WgPVdB4aj2VFAkXm+Ud/XJ1bq6e
FTTPu2r+U528YHGR2P5ngxIG6CCmJmWhf1QXmNUP48P+AXu2lAza8YqzobWI/atO
G304IwKig7lDaVGVJVuXKGbIBd/DXt0NjhirsJLnsTTCHOLsov5Sfo5fkTwhZUuR
lqQ5xzsUJgL6MNKUQlZz9DE3zMEFj+AoTTQOFDV17QdoAjJ4ie7n3YQsfJWISfAI
LRE7qKkqQVHmbKqdKJXtigiikLY6vVc12JtRFiyYJYN4YlQYMUSq/mwKG2fZUoaA
grPjnRP99EZ0v2nl/R9M18RJF9wKrzpMALhty+18WrA2HXNj04O/2cMMzBX1A09b
pg+HGnaMYqmRcm0idoX9KhQgl0iV3Wakp6BvRRSu0KxJfzCzmkHADDt5+ulxHwhs
jAXATh7YloyYMB1t35Vmjo8D0icI8HuF7dastwla0LkLDGHN8DojMsWF1IY8JL87
u1xQab9TtoJCO7u/T6sZMKwRGmwlVsVaKyaAqGv/FxaDvNBDMnqm2AUWQ2AFvIl4
dWytFg8y+ttfiCemD2pGMwdJm4OnuXLgOnj2dK5QV5st95Iv0e/PGEHwret0MOCA
RwHlEJMuEmcW05dcImHRgp6MPFVfwYdbfJ13dsNZzQTn6GOju5oCrtpeSFZKJrVj
19RrLz/0BhCkfFJHpH4eBx5oaoRxyOdfFv1o2q2slU960uzbXdEVCBGV1O4I2Van
nwn/8g16lV+AdeM5rPVtuqSNpSj+HsAUyCGMIvFtTPAx6hNT2ZUEASpOgQUd/aYr
1SplCcyUZ7M15AXGMr2duRiyQCwz5soh666nH+Mx/8cOtj+zE9xPwmVBX3443zyY
sjxGaHuICiuETF6MKo29tF3840dlA/xuAIJKsLzpS9AT/+I7kYtmeN+frhH0TRmd
pxvz6K5dEQZ80Z83USLSc4LBdDQBeBnWW89xR2Xyi52avUlQ72qfIphk47POZ8vy
2ALuu66mSBXxOQAsl+s9OIFI3G5X4FWfBzNuvkrPTkfD5lrYDeaUIaISr4KRFTeH
xPe/WiYvP2unbUe6gQplSFDnGfSm1WHrJv39jlkz4OJvh/lO0FcJuQ7F0JA1bcv8
The8RtsD8j9IsYqhI8XfseESKU7uvxiE9jK6IfqimYJqbXFcKoymorwAn8HlBLnz
fMHnhvmzcjt4fV9RhQ2hLymEGgXxZyZPZqbb5Psn67TbkXR3e3QWqSZsoqXKWvNX
fI4oyU8IXjEV22LuYWzr0rAmIL/UB44t0WJxepaSHzw5O+RMnyEOt2+b/ORJeSuM
BdNKShVszETeuO4WaW08sE8mNCQrn+426ylOdVSjVtub/WmLq8u4jDqN3rz5XTKG
POEC50N47ylz9wgDNJue716FKCOohRY8fEMLcdvPO9zLkQSGvMkrFyRJ3eFXaSYq
7+42/YgvQbKFZ6uO0mKSnNaA6EI1oi8G8iR2FrAMMfATc/XrWGV5nRYHfkIySCUD
FDh6CIvumygrdbc/tb7MZlEgMP89JjJeASDzYxwHl7rdp764bQE4IFz3EK0pDVg1
1Cg45hnOFh8rbL/ETXQ/PESD49XbRUxIGdjrVZL2urmTmYjXvmheJezYMk4u5aEH
dIqqx3gIfYw2zVDXvhF2FAmoPI9XClo7JQgtVGkkW5ytmpnsMNNvBqwXTeCx1J9R
J+7qxzuhbwuTwh8tzkKWZ1g7jdEY94/S9uTgcdFJwiEWNiX0Ek9eRBN3sBzXGaC3
IAFCZ+wbwvYA7H44lQigFIDOaXRScFUmQUyoQqUlAwQ3CCcSZ7kCIkf7Y9CEI1fS
IhaO4P8c6Hj/zdeQ/pdOn3cGnnMbDyqlDGFyEaRIEFMBJsPJ4/hu2meIgNJNeyQo
J7NAe91QpYi2/yyhaJSi1+PyhawWXO2UGMD2aDi3d9kXbSRwClY3cvsH+0s6+Nd7
B23TFFTgGcRBQ3UNl8DEdMH4w2D1FKitRy14GeCkEO9ixjzXI6HHe47/QWy/eUiG
QbQxjp3O5DZdZFRdR7gqx0WCQeXRS49vw223nfvoLXK0eZAKoiwNaXMUL7RJk24E
fn7w9xfUP5D28s40YpDzzucmi+TKw0VNezaJNzeLLVaK+8Il/nJjzG63UIk8HOYy
fIgclx6M16u7hBIpKT/nWNFZ6JAITn4IGpQ5oPubn9SSSjzuQzk90DkWM7T8+VKL
TQrbzDab2tr6sIQKu7BzAfKdX/D+xH7wpwUEb7mCec8erVYLAiKEGmLUijY5H9K4
oXWDRPr9yU5aABBTO51+IlaXfTsCXSsuWvhSvJg825C766k3YorZsOMC07S/a7p5
gIfG6zjMA1RXc/2KYadbxhq2iqnK/+rOkXgF29laiMZwjDjKLKt4gGqvXZGhHWxG
POhEpW5YmQVG8cDg2dTMNBc5WOE2TZ6eRPZBahJCx2dC9zlLDyyxLDUDuYpHOLtS
xHFX8wM45L0Nmbj/x6+G2q/k8A5NP39B7xKfyM1PlXbfp1gdGC1M/mvRINog/zqR
Ibo/8OMyi3D5Mjeq/BOFsYO7K3XfIYYlXtLdVuyWpUkqR07e8q4vJmLoqBvA2RUF
xYzDfT+E2wfIgram92VAmDc9HEAXxoIPbqVBU5ieOXrvpwDCosfe+NDdwRkFylPO
Pp8Wtt4mVNRyf4RDgfscZ0/Xu4yU7J9lUxwyfaIc9gBAhV/aF4JSD3pWa+7rHdbh
Dlh36MWUeJdtfunbdbeiCyjDMDnrb/eTqTYhhtFivUQZG4Hf+qWTgju6WRVm8pNi
1tmI6RlVa0gj+OjrlnQClwtuIoMM/el1UCAqL1M26rVEhMCSsurHFh98JCAk1Ozh
xUUSZDb67mbItconB/+1swXSRuGKpAehsTrTijK1dbLl7IB8Gb+ILCfsbf7OOw2C
tj4cnAjGe1pQv8XypksyLhfl4mBtQUpdfpVYvyhNNtROeBcI2TnjqlIQ5NSOuihU
BowXDOVco03jTfEhFnWY3K2XcXcDlWgdYKph89sKEAH16XkTG7K1DDVS5xNBRAlV
h28ppE8k/TCEzYE5HnByixo6p5eYl/hojELsnYa6sfju3dMnMo8YbJRrgem24JRp
QZDV4La4PSWG19HeeXaAQ8cC7nvstr9PWnM6bLSAYklOUKi6lDP3JnSqPMAquUzP
AIrHZI29ZnmFBtbaEd9QBWyGnjhuY+sFvXs93R71dXkZCPhd5hUY8GrM/ubUR7lW
WGG1EFy4Z5ven/OLAuEy02Rc7eIWpGEFrRREtFQrskzo0oBw8o8T28ET95FGCf9S
dSfs3liETJ9P1/cyJL6C8YgGGbKRhBBheh9qUfvi+zAIpJTtWEtC09VApSPEI7K6
FvDD7Zx4jVn1Xrj1YNGfetsQtn5lEnmGbM577mrjjMpDHDdGXptxvKGxC+/AJFFx
6l76bDMUaPXT6SMHJpIFbyMhA1EU3/ZWLLlUfuTHCippFBaIUY+9+Jg1Wz8r+jNf
ErhqBbxE3AkTwB+0KULevrrP0b8Ym1NOqE+517ILvzVHlLIrLLI8ZK4U+avq3BAj
WJtLsDEcbQ+TPPKZ8+K5jVxYZ+KDcUXTclnbEPnP7u9Cjx2b3jHh+CLz9OYeaO9i
+fmODX9/lajeYIa4Kv44wpaRsV7HFZS8XwEPDCR+07cKa+BQMb9PlPAONgVNkuJp
9hPrQOdlLhJxP4mHzC+xJXSoc7STuMjdBD4KBGApAnRe2+iefX6fVy6YY6SYv+8C
oJXgYBoa9aMPrBlsOdwppNcFhnt/rrIhskrerYv3xTFfLSAQ7P/78EGJ1gU7XPkF
FiFWdkBVQ93CjxjEi8O4PMx4V9j9hsmJDpMTMEFZmJ0y4w+5kheTY3lPM+VIRqWe
O+MqFwREG3ZgzOk8J3Xp/JtRfhSbvqZ6aQdec9wjLJAWLa2+qWggYUSn8ngayoME
1pBXBkN9E0DnFhe73gwrfNp1IkD/uup5G32i0jYcUZOSfItKd+mpHFer9QO8TZq1
6+d/cKGM1xGFO5QJiWQwg0CNuLs9Qe3x52WIgIf7m0xgFmmnQup7j8Kbuaxnrggx
6PbvqCgcNYKWHw5K4odYNdbsIe7c3Bn0oFDsvvPf9+7kcnJodWTWY35cbMs7tgOU
t9kj4wW3ISGAi5KCqQlpLFmVbi9B0CJfhEj4qI/YAVY/dMQVRHNYKj2qFTK8WSjy
4umD+9qvHDNkApAA8c6mMCi2mhloah7EdwuONuOOdZuSQ6v7hKQtjvqvCmUCGB17
sC+IcxjzcCWGiF4wc2pppb/9+LT9XHUC320vsGcwxk7V3UnGZdBJTwL//8qsiL4m
inGcAM7nuhbea1etdrV3b+QS0lc+xr/7sdJ2Nu7GQV5YZB9J6o44DchVzUOMQUXR
T40ODJEdPQNav0GZOh3x/6mQ/923lA7ckaoqxctS/OtFM/fgD8rQULyy/atRhneH
3FcCFk3BMaQU00iFVQXQ41oELx4KoYz6Ffk8GO61YPXk2S84YDNiyRU/GfzJn+WX
R45+eKKj2wrXjiI/Fdkwd7z3z7Z0aBEhLfsJM3sdC0q2vj/yqTuJwYDmfHC0i27O
QYlwulvoPVmwAU6utO/75IbgyNV1WtsMin5Z8Zp/olbGFmif3Zun8BwzW4dsAsxb
0rDqzmmvURHMrSVm4fpN2Wsveuao9IXEvBV/xcbQn8W6yeuWZdi2EETYHAjrzJ0a
QemVyzJpnz111jtInLco2Ga0ITCPiolijRYZNY6/0zjREKntcF2NMcRyFuTwllj4
AZQfQuPw38FJTvrQUEkkDvVtv6tLsCsw2lGyYBxQndUZgnZ0JOwLq+MIEf3rM3eX
NfyY1D7x0mW8UsyAuYEe92W2MCBA8jq52Xd9TvRI9PtSb2+cfU9FarIL15d+QVHw
xRZiEHSapUHATLgaxVsBeVxbCEtzR6UMiBsTw55oFvdjhOviJQKO/uXp3AEqVDUg
PrKl4ciPBV9A7s6SMMFvv/6nstT5/+ORQGrVmaU5Eco0kU+dVhBbHvLHBzu1Zy25
ZbWl586DGIkhXcpBMbJfvEFlLGeAMgi+RjEGxyAP561IkZk0NBFkUOiKEHrk5bTK
go/CIBTmUKt8yi9jkm5fbbyydpA9CQ0pyD4Xis6dLQIT2+Ev9fBV8l9IF0x9/wQe
O0ubPS95OgOyGeuEQcbkzsoCf+iHGH6LUaW/SD0/QvysVWzxhNMoSfbj7uy2SXzZ
hgiDhfqWfHv50cuSLi91Ey65zHRkuY5Lzd8HY3I2igpMiPnuCEjqGctE9ZuJ90Gv
meiZ2zmpKj1ca1ylxouOD/3P3AyB00C8HOvVQOG9icOmRPGgTp5BAFZhtJm1HFpK
/0X0K9cg7/iULFcv+bf5zSgWHifMyu+geDD/No37OQpp3rFTrnA+nWLNO2zq0XGv
rvA2FmoCwFalpWY7tbi+jWDVnxJvvkztagwENSsAjrny5xAGrdJ6fQp0lgVfkNFa
x5J6X0awLl0AvFLVYsbwkTo9sAzhAxoI0SOLr3zkyEYHPuDZ74RkeTjt/7dUsDjr
hiMXhoql6WOsOQpBhqOVg+hXnl1krMiIKngXqu1HlJntXQVtbL2SBUHB2D1yo7df
Qs5+bF+dcCVmpXckqAqZcc7La1FcghVGI7KkW6GAMRLLhVsKLhupfsvyfb6RT7St
uEujErRNRqYZfOdGi3rFNvcJ76qTxqnnlQEF8Oz0VKvS5fl8z4JbshXdtS9h7RFk
qC2HEu/e5x3WYEvyXqqgu+/4ZyQh1YZvYFuR1Vh9TzAO0II2nFEgck5M7WDVf1aV
0BeaLQt5xHJWq0gT69t0Hr8mJhi5RrexDRLvjn6eidCDtWxXmQC1Gh8Z/d5G8qUu
B9EN/DKUTLMl2fxkUpKIuzVw2KPKW0yQcN+Yh6ZSEnrvu7j7LWkx/8CYyIrUSwR3
apO7Cu4ZfgQk3OfMAu24Z3RR++46vuLsWdP/IPLDSAKG/j08oSa88i2dp489xDgG
FiJoUqwYTvr2aX60QPhCSKzxphuhiKkT28hWe5DoCHgKpI/97AZG19PXcjQ6Tvng
gjxziSAeB9kK+I1vdAyIgiKWZVNPbsrk3YM3zpV5YaX6pXa9mo6U1GHlw8IWiuiH
MfjkVWcLBYxCTd4YAS7jLzqTliAQS2+SXSJFD762gbGlxNRWWWGvTaQy+TSTVTEF
spdY/Pu/wbo6enwjuKtpMtOL2hNq0hxSpbTvMBUlLk+be4Ehktjm/lX5WKzOvWdg
HjzFWCRF43Khj2/ZC+Day3ncJaJkr4pXkPhy7IlgUrG4jdek0uSHHjEAFFC5oskK
UkuUM8ihWn5XndCFUbLOzDRIxOFPK3RygFHjVOmWGUWJuzzLhvG5Dwe7abGjDbD+
eGsGR5pij5mIxRJylDzH4f+cet7w8s/didVyWbRThzoHWrNFONKQP9ertLULqMZd
4/xgTMzJXnmyNyjObG2nOVbsfnfmTb4Ww0pAl6ETnLlOlrAKjN/iit3rxUYlla3a
GChMMK3PvL8qxWxPv/H9Ed+TTLw2NTAkHRm1yTuYpv13ldOmpxiOTM4ccSms4n2q
yyH2VV16TxrFsSxK8HZnRnb3bJRhnLEfb3RCvWwdHYOV0KvlLo4PmUc10TpJmc72
nuVBlBXEVWtt6Mvi9gyBYD0/kP/AwKkE4OvaokRL2xRfwV1RG/Cpq/OaiUDyvo2Z
k9n1bR9GzWIsaV9tyiUp2lqeXaWtGSQCRSTHijaHSIx1em518hmevF3MCZEmbDa+
1d8D676luD0oWWc9BfQfBQ9j4FMLv0nisxg26Qx7JoFc1LowV4Xhjv1RNgUWGqxK
4CbJnHrSzMF2AM8vz7V1pKZLuKo+B8wWUfZn/a8yjb0Lfa7sa/G1kc+QBhdF0bIJ
gISxNt0RbQLOTFZOjhQFQ2brLmQzc49ga1UgJkhXPKMUAaQUaZnELxRuZEjpXqwI
JMvRm23O/LuD030z0LiQzvo2Qa08OHpTrD5fdZKm5cv1zTCGwqH+eChfMmeP9tmu
34CqYUFSYnWZ0soUdZm2a3dIMKtUcq2b1zyeESegsc0SSJSZJGCRWd8iXtX51KKQ
NMMjfh1aFoyFFwxQtBVhG7+yXTGspZz2i1mir0VZA/gg4bFZzMb2InfN9PADvkFK
AUNH1sHYzP5RUOV/9yDTTQu2c+/ZX5mQqFRrKoPkRvDI4wPyAqXI6IsZyYmsckGZ
kJBZ820PQNzUI4LY9N3KWELHkH+hMMkDK9V5/X9lZNGK6oe7i5TKBkG+lKosX6Nh
OsNy7b3xcA6xB7qIDALLGmqnrHv8zZEEwtMZJ8c6l5usiegYjYlyxst+GIAyo4+X
VvUkA6lXTPxF2y2mnKT4jQMpWmWC/ya8LNGunyFl+vX31E/eH8+oLWHgqSMaDmL9
k+DJFAdc0T+LnzUZ9gHtC0SD2nU71MkzThQaU87nMcxjhtXqhVbQBpLw5yZfOd/0
UH01Cc4LLUA+icHSYDraKyzyYwO1vEJxd8Q+1dtEldIG5E7tfU8CbEK9+dub/Ici
xWgBk3p54VRCFCrPhAUIyT6Y8nnH4Hw2Ig7RjLgXvOfC8ecZXX8dcFz4pSmWbjsl
UEaCMhvRQlucZAkHS+OTpXYilYViY1HucmFos5ENnCAZ9K62uqK4P65ogtlryFdY
UGt/dUV/zJBjotTj2NiOBiXReLKC+jkFV79oYW5HKIQqkWqee/JKWzYs6HYKqF5K
NBz1mP8F0Uv7iAsBzw+Sa9+jSC+A1mx9CPul7iBRmbZkc+Z5sQnh46EXCrjWz4Kr
AKReuMXVVPJ7jqLkyGcdXFS6riWzPtWQA2NXH8mjTEW2xxSoh8ROWhuwYs4jBHfP
PGxlSxLrfox6mdPIi7Yfl8+1DNXwAy/+5mKwHAxRBzIEuQLy/Fa53dAItFh94p0w
ZETljFaD5RIXaCVp9mXhBjZu5+IZvnBGjqndN8otde10Ji1dQG3QOGURRRlSWYmM
8nCRIPNGvQeoNDR0/pPdRAPz41a4Czz1P7qt6XbzMvg5ZaKema24AMsRTSex5KVF
uPXCIrolIuJ0TOKXqX6wHi8rEszjBUztHumNzPbJkM8o8mHfueSICeRabP9QmWoD
Om0AKm+RAmtQeT9/56XTy5dbXKCpA/yc+OoE2uaH9vAGn77wxNh2/lQ/6tVTISsN
QH12H+RJpy/mAYh6R0VaycxGJI1XW85p0dy16fLj8x2wfRFxXDBenuJanhtGLZTu
/56vGvd9UesSmVdBHl3X/t+sPnQ3OW/DoP9Pgv1UsOjZhLhJsZQgBFA0Aepsbwtd
LX8coEI2zEAxTYWsT9YvJbNwmvKPx9JzpVYSjsv4DSY1oCeqfCYxncvQsUhiFoMy
Xlv68ArOp1I0QD1FjJk3U4t6xctQqQu0GXRUA7j4p8hDUR5wL8qb1daYVAZ8dV8Y
9rpAZb5lkJDH/SntKzuMlHakjsjkGJbTqIryb0lFSsG2ZO5zczRJ3YPMTaEiQmWv
mlKjrgUCE18AMfkY9gLDTKPxTwIMPyMaRNbNOQMLma0RQOqF5zWOIhIiu1ar02LT
SiMqdNJFGRe2ase658bnAOzmNvAz5YrimbxH6Oiqi2C/bCQn/UuSpxPJ2f2lT+H2
c/zIQ7TA9NuLDXOXWO8SRvFaRIcJjQEZOfGPOBtgarW3k5kdhBQGMiHUW6l6oSL1
LFJMu3/HYlxjBOOAwWHaqu3WfGUVNgLIiZiz3rxHx09SFA4B3yTmC1pB49JQdtWb
gFo4P3Mk8m+8PwnyvGHop6Xiv4yLc21qRABWT+5WPinXHv/+Ey7KuVi3xsu5yn2A
z9oGoi41Yq2AjINMAcP0w/LTv+faHV+VpASDCIe/jM4OBUAs/c+JxI8Jfp32y98N
gbJZH9NmCkqoF54Jen3gUP/d47h8GClhHNlxIuNsQg3UOKy+NZVlGuEgNgTKBGzz
57JJQ2z6qfBMxBeUzKwuecdhDUI/osXwAOw2wKjY97W6PNnVFiJoW02ukzhVC2Jr
Wd0fA/vLJshDQ1avLyX5otINOp8M/WnS9ovxoG/uPvBApxk8OSqVTqZ51besxrIV
pKT3f52xIcKXxQ0svqCnjXdLk0oUG/Wtq1C5mdIHHEEqx60yz5kqONpQsVFuFCbu
5AWyyb502X3OyKxHEVMZTTO9kKye+CnOKVmClWgXa7VXqfL64ltE3pwGs3beBr0F
PzuVOsMyVhoaSx1fT0eiJrNET0gbxUqeEFWq0sP5m6Ri40bePbZ1mkgXTb/SCOCJ
RyMK8dMQ8c5qU29F2f986kXOIwBWyS9TpP5eMROOEln0D53fWmUpn2Q4f8n0pGan
N2kyTbT1tIM3WGn8ZRPhaleWlE43Pe+hZB5kmXbU/Xprxrdw+PrGMmHGWA7z8kPn
1rfr6socoxufwqH3+uCnWH08gcW+VYPhtfuJ/VguGvdBPbX8AGeBJQKREjVMkFHD
W5OUdb0zo+YKr9tUnaOwRlsDZA2+WY0w1xSXXm1r9+1FkJAI3UY8e+40nCQunvfP
HwKGj5LHVTpuaIY6Xrzdbuj6eeIVwFyXLKGv5ILJS0eEkFk9GrZ+wX1SoGP+Oxm1
diCGcQHLXyshmzLKTo2p+5Mk8cSbMMqt157Owo2wO8G2dEPgZgBwBe4TfyQ3P+9y
ORCY3wdEOqPownQ/q7+qYzRaEjpoLqiKdqPSMdHLSW67TpgCeM7CEvBVQjp10Zjo
DWMsYEbEgjXp2LgMyEr44ZrtaYMJU/EKM+gTyiUdWg6q40IoBGwsL+5Zm6Ksxbh3
s+B+FAVpEl5Q6cCgSsUQ6jxeAcTdJIwMvXNgMbpn9IrD3LWt4mSgnPfA3LSkSnSj
Jvjmf05tH6t316cYiRNsNeP1LfTrX5lJHiJA4T2NhJNXf19D86Z7BzLtyCpGZVzl
tFiEdoM/MmO+Js4wVqug8vCFIteBpWEiqzh2L/Qfv1UoJn+KzVGLRyty+Tm0Ai0A
sDSCGI3qq10vO/TqAnSWxo9wJ2JRH63vjacgyaSMDrK0/PZ6Tsl9rPdL69f/Mwun
/yr6vGJ3bwImWrHs0iK6i8ovKF3XBreMiPMrOa39pIF7s2p0vsfMbAfSF9RuiKk9
7XLtHhSYhyp03RaUIeSR/9VjOXyMfrbLJOrtQZPO/Gomk0J98sbX6oXpzAHYBGh8
0eNchHw3dmE5s+/tDWsjXPDwFZaxcsy0hOw+iBpHS4sXnEFIbOHTaoboQWf5PsoQ
SvHVyFnakcrFTsJLwhtKr7+pYDa0chmxKPzFOOI1fZ6o0O7IFqmx/wW9a1eXQ+GS
CVO81okM4zzBZr/qi7K99Mqvyuf5Rt92UolYOg5omEsfgYYMztkxbLIQ22Xfd9y6
WOb4Z0SSd808cV/1Ia0zh5TaouTdquTa+MoUAmv8jXeSofP7FRvmKKz1kaGPEMzZ
ESYGJozuPGXJEx+ai8ZeNSkll6/RZDcfeeixlLGnKworGyLC5u3e6f16KPgZWxUS
f2Je0sX4SGD5XIe5BG7LHhmeI3IjKWRjR9JLjyZQoM7b+a9QVcfD9B+y90+R2mZS
c5Ue/G1vxEOky2H5vvuJGL6A4K9FwhS8waZNm+/LqRgsW/+eAHSOPZtEbPy192sH
MmrsHsthBJP5+hFX08jgcYt9kW1TlmI0xT4fW1HCTp2XNTTObCRm523QdrQIyip4
JLP6rNGQOQiARBN9BHPXx3AvMCiGsxIrwfymVXisrgT0SNFwM3gnWutYk81CJEJM
mR0LqLfFhklS2Qvdodd2txxIedDQbwidw1bmtKAggNKdoza46JMEAojDPcy2Xh7p
PmvfOEGhE2mZypgEQRx0Poi9uFgEh8TTPrPJFwFTXLO8XoVjhbaV6JKIfnQ/OXL2
5m5KfZFJrM8kkJ8Xw6bPBDiaiRMG/h62W+uU8B8lKyN6uGTj46efi5pjrEhg5Kmt
yXZd6jjZDSsKzT4ktUu0vn3QGIyZ45bwmifGUqPJ+5ii9BRbJDfIY5cavtWcWj21
KuJWCtBaz7vjmZIHQHQl1ESaxyY/3fIl6L74Xxxc29S4hDxFfWU46WaLzLVvojcx
BBY5HmsusBsAcAd/BUi4hjgc/RlPcCRoVYrdhUA2x2buDYFrgrPnsVPuuHEy64yE
XVixGA8812ICPfzoiYyp8TzW/iWMjHp3OmNCY/GLF2Kcm9f6H6uZ2Wl+blNXunpP
VihfQefp69bdsZ4Pgemmp/aXH065jLL1vuYi8v8KyMQlWrDEq9SVmyJYCmlW6vqW
bxdXAVdz7pUpRJ33V8VX6APLVGVTfJaF9W+KzHvlkydvbYMw/XZ9rmanKDrTlNzI
2bN9UDC954L0MFQZixchIfKRcsFnNgVhRACQlBKdg7B0Shzqv4ywMUcWJNfT5cTq
cKIsqOVoE4K4ieO3TQs6KgUFSA8qZskElFSNHiqp6KJ7osvomSqdkDsoTl0G8aI/
1cK7I3kggjTq+yYRoot/nemUMJ91CIqy7awyVTdGru6mbPTcSI3YkWGnTIruPDh1
W+hCSwZY1acdAmkvqB3VJL1W8iHjBMMEXtK3vCPlzgaL1InZtAMwL0vwsgiFQmwh
NKSP2XSNNMRw7VWwFiwLCzofcnJPImdumzY9Q3NJlI3oHEzYIXJ1L5RYGpIJcXLU
4FQKE+ZApxjsc/23HoIuLe/Z0xYnNvTB+gskUCfIzLWU8XPde2b8WYbB6HfVMLmA
INimA4JXHWXOi9RaCdTiUBd9Gcrd1uCA0id0luIYL+OQLVnO3rvDZ186XSmB7UqU
4cyEYvooU0/5vlDjUsH0bO2df/GDg+AkBDqVuo2a0L56qyxo8VoW/RPixIkbWgJF
6/PnIGERl/SqRX5Fu0DCdH52L1k5h4LKTCo1/kYXxpKLH6CYGDySOITt9bFTelw/
pvCDaYegLaH7LjUr+uUQijgaKXU51Rr1nx33XBJeZnWfm8dHGWTMh87Tn4xvVcVr
FC0SQAKzHb/lsfc4Js+fX8igh/qnjJFKuCVoGTkF+pnM3tjF13LkbkL1DwBAEI3/
mdsBJUfyk1k5J2VuJIAtZuHP/YXwCNP0uhx7gT3a2JfPIaBIOLpiFev8/1MwQOyM
wL9wrnrt8668QEJBj+LujdzUpNWQhatBHJDYeQ+vHm5sUP5j9acWnEtgpWBwBHQC
VoYBGyJBO4eTQmXEGXQIbDbFfFUlcVoGUuTqcrZi2eRJeiu9t2H52oSlDUtgCkYw
tMHPxVuvQFAO6ZH82fun/vVliiXZJsWlixWp/9OFKkPY8bRBt8GuyUWTcuObBvr1
WPURrJAvDrOzx18064te0x+cYsxYl02RqhE4hxfR/eAB8cRrND17tfILKFOjU8kD
09cTLGa01UDxSltJDvRbOKRpT19Y3J+M9lpD1P3dGugCqQiXnvMAvWLaPm+92NIo
/PSQBchMJ0gDZiavTA4IFJxTjCIXPCqrLRp93i++bbh8TT5IU3PRFe4FXxET2OuS
OUKxrOnaTOx8xf3CmDwsRN0xnC3Canl4TxkLlV/jRwIV9gK+j6cXQ8mZBQkyRqOW
XR0Sdcynb2n+hq2/YwnZw6lMFYCTioPFTtFPlS2Rz3x2HkYbt25MhjZduTs4DeWI
pz5PoYAtJdDD4epPm792oGPrZD+N5k0FR2sQ+tFherXESkjQDSUYCnKNgEKI2Qi2
8m64O2I0i0pv2JAB1OifKCmMB9SautmwLI4iEFpSF9u0HNCz0jTbHxzrLJ3fZp7K
1Qnkto5qn2gw2ss0E5gKJyBF2EXhN+risH5GSgp4MTP/Qc8FETuQdsUwXON/CNfc
EQJNgdu7bcxWsnEs9Lgee69Rmd0JRY4mZO6E12py94yan347ABMnHiKOt9ugaGIM
TyBi/telp9Z7ODQwd02FemqmmYnzRyHUI96rptAgKe+n2B43F5jFqjJzAhz203Xm
sVvmyquATXxfuDTxbuEDRepOTpCfNnZdiqY0WEPZaGODhMehVu2Z1W3G8BxVY0yB
qZrhUEMd6rr5ZtS874MxgyVYYnw/4E4dD2qtYJM7bTUT2/Al/0TdHUogYMMaxdIU
CoH8IFnQs8ujq1OZprHWHsuSVOSVbmvG/igue5Il6JTHd+Prr+JEs8j/2kRAK76a
W2RGB1yCtanDD9s/n+gwyUGSwYtkqIKdehuJmVX4Gjouc/6jw0xb0kjMn7+Afsvt
8E5lGdvKJmlpHjKx0/TVLc+Z+bUxCMpyAQ4nqm4DM0LLXmiHm5nGDFyFsWc1Hy43
iwT897kH/k9BTVXvCIJdI3PD7lf/n2Bv4f/TP60ZT5CtETvS3/9AAJvbeUibVX7k
PLtMYJ3UtnssLCBLJ76Jd6O+r9B+3iZGBg//CEV/a3T7IIn1rxo3ZbE4TtMLUCeD
2GFc9sTRBBG496G9ea+UKfomyBtTXXr10bD5gJMnu+Vuyb8vJalKfWeUCiDp1G81
kinNa1aIFbKLZPx7OnKXwh7puABI4rHQsw30dR8aHCm2hrK59QGdPBLtxqlpf/W5
8gS2Pu/Qf9aXylSD33DQA5T1seQR9XB45sI65ou4aG/sxnRVXwtpqbTI8sM7gf5C
vmx6CeyXxTbjAP/ueKUrLXIEQeNLIQPuRA1nSW4BJ4g/AmLevKjnvpnOw69RNzm2
G1U8CyD9LPaDmEeAHyz9BF9HztUq3QzNfnW3Uw1kLJkMk8DA0IJl/7XMXXwOB3Q3
reRBjuvZeDeNzRgMzKzJwxAaAyuKmzwjYigfunfuzH3gWf0fJhhMXCCaEov2Gf3s
NJ8FKnic5OETkF0cAOIESsEtyDBwzaClv/La1n+idm72cludVSIiKCAvSFcRaAEh
+dme4mwf1LzMDQwOV7AeAzLSLTl0QkePPpj0y1mqth1vejVD4zlKad9TXvZ9CAZv
zbdvosjZbcjEWSFT8i6NMJbNLstAENXlrr10QgGB/JTBEAO7vc0WxQtsBSMQH4jt
ITfOmhyJkeWx3dQcUvo/lcw4iryis1+iAEm8si8xXerJaa3h5gHZL+My1RXc0BNC
nIYtN8k/fVGbElqDRXExoF5l6XT1+ijUUcEpsDjBdoveVeti/aDYviV/9by8Cj80
wYgd5i+3cV1fSzx20isWQpLA/gbXH8Lj7MOLzkrYmpkdHpHcedg26VFpLuhkM2dL
nFzQ3uDFpvFQC2CowJ2VeNrD1xNoKoqebqWp+O0jDGWsyFI7WjfxVHmmDd2jJPdA
sE7MpjWGQmHagOLJgnFu3JLcEt94klCXtMjFXmrAyK70Y04N+Z86hSb2MzCRQanc
dWSzT84A9Qxz8oN4kqYOXPg9lD1wKMttruLYR39AYkAYTUoOCdOW+k7f33bieTGf
kZDHwkhk8vkKLbtiOypqg3DEjg/Wp2OALp+hP8hGhna6dxfmY6Z0sGzwRVq6XGM7
zBqVoiYc33iprhv9FL86Rd6t4UYm2sYvW1CJ1vRROylcbe8bgP2N/q2Z+Rwwns3A
E8x/ybX+DE1OCdRcoV8m+seHiksxvNziQ74Tu5n/X9TexAJLuZKRDIbSgdE9ehaJ
by1uTJI9/+tz45pfFGF3vRHk8LzMYsZAAg8xlzQIpBr1cviVVKUHLFT1iTJJfgUT
XFjoTEFGOi/N3FNKOTH4AvTcZEukAOMg26KKt55ehxJEvRF/4MDM7HQ1DPSTZaKu
779N4neSeJVY42wZKh76qSe6cvNYZlSo3jHMtUpVCTuOfODwSEPW4ASpHQrF1RyF
5wuSZp7UubX6BhVw9qmhL2wiYSXq1exaupwop5WPLdQO6iUiSjeSUNz9EAcqo7Fq
OM6J1W9W/T1eK6SILNnoPQqg2x8+CLz9/CQkPxUqt5vwQw3baDDH+3SBU106RymE
cpmA6IjlK6lXps+2CfY0QPo3ncRFrVhqIPCz2cylmAg=
`protect END_PROTECTED
