`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3MVjH9Iv8WO6wtJKOipHyVs9JfvrYmQRdkUZ4yqPCSGf1gjlR3XR/i3gVb0nW6wr
yvcWetIo2vtWPJs6rQ9ei+Rv4AxRKpGIGV4fVxUpVCrwuDu8EHbTDdkt221Kc7bc
C4JFnUpv/RzgtWaJL5b4K8Fpam2BaEORaLkSVDT0wspdcEQqDkpGmzP76gp+14ar
sahEu0d/MYukkuGqhcoSKRuJcK0HUi9OA8qECeVoKrMKt0VVdAdV50C9d2T7Ha+w
66sBBLJUUR5+0uX72B612usNABB+Q2jpRMQYkJiYxeaYbbJsX1lBU30uVPKEuGjv
4SPG5fQFlUiVWsslaLzdy8A2EE9lu+03ax5i3G4zS3xCOBXSVY6Zoz+eEsJPzQQE
dnIoSbT1qRz+bhR62dq3vfXHtkfQOEiXN1mUUIkmEynKcK3wNtU/xYr6GT3V3b93
C7yuSU+7d8Cyli6ipfCAovXK9Sq04794eb/oek+d9p96CvMR2FSgoEhrhzMSEQvM
kFdNn+NFbkrnU3InJEorXLrbflF/5cv6vl9gAYiK905LcNuA7T5gqEnLZiyaLdpu
tDvP8dWOjlCM5wl57CRU0GTKY7uJre3lftKsR3DdAFYJ5ea1UWBcA1SRUTN1dACe
YOhYfVJxINKGf0iL+jrn0lK73ibjSCMKcEdOxYvSbKQ7E1Sda/99rbsaFkIlMx9E
LF+5RUxhEgT/q22J2AbaGv9xOu0TAEzrGgjAy2IWLvzwOkazrEwlEEbSRv8vXl3l
jykPtYmm7fxmeFYAtbFu/nleNx8R9RSCQTd8IATn61X8zVntKCsvvV00h8rjfOc2
pk6VCH602jJWbmXqJaLKQrrumEkVaLI2/MxVCNrzd6tBCcFFxbS31EYtwdc/XSpj
YoEEjO2HZzYSBLu9qzw07IeeFGkVaRDtJK49kgroJABEyHWVGXYjHUZAyara8afv
5EPYlk7cSPYAoKAQI727qNiM7n2cvX595ESU4+p+3zBATDeV97l+a1jjj3hC9G4C
u9kYE3EX5M9mIkP7Q/nVE+Z7BsfCHTnpYFmkxFOucrRn/cT1NZglRMNwCAQBoBDZ
jjbOkvceQWBlSEu3LxnXExt5pVX1E7qqmurTXM7BZsDIs1vPayE3egYdOKJYqnKK
W/2TAguLm827Z6PZY+s5ug89o0Iz1ycMv2nj7yAYYOw0r1yyQxpNg3TbZsuIQPVq
arlK2t6r0OH5qqVQD/O68kSxCgrIoEdooU73gAqQ72EB0SGCofRGEr0ZPM5A89+W
wOCEHrKVutcZhBX8dqYIi63y6HLRxyu4AFeF+n+xUk8VYPSzqYNPYMKyns1LeP2F
k821xsYXkAsSv3EZ5GX7ux+0iqwPTZJh4St7xRTSTl01HiwfMtlkYeVlBPEw+mBK
pJVzNP+PByXaTvgLW9OPp7kM2y830Wu6oSbIe+DZxh8Ed/xeXdX/M6FwoS5bq5HG
Ayeyezr8W6q1/6G2cEzgcYDjGMHVzaZSVy/5scKHyJiwEyXrBv2rkL93TUlRO18V
o1tPF/ePOov3Qw/FfwH5v27ht8Fc7wwydabnk1HriFNVcQrT8fDA3vFowHkHqy1B
lJHbG4uVspe6PMveZyU+0LtnAqhYSnPhz+Gds3ud1mJppwmIrVPLEfWFnvAZnZQx
+hpvVYhTDm7kxitauYFFsMdNDuM02Zw5/irrxqAruP1inuhcXmmc+Rh2eNrtJZux
jI+GvqBdO8xiTbpV0GY0c4p0tRSMGeVcmVEkOx+lMFIKkPnIxCZAoDQDXiffr/Fc
6bAgXy/BgVi1jpkzIh1zKAoJ6rPAcQXsLtlRnW2PLUX9UKk8QbL8Z3LLxQVpO1iG
FSiWwThPOl14kG/GlmpZI4NagDrWzO2nEI2SL1Dm3/D/NzZYVhNrimxMxFHQnVAF
RPiLDMREL3V4F5D4LM8fl0HnRIIGRDHm5PnWbuv3XnqeLgrd2YkhhuDXsORRbMTE
t54mWYNWvgdprl2EKsleiz0YNG2PaQjM/93pJ+jhBZ0=
`protect END_PROTECTED
