`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sThdhulHnmFOpiK+z3c4FZgIdMrmdugMJ4rq7SvVSiUmiZACNrs/NhcvlKA72+Y
Jg7nBXAdnWdmTS6bJ84SvFYTYQcio1Ys+nepF4V3/ERi0vjCtkpR42ktxOWDZFSP
33Z3/t7MFZJcKJnTcTCp27zezzWTP9qeg9o1IzHdsbMUSwStG4H5fMMGr2bXaQql
Mv2ZHuEanfWTSfzZGAuipUXd4l/FniZgU2gDMWsYpOYPIuOM8lWipzVeslgklXem
p31lLWCW4CQPdMCC07hfP2IoZ5lJPuguxi6WZAdNatfOxuZHQ5SuwivL1Dm+VXP2
tkX/3GDU1sgp3SDJQcPMBBi/hm6aARcdhGeyxOCef06nbmq+cZV8gbuOl6Esqz5V
JKArcUHDF9pCrFwutzQQyJfxxqKJ4wsAWde9fEXcDtFIG5dfSliGYOdUBkZkheCJ
+Sx0/p1R2BYwL8t7geZnlfybySExpIp6QJ+yQf4eMZ12f2jFaRT46JCo3v4CAYlY
wuX2EYdpnbvwymdg7DYpM7wn0qGWufqn3jSqmYq5QM97VZl/Yq2GAchLyrb84wFp
fXYeQmnd3ZgJyKrRMk7FekLonxGtQ2PsDwd6Otn2fXpvALcsxJT1WC2PM/+U360f
caqw9Wsf9y+qd/9ggmwt68369kgufg4Xy9ZlZedayaG7TVDxSf4L6YNIRFuZpdXp
udOSpKi6DLjM0DyWQqvWy/JOtAxWzw2btJVPeKFEgIDQrVX2pnSZbd+r5JMjkaG/
muovpjoKG2Au1x0TEN1yi813hDerKC6JIU3DkRhYLeXx2bqFvP4ZcJIduJK3bmLE
6v6SN3brzwyAzohN4IZAL33Zlsh0oBfy2FQKqlfLC2igR+gFeVCCXW5rDfUqpFt2
ouqKnUZ3+rOxdjAHNB2YhVA7Auh6i1VZtmB0OnIiZRDjHQ6xC56vuFgAdwj07dsq
pEcKgJzj0WXy2PIL63DEl+S9PBlLTInWtdh+DwDY9DlEM4EmRV47vl6gYXgZzSOC
h5KWsj5lM865PaPCCbuibHpH877oOprJ6K14p0Lf23cwe24ijKCT7oTzCGz33wxx
W9XNRyHoWBetz8A1vJ9KmUU50EGfF7DlvkWw/tjHNVwxm9bzgYpxcndxtqhQTa0f
eDVbfGdQpb9CBRwjvdxfkcx9IfYpmHbgYJA1AP5Dwi8xrzADU9+ImU8VqXPcyopn
31xbiYstG71vIzm47KFDzSPoV7n9vdCmBRh39eIkQG9PEmcZVU1exFThy1JW9cmR
Ic6oHULqgFRh/eX2hdZvC0OmaE2aEbuSn72W/KYIMhOj/9VOvAPJpBZpqLqiIsvb
rQVFPQ6cURVV0hvfFK/OzbqSP+4GPEzOz8LK+xGmS0OheZJc0hhETq/asnvimdcR
6TiUr76fLyFM+XkznBHzm/WzNLUIO53s3bYJP6BQ3ZWiurxuNx1q4OIFD+Buzq11
uVC/Tas2UBqnyju/TGwfM5+ig89uwSlyy3zbkxECGX1IIc6z8+0gpCtznOfBJJRG
nmOwQS0dUIC3nfs/7gRkdlzNmDWPHa85PzlGSfJr4+iiSybeV9HjMj61TfKEXSUM
xXdzpzCT2SOGDw7PhG3iXgaR6vdIzE+4YHsLB/u7IFVbITBvdQ6W7sakzlVB2kUX
LY1A7qT8K+t5UPQC1TZLShsFJdEROUeqc9OlV6l5XPAJ58j/XxPPoFm3ClAUl8x1
VE9is6YWr/wIx2mWRJigpHZXjwW+ykrJKzqyWIQ0V2tgZGfYg4fi0q6Ki5PPIX/j
/tFQX/hL1WawKLmr+AN4oDB8rf9GEiJXhwNaiMYSFNDTjOvVGIPpbBbT5X8tdWqW
XuBpczArevEci8n+58ccXGO5Ev5xWZ/RsSZW1XhbOrqNjiVnraifP2j6nWmkbkyZ
9qOEkJmiFDfXut1wyEFb4DXn7FGZnsyvhjEGgZLs9YomR2+Oqkwc6jQ8sBjincLL
94kScR46Wlg699YDt/b9XVQCD4UcPhFAj0DQ1v6cviA5ZT8mcDglFhQYUKhdVNYk
jwWe5iu9+tfggfGEg6UaMaYJ4PSm/fgbghbllxS+eZAsmJnTtNNaaqmuSTC/0FgA
cHSBbYeoUhNPd7bHS2j9plnTWWCmmhPyL562Fuu7Wwx+cYoAwsIVxyJpaIJMVZtg
QFbuobd71OYrNDGusUE7e7+qOyy4fqwCUErzY+1yRDoPbrUnfwIJKJScOHENGkyH
lLrtN0h9J6fk1zKR+2J2ZGCXlkKg0iOXFaumOVnW3G1Ic9DcM1wSemlVo6mJxT03
5ZPX7IMQbGglP1jwhEsnJrCTBFTZPxu7ues2VT3KPDdinWJCKHsLEkwIdmeCEnVC
OuAwIN9C4MmHK3YXqNw5VWmv8iw/YEXfh80kMYea4aTrhTpKwTTbGSfFXWUJGn35
hRx2WKgw3BTtroytE8KNdjPv3k95ILK2BZTShM3dFy+Z2iE7eidhnRZXk1sIWRs1
wRKm2/kiZ4xXa9QxZh9wxQ==
`protect END_PROTECTED
