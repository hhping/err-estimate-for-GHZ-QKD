`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dztS15cQfFuTyczJdQwVydEYOQ3vg/LAiLsFBLc8SmdH9Lwond8D7+vjVIe0osdI
SgctTRE67piam05AwwsufwFa2WNtu42yEOklouy3fzY/NLKAmtQMD1FZ4/vQIE+c
+FOAfjRxKt96cgp13j2F8RtZzi0nF4awrZeRLLFRwT6/upMg0JJgzVdjcugpC6aQ
cj1tAVeV5M7iPxXBZ5qR7XIMxA0VLLpDwAa9XaNyOBtB4XhHlHmIfumQngIxEFxv
tVVkp6br7/TI+Wze02MkZ25WL4Oy8PrJn89NlW7dJGuoOFBQllufSosVmk838wH6
Ko7yl48E1JXDhdmOY29Kxfcg//cnMpZUc0XyGChgN5+PT3b4kQkvDBmkPHLH5t9e
JC5gHbGTBqoB3EFtCwjMJcVLw5TsVo6k3d4vCNfHAKooJSp5dqaY5F44zbG7FJxA
UNBwgfZCxuYRkdnCbZNaFw==
`protect END_PROTECTED
