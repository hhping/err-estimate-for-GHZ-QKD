`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2dYYyNYy/T1EcOpRbxFkdlizeK9z7aM5GP4ForYi3Iyoioj14Adn1mpRNxxEmU+
RRa+ENrxDm+QkYMqKmve5bCSRtzhu4Asmh1sPKXdeI9LTiN9Fy1iBZQeo00PcEXd
08Y1kxkJbIADv73zFQU5dbhidkGsuN+P8EMYWPSXrqcV4fUg/8EkDpbsmyLOR4vN
NH3x8qDL2Qgb75YN8crmHE2Fa4bkiwOJDDLwdu8P5IQdbsqkRlUH32AlR5wq4vLW
OLlanhtTeQDDHwUQcjjQBo75PdY+go0rwJD+KFrgxl3jQ/7L08o/OcQaB4a7w59x
nC18uLuUiSY0WNFKnBeLeS8TZlxn2FKggjtmZ+t/t64+FfOZ+zDjxfCKTaKYVChr
zIQ4MjmqsQlcOR/b77jUJcaTsp7Boc8lKLrcwtMf1UbjtE5yLX2g5o77iTXJiXw8
myrBfJWEuxG6yfMtyhL0uc1XpX2POptkJ99x90Hs/96pC3ewJPyDOtP+luUHnEbz
2kI+jTLOow5R1+C6BT3mpWMm0ggSzOQd+1FA1W58b5yiYMcPNU3vNTzQfux8Z0ll
2FCKqsksKSg2BYMWEXMdyNQ6l4357qE2kD0Du22Y/IYKEcuGJUMy9yEnZ4PMrafI
naWtxLdmCnHS0u0yLf1toudXDaz0y8SNsJsgvB5N2mxZ4hfnA/vo77APu5AWniAh
bsABII65a3Bf1lTJ1zlPslyCe7b03ncbp89yARIpd9SJlsMdAt9PLtIJXUBgy7Lj
jeCIXCLIf0SMziEeqWkQqFjESaQ+wHmJjML60X2jhIvCRYuYwDlnV8yUER7w9Oxr
zK5Wf4uVu1DfkuxXDIIU/lK5njLzEN5rUIFK/dOezdls3bhNIBE2wU/ld/dCIiNe
Gx8zvWHVDqmKjBAwxw6/YjafP/sXrIaHonpVgRoIPMNaWVpNWcJViPUqGcyZ8E6C
9EK1kxfuT8w+xeQkOksWTsZ+PuoW1IEHKjv6bhV7yKKcHk4+YKK/lufVKD7VhCS6
5XozpvHnbK4jq/CCgR1OsRXxlQArMR54pc1zrysylDJk1Tl296SgePwzUCQaHvq7
HVQp74jxxNepIc6D9tm58TSbYHJ2pdgl8xduS0NSafaXaYnBahq1xaLLanJ1KTe8
pXdeTQnJL0rofN6kTW0rgEZc3kXUsp9xo3nZqzJv37v0G9kw1whxvJAMz5sr9h/U
wkzsPDBPjKZ0tRJtvE8ywQCXWTB3eMS5U+7zxtbfauVFIeSedw24Ctw9KIuA5xRT
L94EI+0ry8DSwzDF1VclRFt1VTADVImdMqW5PztX6SFkh/BTAKqN6yafMRXPJf8P
V9gnUvP8iHgvRn/d8Q71Qo5gvBGkiblIori1VLsily+g+3u0qRq/vgFgR0gjHPJE
KL4bbLJ5rtkKlwbFeJLu2RJepXcFEDBKMza+5ZNKYsBEQScLSqWcCn92hHg8RShr
XzuuySUyF3SIJeHycZf5//wcZ7ryGRiJjIroclIEwJo7uFnMYq2/HxarpaGIdUn0
7QyRQu2aHmXRZMlyMm5FM2D70o/YfID9g3/xYfPhbZFcvArhcY2C+q3Q2y3Dgo7j
pxXoCBA40Vw4yUV3GdsnY74C/3G4s43T8T5ZztMfNHU864Cd7gDE9ucVuurgoyk8
d254b3fGyES8iZReFcrb32JAHY55GYyDFSrBxw255q8/pmT3tgS0mc4bdhMOc0SS
DvoDxAye2WDoNdcryd9ZMeqTt0yuuPnGOcQOJkjH0Ey1BpdJd6cfWALopMlF//ga
j/pP15XA7JkT1RY0T71NgUvOYIv1zhWyXHxxFW3ErW9ffvvjhlBkPoeICzTStOsp
i76sKN3WHegtSOmilPXNSFSovUfeswFExzcgx9/kxgv5pKPcQFsEXEwpoXhmENZY
xiBDJyybhb5ZDCpPZ9Z5wzc/sJIBiadTt9NulMMc2xboWmrDYJArZvQaM0UtoV0m
AE60i8bMXtrSimv9Q27aliz87rdttf8JK1D0LjtO5UraR/3wY/YCKjHxqEbSilFF
qQyqR11EtBR/QhlQCm9e2NjZBc6f8ZszeXMMK61dJwz8I2QJ7IMbwsCNgwpXI5eQ
blhwnjaK9T5Ui6Kru/WoTlDp7+y7nUMeknZRkkSvGj657D1muAMrWj6WamTG8jDC
BWRlLPyGLK1u/2wpP7YrWCOmueDkYA9E7ZAEcs1i82BmvcUM5vp08ZkPukJcUxBK
aDvzusnA+c+Q45+i5lvot5EbXPCJRZJpF5URUvsWXr45+Bdo/9Yt1JJ2xd5vf0GA
bCVdB8U/wU6c4I2e4mKFJVOn4NCwmZWuwwexPQxQQrn0Uv+6JPtBPshESdmdNYMo
juTo+M1rs1iM2nwaxZredazd87hsokPuZoxMqCDqHGrKbouAINs0k/j+PvlIg9Zh
YE+dOYcdIG0CBk0qclTWgiCwSEg85hoZFDvlKuayisfEO5IMlWjaWHR63xxJ1Nrt
6qd2hfk3g+LssrnMmzwnNYKczpvzE6Mnew9GyJzU4oxNFpoZ9S5InuI8W9QocwV0
XMJB6uV3rZm/YoiUKBcNQJR79pkQXzV7r9lTUUdzsLXeZgUyZqdaFWbECcN8RQHa
KrVD3FcA9cSLKGb4Dc4zLpvr8A/CLwzW0miAyO68ncTkp8MyzU20h8dYxx32GJcc
symI3klki9INZnbQKZqPjB4GGynE098MlZDu3GRs5ExQp+ttM+Z/sULH2K9y6G4h
lMTVhupb1NMGOe5D+9asttgiXNwJ0q4NeqPcbq2afjlgEK6nVF8dlxF1x9BhNrCc
`protect END_PROTECTED
