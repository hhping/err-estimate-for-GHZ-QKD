`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zvFBC3giBDVmLafS91JGUSoiv3UbnwVk1QCG/cEf0HVZTt4OLaenQC7bx2apj2/8
p9LaZ0j0HwGeapzAhkiJf38XuDOPyuiOnbN4AUqlOCrwwT9KJwuZpYisQyN6uhh3
cSVxRECX5gPo+nILrTmN4G7g+hV5X8EofNGvLEkPoJ3igU2LwRkWGHMasSgpTpY/
J218rFVKriD/evFTLImuywAOGIWSxTm0RRS9IIiJm75mCqy6rM/6oTXV7bkz5eST
6qnO4KPa/PywZI+0xBNrxxc49EjLeQKaPGtNI5PuxLI0WtJm6+Rb5Er/VsDrReQl
CtqiTH0TGB3y54NigbtoGTnD/6cLbZidmocDE6l2ox2t9PLEAPjTWB5PThc56nOS
NRfTxRrxn0dgsAzV1rFwpCnCvdn619LbXYv978dBeuCNHqTefmkWSA8AcvYOKxIL
g8lfd+YSE7CTEOTqL+nhr2PmY2LHpz5VOgcpQJpnwTrvLfrejDFcBsMFMDpiYqw6
6Uwbalj1YFdMkuMSTD+QtVQtIUgmyKBkmaeKJ1x2C4/baMeFNQD2smCfiuHQPQ1y
sxRZvmdzQ8cgJkDcBMJpclJJx288MP6cKPnd7aIqhGzBBYo6hRDKWNGhnWLHn5HR
D7gMHi3V/6OdjFZ7vjPICJMbv8MO7ol3jfO7GWf6DOjs/A6PkUS1E6TmlMr2UqU4
ctoElABadWZpboEIjbh7iOmhI3TLMEesEmg0Gau0XLeXXBkKq39gMZLB6LllVRHh
ltb4fJIs1z5C1JgyZHm7k/dTQEaVhU/eU9rPIDaVjU0wWArhg7sshNygdwcD00Jb
pD1FoecFKEwqQ/TuRZ6WjoV0vmVuyzvkySt+sO1Cl34sc2speULKaJL9ma9TDEDh
5+mWJZdaA+MdpQLU7szPRWnmfVeHSm1tJHcfTZH/ZFkNdN6fOgVp+hdumHihm6PX
3d9ZBwm4Qfqa8DC0p2CNUbLOvAkVYZMSNlcAm8QRNPoHOxpaQwuLoDMjUrIJRD72
Z4P2TajTmkbnt+PNYddAm1aMTLCSJD3ssw6CuaIIFg15BGtSk4/mjQ9lX0D4DJuF
dimdVqT/QrdtjizNEJcs4NkYrGkLYhLSLCj/j1XIKg+/YwwBt7JVzqvP4pJgMWWC
kWr6cKbQY1Q8CUt16HakvolGsaiKuPcFSH4F0ZYFQ5W/bjdE/S0rzfyujoTqtUcF
25XFgk3f3R1bPIUi8wcioXoZuivW3s7SaM9nVg01asI6swPkn7rSdm5Z1g3FnTBY
9gfsfLgjWpkwUvhwL0D84Qu0meu2d8swh3UVOByMtE+MzEQKkwdne28OeAnk+AV5
Tf2pL5JIPMkQsVyyHnJ/Tp4lrWmgZXuIUf9Q15ExCet9P46vfIovw5isA2JFNOSS
O1w6iy5wQAH+3uj80RFSAAKqEhcuuKrurCpveB2tg+hhZF09lyHtMFk37x8GDblq
1oUMjIYvYMYdybvymbBSDNgadwgWFErMv4Xd7lgc2FzqMOl7rOJXbPsyrof9ujcj
KHH+8mbYIsYozjJcBgZnrdLMmcd0VrZPFDBw3ym2A7r2cbBwcr7R4eJ7883TuPbv
r71Cd+3FUtWCziXegmSAgUrENNVpjuhkDE3NAebY6aF1EdL2DuK0oHN6iLp0zaxX
adVxGLe3kyBEPHmhIaLQItII58WwqLhRC4bi6T1NQeEvSHv9k7/XBA4PxxsPtYAF
ahCkwXuTBtbfTeCbuWx62rbu997gpKS6UZNthI7lu/F4U2Tmjs6X2yMx3UlXXnjm
FeTWqLPz31I5cGstyd6IT3FbE7kOGXcA89OpuRCC2Ohje1vvhUhvwD/Q6VziAquF
DhouS2hPvZ6e5zR2dNpKGN1pMMgWTj8p24SzxIsut2A1VHsu2q/P8lFKKZzoeoCG
kPWrJYtU6dvaMbUtRboFHGtdireiu0kOc2nOLHpgPug=
`protect END_PROTECTED
