`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3+PraoDdtm8C3QaQ2KmOys/m08wPuxBunMMOoQVeXxjJFvRkwnBgL//jfBWMtxI
NodzG8c4IQKFBoj0kUZvNdYMPGx210n4pyOo9GeVyy3rD/flcHclSQ8uTrhTeqNf
Ol54uVG1IQS1dQt5IrNrOjyuLbgFTJ2QKOt6M7YfhsuvIYwqra0K6pH7NP1LwUgX
1npD2JwuhDEU1YxFOS1EyuPC3cUOlbB3GWweC1hfDWwT5veW3Rxj7DOi1BbD8t7z
cveFEApTrKsQiERq97fwupXiJEnTgIKalWc23XJHx76mXt522pCvwh8kJW3tNZlr
mgYuUH+zTey4wx9yE8oR59KoiJOs+FsFRRL2sfPLdCW0Jft8SYtzRtwS8X/qsD2t
fe9eE6dR0FRJt1eZakSZaaqYnVxtt4f4tDo2qcTc1LqFftwLqxeOlkutQah+RSwB
8Q7xFT00YAbevMu1wZBUuSXc0ZMFPJVBbxdNCy9sWXVvFXWIFEGhyuUfKv0dnati
GDG9aSNbuEFQURsUeOibVN+EmIpAFnXTHDa4rgEPqymxy/PbKKC3aInv+hOKPg+I
pyU+DF2+cUE4nHno6PZ/1xrwQMSZOCWLa4pqhx/rghFFqZPCBsdKNL9zqPIZCume
3iyVWJqpExFaBDL4W7PNbsAFQ0dNTRDvUKV3IKyxLdF5rlq0Tb3UIYUjh5p5XehL
9YXFoqJlKwRR18x17CV62qEe8jsNh2ZHzI3xnS4b4LXnrbvP+dwlGq1YeaJOvDUm
kquWugwHOcmRFjOF3K2Qpq2sYZQ3StlMC+/t5eGyyV6FGqPrho5kK86HsnkHeis+
+X8qSONJdQRyHyiWSiEufc2DOaz983GFVZLH5p4zWeJudZ74FbUsfVzwsmH4dBZG
jcBKVp+jjBoCzqRjk2PrFD9EH69IT7Q6Ve2LijZ4XC2yD3mV7bm8GWahVI/riVmu
xzuDHDHenEpo5SXCS6Ydd/SNtX8bfYQvZM/1zTj/lb7uCHm+AGl8S8lC7AYPyxkN
yPJE0SBj3yHFFCjQAflqXgbH8ggAvZbzzsGBc196Ik1H1vPiXTxM9zSgvldNKoJo
rufawSJFgzFuylttQB3R1B7/nF2TPqsm2n7p9js341Va0tBULpmeC/0qVEl52nMK
8XSY9Jvl/DwxNBYzfwc6ikyyHigvqjdGBK8yBjwpcbMnaagFmzg9tdpLRmDSLk6U
TY+krukkdJb/egzex8j7FFVHeLpW/aZLqHG+VTXFd964fqMYxfnPZR23cvCO4vhT
mMEaeRmN+wIHX9eMokcB9NW934KEMwZEC8gPbPMnt7zCg7MQIM+4VtbRFLZyhlJY
838Tjrir4HJWSaOKjEgBeV2ZpXYziHpKNvhlDsCYYo0clKzfne5D3gWT8Aiju6Uz
kXeAApIed+sSwdi63jxGCIUcU0oIzKi/bBYFLdhl1Y0XvMudXVfa42KsMWJYJRep
oG4g3eeLOMaX1UBF9fP/7unnkLBxSqj8ffy6boONTEd1nb/YOESqwPC6VlR/NO0J
Za9vsVYNoa5hjozxFD4V569f6NulM1fyEGghMa8vWiOUIyv4JSOTkchFwTaRHEeU
sPbMNitwV8VXaEjghgokw9azhYKPwg7U4+5RRPdLZss13ff66aqc0HK4sdjC6A6o
j2kTKv/vQblosngfSCRaSNpJJIAeKI3tGxkTDBEh1xlp94+N3ZcLmzenLounfJLC
Oja0M+FuSGTSVlRLiajSdsZpEenqdBVDPcwwGr5TpuLRszuhSNvJC34YBTDoRX9E
CYddebWW4BBpmXP0BewkxFS6zJR0vx7LOwyNA8YpiHKg0mF2K6LcESI3CAauSu64
yloBrhcn3SDagz07qD+OozqVE3wh+9qebLHxe5q6PvlbUMI3D6BvaiTRbERBWZj4
oMHkGnVznOik1LGR1eIfEpuCWWa4wjcQ87QpFlT6HVliQj4HpU4incNJW5hPqBXa
5hq5L8QeyDlHgXh5JN2a8W4gniYytj1+vAUnUl9TkBOYpF1dKsetAT5XaYM2Jp0J
bckEbFRgSOkphFbofnGhm6aRW+qCuep5KZhMJIsgW4HyiYAfzIOG/FqImtZJwTKz
pVrWY+25l4Vep5K2/9922s9rNYbdQYYm5TqXGZtUju/Sqed6zy+5p/GjXSEhwDM7
vACPV0jdDq1p803OuiGXqb7/R9F0FNVxkGIu8DdWQro98nNI1+QLy/srWJyjpiFe
qOfGM/odmTnYeYjSxtC00Vzxi2TfK9iR3BMEg3K5rB7WZuKWuD14hV9KIO6uL5pL
Y28VuQX6hS7z9d9QCt7Tm+fAc95hPdxcOIZq/+e0XGMXxv0WZIUp/eZpOZAE2Tdk
GbwJurkvtjYs5En9uIKXf5XbK0qIbTtcX51i/ZBKfoZE5p+8ewnflrd4eBu6evS8
qX6Qgf4+zjXtMqfx6dBgIGhPd5xORIgpjtZShCCmE6w0KMx6R7E3vThHuMktYpXj
cUftDGy3MxxY/Xb3t7bKTXGvejev+zoALtTSDzmuy7l8r/kHC3Z8smNXSocxiVW8
zPuJIBZVnbDKIvk38McC/Yq+RyIaeSATyulFHRdeim0OLWWBPIb0GPA0N70Y4LIw
G8I9Tzemb+4THY7+pV+gye54g0y+P59Obuyhnrjti2dgU+C3YDvx9pxf4lVV9tz6
VIepIbgAevduRzW3JuKFv2r12dp135vrXxniljKzXIQVC2z1icSUbhPX7avLnGyd
8CoP/S6v6kOTh7t1h8Xta8D7XMtM2D9rJ6TgeC5LFNlsRf0BdlBhsHHxlkgAYZMQ
ciq9X8vOtOylG+lDT26r/cIbNMYGorkTiZQjU6+aUWJKOLzYClXmYeeD4UuQzLOC
3RUOiG/h00eoInxl6LwmYvRfacFMYwk6ueyUCQKJA4y01/nQ3niH6W559QhLEiC7
g0yplG3yElzQzzO2xvsXhxTpqYCNcNLQCI4scASR+MDHo8qUCy2LYmZuNJgQH1oh
e8fQK6hWc/FggwfxCZRvmOUN3PhIacBGfxycIAeQJ2PnxdRqgE/I7Xp7u5zG53/n
cEIITxDoi3I7qng4CA/9UYEySIaJxXDYcuzVP4Iek9rK3nN/VABiQO9KhtPVcv0w
fsK9c+1fXBaTiyt9lq72F0lt6UNZwkn+C2H4S9ewvve2L7bruPECfuuF++i8ODSO
ILEt6NofaA4yllRQjZd+mO/FOboPlmeXXifVg3zs9GZhJaaIIPki4PBI5/0SMKc9
sK8eJrBmPxQHhxS3VDJaGSSucm2E1fq9k69efkpujHBzn7cs4vBd5e6/z9S1I48F
EmF256U2Y/TLa/fCf0u9q1MP0LqD8asizlBlZTPmF2wRek5CMuuWYRxU1+QPSBYb
wYYJs99JqvvqN9GmWqQzpz6rUXBDbB2wpi7L4nksYm09sQ+B/fVcbyz2XuJGV3Nn
Wne9CZLEY6OrowF5GQ45ilydG4Y/IsKZbUNoCY7I25wFmHSONACvAns/VYsimAup
lXlfYnY9L14dFcqNTSjZJ3I9RiJokPd+IXI747YQeHZTvU9ud7N5I3O9ffdWPhN4
Mz8rnNUaE08qlqMMqTHwwGdioSrYltoPYfzY4fXjqb10b+Pkb+q4RB1Ir5enxYNC
Q8PM81cQyTMZU9TQx8J6PUOuNZpuAY28icoEa5xqT0XL+LaTTkV9xqvXxYTfqo1R
J8bcAVpac+lJSEAKJs1o6qVEd7v+qcBsAYyA2rvWBvyfH2CFhr+LwpS4mKqFFAUI
dHt7+p7onUhAV5tUFISs05dT2zxUSnRPvpte4RrWL6wBVajTcgw47vcrmG2VTqWX
bFDK6Ae3kufOPdjXxlM22QjzcG+sVyQL6Qcvqix6iVGnfaT7oFT+Pi1pcFbzwHo0
MB8CeL4TlImzhq9ZKKK26c+laF954Oga/LlVmqXyqwY=
`protect END_PROTECTED
