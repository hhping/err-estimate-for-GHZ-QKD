`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybfEBvlqo9npzp67AC68rxLkpNzK7TAOH8xFcWoT/9LPEf1OjnAjpPXxZv9t0f6z
P9IaiyBIlZ1Z85wikNtVgcJ2ylPH/EFKdnuq1kkCTMvkDBRP1hdBk4dBtldN1dUO
3jaKNPReWklBh36WdGd3yDENjLzrx0Yb2arIHHu34pJUpFX1Awx3aUV5awaDI2i+
vTFwgY4UgVYd2plqUqteSOcIto2DW8/8+GzUEuFoWAPIxfkcjqpZH3bUkgUPxilL
yqhAGe1F4bIrgeIo1AffY8CJOxDxJHsHgHjgpCepMhdJXCg97hJ/WAi1CYl0dr15
Zv7aGxQQdem4Ft6HbsBWi2Ou24+Mo+zbdLumrkqMKwWVtb9fWP9lwWKl+KUwQSWx
/Cl9QqR2JU+w7zr+2TBi3fn7b+wnF0oFH0gnG8zQLaGtAT+kdN/5/Uns7QbI4/MU
4SYLEY59SScJwQxBmOEGWxUYN32iGhfzoITwogNY1AYpJINYcQzZQzZPJfn8Qkw2
Acw1ot+r8F9Ysn/zLqkEYvSjbALCYMQFQ2n+jFnid/V2Yefs9HpeQJlYIjOJnhfI
7p3iaLHGHR+o/xbFj9AfGEz/74Lac35W2bOG/6o/FJXjMI1h7AYjPkgKUl/DLIqe
n89C6g7nM0u/LLH5tdifiJxWIP2H+gFtIkQ8+JiPJTd4g+Xj/1S1iU0vt9GplMFi
iinXbWGRwoyNKU6FzRSWyxvFuMR8yvGksfF40UlhHVZrueSoLto1DJg0dhFVrtPl
gdvQDqNc3RlZhpXrPJagCaz/46W5haVqVK5u3ii2ryvSYkVm0o5n1JEBt/SyELX1
`protect END_PROTECTED
