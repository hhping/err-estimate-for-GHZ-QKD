`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGexh28e2YgLOp6dQsJWAkQ6/xW2ZO5432mQQavsHHfmrd+o5MUfTInt+QdYzsO3
r6DCkFC6hZXPDNYRhRWFADA+01F4QkjPuNSFYDNgr7EkLjxbfVj2Y5g8/OXDGRaA
PlGUWBJPtR2+AGGDmyuiUBdlbz+QkotYdy4ObPg7uE8kzzuIs1JXq4LMlhCD2gSu
iOxHPTu/ZmjWkBnnIg6MPIKEiq4VPo174ntU60J9nP7BUULHhaC8Q9dy3gwN88Je
1182FMl/AJM89sUBVXX73JBkYlcqK9dUUVLA850AHviqC96I31OBP+i4gym3wtP6
fE9RFXgg8W+3gCSWiuWznbpBML2AkDLmSw6UBcaX9gc2fyXuOpo0y2AZEN1tQzIk
nNq/I5TDi1Kgmo7/AwoKjJr1IpvYZnxjiMNyuf30Ac9uZKLlYSYpFI0zFxhY6XK7
kvjnX5iF3qYvAqlWp60qvTo1GmWuq+AhFgpNJuBGME0BTipZhtZoywH+P2E8jm33
3jHncsxGDZKbXq0D0nejv9nlwbrN19SliUbUxSGXX6sDQZl8zPn9mwShlWodui2g
zUr7Pb2IpR3zRQLSIF0Qkfq5q+CgELAmimHECj55YTBSEkMsqPmSMRrfe1V794ix
YLYCF3Ab5DMkrWW9j6FfqUU7xkwN8btUt62fWPvKYhPGkPVuiOWUAg3P8h8sjASH
PQEjpqKpTgaUEG5mDpPxghABGgisV8UPWdRIvcKLZADpEaLsGZtYOsTgS2E11HIp
r2MMwjCvamHy+8PVF0fo2hU21Hc4X1HZmO+1+BVEkfgwk1O0mzyHeRqAroAP+oc+
8jBuX06kqkow5u5KqN+W11GUZBjKGVbfGers4JW2tL3J9FJs5JQB+ljL4cWgWZ55
hv9whsXcZJGQLkO6bD8VQykoAXxNS7Ieb6JqNzbvCQNCg50d0W6AugEFkDzLy2mG
Lh6Cv3EnhEplFgDoA0Q4Mdqx+A5QhLMj1TDuR+6HjN7UoaThU855fKqtnhf4ZiCn
psG5DlsO0WG9ruSwf6W2qSA8cdlrF7zE4Xe9zv4EwB0Ni8I54KMqxcPAsbHqFLYL
Esr7qQt+NC4cO0tptEuXFZ32LmfBpNnLhlA8J24QHprHwjBrUBBhgnGu/4mnmheR
czDhxuSKPddwxcJ7x+LVUsbjNfzQPA9tj1w+6ESEWKLN6nQeXxuuPZgPwxIeJxoz
lvYj+bgOONIVhoKz/bPmHyGPlUG+MrSpMVefxDI7OIPXuiOhsPaueiC9ihMFk/oQ
9fp4NnhxX+9l9ZVNrsrn3Hn6Gh7eo2B6JuRzWoryqqu9cLGlzXnEbQK2W9H3Sr6Y
KUTw0KgxugunUHKXmwqN46lqBXDVMdyKey0G6RBGhnVk1pn0BFwDzBQuRYV1YVWR
LIRyKfUAA12ZoDN6yAW45flwGqU40T7CrmZugJWxXAREWJLYhcXJ06Aw2i2VNlUC
pJpOaLaJ2zjhLcnMZntvwcGhPU/c6DDO9BMuwGY3brBWv/G3tqxrScQsXcQug49k
rru1EdYjhkPaSBaaIJoBKWqKovMEx/BC6GBv1L2lEpaLtvj0FEXpQtYBvz3R2gFR
COq9C2rfSm0UD2LV7I6PTE25Y3OaPgTMTUT6Lzk0kSsvsc8/4SqkOAx1yonLfKOU
HpmHiMTRZw4nrUChbfZufw==
`protect END_PROTECTED
