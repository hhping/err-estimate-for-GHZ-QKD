`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2K9UpcFm2oupxLoGF5NQ+TFrEVx/fhVF/O/qfjDlCKPhe1zNshPFHnpBDFFQsEcx
X2KjBzcvIS45vHNlY5PYQZ/gUEsU/hYpXmD5kZzFkVGb50qkFJK/iPlFXVUBbamG
XtUmDAOYd/H4V7kuECFhB93wKsf8tC1a/TV8n0QBXsJqaUxlhipXm4oexqNHPUOy
bW/rFlMoXyzXnbb+y8w7SmkDW0vBaVzQfzXAVqysAxxBQQIFZ9nvwkyO0egndq1r
Ncd5EjdI0NYbhCSwLGDQhQAXGk6ZcsTFrq93AOBTMRyCLRamQ6Zz22nX4gOOHvgu
j9fwCLU1qK+bXrVdnmDDzrZluUm4GLnz6+Yl0+fFH3ZIbKw4amO+3OZGawE+bjPI
8+5ojUdZQllz5S5MgPURDbLpa6z5G+BjzQNMT4/GftzSrFnww3LMpkx50vAnIkfg
5nG2PfrvE/rF62M8IoN6gsjAdeHiNo1PDQhRckAGLwh5C0QLDn9Tu/EjPDrLNR7f
XBAc/EV1t1f473xgr27Q4g==
`protect END_PROTECTED
