`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KWF45WGDUFGT+J+WX//2mihAUZf6bvVMuncJQVH442S3M851ly1O69MEHScq0em7
0SNnBUfF6oRSE2fHIllXf3BFGIL5uMhC/KJqVfmd/NQA9UgKxgoIssZJ3hjZNjWP
Ebvh0uikWO6u2MGusjGsS5auhV0OKV2W0SoLiV4/xOMIxVzIX5I5FuQtFtNnarzd
o3jY29V6198DsS+SLv3F28/METW4sEyTQELEPrrY+Opll4+UblyAGb+rgzKPlSiT
VQAkEKh69MxfMc6qG+Mpn6g7cR+FDWjzQmABLm9FxER1mJaVKWKVAyMZAT0qdRuB
/hLbWRxDDel2EZMsQfJvbLksRJO12FFrYlro8aGaBcx2nd/5vrXUSpfgrRG0ylov
fB1lcovqStP7QPW3b6+/w/yVvXhebB7onFt0X1DOi24XLhBbSr2qKvHlXH5Ljjo0
un+Y+Cc6Xug14vYuh0UMmBSIsr2DoSUBnVkOi9pQlZA=
`protect END_PROTECTED
