`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+EkGBR1Pa5F4/wWjxMCmVeTCABJQnSDSw0GbxfCLhmMMUg8kqv0DCT/+XBlHqfy
URMWwOBYbhFmX6smolunmwRHnLEzyobSOKReF0PVIADKzAlCPDVFNJnFJfHNZhSh
UTPvEO51sbFIAHVv5Qc71lE3xhlnwlLr8frE3hcPLM8IE82Iavzbbmi9GOdC6ElJ
s7Abq2eMvv5hLIieiCmnN4+q9XKDLxBCsajAx7cN7Ti1080k8+7+t9CEN6H8/Dex
IGdgs8rJVkk7p4GUXqS0MUnyOnMVIPWnYyQoyDsmSbjuwvqiyXb8VTSE/6YkvZZR
twKuMivmrsRIZL2Eon0kiHVL0xwWGyENOZuN+JrM4klGIaV+t81XcSPrWitLG6cH
gzNHw2h7fYrnzyW8VXlRirkWozC06mYtlyAZZpND6kYtvJb+0AVJ3i7ijrffuDG5
32exfqB3Hz9IHjnY2xevpsNxtdOadJrR/A7tVH60omoUsaGZ+Jw3H0hnXDDDz5CZ
ViGNIHe/ADo94p2YU/Olds9Eu/8gIjVLwElRX9Ox2V5b9saHFcodQbttJjNCYz5c
zjRJAK9dZ2A0RHhLqtrGfpkguSCqhR4qqM2YhKp0SLjGqO8oPWGNA1fiqNPyFy0k
rw5wfieE4JRZx8EBq4VfGWgIqwfNdH1X/tgMHVxVOSFC2yy5YLLBtUxpNqQAexDS
CDZ1sWLKuLqvz3Lora+P6Y3xiRy3Ncpvg5wnOHe8a0bbfT8qdX0JzLzT2TkAcfuD
khwLgzIATYiAE53geUiA3kgKFVbVBq2JfD791UFgNGpOfYxwjBs+jurc6mJ/KxwL
f2y2q0PktZ4818jCV6YyzOEEe6KSnd7XAKM9rg89z1FoqlJucWDsCnAsasIQ5GqE
hdQ/lySDGbZauc8CyOalrCkTx2SZ9HiUF25lI5byccXA2rpfNJWV7++Q/ifgVqL4
m6qnF87FX5XdtAzimN/2kPuzavlLiuNMKm+opgFmDG+AWrm6zsFdFfPWpleo6PEz
X8crcKUxHa+zMVrTW4jK40gXnFcbJNJPVdPhs5Mo4SvXSnpSZdS0tlH8TYJPqrFX
K5468CJi8hm2w90Et+ruCnH7gRQLrtFSq98D4E/ii1W5rUl83VvIO3inlShKTcv+
34sipZCuWoj5Fc8rC7UnJ1FznW8gu9cizfPobFX+sFwhbw3n8lez7GQ8ESdd3mp1
cxYdsc5pgNnnhWTwKYna5I9R0PjxrVX/zRNr9In8spiJtCS2I0mXqx5R7EfOfKRH
zd6RtV68tw/svuTJ8UkoiNBq7qwIBDKdI0x3vHVVMeHv8/jO/aG4JDowdxOn1coI
BiM71RHKkcXw2KZt69qIhGXZ3UXqPkcWrsuUX+wXOsCj89ejvwHjoiwHkws5i7sS
duYePm2GYOK8QSC4Be/l/1gH2oVd0xhXB+hketSnqhKjT5M5zx2ZUyyPjsalPbgb
JiRfkxZwgAFJN/M+4kqzxxOVOc5NYnd9rqUL1RAxyw0fWM8oKzHTj2j6ytnFggWo
NhYlXON/BqyPkbdx2wuXegsuqkOCtJG50ymEf36X1n+dYUJFiXkusSpENelfG0kg
Yis6G81NAH61nrcdbro7BVcOG1TTvfr1WomLFdxMe9qVQegT8hju0pH/mUH7F/yj
XQugrRrujeJ79NdRHxk3hC0OSEGCclmjrUSuNb8xsjU=
`protect END_PROTECTED
