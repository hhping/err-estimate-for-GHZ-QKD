`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dPx2eLmd3gE6/w6hGsow1Bo8mUV3e2ofCVG77+y8KuuX4Doz+CoHVSz7cgYOkDm3
OWw0RTR00fmqmlC8GC1odKdsYtrZTrDL6PQjeaTylUqSFkrIb4gjQkI3bNIwr3s1
aLMbofrmfc6IXBGkw0FB1MZ7gPay4Q/hAcwI30RKbxRxM2ku4dZxGJmbjpl9GaJm
WCkUaCSeq+YvJ8mTktag6/ZKUwBSRwVGoIG4RSKsNYo5jw+ozzSPi4YkzohPbMr4
SMNnvrwUyvlfefT7ELuxKKbJau9+TvwkSewiIVekYh/W2DsTZBJ66HmH8PqtyyVe
YQhJkpJGM/WE5OqJ10xP88FedI4axxUZ2xTALIwu6uODb5DtCo2BkN7mBv3ci3rz
n/mdNPCvAtgGkCDOsouIhSauoNO7GV+zzXc8FOveWEboeCdnXAIpT+LbwoOt5hHG
iyU09D9Q+hqIPVAdlYntvMkmqvZXK1D93XiF8XxsV70v8hdjRozFp/vb50m3cOTw
1i8ny5UY23QvJX7tCC9AQGDT374Ac0Q+i6Gu5c5oDvxCqx43c8Pbi4Ub8HtSV41U
EibDi+POxpO5ltJhfFAdVQrLTz/+pKETD/ErEA3k/PqQ7PGofIlKG1mL0ZLoxI1d
TjkFlWeS4LQOdBVa19ggtOlBOT2efL/8ITsSxlSqpgRn2w8R+bqdxk+9EhJhLXdy
hCp31o66GvPwkszWgh6Aoene7B+6Yhp2dZIMs2QqnqhK3+Dz1lw35WZhrwTyasJe
7vZIk5Iqa2wP4oY5necvK7mWx5yPsK9acP9n0+0hM5Um59o9Bf7aaSPEx4ufZaNK
L6hBeHRtfr2FIMYw0ntjlwYNVtj2JCUYZjn2GU2RkrmcrquxYBCKsEOmLQA3YOxm
8ox0Jw1Jy9L8oTkq6SwG1gkwtdIgxoIbNvJSilmPWkLzHzPpAWoVd6dZyc4E0E44
K4J9VMFscoLLMG2VakvTZZyzo9q88lUPUyZYSsGPljYd4Uc2nkgYojy5fxcyiCJz
+l0/hYuLpg0yma76/vwANyha8Ehr/LsIPINa1xligVVYUlpH2umSkOLd5M5rCZEd
kPwMELh4U9wZ/XUMpboSYTI/N2hZecvtsOtxslG6UhKCtQGy3C7ye+mMp8z749RB
+8sb3lK/DzizDPg2n9LyeuIrSlGiL1PGwX8YWGlSModD8igWL2MTfEI6zin45sYi
NPKxDe0NqiyRG4HNONHPSPEpruxeUQDIYLjAxJGXp4u9PuugrODUXuaRqJd68cek
xYQnFXwstEPjlut+sUh3GpKO6T5KzMtnP5jR404znbjBBByb3rHxqEcPPEB/0rBN
nT78YpOdHvxJdYAyPxrykhhf6MqYbnWAWpkIyo7XJiq9ggYvO3MCuAzTX8UKBVyz
lNyaN0daxmSBUX+4mWGcu5bY2Z+enexK9MEoLfho+ICfh9BsTxalg1hSxmItyB6B
SXugCjUl+2o6JNZfN28cOSGTbYQ1kGH5OWKn1DyUrn++VLIGcs12eapHrKXJmjFs
EUpWr5q0jC2arZgnwpLSjn2npxtzkXrArQ0w8MNc458af9boKWdMUu5ydlCmnFBh
CburLfcNhVtPERK9dQA5HJTjpJ/AsoetuHQQftNznsBpFYTUxuKjx2ZH/k/wdtcW
Ep04UW0X7LUJWtuWgdoZjaXWd7lOLnr6yFaqYXOjMmZiAbrIlSbhC/E0Trzll6Ue
hoU8Bty4o2RIDhImDF2/1fOe3S1YlxSt8rYOUMIUDCZo5m6B88DQBf9FSh9OtP50
9d7QtzI8FtBMkmoTZniagJaw0bxuUpHo8wyQipCi0YVB2jAb9XonsqfId4kjGtV5
5A+e516UHwf4aELBneQ31U6f2d3VtwkGmY8oc9KQ1PRp6qiYA2DP1pPhGBSR2FL0
2ube9SixCDxyQ9B+/duMtEFaa2a61OGZOtjF3twpW9RxxfA71rSiqUxInGfIlrsS
SLPufcPKfxIbmsVKoVyqod94XKZ8BkWoU8M4sy/vmM4+MnrdWEIDP8/wAEG3BsnL
o37xMOXh5GLd1KezxeChBQW+SFDTPOOQ4VkMzSbi9vqRNo0dnmLKvU86Xi5MxSPk
IgLFHIVCqKSDYcvXPWnR7vnVM4BbsPD+8Rp2uang5MYy47CBauNE6uE4I5mX74LJ
GhZmo+/yzGgcdeVBsn9HiPE0YzVmSEOquB2Rs1baTM0/Htsh6DKmGWcnBP/GiasI
y8LPl5ud9qc88lESvVDvfRArDdCNuamjxovoRo3EDAZmNwFlPBSpPS1rHxUagkG1
avdBhrZFtrFEC7RYCQUG/pyvzI4UFR1/B6gy81G6TIusqwhf0nsQS0E5OqVyyiti
r3ptWI7sGHuCA2fqNniML6LdDXes2lC3Dn6+xoFFZU0HhJhVoLR0xoDevtXYx4k3
nkeOxNTlpDVNGAqvLXnIyL2S6RpM+7UxnmpGSUDpa3NSUd7/vFb4An/2HP58jL94
DKNZ5peWuatVtk6RD2utS9V+XxphNJB53EX010MXNw21b4xEdaztYR3+ihamuCVS
WACjTd38+RxzjN5h3RuRYiP5MEfKLnmvarG0YG7hBqSL7ATZsdQ1ZSeAeghgamNj
WxVFwK3vCzNX/tFcKP8Sig+fFDA8Z3eKz/ipZsnTqtbupHRVNzVkzycUInS1+1QU
5vaRIMPZuqxkZOD1Ih0n/f6uzlEKfacOCAqsQPV698g784hkKN+QCZ09zhO8g13a
z0/6ZafKvpJeWee873POKq3aRbuFiuTgjyc4aW5XaPa3FnpO3QyduT95NWflxoe2
Q0lGy66jcqVZudgVHUnoO8ShQkFTxjqTFYDMHAPc2ZmoS7lG3eDcXitrQweByAn4
8JblPH/mpwkzX5FlV42Kkf89Y913eEK0n3thOigvWMFN/Gcnb6a5c0SRdGuWhQUP
iO4iBwXy6APQwuJIqvR7Ba/W2nk3EX0Dar9K+FOT7wGsLEUa5JCj8ZH6QYl9ZCFf
BltRFuUQB7RX8k2IvnF4c0r65e5/2r1fWu279GxitiFddSivudzFiBPT5iBgxIXj
SDv/FMk9Ex/rDcPh9LP9/DvnII+Mk2C+tozW8n3sTHHfyW8TZgh+bfh1Bleckm7u
BfW6R8++K+zcYoCSEErhBFZ6ht9Zci1RNRam9LWhsnh52GTbDTriBZQDJ6Ncmy/Y
8F21fLIxhs80Fs3uS4u302jY9UXpNrdeErpRjhPtFX9SO/hdQm4U5P4Mz31kmJwz
avFXD7Z5GN4U40KDrMhjz0Fjo1+FryiW8NQ9CY4YJFZ/wQNKex7kVM8cuZKhxxMM
04S1kmIfWH6zlAw56hfAOyzRq3BzKxmLdHjODzur7XJBaV49364wuK0rWtQufPHr
J6tGOZGy/Bn4wv3GiUo/TAI25SSkqXk/NieZY/S+PdZSy8k5vyGAEjt5ZWSbQrc+
rLY2XBt3AGl6GtqtKyOs6tEtArOhIKTWRQivkfuTI0mBk+p/RUIk5+nDQo7o0T01
JpvYrRLSWukmHlixl34wytSGlxfe/dASha2quiJgwGdGJygAFOPa7fE2S6AvvmQ6
asajwlS2ei9T8+Xun+cONnCB9tWUOplvcy5SDHOE8RcHgqnw9HZrqUIjRcToFTJd
h7+asmZ7Vfl569JQ3QszKn12Yvmf00QEhNtx1e7jcEsMqyUbpq/madnsIpkoLLCX
hcr2LHx/w3zusDi9uK1D3fBT+bkP9+RQha6L8gTQmG2MUGtsVLS7nctMxVFvoiNT
2A0AcSwKrdPOH4GurvxmSYH8IvpOURRDhkz2WFkSBUm9fRO0pyY1TG33YihXL4Rz
4bdJpkU7u1jSLlOQR+9bvW1vGnIxR2O2ZevE/JFQWoEgW+h8HX8neI605iI2VOmb
EInj+79+RyxWHz0yb4ZtJQ==
`protect END_PROTECTED
