`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sdymre78iJID0JncJB/x7fIWdpiblN+/3ZCn2J2onuVBBfZ9UdNtO285w3hkAh2w
PtCXoJ+mG6YDQ7iYInlJuL7/i9YSQE8wDlwwI6rPO7Tas3twnXNAJO90VtT0ntBG
PIfJSa3IBdZhz8LWMtZbw7oKUEeq8j82KkJASSScrFgirwE5zvX+NQvPcKSTNo7D
gPX8QfgZad+f2yHqitUNJK8tRmmrnZ7UcxGLWYf++1pbeSOoQblU6No9v9ZD1jNA
8tJMARIaVxZSjN2A0aO0P6thqlwdEHuWVZKdz2Eh2MNDck1t41xz9sWX+oxb98vz
luH3GbvCDQP4MPeZAkl7genkdzfgVVRiNX4S4KLBK1SumhhPDbXcFwes2n6V1uBz
4XPh6YDpx1uihcfogtVHNm2Lnyzq22mRKwRyLLC5J5omGIb+V9gN2ZQlQHBv5/Td
oEGSpK5vP4cHaatCbHNoVe107GLM1xn6msmgyrmXpM1v5hj/8kwHvsMiBgAybVj1
JsCtBl8nFkEf9sD7qcFEkG2oSSwgcReZfP9LDWopDrIQsRxoq8/5HDklu1xw5jnG
51Ah39nybFqPZ82lLHl9XbdVETcVxKnXSi5aFWNtEdDUS1YLgVcWBmR+ZSUbMGj0
ray1UbKsJ0F8Yq6AKkKem9sUrPaxVP32/97hYuY08SkqkAKgehaFIxbF6iVcO/+R
nF89M4htTRZOnZdcFLxvBy8v5bPR62Ip/6nhVGaSdMtYwF5TwAUspIv99WGR6eSY
SVCEZ1/q6vMpMwCnykC9mu48clN2x+YoP1rIifi4fChGjh8BB9Mwhr6o3J12HiWK
zSAalta9ImiVWAv/u5PdlesfGlj3OrOgZzJVod0Ycewscpt2CDgTGcPCdIT2iMiP
`protect END_PROTECTED
