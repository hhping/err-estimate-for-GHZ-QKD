`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SXByqKtckHqoVRVr0HIDTe0stn0S7B8KKTqGnY07PkaR46CEdiaeMP1xjEf8Q8M
Lteh1KvUtCe+X8gsAkOfhgOuwnyrgXUemLgALv7WdsDUH6gdBURRIArgdcxHgL8X
rZw866s4y4hPp6894TI/J2kip4V97G7bWC2eLVj+Jh49htSIqCZ/NL18KzyOyszD
O4Xgu8CSNzvZUScnCxq7QfKhDgnf4K0lgUaq+yMnn8j1S0SmTG9yPZSEQzF/Hgv4
VIbXDAlLfx+qU5NUHWXpSeCyvUiQxozcyUCiD8MYe3WX2RziT2aeGtycQeQbWjZB
37BREEkYaTd73cxDzo/vSlGdhlebq6qXvfgpEoArRG9VeyOiaou7s1f8nvCfgCo0
epG/oUb+Brd174T9E6pagxUMvqz1pjd3UMCgPvqXsXyDuJGvJkR6wXGBqq2eW78Z
uZnX/9kTXeBIGeSsMx/FwEFoXsnHSehhlzaBAD25Q95TCvOAUaN2upeyaZwY2yze
RngM8f6uv5qSA6vTiM9OUxH+skAC+wj4F4kR+awmhtMDdADEwENxDUXDG96498XH
BEtIahVT7PzTkC0/y91CGprZNjyWwDFa5llgw8nXwqOG4ZYpi8nPf7Co8mNV4DKm
J/kD7ShemD5PbKBo0Eb009p8FZYpMMoRHdTrkAAW+yM=
`protect END_PROTECTED
