`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKapR28F+OGA+tpTmdcx2Waw4icnkx9lTnxgHe2r/1eSwGe1e0WB8looDniVRfAC
7TtdyzVCNIL2pb3GY6nuo5oA9mXF/CuKg4jDZE90quze5ZzoTIbJpS7Um8/G5JIg
puluvwUG7PrfcqEpGVYQ72/P0901M99fazMb0BmT0jxzI15zks9ONtUN5moBwo2+
L2CoUQaJrHz2xS3RMYcJhEZyyeffkPhPvriKAuc7PEyOW+pE0+g1M4HjPjfRSoaG
r0zEXotn2Sjs+IfTNImAiKgG9A5hjoz7l2E94747AyYZFZ7ydohhMy4ujufepHQf
ygnkQpOyvL/+nb2orQvIEkrplW95SJRtgU2w27SX+AvuoDtr6GdifaHUF/QSeI3U
pIFh/Q6j2815/ZzjO8RkKv7L4TcJ9+YrdqbSI75GhBQ8f8rlMDhonBuAxz3TbVGw
fb44vCB7eJVt916jq6GZBtxCrS5RqK9ePrWmJHb7GSPbmMbPS7Gl6Ua+ZheFW8cz
Po/H641nUui+2HgkCfWawXbAvPqaygbPgYJMevzConEvVy6S82QUjWILef3XBIjS
Va/HSjmaeLYT1n/WrgeeY0SsZwppIEe/lbD0XDMkPrmRohpOw3Rr9Ozmy+zyhKIZ
P8r3zDdAbUKNmne8Ew81IJ0UyLhBL8Sa/6NhhO0eLB/WuyorlvDRY+sMZ+0pVC5r
k6Das8lLQAlYhsx8X/9WlR7+ar7FaCl/Y4EZZ2WL8WWCVti5GYYiOkNvHay6ggdR
qNTdWSinbDkYRGhbdp5xfBIHR2k2RQNZs1l9hLgq/Gw5I3V3S6e3bzOfFlr8h1wD
WiXsE7ZmF9x3bBr9OR2hAOVzgsUoqZpTQPEx5w2T9M1LTwBl/9XdpUxMug7f1Vr5
tl4d4ll6xEKeO/ISJ+Pzos2AmyMlQdpvV/daKB9rC8y+s9qIqZgOBBZ3x3VgHWjw
0c6XWwZpRMe0PAYC3Yr/Z5QAoT5VmxS/GU2ZmvcHnXpER/REMCNp+MM+vZm+I4gA
TM86OaW5BOPpZC5c4ajFXC5yXVHSKXK1p5d51pnSGB/4bvembQ4s4fyjJks7Lyi6
CsxBgzrrwFBs4vwUKNRBhFEnyKXi5k9BBRbCQ7sbDwfAJ5rqt5AYi1iqSknYohn7
`protect END_PROTECTED
