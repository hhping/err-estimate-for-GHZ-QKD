`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuY7fw390l6Lomi4IId6PZUkJQFUxA8xm82UodRJ/I8GLuYbZHDGe4dd/sufa5vx
PaEcwQ0j9pUWd5BtBdX97c+vN+jMkYI6gIM2X1f6phMFY0HODFv3+1O0TzJokFlm
FCUrAxttdp9DkzGFS09BvZTmXxEL5TXpjvQKt2+3B6VxEaQWnou0M0/drRO5R4lw
7FP0oHfDoTz8gQItKzEkhtm8iXrcXr6iCSzQW1RHKmsIBukdywqAJB/8C4hAJHwC
wD301SvDadUebBX7w2x0chtoRlKsmw0lYAiCNnGFTC8+BknQB0i5QpuXxN78rEh+
MrcOb265VKnRjAi/QERKf63PiFKlNjm9L60FJPslMvnL0+qunBOF+d6nfzoX3gIx
L6kLhfbzzB6eYmoUYM1IxS7GZLHN8cXeb8Zbz+NOqKtpVUeyItvUv7iNKHMjT1C+
I3EO6viSM2FE+57g+TtnbS8ktpdOWa0VtJnkH5lvV/BF/jbSRShIHnU5jmto2ner
oVOEkYb0cuuq9cILSHVW3Vtjkse/pEsO10zPgd0rkaRwsf2Tapn/kZoibwYezN8r
meuSkUh6TUlFpujk/+MgWNS2Kf4OAQsTak3ACUleEgda2KUb58TsNdu8+AqMBQH/
0LDRrXt4NieTMWmEo0vkgkzXBe7eyQU8RUU23ZJu2ZHB3BSJZ+/BpgtMQWVflfMM
hHcyhxLdV9NVGJXbcehS7WVMhyz6f3nJyyh8cQfFUqXd5hlbl7jPbKPvt4e1ZadY
rEY1osgN9orSf+B8Nkfjsl5M0UWKzHjD7PplGXTJbmOSDqOYd/u3sqkQMTpTfdJ5
+OMThFFRHdnOnmZBZNG4S5exRMUE0B+t+RQW2SCYMwli1sGp/NgUiDB1TMruzZ/u
ChTUDRDjvqbF0PqEcyzK9mWv3wMcdKqJcMrHXB4yWllNdDpvjNcQG7TeuMm9VhVF
1cOnPE8YfVLF5YSZ7MzA4zQJzEpg70HMp9oAsylgesUITzJrbj9IQdYCnHTAFUNP
Wl11uaw/Fuk1wbbyxC8K52KIV7F7SV7TnfoM4rObN20IQfVkYx+Sh9tsIJlt5dHA
x3b1KNyW2sXOAn3fKno8nDAwzuHdvNXvqykopuKyGbomZJfjLBhhLqkn6m9wiIb0
Jn49Q8QyliwBw4KSyLzKXpj7b1m7ZfBxhc+fNhzZsqEZv5jcDn9PF6GDYDE5ETAh
Bs12uxpypMqyaIB6BuoJX2pTBp/Dj096eP0aUAKh0kqRBw+PCeXpb6GUG6O479vN
8/CMMq73RPB9OW7fWJgU8rRIUoZAe+GnPQVpvXY8GFvz/Y58CjL8zpA2zPjgAfpx
XuUrxbW0cW7sEW1bdVpAXg==
`protect END_PROTECTED
