`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TN9q+2BA80/bB5bMD63ILtbeB5HfmEblHwxrTc7ed5QDqa4iEtfdz+v38PjNpO1b
nky0n5/o0ZcndfCPLqZEa6LnJUQK+yt0bKZumjRm0rGGkORas6rzaB25HW0TO/WH
OmfoJdtSH98coiUW1az+sKHapgZpYVjP7IfFBHas2TGPfWKODCHF8BTDdOA3H4If
peuZuJ9cQcns+grMf+NNWsl7oMLIkP8s5wxdc30jcaRQmx11PwSKVxCVM60LGoSv
wU7zMP0UCSGauhArBAaO6vknN9SlwjxU49p7CXp8yEkJZODLPrJUY4yiKe2w/8XW
/6j8fTiQNjuG8R4UNTe6kdm8kA+OKOX2WKoiSd/SeNWy/AHRGVYgny9HNtWz5fhF
RYRvMkIW/VS3jl1QKUNKcTLcELtCSuO/cJNMDM8ohVH/Z0egjH11c9oPTzSc7Zmj
UUhzwfdfr3H0XXZTGukjsM2sYoLNtTyBjKNd8+6Dees8zkI1hOV5pnNd9iumJs7B
bwdhT1dOwQbuh4Yiu1HMU1cfcSS0BzKX8tTgFSI8vxPY+Isns2nPxt1xjM4xSgWt
PIVicGUbDCDBf2t9pkmUTJ6zQQn+zvEfsibjxR85Ow5DtkHaJHj0i3DfM6vBvUTt
R0T3vrwrzjoADE07wCij91gKlN4+auExljeq30+EBOw9GHDJEO/0DFaB0B3kFtGi
2qvK9zeqpe/xeVtYwM/gH0aowDiBMHxquyy8j174xOFdImWhh/OxI3WUPDULSjyi
kr1ViMPgykBarLEi1RJToQwDQ+0LyJbi2Nn5EVzu8EcQfbSlEdVAE6cB4EccVdcn
KSQ/qD5fvn5ztBrCww8SAjl3cXxELTDgkLoxMGkPot+uOoM21FQ/Du44x/ABpJY1
8Mt6KmVsWLEBEY0nct1AfhWq/kSbAHlnqDYAZLuB20MDQlXdbmTnBFmpsGm6lqPc
qMmefY/3LXQa7FvohsbFPdxdAdPB96JYW5mnKoWujfv4Ep3V1ClvNfCyiavOPalY
9T22MSFsCptHQsVsZJ+PKlEoAFuwjwZGVTSv8QKS0hwp90oG5nE6wF97nlPT1Hat
xYd+eRWvtJVhRv++MJuq30/ajoE6fee9WdqtgxaV2j6TL7IxunaUloeMIxT7YnZI
LGQzqh7MhltuytJXVfflzJ/xbeVpIiDJTSuducaBG9sQwe+eJ3M0k+0VoGIt8SRT
isnSEQHBOjIkwvtfkJQOoKrp1LIrMpGcmFlyiwGcbxgBQx92oR2pKSFoxTLE/Z6z
7t0S7ncIkr/xfw6NrUMnypPG7se7hW3cRhpmvvSzwxrYdH6DKeNU4FG3m5fgpCo/
+8buo4qUheLOQoTk3c0PM5qfw3Vbp/cf88Q4snxhIKkLLCCf/f5H7LNJawsTjul7
da7kEUi7T+MCxDACHaulH8/a8hbaDOT3Qx9PdBdLqXdlCMyykggcR3RkOR6jJK9j
UZ7M6ieCqyMz5I8sir2tTd5bBxhrsHZGAIxZhVxp4B+lOyEXXHb7lDCvXTjs0BNH
MBjssD4qGWBPaqcRJCVAkur/NfrhQV5KKcglqe3hlmDdjDguEjv4NjRaiCbIZ2AS
8/J3ovtKGny7x1F9vTdrJU+ftjIrPwX2dmmC3J5DE49U2c3nVevYrpcoEMiGx7AF
rcidFNlUXR3HxzSOBMXLkE9TlzLkNyVxahKilun3daGOG0WdcRC1LJHrr/lusktK
NA/MByWvOEhyti4fYZnIzzX7GR3XuhaXSt503NloMrXR9Xt7ndM4YP2a0GdxcRVK
L5u0T7/Xj3FJEgHOkbpWcyJwM/QL1w2LM3rV+ZdsPAfPmN2Pzid9pEelTATkfAxW
MwuBZ0tzuH33DhjXFcjYMsVndunlTtTEfeRT7idg9Tb3zeGlWpxhUZDIEY77Bz23
hIG90eS4BwONPI6lDmqb8M1my7iKpCiDckC0hLiEdmK07O3bFQLPP1sWu6szoW+m
X+Qd7mvIYl0OICfGvvp0QSJvuy2d7yYJaUiDWwPuHw2hP0Rqw7MVhU/Fv87WTrPG
b4kAEFWZ6aluADJIZZEdN87lUWc5CgYYk6aX0z5IYT8SVk6qk53ENZDizDSVSPaD
/nE8sOePn5d3jI6ucd9Pzu3etNihYqXjPhlMYlZUn2lLYTuio6cSKD7lzJrX7pwb
SJHd4yPAdFaNbFt6uOaWrEY3Xyi6G9SOMhD6MCuasmmm01arP0I7VG+vosfdckVd
/VonKBHZDLSSUDg9yuf3IlP2YCAuCAsqK0H0Ol/a8maU88boz/Hs/JrwcQYi9iVb
ix1/pc/ZZZP0MT66RFDJi91MMhe5ZO/0mZ0GzXyZJw70TkJ9R8jLZWgkT4gKfxmV
YTY8pQMysVNt59IA/oudnZbx7uhdCvpu3GVV55Zk67z0EmYDyhhduZ5cdu5VRV4e
hMcc0MgdmLDMHLB+zeCg7Pua80Zwc3VvQWG2+iSZRJg01rMezGGcAc9Wrdt1AaoV
O/6epSq7PkrlQafsD+mYmyxa3+8c1C5l6PUUy2lQw7V+tF5FI6EfSwMI/Uos//ej
zGrectK/GOmuLBTfK9nZk8lgAbuMz59XcbulmNyVu5gY+Bo2Gp76Ryg2hb0H3D3Z
s83U0Gt6HCJ/y17EYPru1WaKgpVVqPtEbBg+LMkNNsQi9D1hrDxV4Kxa+mwLEKbS
+ZzxO+F+KkzctUGJb0sBoaOkF/9hHmPv7FDWYuYQ48Fh8WOLX4wdqai5VCivszKK
yhuDeafw7gftc+bSrbTgv+hzea/YmTRJtFNWbIOTn5jVJ6GYArs7Shv+4bRAycB4
f+hLxV0RYyYU8lB7LVwTevRbdi/rowI8pP+slwWPLwFupDMJdQAVcoHNcAddJ3qy
E5DVMl1Dck5aKlFw/3/17zWpCgfo8hI0kYHvSVgF/wlRDsYd97nkD2VQVngpz42e
UX9gw9VHSj0wVIMszU02DPvQBvpRxgDiD5JgFHEjDiH3WEXAC5fjsJmm5yHr94Er
`protect END_PROTECTED
