`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sax0shd5iYMt5J9aow9VzC+drAhARX9Rg71ohbNtcAv66BuXLlpDVspPDMTEci/B
xqYhjYWqsfmZWsUDFm2SL4fDVnt23mqTlqpinkOgPDzqd9EKGH3zDhcI2XJEArOa
3v+aykqsQ+Dx+oS9iXgzG/DJv5iDKI58Sc2fItmEOnE+Gh38dqJJrcuhsdDPZ1Zn
jORtsEtyV+v7s3TxuX+JR8L6SjeGWEjuJPJz0Sk5WwXZEIbL8VR3dm/AqHv1EUt0
6md2rfzLIpQ3MGPStAcUIk7MbPnkEV14cPSWfZ2lpmJtvq13sVgsaseiKeOETlPK
o91/2oeU328+9NXD9IBeEFXCcV8Bf0Yzg9Xta57J0BnvaxxzsMrZWwb+mGBQWzup
3viHBlwMI0RnLxXQsChhX/XK50JvLJsLYAnblvtRD/ODIXyvdISGephyn85mCEKB
Z0vSVc3MLHxDCHhaNHPU2O7qseA3ehmTlO+LhFKJeyKyDj6SpuvNS/+Tckb93Cdr
wca3APBI/VBf60JarAN5isgo6rtKCfB6yYEaSFGZDBtCa1KYWxijoxUiuYAxzPgz
zrh5vxksJfmSoKwZGmNg3dsDnf+daMc5VthQXFbvfY7bSVUNVPXyVlpRk34QsrZO
kdKLMG8ovZEetlPFij+zekuuOohTgH1nrssL3vg3qNkSbN3zozk2BwMQygq7yfWn
ol7e5lCG4NO2wt911RBs5nHAmu8asMVwbQJ8KG1GSQgqke4OS5sPXPBFP6tByH1/
uu5z/yCkxaTi/nQw7XgmVUPJxKxKjSg+60gP6HT6d5sUZK0EPSr8MYizaNQ/Ecsx
9ztQP5fhMzitOU46rHiPdPzyOV9yKamMzJ5uf3uFnjCpU7u+PnA73IsRgtXgi5sD
AE5/KUrXMLWV1YPVVH58ffml4I1zLApsb9Ik0ErJdWFfHPt5erj1t3fqL23SzFR7
Hf8eCnHWBIYlCGslYj6qWOOCmYn6KVgeuyoSD0s4YUlXSKU+y8qTpP2AFOGX8kYy
RkVtB3vICRYrSa5CmMdLt5WGk3G9mD0ac964HF2GbN9BY8fFYKeAfPMJHuUB19FR
YYpj0pLgqyDnwh2gD6zUofnpvuzyIg2HQPs43R45iJ5OmDICr+RtPsLQMo/8Kl6r
UnDnsjPautAf/El+Ufilisp2V51g6SJ92utV6eyJHkMaeHRdaWIc18SXrvz8GS0J
rET5vPOpOtNi3f4ci7wajkTKdd2UH7vK5AH72e38dUjj0HmkncQS7iDPK1hQmEiT
tRIlUO62lVJRE3q5TgTkcr4we02gl52mhWv+Vg6OwDy8Ugysh5WMzOoie5EhKYL8
8vZrcrLwJIgH8tGsTyo4U8dgtUJ2ATWre+ovPpEjkR+kEFZSaqNgq0J8hqhKROqt
Dbnz7a7xJGFzpsc7NbPBXeyITr3B/a02+QmHyH9NMKsDK94Tw7su3OyWYVo9X3DG
7kX+4zjou+/4JUAzKFbFDHBDW9Q7+W6ezCPwPoQ3dkDVdVys+7FUUmIqkL64+OK1
Xb5wckDajwCLikOL1mcR96+bLfnu5fl0KXwTZnBUYds9E7DIz0pJ0HWzStU5aHRl
/4U8PJ8HXjZV0d6Ci8ehZ6VInN4V2p/rTGcJYlQBWhdTd6iIL7aJuLIBhRKiCMA1
dY4XBCb5ZPbfo48VmZoyWbWGSiCW2Vufet44SloEkfMPpWVjNNISPMWdU2decG4S
uqvLJH0D5dP0zizbXOKhnXTj5Qedg32QcMb7+TP5CKSadasQxKnlwyXjyKM7/J5Y
yXUpydiKOTzwNAdWp9NtTvrfnnxOZ6fvHPqcUOovjDqcH0VxKHcjnSvxZ2j9CkWd
bpyByyI0rCX25Pvd+V56F4YaeGRYXEeN49ifaXFZDkpbgWV6nRh+BCoiZeK8woKF
d83ab0u8rCiJ1V3IFd2cbpBtThPFpFBUTiHQy50G5y6eGls0kR1h76V+KEOxJRU9
eJs2o2a6WsyrR1xLDBlnguWEjPTtTNRXTmyMmBavYoER/qHYDPOffSJzBWIC/XUr
Zhph/4f5Czq/jkTb2dmt4Vt+r1fT1gjJBChVN2b0uIQf5A/sf1BYd1eq3iaXtlY6
z4UckEQFt3V6/wC6XrzUfS9B011NLmsEEuw/ZfmfTPz2UcOvwU1FBsS0A7nT/xIA
lRUmR0K7ExFkfGglreFvDiTm5Z5dxKoGakv3iVywl88WWIh/+76CTOstl12mjbF4
UOTN057omWZO07MWHit0vjjjYt87tA+gH/wuVKuQDh2HJuftPx+3eFMFgma+LH7O
ZpswrgoETUxNyMKb0+U9MhuCVvfmE6t7mYFwiz4UL8xyaDVVnW2OXijz/UbBPW4I
M/zcM59S420iM1E/WnrdBt5h3fbMFvaygfNMbo9KhQNjDSSXZxE3iuGUSrwLHHen
zoiSGKuCX8jhleOPivOepTjZaKoVhSVrR5v1UX3hcnkDlJVs6cmfXhNUCmKfSL7p
MEhiAPdxU2660SOl8nVgzLwmc5ElpfEswodr3Bl25aRDZA6gc8TPXcfol/qP+dqm
HXGJMKD+LOfUJNiY5+Afz/N2KpKaIpxTPDwV4LdHCfdXp2ywV94+12c50kp59Ere
x3d/LBEphrngoE0yN4uddetqEeihEIq21y0GSN/jJINlyxNz3kTuNJDGQ0JVtH6K
ipqEn2aYN2cUshJlQ2XNNrFsE54VRy0w8aL6CEyJ6Cl/RZm3kliZuWdRaFRqWUgb
UXAAvLKHhj2OJsKrDZd2J2osRighB7+BO/oPUU/Nu2dzsUuj0skY7I3u9GYaAhCy
E0y6c+VxNrOTPSOF9zgtnsLb7l6dzGN7sKCOrHhAiB0xhWL2kJFVpi183QTtSOhI
NatorGdLhvm7EM8ouqBwDYFULxQx6HKZxVXL5evf1SmZ0XhNpivyFGLMU/QfcVfr
K4mcRRTyGAXGxllDgxdVdyxS2QOI9RbiAoevEf/2qt0lCli+LJEI1ENSjz9hQeMo
JY4z1u5o0v7G0z3nfhpn/c/i0lEM2FYeNIL/JqtSl08uCL+vpOV/2inthkzVubIt
Qr8rIYt+qZhM1V6hnwNvt0ioYb9IaQQoBbClsp+Ci4AONnaK5jM0SODjrpgfFqj1
EtvQzjMwwDn7q/I+2kk7WvUkiBqdqSyjYbu7o+TY2+v1tgq6VjO+uCBRnBGH5O/y
E1tKTmTPfG8GlsFTth2LiiPy8jD/wrqUTVYcRvtwljAxc+nFGCtc3MLyG4r0ERSG
8m9WDZIhdeW8bxKEYpZZxhB2VAwH/XrTmBGnRA1qBFlBo2OmLPfWJUooE7flg9Wd
H/lZ0xM4fAQtxtbL8GnYDthbw9K5pIwX+7/iqmBnXrTTkEHLTeqncSoW+pY9dA5r
yUVXMTclv/8StNFDwWaY5SzRC0os/R/AY4fXORyPToUwyOvLi87zgHgyPW1yHZ0j
+gq/KICoVBh4Z0/k7yvabkPZOKpFxaJ78n9QURETrb60FjROzZmHohuaHtDT0nmP
BLQO/EFjyNR+sjBQIMah/OvDZpZpmCbm4OzIJdG606rfO12Oi9QdOwcgE8GrWAoe
YdJRXutlmokY513hAxQu6xMPdxPath8H440cvt5N79JjbpZ1wnWfylkNCGccdFlG
q/rkmuXoS9+39qMfpxgv44soXhtetk1eE/2ascnB40yCmvgndJwK2Hyu1saltkxK
xOZdc8qit5fjva/ebCFR1/X+IyJjKAWKT+z+wWMh9+kIysmoGhaI71vg6c3tnWbf
3js3ll3Nk8HhRyMB1sI4Z4G50dOljEXqDhTDgs+YTUX1Do6m7hWroCxw6/PfTCLk
Y8QdsRUM3X9WS4wLya7JcIlq9DA9LLKVxgbhKe1oh08mbqwg3vWKOf7KhEVSST0J
4cx3J4ZhDsRynIgXhKXZOMmcZpLZ3FnGImaCrAf1WchqTjvGh4+5S8dnhnJW4AyL
PLvtCcK+HJxnC+RTJiUHgAg0psHBBLY9P8EEufFgY/F0IpSTJex8wk4rxpIbhGMs
0T0lmAsNtvOJU58HH4+Vzt/YYZzn8yTvNNjNStMUvqh+WwUXaOIOtz4bSSDG/enA
2N1Z0JXUMgocv7uEvLGyU3YNFsp2KQXS3ur/6Gx3PBYpe6TMwMjYdFal85nNbhj1
R2NLRPJcRf3oOIFB2I4fWdv2kfDjuZSxpPpeH3Cdje15n8E/kU1yZ31Kz6jGqCA2
nGwKxiq2X3CwkqO9S25TKAOnW0lXF+zogr/0rscuSJXlfjqL7EfeEsIT07c0wHVC
dIHKwwXfy8daz0FLfsGzlehfidhWLnkbwGJKYw1Bgf7DaLspGYpnur7ISqeGn65r
axvuIzJRlyee6XjBK+y2hwOD76aABPFMWWIyRnWuEQ2FHAztUMgByScrqzEVcw+Q
PThP586exLK9HKF2vZxQPGsYqd3lD8XWiCo3dBZRI/9B9NZZwv/qgA7hvipm+xWe
JrFZWbiIaVeeydkY2bpnUHKFdF+tAEMeUYMIWjJKBWIpGpncFTqv6fk74VJZvtf6
5WJO4SvsjEFs+ExO3DhEZKywUQAcuCgZQ4N3AEIPpwdUeWxUOrl3myMiaE/SRSBN
r0PbDHlziH4cDqw6+lK5sfncvGn+spaQl5a58XWEFu36t3oxiv4fQJt++AKQyb29
h7intAfP6UuE3V7zgSTCeEg+VixyGCHLbx7CSJMdAD9iHNQ6knjMsRmYojoKVvbv
UYTV1uLONSHEFzrxMucdS3XuxNjgr+fHH+FYjp1UnfV9EJwBLR8pvumhvVH5HVAQ
3e7MJYtsem4SKhNRjDRnUf8EfeN19YOmrHgTWR7RbxNNs9i8qcwoQsZDG+sjADXD
62OYbv10JM971cNUAPvJuOYhoTMWEZ5idGlR8PT4QsMMR+20+FTDsAtkc1wAK05B
2bscFLvMnZsAxBAXciRKH/ykefj8Fg7siZ9p69AIJgaRa6tkRuB/PxFLKU81FxEx
ZLqF0ng/whMxl6396aXsXXTTJf4Y8pGKSq/nhII3chnCL/XEgzRNN73m3KhunP8G
FzlJmoJ0WxhUYLkMeD9fxfUmXOgz4L5FwtcgE4OQZLuBukAiMjpVOZmyfIO64hl/
HIvG8A2LuDICI3oHfvM89hoSBask8l95bcnGnoeLs1ujK7p53v2MySJRaKUyaInK
F93zgoPYngi2dUjL12jQu1JT4D5D00BAyeVEXSsR13s5dbsJ4JQBTtx+tYX4Gq/D
mjhxjwZ6uBIOrggGsNUg9tg4tHh4mMhIHatHUrXx9fe321vPvibd+DPpqSJlmEoK
Yf8ZvJYO8szhjgSTezdTWO2auYK+M6JVMWUAkDCxxARdoT+NQa1vgfI+lpqvujGa
s9ewuavzlm9ztHLspr1DUumsCviHEEFKP/Zcg+ORTqOlJtb6Ksudq4YjRx9wwgPi
3/HCUedsJaxwu0wZa+yuyT/ARVL73d+elx5Z7wP5JGmG08wEnTf/F6qD5mBbVuZb
/tbpmT0dI/0lOGbYT1qP+2ov6eUV0I8jgQwukJeW3r6G/m+nAlroB5euhSyb8IHt
es3H9hApo+tqE71UN9vDvbwn27M5JDWCd9ujTi5ZA8YYcrBpfBUsnj242rUOor8K
mNZ0Bthi7t1s6DgnsIHavEG8sFZsg8Y9vQaLYGJS6dFUvqODVLxlFD9QsMJnZX1H
QCoQVCaGn/FNICy2svF3A3qf2xPdeRYhBYlJlNIdU68PsJce6+2asQipthXejDTc
ZFD/cH01LnR/1nwtohVFAr+0zGCLEmbCGHS8nmoGeQ30jaTVY9ryP6F/HWIuEr8u
L485wUyY4N/MMn7yHgPlssJ5EIexxZRg31lE+X7S0FsXSoKkBNrbEfxG/D4xjMVy
rLyvorfsn+M+f65Zh+v0sH3oFCn+2/LIEjaUoWEbFuk=
`protect END_PROTECTED
