`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqg9vVQDulUKkbJmxqT7RKYi7puEk67TRlrr0CFYRUEpLha4TAiYXEk8kVI5GKEU
iW+URgnj9QESOZq/1TN9zBoMCBiZNiWbHcXzssYgG5XDC3UUjiiQITUzzbdcPhfL
KFjT2LYEyVv4gvadBQsJ2FPgx56Do+gGfCeoaOTiIq+4JYr9Sqaf4RiDe80UZ0yG
IQenaEXLkjqNSAolDXvaJwqC3yUb0yLF8/cL8vXsKtXHQXsRh6e8lhZwW2ivlKtd
dC6WFPkz2j/tOkONiiIKOBDVhT6p2FYa+/cjXsVYK3hbXr/M+EvZsk00jKoLj6pt
XLRs/Rai4V7hKsiTGX0iSQH1wsyY5bZh7uKTwhh/8lHH4Y6KVvAjVJjnGtulG/zS
bFYRCJpCGT8k00F2MHlvveaC9fzOQp2PhLQNAAaazltHhVF/tKDhOUA6Echl6qDO
/wOu1CrzdWh3RGPqgOTMJyrI1Bj10v9CqN1IMbxMkw+oAASZ4jqfmnzlFH1lVm8Q
gNFZ/VYe9ozJ6kpPie8scC6PdV6a7Dv4cRsaaenTj4hha+AosbN58Lkk0aYHYCou
CLHKRoR1rOha5TpbPKt8kLyt8nTdFDAG/m/zGdZ6Qgcu+J3yu1t8cS61aGbRziqO
XZ+JoJU8M4Q18sZm7/btbBlBTwjaCAz7pR8eE+pg3CUZM0ZzTt3UMvkboGeKR8dN
l6wbds4iXsu60mXp3dx0g+DCTLSvh9oU4B/sT/6QZrZA5HAS1BOhoWKUe8+kytha
s/ck04b/frIsF5eVNLbuR2HclYwvBMuPyIeore4AK5itawleIC3qcAxsbdDO474r
xR8gM2Ajbsp9vT1Isbi88iz3IcxgS1JjR7dhfRnCxCx8eC2BrbUMIRF4bgXva25U
sptPUTIw97Iql7rETajZuKwHSSPTNvj8L3/PvxMsna/sMyexmc1q3v43vvCqxO3C
BQUt9oPZasknsL0Hdi9Si807qJUkljLejk5bRUn7FziJoivifeLn5Ri9pRoYjOoj
dpsK3xiKyVWjgC8/me6DPnizyur55f45UbgZGY2PERgOeowvl4pgwlRqa+FurWiU
ffsMirRL/DHfa49vpboElIC7BGGyxyZyMQU8aiA79/axaSTjCZ6Q88hEq74XGSnq
Xin/WGvePlzup0jmh+lOThh0j+iEPbhVsIv/VKzjF0opeUS+4Tp0Hoa+COnjqpq8
8O1He7T3uyNy0rql2aOi0f1b9GQNugwCHoISLV3Adq+E/We/tYSWISsDkculwNjH
ZG7lF+UWusbCwrcw4T0NfUbBjeCUL7I6G7rSXmpXwLrMdro2EogO/pxrDG+Sm0PL
rkDqzmLxowXvVzEuDOAT+QLTXahMP30/HMJLFBKKKMrViQM8IZiOwSYlnv3vywOK
8Op7wM8MfoOGB2K/5KH3Vru92OM19yxA0zluE5ebce2Kn5j1BKdxUc/h56/qNFZg
wWHbSegrHXxvXoFkiCdXYIMzSnEuACu+QZLdSs79ZIua5UwXb7jVvvU+nXmc8Atd
v8zO8E0hW1LgR4j31LbrTrJpYdSvQAMYdgoIdjz5YsqkHVrOliiuHn5YyGxjWn/m
euNurOCGvBBYrkPT1mhPdFBD/W5YCZ5BpuBREqsJLUHV4chf54FO0JovhyZLNzEy
tS7pQSxNJkq5he2SwZUdwk2QL77kr0/3eE4vsO4hdHj79Y7fChEzpWEAQcRFb+h0
31Oz/7ZcATGHzUszZ7unQBwbq6lzJGeDpNoKNUkEo854ZaSe4QQrnyw0I4AeNLpD
7tFUxgJpWVnO+fwmQ770J2FAUrOFB4+uw60WS+C8wRm1f6MRY7s0hYu1JbyIR9Nj
tIwM4ceXfNWzhnsusy5DoQfLNr9+FvW7zQbagV0PumWy/TBLLUV2nySUwOavHGjF
k7IOnmBJ6fpc38QO9hB+VIYItTV9yuxdkfxPxKrclIoR5P4l+feYKaIfgqL6w4l8
/4jMWFpgZ1EeUCtBuuoyQCGVpZYsVmniA+zTOaLFTd2LnbUD2x8rLKFFyv3svck7
bUW68JXXqwNVxQ3vdQPlwj4Uok5NsBEkZU6ynqGydTIzDGpdjp3vf63PmXJrKE2b
HIXk2Crw6y9vzBCrI8BhtvdWrxMMwKnY9Tjj9ZzHbfJLHPAi3cX7yOZ23Jbuxi6m
Jxs5gOPf4r/r56ukcNCUvrNOyR7VJUd472FcqUdIeTY3CqIHtNudR62o+G6HoI/w
BNvt1p88Aa/fCD9LYz0aRaDK2GQ/h5j9TMV23tU+6aw37GOUfTArG2z6pfpUXakD
H/6RFKYfTJ8tQ5vgixHXZR7IdfSeTFgNcUSNMT462W1vWq7QLoWA9OJpTuiUrFyf
YKvt3B4ugCY25HqQD5aWHIxDnrdhk2x/plJ08QZ99wtGvG5HTHHY2bnYbaKp+VNp
MXN5ZtcOJXF5Tgs43XPMFVc3/S1YqiDC7BKf/sIt95Tnu1u3pdjuj3RmSpCYfv7H
l+TPzKtg8Kh3islRSJ0zYbPnFB2E2I+iKWzzIwU785Fkz05IqqsRfnEk4B9lAve8
c/mdKtb3XYFBfKeEzyE/GvdFi8GLCgk+6zKgzimqbAikvneN6ByJVY2Tq7HbwjKz
NzJb4KvQWBc2Ocv8l+4Osg==
`protect END_PROTECTED
