`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCSqTqRynsfnVoScsLffak3tw1zxjnqNN71tf7Y/lnDsq+FAxVTXrzmKHuYx1F1B
wGIU6WD7K9a+po+O6y9kC7KtgKqCpBMmtdMZuids0vFAW0XHLmBaMKcEfpYoeJgt
gItOZNMUNU4bY1fxOYrftU5ogs+cFF7NaFSXKVIcAUqFb735VaFNAZniCymM9sVb
uggPnbzU8YlSTqYwvDuOKRsdD6rCmAywAma7+Cot072A4qOJVUtvwFeIpDLGUYYH
ks76E8JGi5lfRswjuSceu+z30KuzZGrGobp/4cUaXEmJEuV0K6cpAFYZATDstOv7
iI8HzygI2Y6C7tAHC8/ySPej6au6CEUgDHLTUTRH0ZCkAIz2wcZvqGFMr0GZkd2m
jc0PyAYzSgKO9lq+2dCbChzFY+zrlfVC8e7CVNQOI3dMXQGE2IG4/B99PTYyTODr
5kzW3wxsoEjrqgRlr+pJdUEKZOUO25RrwZR8RR5DcrA=
`protect END_PROTECTED
