`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogB5o8x2v6DyM9aA+bR5mwxPC1VvxKMqiIGX3vT6mLO8r6HfmKB4meAYz+xCkf01
2u847DP7QNVkop/6bi98wEfkdEV9Z9aGARShBePRi0hVSvqplQJQ7HHklSPnp0kj
xRKe1tGORrv39sE8cMBXvjOIe4+As1kXG5JMsm61AvrN/BTb2SfRklxIGMvnUksS
fXlg39hkTAewwlDckiVbrSl0PZjuQnCQc5AM/Un/Ype2SFQtdebvR77gwqYt4t9b
dK/9f8rSbPDRmL2MYi2lclnbaHhndi52aEBnDRxT35EpYviWhobNc4Vg+JCtHKF1
P0q6uluPY4RCnslWo2FmAR3Pxr2dfXn19TF1++YyXZ2By3AkzO1RUCNbvnTtDQyI
oY0pLEwnLrIi+fdEKy//dclusSzk8Gb5hRgfVtpkQbJIw0Yx6G0ozO6HuxOhA6MJ
lq47FTyHNvZymwkvrPjGj2FFpI58wG5rj99ZDTFUbrIJac/RPthP11UBuGIBpqD3
hB2h7Ho3x1X5NB1D1uUPQg53ItStR9uD2uboi/6KCcMd3qE0YGDIWf25L4qpydlA
bm74b1xJJSyZcwyT/1ziH59ennhB/V3npdi5mLjx01usn3lJMOIGE4zOXehTcpBA
hd5ryEzHX5R1CuCDRZ/QnFVQhhEJFFDydrOGUxcDOT5RHzMdjMEHBFf4tAvVIq4a
0QRFKJlH6bjdblBpRWivomnerF3+m05RPd6D8ExpqzJYeKEakjTye9q33SXgWzHF
BnfqMIF9gvJHhUS8MRarPwnqSIH+h4J57HjNd0S0l+EkSX66Wcf8x/a6AAzbe8B4
rP5mzkkiprm1eGENMrKKK1jVCHtSpOsEtjVM4QJZEilAr1hZY/MzsbAa/U8tatYi
ii5HMNlgoFiTwfRshSDcPK3SY0hWxXZ526PeE3WFYMZ/KSEsjNurBv9Twf3XdfgX
D2z/Lz/JlIP0XIiTmREtws9v1M/hjlheWBW4yyOxzXDqpbNU6NDwbKg3lcLYDuGR
1qWdZqaeAOfjWA6vAMIOvTaz/XU873rAzImafhfk7qOYFEnyHpYS3xJgQwFrpwz8
ZauETuXkICJhdES9G2CnzK4lEzrPtsuUMqt86SqVdamlXFVle1TNFbWTE5jLNEKz
37t0tcPR+6F0Gf8H2DhRofjUEUJU3tBGmF59PYNiz57vRvhsVdFyimD0ginhu2Ob
9h5iVuzXe8AXeUE/DGo3RZwyyTE6k7j9ob+5TzJhHtzyBcmDKylLraEV4FZv7gCY
HV4/15NnRUA46mrQ8nnmLBEFqy6cvLvceTPFePS6TlAU20b2ydsXkti5DpH9DFZq
v8Woj9Gm71B5c2hMRFFSdgeVj7MKNheMH+OJUQR5sq7xf/kKtHsitXFakyrftqP7
rj+vp1G46BwY5z/Vhj6iBZyexT9gw3UHhIKAe7rRjp4KCGZ0+Y8TZL9PbohlBkLR
l32BdGYAsudlr2pTyeTe/GGIQerV6Mfn1h6krAxP5AIk0jDhJ4ss1rd/4TAtP+YI
9qjCanaL68fB/6Jp1nQNDqiuKyHnoXfI8hfudgE9IrhhnJqyLSglfbGpjxaGIrJC
dUMITY/a+q0lv1jYaKlYBbrRwV3waug1QmtVq1RlOy7UacbrvdqLamsROBYfJZ4K
ddvPqusC33GHQ6v4+6lUBPkrjGTuyGfN+ynKuFfk6AdTAZ2zyxJ9JJw6OLNDa6c9
sEGMgZ5XXI9dG8VRzOGDLVcSts8eV3Q59RfINl7lQ54CIVXO5gYUx0Xa64+huYU6
E/h6uSn3FFAGchsA0nqyFof0XvfMTbwUG8ePfabkr2x85mk6DySkfmTN6Tmgor3z
OXBtuu2g9RZY+mPZVAM1g4otPyZBuVf2+L7JLc0rbj9GBngEHGgcDTQhGwFqhvUY
`protect END_PROTECTED
