`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Piz3eM1PGq1XZ/DL7AL399uHq9YYjJyPVPEaJ1MqqiaxqvLEAYfeuamBQKHqmUz0
CX60a2TWypymLCxw+Q97SlpY8rpHyU8lT25wPZw0ClEdq8JeSZYcKSRhduPSO5VF
OHgrNtM51TzcrBTmY5tXVDD3ebmp2LOq+Bcm5hAeWI4mNpZz0mLjcFNXFZuLOBEw
x24ACzXLZqtt0BoPAPh8uVochP4X15RHEnsSZ3+3dOhklx7cJ24lTMnCVMH0m3tC
qQ3Fdu1RgWP1KXsluuGbt528R+1XxPcb4y1TZEpVjQFStPtMG9YKb+J10A8WM5+K
jFoKOhBA8XVz1pD0n1fBuSGwE4WjVdMFdCgc+liJ0C6ubK/st092C4v7bt/d4e4Q
z471gqw0fBn3s7X+vgbzN1nIhFV91DEATEMK+z3R47SeQUvNfRVqLHaI7ZSjjy1U
BwLp7MVd65MKq+1HLGKs4K1wuzvYAA/sHbvFd3kTUUq4o8BqDDVCg/dFgCEeJBIb
SnPwA1aaaeXnLuylPIkoCAW81HlP/4HAWt4lydUzQ+Z13wg/CX4z7tz9EoRJpdwK
e5/vtIBvLA1ljOE+YvOIfqKeS2+Vm6F8LsXidjugbZ+gCVPwJC7nloqQqgBJG7q2
XsDNEyK1FS1r31kjbMdFhcElu+iXYPXI5pmvm68wy4GdB3j/CXiZhZA1nBavKzZe
/a2+/1jAJiL7Dn0OYBPCFE9DanP+aQhi6rr1Rrlth+xdER0ql6pnsv4Z9Bt1xm39
c0LG6Sk5XAB2rnHKbbctMxvGUW/FGwKAIj2o337T0mTWyGu349S+MDrtmmfXpnNF
ntrsn8o5W4jMuE8EFaiGeLJ+BTT3a4+J9OAXWN6it1h1NA3zphzYLWj5hbqczUfB
co/y3woHwMWySoRJSx4IDrBybKVS5J9G+rkp/bTwTnPTGAfuw675erDpiP5FPtgt
JS8Wlk2N8ztWlcQhM9BerRh73kmtDRVTig0pDDcA5LxtPlXR3UgKZhT1v7pYYUNN
iEhUr5KfYGXfykfRS6ZRrAnsHnBHsrxHPcuepmNHYLYZANDRa0fhXWBoDbX67jlz
/R7LUiHhyMhOPIVQknNdr5ofHAHSScCkx2G5EXQYKSvCncwhVRUC2BNKYmvv9Td8
0/aURZoCiEEf4i95pwD+lt7FGi/x9mmvo9PmrvfCVOEIGDWpHwUUlZK2ifwbesJc
MuxjotxJjlQArKjqv7eId19X4Tq8QthAoz1HQt38UP86HyLdvkLSaR2klrbKq9wr
xY7R/M1mLgM9Z1KsNgh0DdoywQgd7Y+dIMNZw7epkBzQnY23sgHbT0ZK3ywc+8Fp
DHgFcPFhtAsuf1amZd467xv+RrXxReyTEBGSWWcO0jpRVT01AaO4dkl+hWqDkftG
XRDZY0WboDN3W5jmf2zWui4n8RnYDO4uViA4qm/rz1krRthECwswWwPKkCV1PpxM
E46Qh0dY3wZXiTnoVsQ9fTndNKakW0lneZ0rPnV+czw1EMh/gHb03OrKNvGhKrOy
w3qk33Qfa2iuA5Ha9cm3BQirNlYcvsdF/OaYfRaytBe42cx5vi6Vg0eunCXYdMvB
epJuw0lGIgqT6Wq0NaNnJVqkgJIt5bpexEgeI9+ZHh9GeW0Sd0qa+oMbMujILzi/
orM6kPtkKNt8pTvVewYhtNHK+1S16/reSJLmNjgx0IKC67ndhYAP1RGUiJHslq6U
AnBhFNt6S0112BXk+TJ+WemjbLqQ4vABCaYQckMt+RjhHe1dXFSbr/plk6Yxi/zr
erfryXhIHy9z88rEfZrTNkuUiL4b+3UM0zPbe1mcUQAt2xddCFfM2Thamy9yo0IY
GH5K1HjN1UOJ7+Aogy/6OuRA+aYTajA69q5pB8VAmvxhkAPAzYP3fyNwqCQmEnK3
qpXS/PD2NGy28Ac+CjXOabb5ryk13xjnteNSOExRXKUue+WQy/elGIp4Oli4O64y
kU4qFRhHQRYLKrKTiXezy7DL0edeDZzSnqCVeCcoMQA2g2y/ok8RVepDZoMPDomN
qcnocpLdcDZxD8SAhn1FJVD+SMDDqO7dSLODETQYO2XxgPefTa4gljo/9sn8Orb7
PBT/K9XW4a5rLq45OWP84spItcmxf4aJ9zi9j90XhDxJiiIv6A1VDa7xvOYh3FkX
F59IJl+n4aNZ7QgwNt8NfEvWsfOZMKyT9IcD0zM/NCj9R0cIORMk+eydZBSc75TN
YcUt5+v5E8dkweTzf6rnu/+et5c6rhgrFy1SdD6f25iRS8T6i71zat8spAk1S6+D
VLlG6/FjYNFz/cf92LX2nn9eqmPFTPQJ20RRUrWsniKGukgO2j6+R0Z/ThbJ/w4W
zyd/CSzvKUG4GETwUEPXClaKRyhvd9pbIAtHZj/33DaoGZPOYBu1Kq0Rf/KPrqvV
lMH6hvS0K9ROnETgiyySOuuPax+hSg2DXZ1QaHoIjYkwjdlt40vKNkIw2cz8EUxq
Sh8mVS2tdwZ+YsfqInSf+Pdhy7Jx6UG0qkviwNkoJQwFRem+T9u1IGoVNWtdKeDM
WJ2al5Dnqi6z51jFVea1sJZjPqrmWcaFUUXr++69lJNw9AGcoSi7IkifZQEz5YMh
PNqt8PSs6Xt5JIeJKEwLxQPGbtGE95ISvajsDl7XdyFf2kdd+s0nTjzgctJj+L1/
KvwWnOFt8nz3tZOPazeyWfOIdxX17t9Oyk01FlkYS0qQNNpeb8J5afs88C0GdZxM
wYZWQJB+LXL+fUo0BicuoTbOw37VSp9qtHVL6+HmCFynJi5TFniRoBvsehBoWD70
X/1/30yz38t+t3Tl63XW/kDYaGdER8NziAQZKflDoiIBwPrAk5IqJpPFMyLpMDEY
1L3vpVRKLyfgDJGCWOhSaW+Vgx3U629klV/JoDTsxdYLNxMNqsu8XMLeDXhmAbeb
PqcwcyLHtlqthCV3NaeAnoWrDB4U33U+/CaXCcRpfQ9+dgLTRUOrEROgvyxkyCfo
PYL1JbD3ji8Nlyq7OM7tuxhQ95I+qd19jVn5BO+HZrhhUR7au7YIOLAJDmydNfUr
Tf4Pxw/V+Yaj5j85USsAgaoV47X3/TpCKTzc99uJZHaEbJR9HR85Uym+kFxNXjwx
SjAWGzIEDkHjABja5xfqk4D50dQDggJzJ4GtbPlkITTJd9hfDHR+uvLNXYaf/Mbd
aCN5GzWsTJgBT20YLmbv95ww5vk8LZsrG9VMUCyBVNm1w9N64f8kYdWBi5zqA7ob
eHhSkqGsGQBq9fs7Asupvx14m09SghVtaEdbN+M3Ol1buU3ROumwO5UCw6FHkO0B
Ulk4aZyJWZjHmoqWpf5hJ+Z6tBa2+9dmjmi57H/cwYTfNSLIQR+pRPe/OUEHQM6W
jw7xKBN22ehbWMlIKQGenlATrklX892yPeAEBsaLUkYyGtGYIQL7HD0bTRKV+JAn
E+G6F7eYpgmeGSPXnyPYcBUmBhXXhtxIhPzRJIsdiKqVwUKowJNlqJ9dZzt22jmr
APWoZpKXM9UotNsIGKTm2IWeVv7E8tTOjvUCK4OdBzOfNdx8OEn4rcIItEm+GyVj
19W+v9hZKtecVQsIVUCJYQ==
`protect END_PROTECTED
