`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewMlQpDVXl2bmnJqdREOskcnrYhKXeIEjr04W3y8Lvs0jknnrNM7DJu5j8lFmK7M
RnmJ/fExB44KYcpoF3xxPhK1vYikhEU25ofWxVKOyhnZrr/hTbilCLrQp3Fvrf2e
0vDHLCCyh1hjiXJlVeFZif4QheCeqD5wi6s+/ciWiEXQVGOdkb/v4Od7LkUYJn/4
kF52zOcu/ds5/R1kjePmsdT05pR7GoSEIPOxPCItCWKAI9T7mwuHBA6JTSukyHOy
BwsfybdgD/i2znvP1QSUcSyWeiX4iU3ZSkv8MfqErA3M6PNFgoisXVdEZGX1gJO2
ihb+yCvj8yLpa929BrhBzLXAZyAmqh8mP/xcqfe5Qc4suRp4QEnKzAOttkpO6Zln
1j9OV4t2vWpvz1c9YoP5awog+09Qwt+/jVc6wGngJlAsPwIUZLbiFsNDZit3nLR5
2KtfzKHsqRxS7kWFu3Mskh5G31bA6flCoTQuu78dmwA8a94Mrdnv5M3aTJ49Oxy6
+LJZ/IuiYl6Vn3qY+9ILJ2JY2H1SXBLWInMe080Lvgw=
`protect END_PROTECTED
