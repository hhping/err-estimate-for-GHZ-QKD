`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urculFOOrl0mJgYZ1wfre8vExPyKEZGUZPaIN+ki2iTbmlP1mEOoQ9Ib5A0xLFTu
4fbnkIckg9CCIeyu67s14K5lrGZvjftH74VFBVKozyLwuej3rVh8O2xNo6T3b7CR
uR8Jf58bUC05rfqsI5UgFv2MkYF/uewh6ayPFTioFFHKRJ3Ub+h0ekXI8GxMcIwf
DBoP1k2jDKS9IcOwV6RnXk+F/YYx8GQl8+RWAdDVX1uloGU/OFn1KlA6E5MaWCgm
gQHucau68l5Kq4veUr+eTGRb9+QL5CMhJX030HT59kN4BkI3CMlf5cjHTyWe/AVi
cmOUtFCa7A4Qw3D6s6kN7Um6h9YTp8em9adYAb4h63omntUMurzi7Dxlxy26N4G1
eF8DLarlbrez1ifrmjjK+dWy8QTt83diBpzhOzAkbV12vfmqiHj/yO1IuPT3jnog
s0h05CE8kyI+rq8KX/RnwQamxOPN6L855l+oEfXLPfC8qXbGz9yPDTkdTklBBc/6
tzkYVs05lEmTlxoc/PSlRaSn7Wye2SydksDlozUzX9KobGvBUzFlmITWyYPh5miA
m03n2bzCVU7hUe8ae5lPIT0e3xBi17dG3tRdBXW7yyCCYV4ozkcQwF8pIxqbm+d1
8T4x1Bg7O2vz+sTeg8qTS5dnxxBdvMG2vLvBLmf57uDz3W7oDXv1MJIYSQI+PhuR
5+IekLg0H4N3ZjmGrFlMNNam47E4XVzExpXFvnAfiQYtH12DFXrSbRx5CeJEdqY1
WofIxbBYMIEhzg6YSZR+X4nRlbuHEi/BFLbL5mHJ0D5w03W9rDMgBxsxB41gvQkU
Sij/6xns/A54tAXGkwv67rN6IqSV+a1wECneDz9jV2VaVA4a8YHKFh9/yDtMk7TH
bYpl783TShT0CGGkUy/XyXr0AeDNhqNRceI6Db7PMurbhEkjApbq20NxrK+F6IN4
Eo8g2+hScPle/u95CQ08HdF7NsIIZ+0mtgXHAw2fzBSSdEkybbfu88CIBKPNLV5F
JCoaR/mjuWJjCpOZHG1D6xgtWAghs8/+WMv+wUb8bVw6tEF6KmaP0g5uReLdQLOA
+MfUo3wd7L6MC67PfFyEl9G3wL+af8czQTeqpFd0uW8x+XA5tyFQnnP0jb14rXZ6
uqqgI8GL4ARkpFv8O59df/X6TQFSCjxv2pduYKXND2g1GVDiwQ0fywcr8U0WtC9J
dqpc/v09WC87A0bym+TiG/wNIuoUB8SdDaM+QEVOq8jxJIT/v7k6lsxZaK+af2bS
ZWp8uipcjwi9KhfjemXM89Z5gH/NsDrPBFGDMh7cIQUMCRoOriHLdBX2Qc3tIv7j
PZpgPe+kbDIxpwBKug4nZNRadRNzjkGPJWhKSMQwxhg9zZ2KXQJnLdc/73aL/vsZ
NGh18LhWI+x8u1K4yEtAGg==
`protect END_PROTECTED
