`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1uYm+fOHKkeDrXIui9nilTm4eSVKxqjSMsBNz9c7QXBHxS68IIzaylVpbZZu6BP
od8Ba7bOmCAbDEdNv8dbZGFkVmJwDWDx5wLMLN498oNOJ4sm6GMDZtGDyWzN5UDP
cYz+KcQxbrbpko0WZ+PYEQY9ekttA/qSyKJiXX/v2cGbdiWa3Fh1jKqEQ36Zr4i4
CY7pOsTkpH6jbj7I0idfs9opwP3b0qnaXIXWQFebouv9d7T9W55lr0awxvHZ76ZJ
sOfesDNh6yYcgUCmDH42hmT2mrklJSzmJEa+GWuuNQtnk/jJKRHx7/t+fTc6RVRI
d5H3/fm3i1cKyMKfd4S3pcZ0EY2sr6RoXNlB5/b0BVw=
`protect END_PROTECTED
