`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmMnkgNkr+0egHFLq2yEFFKru3Pp2RAG1HqodpeSW7SXOroZMfhSqLe6rYyu+HWN
j3D7RWv7H5EUoRYUU0i/5kDBgMifw1CdHZW+2X/3djPVclGs6ZepJdfv4OHG2Bti
KOwmZb0ELu6bIHNAGFHxpPzxuLUeUv+OyoANtzn4/HvF9HpCT+3ZPU3s2x6SqpWr
1Lnmw+LrO6TF/jh5T7c/7DgCzoRVq7nZWUpGyFXCEZmgfR4IcdF0UQS19TtaNHn6
zGqCtCmfXEYVYts8xWq3fTW+yyMJ5Y//NAsmWebuAxNYHMHg1sBY3vGB7ddATOkD
gIPIBr1vlRuXfg6fjoH227p68BwGs8oYa6QgZfjvy1ce9i8CODDumxfq0nuYp1db
M3abZGgXYvcTMQQAoDf04rGfBij4gFMRwRFofOXC6BFob1WHw3/mDL3hsXi73Cs/
dNHjTM50gW9eqMUmPR8F6kdYuvRM4L4PoioVyR0RjXYWLFFHVbxBBhYxQ1K30QPv
Mpywzj7A1NoshOLmUOA0TYNvqJpP0L+tgEmFWwiU6r1nZyrevZvsq6Phd69BgZ/j
znXvG+LdDQR74unLaHgBgBMC9pqeDodIkvuH3YdfkeqyA8yO8bj85Gf1A3IX7aVr
JGjKnhw1hLK2M0JhGDLgwNd49kU00epwf21JJF0Cu7aIcY01kD884FTIHI1/SHuB
`protect END_PROTECTED
