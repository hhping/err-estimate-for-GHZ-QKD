`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPmecmqE368IzQc2DaxHitCvhDOvVgSiDYOA8BOrJ17LlKjpnvgHwfBCCSdMNx1X
xTJz4BWbJ97GtTXc6zkosaAMl5JLlekpUEQJBc+ufA/FKlySRdYvJ3PqmNJqmiLI
+Mtng5RNsICX4AvU7ifzj4LuQOeeC6QL40qNuKhmHtttzIL38IQx/wyLQux9p5cP
EecwTLkq1Pnqz34QyApIglBAoyZHj+TusNuG/zFHtIrp4E0Jn7BvYvzygDpiUYbs
CBCY831ypjphGKdRkGPnSzh6w/AaBO8VP1tZ+gMjC9mMR9G0+U9lbm1Rz4B6two+
xky6iK9OjAcfj+94nWsxsom/NTOWIoz2kHDsh/1wJtFxAEtzXJCRZjP2Lc00FdDT
JizbTuSmll9bk57Pr5PeXZWvZBKXgaUmtMiaffkLjDwpK+WvLOaXfJQKumZ63Fj2
705Wx9rRSlQ7tZsjwU9krnw0NZB3fh5KOJbXxcmyD6TZKHa2xP/bzRK5ER6TBsjx
povs4gJvFOV4MGfKIyzlHwWX+fMDd6WTd4fcTDDtorTXiJt/Lu/W5l4H0pDAYfUe
ZZkmkhcQxC7EHlixM0PtTSIongiKZGVPEchGFBtAFxI7UXPRciHHilPhrH2YFpHZ
5b4zKMB7ZTwknwM9b+4cNn4Ot435uTmuIA4emvH3aBrjGJQuYxlWbx47+VV3Etjr
tf9JdEEw5y3oRaqdKiLJsDxl6ca0DTymMrg1mcfz+P/LtZBa8E6KLOif5hrM3u8K
u70OgguL+IxSDF8xyDfZ/hqkziHPLJ+4Td7ur0QOYK+rN+UEK8ijs8eL8y4cWG2W
c9tSBEfV1ynn4i/yXkdacPDyS+Cm6zXpLDWul+h7ZiUc10tbtUZieexZWeLuuQQF
BreeEFtl0/E0Y8DENNnvqjRu326O+gWVxlXPq8KReMTEXtQ7dR89yAFxr3NGaB6X
FUuuo4eXoJejzQsdctnC/TH+1UKil5PLRF/DJTCYqm/o+mwxY3cu1gKYVUbJmMR8
+i7Ch7E8MZT1lfElqGLZMJ2qxI0F78zy5P7norPvV8KlN+yYBI9SQGe4/e/h10iZ
4iob/vWOhdxgUPSFCK+vrADgF8qQNbmhqY6USfqgBepN64cqEmLRBenSNuA4ixnQ
Ip3fpIKVXv4HebU4pTMSnQR6OJEy/YL6pX1+8R99bqIDkoy5zPdnJyK8JYMvujRR
of3JtQ202WwMDL9lhr+0AjlqT55YkNZcFtJrsG3Yaf7j4zDlksvkp9Q39DNKPcmj
Rpn8JmC06oxe+/Rmw4G0rtr6ydVRFh01ElWZUxJlBzaSpxB/xq5SwflWo1SnjzgL
EjFOY1qpna6gume7XcWovVJ3dk/X9ybOXiFiqqxyG0gcZ5BsNG+GdSuNdg2BpUP5
Ijc3rrIa3KvgyVQzxLEAL0ZeABhdwYWrB3B4TXc8y5vCxoQ4YJpnuiXCRbHj1z6A
0zlX6UsvGGLgW7NltBmnWBsfMfmn2z/Pz3SJj8q07CEnlkCo3UVf+tNpwNeTYYcu
GKvMWmauVRnf7YtCMOhM4bbQk2A9MoWWOOS2WWFUct8bw3mLxKGX1R5Eud5vzjcL
CIzHpg5XISUmrhhCj2CZEMHDPzHicMve4AAY9143goTmw6bZLg2L52+9FN4J+aFd
ZZ3NSP9TjIeHjcm87IHNkKUPpeR2LvuEpwN+3W9MpPsoeOIpLLbpW5GMWZPcOo4o
Uojv33mKrg7ig5Rmbe1aFBdD6JwngJaeVoRaiIm2P6PcS7Rm6OinH/JdR6v2T+85
4emYK8t464BcVrVkmvW3n6UWFutPXvHXrScIbJ4Kkz2UcfJthWlmEdTfSwioq8rr
U6nuAbquA5iHFzp2477lMC8XW/voT1anTuHDAPr9f1Uvx/UlhvQHrY8PoFMDaImz
JDkV/RSsVboDGza/v4EuFM2AZMS4UukHoQvNHUbtkea+kD9vyTD1yc4nQuqIGeTb
2lJh2u2pfZYNP3/IwMF8PmRVIK7FjQWCDiWUX09kfPTWWYEYBwtNUuyPNCfN1yxw
qLAfM7t2fSHiCOiJv407wjQ9QhSkEQHfCJkT5WcwfYOaY6Qf3kXSKwJ7o22kc8Tq
XQVPAEN7T5LCG8a47fapsCTs61pY2NxOFQN6eAifLxyMRwjg7xdUnqbMRfPAerbo
Rdb/x1bhMKWYorrOSWkBiJuSTktjOHzcn5zkNFcDiVrPiwjEgsSBcB/tudofwNpY
xbUDLpBiTiIiAif8/1RzrsifFr8L8Fx2EAeIi0uGr9XG9wp+/PNHtJWcr9191eqU
4qJ1C3+QOToBiyT0H2auGB0ETxZWlCV1xwdyXujS+uUcCJ9JIFcETRnBpVGC21Tn
BEtFvQrPo8miBpmjpxpKJbR5PW0OtvFdWmR9WmO/BObXoZFN3RmWn9dbdNrCiPm0
B2IIFVVQf2U9Z1FOPZbrasmMSbFeNtDzTaj9BcoFt0Nl0Vi24PiioQoNeJthRDvY
LU7MsuynE0kEJD7HvTAvK6IsjR2ga5yIZcYODVrUr/vfQYqMUT3PGRMCpxulw92p
UnS3w1QfGYa2pgl1d8bVMnTwKrXBD6Icwe89pklKhmpcp9hrNhYUIgPTITDTZY+t
01TE60b5IdmX8Ml0lS2oLUSw9OpYur8sKQypHacHprMAPv0W57bE/eZPKVfu1LaN
Bb5n//E331xA4J5cO0N9i2bCzVq5m3QzUzsacmO4AWDkblo5kxQxFWYyBsN6nErQ
p+VTR/hYcpjaH8IMs0uqT5EaInCGdvS3yNb0/W3ve0P12ns/QJd9I5eZa19xnrLX
d1199YbREfPGLel43MrLQ9/icTAN0FCFoSuUAFnBMrTmen2M7W4IJFpcBF3dlQgH
NNibIg2RdJP8G66IzX7C/JHB83v2hh8vMGmxWFAiJXuaM5ztT1K0p+ZCU5Qpz+6n
+xtcz5DdBXtgd0/fwTSrUXeuZZ/loMtPO2GtcjtBveYZGYKxVs+oSycfkCD4KNjg
q4gNB3+WMHRyz38AS/MC4AGtgBEVoCgfQyAe2GOyfsPqsizBlje70lFukH5xlqpR
n0VlARCc+QhXh9s7ruQ2lmK0KVtAU4F9c+m3FAmiHn9BbMj7m72UQZOEgK3ig5C1
SdU8afw03yvk+fsDFzhKTua/nxQH2yk/THorAIxdFZqxsALZzcsHQHYum8Ivgasa
2UwxiDvANeybAy03RqnVgPZcn5RGaHFFmZplTgx3fix2yLurwXiqSLE2YUls2KqD
4ndyyfpPt++ppfJMjt/z9LhNHEHJoQAUSh22hXmMS8daA67tR0lZQDlAw+QEV3fZ
ibjGVjUCA3OMVCxk3WEXAiWRa4cS0hYaiWR7n0yrtYFw9VGsZX4htOJbFPlXg66A
T4Ni4PNG07XLZ4znKo2zHcBckRds/5u/+5ED7W6X7gxyvoRJuUv3Ozif2dK8piN+
3TBvyCOhejXzaEwf2oDERycYCDVFanNReozNr1MRFDyAJ97B/KgkORL/Tj4D+WHf
lNtCRmbO0AL0lhSSTaQhWB6/N9DE1VGlblljL/8MUmdVcOT+agKr37oaFV0c1ouw
+Mh05WeIHKlYxAj2xS4d3F9CPSu+iOsz/Wo7nYhrMcztMOQRUp12TLeouAWv8Ugz
cWlVv/R6+zrn9+ckaJB7WZ0kVJcLY0R3kEq0vJ7H7OmeQYFFyyjICc5xGwFE5hly
w2T6pGjmuvvAPjYOHW6xCURWL4m/JA/g5EEeCv9+tYhafAVikNvlatL6bkae/Wu9
V1LWMSsQza0BB9sSMgEocYmGJwJxtvQjbKDnU+LjyNfg/6SoIQGfAPsvBnnam2R/
w2zschRktid2dRqrCM3eTHan70GZFxPIaUDwUmDW3YPOq9efzlcmocEdFNXLPNeg
3qjIOUfq5hHH7JWM0PSoajvzUUqT1lpOrBFet+OKgEEJDF58iWOsw4Ciq6JCdgmU
DiHjNepvbKmLyzz12WpOa9I+t03vOoYCY/AQbI+uaYjTDETI9Y+u4x+YFBpJ2WN1
RTU9iW7b08PvytNgTec0DsTm5YjbDjG/1MsfLDKJYYAK+6kV+NY6tRI3QCSwTWRx
yw6W/lrfLogFHxi087OTMyMCb90ZaNGnovThS/GAoa6uvzjUo424ARMarnjnTO0e
JzXHeghdqcLjzAOIAWqAU4It9jDjFLeV0Z0GgPCbzPmdQkLr9B70T4j85humW0kK
YfqXB0ErbiOP3b5QdagKbrZjI7DSN+TdLFL71GwB6gGYlmAgLcXIv8rT5GMf1E0w
8JbsG8oRzxP08zogVFuM7M1EAp3Nd1ciXyOrmY5rVqEd3ztM99D5kMT0QU1dw+tD
Pf1qNRcP74QqHTBFhXXjaFOig0ByhmKt7LRxdRMTsLQ/rNg0djQytzdUFmixIFlA
E8WM4jLjCbSHcrMiPS3oQwCeDgoRw1lE3BvbAQt+xR0=
`protect END_PROTECTED
