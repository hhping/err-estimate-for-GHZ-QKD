`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
arrCMivJ1NYihX/rcbB1pQe2etnrd4eMhv6pAVoG0DhEOngM4nUd7eYoGcW4a6g5
zO/uUJdawCGYinxWTawMAiS4AL4AOzc8PiXx9muCURRbxUGGk2vBx5nhjt+3i048
+2P6PjThNl5xJRpHYCAAmw+8w1V5qgudbSVaab6GwJz6OyHhm3jDOwH4CH48Z8uJ
nSrhe4S5NwKA4yZpp6lNDhtoWlUAM4sWseJ15Vlvk6w12TxGHKU1NB4mznlLUPtw
8oNAfRmgXpltk8SzTB+OgYREa387vfZpFS3bsOwRy1g0YJYxSlyidDGCL4CDAn9n
md8ouDck7Y5dR20HKdy5EymA+0AyWgRYKZJ6O2FnAgLA61OxFNETa16yXx5RV5fg
i7uxteFn1InfZM7vTm8XOWXZFhJKr9ijB0LmmZUcz+/BRLHjPs/RVekFV97I8/nT
/mEVr59uAeAv1oGHxZgGw+AYld4NgvGEdldDIAf0lIuSzjn/gMPFPr7ePb3Llvgq
XCHL2h6Q8qXMHk+DzEBEBjjm4ycnNRMvk4vNGUQhMWeAW4S+1W5q4hG+yngUbkUH
9qtvd0qBN3PTLem5yOTFjx7jPlUTxl+4wyjGeBDIBkjs6EJYbJhM+A9tRfk5S1bG
W6cpHQ5ikoP7RxoBsauT93NnxM+KM79epgymfQp1VRuo1QNhNY0AYPLMTYhlQRp4
bPkq273aVkiy2/3xrBc/yAZQ2RepP0bM/L68002lqn64+8HLCrZwkrgz1XbuHh94
`protect END_PROTECTED
