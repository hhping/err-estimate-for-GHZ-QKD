`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wHQ1FtWvuoDQ4EzEMLK8DP84eJ8ShYYGd6aeCAuKm16IGoTikObvgCrF+0mFhluH
A/xARs4eMbWegXzc8c6Ly43KnVbN1e1BNsC6+ZFb2HO/qMn7J+pXQLqk3Zq5N934
EUThSW07ubjtG3THkRsnUKFeTlXu8YXUeQAZPVgxktJHivWvDZdB5tOkVJPwjEb4
TRGLiepnJhUOn0QKp770aZg5PIGGSNItuIFGrAuObr8J5E9/AamspVM8/KFEwCAg
EsPMjFtJW1NtZI1knov3qh+b/6/RdR5i3/tg3aOdnqry/QIGWNqfcJaXvAkNCg6d
jmMl9pAJzc+oBSoqZ0fCvfeYcYOnBA4ZJP0K0AoPLbWaIJMLlruiG2fL21IF0CrS
oTg77pXdqZVv0dilzIcqop9T5R6I/nW3zzc++fyNeO5wz+6tY+ouzQvWO+HUzyTE
8Wfb9Djg8GoEM3K2lViJ/4OZKEYE4AuTXqsaFoa+k+k41gB4mhAxcxHRZ3g+gRCi
CTo+rF4eMiuHofTlzZ+MT1MP4Sdg9/Z6s2/wOrjGetZyGz3TsPmUFYLIcp1h2RZB
e3lnxT9Z4UT/hOjX1eULvGaTy3YCGFDabdxDHqEkzlcsCw/vEfmf8lyq8TZG3G2J
c3w/AYByAvWFZSCUcUsR5pG8KmKZdOfDvJX/zoO3qQk7NzwjbWLGWMTcR4MnkqgT
1oR8z3DP1Q6iYlwOpWWn4EOQe3B4JQx95Ei8OQ8B3U8CzBwJBLVLrMJknTcuO4+Q
06sKHTyGcNmdngi2kYedPayntoJ0SB9DuALnt0DBUIS2Ahtevg7/8U4LLdaoyvcI
hs5GJl/IsPqt2O4XK9r4RZbpHZCBIHOAsk80ZK6pITwDTWV3VVJE9N3Lto/bxgm6
EHycZTrgnXCKNaBeZxyoQw==
`protect END_PROTECTED
