`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfAwNXgw+WrIZRfBzSgb7hOt39veRUDqShqmEQopyKGVT8lTm77s0y6gXV3JSsz8
Sc8tvV2uP3zf4pHtu0N5CvadlSmtZMMJRYpepYVWHygf6M7GihWW5WK+XunOwf7C
e6zYmUWLoWbQhSleNM02zN/df7IqOgzf3zL65ZJYwCAFEaJjQUGlgHBoJDCxiIHb
MO5IoV8tIEl2tucIGP9VuA8u5iBxp3MJJW6mkYh9ZnnI4sHPlCxFj9WI1/RsM6sw
FPGUZVa9yEZx1+nz5VUT/cxugofkOVoZwy4C/jVNU6+fqfQPSDJPAYBPdGHvg0Oh
Uo/edX0vnuHJjzRoy7eiMTSSoxcRVRYk9KOdRzdGfhBfnBycBvCiyVTjaF4dj64W
ycDhVMitgMf/mpkMsXgR+3EsP5FAZcSF473o77l8DOEx0CSStiy43dbGJ3JszhRJ
5e22437muuaLJoO45CTNdgatG8prwqk7T0L9hb5XcQ9xVUaNeeHfR7RAlnXx2VNW
dkQIsbKMa42hBzZW8J+HRD1faIP+CtxHPU6jda1IP2VrrBUvwM2wQGnkaXTzQnrT
6IC2suvMpXXs3cDVjshW1rZs++f/aAxnuwEtFSVi5zeqcwLAr0NaPA9x4MFEOYBN
NRz+S+yLozTpI9NECxs60g8mz9ZhCY5X3CpeQzCu9fSlJ2PPjfSqDNF+1Qkrr4IN
9enoTCgOHHdPSfMsWvOj9ejKB0mqMFDtbxeKHMQ/5gWxdQMde6f+IC8HTC9QTaY6
u2HW53e9nROLuyh2/R3wSUXV8eomwvMkjDlR2o8L8AID2AQBclAtz6aJ9jxYCctT
YzydkzvUwZSiz82mP2y9dQ8f3r+Rk141LyKBjd8n7gh+z/9zbkdkQ0ei/GEnB9Xp
DhQaFlcONwS5x3TYxWm+UMDjNW4rdlcRHPZWd68kV1A4uDgcWWqrjRL6kB2CshJ1
9uvoNVA121aj5uTvhtFsAa1W5Hjq131GUwc/dq6kwWbj2OtaLLfY7XZ5PgeHKNYu
8ZgRA5wxEupdFyTWkqc/N7/lI3VOKTnEzD7V9hjjmEyapVWcPLYXVbXFe3SKlNkD
J6H0DAYVGCiN1Dt3LUHiJCA6L/KXj9Z8JaWKDwBkkW/JKCXnU7QWlsX4nJ3zEpze
EOLNgcuFpCwpaJ8u/NvG9pVa/M9yRXFZmAJZoKvMgKiSZahY4tEVvatzugrPtkrq
sgctpvVxmTiEij2bUQAn//dn7i3Uib/T7PiWuKqxPsY=
`protect END_PROTECTED
