`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jfWHU/KeBS4PiSt+2FuxQdcRYhUOQeXaKs+74yisbhDzgWAoPKh5nwmKs16edALI
6RKD901QE0m7tzt44+YWVRCbtd9nIT5+1xmBeS69ChYoMLMuqrXSOCFW8Wa13CxP
wpuD9LWVlWM/w7QHD4icY9U158aUrPx/KpADOc1MHiF1iLeBw3wNaZ9S20sz2oGV
TmwAvzzo1odkJnUp4WQjQ2pG2hjEFVHxXjV8MpxZQfnHj6/mjN+Rj7jtq5lH9jMs
8hO79WsA2sxtFnd9vHAyL78v71MmJK8+KR8wvF2qo06BhY4UMPiKkytVl6EVVH0L
fkPrV3AAo+XKC+nCUKbM6Wrp4uudP0IXVozEiinHJTNvQ19JVJHZPTSB/W+JbFEN
g3fQamrfnyqDNBFvJWkl8a/yNoDPxQCmsYKpiD1OgFkekXRo53sA2nqpL1FuUJ6I
zlcA+Z+3WoGH+mhJaqOJpm7FYfyAZTbV+OmAu+GCTnPdK+XMcMq0CqJ50ZKEx9u7
opOd1A161MniQVAt2JhtJQ2JEhyfjpGaUmeQmqKbbs8hPww7Nh7SJqcu5OHPCF62
mk42baBlawhjOtOFPX/Sfm3c5fCHARv2pnPjfnIgKrph9slOP7BdFWiXdS4HIuA8
HDOsZXw8ZKcV7fmLwzoGO/zUXZ8UR6S1ssodWOJdQj472/8fkHzNVP5qZF2xomSA
SbJKqmpQbkuwlcAR0BjTLz1hBJTaE7ut8HsbWLqJldQ=
`protect END_PROTECTED
