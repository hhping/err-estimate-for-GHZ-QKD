`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkO/vi13XFzvLiNs8AvlRyHpS7J/muE+fcLLH06ftAsZv1n1XxPTnBzKfZuHxEnU
mBsUPlhB6PXvEhAJH1+uSXnUiC+GiE4rixjoDEMB/JMk8ruN7yK7nHAV0hK16aeW
WQv72I9T2D9Guq4fpc3an8wC2fG79MM+D9h0kfpIyY8JPmjZFZihYZbMtzxbbZh9
1dAwilLQ+1qpChCS/YuQjx35qSe2p3DfgEh4VcELPlJ56SThY+9bLXWem38YAije
xkekTqYfsBjFlzlwMcpeJ5zz61s06x3as2nWu5p47x103GGUBJEoJepeqwyahaLY
MK/YbtSByS24u/LEV9TQAf4MjWX3pdMhDc3cTur053Ib6ucovQg8Tla113vOs44p
yMvhVcsUj1a5uxgJaXImltouw/dT+6ZSK0F9rMq7MrL1G3etb52fqa87aRvcU8oS
VMOvBwziR2XB9MFVH5pR5u8yfhWNWbGVF+eeCOkuCCi2SQaYCe4ch8FF6/jDS2zA
8JWjRTz3CdELzy+NL3Ik2d22l0NcWCQtZ8SC1X9PVOY8h5kyjLMmMUFoCPEQQ4SV
qEgi/+i8ETozPUyUHXfantC7wnqISTEftDa2EtJisVsUXO3HPsD2Faode2VIJtCU
uzg5O3io6+Wn5L8SNl9TdP1MtkUw/6v22u8c9jYTtNBK0XoxUEfcYDlB9HjtfXIF
0+YKyb5SxQ70t0qFErOOV2r7ZVURZ7hCjQjWoohUWqcKB43HaTaNP1OamFDrRD5T
3yF7SuRoxPczDe0n93ScgKNyVEXqyly2ITM/6k4d89WFlFfdVX2pERnyWmOCttTY
PVkdrYt2LEpIfqZTHZM1XG31QgjIVhdUaYmYkbPiEeLlB2dQuBE6ok+emOM6O6Xk
cIMcnDcncW4c4MfXMp/UxkjICna9eFL0TeE0Zq2BjXDJ3bLqhOUgaBnZGobP18+I
PR3IvpssHU7sVNg9pDeEGRHzQGG0+HDCxdbdAlTlY9UlVqo2s2ZYw6lhPfq0OA5/
oKtQaLyPf1OK12tdu9KuO69f/Wb6rdg79pT/YBN//EtRpH9mkFzc7oHaqkD4LBfn
t9iJXVLAFldwBFz+4LtxBWyvKFgDaEFbsIWKnnsmo9T5T9kLQuAvSlGJ/NNLmlyI
ozlMOVADGqTJ7rNcw25E6ZeFu5ZvB6sjFVRW8Am8vaGYXrInKbMclkU81oTys6GZ
eb3PmQVk1F0RVipMRBoQTNaEKzZiqPXbS/h4LeyFPt+NQlsCbhYiBCM+b3t6QpjQ
+0BWhYt+wRtiOzHGI2CiLSHV4uIDsz8ZBik3VCaLuv4yGrt7+IMqEAWWqgbDlo2T
O5X1cYzddZ3DYl7hJVmntRsM5FRHohRcT2MS5NP5nVB+I5yrOdhlNu0+RUTLdVWZ
7x8dDVWIq5SYJX/k0iRf5qhzPj+JteWpcrv4fG+8bj74IWzVI1KB7U7C7z2dAzaW
JKUZIsjY65UIdF/VUtGqv3tL472CSCefhKkKVofVwx9av79kJmU6YY3PBwyZLlv6
ZAa6dF8nnY1gAOtMB2pV1A6HGW5AvDiXUdIliPFHK90oBSwAsW+zbnLry6IV5Vff
p/wKUu04pwxUBpM7RT3g5pnpNwKLoKKkT2dYserRbAy4QbElStSeH3Chg3bnHny3
s4l0TcGY0UXTTposp8e/7X//JelBt/XZnkPpDfLUPshZ8vrGh1tMUycvAOij00Gb
3PTmHS2YoqBe/w1xyIf0ZGCqnnolYF16YY9Z6KX48nDpighVdU0FeGKsxW+d6Rw0
FFS+97alE91hIyIHltYqtSycz3QTD5ylhYWX8ufccqM=
`protect END_PROTECTED
