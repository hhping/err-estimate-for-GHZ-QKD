`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vad9bvJHVFD3RCKEH2T6QquVuYtaGvgXPjGjCpyoO9XY+biVnlcY94KDaBSKi1S7
IIRckLju3EY2dSQXZklZG7dIxiHOGtSasxsMaWRbmJh/L4VHUm3jVus0RVf2DaVF
4W0Xly/+S/udWdFzFSv3KCUb1VrcxR5e9oX4gHfgOtpbY+xxY6kQMujcrgJg2uE5
bfKpaeYTcWh+pp64jfAcKnoxR/6sALTXZ4w73BQRPC4k1WCKQMKOw5t3jZfwx6Wb
8RVfDiOrzPGizNZOdoCw0MvnPtZcIwmPc0lYD/SvyzpsQUU1X1+mXFKks+2chD0F
8gmba6yUMBAsuIAzJi0A3AjYypkVIA604Kl+/GrVn1wMAW9Cg9hVNxuXkYOQdovq
Q9+bwjLLSI8DGpTIYMZwmy7LzNwUSJzyX7TX5hDshwUKNH4Rfo7vRsNf0/UuKz3A
EtdnUqDl9YlNLf+v2rQ+jNWJRuTf+UTHF81yDUgrY26XM96iLliNutZqbPaADkUx
pTtdRstP34DQTvsAYilkrO09WhaCI0svaQZKO5Iw6aiCE9k4nWjy7oF1jhKVjEPb
N7EH/k9ipA3oSqkTQHh2kFJjTx3t41dHA5gUrbx4hVJQDC6GNCMyu2E8TCzt6AXd
ZgIBOfAWTozh0ty6iAd4RfiRWr2A9pEzoH7k8BhAirc=
`protect END_PROTECTED
