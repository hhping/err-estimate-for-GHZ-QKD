`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i8DG02sQFHLEVVSNHVrdsjIswZwAGG0SWUXnhjw8tUwAqEaZfOk4S/W85L1Mi8aq
rh5tA4uY4HHtK6Gl5tBroQWBi9mHw+Bh0MLwI/7SdoDebYsaxnW8d9DW1yxLPGsV
4d5KAUoWzLmHCx69ChGu8/ZhqnbSGrdTTfVVG+fP6u7ohTAQjR7cl3wDCJnOouqb
vYIAsWwE7nlXqhZGuyt6lsXqLOB+AXBIeigHBuH6CP+YqDnBOVqhOEg/ilD643Fr
zysE2V6uWpkTXxYUGa3Jp2E5hRmLTxQD8F2NGy2s0wQeTLLP6A0QkOYNcfzucQBv
j8sU5eIdgNknpi64ampkxg3v7KnLxoMPYgVHwHS+tLb8pL4qXkIxbO9eqJ9tojY5
xE81U49ffywSBKU9yvdkVx7lQ9oZSHfU2eEQVyEsLD0=
`protect END_PROTECTED
