`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YHeZEmkcek2Rzq5C8iUst0gNCspQKgYDeT7UPKMoGD3GMqFCA2h0l2ut7omz4WG+
wjp2eY5AJ5hKhKQK1KMxYxODysCunQsxmbGnRfQBKzPH5O+y7KQDyWVz1thJ6Odo
3nC2LVVqLrQXqzoDUtSInxJuxSCs+nPQGgqSegNAFQoARg/zUJ2/Tg/gRf04fAft
vS09pN9zQRcH7wkqp8SvaUpc8Kzi6RYBr3D4KJFIPZ3TB83ieVU+VBNuvEc6LN2N
pfTh2kZPsyLVUMrzkxKHJ72d7BLFDvWPq9nWuE+95a3ZOS1w1QVCl5zFb6Np4hBZ
+81M4MrhgSkjguCHWEKNx2QYbzeY7iDa7Px5bNAyNpJg/5fLBkjjT/zo7a5v95MD
IKe5yyQrL6tpvGUbCBmAyAHG3/VoY2gFuM3NfEzXzvMhZofwRPy4Y13RAuagH8A+
y/CWI35sqpO2rO+Ymdc4jIxrNv+1jin6DnI/5HP9uvwgfDhbyYlPsEhkXLKXp6/1
AEimKDTf93MSmpp4TgtpR3DEsKp+kUdKUEmlijdJUkPWRQKkzE5dZYoJqkB8o17k
Jdt20f0ZqiXorZDqBP94a73YrqK2Y5sW/1TzFrKrf5ww1YaRYQ56Acg+QGtjFHEk
OSFWevvuIKg5Vu0zdaa/+ycRiaFaKu0IOEsZi6R2FGCxUweM+AT4oJF75TJVyPkP
VRSDLcO1jJoxD3DqCZBoqx6f9L25nkeMOdyJHq8Hys9DaWh3QZbNdp0am3Z+OJcB
9AjokU+p9D53n7wHByi7WXcq9qhfQNm8Xyzyg3EhtRr1TxU3WeGCBNUZX59Y8WSZ
TzXhgWiewo3ukKt8ZbXafpnL00EqvfQHIplV30iqjx7BhJzU/q7eaFeespqGdLn8
J9SSMqdU+b3Anf+Zyb11Cit2w+Dx/tD1xpyjQG0JOF8OfaqqcUdOfsWfvoGU1mLh
JixNmb+Oh8A8w95oM/KxyjBySOSxEcRujlAVhhbubaHuf4l6LG0CyKHJ6XBBKYOw
DkBcFApXw5hyqPHMWEoEb1BPRE+4spleSKhP0I9yyXt9leNRvKVpfQRAxP8BHlC1
9lqS+W/iVNGzZgJ7dorJwavAIYo3B0QX5L9mTCsaRN3p9Mitjf/Zl+Pq9/TjLCfc
SsMlQPmaRIznejLhd9xR+pqkAqGENWqCH8cH4JGx5CDyOwgAbqW0CTyZt8TV6eiX
oU4CRDe+ZCXkN6WWQ3uqfOeIWoCCRHMt8UWZjqvol7Qw4vCpo1oTqwIFs/JnR0+X
0Etee9D4P8ZqXqx/04YGmpaDjwvl94mk94n4SX48mvtqHvLvPqUrwp1YMEugG+qU
FOXKhWqL9NuF4fbeF7y1vw==
`protect END_PROTECTED
