`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOB2YF8uzukVsRIcHMTHmXjbJNaDpQZdw2/T/ohS/zg3/17oJAtcukEbHjhJGs4I
KdpSV7+KlhSQJC8QmDWrZZS8wPiS4tp26QS8l+a+xNVQB8/IgohR+CoT7AEJ3thU
rE75mPgoWYiQfUhZgklLzrkXQw8SJm8yRI2dz8vKogYmQUoCrA7Nl0Vr8KFEvrkx
ZJo89FXOxyfeFndWA4YpvQnKS5F4AJHl53krW/8yPe+VQsddpQMuuXKnDwUPYQ7y
HI0Brb20zeJEzcQwECyVkGYyXcNLucjMGY/+QvYFJCqIcyXFBDBoqw0At2zZmTm9
4kFBipWRhJAzR+3syoMFx3vT4Z+oqdn6PYKsWfQKJk/IMIe8781P7tzn3ksQsCx6
QiCiYRePRFN/L9dkHSOQfM5rGot3G1YKZ2WvvH6KYGk54LnuHKlDYjjWbusEwhBU
jRMmtRxmYBTTJFHXDuc1yHD2TsQM2LT+f0ADmrxVCLoEu2ZtqB/aOiLLzeDosRRo
`protect END_PROTECTED
