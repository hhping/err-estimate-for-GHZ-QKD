`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gfpd0der4qyke+GstNC9SY+TPhB/CvuTtYTMWBJUIcBYNiUO9LMSHk45+IeuLzCK
YBZV4ifDSy16eG7t6PoXqO+/dWIggUHIAJ/HSjpv4lq6g7yQZM1KgT/mEt3S0htc
t4uEu3X0iQssMVUy2iDYH8ATJKF4eeqWbq09ghMx5uT1210pHkxKtiLGLDYgbkO2
w4lTkwh5FX5LsryaVK4Ll39qpLo3xjFElkxG2/FtsM5GtNwwYrjoUKljr28OsPZo
/YFPDRusklQXFbYFuZce3LssjWSqLjOSF4eqwUkCaIPa/3z+UmAicZ2lgoc9Fyke
LEjTafYp8zYgxn2WgLOTQJEphtucxAhV+U0T+qOrJJInNzWfOKsryvHs2nCBDDcs
8tW+jBL0VgWFSO730VLk627xQ/cjZNmhIYogDLVOaD9qhMHWewm7INUPd3ek5uWP
/RqJcqZPYM+WdK8sU7bA0/YyeIT0agOSppkQH2vWX+CP202Y7+agU+73oxfgR1Ek
8ADlQzeWlIbN/A5FqN3W9Dc/ryVIbfAREen3c6b3OoEcoRqcrVEIpHZfnvRoDYP3
JUEhJxg15hv86aBnUhzvnQ++/5laCMVNyAekb7oHHB4jrJlQs+h0NCgBesLCx+n3
0bzoOlSmvC58cZmltiUt9aRsyA34oCXfirT54SwJ2AKenD8rclcQNxaSziuJ0kya
g/b+GXlf3f70Re1rx41JvPeG6caUVqCQKe4R3UEtAAuam1pa+J9YyzfNHsSJdHOG
oNCBNFo++f7hqRpQhMsHD3bu8nu7nJEfUiS3/SbmUsISJ5mHQHnzW20x2GofSvon
yFH8zFlKoT3MCvD/UqJByxG0hOWISNHnYupcF5oY+Hv7U7shzt7V/csMI/hAKI6f
yvtTDxfM3+9fuJr4EvNOCA8nWuqEN4RbQ3PoHsWkl6LaDc7aCSA4Eti6HG9ZKegQ
tkogykg/7emwESVSDHeylLLheoVG66q+4XRLafLC5HtMpl7kfjQojFDXMab5dO7p
IxJTKwT/X/uHyalVfWTsDbjfi4DlKDmWDgKSGTN6F/Lk7op4Z5jOIP57rZNyO+IX
O3G2BOY6qpb4PkSzGEZM3zd+I9FNKZ+0lTj1cE2o0oHuSDxHGfp7qyUEB1oWhDjB
II7CFEvyTO7imTb+qT4VXce//m4wsh4t/HJkjkwrMRpvD9I4jPzpsYPbRU8opaXT
YJZVF5XyXqy10IamWZQCBnL4yoNjHG9+27BY10L1hzS0CjcgBQSIV95fPyBCs3Sv
S4cvqaTPtIGu990PT7VxtKNrQpEjEvTXKWDlYzXxTmiT5El+DNIbatU6Dg2GOYvJ
9hZhLy8L3QbVXmKFr2HxCefpq/jayXatN8VQIrsXmOUcwSU375Peozx6Iv4jwOsG
jo0YNMXuA06Zir9FZIPriDlkOO+INwT3Tm8Oo2XQLvD0o+zdvIEVsmD4y902Qtwr
vIw96AklOJTNSk6b+86ufWM57SSlcKze5ieGpMZHvYZai2BYcxcKY6bHAk1e9Uid
qXi30cE3pFCiWhoJWbkad/CyYb88HYO9d5b7JaxAU6cg2N+CkFXP5ylu7xRlQZEi
foZivqvyaGUdz8ggpZQHrFD65dDkhVdTfHF3HZB6YeZU4naXqTqlnsuRgu8I6UvM
Oc3noMPYbKJ2x3sd8gmRw4u2l3LQZ0Q8HZ/f/WVVscg=
`protect END_PROTECTED
