`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJH8PM71P8CaUMY9aCpZEcS/ySDoS5dBepIMB24IWSQdT7tjkr35NNzzCGldHRNb
J2Qikd8NdqGzppqvnj89p//+udhg5RAVL3HvRmoS+dN2HNtN1+k/Da1DEPaNgyce
dyu8IgUtHCxMVREw04TS9XB9Ji6NiDBLpZ3Atg8s0eG11/jKjprr16dcsORuLF6J
bjyd8uDWuoAvifDeOHgj0NyJO/t5YAT1AUf8ukTsWCtyBgBvXPVZgfwITgrSmfXg
bRem3kBvbV7enqKzBjFCwuyN2syVPm1p95x1RwPvlQZng2c0T2VvnMx/fbUvGNAH
H8+/a38+BtQoTKPBV4PDshZxuOE2J8N/m+pEEe4KXLoXK0DUP6CW1PN8JkxqABEo
bmcrKVMaS4kUl0eU9sq/MeGkSfttzQKS2OBmZuPoSTWRz9jUckQDwLQnh210EnUE
9XOZ0zrnzseftLhA3rS7TG6R1nZI+Z4tBk/UNKPDOBGwEq1McXDyGqV5njMxDXpw
tynbSEr3b0a2B8yf0Vs1D/SXEIh9emdzCXB955loNamI7UtRWz24wX1wbx3GsCwl
dtFnH4pJ3u4ILWBhyROi4ktIty/zt8kSryLmZofXwvD6qMbKJWYGINgJnpFSwvcm
i+N2waAVtfWBarbRAUvFB3NEmDIaMHsE/qD7yX5u7SjzvQPNAMpWm3shPALOd+/z
s3Wx2OEP57jQHOk4XsWbbtjYUj3nF9nL6tc0SavYQlLaQRUf0jRf8LGMsyh+rF1X
OZJb8rIQX+7ClclQn5+40NA5nk261vIDLYjSsCig0Xom2gLnJ4Zq06cRIWgloOja
qlqqkUunlcrQNZa+TAAr+wTvi3aJf2JAU/xaZneGsdYFyjQU75EmiEJHuu/0+Jpb
ZjMoujEPs56D6wXd3giG8otEpkuEdTg2jrxDlK7xV0HbGm2fW0Ee28C7TKcftK2i
fh3nH534viR2U72M6uUheS/EIdL0hRorc4lBsgvbeBGJyedbId30s68Sxa/abR4X
SWlbUuTlfzWoOuTO1jypXEfoe510aEYdgPP0v2ieoROHAb7ntno/0IC91Eph7IUm
ir84zjzmX7M3RwOTo1VtSiQHBo/KVyg1LiWKPKd3N7DCFuDUBllWmEOhjQD0S+d9
kH5/UkcJ/iUXUqy/IMOltdfHSSdC95GkEmoEyZdKHWTQU7VDR/njeqI36P+f04yu
B5iH4hK6ZBRtpVUJbLCDi1rL/Xs6F9f4P3w2hcOJviVIqboARwVFguyVmeF9YjvU
kV1z16OH5fka0xu5ZzAGm9k7pk5yDXkCNBAJnHuM4bzt91oFiNYgMCBUrI3tHt4B
QjnCloWmyAW2kizvCM9X7F9h2XbTIb/sb67Uvm5cQn7bfqQzMr9DsKCIyNSGS14S
R/bXb+UltNvEQS6mm5XdaI4siCdBNRyAUXdRUv22CRVRa07v3/Z48wpBWN8KvYZY
WwWQcK6QwoqF06xGw+E0rndoxEG+vmI1bKL9LvRYCs84wgv+MZy/fR7Zp9kMwm6K
EY/jdpwdaY/p5xtzcFGRmVzXID3QvEtiJg8ZE1XyWnNw0nh1gB9J2g3DaYzL+UTT
PhCmWYpREBOONhVFF/jpmNgt7Qd7891ipg9mTKoGFU7SBaorbK+BABtZTrvIgJAA
3GNcYTjD74R6CIzn9wOG9uauk2RUouyHBTl2gGcSkDD7ZU59CSorE1mxMThCuTXr
UoTjqb26SLkHXbes5m1uQl6u9olRRVnrtzCgSVPauAq8T019JfFoa1bH9n4DETvs
8zP2AIji5V86mQPWhXqKgMjIWWKb3UZB2vNRv6ygwTI=
`protect END_PROTECTED
