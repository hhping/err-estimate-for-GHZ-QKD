`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYrycH/HzxaDYTK6G/Oja8AvTG/pceSpq4CxORhBdHJ1qbQ1pt3BT1BtQPTO92vX
6BQ3qyE2r6HxnZWy8C3yDkKM8fj/VztqLuvSIk5xSAQzXt/hOahD/rLKq3Y0jHXg
99vILtheY1egW4gAcNNa6lTt8KliTHgZ2YReKRtHEttWeekYbLzp8caoVPxJQ7bW
U8d6erCGSdCGsbp/wxf9UD/SifHf3bZL49qi4dsZKDsAc9MzJNWs+aMtESJ9ViVz
Yv2ydDZMf/ZW1BIEQdFetTLfx1QAFHj8GCi9EqbQ6++Bta/GYQ3yxvVq1Kbb+zbP
MYwQij853Und9h5WSOVKliVrv6dvuS1yCOsbxlNc7QCWTEnTJuScwMZVBqVJ+qLV
h1pnXVaumFdHkI9NaL2WLE7BolgEdyN6C0h0nmxUFPImam4ctiUW7bzqkyDKM+CQ
s9MH2/cNg9eA9pcocwu28w1gOYWZD6R5lEdHR8ReUNnS3G8cpNFhueVn6yW+no86
bMuR+iLQPBNL52tBoBINdynZa8Y9nNFP1R5D/Ii81sWQdOaU2XmarOx1Y1pikYRI
R38ylGonVtS+J4sXcFnba6CATnnOPhJPpkSb2LdyM4Ylp2dqvD9eTqfCMSz9GkE1
0Fx33GwPr+NzLdBJQxlFTSRWSbmLxXMQap83eZbT+BFjDrMR+rnYHQE/nUr+B1N3
iTy4Q50EDJAZCl6VRDIqyKwTPMbiPq6WQccX54LXz1qoN2UQCaB5aJpeb3pa6FIu
fiFklHdlBtpJLpOAbxpd3SQpCCe6oHJzpFQ7MLkMewDwjsd/wrzj8H4/gl0CnCWF
XUHQquaWLG4PWK62caVWVTPcVwXjWQjiu4mJRw1WxNh9Hdipqz3i1JynMh+9JUrT
FxHiBmXF323e8FkoCEXIKC0r/6JUt7EYnDIBYDe3pK1Y/1xH3wSUKIashDl0SgSo
cqxnD2/6wazq4uADvY5sEkuo1E5ChpRf3meHalubGAT1xekC69W+h1+8SG959kEO
rEGVaOVm4rlvXCTvfO6jVWUY0q8Z33S9sHBJGQjmAHkTPYCr84mMJEKAPcvB4qMY
nHqknytg5V7zQydBbfoDvwNGLGpRqOr3qn1KHeLcrPgCSDPMXBz3i4m3eZV8g7OT
cbvwi2U923wASUmsvJwD1aFEb+qjAY5HX+BFLMmBHDJJmMkaLjg6+2RZgH/wBxDf
5a7zCPX+dtnlh0WqyYOehymD4IuRcc4dOCI1FEAF2U0BPiytV4J9K6hnV+1TLTkC
s+uKd2ERnVxCOVEtRZsw29ffFEGRAP2mf2+BVTqjBlsUlId22jUYNNBqEwLehI9p
VoWP9wxgaGXpjuAjLVCN6G9ac02D39L/7+Sr4pOpMtR39cf30yV6wuUTMWffBKao
CzVxePpuIqMmbchKxH9xMvDgXO0kfO22ajWKXcpbeDko+1s5ftCvjsVWO9q/eB+f
kXkRg1gBIktugRtEnSUzCncpmZ8uWJkZWC+YBVtw/mfANfhORpwcCOMX/huX46w6
cD6LRkmTnrISNT3JGXqRoQHoe3pS74GGdX0Q4vneTzb+m1MqicdcDN8LDJUeHg3i
kkIcvgVuUYSot82Cuo5+MkFIHpXKDqUaCNLlMrLd+6LvQzH+cd8hDX96vS4FAXBx
iGL5awZMa4X538Li4kWJiO1HLYPQgulW15GisMsCUaK1a4K1W8tHzA46JujAd/xK
MZSy1xGNfHNVi5dK/zCeRnvvvSBaOK+Ma2CTXmTDuPWDnwzdb3TS444n+4iPsPxF
pAhTirKvmamhoDB0OnA8tMvr/KRMDohtxP42cahMmkvzaFrhsp/Cmza4vVrzZJtb
/9CxN47yyKjeEPmbfq22Gb9KQqfmZQs4VcCfbbLYCa7jhF87oNJW5SZvO6BnUPJN
Fj5LWxQof/eJoKm9Os9qAwyRMpPCw4oIfmhmB+x2quRA868lTd6xgI3uOx2rmGWR
24t9Mo2B5BELIMhpIBRYQk/g0Jvd4pabxgVzN9pKyjhn9qrBbJGRT2oqFRkq0O1g
5DJT9TXsK7dlA/YeGPNtU7CY6MrVNqwF2GsrRkxk8g7Oi6SiPVEbH/2rXL6gunrr
nVnwiNXmhmrplm3Zp8cgbw==
`protect END_PROTECTED
