`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IarEwMFJXwqas3pRrpnAxP0AtVtsdInEZklem996nT9L5vKiQFfqc3qXhuJ72NCu
xSW7JrlclxhP+vn1DLBpZt66TJbfU5x4iboJIqHigb5/gvh5JqGvtqTF7BQIU8Qe
wndSFuqr7dCQOBNNaiOD11FrUpnNjiYsECjJEWLzQNO3xMJ/dPvFKK9HXhC51/Pt
PBv6YXH4CnPcXzjf7j0btCHX9PImuQvyPfO63ngbAWG3jBuJM2Uhrk0/EGljs2UR
ZRv4/1qbPBl0fyoNqPtfVkjeJbbUelr/+9H2ZT7pWLaOoWHdfVdMSNLKlV5oDzbh
jHwECLMepPT52SLcvJFjeWg0C/6Zi4XCeChhWJHKqYYHT2NAJvp8KwKUuyIgsLEk
eArOrt3JVM8OIhoM0+i0e+qb73i3fxycrxciL7zHwJF6aHt8uCb+zr+P546+F57O
TQyUsIOgcLtikX8RKpfonGl4V2vGgdn16hSC0HrTelmAosC1+/hvltB5+4UYdgWM
or3MQWl0I6+JV85ZbCsE5/z1S+pJVgLFKkoSnVUN+IJgqJO6v0Yx4WygcDVnVY/d
IzGob1uusZln2BdrY0Pkyg3h6YVywhfGImI/sNVkZXB2gRZ0nz6wbg4VFhQMKzpu
`protect END_PROTECTED
