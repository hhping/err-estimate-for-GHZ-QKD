`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTWG3EvuSIr7/sfWsNwtPBlSWGhSAfAZdm25GPyqWCeYJL5enVa4AHUd8HqlWfSB
20LKEiTmZsXFhgHjc9c2qK77o3T6TGiVEmdWRT194DEj9pJmAv7HlfYExsr5Wdy9
qX4aip9d+C10eUm5p9wRkVhmyRNn73uax5UoL6CDg1KVdM8vSVk0iFg09Iczyz9q
HacunKEOyETTJAYCdxo/zyXANJoVVGLSPkmfccjCQYxHqdOLGl2alM8gP7WyeEZk
yQHWSqceVcU6xwXe4kMZ8dvXCKa0sztip7yqqHFmZOxB3BQIrh9ZMoqjqPaUMW9D
v6bdoyhS/3oCJ/YSpN18DxYS15uOPF9pZHpYmuh3Ndkd+PiCKT0uuE9Qn8MPiHXk
V81zWgSbSofmkdl6Oyapd+/1cr21rtVF4Wbni72v5kHhBE8TkR8I0wY+czyprkGj
X11QUXnM/feIqkaZIfAgeGmnZKy5xcNoeDFYfYYefJgsnEQP1h5WBl8wZjUiGzSS
b9p3uDGJyeKKwo7jJvQrqwhz4yitYXXTUHwmk8jrAbNnlTr5axmKK76zmDmdcm3/
hUq7CSLAb7WTUcpbhJEs1pgipKdii52N9ad3GnV+BshZV+9C9CS578D4N9gradT4
gNNfHa1IQGPFcBYhO2OSz0gDvJkQ6lJtomxjXklNgNaVPqVjIJ4k9lBP/iltgdJz
fYDiVEAMHoaJ292zX18ikc9USkx/4248WGtF5v3ARTZUjha2c1sSwb4O1hpLGxk3
349L3zETbwhVi6WIm7b9hkvzJgQJuopCDsXFtw+oLkdfplRZlBRmSc23h7KJvroR
jSClymXW+sYAzfPp9dVRkG5glsu3Zqa0cDNA+j6xVuimUzcvBVe8m/IRqienmfbf
skfPS/xfdyLodohzCtgKhLxYUx1/dyFtvMheq+qVpe87ROyF3t1j9D77+N70N/7W
lwFfAW1oUjZ4pysb3g9j/dY2BT1pVea0/IpdH/pvDiUMJOvYvjujNNwbgV/mvc/z
L6BRWwNx2l9tmV7//wU+O+QYuxceWO58qXVPL5f7CYzdgfgvQxkauRhbrvpDffzy
fBSNpeOi7CseB597VMo1DDVt/JW7e8g18bt/ANBNgolGvH/YbRNbzIlJstVEPMHd
S6eil16yWEKOApllY/GaMOD0Xj3C4Jhc8UoiomXUpNZPz6EVc390BXC59DYW5UIz
gajMicLRu9FZyFYC94MyIKWqowO99eS6l6y00PpvQ1Gi9Zjbrq8cfBJf+2MDS5gu
ngYHm1XoiKg2SiGSWju+t3tWrSctLneMxX9nUe4C09C7Tau1kEvHG9QNZafxHVCE
bQe99mJvk7VRaBKSfDaQjAn6Z0SFgQKS8m+VhNduirOelfaT0LzFHZR53N/yVov4
y+A32iG7peGKRTwZqnBXerQw9wE3rTI4ZfaiBty6T6YRufOe7oXowLPBKWwhfvKM
CPcjXLQpJQR/TvR3Ub73fZ1axWHlDbJGJpN7nqcMhELgAOlcCIGA8FxUtU9D0W4l
vorjUZM54mhBvga/BrvSwddCoXYTO/GMzOWvTVv5GGPOBRk08zZX14iLAB2dgsrr
wL9KkIfmU1LzXEI0kDUC92Yjbw7TDAyfHdjeuqs4zBLHF8Y6xnakw3ukmI94ppeH
g+YbL5cSs/agSWGJlW3xju0K3bNejmUBstmHIEZzuOBoLIGj1zKLA1qEzQg0OsH4
rfiFqx6DdyXFOz5jfLGpYjbKY/K6btGngm2LRncz4WYAR01DXdmjonxM6mEJyTsO
Vsu5rOZ4F7o6kRw0Ma5uxN50vzdm9jSzKgCfhDKmSTWrvqKFqYmQ7fRKSN8LGdI+
CcyP8XuhTQqZ8utRD2xi1I4oJg9WlT/7mDLFvGoPydSVLo2b81eefUXGI2aEdoum
JrO5winOOL5Oqn8JXM9wnXoLe5ZuXOEwZB7LnVRvRxk+uHr+caI+Hd6vhojWPRCU
7IU5Qw/3SgUE9gzDYJRrUQ2r0A+F2ril7X2hfk2z8w/Vcd8nt1rkZxfgxKvObg6v
cXwBWD6i5tYWqSYK8xs4YwAsSbU0e97V46OVYOO/8eETANb/1VjAlY/ROmDl+YA5
O4UeuHGxtwJok46UMlxnR3IbxeqH6zPnN3/+e64aAfo0NsxR1a0e0hi/pwRfKd3Q
TqLS4HfSxZmoApdJwqq1EzEw5m3mdnXCAnUPAtQsrDjV3yaT10Me5+kUCkyliv04
j+Nox/nA25ZkDCw9sTQ7JrnqidpueDEjps/laHnEtTD4bL646o44CSe7QYBE1Igb
AcRGU1YSAkTSTrCtBACJHHbgjKtKJzxHZ/pgnxPBEoI2Dnh1lvJmEqh0/gSHxhm9
dPKahlbV6QC9ghzIHtagheFHaA6q3aliu9luvKlOpKxcPQaxdy4RfgVMV43JXFEK
tnkW6Z0f1noiX32SEVs/l01SD2KRQbakB/Fsj8yzaLfk0lKRLuiKVg6YmM5dwos8
XxcMoOwKrynhdYVdxELKWWQSy56NSzrxe5UdcY04AAycGXPphcVT1WicVBoOSsNp
8gw5+JlW0XbwlsROMxrcgf2H9vtJXSA9BIRkEzKNNjZyNnhfO6ZhjibtnB90Yz2u
2z5X2pJu17ny4vyVOp2WVx72GmpKRmH45Is8vMI6HnrI4+gf7Zt6LHbNvrXxTqew
bR+DAMPmZBFOZgbwOtM9PKml/jYR/bd8Ls9AmpgCn97QRC2B09E2t6XkP5ypKT3y
26jGDRIQTnjU9kLEIYxz4wUtFP5/hrYimJkcsA0L9M4h+C2MRbWsOZs2zxyjVAEe
Xak4xVB53qxM5gVkcho0v1yvu0/b6lb6+6BKhhB3vccqkJpUFByLjy285Yd3j1ms
r6F5IidPBiQ4BA2bq1Z9m+mmtrjI/MvfvvLG9IzxyhG4UoPIjP6zMPNqcFr5Pe1J
PGLRHSgFVfg6+us8uvP6ofBws+UerETFmR2nZe/wCY05xogmCoa1EfjTWtkjKp8A
XhqHhs7LH78GEZzTycnaZPuqiuiuBj8oyYeq2xfadHmXRiCX4AJlmKLYsLtyLLyO
q+LI9PNIbUdKp4A5TKG4+Psl86g45NJf1QN/yvT60BPXqe1MRCoZhSx6HZhOvBtg
LKuRMcJgyVkocgyI4sxqM58AfVoT6WQxt/PzUmDbpOIvMAoVzzbdLfQmQDvXJuOH
4w6OGj11+qUXpgk/8x0KuAR4dQmlZ5GBdmUzFcDGSaYhlFPIkdUXelAJDKTepXJu
i3eqE/ZXKm17MiT1zgWO15gPRyvjxCEdhHUsOiMHM9BXtfy9UPM3e+X7jUXzCCGe
ah63JcQX3fxS72CYqRVDtpTLZS/7VVd+i4U2XdZN5yBADx5BZIklfkHfAWUFBfrk
jFQF+8cKuPJ5eMcLvpoA9aSWC5AtSfMXkpwEPEuhC38pc6BE6bdb4vm7FaydFiof
srfdr+Q6gDLsrP1sIQxyIYgYXit1yyT6WbTK/LHFVLlQ0JFeXsU4dN2QNxa+LOIR
dW/SL78fi9F6gS6X8jWhlIzsj/R1YC2vUeExvIS8Og9Ve6rL5i0DG+lFq08o0S0o
Vg1MyV/RIk+5w1/Fo6IbKACxMQLkQEiTuhLR9hCNqBNvyAom5+We0Swrg9mNKOM8
xCfITyyf4MeX1dA3xc+8C858Ua7x8+gIdupHlDbNtKdvxuPcwIWRKoUI2nixwqWj
rCu6DUgjVqsANkdbYLeyhmaKZmqkWphVUUOvJxkeilBZfGetRRPPtxqkOGTAigxZ
ANfB+hNMNKAEcILMIsom9BzMdL6qvyr6TKrd0mgsjgywRr63yvy4Q711oyd63w4m
SO7rZlhLfrpr7XhTxEWpSK99wFiSADJkbWUPsdQOoKw9e/qYgcxq+ZuImSo/5X45
mzeUV++sFa6EJjSGZu4/9YW6KLI5455aTiz9B1CXi6i3qpLHWVlUhjNgq8thKAo8
czkvBLMy+YLkX4UKKoMqfs6I7gQF1DLtOo1XY96m8KqkKSC738V0kFcwho5HsHsp
bQ/z2jOXLnRj38NJYQ2/ZXPYY4k1ExZN8fEO850FUgq5FNR9u8Iifu+2WnVlyW3R
2yegxEo7I2WNN2oAiMpaaJxaitqS4H197eN0/h2llUYoVpW+WfDdldSDGdClmZok
p01a7PrXJcOcUEpMURw7dUSNKY2t3uM6EeOXWU7CZyWSKlfx1N6/EKZLJnp7larS
yoqmKPt8lT9a+nx4OmKJMKsYVsWzGvCQujzTfGQ6ZSLXh1lEcWW7W0Tq5PK0zNQ0
eSZLpzv9AA/fbt7LifFpnIMhf+aL0Qq/I/cizrOQEOc5rJY4yjaDDQvpHb4S3sSr
KZVuKnIpwzhhLTF+qqzoz2Ql3flrlyJD0L4GN7St3NWR6JeM98k/kezzd+orhiJa
aXTByrsvjkh9Gnnu1cMxLMx8kxDGVWuSlZ8//pY7tQLJNYpQiv1ZqK6HTMpeD4Du
EfOnwXjrqZx7S/to7IiDwcHYK2lWoEkhKrg0R5GGQR5O/ZzqAgGxIyDJrgR9SXow
8EKty39j+lWN51T4w6X7T/LdvzV26M7Si1B4yzeoVQKTpm/sXBQsvNtUciR5aKGK
rMItrEaLLqOpxo3AoG2hRhiGyki6lbKLDIxJ7kP1G9e58TDOyW6oeVlzCbgO9yN5
M61+P+oJC/v608Cb2g/m5F5bonIXIdB48MmmL1rVGqDrnfAi1ARStJFITjXh2UjL
RvmiOHwPYnk+KlzYlAPSvvcjEgf0xd3o5qUb8i9mbBOQIxMFn3YKLSarwOEUkKCI
VH7UI0CpqtMtq53ROECnufc20isnzLA0MmCMfHZw6BM/9MxcLG/mAN1JyWkk0ViC
ZXWtoOReusEF3l9El05krk9aMC5BUoz28sncU7nzIqVtUhQJwFv071TrwSxJyUAk
Mm7WUdRYr0YsBFol/QKbMj1Vi43MuY7fynP6xdf0N71/8ZoTAcFQRPe3X9Ir4aRL
cVxnUUH7nC1u5g9YJHYg7atNPtAZNdeGV6cdGWiaUEcmWT+uq9L33WIF/FrBEoBN
2EXYP9ghf1ab0kJ2Juil+A09RhXHy+CdjlTEKnIJ+mOoE0oqiFTLCi3JRRKwU9Ip
f4bALBUPDjFzo/L1AhgQLRxxRoBmI1MexIVo2+/sXNOyGTgKdEWmPYOl8RjSCKut
hVXtzggr3sQVg8etroE2bX6aRv4oyaW/RrZCiZA02Zssz4jBlapLY4i79n/2a6rl
yxzfbsjc9BU2waxucDpb8lmk9mLaX2koVS3NQwIbPKFrrFUyaYKJZnVU54JdTY86
xK2Tg/Yk/rqrZcLW3WNz4Dby46yzliU9Q6REzNy3X4/P7Vi3C9qXC4FPyvb2iEuW
vQ4rhqXg1cHkh3BTOXaV6GnM5qALrvc7/7niMi2KkqAzDI+dsI0Ovw4EfKGaCZ9B
5U/LPMFgJtwpmNSVPNmD0O63nPOO+2cQ7Hwq3u+KecsmdwPqd00arHaHUBdWzaNY
epbeMZTGySo+sNRpJsL+32AwM8Kfs6+TpDpNrNPn75zA+3cScwlN+FxE4F1u+L9r
ogJNkCZjFMgiNBu9KYhOeWTEk0bmo5B48yWGmdr+qviuQk3D8s1XYiHkbxmkS+VH
PmBI5cVoZwtGhqiq+yI536pMOSsju1zq7wzQv6FYR8n+y7YLK45UzCOUwcvbEasz
0tHChDeqGum1m/HAgI/MLiOIeibW5QmtfyLGCuFOf1HuosJN4/FLZWCd+07nyMA6
9QgZJT1M1QC5wKapjeMs0INL2OpDoh7a5TgoTPj/2CEdSO9lcTjTDHhKkBp2Lv+u
auttWlNoQr/BgJYr5SflRHw4M1JjhvnUt0uDrJwNK8df2RrU1jEePTMmDS4XMXpK
1cs+UzB0z4VYxw2FWJ9ZyTV3fDYgSvqRYlSmpwhTYfRh1TDyh1fW3aGME39yNPFN
XEw+8BVJC4gRkfbXzdFitXbG0GZpdXfcDT3eU1x+fZ/2rd8mFCGF6cIC0KYtSTm4
kD3eed5gDh/BxJDRc4mnFi/GL7aomfLPzhv4yxf5mXvv/Ztfp6bjHSKeuJqClJkC
NWigtWeh9zCHQM7y0XTH+mxdBsGcjK+gly+TX/xJuYu60C6HTHl9EfWCq4G7+f2/
NlqYVqPJfFvP/8NpaYi2aAWgXcK857AjuoOXZmOXxlosfpCBGR+Y4tUbVfZSRVx/
C3N2HjAxpvv1xlj88fiePWSEsp7hn2JmfBfVEV/fJdeRT5q7HSsJzdpHR2ix5IKY
e1I2so/i58zAgtseV7r3AjrJteZzPpyVH5B60uL4+swXIdyLaBqR8XYhpR5bJXU8
Wrt3mbQyFgpEgrCikVFAYcXZv2QUodzTHcETjb+K8iBDe5OtRcyOOdP6HfphIWd/
k41B45O6+FeE7g16FJp9FDRwtg/X9QuX/GNUQoEyyL01oiJG5xrkiEtJuLLEwLc+
nCU5+z1PirSlo5fBWXtw0D+y2t8CSpFTHMpXyyckU2y4ezbMIlUkwjcyOdbo9rwz
3jMfHv/CE2Bk4PevpCp+MgutWelPWUTMk2JnH6GtPSqgVO4H80bAn8GCuOEsH5eB
jv5ERA9C5hM2J0YQvSw6GpDBqmGtCcK63sKwvA5lpX8HMCZafYImyF9Dj97fK0kX
6PUKJkEBEZOX37AtWzJWDHXN54UzWnphdbB75tJWr6m9ir30809vNY+Z6ovzfIfL
TUFRx5E/txiPcLshb4OxdYmiRT1JVzv8iKJjQFl7LGWdarhY9KiYh7UJW3TCLvp3
v9Xo82y3FBnPZqNKVGnvq+bSdqkRUM+v8ic+Z5244WOSPaCdieoIJdzKdOiVSJX6
BnsasFdkGIj8iMmb9pLVukjob93Zs9BSM6YwNNvxA1GbYaNh0S8ao054BAp/f7lz
bixyGyRD2t2+KyGDVU7cX1mQRNw7imfWWRVsir+SWkshW3cnksmYYU3OniUujJHH
7ffAeslw/F5Ljcuepb8g+5XYAPe8/tQHTraKePElL+hk7fCTx2r0xJo8836rzkZd
JhM9FpW3/DXicl3yo0HTAlGPVPAxKhEzXaONw+eubDFNt8Zf5uZfdyADKiKjwltP
GvQgqkiNETXNUumQR4SWXxdFALDwCfqJjBICenFQfwTntLfNyjybQxuQQhk5nPy2
Yf6HSTYJo1hWPngxk3cGK63Jp7mcZBDTD+4BMiRy5X8VkrUcFC5+9cdugoA45Rf4
fEMeC6PXDyXKswIkSra5iptuUkQJ8IJPPH972VBhsVX+p2P0Tgae6nLywHDYvbBU
+rDtBH9/oMX0OQXMYu7Q6tSj1F5KIO5a2L3QKLEY/3LzlnQmwjR6QLdx6jVLztzE
JBBYUx/Msp0l1Fs27k6hQEQdWhrOGvxt26MMeBxUTfwLrgP9rNQr5fnKvWUxFfMy
P7ATyBwRyxTzOCj9JIAGUJ6hOSrv7vu+Iggf9WxN5pyXdFdow8AiSouE2JHpXV8m
Zg3Hkw5CipsNN3Tm7JWy/kZBVzwvT+VVFl+7v9QZrZYMAA6ejO1jlz21sMyPeXr9
yTT5/wV083ZxZ6qFg7ZDInf6kk10dd8sptef13PaUVWBvfz1mL5F/68g5fgE9q1U
BrG6F79h8Gk8Bbhzrbt52tWNH8x29uJ7Ppgy8KMj23o44ViDVDRnmIChLhfgTb34
7inEWtRFZ9PkatdnFNvzXCPpMcTGZT1bafIRfS0fupvc69CBO9OwxpRFGUTyFL0E
aJ3+tkkkvm7aIcxqelLsyaJG9ZBqBLLv3cIrrhFYAQBxFUVya/bypftS57FRwxYU
vnjjVfUz7OB/wu7PUFiIFbILym07m/+Cp2i6Lf2ZRoM7COcleeqPXhbCAtNaw2Dh
B+G8CFpsGVB0uoIDoSPaRO4pKUkwY87HiOe5Ipa5CKf7r4y+vUfnwpz7ZhOjO1Gn
j2ktzUYEzgXZtcgpZvu05EDydj7siVFP/sygRns1NqvNo9a+x1CmmIco/6Cwcf/d
oiNQ/OriHVyQkv54YVCBvHbPJ7UnFtaLBEmUIku/p+DEjyX2Z6ygvOxiGtagOZla
fdaBmlQo10lZ1u88uJ5rqZBaxpwtylpJpA1wwXLb+noDUhjBlH9Dty3fF4nHcReS
/K6CNa68fOF/XTAZhOkaUV/hCcoCX5SXaXkDcIDb093cQpqWpmq9H26E9kszb3+Z
HVnlyB3Tq5kngP5vS1BA8bs0DHopyPa/dSFNtCeUtEimOUfViuwzQfADN297ZcD6
gB3QEab9z4LdxluxG4FU77lTmQSBPG/cV2+A2uqfEuBbWNdOr6paBqlb+yatyE7U
6tymrbIrRqiKHeQ7Yu2ok+Zis9ZG8k3PyABu0uSoC4KhMFNJ87+SspYE2NVmZMuf
2OjmKqkyUhYmzfgILVh9WX19QZHCL3r9OGFx7qciyz58jfWr1Ix3IS4zqz9Ju19Y
NqleJelgQuJ7EjJDdlb3KtBNRxzXaeuVuQHgVC0HyyU81Q1JodgBJhM0F5uTVAOk
GS33GfrJ4Trik83kS5UQVAQweh0hLL5sL+LVjISfGg2bvpzQ18R4IVjyrTCyytUK
yhGCijMesKKgq6aTDlcJRoysgzIOsXM7Foai+wmTxKwsSkhLi0G6c+NTOZQn45tc
nn4quHHQd/gM14iSxZFGtloyFajh/L+zgn2kCYv536o60H15EhLh9NU9MDKpwami
cjYPyLJNpqY0fG8ddAqXKXOT0/0htcipTHY4jsgrE+LDAETat9bNllghpR0PV09M
46grPQZmWjncxHzD40XM6mTxdxvR4uic4eIA6svDa2CU6hvLdE1MeVIghBulA9rW
FLWagghm1fUvNCScA/KBg/ODQiKiaoUNJWmfPU1y6XssZBLfWt06kKhisCjTtQU0
D4q8RMxHqQ198COOXLziea4/HCLoyKccAEZzhpnQB+h/vvXxKpYxbDhOkSH98915
MwiuEToQryDvoF3CM1OWF+p0QbZboyCf8nEgEdO4HduaFs6+JOU0B4rQJEsiXSTU
NqMua7F4qH8YkCMz4LJRh3jQvf6whxI/uD+cIjh8i8o=
`protect END_PROTECTED
