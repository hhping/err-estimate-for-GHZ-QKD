`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6z/jUPnbsNxF9QsnpfZebCfUj1VBd9stpdt9cFGJtTMHWJvdUFfAwrMymAt74opL
KIyKiyUOxdNqmYRXyK1E8h9igt0jZqdU6nxxNwkmvEgpwwMxgWYH9jNvjjo/R1p2
iPKlIMoShPvjGgZKNQQmevTJ6GnVMftBlG/eDqNic4/Q/vM0tqjNJ0QITRIimKzl
SkmAA9U49S/mE1puQuucdUgkME20TFrVHHM1Ce2k+BuTGi2LF7lZ8bqymRVFgEM4
Lz2EWX6a/WkJVUgLjnqS/dziLuEjZgjzyyvRTHHIdLPdnBt4DgPQNHG18+dv6NnE
z6gOPyT32SO11G2YiNqNbffQNPH+w1WmG8vcKGApm7yQx/TVTYyc70T8ZijGNYFY
LKYTBtAi2G8bx8OAMtlL7tPyRwa4D9aGipuN0+3z5FGE3zDzg1gzgE4kaS2BtQKv
8HKlcXQ5yfKrtVz4vzjpyrVr6R5NfC8cMvZ5nN5W3aJS4Wp8NEDWk6G9Y5Rl1bns
ThvleQGlcDzXXrqDYc/YQcrtGPMbJnjuvlssW+ZUEktFkGYukyBei/jvfyQYvl2O
WJHBzdNoSwiTkJY8c+5CphZ2MLcIhmjYO3KrMdVyaxjVqs5il/k9rrPnKD7JLPhL
0x5ayLfJESSvWulEfRkoZixDOlq+XmxYehGVL/rfd9ipETqulJVOMS/blWa+0aPB
WgAY59ZeyUGL4mwCo62xx5o6LJE/PJwXiJosKAGVnYX32Lq2eGvirTiCaMD9GJdq
xHKxwbi/eMiJIgakn/fRtgzcqvLiAgRFSzG0euabouk6ytA8hnR2CrQLPz2NR46o
ddV41pctb/yZ3Ky/WcaL9XtWUsPUDNwkCya3O1z44GEv6UYEEpj2+eU/ROoc8HmF
Pbx8exjeZ+3AxFsSlGzb7oKYCM/oOjYgP6JX7yUa7nMaAASLhk2+k/7nMJ+/SIh8
a1mKRAI6SEPrcJpsZqbvm+dA/0/zRBoPmfJ+iPFznJYmCbltGdflwbol4b7k4Cy3
s/6V2hy5wNnGzgRvnpX/X/9JvtBlTlUnEde+xDTxprMSbfmMydXrT2F/c7atmBld
/vvXxENn6DekYSWZjiZQG9+8+vVyeccfeMPablgBwdU/u/uKKcwaGWEaIctx8OhS
Pdd0MZDTMXZPtChz8vm2wpMIjAE/mffqc7Ycl1XZEv0nAxAnBn/NFVAj2likACrD
UKI2kLUV8wf2tfaprD56KHPr529peeGSULTztiLnNMK9EPLT/Bzn7uyCxNOtwAvr
Q/724oxVag1zWmhchDYRW1YKdzMe7yMHFWQuyX+AWAkuwz2xIB/hlV0zKMb5to/M
`protect END_PROTECTED
