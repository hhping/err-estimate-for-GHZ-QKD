`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nk9eFHB1e/7a6WFw0DDvLDemomijJEiK3EIiN8xbUQhsC5qFMOf6iu+1eBQehkzA
05ECzuxm4uuUW6mUjE+xQs0fXrBa51MULk4Lu+lV/cywr5vdUjqpxBSVvnpM8lfc
uJVCToUHwv8vA61BtHD3f5ml+7ntMx4kdIccVbpBwKpWweZldYK2W6gcBdipa6TX
kMqPVoKO8n6py/77YJD2+uhRDfCYXjhCYOd+6WcBvCvIvzGF1ziUFbN7+HPGgqAq
sFKd6z/E58sKGQhElQ6B4odi+8++6WKQ0lSi1pqjxmMjUG+8+uNf/DwcEiXIrcn7
SunqM1QNCaA14UjpWv+BhRs9TOIDhdCkK5n5V0TVE3YcmoULHjUuQnpOgMX75ucT
dqu0NW1ZlGmohXYkzQjXt94ybd0PeZuiy/aCq59M8+/S0Ilof1ilhuTVBLqa3JBO
dYRZceikiGWmznbYuHnPhy+6quaurZJmC5WrwENYptSxGLQNh1LEcJoIh5ILouPG
ov5x7cJBc2geWEhlpSwhKlm1vrjsapTkVzUmttWUOFQsAR+E+j0EKt7NXmq/90HF
bvM15dF0yNHvfAgwzCjtvOsrUqvx4ShxaZNq0dT0+qNuRn20Rfi4+7tzRfy4/bcB
vZPNHSvFwin2oGyWRNcngaR1Tf4yzdmM6bC2o4NYkRRMKir3sCBY7a52jYNZ/t5W
5EYAaQGpi3WKXWR0PnwyhBdYM02Mbdyc6svCBqUExkwZhE8TM2U6RK1W739tgNgW
uOasRveVqq93rp0SZkSWjNxtQQisV1RO0rd6AIX65Xl+1GzWSGcR9VADzrs/BGTi
S1p2HRVM79UgKeHpwBo+UhghloisHFOBTLI5bcTAC2zQDlZvYh0VAUb17uDoGZDw
yA+Nhjj+x/KK/njJkz04IZ4xwXczjAeKIJrZE44BgIkFno8vd5MB+LixRTamSXBm
+HfjhEdr9JuZrKTdx0K5kw7JpogRoz2dY4Y32A66lFw65Vs8ZjhoFEu27oCtSSMD
k7cqiI76R9OQ1BwCjuSnddcmd7+q2VPV8XTxZX0VoknWrK3mXEsBLOCCWasZBPrr
8/Bz2ysrE6xPS5CCxy01sTlyq8FE17JQbuofWKcQGJg2wcU9r0PZmxHvhs+hg4X4
58DJZtugsHEdzeoAyGTUdOfO7ux2eQ263rWZj6I5CRyo9SBP2c2EnrSFIvuHWpLi
wfTbjV1ynpO3OUh0jqO5q+Qi8Jm0Ia0Pjf+ZPFqVuLQXzRNKx3gBxvE1rkXt8sXi
hZX2+3RisM7+4c6qj6WiyuxkQTT6yRXm3bpb/B2JhbYqZ9Vh7ea3+UPtMYrjVDEW
AJam6N4FL2LYqyFmGG5gzcTWb/K4mVF8GbAvBqHhqqVYXFkS1EFEmMK2Xhm13NVn
S+w7KlJFobQ4j2PxKiiu+rmkUVuwvFc/zZLkYknI6WFQqsyaxp2PW2gkidKM1E5F
TWkDk8h2U65SiGfN+/dZQK+dJGQ/soxVEGe/Yq20XMFJEeGG7NAlVhpjrnNqxwYJ
kwfy5rkOnDKNardPfwhzRXBlLWzHw+p+mLGbJ8GE90EBx6vfpdN40kVNweZ3iKyr
MAvS4gyKo2mpaFuOy5OUnBsSZ8qaVib0amxElArFcQ4c4p/anI1E7ThHnL4c4dHU
TlqMeEBBlGk8olWrpuMlIVLpnYXz2vlk7hShsnSuVZ2O6hEWcz+I4UV082natEmw
oiCgE1+xN39zwYaXqONQhtM1KwScVjq9kaBqCqcp6+Vky3pJfAHkwamJj0SnPipE
2Tnz3ewtaL/JkUDz/+XJluYy/kRKkhM46BM3jgkm6/L+fK8kd2M3nxtnZkLlcSbX
Iv9kZZiP76N0nq/QPrAunANVWnTw5uldlGPeO0ekJKeTDrOrNQP7WT3WPBSodwdV
cNivZfL7XyzWzmvLI5EOppcgmJMztbh5gfUo6pm+Xakp/dszU1J7ujqG/m/h+AHz
3gCAuBojh0gWyU11ErNwU9xh4hWPUB5OE4uSkXmPbmYZDxjLQCxm67Ioc9tYzzV0
RaS+5QWZ9NLreXJhduXeNXcX3MekBlac1WDj7XJ98IB2Vlk+640QNamLvJeTC+RV
x46mpnUgtDC8Dhs6n64UUIKGgzRo8EOLtET7oFi5dM06bAZEelld/BK7Rf4gw07+
zDmb/UcqboKukSsJNkkDqnKAuwym4t+DJ4d6qYxrxnhv9tNDh0uQi+rQhOQbtpys
MnSSWMkxivWzQpzrQaHT0A04zJrzJ97hOPeDuPHsVt1R4r93L5vAr6D+RMeCMNCz
yRe6aT8i6y8WBdtX1h83+Q6W7v7rmhIDXvf1A6SqO1H4yn7rA5XUHQ2pNnAYs0Lz
KYrS67YL2yKEBhzOyt021Ue/Se3uFTJc0qwr2l5vnWtIZu5il38FjiFeChGnknDw
3d+sFuqb7aNKtzQtnrplmjZOshV0J/YNzvGcS5gNpwY=
`protect END_PROTECTED
