`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcY80lmNPFM8rh3fD4K8NMpQZHyM1fkOOHvMG0QlOpIlxIOlDPy6H8reJrXa1J4y
xgp6aQ1ou93utNEMrFffk/yg0BjXgXHdGtp5AenrG9gdoEEDMi1Lf6YrIO4IgHB4
7j0e8qobDnAth9V1WWT+Z/b4ySgQeOQGrErfLPeOi3/7SFDZsmwp7GzxAaxfFflJ
aPXSfh3Wb/03OYI8XQydHxcbFjyZMz711vUG+Am+LUXEmla4brL1eMir7aSKl6gd
9TEPfFWzPJyeg/Mqb4vvBcUz1vW8W+jisYmTTBrag4sLnTTj9oKnnK/OuADJDEcH
2AYcQGDIuJUaSDysqoSvTRfcqDpDomwfAdfdpBLG/16boBI1Te4FQDEzNshsGq5T
pWmwV1HAYXK+MRX0m3Y26VYLV8xoEilGnGZCA7Vsd/7u2L9Jdkfplac3vaCXV3yB
K84ixSXhTHaXTxBf93pfB0Y26TXVM5XHKTdmpANfDSVYpBZ+5MjhxMkYXPeB8olO
s2z3j86x2rrbW6GXOgkIF35uEr/uq1l9XJFyHiS+W2Ss2UtyqnnAFAhXj/yZanZ4
WeU3Se/ojAL2ZrbAvME5FGZ2ubBw9s8dYNo0/N/NruqPSRDj2uG1wdPunyfA6T8I
Y8ObzITLBkqaoAMS7SIsxN55qpIvmVC5gsJDkwPlTln5j0OLYha1B0CyezN7hjJJ
QI3HO5bKG4VWkPLGW++JnL0bmYKCoaYd9dvWdH9cE5c9AWSfg74w/LEAlhUdFYSP
DZx8SpyIaP6T3GH1DNkY7bpWmeabX4dQfCtCxMKpsXmZ/b/ssRNEXlmsOH0JKOCw
Hm/MAOdTMR+C4rOr8ckjiMW2c6r+5ffZXcCYZ6JvPkACxnnCWtA3xk1A0CrAHLnb
z4Ed4L+XmOfWmH/km8VzM0IrlBF063RQdpE/tldZt3+erXHY7kC5EFjAi0xlSc7Z
VRSAaiAojc6Be2H5mXpVqiF4KfJ+myd5nBxry1G6xT+NeNvD47iedsVp58Xu9I7N
`protect END_PROTECTED
