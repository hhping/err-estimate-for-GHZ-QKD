`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldYtAreqVCvDXry6+Eka6kFXnYTUjo1YowHKLaNXREtH/20qrirPNr6HaBKKwz/S
kkvr9s9KR5LeZr5aDSZcJ/Qz9LnyIm1JRiRMmaZ8hed995aismPoZOaG1f3UumLL
BJoN8I/QC6mutHvEjj3UkoHykN7lT80fGN0y5QynR045ry/8v2wa2vRJHcnK64iE
gEWvII0AHxlbFOd+Rj8Rjtl1S5/B7SCqnIkZN/f2KVrJ4OdDxDRcS+bBGokBJqff
WgiFCVqofV4d+nuMWY47VxcOEZbKU1FW2LXC3QCa0yuqjLXPANVyx2Qw9SR2BkXr
2IY4KRqKi22plEOG3bqcz77KBPNgbqUazzYUDrqJ6y0/4l/xdkoQoouTMcmSEOzF
kPoW1ww2viByiRa67cn7STHb0mYGbEfSYysTyRU/t31geXbGEYyo/ys0q4AemLnU
b5qqoDIOGTmqphh7pV2ZF439cqtVj0cQ0t30fYA1VvTiKLRNaiCpFYX+lveKh5/d
d7vsJELZ9SviDc+exjC8T+iCUO+KvFwF/yR53WZmQl/YBHn9kpocbXvh0mwRX6B0
U7UBnx2AiY3SRJDWHtrg7dAv9FyiXjg5fTzJvzG+aCEzN2fHKI4hBSFEMz9TjduW
+jeKmkdzFQ0EDav/4jKOyVHEnzXn0NmBqquSNraLtPJPNs+E/XmzJ+wE8DHLhiOb
NrO/V0uHvS+vzCyztfK7h26f4a8u7yKwfK+pkpweE9GZy7IztbRxc8B6SZ+8NPIx
000QIF48GpEz2PBLUTYbVZltzs9CRGASmIk4WaTBxi3CKVIlTivWhtqZKmrEH6/J
BP2In2AX5GVgzftpSpsgoHePYyCItQxQOUIm9WiG2lp1Hf8NqUins7MelghYqoag
bu4SZxuLFCIl9iwV5YENFt4q/lwWtZqs+aLTs0c8+FVBC9fheFyrVVcM25kD8zys
t+Y9J+u8fPdbglx/jt2pJw3TUPbk2ig5f1KzZrmOYhW0rwO2U63ErI5w8P+8+1Jj
AjaYHnDUu+1l+1zNw3JnsFYHZbhMcps3+5AlP7IOAsXgwqrNNw95S2ZezTSiURp2
Z2f9m0wUeDG+Jf0Wgu7Xojquuro5mSbHpPwW1J4lEnR8CK5PmGBBn4Zuxs5XZXBN
jF29R7yAUPlC0HBx/7uSkMBW6tbRAG72/9aKZce4eL0lVfNWJoNv2S0vMeo7e0n7
I1zycLJo8Jcs/81uqcqVJ6aUxtH+78DlTO0zv4GCPiq6lTBNnk3Jl2XDNaPBxAIE
Ovz0Gut5JzQ0ndDh/zc6tiQwmTHXRINHEJbqBRPbxov5nwjPwcHb3jRVaH4803Vd
WNRpf27Vxu8WuXVAbEXnlRuHdi11umhWBl5wPNgTYxmynKF7I+1RfCVyg14vG6SU
r+IuQ61E0YPYoO+T3c3ck1uisH/GQiQiSswp083C5cNgmlNVdctWuRte+corMZ0h
P237ZLlCQFRzzdJoTcsODTSR3E1B3VkFQalUfJ0gh/t/ZW46OX43ODoA4gAD+I1B
9ELRM3tgWJNzdf4n10MmNRPQ119vX9JQ+DvWdKsJGLtD+M8yZ38rAvu+06RsHRwf
JrJ3ifpkmX1ZmTH+1vV7SLuqr5wRfr5CdvWJeUmg5zBX9aVZrbpZcPgq0poyTGvA
d61QRsGNok27vFDF/IIA8lXIydydc5iqRxAL0KQgFG86sJf4Jqv5LCbHoZUgXYgb
RfesCQ/YVyMDPUZkKWHobbkicMmtKT9GNiBew6JTcqzhMCO22EtprNLDxrCbfNtv
8cGyak1Zb1YTZU1oLuXFm0lF1BxUVDpZUlMskHpt+VtDOEUZGT6iAQRUB2EVk2G+
k2zW8gq7+zhrpHgsQu7VRFwCHnhWfO6Kg7by1bW/XegNBoS23enX6kOqGDIJpmaZ
I5m1oBZU5epv20lqzdcK37atZA6rvLeDGLUmlsXW1ZTh8oRa8MKO2XB27RZzHSvP
RFp7bhqjHknELRsBgZOO6lcqOZKT1Xzd2yadMiBgfHK0zQ3Kd8nXM5OAN7+qRnCf
cA1/FvhzKWFcWsEdTu+ksfV85tt3PI5hmjnBCwWO306ybTY+yMb+Des1kSco4RrX
mf81ivZvbEviMcXbqXaxtmpZYL8p35lpyh6M/B/xGra6mZcjQB5gMWGmKW7Utz3Y
2HvFB0bmNGxpKUmk7aDl5s23Yr5Ectsi60Y7CxHZUL/hRjDzSDAGK1YkLCYu37kY
a78QUP4onf+64bt3py1PnTN5EEpuFRXEIPbuTJeRcSlnOUM4YtW4k+8WDnkgAc0Q
3LCWkszVJaIEwi/l6tOXi1mgDQRda4r6vc0O+UyQE0h4vwk86m+QxfChFW5uzHou
C1/9AMLZn9m42TIcf8tLI12HfnMAJmYT4GOHLbXLSiiWa83fx00+3eReM3GY4Jz9
SUThoYxLLJnX4skLmkuF5s8EooEKT3FkNC5b9/myqbc6y9SxhAMfL5IJe4sqd6fK
U8tgdwp/3FGBu9GX2+yg/ie6mT4TC3URniNvbO1XZ5Xo+e0wNuboWNIpxYCnhB6z
ukgz+k/wQIDyBl59d33AKSGARjMd7WG4eW21lRca1r0yWsc1du4/uawiRMiXH4CM
AWgGxSaMDdq9/wt8kX0PuUXKWmsqM93eJXkO603XztAiR1RIL0deG/7lJckWgWGg
aBVRD0hdKAykjvmedcVx7hI6Vgualt5pm+79rStrwDBtQSLUAAE0ZcPGAY4fQ+bU
myLHyNtaw6APcDv9Zi89oXGf7KWD3LLadfZLA3299iw+3Sx8y2bW5wgBHRCB5xdO
AqF6+1J+7icsDSy8rMDaG3nlMTFreQmVBGEzBY9i021W2uVdYAXLgBZugn6w9GXM
pNk5gioqndI1fGb6kKvKXzLW7Idu5nQxPNuf2biefecGD5nK4esMDDE1HwkPmazt
YPPbLW156ai1sa2f+oI8+hKzDxwSHBCCnCTKxQERj7CF70hkIUFi73rDa6MFRMDv
WVq8dWJjOh/b38+D7qN4+/ND2nX/1+K3DItWonHc95tIl8WshdlfASdg3PfqG9dX
C/NOuVJ2ejrXX+P5BK0l1clpHkJ8yKsGDf34iaBagLoIip2qvG+fKnwPWysxY9sZ
hpVPK9DO52LBNVI+LGebfkRazUXoF83522OUQvOzMjMZxL7uSgqBlmZMlep0M3Dg
/89UlgntYWMRJiOep8soNUDipG8vrswB8pige8bU85a3yywcWJf7gSV/CNKP8unB
Ag5fckkfR/e2ytcibDfcXQbn0zfjWNiK3hHb9POQZmbwQEbU3Ilv0/7XrRzo+6Ws
uZ04FcD8j6U/IYw/zPXxvZnx9Ukskok3hMfH18sQaI0JBMW5OcFbDh31KxUzBTcP
C7OvemwiwGzI69xTDoF37SCigAPjmLnxrqk6tC+QKc3ifXf9HAdDmOuGH2uCkvSy
4jRyZLnFsv4tE84E7fVI+x9ynTzGPaANi3NJVsdhybCIDSTGAlM3HFvif0oz77Pc
78uoTqKmPr00/T05qXbW1/WVHY6yYjeUWjb0Izv2a+n/tfewFKqr7zNM+TqL2YUH
xQPBYwSMCrGYGi8SV/vYekkEo+mkY9GxK3MnmPh6TIgJm/94wfsSXSr0jnpnzLmy
NtnNe/vVEADaEsN+tzwW1fLN1zVfKksqeGQOS9tQxYdELk+3sLCs6lO13jzYvqvx
31hJPdbgjik6QqNtPeiyLm7tKPvdvoXiMT/QGkU8vTofY5oUVrm+z6yquEGNehPQ
xr+zX1GHHdFZK5BzeIDNoAfsUjSPVeq/Ynhz/5Y0OKfsIg2lH4aKmR45wo2H7K+3
ZZwL6FvNS10e8tpz8Dhm70/6UMgqo3PuOk3hbjsEMTctbbXdLyqvVDJQZNNO2db4
pkmjwWhSBJsCdX6nSkLs2xwf7oFHkmNaHEVJN69DozWsJy4Fnm9zPopn9zz4uY4K
ab69OTsL7fJLD+ed6FhdCXpPUy3V/lKymgXqT8015Po5ER+JCWyOulLNl+7tud9H
cZBRMdY7Z93p9xS535+CK6ni3E1wnkNT6tBZN4YX5Hvq1KfVhoY4OP4GNHpUi/fI
+MDGlhKBa9tVWwAKQd+3x/FXHX0/bQgk/H09FlON5kUZmfs9pkqoaW1iBkkAvwBE
nY4/BEpDjWQGgytHSB8AdzNwZPZgUw0cxgqrOP6DbOFjsM8L4n7EM+7bWjfAO3Yi
WCcnG0NF+ncUWul1rzwylz6S+1U09g7MYQLG4OBndN4zPYTq1W+ae+/So/FCPGwM
qtpGzZ6ZSckYlbLKt8AmjDCXfEGZXAbyTXfq+Xrf/8N+cul40gPVUnzzjbwHjSkc
tKlJYeQuaDWPWLCmQy3F8li1KJdu4WEzU6Pue5XXh7+5GfSlbt2HPEkUBxOvo/tM
lfw9fb/aWYFM3I3fZ/xyaMsNJ9dL9bLXqjAqVJIp2Y6pv8ItMZXfmbwJf90qjP2s
/izyvggE1SsIwdAKqsRWG4qTcGoTU+tHf5PCPaIRRBr6Ke9rgCAabNCsznkBeywO
tq094MF2KrRyqsZUMdHwkBhjA4Q2/uzI8Hs+h+/IeC9GXnrD5xl22OmOQTCNx0aU
0FHBV/lJyGSVgJBZ9mWwE1foLvD53UHeKee7LIlSeLgiNTlhUmbzqn8C84NQQOYJ
VASvh0IeeBIMnQ+kgGrjVYTVNFTfTvaE1MJxuo/mVbsXoV6Da2rDWiVLJmIicBmD
VY2Qz5FMuU6wELae347sV2YHUym41dxfrdfawED6DjJmtQLqvNM1jdmnczZ/OcxN
afVhFe3ydDQZ5AB6LY6l3uKAlK8+QqsNaHVWLn5gOTGxDvF8CMq8wWifrGevLXvB
9PXKFDu2NDcawxFgCHciwEpCew0vUtTXkcoegvFTTpvo93mPc42MTYNjN0ObSajY
cch8vl2QlWdZ5z6fNG9dAJSP7wDpRb5tws8zSNoY7NnP0jgdsT7Ci1VK5N+dWAVO
dxunsls+a4iXTagP+1LFkUgBsBg/oI3++i1n6G3RuKHcRPWBQAKUB5eOWxhuF8Mo
NnXcr8K8vsE4UUfE3hvIpjhkE6hh3r88ZVMgVVCr5GC8bHYbJnuL6QqqFjfAUJXz
Bwf5wQQwDgheBE8u7eggMRAFJC9D+kZpx3PsDY/l6Tb91nUCCSfL+gN034YH/R2t
OcvWC1kP20WHhdB4mZRxAACdAQGti+uINm2mhuRB9WKIaZS5z7RwX78fbcopoHUM
I2+CmxZGfrRQOjTS+NTri4E6p+MxOIDNCZuLc2g51bNTQRZ+/+MAZnTpPDIg8z3f
9XlEjxHrLW9swspvC2AQxT4IeqVcB5fMq6nYGdOm4dPjD+bbyWjdnGztxBHo4XOI
lveBGgj1mf2DAOIrWPkY/OBZ57WocJTzb1Z+nyBqTrqPvubk53HCxx8T+m0+IymN
mW0DvvIGYBOuC1+QZS5WX5R2WjvKZwFn7Ny9z4b4L0PscH4rfCFWFTEnPiZhxZ7k
DycRU7+5A0w5987Ucmvc/H2ZFz6jCgdL9W9l/OEBntiNHDYESYAdM6QVFzqTQqlG
T+O4O1HD+7oIqSE/aPGWZGSlavkXGGdq5CoVqcdp1w2cXxPIfWh2GlT33iHlUkLq
2VOz7+uETKOd+GVaIhhzmbHt/TzD692XNrvkncUQjPLaBqJIxxAVdelj3viCBe5L
oObzt/lFwjfyvpza5CE1ylgAqYv0btfpoHWNqDtnXaAJDQthH6GozhOqeTie2EVr
RY5aX/5pNxj1sHiJTTOVhDW8pQ4r10u7FRibwTwQOnW556rDYR/3wD+fUnVpEajm
Sx+5bc6x++EchsS/im7iZiCFzBYzZ6/5VzuTE59LSspDHbl/9AtDTc5uc9+9MQr+
lcUwwwPI1VoZh8H2ZnmjFyBYbXswy832YGwAp5dhU0+DUwfiaOsmsBJFN2G/a2n/
vOAmKyyNG8ZUMGsymIWSxOMPq24wVabLOx5hcwjUYhxxljSNr7/s5Ts3tOqQKFjG
996pcUFUhOjj15I31o98+7YKYgbAz3dVyPGrqqHTUGzFYVYXTd7oNSvG5GMJFFBS
8XOYzQ607HnpIGPud7sDdwLqhpBDT3mefwqHPn9UozP1cRArWsCFw2kUR6O5Pgp+
03cHWb6isysuTzTPOBe6X7/HZH4HvAncb45fD+f5I7YZgANSTnn1rP4tMJzsQ74H
G4SRxL+AcEBaIDlGvB5IN7FFhI7b/AKTe8WF+djO6NZIegQIj5CAlgIvd+wiqqjG
P+h7qRUrqg1DARJiENMEOAnKeQrGYh1oj4Y5rzDx3+DengIaLes0OUpiYZ9lh70D
XRakU3xivQUlygS4C3KB/Vrer90Jj2Apltid+/OI+tvG7Okq6AkxFm7kDBCqG4Ll
+ML+/Eq0/UMXL7s9ux3d+WrMPWB+FLR3yEqnGkQ3UC4833h5nw9GeNS/80llGRU2
yXhC9JfIYqR103u8hECz1OfH4bnOaAJilmFUTTMmb0DrUeBWu7uvPWQRxPgaD2yX
aYMkWfASNlQ3nSlJE3xNsxurEd5at/RyGpYg46QdkMsp3d2fTpsTU1mXiQ0GqjMj
PSqdKf+7dU3pyacZrO2rum2v/nx/aKmlJZmV+mYE0enqJOf8OlkcY0/DAw8GD5lq
jZ3c+Npp/l6NsDb6RlR5KThAO7iHh1mw/70BFu+4GaZNKvTllImLLNhEiK0gqxA8
+kFSLLgKJOPbpca2LYI29/r4qX3U23xTrPb3UqW+/0RRgjI+KX7IeDWovXDUrXde
tlZPIOG+v+4fwiwzm5YBFZYlk0Hd8ZuD3EZgACt9FIGgemdHFKzNbNmofSRqx3F1
4+CgD6sU4Dw0XjqGey4By8xGt/Ey8MKgTcg4ZEI9hzy0pYdE5iQH+QYUCZy21fas
3aQ9kT4e2jdG1irjZftuf6KwAQoM0r1QfcQI49FS9U57H15sTv/11Quo32bAhj7c
PuN55E8z11AyqRebjT+AOubwmQYsjwTRJN/4igsMYHRntsRk3JMKQ8rTGKl6p2Ln
qN2ZgkB4cIbamT4w7dzYLBzEmQfWyl+qBwiXdYSjxiDDjCeADJZkUVSLzW5o6X7J
tnibiXlgBBuvLn/hA8yuHr4EM769sFuiJfMThyQ4/DiEfL5YFUSliww3JFAfLQtP
HWQPPbxd0OvUJUp2t1jBeFTubXF0jlDBeuKmmV+bXX6jRtUDnQj6sdUy9JCXu9Dg
ui/JZXAchCA4dfIRVFMRFrKdNFF5i99VECWbNlTNeNucWeSJzTji3KmtH9Wp2Kl8
jW37LhQGAzwjJiS5XM/0wndIH/4vOadUufDooMEC/PjkCK1VH86EHbkpA1I+b1xS
qluJ7PbsAJV+0Gj098F0wL/VW37CV3NvZF3lsKUdrxOtHuPNROw3ALw9TEBuK0LL
lxRj9VBWUGVlx8IWhD7sbpJ0T6nIJ/ft7dOqZ3Ehf0k/JP2exI/LsVHmN4Bd4I2M
G0Ezuo0Ga/FNQ9m9Fw94on63SR/s1lh3UIHp5J9kcJhRBz0Sn47yFnQkvZMOIycP
W6kgsKgYBbgkFOFNr7OG/lAA+LQ00usXBkQabVZK6HUm7sDjpsL+CgGHa+IxnDue
G/ZcBLMhQpBcAWSiFpXqViet98u8VYCY3BluHDpcSVh2eJcwJpSwJnhb/no0gdSR
JkmW16m45FjhJvIJxortlLAfFUXj7skFXzvjPynsYyMQcar8HYj62ssgHNxrxu+H
GTq1p7FyjxatMzakUA0b7bjE8GObjb47d2ZoAV5baKT3T4T8PROvphvXs2bGowIC
nVHvsG8vnoypl6lfdaG48IxSkjk80kFsbyYQMtce+9pTCEMIRo1dQ7a8ynGNsWny
Qsh0oUOHdu9kOPhD92eUNxZvu0Gte3J3i/LskClkCRrEyS3eucr9Wub/Fjnvh3k4
d59MIFpyHqCiApzp1LauIRQ77LRo5DHpcVbCxJBV20RFvvOVyhqcVlHq3aSB1WGM
lCIefyDsJ66L+0c8lBZMzU/rdNWjnbtZPv2qnXXuzDbtFcobBqHAD5Lz3qROzPk9
pdJuziq4II6/SOINqB5Hn+8AtWkXcgny/UjdKJ17DaNivk57Z1ol/aH0O0Inbmac
91ZDE/OItWuIr1/eSKyid05hOkw2xOdK+kv6ss2ATUZwvSy2CD0zwhFwmB1BTyI6
j645T98om/+PoWRKJNa+bJ8b2io9gvfPFjAVsJbQfPU+6husAdaNNyvlJpmboA0K
f4X9nm1hizjrI9Q0MZknJoh6mzXCa86kTSNiVwJYCDTLN0RJm7ZaXV38E+pxC6b6
94wckmg1EPDHV+eNMQ0q1VuwfT+Q1JxjfRcT+3CrivYxju+huHKtZQOALGl+JNYd
6hZw9gEIXLi5h5pVGG8txMHRzMZBThxMc5wcU7TaccXilH2cagHrf/O7L8haM4eZ
4zAhB54sjsmzIUXPdn+g59ISQpoViFA0GxnuSw1aTSAGwCELsUZX6IThgiXce0FF
YH2kinEMxA1E7quQ34u+nFkw8KndVkoTbIr9/uTuKkNdIP0xJZ4pXPzjgxQ4Ma8J
6Qs7arrFKvHi6pfU4LjKn9rcpv2IYRUB6WRrl19cAJqVfUvArRw5dB7yHEK6VyIZ
3yJX+5IBXU3HuKQv1nnciJoHREKGMYgW8oHDJvzKs+kvuHcVOJEXOIcXHwTDAmzR
96M2s1Dv1oN2poIcQTnXPON0pKxpVOrmyzJzVVFKFRyEaaYV/M9pNKklwia+luGw
3Z53pMf82zOUFjAUgjzZ8LciqR6R3be+YG/WY6jqwuTKlRFh7s0kYrxTt6eods74
smoCR7wyG/++S1jOE3zIUH4mBFkxirKAmOUh4QQRaZhqkgiu8ePZgOXvk1Hj4MLz
bClphi0CmciRkK+RtEd+DG7ZHFPToI/prnY6vbu9yj3VJHRSGMHYBhM6EDFryN/a
p9hqY9uZAlYNM8XAH7kjEiG8dWQrRNp2mt1aWXb6dpEbopbTPABcCU8D9JtJPob4
ymiKA/HIG+GS4AJnl2VG998fWa24kwbt/MpToIsNeT74uvur/yoOBKHmPlsNU3/W
Gc05C0u8KU+8lJGaM8asR0MSfvB4nKkZVYH2Bt1rt7dvDLZZoYjAf6W35Loc/33j
DiYj4208QOO098lSul0j6u44AcI8fVgl4qZdMymlKMhOIc5ot1PCBTP4pjRzowqO
JCIixJGeKd0Dr4r7rwqN0ghm6neFd62/wnjKe1CE2IQbBf+3z90tcnkPk6AZhe4o
6riHAOVPsz0v3g48bf4Fk5nvDwYTE6ZrNRNGC3d1O/igIop3ovokQi/kOw45I2ar
aAOCV1MnjBWLyEOQpNxHzUdTUnrXLuBJXTKxI98r+GFnI1Wfjp/khY2+uweL88IG
bbOnvDCNSroaSVHCllMfSLLF8TFxW5Ig0MVoDrxq7M+GQIPdeyGOnD5I2mQYCzkJ
VmksoY4jr4oI9iSoepvo7VL+c26vy7YXLB0Eae1xjc7V4nIZx0AvSXyyWuB4Jv2j
qplKuHRICx+rJLBWnZmE8GzxE+H9+ZixmxOG8JAo9gZZunTqCWYSh1ByTDkxVnmu
S/HVfZ73LLvGpq/oWP8R69hVn8he2wnHvpO8ZwQD9aBWAn51F/9VDMMWDq5bUHDN
uXialiCrEHwMiJL6n2qlUsSkWmJ+FE6lZb48fDmlyA0GzoPKAhEntOXHBJ2ZCyw2
1e3EXM5Q78z1JfUmjtOVa7NwJEtN/sp1AUXm9/YebgjFEl9MWE2MH9thmLiLblaW
2X4zKmczUFMAi1ZtI8nMZgAKs/ITpO9zx6rsn9iP5VWlmXAnvm5rtZJMP+lIr++E
ROW4ZW7VhxlWQJ4PT67Zw6RTcQscHpUJetbyDkT+FgdBYdfRONsp+GuOA5BxXVh9
fw7AIcb46LDZxUTcmhNxc8xIcq3WdiVzD+0OzK4ssK75iXTOp6+ocpcQAc/5aOk8
4MDup9ktpo0BbIsVjeGZKpwic0UGtXzdqJEAbyJyA5cc+CRioDDoCsbJ725MA/IW
HJmXZc9v2h0/rSmGwSZzudfqasHQkuD1oxwaa7/tjTx0R3RhuhluiBx4+0rFhE0b
4XA3/wQaE7WrVp9rmYOerJuXka4kABmgDddGJn75OELdAin9pBrT/AArrAOeR75Y
Ush3jr60AFccus0KjshfPDMrlaMfUypJE0nsASESc2Pjaq+Rl1Kad6SrIY3KX0w5
bFA+wAV0WrfXIdCEEKeVXhnGSPdWvhLvdkTUwpib4UtwrHMLDkab+HsY09vbzgIx
cY1e1+KWQ7hohvvMx0B8wSNkvypmUAaMsgpbkT9RfGAzq5jIi7RFQZtEG5rje8KX
c9GIb5spX8BQce+PKzRanqHwYd5S5LNb66PGY/NK9PN6crf5hc2dxsHJ9IIMf9DK
S6eMPpH9hvTCk4DMLKjGFKR+2oBuMmYfPHgiLS7qgkBIQY4c0jVk/WDAONp41xzd
jTqg8uINR5i/pgvNwEwAeaNXoQef7KVv0YygkZYgwK1WcmncUE5QJt/khLSnHaxy
O5w5hVuTayQq7dlWD2CpWIgqGa2dCGHOMw9S2mgQb3u/RbZWhdIYOaN3zhyIQcYk
L1XB13ZOd3BQHglbnmHKXrP4Xq4p9/CkdMegzvDy8/LSKzCiwcgUfwOJWbw+m1Nv
7UGcDrQHHEqxvux5RLA5r16eYkjlB20TdpCbXwDjctGKV2JPFYAEQvQS81f2QsZ3
JGndpT9Hn9XnML6Q5XgixTi/PL6YIEFUFOdnTp/EaXYN+0zZHUHOX31fgLbtUD4h
xMlpg9JjDfqQmGfOWzwDMyowPcfQOBaXtCAWNhGXoGrnHpDqGvgkfdQRpWkbQ7OJ
916mSS3w9rmJA+BK8uIWGSNp1vYdAN/3z8e1wyI9EUkJruumEd01IBCEPFK3G/ww
uSGSrrtD7fj2D4BlRMJvDP1gvFHxdaKdh5/RPzOhyoDhNrU5sXsUhkSMg+JaDysU
9E5xmLUn4rdKI68utS9vBfVqNr+0gJaM2rF574M9PW7CokFxYr9xuXYMlw9qYG39
HIxokp0vh9FnjDiXIhEmlvYb4hahWO7tA0F7T4JboaouDLecp1lnDQfbFnztMlSa
VlyUmIVPOW8HDZI+quo5+jJe7pKyVy4Y1GIUrKNXXAz9XbC2LaFf35aNB5nMtbP6
WT+dKe4WIMSq5tffvEFLcjusJ9wsGylWKwar1mBfIx94AoQL2urifCWV4JETE4SO
IlqeDtUk7DlNtJ8LzdG07rHccP4CilLZJcx8N5iDgTQx/ZVpfrW8WrDAQd08MW7A
D8GGqsEZ6riDYJWgXDMKVjlfFpxDu6/TI5yiDGD+IAE1SKHV0s+5aXITMzBtjmX6
YdpRbrwEdphghe4NAfUpWLVpqVZ3TAIP2S4OjwnZ2Kcwnq+Zv42eZqmnNv13oNAG
mbD7pw4i0Z5gNfP/dEvSyzoGplvy/jqn7F0fp5ODSNQCMBSfhzvbAKRY9H1fKRcp
XkvvyY+WFV9PJcdj4sj0il8vZdTvsZDk0RbhfYbF2DkfNZJ3E/2KglUrkP9s6Na6
NP4o1h1zw/nHcc/vFwSBzwL7U5My7niC6nvo76Y3UiouXx38TG4YDoYzw38fH5/U
1gn2eHvQRrl90rzSUHrrfI6Dm15DOARmJ/JEBo52ZUzHUMjdTGHGsfnx+I+cXC0C
VLtWFd0XFsMK/2zukUTcBiQseFUEBGXak/aBAlNIIC744f/tx1B3Wmy0BydtXR/5
01YUHIcpnHHGfo5iOwwmLzl0Vk//RA5uZgTCoHqJ4NcUYKi+MwLThkAiNpLaYDfG
4f8QwH8FmipEeCfRYM98fVAwLP8Vi4276vBRcLO2CrHlvoe7BG9UxwEPONb2pHlO
6urSEv4+8uwGWUvHL2UpP3JC5lsYTPKnhOESqCDtT1IYpvlSdsxv6MBBKUPAOnKo
9J/qbT02+RAlt7dGFu7ZgBghSongim/QwEmks2PvhyZDgmhLESuTH01tGWKd1sAj
fkSKIoNhvNG3yRGXUtO0/8aAajWXDUCQWxjJPfhGm3KRj68noaDywhKUHt+v7S+w
Kc6me7gXyrkHZSxkMIeydmt1joqbbFQ7sCpdPttse/kW2CXU8uVe+6XLGiQjdQfV
5yzUrn/YDXfsS6lBH4ogF8pnVBXdmPGB9SPGerF/ulL7C0NNr0elgM4TolJWs/uG
Q2l2xmf29h6zybRXkXuCB/RODdRiLELCfBfDjI96CaZ9cxKWTMWrLyeu+tdWo1Kq
cAUt2b/XvofwZi+JEt8QLzV4CiyHu1nBOkQR5wXB8aMoMbYzSzoMNua2FItfSaSz
hSI3J6n6OoGuWslvTf8mDb3X6KXCs5Ber6avHMVYwsuRBiqKivi4n0L0GhHAAvZ/
pu2ep81/PHh2ky33f9BBgVGKL9AmFqsre2V3maqvt3EyfHjeKehiQjS3Dv5IS/cN
yAhIej/BF3Y9M3EfltBQkMCOHfhvjjndGh8A167lxa2W3eV4HbJjER2qDHmjTR7B
YFHtdFAkvnXFFbITLHiiQ9aBGqRkNcIyZPTux20bJ0DaK13IDjy9QDIGrLG0SbqL
t3VdoUipBK9eeKPWfEGWtSSlVdRRA185P7OPqciNi59h0kQryRat1Ph+4Y0+1XRF
5jitucj9s1KnQ41uqM54rN8RgbchxZMa0l83G+vfnZRB0Z6pS5liWocV75zpKl9b
iS/BsH/o+FaqH3ybocgin05VfWp6Me1pwsrN/tKIe4nYeg7P5UcR+cWDrirqyo9y
0d1LlufqFUVhpPUNc6fYJAHJuw5ZiUwLHy9P+LJ7MgFfwxs4QsuWYk7lvSryX/ZQ
TVYa7/X7SI4PxRFQwkczlZ76oFU0DY1F0qvJ8NfwgARlHI85xmLBRy8DVe0+AP5H
bXaWnIXj38XWs09zjqy6dDSbv0fMgIxuUUJyMJW2GuT8vQmB5AewqkPBGcKaVFWu
F+R19nCShiy/BmHsA8dw6q+8YrXlcSFYHMvPNrocOhRzyJGakNGGS8vKkhF6BknX
LHLLxr4msHcx1FTt4ZthfkFay7R/py6XL/vWfAaXYoZCCvjsKET1u2kWyIjatw/x
pg3eGXn1I4glFQLQM+bzjJoAbVJFMUKLr9HP1vnjyr9o14aq5vBCCPuJo3v5UGR0
ig0sEF2PRTc5NeF0Xxa1yrHthZh4nPcZNECbEKh+lQtN2/G5TCgvKDFukxcf0NpL
3Up+YAN/qLlLUlplxSBpA9xMLOLOcQ2c8ckNXzjHDNI+1N8eSpcA/T+sU8LMwQal
K0B+D3Gqua7agXRtfJK0gtx6W/w7FfHqPm4XDYPbkkp6Llr0BUQeZyxETcewW3OE
GtSJecYi6mbbm03L+kQtvqybqphsl7gyCuGJVTL5TozXGf5PYb+uDVXpREqokie6
1vghIBxSwU9MLlDvqT2KIzcW1IlCXPTrE49URgd3kU1AAE4Fdp+W4uSHvQtssMjQ
iY7lvvoukcqIiAxH4Siz12E/bepy9WQzn1wCKm9O2He6VoMoGQGsd1guD86lg4u3
/WaZuzFJMcW40+6MJuCSVMp4cxkJtpET0sOrFW5tFeCw1qDye+t12qUGfAQm/a7w
AIZc8ZWwumTiiYekYCIs2G9vcEDV6v2ZiD1sdf1AP+A9xxozQox54yFrF0uYCnMo
PVi395CENcmdaqE8bM08y3QUK627sr7FYTdt2rl+CYQXprNU5DzuQpyqmdN0NCan
+MH9lnONPfOxIXxdXxAOqDD1XV14sHn+5Im1fy3pGoowBb0vKsMhhlpru+BAp7KB
Wjtk5f83BYTFgGo5gRrTQOcNuH6a7Hap/pv+ocPWvcZe0N0+WVx+9opwzE+75OcP
wlJNJsZ9DL5soDCgVsQnRkB+YmkoOPrHMgsshidINZb4QFUVRqqR8xi9PjlKUlE1
5mVb63u/UmallUhTMM5QjweJIWqY5xrQRqnGZ/yPqvNBWsUfZcX8c2C1TmiOXVBK
P8B7ONhF3F69qsJAeJ11ub34LSSLssGQugrIof3Y+TXLzJlu54lWQwFKpfqOZn0W
QqqGsxYx7/0UgTF8s0Wq0lwoTdvtko0Z8j9s0K+lMKthxx4qdKXi2lniBptY7U8q
ouKFexi1fOJ9ZOh/7LPqkLp/JZLTA4J9b4WSZ39C2/FaT6tARk/x+93yjH823zo9
ntaV7YteEaje3mH3a/efXFLfd0aA0W4ZOmXsghdf47u7apRgFc1/Uqb5YjRvAajn
9XlgNQ5Xrq5EJOkr12aA0R9RxLpZylMI0hbHbDDORVCOl/B3hxc3e9C33xbjPKbb
qzRL/5r/p/SDQVl1Vc7ByyfZWCOXSSLaAg3W1XLOKo936sF4Nd15oZS37jax8drb
JImCynBhwb0ZElsBF9x+TZfkZIksreTGxMf5bLOVaOAXyuIu21WghSd5RFaauwGF
TUDX1J3CL6/GXYZA8RhaaZ3HIXVz2g1u7WVsglUxAcyNRpips38w+6eXb1LOsKF8
t8GlJUuKTOHdlK9cL8jOLWCi3wDGhDk3xqO8LeoCfO3VLgs7ojNYGQo6r9Yda5pr
Wp6hujHs+5JQ60yF3hclCGFXJUXudhD60BVrcwfQw8akB2NgQJfgjjzpjI1O4GGo
dVVJe2TucmBcfBnU+BrQjhPXRMiD/ig2IzDJhYH9IFKl8+VjtmcB0P9Hwd7hMQ1u
u4Oxx7vIWSlyGHJFZ2A2cSyqW2E82XVmolATcR5BXjJIs24qczT+fit7yuP4n4bt
kBho0w0v0GI4ZTwkedhC2CjnmI9sPkTFbYmjmWqbXWwLVdgehBQnJNdlsW6JBtVI
xW3wSx7H8SH8YhxewSBeh4oYWqsoE9xnHTl1KVPvQlIVDZ93N74ZyhFsNhr+o3Kr
Wi7ghunH4xpehL6u4WxmDvcIuySPvNX09B5O0RmdTTPfkk+EETQemg+2ZCxFFKk+
Mm67xXLeC8eL6WtfxO+2Y4pVp6K8gmVQZIfomHvnGsPq9oNk7MKvvEqf0jx6W/3K
452WwVOrCbEhUvKuR+Go9CmOVaN7ud60bFAE7M2DY0TZlsgsCNGmfHQi14ozY+11
3KQxVE3dJAsIKUgpfdicWK4RuvM0G93le6XinBY5sFmoznksmsH7lmVJ/gmtDqRY
uAauv6YNgkLJsc/0QwRpKF8PFtZoDvPqK6kh3CWrZepihvWFhlgNsfPO8bPDvYPK
Uq7Q/cd01WIWCvuAsQMC201Yv4Y31BuxtSQK52M3fv0sfIspUBYRGGoGxvcRL087
CehFLCnzokp250VnUx0qCoNrxUId/Vioc8jgJxWB2VOc7KakQtFBrPypOCVuMv+V
bQz6rZeYKkjllFntrYKPfOKv4dBvfHuweY6fplYR/0ArJIOW+VnbhZc0RjkEl9Qp
kqRDf5ecEzzVwqoz28CPurdvlDNdKovuSLuyq9FwZCKtgd5dZbnaKAEuzdzBlLZ/
PyNhvtt8TIHx5bCAs0bm/pHz0zFWOAhOYW0hPGPnzkDzKsT4/l60Mem/6YT4Kg2H
Tv2Xw+P5rIWmzOgeBBFoFPhp7OZyPr90FoIUH0C1LANTSiWdcxhLbF9dhmTr1Zzb
L+89ZHDs3CVMmof63HPnZ2my7bR+tTjjYn9Tl455R+wIqtO9ivssXEUI1iJQiFif
9wPYnVtNcPNcUGBW4v7Jy+SHziZfqHn2r6t/Yg92pnOVfAn0OEE9paGFJTw68JVJ
kqaTu8L+/bWmdzh0TVoPq6UJBiMlZVT/4wn60sHovRne/k1dMXM/JNUzpbpinqeH
NRKLsW5sFJmyARV2XKhTxLfc17VLIR+1jF6TH4LF4aXPE8sVlcTQDCRY2g22ADNg
uus+CuSEw4laRQQuCDEYhcU4FrEfkc4d0M+p6eOdqueDG9QS22uFIQwp4ZWQw+Jl
PJk8kzGPaouZjwStD/lxqbsROqqHrtIOvFVWbsK0KvdcKyhaV0GbyweZie1ymOQY
v+ZseRD87iwUWKUtsu1xNdwChPpCVDfye2ijTXGBh+g0+peTSAb9KzSKBbX8yka3
c4arNDGwETuh4MLDgP22+D5bSF8YH2Xi3Z4UD8wcQhEBWiJavim94YBMWT1mofif
P8rvNtDc/92r3bh9fPUKnehaIKTOV6ohILs4bapR5fJFNKBlq8EKo/a3Q24Yjja3
TvqndnzOEYcok07/4SyhBy/ry44nKaMz5uhU1kjV41sbe7lJxgLnG3o/N+tszrqI
2LZLMJkMEnX4DBsmiV87SOGMwaObMirjgm6PLujy8tdrP7vgI1S4hDXfjwW16AB9
gG3w0Vjip7gk0mORaJHobXoC4qBhYG00464t5Hw4GinyDufEcOiZikxUzH/wh7WV
7VIvWT/RWZc3TUxvxX/pAouUPLlwPvW8ORxj0w820Ieng/HHhtfBl1j90wf5z7Kw
7gLp7o27eLo7ZD7IbRlarK06FL41EeoYyvjSeIEtNJT+zNc7R4wOhu8VY6fssj3W
Vy5jFpBdR/OHTY+yKK8vUVrFu8M6pZ7GnToeSj2zUvlQn2Y8SvOcLgugHEAvJDy/
KMEysTgsZH4wWcWnT+Gr7styWB+BAXCUeOlKqNs5camKNQDsZaVtI1O5+2D/Jgbo
+zM7Sy4X4rbao31wnPOPEAReSbbIeygV5kKtHhjXMZbnA9RfeD+9Y+v4mXTBkhY4
5zoCUz8ZJ+xw4vk85hiAUBoecuWlvbk39JAY3AosZ4Zj9Xbqhfo0CDgyU7KYkNqL
MtLVt0N+Fgh4f8G6S2rB5lgfb1s1MdJkqE/AeEj5bhthqe6aLNl+1U2Lh/fORBb4
Hes56frQTzg7YSe4BhMwNRYQN+9XmR44kXq/3Nru7GovWPC/XlEZcxA+19lenJO0
KGgjs7yfcpv71cumRaumA51zNuYLkuoNUd/2eaMtHg+LzKtXJ/3EHU+y/3JKzrmF
sb2XpleUzojL/m+javfv6F88k4raohAUHl3f5AfyK+qG3k0Ee1+oV7bPtuqHjP1L
r5AgEgem/3Qi1ch24Yp8Xb49HcbP3mC8gLDoeptZiSP7CCNFBBIKbiapC4PmrxqM
OFmHYDr5/UIgzpv6AWF+NlUYmnfuIYwyO540+Suz2t+X19FeJ+QiG1q50nfUQcvH
on672YIVoEPaMqu7+BWofav9Eh7ErotD5vcoFGmcMjWCST8V6w+b90MHimglljua
8nHNzL0z/jWMqLoY04HKfJixPuL8LgmPXQHYVIEcwXZKK5wnyFP+B7nGwvKxDZ8f
X6FxciSi2QFVUjl5+rmPCs+6FnTN8e1to5OlXEgqwq0XNRY3gWXUHmQZFQSY+gyR
50oa1QETBrC3pIc5lS+N+7CFXwzCoj7cfyGHUBeQXWax4rYNbbohr02n5UmD0dQZ
4urP+H843jatEEDKHVYZBDRx5OndtJwnVBFwj+Mrfgdw0T9APIa09JayeWgV36WV
t4VL8BmxKiGi0hGUWn9Ec0Pm8n3Q+16/rIDcuZGJW3AwJwxw25031JIrxWi3bbh/
6wJdJQEE+ebm5FKWE0HNdrPm6a4eCH0GLkw5Yl9FRpjwAPa4u2s+afiRUXpnyHn9
nCfQmvcEm/MjyFVgaeMGWSjypwBJzwSIjdi+pzJdNQHPQhf6yElqxchUtgNM/MlX
uUY3PTYJn6LRS/RbGX3uWv2OreTfv4bAiIp7qO2dX2Ds5+04Vs7TVzbJ//lVftfs
bGoLM905NOD7QWNlEC8zUwWdO3fGgWO9ex7vBiOKBlJB3YLS3mSy2nzRFJ0AGDpy
WpQmY4SXp1C3SbUo2fSj3wcscTRBn6pFZ3ybfusS49LFCYsKrabBg8rh09woS3pj
dcdcsgjVXUy5UKF0ZwOeqH+LOC/3COXElWiW9LpYu+KgaahE5E1ZKO9FcOwxAeUP
zcoMGkJBmBo5FbZyqxpqe8GCj0pS6NXzmB43fOSlzB7ZhpVJ8rZ9qMvQ3a/pMzZz
qOTZMpR+vA84vvuB7UqMjVNbXKDK43OMOumUIY9XeUy/q0ZRQ28u+ygXHpF14bvB
pXUqqpGaCt3/95EFCbhnaXOZJA3XZy/aRxHGtAVwlyiOnnWK2p2Xf5XLvYIGIVpw
5PhC2B+X8jwVZqUlv5oYlOolzaVhSbd5NAWuHAqM9DsozX4WXYLGSxmb072MU3Eg
bzqZ0Uqw1KtYaFLc1yb984v8KKpmWQIjdadffvycVNPkZQ00Hqgv9ORvQKSAJSBc
VOSI2F8bV31TTuTnUu28dw4blo0G6ZhMueBFo8hY0iBWeUQYpPrPtjarf2mYTM5+
Ul9vdxme8Ua++xBGBVvtIDqgkJD9sAKsED+bFxYuOEJhwuDhMpKRmEqoKiuM1WRz
ny3Q5JLJjSZ1o8m5i0ub3D1j3l48c+ALPTRU9bDrFqcf+GHpoEw2mJMLM9OzgxaL
9Wd9nivTFnyWP7vGE4h8wcaYD2eoDobEXNxbyhL01IYOSVrMZOmhUK4CKkts35O7
TG6BzOBVLUNtdgn9voO0DmGAhGNvAA93b2M3MeJln/656vkkNkyFTVExhZZY9AqR
ti717NsU7xrqxk90bWE5zQt6f6W5nXjCL5kURcpfA9mZ7Bqnsr4iv433C4JQ8oE5
kNyDkYoyHpiMf9uvfIK043gAYyIbAdfD25I6bOsR8wmgFFCjfDV8Rqx+NObrv0U8
5DnEoRhAhLAD1WjY7TCGwHWBM7Xt+sRh8zyjSS0GvPZZ2o8CaAWfR1K7hSfNHbES
1Plhmfw97eUTgBHk1GiBH8Om534nm3JtgyGykZt92gt8vDcOniiSvYpeUpWHaM5F
ZTz/+l6HobLn+FD6SSZStq4clHeCKvmgzl3TA0le16H4Oim9PUPZ38kA4o9Yuap+
HFQycZpi/PAYywK0amO7a68gpWVC/oSshaNUJRtBOF3NyE8w4/TUmkNuNZ3fibh0
z671FokvffWSuSO/FpU3jjcsq1Udfd7z8KbraUtmGj8t4nGMKP6fb1lkjlDaB1Gl
OOdTjnzR+S7MNob10s618jZLeNsySK9DGHEmv1Y3oUDOq2C/nYc3X4nyFa9hedzC
Ah36fqTl/fUXaeRlKgAQD1W6ABAfeFXBzJYAFxwTYxehD4cEE+qPHxXcRG6RQOeh
aDCD7GbWXIPjRQgC2Bog4xAYTK7ssf4RbJybXTz+awEyAnm+Dy8NqfwHbUk9rEsP
d51CqoSsGj/Fxy2crkjlDylsG/qCG7ZazBaGj4PJ9ZcrWTEZGC4VpSFDyopx7ow3
Vmbu9LiSoUDQCzcI88JtrxSMeIF0jZ2y1TDf7AYDmzwHAUs4GamosQSxn0S6YPji
H44itC02mRlYf/VLUg8tDqDGHZjw0JWAxpXmHO7RE4iqNx/BoXlkS5D2Trcr9pjr
UuQGmSFJH5BfAvPJ19zotKdmZIoAsDSHTiiobd+dT6Oqu3LtsokHSH3cUy9SsUTc
R/rk8Co30ddHfVPOucXD5jBN0UIiKqwxqSuagAUXL3FcTghibMThfwFcSpdE2y6Z
C0t4y0qFZmeSi1veUmuxegF8pM4zjGaT6Jip2hISNglYKwImmDYoVYGOlBpy4KbH
R/gaoojYVMgkdG62WJzclP7O+Y5TxaP7C0/Khwq80mu/g93TFvQsrz8MJLW5Hk8e
vGw/AV2N9QYTOqMPUDt+Y07aajn0Z15z8cTEr5BKriHPqSNcQW2YnDZlD0o7Sa2X
6YVrVFlqfZu2Gqarp/k/O0Y6ObwMMNzzAWy7IjZnn7Jj0qJ6RLXWQOoDT8F8fXSd
Srv/xmIPlSf/p6xKgkQOfaPRWCjjhE0BiTpZ92Pow52wQsgpZywVO8Zc2swQFc+w
jxL+Yb06NHjPHdkbJAbW5ElLNIrf0mHyA7Shc7jRVT6HAAZXDkcAqbVLBcPpfdYg
nUNrGHr2QFQH6QBUtFXoeT7o1/0eJUgFhnTZ7tXjMznG0cm1z3+xWTpVFFCWVbq1
gp32wTxAEgAFruy6E0NwwoWi33baUCcFbFPK1wlW6wXvOo3Eojfm1+AosrMirpfV
ixjQxZTzuJDGpEri3411Celcrd7TyEtwhqctGYkmnU3t3NYBsMNVgnGgumqj76NM
nTIPjUbBL9dLfFUV+xSTlmfxknnoH7x9evsFgqjcci0QivwU4tq8j2zU1BwLqPyL
kXkeFRaEFLAqqGX7ADiU28XL8M77F8O+svL4n31irAxb+T+2hw6wq3woMuFECIeD
Y54ZYXSdIgQXYd7nHknuljNFn6Xa9nBlUMcEarMxp+DNBjsnXdAch1EzD4BUDIz2
Eev+KccHH+84c8FxbAUDKKNa0n4k/owPmDELwG9LX6D2eIzaJeY6iBaCR6HkDndc
Ap5rHAO8O+QtUhrWw6c5YsOlBeLlT/MnJfVqOeunGjU5caT0YUfBlq34+V7p9SJ5
JTmCVz+XpF8m36r+O8Dd7EjepC4ckIEBviMpMiPS8lptbRY51JFuwzaRXpc7kuaw
Ij1GWfM8TYhoskkr0jf7+6olJLyE+0NzA/zTy7A4xrkT4x6tqz2NGhZkZTJ/1nl2
Ldk1YRQvIjiYeMEd17sKktU41LcDmOsGY0RkJn3IIv1V5ndVjsPxbFQc1iZorPxu
8bxADWXFSaxvYyovRnh4zAVjPkqeojtt5j4WCesgpbQLdhrwYBKnP84xDqdj6qK0
rPahiq0t0+GIJ+EJLZv/LK8SHU9gxTvlX5SeufzT9BdwQ87QnueRXhc979AAI9Jl
9hBoPWftcuA0AUoMlvRIq2cZy/IALr3y2HKY9luGWPlwkuBHydwxP1dMXp75N6zO
ge5Lxl+x6CwObs5sL+NadY93psQfKpBfcnlSH0KCsweK1zoPYxVt/QPgHl931D5H
0OopGX/bbn6emCs9LQ5bIFLWPDDCo9twCH+I1MZMdyjEG98ilTNd057MRBlm02LR
k2U+LfEFQ64ptxY9/2PwZSRSsQ23NZ029JfcdgkaWbKfMhA5Tzjy+rvSnmK6yhda
R56g5W0qzuquLve6a4TVWklB6nLXTO00HgpkPc0KSzF3tsIDDSPp2eNl0tLiFWlB
9QdA8DqY59lBaSY1uMZ3H8FMBTMXcLvdTEwNzducozP10wkDWv58SgpFsIly0smB
Ql9xhstkLkRdJxoUbpOJ01Y4igz7GDa0HVQDfj6ecwR2sM3Dvf4Hhxuv4DVr97lk
+Vlib4kPSylQ4THF3MApgIOIvSFuINZ0P+cBRt5WvChXKUDALI4854crG8irIlGk
Uc6gtkQldRk6tZ0OX0JiobZOs3ooKU0DSHOBF93NHg7s7PQp5mLk155vebDzAKnb
jHCpayAJgej8NwsoaJDCRpPv8jiy0kzJ7vy5rPKr2LgpearJbKFYjnLu8ZDezB5w
EC8xAPK8sk53ypXZqwocrwHu1HP7ItCNRR3lV2/O8kFesMCQd4JNlmA324dNP0EY
HqQpduNBlrU3hgxJSLoKhvX80ffZB8ZhDwnUX8UKwpUDpwf6H4WYrfif5aEWKMaC
NKjPvHEUzAVHl47GIaLyqx2acJ+9cniM8of91SGwGYco5ri8Gex9lB3eUqAE6Gj2
G02LVk5lB95NcznJ7qc7wiTo14Gm1NsiCUgz/KZaNUwWTAV5i5onvTD5B5J4vYQX
rNAAa77b7jj7lkzt70uzDBc6IFsD2SziKhdlD3yFJ32wIJr8uaaJamQ8ENb2d2fi
fgvqxUlt7AbYmRIgKc4q/O0MT5QscYAZjWkGyroAUHyLfC4ACU17PCc0VAlyc+zg
xbi2SoRw6DkZQXFON5RbKEraIym+1/ID28EPEWUZoXH7eJE43T539NQlRy4G/Zbu
HRG1q2pz/eajpGDcyePwpeqHqwqUFoeC4EPbC348fg3LodQ2wfDcpUCGZYF52mOS
TWSua6TJ/q5ox9GN1VN+u2PypFS6hf/jtETPmhe6sZQA9P3tbD1JOD6epwki0rhK
yegl3hWWQIYBA5UD4wQoAN6qT2FrOUKt9WmKWrpgphHsWKWvMWploKeqDkmlB42a
5SpLc46d5Pr6AFeebfqCN87P8d87W0tZsW/Cik4UsHaR0q6XuYzZrLm1g9njyxXS
ga6nlU2nblfEDwurIEGKKD9go2y9lJCatJAbXf/yoeOOwo1Iw48YPKzcCcsyvgoe
XH41wlDdZE/v05gaTBD//8ZFANoxX3Ck26b0PXzA+kuHoIGDbkwfGnZeHYh88hWZ
IyvaFl9rAbk+cA5TlmHLEcjKnUGbku72KWTFahQQEFFgHCY2XTwbWCt0xS/i28A0
DSUWJLofeNJ0A/DH8Zl63ryyLfzFjttEORXPaY3/1e2Lcf04CoLVI6yBcJcsZjuo
3Bmjgg/LoyKy42ElglJN8KmpraQU0Qo1UUPGQazSAQfc2xcQF6M5exjHMgLIJlke
yvbfELnr+1U7KmJXaM2odf9mRBYdDIRqpVPsXImtlna84MKsPxlqRp6/8oVlZvM8
r0GQWNDJLnWxRILyK0Opf0tdDWSxFaBf9TWA8Hz/4sTJ2VHK46GIEu+6fdbya/bc
MNUXl7vK53fp3mHa4pU4Cws+W09ysLfLC0SUYUk6GWr0l11Tr1Pkm8p2X54BDtol
CQDIoBFWOhd7aCf+rpw/p2Fc89fq1eogGZj851nh/TRXdfJdUHNRON4DMpgzFCEB
1QYilWH5UdNjaYetwqTfAheEPCdfadTFejq7nehxcZLtrJSqdQd741+6l+jH6OCe
oknmNb9bPLBxhe+OdRh+xr9T8pIdI/aKoSLYg5OsJTZfO2IPCAhqQN/9oqJFQY49
+b3121IVi5tUjPXIK2TgbcgtYzEyDJinWOAg71L4CM1S4r08IHEbspC4XwIinOMV
TDKiF3O+zLiPt3h3z17Gd6K84KfF0MbupTllhFJ++eTqcrzILWjOTf3Ttojrt+uz
ok2kvRINHrFdr3hy/517vxRMAhe1bAMlXw1njqRYt5SpxeC9hT9675y5Vf7DYBOQ
H+Rc+EhTRybltkifkZ1Kb+MYaDaJqRZHwJRxV4gUsgsh/QdHM0gJMIdOa3vBESzH
50tBUlOZUEi6CfA7VfzZqiLL83VHHjcQwp9KJdKUovDgJo77+GaA/5wg86dNEGqL
kI/8uRMfrDS9YT4SXNaLfe2qDXDcgHYU3H/npnCWJohcxWQPSXbG8igqQLbDR7TS
eOqh3R2/WO8lRupGEzd5GuR6UaMT+1zZ9D12Tm2AhkGMvbCR4jqX2NvDx4v281uv
9GfhgOkBQi9J+vRAw3WCliEzPoTu2vitEKSH0/pE5jVZSZE9EngxbEhbVTAkjxZg
VRUCeCKNNga+lsB7bIsNfz0/KeAVuHeLIBSbGDuRlj6ps8BwCwIbZIO75lxEVzMX
STZinfHMvxOfkTw2VcCfxWSyuRXth4p9hrzlEdtzkJF77J63S/FmV2lx/qgLj55E
TToE6tgkhXUgWX5r82fXqOGWPfjjJxV+uzzu60+Tf43zDXEFTMmUks8qwmq6DTuO
T8ntwhJbQUuGh2LNp5xBiAAh6Cqd1QaugP0982El+IxDPGFf2MERvh4+7va3QKUf
PVzj1L8czaLbQv/ANqINKwIhn+eHvYhonB9KZeX3Qex1iG2wdmretzhNiWQm+vyR
Y2ntY4ft/K9U88hgjlnfZmPdPr/M8pAhE4iUOTS6es3WRm4ha/YkVonCqC85LCy/
V0/BiU30Dm09MnuanmAtW0vWHK5hnrkCAyHpO5oK0umSYzWTJnJV3g9AvRAXwRxX
cDk8tku25d/UXhQm7Gp8jewB+oBZ674kWdgcx/KxNPXbTk2dMreeeOARdvTFTb2c
uz2JQEJqcsLMPsa8QUpb8n4TgycnwvEDt42wcFb8qip+J9JOY6Zn0BkdOd7b+cuP
PuSQ+Pp1nll47J3aueVg3qHBxPl79IpnW2kH3GFaOLj7kzW19MFGt5oxnAXTLU1Y
yajh0/GmVPwdHcSl1h1MH0RD2ZI0TgJZDkIo6bNE7Tpv10PGjZi3QYlRfX0unRVp
3fBZDumsZ7mP4RWtKx7Adj+SN7EbSsaCZZhcRjcYigm9Qgax3mUVkvYBT6cZ25K+
msHxpCOej37ufH4L/S1+CxKLO5klRchttDL2FjQP3r4OE0L15ZwlKwo4QJesnQfO
jNkMdv05dnA85A2pS0sV26OteAhAJaH8ZOofkQTfCdSqS2NTv/PwAk01A3puN2uj
uyOhXEsPN6cGlc1ydT82l1UkvjHM+g5hoRNvNYlQ8w6jA/GAEzc9vapHQsNg69yG
iahud54zKBnnStGBaoyVJY3Gb98TZ1VrMX+Z4lMnREDd/dfI1XwRp5EX8myinppO
+F9Vg+LAcUH/3T98plh61WICXvNmWD9TJz66qpAFo2RgnUrflSEgA++2rv4NS54/
yKZ1t44hOtTtPCjfaMCdz2J5ss6CIt3aUWI7s96OfWaVf8CO+WOk9LK79Ijjf0Pd
cTAnvbVWGHa8/+7Rxt3RsYCO4EyDguYHQx+DqCT3vExDwtzssKRcgB5+DXb9BbA7
7cd090i99pRb2EpTVwdmWYBGUHSMYvQ+YoSriZZs8tnj/2N+QIEhKbDG1okO9euY
p0hUG9J7l5dln9+aN0gqCj+EkcZGza2SkYIVjguemO8o+pktjI1kBDBo2Cr+H9aK
roxGkLwOLQKl1rr8S18kse/1dZxmdOjECiq2Z0ASS9Heb74D5txozR+YtbYB/St8
+BiNTsBNIXc6Y/vlShUh84Tz1ErOHOQRnj2mWTzbJbqGcaqYMeYM+An90KmLcr2i
zGhF3yIKV9EX7sQ9yxkK//uExLA1MtOR2bK8xBKIvsW0gBME2vJTwiaaWpGkJfdS
SJf/ulePCk/iJLwhUm+koYuWfZe05JQOkuAW0O8wkY63rtriHDQgLH4RqBFXP113
HjHkqbAR0NUgPxIDNb1sCGWL0Cbh/DwHCJuAc8Nmm+AMbdRr+STQzm7/HAn8nsb4
7t0DsXgWuq3TnSArIHxKOKlCQHKoABFrato3/bAmrVcIDbux0oZodvTHZTbkfRtX
J/cjiasijVUy6igOLUCwCN70JFiIuC3idqtVYSFHT3xLpWxaYSo3JWgkGYHbdfd4
cYl6RG09TvlulahkpmNWjTKpcm+Ha2Z6mwd+MihIUEWA7CFf5+wke3gnNABzQQjT
G4qA/S77n9321GDpUixaYyorulZJu/Ekn05vJ3mzDy70yv8hVrR0P/HaG8oK00zE
/6Oe6iot7znkVEUi+CZR/w3iiNGNIIBfDfGZoBLgi3jTSecOV2cJ6BMOQu9W7dnR
WvkQWMJRKJMjCbraGGNxmdZOpwZxHgmOGCZ1jWEBrCGcEi0s11lm25yu9bVwDywd
w6p/GE3PEEdNINMDYGWwsAjC4UT2MiDLA93ipOq8U+4jkEN5r1IOwiTJu2CXSJPQ
iBDg/4UbzJ3+C3poqz65yJEkjr4tbt96KUHi7SPHp5JdLXhfxXcCsXLuzTy+gsNI
kRhitr7U5bqXqJxoOJnsi2dnkFtSIwOKZvRnBy23pNyhOsnmq8sMaqdpNSw6AiS2
XIy1nJyZa0X9a7FY0HJ9yhQrYYMT9BJBGTe5ko4lkURRiOdtIlrNToHb2oUMiKk/
sT39jZNdqTXfMnFsl/O0L0MGh4reHxzucba+Fv18AwEp19qmxdQeI6aAjE2jr1sO
0uryJpUvC5kpY2aEg5hq/+GJLsxR9rJyWASfGXom4knnEWWCA5eiUXM9ewgXLStg
RXEg6k/SPo6P4rIca9k1kYzlUcHXpKywLXDDt/bxmkzbElW7vVX491Q1DyklowXQ
NcLy1rmkivqCcYuwkOvd6YPyYjreT3ckdTT5wrIZSaEG1tI+y6jZ0BM5RBwkJ0eN
lBmBRxAgu0gkzs3v/Xi1jdxeT1r9AaaPTQvLdchIwNbL7lvFSwosLGoBdzjalNI5
ho+WE2WqtSrtdA63bEdIePpdxlkJ8VfByUMCeA6C2MEt93k5l0vo/NOaX/2YUCAI
SyT3m1BJLrCIvYW7XA0IYO2f61s1k7B0n7pJZQPg3VqQgxzz/slFuO/7Fz/LWG5F
tGz3QYTATcOd7O8vFl4RpoVdSeIBfN9xujfDTgW/RVwGoFWVN0rsspVAbYAz2Mes
0iDQfCgB6hOfP3U7cP9+FtPmeceCUFnr43iUi7yx4dsn0882gQI4zagksPn7Ofgk
M9Q189yBfklofXgiHl1RvQQPMYyybjOamWc9OPGufG8k37OL0ud3V3nbkkztVYia
cvEpWmFSRCoBl/ic7QcHZlQJ93eLpaSzVir+cX+HhNWKwcv9ub5FJv1I1HZK+9WR
5ocLdXAEx3B49HHrcN9fjNyLV0k2aihVfWZkAMkjyCYsyxw2yk4E4h6liKBP174y
ObZw10k22+ma+44IMPZbxVnsgguUrsAZuT5iQ2KtdDlK4tI678S6J37ivattk09K
VnLm11MZShfiDYmn5rCBPzOj3w0RsFU9JwJfQFZG1XCJ3xlMKLKfa1ANdmeolREr
SY/mWbCKzPQkunhWIG/3mncY7KGJO6K0mdj63NLAmS01CHHlkJ9GgPE2QT96ohC7
fd3gFU2Y0Qf3DlVoDdz+AmDgkyqzB+yKQ+ZPTIGPyvre/cn/NZExkNo6gZ48V7ia
1o1h/QXCtruZ1rwFRSaPkii59jBJ9Uns0B482EnuIOOPxcCBavSz+IxLgOtUdTIq
A3uByBLdU4aO9aBgmCbhjALB1XxOeg/4SoqfPM5BrStyzI4NsGekJ87syU2D0zY7
v7rpS4uUuqDVlimUPB6RYmYe33ZVUgvYOapcc1PFav0mS8hGhKuqgd+FFqmbVs3i
cAKgpBQ99MlCyfYihvrYCF//4NT8FZHIe7NCvKNivn3/Rr8jmN1MXjFYyAGuwsT3
0z0cNOK/CTWNSkjiJxnxPLls5kbrVw+7RcwCBYvVaO0um3/8vI9R48H8Bl7uuihR
c2zSGGKGL+jRbUInBJb+pwW82sH2xftfanp8OUAP0nKYbITzL7oifRhJpAqOH4bv
FQxo9ZnpRuIMrqlMu9d1ii3N0FozZKMCqPE8carhVDgh6D1C3HBw/fAUpXl88FHf
bM6jExmoROaLaauzIxTWtL0lmnoO2K82CC6JaM0bC2q84vo4+tK9s9yt57+Is0Ur
cDuwgs+e+gA3DLyLKwfJ4NvvfmJm+FGzni1thNq16mq7wy5XuPx1o4qPepiloPKz
oL/g53TLRY2iyd2YdACqYi6qbGHO5yqZCta+gOJyZMI/zVvtWRNTUovibxbcaGDG
Yh3Ooa4yA2VYLhcS8xOE0nX4boLlaR57Dn6Wyi16Ajm6QGNu71+gQz2uFIA6brLM
Pq8lfk9XrKidR33ad+G4yUNwX9sVm3VbO90Yb4hPTdeLZjbJZT1QJN7hFF1OlZ5L
bE6qBJ9nNDekhko86CbwNV1SkXDAXxOpHEyOaWp2YiOaR2itTh/nZTzqPqJjyzN5
RSpnkG0XNXUMSK2L2MxXZAWwxd2OPsslk/hkut3qJdGTVY1Gvfgjf4qbpwr0IMDZ
BduESUC+EEpAPqBwhsjPfMVYmsfSz/9BmU7tqTc/pu5mKVTzdFcdm6XxcZRQ0o21
Uhn7FbmrIanbwqmxXnBMvt+BND1C3QlyvHmiZuljMrIb2hSwMJuzb5yIO+r3+45F
fRXVzcj47jKdUSqdCZvYC2QL6RuQjX1gHJwAR7z27s/eGgZhRUc5dSl3WKlOUyYl
CezQ9wHWv2UquNnnVG5cU1fNycn/IiqpOUWMPHRk4QNuYiXSj4FqsgiH3WI3Vo5m
KXUtEAz/IiRn+w/joallDNECy5VmtCSy2o2qdggltzvf9jdd2EmkEZNpSk2SX+Ia
46fQ9M9go42W1Db9/XgD0bNRRYvy4yEnAZNaHZoyCO+tam6ubfpqFWwR5sicXfMl
ws5obgYntQWYLrS+f9hoZyfevLXc2TJoD3NExHnQbSMzl1JDIzkq40SZEn0IcsGT
+sJ15m8FSuBbkzVrec3pQD+/SJhTlZT6Y2Amm+UE/XchHqlixFHChxriQRq9vsdB
LY8P6YxPcOSS5BZjRIVunl7AkFoSZvTvsPPx2kYgyaKH2RZB8jfgtOFP3e8/BHXo
oZYwPpGt5AVneAtAOLgh4UjGYeDsveo8j73/iRGpRGaYtn4qoD6eeMMlAQxVtHk0
iAFZ4Dgj6Us4RPI2BVqKh1wBaJ5cSz5cnVmT1YoznYlpktbwVV/2bfC3J193uDKk
l8+QEGvrjGhvtgDCsRUBkoU3tBJS+V6pDe1rW57AUpcAq2xDXvQo1eF8O285BD7n
hY3PDHW4h8BWRK+fZvg2dM2UCSQpemQvFErKljO3XdM6AlMRqEJ6O1CvRCOGkJdA
xSGiZ2z9ZaRiaiC9JE6srQonkMfJpfTcypEMbCFZYln7zvTtWawskprIWB/i2gFv
O5i5CeMbU4p0LBwzE7KSSnEyE9WD1qaTa4JOHoB91XuDMU2cNY95a4Q9f/LTi812
HgVgPCLGsrrSLfoJFy9XNOpWWgJJDx8lQbBFy3beGo5As2VlsvyUw5Y150jxf18x
L4+n2ERIlyS1/2bamzqP8iM5iNh1Bd4rAlOBFROcufAlFnST7QAetljTBG34uAvw
q4OWAIVGlGM6Gr6aySyNDJyfIE0C5OCwNM2+T4mNE1kZIM8w1H5WLTeTV77ZXHkn
qfw3Ec9kofHCXabtMqbEwbPpiDPiNAZPLOVbyZ7U7UX4AWPmyi75Wv1V3cwpResJ
o4Hkzr7bEjEMKlcrgdh5sJJFJaqLvFgX+ioqkwkyFRQpUybW/uvIPmncANQVKwqF
Gs5eBGEVU7yqLpGK7qfk484EIqGKqYcTjAPb94yyhjZYODA0NCYvZhs63XpKBXYz
oeKRrayowIEPwzCtWFII98zNXFOTMnDEjr5u2d62aKAUtq0k8QTK+rxUcqMTCpzg
PGUDqRb8wznO6ereuX442TctUCiDgLK8eSezUJURNXuDRC4v42xx3QXxedIW2LOl
dr2skuqAMtbHhokRs/NgYt+415N8UUTUkv+U2clC4RN+RdMlLQBC1rQAefSA0Fnj
itdejuODI32foiq3vOTK0DBeDs1i73ESVkPWqERoCBKgRou2fo5uv52yoCiRvIA9
Ip4Q7taUHflyyqeDu7GSiHTVU48iy51qCGeMoj0UHzZI14sJTAhhu2tvGdTqQ5a2
CTQw/5zVT/GSz7AokcrMbzWZqdRXOIovPMaA/UzcTJ/SDar5+qy8kYelYNWyQ7At
vDFJt6eSD/U75bij6IqrizNkBZ/Tnu25mK015L0vGfRiZu8lmecuynJGwp/Kd2/M
EFHGNIerWn6mKyxhYvqjNUodwemIHHaH3HkTk/Ad1SxV0OSGJt0NpdMZQeYGTwft
L6muAcCMgUB+f9ALYnFZPGPGfYkwXZn7o2OZzmEnplB9312lM8evcLrD0ZsqL4Ok
0cd05kDw9b7l6NH/vE2VCWLIfC52z+Nhtbpb12VzldvBX88H6ZExxG/Pw8Qn+azB
IXLAig4TFz9/2PGR6TdK5vOrfSCwQ+5KhkLwYC6qT56MxyI55uCWalNTqq/OzHzE
vHPi3oLL3ktKZLOf1bOhsHhwoY6TA5j2EsmU00XmgsWFXWAYaXHmhOuXLVR++5dS
Yyz93HdehEbTQmh78LzcGMhNENpCCANMOC3ay6yMi79DN4q1+h6TYAqj6kFimWGW
bv93zEieHcRMITm+r2GHkD6aonaxqlsibaUvD8HLlnqZ2tnFj5LEQG0bnKKcxoRq
Npk3MpOROd3ugavixheQpLYYKovTWAKtRpeT87jCuBZavJreo937TObzsCQpe8mQ
Xp9Uh6eOrKMDleFvDneSSc0xWX2oR5SB1qh9edY0ZwUkfu1jEa3Em2QlgP2/t3jM
r88CNI9u4cemqmt+3GhrcuwXtpSL8WI26MDJSJceZSohVbmzoI78wkwBhAjZ9Nls
31vyoUgfGapf3U4GlpT+7d78PhpYjt19ORyFBisauaiVeklPVTmal0U5od4aFBXH
V/baSqb3L8kGdQDYFkin3e2jqrbPJOIpGmrrhprVZkRrNrL5fvM6obdNHwi9ZmxZ
sesWKmmL/DivCzt5l9SW/eAyl8+EElYxLXVHs7Dww7OyFrE4O2bAgk/ZhEqllO9A
/UESfeptQNCzRSNw32d/jYxdGWQwumA74YOANxc0hvjGr7ZjkE2CNKsxf0i54Cf3
kmwcMYPL2M8hF7dEdSOYpUMUU/YpJuB/P6OOKx6fdmPu/F8TjOzxJv9ORp4tiLmp
Bu/8nB4ZduJoiBlEUy9jQ1nApJW5A3Fj3P/oCuTUSaqNwsTLm6zSjEIPkFczNV2g
3qGIR0G/ALOGXAhZSWHePwbPhgQV4IGENb3Uchm2Dn2kTyZBxbO2jab4x4y+4Etp
QeO575f2J5VQsDbGdigZ9bjJhP8KCxdMDNuMENbXUYPVJjAwcugmzrfz0zUcTgmp
eJhukY4fvPqmp9Wau+ZBqeveKmd7DLPQzUsibxCcUL0PPr1S03IftHADjHdbMLI4
NozSMhHlHAkbvHp3iqB5axkbq9Sgdhwi+p/ID1aYILkM4tXxmPHY/M/fQrceXTwq
eso4fR/IMwMqfBHpGJhTZ4yH8HNmkeFDwVoiPjkx60X2XeZgMWC3VyNdYbu5HHFr
RGJY57e0VStmN0VgJF79Kp9JjVhSGXZQQyRnTGh4mF8HA4u5/1z9YZRWsfX7971M
eXt3KGmofDv1c7U0Uf03Cj9CKQGjQxNV4POJZIGMTHE53r/pcoNgsuppZh7ipwk+
oH0Eu+4ooxTNUfud8T116fT4qqdWGs1S7Do1hKRBkKPi0Mq+8uJAT1PjpzLHol3w
s+2dHGsI5wBSDYpC/DkFuABTpVrGgrr/xmUexv1tzudy9z7Kh+sd6SvtMz+Nz2Dv
8up6GpWV8ibc1GS+O+kWysogWRHeL93x4um9K2H/PUWUFOIZJ3ZEsSuM2KpLwe9S
7pYu3WNfg4IXn0Z7IQ+j+upshgg2jq6M69op0r3vsbrQXcVjnU4qVqwtOx81tDb5
ZnjQfdJzpKO/p/5jcmRypFLA3pz4fFMSzb2ZiHEnKANxU2s6RY0AuC7j7gzaFWXQ
uX0jHQtS+HvXr/zlyd1PVGwuTlY1UuwPeg6JVnbkPGqvyb5YMzqAeqLT16E+0dTe
Qfaq7arRDwhU0ffpqkKxeHsuSQY+YChgfA3b4+0pJAlcgN/PM63KydPlFH22ByNv
WrAVQccqgW0N/xVbBS91MDKOee/HYr5bcWIJt0oXUZY7lrC7NOFZY0Rl/mHVnimP
WVDM3yidZ7mZlBAB38VdkaVswDETjmxALmmc4Q6pJf34c1UPr8wucj3zwOe9Dkop
E2immMD3Q2Mw97p7N6vfXEDc028cejLFgZrhfbqM5BALqvjVXbDXSeL96yHNIs5G
zNKy80JYrZ1C6atJKJTdDfUNcNJBwcxAleaunUPVZLYoy93giquhycdcx4Cm61oM
SqHYUg40GPkvC8tnG8u4PdjVpbFXJEsNf1uLpGNo3FLWX9AsNNn8Ss7gspb7aufJ
g/+q9tC5de89Z+9vgxi00ThjPRH+61PNNitNMMg5MTmJCk2puoO/GxseS5bxIcMX
xyHEUvPiWcjR8LfHO3juWFadCz8oL1REGr7KOgO/Mjd4Z6WOFRkVCak7IIFX9VhF
bwyS693YWSVj1l3rivd3cx3Zq2PNJbNmQfMt4v0nzVlbybDixDx9hhgrxGv6j+me
jRe9JSV+jM3cDcGIGneUffFeCusWlcqBYc1Yl8POi1MHS5RAiAqA5NS+gJ7LYqT3
JX/5UQMRWEXkHbSZnL2zk6g1AAk9wDOGYdkn1QxSDSK0KCb4jIbM7M9d02aTY8XF
cFE32f7GR604h3qz98rrqFsnzN0HyGFBKcxmX2XR+//m2ZLuubEJrPHUU8SUbztH
6JGcNeQ4RUhhcNVQ9LIBvVNrWc5eLI1NkWSR5qsWVJDah6lf6PEVZI9zQBSzkfSO
b6Uc+8dIm5QPX0mxST5pDxhPVSZaqwK+3Dc6L29AVRNbvzpOpIpp483Fh6/tq/KK
MLDL4W5BejDyTtpR+KLdqKcXwjEpML5M9q8kjqj4yQZD0quth6kdG+6DWoOdEwET
EY3Rl5Ig8IakRvq0Rchqql7GM+vKHNpKKsl7d+tpp72+Ar83frmHhcQ83Ztgpt1G
u5f1llaSzf6mNY9CVmdPFs6LnlgZl0Z/m4IkxrhV3xe65YCICHr8wRb1w6DaPVv6
QfZIIJe4uwmMqhN92vfF9SlppSi8sXKCnADboE+isFN/OraiCievIbhE8bXsOcvy
KJiplVaJmBj0etHutsdFx0JAddLCmmCOKC+BE5onda+J2v88j4XCzVCfoInQK8N+
t2WDmpMhVSAbf7SzyQuJ2hd2qYExXzAU6Fwdo9IrRzkyEFz5OvnqQTuSNLNgQsKo
aigzyNX5t9E31FMhu9g3guZWLNnoO6skmHI/sbXB9Z5ykKqnpz0JqoYFPvt5Ad5u
LbV0JpXE17IAyVzZsz65Q0MJjNs/9rmfdphpfRsHiKHW6VAwjzsDcaecfITqmA4z
zi51UrEUEBqV6BNeR9or1iF4iFruq6ercMZwtKZt/ZVVZRwHBAfiAltLk8vpeNWg
buCKAoOT4GLG5TZ/nAueweJ00lJ/L9h4+CFSwVr39FmxicnkPGG5Rosf9ebbyS4+
W4wfFCcyLy3fWo+3iWCgIYloTvKXTT331QkfQLBOMBy5n+fWBgJGiaAlkiKJiwU0
QZ21dv5ZO7gPsWjdNEENc2Tba/mJ0QQ4270RTCiwLTfTMYPp0dSSk8GgD1Yy7OF3
lEGwgJZtCZlOhRsc4b1/WzB+GnD+diSgV5jUI1impowyLLWy0HyIWVj3jus/N2rM
LeOMwfD1/5wDGEk9XicI0VADAXqiwMOmLWg7yVOcjvSz02XHfuBvrv3IIJNp2aN1
cBG5VS8V9vsoesFWYuFqh0YQY6y/KEz/auLUuMRrRXNl4Zv8UzKXMXMov1tORTQD
Ge1z7lnx6pW6RnX1joiNIDH4nrKvlJg+0zY6pwaU8qxFEr7jKNL4QKWBdIR1XXRn
PAjL15gKF42IT5MDFW6rcUd4tuLvUcQKylvylDFSBYmGwL7VfF28BdwNnwfXCUxa
FD45+1wn6NGeT7dgOfbgb8kGfG8XXwu5+OWcFd537aE2fBmtNLc3iFEqom+1H5xl
/cGcIr5kGhCh6Gq6csVWs21yhFLg8Sr6TwjGnwDMiHfbSTON2+vM4MhvXPAYb8hr
GD5YDvPqAChGSAROc6k1wXPAt9GjD1QisR0PqE8rOZkjfpNx3cLU/B6B7liOvmDO
FhWlHxuWkYvsYU93uahgPXB/UJ+Aco8kS7RY63bg+5OHv2IFIqDyCBcd+aZtMzFn
TmNLdUQ8AUQpO16zHR4TSspJLMG5c+bfgK9Rn5lFfBs6kHeJ94/J51fA1Kwj/IcJ
LjPbVm12H9t4PM8q0cI06HvkRLntfv3Q4S1LHfcz6hw=
`protect END_PROTECTED
