`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ra0Io7VGaFwictVBMzbaJx/X9EXR94ydMNkPM+Gb/XCZoYfNfci2x6BP92Kg9FCC
AM+4IBlUvWy+mlRgHtHLfJeqflUKUCe7DugORrgQVmkF1iFpF9KW/o1zBZjxVFvM
Rz0BmoUFx/BwGPv5MHedOse0avxP/ZbrlGHZRmUo4MH4AbF6WNtV2VVfyA/SaZol
eMeQbTwenpSQzBIk+26sfkgeCa462nv6uAHU1OcpXLbpxPeKg2vRhC93pjk3MrGI
s9vm51Ph7ZXogavXm4GSswX2C1ANodKj3tC0bVALY8TVN+PcjdKWFgGjELR1X44n
bp+nQuuUk80E95Gr9dt/3arqKPHGPkAncfkHb+3wIceY+9Zbt+xy2MQ+VXY4XVec
8sC2RV4uvHWBdB0E/LbpAsGc+wrgbkE7VpGmwTzReS6yr/1oIEQ5PCbXqOmNch/F
/p21QM8SsC2IALiTcm2QzM1ePm4iaRy2DGKReCzWgVc51Ld+P7UNppQteBLZieOU
mqTPIOJRk7DZARFkR5kPybzSnZ0WYk9vejXar8cjWGEcGiYSWli5P7FpkNwc0CSM
+wlSinjdFBVO9ShWvuHJq9C2QdGFRE2m/VtsNAnZ4h5Cdm2O2Ta2aueQajb9zEt5
TEOgRt7gO6emrbb4sU/+K7Ex6J2BNTfYS1rNMHaA5oOZmcJgdPpT5PHbe50dbcAJ
7DNlauMmPTLui34cIpV8r63577uvK4IFyyYKrRCZ5TWrDl8ee7UAEj2GcmYLIPCW
Aau2AaX1N+c6m+xT2U+3MGMm3Mg28B/hJYM4Rpu7yEH+GwikuWf3PYrZZbMowm9r
26ZxEstBjmE7AJbNRFa4Rh5ulicbqQapZtYfQP9zKVOKvFg+c4y9/4wYmcpPRVpI
o32ZlXB2PvERl7B/F8olisTHwAokYZutnABy4bIZQnJ58DAl7aDiMlbjjQsClbjt
ZuoQBCM8zwkEydw5vQLQWPjO9hJuncGVGALXXapoAmmMpNCyIPxqohiYPcigjfJM
Nk+zpNBTptqDu9K5skuR6NPHYEt+ZB8Kl3qAq3Mf6eb/19JqUpJjJFKdJwyEwRmG
5Zq3/cYURW8Z6UKn7uUY8gC41ZEh3qe1Tp6ukxsUwU2ug3Qbpk3UPQDy/1qZEsGr
7Ir0CbufazPeLGCq+jQd+ieg736w2ZCPy7IVoTqUQ5LxSFivXDVnRuM7rRzyCblN
vpDZxF6FqwnHdW6cweUyGccHYBwCJLVnIyeMXwOnswMMSVZWFZY1xAYjywyP+IjH
o9fNRFh7dU/1nIZ0pbKk9/rEeWMmxa5F+kKFzFVR2xI=
`protect END_PROTECTED
