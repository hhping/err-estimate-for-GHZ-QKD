`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQGhoHJDm8NBP+XEuR5LfY7pwp9mBKuLzMFvXpoMPGe8MudIbfiB8FV04GXAMOYa
n1wkoE43/BBz4hIPvJBWfmtYaI4XCKTb3EfJn6ArpRPuFPWf9S4mIvarhnX7j/SD
3A0FdPeKCcaY/aEfD1XXKjZGGB/olifCDwVuDiefyhYDEpFSm898D/odEuFVAXhj
ZK1EkgZ29vpTvou92fz3xfXBGfN9wxnLypFSqB7A4tJPz7DLC7h8Sl3Ct8ezpeGM
Dk9ngjcyyvdCcfNphS6zyU961zUxjQ1TgbChsu6FAz6ykRhr29Xw3i4u5E2sXCZ2
od7KgIgV+WrD+kEgkEIGB83Y3SzgkEsgmYA4WgVFBfBoS/Pb5g6pOmlrcp7q3IxJ
ryrgsrfc2Ewl62/bKVo/pdNhB+HGvaySqXlZRTmenB5CWdTohP7HC9ZWPcpCdV1r
Ai0aaAl0yDGeSzxs7xeOblykn8ZEE/5ADImQgnIFFECsgeXzTY9YEI/C4//iqxeb
hyuoWzZOcqPSKAJt+7v6CWaUAzeEj7JHDEeLTGMHHIS8SpPme6ZBV9bt1o98nlgD
xaimlL8MHZ7bA1rlA8rE8e/fPBxQBCaf1+eu43eYYWEp9MB3suF/DsG0Hj9YmCOQ
utURYEK1LKF7g1WSFo/eV5C3llYLXydSpEhGxNxUv8UKqNE14ggTdpflheYxH7nK
r21P6La7jbN+p2pPkuDkFaUPca0zzzeyTcUAw5hoeVfIKJgLFRZektbhE1H1tAgm
/CSic5iXgvbJqBxwzQUzG13sXrROht2ibMYwUi/pFwxEtPoha/L1Y8Z/PS/sdjfz
sNML5j8M1PyPMi11b0W4YZa8GgxsnviBiaR6ty+JP07LDaFDBToC/MwLyl1aj8AL
1Ld+RscdMaCcgaUK2zVtDp/JX8GIDPpYBZ9aEHa88NXCH8Nn+abB3Fn6VRmqonPx
i5C7cBu/ZSRWOBOylcikAnTTymkJn7UgIYGOahofLwevH0gMfbI6MBs0+7whj9ed
jSNTHqxH2o+dSt6zmWp2Mhk8ib92c24KHBlaPd5EpkcJQxs39Y8W3X92Md/Jww88
P1qr/YshD16Cu+SdEyzoOPlRzX6VzZ1CWpAIpNY5qGvqooV0BtsrLUsXWgAGaK+x
M85zwRLohRavIl1QpnCPcubUj9BVx1VTu9agwYVdA91y6ZaFh/Veh9lYRWt9Lfld
8mMmvvMkpntrF93XfZhGKXSP527WmXF2BSG+5RDB9DA=
`protect END_PROTECTED
