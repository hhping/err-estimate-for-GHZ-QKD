`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkrCRqwLrcHs8GNvjQV4oP0ceCQ4xoWIrdSuPvF50k3zEbPnxe5j8IPcWm52c6ia
Sf7Zp/SjIIXdUTiyl5OEFh6ZVcaZLwmwS0W8EPiR+BIVijDV7OiWYzYTUVW+KS1+
QYz54t3VS3THAf98gDCf4QrUgO3uALqfTpCXx9T79sKIM1WtFmanxHuyRBnok0//
cgFdJNDrFJL69IHuxp/ISFydTf5eP7d5fvjyLyOBNASimEaw9GqDsYVaMgxxt1br
8STsQWHI62PzIAwfSAPZRuCqs8NEQR13+qVRQAMZMKKWNc/eMSoomrDW+/qWtdAu
e6sMHnzq2ElhaSTdHPZd6sQ7dfcfTWAU9WH3Gi3ZAUFcOImr4clnTRkDeksQdRa/
Z1RdzDeMnIyqMOs4xa4Q4RVrlELt6Iwb/wKtdGUUOYQGaQlte989HeZssIZ98ftn
ADl3rzYjbH6rTvZXfMKmh4KrQ9kiXOnlRBAVarUVd6JWWc+/P5lzHCBHIQP58ooS
ENO+lAuLAMpLyFGR40wAC4Ywe1kN4Gk0rNHIZ6pwSNdb56iXWAZVkFjAA3Spfsud
h/FNkeZFVDW/1CF9zw4zY09KtrKY6G+y9ghOCauswaxPwj5Du1FvvKdpejZNV7Dk
YYHHEV3VKYDtiOS8BuAx4XylJrlm8spVk5SBXQ7DONaBs8oDaz+7ctCo1fPp2T/K
0g2nS/1hys/3zg8FD3wjUCbVX7V7CitSbbSA05FbQ6evlFAqdDiHerLKv9FHpbpv
ZYVsWbLBjX20WUG9Cm+TcnNwYYpM48Dfb2eV6VXsddOs0RpQvDbObFZpnm9QPJUz
`protect END_PROTECTED
