`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojf6Su0+n0va7Vfh6oLNc5J8WBCb3k4loClPLQy6MkS24cVm60WP+iFDR3yYPOwg
8E4EPnRQPWgEJ8ccRSzjH22P+VQqG6QRHuohx48PC0RpLTYVNAfv5tJ7AA220Lnp
iexrBtrizR8u0iQIGZKhiNLbETyu3w/w+9gR/ypmH7kpcPFkO12N3z4qCJuyTwDi
521SzD5mYXLN81YMeAHdm32JEEGZVSx098mwoi3fmE/6ipYZTY3LwFyq6S5mnK+e
eFRtThMqFmTgFczQwM3ribMFx2mbFk2KpLfERs4OYPLkwrAoCpfNLBq8yzRwI9Ps
iAAxv3uvz69W+hvjuBnCZEi//m5J066oAgABvk2fTwhjCWZJ5bPF/eWfER/EC6Zs
zLT0f+2yKJbZVRDeSnNhfOhdohJtQG8DBx7VfP2dtJo9dl8hgJqwWe+EL8AXXGYh
eKDI0Z5uSqArvlCNi3O43YtBkzN9DN9QqMMrBgB+DC4nqsoJdWiCoeG8uEUyk2TT
3W+R3MZg+e2totW5GNGAEdsHUaCICn813iHXxybiMD16j/TziOrM3uRi2L+ng+5V
JIIJpjTLhEH0tQpR120AdLk3+P6crVYWbAGu4SJSYRV/o86zHbrtd0pymlZ0rISG
2NeJOn4ltVCeJEDJ4fJzvNb+H/Hsh6x79c8+QNVEX1QmAqQZiXGEL/bp28jlXCFl
T7NpK4lF9MzU94dHkhSiaNTnF/YeU1Kfs/+zXYinFHCO7XUavfqc2rK5uUE9MmWd
/ht3CMMfgKSPYBiY6ILqfZ3SOucBN+SHqsTuRQSqKTZ+JZNGQifsJzLvUg6aaZeQ
SjFo7lAddfLaRuDyXdq5eAnyCsrYNAnQiT+CxRQuAqO69YauLKKeGeIfED9TEvH0
79/ptYeAts+KSeN1OTRnWg8AgLOpLgaIoQxgNkMLjnJXzAlXPIheJeYTigHuPMNz
C1wMsDHOOnN4wSUfAh9xl7ITaaoQynfsqlGifMwNpxiwrIdRuOMVab3bUuiefy3T
JgCLecR3JxnNI49saT8Hw4pReexn1D4rlt1jcKxcjOMKyKUzmE7Il8/Lt8qdMU9L
8cmFeeLs9vzQBidOlVVktZXftp/FsJsjFMEiHoOW7If2a9mkdaiN1AbQvKME2Uq9
VbyaY2XbdO1heB80f/bGlkmb7RrCNsnIt4OjwkeG7mkCTZWJRg4wkt87FO4hAdbG
8VwCFoQWWJN4SG5Mf3+K0GES5J0LrQ75D1I3x0QtGGIpn6WgecQannhb89BfTMrl
hn/qyvHKh9Xea5yzpYSBsGbYHTfIFMVMaXMKnnbXLG75RFPhYz5qoCYmM61Y+ufl
IfBxmzJ7lYwnfY46SPQpIgyThOZb0twyR9g6mPjytj+Kh6ZZSn6wGYIvbUPuvI+6
6+ry2SOjQAS+l0juN7l/acXuY0PwHsI0mrS1WqNHx6QNWeFD0E1AftX37FqDBSjj
W2OIAfusF9yNnsVDXdL04kQDbukG8kR+vpyRdY/TCKkgKnHeumhVXGwPKUXxNjhE
wGiEW2P+rZjirPLI7haB0EIlv12PjmWePq2iatvDbSKuaHkirJNDGpnoby/x0YzG
Yuo6dYNP4Ui6hp6oEMMcntwzGhG7sNdJFMvKL5wrk861MJseGxOUwsuJY7l1cdKj
zC8R15C7zjy1a1P/Efo/LvYYFuzxCQYmhMfl6i/70fykj+ZAtf7HcCAQWrQFG/Yz
920EyURoy+hGk0MQE556C+7ua8ecjuSUqhmz/fkB5RlgOPk3NOO7214XFMfDWpP8
v5i8vM//GA+Ah4GsSW/VXGakBdGgUbhCpcKWuKjJqvxmCZIflJWkTgteAM6TR7ba
SOQF0DyPYXviSW4ujrY3V2hW7QYf6ts5rZy4oeMzYPLnchl3MoLA7OqIV7UGrL7L
c3SZaK8eAJInhUbifjQpIHzGBytRlbbHBynbL6OZE5HpfEmjwZxfUf+Dgt9FPM90
I61+OytsfFiyDmg5L+ltEjcwyMgmmEZm9tnJ3ahB/RYcPM/LKfNdhjnVv8kqF7P4
ZuQxn1xaIKvymaWpV/cCSH6yU9sP4FN43+HY78PDXvIyVpCCnuNr/IYfrMnqx/Re
ovxbjFOazKBGMUCR3pdNWfADp8mQnPbWYyGEHWyD78joly79Q7mIC7M4fAzXWbGb
2RZPI2XYBnFpRAMH6qRYAKOCqLHxvXdHmklGzozUljjIarU88BDb9lZo00+6m0yV
YMYXhhL6lSgcpHmGGtodyAfyq39Yx9e+MFdQ8q7gBz6TwkXrhZY6SRSqen56a4Tc
aTLgaLy/nkk5xSsRPHuHmjECgt2GhUUdPrecohES1//q8/xJjYPcQBWULpQv3f8f
pgKxK8ZuSSJyRaPk9r65Vum/W87JQLXyd0X/vx/gdOAL+Ejkzdd6YWH7hmMQ8hqR
PnQoedaU5n7rs220AlDiP6HZILiy8CeHlsbeYOwTE9DDaSxIVNYHBVN1uWyIShJ0
VXVuF36npE3MQdtXWxkCaGqayfJEKs7XoKP3+KYwk0RxO/Qlrk2wzKDT2VioXC0i
xxmhwQITjcc08nLVztSQrvzx6mlAm2GNuCHmUFfK4nJVcdFiDcS+lSFOqjmpwqHE
J0fgLk+Tmq7q+yhcpTwcHspQdimi+OI+HK37tT7Xvl6i5+d5t4/gNufvx3WG15dX
BDZMMMPvDVMa4xAz08YJM2GiF/YwSx7xjsOFGuUTd3l9sXFtl4qwCW6pnFMIhfcg
Nq4weGH+t4lAWBjxmRookEMZ6K/FTnX0IlrlREK7sdWG5c9+SLT0UTUvY7REhuNE
jmGNh7mJGAFgpjp8tgJS/EAHofpfyXvN5s7kt8JZjUcEjyC5S9eOcrZwax4tLzZc
uVvEdbUuwnCOY2caq0ZFPqx+4jAaclJZ6esLU45BVL2dWs5MXE3x5sPjNr25qATl
nAshvI2iRLVFMoPcU1FyDV7NGOWVsgWD0IX2XxSNWeU4AJNWqoODhjEV2JfCDva5
JZH++Ewiwv/Gh31pjVz67iPcSwtkAx7k6rhzemUIa1tXTqEMBGc3f/XFf4QjhkV3
jmabJQeSyCbn5OarDc2OvBg+3u4eUJgd4315TZUC1PMp8C0vXk1ciNp4aAwiiD2n
jJjlUQ7G8Q62yvZnbmkctGoIoxUTsM5GcUpxV1I4d7doJ3y/svinBIufnATVDWAo
5Hj3eFsuYrSCDmWWSthgu2qPaLRtmKTUuRInOKo+FgP/fyihfAg6LcoxOr/l0uld
0ncL51igeZYmlrzsGqyoOjDg/vRTJzSOjRNEzCGsRdH5sZPynG13gwKxHP5dclE9
05IYqMKoTk60pdQ/ZbbA9eMaq5x3ZgcXzgKiNs8syc55kYIRG2EygOGwev5bLS2V
XCirzUbbhEuSAIcOG/7n+ieJwaB8HkxzPiUW/2Cz88eUvtYrBB6xglurmT6rDUTe
a83KRas0sBypZZJXA4leBL0+xacblYAxJ6AiF1uc9voBe+VggmlDi0pC4j3SQUwY
/maq+VlhH6OqfPuD/JO6/sijIKMR4uLD7SlC4ufSwnWbEBe0O+VmSCtI6HLpXdws
YBbIddXZvaXdjqNpmuk3jkMx4Tp+V6FnhvaMW9sVid3lLyrfWbmuXNlk6HNBHNgc
N2KrHJ73US9hdhiQt/RpPYuDvuGithPUzkIqt70DEW+5PZ11Iy9YQ6Ujwmyew8Gw
v0laZJ9MxK5A55TLymQnx7zKtG/qGwCSv2dqS/nuZx4v8QC1V+h+rcXp3Gxsn/nO
OnZCGL/yo1bSACy+bDHGiVBErOgU5UWf8SGSk2+egEGBOioBMUx73jqtv0t4dlIi
MQ3lEgK4AEDjJ/ALcp8rhwB2msuezb2g+sFDPkGfgizonOcxHV3gi3ZRkBETzbSM
+ABNNFRH+EfGO0FvP/v+D67YYgdChDLkYDXqvF4eGWf9u3r1oGKBhEKib7AI2x+F
u6FTcqwvsc1EpY33GgMhnHiyiiPyw3gYVg2nLOUsViAOY6vgkCf/KKpX8wEKYEYF
PJDrN7mq9PQLaR3FOEGM3IB1oQVwUostmrxSGEvWwQ8AqeMPg4EOLAlypiRTi9mR
A353FWPf+5KnkEC2VzbUTGdimaMSUkEcFjtp6sIQsdmgwxD0lMYR3cPT4zFZmFrV
IVSqxALjow3pI/gS70xbUlEvx6ZnKtbc456b0DI38WcKZxnzUqcTrkwQPTcgwakh
AVZiCpYC20je0SdR1GJw7uvOYRD2wW7oo1YtIfs7Et28bphZNW07KiZCEnsYVzoK
nazaDNSVvMIXphxBOn6XtZSu3YC2ZOHM4SGP80XP4ennKRibVmP5fgtbrK+wLVNn
baZBhw4W7gNb/kdKwkjBJGP86a9FSwjNnSg3/qNL5yy6KRaW6cB5ip0gFzo4/CeS
Bk0NBNvmYY9/4lZZodiuTQ8NTEKQaVZjYmHR3eTPBFqCgLTk9IZT+DzQrgvs+zi3
mvAbS0rLdB6i9+Z7c20eb+x8EDcHOnls8BggG39o3iyVf2z6NaeUxoqYfMnvNFyp
L2lJUKWw7t2wHTMKVHvYL1NWHU3G5cfGWzGE6CxxEjc5sHXI0amoGfReIzqjBRUT
bfApXZFY00xDs+KDNR3aAtHVGRwh4U0Hg7wQGeMJnq96fAkOJrWYThLLaE9Y37Lm
u4RfpmQmDqXh90nIo53mvwk5o3Dy3MTQ/wnzX5/k1TO+NfIAa6eGhc3ADaHBynea
NG8srEUFE2S8P9yY5biSELFOw05558mNq65KAikMd8MKwI9En58TU1UtLEQG4Dwb
iiOT48OyMrgfHsZebmaWhcDD3H9meyutM71+bZIisISllGGQVbF7xCGmf0U8JKIw
WYwytxK7plZyL203xsMiVhSeSdA8o6mVpgsA7S5QWJyU6xj/asAah73DBMwwiOXD
C5x+NzVprsbXhhQKur+BL4yK3gPVyoLEJNY8GbD/57dADfy7SLuXdr61tMmQkOkm
WHMlF1bCUakCNrWKuUUE1hzS7IH7w8dULjoeFIGQY2SWs9O5FSuHHeD8D+GeKFcM
fLQ5KwGmPCs8B1L/PSu5QRB2hlcsmh9Pf+JJCDj2dm6tjeFbm9FfuHM74jfRNU4/
SYNrjDAmEBnYdId5q+vKQUiw5dpllgXD0aUCMKZV3/XTZFc9o5GhOFNjMU5WGnzq
VyKnRc3V2zRwYyU3qDBMCA==
`protect END_PROTECTED
