`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EoBYUaoPFKmIhEvmYL5wYcjiAVp5B1zowCyD62IoJm5YBAp/PbElWH2LLACoceU1
QvOiHhMNSFt1dqeWQoF22f5OmX2GYWtUUGFG6ndReAuz/qO2EAJ1SBkuFxRpQMB0
9uHMvXZZ+7WEF+XqrXakgkyK+hyYm/aLjnMVe0akippyE7nOguYCRkniayT2smq+
EKu6JwWHmFCncn1aj9FZ9CIZsgM/5IJH5RqwJrcZNNt3/4TEAXG814SyMZPp1AN/
MbVAera1SwqbU2p1AXcCNnkAMJwIFVv964DICtP4Os9obRna6Q/9aRMIWqdcttFF
gQtJ/Z5RpEWwI5FxKTJ90QCTS1bAgYnlsj7tyItYfxiogkGWEC0fm4w6C7SdVqZF
eg8NZup6dlWkhUxx5H+yArHArge3bfu24swiyTOYEYMOTGHLq0RSbcaZzhw8fPyO
UyCSVnTx7souZW4QCDDi7wpeaNDSTUMWFma+D9boQeXE9gnIMA/ucUpubAhpv+/N
orcML9mh51QUiQfGgOpdD8oygSHtf+LZvfuq+LYTkP0J4Lh+RnwMW0XPP0XgxCz1
izoSO5loCObBKoDcRVCUEWXygq30z8P5Uk4VSY+z6gSDVy/58iPX2zeldiOj7O1z
FK+mpi6WTHeJPOpfwQGaRwhB8uQaHmyh8XFP9l1d+lxdOesGnVRiOrrfS/lNT45j
tfTngSkLMxaU5JH3PukYgmvyKGsInUxRgToZqRe2sQRhK4K9WNjHjC5DsXsBJO8C
P7AM1jNtNgsqGCSsMzX1SjkBs+wQxuxAz2XEcBxjZR7Tye0CNs6J/T9gPqATJqqn
YHT/OeAo1TuumtRqHnx0DoqMX8Ov4DXetMipthjNo4ElVDJ31hnXX1jDC6yrTQ2j
UZtG/uNTuHkabe4aN2kHDPMVD0urYyk2j7X3jbS3WF/IdIZMadOAmsEp2SYAr+Xf
6DKWwJ+MDWBQSlXRcwY1zj6JfP77JpgHwBZy4NMpTqmLQzJYVacUC7en65c/PHQz
ar6k8yYmApr4ydbfHE8GrLKsDYtJGblvlIqqi5B1HNE75BL5VufvlaeyUiTXzzdS
FWqOEixEd14qv1qeE2roEm2bczYEVkAdXp52YSG6vcyDIyAFhXkZLIHgNzAzNy2X
UsJklB2dudetoOc5mZtUy+122FC8oFrmPqTc23jpUQIXiKoOBtxuaEjVFBGsTb7K
iV1Rvqo6a3DalwinlOu3rY1tVPX9tR+iSmKMcbCn6njc9zdiqEIh6EI8zK7Kn1JG
7NLzLeBlhehhtPQ/0TA6j9dyHgHYgPjD3crbCkZRV/qTN9w9k4rLeZvMt06mOTcW
fX0YzkAdBkr5fmRRVBKL5tj/lpuBw5OLY+H+Vgu7oqkTU5+IZBIBj44HSpdLVWen
SFIXsEp7F1ZRrAqVxnEejbZdcb8bkukrnnWVmWq0FMy7qrhc7IXGOgJhDqu/NbvF
EEJyKiSvyqO4HRULbPcTBWuv5GNHNEb1HteioBTkzXacDtdvPszrHUq4zi1fui0j
7izewKtetzTynJagvtXDkODpspqEXyl5SkfJGs4h6fd0YcyqMagMF0+1A9KX+LL1
4fhNd8fyNI4FC06dldbb/UHBHW08aOJ1Ivpt+8em3Rpe3+vfeap9XbvLbLCd9EzB
matbcWt5aVcGaqb2LVRNKHXWiriKAKVU556zQ0uuOYxkwdOsYMnmTd3BjLt7J6GV
fp9XyStAbMuITt+lDNAVMUIZ2ZcpaE4goHmuEWrKRPcP7d8JtHxiiq9FG7UNabbF
`protect END_PROTECTED
