`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hPWjtt7hElpq2OKbN4/0O+ThJT1uLUzNYl6gs4m/5/XF/J8K1RZfg7KuJNRanzy/
eSkqzco13cI6zDujIHcORfCyyt8k4Zc9H59D74qiJVwJhJxZtNFWXVfbq+qT8bbT
otBnaBIhQ+D3o6lN7pxABq/pYYGd+OlwASHFXEvRmkKZnWY8r0UhmQCM6KH8Qe5Y
TQ/wjn2mw79XxI/0tXkg8FP4Qkg+ptsYYkpAY7kW/uk860zv2tn5089NUXeT3OG6
zVZWefYeXWLUsU1+Z7uA69eIu85JZXiEdOpag3orjHZk/nRMKZqiaPa/ret1lI6l
2XXrwFfnjAEE1d2MKvi94C6Mnk8NnCFDEK7gA0G0cWUKWFGyYXtskTR1Bas2e9DH
5ToIRdE3O6QM6uztTxqWa8sT5yZ9XTxOxkwxmC+q+Cge3zD6qyv7Pby9wZJr0n4s
dvybYBQdDP2z2/0aChERWb5uefnYG1UHSB6vmzcmeLK4VGo53Ya1/tq/TYU7XP0a
0SwaTW7d8vsehvrxXx+kScwhrr9ZHb5SPXyv0+D9WbdIcOC1Wqa4UujXHHDH69Bw
LC+uSJnNvptW1OF8TZJhCNImQf6/gfxEWIKkUZORXBXfmpH9HMxqpLToLBV7YGGB
HqX2OpB4VaiA5x/01snxJW5jvngbaLs/OlEWvNau6578TANygrkzNXg5PeWT7ulV
LwkAAdZYS7zrzeEOiwYOc949IDUnYBWOD1wLWaDXAIP1oQg6ZnvdP7L2FSmEIdPX
LJ1ZkBtd9+KOnAsZ0RTMg2rr6ErSIw7sftnP4AuVSYAXk4OfJP0Y1hcz+wQSW60u
IKw1wXemQUyPzJPaX0cuhzYcHRO4VJ1dsjnP+klXZHaRIQLZGhCkMWgbIAUgmvBG
26TTdROEDSX+tgaRrXjLt/U7DwF38Vw/EuTaRbDWEkpnDr44IafD7GvW/bu7CsgJ
m24Gw2FtQyKAJRx1xvjP1Ory5YM4wj5oxd4ScQUDwlc5uF0ZLBsfcZOb9alPlCP3
7NHmns+KSUCJt5Pg8VfIXqNpM0pOYgkS6NvM48YdILeNlDjsSL+iZ5YliVio+NTs
SUcxm0UPL4UYnXtH0wnrY1wTSEdb5aA+VzFieZxL8x49apHXZb1NE4jQjebFrymX
+vHu3Ko+YY/P4rFaa9vkuGLTn3h3uWeojibpHpvcOYUKujKcoyC1cj5uRmN86wxq
MB1V9fkcD9pfZmZpho+DIej08q+YUYKbbB31y3KH146uZsymhkEPShd1Wyp7o4EM
rINYuxFfML5MLW7Tmvc71fMYJtPtXeKkuqfzxHqao0mD5ivWR/fvGrpsg1raxHof
YDZ3BTB9mTLTSJwOBInG/yvObiNZwxM4vtBd8r+OhomgJzNodPywXyeQp9PZ4Qkd
43oJacKc9Ch48fqI01rmQ3me97esLY9JYkjE+VTwL2q8TomZO/zmCsmESOnhqzgV
lypPjqzfRDMQ00n9/LvjNDFX/1bXVdAWluNP63vGPUnGT8L2iTxQ1aIU1IBleHnd
CetyN+vKiuQzT9d36yrlhtDJvLX15mvFrVBYUszayzdhVi46qbqPS0/SaQLMVJx6
TwBxYVfiJ4FUcxY9Hicli6dQA0hYUVYvng64eg35+u7xhHauUx/65yvQ4VABy7nx
JDiNonm4gmPKFWFStKVQMdcl70X+OJT6eLfguKs6h4cRaPJVihTXGrkDJUO/T1tB
e7/F9ZrsnEfCze69QX3S5L7+S+qI8b/lwUbTmbeIt2V/Kylh6nzLm8Y1RPaE60Sg
xpiTTPdUrCqr1uipqI8NwDHQPK8RpjgsfZjc5vaKH6rEloTyjWUKtC2ceMBGwUO9
mxaSg94woTn5eA3zw0wGVlQwNYfdirc+rZjg/6LmBELwEqBHIccBQCCwfuy3a3JG
CyalbAh5sRSe9u2ftz4+iN4Y/UxmYUGhZAzcsRot1cr6dCpSBppS1UeYTdDwKACb
MD0Vg7CYX3gROfE+p+cs8KfL6VVKN90iujbwJUd+Lb7513pntxOt8Epfi6/NjAA0
bkPfRgPNl0nLgb/uadrf030G7Jky2N0k+JiRTZC7xt5TC3QywEKzDySRrMYkJzgq
mzyRpcgqx8LQdgEKYsMLvB0thNN/AuhdiEZWWBu1LHsiuYDQ1Lb/ys0RL1SPhwCt
zo35Fu8QAMFAy8NWxgYSrTIKPCys9hPOw1sA0p18ViF6vvoAoXMF0dPFXWe50Tj7
I7bdmBCXrsHiGnxoIhreK/5cvRhK8NYfQmyySHtD9me333pG6MqS46+dRpEYnWMW
+qNqnVf6F3g5o6kOPfiUOdj/G5vpB5LazBsoWK9/zvbIYqJpcPSD9AkBrrt9yFIs
nQl1EbmKD7mJxZv6nvP6lZOGmtJoor4jSUFStGee22syRwInTbWbC0Wi0NfW+Dod
TbredMc568uIgueRXLuvKMMPH85CBdBIpJhFnKwZYQ239LTfGfhcW0Jn3rtWVeD/
pGCSRZbSokVHHzjqEWnGPoyj7NUB+1GCtXHn/C7SeMVv5DX7KCGxeFlh0E5J48PD
alvLmqfcoKInep2+r8Id9F2LTUxCc3dovYlJ3xssgrB0BbS2U0A9Cu0TuYuU/Cud
Occee8hosz9bi7++4my6Wrce9IRQOKbkLqrxoJ8oA+TrwA5V7agypTS2j9uO+NRY
efevvpEjwZqEr2PqhEP8yCD8ycW513+67aphg8ksnCoFUH1mIdB4bgAcknQHjcxo
tODJQy7Cx/Z3Dt9EwZzndwOayd6/HZGHtl1oYGNDGGGxMAKYZDBpR/G62qlCF59r
l1nk1Cnxjb9yOf1nyXcmSbUWBs4ZDk81CH9TbFvSt5wwWKqhHPHCaQsIA4/6W937
0Hm+YfyTQCJWDUcY7VYebQDQex/yjmKUuParepSIl87Pn18QGuqqK8AS2XGd1BCR
KpUtpDb3oIvlncGeDp0EerkiWiyDRRcN66ZXiRQD41VDUnCti12UQWypfi75GwBD
xiUSuj5Z35nCfnD8BbWOU436gB0tz1Ypo8el9LaBSIGwZPGBNxoIdcXJtOIUCkZ1
LVOFXSB7JWhWFAIMzDiGZH0hOs0Z3YkSCOwoh+jRkxUEGhWjJCUdvOoWUNZb+6wV
trVUMkKsBMU1NvrdW3m9EgIoCF9SQrbuwX6KXil/I6frcE43aTms2z10zf4xIjEf
Ok9SuUOf3/f0L3AMQKW7LZ2Y5PYz3UHoww1CDnvXssYgIkaLE05zelBmZKB+oR/L
Zr9feRhMIiNXuxbN74w7ZqmEaMv+e+eM0yGHNYsCnl1iURtONGdJhOCNU/CC8PZC
CDiOFDL5H0NQ5AOeDRPWL/OsPCaPDmC6xHKoo3uIraS9V0NKovlX4Dn0wTI3FuKs
KjDY6rjKNurWZsBqGzUc1HIInE78BX3Umgwr3OZ+PVeODY1m3QE2V6X1qAk35/O6
aZpnkwqC8EoAx1VYYVwvk44FoEzzpIdvTUtJ+PDzXlElONRQD59HUnL1n7S4bldp
sv2Z/XZ+1jTjLCUZGlsQ8vyu4fHW7s5sRsUqZ8HcSOg27p6naORR7wgC4NxzBN8M
FTu8CmyUwbx9BO8dIjiJy+KoHs55izpP11WUUYpvYjX1XEAMVFJD2wOtGspSzGhY
BL0HjxpjRLl+haAS/vSbtDgY1PGYlQnDewCyFCfUm9LazgXntGiP6/schwkgBdRT
yABjb2mBnl2/UZfZsvihoepJ4uWA97oG7YzZxui0Fz3XvYowjpaZkFu5iX43/ARU
dc8cErf3CaFH4svKhWo0NsvElcR6E0ZzOF9z1vs40adjFBgkqyYtwrHn2lLMN9pH
H2bKHwSGKYeUO9RstzuG5Q9nHFlb9TkAf+9n9LJqjvIoVkg4FTwzncVXYAIfZdYb
AZTe1Bkr8rhulsQlsKBtwKWOPMLGM0wimDwumVqxP+xAzhtnYOnASYtEKwEtUhLE
eJPAv9gVpucB1J6WNu3Hxb4fij/45k3WuCqUBLrb1t9da6BWZz3YEqvCXxB73WOd
WlERpapg296FFMEATNP+H8y/b6E3hSOQI6o4kdQFZni8SGIWT/OHyOPnRN5CkZGD
4N+wj+Qi/KSoJ6gFiqVfwsNUSsD7Npq1UOhH184egbhID4FGa1or1pXbZla4KgzG
9/AnSfoXty5Xe+NIpdqj1t4aAC30fajY0yUcdRS2dFVGi1OncJXySpJcfJwb4aQq
DAkKYhaMVeCFkwZ24LydDAZCueI9fIHUlhzbmg9PWo/cocVozUme4vvHWjYM3AX7
MQbWpmVd1ArfSsgV2zPBO5+liCL8+rwxVr2KH8LRA91p7pOCaJ2xkotd+OvY5hL+
Ld5mVLVgxLm5+eXDfcswXQ9fXg1sBGgVVbSFgVSR0l9EFfyXCKmPcJnLSYqvSaC8
nKTW2H1wED2JVEAyOhCypaLfepJckqUmB7ifORinqLbT6moRoEqsTobZk+BUeu30
bpUp715t7vF+se13zmVAo6CTeJ2yVvZXz6d2NHCnK5lvwmXIyiC+fm1qWLmLJGcN
akGcmGIyJ0QhM2v1iQPckFzIlrEzkzp0rPH1QdcTlv2gw71+xHHYe0cvnduYDnR5
ro5XWjDvQEMbFImOWuSsQbggEVE1zi76GDb7Ej+I7wEHCV4mjthN8tVTzbz3Wj/Z
5Zwf9khe4AnJ3f0zkPG2Sm+KSnx3D9SS8TWIeVsIxsG0sx0FoIRNYgxJnMw+KugV
KRxWiI4/joe9T/QjQL9578Vy9kwNMwYMf8h2QHZZUYDfKUxgZJQhSpghVaokmf4A
Zig3MvjpD/SbhRe51g8wliYSyc23ksW7NQAr6tOyEfJUxa2Gfzw6t5lyB1wZ/Bgs
wF2J8psvJ6Zi+acKUngO4XFR+QuLvK1vRzNnCCy8e0LHTf6fTCXVVoQk7wlQHwMI
8LRNYhyLFHN3xl+FlIUY2DHmsluOjFZOozbLjUjd65inGFCrFDjnz54TzULXBzK/
0x63bbe5Ok9Kh7Q3BpRIM/lEutg3Ui3fS2fTgfZMW2jmJfjUtu0NtzvE+rIou/ZD
XpO+C1D4WqlT+WMXPWIQORHxSiaXLRtqQgV6+LwBaY34gPMmRqvTcyQWITCt/t0g
7V1VRT2mv6flfO05SU8BR5p4dSMnZ/GFkQo51AsoxO/pxe3S+qQsoyCZQLB9FO6O
qtV/sy0DY7cg36nuIhGOGeY93FC3Dgc3GPQOdijKEOvN9K8GkJUAifeYnH08x3go
t/U9fMAviooPMz/dL7m68cZdyl4Impw8aGSdf4hCxXfEtOIo7ZhGCETWbH/OEefJ
fOIflgiKWHgGDUW4ve8hxL5sVR/KPWleCbZJTj/xKfWiugDod5bFfp+UsRgvpVEZ
Sd2tWvoTJsG2IWibHdbQIxgz5amFCheU4djojUeAAo62Wq/vo78MQ52SUT4GBFlJ
`protect END_PROTECTED
