`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sp3cr90lCReFsgEcQWUdCNenmK0DZuPZ1P5njlMkp93NFf3ZFIn/eH9WJl8xQEsd
M7pJnCS/EsQWajrw6BGx1cb9ZFcpSJFqPDtygs7CnNnRtpXoX7VW+F3x3f3CcJF8
9uPxPqu5GnaXg0t4dMG2UvDei//01ZtsiSSO6hqI3HOa5todW1GRmOfuWffa1oRV
AvSpr7LeWwugNstu6pvaA4QGG0S5C0+HCyuaKPbQ8A85QT4m8Usl0g0HWaGRbl14
W6ocaHp9SGqvMNlzTW9THQC00MAwz3x1Hwsbiai2lE95hi8FZ9zIMyY1kM82hTj+
e4Fr4GMwhRnA32pstmIQJP6zROc9sG0hCvynHhMIV77uNL1dVQwAAmoamGa7zqeK
FQcobMIUp0nfC2yYwIwjoR1QvtYOCxO/T6vwoNvrUQcpYJqtfSDjfLGoSLRPS3O1
bHD+iWxJkbL6XELPDk1OEUjhWqD45e3as5j7LoPyRwzwSJJsdoFQ7zw+AEctApzk
Ei9aPEk6vV9LUxqo7keCqioNI9iy/woxRIVxtVLQW5EEBkrP77eiTxBQYH6dHYcs
TFszbG7SjoOcqp2s4NJbwZKzT5THfXfqkGT1K7fLZGJLF3RvOnDhLJX5AMQ7AFBz
FShbF24z+Y3FjU82Uh2EBg==
`protect END_PROTECTED
