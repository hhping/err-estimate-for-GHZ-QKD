`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpFm7ewkSJBIhaTRi4CdLWXyu344HJDvrwcawmhUDlpEQP5aZg40ygT5v+L7inTM
8ytHMXMWOcDCuINeRVFotoJuyD2Ac6zCXJ4Hqkbf4Q9wcE/atVbQTdWxWz7AvwIe
QnfDsh+xGzIvav+D1GZ7CHUbYVp32VWnEFoF2doneUY=
`protect END_PROTECTED
