`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FtPRbzhoqXejfFinWRbeLAa8JqazTBoLUL0yy4rWoUdiIW96mFTpMom7rjVX7sZr
gqi7TgAhqEKgsWwZQILvc6jRjn5gDCfATUqHDjWxUTP7QQuqqelehQxWamVRB/x5
9WCb4maDTb6icaGgGmh2H4BvIRSoUykBxRUWVyLuau9TNSO9xDQ6vBiP6bq1vVzO
ZqFTMHCzB5Ghl9J+j5/slmMgpNwFPEXRwYPMHFXGiL0ilsFaW4kfE294JmVWVQ7+
xnsph34zkgQvFpQ91AhrzhYCXNKHqD+vTcJR0UdC0n+zuYZjmIHP4Re9nLe+p2x3
RdkF0Wh8haYu/Bs7BiIPB86H9+n9zsh2ScnnTzEWiUYMgJjNmzDMKMXxJBBolGZi
NW6QrtojFzJrzYijLO7l/Y6OXLhdDDICrnsnrD/ofwV7s2BeXoYjP36RuldDM6+o
/mrb2HqBkWkE9dg1C3p49WP/tsovnc7mkBngbaRyJHZFRNgHVA/eHP+B4zZ+GbYa
f+KlCG/szM1E8P0Oe3ms85oI2nFUhzmB/YJD6xHo0K7TwtXZ1upN0rgLiT0JXBni
Fjmbwp8R4y/b7uBDDmm3xSeLaR8dRlobJNq73CddcBMUa/Ud7T4cNTd7oWJA1IY2
QGh9JB26KDUhpelXCVU+93Ikd0uXm/2DCLO94iwVUoVWOYk0X3LsIBmwl1xUbzVE
g2HeImAcdIQMwtV4JrhYMNN/caT/x/S3haFhSjc8A05GQUyzjYYOWSemIEj5eQ6a
k0iICxJeKOihcagBKkgty5qK/rLy9ugSwCTBmajTSXDXBB5VhKrB1H4C8fIkd0Io
2KFjpLW5uNeF+M/RsUtoFBgAmwm85qQxuQu3rjC33Rjp9OF11nSNhl38cgRWDENq
T/DIRY6LxJSScNWmrxsqrnsGC9xnnCVNoFl5KFUMfXQTbxT6VjqVybyRAtPjLxlp
aJ8/ZA/urvkE8BZpY4o4OVy+6PA/CALgaUv2rksDYaSxqAUOI/i77z9IlMoO/0/f
tpQJQo692rzcGmft11g2NdBNMrgwb4EUmJID/upDwOft/uiptHksV46+7GEed4ur
sVIRGpOsNWXRFCpWAYBSU8OoFaMf/XgzhkBrW43qfUlFWVrfqrsq3APEnD9qEgct
8XWnh+LqqWdRPrx8mYbgLA+Nvt4VIb2zVNt57zamxTfZ7QMuF+g3yegIVrcjTWLn
+zWw9ZSAcOFeBJAbanDh7REySrFjIWR6+D5goBh8kBV57XkIkDGHL6VPeVLlcPqD
Jyi51N8FQiiopQP/XUMnGJXghH0nnK7Yj+1t36B9GH405F17FBHSty7mpoMb6BUm
9rXcClyrKWmSbyCgoDvcNoyczmEqxsLkM9JV8RRm6t1GiJFsLaJoYttuo5QRrUxb
zifLQHkLK9TSiaEFpYnuitZxFW9RZRylUoEGFjKViYW5hP3MF0AEs33f9B08tqiF
Kxfsz4pS+mKJkMF3wrgLEb37BkoptRGKNEcYX4vtUXS5kuMR+hA835Y3C0DcV0em
0yDSH8SJJokiJhRfa9YZT/TrxSALhtisTqOFI7jBEc9vSqz6JeJ2iCDiJ4G2STfD
7eTM/bxio8cRDzlqSm0Oiaxd7h8F/0VSvlKNr2crAd0fNRr6UzFSyhdTT8xwN75r
zM9tyHp/FdSH8yJKrfJnG8Gq1sIIealXlm+UfQYkpzkgipwyETCuh16ZQSHRr/oa
wJXRFFBtAawe7VUGyFZcrULLECLjNQSdLd3mpOGTBtMx5oGDfI14vnrjnkjv2bll
XGuIhla5o4i8Sb7uPjklyMv/WHukHHjtYR5XFCZ3FQ1PfDqf4lHCYco2FaSS8keW
1pnMajJEGyGAx7mNPxy33LJgmPxO4ku+ULFzqsCG/1I7hu7EC0JoePOxjNcM42wl
9bpNvmng57ESiZTgTvYUYKckTMC3eAIYaAeeMgXWM5KrwP3qprkAcDRv15IrVR27
2EKa0uncLpzhp3DC+gicct3HjK3WIjrs5e5DlWozCeqeDhmI4SCWaXOsHjsWqn4w
bnth3nkuRw+BLnkP782bfNbN7YR8TuSH93mEqeKMd/5gg+cQ6LVt4ugoo/VgWz+m
1lZEkd7BvWsXmNKGjcsXj07rE7vmS1p3JAZu6v8O+DUHE1fBTNFQv4xAYKeazDLw
0q8aKXM6z4TEhSPWQvOCKBe96br6eUuMpBSppwQIcHF0WHmqT3zF67V6uQzP2uVF
fYDPYXimGNlG2MJVd3qIcxl2kvXCHYrOeDSJjJXAWMGRU9OZgR2AWZZc38EJ0HlI
6TtjplyQrF3kGrJlQy7qR2AdjbFyNhciVrsR97b9R46TN4WU30+p7mjLL6pZw6MS
MMrve4SJ1qIF8XD/W9Cit4hn5J7Cy6onGL/hLae3yfsgV3Gh3VQRVXWYawWJ0SMy
CFLknDXR6y4uH6BFP6y0aLsPxl8uqicU1Ra5TowSAlodoBYpXQ+uUlxlou2Sv67z
Qfpm49SUnSFVlbuB6JthqTzlkMoIktrWoO7aeesgIHCu3/kWPgUL4QSYtKQohhxO
AOThxS7nJPBoIcqEE1gAQVjNlswgLczHc81MoxawfFoi6zUsW8XX/CfTrzGvb+O6
a0Y3aK//Lkla0WL8CcxkPPq0Bvj/yK2g+05omTURSPSvEPFiRLwNU6BWmVcAippe
9GHEoplr3YnDXCZ88fkmI+dWl67AQkGPDO8H7uDojptkP9RQ0i/xm9ePmuz0neYW
iN7Uz6vdHX/EsAhpH/m38t8Hnn2XVCQTRtlgjjoDWF0Q2f25V1gQyOgX0QuaSQu3
7Qosez8Mv3kQ39AdKaNx6bkBnlo3GCgtVuYxSxAfFOFpjXa6qdi2EH0R0iqzAUMO
kQDWeaai6jZfqnPgUqA1gV7rn0I6Cmo12lZlyia1CpG4NEA2hRtaKexqTBoaSjtd
yPVy7jpDqAOOGABrI35MLMrnqgCPZSHqrDlsTdyXb0szNzErlnaKGFHm2MBrzqWA
7q+1To9sCszL3bRt1jjThF1WqdszWVx39FHAm9w+9akrdeYRWAvrHe38X0Gjj821
7Nu9tYDW2OE0m1l5Q7pzQlN4gtql8UnDfFcHzzkqjrHH69ZLwCiCMEyOO1pXV4Ct
ctXGS2XaZ0Z8+AKtGCgfQciZchPwapcvRVjHzpp6lcIqrThV2jcqq2PC5rzYGLHY
NZHQLbfgE1z2f5a+E/nPlAXZwAcqYjU0FDLkvPQah/aPirRvfMNqizevIriyvyNP
bZqGA8q13257rSJjxzi3i+BodQl9lmKUGsWwwSNzWOuAk0EKd9POFEsdDN1zCeMo
2Un7pbsF0RM9KHbzyAspljXv+dfj53uvrjJoUQcx+Y30c5I/48jBLfrj3Gz1AcW2
029EW0jkBvvEucki0ouCUfngOeN79nISWM4ywUgM7R3YVhqQ30zxY2EL2uGzMTcB
gMccSjWQdonyoBapLmZo/LdyiQd3o2N3JxxXR3MDFYgaW0yfr6JEB86Q5HhalQRR
bQvDyowEQSFB0rZSoBURODXF/bbUXcrRieQ4emiI2FzshFacRF/ArT5ZrdzVm7Vm
I21BNYreR9+7SJ88rOLkwBhSY8QxHGiESSYyR1yNtSpKLPAcT42bhzn7u3yxTXP0
s8phUtHW+zEd0J1Qq/wo1OS7cmrMOsCV7APSA9dZAeBDvlkeCTkJI28RzKUkdaXQ
RDOkAiLSlPToGYreI0HK/WxJwg+KqsM3F+LAb6wiDYKS1LEEFDvS/TW0TwZGeyNE
yiU8P6zLBWowdZhXaYyc5iqmwLv1EOThHgJhQ4z2p+g8H8H3vy6S4GmAnuMa45gG
/938p/q90SLjH15tRj3U3I10HuY62SVDQSN6eil/Dg/jCHODsp2RbBvHL+PYb+iF
CkqDaToktrcFNKHRHK68hgz+j+5KjY3oa1pSsl4ooO5gU13BPQWUqjcf537tDUbF
la68jTai81ZAPnRc67JryCRD3ZkAIwZ6GhO9MQhx78ZQpxhCJSme43wLfCs5cTuo
Ka9junIQr5SO3p3FPPyEBa4VnneVA/etfgnIssyOzNl2YFjtiXER03OWI3ocEJLJ
kIAtLovRmimWQ9MMgCOKYy4ZfKrYk08hinldvbrFzuJ3QKqA0Z85aOeXf06FYCH9
pVRIozRwhwDGMR0Fen4NYp1bcaxaAs4BMXKgD3MQ9G4i8t04qhwbuPe4gFdP2oke
yl4XWy4x+rOC6FQpCJ29tiXzS04+LHblHfOxuKrgAgliUJtBpFFND1MjGseqWdaW
MJL/B0o0w8djXvkH6MbB1fzfKtJfpG8IEgdT1Y0A5KXsS+v5eutIAafUABoa8U/9
czmV/AT4sAC3PWIkEHe+kWEMGIs9CdADRKFZOoJuXctv06qC06E3MRVd35yA+7V4
zzfOqbDVOEL3yg2ssEefGHXb0EgB9KRDf4p/aK9MueqiwAq05GmXbEPBOJMXpZzq
wysgMbaH4d3NUAyHTEzTIX/bBV/xg8Dx63bW0cjGHAES0FCBBMhD0D1kM1QJUayW
Z90BzNppSd4Fp3rTaPW4mEfSSQY7IfzuP5KBCcgFimay0CBIpN6cQQePbWJsAZOm
3infTH0Z7z6T+BDLk+TERg0A/vQhVlNbs4AxfmFI8osHMzM/dLwBmwg+4NcdpnLO
OoD+SdrzIaHVrxHud7Rp/4fHqoVOdFlUzSPv4FDKGCmpFU2xtIgWNNgRHSbatVvk
4PyziYOXS0Kcj/ZhCJ/YT66y65yLIGu5M/PzmNwt2WrO834JNfTYsZtRambLIovC
7n3Fyzt8Ptr8ZLC2LcXQnRwFAekdULZP32XEcsbke7RE23ZLXcueq+NTy/jfDz62
W+AWrIpEBu9raUPMG58DS4oxqEDCanUDkTbGsOmmou0xFOxMnfqk169zI/N3sdsD
ggUFR75SY2ykZSVI4AypZw262XwGQZOsxHkiwzYbDQqtGTQjRpFz5YYfqn9/DQDN
m4ZdaR7AmMwnJViWddGFhyqQE/p0kObhJcz6gKtyxNhl6C4iG2VcCM50iY4bqAQA
V8XPM2GdwqrLz0B8Fmc5SSRDDxCWLj0/75rVDXxKiPUx6wN8iJlq9Jp6Hc8cskW/
DkaBKtrIoT//wfO226RH0pBjOl1uCzjBt1mRydLFXKIIuFx0Yxa8LBWnU/aS8FBA
O3RDEXR+fRjsI2gXhIRj+KxdZNhin77+XtCQRqO9MyouJ/xTuZjHxmHTci5bwU5z
STEEVxzUihVuh8Uv6BXN8Zmkt6IT3auoqNy3lUu6UhklB46bF+pKfl+0J84Fc8Ct
H7K0jumsQ8xGHe65vFxYCYFrEQC0Uqfxug7GQzRorOHFNUY3tr/qDMvRIL9cjniu
kegRT9YZlOfRuIcAF6zoBG8a6R+BkS0SHeFKiVyT8WFhV7iSqpUJq2RKRLaK/NX6
vflxPBFN9QVxg07/9MKXjhIsqLIgwefvwW1HuA1PCTtt+/vQroH3GcB5W3LdtAtK
wMOsckrnBvg61nX5rCIaoP/xrI0ykXIc5X4TKYFWB+7S1hle6XwyW8ZJ7Ztn/zRn
XrPczHJawEsji4olPRgKgleKYr0bQv0KXXSjeGGtmSvCIBQWICUBcFF3jLPHktib
f0ggOkYgKSRLCI6yxHYIQWvocDmdRCFpgXriYosQNXaBO8nFW9F7iYG5zUbSPtAH
0POY4+cbdQgkEtVlvc5bPiokTFzBYbVSSypW4emwcW47JDGueHHstP+jUjMdzcW6
gRt+6CLNWY3+IoK0tCSvKUP1ex+xUaz/vQjhfYO+SkfmZRJ7Tksk0WdpuOzCQGuh
2qWPyuCkC5pQQfeCbIz0z+pUn91nMrPpMcKzG1chBDWjo0cIhjX5NCk6FLl+Xl3Y
IaCsmnW8G9zVduI6L9poYsa0BzKhR6kmMAw+jHuIM4/5PSJ0H2/kvIbkOGFFRko7
xIJSWSSbh8MopIsmrfiXTpNzrVnBCyasDvMkEZ7zQDTVYSUCG5d1RLq+eHbqsHGq
qGLiYGJqWxlNsec/f+vLOd7gIpNNyDjxrv9elTFsywxiIx2NixJB2owC1xLwpXK4
7bcAR62Yd3V8PVZ5Qxfze0cqZrEfSpCx8i+LjvGL+qRuhkeDf2OFTZPPM528D4BE
TgmoE1v+Pv4d5PKlx10bPrnzRsUlRgdNBNX+VFPA0tJXItTxZmef640Kdk6Y+yi5
gPZQiRkLVOrgaWgxgDNRZn2lV3KGcbAiz8jmEQHmUnPwA3OsOKBy2CjGPw7vQx15
zHpKmsPJelSw23f6SFxRTa2fRm4tno/ZMgtrH6xc384=
`protect END_PROTECTED
