`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8b+yxaju+oaj4fzzAWBTQ5VwKKO1SeGTR1TrkeEkHonZCU25yAEV2xq5CqB/RbK
sFp851+Boi8gKzFMKRg5FLbIrwYFe+lOwkQB9DbOsMBQVoQCLHwoa4OQu50H3i/7
K09aleXM6wRnEAfxjU7oFVb6kX4vVzu78+YvEIE/xyTbfTL5GO/4FaqQOT+sXqC/
rGNd61n/bcc18VsihxmWKOZrJRT1YVVmazmBd8gjDXlIAsPUHOUrPnZNw+5nR4S3
jRKei35nhRZSG8LeM77wpe6EDxCiV0Y4NbjAneQ7n/3yjLsdlbuq7Xh9dPYh4qZf
dowYyb+cZEJeMQp1YUUP7VIAq+xx3mk43wY0nD7e/rMHeO8oMuzhWRlpNPnK0KTe
oxBzr7ApjsCNPIEU3ebEsxUtuVcsiTVSKhq1wdSA2FIQf3BbyzEvHADNY1TQibRZ
IksldCR6x7fXX7liaVW3SEiANTxCdAKrkzP13sj1rQ2McG/7AGyQhycw2O98UZAv
MOpHVxdDcGy+BurLRXmtCaU3cncOxLoSjZPXmYm8wiVx2Q4AvSAfwFk1DqS6BGqs
17wHF46J+r4dofaRLQt5T1WrGS4jx4vTYG4owFz3Roqsqgattlf8DdTFNU+o9NAp
nwcukb9xlYnuQ6eLX2YDHVdpaswUEKbXSUHmySGHWsVs77+pfz7Gb0h2ntvSVjzd
dXFGAa/AyIyGqvbmdtUlQKdSdQ4d2qR4Y0K5WTGO+MwAgdNIrZTUkEdrcI6KMqnL
V0NhzJsBQBTdeudSCMC2p8yxsFtRauTe/MBBsE+c5c+qCqdPiA32K8AaZ1WGGyXA
9dMzLl5c1FUbdkp+PW7Rm1ElfjX7vN3Tr8LAwzaMIDHyyaLddB4m2cucEpVMGZHu
RhKRWlVO09/7sYTSTnadyEFnAQdqJV7kIaPBX2dBQYfbL5ZK+2qFTcyxa2GfCjVH
f8vnIT6dE1DqJjcVpS/w0ux6abHI3z1F4l7UrNwuMMexGanj6eM95KhF9vM3IvCn
w56icjCzNSN53+dfaXsxrNY6nJJk5uNpvLmY3RmVIhuGxevRbUTrePtQTwJrLeBk
iehMAphuM3MoWcEXjN8mEKsk3x/5+hbIHQs1ECStjOvA9+bzq5yjEsPnmdaJrG3R
b3D5HEmHZCghOPcN/SmfL1/FDl/b2eErYiYUyR3y1iYqRdj9662FPBoCS5MoJQKW
W7gpgs9mT13ppwPBmtigDTY320cMWnDy/VBEWdz0jYahgZv7mu88pOeA2np2YfrU
PafqyB+/ahC1Z9rWncji9JWNPgt2f3X3zsoAQLi+PlRiPvssxYzdWAmJvVMDOxHc
1ewBxAuP3F7rxktC/EkP4Gg1WJV03uRigJxAkFSrDYSKCwJbq2eG40RCeBKjFU7o
1zshZ+W5fY+aWGVGwYXFbhyraOK7MFV4CbsiO8EqHjd2bLIUdCR+QMvcurjqOXh4
/0GBc3wZsoD4sDGgcumzc4iauabV4fIjJECEYrUJu+15YZrTobPz4Af4wW3isXlm
F/Onz1lTdWMLyJeVaVZD1Hxx2Lr9ClkNQuki6WuJQ0tSriMQX4bpnCmseMW08g1x
LI7tL415nKKuqlkNt5huc+QgUC1aLiafH6wYkpXHFDTADBKflCgyBWc3qY4IyDtI
W05ZaUB7IhrRnAsV4+FEKbozDfCEZCHjFoslW/v3knv4MAn3J2BPSeYjxM80hSA+
hnZBmObYp+Pewi8zi7UIpq/zkFPU53WWLaLIAvKoU5aswMt+hJuRP5ZkOPumnMBd
N0dns41HhTPyG1QMkk+4lX2Ywb2qMh4SndLcgVEG0R/J8SkOEWDW5TPycadrw7BY
sxfJb+Iat2tO1qC1Z8kcH7RXXCB1CVh8CaJMivhLf3P9q5JMROpF7D48j7d5LhcL
sqCldxMSpOl37A6EsP/qt2n2Jwh5BX0zKp11InEOfRoCzpcAke7LW7c3YMe1niXK
n5hnS0Dyxt6WVgnk8cThGUk4R6t/d2vrd9vN6E/vTJZQYtEtJ6ftyHbqmm4KvquV
2H9V1KfaHaREdLf+yrAOvVxn64cR7i1XSIN7KgtOEjzwqklwy43o5FDM4UuIPCbx
Cca0q1bLKDY4YXZfGFW8l53eagf2XFs+ZYerPGiY5CsUC4QpBeLAxX/alJK8U7St
/JZEJyC6WLhVDc1qS0ebbTULD2P15J1VFLTnkLOzUwUglzDHysDWmMYxY8hdRUbG
jrhR9LmcM9JSh2wKjwyRgxPuzBqjMH1xzd+jhpIaSpVJ+qLH2CB5rfy2Acp1byyP
nFh/O4wdLFs0JkPM5x57fQRcn0UyxMOoNpq6088dud1OuEncfVbLStjPoutLOQ54
gX5v33JEdbDHt0AdYMpn6hLVBe0xJD49Z+86IwB/kJjrCb9JxaMWqCOE9/TLlnFC
EmMEyaSIJcqlhhlk4KtJi6SCKy13QbBKgM3bRSCpT8txr2S/ruC3kMfHh/dzRPyt
3ooeqgs6nncBxt1rvQZWT/onpwNcZicrROzvjEIoPeOC+QMQEnPm7JXHSnRePrCU
3Yw7W9K7o+NzdePAyojxTemyw3SS7q2h6uskO+LrG2aYISbwFkr+pBFc5rGYR/yj
KMSzU2g34yCgxv6kfaWb07R7/QuL3AmJy8mJ7nbrjWkRsShDwEPyeBnJwf8wmlvV
PFYauKZLFS8LfXgESjSz60XpW0qDfSDXhk9U1i2vvrZzfc7CHuptUK3a7mx4cael
mMxoPbBMyrH2+Er5/8lX8VwKXVTpYt5k2dZvm8Q+mwkfXbN71Ed9szNltq7nkIyC
+VpyXXwStVnC3IbkPim85h6KKkA09xfVOM9hAaxdmG2/jNlV8lZ66IGtVJVq3I39
FDHAlEw8C1AWYexhVfOy1A0skNA07eqM/4dcrVun35bBHxakluXj0DN0vImYF1o3
pybXjB76cLpRPG05pw5RkcRoojhAEGuXXPh/L5DZjsn8JKfjrr+ul+2/Y6TS0Mml
hQW58gm+6C2nA7JuCdrElIF2ESW5vgNu+P4V0If7DowrtGDO57bicJiIoH/W+2gX
1bTau2WtI+qqMudLaytewYzMV2zOBeNqMyh8kVJD39iTRaWVkL/LvdkzILvnPxbd
g8FPYGh/o1p+Y3GbXGnLcZSkhTleEt2QRTpbZm5RXge3+Gzu2FPf2ZCI7Uxi+Hi+
AtksuFBGTTJVGjQ9f4SbOSDrIzUpgPnw+75wUNtNk8SYn3BnCymzUeWqR0Sl5H9d
IYPTgqnVe31HpkK01lFad5ql3Y9pADlrQjS7N1zRvlOuyqT+/x4Si3YVL4d4bo/2
unXkHNzO9dcwtPMHBzuch8FH+d7IiwQ41hTQuNbEjXRG9R2ToCdhagEGRq1Vz7Xg
xXjPDe9+YWSTajo89XaOFSPY+3IOF+DLJPfyKCwl6St8fPUxi6tYrgVn2w4PzIDr
FqUEl5IxcgE9DOdRC4mxAZB0x+eSRG+UyKKHafXCF2wI1tTUVqhUabFMlXQOZSKp
QMqF+05q6nf1Vj7CfRCJZLK87Yu9O785xvZihShzWg4WGU6ErE4tUXDrtqcw5oW2
2oBtz/t7Y+Nu7LCBEIWe3vJ8uG3+y270YEqA1XZzMVIGilnAcmTJuGNcL3lZnAGb
`protect END_PROTECTED
