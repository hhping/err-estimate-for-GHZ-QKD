`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rz/8fl4BAVQCcf8U0gi0AeqIOuvpaJ1YTdw4d2EXgqvF1Uhz3jhw5VhViqupouL/
XtGDfmBGDPb9xQ3xGYKyviudhJHCLVovdPssGYLGA1EY9uTWI2o5CQ9iL43dNGbL
88YBNDfz/1eEmPMUnOLldEsi5oACg3h1gsG/+TNF7cJ1i+fMHUh+vUnkO4w8C9ah
g+hEgwWqnOEvC7JS6dWgjXajQb9uuZKYkIOgT4DHSgFPMt3tBLwZlM5kUJnet+xa
G++AcyMKHOtnmCgvtvwSUFqUAxZyifV99gL6ZfoXM00cK1HDNqPEul+2RHrNLd/W
UZOyPCEuXwFe3v+tS3IUW52j0fSJFlp6Cn+LHcZsgPfIHC827TTKFxDatxKnXLkH
9TPoJ0K3R/Q+Mk23lUUN4zBY90CaEpsP5G/DBbyS2WgS6lJrPNoK+G8xH7W4e9ed
lc5oZUnJ2n7anUCJ88FdU7wloVv8QNoVbV4rhNw7pIJO4liQ4XPr1FerREY0NMXt
7g8Akdv2DaCecpyVtxRxH/8VPOufkMgYJPtGO8qYFwMrjnz6FDZf1hF9d+gdUZpm
9MuT3fhOyQJPmnAAlQjOhutlPAKq3jOUo9mLyMR0MBnO50eXZnl7tQW5CuF1yIuJ
cu7MpgEGTlA6rZIRAjOvZT3SsOz1sgFgD3oYe0LFnTzCDAXlcTyfWhwCWatr1jlU
P1kr6iE1iawaSWPRmN2n1iuFoQQ0vPOtBF2gPBK7ZGeyRP8S04GYwR5tDxaV+Q5W
cAoWOVe+H5qHh/Bvm6dyGPL+W3cX34ZxnFe9qlIjAfgA4FHaYIYtPwVpbO1b5n2a
npCWQOAbw5+a/bRFo7Q8Sy3N7FkBvHtgFQVjdvQK+yJe8patquEG0gpxIsPL292U
bRlqXv7IWAoFbhbI7Hzp9/htcRRkd9gAXNmWFR1QcKeE6aWVVPJSg+H98055DdUL
xoj8H6Iczj6n5eQebWcOezjNGumFmqPfBoOZ28hVLh2ttWFxwDjgW8u3WB2HCP7S
qfHyAV9x4lhxqERuePGZ2XLrPYuyTJlfSb/xyiv76gU54amdFlsZQVI6yc4/kWXH
zyWnIINnWoQawuEJjbQEt3GVpQi2fgtyJWDqGCaTVwJdedgqhIjFjEp1n+mh2YEg
qFno9S+6m4luUpcbp1RE8Yt24u68H7IAXjjlvXyxirmXWa/3APe2p0i9RsIC26jF
sgd5Awf0fZR/Ow5iq6g4jALauOybddyIFULGkotuukwPCluEa7IfBCwStMncmtMg
KQKSAQFoQ3Oq1CDQORUpSfSezpt/HZzIkoQALJywWWo=
`protect END_PROTECTED
