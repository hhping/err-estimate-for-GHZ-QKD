`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+m7bWYz83JdbJdCG3nZbdAzkfPVM2VUjTUJmTHOFFXJa0XYXR/ObfzLwq219vkD6
2AEPJImrHTiHbz5CMluCZiOJpXZ9ongEgnmA6Apeu32KDM3ceNBLKPX9ciDIy6S7
lOhbVKmz58psxwiwiZP6dxqesarU0Mu23L43IWLOc0b09G00wqG90P5BVT61eBvv
UnYTgB9PA2RLkUBSSkfNefpeOZ+itCvgwW+HrGXatkj+Gr22vJ/+HkdyjDX/Y2K7
u4tj/RdNIVHOlIJqnuQzAXneXtRaKvtM4KByKTM0jj/AbIfvsL1Lgp69KqhfVDn7
iyXKXPn80Bt80j0ihpYdfr8SizoitOCj94SiGTFd1aTqq1MHG0mPlylZhF8aCaTv
PvlMXlXGnSP1HlEUi0oHftGGTVX/Xv15sVaLC0aOSvVgij1BxFuN7vkVg3+46CIK
Z4Nl9c5Ob/+g78FsCgi/XesosrJfQ9cJuq9NG1qbQKCxQBWjdprembGZf27oIGeh
gZgD1k3p+vR9Nyt3d8uynAWFmg0bl9dwfQHzNJjpDj2XGNLnVzIsXB/ep/OofHnL
2UK+nowNOQUqDsHBfXqcjFoSjeBHvv60Ia26HrpGCzP47zpP/Tht3MG94eqLBReX
SP2n8nmprEwIbtkUSsqC2Y1BhY/3STERE+wAK2Taof799TcJ2tSJYJPw+VvCebBy
XOjbQF7XFxmPMsZ/d9YTavBcP43DuwI2JY8tHAGVEMpk982HLPBbxrD/XSIl7tup
Lg3UpeE8ZPBPqrT3bHQpDXcSTiuy5qVzrg8q4FUUYRPy8Y0PzBbuNFo9Ld1Y6u+a
JWLCGjjKJM02Yh6lN7Uv3wljaeDXFVZ+KaFf/RaTAUoZ7kpsXvsfvo4gTTOchWZY
QrPnswd2b95YDRrrwUJbeuNm5A+qjjXAX2m8FsBae2KGqr+mbiab1TJvzyyNXP3c
cqvnJKTOTK5MgZJ5tBtlAn0uQASYVIv5UqoQYm7nQOvbtHHFJbvzvNPtLgdBvSW2
JbgTV+RakKoLlvx5qV/DFRTU8LD6sQ0Kqqmjcsgo308=
`protect END_PROTECTED
