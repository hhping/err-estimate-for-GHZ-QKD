`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiaOpcZW49TS0ix5OZEusNxe7EZnHPFE5QEL5qikSBgwZs/0tC3ru5xJuxPkfXgU
Di4XrUXQ78pApQxXyNtvC9a1N+IuHDI6/1QXwQ7jckKnICKropxD3bCTRV58FXbF
cWN+ru9q8jLAheI7uUgFlNDK6AQJJSDsGjs0o99b+0Nawaf0LQTIBGLdhEgetnGJ
TV/dhhUg+3xfqRVAU5xi0FjNitDLDbOHb6d6dJvK8vsRRGUhj73vPVHo7HfF7w9W
+q8+wwmLwx8vnSMEMZ2Ce0nM53d3YHDLdP2+lSGm2HbFnIIUkMTodEctzy1kVrvl
2PUjtzDr3wHvkdD05vXwaBa76dPx0CsqYW8quWrmZPxL47NkEWRhxlAh/05AC4V7
OkYmWTveswjhkDn0JzfKhG8cDwDox8LVBm5UObK13hYvFEAIWzlWNzfNG38aFXEG
kcjawChcXXR4OSnRb2BiMSDX8b2bC5eHCxQRruQV8rG/poPvLVy5LzCUdsuPfOTo
webXbWQqb3a/emXfgHxsjSKR/9JOsTLNf8OMGuQhlA/zaeQ9D75dg5xZgdfWYEm2
WcS7AcDOCoc83AxzPC/96KXJYZeiGRmVlgzcHD4ksQ+SQDCZ64SH/soAwkGWr8HF
5vu35FWlO+/MSido29jlvHU2svtPMlJGK6P+GJwEvNKiNPGywftR7QpvjhRpjWCJ
HfsUcvtQmYtYMa7oKMDlbqErWVV+lWkeZnmntdrmp3Ju671Sn5wJcaBa4IffocaM
`protect END_PROTECTED
