`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sK0l0iAHxskcsAKWz8k2Q6P/sKR4tZ7MTzD+A4mn+Qn0C3Ddd0NLabgw3r6iZJ/y
kCYA2TB8038FAZIIw4tL9onSmXcn+AyHqB0+iyP506Qj4Je2Cr0aDxttI09UKo/2
4zLWUpMb3yzWdARtIZNiOq8mVhC3L1p1PfmzVp84PXh/Ox3MdrsUkvVWklzwUB/n
dGkspgX7XeE8+w8GM/yBjQR+B1Lo7Q1K6HIGDPPwmG22Nz+mSQSL2JzCsmZWKrv5
o7qdSLzVI6XiS1l33BX/5yxd/pQlnhhmpO9xS/0wcWJsP32ahB7hTeCAhZzKtf/Q
OwTnJkce75wby2lzPK1SeDLTpamqwO6BMnBA8X1fCLtMuoDR61OtGTilvnQFsC5w
fFuoueyiXhkc/nPIb6ONm8CPBTFwrJ7uVEjvG2f69UWbdiG0JHIF4e1Ip0k0bzCS
eJA1KVaLRn3ISMoO3yIEDhtt5kyVtwLM1mr0Rz5PvYeN7XSrWEeSKFvFmcPjtr1y
ldSjMSzPh0JmXSc8v1WIbalevdEXz4V3KHdcj5dM2tIM3euwdsMiermkF5ezIfyY
ryWgX4QAIeEFOjV4KKOdpOMmsQ9E1umSlKzuJeTx8J5AnhSgrGh8qYJ5CcqvP1fn
AvksKdjmKU4DWvnCYqPkNlk16LwlkNehJhyg6FBtbRccYca+kE6DdtgCCBO1b/61
sDMIxp4RolVNnVNf6Z57AOtypsABLzlEU4qhzW3hQtG7nX1jeyjk7n//OVUy1oWm
9pyUWJ2KtTjJ/s5tqbtBsJhwCCPRhEH8rNcpNCSn8EAy+weoKtmzXevN15seAewe
aK4C9OMbGtmONqu7a00klBaCFANlrJNBHomPObdqBJFYX/taXPz80aMDYQ8kSjXs
Awh7lVNcPqIOA6/XF/kwXIg6Tj9EfMbV5oJPY8ePUMt1+fO2fIBViPPtSbrSQ2cI
yzjqZksLO0fj4PzonMlcbf/dMqu61HOd/ELSmgGbCHhomeRqB//A4Yq8LJdXtiRo
f2oM2JpoVzFHhEB8tjJn4y0J4AsCToYvngzWJXiaKchSpnWYQ+3WZu+7aAlGxFl2
9oMURiwk8iDToYMFdlNrNQ==
`protect END_PROTECTED
