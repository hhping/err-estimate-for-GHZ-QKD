`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EG89kctXzt4KSuPWBRx8d1oRsjGjJJeczBnb3OQci0Cx2ow0UV1kDeIJWECsuh+
h/PPHThfbSS9uOvb0ng/9PgZ6xhI+8N1Juf55C7tLQ4NvBd7v8hHNJ1H13h/ClIJ
ouhnOagRqo9ubPHCx0NxLJwVD8E7dunysNd3Ik3e6xAgWNEzwD0jQrh31jXtfJcH
BgQw8RyGnWejN5oMO1mify5tL2O3NaQXFREkgDKzDqbSmArKn6gLyHM9j9mN0NPO
6/Xi6yTrGkEKScUOkcRPlyu16Bk/HovZQs1fHwID7vmcsdF2FcbCNc76LLHfYOoN
o1jY5xw4iEppgO/sUWZ+JvZxlWey5q/qD1OtkVMweBkHJitNyYhYWM8dLUz9D3Us
e42lHUgbw0gSbjtG9ICJrIji/FRKPk3MDqQps87CZ6e5y3gdRMmhxN6RVQyV4LHu
5gDL924+iv/rz4pNcNwojkrDJc5oJRfvooLCNASAQNDxWOwAhq3UGVBs7YsMT9K5
XoRdRku+98AEeyZFwP0kKHLeLZBteEkL2SJhZh29b2MkUBGHEGxgEuB5C4tP2ota
4j9thbPLQQfSoOsKJPiBxuWfI4JU7DCgYjXVbCXPfRCFajZnXQPwodW0ZNrGdPa9
MAoaaJbrHGODOWXIIeAc9LGA9zVgcc+SrV1x4gJX9OK5U2UftS1SdZaK1kek49yy
VnSfKx7oQjcizxuzmxH+ZsFnuD/7wU7swsPgyTodj0tjpUAPHNVzZFvNs1Dz9S94
4eMdSFDKHJ1AMFPT8ZLmNMnqwXUiqVoje/vukbJQVtY2QUb5K5aVBdFg+dlpXXg5
`protect END_PROTECTED
