`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErvgBf+CrygT87mZRVk0BE6Nfgi7kPL+mvuuCVDfSZoyA8HHuCvZe2UHwcKhP2Oe
QII1Wz46ShQtvVOdtRYkMDHTUd+UMG2aFlEuvO35ndcQ5ekGUPiMsyOeiwXxu0ym
IP7DQngjt9VMBHK9uVWbWlc5eHJyK2FaRC8r3GCwyarrWc07vjekmTRRZRgUnDF9
gmsSuv+PWV/ypo1E02srR8G+u5TVNoEI+5raxG4sap1NekBPqK1qL1dLX47J2NxZ
vmEta4R9nbSJcBbm7h/+mbgozIGNHHKW4ykAQseVDl5TyAYybNtKrExc1aAsNxG3
Ewi27DzZYAazqwnCipUBz0JysZAwJswFcSjj2EXXjCcRo7pzfYFBoHZaIqQaGDCS
Qh8UfWOPxz2m3VAqm6OiyoF+atiArE0xrnHaqXB9OtjidLSxIvXlfbTmPP1K9Tci
DWSBzHwOn1dz+T3YtyBriBGEgR4sIX6rbl6B+zgCOiPAsEeq2odbJ4jnSztHvUJ2
N+jAeDTgPZEVEDTo58UAwVZ6rcZU8EfRjRx5I5w/AR4Ln4SYnbrURoHHoIVXrJoj
mOxne2mVfk+8pierz8pFO3cP+UM91iCMYPuh4QkNxonylLFC5hZteD8kmdy4Q33X
Y/Hh+UgsdL3owLee6R6x6kHa2pbFH1x2oietxZO3qnaR3T9/jDDI0ZKU24aAN28+
Y+kWns8t4kKNtwwH/YJ/+B7McEfUWIPu+JK1Sz0OtRBNe8IuDnb3tDh0YwwgFVo3
clJjJWKE6BiYB2Qz9AGh/4/j13PTYU63di16ZFjRI8QqIgHdtFFSiZFgLJdtoQ5z
uYIGU6epO4MgzMdyixyLrd99nzxcYnVIc7gHCCuvOWs/HD0N2gCAQLXQ8py+SqUq
napSoslmeQ3G0bpxentMqMYJPX7nB0Inmy4FLZ+U6J4oTJo6Ud9M/+NHIpTuYEYE
k1TJ1JD7orkZkMD9T6TUV0MiJ6LYEOD4vyiX7bx2M9h2jxMrfExeQhK8yOx2MMLp
QDNLd4iYEIdgSAg3eEG4rFt9/lSGGljXmaTyab8MVPyqXWrhpSkJtnO/b8TZoMc4
36jnXej/jOAUL2pEmaDE/K90hmNga6T7x6CqhkpwkIun8LYYUtbxurTE26ZKsYsp
zHzQ54AsaTNtxo5YBEYSUSu5pJ7HOI6ObFW3rrjPtz6PDoCLkR5E/+JFLu0CWIZ8
s9AvU/ywex1kKsrCXChccuoKE7uTYcObFX7A0GcEbEm1qDvINIpVO5GfS/l/v2qo
qHqUH+fzBhYqSd6K8JylCNYuEOf4AogmerBW9bp4yvwkd/l/2QsT4/sTtC56zDwe
bI4HL3/89vvTqmC1+VKJEV88sDP0gmdb65n1HeajRfW+LvVWt4/sZaPyDPJnRWtG
02YlKX91ieNrLGyf3qp1UeUJZkf2sG2BLXmjn5mKSI5PG5pfnINX+/TBluMua56C
p6WZtldD/NmWhJ7qCSeIwABzx06tB2B7BER6UbQxqOxHJwEauQ23R2i3PBjkoHDQ
ZKXAbsPAQB/kNy3hyZrCv7rsSvfO2tooeKMrswZRhUxQTIr83XiOhadaRMsYzLIS
tUazUzekaP2C1WEfPumHS7EJDRKs+DEJWBVXECe4M6FQaQ1hMd8XKnB7fu2FXZEg
n2SmKChkrmCqwGkO89SJoVqOYEt6NdcKPM+HKUeMcwH6DdHZEO6Gc1UxnohFR2Rb
KJMbFQdcDZsZEMZj5P6CqMQr+MSAbO3lUepzi7cuE/o=
`protect END_PROTECTED
