`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T2I1N0YPXOlG/OMqeUQ/nIn6xWk/MYDqY3ZTVJZXN9fiVPyYxcTJQc9YWUrD4on5
DvOh+ooRo36f2+doAHsmBDIxbpgYsYMWs99xuHs9BgFzA6TJb90zJAKscJrT72kH
i69y7YEXPbCBYxdqBtt3/hxO8Ep6nJqTTNMNpYZofB8zOWFeHFqGEOMAlcxk6kjS
08cE/V2HfhXHBPHbOAxnSyVcJVKG4x6kQEahFTQ3U0Xg2nTZN8sjHh4by31bhqAL
Tr5i4X/lCOblawn9s250P3r2Aq0gbQpnkAn5fOFTvR5nty1IL4FLZONKXQlEuP6d
46angXqvRYZ55dlZGhOxFOB1sZoMQI/16SnrJ0Vmoy6oJTWDvEqKF+acZvtTic7u
SfKVNsg765mOSzroV51tlfy6aeThMgOvQKJIC9hsP4s=
`protect END_PROTECTED
