`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VxtMnzkgydV5ns5PqMyOPAFB1PYFM58AY6SREBdOAWmkWt6SD+sUBKDulAaHdEn
zPCYuTjYwabB/STc5aHBMEULlYy3+TLdiJFEXPuuC/qPTSwxJfa81no/0fQKer9f
apyR8bTliUWCIJGXmrr7Cq4Q5QR4oBgX2sg0KDrl7OF66937ho3egr2ZJ1bs+ezJ
4LnGSs+5RArefDE+vtJGmlNJlvL/f7DEwq2l+rmi+iWcBKMS9SlqHHbxGTpy9C/L
JwXXTgmwHs3N+ZApGfdb2IiAOgiqHNiY6PdAZ8EQ7FWXD+i8FD0vtdl/iP+Nk2+N
s/oqEAuIBHGVSZNlU6zxj9KnaQcSVXdmFKa8YuLRFJeajTGfuaswrccOB40t9V0N
LO7KG9//W+UP3m7Keg5dfX9KLovxlxVtjjwX3o9DKEXjjRq3tPmlN6U41SgVSasZ
R/ruuGntCxm9L0HVhPCeVXDENwcg9EGmE898d7d3b9Drf+VlegqGwSje6WwZMo8D
MIZViWEiIeM/Q+Yyr1nB4Al1VQNQP+ml0rMzBGxEW+a9fjV6i8KBs4CV7G8eZmc4
4EVqU47rORS7NIfEiM/Or+8j6s/33xKif3rpq0dtoX8Jz4iNmL/AHFb9ybPMPXu9
1151ECInrV1HBaO6QK5hoCP2xEuJxqcK5uSWk7N+nYYZBTBPN27AXcdsFelV4ykE
GotxXFljT7dGatQEkmPR04lIAJyEWmB5+Yo5nbgIQdGqJVtrT8MR6jw1xBu7mVvb
5pIBkRKtV0bpxrgJjVu+Nyt4vvLt/MWhetJYlAkv8cx+tB/wFB77UaWHLaofbhmp
BOMBUSCPwdXPZwS9Y9TbLGoYpkublDA6YSOz5cAN/ZE9KEgLgnYDqTyefNBrkV49
MeFgrFH5h5A6nW2ebwsALTexMvPQp+OlOrVwGho44WN4kYdirTq6x80NXREQKViP
mGfRH/EMCo8d/XHJUIjEnBhP1lJvLtZ0mXnN1wDVfpX7SC1rmryAWCttpz3cVwZu
pP6PihPvjCj8/E0hRwgP5Lt8I2V9j4o+Tnx4bhZYSQY44V2ow0Q2LpmGj9ynd19/
oepyZd2USSRaIti57xMS8SrV6fysSCTqOWbUahPUXlRxW6Gzqw+IiNgiJTs6az1Y
A0NM5aX4wKMnmOQX3dgGhUmVwSex3j/+bWRXAyUioiyhkIj8E5au94di2dT07pmd
g/qaYQaMy0UEFUbaEonUpNJfMoELBaeCkT0Z2HM2SuBolQl2wXI5EiLOz17qUGYb
Lv0+6XPksZXiYU2i7drnazuJAbWOmSX/bhkCnKyapvtXQnbjn1BRUQ7QF0AZXCKZ
jnjcZeHUICcDP4JLiwalZn0IzSjJmOO9EPf6z7XW9PJpLhKiu45e0cj1qtEyT0+b
2maofW+f4KZvTKSd5/ycdu0O83lQtrtXNeiuzC0e+w1G/hSOJapjed92zQnzSuCW
BNH0bMr1pV0LUIEHefbxSQTgZd+2srK47DTLISx098S+9WPrZyVyCkLAxVJDtAYB
KW4+FDk65gisaRjqfKYpQ+sLtXzQksW5XUzuCxAomxnYgSBJoWXyPMFmqUmudQId
RcyceSKoG22wdvEPMkyAN1MwIY8U6tPaa0qC0Ig/4Z/wJ6LA2xhMZE/KMSVkUPPb
x3v9D537C7ubCVa4x0tV2JAiD0+8wZgpCt2FjI4lGMx2b7Ryguynf7gGxT7PIdmg
stfia77+owuu2Rnlg1BtLYMCPpD2L9Eqkmbo5ieg8XPicvsR+jfmrIMQ2C11/Z5N
wGogkS+jfXYPWFJqofFlk3XOHYqIjhRtFSED0Ygg5SIjLVmrii5skk10G2/rbvHY
4GfKbquJ0dI0Ce2rU2oKqpOJwi+J8g3SdWOOdvgdSw8XxWbO9Ti4vEE5wV4Rqxn4
ZO5MHJFXA9eJ/vNvNW3ehv2muWxkKQIB2d/qYiWsdE/Gwpzfb0sQOLZVYu08PXBS
fcXNuw//DPivKACXQP+8b7QbymJKTtTQc9iaYtst3MEKxGVxfetsUNu0jzWMIfcq
z76cmDGpfxUYN6e74GhHp0vLFgZ93QIvF43XZWvqNbabiIY9lQAGOVciYUWvxreF
0UNZis0FN3LspMlD18vscPfGAEViUiebKwMZFTqFmKLkWy10qW4RGMD8qARBlpVI
1dDfPg0RIyhWU3LpvfsqWA==
`protect END_PROTECTED
