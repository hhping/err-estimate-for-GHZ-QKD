`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wz+eDJmbm9kjcMjusxn5KaxP8ZT5XDQY3XpUeJP6eOJGaY3fgm+W8djDM50RX20y
tf7oHd+N+SoaQWpw4az0JOhNiVzXhSB96IU6W8weqt0KkzuaKwDpLTQJHansUFZK
c+k98sGJ/lbfBoB2fHaiFkEL2YLi1RpegPIZMPC0CKDehLgFQ1R8lV3mCUOUmOMx
OFKQq9ibjdK20yOZVnmzOAolmU5S9RLLz6sAuQO/fYNxFuEzdkyKGu8XLriZaVfP
rKN7tQtah70rUpTb3d73jaxUWt0PEop0jFXkko/yoK9LlBPj7cNXmAEgG2kqaG+D
NjwaJtbCFzrQlYy72scAc6Eb9z9fVPyQCWFugJfyoTi47lyfP/yC3pnB2DWMeSFd
mPTNW+DXPbM+AwwQ4AD4mnJee4gRb7pSUT4E6r/dzmMEVMipneqpSDfbL1ZR17PC
qZ+8hwiQ5pvzvijUVsKzcBE92VUVGs+wBGS+7RhjeydPKCIQjxoYjgI1+C2hWyE+
VzC3VjtobQv4ccQuuB16RySkXri+k+6cNwrn6cSCYrjjPYPbbpGgTJZInUJyTVzW
ol+VcYx+RZ0dqsQ4mplx62Uule6gJyE45atFY0mRxzTpWRT/mrTYYctZ99jy8EFg
v7+ZJG02DzBt59/Mb3HBbT9xCcaDMEbTjLITKDczeMDKtQOrR92tlpC6aTGrRUbJ
EX9RWUX+CM0jNf2HPKHAMuJc/OYJ2y8HtVI1+mDU7y3hYurxs+c29LpFwvjAXvmo
GE0++nOa7tZaVQzAqORyxq7ovH7lBlvD5KOtvERuTJJm+QibSsiJ5Oa4oCdsQIee
wc+zQew/qjajocdw0QPFlHohH7VwBxT1n0z+4Fldnit5BAUEfop9TyLQEiQCNxsW
qVZWamaV4RtxBCBSaXotJKn0LRTApUYpvo7LgL77rW7wPek5eVImuZOYhZ5lkgjO
3w3Lo7o8qzNhxLQIDC2tn+GDZ356cBu+NeuVS0jgqn7GBmmaqJOzG2gacvhTW9iK
palPUKa+lZzk2ZfRaj0DzYCL7YTkJMzwmLcIMJNS48YLGXcyzrY2cJ/onQFXJUle
fjykFnTixO9tlTyJhNDjdl6mx0qlJP/plTqbzGmXDfCRrPAJ57KPUq2xgIXJsD0I
4wBF0IUCEX1DzOmquJ5mzgFuaqLQCJZUA5sp3DrCqxyu++CCe+EJd1IgWRHVW5oo
6BbvJN9SZS2WDHQtZ25ZqynVtCTl83WzGRtzmYLp0qRbfBtrVtzEzAWCk9WMQkQo
XpIyMdzgNgI85YMnOjKxReObMwYQOBPrABdnDWLdreFhDU99VRBQsJ0ivf1kWmx1
2gBQ3yUXseEVO8uwtelI3HGB2GFXMefJ1BFmjt1CUaF9DuKEuCqffR/RHPIkfQjR
SuZplU5CqzhlLVp9ZE2V2lwKWrMyftpH1DZLDVd+EvwET0ogf5XFSyKlyDmWTPUb
UJqENAceHvv8VwvctDS5c7dQ7UiqWK+Fcwx5IojknY84UXYoChuGHl0klwsLYKC9
FzchMiu9GuLB/2s3fN4xqf+vnCEBgR844iO/MmGOTTz/RrAq9WYSDWG1Se7XHjhm
ABV7x1BkOYb8nYVi+BDpgDNCtcoKHag3eJJPWxPHt1+hn0GfnHrSgXL7CajX9UrR
grBiaYcMWUb5Dzfp0vpL3/40O+K+Fn3jWrILqpXn6Kqb4ytvzYK/S9HMhW4O7cdC
pxmgHwlsFs+i6VbwWI+FOTrhmIsNKbDfMjzmHRVFqYRCssrF4JfFngrwgDRHR+Fs
xftLT7p5V58JuSjJP9UofQK8P9qGgoobN3Dsx9Fda4kmkJeNzFtNix5hyFpIHICv
ilSYxMNrPxwc3iEYx7/ruUcH2CA+ZNBsWxBQ0SEtOnz0VfGmGxF0dbJxrDBStmub
3hTTefTDtirS19cFcg7aHYi+1VKFfMAi90QUd6kr5VEh5jp34PtJt/zwKjONAg2v
Tkm16mtbwoa6j/AVEqoNtuCz/oZBfxSm3zRAJYf638KydvOjEl97BLMOuT9QFU0w
aWmdqaSdJ6Q2CyatNEjOaUEyli9TjvOlVOIrOHnSHxg+Gpb2ZW6LZZLfh1CvXiPF
hmzaZr7P+MVf9Xvp3bp4tIRmRzairV0pH2W6dd1kNO4jn61SNT77p2aYtQ5YU678
SHiu22gla/e5mdwMYk1bc3ESXyayBhb75gii/gEJkvibbYDC2NfEhqFdxSqwQx8O
eYEX59IsBS4LVvyeN+rx3a43iVFQAGkvutm/7aPfSUCb2UpWu51Yr5mZpeU8OPev
TGHBLSt/PXKLauhC/Mig9BAPBX0USISJw0RU+sjUTUwTJTwAhSqNyY8FqmnNR0jH
Bl8RKslQmuohnTWUmtjdDmwddaggh2/gmVLJgCzhzQm0dv2Grc068qUk0xMPAJGL
PLx5xICdHV8zqKdOqVxhdjQS4W/HjUY3PUoMhGDoiYogRZRG03KLVLmhPwYKxZf7
aNJ2kwGsQZKTBERs9KDytISdCbYeMe67mPIf/WNW37VF3aF2kyS4YM21GrVId2Qm
F8tdmLj/eLNrnVi/mAm5E+EvHrM4ajVcKkjWU6fLGteVmVyBvY6WUh3BHCM0Qa/J
a91QTymLLekSShgAN74rJbKhg+2hjcp9P3xTGnq8Tzmas1Urk5Xo7bQuaum6Bh9L
U8n16KHXGrnuiRRgPT8g2VXhlKMFqrxIGOJX6WUWXfmW2ouyDHE/BAUowYlCcPyD
mtsp3yn+gtHPGkUA3IrqlZH5khlsfK6EqWbHsPlyqEM28hAC4WmsdsMUFATwodHI
1BGpmvVriPXe/Wj87a6DvU4Tr0BtP0Z6yfamT9+YpIcvJsIOKLuWNAD/0ZGQ3GJG
ReI/k1u2H5c0LBwzg1Z6zf4IVhGBYoJLy8roYaGkTmXGFxY18rIjZ1wj1tzrCA31
+LtdzbB76ONi7ORlVYDPPArwXF1TOlfDfMD/cG4X0NCXM3t/YTV36tqTzeGf3jkx
qYOay+gUttW4m/FGS4efNRNuTDmN+t4Ur9KzZKZZPqUZuI2ellEt4zsWN75m3U3e
89gZXfMDWgzvoB06Fjm001kgNuX7TO/xYtuoNbnDt68xVnlVSGAtDEjYXw3V3Nxm
HAeso2AMA+4p7R1avn+tzaZEpeW1G/ydr52T3tSJz9d7fNYNqn6ZRV8U0j50d9Y4
IywPy9YP+H3JY2Hljty6hLwufZpHsBZrmjIoTXRS0G+dkrQn452K6CMoGJV9mMgf
34PmnmQZ+Zs6jxpOi9b40rq8tZ1U/4D2V8OMDYHqhknclGWcr/vIq5+XBr5J63Un
Hwy+kwjdWudRlA8hL3G/VUUYAqSspuM2biNHyaGOcTurq3tUpYJYN8k03hWjn0Ap
NcUWctokltsRrLEZ6EoXibHLVzg1+AeAm8+Zgk3rWiM5ocoC+eTPY2JBEBjKgRDj
R4CCrE6g1hGZ5jTcfB8W/fL3ru/jGqErdMb4RABLNwgMW1F7R7SMt5o+E8hIK0sG
DMvcj3Fi6sJQ9QmeLGQpA+XxNDWrKAQt2SfYoLDpgepZ5j/kjmZab0pf/YBgKJXc
3S0EGmR1bJrG1lQW+2eqrwdbJPZJHTCUz192UraW+3PfI6WrVUn76NJv76NoizIe
/+tbG22ZhQT3T6AabREmYBmzDZ285+6l7oa41XxEU8mo8MsTOpyToTm5VZ+HT2P6
FT7wEUtvhn01te1qVsLeOGZUZ9+/2jucTZXB0z24fRMPQaKvGQQWsx3zabChnYUx
zxHEAWD0hU+wlMa1Ap39Peq58G8UFlzhoxjFRjMpU0AXZylip98KAR0oV9yIKOE7
Y6uP9PWYffU/1/0EomXzgz9ufa84Xzr3ceyo8i9jsZ58NO9lkHP1CB6UdNDpdIj0
gmSlInlKVnotrK/sm/8byBFxJuBmd9CHEpy1kVS7wds9F2dUde/Qa9cGHkdhfEHv
buDVZaCE0dNZn1jKVd60lC0FcuidSk4g/GADXDgKZ0V8HTHfmy18oApg2ZAs36So
717xpZFZBPEaiCdPl1S8Kq8eOAInXQjouiuq+sRk6VePD4vpUQ4VW7fcjJAU234T
irtNBJimf4Qdf6VV2uzMYmh9W5O+2c4VEdO+nM91H6akHR7SFk9wDKpp5YOCwmk9
ABzXEYLlsvrXSPckPk6CzbNZvJaIkHxYHp+5eLsNss6FVQO6MQTPUF753c5yWX6G
pbwSuh2ksbK+FQjWjJse3vSCpklhPTOD413E6micVJYZGcAYQF10effyKmHF4ZP3
oVXuP+qpXdUgpXNBnAvSf3k064qcsld5LykTo6QWvIqD8BunOjkivnAEdFgZ4KTV
zR9/YF4ehZ3KZmyse0WLIVccW+H6OVmG1m130szGuYYWvMs6g1Y7TJ5MUHFZ9I2/
liHcfBIIeuFJxvJaXbBy7sGbEt+6O1p2DSZagpLjjZQfQ00uQkOsqPwzJOwzhdu+
Q7Pj0jOTQlteTuNlGDzsSXY+/sXwvm/eB/FfxitH6WyOtTtmA2k0rai8q0+21ReC
6ZjT98+FORQWgGuSXIepTMttO+pK00P3FLimxmOKy1v7vTg46dg+Q4sb5m17KVVb
XozhpSSGznmkVzgdnX5+qOtx+2WCQvMTq9RafGWMxK8PR1we/YGlYJvO8ZPO4hqK
viWjFjLH/t4KH7gbf2J2+T0oubpOBtpOTSM0sGhnBxhy3sc27G4ZTInd57TIhR2R
f3PnJ9f3rUWTp1OzdrpCjHSsExLe0dCf8p2SMM7HOD4QE81hDtzeWcQi0/O1CiR4
IQYfURJCGRwe04KSblJ6dcK5YwbXfQcav6uZlfWS/WtAvNFh40G7n9yrqr/zZ5p2
y9x+5NaiwXXQ2jRflvVT8jHUTD6AnByQ6rhoaf+w1HYYjSmQciMXx2JEQ2nlNotu
96n8KzQ/BHa9bqzRb+IFpZy0bkYk0PX/s0vBDI7qY2iDYcaCd9vd/Na7onx3dX5y
Rs/UGXwleva8aWBSqxDMfMH6F2SeNx5cnMyHTim+HzXG4AUT/bjB2XD/v8GmMAfG
wcCkLY/OGbSjnQf/qX4WtUu7SHEXamF8slvc0n6GyB5YOxDOBpLKSDVmfhaTdFtP
R2bVfItUcne5L3OENuBd1PTvP6Z8JQvTAGzUIoXGw6eQ8cQRtK1RtqsB3FTNnDF0
Do6s5hBTRHEo1KLAWBp3BjGX8Om+oT2A915xA3OnT8LOllBiLQhdxsneTNqVuy2s
MVZbFFWzo1VjPVs51E5WrSiwIyuNFlW2Jr9jlGo0kcEjRzdQIHobf8fYwaKblx+b
49WIwIlgQCE96GG3tJUFiLlpJzhykYOEOW5neD5G+AHK53KCowFVYwxCODZacTCm
YQ9TtZ41/BcFIYk9H71OiH8TBZ4iIqMD5KQ9VYWa3hqj6auWKDfSuSTsq8CIYBjk
5Aq/NfmidELjerXGBhTvwRqkR2GLcParUIpOLYeBfxRwF6A0USFMH4LzUhzvJofA
K8qRwuk09wUVlvVIjKQlyEKSjC+6AOOaqSmgvJlLR6fq7bBOAzbjvvILjUYgFLXh
5BqWDNx2seMSYazt2DQ2W3wE9sm30ubtbN0pnoGzYs67tt7g5l0OdVJgnM7acZbk
xWgi94838q/p5fqjDmaGGvCxu7l1I1upw8YZx0/aEZDRjxYobWph5pCTZqGfLdyz
XaUOZQAxlBvT4k4Cv0jWjKbb9qYFBwRqsWnsDIHsaBxNpHZ6VmvGaPe3whWZnFCD
XcoJWq4hyaMr/s1mcQi+eQSNs2qN7jAhvA5j5SP03iB1/tSd5SVMmTvdPn7ZWTjD
Ssw227dwBrhxSA8t/IUQ/KVhoA3hhIf1tDh2NaCxeWJB6TNbrbxam51EdTDwGRko
y5E6lvWRd0mT0tQl92c/Viu2tEmkf6ajNV3wo6jGoqQOSAqUf1IzXyes4bmen9I5
b7R3i33dUPNeytnwWHXyCwiZNGqiQb5xEWiQejOAJ/Vb6Pp1BBxq/ukim2VKZ2GP
C7HXMB5HjHHJ8DeRXMYqytLJ+Jb/Qc/c5mDACUNwOIGsyNk0UUnG5ZOq4QiNc0oS
Bv4VYNr7OmOaVPtMgT8fAVkmcA/U5yTF77o4/fw3DsT3c6bMvMtQ69ed8xgUBNoi
+m4l8obytYW2iUS/B7Hdqj4t+CEcD47xz7lpBKG9+QuYrrIWCMPmr4cvo17szCQF
D62sGbFfBBAgi3HRJv8qudKbiV0GZeqUYjtUDz2zBJhiRpuy4l3mJ+OBrjYsfXrc
k+2z2WkRG43BikKnvCRsqj54B1Yoo7+frnNkAZqw43H8f9pKezqvRC+eY1zQ0vbq
z6inASVRt3HN/cbdS/8/RltdQBKTZ6pG49IX/5LUvNUf2Ayz2ql3HNBaH9XPLpmL
pb5CSqA/N98I7a/FUSJlGHcZ16JjB3WG0BqDDPFtoledA9Lomjx8x5x1eLhAgvTZ
jDMPlBNbVN9RvO5S1U+EN0o1uYPiojMLgnyV//N5gICOlWb+FJxafsJew78EhtPK
24RUUBq+v0RHfCfQ5344LA0d9wTcJfjuIdjaApECsQm8XEratRGgenzhRm93WoZ4
ckztEYVAIxTH+jCYjEWpYzkqKQS2q2hKPuM436Ymm/mefKL6vyRrDJHDoCCyhpnn
LWiiMToRfraSqrwSdUqs5m2kWly8LhiKz1CmN9xOqZWjvwlLicopSax1+fKi4ihJ
DoocQYQFecrMy9AOxmrdqjUhWBWue9mfTV0Jpi6/AEz834QHQAF54/Z+diYZi+do
J0qwZjCURvymJepw+vQFrSkxalOUkx72ZDphDiJFVZ6Ayd6IBkjgZKDC4lBUodvZ
o0W6mey0ia6W4FI6DfOHhZVFAjRHX63Azu568N4xQK/rFGk8TQvqViGaWX31g8Na
NR9WJ60AhY2vM5nHgtjWcBd4qXocLvZO0dj5/RwR0UNCrznXqL1LLn03gTDqCPoJ
t72TxGDhgvRUKbq6aZVPd/tL6iqbYj3R7yeRdZn3xpglTzBvQpNDPp84FPSB2TEy
mfF43eW+KGvErxcZlkykx+ZG8m9t/gVr3Buwb7Dd31LWkGhCE8xgO8ZlO1Dd4vBQ
8UEum9ZEw4X5ipgCoM+Yrtv4SsPGpb/X8AJOPJzmm0R+Ut0gIRIy38PfvSZcLmum
ojwbNiJ94DAjnP/eUTganLGCotEWuGx3K/Gvb0puMGgp8FRJY3np1LUCjQmhSPK0
qAQmrO+WI+BuyEwJ716Fg5B7GBFrJiDPG1w01P3hV37x9cMiLbEyWXqwuv+lWs5t
Y30Av222DTGByB17IgSBgCyrnu6s/0WAHLuJzBMq5vnnltPxMQgdS7JDJREwVvfz
4wGAOUrfYYM1SNz9D3nw4Qkvf1ioul4G8eh0O5gHPZ7EjLT0ycrO31+JVj3w69jx
qsIpyNGxUUnACLW0r2+7eXwwR6sf9Q0nbpkXUpEbolzAtfMEV66ZyIStFFP5Psn4
YRUk5EA8B7w6hxA/7G+DUt6yWrbpj/zrQMmJQarJZXNboUcMqrm/VazXeXAS6o6W
6ycqME1x/QH6sdA8+Qv32WoSbbPpy4aAJPlu+gFVTF4qshlcTCSF7Zb5wvlbdmUE
tC54ZQJReDAwQIwdKrqS8f8Zzg6QQJ1EMyrZv6qMiCzesAWJ6PUEGwM6XYvFqWAC
I1zuI+sE240t/wf0+AQHrbSnPJaOyVnLRjMZS/vpXvw3m2lMOH3kBuL47OEnDqlw
OLSkfe1NSSK2PlZolgQd2HfU7/869oqYNZM3S8G1iQwdXnNxpPDyU5ElZBjjqbom
hYu0TaLVYMCmlcxvPalUrwlCP5ZmIC4j45nRhz7sCFxQgV5CVT4HOTdPx1cFmJ+q
D7CWlUWZXXSppPL5Ro7Iv83ySpSSv74QfWUx8w45tzrPctJaKDSubITYB7fpQkiA
urcruKD4YiA8c5+KXbnl1rz49wpj0XzJNdnCqhJMBpOOEdSfDCUsNRBGHPweIs25
sg66VUI26pzA2Rb4Co8IarQp29HUgaQ6QPwkuejT+Wl291XNTxXzofid4Vttgulj
9EEjkeBmO3NBIBNtYmRieLc0Mk+Xl443LzQr402KAwWXzfo10tespQt7Z0dbMD4k
i9rpviVKIKdKSFVlbns6hLElMq8LYNX1O4QknAGo1GNSRwW9fZBrfy8xxnvnBRKJ
PSKffS61Sc0B27zFoGDP/kzhv2HhbBMHi7v+NlA3h7QmcLk7xaevk+y2JQ5yOy18
YMcOtZZI29iQYBfgAH6kRGDFNVV83jxrC4aGgig8/qRCwLAEcn3cMElTUyYbBJpH
sKUiakWkBBXx8aKkekRtmFMR57TV3XZYDJk17T3CiEwPp566n8g8LlFr6AJ+jbUo
r6lfr/tSJGXf5X7Pu3MW/8ytXscOsC0x4iFfURbO21Qg5TGMpNbWiYn8Kpi7P+P1
Ikj0fqgaJVYqV+x8mIL6kj7kfDllALCOVpG69R/jNA3vYMNNZv3QDzkH9jcAMp/b
c8AE1M56/7+/BjPPaMJWjGwPC+gB8yeZZKs57ZqvpplmvxF5tP4C038qjRMimniT
jqPf6mDMv9mnEZ2EMyvlhZBqkJXYLzfdoAIlz9B+cBGRqpCs55ST/KbLdHjb2Yyb
SXlpDRIhiiMYdxiYN/wq053W4XQbFodQo4noT+1strOgqINd5G/61O7JVtN2MRf2
DkILPx66M0YV820bm95ihytRvB++tK49aHDbYLVnDqpygeP54/WMvtd/yfiZPp4j
DyWpyl+Pm62nYG8WJtHLW8Zofq9NtpJlIDecbO3z8Au2PKC4ySgB1vjsBcXHJqs/
65baNvfN2jWGkZp8K8SPFK0rLgh+j2sIOFHmGDz/ARWyd3ekvlJTrJvrO/AEuU7k
jcq7g7oAVn0iEX7klL3jzggiOklnsDTLialqmzvh4YuuD5WzGTpYf/k/BVA3SBMY
LjTA9BD0cMBphdR0eKX/hpu5Z9XDoqdmDvEEOl2swaVOMuKw6ec6lKoOdw5J8sZK
UIHfUcYmUEi3YKZKIzgi0zyKOO8CHlwb6VA1tu5W90RiqtHxtcS47/HbGATjYedn
FLTgjBOM6MX+g7NoEcF8xj0R47BCCAbpLfRmgMU5DYN/PURoelMivvdjVtJRAhVp
rShHe0MMEJ80zC//Fid9tTYcv5HtObMLkJwWd2g2zpYqoNozH+2HBn2Fd7Dfhg9c
LTUrm9SOADdQ7Yig2NuTPcxv9cIijDq+pf121R4W7oU0nnCTpGDEZy0aafIRfd2E
GQULFOhEh+4A0uG3Igu3HgbE937zNq8k7w2FAwfSOltvT0k7yPXJ/6qsiR9oUFmi
NUnQ9/SNa3KBzACW/wcU3NvhQxWeyx2YGV3MF32guS6lBuK845ed1vz6iutIuQ2Q
sf6mWTm4o/s3UAHYVIe5RQoDo0jNd6LGsdtJ2hZpVLLiOThsiaYMZbmYX5UHGlfP
04rZmaQ/SrUK1Ijbt6OJg4kvmj8hF2ixHhCB0llRonO9KBriyIvlhoFflSTZ3SOg
QUyb2M896bLQQv4Kmxo+R8uhFaVoIFHddD7JB6UdMB/EA60wTLtSbmjXaksc0w/7
CBPdQL0C1VninTQ3l79Rs4aA2AihsmqJ7wVOxhLAKpcY+u4Z6OcvnCfMeDahJB2B
JVc+wJGUGVPg3xvf72uT8YbpfKlfY/GiwXSzZv/PZlu83delnUR24sjztIx8N800
PWtOGnXjCygM+KaThMPZblnFHIVWGvNWaK5kTqYKji5okaQ0+k6l1yUJVv6R0rUi
xePNiKqud6Sc4JksGSgytatiR8XAhuod+EqZ4APZLOUFGZbzh52r5aYC5dY/cxm7
tVXzmD65GqZtpCG2AFyhYQkM+WbTI6jkBV6Z9IiEMdeOJ7UxxMR0F78qkfOk1Z3/
tFnJg+Jhlv/03e43Nxpbose8Aymetw/nHooUoa/OAtDQg7mE+ygBQW8keyXCalb9
+5qn5p785ek4pe0iOVn4xO6LWmB/jR1wdDhoCwlNpArqSnIOKKGIpbFiBAzqn5PB
fxyG/gGfvDCh6vBy+o71AIC52fFHD881Rjmpg1FfAYX0LDK92UgYBaeXgNxcy4+3
HuFH5ajLcc20t7pis7aF3+LJLz3/QNxKRqLlaUkFgKO961WcTm2MbHYXV+lDE9AX
xkO3/NMGZkwGb33eXZ9Jsb0aPUWiRSFUYZrk3yEsfXmU78F3v9MYCscpKk+/Za3z
6Ne03yZ3NeyFBIMxQkWxkJja073ob5edGbznsSD3kKQ4Y3oseo2t4YDYbDFVIGOW
zI5PXSjjKajUCOz6wtX3O+UyzFsd40V34cYhLFbDLiUCn/vl8imJq6n+buaKNT0m
nG4tU2POAI3bi5Yn0wUO44EKyYtfbXjbagySoMiMDguWrTentXjDtm0GvM5KjSec
HBY6FNHtLXwebHvudGB8XssF3SnFGaNgaMhtzwm372gi0f+CJED/8Bse32K0MOnp
fX3HjsVsWtIUSvqWWyAKkMKUdGASjIPqQq329yIe2j8y+sW+OTpFlNpeaQcbcGl9
bn4Xt9Mp0hCAbwTvNtbLAQGtT7xJZCkpIlm+YCTQOEkLw6BGEwBlkYtXoWlyxc6R
7tNDxE4qmx4kNaXtv1qfS5Fzb4w6tTWIjY9Iu9LW0xvPq2xokZpnFDc9YDv3n2Gm
Vv/ja7nx/6PljNJsJMNvjp7Me/IOwXD93/xLLs1SOyNYQXasccJe3Mw0S22VF8Fk
a+bsDNYbULPJGbNJL6rWVBT0P/UULBi/6X5UH/onL+bj5QiQ7LEaVKy+m1avvQeh
6Z/mFLOsOx1DAH4Z0ueR1utRFG5uAJF3an4/4A+dZd6ks8iLodehYXUDRCxX6hfy
YeumdUkp2hER56HHUwYzfcvsydKP8xmWbdpqXcfhdSFd6va6WYW09Ap/Su0LJod3
4v8lY89kZJefNnNQNKio0o1pcwmvnydmj6qCbK4j6P6Usao1RuAG/uvFBDX3xSjQ
SoqJPucXe06v7gM+tTqLd3mPixNcCvX+K2AT8BnI6AaYNeMoBffRODwsWkXl7XSQ
gDPU4RjP6GSr2UBCYjo5hKuXhoDYMirTEvYvZMuarEx1POfw9UscZLWGZVk7Hkdu
ZwlVK+4jpCJgTPI9WT2aasWCJWpI8JN8V5hxJ0+Hul8NaCunCad77G/feCNWkVTk
iUdn85r7zjFtc+Ey0OzzKoG2oSGgzt8j4/KuSYonXF/WS4UTnTyx0MMyEA05S4W2
wcq7NCvCQAwg1yDjvqA40HoloN1yUuIQm5Gm7xqr8pXkHftMs9iOp7WJHBpJ7bg+
wbP5vcVjPGHYY2A3sj+helHQnf3HPNqXj5MU9gN4XymiE6BEEBobEhBvrKar3Mgw
4xEXsRDZIwoETYz9YI99SzOmTUJDPw/aaJB7iQ/uVlezGxssRErblx/CMYbg6KVj
EyzAvmyC3PRRy/rab4XIpHS0lzDLhIrDfge+6rSPPF1bOth/pkGgeUGa+0iHgOgV
HoCgUrUqYzdsOB6DsRLhu3pa35UNWfwQgxJ0C5DQ/8kpTaQmyF41fn/l6cyKdwHP
hEAnHkIxPfJscemPej4l5IVYb2YkfV4xVNX0Mv88IUJzzCobu4uXWPFdA/dMcYDz
qn0fzRXOOq+jhSHVQYIKCB/8NxiNwJZk74NuSq3akF54ZPnIdZpFm7Mz/0aYMk2p
87HNFudi+ALQeuqjbCXKCEIg//s9VG682gUfRvOW7Sv6tQt1BpXyv0SjCLrQK8al
/vbeBnQX7RYmZh6ynBRRn6rhpWnudgRpGKm1XLytpbqz79es/z14tVBsSmI5Fmum
XpMh/a+yRSGIQEo5VctIzU16R/Xhj/bzIhI0nzpxOqRxH4vWgeSpcwNMyohFGsWs
jrgv/eI24pg4aY0UR8XZk1f5XFFrxi4jj6bpaacb2t+RqSrbSZ4XtM2mtKbtBGNG
62yjDeMbe9IWuBHL+UsDE9gw6YuBfYpBmz0+uXDmHktu8s7/T2Soys0/lAq0FL1N
mwNsfQPtCwc/2ZUAQpmh94GGpofY1Pkovas8SdsXpVgLqNmNOTxfo72wXCjEO0N1
OZlcEqh+TDMndL7UueBOU1CLL9CE6bOKpnCUYmzv4izmpDdhilqnQ00hfnsZeP3M
pkH617mkzaRsdl2XzHeisE5KNefRO1NePAQlHKYz27xvBhFvMa9lUFpE5Z0cBsOA
pg8FdQlXYNRXpm/OZM+oVFA/p1EZ4N1p8jVtxIXWg2wpDCJ3iHzzf39bkSY0Q5q3
a5n0mYBwZ26eFkO9jVYxVl942htsQPpgVjN4DNAaTIzP1j7hH6emIkBWm7aVHj9X
LESDBefim848caaYd6F2hU21ijkL6HPIdSVCN66SIPHuu7JFKnNXfarxd9/1PYOO
+rSKdtDHCLbNW0EN+lrTW3hcxmmaGwDtkWfQMwSNHqNWNrl2gyaXgMtqHcc3T6U7
12J/9PI8mcwtWu+o+bggg3KXMMFeA1AIXfW/rE2VIyERCSPdz5Knfx7boTu3A1Nq
ix89krs60/cNaHjgWk6WY61msSTBSgbN4lcM1AWZIxSTnrdxWdhZjhf4bEyKFDyj
tV1C9KZWoxCCNQNY20mEMJn7PLgFUFIcMgGEpo5JikPtEtWr5MK3M80zC3tEWGoL
443UQD84sBLaiYpi3IvUnfr94Z+gb8pEymiLHZpF64pRNfvJ/0hst5LYfeXyhxxG
eWO8ztxHOQhTHLWbX8RYDm9SYxcsnDJCygh49Xsav93SLF0xN0THYZ2UsaAiX5sK
5If6fjhCngVHKPiOj4mAsvJbu42bFPc20gyWXUZFO1clO2gbLs4FqF0dz86hPEUt
ddcex52mZSFLHXTwh+1hg6xoP6vfLCGxsYQ5z0eEAMLz69vZpUDU5QUAfn1JLT4Q
E/CmwOZJfP9nhOK3OZIVhEBF5QyaFVaEyg65LuaE7Tw+oU3LR+mb9kJjhl0YXKaP
EM7P2yNntSL+4BKqiyzmlN++ZZEE6GquWV3aqzqcK1OjKN+Mmbn8QqVWHbcme94h
EQTx6UCIYlBlSqRKgAJrUX0+J85wnK9UoeZS2gyY2c2SVLI86mjCBJxWQWjnUdEY
eX4gnon4jPAj/ENiAtqC/W40YM19Ej1P6qMp58ae25GIFuMwjBDk+L+i96MrmoJD
gIsDWQkslnw06aybLiD+VWWNK4aiETs+7bknvByx8SU5MTCWyUbVDnqfafNbBzT0
Czph44okQqZFUFdp9iLgTFAHOYp85K+8jg4jLOlSWCByKg3mVRDmLvIDpbAsAKX4
JHT69CvIBuAjmh5kCgckfxyIg5TtEx8JmDj5R6qeDoyzm2A6FNZQh3YX8v66ku9i
LwFH1nYvyvejG4kPmM95gzpZDwP4YFEQ1IOmfrJd+Wtaj5/tzwWEKxYyIDvaMCgl
dnKoMOp+qD+WsE/XCU7pVbLwznLScu1hQ0dixF398CxmjUCxSKjKsMdgons5j+mV
5cKqWeI7/ChPCEPadBg0tCjOZWKA9ihHgKAMYOfG5rn3pOdodwNAFFheQeXRt8oP
JYax/jRxytMNzXxb0KnIURwtkW+L8lf8tWeuzPCRVzfl5FnHysodgrgQ5IQOK/Oc
vmy3jCBuj6augu+GkAUTNKy2uVaaw1ISRJC26BwSE3f5tDkUEEZdXuKtEJOL77/9
hE2Yzz+7LT4aUqX0fBcmRqXdf5Ce3nq+hlBiw/J+8vBZMY2L0ZydTGDKgCOPE1p8
oNcKnyvLLNJwXzahEnrLqI3mj+m6ZZdIQ+DgUkbbHc/XTpq69mZBcHmjr1S4Ijm1
IotgGLa5xLO0hcs+EV+4oShuAny4KJ0ICLlMbGHK1ckStIp1rQb9OPd3F8uNrvSU
k8Bz98d72xC1sAlNKhnJw1/AJcP+YX+OjmMNp48JGYIsIls09K7vMUoqtHAir9pj
WfrhHEw4/F1RIXQu5hlpkpDqY5ODKq8NQceDREFu/3xdUQTV3M8JdqBo2DdwhBIn
PmZObDf97rVnb1K+ELPk/a2qBxVZVTnMLnIMgcLV4wVTclNgeHN5Q1X4E4oWvC46
2yfF5XSRyFdkUWOOaxDYipEaRRxSr6YSh+B4noosz8E0otI07gzuCKJHIcKz41KS
eFqYRdJ3OkVxmnyYKgSthZx/FyIaGKoxSl4buQvWILcxopoph0pdBf6pJeDZGZff
Mwg4TnyYRFovVaczcvIrvcjE/LgK5XdETKzofZ4atKVpTWVONcaXLgOyGiWMJy1g
RT8yEkvSDGan0H2sgNgnYhZgTpEeL+ysbIyXFqqZ7gkhxZcvCkigmQRO2JpxM5rr
nTAtaJtpFLyS1gO2waM1V5kcCBwol29BbMbeDlmwk+MIPcNeT4YrFVyapgDeNhKM
0WetnGs4Z+AXwytB6CY1xb+7WkT5HEv17Lk45XJARsGAWKEhNqn2HC61aAT5TfH5
/bw00GMyJJ4mKEfLCmd0LG6A9quST63Kvu1W4I2+NAPUHeqSP0BjGVjmpMBHRA84
N0r3fPdgob6+AW9Sw2y1NI1ZVrj9ZT3L8kOBkpH21wnQm8iscpW468ADWdccT0mQ
ib9Qy1G1psnj2CVAb9jbmIpe+qCSP/4vpO9RVSaIOOREW6E6+NCq+0iUoSAMUm4U
2af351rvTNEq1S9tMXRd1ix0UO2NZ7ALrFkpvedAqldn271FUgKbKkD1tEGCYeEB
KjbwgDCyq2tmdzAQ7PFwzmjOrq6xINjKIhSqV0NQ/hFdSHGOHX9VNWsV8YRFyF+D
tHyLTirKOvCtJocMeZ0lzFR9zE4JTmoEGZnnHmvnxvmS0U0XPW3JODuBO3TBnFet
4F/CX1azPajIAQsfciGM3vlK2bka+hdukRWKU0/C6+BcwllV/jO1fg1Uaf9AfWgv
xhnvVu3lF9cD9kFuPDACBOd7GUKdYuv3nDCZ2jsBw47G+LJ0HHmi8x8Lrm7es+Df
MlA5+xUkIQxMYV2c9CSOdABFggA7oIt/o0Q9VSDy4gg1MjRF6BYfeQZ7/jrjVAvb
q8dWn50Vyh0u3zYzO/0NaVKCbkiUMDSTrXhL3Dudu2yf//oSXLW85xb/WuB/XWkl
JcRWGE+tdUIdwHDTtsiBujNN49pvTn7Q3eVQCNWry4NnqxbEN2wAsuRHeuSbvGkZ
apdcWHO9v/GT+EvRXrbvAvhA6WSheR3/mIIW47OE2oluqxUE5S9/MemAzEfq1eZ0
2vBmrc5J0WLp6HPVi3TCjhCRyvLXlo8haRDyy+A2gPuMhXuVSme1Y+f25kYGLg/F
oLUix/bbJJkFGL142h52RpuJ8LpoIk+rb/QNJ51jjr90HGv//FfTlUW7C4qLrYRT
RXIDXg4vUGHr9wi3CILIvqhFvWqayAl9GA7epgP90tW13SQFPZz2L3X1UNorske7
yGaZ43hx0LO4Vkz60e+rOI4ySAac0iiaHLGYrcQu3FxhEIClkzrh35Zo5zwLOIIy
9ERHC5+F5DiZ3m4X96Or7+sKIC//7YB5o/D8AUlL+gU7ST1Y9jHDDqxj01wYOEm8
Y/L0mla/RUgYLuPZ1Wwyswzde9AFl8/xzTKQeAuBnuhhM7cDrd+JN/k+jUD6vKRL
SYtFboJoJMTed8Ih5DeBi3HRTaQKNg2EHll2yTN+WE5W/fvQKbOCaCzagLy5H3S9
K8uv5wyzJY9BQVe2fjtsz+zYhKLqrNdWI328NbRdnZjc1bfHitkPtmroh/u19a96
ANed5DjLu5fjLpgPDzQJIKSamHoQd2bZZB2qylQFP/cr2DUNY0u8nwpEoxH0jHVw
2pyNLppX8Q/bZrLuJTcvE3JcCbceNu4ZFXmCmbxxF+4E2ao3uNfBUIcbBccW/1vT
mJyQzHI6yPw2DNYcJpz9QZjN8rSbeHTHg6Iyfj8D1964M7lSj3uOOaY3nDdTsc4G
11u35xta7VWvTB46P1cg7KS2lsyy3avkvy7diCJI7ukn+B9digJP3oHg2v2iEhp9
gOVR6liPGMYBquDqRw5zicqhIr0Bw9npLgonPjbghmfxHkpwSsX4xioWSko8u70x
KzZUwcLBTjs3oWDaOvyN+NQIYToSTRxWuHDo4PplIFhOD/J79Xmt8nYWHmpTgguZ
qqIL/JF8hsT0nKgt9hsfgvNV/g+cajA/Kf8Axa1wFdHUMmH5NR5ktu63PkBSskyg
/TXTPLk6MhWIeBRKpF1oqL1Y3g1VSlvKW/auwRCP9qAMXmEwNX++dvKA8F9YIuQB
iTHTBVcbq/HY5CiVZsO0I1pQP/s1jS7Mk7flKqVZG5wkTcJWw2ErUl5/9o0y294c
mq54eXPsnqzMKy8qFf7PrjGy/WJiIILfwfnm/gZGLBMXWwtNf8cFpZU6tW4E/vBC
vU5tsmBq3Uk2ZBY+2uzop5ZbDxZyv4M+QtYs8jckqk9EC1TruHbBjV0lRfvUnTLa
Cg4nwj+ZDM2A5vf+cTgWTWuN4I7IVnlAaWSxMm+yIlAbjp6N19wxBaa3fKh+Y7Tr
9oP22zlgHrDfmV1J7lpz2xV5QeAXenEhohT2fA5mnyKMkl1pa9wMeElSC0nuYCp1
9u+PP9y4xfPpoW5GcidxXN36F7STq86rAfVvNepscBdEDYm8dq/R4ldXrqDhTrgQ
+yBoy8+5cYNcfrvkaldSPwwXHbjXIhttPKqMDqbl60E5igQCMnwsnMcKnDEebJ0t
wVjpExq1R0CRlpF93KNSoZ44wGwW5rwp94g1QM6Xj+SSpMvAHH/B0bgxyuWxta52
fvWrySV6IYyIlXrnJCcjOnA6LHxl6+3UsrA+u/e77vgHlE5i94MNh3hGHt4SN335
eX5P9Y19vSWC9hBBBTXG9ERYCZ92XNE6dUuYthOfFIVVtKHlH1Rnn7UYpCLFk3sP
J4YrzbLLaacNyrB0sk+xHWBSIAaEG+pWo20e0TnL4yAOz3f/n1wqFeOwKiRkJkQ7
odYy90UmmVTlBA4wjB4+hA8By0/D+NVgQUZUHK7E0yu83ACNVq4Q1efhjicef9mH
emmbNr74ibWPqogu8IoiTtgYOS2Mzvy+SgP/lKiD/ZzhtYTHQcOyvIsxYtmSyZVe
0tckLiaxJOxtHYgoTX4UkdZ/OGSEL12RSX8keFh7dsIINnFqT19nhWiLMk1+AVcf
VLtsVcvu3OH0AaXhrOiWnscWVbg+Xvb+3J5KymRhgccQiKjiA8UYIt6bV0Ht9Qd5
25VWCQsxuHGC7LfEsS9MPVcMyDa0eEIkHooSUD5PvwnWmQqXMl+xgnvmgoRi6CPA
5DToCWsCdfEhR6Gu6bpNf5lC98DxewePWw1cbJpJRT3wn3TNGbeLf4B9zUTM3ZDZ
PobPfQQnV28neY+bei+OEaO9fShmuBYi0MGsupw6S4oQ8z5rDxeJy7Rs3kX91xKJ
7yxcOgdfzahLMjgWvw/FB6b25c9eyl/jfYGT5nKfRJ/1KWLBY2KOLkoEdSyS6Y6Y
vdlKGj3onsWwtP/9LoPdA0GIW/Lr4zHIjHlT7pnZniBVL3PrKX0Fy0grdw6q1ggF
gQybI7e1taNiRilIFoZ6w0xqq8wMP05I7kNVnNFwK6xz5/IlCtrqMH3aRYOa38lB
FPJ8037UOmyTRGPxM2J4gYjggUFqhE27k33kDeY4nsLJN6DJkJBzbnwIzkzOTizg
VLv+B6xaSdoPJBIsFz+jdhKDrFYpmKY2q04wGDlZZQh7vFEIu0atS9lwMurKUMXO
duBFmPqW7z4+ZRaU9e6XcNDLceR648RxCTdnkTax+Z7Th5HBUeBVc9Y47Uc/kYm5
zPS1BOruR+VhgdBpwA4WyUOyWQ4N1Po8tb4AS51uu0AvOZ85QC32EtMi6MqYcWV7
SshKoZIgIQ+wSZPvpU/ySEdcBPcYYZ2xfA1X1xKsNNZvrVSkdC/7uRUAqHcBeHkc
uDWM7IkiBLUiGYxf0Us3pRCfQDrFV8QxKtHKEXqFqRRzUm1TeWYyhXVCuivb6Tju
P6jTrLnRbk07wlzVfyqF1C8jMJNnK4AbYDnV3mGq2juJFMIshBc57Xv+EDMAu09i
kxZCdJ3cf5bNJGrQWnX/dpz+t4lsIi09U7suWuqyzk8QsRpAcn8Qbe2mXY1kJiBS
/20WPxq5xhWk3zvP3c8YAePncP/W+YtjU6Ke7Pp554E3kakqeOKrLkTLVQnAlOoV
jnZbQEN7z4tbMBNayWND7e5KTplNjIeWS6ZEK1zl5fyPGHUNU4EVEMYF72cqIX/M
KJWvg4q/kg3XuP/DgwgE3bnh2SoqzlAdgatOsjxbOr2ka+s1kmJceGTvdT7daysp
jOh3pGu+2R+BOfLhKe1TsqFPTE8lwCD4Xlo925NKSX+RVjX61KmCq7zPvPdWogk8
qJkmY4hS7Kje2se4CiYe+b8M1QIiEqpLjqWPmJvXR1jt9o1SjOYq4Rrzl5vrh9aw
f8jRip1dVMqXNMhzH/1CihDGLCli2lapzZg0ypQLQBAyG0Lmyn6X5ANEOHEkdsl0
R7UxYb+8znGaLeY8Yrx0Mf3z+Pv/E+6NTHyzvRX8knqjsE9bK14fn64sBptWk3kg
LNC41Rm97fxatGC1mt0F0pHrTonbdM1mVsvNx1x+idf3oZXZNdGu9r8r3i+vCw3f
CMgrQA6lkFYsz625Tk4JN1HqRM68biIRmgofH3rIvIJdVx8cwKAOwPcySorfS7ei
yt8LS00NrtWCvdV3UOqEpBadm2AzV812CEoN+nJAlYaaC5qUbBlR+Wz9q1WTXrId
No0gM7SBpZ8wcJfbAIjgYcHMYn8LS9zzImPjC9aKtv6kFBEviF68MqIQGEIaqeIO
L3nm/ElCifW639E6PremoBN6eb5WAGE9qIIvS2POGTALkD9AMRQPTERdeTWmkZui
I1BQvNVovYSJ9UzcjOUpYRulyCEo8duvb4o6J84ctwO8W3UA4y11wTGRCW4MsqSN
A+U+fV8FN5xa2krTwaUPevIKo3wi1zsrltqvm7YTU4RQfFLb9zNx8g4KUUrcjR8U
Q7spR6K1hPqiRdSAwaPGw8B9v8jO2KZO8ZjFeZSM4DSeg/OkZL+o/oJKwxvwlV+/
ibyXmOrImKcj1EgnZiKTQk4A1vLtvlXnAGt++AhnwiHrG1Dr4DhllXvwECEq+llw
T6IdjyjoP2WiJcGidgUIxVx9yzc0oZgUjVcFD1TYprSWTV2OHh+ky1SkDntvUxen
McnV1Swjp6hr30BKAVuO2DzzMihEplGaJK8cTb/1KjOjdvljFVBDsKhKZ8TRTVHi
oNk/Fw5FuRzWnNLilnDO77GhDOG+1AI4c6lcNIqsZKzVu/R/BLpjs/Z4jLcEcJd+
A8FaK2H+3sr2qQeTS5F1R2ZEfDF2/dcfi7hrxZ4nPndbN1Xx0HwSgfMc2i7wtDpI
WJONB2HzDsyGnOXw6h4TSZ8CtMOgH4gD/i1/N4WJFrKWAGn9MMe9jpti5X/ltHHp
N2/ZFBss5RP/GiDCBojKkLAcXs2U7FdK6KG8eHx9ouvLDBewnFPaSBJPFwVZcHvs
pwKVsiN/JldjAwp62hRHnRCpQmDxAv1weJLHojhUwLP3/Nm03VmS91qO2t2qv2B5
3rglx/hu7Xenfy/SpjZra1mmAzm+IXxfbq8rMIHUFLH+MgNiUSR/f5nwgpp31CR6
e0lsyJOos8pmpKZXxE9sTdvwLpXkqZfqVCGgI+/njpHypG6W1K6MiLJYxXIRsW2Y
+LQLLZ7HuMPjrZbk5gq+Ja3oJ1Dbm3yiFexepXxoXvo2UMW7XRYqJb7pPcAOfp/o
PT1AYraq9ahM7i0/2LmQn3KNVVBm+850ytoUP6F3LfZ/qup3BJlevyb1HdIUaFi6
tA9fx/Yo+MQwmVXDbaP2oikLkfBznv1RyO/WkUJHD22rhRr3oAmf1M8bCsjUagUv
mzTGaZDR4hJXpUAd751M3oDZcdwtCCiQyCX5EJ8c3zo/BnH0CGw3oHKtiUO+In2o
NeHAqjCwtc6ZfFSkKQKdyP0hI5ugONCwdh0yshH5lrAgH0CApicyO1LMOe/XHKZD
UUrqKqxc/19hdPoqx/6nC3AEKQS1nBhFC0WWDxtcC3iYby2uMJeldXayk2e+6XE8
BH+ypTGw9ONqEeIIDAM/Q6PQzLSUSUu9Jth4QA0s0eWciNbCwd14bcAawb0FkhKY
IjX7dW1BCjtJBFgl3nORZHe9wEkQb0K5HJZr5Tozpc5CGXRz4+d53/U05nFGvO0S
ES3GnwIKJfqIcmDPD/J8OxGvAa2DHiasUeoVXp5X9mYAxnzKCDWgR0yowUpqimZ0
16itfiORSQvE4Iuz7iDd4edNxBaN7n4GKCgmGySD0/WCWVXAIL/nH87Ei35igwfB
Z2fVsCEMEyQe1SfXFuXClP2wGpgEldHA6BjtNXI0g6PfsWm5ZOVOFZdsxbhOstGd
bDzTilaQNEmZPDwT9FqTlJOfAoAeNTEI4KIj1pO4YKqR8GbFLZ7qeKx7kCPHZJbB
VCuchNggMm0C8nK+VQkELf6HejVop0jgR3HxY+N4afveji5iTp6KIBwJi6bJnTbM
p95GHwmJafjXYaDcoyOv+g/CMyEkktSs+X2SsaqvT3MttgTxA2lSWgEyiAZHKz3w
tG7xCf0NgTVzRxXlQRe3unqYogIFlDPHeZDP/avIH4qmddvm545Y6HCOgosMvHaO
/TzQVqaV4D4QEQW6MS9idSvteH6jopZbSb1maVc1TTihPFylQfffLRaAf2uRlOEi
004UL8PIElMkbLE7Bg6vrHfZ200qfb4FuMoN2EwyHmWbYwBQ3x5joiGHEScLmnHa
M+MeunxHWmQWLV6T/H+Owbk080Q9qnvWLd2Je1ok5CsByoSD6YBjhXYW7hl1OFp9
y4BOAEPFgje1rOx2FrBPBooNiHxro+x+/jsvu0wPNnnk23TgSaDKJZttZaMPbWrL
aRTZB+FrNVUrMMXQ9dFqqKmJKiTALc/8UCuXWYc63T4zOFAQUsDg2B3aJT5s59r0
6WSPvQ4U6ozyMYpz4DKVqmUI42LvdhHGnmQwmGTe6UTrRXxnZyLPWCch9lTdZTXd
Ca000ueu7OY4tryRlFSKw8NhQpy0Ehfy/JoT/Y3h/yQka36Z4kooN93pZQznZutm
tF0Hn7uh6odHWLaM7bncuZheboqgFwa4f7O75mRWvBT5HBpL0Aedtw8YZzpvDTrd
bgSUYZ0e1jj7M23QFiWw/r+SCt36Eg3iCa7UJfFoOVHRaym8Ghz8fmRUGWGEe+s4
n8tspe0HqWBL0ezyMuE/vh1kvBH2vjcyWpDWQ3gRBw3VH7X1z+5YSi74X8fzrjHn
q9BIvhF7Z44wTJbZOjnOXyDt0maXeExINgCQxnsPd/oY6/rQ6KAQxhwvZNbS26o/
F23arIuDlDPpJH+vmOlJCzGo3R67wl+V3vTRik4NzxktcxcouX42GL7QS75mGGLi
OOFU1BliJjWL/Ucaiud3/BbqYjuM3/RYcxKTiRLlocTMo59Ahx/iSlkI3ZdkWj2W
H+vCbyUkmqAeHvnDDEge4kiC7gsePDCDmM5r/3KP3CNNWCGOQF3G34KCg6tic3py
bPGWBvzyKlmoPnosqIim2wV8sxlK7Gcat24tcyVW0l5Nxtok2V0feGnUqIXgSRan
bCQHhlR4OzLkdHm9TCdv2Hr/3/W+Amo4AfmFE2qMpZdJQNs/7guMow7InN0q9OaO
Vqaq9FaClDPI4p/Yiaa10RpQTB+DBcmPXT50ZPaounZPSnh/O2aedrVCjfZrVkW0
xWUPZz0W0CV48nEJzxwSey68Zp75x4r0aY3hxbDIsrevwN2q8Qf9hzxTZ+WM2Xok
Ig2aj2wx+oBpIU4wOmk7j+PthOSNrcPkPlSoc8ad5C7BqXl+jVT2AXblWsKbJapo
G0GjeTIivyNjvXYXDHAhB2WF1EOqvLZtJSHF3rnGEbUR18GyBR7+MzrONoMbFy2q
kG7kxTE3VAMS1UHTUOcEvkmdOo7HhwhS8KOpAq5UhfUzGhprg6r6uAgVikN5DPtm
AdPFS+SKKOWeEtwjJcQ5QTKeoLFlPPHF50ChQWfDxk23H26Wpl+UuqRh7TSzJGzI
N7mrIL/hjA17ErEDdqs2axQWe2HPlROiqBji0cjIvCtEYSGiGdDaH+FTbEE1MOSu
ru/YwkM8Iwq2VdRmZLMfOWfUQmY5oTDwA7kgpFaSbq7mvcWdzaNzOn3ZtspUrm51
yS/jsy7lPR1KNATJEJuZXDV9U1OaCuK52ZMTglsj1LKIcoFPXYbMT9+42/p4N3zT
/w6pB2oyrj4FJslQvnI/lVXWMjOflws8CLFFuGgRbq4rXwHwIrm+xbWYybn+4J5H
OVavkIm41Ij43KGLA4jj9zmhLGf2TSOAA7PdxwSxSn6tkRJGkd8hmasb0EhGNdzB
0Ot93Zz+0sEoe2dMf2AsqnWgTmCa2rls+nYSxMp+quOuLm5TLnyR39j9jyguau4F
Upqat0QcnUZ8+YeoZgPEXk7fIAjRut69IqiwSztJbKe7v7G8zSG54SJn8m5i0ZfC
q0OdzYzVuufGLTAUSrwIoJSsGSPfXxstyFekTjJ2tmaKGMdqAu0U9h1n9bpKUx1Z
/b0LLEk8bz+3xBVvJQa4bDEebISylmucjPCxkP61uQyVjuIj7pJ0nxW/me8hdqur
lNCea5FLjVVGcwmSErG5gMaUtHZKj8tCETQzmXSzfez4UcL6CQZHDIk5ncWtddqA
3hSWZ/80X9E3nzmRewnzUhzAsfdYkmbV2YfxrFU0dGN/JkMbLJ/HrZNkOIow2vOr
26jFMa1xJbmYCN/pd5lRqHQKum6jdHNNgZTO/XYrCPQw/yjPjWVVQSZyWlvcknmI
wQkPuH6yjiA0/XDaUuUkG2X5UAJ33CKnJ80MgMHumClumNd1rgVe0uSylEUfGYkl
IrAz6QkKdnCIn5cRomlfaNVsp04ImJqx/FQO8maCJysLYpc/luI4vSAtg3TxrYwZ
kUwv6f2i/P+17F3NOZWL21ES3VoDyUnz6X3ehtZJYtOY7S8Ry0Ga8xFdztUk3F+8
NxBE+n5APAMgfESeb7ALQkPzoPjaTzJjH4mGaSiIcDLGeNOlCsB7g8/OBOUT6+L1
CEiTbEYWeSQkMvFkzlV0Cvb8x4Id4uc8XW+SS0VDY7JD0fPcCNra3KqP6VWrenQZ
gxYHbZ37yWBIp7nrjMxYdwQR/6MiHna1ql/EbJOQoWmTNtCeYvz5PNX3SsKmyzZX
ABUY9K5X7I62Cch0xrcwvt8DunT/ONRut8tELoMbawwhhk2lxeNdXIR9JPECz/zc
lciXVWGe/WfYAlXFRPgiO1huxU8BLP5NgozFzt6QwV/J+IViC5yHByxlDo3atHUU
aKEyOJLUuKumCSEf6ktNwpMMFD+Yu+VsWZVPe1PhM1FWFX28qJ8C5fl98oa2PX5B
v7LlEsAEJaM9sjMn9KLUT5/ipBi4HOnmQH1F+sv3pY0vCE27sA6uAATwZdV3P5oM
tTn1Yi6zFKtVYIf1DOhgYKAITtSsXHMCTWDctKDPqA7DiK9HzKUTkQm0E6YbMwAs
bOyUrHYClxaVaVbOks+0Z8vqLoyMnlthQvZmLvk5feSlURuwHgToMMDrYw7gYPPO
IHf/FuBx4rDvJZ3e6wKrTLd0c6ZNh2CbnQB4fHqEYQb6PiO6fFfrfxDf5gu9oAhj
Cd9ZD9jMyzBvB4Xk9bgi9a4BxlhB4h8czT2h1n6xWMfw1OO6P/TjPPnbBlsw4VYw
Ee0WTHmfR+28GTLUlSjsb+CYMp7fdRBDIpEgyhcRZ6IaQAppmXkfpWeEG5Y3XD60
/s9UkqzS5vSuOOLcEaQZj070vWRssMQtVaKpDmaiSdtYZ0SmNgYTc75tFSnskUqO
BRhw5amgTR4seSehIuNWSwP7VI6mokbQSf7a1anG1D0E5Lr1tiZmB23nXXTAZXIX
4Sy1pQ0RsWwgwu8xV+F+mQgFC20TGFbKZDQy/QdP4+J9uC6+mKcc8yE6rPEAZeVE
9ennvRRdIhaKddbB3jP2SNmeCMZgoc7K/C9o0NNukVLaaizJ5+34NSCxqF683mZd
6C0C/b4Kz56G2VMVLcURDzgeYuJbmrxR7+Yj8dxadY65Aiil3V7d9n/aS0jvR2BE
X5jhQM9twnEdipp/cu6vO2vq50dQgqidQDi6KwB1OPDxRrFHRjt3RCEHJ76GxNyA
7QKf7r6nTrr5ZKhcSOgHKSSpcgoiJBePYf0o0TS3Udyfb95/i1IUynqDKb4d+Tv1
SwumW7Fn3C0QRpr1iai0rQVYQfYCAfy0JYXJfvPhSa3dXSEOJ+lt0Dz9EskBf3i4
609NlzZDwT01uGtvmfvUnhBZYtIRaoMgeyDXZvR0sEvsl/jX59qxJ4dZQAtNFKxJ
/XsjuFEEpYweOAXpd2WlvJLR8mC8pz0ODKGDzYttkat+DCVSdcRqShZOr1gzmSQb
tbrAipS4UEe1QuNXhIS+XrShA+7VvlNfTlzaiaW56vw1yBVVOektK07y0hyLek9g
zkZkm0Qd265GQVonMGdSe1EqLjrtbQv4Dc4f+owumDGE6eTSbiyeHAm6U9N4WLZn
9Hrfob4ldqqzcitT55tPjM16ctp6DRfOICdy8PA/Ar760Bvs7WwGte2qdWfDraVV
1fE12ywK1WqxL3LDIZkCfyfdndISGXOhyROVsTUSczVeD/ArmgpXoY6ILrh5PBsB
Rh12dNrDqlrxtURItYQtz58w0Yo4i443N/LK0eTWCaEF96i5cY+Pj89KD4AeRH8P
fcTMWI3Ie1N5JldOQCzVF6v0p1c5fVEt+GgZ5E2a9sCS1jRfi1SKOzY7EQMEKCVC
cUVCN0hZuU4OU/vI/Ouk9OGh9ODVwFmLXWrjs0nUOnw7SvkEhiAlTMwZe+QZ19H4
RJFBKaXTjFLSfUGdTHORgzJ7qfqQoch5IcCyFywjmzuXqOsken5QxHIwQZ4TPbmv
y026J4MRt9afMMgMVphhXLVKHDjqt3omHaetNXpArkdQhNJxk68dwVkm/3qtY7Qp
KuIzQgI+SWkbDdi7M6Hn9D+f1J6uTuNfH7mmh7PIFM+mBVR6IaruWWgHzl1t+c+K
JHIiQkujzo4SFL2rKplBJGsnbjQcV0v/gMgso+ZL4LRZrFBQZDbWKOyn2oXiwLBB
0ipFxLbkRhDeGa1dL8amYwZ5Twq7sLzzP1DVNLWGEszejDCYeeaZ0FzJq8sGN3m9
QMWhqqxoOkElapiiJL9neXnRH5LDVRBkMn20ylqMgHj9mg8Su0miLNsVEXCvsPWH
8iX/iLEzTOiOSiE7LDI5poC01lSVQXipvlO82CzkBwcb33gcrLnFx6Dfvhbshnbw
6uInHa6QndfAWuCTXxlWl1gLmajqSGUsKeYAWnnCjD2/LFE6Fm/YxvZMh4Mdpzjk
z/gDSKS1MjQwEMnsbVKhzmWvvdq/kF6tf6qy1o/cvaxG4sO1DGBE4xNZEdvQxdcT
e51Tl6IMKZj7y4QUTL8eabOUMCDEi0hEqUDZWZqGAXjA7F1IpbumQGdwEAM6DsIw
m//O3ajmKFKxLgI/hgGnRQsumQCAxv2ZJH5qa0ykeRN5N1JHVO93p8trqQDp+DMN
kjS/tvz0pAkar8x2owr6Mib78k0Es0R2pdF/uIBMQoZGyRcLZ7CIWFT9ksRrgqzK
hyBO1Mqsdr4xCZMDFedsb4r6856ZGIqKFvjZrd6giTqJ3Te+mr6XlhU+ORPMtbUU
hpXuUnNUGBVInxdfDdlx5lj7vHzMDdadAj1FYAzIc89bEDMU2lv+JV2AN6Ua72Kl
rn4Vu6nNxxUgJ1c3JYV6/9gYwKrC+QAzDeqHh9IEMfpUNL/QwLH27RYA32cTga7l
+D+F0htW7GMk8ajtv7YAzo98MjmXDRo6zL9Nr202zUJXmL1Zif5GkGJ/6YgCj0UP
evgKHIbgPIfeEAezr0rch8krdaAq+1OqfsBw3kDYe1jDYGrUivVlqHtEkoLy4TEl
fJYb6aYQcy63qZSHdYQEmvfG4963pytPL5HQKaNGBdS0scnZxQ86hYIg36YUekmx
HiVwiXbcw5gWt89+KjHWWbfY0nk8z7kyh5cwFK8YyF3kl3iApNmSbbwKqrCDoig7
CQwdH51eEQunWjfMqXuHraBMBV8Ev7i22LZ1YNlhozM42fTpcMpkEFHxPAtY3k1B
VU42L4ZpbY93VZiu7oIh7XQM+EwBXjVaoXQxLHXoPvpevi965Sd1+hehtb5j2qlr
KTPeB8vlFxTvP4t8hkCS/1ZKQbcG3XC/QGP1sX0fxEr0At6udpRPIGpi1CEo1Jnt
Sm1Y9kkf9xdn5vDIBML4FcSAkonIpvOkf0gfpeWR728dtDxwZn+53iW+p7V8kIBh
HcGbJ2lgsWyH84Gldoa076pLVbcCrIZ7pQfGDomHmVmEGm5YSuheF70b1DAZQJyD
xwHmfGcTFl9J6a1sfV27JILP6Ub4QL+gD66I9gr7MB6M+vNjprUgrYTCw34WOWtm
PnIn5/P7PV9XwhRAA4cr2qf/1PpUUTlRM5fZYVSC+PAE3yqaZctHKGS0954m4xhc
OhijClvtwfCWHLPnDQKeriIwWaTUH1yU2/Xaun3WoHbRuTF9disD0Kn432K1lh8Q
KJRLWoFhu8Ey6jFuyKOscVKi1jq4F6GLdMZBX2m3zVotZ46Wg5cjpu+y/6lpfabn
dFnN2qaQXlLMV1iw/bpFNSHT+nlQB05QqQ0Gh0zjWDzlw3T5G3batfEr0S3jCPhE
aQnelOXkBTpI8+5X5EO5t51t4u99NKDpHnTg+zsHC0Lma0tnrMJHgNSIRXZQR/Ut
78Us1Rysh5qJ99g5F9LMXMbtQsOHpOqNcq3JebKPw+Lhl/6+tDYJ7fPd4VVhB4AJ
Vq6noofHpgcYWyXlMUQ1S3hRig4h3NZQD4Oybo8MXkGQdPMkh/cq7PKmx8uCyGYf
tQ/ybEfECduBiEVhJrbC7tXNaKTiDb3+ngBrSf3W7Lq4hsdngcfCjOpcuaWuTNnY
QaockHDFg/JVhV8+93T4R7GWh9U89E7fb+d/JcyXKvzAAkm7kZ0jN9COirFNSbFb
NrYy95DChZsLlcRVgGXfKclxtUTOxFArv/rWcFXkOIh0YjiGYFq7q1wNBqrIyj31
ilPvvTi42VvPEFcEFGnwcpFeZrFc7BUZosnO8tVyEPENqVpSp97RrWDKeZg6QtPt
J+DbdIWhsmXCnzKdGoG2U5nEaf9eRYUeLxKN5Vn/Flp8lybpEkQavlg5TOsbEmb1
j9DGMjVqeohGGb+GWRpo1WtJbSWbEIYAchwzuo5A38VAA8wMTNINeDd3I5cbxHZ1
ADiUjwXFowwZ4Jb3oP4Js/5N9ajAAYAbLCPM/NqlMgJmGLDwqgJNoBbBN0hxpPsc
TjbuI7BdcjkLckVckK9/SPO9k+asKmtuO8VhiB8+7SinM2d8BcImu2yMA7RWHq/I
hLz1uKjo/QCvvkNHOQg9hMz8+ECzIFdHJydY2BNV5Qopw7frUdD94a5C/XZQzSkH
1V0q2ntVuCo+4KvHOTY8A0FfBKq3ect2Yqd3JCNHRXY1Q1wW1GX7AmXbjbrUkcof
VjtSSrbmXyUXThA8y5v2E15iK2fytwUTyyO8Sn7IuGb5uVrk7J/alo28blM4znRi
XHkPP3RwEguN4IEWXBYTSvPRzdKsQH+omTF0asAOjknCck22+iY0U9Wk9sLgM//G
0oV4TVNT9HzsD5O271gyCRbfbSc7mKfwfBn9BZzcl7LARbO94pukl2cIw69JzTm3
jtldbtJ/dIO0ZX2WO5yDAaJTCnWD4hWuR3dspnmlbrouZCg555TsxRSKCDVE+NJM
llIB8jlj+sVlOsdTG7KdTwqN5/Ve05sAhiXvX7UFDpK6kjmyPQsOwMDRG4C5LdDS
ClHc83Sdq3ZY94nUxxasQiiZxOQKxO6rfNSo70d5ve0eQI84taVujimA66hrRg/N
5I4/YJfdGfpuvqcoaczUXiHmMu4Vw54p7duCoOrDF/XIWFAp/+7sY0WUoExn5Y3g
HA6KlQvNkyG2Klt/3QvX89/i1iGfsgCBa3S+ByKNwnlF0t2HC1qi1nU/8TBeJesh
r1e56yf6WXM+LNVzVvfFUT6+cBYFuUgayTGhxqYdZbZzw1aosaJVqHMX2OtqTsl9
q9Yk/LYXvGxULkzZjqKfBM2H96iQw4E3nGAG3NCzthfc2eR2ptM8R9nVbCrO6YL4
iWrLWhloPdfW+fPGDPCDqDJjcPUKJA868bOgOsQCQBRVA8iw4MCZHLTAGfY20YGl
D1mq7RoUnzvpfcmmwjatVEjMJ0wkLJgiSBhIWBB0TWUn2i0LXWQ/4KKaLXzti//R
EewPKFVV9VxI7POik6ivWQW4J9vJ1BjJpTGV/B5qWgzz1Vhsrc2VqxIGeoJn4Aab
GNLrBPwGVtU5vRbDXCUtlf/qlqrc5C4w9VOjFXVa3PXNkZVaeCGFcBvA71SHFYZO
uu+1ipt1Q2DiK1aS3B3xl33FB6KWgisW1mBvXGgMJm5UFTjz/91DzROyqoPU98pa
mYW2cIUsWpRfJ0Wb0KYsRQRr0ebW7X7vnO7wkaIkygZkUS9EQuNflgbxEUFYFWlJ
9m/GiWBggGrBZL0EHJUpBH4tCpI9FXc6OrfUEAF7LEstWAFGJqvM1kt/nyj6VVnW
rU8xr3QGnmSU742ZjnpfXq7KmMQXEy1K4wjiZbWPngZ4/ZOTDC6MEV7BSPuM/1RG
Id2iLFrbUK5FA+txN8gW+JnT3o1bAk7lzeL1mES+jYIVCbQOV4RycVHyenUZ6JtV
6uNINdw7VSYl7liw/22C70cPwGhwpDIzBOzKfmeJSp8vaKUsu+x3zORi/TrZohgV
qlnNrlRXZC22uMGEuT/f/n7UiEn9wYOLH7JkJ71FNvhDzUznMA7RT3HpSvlQcgDI
JU4ZvWkdsbAy1sFvLGM1FKTbySaIjqt4x31/gplzpryNigy+REZBgmL9FbUc0qMB
MqFqtR6V8cstXpgd5UwjKG+LUVKdXMfRZitK+aaAY6Q7IYGsj+mwNapP5vLi2MTP
RdU0l7qAKFEfMKyFYOPqGst/f2JZ6w1Ln2im4tBRqy/N2l09pWpAli5lDk1GXr4R
JTPtYbeU0IgGPzs2qxgnrmB7PinFyHwUHUh1005aQoRWD3Nvp1nQXy8n8zEhNAdr
QTCHCJZApBr12fVIg7iw9fMSz5wSfRcGOMBAAziDXp6O+qK4946/3EkXkAJ89lvl
gvKrhjXAMwFD3oIj/QFg2M4Dpl9F6wVGEg+ljjc8lmTfRXIDjEkAywnIEpvwuoFJ
4q1mNdkS4rkAehnrDrkT74pZ289A3trYX1hjYVMPcv8iJL1O7XH6Qx9eR66nC/4o
HZKXB2JzY2cG8AG6C36xdK2QJNe6BuCw4JScnugh2EzGLPgjYgdkwTkNyA/CTr6F
3oKKDHFAVIjjuuyZ1oaG9DhUo7dA9SLpYenQ1YTTfOP3KbpeWgeXR1saSH7jKaVn
sww25y0gsA1FJagPsrG5Quoz1+QnqvmrJSdSJXP7uaHF8WUXe1Tj11q0OcEckSc9
GPcKgJBI2LGZQudXrhFn3h2KiVSzsg6dR8imeAwalUnwtWpt3HUdcU+syZSo0hBW
nE23IApuYx/UOFrRhEOTMasSG8hv4z9KziGTJoEkN22a9CBad5PQS1mINmtgMRkl
feiapNi/u2x3MoGP/luYVEFoAXAnLxS0aQ/1GFeo/vJnzL8qkGfvMLL1dAzwrYS+
OZZ4JqddtT0hPuh9BG75vjC1Tbcruxj+7K2wPjZ67uNdcESv8WziNHhBhvz6OkZF
OGnauvUMQBjDsAGchdUOk/CNgGzi5J1fCOk+Yp3wU8LTpE/P68ON3T/GIMxI59Rm
Kc0bKNEJpzzCCZw+CSAZC55BBFt6nyF4zM0Q9slqupaqB8qGo7r9OMBIvuwIgTCL
sN9XqSdZy7q+EQvbDFMAcpcBVjR8rurQ0CQ8xL8/HOlNZT0anC+FbeE3I7cLskO3
XODkoDD4WY417PEhvHtd80y1v8mruZGOU2okITTirh7SRNogtD5MxDMbk4Mk9ZKg
GGblAwFVmsgu+SEhIE+j/PqD2NGiCZGLpRI0Lkw5MAbEE4yzsSfH2beCPNIf9N5Y
fldW7qH20os1PGTPnvxBJjli+X/Ko3Snkx2pjiU6ZLp1T0xV4geA5ADChA38iVXa
iVj+38qY+A17gdHz/9OILGZg+Ecj9IcY3qeceTYOrG/91Gwg+oBs1c8IvhS2b/kw
9w9umnTDOUYh5gFN30WyAQQgB9rzRr8MDUiHNGOj1rwbSpfhxiStl+3suy85oKc+
nYdHjnRaO0vaCuGHXc1yyF4Z/EWUa81hSbonxTBmQk8gOzFhUi4BB4fUlz4wdNQ8
YCllFEdlh9v9+DwmNInJwmNFuDPCODnQ2qhv9xhgMLc5Rv0NxRo6ccRgpP88sUjo
/pOC/x/Z8P72L7JnJJ+Ow/lcneWM+fyfi8Puj5FEpWVjGemD+FkBdozUGeNdes5l
9e8AF1fq99eqB9ZnHE14zamRM1Y92Z2nA0cEOQKTTTdbbOLcYXRcWVUVqNvpHOC0
Kw0/XGqPOZj3rHL2wdz6uGRs6qVifNEiQ5+0i+GznQbygO18rhS2kYLEP+OBnV/I
g058vQ4XkizGMHIJ4EBwcvWneyJgGBi0TRUSARMWvIbhfXRLzbcNQ0acj1rFnxas
a/Td+UIgv65pt0YdcpcUmDrmcgvBg6nOCJqxxI27P9CaIh8OwkVEwpU817HBAfyK
+Ax1CeyX0sHzWujcqhdFzZ2XnT2TLx1hpGP/tu3DurXzAzgHCf9V09aLOueD72bF
zotE2mQUeW05qrqTOVdK4EvR5AnjA3tgvGZr444YHZPxzpfhn9Yt0E3zOXLMgBrX
XqZfr6dj+sqyvRouJ6HNFQlsFlnvJvvpFXvazAbZyBqbJQJyLcWbcKLLXkook5WF
C18Bmrn4L3yZOeI0XSrL4nArHjtfCddVD5jY62wQiFu0gRu+TyyDqC0rAulvfi22
ZjL4exGkPzaubku+GBMbt80PsaeEpkORRzGFxElLAobg+Qs2wypnuZdz7jQotcmW
h+x4ithM4d2nmN7urMQPSCAEc5o++xyuokXLERnoq3uauFa49bCNlpW5mUZGwpwb
QDDaDbXqQSulmlCxx2sQm+dviGdQQAXAl2Vqsj7AMsfM3UgKxL5HaIW0C7YJCYVe
NauECAuwcNHc0/WJuxaA2WQ7xUKG7nh4EnjgERy6H5hG5L+kXetm2ZwzeHugnQrU
0cEs59LjTLY1lwsW+xOa5yxS5vbxhwJB1Fb7utRB/89RrL4O6QUd+1MPU1C6zgcy
1W7Bg8f0z5wzk2EV9OnJ8idYM4io0waqCgTWmKKeJ/RdF2kCVdtyj9ogEYKqlPgJ
1z4m7HPbYcVlvqL0opB4p05FUsDVWFnsiYy2HLl7BLMrvk4kXjWqO/f6EBo7yXoE
3d7ow7657DO0RXjG9iIO7iedrB4h0tjQBFYVG1BdMr/2nE42aarom7oE+jaLWFPN
jj98JjfSGc3ZNKKqiHhSTmERF7vMCVVr39L2qqHh0s8HkFLFjV0mbBPTLBpSpoor
1NovL9EfCNrW5kUm6nC9RpMfU6jhs9rER5hiokZwS9xiIqtOCU75/PvLlUYKbqcQ
KYu+BbYxxWjpyjvzkZUFiJ7Wa2tQoPwPs7jGVY5D4OyUyXzr1Kw3HeWczzX226YU
430QbRl5j/tPf00uGcfQWdUxjIy75mP+oWBPUE2erCN5iI2ALKv8xNhrZ+0yyG+i
/kUt8ZsTcf6Ji0Myk1QpfS/P0OTxRESCdkWAB644i8PhHzznktuJDfZotlMsTBVP
w6mLzoAQG5q1d5kWg9nt+/WHTewNLiwiXFGqdPvsZsU1AmJrywCBss0oKKo734EH
fRwcy+yStyOH/Y05z7FpBX3rQzxM3THcVgaz69mH8Tsbao/AdliuX9mJWlZVHMYw
nb97qUK+M3l6NnTwHRwJ8Tko/BrbOM1iUvHtEwPLoc+ZffOvGEU0caAtts6wShgV
m4l3b/G27MVCc450ajDU+JdHLTEVHbQrYIOKqzI6xN0xP3Dfk9r+8cTLO32S9ljt
owvcLVk3RziuLC8AyvpmF9k2XuGd0UymG19GdOSP8+1JSHxtnvKsqLlAVHzxoujk
hJK1VBO2PyefIvI1YsZ746m+vhxBeJzjBf9947tWDpq14YzG7g1fLAKzDeznRjuH
lnvm6CSBSWn97DPiQamt9RVVLnAD751UmvHbZVb7WnA86XVM/k/ePWfAwH2eIW12
xiGe4zK4wOcLJeX5w6bpdRBbxPJtky2QtxDPbsa/6beYOdIlJZRULPwWx2WJCqP9
eptTYmVNSEdFfLgxrljFXqWPAPpLxAwR5uCw8Nq+Ihujcp+dXeJP0yDCOCilSzrd
JeobMdh6DXVHYMo0i0e8KUV2zfKQnpmbCXQI+ZyK2pLSQt8C/tV1rtIem/RyxDrn
EyUzd2h+GS8wPrzSOXUJVad0iXhPDBItkWod7NRsauCGGej7ujLBEsI3iHQY/VUc
fta0wOe1MsZ2bRKplBSNlz5UOwLB+YNorJEuSJS/6lyvxsooxfyM85TNtxJFItAv
kEj/JRmYNRptLvE7XpKy79IiiXuXlOP7pXEWRNpCD7nJUA7t3gy5Kt3MJi/oFtho
IWnHiMpKDo3xYTCG7Z+kePty05WTF0K3LO4NmE0odFPIEzDKFI3PwDcqwihGD8qN
Gt8arleLIDYBH+0QgpzmfP19N+W0/HtldzABPj6s/TplBvcF4uITeyRv9B2KcOLx
9N/Z/TYBvaY9zH4zSSerKIP/T8Px2vwQL6ELCk7ALGCbKmQqJlQdUq8n7MEG5sob
lfvumg2YEzR5N4x3ZmUbscLl2RYGJNOoQKo93JL9/f41UvLZ+P22B4gMoFstsJMm
0hERwjTBDmZaIq5qvtfAsDEZGLSpcq2EANnWLAnyhyi5vlZbbSthtERot65dOvb9
046jWPWePVnq7nGn/UkwJJKXyNKt57VuRzEtOI/HM3qQQEEGVJpjvKtsOER1oF2u
TnOpyFxQJFcJWaXeYQCyo3JxSSCgIuWaRt3+dQ0Cvy3ZIto9mGp4YwYU3Dm01B4J
FRmOEgdVaWCNgBnrzbhz4yaQOclVsHy+CjIogIg3fWtzO90Sfeup0yx3U/8zCM2d
6N2R5R+m60GJKaXuUvXhQhIRwiZqWhS/eTbx6uxuBQmvqdLb+tGULSRqM41/6E7D
qwNDCMmYQ8son9R4E/gCB1JISzs9ITtFl728nWug+Sgbw3O/CYamb/oOjSuwbvoS
jNS1gaPY8m+niS6pvfxf/3YLfU9vLzI7HlvZftTZ6eKk6rjsfDIAZL3GZj4FIHka
8c+tDRX7EAGUsGYqaideIVJY1urO04WtCP2Ton2W/dDYsY2jHGULxrt8yJ9LVUJ3
nb0Zy9tzg9GR7RMFr4DSh7sNrHn+t0cvkGJWgUIMVc7KBNqQQ0rqOVJuzlO8L4VK
bHYtb48fiYLJtCF4jtgMij89dyWjSx5xKRGnkYA2UxYpUyZkmvugBM1mHvs6463b
WD3O00OD5RpTIjN5TECbx1QBbfGuMqVsvW9SpmHyyMCg5C4k2PsEjbyvWzAW7hHz
1TCZ0pCIjikd2r17Lx8p/a7K+mZjyr5IEqc0T3G1M6CxUAnfu61AAVgSIz2NOpLA
w3zTxWuFXHjKbRT0tSN54TwV+c39qWBcXPJA0pkbibkA9O0HfgCtzWR9PIcs4nsG
d/JJNe3oWDit36JiorOVs3TaCjQRUomDNBKYgc6xBZ6HFnjmvoMYVkYIbhAaMrq1
RhwnSBCnExsXihibpycut08ay31lYx84x66ofPTI1CQG6nwKPmp6LZG4CO2HvFGQ
xT6QtuHp90uV4hc9BFyehDbSZkJa1rPMsoT00X7kgSatRHQ1Z6Zpbb4+JsuufQn8
Sa3MR88Hi151wmUO4EmW/DhY1MnXkFiwayW2WkrFCpSH7IKidZqbhBUIOjknTXEH
hJ/5ljoIvd72W3KyXTjRK3FfdMJu3nllTLhu9bXJ5NBGHkPoS8UDxp5OOgyAgFd5
RuRA+OmzeetQwEb4Cxe1GHkF1OylRr9n0PNpG+HZDA1ZEXi+66v/Mz3NwBEoH+zp
JXCre4Ux89A9zkJ6oXtQBhtSApuEtRiMo/dI0huN0NknJf47Id6a9BCHjRXANADF
A4DU/FepXfh2J6X18dtLUwMotj7GT8hctH9MVDxiMUIisW2iUNMrnm/KVnuIYSta
24fQLp6sGtdQ1Ezb3He6NLblqY8DAdAg0KHM39axA3PZFWDvhudP9KgTQ3E07wsm
03duQe70V+cNf570t/c5W1V67cUWPt43dMVBN1RVVIDjMUym7wiyZ9PidBmrk8Ye
EB6kSMABJc6s/cLLX7kOjaaQFnVNE9yLBiBD+WkpFMaFtWMI3bXhsxmWJO5v09eD
4k0LFAtDDU6UTW248ODoDXOeT3XAFsJRVbbdDlNryiTDyD7Xw6iEB8B88sxyT1zr
iOLnBcR+bOslYaiQ8Kp+tzDyQn96LHprS1LXCcO6nlGMUv0aeFBPVI5R/VxsqgNT
UwoiFMvXuWv6chPftpPGQzA1OuTUXUXho5TAza4FLsuVFfNdF3/AxUUAqOCX4szs
ZlEg2sqpaXiukyY1Iy1MasE2WDuSGn1Rnsi15nugGMKudkJ6E9MNyYGo5QuCn8U5
IjkYryQb4tnHCBEj56tkW4PgHMbbcWj3f+X8p0N33WuPX/BQ1i08hthC/dwZQjMX
8A1h3M9rxHovIfTEIvULOX6flYxHChkihVAKjVb+q6eNVKEsRS3LvcsAQRHl28jc
tfZr9wkfNz7FG96PnnT8on+cdwZwj/7Nk3WCSoe6KYMq81QASCm5+vTOSKWUoh8D
32phiGulnOvvykqHY6sC7i2GyA6gn7s4DeLhah9tLA8XzRFVB8JCQ0AE5Vgrk8h9
ZZz7vp8XNLQNVWqjN9zYmg9xDHUX3xhijR+DAO2kXLhxXO9/fV2zEaakefoPvAFg
v4n21pg9PvlzEOAOGgKw2ulJP8okLLgnDscs07trRxKvywMIaLuxYT/4IUeM9vgu
ddI+Bc5rnpM3gm+VUfqu1lNl8ZhdFvpJYKX3vNC67r7M5iFEzUMaOhrFW17GFCWh
hHm2nBCZGFr+cH1KJAoEDk7VM9TkOtrZDULpM7MVjdzis9qZxA1A4hXwl3av9OsZ
4ASOWQ/0tc5Wp9uwHEd19TVnShTU6T6jTGDjFpsaDXarRT41v8O9y4lbvyqtTKT2
WFtgUMnCjnnkEHpuEN+OYosNnefyFn87roIa7rM9zXjqaygWSWMcXExuMMrf7QyC
kW2suxRzS2Pg5g1uU+6WOVIcwPi719oedIV9fpUXgUnKGX5mKViLpRuvIml7A+Ek
QeuRXuvDbxt+6x/rSiSeV8VGNB8z4NG/DAnWumUZJVFDMXo4wt1OyXZS+Vkm0igV
wMgaFKgYe9mfhJv1UEb5YS2lnm9aWLc45f/tHbquPQPEX0qh8lOzLKW9zbFN62oQ
Elv5G3lufGk6jW9SGfTvyUq+vYWEQAEJMF1aPwiVDLtSOit93aj8gwI2E/AoF000
Vh13ZVhxFJSQWaEy/lOL585FtNRt9amWy/hrsgAcXSoCCk/jlH6x+iLW3tPf2syd
uAv7epkjGrnM0ky2RSFNstRW/lAL5CDlr5YhMe9wLzfJX/jsIpa2lY5+6O79Tnz5
O7D6EETduhwVp/zdIx0a65hQuOQg/bEFWy9H3JHNBaqq82SdtHUlZq94EsZB0CPn
3qAQkIROA2Q/iP4oCTDn8bSUFxZuIZyT+a55fxT4zTwitwZnLzjvvxmVDbKIfFLZ
ibNyymgBwVS5VvyxxqGfqJhame+6NgDaB743n7+AvrlmMliKOFntWTah4Atthmqk
VI8SuDiDbhd5mOBCr1lNCzzK5v4exVlym1KgzylvhoDIN+gnIqSmAgfJJEnax7fZ
HEIRkIP27ZKAlOzFLgbD8Dkm19snSbCO4+7WeXXogXhvBEinmPP0ahMAG+2E8d0Q
GMx72h0ZuE0oalk1w0i4gpp0Qfm5Swtjx8GZxRun0X9JMtJwtLJmlk1smS+cDe01
6fcyJMGGXpGkgkoMEM8caeKket1gwNYvldDP3XvHWb3iIelKpumXzSgjltwEbeqw
vR4usRx7uQXQ9j/h4gqc+6nvUjPj6cKM5KIlQeN8vXygXsIestKbgiuxkiOnMEkO
dMP7BcLZoA08MZYnw6wYPZ6PMhlnHnin5crALWytox4oc74kFBlUIeo3+eRkMy6U
qpOK/Lz5zoxI11AXivoeUjYqMDGR4E/GvaiJlwB2EWDa5sYKJlLNJ1TXowZ4Haj/
f8RLg6C+pM8juQ7EkJfFLGogxJrR0L/T+dAk6UY417DUoof1GzJ6BKwrvOXS7iBl
FP5AQolVM/LQ75dAj5ISziC6/saBEAUWxJO4D1HzPkuRjqlMlHyf7jatJbovniB3
ceRzTHgqKtGIF1AlHyy9lrKfWYOZGuuHbwh/BkWrot25E//Uk6tj7xd1nxsH2LFK
GQt0Kz2VoC1S6e3P7+FLh89VgTqcdWVeD29QIzGMfBOZeY5pyECJ7OTQybjW4uBT
0iAqIuqC4vYot/2XtgGUDuUGRxFzfKkJBnKocI8wcAbDoA2nkYQsNhRK/zydDsYg
KJb6Q0usVry/qk63FezRRHEATw0u0T8E4YYv+9qO7maRxqpg4jpt8mwm1n+hOvES
Qx+bUtp65jsa3cLvwdRPOgXe2BKoaM/yLUTwRCIxcpghQ7StDYfGZhK6DSclncBw
CgovcVAfY51DFXBsQtMYeCSVgMnjYoT1S5e7RpgfiPk1+tzOrPgu3t/KF6l09B5p
fLqhpMdWzDlLx+GWhjVawKEi/R7XpXbNS9h55jh+Atk2HYvQkx/O6GMj1QJJE4MC
SFZ+Dz2SVD2VGXavcreHD+TSWW8ehtJLhtWZ1oGnEr1JBdMAUvIcfwxAkSVy3PNy
6VfrnnWsOaA/DkSaKGYtIUeU6m96cO2xv1MZMyFiDsQa/Be8sUs4vMnhwlg3EcYP
LG95GxStVTyjWpesNMF17TqXV+WrnIkEJCC/TO1YEf2vIIfQVRE6qA3Un5JuM0P1
Lae85yxm8d2yB6DY1sCCbr1HBnkzQ8qmJnC6NBAIX933AQDjtPU9QmgEDbz8uvOg
Zfqq/oF8VnLlUcvZuN/dzvNE165XNbGk47k+83EdKxypUxvRK4ghSt+s3UcxLUpO
fjO1n+pRF5p05dvAVVbnTVlbsR9WgZn82tzArkvEM1KGL/APi8wOWs4oh95dNuFG
FDRWrBtCWZrRdrxv7PgMDcqr1tnZT8DxOUOFQJA9ME8h6FT/9zCILpwG95dt7ZBw
uTcGhJU79nTGcC9TMwWzCBIRflBE1CABzI8lSYYfU4xwSVSpnD1wsucjseXQABow
xNtp6c6KaVXcaM24ziAIvXuE4Jzig5Qgpha2w8XiHPoXZYg/5eSQ8kP+I/9zCpRz
Lmn7cxNb7h7uW5hCt+LTsioMo8UD3/dQvQ9hE43hmOHWsLq3pfn7hDxjTzFHxib7
fcdUiElo7qO+ErLvSSLP6LKK1rV+kQ3Q8ji0DZX0nY+QLBBCkaGTQnWhtlppclS3
+9TO/zrYPS9Nc7+InK45b5EfGVCRcHV22U0dn+JJUz3AK5oZXqeFm31VQZKNilgq
/4jcAbRTQPPf+wQSvor1iteQMg6WQT5R4J0KuW4JKmR0hwrksthcQzFBT2wfCX6m
P4sTZy3mXQr/Yi9csyv0TUsg3WHkpJ9xFcAftBsrQEXb38oA6bypZC7rwk0QwYP8
+WD8LcgIKLtwewiDz8zeEmWJyPp2Q8vhAaN4fefS7abv89OXsWYWhR/Y6SDtpRwt
bVsE2fJWfJxOQIlzelNN3sRapZn6+FsI/WHPqOG30XtIdopurPltguF0sOCIXZEq
V4i1/5hINEjHxvqBByi7n8AdnBHTRLQybCUkOHSH0LzW2gXknfszwJMoD7xJ8aJR
m8HAUvmEBcymtGKG6H+rcVAixKdWKLa4B80waEyXUSamezSDVDtYKt94m6N4fv5E
NCLV3/ff91f2htERPTwHXjFFSyaf/NV65YSwy/2AyrJ39vYWQ8YF8S0T9r9IxIkl
kgKQWM7Iaf0xghaQ1CFL1C4UlTGM+28nGDVacmZXIqU7ecggfi/Vvb6fARLLnmKW
ZgnYp9P5VJMRVCzACZYJdTftadeC5v101znljtI/57E1UI9I1Ls96v3hcP4ruQNi
kJUKGaoYO9eF51Jp06AC5Fo0XuNtJwRlRqe5icQ7vgFlfDEYFetZIyV7P9oLRjlv
dnBWEoZgTSx+0pVmQgyot4sk5pnjNa4NHxlpqeHjRnZh5I28rGrEnqXc6usnmJQ0
eZQVVRqhVeQPpGoX4gAT6llj6G2ZGnEQz9EVCQJyHaNv9NYZMmKgvX+VrKD3bRwx
oJZAhthxn1Bz7xgU7zx07G2avKKviHar8I/7moGG5pIcZ41nrEXtsTJiKc/RjHXv
jyTOh4qTjbB/W6G5wMpF3dXHiGGTSAMtIOTM3UpNy2cWjqU+BWennIzFzpAk31ww
S8fdq/8bjiQoiIMQhZ7EFEUh0uHYFJepGA7E7G2fkfG43jloMNH/RaqiSk6WaKeL
xCq4iSXBmFkraeTEspOu4AJh+0w3tIAnEH4REULWnmCYZelWrsWhaZydWfZr5TIB
gwO+86KLdCsMIHAHviptT6owSfm7SYNVbEqAkqa84tqA7vjIvd8jRWLDF3aP9ri3
GG7VpWmCwfRoFGd241dstLbksf6a1Lv9cdoavWs9nLxVEHGes3DsThU5W419ciUx
a3G9EefM5rkABHQjJqbYkrzl5iV7yfXI61kQZ8e0ZSA3UDe8vjPRNkjye0PnaSiJ
2PWM9J6QBBp7p1CwOvaX96M2VRzEe6zeOASzbxLc32Q/9lkGcYgrfTadf+x2K8zc
amlftCyAT0vhE3+LAL69wCE9H/n9WeKDCzDXWTYVpHezq2MxNAMetN+R310CL8cT
hDSPYis//oAGG+XE2UfL5Iq6Bv2aebDN0Bj0dw6bwrpkAOtqrWXmW5Yxc5ZY24+N
tWPF5iUTniZ2Ql2fiu0ZLmn5MC4yveJtHrF1vfzpmuktgbBIKLi7l3g+dr16fpm9
boclKFFteWaZEoF5uAd+Vk4rQBZyaJlXmze96b8mC6BLXhCF34RGA4ABTy1Wl5tF
cssPgPY45a1eqvwRQSp10QmquGDnKL8aEY5uH0uZuducWuhmU6oigOcCfKY8O9a0
8qqDyakYf1CDEglOyXRirjVvNSUHONVBX2Qnm0m5Yc+/B8vJZ5fC9uzXaLu29t+2
uTmn0ap4nCAHkCsGvQAaby/RhZrR41kTvoKecgId3Zu3ryUkIKdJ5m3jnUcXOGol
mMcVAOHYsk48cfh/9s2O6BjdE8JDP72tTtnWbk1OyZu82vIJBBCqQf5i0wHl2nY/
ZAhrcGkfgmGMT/QhHOUq2QsJJe/Faqq9bZtouUH8+VjAkw2wNj9rmcXSNEHNKcQ9
5A8X0wsBBVldiUF1feayKL4oraYzwmVESPKwgWThB78YYQg+E17MAGXT0VlW5bNE
Eozb74PSPLEZTXxtS64X0JIj6UCtQmCQmwmxIgCKd4GeNcqLx+EuKmDk79pwvBvn
ROoPmlzpd2DeclzpiVmcSnRTUxcVXZBeFBccMpQd0X2MsNyecouUHw0bXkn88jhT
jXoxJ7u2R9oKtjK0Nw7gQIpmmMr7aaYVS6Inx1JAh4XX/kOFAsiXfozV030h68hB
GXNukIP+n2WXKEe7adLqudQhOWG4OaIIQUdvEUTVBn8Bbvp9buwvwC+OvKs/87zN
H08j6VoCmAHFMvQ4NbHZS8tOLu5mJqMEUGxwFZH1hO1jZ+6EmDSG9TRzv6+NouHE
SM0hdXVvXhoVPpHxY6gGdHTxdE0cldsoNGsyT2v5dFA45ps0+IzsZe8/gKiCmXIf
cATQ0VZ6GzvLdRGapTkDP0PD+22WG0RsUmTwNfGi/Kqc66kM5gsf7ca+SE8WU2kw
x/o4K2FRBFlAVTf7mgVydGl5PyKMgHfzQ1mPwvuuwfmq52WoIpgZjecJ/oZsP0C7
c2URcfccnb9U+xYrGXj9jy7ppTdqHU1ODvByl+1jjHY7CEW2e+tDLwxn8694ffLI
d2dhXnysleMPpJhh34g2LLsWeCuz8oXg2zfcJ6URnTraloSq/RZJdy50T2lp1Epp
+xy2hC6bY9ymubychwN5qlK8ii0Dd5dLpBKMyIgolGlJETUgumxz0S2tEDOq7r6h
uiOtWdou64NjhESLHr39SS4Qh9xFt49z3gBHWKreyC0dK9S7QMjP6sMFDGyUSK0l
22BnR6kcUon718PEXqNAu+C6T17PkWI6vByuCJYpixKmIBt9lVp3QVDZEbxPyMEh
yrirM+RVtyeO8b9ELbGE2phjWp3fVJHYFMPP7Q0v2W2Wnb6p0PJ49uFBGqj7uT3Q
PMQMi0zKm3IXUf0V7VWeL/ig9sfPk9g534t/nNlNWUEc55yygA0k3LqmTqdXTfKs
gswsi5p2Ph3Kl+6kkbEx81saXzYAa54z4hP2jcHRImvnrU0ZJfADntawZOzmkD56
VDts8r98AFnAXM4yg67ptMpiZZOe1Z3M/kNEaLsSMjhgu3nbikVeNlm5uInaM7R6
CrVegPRVpoMkuoELz6ztc258uSVZr73pAsg/GGAU7Vo351PCjtoTRHI9F33vq8Q3
Mju+eky4671cCTUFdHSrw/V9T6H/NmJhS/Da/XVHHLsalhaC2S3pQxpkZLKJvBPZ
pCBsVbZe31s14Ud1ZjX8Z1iomSDWiP+fjbGWeKnnZIoRaARH1HF+8jyCXJLeZTLM
mqEPazTjs4HX7o/PBDyYkQ0/DReR+Fv+2Nt/12//28xhrq+QM8CuVnQbTb2o9esw
uYJArR7BhB3dFy/+sTt5AbCEnf3If3b5XA/KY2FkpX5COUaLc2xylUEEE3D3NrwW
iCFKKDsXDi9BUaDADtnveCadMIH/+rnk2K51jkffJkv1wwjngw1c/bThjmo90+/7
Tl7xtBpfZvf5tveWYqrfG1EcRVXwo4BigOLEWsaM0cESWZZN5uwtQ07nLNtY61kx
/ekKXSzg+bIJfOec9odVe8lEfAx3oc5CyHOd45leKCjoKKsW0NyTFLTAdqovAmfi
1SF1t//nq3FPaPJ3Y6PaVogIAB2zjyYIz3pC9Z6gMOIZ2xdzm+7O+jJ31jsQDn+d
XCkglxfa7sYZ+9RG3TJ0tAENQcLZUO+7VGERE2cC7AO6L7qXfF3e+19JU+UIw/Z4
e1JgTOpFNJh9suIbRNYoC3b4jTkfDVpR4bfHVbcvTrAnnR9OAFXDFGwMSdgzO0+/
ZSGYrr4sZ4o8UehaadGpebh9glNiXfklIeTS4wYnMS2JZVuBZcZVTehDt5dHz1Lu
wgqZepIIiUGGreOTfO+yC8hO1729y7zae72j0j/0G9nbsDfvWZWH80Y0Vo8j3Lag
xO7C6L3Hodr8npALcHEU76Wy4vjyC18nL82QpSmp5E4FsXls1ORLX1KGvAHCgbcP
ePhcOxLbazoTbiw/X6beFLtAvtQuo3xjLnL3+lndOKR5arCK+uDF/tFwZl5xKIhr
2B6nFeHscs8ad52fDcMGdPIoESit8I+ZVfrSzG9jmG8dWKYvw0L+yFspSMhvD+C5
QURR+ajQ9V9weYEK2uo5x1pNVec0Uw5z3pULcKejjcskr8a/70gwOeUfaKdxUh8Q
JNM/8gWtFG6gNGzXy1qEupJYQI4QWEV+2mFmsAIxkdxY5pWka9gNlsWvKPLCfW3e
IzA0QFC9BqyvZypCET7rO1RSqgY01dYfD47UKxTFWgvxlpT3KK7tvCRjxBpjYtZa
AJSVthZh4CP0jx8Jel6dfeDYKYDVFZTZ0wrxAErLBrq2di4Tw4I4Uft2d+UHPYcg
8wYb5yvUsj+5V/1W4abRz7CdPa7qeFTG/7SeIyCrhH7fj/tTr+WhCkX8uBpPaPP6
LS62E69JQH0eK+UrwpaZI5SRFPhh1dG8+d6A05u85isuQCU0w0xSld8RdgKl1WiL
9YH0Qv/+UlxQFhstxefc9KdKTbe/9rioVm2fMJdrDvVV8qEJmfDiYWq5uJBNMRUb
RPjVYa5rN/bVqZw5mxkm5moS/D6r43E0gFlIWUgbf7Pu8SEH+d5eGcmlIhNQTrLr
YugDV06WmhTgm/usBVQfH6d0QALkhbeCOr6ihyWPieNuclSJSJmkLm+uWYToebUj
LVAQVOFfltEcpgQsW9/W0cEwKoHUI49aL5meMH/rA+UCcCHpwBfwhghQHtOfhaLh
GouhrZMEgrhcKRfWhSYruF804o8MU4IuIFkmrut9H9vlExAGf6pKQx5OG6vxtL3/
kEShvW2yQH5awXmyuw0Pm6R9tu2VVr6l+YsU1SpBr/8iPwj77DpV1X9EKmCGjeia
1/0N9+2xy5Uyaz5ZqzrYRveDBFTgOCkTKiKv69kx3fgem6iZ6K+1px+r25rRWyzJ
7bcrzpHfMuFvzBiPfeplx7KhXIS5lLznO4apUHJgepsug7UVJ8nXN+58rb+kQCVa
HuDH1XfhdztBanGtZwDZOoKH42rJD/swzmUnHReRpZFON+kbtYJZ/QLvm4BCgiJW
U8nU/y+sqfaRGfOy5pfTmJc/THyTWjB1eX0RzCkbrQg+sIJBQBYgCXWfozPojDd9
vGHdQJPvm0IR6rXSKsrO3mfnAJ2VgAP2czccO0QhLtwUoivwMNWPC7KRkw2vm3CO
fA1lo+LKS+ASEIxMgUsHajKzew6eXHh7rm14a+7/svIsoYF0kRDt2WRfFbcRfPXL
U6zev3tp88H/Gq3vQ9zs6IBRs8a2a+DdZjwem2cvCRi3SpI1OEY5QQZFS4ikLcYB
j2SsxV94OMQuIpTTZcpS6WHK1H7NLq//mXsB4wShOqAz7gnStNioxgw5LabLFoI0
nJ7NtG4PEJpkqdSXQv5vsHjq7TRrA1MkqfUoUBW6KGCZwlmUz5mycuJA/ruLkDe8
v6my5KHC8JrhyN64yYzLVqXW775jU9uEsSxFrEevq9lVAhp6gafHzUP9ERb+1cRj
54VfIf2ks1PJFLzTnDyYsMq7ZqlFZfxGGB42Ypl6AbJxk1SCCV46ddtpCvZ7+sUE
Ip21IoMT0yWtjYkApCSadIMBzjuNHzBBQDF0IEd7kW4ToxNW0h/3it6KNqqVtt/8
GbdHuVjT5IkU1UvXBYRWtVjxi8ZoHLwMbARjMsXBRXzGXnW/2LN1DbtxnerpVMKq
KaxUuVWGIlwoScAA33tvbhJlDD5ZmJGJWVsmehSyfVnkXAAZuj2brZrtyzjRD/zN
Lnfh7AN3L5ZPZ7EwuV6X6dVbveUZaP39UblIMdjeWDaJsqMowPx896ZbvAdKEkru
qJtAy3hpmiy/BP1B8RGHKkfS1g2LbIoFZzTUQFFdZJDG5YV+ERUUfTz5rWaed5WB
Apoqld/uHnAHKmmDh3XxmMTM6iV6Mirdja1pYY5E01dnmLTBTdtZLVnWQvfPJV4g
h/j7k9YSYBruiNKqgc1tLmTwdUOcLhQcNSJYIu4pQpgpDVclgdNythY8az+nx8YJ
U8uSxu/66C1e/m39irS+wgeu/+fEo5ICKUhZgmYZi/nlps9hLWJGRALT9UG1kmAb
X6ZDdbIsmpxlYDbkdMQExDqdoz4whBS0pPT8tYb6o8XD/KQlh4n0NvsklylXqV7t
Fq0Lk6oxcvWH6nOD+xhh0aKos60mmdiyN1Nig8b9XG4ipgM6LsI8j+8eT9lHEy4N
kYo44d/hdexXTp9KSc2SJMDHkXu1wg65PIvKsYdGA0v1otvL5mZGe2qrOb8Wnwv+
z30G8D5DnN3fqCkk7IxwGHs7aMa3t0b0U6eMth1Q4H3BRYEopm0ZFszn5f17Omkg
2QZD91nkmbfUqgCEZfcKHQrFoomjIXnl9t1QzxqOar+Yvml5y4QPHQ8LrExNnbDE
SeuMQav7864OwSHC6kq7bJ10O/4cCWrr0cS2g1ImYTRm1jUh9gT4xm8LwYMmorw7
rsxcwfS8feVqPJ+Sc3gIcG+EyLwpIrrZSSoxPGEofbhJMQfhbV/IFCUYuTrJhWPV
AwAd7gJ07+fQAqXRe7gwtNVN6+2L4lM1GBFm6zEFRzCT9kqdKn1Z43MBO5sqECVk
764+Yl6ZYHsXPjbRkkkuR53EAfKYAxVuTsWHKAulDEvPDy3agIyfCQCOUJfobCVc
QNVBFs6/1W90cdcGQJ5/dE4pt6WqXvdO/1H5ytkLJE4TT4r46LRQVrvJmRCLZfni
eSBYIjG3KKM/jSSNk45OSZAPGndO0nIq4VZ6PlKD2r2z0C2VFXTwJXXEc3cz0r7S
bkROZVQDE1H0tj/vo3RBlL3L8X6bmbi53bi8Eodgg2fPbH42gUiofw7ZQuOiquQN
dG3rFeNMqjkB+raf7OqzYWh1jWHWnm1BfM/dH/St+FZKJWny0zOSX52cOwD5Sahi
200/WXL5qQXcuwTkhHhHX2wCbAdLXrGpupRpoxyKy9f5vTyeV/xjxuD3qMGl7avk
XGUAppccesxXMitWZ5vJ1x1fxa1FpV8gsbqTxhHG8Js55/QYqzlArpXBrWT6DOdp
q1kmvAXg+80b4KE85cgDHowfkVFE4C7OAW21+D8soXsuZefmoKlLytmZkeVlFJH4
CZniF/v2TcTgXtd+7wybzXDA2YOQuuPkHuP7Bxr81KRMqzV1L7gfkJR3oTM7r59j
eCtAgEgTgRCPDT8lwULTYH+g2VzfwRovCP5vUQfk6BzoZfWyG425dp3bvI1o7cq5
sbWEckpfXxR94BtPl+JGQ/ZITRo6mBSwStza+ATPvy4iylf8do4iVqFPwaR8/cNQ
A7n+TACx9Y2aSWQZD0L6r6bRb9OcpRFZDJveQFlxtMCSGGD7ktX0P+QadMPljQy6
ye3udoZJK+D6JZKpxxSrmn0eagkLzFhjerii4rGMHVQmcY4lmxf4MUJo3itYTG6c
wwJxMjy7b9J2jS/srxAfjOqgF8KHf0AaRYqiPlF0xvgAoNHfE9iS9cdnSv9o7Hq0
UZlDFfvOOceDoisktGzMNmBQ5CAhD+PBOICu54HotwGm3E75mjbX3BvXXhWAkAtB
iGe1mBrELKDlEtU01TVdqKi1AoTIrCyTry6nsy70DXrQi2J5ialXMXLHlxG0RkuH
yXdKPtm/YHy3wa23NnvRIabPOojp92o2n3eU99Ivve1uGRM9I3DuLV/k5Dr+ppWd
CyIKGcvh7RMriszMv1a9qrg0u7gLuZT8RZDuI58+KB6mvO8Hwcez4IAb4B4ngsqe
w+YtHlPcpr49enNANXj77rcJL9SZxis330+qjxIslertnAw46kOD9YBbEBXqyYR0
jr4jSI70lCx+hgk3045O284Txoo0PDoIhM0VcXJW1lVbF19L8zDPHohD/H6T79sZ
xQGNoE7UffDyzbRA1hfGjSmsQ/ATihJlKFzl3/C+gTsSLa/bw5M6CXnr50KYbKLB
Wb08Xrymyw2OXxTT1cpKmEhx/Cz9uBGSkYytdq8/rqupcLjc0LWNf4SxkuXkCK9J
LlGgpZK76P1lsL6lg4o8n/22x2ZgnvOTxQ+IeaCP3kLUPDMfBhdpIXbMozj6y5IM
59G6q2Uvi3saaKtjpEy24HlEZoJkP8czE6MnsT1bQwaKRUW5EnhiaJhS4bjLTYCq
HWHX/u5ZILIrpqvIQ3aYpniWc6ek4v3bhiGy9Qn70ASDSbY8bf8X13ofY3TrQpVm
cOLX92odrHSxWTySN0hF10IVbl3GcpefnDSHwfTnL00s6jpusLFdv67n7zRsZJ6S
1c94VdyYFMrAQHL8og9tfThoBpAfhTrWtlVuYFoIjE7lAMoYhL0zHjphmdK8rd3m
XIzJ/8uRS2nX8vr6GizbXCjLSi8e4fYpR1txPm0TM7KJDGhFbzoWk7x50OUe3GWq
cdMvaYEJsfUJ2wVmMVBenx1bRaOyKCA29uI3sBCMZwU/xVzMztIQkauwB+rPDYnw
09GAIiDdH1G3kTEdFl38/kHFaz/hkP38V9ZSDwg1ZBbiQeT2yh/51lXA5YfH9RuK
Nj6QGx0p6ShCPvOOb1FS4vgeq8VZKtITkbrdyUHXp9EVvZrZ3MY/14w2+tfhMmSX
TrFPdJR2M8TL2plOCfm0V3WWzwcXLItAbtWF/lj99sXgzXhhFZZ0UWZbqUkw7qaP
9hU2vIvVMd+ljNS/g2wqPAMIZDOFtdNT4PBI3WEzoW5eVrIsWojYBPSN2i7ZX0rL
TE+hDGxaD1L+fgBEkDMg6YePrmv0arWFVNoZar/GUu5YCTsTp2Bq+WouK+vLw3s+
AQBwiA2jfExwpNk529T3/ZHnKsN2jprDxzl691cbQXGpfe+3YPyIwKDtTrDSVECI
QwF53eiko7Ivf5TKCbnaz1JcC82tfrxBTuIps0Ze28vN4YCLuBb8gnCErV5p3raZ
5qBor4j8x3dZcLyo67LPafdHq6A3MZ4pKXJgVQCx2IssoVsalXK0yaKzzqXqV+Ou
zVPxSRJ9LBWpEFfghIjOverDvI6dQl1nBJrebr3EIxNQ75SXFJajarmubyJ4lI9f
Dr51BP+FQC0MDgqRER5B5mmhvUg3MNx1pe9epNv6AYE7JkRkEt6p0aMVk/C7SeYN
v/fzX0zUj9zgQ/ounWifBg71n+AQl1Qiuq3/x1VtrQB+b0m50ZchMq/4qwsw2mIt
Jk0yFPO2nMmRMqawxVEsSDMFWOJJFRLqwhTx9/ZnW1UcBzWVj2aVwMKvw70fs9Zx
AlTL8VzUl5nEX0rgst6i2WJ9BIZsG0p69JC9NbkOmWG6f+IVQ4/TjvJXg3kPm5Uc
xlOODkdVlA/upqgL3/gN82ACu2g7LBSixRSKNghEbzxgwVVeJcfOKstJY9shh+TW
SGi/Yi6qfhQ/zFqwL/bQ3iPWt5uUUrjrdsIDEzFZBlBcH9OJC3IfKLt5/D+riiJR
NddPHmZIWxx/GZoxZNApApURuZj7w/TXFyWEFiBQus/MaOyH0qa1z0/tYWMev7/X
4gGGw5ugcUXWW69wJVBvE0X65HA5290yhwb2vrJ8jJfFhypap6OsZnH6Hfx+QLqp
8iM7WdpUqJ/7lR+cMU9m3ioqVxKb7cCpKfhSmL7GBHUwpQvnVXwyz3tmrYNt16fs
aXNSwcJRF5eQyoo0g4p4Vlhn8ZIZkjcRGsYoh+pVvJd4LuiCowlzFTBgAAkcRg29
3qzXzqWFM8zMzma2M6GKX8uhvxOWwFnMrjvRPpj+t/VSGx3yn3kJnf+3Lia2QNEG
TwxxCaWZbWY0HttI9PzAHktfJAZux++hjsHV1weCBwfaRx9Kw/jXwzvyn0xOe2yr
HjvPAJtKwkDd2RmmwGDDbbjg+EMfidV63lbX2GZrwrYPvg9Zc1HMSk+tM6SGoF6Y
SSsN50wLNnxWDxSJajo1MKsDf3HmAR5JL8HoVPyzSHeFzc7OfdX911Mu78T+d6Gi
AAi60pJJRSVPYWT9A7aYnSCnPu0qAkSpPoL3TTZwwwDTlU+7a+J17v+9FaDZziNP
Y9jUMzWKTMwcRSuFnLZAQd81EGgxpqk82dPMCgOsoAhJFusgZJROX5JvJOmTf+94
tuvJBD2hUuZbsSHNXvujT/sSa0YzBzBuRdTcJBWZGQF5eBdkR7Vn0kSgBcqLBuX2
ZYAghN4RKdivob4DLXBB9X741xjW2F9jPhi9k4sQm42ogIdbmhJliTxS7UwIig1t
aLMJ/z3HpnXry5GF3iGpumXKtF93uTDRqBdNRncte4/0KWEj7sB4PADhHUy3LHm9
EzOVYQYQUvWPlrLEMJFp4A+lZEcfKFwbZ04vVQuurPLE4bcCrOAv/hZNvvqg3VTV
QqAAgHavSHOtb0X16PZwi7POXIVaGAm6etUSZIODZnsPbbKrrq7RFFJTFJd5s03T
Bfit6wWQSMPKHAIILyn9ryw7qN4e41XHqjTsaAqhTItoLjAEeWGOaev/jCCiy6QU
Nw0s5jYsZjiytKS6igTACpRVeqTL6YHU7ynQJpK3UGhPrt52Vygd211SM9DAkH4o
HQqnjCGpLE61X3xO0LGYiRwUxj4xHwrkb8+O6J2XRX/b3qGkdNs/IY/sidB4ZVnT
myb6aA/S6xRIVu/2bOcN9KnZG39sS4VBMHaX6IRZDk38QRY1bR4dYNtC1+FqrgDa
Ize0hGGW4z0PG4Xhw9h/wnT41X6F3ILnzYkZAK5aPg8zcnzwW1A+UpZ/jWfev5iv
XYkmy/tHdEhtU3Q7ur0mJK4IHr2Uwgl9YSpqHETMOZZM/hrCEaZaRFtKpCc9jJrv
EjWUde+MhelQI1JkEzKYKs+ezpkhCiBTOF1z/6udU0o8uulPkvlv2oKTXv2noD6H
Mck54JxK83+3BfP7EswOG8t8JwbUlZEW9Qxaa9lGKrhttr0D7BZjKSRWtANINfmy
UJ4kKB9zvEhc4xazST3KQEUhhcsIqiLJ4jz5sXDX5ENGSa0t9j1Kf8PDnYUqQiH1
dxBPvXd6jLm5SPB9DeHlZgH0+rQMW6X/iy4z1GIz0IzB5+unRyId+F4fzmDCnyjp
nE7jQf7RCLE0aLKpU2WAgvMd3EqgNrujSqmQacuJP7sZJ8U6huJxa5LMCsSoIx0z
1st2TUK1cg/5naFVgsb1g9FWVKbDJnqINxKkEEzg/1k3u0dWq4WYjsMwPvGmlW/T
k+18d/wI9vftXWl4Q/N5p2AEdN0rMRsba+5kC1pab5U2SNCUG6mbRqq+eJkX7Fo+
6Iup9iL4G4BQjx74QaR5KZES/Dn1HoR3LQcpWbxgT692w6lUbRImwo5/D5+YOqN2
T0hXWZFM7CPQ3RQ3lVv21tSLcVNetlkO1aSzKGlcTX2JZWolBu6vmiK3IxhyLH8f
639MxfBB9YuqxoQIYNXxdjq21zI6Dw/cUe8Ancn+12JnFGbRf4jJuzpuiT0Gs6tD
+ImO1ba/drQUwYO62IK9ZcN0wn3QD2dV3Whm9ojo8kB+0SC0q+HseRf6z5fs2srG
w84qPFWRMNUPFXZmXdaSAQk1LUqr+flmauzFmc3KEIZJ9RyXOdNsG2Nu3Ux73Rga
Kqm29awX6iAH58USmBVvspa19vbCMot4+aAJZK9z0BsABYadT4uFvkgLh9/9TzO/
t40HkWUnnAqEtXyRrEEzhQp1jp17rdlEifi3oTTefqqC1KDpjCs2VhlF5xcR6IAk
ul20yt4xvmJHBtQ0Bec/QViw/su1lR1uoYHZrgACPtZQNbuEQsFFDK3qH4zh/qLX
gX5vDrEtE/vhaD6/0x5GIF1GopfXOUAQ/LtlbpQfVa3pYVaWZ8DMJPd9KIEARoco
qvRHQv/sNwz+yd7upTNbjw4C3UlPUCUZaJsd6HNj+rRbgJ/IFEDhQAvbl7ZhOyi7
KLeYmJTn0/ccqEOAInR/18N+0aoZCcRSXr0cPRDPoA3RYuF/jMyj4TwMrGMNr0D2
FlDgSsMhur95AqxxoWdpaHaChMTxvLztV6cF/rJA23a7ah+7yGBGVwwMbN5dBMna
YjCtF8MuUAI+zBTK+iJc1FaCj1SRYG1vcmrjJjcKEjhYRKV6xUSPfInq1VGAcWP/
Pc0Kq/K8akcH+1BtvdGWi25NvoakrhwJCninF3HSing4HjkhSHXxu9oxGDAISxPC
Bv+PIyb3KOvtuLuyFRJxe5Yley/I6LOjsdPVYrCK/wfdL8cPhuz4tlx+xHfGR1d9
LoG58JvsR8m1YRDa3/CanCYYgBGvWaC+Rdv62r/C44sQ97mypg67itaP9ZVzqzUW
EFBtFpndzz+CzeSsU8ebXQVevqCFEEWIyGSdHP2ZzXFQWiD71v6CbT2s0TaUQv7k
X3TtGutr/l0zOIF9n62GdNfsxlEp9cVbbIUmyeSrlw+o9CVU5or/7bTejC7Oy5Wa
VaypQzfOKiG55ouncjmb5zQx5Y5YXEjyfsyUqdAbjY3F9RdZpSw9IhNexXU8EAeR
VwG+g/g9AypeVdou2GsrG3BFGIPnU56a3b5myR3cTrnKhuqq2BXMKIyveqXgbfUf
k8CeL3ow0vkovfaKpR26+ZFGz4GiHRDgga1bkMQHTCihgVRe7asCsqqMf8cu83wl
jLtXb2SvM3gavyheQz0t2GAyRlJlO2YLaWiwHGkdhDzEeWhujUdhulk1fqSD8wj/
Kwc0CLdCo/6Q8sV65p3WEbctKVg7T1nBtlSMwbQLm2e0vh49c3uHVRn6CHXmdQno
qUsJyWJFBPRHvnd3e+h6dG181CIDaeHYb+kS84HI676NXHwNjdyYq2kMgECMnZFQ
HytzbUL9mdPkz+cvdLAE1HwBbWb3MgGL4tU53j75Dx5nnpOi9VHRNGU2y7JKZdLI
zVUY/1B2H9iWtd8IAtUvlxVG8k8SCR29VSVou+iN316QrbExCYGI6RxB1RxNF23C
OJDQjqnUNrzdffjmYHZFS7frUcDO3WxBtFOPUMlqtwkqs4nvBVLRqbsaH4ap2SdM
tJoNuqwbziFsiV0dzhxRCQhGIJmq2X6evcunANPpT1ddA2gUhEsFFiPutes7NKSc
CVvGXYh77gw9Hb2DxkG31L2fZbbaXtWR6wC/pujc9g8IR6HfixsIRA6nfxrwjobs
Q1QoCz08JpeBHIpRGvK3KPuKqk9RgUFGD/a8zn/TcPhrWZueXgTe+/G5fI6qpSJ+
vAU6sYuTCaCAdfjse7mZVn6gSfEX6E38Gg5HUg2CYPS3OV43LaU92sMRbLuwqyLM
vZWocnlOJRlqmjd7USxxsN4YLIsQvnIqNA82a1xCsCnV04digxL7h8K6SDRe7l1Y
s/uuu6OjET7BwEfkEYqzVjbDUSu2TKezUxR1T5DPRGc1Dk0JYoKVKEnaO89F8VcR
iBT8H0kzCS2dDS+XbhUfvUCK4hfc94jVpMDG2tdJZF2nzgMDDvtnjhjinuOgf3nW
mPbv2ikgaV23aB0pkaBiwyyfWMLL9j2AkrFUsBJRHkhG5AcIWKhDG3JOIMvhrCUM
BCojPr1BQcb38IJsnUiOrAUREopKaE3El4CWZ2oLV3AYuJ2kBENBNBtvyf9IvUJq
NT6ZJitDYwHUDgKS6gU56tmvDWCtx+o2z4UHsbCctK3R/LGAhp33497hTFKYUVjH
F54X2zHhOzlvJkQQZmkZTL6mSVwL561Mp1rSVC17AfvCO8sssEKIT4ssEhtR31Nx
VrqCY/bwbu+o8DcFuLPzZafdhEB1PM2+G/6YJAnEo+gf4OQTSWy7M2BTvE3NPJT7
9+G0WmHWNRwRylX3GJCkGiYjdcv5ldPVkAw2nUDE8v+qhiEVEjOEiN3ywEwmGGm6
3Q6oqsKuY1z21fdWK046qzTacjSHKQxL+tItBhtFDJeMTS94UFNsQWq9uFCUsUQA
yesGkyiyqBoJvmWG+Phc2FZH4GmXX2/ikW0RV0kmOKDPC1K2O3IWsBrffpaMP1JP
cpAGJdVznNkpx4MAgYkbDuQkFHfrWPQllxgJSEeyLTi2GSCbP1ykdn9pFmixdDiM
9ygdMKp36jKyXRU9F/JJmj8LcwXLk5BzuvDAH3xu45zpfuke9SKh0NGXaExTNLu2
XrfUxAfObT+JjRNyutZIWmCSCxpKb3q2GgvFLYmTNV2txBv38/IfrQMEsCET/VoP
yh5Jz59eqCXEa7gWV8b6F+4vDS8vwpoX4aefRQpFr/5F+0Vo9mGTCyyV7GdzO0bl
msYdygnH3T+oaEuX6WhMHfBzESkXdSngdVKQV9VjRbI1/Dy758QCtVrrBtzLnBzP
jS+iyLPGc+wUc+JXOjYkAfzmrg1zmguFww/qlm/wuXrLNjKhC+Z/NMvg6hg6yc0o
HJGp8tE2yNBIsEKdS/FHdksTxvxNz/aGWciNGsLDCKjzI3Oo5J8C39av9FBHIaCR
GU6ewZLH1bq1n8+NcUh6Yp1Ln1vH9d3ROnpwH4QiHK+ruqZeAXfcDzV0/6eEePTw
l+3hJyRarRZWf/jSf5bVDeuHbV/NaADEd4QYmO5KnV+A7lGOSHnNVXKJlvnm7lu7
o49Qu7znIzrsDggdoTqrE+6upuu8aLGfTrz/C4w8mZ4Gjcc8ZwPqkrqkvNGiKU0G
11LdppLVkacCmPeL6eeGTOyRiewOpFZbVu8lC/nr2lJNBZuumBG5Wje402tZMK2b
9P321LY2v1x+JClMBHQQFkNq3SxBwsC+LXtiCOg00w49dJJc6BMdv2HIyoL9qQzB
TEjFoNxDMmaqG7TuYNs9hJ2uYuHR5omCCm78g55LmFk9OuH5SVY6+z4pNttkhVp2
OqwBnU1boG2niP8J79G4/0L7D/K5LeigzsFe6Pgz2SYRr6cqbslPXUcaQRf91dQ2
YdbX+G5PWMP/piaWy0QoYpBrAzPAd5vaCI1IfgNhEPTHzWAOWl1GQRgLs4mKEvCZ
2udhSqNy9PNiH2RMhheBS84KL1OySwRHzDI6lbM3RaUiZ0CMaXQYB//Elucwt/9g
i7gnR0c9v66tqCMssqQlIoh5XVgHeX/LBiWSRXTIc1G92DezSxX4CX1pqopsUSVm
jVFRIlXzmxl8dzoCk1Qk1jY8zhXL2z1gz3xgMGSmrCgdfDlxL9b/Hznz5u08+W8B
db2tjGfX5r3LdiU6DYHdDAvckblbOJyH0wT5Tpo7MBxtmu8YjtHS1yNCPFMdQ9E2
llo4JG9RN5PecJfOfhdI5vVsg2MN9FA+nlm1ZC5XJcDEnPXVTmg5U9a6FQspwhKB
GmYEGe1xmbaT+UWojkXoAgKMcVDGIXlx6D3/dmjBVgZzyyc0hcQGc3MrULVXE3g1
BzJNyC7J58WHFNLSU6KfRcfuIxBxuz+oSGhwREO+llreLXQ7IqHTtkCRiKbsecM3
y5YK+tQvWtOCLfMFoHR4XRIWY+33ZE0HBGXo+9leXrHb50ct8UAnKjBjSgYCxP4H
yYWqIlnre98wGL8QOkLyGt4FJ/qaCare6wwbdLXlH+pusrHsln2wA4PWz+hS/jss
tew6nfHb8kJrp/eOeOxGx/p7vMzFX2+AEYMTX8SqOyx5fVoBiADBjuL5DV4EGLcB
1g975eoDhb8Uj6dX8Bg991tWowLl4XS6dpeO/O4qLDwRNP+zrW+uQOqo7RP8kTMs
BKcZQUmmHHHcRhECq0s0s4BBpeuKtJvekMqCbk6yRELB/QMBhu1VB0OmKztV2lNB
ruV/ed+EnCNWqzI16VcNAxZgX+gdlFWIFQssJArfM/ucP+zA+CLCYyq/y5oaGqRn
mmoPIwMdgR3SGVqpghJygVbGFrFsGGDl9r4RWkLb/G2AzeHBvGbj035//ELSvdNk
a/wykPTytBK7mzIAwvv5iiSKLV3uawU+S9KKtIYgjMqf5sV8gvSWUDJksMpTq9qs
1T6TdxnBRmGyKQfprak2zNLs92bmFhIl4ZxmbbfaOgCUbDKKIYf5yBCdqZMWT1Vf
m2pzrjsiPKGlypu7NqUohlEDhf1ZS+dtb5p8zM20B37BoDRiBGX/TWFVpBl+cd5x
BsHL613kpKCm9jaJbM8lPFdFhs0PsVfGmPnPW/4EFQ6x21ickyyosI7bpLcytuyp
XJl+DxULMcFyhBr2IbYdC5eS9YNEcE8bmrZ6qqWVgD1b8Qd0qoorkWz2cTXweko6
yFX7nhfpHQJxCxb1558qATI/glOUT40zEKYknio1i3mz4Wyo8Fl5jjlLKZoJCQAi
TrL0IsBoURKTng5X4Rp2K3jft0E2cn/0REzW1KC59R5+Cm8FhHbfAHS6cTOE5lZ3
meQ7J+OWQcyQYJ6lZ1GHrFN1yAHFt3VfP5KEOtgexT46/7ZL9QAhmED//aDKL95H
QAEHjob8THJ8i6rdqkbfrbEzIqo4R13Tv5RKebRvk6MPzNE4UU4hjk5rcMD093cp
UbQIEmXwmlG6IcXyuKDZNQszjNjJ4A+dtlji2/bgpdiYPusWtrDhB6nwDjhs9oP/
CkUe5bXCuplV5IbW7esKOMnqbXsFwg7HHKZZ9bJcAvFXDMhtyKoTryqlRaGW9EvK
5LZhRmZRWOdRvfBDVBPt9+lgO5Dtn3C2M1D/sdvNh9tT1PP/rTFnYVCLcxzDT84T
5x9B8ykotLNFI4TfYsZbZwYQ+5n4EpsOoeob0ltZuTKJMV0P80CKRoecexBH2Y1P
aJq9qys5VAIn6DdFwDMYuwQ4RxbpQeyy+2/2oaNu1L3z8XE9MAY2cl4srOK6/dLR
kLULdi+t11v0tk+iPJAspokhRy1M/+z+TrKZl5btqOAQIkjumSoApdzyxfI7wZek
yLpHu8hkjyOjGcsuu6bJ3U1Gd1S3fP6+e2A5baHDZxqfs1BLYL4+eYBa59oV/RG0
R1nj9bVPUoylYlgWlIIVRoEZ/kPib8NcDmIfS5qahD8/0mEx8d5cdXopEBdqax5k
d2rTObYYbcAP7JTZ8kXV0EM4A/tbObZ2W2XsgtPiVxGmEFE7B6LdrnhEOc7/VMtO
DeJNVDMwWPENOmuhTVvvo6x3Q0NkGXoZCtZrQ/W6LqNtK97NcwfgLVTzgh8i+0T5
oFtHYUJKptip2AXbMmuLUPksw//1dB2ou+QTzls1JH84W0dtsIN+gf/uQQtP4qKb
VIoIpTLQfwIEJtNyYQ6E7+w6HVLlAATUnXUHqt84dE6aYrdIz2x489rUGamCYijy
XA7+hzqyGl7yABJYqP+iQhX145HtddRdc56JskCKPhaqbY6ZdYsTc4wLwb1Fbwax
IFNsK4HflqZvI8cyweAT7+oMEi8FwctvrJ3KL2UJ5SvgZC9f9a/Yh9fJcx3JPHf4
6bdJ2mHpAsE1t/nOXgFIIPH0hbngDaLV9MpaxAcGIHRa3/iqUq61K9sBtg5Hj/9H
EouGjHAe8mhHc8eV8dNwlEwiKvmYpoLLZxSl+IOu3LLathVsVxA8SOIgsTHUQLwE
hsvFCxax2Fjm173Emk8YPTfxrRpOzVhxlfhF2LNDU0EMWVhoYDvVkN9r0vLgeWU8
RwQg4Pbnw/5xGLawDCxcJcPh0dCs0qzW962OJDXfvlrxCbf3nvG6iOLDlWjAsuwS
tgRKL3fnDj2xGBoNK6Cd57IL2DlQcOtXzhC/6mHRO9thGlfRNAC4MmXQ1QPXcCkG
QqbGF/jToXHNosaR0uaMTqbKC633WbtQnIBgTmy3XCMJbLhIex8mtnBcY67+brzo
OQ7VFhMI6kSMokbO+CvIGdoxjt1p+PY8BrarDiMKUjon+PvZRUIxiOIbSw30TCc4
`protect END_PROTECTED
