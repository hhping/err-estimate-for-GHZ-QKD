`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10Yz3MDfLkRQqtRWnbgB1os12dzLBFwIolRvUcwojUqbZbf06G/fRF9aCOvzr/8Y
wel/gTjv9nstWA4hilpp+NnxAIbf4l+kLNrM/JHyEMChcLaGmLZyvO8ZPoeWU+Is
01IwulPX5VmzHo2cVIUqDkD2fOhy0UtN2v0Uu5Gc0P8X5SRAamtNlY/4DNSbmZzW
fdN8enJkf7CEbw5YdRcENuNp7IvvtMLKEy/MnJxCT+9RTQicjd6vO0DM3Qfp4Ys1
hTFXk3A7SZM/wJijic+es00l63U4LArp6rBHP8u75kHW1+kzFoLqXcW+LyjN6ed+
`protect END_PROTECTED
