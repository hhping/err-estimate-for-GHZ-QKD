`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sh4nj9sSWULThIzS5c++xmIq30815I2iV8TTgDURJ4ttaqrRcGP41v2rySEhmqIu
xAgWkTIKUS+kFB0vuQIK3e+c1FmGxpHTG6lCOGvH2dBnr8iR6ffJoofFy3RorjIS
rZuJko4gRtx95oGuP2cP/avAhWlxjBB5ZtXIuGxBqPh4xV9Yv9EyIas0IwG0BL95
N1f9Injd00vsBpzGLiAJ8+n8ystucbLNI6jAK+9yRVOISURSKGkI+7VII2OgMWWR
IoDUThTctN8mJObTs/A6feNXAAjrtqvQ/NjzftaZTnTTEIx4kPdW06B+gAXUBva7
HnlDKMZs27PaCk0Eoq6t6hpZNRyLGbm+czDcY3NDcdOam4Vybe9mMeoD5F0Re8gD
pnWwBjJoJYKvgJYdZ/pgQIeTIq2h8pNI1k1WUaILLPzXY0wx2EiByIWu7EN7FN9v
SjShTXc0N9+KDBeeIE2jsWt1sFvtTMoHsN7XR89dSguZR47p+3moENyAYBwrk2dQ
nyS/L/nZ4XqYWvwZXzhlCdyanEQ4aeNifDg4yfNZFoUKFE9+Q6S1s5V0CsEy6G6d
/LgWQFxGRUi30na1z6P2kmRWOQk2YtBsbqK2UtURXMQyUpsoTA1VOc6yQyzey0hq
+Vfbz2koLyqmimwZCxq5XNrs2KiehMdsU5Atlbn0kylrzFdTkSG4qTU6ANVrRnAt
Vq8Zr5h+Tcz6G00/udaXCu8o+2ZZrvXFz65MgRCY9eCQoPbR7MvmvLbt9HuOuzMk
qa8UOy84RMZ2MiLMDbQpnb72JUtPpauAVbwPemKwQag=
`protect END_PROTECTED
