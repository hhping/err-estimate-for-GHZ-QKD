`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBgT1Yp0Wcj1mShVDrNNRzZiCmZBdmgLhrgJBhfiwtkcJqI5uzwJNHTLrs/Fh8ng
ivdiK/WH9nw59fLhQSgpxO8+trDKlblLdXVUtYQx6GGAkVmTXD/lvFbqV84Gf/Ge
c0561wHnMry9eER7cuvXAcdD5n/AWTL4ICT6kyetxrRppM+gOP3EVoEUvGItlKAb
wjN0U4CYCRI3kqHDR/r/gBJh78ZEn/TLXm5UdUNyT+BfzWbHHVHu1H6cc2bZlwj4
RxHgDt504K/nLkdZ/w3QQ9wsQDAmIE78ig82f16aL1Vgy3trLG7+RiEzwvJEwDVs
8lsjFSUh66pEyIIYBuViFXXntuPDrqrqoJoWr9k2SOQTfTl4+jgTvG/OwzZ6uE7d
oyeiZ4aeh0Tnw6xNv5E5XSbcOgYdMO1F2IwlVhj45CnqXeNp8bO2LDW0bdqpaosk
CEyqtKr1FzDueSajqPkCGFggq/N402OVQ2QijpcXmYFHalaZ3Q5kHlhohrUdgIe2
hjPBbwFt3Cmr+Iv1ESjwjkbA0qVzzLO2IxbS0b+wZ3hO/l6u91hpkgTqvfGjDB3q
95OkdkfevZuDXK6DSXtMT0N0ZqZJS9AYtWC5npUDPcngRs0UxLoNW2tu0YzdjXh2
FzzevnDgh0Ls4QzfG5XUzddwD0P5ULJFali78XrikwvJ/hYvaWZ9eW7LE6TtsvYu
JjXUtLni9HaBLcbmfpJiH0PMXcnhQ5G3jDwDrAHp8PDZmsQIzpj8Ok2HjkrMBlVn
xvLqvnyL2w8u12RrimEMUA==
`protect END_PROTECTED
