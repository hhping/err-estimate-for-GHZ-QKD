`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JxkcQjmuY0daAy7rdkkC4uxe7ybXPloOkD+f1mqZ/qBLgWPQpqIY78PFD4UKG2Yw
cHs/8BhFm7Gsq+q572VCLg1WCX3OCIVJzUbJw12813DUp7oWeUUsESnM8m8NefoA
d5K9ye1e2MG1yeg5BV6RRej+akhf/JlisiVCrTbcRK+BEq2QoIu20fZsHu7egjQT
1T3O7xyKzWJ0ofSL2rCmSRAYG/St7drtpXxHjpClRSn4bu2QuLt+t4Lmib1tM3DB
A5csyL9cDLI9ndQJA+uBhuTTmlXFAWTThkGY6MjKbQh/CHmC2buVuL5720hof/PX
Ql1hEeg0uo275rritByyI4afbk71/om2t9auc6omS4UIe5liH45akLHFINTELgtL
Nu9KBvRrI91TWQaOZNjTc8kOmck1Q+X8XRVkb0fVkyc2iEpNcKNi6mVmhs2W3DTr
townrTrlijoPIyw4wVEM5K/85KzXAGvNFEplono1wqESfQuTSL4Bq6W1f9gsfLjT
tmpdB4MTZ8y8IPTGs+dzf9FyRmrj8MrVIGlgVjIKhIG3+2wYDnpnreaDJ4ZkPgit
QBfYuLILOXQX92w8+UdU2D4kervTMfjZGmT13vTD35vcgLsv8KuJ9obSMxZwk/Au
4Nhcht8VsC9JHE/INBq3LGCHgPAwFmZRd+JiEbPiEx7X0b3McahAsiHNKdj5hDX3
32ZTtGQISLhIvE21W0RELVtNf0B2hVR2HbtMeXU+l3crUc6IpCM0kNzYTXWGlWnJ
SGLZPKd4JRrkrNZC5AJxXgE8UGBs4sBjrh/rAqSNFQHH7HHecIVFIsXmk47Jb9Uf
VhOYzMrU6n9M175Zq8A+YOLFHnnMUqUFnGHqxjkqUZ/YqPebnfySfQi4xWA6uTz4
0f3V24AF9Qb8VTb8eMbDVTTBMYy5aODoUeHURDhRojq5nE+LaCUycyJ/TbuISAp0
W0oFc/byaEw2IFXxplLlQFFM+oNn8yJ60rF7Xcw6ZX6UUi9VbDrD+EVmX8BKuadE
Mi2R5Cm8ovCelcRQEfT6/T1Dt3pOnBq9IMUFIwWE/UX8WPT7CW6ZflX5y2JS39V8
tXIQ4Pe1RJDDdc777WeluUOKE6PYd+2zlTVkCoToLgyx91wxsA8h1IqWBVOiMMt+
MF4hnl9uMboX80Udr7E7RdjRIFtSE9IdiyIY3iYES+YrDfocqAkSryQx6srEMpiV
qo5aG6vGXdTZcKLRkWyMQLpaGYLa1xnKXnq+OZbbY5rOvJW47ZUsd0SUanggYYil
JQ69aNL0djqlwrDnprfroTS0/Zo0OzoqljyRrv+I8zSclF0Xu6CQ4gFcJy+hYLa8
UuN3KD9UNgT7ju+Lj57Vg0LAuDZLG2sUVt+P8c4dnFQsyOziSohDrtPTk/lkaNKh
XDdNrY/wh2tlDoxsQ9qisa+dUKq+rjXOd1WVhAykl98=
`protect END_PROTECTED
