`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uzdcFROPTall4ur46t3p7v7TWXQXeVYbJRl+aCN508WHZxXFhBIVl7+Zufzi6Zr
Ode1Lje7cGgcp09QgAiZotrwp+rBzB3NW0uA1JXe02bz1xZp0HyCJsN0A2Tl9E6n
xG9AIp3T9RQQxv/bbdja2vMHfHKVG5IPmtWcNLLieuvLttIH/CqEfXLMkNLCS5YQ
8SQeHNb+g5svw8AH+CIPgeL+zSJuvVm9v+zsSRpMggw=
`protect END_PROTECTED
