`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrI0nKkFSVlYKgkT3kh7sdsCSTfBTzEYsBiAou8s2hKX7KnDxPZlftosOJ0biDSC
17cvaGSfZGXjl+20oSZGKM1JKOU44W3ZYm8XzR8eNFWGZYC8q9jAvbDqTesgEET/
/dY0PX9PLY1xMQwERybSa7T4MP4xHU8/KhS3Uwp32yvehZm7qt50AemcDcDK6ybK
RgNbY+Wj2uTfLLKGw8I5DHnrhwmIxpatfHOGkY/5LpUo8w7qvILW1LLb5NuVu/Lc
t74ncmT0MxXJUoiSoaBRY2TsU94T0fHdqd0CrS9ZrqoT4mprAkA2YW1+SJwXhnat
tPYYnLPjuo6gRl1ais63bWjWDKeKJHPF1Mjrt3IneT+M1sTWVFM4RSlivLn5WHwT
MxclcA+GJjKqLD6er6H6Ll6IGaj87AEstG83oD3Nd0Uwof0P7U/yNFi1EOB1ErCL
/B8MSwirAEbw0PjFFrHX4GI7/DsP2BMSNIiE07yAeOxVEntBl/IioQYVqXDYHUNf
80fbSsoEJrV3+yh914euaRAaTR5Hd8ZaBhtluyNMupFKp32Gmj3WUjtjTKr6ApGj
ejRKNyFcpLbCOE79fxnE8kcJm4gyG+SVMc7SQlirxve63Fqfbj+XPmjliquqeUkD
t9hnvfp211VpVp8jQbH0NA==
`protect END_PROTECTED
