`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B5XylP3x7FfnlajIDu6D9iBlnO/709ln6Wc++x8IkG7dp8rjlN5zRAJwaDT9cjz7
2psRu7WQ1x+B747gSyKNYI0Rb/s292+adPJUI7hM1HOqpmwz2ggn0ZhXTmMaMSvq
EVTs7hhnZkFZOMPEINr3MT4oh0zTNCJv4rywcvo11kVfU0b/pcZQwrS+PFhV6S6v
HLuMUHzbNhk9SHpWwEt0hZXWTN3VY8AnqdT+y5vSrYC6ytPeuVKbluYmkIGqdpM1
msfyzGEsplHWJxWvSztst75wMG3npnkpW+Bkw1MJqD0xLdBT7UOckV/THAQhX1Tu
b/dAGwKIUL46Httwn7md3nXOJfw/YlRwONETEnUT+z+VHnJTRZAqDwaAW27b5pt6
ZTAGwb4N+8uOJP/8Upk1Bp1yVgqsRjUzm/MdGAqSX1flDKDnR7VhFKFqu+6EVe3G
AEcDHxfP8xkN9R64Ev+AUw3beXi4XVU5uJwSct47LD6JZmbyU0Vgx1ulzBPQM8rC
HcnYtug4ymljDQvDolMKaDyBG/3b3VthOyfeVBLzmZJEdzyDQNvS1hJZ+GRh7Dku
FkovWqNqQSq4VroaEcUpi5RlbeXeOv2dv1hgcXKfb9O4vrGjUzkX9eT7b4zNVyo7
3naP87LkMCX2QR1RRH5AcXO46ooD2SlqeVPcwsYkJk29xpdhYbn+nHs7+KJSJrXa
YXUsTCZCWpTd9xahvvUTSEYs0CisMLK2RDX2MWjSV3yq/ZxcGeShpAzz0wGgE6WC
7Lr7IuVeCRJQrXO9mgIysWmAuqRoWrobsLDO+myo9ePI+woGXd88jHshG5A4LQFb
gGvtmqMFZbRHoTiMK5X49+tj0arj5FQE+6yjLB2AGhQRR6L0vf7k43QRwjtuYDOp
i0NJUauSVG/bYys9uKaENXoOV78ruEMmsz/FT1AQBGBoaBbcB/+kBZBepLAHM4F0
FCqOpl//H6hA5V2TOX4ksm+uJItE+39tT9cvwuHINfwIhgCI1QqGTcAZrRGgCBFq
D7LdIKHyn85F+pmZ+3Qa8WkN145iJl4Gz11lbcclmOU=
`protect END_PROTECTED
