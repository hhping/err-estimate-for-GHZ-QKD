`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+82qg4E23KrSDgHMkeHh7/25UTUnzVHD1Ko7ivRrMnyMd0M8FG5nS3kYlCjKTT/
3wX1G1ZVd9QC7XCGBv3Gwr3J54nOwNKuJEP2FG1FM9Rr1aq9ZQeoadXzsacjEg2m
heUwmZr+MEfp+gFF3cBMGMeUaPLOoxP7MP2vv2itkucUsk8gfZXUGxU/d/ueIgjV
plyZi5CLc9z1a/JFC3DTe74SQoDnw1SSU6lge4Yvs/tsI2Vhts4ge2rS8IB/EMNM
A36QiuD9KeStPfiNdxzan57R94yXjPF87Qzl7my5udg26vXd8yi+XUAGY1/B94yH
zPjJaFmZR/K5DmgvLwbpExfBIr2Ff8uG9LbBnl62If67q0GqCCeYiqqq2niKcORR
Gqk8tQwY1qN/x1gJdjLCYHcjR9tL4JJBjwfKjphhxKEoVGlw2xA4R0jtnXidlPfu
5NbfAIKO52lOnnBkp9bHm2mB0cjE8e1Xhx0WQwD4klq2ef/N/XHVHuDAXxFE40J1
6PykHzIc02UOrGLzYYep/wcH5osBxkuQIJsoiob2b6d4YNj/h0I21hJ5LBO702Tl
BLXT73AceuDOC10MaksbDOHsiQxUB115Vy1bd9Mdc6u6Q6CNDLZDUP+LZgQJUVbH
jfytxX3+29H1W6R/WEkhCNr7cGz1tl0HJMTkP3WH/RPXwqkSIgKEqZ/1wsrumeq2
bMEzZd/f3uzKkI5qR+plkAg9fQgYMmSdGDob5oeCz1tdyCggWW+2OB5RSiO7F1PI
skajZNklIxR9dV9Gp7Zf0UpwsH/qJja+q80/90RPjn82KkKIGlcs0l5HcwlKiRSm
1jHtLOqHT3Q36qQJAtRVNucvVkl82IPpzklS1PhfUG20ns+W6Si18A/+AaI8fYGU
q000Aqk7D10qXbbzXSXKKAQradj89UwG/1NhbGXpNn0AuGM2c4Fn/q47YU+xibzN
v+UVbOSyIBshyBUfodabJ+zz1w0O+LpdyfzYUKUQElpSx6DNGkT0WzU8+eEAqYCQ
ct+1INfalf9EihLidCDVxhHgWQwmRIjdyJt8AaIDwnLuEBfmofY+A1xR1nLCI99K
bu+Hr4tdDRJwY7QGcWN61jiEx9cQR1tt2WKNaaQDHOmiqeukmeAFiJ+O8CT4na07
CjbMQ/iSWg2iCDGE5KX6TZkVvu2QAV8fBhsz59VelGJGjK3BI8pcQ34hEmBKKARz
1uQ2sbkbOhIeqtQ3YEVsm9VeSxt7AiNL8hnAeYEWHLsJhKekSHvuq0+sbClKJxia
1M8qYHfT5rhZ1K2PsyhseFfIJ2eVPDm03Uh8Zz45nbBynLOTo1w5pimX4QG7s0bN
HzNjbb8JljdRfmG499+0tXoNBpWYXKBiZlpiEIqOk4hjVAA6yxrsTVXDJB/OdeGV
mNNNjt6EpxfxCINPAAg/mxK3znCv5gWnOxybhcC0DgyL/C35bY8OjYr/Yhnv2XRm
VCVMF3Ixh9Fk9waXQ4W40w/MFEsj5MoAPgdJUKswAgx35uXn5BYibYpyjTQcGWyT
zYjmrW78dNQI/70Gej5kR6e626gQ5L1vC1Y4lp1SJMcWUoljJ6ap0Qhp4j/jhc6E
33ulfmXhZfEO5smO0Pl4xIsX9ZEZhYgJTDCeD3x1R9AYOQctmhDLIqL8GNyNH2uf
OOpQsRWpJEKFK1a8Q+RdjZhdM6/sp+2dGfYgIx/SyAl8eOzs1uvmPxPDfvl4fagx
loxBPWzXtf6/YcRBY+1y3HlSRbbDO0cFGAqHWAOsiwh5lXM6g97XlMNeZuMLAVyk
GztYbjXjsqYtau9F3X7fFyVOozqPqkfXzqM6hzExu75DNE/plSnl1w+dK/z9FNCl
XFXaScynuehh1yDA9h9cZhcmmlSCz1JBkhJhoAuSpPHoraY8btNYqKI/R+L7j7cV
UXI4BQvzSrtKfNILBheQaKNx1UncwnS18HYN4AZFKw+gny+fN+v+jQFEuArWgRvs
xYayFeKnPjlAqZHxrChcI2c/BldRlG81C75MJXGCngMjCo0yPysT6SwY0RtDyVYr
NF3Sk64t6WVUe5czsu2bfq9f1K1n2m+KvN+Wv9s4NXjlv2143Fl/Hc4rKMX4FQfT
j4iXBlW4LL9TXwT6i73PJ0//WFaTRh6/pi7l1l3gINicTtGUsFTWmP1L3UmNPCwV
W7OYLY812WkDYWmberEvGRoXGcWSW8XuQNi8yPoT2oNOZggDcew3It+6sDFwHadA
RJymWtJlsBrur5lxVwz6A6A6gqzXFagAAIIjVyn6PEO1gMIqs6GGvL/xJcf0/2Lh
rwh9BNkKARHjQr9Y0eiB4ZgKdfDc/Rw4Tv8AS5TtrHHBaTpM2qayWKt6DVAMy1lF
QYGyH6HBCXg7+sNjT4WspEw8KjNMdkr2LZlUH9UK6L+E8SDXSiE7xAhcQ4sM76Y8
y3NnWnReh4XBtulXqxt1Y/gl5XBsCNt3BGN/BrH7pfZLC/9RuQIsgw378+MUiDRV
A9mWUlbNUiSYUN9RUuj9Ae7stI+02peycJW9bVCUI9U/gKJoTHeLCk/v6GtkyfUu
bpgTBLT9UHA6ZvMh888R0D/DwATAaed/D+t++QYsqMrzi3yMf1xqnZVKKXtHMLTm
QJk81xdDNmz1S1s0TF1Ve6j6E2TCOOfFXsRhswN8AeHN+mcO2vZFkiacYb23SP34
sGcLLS4Bddc0tWBLG8OkA9h2g3GSUYNd8r54R4aVkTaFbh6yKhag92tgglA+iLLf
J6geKS2b07RTVCaFrmVi2LUDwZqa8e7OxVKrKgwFgfigggA1u4MG0ncf1oxlnFkh
kRElCw9thbcGZ6Vs2OONrfZa0Aa86bWSAi5BzXowhrJseepX6rBusrqsFiedA8jW
nP+owWiSG062Uraant2p6fJ3Elkqybr8cjjn4uCrQlLMMgw406y7YnIZOyKYJ7l3
3to7dU088w0A/J6Hg0JVUD6HbsnHDVhzqSmXFu/Ef2vHZ4Epasp0YOhhUr65HvDQ
BJabTUMbdrHM9QGmyYheaL11QyyT81d1PE7sy2ZBs0KuqHVbgwVNpKQcKOMo3192
eisuSqzfthBAi4T5lEVHkiVMe2JARiyW5qTQVHY7gY2cz2v7Ql0RS0f3zHBmgaTH
KXF6rx7rd1Zu90OhQcIQqr7NkbsZKlwFnwvE2LgmpSoWXtfQtYlgzfsEuFeIOXLp
4kS/cDd2H0nN0jPPSslSN4CCDYW4Q5IPu43oUPcjax1Un1twGgdU5n7SdZX+GzGx
fU3QodNNgd9zTWkuNSxeXQdp1qlkSLSHrjDIKxMTt+87Sro6DKpnyQZ/0Kr69LCv
DZMMm66eXZ9s4xK+gjoYJk9cDaWuz6peLOKxkbGrz+wbxdm8lgxNeWtZEDDfl+wp
M3MujuVSG09oiT3NIZdwYwZhRkkOgX5tpvNNF0hlrLli6NHUCAIOmAazcnOa46wI
RjP7aZmctj310S6DHxTQZgDmGZZ/fuPdChy+TkI2LnQ2xLsLcrCKFekJnmLfzmdv
JxasrfqPDXo+YW0QYA2oA0KA2XYUb8jJVlbt8cA5oP9/RdbLA8FsEmufTDIiScMi
B8ccSkPLK/Ehv7UurBO5ZrH6CwtfTxtyPOzKzkyD6OsXSH19JzuFcOipbOVXV3ir
JbgAqQqzJAp97qLZAdmX0TRptvS0waV0Cs+GmNPzLUH9ILXCBZ7PwzNfr6tIIezz
j6N5z0Lk1F5d2OnZg265/6TvH5saypRN1E7KT0hu+nQo+7609LxP7Foip2g1WIDd
nYR6Plc8HeD73Hb/iSZJ/Hgo6q+e51a3OgN4Dkyp+1Knc4v9/jo9bf4o6r02IHJy
52NVp7r2cej9oLJuqOf4rBQ4BbQ2q/0iCg/cv0yWtN87Gw7iNMUs7RubWpDE8IXH
T1wK/9xurOPTTpmcszSk8C78uBFr9jXso/TJq6rhLseYZ4+ZxvDJNFNKa2FzyUdW
7Ms7DEzgOVcALeHVnV6pwKtwQNq/jrE2ge4TYrok5EpgLQ3d31cY08kN018RU5u2
rv6yhLljlh/Y57ztfzg5HBwwxDvMKkx1pKY900Kw7PeDYb8URCt7xkvLutEEfWqI
C+R3eth/Mua1imBf4Pg9uYtq7+sYUxL/20R8jh092PEKxLoPutMYanSXLtoDLKgx
x9uM90XRSoxEi0Tvx7vneex2Hq2sCPQVvAX6ZrQpQn10esLKq/u8Ep8Utg9r6pIz
g5nle2hNyuhs0L+iXOizF1vtyuvXBnIGyWLvf0ZhKoUxqw+D1t9JOjNc2+YeM8qF
a++jBdTQyEDFv0yEJcfI96WLEzxQMlo0zh8Vd6xkfnesppBPJEo5OKXTqPKOtJqQ
DbT8hGMV4qlM3sB+uHyfdpBEvMJO/c8gQElp3AgyTPO0LmMI7OnyCmjdjRes1RsP
5EB3cNaySorbCfKktrRlGiU1pabL7FPUbb9hE+t6iV3+/IP8NFWFuusngNqq9XEE
ZO0PQNHxGLjcncYcmL1HR4vkobrm9B4mMU/eHFkVSARRiQ0yFpHEkbMB4DE5Al3z
zcVOA2AJY0n1Quq0Fv/l/JjwurlL8eEBihlnU96Sa91nDkpq57pnFwXPv8DEfQC0
pyV/lusuVjJtipZ/UN2EMBvE1/yXz11m/b0HZK5PbwkmAKtqPtusJnTSckSQhItE
mDXPqT804LRqmM+MjALRctP8otdcolRN3VrmWKrubHqVS/16YszfLH3g9ysuLIKa
poTulNNV6hUNJ0a/o4o3TM6o46q+8nFJWiUPf3Mx1cWaT/tT95iMbY/7cJu2DrKh
2yI5bnfyGyaMi/ReL6Yj42E1qXosi3LTQhiUr4YHqBKYjh3OUSCn5VfXT8FKGahN
f9xk1aWYfgmJNJn8OdxIWbCUrkgdenjXbfNLdOEhSenMiaNEdzbNRgZx2J9Yz2Zz
4jqLSEz7M+deFARHH/nIrePsRKiAKojXa/TeiHwWamtZYN/cQ6gNlLhJdFsqq9On
H5zYPW+Ti8Kw6KNG9iK48T5ks4JG7IEPK24tMLgvIfJAgtChEyBsYEEO2HCcfn0h
taTxJLSv3bisgpg2UhsTHN9Y7HC+0UFgvglnQ93Ael38kwVwJGwxQr0U8aNDcbWa
CJxaKdK3eA+qWVOVWPvykU5rgVyrawooesGcbQKzW7ccGkSp3SZ8Vcd/53shfViL
pFKZu/4cWWx1EjEuEMTHuGY2uA56uK0hZsLL6UWN3UuobVLaV+Yzpa4rrnY7RbuF
b8immOHGQjG+KrclyDXhX0Jd+CT87pfyemk3chspslfrfiny2tgPK7XT5zZJ1MJX
LJ7LwEfyDetChVcrKrqDHR48qWBC9HzekMIJjK5ZuEMR2nsKqkrPUbvu3rJxt+Qr
93jhxlksuAtYrzhwcfj1trbuGVB4oyJLjay3sFnCo2UA9qRBjmV0fDVFl7M0svpD
xGDaaGH6j8N6iyQrxeOz7zH8XnihBJWcJ+yv3pWBU+MVaeNTdLGDBkvK7oHVjvXh
5OxELornTYHEt0qK0oonwu+SmDAbOpl6PMtRVWSENCYmM1jsH9ALAcutz2NV8qb9
R1YysMqat6iuC2gYXdBPCtuCx54mQNS/VgZ/aYkALDS/J4Tdwob+tG434XOX2bNw
B6uEzFchDCO1BiKSJ8HNWi07IJxEjEdcUfUvzb/8BFwewzfka76GC9Ad/TtWewTN
RrCplwmdnQw7fUPjNLnMYQNMhlG85uQQtl83/Ls01FK0W7K/rYC/Fw5AW4VMXAyj
Qs2NnnfXuNDycEh+MMq9WrNB4OF5s2SI2DB9oqH51iN5ZroXJCEOytn1t9PCB0wu
7rttFsx71rLk2dRW+oTsI/AtqK+WeGm8lNpoN9eIEn/LzLS1ZH/2f3r9+uLCBzUc
ty1ntuSqAz0s0pCxqNZTPFBkZwmipJi55kHiT4Tp1YnWRy0iQP2/SDN4QM8FQe/i
qAt4vE3mRS1cmJZ6oCx9XuUiKBTCjo6NHnuxa9xF/ygZCvNcrbyTX6IIu7ceXx2/
mAsG2g+dl133HanQ8v2Nu/0soWvyfqhL9STouBVu0tg+HzM3CcmgT1j03cDnWm9I
Oaw5Lt9yamdKv/exXXtiyYQTu1yzrFW7UKdyoy0cfQfrOmmTYKjHMmsQq8vo3YCs
eGcmblDHCiCtucUdf/El8q9zg/+EJI04/r7F1brJfv5jSIK/WvU5QsnFA226VNYI
dkY4zfo24WINBq3zU0yitU5GERnPxBqUSDlT4IGsFc70hFBC68IJtBgg+9kt/YZf
V6XhXSGJHnLCcEe5fozBRg6vGzceKAUeRF5F9BCf0wP6QbZMvHgfbeeW+R3kA2xi
UXfynzpQ8sIvX+sY/xwQUNX8I22jJGGKlsRXLqjEoAosJbNfZk6LufR2C1gbyxCo
zUV76pv/ABa0nQ3Yc0hHugsUkThbxpUR/3o25i/vn2o29Dn1om42ERSnMFZgwauG
1WPATpqcMHVE9G6Tl/fxdTn+o+wGA9rp3CFtuhjCRqaA34PXrCP/3IWtuUMYJXBy
+ZXQzgWqsBhfigbim2TbCMiqHkXj7ha16O9z5goWai/hIkEn4uFJzH6nIzM4PWHQ
fSXiAfj4tcqhJ8gamardEt/eCWMphF52RqU7YMYMwW4pdlCswEUBiPSLCT+EIu1P
xZWP4//DIZ87cUrUg5WQFPdpr22upeTdydCAED60mcR7Dd/G0tPWQ/eEeOnV+AuP
k0ik12Vbfwdya51epxPnBoUzQ8fVfmX+TQh6zEAzJKGDsOI4X/1dRl8QVJNSYFTo
HW+NIg6yxwhK/lV+4zA4R3utKbvMcnB6z9IszPY1w7LsDMVkm+QG21VmMxb0tExh
urd41LGBLTuJRWYoaOt7aJL4Ire+OgR0yBSMvNpUCMwEpOwYFCP6C9QjnS/wgq+g
1Un+olF4n8GvI7EYlC5sO8GtuwGmM+W/ZiK4OvEKrL2DL9rZFTDy/LOy5nnKNeoy
1XbQnliN/+ErCcq1sa2iNCktkiOCawDMhyQXhjoMuQSqict4j1jQ+23FiYl+G3KN
y1gJonjmUbu/ti4z+xjHGU5OtvF2+JcCHzbME01peNuw+wjyUKxx2pzAMPGutYuJ
BjuVHgoYW5hAdbfszQVx82NDY8VyOab2i2xDgkO3bd+AE3w6Njhhij6BN3fLlOCQ
K89o5cfAAnXavURByna0Rfcu/HNWMLmL01+Z5CmKhgkvXBnzRU/q5W2AOqDldrhw
8O2DLsamdAdQs3i3Ghmre0CLQYdGEf9C2KrVSc140QkWcOGYtDTjqga0KABZU4Yl
SzX/vu3cxfaNJwSY2MkCrswjuK6f7goLUl/fz7ibEgpQzRDPC8kTW90T2Wu+mTfL
J50ZU6Hy8ABkdGtMb62x5ABJG64qkr2yo3Qj4qvqPalML9evtY9T2aWLzOZSg1r1
flcRN22YyRqWYaZr4nwyT1f1xh2i884+b+WOqDE1i0UVHxrjWSUxCSNTBF5YAiSb
L+ZJ1r4K2mHD5NMc9Yxmw1ZHHuARTV+dRW6ja6uPQBbn+oWrXD03s9oNhjvBkn7O
TKgw05RxaLiKnwlpoacxzRsU8MvpCQ2ujHvkxjBc/yPsIQJpMn7/4LDrAnAR66pZ
TGcdQ17tQIl+dgi2vGs5QZb25o/6+7UvyDNRoto233BeqwXB5ToJnG6dnxPUSpI6
nT19myhs3l+cwBu/MR0s6QfMt3Qc8hwey2KOHDnboXIcgIqNHejEpwmXj9B/aykh
jd822H6sI7ajHrlw5SrGZhwNCTAe1PCItYKcXHHt7sxz6SxTcgv6XF5zc9tly9N9
I7HwbMNIHOL7++6FAfvedhrvW9Fn1QgbytfjRe/4oAHshMHzLgk0OuiYT/VeT8ER
jELJTnw4YWo/5A5lmbnWEMM7snoIcSdEmtIuIWj59bYFKMBJqzOnCnl2YED+B1me
wTgxqubUOJnqrufJqZoGauprxstazlYxJgHpoKKa8Fh5lwHM58Yk09x/jUzUKgpH
KmPJjyarPhdhMcvjSTciXj6HUyq6DueXYo4tPzceiX2/+swy+y/vxX7yNUf0sO99
H+OvlqVSt39d+HeHoOHVd6UL6r8NiXAmW8sFg8PQVbt9O9ekzMZEc3y1I8k7NrHd
fUaUHv9CdSiDC0qzl4A6d3M5wFGbT9UI6tWslgy3iPzNBvm7sgbRqjK9LEVl0oNh
PKJQuXUmaDMY9HNQkl+9uqnIOC9kyQcdwnmkQR6dfhs++WylJ89oAidYr3GCa/Yi
YrhSEKwEGSrzkm1kkwBxrUlPADo3E9NA0jWMsa41SWHuOVJzPcktyZWnARpRq7e4
B71pO3nvfLj3hDjc0i8NJs4VhaurG+0mTuQVOWaK7ZZa5zX593NKQi8KXcjQxnKX
L5GuxUNeHju10AoLPh/p4pSsDFCzBOPjdNcaomr3TTNSUVPWasKl6eUZP3lWMUqc
D++RKydzTA0HRo3PcafW/hQOXpZd4aia9AF4m4so2VVKoMtV8bxBETZyZPV5knzL
yKtMI1G8YMhG2Gm+S4XLffxnduM5IPrREul2+1G3a97K728a9a8DgaL8EbBiwyA7
N7DDiCzflObkK8H1+UbH6dgDaZaL/B6xa0bAukcdBFiccatqi27pBgNJ/C3SJERQ
tO0cIpxyXw5i5slk6O2h6ZHMl9yUyxOLhy4xHWzWMTCC7JAukjVvbnr8DKG2PPRI
3L3p3s8d8irmGpQmrz6eqZ01XKMgl0nxvD7+5KmOMoErmz5/gG54j47CoQdoo8Il
gw84D6eeSZ4llAMzRAEu2iugBCfMUJsSoMullMWJ469nbByLqPspiTP3KTVLPv5+
d3t5e7i+x2qe9qG1k3tUESUJoIEvLr4yWRKl+6xK2c0+onarionVq2mfirI6NK8/
NKKjiJd34CXSlvyrh3BUp+5z0LTLBkWU9LtHBUa2rw+9ccm8B8OJPjQf7+UHx9nJ
PMEbFq9TSsRz5MeOX1JAR5dyzDud0t7y1Wdo7rM0mEnpWDQVSmDol42YtZ9gwCJG
kYpjpjlDHGqp8h7fYMkmlGjoGSWg/yyc1o42Awl0SPwH66WCgyMMO8eZgoqlHDfS
4nu1NQ1Z8xB+dGDjxGpWfR7rbhU76M0TEjCR1v3EdwWlf+x+Pdp+hsrTGNjiSAt8
Jg7oLWrJvttSzepf6+VBm4uGQPkTyWWgOJ9qkdmr7OGiID4sMlhJXvMQ6E0yjXqP
FrBnJwH3rFeJ7chxHJbnD7f1oMA1gccyqw1aWjEbjIPTwFAOEWCbQKCqs4e+STcT
v7X7e7n1LzcR86nmAXHpEl3q3kQ2MskeZXSzcVP708CD9FMQADV3U2QGc/JC2Mzm
7CHrp2i6tzvMbuOsci1h1xfawRBAKgH309V/BdSZmlKT0yOuIKtaycBbfPA9jbSN
qLHIAQymunGhvi19SxIIyRXJvcz0DAEiRSt+zcenKzOeqxD76fl73NIWrtDC9F21
SzDoff0RsB6T6qTuAAlCW3i8xKDb+4HCjnjhbPqy7rzaSWmGYmpUlIyGkIlnM1Rw
jjfwpYe5J6fEAGSl0wD1BClKyiG3Oo5ZUAQ0q2UXydZenGMnlYp3kvbAUVATyduc
Z8zXbebPg164wVUpPlBlF9awHWFw5s4mSu9jPckzs/c4rWQE5GZDvARJzlc86Dq2
6ctmDHeqcxU22VSD4R4f0XmZcsrHqjz4m6zQO9ndkxfI6nltwmRVMDUIXHHE60TC
wE9bledxJy9dE4oZnDyOKOLeYQ//xNhRwAzOkXvc/nHvO2ymDChTPtCyfuo+70b2
7XaWbR9StCXjrh8NeB8CIV79BQa2LrckKRBEEJX97536uwpGZbNnDB5poxXtakyx
5xk5bD1h9pvtktKwiE3JNrAKGKRK7rZ9KBSGPEQB+tADgbeLH20ltvonrVmwhB+5
O6f6czJTTAHJ721CKqfo3+clyL/aN3lbnrYXn7hefs7GSFWEIpPeumWIkSCqTZVx
F6H7LSoiYhPXOkIrWskG/AiGfWP3MHq/IUg1Sfk7XI/1z/p8CbN/Oxs1T0gtuojN
JSpv8XU7u/Ruc99WT7F6PmYbUun6HZRDRM20n3HWdmR8hNXT7iH90bf9oI5Gv5JQ
V57CO6+lNzGYVRJnseaddgu5nqrLP25Sz9TzELyWhEPlPLGcWXKTnmubi7A58nnr
NXTZ260ojIb4oBg7x/qrqmgW7Ks58dJrI24wik654ASiSPFkiQcdwxfjxAwguiph
Rf3MHYM4zepSzBqcEGsvw2mx02HG29ZJMfDVt/qHC/fbWfiI4GzBCVa204kVRbyT
4bFe9Tc2CsQLb7jzZHDcwUes4o3V5NqrdWa1i9nh7J1lkFtsTZwYgHFJfpHH6JPM
MYeGl6pqnIrWfLrWYU1h6bw6ZBn21w4nxCBPHg8ywE2XjTanLJ7aPmhUc65dMgL9
n61u8m/+lB9NLjdxjAvslxKW3mMb03OJJFjh2xmE8jRIh01jtL+Fymb/9FpvbexY
fy3wDpt/+lwTbSvJCJwhCs/T0RPG7EgeexFNNEwYyqo0korDSP0Hx9jeDPBj9vdh
z7IC4Ra12oC05a9lK939ux/NV70AWEj8kDsfG/lTeYWVwlp3ZgG4Loy/fOTaD/VQ
KeibujDHQPd2vIpVmcOoB2dZkT8mMqjxRTGYgVKSp36QY7nVcVqsxvagDP8ZDqMS
n+qRSsOUqZc+aCduSHsMvIQ3fPqLMyO9+swRxoo2Bxyznv4NxBkDrMvFnBWtP2DM
mg26lerv5QM2yzPmvLygOCQbLM1UchcqNbGASDcUQC7AvQEEX4mizYMGhnfibGZL
BFE7bqQXxKBVuz61Fo+GsvWZz4dleI6T2hkw4S2DA1O+5t35gc4J5S9kUXZkYh7o
/mP/J1cxT1QMXaMsrm990TamyBYjckb1o3R1aY87iV/nsq2L6nf9Qn4lp5TXcp3p
oAlFTrZmvWyW+CNi3CtIlYP9PjBEFXsJG9DLzXFY+ndPemqT3FgqrX2uUni4YmmH
K/BhvNJ8dELEQgsTsTUaeHY0o9/+HvbDcjVsqTYQsX1f/1xgQ782yAfcmMSVhPzH
kKeUAxJT5wQ/nfWjauV7Agptb2Z1OUIMax/jHF8t7ygXr+KaBIy+6vTwKfI5Tyfd
tRSSscDtVDj+RINnQnyNV1ON2B5Uxj/zlltFQ6qva4DvGT9psueSB/uHxk7eLK7u
QLYCwiEPAEVxGtjJ5g7Hz31LOnUYgM8LxDsvUrfVq0foTO3nSgQ40CTwasBGeM9i
w1MZKvhvteTx95Fu0NZjnb52JPWmyrvoYKfNTjQMEuTqZkCDnEHOH5QmCBTtOSo9
xJFhJTUCZZEHV8319h0j2GHFWajokEiRypF2qk/43Tb/efNHCluTi2pFyRA/U5Rn
KUBxZ9GBuDgh0tgcyjVJOUehgg7C0EA0KXThRnLIM6WJK75M+DIdt7A2YcGu61ic
Uzr6OSwlAoGf2sRbhEw1dPLKyy5GQqt1CArOnddFjaY68/OVyPvr7zYSJGAD9X84
4kgf+TRP74hoNXs77j/eaNT9VmHSICaLJEVcRh5PUhXG2VCQHn+wfeJztD/ksO/G
sPy0APhj9x3tEs1+rrBiR2s2wYOkiw+hZxggnhg6k7Ftk46mZ0xeanEFEVkITaiY
A5cWtc1aW6DOzts9/K3x+pwuNtlHNIh2XSHbyZD7ObWeXVUmgJqkwTFe1JJ10gyy
cHQAJoajrI8oxPttNbtbf8FWUfWRQ0Oomme4ithK9JoRAcfFWkwwdQZHFk8r1a2X
JM2cGl1U/bIRTrnhVokMuRFHn+ujlhHE33nkaCPFlhq/FsN8omLFsWktcnr94cBa
ufs5P/ht7P4J98J+thTfO/S2Gz199M6/QIxUO4evDiXjMpC1AnX2l1OUA8sfb2Zb
E1nQbN8Aa5E279hQTN76AhboyJMdNzFb1hJ+FMsKgLYSxZjHcU9sCdwideO6ZrGn
1ECq9MCBItLBBJHmXGtQYv2obaE7Q8iOXtODU1glXPKuCOJc/bOfaVw6Yi3SLyg3
o01b3q1NQZXgi3fomHR5eNXFY31EDu0enV5bOw8qbT/VUVsEIzK5NzcpCblHkUzP
xsD166ciTZSgqdPJqLH8QkYPqfeGb6a1lipohlDesc3jZzOYRL2P98n1KE9BA3cr
Cd/AwFsRK1TTqQGxWOQZl1Nfvk+6SpbIzmhUU7NAHh2XQ9Vzo+UD8CyuRz6kyJDR
JAz9p49G6nTEVAeFr4ynZXwDlxA2UvYmI+1R1yuaIwMnmbwQA7lBdBgTpNpmiphW
biLEBA69dA9SaHMutxIRYF1z1rLaMKv0d9sPc6r7VNQZ3RTjwjQMZdp/8uXzU0Ik
d/LEc9IVnItGnlAwvNF3NVcltjuj8JV2XTOHD8LeqvKBVQ0mK4lmNEue6oEyFceO
VkVoqmmFiXTPzN1LTU43bLGIWxNSnsPj5/obEEsik7ExHoNPRpd0dTnhMjikbm8n
o19o81zJWD3mGMIW10vLMoYqNJHoZiBct4s53KfCdo2CcL1waKgmQxFNSFANN+WA
uLFKQSoTi3TCwGfq6u1u3gmnzXMwiaSXjohEN03uNavgvFnyz0KwpDZXDBZyHkLx
KSaX6qmhkZL3nH7ip/kdtZZc9XjI5uGfZZjMVYR95MkKh+UGcQcVpryfRse2o24F
jlRu1stnP5N+Miszpo6WO+bxLYf4+llWXRHLm+SgoMjasXvuyUxyQl9IDtGKC5d2
hckHsRkoMdRu+M2yTqP70duIfKb+LmmHtOQdNHrLUNoAFrBHDDS5/xX7uENloqFM
aYQIsg3NTyzJeuTem/83223WdybLW8sAO0XyPH69xzhx8L3cX8OPWXIraAHF5y7R
K4avXlkNH+Um5qdzZA63Wq46E/KszM/E15Uq9UWKQ5rn+QkBDZ4wufh82QBV3urq
QLpkWAhH4bhNaODeCM2nho0x/72RDTySFGqcXLxorm4uqvyI3cCPemr4IJJIGBh1
W2g0kKLMOL+meazaymcMQNrd9OCRdLJd+DuVvB4/7+ELFQwGzp2wjXOYdk+U0znC
YvC6uC0bsyI1vXGloAxUjDm34UwZzSI3QFur21U9N5m+l2aqY7fRU6DEh3y2wzB1
E5SRSISmVZu/48nvTNt76kRejZOlg7seo6dCxND3/TLQJsexfyeJefT1lyvsfp3s
AJ6LKfzoCesHw+6SA/NTgPm/8omxzwElfBkNZOqfb8n9p5lJhAfgASmIBhBKVwNw
n6zkm82pQRfgqBy6Vup9UVP2V7HA20cpKwqSTRM45/VhxHj2Uu4jKUKBOheAeFO+
qc3ejrxNvjxJTMosgNkFfBxFrEe28G4gclhRsUKRaH3Ux3nfvJntFOwJnAXSSbMY
XVkLkAoWoDTemGWxwLCXhaUL5uBgXdRT1cYpGiy6jbJGlN7is4tmCHv9JNonahe+
6kPh6Avx9VHZ8pSYjzHkgbgGN1KmZ/5zGXWL2OiQx7ZMkEr27CrQ+tc/rzkJCSfb
+ZUgM1d13h/T8JEysi4IqQ8AURZMshZdPzceTb/xUISYq8WRQcfqiUt1Mc6GySZG
7gGPGrKZv25pnImUFszv/IlfjdBTOPvZ+4LRmWWW2qKlE0gu7GKZYYTGxbQdRN/0
eoORkJ7xjkIIkAIa+AqYoic8B9o0E9F28J/znUzmgYKHl6ycp9FaFS6zl+TfUneK
vVQjtT5RLNEwa3h0EtQsyINWq1V3mkGrhUD404xT1aql8QfBlrp2hlEf9No0ln8p
wTALsIY+e4Ke+VMgrOj3dxRAdeFXX0qMGyg5g8zk8jlgyYF+sZNVqI13sHrUcc6D
7jXNrQDUluTjs2+4Un3pL/RIbSae+KsgLmigL9R91Tl0Qo9DBqorh9R4hZLFuzyX
7bCJzbiCaq2neQZd83HASLsURTMLdH5i3kFDZnl3iD2zTaQQc6ZtPDxApo6fob7J
ty/yrveTL30KynolQxr3hizdFb86xH9sc3JacROe0nLXdBjloygt5bYliWqz4f5M
1Pb9ADrb352rbSlrMZ+ze6Q9dmGKi0SKOX9Yh2NRQ2Ta1XHcZUyZMov6fw6TjhqT
Lq4039074pa6vjVyBhhXi4xQLM4lhNp57o34onSI/2qk1R+ciRm6mlnGbSDufzT+
+ZRM8EkZwNYAxVrdWpSMFaj1VJTlQXNfxB+BKW7IF2W2hm/tcvRw///EkTJAn9kr
xlxpRcr6BP1fVuZbVbjukyF6ZNYXgRylkdKuNru1fR516EtAG8FlIOsN/zUM5LFA
egNkVQDrZH6em44jQ0rv6JcLZNI4YqSyKeac09tob7bquYUzWfOQjMufIon98vzo
6zoDEkQYoswaMAVdmauaCoEY+vJA7SfylNJAg2C6VKN3W7YB/26HcLI0qt3NQNdL
kdDlodmWcSMVYfvt20wP9QHLdj99iLpWJPtQiYw3ZL0R0maWRF4DUnAOWRGscpRi
tTuGYm+cqFdlYnMcmDR16YFs2sO7JuClCR3AqNowPe7Y1vEkSmAOn2FZtGnaxdcq
X5xZQXknd/cP17uCS41p5Hv3gHcQq4L0tVKeOTg6v68wH7/l0GKA/GhI0Fr0Q6Pd
ENC6oJMNirtkRqdS2CJDm+3L2DwmPam4IG0DofEZbGEopY8AGKtunqTSmlfqUS96
Uey2fBhuJH3yK58KL1F5iaWdHn5z+CNdvwhMniE6ngUpPHmf8Lu1AzyfvW4x9OE+
SsK9zpifZlxQGLw/Cpsk5RrEuxSpNkI80W1OGrp7eQmfkCEKPYzwYKnaJ5ut2vUv
u9MN2HKg1IJsZs/fo2bfXH8Col36/4m85L9jjvhAVYsV9ldl4Qfa5W3ysDj0hFti
tLuMS+4E2iMhSZa13Q4qVfNbKyk7WUFeSaAiD0P93fHzO6f93tvVXeJZmB529dfY
ewQFKszY3dagAmafQU96x2cnTgzGvlRpSMEcJH11YurGm3/MDwkaNSJtI+Y0OH1d
C7DavKh5OINJuruc6cndkUHLTROeC4qBjjfMSNL9gItUmRJJxHIiG37fkHpom5rx
FunHRznTza9+/zO34h6340qcCJb2k18jnrh7UTx/I+S8dpd4YtXoaKOjZnQ/WmzO
jyBI61aUcbiq090EpbYWSbLzKCHlv0e0M0HEgHWrnuiqgrDNJX+iUitr2PnMSZQR
MuIsgZ9OwQz01Hf7j13TiaQ0U7yGOK9TVItGK+U6J0v9AOBH06Khxo+dKdywFf6K
0y1CSzDvjB0dg9nk6SVU1KM1q8evt2cPl1Y9Pi9c8nliHrctARqvUGYZDjZxqLr0
z9XSIMZberbXteq2mZLlPnlWaukTdXhVZ3/NhbeAjJLKa0RAXb7s2xxjcj1WpYhc
sRCaPVR4xjjG4pE735PXNVbWbxIXFmzIUnApeL4olbt09W1qZeVejSRvmKuzYA+V
KMCvIeiYEfJT8m0iMcrqxjHmE2cB0USViOcWIrLycvnLCK2TvC5SSBDphS2UB8RS
r5peBh3OrJWeuT005JyjIlxpcAnFLzX/H5/0URAv+6+n2z0bdsBR+rwRTYG8Ot7m
qsv2XV1OAcf86UgH32wI1e5D8HAzzyplDjLgj9zRC/inLkTNElOHRrlfltclQF+l
EaxomFUEPzASwkVJ//gj7bRM2PpSPf+FslSuKLPJngfuD6kszCA+NwCMAUHeQE5N
iaJkY7mPZvNOm0ItjAva4r8ZZKYClRzVirOri+3kJs+mlBG1giDOLoQDzK2XrgaM
+VAnV8wG05ul4tnuDuaWG5sCSjU0VoXf/lXnS/KwRdOMaQn+CEYLsMqkE4RUvzBQ
CQKnnUoPj1N+CmKJKYjDedP5P8uiAhggy6HrmC6X4b+f5xxvvYcEsFRXLCOZGdKm
g22r74DVbJFQLqROXVb6D7GoTdXC7SFSKzqUojCjHxPbk3gB/ohdjebO0U05hkU3
sXQulV+tP3e4hOo010OLdURd64KCETSlIg1ZDPrjgHRXrofux08L1QPrQjpQpm8P
ez2+xNFq9vh7BZhsusR4fUkaUWWCr3HQsa13FzfWu1jVOdrT9+Djw7X9qJbgD/Ib
2NQIZJKHoou8y781nnGnuQANG9M6Vsfj0IAOsgM3NGT/XT1sdJk9qLsjDuClRsqH
fFLgEGdWIZ/RZvxd6SJ+PVB+85dqNXqYvBio3wvcK61B5TUH05iY1vFxmakh9G2Z
gFR8BPl8mNd6zMlkJR4CYQkF/SX17VBA1kKLWmhIJkWwy8cE1QgOVxH/JfaxN2ED
83lKrAreuJRpT1ebpS5YiqwCN2G6QEz/lWKR1xyIlgGiA+/BCCGALPuJfKJerOQO
wCLKlLG97+cxZMtVEAuBzJWV/EX7yurVRWJiW+ydFMmXlUF06uWVMT6xuSkZU+8F
QPVMEFHypu4TIav1/s5h4BSJAqympHH4J2d9DYC3JPujruO4atK51oyoLz0HnvZf
N/U5036Jf7679On1v9nRpWiGiBdgPtgMdYo73+27MIOYF0pVr7MlL9kPyz8HLZlQ
kLUcPD64aAE9nXJ9wP9A57FX9wCAm9QdYXYLc/Yo1NKIgilwUntqKRuAo7oTk5bP
kdjDhc/3Z23U2dRlC5okiIr+jViz1npp8kw0BWC4G4110VsvnwGVPwTGsmOKPItg
SoIYwLziFDQIJOrH7s87wYgzpoaDmjVJNG0zb0grg2oanBmcX8eTln8NjyNEbVqj
23o//eyqNEttpOYOb5lu6EGbiYv2MhbcaCwAwAVuBorGGx7dGBI8CQS7dJuUXyky
mhSDQWGNorRuzEWIykydsBhrfZ0uetLf0VVKs2W191NUFbli4Z7WD8gFnK2f4G60
lbeG7vzEjWcbs9BrfhBYwEwrWQ00MT09UGeLJX5Of2zvN9Aly3GvWm4iXMajEx2G
8kmt/qbq80ahJfQKhqPdNnKzn5a4uqqnBgV4aWzSAIJwgZdJlKTNvISiBeqhAO8Y
pQY7tyDJ5DxOvtX5/Ds0vL1CqQVgP3YBNmp1eornr5Uk9z+r4Pp1IP3WDUQuqIX7
BW+tFxI+nDlrTjmasvkE5rGIJhIh8ngMgSgPoyAmdAvXrehw2/KF7QgPc9NGVGJx
47GFVjGqF17H8J9OTTmOerSiss2mWgZwOyEiZZeJFXRX+JdNlSOw3lqqGJa4UGAh
CWxqPl+08lbNwz01uTjK3IoSo9rzTlNkrGnT4mQTolcCqFAqHgdahSEFx6YrTU/y
qbvbCNqTaUijbfGG0xf/7uK/r4BP6UW7a/EDhWH/WoZLslky3vvxkJ9npafhCoZp
+q/vw9fKec32oDsY2ZAczsYcxtirmg8BVsdIs8E2AHQanQC6vVRAtvXN2lJy2JO0
iMv2TfK9HYw/C+njkD4krdH+T8DIOeatJe37z1F3m0+0TFE5aj95omWcITlC39GE
0yVKmEEQ6W+tVO7Pve8w4DeKFbMnbsFID67ypo95t32IhBBhJBJzVtoUYyQMQm8E
IoH+3AAT8GD1inf/WWEvo+gc/xeqOFMUZ920eiqjJtVtGmwPCj+96PoIfQtGMHaq
RVTU1wr7oCk38vJG+FCIepo2Gi4YxGP2cZn21UMJyl74bU+hszfCLykCiF4P7FFB
1pqF281mbR8Aqn2okKCAVxiMKHU+RDnBJRBK7aTsAAYIy9z7ueiYUMFZ551QWG5Q
0hmeidtXMVlgjcdZPMWeRMvu7vg5wVV374AsA6haRU6+aEDJNptTyrQFGKMlavL0
H8C/1eb4VDvu820YBpmrpYRUqh7PoKbqU+fGaNHUO3m45dj7t/aqdmWiGq5QmUAn
uktODqji3xjNd3KgSy1rMibjh+wZrsHYjfLTGV3LlKwAbZMSWz0sRJBhyrpyzg/T
JKwLUJJvBl17TFfZPw2GKTgV9HyDfdkxcVJ46pGJAbsixzrMPxik59Zb/w+uQn+R
9rAGH1jyp3fWs1iaceDUnrdUK1JLjdRlrxEVQk2JGrNuMga99+6q9f1rvWCs85CV
/73rMugW7QOyrrjIhLegc2ikLg7WQC4LXo9SMQOuZLcu4686XvZGZCeLPF7aSdia
qpPI/vhXbeyHWfvB2SHTVcKHaNon7PAy0Ch6uSdQuX00SDfxDd4JrkLFX9geb3Cf
4bYwQ4+sz3YwIxAjC5zTI+YiFgxHgtoTJHc4Bj0qF/K3Q8oBAGLAKVUDymx+N/14
GGZiDwbmTQwTXfsjJ3a8jqPPcFODnoUaJ4Hfyc770yVEXlR99crA7bqjI0mOaScp
dJHAXY/iiDkmJ9cHnS28HEnJo35/yAs1YWxDm+1bNjDpqZNqaMRsVdE2ezSR8M1+
PGUs5JZqdlepbi1L24zxIGtbz3VFhkH3xFQEafY0qkvzgji5qw3vy0N88slFJbLI
+5n+pGolTWJ9/CqmH2UtT8Qqxyk4sgKbGYJdKSKGeX5JbTqYBPRdTEvuanFxwD5j
+jFhwNBR5WYGbNilz35QY8IA7CCVnXwjXc6s6+wUuHHyqbfbFTCe9qO6qIf5rFHp
wU6n1NwfuX5lUcvXgZHK+c44p/+W5ZXtqVbvK+0tlqxHOiryM5Q7Wm1wY6eFZX3s
qu4TGLHLRKDncuziGhxCCfOf1ezrpC3Xc3twWUhgKVbxmBsQFuFwauhSBrC87h83
4P7GXox+XKFvD+5HmNIXwAD1TQm0WtWT4zFj9p1z441HJSbldP3XQOIWM4vUJQgT
5tDz3Vbz2M9CfpUkxYtwBu5crxJ12Qk24r2f1Gq2k9rRvoiYBhxl5ecSHtt+Sopk
y2HPVYhPLA/g+GEjq8iayHrS6NvSqTePIUkdwuX4YxBgvmRDk9iX6SKQZe7PlEz/
5+8ksp157lo+sfR354Y+rFnSHzcmHp8U3CjSJK9ZlgIm9rc6qf706E3rk8DzMRC+
N8kHeU9t+7LbRiy9RAI0h2CPWUH9jhXY4FS2Fh9bAaXdWKoPJwBnk6zfxgPNvOg0
SMIfuTAl7xJzvCdmbHFoqV/2Brhx7kdBGoicBivd4oy4dw+IfeslLOr1aiiZdb4o
zZqmwdykT5YQMA+SzKGHQj+Hd6iiqI88tberih7jgXT/eoI9H++08me43xBvk8Wc
X3CWnirE80EMPLBnPYqG7sB7JLUkzVaNg+Obwkm/qWuylWCrZWKz28w5p0MnhmBb
RLVZSIn9sno78epG852Cn3LdWZPdZ7t0/RwkZExuCcN6siiYqjzJFRpn1SnEppmC
nU+l43pzuvodhfku7HCp47v5/Lq+MIm8Gb9XyKhyc2abi2Vaql5ToLWpMTjjIxto
/+8gM32ZMwPKmwZF/ZVVssXHQC93ny7yNMbSEf2RVled9x7FJ+wR4tCNxQf6pBm8
gMIyZNIBkzeEAFaddsUVzCmJnTVu5WZxNtK+5TwGb0jPwiDswK3sgdWyO9QWUs2w
MziXy6gwPBkDZ4vFGPxByu/EF2mzxHTah1ooL7qUM/KUpP4cR7v1EuJ3vi63XFYa
jRrrcXAGZG0suYYyVNOgq9KStMqCjmb9uklzMQwxrBWfMgOt2YFt1+Xb4n5XPdg0
Pt7jXHd5RNjOkvTaGOnRDmY5RY7y2wP7goCN4PdR/b6olcbpiH2DfTD1Ptb2b8Qw
g6lRkzROsMbEnBLbOaj1XQbuR6hivuCBe/UjJGj+ZNqPV08TPW8CeSAv6yJ3UCTN
6FduUryFpGK+Qs+ArXacPuJTx+9W6Ae+vQp4mK6NKShGZbNuzq2irQZQmIR0+tsE
vbDpjfHGGl2qPYOj9TaXT43MbMx11nEaiugDQkSTXss1HsFb6ZyQsk/jp+s0Utxv
U3Za93NH/NIvDVVbdzIN0cqWNybw1F2um6PBy/eaBmzSAIQUdMsxzdCk0BYKAphC
BEMPqQcSgrXL94+sqoqy6TzfRhQNgnBkxHT9m2toKQhgWkQGqa7xiLIcdcboMuzl
Bdv/u/mvmzmvpdKg/IeGTzS5tJPMtWJKjHMnzakJwCn9qGa9XWQqcBa0k+ceKhqy
oXZiuLRt3bHUfn0nHbp8fjj5ctTODCzJsnD6a6pSpxP992W9YRFpLUB/F6OlmITC
QVwtFTgXlthsx3sYBSrqYUvZXButPlT0fNRV/QaUp8T82mASx1UJ3pllSrIlNaLI
Ax0gZ5mAgyzHZkdJ/cqIWNAIHjgrwf/GKhddi/OLJRQFgIgZcoPBoimOr+Jr9qa0
9j1I9/I8DrpKbCRFpZxosEwSzgo7qh5rfRc+pd72AyoEMKgprUpXAjKWlbaPG/41
5wGje19ldlGF6GAW/OIX44CqislWKWHo1XXlUu8xwNIzghSF2m9k4JoN1mSfcNrF
5SoOu+9TnxnwVYeJua8IX0wDna82gfVygndb5OpVHPdZvwbbhQl1w2zAED5j7Tv9
j8eiFUpzk1dFSkR/PcKYWXLiG3eYl6xm/TbGiQZsVG6AddGkK1fs2XbmazSfB/tH
/R/5QzcjZyFtdJ3qDpoK03vxq3oPsdsIuPWNbywW2y9VJ5HxH7l/TLYOh+cSuOEo
xgB0UfsmsQl1M7XyoqgCrj8BxcNqrjOusdqFI7qKzfQw7Kr/+B0E6M8esdqQRFlW
4w+jqU8yWhiE+9eM4I3DKTb8QGaaeDWjxzWcRR1rzh1mk19tf35OHnV7op2/1GEx
jCJ8oBQx9M5Y5d71EdEfN3fq7ukr+g3Ku9BtOm7Uq83xAjsu4OFnfAVbunJ2MBub
tFFnEurunXzjH2Li0ktT3kbwCkRPVAO1mTxGzTeqoaZqSSFTQG1psW/ocHVr6MCx
V9h6lNYImfwv08knsmeJT3jiTs6Rl7EvVMXEsxo5SSkfZtvzw+zztXWBqi8TfBXY
cZDuoAUC5/wsD/ooUJ6oKyRGvQW9QrhDl3r9sO5Ms9/1ZdHJhGOcYqzc2goMabZk
VPQ57ejNMMYDGVzBnMSA5emTXKEqT37NUqKdV5GcmB7z2eMuoJDpxpUeKT2+kal4
OyGDC3HKXi1Jb0E0kG2VZz0ntBNYkER8HA+5n8+HzRejCHYL/ssiT3n/GYQK+zT4
PxKNaxLDtfKGYWPodvNdQ3aJAq4+wg9aM3Cfvl2+TIZHME7NyRh9a3eZVA2un4rv
6xYc/ipqbW4Kfi1YWBtV2luWYu2/PIbz7rv+HPDi0KPW5fPOpIBl6aB7NXKFAxth
N/IaAHe2jIANAO3nKu0cqrrceV30gLSQyBiczOT6a4GFN8Y3u4dGu5132k3DGh7T
FJpztHhzNY3Fu6aRE6NsjwY1O0wPRG6BJoYf/b92Q1hsYvA0dEqnXB85VhlhG3wl
3vS3hl4O3jM1eZ0JTCWJfaYRv2WSYBzoyJhZEacw+lQo14YSiRw9f5PakHyYnd/B
hI3gXEGMQF7hc+oGJqQXo30WzetvUGgw1JmetERYm9WiLQ/PygTjqZx8DvlDz3sf
y37UR49a3n334tsp9pzbTQx4ceX8YDD2dcP+FZigvpgWTwTZ4AGuQPY1+oLlBdm1
4Z+hRgcslsOzic6BY/kVLu8oWQ0qfa6jZcWOhh6bT0hONT7FJeWhRN1qji96AlRz
BIO+FpCuyfKp8Fg0hBt73h6NrFM7UOEf8Ut5dIueeWqFFuBElhhi58o0RBYXf9JC
PoAZCO6Kp+4GA+k/Tf6XpetBoZgyZu9PCve+n6rAqTKlMTdQJFQ33gaXFS4R7egV
2HouuImjgeKt3Fu1F79XtnWBgtS8dtc6pEOvcIjpDQR9X/IwA0Q1LPG8HU+RxsCW
sYtREqfrOklLNRfYI6CPWdrLnZp8jR3d8zbqZxjuumL62EhfUgu1ExOjxbvdFgRb
Sz39v8Oh/LpNSXCBTtp7Y8W+h2JRohe/j6pY1X+Oc6Mo4Vrv+IPESIXDhCr8xeYl
hI3eUpMZQYNRT67K5uAPId+mzM3Uxa+AHeAlRFaN3ztl42YKepZmcZWOi52MaKLl
xZHkrS/HF3MlTE9tCuEfhzG1bW3WVgWJoiQbWkCgk9Gm58kaKytf7kSlL2qA3iIL
Ao9yq5lKzoPnH+LeP35F4QK8YQD5LsKB4lpxsuSCfEwb1JQwx6xLYVzsXOiQGAAt
T6e+j/XDdSVO261x1QFih93g6RWMlX2nJkA8ZR+bYY32XHQYqbmRyrtgRD1zHHxU
guh+NxLIcgHkQ6biLYpquI12ZpFUfTX0lQsmCcooHmhZEI4Q6Ve3zViBGoRWEFIj
i0AsDJU5EFd7pxelsfX0o/kTjxBzI72lp/nnixNzHJOh8KM3bbRRKkXjQkSREF2+
je6XRxOfT4SqAZPQWq08rPXC1mkIXiQ+K0Nc04goGu63d5Ss/1S4ABWISdh5jj4A
Brtg5RDOFFP3a+UJbAfWSe73vM1nCow0G/XZFOfu6fqJJsfZyWWvn42Fh7s7MzMb
OAI0pz0ds0BCuz7k6tFSWJ3qNbt34v4kPzg8MA0/cV6cyLjZM9HBN6ccpw5u8uRK
EErwEY522pFkGC86j8ZEAZpdrxwLcHFLO2qX004jG3NmPIdTD1jL+H3uUCf4VW5l
hhBUmtJGsMjCj9C2QvWHBcIyMcLCKWR8mL4HyDTxc6WYdwbLyDEgdAQuJ4bXiDxF
H2Do445b4C604eFhFDNlQjRNWxVPKzXTGR73GpMjFBT5fi1zPhjjZhlUsvsDkLxr
oil+owBZ4FPLn+OgX++fnPY+PA5y3dIJso1JvMK+swMz+wBHnIhmDCKL4g15IBmM
vM9vP6MzBJ9c7m5JhWmKuDlB43uzuBt2hvXIujQoWm7P22ymuHT7MhxaZKjfiNSm
0O6GIFRmI38SU+FXO164CLaqLHmJW+Fgxp3zPOZSr8p8iJ5a8PC5JtsJRfWwp/qB
f6cuyRQydWl2U0y/3/taBUZ3fFiDsyXXQSb3+whP1nhEdkBchgUrX89gNA+UZrUQ
ypGNIpmxfYJmucew9vQzru40m+ljuevI7heScUpaW26DXAcQmvaPzQ/w6NOJ9DBW
CNVIT4XcCZUCCjaUEvnTQkyO8wNOA/UhK0Vkzj+rRB2IZ2ZYTff5C5FenmMjU6VA
kfvj3QywFyZudzZ8ClAfWMP2f5LK2ghrpNyXtKpRIc7Lk0C38z+VzCvU7yyNBmmv
VFHuhqZinrTjaRKYWbEIzJUWexXHoLTQxpIwX8Xbjh1QieU3jTUep2HglSBwxt6V
f5wRqWYIJokMzZ1IGxCdNbm1r4Nl14OXWbDZHnB45mWodyIkfdnRHwwBBaFRXUmO
0shXvRtxTsrf0S83N5j7oj0rwyUZheHmAXliNqqdYrEjeXgZ7HawrrNsYlD/1Ktz
CzvUsWFaxZ2Rg6yS26/K7D5FsoGkDGs41b3Tbaez3uEDHuXwy7PQ0SYlB0gHVtq6
8nzeHD6/T2gv2VM1MsdkhyqvHfmgtSNjMAqniICZ8fuOhvNZlqasE9mBgnrU4nHR
HfVany++BUzESvfUYOhMb3DgObABFXMb1U6AjimH0ROtmw1EwabN+M0BZ0E3Q0Ec
eqBzhS0TJ57cHMVQV5woLAHkSBgv0QzIiYUhN/Kb23gE9luNf8GTLf88v+lQefpP
AnTwSXB7Egf8+h3RhIgUrzuYM9uDkWx0kgzpAWr4FpbjfEjzg79V6PU0cprLQhqR
3EsykP4Ds4TPDZFk8Tv7XtJnzthoQMkboqX5lFCkgJTY685RPORMYHq1rgFnczNj
U1RGOa4b490wgfp+lPEzpqynZpGX7t+/8/avTRJ5Z4W79J2qicfxkE0ME7/UnJhF
L9Olq1iWPYJJM36gEq+orma+QYyjcdWQ6zB8SeUDFKigiFW9Fz6kVB0qv/rou8tT
iA5Lk8VUDxwhSZbGphtj36zRUNhB7v0YaQjjO2Y7W7TAprCjle12H9uK2K4383Ns
uivsrUlMnDlfkVR4c8Upc52dfqo7P2qgHjJn5kL6HQK7raydFF2olWNFg9xQ9vQM
pDxEqHc4HobLkwD4zzaHW+pUllzzucubtt1rnwQVrY029C/tD/EIT8WWg1mSNqW6
WKzqA8G5oK5omZX7IGBAmebNe29/UbXUqXzjLOzuqHVDf35iVGniT2qH07Fewc+i
qQk5qFuNIGVThV3+VeW4V+RxLKWtdC5S7rp0Z+eAiDY=
`protect END_PROTECTED
