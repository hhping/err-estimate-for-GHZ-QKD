`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T1zeKLTo23L+FVb9tcqQQ+1iYXtP7q4hN9Z1tDNvqsfYIttBJXJnWTwHiGbD4EBB
lhYwv7se0K2jIm4zhO/EhXC8qw9nEDBRAHO1K8BQbCagAyB+jTQpVGurx3BD7ZGO
F67zAAiCvRSajeUFeCntBV3WT4iNw+2h7bccZPCADgGz+qAhZhydeayFN8kLA2ZS
SOF/Ra7ayam4Hzrr8lIrti18uidQb/LDPHsOqGlt9D4qmaUJ3yvFBouny/W2WcM7
r0P54ENNRF/myEuQcd0+HPg3ofU5FZHiysk3rEszgL6fHNRdpv0T/jbNT17pUpkO
xFqIU2oTwgMcmSKU7aMil5WKkINsZOEt1oosgAJdYwAFdoAwtOSy3x+mKFeETdDP
+JNFJz6OcKY5xYWW6Dckr505bgzkfvNaNs6gFTvgD2/egtu7SqJfQLVB3ZIHzx42
WFc/Xeut265zRlRFbrb4EYRLwOgQ3XOL91ax91g4E7QxzHj03kyhs6B1m2c1ixpp
gKeyG/Dgyacga2JNIqfZhjv02vT6RVh3s8aTG4mG6HwOZAwsw9XkTvIZF8Da4NsM
k2lbYxfRh9u3AJzvk4aYAovDG5iSoMxZqY/mhHAmPIPxVi3dXsv6q16dxVi+qfLB
MWunG2ES2HK+EB0fvjrVbcM6xKW0mCr8RHefNjyQ5wwiuabAMODACmf7Hw5Kk/DM
oFu+aILFp8kFPedUOjMiSBZ9jb45odC6egM3FopR2uEb0r2jwkWjWYUjuKhNa6+U
jo4ZlQSvqfVhpOJA5YRrmw4vvOpUf7cSNQama5fnzUMAPG5JzMZVVHST9m/oJNDW
`protect END_PROTECTED
