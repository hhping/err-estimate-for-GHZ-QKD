`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9yz8/qmHcWgbosNYinZgtTdy2O5AeE9vdQ4se6qFmt/ZaQuiqTBU1bRLfa9bkrw
GPB/RzrMjtSZKcKn6Dl3g1n4S14chbzkl2ay3VPpyS0W7SbtXlZ4XccaWNjIseD8
0mhVqo0KxiF9bA5o1DR0GuB3W7R2EVOMv/NBnVtc02d0v0UBop5SpPbArlmNbCoY
8yOp6W1wh/pLjc9jXrQYkHzx8m+jDQHUxcEDk+6LGpM6DC97YT/V+sqBvr0sRx7H
px5r1yfAvEj+vC/BLHB6kDEck96VXMjNsxbAMTHKgQSuyP1u5x5PxY+YCfUVgWI/
iBeqkPOlTTo4dick6xDZ95VUZHMYz/RCkag1/imnlFLMQ4pwKulDCt4KFWS+kHb0
FJpmbM+UEtxgVeRY+/qkfre+4Ru2YGfdC2uNwgG1TcfTDzHVwOtgTDnaaYGDnkJK
Fc8YnOGC3lDg14zns/z7v9uk2wQoMuMdsQoZKg6joAW0PeF9rDYdqZyCFPnDNrxi
gbTQfblXuQ65cIX85FNulfp1yWbJTpOrzH81Dci2+X5+Zz0AdxLOhFWNM+FBEOph
5JAOx3didpBDfAVUdIIuHhHpVXYlW+winlo7IhB9xzIFxyRCq/Gk2D5nMKAjiB/G
lPubOjjTu9vtShv1NBVlMp1JZuB8wA0cSe8nLiUVOdIPvfRGVmliY+8ICpA36Yk9
WBHrpC9C+OuKIBuTBEFM38F3wtvDDQGuUxMc+T2+67ljDZyiLX7i0MkUGYsYdDXK
oWVg2ZiBwhcuPcS/U/uHI7AJViQAxltcPlwtOiveKk/xJzK6clXYWJBVrO/pADne
kPzY+0MSJCnj+nIkcVTt59Q3Tkl5E0sbYqpEQb01YbSBkgOw0m5rddDgoYLvVOZu
Da2sgHTZUvavnJ+iVFg965jENqiSqle7oNBzCGcWpl0dwuY8XhlJGVMvxDGpVDZP
0UxJKInTrSXxATH0Gro6yB408QCIKnW83mQBXuIC5IfO6GO+A2YemRiTQ63c2Zko
U8cuVyEM2bDyLKAKxZJczvIqLZfePlQ0i9ekkwLLJ2tEckhvuL2HGrhWkpfQ5zCi
fCjHOn18+sGfo1tMhX5cJ/q0PruqYOZPwyx9tJMZXan1koaQW3tJmpkzjCTWmEkS
Aq8tc3QrLjFWmAW3UlS42wq2SfCk2l/a5PI+pWv1XI7MxCUwESAPsycDEss/TpYM
AWvBEfH9UEFlfEXyWFMFnDJxVF2kIW3g5/T1N8iIke79bLn4D8mhec7r5P+BJJLW
nndmp4TfJ0/irQI9a7k15xGGTJXZABrygjHG8/JpB4iWCFLVzkxoOkeE4ZYSojC6
m8Sw7r1dzX75Ldx0V3fhjgF9CQPlTDMUvIQ0oQLxlYvrnrs/WvZ+xN5slqAaWjkp
EK+G1bOFSbRiEYUYDojbKsWq68FV22YQf6XC30MzhQUhGz46iIGjuuCageKlanAT
BgALDzTUCIUa23IAW4ne4W0em5f2SUw9OtRHm12KYYOawMhFEbjjUS2PGRsvKNnY
WHkRFDcUGT5TmtMJXW72VOpG9o8E776cCGOBhlpB2nhPclXCekWjZOQgbe7ELKAy
/PgIxJAS1j4At9eerTUUBwntaRoCXFwI6BvMu2xLg7OsOi7cFK5F0OsG2CaubtE6
ZdUhre29ZFMYj9nDlchi5A/rMSX90a5cQSf24DSXko8Ajn4tkjBeydBbXr+IfPSF
evmFKfzZ8f1UntVtOG3v6DfTCaJFITRiGVhOI6ZXszBk0/odnEBt1MRGX9pFunu2
q1hGdjQ4JhBOf6qipS7xnEHxUDEWQBDldgZxEDtV30zhPRtlL8h+64npchBXH00N
itiV070aFfWPSeq7aCG2HaOWcMwTR5u5zqDxrCnBYIAoT6Fd5o9YQTZNV2+XfjiC
R6BJ9XomgGFP2it7+P6u6wb6eLyVA3fOBiGhJ+M7sLNHuYcx6JGrCG2vX5F1yHGr
YlxZwUKqls8aB23XEtMtlEilW2tjdQluB9wHXAbhvKtfet7d0JAkHwKA0uO+PMt/
JjByjx8PzVdMT7uHLb4hWDKSX/VWYfYdNMmChbOoFgGoqkkzzoNIv28UA5uCPXe5
zurFcm7Ffe1olg23V/8UtAwI7BlpJU0sqczwcF6McZc+c1mRKYw6qkZicC0ik9/H
5+WQJVvC0N3KLjBiJmAUlSKqKWE2A5+PjbO+AxYPgpGmKh6BJNFOrERUoDOvuY4E
15BvsdZfo6nVIpJXeaAloSy2BgeRUYVbYO7zsxlThPRWPsSCMVEy1EX7hEMa77gH
T57SIEXPOLRXr/ZApMg6yP5boypRInF7wfrhnkTznoKAaaikpSUlmurdU8Ont+iD
wSs4LGIOJcwDpgDdwDbstEL/9rHJ6GjOBa6he6f/aRBEWaxUZxoyno7qh921Ehpt
pBdid/KUrEzTBBKYxHiY4Bu378cPmb+53Xto0ebn3jNg7+FFVaXHy00+UZ121W/G
4Dg+Na2XM4EuKMw7yPIJXUR5x775chAxhEsTeGdOIXVTpJeOGF9d9guATt7sLfv2
67qzsovc+lzG7XnvtxX6ATbc1HTOA11hCtM7y37w0Kg8BE+27snNeY9DNdA/m0B1
Bu1TQo3EiA47XqnlEMcRs+Yob7+9CW++j+XsX5j0kfBuzcQPyZ8LM0BHC29WabzU
TpO4wNZphORIhC/x0SAt74nm29JSv33naxmAmgw2osWHhl8dSCtFLrdB+CPXIQdv
00QlL023sTT/Xzi2QFF5BVrSs2lFYcTyPwkzo5gcsEa+Y+7yhWxSjapmjufwbsN7
CFIUNrMax5+FmS6nOqng7PNVHTodA8Tm5TYfJOmvHttyZsHgQvGJZuFwk31rQGOQ
u6+uAr2e5nPcIoD58Q4MA30gZ4wImO5HLsBGRiDhAHwQU8b9rui9UuzIChuB4HL5
M32qdTAnmogE9CSO+auJ53s+yV+lukSbUuLGzKJM08Qirv8RKUlOqu/70nFzQjtQ
`protect END_PROTECTED
