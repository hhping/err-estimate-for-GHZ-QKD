`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlDXZQuuHgyKHeMlx8mjSoJIU0AfN+TmFBL16DROpS0MypuYbJd/pvYyTXJ/7jId
G0aAZBYI9j13wdQ6D+BDy8y9YwObJfxqqvKNwh49+e+xdNpaqYGHP1SXbLoE0iB0
ZmS2kqit2zQ0dboMIo20+JEoENS1UshzMLYxBU90FpgEqh2tl0G5hO4TkLE3FwVX
RNcYy7Sqf748hZCK1nFuu9LcJSJJ0L5s1RKrn8novnAbz6r9MWhqyuD/VRPEVucy
x+FSdjhQo/mxMk10j1nv8fhvpP9bdBZ/OOAwgJT7oZRXqG3KuYdTlk1ZZpkdJM6p
QQWsSUNICe8J+ugWVLTZ5GNd7RNEtU2mwEPhT+a1um/xEGIgDdss9soWy3xwM7Pd
QRkSt12O4dbDECQvbKgVlF7F8A/4C4TXs/ofspGlb7dUXzxDnTKYZLkj3LXaNffe
B2Hdh2Mofw9px4wlXwEi4cZKItUr0gRjF1TE23h63yr6dgTykZOyjhbwlFNAlfE+
fBokZlBh94OB7Ro9M2P8M/3bOnjp172nF2CdmqSQTRxD3WNnPQvkjEi4raQ151JC
0EtAkDsElkMjhFFSZbTTAxRzN4sLrE+LFOaRiIrXfxNwY7WKHmFVZ86wFUSpsli+
Kn8wAf4EdVjC8rzAuF9ybv7ZBfEv1FqoVnjohNZgOuu+G3kVObdgZBfsUOqCkYw8
sjRkKjJRGrDz151EYN/tB0Q0qBTHka+bleh5LvNs5+sqx1i8hTkrXSJ0FNry8pmL
Ai+4ewYb88SxJ+WXKsMBp2ukLfnf061CO5EQ5S1Jx5ufZvi24N/12KMp6NimHFD0
4kzVtOTLhDQ48SVuV2jGV8fhEAsMb8R0jKvCud5QdFBcTCvWKXhqqZpwXpSlp0KR
DslfsW6nS15sv1wPqQ0CGZ5bzrxisKKiDyqW5vPf9UQc/CSQ6v99XaNTUshvzC92
GLGqynIBUAm+Xeflva4PdfOxBoKUwNazRZndLLn1WqOO8IYG0E60xWhoV88Qiyow
2WzFoA7qFlq6GLQ/mKWNk9JBTM69IMeDThGAkC59sZ8nRIXFoglUwSie3ozNmdgy
m5B73Qz41LOVnSsP/wSyOGp0qtql93afjX3EwID2stqBGxcqCnQm/0A+aE2ib+XG
XILXS1q1ieno/pPsIs7EVzvkF5VnrLlT0uoMPvRcXAUtAI1ObCuaYrojp9uUL4F1
XHZ+WH11XQow1vSXocOI8tRK6MfYdgicPlDVBg3gUblget3d1bXvUai3mLrzTYl+
zXYqLhK0PVw2bATTf8WIhwD4W8YBMVzft0xaCqSqAzJNQ0rfVFc6wbp25qr/T7X+
DmlCo52wDfXnmwXNnzLyS/elJc+LE7v+TzWX03T9hlGFp0aJG2IbjG+Kp8x2afDs
fyBm0bdinPaE69NCKE00vjZwg3YtMckkZZ/05a8ccZRA/XWLM5c371aGzwbuENkf
mx2udUnu7GYIOz7CKnSSQ9J0YMfnCaYaRbjRSKLpNJAjXHw9HmekEPd5jGxB/cVy
7t/ZgVk/9qwSjR13nh5m7Q==
`protect END_PROTECTED
