`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDbbIjzSHtWaNKF5oI4ZMPxiPByZEKrY/Q05WKXBQ3ufgp3MVrA3BEFEB+SbRbT3
OHHHJd4R99Y1q9pUaWSRhkh6LkOKhswD03adP8AWiE2MdW1uKSnQ0u8pvTQ3QznC
D9F5ZnuTbg3x3RPxlE47VpmXzja3kLm+72DP6ceVmhLoMMb7iW5nn+GZOPzJn/vt
EQ13/o7u6mCGcjB3h6QKWkYggJF2Yt6vcWSX/U7xNLKDfbdSXK8HiW3lt0Gb1LdX
NgpnQgqki53g8NOfvPpgvte0E3ND+y19ppxGNuE9RUqqpRAd8cVOceojjTkin0YP
WcaVOl4bhgWZeiMtwjhlfMy84jdadqpJvnXeyUDTjWY+enAzFhpw0986pptL7sFT
hB47jCN0Jp3hG8Yshnpn5Sia4HYhqMb+T0Y4duiraYzeEf4ElPlMoE45aJZe4lKT
FJN8qoyyPGVHyEqisCIhf8hU3656McyhZ2VWoHQy4syxqKDzotWFHCsCFAMUIV/2
IFsgqjbwwDOs5ezJEpGPgQ==
`protect END_PROTECTED
