`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYTVoOLkxDn9jlPFdgJ3H3rS1lyzo2/ChWrMv4UFlutfB2EJ7WTni17/Mu5tDyDZ
2uC3F2jvkzq8TylYQTI74Eiv+Ux9vTqfB2JfiQoHNJUGFoqTxghsOdMXZKOXJMGa
HAhSFUVGoUjUXu3LnMAhZSBoVT+oRp5zLYBqB+uYEy2CHR2DzTi5Ox4BVJDvWqjt
2F5RT+E8xEI27x8ELQx+tJMoF+MjU1BThADa8DytXnLaeHYdawo1V+Qe45HSkWuU
HbAI1CTQ8F90huqdBuqJIsypbi9d3Ur9zh3MObhPfyjaer2sixKRL9G/KHpts+Zg
3wZDpQXiW+s7tY9gc9XHTl5nh7BZUYylnB2OEN9zSB2l9Ea/KQvuPLGnzSyCWZlc
VZXghxJFW+mCO7kg6AXDAtF5iMaEs8QU4tBNaYRSquWnotqDsrVSEsHh9dpViGJv
Y4LmGKR2eh9K+/Q9siks7pLacK+kg1plzDNA2lafXVogMqWW/Vta/iC6gTbiDD+S
`protect END_PROTECTED
