`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mELhOKwL9mQWQWpL57R0iSpB87OqZIJYoTEWbNznDqjVhk1k1U/MweIXEDO27ln
9JggST/uZkL2quoA0ghA26+1lEuFqQ+4cTbxnt+nd5U3KZeb5gR/GA7jrz8SRhbZ
9QVTC2dxT8HyNAeVdntq/VrZZ0aMgg2kSMaJY9y2vheOyeGT+Qy1HmwWdDlvKY0F
WEojDG8eaZS3CMonmwkOle8PJpCFWY2lDrlTye06kX91N06bPVeCkC5C11ZRqibc
9Dn3cjEaQQusY+6eGlxsAcESlMSiccXnnopBsxYIn3mddmlKgCcSGLQ8EfZKpB5f
YHUK2MTtxrZcAF3wDdKYibsQeqHmloWmBPMgBTFMyQP4aQzisn47fIU1VM5kgaOe
DYGvQ5mPwrep3265BF95rbYAvAPAjd14DOPucH4gewYdti95oUo+4DLiBVZZG+m2
CPZHlwt4s+gjdDHncQV46eIGjjrHtaLtBarJbqPP21vdvK0m/doqiY8h6hQDjcne
J6D7WdimoSBpRoReDmT75HaEbwEeMzJOFJqGLkzV0VBMw7FR7VyrVGXAy42cirg7
Bt9FoQyCJo7MvH0FChfP6YZRwNu64RbfHLzMQqVsTZPeyePSg6O22Y0JjsGp/89T
CaD4eu8vs8BtbGm8G3s4S4qSv/kZ17WPIFoDCtJt1KDj505pl57whMDii8P2pIar
6uauKQAWoU3koKnhC902DD2J2DaP6WqxCQQKbknarBWK2A5c33ptGGLCCc4Zs/fs
eZ9otKtlDg9HDKqyoVIQoHzt5LI5Gz1QrE072wZWh/f7bN0mDRqk3sxBDLfcy4Y9
K2iz6DOUy4PLNn03/Ah2/hEBXzhT35GeRzu3B+M2h2ldau75niAz8rFHj97iJEDW
U0t9VCtzllGHw9fTNgPBNbeUlGzNiv7fnNiabx5pkNkuUuX6FrSq7GekEN/Fjlob
89YQ8DfpPetg0ItFYsLAkZAJkQoMyRSdTx1nh+n/2rIKUUL6KMIW/A2EE9FNxEB+
EHWnETlWkPbbDX8BYG0iRVv50wzQHCbdC16IzxiCa5FVmTq/HbZyMlQKHjWvGzWX
irsByEGPgC85/RXskovAexDZDjKte2rtsx+0YcvX8wyrdBt68SHsNdY+VkwLrdfG
I3VDw8lOjpMg9J30q0iI5s8RlP030niMkTVYA3/Rnb8dGRbj9DoHUda6pS7tS+kA
fCVHhohOlyncPBcEvtrjcVHQg75kCZzGDoUsFQSG7P/Rd9tLS9wtt3YAgGVQ5icM
l88Zu1xfeuf5ih/7R5Uy67UdvusuKJY+ltgS062HHAxhkRlUItZfIaSun6Oxl0Hy
qERDJ0XMhJ8Igb2eCXi6LauxX0SWfQzRICYWHXHuwZHx19HJGqHHzlLS9FQfU5l4
RzFGIpxXKGEko2UP/5BEGy2bRH1vS8fOt9bR/b1k2j8mnViTIdToZNv4x5+iLI9Y
CSA+wVRDy3DSX45oDGNoE3tTonSEOgDnR6Q3UpPd8YE8zMTMYmu3MOouAq2JqBua
Tq9OQXgym2nWaUPJh+PorC0uYPsBqCOXJj6C2Mad8UMMNagPFUDELuELV7esX+Gx
A9PQfwFHkSBk5n7EoX6bLuG8Ls8IgTOMkj68TNq8gYK4R0SpiOEc96ZbR2OLDz3K
i4+nSLEnOMyoe/S4bePhviDtW6NHvl2xVw0eq5A8uuBULipD6LZTAR09Raza5xnA
LGSqKk3ecs6GH+EfGgKyVnHtW0LUX59EGBu0ZRPqwL5jSHa/+SH138vlxI3mc49c
qi4m0SXOukBUT5ysdj3D3ejvBYX+O8L+g8vYX6YwTEQ3Bg0O6JMq4tyOdjgodSAC
WwFnFw99hLZFa8Sj6cbwMI1AV4NcnEMwyHK2NZvLQqjr4bqxrCTsvosqALJOyS2N
jhNPePLFd/Ugsg6RtiywZitV/sjgY0Z4OLvK7rTOe97RII0CJgr4t8zQPWnZ3aUl
hvDWb8IysmjBnQg58O8VTpjzmMIv2OoD6eSZ90ELm7Jt3xDb1XyChB9r0w6UJo93
t2ZMpVyDP5Vj2TzfXHqE8zGD6tLdSA9XjYrs+KArD9QP+1dT1M0GLf04WqcySOCv
NTQekGKcefXjTKQqFNZ+lNO3PRf0WDGxdMGy3iZvae8v5eqVSt70IdhhSEiKaq5h
kPM6QX8NTRZEvbONyh2XBCvTnSBLSydtIFgHsAzxnVkoB47EIs7grjPOEH9Mhjea
8R0RmtWHIJ5tE9KM6CHygYJz1tPWtu63E10vdEaYWrzPfKdZFYRKVuQyRWhcq0O+
y8Hic7m1gJuZFhbC3JgZ1XL03pLpLRn2cJNZBX3HB84G1P5RBXI7svWlvSE/UGtR
Y7GAdjGzx1FC4SodGM9jAJzzTTH1Xjy5e/ioY6qG6MeWN7lbRxGHT6ppeK3Y46gl
4+suWpMh0wUwtCHAroCbXAIGCWHJbVZUx/4+SHJHcW8cACUdh1fKUHWYlq/lf1Fg
WomlONyzN5p0e+/oZR70Qf1hdUezwr1GXAfOl+3Sv96yHg6IfSeh30lanZznMx7w
wMsOCgCCusgDu7ffg/nfxccIdSqsutMHkcis3UJDB4RkXGjj+dTkA4dsV1028XDD
RNzHZsdfguFjDkimq63wB8LViwIfwkgevn4lBGtrt8ynQqGJvXaWhLFyybtw+oJd
NH6xHirlj3u5+f/JlWtN5rykb3FfS0aLRJLFvLjE9w/w92K9moB5YB7e+BVHc3Lf
tbtZt7EwsZ3up4lc7Ja3fYbymPyaHGqgsB1Lavrqb3cXAUfa63FRReQMyAJeXL9k
rWmeYYFQsN555z4uH/+wIOEQl9q/06ZPGAj1PLEWqu2Tth9WAu1KMKgxAuzO6mcR
npDy8+c5aIfsqh5/iMlCsA==
`protect END_PROTECTED
