`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7zcY9Hkqav1wzbeZn0TnDls5cRfNn74GChePNbPuqsxGmsbYwHCIH2WimshPovfE
1OS00lh3PQCbKzAn03eIiNkKF7Zo60OGdyve89uNS/OS8LVblAvPTrSbm9pa5Wve
I2nghXP5fvMJuX+BV4dmqYFWwPhkc/gayH93Z3wDhKU5J/qd2rj3p3P9LhN4iRfo
D4A41b/amySuzATTmqUIuBZw1m6wSbomJDOLQOOxkpoCcd6OadIYqPmovGOVr1H2
1avFbNMFtyXFXsyyDcqryvyAwtcjUQ+4lwOvgnlvIHlQAHRp2w8cXd2sNEEM12+i
b/gLkb9zAB3lgtiUM0McdHjAo60dfUYb5tsJMocRLbVOm3fybAhT83/WnEnLkc8r
mpwxyoVHyNBmbaNBCFqTO13WoVUYpW72kC03pq9b0MrHOIWt81ONQKUUst9OpRbq
qmRE4Z4TQilottRKG79qcgPb7X7vEGgxhp5DvG0HCg3dMoOnEfh4Qh92P/cOpMAC
M4NCOd56Hp93qW9FXTmufQXCRFH8VSIN/fne21B65TIvXZJJfMxWx72A4qsjc68r
BVPRZTmmWePsVu3+UOHWFmSq75A85rH4ClPoaEw1gTuTByrsK9adKiz939ZZRGHw
W0yU55CQEM5+M30w8PXKNL3ZSgGa6TdT/Ibdrlt5TSWib1uiGi2ZmyLKpNvpiRVy
zqBnlfAizdArJuo/MDxE/U6iIFxNQZf4SVFO1CphTdigbLCE3Iuz/eBHiC7UKla+
XzuN59G7mzxXRpQ1k0Xt4GaPynHhMJN9jsz/2IxIVvK30Gzjet3FUasLUpE8JsCR
xLNEUiJPLmCIoPJGm3zk7jnfNF8lHmX8OJxzKNhgqAdfD+5UEGrVmNlBiFMFyQly
0mQnM847eKgPfKpRAYiwROeOQ4SEhYaDWnFXF5duqR12e5YWhwbm5DNwlNWvdihg
f6JMT1XNWFovBObuZj7icyyFCixay0CLvpmEZ9qN/1ZFmhxtI2hcTtXrIpaYdBD8
/0JXDJKb5O+xP6c9FGtoQ2f9HN6mPpsXppZxtZXzzDGS8KktdtKb2ckQ7AY/62wM
Foa5XGwy8OUIO6DSq+snk6i8KKsqFnd2GapgPFOB/P6Wh+jXyVJNVSACZZwXQbUy
DK9grNBQi8LEptz1qja9uuYoeWlYNbsUZ/EfWt+sgEflC+6VUUhdV3/RqFUEOKSt
A0CptgDrBDBpm0xSOX/MWFHngrijME9/06UJj5Dp/QQcx8CY55NK7q3XfJuVwF3u
3/SZd41ILy25ClfhVlVSX8FAngM02e/rhzTuAVvU5rQLrHk4vJdB8cBYj0n47kuA
emYAdAVyJBe6Ht2/253QTseXetDM+ez6SAVhAntz/gmn+tzqb8klY6UI+YQLuAi6
iWTgLF1G0peQkDj8WTnuv39ZFEtVxXihNzPdlx5P8lV6LN0T3CgvAHghMi36X2iT
bZYdclNfvuk6LSZkFhaOh/QFbGuFwmO3I5Qc/CPTN4YgfhUTvXeq5gQCvG0hunzH
rGYaYiHGm6MgsJMdAHSx+VTWlytYKkD38cqnlZblMKKnjmqx8t5gUuRMeVOFk3tP
o2osoOxhqqm4fOiekmPN9qr+QX1QcEofq5dJHzcsGxIBe/OFgPbCKheJqfehj+mE
`protect END_PROTECTED
