`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YEZugjmzLAaQj8H7F80uklF4TcQ9d7vLL9IXJCKG1GIVcFRQilIbMVKzCPs1mF/1
ge76fmp18O1ZlwI7hWjRKsFu2jZyOSeyYzynqU0Fr2XLyFDTZ7RBWn5XCvSHXjMJ
guWppBX8AACq5F9/vyZtalx5aVScOUMfLEd2GGBHaW/eujoOfSu5l5u/xIC4qkfn
uB7fM8Pcc/h95AfVptLbvmFsV/OciIURyhw+zQx//JsQGog44I+oVtT/UTxauVMm
WgQlxjJwRLnEE4AYo7VShod1DHcx5zBzD0NZKvqhFWJQuPtLwgK9v+CMZGcAmTQq
EKncC17uSfSjzO/sIluuqu2leAYhWG2AZSzjhcBDPbuEVUuaOP+58MwkWW2cjcAj
AnliDbwxbZ0YYSbPHqkZOROiIv0PMzh5RMOoFWm+cmi0dOdAEOoGWpJmFQdkuCh7
lQOBbDNtRP4BZlttBB+hoVVj9itUvZnrm9gv9Ujx0ySoXjRLFsN51U78Sop63UQR
ddAywXg3qZPE4F7V48E+Ok5FH5KjVxpAEJvrigc/UDPPsduPlxR4za2XEu8zUY/t
huUBXEUOpK5HRP1+srbrcsbIdt36k6/x8GCOZjzRRJ6QCEIgXXXhpOcKNb9OBeMS
BQ86TRgRlB49i7w2pM6uFzc8Y/R6X95OxdZSbvyo6GLNHhRqOPKoAe3PEi6/lhV4
/09EHGyOaxW6z/T6Hr+j8Lxnu/Ca0Hz9h8E7tfqR2OydJGjWy30QCe0B3egLd8jY
bJyX4FiMAO1yiV6e4x+5h+WmEVCtMf+rRXoxAjfLzkq7mChnp6E93jKeBv5cqG7V
UhMmOvXQ9VKw4oWBYIzjfuwbB6VA5FlmfXZorBRRMKYbWVQvLTgUykGTiTjE7BoB
v573KwxuL4GYiMojkh0n92dUDda/VWzXPXQFJWRRqWVPq3UF4Tzbt3oDlV3IASud
pgO5Iv1G9iIJmyJxlxuDC40d+0f0tMKGTwzgnWIFhzdIdHlUgAtWlShNsixgRCAy
YCOMuTJHgmDvJger+auVHM5vRkWIeiBW2+KQDy18CGKateeVw1TkU/ZxMcaMRkhy
9v3QRShaZlKLu7zedRErnCeEAqH06YQvjpgLy1ar407SNL60JdeGs+BdIciVsy76
2rKJ11oOXIY5T/AatP+jihrKGVRVChmLhWbXtyJZ2MdxnpPaTT2byga/BxN3cgmy
ygWZ7MidPo5zYAS8Xtt/F6trJX9j5528bTHaQGXtzWjHRqldydQidK20umGNJ8Ia
iGN7bfIafjhi3pAN6ryj8yn9gG9M6wI1ITraVzwaHncJjqoydAB1izfKu7ot1U2z
EhaxNLIb8e56yvslejZQUiybFfb0IaA+OsFQWnwdbSqFpBB5JQC/vuE5b9/5N87I
4XJzy52hjtrdWnfYC51Cnk2/bUQvzsNLxXpdNlxk/E1FBKh+mmxld9boML3S1F+k
A4mJjlhs2PrZ1I2+oAy5639d+5bnA0L5gLlR7tMy/uH2AdqDQa2OgkKsgk16c2dM
j0ZIX1GxqLMZ8xzixmmnHLzJjC1HE8iIwQ/5QPhh/Rn7HgaBWqt6IN3AcQsUFIkf
/ldjVtScFzg4EuFYNif6lNyUVgNJ6uROwSf0TtReLuDZ7Z6m78wvDxjITjS6BP5X
+73CT3RtKdUC2gw7AeHdT3hDFYVySD7SOlNNZ8fmhR2BfWiJSMUMUklc56PZOJCZ
3Sp+si5HySp88osoU3+qAVXNWl+YonDZiRJyeebxSjJ8lCT18k2yKopcqAT1aLBl
q9Csrhf/V4YByiPOjUuI66WXN8J928RmBrGG7oLPJl8MssI8y7HfsJQ0di59NHyU
0Y2s4sySWdSr7qYJvLaBhSVLoqXfmg8JU9fI7jhAXtUUnvQPHUcwwlksef9SeE7a
zHo5vlfx+KvOuGIo0ErausCKkdWpKZRoUf22ywU9lj1j0ouAy1z0rHF3w4h4ZNCj
YOLLKMmPUFwspZkfE+1XhV6+YWct0Q1nPqa2GDgzUk3+6IUDO1HWF3nnEstvK5hP
uSEc2u6iJFdufxZA1Loh0vttgdy5eeNU1RccDh0GLbXCI6mwS3VP/NyEZc2K8fZG
fqvCRmAopJA8qIVVGzJ6T+6Vif4E6hDss7UMa3nmDNx9/2EI/y3vxQ+qpsBU9EEl
Er2JLvhr5GVPBZ87USlNSRDFnemzJJIMI8lDZR24KoRD25D4NhMQi7SfJwlg2xzW
1BY7D57RykdHgTpZt/aV0El4yuDvjO9+dhcezDQGSj7sQJlt9dP9c42PQyLN8b1I
RIuXDT4CUWT/Pa6g8FNkvvJ/bGbqMjJa5vlj/MEihKJ3sIdrJ0308D0gqrXnPXF1
c9XzRpvUtB4uehUy6i498CTqP2hYseO0SyPCK4H8+tJNvE5k7TsIX7Dxa/Idz7xg
HecEsjtIAPpAq3OVrbhKoo+Kn0Mu3dgxGawheVLnudaII9yxL2KBYzqhIiu9Zuy4
FhTDcKaNIMelcsOS06YDnwmwdK5KQww0Q/rHDkgYLBVeCr+HMw0HSxd+q+MlygWy
lF0ABT70vF6GGoUMSWQaw00Tt9dt+vpWEcyr29VJD0avSMNu/mBtcTUw/wwFblSx
5wTct+imhFqKK8jL9TE0xVoMw7smuf+2sBzapIDihJWr/HOq6xrINDKL4CmrGjbo
Anf48AZkH635X7V11RimFVgoFyRvb0Z1tgsA9TlBQjiwwTok9WLd4/guz48QxqOD
cj/jUxUCGsutBKmglrC+oUNQxeA+mP9oB39TmRbz7JI2LVO8hYBnoq/jLxh3NKP1
cPsJ/De+jaoAXWhEgw3nFB709jRULNm4F50Q69wrvJfT+6ln83sUYxbl+v6AjoL7
ebBefxJWeDAAu+s5a2G+HJ2Cbic9JNCh5Y99/b1MXDkKZvmeBbwQHxIjTTP6OxaE
2GNrqjxgxfU/BYTct3O/6uB06i8wMlvy4PdvQ8SFy17xW6IcWMdBLbzulJ/56mM2
b6WMs3vlCUIBV1tbONEGIjTKje3XUGsdkYAYkzdHZJ9q8cUsVNa79skENymhPze4
umA++zVicmzUk4ESM/7tEAX9jo8Ht78lXUtCDxlst+7Ogt5orNVuRICyt5WUd+uM
aITMExT18hPI1GU2aGx9QJWjNhv6CLEvPfx7cgmANygzvQIzSUT5xo5agFTcjNNB
e0hD4f9sKcqgeXtObOcG0p+GwgdwkH3Uer5mG6EH/5sZJ0w7i3hMj0yLMGSNGFn3
2SGF2UkRc7QjFm5h4HRYH1uTpKftJSWrN9GaKuqRmFIKhpyk0xshu8mrCn/JkWuA
C+Zw5zGaT6e93gjpK7B637PUsnSSxvEhp2IW38RSIAm0gSDkGcskjDp9NUahLd4J
mAQmH6HPwkExeHqhLrNNpw64Ma7TRzSM5UduX+Kei64wHFyQbKZpONAWT7A4J6KA
gXF64iegzlfjuyINw9sD29CblemBhof7vwFJgVUtdcdLkMNCC9rm8OTbN/XIco5P
+Gj4AuHKXxJ0MXGCG2SvRZFxLV7ehFWKsrRkTMpx9wTrLryOnUb9lgMytG1bHfD6
yk46xhKchIK70UOvNp9MwZJxcUEwrRk5aSPHveksB+y/a5Dgb2wpmDVs3r9fPO9B
68TGsaFW83//cQdnhOdbKD8hPYGnQflPqGCyg9BJB6enoiAywC8KYCq1p/MTsGbv
Y7pQSLDGuBnflZ9nL0w7vfV+LIr0lxnI9WOaX6MTHGm3LZQhBtF/ypajM07a9Oe2
2R1KBwHjgU/J0ammHoz8vATa5YRRLoIvSOSSO7LuVXulBhfr6YgR+V1WwSpujnTQ
U3+npnR5xe9xs1km291XIwPsmxE9ukSTt1UiWszD5HpcIuaAUnRJXLaCSSxYm1Es
xfYZVo2kmy0AoUk0L7G7MoLhzyVxbvvPmcgK42Etabuft+IZAdsLAWPzFGRTa88T
YGTaHVzIrb2YfxG4L1Fe3pYo99gwc/ioeAyVDHRrOryxgcXdj+F3lR+HyiPQhwFb
42sN7Y25yRGFZ7/yMPQzi9TWlkbT2V9KXAZB9GaGDrYUCgyfzLgjSWAHpE5OjvM6
K57Rjtw8bKBmIilKPmPLt6gAwrB/cjRzvsheS55+ULt3zYQy9CpsgLDcNqJq1D0m
DJ9L76qxDe6mArRTANYb6P+/9OWOPAcNufQgbgRcVHIGXP6dpmxoK0l/YvLe4z8V
m2RN42aN1GBHlGN1JmFScdGpxD+FyvCvkpTkZA+Vd+dRaWnx+Y8gVmA5ULxYoXu5
x3Mm1vjYUTzotc8q+Ptlr+2eWh5WeCsBF+lIzkQxB1GMtYZSlGLxQcIZlnQn25El
gApgch+ZHFKx3Q9p/l8BkB1OnLy683crFI2UZ3cmJtsu3JUo+BEX6PdkpYtz0/gB
VXWn58mFtK4Zhy3/VuqVExkAiQ882vkNjO0gmfeUolpvemmXjoeVlVZEOIqBFglL
xyFE+msWZEz6rAnE5gZ35q8p7oKJoQzx2GTuCR53BIei7pGmFdFzddFODC/vCDDK
OLWQR5jmr0cEFv+HwtTUaSusqGebP7EzPR07LmMEVCSdVye9FCl8AKHTVnvSnL1X
wVK3Tk2TEHFwCo1bhvHENOxn+xNgHrw1UBO+Moj/0RhLI9C+luDWokz6yURfguUR
CbMYKMELDhvoSl74tWsCgptbFT9zivdBbrSqNAjhtF08eSiq8szeg2e9FoKwTYY/
2kWZlwcAq+QJdN7LAFopWLdSxqr9dVcp1Ut6sLcWin4QSw4E01bkFgWdlXZXKvDS
Po5cfUPKSfHe0lHnOqJ05fy9vl0jZ2vdFKXHcq//mRl38Z4DGWsmWuNoGLy65Csz
/RQLXWiZrL0lHtLQ0jdGU2BIvqO0dMKx8mGYvY8Giu83WY71CfCDk8IJQa8sXzxO
0+e32L8EhfXDENM9RACmJKyWTcMDhUnZdVrT5afS2EJToC6BAZHh6hHjpxk/sCZp
lYPx1YsLMwxb+kGV7v8CbYN2481KpNPRb6YDLsDM7L3gA1EIlbXfUAm+yxxtVhpN
OiQyIapbHmaS2ZIaQz8NsEQrZ49TypO9U8agDkMnRuvp+FviZoAWCT+CXhXCmEQU
Ff41+T0KpR2emS3RoyT8EMsLsUQVXZB01T3DiE68SBd14kodcQGRsd3AlIuMrA1Q
gxDwQbo2N6YVzEWhLjq+up8SdV58YaVR+/BiyMSrRNEjIAoGcC3M7uIQoZiALAH6
S8WHteK8Y0/rjKZWOOC7/4Dw7LCq7cMmsJ2Lp090SZrRZTf9cSh2MYmvtT4XVjIE
hXosC0A/vgfZfMsEjtDaKWrpdPia4t/7oAClcbH5FJeKtYxRe9xHLNTl/2EZPGzT
4d/dWPS9YLwFTPMiRWG7BJNkOKyasI3RzxlzUrS4JcC6lQzznzDBPLdg4ueVC7NB
nalQOazwHdn23EpEH0M8g9DQW/DHSLlfRwNDM/rUuVpm2LlzPKNwl12gUZCma6G3
0SOk/02MXM59xH2Ny0mcPi6zh22icMubSb58dXxGEZVDXpnHQOEkTngU/LkVF8IW
MpIbz7hul6YI+bFow6Q1kqcOgVJ122vagikS9Wj7H39w0CBk37NNv0FJ7p5udTKj
h6wY0+vxVoLa35MEbaQK2fpTfyJO33JZJ0T9jdiFxEOeDZv6X4lVFEI7K1std41e
askst9+6T3t0xrdEf5yDoyyPIXbUxTaCczfOWF8e+sp95owbtBX+h+xIPUOjN1LW
HAyAik/t6Pznpgo3sk3yZ23dDUwzaPK1U+HuLh0UooSMfDNRtVLj0M4AoLbI/hT+
ol+gEMLzFq/Eut/p2QpPgDz7SYhIYy14IUKbPk9r+or4jM0E3kE44Y8QhiX3CyOK
I/b54rysU/735wc4w9iuMGarD29PfFWPLtNvW1c6okr2nELlzjNSkWm5FlE3hYEm
WFJ/OiL4CjUkMy/NtT4oc6I9RzqV1gh299zxtOqjX6kJu6iOHVSPZJMDi/yGt/8d
lzx+wu+dC7b0GWZ+9fJ0wfkvv0PMuMFITag84/1M0CvTvPoh+QRb4hQtAQxqvYco
eJzTQC2f4mzcYDUkqN8gsbzad7S+BOnEKaVHuO2ho11Rm777YatxMEDHWxwYRZiw
byHDUboU2uwn/QkxCu/UjrFWuU9o0M/WqdoKTpoUq7aq4Hruv3llJyGFNGsWyJrD
QV6GqBk2K/eM1nwzcq0wu2EHWuR65FRG9+aIrA+W+C/Kr3KGXwm1sT4Yylbzoujb
p4aW/2kUup0iz2rontg5JeKnY+24xXAzjMZJGHfjdQ/eGBr6Yu6Ehf16pWolduPF
kDsQfnsSz+WXQqh1WDjrkaKBqLVR/Adz0A4Eid742hyI07WfzIdtGNCiXErcXyhO
F+ly4WTglvVmzf6VK4EFIp/WzHNNZxemYuODUI/Wd15NQuyKh5ScgGMjJ2Y/zKmF
E1doLPt2qMHo2iBgG0A/2+ffTJU75Nr3uHSswZreF1K+8+lj6823izev2sYdVdlm
NiuNLzzHc+o7dKVDi4XbfHDHzOrRtxqU21pLqafwNcQKIwypE7RPJlRUTKQgvF7J
Kj4urTpuLZd7dZNtmqyjMd18GLTwXt0v/XQLd3MM+pHIePi0ee0cEHZW4reIHeRd
M7dT0Nd4XRoOrZUAMmaQOcIx+siu5qRqIDQK6cmduPi+PaoP1PdF/jb6rxA7Lg7W
Cq0LqR4+V5ynH1kaSV7fYL2E1KjvjHj+VgZRAvve0egp3RJBhS2VS9v9hqsR5IGW
uINnHgQH/QNRKgv8F6+XE2oa68a1K8cxbhGDM4X1eEXCNrZ+VM6LbhETeNB1Ky2H
W8QhwxWF3HS1uW56OWW8s6e4mNiC5fe4A/KNdNVDZKlmBxT41iue/MZ1zCxiSMZl
Flfn3BnYMfkIkprzpCWGNCCRLBFZmsIHrutHKpt5gtZ/PxH3TbwWOuChKZJPH218
Aysq5evKKPtIGzZMJM6mo6epu2GOJJ2XXgvoffbLIXCkzuFvYQmx/l9uQpkDPzcy
Qac+7o7cUJ2u8+GxJ6qyqlKkTuO7XG5koZi3s4oja1ln0nJ2y+m5WqPnqU7fHpG2
zt67PmizynqSUs9A584cfcdvGCr+LsLKdYBRMAPAldJRw9REMJ1au5KYvxxTiUyB
+AOf5U1xUu+lnQg98k4of6wHMQ/W1GZbAtFC+xGzv0H1Si5uHu6dz0rfsoVpYE5F
kn0hJa+Ugg/2YUs3syO8/pX1J4J3nre1VFHHHHdZ0Hs3KTFHHXhXnZxRbW0EO94g
YvJrMkCZnAPsylSKXQDW8A==
`protect END_PROTECTED
