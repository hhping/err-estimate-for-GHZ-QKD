`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
px0NJHbVk7YATQk2TQxNmPYhjA2VZwEnqdvkQmiF+LXogeA4F+9x3P7DWWNBk5CM
xMGArUa5jkXJXOC709oG4iknh/YzzH2Tr9DV9Ln2VKp2Srfc1LFJyt8O1j0b5DTS
hGb4qkC3fC522g62Ykj03vfpJ5CGZrpjIaCY0+7oOV4Yu0gLuTmI/OmVhms+zt+w
O/H9wQukhFCyS6o6liFeofMoFxI4YAQa4DZMMn5bPaeelSQyN2XRMPWQyYdmIMoI
nqXgn7HForN8MwFXCT8frDftfB2prTfpp0LTeFDFayi8r+eUVAQDOU3RxxRVhA4A
PC5L/MC94iSGyIIA89sUupRii7oVmrmTv+9wZ9betZm7WBflS16O/jZSmCCzr9G1
c/7v08edHUJgLHJy7DGe89bOu3pUKMRFK1p3hu4MyWGgkYiZcwVoYUJQTJ8HHwIh
5ThIuiyS7eShr+rIGs/e6dfiejcczmxAMhrkUGbdvzGc4wv2YRftkbMY1bcgXHgW
lQgMpIK93XPX3jIqozdiZgqSmbozzcVCNQUqTTqsTcYMSyDRmeXpnQZB6oMQxSqm
L5gskw9dPCQMX97pDk8ZC7vNOuIvu79Ex/63tA1jia47FGFmmyxg6rscGAIdVO+q
93Sg0caL4ABe19/VsYVy5RU6pPl2rWAeDQUqVmiN16c=
`protect END_PROTECTED
