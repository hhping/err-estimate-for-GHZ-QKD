`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zz2zddTCxtd/h9eoA5A6Fxl/3xqGMMfHBLs29ppGP3jgn4Bax6/KGFJoMmKsPJN3
m+TTFL1lE6DH7kxpPDuc0o4pNQUwiqHHAeoyLUFzF4OxKAXi9EXjx3Sb4uFieyUA
JqGMZYId01lXlQrC6mc1qgdih8d1uIxPxjyyNSMRVb7yCKmt4SvoZ3F2mM9h/EHK
RHS7dv1pjQHfClbUxObKI0RnjDuuKZv8bGDKaALQWU/iZLp7JvzrTD+bF36gYzc3
6yy/iL5RSqRcoJg5xIXuHZm6t8rfB51dQU55FfAdoZPuGY0VZ1j+HLxxD0ux4Soz
y5EcmV4gtSkD6l5Aa87ebfT+Dg1MtyAA58wHLnvkXfc44UUxME+EuDfj/BAi4a57
yf+mH6fOQA226sZ47xWLkHvds4y3YC0G3pSAUWs0cAev36A2Bpjh3S6ZItn/eJz2
Af8nQUkiWJaqxJfvwdzai3Iru99r67XwOkQOzWAThfyH71ASDbFT5v493oqtgW3E
SAK+uYvuozU0dYFiu2eH6YtzvvAwQEzQXG0l73LiwJq0OQP4DHrZjGfmH/Bfr3XB
huvip6AtfTIU/RKiOYDH4GhK21U1zne25lAg+/eJfHJ0YJqFMD03DI5Mv09tDPce
YzYemtOD47ktiFIVAiykU3timQOlpstFK5zNfj2b9PN+uwMkJOBPWEJzBG6UsCHI
O5mKwdaFJi4c93rG0m0hIrTeHglptrrHxH3eOGeZkh5WUTAaVeVwvhu6oRsmDHtx
0Fy5hvvO4/VSRIkvKFCiMzOl0WWaeJopZW+bV/pCuNr0GV0GdH6TkqkB7zRLwsmn
lBr1IaGNx10TA9gZ87uWq6fn+T68gbOpEAafRKJH+teiAM1x7d4LATsPH23B9LbL
KwMhdam0UK9VCsWKcYLroznJkzn5MkqotF9z94gCw7sSvvFCZcij+Y8kREN5hyd0
54sOy8zjMflTDuRCqCoZG3SaJMxGJzuD0wz5phh6ssNCAW1FD5azc8mLfG+N4ZLR
MEoBvpbyhtzLzTamcQqxI/kCRCseZiNB1r5iDhh1ZStmfFFN3xZMmRrEzONzLMv6
eWXqCf2WWqpbQhLEKu7qR/goykoCFjvsP9GtN1UNH46ZY+kaJRMSqJHcMfCf77HF
163cfTaO2XbmN+9bWHgWmWTr1P1xWA0S7yFcQgLe+KJvdNZYKVYh7AFWM9z4SX+h
ZaPLq+nojCOCFIGOgjrTplzDRRn4xjfe/nkmIObzpNESs2jHa98CZJ7o0TFwQq46
MWtWjNTHrzC9mfqmWZ48OC3DiWVhBe/YTRBPUFurkApfF14JxnF5d8+QY1Qthq0s
w8dqtHjqZfWRZwJ7X+zYvbBNWFxe+pJudCJq85Akju55FefUNVH2vDczHSNFMl4/
JUi7JyOKMLBdoCaIjQ9NNql4zn72DGsoz6LYI8pmJrpT4HA/p2LchFpKaaU3oSir
KCoOUziH4IQPU6f3cdEfWpW/E7sqLQiAs3Qovl5zSRYYNDtKqUe0s2V6IQUeL46S
yboriA15AdoA3cu/L3oe5tcSFwvK/JD3j7jOVFMEX4u+PuzPR0O77hWas3t+nx88
UFzudo/XAOae/9SrgE9ZelXO4KxUhlFjIqvPCaV+mGVbH7tr+C2qb0jpz61McOBv
m/kxxY3JM/KOV0hKbN0g5n8nj5uwDdNuFZnqNGn+EaKO7thTuVeVCUvZSTJ5gBEI
96BXar5A03apwibT9gi3A6VVSkEOdi7GxcY1BCSFEUYNapaKOdg83P6xQ7z4HMoI
pm2+FFQNVVJdA1CbgEEkVLxBktX6dPeWoUi9we8TykEaIBqmCY2WMOaxaOoA6DQb
Brz2VE/dG0o0i0282Sw4nw==
`protect END_PROTECTED
