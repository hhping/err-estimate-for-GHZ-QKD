`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9neHCEKXKt01vEXvzun4/SoX5KHnm7hPgVOaDFoeeWLMKUymim7/hPPABU5kEdPl
IIFLJd4TCcM0Ao2X0pmm3zHq9d3RGwxM0mbx1ZVq0cIYn7hxhZfB86TqYkt/WoAh
95K1VoM2HjhuzLmKLo1fJ3AI+E3d4PkZb72WW2E2tOYLSU/PJ6WBXZJj1SL5B53s
7VfWD6b8vjFVG60Um+Eu4LfEr90Z1ozB5CyCmwYvpfy4YfsgKJ4wuYhM+lohfxpT
uSTgd7U+lNzyqG+Lq/5+PRWYIjSwB2Yr2Ag7pkT9d3FGYh3vCijW8x64bo22GTeJ
ELjnPhqXDX/JNTcbxYSkFtWNCiydCuRjgL/Fe9xn8S0FIlwhzXCttWqXnp7bq1zY
FdK2ekeOgAkvK65g2iKZGnagR+xzzfDgeenJ8f90hrqOXSDwKTCaFq/yVQ7Wm3h4
lWSKexseKTx17ROzGsNXmsuq5O7Ikvc811xI0Sg9M5BxJTDlFbP+PzTfv+mGSwV2
1sqqRHM84guA3KtexnEH34ypqp+PAll7mb3kqd2HiOKkSr0yEbCiJVmJoWZDoWHX
qvwXnzKi1AIXjwcukHSAWi/yEiRiPws0vvCYWc1cbY8jVYGoPdqn3uakMCEDN/u/
tWEdWFdbMNTOlnIY6pJ5jsubnyfOesBYW3GAdaveunCHtTVJwISRJ4EO33c56MaP
CxbV17ol0hv/PhPO8AYYY7B/nAbwM6okQ8gh8oByOm2bq4VIEuACcWrLz4puJH0E
jYDYNFKUuwv4wFdVTTlNhToIKu8ke2g4p4CsYeAlQ3Klre6l5wsDm5MWWTTE9nIo
EwE0oR/gP6ww44TXSPZDJQAig6+hpM90FyiP4P4ff8JZTW0+/Qhch79KsIafh4/N
/CBHPlxEvVQrOr0slZcXbeSf9aMfVPr3DVFA6RPEijnoqAuiTJy7SN1wN/E4ioAc
tVX3+gYAEw2heRB6Kj8puweGORYKGHic540mzfl10VnPwTyWENCXrhvgql6iv7T2
ZJqyTY+3BRheG5VgCRJd6SRhEah2vb7bsdwOxmJ0xPmFZyYeWK/iI/O2igSaWRQf
m5rkbaquZm8ATDPrAXzTGd/7m2gwlrolTkzFeYGzUhWX9gAHoTMnZa6Ez2ZRsGIq
jX05DM0k5Rezf0WaLK8QAMYDRQjjWKT5RPiE2coIDCbliGrQJtYXz83AECtCaIDI
OQyyFw7/4x6jRxuvuX55dcXZL9ivkRlg2J4ZnDhpm9qmVRzxuoU+Ml7pUx7LQqqS
O59M5oSyPEt8SGlk7GKg7SfU0Q3SjGEN7OKeNik/A4smNscrFa7MAgH9428YZMk1
p6gASE9vyXcshjyC7boIqIUbruluqDr6sH9DQ2D4mZnMNI7wHEeCXyavKW6nMsyS
`protect END_PROTECTED
