`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hQ3ZUPbei8huA3I/MTVhgwwoSbdOquu59YyaeXU7QFs+vPtfpjpmQ5fQ5u32x+Q
8jWLFgMjdUsnq5pBrBIYo4YiWH8hPeAKHEWcqOiAU95BeD8tUf7RSo7ztn/t9Jvd
TksnIYisXflcRrfjUai2On7XB5qMs68RIiVN457BzjeXZjMY3AFTzm199gmenNd3
0P1lgQ49PKXE6SHOQfBR7iAbBQAjOxBIbXEpdGBT29RrCpP89KYn1zJ47ZNowl21
CqE1pQtlqTPkwpJ/BbdgkYGNufUe0U8PjlOhUx+xduMTA5YcjhgSbTm55Wftem6i
qgT2C+1WJ3+jb6tLGRszphvjdMcidprqRT1oUU1l/vCeJG6hykM4T9pA3QAmlpbK
D1oG8gtu87/tzKa/e2htKSh6kC9sSilXlbKuAd6nAJA/nmLQs3fFlFoImBplcDFJ
GsF39gYt+pVNnZTc/7EgAAmkrbPYNOKcvPY+KdXeHs+3ullYv7cUjnqCLHf0tk+v
69ZKgkUKSG256ve+bIh3XiavN6zMcfub1XOzy9D/k5SYqhsMRkOXHKr5PW3zCPcL
qIZRN6wam7Cap96VDOBVDYlKdMXpIrafjH3RxpUkpGAjEVerOZ/1J+nrtafomcEK
O6+mKclVFv0J9R63+sWp49MJQzzZxvWi/PDP7qhddnTPPDY0rHvRrsGvEn8INjyB
8oMiA/ICgMIxBktNkgl+Vw54DhgMrfRimUYQmNAsjr0tFYkDyq40N0OguVe7TdKg
ACoNz09w28zV/z3FSIfNNNOCmTLzGbymuHn1XoQuhDE=
`protect END_PROTECTED
