`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAqBG+Ys2GJkqpq2ea64obzQnCovqyaKOquyhr4TerejaAcfBrMCFIBovkIR8jt4
TE7RCwPTZ1mVtdgcWvzXot9FShStp4NoBcRpADh2F9mQcwEJY5H3d/W9yIa3TKWG
CeIAvbunlb9eMszdsBXWSiXtoNJYkfymArvG80xFTJ3qcWlzyOdi9G5zhES9dEvA
87OHnnMbKbxh7TmHAcrGPyx6nB2K/wT2r9b0AvuZCzsUWS/hNMJdt320mjMOHRsK
hYlENNLEM8jPM7Gbg1cKgwQS79jAEalRDqR9Cy/ZpIED12a0ScRJwMoaYxCWz3SR
M0irxSaW52f/aeE60mAjgyc4GLqiVPZX+neC4Ln1PDkxOq8aC9Tjp//oTQI/cWEW
reKbT6anTsYO3eIUV7yrksojKixi5wqzOdBxpSutsOOr8R3pKgzNNy8VQkTMkJmb
u15vVGspMxT5i01d9d031ieh7YIB749fMkr8/fFaka04Y89m8iXrhv+QoKRp/6Oc
Fb0Ov13wh7vo1mU8Pm75fg==
`protect END_PROTECTED
