`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQlKI1qcFi4j7Ieh3XWdBlCTSQcjGn8JzJa8dVrrGJE5YWWeMXpWpAT7d2GZBdun
qNdpV7ijCVreSTPiBY3hPBMdB9wIAdfjSUiQ2YP0UH4gyEdjXfDbJZ8swHrXhZ/J
Dhl4+kgTu15RBPfDjZsRe89P23dkPOW9rGX23tANADZcoPdBhg15cp0EQlM1ZfBh
GwK18USuqH0DcN/6er3pQw5xoAIQBLgvy2it7ci2CiywM9u563ALtewOV1EN/+tg
dlnH1/IG6kISNYRGZ8z6QlPtmj98bttgGi02cyhEDVe1LoWN1iN8MdnNU6pQcbNh
o4saVbFSMjp+RAJVY2ygjP/NqI4pCjibt/W7IkI+n6E3HkyqZzHiC/opmrUm+795
gz8qjRcsVlHih9Ed6fomiQ4wcSVkfr0ui3TE7XAjgfuDJWXddHBwy6QqzXU8C/be
QyST+J6A3K+3wW5aQoMACeH4+XB+C9NMxlvkYbqd5A3xplvUf07FbQ0B5o4wMSJf
46k0hIqZeL8c1GDmnCXHfBmnTLKG95sjLjOW3RRLoMJDX8ALbBhdrewRG9D1DdjY
InTU1Yq8gTnV/AfSTlpj2MVjRF0pMZHNXIe7j+ySx4xy2E4MIQn3zHeiwA+cro5D
IJ/D7pcZ/Z3CroU3EBQjsQfzyJVZgNkhz5bHNpQUbJQDSUpsstS5L692A4nY/Rf1
RkKqDn5INRseoXjUX7/WIdAKp7+jcRv34D6lMsGsmaky5zC6CRdNhiP7jvogEJKr
`protect END_PROTECTED
