`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KPg3ViUV8Q/yhZFPLE/07MlPBHlCqoi9XC0q7UXWJo3OiSuQkuGn+Q0Zrn17muOT
UwHSDmnQWfGePKohoXpjuhKg5UCFYvpliL0YVvtHv1X0gN32/WoQxJJKSg5a6ugP
c1wwUVlh/0cY6nUpd73rDmBjgovtjt5PAVgOgLRxol8FgO27CGDPBJw4EEw8O7ci
apj12DupCV4zaY2oSoUDH4lp2kec1T8lZl82aJrPHL6Ut9rlyDfAiMk3bkH0tH92
JdyJsVP8WmIS0Jl3209radDPXl8ABu6g7RzdqN1IFHxs9WXnU2Mklwikv7u+Vubo
tPGP4kUjwlNFVrNVjeHuWetAWhpMcEjMlCQ/oiPnlzSIpJdjOM1TUpOYfKnHWSRt
FEWyjM1bkgiXR+Pd83rooVQhXAmDqUOGcm6LZAwnFdQ=
`protect END_PROTECTED
