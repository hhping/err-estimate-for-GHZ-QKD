`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gHc/Joy6bJXs9jah1EDKPPvWXW4eMSy08h9yIC/K+oCyyltTklHafRerGJJbtCw5
4ZMsT4KuyxkfMW1Wxy1rlKZQ5CDIK1uuyDH+NtAPBIhMkdBRbdIPAaxJp1ddU7j/
2wXuUbMowi7crXVsgDiHKfbXOeYi7VffXUo8XDWDkL1WldepO0+UnvhJ80rmrs4S
m/oHwTTnijFfn1Yl/rLIxKJLCMvr8RdE5dZeEHVvs5iN3fZXiKjRi9dJU0MZ63nE
LnmcR+ZbQDqtbfkkaTw4bAGv2PVSVXLsrmUZ++Et1U5mEIQMPYFBd6N9HXZy7YrX
LNRH/3iUzu9cfASzqKc/VCS+6MZvh/dvN2OUTBCoHgj7AeQsdFIh3kTD3v4gOdMA
yStouTSYaXOYRYs/h07hcyG4eRDJDeBNXE3awTIALpzk0KedhMA5ssJY7ogSfgjE
`protect END_PROTECTED
