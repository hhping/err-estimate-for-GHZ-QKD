`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5Q1Je3NTe30tnixmnk3Y16RAr3ll9N3zL4EFYL+ErAU0C4Xe08qaZFwFOjtvtDe
WGvayva2K/MwVlru8+CK2jD9ytOw4ul9crgdBLczH8lmgLoSWe4CfMRgJDFJ2x7G
kK5WBgXLBqY03a4jdrnH5LDV5jADR7JINIQJjk3+5NpY6XMQULPHHvGygTTszHLo
2GlatZSbsdSaYgxkXXG64x594F5AT12EdvzMiOT7w0RaO5DONeCKkvLy19959znx
CEfMjTm3hKIt4ZUMbmpnSPg2DaDSDrgqtLEOzp5wf9MPtmEnv/ftcdQPmN2if/Io
9s/Q1QL67j725SmXu7LkLvnrMRCPkwMIkh2gfPZ/MWgGUFRnhTF5bNrhdPzue9HS
nBptaHi1xOJyEBze/fGnJESQgV1YaSOCvrNsg2mjp5m6SJqyFxtAURiPNuH8TKKM
gjoDDP4fyvPjcCZJaAW1BNaKq5GqQnQquLrsAuVsA54qo7ev3CEe8zc6cXNZRxZC
l3bejGL6IteIi7VU66OiFsNLZw3dQDRa520Ck3fPqFvzQhciirvvrtFK75/OuQdJ
SHQkpxHKatMz18Yg/lgkLdFmmuqq7mbnWi7MgFcpJxJ/nMCkIMVE16emjSkwhntR
rmhHBlx+v+b5m/+OTidLlP6u1sSK4OesOP5hhNOFaX6ASkscibxYG8tvT6L25gky
7dIP7ZKNrczvoNcnYdS6yxpDcUlIO3q2mFt4Rj1SY6nzm1CDXT0PjqYhRisfwFOa
F/2/2Hw8CbIzSq8aC2PUsYxvgREbNdhOH0nrLeAznCbeJfEHOqidWSNMozA1ivZJ
88tnCixukvFD9LmgqABZulcoWVStK/v0IXxdQz9vPKCF1m0mFuno0MwWMemBFt0b
p8TUJ8P5db1oAun8fBUDcT7DCZHXuLBdCNYV/eFpIUbXrx8MPTDoZx68lKtz4shk
7bNLTFS5K/LmuLgVB0g2Ibp36NBQp+5O98n7TX6pV/3VsmeMiGmv0WGsSBh6DmDX
UwXk1EHYv237zXG3duxE4tapwmvHUN5t0iCescRarrzfeCOViIwaDiwdOR6HMB0R
mevIxOB2938NkATWJ3xbpuRndtcJul9AoryTs74jMSLEYhA0BEGpleBgIHPi5TAG
z99ljDX5n++HqBQSfgYmVskNUvLjTW7k+bQezwv5yUu6VwwxbE5ZC8u3cSrSvLIG
aU10VStD1dWcmTId4TUcS1isBLUIm9wemn6QMFj6SrH7Of0ZGR/jLcJTkt94Jkzc
habJOgeU07Ttkm9oopK5zOE/40xvcF61cUoBILUuFfV1GKIZw0ZzSCkNMU/aBrLt
d7UO0VtoTTaaWuHPC5XPKRVOjhdRIrIhrQG2kvFhXBveLIqSRKlsm3qvmWpJhrZF
DpVG25B45rlfFEPCT+dwDbMooH33C6fifB2yf12uVzffWiqTJlW6wUiYO2FbqJEM
nU6sXDJaHlhzbcX/g6XrOnD4mD9fZBFdAuLRnAq6wocATKhBbpXlXs06LVlSMDpm
RTG6iE5OBikd9pm9me5AtzTfhGRYZp7W0NrVqEM0sE3OFT2537jC6UyqLBgk6sjP
PtUNdPcW5FzqsAgCfK0vsf9NzGI5HO0e/y3KKE0EOwH0bOqa7IR2aJZisEeA23Cz
3ahEFe3Jx2R9eSy28skHlmaHyUXYbvdcp2uj1qC6rvuxFgtP5ZOjO7BSHaL7lS4x
l6oeproH4jlr3PYbnYO0KqjiYs2Y3qJeqPXR09NA2cHVWJI2FvUVBTURK5afwes2
+BN539T7iqV9dub8C81TFD3Y2Wz+OXnT6wfuBqCrFgvKY144DhNK02mgP7y9Vw4M
R4l1MnPZp212HUPHcMB50YjonDU3xW8eNO5v7dF/SVuu5JKwmvMVUPyIP3OmTook
jkoJBOgl/d+BWlySERfXA6kWBVdctcWX8A1sTFYhgQ9fWAIi45OYnzqou+zUY+XQ
WyYjoNsBbFY4iDLl3aHzfmnu7QaW/a5KLV0QyhcGV1VqCezBmPoSsCz1JxwMuP3Y
bOkR5aHH5AJ0NtcTglU3BI9xUJDsZB2g15D1tsE2xbZd/XkLJl19W3gXeHh7taBH
slFWmXGZ+gXlmIO1zF3C9o34W1TDAWnCTGnkIV7FwykDi4m+Va1f/gDyENmht2ev
AbbFXgQirY3pO44fQ83CPqeo8MSrOzyu6zDJgw4+rqS27S4DPQDxyUvhbfFvr525
1IaGRwHpzcFyn1DPgdESe5Kgxx1e8lPivSiWksJ9zuuLY7lOTGbSj/W4/RAcbg4k
VdlKRODh4kohuZ2FWyNDeKJr6j4LV5nqR5Yuaf19eKYncSPSc8YB2C2A7MU2tiGn
oQHfKRPUzB2FU/Re5+OKUgWWfnwEdFShfixCdfgLoxKUE4sN4W8iYZwGIsKmKZ6A
X6ju5O26TIQNDnPU1RcXDbpGAjxbBk5mf1ZSWEfJ9Is32XhvOUrbbSzG7NWwll9c
LOGkCVIswUWlUZVKyz6ONPr5is3yrhWGamoDhfaHTyMgTEHpQQU/xnkgMEjkw3F/
zbBxDMipUUgDC4Gw+BSsNTmGb8drWALvjpHMfZD8MDxTCEuQnNT3UXmNIuGcvH7T
qQBBL/9LD/0RJDlkUzbFUQN1KuK+Z9m67KAt0x/5mb5MrzXdButSgZBBvCnHBS0p
qB3MNMi/iEvIrE163NOkmJKBcsQD88JhaPZqGuxlHIaJewpxPyUgOaEAa0dsAqTb
+L2v47kXkvOCGnvqN9MGvTh5AxjMUP4SdC37nWlI3o6nw+JxIrUZn/WiIQBsoCbl
ofzN9rdQnb/22xt4W7xr2eznkP3KLYCG6qkJ0jl1XSshVx3jyHEmYXpH6pkyM9u1
JsMJFCjSkHMGvuY70RSbbY0tlWuPVQRqP9qtPK4sHmomBaZvTTMiNLgTEzua0cWe
Eb01pHsA5+V72KYxysAdTQDFtbfE6VmcPu7ALXpLCCs05r8QOjDITU+sM+eLylSz
TxxwQgLra6+1ec6QUbyv2ks/iI44p9rpORUFSbqnCWIKhBQYSrPDrmUkgUxaVC1s
Po8l18MnLsKynT1/hJo1mygIOzUmnBqOGmZgNDT81wLFeGyZ5gWCqf1VrCFeUerr
uA1tCZ5edQ9AunU8T7uyXw==
`protect END_PROTECTED
