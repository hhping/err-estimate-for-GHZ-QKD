`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLCsgy38B7iErXzXRuFQ6BvayLTkltVO09xkAyGJNB0g5jdT51+nFo7chXpzYzz8
ezcmGMPLzs4evXZ5dOxqIMxTf6sD78aKwaZ6xXOykkO7BGEeqCtm3yg+WMHoxnT4
mLYW5QvbHuT06no+fnTz8W/dw71X7vQhdvrqTL3nPdvIfCGpqPOaEXeXeRC6aSaX
90tQb3JONNfW0BEyy5/q42U3NPPG4mmL0j2885/tuD7eg5KWBGgiIxcxJriRfu4y
XFpo6QmlJqIqGy2jYOMqKWZqMQdmvvand2T1qnAq5Fq6QLCi4bPpqipwWxxT7Hw7
c0J86lCu7nr4t9OaLV/9i9hlZFyv8RoPN8UdEG9YB0NM/gRm58hOaULzVn1V/aHD
//QPqdHhAgGbHADNTNVe5yFF6ui0uA2HMIJG/PF65GwNuRket+gpILCDBWjay/CG
F7Qw9wvNW4R8sWHmTO5/uMwfuC0qAq+0lafpB8xmEdE=
`protect END_PROTECTED
