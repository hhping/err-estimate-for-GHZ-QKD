`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3DmOR3pNcI5Fk5sVY+WDj0pFBHsEe3tuvj7VnAwilrLyaKdysq87uFEPjQv2P7N
wK0Kx5WRNKJIZvKimkMRNtgv93e9DUOr0tgfzOxQcs4irV2676/DNcK2CWysOd1r
q5z3mXLsN2EdD7F9L+4TVsa9GsTlZyMHUgJXeOgwhe1KIQeCt8Bt/4BBAQ2HxIYV
734NWVvIGZFM7+VXmfOZMlBBOxQRs7w2/3tnyDO49ODLHOark9TW8qh52irDrmvY
wac+cKFriwOiUEoHeMtKUdmZm0W9sC6xlC4qEo2mZlJ0fJbFp8jIDK/IGxxi8YrD
xEN1oaI+yaq1g6Qkvwps6S/Ujf+y2Iz4sxK/vfHdsFMHIJb1d7vdxVvxTNDq0Tey
3cobgz+iwqlIO+3ipfWVIok4rL/394r5AqWQyeq+qiGpu+ZrYwgixYwEfHFpav0X
BCqIRgcbwdD8Qdndym8ye7KLj9K8KHJ5ZKwxkXJ2vU2SU/a95IIpFXqPkNttwUtX
qFaM6JaCtsNuKMnP26Xbim7HDLjT7VKUBpCn4xehNe/DyY4kAf/8natxfrP7c8JS
8xMTbBvD79EBCWhZMoH3XnnkE9/1NHnmA6flrKgCnpB9cmhxDBTyj669fFbJn4kB
dQZyQmipetO7s7nmUKItXKKcedeAJKzmlVd8v8CR2cEk9nyGIwwG1hnzCsNgVYzN
XVNy6fIPeYL1Z8d0+xbP7ck0zNn9UBnKvWYCKQ75n6mstCf7E2MhM7EtrPYyQRLA
mjDNuimaPJh8pie69cA3p6E2Fi1LN6w1KGPQsEWvuqY+UyVJaj49oSjF2tH0Ocmv
wWnwvLyFK42AvTlEhXRIzI7oIo4Xspzff8CKOhIO9NaOpjeLveluAXZ40hTYQyGW
TwuFLEvRivFZlqiNKBFX9K9SGCJ3uiaHa/Ur9YIjWuw=
`protect END_PROTECTED
