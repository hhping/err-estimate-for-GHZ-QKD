`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWB2ovLjCf8ehUMDSojgwYv07jIpo3iu5ocTT9m9pJTOkP9m1Yi5aXDaDDHuCl+f
mDP8KFHf69GisFgXp7NOjjSeozrS1FQrVkOV/G+PDFF66kTd10x1WQrX2b7aCc8D
f9Kut6olcYofa6Yo/KwT5CT/H4c+598WAM7Qbikrr+juanU6gZULndY2owFpZWJ0
cREvwviVaoidZ909aUbN29S6LOTDOpMxZ0oa6fxwiCt4vCmGGPqnvKFkQZ2EDM19
kBSaLefjzmgtNC7/7SknV8NgifUC226aKu0atthG9cMDtJYHnfh8C8AFlrJiHSxZ
UMfRnzVWayrLcJ3EsaW+NPC/rqUtzOLGTRF+bImd254GbxyBuMGsE+HjUghAKx4G
mFCTAprrzk4WVlnD7101qlFiq5mVf4jCCc3pHV+eCSoondTOdEXEpLqm3QaRoHrq
IGBYNfVNSOyJJTNA5i998WjflvoS7482/D0KYPUf6tgwnSD80OX+hJmOOnSQGnq3
FHsa0Wyo9MZCyTnneCxla3RR1KC/wFnZ7TJRbxD6PYa4eFfnspzFlINws7852imo
AClm6zffpT7OstQtOEXpG/SSckOr5rffGM4NkFu8v+uZ0+Zadmm03W6BQa/2OnMm
3BwBH5T4gQI5Cr6eTMAHPkI57Q2VNLxuQXucwCpy8FotdPT34ejJ8QSY74acmOW5
adbqyzlISGcKRHWIPg2t7GJl+5KghYOHkt2a3L+zyHDi43FxtOl9W81LEbw1J7Ov
qvBYRAY7EN78OIDoBVEvaIIjcK3ps/PZGAIu7lv43B9yXHlvJDYUf70dooASsOWB
1hKiWREi4e44eg+2AHDjoehsmhgrdFk4JPNt6M1lIW2DjJa7/5zcNe+tvW8gaob2
+i6J8QIw6O8A4hs+yvwRR2oi8H6+Mjo9FVvtvcMsSEOcfuaNaN3/giGiMgf/hSfQ
ukYuS6KrNy1J3zmVHnGylgXjZJswyBN9+dW4prBmsfV0+HGoRamjqbR0TfBZyFjY
ayqwKy/pnhYIFQqUCFnq9E7LSyO2onf89rDv5Zph5+hJVFWNHZLf9ZkakIfV4mKM
WYr+UFra8qbzzSXEL1Qp7AEKr960UeP1XttoowZMVtuRYBkllFPDOXFdTl7yvP3b
zwE59MMA9Ec9geEct3WOEey4PIpKhIINqJhX5w+mpkrqtxDb/VULJ39S/4oXWQXN
pd/WeZ18w5RGd2z7s2Hw7QXj0N1l6w+4OWGTwOV4OEelPG9sXmaTOO07ix9GOa/n
iLLivPCFXvU01GAHSiso42YuKiawqYlX08tYxkuW0G2cVgbCKRcWIVGzYOM5tyXV
qc7sQEVTgdmxOVKgWJ18TTOuAwUQoCUYoAIOT8HzHsswBhlFIxcKxqzm1WiiviSi
ty/FXrPHe1daTFaK4t6JVM06JHzEbvNpidHT0yoSjKQybsK41JLq0rzlLwdyPoDG
cpTJrDnhtve7y2gfo5pp5viSd311zNd3f80RQvY4cP7QPjAKftMlMl/WlwEuS2z3
rdcT5QdEqMYpudS0wDyS7YzA8SDFQszfq7j2C9YE2SCuuX04xODd2wwJ4+Zp+OZw
P/pxuxNR/wATha0f0gEZge4WU/CvurklnXSehXu2CJfkjsdqpnPCISLGGypp3F/S
vHGq9WzJQRr4GNjMrCIB+mD8WXBlja0tjnuUo7El7Jw2QOnnO0qFnmQifPB/SkB6
oR8248WfQG7PCHTYot3ZviOxUYElIiRgz3JCAxyvZs8QIFNWmo3A0PhFORfeH3S4
OE4Y59wOh6URLW4gFyYdLcx19CUx6tg/+84zFegy4rD1qMCSmLZbq1mmSmnvz/2Q
kKlD3kLPjlVGTWEcbSStyEunRfhr5hhKTg44zzPRdcfsIVQ6k4oqQ6wHHSmfPqHv
PBPsQrc+fDm/5RDWX+AcgE988vb9l9Ov6h0sirWoSJEBVgViL+sN8L3KRY5L22/b
zpSfwYRwHXPIsctr5bMaOZQ5qYQrPJLQf3EjkjumHnfdHMPARaSaykM9+0TvFTD7
DiH3FjrOuz8Y+Vpvd8PLpBzYdRf7bNknBL/zHZ7l0qyM+zWZy3rnJlOJIvOb6T0J
zgE5XekaKbp2VAk5KqN3BJAH9N/mNEwtrBq9+GN+ub/Ut6mhc+ssoedBUpS4xSgX
bqivsiN+Z8UJJEEfZC+BNTqPPII0f67PYfWj0q/Mhs3jn+WCAz4MZ1uPwZl4J1h8
Q77q2ka/cugn30i+AEljN08Wd8HklWn0rVMgG0am2jHIT6FNIm24c0enX+KyWdba
yDaMDdkSE3Vmfi6103Rh0xsFfbrIPnO+tuw0W3RgcGV81/yDl23hJjE10wnbY0fF
/+rwyqfNarK5x6wzFbYgPi7Jddj+d6N8cvKl/hayZU/XOtoh27zIITslgXCAKqdu
z2U0JIJ6EjkCcd2iK3OOYIIoHdB/FOiFmTtlifTFbRfZS8Kzmj+HxmuHNDmuoVXc
9GG4k4XFYJ1nZib66sIvbqSLp3A3w43H/B3xt9Oq9rPfg+fTlMWvFIsHFxdTKt76
jDI7f7YV18RFn47QdLfVdKFMs4H87C/ImhXH3W2gXTZ9P1uUCRpJ3LinFbe4nsIL
ftCL4xXxd6NtkmptaR/+EPY0EFGwMZ1qnQLURQl8W3u/zX2id/sZJ+DSd5P2wszM
IbuV2L5uzzoLlr47jJ0GeoWcRWyVjfWQbRW68JOSFu6c1cb0cXaL56t0UWDs6Wfk
Wrne8Lr/86pYbF1Ky9kiRZdwiwhjHO7x6b1atjB5fCpqd6Xq5MqNY3NZi4vGov5l
wYfB5VX9k1AeNt7qKXIXIfPSTsGWvLC3EhzQDexFSZCv2CCEE3L+C3CoRUDdLeo8
g6QBmLdWLKmblUwjbG0TwkqrHsPBk1ihLxEiV2Btl27tGtCXVrhrFro7+gEjetWO
vlWvP8PXBEA8DRx9CtUxTUmJS27KtxBPC1vFG9ZeAPGIvPh7jzc/JjY0OOIWiiK4
R1pFuSGqwK3XOXNxvVkq4HoODZQRpe5J+aeyFoAettzkKTkV8mcrNuTcRGm9uJvP
v+CPlgzUtbRv0mIf80FICAN0wSm0h5qNTT40VKQd2qwmCODZgeYXLtHd88bvFTl5
IqTWW6IRuwOb2k1qemhNIpbdI06owJdHj/oBCJYirDIRs/Ddei3gbZpvqP4bjU/E
BajGQUYddBH6TN2UyspjRmMUNeoPe/qDAOlOAmzauAQqY77qjTWKf63dy0Xk7MA9
deIEf//DmvsvfVhoMwbBbWf3Sk5bwlVj5oP2rEFbCKyeVTSeDuF6OS3kK565W2Bs
pm4nIERNC73FXrrG7GXY0M+VZ7AddJzZvhDBQeE5Ry54icL8K2rleZVg2ouwBniU
/+M3vniNJw1ZTkp51yuuaHwIJLQ8UUDOKoNE66oYL5GEWR59s5cLmvte9rsD2ZRJ
qutwMlUbaaen3+sgByVfkcUj4y0OJSKZWP2BX0WRUNwsvuVhvQEs2c/kxYZj4uVk
DQyVhzMs6fUmN+k7qS4ysBp96Bl7m0oi76pcv+5Khq6XbDcliok7XllmS+U53YYv
OLp0WL0xH85At/WMTyRIo+MIIcA5wnaa26DMpV/Jyc8pQdcqW+1pQMZkMj2PUaxR
T/LumjKHbRMoXaYHgia3Rbreq+BXXTLvGrPwpHkRDsAGrjx+iLWOUU+FaFeSb351
7yypOjnXWReyhPnNAkXUidqdnTb5wX5VDPUoO9jVPSo0rSEwd/F7rkBVZfH0+54K
/jll5ZMy3So14B9WmiaiEQ6xBT+XfvXRfZIx80fZjVFJf6+gH35NH4cE+8fY0iBw
a/hz7BD1WoyKdKK0W5+Q0BftD4SEthTBjUGoVS8kBwpNa70nfCOy7TE2v87Di5M0
bu9WV4LCD9TfI2z9tm5cAmos/uYXcr6ryV0Kf8Rc5YW930dp5LocUkb8Znbkl1/5
aWk5LWjjzDrgXo9C2N5oV8zeorAfr7UDN/2e1lyjTTjhlIxdFDnCsqWh6hKSu5sY
dvLWVutumv2bE0VdI17xfLnYcUPzNq0nWMXe0UWnpI+7fKVv8DvVV1vor1nlBJtn
CQVoFkhNeb5r0ODfA1SwDOSex3c+cUaVAiDPX6oJmXGrIur7uNZ2t/Q4P4hJozSN
6H4TA4y2BwUtjDO2pt3z4ylwV/d6mig2sOrqw7q3pXUGo99oGP2CJXqTv4k0D7We
/LMc+hKw8cqNLhKukyCC8uLwL6B6g2k05Di9umSd3LNzK7w1yqNBOKGG9o9y2Xla
JW+OwNhF5QKcbh+PDT4Qs/h6VDNGEuvErYybMn8rXjMar/c2nN8fY7BFpVNEfsLD
N9M8OQILC+vdsEOifXgI1D0ov+Et4VeTqVKqDzRiL83DUGtdaG7Lgh3j2GmON0Wl
VpORlcOYsJeSfLBzmUqqSNj0H9z0gSH6pQ5jLnhiOr/1PjvEQzKwfFGLYQ6e1RFc
eLphZ5+Xn40I4mI8Ashi+qWrdWQCstAvnXHgSOzausMAd35WkacSWIR1AJI2eobe
lHQqrlXs7FO+gHx0/3x/qYOnpPiSF7dduDFP7VCa9mw=
`protect END_PROTECTED
