`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kan1jrG2z6fbOzZlo5ZPEcZg7kxjCbBadaa/N4QNpvO1NnB4Tn17RPJBbaEje2EY
sj+1I15r6Sw5bCGQS2Sr69qD7ozrf04VuDYw6ppyb03N9ld9AYgoA5sv60HdvLtW
uZYY39DcrrRuw9gKjrDY8yG7wuaxR6eT1cfeyAG9OpNhumAsoihjQgLJ6Lpo/ovW
uXeTety13RMdqUeyjZDFDSpuJYJDqwgQO0v5dob+ihTQtqjyc66GJxnmxr6dnZRG
NODV07g9+njg/CUXPuX3EBEiW+s9sGIXoONIUnetqW8A+9dcO1T4RnIB8RsQS3eY
oWi/4vQtrR+oeHHi/kLw0P9B/YxK5TMC7qHw5cDQtObxixRahRlg8o3aDGRoCWre
tjJJuOQN2K+EUkU2Suz0MMAqmwb4nhAP4hk5A3JsH6dYEpe2a0/eeh+qCvdbCacE
kQl1Y5nyqD0IK/88TGkORS1b2paRiCx1fYmKMERIaQKXRALlBx3uKqOlk7LIqTZ7
Q1V36SjaH+t5e32DyEn7W9bcBs/mia03YnLy9I2ejHGA0kA5Fp19mnFc4aG2FLLs
HeoGJguaPVZbNd2CAlDRRsXCJ80V59KYH8JCqSH1aWsVfBQzbI+DMwN2oGLFdGMR
gSHbCWUi6Av0Sl9iGoyM02VurNpwU7iz2w5MlOLHSfQDqCF9OKecAy3fd+NfEJ9v
61bgXtsa3jZRTfT9mcNRvcmvFCHRwVM+UCUFmvvHt0/PWNqbkzqrzJVIiegTtXx/
3CkEyEGYCqQL96VsRhmPBiUVmVnfKrir/NDYJMGv5i+z8aIMvOMKqZrBBgnKmnNO
A/XEF5FcTq03nCR3mcP+3MuT2gXseNwV4y1MGfj5lHLkex5BIAHvaD5M80BnFglB
aN/9bSb5/vrvNocyyQ5keffOOQ3hoDYK9yUdwxnT1Fe2uMGok2aUiEoecbpzQpMp
nJYmsaPQF/vbU/iSBGZ8HZV2Pksf9GdxC9G9wX1fzbXZHO6pcszpGwRcWjXrpDeP
MzzBajamgcntAt9YKE6YNpM8xuDCJT1+hcT4CADVYyThWUAXqEWhILS9vuLIBVlv
uth2jED9WecBtZneEWa6rKXTAxGeZFcd0viH2zWDv1M0XZV5kDq7N/beNV0T6pk0
yxn3uSfFr6019mEjgeJHOO7PK3967IP/GtoMNret9JUPN3frza43naAlAR2AEjm0
ycSjKgCFmYIPkHnepwO1uMc5s+YSUN6EGH1XpzGyZR5K4keVJUot1DL93+xtTimI
CfFXCLtfuh/VVaukU1rYHxai1VosSqUhDlHdt8w5wgnO02y4btgxx21p2ZblYG1p
08YArhIQ2QVjRqRQdQNaRjKTQEATrz3ObL+2Nv7qfg0e0HemDbnEF6RMmR2Q8j+6
PqRG4PhZ+36DFXjrq3uI5DC7ObdDw8m8EBo/pTDJm92sYUOkB7Bzy5/nSHbAVOjC
BncqkiqsWdC0IJ5Bt+viFpE1k94Lq3TlJeiE2Tiz7idahWAkfoxMemD4wA8vWSse
6Qe2RPbARnrYWeaJD+tbrVWk3dAdGp8dS86Ne3/BI/NE/w7gpemJlqXpr6wpmbfz
QqyfVdIMm1jXe3Lfuk73JsIx6gLSz07XjDYeVJgmrzlTIY0I2iicnb3UMHeuugjr
8R6z+7xSZpXdzSCdzhujE5r7ae/FBFPRYsw6JbWEr6zhZbJj5YUz0TDM7XB0/tFD
x79Xk0NZT2KdOT24EEtxQZAVTTpJAbchE7lZqFksWB+TAPfWjB4aez/tSoyqeNQd
X1qAceM5B4oOPE2NiXKeqdUMKn9gL8qn12z3kNlfZCTWYquMBNn2JfXJsBGeWGAa
zNxBpNM3fVvyiso47NMY+ldpCk0mnE/Ol4XxgVHN3JWiu8s+uR5oK+EYz1R2uNLw
xgEJOr6MV2Kpza3THjI7GHP84tcuZpiR+VWczW4xXdJA6+9wTDoIAM4uTn9gRBX3
iRBA9s9Ew+pNx7Lv9gwezF7Ewx/MfXr3HLLjV644I4sUTBL+vkE2vnLD2vknvICX
7rAXEh5GfztWqRM5CqQnc1mfbiPkc/AZikLZesxLQQQWFbkLjwM+TmAyOS1dAf1F
WAXhGcLl0HMqGIoKGGomW8NG53EfduMALdVCru4cuqDTd1/zIGmXh82mgTlHSz+H
v7ykOgkfxWuhZsPhN5mvZBjSGULsbzO4yI6XMUA6R0MMxxrFPnf10qRk5YPEQOJF
zRsJ4owde2stLyJp03Z8MNOmZ0FjCBCvNFOIeh/ac+6WF0qPAKdJEYacevF7gDIr
fTmt2co8QBQSfq2nSssgWXODnrgSXtbgHcCPQGW38eO6kEn4xe77uflUh9/4ZkEa
xjl6blCmqQQp63GEx7Sj3P37QLs94e8jkp4kRxXh4rngWJN2bpBon/xFS9l7aWzm
bu4fufyQS8IFWLQwQ6xPfSkwpzD3qUorpmwFBn+IZh+un6cJlao71EZ3rAlYnIr2
VeywNTqbM0dfDArENhG0B/MKRGtuKMKQPTO68TmJxavE4k7qGS/PATD/yU67F8xe
jIJjSTilP945dwQ5MR9if3Mr7ljMF8hm9kGlqMFGGWg3r/q6acz5IJnA6lqS+8Gi
GWG4zDbo3+6goiFLEait5SjPgieVeKSErv2PdkDdvCUVeJnkZW+MxJWec+b4omyf
EPUI8w/auU1ORSIit51tu2dpatc/y/zOkGJrgrmlHBPGc02cvV9FTMB3nT3aXCE7
ceFmFTl6pXlenQZgJ6h9xAJs/URarq1FkLkW2ZVLbIklKrsV1u7oDEEToEMAunxv
i7thoqvCFXyqQXUdnb66dZmVhzNoUlCTqWRVzijODqChEwoQOjFN2W3nX4CtE+kI
Avl3LexHVYzDP01ODT3EEuLpeVA7KElsgntudNcLn8QoELrmHE+0IgLryh8gnrnX
FB6IbiOfVdL3nESR5/j8qMFY6M5tO0SVS+xp3C2Cln64dfXU2fgdDIzs7d49XWFi
QIxPhSnInJ2GfySNhjjVv1d4K6EnW+1RvZfJWgi60nppL1/ryE+9TfuDENpWhgJe
f3SjvluoHltzSF3SyVqj6vSuAxAecOuiDxPL9hAlRXgTkBzboNTHiMu6PolpzVK1
IwA8uvrsGDhrUjBuzXPrx+RNIZFV0ucV1YlcHRKI7Z8DNGGdaK6FZW7jrVd3xUAL
MBvc1P2dhoCOWmx5MYtEoidTAC0x2wlo8iNLJPk9IBvP0oY5IYGic5d1hBD93f7I
gSJ5Fk2Wj/+Hjuw/CqgyUl9DLZc3gNm8YR0+x263c5rfttmrhUElx+MMjGR7xbMs
ONfNgTNXn4axrrEji04IPlGC7mcyDEVSbNe0vf3qHzoa7FoSfGB1p51Qjs+Uyram
TisCKcDOmvDJO3P5HMi/4tV+YiwoiYRZtTqS5orewGryFgXydASNwuB0CQ28ZTdu
940I9n65UNGLhqrHWWMKlgcC8WHIsFuQSljTd5FAML1jiDfj7khcVss8asOso/kK
d1SxtYHVtCi6mOVRa+yvMc92PEhjldracTgNYwo3KlcrTDL7hObV9gOnFk2lI8g8
4d9zWROEYsVK1VvJIFeeWjeHr40ybg2AHehNNPcntlQGAYrFyyEjI6c347Oofr93
NVRfP8n4TUvKozXmOUncopo9I4atdIJGtMCDyyLpLOyKsuI/tPjQZ6pogJcsYckA
k9CUk9QAsxOTc+QqWyKqlYm4HHXFt4IWXCAA3ByaltQIqvjhzuufcBMdRJB35LEn
RQCfJGEgTZDhdg4U9OYNamSETtP8UpCA7fhKRu1a3/pXDHi82wilCZi2fvbEy0+N
ZeOLhr51lHGWPKqnu4mjj51Gydvr8OYIPy1UWRSc0WJ7M532NEpsfd9OQ+LBoOx4
LLS81Wn22F3nZ+3y0eSXD1ew2sqrFZwKNmAXti6xLmg=
`protect END_PROTECTED
