`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSK5YekHub/PxeXlMMcLB6Wl1UVFgdB46YNv/eo16raf8q05TWT2jJcVMNDqq94D
73lrA8LBMA+23JiJ6dFAxTazLBdWr9aI9WQqYwSvrZo/JnwKOFcSBHwnK3wX4fo7
Y2Mc3ddPNMeZiB5II1pXUMnUCbPKodliyxOcD6LLr9cOsVXRai7EoPJ2yDArG5dr
EKps8Qilenir1pnxRFEOZLE03LkQCJB20YfiaNy5r5YW0BprxNwaoOaTvXkpA0wc
PtTdmEDRB2HcrIiCXFXf8SX4ueZa8scfIBYgOSOJrw5RJ73AYI0j2buDvq8HU93v
vvZaHLlOm6wK7sUVUx9SBiMyJXW/60yiu3kQ0eRJ7c+tloW51idPVGCdjPB4Zp6B
Ko65SdnXLxI3QW+rtJPca2G1VSJbz5Gg03sjn2xNv20ruOoRaLJgp5yLyq5lSYbo
V76cikI2MspHux9LvZGHXTarvs7FJiBFllDeKOqu7iuNR+Fg0MGMj+wT66VfHJ4O
W/GsifeD8dYn4Xq0J1BAeLjJL+Yw5XEkrqcNFUs8vYGIbWJ9yzz3CkSipTV/mH3D
W4SUBILXbk7bOb5TCF27a9Xp3HRXQMu761tTd2Y+hpuXqzgebDlYy+iN2O8l03EW
KVpN4kIWdePOym1/Vc4oyKMa/S42nofpullEqzNTfCZmId7ihZFehjq4cxWwykuk
MGNlu97E2hOBHHyg2MSsWHmukve6p0Z7E3oL6jHJRzFZuuU6nOk917rLu2QEbcAp
ZNjJPByIhMOdqxbHy4tGOsix6fuGeY+EoFCVbcKWdOZJETJkeYFFi2888BqEgmwg
MbCh5T9I79MnNeqI7sQEUZSfPvluujkYwMAzEnNDuzrqqjlw6TjlGdjuq259dS1C
BfeZHwDhSnMchabkBkxc5gRm+ffdhzXCNA+9dJfjaS1n4i1FhI4JJyfwsk2uYicA
LHR+GPnsVejzqrAl3rjUB/Pj4PXPGVZSQ8VYpr6o1E1Y4/xdLcoNLBh4fdVoVLwc
i40MBscaT/oWJdjENwlP70UnG68pfJMCfz/KKqIOsM7/X1VJT58R4Q5HTr7PnBxu
l59mHTGOm1DtXnd8Ra5baVYqDe5eQq70dN5EPPNTR+ezaSVnRZbkQ9jqcXJ8GEXH
+wQglHeLdSZYjbYuxsoytG4ZR3CRZCrnno9PEs30oakKkK8bmgF9HZbNvP5hsjQI
rePdljQ4I/GGHnHbZnl3Rz2qUihAnQ8yctqkSLsQTdweghKaY0YpC1bE+XX5hS1j
kmAAEFRLey1S4RQHua2yM8bGqROWDQ1WL3xz9V8o2x3intPJJrEHzhw7r8H5gRzh
GjOpqdaWhxtcMskTUcohxfcYVpmmz2pB6e7qfkaGWPTubvx/4v5xULAG8xnXaHyH
G+sDNqQhjfrII1NDalan2+6pPGU+MR65pohnofrbQ/NblYLkCPUwGLmGtF3YOHYV
M4SXLosDwyY44ffPsoo5Z2uhuSq/A+aog9N+IlBM0la3q4+1xaV0OuA5omM2EZiW
v8xxWIkBzSlS5x26iM9hxEgdj4Q3pVivvobDuWwMvB/tkOJPvjt5wz5H3oRLUnNp
EceBiWVD4dtXxPrUQczR7rdurOEK62sxYP8pMppSUieSrIfkGAmlhpujC3cTxjzB
wAuHFvf3i7devKUyDQCqOHRdG3maXOpMP8QcY9oFGoEPxVlnhIQQb5HEBCGuwBL3
zXCnqpDhipv/HyclEIdRMTJCm4j4DibUVpOTCyF7fssIf//Scy7K7R9QBc1qtpQg
j3+bKLH6zM6VhbOm2kXzNcyWazgZ4NAQnDjtXa2u4TZz3ObR3c+nONUwWBlIqYsf
rDt2rllVBVvw6qqJ2G0WoE5lXeWrEOn4lyFLuUstgwJhlEHW4MEU/3sStdH+wKs2
MwPj1Plb8y6cLMyMeGTqYTgsohL8j9A1u7qRYvPWxe2fvmC6tVKbKl09bhReODuu
wO3g3e1NR9Gl4LxXpCybZN/08QFo0y3di1xcHR25CIfUZyX5z+8IJk9vGd3Rm7NL
6CsUo9QnQV8eToo9cEQ1qI4xJEzL379TL+375fOdZmWZLPvrrXzXNHOXu9jqPQsg
Hnw9wUvsSVxqyPtuonB6VH+jJ7Y8GKtCUqSkU47Io6B73PWcsyMhYZZJ6I0BdjW3
fdFnPyjYF815F3iWfsQf9dixx5kYV57fJNSBIz7/Xzhn2AA2KReCVjE7bLqGE2BY
7SkdpvTirIXv+b5bD9kHr385Tg2TqF6Z/ej7VG5YE+45kZMAjWK0D3GxWZDN2cjS
6NEV6wqYtXOzipCYGZRm/H7lRPj0+21jMCKJbKWSqTDvnSaM0MA6n4NzNHwIKe1/
IifoLv+UYiRsCi+bVzLLU5k12K1yo4bMZnPWx2H/WwWW79pToRm4atlQDvKSdSMB
opCiNeShVxEzCdx12WjwccZAIqpsucc3bnUIqsLRWDgKVEg9QX90cNxQUG2GloOW
qQgbGTmQ9z6eeMw0OVjoB7nxpu1rr05F0c0tCKTGaDPqeBUFuer/yH7YXs/2zzA0
IOV1etzrxHG8xmnnKsju5hch3NKhzyTltB0l2GunC11hqRm7yzo/IuZWTn50aIFV
B8qJp0v2U2+sZkFKfPio1yLx2THX8bKbpsL3kriInAJzc09qkpWakbV8A8u/GVCS
wg6i8AN+mvpBIEFglJ+V5cT7qM3uWYXV3z0WNWIYeyy3GmneJduYi6038YYKWocp
dk5ApyTJokRIOGXWWDjBOw==
`protect END_PROTECTED
