`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0TOxJoHeemO3nGk4LDA/BbJ+k2xuu+SgLkObBepfry0QlYWzAAsnz0R2Lqti4Ay
Z8TZsOzazbre35FZa9xDVNNFqpSt5ZYSGMcWIiXd7Mme2p3dcli3z5jqamIprQ/v
oWKvCFhui7MDORmb2ts1bvUClmjBgl22P3FsN3KfAsXJW2Yt/cX3Bn8iDkN29NJk
x+OdillWcEcQDzIBICts09v085LtMYVPQpJph335RAUkOkaKpBIKR8o/R1Ifj9E/
+Kz9zgpYFdNOdekbkRNNjV38bdD/8ogsektcK/160ernHekb3A89OzOWgYlLBYi9
wt7TkQU5mRLrHAwKH3jxIgWJ7KlzwwZ5y0I8qNGrerGs2Q9tEdjPROUBkKgpCsEO
sGn0znRtOsoP2AuoWRby1OSvSwjEKMci/CFVE6346a82nK6Dq9dGD1hGlKXGfzmr
0tN2Skp2022/L7K31hhBpOHtmdtCyp2GjpDddGkJ68xFEhQk03sxKxvZwe6SZSGA
IUvcjVvlKfrh6IJcrWfvMnhmRPmnxtEr/Jifc5KGJ9IiK9rhgvY5/P2KXgN7Kdwh
lMILTrf3dKcOwLZXfMyJKPnTX9oujPtDRYwEHQ6igIqmKntut7Zeps/6Mt01S06A
V4KAbpTqqciz+Q+/DJnj2RCzWyiFai9H4YuCYBjKPlJJK+MzvF/fnJx6HDpMh4KH
qmd5X3Ug6ZoyIiZjz6TLnmdsYGXYsknNGL6g9adJKEioGfcX7jVhVVTvD2Hq9ZIm
6Xs4fSXMkYLUtt7H8cYb9W/Rrwj44XnRi+LfEwnpyDJuwOD88Sa9ru0KfpxQlwQn
EbOIjArD6e8B0T2mYS1+U8uAw/egjLMS/Q6Idq0/J3I7OJiG663UL+j/F06COKGV
KwIrzJiL9G5O5ObNy8iNwMDTND6yZDs+UCbKF2H/CdXDVqLWkZD/gt/VQPFvNB/K
20ALMG3QGVnSXcdh2MvrRWbgq8XxFO1BZplZGTVdnUrayyqGfhRbZpLe+yq//0Hr
a6gxeg0uhdkBlpFnleI1T3/8OsBurOhpraItHfsIIexfMWEgEe1px6PjHNjmm0I+
9Lh5/LlhDuKZOAg/ILX+GZlNBDDzqq/J5tyR2gC8o8FPwDeFDtU+UZ4JH9P+hFTf
YS7r6Bz0C5VtvxDnDdFdiFnQ+IzwZptFq29bvZQkLtcMpGKmFFZw0YMyOAHGdBMd
jP3TFL4yrmrECRrUiRw59kX40hJZApkdbg29530zIMIGhXIIMQ9BEgn8iIKTlyTv
cdnXF8EoW0Vrs7Bg0tlVlbhDfzf96s/jzpuKjTlfWDXWelXxfZlaa/cVJa1FNhzL
soIe9G2VJ6+Li87RRRx3w4u3etKbk9A1XQ0GZkN+b7O14Zgffyw5KakWzh7YOTmp
bNPQAujGNPp0NnwgDKa0LQqoz9buV+bIKSMMQsuW99S0HNAzse+0asYbS29SmbB3
/yQPnqKlnuu6Dta7Unf1q+dIhWM7314/cXCIeIaLWTA8IxvfSv0Jci1pob52rFUP
XK6UWtpKKWs4SI+Rn1JzXBnquMQ7Nj3VO50cV61+1aR3B55JAm2iIDXWyLrIyQyZ
fAhutZagjUh0O5rGjXL4PD4l/wcg4+r0GtqZwsN8ioyDbvT6owi5oDfNvbaRtnqh
cZ97cAhTFOclm2dxYLKV+f+IiPtRsg6b7EpAtqtrPbOH2jl6QEG5/YsR9pI3NcQJ
Iu8MRz/OERS+bu48a54/HwopHlidI42gLxHMD595CuBfo0cqqmu/7QDUJJw6TaaJ
tNk1DCms/pLhXo8Lt3t0mn4chNwTu+hQ8HFMNLqo1MCQ7HGhkePPB7PBVKs+3R82
G6AVY1LWEq4TGnYcn4+4GIjnW96JREs1x/VSSXuoFIxrW0cqBG8upAV1g0BZum8l
KlVJqS0xEzUqsMF6u2cdYnymDIZZ16xvtcIH3mht91TWos9JKWfdfwyfzHa4VY37
V4g1/W5lcEiKViPKy7IKsylARD5ZYrrT7lrI2JVnMBzjnmMxuidC4QHX9Zimy8zC
VpyN5OUezEuhfQ5+/nRD58hfXIyxexH+CowmMlUPuDygGuRmYjk3+Ot+ADQGkwtV
vWgvgmB1EIoHCUyiCXtrJH+t74At0n+fcAnqxit6MXzMi6O1OdugJKNWFPj1Ukum
AhumDDpwQnbSWUjTceyi1uJMOeuujJn0iL+FHMrfScqwp3KzQBIcFVU+trsMHnGi
vEwEOpAnFnH0bbT2vmxpSYcg6E7Myj3tEyk7QGUtcdGg9GdM6PR6Ck2gl03/1rVG
x6FMm3GoZ7TCANrWRoVeO+V9pbXTRE44JCNcHojWU21IHToa6OdakvR8wW5i0xG7
9Wi4Se832K8vVOY9mzar3CDtSLp9XKb05TH3/mmLoD0CcVxWh0qST2d4ddx5P77G
vSAI8AK9nl1Mao+t2po7OH6OgwofUxwdTdhatD17G529fNOfJAHUKxx9JrVGDOxe
SLaIlyr/wJOIFHDlHO4NyFNfYjhVCy6eOTCwv9Heyi0j/dIt2V+ZKP2++kaLDq8t
jpJPxDmW3LfwZo2giNx9gGSVA/iM1l0Nuvs9VP//TtxA+nPPBzZVQwCesW/5UZLu
4Qv6EPxVR7HeQNByE+gna56/whKs5py+eE0jz51KjDb5gkgCuvJKYgJpZcx/E4PJ
z/wYjto+2X2lz9r6WHuoV2wJPL4m5/vS4zqoZHy0s8aOqIaq1sVpVppTxMYyBmhw
Q8aiRgiiUX8gRp8ImWe0tIR/cyxNAlr0P4sQEdB/kCtTuzzHDkg5tmjdm/OYTh+9
u5ByjbVZeRcCld862a/lWsy3bi++86nYuRaFc+lVVMbqYXssouXZqDmg5ZEFPt4o
MzHokLf+0ayc+LvrK4C4QOVeCMs9xFd4I6tG1m6+Jm79OssU8y47BJZ+Ub/xqpOu
ZvOjLIM9Qo/g61nSwCmyw1hMQlwJVz3PCLRW9WL3BEsWscbBDdTP4risZgOe7lqL
R8qBYUsrVuJ+tGtP4ZEXwxQrAyISDdz+EvXuElPLgKOMqfRzpGuYjBnBaYN8VU9D
alVshwQWPdYvYEdRDYWfZ1e9rS2HZVj1nDYlZUWhZXchwTsYeGT51VNRv65S5p3m
k1rztjYkm9xipxY8TdOhwL2ca6Nc8Gpz7zHD0hq/1Lf955ndH83vZYL/4ndrAyW6
z9BXdfnf9kt+BoIKhCKqZeVhRTgT+XZ+n0R6lG5n+l6tNHP1cXm3FY41+Is0SLCP
viQaHcQW0s7E5sl/sE/7WsNtVzYOiGv55H47K/quCU+Wxhm2OeletH0IWjL1JDCW
Uy13PPDNi5at7XZU9Sxize2cjeYbi02cMZh7Gbyklt1pBIKUvHHgWDweGzj1/BKD
3DEYietRA4ZomJp3DPMcJz2I4b2rPeOrdB6RN2kjWQPQ7V1B+WeBjUU0f58DeNoF
yzj0FtrUH9n2Y4YmxWjGcBnupYp5+sfpnUVDYFv4NoNgZCQixhm9pM9nT3zXt7ue
TbpKFP6hOjsai9O6L0eI49v+t3DCiePWPhhnxx/bSwKrZ4HkT3Tw51De2A0kwTC/
7r7yEnju6CRqdBKFRUjrq4vOjM0fim7OZKtleI3kF1Ps4BxhV6b39meyWoz65eA6
QjEoMxAJNyrrFh6Cunyrfx1Kpb9o02Moom2dHItNHVisKmpFKTQX1kuYzeKZJmS6
ZcNY+hGoGPLQc++RrTngriRa77vOLC/KaRYH0MhsGqPZKxXVXgbYRxsoW9xqGL15
RPy6dt8d0//LkKypFxmYO+vV5BwfHr0eXPnWxcRfxAqtNHBV9xPvyVS2UQxcHwkK
KsvE9aiaHlssk9eYSTiv2OM2aSPl2GPV24UB2GDDZlJuS1idDw6cXgyXy8qtvg3r
cgynzhAtwJUY+qI9xmOGP9rqktOQm7fxPF7hR11Ue5GujKdAImEoXF3vXLYotYrd
iyiAXSOSLKqmS+XUpEFwBw7jYNDMRtybDwGkxE8126kNx0MmwCXqMoI2sZKrpRvS
eIBaoPxMfMQ10/C81iMFwKQo+sMc9ZAicb2JDMWkNXW1XDa+jPBGfXHmYXm2k7Hb
cNi605087O1MbUyi6a4sN/N6Z1lHZJvH4ILszY/t4KFRyH0GayxtlaS89ZD8MNeM
Z0NLuO6pRe39n1COLtWJ1m9MQS6XbCZovEkkFD2hs0z3Jm9uJJzYpDcJ0gI7lN38
`protect END_PROTECTED
