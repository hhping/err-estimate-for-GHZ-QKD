`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7jUgeCsu2QcvPc3oatu1nG8DVLbV7yfEgV66CqqqGvajokCYVDFpnh2bfymPvy4
644E5H1xBEkZpbmhZnC/zeVIWAlbdpWBp0HL0C0doOSSJJTbr6yvsSMy0Ly/Py4L
XWKGKAb+xYMIFrvXuzgePi46X8H2CLN40hFpYPJW8xAbtcTJCNHt0rJIthoDqY7J
PxysGTCq62O1hwTcofSntdftTCkuWC2lizpBndfOpdFWbJUWgWmzD4DVHNfF9kkv
knOlCqEwVBRGA7ATf5NK17Sv7gZhziwhJiW/a6K2hLQuoRmGzzmSHsbX7/XAwMds
hcD0vTCAmfYoQm/lO4igRucFya5o5mmtsJMK4ce+J2skfDzrVs3tlPxBqEguqS7X
MIdplUtTRMcjvA0IXktW1L+EAIrSC9UGpdAg9A0aiR1ynanyzy+Fpz5NvPnBDHWX
xGuwIMAN0ggwPdr5zjzubEJHKlbrH+HK70kpsOe+Yr8fCX6pv3668be68qoj/MES
hBaUURSTO6dx1fltjmg25kD+yelWveHTTjF3+7UutmcvmQgni9czHUK1aiIxt11O
N63udV37Kis3WSWvWJK3sQ17HldyA+z4+9D4LihybbYCmTTd4+X3D3656fYNZvpd
IM0SJz1QV8UrRpu9wUMiWaSiAoJli1D0Xc1tSegnaXc4ytLg9gkcLULxpUTZyRup
QTWEJmgUMLMN8sDz+nrA4ECNr+20YnKR2SpcYCn1oxoLfH5/f6YGkyFjh98OjJPA
4zUxNdPniyvDXg7BwOmZYLJzCdxlkPSRv1+lR3dKtgEF91RiCv2dHI4o195I42se
M2xRctiqGNqRenh7mSWbiuinwBxE+GJM7FKqV9zwqi4=
`protect END_PROTECTED
