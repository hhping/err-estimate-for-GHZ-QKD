`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/9mn768NTd1KsmmQr+sLZOOpdDNak/KLxtOB45+9AgRSEiS2eu13LJmDtvF/kyMr
OuxI49scdW8WlXTEB37ZU2aon77OjHwJU7GFyFvLjLKIBkz1RV+7MEbt610lUm5q
JkJUaX/sFsQSZDt7+NCDwgE5G1aPwlfQraEoPMt7FdxvjsocWMMLcCTK5T0VFn3U
3VA9CxAR4wZWCqmyvKCzgZPrda7JoKGNJsExruSI2xr6oklJLupu4vADc02SfjF7
FCYvc7s5Phd15e20y9QfduSHzORWBxePtCRdlXrriCbjqJ8iLuCnpKAdJKPrwvSN
cvGc/UjdC/293NT9uBkNk4VVoQjB9aO7QCrksXF0rPKfrGis9Pj1b415jXSo/aED
WCdu0muURZqkhjUnsIaDD5vohb2SKzqFPX/RKCAWra8NiWeH7ZrIdUL4vNIhC3gO
V/S+y4msNGIUdhOZckED+h0lo+nn4OePHON1hNw/zR72UQdM+yYDM7HgoeZfol+i
s4Vy+M8EuwgaI/V/IrhV8tbHQ1vna0nlRgofVkwfa9SVeLcsi2doYvmE/iPYXuda
Tyf6PBk5maKSz/Qncg7RDsXyh0v9QLv1bHkM2grqkw4g/eocCn5yk0oNDr7DcUsp
Xkhahy9KRawwlPtDF8AD/5p8wagfFzawPMxldOtikgB2o3zsefh0h2f3Y+XO121V
lBLYC0gHDRQaEVPf39trLNS5NjaqcwXZhR0nqDhPOXFlZXgS/j22hx+NdZUDRpFl
B30wieJ/YlkaBvu5b82xmd7ky9QraGkW52s5aON/jSsoXNECqxvhie7mnYfgCl/k
O/o+XZVXk1syhUUlZXij6SszPqv0i+7TFSXGB2MECnapX9ugFenq60R9Q6FNlUyI
ZiuiIvJb3CguVhPmjVkyeuLENJZnwDLfNeA3/s0JEYIagBlCRbu41d641SN3SCW5
anSRL6A/tPGXe170n5WVmxnwDaDy9OUFV7SIeOHje2mfGhrQqAgsFezBVncAAg2t
UaMNil3EsYz34A/qCfBhD0rP4/usiY7LAJqQaNwqX20aOZdJSMaTFX4IhBsBzqbV
Z0uf1OvPT+7WGB+dkEhBEAZg4mdX1tP/QYGD1R1+4xbjfVAOeFJh8+qHUb9KHatC
iwBI7HXoU0JyMw6Sqh23gVULmw6j0/iflDHwtn7b6a93YZ2Ib0BU3gzvlk5p3Id6
Fs/Szmyc8qqeql5cByhBdyVFsZD0WZtsnZz97GrwpTqLKKqazK1w+EnrB8V0V6Iy
mLI1EnD6vrUHPXHG8NxQdPGef+SSOI+fRAF0CUeAiCJXIe27F67aVfo0oWu+9ute
Vv/oYnKbo+M7S6jsxe/A4bsETvzBXlWc6+wKLRrFf1McioJOu4fo9FsdpjT3aNVa
gyWto1O1DTKSzBFmfeDbAyYVsEE1uEqWIvNMQcP8IzDQSFku8sjOvdwjrjOrCfrQ
`protect END_PROTECTED
