`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt2wRS/ZMcU7qRR/DFSQXiTrMV6TPdjd8UhNfDxbSkz836xYZ3OAqCEaFfx6kAkG
0jlALBjIcFsDnXEE3Ifv/MhPbDozL443g4AAsOUZG9smZxF1MnK0r52M73xJdtRW
gjVa5BolToAKtmlerYKpZvkhbkiM5wQqymaNopu+ZxUxzgMjG3JklFjx5g6RrMqX
YdPN5y4R8TFhd5BpZUmxYkKuaBKm+qwrCEU50QkN3QNRDodGbzzQMIk5Fcam5ZS1
LmzEeDuNdJJ3V6u1JeDLmp5X2ION+tip+JohEqyJN8MplTWUzr04y6yyeSIdRjM+
AIbeAr/iWW/ZthO77ry9k+E9nETxTFs1BahEAOtHzE50laA7p5duQqSxK1o16VnV
3D8bBsRYtOPtTLFJUfTyXXGTR0acXTIlyaOoLcDK/tPmeAstazENey2jj9jPAWoW
6S67KOfAeeGcBOYa+mPWUl96paNjhtJptFz0xfPRcWtXIxyhrGPTq9/7W87T0ZOF
/GKLK5OXXupLuz6/00Py6O0EIB4Gqq9v/jwWY47cN/lvia9mt+/ambPt5rVMnmP2
/46rZbIFFGNbrJN2a2qb53lOWMY0xiyVtL2aQjO7L+QrtX/KqzgJyOB76Km8xGre
huOlNLQ6Zx6ddCANTh4JWgZm22V1polN/67nkEzyeY1HpwGQ5qsLKcv64YGWkzif
4SvPhQgxr1605uAUhtoqSH2B/YxRSDHQKYPojfPpv758yXcZUqGZ+HdNBI8hEBdN
5wWOjhZlbJKBq8sOVlh+G/547D2S1LjvxH0vl1nExOB+XoLRi4C9kP0miVkbwuys
oifT61vx7N0nCVmF5NFOU/b7vlJblZYyM+UVDGtC68OUfzQMYe20GZ3f2g48H87c
Wtt1UBMgzICLt0LDb2zwuEiL7bPKgxhuhgBoWK+s8/7G1iauZ1fhCYOH6qVzoPR8
GC+yxsGTlQI3jkjgG2hoydvGrQtez7nhyGDzdY8NLNpMCKDe/HtW1DTjcWhsnl1t
zGw+NvOGIzxPouiPASw319BWt6eYL4JogDbnDfUAplGfzpEVXgNb7iVrHBs6hFE0
XlZx39jadFOiI+yh8HaP8B/3tb57wBAfRGPnpRhwoITmbWTv5N4Ml0a54lQuTKmS
MmwweHohDBNwJP8U3TJn8ZjHCIleNGDkhHu2C74cq1N6wI1ZKWFWrrp1mzP9qW5E
Z3YZzdZ4kRgAYOCvBGGl3+Q4nRPzPnB8B12bDKFy7V4F8h26xAYKKa5okWtyzqzV
hmH+4snUTW72mzY6zbJx6IbPo/xxna/4WIekrhNMg3Fch9y3aaHTD+eNLc+1bMvK
Gzi++hZK3RBg7qEjYO1bYargDCCcMk+byxS5so7eVBSHCVZjskwTdD4orgfCL0Q7
XyWW0khS7eranSDroOxl1sR9h+H/N4FBChB2dntZJh2Uqab1THkbsoOx8c/33RUH
rnrrpNF6ukUg8PPB+vTvuwNcNPhe4Bpe4s/DvWNO5khA3LJV3w9DzuUgoCLqcfph
95aoOG/kdHczl4yTPAfZzIKcQH6wLQ5gnUbcDbNYf4ZBaWlMawd8KoPDe9is+wUt
8VxG1uO/4CYtIKwjRa3yOqNZywLz8/VBl6nM4tq+EkW7gysQCHP2KUscTUiT0j4g
tvXYZCZxOpq0Lg6ALRTu4Gp+o3ddg7onVxrEh9lbp3qcK0vMR/Wh2eWGmv0EU+Xv
8pryzmebsWbfvygvYjtfhsUlWlSUaG/uUNoYfsq99EGsdpEsbmZ0gcgv9vF15lLi
QF4j8SgadknACLBI8ohIjZZAMD5NNrfFdGm/V4WvanKNTdn7pszN17mcQZTTXCiB
9mWVT0Qy/Aa6CDDvhdEk4hK6dEbXX+fE6jNJvqY4pic4BCooisxRwiuBQS9GdPpa
4MVbicr10j+hozaZtOki9neinPftxr//lcHozk1HcV7mwDnwRMh7ogjDu9CArPzt
vZGOXBdqqQUJ0JsvplMMuu2ONPl/1HcutH+a0exn2qHKL1pHQyJv6xsrOontxCIM
tX+rH51bJ2M5m1centVRPz761arrm/l4467LDLZwnbM+hL8V2Yx+iAxByFZwQTxv
8gscUOOtuqiRoPpmV0uUlK7ZP2UE1oNAiwdy9sOXZuHKauf/JrkmIitNjcQZenYS
Px/5zR/vMB9n0sE+ITEUAYaDF3KJrtuWUJRe6dMDtczvWvHE9hMRNBdoDQKNyS/Q
NEhctDqQ1v7hvjX9xTfCRcBd1rEN0qmgvTmRH5uZG7CK0M8IC37Q02vlFdnXSBN7
U8tNeYZAKoSVn4GRhq3pUTV4tlZchp18l9HBRkyT4pYrPuMBjBpVpfirYHlm7xNo
njm4jrgjBT9PSQ+ATDD3s3I4YP3upQljH4JLsBmLxtpx2K8HU6TUy70TytQr1//P
k7mJhQ0BpdxwcMUnD4OW1nbJH8NJk1FWGn7ayO7JqBtlnrAk3Oninw9MSccxk8np
bE7GaPgYem6HzwCRYP04w2CXK2u0Tttgjs/yyP92jZ8W694DNhcw0KIRO2YgwTQc
1xU564NykKNqXIA/ImbONmTAtJshR28VgTLEoJyqMOLqxwNNJxTn3QfwfsJA7894
+xb8CGgvJWPJsxkn138Rhqi1vvoNFAE5d/A45llBWZWM/Zsc6ReP0ZXiQ55wU5Qt
PwPRZekZgrT2hiiPkSRD78qNpN55IAmQLuTsmlL6xu37CRapgrDhGwG6QQQjlFIF
B4htS/x9Fby+GTUqfv88e6Y4bNsUhXy7BvHrDo8gZSTtlkh2a7kFehIvtqfu1jZb
klXLbtvDaM/vkOg0IdTFTUMP1n+rp9vLxoGwkfhkNy/NAYJHnoJRpJIOFJqZgoXm
jS986HTxYxTUfI7K1o2aERtMdMwFNXWL1nwrfkGlIXofG/HANT+UGKGXO6o/GxMj
VhpcCvwD90uGrnZ4DFlvByuhqrokvLWylWHTjP2V/QzErDgFCt39134+CsJwywfV
wceyZMksiybyIFXAumhe5k56iJ+PnipnFt+OFN/MBQqxNZvbjlSNWilJhEFhCF6I
VTV39PFb4snfnMY5m5ea1zIyMihUtwWv7UUL6uODTk3DXd4jQdZQNCoh49SQKygQ
x/42NshAFEuAQUwcpU6K7wJGMmJ9rNSWjL1nH7TCb4rU1dhMO3f1W/qaXzDgrjGb
Fg3RgDKinYyshDd2l/Kyn0GJQlrBpSISDPgs46wJr211i2OFW03jlTKnR7qKvwRa
cdvdQyv553TVavJi/IdA2BCnTsbIBC6apDviHMLMJG/3D4x9jp0PaaX0UeFxkK6r
jfAGBIZt3W5FGhqE9ZQkYIJDZPpxb4TB1qClEyK9ulfMz3DW+JcfFDJdp/mr9Z0a
cALCMjXxeogVNNH1QjdwHkLhTP6r/VH5axzVdUAXFH5X96WcGOhzzDYxssHQA1Eb
UTZt+d+e/yvQJ5i+MTxzJfiiIzLB5XrF5VYsNrGwancSxCN3LOEqtt0jg0Y976DR
ZYGVNCPS5mys9QP0WR8T5LqRLKuVP+m3Yhj960A1K8n2ish+hUhlV9+ItyoXpZ5p
UMvjfO4V7e2jgKVrwa9RF9Wja1+pK+oGoFpLti0LsQvY8rwbyDeAcso2rvwT0/0K
l3+zaCQrTSMiFOtrOG3V1E/C756uxzGe2ffw/7K2YKUe366CxD1KqBh3SANGeBCk
QDGZ9CIEpeoeSHZ6x8seiOgK6OvhoPCNrDX5g4nC/o6V6IP8nK8E3VcRURWLl2jJ
9wrejRhHVvzDvTZmKOuE516XYIwcHBDvQgBNryby0QAHL+Syy2sdaGr971JeymXi
CkNdU/zvZ5oMVKj3mBioBbES2fM+6GHBCDhINO01G5HBuDYYNb8wBe/vvyDTDykB
VuZIemZWdyNARJCggJ0qh/kef/o6XgO3e354+wLdA1ADJrhqNWcSgrG6cJU1T5N5
rp1Z2gUoo07q/GgA/zAaeTNug8SKuw2/7KksRPwguK3CjeYZhUSHpanC3ormuq2G
beuvXYhSTtkyJ/Nc5rswCrY4BpKqhFeTz++hZeVyRVzd5fkozBKN51MsgjjPg+Kj
zzLl67bwnO1kLM29aGsf5EB/Gp23I22P8QWYR5uilgzMtrOT2itXDU/Ck90EGw5s
CP99eM3RRch5E/8EgB+GfqAFZsKc/UITPBh2fcPlAg9lA7rvApS1gDZ0RN0dt3e6
orQP3eR9M9uWywsu6IpK3M7QwCm/pcF49q7hOQBrM7M2bOZoAXxXjttTAJW6XTil
6P1PeBuXetKJIF+CqCDWZSB+TVXTf2Gvvy07iJ4KvKluMe0RlA1ZoByKa+SxOxgV
tFupSIgly7ugl4YoKzqWLRPJ45Q5uWtCY3vWT1tbLE0XkPpL0MSI7kl5n4jcboUd
67LT7ZD4yi2f9PZnpXS4/Un4vJadsVh/VyiTXrX9UR4hA9FPub6tvmN8ESJXzuuQ
391IG0zRmrtRz9jf78bRkoICpprZZsmpAwEOihfpltUUYGTN8/B3Bo2oPHxN+qUO
rSeEiUfAaIsALgX/dcfvLTdhXhVwSKwrF7bluwItFKpO088LAhBdqCAb0zprAIHT
7UyXNFh/rIOG2bghsIOn0FiSVxEQ1ltoP323ghGcUIhoq2K/K7LkbXgnVfodrtOM
vH2syvTwXwd5w8t5UBaX4AK8B/lbigAxtqw9/8EjifRSfAa4h2Qv3zZ2DfSzUVAJ
uRO3B7EjtxcRPJdMA3p5lk70XivCZ0Pd51UWG+a15+ZYspeMmMvnUZDa4m6XJn4L
hsRIdz2ZHr2vT52NMPJDe9RDxyKwqlMLLmaa2fjn3oVyc6UL3+NoGIvcQiGFpl/1
F/Jt3Nkxa5IZ5ajkbOs9Tt923vmLxMiltZzfSb87TYj6tj0q9wKZLLHovLxVYbI4
+esyhnPMQ+d6yNhOsYgotVAWoWsqW8XkS41nxGtmmpc8gp9B5QRfyWtj127SZtYp
5mXRxxJNkFZKViVmDflAzg==
`protect END_PROTECTED
