`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzzsFdcgsMPzcDmTr/GER5oxwG6/EHfk2U3V2WauYrgGzgDSMgKtKKOGQ1BrLWKD
NLqGa/pyh2jly9WBNY7nPB9ajeOJMyHmVfPwLSbkFGWJw3L0BorUG7MZsheCJSbN
I+j+nUP6Mc4aQ0NAWFihBsAlabiqPJ0PhS23IXmHHmg08rEZx/oJ6otG0DomINND
NFYk27Ta2Fb2GnEvR5lICFw2k0i3F+VaiL8bVTRPnMjqHrzzEB3mE/WcfP/CtnLB
MKTz5wk4GUw8Gnxvu9LZbR4TKB1YnuHVfD4vSE12KWg6WB2RYZzNDtG7R+YMRass
hhWDliwkAxLQcaBtCBM7hNznPo3WsHiT/7zxmDdz8Dk+iITaz3O1lUGMSQuVxRwF
lZzuMTl+Jylu5U8bMHmPjNUGsqTYeN6QsRMyvj7AlsFVIND9gerxlu6V1rRoKkQd
4PJ5OBghgAbrlRouP1vSB4zDPxm6tLGkTuv3+FELOa66ee4D8M8qUE+gQ79xhRY0
qpRh57dRdUYTY7D3Juu6havQHNAc+n+K4o/bpkk43RzgqXZmjHJT19NAqbWmET+K
vH9SfOu/zYNDl1BgF626FyouJF3PutRBtzd2CjvvxkQB/MkmWLzjreD1dzSp4wUI
7EwFr5+2wP9VGGTOFwmU3rZIYENICWahhWUhydAuGVoLM0jE4xyZLFq9UJn3PJn9
9hsAJNQj7zBP0bCvcTQ/JaZUPBWFCtMTkTPsNZZCZ4BwBjjrJh2MXl3cZ4LVVc1R
AFq/5umIMuK+dft4QwVNO8PG/3T3M3uQjEMX+NpRP0y9cfNULODsGt2mqKcsyt5y
ThDvbIK4evuYaqPYA1iLpA==
`protect END_PROTECTED
