`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5L/yMSrGouW3PznAdmxKX/GhBthvmIu3mW/ewYRBoPboVMKHF343QHrieaXIpfso
dLeS7dAMtQUJyzTys9NDXwwaAksy5Hubw7S9o4blAo1hPB4bGGvlq16FvlpG2co5
2JXP4ynnlKuLzMW+I29cmBmX3p0HyRvukdiG+7PNkL/mifB4qRX1OX/1pGl4XEp7
3u5NJI7SzjNvMr6Ili5tFTRUfnpnhuUG1asQsdYFzM8mBTJW54mH4JFXGV4337cL
TNPvjRySUVcPCwMJ4J8sestqKqKFOlGYSBUns2FXyp6t91LsNkHTVcj/rmHZrkhv
19HaR7m8LftOUgeGJhJp/xqjD7P8P9L5PZ2ojsbbQoqWhb/Tz22Js5kzbx1XKHer
Zy7rDwDr7nUPi3LPlYqiH8gpataZ+QY2Q+5wC0YV3R+vzeuGSaRztzSfYBhkQonq
5ctZH08kM0QT+RJt7nutTTkfDrgdpkbne/M3bxEx42IGPFdSBxPfkMtGPRg6LZ6I
Pd1DGXbo7R/izZQbwAfoRVgDPlLfMghvBXgaVVD6etBKSUTCPOBj6acYOE+7AJGW
dpD7rnPOUC61Yce9WG8EDvXGhEv2HV7tXOCUq1i07816WNAUb5aDVKCZrqrTTXhJ
izd5b/flRWyK9377irdGVwJJthlCJ7iUTWljCv0ATf7wiKCeCjROBJdRe0vhvVAf
z2c5pzr6mCl8dTxwkmTf5vVDC3x73RVRP02Nj4XXkP0pDS6h1lf9xaq19NgNnqtL
Bz4NcrMK3uYZkr8vKoYZyqmbcUK5NdxmCptcPWBVsxZNTjcGoQwLU9RCSCe0gHQV
JgGoqfmDmrNpdzTVexLMBx+ORu5+6D22SR4TF4Wk+qMUF9YTsWYHpJemt/LSdoDG
2rrfbllmI5+6o4YW4XEi+R4vM8IzBi0emcvKEf8q+wIf5yjzuoOUDer+8X8oZgxE
GMPqYgUmEIW7LtXKcymswFzRvyQMAbw958pKqPf3qGWbs0/pbjegLwGKZtoWJGI2
A7+bNYZoCUEb9hguKO42OeHQa7VAOiZh4QD1CM9qCBKnnueN15gkWF42GjSGwluk
d5r4rBcbJ6nMPXyZzlubluMti9zYFWgWRfFy7vm7P5v7SyiiPl7M6sHDpGBYCdeZ
wv/wAC3iXPTq/DaPjLAD1tRNIv5uDP4Lnv3FqxDPHnM=
`protect END_PROTECTED
