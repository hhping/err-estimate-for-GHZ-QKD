`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SjHVcU9nY8QjUI4NHnrNiWE+YGhgOmkT6pCElpZvkUgCcU5/Y+crCB4P+GKGxnlN
k4W6zAfZ8HKOYV16yUiFhGbavB99y1aHAwwWed9nz6lC7UCfn5Ea66JA47fZhOTX
YnRBx7iDpNclhJvvbNk6yd9rbD474PmuHOva8256LPQDJUK7X9dnIe81r2uWFDuY
5FDeOS8ULCEC9iG1jj8NbDFaoElvv0LXX6O1Fy4Bahb0uQayGlLJNPqc/LBHlJ8a
2tccINcOJ/ydndCvTQKHdbmPDot0PwvtMlmddBb1L7Luo9VeOO4pUEhx1sFu9uQX
+RAujBH3EIqJ+oCAVlB8wBhz5T483yZec0vI2xDZQMVVE2VkJV/OOF0vxE1S60mY
NOc3tGAz3L3BV5LszaFWDT3D+nowE84BuFztt8E3uHeJWkXPJTyV3Ptm34v1LhlL
gsl6TFKAAIPYXZpQ8vwS8v54FqjdRFPZHDqiqVilfajSHXDsJRkriREL9gv7fY6t
t0p2Ab3BlYkyQcA6Bq+RxCh7Mo55i4x3QhAsBwCeyRB7THSkSfiCoB8dbrzSss3S
XOlGXF1lFaN7PTff2Nj1ksl6MlnzLD2dXW91wPqwBmUumcVj9O8qZG0Y6sl1wm8e
jROm8us9JXzOWeGItSVAt5zGlSMdhCWocXsUIYZFcp2E4pRKIxn4k73MrhenVkNG
+tVcGyeckPwrc7zchRJZ7O10zBF7nNLBSVJfjWWDpSKGCItK4EsrHS51J7MH14Ml
E20MCeQlhhEn+KH0l5unccLLHMloRMSaXTta85BnU7xSzj4VwEn4h8i7z/3TJwH1
K7LnXHWmF6K4FPd5BldkCdCLT6C6GgTzK/eRmTgi1DowigxcSu6XnZYmTzvCPaVN
ouU4WD701PlmvWQH60qKrNvM7ZOeMmyMg7CSCSUnVU5MAKPzBj8GZCMCXlD8pmYz
1fHN/igodSqJ2JXjz9ZyGid4jN2R61e0/xeyje61UoNntJo3Dqs3Tgq1ndc9/XVS
UzPZLDjp5UzYaIJ8xMreyOgoBM4dwYGYTnIWyrqIKp0METkrCWiS4gLy8o+j25HS
dvVBB/MR/f28s6bkkLLOWBo6KQHy8cTgliDr01tWvS+sbMAqvwI6ZG/RSXlYMHm0
i20W3/lF3nX/SbHgox3tp5tvdisreaWZhpsvT/bVKc03VtQ2Tp1fGq66VEvXGVa4
Alhh84nycmOfqUl6cMZg5nNLFnestqe5npLVHZp1gd3WZuhHs6M11HE5acs5cNmA
HHfF96twpF/NtwTh6GNVp397GxYhXhze9qoNKpuG/aEyiWEWRjgsSCwhG8z7QMsL
hFjUQ+9O+bbv9lmojuCFAW98vNjep79KVsAgQaXnpfE20jMdpDv6sLRdfeEpTtf+
U8H8oMSSRM87ZOJSL2QfKZxxac1Ym8Cgeok5w0+jDcAX/o4NQwx1xULBlS1oxe3h
`protect END_PROTECTED
