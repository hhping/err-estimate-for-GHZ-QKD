`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ycu9YeidU7Chjn9D7Jo0UMhUsNfEQXhGG7/Y0Peo/RHd8Tevo3nxoGw+5Uw0v8Eh
yRGDUQ4yGpV/U/183sWb+44J0HIYVmXyFfDk30TUb4WG8Yyz493RR1335ZrzahI8
YY+BSybz+8JoNwWgIiCKLE2q9VFIQk0o5ajfFVCJQ9qnwRRo5SEyLEjSu26/qkiS
sLmpekVyLkJN1vT4shj4aS68V4F/doLj5yNg0XmKTDwzmBS3dd2zY+3kb+C9KrHW
RvzPICDZU9c49FYEbjtPUuWIFpCvIYw3JuLFGG1CCusV1pQh164izIKaYtinC4Ul
6BrPy/QjdrFYI+bOxArLq86pUlZuQ0VKEBOPUPCFFK1OGVGvG8fcJGXa3Zzov787
VPDOrO+73Vp42SlL7yCm3adTu4Qb9X5zY7V5Ikn5Ueg+zREfoWc/HU1JuNAGLpWP
4EK4PCjKZ877Wx5jZim3/MPO6kMSKlw04zPsNSEwgOtC8e9WQ3haaqOX6IAxsQjd
o8C2pXl0bgdZ6Ac6oqdScJb8xG/4xIuI7ubpz659aqV+U7T0HRgYTXr8pdsCKcXP
VUQJeN3QRB2tcRazKhiKPyLKrFs41Z3w3BsbZhADKlaJv5PjD8HCL5s81oImOfYG
OpXb0bWGG1TrDxoh4VZBB9/XNEJlTMEf8+zL2FLRbdEpclsPBmZh2fChGAzlUG29
F9lrdlinK/qn0mZxtMnJW9yhqGzy1HWYHEZAX3WroSABvhN7kFyjISstuHn9M7JF
Mj6jNj4RlQw2trzoZi5QlirXUDKKzW7lYAxYPldfmkCnHiV7/n1fS/N4Lz0lWj4f
LCcRa32yafgSkdxjk6xlXnNH4DaL52XPBYP4FHJGb/f5nX+Am+PnHWFeSRNgQRXC
c5cosjFEqTFsAVG+AWtaZWrgy9US8mA/kVHTQrUuKVSFdTNxBLJsdW0zbTuGJk2Y
26sgDM/Ys4paCssM8hC+Iizu+gBmbulK/8ijWnYjJJr57u3cpI++Ml3QDWIgDHyD
dnm4Yc9m031A1OkVrjEBBNpV8NOzIGlO8aiP31e01l4A2PVUUfKtzTgA6MAvpnTx
3232dnfveOcLDdk4t++vPUbEceVbgPR1PPEfN/VzYgowA0fDJihrhuFbzCd+LPfE
PdKYPFAvmiOPkGLq2KABjIwk97bdVHMUr0EPZcWiKXmVNe5JMFwMFmOjY/LTlaTz
Tzz6mYCQr7ERzuX1NBSMTPThOYTD/Bp/gJXQBrX3MZG1vGzWBNDO/5DSzFdDoJRL
wYQsbtYmDgvBf5ERWPr0pa9VvwKQv5mLFyQxQasaRxQ2ZCYshkAhLdKUbwR/+CNN
ixX86m2nPTsUHtGZjFPpLvBXVTLB4xmZdifsHLYfpgh8lXgnk19StLr1NkudPcoJ
3nf7ALYZ6XnszrIyFR8aTvLhwke78du4NaROBhC0MiwI/kRUNfm7Mgym6SfwqWpo
l6rZCvgewbWOqGPTwoaOwxzrStkZp2t7b1Y/uyWfC1V8ae39b0vxoDR3JS6boSEy
8JpGyICzW759jKWKVm8Yz0TreHERlZHnvXwUErOCvBXGsLXOSkVwzgGWUXBCdKKF
K1d4E9m2r90OXGMjHkxOakEeujqwNQvkuOk0n6tgMnUW+wrsYB8420HRDKQ4t1pt
N6xqzSJyG5DT4qaY1nXEHtGhfi7vlg5JyTbEnP27S4qtXZN5KLhdkASRUzHKguqr
M2WeBAf8AqgQa6V6xo3+JNnMk0KpDiyeSoP5x0ojRFp38PJ/AC2uIvJFGGkZMHH3
/1z58ShkZxtig4hUVcNMr2PnBazC5HhHOSaaeUqEr7qILaT0tTeZilMAOPLmNkZh
sowrZuuoW8r5rtnhzA352V7VKI8Fsgx6fit9i0hsFGZPX5Sr9Da2FQSt6tZgSpJW
swt3MWgcYyEVK6trBKG3HTsYIm7qKSo5NnTFUYVktVv2nMCD5pgWE2ATfAzuVY1A
xOTONnrhsbrH4bfECgKFC384ppf0vpT0UfcoeG62Ac1MNNaW7ug/HVH7SrZIs+CC
bSwQpw7kYiZOrCKzn0r+WHrrzePECe+xiR6UMErliQMBIgjv0IbDGiSSQTGlDdof
wR/ThMnoWs3HVMvmczmZMkT3PDQCeaDxtZ68jPK89COCofuoYr8x0nbyWxTt/yLr
+Iyf37GuwnL/wH9iIVQzB3YAlXaDgqNNsFzt9CT5PVGCjHqVmqiStLucJvTf7RLS
9Z4slUIncubjSeRiwb2yVryrADIiMPCci7z01eiAdfxje+kYXVo8DoRINcHdPNCG
ha4LI/FSVTlcyw6wvHht6iG0hjvZ/RVO66M65zKvP+j7ECudpThh2lPTlQMnxGkR
BhyCZPU1Ghk6UKNWBxl9h/NEOXlE8WoscdWfb75pf4HlUAT+ARcjQWiRX2oDOT7M
jO7pR8C83xquL6Ufzrh04Vy3PJriYsSwc+gO0OMqAsoVQcUKUkGOrqHULR9/KRL/
3XB2g0zVF3c9NldLXqNWyWxjStQmNAplh7ZNr83yNaARwyYSXP1a6l6f8El2xoLH
vYTKsWSyZF9LFtNHMozeFMtOnHzhMbN+NmZHM4VAx6m9xpWTZY0yUKJBZn43uHLb
xyJTuQX+v6nCTDZwVqVmZuQOZKx5eyw1OXnh3moyzG/sVN4s7cc5AMgfh9Gl9a92
BccgolSAvlJvqN1w0gqJ3UoA2KbfpLMl8ZNGm0k64XlN+mgh7nutijiR1KHwwLwq
NNHDm0ct0ytmb6PQPe4fF7VCrMHOPm+ZDsWnbTmEjqOjgo8lmmPlKGtC2Fd6MtXM
VksGw40XpS3RI8FlSUjknBAT4m0VPWU4atvMliKWtSeVJhErhxQhA5u+ZdEuPgRt
W+jirKTzL+se3V3EZcA4n5Gcm5D9Yg3l0Glb0ccK3iaoV9p91448b4RvfmkUCTsZ
FABI4JWXVm356mXDYVzUUYFT3lC9qGCNIGQnPvuSNKif2rzip3r/gAmUZbnDWgCa
OpYm1kDIRuaYlftdyQBIbeY+gaMVPK1XtHQ/i6Y29p9hUxbVhkTXVjV6PJ6rpI4E
YcJvZ1W5fmQrBtw1riO2oPGYJICSi1hcZHGPxT1apEZsJRadpWtsJKaFRxsHi3O5
tac3ZnRnS0GFDKWUQuDk9YcFkif3p5QiIBt+hUiuurJ7YG6ZSuXMzKFHZ4hzDosN
dMx4SxoYTX3FJ+grcCFZC+6EXd1nf3jehKPe8TwN7SBKh52wH93J/uny8n0mnib4
ur60Dj5OKnpEXkI/2iv1GdIPrB96CYsDB9cSL1jgk1dyJ4spFNEm/ZleSDnudDKH
KOegLwXMsIv/K3DbSwfVCZyzAJkFDT8OBXEoeae+ssdjwR1Lfd9BFa5AxAQiaUnY
tsv20rD6kWPJzLM1a5LwSir5XBzKzO+py5QZiwrIdmdyTRRtK8BN+XN0M4pZra49
g7tZO/oRZSYBDO0VG0kno2c4BcLPmBHiX3y4AIKeIpMtKeayYX2bbFvrne/v3/+/
Wi8dceMrSKWOdt3dq9q1LJwbLwrP65re5s8STJJjZBM2jNpYkXOcmrjSSrqaQQ81
C6pLN2oZzBustAToQmrZNE0HCshxde3AMiMnlxNq4qqaDnrZXXb050hUkvnETVqI
tGVs5cAYP2rO2ZctYWiCsqrY9fhQvEfvbAMYu0nXMGGzKNLA+PTuPOSuRki1iXGF
TPzYh5Im72ogvCYmoPOAGGzoiVXA6Dsx9UG2Is8mFB0s+EHTT26yHsIFPmFOOyzj
HNvZIDsxcA4aGix+dXKpwikUNVbtebGCyFgoo99ZR6k+KVheO8lK4miGHfIz1hlE
h1o60uGt5hshu4pWwbrwBpq89X03BJwgx4360VavK4GzcOEYSmqUTO4exaT3CpHW
a8qb6hNSbIKZV4eeEVuVVYCmLosY36YzNQamRQCfRl3RseKWICK27IxvTbPIx7hD
YZWx2Eb49e8j5iUroUgGCfJBb1XVTSna8UtxKVvVhPbqg5irW1E95vvRtucolaXh
FJ1//ajII8HfiHkrx5P9DY8wTkLaABEyINdL9zBfogkL5dR0KzROhHLlscXStV4Z
QEzyKBXTe8I+X5ZIl9GVI9XApRuUWzVbqYcuyaZ/f6uI0fABsPxHHKNIFDnLHLyz
cZqKQdKDaNgyj0Y5sv3E1U+lVqbNxJsiboIQvcTSRral+dnPDFGvJiVxgl3akuNj
1F91L7iQgOa0QxyaFwnliMtVrWM2I66jSqx4uWlt9DhmHg44V3gjRQ7qjEGCgOy4
2fx3ar8dnZmpgGbw0go5latCmcvXfRUUEvT8LomXBr76dlvgQNpEg5+7o+JShYE/
mOHbukep1EzbYsE1zthkxXYpvNBnx2rbZN7XYfR1w5LS9mSiz7odRU3VvdIkWObN
wihcyOwKzRbHUFzBcLGZ4lWdwwjZw/sHc9+DZyxu1YUb/z8No7A37PkG6kdkwW2u
MrJyEl+KIkQdaHXt09Be8gKJ5u0S2jmJwuR5R4GQ+Li/zaW3fBe6/Q0KJhdtj32l
5/+eFvGOm6Z5ywx+JqzKKvz1P59g0qhU3CzB0PMp5SGT0bK8w9+iJfNDB3D64PSm
dmtdMKNCQjRK8yRtliV3+KjTYAuQH+yMZ9pDek9v6hmzOYFnm9CqCoG+uI9o0o97
8MP4NntwHCrL+fq2oj6Ie+MnnJYmSLj98FaWB7h/U0c63dz9fjVQpCkDv9KZv/Rr
n1DnJkzOVWe7y6Cupshl291vAvanMDFcMwOsbDYsjAEBZAR4b8T65GAW7kMZLfhx
k2AZjS0yieBia2Z6g42S8c/l50LgioG95EOxfMSOkK3z2W4cc6Ge4W0vqMhFEbU7
CY+aoBRiaEiNxp06tRhTsnnEFJqolw+mt+wWmpA9tXyY6/BWaR3bFn/xbALzrPSz
K44KUsOyjxzXZTJ0EKmDBEqBsyrKUQpOtAr4V7AN4tWAjKPXz/5KGZ2XKTHCFUli
jXIm6A/+5q77II29byvMAchpeH/RSAX2NdzLKgHBQ4BNC2VpRxDEKlmXMscXSbFm
LDM8e+XfpDIJW+B8a5apeeEhyWMM/87xdnCkiqXm21BzWv0QCu340RxCWmu/Pbqj
u54dZrNJqAmT7XaNE6AORae+qz8MO/3bXl7QDR3Yuz2n9hL6wkt1ZGOt6s7lrhzm
6laO0t8s6ULn4jggV+UC3JMjed+MJiQxSDYj6lTWRW8BRbunyhRq6X5E36dWwtFN
j3qsI9fJWX+MK4EXdratRl9Pw6oraQCzcKHJ9HkhfHKxt3mUM5a9DRgE9bqnH9jq
3a4lfq709XtWBLcoiclROWnnok4ITi3dON0B3+H+kDAZXpvPHwceYyu5we0BLrKC
9H8c0Q1aTcelVFbDu0lCdGcw5MSmFpjorU9tNUla73ph+PuRY9sJnZkMTiR77WJP
68QIkolMtQj8UcVaGiLXr0nOriNS5mbZYGEQPwTxkzfSCF94QGiuBi3VZanWoGEs
qy7szOeItuRGgR7EC7E7YsNAcNYHoVU0FTOL5oalfTAR2G47yGGqHzyO8HRDezTY
ctEcFjlHTqxnFwmtoH1xTd9IxeHoB+w277oCs/hl5tcflOUe8IsWK8RqqmXiUIeC
tykgyQ0dM11igBO6cFa0xma6nYzNqMlsZHYQG9uD3Yj7ouu66b6pEv/XFe/kSVzM
pjMszHdZRK2PNF32EFnCheLV2/YVE06kCUhu+UCzuhaqwzIxJjtRU4MjUYIBnPTZ
VecxP+bcIUVeiU7x3/Ekf5EfpQz9bWsHpKwreG96D6cu4C5Yd1JPzh00DW8204ro
6VxFfvlaFg2QHP1AWG+sYXJmEEd3xZ/ZEQrKJZNG9Ji0ds5Njv/JBDcSt25wV8ay
o7XOXnFKsK9hcVuky2ScpUSRevsUlYj/IZaluW3R1pgD0rKWWxCJWLJBfQ5AoLu5
KcTR+yoN8JTdyGOOMNRleWFUPLEF+upfbzWetx0blwfrS4BeyN/W9mtupt3lSBtD
mIFwM73NX4yVeiVAthNjmmbrjX90HnnvacxmjgiK8hglZfBtW06rsDOibWuqTG03
`protect END_PROTECTED
