`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5wPDpMqTnYtTX3d43HhYu6sgfUT0PKlIIHAMYm8i7LZJKL74tYxALcwGWeZQfj46
I8MSi+xNOkphc0XnkxgUfd3LFS/BhDDecRmQALomE4ZsiMlCezo3slia3xrl3Fkt
8bxE1hRdnApb8fh7itH69+OYKJ5+7tVBoIvukJj5DQ8jdijexsPsmDxiIKlFNUIK
`protect END_PROTECTED
