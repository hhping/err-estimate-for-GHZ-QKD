`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XqEsT4Pfp28zi8UGc/UPzdB+HPe5+8370ffKhwlOZES8+/iJchaDXZ6N432TJ9kp
Go1suSi32aR+gRUfkNJloLSiGZz4cq0QJ7HZr3iE+nM4pCy82aUDceLUBV495syP
qaMQ14QXsAW9ap+apkkWNwxooxT3xsbXBtSN7Cj8eYGFuV7jZ+cVGHLtfcf03kQV
/uLoK0v29PMcH3PoD2LBm9O3AIy7h7eKKRjrBBn+/RFjHaoyEC4953nIa5ZdEmcK
VSga4VbuSTmszMbXUGRB495s7UxR7egM5joZle7FBPrSwGfjw/8gdRTrRXs279md
5JXrf2V9XpXsacEpJYNLzhVmaCsGi3h2p6dywgPW6+wM7WXviyizcVtj65KmniPL
2P4ETrkKpo0+DvpADBommLYoYB25KY3LZcD0y2MCCR9hTCHmZ4VRtXwKqP7B+9lr
WzeCn2ZZowuJAPHlgkKEPJCFaPQAJWf1UvOoluSxerIV7/EQuqWyaOCL9LvJjvjJ
uFtt5Ei5rEpQxgOyP8N/QFK3Q7bVN6B6gxvnO7vNiZMG6wDDM3osvhpUmTsSsEre
IfzkOVHJGIKgh+BX8hMC2sw1KmCHMRKLOJWSvClBI8yaCdWqL4Tx8m80uMWRT/DA
A+wIn/v01jneBq/msYrlNMomjVxnm0XQdWzJgdf/i8jMghsrUBWQfg45f9YKzQ1H
PtrkOFwCVJRDBnp8SnB+ds3eNs0MEfy8RB2P+7zaIInXof3yvdQjULJY5GlWIiH2
qifTsKmFjmpPYNLwtQjeeIJ3EzvzvuZA+Hn5irfVHrnsWia9aP31r19OiGm0Awg3
xy4BlOfpNuPuuS+2bkaTMMQa+05PA/CXFe8Cg41fleM4XAQ0hczaZxKdrZyGeeTH
Q7WDCe3NfnwDRdaU/wenxed1KfBEpTy7oJwDV8Z/Of087gFWhySJFXTlq4ox5T+5
QoE91UKG7x9umtilQjqi2dCkebjTaEFXXsy1E7Rs/JcmjodlJFlGEwG0byjdH/BM
+JYsIcLe2bMnwSAt58ym+latndhuZovRuYQcmyqifIz4ezFv03PJoBIVALw1I27r
jVbsjvjBkyFsgYAfvJBErOuEYhX9tDqinueFTbOIzpnK7dYo3IhYVDS4HPkJHr3h
6RKM2iY4jKUmF52zQFuPlYBDIP9yAkgnoTNd2LXq1MoFAkUC+hgeAUkTU6GB/jc6
j8JQrXC94VS8vA1DVDoR9VSpDc+OPXJnlEZRLFf8Jy1rtDn02SwkVYpNBrx0bYT1
Dq3GrIPD4Zw4gIHBXNKm243bWjLzQqdkkDCmvxyq2iE3zwloNNnKCU0VUBNZGeJX
6qzQSFn7WcqGsu0PkJxnOqVPts/oHm5drs2zzC08/QO43oYPrZimEygyxqMQDFx1
GgM1rbrIQKqzAdDqj1qsbH8W4nmrnl1zgmAkt2HabVuf7+/TcKVvINQgbsbJNY1Z
o/HtgQRJShsBQsc7oKdGVdLXXp0NAa9xZ8Y91+a9uiIe8iYCnuc5MqfqAOsqA/v9
ePoGRTXijPhR+wzUkOzOziRYSe0EW+6knAwMQWYyTHssR6JjcktwMySlYp7twgsK
AJlML/RbGVxYx+6ASrZ7XEluf2E3RUpMrfoeqHXpzz2YDdd+7NtvksSFOw2BSXER
sYHYwuzA3qb0xwcrBD2hor3/U1uPzTL0fty9SbqbLNCGFuZFRig8TCCbD6hU+6jZ
D97y25wSOHKp5kwKNxR60rClo0JoTka0Y8Bd4Nbh5p3kxo1pCHYD8mvrM/RY4dlr
U75KVrtyLrtKisrgAjD0xZsCmnXEaINYX8gCOOswaqoRYeBIETwruvHYWNfVzkFV
7+JP3ajhwxR6QBs2u+oMFgzqjHTsvlkQ3hal9VJmUEttx/09rOdYHG+tlhu78Gyw
THo4Yx/RjHxIpPTfB8HjnkYMg4jME7EQWIYlS8TSBFwVSmv4TmIln18Hl2RvgSPp
A5YMRO5VgCxeoMO/LJ02KaqqQn5gpcDePmvdTBn89oHoJLcmzXqqu8HUCbAe+L8z
s8Bx4xJVEk4IKrF9vqcxmd9W8DSnwUlIDQrDDoku8TiSSsRQoWCuwYM3TCI9h2eN
`protect END_PROTECTED
