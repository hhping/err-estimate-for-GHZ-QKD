`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFrzR48Ccw3VrU4yWpvBpfb7Ln0bOyrcMd/9wJv3Jdcs1UlwrLd5HV6TWMP4g1Q9
RYQzEMMeiYuqy/zcBkSC9CwGUeWx+Ux3Zu3qOXN7/KNX4ssKGZNOsIgd9kiz00Ia
ym37jJyDi0MuGaYoCJ6PpsUck98e+g5d3Gw5Xhc/9I4OeQNcq0fLSsvnobCF2TAn
PSBB0S1xmM6MljYOD0ufLLyeZf7frgUDoUeHtFtRk5c5bP43+XFZdEZrrB85KcQ0
FaiJrXuZUF2a0N92M1+0wtpAHQf86KE2koIBtAuc49HVfKc5ayK0EkxqrBUsopH5
jBfQgHIDX5v+PzuqQlX4ib8823BmWcWsz+W0hlz8Ftn5v3OpAfqyr7feBXqRnKHa
SrS6g8bF53jw3E2lOX4B0QtMFN5ONcluqGauJ319osLHcACEOJlgvWcdOOZ3hCBU
AUFl49YT/6vbufkSc+h3ke2jBa4WZuFIJd8E5fiTrFvgfRWC3yJB0B8dz2zv2Q7c
SX0jLL10GOcveAgertHa/ijGuQECUVjprAjwJN9wXCFP0C/OZOrQK1ExdcYcjFka
rsELvNS5PZqcql6WNj3XnsmZJ3P69igBy1ya+KWRPXkfl6JwelD6FZ1LtbK8mrag
FG7rhau+mBTaRMP9zafm0zGVJQLxW2wbH1Gs+73mFabDNWR1niX4K+AY2/1ofLEL
V94AclvsTh4qPwr2h7JZMHDCjlq25Jc60nJshjxHyI8TIZBG9zDYp+IZ1e/cMpNl
RlOV3r5u4VOBgipJ6RksT/tlbvqkf7rz1/R4U9y7nbUt4irRWEQoG8GTf4/ypHCn
6E9ykf/xe/hHPGpHJYAwq4PJLftmaNItmt/WUBrrL1RXbJRQJu7FQP7+xycyYZOu
m2bRZ9ypuMxT4PPXh2QnaZELJcUHcv6UH6v+QU2nRQ2NUZDbeUb5E0knQEHEqXLv
wSgZCHap3Fk+pe2kwPiZhTndbWUZgE1M4vP59bR4r1vzbges7fIEMzSsXCNFgm7k
JSM+/QqRiMdqMPfzbIUR8R5G9W4ANulWUFmOEN2AOrYHejkPMTj9RC+Z3jQbEKrQ
rIexsALFqhzmm7uDuNJ5IL6cAUtAWG1mUqGv28mxR9hX5f9aH5WeyrZ9PKErPZaJ
EPCZf2/OlKtKy41uwLCtILlwYP19Bh14VUfjAozFu/Xbshx/WuJ5PcEIR1pwMCJV
Xkauw6Kxx9qkTZftqUFq2jbYxtpd0Ivj21O5mepBvEgFrLM5Fci5S5sDMLQA1Nz5
z+UVIDsCubAPzIobeWOn4GpFxK+rY/4Ern+M1wkfXuzwrdn9h2VS13AqpZyTS/r+
m9tFS7jMZEvSpW1gKay6no2dc7VxNJLoeTggD4k6jbXU+BXJInkH6cp4qHsQfi0j
SbX2td/uhGcMJ3Yg+NUF868RNdn9YdYvMTyHWPhGX4a7UVobV3lRAu9sey89oI1r
vLi+k1htt22MN03VPhuXMLCMBtvKCFGcNFbzwS+VBFMqQsi5jJ9uACjakCC1/113
DylaLAf9kH3jBcTFf7OlD/DaGnfxwUGcPx39gRfxjT/988+GeUiiilTf6F/0rYqB
glEKeZzc/99mbeE8/bv748bojfED6bFfkJ0bEvxx3EVTsRj5wj9d+bJxv3JeijjM
HT6MTwhC2JjGnPNfZE26RgAMlMSADdw2Wj9j7YaY3n2VeSwPtOs3MoyF/i0hJQTO
uRgOhM+qyzjfV/9NVJ/BOtgLQg8wwbg3oUQePe6vWzeaeLPTLQnexvRCM9v+po6I
TiQd72XvvR0LQxwcQ4Qh2EKpuwv4Jb6u8VDq9UbfZkg6W4Nvs6ZpP4u5NsCqKnvc
F8n9HM8WwhtZ4cJuTbqpn457EFnph+AM2F9k2kEj+o0mTwuawRpNqcsX0zqmg7vC
mUIzLDe+MRtuur9iIX3agVC7tfSpqARaefy237y9rWDVmHYXc69bgqwZf7jCXgS4
D+OWnMBwWTEZ6NvnguwlqUAWtMB6HBLYvw7J8Gnv4hjXvuQXa4a0oAaCC4OsyAis
DRzLkU2yq+Vag9+0L/l3zWGmwWpBiH8FG18mDv0bpScHtH86zy/mV9NwP8WOQr5Z
TWvmNIM08IEAmlDHg0BLpm34cIxl44i5zJX8tA6WJDJMDmpZuwoBBzsIg91KHo+T
WQDDvAHY8DFtNs5IDivbm25PF+5HpotHEDWVqq40uPiJHf6cXSOPaD64TstYvMSA
KIwBOlGQxiX/HFMdBHIABSnOsC24kvRcikxbobc9znAKGVzHjHzxnMFGF3tCOvTC
64U6hNcJhXDkNGaoRZv5kavhm+cc1H4qEvzF+vhujEreg9pDzT+PQtXpBD38LVTa
YRMCh2FuU+N2+9Hs6k14SNbKvbPEBgNMtdEyAb7Nl/UvfF/pvKYYAzxGhK3ylkL8
DF/Bj72tzwzP+np069pXCasfplBMy4gPae9LOQrQStH95SfrEDgRvYv6prOzPRZ1
tlwiEprcZ4UEY3LNr/ieqCr+pF/vKTHMroaH3s4uIPYk/rbu0OWkFCEFNZvN5GYj
YwuZqm+m1kT2Lgn6Dj+JP3Hpgl4kK2jrA1m9nhI5gB5WjhV20fzvFTRrvVNxyEHe
lKJ9E83cdDt/4rZGckNB70Ocye9h8KfnRG5USgxJamULMTARsrp+ou7AlFLhQ01h
f9Yb4KspFZYSU4+e78CTTlmQXxMqShGHakv17G/8eoaXUusDXT2ljpqfvrZZ9joI
5Er1uruieQsztpthNhpRYNbDbWh3k3V5fX5gJY+8p6c4y2rhu3d14DtB358AbG1N
Tbu3/A2E0NqGEd36iwm9cvK4Hd7J154OlebKChYtSebA52Ek5SOPUXOOp2llHmDj
Jhc6lir4UwEO+9vf4vSb/97XcAz1LYTS10wIzB0UdiCKNupIuPVALD/Pa8xcN5nb
HEYIPGHqE9xv8f/wPn6fYdf7d+HM64XL7xqsl5vHI0udruXae9/MAmgm9OkrL4aU
A6KoHZ8btBTeF1XVcGtOEVfH/Kz4lcMlqhncLQn7qQ1JJJeZYASqAfLEaH8oTnLF
sQN/3/NJM8s+PgmVGJ0cZiLYMT8rF9/1zDjIwzUQELoW+iWjqJhiLv2VGDx626xX
fCjIcsTDNbqKxSVvKAn4BGCkLX2pjdOsH4G/HXQnVsOymDK/pNFHzjZEN52/Mk3x
NdOL+eB31/rvR+vD5E71BhLYLYSaqKLCUMNYormV5OvelhoDgh/n9kg9lv1dhv3n
fFGRQqDTacGSpbDmeZhjv6e1iLaljBG3GjHyGyQge2CZTFZOg6QxRHCZQNqWiL4G
jF392Su4ZgqDfLAq4DksYfuhsn50s/zH3HcpvmsRKr8Oo6CCIhWocuf+lBJSGXe+
2MJAM7KcR2WZvXgp3JA5SyYXqh3DkQFW/U1PeindC1Z/JOvXhY9D5/v9VW/NsswL
jj8a59LMrrcIwNNIV57eP1YR0izHPkfuvG7oMtP5OfmWYhDduOL4nNsKdYhXhw5x
l5JLTnpo4GtZupJJIsGggEjW2L2uhHBXQgILMH4h8+gf6pCWgbkbEfkxyohrnUi6
`protect END_PROTECTED
