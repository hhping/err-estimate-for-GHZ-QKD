`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9uNHsCpAbd0gmN82jzyBujZujvL3/WNOGF0g7pWHlJ71Dlo1LI3Up/wPqi4j4YtK
UUD1DShk3NL0BbxF4ywTyRKEkQWICVSzPKjUvDapdThj5T8cJU2TxqhYp+O7HLHD
aqO1VyyeYTbB1PDRVoUDmXziM9/Gq71yMl3uZaAnSPXm6CTM+Ea0DHiDzDs30b2p
UAwy3Z3Mx2smXkj6dmcM6puOldjUeWUQ0SbzqdHa5DO0FJHveqqRuIOH4+ssG0R/
QKem7TAr9Us6QrsGUCxM6RFz1wcHabQ6pVo+q8G7WluUaYqTeDwWcgQyipg2moIs
+0skgeKZnBPHKQL4ppwHHJhot0t6ta07gALbM82db8YaUdTjLFdSfauId1oTS/Yu
XeBQAj3ebFkNkQgMLYdSi6wgd1Hu6yocrW5RsjW1qzkpCiRdGWY3OvlZfU3ymufX
yvTueaH+VxeLzDC6MRDO9ZwynmRHdTSBkN2T1Ehej615z/W/Ym0/40uAlcOHjUng
h/aQ/IwFcltkCwUPantQt9GAcSxBaOMUV4+YaUvtr2Gbs9J/QcMbEh03TWYgkv/P
3PaeqceeRtjND/RJhxAoUiPmUoSz2zSp4sFCvG0fK6ZMirRusH0gmgSkbpb343h4
0Xs51P9KmYetzZ0TUcVwQh8KnMeHYdMnlpn9H67Tk8biV5BY3ZpdY4RZj7dacyc/
5MyPdKTr0wspYSwJss/HJGNRFpC3gT/45S++pbiuWeMk7jB1h3bz99aalYp++2yQ
Xh8ChDgZNweVp15EfRZk55q6UNXdvwwyy2wMcZM3UFFuVS6TGtuX376Ue2h5xCHr
JiVjBCv/62VPa7PhwGYricfYQEyKWhYiy5flZAHKtBTgHEz7u/1wj6ALwLQnVgZe
3ZV57bMSuekn8HQyZMtEGpA6alf1//kzBEUZr9aI+dy3TJ1RF5AIRTV8XXiACmoZ
MwUYBUUXFBk2eZT92v0aTB9z3BQhAbCLZxZfnDf2BUD3Lrd/265GNWbUaoGsmnSU
fX1hq6f9NZLOmLN+cC7DJOEwHX5gkoCFlACETe5bXwZczeJZeoRDdmcpcx9vDm7T
LdIXkGayvvscAfOC/rFZdgk5reK9eAEC6Gex30M8g3jPg5jv4aly2pqrPmlOtzg7
ZKz1umMxmJalDQWmLTXC/zs5Dd6PQxXYEUgwGoMFbryr0ojGkfZI0xEdoJ5FXeTF
0FRHd5TeahaKWSoeUUstVvf4X8YGNEJfKWG5X4ARa3fXzQGaY33UQc/G0C9rzi4N
UoZ5leNQkdgJyNXoE2znqJ7C7gniAHPbfgdVyKqXnXd96LStz7nuhoep987wwddF
2PkZorqQx8t9PUetwCis0KGMBVOUf7gtwhoOh1+8TYWKgG3NdBVT/Cjt8oQZU+AP
HdCnMzVNpuE/ASAHHRLZyTX+5pIuiKqtqDSFUtGVAgllPBrGr3SF0u57ZlPdx4Ib
nxk1+FRAJMMmGC3qjlvYzizg3w10BdHzHQGEoZem6o7T+NPkQtcryv/18y+UCgU9
G5cVIBZMXoi5l8bXOXmKB2aix5HqiPXFV9X8cjBGoX3k+5pz8MeXlm8vnfktfPj7
ZU7I1e6UifQvF0rYjcYbob38dNmUxZU7FWn6QVyhO4mHAlY1A4vJF4OGgUGidaGd
VAxBE2Y1K2WoxoKG0FD7xppjfOrwsY6M2M3PqUWGi3qEDoqZFyWuSgu+40PVYgQg
3OMDYAjcmWT6ljC27bppaHE1IY6rW0ZfGC3GWVWOkCAHBEyLww2WnzpB8nxZZ+tO
+ZL06UUm0r+NfJMLhzmhf4EEkIRuIfGlhlZx0+wvIK6E8Jnxaq+nvyTGAGCrXriK
50Ue8YMBCdTKBI3pkkj36ahXcstW2oTqcmLVMKlM4AVEtowydFnH9SUQZ8nHsmVD
oCyRS+GZdMnnEO1t9jcFNopoD4/QuPl5AJvThEhhLy1qT3YZ97AtHNztC3Nbo5i4
EpUWQnQ9hzQ6F4y/ffnTYCajejoNjMVOmidvaL4JFwRuuifqNH2oXIYY11cvLXCd
SZPmDx1bSMFimd8pLjj2dO4CoLjuhjeR9jmWA6JrTquQPfrQlU171dI6SOZwa9FC
QD5U6gZeQw35Iwji5fi62H8f/ev4Dwoxe/0n+JcKStydPU5+7VyTW//9Lr/md7kD
cAZT1R4Xx74beg8c9X3qVOACaYHZOGGJ05nKKSrxmKnhP+qeoluWkZVN9zM69ObV
PeFqbsjyYVENSC4HWLWs3XpA+l+dbUVv7ZUBu2LL3xEtqefqWgyp9k2qjn852PmX
44zlw8ZLTaGSrxP2CxXEzU9FIo+7RU/QGFUzx7PfqEXkJoAFAW/2TCYnpHzUZ5aE
zFsnXuK8zRThhK55nb0F0s2q+13JBIwsQG4zhVwdInmGQSF3Z9rqduHiMlnx/siQ
P7fh6iORXmM7Es64cPQKNTcnx2D1SwU9ZIX5otjn0FD7VEMimC5sn1+R+HNwlQg3
4vd0UI4t/PHDmCwv0IE8Hehu9+OaJjC7Kbp5csaeaFtrLA3gpQGnujwthdD9lKB0
D1XXUvig6MdxOOcD4G+X17rjAaFmfzEkKfymSR8G/utTx6Jwae2erRc8SDka89nq
LHOtQdB5fVRD+AGAwRPpWTeHSY4qKedufI6OU0pwBxA2c4PCeB2ROJNsYm22I/LI
X1sGpRsOadkBRDMD2SetJHcYEBYRcJmUepzDEt/5ej5TepWKGT4UFT1uqOc5x2Md
tNVSRO4e//7YYhw8WoRmkU+5iwqv1N/KMom9jjQuluQRrWCdErnMwxVFXq9oFHb1
tmC3FxnTCgEInC7vtQUSMcq7V5M+X4b1ctCVBBsqdLmzKAVBkGdqKySDnJMOXffw
jhi80TVdNKxjOU6A6ZxSZZPDq8IpAVXiMceSLCJ/RGg/uGUQXFnWlBLLptIvFf13
kkMRZ/AgEh/gugynZzSBSXFrNZowFhKFPct1NISm5U54QwLMQTCBvCnLqKrmXZPO
IMCeenkNbKGuI2kdrv1mlM6HpyJcrymx1qB6f1AvyQTQHzfw/Y4jEZjdidli+pCx
0Np8N0Y/495iYKczGdBHngfTqWGcEBedJHcCv1I6RsrksFyROjDXM12nfGGRgq11
Ww3NKR7H12+yF4cc09h+9jfH1xj90mECFGcVGWEoM89elKKQb6lON0P5Q7mF2CmJ
Z5uD9XT8zJmeW0gO0xjW9hXW5SSWKsW3OuDzyP47I5uDWZ0kmb0qlqOXaMczJn2d
JX4wAWa9vctI2JfPZOpcYL9tAXpaJAG2iMD9kA6wczupwK4XCWl0z9I1QhlW/mCq
9d3WgxHDfCYSwY7Caqxhg3bRNxmvXTOX9wVWT/+3m/8V2TR+ZDcBo3mL9owRn56o
NSUmXzVA5GlyiHSFPsVsT9nJPjR0FWGKvb15q5pEnKWn9WI5FoZwjfORvKLnK+j4
XeKDlRU0A0GAIhpLImGOd81MjlWFl1B/qj06r4rtiPJTUPueb5x4tgUzYbaGfMLg
bgFHY7rJWMhhceYQcgDgzEJ3axC6dSyzFaaTG0OTusB+usRG9ePyXQi6NuSzkwZX
jNFjoghwRqjYQZT/LYP25nVPBCwN4cVXfgGOTthqiQmmHmd3gCqOWJm0YAmyesCU
QKQrhxL1eJigErn3yb6RDAVGPvWk7IWItbn/w/b7HZkRmvPlISWfSg9PBwaDfW/2
xgz5LxyWosuem8tJFLUJAaVhvny0aytZHO06ORwj7MAH7Xf6jQmZAlSBZUNmnuev
wBPro0Xw/yyZU7HE+psmXsGf3Fzv+OJidHpNUoeizn7QBl7D3chsZ5OMJRc9Kyd8
ha1ze6tsROfSGoNL0OxGtaZEj5aXAZ/4rAjjW58sYZhgmqWfKPiS3maOKFDqoZMB
QdSAVSAEeNLCW96klrpKY6XnU/AStSW1UBsC4b7BHAPvrL1NMHyexFI33qRojqR6
czUBvsSjXGawZeB58W48X+HYllb726/3YUfcK4KAzxmTasrrREzGFaC6tfz9EOz7
6bwSqz4mcXdF1Sw1+Fi4Ta65UYYeiwAMaV9TFUP+7P0SgN3eyoW5a3QmM+QPREDC
`protect END_PROTECTED
