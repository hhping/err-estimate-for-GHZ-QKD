`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXeuWqgUH+yF2Z3dUtXuZGyoSzuxVBir3djYt7wKQ4yTVZZMlxv9Gqfbqc8lrQgZ
7WFlWwN4bnGEvjRcvxMUFb6W2aXtzC5+WgQO9zXnCit0yY9bkRg4M9qNbzXqFAIb
JAxAMzMi6CX/U6TFyZ3qPMVN7SGfC1U0iYZrW8Q88kuFREGoTSHJbeoqe/HznOh1
oExmrTVYRAnyuqDKkRDlVauHAnV8c0YIVbOhmbW7aQ+MA5NDQ34JV/9KQs61ti4+
TvZ50qlBJCPqWVFpiKGPl90AUHt1GA1sw+Dc3KfAkQ2HJUAgYnDyPVKvscqzb998
5v51zYRhRnUMIA8TCVMzrgmFA05jry6AtbPpXaG8RqNbsqz+mxX/hzIrUu8yCGcH
fSo8Wxd7B50ekgiaFdUJ3WCBG5V1sS6UpZG7AFhhQdV6DWSMwcUeRMGcjU9r5afD
ohe+JZfcT2P4UBuTwmyuCoXA8uvUHI7kFNqtLPGZGdv+5ErU4NCaMB/Uaursi1PD
icJE3EMPhGY1s2csPq74ejXh1W0DSXaX+kf9CaQOf3sBMj5xRD56NHXN6giD9tVh
6gIX/5AzPcqUWBHha5KMt45vEr5630MWw9oxQb/dX8Hp4y221riDu0YOw3NwDvv2
jbELAOUk4XJtCzPU+mX8ERlfwlXat94ZlXfR5YGzP7cNbPcmhxWqXMMCaCzPaDTj
FJP7eQ51fWziI6Fm9+k+Iw==
`protect END_PROTECTED
