`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEXoFNUeY/fMvs3MGEAAxYbo23Mjh9nIbXLOMoJDWLNqFweD52aiyg7hzrVlHmPm
/590pXZh5qGN6dP70S2lmDE5XgoZQYn4XpQ4UZNUyRFiKOTYlUsyL7vSq8prI4qN
QF5L/QQkcVppijl75sxohQF3I2/BSIqToWz+POxhIEn7PCBkYzcVr5JrqZ6Kr0Gg
XrE/ohpO+o9vv+XRl1dAPKIQuWA2z2tJrBXS50IRYqv5jCLJj2uVZ/O1nKQRlrtC
hhv1owtyhXpbM0WD3/EdrMODwNqBJ0iGD9XgeatezlhA9a4vbnpGsg3w237BlwJ+
HPdXQ5cgDhgvw6hGczzKk+PxoiCBftW0tXiv5ZFjAhMeY7SKOlbx3gsdDv/r4XvT
6IwKmgSqu+mPbA3nrdqYY55HkfgfT9ZYk8Yv5ukc9C+B7xp65NzFc6DOTxwA7AKy
HxepTSMkwIanYace2oodCnRi8byBiJhsKFxDDjOFWC4CQwoM4AgBRdETueSa+SMk
zgqubN5DhGsvwiJZoAeMVBZUaaqPi3ZJItbDb53xoQZK0RRxQDMnpNCCCvNdtFDE
`protect END_PROTECTED
