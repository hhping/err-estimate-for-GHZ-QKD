`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8Y0XPfbhf7Cv+bJr4sSgnob6n7WiNcMKzApk//LYyD6kDo5JoNddmnQMC99JAef
phvALEIYSO7xyaWFvAIfdTFiO6GzsBDSokchXDeGQpMSwjMoejSkcMvr54PJph3y
WA2L0/xLdy4tMLYG9TrODo4DZdsZhxh9bsSie2CKHE9HpMExfx+xXhPqKVomxUBX
qashIJZOkK0No0QeAG2Ynwip/qMFF396mseivt9c5678ibDvupn+llBbjqRs8wNh
hWJ4c6kzTYiFDU7aWL4jzF143Wvii9fMBHXnsJwmexIewYFGyNtcaUxjOLtwfOlq
DM2COfgyPOq30F92UhKaU3Hu9hFIFW0kJv8++Y6CNVRE5u1nI8kBXFSYKtcquQ85
MxLTP+rrPSlHYTXat7RF9DrvrstZb3W5tYPWl1+ApD3GNIJ12ymGNy8iHVFtKomj
mZgJS+sVuslZjx0SD34AdI3orSN9mnZl1LpvT2zMrTULb81C5KK9BbjdqTGGsWdg
SMP+W5y069/BsoLvlnFZ7JbOK7L+T8fz+lNo1V4uQfye3ANbnVE++bRO3AbQvdsU
fy7RUW7kMGSVhfM2YHFu6ntca9nc49uUkXzKS+Sch5JhiXbVAUH4H6WyMXnz90Mr
Md7LLayZk5d5brNnbbWLJg==
`protect END_PROTECTED
