`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrDwz1uv2wfAa8250Htpll1gO5RtkrvYSY1BGP6cfBLD+Pb00MifSlv350FqM9mW
C81sRSN/5UcNr/bc7waBhyW45NWFlhcqZG0TSJ4ImRtfR2IWZaw+evJWasZyF2Dg
7S8iylUmNmmB3FEBDDSvDGfV+8WOnML7ORZ2krgt5t7o9XqP2Zk1RmUp4CI1+bz5
nkQyoyA0HgfhNMUvsAJV2xGNdET2hMIoLOwOMhhu8ZOAPQBZ0XlULzocozZiCTj2
2tR87FieJYzOdGJJXGedOf5fCs+AbLUzI/51IvEdKNw7akFLKQS5B/vL5Os0jEMu
JB7vfUWKLwz1PAt/kMSr/7TdVM3qA5mqsPaR5mpfrBaTJDky7zdnnG6ksHKNRCcL
CBU1KGHRDTcLy6Z98XVsibQSF16U8SnjtkJSq0vJPtb7VtwT6705binju5gkviKH
FhNtzrDQKTKa3W80BiQJ/LsQvl3fZkHUkgYdvxE+Voty4FkPiJojwhlnr0WgdCj5
NvbFUUfZkPglTW82m0/cSqzAvLNnVFSkyUVqHJTL6uBp9lN4zjQwzlwNQRfg2owf
vojo5BDfZHwDwzUrvdpc9rfyo851WTJ2NzmuSShDWh7Er75vw4/IjahbzTb7p1Db
D4Hlh3jOd7ombixydK/3pRwzzPVPPoLnGTfdsKxWMa+baJJDUjCEH5xNBwyP8H1i
dZKqTi+8QwEUVqreFuYZ1jBkNLiEuOrZIEUQCq5asYzlFoSBUuWikRuVr5TgG+CW
PGk4wL+zxjUJHiQOqH/hZ6pI9x9FSYuAS6NuQhrZfILnj2GmFcFWlE1eOsDQN0yz
8C0glCaYVQdNPyEe6yWP6iQqSkwfvRZBs5j9SYIjdbcEB5qcS6XltUpbViIooZeN
5lyKtwxXQQizTew0feRSuR5BdRRlspJ22TcShIa/6BhyhMiBfo0GCf1a+cGs00Pu
c9E1zuPFomzXQT0t9UG209z5VJ8omDXHJpKtXZ1mktvsqVCEeU1H1aMVhM9+Qw1I
IrPy+93c2v8jYMRk6UPdCR1kupF7lMqGZKLZX+F92X4YiDQ7f+cNFlIQxtJLRvhF
4RkPQEf71Dnx8XdR2w9Kq7Khk08S7K0TEPR4JmT1aDbOwPholvptHLkHbSq9wOJG
yZmNVKqSEr58e81joNDoe15oPMg2LZAnPcWIR4YJf61XjcKaNiXiol+FOOuetTTG
GdUXafjts3sni7vaAlTC/F/gus3tChQABcEm87SsvkJcfOixpUIe7V4Ry4omvs08
`protect END_PROTECTED
