`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A0z4uU6FCUfuwC+OzdgQxOyFNsoi1L+fNqhaUA+fUDlyBgQWWa8MIAugWG/k6yJS
99m0KndMnMCNFHsa6RDVDEhtePmT1dNqy1MVuzAZ8J4u4+wFP1Hl38cOroh/BaMm
7qQ5JDbWSwR8HgCtX+g5Bjya7l+4X8Ua6t/rFULSKPJOkE0chZ253E4yvXzkfAlP
lbzuvwCzLHS5OuY+WnacOh5Wj/OpKh3DcR5HaFfqWHWnXdZ8LGG67QQ6B5pevBP9
l+r8sWKYOiRleayoJWwyKiqehgL9cRnVwDC2nB+40i6xrTU602qKkGRfNSe0BV+j
Bc6O6ru5xJH/Pf5h2z+wo3FKz5KzAscFoz8BUopAhYwPm2JxFO/0Wle49SrqoFsY
3DBS7acmNbI1r/kYKpekXGIRPWn+Bb8jGJkBTUJ13mXwoHJxFv6cpYEzAqKY8nfK
HQe4KIXbDCC0wJjdmwzSySOnKLLwWTRjL+3pouzaB8tjR7VjHgQXgrl8n+QHKEyC
EZz9eUCabCF/nBwI8q2Bq5E7aJ0s150SBw5givaj3tCWKiDQOGjXUWTY6ikbVDD6
+mkcJB6muEHKk+C6ef8oV+lkzv2QjWdUoHtfgzSAmSLLTTCSdyTzlS7ebsKACo+v
iVou2WtBGPmDBnPin+cWjHez03qFf6OuFJW+6vjRwB2Ki9125EV0CfmVniOygqZE
M9qw/Kk6JRjRSTGmSj7ofc4B6yOgFtE0fU98VUMYhjMnliNcjGNNSXRZFsLIhFYp
IgbV70lw95sCyAisKl94brefZ52asPVcZw/Vr1kAPOm9ENnm6lEMlyyQHvv06zUf
oVLkIVMCwiLDquLM4R43AZFDgSIJ1GQP+N2D73MuBWlP6LfFHem/vD9GK5oTpIcV
w3KcH6F2+CBDvFM9zgXWukLKc22xQ45x7vzmPaoSqjqEEBrzYl80UP1M5NQsfSvc
QkMKaStSlHsn1u8LMNnoM5vwMyVrtv6jzl0hNLUjhhudefT2JWsnRSVPteLe1+4f
8qlzRBAIa0UJ2DRQkrYHQSt1R8C2Zi9u1DcSU/wCSxz9u0LJy4H1Dn6G0o93+Tm4
nW03zGr7IhA6CvDruLqZf8q3/0Sd7AeEA1x93jZ5aomZUBT2ENn8yNm7a95AFc3+
+4/quKZ4hij/IY1gIK/oQHWuuxSLABAfMQQhFdXI4nrPE/W/GO274+F6uz+capGi
sd53XGCYWnz70SDZ+DpW/TbFqHWevnfEwtB1gQQVrMSYYkvT1Xl1r1bMn5OWvE7i
GLEg5fAXAXsRQnT4FYnzf3c3or6RooGLuMpxFozSvJ6IeoR8QzCSm+UuEL0Awmj+
oHh+8IFxOtqXTdH7lPzOI4d0+3+9Suc4xNkwl9agnyTolwbnp4qt5Lys1UByKshi
RyxyrMVi67B2hTVc2Z/I0/N2gLY8Vc9A7QQnQcq75Gwcjy9rl++c1ukcMQ3zkm1+
YAo4LfZe0qi8UXsYcL3Qcg==
`protect END_PROTECTED
