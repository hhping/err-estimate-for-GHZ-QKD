`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqugBMIPuXYLHVZmmFmcyxHvXIjQZgTxOi51rSPBRQnhVcK3se+CLJnqkYlRuvf2
t80lLZkv6phq9YDUhS5/dwsuWkKw1PsU1n0gzUbArLAKXsxIRZwzwAa3j9vKy1gq
YFyIvYuy+ZuBv2AHnX1qm+chDkYNao/G6azD+P62NeDI60SJ+V+AWUXOGXTzEchu
H0mtOiC46WlMluACWq6k31NLLJSYs9fPeShlEB8geOESTZTjvH+ng+8e700EJmY9
a+oAKj7CuIsZx/12onu7BTyefmG4NXJ2mfQ9Zj9srnhjkia/o4SkPUC+yOj8s5ow
nyORaZ0q56gEuWe/7+7FyLCZn/FNLxEAKJsSHjemYBeDGDfcfwNBzcDEbzKmleJg
hhP3nkje7sB53cO7lw+0PtHwAnX5VOtNV19vGP19lAjHZziB86l7CACNwC9HTiHH
+3MhRTTPn2lEcM/LT4kR4xca1bwTmAEaG3TRE9glfzKsofeandVcMX/NzgqhJiVb
fCTDr0raa2T9hh9NWiNZJanu30LzI3F7pc+Zgh0FsYl+kW0GbcglkdWTv+aOv2/Z
sP5yJ3CWBqmH9zzJM3Sdc32SmVOTLefsfsKux40ho3GIf/BFxs3p7kAxdPS+BEs1
dzwn3dHkjg5EX41Y75+Gb7GIwXu6m0BwI7RRTbWm4RvPX7hsEjAqA1FUqZHKaav4
t1tdGfSZNBVD49LQZun0hoFbd9n2NplNcuIcNWeSR8Yvu+e84jGanNQF0uIj6VHG
Y9Yf5EKQDT85xEtKIwMj0fC7OR+xS7CSWqtGOmomoVgJ3i7QNC5qmyhhktf7u5dr
OAe3l2gIiIudsrxH83nAe3q0hOEsuG75Rfql6ZVUAx8GeE3JltB8Zf6aKbctzRC5
tKW6TQ8UReN5BrssZ+q/I43enLlY8Cw7Ccm2jn2cGG1gYqnTvuofnXo4QQeBfcCP
FQ0s+qAbqF+8amMpij4Qu4U+9dqbjaTc/tqFbP7JmLh6GZ2QLwF8uXROauSEJwl4
kDO79q6bFD9R7yU+CTbqCmEqVzZvxmjW9AXdVw/x7XgIHOmUMoZm/hjTrMeabdAY
G1uC/GLijA3ttz4aizVanjMHXfwn2Zeb7QoLbn86SSRYbdfoCTyn0/Cva93O4iYs
fHrrSQ7EVGWOf2GH1LqJKNFFx+WSDX4bXLYddaaNTvYLLztLryngmvRQqtYzm0ke
LYf6eTrTbKqkPKWOlaHshYrKbx3yLs/0ibLi2OIWy04cW/ljEs9BhC1Ug9m0w1K/
wQyWcubA+lKU0IOnppwUYgDUNB/b/ORPDGleFMCMBkvh3h0zh1NGY6d7QeHqNHSV
Ov9AnLuyz3oogaSOnbYJA/9pK3V/sgjKynUUIVLxmd3ycIlh8ITaBndiQ3SJHfIL
bPteFftwV3WPa9iKVA5+0VuY235zOts2YVJ/QuUJKJN1/HKoqrz8xAdJ4Z8KN3Tc
PORMqwhALJbGZ9SZudTYpiukp+pEJTC4+Wz17kf+AzlMeWgQrTGm/l9eC9uXE5Wb
0Si1DT3MKfRFXAQA4YcF4tGrVmtomUTppdC5plrbiz9agtercYWnKP/5w3VT6GIl
q0vPI/OAUY1c9d0EgVylKmlUsVv/UCREzGD6nsB0xWoXtzaVyPFFFsj332dIuR/0
XeBTLt/E/FI7JvWxleDgZzeqHJOntu9tA0eLRHrUZG8=
`protect END_PROTECTED
