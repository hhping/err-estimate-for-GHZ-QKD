`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbbqjEVJrizTGHZEAqIKuO5R8eQOyMtAHPU6jeXbLSywiYKw7FCvcqwbhCKS5uVm
rTvslZuOE/KWJ4b6F73b+7l2ygnwA+a0Iqr7+k77/+jIgLgIooobP1EPnUEWHUKt
s5v1CrtirJcM9vTOoLYIMuEHdOiul9Zygs6UYqU1Z9v2UpwBlIThKx7kNxZLNuFy
8PIzzdIS+bEEIpGcI7zf6MxzOVNC8Ov5LVBAQPT6gew0JhlrqfUKZECvtY0FUMus
5dw5s3lj7yobj4sPTLbwjKkMOR9C+XQLD3c+ARzXOD1EiE2QTuTfBhmgp0NavB4B
QiHncJGt/VlLI9ugQdP8lygiP3iqkpidZWvQb+BJ8aAjCLBfN9hnglZoW2Gi0qJX
OWlVgH1sCCJlH4VdYurjTThAQ2etnuV/1SpUZU4JV2jnhAqZ1uFIN1PyctLfkcpG
qPHS26jeo4kI6ga2Aqqgdurad+R7uoV3A8dBiy7S40Po1RwB5/fJN2zcJF3BG0Gs
ZjnIJp4lAX62YWhIQLdPldXSjv7cZK2pqoUcXkybxgobmIlylmPwiFGoJHqUO5zs
lnFU1KX3zn0QL/DXTrfH8hEgHho6EIySCgX1Kh3HPHV/5JIFfpZ1fj268eEPLrhG
eycNFN535Ll+WitxqHF0JlT1Pz7cKUN7NJI36c0b6DUPR5fdi+W2kIMdHJZFX3dQ
NG84v1htibIjD0jYdw6+KEDNAHPG9Y5icvQeVweM919NPEelqt1OP7hdZ1eOMfsa
ddAz6KodDkKf7v1PT9yUM/hXGuNo1o5NMmGEnR5RnqRJfv1CsbBP8dY1HsIFr/e3
e7ey0f68PfcVWcjE/xKReMddWUDrlMm+FvoEZzz0zgWZOiaFdcIS1gBxMUy2vB3U
R8tqDR+DmpDC94zug8jBTryl3q1IollmemVNM3GNys1lRqZoppNhzrK9MTofUiYl
qa5WAkUqo4MoULuKpRJf+L/TKNWIcX5PaHi4l5+pHM6BRw+TdorcK/ix+xQT0Adr
HOgEOo1dxZ77WFtFmIzleIC/QshCrTiKGGo8n1WWJ1mLf05QdkEMVgqhBspd8kRO
gjXTzVZ/tZQnIICJfe397mtSc7D7MQcfC5XuFgG2eqh61vJOtQvMtoQPE3WczHyk
1u3qh3t5C/HhQiupBBbUbQ0nf0u9n0b5a9++X9NmWYwvyrfFFzniygAuBq86YsqY
As8JY5S4FHiZ21KuBnfMA5amY7V/3flksfc0CAgqweUu2+Ll8VoZS/L5nMfpQMCk
RHnGeDcUwFDzYNYS0zfZruXQSJxiVtg0Rq4idePNVOrP8D5+VOvVCBTGXYx44ufN
yu8SCpIpuaoVrwr0WDMun/XtKynr4jEoZ7rCZvC57ykMxvxBLAOwRadnFPxsJkZW
6s4VonKQgC3yZh12ruJspHpbFTIjFzu2i661ieQefvtybSPqlY2kEgHP+6CkUYng
2fMW4NI43JvJ9g86NQSj9ZD5143s1DJmrbTvAbxOie6JdnfA2rG1ZVXpDg8MWKYV
MWVPf/9oeptr2Lv/hmDUUVCTODlGAFByHSxo7ktcG/kLBpp++p/1pG9mV5KIUGzq
4WVl06tM6Pz45rRBI9j03bRwWbGUhaBacLT5If0iB371ArqVCqbKn53kUyM08w2C
EBAp2UGpeP7zT41GANaXfB14Ed1NKrKCuFzMfP3ZFqX/hHMKloN5ipJ4CISXgC2n
oEVBQilnCjWFYkHfYZwmcdWDEcbtAYzfEnNSQ3lWcD1BgKGDfL3NbHdl+Dfb0jIL
cMxa+bFr/IhBP4DQA8pdoBHosJfTd4I3OffbKA3AF+RTUgA2/Q42Atq4/3OhOP+m
Kqc+AqnY23VKFKCxOIdo4SGleKbNm9ZheCR3ad0xSqcLhkqDxHYWh/PxnSe00KZU
`protect END_PROTECTED
