`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kK8VGxmjCUcUNx4aK2DwsC0c2B2TSVk7hPucyMoS6NpALii3H7S/uyqkT+JZIF0I
f1HhNxTqOZhGSQgzRSUZMXKRGmUInT2/Rf5RykGktLeEoJg6HPUpJ8iTWtozz/wf
hMFVYR7xpV/FPLuDJHsEpdQrNw1DIWJVGeMrxKq6/kKT+UO7fWPZkLICbNSqG2AV
d66z2IpIRezq5WtcucnhUDcSpQ+HSXwVhIGgiXDC2xAvhu9anKfH0OtFhGqTtFUs
xt1wctxppiudwFxkD3iNMTpV2DGLuivuCqduR3ZTvG23IdtnVwVnBU7YHq8Bv+xd
EitWSMRgkaPIQI34tSCFCJHIyMn1wTuQjSE9+csa5v5UN2CMMS4rUG11zBxIQZ1B
Z+qUUHgzyp3dxEXcL/33BNO3Ja1RogsmgDUD+j4wZaQY9N9n2uHxGq2klyHdfubx
p3BEBMncayuftiR8SQT0mlcNjuMQo/FhpiMZnHaBLdMMjXmG39qSdrs96U0DcXpA
Kd17Jw9Bh/j+n9LSEavnuj5XS+8WLpqEGOcgmRQGFrFH0M1VP1vWEdImIFxTaJS1
ltznzjUl/lrzvQaJZm3dEq/rsHW9gCPWSFEE5Hrc/bKcz/CiFvuLZgRAO2Yao9Fi
sugu+S/1nHDFfu3rf+jQY2a/oaqjkh9mi1nNKuq6yVNDcP/wQ5/4hCD6xIETMtxR
c8R3hhntRG44ZiiFnHbCX4JFjifkZsmUE3EIgLeE83jHtaZa74oGSeZX3G87VdPx
j0OoEiJslAQL3gwfWRAe8YQv20WiPu2dEPvd/WUmE1Kd2elDYPpjGQTQyTEY5Q6v
poI5sYewj7C83eUQ6kYOBQwM46hXi0w+i6GmFnX7X1UArTCJMkJVIbNNhFEt9/SU
m9kdKLA5eAg9SPaLnhi8VDrBmr0UHZ4v2L0IIx+T7h01NxMDZz1b1lrTb+ZoXjd8
mrEk8pVlcPrrJ1dlyOiwID1WDno+ySZaX7qKGa1CC1seffA/PUPJhAkStknOADur
xpDwlhRw+q5p9hw+1f4EyQ==
`protect END_PROTECTED
