`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/wvWxOyekjojsZCBGlkt9tXa3gwbItH7nG9gfZd/AnvTydzbCLaYrMMICpHz/eW
9QeFCjomDTNxWY9LIx6KoXwVfdT7iMjtiNiIZl6a2hDHgO7qT0Kbb6s05OTfmqiH
1UeLYNPkmkILgRxkR9nPogm1ic3RmfXeVZBdn7tuMCf85pJHEyoPEe8v8kl+gY2u
nTrkCT+4pwOL77yOQCVYpzXXebVKpLHYBbOo/VphDOkBRR/CK/TmXS9aOlwFl2vu
IbY6v1pxiTR8j0dgrNnvfDrpHVYKGXW0vXlydc6usMIdH3GbhkzvyNyVrVLgWc1J
UteXu3xnhLPXslyOHuZ8JBjk/VH92HNb9qVifN+LEAUguAoF7KvF9TA/WE+KeMFf
QE0RzPACiR+2xam1VTeLedaWuoJlzRsE7TjffpvrWPS4G3TRsz+Ig1Nh+zZdMRbo
qIY/+HCE5IkLRkP7xXodTcc1LPZNoOPfDwD7lMsH/Hd9HTWF6C5bT3fpWnt78U1L
bTf0X0slrQ8Rw0qeZLJtyg/8UdY5Or1nmRAk5q8ArNMshxt+QOeKQZxuXUVgexeC
x709iRgjmGYuyuTeoMdfkYGPXoieyQayJqd27Mer2QTCWPTo09WXIUK3p53IQVEY
VcghaaMqMXlacePVc+P0vf5QSYyFS8hrPegMgjO5+nAuN2mrJgkYdp5Q4aJX5eoy
pvXEQtno0cHYPgJpZpJrvn4vvAMhEiBKFLaNNXDriaHhxShrOHQvkDuHCGQ5f4l/
PQVTIOTqRG37V+pBr8nREArUP8+Lh10rEvhIqhrJSiozSC7re+oMti9LIrFj6+Pp
ZrnN2Vo2MTMzoAPboj+fLVX4HfnlD4ogUyPnVmxHhDRuootGGF5v/RGXl1QMfx7/
Qj3m/WXGjBbL55968hKLd9qRGxCs4xNtcbOsUTVWCScUyeAk4rdS07pOCln8nAgB
tJtlybqEaCHdRGAoGY7yKZ19piHpZ9nzSc1SHcnFfGZZmEc3uz8PYXNPAWcNmtVM
opdEWtsag/UvHmJdpdpsJe8xTb0UlfYgqK1CRt3uEvYA3M6PREiieaocOat7NbNz
7WBGkbqpJoehv7BWut1j7YTpa8eRDssWZzE2Kvdsfgc=
`protect END_PROTECTED
