`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bY54tWszKw01YUWJouEq3U38LqeGhPHwNJz35OiaDRqQv8261o9JWYUnOq82JPLa
23qJpYLHKiuf5mXY+OLx1r0WBzM2CE3bOuQfkLU0iHNAsnZl0JWmRKE3G2zKf+/6
3BN/uqtvYUpzF4SPXJR+wBfKCNkI4q4nueTFsNeEtJNhPuqb6OuieTuwavDwjhSj
1jVi0qPe2slKuQDJPHqD2vE/ST2VXevIRfqcZ1Umtd2ZIbHBKC5kcQnCbGUuOtB4
4A1qkgpnDGCczh01wy6yerTHZDZFH/Xwwkko19svJbAUtrmbJYryC28HHNVZEzJ5
oFKW0LIFSf24S8JfEGgHKfsex6ZR/86YlHblKl76F3FFsF9h4U0Foc8ohuPuIPRH
8q/q93Qaz345/Uiz/Prejw4WAz8xXLDhPvfUW9BXn+c5QDHxHWAtBVKB2QgIRdoH
+JOsp7W8vP2/frFbCvvyYziiJX0G+gLPfnwVNMZ0QuTxN4XduUcyTWpXlielmrMf
fH6/ciig1OiA1bnWaIcnWjgzrSaRzHFN1Bt0kL05Vf7dXU4aV0KrLwb5iTJ3fDV2
H81rWmUbMnovi78/nrQcDBxgOaZtD0UgJIVVF+11zhbtU3tKxcVarbiTssP0/w+m
`protect END_PROTECTED
