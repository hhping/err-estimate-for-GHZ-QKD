`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrTzndc1u0/o/VmZyscfYe0s8v+YPV//MTKMmoh1g0ENm2tOUUWeICAks4lm1cU1
gYl5tbCyR5LUu015wRSiJNPFsUtfJVofB2CEuFSjfn0Lz7wS/lh8hnhyAkkLXyUQ
vKFL1WocdR7uRbE8W2ZQpYdS/oNqsvMYC5QmiE0mj7RlOxZlGRsc4feeOZ4xAkGq
AA0qeQKJddFrHm2HZg1eoE/IFNYF+G9oyZtyRLbYfP3DlTpYUeI5WH9Sn4LIdG5b
/iZCYDaji1bx7DqU6SRLnoeses41OuxwtFaGMiqLee+vMecpqo3SU0fUrL0WxO92
yx/shSnBIVp04ZxUEQlhFkBqWXXfMxEJ2Wp+yaI9rD4SGDD/5oCw7aEfvif6zRf6
bYIJni6UEYOb9rMw6HD13L8zqmKS3ZX9bEnQQFjE8jvdOTon0aasVh2M/4ttWbpd
ILOts2hdTJLVeYVmbmh2IU4F/Z5TVI9AWU7WA0vOqxVAYsMVQzdVOEE5EMfjswYK
WaIikYkn6f0KcgBtelDGzXhg8JPApBYSaK2lTnmNGVD2ieDRuQ3n+GnHPLKa3WiQ
NbgRl7O2yl02e3F4gkfTUvZoE2bvEXof2A6ZvKEkscMwgwhuCD4E7JN82QH1XIuA
jRD5MKSBDJ1UOtIznNOPk20JYDx/wB3SxM3AEfAvbZXKDZklagGt3nh+QWLAkoq8
K2Nf1neGRQYDttBx/Bvajvd5BXaIT1eBUurKefIjKfgDhPM2VsKMVlgFcWXY65ij
EOMvOgMNH9NcnNXTL3k7tKI6gBsT8Ib2mysKBivHScyoiKTiWzzbfYvY7jlvceKo
U8DL3PoS/m0CderFF8IcqdkJhMr1nmdHhJ4n9W++JRi1eBgSQc4bZSw2shxRb/mj
huWR3iGxE8TRw++guJEtoytn3cVUS10XB7VbdTTxAzq70ZR6UyYfxdo+1WPnk2hP
OWgR02Lsc7Pt3JYDmP18ZcA3ZaJAFrUhWJHW5AGUc8wlbKLB52H5nKneUxNFSBKn
tYMHMjCBnh7bjjgY1mvwVFBmk/Cej4dptvmJaXI3a6l3aUvHn+5Pxn1fjiTf+HDR
ZlL5UpgQv8kJ8KZcCGLeU1wnfhmtlV/GQ8x+UsO7pjJbuVhNFV/5a5fMbdKDKKDq
EuuT1BP+VGEhtuXffGOCcQ==
`protect END_PROTECTED
