`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQpAKJFGoVx3BjEw976rR2fW/ZOnV2ltO7rx/Quz72GO3WDd80x6AE76+82DGvLA
de0AuZOa/K5mqK12rFqXIdXznXsAu9maNhH999qJUkTJoJ+FF7ZskHt+Lpur5eKC
gbW4VYCqOq1CzMIa5D5jrivsry4HXwanJyEELqS0nXPGZBOW6T0bqr4sXAqhfhaJ
jOV0naitF5V77JYT/Xv8Omyst8kUWtr1T7byHFVyJ7jwO8yjrf9FxOoOnUd7LKpb
kVfpBZfiWbZFNqf2uTBXrnDnVqxGWVXEWwWreugh8OTyJTHzpK/k3VwAg4ixeftb
HynSAyRR10vY2CqqzDFmEG4i02JAMOYqVOnoTmICeMeihh+TPQGA0zMlSRI17C3N
aqhcrJySEEbAaETNQGcLj0f56O3ZiYd5I+/45tZbzc3eQTGZ81xf1MkGlNBp2g24
Xv6OjQgUc7MWCJectTcAICblzm9Oxh5qRe8epKmiL0KLIWwq78+ImL3NUAo6wX3d
Fa6wF0hQUTRKIEwZjssCyc9KyCQL/7luJEM41Tp8JJchcSV3yxgjDN4IkLVNVLGU
RjA4156wgSc5lapt5dvrfxJzJfeZ8jjBh8uFZAH98Pr434/ATuBYrhs0EJ7FHRPB
AeltJaJYtnfB83pjk8RNkyqNKLWm9E252mOpsn/RKbOqthqKhn4WP1YhbqgQiKzP
ZQ5NvN7B7L1Wnno65o0+HmYdSddYDoOvHLimhXTBSX7O2ZkIxblzAigl/nw84h78
YNN5k+4JcNku6ZM5sj6yCA==
`protect END_PROTECTED
