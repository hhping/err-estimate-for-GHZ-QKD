`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n37cRCNHGrqZ4RYr2taASnaXoVlrnhHyAVHNZFwQ3cJafiOqwgUrrfTtPfQlPF6M
3HlrIcnhlf2emw/ViL6sLWuUaCacPPzILDoLeNXcZTLAvEFbY6uF1aQPFjtND9kk
rqaAVZEM4/iYfMiIo/yDkxZ8qOxxu0P3ERZKCOjzwo5OfljbibD6W7zY+4LhzD9O
QZjnOh1n+NXq7QlUjrusQ4Gc2hPklxIJzL6hcjyd678BTSLEalvlq97IITasynhu
W+o9dTZlQy54c4bhjF+1nUke8VSAB+lLEm+jLr6d0DnUmFWVJEZQEIRVu23sFuBZ
wHlKOmRKAZXg65+euaa2WmjzAgw7c21CSWyKvalkOcaejDtLNtpEHjtbIdVO4kMx
yjAP9Y4PvNwqSaSBny1q06nf/bq3ZwAM+eiBP04S0hA3s0QhccGceVn+bDHkpi1o
RAv4amNazVFkS6W+o78lHvAGA+Api3O+H2eUAwfmjyBz+dx4Vv97yvhIuuaG8LV4
H5FjjM+uF67krCyAnLpNZmDJwvdUoz+N9wX6PvyEwKbFczi3XQAInRaN7NeJOg4e
SR+kigbwAt8IvgNwX8+5IJW6tl7gihuI1HVU6ouXTUVOlpOyikELmjFijrcpJZXB
fxFmyuZSniG2v3pqsbqT/UM1vgZnZ1EWa/3ZSl+MoP/2AAa3m5r43i7Zi1uU00qN
tUP1xRs1sWAPNovPEWVkf6TUEzlfAltGtQAMSWFMFi9I5UrW9RlmKComLS/u52JE
EHd/A3WCIbdRGDSHiqffx0094OshJA9RsxBS3YNwS/pmMpc0+32FvQTJlYPBB59Y
Jk0XIF5EGPVBWgdeYyC22c2S9tKskVUfOntEvglIWnmLw+R2S2vb5sXMBUSHWGmc
DdmrNjbyB5MfqlzqnuKJHnNP4Fm0Y4Lk8rjbggvmGGjbKZCyCdQnQGTmlJ6K06tw
DHfO9eJGoTHc1xIhqGIpccpkM5pMn1Fw89uhJW9iIN7c7ePcUcKOKuaYA6SCYsuw
4bAiW3ghVbupSjonowVE3tP3ul+vIKByILFdY6dI//4IOstV8QIaeT/CFHrS39pH
oW0H4VCMU47Vut5+sKWLX+eeHfwUA1gZhGNAo/rfunFhjOM4ipHy7+wDbFifLphA
/p+l+tr6De6g5eib7Kc/CCpe3pjEHt/LbH+693d4nqg5W/PRMH12C/VzeFQSDWPd
hrbUmBT/fcIvC7N//8aQ/tAjC0O9EyyzGXpE9VsOdblYfyYJFjUo+oQmaCS3n5gW
`protect END_PROTECTED
