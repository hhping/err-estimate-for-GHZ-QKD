`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQZwoI/1ghMQ3TQnlo/lWgyoxuTxlOLG95rVQbsfjhBOD18f4B18MLIslIgWotob
AADdSPR2waT28EX/1TjhqhmhN+A1alW48UN18vyIOX+Ypif4AGV0wPJwkT82is5t
+6LGIlJN8pMwgY0puW16H8NJhiP/vsrgbb+TF35ERIxsyf032kyQNiOT4Q7LEQrE
hwZouEhPOyN27z6B7bnbAdW/9s9sHsN8vCfxxkSZdJp5r9mOVv/Cf1hQwbh6zR25
I/PfNBe4vkqbrRBYnqJyRkHTc2NnaWl6XbC4KBvaPOpuDo5TMJnwGVCCnbfUOUcv
jgfj3u4rMMXDomR29gWkVgzpoG3lQmAxHDzNWsWt9sVbr7y/HgNO1EhkDpXnwE+A
srhIJX0J4PQK/ZGqG8Zsf90gsqQJv9+8LFqPJBNAZH8OcjqR3/CF1eBIAxyibBMn
kLZtpT622FRnJyuCEDRAHn95uu0mZv/IVlNWnoMuBggJYDceHTOLMZQuCSxp/IJc
vMQbUAyIpqrdlz77JP71H22ZhtRP+5HPDJ1A16kCtj8DfU9ap5CUaJXpCwzRxp37
EZ2SiEGKKo3k37o/+juJUDb/mlPL9LRS0XiAmAYp3l1EM3vSeOvxtCc8EqcyCobA
XsAwxs7scCuBfuiETKAaKDRVd8AqZhh/p6s1ZzszzuYQ8bfcMPdiVl4qD/5Ml0CU
pDHQxjbnrYTI2p36VhW4GzsipSAFyBF7pVe7lNjABNwyVZkOm9dcK/iObpJOxpqH
0HeX2+eX2le79YiU2R/SXDExVCRiLyAh80HDTz/maNGuBh7WUP1Aeu3uBNsZvjSy
iYVXACXudh1KIj90zOqF2ySou1c54ChON7iGSEv6BC9C1DhJuU8mZC1a7FzjeOkj
+lUOscgwzhD0dudC4cRH1X93kxgB2E+vQUQt5r/OnGTAWMC9q4dgWktT2QLiy0eA
U9guvbeseutEkfsGDNQyjj4xllRfxr6YlZrEhdf+AEuqD/B0771yU6kiGd82U9OG
SnLiwBE8T5FfAOUE741kqMCHjWWG9b+Pc6Qi4s2j0M0sMTSpR3FoR3qF/n2w8rIE
kFxp+gnrbGpX1Lz1LJgBsF29hx46hQh2+ap03pO3+A0IJfAxI0pJr+I8rGXGOIDy
3mF1Pembu0KiPA5lbtkt+DET9TTq12l6gsT3TR2/H1b7bNOZs/88opPtUGhq58Vm
S0gLAhOaTVMc+KNa8yqFrZdLucLM4lMCKMN+4xXOrIKwxwWV/J6tZwJXZPfruKcR
pOhBZwvRwe8hrQhhmhLUzSLFQ7CLZxHuUcsExKmU2YmV7VXydCFpUZ6o0auWz2S3
P3L+r3+Y0lboHjqRns+PctfKDa0VkUXnmKtOXpj8DciLY5IYQfodU6nTkN3Pv4NK
nDk0RgbAEJBA7yTlo4V/L5siiu1urI0c6usGWR0mZTMP6bdzBXVJ21X4bIAcMce6
tF6FtDWTEMeXWAKslAj1bFC9qv05RRfWu0+C6Xj3S14MJNC8DQj91J+VA6UnwWKf
sLZhFC71MDiCsmkgOG3+Od/8kroL3y9Gz/wAzm1SBvEsyXgo7lYifDGAGcSj3aDH
x8chMolGBnwE0rtgW2QmzkjoJGyu9ct+kiI5C3UcPNr9tHS5YCtq7460sNlOP4v3
B3U6Z0io3gFT5cKtF/QhtaAq7JPIi5xNq2sa3Osgl+s1TOKcrMSZGfHZN/YxA23V
5QDN9Hyn2bqoGJbWxQwMVjZdZPZ26C2w98pNprUOZ3Aw/nMnw9giFG9baDpTjqwM
26PiswEefR+MnriwvvabxKLhV1KLax4OMtZBq8ogV7n21QOzE1rRXKSdt1XhORKr
S9Sgjm/ruWMVA+wy/fnuWj2yIKJAxjtIeiJgIgK5GAHZ+u7regJscxGhhuzAA1rj
gCNRL/B/zrAkW7BOJp/GP5UOycLl219/1LPdFeOdCkzVkGWa/k4bKz4F0Gp6CqOq
2VlFDeJsF9ztGcDix5u0ce4qJ5L4SjnvOH+w4UKSGczcal8HYK/mQQK3pgTlpLHx
SpSEq0+6WmEtS152jjGCz4sNguhlnP+a6MkHTPgNnZPXd61mYuxFVHZXUe5r0HZe
jW7Rl5J+MaaDeV19PsTx2b+DFIM5WxytukFqd0++0tOil2D5EFmeeLswDns4VWUi
p4o8WQo2Dqs9Y8tsD5Q8nYx3EgtNdFP9S1/fIet3jj8vSK9tlFBiOlLOflgXBzkR
hZPNR4zLCXuHcsc8Gn7s0zLzOwfFhUSpbIDL2U3770z0+sKF1d0zhdeMdexP553u
iyu3s5Yg34mfI5bC+GP9y+7oXAyiIFi502dHsurbLptZlU8jTBylbbzimlRZRBA6
3R2jcN1+uspVkygh5kiV/lPH5WneBkNry9RH1Cd6GvVuADTTW4ipBXF7KuKk5ww6
6RpFm7yRpQtqqL3RmEQEU0T48YsF5b8gMVKqn1/SGMQ2ADG9fn9M+d4qZhW8wTYH
A5RlMx8EV1PyJslpqU63eCwyNZtbJ16bHQtMR3Hp+JRvv1ymG7iVm9C1uxbgOGhv
iwae7/hOej2ESi5BPH2Dyw/qA6ct4kGcpUOhryb64VvEOaBNndteVpfWSS+M9Ewm
z2NBhImyu66cY3LSrBrxXXp1ypc+xZNOo+8IkFehbZUorqUrUztMhPTdDnQ13P8+
LIYv2Y7bADvmnScrvXaiodyUL2GXiBdi6w40KBPkVprL0Ahv2dw8RaiXntFYPuzl
bioG4JOIJycvk8ii34QUNJSM0UhAFUemEp/tm9rRtyFdSxKdAJG+yIP+D8itPZOE
IMXHncVDJPGK1CNRnYuSTigwlJ6IOW2dVwThR4IWnYaXOc8UGMFZVjqEDpW/Mgnz
YLryArZKCFbLh9AxNO56sg==
`protect END_PROTECTED
