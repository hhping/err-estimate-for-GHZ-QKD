`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XyEoH70u8UwfidiKTeRbSGepQeTMX+bfkY+ORF0cAyeLy8FZd6lUl2G8fYqos7d+
P7iEVp6E3ZyChvRJgR6BvabKttYGgO+Vxq5MC8OCGWb1rJiaYcCZXWJn00iqB1ZG
YpSTVDSJAUA3/LPqzPZA0EMHE6FWdJX+An17KflG6UZCiyyrtLJxthGRmp1ehECq
6FNh2bsX5s5XPJnoaEOZbHwRgbE8iAHDHMnn0ZwhhYaTdd+iKgRT3umZLp4yy0+E
8UCBtOd3xSGz6+A5HVttCl0pBiLVHO3nnkfrlXq8VEcq6q7mLHE9JN+RCArgB3Ed
8IRh5RvgOvS9yQC3iGZSHvGBnHXD3M8mV9KfwV8K1FRp0hJEWY6G+qNzE//7WTzb
4BKjyzolRN7YdRPpnqT7o/uNJphDjnyUFmYFHJlFp3s0FSBXCI1IMWiDVZICaGaf
TXnTQ3GCa8ahIGIetgzsA6VaIJuF6cpq/J7D8931cmTGfJG1hG0gV1t3ZeY2LxPx
Z55gIDpRcF+MQYOZJ/3fLjxpeLwQFr4CecBLiEwAWKjFmy01Xxi86Pjllo+hXKuJ
Rs4m6B44vQ3eTe13FTyOXf+04Np4XqQvUBohZYOCjst03PTd7kW19BznM5xcc50R
`protect END_PROTECTED
