`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICOlzz77vf/7rL4rZWGz4Sh5mlH+EwPKEVus26DoFzlFm/zive5IYxVw+K+HqFhw
W1LjaJTNLPI3LDV6UU5yBw7THJHdBjjuvWPs6KXNwpJgcqtc5UA6o+6qRsAZGy4l
RsTJJRZ18JVrf9xm9oIpDo3bBqRIBtV1m+aAjqnHCtumDhIJO/GiwYhf0McntVN0
gKO45cZjQ2QI+ls7bxcwb9V11P/+kTXNrOiqMiaoQ+LGNX05i5c9vQEMymqhMO1E
8xBJcSnYNFwIbmRxz8tdr66gODS7+/T7jdXikWAEASwR59obzOMzc6kynIsABwIE
vaLmQ5O0k8qxw4W4QpUnjW+Wb2gcr732QwToQkfhpBEc7uw3swnpZuEpEQR4vFiR
qluIUbSNPXAyMglpFm8WehNGERSqW8l5cJB+yFNWizJvyEOvWxglNh6ZfkiVgusR
NMe6Cl+ZySFBdQETsYRavJHYayYFqs8p1mNE8uF04Hm+1Ye3/YegVFI/z0tapO5Y
qeR2GpzhaNCim7S9sHW+4O42gTylsbm33kMgjMqvO+omFPY/GnKdQDv8fX8+/Dn/
ZsApStFZplAkhMxEj0vCunftLsOBKT9jDinnbMhzHYTo+jQqnicKAoQlXrFWbxTs
`protect END_PROTECTED
