`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSfw1yKG7PN/+unsmxvnP3b0klzppqzE/OOdP6tbD4dKo4jjoU2036MUzOUc1xGs
k1T/rE/HGNPT1SrI7RngKQ6W+RmqHhoye0+cOUyZtamJg7lbac+vHI7yXoWW7o2Y
kCUzP1kQqPsjaHHmLquWM2iQgwoGD+thywTo0Zkovgnp45o0MM7SjI+tXke4oUUA
5ntErpGdzWJsTnPOMcpL+hDFgT6FpHSD84bkcFF6GjmlWFpr17Y6G49km/b7kYbE
CuKvFaLqGS0Q4yOAnXClmbZvg8W3op4nEiC75dG+vOnHSGWUXb3on5+0hggUgf9P
st70LAI5Dbm0OpL4BEpk1QqqizdaLEwlapZfVR1XlErsWSPq8rk50JHlgjeKWusr
Vjg38UvvlYsJmJiYmzuFwVUUVN4ZvhZLWz35uKNxApPskd23HEuhHWKnz1FtY4g5
SAGmtq5WCKMGHX6hLE7QW8GxCB/slkilVjrSWJ+jltXQ3HnuuzUrDwX4jJBJyNpg
I5HtPI0iJPSwHFf63RKGQMc+bA6cKegUkhvoGSf31LJSu3VjIYl4e9f6TI6AZs3U
i/Ja0iM4jXeFdH1rynMMlw06OHtJZgfTs8Z39cl8JK24AE8vIVSXaD1GjX9vaNNH
wBQcCJjfeUF1oj7i1cxf1f9WpjPiZ5hWOWK1v48i52dKRj9eEWCLXzazUjWx9WA4
OPJH3yUqaTN7NVA6D15WE7frP5xTh86O/0z2Qi9Ym0Gc0eN4CTu2/Mb2bqHX14GT
nJPyaG1sb5xhOSvHUez3JVo1ZRvmKR1kbELE0sIgmDhmxyZvAB4NK0kqwOViHgM7
6h2Wl2Tf85mKfuELEnl2A/LM/f4C4Kf6hhghj23ls5+bd2Nt36j0l0U/WpwtRRCl
RwyVat4Vv1nRd5txsR78s5GMU36cSHVUDTNUlBO78xneBAKyCL7VUemClbYVAA8Q
q0m+jYfv5g1LnnsPXDcXyOIfBZUh5KPtGzlAlkBnHTED98q+wbLRl0ZyhxtnT7yj
/VXuSaOlZ26fbaPrFJfIlTH9dHrDWT5TUEcQIm9j8L6EIb+v6ST8DnGhnqn5uPY3
PUatdxFcXXlh5TUkiGHtPkMz+GNtYjrsn1axZHpBq4CTfkIj8TOVcXFXeMa6/eC0
nXOs9NPWBuYpWnd2jiGn/iNiiIQBtsO49lsyiefeQ4ljw3TC6ZhRbX+C/rIT9rij
7NE444ldIwsOzRfhC3/tHC1v78Di+e5uuQ/0AL4ItlRB1/HpBkeMrU0B4EkqIkJQ
AJm9g+PeRKkBMEZbC64q4Wrhsdwy1TlKSeNNnyTTe3r8wG7fyH/OPq63hJzo4jlB
NWGChAw+WZ6vGLGJhzanzT0QO3lK2py0ROCCbxQ8aiRHEMEMq+b2+aMD4UEhkfAM
n+0eG9kJgTrHWBJbnyEdJ+sGn4exvNfvo/ltaseVrSxprcp6taD9qKejsik4T7zU
pdZQKAB3bTUiLWeSM6APNm+3e9hbaka+mboqWzYV9+zE6MB2PHRDxQwm1mY3gpek
VeUdXMvECV1GF3EW+iLExzksSGxnYvIF7rB+lyA/dflPmRIEPsK4bSRtroeRkFnu
+Xb0Ql73rFUa08EhINJpGAEBWMvRIB0amsq+mgDA6ftzlRiiiw2hv9hdcTGaqqzB
vA1F4D+ntIFXbpQfrPuah+YGuHmniV5oj2YYu6ufOdReci3WS2IFO16tZ2xetaSf
b1eyUNFsioqSNJTzwgltDszo5jzKgzfYI7OD0dyoOkW6Aj/8805wvdMbHuN59tZm
orarwgSPFJ5YdZYutJX2XtUDNbQNof8D+ytEUJZUfI+CmAD19KjV9S5bo6LC7bHe
t/FkIx4VoDEqgQ/DDVRCyiNwCFyNlEpp1eW7rRzh9Xx7aYwGWXjeMt9MbpcdGIOm
hY9s5w//SQOPKx/eV6xK3l6mrFTglYIi1ZHFvXtr+bFfDNmpaZC1VwHMynlKTCRh
uYzmqVeDA1pznNxGVqX3XBZmaN+Da/wjPZuXvLxE8CNa2ZcgMfpn9uJLHVYZn63x
4b5pXoGS9yWhNknanlMK4558sRT0Mp/G13bOlfCXiH7B86Ta4Z4IbLswTckcqMJA
p4fluCS/xTNqPxQDE0ltToWCjbYu03m94wJAjwN12ZpD9h5KwCSS8BxkXxEcvsyB
mnK9oE5lPWbyMSxVmWMp+k1BHEuKZdhXzmNV3Nf2HS3EOCIhhTbNvC0lxEuZ97pe
hWrCbQM2eOYd80YQNMyiarQ2iFT5DbzYBnPIJ03RDFvkyr/SxnnCDrIGYtFxxYWn
DyeiClkgTDv+dWTWwFhdwREkAXhbvkgHmRgql0BOCOY00EPonX22OksVq5lBRVR4
IlZrQw+Uv/J8LczdmSJSumP+zAZhSm3BKQjjL0k+pDKlLdS09dM1B/5rI+Db7+Zm
3Hxo77nE3fJThNJ4z82JweZdoXjCtBivufl5tS1KLpvirE3hS9QojJ/Bbc51t2XF
KpIe6lbXPUzx24D8nm9++b0nWoUWlL+uE8kmNH/b35VDn/2ewCkKE3NjqY87hnm4
8Y6maMlIAiX5AlUjMM5pmFZlNdI3HOv2hErNtqj4/xzvK1mtFnIN4yalZQALN06d
28j3xUfrKAaMVIZ8oNqgjaTnrrtewbWGRmgHxh6eVg7wgA1ThVKL9qRB3fbSGr0z
A2cC+wYJRAhtKYfWMz1Yq+Kz6T/LqpEuXhEExJSM36BtomoU4yGgHcwHbq6O1HkS
XvC4FPIvuvN4hRqhjFwpLFCmxGiRrjCisgkH/uhvD1F5cD6gqzIKBoZAuteFCVqM
TYGV6OL8D1nsapHhsaRL48un/j4WOK4VKMOgQ7LdmREF4UAcjwBkNnCzppW7xmfZ
rZwfmgWb8q3/G1p655lZgvLQAvw36FC1CcPMCHxNZJjrgX/SzxUA/19nRSU28Te9
AXE2GFWV6fjLgkDuMAm16dGCFB9pelfIxNwQ8U4HMmRl37e7HkOUeXwZ6nX9iBvE
3JeDQhDasRaOOI+F2Yft0UFgl/3+ZWEXIxugQF7U7ahIgjEfaOmveB1oeMaDuXcw
gh/ntXpohnbG7D8iC9487uqxU9+DUfE9VQ7pg0/JDJ3XXf34Ss+ehpMHi2oI/HZV
oHQRBtBfSAEzVWrrn4fg3vMOrwd8kVMIDFUhCM9Md11kGsyfXqo/L/zJhP+8WEt2
6M7e7ZqbEXBe8/leOmUlbALczLyDK5x2WAdrA1k9fK9SWepkR9DiT8Dksl6QI7MC
qXO+Qtdw5OJwTItZriP18jJ3ScdUZ0E3hCh26K1CuEta+J9ZgvCxNRGbQ5Ivp8in
tvkH6qbRJpGNsQIRsSKZr/6emTaF62z2CGFwgQ2uuogFFkko8J54oQ1acRjzbLzI
mrbdIQDhCtj2A/3uAUEBkcJW4sj/vBNV04GDS6G4NjBgx3fS0oP15NOR8aEg3GEv
Uqx1kz9FYEuwu46nDzeTqzEYbGL1xqFCnzG6QH0gWdaqgm/qm75GxGSZkCfXzslq
uFoFoTR35cm9v5q2dWu9nTa0OjsqiRIlVklSvhtWdJdu0Z5A2On3kIAhf8R6dKhW
n5QBfN3Nw8DKQpBT+3V2yVa4WOt9euW8yGiSFpufPUPz1vaQeUnANzZ2vPJOzODC
8F9l/fvYdi4F67q2xBu+xWSQtY4X8apUIbIDt+crwBHUJwCO79un4SSsHfRm7o8i
8PbrljcS05XqnJBI6bvjxXmHZCPXoHRKoGjaHHylyd8+Bbv8duztA0S7anTafPEN
BiNxPc9BuiL/ML6pGxgZ5lp367FAysdyVySz2RQkHC9qaomuAfAEwAqKKKtin1Kv
ERPtdM1R66XayDpHVNya+pjeYpe67102RWsczWb+rQSSEpsRAk7ZouMkvoQOhTiH
jVBllhgBO4SuJSz7GVs7T9u+tFTdZzWrKF42br17eAHMzNIzxj/nc6E/7rwKcJu/
2nwP6ie9TD2h7Eyycg5xG7DZtd0FgKK8s0Vd7IQ+2J5EczquEuSwhVOK24JFHZxU
1Asyf47NZFvNXAfEBwgywCLNjzjoCiYUIDWW3PnGaT2dIncLFSO9p7A9cvB/5CrJ
vSN4s9aaZl+WXTDMMDxOdlTpeNgIdLziOPFFRGlu8UQCjf0YEmARNLyIrj2DEnk5
2z6ij5kV47BVYa9yiV8jP+omYqGlZhHSJmSwzZkUxJFXzEEtgQfeoosS8ouhqVdr
vQSl42rxz1izS3b1gS15EO1sVN3vc2592ib8Mtx6eDtN/hCkOFsmkPHAU+2Rk8DX
wjvmc5Q0fN427M2CkdE54lMTyQR5mLHTJS4jsokXG5IVmZNfYyU4Tq0lo+Pm3BKw
Mzbmd7V50ZaL5I+KffLd/trsLyN7Hqu8Ku8V2dfNir4QaTFSIHJnuxnGeAQoqMKX
6tRll8yA/1kSs4wrhSRZPPIhAHWjhSLvo6qZlMho6nuU3Xkb0DvVUpynLsVSvCjz
y92wO9jpN8oESAW7nFkQAEzzq3b1qB0l86lGWJ/Nys917hVrfyPbwFXkbIhDVfSB
HQVWW178ikR60Xh42FFvbXalkY1nwKieBKMx67iX1VxJ/dWNjKHZDpFFwNrZImDJ
RaBIbPjdIaIxIi2aPDdRnf65wLsNdYm4U0nvOgIZiWu0VDodyGfs2Y26I80t4mBA
bcCMQf6AahPaxlQ9KKHOPHY3hfURaOK0yiOCz7xeBwUkVVqDKapxutKDruyWs92Z
NDi2qCt9HcbPN4eXEes7DJdKX1UPjdmifxuGY50bc7Ggy96CWmBtnedsB/dpammo
6eeewhCyynonLepOaMhjLSxwD5DjRGf9XjNEl0RyO99eCptgNeBQZChPjRaM+aPF
zWTCh04gibVn3HdpyvPvFt+mh/EnN2JcfgP0Vr6JFgO56g+RnUdIXBQEkPYPybDG
YGbBU6m4warnr4iMORJuQkQcUm2PT2CJydCWwopU5Ttkra5MFQJ2YwK7XSlHI69n
8c13cqHJi5G7HDKeUeveQvy8Wazi/xW1pGpyx+4+MT/JSWfKsPSknMzZNp7TaRvB
NNgWDcgxSrJONVoa9zmu0NCpWjlPPJAhKBdVh8qCLwSg+xJMFlh5n8sUMfrnAa1d
b4/41nVlahYKbrj624FtpbSRefoCDnaeD/5wZ9bqOlIwJgfXsa/qBI89z0FuTD/b
`protect END_PROTECTED
