`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSlj+5LfmpffkD+hG1guEq7i17/Jx7ICmn3mxFYUnDcHHBBkY+HwTbwsdzwfa9zk
7Yxj2xSc5o4/TYvV2hlPqp7eDV5BVp2QBVoXh3PJq5o0Q/9GZCwUZ77GstyLPxeD
TN3x21b87E4kB395E0bPjb8kZft/FFYlFVlI/1tqDp2CFq+0UOYEGhLOjMa8/vFN
ZE5MRWIeV0nq9rJUMgQRkHnhF8B2ndm3KhwpTnIJ9zpdQuaMp3dHFZ/W9qNPofuX
hrn5d5TVf4+vuTbvd0VxyVASY14C8aPBwnfnxeZQC3hG8rwkUmBlFEL4kBiLLwTN
eZZJY3Od198Xf/3Q+8eyVZWd8VTGn70wW2gnlny4I0MVqQB0J0tN+/tGv3bG3McI
gAj9EdXrpEHhqYju+ifDJCh0ndLZNn6sQ6jRpGIgSyvZI/gsg2EgQDVte8kCwZLn
NSs70B5GTkGRG5NWafH7EF8osTxHNG9JAV2ZoJDSOZkQMWmjqV01mKsgrZ/tn6uD
zZTAcqn69Y8vBmvyuEbIrByjhA2j9UeifyRpcK9dytXVIgTDnLmNzDr1RoZ1xxvi
LeQnKrbcCfpTmE5jOv6suKkHPGwKTuENf0ycv/2MCGS/iNuAcn0FRAxYzNHzXce+
KNP139dxMn8/9Iq+DoHkBvOPmCKzBFN7Iewlqg3i2Aexp9LJBeZkwjxKpLAMWQbe
ddlPNxPt30BtrWw2TV2kTptGkRTU2rSw6sFc/WD1S1ftKf1dFtXTaUMNy4YAiO3x
0fMRrT+L9DR5t9GyYdchFClhCG4fugAeJHF1yyiA0o2bUiTHtRj8BrY8uWW7bmXY
160UDJKyRlddeEciRqJRVsTA8rryjxzMjfzv+RrPlJ6nghfrYhCrQcG3Y601Nkup
GV/aFH1YituR07wd60OBHiCgKMnIWy3ocnHRKiga8ZiOw97LxDna0NTW8rKR+5BZ
kKCI6DmoqF9+fJ/NNpVzmqsOq1SzUA11a7d4SeIfn+M=
`protect END_PROTECTED
