`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rflxA2HfYWKrcmbX50lYr1TgW2N7LoDHfgUe1PpSSzNMJnt0htiTiEG4R9kdjLFk
6Q17ydyL7Z3laGu720frrVH8MA2fWZpY84AwJ+PhwqxEEw8H+fHUmrFNMEoS+XoZ
Pz+XqXRn3U2kTyVeoDHPx2iQG3Hjnyg5Z3UlUSLZQ2qQxqwbnGddqQwU0+cUFKeg
LAHH5Re9OfnIDVPLB4TVhoLWzTHtzP/qqzqpyvTjMLHeDCPVDeLz4iJdPlBtY6mc
8T8/PtyaKCbTCBtZm5nJHELIRXIylHGO8P9HO4SlvMOsluyyoA4Uv2KFZZbgFXuK
NQgnouX5BaTu1AAnp5jZ1ETa3mZZye77f4OTwhIWaVq9FJUjnHgW/ZfAB1h5NYF0
pjfxm4DfipFzMWngkZHW6igjlsfLGFhutEpWGUvoMEwGLlA5FcXR1bb3tUc5m4jK
3YhBJHs47HZ6p3m3i67yPrQQJp8KX3PgL3rBkvefumnN5cwaEAsVoZNbbyfddrRx
hMgEQxd1ZoTHSSoH/274wcMjXRxpXUUabkIKfIaoHWfgq5+2x9s5C34cMIqNHVqT
NGlfvDbtWqEfAtn1KOLps7ELTbkKFBBB4iNOyRce93hfsA1Xwj0ZZDxv5/Ewqtdj
wg4QeKEGag9BAyIQKr9DcBE3t4CrFKB5wPxY9v5P7JEomOKlEPUYa6ryCQACCInu
K3kE1U6uvTJwMXjwbqtuBkQKEv/Mf8fnfBrT6XNK+NHa1EyYOEkUVEMRE6Zr57Uh
g1dK2JKHAniKuJW7tjWk44OSiwqOjBIu001nRGEjmWwkfGp4wplD2zr4WVgmtcWx
OsJYdYsU2vEwoov7JEwxH/DHcyM6KFgwG+f1I05PEUyaOl/qOi2jzzEUpJA2fQya
rMjXGDO9AHKoV3YyVxp4KeitiXlRY1MiH467g+9BKxkBATe6FekE2Y/6umKgfXzo
pWb+P+XSLWNsZ1U5jI1B76vR/UDtIMDenhxtHuKrqoMvIJGHNla9UYsiVk8eYV2H
3iGDwxmY3PVv+bpXCz9X3BTUn63IIfZpjVdF7md+d7JrzZ14p0btfAjFUZkZ/bVp
4BXFpEsYQnCJcrKs5J03i4ZWrqqSgZxVE9KLePU74j/6aGhDl7E/79/27CKlRMc5
zRHKiUXHn6idVxOf3JzGofafjWvh37uNxBXw0YIQwt3O/iBJ+D5RIBECtQ88E3Ra
wIBA0EEPh2JbMRBnZeSbTAbBd+uYRGTFgggG0ZNrX+6SLeT9wQS7IAuJStGNO8xU
by69B6x85khs7AbacVvjUQYxnmjszxwa6e7E0Y8NVVk=
`protect END_PROTECTED
