`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XS9fxxH5AnkdMcl6JQ/qkw9PN8gcelsvW2LvC86YfGymyzsBec2blRK4xSRXivlY
/V7JZoKs1M09gSMX6wvKliHfzlSN3CpZ5qCH3MZOItulILAMiin1Eg6554/THDkt
2OBlS90rGazVQhVRW9QfvcdfF8f9+KJaR+26W8ePvygZ8YGSRpdp3InIP8+/ycp8
p3RrGLUCtGD1u9rhSi93vzst/wdvpJQud6thLaXqMm9aBoCYErsrZgQr5aJAOYT0
TUfCOidWSYVzYrQoMzqG9mFgMehrOi014UkO/F9u8sGUyJHBswqW71wqpPuB99Uo
BiKD5XSVkTiR6cf4e1Yfy3qDETQqJ9HP9a27fXGOqyoKqYbxl3+AK4VDAHlSuVKP
zSh6pr42qB0HFWldhLQ2xIDx3qf7/5SvXUkfhj7UKss22CLsinHPgsuAmCl17pIK
QxmO9rIkAMivl9F192fbJ84riJSulnfSyiqpGC/mrw3gX1rbYcEtqNrs4D1YcNJI
7Zgz6g5zEy9EwRk4YvKDMSs9jnaq6vtcxhHZdqDzm6z1RomDrWuo7uXtnrQno8CC
Qm3XzbESe1mMjF/fefKB/ONr2X9Yvox+xrWDj3oWQ1NDWqV7kjkYgMvK1KueuN3+
qFsonJKytahn/Sp/0v4XiZ2noPnj1hPJdmDVNwi2YxN9KDPyxSGXUs+go1Cqh04n
+nqm7zfdqfYsnj/4VTlCGu0FzyKjnGJbENsUKsHXCa4LJ/NiuAzyWOf1mf119+8E
`protect END_PROTECTED
