`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+rjKUI/CgDfKXwlBArcl9QTr4MLDFqgoTWRyuCKQRYGJtgIrrlzrxzjEIV0pdbB
pcrkuLeeM2ZIeJomUgmDNhiS6iChv3RFVrbkDCG00IQxV/qP+prNHNUkKYMl8Gek
5zXksziZ642ZGMSqJmhPvq7AZ7mAPY04kDB24tHYGql4HJqqW+sNicBAP2s7Cwf1
UgjosBqb7c9BDaubN9gD+5KzTp92LLEcaUVaq1Ztxzp0U+s+F+p5PhlOxGoSofXW
hDA6h7O8lRhY4MwDGtuPaSo8h+U9MILrXcJBnZor9tazbu/j0x7rkE/DkRlQ3Vbi
61qI6gNewLJ50hOnmDvj2GE7ML4+YLvOwPYHz6DyQHFOV6JIqYI90xhCezcnN7O9
Wj3T77UyN+17kt1iVJYuSE+J7kk6kV58tBm8cQhx2ybul+avuHIYEnA67HCTIF+Y
8D2vBJM6ANbBmZ24+i0rlahPIPPst3EDYAOfkPuKYNanBgXuu2zhTnLamAEUuXb0
QdTqMOHby4oHrZksxhACSniTxQ7tcrT+0PIrlpEIAW+VUoOu7O2PnW42YWFmsr8P
a6zV2aERBwugncAIuPHHFw0olCBqEnAHthfcX1+taTNXFDilzJeDELaXQkP546pI
yEWgR7wpf6XwXogSoXFWd7tuDzAjmElTIWeKAWHQ3Avlu9T3bEHA9CYUr6RWEPqw
K7zD1ImwFd0oiU2yvdDNOhzejLEvt1zcDdESCKkJPEU+gbGVfuuv+kLzmazfr2Zf
R0mlNtJMn3n3brVHiFFbR/rnri08q4LJOSNg9ekXC1EBpwohioZTduKQ1CT/pE9A
3TH/qIHX9mhKF5tcHL0R2/2FXBjFgZEH/0EepJryvxYjysNN0oIhtC/zgd2J/zJK
8AgnbhzxOKdX33onn5H9cbd5dgZkUZijjH7jvfVz36/mYazbXebIRCGfh9RP05YJ
3bjcERHy4u8mB9mAGgujq8uzeDzY5/BhIxmV7Z5k0ZQcHfTpjlsT+j51xI8IsboP
qW7qwqvV/mw3ZGn7tXQl6mgVij+k2neho1Tc7Ft74EBv/fRPI/Ch8C8LqN7fx8ek
RQgwy+r4VoaIMQkwYRkMmd8QEZeTdLtnw0ZTH7qbRiuEGdIMMSj+tuNyPYAyEmYD
cYItVd9xNQpCRtv4GjpYqTbdE0G9BnXP+3zbV5E2Kt+gUglqdUWfPxBEQ4MyQFoP
6l7Lc8vVyYNehcNV0hp9RZrpRFhJR+7zmT95qz75Jv9/MorEzudzWJFR1OtSy5Yz
Yr79/Sq2m7Jwq7Kr/2mULQ==
`protect END_PROTECTED
