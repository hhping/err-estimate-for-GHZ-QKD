`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cd2nsURAlNMP0qlTebirJ0aOWW5AvAuAL6Qyaijr6yDQBoZbgbd5XvoX2utcyLJR
weRYaDQn1oYuecEPbqdod0uPImBVIdSfdbATqVPIAuiH1TVAJcY6a51uagh6hPjz
V2M3rOcr9hpo4s4CgksV6KnQrkXwtr+XavAXqdn6XSKwpewxgKNJMRM86hFQ2+h+
E1bGkXFMGDkfJxJokX7Vey+0STO0s3U9YATECChQZtgJftkEpHTF3EHUHRMKVNTd
gl7BY02FWbl9xaNu3FEVYZF4RYn1OlZbA6mLxTEYHqAQliNt+O3ocNdJzwAXKnbC
cvAiaNDoaAEazKOyNOf1B/xFN1QKyapmHTjif2hYZ5jJipZTwevwtckEaIFvqTOa
/eZ8OcnrM2eHIStcIVHCttPHORsBRWwBDDA7UiPMTCSrdLUJ5GeBdWufIgsHlJB3
8+WcE3nhYxXvnycO8D7jxuBfd95nHWp8l+fJ32xqMPpax0u5t9Fg93s7eJu69k05
OpdOcVvRIwm2kAp0jJDKpsDEcgsjv5Oj1Ui5UavK0qdgLjzcC3nTpJw3WFe+96hC
UEDQ5nsRyzBamuGRjswLh9D6F9Dy2SEBisRkfuiTZfW4MahiuQW/wAScrArPWX9N
f80TXvmIvlVTunpJTTU1R0gpTcGGSBYfy4f8r8Ozp/400aFGKceKLtl8SJZsII8u
EGdTyx4T7EfsS30pI7JKMMDJ6L6ebFzswR2Kix7eQ0CAJ0oMqZKivXlEY2QzWPMX
DCk8Q0DNqxaASIj/C8WVwmjbLOSvf4vuDkPP6gOcEKZeMJOV/6VxJHVlry1J7IRw
giSVATUbWWwanxvpe4usXhQnxoUheqJFM9JnWRPFSOexD+NEN6U6JGdSVof42iEm
KUntDtV7ILByGNnLexIpAiZCWckCZJ7CZcg/2UIMCG1vgHpSKTjGPe2GgpJDH3Ls
38+ncI28RgcSGXmmUUHQKaXSKTUY1Vv8BQmk6Srrz35qs0IV6+Jz/nbMlDElw3ks
4MqNvwrnSf2YlqdIMugOEJX/ZHwBQCMX36IKDPGHtwX2T204Keq1PedG80AFCVSz
7TEy8+ze27Yc7Av0qTwI15omc5qVbm25GrLM4yuApuHRvT7p51vKhe15abTIcaa8
ENuvYxky/lwSPQlSsHDJKviF3Qz7yC739tgcfleBhigbMHqmGgGPWU0aYmUmjmRA
tZ4PUltkzDW3BR6bVxxtr5yQzI/tkgzNr++tWb5IxO+Zk8VFkv4vzP+r8h3SOtP7
PlKMHYREIeXErL/PO/+TCirE0eMkQa7kxqiN6t0k9d9BCXJDLhneTKWo8/AsAbif
EZj9rVhlpPfzBf16TmDi0rgm3t4Lp5PijB0dhEf6AhIdL+NHhafWEiuvxYTZa9uI
ATC0rXHArV4iPLCPtj65QzHRJznI3Nfv6jF4l68arxkVd7c0hRcbP39Xn5hPKzgE
xpVpJ/kSaJmPPReRGxNicUdOUZigMXx+R6ptZw9WGdwNkEv6xB8PoPnIcT1YQpX2
IdnuRHy2NXrX79O/yp7iAh1p2fs3zWWxxK/Ny812cQE2UTtHN460a+1ZPhEpHcj+
KiVgm1KdETpc3uX1PbMP0arhi+JWEjBRpzD4Z/88z1Zp+L8jIaXvOgTs2EU2hESc
SHS63EG8Cjmt2ULyp60y7gpYQ9X3QQ+dHIMgAP3kxhIyw6OoseDoEAgHU5dddGs/
btm0agg+CDI17B0N0/ftOE0pmVMVztEekmPwYr337ZoHIURIrWc6J5P3qyk0IA2o
FuAcqmaX8SH43+Dw3sbPmlrLPbd3ByNoxDf/4I5cWWlzW1UJi9ZupvF/yEbcZapa
cIAIG37tjhkujEu8ccMe20ujbrGKkovpQePwWE3pgg9WRgzCTmTltcs8AzE1gfOb
p0oESuVOmZG3IJpLFknf+++EgmWIUMevZat3hmqZQlu4j6nVJgULsa0xRdkkRjLL
HbGiAivvi46OqWto7AcB2zMXvCoZOGnftziy12O9UAcuu1vNRodDgjrLhrkk16iz
TUCzQcXXzx2sV/cwK20Ia4FhEycavuTu8kL5NWKWni6MfaD5fSOn/EXBuWr5bB9I
Aqez+/ORw6gT+rNAirJErHJtAYMgvGCjFYXJNNgHcYbVmW1rirM6W3LOfaWEDCtw
y6re2ZrvFULmTRZg/xX0HqbE1/XdwX1EBUysmitvcPto1GSheqsHNz6GW02yyDyF
hvYM3pSpi/cDv8iHJMvAR+wzaSBnhKvbAGZYWfEusMqvGeR87EmDiGD1LGSofPEx
hdnSJukWS5RtrXhgFLXhCTj7l0pPRs9399E43hgeCDQciFe9ZAQ7qNjhSfoqx78H
EV8YOKMZ/tyE6cKyqQ7GbjCBrddZrmFZ/bIKrFp2oBrPCXbTwwx4i5lYrLP9yteU
8SIn9DJ71MwcburyyOp4/QbG0cvjgRtZDX0aWT93NLXO1fzaqkei1IajXeOFM9Ua
9nx9L3cCGaZ68/BZUBeH1CCSsTkAG4NrSuM9/c1CLOhFgYffXIPr3iFwLKexkzSe
1Smuc84bFZSMvx1RhWbEGz1UKuupABPqntCP7ZUHmTJNyrsYj8+H/KGIFf6YtIlU
4xRyVtAoor5yX544EF1j437hIiKBbdBA4Pjpug3b/NBUW3g7vaZ6BWlooSrVMo+r
2aUPPOwys5njNVH9ew06iJPeeup79ib1ULIITsDBWdJv6sZJ9ZzOXKBgPyUs0dpx
jSoF00M4Iv1FaDd5Z5h3t6SQBEro+7agdHSVoYG2zSgzQFJId5dBhimBU2Ofa+3f
4+ZZ7t60mweywiAkOhP+XlmGj1o262DwuE3nhKvvV3uPU5Lv3h7VtLeMAqSlF9EA
5/9eAHYWIVRZWcuBmTTtpkc3mHHiPTfIKW/nhvjh+cP+MuiMBmcDvS99nd/5AA7P
pF0lIQGsOvFzZDD2UqTw3e8FH7oiUmBaScOh+FgkWrgxMe6K6f6Vq8Wg5X4eNm91
A8Gz3PUFmAgD0n2HWB3n8Wbz0BwqFOWwDM8qRUhXKY0kpfedlHMZSPc1s4yaPgkN
eK43Z22Fw2LVKPfPq/EpbW24jbatxxoQiLGsoya8yNT9nyDx8qf+HisG+IL8IqCw
wK7w/9KmKoHmoYb2f9l+7Hrw/Twb62OBzrWsw8QSWNeb5xG8jW258VSaiieU1qJq
1ZnHD0nm92AhF8TjZYxnMm96iqekpADz63wDBK7kFci42+tjR7Ek9nnW7PCsZeRo
PhhEOoO5GVm/XrvsMx2xP/IUYtWv4WbfVrtQf1LjKQfIWuNNMQt54xCkkZXGXVkj
dkpnj5CZOf/IdsAWOyRnNQyLnOfdwFh3CDXXbFnQUCgXCdvUXTaYNETBE3QFxzE2
zzY5s/vz/kmuTUUKg2jSozt0BbV89NwVP2SYiZua1aiql+v2OQx2rKCyH3F4zlWm
khL9X5bAV37P/oLR4rPAKap0LlQFMH/ALIDEqKl5Evzr72WZ4nLGAN9fSCD0JtLZ
NGy4JEenDObE7uDhvY2LPYKGhX3NbREqO6CKMgq2Go3iXedithE6TdyVt1YVBqDw
UNfiOF7tAJg1RfDzqgbWk8fbtOU+aWzGEoFLRZMk17JpWS5+695E4VrcQIk4kQmh
UVMA62UykV+UFW1ZjWvkGXA+vrXbru/WfYKzaK1vO+6JR8nTcLYM1xUZL2fMChti
ySZuQRotjQ0XPjMUmqCzZ+7RnV6wEsk8I3dBNjKLlpHU8vO1IyCqjVxFW8dtXyay
mbktm0stArQYsPeTHeT6ukjwNq7QaD5InQvPw7MffTXUpPfIGUMS3NLiDj73wbk4
ydQsHd0rjhOKFI7HU36UKHxc7xUlLiPhsRA53MW5x4cC0y5hI0uUj0gI6SjFOz5Y
XK8GdApiO1TV1m67j1Kzzdq8NQJcAWtt8mMDwCnfHtYkDR27wCSzMuvAE9FyAwIQ
qJtNtnnpvjq03QctKZR5cVOfg4e1ZFkWl3x5AD7RBHJilWSQ0bFowopNHWMi2Vwm
18VIy5a2NfFPyW7GvJkcsbl7yNGhHdPXBOHkqEqGdVXEV8vBeTE6wf6rAUBOcL/Y
N76qULzxBn6a2cANBI3S8ZwjfxtYGxq6jUig84eTo1cs0tlkCYPetdM92bg8V5d+
UULtneMZV9H0T+AcXgxts5vh0ePyDoWzpFbR+fpK4xrN+qVlV+ZBRZwC2VnAdKTy
NPXhu7sv3F+lGF83AniV0ZfVLTZtfolkVPdPRzBH3j0MXqFeLfewOK5eP+sTsk8t
xfcSg3HNfiupz2SozKEzRdHlzknQlNAVq8lCPC4AkEmtwLiIz+jQXTd2kr7aeC7L
oXh83KvqAesKkchoN6ws2K1lmAukca1J5s2UTgTsLmLdLlRwCY4KPmXDVs6EkXCy
KO+LgeD85SJWFTxF+ifABGX5ErQBlzF+R3+2wkXOeIWfcwpIbIvr+BAXcQqgLl5U
x7j9UtvYjuwDIojjZonJGBV8cN7zJippwVMcmAdoRQ4urscfwaFqEX/DkiHFA9z+
DlwBnWrfz0uqT/8xnmQOYl2kOl8YJZ6TAR8S0V9L1m473r635VouV+ze3slP9Cpf
eP8SifNK7R3yURxRZ3iFWhztuGTNGvTHYPS2/E3r8liNw2a7V7REDFpbNrvyX9tX
s41dUXL6qiW4cQxNZHVgIh4geShLTGHDbsyTw7rw6BuV+O+wh5cYwllU8MG37ggR
+N9vvc/R3e6q2XKAHOsLS4mpkeqmgfuyF+wmmMFno6Le/IuoEkIox94lE1o8G52C
0tjf3Q/xURx0OaROMN7okGRr3odTJkHdKTgtB6oB1Fpb3tDRN3D8S0367B4oCVnL
Dq25kXXXles6HweFm3IL1/EBY1nawyzXupaqv1hEx1eqroo4HS840X7hrHEOtW2y
Lld5/vYc5gtyxIYPYJTX5ui1+5NI3mViPqpVBTEMbXMYrCDXgvtkhb2ry6UXsMwO
1+jloQ1pWcn5eZ3oxlaVxpoC9zPkQmhr44vob8S7b1dBxg6UhIQoe7dTnu6RoRLj
z6N7+1rUXhqoC0hG4mHy0StYcRk673rlFgnqT3Wp/RwUDCgTM/uU+ir/XlRiFNMY
e/CjZBt6tOcdX/HsJIATrk67+ThaFqwJ1CcWWw7hCulMt2pXP87pdzmZndioVNRe
f6lm2XYrw/x8VEevfA5OQiDPkJdmQaVSduIpbTGt1f38dOuilZ/KODy4g37oeLHB
/zhBk9ScF/LQwqAdSlrMuuRj6ZmNDBczWpowSUO2u1O21C0URs4WWJewn7lTrswe
TMyoH4UyM7BzF3CepWe7fPlE1E1aGEB8vwpn55PfsR2TjNAB11A4NKmvZY2WOK6Y
9uh6STBCAdCgL1eu3Gyur7Qnw0vhlj+NE4s0q48PKi3H3dkcbQ6qMt+MLrq4hV0/
PvaLRXuvn8Ufw7XNDtJJ/M7Kq5YCeJ/c7qt4Lh7ocT6Enqrmy649qDPTxKao06iX
vBBKq/gAiz1kMJOyZ6WYitwnKk4WGgPTLzi+vIRDOuGwclV1UkPVkv2/ZJn5Qf/Z
9o3Yi/eBS0sboJ3aVcmcxy61W8ZpZPp08erF/wXMTjLnLTmRxSva/mWqf2gVZVP9
tmkhqtvJMJzvMkhfrnvWwA==
`protect END_PROTECTED
