`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7+LbFsnC/j+kccpaOlX5nkcVwCL3EMQCPwx+KaEcj37YLQ2cErfEBlYcQtMO9ko
uPws5XJqFNhUV2qdmcNsY/hmbDY0K4Nur4tupGxM57Da7auYMl4IHSUNUiFYaO4h
em8I0GRYr8NQF77R6J1lSgv/CXagyVI9qMhn5tr5WLPhiba39lB2ySmBDWxPRscI
qYBypn0ckethuS4sBgE73dTVQtv5D/Z3O0gPXCTuL3/sG7LhPecbgTXiks2znar0
TRavZvskajcdjr/XHzEMdTorkhgdOCz4apLWef1UFGcDZvnwe+BvbU05J/SNqgAj
iMIWskhW45ior0Libpy6XVCY6EYKRyk6nvYQw7a1hxnzaPvrBoPj/y1jeZxRkduQ
45yUHYsjcKoWY/tHIbW0c61+xB0ggtcmriPr0+yhA6QsAcFKl+glB6TmxQrzxhbb
Z1hJJVyJ11hQioF42h0jwYwPO/jdkNdTsxW015IgQuZaDL+E2wuTaIyHitdybTwu
m3F2sy4OZ7w14krC2giR/JPSLQ6OKYbxjZPBiX86XjAy6NOZeQsBNoBRh40+2vZp
XduCAF5UEZ+a0hliTkC7cgGHNkzCFFRjpQ8ca4Dm1j4Xkvftar9AB4kd9PUCDcvj
FpY9e3FLIkEyYWrnqNM/F5Ziiv55Qk9Q/J2apVY8BodjgGfJhB3a2cvih62eWcv2
bTk/9wIjIGlUPLGnnNOrTXQeRUDnQkf1Ca2KbtFELUOLILSiUODUaN11SkyFou3F
vGytQygspCbRBopne7guufkjQXjPWue0DbOJjk6AOUdVlPGBuCXlWmcoF9hhhp7B
QnhW/+z3MpnZZMiUBKvvC4MaKSxrayunMtZYyS0I1/hszKtd/zBE9gHTILWIlhmL
STdMhmEouUgQNYbLKabiZOsbRr+OO1JYUojw+wu4ie2WAm+HS/5i1JtlqdLF/6K5
wuCM5pRbkjwmvWOikJi2x4TvSy/II38fBWMidGUyY18n7kZ/FgicHh1I2xrGrix9
MSc6UTPgK4bw1ufFt5gB7m+dHfV6XlZVGw8A8p170AR5QPMHYTB/HF7+A9M/7JRL
iGmd4VpJcLI9f4uRFE4QZaq2Vd/xMe3BcQej6/nK8FQLRyqwmMAN7TkEFSwWRfCK
oAtDGV4tDdJCPXb/msVhPqjCjHD93mz20Vz81bk4rqTDijBVIqUpCX26ctM5owaI
gY8H3gSEhOex9/le24kLSaaSHZSABButMQm9VaZM28qbIOYM7TKG+gfISdfiHT9m
vbQTj/WzuZQEDyybKJobFzM/QjyLQYbhWWXJMnu7nsaNSzjzYB8XN8bTDp0v7+Yy
LD7oiDbf3LURk/ePeDrfqwiKW//L64LEyIQY+gnt6yFIBFXigtktkgQP3IwmXxx/
38c63pdAlesiKz1t9Hs4myTLq8TwnqK5WNP1zWX2xEDalIvG82Zkadkxs+QzuESc
GvgEcJfg99Z5rkoxJ8v60luCZHXl01IPQLIDOl6JSSbFp+M6i7IRAuBDCT8/Jo0h
qAawBE+w5sC7nmc9q5PbJRczWMJObib/tvxDUW4a0rY0VHVJrhd3Bu0euxRLlvn3
9Nl5BeKmX25ZL8z6r2CGgnTV86ISiEbw9adlTdoAKFnvj1OpYnIxk4JlR1CxqXMe
61kyIvQc1ieteMRVRlnbeOY/R+XUQmDmlavqw5ouX9ynSKLwqBVmT9XZke0OdbFU
4KDevYPfhLH7XRlUBKPMUdMhC2mCBaO9vzZBc7zXpybPUbM3JZUER5/K1hoUpYnP
iu3d2lu7/q9J49WBd8PR8L4VQb7I2K2US2W0P0f2QgHtnNhBFHR/ULCUOpu2xxJ7
gjrcRRltITWblmTiF7EeEPzSdCZHWHvwkF8mKO6RmTBvgQSRvUTovFmGD9wOo8m/
OhkO+tNhK6fbz6SJalQQ39oQ86BK9OLuykwfJjuuJz7yalaaLXl1mxZ9k8uaqggu
xGIo2TvRt65HncREgjBpKEVdsSpMaGhPiIQ1tzRkqRZQkIY9TIk79PvKg9hv0d09
4VcYg4oRthglwCA1WkN7NP847BSiwubm1DSat0Cu597o8dUkQCVFUg2IoxFjb4FG
pPtKNaWmrYgWV/gaFKHXw54cbhMCkRMcwFBddHxbPFj/Nesmcq84rPTsOS7i1aoA
1s/1osm+xhLviir67mdw1QQq9pG2YtBPTGT2BgL7aqp4KRC9HVQehp9L1Yaz7DAD
9tFxM8ZTuFLAwhwM2AMIId5xNVxGR1Y2alSBm8RU2dMqTG2bhav47SylEF6/A9qx
oZAMcmf3VtzZ/zTwBiOv1mxkFVL25H9LLkegpT5zoEumlnhHMJ0R2pkFPUARBxnx
fBYI3Jg5i8VnHLe6s9j37Z4YtVUHQiNjX24ruukan56E+eiJioq7KmXG3VUO6HN/
a9lW1dj3kGQsr28tzYR3iJcNbffPbZSVOrpAnWner6GQ1zVNwnCK0mGqwydelcvl
VDKLNk5Hq60+7FziXGzHlxCPOCOEm7qZOIorLNO05LVTUskpY8IiNVHHbx4QeMML
nRdgFTiejQg+H65EbtwbqbOfUCg87V4DQlfUZ2X/eLtAgBJnou7/6/AW9e21sDuz
Jpf7TVfhfaNuyu+u0qEeBKNqdFe4LADcAN0iyswk9dC0Lvsalmq1uxUoLH6RKkxj
vZEPqsOY3w2IDhAjXhd8U2uYJ9zQ1zQzkz59Wczsgp6tFNa+67BU0PJnZ+7faOWJ
3Pn0Zz4JUvxve3uGXunLw3VqqDdrbP79gEGvTLIFso32YiR9nl2hwLnCQhGQjan8
BnuYajuE93tCEd9L4asOVeJ4o2g6qy2AutnKHtT/NjQ+xeqMJRnLsSnVgTfLf6ET
0cseia9iBUjt6vt+2+puiB4BNYcFhB2mF/fa0TCLBYAYxahvNGah0LXrre8tJphE
khKH5G8ti+TxNnif+YedapNmDBNAyCfxxIWG+OBogGGVaSX9FD32/ZJj4B0hGARw
HKl+hSMg8MF+dNlG7YiV6eB5j78vW8UIpStnoz+vVrQqTsOMls2X0a5UddkaS3iY
a+yaUIn83+w3CuCjzZX+u0QPnB5jJGpBr/RayHqyMqtSD+g7VLV4jnpMDCnvk7Hv
6Cd1Y8ewQjxhyCJo//hWV2byiLpzhyzetuN2i3gYpubLAuKX7aZwqAU9s6UCSiJl
7eJXd3OGEACcuxK7HqcgEl/E3E5t+sSU9EIs152HbqsNDIyPWRcVohOY6lL9uBKM
NjtTbonfV2lXN8nvx1cUh26Gy+a81AdZgkHjHrXY4x/1W74bZPcsIFp9OFZCt3nu
oC0tSSd08auyeFG1h5LS9GVcQd0sa937fE5z4Ak+O/zgcuyW7VSCXeDyzapMIcFO
YouOZl1wpbF69/n9OIDx9L0kzQrbUpuMGhilnpuziyb/UKVm5YKnUFE0inJ243tA
8LChOajNaXpimizyqDbM76ASlA0tZxmpoahyN181t5BTd9tqThHut4StMaOnGAyL
eg17VuUCScRdk61fnE7jZ4Ul6o4xEx0wUKQmqRp528MGHbXB40EJV7qXClNY24aX
xat/zXgTER1gF8PSHCm6JFlS850neorAioH5CBgje4ga+376HmNlPUxUvBB7RGWI
e8uYUglAFUXgeJOCVw4kKnd0vrkePDr2PqIVI0eIgP5xYGeo9jXbu5DARNTkkWrR
Hw41xYF8kNxwY4HMNvWFjGkLGv6hIZH1UqjiGX+NU5AhcD2QqyDSwpdUHm+/fvO0
m3oh6hWJoCLntHidKj9Jdy9dIRkCqqOZmEpVL/6coTLrFGzUTlqSdUAVrP/fRtyA
SKQQUQOz7SFtB2BDME6k0CM6PWV+vOJH3leX9cKOHKT6zgjMdzvKxMUIC6qRRIcN
lsmN8bRxxoNC3v210qwBkCnpyLNz9W+wD7sOCj5w5CKQ0OP5HvQHQaBdcMcg7dwb
/wAdoavYk8m0xePAx1h3iP6s3pYK7STVIbFwPMfABHLaf06YgFzoasrrQoJ2OSnJ
+PrFP/ulck4NecyUG+iARQeGky/KwgNvwI/nEmXLK7nxiCWCMh4zSadl/mmTU6Kr
xCWPOkPrSbpFBaUts13fU2+IQP5RSRRYMmQNI8etjOj9gsV2EIpUsdhH7Gi9Ac5j
Gr0/VqQe1Z4R8MqYt59qLg0/L9b/xvu2RbDB4EXfQVMrXXKfsvPVGZJpu8G8rN4F
C1f1gjYkm3foMQmgQVkTWwbfqHqyttpqWSl1Fl8+O/id7B9Hm7lk57+FoRhyTTjU
tbBiQk6hnzd+gRzGTI/EFl1gPi6cKhSfUPbIcHx5dr7cIcx00zN7cp5T6neqytSD
h4DXeHL/Temsdrgsl4I6stPaDXeh8q/waKEH9op/z0CH1KPZvy48R07NH6jivlNa
dgtic7R++Ng1dylvXVDol6kpJzjD/v6ADYSWbxW++Nz8KtA1/zCMmR2wAYUjufka
DDL4Vf+wIRHsdVU4vJc1MTi3CaMaGebgFxPVLYQ+KKgzf2R30it4zsVWrOImq3Tr
X+dZaBqaMeV5OZL6fculSGmWjMGvgSpLPWYEIHQ1NOWvcg8Aj7v7PlbmsroecQpu
JsXtWbHCf0ruAo3Iynx75pNH/77UVzQ9LF6SSm/kbi6EEckEUPRFI06xuFX4E8vH
WiZGyW8z8oHN68KjPsHNrBMBSkUOiah1pMUxh+Akh08hoMX0bXBIRg3XtrlJVROV
uade4gktU5I8Mzc59ixqZ/QAQRG6/eRTF/laJ66jZXOC5scViG7/ttEV5p8xOOsp
hWIJ18plb16q3pasRqFdUhw3WY4286ZZ40J1opKOIVGnMoox+t7IgGhBYgZfMJVO
objpjXJ0DtsaH9AuAQpDftX+nulERUvTCyhbAuxD3wpKqj9wLNx1zyecJADauCFc
LszUR9DSeq/mPY/zGHJrD1EeHooJztW7WIqKOcXHXlW5HukK8f6TEL2iGyVRPOHy
e7+yL3Ji4dc5+uyFXsfwTmJWJAyYrs/eGnZv5779GTuJY/XZ+U4DTUuNwGQ39wbm
CbMhZ9cl+XVlDd/dqvu5XRrO8mfZYFwIJwY0An7akZnfAXPTho6OCrBYaLcKG43F
Up5kBw1FJbWTlLeOySrle+o0C6LMtCSXPvhQTqoRjQ5OzUj8VICfaTFvO5Qo2cuG
T6LUF/t/WgexD4Xli63/HMI3PUMCg/Klv0qt+hw4677QsXY6CJy+Yp57GdTteR9m
gBrnjciIaRS5zvFcWlpt26XTbnmqfQAlA2lq8dJ18FzX0koMVCxgscG6qo4H4bgh
WQjhs6wJFbNK+/7qPT1hzFsdEQWWQhQ6Q0WKHlG2pFjxvivf6MLHzNgAkhaPQmZq
yloYMB575BkcFd5mztnPWPRCGkS53QT9E24JwpMOQENAXElmpISv98AIokIgeHYQ
P4IGriOy3iUn/ZY/MJJ2rTK3jQhDipH3tLuY8noug1Kxy/tZlgy7LKl0svbv6Pt1
YQm4lrt/dyX9/JTfKt+uxV3BECAruDA0nyDWasU9RTJYiJdJDLV/UBPnrk/6YPaX
KkhHhv5M9gY5eAP5PBU7Z23f0ASdexD7+YxufDlvlr3X6pO58X/D+tnPvRX/j5p1
FbP8oReG9joiTy8Spi8LXut1FDM7tPhAS/zI5JNmr73yRsoSJWigXLjj8+K1uj2l
AsiipMdYmxoVePLn8QX8ef7V9tCekd8JDD78jGZy/vVoNCbBM+8c91i2d6U3qPh+
+8WozGOVNSclmh8frr3xIDxnwvKr3duZXs9mFf1CMME6NX8N0ehM14Fvyg/oVDX6
MyhdJQGYRvi2AfWlbNKaEwCQu74VJl2GQDQiZh+wC92L2O0FsVreCGv+vTgE0rNA
rWXVdlh+ytqeiNtYR/OT+4JieBJPWeKD3JrsjPEhDmsSjlAOB/ckb4/vJTCo04yP
hcl1F0lgqcWJSElnAxC+sfLKqMcI3udPSpZTWYSIargE/r48+g38d0JKx5vRst4y
LBNF6NWnYFT9ssUs+ebcrWWboRpyjlUAJmK0KkE4mTcZYUf4VaVLzXfmF0Dgc+Yc
meXDvtbPqPn6htM9XK5XHOK3WbTCTdOyBhctCWc5Y0sfup/gYxY2dXW9A2ephXo7
9r5zH/Ej5jYoG0aP/LtqsLxLx9wqSWdmH9umNWqG2SGcEI9v34W1+X480m2JaZsK
aPVsTfpyAG1+mmcROhvWo4MkDjpK1cm5DA+b8gFGQBQFCgVxRHvPwQgJsht/MvNG
XCQ0juw/NOZxR0Wv0fYv7jdgD7lvr00Xg5MZh5aAvXfTRLSHxrXFGhpdGigfLfb4
yMsc3qdJS0fy1tlJfDG6014VahVYtSGjf2JehafpLjKifpNYdtomCGqlH1hQOZGC
Q99No7BLl/0YEs6ZM09+Bgl9VMga0STAOP1RnbDDF2hALZIy8y+c90ONBgp9FGJr
ktMNnYGE+ouOUDLjz6COcengy4bIB2w92lc3OJEICZq3G8nsMo6gcPf89qF9IREw
TjeXB+odn6ex36IfUcymZHoK3SFFITEV11oG1hxUzD9JJWyzZE1q3CTs+o5sN+pc
AfaI0I3ztmDS082AdiNCm1ajAuhVsmOIa1ZXcg8R/XplHpemgb95kLyjKXxZDn0x
tict4oBTLC4AXuQQ0g4J8xkRQsVIrXyyumxwCcT3W57+Tqmu7FkUiZGQTioT1svi
HaWHxJLvXSle30W4OmiBQ1HrS0xOmLfYoOtvyhNaI7h9QYbphjoZhaxZd/OhecJN
zhZL4KpR/N/hTgHhsSWlYo7OAyefwhWIVC27L+NBLDBdWZZvhxepIN/4gpBR82Nx
Ntq0TNMsk/zWTqiVu4u6GC6+3RO6+I176/70qFkpZky6H2mjSNh5WvJ4Rhyeb0oz
nhPPXzjgkgBbkV8sqlbtQRe7s3ZaVZHnBxBBfU0lwrIEJ3I3Bcs2DoyNnA0WAkwr
2UvLmcwWwgIBQM1low5iCJLKFENnyvzX8d8bktHnfcQR+frjsd8CYVY+n/kVb510
/Yb6f0GuRfDaVCKEz0HmH+v/SlCPCL7ZJj/sUulkRDOK5lEmRcyC6HijqPdLOu5U
49X5/ycc6kdGjEVJj6LSvwbkXYmTEcADlP87LVuFXrgwo0XDegyi6waHgiWNyIxI
FjxwIoYhVwEwIllhtx8GF49jaJ9fu+wmOjsdIVJbXSeWbuNAaa1nwuAc/CRkaxOL
Y10cpcYkJRGeNQ6WyBQh/Q/WuprAiJf8qFCE+KunXrGSrNvSPAZdv+u4C+joAgWl
hcZ64i+exsA8gT4qqLdX31vYEiLlFUlN909olNKMR708Js7EEEgf34M4+Z85+TSC
TsnkbVyC8LTmZAzA7TlZoNwpizvVgRVsz3zCrUDH/4bio9KUJhXw6Z8DNahDcUfK
v4H5sMAO6YTMCH8xU8CRc/Z+p/v7UwlG6RWNs2p6QbEAtJ3j9PY6JMTR4XS2HNcp
Y4us3+iQiQjk9wjlneF22ZrZJJC1db14OKqRdPiAYdfrTVDbLtBM+0+9n7vyP4Nz
g/KJZv+boMESS6H4g8lNcBbbMxa/3j5KIMTO2pahiltiFS6+cp3M87vxZ2lMm414
1now2h7FYYMRpVv3OI01P+4QozxBpRlR0dnnwY7alQDBs5hDxh/ee3flbJfpy1Ws
PfBbrZfvIU+WqN1QDgYYnAy973O9Ulm5dZhF+srLWrl5S/9W7k6zEMrObKXVoH8d
e1pm5/ftEFdnNiuzRvX3aotaP0ptz62x40c+fztnq3Og+aah19JG1h61LCg6Kk70
/YwuzM+BM3YZYitcfadRTWkOSL/+OC3qFHbsSo14ehk5tSgo0DUBc5JAbywhgCDA
WHjaNPNY9+ZVTNVCMTeg+4KCOY/2Grub2sqZvJ/O/3uhOSXKaGg+95pkuUqPbylj
yzDSAY0iiKcCG+jYEIAS0RfQ3mfGhYLjgOVil7mTK4k372eU+yX+3YRvcge7zwW+
v4AhEDcIoLJKZnJX+0ysfWoiNlEqdnH5YiV9h2o3heYKwiFjdrA//vsGdvsAWAOs
HhO9+SgI3SQym3gNYJCG5m8xlHcjEMEBmuTFeNImjOoVKC1bcNMEi3y6lwKOsszI
s5j6X0cUhRLTwxAN9m0Yh95SkVgbjBXwa9TVZG87T9NhJgAA7EpCC5d0hnw4ttQM
D9r1SXgJ2Hvn46Z6VfYIMkKyXzKtkxeaZXDMIgAMmL77sUrBwJdmiPLoXh712k14
KZb3nleQnBpC9mRfCjq4XwYvZUIpHPYG+OyGWct9qPIVh0b3R+rD6TB46THtXNIb
qFk2PT2twogYVIXsglQVawAaBcXlhCFTaCgZNhipON2N503pykAceK/bPuaCF1W2
tj9sg0eBeRJdu05oRPnbYVIbLVxWfMe62f8PNpZUtz0LtCG2IDsl6Vw89rL1PdKn
Y5uPNY0cPf4INunNHumCJQkodSHyme/yMrKJfhpN4bHJ6KSgVr0y51kcegewscUR
A/oL/dnQBaNK6LuuypgqrLxKHOYMjhPiQF8y0WGUkwidY3fNwSnaDJ9qrNHbz1B3
U22dVSzKd5MK1Ksi2JTpZFq3Y65km02nFoI6brbANrXav0qF6PYyiuvSgPxVtCC0
j2o8YfSKm2dW6CQ7im9UlrjjvrTx1TGC8o0yoBUgS4Khubw2z1GvJyx96DsTRa2T
nBeqbRVmRTGnKz2Abl2fXSPCL5LmGJdFEcPBLsGO7BWjN/IfcX0dpL/Oc2kretYF
9UTBXBxU1v0tsAUkBGLcON3k12VoujNMU1cl9pC3N+cAxI27Zw2xV1VM+wKD6U67
0k9+MaYvl+v8iN1RY6DbBEDGczt3acize7UDsxTlYTzzfjv/UMVC+2vmAa/kV1+X
XKlEPHkXeAFCr4xuO9hN0lcw8Bnw8JBPVlluYkrHKXYJW+RMpZBYYuW8Doe80xex
awGCz+oG74kfbnbiJZuMLbLPOXx5KSqD4uOeG/hBPudClBwVATjGq4ZNdehAwMpu
ezpQadVfGOpIqQpUB7GC96SXDbbFEu2chfzTGhX65YPBD1F2Sz0pgfjuMp4LpyjQ
5IVQ26urZ4uTeCmCMARsFNof0Y98MyruyXfSAq6e5NrGuPvTzfsljOKhlC/80rFT
VAVXXbJnQwqGW9IC/PgLASC4+tY9xYjwALc+4yV9pDLcVWQDLSsTSprCcW/zDga2
18yDmZVsosj0LphfkV4De8bTjCKSorS7qjn3ibdislpnQ6Ej8KtkAMOPAarwZwI+
6idJLUC6oIO+tnS/fKAcyELxe0glljJFhKVu4cMc2oub89I5lgH8PGqIvPLtlKFh
RAyzIUddoondZDI+e/ZU3N3/ssxMPD8H/LkMKkx//oJr0ZEKZhWwK6Vp4lHExnI+
sUlpt6ZMhaFD1xToJ3PuSWXuYzLbowf0lGpjgkIDrCSzK+teYzLDaHZgmiPjlr14
Hz0lp3iDSerXeL8HS7LIB8+MXxR5hYFSeIM4+adfXXfCd1ifwv1DGj1OykTuctgP
/izO60yLCi5zcjwhtrPvWkjYl6yMu94bjdn3zi6Y4b2mpa2BY0URFk3K9wPo6OYM
El7bQjvfSi9pEtv+rMwbaLLwo6xTGlofrUcANgvHprnmfe3+cxCrjuKMPqP69IHN
G2lB7dEDrosHBNm9HjIQH6rTXRPvbJR34KKWzHCBcGC4NzKJcSg60fTJsR3rNSr+
ItUXAs2VEXg0XsQ+GWb37iLi1p0P2oSBaEJCGv9/9BjYcQgOz7Ebq7aPzuB/mgHf
LdwziUGUch2dxbYkmF2B3Km9qkFd3FMaP1v8urmn/Ikp02D51SEjeOFtMCp4KR7c
5MbMp0Av2RBshf4XPYoeCXSLKt8KJMKxgkxpLAIM/zYDfJqIKQN9q6NSdMIkuh4c
YB+m6nFQ6YTtsYbevWg5+QbVCO3w2An5Zk3oj04M5F+mQJlR4YQtSDDLdCvDWZ25
JBVriDiuo+BMnvUMZVi0U5f552Kik4UJLzB+sP6sicZhOSlgvq4VTztn8kpV7bQb
4kOXlXVupNQ1uwB9QJeb1uLNoD8OICOryrBeO3jn8A0lTcgPcTPwgr/i/MPVKRJK
sJQOdkZ/+uwEqSp4HzaryVjr/D7gGehXKq7BG0nsREDCprZUvq8NUyXqBQgJvZBd
sCYBFevRbdbzX3yC/GFWsMzHp8b48gO+4/8TIHPAPLbNkZsOew/hOGot+SR5Gl+m
U7ruXSHJGoL9pstwjuFam+GZVEOPL+o/xuldyPO4VczXW/Yfm3kVQolb4Iz+0xPg
26F7soY3BGLk5v123rw1603wbTyGFOU6GNzdvvKxMkYn9VxIMoPOZoj31sOAaXco
R5V2SknbLu12FawspbKTmVHrNEIkfWwHcGjnBFtoHp90iHH1H51b/NTFew4ImRWw
Axo4dA3HKm+8s7AUdYXKopMYrsiL0Wgz7/wb2z0iJfshtoIMP+EmbCgh8bu6/6Me
iISWYUyGPyHbKic1bpQH7Ief11SFyR00ausrlZXBoqp3c1qkK8wT2KJqNZlDMUW3
PBrDPyUtgqLiyqxFjUkLK8NgX3YNA9kDb4KUk8ikJJiUlCNPpfilqr9+vszV78fU
OXQUc3LcfNbRsmmvIFtgw3VbPWpTeUqGg9jwRlOQpHFjH16uCklkCIIX/cMBKJQ6
60EtzaLOa4T1M1gwMkrrSbwCOuOd1zXRbdrsROhwymVt2ay+cHfvgYxjNOyLgQuV
6h9GL9/3vz8L8tdmq8duRp5E4mKuXCGdvVrWOTymVvs92mjJd7xvODFFiBUAjB46
3a1uVPsg8RkgkF8iBoyvouS62XkgGA9l/sYxOnnaB0rq3LhaJ0d4KntojxXqKEkB
IXSqkY98V1pNamhGEqXWklkKRw0l7TQYFGfl7AaMF3QNxkhKpuCn661Zvd10Exn6
ZvwHG5sHr+bIr99MXTRnYXR6PZbU0GSDL/nVIpbmzCdqD7NuZ+Zf3rXLrtYnz5So
8juTe0l2+/6oeOFlQHKAy+bXhJDuudNFj/BeYtdYpMQLShBWW9ikMHb2YmP/QA/g
0YHtpEutjolksGiJPvU14DqEsvvOYpb9gdD4t8hcJDzlh0Yoy3Pz0lKGa9hDmFEt
EQVIZvBm8GuwRzFRKImzdb46K+6CF5PYpmWUp52w0rVBnRpYwq3TVTKbLpUC3kjG
lxOXEyHFeQULlRDWrCmzRF5sok9YBZ7eQvtQocXz1rhZbjc3wG98PYduNaQcpHD1
3aT8If7Hk9HLDLRtx/L8NQt3eLI2ItD97ZJNrYTT3oPmozREXuESLzB/xmXfRSYF
C1JMzKYtCP1+iBea/pCgZfWxy1NJYdGpVYNuwRgo0g/EtjzBUUvaOPB8njJK4xO2
jnuTL1xIgdPbo0GiCWLl3PjOcifc/Blb9qaHEpNhqYKJgzDbU2wl3ZjAlN178VWL
/2yHV8nBTU5XPiPWoNC5KLmkfR/bqkXgpbM11t70CP9Vn6DzOvzlSrO+Xa7h8GEy
1sqe9jwDsR85GJx0MHsEA2Zc0koPEAsj+6yzOVizAXr0ejP4vUM6K/CNWamhodMH
gxFUyVMgRuiTpUIAQV2f+j3r5hrISCaG0/CqI0UztytmtwAtanJquQius6YdxrJZ
+0Kf0kLCs/DAwsEGr/UvLsq8vf1wGBl0eSjiKjOs/gz2bB23dZytSijUkV53xJHi
gnap/EUr8b/a5S9m+Xk5ujuX86Ry1tqd7cTRP1av3GQKra9UlMedxBNWNYcz0lk3
MfCubxOpdGpHAr01VcgWwJZPTiG2RHkZBI4XggyUSvpn3kHVopSWDupkNgf0/hMH
/jqdgqkE05A6xMMZGo8XawcCEw984gy9ltDTXC1+vSJifL0neoqwoseTW88N1ddO
tLvFXLpetRV0xcU3gRA9fNUNt8FsbPYFmyFyweEFX/4qcFTRrMA6lFLeJcU9zquh
H+6U5ISI96PdR1xofS5fzQULkH1iv4ZjAXpvuTqY7GE54hzj6FXcSWvhfvdhu6YO
Gei6E5TYx6z4zg/oR5C1p2rRmJqBQ46wQVrKzyOhiKSKpfqs7ry2Rl+5f7AxcKz6
RZ2FApTUatq9qZjLKhpRLOrFGmP/Xtz+XEIw4KcB+zVXFFWvom0rYDB0gqC3Y2Sb
vhqxPP0dTX4j+TndOdhrcVu2zOsOrlhp7fvkG1R3EY8zkvX+AmEHCr0AzlR/S0GP
NHDLRgsc0cfS9cH21eNDjMgYY+GH8rCgpDKMRcJgcTX+PTKdjXwcy/H2fZIIPpPM
1rnPIMG5CVHGlpTEgwDpwuw8PM1DODHocnoO/8AwqpPvbAlSi1DfaFdwfD4Cu7Mv
Xp7pZy4CaXsrB3XNwpleAkAUq2JHG6tWAHV278udSpEid0DyXp6BWeGpvbMTp3Hr
2RUBTeEDe3VWEsiJkQd19YJZuBtN1VQ4YgP2GVzEhdFTD7VNVhLHRfkIkFa5IiR3
L2l3DNnR4mxxNvH4L4KkoCArlDsb4ESotqyAo9Sv5HQpXIaqeKzWTJy6AG9npsWm
x3n/LT+uhXNcWjukxaT512948Gg9peOzbBhACsJAB9q+oaMe2VHBR0QmLpePQZ1F
K72KbvNSId/e+ODX0/0+GKL4hz6qlJM5oL57es+1AEfdwSetQyRrH46Ht+e4B1ie
v9+glM/fQENeLn6MCmWODtnb/NreTKcdsqP6ejU44ymiPt5PpeHCOFMXGCNDUCVG
ZrgCtASz7HLSFpUN/woyyzWIjycQ0LgqSMTPrfm1d8f3bLhB1o9wQD16OR23cYuo
Y9OlfgnnyXJUMd77pLpzv6FnbOBPsMTpSr8LDgbmZ0fD6gqjJQA8k5PLmr7Mxnjw
2qItff396kaQBI/atJglECVhkQw1pKe8urk2sATBemE24Nkw8JPneml6NGaYL7T4
iNHbwcPgdstFUdjxF6HAqGJGJaKpAig0Hj27/3P0+QHgwHGxi4OOGrfN8VtNuq3O
ceSRE2m312rRntvOu8GhHBJ5wmUHeNSYfSboZcYSITQ+jnSUS5xXJ7qH+TbmfOAx
NRzTlrownRI/67oqbcIEQKEX7VkbzaGdfB5fvjUz9JwqGUtGThMfkxln5eyo6BHz
BVQpr7fohqkN2WuDnDqykkJ5/tcGIQ+zuIYmKLMDVEuk7DgGI16DrSAEyn+vJKi8
79HYBeYYV2Js0sbLdG0fLa3oInLjJ8ZGncFGHdL5dAyaSbNR+bJ3bewOD7n0QgjG
cAs2QrihadkhpT1hCo5/W4uz/VVca70iJZL2MK02mWYqazfkQsGTDzu58wIe8T7P
93Sr40JZH+ojT0ZZIUSNqPrdonPMPdlG2rLhu1/KcdrUmcwuS3sIzmmzknJcCjY+
I2SePuc55bVo4OllUeRCMtVAiCex81rVSUJlrCV4Sj9lkdDaKS7JN9Pb854ZOPBl
3IsUcLAHrfkqoR7R/5HmLs2sgjv+xDW/Jhvu1giMDLL2SWvukQ/EeQSDY53tsdP1
Bq7Ka8ErUJDWnbZGwQJFne173aVOcXQ4B4F5wXs6rf4YWQ49924YVN38wplaG0os
fDXxfG/Ql52hLpahaZYjM/0Z+PT1+dXz0dCr/PiOdc6R7okI9K5/EpxQYqXvrUJ9
jURDkVmv4jA0iTW3RAOgrYm7D/Q/Ox4fzMNfzS1s7XrtjnyWgVgB49lQO/MHJuTs
JIAR692JYgDNp33U0dhwljCgoj3um/AcnJNRfH+M8QCkevQ1rpB/43r5OOOu7Ure
RVYJL6bkO8s7WFrmiodaGK/KG/jcp/O51UGE7/A6gZEScl3lvW11Xm9urm4dfAXA
646t4CxoHqbaGUYL0KLMQ+mSo5uXq2/4J30qTykfth8kKzSV+Ct7MM9NnmkUbN1z
pBc52HFeJ1AQkm+46z8nXeQAl4pa21mhriRAtgCasdV0EA6ORYy8bHeQgM7KImuC
RN5w44kX8oD6E0cnYlSovLIHzJicjufEhJB8w/lwv7/zRibsJw711x7vCrazHZqL
u0XLVCDEoF3bBhmwb0Ekrgxs/eJeAoSFObcjQb8aIcV0cI772Oxk+Xqq+68BRYiH
mTQdSd+VteleNJ/w/hbyhQ0joA40kx5KwlRtyngp35B56b4v0IQ3uum2IBkzmETB
Y4U3eQWEGdVn9fO2s/vpYr6bKFZaE+iAPg4Mj6v4RYjH56Y5A6c4gZwzI8LH08hk
jTDkD0ICWMs6XlBTv0lOuL3ieb/QHoAYTLRwaj1TGfuicqzTgf93igiUMOC0NVB/
6XS8LcKd6iuyxKeiuLEBwc6aL0QgKwISpl5YBGb0+UKkC39WSzJrX2vMAR4GxqGa
iSnsQ0asHCAMg55wwNhKk59QGAbdCGewK7ewEB/Oz6kv74N/ahKmxFBzHdfU/LI+
7Sri03CREC3LViDC2WiEHVAeq5zJoKl00hVYX6c/vsvRrlqXO9MXteAhn4Q8Wwqr
JTBbB1TvKytxXzZTaTdYmgPAPwqG4R1Roi1XFnyF++8A1XABpI23HrFYN99IVwbJ
+X1dOsohnA/aJpuca4jRiNthrGPAV5F8WwV3XixCUOGrkzMxIh4yX4rAghfwXrwO
Xw0SendBIjQ/JN7auu98cN+LZGFUhIsLb2yORqjanl8Lj20IMQp0MA77Wsu8rnXV
Yw++kloVla92pigjScr+22qlz0b5a3BnHkuKsXM/khC6XVeErpjs+M3L7I+dA6Qj
UEgiHYr5epfLgWlZGybwuPendjFQ2+G4v38Z3MQQw2riEfPZIKg2hURhVnFTx8jN
vtVZ0GwnZnwNeDr4gyoFHZC/50ENlFKy+iE6YRez2Qhyb8c6e2H8emPKyS7YhltH
0DeXFYOpI2BnyIQwcpfLBR3W9s69pjXW+PDQuGLaUkaQC+dIQ5DRR2mAQYLtT9F1
nzOplRwdVO9HyvuocTgAhNf4tg6LV8Pni5Gh2lXL9X1Vwt8sLwQ6Xd4nVkmVEsFh
D0vYWJ5batKRf7W2aAdARbQpvYd2455r41BSmFsH9mnPmRFQTLh09sWKEPlFB43p
fwqH8k010mvDS7sEDKb7b25cXjjxayMjYBZBJxMCLtjPN7pGEo2gAhmKY4E2a1E6
HcCXLBDoeVGI3p8EGT7dgOfKV1TZyov3CGEwkCl+AVBPmD0y7zu8idGUhIFJx2Wk
k2iWTsL5zdWb82IgN7WlnZCT4Mfo/+88Fzu0vvdi1iYzXabVp0E7yKVvkEwpItJf
ry2YEZ9IVmiLdr09GkYDTxqxJW/uPlkcIgsnkYmDR4yH5HT29tF76HznbkgTb9YA
X1Jyo+ydBdD9UhhF4pa7/V/lCg1MrA0zzMJ7a+kqoOqq0EvB6rPWcCP5Lr2c6nrm
jgTsiZ+Qvl4tQxnxaztHAQeEbD5nDPWjuSzMK8dvFKXoWPOBKfFjQi5FooSAlIgr
9HM1ot9OOpu8scHbL2ofbRcu3VZp2R23Mme5S4sy/YatbzyYX0J4qQ75W3UeQ+LH
thA9ySaz5q2v4Zgi1WbYYj8SK0uExyNyiBi3pOdHRjQItciGKwpFhBfxRA2vzU7D
0V4AK01WmBtd5OPTKvkeg7vX5jYxuyRVQoPhSzENOB7+MIcg1YuLS+bbKjCGnegX
K6rR719NbdCa+AjIPzX8hCFeY8qjXyDqF6fnBH5kh+gw5z9Xw+QzR+zw42YGn3me
Q598tt64sZvWxcaYUNp7EfLDRkdovDBOSWezN+cVylNU939MMhriuYYkcA4h8zew
girisd+mIVPv5hMpTYBsr0S0brPyhTbL9wdgqX+ocwCe6sFpdPw1WI7hHuzcR68I
4PSaKrbaKyoTRei/2V2Ar0q4hc4be0BATbV9DQcaHus5Q8DywJn4oDRuS3Oum8MB
HxxdC5QN3sAkL31KkcVhqAdFxZlaHjBZpu6twi4NEgsKMM10PbVG049/mI2PayVr
jdQ5bdE1XavT9/YA8GVPsJNWNTmFiz7xC/0bC28I65+JA7R2YhLCVXNG04sOr4QC
r3Zx83+QUf7ykFQMrsNCg5Mk4+E/oqXoR7hozdguzhHFfgmkqGNBqUSrU6BPffPj
P6nYheKFSI6vLaUPZgvMfcYSQxaaujrTiIjWLf37H0aKP35gUCoIvXxyKgZ0JUWV
cnq93jbw1l96KW9hQa+Yc6PbVA+lxQDsDdB7mHxLYNuHLZOMlPg6v0JPbwrbkLXp
mi6bY5hyxXjZUvD7jBb8lecpPSX1t5Pu0w+9xWSfFlOdVAnwMQYtHM1T5w8SLzQG
rvdcJZlQ8gbgZHtSA8surnQlPUMkvB4k1hS5+aeRHMEahKAxbi9dDFy81W/4G0Ht
Zn0vxiw2BpGSfowb9lFyTYef/KGKulmS9NKJGuF48FZklosPOjMnoPDcFQbdjZEC
qjtz5F5mflwGo8xw1JKPP1KgUKb/bh5fvHcECuN0aLaIYtMxfi8XSAzPc5zujtWB
+gF1i0LjxD0eM6V5u/O+88lzg3G/M1iLITgo+m9X/G4pUFMSbc1Ezp9VzQ0G6nr3
Nm+DHlt4guR5JW7Ggh0pUgrd/nzmElw2UD+o39rucuUTxO+7bFSdQPg6vQcgQtz5
vp5sFdGGrQNdNmmOM7Cn9POne5AvJO8ILhS1QLJhmsPuY7Xs6YS70eauiJwqbwDy
UDLwLGi760LbSk7d7RRNDhMb6f0pH0G0v7RNjvEGOSiSmpV4J8mL7BF2zx2GklgD
0bWT7I1B181o9pMIUkiIfTn1F3x44vnF3N6UoY5grcj2smD+dbWcWoVWvJM6QYEq
J6NjUTLYAtuQqTvcYZluCCQqgm2Kd8K1AiAXyKSiyweNdUxYroL6gUNbE3XxuUio
qVhnJL86QOaAx6PXEgQifwD/O4OwL/mCv9p0637+r79cmg5yk2idu5qqp4CuOmsX
ibjfRcXjwC/CNgbNABy/p7x+ZUSxRWhowl6MKzUKaoU+6VneWFnx1zJeGiC5u5Ye
590djdjIt4Bhvwud4pcOlL5fnCGcdadwsaGzjYbKYHl835H9xzop5Z4Pd3Q3kmSk
3cjHtPXAppO5GJ6k64dao/9Hx8tCh0TxaT653PuH5bsrBebqsEbRNveCWHiIVUDa
/Mk8hXK9CzwN2ixQ+mpjPGw7tiOOMo0OTKosf9F5pWPaIlVWkQON8S7rGBeiSlIo
Raz0cHDyERmxBzDhyh6UikqyZRg3ldZmQlTb4LFdT3KwzDMT3Y9oGz8ODXNCuAaW
+nYb1CYJoCniEouusPZ+3nZLvVy2C+Tv2hVeisu65mcWaYwH+VVNNBeGagdx3Cs9
xIwCfZLyLr3UgKHap5W8Ud/lQwusYs4QmXG0GSlaOsl0p69vU1/UF7ij5uY6xBht
GS4NAK5EXXIiKe4YXZeesLlG5q+qcvs5cPpG8uGiKA6LLgXsqXNW2vuTdkwrm4ib
Yq99Fayo5IRyeH2T495RiE5AaqjWk9R3sjBygk7Q2lybIeBX9Kxf1oWzQMsLOdWW
9VP6FXLcd5+hZ+Xd1kgmNH6z3dd2bLsNb8fFsss4Lqb4ELJWQvkRqlcLp7HgSOUT
Bm8Ftu/ofYD/QSQP/aerDY7mZkF4K8AB9HbF0bOhQ0VVXghWKFLP225zp03OblNS
CCf1l0pult48uN7AuidkrGxyN/AazQZqmVNZ4hkasqLECIhc7Uuo3DfCaOqDDmA1
4QQkHzq3vO0u84bXu+R7Ni0bXoiCPES4o8diCItb9cj476uLyjbnEmYh1T188IuJ
uzLvqMMENe5nJHFyKVAUuwKHy5ZbJ9P2iYSkvWSFcGfU8w+iDcG2tr3XW7QwxJvn
r/7T03hlYp9fnypQ50XInhIfLRBD7O17vf4R+IorpHuZaF9c7Qj0LPAnAzWBm6+h
Xd8jkpDX9OeZpgeCSY1HYdrO7X9IqDzPB2XnmHc+xMRsOoqf9DNeTc0EcUVfCK4z
KcbniX31iFYTxbKHx586uKBywKb9RStmpIX0u4R8q9gBJcMY0QfO9RK1Kffh/v+e
1HnJ+svHCvVrJkqkSRnXZ2OKhETDSIhz4zG5828S9UO9UzvVQ4k78J6CJR3HAnEW
mjw2HIj7fjKD5gvHEZLi0Ve6ZhiZnQ4lZ+Vhlyxb5UJtNMzugKQegr3//WgbGQOr
i14I2DkG+FePnHNo65uyW/rLGqfTdIPn9HoVpCIAMDmXdE2bTBuN3fnTCL+CBguB
aAo6eJ0Er436zcXIVZ5bofSZ0/iWK9By5B5/vG1+pNA2YMG1SeUZ8VmSd14xxSxX
s0F+CCTFiq3aZIlLbEBfyxv5qUO9yR85300uj3DYpkRDdqk8ufw+3L/nkOPbFf/E
tf0PkXE2v8DBCNZbpgLK621jH8u6FvnwIilneWgrCENgpSIosXNy4fqB/I3SHyMC
X7giR+TLUb85MeZq/+xTC3VLNG5KLFh1FBF2i95KnSPurIouWVZpSdJ6+hl+JTLP
MWqcAVmD2ig5AResVFiBSm0tDjpjLisHEk+QevuVqvW8Rbz8/Yg7x/wMaxwxEb0B
UaiGNJYrmp4DWsecKWwuWz1kqDOztxOZjqBi3VgQOWLlzNnqOrw6401nn6WbF2ol
UGookdQVK2eVmxg9RzHeafyw5v7bklP8wGjGGyozxaXgag7Ykvh92BkHZ3esCihN
5WZ9/tFvYqHZLffzu9oMi+1ULkkwbOmOYCHdqu0JYPTn6NAxwRcDbfZD5ldTgH0p
9NvAUX0O/L97BHRgpKpOt2lTOGor9IX5e48N6NLg7Ft42yfLWSpbXkTcRGh1iRMs
Of3y8KYj4CBI0HuCIIbIMby1wWZlOb4sMaR0IaKB4Pog+ogMYJ7hUunf+MZ/SXY8
BiQfodIaGY0/s4A6nC4oEltYf3YOsESp5pGRuYlhakSUHJNnnnSX08FX0lv84bjb
6EedUDf15l5NFryr1qVGGEOupYM8rYrykxMgOXdalpi4oTjkbJ67e6ZtLtKJZk2N
loAgfC+g2vPATuZQO0pfGN6wCZfqCzLBFotCkvmPI8crtYrEKTTk3n5ZEmGMyZ2H
zvyvMWeLQRPDLdFeVts7ww4njHqbi0vvmJroTAmHw1DCzppholi2SScpmwQTEl6V
I+2sj29X020mfeUnKSX4DRLcCN1GWnd4pXIRmwwL6GagF5oeFX5WB0duD9jNz3a5
Sb8sfGM9G6+5l1BAxHg+71A3AVor3cxlGRUfpbjf+wqSENi63IkZju2hF38/cCtY
EBraOVCnDFVsshcG4+JaKeob+meqWOYTwvi+h2HjfUBPnAAUSm7Efx0FVgVbXR0x
rSDTYHuOLHCNJIDfKMp1RrCNq22gBQCIrtj1Zave3G7I6E6AOwLW2iWb5Xulm7bv
/opFkNyz4mXzJsLxAC9rUEIlx7qqhu5uf+f0DOWegz4EYabWwDKkZB2JVnNxTP29
TVtWIShRbDljza/ey0ok0QAvmXsIL+fiLLynFQcx/glSj6rQUL+s8zoDlBotjluP
4eDJJ6sxXa+8Gkf5jRzXMn4USar1G5Q/YVTllSUzJsEDxeVMJOuGTh7/DH+bux/4
xT68pVI2fYs75sLmcK8z6xkuYLueno0TTbtUAfncW64U5bBapu0bxIUnm3RAPrsC
eVcVEZ09vFpoH3VdVrX62TwZ+vfPOCUVACmCq60uLEmaBN1Qm8wAfcDqwRnbB2O4
VjgYuBYNFri5RJiUv0KHERdj8PeFw2LCV/rLju7mQ7bd+izI+j284IRe3ELgTCGt
+D8NlPHORzrmSWE8YFkkVQa9buLvChE0XaYIKNPb9G1HtxSyiAs5rWE/Hfo/SBSK
qudehyhyxtk9vAu9u/cf7jKnWO89qsv8l4DIICp0sq5iyNSi5rPLTi9gBdnJRj76
LSiSqKbfrRBLSA1IA5mwpn/2CfdZP221OFxSsa1ySqqBLwhvnxsTV/+6zWidC6pg
w6lk3nWqw4d2RnDwaeURld+TBVWZQpHUe1Ld2t8l2Q/p+R5XWeG7NIe2PPueszS2
6ZyUjJZZnW7zZAnGrYaA8o7oIhj8KKDZ2qu4oBUeyB3FuGcX1c5tymNVu/R+xAQy
N7eXeMC4G9ItihNSpYIkZmO/nqzgi+YjF4a8X2yPsQDyZtSxR+SQ75ZNgVQCDOl/
EWdQ8fiz3Ca/MTVtPJEdbBGL50OmM7EzR70pJogbetauzNkGGXhWxthlkn2msWDk
0YEa1a+I4GgVMEdQDobcFhDVJqfzWci8UdJiR2BDDChO5JeZW4CtwXCsaQSjYnAr
QL4L61NyjNRczDB2AygEOk199F5iatEUHoe5YqTPhDcfj5JIJVFckI7d2UMo+HK+
isgcEFy34NNwHJ243lHegw3qsQh6NvbbcgnwhDnW1NS6hKsJoDxEbz9zjo21Ppt8
ObZq4sMNjtOB2xBT+qPfl5YB7S6PStFtglWwGAGR7JnE6UsP57YILorgGZiaqmV0
aMgOocnv1KE4vNGgpS0NSY+rRyq8AbeHMgYYxUXM/xRGVlT/xjqDNyDS4sJyZOQx
H5QWeP8vkmJozNgjOmi7ne8TiNtEKtYCx0XpwpIZJgpEoHQjm0kZW9R21PC41RXA
edFumZKGijTOpQCm20wvGbHp08iy2I4WqBp1XSp/Pcwe2JeKpvCW/RON1FbgdGgS
dCzdlN8nKOku6GxLYkgs/kbkZZosIX1PhYNaMtd4QnAYjZ3QDQkpGtHxEXwWmU7k
yaWkxeqq1bxcw/0YAt1pVK1Lekb7FYe5Xue5HiFlGP0RCKL4QPeg2BWKMv1t3LuJ
wmO5pBoPYAhjfFat2Xj1bV5Z2k9NCUvXO+pSdGUqC03y7EVDipLJ1hNHxZCglDfw
D8ptU7BImzvWPfxCvDlF+BXP0ucn7Vdpph9ce1Md+WiUIOPlTAVu5u9LW3d8XuoR
myqSh/Q4/p5IKDkJbpk8jc+NGZqqty39bBaX9pFBuq1EWasHoZEmRNVg9RkSfzYO
p12IJzvDrwbKJd0PM3c9N/XLmeCdHTyJ6tcWD5a/CHjSpKICdEXYRcuizqiqQIJB
MhP5UB87E23rZuJenK8/LHAW57fVTQGiPcVgIqpX30kNP9J0Gdv/v9aO13n83Gaj
bz86ggk7e60nDZ4ThJ3w53+7Lzv4f2fPlfxIyZa/1zXSjDdG0vpKRTNvfrwAsMAg
C75iy+Dn3lPGSIxWMIOr9+JCVYLVj9pnJlStI7B6i/AEfp4/NSqmWfnL1KCStdlo
Uw8DRgoiC1EmewheYT2/7KTyl00+x2BN1NrhzpMBNhBCCTstXf+q1lZf10WJqDkq
Y2ISBCAvjeiNCRDoFpANLhbgoKpncy3OvXE/BoQQC6SYpAMJAi+aLVXYvYsojxZZ
U5OnGE8NJLUbwzh4iBlFGpiIpjUZU9YiLqIERKtDeh2YpAjjah3K40HQmmG6h1vh
TQjCCpsmmgBmS8xV3AGSjfgftJzcHQHS6QogXgCZ55ujp84dRE5bJubLOyRlSx6r
do9mCjvQD0117BI78KH/ny0tTn1jl7jua5gnpfPrhMg8omF6ekcI536dfIUY/lJ2
dyCYPJ/Me0rCVvJK0lkhs61kbq9oJS/uK9PC+gpwCfKZx77Yu768Hs+BQ0SUvaS2
LhPbSHAEzH9ARZGwu5G5A0cmX7kX/wPnHo3qOfbyOd5pG5CrpwxmzzhNH0VszZYX
Fc18jEHA6dIIKCCXn6+3vBu38WgowU04FaR8MemKBdp43nCaGbm3Md4qwKcb/x7h
JJSDKAr9DoYQefF+2IH+D00u9cjIOzingM3rwKZaJabTD061eKDsfuBEpThZ2E/+
TXoX+SjUl+zApWLNsrJh0RjTlI0hB2y00hRHgRlTY2wdWb4C1ysBL5R35iUkR6si
JKGT/e4nGpcBIovJErkSgiRW5EpEI4isfnx0KzLye+fu0YeqRVEYOEjT4ArkhQgH
JkaY6p7k9BbyG5Eq9GkhT0uhDD/KnV9Hm2DpNcx+JOBA3mdD2CP+EZrI0o2uqXOy
0TRLqTN6dNPnzEme00eQm2nZEi0b2aoCNF3qe1IU0XTyc9io3La+oGFHRVlSmXeo
643QsZypjQzLiDBj8RPZj7Irx6wtso46CXblUO7J7dbf1g2NLUL1RRsI9YPqPMNR
FVmgYVjxklegFOrvnJQridATZEWBX7l29hR0OtsX1cnmmt6a5ihCCr5+Q208zsoN
XS9rleJ5ioQlswkfMlfi6vpK7WmdDc468cu3EbUoP767Ivi2zyQEIaJ7WlJVqnbK
Ko1TsbbsLeNkZ07rvGwrkP+zZoo2K+54qRAAUMsdNuyvJbO5+JmpUiWqV4UU1dED
gM3NkqxQuXNnOy6ANeIslBLcxa190mLzZ97DjlxVtScD07w3AAbtIIQXs7/4czEd
wJTQ1HFc4DL2nAta69vUvgdFbccbyo5MGNlMDTrtoWsh1uuMGXeoOFQbv8YEGqCN
+rpUzvivjIj4GVZVPcXqOYXd3nkhRRlpQtLl/lMxkyqMCfxKUuHoLha7/3+tpPAL
PyyGPbM+gzz6YzifMrzbvdIUmrjBSJJpy5bPo9cBBHW+Vac1wi/7qD8w7FxHFIK5
ZVIwmGEprEaQuzZHXz4PtakkGMOdptkh5Cjjq9YGzYIKyq2esOX1CqTHut2Dkviv
pdOj0Z7hppnqorkiJgcQNAgNaDAkwgtiM+e0r7DOY2Po7ElDR/YWGbwixqU4nqs3
BJxd9hQ5TVU6DdcZbGAB/qb57q0suvjHVvY47m/UmwtJYLf2pejTkou3Y7fLs1xT
aVS9rPjPn9HSJPirxRXQKr7ycMLboiwY6qd6iOzPZUR/3Y9UA8vu4G4WT0dMlnxO
43YGuHMwu8bCuz7CE3CYWrdj6zlXiaYN+qACVPI2FlpGn2PtWkg1CpIVLyDCURyq
uSLBklVYDRvxtTHQgNDciaO+QnnU39MFnO/3Qv9VhuOJEJRKY/rYgRkxF4F99lf8
LOf6JB5XFp9fzoXQsMVtXKIqbs7KHT+9HT+F12GAAtxHUyBDwg3bpec5PsnpHik1
g0prYAyi8J8u6uYXwLoIgP0tTGPWxMQv/9ZVWO4+U5o=
`protect END_PROTECTED
