`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHlOr+3uEMA0aXirwpBI90aMUN7l7C036SDmFyVaucBhW+4SLGJ0Qfb28ttgSkkn
FMKe00fp7JuN9IdEucb3hK57cib0MIOeGwE2tpJZJeio4vgxr1OsgrQ4J1yCFkwR
edKL5g6y3sg1z/ZHnA+2Ejio34mYHFbdDIit+v9Vz7ZOiFXT7e4jrqzROJ4KZ2b6
8RMLdrWU+qz+GuGxfVhbMc5skHtHnKrzkAjM+Nt4LF/Ys+PWEPS2Kxyp4OpQVFnq
GV2kQ3BQwk00QdKqPH5/Gqr5r+YpPS4dLStBc5b9agUZHXrIe3KGDeogkrU0yEjj
Cih36Pr/WaJHAavTUEqmmbvdE78/feC0pkxTTzkH8382ZmKn3Sum+CkytxdgY9I5
fnw1MtVTwfUkHA2sk4hdOCiAgnlH899h2BGZUp7dZpKuyI+Ynmpg/Gd+D57W4yb5
sQUTOIsB8yBzfth2JCNc8ORzj2UH7z0qS4RIfv6AAe3baYvsZOKOO2SKuWofxOis
nBhyk8JQTCxah7/GS7DYoWD+YKRdFiQqGp5PG5wAPbsqJmvFrN2BwLLHuylqtoZ9
8NIM1T2sV8l9QomABh3wAGE7M3BZQ7+p/Y2yPmn1uSjYTuPWrXgQWTA1S9ufAs5u
3p6z5kWkl5Wh9Ovf5bqBftuMQ7czYcRaS3gv7kZrfk9PUt8JOq/i8crD8lcfo3zq
6alYZoAx4BAx5rW54KHXHcbpyKKp7DG/Eq0EYrqSUITdB0jAK8dyDppO+UgkxBb2
ZGxkSs2PTtU3nIU10iAcuz9uhGuL2fHdhnmgX7XJA6zHRG+HuWfzxv7jA/2B7t9s
In+Wtk4U3QBJqJFlqiHbW/Mr5Nn65Db5gbTRVaqUwZ3u1dl5/YQnpIjSgHpq/n+G
jmIyKHhDd0PkviftDOKq3hzvsFcKd20N3ypNjaZinK+nv6Rvc8O7G2j5DZ/frvix
w0x/FJG7/HTKQ407V9v7tM+oyNe4NGTZCpi+eFNvEgsCI6ooBRLiVCMz9Dy5KyvE
/cfNofiSgTrLooYKbE7cOYEsxUP7LWP46ifZgLDd61kb+8veSs3hvJd45knCPtD1
KY8j8xHDy6YvBrBRx7ah8DWG2qYTT3z2inAjTfsTubk5zBKfLqtZ8ytk6XNUmpMB
VSbguTk2DQ3dFddLaUi09doKelrNlXE8DkdkY1ek6/hkDrvkJuJl9ttsDfrkavTx
zzMGZHMs/8B6skw9+RqbWJqBBt/8BOYAEIw2lMJ/ofucgSUIIfYuzrEZo6sz0/iO
JCtutyU2ftCI1ftWk/cWH9zQPYFUdVue/R7mmZCSR1e7oYc4hKNiFx3yabPXoMH/
b4bFGCyXPfNAdIZQGCriT8vHll2uvZUHzGIzOZNVRfr9HuixW8dTfjsdZmjMzktp
FEB/9i2mSMOV67vKPPXIrVAfFkWbcDjPxeiKnP0RrsYNDcNKvfiVc7bUNUQr1aEB
i6FmkaiB1NU+fCmNZXXs7ACjEWysJS/rKzs88GBQKiaYmxP5JeHImWC9HQ3nxvAx
S2AuoHZ4Hm2dcCevMGYueKHaM6BbTreIzemhDOM0JhzBApOcJTNbSSEzhXJXIMRI
OH0u0NkWPQ+fxcg8hPBshgt/3qjzOFg5WAHZJoFJphi8afl7VcgzkrnrJpbWqmtM
QQU1wjo0uKWMRKKW/VtRFzL6Ydzc1EuMSlwiF9dND4GevbxFIzud00sek7K5BJT6
vEEWQ9DYxmQcubEBofaJM/JBpevUNAM7uxXxTveMgo2PgQEVBqZgVcMU3fTbEVzd
qtdCx+HxhVaquYYr3dftFdZcEK2UlwY0caAefL/iGTSBmL2gPOfZyzevdWo2a3X6
WKD8kB+ZAiheJvOGFXalrwLWWCDq73BH0rkSa6FRdAvSq1tFp+fnnzJxerPodvBR
6XiU6tl6AYsCakri+KvWmkdH6K/DaKWoEifq4jQzSD+OOXfcWpamgfRAKJanxiSG
yJCEs9Keaa+nqAhmKVzzlxvITyn6dQfrZ/tHNCFaCtGNzbGbRBYp31X+4wbsjRyp
gjItfZHTlUqUpHxiZqfD8mC8JyEcjNutaBOjno6ProUzOQuwJJV2YW+nfuBPFDjv
OCJXCYbPxaxVI7Fv7Nfn5brY24Ycegu1bq8omOSmpJUBF1foEKtL9Bq4d81DIrxo
iqiVo2f8YEq3hV8H6kmA9MoJkktvyyyI5g33KYhIGMYxQUlMrKiTu+jdCB+kHSft
EeQAurNKlT2BHocehRU8DN1D+i/dX7SpTr+WlBxO5/IOwr6ZAQLRfRmOhQnsFr4W
puFsvS9a5WCt1FS0+UVvf/ZoMK96oyWlcznovou9LwyaqT1hmUeiEPNfzJSQghRZ
KFxcJkBZDOqUblJ5rHEoSOdjv78Apcn7rXiHHpTi5NgWWx8LhMQ/R+1M2Nfbzfyi
/p8YOQ4HhQMcwQjoZ9mD0itQFPzQasl3yemJpKuBOh7gqET6VwAypHQRI+HZcy/2
+PAuSICGImMK+HYzxbZ2pegdEY3R+roJYjA+9BH5Vc1iLPjVZnwIuEWE4SKSw6WB
DG7zGgRFeKc/l7d1nhN1t1gQ3hMRlWEcBZsW/PU/N1RyTWlnxnop+MFWhKe4FhB2
bedw3+PuaypjaRkzeTRB2m35DvXMR7NdZDARin1zIjo5CVriPbt/dE3xKulJiBFc
88yYxGesCNuHPIi4rEgbd5XlvN60O8T6yxXRgXgyKHWPwrc9NUkFU+mD8c9gbpda
vIjXygMDxLmtuXoKNF6i7wPGRf3hHITI5/Hmwb2giWpvroaJAXnB/lx+Gd4zcaty
MYTpXXup3nIAKBlc38gp6boQ3uJXk1CzTon8jWw6GpIQub1G6RlSEKalwdwIQ8sF
kw3dtclBZGyrigPjARpn5Ig49mXCpjuWbZzf9/ehNZu7RoB/CdiHkeWe8gyQNuB5
Hu7X8V8/WuKt8Jk3i/1bVUjR+jR8wPuwWH3AuaEGLZ35ZmTtnWfJ9/HppbSIGjVh
OEXg3a5DIvAdO6Zn5wGpdDFhIATEbJUjHE9OlceSGLeFEVjFyho7GkVfMLC76kwx
kaGnYrnW+KciBMrUfQVUdfv/1Yp4ejijsXAsr8ONmtomZUayxfSXj5O16rWWy2tt
hmc81+ZOvdHMvEkbqPnW6YFUaHQ+PGocH0vjuX72hQy07IdmCZHx2rmgT06QM76i
e9xSKFN/PUZepO0HMG3YXI5+K5ONIcgOjBhuvMwykMNlCP1d/6KSI77USgiXPCbw
m2Cr6bmVhu0/mkCo4swx/JBK6BBoYO1r4/KGOVNuupprklja0qGAnMmcIgjMOY93
BuYKec5sQc5HZLrQkfUPm36c3sIMltjxxWy8TBRgu4/S1zkcLLHb+WEYh0SK+YcQ
ILErdTFr/54JUZLZ1sRy+kt3gwrW+gfk+TLHxWYq2TWfnzjUeJ1QZKmhoHrqs74s
EZS35lzXI7qa20Mgz5KZ3RSyc5fi0F59jV5O1BxZCOU0j6ttoC2tVt1JChdcQsef
v52gtaYDlHnqFQ4TnGN/qU82nC6t66Th/oPgGSszrVPxX2R+6C0OetW7r/rge8ve
0Zd4WBeqXAamKOgSIuDg0bQsCImc9FVFgFjeT//9JxTfXDwaL57JYRBn78r3PBZK
flZ09W+02W/6JnAqrn6lAnoKM+mPJKdEHg6+iEooxdnwiLLlA7Oks6nH3KNqXG0A
qg2X696s1YJGviRo+ULz/wCFfy1nUoDvQr1RuIPVoS2IuwfQze+lIRdxUaBWKQsF
XJk35JT29X0QKTO4qhiPwmU2ar586FYlJjzVMicj6Qs1UD3jqCybnBHx4uYhJcM+
s2ategt0Kq/TiJejFrVZQfTuaZQkBpNsHmaAu9Ng8ZufOgz2e5kYInTMMYcWsbK5
1QT4a6hPHbOvXRbB8di63DTg8IftDEKGHyvpq3MsJfEBg4wBh6QJufayaGnZnwE7
hdUOwF5wzrrY6fapSsWkqETwVO+wXzuG4H5FL85VTUDZW9bLb3B+CdtPbzf+WcNw
NRQx6zddQyC0/YErmfooQwCIrbkzRORL3nV5JX3XYb4ptQP490qJwNFc0ZqpTTcO
UPj2qfGlSVGi1G5aF7yLwqwuV7hM3+bfXzPc1KYYNEW88dyz51vrp3AAoPj16l0C
VSeCMd1vzXxqQvANADtyt8Jq6Uy3LBZwn67sGFx/HHsRCXSdaaLjQME6F8Fmq75R
DAoxDAwv3/MLcqS6a9gOWSvSzsu/FKmPPvva6JKnneh0hLkZ5yEEYUXToof8i5FZ
FoOtd5sklZ6HGTvxKCfJyy2O7Jq9u9Lh4iVlGn7RHSi4OXW9oUop1dY/JJBvPOXc
4RZ4nE9192wEaJIzfnP7YhpdonYyXcX87F3Cb4DvFf8rhyVzrJ6LEZkQxKpSpAep
hzwsGHwaGlkP+3h2+WSP5ZnkzTU171e/rguyJjFjgLv6JHLMdcI3jBL7PrKlXpUw
DizZ+HYPp5+9FkVUTnBAdHPg58WJpjGm10MwOr0QtJC6XiczH7E+RM1wTs5jc+Yq
/x7CsQaxX1ayyFqDTYkvJbEAmJtZPJPCSAjcgPVda9OO5HkiilEDkgcM30U66JVr
U69obV7hZ7VWcsQfkpIzkLGAC8v5Ul+Cb3aohT24CtxcS3W6zh5nQPMibewEfepU
8GmVr3GhEIXVjLbUV8dHNOqqCF0EDJCqJYZLR/sABO/jIjsVX4up1xvzDj10mwbI
SZ9FqXyc77ZuJXalFXNkWnKXOHIe8nKHyYEhUyDTqHZHXLUIkXRg/hLDnhrS0I9H
gmAZ7bEUwd2i9+PLWSJa1JYfRy2MBeKMW+M5PhYhVVtnsHnygo/rawC1NV09FWbt
J1lUbCocn+8jN78gh10s7AT9JwUw8sH+OZnutKpF9U2CKqHvJAD90i3qjj2jNf9e
haWSN7uHPl+eTsS9/RsPRZfqNm1B6NVulsZFjnzuo0+WT4WjP0ElAI4EnqqcvID5
sSFJ7lUB1pwEiTtUMc209ylQRFGe98gxAFGewkc8GBN965/2zE4jG0KV66aI46Ew
oy9KciMWjhFZ+4onyr/8n31L6njGxUzH2I1sEX91SBDVCNHp0kEwHlishLtRbKnA
2Ct3OEQgpg/1TnUUerQJNRpwHP+38yUBBfBSUdTiv6QocTYMu+9fGLUZKmwMsVM2
qAexP0n1H6HVsbYSnkHWMtqZy35YEi5YiWvj3sd2e9WF+/J/iMkhk3x8bsJtYqnK
zDEtU+rtiR4ayg29Prfk3puEOr4j+2aaS+T/1vbRUwGRvnP027IMVvnzjGQ5LSUT
Z+Hibbua4+ewwDd2bZjx8V9qczsP3r6uryXdN/IJCZ2rZFWgNpYeltsXfpC3baIi
3/dvo8Lr4aQoRozsh6+5Q56YBoJvfFiI0o6d92M73hfswPTJqYGyzkNfaaP4xlvm
Kju18EjIWyYd3dCzvb+0qpdnIglX9Ikw8Qlj+Qh/IajqtKsZRp3xVoipXFBCO7F7
zH59Rs3AyS9emghmRPHL9GadumxLGRgw4Zuybd0Xg9upDSpb0N8PM/zi/4ks2H5b
D/8gX4Ouh4SXmq7351Kh+ZccTZuslVwyGMvZXL5HwsCXPNzLjvWnk99pzs3KRYi7
7t+r7dxohOo47VFLgMvBKNjui0L2EXl345iREMuJZ+uxt4q5pj8yhkwwEX6R1H4b
b9NQmq2hUVXR/UV6oQkyMCJKFW5xmpGARQHMTaos8wph2qOJaQudk1OCy47N+2ym
wrnRLwNLKspQCuanaHlqXq4F2p4i/aXvYYu65I92pRaNYkXCrVVAT5aJ2w2781Br
ChbIZbrxb6M5+Gi8AflqUs6m+gl2nQUCmAhra9VLT4Co81TALDi47UiQgInf6H5e
2JSCesXXHJFjp1Ge6Y8S+XmXv4qxkVPNQB//Us72pmgjGvUtMmor7SOh4/Nu7ndZ
S8DFxXtnlVaksn73QuyFb0403aWybSmnZpAdaH+RBdQilsGKO2efcicPTWxl1z19
9IkTk95sS4rS7UAVBpDVqtRPpZJYtXpmkugxE0dXpZMn9dk1fNIctroNR3/nhLYr
FzZ+ZGa4iykHuukjGShtAH7+h8qmrqj5ctvLs/EJlUAtrTkf8E18bE2DMVgqtbIy
YGqt4tVmgcy0f4onAn34NiofzMFHBi+arj77vIpDU4tp7QUNdatRxe1CVnf+Diqd
sXDGKv6hRbOiNTG1sZH+9AnERaZ6iNe71iOxDR5jLfmUDLR/dHYqrUn9kmHSVPLw
yq8eB6ybThx0Ce7tIq9f+pXYCvR+s22Fq4FhXhUYvjfoexsN6G/39XWJjcUVDu/S
QsJM4pv/SGODE9F6vZbcvHiWuzXNgP90jlvNJOzovmZRQXknJeexrPInqFtG1h7d
AQpTx8SszVZPsjoD5fj7w8s6MlgHvxt1TnB+Y9ZPpztm2viV/wno9n/AcGaX2qKD
9kqzQmTGbRnLeTBOdhtkhJ4Hn8lYAWYnD5w7mzRRlmSjKpStTUGoKiF3ZuiE8TSM
NT8npiya5i0TYNgefBnOnYeA016+Edp8uT42yD7vJtlZ4pJZhhYROQYdkt1Suz3m
5emFCgA6qwxlarscbzjegRQpfAaSlCAY8sboUVeQrviiEIuSxAlVHEjRCtytnQfj
V3GlIVv0W13W/2maXTHq7FcLBvOk/B2SyJbC7L1klPdAprZZp0aTzrLvyEukpnR+
NRadVebnuUIXPP4nvVN+tej6xHZJIoyJVcyaJLG4HpKK4Pc7GPAZRuV6TEaJYXqR
zD2+mPlGFhg1tnfTU8TrgooEkSPtUhpY7mDhTQ9Stz8p5MkU6GfOubHSfqV+Bb4U
kfJtT/Fvpw+JS9zmq2RZHqD1XC580YlEt3fqo2aQIqBHbONRi9rYnHGbWLOWBECi
bhfuY+P/05o7Ck5uCvQOmgKNszNzc/t67+lwSjh8YGrg5300cSfVHZRkybdtJEsS
xMhGtLmk+2J0ajkqAr2/Fv8U2PXPD0Z6PETC5SndeqL5kRlMeX00aeHSI5FXHYWJ
mfMpPOTNZkRQrBt1OWqSavza6TxSlKfqSi6+U6uLuXWQMPvV1ryDP4RbbPZUwmG3
MAEvb3u2svCcZ64Si+P9Hy2FlzCl3isD6BGoFDHqXIW0vRBdIlNo4x26wYRI+S5Y
FtBVj1mrubWks4ICzdHUmLw0Pz0HQpIMBSFRN2F2EzyxJ1cxB4QuSnWFKeses2o+
L/djPjp/9/M2hYLzFVfePxxaGIjdU68yXd5Ao4AObP8cqyx5TnwrmwukzuUzsaNU
K+Lvg+RVrBax4OgRQ+7iGmbZza5HxBoZ/Za2oTQBWrNQhQyoZqozCsUx3/CSBvVn
iNCexkg1Nq45SRuk6fyiJN6pS8vn4+DLck99x0QjP0hEXQfypOTnR2yC3NF6m6v8
18P+uc7D4TV+rz3OoC5rPMjaaqKfXkwFuzBU4VriGMaflTkxXiIh+1vCxdY+Use5
Grz2wXRFXBZj2sEqlM14tKh7BZT5hp9ns43W60zo6IUgCA6pfKQ0fkbZZaOQCQFe
FW0drXYiT7G0OBAAB28evWK4Mp6v8SOMgeRIXIAIj9ZW873Fkigq3GB313jxrZFn
eaOHDcS6uPVnKseyTHh/YHkVdP0MRa1wNMiAZNuCN984hj1wvYheUHFqwBjFcNEE
ezoyhoDnkS2CjHBEvPCADCbCEDc2nMzhtNyJzH1blvOtd8cYYtf9HPN1Q4clvZAa
+P3gxEVw97B4PASkyXloJ6k5sd6EfsROFg5UY218CH3bRVMdWHBZSUsh3eMTJsVi
ZkU0zUsM2Ti1CsvaCrN2gLsYm57SDDMBZKoPcFMJqGYuqIX2poBqvBLN7IeU9AoU
hGPDl/0JglBEE4WAN40UnweulUPGlb09Plfsg7mKxNAxSMp46M9OQkhtYYaOWhmC
AP6maqXBsPs7vHqza5aZej4IEdxKv00w7AG+8OOfTGEWzlvoIiDEG7QoIilvAsl2
06erLyC4N9ZbonHw6oRUAa8+4fomjBPukVA3KyBSWuLpvSI/FOafLePG1529khtg
nUSnhbGASCfTsZGO1Rcn5FLdJv96fGm7lo0P6OIRAzGAerWq/EmfyWeZgZF2RUiO
etn7l26rmw8u7sb62SLYsLQRz+M25Lk5C4BcLdz4VSyrfrViAmUUplRA6nZ6syaa
J8NvEU7IJaRyycIVRa7G7nyPxa0ubRKpU/6ixePMY77cIwgP1l8xMc2Z7p8H7LUX
46gyrEZRIhvEBkqrd0LjzIZR941hoLxTy/g2qXr47G0Slg/FUMMEEScQP0lVfJiE
/L7E7nWo0mj8AGLI2rmSv6gjuszzHb/5b9Hbt1sAeLHupGYo40c5dRaVEdkkoeqR
eDjvIu2HomKOlXi3jFH7ugVj1Hi+e6gicRgQ1l2UNrceIs6Ce4g0G3gLmzx7UAFe
e/YZyqC3dKcVnhZvhg8NhDwigGNwdJ9US/D3OUyB77Ivdfwswo88hJay7RbTm3oQ
l29Tz7eoTvTw0kzZ4Yo1NgCxzGDyXnY7NxCh1CkTEYD+tQNBZNyCLyOPFYXxWTR/
ra6SphY55TnCSPFgrv42BiXmIdOLDNwY6gv+RBLEgY8tUd4bCXdLhi1IXoh4jgbf
QyggaoEm0Au2tGERsZhPd8LN4fF6qVh2TaTjx/dGIS2oa/1csNCEhtohG1ltolQ8
Hthcj0OCHozUFmcSzjzGfioYv6NHEKrZNyf8PqZtx/Lf66TrpoI9VzQJLfTAquSZ
aFXOYA5SARXrpzepRlFp9MMmW42n7RVjmJyqVAfFzRpftOVaALAvjhgJkN/EHrGf
tYyRJkyU5afBh75QA9lrx7KHB8xYo4wNs77oaIxTwp+ettRtTAGMcOWWnCkEtPFL
CyYUhph+xXCJBoPWDqm8lAZLWU+vJnknPZ4dZZLFUTzA5pVGpAU8zTS8R4yUGpU3
cqSXz07ARuMyG7qs+1fiILMLDOYs/I71jky8lVFp/mYHHuaL6Bq2gr2e8BmBjWZL
jXoH5lPSv0JR5Zp5SymuhuaS+6afDvLJtoT4vi4lH8og2ma6XdA9W+UzAAAriEIg
YUubRR6P6hSohWfYk2UPZV/q1oegme6sraDeP8rY6omLH+jkSMZjQpaGfoq23xyo
biIqWuFvySYqcChRp+xqshnyImi9nAdtQeXqq4GQME86v3dfT2A7VDDTeRt31OJe
MCbYAN7cw8Vwht0xGGhQfv1DDDDzLGzjpPC7HnQ/cZUZxpMItfDthxNrQceTx3wt
Uzw+gx8c3iDaub5WfN3UBqAQ7akmtNRNh8aXJWfYQpPvqJ7r3PpJaT3xO9QnWpjJ
1LfbAj1rMYAWwuwWZUYeYljy9HGtCUVDReM9zcStBsar/wXYvw8O2jyu0NRWiCj8
Z0TBOy9/H3qoV3kKxhsfntV1OWMheRvIDoY7s0Gc9+zQRkZQx7YW9nZ5leqIrX1Z
7d9HHL6CGySqkhKizujpWrYmOTH+HePisQJqkuyhTwb/keFRiordfeKKCvnQaGjt
YuVVvGuCL/MwrA4bMyciBqxN3ScywE947CUWAKa9HRfMPfZKLhs50SgleRPQTCay
mnr+aa07qJL8++3owWlhK4Xktvb7vz2rH++0Wk4YAgbDvnnWJj8Kl/lTylALtVbk
YC4SxiNPtivtjNHvvtVv2eTZa5sAQaoUoNYCrxXkHSzFsvREBS5YGj4fTpLFUuat
+gArrnYI71BOQS27GBKWRAPt0tOyPWYxPdF1jGvPs74NTTV09TQGQY9hBFKMpatV
CCcHG1bUuk0rceqnWjeS/Y9SgR5W252wusx1TgD9NdGH8+Sq2BrkuxlsDFtZMx89
yOOHTS8yCG4fDAlLfmq2q5lQdKPIx+XGZUKz7EXkArFkkzPF1fn4fich7cfSx0ZR
dT8Y7VsCzbiXFo/JoOAi7hFLsM1DNobQO96igCPfqu/hHMeBL0YDzM5H833iPT9H
N7805NndI6wEOqWOVSDVxPUpL2nUvXXqJk+GWRuHYsqfnD2YWteSEbSoKXVJfc1R
rlQy+UNi07JFleYGVHvfgt/g2SfozKeOYcUPMEB7A++SRL/WwANqdPq3NLkl5BMb
bLwyIL+9kzC9oNWKuRWv80lKaKpdOxARAX62WpaEzs3znWM8KdXsTk9KqnEVtXoU
FxmhhwMyWz2+Rl+fORM66Q2wKk8LcD7oN7nYJAJ1T236nxoHS1fb4upEoqrrhgHO
sY6LOGkjxIPGHL+WbrVlYBB8iV1zAIsIYF/ulvsn9qEsWe0vnkWw5V5R+4hLvQsa
Xfnf82I2FYdA8WaN4KH0yJbrE6b/rexvUqjlYcBTJUOxEWnlx+q3rPwo8OQynadT
rsS3O8u7ct8DdpLML9HqMcQVYIdemMTGtxKLgdgiK4us6YZ+2eq9ww58if3uPGVK
gWs24UdY4hdoDyJc6Sc/VWAK8YuKaIBccWA66/mcM/Tkruy331e02WhT1zlCR4if
JWa+aOynDlbF8P6CwVmK9wFEqEBi2hwuJ6ZWXbinkM7YBT2dV/3k/k5kkJNzvtkH
8L4LJ7sztcPFhnzaXDoUSaI1xVWyGWPjYSpulnb8vzYRNkUFXjpeh/qPwrcUIS/u
U/EoS0dh7KxWIhGLtj/crDAtPBJYG7EIPWBqaRRu0TJaVrDNuqRtr20PJAKwZR54
L9NrsJfzNHOwXQONjgDRW4hIuU0tJkqA3QXkRbO11IqaLPH7um2qZ8Z5ZVFQVcqt
owCyoKgDQ1+wb+6Cl105WFeuL8GE/Y+Kn9toOY5qbHuNaFeMNYt3aHurCX6MFKxI
b4GTPoTU2253YFUTuOaia2GB9xvp5p1ZrHW2CE0mbF2TNcsCqALnx8lgbsJAIWfk
piCRFn4f2ao6PiQ9lccB/Ww5+YSIr0GmqH6PbBPfrr/ZnDxItA1nbhQhIQVDqSYm
4cmOyUC5WbLr2uUQQuZembXyBk3hlayWjp/+aoa90OsqILBO1/KRkons2KcKxlER
9RoQJT6jXUODGB2CkSsXZWvzKapoBguUSlRkI51RcxHHW0H3O79ruuRu5l5+jC4a
DZIe+kQhx2H02ADxOu8cpuOTIUQoAT3LxkNgsIDF5uo/QyKLj3rQsnTCfzVOGPkQ
/KrLjCuUeE+fju0K1j6pVcDq16yxAA7WbAmcAYa+n2KPTkASri/g0lxXieDJrXUT
pudcgEpKf9exgE4rkAee0pH95zR/9VHSdBU8CdV5JqsJ8chr0iwckum97iD+ruCI
lIUbc7M7NGKRWS/i/3BQgHiR11JnKdQ180PH1+RpXdjeprHqlOJG/PJi4sL9po6d
XfLBbhIKqv1yqB7hTUV8rvgc+GcJ8/LO8zjibKt/dn5F7pwaA8AXe5oZTN27lSdI
b63ds+4Zpioz4zxgTT9JEwA9G+3KY48jyCt4ECTj7LvQHrLZUEfhSNjMt/D1m8DG
fsZ69wODIRNVC7aitkJA2pMqtWXWOXxrlliIZq+wEiMOuy7oDXl9CnkmV8DA53Qa
ilLQJb1Cqx9M5Wdw1Bxm8aUACwBVvXJmWdgAxdPOw0G4BWEOVnCUgmnQHv4uHBld
kXmtND3KL1vK8bWINS7FL49/KtUQz0kB0KHGzPL+zBiLT12LZaSp2gQ0VQdkSY9y
9sI8whmmQ4ybLBZonsduvhQnDRS5W+iSQMJfs7i3wLD9DcY7yPmTVXltWcMyMwZF
EIN93gLkf4NXjnujAPwj4gUX74FTnVoYPAQAGgFL5z+e2jLU+jhEiDrr6G+zcdg8
jy0JB6WwKmFhF53lFvwFatDpblXfR3hJqZwLGaganjSq7HIadu3KzeBsvOY7NMzu
JQ41UaduXm3Z0GXM2cUYxAP2WYmPXQwH0Eadi6u95AsdoFePxiIbrpWUcSR64bXN
zTPyxrpIKMMh+h3kK4A/voA1sLFtEYjoDTy+Hto5ytuxc71Gm0g24kWQwwF6S4Qu
/FvSBbd57lBu4ZB1fW3ngUe8D3uuW5Cs/R8b00ggUB6E6ZX9ovt1NR0za2qhukR9
MriuEHBfqagWn8RqpdP240EyhvI0MthTe1zKf35hZOIaw/BHlXrfoT4Dlhh+pFDq
IBHV53II5q+RDElnjHMTZDtD1zZiC4NFD4hqjw/3sXbtrT+2awc8XptRpivBinLK
RYMEMNoIcl8XAXHY/j/4/FpeVShEYgOEGBjxWlbBU+MN+08P6HMn20e/5+5lmtBe
c3o3J0ugTCk6ATjBEtqeoYBriDZAlTKqHw9Us6wJlnQg9hK1+SyMbEAGNsVCTG+z
XkLpK9P8xzR+DcqwJh3MOcW7Vc6qgxv9XDo5RlZAqufHJhPqKXYN3g/mxebNqqCP
ACRmDiEj0/zsq7nRzHejJABfknO8kUYUknGW4/yLU3Z3quvGEH5syUlLq3/plqVq
AHXKDGy0fge3wINkq2QdeKyJkYZWNVsd9nN4vWfQnuKKlO1Khr4PrkslmhiRNiXT
8WGiQ+StFuyeqZQviphNCHVTCw8YUZukk4MONDBj8ydH4AxpTuIOi/eTr5o4Lcox
hMXCdAHZ+7LaZwS0QcrZmQSO+fbi2d7lL9r1yOTrlryN3b5YAl9WYhFfg69S5rrh
q9lanlJD+z4lJqmaSsCpTni/5oaM7dK9Kxtdvzg4q7bJJycxrhYocLd8MBAD4FfM
6sXa7BhV33ryTNjz8E9MKepjFIhdFeJM8CzRzHR/4OqA25c+8xc3sPp8iAkzL+Vp
YDvqYuniTtD05uIvqWGr1pODmK+KLA4k4LNpJo8QlglCLQ2YuQbA1rxgq/78rHUH
oB+8iNeRv4jUBzDkTLQD6CCye6zgG/Z3C1VkAI2ggO7Mh0Np/PskntdUaxWlnqHm
uZEwxYMMh4pRktO8Hhylj1wq6SG7Nc0tRIn3ONezop2QoV9ckco5mqGscoiL6IkN
Je2dc9+9FrvAXwN9LwDrkA4LSCl7XQeXU/6v4WJpfqJKhpuo+82ZzZ6sGTmMT84w
haiKdx2cyqw1t010mLNhbJW//Gk9j0FodyhWI74TzZRMKrIwZhQKknlnEjyV+EyN
P4mTCXE3istU+A+Nso4FAzAbwN/SqTxKhCAq6sLZEuXKitd8SvQFvR7NauCBkp3I
IaYROIY6uWD8xnqCgMsPXYAIjAWAb0tQf4BzTx9ac3hgKg4kNbEBzP7CbHDqRxqb
ZCc2YYswvyNnqt8YKxYHDiOsZTCMCbNhosMM2JFRF4hUGB/5NaEjFprHZPw+LePx
m9gecQtQ4lHq3iG7ohr3XyqJvqE5zZUBQAg6ae/y/sw/AqIQk7H5BDfkk2sXFLKG
qQ6/J5QEDquRMYTZG6n9Zuob0Ichn3NSIsFz9yX1PnqeK7SeRXwJCM2PegkysByf
9gNFVWTTXwFbwXRUQFtWdGClxHcpKdOSuXDGK8a6jlNXkDd4cg1JqYEBCqXu8kgp
FsIn0VtrqGMJBXx/+8iWIkGZdimtS6FRjK1z/3cW8BMWAk4tiBUJAwXkHysjCDqW
tqGyjO2CqEVpMyeYGobCPVOB0MLSFUGuxF4W8rjp38cdT5AH8/+Y4WUTQ2ELEYRs
qqbsQ+HCoQiNj5lqHuXnNInuWl+yiWY866X1Dk1Suw08rR/BbOwkZoTowQvtCaNX
Lr5DZsnGDIDogTJDIP5+CiAlbfKEx6c3Kzao1ZGWI6X1imhv75s1BcvZr06RPcB4
uvtN6sAVgzwpxv76qyaVp/e1EskjzcxH0ZJu/uAWmo3KYri+7at1khiaW7d/Tl3T
JaRVEXh2tGt+J7rgQlvDUAfpw46DBCnHXgq0XqzpHff/21ymbNkrcozME1O9rXwd
hST0tQQx45iZC9kfNKuuc+qmV0NGaUdAxTEtkQi3ecuwaoUbRcJYtXkrCwUQF3nr
K5xi9dLgJQ6OJ2ITrY0TtHXDu/P9dYgqIYeVNOiSFDWLGe18TKjKmcMuOk/qa9mO
JbR7X0+65YxwqjvVGaKooktVN82LzmfO1ybKmRNXXYfeVgbCX5VcZIG8C4a/NQ7/
OU+kmIlwcEdBBulAb7U5/iuRUimyLszUyxi1HiL3EtBHV7k+fgeludB1Dtvn3yzz
COW8StL9DEjX8FxBByTr3IJvMmDImHev6RKHLSS06U6/D+4jLcSI7MlSZEYOuHKN
LcJOup85pAb0EgonLVTuQ5+IW2ufiUVjY2McTo8igMZLxhbxvchccBuTX3tHhyLC
WQe9mvdhBbEK2kWyMRKZK/4tbyBU723upAxCcDhG7xm5Cb0f05B305ltVHvi43SC
VfoyfDxC/YAkVJ4CZK1CSFrSKe9N+uSWOhtENytZKVzpyyyEGsPPh670cJuJB4lF
hkJDlUoBx70+EOJsL/YEJytgCs0VxaNdwmF7OeE1ZvRq7M8RpHYpphy7tPc8HmX0
SWhUgr9V93au6wd3WuBTYHq3MM4jnZIveu7ne9hlYT43f0mb8qkkUbPXcr8pdeiB
+BSHBYdpTeYpbh+N4yaVuDu5WhUHj0mBNHhCm7C11JtnjA51kFUkdFbNYeOzx7D1
MuK8Mz4BjQPfymttX7IavxB9tdGzmNk9VNvqNfvZ+jpuEmsQPShqeBNXWiDI//V7
NHbX+e8nOccjhCdJoNAIRYj1dnHIL6RPUryNqDOHX99QkT3QD2JNppTtDTmUIHDn
r5jumDGxgZzkb8eSk2MGgDdQpC+4b0iepukV4oXuJim69TsqdPltPgtVgwVvc4cq
1e9cvHayUY5Sxb9s3Yu705c6ywNChh1rrNeGmsheUzhuZQ19VhshPBrXb8rTTTp3
aHW7G8IE/24DLCr+JfGcpMWskYrEjn7ugmLhhzJxgFIczbtJCxbrMN8cX0qArZxk
VXrb4UXMEBONCh/gcu1JDz+nofn2IVP1Xzss4CPl+3fdDur3zJL0y1nEc7tEU+C8
zlVD+fv19R5fYCgDPgZu8gtgrhSWAHjb5vlEhlEQuq3oQDkEbHvD7ZiGvmole3Wl
zMeIrEN0MkJnh+IpA7Xx/CrGncPj7G/OxH+kOSk4Z7mbtZgFDKdmCMYl8WviubNd
rEvkC/dt9JRatXsm85OVQTSiydABlHBNjAn8T5iyyqiBvmKKb15Kt3z6Is3XFTUF
IGZ739/mgtNupdf0/0Rvuk2iPfrgfDAQqq1iKr1U1o3KNxyXAE43YFLssjNprD2Y
u21IA6hQv20Q6vmBJP7y3Pn3vy6Unis7WDoi5WsbmIMiAp4LNB0nzJ9vIPX+Rvl6
MWAOuQsQsL2NTsvsO/lVA9m3MycZA/XjSgWFsonqGBALctU2X0CHMuPNY2JFG5hO
dza71t8+7uI91JYnT7QI2JLTo2fBnIln0UHAaZjNdmAFejBMkL3+kfdTA4jYmkpy
pMxj3hzPQakAETSLfGNlsH9FRXlUnx1XWCOlYhgIKGKq0XmOdQK8HmEsDVLhy3Dq
34obz6vWa8WHAc3aiskLobhc47TCHNaP/0rE0xYjHfcA5ItWLsM6/9V+hZi+6GKH
2CMP7fRQElO5RKEyBRHGEXoE/urhIPz+92uF8Tn0+nqkYkSigBVhSyBcKydy5Aut
fY5VYobuFArnF635O+OgK8d7JK83m9RVNuuP1kBW73n4bNMmlMUbAKm1wHuWLsib
C0ozTV8nyNTls9e98I9Rf2Zj5+Nfmtcp/J55T/Q4046tLJe2hCQpGIDeDh3UcZ06
9/7FvtXxuyo/n1cmqrhS4F0C24LOtm1UCjwJJ+1zK0FShjqkQf6FsZJgbLeAoShd
nWxaQ/sPhV2oZC+q4biNPRiwcPSDlVBEBdyMAcqUf2ICAUZzF+UrMnbVi221E5tJ
UzVHN0n2U/bcOqZBPeaMzENKt1bGG3kLeOPtjP6VPnCDEujWkb+7Nma0K6/ZwZRN
2AeUjnfwERid1mzj8sjIHc3rWdHvCTaOP/F2Rtc/4w6pB1HvP+F2V/htpLPH/4Ev
MGjcG6DgL6C10zt0KLEqbL5Q/inSfR+mape1uYkFnv64/ozyaFit1Klh2R9ro6ht
5rWXkbsfr8jinAthqs5X1/vdO8gCBZe2M1gaAqPGh4NxoHeh5sHYAgeqes4Cg6JT
r+6+GuXCUTusJJ9MUx0Vws0mBO/awC/38h4+jb4lqXgfggKkjywCtlGR57ZF04J8
/uHpYIHCT8v9MPPxzEJpkFqlILGpQmWNuii4cRVJSE5HSNaGmRrKyLVOCTjFbVh1
HN7mxyqFc2FoPrv7rTdjDKvaIW+Bmq7emeWrHTp1fSQzEw4KokkI8EhAIQlYtCka
eQ/xtrIvJ7Rqi0Lgh9i1bWfqLkRHKtKYOqrsIPLTIsoaompTQVuurAsEq8Ozzfd3
8heEGe/kjf+Y1UUplq6WAWKhU8zt28z4c9Mbk8NGm+2PwM+h5zM2FKTkg6mKtjq7
89GWjlm7p68CZV/SSNvEA3JNMII/t5XA5dFfN0dylYzUgCaOL706MAdX3HSWVfOI
1eaPhY6qgPCWhIR89FQwAcDPeGFNvKgy+KenO0molQyWHJjF8A4CMvU7WtFj6qtw
HlJIFApMxV620Tz2WH/1KbMSw297aemsW1T2XZbQr87XBTYkOEnw13hquSmcqOyt
tbnTTCC2V4diwy8Vu7vfp6s9gl7e7MpMGmsBYQJIVKDYu/nxqTeYxqhvD8RN+8Jj
rKqrO5PR/xR4Z/s1aD2r1xP6ZgmDZyHDoYugTfYtTBShlJG4RbppOLFZOvP8vHEV
Nrice6iTwn/a/MCtp76JVNIVRE0JCB+eZAYs98Cf/1Q6iXatdxag2oh6gK+Mb+Gg
INHvBn70R1ZElusK04tiZAGs7/Ra+oWienfpxb0J0g7xE0A17b5tu433f/PNmg+c
I2zSP8J+MNNxHXCiNIdH7EpE8EyBSbnAEs1qEwB1tqzNOlNqgSFjLXbqG8+CtmeL
Xebpuwk3B/Km4huGKivISC/BYd5eBBAw0Z9blnGF+A6PeUvOncuoYMUQGgr6u8H8
f24ueCZ7GFu/KB22p2m7ZgLkjcipKNwMlnCzqHwlXWUVvQyHGvjmjRf5tRVRC+9t
/11PYg7ZvbJ1xqS61xYwQMMYmEvPlX3eGCQetUyIBUGXOn7u95dYjAjRsA8VioHf
hv+1SePfeJdP2QUNzX40uTIYKKesx9SrE7YXYEqd/M8k/A38G1rdRpp2gWPxAITx
pll63RmLbJF4t+ZvRt5rFzKzdu7uKt5XSgQym3scxa88AVn7c65xAOdZVMPvjqf+
N4NzvsRC8oELtQf2mvPcw9X7TBWiDrKleAkmxgfWyqN0nskFDXV9KkpuYQxXm4jy
kY3UQ8sJMsS2Aeq16TKt7qUSoFZQ3GJkFA8WNAZFoNnx1kawZANjleD4IoN8Hgbi
bGW76cSEC6XD0+KxZvynVt/OPCxmzfqg5qp2lqWm/1+Bm4qDusHFu2xQfLEwsi/w
JodRtvKY6p+5gh0Scsp109J0j/21V0MkB29YC50Mvcr9KLS+PoYPYGHF7G4HRLT4
axx5KcmXoU/Z8hbSH6hBhRn+Cfcka6JxqH60Q8QYjOsyhwk90D8U0YmXQt9hmgAH
WyZYZrKDl/6XZNjV3uXawOjmyBiqSpc8k3WDapqGiiNnM+pjamtLRQ+zynI++h7K
+iTWNn6tRAxNZlFvq1ux/A0uZPz7xgLYicGmO9Vi+he5n+QlTpLyBKznPpCq9JMA
sSM/+ZaTyt2KpggEzT7b3/LXlaVWt0Q6PslycK/BPhKDL+WxFGbOCMPkfQJpiLwB
jz5bumU/EiuUtxjuTQcLoyXDQTli3Bkky9lG/x4hdYXqzrg15bxgAfkePyO/tWSf
sS+aFQe2s5Q6iHqv6s8kLsceVQ5R9jPzUNGXQWtdHUoxNuHbNJ2Ba7mX20Ffn9f6
wv8/hcj5gvdomoWmMAqQIA35ApHjrY5zhJM/5kBDvXqQ+/JMgTFtnFOQwKzcTExy
ZCwG/pdS8byXIg/2BCOrPpy05xWQKJe6RRkqfE9JjlJtWIzzDQPzB2w7tQnRUjn0
qygImtGBqFpa7KYyUlP+xYN8oAWOMDi+jymc1NlCqoBBI+bvosbP215wk4CtArXL
4r6UunVKvf776I5xL8XMvv3eNUKzvPxHeQW0ZH3Qp8289Ipj9XGcTtxYM/c/dtFV
PZsUOO0sC23CxI0XbCoY42IZDuoyFyu6o6W2/E8P4eqDMZzIEzY7AfhWVMgPhtfg
ae/P7OhxLamNcobMqEqhHmoIA8A09RlPh48QtAnfahNgAT2oRmVA0dbEA20OxbBF
q1cjbypefS5O1Z1E5UmqEWv2KacNOpT9Env3pHb/q1eykMfaS0OvVRt+zNs+1epW
kgSo4C/4ycX6U3q/ZlpQUvCiUFbxlziTUdM3YHdzDvWBN2960t9IlsMrkWJWm9AQ
MYorilS55Y/KBDVL00Lz3rnUSQ6X1bw/dRkT0BlXqPTmEet6/zhLXDLAZCP5tlbY
VNG/Y3UkI89jWPLgwzKZZuY4ErfxdyGy7ii7Ertff7A64eIHh5pKp3c/8xQlLRjO
6LYDp31mU10gywdK1E4czjN+a9AnyFZS6gWcoh/i8ZCF7H0GV3JXJbZw6JRAMnhC
cs7avkPz69Li6AilqeUOIFHia5IoIYag1opY4mH0G5HP50V9Tiqi6f6TxB28RUaX
AVfS9LQ6SSV6nWYlV7R87WZQ8TPmgg9Y/Ibp3WGzy/GgHsFemmxv+alhmqMB6d1K
FuKSZhRxa5juuEaNjk1eCrwWn0PFs4LyT7iW2qPE95acWmURfbSE7JDyhP3tSq1h
tLxI+jeslpZWZ9EiAcFVZK1dYjGv1VXEZy8lAtN0+bjXf0AuLJEn76Yg3uBRYiVU
AQmqm6jeqbGCf0DMfPTQRmtKkuztNbRnwe1nDfBwEV6qcJMrdfsblnXX8izaO9RF
Aigcl/VqlREDSZqPEDSZ4D1nA37LIOoUqCjcwH7oLmR36dtdP7D7EC7vuIgkfgCW
gMNRwunQRXb6vLG+NaaHtP4WrtB8UiJbALlmJnyEKKT3oKEUP9gohqCowACzNsGj
8W+/ylNZ5H16CjGufVzrZZ0S+YlIId9YCGM8i/Y3G7/RloP6T5nQaImKvfaOlhNk
Tm/zIn7VHZ0Z+c4/jCpC7G313+KI1CrOdqqvrkOc9wzqqoU4tWX76Ovvxf0qfQXJ
/34uYiQWpWj3JvajZrV9uWNn5iqqbNj0QaR3jLLkC5N/TnOAyj2vBuhgxXb1++rn
GzkVP37UUtOZts/2R/fanZAfXOZdwvtAl15Zbl8Q3k/d/DMyiRQiNlj0/ZIg0jqf
e/Q4D9QB5fTFkvAA+4q013TEs8ygb4ici4lp5I3fiNmuAOcB/CVPNe8R/Zr2SUy/
Op81RVQlW6lpi9MuAI2l+nXuBXc0PHAlZAKOamB62cSaM2DI8kF95xuAvjOkQwcZ
umx/6PED0tBX6Uq6TjYcaLUyKojsbvdJ3Z4NuimC9qzv14sIN9JP35M5m8kWzzmT
M1idyJcOERmf4zXU/FkIS9fmigY2jMPll/E3icTEdzB4nfXzskxuzV/IjRFN3PDX
Aft5rFu7HceoVmHvZ70GNsyyB+LIUDewiUX3KVSvDO+cYIxib20crG9ZOF6Dt+SB
DtlIMGzb9Sln4b3XIbyp6KsRhDXWv9aH9ComMIoAEPEzWTcVcCj1qbxd2xlUlqEn
aUfurPgBsWK/2Ujw0UgEqPm9nUI5phpsKQuNdL5VD2VhCWfDZ3dOa+hndPaqPoV7
fqMszKULwuJD/9BJT93TepDfQk3GykZ8aboJ21Nmm6LuwOvSXdSlkF4fQCYverfe
LC02eC3/vtnzW6zmk1F/ik6pUnnGyNrO5Na/Xe/nn4uqk3EHoTAlqnWGuOfFqgUi
4T6+Gw97gshzheKqq6v74YQtWhvW1orF6PynIJ8tTfXNZw2e5+/N+S4HXbv363Um
OXCBlKcW3PVyLTO2CgMD20yu5a3KkihZ7fvi5wwdtQQpRVNJwYrTZI2bK1HxgfN6
1bmjOeFtJDsPrV8nhzRT8hL32wky8MK0n0HELrOAWj0CtDKVTG8zNju0E7KEmMTE
irRYY9QE5Sb3sKYl2qzzvRsOSGLxu3PxpP6wcb60hVs/9s5KuMWe3nLw9QFvmPeC
7FCFPEPvLT0R1Cjp7V6VE83mIVFC4rzxIaSjKzCmLGdsilF1qb7/geXqOiiifSqp
qS9YRQl6UVouKrNJiNbe7iE3E3pn+NzkhNFlxODue9h2I3kls5Uc07WHpTGcBbv8
`protect END_PROTECTED
