`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knB22OM04i8oFDcaR8xvBNtplebu5iojlGaIu97QIPZE/UZN1uZMtuDw58z3z+lb
s0jgduv/29S6+M4GUxBl0ICl8e6ZbthPMQjUwNJmaLhKk7TKHUSEXSmHjz0Et2p3
9TO6UvXBOartD4J1vvDjDUBpt97KnAxGTJw3c3FtGzNcDDPl3ctPRlJ34OrIzxdG
6bUHOAaNRGBcXK/8kXx3MConoFnBTbCKRqAp7Ikr1iMdKHND5r17hQSHy7nm7t0H
y7excu9A+Gfh8Yh5v/sWxZueU1m+XJ9LeNEK37CZb+wsHBHmyvINRoif5pwBUCLa
kBIS+9r3kxFO5QjhshEUYc50HPP0RXaztVReCoawLk4zoK89f9LNd1GdxiNDFkBu
6jMMKopWnrU4XUCpJZJZ8cCzYYgWv6m/Xr4upjTJhN0/yWFqZ6L9P8/1jjupaiFP
TAjZYwrb/BcrrFXE2uapAl+pOivevSvyXVscYk9KJnxWxiuikXolYo5QaTLHB2rQ
P1iqhMp3lbPpW6X9cl+/nuuDXjWV7kjjGO7UWRQaJbqtatMNubWkx10/cNCWtEFo
tZ9rmCESHe3wmF1j5c1H8cpNBmgCMSBZvD378v7HBw91qmahyylR1N/J/YWIxDGc
uHrTzjC9mjgidTjz9yxQrnDesjhTgu0T987bnTOfOH0LbLwjR2Ld6lqseuPMup4w
qUxoj1ZfqB/hfKoGI19L4gtBBONAs93J3jWVszdPwV85A50z74mhpEMb+Ru4asO3
oD3ycACvbLAEsIAD6cJev8ee9GORIazpO5DUfAEA/8BpS1cqg2no/V0qkxRw3/4e
lr3r1vNtpRxdCCMWeZAZN1FDjvh6r6CxS1/PaDvzRAfzbHGAc89J8sD0wLgjPbHS
wxPspcDm54q4raE9pZ5XlZf8LeCEO7+3E7AAKQ5FK6aZ2Js4oZe/IjgvMDWOxf1Y
auv2vIBk6sgRNQVy7jaCC+i8tE6h8MG6Pqg08xtszXTXnBl3pP42iv0Z5VV486cg
8oT/30ZxJYxM4ak25u1xSYzF/xd/F6gB9kzk/LURq1H5Bjdy89xPPeRL4KJmScAm
yotTEeGljnc7VEVuuQ7TnwB0m6HkpFcGXF21C8UVbCgc94KeQAZQOvaSu2TIRQY5
IqEf0KRuDr2in2JgOgRwk6545CuuRvzQeQxZ9tvON3Z/TvHdmxb0RscGTBjLn99I
vjyb72Ge5KMH2weeOnccwYd/4cups5/p6tshhx8pyKwb4JDegiPi27RSScwl7ULO
L36xptK3FxEKQpZ1TlZRFF+hNXCIA/EUfWvTjTzxC1vpDJdxo5uZ+uIsXnnMaCwo
gOylFyYj6yE0jh4DoLqZpVGFTeDGCz8xRJ9crZZjLsc80PwmiVaZc5QtlsniAVIY
2oEn+K7dvTjOoBOqngjfXyjsogypB20E0DXjXtF3JetpdhqPrCCp0r7dUmtP04+E
d7GKlg3pfY6qoPYP0c4TCjfa27/Xs0JkuJ4wCXvQlWSJ4M+6jqy1INPVJToIL9sh
OoL9h4EAhIK823rd2+36I1HVjLPvs/hLgvmJ4mwMekQHGVf3jIi9vc3qURzTJ+eu
DOPgA9YG+wAPCdsbUe6XFfhg2ERpvY5OeWpk2xlZO0HnPrczOUGoep1fedXrvCaa
dnxE+y1eqjOPXmUNzjUY38lMixg1a27AVoj7thF5Jau8HHyhc9CxgafAJwY3045A
roc5zoEGH45ObIj6j/uE3wi6O5GlkIpTQtf4ZHy66Un+Syd3kGjtcV4iMSts4mRW
gZlD8RWxHo3F+LN8U4ofefem/YuGPzmpHoh7A3v6M00aCZ99X/sAgyr9A5xCbi62
mNSvPUYceEAd3vkot3Np103Fq6YWH7cBRFToKFsyRx8=
`protect END_PROTECTED
