`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NlYY2CcUvTxC8rHjpxDMHkKuxqZCpLdeTjbhYRtpudUn/dsmZ4IhhlJHEVQHcXEh
Pv2UPFDzbuZHs4t7I0mLkn3t/z+R8SyfIj183LAGkoLGiyG/XtOC/mRS726jKZFk
8QBew2vNvRuwRHH+a0VKGjMxtzPhF6DfreUeCW2GMP6N/crBBFSIcxZZ1mG/WLln
uqcYKrJgLrFztk3pd+Dz8lRNfDSz7flffl8nK+A6s7E4payhtxJiZPteYynviNwY
VZcszOTFQYQXjsrh2+jKB2I7D3mWcX75Q2G4xQ0HFwfdHybyTwcZejjTRWid6S9P
nqNJnYHzWSb4Y+5OBVc9Phvq96O1Oqflt2dvjTWBuygU8kZ76NcnYE1LH1idxjjq
`protect END_PROTECTED
