`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9OwShk9TEUrUkrX8qup9DVaUiWWi6nrRYebzkhA1rjCvIlgEmX7hHnNT7SwtDEv
/0P7HPcnZTxSwGDfGtk+RdA9nULelgryxvfFAqi2dO04TQMGnCAeYvOtL1fl1fgo
3eERGhMZJzwis6XkBEIwYsOEy9e12sidXpXzyKVtPAl26+L3QBKwsOM9YzKPdVX8
TmTETwwwa8sGUMkYOS5reItNK2CCftjORQhawkDj7jW/LfqG4dEe6Eptba5rIx4T
LEvcG2uJOo6blAiQPI7nwlvI+wGnysLysAs6v1k2PXPWVjiGNqlpI4AjvoKzZr1C
FTMJY/ZC6biLGRmEEOMxWLjCwRz9aSXG5ttl9yHrZSarE8F3c1K0WH/T30A96sNa
ei10VBKmgfIJJk5QouKRGJiXwDlsih9ISQsJ6DZqivvnb+zfZS1UhIGh49TISXFA
nzL9fI3/vxONiEUxkcekS+eAfWLZYNptAjh7KYnT4Oo1ca5IrjeOcifnTiOeQXTb
XE9SBR5VpcDG8bPuTS+ick1mg8aauO0W09BrppScuul2x2TdP1db6lh8x1vbRyW6
Y3UOo4suzIkIxH54hE/7VE1u1teFQJnjNLbJmaVPNRMfDA65TFgw4uoisIVYbN/9
2rZlNi9N9Il+vx/uhNxXhQ==
`protect END_PROTECTED
