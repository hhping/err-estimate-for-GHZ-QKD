`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKsv/hFqWi7onaEX+VqXbHgBD02KN1uPishZ9iEXbEOVPzT23blM48PjKK/Dk9ox
emFaBNhdat4dFWdU4Oq9qyqW0Z9X/YDlYwCbhcNFcniibPxMtoHZzQH1iXnqPDWb
u8qpUKCCck5WcXeiLlzSQXPgx6lyHzh887HmP2qZm3+a4GA7MwzxmyijhjSLFG0W
cVu/bTcuNN24U4wQNEu7Bs/HK2l8wZOWyyhAfo53boK27Q9tSDLiXKJsIzEuwqn5
VuQ89dZGv6ZLNslAXMECsnZZ1JR3KqHZErJB6GtC37qSqVOeK8J/hsHrxR7NLshv
Gqnsvmvk9bzOmDZqfWwJG4DdzmW8E7+o9tfi3wf08ApiidQmtNJQP1dtlOaHFF/t
EnBzlBmplSdGRl9Yg2FyonB14zkwZWV4ep2I7o4/tqztkjzKtxQLGsJcbDyQi4fj
QEvjENXG1JLTUbayhGg+JR4XHcIjGS7ZQRiUiU4yFbvJy8logvDlej4vw+lXIa1e
Nob8RgwIL2mXfilbyVyTUCEa2qp6iIWKa6HRHJke1Hvgz+n/y8TeFb+E6KJbzQLe
+JGX6KA1rLifJ4kY+CTAabBu/I9jciyMpeZU6qO54BTtBiMsyleV6viYkokxr6kA
xt1AaLWU4ZVljkAZao5D9zyOgSlT5G8b2Dohg5hjg7Z5BSM3ixpxB/pDxlxx0THi
dEwgE8yAVuPedFLmJ5n1+rmdXI+WlZrF2fKsBHGNQKcJEJuA5tcuvrxTvJVsWGVl
dpwlhHZXsw17VPYxr6CjXGijCf09jm0YmYxT8RBQyhLR+kEX86YpCxTuce1/+2z9
Pg/OXQ1zXs5GN7dplgwKp0EvuzTQ09hdDk1bUxQZzNV8Ok80hj44VAaEUR/VyFjE
+mTu7ScUsubmCJmrcoTL3Fzecl5XdblOvrGmoTQZfIo8DE+0pmkBDbbJWKXaSYKs
wyup3YpPQOCzQb9t4lbU+AmaDe1w1/ZV6ovCcxqc2oM3VOLUwNgiK+WOHKPH+IFO
O4ewOAORTojNg3QA1vzhR39x3A+39pERyN3Yk0kpEA3S+pnQGfKRk3jU30GccK+R
MBKvsxVCtUCMHmDOY+cCF/p0iqwcDby456+ZEf1Btoidg2RDb0i+dyJCiCxRzmCt
`protect END_PROTECTED
