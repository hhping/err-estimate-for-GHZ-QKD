`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJZxDzcMblA099X/WlO2n9p7KkwepWHCX5HVBVzn9chfjJ34N3L+b6vR+guvH0Ge
JaKxu24H5X9OIr/xBy3x9tejZAb77wbo7CTveSf+dqDmIw7NN3SpJDThbJS4VBHX
yjQd5pZmupCEg8W8SePf8ItgVNOHxZzluwu65hgwwG69VyUwgah46porC6dw5dhR
WAM6dKb6hdsz8PvlcoD1gx+Q/6eovWyf22054MSnYAZ9MJ2HxqraD/zpxyEX/qGQ
M+9KgDUL/uk0YJPe92UlxRBsRbeBnpjqXItyDxHWswn7y66WAOGb2g0y4vqCVh65
FBwHKv2o3Z4hcdQRXHrPO6TKIZibLIPzCOL3iADJeA6bJnkr23kFF8PiVzNciHHB
0pN7D6dNk9nCURPXKDZ4kXsgHNrKElqJF5WOJIgaCBvS446CB5baU0S3C9BiOqLL
Dar4B9ztcBj7A6YXR8CvseMB9Z8Ax8ZNbtGwnFf8/mu0PHnAnuPDnFZO5DdBWmeJ
CFqaB9sSwUaO1hVHZ0hpPZUKzisSMFdYrM+O4Y2+BrjB8/ii2czeau6V3j3TqhtZ
Sqe5yPxgmvqcsS8ZT6RYZWTtoyZcvUijXnEDiwMIbseXOOyin4lXkAZzBBbHuxV7
IV6BoMUQrAF+FZllma8ATzQD2b2H4Ys9uG4AHxlH1D3WtAzzCyoQyWAXlK94y/d3
7Ya+2k+PY14rwkQaz5FJ/dE3rGcjJ7sX2I4cd5d0AknLPQseDA4TIwYf07aNRhYR
MGTCEgcTd5Mm//mq22TYm/NMusif8GQ1NrfjCnB1sBx6NbfcopOy2GRm7Hclftsi
Dkh2lsIbxuCRJYh6snMQNNxdW/Wcohler2XYNoX4imM=
`protect END_PROTECTED
