`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+Aj4RqNlAh1FEBXqwKMBFLu3FlWR8bD4EylAkwyMqPrkhlmkY0YE5o48qPaSEF+
m0rrc28YhOf/OgOhEybcfi9VhpxSLTk0qA4zKcGaAG7rPPK2F9fguxJCROpNDJWw
S4khYrEoM/IPs9XZD4Hdm02Fss9KJQZ63ReZQO7FpP6eNVwMNN6UQOqeHPhkXOS8
mR4MS2qwzfD3ybbwGpqWX/zts7j8VgenhGof4spkDB1pXf0J8ezU29Bp7VD4NaXS
zRgE7q2EDp5UcXD57qH9R1kBkutXjYcI6AYH9/CTauOzciQA5i3qnZ7TkjJGc6yP
VlEoHabozLbs+C6wMvu7nXO++B46kXGOmcaTMA17kShzhQCryK4I4sdJDAAnHdnR
XSw6RedmjMKcZ41r0DHYJq23wPxLT1o52tlSW4G1ZkEhcm5vP5oCuO0gw8XZ0JZt
V6U7O9GkZnHaMJ0fFlAEHmR3QN2m0JKzWknKM8oaUY35GBiEFcmYFSsqgZw3MOnM
bW8EZotdPnlgZvZztSb0S+QzS2MnETLwITCURRGq6v1HcUE6tm1O+v85VGAIYR0Y
bgbOD+bBbUduJX81OeTk0aQKABXV5l1KfdCRmPHNWSycUn/0V6VhcI8inHQzMzcI
X4JOFuS4Nb0INjoxozED+11APWWJZilbU1niUz6T5IU=
`protect END_PROTECTED
