`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XxfO3yvi9Te/401EEVm64UvGvtFAMEPqCo6oBFnJB2X1xYOXCPBJZPobDamS0wYA
W5O1cSQYMk/jHn7TKkYRG5w37o6tJfOURzHkMNwV7uPfOgCd1UfcSIuvJ5dXJFfF
mda14lKcRKtKU86J33EZL28kvyYZkT4s9FSCB887SfIM5VMFy0zMwgO5Pn89pjIL
CTvRntifm0XE2FcYWEyLef+cQnOQ/5cOj5cEPf4Ats9ZAaYUCLAiNCxtnHrXPk3B
cSfGsz6/fAAVTZd5eaKWOXeeAQs3hvoU+K555aW3gSo/jfVWB8sBg9HDWkt4FSQ5
JYluo6A5WkjfxsEoQEg371RDFra7q4aQp/7C4Q7EBrYAn3g0VKcqueADCm4CkRbi
6riPwfN1x/7w8NuTem6Beawp70eDhGJRmJsxCA016FxjayVZ8HuVod4GHoViQcil
JRbcTChKh/mgR+IG4l1uwgVHdmOuDvesIXsjErAaTaVgmpTWVp7wsVFo9vQA9x2E
HnIl0lV/0SidaABm3d0sBx++M6QjwCMcdgxDqbrtGV6XQZz6n+FPC+xPzD9SgA+G
KeZo0zPwzTNkJxkhGX2uAiahg4zJbHHIGgA08tVWe3ymyS8bJYAN23GLeOTFYm/J
ufJfBZa5JOxuVH476H40mm7gLQpyylhniVEb5i3tycY1mp5jDig/Wy32vudfcNDy
xMEIwtE/dOEOmO0dJv5xtiRXFsTMxopr2t+RjBMVDo2uC7auUD5cOu6zT8KZaQVs
`protect END_PROTECTED
