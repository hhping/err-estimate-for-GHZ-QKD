`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCAOIIw9eRXksf3FARG9ts4nZE+g5zNxzeO4xQEvcdDlUsGKuIzM0SkOHX1PHsA2
TM8dTuQ0PcGqASCDp/XqJrrw6/JRdDActebgV5LenKP+Yy+qBR3V8nOIJWc9t2Lw
kawKnvlgkthBbMyzN3cNr7q6F12ETPksTxEvNx/clHlhCWtCBDUz6fB8ZPRVzLPj
zlLrBMvd73tXGzeB+Z9NZGybMIVlYO3X3LNWrxmYWrTcWdUY+zMfOFlt/nRbSxSG
GUwq0acZeg+XdVWYQNzQrvCcznrVMCrZWx4PIbFQvl6jBafVYy7ZDhs6+QSmI/EF
F3mIS7JpgUE8cgObnQiXFdpzfEenl1pghqXgKu+lvbEYqDA7Y6EdG4Z8rWYw5Xh0
tJVjGYeBBQ0z9Wxs2NSZ4Qj3S8pquKIAsFEAxDRw4a/P9K0Kn0YxZNnsHe0Njgf7
bsl7HJ7+iv50sJAVgNWSs0KiMN5a2RVY+5QNSf9Abd39rQjtSchhNpMuKR85h437
IXuUFwcUEE4odjsrGNUS5hRDbm3JSMVQNfaWKL+UA9YrXDwOZLW0XIFWoKUZ+79R
fPlH5uA2MLGij0af4I1mCICffA7XqydAGkqAv1zUHWc1icnqpm0njJRGS0XjRH3I
Awn6WVe2n7Q5W8grLqvgwrhq3JNcvtmrX4QlmVhJtos7BAA0RbiaJhX2xHf7XkgL
0fPYwaFmLfAJUdkjgBNiqpaBykOzA+Eh3pV9G7o+/7YoCV+H95HL+ZeU7wZQfZk8
HQ2hwLGqEon9ngCQDHLkGuo2ltown4mpTuHblu9faxfjeBhy8TRgnKiiQzLSP4nA
5wHx9iqnCXXFcPUAffhvV0zCLh21XMGSebH4Nxu41cv9g/RPesL4JeShE39T9HpO
j0/aoZ793tQCf+iNCGmlwZ9Y11ogdWW4UA0JzLvGKL9kPfJSoPsMfnk0O0S3STDP
m06mUFkGrau0H/LqJMneEuUai6klXic3U0m0RC4LL81m6oGQWGwNtCfQhq79XheI
w7tgIx0T1jdSL9Zk7zqGryLSe6hDWPjcorrJ2tSpUVauISkJVR+XVvdcY0RhaODx
wD/Xcj360OknDKQcgx8vqur8t0CyQPUgMdO6HqB6pASG/igEwcGnjAwajqhTr5Q7
ZFxbO5L8qQkPz41q+5q2VVJtWlUFXnNp0zGrd8tfrp132GWyo5mWRy3c0jTXRG+9
P4zYf8pWIiez4hPHm5tQEyh8u7x5cwNGrFLhSTyLoxBSMw5dUJJpQZDo4xV1KBuf
4NqaQeveS4jNeHahK0PQRIsgB7TxmBqngbAn6ZE6NKPQs02xG+4TQOw0OP7MG5kT
JApM+9QDwUFOjw/DTeOfIIPykOKGzc8VoG/vlt+SlSE8+H2rxK3UGVSMSQf2Hr6Z
R8KCTVGirNdambiLyLZEtAwWi5amDPSEUUESCRPQtGDq20gPlFxtsowhFHtBF+cH
vJAADZ9mdC5nEWJK2dop4PN5eiQd/8F/DIFod7+dxOqg9T7JmH3FqWb22zSyLr+1
yh0z8gQRUvuDck6NDFmuDrY7X6vtpF5wlvSSh7XcD0MpBlF1uK+jMvGQfVkZY1cU
9iAFA/BCKqTg0rYu0M4F3Nf8i0jAaXAnSYT3DQurNjkPOKyh4Wv0aLgjMtqNESxT
0gRwbSz7WZRHqB9ACpKsld4pghJDUwE2yLbrt4nx5Dl4WGwVzVwxIGa/Mri3W0UA
toOqdlUNDLO7UL4O6Mp1TN182yHY9DVtTlFXXnBaV2isS9Sc05HwsD2NS+E6L7L2
ETULZ7k5dINKwIztbN0IjUB4mXsuSn8CQIF5dSmUA9Cpnqdbw1CogiJhUgLN/yV6
glZgbaUTR/YLVT/Vi7pYeJE/yDQkevTp1un2IOsCCKnTQtUk6fsebQsTFdYHPhye
N5nReKOdRx0tlMMeljdjfNrBNhKE0+GK6yP73Gri+sT0XgeEwER3ZTGQa7yxqvPf
wqGKMvpDfJyAekKYx+SGkoyVXf5X8RIUxOeCJxGHjDusZjatD2ry9I/kKF3/siMv
WFPhOYDsWxbzIouOy3EgC3rjbd7FMF4EnNP937qtqwlNvj1GuFwKmrB1pA/9GxuB
x+8EMRrPkPFD1r+DJPu7L4uHwaGNFp93fakQQwJU072UTySyZGtmW8jmqcw/fOEG
91fs9XxmgvfP1BZZe6b4KTQ0SObllPc6Ymbg8AImJaT2Loyr0FHxIX8nHc8EMDKf
KcUX7K7Q/fcMtCK7PqSGrp+90+DCUdXSEMjh3XQaP/Mg9xF9mepIC1n37i/l8ue8
12ajy1HK3ua0Q2FyFoqnv0rAIadf9DRgRz6gUFdCMCoPzRji7yqvYR1zvtglVSSv
hXT+H/jCmrFWZgfoMt/MXwNR29JkP/3GAHVeMUl5cjYkSoJt+unJQHkjtsOHsagy
cFzFnmRrxqN+Rva58jVR648JD6nnBG72MzHLiP/Mbf0W1jCOVtGOPf6MbwNHkuNF
xG5hOOlL4rJ4pd3Gyza9eI3IBLJx2tp2fvPaeBWB1BPqdlAUHySDvS3qrxm5t2mY
T/GhYK/n8xHobhVfChP4wT0RWnewAvV7/8doFi1UInJYZkuwSwxRNGXqYBXJrX/h
saA1Gbjlh2+50Uei7dcFTpD+P9YOmiuHl2/rTOsVZB1CHiTJwfULaNaIfxm4e2hg
KNs1aQOxNqioS3e2HhJuMg==
`protect END_PROTECTED
