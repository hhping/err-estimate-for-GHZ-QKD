`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndQ3cRKG2flwcXlUBbKwlFtTROjZwQpCRIfuxZp0BIjs+X9OZQIo75hnf20Vn5Zt
FRXsobLCMosfxHOldckylMpS592ni6ziKAwkF5E2w4PtBDEifKDaaCtLFVh6Nxs7
q1OYgIvOnDK30TY55Oodhi09M8L+Ta2f86gyqwUFwSm+LLcw5B/gAnh3s/3/C2y6
3gR/Cf6uQiqBNW1k9Jb/YjNxOP2+Bo+2GbJP7Tjle5c/zMsq3Izefqb5W3y+39fQ
PrT+wKYKDoQ73PBhAHSIsTihFUVEggCtMAZSYoH4xCwofGHotquUZPXjRu37bNXe
p0DrbZKKET3P+MDIkxI6AfQJVlsUIYJ9Zsnc11boGqNYM0dkDHCIXPW4T3oCqZlq
+6ylUpJB/NVEtQe6oU26I+6epuopZNaZ47EVSrrFQCFeryZ87U3/fQzJ/sZM9HPM
bs6HRfldu2lRJyjfGVRg9LWoUKQHCOnWs2NWrqcO8kiuJWtAC0HI0KqPiwewPp/A
O2P61PfcREKSisJWbxW9RdCldiMPDuAXwMh+tnEXV5UYgZ7TftVUmKhO27lWCLQA
eM5MOmcTjKn5K6O9TNBuRKcNaHgvxA/vFmAgeqqZtlLzvVhOcOSeUc7LfsxQZwZV
8kJb3SrBpAYVV2NatpInmPW10NRgCZkK5tlzGQUBcjF+W4Bc7tkuu9bM7yv6XiH/
w3Pzl5tTV9uVXvgDOJ5+NWyw3piDZqnfteE2w95mZb+DJI6m3KWHsSJ1yDitDy4W
4/tQL3uHzAp6thqsJNLAgeHfgTGs3Ek3EEpUtabwBxls2YhDp1BFi+/aMHUiZqVZ
D9qeLyKo5dMQNVLMOMQVxhaebNmIjkQ0h5vcOTsDLA/cGVkW6YaCtomzB9QvEe4L
iFsPLRnAsG5Z3piFZaixE9KbdL7Vyx1SJYt4dHfqfCJmM0d54T6bNOWwz4WFo7+6
jFxcDJMNEX6rn4nXSlTTF1uj1p5yS8c+V4hMrQfknFcMUbq1WG7WloIUAGJFKxb5
8Ce/DhSIvVxTEE4pfrqCJuLe2IdBZhyuZeN+PhrRm5GciBBnUzBl6N8Di3Tn0EsR
KmnRqhgyNGBt3j0MvFNkt6PmIh9U5rjAWv6YrB3Y4JOY2qhpDHylt0R30UrhGxaK
sEuJm+OhLQJiFH+eQoQI4e5gXhOeo9Txx2re4YnecGkGQe8hB2zHZ+JBtoo3zZnN
zRrG5mQ17+lvZ4lXDIXKIFlEr19HxDEUQnhSOBwvQ9olmtCpYVrWhWQ5eg+EdE8t
mzeRJQpvlydcBI/7Tuc/ER4er+p+hVvCE5tR6wQigfxr6UWETYuYvOMBkxxIv3k1
gsfy8F4dYEjgT2m+fjBmznqMRAFmbHDZLqP1NXiy0EkNHeI7lQFtfazYdGwkfsF2
izUjHcFHHjWZweSDokLzcyoeJlhwCO9l6yb9HMPblKqpZeg8NM81xPs3VEflinU8
ojsSg3D1aQ1gxjjyRU8WPWTBAOsBKAstvZCXsCM0XqkTnAOahtuetrqioDcKJ9fL
rogBWjPtSB+O+nW/RMASA6d2bVmIsyDT/e7kAG8j75ctUg+nwfLiClAwPSfskRe4
cHA6hvzR1oV30KkpPg52Gg==
`protect END_PROTECTED
