`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wp+WNSECCs/N/NMp8iNZxXWtqTqWp7r84XNAc8nmD41Ds4w7/LNJ+ZTCmOFjM4I1
6bM/WWY6UeUg+B5uMlYzkPDftMPm2BfR6K62OFL1LCTdJkGiWajrtzJDchqA2xmX
YzWCrNjYURaBlVN91tTOB44GDdQ3XR3szj5qgVnnoJT+xogoKQPoC53OiWtiIY8e
nxeNepfx287yK9cS1Dr7ARQo3PJTIu50pCLqyTmQK5Exmwrz8wSsexMdhjj+LSvL
3LsjgyMT4tW6DHgL+f+1MXHdCcBHiX6087V4jwJLGo6VCYzXM9SYrHHLV7+bFb5Y
pgJqc8E1Mr4DL2FTXlkUeubIk3Cu4uubq6dWPc1mjLLfY3sS0+r083h9S2cvojYB
6RlgGnz/hffVaaTJHOTANKHh6ZlyT6ZbWcy39TB4TW0meZp5ZRk1JFZHsa0ImqbA
pX4rr+OxgmuhWjc5JaRm8xzRCHyRGdom4cUbYiYRNvoc/sPva25b8D7/kL0RRpCJ
L/WKcDja4hWR7cvhiFU1MqB03KhggTMFDM7cI353Mw0SnfRDoeL8Asl5DnJoUTOW
qjxBnE4Wj5sHfzPZ8xFmcic1Vj/IGEPsR5WpgeDp/KbW9mrt1Xai+KkF4WLbzUR+
aDBuY5CC7twraNDNPe27v1QF119VmL+Bb00BgODJSqSNNZOG551w7r2ssD/zB/xy
ZCtG69nIXzYathscm9v5ne1+2uJhvt7P7BIZTZfisBa+97hGShcMFBtBjQRiPaHj
7Deq86x5N0yvZpE+m3tMdy0kmJqERPnN7wJ+ovRuhiM=
`protect END_PROTECTED
