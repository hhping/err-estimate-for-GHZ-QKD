`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lA98z+a0jVLMDk7nROCC4etRIAphE41qnSMDT1ttIZIIqSpLCN2CGR50cQrEQjrp
Fwr+JPy8fmfG2q08R42OKN45EMywNIMlOgJ/aQHzst/3zdZiJejJV6KXlWbhdMmi
PH24DmTQ2VcD/Unwey9vi4Z7wz+CCe/mG4KwuZ4R4//2hbc/+jQunUYzMEoi/dut
SdbSOkTv4Esq3DV1u55r305zMc+/YqqAMaSPeNV+FcxNk8B0lGp5RpWQb73NfVsq
8VDAPoT34BYd27boj/33pGXINGcUGUNt7uJOTrnniXQYFy8yldkY3FCVqcWhSDXO
M6Z+FMshW2a7FwiB13oZaBqvCCKLwYEbFg7H946vffrxHggnB5ATn4nRqRAxzGbw
HFLejInA/FBXZzYRyd1zMnAegeWutz9WCioD6g+ITv0t66+S0GE3hkoDlcxXGqfz
5sgyLsME1p7Wz/x3mzkRVz/YjpJ+zjKjqFx9MdM6KolbvrneZ+7/PB8Nvy6pUiGQ
9dsD8ByAT61Jwlc4Rm+BpwPd6aYG6MupUmtcRlTTcBT57qCbKABRaj3qbO/TBpuT
pnK+37wEMY4uBwM1y6A4EarQskcbRI8IeFUZHgKvjk/iECSjD9MUg9pN3edQFrXW
JYAKJV15pbdxWy4JRAxkZnRO7ao0K/VYoX91MxlWCt81PIRKkeFMFuZS49AtjJoM
HTsXFo0KgOMOLIyyZuMXmMBXU8RoU4jIkCkBqVc/tMZU/7l3TIHu9bNFc60Xy81L
TRlnjWhwOVHRMAqt2cl6rn32J5en687b3GuSfYyTrHkIX8MslfpAlKyVfQQvKGjV
hcPrLLtJUEStvfug/+8/mWVeA4Naz2Dp4Hcnz07WqQangQ/TYms6lTaTi5n2HtAZ
A93xArIEy45faA7QrdI62VyGmc29825lrZcyA1kHrO4qLUUJf73XQoa8CBowWQsP
YcWmCc5aLvyh5cVVjz4wqTT5M4iRuc5e3+R5OZFRbxplolJ3EvBt9w3aRLra4jDw
1f+Y0hv+2Djxr/pkyHUQTndxXHJyjivLPpmUNKDthggFi7bcLRNUuaTmmA8r281M
OFegRteTgj+YQcyurF5fKyFAd639Mrngzd4XSfXClyrBrzkJK1+jmOTn+Qv4/AKS
Fh2VSxEIkZ4qcHCs+3L1fQ8q3yRqkXFN3HgRC7pQrOVlUuGa4ODL35KYshbKxQZK
prXaXxf75ADwUr9ELnc8jhtXiBUu8mbiSB5PiyONLLzY4mTl2Gdvxz+YmuupK08c
/PbJHCYD1hEZuBU4/Yq8dv+FrWTEjq5rPsCe+ld9nq31j6fYnY45U6BLXkaGRQ2d
/I5nX0guxW+9lL+LmlbG71BNXN8/IZhLO+leMIB+3ygFxSqQUS9qovIEB6wFJ0rK
L2SGTIIWvjIC9Gsw2Rde0h9FlYoPSh3nrViAFnWd30yIP9KtKocZwBljVY3PzEJG
V59d2H4955nI2SYSlH3/O8VCHkxEJLlzetBCPLz72PewuDRNhu5DV2g9ZrOTTFKp
fNPQB77IErFys75pYxFG0Q==
`protect END_PROTECTED
