`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzJ4q307URbx0MC+90c0rfuQWH4V4zWgVuyPAQBeV2p+uSej2sRFiYcs8+/HrXkd
x3MjRu/H7hu48mabGEmMpw/PTdXomEj2+69bzm4D9RVqkC3n985hAXHWoDjX6KW8
mViV+iaYZrM3n/aHjvgl/TErlfFrNitVWiiIdF4kpKIbIOKIDdLlChX8lX/ckM91
9kP4AexWWjYrk7gEIcNlaKGEEUOVfQWb1sZ9tvHsB0K4CYqE7Js8spEdjIgOKNrk
2S1aQ25hjHO8fGTqszCsdOvgAmMYxfbIWCQwEvqIgek6rvgvxfZSFu4he5F/+cge
7DbtP4fbwky+RlRt4e5zlDVVGsDiGOTmgupWFKjAvJcIPRSntozml9cWWoGimROj
PIjt3Ar6jCTxNv3tU23ZnYsovYI8o/kvZtWuQQ2EfxOIfl4daWtmir75qMeo0pdo
7mEoPv604BCZKGtkd2i3L0nI2ZCbksONM/A2JW3N2u9Y7/tkhBWy4H8H5C/AHUBe
gBar0xOeG58koeGfCzE8Qj8+sLy2pINaEuHuDNpMEvOFb0K0TsVW4EXIEIE0gTqm
NNZ91bbcGESBR96o702H+9y1DMWrRkwTZxxf9zVv4/4v3rNoMfIapLvEBAiasrn/
5MOYK44FpoWtaYx2pCU1RB0NzRij8fXsptKIFKq+Z3pQt1qi/JR8EU+ylL/Y0GZ0
tG5e+0jT+N9Gg3i3wJJ9/4wnqkcFyXy9ui4qneEyD51xVL5lf/DveMiKo6Mi5vlk
lTL3CKqAiDkY4VJXeWABAWRuTxE24JgdAkHl5tWLNKE1J2jVZ5v7kjBXQy0nNfII
nh5Sj/zfPm45xQNxZeODDmEfyzesWgO1kqlBHiJueqU1SKTEkSkkk1HCR38K36NS
5zQu5ThEmSfmhYhB7VeBbSRSpAn8ragUczgnObpbqtqSeBDiroRiDZdPF0kluV0J
lsHhHbQlXZJcp2EfNjJD23sdOfyRFYl0SAHMlKvL/3svQQqr9EZqyy/+sHYVzgfc
ICiUwcmPu2pm42P78QaAV8M8N4zVVj/Ha1nmWnezUabyt5jwZbh1SvBr3ItU9akd
YhDYpe92v/fIL8BAvsdTivUYLRxOwu5tgxPrDM4GfS8vepdd6LbGSuw4Qy+5w/zo
TvjCiPQGv3nQTWZfTrLkLOddtIhaFbRDRCW0Bt8D2RTR8VdgHdHRMqMkxlaBpmGV
SgNXNGIOOqRphIOfffau4vI5Qsxax5jcaoA/2ULZny9azKwCMPDF+ki2zcOZQs01
3m3eJXeHgw3EtsI/BCsLrA10qIDMuJb34RsfsajcSx2PVO/JQpyL6b0C9KT+YNfG
AXlrg3JYnHqER+JUpuq3dJ6Q+M4+rjCJkFm0h2R8uM/jsFC8RdUZfm8PSm/0zd4m
6/R6qd2IQlANlJuM+yidGqx+acmDGhm3sS6FWmUFjf+WBa45zu1cEXitBLrBdot1
BczGg2Bc6FoqkKba1vgu/GK+1GPvACFSIsRQk2wfUsVCYJvt9wBBbGYp0v+EYKbN
3cKvEi1RqhUP6tM8IghqXSsLAnNiBbZf/ghx4qWgIy9I4wUU0UBlJKSZSTg9It5Q
kU49aEmnLtTI8iSy4Cw1dDgiPONIGfi8pX9P5AVVucGVhKUePBgJXumXtgMwsRS/
ywBZ5l3tYuYu5ZLk+KowHQTCEoGYNZsyIaBT4xHp9L1hzK4a7HLsYyH5cS9QiUK4
geLcU8dEk9IXg/3iDVPeHfbmtLioifs9ZqQzGVE34/8dckCXffTDtlhT9+KVfkHJ
95zaFp29PzScvW2DoyWEDc1RIuKv92pwIexRjz6ua0AYlpfLUfaAWGf5hv8V0W39
BupOpgfO1bUjGlY3Tb3W6VXIC9nA6+35eZa5WAlC61vAwXh7sYZK3fVTxMHj6t0R
hJKTfSxX4YYyT9nEPc3ojQufWLOIRfYpIoOZ8FaOSJfZ7iK3aGhUwHlUw5+Nr2pW
Uo5O99sKiqkQHvQDq2/XP+YuoaWaGVXJKJJw/aI2xlvGRffXhh5NB7ybxHME8ATg
szCkSSrrF0lYWqfnO1Ygy+MjQRoX9DnGKD0WSkOQwBCvt0xmbkm63o7ulz+vfbMa
DFN25LGsd83QU1d3yNEUFOVdgVMLNJd/ftolDUkiPFU/jhBVkF35Tpxz5EgjDY+/
V+eUxYfJ/uO5mHDkEJJXnRi/06YKlhYkaxgwj/ONyFhef8oaFL1wgEP61LZV+1X7
NS4QkqAv/VU/44N5kDyg5CEOLUmkxFTrIfiHMq3wppW11lVBadHE4O7eFPWN7XrI
ycDVMDLTIQF0XgVB68UIPgz0KAFNmbLP0rVPMKNYtLgatWmGpztROpwHimItHNZO
hPYeq9jeENhb0S8IsnGK1vrdA4ZO+f/c1xFVqJUchqAz/PMxZNh5d1Q0W+RgAdZS
/S7uZjP2uce4rWS6UMXQB5lDloLuENnbskgQ0iDL7NJ4E09WI8FWyL1W/nzZa3zu
c6MaU9D5SE2YSFjGWVqyhLi2sUYUzPMGLgM7q9nWpydVOybzxeHPy1UnVgKEUu4F
dj1TQeFZaiDESWrvi/qmrKbyrvwa20ghAhQA+FCxjKC+GtesItXvsoMMsPWkB/m+
NWT0z38eQF1yU9bwPz31Cns0esL4b7214LwrTxHtxuQjwuBD6ENF9wEKspKkDWNZ
HuX5FUv9PVb4dOFhCAiLD6Iiw7mDt15jPc2uJDfSDIhCPeiXKer9Tn9+VIWaMxHu
TRaXYtBRps5Ji5/cObl08XiVXfNj5A58dsCpjyaNcnPzqaKYlxN8mjTwdNJ+dBUU
Q9p3ByARw51Rnn725Jl8U5Y3Hm2doVWfP0HU+Cv1qIbJxsnLVZhpLHGT/4mFA6X1
fU3OOfkWwWcORmj+NPYSXnz5SlfwlU8VQHNzU611vQdmhmUass3WD7rA3Yyr8bCp
a19Hb9S+xWrRfS5orwwtbhTklTOygW+n7PLp8tAwnoHPvzf10e0pjY2Kb/X3T6Be
fPw3jTWkQqq8GIGJ+rzX6XORoFdEm13jZhsq2FsrOQjnqCT3U7MChbhB037pjXFE
0H0h6ex9CU14rTxru4yzN1/OyBuvF3XFyVnAlEAPrUEcSBqC121baJLt693K9NFu
N5IvYGuqr0mapCN0dujNzgQhP8AjSlB3GKmpxwnqkk31HefeODo3rysajQO/G6ak
P2d79l9ljerTJXBrDFXTVYl0CpCXzrhrQg+s0W2OLZwoVr4Q3lwnghPC86QKYi8g
bSbB3ibnOKUgQfU8K89LCSv/lXy/iPDrT4c92gLAhx/mD4okfCnHDzA6d0ZEMDZQ
USCO55ioMBws8r9rf2P5zIDC8JDaZRWSoY1p8nCwuqWHnXlx2kXfe6fSs54LWz9H
tVnOlaJy0JmnUd1jZKRr104ppIX0dovB0AskAfm1WjFPGxc7PP9Nw2wYDtrGyVqB
TnGtUGzGMazvWyjYqBcneYaZMK4A9SGNF9LgMhJpHbgHv8tRju24QcUDICVC0lx5
hyH2hQk/1Lg6L0VRy+DRHzym8zpKsxjkjYeonhz/CG80pXW7M86xBVNRq/fPjHzU
KS6+LOX8zGHhojz0UJCwLhI9ZjUoq0vZcSC6ZJSb0EHt3CDzfJnocXUhEykFOI/z
/hRV+SzO2m7ps0k4A08IdV/2ZajqThjbw5tQB2ufJ9d21zAg6zf5QmOvV/TBSDLU
gzWNBVRpk93alAdPe+1nhEOqELaAr37NjefVmdZuXkc8WCj5Q8D4Cn+RiSh6PSWN
FlG0P8zEGDsiLxkrtog4NFMr6q+RIbrYhFimHXlz44jkw3uUBTSWz2dc58UFV9vz
jtuUl86KyjvdDh/X/xM6WD7WrDvje/L0ydne0zD4x1MTPFv5nN2F6m4NsoN2dcPT
NDlN1es8AlsksGjhVZfZNAlzoyks8mb0FfMnSb1+XxaCdTSOvdWOgSW9MZKT5QD3
XKtTg2Dy33eYSiHWIKYMGsruIx/ROUFUr11tQ6oHfOfoGYHXB3oO+GyxqFzXO/PB
Bdr6N+/Xg1iBI1AxBvU0LSCMxV6mlQUCkQqiUZq4JpNhpcJ3zSiZ8xsKnhylK591
vOu9iJY0W19LMP0TuzmWNeeBD/Spz+xTh+tHp9L0WqXq8WDS8IA3tRK7VobAgx74
yHTJFv9vv5gy47JT/4pqLs/Tx2QveXtgtk2ZvWri45s=
`protect END_PROTECTED
