`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbyPeb/P50aQDF5JJb/LpGcV4mmEogxfYHE9ZsitbUiWq+syH98/xNVdmLbaT0Ul
mLNwPUggC84hdSCbcqikDOaP2T0D6VGMHwvOGoyBZtf44ab65oNmk32KS0t5OI7Y
rPcg2komh9kH8IVUxgxGYbefILJHoaxUj+UTD5OszpwDgJSNBnJxu5skTmiSOn4n
aFc0901O/X5xb9+pBToCpt4YhC5YVLJK/u2/oIoPaoP/LHXVueYs4VSPv9Wvf5DV
ESo8Na9Qz6VFqXBrvYJsUsEoKhZwR+32TIGYRHtEL1O/X8Gy1pj9VbdCUpQOt2iB
g2gqPB0cX8U9EumwpX/6qzkS6k8baOiQWEE/YsA6cYakudJejiRmCl6X9j8Z+ywD
7TGKsnptruwRbsSOm3lqQiNypZ700+I66EgWBfbc6A9M6U6iZkANc/GjhwhRNUAJ
uuCXIaAotOs2KmabH/RmX/rO8uMToebS/TgATXUverH6wLfYOb4BZjf7qTo6WORR
LRGavXs6B6NShg3meOfD6QK6L6oZaeawb9Hwkbcj3962E2Z0FnKCKrheT06lsL5s
D6qObrGHr/spa/wjXz7x9K/5aq8OX4bPSiUdbQ6MB+Q=
`protect END_PROTECTED
