`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZuLd9CCe+CdL1U10CuJbhCteZhIALFsBDqelyrNjrl9bvy70Cy2vJZwSdbvbKCb
zflDoDwoKfsosnarqTdqntiLXx4Xx9INrAuPiHP/sP+SKp5ds4nD14ob1PGj+imt
ET1FbJQpigRGtLPvv3LGvoVH5lZ12X5WZHhIW1M3HOg/dWA8dTtJQs9T94dW9Vt9
qbIqIDWQRW7SjdZf2ujvVemOyLFzEsmlCC8vAnLXSHyXJIfUpMhpge7PpQDAz+9O
MPgg+5Kba5+I1iYwMRG3YU6fCxNZC/SuESeGzQof2eHoENJdMOE6tm38Q+oK91lG
E2Ni5O11LeZB6wlgGHtrBA5qUDHve4jky1u+5GZATMU+r5U0CA75Hf20xchRNAg4
eJf1RDNPueGiFh5yWCy03+CMsZm7KW+qfbS25ubE7INt2JO03UXF5mdHHKv8aJml
gve2kfDlDwNHRilrKbiyHsStBSriPNBYamQI55W8OsOBZwpXz49/lHZep3yMZy56
jJadzLomDU/WF3/+tfCpxnkMnHiC6m9ICyILBIFLZrcwCTaMRo+AWnAWpr908Tl/
JcnXeVWcJ6ZKQguanh/vjFBQnhZYEMHi4HfaUy19gbm/6cqre8dURrBW/JwQ1eME
C8OkSamAJegarrW5OoJsgkK3szrO8vgR/LSpN7MrTvXilJcVvSB4TxdKiwuFGx16
haz9qViiobinsK1fV8ht2+dFb6JMeebyrS70daJwSKYIY37GGpqU7ZgWd+8V2LCn
sjaWFy1VQ2sJlDYC+/jtdI01YQ8x+o4FmIorqCe2t/f1xBnq33NX/G4ozbYTT5SW
`protect END_PROTECTED
