`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BYXf1g5m/XRRDOn5AAS8E5Pa0qYKMJGJxMFZxxlC3HgKOLJqogBHyq3PJNVBat9
w+Pmh0WYRV5RUsoVQ0L3WlSOdGfL56zMRq04jKDlpnqglOSFNG5GRatEBzkd6rE2
H2VfXWy8J2SfilkgfWAB29YpymT+bx8JXl0PiMKfV20LjJcErClK+qe5GpKuL3mP
0M3KT8uch34YdPgcHNfiojmqpac7atXdG0ZtTmLhKcfTZUmR07qbZinRfQDuCGpi
3C4vXkJqYwo5NJ/hzDmeFswI3DTx7N1pqo9ub97HM0P8WfFfmulJDi6+L1ihhbw1
/6Y6UyYtPrhEy7JQ17o1kDjlUObkRTAY9OnGfB+5LIKzJZkC0UUQ31H18SMKbm2m
8M1Kq/wWSE8IDA+CWPcpVmJ/znR7ulb5t3sPa43C4jqHOmXLdQA84x7R7xjv9t53
yGRIMP8yM/sAJtWQ8rcksP+VxTg+d3VJpz1Q00Q//iaSZkRmKhv8Doc/K/NoJYcS
uckmKELdecopvSSDrvVeNb8lQ6FoE9MErxU5bzJTHq5XxqJD9aAn1XIP1k4U+QOK
SqXcGmQcFc1ChPj2ucKxpZQVJkNKjKOtHJ1oVzCOWm3oYLuUnnumdn3WMpekYysb
rFuGMpDx6SWT7Llwk/4vrNrMfBXW3+SC5Gz3/U0oxLX4PUgbLUO08evVpItj4aVC
PUypA0IeRhFLGO/htjfGR5BSqx9EhYV+8ix2zMcAu1qQnCdMpclfDMolakO/SdFY
0uXvYGyQuOTOM6TwqDU5JCn0mq1C5704VLwc+vDIP6faSxL6c4btD24Hsyh5lGnb
IT6IcDf+eSDYbsV9lh92NrdTf9FKYFh/mh9sRicO5cKLOc49JPwCSQo+K1YEZFv5
kfPBXMGgwX+/huDljtD+0neWROKwpbafxVZX/WVYwyVNWT9asP/fbuTdkuJdAeG1
a2vSocTv9hfVNZ4PTjSPU/Y4NLhoSbwSurVH7Grv3n1I/sBRDxtGt87B/exejpMp
mG6DDrC1sWRmAUNSAma7om0nhKqyYNK+XpIrDEL8usw=
`protect END_PROTECTED
