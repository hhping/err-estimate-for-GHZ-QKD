`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2I0ztu4uJdsjnfBgMoM2q1mdi23o4oy5h1M/cqKW4YmPiWwng9bxvPvd1FEjp9/
26QW7KGj+/u/O+5U/tW9yaZN1rnmIlomwpWe/CarDUAMBA73L542BM2b8GkdTAXv
fbSqtqckI/6WQ13uDCSsPocQROWCacg1TQPDTQUBYmWKXzExxgZhgkupjgN2cHRb
5ch4Vj8gCUM2nJQcN9UrTw8LefqJrmVdF2a1Su5TZjLimV264n5+/ozYQODQVf1W
fOblst7nHQXB4+Tvg49ibiXpvKfhbfbg0xtrErv0hXc96OFyBGbyP9m3OEwtEWH0
Xse+zBuO5o3+HtuTPvRduXl3RN3nYuK/fukHYyd70hALGQDYDm8yox0c9mb83E6s
RAVAUsGmQ/dQtS1NTbXtNlGsdJdwxXk5wbABOo/mVDsZWDTF5g7XBx9n/qkYaadr
iwKPsDJDrPHLpcAUv4sGkWehdv25ebbEf+Pb404aXkM0iD81qmEOu1aBqLKUtBlk
typ1Ti+DQXiaa/r6tIXJ4O2Zy5dMZ/tRa/C5zBLGVoOF9yOK3cblkFt/4C3pUM4I
kr+Z+6SXZ5aHIkGiVzuuiybBodIFJKR+CXqN63MOUDV674SxlGkGQxMW9C/ypWTj
kyK3rZZ29WE4gCslS+T5dvw0HpKpA2Hmpw2ZxgUaN8Hj0rsVzWOrYCG1ITtH2FtB
+pIuuhG6PfH/1w06MEIJpGpMy+97Z30zN67rDncwBvZRhYoEuAPN3JVKtJE2wt/m
3zWgO/EPqjvxjMgq1eeNpLaVXgme2N7VlXd4nW9YMQuM2wTlZ/k42dZPIY84u4vu
NPUoqZux8P57oIvtRIgeb1DDMYqRucjBUw2KzUw59G2iLH/RLRG2As4dPZzrg28r
bKjzBGxXW77umQv9GB8gYGl3kjpTIcieVeGe7f1emgt78emYjhDtYMDkCdwmp0po
I/rqh1OLnEMjCdeOh+uFAzr2HHn42cPzOZ0fI1ETY7ZWnFCwN3nhr2iXOYS7A78F
jCIbp4yJekz7xj9qmNVqG/aIhbYWM8WaL9ZswiFct9/d435PrZZ6BsfOO6hDi0GP
BecWgqOZI/TBrT9cMgunMaIUowN9ENtGQqJfil5uhmTwTlM8pP9RSqzk3jCODJFt
etXCCyqlRUuV80hvDJwEvil1avgklaH1WoQgHhfu8zU6Px5UTob96lpzmFHtGCDT
QEtBFslyoQPfgMNOcIhVSZgYm5wZe2GC/yyTe3AbNlls5PGtAT4sCjzc8i5bY7ia
YA4sN9650jQ1OTMc0s4FPUy3iijFkn2tRrVcu8pxNaTTzinBrTaHe/UAMAGceouW
2IcH6BYfp/aM7un9t7ZoOFRwL+4y1OLRgNXmdCM42g1+I9ico4DaGqYYuJSjWhpi
2f6+QejrllxcxbLrUC7YsC/kBNqoYYZx86YLkxAI2gYV6aDDEziXtNdVaWVP+W8M
ngPRQ8M0j2UTRfbZWSvUsLwPFZZEMWcjNOq1WS9dotDiuDFaBzPyZ0p+NSnUNoCx
y17IlLLM47pmAXP2BVq2+XxSWMS9gLkO80WafgkVGAB16bmWBEltoJruMDtnu4G6
A/5Tzrc6ARtXZLcGqWEm8NqOe/kQrr9QxYWWBnyg82cs9G27gAUD4Wh9I68oPnSz
oqTBNimfdk906yBnENyawU4kWan76shWyHUnNdDdORbaDA7oYSKeelhCp8OElMMK
E86vjWVcfdVeSz4SmSEqsjjLCmQhyM80fn0fLlbuwMnp8a/NnqoLXCIGV2d1Iz1t
2lqPu/ZSkt8G+P4zz9zF8Df7YarmhSZtcF6I7lzrgZf4pijhj6rpA7u4CUfVoW/k
wjRhbUBUN5uE04uarw4CJQ9DXdaKlw6uKCEPQ1qTnJFQUXX6WlJFSkMFO4HMaRbA
FxUB2/LKpVYoH46RHp0l0C3Fv8wHpdNcnlJtJ5TFTzwPsrBdEZL5MLD7MhkGRgOk
OE8IHQFVRYeQ7flKEMtNtpxXwHaDE9Cy7qW/nC/KS3fwMmtf+FqEdE6qB2JT4QHY
fzUrX3nFHhTMgTyIC2yLoiHUiEBbVQVJ5eqXPxvRzpZL08W2vPCggRn0lJoU3umg
H+JiV9BeBy0N0weiILXe3mBtGImEltzVQ/9B6vHTC7IhuCd7APHlpUQKAjtYTho3
r3hrEN3KPRx7sCWbMthKfeKMrKyXwJmJAzTnIYGb61ScffdTfFFRf1ZwUW0H61Ow
RimbtIZp8YrTtdJBzfbw4ymG3oz3oi17X4Us0PNSdBPbPuR58CzVnt+f7AeeIAOZ
yqI1781XlzkR0y7H64EuKmuFcYg09uELPshI/5oiKMvQmrn8wvuLnk9cqb7eYwse
VkLOtdRV1bjErUVdRkPfTCTJgVILifJMRVGR/a4N3CWZjBxB/yuV7tktA/zDVQaL
As5AjZSABRUs0FOsOvua12uVQ2hMJ+LaCZ8JSSym+8VSZ3CDuv7UaEnZIjxRhup8
ht2XrPBEaWeCiKm2576d5olTxfE7ror5oOLEpeyD6rTvtxdYK3U8GkQBymx+9Zs0
Qoz+RKg2N9/akiaL1gn/qUCKfOL0Oj0elZhxNrpP7TRIl0u8hZxSGTBTHIjL1Mdi
STuxwMzgTm+tsX7jIqWYn0KBDcTDhsOK/zMauP3TbhrJ9DuVY4hlzq6b1ORdGXNF
UOwkETkyaSdjXMSY8xJfUqtvcrxghSXenryi8SXkKmq8Vi9ly5yRc8rPUdDuDoe0
sxTHnvJu+1UZ9/4K4DFalaGPLhjQy1rLEzBqh1RTHCA0slO3j+JmeSTEg3oFhdPH
7ALQhZN0qZA/5BSwohS+op6HlSxm/H14M5eCc/EqBU05J6ReB+U5p9m25izYM6v4
4zHBchziA01NjSGOcWc4Hk+C2h5j1S0XkD7fpXbyymDgde6AEATELW8F/8MG9SVk
WyaDdkZIpHzTpAiDVVpwy1ycbZVtpUticZNkUF4p7+jIG07PwGIADzzF3Rx+dTGk
tfa54hHrqGQL3Qt1P6OwSs+/Qlu1AkDVzLkZQA0/UZ1hr1MDzGcc0gRAJKTdszCk
KPzp0lr1qyiHP6/3paRhKg9xcPndSx7vYnAxouRoimrOS2hbWXSh5XIQ9a69dG4r
7o2ir0+GJ3m+pIWwAUSyXmv4xhXtAe34NbaaDcoW8Ug+5P3/iFNqBFAuFb0hwGB8
RK9bup1YdDMtMoEK/9cH/fD7TmuSnRe8wJ2eC6TudM8S3bO+oYRg3hD2oo855GTH
jISYm0gynumbc4Uh2PaelXGzzE1Cjt9I3QAyHe4FRPIEWB3YzW3tID4vORaF/xR6
fjGHbCASPt/nw0YwXY8m9y7Ey0qoIO21uOErvH0BhB4JsJImoY7UpyvtuDUToCNT
0Ui0TKvf3EtBBB6wkoZSSYLqsRRiG5xfMX5W9c2shQdNaBlDmp3Qw0boWpxlaQil
kpC/Go2oCGWttO58JBF7xqYQcUgmuzEOn2E7fCyDWDU1DzHn0DQ9c32owP8QxCxy
H4AdVqlMXu1A9OrpqzI/rztgTs0Ur7TlASVgGgOv4hsXJ11obEvjVjVfx/xXR/sr
mszBlpgSYbUUHHsLaMQW0UZWpZyzF05GMl+kGHTj027fA+2wCrEMmZ7/ZvOSCZb5
+RACMWAJs8Ow5NlNnmoAFriGfjBLRGtIMewPVvTS6KOfqOn2Wy9CIoeHD4OZ5exk
jq9zGO2IzK74UIXpZ3qhlTtRRNRPR14AqD3WcXS/MjEhQhj7BZk2O+TSmFF6SRvY
fv+FmtpDM4Zy5m8bkP372V228J1X1+PIpsSqP/but0aQxJDDNlJc9/2Jwt0I8iUJ
HrGDIFHXBJmLgaPy1rXR297mEhNwCgoCPY54zBlq7SelmM322kF6AOhP+oIUsQUF
Np0s5rlvskbDIcfK/6JQuyEYCCZBbmn0DUewHejvDgaUlBw3BEu/Tv04J1fw4Iee
RgrkYfOG4+gPI3faECEg+I2JHWSp9f6NdzfxlBtEVnPu/AU239Sgx6YFPMiRMtTD
cp71Il3uXCGJodXv9uW48UnpahLMoVauyn3cJImWudPoRdlw6bJ7TLqAQNdvdzSE
tihSI+VX39L7qWqJX62soVhAj3dhe8dm2OYKpNHaVd6OsM2r2Vll9t+1V/9Nysbf
tCsM9wyXU5WJq6xFa7WZvIRp4iIbjErOgVCDqQ926PRKwUlyTS0mhS5VoIRtapXZ
cidyJ6FY4+ckwBqpTIfffQfEoPD6H+d3wfQC4vJI6pFcV05vz9p7IjVstIPDnh+K
0C1+yScoRU9Ue22p81GPXVQYuO2045QZwdw3d74ZseOTajH1GOMPJdlj53+ZrowT
2bUS1NxkYmOjlo9VRfjKgW7/RarU247HysI+6Meo5NN0YSgcXKaSvLOwx7BGdPAd
ZAa3aolVhTH46Hdl9RXeXqAcSBKLZ4DCYhUl35olUJjQBrvA/GEcojFJ6Q2QjrgV
EI0+FhvxbdDK/fHz+A/g6GKxiiiKEOorndK1sBX1UOfBw1RlRDWEAbPu9P2Qq0+6
xokhBAVFwKBWoSImH4DTZT+fVw3VnhR3AU3at4HynGtY7LVy90Kv+aprqA/Ihzam
z0bnRqK624x9z5CoPxfx/aPREvXc+aSb7kvdAPKBYciHA3xn5W/o4Hkkxr/vjnuz
fJqYXGp52HXJ7uRrt3MlEHrs+pqyFOXNWpgjY30jQJG/HxulKUF/jWjttOOb3Oj6
84obJwOwgp18CFi5Htx5M4I2JkcQ7rP6LX3/jnwe9PjzG87khw8UWG+xcKqRU5fi
o5ZP8doFaNKU+ENiTY3bYwN4bcj5qWaLKwzMa41x2QTNHw2Ut2IHIfc2NSgwsCb5
KGl/TD7yFWteGK6OTRKbnkHThbrM816YwMfvs7MTpw/WUF7SQEIdChXLPkRSoBy6
qRDgjIePX+/vXGjE5vpyV5ldbEEVWUzFiWfMb4B8qs3sD+Uz/3F6LCP6t8c0vGsD
Yw7V9n6PTR65ScDiG+8wfdcrmcJwR0biJG84XmuFfV75jnQ73+PbIAAL3fCx+H5M
Xfc+3tmx3av/3vAOqiY2JCO7kX3OGZGnIb1qbAvyWjDupR5m/WGaDz08j8vBSQas
LvsybEBaZ9sXkNEYPxds9J7kEWFt6sWGkvlOrlchG/sOJhC7kvFnzgWOHik/sjFp
MUoUAgZhww3rukmNrSsKTYzcLUQQ6RSYn38L1NNAigEUunzWSVgS/Wk4KAuSsfyY
tuBih/3DVmCwXT4a+udVlpljVs7XuEQHgwoeVxcPl5Mrdc2zZJE9tCtaYl9xSXUA
iLeMfpcTQlfr1jO1lz0Aydxt2oNZEksd9i6O+WXmfukyrMF/sglSVbdgNg3cl26V
6waLx/W6/dJ2UUyNRhCJUfuh3zHb7PoMcQCP7ZC+oQuN5hkfuExmfJgi3kT3QSfm
XyPGiEY+zSsHup7SCwVMFO0vcbPPvmURJ7ws9Yk/TOioyDI/PQ+h/HXfD0ow8d4V
naG7Dc5oVqutA7pG8FNfxFmp7yB3qnmK28N+10sG7pJCoKCbT8j0v76pkL/admRS
jqhKJDnWu4N5IXS2+qaJHZgbha0+xjmhAvKx2o8OjySzY7A6IGe4ldig2p2Bbtnh
WR1AYPtSZGfVCdPBHYmkbT3xQ/wzFfOMCpBnCIiQDM53ZnoTlcn/BK9/4+gMnluG
3An3lIOaCd5K3HRbDDpCj0pj8lqYHrd4eK9OwgkGtFPwGtX3D9cR5tqJ3vLc+UAu
bovSaf5r4L66Rt08//dl6HFX4OlYAJF5zOUO8H7WWByTSQvKLtuZxZZRWZf/pK9m
drdXBKNfHocgjxDNjWfggyjlfVx0SRasmUcAQA6o6Oa9CAZ0SQgI89D++RzTyQmi
DJjMK+5QNYs+sx6Dy/SQ1QydGPPcDJm2JCvlDm29eVJOUVAOZnQ39Zk/SqSlbtR3
7KTmA2YFwY8xLmHGf0IxrFfPyCZhcP0Kof/p1cuesu5q9iSXLUfp70/usqPz1WtN
/ixf8pSfsuzgdjpAImuF3WXJRflMkqW8TQIE8VAmx26oGeLrujmBQMgJcAoucmaI
30drX9Pl67DPOqC+s2ZvzsGeVsPJzeeqGrS0OULHMTsjvBmx8ji6T8ocTdBXuoB5
sHLpvVrEgyG1SYH59TWGnNZtwx+qrOfIUzYBbM95WpklUxsaWpDD382NnSu0/hzT
b1eRCp+vnBOC+LW47FD5PGNgnLwS95TOUMzm6SDzjvByx0stL+0+ZoeA2febU+zH
erlUJgQHunEHl1vjha6u1k8sAQLfsQtgqozjr4AVwvzrM0q016hUR1drU8gYGsM4
nRw7JLc/dfgBdTbZ29yHWBhG90hbEtTetHKdZ7o7mPynh6Uf8SCx75YDGnnehYjM
wT07DD7fTu6ZUQNsLCikVdlsoQ8fdgzjhQcfntt5d4eIyZNDFvoDEUemkIX3RXFU
nOQaAST+ArMMeagR1o7SyFBaXB7+tCgDI5sVvzGEMeCqxPe+v0WWLUZ1q6gLr3eY
Bx1l+H4MlFdpHLL60gUxl5Rxf6QgSW24vfwxFYAB6M2AZrq0c6sybewhu+mcyUP4
mJx8Y4C0drEJjncLmlwAFib8s8DCOnzLdm/hY4GOwtm5yjgTZx1I7TB7gYs5iguV
/tnpSbIWGmcpBxW79mWO3jzBivub4hyNCDrn21Gsym200nWppFIeILG9TpypfvXf
uI601JLiP2ZDvPZRaYIdasUEIfFY8LjICRxw53jmW61Bu2l1lJzVFbISh11SZeFF
0/hjuNuF/8V914zm7XdTN/F3wqS+qdElBX8R8PZVxCQBDtm7EA0kHv//b90+M/Zv
Rl8US/iqDwxX7cb6dYw3HMrfDd/m6HzOnEHwyCedTwCi4CU9nNfiBZ1K8zRUfoaK
hZZx7tdDrUOPKaKhB5dmezK+PRS2wNjCRUSvFyJNnB/EZFLZPjK9F0K0vb5Qotij
X/qGdlla6wO1rZMCfsK1fKBlOeOdZBgvSfnb7KYMQtmIi6Kyl7Nw/X9QvUvHwfPS
7/3HCW94K4hwD0qZ5oY4HbMzUwsqCoT4OhjdOnAXAFRClHE/6rNEcNSA59WQTkYX
mevPzZA7mMhzB1K9kW0A5AtON98tmOVOZjSb2Ev+g5VPuqeM+VwrhM4gRkdQsP8l
dWUuLtwNOq6esrQGsZQslcZU3cQQqFi7PCN8fq17LHBqe1FMztdeIVEOquGVWMu+
azl9nbN9MqTMhaoG/0BS0KoKHgNJbVHPwOGY5Wpr/8rm2RzZkEGz1SeRXMFVCjT3
iQfzdMiBZUgNoJfVUeUoPDg+ajkYD4qDAXGFJ+F2otRGB4/kr9YJuaKYNSMUvdkt
7rX+9YNM/e7SGC6XlzMnE0lvm4k7GNCpL8FQzSxR8x2TFBksCaMDo9tfkP6qPWhw
K5PbwdTjWk01s0cmTPxrr8YFX365j5UcGN76okCbhkK9NaeUl2dYO6OpEZjBCvUu
8Pi7FjkXXP+H2PdRfZ3c1m0GoArpBC7hAPVLUCM8AaLEi1nmwZLuNG98Ow/upp/j
+ipxLtzRgM/xnZp09b6RQD6YcKqEU7iIoqWIKOwQ3mcfIz227sMM3DBk91STJQ81
1Kvkl8e9UkoIRp0lf0RFDrwYduE16sVk+pmtPg2BBuk8mAZi60luk8xe+UoXI21t
OHqZvNR4I7JfDkpmGN0Ce9mMV7e8GmET9FIWeV5IaxpmEcB3l1aUTnMtrgAbXIEv
hnHin2MuDsO8ovPcRqN0ItOrfMkzPmdHPVb9pFiHFunIcvkSkt8s3LUhvrOSiC1J
HlDs2peHY10V15uq/4Nu4l73+ABfmYGvtMSwIqByh41Bnde4Gqv2zIxpGwE3tSX3
qTRpKHFBqmEjmfDuyhk+OtKYN19VTjK0KmPHPc5EVEFWc6D0DbVope2OyFzxKI+V
v6gQjvn9GhARSfr/P8CxJ27eQCDqtqlTBB6u2I+8CK1o7Aii6wXVErl7r5N/yS6O
oBZ9SdhdrYEHBHO1NwGVoL+E4K9CpR0h0x1i7km0i4Pf85g+fEdf6bx+Linx41k6
er/RK2FjQ3Zwr4dNd1Crqd8YP5wFwJx8aoxlX4JQA0WeV+U4u9zsnzlbPR/IFOpW
ksyBnLmRj9SsDAK3afThPpwbKDwE0EXu/tYvzjU/JZBw9AcxmM8M07HbgpFo/LxY
t9cDrlbgROyrmaz33rC1wF0EgxDhpWuNVZguZI5y8tOcsxKmEAX8TMcDbyi1mXRZ
pD+MjDZTLc9jSJX8V0DD/+o8ev+NckQSUxm6PvGHnxS0GNfz4RO2q03m7dQm4msf
PEG/Io5XKEJLG5sk7oSxqFLj1sL11J/QKs37dyJ9vG3JVMOH6KDyE7laTGEkqm2T
ziPYsgqOtT75MDu7kEn381QrAkk2OZlBYwcMwW5jmHYosL6EvqRPwJdOFv4xslG2
vTs8qNk83QbYsUitYUBYUjlIWNvjK8+Ebbqi6RYtB6XkbqgsXEOB2KCMzKdcwuZv
dabJbGtaLxIOVkBSnUupzCluJFyKsxHYMfsx6WJ10uqFN9Qn2RwHk1VSkchZ2I17
V6YpBXK6vR03iRFoOnl/+lMkEprrYdMseHhOFmyHpTAebvTWae+yegHTMHTrc9xj
UCPcxCJMHyA/sWcamEKUQ/hxhWjBw13yfVFEyyW4666E2X2w+xE5wTr48fDCRfgs
8tZhvbZK6RVAyM3/dGPl8EeqbwtbUb11hww4tLCN52SHuWrTlTmMePClbTUWH2t9
KLhcbrWkFMF9+lKu1p9oM7R4i/azEg3UBRaQKtGTY1bxGGtTYa2J5ush0QzM/tzS
Chi+wCg/HQ92R/awhUJz4l564jb7Mqb7GuWIVJ5XJWWvv7uonNAmgqUkapVloWcn
rFN/U2r1FcGAJEw5UvpHV0LCfy7ZPww0zflz3omVMivcIzG67RH6v1C1a341ejZE
aPY9h0kshW/pD3BIHZjQjcajjKjE75DdoHhAw6+lXpUbkl6dLqM4zRnhLNMV1SWI
G8xFynjQY2fk6uD7eu23lkdT6gIsxjjKgJNBit9qCPI6OPcKso9BYNCz4ThXAqdb
sVpBBNqTw7eF47OPNak+Znd6lxx6tcP+HQhc9iNCN4ENAcMdElSsbJ1UzVJ5/oIc
/09G/dhYEyuL0auFrHnGasw8cYPzHFL06ebpQk1ZVH9EOW31kjK8BY0D0FApnqRf
XMz7BoJyYzyjgPXuYi1KV6lzPIX0an2n3MKcaxAeBY53cmhebDpqnNjhnBhHmrJf
ICH7AWEEKERVv//SNtWded0F0UOEVN9min4hNKycwGZvPzKTbGdbU4bY1nRBPhiZ
GoDxfoREfmcJr0YJ8VKf8RFNq97crHEiWc+pyZ8Oo6I/klhW4Rm4FDpDhHrJaD8/
WcRrKRPMgP3tQi8nvs/88lVPGHACNyqfMDTfTlSrVntEkvsB6dG2P7NNs50iIWXz
TdN8x2DGISv9Ob+t1V1xrrdHIWvgI7XJkzfKdcuA1whroy22BevOZIAM9V9Ni7Ep
ddhYDwEQP44QXgyppj5tc25MUi9W/+anslCKY3i1kdLiTB//WcBJZ4bS99Y/IuSb
5CVImfs9MZ2t9HBg+t/2Xym5UybHBVfggzbsbxBbFyMHIikip4wutC6VtdEV8/rH
boLDwJ9Ktky7f2ntbUphAdv36jo/eXtYWVYBdvtaA0tkOdo0ST4ZaHXbtP2LCZ8O
EPJHkPxmlw8rWVleUL1gNFop4h3jqNc1aisU0uc8NUkDPQKERTHj/v5W/RynK6ev
r3Ygg7D5AY75/DxIIzNVberPvh14tMRkhcuoMJwwe4NRUNczobUlCmwrHSPBDckR
dezlon1BmNF8cQuehaHRy/LH4JkWfy80gB3qZ2LVKFbhF0kY1iKbQvr0gk7sKt2b
05Icwvw3jWiyCQqKoC+BfYTRN/Ws91GCilE72KKrOHB8+eyMh4PbtL3u3fx0Qfm6
b0p7/a/zWUekUSlY7C7CZrAuIwaSvJve5GvevmPLmEoih/yWMKTpq0IVdFWqFHqZ
YFlcsEdoKJlPEk2qeigV/NCT/HDqaX4tgVP7ZpOWVWjtSvRl7lX/+mjYSIa1PlYk
tR5E7d7fo3kdl2cxdtiC15yghAvD0mtjxWX87Y9lmTZD2wr4oefcFfpKiPh76aqi
AsJz2si1PsE4K6VaARhYmaQ4g3YGfUzCcJhqbjeXI1LIgaDfO+J3B5/Zxe2w/0l7
JYY4RfY17RIDUurllhpEK+WwxGOijLcDB+3OIduNioEXtW47Fm8R9VXipIs+Wh5/
N76kl2ywLm83HaXZ66gL21fEeIcKwW1OCgQzdcmUWazqgr/kY2/lceD6dtypeG3G
UIWTYH8u81cXge8wT/HRGu9HLAdUTs5onQDMIkdNfHIRPh4e7iiCliNlwOsvvZzC
pE3BmurJJ0URkUuf/YcuO384EgguMxUAoTikLwV1T6lSrq4lb+7UWPOA8rohi1gD
dWeTN6VvQAQFOSv4j49rGkEe2X/c/p/ixYUk3DaVB6pAmgZ3ZiHg6hQdxOlyYUWP
REVivazk5TzeCV5qY8is7VzqmRZLYukOH65v6cEQspoDqCmqTOMX4+qMevC/CHx8
4zxIcnSJtSu8PycMHOLmjygx2Ib4DAlo/KulLxteBMG556aI8MpEqs8Gecz5uY1z
KqoCu9JDKX7XwbQ4We6p01gFeTL2GkpBOBEB/hE0bwAl7eTnhSQsloZBLi0HYDON
rl56DDtWHySeRVAedCIuiwVmlQ0Z3J0/G2PNM2WPKEDAlzt+Bt0zqOTTDJv5xeq+
OwOIleQl21uHhOs0kqPKrtJUbti1A++yT/eU1/dVN/dMUUQn+dZcoCXwr6nsmN1C
lLLUKbYjCPYuVc+Y5VvD/7GmaRsqDHeViY2gzJl27wAN/GO4aiqVvrbP0ByFwv6z
u3k9tQTiLGthnNkt+ww5Wq2R8Zuk7j26ErnqL9jng6OqqbIZnBIq73MIFYeoJrmD
8e//Z7HkEIAYf7cWaTsU2EwK7fNcREMTYQXQO29jO9yiiW6/sYVHOLlxDdhMFADJ
l1XoU6pcX3jj6OOtnJRySUErqyXKqpvscEoW9WYW+9QBwYPIMNqMkx4xTxaxrHy0
ERuJC3OOz05/haucffle+U6gzQAp7nqQF6rR6btshbUbZfObawhcEZg7fxEaxVCU
ax4LbO+ivgAOq8w+KiAIEwKcUIXDVsn9vRsz8OTsF/9EN9ra6N6l96GC8qRt/0F5
1gGAXP4ydfdOWxRRXXPiguTVm1972RaulMrKYDzvcNi37wpaCcpQW8zdusnIH4Ru
B+4qoa3ed69ROJRzN6ocZ70epCBuxbE0yWm7+HNfARMB2EfgICoi/7d4PLjfD7K0
4rx7aUb5RncVnH8TiJ21RCwRxAIX5/5vYbhn2Y+9D3P6GsW687YHmfojwZVYLl7Z
WwshRJoQ5krpHa0kz8BQKH6n5U6PgdzmTUMDCr2G6IESGbOEvSuYW9iUdBIKN+Gh
4Vibmoa4UPw8zXvSoshAaM4y0GwfW6TKXaTaLI2+JEpE5E2ubB+7tK2qG6RMGrZ8
OU9UuQn/2XQ5x1P0plkfrvYfJngSnnM6QAIscc2ybsmKn4i3xnw5FPMn2NQnkhDd
VMpL7mogj7Q3JMNqEjz4qPR44/Lu3KPvuVfWdew/g5fMqUcLN2qUYKm67wFOJVZK
5IMjocd0X1yg6GMn6TsbowKF/utNfgY1stM7R3Z70uhY/GCNCD7qyRvcPuVIVhUJ
2CMmHnOtItojrooTkUIEXc4CSDa/rQ3xY+9d62zPgLt+NHpCh29oNX3YZrPGShCh
+DKjxXzft5O16C8iaAV7sam8Lc9s/McikAGAWqmtBlFnBmMOvIBbIJAvM0AUZA0N
vH7FUOg9jFSHyJ0pojtCTDGJkVP5Xr4M9nFohWWLlWfrBnCxLkTraXPXsoL/xd+k
Vn2fgGsHDwrX+q/ZPXIMnrm39D3sNGmZEEhh4H2rioZRRU02F7x6VO6Ggm/vxtfE
nyxH5VbLF5kVHsKwc97AuP4/g56t2YZLWFW4oLR5vwppA6tq/ciW+krtT8rnC/gR
TBROLf2yJ9SlmmRMzLjbRjI8ZvVUWMvhASlCdVWeQoSxJx6h1Gf3xv2LE5wqjees
uPr8zSVKbRuIgyMJz+N7P8ZQI+XAPUeOdzYE9llR2FDvgy0vqb8Fx4p//pT0Br8Y
KtVYoF5cFFpI6ksSBurQfMMI790IMxqr9rGkJLqVygyDVobRkYpURiUCeN6LkC7d
d0ihRW6XV5v7JnJpR6qJABagdj4zS8jxUlTS8IWRd6hKnmHQyGlvobgKD8mDTRvc
4ZrDKrtq3o20sTXxxQ0vDhFbygGKw8k8WXMjifIuF+iiQSi58MJ3iLpg0VjMe8Wu
+13u4uWsS9PRwr0AOw9KUWlUnpWwwYlh8luIxwl6jrnNlv5xZFHsAHlAI6cS6mNK
i7ZFQCaty9K8mSNOVFKRNNFzGpBIJIR6mFfMBq5a6CrK3fG1oMx6WSkA+lgYJuQ+
Fc0T60l6lOSJJ/XCUL0NKbdEaxkyzKTAp4di8fwx/qxCdRw/VxQfMOk8DOwdU1i7
FMmQVimzCSyIVTB6Nq1M/mubCLhi3ZV77I3ibY9LdyNIGQ3fp7XWDo58AkAPCvAv
RYUsQX9Kp+iLn5sgn81XaZgLWKz7IcByenh/6e/WCMiDdmcTJWvEKBZLMDPNnqJf
wpLFpE0X5PvbquqFJxr8sw13l1MpkG6pMQSpVYsMUior9GrUCxwH9lR/Fka7+FkW
lbThqGodajE7S+WFTX1jvXN1rKxAImlQJNbF39LpOPIlm909dv/ZFxeJQ7aNfaBd
j5htdDAOtW290PnC39kScTmgc6IAexiYIKla049qgQJqEa6wCSvLvylvpo03B0xs
mXAhv2L3OboexXgMIMYxDMR8CUNEd/IiXCxf8tV2SS+KQ7hM2FugvVR7oY1CPlPc
2Kq5A+EMDmaHNrmk4VFX5wlh/YRIu2N8h73CfQuu7tLBf2xmj+S1aOICWZMGzEQd
1exa6nhrMPmt2l4x9hnntsfR2m85YfBcV2gEDdIwM+O88pJt/QptOvB/ZyPxWFzn
+CADVfNBXd9i/nJ+N2x6YDhqXOJoecmi01cz4v3EHv35/Eq95GCvtv1OWr0ADFPY
m/kG1zfPoZsCcM/FVyReB1hU15zZ4ReQXX3FtqGwk5JzT8N75N+ALF9ZO4qM1LLN
UaZ77x/hDnmOGKwuOInNBvJvafM5B7GU7ZjB2UFHJl85pdk03E/iXQ4PPfzm2HbF
N4otgUdpRFeig3m/eV1uaCx+9nfzZJ95ukY1xrxV4FO5e/xcyNN05v7ooQWVP4Ou
kJzW3pci9JFBF3ijcBjiwX3a8i0bBo7bOFzIibmwooCh0FwZydg5U/RVlLOX6Pip
VFAuEV4FDTxQYa906D748J1eZfi0tD10pfrKh/38KLNJCt2t8sKGvWzTUbAsqzyt
KyEFKNwSDPLzsNwxsAAt78P3pSb2nj/Eg9HAVudQBE3o6PGJ6U2M2FpWinE9NGH/
7EXZCWEMWpR3CE0W3wgx/jeMW7amuvzcNfb6G8OZTiM1mht+75/eshjCGD0irszc
ciLyGV2gnN7eSp4HO4SB5KcpubRyyM34oIDbirPENulZ5/Plln92HuC8pxmIVHyy
podYWu6RhaQdYdY/cEAOykzDCyjp4T1KtpnJ6OVuIq/bkh3i4T1jvIXfw4eCeiEn
hZv5frW2czzxunnQp0SI/mbRNbLTGSgaONLqrstucdV8xDqlo4UbirfxutI8VIhV
0iMzYZWPo4sT98NYJPgCguak1wrve4ZEnx8locBQKnkahwlvdCnm+sk4gNnhTUiM
RUtJ29rxISgACBVloWXNFZklgzQLz9ZjWN1odJhkCLqZHCu/0NY89bxmfY4i+SKu
gOAhbRWCn82pblfauQHtYD0ITHsDTbG5LNklZmIc+4YWtXDVoe+FJSink38/+xdB
N2+E7TQdtXfZUz3XUN1kdbhIr/z24MOY0DhjkLP7Wo+jK3n1sYjlu7fcitgpyI2i
bgdn3xjqLZxVA7OyqVmRPvUZ9mFzwxH/ROc2TWUgUfpm8/gDJy6WRMaAZ2bnBzRh
tykV8Fxh6jk/sZ6hjb2WP6HDrDdYSvc6LiibhNYStql4AHImRlXgYnswkdvpo2WM
ThUZjTjq2W9DWZL5+sYL3I8yI0Ns2kNbCww+44h/ysCiit03wttjcf1xZfxlmRJf
F54e50YDZPALr1PzN6lbYKb6c7nOTmhUzcoIAVNYxtjtLr+zkxjY3iZKDEJwBjeQ
EYUO3VpNT3sYHFovBJUcxNdivZbj/Ige2bQ+3Ammg+BSmHmQPkFlm3KwNnwNMhU6
hFzeGpcrMRXNR6hEelwkE3vvEKX1xfRSVufNJRV9y0fYNzw9mAJwCO74QUl4spsn
RiV3DzcBZrTVL28CuRBxIGYM6POG/FmRvNFY2RpV8YxHN4BcL1T/8cdoPmEe6zzB
0oo9G27G7I4yAR9NjFp6LCc11qkMBcgauH5UvmkQVP3ua3powUtAlpo5LqACBTJz
us1Zm9xlCHwzo5wZ8vUWhhS7EWczMLKiR0fSxjvi8Rnal5GVbtXdvoeGefdOa82V
xNrQg7/4a0av24kiHHKSYLCmAsuCwwRYOOqT0hlCzx/Zzdv8OP42cR2Fitsgnnqq
O3sYRShiqrS1jDITf6W9dNTQqeyOvHVEfK5OTYdwzg/xFzfW5uKa8QwcSULqCUQG
lJ7UEQUabhsUSZev598fX2lwDO1jzntl8UUxRTIBiXweI/dqn8xuKTl2r9RgVsyX
VYlohwl8uC6cJ0igeoLJg295JmnJCs95a2DrRmobvSnJ+dJVeO6/uvUU30LiX4B1
owN8gvo1755nWSYCXMofewPNU0KgQsdIYGTqjKOOMkL3gc5nyjBMWN/v2nTvbhHg
6+20L345GOSdQgHxsy7Q9A5trhNvS+bcxcbsWbpx/QQ5KM03uXl5Gxdu6cV8nU+P
JOG1RpRTfdXtOlYqaA50+kU7eBLDLk1vLKJOEuBgiQ70uDS5DU4OYuju0uS9K5Hq
VZAVamdl+0VsXzULy8f1+0dexv9yjo5RwU01klm1VGF73gwtXa6mpxU7ufusOTk2
4u9GQIWd1w3OZgUh6nkR4LgaJLEw38B9+qCD5U7gpy9Q/i3o5eegfJ2OurAgRoc1
+AqlK0WcgEf0hcnuUMczYnfO2YYtLW2CggeVmulG5kIOlo6GxVaswSvKK8xdfPR8
wITQYiYM+2agX80W6tdSkHe/5YQmnCPhJNr49naLYx7L+d9XSnWX2F1V2rMKalok
S2RVLbNVkpdBCKdkVhheBMeyiKgwXQeusFIY0r4lj6SsoPcO8KIguGsEa4B4UX+P
RLE+C1Diz6a/9jRimMarvRilSW9wjYM7P40YPkbW/joDXNIQpJnaQPt1/1hEz9dr
qQNHgb+gkvV+KmN4nlFGsaVvO1NZoHPNG/W4nIwDlvbd0NdMeCD6OK2mKu3gdK2V
dNNkXUmLMRy7sglylN7un9PN5wF79CIF1AkZRYyH/o7hPJ6QUC1NDBi4zCjM7xJ0
DxFrAm7EcWdi/1O1mBVf7E4Hz/aXJrYOvtQhcKBtb3SVinzj/iPOE2B2P3C5pLAW
TCD01ZGcJBEKSUT/8jqdQV8Ubdrhka8aH7mg+f2/5+GdiSMUVUEudtaysatjgIIL
KnO1R+v/1S5sn5RPtk9otw1rr+E72fuJZ4pMNaMM2ETVUNCc2MTL5OEWm+b+fyru
bEFc5spw+YFXOP445jRMtvKmaRa7RI+lflU2SjY8NzGaWm1pNR8A/yjqPfB7fXLh
R7ZmeUq0rhbAEv1lc/vdVmRi4+j9bIupBWPWdWVWKcu6i7sz/jIiOLV5YS3gqNWt
qVLedVY3SEiZ8TyukBZM5vFztBZXSvArekfLzjFkQxryQiZbtEKPOaMge0T94psA
qe71TTZ7CfZzwK7GSVDxXm36jD0oDDrAuJwpD5BYG0+kwu0hjt7vHf3TplT3PFDw
KjyLR0pCiYgbHKL0Qu9VxMZDL6n1l/axasmQKnQEvWkBp1/lJQTtQy12jrNgZ0yV
wxemaB7vgrLqTWNwIGHzG9PJqo3P3jlkW7rNRqMhfPPztf4941HgqdHgVbZLanyx
dK9NCZZnJfi6Tem/r4eyWjpW5YIqvMYrT8cu5HqnFW5EdKEZIluIRW9hhlEhf1Yx
zdknrWoZb4HhaDzBmBx2P/nvKCNGYjvoRdmiRlG8bhIezTxqurL5cfFKK96dyxok
8pVDryvwbrvZxUBWUJhGbj3d86VFnA9P+owuivfOX8eU6wrtq49rBmhtkxGzlbsl
zF1csZhiUJEHPg7XiC81cV3CaNieBNBE4Gyc3KvfzFINMfb1QekqxBJARR0VcAQm
1WRDqb46thaYZwkNNP9i14duzmAOVXmVGP8xXp+H7IHS+2WuruqnYgVrhbizhjBG
m503kb6rUNYvD0cg/S1W1v50GL/oNrPsc4ZTfWNKucjYOcJEnLLx3lP62fg73dbf
3WnMhKvoKcXQsd4LeEGo/KgMhzeZjbqPeIwdizhURibAHIbjx/1ldDJjyoAhKCV3
Ci1IHR3Mj4+YzrMsGc7aSyUMIQeQxvA581+ZO4GCqFSFIx5RjvvGXXcQr44yjR2S
jpdZldlOc9vEB5ZMyielFbiqpFaPm3fylv7RK8QrAbIMSHc43D5fuzCpSxaZ4RTD
z8B4q1eIxSXDISjb0kROlINFhaxZCYcqglGiXxYh7YYEqi8Y+MOiv04qmv0FwH+I
C5k1nN5Q4LQqHbm05WcOpADws768joAIA1v0GptpUShiUl9K1zirxVYanF5uJDG9
0SYAb3xRTHk4KsEOmpiz+dXSYQh6y7VDOKGJeu3jILlIbkzRiAzxHt9Vt87UWZf+
okzdv5uiQl0eWs3vuyeBhS1viY+e7wtNUORQ/pCnJhZW6p9h7CIc7hM4P7bVL0lZ
76zrqzSXfBAHgFVOz8PfaAjieOarHFjGWdemM56OeuedrDtkUw2R4jjdPkoLab3b
fDrTgxOQ0RFCG9v/2DZrbdSx2A7Oh2gU9UZSq2zJdC/rd/1YunNisXYF9pF36HnK
7YVEG2Fa8Jv2FNTk5SPDj0a/A7XkKAIjc7m2Rg7sxT4S7EHG2KhS7ydDO0UqZSfw
6lFi+7cPGCVMQOBD5CmATa6pmKfiUl3uMMQjZKj+Yzcwi5hcbDB8Jyie5x0Nf/bE
sG/Gn1xTi6xPAmbfXVmeqkO972Z23MQLrRqFM4pU70HDUs7YKCtQxO+iSfwgy6jl
exh0Q/GTF7UKaOz4Om6ibxgI55Hs0+LI4BvQ3UmbPXIIJipclRKMl1bDe0PunvBK
Yg5388z4EOnUQC+V1N6a0+VVnzESqMxUvd4P+8MOLyzR6eyx7Qwxftg1q0BPEEgt
nXu/cv1SFzSMezw77GrHuvhJiIKSAXqOS9lAmQEDsJz294KL7EnhyhKipphjeN5L
8zhTFs6E3jvLmWMq3bEa04tk2ZAC90WREpdatdBheP1pMpAXOfqL4MUojmQBUkPU
8pLU6RQR9gLyEijg/cQw/L2F00xZso7Pww9SrBt5mYK056myvwU8PznLYs48Cdb1
d3/h9XVt5pNLnLhc1vkWR6dfuIvSV9cyhXtC9IxShGYbgsgOv2+dj4amLer2/JSp
clpH1aS7bLh3156frGL7zN3kT3j0nJSVvtzqG2Cpo5gbEK9fRTpTb7BbL3svV1CW
LoyBXmArEnFjlEuDg0mUslmlvMP4gUw4Aixg9LdUinpO8tvZdImNe5VcW3X1d8qt
QhwbV1Y683Mthvo9HESdS3MDDxmO2TMwGYnGOpQXDcqHMEJUSqHtML+c6ZP4nUaw
zWe/UWE4MzIxLlzgqO2VklklmkOYyF/GVl0plbXbpnccYIHd9nrDkRuT6qchta46
4hrLk582+rP4YInsDMDUnNUsKPi/I2pTVC5MsAeftS+JWuIKv09+hVr9216A7z3b
GLLiJwI2i5F5Jl0rYMJ3EOz/DFgi6negNeAwVjinZY2AVfHlIBaQ8wlRVYEpWe+a
gktRN7B4sblKiOF3/vpNVb5+GBl0wzgzCam23QPDN8hd4vcd7rskuYUJQAlZcKI4
Oxb0Pzm3x2PNwSAPz+X0xFg6xB57xuhklMMraeRhjuoOTX62HEEm3ynPle2PUs9C
+w3uTu5Nsrt/KqNqR/9uZ/S9/SCHzmWRMXqClyB5cWIEJwdAFNmTm9KrGswx54e/
PXnwD1yp/IpIoUptpp19DMURUQ6oUg2Rmqb4+mrxOH3GaLj++5xpMUx/OqVVxuYQ
Z1gfs+gEtKxWYxjloXEGhyqOal3RrBEp+IZoR/vZFvRR2/H3v6GJdmnoE1aErp9E
RruVi8UCNx0sJI+KqnpBrz71ZzFKtejB8eh1zCt0q3bynMNCGFyMxnASszsZfZq7
kTxlcJXiKO9eDhrHDeO48xav7PgD3oEAS7oQZHluO2Nlvo27iBZTHMo+w47VoZWQ
lWOV51ayIDtHtlr5rW7C6E/qYSPx7+HqcIHjhT/WDTZghfATaF0eRuO89tjhElMg
uGl4u6LaB1UkvO4tufj6t1WixM0YI9HNjmBz07CC30wDFd/9+1MYszLuvk+2yrTD
EmDS+XLYt0F7lsnJJM5FXE/pXHiiXcfxyTw0NC5D8zRanKy6kOSx9hE8O3xIgdiD
/mwn6Hr54rD1YCof6HTwETy3/cf4eeE/h10FJ4U3aUYoIG/3of0IZPG3B0rk7CRj
elax34IrqmbPRPOunRUDLKG2XWZg/zhcrCMRj6NjLVIU0R6+agP//PGm9H4P5hGC
hkvXJqM1kY7gORTrZpOhNJnsAlCWasymzudZvkTJuJkgDbWhERTnzP7gP617aW3w
0RCsDSDvD6ih3Dwg826IciHZZL4OYJ3oJ3zmVSa8gCWa2T9z/QHo3/9bg6O/TvPj
ft9RAgmWt8v29wVmluvCQ2V2MWPtJPGRuOxKr7BHuoGBSmZ4iToTbpvLFpVR3GIc
jzbIhhlyt0vwcUfpPOoYSGAO4z/K1RM1tIPMFhYV0AOpAC0zAN+h10B1vB4wqRQR
Y01iQ6i+mLOv/DmKD00Bs+ufdX2Uncr7k9ggh2r/5DqeD7mbY59mR1NdWJNagj1H
7LkdLQE82BjyG1s0ELC4Z2iAahNds/HPh4sqWot7Kr7A17vUc6hcx7UwmK78nBz4
FUZ1pHu25Ue8hVQAQG5e/8SYALXh0ve/8SKBL/h+7vFA+7QPH+3FSJIDFQwr/wJ8
xsXGhoL3pTOyFBnJZlwRYggBh0BT/amZhRoP2pOLfvSvwXvQmhAyzsC2BH/OWzqW
eCXTxBUu/m1qj2RljRVP2p3JbeTFkNJl/2ONPanpZ7Vh7+xYlWZUAf+KcZkX/pn8
RaEqcXiz8RdpfIxGllxqWvpMPNbNNc7ncifp696hI9lEZMv/fjny2S81ZNiHGv63
30PK5U/oEVPrOm/VeKz6UW7Co+dcCapXL0+dLDJsW6KR2KSVuZevGAIhFZHcPrOD
Li8bb2c3X5b4QTNEZAVyP+gREHwjm/mmu699JgwbLG/h87U67Kl+xRjKLX9fSPEV
oaMMDxmcPyb1xirCd602ORUCALAe2IW+CNaDCNCqENynj8j/h6ROMvl/Fsx7dXGh
BmAGhLegMZhhvRQ/Cvl5JYpEoz9E4jLKkXgPVLva/w7je0ZdFBdK4nwzTtDiE/1x
jzvtkHPRpv//u9wX0fSjBQmsWucoiwdw1ii20RKkUyCsrqGB8ua5QeeFFouduKdt
zVZzESF0sBJET3JLg7RuGJvsDpp01Sy5XhN9dF94JEQQ/dWhaYEzpK6tPcJeCHLZ
Tm8NN/ZuNI07kbEkojb8WEYnGyICvAHPWFHHhJEwQWgtJgzvlt1bBumpBjDlUwZG
l+F0gIgWgMGfy7b/uVdQZYz6EdcBCixboDkO0C1pys4adxLKikQfxkaQPFhB0Mai
NjYI1Yxr/Q8ecHTMKK3FMAEHRc/MBYD+9JHqB7zf3dZ7lD1WS17uuoNByo7kabOu
RUBCMlso+xL1NQF4fkSrVRxB1XA7ZZiMXDovsAI9vItZE54iLUoP+hGMmqx3PNJD
sJEqt3E6TASy5ruKaHy3DYBHajlpFvNcWPr7Kg/nEnfxFx+dL4qUbrBKKlTIr8yF
uYrwpq8BrhaFLlF3fyxHnnyrTiNVKG/7I6lMmvPQ0Rqt0VBO43fzDGdRgK7ZMNcs
x1pYgZ6TGbsCTbVqKYEqvSs95Y+2nGe6YOEPVZtGvBfEU6CpLcy0/Q2TnFm8InpJ
lF4Y/tzqlQ7uFX05teBwYTJ44dZm9AzFDAhta1wXb5X3YbzqiZIGTHM4/aWbBNNW
krOAW6mm2cnbcFuDmgC9siJi81kuJMcgaxEgfSXrRFh++BAq2A3I9jXtVcH1WaAU
Xn/ZzmfH0HNrO68ETNBYDzvc/FiCMntVm0GUY8aeS8IGbJ50blwsT9/mmG+8hLeU
McYFKVgR8oDQD2JcpmD9yflxqDwvlf8kc86nCu7PiVvECOB5c+rcXXLWeZVuNFif
1PmRl/unjF7Ly0PK5RNeIw7U8OOSxmZdXwOqXCQOYJuN8WAheLBTFam5yAU5Ddjd
BNu06V05MX52vvUiitx4cvFaM6Z3tHGNKLq7YIPi2+dmilPkI+rqfYruNCYTHDJ4
I3XnPRY7iKE/6Xt74jFsKilrO8z2EWTDXC2iBPqMXPR6wz1rSd8DIZWPSt1uMc2X
Z9D5yHlV8ob3BZhCPlQfKCJdxJVivSLE0lBtk0OpeNFlO1ou4pySbLCn1Hnm8XJr
Xdzct9UcawZ67wLBVj5fRz3MmHp2OQgfz6LBQfvbL+quVtcPqSOrBUK3I/joYR94
mS8fZ3ptcfeKopDoDFIqVxtJiFDiJfp8fGQAjLcPQ2EPzBdR35qiFkL9OCxbwc1l
LkZmOXHnrRkUG9GsSRAUT5m53v/mIYwzIq+qBYWqQ24lJ/XhwXtkmjhY3/AUs9TI
xsP8PxiWtlsrvT+2m34TxoTyQlHe7ESGYJk5Q7cTqCVSaDHVbJnkn0hmLb4JlGXE
xjfpDxGPk12t9/hQnuowbz8TuWPC83H2eBYJIHHMPgEI9eQAwlG8eHXAirkTPuEL
JjBytUVyzN3J5z7+Gue1p9WTSnUYmgWP/0SkRrltIl8J1Ow14ZNhhuRbNpMmBMu4
WPSwXE1NH2sO8NWVwJCLUnNfEYrJlu0WARyiw0hxyDtD0jfFoPZaglWrETMsvaVW
90Vhe8F4xZPlrYvi0wWaMI5zC2h47pzQgOdd+Cu15bzNSHCNk9Eq/pm9TxYmq9c6
hZ2+uevZLN+jfFB5Ud+oEYTizufKtosPM/xDmgIihBsBoa77ICc1CrqTgb5hmKHm
JC24/N81ZxV5vEYqHhCkZ31xsVwXAzMEAFJeYOSlH5VyOQLoSrxA+/5PHhlSw6WT
mgvvbKaa2yyNyznhwcsO0aIy4j54ug3d3ZmlfLaa6oCtPMgPAsCYb0Li430WxKiK
n0rsT0Ry2zczWZ9vtHZEiCaYYxHInQ8H1Pxc0xcbjFCj2FocNBHQ8XaSvmWIfiMU
yhenv1cSiSMG5PGRyIYlixXeD8HNWv55UyUD4s0xcsJxQhSjHy6eR8PQRfmzMeba
ZlllJF72Kx7DLr/BqzCGwmxfVXhv68kRXiFzfWNVvBQcL4aA0yKR6a6a5/0a7TZV
Zlb35aon8zRAqoZXfzACukAzgPX3VtVEneZG28wbZ7s2VMI25AraRS3/If5s6CwM
3izkkkWf4jk2yIaml+Qx5xQn5reeO30+/c0ljDdVnmIvQ94FPik7bwDFm0XJNx96
IfMQPN9qoJ8ZsiLzDtGXQNHdLTDjqKMTGoLy/REGfD/z3NV0mPfph5+Say29X1oO
th+pKKuNQgPTC7Cs7mzEEl5mp5PWjxPqy4p59Fyip+5mT147sNfgMV5nEF44bXi3
Q3ixRqS2IRz4CFdzM4COTx8r/6Dg+Tq2bWW73/3GzS9OK4LkXJCuIp2WYdgaD8Iw
sv/pPZIdeBCXtlOETjLc5a+iuY7F9N9PBhec2QEub/70PFf7iN2j4ryQBcGsskHc
g3T7CZKhKkbmi4AVx+TdnwZN7YMPJaL4iI7L3HOpMSS4E0un4gRZ1hdEzPZt+yrg
WKw8Kpa3yr1W4t4AAmRBlJycbMIJ+UFIHqtKOiRumNaK/ehe0JpSd3itcGkE1kqp
RS9aWgiU5rrf8C68Y+ERueblMNCIR+8icdlnTJsrY5niPJzpbX08Nlzco1zr/0xh
zQl5HrKisHYZODsftTKsS0rAZkwuGJtP/xzRNIsr4QuHUsW5jvwBwd6NzGkfPYm4
zbH4ThvR/EEd9aICn04XiBSEKEaqLDNAj8Whb0kkkpYxxmEEwSTYozDrJ1AGes1W
EoXk6y9gg8qX0V39ARFbK0QOH5GZCktpUMMrO7WLbeo/49uhdXWNwR5Fpux6Kb+d
TQPjBJKSvRjpnXT6b2JkiOLN1Uhpv3C6j3N00iVlfY/fm2orbuxUulvzpDFyj+Tz
6UaFfiCZmPPPE7V1CSP26ZfmxyGVJxaehc745Onfx6NBoOD4qp5pLq+MwKM0guNl
0bmX6yjWiSPV8bbzCQOPxbI0NXVSRd0cmjVerCHKmn7mfqlgAwWTLG4BGVW8fPpd
QgXpeQs36Pbi3rdxtSsuLr1oThXeTFLckMJhix0z6BlD5VHrCmpt00OAiG20cSsD
EF/aqIbZyv0evnQ+pYa2RwiIHy2fILukwlSTgylkJXsCBf20P7PtHy/q2z/enoGA
+y5x5ro97bvPU/w04rJ5l8it/i0gFrsiXMsfWlmWz0shzPhV1EsqDzj0pJ6j1dwB
cWhYvG2PuBDmoSkKygjxjZDpLJ4P/jOWGLyrADUssTaFh8SpcZgy0/9h4f/Vnbij
iw3iDyuVB/3Ic4onFFLJWbKIZ081Z7ROD5Mk9K3jL44xUjwG98fRRem5kmwW8XJj
awC7A5CRrK2C5P83567Jbn/ZjFaP8fZAU2iTT/JfTERZ2cPnZ7SEhcJke+bg6tb/
bfUMGQ2j86X3a2SN2e6wnQo2N5iOybCaEYFU/2+MoVHQzLKUHx9ikXnj3+Igw8UG
/7Onxd5MnXo9jclZBkF+WCPajaMKr3PoWUodG5abnPZpKKIJ6Usa9ZiBAduk6Nf9
ohZ5d199b5lDSJ78aO9rmEBNJD+QuuR44C13JHlATGi3m5SCVZo1P365gzhyPkYc
5BWEyxLfNrCDBtgGNi2cPC0Ub2yBM1TAmXdTOcXZTjVGRsRVGyf8rDqDyVI3DE6L
QpSD9UPv/2uHmAhO86qzDQUTZZg90YFCFdy7cCBOwTXGWmA+tpQVuunps/ryNqGQ
S+yKZBbB5MvWjCPP9q9QMKqQQM1Gh0mkuXnEB/SHsSpYsAV1AedWFf70bp9q9pbz
6MkL+2vpS3/FlUNMTzmfQzK413vUycbPAVJu/ZOB2x4496Rce9uZRno9VAVi5GhW
qo++ZDOJK+w7x10eR91PIp9vXl9AZTXboSjd/awdG1ZiErkwEEZpUpHaAIqItl16
HYi+shU008vkJH0yeMMC1RGC3xfC99/gofaLQ6SMqDk7tplhvqHS4g1wihQIKPD8
sjim8k4ADOKSiEcl4wgC7UpDO9HUzApURNGnijkBnywH94HgayTXMZ4fNm06NaKK
7LZphvZi//AEvTmFLPBZ3zxRKjhO/2LwtOFgw/knIFkYgBoFFVcvc+2yHSL3o3Jw
ZiqSt3znbcdl9hbGXPUyLP33/vy8s3/sBBVbUzyn8V3+0s5iMsx9R1culKtLdpcZ
WBeWIJ+1LywAKnEPo+oEHyH/S9VQLBnvy6c8meH4idxB/Ga/w0po8FPbehEnx6fo
ekbcC3TS/k6qSU/nYZHn/1dzEdEhJG1/QMyjecbeGBz/q05kD2xnTlqFWyEcjYL2
mWQs3uh9FZ6hNW8m7vRvZRn6ol3JFIBCLgylRj0nfRuhoVG5dOKYCqfz/C3w0b9E
XgUxzM+Rrqb/iYodMWROxt6rMvkFz9N80O/eF9l+vYZy0Hn1v0iKI7Fa8XoaRnwS
vH+LMxkeMLv0Nq+5k6h5uqCD9/PUV7LYSFQqgweyArOmC4sw7bN0rOyQndM6SxsW
Z6rh7TG0tPYFQl4tEwKIpsaev9GGOio6KdKGPokhNcfq8XWZnNJZ1qAm0fGGBnKH
xSd42H6xNBlwLPtCytY8iZ8qp5EQoBtys4RlqIba5a9/jYk8GjAc9gKkvZSZ/WJB
80oyGfHlXCa+XG0aM0g0a+KGbPAtldcJiMP1lnw98dzPiYg18cRceDWC9R0INuso
CiRMwPMaYjhSmMx2OiuvpXigjZJAVysHrc0eEWM8n5etKdklM3M6Ni+8RqPBWakj
t48ndOoAoQdZJULBclftUd/AXdAti/RDXu5OcsbwDOTDtPKttVXlqPVJIgxnoogI
WCTzY961MEkqyGJjsNMrkfJgzXjK6FSqzHfdVOIKRXcNPKErC0TMq5tDS9zZKLMF
JfOTWTLdo3OrOXIfuYN+laAXtel/xs0tEsg1EG36fwiBqIwm83zBrJbb1E+plSqO
qZaz8zf9cg6meLdfk9Cz36s6GVtGs8hTaezB39WWBpUXe9LlGEC7iZ/+A30GVEG8
oKxbIwe0pDFU4HHpMPUcKPWYU10IBze+M1wY2QLgNI+AZGbzEiXftmWeqDJiC/DS
frU5X4IU/NoUYckG76yZhR3PdVPAA/R4HwHeGojSpyZV1BGQuc1T9wfnXEqt6NQS
VmVAIx0irlz8IX9rUbaTTq3YpaKKblYqvqxdXx9ZczKkQD4LNW6jOmpdk/jFeBQn
OVgXamJn3+DiDieKZEmq7uOpYM+galT44i17iC1D8yOWbkZuUCqVYWbeyZ6IKumT
woIq90opBjOfXikHrx1IQA4Z48YTQ5Q+BZQfYbr30SxhaPMXPcXqLwSc++sNrx8G
ZAUjiQ28MegJuTIwi4aH/g5xU1j6jF+KXprBHj72QV48qfBjophc6d8rNiQpZkN7
ifJL2MEVUrtis9D+yKFIIIisbds46bkAt99DO3DKJ2gTcQSGPavNvvGL0v7OdsPc
Mw0Ci/XPqVjqnajgpY74x3XatE2UpYpMJAIv93OzMAek4BSAlQUB1g7gM7U0/eKX
mLHCTNhZuv5oj9EWhcOWd+3x1ppw6OmJaXbJuPSM/MnCOsXLTD+rq5vVp0zApxAq
GJFbC+fjsxbO3e/zgWRN5KfrTj109cp5DBKy56Yh/r7dsrD7dP/G3zS/rYlVPaG1
TqBW78cZDR9kYvu3gP9BICnGBtXE3VF5qDc2rk2B3rJb+918Fwh7QTiOK16ZvZzY
1KO9CJZSm60cS41AhNoId+BdLFRBocu154pgIVderSRYic2TwZWAw2mRDsfxTtc9
yr7MZSTxRQfCiF3xjBoj8F3C1ftgQY3LoWUI4Foohi6oOHNXMjhqSJeAFEMB60rx
4TtalFDqATVREdK3RZu9nFi20VFiLZ3rpVf7G/U3Kplc2vs2e/+s8i59sDNvc5ru
hiCsij1xc5yXY8es56UTOcYeSncobvygrVf+zhLkd2EPd1XMBXsKKukJY2ySznyY
bEn1JFiz6tqwkO69n33cRAoQ+i6MJG4kemOo4nBU8w1OIROJpbJUHePZLNwBJKXa
xkd9BKsLvP2+saovvj3zTdjjCemKsh4X/uOl5hRzjsHl3Tw3OPRIvjbUOJV19iNl
iRD+VZ0QyYKXWAHBOt93ubdaMQv/FNszOShNbXiynGGIKYkOjNY78Ny8nsT+e1/L
fwWwqGgw5o+rxaFSPWHDxTkSsIQN8fpJHJjztGbgJoFxWNndgMGk3SgCtROmNp19
UCqRuzxic94erYCFVuy75f/ZNfgWK72fQUCPs4MepbZtwkIqQXktj1V2wt3KEgl9
LdUB/DHQ3g0XOpnUzmQfr1sRk0WQkXACjXgIO3sPFOfzUYkm6UNs4MjGNwFoaDsT
Dzh9uZ5cRaSVRLb1XmuAXzYwnOCMCnI3twJKdaGnt8a4K/FEpUb71J7CSa38QExv
D2LTHfRyLSjufVkkZt0n+U8OomRAtou+E14NLdvtD6+SEjAvMzGl9XOoXgXMWZHr
TxIZIwKGUyJGzvLechs0Dp8uCmh+Itx4+S2QO4cn/v57NwJVHpvFMyRSMNhYhm0M
qe5JSl4ZEZamhFpUTPkm1EVkCn9ZW3W3szQPQzxPbkrRP5KkFZfaEQHSgFUcWWv/
Xxh8WkOKbo4OyO2t+egqxIC3vVQm3Ua/OPbaN5qPSixwrXbBKHRIqPSucQLGd1FR
7qOyF3nVOA/OyMtmoXoMWgUmTbM7LU/5cm8QyFahtKjN+mfRn43+63RTCHzPqltC
YSe631q40nrsHCcM9vu/80ETLkUuuXmFjVA9C09z7k0G7lC5bpEligD2uyLGJlqM
XFMQRcUsbr/HjvW+iaoHs6+e7EjUGeA3IzmlX4KCKyTPcOBJjMOksyPsZQ1st96T
148nMK7qZLpkl4UIxWv15TX+v1RioAHuZeiUu1HD5VUsZMEhv9tB0zvy7p+v8gfh
zfEGCDRewnmfcEOZ6RM7C/ExkMefPveYltf0XCcezxIVWLe4AzayKOK8LpOefPI3
jF13Wf5if/6UKf84Os0ilMS8eRB/8RrB4vb+brx7ucFYFU8anOeWSVahgioaE0Lg
xbupmvOLJnFAzrJQyJg/fcRcb93ssyqCGmcZ1kx3SS2OamcHOj8Si8s6jrQuGrxc
3ffUMkUgS4d9vLQHWirgL88DFhDrssdI+/faPQyeBgk+Z9K7O3Yc/qV9RM5Dbp6e
6/4iievHM2iVbfAQLBIQj1Q3Au3UZagc1lRt5DAKnsAoNZzLTL+2mL0heon75Io/
LqT3goRtXtlGry4oS7DPyQPzoGCN8oS1HdwineVYyKLyuI3zW5x59SuH4+uGPQEa
BvGbPdn4QiaVA9ZwWGgZCkxSjqmQgskGX0MtHMnmMhy63Y7oy8qfdgaAPMe0jsu0
DtrvT/w9kqrGhI93qbp2DcocuAJy9F8F7CxyjOAbhhYcFZOGc5mGk41sBKeuOAAT
t8WepGL0tZ+RPJdsCuVDuRrjmmaNliB8dBaczL3rd7AhNPyRe06pW4ncM51Air4I
hgGApSY1ly+9srvGBd7eD9dG4rV276Vw8ekD4Ay6caP4gaEMvWLFJv0JA5jHZ4AE
Y5cG6fvSdSZaa+3AX81fXj1lUSAM5IjzfRnTh2SMLvzC+qaADAGAcIB3S0tgfvxv
1+9cha38Apthoc9Q2PmpcU12782hiq5dy/XdFCqG1he0GSbmuOgHZlflNazM2ccz
E+kACZHkWqgRHbMsFib8d5AcPvuoACqiOBXLmp4N4B32oaDTcvGaKWZuBT5qAhOx
ox2Qcb+kEZtejlI/ZVSdi8U7k77jrRxwiJTMhcQI7mxZvySnoKiFFeDbVm9pZmNU
93N4wjuMqRPOQZwj1HOxjIR0TwvNyRbPTRTdc5UTFcPPV8F3PBZrDCb8pqSyOSft
pnTxDy6ys5d9w7IhCN60qv9fenDu4QnLcy/FOgqD0eEj6HvFDzgV/ili+p1qm8Nq
KpwXNLWvE77UwOCi2oTNzcmckPkiWUMOTdu+KUikVGuS01z7hJgMMXc2LxNh5zD6
iCneqN8dr4PAUk902ihoUdmxGVXzlCErpavfNRTYNSBoCqc3TDnwPLRCpa6RZCYi
m8KVlAe5cnk3yk9phICwtYgIAl3DNYSItf3K7THBRFyxuAa1kFJzO9St0p4K93SJ
Kga2KVoJ6Ja4jJd+ipcrZaYYgDyj7QEhTWT3MdGCHICPsxyPNdZkZ1nU90tejv2y
Ni3K7S2Z9iH49j+uhIoPuHfhk0KCJrHlq46Qabu0LtyAYN4nzEuRhlyByH8gQguY
sbr3k87Z0OALygaOiVlSiqfpwrqWtB+pmHAUW4i71jgvE7NF1o0wrsqZBfsrXUbd
pI6IbhOChMh2BPeeVoZT8HmpmtR6h4CjtHYnf9BM+TS58vrvl3ZQjxsBExAqqoti
TcNDghHDwfae00dCNIrmRqU40tTwj+BbvzWRKpDuxIS1+hfsUUhD19hZ6lQSAQp0
5lLlCE2pMEBt4LFcAs5QM/uJrrRtqnGWatoqk8S1DlDJUE/pU6bZ6KKCmcIncTBS
okfvuS/2nDzywaoEGMjOZZTc538UjXtj5mnbLSUT6qzvxAa9/0JME3b1hJDfL6FL
OW2qRItTHKSckk/z3iSArvy/quQbwiw+f1AmhXLK+pbNS6rx1jdHzX0ojlqFRrgm
sVunw+nSHYZaUtaJFP1PzF5JQo5ACT7Iu7cmlDNcRPLL/bGmrfjakn4WiRDwwO8f
dyYVNRpvCy/4lf34QGyOMHMkp8Jrm/wGfFuzh8hE++FN9C/IFZgxHChPam3srL94
e8T0wqhhwfsYPhiboUGw3K95S1PuQH3LgAZsjj3V1/qDMiu1CxGRQzEk7vzGSQyQ
cwVrprJfblxdedbv7jpJLtlLa+kOp7edigCtotQPSCojDwE1+2hWpYfUC1Z1eU7I
W7rrKHgtcGPHrH9W7DytR1oSrM23oHDF88zb9xfQtDVLgbBqH2gJHnIbVaThDpAB
B0TF4ZwnbZwKtjKPlUi2eID8CkdIRkLCR2uxjlehTKgVGi8f52WR/KlQW+DK5CbZ
xnAFQe7XaAJLcim6JZ4TvQwcxnUUkB4pWyXgmFgHi1YHEARsRRSI+XJPW5cM8zkY
a95utdh1Wf8bl4mvYiVXjyjSa6P0ljY+XzTCHzKU7DJ60I0WM74bdTUqVeEiBC/R
yb9uUymS1wYC8B3H6qCF8s2cVpJruulXiJ2sgCNF846cF5mOlpgGi2aYsLo+oSEt
sjUlsok0ZpHR0fqub/gEQ8Pw+En2THpbO2j0TNcOJhrjc0hdhFEqImoKyW4OtG+R
5u7L9li44V84NE0BcU7qTK31VwlThtUBUwQ0gvdmLwMBIvN5MzSZaCZnYMd4hmx1
A7PWXkAcbXVOVZ+JPRNr+NMnSBtnbh370lZkrRLTmGFLuSM4RBVQ1VXTODEWugSX
kovtntqOOzNSwMFyyDt32pRJwQvdw9dC7J0+HeNfxL85mXyNQm20RaX3cAsqHK7c
jnVD+gj6fIy7DOus/0INnZjQ16LHZJt6Q+2hVQvbOMM2lgxH9BtWvaNoNKHlgYRj
h0onQ1M4TPPDC17hhELG5+ESpUbUsrnKBS9AlArohWD9uUfUOi2qVisBSf4Zro6A
QNe/PqLP/3lVz5E3eno5Ll9HTG87zIPX9Eg/fDaTrSsegixw626UFNylO+R99qXa
PQN8PQH8zmPLXH4w6NZvAF+R76ES2hGfRNzjeKbJnoG8CTyBbvRb2uqhTH94uL4K
uv9xkwWCcnhIVjq5XUPX4wSmSw8E4FkUDHBB1G0UPZMLSil9lQjOfzkM5qGWSOsE
a2gQla+Bf2N9Tv5u4bcfTDlFjontc0sLCmVSRgKtjio8Qg/wGotx2Zyj6NxjO2f3
0ss6gVmtzk1d4ZHAKwW7Y56mfFPbOtOKLvMi7OAFB/Uxblm4Us++83V7Ye0vnwfW
k4IFOFgeFEp7vL5MKx0keh7n54W53g0SJBsbDfG+x5c=
`protect END_PROTECTED
