`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKKq9xVslEHcxFKahX8/cXxxmZW4Jcvjw0ujo69L0nbq0RLxqW592fCdH9OdyWA5
PT6IRqTdS2iB401g+fsu2w8Bk0BAG2C20+5z2dWz5SielYZzrgImamfqakXszvfT
ljPJP6/nnjgyG8LzDs3zu10cvkkzEVFKVlUwWoDbRiVL0716MJYKt4Az8RnuHM/M
FvD72Y6H7kqFSvqO7oNZC6ArHfskSMwf2cu5tTYbS8kx5xm1hDk9o7SvskdA7/9z
G3l9ZxJXXc537xSpgXRIaP0R7U/gh9ga5BHozKiZcfydXXfknJH2A4cq7IBWuyD+
Iv+OXwzIQ4dVkvk61+rFe00rUUqUQSPwBAqQyCH713pFGsjwLdWQrm413RJS1qVM
IhPPreZgQWRq1+svraEmkSqTeOQGa/KuVpUZBD6EmN4mnDnbVH0k++9PSoiVEaaA
dW/N2oPUjYSnNthUkqMc1K+W0rT2KvXIZ+mk8ysyxlRZ4kT8594xclDDmxKvRBps
vlpyKDID0yI5wQV9tOnFzomqBab3n1gIqADF9qZmabY5dINptvaXgoNpcFeLbbVS
WshO+68YN3jNDSkXkFYpF3N/cT2EPaqldHToNLJsCl10m8moPxq1mcht5F/mc8G1
w787jF7Bva4r63sJ6eaJ0ONnZxbfXW7petIs5kNXUhB+ZZGncKSyFblKNMDGDFdC
GJ11kIMde4quyi0HUts5a3TM/AkWx1yMcfDqtZgqroT3mBHePThKtQbHW7lANGqt
kQSRoZ35tGZqxsAWVFGBLSFcbh8+lgjVM27ju9pqoxd8+U64lA30LFwDK5xbH9VW
B0pMjvcN+hhGrsSRPHHTNpNOD4lFdxtv4Pw37CzxFn3Y4f8FxeiEFCNuJCGwbjKb
MKL7E4gSPodYTASOgmgD02Vc37HIzwTXisCRKf5v4lmCmVNY+kF8E6Z6pJfuQHRj
oKarlDX+vxzE2y2ZYrR8v/KLI3dWhyVlsPCS9l3+zbIBHz1uZtl8pgxe7XJ4S2yq
5AmrSfEBcZqYjHRMPwQfPmlAi9dLNdAGt3FnCPMi4JfgGXF+Xbnd7/fM+57j6lyF
PysTN07QPzj/k6IWV8oeXFEWxEE4GR8Ph4InTcgsHM0v/bFswh9AgCTjPGHNlick
hGtF/kAtEL5Dz0EINEbB6Z1CXazI8sm9ZLUlT6cKkikBTLIVJzTzg/393NRjm0C7
AmpMOhYQHvDE2IeGhDHfwAnXJBKAnt8HN9jmp8Pe6UVwiEQSUnDBreDAHPF0P/1K
W4ePSoVpoJ5kiL6+DMKu+w==
`protect END_PROTECTED
