`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W5qKlobjXKAp2wD4HL89TMNWl34xmDfR/pEukPijcyoldiYVKREqNy02V2uAYYdv
UI6HEzxvpAq+obMbp9x+8Cg+5AXC8R9TAZa+n/FXttjoDarJZpcx0cgdzoIZqAeq
JvIZhUhyFEICinQAuLQZlZKBbT2gXFH52Ci/SyLthOn6KCnNFHL+cVnrDTbRsBHp
pbAkpz81b1v0fvC9J4Amb6kYzlXEgwgjAqXO+3R6aA1fo1Se5p/7pyaB1qOvNGwO
NgPqxq4z9RDk7yR5P1o+HDNJTBeN8hCjlGh4hgk41aeMVlINNTNfYU9N9oyXLTOu
FpvbVd0AtgVEI9/jUNXUPav4ttSG7f1lOZik8CDGSSeU26vHlaVQeG2xadhJPFpM
knpgnb7XC1eniq9O1qqV+HZeQWTA25vg152OLo/ZE3ePdjNXpM4rcNrNmyN2LfVL
yFZagiTwxiztzu7xGQAS2worag1FLhTqGnNMNz2+DxTz2oQJJL4FmQw48UOJdYxn
hTiR0sKl+GVfVpuzXgoTKsq9P+yzCVJDpD5k/ojLyBt8HTzKl5tCnp7FNJ4JTwPT
OHWdSd4H/UHmJvELQRBMtYr1rJTi8m9xeM7sq4CtYi19YxIPq2Z5cxVzfY/CuoaI
s1UAfZ3kp4wUfMC6rTsfbys/mYr60NiPO/4WEzfbfcbCATjaNFcOqiL6L7lThDkF
C+/XRqeTKsDzgL9Z92hW9Vbn0oC3lK7acK9uOOwdu6ClrrFkr2xOyYi0OomU1MIy
PjztlbGWEyLzFqvNcqMqmFTzwQwjmzyEdIXN9xAl5HGW3UE8j1mTKc9SQ7DyG+y6
tt8Li3XhKgC/lSKqaK+I+ByV1HvZomss0JGIqetPTeFnCHLeRxgwPEa2TUvwUPi7
CUBoW4AZWI8fxRjAS/kmOsceMva7AEaLrLWx9jh2pOzSKtqYN9HF7i7ta8edLhlf
RsO2SMNDDU2FLXM8d4c/QoZ/p2aZQiPIl4VGXlpIpkdUETmFo7tYxmoNXPDqOP5X
K9aLaOfaO941iG4otmBiIoCvNhlCYlo0kVukPj3kpY/5tOV+Ru9gWoN6mlwPCe3R
HAHEkg5gQe/IPe1yedw0WBirwkSlyHHCiXemampkLUD/477Ey88BDvjcKLTqDpqd
eZlXIrzODgIz2O/AceYH/ngaH/s/KAxxQn4A5xJlhqTRBEN4s1BML1u9VO2xUNql
mjZATT/XfrmNdU9SRPVz1JNDosK0Y2hrQOOWoaz/4qRYTV18ElryjN0QFmv1RxaX
xW2AGqH/ZLMu1npw6C9bYGrPCNcbgFXLowaK6MUV4xg+QQPdYjvWrGX1OVMb18bU
422QMU4AEYMACQ3iI/HYZQrF52ZhEXHr61IUhmMMbLx7iTPCGJ+B8xdIBUs0iMMp
Mb1OmeIRMr5FrwWX+05LcSYbbfIe2E/teEBgosG6RsYLdkXPcAjGaMSmbdKFQdy9
bUfusg1ComipJx2LK8PFPGi6nBUgsSE/Kid5aKXduQFHqC1WExymWOSGYvo+hAgP
erDflq41k7sMjh0WZcQKj6LYcraOcoxbwhHwJ4bBAi90mLiEAl1Wxa2flSVqjjFL
4YvCeFAW+cctpMq+KmG5LisezH3evP8wDEILGy1mMdD9NvLpzYVO4Gm5U1wCItdy
ANNHXekAHvxE6zWxR+wo53UqKMkESIp8sOBN899cy2U=
`protect END_PROTECTED
