`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYMJXj8JGwL8X3XDWqBRXdaUWQCkUHDmz8E7e/LC26Rr+wnlLGWSp2m1k74BDdBV
rzovwWagjfsNQyuGUVOi3HdgFoVA43QCokYivtfZvHf4AJ0qWDDhqBFz6g2BVfP7
Jng/i5W73gv1bdhSaIbbRVEd/TSz3k56q4nRNcdXY5lXLWFxppAMjQSCVNjORn73
lcCrWNlr31Ho9xGw+4t62V2LnvCVY3e/UJ5R4tXj5/YPlJwdfr4ts4uLXsd1qPWy
or5WDW0TJ/q1Vlz7a6WJp006T+DJJTa4HLXi07jTUaVIWTuCOBNdQ+QAQjGREaxx
pIcy8Wjctitso/+i2DKaFlooDph+Y1ee6ho/hofMUJGSqysJxA0k3mHdjSwN6ZWv
3kt49Ob9gAbTmx3jpPr20iuyvFlDS6bQKUirvQKOymErFN8iSGKBr7p5QT+dNBw+
dssvLGgTE4rR+fcTvZIbSy1Os8yWph2Fjf8Ez0KxoUhgzNUh9S2/AFCy6LTViEzE
0W9EpgWXt56u47er0gs+0tl7zGe/V23YPyRmMkqCnQ6DFoXXq17kYfLrfkwF2gAS
WSQJ+m/Dn9qPtA7LWV8abr47HgZpsmFpH+twFu6o/8nKs/0TJgcw0G4NZ8ZoxCbH
RLg/N3mCiMunkXYq5I9yywOFxxK/nS/GLnhTZKi6A0hBGsqKZLt6QLG2fjlFR8Su
yaV8/FqCmCmyGuFGaq3i1/XfHzPnq9rAPjALYL0Toyx9Fucw35pKeUnnPVwZ0Pd0
Qe4FDJwxWV9O4GizlXYAHKrmIBteoOGwYUGriE6FTYTVIPheOkxywArgIjuKsEVQ
uiNaH9wMMHdhppOFNPstwlvfhsPGWpHRAZpSP30jx2FQcJDFu7JjK3gCgDgI1DoE
iX7nxFI3Fo67qCTdrvskc7XDRpJojSULR+oppllGggYP5VNPN78RQK9dmj//35f7
gSrlJ6ZK+ZREjQcNlea9SEP5qYh5n+BYmU4rMZxhpOPt0RTAgAZyUVfOmGBML0Bl
9dt8uhYyvuMZV9xszwbARhu5gsaDyIw0xkD/bMJ9T6tfq8Q4D0VhhvOX9MNxZFEn
TPE/q1cKBybtQhcAqjoCDxPnBokfUkSlmZN3IRdlk+Q9AZY7Rf9VPbZHmNZ+mQKz
yQzqjfc9PGBoLKKCZxFP3y1xIfjIRJmfcEGMzNnoYVyJZZw8u5FpqDSk+R9r0nkE
NGJyOSSyjrbwP83REDFDvLdSyKHvkd7D9AFZ2lWBhYHDRV9RRaVkJPhaO5mTArN7
GaZNPxMxJY5XwmGWWnIvZFhdUdYOKB7hKIZr6wDZ2XaRFdMbGhrjSIRIOF+YLxj2
ayCpqu0E2Z/vPoKmYAkynsG+Pf8z1n+aQoPx4XNjhvlIR5qjE1M0ZyRpNlYLJTPl
o8I1Gtn31iK/Uvt58xzJVYJ51sWy6svVGBGXEWJTx4MJVIB3CZH10bihiU6WPvaJ
2FUbdMzewpnXA43LYZKaYFUYEYqHcFWAlA94B1pPVQVWNHQYMVUzVHDl8xR7ZRZq
dkHbIqDvOt6LkxHArvfEVkjkikshxNv6aF79VwZb0nLkDe9ZlweNwcV3GtW4aNNe
dykEwnEuuK2B46FzguLq4iVT3XBn40eS0fDWFJCgRtan0Vwq5I3lFz4hdatlJwiW
YDIoeb9223IYmrPhpxXmQ92Io0T4gK8A8335vU0VDcjRmh9N3m0I0+TlYajH5pmU
bMshgtExIv/2XcTcba2eRQ==
`protect END_PROTECTED
