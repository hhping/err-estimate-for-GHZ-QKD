`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCbLHQ/eiMFClYvjx0vzYxFmHzrvTkHilyWeQqRUfzaEwPhHpehn05LeGCY3Pndd
0B+NeM/xkDUSPfz0tpGr3GsoIJc1+pNqi9HCJM1weVmtpxBDJAo1nvpQyCktMFMR
gkfaHPhiBFXo5dQIPbsiNsIO+VnsS/UtCOtDtK2tGhnA3X8suGAqNMPwuaRBvNEN
0ZWDCj/TtESB6Suu4vvTxF3+/XXAgg11HVPmLTsLrdjj89RXmCDFhzGkMAINWBCX
5E9Nd/9v38nuTEy47x8wPmXUSyYnlRRFRpYu0WKmpqTcJ2597GwFdQODuDoTyLOD
nyq1iX6RVRk1CyZl3og28ljRXSDWY+VSycwIwyA9M7WAYyvUxsRq+P7czxIPFfHS
xh7H+jlbVlemHi+WgQihdF8KXJCMJMA5AxeT/1ZWd4SiU3UV6g4zZOKzTs7KpbCG
oPaRi+lonQFhlHrTNoglh6xUu0sECOzauIs741yGRy16G88rpG5C/KDHEJf5nPut
RH82fink9oAs+TO863Pa5jyWyml0LotJzKhizR5UkggzAXMsztIpH8WqJHpIfXrl
wf6GeVKnan4KcKS4fS4oWLV2bcy8Lr9W+jWWRPfJE33OP/Jwp1aAMI1KoSnZPwmD
Cwf1Hn9gvrnuK22yYqZ4XLH0gPFuZ5vw86sJZXgMf0ENdmDtMxR1HPTOc3aJTutP
3nV7phe1Vn8s6DzOshtcdTRAY/NZPA+eQJLOPbBAJUHI8XEnVjiYRbFdptvC9cKr
TPEQ9rr+8yaDGyMTuxnRm2gOhuzPHfxXzlnlsDn+KTeZ4ebwo+9pF5kJFX4F8HZQ
30ckZI8yD8K6uPD/wxzKN9fVVqXLhu0qRFPsEtUy9wucveHtYX0lSwe6SFCRuCeU
iPWAsV2Ecb64ebVDicLfyTtX2mD57r1bn1Mf/doIRgG/0jXL5E0LY3+Qrmtme95I
HMy3ZImevXoglQjzEZCtI+t4qy4lTbLWOFHYCfFEHI6qDuuC9PlDjq7GRSPeYXrv
hJAChHuFPKOgBx5T8PfPkahzQT1CYDnEMWMQmFbPdjNNvAbdWkX26gjsUieT06xd
erOO9PLpZBj+n3UguZJqF/MYEta0fkOXqkUgsCOAaMsuNVBWIH0cpu7zC1Sw7lDh
ikWO2SEqPD5hzrKVA1Zidr0n9tJYWEEeQw4nuwHxdaExUOX4rxInm4kd3YM+mrgR
hwbSogboZU0h26el8NSkxfWL5gU2XPIwSYsHiOXFJDCdo9aT6hmEOrTKzGrq40I9
6TkhyuhKb6MtNMvb3KjFkkbNwfHRqthReYWYA+TodpWAc743v/XY2fo7XLU5qnnE
q71VjOBewImTxgC6xebvZHOQyCCWlGpPFQ5rIytRuTbKJ8Mc7l/OLurKi0jmZLOj
PPu/jRPub8AN4mmdeSEde/4Av8HlIz76Gc4OpKLpydLOEXO/lsJwgoxDXnRkLnos
a2i3LHw5AFATiOysSoZqV4RxP15qXa0I6GN7bYyurIBp4mQsgEeWFQsEnt9He3CA
a2f8M6alsjhGN/a62Deo+e958sVolDPn+uV4naWAEQ3MJknDaQnYJlzwfHP5Pwk0
7XbJtpHh9BGt2GUSHisieLQ5LqYLOuVqa2xHzE//D8Ef5kOwT7yih3VYtD1wVe8Q
hw6DyvC5xC+QLJ2289tR8LVwfRSOJiqGGiiQTI/peT9yxEEQamn1HTD7crhrKCze
pP0YJHIzk3328o3B9pIukPRr/vmcb5a2gkK+r7Y3iRo8hegeH4AcME9CEwBFqmk0
sH/rFriIq468nOQnVgv4aILd3wkbM3W3q2Rl1QVJRtS33Zzkg2qU2lvgIb1FCjGp
bwmoOBj09yJwJe01meFOlG/88bhBR7GnnrnE1C2iyAHSvZyFhINQfu5FM/NpTJGp
9BSs5IN6FkVbVm3XYFytgn8f681HvNQPS+dFjgZf8HR0SMyHmRT1bvrqK6LjN3+S
LpeXMCbZqWlGrRdFcAtctlm+ekpuU4cvGpO9ai3yIW0LLO+VMYX8xJDue6rfWNms
HsOOKPBCMmZSE+BRA4/3r7/Nrmq1SqynCT9ZVwBy0y9DkGvJHqOnFLUqNxc0j+q2
ZjtFS9q1jEGhIK78LV4EI+SXBhcJ0axPNET2mBmbrq04byTI3+NTKJce+qtwqLYi
lwe4u0IBtqJWptJUzyDy3PrtbqwiBPnMUMJQXUX8eyxLV2WUmQ80y/3/SGcdP6Fb
kfhC/lExhxVO0XGRoXVnXGJZ/WYsb7drjmPZq4nV7XmY8hJxegcviuYzJcKCcen2
r07LRI2V+ZvI3gLsvm3CDxFlMW2kz3DIgDEVZUUJAuM/4JDej28ENhzfwbQxAA1F
yiVwBStarhv3rVEJTczpVhx1fSWfQ8nxa5uN4Lf8/a+rCP5fK/5ssgoKoErKDolD
/3MEJVQhkqOrvH2tNpkcXb1EuyjNqE9pgIRASDSJ2fcIg48DmXxbvjLySCItrpaW
DN7e1uE08xWAGQV2AYWVDAdYb3othn9tBIWrbDJam/o5aG7sg9aHKok1eA+LE7iC
NqziN3nLqdDnokMfiOV0H+TSVf4tADccRojhP3peNPZqrlxJU8FluM9XjB1hSi5f
+urtlP3ovXhYFd7b5XQ+7vgxeLqNQkzCxtR9NyVdK2eKJif01yTd9G1bTlPzH76S
IwtefSdqDSfWaA44PdFZowsxgiM2IBLkIgmCFn81zSDgiaWT7H5IubdDCm3uF9hB
WKV+8zg34262X45q37L0oqcLx1Agqlf6MG7SIDi7gNknE8SSxImaItCqK5y2c4AD
7wVIPQfK2vCKcVGZ+JTpnqZyoc/uaY3IS2s87hsYFtLtqnro+LDJ5uPTXPBdIB2I
dZajpRvBwVOKRkyqIUCpZWLXa18LtQkc54VCzqHZbUSmb3d0TpiVCKVynj3/YVJ0
JrIw0RhwicVFhmc5+EOxEMj5/d2clIwa04rNpqh5pnnUKctRXWnPM5JgaRIcaZxw
nSa5nGYeco0s4KotzY8TyKc52pKJljHrS3ATHCQRFdb0G6xr3Mqr6zjuL1RiBI+E
EN+nxgDWGsonQI6LqHDhmuYgxkEINmEy2FOjIxh++JyI0RB4aybJYqFjWaW/h2MM
fc7vjfaJqYL6pDBBuekbqfGkDsU6Nr82u/WL32W2Ir+c9vcvAgKHLRaj6OzeNxs4
e5cgIzKO2Rgfxd1Q2Gf+UrE33yFjmXw7CeOlxXpZPGdP2axkND1CpV2vocftHDWl
WJ6rBQ+W25buV7blEaD1kqdHf2aySnzDWSipvoRAl7bbcBGYvvSeTDWDM9czVTR9
YhokLx+IomoAMNEVqX0TNFzd79pA1ul3rRrS6JBMwmn6P8jBrlzT/qd/pNUSSXWW
I0MVH2Tz9oU+/dDdMvVbufTyHrQYFdi00dTFwx7o1Rv2zFi3hBRvXce/Di9E8JMk
83n23xG19auPGLYjp6uS1JjGKp6zBACZD8A7iBr8dyrDNGTCJeMT5oUY+wlBSG8t
D755Y0QIKwCXrYVzEQRgVCDSPstm8tjX4Kcs+d6rGHqrumBBUlYqswA96euvmAPG
5ZJiXwNjhDoCwtALO17MDhVAO0f8PebMwK+kKPRvQ5HsbcQIi5iYqs/WuR3+b8b8
a62bT1DUoA+hWIKys1DB6Qdzv07O0xjYba2yAGkVuLUf1rK7Ic6JuT+dGXin7KI4
mwob+zQhb5tnzur1PaKNLwkWMHfStxsqrxLDP7chA+YI71eaKoIuFb8k0Ea87Fcy
u0ZJ7r5KUlwYd+nKJsPACyamX99h7JaoepslfVXONig5OT58+RZVu5AzSbL29pWo
O4vx7kjWr+h61DDdqpNaIHbnPtqlb35FUAiq6Uapcc56inrFxhdJVJyOs33jIHx3
jliE4n3+hs7MNoUxW61Qg9YbbJ2n9JdHOUMk1JWKy/7VMkarAsUJjySj6LsFICAC
JmJq1nMxOgtdg3z5FEmweRGE4IU/lR9cII70NGXlHQk8IEif6MkvUE0qLru9mC8r
h6Gvsb3iu6TXX6tL30nGhCcETsBVC7AhV4rEYNTVd75tNYWPF5VG1iGVe1crsTMh
xPYAp6a6lxUL4a5hTnYxOvX75m4BQC5YGpgxkN6jHIJaSpkcUjIaGsHI1iEZKKbZ
bBma0BJmSmBTMUYu4nLfWHTrJIGFFxYB1XNB34x0Z8qnR2h0Z0elbNS57zKS7Dqg
SisnGDBQ4gI12Qe1MKhOdlLlCqSG53bQIwW3cg7tENdzIDqPKTvCuR1JXbcAo8pA
y+r2nloQ0M24t8AZjg8U1Xp+HXSujJPxtb+0Gt3aXe5T2Pzq5eIJCFtDo2djzNl4
0+hs/aMBD8/nECcAIkjWiO29aPAVG4Yg/0318fi+jY/IQEsVPX7YMejURxjRqpd3
T0NmnNU+rRd/JYR2j1WVNgakAogpVnLj4ecL/IqCkrJPdjX/82PrIBK5BqDMrg2j
RAyhHvA+tAhHQ6gOm0ZvPAkCYnjUcyaO6iTqIEEOznkohh7K94LbBjPc1fE3z35P
yKr4FFBMljcSS3w8iVq4dWXMiUd67UgPp4e+F/Znm0V4WUUtFTYv7KlQecvcwrQp
W1knpeXxGCJl/Gjaed+BBogLS+h86nyhGxpPkTn1+k0=
`protect END_PROTECTED
