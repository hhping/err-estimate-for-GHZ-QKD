`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UnBCG99PK0fod7aiqnDs4jCS9uxI+hI9wL8JHECYcTOOZokPkkXDFUCtqqhdjQo3
UXRLZ3FrHbEa/GCVcOnUTEN7oixnqQhNRD309uokK7+nu3ad4iFyyQ9g0qOJPRsP
UH0Gn3JO97UbMQRxCHBo5BcDEm6t10gEviPB9oyePoOOJz3KDQ0y4F2pe9H1pXVa
UIE1gVPqmp6Re5+X/0ncxaSnTrs7bIlbotIQxOfo1E4el0xxxGvR8WB4TtvpTbL3
fChk3wHxa3BQeHN5Sk9HNE+Frrzw8atslNvt2NQcFVRB8U45FtXoUxEu3xIaIKsT
ByyZ7lZOJEr9dkwNaB86uCIkK1FH4w9DwZk4ukPySuUw3bW4HDNoYojrKuPsb6qZ
N5j4VUGHDBpLN3KqhjNe+Q0gKcr5LKLwjnXJ0VQSoRc5JdzbuxVijhlQw4ElNUXD
GBjfyxqTA30z1ioMlzR1WsD4BYPeW7ZQ4c8GKrNwhjyVbsmFHCm3/dgLYGs9CQIz
g+dt/PdAmq5obHVfFxh4GriLG8U8PtR9xMLO4UvYUeFrkft9t42e9X8rBGkViDd4
lqwVrAhNPiLBjulVCk8I5zo3OAdRtASiBhPDUpitr++4kPOxEG2sxU/oYSb0wi1e
pdoxiTWTF13wGepeveNnFTId21VC2Rud2dPojP+G8MppvOFxnV5trulf+4OloYey
CFhAoIZ59zjNaBsvwZk3FKx0QOltiMUT3ti+lyJ+lJhAb2+FNZ+zXnwj1+j4QjLh
N9z/iPXl/x9e6paw2tQEvw==
`protect END_PROTECTED
