`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MR75PuP20J4veJKEcXxOiz5DI68uL+W6aEWtjSKJsIdj4ahasPgZGVLRRBnUKREg
Z48pgbDLA9f3JpYmrlJBPKWlSHAZYwp2Mq2YZ8JnZjkLTJO6tOHfpUnK+hXBEzOh
q2WkzcXXM1qy+tecOn087CqVfOrgY1jaMjpnSYI2nmFynKMIe6tw25yc9jpFQEuO
Te1Y/FkhcnBuatHdqG9IerlWmyUzPolUQDNZ/UCVXnJpVYPL0ST+7Xv/vEt37C4G
hDpmhk3P5Ubzu2shcyF/WMu8Vx6HdfjFNrivpxv6MqXVgY7lTU91VJeJ5Z/mBGkU
e3JB8iUmrhjfAUtMTbyokFcvL8/JdkVhoTqzEGsmT0OMbSeTB5BCgGu2L6lf7E2+
jMDPJn4EpConO58O4MWaRLNS2eIupbQT8W8bSe6/cRwkSL2PodaY60tbJHYjnPV8
EH7sxqcL42fL1xoAkggfeOBJzMkQrbU0TvlvVDgED/w3HwcfZoqDcYfuHpvbrmcP
WMeeuODkZyfHnEisQItGk0cCDpdbhgwmBd4fTSDPqoQcJeO8E6obLUNrvMxQkZDx
G63jAnlwMaGA6jvSbDGqTMqjwwf1SdYc88CqCZjvnUdzF+XC1WUNhLz9CfDkUMwl
SmHN4JnhNnFnZQCDugb7h4pGFegZiiCWV7O+hFIpAlVwaxtMgcZN1zcndLMTZ8DP
bqadpW3ebJ1SFo2cxHhLXYPh0RzX5PkW4tEDBZEgQgM=
`protect END_PROTECTED
