`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUlQwswqdYCzxFy1Iy2E5eC3Rx8K8nZeXXYAsqQBsEJcWgg0cgx3O5cZILLj23O/
EvlIzCOUb03BzvvUx9MqlcF2d31msYs+n5PpDREkcHOcARgH6/OPp2Ecl7+1HQnJ
cbpD6dD/kBu7C30siqyIjC94AOT0snbjb1rpb6uWUnTkPAVjRRiKaBLfK0qD2nXN
46pxg0h7EYqHIezl7zJJerzLmGWbLNa5x6ffKuj4fRX2HsO01d68OySjQ7GUVj53
u63saaY1oiHwODafiCxagB3+DVMkV0NJjg62n5ib7UhEy53ldS/0XAQt+wjbDY59
fvuJuL9GvtGr5lXAi3gHhEK5GeMcD1l8cEezwrBI3/jbkBliKCswgJw+Nj9wh5v7
mI0w4Ad8rLzz/4WquuhdcUwpMeY5hbUYprKS3cBfvIhpX9ocYXeLFzEARd/xafqt
kMOmFECkLhAvpxX/WqjzJNEphuofoVkjzhiwVqcUtQJYngatn96O1N0aUxMXGZl5
puXOyPm0lvVLZaqSbUe9R9Axr5lAub7Rz52hlB5j8Apr+pSRXs+VtVcEqGG99H7C
PNUHSJx5I4oAIsgJVA/KsHIU9o52++B7FaxgpReNfPmObyI+U+r4Ea7nZ858jwZU
kGPj38psCQo9XKrTpD4jLfs+FuGOXpnaNekNfHUwS8X+K/MZDFtFufWFhyKvr33I
+oYrIsYGQGrFBv5krPOxxhB78qxJwHJdMfMbCrRUaJGhxhI05wGk4jIe5A2LsK0w
rxYZE8+DDTc2sftqRmryINJdSwvtJ151TvPqc3gwjsyuVW/srL2XNNwPwoxq4LmN
R+C4AesHkrNPJ0GSH5naC9IEaRHfRhfSk2Mm9ECpMeVRBHwBkfWJfxlfCEuqBllp
qBdHrXFn9AiK31FfUzFhJHAbegFzBEEN1guQKfkT56LvxvMJYCRmzdFIM9S2krjC
6L9S6BpDx/kdme5k+Bx6RIQmdbnx59lB+MCAx7rsISh61rbtA77Y0qJ2+929pAYk
moB665Lai6uUpyKTfcNZSpfmh4CnpV+jGqlAXfbTOG1tO0w6WG/YnIREpLbgLA72
ABueJpAT1AX3aMVacOxrk6SiggRWbTzYVasl5x5XyVtaukEPsfx2D1thdCqiy6Uv
/CAMwXqVbjkna9krHDFK08iX3cTpCWKeOdHu2Bw769DDA+9vkwE8EnSbbSyxcysl
yZTdn3vPyTakGDlWFGC6tSJ3dlEGHrJkxEPH4On7P0ISIIncPvWQ8wg5gE7FJoIP
SKCW0eCZ7ObVMsCVSu1EO2a4FMIjzQjoShrUvrKKi8LrD/yFjuPVahZuRNjPJQ3q
OwpUY4+tREsYg8qCMHN1JLwQNXAQJ0lOpzvu3EeB6QZIp/gcNfCOYJODJe5qb38y
fbz/RHcNWoBUVKyKJSCKAbfn6um4BUMSNZcn+UN/AIMApN0X25WVjGLNRy4lytrj
LGoX30qwVZRnfYv6Xc/jqWHOtPc+xwDwzw0uhJhs0Kj40DRJq9hxGzxwZA6+tsSN
zBIG+wGszgvHAKg2vWrjucU5yEGQYL2SJyPU+CJzXtynhsNgHl51TFQhwMl1a3Wa
ZCGwTttetpSFPt5udsPA/5CPdpjbcqRRC64UCuxMebQfObC03gYqiioTOX2qXsB8
rylHuFryLHHF/SfahS+Z9GZC5VESpd7BWCqF7eRJGi4gn1W1+FF6tZlSXm5bx9Wp
07dPAL+ldAmWRFJAff8EMwoV+Kc1QV9wHy967w8IndFFNbK2av/orDTGjWAHz1DS
MIFYs/UJL+i3Cat11utFe5VxJFW93Mgay8glSh0qk6CFIRzOZHpHm8tU62PdTFiU
X2V/gdVedDdKTlak+sSq9+URbuT1KxZSl60Bk5VZ3IeDFZdBOm5jm/x76sjhcnt3
3JuXocAcs4vmkGCsBISu7w0V1ogFBNYxMUjIUzDdBckDt92wE75E4ObqsKc7D+gU
aQHJ2LTwpoz3OjPhzEYPk20sy8bDnLmSLLnYCTsrjHTBqR6CSvP7+qyhe8ioZgRH
LhFflbRpLvGF+aUgJdTDF/HE+roxD2juijXnu3Z4ySbvGmkLt7FBa3zR/15SZuRU
M3J35Teq0O2lIzh9ceqXLl/S+B7fkMxZ2KM8DJCGJ4m2fLidEdcWagNJdOEq4ZdT
PwSenXsQPvg/kBI0gg1PBCs6lu1Ql7bMku7yMsbG4aX2hzokmHTI5ewEjhLGk/V1
cBlJEnsnj5jQspmJKr6DB7mNc9jpjV54q8oEKR3COni4xGTRai6OCvvcePuekuOB
OT8LlWCwdK5Wj+RxWXciZVgaCgNVz+hFwX3WDzFHX9mXQI1fXgVPVxhwkCLlDJq5
pdMbxTHvEQqvIdrfcuOeBAk+AMrmWistDqDZ93UYw8QWHcXf7r0jbWt9rwtSVQH/
4k12yaEa0OTkCe8S9SfpfOVR/Tm+SHAKtFs5+t4icuazw6lWYzc+4lOHd0oz3qUS
0qoqQu3GaBhh3dfo0yyyl1DamGDSnDIGwWPGbQA198qy8zUg1vHSTh+UI7fTkkHb
vGhYI/CcKAMGR7aL55TmGXhDYSNz2h+a2Ime08mPvTej+gSY+CxzGpzMr3zgtBSA
wjxIDkVwVMDwHg4Tc20rp2Qb2Rki1o0sV4EUZrCBezWOYvomrYFgdl5KBKoLa3FU
Zyt5A/UKsHNHXN824ZwezBa9QTlLHdF+d5uEgSHBd2wcR4nxy11Az7mE/1Ab1Fa6
da0bLqEVH/wSVLnvcRfx+WgB809c2DeFaI/TgVyH3R15nYwGWjmGbjIOcFkERhUs
dUc3TOULOsvlSsPTzVdkJUYWCX/0mqzU25m6g08u/VpYCxJBqaYeavhgOEtkHS8m
qLkk1tZhMLw6pBj9yRBSu/eGGI5CiVSnaCeaQlOaKHTr3N+zh4b+Ab4wBxt2GvAZ
NVBrBjUF60Ipo1E/a9T4e9G5guMdCgQfdHzmpMgXNDRVO3rEqfoUwgSC4ZKpTAI2
Y/auhTS4r+B2Ic4E/DnNwzyl5WVr7aXDBGAFGe9xam8upFFuxnqi1nbpGMeBH2DA
3ZYrZKNTcKk8STX9VRVmkw6D6/NCKufC+tOBXmxbniVov7+bVHE2TDrVr9dx2Mpc
2o3mOFx+NbReEJzJCc522kLbRSOXX/btsu8nviJcrPR3XKl9+87bTQTMOx7hSp5m
yZoeWXK+C7RO7F9Hp5n91lTAV5slAz+qvLYHi9krRBk/vXSWhtek8ajVeDgQTZgT
pIUjlQdgYbGIU0e+27swHa/RVbKWzxvDp8b9A9cjR0/5d0VXPcPYm0QlMeaUPgCK
eNZm5Av6GkBL12syYwl4wdwIA9n1ZuuuM357hpjjfq/RGK3NfTn+A08lJt9M1z3x
k988qwF42Bg07ggi2dhaVCYw65gvYbT317VE1+UChX7pL1eI7v3b/SM6SOzAE/QM
HI9qidu8Cqfmd0VVkNph+Ip9+Utg1myRfybhrYnGLGrUuQmwMt58nv03rxraT5O8
a/IR2wR4Ck50QO+LQF2V/5MbJ+yS8OLxGT0dOuYqk0rFFW2tNWksygbJXdcK5jIn
3pcDudlRM2/re16U8umj/am2OxW4wQjyVL3y9elLKKpd65SaSCzKrT+d8oN//fqH
3n3CIj3bd9M9O968bCr5JGMzfI6UmJ/z63E1sA1A8gWBxOKXdb4ocOfeOfGVWX5O
BnBWyptwzleCDN2z7wnjT+D2HlOpCfMJc370jqRygcETkiER0y4T5xmlrA3JE+Il
kGgo2pyrr5VeEMiKgHygVUCYsNBXeDxWC/vl4I2NWFvzkCF5z3/dMliHbpJlcZzn
J6mDKxoZrUODba+qlw2EjA7nZw/6W3J9kYQwH1NjI8t5ERb3kPjd/7nKOTR5fGHU
5H4T40H7Iky7RmT0YkPDjWV0MEzbohepNLbFShD9CXHfzjByaDGFcAiFJCD/JVCJ
HZ1P3mx7ygjcejk8m/TE4JC6XJziT8r+V7n4wkbufSnI1jroBEZSxmaYdn7/SiQc
WW70x0+BLIV1FNU6Vd4hj/+2DLWmus1aU+wTsvGwHvSda4/a/OR9Y/Ts/1LhLa8A
iZhUjEq9l1xoIvlqtM4Z1dg1tI+Y3NmqMzaq/SCL+llZc0oWU4GGwQ08RYs/paKV
D3FWKg/gP/XMNYrlgooW6g/QfENO6EBXOyA9LhcG05jwGk3VdeOpSEzlI3iPIglW
XKaBgB040hAnFHedrpJMnBiQJYOixSHd0tiYZyVlxfaF4YJsUrhivECxoOOyFk0Y
8GHD8qq3hX7VZzpxNx+NiuVL0xa5AYS/qHEb9f+xbEL9+GZd+O6VDpUVfwim/Omw
FcgEGG4eO+Vzj3FGmxKO1u7wJfTiMg4LnTqoxP5fe0OfFItrLJDEUAMqmTocQKV5
g5Q34xi2m+HSXcatRdxbsUmmdlHhFVV01SPUcSZD9nvcxvdDifuXdElgusWg8xBH
vzjMTS6AoQeq2XPmFpGv/iBHOMf9doWZqBKi08cQBALO2j206qcMcS2BquXRJW+a
hpf2wvox95BsHB2eMWy0kiu7gjClq544BJwq9eEqG5D34NkR365ALBBChVyJ21cj
9XcYvtxYDi01JJ+DrCbg+DI/32sb0NdlFsFMuz0MsOnLXUdoWzqRF1cgZ+5z2M2v
wdOQv5PkdwJcE/ASjbfxotjtwBwllgE+v1Q84TiKdTunCT22j7qmlyGbp2AwgATF
widFHLyjbY9SgukT7phTeqR04m5AgH8oa8X7jAmZltcS4yZX8/ny30lgnjOjpqDr
2nGY5NYDZ/napuO8Hc3P+EYbbxakKikGsQzYoiQpEYp6pxoLgZx6x9TI/hNjdgzr
qeprjtJ9PLBOAhY55LO2FSxaJ965bhagc0wYNgKsUm+u9fwzXJw9nZmbCNa6i+HX
OoEnqJzmwKzkQl198Od0Tn6KyC77QUgxPeeCnm2F+eVciRuDiLv3Fyf8f1Cmnur+
ce9SQE+2zzXW2wEC/zHooFrm84FwKQMWrkHlzDPFNB7653B+PK9qg0COogQ264Um
sroYPOkSHYOndBd2WEbp6rOrSLM80aj3af2ZfydeDU66nGs9zSyrkaekdY7Zv/wS
Y/5o1DZAHQ7755oaM/KSbCMZXS9wBHvbVv1fEJDzqqmm7MjVrJrDce0azmOpHJPk
BDbYtCA1/FkXSSYoVwA5yYFlnMtjSWv7tzd+4KoGOmw6uiruplIZi+xnCZm6xuSZ
ll7RItG27gpYQX6dYdMR+PVIKgIurhftTUGeeHXNAm4bxntBgQPX+4vDBTZBrPFj
sJCT+LpaYYHHLn4PRq7XSU3v6G7nOn0jGComHq5aT81gmUqWQgZwS7cXG7tceLUw
PLGSeAo6kzoPbftsQXWenMmo6qhONlmF+4VLnWdcXtSpnmiGubAr5yIS89Ld/70o
adNIbFuSMQt4S5IE6A0J8pKEM8KNf0UK1C2WeXoxjLVYcpqg49FaTasMiGwyW4n+
mN6LrRSZZ3NJjYZ+Z4RX7y7cmRJe197Ly919qRmNLwY2VoK9/Llln/m6gOuqWGOT
Mgf8Im1Z7gkkKutKZ4gIkIxipSb46Wg8Z0q8SlWkzNLOvfwlZToB/lz94GeDTiLP
wvYdabzSkJmq9P1ob3/ZncUSWV5BA3Z10oS1roYG4dIG+IM+2g7SFUMICYHElZzL
oqhdZdgHSkEciIv49zK+L5HFoTCX2Ye/qz+MGGwh/QiE/L3chPJSfF+dEQflWX2V
bEep7XY8abC1uV6iB0SikEN3FD9wpWMhvDJt8kko14KlYHD9uAPN365fs2OTprvX
n7RbN629jUImPSkhJr+TA/QOKgH3HudfRtsM0ZT8mPQmgx5b5wsZkkLhVVWfRyx7
Lwe1JYVDHdzch4KqKEWOYU2P61sANffw9xOegXWltePQk5nbvHPFOv6jugoU87xt
wehUWkmMdDg1nohBS10pR92Yey6LtlB/nwbkGKKXBAjFE5iPFgSVDGqAFS5BT10d
dAyIhB85P9qPG2MwhRLUd6TbBgGGi/d+C0g6MQJ/kOcSFYYKnBLZIXiZref75fHH
JbKP8FzUPWouLoaDw3jeaSa4D9Xx2CiNHJIiAP1mfIsHlC8QiVcY3HQamvpohTo1
ZE3UVNE/ByBmczye7Q0gw0qF034U2ljxknP+K7MBk+/X3Egz2D6gWiKdJsvznTeA
kXlS8Zi4gt68b9HNKCkO/TeIp6TzQkjkKyhbC8suR1PkwKoFYI69M+vO8CD0TID2
xikmnBfsWR5bvD2HuE9wrZJqKZ/0LxiT1vfo8zC98fTxNe6F27/aEFoAvpcz6lGB
sLxVyED4NGVLWmpJlcqs95Qqq3aHOg42M30oMG2lcdZb+eH6jTU+mzGb6hfMf+6d
OlKJgjN5yOr1zsrCFHnvfqaP7Ac9uYghz6TM45MYhKtCTa31ZIfqlSvUrdblyN5u
Z/0sHCxqE+g2Y/iVRr1bxCvxwa3dt6A+5zmkmhHD3S6YR2R/4hs7zLw0ZntlkABG
4F7QxwrSoKBpXmR9pbKcFoPuXzmJx05L+0TcuT+O51qJM9LCKgv/xwtPg1fIjKvV
`protect END_PROTECTED
