`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZHmYQKNEoaIpzo61CvqK0eVxx/Z1grEbFYxKa9WBOUB3XmX0CVZc797LCgEU9MU
UT5vx13s0oKiOCbiEj+S5TkLCzpe35w3S2gd5duY1vjZj0XgUjhwj+Yt0pC32hZ2
lcl7enqZfm0cpRm61s/NEoZs7secrjkzvQk6pF01yfCuPzz08SzZu2MRQMPaqVSt
O2Qup7JsDz4DICApSWPj+jkA/FpPRQcayu0Kf25553JRheoRxWtYz6CMqAFx7jDW
DWFwbugAs3zDqSmC6WHeDSObQFmjLwz01jR8AAndDgAKlGtihl7kVwqxX1JrszfL
6Lll0YWI1kHf55OBKVToB1cVl8rR/AiMz90Tb4+uh9l5GTP7f674GaEUNQNw14W6
la+fkn6AR/1k6zwS6FUz924MDP0N+0SrlwkYXaq7pF6M0Fv03xYxSlfWb7X6vIkM
7arpyXcTaA2ZCo1NnOTEmtfi1aM5JI55TEP5nJ0bAqXYi7MxPNTGCMpwcCvfBLkT
Z/pDI7Un+1xAJYVS7dOgcuRVDIq+jXA+KWU/KGkUX347NutNM5Pgbf/7lpgh5EzA
iL3Q/Jg+sijLcQRca67nyibAfcgzKKizxTh+xK55CQjFClhG90LAgWaKBFPSw9tw
`protect END_PROTECTED
