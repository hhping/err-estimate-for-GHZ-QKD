`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGWejBMLbiOId/IoNbNEOZYbzFk7+Dn2EvuLcMYyTzn4Uwz5Tiv/Do4E7k/pASZp
05hZOanJ7gkfVgwDJJgFBhzUVcI38qguJajesJ4w8PDeecn6upMch0pI62/mJclJ
F8ihaI/xq8mBVzUy/VlLu3lGcfRSOU/Mi9KpEqk9m34P9MgB8yrX49jvY4y9XI+H
OFDgw1h6+axrlWc1JoPxMkeU3C3csCV9kILnxky4vOM0w3LDHQQkxQlSBFyUCUyj
xJel1nNoNefkOQwLwZKlYK72GJ7AtdvYVrQkdIIM+oOT+4ay0cm1QPwfndO0PzHP
3QpsjgaHD3JsFeCPTySFsmbPYkyY/gS1gVzE38v8kTmeXh8yAQ0juF/Js6Ov5vlw
GET3v1GvJjloZgox7wCdjBmSdjrCwwdhGInphGhvwNYatu55EKnCW921xwNVu/Xu
vYBTWtjbbKREdo9sCf/Wh5sckM41pfdM3hKeVAHwmbdetmHfnPG5DWsBMIfqWYd5
1kq5zCGLt+9QuCQ8RcFo1+3R5q3RePybUhfUNig9MUWpQNJSA3EC2y+3AIy3D4aM
tH43SArdW+L3TH0w0FYpJieo7vHCc68arBET5E8W920KuxTMM7Ao/QeF2y8cjLmq
U7bvTx0MELhbxX5/++5HjolNpEqMJVCdePT+yXgvkF4fIOrtHFD5TlfuyrLdsMSB
O7Jchog0WPN9Sz6d6WmV/+95FRl+UM+teZJBnqPzONzHfiOxcQBzbqoNiBZxr3sr
2ZfVYwz8rnqisn9MUtWOwDxkLFUCHxg9DWC9v+J38Nj9ytrS5roDPUyIQyp7MdfD
oYv6xzuKFdLtaVrSJI/jSA==
`protect END_PROTECTED
