`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjFUknThNCT5XMNNrlQ3BkCZSLiEe8EbytqZSsYpkoCOZHxXVjQeaKt9yfHasefh
Hj6yHdkDPGull/OGDIeQXnZajn0dUCuP1PoorWvyKfsRZU+8UeUT0cnLeK76QC1z
TSGA8QwRQQnaeFS/8p5WGDhU9CQY8O19PFB2NKVUxld4IL3Ksp3ag8vPpkzfDeDK
6cky8p3XA+Hsys1bmnHf+dEAITK2nHjlzFqROJ5ZgsE1E9GxnL+Y4ToAus8KJGnn
CCVXyRm3vEGM6mF3nv4LSOMqBeAkNIK2fQWSD2Ss1YGTBrv+X7LPITvQd8Xml1AF
su8n0FAZcZQZXcWifc9ZTK7nFvEPjy3UOAE1gapWYDr6c9hucB+fYb3VE8c1uP9S
kfb83fleT/ZULhKVwYKktPkhRHmaHVpeiy5hsRxqZqKfm6miOs2ccHVpWztDZdeb
Ockdcn0bTvjrEvY8+aerYd0i6+EhRpq7E2lzT1g8JnHVPTMB4M5puhctzsT4U0Mh
GqeUBzick8Za1Esxl2kj88aEpyDX5lN+l473FQzVS+5z4lCM/fl5YTyVJOa40rj5
IgJoix5iUmFIchZaUv6URO1ak5DFnzqAunPGXjq10qE=
`protect END_PROTECTED
