`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aP5Kxi5ojoTB1ylt4vtHv9b7xIy7w+3QE/Gkwc/ALSSYUSqwURHg3zY6YAZf3FaA
4EVyzcPUpkwVxWhgCISUmAqv9avX+qjWWlzCwtChdSKwz0y9SiBSNpypBM5Rw5df
xstNb8P6micYkvgeDY93F9XtlVst3Ahvy+bTZ30W85Bmilym81wzztVs4upKPVAq
RE1kpoAJnGt2/wPYIQpRZ+lbgR3BQSN23l+mLaWHjGU0H+wQ7RCUXSniOYi3pN/t
fAXy28MYLaS+ES/6xG3QSIAzRVk160m10q/XOPj8H0PuwTndXJNGU4vOL+4hTLbk
Qy/d4zW/eZfp41jz5yaCpqTEd8S2r0/m0MDyoJ3GCFgPbxVj9UMwDy5xpbg+8OGw
yFjz+yghboICRtfq516zqfQ+7Q1G4Mv8TH/tjX9ldQnR34VXzmp5ld065yPRgKOK
hMRXrbbbt+gPMcPO3LAMjCTDceyJcLxX0GJ1azGjTdR8HFM8+Wxl3JM1mV83InSX
+5t4j42BRSLroJkXhdObPIQGT/SRhklD/BAw/YIc+4UZPjxOinLnaBWHTFiosZU+
evSF2rZL/hiV/hIKtzISL1N4jTHk2LmqOTvh1Y8bcKYK5PPE9R9Tqx7zqcOul4Zu
4RUw2idTEYTbqx5dKMFWkA==
`protect END_PROTECTED
