`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iv8b9CCu6JCBb3+ofgJjLYIELLNep5fZG4oTYvxs2YO4h2REHUOlnWoNSgdECacI
sOawd3/DFaPSEUiGirvbXSnwXQeDsjkbMi2fFVNKIzd6NpDSQASdYs9LuNTFvPbP
iqVOpLxIp6mXWlFpDQeSqUYEEAjxbhaX0q3O+mk2GieTW/MLHVmdJtnJjFjGglw1
TQhsuqNd0OfwbwzdsiE2Kt3xcFAc1CC8q8YNIn3qJEc4HyicpdnT126RzH2NjLrC
qvd66f5vdyJDeGB/wuTzRrimiTjy4Xcc4Ex9X6zK98znN8ay8/7HiKaFVCmay3Zz
7sUv52CUJSWIMYGY9WEwhMW44dpUNRDFd5xjlJlTp3CPF6UeT4fuxOX5+IcoM0JY
oLe4juhOeLaSEW2kWE6QsDPjbEf9eLjoha6H2BDETTQOB49iamsKSIagvJiwuifN
fPsM3Ag8TFasHUcCp1sNXl9HXJw+IsJfBT58zuu7HVpgxEzNhfBRwjk+5ek+pp2o
xuW8LKfPZp6ybWPdhVZ11qzjhw/4amGg8kHJWmuNwOj8Ll5e2Kvx7ME8SmskcnJm
91Qvghpano+rzYJ0S2/+gzrdyqtjsQKk0SRGCNFAXU+RvD7pI/HUeugq33RHUjnF
SWlSzqU3/4cqFQeegqbIYczg7ef3D//VJtcErrUMnApkFA5JrYPFMaNDhqjozyb/
D0C94CCA2IPuW2QHY/yRR9tUBFVhCs4Kgcd74+OhyAwbBM5KcMJnXtuEx2HlkAgf
KzfUMxV3J1+EkWXLaZxEdA8pvWFNiU9vYwEGAqE8tm+ZUWcio/OFOZQ7Adx77pYW
bSvPaOkYQ25gw4n5onjmNaPYIxb0X7FcEp4x/3yQvuqtTKjsUeyYtnRc5iiWVCVw
fE7y7jhXNUo/oNIhpQZeQ6/bB01INAx6JXyhN2VjI4TMcigyISXq3SJVDtavkpn9
+1b68cBTYQx1JebWScxqNcje+MBQW1UltOPftZEPrVD29gwN7qEP87E51aB2s5kA
lV5HL6Uu+w6yyrKi05pZeEWDmUfinSMvxvbfA22ro9+I/VwQNimCE37BYQjvU+mO
Zaj9Nx6nVBXXvskXqC1uHrhgF6GVJxq3mrVGREBj/DWZl2BJzvCy11tHRjy76hKT
C8ahnkHhbkO+4kK1I9V8oEW46xhp9Mb2G0guSer5E6HsSQI5gHRsIn5kIMWJgk36
3KDYuZVdjoi1R/k/EdjKniLA1+wMQBNxCPzyJid4EM3llqT0iHZwXeMZLUXbWEag
0N6jJcjSBqGjJkhk7/W6PUGXKiEgbHrwhDhN0Ai1tUdbkPvl8pqv7TlDKVtTYiYd
7OuC1U2vxG6N4V1hO2zRKOx7WxBljqjhaSdwBe9YHRWaJK9QLqP1TQJA9O15SkK5
V6L/M8j7254sN1o1qTJwU4HIA+YVYcVJ/a4wBr2pS6lWFl1pQPVdlz3LP7h+5hkk
8qc6XnKEHPQ7QAiOWrhwWw==
`protect END_PROTECTED
