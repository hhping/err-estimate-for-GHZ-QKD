`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USmiNobw43l1ohu72yd2ywhvwF/VeTmxUviywRSumVeND+BkEV2LjR0WbeGTm+6H
yOG/pAlTylpgMKFRF9GT1qvZZYabA39CF7nkEUk80ANFJPxw/TAJ/MZtcYsFUvLJ
HIyULY9zG4lHidF0UWst14FZmeQTfpvfWxVmxhM2eiHiRF0XVAF6vLnn9mF22upX
aUO33VXnKUYbavpJYDtyKAx6Tw5HoKq12deSMbKAuzwAmZCzOytEuC0LBr72y55F
DCV4WUJBYCJ3lQ27cJA7ed+fcfIabjGE+NWU8rHKjUsbrsU8XKLJlEp6KgpxVQ9M
5Ot3rM+PbWPXEV8bmegin73vDbHJp0950cECJm7ySt3CRGxeP1z6HgiMEhIn2fjm
rCLL2zgCwg19D7kUaZPkFExjK6T0G/ItZisZBetxKuw6qsVgjXXZmE8AtaWZJ9Y5
EFwRIE9sigo7vtcFf9/r1ar7japLFMMGS9RwCiRysPsseayufMpAW2bpjhYtr1eC
NjgOI4/Dhb/2Dv6jpGppjmLtr6eYoXEbF4ufx9DTI8l1JBBLLSMUZfgxn2B+Df0i
`protect END_PROTECTED
