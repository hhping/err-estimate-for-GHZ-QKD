`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctQK/9+ZWFIKyfR79w2JTg5dogxl+BVT2c7OsCpN6MJwM9qkL1vQEoBAgpH/wMO3
PKVbFKKe6b6dOxC/i/To1dVtGQ/Xsge3y+xxiEuTgbUUQo3TrYtRp8ekHiefjDJL
M8D8WKshDmtP2rbCWh7kHBxz5GbJcXRwuLr1FAvxn6CtzjLRWAIlml0yngVrKfhD
K3YAPtQczXI7v5691l67RSNwk/QZoUL8EdjDHqaANjiYPwnP1zYrOjVGxIRSe9AK
GhcD5DEuH6G96dc/yn3EmlMt7jAVP3VdQ3QxJfZm3LyToZDYO2f5OKwOWHtcBwUn
cFsW86SC5oqc0MiFtbGUdN4EMApP/0BWSWit5b0J4ykVXcUqMe5QAHrhQl414ZFx
CzzvAC9NxdJidTnmOrdtpvOKd3l1ayfQTS4G9xzh4aoC7EXHExjfnTzFNbS3z64F
wQZhQZw6twnvJUPTe9nv9lFp3vUBXfgIoX03ZgLDLz0R6+KbI8K/SK+NTUqgtmx7
iK9fH3WGqBaqCo5OE4mZdXLjHcdUfzR9FjCD9dYzPZm/QyJzYUHJf9V3bxm7OC8W
dnlY33sWWK5JZrsuHzFMBWo3PKYQcmzAMJoJJDUeZiMvCdzQYwwfRBX1oY0/rLll
vpt3YRA6HSSgia5/OsXojIWis3lpBvA2OVJp0H32wPWGEmoCmREF4qVLSE8wFyPk
xbJLwzx0IJ545wh87dj4BzE3Me5G2OP/VzlHHVt8rfb5R1TVnCggaDT+mbW/IHbr
sNnbAGdxQp75IYa52mFX+w==
`protect END_PROTECTED
