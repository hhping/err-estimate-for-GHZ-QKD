`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8F02BB0nHIZFB3bH0S8hmPtPWpAc0YxTsEcuC/Q42AYVvl4uhF6M3X1e/npaYeM
D7A9LquB5SdPKBPwLBCoSnBHs2KyyHOxCWoBHDuKgipSRRHsgXXZ9y6MLoqTn4zH
lQp3ln5AXbFEz+uHITRt30+ttNCxQ5JLg/jVRqTGD2BssXvMV3lQvDwfPlwGV3uc
hMfZznK7dB9VMF/+/oc13OEDrIE9ES1s0DU6fjswqxF3osn+d8iHbhsdFbjUP7wI
WXH/D3aU2H8iOg6v17aIITh7SszRxX9k0i0Aw++LDacVTs5ONlbSIsxbdH6+ySY/
z6CcBcd+FEdGmT1XhEa0EfwT6luMBXBEi2oIHBdVGTx0Q8n/yacCThWeKWCQ/i0Q
clOH0LzQLkdr5dvo1/k+4S25UAESdmHVXHyZLQBbbfTA0eCaCzlv9bRfvoVOOyxZ
Nn4AfsQDWzAIsNCbwZj3G1oYW5cVxRdx8+F0N5wdkyMlh/zZwm8yHMVsEFue523L
AiBdNQ5ax1m66OvxCYDiTOUb7HEUUlxg0+zUTsdGuvsqkVXhwz6Lj0OQADX4ff0P
YxNHDi1+cIdVC4VtegAxBajGyJVK/coVBZPs9vJ29iLid6I1TiHFJzOO/LJTHJyb
WH4DEAlrw1Shcz+/JutlM99miZw6gyZFptxH7cBCdN+/RR6qGjuPNQradedx9f7P
eKwkXLqGBtFkIK4DFWswYYBebZl/nLzZ5Wdy7KklrQ0=
`protect END_PROTECTED
