`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
orwWjmKKCWiKiiBAmOBvJWxgLWwNiRVzMpXn+rK7JKb2ncVuOsWK5pSAkRftOIPY
14uzMdnw0ZLqOd3i4zpUBucB1fTGGJcjdJ9HN+Ubjyg9cP49NYTJNDe4mIJMnp8Z
HQEOn52CvffiFAsWADWVKgQGmyuI0S9uUm7fs025CYPMLlwq83DObmO9MHhx5SHn
WbFmY8k+dbCFgoAZIs2+J7eIGHiClZQvo0PKzd74nbsQlvPSOBb7IUbQCF6mSI6m
1g98KlPwq6FhdsbFUHMA+QFaH4Ft9y2Hamt6uh60Astw8gLmADgKOcVBeHNAHrmg
fIs2aKAMcszXIN7YzZ+JpDcJyZxu9wHM9GIzg0o4/rZ8/7KE8ba9S1wFj+pSrUO5
AeE8NDmfiw/gI38nYCW2pNFE2YLpZGwJdgLcbm4XNxsXzGHvYI374e+B89R4ygxR
pMna1HO7L+qy4gIhJwNHiBsp5NTOPGggBLh0fRi6MnO+ZNhbhw7AIg/IeHHausQo
FmeKl9T1xc5UJXMjNaJYTRBtMMt7niymDMqCxCHLmjOGlKZ81DQj+9UKRJczD8eX
otMHBo21CC1Nq7uGOoW4omHX3Zm9qLUakqBZ4mrYBdIPyDETpBOG1fEoYaEyFgi8
`protect END_PROTECTED
