`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRHu48WYHiVeh4PMFTBLew16snGwC5j47guVdfPLpuKmsbvxNWtNieU+TQf12+ky
fK+WzGMKpiOn4j0AAilv0kP8Ua5zv95uaG4MFfDZlBMLbGcFG5T4uKFbyT2ZIWwC
RJ6Wt+8EHxk5lxjIMTpq9Ba0jyToQ3+N0hhoSGg5e3nNv4KP2K7Ux2NhntCCwKwR
pMLAB9MfrojzWin7TrdN2by2D07b3us30GKTGgO5cIMZ8ix7zirXIIl+7PwKbwrY
7yDG34XkbJfgvECp0th/D8F8JGmxwq2ViLH+Gmy3SJ4tsaUusw48UVHgrVoV9ZhG
FofTNa+BZy/qDJuhJZfRn0qQD9DrjXo/AYfYIWY27TVewejTpagDfQ62gBAqgba/
MWvynbUrb29/ceMypxXg7CHdUVW22qNso0dn+6TUhvxdB0BecY+bvhh29YbrDNAP
tJ3NyS/WxjDGIf+l40kcL9LJCHCkURlB6EZI4+3b5QBxWF67V6YcYMvKSK3W/2Kx
cHdDbl6WfblN1K9c47ptMl2hklHQCxhH0ijWr3Uq8xPEp5y9/OzvN2LO4+NAXI6l
gVb67hxK+gkN8nSJEnQfSfe2VEkM//i/cvK20ol0aBmtKWW+1EZkevWQk0ZPbLx1
LZOWk84pHOWTcjxqBp8cCr9Al9d1IhOkExVkN/Yro4/956xtZfYwn/8J9W00hRkC
PfSoIii9w192SW8r4oDgPuLko7bDoFBRqAdcUMMWSfKHChpZZm1xnFSSgBiOZFev
4ZnTGvX1HuNlNxvcUjkjPuxhdn8vbklbUDoTDIWcMalVnOA6OoYCZJ9HMl9LonvB
e/Lr6MJC6OE7evlGUgnYddCpU3h6Zo5dzNNat4R3sGnFWylJX/hPyvbQ3YUC65Hf
2A9wBpDjibUWgIuKBAlBmUBzSaoUHALsDQporfEqWd62MIxWVfS4wfDXS6+FLru9
2jck2IkjFQf5uNYqewXyhocdcP9rI6IiSQYzgg49rRE9Ga0rKMltdmv/6M3H0cJX
clbV2M0bh40BP9yFNT8yeHUPmUY/D/l+Yg3vvvqqj6/MnkFSdRzn5dqzeiKpmfnC
Y4NVOlkkdCiouwmE74T+aM2rTjI0laSzWXEiQQ6JNuiYUvJGLbstv1bzGk69wy74
qWtCRPcQwX3oWsC2Zie3524g7atCpztXMPt9yKdyq/VlMLmzz+uM0Q4rn+d0oViv
bxZ3yKNzTzbAgykRrGPQgnKY0yZSUWJ9wTz/pIMils2jFWEVqHK0RJhA1vjNOiHU
CLPztC1ivTRxZPFhqeKekg==
`protect END_PROTECTED
