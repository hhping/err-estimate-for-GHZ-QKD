`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tB2XSw3QOtet9qp5bZC8rtxpgSjoxUnEJuzsJX2aQyWKV3b5Ij3FNl5ppHeM5qXj
0O/EJxuEGxhoVPe3Dz14NCfrBL8O9hIAg5evD1H8lcFAfC0CQPI6H7+PqeF6B3gn
mnX7UkCW2l+hKsPqQ2ZrRw0W8n3iVtevUCQHWUnoi8MxTSky2V1Qu8j9kxOHOMeq
m4NDK9I72TQbYDy7VT8ffr5ZTyYCXyny6ZaMlWCu0Unrnggi6Pgok/2++xZHGRyo
UDDWy3B+l6iNtEEO6HjVmss6XcWjMeEup7IJ7qKpqvrWo1ltoQmjwos3xSBhiG5Z
VGpi7O7etiL96ISVuRIditWjna1NgraBAo5PubFJC3vDDxpatkd97rcAPjD8uGFp
llNT8KjRAjLoQ04ll2wMGd/COV4ueYqipA2YAAT5FJzMjr3dg3ZqORGENlOnSBRa
CmAT/u5Vpq4LZRUnrl1MhTDG2BDIHBRU1G83PRYGPcZueXNx03ulgHE/ngfJQzL4
B4L8+2bpmaZUSh7ArUnggqQbGbsOoeLVVyLGLKf+em8D5nExU8gOG1mo/htfdZfv
Z6cdm4jnhEA5/738T/sCHvuWQYNRnj7sQTy7ZWAD/13IcOBdIn1kdY2uoRp3CdM7
qj14haiyOyRwEHb/60guwDqiOGcGlJRJ3ADNihfw/i/DwB8WOfVp7qGrp6vxnYvx
rbBBIrqHKz9a4Q/6uQDKL9bfT/qssNEv1mzgxFxuZfNrWl+orRlZm6wi1fmTkZjo
Cm0RftWmHhCBskw4qpsd3KnSh5NFdnSz9V1335S7OrpyOf7gD06xBcWX+QyoUKRf
aGzaQoAyE1+Ftgm2CqhHx6UvsyaLdnpDuM77p0fUBhs=
`protect END_PROTECTED
