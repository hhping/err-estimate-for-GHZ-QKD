`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K08XuxPxcsnsnSAXv8LXdm+6N5UI1bsz1jtMcCrwz1Ydkkb5w+LqrRa/Ob5UlINz
Hli46TFnxJ7ISSqn0QSWluplvMJjnLTL9ioqmDyKr9D1XWJVOdkwLR5dcw3GV8R9
EgrUs5ClHo2QHYzD6b2v516ZTY7XNZXzspU/K0diM9EW2d7yNAFB0tIHR9C2da7a
E5KJLlA9p1hbpFxIx5WRD55EJgRDHNK9RUZruc8VFIjaKt4P8NVxpJmmo1b2Vkjz
8eWCZrOc8WAXCdqNwtfQKGl3yp/w7fsME4gI0ZCXNpsWlP2CFH95ouhn0Iyens0r
UzV+GqlsYXb1Em2c+1z7tXMp0nzP8HlnkJamqGFzst2TEbi6fExiO3BdyQHTMC1C
CrEg9w8gaBGkKeQgzLDmO6NRriK9SRxROh5eszlxa6H+EHfQLr4lMdvXTEE/tAIz
m7khUZZ4k9YumHi5h3aHYw6tL+6eVvnvyFzQNGvQOL+QlSjN4qCibcSJtSvm/fT2
wY9lcakon8B0havG5s5LVj8y+RdCTyO9DZcTc/SeacbT+yNqMT/AhiAZZVWaisZY
7sZb9RjzEJBTet5rLgDcGbZU/QfqLiCUkm5w8FuRmZr2P98QVEcfNeXfSPfqNwyw
YUgReu0YyJGeDVPMeTmFo+7I0kHx2Pt6TlkcciRNRC2TkIzciVfC+tItgpnoPyRc
r7J2SnNtlKncaNzzKD8JotS8Pkbs+BQBi/8MUFbospC1mgWaD6pMXUB3vTKy5eNk
XbXkbGQ7LO8UdnamroV7GsWfN0AiyFAXbdS5ik5/tpF/pKm50S9iEjD/kSw2BMc4
QbE8V9rrdIaA5EFqX9Op+rPTyxJgqSkDTOrVJBmA/kIn9n8WeTkCPhV7bVL1u81z
z6YBA6IKVPAcyzT5YuwKkNFntQ6oL8EF87xkaxZCNH7nK7nyRmIRiNWNiWBYlaqG
151xCrObKPR1hdRPztNVrair0OjDKglmkXJEYbkc5v5rlbZARx3nfBkFdnHBTVba
Bq1S7+Vp9rfiBfm+sSmDx6ZtBL1l8jfTE9fGOy4VPwTk9qQ41ww8hnz3NkPtCBjO
F28OF2bYweErulMAB3kMLRfnUmdOgtdli3hr5iI18KnDsC0+FI7udSr3+8EO82aI
3BdJXEdlVQgF0zi1ofPtNPnDLg5xhVpiVYCXjGIGDWmOm0v7iSy00kvd6UJwoXO3
ePHleJgUNAbxzMh7kunNUUGtyZQWVZgbu7auz66OH+6c6o9Q+3ipn545cUzYGvdo
NrYwM1d7r0qmf76SpaO/iBNgxGRS5rPfkNXCaIXMQYz9/4AG6Vupab0Z6kYSEZ5S
9hTtK09uDXtrR5kGeIy+78sBr7Us+MtISBuETcLy7QZOrI7nTeHbOsCZIWhj9I/P
3bC6k7KvNjD1uOUnToceaH6oc/kumrV/JN3icULlJOIdh4yUKpVJCCKZT60+tSPP
pIbaMWH+K/OBKLLv15EwlRdLCvz8nwRUh4pLUr0WC5x7beywDmdBjKrp/TOqjMCq
JXFKuPOR1X/l0eM47qLi07GoeWuGfuqIiJk0tLKrKq/2Aly/wr4AAfB4cSUdhQTZ
dQkY6t2JYUuHW2cAticF45eHW/cDSHrg3WbZwxNfd2a7yfxf6EHvdG9bWhPm4Dn8
9J5zyHlYBBPPIQ+P1sgPKGomvh+TXdxPHV1x35tTSt9G6RONXWN77f6foq5RGqco
19GUFU67o/nbcyCUm9ny6km5lTgns8aZjY9I7sCYjtQSmaK3eF9edeoRjPadN4ZH
VkdfFGu2FhohT4GwcAGAaoQM9mdh4Gkc4MQPTMWeJYMYvr3Hx3mdKZIFTHZq46He
/ifeHg+FLT4LmMk4ubkHe/e94fe+U+HBVyM/N7umiEks5hRC3woMxEG9xDtClW8h
t5RWlrg6vfOmF1m536/+fg18ezv55QnTJh0fEaodcKPoim3A9DKaqjly9XLmwmSd
/NYR7ICaLgQyPd3zWowkUA9IC1HelvvcdB7X1I8C7rVwQXUbSxz7OQHoDec0Fz/J
ziK+KBkm2hH4V17EFs0H/oY+Vo2DtWNjHLHCz0RsFQ7/0xJUGuQZin6NOpDrJ/6F
kY7BWtbM5Xxqh/oIMbzEXUafcMDJJ7N28Znn6FGJVYHY+i3ZyXEMQz014OA1aSAy
vjHRzFX3uOGTOYUy2lMFqWqrrFA57aD+FgU/n/q4RIYsYmkGHsoEr5jhCWjm8v3e
nJVeaUr5oIum2xS0y5TvJf6J1buRDYffKm1eqI3WWGGppisIZIs/WEBJkwMb8QlJ
X7TfY68776m8AvfFqiTga9TfjDQ4R674kDr+A9bQnTAKQeTUDQhxr+3ilp6hID/h
uMQzZdetMO4AUnpWcJP7NoBlb0ZLlT0HpJA8gMmzZQH/TX1Vmn/Kef5Vqu6ageQB
9SIrYO38q2kWCrf9s4BftYxcwe9Nfu6DitEquOkdfuZLM6ujipPw1Rg22WwkoiFo
pc6kvyCcZ3IMyLtm3TNjB2zcstBsferB3vfhBniqlFWYCaN2YY7wvjEbb/HP7mgo
r9bVFncTIyfgh9oDO4LbvYuH95e+KBQtMm3CeWIz1l1lal4lL54f56FhNUm69dcZ
/j0mjf0QdcxsdkJwZ3Yls+XJ7e9DKDkXyNppLsNkWK7RhHVuVGzA2jfBBAA9gRRx
6+ZryG+U0Wp9jvOlO1+OPg6gw5jAPyF75jFNICz1EEG2hG3mO98hk/7KcUQ+wwvb
4lIY/aqX+hGFdzNaWJDAGwJ0SIIgz+iUkuRnIyofrYzkktOOx8tphiKZ2mDG7kKv
Eec+UcAyB8w6TjhcDNyoF+ZXZtQL8z+FI9mCS48fwUZJcyk0CSzuSeoFaCbEU+Ah
Q0Sb/lEDAqjHUP+341pQzbo/uJ6KjA43Z/DYMpz+iSzqXE7ppL+ZfZPvEIsp64jk
LztTPsB8WGkNN4RS3ng8mnMm3oSDFIekW7ujwVOtGP7sVE32NUj7UTUiHn6CCitt
eF6VkqbYzu/A75sWhRN+5UopuF4cK20cKkZJY8+Z1CdZUz0cAFiVKtyeOJXA/ZHz
5jlELsAnMwtklxb4PDR4M3I6608mc6aD3+sp7YK2aiVFvjwhaKOIP/aitlJsNedD
TEJlTadgo1m5htmNd5ZfEg+gYKpA16UxG0PfIw2TaQFzdbkiSiMwqXz/XHUnUyqU
HjO7MLGvJgsT4I05Gc90hm3nwwmgT1Ljr5eqzxuD/iY=
`protect END_PROTECTED
