`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
snmRPvedG5PZIADotfDEOhtyffgd/xWFzw7jfN0cHYETYIg6vrPAT5zjjsCpfDwZ
brSFVgJM00O/GUBiO/MHzVQmUn2Emt3jazTW9q1IU+hKWYqPrC53UUltAhcGIZnY
C8QwLUcceNkEs1ucXLN1hfBG/emqR6thVRiAjgDLo4M89wj3eBy3kF/bLL2rfkZK
wLNuOSq4EIHo3S+rUhwEOW1GMTGTjm7oBVfkpPIFnHBzHZNfHLqK1fcuKU7uAsPu
PYpLgupD9LdoIBel+fCa30LPM9eeDkQJOboTTR01WDAfSfYr5AsOf0OWM6A7dImU
yJ59XIn9UNn2EjwZUiEgv27YzveKNN+cxOUNKIXCqadm3HgWQDo83Gk+GiQjGmqD
JfiRHVCbdsRwvNkFuaV7LGsTpc0+IeXYrKiKfrDwcEPnC8dONMWu/q3dQXhr/ow8
vq5fHGocy4VDkMH1OZ/H97/vB5sznz+k5v6DMPvIpfPVtZpJWINUyuT37N5HyIwz
1RiZvXI8WADOxQJ+UwJn5+AlvPN6CfFwBAXE7jejUgAIPyLjSyxQrXR+LhKKRjzv
+HPGS6TWYeX8KK83YtENLJbIa2j0dZtvBgUyxwhp/cYloLGh2C4WaSTLtqQZSn1A
cXQ/+5Oq5OUrHXrdRR6BJQUUlJBbGQFkNhgDVoPIEzdeF7enTwa8geAxVWYQqh3g
jj+EjdpxqBTOJGm3rGaQMdroVOADbfBWotp8SAqYkmhtnjhN/rsbw/kDc1YqXZkj
8Mo7EEbJ4w5uUcTY7+yQKtbmkENj4q3VtosA9fwETto=
`protect END_PROTECTED
