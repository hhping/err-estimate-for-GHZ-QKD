`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GsU0ehU+bDHUC708IBmbKJC7NneX7G6yZCsGwNlMSranDJr6qpq3arC1O72QdHCW
ghq+IehoHby3R83uSV23AOOdeIENFeeODK5OR+FxEwnw69ezhozi7J3EJzTVwb4E
LAgBt7gxiWoGFvCPIRUSTPkpwt6yzqq2ee8X+K4Vh1uaLm9t1h/pXsMn1RphGZJF
JGROw4uYqa3rfCkMwSLaEH0k91MDewYL9ZqNoA/0OJi9u3Y6Ge4mF5c0MSV20VFO
RSVkCi328FnFVvZH7QG+79jR9BaY8aJ1EugunH3HUHiW5oN5UfH7PdMl1QzA/rVh
QQdCStGw8T3DfN5zYgcQCuXfPSud1ZjSTnZRAtc9optN5nHzmkJ6C4V7eZyIlqRS
8Ho69l/8LPgxIq/I3EZ3m7RdfPZDEk2KVLLPKo+5GzR9jB60xeJagVAK9pARK4pV
vA+2efN/iVOklH8/2XtsboINCrb5oh52leBR2nPgJQBy6SSVgKTKqsJ0MhijSwCu
8l/CnHmQjlF76ci4fwFPbBG5VpGCxjPScigHFg28x89RhmCtYvJcRmTCTRZL5br6
vbmFOpEMRwa6+0N5C9+AQg5KqiWZ4Tt5bQgtyGNTo3RCnijNsvkZ2FvxQ92NN4fS
eBkBTO2JENE/oXl1w7OgYHJlhSfJSSojCTrpLZIeWLravROeAZLMpjzuA34WrOWK
8hp25ZqcfaAVpoVWCNbT5jqh1R91dYl6TS5f0sqBHMuQK/+ZExebnRi6ozSciP/O
R+KdnhlEj0Bt8h1/mAuac4Ya+bz44ZllQj3iKrINjB0cq+rxHhewMjPY1pMVKKv3
lyk/8z0Ktf99AfBc/JYL5pJ5uGO1jACg884cUev7EMfo/qcnoCgVB4e3/01VUUz1
K/WeXRuS3SqUYTns4kBCDe94F9a2SFM9shXxzJUIX3aVMjGe6U/yJw5vNBRKgcrf
fmLkqGYoNu5ldGxX/phwbjqq3IGxFghba4ICWcwU5DU2qQI5RN/w+RfuVctw6zUP
o9WLbStNyHJJCgO9J8T1DfoWOse+HtQZQGdLbtDFTHoPGetHb9JML7DuSjG1ZNJs
jB1MFFiVFv8if2mNmTUs5pSTwG3VhJNXDcuzDLIrgFaULQ1cyiPBgFbZXZKcXe6k
BGgFeiSKJwRDRRA5rq5N2sgDQoNvBxzcxtzWVldb2/MtC3kZ2sYoXlyg9SH2wfIc
1ssyAbiwDCR3U20vCtC5dfnzTTmh1qe/K+C9g2bkxbAhvtHuMaKtupEj1lTNyqsC
atACTO+NiEe7L+MFucq9XJQOHhllMTbgwhZYUVdiMR8=
`protect END_PROTECTED
