`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
344iEcx1yx3kFpH0kmWs2CAMKS/k2ltGl+MGx2FoNvfFiCSpqND6GKSjOtp8sUO6
vt8Z8OjUMqDkChPNEDjr9gMsU0ZlCWN8WlvaO3TwIDO1GpJ/kjTqsxTYSnIZg8Zs
PPAhhKW+p9xxBdJwCkntXdzDTcl3GZR8XEW3p3FOcjK3cPi8PlgXlQ4ag3UAYwZC
pbBkkLeWJh/VyKavUdXvtdqq9iOqQXSTwwKZeiHt2ctgweG3tP4uAxiedZLceDGF
/AqyY3EENPYFThpCnB8VRPWQV6QyC9sb1nFwjw/0ZGw7p1TXIxNlznYn+n7RsISv
vm+PgY/ubyE4bIutSvGn+W6nUWN4KzrNM4BzpuO4/Ph4Cd5G+gzIKZ9bnFuuiVf8
/V0BM0yU8VYbXfsArqiW5BRaswG1GOEsml1GNrViLDhRZ4ioVKBji6itfZ3gIgy4
H4BSoER5+9CL55tIdqM8g84nCmEc+FC0zwAmjb33UknC8wqGYYpHgnTGkBE6U+pN
9ll4gQsPqTl8kjqgUpiWb/CTTNpgc83UXJ37CYB46dNrZ6ii5wbUDOtYundYAFSD
oQzxnuqasz8m6ztjmCmyZfDF0Q7b2tKm0UUVqClvqq3C/AqS5iCnq0dSo2xapSms
kXwaqnG6M2uZSdTUk6DS6p4F8vNFFLpb55k/KjNJ7FDGiRJCT5TmGQObxZ2nJPIr
Z5dOaWm/fSrsD+zTbHHvtpnLeyO7p6Y1CYOo3d9FZHzUHT3cPpzqs7Gmtjgdn0Vp
8hha4aVgJ6HG9jnhfZljj9WeWX84SGhKRg7yDvJheG144NgE8sst00aKNxKcpiza
zOyZpI4ESvkmtIMyPnJr5AnvQd3Dqukk3wu1dHYY1Kv0K9uhOTJMrQExfBDDLWWo
ruLU4dA8ZW3va7YSrGHoV+4zMujkWsZnns2VDKBNe/PPjnsnkNG4cAyVniBsctjY
gL61qBILosb5LnVUUZQZ7K6ZTZDdmZ1KnT/qotFwWyK9U1gNDCu2Pcwxbdse67cv
7UFJqMfPQtGwzSvPuDRfJUuoQ76XGrnkjmL+K5HZ7xroUkIInqxH4RZc74ESTdRl
2p0PMUIadtwe89ar91zFVmvoQCHa8esmnEzNauha71Scv08EO+rN77BmhNHvRUIy
LubxbYOIDp66lIQpJ/yC1EWWb6ZDeReAf9+Zklt85lLlbl8XMaTSxhRxELXWgN+S
VmPepK1YRaiOrhiX8mNKKKejgmpBYOKQSJaARHt++d83ISRtJGs+rEbqOqJBWV40
77pBFN2acXbIMRfBE/YaDSkRJdUz977Ml4iSgfGGjlqxwjO/WAIaWPYPX4CtGd/l
w0bacSnUElEJoyQuylLN/z80sPSLMtktclkb0beSKgX0831ziWtI8LrFAUfA2tCX
nQJwFFhDB2HQJL+UlPXCMIfVHCf5n9CDfR8qAQhkvXcyzvyjKP5+m/1c7TsV1P2L
74/ZSXZzWMs3igOH7d0x5Itdid9ptJmikSOVjpmbgsrsAVNuD4OyfIZNKEoVdfqe
3IrUmEpRQmMFfEArbLRb35ebHO2eoZXuVzxKllQR4zzg/F0FTE9nWuiVrkFJYCY/
KINEWgv0qxEetMq0xT9dnqn9kuVIFmYSHX7dWvy5nJjXIyTOXb6MNIOmA/37P685
RoKxS5ttEAyey4oNYzeAQmFvkV/Wu3Hf1r5sNu67erARtZvUA3l73a21Lb+KGkm3
uSrXJLF2UkFq3Ff5VJNcL0qx9EoaPdOsq5VTzBdGZoF1e0ShSCEQOi+Wy6N958te
43zHkamIboXzAF+8s5aUqaC3g1FqnjpYZ3P+tCdF0bObfR0I8Xg3SiDN1u1kUbku
NNDryPt2R+UA4jm0vgM7GlVsmVTL38VYnyyXIvfppFBEJbNqdYNQqw0x1TeY+O8X
4w37+Hrgu4rhjStBm+WIf9q1h73OxkDbQvizZKBkuQZOgaT5kP9b4HIh6QtMifcw
2waapWJGvkTZBh2p9JlhwZUAjPzQKHQAiHBsn2xeqBzhRkfu+0gSclsQpURGHXH7
BItuAPf+cYii4g5mWXPwhvGGIVnRFwz5YqslbxshpjcukVxzam6WV1zRix58lsRJ
9jVqhVecA351DpfRRSys2BDh5U3l41D4p+j58uCKmoIYUutDgON+i01C4KtDu+Jy
X9LbrDG7RzDc7V0ww+hLBFuZTpeOaP2FSAjwsQcy8G9zNUjxqpU7XoRzY45vNU/0
yZquB/m4xg8swTfeZt054/qI/ndD4RGNyFhYEvXTA/U=
`protect END_PROTECTED
