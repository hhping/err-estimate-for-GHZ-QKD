`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+8lYDMWyjDZbXRetim+zJfIeNjMoyuCHRiNbOZ9bfUjIGovhBM1nZs6U1bwtjyO
Fea3a/ieDRz3X9BvpEtOfnkafl+3GFFSj7K0InXIPotn6zs5WDjNnht7KtVXW8FY
NBO3Bs3y4E5gjLKs3Sg8uaZa1ubfgWDfvWpL/cllGRBYNSLTHvvbppA3b4ECqCGB
Pwh9I1N0bLrb6hkVdwfjLNOHnqiEEaEmXwehd3Ybl4dTlZQcVLOFT+7fzeBVsC7l
2iJlrBmeeuM8PUzPhChwCfbtd2Dq2Xt8yjqrkPXK9K7YS6G1oX5UHf5+UpE1DaiF
bOTrHauzjY62Nam0ZCbfrV3AtJPpaY4SU0n/tjVvENqu7ubeb58RHnVGJBwVGT+b
7hOG6osbgIt9XuNXDI9eezFci7PbYKy21Gre4OUm+3qKId9e7m/cSNbc/N8cijan
DfDZXljbcjaL7JN1Mlsmr0YOCNlqHIfxQ7oA19Zfwk6OG1rdjccK8yiy63Qj9yTC
kreIT9QEMjCGWhrrA2URDXj2oO6IFNAHkZW0J1nu+cilOSjo9XOLm5OrARHW2lXz
/p5cnT57bXlkDJRUnhleNheB1zSWM7ibsc6l5EZbg8J1UoHZNXH58Jxw5FoWZ1E8
QwYpOljIEbQzc/hIVh08ug==
`protect END_PROTECTED
