`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nqRTScCoUL77RPkh+I7O7+FmqeBfgedRuImrXDpbHAsJOzVxR8Ig6eFuYaEHeS3
FrcFniIkzBJtCyZoKB5982ldlx4xsCPNW5it25+ZzS5Xx/xuievmVnUI9FW01V9Y
sC81FSuWkrxlRSE65vawXPTbXUOIoErFiOqgZKTpawDYgwXQCNBoztzYDJZu3VXq
4VKbvqeS8eQnL8k7pDNbWhWvGX6FNGwKz93Bdg7qgAIHAC+F3BvzzJ4LZBh4vCSc
onU3F2uSndTbctn4/lMWnolpSNJVP1BsBXzTr/+o9SdMTjgz9OifDTVZz6HdgNSk
s1aGwDoiLTpo3smmO3KFR/m+Ern9U7tT3ycl2HAbnHKPhYJt1vRK3ogrzsD4CsKL
yaxS7jDBbZapDSRNYdY1z37upzGJzTCMCDyoLKT2YZ9/oHlQ/MzTpBAxhuHdSCMv
Q7MFBdfLFf4ZRdYPRUjb+3L6berX/nAD3oyULam7JQxPVjHeWVFFSRjQs3KMb7vB
ckuErbnm5Vmgn9trdwuZbyYn48vl/c8XbV03mo7d14GkGUqxFKXVTdGC70DS80Kk
N1YmOGbqP04KgR7oGnM6utlwsGxBZmKwarZ9oGkgmB08BuhNlIIfmCQ3bQ7bCz5b
c7jQSWHtgd6gqMgonn+i/eO4HNJUmEWej7fvCwLrrQSZvT7sP4nH//yjuYmVdcQs
sGQmnnWXueEpXrl9vuyjIedZ19++W60TlpvyvQpGWOvPNu324lMs8GkgdbEOR5MD
PkIF0ljAd6Pn+OdlTOLTx6x1oox1Ti/h139mtQwDoPHj9mUYKSorL1023EZMPiO2
Q+x7BLbgjupSCb1qY6JoajqnPhP08Gq49i940ekiIK7LVmznJfMHF7bQAKa5xvVc
jzxYUsBC6oxHejrpR8WmW8lcrkeTfHLCJAfuRqGZrORbU4JKr9SP35WLH8K6i+ng
xrtWd7dOnP5mly7kOVTSZQckwdZkQOkSrPDCX1XZZhmPIiN73uH5OnaLlhROC6J+
Q3es8pWt/VTcdVsn6nbCnQNPYquet6ArxDThyzsB0SAZsWXq8YDII5HT6/tARucX
wwV7455T3VZYV3zR8PcIR5cYLVF7uPHbnRqbZ5zb0qQMS0tc1jcgyryYFRsyWygU
AKULGPNzPPpGRaNlnLhvCNO6GIFjWhgz7Z6rT+65bCMxmaCx7yJeL4mVQ+63O8K3
gJxSEb9ivslaCquGpq119OECFrmVhtC9P4jPwqHLFihhDU40h1WS4tKOzRwF55vG
Gytp9f2ywEzmZ3Ji2HuPlGEoZ6Mibd7fNA9AXo9FmfJOBzQx+a/Mw3Vnk21xVmLm
G3W7uxc6/1N+h4PQl5mxQFVoGdTYN3vHfPxVJd8sI5LwDe6vZGJM2aNVdPPQr/q0
J/nyiT/o7zSz3eRf9m7S2vFbMaDIpVIxOF/m+IoM8/DxmQCsT1glZTt2FF4FwGBC
7gtmiDCrI/hU+OMf3Jzzld2gou828Z5EdbYHx26hR2bRZ56KumfL6w+p1AIM2RyN
cYP5S5K2xF4D+gsq2EaV/0Om9qgA8lnUJORLyuwsqGJLhzffTPoDp3om5BNxP+QH
Uf5QXRun8w6wWmBIpiZcic0/M2bpOMBSAvm/g9ggD8bHb11GE/Ydw1VBSBBiD3Av
9VBNYpkD1nKdAZKl/oTqxw+lUiK8uVOmN0Gj6Cumhlix3/zhU7a7SB4v79UYB8YO
AxzmdRlADNXBok8rxRksn4BSxCYs6qLKXaUXelLoSwSknoFBHWkXRNoqG9vPp4KC
tkwCweeHO+yB8zrtWdxlO3ztuSYVXkkqSFINaXzSEwU=
`protect END_PROTECTED
