`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jh7vYY/1cdctlW9cs1dX5OHMbYcFHDIyoyN8ZPjaTKh/ShTIRpHvDibeuSjXjRp
Ft+qRWgITjSckm3hkKNGAWou4UbvbN2y6l84zbgErK+9w/maJzfkJLKYyOde/247
NJvJkjJTsOmHm4RAecaI1son7U0yzHVeZsG7Dpta/8k7uyKbeTPVsbI8BwMhA09W
Ou8M3IweWPF2UhOf6t4z5OVLFXLEh/EC2BtNR8SA3wxeZrvxRoBMhYQ9CmSP8W1r
JK5OEYXu8GL5uwFAGqvG12Njmu1KNmW+Cwk7tD+aWN6JNO4zYrGeWo/GBhhiXJpw
U22VBIOKiUpmv0zB7AmRao1gnWDvYzHLyg1BkWplClgFJwr6Kos5wd9D/oQ5QqHQ
2giuOJce4qYY7C4KAx+X0Oqyu3K6Fi1NIzK2kZkGE5GakG11UAfCckCu+vkoYLEU
iddqGDhC/ed73BIBXEMVrC19Q8B47JTqiAsAMeBfZFAFALP4V15kiD9kG3Gypfup
0E3YK1QIT0hf3wD4JUlsY5M23ddq70Xboav5dYEDb72aUH76wXO6uP1CzAotDoui
nHZL/l/qNNFeenEsZOJlnseNTs3XJKZAF9yKzgEf6KJrCAk4zNCWBm5qgvTjo1wf
VQUJ1msxxf7NohpweyAbNi1qA2CHyJVIOq+O/ivZJhHJ1y2FjnLrGl7/wEnJRoOC
3TYR+KmHcc5SxNXhEUmvjhmBGofHFUBxVrFNe06z+aLLEbKtdKTcS5TIAnktbNIf
EvZ3dzmDRMs5KLnfV8rMhmcmM4mDfhnW6xjlyEN9ZlyGb+Jbd/RM1Z/r+lqxpFnZ
dELFxXHu05nyyFV596uZeKdNZlxuoDv+TaSvZtO2W8ViLFNQmoxf18oetBOy3RsZ
cSfVb0uaJ8LDn3DxX8+mKAIGLIICSlIr0YdZ4PzIelmvaFPZhBwfhPLWqRmmxlKx
zbgfPxmsZ9BdLAq5a8AjafeG2x3nCvUSneYZ2vnd2UJWRNHVUWrxEHS7dVaLT8Hb
ux5xsLU6QS5pQ3iniZKTBRTrSJCKXobtaXlljVmfex6u0orcJaSEcGS5jVjNB6is
MHXpPoGKc04kwMVWuzHldjV2NkhsUa+E+Owwk1Er03VZQLO3bNC5k3SKX/RnT33P
6KtFNi6ofrrFmmhAgwVLTkrZKSahRrU30kVuhMALa5iBdJUqcBFTzT8IH4oX5btf
GCzFy85yhW0POUEw5ELSphahwwdEO9I0IiAtffq6tT6Vogy9DY3PX3tgmbytyoYb
Rdp6ZZRHUUTyo9nTZabotS7ZZKBlkck9c7wUvRA+TptKaw7j9PseO3qY7gG35Eg6
yq9nWaR3JQk4JLaa0jrGS9Hn8c0YOQwsfKkZE81dcYt0Cww1isNYL7XygZ/bHpvt
j5jwnZmEO9o26w1PWdWKaNcurDp+/M6ctEaHWGQdhtv8j97AwQRU9Tt1OG2ebEvJ
9nx8RU5uxiQAuhasfM1Ejf965RTyYG7nUfp2NuCcUlw2L5aWme1obrlBwU4jiDHi
p8OvegeVTgfGSNHD/vkWvNrB5gYqVS4lcIh1QQSEroPDtFrQGj4hRTDlOc/UH/Eb
KdIPPqeOcYjoAaFHcfq+jRmKZG++eDQo6qiaUvsdFFrOEW5ys3LBp++r3JSvJfZC
upQcVnPmABAzxBJAXkliwsj/kyfqTtFZXW/LFADPdo8TkqVsASo7425c5F8r/rDr
lb6V5j8vn0fBdIGN3b7mJe2+tBqvBiwh9ZtRzOVqHeMdamMDNnUj8RJo5yW8FZs9
zZNIDcAxJdrTbaeOgDlc4sk7HH7aPinUE6WKyqNqig0BjPEpJ1jy1SXdI7TsNSJM
6OImZWbCAdMdMOm7m/V8adWkgYYp7S/00BNM2HUJOBli185QEvDa8cMo3eeWOM8k
l/UBUoO4cTBzBY7O7EJ5I57PyGtmBs+u5yXOQT5HqwikcqzTd810gceRmTNqw3jt
Dz7KpKxiFktAQ3FjZgU9jw==
`protect END_PROTECTED
