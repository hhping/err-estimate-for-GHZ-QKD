`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBsYJWWxPXRi9OHVbNKv9DyTB5mtCvmq5NHmc5Yfj0NJttvWyUb6IiCRlFR12xAr
b5sfatZ/BRdFq2avX2FEXxd0QpQakeTOZHcEfPuHtexdjSFaomdJiYaWWnxtT8+2
SCscm+7NopCSMlpWuw46XyS8F7F06aN0kNFyxv7Q8fb02OADpTygJiRR1MEy61wC
dYlJlkl7Q4Uzzj8t8WOi7Km4+ZMyrzsxavk75g9oDle/rMN/X8Ojfu4XMyQ5rzPW
zYD/rFOmH2a2gM4FxawhmBgM7J4MkHU1uWZGFjeZALqn0FzN0xsgMGfuSjgkl4km
r/ybYDzCUQ9wMHjxVlAxkWGJiedmCHaabpH/gpz4wxR56hprQh2XdGQ3os/sFO3k
k9JjTQzcxecRrrZaUmp9texBqSXrM7bmH3+1H2vOoFuiuTJcLCms4uUjcOlki3je
+Y9zkwEMK/5LbkZ9Hm9tkdu+3V1S+Jj7IKAYDcdjJfLTuq8ZXfraJcts5xbW/YHC
QSsBytmR6clVOqfqIEnXL6759qwNtCa/dQvOEw4uc5hqhOcZqdEtzzIrqFzec8El
DK5lj5VhQNhhTHqiIB3nnWzyamClUErqeF6V1huIyIEDCSZeNWY8CmR3/zruWCIU
09y19uewoyvn2EXkE2qnMw==
`protect END_PROTECTED
