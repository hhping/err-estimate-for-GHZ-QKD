`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pkqhqrA5zDD2rw/JvXS7LkaaC3ILVCpGSSWBjMmwwPg+3e3/RcMdV1CPKw9Vw51
b1wNgggLJx61yNUDO3txM/tMAYUF0rS2C0Y1Us8p55uWbpQsI78jUwwtMIH5SE4n
ByWb8vBiceCPfrZfUSB0hWVnpBBPoeVUllcmBNtEL9z/zjYczxD+lg1KRG0jR4sa
SGs9XUfLw3eHh/uQTU0aEeycX4cwlGHbnbj03CxTuU/aY91s+lSzuH7VhHUsr4al
PrjH7iEC1flXiWmDjoGbYFDRGPr/aWe5Shx9E5bhzouAK4ctrLJuNFzTwZJ3/t1A
Ji9Ad82ctT4nKIfWFqzHY/85aO9y9KGnyDhqYQoiqZz0d8tJi8COMw6lAi+qlRja
jluGlt/0qrLUs5473TMgLZ8X2HELqkioQ50fogFiO1PtL6iAHrgUKIXFGIlJHp8C
xo1IoymjATBH51kCjD7+swjHBJ+F1vjJdWljNDHTOuKm0SeehI6N6k1AyzXjtjHC
JC3IZAN77/Lda9/4Z35oHX6vuj91XunNSHcDGWGlk84FMVgMgYqfL66WwB/K0QfV
iahO1QqsJjPWNwAxqC0jgVFfsnp3VUg4R2PNOia5MX3gs27sZrS55nVSoGRv73Fw
J7zRobJBBElKFmdQSwNLY9+09sKV+VPDpnGQJ9bufHW6FKU5+jC0MxUD1jLNs8as
L3h7oh1gGLT9IHuYE4l8n9LpBX0n1bTyyIo1uqFT0bz2CrJqCVyJZ5MfYFsy927e
RcjLP5ReZrP1nbvpDZ+Tkt3aHXHL1xBsVquuE/Yw3a5JNXfDQEQqKZNe0p50QdNY
QLhlFi1gsReOfr1dRBrvUw==
`protect END_PROTECTED
