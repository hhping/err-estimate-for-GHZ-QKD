`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MnUXlDdYJHbKWWQSmZvnaxnsbz+7Hfp95UAyX4Dtr8ZN1eAGVACw5Ku18A0uTGKk
tdyBK4bvwvx60NRC6fGkiiM/BS9Iz3hH0si+DzGv2cExGEuH+dLBLtt5jw5P5gZr
k5MAfSYBPwhf3l2XM+vXbIUKqdQrTMo7TI6slJHYbURWQMu0VQYtZz/Jlyh1Olys
v9vK2P8iEhzVFQMsGpefjtUiQBiR85WlpjAnprgA5dc1JO4aYBiomvqRsOQYNz4+
UNipqBi+B4wp7QlbIUSnFFPU7p6jBmeN/t9SuTMY8HJp/plYAHwSI4kBqUkLDERJ
B+aKqldyrd6dpzLVyhcg7LCD/ZD4A7nlpx9Ku0RQIXGS74/BYAPooxmrF9dtnlcX
dy/9sZqOcJzMuKGSrGTlj2nZ6l9gQPn41Hk+TVTd9bG3HAeBE1OFHIzbk+MGOdh1
GiK3IrpyF3wCC5IsPL5qwTvTfrPEOkZQhAwE6kvCZ/mt9psAcFju9yP/k9yGW5PQ
u3haU/mRAbMkmQPxB59PTjkL/PUtA6RQWFXDdC7KsX22YdpGQLS3C/nIVF24ZRdH
b1SFIVLdxxOxRO1feoL2UYf3T5DDzWyl4ESAnufTIHAlDXC7gU7QNpRjD2eLfPgc
eaDA9T7MYWOp/KIBGmv67u1ZxMmLNzzqUmC/3f0U4vbcP8upkJKvN6Ew8U/owDsJ
s6ZttvpJdqZ3NHt17JQzHRWpBdB++IY4YoNZpLoEbRBybxw2eS06mnQgpuxpaS/5
jnWnSoJsixcElNx0GN8XUCwuqfyqENZGy0Xx0Sxr3RTLqV1i9NW6BlGkQ1vbInVD
`protect END_PROTECTED
