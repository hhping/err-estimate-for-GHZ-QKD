`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYvEmN1FlsOxsxftbEOS88OlhVBiBG9cP9zSjj8MBWPUuG7wr94378n8ceGuEXbb
7LmmWFUgE5SgubvwwpMkurXsR9duNYvBrQkUrIGdkl/1Gjx3OQTqJSMb7fOnGhtP
RyEnR9H6RyIH5R84BACNGL+uwdXGwb9Qg0IPMRRrSa/XGX5sWaN/pEjNVWVQ+moq
bbDeXa9vgAfOko6GmNv0teC4iua1O7zg4V116nEe1Zrer18pkRdn5o8XYuEGSKgl
dmWvYEZhvBtJAVZgfURhMoIWThq2UC+gp6u/kNe4vGqWIdkHFwFSVcONqrKfzZzg
njHRfiNyVK1csJmnRqfS4zqqKJfPyKFmbKTqWGzQgVnTfnIFhq4deZ8w6vtG1l1D
syM6VCZOrx6W39Qhzk7ZodAQYSlcd0iMX49UsIijrTfQds8p43BB2qEqEHzkPTXH
8TUQ4bmqG894UaqcT/QjYmVXevUyNKfNzo6Cm9jQnvfeZeJ+4ioxzvLnlkImOvSG
RVTMALny4HqhDMPlIOL+bwHpCIfwukze6vE8oWuSVDDo1EhzRCi1nCcD+7i/7t2Z
K6GUt5tQxzAytiszb5EdtXVXgq2pG0RZPQmjdY9Gi/S0AzWGJUQ9Niw+61HqybL3
`protect END_PROTECTED
