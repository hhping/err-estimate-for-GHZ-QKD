`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/pdbnY3N3MGGdbAAfQa6hBmPtCCoyYghXuP+C4tCpyV8qh3j1mHr8hyLyNZgj6Pt
yg7w+qoLxZH+CIdDkh2BcQsLVPy6xkjBwkhCjw/UjDE7fSK/sFWlmVpt9i7mG2lW
LwrQUCqGyEo8ouk9/UrTwzb+AIamZXmHbKzWF8E05iBKesRFOPONxmxbBRahMb46
3Z7HB7cXYu/JFtBUbvvcDsOUetWanFcLwBJvV59M1ejNP80kilqbJh46dGY+ai0j
Ck/JcUeHGthWmfWPTTOEbs/R8NZn7zOHnmSIGVdygMJJ4J5dwEDve2KWgtrnbOx0
MDQzm1CCTAHEyygwVrJk/urlBpF6w0l9eciRMAoU3e7QzkZnMjnjZK2AcEGnTkmL
uqvO0iBlZHTcgJQ6TcNnuvpPSw29gL6TDxWhKS4KPqRVWoV0z1ud/tS6sgMjJbjb
GFlqROXz33KGft8rGlWzGG2zlbLNCX8e7rAjohDe+lhhqDSwy+0GsANQt7Imqykl
L5j7u80Ztk2ipubtC3fviYuzOiMgOsR1eu0z+k316JX5WkSoEdFqQKk/wo93tTXI
otRHhNu4Zap9cDNKnQa0fvnxomUY50YZ5C3bfLWagMbQH2tZHNBzYuzxHCxpR4Yg
MH5VKfRPJGO4WiGDPCtGT4vDBxu1hurI2PsdezBzJnh1NhKSkf03b7ZM/Qas5tqC
QNgu3LqxqiAupCjOXp0h8Q7gDIsteIDZD/+otZ8CQcwCULxXMu6vjOiorbjBZAgK
IQ08YJ6REzG7pGhh3aqMgVcy1SUFzxhJzRva3nsLtkiRAG8ghlQyJ2JjB+H1bSWL
H68S2k5wIVjRJQkeQ8wC8dBJ33uJlxonIZwqFq8xgh17GROl2k2IqkUTtYaPtVd4
GOhnX87MPkI+SdG3AuM19fWtorve5OOVNTp/t3pJM/OtbrQP5Ldvh2o/W5jKkI7l
8YRP/fphdQHImG+k6w+hiLHpBsMmw6TgH1/oDpCwIDCthIsxdloGmwLXb45OkAnW
gMfgR8LSD6ae0BPQD3JUcrwIhgPYNL+sv4MQIlOOZtLTeIy8ZkK6crsmVxh24kSQ
j11pMPtuDFGjfVDABiiasTwnI6gOl2uLINorcLg/jFOdFlts+xAVG/AVRiQFRGLl
Ik0Yfvhj2awXgxOSiXkz8TYWap0NXZ7AszX62hvROVRsS24mOMCr9dMftaRMh9Qp
rfUJtEpuDdbWhJANTF9ihzmX+Fav6fNyq8mA68oP5gmlSacSl4EBuldCv3TjkoKK
8eNbPojQbLz4YQpj3QrDibBOZiqUESbiRQHLozFQd3j4Ui9MOCeyJghfLCIBZsGg
WmD9OhsLN7n3qqoYq3UlpzTdWFCdeFX4cIiD1UP79YV6SbgpZdjpSd72pGJ+bDdF
qK1wCQmCuKEI0oLvK/xutB3j2QQmopkIAAcv0obe58hOJ41whtTbthqYdFX7FIxM
G2wx87btgG+1nxrpO5eyNw==
`protect END_PROTECTED
