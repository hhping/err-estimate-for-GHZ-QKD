`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iCE9z1a8edVkElt1EUVaJGdeN8N3uEibQzPAevDjWQUzedeQznJ49wfGUlqRDgV
ZuFUFm8Cs6fYDpHrg2Pa7IXjI7PtxOeZhsqGMS8FFCBxEjUC+Vu+7MHrxgZOgnMy
PeDdWGTUgvTkJ2MB1RnPo3ZiH3Cx4sPI9f8tAiJ9VbZjZxhRyo8JeY+pF04gDwgO
tx/jCINSwkwwdOkz6YAzLQap7x5LrJwbNNoK6/3t24ZtNYDdI+joISjTIeMMzock
R9DDYCOw8NItj/8V9lkpm9gyKN7dNAlmxiS8vfBWjDApkKP4KozZkQnpEmJGARlv
NdHl7NXJAyyo6+uAERwIu4m+aDHavaPLoUf/Zg3s7wxcdKNGhm4JVyOFiHGjeoIJ
fGxfSX+SSbQ3DK90Q4NAVrk/fvMLdEL23fnYFU+3+eqWo7sNBqppjH5crdE4FE+N
PfYGGsxT9toer+E2tk73pXtRPTu3SH//5j3R+w8WLIfc2C1pp7rJKN5RDnJW3W5h
ZG1RbgGxD2X2F5Vi4MzwrWcojtxZESytP7S6P9eVXCM=
`protect END_PROTECTED
