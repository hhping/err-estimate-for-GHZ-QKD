`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ug8ZENGo2k0yWfCf7ntw2y28/ISuvCk839YGNLsGSLu/4WbSS4oRScZs15zgRH+2
zQoQetGxO7FuyPgF/xbjPGfpoVHXvge3VduvaSH0wnmqqiCKFuAVl9tlmXvJtRC7
w5MvqAl2twC1I0MkiBI63P0Yx9YSWYtrK0+w/EHmWlv+Deg/S5VqBKyCs4yZ1ZaO
z9pJK1yfQ++erbQXobcYL9l58f0IW3TKJykRRT8VJPlVPNnzDkiIyavaQziymwdy
keBl3HEyJH91rOw/6ftsaZjZi5TLW9vBmIECk1ElOawyOKdMRjTc9Vl5R3V6Iwkn
rWWniFsfZXJdaCOlxhQJTFHGOryRcJZC1IrjUzRFHLhruU22RQViJcmeftyjLiOd
rwAsUWpxutu3ptI+8TppsP0PkWpAD25gRB4vpZi3gVthAyZ5t7N9HJUUKoTS9QA/
tPohKFhCvOimZHCFmv7l538EznBWGVrsyUlj9NGn6yPpECjc2Nej0zuFZugZODt9
KoR3xKjgG1fFgD5lKiPZRh4PjWZKMJ31y1eAU65u8bG90XCNL/OzzLuOVum0arPP
08dlTYuGzxA0Xa9UL3JhXqkOaFpASyfw/8W6D2/C107M9eQ/OZoog1ICrtgI+PD7
gUCPElayLf9zMFpkZBSwqPuC+92hb/8n4nsvd5rLq2JJRVtfWDsNntBu38DEq+EO
9HBCQwjWToP1YwwVCvBAlDDgM9OgLiBPErQ+FaX932ZvlIVMY6pcHVOr/9fsptsD
SwM7iRwpKTBRue7lROR4wo49D/ZdRHrMHNpGSzhv+K293sMNlRGby0k1ns4tqZyj
ODBv3P+l4Qgd21Pp1wLdxZ4zbUoxb2EP4gal2+bytSA1MRnA6+7BrSryYS9bRmi3
6JWACaI2EIkdd1r5rqZ80G/IR28qk1OI046zfDNjjtsQ4nMYHQYGIRrv8ls/98GD
bRqNAycRQYXT9y1D09DaUYjs569ko/RIw1j/6t+Wi+vqoNkCjgRE2UDmv7gkA26T
MPo+blpjQmQ1ItBTgWTRs1Tz6EaIzpVcMVDaGKmhsLBTDtC73AMrNH6z4N451VMi
`protect END_PROTECTED
