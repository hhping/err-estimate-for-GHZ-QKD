`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
imcme26q5RF3btc71a8hStufrqWr48CWtpW68RdZJH/p0hdAmi9cyLJe4lQ59jVV
3NjGWC9kphmf4SE8UBIlvQW9ePK++iMs4kuK4/+ANULnlOpJrTuY5jYfZN7ROtqC
GkbVN6RQtML5GtyyI+LArtaGqglQx83hVYcMzC0AHreHUbaKUtugfsv1onjgtomb
t/1ebeZe/T3s4MC85jeIZ588LCetkVfJIP4xasYVEEIsB3hc7zB55Pd+ap3NPXGB
D4SWyycRtuJcRDjP4CFh4+SUA25M6AzjXNG+FfBKI7Y8V+9KMxSN9WI7zLXfYkQA
chy/VvN4LdXuDTubMdhU+ijNYB9OKkgIA7wyfvDg+SBXDsGsZcNfQrW0JRYFa4KT
6fpN2oBqZ+LzSr8+tSi2vLnozyhnSUyeu/uDjQmCyV3UGb3vj9CLcMRG1vHyFJLZ
5VYGk9vkDzBMHwClNGDQAos/DUQRXdOLbUvRrlzlURkcwZsr1KF6gr+OIXsOarOS
1FvgZdyqYcyP7e3FGpeUH3c2gcN0wTao8VVel1dSfg1Nys+sOoJada27RbGHGB9D
DFEliuxml+xGtqZODg8qto1Xj9QpqZOgb8rUSSWMKgBFpeui67z80jgYBfDPwhJo
7II7HUVqAjvSeancTV+rzvKQdXaMeWhu1gFHpp8s2wf1VV/D5+HzBCn9L5WWuOuI
2Lv8h5IPH+KWVbiwYHsVq+7tC71uP6x8FkGpB/1CML+9g1XqWZhDzOyRslk23JtP
Yr+ip6I6MKJRA33+SFWvzwiLr0P+bq5gwe0DX+AWmIZOo2Ow92pejJ2sOqvPvps0
E3dYkhVQRwf1Ko6bcvqZrN1cC7adonJTmQVqN85gtxd+i/R0FwjDgVeKMlzWajNH
+IUCz/SIyLhtd4Zw5LtUHO5/Uz1/xBQXeM9/Sxk4OKTYf+IoEe9oe4XewsaBuGe1
EvGNg8adwtaw2D3sYp73Nx9HlbabjsSNwwPp8+mQZUyl6S1ccmpUXi4caoqFXr6U
KUSyLuaOQGJ3B5GhRywuwZBxT7ka83QwaNVOYg1PuvLKORCxAr2ul02YeNmpEa8T
slNRuZwQBkmyfEZBiC2ZFFeUTfVV2F7X5fjyLgJRY7/6AOUf1bGUhR98H2myqY4Q
KuenkTDOn/Xl7V2t2KSXGzfkM570/NVJM/PvPJYta3D4fpz7rRfUSorzh1HISE6I
BWI3LPR2VXpAlafLHu+6ErRaEFatrsfaNnkMhWhgFTV+GCoOO7AX7/aYWYO7PrCv
9NPGodL5X4PEJ7RfLsD+RA+MhPkm2Fls4lmH09t5MZKN5nlNtR11bFFe/aztEpSa
q3QUip9PCVl3ErYoqF828w23NpfXqYoESoOp7p8prZQzX98qFeSn5ZeoUFuWMN4T
CFbYg2e8WgZFJMTOVjW2HA==
`protect END_PROTECTED
