`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7oW6Z4B8yfZPYsWL50an/ouHG6qfN/4R+HOATKi2C2txg1SMIMkez2Wc3PlLyP+
AQWNELr5u4j/zh9+TWxK/yRS4NNwCeuFRDf+oyStcM7Y+ir/WQFNvdvxJZn9JfBe
FfHqsr0l+Db3CqXwb99GYsr6sae958NCGpeSejxPqAlwn92GwOmRLOZP8NyG+TLX
`protect END_PROTECTED
