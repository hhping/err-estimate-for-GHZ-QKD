`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxgy6B0h3XQ06YjHb2auyIA0e+ieQIT8SHLeJbWx4QYvXbZY5I/lh/tSAdl14TmT
9l38aH6PTCsIeTW7V4CN0DhvD32uPh/A/lVmPTRNseDvariSRLU4IuPpswy4QdL7
ZSZUAbaMhPtbm+qFl1Z0rXMgAg44PFrVFw/6YRbQjekwGbjUO2O3GqFd1ugszmYe
TKoHU4gsmxYQQCt4TMwoWQRR3G8t1/qi8XJyXsJZNDWWdSMNHLdr3iFdHnSqjUgX
lFFQESPTGdnuzOzFjsi6yHDyyAemk45stRfLNLvsGiHbjh/nubDXsgLnP8HgjsVJ
mfWLV+lgAbnTExG9GWhakoXGtFvpJmPlBI4o2gZxPbmzEDe/rcoX23qmo2+Yluib
jKYpy0Gc/czd9pTtYgQUfUeeE5tqrEvh9wSU9igGz9GRfCj+xjz14LYoEyLY1mwA
GzOx87qxOyPsjauccuop5OeRgJc9smzfqHCZTYGM0+dsbW5gIS49gm2LyRlWRICW
`protect END_PROTECTED
