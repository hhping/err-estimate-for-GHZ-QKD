`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TDdu5OcguQxCn223jLwadDGIixM5sFJYqgtoRQTg0d0faJ4yVI+NhTlc1+r5/4rI
IZ1QF6kq/8U4BK+UL59EhiySsj8iRWEJS7yEFJR1mEVkXgkL+RYdP9ErS6SUl4fs
HjtcH6yxxGmHX84kBUC/VKwpLgEI/QKCHTFepv0r0nMpfXqaTFzliTOoTdOYEfyz
BXh0xNCofcXAUdgS1fryUt6DwMsRRED5hlt0ZzD/qQtJHmrfbduATveUtdLw1ICf
zWmUuvMBuLKOY3sM0P1OHVIv9OiFcP5v9jRTmv4pBGdXB/vB59rU8pE0WKS6Upli
2BPydnC+wl1r+ZGbZ0htoiOtGX20P0Z03TE4cIKYQHPQLZMqZwGvvkroDbMtfP2G
Y+duEzAn+ZiwvoFSGweNW8kjjPubyL2o+wGXl58h4ceqLzQ19fyaTGCkKBnt3XnQ
cTT5dGuVSW2aeosDlKAPSl4wRY7AFSaiBzN4U81KuKBwpBQM/xw8rsnbHF2jum+4
lwYG6CgRDh/CM7fEF4MIYGHVKKsn1WnHwPWN8GNAatzj7PtDL9GBP6bfE6Vttll1
reqmjxyT/pDK8P9MrNWCxbgDXdk24WuCB7LHpy8wNEOw2/+01qGKcT3CsUcnheqx
QRoCmKdvknBvA3CO3ScHXVZ+ULc3wdd4a96Jrfn3xrASsb8Cxs8MnmDkzK+6pGol
9OVnv31zAnOAk4uib5XM814JXEpHOvIqTTLijD4w6O0=
`protect END_PROTECTED
