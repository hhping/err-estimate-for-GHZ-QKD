`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+x8gkOGf+xH6TjU+CBJ5iW3iQVHgIe1jKgTHKLrDjcNfbYD91wUqK2WdJADOc/9
ZCnW3/F8djRaEej2Xilm9tWr46AeE6BgKW36Fv32CgWm8wDVhPoaD2HyCddeXWHR
3ynGoSXx38yDl3Xh4tQ1LhgZ2NQEVkGr12fgc6/rt6v2brwbf8DZKtD2zuXXxXcr
DnFqUN/rio9FLi7IwI9Sj714rWnlLtegEc5oKkqYXILbREt0Djs/rbXJNzXrYQ/j
Sakr0wcR8rbPwy+2ERnammVro1wNEH6xEhOesl1uZ077JaMZQo8KpBssEJrSTzBm
8/q89KNJV3CaBjv90FEcthY894wSL9DjUMGKGOdcyn+oF1e1F0sHOm8+iFDwkKrG
VzS3vauuJSCb1U64xExPoAPZ5xBCcc/ogLlNZ43kN1yS1FZVtOf50awvG1sfdgIr
/ZxWgdechPM1a7Zy0lUvW9KbLSaWpgLGzGFfexReXEOsq/tevdCIfn/4zLjQ1ZFm
zQa/wmMpa7CAVYLa06dawpJmV/XkLvpTwJ78I+W5urCt5D6d6FvZlDu5QFLGd7oH
`protect END_PROTECTED
