`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WBU+sRuvUtP1hepDrwZZGfamDKD8JLEDQaZLV6Rf2Nm9T+ZowztkOoLdMymnPHKu
ypEc1BtlLVE2WqqQZHGadPyd0hy1vL8odF7OuCsrNW/Ys9yaZm1Y4QlvkgJfhpqW
Ea/KzVjV26a9xCmzQ5HEhS3zv+chN8tpAfXUGyxdhNmlhzyuIQnPUUC7Fi2VWj/s
lyPJ7+c5nDyUNpzQjalQMO/+mtJxiEPXwTfqKdJriCR/EgoEbklSJE4ScP4TIpa4
SBPAykQH08s6cHw9Sol8zr5V4yTN3ciYUiz3hZdHvSXtqKrtt9+PFaUt1kxo+akO
lu/eIbHgwdMP2y35M+g1YeQs1v8q0KEYhtFkvEcoq5wuAaBAI601dyHy+t60efhm
3INgnt4x1vMIP6m8b+74e0LKgijuL+8/WmXyD8Re5eVY8Ihu03LlECRp0XD32IEH
uVJhyk7OrXHjj7PbegTW6NHm5XVmq1V2Q2CvKebuPIg=
`protect END_PROTECTED
