`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ht2BOiypTz9nFbSVD6j8fP3V933nr6puutmXgquIKVV4ecbQdDsbmRKmfhbYRRE
W2I/njZvaGCWjL+BfvMQf+LRgZZGZbkGKkQnlPV1GIC+NS+taOHGOf3EC3pm2FIM
m0tEpuJh72IZHMf9nevShG12j0Y5GoAqFxmA9QQs0c4J0siGyC9BsPS8R/ocVD2S
cSas4+KrA7m21JXKcQCGX0FYfla1Hl6Fu1O9muNyqURQ+58mXlQntxdoQiYlc3Kc
D54gyZ8SJfC1seT3jFOCKLxMiGpPaaa0/7L4ZB8PUXAYQUr42xGPMOePDzr5TM6G
yZH5CJMw3KaJQVspUHFd246B6rSyI6zjbiJavgdeyMd4hOhx7GwDCeRrawFrotpB
DqOXWYZUFhhMUFhCm5ZcGSz9n0LgMUQ1QqvzD0T8DXcWu/HqwTfmsm53aKvI9Jtq
KF0mjYJWBYZNKZ03/y5dSZczHwrkLBe5sfBgprubDZc7tQg/gHQJUzRdDo1kXKAT
9HfhvxuzUXvh8s0vNt9vTAcR1TLyaOQwFktIe52xFRG9aR4bJP/YT45dX9o+A4mU
MykLc9qAlTEjTTVtGbrNS9FJL+IxDMaa91cYGD1t1aBBfRj4hOFPIDdf2sgi0z1U
2y9+t+ysrutqqLFgIAhKTX5tN+OesSanKNxCI06zXUc=
`protect END_PROTECTED
