`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TRoRf1mdTPZIz4/9Kk6N7hfsqZhGTy4Kor/2vPTUAcH/IuzhD2ASqZfE8JnRRJWX
h02KYdGStvU7tDorKN3S1noLZFG3ePpDLs0uOge2zzw/TLCVMWEnq4v6J8cetwKe
z+BwYDPcmOuP5lgmaNM+nYJpFCUXkGQPh4q1XwhkpX+gbWbiAqzT0QafnPIHBLhv
wEY2S7W/FN4qsO7DVKtRjiTOKeKcgzv/NCodppIRKXHJ8oOhrtWrtuC/KdAl5MNx
Q9ABEmr5dUhNbPh8dhg3IgUOqGSzf1E0KLWGPvsVSRLF+jdkZnKZLFSJEGld+whI
qfeUCtT203VmVYNteUBVN8bJVDTJx+uw2utCGS0fjWRDNq6+O4vqg67Ab14ZOyGe
Lylp5g1jjbO1WFg61pQjZqXy0gjAnCA/Hp0cGJiazNX8IuBlqQ8YzO5JMpm5OSPx
EgOyoD/e3ZMKRf0XnrOSrT/utkm+xRYEZA8wT+8jyonZZ7E7MWDbo778iYZiMNLG
oPn20XkYrcMcJnWCWqe3hJKjg9CoA4+U3ueXHIp+oYI=
`protect END_PROTECTED
