`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNF3hYN55QaeNQlS646OSIt+55+f/90xksoL1+kruPOMtRaeHh/J9axajXQaWTnd
mDZTA3Xgfu/YoBLRWTfsPKu5YqGC3KnsDmF0FYHcB+N/TyA0L/86sc0z4GMGi6nH
Fv1MZF1Plt8GR08CAHWmEEUEMD6c7C5tkmrdan5sGesgS1AlCEvLIiMaXGgadpWX
OCd72iHnoZqIDole4kNPHDn46lq1XEFjWBdoPU7b/nNECFtx3UTnOE206yJMu0wH
ENpWjDw4agOVKSxjc0ZfhrnJujT5O+JzBUbbEc2CiHcK0zRReFwFYOOX4J6LqTOs
95BwvHe7m1tUidlN+oZj3vfTNHHpHDlcR/pbYcD0nUiS8RB46w3JMswDQ1xikggF
bxnKe20IQFCD78NbjWGVTUZkw9Y8XG/8sERcEeqMFLmpvMSEL5ZS0WsjjvRZaUru
Xzn77BS8pNTAz0Og75I+wD+muevNgu0Vd4UvwT+ekiMkc88MqaAUfM5d37KuqjJC
f5dqEbM7HKvDNRCSZqqGnwK1zfubVRmb/V2dYY19CjCdVjJJPuXZDjphxWohXGlE
tOUHWCeZpzwaCh5nUhggxu82K2zL77U+fqedmaAUeo7qXWgNm2r9lzwpMe1uGLPt
NdIuD2yXqVfkG6TR78yCCjluDmFxV8XPKifPnCMZ+qRW5bTu0gnbvBfitYZwvh/S
5/BtgCWj3udN87qZOyFPUsVs3sWGTJseJbcx+qUWjulVgyXD62zrrvxhwqZ0Wwqd
5u66HykujjPhF04ekcGjuIx7VCO6MWB7vQmNMHVk4sC/LuIRIquOz/vRztAbpnz/
udV46rMU+Gjb0Za98FVfQJOiG4OaxmRqR9N55/fnPHhbBplZbokiTaV7Hfey9WYF
hQr5DlJp/PMN/9kY4ASH+uqkOn9hB3wWifySkchIZ1/lbciySnlTiC0RT2OoMrV5
OfoH8DfHVbg5yhBJvS/2gdHaDLzQb2iT+Hlggk4j6iYIyfl9fJhjrECzKm4BREzy
9UUaghvFwtcSuEnPKl0Ebp6Xejx8d41UgTAPwNc14tAisP4eC4LyeAJgXILX2LFU
N4YMxXeMqJLEMNjpTOQAOHx8aBd9YkDhaNf4bPbspDTgFt28LRfKeD3CrpVJACID
agO9dWg2xvBnBfu+zHZ0RQSf/5Ry0p7LTRXA1dAvnmd2SAj9Jw6qu2XOo0jqK/J9
fgS1YjXzRosVm9Ijk/PRNymzkQpPpx+IaFujTuZLAU8yEOvgJVPTY1QIMzrZx5A1
jQXxqixkPSc/C/Ax8moe3ZIvsVbsKgvLEFcIIKMAlLtw6Wsj0GUsUwDKtKGV62Nb
`protect END_PROTECTED
