`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxzPSSiXb6koVRkMhxhocSYGk/vNoYzngmp7jfnExr8aGrDFjfah3LR0dmVQUM1S
WEBaUFctrlxk5tm6ZlnL7+3Eps7YLb/aAQNYxfl5SwX928bqHnNmb5+PwfZij68b
4u1J6xSRBfoPIf4Ss8aZG8h6Fi4+eHNPGAqZHcC8fhlgxu7Z6812/7m8ssQ88oPQ
gxbLP9qLjXy9aesQG1OaFwtm+ItyAzjAh9iKVQepvJfvwFoOYWBlG0AP7UTTYzBl
SXlVXm+1apoKnJ6laa+opD4Zh9j89da9nVQUFlZ1xAH/3VdQ2JdnDdXkuuiOXpa9
YFjulQDSsqrZihOEDOCl6UDrApgHV8QcSNb6W4RAlURG0bFK8+f7jRb/0U+wXqza
3V3k5gB9IssMgE0lySggW+xkCPTk8KPH/JTUO57I8rH/KuQkdNqYK/gG6pL390Vn
loWcf0QlGRsdnsolpd+O1ZIKh5LU1Cnw9IRv1TKGQ9gG6NeknK0Bv8p0J53tMwYb
jHLUjWLmQjZGOXCAyF1YPNG0Q9hCcVb14df+6atkl41VcEWWwVt0psV6yNAzLYCR
nfNdlJtSSi/2/t6y3oJJIyG8FwRD6/iMiV9S3++c0nX8Omdk8eRsfEqmdzHAoS6E
1jqDqn4zTQ8u7JS2tsNo1/9PtEB6WkvbqoLyN4mrU0DIW/GhnPnbgqPgVEWW3gIF
9ZOqyZ9qDIVmR/QMjVyz/+EWn8CkD7WR0+xxBPbyG/+ql4i7mUZ4smH6Kyvj91e7
Yr0vmjxyg5DTwyVu4IQDnB1ZPqU/ZMT5uU9I7daSs52+Ppi8oZ/nbkoG+3pmb1QZ
PkwSCg+YJxRDDDgwGd+OZZTB6Y91jsONPu4ww5AAwgmBZk2PhwNE0yJATvWOmzjm
+8VC3BGQXLlzibuEU+CJYORdFiyFoYdhNIuiPCqBRtsp/wZPcr3g7k9utcJCw1eE
0qGi9+Ncu8CexaEQPrzD7rHoG566fGMhpagr7d5acWkCgcVSAvDIUxRotCHG+kBJ
CzQsYDrgpqiw0RuAo0g8NicQ+ZTlwrt/h/sf5grUOZgTjY1uh0awBJYZcZh5lxdS
F9ahE7zbNK6q3uwHKiAyhAJn8dp9dY0byzUurozWlMhg9IufMrHMUjuklLof5pRO
MgLTJJQXiIK4R/N58GP8O4deyfr8UNccd5wy2rnSWunk++cDptdQKAQfaZHc1WsP
Px8RqeK+c5Km3DqVwy7FABWshX9JnllKuSSrE9gHqp6UWf3tXfMwPxQyFxRCF2av
EJHWinwfH2sydW13ltmsy+IbiGlb9C7rqjFxSkgp9XJGWQxyaMLWcZcAOjLGsqTT
Y6Hbug/3/56raOnideAlIlELrsbo6jzPYZ+GC6CdHTg=
`protect END_PROTECTED
