`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYJwAuCWMMshM/NJpZ7/iM3/biJfs2QQgqnWvbderkfpjOeyrdgIb2Eg0in4fei7
CUExApx/T1tW4CJ+EzoU1yvhTTdK7oDn8E73myPOJejOSseetVhDsAcCaNIuCHFl
WA9ihVF1r8tLTWrxQARD/RW1oWUF8mwEuCaqkngBRoArxZM32l82bOvDH5DQAmTb
e1GkGbFsg4HHMv9JfHVctTBR9FUc9mcy6acFOAsYNLLaaA7R8FRxakotzi4+JTqE
6arU/+0TkfCH91R9xDFXbtvG1OjqpRU1VCvzvoPGFjbPeNrM8jp7yQyRwVNYW7Jd
ZRmBQ1BhsnVK8BEt7mTxrKlXcGmWjB5sBp7Fvf6/9KBbSJOlX6gTkAYOVhlURny1
oRYExuoa42PmQQYGUNhcpMAki6pluB8IaYnXJOkdQqXsG+JbuVTP9oUkCxmCgSSV
B7QEgrEBszWffrkqw+ofzad0tJimd6CY8Gv1qpGlwEtsJDWPfMU/ocuGTP7mJhNw
xUWir+aOwmGm0xiEQsFZg4XdPfC2CMRer/PzRcm4gpjmdtaHfLUpgHNTz/H7A5DP
1ad9grBeKC9gcYLk29lL0DK0++glXvavJY5M/aa0E8uZmjUCymCDoGj1uGFhmNZE
s33/JXcTVB1VR0+qSmdCNnNUACa/kUPeT47B3qg+jUbzWcavno1mifBwCVm18kJZ
4BRGOTvf5E+giYGShfNAlXZiMSrQoFGZ8Wt8h3CEOZZqPKq0/SETW1qxKOaUqgwW
7V/51SUVNRDxFetMktEDdvJJfhl0xBTZ3fE6Q6UorkMAsoMTKz3CO9x/WYuuIjib
WSh3Xb8PBtyONwHCy8zD4Z6MK/mUc4wUXNW7H4e7GyoYAF+B5Tbjqrt0z8Bj2Fb5
hk8y57UZdURrikpBUvgpjusuModoD4HRV+YClswfPyLmItY/Ei/7hEU++G7jA8Sx
JzhsGreOXg2pdNaJt/kNNBuYSQx5+3eg96BaojBdfk8dHQh7kbromDY3vaHD+/Ww
q/i4R1D9zuJ9mHJjknqOtKjY1lQx9jlAPmE5uH+mCoI=
`protect END_PROTECTED
