`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16O3sZQI7ExdR83yICQJ5EMRPbXhPQP7Q6LwBZFT594P4GKDq7PjYcl5Pje55GVa
THRq5+SGvR39b5nZQhNy0EoVVi3Rn7WI59gxC1aav64NJM2VQwrrUMnBO7zpO/wU
n65gmclPRQ3yz6Z4S6TjgkQ+BFJSXnhfSkfoqgfgTbjT2WGcCLBiWLm1t38QQ3cS
+CuDn/q79FbvuvM+6iR36VyWuLsoPLX3EY8uKhJHmx4kKQP9GXFHAuxkua6wqSnp
bdmUSlxcmukdbtJDV6U0LzmxSVhHo8AVKvAip083jRkrmGXcGrfez46pmSBcX+AX
FvCOEMpjsfmYrtk+fmKoKcyjEGMIcEVSU6fU22AduO9ILMbFITXeIP1FH69H4Nhm
xuYB5zmR21BTHFH40f3f69uC/6X21dXDi3CBJIiyC5kZydZZIJEQSwQ+haIdztFj
cYPCr25LqvQWA+otpFwuoS3viU0uS++FlEdqztkM2K13B6ajocHIRqNway6DzBhT
Tppywjoq5X5LvJfnDeqvc1WEvkb1Rf4nk8e6JQbP9/F+V3YY9NA6e388iF0mf+87
YlT3gGfm3dbtkpvHtu2NAxFLvbqDSgHI5Tap9j4vpdwSU1CiZiA8zWaiLaLN5OTV
`protect END_PROTECTED
