`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0isEmm6i4vxMlUYWLALChNtwgC3SUVionoJ38UxYEYPmGAI8yo/tMflqe+o/weun
33MmylawA59t0ZiPlFxTVHFGYOndEnCrpcZ6nAPUixtKDczCS0TCF4oNUbOeRYFV
15Nu+o97eGBuEOh2VVqF9b42S1UwQejf+I80uVEOSPnTlAkA90PLK2D7NMcwOCY4
MrrEj5vvLCUPzu1YhuAzGJMG/y6V6rAXk+r7EVyPy3ubGsyv4m8f8HKZhFKd0eFm
Qs0k6Uf9bJPFlp4vQT0ytLte0AG0tU7b5/aiqQwfVHTh3dS3NywZpoEp0o9MEEGm
t3g+I+sRmFQioaamGil5oi8FdV7qtI0binZ5RKUN6oG1ddcqiLL+oPe/+zKCbRDO
AAaqeV4kqgW2wOKbJGtqxPhusKjxMqHOY6Hr+Z6wmW7pS0zfO8Ij8MuV3fYevU+K
Rck2e9RDH1puNSPar7S8eoNjxVwPayw0wM0/QZI1iVqHXF6ZoCxgwxc/dS5KCzYG
DmjCsImQpQJ8GsV3LPbhu6oQmWd8wDzs7gq90d6loitoPEYBAxR/YruTJ+qWeeh3
9D58rF4BVovtOUh4cat5g4eGtGWBKqr9jZNZCh39em622/LdmfG+HrUaJxPggS4U
G+6RFoisbHAXgeDbG3ke9bpvLjVRO9SsHEXoLayHgY5BJhjgWEBeYJAYd94eApwP
BWE7hjbisL5akz0t2jJAh07W8ip6xw6iRqpIRDzDs7G1gI8su/jLMDTB7ogc3hUe
dyZRWSFUNOEuVeJp2p6gG47myP8XlI2yehs0+bPKGGLMEVNQGCFue39XAggcwa+p
bwYNC/MjoeJZeFHenvq1zuEr6V7ro7xRgor2hy00TOOFK7HtGy4tTH1PGjkRqjwN
vRADrM4poHoKqstZU2F4kO3rJq5ukT5vnrnz8bEMpbve44t66wZSwPJhSTBGfhdM
spyQoTkM3cjhcA8VV1jKmLvd0vEaEVS+wcFF7EEX2boWxSKrPD8ofk+Yal8tMsCh
NUNp2QF6UHxZUTrGtrb2Pbrdialgx0fEimmYuvF71Wy9MDYO0WnmnxvVTtnx2eug
48uY8rLPuBOSm7T5ZU2zF1HjJELKvWeHe39awhdHEzOXKwo9yMFzIii2uUgHVOzc
fEwWttZVRt8cG23bpFy2p4qFYJzGuIxrDbZxX0HV7gs5PLTFTTd4+kC5L7YJLtvV
iAeJ2gtQLNmxCVcIBwJ2OKANKl/jXNTghSCxmASQXBHa1ggWutJ3IGAjnZLzjKGW
5LBt3xL1ACeti7Ufv6PvitJvZh0DF5rRqPvFT/rjSaBTlTmzx2mhZMgCfAvyc/Ya
nLk/6M5NT8t0YKVzMZ8b9R9ij4A+1hti/MVJrTsjwkwsr7SmggXb+zICUvtsduvs
vrziTznsyz6hJfHFheTEL2ut9rcutEvG5AHbE4m1DQZVOa8MyVFdkjJh17naRRw/
qlWlWcJ58GtXScBGFpd0XPE/6cRfiQZQ2jmmqwgUd8SQno4ZfFiBjCutIyRf5/yk
tA72PSG7LJ4umaLcvtxtQHwdu6DG+eIb0HHySguIqy/UluNyZKMGWcu60wUuYpWd
GHDzS/M6uI5yoCTgY7y8UOm1Lx7CSdJgo8QMD6QAzJHBAIe1S2V/FkpTZvyCVTgQ
7LgF60pujvlqduKNlI5z+EStPbxJdBQKtG7M59C8JAgQXo7hNj6TjFrvxVXYUUca
mAasZ9IxIirMnJRpycfoMeZnaKFkRSRpwSoW/QTqeMBDHWIjoWOEZocsf16jH5IN
8vp3GcTaV/UWglBYAROUNSZU+t4opNPoS4Bo/wqbCEBqlZYK+MkBw/W5H6EHiN8W
zjcEK/VoYS8eC86xtFHjB0+aGunVR4fxBMOcfNQdMVkGHzkzXrzgUIjsH44bCtl2
sTsyaaXrhdiDulG4s+eokZJLeRdck/S64vT1H/vKcd+4F77Z57vFOimFk9hQQhW2
isQueb6jYN3h9pyW5fPY++qIurXXclAJAIi6QykVnN7s4jHRdSfzXLoEHsTBpjNM
7Nhve743eNRsB7YEbzCICIBXD00MWqf9Vw0VIRI3IT22iUTFrQPYEwAeEcsCwSBr
f7jN55AzeTrkl5p9HUbuJ0OvdeY5/gZ8OY8+lJOqt52EZ5sEomZ1exWGrjHunVkA
ftYpmq1/b1p9f9D0LsBdjhko2hT5EZk/HlmLxPfdva+JtAEp+bsTVmeSvCk1FWY0
SlSxTyLRM8BfCpwhZ3so1UMBPtI3wK+5OAPNESimPtk1uGCD9PWOEFZbPhO9+H+Q
`protect END_PROTECTED
