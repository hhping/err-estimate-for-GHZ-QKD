`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqX2OMdDZvYNi1Zz3GLReyuenkkHgvBIDk7KJ2/zYhbORy5krrO6Gl1i3wWBf/I8
Iw6ZGE0SyNqJV4Mg3kv3zoMSCC79z9sRM6lMepJ0mDYTui5vDxsA7aAjjsDcMKru
JwiHUIQKpuVHefW4zSvde1ZfD+HNNmzAEAs/r6dyeyYOnVbqkWkcV5ddXx1+RNA2
CMSkHoPh7BEQ4K231rHgNzYkqcnd+avtJPKd77TlCnqEOS1ZD00mf8gQZEgtGklo
D2G+RolyQ6qUCDaaMuK/P8Gm0irn3R8jOu+Jovzdk3jnCN0jm7HfGa84duR4PZwv
zUV/spZfuhvxH7XaG7fj5HwUD1dUvI6pzLCv2ITDUyAPVaWIYCv+4hDx1UZh7TKs
NXCjmET1qMSMtNSwIdRIRFFp6I7xJV3AwYscLgurNMNsL3Q1igB8/RHRqECCLCn8
gheAojCSsYUGDRvlzn5nLHaZXxt38oPMYWecg6y2EiuPO+gnx+lvXsvGHJkoRiaj
`protect END_PROTECTED
