`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YiS8oSH1/WwavAJRiOliGg1NaXMf9KSDb6vBgv+XkZkHM8obGV+zJh6JSrNsAyI
eAz6X9y10KcYRSBVk9OBYLjFP64aGxre+6ugJVhg1d22YLqJlj97Y5/v8jaDPoi/
X6uBaWF/ntAW4rqDULW6Qdxbs6sbnWnIhz1pC5JjXHqo4K5M/cI8jM529XXwByXf
J0vsS9AuNBBJWjyf/yrzWwOQwF+fUIBiOI+pqGvFRNKfw/DsNJP2dZpTswZspGEa
1h2cqEayJHS+MjOnhKavgB4EY4FFcryxahORY918yhv1VHvpiyHurpy9gT9ByGEY
DHjej+D+c2jiz0Q1B445TUZiD/SS2JStriXuMYed91rweRKAoBlkoPzOqI3xjn/4
zmq5DfJROTRQVY4EBu9Xo4pwtv6mql5NUdRgsgUQyMgN0QBIrRkb1eIewnbM4xHn
E9+peD7VBa5Vf0MtMIBrIRL2ofmzOY4KPi5ayFk6Y3zLTrivAw9Gvpvl7q9VwXRq
cgxFBCwhwSh0IrRtinrlkB5s5NdQKQy+TNTuzlZju7OAFwpcIVQEzwnR6yBXItKQ
WvpwqJdD4/zJBBD3OyFeElgaACVxXx0cd45mmv+nmseCInFts0QQUtNp1lyijwxn
m6unFsSdmZpxkiqmu4kcl2Zc9rhWXLn0H8I3cXgYoGTYBcJreQVNSbH1M7fKR5Dj
D+zRsxY6MwOlurxfcBodzw+m2h9McSFlO/riTs7uv0vc7SKsLxTO5tMIRUshgMmH
Aqv4ObDHRY8a7pe87bg7Iq8L6lBnZ8SVJ1RPp62yo5ifLlxLNvn33UCN5k8QxiJB
b1jiHl1918qqpLpm3zJeEaiJ6DYkD58QyCdgX9CF2YOFppqREIx7vWrk/Lvn/MIb
ebSsW8bVMvJdwxvh4w2/QUICZuPhhioreA9CoiEEooTTGx1vBSjv4gXu/F9L0QKw
K2kU2eTY15ssaKHFxhtNqa4I7DsPM3tnaLbEYZRG245N20QR3Lx/mrQJ32wBlCGI
THb4mTwnh5nuoeq1bAhM8neXaiCrUbILT3H0hWmE2SXcMiK9+DNnsqf6fCMYa7Qj
4y2+hYvvlBZ24MlO695c/pkAaPz9aab4LCZsx1R41hym5uKhaggogayTr7LjYAEg
Msz1icieSFYIHMqUdTDao1CDccbku7AwbuEhp1I7c4lm22XFGtB3uSWAYVJoN8UJ
nnAeAO554JOjrEGHzjz5oyhukMyjqvp8wmY2YLC81B3QD8aQ64wsVgZzjdf8rRGA
lmlF5baOBcaisoYGKgzsj+9Q1i0kSAgeu4RhppuEp7tXnlJRPeE/xR2ebXfESbiB
wIqMDVaoPNkuvCm32WvG2TmOIOE9tZ+RosYLbj0lkRBCKUf+jS9YlWV3An679tQO
dY+5HZ0sOmLmP6R/ATABWtXPheWTOQ3YW4l6pOuazU6JlvcmtNeUOu8qegfEPZE9
rc8XmiO/qF+Vqgcq9ukuKuvxJ+6kmIEf/kvW4lCmq47A3a0UUN1YR8MUsJHL1v37
ffRNF9wJX2I4nSu5I5Y9agyvAkz8G462mmOzD4SygKvZAPYJOnPQVsaAOA5leKHX
7nUqRjMIAuqPTYKgycnPHk1eQtXArbYrxN8Fd/oh2kSqMiVGHS9dg/ydFgUo2EHD
O+tshQb2oFyVbJisOOtke6QFjqWO6k+nezGUTeml5s1y6rz/fovL3kWz6t67yoQf
LhzvTQgqbB9yvArGyeH59Jpdt6r/L6iGy58YjcysdblLGSco6z3kRxkcl1fRopnz
mbVCE8jDy3dNnN0myO6HQtXdYjbavhoHFyu+b5KgfOR0S9KQCDfYFcYKAW3bsuNw
Tw5jmmGVM2AylTDlVMnRT8QRB/K8JTOl8JEIGZfGJgwS3Fzhu2+bSQFwrgWLazwI
w6uUx/36SY2r1qG28FnMziOkfk5eWTKZxvJw0m40cIXrkxgLq/JK/P1e6bfdLl1H
5YjZZHZgEgeAvc3XTqL56W1CrjZzZXWKp/WT++XMmTRF4tkTR7HSDb/kVNtnCLgM
KRdcYKW+XgYBEHGcBUnbR6Sx4acQyZhlw7D7N3+w1EXGIeswRySONb3N4JWVTr8g
q7Bo9R4mAfInXJbA3HXuSvFlo0y9IZoV5EnEsHVRf8xFkwIPtI7MLpGdWk53fWtS
Za8WhkMukiisBgyUYvdQHwvg3hfpDK6IwxBQNRiQzRxYTzZzSjRRFwjITeybnCHf
t+qgOuwQqj/qrs9WGZojug==
`protect END_PROTECTED
