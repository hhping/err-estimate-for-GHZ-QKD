`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VoMUj15kiby3kctvPeNqVuheF/GFirURmjefSvKLBYjAI5X3LiAr5AmZi6ntBC10
3lDMIE8tdp6J05tvmSBZivEAir1BGe5j5W++YPWyDceEHC7MYiWwFbNKmZ+oPVmW
HUiVPJhNMvfOI2TDfQgQErp1xnzNY/4rbgP/e3mjmK2c5Ya8Gu/PbyQN1g33P4yr
SwEMd45ZY/TUGRDgig77TwQj/RL2HiJRJFLXqvSys2Qa3WpMksXsHGiIDoGlovOK
nTw/ZLaOubsXZ7U8z0Ech1AoJd3pMtOJfKZt6a1OpMjjGyLGKjnhpEkn1/N6ZNEW
csxxrMOuxb97swpBgYm//mtXQbbyBKYkpmsGNbGZCv4wQxh0MjJ7cn5qp/2X+13l
a/6lfkdp/Nx6Wv4p+QY93dqAInXgc/aGZIKRjYdfKjqdz6r0TDytzQ+nEw9axXdN
hJIukmdH6VXuX0utPkAyggviJtkAp8pzYxWoQHSH7ONIUY43xQCAQkq26G/E549X
GWcFZR1cp9GOkVwTHLX37VlOHbClPKTcVd398TZ4hz8AXTJNvru7wh73jFtEHyNV
xGTOQsbuwxYCdYS45A3fJdX9OxD35KYQul2R0cJkX+JdwyS4NnQ/ltRhB9B7MTHT
f90DZ1bd22X6fohqL31a8HLexbQPaopSv1ymOcBFb7VZaiE0dBeuQ9UtJiYHc8br
hMMdpynXWmOPE9Rbc7Ezhn62VND105V/XTVJiL608pITwgQv1PRGLDAiq1El/IRF
930DDuicmtqOYuQSDXBJxn7+UIUQcopKh86rcvgD1lqW9eiK63EVtf7QOXv5LttA
uzTn159aGOirCO2vm0TIjRWXULJew7U0rFzxVMOIBGzOfMoiDbY36qEOd8kO+Khx
Ghjk9w+R9Pc1DERmdjmSCspmea2Tq2zTohXZ1iSJp0v1IO4NtFxlzVjZ7rs35Tz+
m2f+LxZBouQiMsaktQoR7onuTFWN2HVupaikd6mg8uceX/AwwSKHbiqmK3qcDmrx
aG8I/3bbmDnydAKMSyXfFw74/8mGj4Fhve6DxMNjgtR2sZAV8TNjDwEo1HNlec0e
eZox3DdUmItZl/j2uV24Mtlb7FbH+uf2hxP/OLa78TBHdr6aELDiS8DgxWhqr8EA
stiPgiw0OJG0jJo18ggd65G6lv5YI6bYWgMw8er9TY3us+tjQJYumbppyOSEAOOz
fJYxSxYU60GpgcbgyqCRDFIOpudQ+oc6c9vfQAzgvj3eKrnNNr7AkXCmiGEdtV0d
+C3LPvMfNPOjyyq7D3Bbsjte+BLFztrrELrfvsa6B+SP60KYq1Bnw4uEPu9nqzWV
PQgouQp3qWuOsjRokQqGq3Urv9z9sf85ChcsTPc1BLHKDPEvKAstYKyE6vVHjmO9
vyoUkSN42qyaUvhcOWujbKWFcrd4a5dwuDrAi1SguKp6n4qIcwRDLI6IkMia6YZa
N+DMgye/GJ362rnx82mbZRwurTFaQPUkotdNVxlRtXNsF+oMJMnmEmsfmaO9HG5F
IR2kH/ZCAEnthg/S6dkEIQ==
`protect END_PROTECTED
